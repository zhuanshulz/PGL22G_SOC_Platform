`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AesBCkyoSerIjtXE6UCvjngh8AHUmz3zEMvyh+thSE9j0mw/bTvw94tqSOQAV/qH
1BNA1Iwx+Eu/KE9CclMDpq7rjvdDbYeIuxjUsDRwNbwdUoGxJ4PhNy3Q1lB5HY5S
Z3L67u0HKwrUgRd0iRm4yXZOcCX8WMG+yXEjlbef6RA86of3I+3NKhjGLpqnOWNL
KzvQNlC0ocAu7GU1iuiB8XEOL24zwZgJ+saPBJb315uUUidY6fQ5E7jsXvcGJe/W
IOw/8hShA9EMvUDIolJ+SN04eHSx6+4Uh6wT1LUN2YrqYSdPbO2xnSEO7aV55aE4
JoFxM79laBNKhL27JisOtTjFVhkmaHlTx3P6/0xIRyJnZdvPl86044+kQ/nhmj0V
o940eG6zjSzh3HT6nxpgUl1HKRFS19U4q2oCd1A6gEmaT40NkwclCPe+I5V2I+Vf
Ajw7Iue5tvP1ahn5neOptTv8XauL3NRsHFYSUVmZvhCThftozMI3JVqFX3S5+3j3
bJxBp9NvHBEp/qIN8Qe4oxsAWUDD3w9vtYE+JbKZ/QbGCBxmzpJoOo7iP7vqOL9J
B5EoSHJHYUpi7ZxwKZaQNEa3cNdm4f0AxoArg4FZNYqTzL1vNcdYDNapBPyCOuyJ
NnRIJ+w47Op3m4HEO9RzMgsQ8HmX1uYn5yc1tFSn/DWi2dNQN/o/HiLFYOmChBGb
gkB5M45Q6rb03bKQW+kRJQ==
`protect END_PROTECTED
