`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g4ySO6TxIvW4vw+50mt8ny6bfy8kC79u0KgAs25P4dWoyb0hd/v7VprNILqERNXv
MVsS1MslUBrHASDM2YKyrPyxp+ppMEHvpsuBph9KZR80Ydp67YPF59RgtfQ/c1sY
7sEeWf+kVbOhhlATsv1DGn8yEk6J+Wzk3eK7VE3JdZ0Rtbd7qTvU1IdJfjo8FML1
6N59uOIr5e1qWtPvQ3iDbbbfqhTiLu7hU/ltaA8EgKE53CQjqDqA4ihk0Tdb1a5V
a1uC7nLTrZhM5vIzg0oJ8Al111OCgFXqiQioy1BSPQHRFGglw+8peoO7Am/qCw19
ETJV68OlzbUPdv6BtJLFXlHt9+TIQ7uIBRf84pcbR0/HGL5tQ/fthYkdCSO1EwIj
uNxVZY/oM9ME0QaeWZvcUiijRDg4XSc9Wwz/9WBmPo+CXj2oWrR2sWRkgtrijFR+
4CLK9MMO49DdsaqepeQ8aQ==
`protect END_PROTECTED
