`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rm/nEs8jyINBTL6wzjtyxyP8nwvl2kGTa7V+FH6q8MAivGiaFdjG5M9MQYKANS7m
jzWfGRIPGW82C1VRlErJzEKkBOeCXmz03mnHKK2bV+TI2ryCTDORz7qndAQCrlla
2ehu5ikGm/BqxFxOBFmTGIHxjqRlsf72vcmDmW1HuwpFlKGtZF3oHHIZ5Ny5xE8w
Fd4tJAE0q10eC2aNxpN1qPgv+SNd2wG6jBJvgFYcHfquTcgqImdi4Q8whmVI9mcc
ZQeiw617xXkXcqjkY+RghScAJ+NnzmCZhOPVfaelPDyxTLvXuxPOQPzJHQ17nWOb
lKxT1bYgIFAeKA/M8KYvMtKYR2pXdSoFZVvtMvHG0vRsEEhufLXxl+VRE5dDQlH4
a+YseHoEsPVYBcUDdCR+UOXnS0rnSRCbWJjkiWHq02Mb8Q2qnxFxURLsOOi+f93/
CWEkcKoe1j4bm/cq6wCbIzYQ7aSA1t2sIzQxhRs1c07JoFWNpwzozDoo/yk6/mdy
PXdZnux/UIM8VLvp2/hVoET4phy0T14G6vNrROEnmKcHbT5vYqL20oOPL8OBwIzu
KgWaE7+FV3DDK022SMdmcqH0F9jtSvdtI0gA9TpsMLY9hGtfNdxEPS1gh+Cx7Rao
opI0fF/TAHVCyDsqQs2OLJMkmEHOVEz91FC4StjzjObbbuDJ1URuzTcW8+JTVWhP
bn9LuBY+LzOiuXASzsBbRiUdLqz3YQrxOo54jB5Ggr9Lt5cnyFQp3ZbJNO9y0O8d
kg2nKUEyVq7/8hXeehzL9DZS7+ZCICnVGA6yyz5c3iTzNUjmp4rhIleqs2AflLxF
1AOlYcqRp3VCVlZmXIGimHmBxFNSQ4Dt54HJ/sGYbdluv0s828CzOEr1gIRVMIY4
MDuZrCk2pJQ1WVdksPnn1kCzUh6ogaMSkKbwi9Zs/AOMVB4Xkzevt35RY6DQuM/p
8E477wCrbWRsKKGsJq1OXnb7rU4wv8k7+ZRZKgnlOgyStkAgRpg+mZnUR/P1YJ3Z
gcL/CCK8UVUn+CCPsLi3YFVXmzvVvjY+U0FW30Y5QAJaQgVA9IIlpSWh5OH8QcRw
`protect END_PROTECTED
