`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+lbU6gJLKyiqcXyHDgAFxMVQfV4h3bmKIHepvXU/6YlZBtIy/CdeDOiD2QU4UG/m
hX6bF38OUyxDPkJ7bE/EQ4PcnC36CgBPAQ7kzleDAv/fqIINMoD3mcflY1HpoKSn
ZBP4oFteLNesl8KBRUyD4r8iQ9aGeEqzyeIY8nIXSYuII0buhvGzpEAOntg17Vlj
DXQEtog6HLZjUfllLgIChOhwRx08RSP3fzSYslY3gV3Xf6r8AsaDfargsTIgahj7
xz7RT0Irlnb/I4lfDrnMVz5lWvjwHluCdDjUjRyp55IwAzq2WFne7iUcYE6JBd59
qMYUFwEA6M6fxI2/kyt2viCCqHWd2dRQrSdHbp6X/7W6q3TKeizHynbd6609qfpo
JT4V0gxIILBweSphHCNZkdXmKq9YawkGr2NO+Za17mo5nNMZkN6F/HQpXfc93fSx
F1TbMk0wgxMvre6jo7jNAJVVF/We3RFejFS/YSZsVsYFFlojwDjtTZcdwvzBkEjj
LDNbLFT5nCqb405YVQWPOF6YVru7FMrIz7YwRPitlNaXjwj20ef49ar8wM92rtWy
x5bJfhV1gWsdA3RZsaHrFIJ8UPgHMWRZGE9G+waAF/hW17jKo5QsMD4klrhaK9BG
7Rm/T48rj7vjImy6fBezca6owSCpMYQqOofwOhpgbqihOstrhR2doFpm/TfqMTw4
60K9plngxCF2TBsZ3Jv7hAjrKwY8P97XHDrwHFrtF6sQKdw+ueb9ofoTQ5FivGoh
ZKDZKyEKg0ClgxeVVqz+eyHFH3+DcoPZJEAG3IFxc7zkG0HkkwaJCLFhOXROog/O
hBEJ5ojHXwRNO6/sgEMJmBMvfwRbN6q1F07dFHpRWnDWaWe75ClYZ9THFw/T8BKy
YTXT20o8AQzTSY8AeoCE97YM0b6vfM4WzLGIGWzwODxI21GE4RHeJDlEuOhg/z2G
jb6rYOSox2j0T902DedmRrUd9wAsNNxLXTouSP9Wd9cP/vvebtJbFJxlMH//V4G/
CrQqOwIIomLAvjbKeixUXxPrOtiAhYSXF8lyPzvrZq3ndIemcW1yDPqRy9pMcIgY
ZBFLGQcZiTsmhcc0k34fyWKvaeyxP1HnKvK/RCN1DdDVZW/5ytOXb/VG8fHGtfZK
ZNBIdaQbJ3oWBPPnOS81GiWVJELsOQ6/h1mrG1Vckpm4NTDp9/BO1GcvGqB6q1F0
mVhIc3+q7xxp5nJvYRfvOoObSGiEbe4WmtpFWVOf4O1K2//ioh8MTzlFA1yugYG5
VE0q6JFUqg6+HAmDVoJ6Oo5YPgQksWv7sWJqeskawLWPGRTXOJajlUis3TQkEQen
CBvle2XvIXL6+z/hfFu/czQeiakdpFbzSzwDLc40y712t//ahG9ERsNWuB6bEiqT
ZlY/RbJ1y0Ishk6wJoOXIocAlbyn1M3ahhYushlAv/GcFTBk+uwGhe7G2w0d8JqF
VP9QaWv+kFKCLumdqWLDaZAqxRXoi2HJBI9Cz/ZWa2OrjlhrvtacaxT9WtM6vGPX
6rGCpw7LkrbMvtcxdyyVk7MbY1OVUzc6ryq3K8/1407CK2DVTcALeeAhuBr19H0P
7HDVb6zRz7IHBRXuwYbhV4n/3CAbXI+XCmy7m1gQc9HUt1zifH4rRTNyypYO95Qq
ZhUjIgcGPoQQgAC6mFXWmfRdIOPvEQi7lt4NzIiUzw7Rg0u0Sv00FHzaFdbDxRtN
5O82REpT6VLaiIzRuztbmqpn1HuGgzH+DBdovx+c7Slf8sl0TfT2nE8Om2SQNi2E
1cAfnkWt3TVr1JkSi5aZ/jXWI6aq8G5p4CdWJQVHp6A6MR3qx5U1M8Uf8YYOeas0
x1Qr3T2ngTOfAn0CAPIEHOVAtwfoFN21KO66CXaFpGgsWiwqkQoNR9Q/4LB0KzZ3
Ry1W9z/7uBlDSO+BFS23S0hDt+MIs2UQ0kRQgQ10u2jWE+JvOG0MEb9AJgVDkfDR
66SM44ERiHWgf8KNXV6rTZQploZsF5EUtgkOJiIjFrH5D2wzGuAO5Lg9SRirZmpr
wNxvDXv7kKsHGpw73i8knDNRaM2afb1LPS6pYJbvEBNy/Epcp8S9tpk4ruez2ur8
t9FYtYB/kCYVYHzfJWfYXGHQbL7sihH3GQsmn2oltK5MTxqDTvS29uTv1m3CpN3l
l80wfDgYdY2sH0gg5rFVFm+t6flhOnVSHQx/TV2xMw4rm81ReQnU4oVOu4kNp9Tx
PJqXW9Ez+C4s8LtDPkAzEku1EJvV7fy9h54eTmOYONixzQggV0LfGbNRIKvAIIgO
QKvk1EbVmSbq7izK0PGYadE9+QbsWdXunU0FArTYNtfy4sgVrQuHmt5chta5Hu8q
jvSUcG7LDPcqHSGg3To/BRgMJyNAjfdJaKDnrfSUw3Bn7Z1wBkDLJkuFT80nqSFb
B8NGCd+sGfuJzVOXMcGWriH8GdsFTgEz0avsQuaoGJy+bITyoUzSQ8T+QQFXc1UD
XsibZvUeROzOWo35PhHTDJVmC8gJySxHEGmH5J/QAhmpqSeADqUvLab/LHJ+liZl
oImeS1OHTBNUM7ZB4BMGN2OGuL3v1p9aQYMsO3j9YUBW1KEHrNq+K4n1RWJtTvWL
tg0Khtxe7gJgKPCyJbH/lzELvQ7Y1PSzeEU1/ssOueZKWrEW/Kpg8ccctV5tpBVP
V6FlEytJ1Nh5AnSSjRsxj0pYG0SuAvU8UA/M2MkUwzItm2Mfd5CQ8YBeIZQbXddg
bzgGQkVh7MzoZu2n5T3xd+JSgfrsg/sH8QyvwUFL7bMwxgAMfjsZ6NaEmm2tW95j
4dWu2UYGs4W3gHF1ukDdoKvSRdM3PAEOxCT3J0dFcw7/av/nu9HreNXOLZV7sYfX
Rk7Z9AqSFcc/xaoeF2ubXEFAFC6siF5OfaYlS73s5vvUkXdlR/AeaNcskiTvh/rx
thrux4e+5nY6D0MJLntwGx7hrPaXWyQCjWnkMzirlBTt1ysewGRHotvMvBh67KkR
8MYa6GRe5s/ivBSt0ELO6XP7OZbLA6R2u1buiY853cZLYB9aBm43uoFoEFQlhvAF
zHSCAG1LFY5LHdb6JTsddHQtOenJ1nR/ukK0ExZSDgqkXOCvbJWJy8i6kDyThGQk
3vQdBwHuNP3MXEQ1ftqYM7O1bpj/9wR1/kANWPoOuOv1y6Z3lcyCMJCZf45mmlX1
YwdtNstRWZ+BEL0rWRsVKCPPLO+WDey88WcRI91cfR4eehDwEghve+sCvXN3OkN7
qkGrcatcuHmGye1ga2qd/G8U60ay9/o6k18h9adsu51orOARt5+5tI3gWqAzCTCX
akTuN+KzKYa8T2Abq9MlEqu0/zEGtj9bOKBYM6CMuZcFYWK8erZU/wAsWOKkNJOw
f7EPQEsqcH+2uBg5g+psxz8D88+OPpNOpEMoIj7DOwxHqSGoEtJyXHyS1+cxdDAi
el8DAV3bTqi0eMo71LRfNNktqr1qfvTsncf3fwc/q2NY2vgglS7XwriWWblNlrSw
YjpP+sSn3M6eIs9RfdfjhOtPvXeI32cRTVH5pqLXb3pHdlXdsmmU1JFX68mg8H2J
Bh+FMrCD2YQ8xqb6YnoPCmrJApyzC5hOtz1vjOdlsEpUg7TNQhcA0wY3xcfDPyk9
h/d4H088Qi5Lux6qZfoZcUKuG4XU1u+0QA5WFOOYTIefuOqK+uiribSVtj0K37Xs
ZaM91uaqqJHClaSj8Zf0SJWjtoROQJUT6xDlbVmXAHSg2c/8iNsPFZfZNvRUSquW
RLBAL7h3BsJCOPozoyYVr0U69Opw/hwa3hb10lGz6BlsooHiORoY+RMdz9nboCNf
mVXORBtF07BwlHkto/65cOMs0B1vCUVD8F1u7+ZE1BH0y51VyiVsRXWJtFSEegUR
TCP0ra4+dQz8J4J7kcVsUSiklD0+ADGmI2vqiAMR8jAxZzJ0+8X2yvRmB6jtyiz2
yyUaxSQEimPf0lVvIEy57RL1I77lhV83JBQmhHzgXu4IDZ978P0hvr/WkSzxHTzN
CT0Zde8AIYQfsuprFtZydqBOSDlzuxlTL/8yWKown/LoY7EWtyQtJwfMBCnUOVS2
C9K5/5EMxtohIRmfo+NKe3IcWIa620EhpIU02bnSFrHc9Co6zYvOSd/9d4WqIZe/
XNd/fBJ2IFZeLN4pLxFupg2b26i1HjnhgombiEJj7sQ4SY/163PRdK3zOwJyL6Or
MNP6MgFRqzWPutFHglGheBDmavSkUwUE4Q1T4/sU2+KVLeIlixvDRf3cfV/9WBN1
55RYsqZfzg12cRoB14SfqE77LbXg1uQGg68QBIiWP4v3TC3sOfikmF+josAX9Xrw
14y1HXURVIGYFKMWw0xzdZ8wDhrB4tA0FLXnVchy7dS5A6bNuMGCOlryojtQkuNs
r5yakkogVA52CD065hZmt2M1L5LfScbwN0mL3OytMPVKCZTnUjDvS3hguGLsQ9YC
Mp+5d53mc0w+aYQ8KT5e8M5eDVGHRn0AYdlhY8H9xoAp8ei8UzNC+Tk3PeD7CseA
ucGUx9ZANaHcc2R61a7Nh3+wFTKBT7m/8zvujKtZFLWRKyBIVYaAeAhffvjHxCNg
Gn9awt1uLxnp/s2RNUB/0A1N8uDvv88V7QVlDXMXYysfEEycLEAPbsZg7SfPZDTu
lp5OlzW8t1YgbeRPfBkDG3fi2VFAkxUTJ7eg4VsNgRsvb2LVpqCdPhwqrwn97seZ
ewpAexwNawuSaYNvNObDhba66BJLzmFI9SYxpdCbboyKnLnE4WG7Mae27RxzOTxN
1wmtcdiutvWeIyUk1LEamWAVNzUthnAjtblBEb2Da4IOAGZhqq3J3XgRLWiNN3IY
oyCv5Ah2HCNuwTbueb3L153KeWYUcKrnKz5vFsWMRmVEjgQNH0dpz8JBD6CnTeSO
sJlY8hA0p+GZtfXeyHI4eAVAE5hyLtv5RUC3qHkMalUp9ir67u0Xe0RfKn/xh7uq
ySUclXuXejZGY9uiDh55+4EJ2hUkbmdcFaaotrcFSeZP9GLQZJk3oNnEsOAJxc15
cWTuRkIQ91bY0KUcAr2uxdFRioG0lUygjimf7m7BTFpwMCJ0KOH+E3lZHuUaXEx1
a1OYyzwcb68nFr5HPvI4hIhuNSlv+WSJtBZIzOluWEQyYtQZmAmvuePTGcX90VEK
szLdIGYAyMt44k9d1cn618ucNA1q1QUHnAQ2RO3HuYYt3yI80dVLK3zZhb6ASr2f
Hrf59I3+s7v2MOOKWzc1CH+XoJx1s9mHIpNqsHMbZalEgbIbtZnQJCesBNrRlRN/
TxKI0bhEcngNb+I+g1DuSED7OxTROWFk9vNqvMytaCOqO/e+l4xuYAbarJLKq/ws
VwCTaPkD77VT+bGZCWF4193oEjaY1hc0XgDCQDbFkjsfFidcd1ln3PFnFDqXH+V4
HpMT763A3UqdOVZnAKw8zndnZYYA6nrIgiF2NSvfLbdEcehdI5GBrzw9x6BLC81+
8+rY63WLosR/yRfSpfJ5ioCkSyKckY5XSrL+FE9v5BeJRRk6Oef0Y4yY7wn+YMF8
i8ePwdgtQT0bHe8e9yegf4dwZsYvhJrXVHoh/BMlMEv4kkcB66zNr7tVeZnTy3YL
5R+yDAz+iFtNOYfztlyIFqvv1oGZHjilisLTFI3KEE/YcjEIHVOCY6bdlesiMuic
el6HWOuAy1lDVUBdfLJPx6o5GkVV/TBrKNa40WTHiH6OEShq+pNjqbRwQpkywECX
pYmGyKsXyvazzgsdcSFnlA==
`protect END_PROTECTED
