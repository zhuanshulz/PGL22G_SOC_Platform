`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UIvhfv+HvwlE+yMRUb6OwAWrZrVTX0XFBnIHlawxSqv/RQAbUvlkdsuriRDy19Sn
huz0WWKBX7mwMo/NednEZRuIMUGTxL2i6IMH1X2jBn46Trx6K5UHPoZsUiydrbvL
hxlcuDjTAekkFxYYM87USrPFr0xx9fh5B+GljroLydxq6j71FSgLbhzIa+dwfka8
JZKC+VcpOjoSoSZoAy6BgqmMb2/4paGV1PmVKPIgiIgYGLQygGuyjxDwhT/QtmAi
H96cALgxjv8ub/9/5/ZnOoDdbpmCV0DRvKarEEWrivC5mk7GR+1j7kWQS6n/yF0l
FPcz9pQI2g5cwFeFeAvcO1FxoG+nKsHFYZ51ccsfNoh8Z3n3vVJ5VMANnNc0SrPF
lddpirxx6TJ6Jd+6bop3tu0L9dPzRm+0U2mFdUJQT1g2jnFCHa1lfgKbGiu1/rcw
HP4d9PzKkzo7eKbG0HaGFXTmUycNI3E3y/PFnCamnv9V2mbIt3WGZYSgf4g1UrRr
Limh3j2uklWh5TtLWuTMv+gwGSQX+JXEY78LuSNt+PLGp1GI7bx5UTewCWsjHCLL
JM/sNph0+lT16dncVixSUC9FR3LUtZVSvmcVOWlXx2n0R64aQnNdO8g0WxNcFQqh
drjqAhmLk2UtH6kStnPOr7cFqrsXtpdsGaB72fUP5IML9536XIiPe5opHgklu+wi
TCdRBaA4DILtr80oUVAPnDfZDroZtAh8LLifdyzu8lBCq7s+rSDaRM+TFR9aqn3Z
zRrZAiUfw7lfSxsXIN7VP0krvBnL7z3CbZWvAVypn78ts0zqNHHWAZWxd3E3xymk
+ztIMcv5bpyIqTc8Jjcgv2LqYIhvMEMedMWftQxv/8JU5mk6kJl44ih8/ns5HAML
ulpCZDB9iHSTnM5mxx2QVMp1s0rTLV9CNOclaIVD8gBdnnCMFrxm+4FzYJOl6wjg
jhmeZ+puHqPj4kT2oKAl37eJO+J9tlKUDpeW2n4rjje7s1uyA8zsmj8EtvXX6SHY
q3HMlWdXuxOVPTHlLYHlNPv3MgD/ygnqtN/ckPq358+piHgNE0kTFqhCXsFrNxhM
bwxYY//X6xgmLBmFQBCkZCFWySe+tNyAbAJEcD/KPktDzlesGTNn4IvVrri+BxzP
zLyP4SEo6IjgR2P0Bf4Kr/4Nx0e7dxcfc+U6q9pR90y8NN/kSq8axiAiS0HnP78d
uV1K2y5HnmKlP/aHwRFVLsAdmDv7BagyrCmFLWYu6wbR+Q+gsWrnoAtgXwpwa5Tl
545MqvQFJtJQklETbp3/MwEPpzAYcqWHX8/mNbpSD7XZy+gUN1wvKY+X8lsLGkOx
RHQvRDTDiMLWyGLQSIs6+Cdn5/pWPtR2x9bVKcNqupJmrOc5IfJ+tlowkqH7IDXN
iLXnLttqX8zwR10NWRd4Wgs7ugLmJjxLTHKKD8TRkW2C5vrMYH2ibkfI0jU0JOfs
zyKsrasVX6pW9U84bTsWqxiKIdqytTWb0Qzd9/TuiywnYQhx1obI4iuKGV29qY+w
647vNkZ5+6MRXHfY9DGM6ehc5z6OLOER6ds2omH9B7wGw+jF2uJpNKayyuGqZqWx
5iTYitt2tadtkgcRHFEB+1oU9OxAOVtU/qLrCv2sLDeB+TqDn/6d8HCXlNmcerXd
KEbFsbEaw3dqL3ZiS92fivxyqquMQMPAuhfAsHftgZYQujtPkhM8xeM9RLJ0Pkv3
E/HbUFd9iEOKpJV1I0sxmdI52i4zAE4Fby/5UjHyzymhMuQgVa6ymz4npsvbUh5w
P7ATZ1Y2Oif9Tmn5o0bSy2T8/gc6h7qokRQKhs8AVcO2Y7nQMKD9e3nVt/f53ft0
CzUSBRxt1PK+gF4cnaVHcTLhymeLd8E+LKE9Kqbuz4GWyXPm6i8CQ/RtlvZNeArL
xK80Y/Kvo0dqlez8J0GCYC0obc/RC+mBSUc4LIaT/2uu9YCpKGOkxdm6Wm2m2NJl
mHM6L86h+FWFsBlXfhscClWx7X7abkKwh1qWxgFlBuy/FRfS8rVS2dY6WK2AIYqW
XDwPtBQMctKqHk2JsLBElHCJ7S81jLsWUwzLC0upA1J+YyyFfM9jLAwedcu8RUTZ
jd7HIjSBAoYP5g272IWQEXhM5jPe4xealSK7ocmDA62ZKxDcB/kUvEHC1Lw7fSdB
iiAFSjcr5Uglt8RvBLCTE9jg5AvWxD5SKiUc7uFzBcH+oscRJp+E6zDS2QRznixy
eyVH92U7Y4az1Cc2CkLu9wu3bHbhuIdV29kBpVB5ma2VK1KS04qwCCTYMrZLsIFE
6n3wP5GlK3OeGkQn38RCxpD5wWBXuzEaXjcLg2aYFVFIl2WqrROktFEMQaQIaNB7
HxA0EqQPXKOkS7Hxjbs5cuPG1otw7MFE59bWzlT1QS2G2DNPhAVSjqSb34G0xjLi
NtwYdeExOqBr+ARUEiLXrkqs86c6ZnViULLw3reCAjeXvMyYiU5MKOukbPMG9qdJ
A5Rczb6tjVqb2p/0lb0GK4AlRbDxa0iYkHxR7QKoAR0=
`protect END_PROTECTED
