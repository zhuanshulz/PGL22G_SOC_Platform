`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AIYeBRtBJwfPhJMrgyCUZLj4GN3sUveNQGUKW3+48O/8ZjBU3omA86bW75wo/qAK
4OmD4M8GGk+l33lL/Tck8K0RuPqBswjYJIW8Bel5ivc4OYTVMVPwF3NDUE+aC51W
umheWyc4NWll6HaFZzbgv1HRX+BIo3O04o2GDuCD86howwwkAAaEiJKRKQnD8tiD
bS17AjA+Inrj6mOOrZXQkdviZszYFWoVVAh/W9+j3Yc5ddGkaePbVv8LTohuGlC2
6hycAc7DEe8S68DpG3rix2uovXXYp3zXT7CzPoZMqjIefzM/LoMjXQ4Zv2wqh89+
c8ahfjNH+ZM1/bKlBN2osvEmfS75L7ZdYyW/mprgkRmm1cF2ByeGkebnaM3oS7B/
kUalEar9QS+NmkdC1QZjvoP6+bgDctLWISVvPUAj7do=
`protect END_PROTECTED
