library verilog;
use verilog.vl_types.all;
entity V_ADC_E2 is
    generic(
        CREG_00H        : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        CREG_01H        : vl_logic_vector(15 downto 0) := (Hi1, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        CREG_02H        : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1);
        CREG_31H        : vl_logic_vector(13 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CREG_03H        : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CREG_04H        : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CREG_0AH        : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CREG_05H        : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CREG_06H        : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CREG_0CH        : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CREG_07H        : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CREG_08H        : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CREG_0EH        : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CREG_20H        : vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CREG_21H        : vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CREG_22H        : vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CREG_23H        : vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CREG_24H        : vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CREG_25H        : vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CREG_26H        : vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CREG_27H        : vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CREG_28H        : vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CREG_29H        : vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CREG_2AH        : vl_logic_vector(11 downto 0) := (Hi1, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0);
        CREG_2BH        : vl_logic_vector(11 downto 0) := (Hi1, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi0, Hi1, Hi1)
    );
    port(
        VA              : in     vl_logic_vector(1 downto 0);
        VAUX            : in     vl_logic_vector(31 downto 0);
        DCLK            : in     vl_logic;
        DADDR           : in     vl_logic_vector(7 downto 0);
        DEN             : in     vl_logic;
        SECEN           : in     vl_logic;
        DWE             : in     vl_logic;
        DI              : in     vl_logic_vector(15 downto 0);
        DO              : out    vl_logic_vector(15 downto 0);
        DRDY            : out    vl_logic;
        CONVST          : in     vl_logic;
        RST_N           : in     vl_logic;
        LOADSC_N        : in     vl_logic;
        OVER_TEMP       : out    vl_logic;
        LOGIC_DONE_A    : out    vl_logic;
        LOGIC_DONE_B    : out    vl_logic;
        ADC_CLK_OUT     : out    vl_logic;
        DMODIFIED       : out    vl_logic;
        ALARM           : out    vl_logic_vector(4 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of CREG_00H : constant is 2;
    attribute mti_svvh_generic_type of CREG_01H : constant is 2;
    attribute mti_svvh_generic_type of CREG_02H : constant is 2;
    attribute mti_svvh_generic_type of CREG_31H : constant is 2;
    attribute mti_svvh_generic_type of CREG_03H : constant is 2;
    attribute mti_svvh_generic_type of CREG_04H : constant is 2;
    attribute mti_svvh_generic_type of CREG_0AH : constant is 2;
    attribute mti_svvh_generic_type of CREG_05H : constant is 2;
    attribute mti_svvh_generic_type of CREG_06H : constant is 2;
    attribute mti_svvh_generic_type of CREG_0CH : constant is 2;
    attribute mti_svvh_generic_type of CREG_07H : constant is 2;
    attribute mti_svvh_generic_type of CREG_08H : constant is 2;
    attribute mti_svvh_generic_type of CREG_0EH : constant is 2;
    attribute mti_svvh_generic_type of CREG_20H : constant is 2;
    attribute mti_svvh_generic_type of CREG_21H : constant is 2;
    attribute mti_svvh_generic_type of CREG_22H : constant is 2;
    attribute mti_svvh_generic_type of CREG_23H : constant is 2;
    attribute mti_svvh_generic_type of CREG_24H : constant is 2;
    attribute mti_svvh_generic_type of CREG_25H : constant is 2;
    attribute mti_svvh_generic_type of CREG_26H : constant is 2;
    attribute mti_svvh_generic_type of CREG_27H : constant is 2;
    attribute mti_svvh_generic_type of CREG_28H : constant is 2;
    attribute mti_svvh_generic_type of CREG_29H : constant is 2;
    attribute mti_svvh_generic_type of CREG_2AH : constant is 2;
    attribute mti_svvh_generic_type of CREG_2BH : constant is 2;
end V_ADC_E2;
