`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vrbbqZzFjBMMy+9/B2LRs5uqHwy5nYYFj2ww9djLNNL9dJra/w1wJB7mFAgskBM6
0t3Otept7peTlpSzzc6YyL5y/RSIPKiLOq1P3PNBmFau7V636f/rqAaGrKWN5HzG
JbwkVpYu0rD7mzURuAQzuY0EGmA1DUa7yJ5H2JAk7QdZGGDvICjaE0V1bRMLpVKf
9562iC1ZUgPcevkpp/Q5R2eFYVjZQjTwvnEh9RHm6WT1ZvtZLnVt5+5PcQDYZMDu
4r846To0W8QA3zOmrJgSIH/P5jVielHdYaRhkBopMFtuEFhdYvy1gwisHzceGEiS
oyJQL8VHlpSvXrNNbr8iz6s4GThEDOSB4XX9i5XA6fl9DVFEXW+jaWwcgxN300js
TegMk96AqyGDJsL+FPqL/pNmhk53XNVe/YNmk5ty8LJY/JTBVTsKr4qXRY9QpwAf
7iev2WpQbkAuNBQqLEbfmQ08pEiDWtfS+Mfc9SJk6UWK0VhPg4BYjr+/o+J4Ds9W
EEHKKns9OZcmCO0BjM5cnvZgWLRObvkaLXqoH1xkyw8B3BfGyK94fvPqrbaT9C3+
hXsXI9pvYpuZbDI6M3T6bDWrTc8hZ5/95ZvZQub2Xn9DAlcUsawAG+HxB3mBRzwl
Vip6dxQXyHUkU3UAQXpO/1a+vPPFyjcxCasweNwsqZp4NB8n/LKuP47tQN9VKSUe
60qjk/KZPtD7Mr/Fjj0gJakJmhnKyMnsnjY4r43oas9SUqfbYYTS5MsiBXKo+eg8
A/6uccpZRKgF6OyDY2mIQV9usMyiF0tWjSUkU0uFGcjh/a39H9qhKBj8/M51v1mP
5Tr9xRZf+ThJvHllWbpMyvpQnQSTqhqI+fUP1VaAawIMkL5WFZ9llaltcgQXeGcm
+q0KK/YZRTZKGRjRT7ZKZ1ON2usZQqDfE5R66GGGbMsR7P7nNx+bNSFVQJS9uVF3
/PQEwK3hK+9/KUTKAlf0lKGBIereBu0goTnS7IUasrMVt03SKHcmIN/1ATamWUwD
eJkE4mNHrPeY1dDTDnSxPMMXr3ihz1BCgZVGROEXjK1YLHhLqWbOfmczG1it26UL
Bj2F0sP8gdAxC3qbyc/tg2TV/2MM425faiutPUSLLuhr9iOeMma156kL+b3XWJZn
Nn9ZxjA40rklrHN9PcCPIR/pGR0stKXbaWqfydq3MAfMzsfxe33ijd15pvET/R7P
yrQMd9/u1mHYcrqWITiUBxs/9G8ntWgDNzuafJvGRsJ1F7Hd8Jl2iXag6RAeY5pF
r9iIPKVLXwsOJt31ke5S6Rv9eLF8SmVowy08bxnZAeY=
`protect END_PROTECTED
