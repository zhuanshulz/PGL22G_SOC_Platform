`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c0o9cYZyGRfATOyHbkVPcDkR/AXZKzz5z6I2wxa91or9FzPdDqKiHx+MHXNcwox0
Edblmqt0X74li5V9sy8Ze46lU3HBC3VB2AG8EA3z5J+bo/pWLytpR006juWLo5ao
qm6xy5RqkNBd9YAUnmnRFgFPdYV5TyZ3hnocHAhpfJVVZw85GZJ3aQCZUbk9wbWP
CabLRypwsld9DwKILQtlCYdnJFHxyPwNJZqYQMFl+607+1nNlSWKmDmSEahp6ZPV
WASCmYs123RhzSDlXGjtfXf6qVCu+mBwFuIEopxpC5xMk4BkKs32oHw0cld7oeRf
Vox67Iv7oF6L9NoVo9PGlb+1BbbaXDpy4LHcySW+NVVXrxV/coB1XoPtIFyuuKNf
nJlIjhUeebgRkqfT+ZySX+vOfp95w+uQ5xgrgCcIqSoEDM2OerJScq8BsmKRPH89
/Als6rJutmj1kRpXsLGPF+NQkE2SBv6PWJukAjQqp7dusRQkEFsyKHCaMYxGvZWQ
mPyLvJfhrgudfcPOdxA5YjSznE3Ak5RKPndMuGndFhoiNEr2XPraaivx9aulNgKj
tipmEfmZv0qFPu7yf0mXgnaCPzRQMJLXD9lRRuC0IM7z4oR+RCHAVobBRAm5jwjo
9zr/b7t2rRSY3JKlwKVsuAHX3u6aSjS5CAwk9H3o3VYc5MwkoLBRtrX1COeanvRN
wp44s+7HIifBqLGpnwGW/VzjoVu1H34Pzt+lYYmai6BG/pW99o5/d5t3BUSHJUP6
9c691SbVsjlX/1Ox2UxMETQ85w6G6bfl0vu5AUS9Wo6cOigVo5++p/EIx309/Tuv
cz7ZozVNC3ZsM+2trGJsG15Ul4y0XQZgw3QYOBccFbNv3HgmX/ZkxalhspyZnaBU
YYrQwohBGoerEy8vBJDU8yspsteIzN7Lu84WPcNr4fp26iwfxF2Vq8BnXo6t6vCV
9LWNaVtL1wLg28xqIM6c9DnQego9d6yXILPf1BURMxiSkGPfUt/Qb+nbnBpmoLiA
OPeU5NNamzQiBy26cHRFvur63iWUdoezHxcsZbdyAv6ej1wG1OXSQavtrCfDUFY3
Mo9xr3rK+gHKkVoMZj0u6y7ix/487jQhJS0VJNWKMJAMa4yW1QqmxVP0Ot5hTj9J
2cQwmyXftcOSyzTPqAwxN0jZjC6KsPG8/qLg0Y1mdUC2/7JJfAVuoSP8pbu/9Z1y
DF8tEbgHeZd4BgAgCAsVJnN8SvDx0xrX4JCxPYlIJUmyoo9Vsmff0Iq45RuZdsIh
x8Wr2/Weptg8mBBxP/vDzN+YErbyJQLf04X/+vCUUDEcwjU9OWNFIhf5tZvIwOr9
dd8KzYykhT3a7zsVydOf2quX3MHnV8uphQl5gfnFEcXMoTy2tHGCcK+vUYylnNPb
G0G/6V5MLBRra21pz3LvkfZ2zz1hjk2ZIIG8IhxiL1H8w+S7gSASPA5KDzkNUZ7T
NuS3870AGdvRJdnd+GTB8kV5Ljub7a+81xetwZBzir0=
`protect END_PROTECTED
