`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7ng61vYuYtupEO86o4cHu/gFzFFtZgJ0ZfP9GBkhzJVYa3ij9Da+x/Sg8dZIoccw
TGNy0kjoMRO+VZaSg30cwjSksMITONdUeXsNojI6gEmjVQxqyhIxwZ9rK8VIU8Qm
vf+58BgMIDwuClVrP+Bq5JupCy3HfD+bPxGps95JF0L1Myal4gyhaTASzjtT0JTO
i6mWBalhvJzdiqAMwMAYThSXCOkmRHX8Gv7da32Jm86DjPHJwIYMpUxdMqKI0yLz
/Em8obqPYf0xBUvMdm3jpt1BlbwAz3TV3vbcskZBYLJC7dTTnX5UPEdQieaj/yg1
/ni/3EcMz3zAa05X+64UnV80MEapbUajscanupv893OTbG/xnOd4uvrq/pmJrlSC
K4UibEoHrsH/10reDFJ7+g==
`protect END_PROTECTED
