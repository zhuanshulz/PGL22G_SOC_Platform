`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f72wtDQ4rLCDNKw25ISZfRlwvhAtPCFCdbjveUYaiFhXcV0Pxi2zW0WLBZKeXwv1
tZx5Bx+9dA5kYeveC1gE2SyvccK20fSnDgSvPxv39ZB6VraOKQCKAOgRD4U2HJep
aEgfaKbn9bnkaAgXITEk208rnBhOKEBT4SRcuglKd2qVSWXBymq133IRKMCfiz6h
zmmKbnS/0NcBSgPz7eDL4t8pMt4wbmv5WXNf4bPN3J8QRnb/iOIFgqBjxhiAKcPl
OXGa50ShsOhl/gFyQGMjXzdfuu2vLYDppsOXSb7IIwJO3EiF2slzU0cztD3hE7Ep
gMnt+kVjQpuPf2vAxB/bDbGBm2Q5sKEzj0E+2wOamqfXS0IjS8n86lnuEpgpm+gg
nKt9+RX0C/TmmlNQf1hXMnBIiTNFnRtpVDpEz9J9FSsKXrr7Goo0SZ0sTZRzl6gc
9eBzqTuT2zyhmc0ahnQ8VObwiSnMqKlRUf/plna7sdY=
`protect END_PROTECTED
