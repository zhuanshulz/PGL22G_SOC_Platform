`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tQUGwGH/RQDiBpBdeI3ZvsWATg32jEGDYzwOu804JD2p3J7Uc6T1yR063dq2XcNi
HUztS2G3bMB0rujr1oLCoJjw8xWLNOYm2dNDA65evhQPfH0CmRMGRB7VY437S4Iu
cGC8ThBlbTg3rslK8VQKbR+TKljXn2K34tB1YD4nr0mJeHjdkXLEQ1vls4E0dIBe
P2kFd2NK9KuO+HcIWd23n6nSxkway0LTSryLxADRl8+6rwE3S6jwGrDRha5U4TVI
jG9G5oEcK17oaP8gXSkyC/IsJ6/N6V9ByP7pZ1l7GMi12Rqaf6h74cp6vpPVbAlP
Ha1RqIjbdcNaq5CHbIAxXJTDZ7pNBmk/E7vTf1fLE1oleZh/0HUn7konss+ZVtZB
2ujxSIX4m82OelczPbOrtT14/8DaghJHw4ueQ8g7+ZZRQLBPwhM6UbqN2agdn2UB
N2Zhdsee/1VbsV1ZSkWydeoDS0GGjEVpCwy0WtoZbfwWSpYoLbUG8rtyD/beSzH0
iYYUWYUhMOPOKLiiVM/M/Y5lrfyy54EwTNtl1z0GJH1wIuwTsRAHcthYHtEHIJWe
wiBXRZzv3koSDCgbXhGgtZczCQR5bLhMp2SJxQvgJ+U/oIoBMfkRcCQ4lDntZV+H
M7a45Wqdnfcmp6FZ569TEXcODtc0GOwP2YoHHhxZ5xkhxyYue5yBYATVLCoh5B1W
mBpz7FxKsI70Q39nWJSGCLyq5k+V5zinh/o4JsJIG+k=
`protect END_PROTECTED
