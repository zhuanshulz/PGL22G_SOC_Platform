`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XWGzYOhu5ZkXxsW6M/mwcZ42A7WHNH3y4uIEYKgTQcpzaAroJ+kq7Oe+N+JzD4+9
I5lpTdo00lhMo9+8E2ATNKSa8hD5EKBNVMZC5tBnCUPIaDdEIUZLAqWkuNsVfoRl
CZ+D7Nlpy/wT3eNFYlI923S6otwDzW2nNt56+8GSziwpzKPn9NSveG/ZhBpvVHl+
zd/ARxiuTjIeiO+xnCLpMEvLHRZ3sKiQlpiMfWjSFBOldnRGExUZbzrjn05tQmel
/LG8HXIUVfbk7OFdtelrNCB6rdzNERdl56uzn3ofiTSsXWRYrt+aGizdlWQFtSAL
4FRAfRd9+CufpKAA/wRk5W2SvQut1Mnbt65S3KKCfgtjNZ4E5FOUr6pepEJzXdVs
+jeCYLyC7LmQX+U+IiTL8GTJJYDqGluarOlOMyzNcWtRcRBHLVcdS4Jx+jWydPcB
H/JeM4vacY46fk+cVaJs9MJ/wkV2RWy8gLVJZ+WbpaEOhkXX6GOtPKmjxPIl94PO
E2a4LEpPzaq8i9IObTQMfg==
`protect END_PROTECTED
