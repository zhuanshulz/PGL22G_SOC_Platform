`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AwTdRqOFB5AZzPsB5OdUCdqDNi+yXwLoTvMStJmluyWZJlXZJ2huK7y/MztBt6PT
yADzcpYzgoZOCsYuoVXDBa6oPXmpuaXYvLGsp6anuczi3jn8dn0HRLKFtRELsdHT
aZW5Y/U4g1iA+C5tRHVLrppz3xvlU4y+AqCqBDAgBP8vwBxg+iSvNBsUPOJbNr+8
PzhtD568edp760KUfEWZEFeUDSQHAFWp8a0PzU/uU6RBisncqbOP2352cxtqkk9y
up055jPOyHm/aQefJEZ774LnTl7yyDNHOtLSdsqEnnMEx80xIKjY7lM0w0d9I//3
i2Cw2wIB4ylpYsoIajfe2ZbBGS/y4L/+naQkaYult8xyXU3/lu6JKQBnQQdCE0Q5
B7gUfz8qJqUZ8TMoGw2Vtsd6+ENL9NKXlvwq83cAYTCxdGTrsg4D1CkU+6WTRLwx
0FrnGfnSvOIvgtxg7O2uFpqqtPqMCosUuy+gXeaAik3YyohZhuRo0POA/zCUf58w
eXoQo8D6/q6nQs06Rp0ApQItQOVTxPtkGGC020bhDhCPZ5EYbm2jgkVOiXlqlkgm
cCd8iK2eLkE+buDg0KiNVg==
`protect END_PROTECTED
