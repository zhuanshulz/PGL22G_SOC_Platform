`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gpKSz9cEm5YRYwE9YXBed4gr62GhbUfsfhwfeUfWGo2UhNm+j7PBJ7t0J52xCfEO
Nx26NpyXi0w10BPRHCSDrDN69Ux/Ep3/bCPcyJKFnWEe53zgqYS99Tklp5VafEM2
PlIoAFaa9JXXmlSjUSfUHoPeFMOxcnsfAyG3wTvCA7jZeQPrwVNHtc9b8vdX68qj
EvKgo5mBY++1x/q9MIJ45Qm8A3tB4amaC/79KXDqVwjN4HeZeCvNfxn25IWRhN1/
8hDa7HpIAsL7/6vc02EHTA==
`protect END_PROTECTED
