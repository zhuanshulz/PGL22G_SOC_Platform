`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MiRCs08A7UiLss7s3HFOAOhtt/CvIkviE8rRaAoiK6FjXKW0SGCe9iHKaI8fvfcK
7tIsRtpXlBY0gu20l0Yp+o7ZjP6H5L+pyybje3jajbRJ7YMDrtJ1yHbIEpOhEQ/+
93lV64sUkIg3bTgT06kxUk15xsCDu1SCSOc00TH5iB5um2uAxkQR5HQNngK3ZxFo
BISMYnIife4Dr0Is9G5R2GrQzv8YDFo2V8agUD1CXcTbP5dL9Bgj7QxpvutmwPIV
Dz53tsPup9jJK7sTiDWJyDPjFJsaYAKpG2RjSdKKshYNadnWI+uTUbdF3dJFFFBZ
iBkDdyvQGK9r7FyalXtbh0MFl8AOvoT/CBuLlem7Oy5gGcIAPA8fytASLdCK7xFB
wQfLhrRWwBwUDPtd/eSh9IaMxa8jSEhoiSqHxeybj0ErB0o850SxAvrmv9d3pxAm
EXMcvHyKoQLW9DL8fhkWMOTMZV1+SpbD6UoE70moQ5eE6p9HO8phTiQDr1iYUcbL
Xh8phR2Lo8f/WEynY6BBne87t5aHjTOch1l7nLmgROu5r4J6X6ETgXhoqRGCWYUZ
Nsb0dgFOarBjwcn+z/gqU5QJpITnxBORb4cmpl5CSIdruFNL/Fi5piv4Nt0Y8ptR
08cPCAPGGuY5dXyBZoh4JR22yDygKuPx1wARGytveHO2r/sKInwoa1WLvMPbo7Q+
xbJ7/UztM5RfAZ6a4lUya/Oc2abDKLUoQZ0auQLsvTWv3Z8Z4O7Oi24/xJCPdTsv
lsCCFXUEqMIiQMkRwLVgzXF2tjk9/n2e+QXAtM+2vO5fu4nhTfzQ8/PZWka6dJqc
ci5E7aMz90qs+D43jcPKwKJbhSXL6P/E88kYHAWUbap81DDyCJjDdjut2o+tqF1o
9x4Gs64M2yZcRDlCauxCh1XNuXxXBPZp7z4XmPM10KLQwWHjibJh7oAN5prcFXMY
QnEAaP8hFkf/hQtRh+0cFaL1krGlbDunCngHMoWlfR0eqkFCClyBb7+uosrSsJ/m
PoBwUt5P5OviBf2CKitZKbJ/CdJLdvF2EzV0AhWda0eLXhZmxV5ljjgalP1NRNdb
I+mMF9TKxI4bVj8PTeUExzLWV0visM/Pu2T/+D0PXeQEj3VQFp8yZfQ/w9UuE52X
rsxZcG3SnmoMjayDW1W8L+jwTsSh9LSwsUAeI4ES1TYaL1ixmxH5EhZ6p0tSThTC
teNMpsobNiTIIeExVMKFgVOt7X6y+c7IJFBObL/qW+JnNtei+1xR814kHbBHvU1Z
AMaVsnvYPWY3K3CDUN/FctX1buJUq3F5L82WW5qIxhCwBzD5DtbpTkZ6xFsYf1JY
+y6uX69oFYN5aCKT+Y8SEHpTNQV6Mdokj9mzBkx3NY37HM1jKS1aV+mHf4jmC4Qz
WQlUpb4Qv23Y9hQnqaNEE5YFrLdcTzwlEVCRVk/LhI4JVbgrDgiHbURXDhFsP5lh
val05LXIpjgJ2eXFLRQ/Se3boSpI3udS7C7wiCLwMYhAka7zjy/LzSYYqVK54KOC
HAWldCGrhMFa+eDdShdDAWgc28sInih251CqPfZOQ5pxlC4sNn3ctmKtKNaxQvLX
xSDxrLy4drRBd/QOlMt+nPx51Vs3uc/9dbjwsDdgLKx77NR5nqujdMIqKuxDFfM+
y/28wPRx0RSaxQggrcQdQMQB7UL1RmnvEY1EkdcXYaz0YsfUVtf6F50u4G+b/hx3
YapbfLeYyLMa/0kUZ9s2V2k0thj9WGBg7gEQnYR743cLWllvoeMQEq/K+ZVcIE6M
jOUMJCGsCm/hyq6mnX84wbCtMbZ2E6/V69Kj0tj5NBTrCChsBat/ff3yNe/xY4RA
v+ztkHpp9plRay+qXosUPwPD3AcE9ifLW3VA/iSJ6jj2MyBlsy/dDgrd8l/PgIKF
tVRJwGdiUha/2Xf7iiBf3+mzOJ1ifaVoPK0NFeAumRjkTn1a3yYSBShIZlSbnNuR
1SBvDt64DWJ6c3y/+7tbV3OIVH3YsoTv1qUrzIYVHbAuymfIc/nE7mh/awZfXn4k
nmkqhCxI1Y4P2rpgcsOh3lvXXAZGCaO5md+a96XGVt78NVu5f6N/pN2LaONh92uw
EyaBD2t86gR/7YRHPV2U9jLrBGR0OJvzukCFQrS5D1eQj1JdhYP9uzQICzTL+GbC
xB1G5wzZunF/gACUe5f3arz+HNMj18p3P3Xban+kHMPSZw9hrt0CKmHMFKqXrOy3
JWp6zDdoqBz7eBvla2ibiPz60tty8jkJVAGMZbOQO9G0nIz1qqUoZAvuYgwFPe/e
aaUDZbis8lxghO30IVZwU3DKYLPheRW8NkCYk6rYJqJmJM9KFU6e8sLydAEpWyX3
Vp/KeOIi1hBwQK+EiViUMu6lBHpY/WMWeC/nwXzRecEwI4nyRASw2xA5zqVi6fmf
96EiDlZZwec23WYmaeiTNdLF/4MtiEnhyetdocu4n2eg5UBlz3cAHDVkN8H+8DtJ
6fguzwPwBYOf/YKWTGltH4tVt2CY9LbnCvgNU3RWPTbl9Fbk5JrrAOtV3Fhe+prn
rERPvDb5Ca0PaTwsXNh5wduA4Tf/Ctp0cPlWtyrm8UyQbyTXw65bIPpbLJazbwCv
yFrz9jVV2ktU2DC+x3E2SJ0v7LuOf8WUtqDQlyLae7yay5rdunzCWK4q2wtfpMEc
6yKrsc2mo40+5YA1CLfsyN6fp4dVuoAxAYy5IQ5d4ArZMK7tFsZ/KudhmUKt/N45
u+jdQpTwVZfxUkmzjGNHvMKcVZCUn1N40jmZY5zOzS0/+JQr8/0in91SPjEsWgpq
UrDZdeMzI/9XRbrPV54fJqV0TwfpNG6S6d0kPR9vV96xUOgygic2rpwt8StydW2Z
8Usv2rBBERScDbV2SycNMEOYBnkpCgK5ebfozSHa0ipEOyD6Qm1CDnvwTlNDhzXe
ykY5QUQ9iVsRTwIJO2Lttu2KGutQrAxeKz3eyZrdcn0Qwt4+w987hdJlthV6wZVj
GvssXat6ik/QYp7E7RZJn9m71fe3k9Y2ojNQSIQmv7eR940pNSp9greaogMqUf8c
F9de5AsWPs5QuUlzFrd8jqUmcVJQaEbN6uVCFGBc6ZyO1bgu2oDj5MQ3h+RAsWR8
85ObB/VsAC7JkPpwy3/1/w1QlHHtFLsyhrHSHs10LjPZ6PCY/CtpSzG/WtgAANqQ
wF4J0+SAUQdfRAuQvma9h4Vg2RtzfQVDViA959hEau5/egep+8bxqNU0yPO2bEY+
iAnjrbK6gFoWkv12c0LaZDzgrIbbNWqWaIX+JAxq8/9Q62CDsr2jhOoON/aT9krP
fBBLnWasJtlgs7tUSy1Tx1LZyhhaHnnX6ufTnYh+BDY1XWbBeqZRcwqx+5iBy64w
xM9UytC6LrdhticJWMQeg7d0rVHV+5cbCHcjikZtfRMaxMIV19vMea17XBljNG+V
ExZ6B6rLk/tje4RxMX553sspVPXau1vTLV/6zOJu39IGhGxKL9F0sH0fhCQ5RzM7
sO1VychfPOFgQTzy/TJaSaqe+Zg4ZTDmiMKVjSctkjESMj9DKyZ4/LSVEfR4+fzG
wd7aoYNFZNcTVReASKf5+tO/qUdzDKPtl5D4t8F/2Ury1UcXmw8gSLf5mIJPljBb
WplW8awph9UvtEO0Ipz2gbq26zpQOGOxgfhP7hozStguH8un6k4rMYGYjHVi9C/Z
lRyyWlsOdz7o3mPf534UOyEvkIGUMcBMID8vJaKubMg/Hbi0jfabd0LzBPm1gXCd
WofM+c/NPh+eOFY4o99dVCHyWf9/1WLzuaWgbybl80ViSIdnIVMEP04egT2wU8OO
U+iPg6PDXTr9lTDM2L399cP9hQpLoH+NHMkVGNMLWwWgAWAj0jxN2XYF2n0fSocg
UsBpkFC94aDZz6YsviY99wJuUH4lmV76YVlODmk4dIYPZUDUHGeOY4z/yJoN5nI6
87J4HvIi9+aBI5rPGt+Zw605HlL1OT9NuqbVqq1fAcPM7zV1iHvQMspgJvxCZ2CW
KWjxphgwNpVOEEjGSOPnP5WI6TQI+iLqHkGOeUjOwCC91c5mOWg1mM4bEqJ79YHl
D9kro3s4+qiScX8dIlKAsxzheqpmRO3SK01PXjbrjINW75QaVsU4LYcNhtGW/nSv
mMf+A7wFudzrUmKlWEEjVt9BzyQDzhDcwbhPpicwn8oZ2u7jr59R8RXQI/ClqeDC
tCoUmUDKaYz2JF/WiuAsWKAqFSVx0oIEhm2buahQWtLYNCj6iOkY5zvCgPxjAWAu
43UssXcK0gwj7a6u2qOxCyYJpP++Mh54y/m67jC4V9g6/HeL1Av9mRgG8YElh2sL
XE+xhL1cCtRphFKRexJC90mj9xhnbpjm2M5DYhTbtbHk8uGUx7qHS746D2oOf3pV
6HdlR6QejtUs4WdtoUY2qBD4HeYp2e/sLrb15FFSby09X1JFuNqVu1qvo7IFJ6ye
KsRLc86tT5qNZIVo8EbBTPH4B7Y/l0XPB0r1Ra4EecpUZDjDUW4wghWIhmaDjLy7
NryK/tSHPVFSf4a5lmofEA053NrZ6zm9LM8ml0OAUIy6hw34mjKOHQbiTfl1PcRt
+oGwYeKDnf8tR9JC6VbYQIWZcsHfCNrdnESZVyX+ox8ji+8CrosA6WDFOESmRG1k
0VjIVxEnq9OWNW4RXzZGN3m0rD9wvcBFTqT9TgvEJF/W3CSbMXaztMOQL8irDZE9
CJIjynMYVT0qeU/H+F4n3q5KsCNJNP+t8pv2UD6b+kMJ5ihspOYXs3bmqB1vM7OX
yAia1ZbfF/9YSsZlmcNRq4X7Rnx631Ubto68K1zdAO4UVjRMHQ0gObWFj4ccEv7U
C5RBJY1n/zfmZvTU3K2GxRpQv72Ik/YDAIpRcmnK1GTTdRVfVhss4srDrPyfhHHk
Of8gY5YkkhgL2qIpZKNaO5GDG+zMz+rz83gVvcky+LHsyq56XAyx9N7nMDIE4yl8
HvgNr7OYYexvZwfA4ZO3aS+KDxfH/3eTiZZ58f3AC5kKk2DTqmtN96kGaVaYneDv
xy8OTqEyigamF0wwdHzY86FUj+dqnoYIBIwpZQcpD20ycWgf68qtjUO0fXtxSJm7
BenKy+M3CFqwc+v7KvDq1FocKghdpkZr265cEmlaHOEqFSWnrAwJqe1iWupVAFOe
ONUJG7UQqSoAVzHYZQ4Jly0jJx2f0kASWCdJ8jis41t+yUdPam6u6XNuoLfDRtEX
gyF0KCBOSmK5sN5ADNhNvCJ+Q90nyKsV0ENwd+fIVeAKYTeQGhMV4WX1Ez8rHmQQ
D87hqpVoyQGyquMurUNRoMdlcbiGD3JdmvPTbsgPbkch2ikj27DK7U8W3rcv+A5x
2Vc6ojoAOlZ7nuo/qAtaFPIuApMqqDwrltTQz6bwyCMIIheLOoJwBNGjnK+kby8R
ocA7u9Y5EszR7Q03dKIkEVp3f58r8ndA7SNZbnqP3WMf6/H88CHgEne4cMuzdm9u
fnazQI/P1rBjiGZaieXkavC0C97lr7ekZwd4sIkVYd83Q+AE7uf+NoKpSr9C5xs+
GyBwfGzFMw7lISMDxOdCHxnbFu8wQQxQmlhup7yUimAs/WsG9nsq54JHyrz1ypMe
42FC3Kl3o3APb0yaO67hDv6damiZJynuobl3QwuuZqYlS8z59g1MuXKqXcVPFbCo
UhnawSuALVvdK4qLbbHyrYj4fXnA9UDFzgZwkdK+2AKujw5EO7uNbR5Y/YApyyem
fUVpfZaghUQGoYpj9UktD/XgG9GxMQ92o2H0Zw9Wzi+fyHC5foFfT4/BYaKg/Ly3
cv+eirUIXD6MicsoE2LwVhfjL0dBKdpAC7Ht8EcuZkl7Z5QChh0yiu03CHzlRq7b
Z+aMru4QKVQk7vvbfAMfEAXZ6RSYLOyVN6vhrAxdIO1QRBU0DSjfJLBV+TaFRlSs
2slFZDJvF0Fkhap0CJtmmYUxA9Pnqy1cf8jJRiy5TqqmPMDYIgS0jjpysYSXkOXj
D7lz0d+ISMaUHKboh0DOxYltIwsx/DfLaPU9cdFwvKz/x0dRtV8bjovvpS707K07
lZ5Jl8NaBBLL9z52VXjR7IIOVJ5vw0pBQJRa+dPiILoQ7Q4IEg8ZOobC80NWzC+5
xiX4srCkHjB6ieQRTvfwDVi5G+sDtLUv438QjGY11C6XnDBCcVbq1swhQbbuxoO2
Sp4A6tsOoxlcL0NOIOF2/rIj7QNCprsa7nJ+sm+YaXc10p7qK69z5r2N4pIsBAeS
Os/UWO7pbRQwPqcil2tdTktWjM9a6I4imvVlw/PzizsXoJvTiDCVCjOiekYnOGQ6
zxpfsn9dXu+MYdZDZgs45qkwUHqOk8XzEJ2o4hmhW2VY1zPFzN6b8J/Lg8L6sme2
+6XD1ggtlHerTkyI1effLwWaWBSFu/iaJ+gNUchLVJrzdyd6yxEORD3IzG0jHVT5
4sL6i9c+DdUzZaorVsIBgJHo9eEMav2qokPGqObyF2OHmvQl7H+gdyowmuRAtwvr
V+3joBpm5PwMU0MAmD/bwW13+DF1eQOmxZM+9+mhnbw5tRAwKOKkrSuM5ALahzav
bsn+zydEX5gZRkbDz+t7DqHqU8ZpN8tGrfLKjyG6X8+f4qg+YwgMZDTazSgfR4vJ
PkAsjMKvBCI0EONVWnMaM6GidiiPUwvItU2HjHkFcieVznPy3q58PIbDjMWelpfl
4CUscFfW98wzO+EFRaIXstBdS6sPO+hmNziB3GKtScO5JViHfacxpua9Kem1E1qO
ltuEHpCPKph9wgTxMe4GV9E1ZOott4AkczoseCcso2G7YoJnxHbLkhoKpaUsHOe3
pCnCLid00eyed4j2rArQQAhUjmxP8ns+Vu+qnHkwEV/2qTzzncJDhQId7acgcKoe
u9hPcSZYf+8csHlM4vlaQHOd5tPpnttRSmKHrsLmoxxk0eF8fuo8p6HDA3Mr6nGC
5UHIxjHFrNpNPL4/o5UN8IVZDAdzUeRKjwR9G7RnTygdGW68lwU2Dsrf7kFaBgqZ
KJG6OJUAUzCmMVoOWslHz2MVnDypQPd10+20jvb1q9rAeY09BO1klyVhfoKhSZKk
5Sw/wmKecoYeWpwEewCZ6e/4KptqyxPblrEPgQb1VtQ0lw0bUJw1LX3foeLXzfqb
Ge+u/8SSnlPfEPtAZHF6c3zPblpwBtCJn8jj310X6Z6wVUcijnRlmzSd1/JMTTrl
bo7P1zUVTSMhS+aHpJrtJ/fOyq2YHtepzrnZL5nrpYQ7dTC7fUokdeuqYoa0g4w0
DBgx7+CJDw8/treBv1lzI2mSBFI+KCQRw3Df1c8d2L6ZQZss4UZUXd5q7+mqpN6L
QsM4wPb3UbWQasXwShn104DInnZTtfo2xE8lBYVJL7glFJ7U/eTCyLgiKH8FmAbb
jcNtEOjLr8Ogj342KUwBTdQp0rMqQwmuMZH3SR36tkjwGA7NCRN8J1uen/EANSzM
vunSR1RfABtt90bvnqHWcTTud93wrtN0ml0IUVGjynWUc19rCRPKa9dvKkR8lqTM
d5n0gSu74p2PEiRNQO04jKWO5BVKBBA32jpr8lN8qULk6jAYRK92I37fsGNAgLy3
UNaxgloYfI4lvdz1ASE1Arf5lK8nDIscZj5nmRh+Rh/ytIiCV3AQHNxwA23vWhlz
fi7t0Rsu5l3PGvgv6ZOy0eTywcGuRoUOlfp0XTa4tgLu2bKQgCpGI7m8nbmFWFRC
GINzl9WoObXsUvNfy9E27QDrZi62tBXHbAflRP/0GtCq7jEcfFWQB9CxXxfF2AMw
fSpsKfLfUZCnSccg1WvhlSMnPqxvpXj0Zw/ns5UgUfNnwTrCK802Y8PwCiNabeBM
wRHoELQApFNzGxJE1vHWB53XqPZUBvA8s1a3kB3GUvYed3EQX+Lk9qc2wrjgEOSu
FgfNK086DRF66Le/dFNfag4yVbUcycuDb7gG3j2IbIIICGJrdDVS3gMJAGIDu8z6
GGJVZdEOOsbSU0qvRenMbTVROjzklVtOynl3SSxyfggTKUjk/Je4MPRvG3OxAdwc
p85WUTTw6mLoDHNmGhpaZVDnzJbDtjJ4bMe0rzvTAR3zVarup7DBMZ/4tPPyf4vu
9OYD8NhK5T7sdERAG4n9J/gmXEYYzH0+Y0Npaltq94vxM5l/OavBEQKxojZtTzWF
bIeWXjWn1cDLEjQbQgZ22Z/ZeyotusmdVIauQpyslPyhrjhrhNdgZT/zps+o3dAt
MwPIGPI+jurhxu1ALIZfj9Kc86Nen7N7wn8fmI+o/JMV45AL4z24Ho/1NQkAO7Ly
izLgGYqVtV9hx26UCUBLC0Q4+jlAkdUGug5rEp0AeSET6/KdQVZThepMrn7yz+Z+
DCAlpSe/CUcc7+fFFLp7Y0cc8pbZMYw1m49wWKgN/RR21tj0fNqSBkXBkTkC3DC6
HhRuRZMCBPUlF4rY7WJcmHjx/dWpY40FLiNocoalXW6GLhOIh7lP84mHAtek38Uf
TT0VddH5ps86Yis0Asso5KffUIJaGUlfKddtzZE4RRQR1VWuGbxTztafJab6xR9l
7530g024lf9Y9m6f7S/0RIAJHPtoRn/5LUQbmzi/Nz58WGt7MpJjM/SFB2Lmaz+x
HCdwtZ0hzTrJCw1Z2TNVKf+gMpT2dt82BIrp2pJrSmjtNmZspEyyEfmZ+Cjbo+3p
XqTKro3b1dxzLHFpVC4uixQf2HNtTbJ6mTzYkLfKKUayhlreSxlMfRIx4P1/bw06
cMua1hDuAVGqcMsubPvuVw3IzDmAcRDl/S34f8q7YGGhptoq3rdi4082ayYw3gHM
UQ/xOAnEyHQACKaCcS7yJi8FH8VxXG/7pKAEsGKp6f7SJKMbLv/PGqlS+IOb8VVV
ggG/DCtwS85fKrUbZKrCW+ypnFrEdyXhPw6Fc50g2N13Zec2LbW+Fi/gTWQLKcJ+
vYPp1DJmB6LwrmoIbf6uvdZTdVez7k/7verPVolVf59X5NIsFLT5UmB/ZS4hezWT
fnvMqW8Z+rba6p7BJbC8MthF9D6n1xOfdgEtrTgwvb2Q2kUCZZ2R1jMd4zxCQ0iK
mVIH7w677FkJZ5M0ksLev6MMQz8mpUuPmXkzONfYqPF81gYwa7w1AmkjeD4BmPcs
shh7lyaI9sbpGf4F+9s3PRVneoITHEm9rKZACMPSjFdYGgy3WzV2o9ufm60OUCYu
IRNz/sunD0HvPVZurOCFyHb2FXezT7RZG7YrHXtu/7NOHk0MfzI7CSZEwWn4tJmC
OEaFzcUZG2A8soIdQ3Pa2F6FwR1KDxuCQM63/SM3GKy9Cr0+wPi2LsXcMnUPCAyO
vwPPBE9emMkVm/fI6d5UfCOIw6WkOiAkY2rk/Lcqq5sLesc7uCEMnCGovZELgEmr
ilQvT9du2BFkg4gNZ1h0bT8I/XBC38zPjcawO4Wtrtfz3LyqdudcsluxRqYCj2wK
dpg78tjcfsxyCCjc3ih9gagYiHDzDqscn0XJGyDxuV47r6Vx5wColJZxfQMRrzK0
p8JedKTjDr+88WHBXKtkeRlhAqHajhjUVL/eFufhaRQYLGpUrO9XF6cj6Gsei8DW
2/sBq3MxO7WuLcJMy2fjGlzCmWwqnsjTI6RTYZA97pmzYqCmPBnfmq9LnEr6aVRe
HkduQLWhV7Z+82z6Y0SUyy1RR2kAmlza0xVDkdYNcMGHjb+ZV5NpNnYs7nrRJKNr
DC11MjCQ9VRDcdXIhgn9b0kIaHRs7/Iga6dIABzl227lWbbguMYz8p6fzVlqHYsL
o1FmHT2KVDfhpjwDUElfVksKMz12CEl4tecFGPb1U0X54kCltKzLPcVX+4TjKnwV
cw5EJ4b7BQE5rjuDtyvrFxm6HFPEpJMkxcM8H8dyA90jM92JDidxZSP8yig5tdid
ZBM3srmoa2wAo8kraeSb5ZX/DDGmDiAMcxH1zMa16OLpZkCEtzn7HCzmQdaYcOoz
EOPMrJ1q7t0udXjM7qB/WEwN5g5TxWqnfpI7yTMim5aCCVUmLpsV2Of7al+IDnHZ
jC0ye67AgHj6GLNusPzbNeOEQFTJqP3Y+zM7hcrPNi1MfaDPfQsyl3C6/lAaGl53
pK4Pdz2Ga+GDc8cCyWh3haet2LmJJ4R57sXQw+8ZVPlk7CKLBpqNH1kycF1SgJzu
/p31C8laCg2zFzdya7dXPhXyXLUMiQqjTyoi/Y/9qLaoSO2jCrep6kUJkv6HIqe/
jVGoGedUxLhXKtNC2Z/f6gs8Ay541AfyJFVH0eVyB9niTK+Nxdtmp6+TBtw3l5Xv
MOfd3PISupMKgs3FjiyBfVnuPlrxnvxcbfSi35XqBvrR+4J9QPUbX+D8c5sy3sQz
efOJz+KovktDAYMGDBSon/Pw0xZcgCUuOORrkKH3u5voU5QRoL+7weJ4/GgZUl+0
Hja1Enh50KE6uDylftBZGIBDi8Cg3iYDXO/DSN+sst4aelsJJnwQYkl4/BGoW2yj
nfqNRMlNA7nZPLoQCdLVBO4xm4uFZjaRG7ObsYYLXXUlnmvCG6DWNk8u0+w9Mj/9
vQR3OrhowdLapq4fYp+aR5Of+iGmzFfp0XPhcDUYziOuP46vt8jPe0yL7b+/1jD2
6MDEwMt3JtGus0WLdQT2DPgPTQ5z2vSLQzw99sP9XKHcMARMIWB95EdmuYRp0O+c
j2iYpdGucUo5lscrC+XQ+D7CYmY7i3YSKn5GNkfyWdhUjQ99CvGQ+jvUK4+n6toF
5ZOgP2K+xczocITnhIzcfojYiwLJiynBXZpQr0+X/Y1CqaMEwRflzAN0J6H+vq4E
rSSgEPdUQDd1/0xJkNun0gyJ7L9oNSObcinEpE5Uj3GcqZ+pdRUS1WBxfsFfgaFM
4V+3hvVCrdlqdljAinRvo3YkhP0Zr84gtCHMcJ9ZOmghFqCjenLCBNRd4K7yaTbX
Yt4ghU/7q2LSA/t9ELLRcbXuidhTHAKpMyUMosMPoQpVKlt5S2JZh5j7mqk8R5SE
YXNRbdIzHtzRBrSTd0zWUd7YQfQ0m5wOT0bx0VJdwxCl98IPklQK8UCvs+gCsvEk
dXnvYYZauscisy1dtv9MDwY6FrAnNRpGLQlQphcR4sCU8dq6/ZmR1YGreMjZXfA/
gPDqgvKZNYm/8Xz/efS/PPTQwv5wrfGLsKt4IjJZhxKFnTahfJN7vu/g1c4iqHQf
piM5nE/XWocx5/EF4x2TQoW9UGOX2aqn6TP7PlukLUCHvZRTbs2v7yo8Tr1DFHkC
IDuScQc234/C6wVs039Q6aij6MWDxseiHCgi2fB2rbUmWcV0wzZRQ1kiS+bW2UBs
M99B8tbxKIbgtB+HT/5Na5CMNRSv9ST2uu4+wbreGRrNb6lxqizOAXGk/iHjAK4x
TDci3PW5ZhN70G5LArRqWy70QhFLvCJq3mNfOHQ21/Oa0lBoRowtvGMaIpwrfiWj
dM9wdQ5S1OEN9RoX9BIoZo1niDM4wW3QCev7bpryl72dPaGLvGpHiD+JSNTZPLa+
TrmWx7hwpTqgyn8vDarY4Z9ly7se7fM5btMxYjzL5uutwpOYpC/phZNCDg6BrDVD
vUfhcRcokpUg9xk9vEG2v+/GVEnumG8W817R1nzRfki/8EPMTg0EvlTOG3BUKlLE
iz1i9JNDdCuoYFrCVgn8qJJ1I7sBX0FXm1+MrAx0IWIPcqKvvy2qUCeS3FZtnXkl
X/jhTKl+SxDD1curFBoE60vhWODLXeOXzTP4q/SGvY0ncT39AMICAkSAsC7kJen8
OW511TxJALB0QJQiamZ5CMOdQ5lDQJVe4LtMjt4ZW8ygpt7WiUlBaKQitEud/Geg
mRi+zZapn8Es2mnvKmSf7TS686yo5glr/BWBR5PVv6HTvoHixMjb1jjr+MEPet2Z
WduMWgeG6fvovn66cGd0KzzfD8WsnlYbxONSEmxq4HTRqhj4mrHat99cfz1/+eH1
FniAew4+B3rquzvyBRME/4Upyhrq7o5gWOlRrd0cRGuMEW0HfMhr5wE9RzXFx8M2
kGwNyD2SJcPFD90NaQ3HYMGjgkG6ka6s0XQzLF0up8DideCg4mOnMoHo5La0U7fA
JC0oc8SD6R8tElMu/kKz4JuXsyhaKjhCyOEC8fHK02usGMnmIw5harleAueCph+B
LUL/cKd+p+Ul8M2iZtjQpR5etTCwe9mj8Mjb9eWrzx03RketBfVB/LP7oebSGFpQ
BWNUE4e4CnuuA/kklpc0mz79IdlEAOn9HNnmGZ649CykTp1e2zAz6W8YBwkJzqWb
ZJ10mXrDIn61iLxL9UI+eFAz8AbOTfMllM+Tg79SKW25N/0DN9sMuhUVZOJ1UGbi
QbMMi/N9RGTIElnw1o/mjgIffzNjxBtzNBIGoQDZ5SWA6p0WDlG+9W3TOX/EtzwH
iamGeD+i2Y3C8sEFqouqnO5cFPRwem9JeSyRyqJV2sPqKVhS7el+eukKAFhyInDw
bXwwPNYkYzgv7VohEKzc6hJKU90etrQ4RUSM5Ya6REVraN3C2KPf1EDbKPHTN8HG
PmYaYqOrHZ5W1N3cegNzR62BZjLW9o++55onw56bmvjZUxz2cbRk+YOf712lnXBa
4wgd4xz21iuvVipp0SMX/o9OTM2Xx1a0ieKXX/Ket1FB/5uqoYolNxmSfSNniWxA
6fHhnuQhrmXvC2EMjUG/3eZzVBdY6+rAIioHLm2kD/jAn4FxYYI9vNEYnLw0EV0L
YxkVydumeqx+94HknpwX/0rLgLBhnxhktZpCrGo9qCqElWPJcP3kfOjOXhEm1cmR
dU5+xs30vHkGZSQEjXFqGKh68hAFFMsyBlsvTfaO9QNSGDp+kbHiP1dsu6nwbDPo
sWBEdiC3j3aD5vBSXaCU/cbZg8nM7UnjdY5k6mSTky43ZcTEB9PVyfHS69QXDb82
AxYdEbYbNZyYICkE/IvS7vc5ohUpmLAPMt21+fV+schJnLK9ydDE/ttxcrrlHX52
qbLcYPE7uNpmBVZ4u1OWkOp1o+Sp/587St4vRAugHNFI1Ltlfg0kYiXyau4MnhSW
WYWYDjgCrAw60QHqaxq1gxlEAgvJd4hLPzt8R9BMs2Pm6Te8hquTFTNK/1b2qNP6
gp2y5/lo/olONHb0prR5lvB9zRdkrcPouFm88bWl8jgbcy/V56wVy+eSL2+aUXTL
8+SZS43KrWwk13gyydk1+hP3tUArmWGywhieCGA3MP7Qvea/GIR5F1MomZO/z0rh
4xxd59fmFwQ/0ki34tsCmqIJQSwsgnp8gnIXrhi4NzHnkDwLO5LIH1kryVnrECvU
20XVJh2aeJJgZKP5PUogQf5ti8sP46wxv8rk80M9Byys/XWQ09j09/MEUvQyt4V/
RyNerOD28IrS272Qzt7w9h0Djw1awsJf46pgk+GlQkfioROYyKyoEoEr3CVVzhgU
T9I3XlUno40t39Cwt/uCntb5mtkne0rGvc5CGcbbfZ1p1O9D6m4zrLBn4UVxw+aR
kqtvdpb19U0A50gLA/GugUsV15rpV3JcfGRuZxHjub1gs9IE9Gy9MA05cfX1raVO
kzPj6V0y92ocIxvNnCq6dhp75d1XT5QObQ0XxGjtL+S5J3qacZGwWqAS97KccEtt
C/gDjSA+ZoZK5DNIqBVrdz0WNoQv4kIr0dbu1mcHoOh5jb83NVeaVJLG87OeTs61
5KwMSST7k30Jl1LTg/AqFQkJhH3C5PB0uh8ENm0TN67JIWrr+Gx0DNW0fXwGWfJo
qv8VDMsr5ERtAvBoRCCTbUL6Z63cgSEz9G5FrexigamtURTPbJnSk3mBp8zyMAUM
PEQP+a8acWPtyDyq6AqHBkdOXQYFrbUdQwnzZGKRrkhCOIFZqyJspzJldw777NTv
DSVUTmDTJ3n+1ICZ8C4BqEeQ7st6QIjxJY2Uvk6ozHbiZ0HnG+tuOyjq8VdbiWrf
l3cgkvT4F/A49ozOm3+DGtxiZlh4+7rcOIPqa3ytDp5bojyAUU8LCUxXs4N0FvHj
YO1CK2MPHiWcpOTvJO5NDwvFgry/J41zCQpTmuirhe6UP5mFCAhyywmvGleB7U99
z3KZwPeEAuey/SPOg0y4DOMZiXOXEGM7H4xZx8chZ9ZdaZ6I/+3bW4jea3cqBTrA
+QuJW9s5E0SQdEUK6Zp3ycxJhWG3jUBNKRdKwGCWNtkaJvU6dVetxXavhQl339QC
EhsPvxfhdXiZur1p1M4qEjSOMn2/qYHIRusjEna5KD1Ef7WMaDzMtejK7oR00SR4
PqiRqKGaa+4teopE4gEz5J+7/QQrqbw56FQESAtEShCrcDJYf0yzDm+zjAD8+g7L
K52GpWzJMZAN9CNuSqczIS2kr6xS7layHbyz9gRR/9K/zlft0a+XQytFj3QFxEP1
eW/hWGuSSbtb3ym76kDqnkizIdI0wYhup+1uVjZTe5cReZEPE63xJCzkrZJ6gSAa
FsQVt6TvyVFb0JK8qLvCNlR0OHi3eG6XeglHjvKsrO26Ly+AE3YmmskX7AdamcG1
ZFQU/uSxaG/LpmaCkyWB1auHu4hSTGEErFqb+a/eAhoeWU2/6wIKa2Lr6PicHUfX
LIckOGWh4AcsxWEzGURfExloClAZd/NABhnEXkiZL4P7Cp0RvC63QvnWefVFZScW
6MQTJSoaoeXum+9BMBYRzPr4YFHu2aY0/JrcCs8V3HL1faQ8pIwL91ULrXWdHDW5
YVPrO+OZQ7cChxKz4lJjY99zQJJ4WdNqHXqxi1R+OpY6AE0WrBK7W+n2n03/MD3i
Ic7W+0TU4EFOvBfL0Dh4yDpPZK6A6QfPQ5b9JH6JOvWTPv/LAWjSD31mQ0X8hPw9
6wqwCmTv6EGZ10LiSaaAUh1p82Pp06qeIyxA0RFLMb7XYA8LW9/0ATbRvcezQWTC
PvIQda2SlRV/8wPqt/KgUNcz8KUkPQhOhsRUr4egn9hkMGHgjjvST27sJPfvoJHU
F1jrPfQYMe2j3WJgOKDB6ByuzUHN7jU1FvEC07J88qKx6TIMgWxJ+11YIAxgYpXN
MV+e1gazTqsANJ1UBVMzWDtr0I1m2BN0QlhhNunU7TrOn4/0hf3qy2HJALuQSzuS
0UZPW1iKo7Hi5JbpXtR44BXd3oCnt51c/BY0azOt7FIGdr+eAQ3DpXkbZrKWCQIz
+dGtdMq5hG4kp6T8psqryrSuauyEeSEe6Xcv7S+ZhKfHOgFHyVYj3CR1qTkWoI1M
w/c0MXk9+8K+31AigRu+hAkQFyndMcZikFKaZsj/lNYd8s9bk4LQCjG29+Ke8h6j
40WLc1UaSK+ztu9SxK0OsnF6sYAYkJQXqw+1u1vP6UeQkuE3QjgXEpViYtaBsP3F
/MLmwek6UNRa8ySIw2B7mKDlUx8aNR3JhQuB7t8Qpkm9WppZINQYalZBTkzx5sBG
Ew/EaNk/3C9qWuKH071MRHbS2iAe53s+TsN/ayslW6Ih7agSCxzigOnwl2j4sgkt
NTsp+yapkjkZh/DdfVhHWtP9C6Oje+qdQbKXYem8oKgTyHPaD13PGKhnLENXXJnt
3dyT0Lv5kxLz/uh06klWyufy99h/kVPMrSmGpFt6Q+Rs1N4Of6YC1FAGBLcYtQvl
gbu47YqIYbLXS5AoKX1t8Q46dMkl+Gsl8FanG5IvWUcFcQmx3XdK48zpES+OHrab
dgA/DfJemKuygOISff1bwCAozeSvv1oojF2l/gFNGB/P3hGT03TWek9rK4Bu8XKT
BUeV/ZyJHd3lbVpfnTa6FqvRaCgzRr9xB3i23c80JfXlae++3VbocjWFMssZ3Co5
Eyr2VLa5Q2IKpLkwtf2ovlZCmGsHDKHQ5y+0w9W7W8eV2KlWTSdyWxeRLpJvPLFq
VAwBW2sxj9jB/EP8+2KoWQDOTJmsHCL3bQ0gXdlT9yQYkXlsdhyYI17TNVdN7H/E
X/+YvqvobeqtP0uuRaNIPANxPRz7a8XSRcAdHW02h3d35bAVKI77YER8cT1J14Z4
ZzYI0iJQOq8gxnrzXluGYfzwLed+ZdPMN1WXl+TtE06Rbzl+vdTCpjW694jFKvxC
u0T35VpuGg9H+wCwCxioYp6sCv5aZq/FNczo3C+kWDFqy/ychGzyCUcDgwyY47Oh
7YHX4jbM1gbWZXsFqTN7veGOUfm8fK+zv+6c2qOcl9CJdSKjWUrmUb8FQhgPnXkU
IerHuHh0BflflTVpjalrGKPzzh8cj6KfIuQHtjjfHJN0tqD56PIjdVyOT+kOmzgT
XjAXKow4/pF8ebD/1raR01PBRCMa1V9dnPBQlK8sKcAMj5iS/3k/MTWQNke8RAd3
ZxdesQL+G0e8wgso8l6Q+1joxZ50zgZaFP0OmYnFvMWLcM3HMnflkH7Fd5/kDrOh
AIVGxnfvrmMwzgO52oq6RzEHcMWda3FA0qBXh/HK6yrH2bP1G/PldDVSOKymcNuV
6BcSklCqJSg7f91fZGBNlAvaTx0kKk2cmuljZzB0VzikILrGdOYhsMURnX388VYM
dBsMyE32ypcy5hKj+QIpODc031LMfEciTlqB59WETSm+p5qYKQtiUAB74hE1Gy0v
Jkl+n1cOr5tOHkvWN0IJPN1IVnYS2RaemB5ulpql63drgEhv2v9nqPbf81RCE9GA
VQq6+UajPpOPSLjlMae2ZCMT2h/uqC0nbXM4FkTcMHMg2dwsB/tqsmgYjarHI/Bz
8L2XU2iF0sFrMuKAeIpuqFWNnfNmLrYQ2/+AH5IJqDk+UzNoHug3sZPnoy7apgVb
3bD6+T5rVvNPMQrXJAnEgCPGkppQRBx96WGYkxaGZYSZMas6WeOp3VSQUQVS6PNh
Le8dWZj32JeO9OitykLSwmTEiH0y9jsNgg6XwqPSGEk8RNt/7AmxCYcCU6nNjvnF
Gbitl9TQ2c4sekjwE2XZvBRJ/SPMzQDcjgjvkInhKmKCtG2AesHdjSSJOE/bzh0B
D/M/AAyUMeYFPUPkzRgQrOMdGIs1DqCCJVykewkx9nfsxzgQDMrlv2t6BjFLkAEK
BiGLvrMbczb4YvDL2suXwIbemiVwaJ4q9w3DAaCLdN04hpAX6Nt5mj/WlkdnSDrq
wB1L4JtQDhZRXVtgCaBbY2mf02zP62WfZCS+r+ONy8hVXjaLY0m7T3SrfDGXexN+
/OJSsVspt48LeFleFfDcCyzBmPj5Pbs7IUdBOGDx5+6rpoKEG8sgqOkeaDS/q8DQ
ZzuX6NEA8RXl5821fhSZz2LJiAFz/DOlMkIrsIwGJb6B7WC4wOPorCOrla9ma3VR
NWlpIeJOHJV5mCC4jaAnk29iCK8DL7X9P6+7HqZdX4o5yIYAh2wL/JJwckDEFY36
XlUs5has6F5eeDu9yoRkCR/6e2TjoXRS0D13tC0DeCPVaPuwRUyG7NUbDhUDlTFH
RLCN5E/UgCunqYeccJZt6rc81a4xDxV4yMwP0cAIzJa15ybtr4fHfZhufUIf9IKa
jzLPa5srtfdaCiReATwwnV7676WHfMlzxxxsoT8FwZ/kEtmpzmqC5xmeExTHhzn/
75Lwr/EpxzRSJAVAfrUtZypCeD/b2j1t02oErn6HHJqKa4kt1OGtYOwSl7nK4NXi
68aXu1Yb1YLydDpPo13IMNCJX2cdN4S3871Iic5HPY6EpXrHw6Wb4si7z/lf0ios
H9JfLzIPDoclJNuwRpWhJXXm2y0NL+S/D89oTCnbcrpAb+xMSEUAtMYh8K6kZ4Ra
1Moc+rHM9OY2hkCVF8H6C+M42YDkKt1mYIOms4/h6/4Cq+eujjgp+IYfca8xzF4i
QW2qXknzQc4tOj76eRKfG6aqfY4dw5N9M4h2j/Mve7ay/nhbKWz/PQmELCBy4p2h
5ufQt48lhNXUFgxTHV26jgHKl1ZbFPlRJpkbryuLXYVRH0hNw0/qmJH6jbaG4ScB
JC9hPnBUMjM7IuvgXcrDv/tlcXPe3jlceKcoWZE/+vj1G6u2VeGw0NTCWCHJHUFl
OFtpIhZXkt5AvNnPaX7b3RdV4O9La1jo40qvqVMZb67ALTpp/4F+wdtyarA0VzQ9
qOfBvuFIfPexb3u6rqbEWGfy6X0DcKQlb1c2LUKwv/PEshJGMzA11b2b8b4oniIl
e2foC3lZCGsHlb9xViO8Ly3diHf3iY0yJR5ir4ionHezGjDy0n7XjfN4OsUHEYoY
xyLHdc/V3Xceeq4Nfqy6KskruUrgP3JpOLBg3JXx6eFiOI8j9Z4x1UsXfWOwp0Cj
vLGuQi0h6IU++LqCJNvadTFv/RipgFETQNQLPe7ONLdzG0WWBm30nKWsXF3NPqAd
WC7ZKmWEFNgOPg7N1eAfFuVqGTqaS9fIJKu2jkp7CfLsyXRxq+BNwNQZZ/BngXeJ
fo2vl93kChG6Qact1jvfV3QpcSQIB6wYCWo0sLqYdDTy5/2P35kf3Sp42E5HKp1L
Zc2KBLKSyPH2Oh/mB58W4NylpDcDZaVahJJDrTvQuMznDhRn7g9Etj442ZyGWizj
SVRZgo4YU6SHj4EzPa9/GI/tM3trsRjN4ut6eyeQ6AYiwqAPIGBThMprQMr+kO5u
zOheqsCPl7p/jJZCivoGiFbiZ+l8uUMkad/iyix1Tsw3IB92SEpjzunQLB6yfM6v
AlP8Bvtp6B3wkMqTJYyA/Dhb9x85L7mrI5JNvlHRloDcT5g5gIA0kC8JZtuImh/E
PPEESkYSr0C6RQltk00IsGWgCjzFIoycM3xNSrEQI2E/WnzSgtbf+ziRTCCm9HK+
uCfJVlxBHm8LKn7FKddzRnslUjXDUJJ8CQ4HfR6cWU3iL6AazuC6tr7hb/niWHHK
OLHA6UsZ5FphkIOpqbuhX7T5NW5LX4U8SmimmZTk8rs4RA/qK8T0DMfKfutT5KTN
M3J9GZrINfEvOb/TQ5Di4RQ9w/xb1WnD80g5oYE/3CPiNJKgJ69tlbYV29QA6VC+
y/16Zi3BhSDTiB2ytH3Fuxi4W4euGley6wkhIBNWxm0KzuNxj3j8Gx02UrKan2xC
Ntn9zz4XfTnRIudoWeYTW4IZpmGfiziegkBR/TEOiSNKNac12czT+HCWOuQJ3VI7
8lJodZIXd59YWIo/XGZ6hj5/QqT7qp54vo8NEH7RDQAcXzAZk3lD0jWoL1hwpanf
XJcVq9zG5wYDxKVBkEtgNr7tHHKMmWuyJPFnXhH9mjbBAA9JJ6vzfuH7fgRp/Vmb
FcEBzH1DPMBK4T41NO5d6QYdEmN3wpLw2mPqCSeiTmVOYM+vNeFOKyeh6w0LQG7e
jDnKK3I8YnAb9u/T4PKkj7H5tkvgkb6ONen2gmsxRY0qNwIh+RoNnHnCGdRXsBjL
jKBoTHKGX9zMHP8vZT0RepAJ7ZRa7Du0s0vTeW0o3rI2zO9UZl4HWQwkNKmEHR+1
zao1R8N6s6OcEodVJFXnKOBT7+ERvF/Y3htPf7EFPOqV9lElBntWZh1l1SJeHV2c
aP5YHYDE6CD8TkyrCkyM0wIEWbUfQBVMVZyVD8jC8b/tD4lgXI+nKdTRv1o5z5gJ
BHFpO8RMUXuY+I97h1677EMBHh+yozqfwCiiKRERcQyViHxjBYjImSVUq1ZwAMB3
QNOik5eJE7TgbXi2Xup+cZWr0n3hshfOqoZIPu282YIuYrmo1PgkxmU2xwCFvVf7
5k1FfON54dPcbhtDB+I3Uapsaxwl7rtKkABAJf3z3mDaFnGY+Cqc7vj8SSy8U4SQ
oZM4rW667ojCPFeWnFwap0b1HDMsAsDI6Jc5xKJqCX1TI8sCiSq4RF7iY3TRFyaW
LzOGw///WHtgPNohUZeOL66pA+VEyAXX2z8iwZK7f5Th3MxZ0rkEQcbLsnSVAO/F
Ju8hGMa5NZxznWhbjRDI+F+1e+MDSn/gcA/Kn3Xu8iP8IHru9PlzE/DuL+XuXv3z
AJfjpYgrLd6Yg76a6lz2gpUoo0k5vx0FreCLlsrCYc7kzdeY/WccWX6V5bbJCZm8
5N4d3yuLP56wVAcTMxPjJzs8Nx0cVgtA48yvTPHbbPVU22kbj4Kq6A3KhPOpT0HW
qhwJ5MyqpyEHdkVHE1sMHvTKb3SIiCsWsEkSclYThVhUZIa5uqkGERcQR/6xWqRO
jJT+W2qQnRSQHHryvTQbGUfxMJUHhlt1dLZgHwzppLR8bJosMMTPkdY+u2cLvxYl
NQrV09SNVcm5NR9Pdry4NRu31nqJtHHzIbjrc+Hlb09xnwtYt7YuKcE4Q/uC1KMW
NCO6hGN+dwfwryYmxolMAX+9elmkeOl3ZU7er8/OcRJB1bEALGyZdW0dDCaQLyPK
aKo30r4+c8KmyCvCR51tCT590GawsWgw80vJ5QpjbmILG+Vog+KSHmTsjCqZ7nis
4EB7G25SUw9Dpc6oIRZoovzQaXJyDE2uLNFkv3b0xzdM6yw+1tQdjuejpbtfFOYc
ROJHPNE45zoATRiy28ffjvdgz+ypcHPQ/VqgXcv/4lXDaonaeWbzhkcpvv68zL8d
A4f9yCBjct/2fJs0GRaMDYAat+GtgpHaZP+TcAtAQy6tfXSbnugwfeles99XHMr8
ZYWBIfYi3fwWL7QwjNQBABv20afJG1NeDYNydpNtJWXzWRsdF3qRBmNsKITC2uCC
GB2pzybwqEzCsIF3IrB5i4I+FFCMHJhXuOU1Hq7dUIB3de9z4eFIYvkGiMfMbBC0
uvp5iTcegk0bJLZ4LBLf/L85H6KdDb3Z6/2QeABO/pbOWZc1i+JMW7BnKpQsCIPZ
3xyua5P22TmlhbHRuDvvcBOWRJRqvul6dnV4a4CuVpCNpm2y9M0pwMpt2bj2N0oR
WQb59oGe/H70z/kaFSkJrjzfxVspYHU3ft50C97GjMRRf9GdDGA7OcrZAENCMYiy
oPjHkTcQkTf9eCkL3oM6tD5zK3LhPSnHO3uNfK+f/N4kID8lBLUTJpKjWlT/ELKl
m4f7Krnifi6SIdZLteulyfsuD7VtloNjW+vUTW2/amWj+ilAoVyDZSObAvrpKYXs
vk82LRjKsgsH8im2nHoAiLPxUjWTWftkhsXmR8Sh6qavNOIQtlDgiDBGc80OCmHv
99FPCPHiseDMSmTjbhYsg+mg5uMlbdo+oakUK/buXCVIwH5I9QhOZrxRxQKB5TKw
Gw/vtmFl+0eRLMk8JcFA79G67QgBXhDDoi7+pRVAxKry74RurabSCDrEeaKWLwIt
omgvA2RaXjVNfFu+MaXZV/gTDB1p4E0NWj6hjUZwFNCxOjofTYltfETYFXEmT0RU
XUWLIogdarl9b/OAfn3a7k9FvLF9/em9dRKU8vlTDmozyfMl5zlwfiHo6rmjQ3K3
pMUAKXIqGOJMXcKzWtpj7UqQZ6B14Gu9A9aG3SPAAp5mUMj/O9JRjlhyeRdEugf4
Rb2QgF4wh/q6RTOIAjlv1wx9WFlnZr0z26z0erlWV6/jPw2WU8VvHCSmv/6fSETW
plHbGj7SPTwiLGrU67cVDKnNYAfT8AVhvtBcCkPO6gdcKTcn3oAuRj9Z1f+hIWcC
aS25h0joU0Yp0MY6fQ4UDNZDfYZThgMYAY0g2h16psFWR8Sq9sYm2I3XuLTPexxY
QTnHTz2oEpHanhfLoPHSRDKxKZsxN5rkzEczizufG7GzmIuq6utljP4vTb5yU/4P
jK0M5MBsPf9nVZOcaoKXSjEsDn/Q6+1Ic3fzfgCYkSRRrfFTrz6mCQLCAaE7HnS8
lnC3GMiKHxTK70xmDW/9GnBqipHnCYSg45MRtrb2y8faPx4OXGjdbmI3qe2E3I4p
qbkqTLPkzOELccS6ovBN7putXHe2pEnT/q5CnJdJUu7LDUCcwL03lULBwQCk7KAL
Z3vxRL+qCeCJyE+WLJpO8BnjfvbBZSLEv12YURm43NfxACyO+n+UKA+wox0KPxkB
GL8Krqe32DNTnOYvNb/6w0pjedDxEAYvcRdeShKanI31INpy8fc4YyQ7nmoi7q3M
dv+dYSeyB210G7a1LRBZiwBxeei7fpuVVQ3tcGT/9gkRIXWzTmACI0Dtd61+VJE1
xf1h3VzDgADDUsuwYgCqT3bOthj8Uk9RvZFBwibSGFNoRpMBF3FbRQd2Ailz+XH7
rPCvplnxGMqgHgjNnMkExnDW5r9l6nWmNNilIQ6m5t+wtlw3KVQ+rZNoylL0ujyg
NhirjiCPJEsYGkAkd6JOdQRfiY9zV0+tReiXJ4wA+8zZ5RYUpgzorb8JmRLnS+KZ
8dQB/uLd7ehI6/j4lwp6sERFLyh6gPQ5M1HQexnno0kzMlBk9sdd0Q6hPPGjwezd
bvvBLkQRN/VHosQgk3vI0KMqprn9ESC2VHPlvzaIpwIYHk0yKvj7MOiprsXHJs4C
D7eWl/ufOZ2J7D1DuCEdHM9qsywC4L6MpYEvX/EtITmqteRoN0hZDSwJlE5P8q3Y
ziUdMqh+HXW7MUx/aJFx7Xnu5gajRMRv2GAmxReUT4GNJO3l5GSSj22RI+GYxAgq
+fsPvpEhpU1CZ3nMPMnjCSc01g3HDIk8UNbiiHR4A3FN24vzICjiYkguQjLfhy+9
CVUGS8At1I3UkH1e+T4wfyVA7Zs3QkSGpiAxbcj/C1QxdEKdSuYxKj4XX8r29EgG
a0yyMEeMT+v9s6/q7NE3N2KrGpzIUEN059LIi6kbQ/LTA8NOZp5+aphC3h4RnX3j
mX4fViarrHHAOw1aYW0KByEXYjV52tAM13O4BBnM3gjIyCwxLZ2s1QUmUqNL/UaX
C7f4vnkt6j2ko53h5RM3AhjymYFyIEuFsvxpCgHJl2/EMYyB2I3INMRG0eyoC+Xi
x4b00jjzfFaihzo/yLuV8lFRB39GNsrIboGixeVyTBrGeQdmJqiYlF+GxXucxrqo
SF5GxrbBASfD7VAkBWwuVd7bAEecpCzhnJT2fHWLapOKX/UQuAkYQvmzuqm3Hkci
rbY7MjwLM9w3z3ni+cy1O5QzQu0BHXuw7DPTT9cRDQYchkHuwHulKlGCAjYLul0C
iKsgSC7ukmSNrV95AiXegN51sHzc3Skf1F2wEP6JnnuOKNWXh+no5pGJPafVVm21
oRsMXJAE02jK+BKy7b67euVI7zsS34WZzxVpJga8p1S21kGsT5WIDyuxZ+eXHhHq
DFqZvl5HrK65DxBiAuQAYwROVK+QEcugEFu/0R3Rssf2mA7n5XoiWS/RfUM57BoO
+LqUskUWLgXOT8ySnkoir/ft4Sei8pxVmQzYw9Q9pDvKBXsg+hJZ+dj6qoTFOx0E
j3EveQQjNB4wwU8jSchYg87NcyhcspD/mjG2hmpxbyR/TQUEHCse8uttc0gS21tn
hiYatCmlKzGE4kUYHkn9NRTvzAz73wCqDFZRvAm2FBBYWiiduHKE3NNgE4y3hflc
SMCraYTe8YdCuy9DwWeNUD/SemZUBVg0/Lz4aK8OTSPXv9OAOHpry8A5RakVavxg
rcrIaLUuKfoGIpTRFWahOVhC5cx2ndFnkz04yjF9cGba144BMaj8w+QPIsJeRHYi
WM5DYITMgD/dZU2IngF5MbGnpjL4XFSVCcuYgJ2C9JF8gWOaWbBXtwFQrL61xK5D
5cZs0DQRqtF0vIcQatH2M/eUqFKBZNK0XKEeNLZPi9GXAOj30wgs6NXZYDRDZwvT
ycRkwE5x3BJ2zgcTvAVt245935daPXDLrWh3xMmeDxFGHUE5nLlQMq9i6OzpgheL
EivG+7sajbv0kN2nl2MtTjI0q06uxvVL5IxVyCapgJYlFAIiow8e6lfl/8KPXmeR
CoVkodGM9po0SXPACc8eVPfCs90mbazNHEPT4VlTsV1kTFpQflH4pd48XBOVAF1Z
qVSSptyWxDr5lD5876EJ18+8wCdy56pd+UtucX4aVOtoFf/6gcbLRjvFPBDRV0nv
oNGu5gX3KH6SiHd65oI9uZVCwU4QHlNKfiRqQelZOTymlUV63q4adiGCGdBn/FB+
kszdR9PxpPg3X3A45T+POtCoXpC21BBizz1XdCugM4kQXNHGfYT00tt/lCMwD5Qo
TlhkKuVHOfgfCeJyx0ox9E4ha+m7TxVhggwPIYh7Hj9IYaQzGE15jxF5EgcTVo2E
1j1E6u3P+xtU+l+Q8W8PVrJI2jzL3rD8JG0/czHD/c+4LQaQVYIrfTb8S3W4naV5
5yePFMEwWLbu5k789QHttHv56tvFOb5FhmvptdaJkI+F9zhkMRnST8KNq9M+1uzC
YjHzzBX7c5197GrNnjTa/8HApzInhYlIwu6d0TNRvphAeGO8HBGnSujvdZs/G6Uy
ZbwNwP5Txvpclzf1XDnhk/AvlMnPuHMNnvxhysxAJw6PQsW6KYlClanLIGvPACAt
81yLtA/fHGZKjpE9K1dfuZuASuJxRAEJlmb3NmqDQ7kyTzhxYy8h83dW11E7GdUn
nY0JIwnGbgke8f8T7eNgBbgio4vUepP5SJ3+ub2B+Je5+XmRM369pkxVOxJor7ge
lH+szl3f2KdoZ1uICqTXccKGBHJuHEudm83JhaA3/ywND4vCA4jxOwqGWhjtvJD3
m0qEiq7lv9AnqloRJ2To5u+UWAZbFkuE8v+BdECgHP/iCxWYwLI9mdXgbr1FkhtG
ma3f/7YCWcEEiIzRJj2E0HWRgtgc7l+uTtptHHsrlLKHV7+R3IKaC18mzvSyLCiS
1oyO+L5eS1QFCUsi6nmTbS5u7olw5KIPlD5fLkDKB52SFE/ALPskopFDt0SOr7Fl
d9e4A9BYbn+EDjf+KTkHZJwx//aUgDclwoGo5kbmYN8xHJ8o3xnnuVqQecAvnkYw
JHKXBpfGOJUM9iWXG1X+O/bYhE6Ph2NggPtGk6zpOydRMhcQ5EqycOorDwuygCJf
CobYxCm+Rx4Z+uAc4ENTz3lbf4+CbGwvvR7UIV2am0NzQ4m3IEu4YQkzK43mLL1b
fV2gO5kx1+35+pT3s4ylTbr/H/KqmSI6o9MBMkuHg2Iim8wK8RifxPj8ZJEMazYO
6ay6rlraJ82aSL3wTdq5coiXHQiGql/KbjKTFdGJH2o4sd9i31rESi93Taui4f5s
3fOtpc1CH96kEJDIaQGpYj8kGEMmmYvSZr5m2Ohirx73ejqqC0nx6v8mo9YbfTxQ
UOKhbPUzqq9FQi0KPUfkXdHRXuDQvZg9QFE8MMDmH6ZX5eBCweaDlr09vGNGBHz4
ELyXUeAMX/T0h7vftMjzL5n2NeC/RWd9cQ6LCDt7YIX3D7LuB3nWNQc1Idl0IQ5e
6CPw2+rF719Cto9XiVRVyxX8Ilr2fjtWdA1sFlLvLNM6R9p+d1mYd0Wj3K2RciN9
4XNQWF1bLy7Nd/ASli9uqun8R4YPu39NDSoDMv2vhGWH6EuGNUPfoN+uByrvbykh
W4cjrynFCBug5tyTd6KbgQDRPJwLYPzjBGwSG6YLciF7YjsMoiy3DVisdcdrshyq
6TRwXK6id+uaUDe5NPG+MY/VU4Tnyl9vug2r8Of+XUWu6LtX4dQ79zpiQ4szMkLv
8mRQALgKj31okcXgVNYGB4ERdITMe3myUOOrk3asoUFEc0DhtMZ2uzE5UOfq1FwX
AKU3oLvfNvPvqedlAngVGDlbgFKKyF+k/ywl/9rTAEeh99/NOklaEQCKmNmIhOCM
hHWIewWdB2cNExopcEKv/SxWos1b9ODMz6uI1hWLOpwT4PXo4+IPxZ7hYsuab8Vc
6k8aoW4ODWK8Z4+Pl61VjOUwvrNXuY5Ay1tJ2NaN+oOwlaSZW95FxxCbukkMUtwN
qASKfvxR96lFYUIfc2JgYtek8UCedvuXwPK1BbSZLnEy+W0wXwdHwg8/kQIrzQPZ
88VpVIO4nvD5WaOah+0s3K99nUuDigbKCJHhg1uk7ZDgfr+RI4Pd63X0qDSdNvBS
0jbRmhPak2FKse+l4T5LGLiwBjQZtPGev/6+Ffo/6gjL99P+IJ0QpVnxThENorpw
RA8fP8d91YkqtdNXVZWmuWIdvjryyBZuWQtgdoBhPYZHNXmcDK4MXupQYes6KvV7
YkRBkgeJXuhrQqzj/yEbGQOD4nQM+vZhckCbrIprmUR9njA59HZdKw1buQKfZLne
eHt+lb1AEkyymxomdRMZaJSmvegZFdG+8qGZpNg3BJF6t3DQvTEv8sIWupNh+WI0
h1EM80yEuE3B+lUK6P1fXko5eDZ2Ah+UptqGCCO+ds4QDlWMPldNgCO8JkPb1b+t
9/0vRNIhLZqFKpo2FcBVdn43dEuokWVWJZOOcPPsxgjFDl50bYgxzDiFdMfyAgDo
fcWtis1lS6FexKDf/UWUSZE2NkuYDedZetrbu7oJwXorDCRD2hj52iC9ejKWTHhG
zhtA2QfpzzEqVaNuuHtobecN97J8xvEX8jixoK9IyktB/+DodgY7PNmGPNWf2ge6
Ei3HXixP1T+WDRPGQrfQpSK6oeHa4hedff7venwKVnk1Vd2yLri/056lObZL88V1
WpCTkPrDGxoncCgOAM4jOtJqJnsV9FQo0hFfAbby4llJFhcE3tv0uDI9Mg5Z3JP5
+Y/brocVZdPXOX9PdticnZoQM7lic1s5W2e/JKUUU5NmieKELC3NKLMmUizKtp10
3x1F41JKi4DGeomMMwH+95JlLKnPU2tiKHuvhhLz8IIz3X1gIziwHEhxPsZ7jFjJ
i0vdGa9inggoMcCu8UJXklV8SIeSLfqxHRUapZNa4NNX7AtHb7pZJbI58t6/wqcA
nqeAiJLB2zR2EuyGlhR2STIyjxtubL9HDGdhz+LubhzR+dpwe8uuuJoYpKw6WSL7
Gns8o7rM6bjRnjKrwSFhFUFZiQ00+AQnEVZ00wrbY0VDcZGCCgbgDdxVUbVdCw5G
JCMbDEDQEIODW7/WGFHKTYTzFkucfTersKjua1L8QpYANEHdlai59Hb98NF6Qzs1
cyQAeBRDtRjdLk4bW4GhLjSeQqKXW0FJWJSAGHA2JbI9HgdrcZZ/AV83DkfyO772
WIPScua7wAxCDekVk7fkDVHsXOt+grCz2e5qAYe/08zPSp9lwNNb6HrNpGkHaUBx
b50Oii7chtxTXk4YdfYa2Y6DvLgBmNCYLNgYZlC9sNIbR1gKGrgG7SnbKkt+kLjI
SfuT1zMGXxweRYzyiFWyh7r53cQJCCqZSwqggMH8ln2zQ7OnHWbQ/2RYYptZcA3o
P4uZqdGCjUbnPzGGF3O1UZ/cEDn/xTR12kNCZM8amSIaEEr9oa9dblCULJoVXnQl
sJIWKo1zbC5keE5O+yVafbio2w5mXdnt8o/A5Eg3D0N4S8LkaXkSTDyXafjB7Cqv
48ulz+4A8PzR5IQw7Q+b7JjFRVUERxONgNrdAVfx007Tejn9FdThcNLLwApEH5RR
rrL1srZ1d1rJ2Q0Oo2etMxxBPjeZIZHn6aCU9LqoRCNv6OTNZCFOnZs09BCY5BsS
vbEbe1Hrh0SpuW3j1UeUql2pXPbO+1zlRwTh8ZFALOU3jSXdOwl1rcOmxNoWJGDA
etvvaXQ8vHVb4Z0IIrPcnlW2UA6sBuOjms3cNV1Xy1fn68cI4DG461nPPUbieM5p
r5Y4daUjLJleWVD6BjvbQDi5lEB7/zVQh+1LVXVRT6muU2KUaTs/QZIlrZ4RqIIN
9YSIqNe6khJuC4jo8b/sj4Akr34SjQFRSBIQhMFD423iMO/pDbQ3wvNDdMD/bQKh
XMLocbqwFeNxVFVs/p9XtML8CPX/Odla0o4nasf9lfygOSsvYf+gTor5oLPqIxgZ
U38mC0gmSr//oPb3PbGGt5p0e4YC2X/sSuv14l5SXz7z5XTSuut3/2L1irkD0Wj/
sOn+yBRlyJSam4nsOKdlHZ2lIqzjnSG5rnKbyx32c0NNker7aKrM23rkxWSRP0/w
gG1o2eNm8321lTrx0HfztrqWWHSmHLyM8HnP5RyiuRBoZY/75udRkDj01GAfp3mn
EQ8wAFkWRWD2YkVLjhFVYIIHOvTTjBV9VU7e27ahw//M4vh44QYt91E4atacW1p3
icfxdkYkxge1FoS9MmViVUhN9VLfbrXcc0mTzGsfPjGOCOEr7oy0pSfnDnRnz9Cd
3ppgKY9Kgx58ZTzpBykekGI/SI5l0r5OTQ9BEGfsSYAx3Tx/iK6jygF3Z/ocm8gR
GNtzRJLNRf+gvUnw+vbnkdWwb4Wn6pDZau79PTnGd74UZE1q8ymj/7UWeZgZq4z+
VN9wnU513R3p9x5YfIwUMTtJESdOsy5Q1tjzMnvirEAArlHo97Lv99+HESijQFwC
Po3yrs+gwm7m9wtVl3a3Jzpj6WvdzzkqeEBJi/25HqUEFz39OpQRGeBhzXaYdZIt
s8nlMzyoZqFbD+RZf9hKTAQUAhTUJG+SMEwIOhX/PMKxWTngLh9pfmC7oRuwQOb0
jvE19tSKSxDUo+Mq+ToqgXo03grrv7nSQAJdj0iZfIXpLicJUIBF4WXemMzYde8b
R8APo7x2pYXEPzQq8HB3SfCbIHfdmgZOpHNiSRG+F1rZpwm6BAtQ3KXV/oeaU+Qv
G/uoWjZ2pZIKvKm/o9Bguzp0uFPJV2VE/kC/Lg9Gv2bYYufZpGjGmGa49E0FdJk9
S/YKM3Dp0sFQjyjQVAFMfHTjXFvz51vATLYU4RXzsOlkoCeUxsEKkxB6XKuR/Jyr
E4NL4uqfs/pvOLNKwv6B5ZeMq6FAnde/G1R7kHZIM8fDZAXdWRg+6y0zhVBQY7cl
y6HI1nfUJk7nOZeCRxZc50nwcRQFYOyU6vUn3437cyd/rC1WH8o//ThS2rqtkz+A
2739iSGWQDMG5jvadV0/aKNBKxHJqPIFvISfVHrSE42L9xLwtcWxB6Iera/E4MUk
8XbaH4CFwcC0cuGwuF13CqiZwXCjssuMKYV3bAiVjhU8HF3hUlXeeE0J+LXxLSsy
pdEdbDu3ZA4zKPPmHwy9On/XJoSkad5SWhpboi6Hzh5XjTFu2BH2lHamWBZXaRWn
UBAcBNxKrRBZWKBB/hNEJMghijvN838aWE9GXwg9ZJC7eX+Svbcdyo+/inXL9TUr
dI1qGcCsEWjUt1diwd9ehw+Gxi2r81D/g1iQ4PbjFMl5IgCkM5FfMAcLVoMOcdnB
D8Dw4fcVwwMaRlLGVTOABqHSEF2JMwxEYS1yOz/tQho/eiVCW1hbuDbvtbt6XW0C
hqwkbcOkLIfC9dlXRq2jGRYBEcRBNJwmBKizKRQd7En4WhXung4F0vWRg0Rs2OU8
/IsQ/KPKnLkjxqrGqcoI9EIKqPY7ivulScEOyARcHGzMpvt3nBurgkLZyW4A2Egd
Z6t0w/NLyPp8V3X/HxTERXAbbyp4Tw56KS2cXUuEjaqV1xjTwyNQ1EC4wTk/UUle
Szbz+Tcgxq2HckAPl+AqbLSao8rAk+NSqOtiVLZcDw+lpNPCmi0PJb5Ek1BVUGVI
QTwpk+k+bDaL8ao8arSpaRFdYmmipcpxKs6wBiTv8cOVGsg920Ia8OjW5wCczPW5
Erzb020bB92YxrAl4qzH86OcZSXw0baJpmYb1j4rzsW8qFRP62PVydWvAtNq6Bkx
Gplq74ZXvb58Wwa+GvxPOC5pVjh38BoaQ/WCN+sa+r7l5CNdSL8anJqCzkz0Z7Cs
GYgSXe+qhoaCvBkB43A6ZAWXovJjsfG/DM3eEAvBfVYuIwXyVDlOpoAL09vytDK9
rMtiyYkxlWC0xVTVpDEdTrIkyngflawxpfx7N6TRX6isF+qP4Ow3IInVy67Cc2Wh
0IdedsfUVqzkyO+MdB0oGUpBNkA/IV7N4/QaIJ+YKqWZJx6VhlSu0wTuW8fFYP9y
AMUeIxQkwQ+n+LZPJNu0b4EqAcqlxzcL++652ftM3t03c93p4PD4lvrFoy8VPI0Y
8dNDYjyWRfiLCBDsrsrfdF5i6wD6nNiTmLxyohu074pojoLuYmY0p+ziUlW+hKsK
5NoyM2jKyBFVCadCuoe+IGiR/dznZVDtW3/NPNoAl4I9GrYyE0euxcq/zXJ4ZtLx
aAGNMiPtJNJiPEAvAno4x4/jfptUC/k0hAuHBtIhnra7WkV2vVeeRCFPtzV6dyLH
cAdsC0vF7WL9O5GAfTr/OfUUWpUym6vY1hpoRhY3yFZjKLaRfq53Zs0+9xyyMns5
ybQ0huIhveQm3+APP8bZfAc5ekCFT8oBtz/adsaKLIhsT4zTPRieAnW8XxcZe0O5
s0yJQLzBsBtKb3OkHwE6bXsV8A43bFJlGIhUom9PWyE0JyolvW3pBeEwJZcGRvpZ
tgi0o2Ldi7rCIAEmLOYBFz/nqbs4MOzPp7un6vSFGz4eSvEZe+nv/ZYnsledMcql
4y1pChYXNUpUvHw6uaCFxluN0Oa0wO6R3vcbU4w4M5TGVDlI+hcwWckjC/SfrazF
3hDpZ1rSUCKh1gudikEuuYvuVZgQUkbMDAxzgLMTniTaB9xraybLV3zWjn5Dcarf
usvVyxSOqBYMkuCGaoqoIvxTazEaUYgZR5fpQuXKT5UwtPmYb8UoP3fqSGYlRe0J
3IaqPkiK21IOxuhyqzBW7tvBEXQk17vqPNy8ZChlmEiuhyw5+vL1kLQ8wvrnIK5p
qNnbChlEZ6ZlgpijFbMLpxT1tYcvFTEsCtH/WBIJ2BfnYqs9umi8loz4WbFTWJkb
50fkU6bqN+qRZNfQoQhYcxp7hazwmJSl5C4r0UBewSC4K49cu41+1pf0sURs7IF/
DvFTd/v8cJVbW9IWCaRXLg77cgi3CNFMY9KbolxM+TZdiz8vs5+zXYlVYIOkUL49
YRdzyKyQpPK70C/OocinfGF1QHsxxSjyBmHrsio96i85kLibPSufrwRst2EBQNPf
CQ//j6Sl70xKlid1lun8cbrOYSn7eD6EYwK1yJiZdJwCQD+NgFd8V2+tBbvrTyVt
antIZOrARBoI0guqtnf2tGkMBj+uHzbzutiKGgjNs766X5vX9Y5f44Ec3ZptWnRE
idUtc8uiKW1uxF8epIWEhPZzFVTMiP6QKSxqI3WKbXYhj9uVCE8nZJzAy2JKkYcC
ijO6vVO9JQg6hTqyw3I4Ha56WkjQ6ELB+2LpoKVAlBjnP2mgFwGNkabo0RC4cfGf
P1Spp62ePXwqV+1qbJ7+gQuS9g2pvQSQv8QtNvEdQfwoh+Mjc8R8hq5URdeLz4+G
1R20p9Q2t0tR3kb/6qKeT125M/vQdyBwd4pradQmXalgyAGkSULklrvdFM6PfOYW
VAr6aM3GYe+qiX8kr2Yyvg9mEZaZz71GuRfJlCAu7upzktpC6pD/jBOPb4wx7kkE
+6RuykRfHodiSDik4wrQl80dZ2RvcUofeEvO0tsevq13lVKdWfDy6sfagm/R218G
EszCKSGrcOSeuldgB4BbLM9uovxNXv1MxvUVjh8HBYz9NosfF8vf/CNZt6NXDpCc
pi5m1kCxLL6DsICL2t7DnqSLEkSVlIuG/g8M82T+ndhAh/biEpc/RWTCfc40f/l+
1cAoyrrE85KUoaEOCd52b5El/L6lDi9y4TtriAyXb483rz+LT769pMCK+2AekgZt
SxU/LvmPpjemgAgaM9SsZaZzurGvOQpjcTeZUFTskECtqjWp4r0HpG/YBNox/S9z
EMbWyXnlrsVl5DmRZF+akvCC9bxm3au5eX1oSsaIG6g84bAe/v62GdzO+bd2kxO7
roWixmf60eHrhNydlsDlULfuXZzEVjFnR1HLynyQFDikHJ6z0n2n+LpWKpkmTNHF
fHzOJXs9JDwh7K3Qw3czCTkF3cllD6YIPfXtOUJkFplYtTzVOFw9q5DdqOYc+1sZ
xUmICgZCQufHyDXJ/zSZDhKrLi6MMmllweXWfCV+Yi94bdD69wWQhQEOYEf+NOB2
6FD51Td4U2jbYWz1kJZR1Gl5yY+T3T9xS68aM9NfDcyTFwtW3Q5n/HvyXE3E/wHU
9OVmJqLRA8QSZXmTT9CtlgMNSLTp7hV/OoMnmnitMUWWVbJkPApcE1IjQtUScD2j
cTW0e3LN3BXNZOyDeNaaPXifhjmqRy1Z6Vb8OUSTEjbgHsiEo8fNfzGMSQFQapsE
vGe8uvJnKHUgKQOU0OIh3+6hDA1YNKaPT1TsYyQP0UpRFhFDqSG3cf532ZnRmQrK
qZ0G8Zoc3BBr9xSQ9fqY/5ZqlBgCzi+HQx9M23vWAEpbN82f0BC/Xx4OzGVq1Y4M
TmsJG3obcgoBjODJU2qCLhDXR5U3XXq5GsaJgXr2bnyginNNRau+BMyCWOaNoDZJ
WZDpIvM42mXipknxEhMLsEEmyqja/oX5ShvMad3Re239Cs04LPm7FAgjl1XxOSy2
2M9FXjizzfR5B7oLkCKn41KA5w68JV7FIrPOT43DHkacwUz+d5KTn6KR7CR3/EoX
tKnvN68lL4XpnIaMV5C11rBDwX0WeMYgLDtAdEPpUe60YgXRGohIhujugvVMD9dy
OZst49j1XJZZl5zpThQYD0lZe5KDkqW2AwKkahWs6weVMUV3WBZ3GYNJs5e4qcs/
Ln0W+3vTETVEzJghFU1yTexe9e0plZh31Niuhtc9gDNd+vDYgfrJaEYVODyME9Nc
heCNXE1W7+PDMze/w57NVV860ZsuSJskc+Cy6+qlDV0LyYWYAmG24MTE+XxxH0No
+/kZI214hVgpDcH+FtdWhv9925PsyWKrmkNZhHOz3CA+0tlj602b3n76lAKaRd2l
k1OrMdtsbTJy/ptjTmUU5z9THkTFRclu/FZNRfQD369gBhe41UEPxiQ1MYuRmNLX
oNLHrXpSk2l30pwpfgwOHw/e8SVyCaBYFvisYZJsgkzJEV7EuQSpJ6F3BXHcTQHU
cy1l0bE4MQ1ZEeE2hTOsI+dSh0rfPfb0OBavuZvnv5k0bcU4/mkOJ+/jz2fU+XQK
L5oC89VPhVqUmFuPkpzscZ+AbNii4qwp6rNAvyeCj4bdXff107YJPYqgYsWRPlv1
WHr6ML+bkbksRb1/zQ+PBmPA09Vr3R9Q9oth6RZlWpIaPM118gqa3dB8wa+DZguY
kG37eaGHDwVCrjjAo5O+dcKB8lK9KHe1pO1BklETVdJTnddr1MEcxfnA+StJ/FzU
u3zFiDkIrhboBWXwwRqqL5ZxiWpvC026Att+boayYRMCty6E81+aGNYtOdjz42M1
1/zmzUXKSSE/d6SCunvO1gr0VcuyhP71ne2yrqIyaTbKx16GRBkc1JISLvZ29oVr
7jHIJgeNcWsA09+y4t70AXRc5u/CaINDIwd3W068FaDCEAdLeYyuINIGPvalbz5s
GSO+lfYYxOGYZy7BsPG3woE6D9q2JrHjp/iaw0I0sBqXNd/rifKllQovwpYTU/j7
IBv3tOZll55Hy6OEEaUI3hIrn0dNPy/3N2zIx3ZMv6kmqiuNifTT2TLd/PoPlaeV
vZFxpU5b8pxNZt7B5Ljo1ZnWCUyiJxARPrjuPZJMYtatbshJaJdm/0IPzMWT5AZ8
dGvJ0nPitPMrVaWPnOQ69MgOzu28q2G0WW2f0CT6vyTHH1lwcZlsKAkijIwbgBLn
UeCURw/8OU4Wvlm2JIo9ro7b6CtgabnoKm1vf9B+2g6TonMeyA98KGA5ycwu3wo4
8lGkCYHV+LCv1GuXTJ6dl5f0svZwq38Uy8Sa1BDUKuFCzIhxh1ovT5x3kvYfOU03
MhFgD3cqkFlBfAZdkzWfT0WZe0rY2/BtINPFKg63GsO1wSgDOw5JhCv+wka1fPtK
SpDC2Maw9hsItrRvQznM76Rvi48Sy/1nJbPvwmsJomeKm2hCS1Hgrx6pXWsioQiY
jcAn0ac5X+qVB7Tt/zh+hxY3NfCHB1lMCh2Ycc4mKy33dq644kdq7KQ6wXETkwDI
WRieDAaQm9GQwcsKtKcfV9U9E8+lD6FajeNy9rYzPvsGTv8ueVMsHAiOkscL5Tda
GXAgOHni5duplDKUNoK022zr8sEvyuBvC5rWmd918pNDMJWzU7xf8G0l8Y2fh3FS
OZANEcToyxTNwNSrfm6SpO2+xEgvM5QhXf9EaQ3Nmur0Wde5H+f2xHG9PwWg4YF0
qMi33b9ghHZqYsbIZWaTuTFLntzUWcTRsW9OxOOliRHb44CvlzgtbHE331ZFXeV2
eqtlI5ZaoTK2uP53H7m8bSzoy34uQlA7JbkOgAtidDmIIWUUjgNl0SCM0yPIsBrQ
yxYgIWbNxlXJozT7dHeWTplAjP1cWZCYur0oJ3odfaQWKdkuzJofOyvZ3Wf+zV0r
k3M+9D6mY1tIZDIWBaf3Zn5XPpmpqbC0S1UAehEpJPLMjNEFzrToqQPST4BJBipW
6NLIUDffothfUA8YqWw3vikfVq2hLBpbP4R/ihwxP1iHCKmxftK+u2swbgN66leE
U7Mn7kD+PE2tC7CGHlDT2W31oOKtPsTjygn8r0JY3vANTLYederMK55m5/Ppo5Y0
RxjHUlmzC1nsF8tJGDQoMG6denFWYOwegFMMGiGNC+NCgU3jtQF98XCGcQJ90upN
idQPbGaXHHV8iIDK6ASMZNDXVZhZPKFgUDJT4ndQm3L9jYo/C+0uce6/d4nYhRPR
lnsveVwsQKE3QkjQT06tuzySp6MQNEYXOqF6kjlZLKtbSLCLhf9f0F8/b02qTy0P
14cAq/K2ZqDhW42y8IdYqNHBL0qGi3fmWVUCM9xn8nlxCupfa64AiXRKK7iwqoft
`protect END_PROTECTED
