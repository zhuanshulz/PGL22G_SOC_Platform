`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wClIOBRj6c6Y++i6ZcLMqiBq/4mT1H90FCyxxzQLt5+LGFuXl+e9aJqJOSV74iRQ
fLaocqY3C0B+MjLLUuI6sgwAL4Pf5NTiBmv2iNVEIUi57gZrnqxbOkf+Oh9ay4Np
NOVP7Eya6M4hF1pv+sUcnPpYwkl++dtEqOwwSWmOPTYRRRjSeiKb5yVeqNk/sURC
aNuz3TiVK5h4U778j9O2jtonY7w7ciKyH5g0ckEWbUiA2JDZbnSOERA4B2PnELne
5keVQ6li/NZwI8wbAAgs0vGV/zWUJ7sPnuJU1KLomMP24OVBcsckW41EoH6j29/w
1t9LMgsyYnQNClfasgi4e5Ew8xFXajzLKYtAX19q/c0lQPfOn/lSAUIw3lvWdI3b
dASp3crRbvwdstUTx0fgoXZV6tE6Hr+KYC0ocvaXrSQ=
`protect END_PROTECTED
