`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9lIqaAY4jB+dWOZVrhttGASbtXYTA1qoB5Yjy8cPnMS/cLMSz22q0rUxtRTz7U82
QTMKRL4bQUXducfQm3fHHzkm8VD5XR5PUj+XV/7FWQnwqvY6fZW9AYVQO4nLDNVJ
IWCN2FhSRjXkPNcpqNWRsWRRB+Gtpf/yP51Pcu/TsuzZ571Au5DgDLhr6V7EtmLI
ybXhV0+Q46kVnOVou/YicS8iQlU25ZAIjN7Kn93siTzUAS3Du6WBFR6QGAP08YDh
Hoka7vyUupUl/6+XPIX5KoluxwoWJ++B6iwUPtx591gzlATAGVTLiUFs0pj9fvDp
kcIhQzzCifJ/mTvjFQmcDB7VRphRUghxH4n+ORNcg+hIURozcTX4tA+UrYLdFthc
rcT/zm9lYoJyfMPzJoHJfna5SzLdZ6MJ4dCT/cDZZe43UQ3/Ey2TZG7jFnnmDx1h
0MKzXzk1e/wuglysW+5VSFJz48YvA2p1oRotullBFI1GgKOXkcQ2Itor7+2HXFie
13tGC5XyiOZFbdUAAzZWDVsj/1GDs6nqrTq6GmU8n9ZpwAXKylh6LdP0Z6vCFaF0
sdwPTtTQGCcTbEph0CYx8qECo1Hc/9YL15KH+4J66dBG7qtjXuq3+eJ8IOFjNLdF
vWCkSU4palVmOjKtYEenMnE6GSyGIGkxTVkSZrPMaNTOVkD/1frze2wJMCF+K8lw
HY75VsXN2OJbiiXelRnUH3KheGZjHnckzG7NI6TthwI33Tbd633UwzDgainom5Q4
fUT6SMH5IqlLleqIVW2JDCEFT68Vs7KlvfNI5IXtQZuYfgGi4jHY1+PZ0zCxavnx
6/fsIroLN3YCm4j2LerDqzOHTNyPQ6orc48/xbTPYDPiJ1R5uhYv/lJ589YqtjiG
TAzIpJc6APTCKRvoj5N9uQHTZxSMq4M0ik98zARaRqRcPMWodJeB2hDC7Bp+JcQN
I0BeyvaCIgxtOr9SvuoX9Fq7lmQHTNnUv8p2vQdlGHIAepgqt5CDWt/cHIswK6vD
l5TUh4V97gp1Wsac7VPQdpLJ1yBjJKpuG46zd9p49TQv5NDKLhOzBQH3ekzblp2s
vmNpxDfgS2yTKSpSQhYONhDsvL4x3xlV7e/7eC0f/kMHJLvSM6bLFDrtIpHOZJYJ
fLTTRtwTV/LSw4DjGPSJcAsafKq4YT6wtGy3B9o9cutAc5vFlAEXTUyUzK2fgxZq
ymhFYE0xKNFvT8Mfek5XpiQbYIuzZEnbhIVq/SxzKbkOASukS3AaLFrL4q7pQj+E
XWE1NPrq0NV/zYZDNdRZ+H/O9ao/jkLIpsT7fpdPoWM2v73aWrV/AUiFEMtwD3Mw
msDgtncTyPaDirqqYCU95mOCKaee56X8nLS1szLNwrTm+CIR6tgpN7LYE6qMlg+3
NeoSeEsg////kx6D7CX2359HcssK6PBC+IoWJb1pLNvOm5Ghj2M4PkfkR+B5Ad+8
VcgQEwx4Surt/Xz8IyHsMhx42IbDVSjOKD4xCWdZFGWoYnkjEslQ0NOcpLkUluU5
p08dPYBYP+e3L/U2TgKLaWCk3E1NvrfJBB/3TXtxlaETRqGhWleoGd9rZYfLBorf
c5eP7YCzOvdKdCbYCMJrYc6qnU8EKvjHBOT8a+lVK+z+8480GkSnyqUeuvYxR3yS
mC07itjbqwtCP8/6LKZ+XXruVXXPY6RZN17apR14i0/D8yBXxbD5odhm5jnHAWfz
ZeQDcmUpEuF7MtWwEVaHNCHXFJMuzA8LBkyC//9jRU2BEdlVxmY6i2SedmBOzrOm
7BYrwx4ckMWN/67/MQ5jpPSibTJRJebIHbP+7RG/eJ9ABecV/9zSHwI8Frsz61d0
dOU8LTUtyglFzQyhla6U5zWRH0Pgiy6XvvTYmTQL4MjMsXRhuxrpu+1PBXVfqX1+
Pb0TIW48w6MF8VjHmXJK8trSUnLKesR1k1KQfpfk+cnWL4z2brrhzqtZ7nikw0ol
TLHKFcbW+o2FKFbMnlwwZynvqfmn1pZ2pOidPIak/I70hCqdlKC25biflMg7bZxf
GiSlM5elSsHR3SvAYF4yEbUNX2nU6i7WrjBKybB6oOx0Av9NqTkzVIjYBqv2cvZB
D8VlcSCCpS9aTpYPARy1zlOjOLtRoD8n/gyPRW1bI/+X8hrZUr0lwntfJmextnTb
+sKgw33tZMllMO7SHV3WcsbnXDLCu3bslBPUhlodZZ8wYPuhMZDuumXK7LGRsjH1
4Vdc6/Zf7mtSTGIewv2uHhRDN67XADLVtloo1zIh8aInHPrUsNvCH7Bo+VIWs3Sp
+/hfdWVhzsZLA1vE4xHPOd1FSECrpU6wA+aW05Ddzd6lanHDLd414FBQWCD0xYA1
yTtAXcqKBZfKjBi7HipF9A+pKevkVWPWijf/FZ7N9cMYGNRrGlEsydLDvdgj5k6H
5fHjD0c22ZqhsugXlqaNVNfhrIENd2DeuoG5Wkg+9EXQDLQYu5yE5e6/3h7JXckY
eSJAtxzeY2YafQNRS/uLCerdS95xnYR3BHA1MtEl1fpxIA12DxqhqUE7OI+DMs+A
ZXOzmpncSLAh7WJui8nYIy0KYpmfXpbb+kFbsBYpib/Dmsap1lb421Pxpr8OW4Ml
7YNWQlwnXZ3ff1xzzBNLdHiBuv4A/BHYuouWmBv355toUiSW1FmVLmbdoDo3IHhN
RoKFx94yqrbThki2fuMS+m67Cdycaq0sbwDzN7vlHX4SjvxUq535msGNTmZ6CsI9
jjwE4iS7hroTK09cHVUv+qhQuSinKjX90/Ilcmhnf+0l1YBVGuLVtWldlRrEYIkh
vOF0h69N47uTG4EwTQP6TH+jouxaH2yIdQR5RJ4Rw52hNx5c++dwEk+cDRhhdedp
4QdhqJoiBnqsF7Divl0mR6gify2W0uqqxVeVQOAnZT9l1jqhRxkaPKQIwxkqlRkO
n/31PCN/NZ6rgL5JGqUy/2xFUyoaEkLN7dtn/CVccC2vDuQIYg4g6XdFAHMjTaLb
HhpXou8AnVe4HZVWB3gY72hAAQeXTnO3mqHgEpS8qFkkbUR2qFTpGCJJbBf2aqaZ
OHRL6ccj7E67J0rLWyJgDyfqHNatXyxgnYuOPbuiIQnTvz7UMZK00MniXJ/0efIp
vafRRODZTeCeWyK29/SgsQLeiHsq8b/xXybOAmtKFc+BnykWQTfUuGS4yO4sH8/J
0zbSPB6QoJJ34kVOkmnp5XDpF41du/yH8CsyYcLdybeCuuaUxqtqJncqM0lKcMX6
C413opUiatjw2R0FJ8QwiJIO2cIBoSSPpTFLLo5ib5JB94NEEqUW2cGznykK+xlt
QiagKPURVf3cCLeDLdM98qvudIGUiOsgydZHsmvR+DPsGrbp8AyK7JI4QiQvDk5M
BrGQAAbwthJ6zm8/GTv/aFmFIXV5hzAa7xiJpgkyy4N9zuS4Y43SfPHAxMuMMAJZ
iJ4tXWsHoeTtyUVBwUmBJWrkmLfHexwvbhHLM7hIAgwF7KQcYjAdKYSCjRKky4dc
h99vl62sEcwq4qanvBqwTDa8ls49u2u/Ox+nZeHd/La0geitc4pxGEQ+jHguSBcD
SfflGfGT8dCZCPgOAKBxA7niELTVakUfQJW07vuPCnpmtkI+Y9MGZHbkIslQWPHT
aLYw/YWJb7CBRYqjbIi5tX10PiPXOBetRyLvPzvviNuEguSsBD3uxHyCEi6Msu8h
fuIGQZCdFAWDJlyLtk+NKEQ2F8QP/HWldEG6jhqGg72QNSc86EP7FlU3IIlXG12m
+8X/MMLmcAvbBdW/7ix8OVQREAB1sgeY10FOZNo9Tw8afiCaSg7jaiCHDzO31VyX
Q4q4DhWFg6NRzgJQAZZMjGerIynqGxmeycU5OFXAM3dufQTCtgXP4YqDSJxdRs2e
XARDIcNIWJvzjezioXpw85pXxDKZwrJtVfYNY+Bm3lf2pE2bvtq2PLCgdJSpgdxR
9ab88wDc5t6q/oZfYSfaEp7bZkE6T6z5KfclfEOQ+R+rv1uziIGPlYhb25v8g1tP
y/2zbJ2xAWWC9FcTFvKUCFtY3W9C0uKRQuinfL7igui3ghsRQ9w8nxaSIVTNREy4
Ik7j9NrdRUYca28MVmxtSLy0vlKXsJvjCJbOPla0xZbcGFAUHKDg9jr61EkvZQ3q
J2GiojYHovtz/iJ0AdjE3tENsdJlVKVLXvYxPkGGrPec3HPL2r6Jr8MQxP8mvKLC
RzLMA5CDggV4EHhrM7Oegq1Vue1L1F8Cjw7M/CXqOAKzKrfHzguIfhMpheJgAVL5
INL2X/oqkOW4Oc7vtbq0MbEyARteO8PT1YVnmsO9aqgIctoJBPX93VG4i57eFcHb
F1pL3RRkgMm54dLCL7T66phSOdab+BA7CkfunPnbERUuyUK9kN02CBRc2SH5BHru
IPthjZFT/kUrgGHvcdKsqe1i1V2peDnUJSxMNUqQusJEDhYR7CHQhEu4k7cl9u9L
nO3Q6YwCy+GGh3pJDTDKZKloibzLvkByAIzluE+ZorVdofJfRzayRmt+7Hj6uV6s
n8rNH+vk/l6E58Tnf9fqcA964kvrSxVQAnSSxVNJ7TkrOpcvrZoRN7rVtVFFT/7C
cBkCJndimv5kZ/hDECW3RC0kGLdhj17bR54wbRahhLN6Fq5gt3qDqQRsLOs6Lcyf
uGKuOjJB/YgFSWT9/8ym/V2QKn6DN6ZWY3sHMaaANNlSQwvWeJFLMx1Zds+xcsvx
FC77k1V3S/zHOSrqmXhdy10+uCLcSeRHr6PiAhKSCYasTDTeq13mM2ymfatxdpyw
X6vof/k/y+d5ghTkcIzu3QPXCZxFDpiPyDkIAK9vunjpjATemIDF2yPrylDp0o79
FXyoxjsAhgFy7qzpwtbKxX0bzwv20Y9w72dCBbMzRj8BWdCNV2R7OdwuEU8m4MZm
nOpFGi330vJbf7HpKHPJhunlfKa1yynPjC+tFAUdrFuslZ5WDoErzQVpopkc4JfO
Lavs7OSprbtwufdKsZ1YkB5AqJhBGyuiCVbwKP011Rly+C8hod7jnnF+9FV2Kn2O
yMy7iklm43KVff3XgXFgC1H4EfZ6KGqeOXZoAtca0FOSSAhb0s81EN1VSlhw4CD+
ZbtfhpJA9nXgEebzhmFh/4muBd23J50idxC1BlPAN724QYfmtjY5SM7QWwvjt5om
wqENUvikgjPPCVPJ9PAZfeZxCMmzhivaaDzwvmqmRRxPfJ5U6xU+GGtT+pzqyEaO
vDfO1Ouh6apKVoiaArMZtqVJJ76poClWEZ1dVydzza8qe78zx5TA0FM5WQ6EBAfl
YFdOvrfAXsTPO3Oisdd9zK6skXKaoi1sjrYR52AN80gmf/EskPNclDdx7Qz+Lbit
OvOV2I+twar2LqiaOFbjF2txy7fkeq57uErqD9tgxLr7iIxBoPlkU9mc58T0Z7hm
oAcxxH7iQ8ZRINsyQvT2fZET8HE/YK18dTZcXGq83Q8lAjAVLy42DTLrHovbJ875
x29Z+QSsV1nfurnNQi3Lsj3QnRLk/DlXmOUjCphjuxOpLtU+YwZnzFp+v6P6k+Vw
s6+74Niq6rKnQ3SzMZi0bgbizcyMtd9rAeUeMjsp6yH+5BBFEBUgeChYX9yVXfDZ
ZUs/vTonD0I3PA8F0FKdWw2843OHcf34j8RqVXYUIyXOc8gqys6mAQLkQzy55TSJ
dTO+O6DxRCiwx+RxMfsMmrwwelig7Bi3e5AJsXS6Y92YlFwIynRPyHc3mdfADLqs
wWt623tUX3NJsDKF1cQW+xMce1k7MQJV+rttdR3uMHaKlH/n6gEGbqviy7WQH8jo
HgrL7xPcIaWxad7wW/57Mw8WAgZKyYl/5ia9BbSMeEjDaM+mpSv3RFYWQ2296ZxX
1k2TiL6+0rsixBqdXSR9c99KRZzwueBq+nPXC/4Fd7T+vdhXfi0FD2J2wKBbtjR0
LzXgfJxWylZtYPpRmM31ybUvDVZ6BX1uvWJjLmX/xHbPp5YubXft2WSuR4H1B531
U1AqZABbCPnbxRgFrwUJs4vjVi9f265Ud8sCvuegu4i+iNrlBCjsEAK1mUyEp9us
hXcdZ9kglwld7Bh++lLxnPhEUzLmnpE9w95VgKmJhmRErRlHrxWsD2tQSgBRrC+3
TP+q8Y8z4Bd1S+evTkXIq8oJ/PcbGa4yTUEKEYBWE1XD+BK5ZCYzxy22EE0abqfz
GxEmtkuwZPYxv+BZL02Vo0LArzpLdmAicWXSK0J4ep5neCVK3iferqoDnqFJffoS
mXspe4f7Vpqr/f4T0qtdT9cWiASNgICap0qzTQrUfbNx6QDLLK2+E6rf3QU1uGPH
u+RLEG7KzmnOEc/+xQ5tC6E+nPNnjNZoct4p6MiT3Ce1h/XQVdboRydAn0+lETNr
9Ffo2xj1XnsgieoQmr9HbEDo7ViZnJN2YTEjq+/0w7hcD6ivIaaHja4G8UDTKOur
u/oHFDCcklH+Us5aHmwqUOc3k1eFtYaEJb+zh1Q/CtFrHtmEJmkXTu9ddXZO97hX
98kPJMlcz4M+mGHTLR5GltTBaCxdceP2pBoRC3gAJ3iPksKS455XQ6y5eS2/SK7J
guNudUrgpr+bnDhQJH2DMprpFsyXK5LXq1rkc2pBS5rn/tPKD+zuGITEIa6neajz
OoNmMNO6WCZEZceqN9z7eHCaYIYoSUyqZ1/SIcFtYukgaqgHivYzB/uKJgpUUqb+
U7MKXSG75Nov6EYvcVxsXGs1u4fvtTW6xVotszaXRt3XqfIQ7EVobuUem7Gv8e4Z
XIvJTXsqn11s+ghtABKctbSZDLKnR+tewtlZenfs2R3V6AlMUt0ECBCksOE0dMnc
tZbLbZDsCHHjZoSGsDK3ieV5qq2jcCTxPxoz3tHzJtDDMv4zvvqAXqretS5061/W
ctxJrUSUdj/0g/sm02xTcF1d3VuT/6qmPsZDDsCpScmxSYEWR0+QxbVHJp1rEZoG
0og/cJYorfWiuX/IzCWtb013YJx33DoMpEFIw501C4i9EirpaedengwDaiilfd24
ksyu1rLNxqn7bRCgX5+puuqCczMDOEkA4liHaKW+ubbsG2lhov7MLvSOMsZLct6T
7a5LoitzvwriywZD9+c9jHBUSUOibugscDShQHPQuGdzMnfTevUFPD4vfCZQCbfK
scoXVBlBMTT1Dt1X47wGEVCsrbkHuQuiLG9H9XvHqQ6qgO0+pyBPzCMQRngXYk3l
LVvJBbR5X/w3E1LR6Vuy2dSDcJL2EfI0V0c10qXL308CPc3JHXPbIW+kfUCD4xG5
C9FvCeqgASgriF0bYkVmlqiztGVC1XJaknbeWPNw7kBkdevVEioE1WZFL1zt6IYN
XicyfQf+Fs8YfpcHb6ekMVSqUIceJ8cFRRQU5mQj3rMOXfetI3/+Fmy+oz6a33Fj
rD3icVzkX8fxPcaDfoB2JP3MY+UH/hv5N+DA1ja3SCXJvcCUsds0baoiBtk7Ccxk
xa+DlwenpRB5U3p06nToLtpBVlS7fV+BQ3Tlusq9IM6Ieap2j8uyjGWM8cr7fXP0
0Y7ZttRfhlEeBfAAa06gwO2ByLA3sCxvSUIEFyFcYzFdfY6kAOMGeikn575Ae76n
Yb4BLXsR3kzGNdIsJovU1Ud2iek1kFj/03tigN9S8ZIzSZuVVjU80+VGkvXUGL8m
+NgarwlE9Ac4zw3Vx6T7wC393FQLWGKhtWe4tKEPyFmlaQOJF0b2qZSfSxnN/eEK
DXimaHOXflMHgozPV0t4hnldin3cUSHkmFxdjtx/Xe7EEaiUrVgZ44A1yEWEH6ko
qr0jlsm1uDprPoS6kwgkWV6h/k3vQo3ncLc5292QgQNvQHSxvtGHq6pt+fsxDwjQ
HWMDsZ/eDyZTnl/dT0TfXjg62bAuh6vIxYc/tBfuE/GbP8yFb002ngwWs520G/14
HPQcqvAvsPo4JPavN1MvP2D1Kt34Xr+ESkNgZpbK2A1X6OPG1Y2pFt6i6bQIvbMp
IMEr8LYjnlap58ZII5MSDcMrej/TYfGO3bVdG/s2Xt9z8PNNq9IXs0qpzIwOk2sF
MU8h7U17oop2Q8bE9UsddHFsF7lVCyGN25+Sk4ZXV3C+X7fhTPqpd0jj8K9dGHBC
Qc5eJDDU1e5adLzCcSB6CRCTVkaU3y7iq5Fa36QLpDb+Vyfnxgqv53kbxQOoQDj6
dKfVBXyHVuLYsDPnna1mbQ==
`protect END_PROTECTED
