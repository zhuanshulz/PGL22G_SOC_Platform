`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/4yZkULuq+ihuTsc7whaY3ZHPQBHtQxRdjVzSwjoHd2fgBzGvmjE9NE4y0ebZVJ1
Bc6joo215sneIUsa8alC8j/jIJ6Jl0W7q5wDtXtHL4zeKOMTLDCRi+x2BQYoXm3n
jD/8/kOin2xeSHLzgjniC5qYlV7vvYQfBtiv0W4aTTsAGI0/XMB4WFUv/uxJb70U
784O2XX+hp56eI+4TZip0Ikc9bEjUmdQE7RZoGRsJ3iQmMTji3X3hngl2i7eGkVe
yWUU/oKfl1OeeeCz6+NllvNkVFx4aczDU8+tqLREGO/Qze4Cvxb3zVurNQJu0Ybx
BC8YwSIKOaMZY+fS+BxZig==
`protect END_PROTECTED
