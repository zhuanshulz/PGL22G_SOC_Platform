`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IN+EC1wU9f3MLw2Xjyy5ikHgYbirBUmEzajVrEKAWAZA2LeQeNUP3mMFMgN4nJAl
7sFxLJf6tP4KJLApeWHJ3ykZizaZUx7a5VputGPrSIwCeftWl+SNZ+lQYMcRcshU
0raIwJ9lfdpj5lAzqz1XykHLVdnRSUXPGiDNNpBOl6ilZpEQzMD139rqUIErnXi8
g7riwoKWUneHNzf1oqzHHx8mxLcndCATr/aVFjZM25W4IJghfxepQbv+47XCt110
ogyK9IX73PG1tVVxj6WnVnsEOkvHtfRvvKwoK11f+dl0wK21bbJ32b3LSDk/oSGI
QMrx01UicqMkcXwExSZsW+b3cvZP5bdo474S+bzyJ2dddWf2O7OFb1cnJKl7QiuU
Abk616ByR5xh7ly4Aeo4RD9A5Xakz/He+vWY6Doma1mTk+QayiaFEMF4ylSLRA/9
xlNJcPqW41yJoBTy5dKShNeEGQzPBusGyqSb93taiS1uWRAyAVXpRtchemqxHv0O
nza7Lewq+rU4DK8Y8Ug2l0GmVEBaB9gWGqCNReIRiuquYcjKbAMVc7QgeHXDg99u
/iJIoTk94h3Zva5D7y5hLdxxFwYY9zSXFDVUTLMof2h2dScki+N3s/IPU3YD5dhu
7DTKM20gx+ZTdz7AMowP+nUtacDXV7mP09+xg6dg6iMUO6byMdXePNGxdukYvvFh
IKTyAu7fmKm0egAT4elznCc2+ll2fGy4KRmdjBroeqRphO2fCG5fH4blMJb4aUGU
4K4ojzuZ8v5wfrXy8zw2ZX/HPvNXV5l+4eQt3sS4WMEG8XSbxKX7h95pHEjy6wYT
BgQndtc/vE9LdvrTmNguuE2uGOicE1CXpkQNz0NvQbM9nbW6+6VqoBPB1YS5aq96
G4PdjSqXppfxsR7Oueby4tbSnmg6RYWgkuvPgntqb9Uu0oZxDlTTxAEwY0wPMrmQ
1iTTHFj7EQEUyYD6iZLHzOwXeMJkMAmmabrZcL7DY7FBPLS5WF8GFohlGRWa8SJU
hJAZK/AjmbKvmbUCA59exr5mZHwCBaRLLdW/d15/uTdwbgDEh5Ig4vEf+ei/A3yL
j4jrjZhoGTTH5dCiUR2kJM61q9gKhx1s7cn29DpjL97707BfEB0GSMe/fpAh+v7v
2NgZA8amalBQTdgTNDe9MfuxXL7E4IGsPj3bZxicZbtQg2JICX0QhzwOMvynGRc/
9M4177Ntj8ekZGYT4Kxwq3CCWMsAaEzKglujdfu/thRNXfGLWk6V1XPY1wJu0UcO
lV/4/MrfWA2qmyUDjytDfjlGs7f52Qkkn76r6+l/UngFkYzQjnxqBcJtnfS3BInb
BjM5IkmXwIglN5M7e5FrKGArLTduaR3dy/Nw54nDKERLlAJvk9Q+1Li8pvUtnLcT
FoETZohEDMlV3B6lOk5/K7Zxdl0orwJ0w56sx5K5btprZmxG8UWA4SVwu8PsRYP3
mmJHrtEqzyxjC4LfIp12yO/u+XcdrgXSah0kp40Ssek/Qrb7XjpTa/OnlwWgrq5Z
+ixJkdVi8zzSNDSkVKNTdEQbshJoWItpUZMWBVh8VA5sBImaJoxZEFVZDRbsn5z4
0juNGfx9Pbz3tO8JphOe7CZY9379FnIS6jkoxuTi+wiqTaROStbXnhMKB12w6Z9h
RU5Ll78ODa4R9XEwhhCRTGCfRUvA2I3F8n3uGBRDuENwbgD93n27w4yFknXzVqIi
RKboMuC9m6GkSmlWjGQWnscsAjIEd5yiTDjLHBUuKvVH00yJYxV4LrzT2tMJYD4H
iSuaRkCHm8KRVY+YQW8SNaIaoKeSW+wnzc26LMZkK+kvkg+cI1JxjZu04Dh7VZ6T
/OZzW5Y1lCNSo+suObRAKaoVLYFOzU7VxZCOACLe0iMomB22EcmBdrBMbnfJfFE8
TSFLFRFMRsbeqPE/r4cH5tVtTUTOY/dFwZetXRdTaiypHt81KfnJ1Xr9/DQMnB2U
c1AKndKpii5e28tVjHojSRz2rxmZlu7FypGqP878HZmzb0ksXsxn79RKo4FbRoih
aFU2i7ckdevlkAy7JDDNzAQzGloKyUT6vyo2w3W46qWFrjakjqIqMTjOKX+1HEi9
2eMr1UTFP/arMSR38zOPGFkXU5NaUjGOuEBoD5IH9v2qP2fdh+yZK6FILJrHAGuu
0oLUUWZNAqwYwxAYTWy5RLKkiYZilvQ+gj+ELFP399uUi7BINtzGCeJIl8JU7Ohh
ouAS4tut3QbF9H2r74cLU84WfaeihgSemAsW9mNTnCK56PVjAuxEVeXG5DiHphpd
6/4oGtEBaCoNKGFRLb+LQO4W1BOD4h1hsLUDsZ6A3ISjtMQ126Rr79Sgef8G9Po7
eB2zk4I2Yxu4T2nDvSC+raTiyZFu9CAE87DMYnY743+4iBeF483RnGWdo39aZFVA
ZU4XRduQHRpvhi8TPSph9scaBV26ilaUq4Ty9PU7WFwXaM73kVz9fLpWfqa85BrJ
pwem5rfb0+0Tk7cTNI/qF/HEsTEmgNJHcrtMWKKEXw7HTh/7PKbt3BcrVOLbqHRD
tsC034g00LPVK/8MBfi3frZTl5/Wa8coN61swnSsR3nv7WL2Bb1SrI/z3598EOtY
egVNvw1QBKEmyVpD8kZ6Twrl5/lklkmD4ay61gyOAnqrnDHWnKOinMFxcnLgXAyC
7YXRDRk53Y5J3NoAgn9AoDxihJPg7lPSEXH+5/qJgTVMQqOCO4JTsbJQ6TnPmFba
tIifh66xWd0iLN1utA1H9mJ4BD85G107atieBH3O1CZEAry3bPRqG3lmR93mQdbF
47VVORuxUOZLzvVSFspLka20OLVolUmsIaRm/pt2IIf/pvVNrfl2wCtP6ShACKhU
es94RyLA5yml8guyKRwj3T5Y02msvaFSG9t964nDDLR/jOv3j/vaNCNFI4lxF5qz
uzUIVzuzJKiH9WSroB2yBRJSR0vOHneOk07rYvVkOpS8vXlQo+77cHlDYivltIOs
pu4yLRhQjwTikuroNu3NQsigXKBLf9sIwLTpD4A+LGu55k5OuBNIkIX31M3rtzzv
cQIPVp2HxDQ4qPHTbLgGeuJyPypBbuCSTQxnhdciDr8irE0yirxNi9L6J7KOKUj9
yBlpX5tP4gsRdPEbOX3ce0IWI9TdFP/xDhI3Icl0wfVTj/FI64IUKvJYldWXL8td
N+W+UGhbrTCtv/i9fJ3vVCxQzmt7wPiNS9B/f1htR3ivwClinjPVLjoiDhEM34tB
H7jumZtZ/TxpoFiVNbB9g4jeEEs2VRbdKS1kZ+X40rlQz5w+hcMY/lKgYHcaAmnO
aljz8h7lw+a3N3xg7bkc5ELg0dsZ6MeGj+wAZn6WQo2zdae9CwTl9OYgzA4CoZd/
O+5gCao3oC4dFwm6tscN1XyWdgGH69WE2iPB06es2LH4P1lEnXj16gtCL9F+AJ6G
AJmQBUUdGMBRFYkMI9slfhpW4cNq9yLnY7zLZ4RFAIBiCD+thF5U+ot2urcEOuQv
kbwJf1QyZobtk5war6mugOioIAhV9OWyVMO4ekix8zJstrBOHspDAnDd9vg0VLGG
nFXXsgBeHPfeSzHsB0+QnaFCnj8e5MGW5TdcDu37cqnaDvfIUdHd67PGvvla0GTY
lrGbPlTy6dgKl0g7dkLNfTwWLL9epKQz79snbD6MzBlIftPPktP8oV2xS5vcDHjM
a3HjEhm9WS8FvJJqyriEcrd6Wu6UpOAsJTOxf7KzoGqho8TPDj70qnJZYQ1gXbAU
4XEyckYQBPiufPT/yFeGqPYscTJ/tu5aUqO1nNniYH7tx51Rgy3MPRLYaB6mgcjh
jKwkQ9Em6grVtC1VupyNvnO4/rqiz4px46KOUZa0YnObrCbnrjYUmFjilIJIArFp
077+GJXJqki0lxWNMGMlMvyLsbbTk/km+b/P6x2nQdlvULQns14p/+Lqi9refpo5
E2snFKroQIaY3GBoi/srsdR8JiMyhZzxZKX+YDMOiRo1dqsGBlyN/owQ/b4PFOsX
XumHT8l0KgAB1IAPYr2gVrDJ3325uUTw/3OYESfL8wpQLGkvW9FZRXVH0VZFOHw+
lEwIxTAtgZ1fRiRKf7kNdCTd6BUpz7lNRBrCcjg343d0RPKPzP+KZf8NqoW6AHM2
tRWgeSEmr7mTlakTep5n2q3Gy3WjEhzMSdMcgtnucEt7NhjLWust6AvN1YKopdYs
YJiivcOVzIFpIUNjsn4gA4UPiBiItFPNjDoCvLtfHYa+LkAjdFThVH3wGuMrZkId
d3PyePgeJwOCIFQiLl+Mc7mXWiaYsAd5+kOMJSk78SgiPr667uwg5fUsIED70X7W
c6kpuLPJl6cxbf6n9FkvqMZMrcRP8DYahCDUEy8qDzKtu0FccOofMVTNH98emb/T
4BhiwHgLC32sUp8ipe9/U5rtga1iTKKoOUZM5KFV8NUpjcK0Ki4raZRGBW6zDZzy
8N9ExZJBHEXlCJzPMp/BKTmbolGc+8zQ3qdZDj3Yt88JfVTbb9WUsuo5N5AT7ZLA
kHXYJKmEiESfmGK36fdDps32200jDTLZVKLy6GVdWw1zoTa2ljyZ3+mRl2rNCZzU
UUOjylAOMbA0qdzjC6oR+TVr0cebBUVOyQsVdC298rPmIodgfyWhKo0PQOT90Jat
nAG3LdT3+DF7ke0z2gQM9fbOgPXaYDY7V1AsTOt0P1Q01ZPZhNRrtM14lfFbolGw
7s7drhVYomiKAkzgKKbmf//eW+QgjfDhiVXdgsC3yhph2QxKszkbp2XMfhkeCIWO
7Ec0P50XIJR2A2Vf/15bro8rP0dgPRfCxkDhIaz5NEKM9MyxIs+n1byy2ADpKaza
H+aCyAiV/OOO6BbWm6/4WIb40kWs3OpFY6ZT4GpcQGDRnRURl1XmdvnvP3brDS9U
1c25WwFKTsorZAhp2CGsdTZ1DGP6Xistym+yCkmDas1Jpt66rOVlWD3Krbgi04HZ
kZBCpUFjQH+FUgYum2S0CWD4ChgFtPq6QwNdh446zQYbZPyEAr3M9cDDy0jnW4yJ
AFf5si+Vd0swwDylfEoMreaghSJG8AU9bkqwgycXXAgnMs0SquHy56JbWP+25xj6
6seCl98sV5J2kiBGGLonEtCio7GDbAUrceej6Fi4RATRcqBa7knB23HuiTr/v8xA
5DRA/sIv7Osh8klPQ5X8vJlR3MLViVDRXgGchjttbQBksBBQzVbv6GTorGATN1EE
hivZ2lpjKlw3+cI6SuWb6dGcXiUj09KGVrPgQPksOUolP69HiwBLLdKLcGn6jb9t
T0AWVgLzLojZ7cHA/N03M4bXPpg+oDwJMbh1MIv8QbCkRMMVXZ9Pge7fPlVmglLd
SEYY6zjL4oHRV0X4LBE8EzoGUNjVEb1qx0A6+vxzx2heHQZdI9i6237aDnQYQfGA
bFeAZhGvPaOtVwbGuyVg9BKTwUx+m/Dm/ose4DXBz8oXOcxHo/rmIuq4iodJ5y7c
vwRlTuRIlfI9cseeD6Kbjg==
`protect END_PROTECTED
