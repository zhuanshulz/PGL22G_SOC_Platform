`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hy5NyUB3YTexi+2xQOWNbtNi126DvmDxSJn14Zn0lsCrV6TBpKdUjA0A/+M+Qyz1
vdVMUxY7gWW+48HSvApRlU8KSjbSEOaM/EivbQk6PktL4iNDzbDs14U26H/Q8FEI
YsgZCYUmZKodvCtSuL4UVjjbeQT5B6soS7EkrIpfRozLj4Gv1SYNYY1HwLx8ybkx
UVjIhN19VeODt24zwqPQ73TiU53RpHhG88au1rWABsjtc1DaMgGCIR7lUd+nStDq
ws1PoGhAGbw7zevMFIVCz0Zbh/qJYIHGLP7laEkPRrPrdpY3G8Rk0EyDFernkrV0
0fhO9ihF6AT0mJ/YQ/4ARuRrQD/CeT9nalMTn0yZ6//4D4/RFX/NM1mRdqMnvvk5
A6uhyuay0ARaFc+fKguaLttETVwvjuHpKcx30aeQA6rucHoNC67QYouIqj6qMzbd
`protect END_PROTECTED
