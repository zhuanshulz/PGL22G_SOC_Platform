`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R4zEEXL5OIGSDLZ9iYuJRtkp8GdFV2vQAlka+iDR8ml70JzsOEYQ3tRuXV7G9Afy
9yFiVQIT4d5qAjBJkjBVj3CTSkFH9YIPBEdj111/tRo6/xoSCSCwAX+9jJn2w+w7
dVCZ9ktwR4brLSok+Qdg7tWRG6IU56U0iIAtGFelflPzBi8oF+n5b/YaHTSWUtJ6
ccDPzul9Sn7E0O6nOsn1m+YH/DkmikUyWEUkS64xuDvNe0YPnNPWByYOE8P5DdY5
hpiq4roaSnOLsR4V93KYpwsWl/OH+quCnp7rHtNnM55FQgujrHA2ZnzRqoYIAhl1
IxPcLD0/ALxIFryu/Shk2b9ojTHwH23z6BNr/Ef9zg095AaYMeAe3lwAeDeutJ/v
95Y9FuzdCi02le3Gvw3D/VkrA/AO49o5jKa1pbli3iN7F+zuTy9oZloOr1X795Et
`protect END_PROTECTED
