`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wZYgWHfsUG7nDKhmKpSpKxxFXuRgPS5ZKZw8JW88JzkeUH2Z09breU5TxJ5t8Evb
ybyly/uzD2WLgvY583jfpqwS21fE3yBCwEwh+uqE+gguYwPQP1L53IP1rfcnsaS3
mL8ydkBwSyG+5q1appvlEPbNQ8rCy6DpVtLbb8d2+dvUUTNUiKEBF0BapjWBQRo+
IWtcz24j+pMmWOAQaX4wJmfar9svtwAg1FmdxzMstagGJKWUSrV1XIxg+GacKSr9
YTKHS+UoNM9Yj9uOrs4GOPqLHUeOr7kC3xf12LfnqH+0+2nUVTpUnlxf35o83Ng7
58XMGi1miqQNL41GhfhbSgaNDfszbJxoZyTRqvnCpCGvsE0fYQGlF2NLYGENaBsU
VMP/wz7Q/+fQpzT7QJL0tow95NnNeb7xGA1FfckqseyVtDuhAEgHD6mwpVmQh8un
elIvtcNPV3FahETwbYxZ5HjkzBt2W3HFmW3IIWoPJNLB80RVqtFUc4ZU3nIc4VEc
iG3S1rRXFD7xV88so6IWlXOwnSKppl6RqT4d/KZfltBGVR8hnKH9Vhk/GRz7ER3E
YnrXPaW4mPb9YwmBnrkzynrIGwT+exlNPOMqKjAtdWlnpXs8Uh7X+QlG7RAmBt4r
OJgjZR/tKHiHMODXaBiYzhmwZ3M3l+orOAfq3JI+p7plSjBZ5J6Txwwqp3S/xGua
RKtVSabY3y6FFjbBj1vow/YSlZvPp4EGWLlKO8jqTgq3C4a4P6thgOiYYKgrafy/
v1dKmAUuun91uw8HucuSEJUUxMcoAOSQ7XiBQTGaMJ62JELHSS6dUPVUxu4MB//a
w6SKvi/Nrhy+v1VRBPRqfciRGTi4A2yfihffHwEQLfCUw5qRNW7uHoslAYw4+5OP
9yb48qgpcTnH6yMlySGRCzm6YjyuT7hXv2qkctxw7oz+I38vLntc74eIMiCqdc1+
52eVhNQ/FNJuYPHq/BUHgC2q+MTQmihEDazDJESyGuMZ0ZYCWvbakTNRj/5ieKRv
jh4QO053xdg2ihGysKdpcdsuAKANExcaqfmpD6+P44oLMh7xvAhmBGkD1qz4ssZ4
U84u7i5V5c3WFikvsPEtWGv6vgVH21Tf5QitPsYgtFvOeyMaODOlr2XE40ZDqYHg
3VXa9+yJAKWapHhD7a1FVp1exP+t/c+maLIO7NCdGrdIz5TPYvIu4sqs1Q/jKQqB
0QOQ6rcM6WbU/wFBacRQlzZuZavOsM5fl2jhrGRvHEu56UN1L6rIcFeunyRmjteK
/nF2/qkAALoEcCSELWH/OrN+cQdaQrjao6O5uvE4rFODeD6CNPx8Aw8VnliIm0U+
Fl2fD/WJE1wiTD5DKqODDq7ZAvrftfITfULuYLigZT60Y6TQz1QlaeJQqaUC9uAE
8GA4HqRG9gB9cHiyagmC/Q==
`protect END_PROTECTED
