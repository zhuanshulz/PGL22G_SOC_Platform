`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oxNOHD6N5evgeWSQojQzMka9HwEUFFOC9sDc+c83C+nPhC6v1SfibimmNnPg1dZ3
i7e62gmbqf+LUtB6jMw+zWqjRFzrmkqvua1oR6yRSpHGZW0XhoAw4iTbs75SjR26
hE+yYRcC17lMMJhwUqhP9G/JdUEFehgvlLmfp34UnTbCR4MU4rs1mZsd4SY7ioRi
CTmEJoTnoWdI6OixZTsePiN4mYfWcOmuO8oSd9Pa5LNAYOHRyKXePhXvIzOoOMVo
RysWweiMHHdoNT7IZi6EGRGn41PD4zMxEW6CimNN5Ih5BGq48eEFbmWxLx/SOxxs
KR4vlsVSoF3Yjksn8v8Wapwoh47hU6yPWmZIflUuRzjDlM1pAND+fW6XfYZV/Oo9
fITPCEv085Er5ZH9vhO9ujrOUi9NcLWDVp0VuW+5azenhUa3wI4QdMrpvAlHh8Gi
JKQF7w6/RjEGcWV+DSy8aKJ0++kyz8ep2MBCNYDxC+04SKR9T1avWp8985MOR63W
/GdNDzvogqz5wrW2JwfgP91Id4SqXuLC2hGdiofFhPuwxDLUCxTWJhb/MCpslOCu
AuhZR4t9YoZC3NUTvJ/Ja9eLBKHHTAadgN0hmnv/2T78IL3+8VgzEYqYEU8sQDNl
+7aKw5AVRb+P82coir1JocqC/O3cXra3pVl4A6Wlb9fR280HDfbG81RfHm/T82tn
dPTFsBQMSKLx8FPsDSoWg/JzXiFxFhxm12Gl2dYHsg95jA0/f0n6Ls4092m6FOcQ
tAtWk/vW3pHJnJg7GWxucd6JmIVNLuH6rvTNQoWENeFBD2mF2VfaRWUCWkVovjJh
kFzn8UCOZHQcbogpm+qMFJj2NKukqaIlyTsPXsdtHHtThi9as8TmIDw9ZYN4tNjn
`protect END_PROTECTED
