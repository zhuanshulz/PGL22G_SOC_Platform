`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cSmkaHnX8SUo7yxl4oVjwI1eUE6tPgIbXtXtz0M1MjQdJwaiCego/nhmTi/5KTv+
3ufAUJ1w60NmOTu0McEI93/ZbkZ/IZT9eIp9vIceRRPB1ekMD0B70RXSfUoN+M2d
/JMxSDFKmd6J0oUtyeJZBEgWPtktOb/aXDN+ZUgLEmoCmGFwMMKoZlCrdK9MrslP
bzSyrUj9TOb4rEHqlN2vsmRM4SJhOH1Pt6sJtclUAQqvwVmedz+DH8OdfO/MYv9H
NTIUQp1FvT6E++Ryri0CMFfS06RpP7nXy0a57fYlGBSWUqhVQNfIw+cvu/BjMrrK
G51VFX+zcvNwk3e8BYZrTjgJyiXxY0//4Ju/bEtfF9yPm/k/OYItCo4Et9eEZbx5
h9b8+EGrqsSnX+dA68Mann3lrDdAeInVmkWwcDG275Nvnhhfl4kxet9H6t/CZT6X
J+QlY69+VhcOCJf7cictnvxMqtl8toxitPzGVO0TFBb/3i+fP+xdN0rMJjvGG6xd
wakJa2ppjL+MpysBXAg1lbqxhjRX8Dc21E/cAIbbxXw=
`protect END_PROTECTED
