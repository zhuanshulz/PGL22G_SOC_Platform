`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rufwdbpojKq7hcN/ACBOKjSY6ezJ2oYilL//OjG+bb/dsxVniWCgUCl0iQZMVJ4K
sjEru2yvR+jPRbTRph48b45s5/o0rmH17hyoaDN6yJqjlt2Ksi3rpiaD8EKN0/Hs
MPlcBbGEKu7IzoYhCMaaNgUtI1BPmQOXaY4SJvbU1CNfg+RKUlbTVpw8WVfBh4+v
yK7G4IN+GqlaFXyAb0CqG2hziuX5op2WFBH5LAtq/PqnAIy3Cjypxg+QgiPp196o
PuMO32itvFYLofTKWz8KtxQALv5Nrix+hKakrXcTRnNdZ7Qvf5fA35atKvjyzvxx
q1P+WCuONszjOwsYeYPm9ubQcr3AOE/jHqIFywR3DMhmPH/N0gnNRctH6lHPdhMX
3QDIl1ISfiBn44YH/djdQm+hgf7ud2qB8fwdjiy2J3HduAvRdMVn1GSrwi/r7LEf
sugoAL2w2ZC5D2gWrhfApw==
`protect END_PROTECTED
