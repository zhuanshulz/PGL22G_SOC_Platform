`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pT/1Y/rcY7M1KMr+aTz9irVnfn0Bd/XqYYl6xw2/9MtzmDOJIBsjQLMuNArAX1HY
ZW2SuF8P/5dL7ommr3OR8ahiKY4NDm3q9NKt9oQMOca0cPJ6+y1uKCQ60UxWwDxy
LmBbOvwN6TdbJ/kTlP/VT9ZMic3eAHYlnOIuN0N8KSeFRk7CoYub/HVO5FVJZUdH
BM2mFSpG3fdSki6F50AmD+djtDc3eZ+i/5OYCLIuZC1YQ3Kzj8LgkSim77ur7mAX
IRFQ4rSofsYGIQDn8rTvEYSA7NUw5I3vkN/IJP00Qy7qcAiX+rpp7q2qvMZaMvmU
R/nuo3uHDLIctUFl+Ry9VrBNluN63WdwBzNJurpn60CsoThkkoaTl+/VvEB00jPb
g98rLsoZEDA0ZVW+aG4/lLMHNcGPLYnwnmjwY+J5eb7eWHqCfWJKMhlCPM5f4Me/
sjfhPhNvGaCBFajQeNzmnBWyr73ja2CszbdvP4+Dd6wLFm/ZfkP+W4R8QK2iGmA+
b2GvNWrMkUX62WpDV6VwPMDchcG9K3fYzPEnyFkjlCkQnyoeJXpeOdAOcc+NzgZ9
vFE4dVYZP73tjc0AcaXTYj/NElXksGC54ozUj/sMFa48d5bCZXWhTN51P8kDKRbv
A48wmYd0KG8PexW1WjhnZA==
`protect END_PROTECTED
