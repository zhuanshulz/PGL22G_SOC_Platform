`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yxPG0956mmBjCWVN6jfA+NILaKltx8UpaATDPz2KiDC/qz1ZPSwPdFKYJKJgEnzE
kGSheab6vO2jTd0PY4zsJZ7cC0PVtjJhQrg16HbkBqnunudDgTV/0iG4GHh9bn3H
B3kRLiR/Ho5PmtFmQvTsDG+f2XWUu13zYG1RZV1syz2M2zGOPZ0fz5gwWkLGKkyt
T8ulyLX2dOmhLvZCC17qkIQ1qYWSfiR3NmmOBCq49N1O4M23wFSn9C41ZLxcSSUf
BsicLed35WBzU+HGASXop7+Oqi0VP9HQZXiFXO1WzBJRecGVHnLEAYz3GmQvJ9q/
Z7AAtjEyRJGygC0ty2RGTlOqiKeZiB9bxj+IPSEm6DXGxZu/bOrSiZxLNRN6BbIm
Txq7h8sMXRLGpJQ5crCQ6DqgDgQFPW1K+dV5ZtPSdTcvmMTdIQnj0U4be15xtkPP
Lda4feWmHHJec/+/NaktUhUWwnbZavqQGQ5yJeTmn7UANkn0P9o3UDbmfOntq/pn
4DDPSxJ432wAbSengJLVbA==
`protect END_PROTECTED
