`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sCX1hYr369wX6PX/Jp74of5RYrVbjHhtoO8sL0Mv2FRJKWARzHsJw+9TxNMLkkZE
x6GdgQ7MRj+jeoL3UvrT8bJ3Pv+bugdkrg0UOKk0gSGulsmIj+RycKzoWu1BdkHK
ddTDZ/FA5sPvjuyeflzbrCOTecjLo6j+supgozhl3WREWlGxnuiNuOPdGz+ytneh
zY1g88rdUS3M15TR96bj/3H/A1/XG8kUowXYEUC+ct//Jy5owMKr4PASu3Hbqq5l
x7mDvxEktNSi2Hw+wUVizg9kawBXnR+lkkus3y1vdNAptjLzXcV5UlG0C31DJ6ft
K5zOWe4vfGi+F+751qz5dMdtQayBFNVLePcWMF0j61PSlJ7sbqNPKY6zGkzGgpFz
vpgFaw8VECPx/nTyf4t/dQ==
`protect END_PROTECTED
