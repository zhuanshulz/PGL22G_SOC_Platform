`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jeeoaA8zuet+7Uhu7FwKPIVBhSVsfSrad65fe6dI9i8CCHNMqhHk0qaJDYC9zyS3
CwHKx0PJcoqNyCgT1CfHLy19gOvYcncNDGpfbYAyWWfuiOacW4wdXTGkSuOOQycb
CaEWqfHF3cMymb+yW+w0/3fI4E8zrr6wnX0ZFC4JM1LuxUvhiRmzGz7NQ8NxHYCX
KWkmQFbdRWG9JEORd74kPgy8WlG27xB4sNtm1eNIpyHTBqX/13Xtd1epdhFoNL3t
Dp31Ib9U8CX8dtxCfQyXozwio+MSnsOCE1RO/4IYZLo18i3p37S9W7i15jepcwa9
77/gP1FPhy8mMD/Q+xgmg2Zc6Mtq+D+DmZoBWQLwloj09RUApRhqTM3xE9bDYY0A
BEfSkuHqDO3DKsK3yRGHQguVLI/cdQSNSHwL+hEOWGYB93oCgNowsy1hTNomH5RF
rRmHmg8Bb8Eva9kYelXFBw==
`protect END_PROTECTED
