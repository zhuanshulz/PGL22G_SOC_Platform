`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OcCB1CJ7h+buXkpROvHml3UwHJTgFzbviTFieFiVVz+U73BtB1/D/1bOBuJM6GDu
7JaoTG9mbIPIUv0MRL810OiC/tHz/N3qyDVkQbDj5sQD+BeaOr/ojWar4rqc806P
gQdH7rhWlP38qd5q/uAWlJpojDmKW4+T6hcZg1sCDixHPcR+NZLbkZoFte/dq6p9
Kg/jx3bjuwML/dzX/IJlxOrlD84Fg+4+0FNHP8qklGH5Gj9dlHEyc53oV0TqGesv
DAvyzyNWPZg+MbAdDf9Xohg4lItuh9vFexnweMhP+34C4LeGDpqDvIUfPPHgz3rA
KHGaegd8GdDHi/IhkwC0fXdr63gnd9lw7EI36wryMxmhFtPB+EnyiRnW8zhCFkFf
zpfP5ez42yXfxnpBDFWkyjA+aaFDPxK/RWaL5HhafszPGRivvz+vFn0TBPRTcxN2
pUVXOiE2jx01Qney4Aww8XblpS4kbqwlx2GlRgGLEW7LB3K6He0r6RyjRZqKvXeS
Qy4cUp7BapkOVLQJQ9ol2dIhTKUfQSdvEZG33YAjNDMaDr/+4UYVzpV/q8tvSl/6
7H/Uac4kTqKIdFUGzAc+2PvgyjiAWGI7pcGyxRJtm0P19tRQadzSqRGF0PWZgncB
uvNZwe5WrDQc0gE/k6WoJylTua+QCkgHdhrKfJfk93f84yTwkLTBO6qTAkqL7A4W
yQwSU/35x2HJx/vZXuaufqtQUAPTB0HMHVAOzQ6NSJtoSmbAQGrHLpZ/2R0SS7X/
BBcwpxmrPcjbV7Fn5WWIewqdaNoZvDQZN5zcL4CGdYPPuussTDVAdHgvVIc24uQ3
v/7i7MAkGQgm1YQBsyAFZfXUDnWVGxpjH7Tmc7EtFSyIEaiKjt9/zgnt07L2gCc1
vGomJPLuJ9X41HiBYXrmzZpXEzPl2xyU4T37TzX702TmhucJl8DuitDEe3QIomg8
EZwMjcZeykROcIxqlaHmiqKVgiG/MpKFRhtrNe/CBz0bYOl+RJt1q8ulR1RuTGfc
cf47irFz/pSi3e+JAkRL/Q==
`protect END_PROTECTED
