`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qSbtqG6x3C077We+pGBdP9J/5WODs3ejiqOkIksqzhH0RWU7j0EYtdg08AjMmE+j
NNJMQi1ZeUCp3YnhP09bI2TpkX7kxr8pwJI5AGQ4rhWc/N1zQFHwsvYAPh23ldOC
5nQhyJ/jXnLkoSuE+rC1yPvdnSsyL9TjITEiAP94IAkInKq0dnDvAuEYVQEvKoGN
Bry6gmSHyC/iKlj/CGXCqXGIASid66op0gw16zWJi94HRdUD7RReGA5cpeCjvaCz
Ge2xvwe247rMMQFT0h+HCsi1FOFlj2gUgRnK/tY3ysbshDl3h/EtVDcNVOAPusO+
lggDx85K9ad0vA9TOeG2XUJXmU5Acd+3aEvOcJbJgd5BSnf7wH/PdknH0abP0l2k
NjLFiaKxPDt84JQ21fQKeTc71VrXH7CI22WQq+x1uVdNIuPPIxzcdTV2+DhqcYLf
fah7kr12PPyMqrDJMZ2mgsujNF5xsrm+CnO3eZPruTjqUGuSkJ5u43x/E5igL2dr
`protect END_PROTECTED
