`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6rGOiSfblCJjIvM4M68lE533CwhG1c5StZKQr4O1o39oOg+TAvaEb8ebxrcU/VJe
ztDLv0RNVvKsF2Z0ddWTiqp8fDLpvSzF1Qxn8NgyIJ9mt0n2bH+CR4VbrrIzCEBc
LNT4M3u3I4f5TrKeQ/Uc70AShmKsLQrKoyoRi3unAcJONIhFmPjd1QB2gAHjNXrv
u6+n4Ilf4zXQ2KQ5xwhTkZ+mEtWHLv3IMO8k1oTqfNslwX4jozuj69amOz96wcsG
iqF4zz4KCdE3/AcSd8OBHCKiNh7DJTYGvRzM6JZJNzB9N6LsHu7wN52/1cDeqSKz
3xlFJQ8VxecebUn5Q/dc8R/vAKA7X2c/1TFZ4HTcTVo=
`protect END_PROTECTED
