`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3Mw5rlUZtp6rgV/iNd2P6k88sseYvLGDJeYfNg8n04q8fzqygl356DDlPfasaNlb
ekYiuMAitcqBadJaMxkBXigiAGrMzlG1CQnhHPJKOWDQL57YUdrlXcjQBBB2+k1E
48BWDp7DjifoUjSbB7tvHNDyngUHC4Am02lfY142KV+Zw4uPphLBWmEHtRnrm/Lx
mSlvukmYcHir0GPgqiYWxLVONDdQPX3b4fViCBM3ZhraAl63j85Kb9LTfjuujgg8
`protect END_PROTECTED
