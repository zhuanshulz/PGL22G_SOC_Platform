`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ndUbvUyLY//TNEvgAZbfunE/+1lWsqNtvvaKfpbxhuN75TrxLMt6dFAjsOuwQxRG
qOgaEvz3y3T0kiwlpKGNrDn/1r9KbUN0fDbmj1U58Pi95hJBLCU50kMR0E31cj+h
7Nx5EAUusTwWCJJ+khhLBBCGUXD89WLCTxlhxVcOY6mCALRtXS3dvXDiCg/8jAX2
aXkRXYOosB+ubaMw/oLMj8JAsUxws4X4ARLoJ1ryExmfDPXrCYT8sqRBRAQDbdQE
yjiUuWaCp7u6916pHTcImDA+QqIpM2su0VVnBc49keZGjAnwAT1a0j2JaALLKyRy
Y7sF6l7KGpmkpOJd9pR4SjDT6hKSzqpvuHr/zF+rsSA24/pZwHIaVDjwDskn8KDb
cCMAZ92CHkaPVBi4DumkUz7AwHvjwDZlLG+NtQxg+wa7rQSkLvEamxEHMDrEWrFt
pZqRZ4EJ0Tjt3fsjWt7npxmNAyTLXhcfDL956sBS79f652sbcEGKtx2vPfjAkT37
SpHWRfA2Bl2DxlHTlPVw/BWd9DX2c4+C9Q17PIhmMpHrZU+mTNaG18Dh3MSHSn0V
dAmLBKt94r21Xo2WE/tbVoKD5RT1h0B2jWeYpVdw0ny/mpGMQ687jmrcUykVcONW
ASLTGdv5Kn/499CArITfvBp6jLtgmI6GQXX6STjgU321FvrUor5jumUQKT3pycYa
cjlCYLDTVAyscnuaDeqJZIfpyb/hOlEa7v3iOHPsfMCrLrrvzM65I6y+DIPBS7Z/
49c1hRe+gt/hOjxnZZ/8HaR5nbHEQBMCWm+rX+nEtE4RE949PeePoKk3OfyFtjF0
I1y3oD8Yewe69waIwttNQN5Q1cpJejZs0gI9F4ziEyUcFrlwa87KBOCAKFpa+FPZ
XBXPk3xCmPuWLsmQKa8Q1OJxhbpOxvAjlgFpiRbcBF++Q/uo/PkMmXhrZ8V6Lzqe
V7zqHYK6aLD8BuTBzDMFHKGiD2S/Jdo98VqQlS9Tg8mie8cK+gl4cm03GjGrT7JO
qn2NLEKl2Q1/cvjk+OFgzDOtoWT/6nmpPooUVbBE28BNeiPXDzGixNm4rMW6rVJm
B6GYfqbJsM4zmjgo4qhgnQT5mQEd63aHk/rf0LsEiD0/HGxbpc9qgfJg2f1rQA1t
oo9+IQASggh+hmwGF0E0oDa33X1GfTZEWGeWrHuAXVxUsP2DE8ENnRuk6sMLjtFN
O/Dav0HLJwhGBP/EYvKgTLmgFU8KAmWtBHTy82K65X5TKotCZRZU+oP+KFONBzqM
tUO5zuHF2tRANo0OqPTJSv4D42HVY8ZD0P85Kb+8+37dBDlXpdXQ3Tc/TW4R7Djb
4wa56QPs0Hd2Dt1AVV51+9t4sD+r8I8uw94chhhl2cjxUg0O+1BLeQN1IdRtD4/m
awY1fBFH6FHLj8oUX2oTaZ3x5Fr/WEG4vRvwYHG4HHIkn5Pfu5pxkwcby19mpPcr
Bco8I7fWuNvLkjl+i6bZix2nC4WM0EWXC8Kdn3Bq4u+9NGcZYCGodsIyVIqessqo
fqe/X8kd84tN+3ENz0RT9V9PzkWaWBeMcdVXMSU0NDWhaF6vvTLj3ixmIKyohC7T
2FDCV65OfpVPjr9ILqzTSu0gocz3ZjhKYieI/3SBN4Nk4gdI0pNymHlew4ZuN0Em
JzXYzoKpg/uL8JcXxB4b39VdgRTgyhkuHlJdCLR7BaBPKDa90PBV5zh1LjVEIhx2
UI7v0u63esqgOG74EFMwih8e75/If2xzzOrta7xMJ6ZyHXy5tRH933YA4wri953a
yzj5eUSR8ZmPD3SDm+aBjAC5JPP/yAFsktl6dL9PT8g5K5o4dbBoCSpMZmaZYQme
K/hHdHC5wZ1fR8JvfTZlD5x/XRIu0AQ/K4C74tzIxK7EccafppR4UsbsikgXTv/V
3DT/KNjXC84C6HNzvRIIEM5pdJSRDeZomNpdOOVPQm94u+gCZn57hJHtmaNegMhT
Fgav0BmdYbE7uBBb14dzu2dA1yC0bcb3Rq1K+q3B08Ew7fXf9Z5V9o9Mkcb8LCV0
/mE0d3CrISvFHd4sTCuJIwoQrp6yHAkoZzoDYmKL+jhJmQJSWeT/l84BgEE0dHGU
mjhTe1vrDkZ8vlsdwTvn3wAv1nrRzwdupxDHThTfzsCRPp+0piOzZgK+r+mjxXh2
7WP+pdggFWWI8mHOLStm1IATMtLa65rotdKkmXOURqFKEdiOTY2ceGCConGrqQG9
c+cXVNIqM51nw9Hr/uHBfgJEeb3mek3posKPnsYEzjNDBU4rd5oDvXewJJyLP2Bz
aFX353foCRFQp67f5lNG3/cwTO3I3IqZmsK9B6ofLEV8Tm0W3ExoLlmw6Y6wssvu
cOBQTCyW56SqNPLA+oU9YLKiaVzsaUmKmNclQ9y6QeP1TVeQYGELxz2j+KBf30vp
HdstpdtER978DXguTsYevUsA3a1zpUOfrXY/xGNVp4RHvhjffu/ZcexnsfRfdscd
jtoOEnrPsJBkLqv83SgT6wEPtAW9FEeODoJbj1w9QiaplbR2ej22KkGxtShEKtui
HtsAPQgAImvH8nXqqY3YEDJ2HfdB1KzPn7I9cXgr5L0bkfad1prSGkENjV5IsC5w
n1Uz5CrWsV8NolPTA4diovI/flQag5agqe2Fkqu96F/JBAsHjCukYXUI8ZHn3tDF
bpYiq+hpNWZxtbCgCmgNDslM6qWk3+Wy8bx0ZxADzFnTe+qYjyCPW9fixFR7sjdU
I5bGZf1G63/5tfz1RBUiNgyizGHystVY0VNVOng8g/ZQgVkTiXjcKyZdYus5/nQu
dKqmVR9QO/mYEI9jYLvbZ3oBkXt37Ie9PKvDg1vdZAoHRz7LoLiPVaTDFConQhCw
tBBoCAsUSnGbEFaJsNvuCUev+2J0kbg7iqF1YQJHXMdpr3Ia91h3rUVkcim1Wl8h
RM8yq/y4NjY9LyCrGBtVctjHQFZZA9tJekO8h0JV72fHnnAMXrlZXm4+O/9bpiHa
ellpRflde55NKkagLQws1JVLPdUNsYuMxodYnq/GGdFVKky4lFRZYum/Y6CYxHAx
jMBHQDrRrbe6cHMZ4gGg6zwl6lI/xchWtAx8KHJYSuDq0PALa76QVYGeDwsFQINL
MSoFRUkcHLDiokli6f7NL9UXUdrYBHku5eSj3B+gO8M2QGiPNJMvxo6RjH3zbFU3
XO77P8FRvlCPA1bcbKyjOX+ph1bv+8aR/hrcxrC1lMRbzLeYIPZX91cEPBmgNmTn
`protect END_PROTECTED
