`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mkfe0bW5HOctRVFNhJoXKbKeyKBGaaXfrRjv3gao63p/ga7F8szTnewLl0fzzc9X
EbNZhLvaHM8ONRHlcKCTExWX7xvca6hKv8h9jbsBNCBaIISM0F1dQYA/7p8zRQ1W
MxDoReIGWDmIaep7ehw/DgwcwHC3VlNgSmp/hp7jOWaHLKm5FzaPdvSFz7AzPUYT
iquRQADIR9HE5F8LnkWafQenH9yl7TSqqkD7Rv6k8KUXTbs5rfFkhvvLOpxyw5Th
/BlSQC/jGskQru0n7Yp7HgDCRwscY45aglLWf3GCw641h8AWY7tmgDMsCgM+PLts
yx0Ua3idjvh8VCoKVPmX8YNKis2KKELqkbaBeiMxwGOdg0lX6pxwsA3NELXiVB6S
KOJ35aewkqX5z4y2NNeiewNoU+bkecMUvQM6FbDewTZCBJJA5WKy/DKXgF168ZKm
bTIMzlphvCXy8QutLKtBzifxEJ+xnsIDZ1585VESX+5KRMbv27e3oluSqN3qWj+G
1RB2pab606WJAt/g6YUDj0CFjcdwWvlmmz3imLwB1jz+w8EhLQpY9EwPy2uxxDZ9
+WXahIRRxpQjVWcq8Ee5GOOfuHNCwj5KlYaeZcUiIC8o+4PKt/24f6ex/Giu+JOw
fijebKJb1i963r1Spjk7RSyMqmyspOvBtWGTYGzi0M7RPUsdvcs8qccti0v9sjcB
KfOa62Wbi5kfgSe1SNMUleZJCNEuvZhw7c098UphPXqyX5ybeKQdzLtNtfA1ge4J
PZAK1GhgQUi02GX2EevYKbqlEvhsLvfBFbFFGP9nQz8fwEkIrlp4xKTpQG3jLmYA
`protect END_PROTECTED
