`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eU5MpJ1D5fEC4cw88v+nXCZF9YSjaAA4zWnd8HPM/hrI35+VjVHbEz6kalJrIlxq
a68qNWr+LCGu2mBA4J6xYD4SC5GAC8wOAm78c7y3DSkhrqo7t4FVcXeLZlFFpKVq
kGb4y2D9OR1Ic6LD8KY97M+W/JZdqCfMM5hmlMIwZzPbLOPNw90djAaCVAJ/FhSc
4GQgGfQni2l7/amurgpvNOkVLtZVDmMwbGncRLsaCNLDYYed/rJpyqkzqaomoNgI
BSFYVw+UHeGI3IDiqiXMI+wkuN5/nTA7A5NVAT5DYpuzwdUssLD0C7zzWRJ2GZEi
Th4m2Jmi5qFwluk0a2SQLhoGMokmMK/hu2gW3tb8d8oBBuGXOFzxZahMzs68evPR
JZ58BXiA4E2z9ssYgxdaKzTiB56V/WX0P6FVNcBME2LeLGbSIsm01bLqVhvUN6oH
ThV+J3LddO/20sYYug8pz8nlh0No8OFSh3/w6t13pZDRmIx8TpQ1WPqMFNk33t38
uly/GjAwQtPn13oDmplatWW5LC7jH0diVuVteErbTlHEqzuzPMpZpucG8RhvLv06
P57KV8C5cLxxZyLMiW1e7C2kpVMf1RXUTZOksMlOb2TEuujtwbpnibyVAGF6qggY
BtZG9VjKPMlo2OXN3a029tY//cS/94zgXDjrpBTxZgZGN2FHhvAbgclJLGBM7/in
Ky5OdVj0iyZNKDBjx7q1mpsAfOThA2XeVob+wU/iSzgB7DSmtF//6dKcm7G+D58m
f96QV8rImna/15zgNv+L8Njonvd/0KxgkVYRFM+oOrwpRwhRsFlbYGq6NO9FYLG5
TgwqSp+adVD7V83MgPOBD6GVgigqC6PSqr4Rd2Wq31EU+O5DEkO/X5HmRJ283cKy
44gCrNSYJGvPyPa0BgorgYHEKvfaXiVVFaXkLpLzrsCOouqqAVEjjX6MgYYSi0cs
VtqV8K1Wu5V96iPB4tVwNgUzs6Xihu9/gytkToRtZ2C+mG55FyGyT7LD//lGe1rK
Kli6NFYVesLBXkpbjbDvGHbE9/BUf1bp5Et1e24PL0gMdq5VErN7jXGWCXjeZvpl
vNbHHyWqHfIgb9tHbptvK5SM1P49JiMHpMuaQCmSzEhh2sKrqJdfOSWpo2bUmmCy
q1TQfrPy5MCQop5RhW5G2mOsmosppOb4mXyGd5lTHThhUKSDmbJRqC774jjETgp2
Eel5+AC4uiCGgzBZEXGhrk9Mg6HjNUINUnwAfwfKZcPAMa+VHGObMbllensbBSaq
PBx0+sketVMnruh0L9cWgYgm8U/bEcEzNrCbB5yjJVE9rOj8icr5eer2T64X+E+I
gRqF0ewLug21fs4epOZv+XBcQao0hkwOT0LrYOAFSA65XxbGIb30iTAPi4ewi5+r
7383VkYOIrIMsVi06+Eo6q8yb9wBL5DscwudqiT6vieGpbWEKPLsj7qtmseFBK3h
vuEO3X2SnW+TFiaemuLNHjonFBvsiDQKw/vovgrMx5R9d+drLm3il1GzrmLS6tn0
pU5UnGr0cW2XSnn3rcI8fv/5qYHJIZW9FFVlmFMiP9zz6jM/g0nCPIzWRNp4JEtx
xrFrFulsc0sHrhEximffZSlOFisST0WS4pVcUorKVngqSVX+QFeqlmRDiz4OfCln
i9LLXHLE+11w96wzOzkrAhevzcZohzGo0+RniuAi9sSFQYBI2/iYYI+hAaZRNMY4
z2IPJRRDbWoaNjcLd67TqakgJsfJy152EOuZw0+vuJzeXBZ3OES7EkMJGpB8gxgX
0jyYrATF7HyTn7JrxF/iR7GGFcXYFDYR+TmUsxaTultL5QPbotlc10g0D+SKjjkZ
N7LQjH/L1xDeozWU1u3TNaYkcfjBgy2DQotC+Yjg9DDK/LhmcNfRHcXZ/FDGOR6g
10vE+zZsLvU7EwO2z9VefTf4NaQzsAsYyt2HDXiW0vPz80Husd1sTM5iNwnvUl9A
MEm7u8VkCJMIX02/TlTsK/J3rtNOjqRpQBTnpNLI1R7nj6+xJN3k3KsSnfcykinS
2YsrDOUYforLGhhbg+OwDeNxZ3QTujV+pOQCj1IiOzWMmeHMlLE83ePka3QOCIoE
eNwQFadZ3aUp/vi0oa588g1FQ83sePJl4enANnR3tNj4AU6l8+yPBlUw7yVavBjk
AXaAJrfHGC4TNsZ54Vho/Hww+OFoXYdnYJg6QVQIAGj6Ug4JJcAms4O/QgPMH6+U
OYlaKz5lnyq50o+o49REtUlEHvXyTgWuF7A19LVNzXoF2uCamo+r3A3yNW9Bixji
ImYQ2NJImjoc8cw+Pt9ybR6dzPTPNrOZE5pgTRf8TPWXrtbudfkj+ALNh8Jjo2sJ
YwrPabIx+c3ZejGL2D3efpqn9lnlU7BFyP9QuJV3xBwxt6mit/dkFE4FWK+WeqCc
RiAoiZy7nUSKT4URliFHJL3UN+LGKEWHT8r+46pW/d2hoGgnvm5nvk5aR9v+mO0X
X1ldBDYG7RcKEkFkU6SNNoVn47FZW26IaKtZsumfsE2M4GrHEovtby2XcGZ49n0x
fDRWT962tkB0OSqwFGnrQYmQtpveFrYIZaGiGYatjoW5OoegoADEBRj4bsownsUk
p6wpV3HQ72odeD0HnLSNQ8ifBuCE36QLJnFvMO2DuC7QM3HRfcmrGzsPSC7a5Dp2
spH0M3B5qjWVuq6Zm5HX6Z1G62qi3rgNa1EvGZ5vkm0kaQJ+TisGooA3BONC7fS+
flveBRNHm3cn8/xWCo/xshkq0TnegZ9zqB9CaWupiJJ6oHPtFxZj89R8YwNjHP2H
WnNs4XaC16Rv6NWj3zkDMcS07LYavyOGpAFojUzv7sQRgcIxH0URTwAH2K0CgOJf
yiYW/yX/mo4sYzZZFgyLXeCz5axxM1Sk6UFjuIbAGURpG2Lto3pXI70WdZjN97px
Jv4V8lNFtDCY/CoYCUieAGfIgKVECbScSLj+RW+Eiy/mxwBBNSjLg/Xy/zBQjVY0
Xav/axXxxK8G4ZAgH9W2t22qsb7LzgZ9GxyN9RKlpvl5N8M+tbCjkrgpMHc05EjS
HQ3ESUrT4bDdikmg4HDJVcu1yjTYT7eiagz7E0hvx7fiMXBAkiYBSW553e4x8kNP
FrKlH8a0fHCi1Ecp2FNonK2Yh9LKKoZBDNLATa3uipCtLufpifRRIBHHLQ1XDakO
7bvInLZJdr/GzqmfxKwO2vVKk9wzREi5MItB/wDppUL2HVAa7JhH1S3zqcP17Dj/
1UEzBsP1rTu1qIRkJ2WTvCokSnkt/j5rsjjsI35ZttCaA7JVGKaLTV2lhhONbV7r
Ty2BHetfFLGzVcrEgUSPbHroqwBpSIspc0bkimy4xcSLVaWgIN9/ifHLyLiy2bDh
ndpqHaeFtnNTDbA33v896xWwkWh+MyQdCx8nT4inkG5hZXW4Z2elV3Hbsrov/v19
EgDu0RY0X2qbWHwXXDsYPaz00KQCOdKBT8JYZeSJhB3x02qqvlKIXFWzcMLz1NuS
PFqwblWFCRXthcUs621oNtzXMlMOxf1P2DV6cG8HBixHCeNfXKEd94UAswf1TQYB
evTMLEG1HAzLIlhs+XLrxAhFntfWsTP+8YDCP+USN8+j+pWqECydS/AjALM9b3w8
ZUXfnnm7XNh+WDqqvsnkJ7J6lXr7z1tyx6V7F43LiE0SMKAqnd6y9YjU5UMl8DsR
n+k91pwqleDXLCMWYt2ve5tIH1+Xw+tAAi7Zm7fmHdvvM94zEaujwMP+v68HYZan
F/5lOMoSHLtJig0lAjZpNgqYasx5BMNQtJVMokalO7B5hqshfmY/5yaEJ5/iUj+L
GOj2mocTTEzCdZog5itJ/6q/UzJZtpRDLwC0xEvq9EA3SgmyvYccyrG6WoylKNRo
j+nNs+RoMkavnT+kWXbP5LAveRFcI0hvU9+QZoeCcBBozyFP5fx4spr+H6G81NNj
BvFqAn6VRlZwcolQ5nCm+nl+GDLR0FErQLTw0+3b4JCZS1DkfKwIVwDQyJWSKEWa
EzSKqiv+IU3mD8yayiLEotDl2sr/Xxu7GuBJfC2u15uuwbMNiko4o1eXg7kP8iJ2
Q9Xr92H2on4JOHLpj8as2AUqHkanXAvqC9pmetzTpnTKMZj6C4R7gn5plY5p3nY9
38SNFhmW83ysm8O2ZXW9OWb+/cb8pA1FPpTtaa9+1Lh0t+nO8GyEGTAsjbT+jzoB
AmizN0TkXyMCqdcs+b77+B99qIrLwt9I7VshAZ7SlGabbG/pJ58gL2OHpdOmRDyF
plXbOQGiu8jH+yS/8ZCkVb5ibFO9EH3uEOHUWLgT6xhS25ox9t6rgqtQ29AGhVMF
`protect END_PROTECTED
