`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
88oNp6zHGGpXoPS1oxGkzvq+7e7DrBC75oGbr3Vz/4gi5NJTufGKPW/bu+oTE1RW
qyATJ28Ee+S48mYz71682MyQIgM5/5i+MC00qCL3ykkG1220pYRHcK6ondzrZFWm
ki7YhXo68FgAG+Fs8ejyq3sH8tbpHKr2EHXXMf2hrRu1yNNYR9VMlH1gH26nrbQ7
MkGIWQG+I3HyCI544U8P6/CNr/IybYC3qB+f+s1TCPDS1kxBCTK28SPyI0o/AbpO
Sd6jQoMhZzo9iIZ21nXHWxw3xNNK1fBqpKcXQNo1zP1dlU5JEcz2kdnVDloKj+TL
SGqN6c6Aoj5yaubUZkh9zUxwzkYPGamr8wg4oJs7n8oej2SmmWyUNQlaptAqWxKT
WYnF1OsWxGubjqvv8k1tVseIHQca+uOUsbd2gnp1cy7om/2RILr80R3CepG/8ho1
xra4cuwU/2Tek4VT0ggrex69iAfZBt6L12nT/YkgKqCcT3gl6IlNzhZ1FDSO3aUo
1Gt8SFlz85ZTFgOunPgVYEcmmlctRuPi1BI0uHDJEtbwk8HV2wS1ri9xsFaB5z+X
LAtKUIuNCVXw+5QVIQZWfLagky3BdAzlZMe5tMixD28p6p5SNfoBjbZPicb2ix23
aYInvuQLp7o8dAS1uw3RXqXFdtBRLaCa0JGsekmE1PY6PSdlOCiszlVD0vlJXNbL
6Gc3uvOjsLVzL5zzfoQz5c285ykRp6I7nh6XRaCumwmTU1YQEpwtWUGTq3gzW++v
Tk03c+AUFucIDc8F1kGbJJ2KUhtxhUznob5Qa9mItGYe9ychXvoyCDqyIudlj0C8
WvXmUwSXzIN0ZFaN3A96HLDHl7A0AxzGKWTTxjTDKJdW55K+C2+R4RL6SbvvJgHh
lS3KUCgBkEqq6dlCbzAbBW6CK06XMIEx+Z6xZQvXnOcI/nfO+Pmxm7Y+od3W8DHp
z4n4QogJZajrANFQMkWdqsJ6Bgr2biJ6OURFRZ2vTzpPqAvsFvv+mLKM/rbH0XAY
vS/+4ydUW239x1WA9HSrxQwLpDUrkeMeL0uHPjKUCZeLinXg49dzuF/POQy6wMAT
VrI3mQ9vJf2msWtZe47u/RJ8FHHl5h35FvpiC4UGyOqzA7Fh9V7cdKItayYK5fGN
`protect END_PROTECTED
