`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MEKlvSlDfOcDJBjsZUZt7vgqK/8l/pA9mBIrfh5m2vzw5AC5RBDInpBi5m3MdMM8
eB/rh6wSKN2dtL2hGujtVeYiPN3TYoxE7eH9bLg93I5V06L1KAMdYPLQ8gTD+nxm
0ZzDaJHF6rPIs5QmGxYLpZBdUySoUmyb97rBIgjZPUZutBVnRk49mmJl7Rnj6+d/
cIFxrCvEmkdNsdXWhC9HIONp0WKxq+5MVQKHpK3Fh8wyFQbqZrNXUOjeC4FLC0bb
AyeesEzmbYhIyc9lN2z+jSGxZ/oimGQKnMJFLIzcrvqQc0sKkJZAQ+FGxH69Gokv
qwAua4zgwiIO993MyS7vLPptRce9r2bPXx6odwqgW22IcCuXizH7wARxhUkc93/w
5tP8wfdsuF5lZ8Z09EjiF1zfRTP5TG7Q/RvsW0jFg/oU2NeD5nEwTXj+6ja5Q0lq
wzPZB1X6ncHWc+rGWA2VRgZNASoD0Fp4sowBuxubvvRTMPtYmftto7Db9kEq3ZJz
GpujpIv+gMwoKi1S5Y3PSxmumvqm8Q3cKy508PNe7pODOwrDnojwogIRmK0tqInw
p6DN/gi14sd4BRT0UnbyU3CkM54pRw9cgSJqsWIKWR+t1tyyhwU/mxtdTf0qgjUh
FR7sFaSVct4blikl2TVYBVvYIUOh+AmnJ0jRvSY93R2R1UpVNNI+GT90582vZZXy
1RGz6FbM5CaQpcO3Wf/FHciM2qQvius3aQX09I47qu9Nja+O7mkuprBbZKy8nkvr
LXQEYDD5stefuQ5d8BT9+IW0ws4aIRYUK/3xv38rDWUjcRUnt2hJLLVNRQ+1W+ux
FNWKZNKciArOBIzBexXrPSpLNF+g1gYNVznc3gPEhet6pjaAnD6DJTgtUD/hD8fr
bAxj859kgftbceytYDFSRr7Qwvk7VPLn2iiEOvuqIyk=
`protect END_PROTECTED
