library verilog;
use verilog.vl_types.all;
entity V_CGRA is
    port(
        TH_CGRA_CLK_IN  : in     vl_logic;
        TH_CGRA_RPU0_RSTN: in     vl_logic;
        TH_CGRA_RPU1_RSTN: in     vl_logic;
        TH_AXI_ACLK     : in     vl_logic;
        TH_AXI_ARESETN  : in     vl_logic;
        TH_AWADDR_IN    : in     vl_logic_vector(31 downto 0);
        TH_ARADDR_IN    : in     vl_logic_vector(31 downto 0);
        TH_WDATA_IN     : in     vl_logic_vector(255 downto 0);
        TH_AWVALID_IN   : in     vl_logic;
        TH_WLAST_IN     : in     vl_logic;
        TH_WVALID_IN    : in     vl_logic;
        TH_BREADY_IN    : in     vl_logic;
        TH_ARVALID_IN   : in     vl_logic;
        TH_RREADY_IN    : in     vl_logic;
        TH_AWBURST_IN   : in     vl_logic_vector(1 downto 0);
        TH_AWLOCK_IN    : in     vl_logic_vector(1 downto 0);
        TH_ARBURST_IN   : in     vl_logic_vector(1 downto 0);
        TH_ARLOCK_IN    : in     vl_logic_vector(1 downto 0);
        TH_AWSIZE_IN    : in     vl_logic_vector(2 downto 0);
        TH_AWPROT_IN    : in     vl_logic_vector(2 downto 0);
        TH_ARPROT_IN    : in     vl_logic_vector(2 downto 0);
        TH_AWCACHE_IN   : in     vl_logic_vector(3 downto 0);
        TH_ARCACHE_IN   : in     vl_logic_vector(3 downto 0);
        TH_ARSIZE_IN    : in     vl_logic_vector(2 downto 0);
        TH_AWID_IN      : in     vl_logic_vector(3 downto 0);
        TH_WID_IN       : in     vl_logic_vector(3 downto 0);
        TH_AWLEN_IN     : in     vl_logic_vector(3 downto 0);
        TH_WSTRB_IN     : in     vl_logic_vector(31 downto 0);
        TH_ARID_IN      : in     vl_logic_vector(3 downto 0);
        TH_ARLEN_IN     : in     vl_logic_vector(3 downto 0);
        TH_AWREADY_IN   : in     vl_logic;
        TH_WREADY_IN    : in     vl_logic;
        TH_BID_IN       : in     vl_logic_vector(3 downto 0);
        TH_BVALID_IN    : in     vl_logic;
        TH_BRESP_IN     : in     vl_logic_vector(1 downto 0);
        TH_ARREADY_IN   : in     vl_logic;
        TH_RID_IN       : in     vl_logic_vector(3 downto 0);
        TH_RVALID_IN    : in     vl_logic;
        TH_RLAST_IN     : in     vl_logic;
        TH_RDATA_IN     : in     vl_logic_vector(255 downto 0);
        TH_RRESP_IN     : in     vl_logic_vector(1 downto 0);
        TH_CGRA_CLK_OUT : out    vl_logic;
        TH_RDATA_OUT    : out    vl_logic_vector(255 downto 0);
        TH_BRESP_OUT    : out    vl_logic_vector(1 downto 0);
        TH_RRESP_OUT    : out    vl_logic_vector(1 downto 0);
        TH_BID_OUT      : out    vl_logic_vector(3 downto 0);
        TH_RID_OUT      : out    vl_logic_vector(3 downto 0);
        TH_AWREADY_OUT  : out    vl_logic;
        TH_WREADY_OUT   : out    vl_logic;
        TH_BVALID_OUT   : out    vl_logic;
        TH_ARREADY_OUT  : out    vl_logic;
        TH_RLAST_OUT    : out    vl_logic;
        TH_RVALID_OUT   : out    vl_logic;
        TH_AWID_OUT     : out    vl_logic_vector(3 downto 0);
        TH_AWVALID_OUT  : out    vl_logic;
        TH_AWADDR_OUT   : out    vl_logic_vector(31 downto 0);
        TH_AWLEN_OUT    : out    vl_logic_vector(3 downto 0);
        TH_AWSIZE_OUT   : out    vl_logic_vector(2 downto 0);
        TH_AWBURST_OUT  : out    vl_logic_vector(1 downto 0);
        TH_AWLOCK_OUT   : out    vl_logic_vector(1 downto 0);
        TH_AWCACHE_OUT  : out    vl_logic_vector(3 downto 0);
        TH_AWPROT_OUT   : out    vl_logic_vector(2 downto 0);
        TH_WID_OUT      : out    vl_logic_vector(3 downto 0);
        TH_WVALID_OUT   : out    vl_logic;
        TH_WLAST_OUT    : out    vl_logic;
        TH_WDATA_OUT    : out    vl_logic_vector(255 downto 0);
        TH_WSTRB_OUT    : out    vl_logic_vector(31 downto 0);
        TH_BREADY_OUT   : out    vl_logic;
        TH_ARID_OUT     : out    vl_logic_vector(3 downto 0);
        TH_ARVALID_OUT  : out    vl_logic;
        TH_ARADDR_OUT   : out    vl_logic_vector(31 downto 0);
        TH_ARLEN_OUT    : out    vl_logic_vector(3 downto 0);
        TH_ARSIZE_OUT   : out    vl_logic_vector(2 downto 0);
        TH_ARBURST_OUT  : out    vl_logic_vector(1 downto 0);
        TH_ARLOCK_OUT   : out    vl_logic_vector(1 downto 0);
        TH_ARCACHE_OUT  : out    vl_logic_vector(3 downto 0);
        TH_ARPROT_OUT   : out    vl_logic_vector(2 downto 0);
        TH_RREADY_OUT   : out    vl_logic;
        TH_CGRA_CACHE_FLUSH: in     vl_logic;
        TH_CGRA_RPU0_ICG_EN: in     vl_logic;
        TH_CGRA_RPU1_ICG_EN: in     vl_logic;
        TH_RPU_0_TRAP   : out    vl_logic;
        TH_RPU_1_TRAP   : out    vl_logic;
        TH_CGRA_PEA_ARRAY_START: in     vl_logic;
        TH_CGRA_PEA_ARRAY_FINISH: out    vl_logic;
        CGRA_LKDT       : out    vl_logic
    );
end V_CGRA;
