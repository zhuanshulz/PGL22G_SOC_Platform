`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z7qRxpiaZ7DOvqQIClPD3orxaNZqM9lFYzDTGBunybdZdiP0UAnHRGcTh43DyMbx
XH36miksONVjDWcL1xmCnlvqNqSvPy0+cOO0h9drbZMJdgN04YkRIK7FUOsdXWcs
dgm5ma5i4frumT4b+iot1TsKsP/VdcB1Kj4ZlSpiSl2Cd7tVd+MDtgFox8YxZ8SR
+caNutKq2y+zGdGbdAGV4VesLnv0wFA8s8lk3PzKUYKwx9i/GH7oFHapkJKD7eN/
O+on6MkRBoPT/9JhZR4ebv4INVJYk7zl21uuFZrd7lEBq7AwEfFR7ZPX53Wmo1ez
aCasYgzeuzhWd+sA8s29GQO/WpP0WRZgLQnJh/E1ms3eECOex084OeNdvlSSARL0
iWRXDJRNApi+N491DTLtv9C2k9mjdfFcfGJ2g6sk4USJvZkWFjgesVD7af3fLOHq
X73x3S7ndqYSZENvaBhu3d4JrA+IRGIPqbPhj85Xx6IvucSCYwDOdfF1ziJC8r/R
S5FB+hRCYiMh0uxYpeixYEWy35dxjNnDpkYfvtlpQODNJ5VWoiIgUKAgmJnsNMen
agjdQKUdHW55vyEGmw+tz4C/fYa4neCX3GRR/jVKwwwa7O/1W6FwxRSfUEBVI/Sj
+8CSnPHr1kQXcOkxnZNNERD5diWD78N/HWVMpNb5IPPM5VGBiVwvxAAQaCwMkQkw
AQrhByCBCdAbMsaISq9N+g==
`protect END_PROTECTED
