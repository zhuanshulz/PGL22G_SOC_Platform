`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ER4Uls/ehi9vR/PJL0xMQ8bC31ggTyjYZaosxbf8cxK7CKnDE8/NHFwOEp1HcCxb
lQomYHdq8drVw5s917Ssd5BEkHUoXBfveHO4Zp75+TxX8ClXmtvQohdIcRG7WnMg
TsZh3rmB5zb2np+sY+ZGNpS2tIj/dkfCuB+gGaIBGznL2DwQ/1uTQDVUxUKGDs4u
l2G8oxT9/gzu8UAHlcEATWO8tfxRif9Q/f1r1Ts5Ij2eHrcxyHdZ8WeQSbDuuFuJ
Bh2N3zbnTdHQkOc+lKHU8eUS7karTJpN97XHwH8aS/BOiSiGcr3zgdx6yPImrs5H
uTWpEQNqWr/gpl+vg1dmgvs+joQJinFYsSfk9DLN1KNXr4O78dIQll6AMygRcfWt
jHD7KpI6/giWc3sGuwcNYxpiwPs8OHVAHaFGvEAJFKEKrcEKkeUtqFPEseZOHGxL
CpDILuX0SC3UYtCaFeyil9No6zZuJd5iOiGPirrfTjAreu2IFDp0nmw5djiaL0j7
qfn8yCfcoY0pxukuR6BadcV2236VBV35htLZhJO6KAcId/54OhU5WlaDRbzbJ56r
opXvx4ediosDAebxpGxM852jbFPw8L8hBPLRQq5NYeBiy9PtFVG+03793O48RPg3
`protect END_PROTECTED
