`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3Jeyw/Ro9cVDPHJyNz6pitShChqggpmYhBBX5NEm5gOa5qcsMcl0n40d7URnK1un
cJ1VKUO4wgH+urPTLZgWKeEFtPmXF8s2me+qdIukaAUpuVkoIOEuwTbqnuLnD8ps
dL9rQomF5fN0Wykl9V0xYf10LCkRiNsy8kr/yUElGbYXtKnabAIGCHC+k2vCeuSM
18KK3MNCKyESFNyXIX1MWEb9vxuJJV7pWSmgGJLoEn76yWPMSxRPhll5+n4UAlyu
ZDw8rocYsCZQ3zLzTxf96sJw1e91Ouveft5fbVd4jmj/QjaJsvyEB8nF2YsV9oHG
69AF9tB8aGTevlSVPYLQNa4dHbDuH1k4nu1T50XOLPArFMRUPVPOA8/Uhk8O9OUB
VhM9YpbqQEO5V5AhAQuOnviHm3bbQfxwB2ULi3/CVA+WX9M8d7Nj4C1b9u3QhQ5O
tUscnxfMLs+a63b2tCE4KKyXMMcNlYJFWBI4r+1yr2hPo2K4LPEfKcKM0iO/bnn9
uw+j3YQ/K8DYNJ8ht7WgbMeOm+ZMnbFHvfN70PKJ4FTWPsB4WQeZIpt03UcycXvg
AI7/VJhiHtJKxO/5J4xvQhb0iQenUAdRKlNIp3+P27yztSk9uh041MMfP4eRcfrd
bo57j92Cs+qeyZJB8DqJkxWhOn54PGKPFQJ/M4k3smpoe/HtELSCrUro4po7ovhR
hiEopBTsfJ7szmw+CZmqsSYQeWxpJhVojbkOu7NHAF7gMyIzgzCtfmSrDn326cT9
eb8vEekOr5d4I/bBa9I19GQvCPMdv7VkbbxlG8scxtVf2jIIW64r3cW0kA8liQeO
ubiY9DbrPJAGsRzi6j3+Tkq6cDwJvthNPA15dzUgtQGmiKQPnI1fZUXn5DH14NHd
9BsPb5arenGSda/AM7jO0FfMjZ/l8MBrotDkfAvxqmGeokuekGHosWtDWqH7NUL8
gPKKQ3r0STU7pEkbfXMEL7DDeywCFc4dPICCeqhssKfU76b/GI7+ffYGtIP94/0Z
iJdNb+trp7U2kMR00lbt84RMZQbgHg2CyxR8vefTcvYlTjlrVuvbSzw8rTQzCHLX
7TFozOGLgUdLDFWknqlt6Q==
`protect END_PROTECTED
