`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LcZJO1IeTrKJjek+YZPOUjmuOPYNSjXvFxaP53fPwIo0BC0IOeSx87wSt8FkSZWw
jnhdJw5mDOlZU+G1uMh8cuTqpnoDYTNWp5bZ1xomZWf5aUv3njQSnvVjDqHLW33Y
QmTaeQbcNYNvLrSBc7kIz03MIKUvxFX7v3PeHulnvNH7opyAdv2KtVI6P6i0Gvym
F8LYoQz4Hd7ze//FsVcCWZkhArchMPptJSgtfddAuCCsHTybgErZ/Id4lWAHPCnL
h/rhEuVYTYteRuDkELGzedyM07foBqYE7K52ogSTSxIKhluSH5w+54Enji4dKXGa
uj8NxvtAcidPxs9pjJkkkeQjQ0nQ59he2nqZAD2JaMqHx3y+pMRYoRdgWqXUFm15
kh3IjWh6YEvnvuEVUHSSYOCK6cuU9EDBJMAtS2tLoK0V4mM7d4DliP79U6m53JB9
Zg9Zalk4sRH79Qte1NROkk/AfRP0xDb7neTaq1AAZf6DvIZrX9SL5hFYn/Qvqdnj
lYwk+dKQC4HxST8ggSDeINFfkiWGvilBJV356skW2Q1PxvNLxiBHQo/EaGiu6owg
6xYTlf0MzFr5Y1ym7dpfDCWO0LSSdglOykFVYNdWB4uC7O0rTh+mC9UZFfFdx3Ha
rwd8yzjT9Gstz0R6QLJUPxquANFtjE9JLuBbtxE1lAY0jN1WTQiD5j/zIWxzmCZV
tnbbnCR4vW5bJNBNcOuzOTPWpl0E2aCM5F8byzt/Gia83PTGsAsDv8KKmvQN7NnS
+iL1ZnVrmnmRaFR5wKkVj6SY7kJuN5aO59+LcQtyzMBrHkEpsW5GRT8lHzgjMo1a
xlliciSjmZ8yeFiW9+XG3+isEYueRBbEckTRxbcgPyKNZ5mh72pnR7VgBlnVczva
Gb1/xy43/k0prqPocQ5KEMuDhCgt2nputDAvpOqspjp9HzDEFOnvgDuu09BZ6sy8
yEQfvo8a6TzYxY7g+IMxk4M9N1VBQmRohTpL8KiP5ymreIxAh6uH5Xm/rZL+2puu
fXriSZsNZ+V6GBD9Eagy/B4LcTAsOqijgAFj/SU1iuLE7nNCiK9FcUQq6xB6ayi1
Koo0Y0JphswV6yc2/SK+d6qXmns+KqZ6jgb5JmzOKARrNm743YJHSp61YaxVrRWu
Z8GBHMSptplS2xOXNd9oM09FSsV3SDVKIQ2r7/x1XuJjghKO56nuW/7t6s0yuhoo
OArHG/gKo9D2T+t1hpFr8UYWtJPM34sjxRPQ5vXE2fvYggkbDiqEQ1nvngwWwwR/
Err4H9XGg5lEOR8jI0xEMrjRbjOB74Ms9RMleJPZbrwiumUJmSTJyDdMHU4/4nOZ
c4RvLGK8yUwD0oHdsO8z0kfiaLFI+Qki6BO26xKalSjFQo5SNWzaKm7gl7XxajeR
eShw6/WTQYdgsZqHa9w6VapLNYZgzjef/wng3LLQgBmNiq3LsYcNaKMVLpN6jfO9
xLVvMk3jAmLlvQFndiEuexhMG6eLX2zIPbj5o8XYBGB4UF+N7qEWHg/IsxZWWNUd
pZ2o1iIV92Wh77iHK6G2/2Yk+gdE/UOT6OlIXEBAo9qBDD0yn+dd8L2/Pmj3GoeW
LHsgndwAjPjWdEucJCvM/UG2Uo+g1IgC1HYLVS6xJ1PgHdfP3X0tfpWeQMy3hPjG
5wxgx4D5bAh4NapHTSzy5zcd31aI04P3gb8PO1/8gjQqydpajCSseEb9SwEqTeCI
2AJD0Bruve7/bVTlFG4SR4JjpwDT9f+NWO0U4pvawSp91azo8RgAq2d2qTY8mINk
ACQ50R/ge7bxL7HiMmXrWjPOZus/3W+EsFbKpEdDo1gkllt0DRXtb1rms/UtJ8qa
KQJVzl8apC1C/36FuOKxyW3T9NltRCdiTaABJr2f0St7WnzGjdgweYO8n6N5iG+E
3UsCVjkX3oMm2XC2v7C9HMFXWP9xZX91u0OUcyHadpXccz0xUR+YG0YH8CWly1xh
hJZjBnOkxDUouGwqQG+klrCyg79q1SiKIoyzg5WbwrFzxHtRyur8c289odn1No6A
I20n9DdvFUcZNIc+h2I2SORUG1A3boZ28+7VbYceOM1dcyM+3dvD8qDaCRdgHiQP
eyAjvV81yKFroGck4CtEF9TOHM7C5aNk9aK+nwGRCU4szXDm6X/cyKVRocFmcPL2
I2OLSfedEbPzFZhTxAXJKYo9Ix6u1nu4EEiXbk2yEE37azeabjYRwI5jCqcb3INI
hG4Q9zG7YVWRLyx7YH+BBoVkhRGclTGwLRXxS3uJl7cF7YgYg46q/Djq68qCNsvO
M3cpzKR5/sZgow6fgTfWKh8AuIkq7RYsQZcg9uD6j2gHJHeIHXDYEABPRgSXCmg6
MGGiuYbAzD9YpaIq1qd76dXWYK6oNTBuXNvAdjIjch8=
`protect END_PROTECTED
