`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RDlX5IlNI3kxcwT/GAP25JkffnuXwdpznLYUk8Re3rTfpf+2JUA/D0RMvDzjEGEr
tsAAJYiH0Me1XqmJEYdCrlbDSoBwsUheyflt0rDxGAmVAW4zE3b93wGcke0BqqLa
CSThw0OyXuRoCVoG6FFxds/65yJmSAtthtImb0hrblFje17CMPSAWW+oSrgY76vb
ETAymHv3WFjIfOyYv0ftThdUcdyhwXS72ZKeSFFA1Qtu0JOF/+4KAVtbc2Hus0zq
zif/EJ5Kd9kJHcoSVqOFK6Y8mfdA5/6SQy312OhFEiFKkOv+IWbbljKJnnbXX37I
GNReNRMw54XOqn9jH0aPkjXIJBcgZasP9HoI9UhPybHzNXNHglfjcZCmr7/DTzwN
d6Io8udgWE/jl3doChUlyrbrppOg3RdMz9NEmp8jPBjJV0uK7jezgsZCt4RiYEP3
yE2MC30B7T71ap5gnQJUW94jUySUlxpNTBt13XbSR1pXu7N8jDuXgcXKgU/QtDjG
LcVdfCA7ABwzJ2DI/2Y9SRS8U9flbAwNBXkKpbhhwBLQvuqa3E/TlE50PaH21odV
6Sgc/nd0FArbA4Yx6wTPGW6h1WoZLwwxPoWAxsf9U0fsnuE9nBL9HTU6CLElauz7
RkYnlccviyIUrTa2UmjrrZJXW/02GwZvF2y20xL/Cmvlif2J3zpdxrwadCAjQ36L
bcQvUJI/ujl/hz/pE/snmSuIaLibvBdFtoh9qG1LsDR968cO2N5zawEUfw9xBFzZ
O1YCMjlVCOvau4VK3EVG2Ko9UYMa0UzF5Dg0yRPmQmvlu65cMFux7Du1DKcmzo6a
bTj+tgAQNsUKQiAo0zu0IdRzdee5/N1qFTEuw87IPKbtM6mbPXhQf0jmmOj9fIXM
cR8OKLgKgtof6Dk87zIEzcKtbv51PA5+FTtsXnO9DfFWXT2n23hm+OGEYh2cZrSJ
B60RS2SGS3tNtytCMCfsIFdQBvdoLoc65sovf7YV+96Pr3of2kXketjjzE/V9wDD
mJpq/b8UiQwKPDO4S5oZ5m1r7Rlbl6yf+XlrZdE0zsnP/BSTspckPdw5heEXfARN
N8VrpkuRMKBFUTM166OlbpooYKtC2FaS3TgDz5lP8OBrGHYKM7uxqLyGJeColNpu
97Fdu7/IWFYaa6MHY7thgKqcP/s5ymoQ00j2wiDfrDBhbj2Ejw4mkOKcIBuWZV8M
DvX22RpKiJHrYclwi6f2Ndc/duAEGaZ/nU0cpig87T3TWWhfbt8kYl5j1TbrKf2S
cYPyxWU+1pDhjkgL/Qu824by8I60myEUWrtIVhDul47MQ2TxLmqE8PLPKwx8eirW
k8idqN/VmwwTblUijPx/uLZLoYGjDbZALyP9jCbmadsAcubFCgYeyXFw+zynckOe
+l70R/uJeNF/UuTYIvSvalZg48qjJyW4f58LGPaNB1HSLJnouA4Ur1zyZIXU43G4
z/Gpieh48N8bwvbpVzVMKdM0kq7ZcdCba3LZYpWOk8KmhwNya9R8NQpKutHKeO/z
/Cb2Dgxb5H958YKwx04cku5YpZCjB7zP37LqOoN+AW8g0fS9Pcghq/+Wnx7bMYV/
gdKWSXBO14w8Fl3oy1dHT3FfJXFNCcL3Xm3yzfA8P+R+FgmL/jqRj6/adbqlFSzp
w+Q/86yFHHELUzmX8ZqHG2AeA4MEClTSH2URND2KFbc=
`protect END_PROTECTED
