`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vEQC8cDF9C+f5iTRmutNAWseZ6VzW74UB6fs9Sp4uiuvMveET9wGB9wG23jrqepn
3KL8ufJZjg8o7qY92UNkz4NKG/noo7VwGpF4a4RA1zFYZjUe1fqyUuw/UGR2KOIR
xT3oOlvWlXb5hMJNn+P1u31YId9xfwrRYiVZOyX6OxWo0zmMwBu8oRhHwApPYlz1
1ncjqBWS/7KmlWMACE16ZfeMZoQJLw80ysALWQadBmxGA1ehwRgKMqJew8qnQJsA
8B/9M7gREZVNUvnS3P5Zh2SqbC4KdhtKCm/6HfZmB9TGvD1raZUt07FdVX26HdTg
AtC8fixVKHMUqz5fEosxGlKQiagEUZZiAKisbOQFHz0oejptsk9QJQanJ3Plpth4
tCZnq4IMBt533oyFi6A8KKn5Au1Pl2bRTPjX1N8ZE/ZO91Q/vFBfOFHozrxVmghe
BLXCH7okNi+CprPAT3s9WWSjhYSWEqxHp9+NdO7DkuBarLu4PLMBwwrrNXN+z2oT
sGsaXZClb/qWYjGtGA4IrC5FE17jq+laOlv576frB4qkDC7ExAlR9i06qqVa9MD2
JbJ0lrVOEtFFcEE2upm8IL9UXWPppEPm3S4FcUFKZ8c=
`protect END_PROTECTED
