`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xllwwYgFqcqc6WDP9530d+tsnOXwDEphBiIxd+W/iEFIhJpT19ZILuS+jIWFFlRP
y533obQrqdN2R+NAjXsYitfnTuT05/zosMAJYuNHiItUGCRP0rnJkQbou31lnRpT
c/vyi4ypES+00JsqrseGTua5kvZB22FkVtuSM2kRLQ/jVucdTZSk653bun8BsZRf
5K8FmmI+DQsS4K4KFXRsxuqTBFGJ2Hti60lb+FKgy1TEysWZ6I/vaJ6p7IuJN2RP
JAVb4mvELWy5oiPTA6Aw6StHG2V4vOeAcOYf/rJ8O5lcP1HAUynRJtRjDpON9bwD
Lc+smRZqBaNQ/CkwBxQ5ohmlY4SpeeRxIfgH8WXkOBCzoC/FgZY5WlcN2O9VqEs6
s9xKGkFzHqhPK1e8vcK/nA==
`protect END_PROTECTED
