`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6IXrtI/+dY6SyOiXA7Fd+eEzD4Wdnvx266WZnlc6Sr92VkyuXEwbDWwcI2KjBohB
mhlgdVbLTMhe8AT/wYW4J7CSgHHUXN67OGelPExV4Izik/nvm0yX/jigCY7xZTyn
vmZtrsnkVcgQWUeXdRgPeSryLWFLtzxLj+Z18WJ+XyXlar+N2fp0o6AsxQuw0SHs
J4G+0X+hg9GW1DkqR0ndFNnyL2RHylaE5J7cxpvW5TkUfs+E2eLcAZxlEa+w/WDJ
gZpMWq+ruhsd9x5aKk1OS74csxRrCOnOIxGpgbCNQI0bvBELzo2CFc7Grk413MXC
jGXqhRleC5GZivwErD398kkli1LVcrje/8dWnehtmsNx9er5ag05YUIM0/ckU4+E
pkFP0TjYJGCiqKfYk1ajXaiIUlmuqz7aEHyn2/vl4swoUU4LQHi4Y7DqNsXWJkXv
rVhLy5PI7HMJ9FyBqnFKtn9XoGi9GuCzUhOkRVXiJ2N05rDjkrqN3ok/KrnITIxG
6tFqWgVlYij7RKJk2pfLL8LHgST4zH3JrOYLVBmAkfb1B3ZMyR7tnsEHrOHMp5c4
EXs+4o+enQBCCj8xnnZh3Y4sgFtlv/BSCOtBFrRIIMn58vaN8vz3LEN6UZHwE1wF
MvcNYoIgkyUAliTxr7yldLgAeK0w1LqFH4si0ExO2/soPs0+qqhHzBAbzqp+5+ov
BaEKJlYhLcmOZG3TuLFNuEc+b2AKbRybshxkmFhLqz3bXQhEx0AEzapSmjezlqsJ
P7V0AcZw1rIysjiRQ2IuP+k+43hR41Hh8ZEvwaP/9tKvxle1VcHCiApjaNLvqmPN
2e3NqZrLY+qa5yBWS4inXb9qSrKS3MsJTwcMWZN5Ypleh//C+3JubEAs3PwSsJ4U
yF4sOvveCD+1wkGXW/XXszVKRVrMR6MG4GYjydrdfktEkCinz4zhYFMqzCS1a0tH
K0OTtLDPWk/Pj0e899n6JBtoV5IrEu6XHTA3s699AkDJsWkKv8GNdKOLcXba3jNX
GVjr0akqkKW/nDAmwUziY8IgYtyGJokbOQwpqQZ6zenCDcMlbIZWJJSsfHOYlWCM
G0tfxYGIkK5HQZCuR21nrsCV+zp8X4MnrkofLzIfNAQhjasm/jA3pgE720hTIvh3
LFjmunYnZ+JVl9mO4pgEN2nOlSQP+TQTCnU4d+Zb1fokKV0VN5o9NOpvxmLdC20z
z5+NYGdNcKsNmUv2B9RMMi1pxASQM//XbI2M2VJCpw3DL0kASugCtkuBZyISzXF9
`protect END_PROTECTED
