`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UpBlb0q/EosVmSRhQ4Yb1WwsANsWYTvvYbUGrTGfH0xot30QOLlvOYRZYueCq+T5
RBJyrz5rDH+zhrspWjTmbcgS0tF7ESKoLK63to5bP+f/k1tyAKZXdxu/avrfYsIZ
lPJByy8e0qeqRECeW9VNBVHYlO3TDZhEtTV8P+Cdy1BLfIMa4WCy0E3swedI4W6E
+8SfK8dwhy4DLXNJPo5wBd7YcjWvovmqiaeunoWpClhNsLzeffMV/EuNRuAPjxCy
MvPXFUoauFJSC5ICffN0Oryb4phbSsvOZ8ubvsJ31F2gK10/B4vJSgp8vg2sdBDD
B27pdfJzom7zoJQhFSB93JfEP7bVrD8ZuYSXRdMvSaK9uJMg+bhO8l0q/9AXGRRp
vzwd1z8zgfZOOpRDpJrKuRCmTWFCdlJwgCUvQ8OqZ0RuW/Gyl2j6n8KR7zjYUz05
o8cIYiLgI5QCL3Yyx2w1AsQwqD/PXR8Hs+rtZ/LMi7WVTYzIsO4BfgJ34zvw1Ndt
FKffrHDKtx+kUfEH6ASfWd1Aurem4knXxdKMb8sLaDo2gRhsvCW47OZD/Ka/pZ18
BXwP0ccrTOMTLEhWVvvQ4ptkEpamVuw2Na05l+PHU9JXQwNnfoxSqx45wLGmn278
y0fnhSHUVe10XSBqSElgnpNtuOO2VcCUef38QQE7x+kz2TDXposvPMijuupXtFEI
A6x3fNo9OeBdUJ8pskYLJ22v6Sywc2jxybsX8czX+5pOgrw/PFksJ6o+E1ftG9jn
HXD+Wz95vALgaBKQYq6WDz1oHy/A/WHJBdf79aMQGqpRJOR5BpD79aXZpLpjMdHg
ugtoD+mwSe+jJQqa7t4opUTm0/LLdy9xDPRc1gtIMJv11aC3+D/XkEOBzf9q7vwz
MQBorevVH/a6BI0GmFuNpfh7qQK4iN/hjCF/DrKu/v+604xAFZ7QDISPyEiPkjDZ
3BG0p+DlBW1FVgyP1xxovyk4mLzRDksYmexledh7qobtbskhEQTuoNMAYRUl2cW5
oj/JEmWauORfoSlkiI1ug4hX691UOdEJgTsci9RUWQB/fwO0SED8w2kL2lXHCAte
0kj9PShEn6d+MLVU3XgYybaBYgX1YHIu0E1IAHuLO40GGrKr5lGFNMLPtBTtYPdm
J/Mi+391AkqipfzEpjl+8BdeZw7XRbQEFPsKo2hPPTH2VIT+0SiUdowKvggrKY7D
sIIRU/i4NSjEXTL+UOhOOolIwogJs/HTXt9ikzFrWyqSsHtVQ0ceDIwz+ILSzn7i
Qj9Opi+VYfGz5Oxo3u69NVKNYaDXN8tTG+mbuijqucf6Z3P8LNk4EWL1NzyF9Vbw
ya5P1Z5LCPaMelhnl36EdIh4NG5I6bKEUEr6v0vQC3o02yQQVKOa6/alZhp6nnaH
aMZRGBQAmLSfQmGfDTSntzs2nBxtLuB/BboKSnTy9XSwGrIh1mqFLBn3vKYhiwkH
KFHe+hY5XqpU8S8bHjJFepC+UZP7IJrcne7jcxd58WI4zv60Pn5zreFYoV0azxKm
Ltl4pnS5Oso7zE54ePK7bSsAaH53hZyUf+cVEbShz+kT98I7aZ9q2zm0LtvQtHDx
nf7A/5kFT0+sBv8JUypiMnN6ISLuKRfonLnyNZ11hA6oDG1Kq49rH6MEOpIqwosy
Yn32lfULjWvhsA75s7H5KUYJnowvxfZlkq2c5wOrRJtmb9F524jIoCP2uoqdtnZ/
oo12iwDfF+zwnwPUOuUCn3oeEJXJ+B2BmmesVnGFlYBPhyNsGWRQIu9sQt9WVvtb
P6dEYU+fQ1hvtmocqN7w1dgE2AQXAUemdqgvNTkUT1FTrFH+MQQ4Ecd/LDbdo5UV
x7qM0r4GtdnH7aOqqv38DHvHXFtM9gRx1FVWAjF5snfu1mxRf+pie4G77SL79uD2
ObIL/x2ezg7rY+6LG4C6iC0PAQOpOMC4FufXhV0zErX/VhiHuS3kvAUD48Bfuxf+
kQeMRE6c/nEvgqywBaAZ1vJAx22FYJkQceMSh3ZewzVoBjwYepamB/1g3w3I/VT0
WPkNcRJ3zE4ROfQqDYkS5EqWhdkLzyXmzJZqt1wqTnfZApCofh5vJFDfQ4f+3cgI
Rx1NthwouBghPPP9pqKRJ8xyNph5muscfdZZycPjIrIyQ94K59xtk12pQsTP4phT
SWqgyNzj4a2TKaWa0IZbRvMBgCauTusFK6iZq5fiy8OGj/4jCeaGCaQ77WZ9RItW
9gf/tTb3n1bmzbizvlmyLjxwtVeTecK5fAFx9ngS0wQVO3SjecYpB1VWZjjaPYZc
MVdHFvvl+9w0eHtWfolscZ99k6wWKrQdk7MGicOchb+N8gWsWjjxrKOh4+vHSZ9V
k5AekuzDkBg6Ud+lRyVoBkNkSrf4D6VrPCHeFSKbohnzQl3Wl1SwRNT5h8hOLrwZ
5KLuoKVeTbfkBy6j22V6BaxpeyFzQjiXZhtg9M/7EAqdWKOWk+JPf4UwXwdcWXxE
adLN22KoIjFhWa708+S1vR4VsBtwtfc/QZ4pHisDWsZc63bOn8RdT1IrQJjs5REY
3zmymISzDsTd/7+MgFQ7RAgIM+XzfJIPXiODF21pFC90cHmqeU/l99uSLLyX84ow
7z3shbsXz8s9YdP6S8WtLaBzwVcCF3YktjoTXD7558PI1m6HXNbXcKQ2upK9HkC+
icjVSpGtJ5UKIltORKbc0sT58xyZq31Jdip/BJxcpeF9qIsmM2jL46c23adjluxI
qUn9ZoIqFqWGAR4cCx1JaoKiZpzW5bBBDAB9qIZ+tj2sBajWJbA8uBjww0W9rJR4
bItki5bJxjJRXt2WphlqsFKb0o7EZkniLWauJPMeRihQkgsyyIoHWRrel+o8/klE
NJPM7vrHGUl1ZbU6B0ux1mrJVsQyM34zy2S65zzX+SyVuq+Tq6TAzfsis+chTifC
MHr6A8P0dWH9GmugK9wT6t1BddeBFqKKKnsA71RbjmDYXci3DmdyVgXGRoh/Syut
iCzjHWpHBR1X9vR12V7b1YFAz+FQGkkHtdk9O386lep1ngB535re7UM91IiX8qCY
2dF7ltVSCJ/rvLVYkKzl6yZTJ/PvEW4B9wc06WbomcIC0+n9KC5Ti+XRy1jGcFbJ
6xwBlWFvV9NtHf6Z5fqn3EdsXD5qZxS4RXKzSDDW92faTK5sOiKysUbo+9sOiGCq
6hLPo7gtu6Y6pB+3lgyel5p+h2xq/4FcUjNAoOiFZ5BJX4ZszaEyPdQoMPASLCtu
ZxG0jTpmhyzFRBVp7ww0W36xRlxK+7H44F6Mie0rcVVFIR7ydfn+z4UMKqDoQZwF
RAoSjK7zR00XxQnLA5eu7/5Y4WRy0ABO2QGv+8wzqjwbR7Kt2+LR+TSjv9Wk1cfY
Y4LjlCU1Dt4ajG8vU8kJyxq6RidTYV87E1681XpSYycTvJkPb7om1/FaMoa9u5YS
oXzxHTfSRwqWtQcLqc/urhv5XO7aCAQ5n7zcUFZBZEs7pI8RVQQueHNmtqdAKbzX
wdOVvL8JhnJLwj6FrnSg9vRU7jhe/ZCmxoRLf4LnRkA9KCWtw/fBFfrknNQZBu6F
WbuyrdVW8HcoZoqt81IhlPT5eCTxUChK0R2q1Ai6Sg+6wBLw3j78BnsstkkngnIi
dgAgYpYGPlTH378TubY+CfaZaHwaxtyISkEsg7EEQHM2p/c9P1A9RcmiFZTgkIF5
SLfYoR5at/ZKMq5Pgl0M4NRnogyWh4beb8lA9j7bE1Vxx6JhRT+sIlVA9H4tARau
9D/t/lu2ncYCmfEWO9SS9a9fMRIRx9+kIqmEWpIt0TEl3kFJMgecXXM0ApenaYuf
sFWs4jDgKjOYNd1mHVmiCcr7GQLOn2k4+dUblqBE/InhW144QP85+jV9hdgpogxK
QhRWdCtUdG/NCIRdGvYL+v+e9/EfoeMZasEym+fX/9ZHc2dBMReP4kA4/axeUj+U
pKdHyUOGi6vHSAZRpem0NaDxPqsHJKQJkr5pCm6sY2Dn1ISevJxWOb/sDKlghyI1
6LB63Y3wloF6mB0JvbseBqDC2syYEmYHnEq3ZUa6gmBQ90LoeJXkSHssEDrgJAzj
g5HcistrPNkAIZD2q75mCztBRjkUXjLrUmubPGkx9xlI2EJ2vd0VTcJt13qNWHK+
VRvXOGaik0hP+fiXqBwJd6w/cAHUKQJ3Jly8W/k7AqN0cw8z3wa7FEjYDNe6oDcP
9TieVH6EEI10QTqjJhi3MxxhoINAUsUnEyipGmoXz2XvzwFbarN7wj+m5GtUbiHN
oo6TPFJjQdrIvCXWqNtrgnbx6fD90Pn1HvqC1t5Ywi1334hCitFyic6LuM438DKP
WM3Oyn7UaxTvYD/Ivk7Dl+0Ra4/fo0LHl0aGvHvqGaR4VZuMGE12cKnB3qrSPnYo
RugJEuJJeSUomNq9s/sc1PDhQ8E5mlg/nSpyojQNOBYpFRZGQPHoSSqgcMHvMWes
ZUcvb6ZFwZ09ZzmuN/tiesGbx6m5FubQIk5FZWMWKi3uDY22bamEQBhk1zcR21pv
sgqRBKPabROm957QBenRU596HMqY96DMOQeDa1qWHay3Vj2IPKgjt16oBHL+/VOr
gRPQJxJetX7Uzws1pejlTlzdvlAJ8nGirg1ji6o/kh/gmqyaQ+mXsClP0tdb1BgN
E6ninhfrZtP4HorM3zPG335BFU8lCVy9uJjS9zBl+V/CdvgUOJzho0G1AnOYh4mV
dxJwjqiU3IpqFkkoHpEPAJaOIImrtPMQrOes7IzHLXwFSWdVmjw4LzJuMXf4Mn9c
mU7N3At/NCtKu8VHi2FdF9NLjWf57GLQbxTKldnD/+lLBVW0Z1stK5o0TFQXXebp
uiOjulf9fMZUX9yEV3fba+7MDEJQ20H7hzERLMLZ7pZC08e57xEYoMRxNiqZTE+r
AgvkX3kWPyk8lEAPm64lvRaU/EAJ5J+5gZwwmhHMBw5uDlF89++QpYwfQGJIklaq
eyjKhhugVkSl5B/8Vc7G8fxpQa89PXZbDnQmd3J8lwMOfNZ7nYU1gnFIjf+aTEBI
TN58cezRlJzGv4Ls1SR9itsx5DGu+Q/gbMVGIkh18ROlJ/RxQaQreU8hZHXz5H3I
dOLZlTW2M0ONw9sQDZEzc0MDlp09Gw81307sCQle52I9GWCIHAkIIc7oemuxthir
4gex7Q9Gg9e87QOvqGlPXcbzf5wFRZxTl1JSqg8CmTjs5ILFCiUjPPoy36J43thl
YHnZJLdPM+4sdYhgbgzz5WzTNMolSn+3mkmSFwDo15kJuKspuDE/hgkrC/0agev5
pf8zMxw9seJ01Fb01Ct0/VtPwEWAEC9ufnBsf4k3TiwIFSlsZlNjwNjd28n2VfHR
v7zrQHJUao0cHoNPHy94OZF7PssBMgrrVb0oXtqQUYbomRxEXfvVjHb1iM+p26XF
tHCHIuvn4wNkWU+DpH8WwrIvFua0vifJghGFHH/YXqaI9ERGo/JFly5ls+ioXia6
Rfd9cm62fdmrb21TmYAIwNS+uYIAAA/PYdSpnLfK8ktoJtI14X6x5eg5MF8kLz/w
IHxtxuY2aHSrsCgxfN4KI/PBSEzQx8b6UCHjY99/FgI+MjR9QvL4J1OQ3Ive1gd0
tLhlw1SvGa9fmH6aOlncte8KyrkK6P5lT7sxa7C2EKGV/guwrSAMjoJJVVs3SBub
JEIUU8rElUhIQlneefzd+5vgvO62zznVLczZEvKGqNjrCGimwvNamf9hK+c9jNZr
LQ+ILrJcJ8HvpnIfhGTciqLTvLs1MMTrnDPhm9Ct/80AWIb+cLywc1PyI0rkKFT8
3ui4w8+yzRklp+0CiBXMHC6ydl2+2gRQmY6zenXg4EzkTB7V53yRz720NQRiL+F3
EcFRlxARNUdurHbySYHCqmIE+fR6GX6g1D1RYJWS8q1UYTGJjZMlSHOldH3ljbFi
nMU66Z/uey8rrvocSZovf1BvZBofuyZ43n34dApz+m5euJY48G4Fp79IVQc+C6yO
AQZsC4sqEcRkItFfmbO4XFCUGvv13/Gzt4TVynGHvLy0b4t8YMw3rTFADeUMgZdf
gl8PAZ1GGuxYG2pN6z09uJN4rcm5AF2R9HgnmYJUJyFsr+0ZUG7q/xfkNdqC/2mO
ReM59A5Iux09b48SN3zgQ0DjjcfMns1FJn+stFQavzQMrqe7DfBz7ZE2rgjiihPK
Rjx5m1MTXF7e9u6zAyuEZ8rVZ3PRnlJilaK1Ulxc50rZYG21uhYM/lQrNxb9elm2
4tz9uvJnnXz1uoE0PkGevFpuO6/xymXkz32Lq+Uqyma30Q4zeKi8I8pUXipmjBLD
`protect END_PROTECTED
