`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OmRBuQhmE3Z/XGJ6qpWOyQyU1Jn86VgeLeuM5XfdqZjd4owdjLmV9uar8lcDCEnu
7whDIPGsPyzUrGQ8qiqvfR/BJT+L48qo5vtpMu+KA/7IdGvwYn41bgMyLhbX42CA
otL5EtF81+rM5EwssVZmmD6/nqkHBfMwsKBXgOPTiwkSgO3S+IZSdxRZt2SPdIWW
vwlvv87qmM0jltTcGZSsbs+R7qotTToGyPhJkcCkKpAumj8iRh/Sp+oIqjQQvMjS
rtu4uMC5kc9K0+bAOY4LIfEFZ9TPGilKNL7iWe9m8J86QEuvKg/j5wUnMAJjuoax
rkMBBeJgzSIKJqTZeTW6Ltd3TIX5p2+j7uhSKAewbjH26bDhKmJCsGi8LXkdTMJx
dCSrTSYG0gFms34a1d7ocrF29LaSn3TBiB4Tagth3UVB82JZzNlJ0CW7EEevTKYk
jv8bmIlxQ5nFAb38JcB0iCxORfMntf17hxw1jm3L51VWNGjVS21bXqzzaBVeE+Vi
mr125yexUOSmuk+ubSTa3agi3ygROsGkUJhmElFnVgwx3XBiiEb6Fa/kwOoGTn/r
6xjNK7kgB2hHzYEzoesyngjeHu14esjR0WvaVrfP1u1oMPnH6t3EX0XyoVTVQlga
TA/gVlYp5oBFLdm0KbZOVN0xoB+HaJSxgL4Tu6msn2GKU+qCdnHdo9HtRXhIhsoa
0oCPJUpZSYIZhFEQaxTi1ITzuT97T5SCpjNk1EznpuVJuJ5AlCyOTrBK472LjVJo
T8s4EAPJJe2MtWgS5edNR/srvTAg48EnsaLwzxfizdamGzo06H76lovnqiON7sqj
ONTBzhn3jxrSLCfdbqMtqlMn/r1xV2l4n7boeotDVcva4u+wEWtbdSkXJI5hj6/U
f0tNTLeiY1mD0I7lvl9QnDSLFwRaun5gBZK7raEno41TmIkyR+ntwlHkYC6aWPmw
PVXoyyCBiOeCNeeWOCFuYmp+AHtx2QR/NCDP6U53TVxRL8F9VBIS4u4BCpiU8tRF
bnhQ7mr8SvCDq3imgDmxAVkxFrC+vlPcnEAjy+wGu7Fc/5bLKDvUoVKf3vboXIrp
8gbLshTuyZFXn6gTKHXFsQkj7A4kdk8uQMrjb6XhUKfy6TrRFaD9F75w2RKx3lpj
5DA4aIvAajVivqNTO8BoXdVrUMi3d1HZ9MKwqL4E5vOTh4lmDwdHzMeu9AJnJwgI
Ouohjk9/51q9eMOWX+10N+XAZ/yXjCsnAMGhtjD8VNjyTKP8xcceIxSQLl2dFvTR
eYZC9197mgqN8V3ctn2woCqkKFM5y5YqBSU2vcH8nZLgScPtwSct3uTuIhkqYucJ
HrWmPCfnUiSYvmTp1ulYtT6nn9T/bB4U4R1uY5A4fyJIABvKkXwqFFqmFEbLxfnh
2SQaXHzo4NN4PwO/EOfYot8wG+edpgem0DRj+1LsHyryVLZWlGvBD5Isu44km35O
rTXXcDuf4hX6Vajt4BZz3XKjovvoMQ9lPe7qyJ3tMJX63UO38ansvi7VhJGEX6Tg
Pk8TNxTs48Vs0U+ypTAk8PuTagkibGg5oVdqFCfPGigAC1HxLD3OsXM+g9UCRzr3
vNzRsBgNyQCTwk9huWzcJrLHYKbGwepx6BnnsjHi6B/lRFfoxbqRIxpelVQL0J3O
GzZwKhat0uUMFouiBZ2LhcVXduLeyM4HSjqKoj3k1b1y/oSe+h/Agh7jZaPjJaAZ
FtUoO8qUmifx1HMfepJbziJIe6CR1/kvu6WbgBrQZMOpS2OZGQr+19YUognXkOYp
xEgIsGtNZ6hLzhtMOcN9vnJYkpE+YfyL/i61SzZBv7WVGUpKvISRzvSoS8Wru97B
WHatGjLYH0cyHMoUmzI47p4/un6m1zrm33QcQJLS4vDRZN8CRTwu98gsa0Ry5KcK
aThfRTAQqOKK6KwIYJvwpJ+efvWmbgVivwmUSecKEyIMXM7fiKcew0ycxFe2Q4Pg
si+AK5shff6IKB+CIs+Ojewa0mFz6gCP1FSjlyhNV58rfakrUdCR/QPXNNVfEdHK
OF0vo66hkpoAL0c4g4xEQ/gOSjB1titUQfANKceOlLJcBSgESuRnVMftXChWEjBD
nakbedYjlzjMQoEV1kWpEtBXmrDXNgu2aObXNKOEX1lzqTE/f2p8dAjIx50AFjnL
BKKHrGdzK3QavCHysl9SQu0QDH1qvjslGhmtjhsSVkXn6AA5R5HjiT04g9QiZQ59
hSbikCNHm7yIVune2G2+5IDbeT3uYAHOljQ3YSsdyqKwLgZ7X3mlnAc0FY71V4mt
n09pY3g+JHfEB+cLiTLfI4LlGKqxqvHkaq4wQBRrDGk58tdAD0v6zyPC3V/ficAj
3vynpROPQiXS5GJKDF+e6Ra1jLHIE0kUT61iQ/Y0xSn8UAqNLoSZJg3yDYf/t2rj
iYQ63MRIKUDYQ1hxy8TwQwspm7XXt8GjQ0tz9D83apGhDyOxDXYL7/GkHtkbyF+8
7Uc7FLvtoZ9nSjFgfuzya9MAVyp+/gDSIjiTbJUZWy8j15gPIEp2ULb0HbVZbIOM
9Y2dzZEgs+4D8cxNWweCz7quDlQKHzyTGCJumha6hVKGlxdN5dWyX6Hkj4NEf3CN
zI23VPtc/bKW039OTIllJ1/KChK4RfRuh3YOuY7CKt4UAmLcKBfqOs1pHwXLH6mj
qqiVND6kz55Jh6od7IpblGJTW1DiqPW/w2iVYNwmeRKOGnHPguHQbU/0moVWU9/0
H3Ekx+Gow3CbcxEEHXooxp2FzH8ihCp6VVZlSQFaM8LqfpXYTLRtsiJCpZVpcFA6
manZv+aiqflzc7mZnfN7uwf161uYjqHI5DeTUrbp4MGAjmreATca3qedcrWwuGXK
ptjNveBbzB+U76Sg2AXQkHtzbVXdAAkcTxE7URITcgUHr0mP29cAqqLcLDfWLov8
5TImec8lQEjxe4zfyWThS8Iewl4GnOu4rM+/72uUI2en/uzjg38Nqg9gO3iCkNTb
SsUmnhd5Zb/+zfys1xLzMVnVWW+LDBd/cOHR19urCNBd7JbWVv0i0cJB/UUN3bn3
q5Q//z80WiD9hNfGkGkOsI4STHpPjYb5fRhpKPvsHOMzTyVcCKLXvooe2IdICjvl
pYFm2bLh1W8j2f+bKt2MXipR6m0UBJg9xb84zbst+nMKRAMIO06X2YmeJFDPvNTV
1b8aq2zFmNSvsWopRfmu+rHpApxXUflQJDNUo71oXkvIM2L/kuTH/T6I1n8CG3F3
8ic193njwxQ8Czu73XVn6MEiAsY54LiBiYO1akdnL69ytCR6GFB0TZF8Wjz5+uek
LJZdVSPvs56tFB9nKss0ugDSF8SKv8/bTcR90hzh0BjYz1IoNFN7EGDDM7Fu/nEa
m6+rXqH8AUM2z956HYDE+tE89ekH8sChvZGo+mFIQB61ZvapZ+Punhgn0ENDsBUh
ZmTnZNjuxZPRYUc4eE6HcliKPH/Q4FiMdJdzSHGCicKPxgho7MPvhapUgYW1JjzG
XR3S9E2MvWR4pO4zDbSahf5nqRSNzzwWLsWOpMfkEPY4U6mv7PY/osQtWZ+XN0q/
C9U6sGP/BoEXtmRXaeZNZrLdnbUzz41NHxNXjozyF6otpzSv1xE6MX6tuzW0Iw1e
0QWRjOllnJFGzPKgC8iGYLDSa/OajsIijl5IC18PyNMHZNgVmEvQq+ulJaSBK+nj
iO+GSK7o4R8BtVytxhfT0uzygjyfV9MFPwVUAp9LcI8ksh/yHgQRL2lhkqmgaF6/
yF5cHQonkOmAV+un2XvsNwC5zRXs8g8TQsDixanWiNvQQEhUSM5jQc4VSpvw08mq
kpOuaqIKq48oWnHgGjOpw5syzkNDfPJsKalZum5bF3w9olsRH9QJbLcA9EdKe5kd
JRowfQ8H6dVKbzQJJuhuVALIsHkwklcbnZTzDNHqj2wi9UaeIHGOC+qtMIt5k2yX
lKENWAoyTulPMPnnfxQi1QhoSUqTdzEAeJR6ImYgPgHF2GirDrisf9qsi2LIm/WM
u8dUtM+Lj94yQ26x6lNX/azcgKthP7uh0N0+Ejxn8JB5fC88uFf/YaaFvvHft4a2
F1sftFwVTF56ittDpd/vbsPRCkqKzEfZDHcgSlraDvFzOmNZ3QuTAMSzsKExeRhU
lz9w3GdjKFpVI5YWfEcy45wgDc5pDP7huJf92khb7FcagQSBodVd7Fif1bxEthuM
M+slGCC1OjGB4n1PIRKVbS9DgidBsBoWPZQ2ZusCsbmcSyNECAbO554n8Vi40bdB
AMsJZSFMsJv7zXymhJpbBee0B1rkS5Ot3k82uPwbhObPsbWfDnoLvyypSToaGN/K
iRj/XPbHtGEzE1YkmIAVIH2LoOA8JyjTS8PfU6z27DLbjwMp94KvR3t63MM4MJge
IUnW4KD1QKjJ0DdTFNvYii4pA8X98qzA6bpozWIAasa6/f0nXdBnQgvOBMZSxK2Z
PGBDP0IZS3Pet39YxjXMztISjviMhejwUVvJEZepBAMsSCVqDcwkrbN1uvJhK8ED
YRjkFZigytWkxvyDwhnZxSj9QZnkd8VQmlRUI3MmOaAJZ38xEFhKTZ9LBaj9KGJJ
BqLU66cNVGPJIFUat2S6eg9XtQ/u1sGzHQSBP9dMTONrt/B10aBd3CJdRRbi+OVT
LoSwiWjcg/dxbuFbWfr3hGL1SNKlQC6nhBpANjOvPJDnBGurBJYhpYuomcP7Ssmt
ptKd9W05+gaNNMRe+Ssc96avrRzT17p3o+JKdFvI13ui1ic2YwjcAaMelMBjypqk
0K5U9DTtkXSLxLLSnLfOmwNMFPBEntaHGgZeElP3zyn5/X2iui3kU+ZFoSG3z0KD
84YOA1qP0fOa2a0pzRZKuKzllF4lrdlW3k0QXylW9RV4RcwH5jJAZ9a7Hv71/UCk
k1PAIzoEQTPzKJ+pQJgZ5BBTlHUYkSK2Fb72mpySIJxZlkwwdH4y8MjM1+c7iBtL
V1B1qA7SS+PlSwDyMNNAICDRGyN//CycLTFLkmJYJxa9S9WJc8GZFAx3fahJk2wy
Ggy9iYdLRkfH/bFgA40sY8MYgtPgmSKaMpH8TplukZOwOipqQu//lgbnWDY6o/FP
ic8A1Rgi3rdd2Y/0HUIMQAfJT7MIynMepLIvUkqv38ljYXfKRgDe5fL7YDwBm+n6
4K4Swk7GgXJ+CuqTkb4myXgwhSCRefqnV3LRwMwT3omx3wpNIIkBdy4KnwTXw3LA
rGZFDPPU9vlj9szMIXK5RHFE78duHRYnJdmD1NfLtcPN+fJomcpU49SerETN9rOZ
laZuz5YeKtHSrdav/+nWEFhrhyvT0300Jxs8zFOMVN0I++/eaRaTxAKna2QlPyck
75tbrKr3Y1bMGpLIZKtWBgde+IsIK7/Cjkx9v8XL5vh6lmiheLa+zzynzxvHEqqj
raIDy2ttf6CjBHIoGKhIeP+lCRBJZ1iT9I/wYPcVvl/OqYeVuaRUzzKg1SuAK0MW
ZZNfsI3b5FC27dVTMmeucVDFqNYGjI2wZ7Ejb5DEeQZ3xsH2Nq+2SOsRTkTe73z4
hpx+fA7L3ieXuJEJYhPEddWBERmVH7q77eMUidI74gQGCdlbSLQ+94q4ppW2A7iH
0WEB+crUiV7vhTQ1TqxEbI+aNNOKYYhIg7eI3aCflu5w4ll/o3f5LCceRon6kT90
iUmJnY4mWXWfkcvTmKPziNh5QAqT7Z7itk/ZJ+bS81Lal7uTPrc21Unx254seRB8
7MZrxenuh/B4c55qu1AsAunY6rbGa7Msw5gIK7lX1qCB3sxh3GMaGZ1QZloZOlBq
/jMDxmEI4NMWr8FihlOaC07SWRb1lgUSCyfT1YgwoTB24CTCK1m5qVKeFHgjTWv4
ZB/K6ksQZ2hxoIttYs5ZAmt6gmno3EPtKa94eYUriqfizbp+9p+D12AD1pWJqDQh
7ZbGk2/qrhgZuDu1HeJG2FaDx+UKD79w8PR7h/JglQDJ6TsrDrAQpzRS0VbOvLXx
inQF+CjxLlrMwpgtXLtH2Rk/tZ2iHzD2RNxBOiTVjQsznTkAp6tvjUPp1x8Knemq
4+GLBAk46w5XuHfOTc/sSoUEoasL4QYFN73vMGP1L705daFhw0w6NFq2kuupZxWY
JhJjnLeNsgHSRxWUgdqGSpLftacMsfdSbItzxVQSjGoGtiLFJRhXy4g+P8Zqwc4z
yCb+EZh+kI9kbCNSpsWiprF0ElpzNTvVHywJzGm2CmR45GkgykNss+I7Bwxutm1F
zrHnJjDxC/sSLhxwr655PVBSAw5c0ZszQPuzZjN6dHDsvf/1UthzLqu+e7MOUB0K
OGWambMw+VuUCIUl0e4K1GAxjKRGhLEMBQmxwSp4qpmTHPM383eJB7u6kxEFKDMh
lCcGS4+5dwXZC1pppecZRoUdCWRf3zvP2EfQSQsKxU5wfbRoe2BaN+j30yjlSjT2
zzgMNDkIRJL3xxPbvRy5dEjhReduHN9zwAShJWUAz1IpbQ15CiI0hcbRYm8gBe/5
CHGpOAS+840KadKy0WAM8G27Kga/MARrwBuo59FLUdtAeg2aEmWkH1wjTl2ZM6kf
rUY+v+a3qkgngrEcygnRCvjxd828UokY35tWzq9xlPCD057xuXu+SBDusC8QRAH7
FXRh6rShgq1ke1CO15iD1WxJK0QYncDvnTw/R1OLV3dxUmqqnjEgl7VpnutoLP8B
GnJVhrUhR1PWP6RyBD9NZjTX2L/3i6ADtFsK2UYp8yX0GsUtdkQAv3ecbDXJ7b4d
RAt8N6G3fffaPqANedelpcdrK3uEFLI7Kz+672gVtVsl/qTNQ8NtFut4x8GB+lmn
rHbJwK4MvmDE9Jb7oZe+DMPTNabT4DTVxusLuvE60mbpFnpzvSjg1rMNT/gHgI8r
KFiMU39DlLmlYTwa+0xbdnK/LCgBRxOeL1Oyid36m4P4gGvew2e/YDYP8bNP9ywa
HN/Vi/UnLCVe2h77Wm+MsuYKOmnuq0ZohuPqdNKShtIzwbimgsIuqKT6NgAUUBjJ
/zD/SohQKquslgm65rNmGaj3wZjJ4QZI0BiETKPvwSYF5Tf9+JMfOdTL8Gw3HF4t
V4UNSltGfto3tqrqXCpNLaxNoAOlwfLSZYRvDrswm8CFbRu68MaBz7i3B+kaVPUQ
OycYO+nu5uRNwyWVr6+b8Gm31dMOcML9zZlulME4GPT/wbN8bgcoYG7HAiLWKjfe
3f2xaQkXXOWkZ5uWdfPDAlp9xyE7FaZKKS0i+I5jCUgI8MaiuPyTD+Bc6gS2tKqc
SlWtZTT4j/b2HUeHU+rLB2vwNZDrtOZRelynOVovd9wq+fsFadsq5Bu0Ci9HnbnK
8jBMnHn2U+1dzNYPtwxSTeHAEBhCDeU/Rwyoc64FDV0wFeehf2kOYrpsBMy9YOm+
R3cNo+NYOkPfTBaTpTvKMWFfmXZqJDF5DyeYuqH1uyJXjU9a8ViZTTQ6zr2sqvTd
tNBJbsdRsSWExp5iD81msTmeEyvtIl3EIbnhl/sdV40g3UqmWjD2vpt/PkWsUAdE
PeaL04TFYAisSGjvzAOQNa5kWm1egVCYIMpVKq5N3/nFbacKxDbsb+uS41EqzGG3
xPL4yLydXjrEBAUij7EAh3or6X15qqvZuLnwAqIK8H8U4Oo6cFk7hPQnG0YPcJY+
BU+2hPrb3mh5Z8urCMjcuGMKNZpANmpkp4DKyXXp2OY+NfLcL+eR54wwWQKAYli9
ogNZKZn5f/9G6ZvrwYkIamx2GjxzRkKISo2EtjKe5tOJNhM+klkL6pSWpWP5uoo9
hTBvsfA7olFpgNJFLH90lUxHwT5LBgg9O0YzKwVCw0zWZUY4h6xgLRlEQzdPSeqG
00QCuq8Ydd9WN5aUHoH3FTcfgWHPi/fze2hR0Y6EkL4YJoW0XBrTLZqG0Dz+8PGD
6toyjseig8ZuvgYT231m3ae6Lxvn5IyD2QqPxHmhg65ZXIZZKxXKgE7sXHtMx7rx
FEma9YebrfZ8TrJOr7FkanqFHNsQyMs8Ms8GN7l90bMYQ1X5f6QQZV7EEsE23wxM
mR2yC5A8TNq0uwupjokt3VK16bK6e9UoZhd/sDHy2fcDt2Th1/W0abtRHdC+krS4
mib6+Mlsl06FFfsoEMWmzulWFixAfiqDDjRnK/90uv/jpE9cyelJiLJq2jo/2lmz
rhO6u3mhlAogSjEtCenCPwgbdYKc1xJEp8Qy7xC4TEtbSxXCOQLQ/7Z7eRw2TonT
cgqtaQTn+xuGji/uS/VlJnazSD+egslFynkJHXMxCGbniZGimvV5idj+T1pnXRNq
rdEisIHvdAO0ICetx6p2CSFGrHKatraulHmV0Eg1kCaDzrRU3qkW6/rzY/R/kkw9
qVKLRcTKHkxDBvTQLIei+ePOtQk8FiT9NT5ahO8jLVBIVX0c7fTp0CYe0ZyQwHH1
pO5SbWnzAWAvefCsUsQ5ClkuAiGEcFMUiiSfmlifoDAFq3y8EjFY6ubE19/d9+Wh
9K8Rg2ps2NYszh/lHopZtyd3Pn7g5tiXIQKTgJqc+/ETJis6Q/hGqXFALRrz2RcN
C0Os9+DouQGl5Kfw+PlfwvVAq+0gSgglaTf9fL+7kX8NdmMEhqJu1mxgxkehrJgu
e3po/8rLznv6WvQmccdk6ijOA66tJ4zWOzO2CAi5pz8Hy5wPcGtpXjVtLYcVyUqR
SqTMHMGVh8j1XwT1HXG3PotBiUWhqNLg+2ymg/4Te/9D1LhkiBzL1D0KVMCU+mcN
IjF+9hh3NEgap5cvjz7Z0jrZTA/q19KsYkUa79qtMWGzt69Niqu2W0loxtRR9/05
6zqRVoX2iwBJ2WrgV6hidqDcFJ72uztDmbFKUCYq1yFJ2w6WdG5rh4vwSElTReEl
WhFkaw7TZpYruiclQGZj/dwrG7cRKY46E2t8pUx1BrT1rgQQ5dmML3mbL2E8Qjjc
t9rnIQ0LfrJ0rkiL7/o2HE/LX1OeRa/WWNDluztZmdTOueAOjpwZsz59G23KUvWm
V66PWa9jSQJ2tgbfFyns6dwVvtW0NAGmW9G3aupiGIEeEk1DTsDDPifSqM0h5Xe8
Tb/IQMDVNjsp8VTC66bJZQtIJWLzW/zZy/Gk4+Yx7x6bSdmoqzHh+0vOvEPl2UoB
5XY+ITYaIHbWCmYk9HPG2bnOdQdhhAjAMmiULygiDSE+NeIVsggAlDokzvj9Ip2F
KDFZmRT7o53dPGEbg/60dbwa9EyQIAPPZyd3MsUUUGdW8ZF5nL7TXplKtcJ2J34F
9VGyfXggcjsTQjBRthIWgfKFxQbkWlAt7TlmNLj6yssNdqdPN6u54akA00d8z+zJ
j9rqduhEdr9hnI+rUlKo4MJprvZowEu8htNHdKpnNWuuPsoKoRQmn6OLOUt5f6Y6
V7gklPiYHqlXa1b1P0s7bojXy81ZFvAgFDuq3zyZpn3bcGsMGBTlyKi/JzgkXvUg
VY3IeK4tpJ1sJ56+5MX00HhhiOj9WJO2yJFpmMZSrFD5fSm8b6T8Ee5UvbsprCFP
+Gxi4D9J6bmvEuD+F9lhHYXOeDot3ehektedQqzDF4yH49AJTC7bYlhKXBXJF1an
c3ZvcOVOIxIHwkuBcK9MBtEH0sj2zbEtSy/y2ahE3yyvL+zvuKKu7eA6o06PCv+Q
NB4+b8VoZ3ZcsKMRhedqv9KTEgdMXfy0ZkPLTfQHpb+fqRHfg8smOOIWxkD9UuYD
l4Sq2V9O5eXXPMyBuKLtuli+sx8rLonjLUiWxuNHhXFJA9JuX2veAnW+o4+OsZTl
TLzXiuvAud1OYaCpRFU5h1CKPuVBda2rnH90c6gxICyf4K48bBJgEh63biRCjaSO
8xcn7ucPcQ75GVE1okeWQhKSbuT2gCWpZgyxQPTJpLjWwvMayy386e5BSNYnMHP1
IXJAXAI2J8TvxkJSNtgyKSAEn80+V1fSFNhX2ZqkvudRwVFNmP3Nvret2G0md8iT
XF8KGDRIl6iuRRKRpyna6eIrm1pRCYI5wIg3gfd9lCIL/QymnTlFA6i7nfKf6vD4
6ueL5YRiDU4GaMDKwuFhS7DjHyAzg1rqI0To0itJqRFyGsJBD1K8jdQBf/C4hVIb
3xO0d01OSVPKTaY1CFpHG53TTJRQCIa9r4LcDl6Aexjw0TZ/rFrrU+uTefDTHVZd
zqh9Nm1EfiupkSxuXMNmGJG48Kl7B4mRr5nKWvxAoIgLpVAzaAH6fzQVelxz7+Ve
19dLcwvtu/qSEdoU5FKrWQ==
`protect END_PROTECTED
