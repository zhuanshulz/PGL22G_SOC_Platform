`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bWDX30EpgzyZpGX53xM4KLcxudm5rCTxpnO8YqD7Ml1f3oT2wXmJ3IPFlw4CRgvV
Of1m//3l1mPNJ2aBGu8gUosUA9Ubsrs9IONxp48KWZS+EMjeBS5pD4Xl3ChAl2bg
Yn9WBk0m/V1ULOxvDK0Ezns2itHVSr2owI4/SuxqH045vq6zyCmwfkoB8hTxoZHY
eHqnh2/Iy0ge3R0WRQAxhUYJhkb5Fiihsp4EU68meTqfod2kncovaCE0QIJqcMTc
R77UdWsWswWs1hsvjKp27QUf4a+t2Lqfb68w8auFe5KrehKYVmV3l1n7jx8vW5Ux
G09G/ZRUu4jpC5WJXCoBS6B9o7cnP/RDVbIjoi9LPT7pi9EI4OYahfkymCAv7qlk
teDZ2V2YHCcd9ks6keynq8sPZQCB1ru/zRIwaWmbZkDa6XLx0bvGWlzZSUnAihCU
Q5h7Pd3Z//7Cx/WuMRFDeBQOnxC61sMcYXwugMop+ByimBamIuoJVjsocc+iUByc
RT9vtLm6Oix3ID8rV2x/7kCb6JFvig/owhb18bXQIiCn2JbOaO1/7LXwU1zUJYZz
95d8qN4Nf9gN1deAXyDJo+sJkHCtT2Y9ZeeQ9WuxYCxZmJAaZbWMfoYBK1CnvTWg
HBerG0jfLshGmPlH09QbXV9VxXN/5/1BNLpKEWegx4zvu1s/ER/3Rh94slOkCK9/
WIRpriKbesHZ4OkYo5/ikpWD2dZFcqlxalAfm3ZGEyDLA+ceUKlDf8w/j+FpDwrD
sew6P0i6yh33WO6bwYSX72fluljMRAp8Q/rlEinjycQ3zh+nsLVCGzSuqcHADNvf
UY8uWnMcjBOPCqsX+xha3sZEKAfpPrhosma1CWtIhlW0bOaMwjf7ZDKpOigvHw5I
extU1x8cK1+oxtXmp842HGbtRG16Uqf915J1xbgpnpWZrxb9NiUCJKeFN4m57y6U
XtM2yMRWHGShg8MyRuaxMbFjlgYv5ZNC2aZVb1TQiF61m98ExLfRKWJpdnjL1ir0
wEyfxDaCE8OeCP+WFfzoapp+br2NxbPddDTychkYDUO3GS85rVx6w1GPA4Tx9oM5
m00WTuqaLQBmC9FLqpIxXmVSqAfugHwoidfq7PkUPS1/MujK/vrdDYCkCZXw//w5
r+noDNggLsvBE/i7/FHCviQbdFtB794j5RXUjkAb+8+8voaoFvRRV/JWGTwEab2F
m+63DMS71eTYtPk14rQp3wUK3FGBrbvaUNIejAoaZAl/OsXVVP1DzTZbynIG6lhB
ezy0yN6KjCqc561z2/0hpX54FpNZiAjX398pbPUCaTAfyq7QwS5/SQZCx/fnjgnx
OT1cpE6+ceyG7ErA7Uw+jmhjiLRgc2yfo33yodeC0BZEOyLKdqHsmNcW6yadnMnK
O/Jug7/ZAgsVbXyAt0u9rt+AixqR2FTDkdmCHXq+Ko8ZkC5yNqOLJU8/XJgPf97Z
XRX0wEBkywrtJjyu9HNPe7yCyVGWXOJSQykGbegG8SQtx1Jr2QX1QvTdranqRt+K
b3RbQ1WxpUeZj0NiyQlPA53wiUEp9gHc5BpU7DHvMSuukAJPV/QKxVXNK/Y1mAxt
dzUHrBRH59tGLUmanLAj4oAlBnQ6DEWrloP5vBJm/++LpRbJ3aOQyXucRU3T5STl
FzbZHI7VPIyTLah97W4272rw+AJU4VARfjTsit6Rgii49ZtBIKzZDWwB8v3c6jrA
4Asr6p4GDCKYimw/Dxeg4Wc8QfdzBjM/svJo8t4fJv65qpP5b7uvwK+6JMp8VNf4
+Ji2875fZp5OnFD5sybtZUz8KMGWuuw2Z6550Au+hkw2y/4Eyyq3ofOHk3OMWC8I
zvV1TjFwY4CI9rgB0/wcQle6Cjbo1NId6quSsKsTMKE6Vyp7+64Mokot8yM2LbjI
4Rap51IWjaw453b7ubSJEs5QshO/OLiwwMsABqH67Y+2EA8tHy078dLB9ZHgd3+F
An6s3NGhevfwguZF8gFfhxYFw2+H0oFVagLMR1W50xrOW7ctomaLwDAea9qZNUjZ
xu2kKdOA4BppVl2gBHZNqzgCSc+xnpYuSVNpmx7ZvhmIFi8AZ8BK7iaE/wn2O/jv
2FpBH7HRAtU47ySHWorc9FCuCtyNrSzNCYv46V9Cd19BFipRVlMU20X7NlAL3RXH
xoN4NQ9Cc52X1TOsUqbPcu+f4gzl2XU3uvapc0J84iEAK0FGjzHFDSWxghk2D7Lv
M/payEp3eQ3do2oG/xpaMr4inwLOHuTWuXXLz9ZH29cGTIJhCQ4dBvSGTG4OXgMM
j17wxd2VbdNvtYiv4gr4KujUjV42cLWmFQhPYmOfuSAxY86VNWLWK8nuh+kyHFHS
J7cxs1Uu0B57xOGsh200jIIrQyXEIUO6YqY+ygcE4N4QeceNSo2CjmeGgC1zPUrc
H7A26EDT1bWE/oSuB8GqW2JzZX/3v9bZNE/7xx6dBZfee1PgiEdRXjaDFrZgLgwy
VAQO9lpeaThCq0i9ZdraLDXsebfLvO8yQoHTYbQvgqFeq2OMKxxCCybZyS0JYRvN
hgAcddPo0gbVrgdb6MZVuF5PNSdr0IWsMBCvzrCOYdrGuV9XnFCaZHafrWw8atq2
BYp+eAeEIxoVRoA8FwMp7C28kStK6UDq8fH8hQ6E0iRWYCdxJHVBWgHqSCvaf0B2
pzZj6GQKdTzRQfBae5t+QrojVgj7YuSwyvqRtH85oxg1LYwFkRIOA8Pzfc2eHGAS
UnfufTnKcHL0T9s6FnSxcP6AcA/0LF9AlvXJtQ97bYF6IkSxw5KcJCRHCv03X+T5
pN3i6cG65n8NjKgHRS1CivxJ+qKg5DDqxnpPqcvSfTi3mzOskHTh51z0TMsUBuDo
KTxwOBtnKtmZ7zwYXPaDgt990LXiInnt+W4G4ckCac62d3h3O+cUZ3bXiK75huyB
hOLsqB1B7fsVR5nuLcgeIrdec34eBY7Z+6m5Bcx//In3EJOz6IhgiWnX4SoehcJT
QHTeWEwiHhUGs5urPKGm50Zevrj19rGxzoA1xnNCsG7zOCRe0K8pyso94tQNgp9R
qKh+3pwmieMuSCn+l2SwtRAOg+C1l5JV4WIA/2BlVZCeSXquCvRjFPvzNZNvspph
sbUSGBw4g1bSkGxnbqlDpZtaPOt4oWUP4SzIhc1P2T3Ric8IZl5AmK37BM3DEA//
IJ6dR15g4PLzADu6utxbbA+iNYhwcQvjeRLWkQXu5a3nWRkMww2MTxkI/V4Drm7P
dn3A26MR+o4Kg8JV8/pSkgTIgVia40WVRqPAtXt76MCQYIJvsILzd0w71jke2HpC
LchnLHgUkRKcdnCLoT1bIMoTLXep4Ryw84Qo6Is6RRrUffIwTTmNcn1dzZHLfpln
/P8CLxP6lQl0mAz/Qsx0UdDH8tiu+uGpbFlaThn+Zg4b1EdHKLPuW0TYOwwQOahy
jCH3tCt29gtbc3PkXAEFtG9PiIoRrOUOXEz6ToKQKr2UncnfwVTxHH0rL5XNEq+8
4RdFFf2P5TTpI5J/vYBBLkQbaBsiTlcLKaSYoSoBFCrTBlBFZnTONqtSHFCw8NKt
mM/9ZHHHifhKjJhj9iNs1DaxTe+mEjDlgc3gNz3WYH0m4kipJC9ZKuXp3NUnYVqD
v8o/18C+Dzfhxq2/yCCWpKzXNJ6chVuQLEuDKvg+kY93u0Q7+HIShf1MR4bu+E4Y
O1U7xaRLJuhd7SeiO4QwWptCbJnNPPQOOTb59yQ6MafYcpaR4jbuZKdEnnFb0hLL
mBVeEAC3m0kXwBAtX9eLe48JOTxryY2tAAHpnJvu3LWFT/sWkc77ewFVGpdDHcxG
Oq6KNh5pBG35KC+75N6RapDets+C3EmHGvKK6cp9lC7UABbkMGpJzvpGNta/zT48
yGQRcj20+oXvdQVTj5qShVrcB028ktebF6tbRjo2jGi/mY0QgAS2JahDH6JsDadu
6v8sZeZc2vL96FunC8XELrf19KWsfjI5PkYvUxam/KAAHe9lMToMypkH8waQLGsa
0cl2km5BBWi5FkPFyEY6rcRezhSlnXY3E9k7I+NgpR3jJSIupU2QbK6jrqZUXQlJ
POfkwuh2843oslmpmBdhzhvzHG4O0Uk9FGE30Q51FlaUMUS3kcjx8kmgOD4mENvu
03JFN8Xw1mLxYt4uEjuf5hPfjWn2cYHNsZhzZjElz4/pKlB1rY1xnUX3YvNsNUkW
tjYCiFd/MBwBWA2wqkLvoWX21BtTPHSONcJx4MVF8my4tzmSc5YRBnEJ8ZDOtJxO
41EZnRY5SzLA8P31n9fcVNumh/qw7VzC3G8gKmOzq02xK/CDfIWma4r+4L/VZ2tT
eQN8fu4JDsWu472qR2ist7pW3+N7SVIM/O6xMXzbcfO3/Fp7/6Uhe+uZnptrf/rk
qYdkrwjn57fbeE5HnvYwEik7zYG5KjL7t3V3vrQm4MAkmXohMi5A9uHZFggbYs02
KuDCMQvI4ymG4mwrkyigTVFXyeVtbhpR5cuuDzJlG0ftYQZOv4dK9xUAgl7FnJd5
3mp6o8lWgan/4nqPnEK/r7aNoWr4y5DwEHKykaAPgeyoMhpKqDacpl0GdKsz6SIz
YyaMN9qbxLcbEmLjs7cKpjiQlVwkNKCf3J5mnIau3BRWxdzpFeD4scWhxfm/zyCE
4PU2ZCMosduWE8qvjl66VSRjJzNt9V+teFbOckFtBdMnb1b0w3hYC40URcpq/oHX
k7fPZ6P7e099i3XKumFzS5LLCA5QAT9WUVZyogO3oLZ0S9G3E7GpxPjfPBIqu3Ls
KO3mgN2cVWsZqCgJIKwl57c3ISu5a/Ih1VcT4Um5iVIWYNJponmQnrk39dwIMZTI
6n3RO/1mZUisaYhUzmSfxC7lFsa5+Eb271tH9aEzBl4ZG0OYihPyHHLbsmckraMa
DztztGPqJOc/p8SpvOGJdJplMBz0zMZwkysqUhvn/H7F/BPK3wH2NYRcfx9yk8Uy
jOktbAvWendpWJKvlVIs/aovhD6Nfmp2t1NXU/Q7rEOAOfbuhsqbmQOdGBP3xNE0
3lCMDcDSo7nppEBgZZRtP1Jf4WYQQNL3f301bbYV5HBUlWEGnjsmbFgdqo76YX1z
dya7YZcHlnOO4X/HFAtnZdxP4JL7sM0T212J1Gqw5RckYT3BEfFgo+mpL19bhw82
ogEInqAHD/4jz8bDPNXrI1TpqCqfjhtt3voZo473wW6wmXL6ztLb5y3Au4T9stUE
7By/atTtjqD9FhdZrfElpioUYNZa8GDN6dxM9GRWGCTgEm7Kp4io+6UHXpNOjvPJ
LHaOUJYujUDlLfiuICc14rEQVQW5pQB46KVAtnMrXsp3bNnVRFiedK15ni+VPrgH
29k1fQ/3vEcrbRlg4MA1T/KVOr9vR1ou89RSssj6BNuqt4pPPli/7+VeSDRgiuB4
0oj0E/NWF+7aXqHHfQ6MfZAs39luI4RQyGIdD6gZ5UwKstlcnTTjL4pVOUjZ5dNY
59ewwkLnQVH1Yr+xJwjoL9FQubdvTH64tPAoYmQu2D95M4EoF/AH+VGI3kTm7yWb
f/AZwDH0+Ry45+zItooJTO1AzCEfAKZP37uxQ4xE161hSHh7hhf/UPmqu1YuqYC4
LlRgqv5MqbSE8gIlHZG0aVeNZfF7LWYUGxFVFVyc+GETGkuykQWQ++kRYUFSCa5o
BRvfBxzRXpKmYxke1jatqIMCupg4hZ17080bGH3FGwtkMzcFXSu6N+h/C7CTcm0f
3TDScRTruWcTM9vbCzoelE8AYx9A+72mU4RFP2L/czYglqmlWZteB+Mr+1T+Aam4
Jqoy4pEqsbIvkRHbJAPYmyij5+DSFk8nvCR/Gb4ahvo58Rokf6Qf2doKO+RQqABR
siCEPnsGaKyFdH7L1FoctnMTznfaVgefpqZIwK8TFY8I9FJINxfqaY7FPTzFS2fE
IBzNRclZzhW3/FCLiY0MHciv+ah04x4J+HYvSFCHTHMANgIVhp4v45xs5yFeouKq
Ttcv6DUnyxT3LDXJ+IMGKY0HLyLRW1T/hCdPK5ho3pmdYNuAhlQQvcrw9I7nyG4v
coc7ClhMRCdja+yxYXerVy1PNwEMdqnqIPtq6nVzmiAsAUkBzgzVOh0Zb3l5LcZA
XBsGAzf81aLM3xRQT2I5MiR23klFDT1cKK2KMjHD00mLkjsduEDW/gDBDj7zM0K4
Atmq/JMDR1c4ddenY0IH8ESu67onWZRFJzJqeI5ybU8rFLjYj3tjijO4p+X5OecV
MP16bpPeAcDvnjaBwHZHIrEhZLBc9AeziiOooVHoKaBZS1QhHGB6mcIdSxch3w88
PIBtXGw9AB/3gVJo6kdLPgM19TSfNs1Rc/3ohnOicjwtvSF1a+Q8nB347CS0hq/h
r8nIsMxEHH6aejVlme7T+BLd6Tj6b+ecYQbnZVlE2gZKqYqttvVY2AG6Kn/nsEq8
TlcyiCyaTty4+sFFC7faeickDl98tFD9z3uLEXFZmhWLL7ARUFHQDbaRupDAQpYe
3EF+QD0u72eUN60UCxZpg09YbC81y6LStKzQKe/W5peZ+OXl6BUAZ/MKY51wsRMU
hAPDNgVGwYBv0uLgqQLeqvlHbAa/MLtVkthGqfIMLEI0ZPWmbijB+rieMn6BxdC9
XefmK9vLW09g9xCP+wutg+u76QvGsYDcbNax72jCOzSOZsxzfUgfNWabYqX0a+p2
fiWM0nhk1Fpf1GEax9kX0P7iDrO4j1OIfHo1T5toR8piun1pZekiNIWBh2H8GW1z
VST8h56uj/xxkzYZfkecy6AJMMqTSm7tGr3dlrqx990uFN8fxy27kh5QzrzhyWZJ
yMiPcdPoOEs4VWz8xzwJzI7KjpKSDgxBqyOgxySqMoSKbwPeuqFvbnToUuSwdZUW
y3r/Po8NRqu7zMNrijS6QB1wDTRXcXZJpEmZG4m2MSB49co4yU7Ralrm53R5wHD2
0SSrO7DyQD1VR9W68nJgQA7f6YCSH3I3Xl7ce8rlzsbOaBH6AwXf6xnuVCcStDLR
fmvmq4XREHl9MlOWvAbwga8h8RrEOw57G8H1RfUSQZYPcmLamarfrjURi01Vm58a
0lh9bWVaNQQT63oFsVmA9scXVgu/FDVY7xULf0rVyGBZY2Is0XjZPf4IZRiRe89o
vmKRDaJJk8R3+ieO5bU5IKsQP1UcAL7b/3JG/1MvB9J05fbrf3lAhngnfQ8nGsIZ
V4NxPsrcl8C1HqDsMlVx4fJXR7dDi0BWH5uyi3eybv/iTAS/E2pj8cD+1y6vv/jE
JoypdYeCLwn0sGt5n5+5AxkeuP+YMWrSNsjao4cE2TF9q4I4q81YLVUGSasDjS5d
QIvWfXlr3/n80Bh9cfbBFy6HYqvsJ5FovOS+w5n9yE0Ou2G6Zs9jh8aRBgQDxDIb
Hj9qdFyy+VapXFmUob7wAHiecwtACn4Ht0pc0YT9m3d21t9Ql/+FFxt0NxmE09+I
fa/MC9wF+6cq/WS258p3xPN1YILUsUvGvr38TyUr+RAvdMK06ttgg83GsS/4FWrB
9j2SQNKqg7hci6LFxm+iM7gFqQ0Sdi9tTgAnE/+Eofjh1rI4X1K6rXxXenD/8rbp
jn2nu1VC9rr9F+tOsAYhnTWRywymooh0Fo2bJKPIG1UH220XB9WoQxexBr4MxhbA
1IdBjoX0feeLdXUodlZXsQKvLgtlb177C5V/SgEFnjTKkY2E8MrNOMItcbwLijqX
uUQyxqhAySk4HbweXa+EIJBp49N5QVCtXVEMDhVhp4qavKsHsL13yXDvILCV3qh2
zWMeo960v3cqZmdLJ+tm84GnYZkd/EB+t9t3by6ha//QPWSG2ve/hEwh/wac1PKm
o/RQpHUHLXZ1fxiMXUc657QbDjE0sc2Wr1A+XXQKlkMzDpKfQEO1zAWXRqXTJ6sQ
zoSXXsnIhgnZIw4Bf1k8lK2c+yps8wpi9+m/VrhIDXyGCXRAOFzyqtzhxo6Hm8Ud
HBA/pBgpV19jC9tn7kj7SDNdzZXalR5kVVY3ssU5MklZ6xZgpRa1XANv5PtBg6uQ
sjRlMuSs3YtsnsgmKZzDNbgxrLycxHA568mk0ZblYx5qVNF+aCGyHpQxoPbQofq7
RG2GTsfjXDgDruMhj71U0aWEqIDU7ZBiDGfAT4F/oYY3GG7EmBZrRzhJ8rn15jG9
Y9FBl+tIfpDt6DBQl9I6v6zWupjTCDX7bMiM8vbdD/QWRY6OhTCQ6ot5sCLp1L3z
Sv9L65WtzVd21zf6gaJjj/evILLroyEC1kO9h/CfQiizCSIjvd5tV7ImQVLcO/b7
poU5/+DwDb8wUp/sRxKN0Izra9jWCfSlzECrMiz9FUiq46fjL0PlFCnJoMaA9ZE1
pNwiRiJtU0qt9ijBy0nKmdOkucO5attCG/avqqboA2d75DdxyW4XuUTQKk9PCt0V
YLywMdODfe+JGbfuPQyxsF4mrHfRXSE8mSJuRr8mZRDVxrwkgvpzNXlS/X+5y1Ao
DQAh1ZN8uE/La6JSyo2JPETTqnBsoqD7weLdF6ozyRbKry9D7MrVt/EzrlRA7kRv
WhJXlX/uBFw01NEEyOfAPcA5bmErW/AL2Aq9QpFWw3wMjAhfYH82JkRrhFP27Ya5
1HnW9uNYsNtY34NNwizb/1CpTb7obGaaDgxRaZClxlrLTCSu00BrvSidqX0LkA9y
beAtdh6KKbKkf6g36HFughKLcqJIWTnRX1MuTmgLA1YOpSoaCIB33dCHcCU5R+uc
QaM1zEPi7SPftcCs2UNUFTeRSTGww7FzQguXgm7DF/eGmCbRV95NH5cOmvkDK6Ak
oTJq+ULqoCaZRqKHq3K+REkv8vefTEho0ineJecMMRnanI0Se0Fmoxe4G990FjcN
46GppgvCRZj8fppyG6DjL6YC+4KccpmtCsPArq1dcg0OH+HH6M1PMQY708p2z2hk
Jxfh7Lca4/11WrgtUFPyOB7SZboSKN2rbL/3vH6RSI6hoGg8939EOgr2HqUmg+9O
yh/ZfHdhfU4z0J+zeLDvUSANy/IAwB5MW0KYuD6ietZa02fXR9/0SOYuFnJ8j9Te
ObVK48fCU+ZyA0+CPSzu5vw5cwQBmr/krfG4/sVOmtEUXstJuX801KD4WFJaWYdd
BvfPernUhGu+feDuc6mX94W04jJ/bB7zpfao/kdSHI+7Zg+BoF0Uo0cJxTA8kntZ
GbvNdBLqbWcqJw1xGOn4tFcR0K8VJAQQZ246xW+QdaUZSDIvbhGoXzATZbHPoL6x
lYXbL69G2aA1L+sDwINdEZUDAyYTqbhp3nUm9at010slbgGntjeUzZyzvIWxVjaF
VQxO7m7mFzU6r4/sTpRASQP9cduS8QZU7KRX2QFkHgUBTDlmkt8gc0ddjS4PCj5g
qK1sD/JzGWqWa5V5qQf56EcjrmDdaH3t2jwXJXdZwWZy5oQTBgBdQtpby0yjLAF2
6JnG5NaWLrX3z1SVHMCRQIuu03mlmbqxbR7TnYUmTd9L5JWfkAe7btnQeVnw3ZMB
tVC5cjLqerYCjm2818t2hCTpO78xRX7q7sG9rtjXCT0gIqV1aImYuQdzNiLNypyq
KHp/7Ssy7gSmG8bBK3S0p9S7sU63xHfUIvpE39iqreH4UvwD/0VrBms31p4St955
wjUkTuuDHtwXyIuOauHccSExxdZNxr+tT02GTOkdiFKM9PJUuuxFWSEg5tQOCUzs
+uISnPdZzufEOojvTLF9m2gPXdsrUrsbnFsM4FOwqqgs+N8dgDlwA8E33bksniNA
MsmJQMth661U58f+1iqkPUyq45lRoZf8o3pqcAn92F3AmoHNPJZV968FYr46j6X5
J/Jvkam0C5DRn0KPMNdHe4oqDMXHXZC0fIMUn79yAoXKzxqpxI/97FfFtLnqVVab
L8eOddZplz6Qmug1lR0YzjrwbEYm/G0pEZAHtZSF8rfOBzHEN+YS95R7Qf/vp8dS
EXBjYz/05CxIUYBqggxsTgeS0duOkzW5STEndCbvFsah/q7UhEbIIT9vMi9UiTsi
dvv/q07IGu16kyhYrBcPIOJVCzncsQV8oGAJwkbWmVXasOPpCVwC2bmIoEPo9IuG
n+j7gNKuvYDW0MCcfxv4z/1ivPN1Ulk1d+NxTh4v8yCu/fl19QvIC4flQcRJ8UvY
bqMeVipo7ibo2UmXRonyxZtkGWB4K21dtLPjmos3RLFoMU/79kfduppFfE3wR5Cx
X/+VaK/ruBmosmQWrOED8Q==
`protect END_PROTECTED
