`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l0BtREDpfM7k/jFxLvLzRhrtjtdk2r79JgueaaXgBnZE4CirhvPcr3847P1WdJLn
mNS+6ovYBod4dB7v7qpogbfk3F0T5Jn/3AgF4gwXSKFMPUvZxcN+DZhI9fBganJg
jFWUGVIFLIrftTICV0X8b5XQ1gxX6mO0y1/Xfppvpvq9QLVVzBRn5h6wWuwwUccB
eypZ26jJfNpVkyq4EaeNWTcyok6+bbZYXGWEgQmzIIHe2RQSRFrm8rCZzF0WMTti
3LlL1LhmKtiJ3ulQLhPOZzjjnMkiM0MfF0vUzvGBGjsYiiWnu1r0fJwJfz4D/EnE
qEdo5NCBXcg2pmTi8p3dVBC/o9D16H+EiNzHXMSHpFQ6L3ndb0X0ZZzAdndxd7dz
lmq7qiNCnT9j7IzfgYCWd7uwIvdURAatiSKAKaMNAPRUByltEgvcPKf28C1uhygy
uGt0to40vMLpo14gkFbKxoH6iOSt7Ldo0Qai0VGb+9SWzqWqFxn9Nvu4uPSnu2G1
UNpWPKUWr84WMuPVGUszvprt+Bw3GDQdbyYA4t6Uko+bzOxQ8fmT0EfeuKKup6tn
NByB85h0xHuSe8tFVxNgydfla2ovKlLp3RECvykeGCVkYZlUxWfpRVMGfENq8IXe
cT2b8H9IX6heqkgDXhQfd1dJonwPou8PgRTMtJnWhnlMjDCbtdQQV5LxG/vTbMrD
QVAnFc4hFReryWF3S7SYtvKe1S4s/QopN9ME0ZIY+QwMFy7amQ5RwgTEkwtO1qAg
Lp7yCVOPi3fg4T1sfl3jSIj2l0v/QqFZLDT67umImpu2WgqAhuP0/XQZiWNt2BCv
swgErWOTNF/cV4YF6EpzhgGGv0lI8YklQQLf6g9jgILUQV+m1lYq8Z4/yPK1xOQb
puNwcljE/wBhYuuE44L4xoM3DfYyNX3g6GzZtTm+QWFkknxqtqeSmif95qcn05xw
oSD7Oq8PLW1iXRfmo+3LdoaqG+5WqUV6NIaQREM5NtS+ByLJV7ZQTJM6vkZGFIdI
b66L55qNoHLIBHfnji6TPfCtd89nafyStRZ4EV5ZoXs7axN1bC2fT8SU5mGNxVyL
+RffOuMPCWnvmVfp2saqwksnWAhVUY7bKStvymU4o+PqqafZGu6vy2TC5aNLeQuT
+w0cfiFa08mag2sks0/LoCw9udfRpSlXLcfpZH5MQHw/0MZ0+nxIW0RFww0qttV+
qg3HYRdLtiTnV9WkeAuLQT22uLDRo41/swRF+NyVcFufG5t43xs6pyBmMr1hXmnZ
jxR8OnxREs4SPstr/KN29i9Uz2EDoSp13n05GGSghv7qVcy5ANmimiKqdIx91KGO
72vmBLLeVed8zW5MmXfUI3ohry93xUkETSkbnOa3EhKIQkzs8PQcE8Xe4bRsSPlX
vhqWLcdKcYpe0Dh6T9tuKvKVVoc0sNTuI3ZCNkp43csDsLcqNei2/pAb4RLz8bjb
SSs1HPXsmFhPF/N8ZHA0fE+FKzczGeLGOLuWVsq++1wua3ippZmTgxg+SW5BTE0/
OJpdU4IOkRBdgt80IABp7aO1/NEmgLpjYnzruM08tusyUcdVyZWirFq50m5VSB4B
tmadQVYo8d+P2p6xdDAudQs+zCUu3H5zClj55rqCojZdWcnsSuGr32VFmvhuYA/x
HcveY9NISOqMmBwFe7jUdvdgoV5cm7TLZ7vTp8aBtFUUbfCyMGc1+sZV3zXykXFl
VwpYPD4MfiQ3GDxYdcJF6PamqZABOHBmvM/U/AQLoOipdfZMbneiIqNkyRz1iScZ
rGbjq6g8IBSJptb4n3K77NgFhLPZsXmta/pWC6LRu8xLJXRig2h/NJp6EWBXh5SD
l65dmLm5K894bbTYGMEyYOuhCZx9jBhM2gsIOlT6j4Ob+Zk/6wv4WOn1Sktje8Cd
NNzvZiV13xTssqmiXi5nqa8UNaA7Y/DY8j7jAxcFYhewGTUz6TIqzWGq7ass38iu
8SJGs8fxhoa5fFe30JvLb8k3JG5V/zTPncTEowkVh2LLnKqfQ1nCpTbEYgQi/x2+
LeGiGCtLz9HRxCL7QeFoc0gcqjUHaZGpM23DKRuThUVXpTeehuEp+iHR41tjbnh9
/2FOoh4Y9UTQlVjUU6WLBtxeT686vEOrb1w2cCQ2cDLjZGzFxmse6iUnihV7IBXm
XnR/CeZ5SRk6TBboqLKEA2cKzJJWi8uMjqOVM0cUZD5T5AJA89YBWiUoiSddA0IM
cwNDQflPgqLjrOXomWPHiNf9oovHtJ+5CmapqaGU00t+ZEHhDTPgSRJb7/7LuAYc
E1cQJLDIoprxRA3xQihx47i/0dBj+lYRu0/sRZ8t0dnGINhBWMK2f7CBIrQxZ2E1
4ALOJAtcukS6/YhEcKVLhaLD2/0uwVCFQp+EX+sOQ7kvFWkehpXVvX46K2Zvn5Fy
6+6vECvXXWnJp/4a63IXh6H0W5dWC4ZSIZMnK1kEHMGtxVdQTySlFEFT+sZn/c9n
iYIpkXOAMYPXGgZpXjs1h1F0wTo0km72mTNpwZiMGEOnZwq22ulOypYznRJ1hkst
qSLky6kffK9h0CX1Y4BSPXLWNf7m5qUffcJPekoIiGiev2sxAQanB8YU1hRavDtM
lMhF9XVPMOcHSxP6ivWu+5RhsONaCrpL7kWs0VHGhk2OKtTht5cSzI6k2YxEdTF8
mMvZXiC5NMphKKNy/BGyW0vWCpLOAkos+SCajwD01aa2CehPMcRN+0aGF6dB/Fci
0LuqZk5ah9p/qh8Fd7t49sLwrVg+D8lDOF4MUaJMhLS9wpCt2ncK8hvr9jl5JrxD
opJsqYG2N0y8EBRfwypimVR5Z6f5z+Vl/ZMPmzgPuYVzgjVnGe1EHJnuATpekA3D
WHuxNg7XwW+CBAxAzrzxJaX3Sm7MMTRspUxdvGvTgxyPRCuG/1BhpuPQispFIaYe
jW4TnQZ2s/YLy91c9M8DWNKvoMNUYUs4HPDVbnq20kGsq7bdKFFda/IbOO/65Z2i
cgIKmQoe334ObJz7bWVe+LKyDmk9rPUWF/EZlIClEfEn769EcRHPdBwW5DbZ+hG0
69xTDO+s9NPMZyKuu7s/Elst0VSf2aK09ttPmxS6kU4CKxF+u1iF9GdJpBlZEJmK
ARQ5bIu01qSYORWwNYoA22KbKRa9NVDORJpTRZnLpd1r0O1sDPhd5laFO/Ab0Jh6
Nfg+bIN3rUnZthdF7WHJYS4kbvTM4yiVmXzX69knVJGc3DViqoMJsa+w8s429ZQu
/9NZfUhglhvRGMx6I0U9C4cu3kpWH1oYQqMQAmgMz0iK9k639C8TRp/A4SsUPg+2
3QvlzL304+n/65CFra1PauD4y6ZfDTrTXY/9aHXfIjF4bwyK38nbT29aMZDpKN4L
BZA8y9GHnaMKLNJTYHQ3bcZjvSSyy4UJwvfY6VRmyNSsGH88onqRWz7N/0W+TJrR
cPTj+uhqMpuX8vlRVvMTVybtL5c6q9do4E4jw/5PRt472XxV3XC3VYHf5BFlU76s
8m+Yg269C2kAUnzEnQzS4JfCGooN8HwLrVlWIsm8A1LIRM36DRpkrJt6y+rtn13l
ZHeubMODyJkSzxRmhmPoFELYbow4O2UDkOIqMpXtQl9G9r6OBG9IjzXAmBqt4tTn
P1tIJQQA8kC0Q+4swcsilhdd5EFTZ2LnHIidFaeh54hwmlXt398Y7tV/iHv52g5R
9UzxJZ+sPRQA1IQW3CM6ry2tG00WQVKB8RL+XBlgsKP7hqQ/hMGRazT0GOnvZV8c
Rt7OsTQDAl/LRTwHYgA+0ejjLEAnKUq/PJPgttkANMJJsYwLzFkPF+hLc+ZbZm/n
5ofpMVn2FklxgPqkDhJRnX04qkLgHwa7KqsJidS/T9Hi3AvghUb19xQSQYsP2Ask
1/3PoZJynFRSRh02kCh5nYgBC35E4KGZ4R/oZrp7IlyjS6PcvFW/IrZcSVaD7Ouf
ukRJq5ksSm4oKYkWw/62RYFRLZbLT6kSqXgfaMQ1z4P+p0WByHjQ7LnBsqphVYPT
BMn65Z7cK7VCSLvekSXST24Av52Xi8npb4Rm+RFkDA9xqeqTGFUawybhNfShcwAO
aoKe2M+lhbEFeEx9otm1ph7Zk7fkUGs6aCEUzaSj9bgsI8kFJoKyzMX+RWwQSSuX
kgsebsJ/I4gbZY7ORd07Ye74xndxN3t5CxlQbqIqfyalMvBuzM+BFMjFN9HC//JV
SpJPwewUw4knCPyIzsmNvFs5+6aNLCCUt7DqJZp+LGhF0NWVx2wIKlmfd3IUkLBN
GKL0rYgOJUKtWL7t33eZQaNvAUU39vgwHaeasWHFANVOZgVEj2eZQm0W029ruK3X
TqFpnpGjeJg/JBST343HbmF1Lap2SdJx9+kARzMYhmcS90od2ezsidpTJXyrBZEu
s4GmAMSddaVRJ18mujgafY3tBaiEM0TK08PrdmLZvZUNT0rLjj04umnosl4nU1k+
kCnSkx3TtqwoqxKEc/3jknCrwvOBU3HkaRZh3aoPBiRmvPQpl4oRCFtlw6+K2KMf
0un19AlLyOswFUxOyaiAb0qcTrkRKPCKn2wOMJWz5weB8axHtbRXhhYYfs98lb+7
AVL0VAL2ncfznaPBR1nTvutc8/TLCXhsLXX+RdvWCACpIPGhaiCO1cWoQNIhZyIF
x9P09VswMT6spsmO84kt2SCSy9AIhgKeIm8AtxWNIuGQxQPZPx8e0bGRQt27w/nZ
B7Y9LIR+eWcfP7kJHDxH11MV0qeAukzUNwCWtiT+fbKSn8/73PJdm2LkmSs3c6WX
GxjsjeriYtom9bbn07hBvc4k4vhEkKXxpPU6thKaPQgbwV1PD995o+QYHVDC6PxH
iEjEmoduxBAzLnT7znAHQPON0CLKBe1IXxi4tx55W/GQz/rcUJTeU37JlWuXWk8R
OJxK7WOe0SV6tL29PcXrlRMgNPlBI4w1ZagmNWyi/82LfebfnjR7j4DKOFRgRUa7
22TLzXR7yoZ8d2CbnYcObYfwQ4vxDLmPunjxx+F/Vyu2JsU+rmVlKp5xCYo2Hqi/
3lDYkgnTXThiPis6lPkVPJewCkm2iYiPd2c3t/Q7YeYO2x5C0Sa6XAMwkD6KEahY
nfeFV1YvvDMleXwDUogJmN1DdUBdI9COrVUF9o3Jo5Fi5UgntqwbdmyF4Ipk2DoH
i0d2bEEOlyC60NKMjiC8cKYnNCK3gxv+Am0ZYoJzCNxT7y/3aV4Dkn8deVWG0vcn
QVEXBHiena3tX9+XMANTxEEZEhZufyS5rE76r6kQYR7tzELYpv+mO+hnRg9UmM05
WaBZZcx7yxwZbwhMQrsQdLtO+oLYGUX6nOgmLWYIU/N3Hnmg+Kb/znVpoxUDmNpR
3N4Iy7zVHPD4/A2W8TuP6azvxtwaHsyZFl/L8/IEw/uUozxaRueSG4NZROfaM859
jDJV2au1YHGaWoicjr9VxBMg+ilg0VYuLkEVo39YNKTzvxF5bdbpVQKvaP9Q/rfk
1x1CqWuBaOA5J5mlHAbwS91FnXmsG7cP4q/ntLwzQn55uy3BYRqfPnIQ9D0SJi/9
8FF6gnswUzpljP4R573c0W992LmFbB2kJ6QxnzNR7rkTORttEsRgmt2YWje1khqN
/s8YKzuMLMV84thwekmFMggT9EHmTymApGrqo1TyRZqkj9NiSV0Fj/CnIMMxDFM4
WyiYSwnszvK8FOOhJeZbYcMUuFd99wmCgBJizAtmESrLD0sRZmo7B+8QQ/nfIQJh
ihw678Fvzp9XonkT/MjVa8gDXsAP7xjrVPOgEKUb7huCh30OcT7BvTvFM1cC8xk9
eOuxQ3/zotp0RFvX2WhhyCfMmjcfOpAbPA63gQ9sSwtXD5Drqux9wqpEvdygj2+X
Ozs3tqcyPtB6wsLNm+RsPBQElIFY7EyLO6qPJlpky0yFVIwfH7UVS1jSkTllnMAZ
or7/J8ZVnMUvAkUYkaPZFXP8lYOQ3KUDzpp2IX7QhTNTtpsR6Q2DDHtxs7jVX4CN
hmzrjKwtY9oeALZ4JMXOiNbZWO+zwP8poHvgIEc282rwKwydBlsE/zjEF1aYn8G4
h8mNxPzNBgcOwA5DX56CgiyNucEBVAFClMfj00ewSnM1zBJZzNvLG+UR1QdZ8Ez7
`protect END_PROTECTED
