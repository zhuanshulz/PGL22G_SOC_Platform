`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5+tAmTmy4wOBoj93qZIoBIkHMEu5nAX6y4HxnT63Zlw0N7NyIXGmCzxpfiMDKoDw
mVbF7k7pTOM1m90qd7kPGhYc3tv5V0WBH9s6Z9MQPPUf2WqlHKfUSeEthscXNQgR
bTojpCZ12vTwC/EiLGT25I/8bVyBC0ggWJE/dTvEsVDc1kBVHjgYdj0Sawye+H8i
AWGXDWrUtvL/T+Iv7y/1yF2WBJmU/tqR9s2J32aq7D0ZlPdeF4lPwpKZWClR7Ull
lf8+30y3Jh68u5Mf8SjYOXRu3BPnVFf7EWqUOxVzoXXK19sr7z3dnB9O+apcSHsl
9kYa9WVAC24ME0B8Yr3/NHdNsok53k6vncYMHr14MbUSPmE5cGXdDgbhOgk5J9Sp
UhzIUOyH46OnSKvOFIfaMor48gkaSr12g39veaprSOzw/G6yOi6l4RIFE2L4/S/A
JgL4W8SRz2A9zTBu5EX5RxHacWI0MQIDFYrlCQcGRSEhXukf3cfgijjzXOpCnB+m
XVDoiL8R/OEg/2rzau6Je7VmtGitRkUeREEXrZqRCUvOETCNPpFyTbCW75YnjH9n
Dj4M5d19YuN/eKtqC5wkKlwX/mLnGTDG0jqdt08g9N4=
`protect END_PROTECTED
