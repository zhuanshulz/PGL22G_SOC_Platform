`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jo7wcAtZIk/qD0Va6CIkGSFKL87nmgdqTNYRKejhb3iqXfjSLEfvdVfXhLixCat4
OQ3uOLHif5G5wTOA77ROVD1sL02Zh2fqDm5qe9ZcVDtrQTE4WaXRNqpEdrpVzDLg
T/LD7lyDYS81DTtIEDTLa8fUCS6oVJhcmcxgE7iaCsJst4o5lH4Z6QZ/bHO5tbQM
uJ0lLckDagGn3QgmXJsErMw8Giz6SGr97D6Cn1/yvtC5sLChyVd4uMIl1YIorywt
5O0dWI4jkGCxeKhp6KPqCZJXxSYzv7lfy/O8d81DrI1zCMMRdEpowexX6vdeCmEa
tJtiLAnaRpv35Se9xelmoP4ilHQ1lQ1p9OdODpoO4hPPuBekExiHShiObBxsQwRw
T1C4fPOA+bhgYQPwXo5BeczuSwluxw8gN/qCRsvfNeelnSzoIR2f0K/8IW8os61F
HS4MndEFi9d5tgQ0YFbLY8n6ywvOzUOMSJ59lbaZwmN52KEtyxzuTLzs0tU/x/Ze
DEC2M5n4p9Mqpy+wfU/YdskOVnqmjkl8MUMbEQWZpUfi/SL43SUAq/KxG0bSKTLD
4FStuqYhfHZ3gbnyYAXH166+0hQ52Kk97vIxCGyX1wb59p8oAV/fuRxYH0PrrI1t
ecrsTkx9S3NMfwyvrwY7oWPOQo4fwdRSr1IKJJXEPNzzjtrWpvkYu6w+U6ut2FWB
WkuvqJCTsNgV7FRLEFnhXkm6kXV4PohrFxXjvCMZuu+L0v4Umes+YfBBAUhkAWVt
SLsT0N073ovymxYLdQoP8TTjN/vP/InRUY5MIsDJiLvn5/PQxl4JSbcBtJvFiToS
AZ5pubgB1VlxsjYPVH0R6E19SqyVDcPQLKGeZOIQq/+lbUfkYE0aqu9Tpk7Xz0++
7L2E2VxqD+TAY4n4NFcWmphruM+hQ/Xa5/N4pzweBLKILsK9qDH0Nh3uLjeXCTMt
riZOmETCha75uGQ1uA7oW1CtawAWXjVMzUEUufYbOyUG+x7RY1WC1OkhNxwsXCVn
KQZNhXA56Q5Axpp2ixGOvssvn4QfgVblmg0iEkJJqDpEb0/D6D1gE84tLAwiLQGn
qmqfe9nDJMjvmI/mFzjwBxOCDYks55yff5kOOmxKFsOSF0Xu3nbMQGnSzm6qbYsW
sVfWYy6qcFXKfStECtdE/ND54cZN4N0+scVZgPDCIzGOvRnp8rNvBJCHYkTR1ypH
fSAEyBsr7dZV3KpITkONNwgIRCmxiO9/LU6O3YwthX7JyvTa6b9QiAfGakI5atlh
OvUCfbYCruqace81xDEaPBJxU1zW5SP+XvjpfGwHDn5es5qEcmUKdcnLiOdqlc/L
96hUpyfstH27n+T29hjqYQ==
`protect END_PROTECTED
