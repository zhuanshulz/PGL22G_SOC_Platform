`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PWMk8CgvKj9BFM7iyEHFQg/LKAcI7JebMnvUtg1PvnED0wV9+0vpd478nYervSXH
xiS0I6jnwht0HrE2NWxcXZKsnVrzsC02hgkoZ+rydskZtNv/9j1oZRUYYFgAJKy4
FnP+FXpNmlycG9YLuZBjNMuxofwazNbNdL8w8vAvvjihDKImUZFZveRrJEwei6gM
pNWud7+tCB1eMZ9hEJQ9Fs6MARKt9uJm7H6XkBznqprk1rO2Tj+KGHtEpM3YigK7
5Biohjl1Wql8HkrrkbAUB6af3OjWmYP1J4qmTHDIj3Ro7jHAmaCyzqAYwxdPnnu2
28dnOJ5mRyLMFfVNK15voCJkThftYBDEt73ui8oRyQfrrx3dE6GddkCWwyV3g3b7
M+rjxutZzWVNa8zgoLuqjw==
`protect END_PROTECTED
