`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Kwjr+rrtxpe4HZS108lSkSLImsUA19zn8I7f3dpg3qD2GV9mNAdz+x2tld/v5a8Y
Sc83F4lvRjmOPmSB2kyFChbQV5vOoH40/KdNLxQFZzZXI2XchbPepu6vu17mMWoI
eaDIuvYyBpilhs1Iim4wDp1gLsHNjiliYIyO3DGUz6xOECdHdI+2vWvQTJhFOs2J
6fH4ytQJbSXimO2ihT1c7pz9Q+1x1hPpUp1N/aqPBGE9nXh/vB0FtD6BU2KmaDnV
WGAhlxE3mK98D+XnZOpRSEb4EPbvKMCDK6duRar2AF4iOzpihOOmRXdP5ULnV4fJ
UewyLjA2UPLCYfdsmHYRCs7XutIOAYHQ3ql0oYeb2ehNqa/R2TTsaFTMt5IJp2Mg
EVDQJKnqWq6zeiKMNlGydciOfYagP3wDifJlQCrYq+gu3ja0JYdEDw4qigP6n2SS
vEBGpclCyues44hg8umShElJMsPDH75ivnB3DqEWFFPtcEM/+W7sFhQ04S6qkPpc
TkwPtZ6DyvriHlbXCvSghC6iWheCuqR+tdnEx5En2qXmPDjB7Q3GepUlps3epeA7
x14XSn1+MimmgVvmZPkGmB/Uj4btX1ytHPVf/37st6VDoUqCCeuvRW5xUmgBUoYh
hxPz0WF1bgtAZes8KsbbxSz8zQ4taWAAKX5MEFZxD2R/z41PuWI0UTuBm//coo1x
PutM1FYLh93L5QMgW2SFxw==
`protect END_PROTECTED
