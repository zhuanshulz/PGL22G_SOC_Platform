`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
86pfxoLsa+uBjZFDxbvSWB4VjDrC2hUIWWMTrnqlrNzIMzwcWFVqU7SA3hXfkBQl
itK6qHR5B/bOeHaBa5Tj5syhv4g2b3iQWXgfkstqWmFnmNdveycZWICZRomhtBUI
DaTTp8y+m2UWnwYd2YHc4t/qqYuBZPrKTRG+XmL38/BeSk9M+ql0NIs9K9Nljo7L
siimjw3t0ZU2olkgbsHKzVO6N3xfO9g35jsHkuW2p2xoQUrPjhUekwXZ7xq8AOid
NlX3v2v0edpctd5EXrHmyeCHKLjQ+XAlETVhjwBHam1RRJMJzkkunB6Pseq4v7cB
QLp8i1IxnJ202s/Zx4UG23lc6MJgOnCT3SUb+ZQaXOIXoXzRP8Bc/cO07A9MqypL
PIQJpNujanP8NwyCCUUhwg==
`protect END_PROTECTED
