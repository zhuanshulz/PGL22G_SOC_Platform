`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1L5UDDOeY1hFZuFHnojS8+q2ESFEcFZ5lqnr35+EzYI4FBXns2goNK9dt8exZNxw
RfZ/rGejunlykpmqdxBKc60EIYO//uohQ5witEhL3TztC5TZlfmxpHA4zsZW3qq8
pZJZ2mrwR1oYEiAvFY8kxiW4SEcMt7HCaTLjlA9OVb8T4MzPt0W1Mz2YH0NaUVFT
a7TpWgXU8Gtrg5UlpVbNL7Uu1MQV2Z83FnvLyEubGztSPIVPZqZU+TFv/aWTLCGy
f07YSqaVRFQ3ZwyIjt6d1noSdYeV2PEg77FRCeLaTMOPpn/Bio5h7ZrABRETcD0N
qr9RdUnBjjKi1ci1nTfTpSLE2xqrE07kI9Hg+4AS1M2M6kPCLY7J01lh/5MVg1x+
OElsRZcHwtOte2Ib2Udloc/G8w+vcKHFI1THDkBB4wCxd8tvfBcfpVlmY2uKr5Cv
HAZF495ielNcxmPeUW/+7HhIOm/397guMkWaosG7a9PAolGfhO31OxwxSQdU/Bpd
THiTqlIZH4uwhY1djf3DWr+FA+FFNq6HNGuvk4ZZ4/xntH4jGgiyNOohtJdlYpUe
J2YuXqWAShbzUAB5J/8unZT0VALXsNW7Q1SQTBQfd8+7/1OOp9QWA+qMW5J0Sy18
oIMfwP4AvgrmwncbvH3icxon5CZ2vZiQBs136tB9AB4Sc5xjbaPRLzQIJA3hhfS8
5klyds1Cg6A3olPM7bpSojArJ/2803Xw/unGpzoGf24KoRvU7OC7M9v9z0+QQKa3
bK8PFT/gZYP01XvIbCrqGa+NFVdnujvzzlP8+HgOqacTE2ojEfb4VbnJ0BPKQSy5
ojRu85wg0+1uEyhtOdV32cSHn4IGsoB1Lw1XZyRQik6uQEE+Pe1CHPzBsAgsyzoL
/rCKy8JqHu+Tvk6kEns2dEGNqXPpphJIClnnZsAEu4CgVT17Rnrfrqg6SCU2h1eM
L0Y5X1g4t3sYd2D5c1VUWBEa+rsMyLqTWi+yUni1GVXTI2BCFSGF7VMKMYAvD03a
12HjV1z2GSnwE9s4s7qlPA7Amw4j/up/n27JVrA0opSgEqEgWpRMKNY3x630q1w+
yfBp4k4k1BeCcLRovdk/FonDAqpdUtYRY8tqoHeakQ42gV1NRLu0sqQtGsMM4VQx
laMD26QRgyGPDhgwds/eXB5+s7O5XnskpzDeW30jVGKl7yLsPuJKDGkEImE9Hgeu
y01nKDYGCS7x16x7BlUzLMlO8r4WWSfHSyeCWxGsdDBvBZrAmc9Axhng2I7SIaem
9xFLeePMkzkI8pLiKIo9g/Nm0Y+6Vho6tI48ILT2d59wc9o34GgYHRKHHyGFa/hs
OJZjQJiOCweX2LHTJQG16PcMvyeF6ugDGx1XI3ucZszvcfshHNkZ6V1d0KCOQPxZ
4ODTVYpLeMXF3mQRJHXYGZEsDtKUtrgRqV6vQXqRDbKo/vG4u3rUxUPfysLqx1zx
vun88ve3ZmEckp1woJrstCoZOa24z8vniUI86QXqgqSkiT2vxRXkFQk+BKk9P6uh
0hdRN0tgKCv9JYJ+N6kpJjD/lkKbOqO6UKrZw6Cxz8THd6Mv5WqTdBHRppMgSfBh
sRoqD+bGziXKtsikY/7Ay4zY6W78UCPb6zMojLVX/qTznrJNkT1No0kj1Pq+zW2n
+AQamrGWabtW2KtmnuJscDLwPDK3ESLbJ2QbQalPpNQWcGroZbCpfPRm0RFjR0AP
oFYeML7L3aK7VC8iRSginw==
`protect END_PROTECTED
