`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p5WXbvxSZBA8Q2SHk0hU9LB8zrZEe1i4bWKr9BL46T7a9wPOkBDFpTW6XbmqxGxc
ystZsG6TwUsm/6jachy3Mgtz/HMcIitlJOdxOZJbOYOWuCMHeNRRXIN9CMiu9OSq
5495/dGYN69BPpBODBILseXZsKgpbNdtqh6QekzVep66bs+VQ0SJjTazBzrQbfri
9MZD2ZEwcg73rY6k6nHqrOfGXRUZYtaHxAgw3uJ5yU5XBi+uGUyhxP4BKs6AKZ+V
juFHB4vqqf+6gUfz9ZHBbqGHlWMZHs/FByWa9NfGtA9RUYlLz4T5rtK4PS7BOigj
9/OLL8NPk84E0bbA8B92yhxq7Xaiz9pvF44I/iC/aP/+Yy0RdTQKDwMxrEniod2v
xigKQYMExMKM/SOx8PuxUKfQQpQR0MhBvNGVdVpFLIU4xace0leYvpIz0ujwKQu+
eGdikkl1YP1ecasNSz98MQ4AayUoLK+dVWr9hhkLdbaIQKRveVhiTEy7BmbEOfPt
11Src97f28RswcXqKIpMmDNF9Q+LMm5p2P17fwxzCObImnG6LyvFRIt+d244+6vt
bLMcKstP6fqodGhvOHOvjWawwWo/rCdoJawTUbblitBEj4D66D157k8JoUjVvfPT
s6NYQBMFtkPZzb23eDsD2kjwpmLuOyqeDuJ7E+oku084/LoAMegZKd5bicAb9tFk
nedKlXl6NdbvpigRRc4AmG4pQfdElOZS9tS9uXqkQFQmqg9pIxuEkV8OKEKc2roX
qc1QK2vyHgU7UKfye4DXBW6h883peorsBhpLx5t8cPmR0mA410NA2yq50Tkmnia5
Z7IMjnQcMc9sAssGZonHm5JqgNEugcn8Beh/CcRrkFc=
`protect END_PROTECTED
