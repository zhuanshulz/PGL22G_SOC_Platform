`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AM54YmMvW2+Avz4iWb5M4xFFa0d1p00bXw2JrselScqrLrI3R434sw2F/AzJwaSI
mtXhn0YEqGDCTqELuhz1kjVN2tbLPVLCB8tpvW5CEV0hkLPFPPjbsJGDnFjJUmDE
bMolFh3KJ1gZMXhvZv7npWFw5HtKYhdR7ilt6CpzHqKsGIVnCA9EyxPI8jE1eDPJ
edf1mFECQ9XbGtWCzxNsKWXU/OcpNpienCE6sF3eWTgy4Kmn5gf7GYm9sbpi91Vj
g1YZmLvfmyQXNC15voPKChp3Y+/g1cvySI6gJ9IN/RuzMhS3JVZiM34DkZvvN45/
z/MmWUIzQQHTZMAeaDSTjGfeDiD/jNzjr6TFG8qkEhVvj32J4Kf7jKyDVwCiMdJg
tCNZSgbDFzeURIKg3avKT7qRqkmRVXePp5zWNjyxjKbjJh/SsdMf4wruTCJWT+Bw
eFQdAsa/Xx1d17ylkb60roPjJa3O7zGiLh05obBAvvHFu4Hk/2Kekpin4UDvxrjS
rJ3b6gau1fbGhgJZj6bTFhc/8YOWWCR8MfS48bYyE2lwOP//tZIf0VTlWfS3/OKK
YwrfqU6RN4PWM9+Afb/AqT/uzrOHk13gvLZGVgqDaTbn4IuvT/U0OxglDfA6mpD6
Ug9NMxNhhnkVBh7AT0CzHQ==
`protect END_PROTECTED
