`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DY9iGMw5Y+6h7VfmmvUJEsSt2w9afYggXg+TNImgRQRCWCoeVhITAgEPfRD1+fVb
8ce9UmsMG5sKvOKAWcrxbvULTwFH+7fPSjfcpeb7/fIH3jam5x/PHKDGgLH9ggae
ZqfGfMLiVLPNaBcquLJwjiIFLeEUUZS4CMSC/dgiJLEvFP+dSlQRUp029c+8EHbi
TDdYnkqG0oofZOdKrggPLkVfY/JmtFYpa7qJ7dPg/ZdP5TMWhdYjP8fOwwsXHbmL
rmtjYSLCBw4aK6cCBampOJyaSKXR54Wpj43bwdRg1TLQsHZjNff4YuARYawOtvFq
HlAC+XgihZL7sqLBHpYVoSvopmEoBgWuJqPis+UkwfAD+pNb0GxFEnRR++xDE9sF
BFgeJ5Okut7CPnCbqWMwCwfTTfa9v8xv1OmKDe4YSQI6hysHSnPYzPtMR2i0bxTa
1Y1XUxhoOt1qQVQcbEXCc6cScasB5yNGv+Y/ywv9SQf8KOH2XB0SMfPwypH2Wjqg
/CE+f6UpSUQzmmjyTna8xcb1ee5a8X6YmwxVq/PO/cW7iOEHaLcbe1oPwSeacLmp
bJ7Y2E61nIK0AvglDCtsiAtDTV4dBpLCc3Y36dryZShKsbJqXOvTwrxS0ERLpzGp
HNGYEpR+HW6MzOE5q8Xji38WuCuea0WfLAHBIlXdjETLFmrNJmVL6l8dAt9TIQcs
VjTS7+SeByHY5Mong22BfLNQVRStDF+HIExk+oAuSk3gakaMfxcsnLlcpX4BzYp4
SzL2xZVqDixwBByZQsQb/Xt5ou7LtU6M7mOC4rl66NE01OuaIleO3Et+8E06RJT0
ktC7gsumvzFAZL+sLxqHW1eDdltRu2sNZrPwjPLPkqpVVXB+X4/mdYoUYUK450i9
W7A0p2i+FbqymWdpN4V5lTxvbuFCDUk7F3Fn4S8Ujt38PXLvt7cH5d6Qe7N4ThAo
+6RQ9sqqkKIfymLSDnDyn7YVmYG4xkPwxTAUoZStSJAS/+QpOo7eXwEfzApOcDxE
e0rAFkZDbTvY7PPr1o5U6FBvUtahn354d/74OzwFgOpQ2Xh/LRTLQTZxKcL9aHUc
B0RSgmECF83N1S9cMi+C5HuLE6uP7MnJQAqBJbGGhYj65RcsvczqvEPdsxZozlS2
ciVwretpzeUID1KW1QvU2BunC+ign+DriIVDLbprgPVlC7JvPuHgtO+5ja5TEYeB
uv5VcTbrQw6msDgYfVJ6Uya40dzGJgnuUS8O7OZNfEOtfFXrHJ1fM5ZCH1bQIpFK
xvQmUDJA5F2kkSOvYWCQbiaapBxGlRCrbUmeN2NKceO7vgRdjPhNQHG4sO17ov69
ooqmfCduvLZRpm2cSJgdEK+fSS0K8eqLiejnAjygr+luv9vuWYNNgccUfL9sjlyq
KDKXp8kzz8cbUdjvoLuHr/66L4cj+PC1IhURgwYOoLtXddOUQgcHOjSwTmSod6Cm
K580wi7+cxB1NXw322B6qqW0DEOQY1W9sxqtuoKJw6XtnhYHkwPByowwaLRo7iex
i2ttynjpNcQk6ewhQsMWszPf0g3SbirvFeXKHgI88UuHuSJeXH/deHfngdMUPu7B
fEpTNeJtYiw3NosS6cG3aQi1I97y83kIkZ+zoJmskvJ2iKXH9LvFAEzcSsf9MYoM
yQMjX7gvEErWsd0Vw7d1CwxnVCiUkCtVqFpii5xq7xyZzal7h69X1edUZw3KrzsE
EGtun7LkBv9mWzQsQlo5eWS8btDnnHAy6GpXWYc7lf8HxpTRaf38lFmFMxxAtfzp
NsfyCIqm2WrU7ROVj1paPG2j5D91UNJ8F3vxZqM0t2H2QfvoshTySEcUDc56oxLN
ylYua2cLQQ8EDrHA53/ZuyMVODfHLXsZ2rVDQHfrGcEwxkRWltf3QtK3b4WQmm+z
IbBkeZ1wl9vQIYIeoCmpBsbtltbMp43QoJmXFVTmqVvgv5DHLq243JtogbBxIvEQ
cK/zh7pFjx3+BlKomSLOqfKaqOGvrVSc4BWHta41KlWP3BMsEsO74M75aRqOeGrk
GT5poRmMgnPcKcW6QRYpOHIxeyGucij7xcNGrUJ4tE/MHspHpTGz3uL2tYm73gYm
4Kdetiy4qu7ur2H66ZHWv2/Ik/p5To4XGiBGwkcrWol+2Za3icbi1g5BB4m7x+uJ
WsaFek6IChw4t55ZgJl8SAH8On6Hw+Jpz1tIESw7E1Iy2qhSb9zDOgViT7F0eN36
tDjPemUWdxOYpn6Adl4elMOylguNxDqFXhNcM7anXasf41I0LrIHGw3qfNUgk2ab
KAr7AL8AW86TRX20uMY0kFCK5n+6PdKN6TEssxxaJJzBsSeoSpxBEwcigtcU3DWr
QbJ0uNv2ABAUiG1E0pCCFNUCB1IvoQUJgla2/nqDHz/UL/Hvk7zhxoaiU1dFZqzt
T7h4zNs8Ho9NtO44jGDQOXtHI11uCxtdJ+zW93kPZqp9KxTmXxXktSoA9olWK2nH
moVzb2RFiMOqKVAVaUlBG6gMGLRpp2XkLJBqAEgDTGTfaw4CUwfhSiPrRWC7wmwF
MgQtLRFwX5tUd0Mo58XoveAuegHzaNijLU8EnJWFHzMOog7ry9dBgYNW5oTKoTG4
dNCZjGpd6hB3y1Cw9oHKOo/areNnC1Kx3nytlz7+C4KVEh3F+rQPEe+NyCyn4Iru
JFTMAwB52DLL5AXwLf7G6YL0O8eWZNhni4c4f7Xs1RdLFz2YW49as+/60/HvmS+r
lPf8WZEtiFKTI7NkcNemYxP72of9q4LvdHCHqvqcXjbtC/n1iwtg2lnm6REoxJtg
bgm3aaNlIQ2Np+r0KLkvs4XaQtbFO8Mknj/qhD+0YQc3lMXukKqVYgbgAi7ZJZBh
fP9zx/VH67ArEvLs2T1jK6G40+9oLvrHXuT/vwR/8ImoSole6rkiK23Y3cLNxqkM
YmR94D9oWSkkvGxUD+5bjfKDMtTnL9TQ6IgiTBQ4sGn5E/5GdvIFUMSn7YEu20Qu
903LQXjjqsTfOBoy80uId/7gw/8Tji3VwRRiEteIlBNud9Ec53tz7CROBVwJRQpE
jr0Kr/44nYpjFuDOs3LccB/v8dYp3Esdwm7KgOpe3BBXqsFSXbaGALu2yg5XkGAv
zwGE8CL/RWwaRbIoGgWIMK5EDTQTGQTV0K8+CsgjgcV6eqfdTH2LZc4FB1544/Qu
wgWYAdVsPbwLIxSbJ7M/wUPS/dqnMxC3nQjHaBmzx2zE8n8q8MAm3j55kTU9C2lT
gJa5DexMncJYkXcDvVeHTJIpQ738xvo3bzLYdD5b09loIWVS7iqICfKd/wZwGicL
xFVsiExc6Bq1h5kF0bZK1gIvM0hEBjFFdn4auaAW5NyRJYOtW/Rq+NjNm8KxvNSE
dUzCexpUOTpGvklH8vlVMu9VWgVrM79cR5rObhPRZ7QZoyh9H1IhjCU37F/6InmF
gsZhn8BqcgcVlfPJNJ0zNpVo6LBh5pdLg07K89JbZsh32L5yLjY0FMIuMlVFK3o8
YUFY4B/RWaLcjfLttP12tbYX1HU2QBLGq15J8q3iygD2cH7M/a7iviT0FDhdR3G3
Gz1GBQNkP1jlds0M4VDiHV3y2NGZsB1UUQJQP+Z07A2uLg7X+NsCD58uCSsIveVt
DzhPVNNO1UnxHer0BmdGJLzdU4FXjz8GSKYwLArvF9VbM1U0cvO0Q7a8k1pcFPyd
ARYNa2ewJBFc2CjQC3mxINVB0CIa1MM1aJH7pfNrwoY+VPdxPP5B3Hu90XUSLvdq
RfATmhiYVpc4rCwu8LIfRSUd8GjRHQOvBiqr3GB0NyfZFB02OcwjD4EWy2vyVS0j
7lZDoOmAOVqiJzI2IdOtjn09ntFg0rz5MQFypiIkRM+0oLv7MKZso9Lze2D8E00F
g984mcVgieRNRwP4UJ4TrzXSSFFcM4e6yfix47eaFN3tRGouQV6fbD+HEiSrYffq
pVajGyomjlgwlCxtCmdROicekuakwvR5CVKHx/F/wM/KlmgoqJ7lKZpMx9qhVt2j
d6MBfWu5B9Gh/QjTY05CHXhLM8YLJrkpOQRMX7ivjbTna3hMN5NmWZyz+t77w+UB
Rhah3NB/5KjXtvciiiZdjgWnmeffAy7cily2qFoHvQAcBrk4atFjQF81kqMSt7TH
jKfke0Gc00hECAiBZKz+HCdoRzJrpWa27sWoIIDnLm0tFzyJx+mnRvfdG56yA/13
444uOH3NSsK9XYJ1Lm7Tqet4BT/1b5sqFDdd/xxaUhWK6cUZwwWeKd+eIdVNDzUK
YL00DKO6xgE4jeveSrHGx/X9w0eMiaz/NUIyOKyKClJVYBkW3KhILCRcaQou3krE
LKeCEOmGduo6+/WEB96toubgtzSROhADhALNjc10yHJapYfsSyrSVWTDZ21zv/2c
PBqX9lo2d7ep98y6aEYqnggO/QFVLjukPHR9DLmIhRlOlpzE/SxZzdw94+pMfUjx
yHSSIalS7smvtkSVzEvZU3+dk9EG3R3YcbmDGIY8Vu6IvfdLaDUB4DzG2iGZ//+6
/3RwK2iGdNqvw207Ftc1xYBykE2JCUQyj9q9t+RtyN1LQToSzi8wKp2GIr59uH/2
pSAeNd2z/wCzzliM0J3iZizT05LRxKBZKn0tRwUuZhjv59HGxR/jpJZW4qUtBXaC
es7wd+Y1VcIvgZrxw652cTktWxy8jBKNAJGVOMzP2Scq3Z7L1UInXlV9qpcdDsSy
namSTiyceRpGyanbX4xrf99xfUdyK6aWvO3MDkuAUoVCv9XXa9wcUJ34eDkis1r1
kajPu+MgoO7mwesnyOJTbGrCrYZsLYE7maeCb1+dlT1qx74cZembVG0X07RlAXZa
ED5NuE4k9ZeokbpKXieFmMOyRPVAIjI1h1MMM72+pd31jzbK7DKh879WsBdPJTIA
6ayzzvnN00TIKr98dKn9Kv1cdgJImRMHdXJspDSNtiY3BMhO+MxOwRsiVQS8Nubc
IRVLAg5LHpPDxDVIScUa6Zc9r0YsY8EqJzslgiYFd0qZu0Fv8MohI6n3Is7wtyEV
L0Ij5N7q6Qp19WO5mgHU3W725c0bSzWICEo/3ZHHTT5iTKeMTtqV8Z7zZc6Ab5Fs
DYXQec7Ke7tMTQo/j3OdKLCPFGk9Dz5DKJl5nvNnEQdOwmOm/qw/XxEpeENzJq/2
Fz6tylgOAMQXffahGhTr+s0ZENJgFYKmEKA61ApwaY8QY1hbbl718MECqye8hH7M
4ooQsimy+CSqtkNibRFM9+LngsSt6hV8ZL9MuM76pidnTmfZcOwudXLJ/AwExc79
yXlhqmg02ZO9aEMVHTH60U1SCWevsuFraQjJraqHSJyLDuXzOhXJQD8+b5ertF8/
QdVfr+/O37oe4A/IHwkmG19y4VDAn3J1AM9QA+7LhqvM5udfX5KrnaKQX0w23ZCT
ojdb7gZPNjYwD2MvpoUBFVeOLMuH5q98XnQrQU0hSnUSJO4ZQV6vWVULcmufbQZb
BR6M0kYnpvSz1czLiKuze6eLxKD1Ar3Hd0LKteu5ovMq8tVZFByPcuTmqNktOlSJ
vurqSv7CdxkCNkFxVrkeliVHvw/5n1VOg8wjPhgTgjwBYcGUU682SEXvg+nb138B
zt75Toq2drPc5NH2CF460LfZWnBCdVErO0Udn/KVco/UXUC0m5CrhxHRzFDpTzZq
2ombXXrrtx3IvO10KwuS1bsPH202zURkN05ZkPXf5BwwhNCAmRl7HVBytj4i7m4Q
qfT9+ZpbuL5Vf2vQIKN3hQEXC6j7ckuB5JhSTwsylUk3XlHQW5b3/EJTMyREwK99
R7AVRo/7dMYZBNM7tsjeJ/Vm1woLckyb89N34ObEl5LCYnEtKHqpMD7q46xV7Z4j
w9f5PppXzkylr+J/L8fbpDybk7DDranmV2gq74Mkes9XUm9iNPDQO5XCqaIG5ifw
UlBtJUuEm3xkAKEgC5gHs9xET311wDduv/fMdx2SOniwTcUwwBrlQrbbZ5POUn7s
fWxp5YJS/2fpmEUqaBbQc/ZUzOLUqxXAeiq0K3XlIwg3GhoZFtm6IZbKirGFymwB
Y+uJpysqVf3H40rgJT9Lqq4MyYZf72asoLQnydPaLoaVLPKo+QBPs2/s9SljDN7b
Ay3Sd/3KfyR5EgrAmcCoj4lRJdMpNQ7LdzsO3VrEueXpuFQICjY2TmxWix+yU4H5
HnpXoc0QJW47+0iM4gIkza9NEkoJ8GI+UPUDhFjHUMkbM6IG9gdIoQFHmyQKgSKW
ZECvxBUPuP0+aGFlrlMvlJS7u5X3QI5yA6USnJ2QimowgK8o24N947KCc/g6rHvf
AQMWkV571hAJ9zMabn/ueJEw9cSi5jJRS2QUnKbr0W9ZGqEZORaV0RNPmhZoSJGz
XqWaQgsnGJvP1GQd17FqkWqBe0WF1ELvk9KJ7pVuHayKni46HlRMjoYejXVEM/H5
ttu3uZP9B6rMDfoJjFKI2D8c8ffBrg70do14njVBWR3pVZ1LNGi9woI5UvSudppk
Yq43EzQLBXXjlmEN4+jpYWmM4YrFhg010zqvS3O9qvt0+yPbLkSJzKOc7G1RzOKU
g9sExMRNjPTqxVSEgMOKWhMZizSo8oNJmGLE73CC3zXr5/JTIyw1exI3xciP0n25
U4oy2siBGoe4LBuLRPnjshpq7FHNFviVdz66hAvg7jrsqy7IXCQiUMg5dbUGJnsy
Nw7Sk+AdoGtSOK//0RQKyX3+0NgWvhFFp3C2SY73Btp76Wtvk4kGrUGUmMYpFWSw
1H4IU0mwXlQ9fyzXeJSdVgv2szZbfyLTxF6tvEf3xtlZ7xsdToTGiASOnJWQaze0
o67brTWF0L/Cndm2sBArBiHyofiG0nTIeY35KprXd0ppA+9TIwtuKCZoUDGE3PIY
WSoSQtAEeCkvW9BU7jIhrJ6KgkR5C/6dDeDNn0DtpSCAT8TbKspQXNSsYOW7oSZy
xD8sb6ynfH6xCu3syjgUwUDZLnQbBjhdRsU3VDONoaNWTTPa6Txu0TamvQAaWZ//
Vbjfny3Ja37Qt8KR7nZJ9OtEg1F5yNBZ4idD/gCAnpt/gc1yGRfjqoCR4jC6b2m5
LqsUpoDNpWBPIoioYuvXizYmXNvc6wj4r0+nuxjTwVcymuU9UbNbHdzCnVA69PAf
yN4WMlWlQ2BqNTlOZmtwyXSuC3V0CN/V4TgK4kuZZphEsnzgIoxTe93zICMyQoTt
Ptna+cxk8vL+eMMWcfI9Qcl429qvkupuih37Vhn2GAa3n19myL+UX/s9k2kyu/l9
LyxKmnJR0SfAbbYWgtAcFsnNMdXQKNVDu8bOcNylPgUe9Wc5ro/ydOkZQgb4hcGj
27KFAA4R5RMd8Oseu5AbqZLHUlWRfu3iOwXzLgfR8oBRjCIvcBuHod8EJ9pj86np
YbSUK3C3LWej/c3ma3nMQaqeRNymkebenwxgY31RVJwy7gvto8R9QMKL7rfVv8wq
g18ob01/VVgV5UGSoOrprRxURbOK32R2P+eYXRBuXj+9KxR/66BL5NhFmZRPeFGr
pFt5oLEms1e63+xkNJZK46m5nu63drwrpcBvyj9UTEdE/hOJdNJi1sxWtbcictmN
cudfwVq8dQB53JGGf0+e6JTAVPH9qYI89l56QqHokpEFZnUJ3IBccwFh6jGIbLRJ
BmTXQ3tAtpH4H+S8Um3AN3j5loLhwS8SqVXEW4rYvHxm0cc57mKojK7fsySQEMIT
060DnGHCQvzHPMDlMt9DPA==
`protect END_PROTECTED
