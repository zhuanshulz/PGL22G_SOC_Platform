`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VaF/iP/tafbyjNbDqv5H4iGY+wRZmlfthei19PRk6bkdppRMplotu+aMTlj1l7EH
CvcwLIY0OkogPr7usfcFOJRQJViqEQDG+SBVIWBBpGiERppVK0Joy8GPe6Q4LTeQ
r7eyZ04LHhZb76R4VUxPnvTjr/yhsJCmEb3B/Dl2a56VZbshp2FDO8SWlD9/AIeE
CeR5wDHyGVr/JQmqAj+wgspN/hxYvTfyR5QImy/6v7C8YzsvzDlEC1ESJrJh1XO9
uVTCGtiDbAWDb1yn/NH9tgKjTNP4/xE6hrsA3f2mXl29eVkCgINq1yh/gIn8NQTb
b0n4gSrvRFSTDa2wY0vXSE34dqPrDJiByvmLvMX3TVv+TiOY8/wu5A+NiXbrEG3L
ckt5XGEPDT2wyTXyrgecs5kn4Ksm0fLOJ0sAg6SlDd19QxUzHP303KUkqf/kl/hi
tHX3btj9ziVeVS+W8l/rqRYgEPB6iWTdiCGeELe9cMd9wfCSpS/chyVuoI8Domxb
2QzFgntxvDYoKy6ksfXHIhILgy1hByj/I578/H2tl0RJeJwtt/Lm35AWO8KXhOaZ
+ctFkekM8fzsjs2n5rtehjZz953dSGMarnpesEKf7WMRC7l8LH7nfVdHi5Ava/4U
fhaDgJbe7kA3+yvtft6MMUylNHz0AeBlt5Hnt25KYoDcZqGdfqCXPpp1pLqpaVDk
0FSC/yfHBaGMN9oDZXmmd4Xb0ip4fLmb8SRZ0JqI/bUOghc1LGZrhZxhOogdMJdy
/yb4F2iKzSxPDgU64EVR++o1J5aQmCSfiCrh0yzoKZ2918aNrFmyaXEH8WXw2fCS
KHot0VzeoKt5qDXqYn6BB3Eq0Yeergo4ipkJ0K71mfT4Ll+4i7lJLpK1YHfyrvcI
G/AGSV+la4XXzENSbqGnkmGTNGuYOnudgtezBSrUs+yqSZZGFJHRZQtJjeGv/K9Q
4IbMnUMpyGUa5t6sZKGjgipFaUBTYUwwFSUAtIflJWc7RNTL6EUo0vPU0n1YOldh
rl66zEJUSr48yr8YpNxyLf/Pt0nBiQ5gP+bVuSqUc8PjGz/O6s1ZowpFkbj+uuJY
IR2vChdrnxVwEG8Dz/w1KIZ0LAK1jNskqdlvYsZSnZR89oq8pPtUvxjYwfIrJgC2
POMm97//HRbrnCFUatfcluk2cLLptE4jkWvv1N/kAF1UdkkXsqj2Dov8oQG39N7B
C5gIC/RpZEw2b1JEssvHQ/VRrvUH/+sTbJ1aWtedUSN048qo5woEved+UjEWBHdu
O5Zl/Wlb+S2ienwxiJgOzfe2LLD7UCIwCbi/lN7YZBqwWkolEGhUcgHA2kdRf7jq
/00figPLjbE0LbegskdA9uOzdTNQ8EEIe7oE/iw2rvT/OIG2uuoMeNoqrtWDGD7j
tJIQwkfElu/ejhMNqIjt0bfyt6AZJqHsiyvrpVc/Us+Ae/RwwcYJAMZn9jfwHDrc
vB6sTPCmqUPkv/cDlGuAOgDXQECwK+QIDyi9GbGkFS6JjpemrrkhdNV1GFKP7C68
eUYXRlgNaAuF4qQVsUUPlLsDybCXbllJlk53VFg5utvXYnTVe2tpnxTnGbpFAink
mAJw6g1EDCo+sQI5Zc3KoDqrvuB3uoiDTuuw0UuecKwFGlAh2I6qjprEKvF+rS9t
hpUArcNrNNv+qhmpIBvZe992NkS9P85qjeKJtRKfhvfvzP26Nuc403HjlU24I6Fh
CUpchQet5BOjmLacoUg9Quj/NH1e21fxMjU0Vs2Oo+5kgWpf98r4r7eyxyvKeJ5C
VG+yeKMCVWz6XfH/bdA+Qi3el8o68uXdAYW706HLZlgXD7igxMcA1lvQ2W0EiWrD
f/1Gf+Bij+zN0wgSDOWhWYnyLP/ijAwvIv7b4QJ2JvF2XCy1/sxB69rzpwu8romH
3rx++JQg8/u/L+Nv/GodfyiYV9qTHmO/4O0C7ywtjjiLsMUaIVT2Ws2qzy/+jrjF
EdakOIao+iP1FjQ8tSVJ28KyywXZAtEprJ+9Swy1j4bWiC4kf9aiu2iFafQ72hHy
sd26wHjMQlgxa/zUA0kIBkATaXZ4/53zq12UzX02VfmuQk5ijgGC07G+Bq1cViCl
MCkh14wAKmhASu/dtvUzK9WXocJ1/SsbiBo3qlgNDdfAkV17KdUWo+G22iXTLKs7
1TG7X+FlclilKtQDONChsc7YCUTpBrGPpIoKiyW/tgDZex5IyaK5pz+j6EBnqS4j
Sd/AkfGu+7jIgEUc1nS5ZjFkOXLQpKHrTyE4EEa992FpMiLURKRyJ2Gtiz9YmAY6
IXXzwWBQ6ghe7mwnUdb5HiDSLjXn798IbzJmwHkQkBfaGqcXI7zsxortwzWzzmzj
oh/7GfsyIa5M4rp/1BhewRTZMTK17GVikLhedrdzCS3Uzg+isgURYTno8mPFvdh3
OnvKNL/U8KMy+kriyzlg+PlZ3eBJZJRgZhFpKVLA+VTC45GXgl2RSKTRCq6iCUWa
J7m5Kof71aGSu6vuqRn9HI6Wmeg6vNR2nwqulOUb0GYYi7/E2SkIqmNb9uiCBFot
alMAhniBAKH6JWDEDf8NnvuzW34OcbuXPI5SckVynGCvnPbbUDB97aZwqKS1gLVG
8/wNeQ4Lm9FMQ3dVXL5qQlsoHq+SskFCu5CwrvvvjCBSlVXjuStJRuIx7b9MXAcK
3q1eNrQBP592Mihf+nRJXeAnnSrNUANwenqlaefrWl9sUxlKunjUPGi/9HJ0gvmm
wckhpzcAOGdqZlCTxmRLHi3HCi6Zk3a2888wCADUsij2wcKbiZQvcNTaqErvtBgI
8FDLoTh/LHyG/HfGz3oyDWGqdNdWq27ESk3axV+yVHQwbJltwteY8ICAcdERzGol
AF5GMljq1VhSYos2ySh75YXoIO0qdjNg9as6YbgMlcCDE6TbNd9hoE4GO3hKJLN/
2LCrKqbEFYMUb4eBcRAmku9S8HtMWMaWeK3L3Nop+Y15hhEPp8ZkX07YTDTA4y95
eiMmh6uw0ZoVIvZxtAw3PpvRAJwB6jhlxJc/zFNNnAOYFEYDEGntI1r32apqNXPi
Jf7YRHifnOcMKzLBpesrdqXufNT7I/89WQ3LfB0q6eF9eXM82bpcIqXqAY5SvxQ0
iYvFSmVML0WL9su/4KEP+vcl8uqIYICd7X32fHNPtttLyuowSDbN09+9PwC43YRH
N0CP/N9HBiLEpJMrXmCEypGfQlPTv+3Z40bZghPc3hz73zwDCxs4oUkYm+jCoo2c
91d+jxoKC9na2eqdkDgVqzA6LZR4t+Gp+9+aRxkYhKgejewhCbYFU5rQrGb7SpA4
Iu23U7orugOZEZ5q9hyF2A44kvKIMp0KnjXgtq/SKdbiI3Ff2T6BJD6JHp2pJoVd
grJRY0/BRSfpFjGb63d2it378t5l5pwcs4difaPh9bS83Sm6fQ4IRjnBZJiX5p+P
ajgELVVpxQuTAZn0EOtMyrNP+KeJKdtfE7diMroAuNzEyh1ELAZBW9PmyugH6I37
9i10ktvn+8fVd+HRDmNf3eI7IJA7GbLUgmakGa9oEe06zVpnMCLMjXD/rbGmwiRn
pZ/EiXvCC5N999I4ax8AgW4DbS4wIGwpxip/7F8MZhZfHo/C2vtMh6xSNIQkFV2Y
/tspa+knR/yohd3JGrGUP2YPdi1wiN1NoJeI2c4YBpTx/CQFvc3YQ675vWkMez19
ZVwwxw53RF/GccvNTt18WBIW0X+vT4OiSC8xJQAZaHuBDi1cppc/BOxftybVvGSJ
kNQUhjNoOgq/4mytaRV42fylyjtQAHCCUFgp2FibphZZ3jNRpQmwSlRwXOl4WYVT
mW1aqHXJY9wK7F+t1BxFzTDPsz+dtC+jSDAsXfJwAdz0B7v9s3e707Bd0OqpkHgN
Nexzf4CVdAP20YYNAzdQNLSY+YXgG0eIBWyfLkqhKQyRFcUMIeHZY5kqFMWhRWWk
Yk2sSLzv6Zr8xR8z33ZiyV+01DTpSiFLgpwvh8zzVyqzR7ZYaKssrce9os9pi0Kg
Ote9dij1LX9QUUqXxJCwowIlP/0ZP07m4+8SVGEefAM=
`protect END_PROTECTED
