`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G5Aqd9mzbW156/msbDavxqY8eFn879WNxnFUnJMcSUjYy2AHfs6gZBXU6Dtt8YhC
1XxSHGUCsCWLCgDYynRBKG6x6Z+SEwDca5eVCPsDIUzZ4/oJYCs/RGcyxhXiRE+q
Y4EDtQ/198J55yr5rW19u9RiKBsQPDhaVCBK3VupqQ+eenQE9JTrbWF/t04k2GUl
a7tpUHN8ERQc6+WV/fn5iPStsuLIu/FwmLerr5DM24B2JUCnNL+7Mkx/xHAM03WS
rZFNoyjDVE0eYzBsE5TdCap+ZQIz7Hp//it3pCSoa3R5eew3jOHWGkJhfeVwMdnG
9A1NxeRGnqsdLewi+BSBXBkdV5DiudT89cizDMQB2DXh6ekOT/1S3H93VGU3juAV
Af4fAFZeemyRwjacqonIY4HsUhPu4RaQ3PKrP0kzkA4=
`protect END_PROTECTED
