`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3tcxjxWiAo24kqUixA+4xTWtgfxYvrNB7/I6yC8Qg9VhW5rRh6AA9BPgNvpdH1DJ
EGxgYCauryVlt+7YX3ynFW0raVxAK5GvwqMMKTUYTNHVGEqIkEL9bk1CCHxzYH77
veiUjM0l2cTiR7TYpC40XH5c11r0qyDeXDSQ4ySKUQqC381mAZSQAbVf90sdjlZN
P5TI9LNzABd//DTy0fleVnKAG45u5n+ulxxWUUzRKhJf+XpHhM/d6aMXwz+2I3yV
GrmoDE85GO0HeWWiqvRknFz9Mlj0kbRLZQs+M/GbAbtrM1+mFQBFiMjy46rszn6c
VP08Ood1jT7qEMtqFIcDqg==
`protect END_PROTECTED
