`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oXs2irZv/p4xB61h0ubeXKLnxrztWsey4E4VWWvZAV5DLuUEpyCHt837z/ZxddtY
WzYD3hyzOINvbQ1CjtBBaHO0DOZVatiifOSQmT7D63RTcNxJ4AFudfoHvu9m9xMS
OqyfvlkPyCthba6ko/zM1ScghAXS+Yo6cIyaDaTkdM9eKqVTfBCT8z0B8GGRWsfd
3KUYiZF5oHmcIx735bnWiyNL5mkYV7nbb9SAXVFpzieT6k+YsJ385yxzKedtOjUP
N+uQSpCdevBjkoKGjKZvIi/GM7y0Om3ZCCM2qpjVcItwmSlWKQJKEEoWH5l5dX8A
6p+3JDEjylKCFjskW1aeVwydof/+tlI7cI6B+sM3O+/Cu71masR4VoJtrPEjnFyC
ZCfdpvbooE775iofyox0tSysCYfkeXQM18mZu3wmQL+gpU44at44kj4nhw8EAlxQ
aJGJZMRbOQSrQuxQAkCFsUVGNPRZ+7cjkLEsO2f+TsXzmwmEj/nA7Wrav7r/CN95
0LlpZ5VexUdaYR2JHs4F69C6BaQ5EdhSDPx/Rgq2+fFdyJwJesTSyhuqGfJlTpA5
tLmBmb4Z7lbT8a47RVSmgOowLYSb3YnCkmPVpQ20wrJs+MEAyFW+g802lsq/thxm
lVOqMafgWeMZvyiSYG54kxLUWF6qua1/uTQpRgKXVPZ7D592d7hwHdhEKmOqwG8O
Ncq22jgH26lSfxwzBK6uoIL2HJt71HITJvprySu/90zja+CzjYMm0m/FnQeJt3Nb
n5Ogjri3DLOgorD3rT95bqYqK9NapN5MQhHT/Fpqd6XLg7NtzJ1BBDIt0ribfhvn
7ixc33l2uq43/muTDDL8G4f9RHjxOwHyy7I0Rw/+NQa1w5ge9IEoSTXC7zRHLDBr
qWKg48hulhE3ly0TSjK5/OAUnkWHxMREVB/p//ViF9Q+3xjwxRFoS97ipyRJul0y
z7QLKZTwW+kg2qt8xSYJap47BsD+OBeXV7pUXuck7djMhVsNmhjbGRDnGKUvFfue
LqPvfUA7TYlWwLYep0N7YiUMK+Ia+bprnJ4nl+/oo4FA/mIgLXrXd4MmI/DYqBs8
rpXVv2KbhaZkCXoJbp1neME6qokifth3TvaNTHzDJeejjjE420b5SWWuRuDG3vhP
JbcCHUGYrMruRgCqC5WCSrqhsyDxCVW3VQZJNPTPGe0oLB8bgvTlUPD0ZTzCkI1V
l82jTLaucEX6uoWjT1Xj38MyWV5IrVlunThvrHXKC+S5ukzs5NCxgqWLmtNyksWU
u2k4MLh9chvwml0elRqiMNKEocAgOA9OYO3ePAUOKh2P3KrTot1oXN7PLsEO+BXD
++6zIj0gWwXfgacKegGEnO2aOmRDAs71OhbTNTlH0Kx1gPqocXSckJ2xGy+0lJAR
HqnCo5cW+SuV2/N+amCQWcZrg+TQqdg0eQKyxqS8xcnxFFl6Fsx0nN79P9eeb6uD
YkoH0OoJQWdmYZQm4KTFj41kkoMLY37SzmVlJXF4/O1TX6UAGBvYfZ+bbJiTpWCn
sAIieNU8awa+1RZLtK2MYmzXNFbdl9JroQtjc7hyEu9HLvNePb7vdfVmbmIg55Oe
ei3kl5rXcWWNXWYk5BYV62A9AxUhakt2OcCqLwj0V3lnTo/W6wRsvH+5si1i9xzQ
4RGCg/Y4JMp6JRpzBvB4WZMTAIvcj1Ef1HddiQ6vdtj/7qIORWIbjC7RhhmgZK7v
l0rtb68LYNrl8RSeDweo5PMog14diH36RaLEfoe4XITiTXvyHoxCAQLahv4/aqG0
QwcMdcFeNvJpuNna58R3H4sAorUrj9suPGCgV9JChLYRK2UFrjb4Ada//zu/3ktW
6v8ee73NMnT8kAtdDcSje4hyV5wuXZtnw1wZvyxPgHfxSEvpH1eg3velI+oCqrCv
ENgzUfneyJscd0fp93lF2dKoRcftSBX1h0uDSA/kit3F8PrR9Se/PmNj1F3RtOMM
QdiwwQR4lE7vlbEOK9yku+xYnNNhJEPrlOixBeNSp+4YUaurOLpj6jpE+8kyTjjH
ayb5ADyq+OIqNXFv6dMWZxwZ6U1NdAnI1JRSoC3RXf/FoKb1ITyMvgyEgYEM71GA
9ZqW5+fdNunJi6VHe2GLgvfhjMtmOEzgTs6lxtSr35s9NoJVBmZGO0csfHbxQnE+
mC06Q9tBuqStjnmrSBY9QlpORdQGd/ikfK8VL4U2xpGIcspPO3U8RWPSTHT8Bi+y
czzqQvk7IbGtYCPKqK7tZhHcK4s3VbqZXelyYWG6sB20EG4oULBf0E5n1xg9g1L0
Hv0FYozlZyMINhJKzrPLogMJfq1S0iGFhJIJfBSFrJDAuPIblm84QOvPRoO4O4CB
a+iL5bkv31PuayaZ2N8Z233oUhjdI51FBa1SuawiDUY=
`protect END_PROTECTED
