`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YxpwLqBT8fbo5KPBZpuoCpEHVS3LHJb6+9WQl+M+nBsqWJavJ+DCEASdTO0cniwF
dYJkZTk8XFQ8db/ByPL6F3bm6cn5e2x7m4OMXqScdAptlgRpz3kYhiLdfgZlqDsZ
yyY9aGXMP+wJVNghULxELzmeN1EGrDxihzYIgf1GVMosVDiPfaOkGYfu6t9M5LkF
tzZz2XUc2HG2Tp0fNNzQ4EU/nYtLfQbXOmWIC9elUQhaRby8kHII513inw+RLsKH
Bq4WH8BQ9sO81ShX2qZmwQ==
`protect END_PROTECTED
