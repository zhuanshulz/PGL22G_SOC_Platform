`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6qECz0mQkCxaaquLRqTkGV1yFzxW5jwRR44KkLD4fvPD/B9Eqg58ObVyjatVlBS9
E4oiw+ul/eOQtaYf2sPrZvSrwAA7VOm1ZnGQAS5y9bSpbMelSeMt39X7cyyhWYSG
QObZgrKpXz5PBOW0Hv2oSdfszYCh2fjZu75fajfs/pIvLq7yD/e+V6Ux7m9jcTAR
kICC+u/mjldPgWkfpUOMs4Z7cXZDuU5sHVI9QlLPVaKVx8e1Hoe3Nbfx8ouM2XEx
OcSNXrVHTCe/JkRE0xvbKokM6Z48d0N7ERRIEvR4gm8xenDfaCBqdclak5tvULqx
J2yiWqUUucG22IUPw9qopeVCWTP4SU7aWEMnjUK12+CeDLNvrkTicdCcYGn0yu4Z
MksZVQ1FcbKEIHjkKTPAcsOuSdsdommIz0N0d7NU08JBU7rZvPRyaQsqGxbBMKJY
1xdGZ5V7tvOWSpyQATNGocobYx3GPeCNWy+c2Ca6XNrJpQxln4L6grNbWvo3sPhT
CLiLukK1G3iGTht5lE5ok1c+TejOEMPHT5Yf8o8MUc9ztPX5g1ihHNnzhmcDjZE5
6EEX2GCBQLqBSqgq5GvfjRkupPij1KJBXs0t4zeuo9Er1KV7mhdvOpZ82xNGS2Wh
c14kw338JHQTGd0OjAa2sR3vmuYgaEeTxG+zmK6OgVpw46qQrRe2QMtskzXwfarj
DB5e4+Eyz/yElsALgQAhhsWRPsMHzoL5P1TvYLm2SwbTYCd+1R7WUhghVoZ1Mk63
J7Mh+ACAIHxiv5D2lnkoIw==
`protect END_PROTECTED
