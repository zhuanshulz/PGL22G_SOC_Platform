`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7BOvCr68v43FOweNp9r0VHOfTm58zd+qNqNg/s2/tAiV3WDXDZ/Qg8DbrarAqFMO
XxC+gSt3i1d2vecBNXMulTvvm3QH/yi0flkIScSQR9q3QRVoUk41tPsF4lYEnXom
EJVmKlx5ihynQcGpjo0z1EpBQparRpH4CYA6ElbN1/F4o/3q+KHutxiuWlPmDS1w
9HFos0baoD5Th6hKTJGdCoxew433nN2Qh5KPWKxqXM9ag7pRSaaZ+ByGRJRzySjw
bLAuPVTVUCMwR7gxRGE0xn77Q0t15M1fuvCDytx9Q7V9VwrIiIq/mA7qlKIWSMVa
+l3GKFKgjWULdPECVYeLEoIZZa6YGfRdliL0lCgsi2Enhhb8LPjtmVuynfTe5Q/b
mPz/Au3BWFbpQ8Gh/RULRV7cc8M6BnoH2R8aqguVRjgEHSODCi80Qlm6ko8Gbm9Q
axy0Mm8Fg9TVOKdHBXNLB0gPkRrnMmqWBH7KhIGpAIeCU8iy+HMKmalf+H5HdJPZ
nay3gRq7q89ujOGb+lEKjO24ZjXl63XAvYW9pvvzlj88e8LKc2kk4eR4cUcaBEFN
cZJy/IyPjAcN0W5hldIt0K7hoPppxoosNIpIeKlpiFTpQdzQQHQytV3BbU6nIGUG
EIxiQlhQkGVH+WBkAWhJ6mEM/hkxQTtFk+UuR3eC5K6ZS4BNKJhpbuKwPdYzvOU4
H1PlZbBcTf1M1amZ0+gM15C4OnUpAcmsQaUfwzxgnv4dywntVFhLFCr7dpxYqAlC
czoo6ZL/ICd++k72HCzj14Lo6cUU/oauHED67ywNeyTUA1bWsmR9Cge6lj0Z9y0M
0//2VcGRfmgkbQe8jSlbDL8x1i8OKO8tziNPJZWsP+WVuuDBsLnt2dMnk6f570v/
gk+8FFxGx30KEAwvqAMwesqk2BqTECtKNlSMKrHwJuYqLHZyNGQ4FhWKX8dSmZrw
IXBUxs7uQgn4Q6L5M+aMNVA9wzeW8S/zxDuMuojioEPxl06qMfaPvhXjWdW7+N0w
FYP4fsPCvZK18bGh2crH12MiwSeKNN72wJ/IKn9HZzbR3nJKZ+ORLXMccRJ3O9rD
po4jo2/3BlOdA5inimzWsXUHsY3OjHJMQA0IIMtClHxs3NCf8rSaVFN87jr8ybYC
rSH+BtigdEFVlAjRLvkd0Px+v9GrRxi0pfeNO19QEfykLrEUikeUWMoTQAdmh2sn
RZHBUMt/fBD3Qewj3EdtAMCTMOwKE2qEG7pEwln+frAxIGwONfYrz/4WuJxKDpau
hZO2Kbi4ImbhsIGKBbj4Qxx6DAZ2PWvH2fyuNXm6r7kltHHph15DcCZ0Z3HBNko6
pMc4yEdGE+oC7eFyhp0KU72Xjz0XDW++RyLF+ixQ45Cy6hatT+EGJkJHVnIusr7c
oK+5Ame45Haz3pOyY860hEPoCS2DX0sdB2ERVPTNYWdCU00GYvWYcQYeT40KSw3l
E5x1o0cnMxy/Uc1Slvg77WlQbgtDdR8LeS+FSqZ5H3VigRgglwp4hVWDfm6emP0f
W37Wtw8V3klycwnBVXxf/nkxm+MnFLBDx4na3LfkYPTiD0yIv1vgI2QLRKINe1si
TzKpNjASLjSx6dzt9FNV3XR+G8ToOFEApAn4veP7+hDvJaFG2jwZBoaI2VirLGu8
I6DxpCx/iD+NJMISpfPCfmZA8fWKhQpZUeofkrZ4UXwBLfTT67AG0suv284z9eds
Z8HvIsNMjPAUylNdkyPvW5yv6Zbz+kTAd3buBUNLEj09DPaM8K5s4bXIU/i+VvL/
j5/izQGm99EDHVsx/00GSBFNESvz/gKHEXIrH2qyvq1I0gZCFnaykqxs2KnS+T6b
MNgwS0EjVpEJVjnR2qHthxrN1BZ7LaxKExNQfEMcxlkhdgwQH7jy36/F29zW+60i
o7frMfmoB5Nc4X9dUlSaIaECAx16FAKdrNo4/T6qCiDNPuUmt+4hPlMOXs19PiQk
Cx7N+wwlp9o0htiUD1AKCdbWS8sM2eLYq68XMktcDZjVyp5HnXWJnrknzuDQFLrX
nucriQ2h2soyFLE1ktR/A4BTuRPY68xUkMNSfOzh0vyC00uqQ8xguj5G2/tZWkGI
2D4LyUz+lf9AX7d3o0XuQHQd/VhyJzoJtH3uAh+aw2uqFYIJ1W7H8MhGgiTXelEf
qE68kRzUkBwFviNecGAtyJrOFJNDKXFJoIN/DAzzeoVZwKClE1v91Vhq/xThLp2i
s52v/mlMfjnWF8ia5iW5XKc4Nc+ide1/zXWLTDRt5C36j052xME66ovSyk8+mFk2
Dc0b/m6uptmN7vyS+19TsUIEyDQvNwRO1POsHCY/xd8ZqHLVlAv9nhJW11F1jOCd
suED/12k84ZPOBnRJYqavrpuRBVeviuKymF1EE+c1XFq0CuFI6SCT+r1uhU0Rnzt
NQDrpj9rMe0zZs+4Uqsr86Qccu+g2PYgyVynFkipJArd1IrFKMM+4s6SM5xxLJZm
J+SB+IB6IyY2m+9iP5vOb3JB9v6PENGq3JG6nyw7ni+4g+zUSpUK9Rc82iwujAFZ
`protect END_PROTECTED
