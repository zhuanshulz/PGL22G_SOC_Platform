`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e6az+SxAqszXUMIQhSGU4Ob6EY62VqY/DntaMyGIXN9UZrbWAY4VTrBAmU+zbZCA
wz640Vnuvar1wS5U/3MAMHv3j/+gezO1A3LSduyOnxQevThfq4a1f4MSjcogwH7r
cQY+ROrJ3N0qEwM/Eb4wojzzsFgpInmjLuUNY0Cqae99R1ygukD1V2Zu+BPwM5LD
fM+ATSzOREMTz92ca+M4fGjqBlU2D397nhYf58F4lYQaRFMFakscCmepdp3vRhKY
21xA98AVvCVjOnvG7Gk8M9d4FZU7xp6srSGjBE0QEpFvrbaHtWzU8HFuhO9pkdU1
+0Zdgrd7mDLT3n6M7ny8Y+E8VSI4Mv3dvmwHrKERzwawYRJzmR/QZU8v3JHaE4x0
ZkRcvC94pqERi0Hl+hNSpBTdAUup57j62G30+myLFWaTyJbkGMrOY3/hfk4CX+Aa
7bnN0vtcWquHXOrRnyleW1Ys1SvVA7hQZ4t++Wl8QDTvVr/xL8A98zIDga91Pj8n
dgRUAkRsn1M/+KbbAEB5JH9f/uBK9gjWofAYueiMDUWblwf1fb5ujh5mRzWnSS0s
jGNc0x9vLms8SecuCf8+8T2loXAJOK0R2lvZCR1Dlo7tJ3ABJadoTG7wIBJL9D0F
9yC+dBsV0SCwf7dM8w8xJsRIHHT+VHaPcuSENU2AQU5Gxof3X0pg1VKqKC2rNTzi
KrYjlKkfNvT2XpgR1Kl2JhFr2JqpxMpXEqGGVRsTcPk=
`protect END_PROTECTED
