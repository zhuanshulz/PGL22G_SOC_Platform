`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z/OPDiezsbMlu2dOyaYEb+x8mw9uUlDd2YEvM9vVe28FbVM18KSbFhaz0ooE1Imi
baUKz7jp7Yv9jMtbaFBwUkLc3vHtoaAJwVlhKrj2AdAFYFnCu9jValCNRJNwJVVJ
D9Vh6Mr+Cy52jB+HzMpkznsZwxWaG2WMlCp+4nMV8fbCdxsJbZ2XZtpR9lhVYOIk
9wY9oidVhbK7QxCiXM9WbVZVygOabS7cwx+obCDSr/Hw6QXaWLDePiwO4/zzgKFG
Jq7GfnGBPJlM9duJPEpPsopkbMmdQbCKWqclX96ZohNJ0roM0slqGSieMoHgQo4f
58Tu4muYuQtCZMYekQCQ3wYtV66k2SSCdkZ7xetCbifv4Cvqdr4o0S1tk2AlAKSR
y/HtOe4YCvbnM6Q8mcYEvNyx1+m2jAntQ7wp9Dw/15Bwn8A2Y0BKFrIgpKxdnnqE
vJQggGA4bBPxj/gxW1bv2RYd4sVrntUBVg8V6YOiS0eWOS+Jr/ODlKDEBgKiTMUG
T1gxD8p/kr/5dxPAnd1TT6EUZ14YqTSn7Vnokn98qrCAAvMfgzy2Fz/FPAjVdZVl
E1rZgZv9/lyI5Ne4JAUATdGe+cCyXnI3o4E9RZ8+MpmsbIDBdchZx7DENBUpu8U7
GkdPZz4/KZAWihDunakjbU5FBo5TCKGOdypzoYFlxeZhWRepP80fdLdGjlrnsDSw
SMgERs5MhNGhni7oUYPV5Z6iPi66Q8IVY815X33vYgjCnfofmZYuFUeGXyYQCn9r
J0xU2Nq+x8fx5zdhRbRyrXBZ8MTJbeeRsa5OdoLhAgMp7b48+aG9lzpaFdcO6Rjv
g45WFZxlT3Vc9WWfZIot2Jn6aERJio/mbXdGn8d87gJOcN238A4ZAxPld+ovYe1A
4O4c/5A0mgjaEDFv2pVTaCkSkyMPXaQnhWrP//7WilH6/OqAw/fxIVknjOBjfIRG
4vyjT89R5K6sE9Kpkoy0fipdtAEWKtyGgOHx/RjY2Og684OtR9tl7hp791tfkr51
NG7uE7aedBJZ+5ebZSdeIeo5skMO43sbYYkNGzZATCJz51i1mHNNJhiaRPqpEXVY
lBpdW/xW0h71iFSEOsQ+yeon4R0tvrcGubVWSwogJEZLwzxlsSNgg6iUQfelnSCN
AddTnBInf7EBa8+MuPDhYdD0+7HPLahsAd6ArWAqheajGKoqR+fjeqPmB71d0DfF
4tUenYBEyEVjPnckCTWQOQte9WR+v75fWMBqz4MHDBtC4qTSF1QSdXEJNBD81jR9
s3ETvaRQac32zEGxrUs3pK9sksHIwqiVGM+ypROGPxuc1j0iGsKSxrmpkjb0alu1
19Ddfz1hsVXBvWa8M2RO3qNcBlibuBTt72zQj5smqGKxw5TuOeBHCJAAHRsvBWAY
DHlLYYikgPlBG4coLcv+ms0Xe1ZMIcUpzehbrB7mZ8naLW/x6oLic3g3tmX6AR3k
X3Afs2AXemeL6TA2ifPErpMH1/nMGJsmOIsL/BpZ3c9+Uw8yTK7sPAZCD4kRskwQ
mjRNnS3GKqqu3Fl0eSmvISAD1ZvhoM/C9vQkz8PEJptto7GalsgG/DuymYvsxKhX
eBo2fYAUntVcQ93s6mqq10qMiP2BfFHpDtBcIq0aYo0OMY4xWY3BsRTotKquTU7J
Il4sc2eyhmJpxHCT3IiZtMTEpQJwPFC4Rj8M+Q9XJpPRK79BThJbGWJX6QufWA+g
s2TVon966cUkgpYPEq9R3WsfvUY9XVsQGtnT6qPN2pazheukFnzGhTIX3+PN7iZO
8tf55QVM4+WxfZT1eUgDIZ3zuvLWVyok0EQWZksWjQ3/Rpcia/V9aALsVMQZTgB8
+w9Ob8e/JVi6zoDeRFT09kzFNx6rWLZfCfH97n6KBvNECFtAyIstiHcrN2DyfoKk
YUjk9cxab3q7v6esK6hnLVyB+RNinhVqVhSaIwFHf+hJN1NBhIpx8ZianlVcf46G
Tw/ifUXup+aAtI4FM5PecP4+//aOfbqeGxgezvaCnWXOZ4WzJx1gjnijrszr3P2l
p1TaB6NtxzmB1OiOhxEJE4o2zzv4PzhoMRU0cN2rXEaxS5PORSev0tLSeBWQoMoK
C5oXJ4QlXpVnG9Kd5bSjyVCAsWoOVs6rwMsm7XOhFPOi7JW0rZniU9oC+WTySzZg
tcXey+QX2IURYxZqvNt9Iv7zNBbx0D6trbJwdz95KYQI7Yj3+n3XYa5Ij3QRa9se
+tXNEmfNiSecRtkWShUGY5U6ktTwrDLV5TH2Wr1BCS0O5SyEGxxQJ0zwe2oeuksu
moVu03TmjLTADZUn4CJiUHCwZsllnub3035LwC7qJtRDmgURWX8Mq2z+i7MFcrt9
AuduOQWi1ue9bte4vT3QQjO/dCiadq+dchI2u6/kdS8qjAsRTOSKs8vymsPciPWM
3B5QnCAIvtvAgNdDA5qoSMNM+562SDkC+Dly2GQ6ZVBN7P3M3MoJsetn0ASCdBu1
52MjZGGTfbQRYlQB/qDVrDXdqJ2RTwIOHchDe5DBarzIUO5qniU7VufIRwy6wnFE
2yMV/BeB8BKqeDq1VWPdMlFEx5HyS9j4RMaxyTk+7eTMX5ZTnL+b+bpN+habENqF
IMt/AbYgJztVX04VYGKFRmTqYOpV1qIRSRgu/70SFxnZ8ss4vCWo8wiFF9a5iehM
FoNw78neVrZnE4PBq8N8YdrILMDheC2cMPcIAgd08/tOxwfF+FB3Avoq2sTrImY7
PAzQSK14sjExaXEnAGSeT2x71QVt+gRVFF7Vjt2pU1CjGs0QU8MZ8Wwv9T9l3YPr
BnkGW5ZTJnfeT1XtMPhnW9lwCmwaGJVUyDqgFXe0GiUrXAoBRtUQSha7vgrpKOuP
1VUJ0/0MPoMJv0wIPIgjy8nRe/aiTL8scq5koQcqR6KU8/OXOz1qcMMD5NHfavvq
3pFaNjBHFQhqB+4ogpfelvsX8Pp73uVMHgXQrkpUDFkJTdNGi5Dzu0VM1zgvuLth
wLrzB5YD4NpT6hQv9fPtLxRTycFkKvcBxbXsvC/RGWodb9q6PcH2sazLlkp/bi93
h+VtMBeDODt2vWhkfKnbGuyf0BIhZrzMUuraduGc0kQUqXMwlDfS599wYOA7I2Hl
1uQJfPrHMb8kotwrFV7ALuXB+hcePIk9DUYWdSGVlUJR2fWegqKqbs9bTyyL9an8
ALx+ZrcB3rgf5MvPBLd9a0MHrfurjI4KzqZZYyq4H5H3Br4qXK7kBVlc3IFS5jPk
LVM/YjmzMeKBvK6E3MjEeNwyw2PoqSKfJnsEpl27SJ041BmMJswTT8uyVGTso+Kb
Yx+2P7Tn9QqEfRIzM+pRcPknKgYeRANsqeYAxip3AcEei/rYLxGRQVwA13MAj+D7
8eFgliyBYn1moQHE1pfdZQ==
`protect END_PROTECTED
