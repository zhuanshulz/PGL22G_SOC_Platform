`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y6p6Rz7kUGFIZ+j+2nOpFGME6mlft/Nqy30yk8P+PMQHiGvEXbV0WRkiwc5qdI1D
67y5CkjOOVyYfo44uxXuFLQV61ZWvnf5pcEChtJxDlPfjkx4fOAhag84x14/y3lf
UUdSO4uZoJuyZ5fjHy5nyYabKyIhk85AncLu2AoHhDzSiiX1ZzEb+liqy8VZEYse
j7YRA6MtPIYYgRkE8xpPov1aXFP05qZMWl8fKoppyrqlDeEb8rxNds0H59PLN629
axfgvG45TkEBlDb5NAmuFtbvITOUpYCt2IaSpWi5HZW9uwiPe1hiriwy1ampMCoq
omOTb1wObswi1K5s2kvP3vgwc5+gPx6CkUzqc6CN2GVDqJL/VsxAnHYRDz+s8wI5
fc5//ezlHrL/ODi4ordBu58T51D2VZhxDVgWDmYMpLlP0g9GX61XobCvTnVwpwvu
HPQ3097lNo5UWKL2F8a6hoJbtcDYEzGHNfAfU3S+36fOQTU5hIeZcTGij+ScbUL0
HMzSGXE33Z0vK8VFFat8L920C5Jj8AwiaGBgTR4tETw=
`protect END_PROTECTED
