`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oo0Flker2GyoeqqyqPpIsqPP1KwB+uMpKTgaAYqTtut2ySMPTRD/Um/w/ytmfm0l
1jy7KOUNh7UqoPyVbwG6d8Vsqoy75Yb1lvABjUlYTM2JQuIWdB76DlulXUKz+X5x
6Qj25mCfrLz2rwAQ6iWsO3DwxUVhWzaUFlXNWud59MzynJFmj2ergDhoxp/kQHyW
y0U/9e2cy0A5y2owlgRfEtFZ4Gfkdb4Gnbgdah/7ITbbtttf9+/wOHh4bbCkcVf7
hUS6m8hg+pEWQwZzp6N447kgD+h7coxvTQJs9doLjPtwFh2wGoDDtFulvG109ax5
Si+U1w8xT95E0wXF/vmTFgp/jCa9AOEdG1A6Q/x+ljq/L8NZCkt7XK7GrvGNUKhN
XcwFvxA0wsNSUunL5TiaW2K6yeGq8sA36dzSPnWC4Y/N5PeBfT3RlXQGk6imHYdz
h7TudTPekxrKK7h0ovtSjBlf70n+K2u/VziXcp4/NhzDWuIJCeuCbCgbrNRkFrVB
GMCpMA0GjT9FYuJAsAJu2sr00s1YblzczYwhdDhaMKE/VkXYDfnYIH3QIC7yOKo4
pCPA6yXJosCdwDSC57VPwCwNbvxV30hlrDOUAzDhGMQWMDhgdtForOFggJK+ykmE
TGv3cSotrsBnko05CK7VUNH2f1Y14uApkGx0KK/2G5RNOiqcU1fJ+WaE2M6oskot
JCf+9wsppbgnbUxM5ieYBo+BfZ5dwr81WDdyOO1R8Zin0o+KkRXt0LcwisnYj1B4
1/BAcXIDgzfXd78BEzPWYSuNakleOz7/f/v6k24uyKucZ2DamIBgQ3U9qvr2n6aq
`protect END_PROTECTED
