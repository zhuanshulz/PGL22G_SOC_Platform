`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dByYG6qURQYuUt6fxlJ9v5l3teLhBm6lGCBuDAHo75m/geBckjmgvDLLEgYiiQc7
tXFQN525BIIB367l6ijiEYQ8rMoc0PLhKYpOC/QhFN+ot0Z146QAu1ZB+qLV6LGg
dvykjOZwtcUJew+cwrwg9uiXiE5ycbsbaZETMi4dHCfawrF0/f2+utWDK4wjeoY3
SdyOJf58k3qn1aRjy14hDJOIXNW006gaoJCKBhfhPWMHWbRkpxv/IiN+0kQu4NAK
jfG4VP0KTer/bbVO/uLV7LP28shZNBMjHiUkx7oDZPZNnS1qduergkHk6S086msb
SMGvwH4uQV3yy1E5X47z3tx9FdW+yMlkRhKM8QXXwSPvlDKZYukpTcXbBdGq/XYO
7sjEhMr4dGkP8VyabktLaFKB21F1W+qsRIIKhMOUOrm6QasxaG9sS8FosG4QcyrP
CrWaogUenGjzBXTOm7o0KdGPEu04ATdpPWaBtSjhWm0VNsoHxXg6J1Dk/LLlZQH9
YOxVhgXc6ZTslksoAtfTAdbdZ7N3PWIqKoM7nqioAFZJxQ/8slx811TS8gWQ79IN
MizbSOnO4RSARs7bXMbHy05VmefXx8eB8e3F2YtvupuNdLVBzW6Bk/fVNnB4kxZ4
/sPdD1J9ALOOzMH/Xzcr/V4/NWuPHoZFWhYawv9e4oS9bHiuXnwPB8zEMA8Jpmzz
fHFJt/X2/q/EM+9XuLp5TRK8eQKc6VErYo7+/PRhEH4dfcjgLklG8YYDtjjUe/RP
FbGBlvJ/5R5gHTBmEaQwFoL9jHzBdkRpLyllD567KV1gFwzfhhF5lqiF6Au1xv0n
fk2kp4wB5rAOXmHvG6rg9uK55vv2dWl/dPe+UbRLYcM0NlfEqqfj7h3h+XhL/+cj
1ZvnB7TEVL+CE994DHY2aU59e+VBMk/vpgngfAsZSvsNjdG9IXiWI2qU2g2tXE/f
za6TOz5Z9rV5K01Q2lhj6vNyxfTIBcfk1Z56mbUmkoDdajgkxLV+WPmtrgDPJQ9R
8dOVP/qML7+G23MB1m1urny+gNIF6HnJIc1W+xmEDFs0BgNrbcAQ8gqSV05HzKlR
bSzg2mc54YsPU4EqItefbUOzyRvkmiLIPSTQ05L32um1eNOXEBb8hNZHL/TuBoox
obfEou6kOuXBxZUDY7gGe8bK8cvY4R2E7Q01QELwGjAlwiBd3OpQFy/mCS07qR+q
9YU7ziokicy7baNf596zH7wiQIkzvafQ8RYL2FCWdZHRXl/e3extOlpDlhBsFHpF
68bxp699weohC0eprqYH4em4s/7w8+zV2q0VGvC0WnCznbpwetpBTeLAS81XHK0s
JypSTBchaRQyFV/m9UBAhXFAxj6ingHlLHb88lturjRgmcR+7firhTsmxT2HUDFT
0OBvEsKAQe4VQP8BlUbcfJyv3CCd5LK3JNJglit9zzWltrhPyAw4cvKp5h7eJEss
NzbhbBFQSDBGRxdvQd+le2N9tG6pSGs2L+iK5aCLjczMvKwYs26Lf0pcXHAzo1Rd
Paf0/723hri8WRVbEZ+g99Fv1gmacX1xaVvJUHaPGX2pCy3xWRFB4R0fbxWS/AcT
GBGg7S3mIry07DiQEuzBsuHteQEt/cj6DkyhBohAzINXeXQ2Nd1mQ+3duIymTGUd
MlDVNX/0KhAaJ/aZUCuGMexAVKMN/dZXDHD0nZNT0MpJ28gjYKpEwWAGIcw5k9rD
cItKcGTnqTet1HbLcfkkP5N9vMwDJdlfgTOcod10dVdPgKb0vYoyWNJqBna4IQaA
UqSl7ti7ze30DwY+OUkjKdQIAKMzr8TYetEWWBP/+t4fXbajgs9A/sYp/wHn/jLb
5d9ArCgkPdZLdiiSD6plDsBse8kiheIJtbkEj3MDedqHRisKgUQPgf4WTBD5m/3U
YOcu1Ldx/ad0l9rwhxAfmJf7qQrJ7IW1nbCoBBQP4Y55A9t0LzutfIGfhqmUFtFV
R+Idg0aD4Hl6gtePsQgoxvkJp5VP5DJ2s2TnS7HYF6VVH3XfpPkpcgnhH0HpnABL
wX6hMBbt+GE/+quVwiiRrvuJMJoB3gFgmv4ZhfEVR7wPrXzTYiev5r6y2WCQWl/A
hA1413Db5qkB5lEiVlQJ2XUKGP64mgimOZ9u8RXxuEyU+/vcKROmHb0kAbhdCTcz
z4YnHX3NQnBxhy+p5gWRxi8As0dS2lD9wb4Fzd3hZO60l5gd34Vkn+/2zJzjWneI
fU0NRRu0Gk1JbAbZuW0A8UCYEoFw0obuceNSxCpRC5ZN6fOdy6Fb6LIGY1n2WKay
d9PblkGfs7rV2PXd/SnJmaH5cih0KuGFtzipC1SxPFeTrtK5ZpVEyZhTXlPqT1n0
2M3FCBVRnijDBDil5BMhvcfdQg/qYPbk1zaIMEE4AeSw7taGy0tZeI/m1Yqw7fZD
buHUq8y+tW2m21CP9kfZsM4ksRfw+4yqmzEQDY7zkY2VcgPr5wtOkId87hOMjy2n
0iYyTJw5TbgdsAdCoCuzGpXY4Yhd42f+EucXn+yn+UmL3rEJvxbRlx3KUYoZlMkt
t7NR4swTyAvTSRENtDSTYCt+0WLrUcOOJtAwbpfQ8WQa9W/FIcdNNAGlpakgExvN
1oRTi5Yrca785EwQkM5ZH8GGzBLO6inrg/Ns/aoF1Ik0mhHdFpYA3IuctRV/mEeH
LTgFVwmFX7cp2k2J49aU7qOxG0fLXdxxzXmPE7was2iSotKNWLErkPt7rSIKpU50
378rXHLyiMRrE4i68OnyCLnOhE60Tv396JXblWU9ATxIpJjG6+Y81nXf48hc0eXW
fK07e87Esa7Gx2zWmJTxAQ8rEHAY+ObgTKc4X8bmlvS1QDunF+0tgRaUEBYBDzi9
jq3V+8SL5YRNxKWtgKokZWGuWHg4U7IxTEVEc/foM1eZTy+eaDVYffwQKxSGZwQw
VgAe7N0Sj2p/esp+R0dRFYccylw9Ves+b2lTz+Gz1R9ip2nXUX1myivGoYiK3Z2T
9M3/deylzZAmN58+w38dbci5RJrPXYqlW+xvOQA/qdjj7+Hj15x1FMf62OgnXVTO
3YELK42OVa4Q8/Bx42N4PGzN2/pHffwksZHrsA8YE1OPy2uZ8+cFv8U7oxQyBN8W
JokJzzM5+Esyzqdbv4qqsMd3jfjbyhQbT9m2gFbN4ut3iWZ3gMnhX7AS24JIX1p5
9S+uBd0xSBQJwUxRYiXOZAg7bgG3HSB1O33DN2wk2fgV4cJCwDl2r5f0oYdmizqm
TAZbV1ixvaeYrGRZJ1PueE4mD+/Aen5znmzo6pSVCO4YkzjtUb6Qq/ENae17y1zq
ZBp5IYOl60UxrVWn5FH8eX7bX3BazP2uYsXLcyIGMGjrvHC5Fnfkjdxs9czD/WB1
WwVRYAzFSUor60YNu5GlYAXgV9S4TGnD06eRCkLnhk41KNzQVmZuqsFZ8qCmUhif
egEGN/5x7LEutczEmyTZ7h+8G1OhO/qJaZe0j0zFy11C59MYsqAja7RmvUuQ5N/n
zdJEm0BTroumtYq+0QTxAXvW2jSw2ruYm7A28I95OxisY+5kI3KssaC9wz9+kku+
0c+4/2WkRRbMCnVuBpmJgNLxoRueZiB0y7G0TuTw3HSymMHbFP5BQWJcLTQGDB58
qlmh1lKfIdqeeF34GlnLsWdwQq8gXZculMGpGpVNFjzg8HqXlf6yVvWeVCMh0N29
vPVNYppdwK4c1beX1xdG7gw6KyXH0vIgWSwbI5XIZI+E66iMMA0hxIrQqf2e3JMR
c1liioqDHU/z0Mo85W9N8z92/+Gb+THqCLT6C5ks92ChWkGaDuR2lQDlcsd4nLIA
e/HV9en3CsJNUmdPKJKu2XUI1B12/C/OE6fZiuaavBUdXPoV6a2x7RWiHrw4G0FY
6N3LJzwQLcJaDkOOxw5pa1hHUEj8h7f3o/IhCvM8QMyuDdR9YzP0AYtpRLwmijUu
Iw9CFHA4cnWWzWRwOIWlhFxUqZgnuoWVxwGwMvU6YKfnPpluRaJvzChB9R/89yGE
Ht9aTDFqdTuyAJ9u+QneVt2ACDFAwlm8oexCVvZSEItKMO4FP05F0UWP4SExld5E
Nt5/22UYHb+0FHKGB6lVs3mZA1mAbGngbpfvPGvfU15yfOaQra5AuE0P2v13P4+q
EYfMnd6a8AL0pA9q7RTYQzmIxelCUyFAW3MI7xV2KzUUdw8p80yNHzvVCZbaQmBH
qoQpXc1S/tdFWvVVqrKXWX4LcohgYsZ7QrfdWpXmH7QUpcIVAtn3xB4t+VrAEZfZ
hbDthbB9Hi8NJMQbBXzZ7H/VrngN/U2DCnsMptxZ4OtDzE7cLuTyxBzPjvQ6bqVH
43UPOgjCz1C+YYlyNRLoZufzc4DlOaLJmU8E91CexjH7EVccfOmid6T06V39SKjG
k6Ql080vxIaCqvAVAtiNOaEAUcgJ6zR1T7A0sIlfK0US+vV2VJlfcspjD5y8sMC0
nUk9IoRzcJMKsMyxjWrZnWXcRG3DyCKufI02e0pQncid6N7624/23I/NN9SI4Hqf
R01Fez8A4qaD9jp+gFlny15hugSJ2g8wbdOBun/B1+bt/9qCaglLo+tT85aEKhsx
Thj4W0/AqLcjPkP1xSiiqRlj2MZumTBxsO6DvwtXVZfGLdZydQUIG2VaU1EkoXd7
xM+vWy4XB/bVpFk5qUyOWptDt4QAiOvSKGlq1y05UNLOrhsTZ6kFf9B9AsgDYYM/
tUklFoFBqSOwwvJ0/Ala4WvNXgnSWrY25N+B62rjpcKdaHKbLzgUndm7tvUthKCX
cRT6A8KdY435p75crb0jeUkFLXlae38GGKtBmaB7HtJqdSFXrXKIYIC5CzsDSiGD
gX20IMXwA3PVRBJdTod1wZvwOsBs+MPiWehydjr5pI9jsH+s+8yi3i1Van2gfSrF
dq9u6L++Aj3j3nSnFVJCEkSrsA0fQ0LZ+EwbzQ4aOaZskexpBAsV30ziYqiDmMis
/JSzt3RWqPtmzrpCzaIZ3eosHjs+7u0q16aMqozrCKQnxK3gqbaEHckR4prq9Ew2
YfBI/v9sik3vbeB0E9sZDJRwGApf6hEmp8GUN3r70Hdi8cjgT3JGrOR5lW3v0x9n
+kkT3qgQcScHb0x/TVy2+CiPsGEiNCkNnKkSMofwyyqP6OyGc/pEiM1I1JATG/HR
U+cqAgHIKYfZQhlToEcLp8g8aIa2zEBC282X9V/LlMzIspbNrWloo3l+t9zH+lmQ
c++6KAufkI4cb8Ao4gOjwcGOdx651UQZhxt54fPjgmOa/YuuWzX6AyBruz1Xaep4
PUVDYrfWRDfOZLE8NbcbgIN5RPwVSMLMIieZo3kC5VCSHeWotKq0v9dIK9N7q1gT
bvEwhByakt249rJG56I8VIho9ih+eK49MtzwjU9YnvdhpzQYtqd92MbxY3TtoX/A
5jhH63lmI3OMRiwexURStM8GFvb8yCAimV27zMppJJ94Su5Ptggy1ppWiQA6Q5C3
Nulx91J3UQqa5tA443bgMTj+ju7kGgM/Wkad2NNTZu9L6AM2Qpmh23sPVsveitqd
caOLf5y1G5I995U8/hiM4U/+4rpdaAF98imNOR+7uAUYZN1QMmAiZnEtg68wmFjc
T/njki2GFzpueVNRgEo+5soPMpanv1UePSIGfUAdMP/hK3Ar2LqRhchRdHHf8hsU
0LSNEUFKzEMH9pMUmFhR5JysH2zYi2ikDuekuES+2oUMo5Ghp9T402i/Punlwjrh
v1c9OZGJKa4Ys+serCp0s8O8yzZ/E+QMxFSxmy4/t6krb7j/y6ociFvyS/wpcG4n
jFujB2eKAHwimTng5M8bvwc0PM5a4LA0cnUqVd7eiI81kQYaF/qB+pG3gi5QthaZ
k4stwiALgRaZmGCPts+2DwJWmzqjOhskcCOTxOZKmvRvjvpS5U0jfe7RBim5vsXS
ViJzpArfrjpxSonijCwdioVOwe3wRYKt2Pg05nH1l2uWejPe4r9BhxbxgkXWDpwI
9gd9yTTn5z/vmttWYL0T5AtEqfQYBBK2dqG5Z1MhUB765G+3R+NpA4pNYRv5th1T
nUYydC7GJuRZ9Ls+sI8uooe4VQw8eSDknsxjtOem2BvzQFKYdu/2t1ejOkC8OtZg
0Bg+1Q/V5zlOHBbC7VpyUqcT+kOIDTS4PTSNgsupIiLDmMJ4tqwIQBnNwT73P0Zi
27rOaXC1ADmng5Zaua2VpPGuDPmX+b5l9vtrOmWsrl+GOwf2do5LmbzqGHShdpM1
ZQFeFS1ZIX8vs1/YpsOkZMnWw+BlsKk9YldX9UJSHsifOcjJmeQYkdBQW9OxS8Y5
Bg4lvBZJpsipZYReh9ss2uvf632u8VNKiORQo4nStZn13zWEb/vBQwd6jE39bETL
QbQ+/PW+eYp/qCATN3VblCmPLOF8eWzzHVBjNJU0BtM3P1UGSkVTnWocueLvgyAT
BNsRMToHkz+iTQCIGsnq5cT1BxUUNud/9oBh2j1pCRv1O/FtYnBOVjBdtywbn16N
ta3cmoUAgVaB6S9OC82GWxmiy/wJkpi6MCB2leZMm3uRjHN/AkRjU/QecIlKyRsb
ix3Q10+m0IuZr01Ldj8zoa42IuZzFTCXT9sov2O1FMFWC2h8VcM66LXQI2fw4LvT
xYMYffxlVtdjkWqK51fNBA9TSbSknJHoQCKGIUhGjOLImcX8KFf2fcSJPkhvjYIA
T12IksgbVeBIew/rvo+MutVL60lC+GrODkLAt7TmAygN8At2+gjSC4tntK7WFTci
YM7/9PnohoZry4TReuMkwFgmyT82hPTp4oaLiVv+737VuDu4ZwvfIMAVHySJ4Hmh
TZBlHCNlyERJjsDvk3cQlAy8JgOAP+3dBGcvsQcDRy0WXPlXE/hrpJPuVWkIx2bu
1QAEtSbYqjBk5BAWfWfEd1uRUR5IKjrwKgjnZ7p76qOr0uDGxaHbW6YKVXb7rWf0
FEBlfn5Yj6IKWtsZM7/QmEmceBoqWGi7kT1Qxpre9uN1nUTtOYqG3epFPmPOajJA
GqjipMBIU4ZblRWHqAGfDag1Gpj5qK8GTff/oDxqOUKqBC43YwKkmv1Nh8LVZlrb
ro/ntCj9rmP+hmVvs0NUG7lpbTO1wWRX0rMRn/eVBH6b0g0voKUoB+ICSsiU5U1p
50P17xbwnmsITchDT9jCmhDQLs2Zx7u7MdFQfU94at3kXaAZMQbe13CubP1FzmZT
Pd3uMhpcxwuZUtlJQrN3YsA6dY4/5YcapaPdOchcCWHh0Y8QgzEGjfqodEsB0Xoq
DPwAATZjDDYW9y9B1li7Do0LYgCwxau5PEkllkJRtaHGbcMa/lBFZbO30cw+/d1v
l/oe/YXZZ2/Rb+/fwJK2smLRWJD/tNwNfbyVUdiauJDidK9GEhrHdcrgrOdlILNW
oFs/1hG3Vr2vkbiCeaanGyoCUDscVaJcPiO5BSgxhb97G7+86ibgAlayzsajDfUp
SLtmNvasLvsdctCX6LovJcGWE0T5C1oxByT/16EvAZIEVdN55C/LCjcd08Iqoq4S
BI8GNxn/ueybg+AqoKFCvhfHkmAJ94c92pkxJangXazH8qZgBM9acQaYnwDHfmEt
eXtHJ0HJT1j+PRRAyRSqSRPugxnAwcGHZnCmnGggVsr63iI5qalBIcuazZc1niRb
pXrHlov4LdKGsMvuZiKXTSaTgGvZhyTmcq2Z5OFDQ+cAzJyKE85U+4Ocf3e/JjNE
J8WUuRSKbWvzYdkUvIHk5mux0UjtWQleRlS6aoH8OiUiWutE5R0m4GSgIhil4vZ4
d8pVMjPxGTaJhd3oGYn4crHDsLqm60igoSAZo30rF8rGvyDFjD9jOzbfJB/d9JGS
MK0eUipCxGvfW+nuI2RR0Ka5P1IAcMbXzBIenKvDSD0NkUgmuScAn5/v84n7Sqc9
Ws9nhSlFRA/1vCI+uHx2yzrOUPMvoEUL4/KjsVOX6vxtZTV7SE3xKn9mAmHCjA+d
M5xmGZENIH8h98pRZFU97zN/aN8clvwUlvkk3D0jDe1y2kMUNOFAtwy8CaKD15Yu
TbONY+qNLulL8uCnNNZnEbtcEDXur8v15Wh2ghFJ6X6ajMw3SNDeBQtW6E//W5SL
9lf/x2MEaVS7Z7Lz2gYemt8ih6PyAnX/rGRed5+8c06sf6OciT7OZMGMlKkr15mB
fl3OkebTRICYKMS4z7oBhc2puHbKBidswmQ0Rr5BEYex34vOo7RQ6k3NWgh3GGfG
7NfTGo2MlrlfQOErEEyzoELHHltkFpA7Bd+9k4Tq+wtvPelrVuQIk4IjPARgItG0
R28OSnmEhnLKkXTwLgEZOnUqKA2WpSZ0B92hR3ls+0x+WlhhiJ2xasdmeniw41H6
nDUZ5TrZqHEp+jC4are/vkW0zoVp6NBqOLfIF6g3fvQdlYitk7+daZFtlY1taAqQ
X1nSZ9dKh4BNTo/ZqMB37Fdh3ylaxegCg5kmKxS4aPjQv3m8zx9ZkX3+nIabhhlb
93OFY7JPIlx8n/z40lss4ARx5Z81kg/UriXvACmADW5Z/KNp6IT2RSfEhHHXOF6A
AikxxQlMhMuOBjBCGdQzuZIisrpiqDO/+ZMkuq/xVCC1+HwhAoD1qbt4wkccHWjz
wYU4G6avu2kWumJMPDjy5rxATgirmzBSJ5eTYifyzp9jOSmPGG2gQR6hFF0LYfnQ
2dB4Q6vmnWz/nWUhIFGIdzeSnWTurSFrcbPuvzUunhQvUp5V8R/51XbdYeTTXtNa
Wd2rtrCYwOdTozMXUjWFtQM61sZuygWsRyXbxGEaN58XhRr8wMxXYbUvho8MDGkV
TdDkUEX7QVsgj05n5v2v2HAr8IguuNb+9l3YKBfQtdxGF61QHey+KuDaMVOy+wxA
Q0uF8gMfQDYT8MYtBtxA/Sa9lpt7DQaitfLnpcvNbr7GW5g+pIGTnwQSS35MIWqv
GSMff2ZyB7fmLyxPWXSuopLIr6yDdKtyDXWNBlJ8dr8HG98RrXvyWFji4r4Fio2j
+fwoCoqD9smhXnYOiVQ1OHeWB75Uwp5Wb+s82U2Aqq7b5f8JVdhii1qPgZuqu+zR
xwE/yfOw3RRNThYUgBd7+7U3927wuMpkXvctvn5cJaMvTT2Z1D8HLCrMI7poitz4
b4OoxlseNV8C0po37IAeeak6pJBKTYmKchGyRSIjjYMTyu77/82CA3kX9cWVU+K4
d51x3v+2XsYrzSvjufD8auUexcSHW1iQZMXnbwM5Cfkp2m6XXj1R2S0GZA8m/PbQ
emg7yNQ1eWOof0+ARuaCxxX/YVtXazBFHqNexEzG3mTe+1NRJ0JRMEJB0RI67uwb
A17XzLOH1UIwMG+GKEzh0xTLEC55lMUktQkE7yNkJUnO/yRq6b6Up3ciPd6PGoVz
xr7KNewUJH7pDHUxEdvUPgK6cGQcLhP3wy4MmWYBVTWR3dvYplRblTuUa341FTsi
gXxB1Y95bmljIYURm1IBaD89GMaJjJ3rBWkLtMovN6jSHpU2zBiIbBq4MCLAH/aF
MIBtydWW4jjRc7dLewmMg0QkvckcAcMnM3KX8hLTdGE1wHTJZp38fwCMbBu7v6La
0jeO+sj+85IDCwUxOFusgaTSW4h8hR+GF5tZ48sivzIppE2SyJIRRn3NAjNWFN+y
k0/8tIyseT+7ilUfIeQDB+LRWQJ6Xk3fd/KKQWxnvwCcZxQp4BaX4iDo0JU1taAt
fZK122cBBCdRklpqBUi9GP4ycFZ/icGt1bbO85ES3+Jii44taKJd1sD5B0JXjQG/
RaUPJD+QHw40KuQhA20ozpFKS+fx/rhbOi8jPz9fZ5sG2es44gNtWNwuW9S1gc50
zSxWd+q5hb2nfs3u/IcdtF3DrKBRzMLap0im4e2sjkegknA22mMCId0BjXK19XKb
wH1YsTYRXov9I5w7vxcRD4Vzc9KzweWCWL1lzA8HuFsXtqiKpA8sZ+L+upgr79Kp
YBtdpKc4U/Coaz1bE7aYfUyGwxnW7m1xTSXczns76MAI3LK8/x7dCRtuXWbNp6ca
sJbvALLZPKtPmko7oZan/o1uTgEkuzZlwtQLtGya4orihYgMlHlfMuSIuCmnPqpZ
9kfyURXv46BufdwfZPuHiU6gqRZ/+SdK5suMoir85vnyxfExyAkIymucS0YyqHur
JaWNpxCmOEcmCzKRajJlqvBaesN9PvxN66KQU1wjGfOLxFG9szEDCZjddeZxZ244
BG+lyyCP5LNWdTWlkMDS/mKvWpEXjfCMYbWTxTuuc0Z7qQ5yoLsLh4xkXscU5WEb
fHkrU1bDRhkMGY4DrPtOGdjnIBxB7Dol+FKMQTILnuNN97+dzfw1GYyc/A5cXyJW
xjfY9UKW15KIqLwb7fLo9eMVebFZVZrlDXTqXHEwqtJS2zfQGBuKupab1hhpigM8
AFSR0GlFbdk0vrIi73Uhxheub7F+MEyEs78rfQ5iZaLOwTZdDv1uRvRmcC1xQ43W
WCJVwPwbptvghDqrWjqSQcduOPpYdoJgDpPXG6Yv2KOnLcK4mK6FIzJp0g0Ps+Ra
QkqF6v5fTUbBOHjwV4lOhyBg2m4iK7m3kHd7VnE61bdcciVU5VJl9m3Lpeuj+uYd
HvRP7hKhrV7fumAT6FnSXlvQkjzObOutMH1RJ5T30NxRvlF//GX1ZA70J58VneKM
Ssxz28/UUX/Fn1o9prXCSzvxNnS7a6MwN/FNGxzB8NKSz7jmuQGOFHDvjABFOujz
UYKXlJfTZCrAFMwa9UWVQvNZ9W7gZEKwwQ99ftHn6fHb0/JmBL5nf5EgJ51jnYwX
AVLUkKXyyykyqCXmu3VgFH+ym4RTyz3aF/zHBS/fwxQg97W+F9S3dRrKtvnqLSt7
rkML3dCZ305X/okg1OstTSbIKDgOj6TwgPEYU757dg8NSg1f9YiL2wpkAf11VVGO
1kAutpn7aNzDIBq8kexYlE9ikU9Pfpv3CGvuu0kJFL1GF7UWqR3Yxkaqjt6tKKKl
XtUWm6gs4jSgPQdSrMyGVGaNDiDy7z+vIfkp0I2YWzWXoRlZcS6QkgoYUDRvPvvX
rI3Krq1V0rcnnCi4yZtUFE51phrPRFN3IKNxFl3wkwZnqlXTO2fHeUaLK7hRd44T
rivEmUR0vSK4cjyhmVJGVSXRLiil7o1EzZ040JdjSkfzHOu5fA0q/3Dgk/iqshx8
/6f7Xla2aSOLIkPcGWMt9CNA6CFV5L8y3f5uOml3yy5WLcol6rKrM/0mhJcertYd
EJHStDEeQr93VsBw0CZmfCK2zEkVeR7vyLTYZYHVYBuYgBi1J7vR54zoCyCvxyqk
dlqNiu+7k7XrJKXj/EI5kwy/syMzdz7OP5P2LFLgPHVHuOZWgoZpuZtXwddtGsBw
r5muXH+PxDgT15lGritgrd7PKfK17qPfBKN0yaw8+HB3mVGIPL3qU8VDKy5PMYCl
AdSU8680Y8w8NCjoEeOskOWz+uV1IYUZT2tMg8h4U7/ey/3CdgqOX12uUPe5mocq
PC9/xvQo5KG2Le4tp70yucxSvlQiM0czS4Ujc8mjPDkpfVZaBYdfHE3aJ9vuFb4n
nDbuTXpNmayTfVxMxDgXk6n7Cwgr3GoakRfORkBhOHQGTiR1Wnhr4WKoi9NGh0cM
Ur14yPMUgpb3KqHHRJbl9WG9SdGz5fADq50cOnscMnb0nkx4NvDW6mApyUCS8kKD
u0oSqGJo4c5YAkBm+zqjJV3GADzSMXpas5ZzOprlAjrInlhHWhhx5hOMHzZVvsDa
IazFMMce2HZ+vA8DNdBedIGQ1c3dHfBkCVPyPac9D8l4AibxorvA8htaI5w9eVFF
35QWq/BqcBiH8LTGXaHRSSIIid6/mMdJSGwjCFxwsV9h5bFtUR8l19dp5muz2QU/
xaaWzfhUi9RdzXhMy4H2IAYTswN3MdRfYSwfEgfWYmCiRZ07bEFWSsxnacyFrMLw
e1b67Kjnq2kre5BCYKDn8MPbm4YLhnZ97LmLOxyBVqjMSKhe+nNGdyPsxvlyXNob
W8EwGRNERkOoK7ygiKRZxDYesAXBpUX0BiLN15N/77oTUAA7KeCFWNXqYWCSGpRw
KEyc7p5b3xXSlcPFsp42e3rTOfsUEAU8Ebmn4Pj9sXBefM48sUItfyD05LDpJs7J
Cn1J/f8grFxJpS3toH3TWXcnAc9Kywx2EjLAq5cnpixPfba0MKwdziNzHzW0cIjY
8Eb5bxOWABRT4ZyjzdoB4Zm7BDSVmSONskBwAWASLgsFACvROMy+KBDmBPq8Ir7C
CVvcEKNtTo8TA5IXeb/oBXDoox2rmgqdlpy4vDQK/Y8pBbtQ3JJohnelVj7IVcE0
AE9cq5Bry7BIVbfcB5dxttM5yRG5dkI85w6vRryf0W08FGF0X5RO4O/NEPs7Mapn
3D8oWHo/JxTGIJu5jtF/uY/9uZvOr9jCeAESUa8t0onN86oEKS1PPpaRvh8pMXKE
BSAArK/wvalpEpLlcNHwGb713h3aIpJpl4OmEcstLgXdgggrjJSQnmP4Ly2pEhdI
P9iUQlOjCFsma70m12A2QrqWk/EhoPZhLzkJfA71IqIMeVIuiuhA37QglOFMm1Wp
vR3WyapEoadms6rWbh79TQL0jtPMirtwha2LULGh6ZPU82SWaDaNS2awskt7rMan
EZtkfhm6bdGbPg5ge6C0GkFyGrxsn3Xm83th2kbjlmr5IUA0qrf1EzSLPIknOiSi
JQ3PMyImQH3ct158W43Mq7yH3cHKsBZSqj+Q+gj698wfoQOg5C2EZi7fJZZeRYpd
IAAocUJe+ZNePpsuwkXRW0b2k8uFaT50CBJr3tDcefSZf8Rp39hDnkrK7PCSrTW7
tXDF4M6GaBzkiZfF0mSvosF+kABJQT5v68lqh0NRW3Emqu50ZBcO13f2V+/wFCA3
zGDgwL54o9CC9GdE7PdGjnbA3dWwX/bqTtD3gRgfgK/J/tAEOU6CpGQT4rdh2QrO
lUKwRTDtn0bxugNBLqD37QbqI4D4lHMnwsGZx5z8gL8jL72sk9O6UT3XqdT/JeIx
7ARHD+H+PowGny76HxLLqkriEh2szuEFRKz/4E+Wpr2H97On58R4itJPVY8055j+
lA+CdaWBLUlxJKE4GZwaOa91PGjz4k+nrem3TgzK4+vGvgx0lhAraDezcFh1pmux
8DuobSWF0sg7rs+7W9wEinAJpqO8NU5mFLEr2RE0sO9UOA5Q6Rukf+hOFsdU+0Vg
tH9m27SLfJXjcoSBUPmWgU62LM5a0912ga8wINBOE5bdejnjcJXzll6dTUm7Q8wv
FcvJwa8XsY3bcQWjlcwtwq1vcbeepMiKX4erSgkzVYj8H9D1zvQ9JL9rD6712I4U
A6ojXxBSWY4/LMNXQdGELDlLtr4f0t4y+02pelzWyaXYwkafsGZLHHvtVDZB3aDk
cHbne7zv8y+YnGK0bWb0F1N4YdhGSizrEn9dHSrcfvKHMvR2435bE0GGSHUJG+LY
mSdH+NBEXJWs9H/460DJFnbilnx16rY6JbyafyPQgKGcc2r9vo3lfIoPViLNYA1a
1TfyOQFkwbG0T672ad605Y82XSrRH3i95FOoEDWxJCbEb1fimnSMyVXem+/pBQEu
YgGl0CT2vXhb8IaKHj8skCrO4zCJQRtchm4ZxuqSuyFM/8A2D9dpJVYohMQlVMrt
R0e726aP7DK0kO50VNGTAtvyPfAyqLVqckWKOSKAsxSvq3c7P6rt99osbgFPyHYG
/i+uAtRBA80IH9vyZwEcT9nQ98AIJaAgtIIaUmFS793+lPlkk3CJVVOAG5eJMDTC
HkGPpxRYSPLVK9Xry0vq6nLGYyZQeiUwgetX4R40fGak4VuQFImqRrMqebAQJMJ2
TvAWoMR98TIFrNWgQpTbEPeFykow3BlOF0NFVaqylrL/fTtmGJJax8Nn/mK35sQn
gFtyR5qe472z0VpOx9aog5H5SH81IFxPY8B06/5gBI/b5BgZT0NnTPrpNV161FDm
m1uYDAurK8H2/WUOlUQide3N438IOFwhEii/Exacv+1icLjgU/er6l0dMFTOIz4A
nLwXN6P+B2DigLnGxuQ5nX4n9C6PyMwZQKKiZyc1HcOUiRNMhV+bCaJBHP7twi5T
E09W4NMXpyaRcxtIeFQ+7z+2MqPbLoQXtRx2GKX68yCHSr9SNOKmcMRNsb+WxLo3
tYrN2/ZB5sN4bbL1yRvEBh0T2m9TTT8jvobV+f+MqooG9gFZXtaiS0ihkd26Mcmw
YubdJKImNgt0bJ9kk0asvbzBZ3F2+Eav3KQVBwwknZTxi+HJz/p682uPdriUj+dj
s5c41hsTSRy/5bLjWy+CzZda/qPyGJWeas/hD4hJXU8ePhPByf7nWPdOIgLpqXbf
8twMe82DdyCbcCSjh623iNF3j0NwiBza3WDZqYh5ZvoYiZFDkzpDHc8wRJHomBEi
qOFRA0oQ2Eq+9RRk6m2iAcWrzkg4rXd8YOcMNf5YUfA=
`protect END_PROTECTED
