`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IrCeMly7u8QRnV4l2GOBqvIBKyLfQUXQb7D6Pyn34lwqr5IOwlX4AzKZxoUFmREj
G9Do0zzmTr6oarkB+bdJrZjtQ+Pu4nKFynDOCXwf1F1ltC49XjtN98nffCffrFV/
UHaDZEC0+/pZk7C/WiHz7JOcFvNgsT93QsPTc7cc3BrkUV4kMTckH+cBFRiZ0RRx
zhwMY5fo22AJ1MaTcGcgZOAxNr8qZwAm/i/AqNF3C7dEfZZCDtIpl/DtUVWwsOaw
NFKFYnCFZXeKHtI2X+0TWlcFXjk+Xd/B1EyDSt4UsYefwCzwjxw7F3YV/ze7QhJV
zfzRICkeSYOB85+l+XJUaQRnxmFKSHtTM5SMjG018gDV6YgsiG1M4mQQ1nDL05Q+
m1HeGI/FfcRV1UmGbc2DOw6if12dvFLxonP/+Uyp3u3qNL51eizkJQwVMNiz8aq3
84DzyuxSusrR+7pCo7Ho25BA406oCaW2cskt9mBr6cgAjmvLERrybJ9JOx4kjnXx
vF/PlZgQLFrh/jBXf44XH3gUNySB60DQ4BKzrivAj/NIfvalmiswwAMU83dAXFZJ
Tvuf1T7Mu8ey7N0KGiHStkf46P6v48OP5DtjHdLndnlFiRESk6r5wzQb/0jIPR3s
fC6W3xUj+EERpMzkT9aNz2RKX3xy94S9ZH+uZvwiiS8VZ1tuLtnajG0LQHK2KMoR
KOz+jq2orJhilqDZA6dqzcgb6x/iMJCyyWOosHUliiiQmka/baV0CO938Q/Ul+/y
aa/0q7ensVcpj+metOUuhm62PxcZ+wzFNv3/b4uf6CS8LWXxMzR56J7nqw9os+0R
F093SuDJAEPwoWgWHIwEreph8GNYgDwHjQfTgU4PPMM=
`protect END_PROTECTED
