`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZYe0ZT2PPhyKmHZgWvpP03TqTibGofUsCxtwpAd8p10xgEWbjXmFaqYdBNCfOtmK
VQYKSYeSgfVD+fcuMonw3xZSN53B6MRPJsHFauq8KNRn8fs6bhuKQElqezPqJnwg
p1NpmiEjoddFoxePtl5wivlDUBenZQ9ujOkzcYjTMU5tKpMdP3Z8NGz02Kcn2TSS
G3cSZILfXQC9v4DZKyu8fp1FpMipWjRIoUi+8k7yp3cMDNi2NcPbASkfiWDnbB6H
iNWIUNjNdBt/F635VArvHXVVWOg9uTaoDskpIcuMUXJkIv5mh+F+bX1F3eFcY+F8
AaUYFqTBFa6ZI0OU4WHD/vseORSkEDCFCcRZ6ngGJ6jClZaIk5n7Bd11+w5J1z+A
AOXOQIaSXxQ23nz5om+9f5yaHH8k0CU9ucaNR+TQ/yHeTcPzbj6Rhru7613mTY6V
nWLFdPe86Q/jJDkwDKF6fLeRXT8tTmS1oW6XS9Ya9V+bfhkDok05r3JM5U0lrB3b
CvIlbKVvl1E0KDolS3dJ6Ax4q4aKyEv4P92Shso0yrgxMmBnnAcUJW3Xbpgp7RXF
Qu0jZ1AGYOOvCP85th5MsmpU4uqIaCFvCWM5THcafc5n1bIGkNJcKptLxYONMBeX
hgT9//N69aXBq3WgS/WYrQ==
`protect END_PROTECTED
