`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6kloFx+Ijdkb3co3kPsQKzZtx6Lk00YHOJ/Qan76EzGQnFjs/InFq1SfKOHL1wyu
mnalSMnjmuV3/EvmCR23bqXGLQQmrJtuDqHahFNB99C0ZghMYzIRIQGVV7+IGYCd
h3IfnmIMr5ZTxEfEoZygQeq6CAORE9f0sjw4p4Yr9Zxi1FwfzKwo/EWIMdC9lHOI
7C1sqNQC7yairJVeFFjjhhvc6bEk0W6uKvhw3shWozLJVzWWwJxCmYDT4tACemMT
EqO/ODODxDZfs3/rd3Sr4Y77H5PkKbEdaZ9RUHSY4CFfd04PvAq8vEuBRHo6fe3W
8ZorgY1mO5eOJJpHdZz2KVsvDugLdlkfXkWmHCFWUSMS9hinp7B7i6lW8Oh0lBF0
tymJvmqhvVloxJxyo5nZBPniTXFobGTIZJIt03LFSnj6acYY5+e1+vM0uaZ1tLnu
co4Y6xwmZovTmon4yKPq/DHB7dWTfCtzcT8+o2EMd9Kbo5bewk2nszGXoV6h05q9
xJYWulR5v45eM6+EQiX2NmtunnMABMYMeKQkiM5/HP7t5fGY003kCvvfIG90gdQC
lgIv1f+QnFm2fkbdAkhjZBfm6z5nejio4UYJfmvsK/xVVaHlPnVHfftrBbHFprJf
yAOkOZzXa048AFZHvwufQsqEYNu1DXx61K0+2aT0GftBC/BB+S/7TtGNgy0tX4B3
0lp2ndFAep6eqGrSPUfncg==
`protect END_PROTECTED
