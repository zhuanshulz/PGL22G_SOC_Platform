`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1Z4WAn38TbR4HT01h6ty4d+N0m16LXgh51DRQ9upghpunh6RU5kNMEpSduUcQb1A
8ooftk4ktCK57ifQ+FmwMNJAPBvSua/PVnoTnFzp6ZAiB9oEEoL5JqZYjMFkNP1f
Xh7dCUrfQzhSqjIlVM55ZR6QXm+Moiga/81MEf7WJMFAsGK0F5Da9wGDJ/j6B6/b
mXit0mkHvKRQ4l9hM1/7VuTz4UOf9mfqVdRd8l1hjfvoTW7bnQwsiferl0wGA9GP
s9BsSVoW9IvXtqyhw3/5R9AjrVjJjRJ0bzHdPmVc9L5fOdoIOMPzqDLA+E9eoLKP
+RJIn1rJBbPR0PgMhO1QT/0D+FAsZT3xELMzfGtd8SlLVvSmZbXdNs591VrrGaRY
qZ5BTi+5nGCfvE4lIrL7U+Snox3O3xbud9EcVhQg2XXEUOMpSR6whunaYnTvFzsJ
TK30SJkWGkLIs/j6UFsy6jCETFMU8i9x8PeSap59kqA=
`protect END_PROTECTED
