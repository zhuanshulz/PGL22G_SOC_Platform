`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6qJDo9d6Om0KOpmUl9e0tzYerxZoojKXiLMZRY5HKumbro4c5TEi0f4tScO8XBFd
kpgK05941f7tRUP31Mv9HrJnZYARFxrRE7E5yUYWrFcBAGTpygCGUH0d3sPp7/4i
DQUNzGIiyNtOyZkKtU/89kuaYTM9ByjHmRIOWCJhdBx95zNjRrOKYsZ8G7BG1KtP
xyF8YtFRqxiieo3M0owZOeGgRwkkAAbT+phi5YBirsTBKaJ54DviaA1jBJUlL+bk
dOb+SLz5nI9kDf8+kG4KxEZ5RNkhiU6E5TgkdKjNb9PUwAeu7if0X+xHy1fb/mRO
fe8MESYG62qYdzN9fHhyBcnPeacxRxpCsLhQ/jF4lmjR9Bg5i1tJt2j+pFYLhOxI
qgQJEbEmviEOXJFAwDmyK2BJOrL3IblRQkHlA3J4EVq1jwaTRTkySM7A4JB8qg3E
TOsrirRm+4TSirG9iv1sg+scKKzAvQtq53dz/o+QShnFMp1865+sIBHy0FBnkgwt
E58d4YTEX+P2YRtjzYn1SnuAaaYAUVdKk8WHiUbhNJucLc9pGOxMcWmz49ht6l9v
m/NtqEv3PzqaADG6xPZuHLs/YTKU8ZjqIL3yeGGVcVVPT4zmhOwNPL/0GKz/KbOi
05D0WtithGlK4M23N8AdD27OMdqVRevDg6aXiBFrPYSR+IuHOUgJXvXsOB173llZ
q+lL+9L8DIREoPB9etdYpmJHUeToj0F5feeMLCrYmaS67eLrF0Psz+I/i9QQetlr
LIMnxEYdl8fi5NTNMi5QNjC53DqCXcgq09ZSAz5R0Vk0TpPcERkWy6ioUTCGTA6t
JmrgiAaMYqm6tBHKS5yiqhnlywBGupxXVBE11VpQmG4+RCACflx/ze4ySVBY5z5F
f5SfdX51jeoDS+iBvuNyIZ3Omrz6P9fHEnPGaC9YH69FxF5UQbpiwmY+ROzpG8eT
/LlE7wSOFkXIUYjgE7LqOEqyZNqiaTd5NOBjbTRo6t3Vn1TdTvr+wwG25TTJHOIJ
uH6AXD9tMqGhy0rBIEXABj3sN5oOp75MBnq8Co19gkylXbIsD/mWYGlBtVy4S12f
EDz5jeJnbf+cCNqtxRO/0EtWdiqdbMBEsP4Rydt3nxeLWS0agCkcp119y8BsluCB
nKxALVytPA4CFWnbNEY0arLM9yRnJfRKaG/B7ibbzedPecrc0+t2UbpyqO9kXLiL
L3dxliLb0Ted3SFYjOVMlaZ5M+zI/0KRHFQbp1iU7uEcQiqIVWf3haGG9Szce5cy
T+JyeSlAEdeOcBkb5FpQManQxKPlkHs/HtI9jFbXXkruMiIzQR7U5fGHsUIxBPC4
dT5GfGQ8FxKmvqTpLmvj1n5qgHrPZ2nboRxnHpl8NShtQ6WZsKn6croXYSvDVW2j
aiBkYwTO4WhYrLyUF/fILPtdUrN/ejBcQHq9RLlDhZLfZXNeyoZxHjlDfMJ3810A
jc59RBM5ClgP+2xnIaMkHiJuTBgQHe58rUKkCwggn/QI4jhlxX4yVjVQX6KIqicw
eWmGxJ2CgPtr2+tAAacb1tyM/QpJEJs4yH+dfyURje7RyQqhJv/1mz6DR2fOKQR1
T2a3NHR0Zu0WkKCobVnNiLmxq9LhNbfe2BRU8rxDDFm4zbTDE65DdiDlfgLKSG9W
9+ZfaChhEGVWfFbOh1m1TeHQWQQtjDnW/e+mxvgC8frcXvnLSntzCI36qF2cU87b
j+1yA1VPb8scHijEcg3Ng0rO6nGxx5IlEKBleKZwWwQKVbS9TmDFLVK0M2AGxClQ
9l+XGmh5lSqtpIiRPvw6QlAIzoI1bHUYYIHvihO759tXnFR0K/Umb6yPryMURI5P
NYku7TuGh3xCj/kzAnPlcB+P+1ako/gGIrFNE/7VFJngRf6JvWkWAb+ROflJzs+p
PyGI7zR3g1wCGxsjPag7Hf7o4vzViDdNWaOKuapJPvjzDitkuNNOAfRRRUrSqf/7
8fT8a7yUDJFmH/B/5LodHlGq9yk6ATe8qc3Nv7VXddpTdHdPoiT7c23kROMmsPF5
pl6QrB3kb18lHsL/YsYwIrpnBTz4knmzSe83AJMZRCxqyqm6j/GE9NBHdXIfqirw
WUXVWu0ot0DqL9dFv0B0E1D8Fq1gFsVzXsJ2mO7ov93BILoOuHGPubxY0oKnOSvd
8dJGrBDAiupHv1CG5XLI+aXZKMlYeYzeK7ERa6PgbI3oFyv9ES1JwSKwD1phDMXn
sRUyLP08y4JFUWwzpofwc3TK1AXfMPcLmAwVYUWFPevpaGi2B5pUlMII/V8lBU+1
zYZ2Cs6KfJuKHu4G/inP01wGc/9+Rtwrl/j96zLbu1ZOPCX9w8Y95CfmqSELiUSK
e+20TdBjewEpThMDNg01qeftj4O1baqwDOe/eaZZBrybn6LBdj1vB910VQPHQcCw
0X9hTGpTuv45NrDIwCLlQSolGqDERHhNqLNJHH1wRiAXdoX285Ra+b/6xDBXHNaY
Wm7+1jArvxJwui3Bx1oF1EY57uhXcRxvtqfiLytPboSSAH7uvhWFdMiqJrrlDNwj
hPHrH3EjoOWF83f/2c3F+FlHUsDtFvJSx+36/39rhxdNbPiDaD++c7fEFEpn/BLZ
zK0n9qgCnIG0Y2ZuWCThR8H3AXoWfDywTHoVmGZC0sGZtLbnZjBmKafDGF1dMIgl
MjXEBK6sDQDTzp7FzNEJ64v/tES4kS2NVVMqJditVyYDAoE+J6ODG7V0Y52wjTH/
1Jh0WdjbR4HjUpYtZTlNlU8ygY26OkQ/VjrohbvdI02Z37nCudPCQ+8T19TLBRnI
wcB6ve4tnBKcyQGrNner0l4Ss9wfytdrvLul+tCr8uB3D6d8oozbzu07MJWSVddx
ZITwbgSi36dwoaYOX3w7AsxP7x0Sfjk0UY7XuihC3B3/ZuZO+pkLuyPVUHrMgq/5
EApt2Ma4dPge6FDYRip0Ls5coZk+5RjXA6Bw8ZQGMfeVRZn7D3l2Sg0vbOCzZIzt
vWpO0g+0f0wwS/34aa/4fLnpAzw5ewHDuBFoEQxj1ewLEwO0zzBlzJPoHEoJcoom
PMyDrVHV5mZHzwesMhLdiWPwbk3/B0N4OEHA3VxRoGf+W3zd0k07wSAempmSmoqN
97ZyOKXqSi0vo+kD80jiNx4lmxiZT1vMurz71TrVahRmUoGwC4ZunWqgkurXFfHt
2peZxYH6S+LpFuWXPhWBvome+f7pdt9kZDzPh18iULf5I0lpwKtrfni/+CgeRv4v
0b63jDG3xu2ieQRpfzMaUeIBdK/oTXwK8KMMnA2QtVlkYS5eoUnj9/rJEGc5Z6GS
7XUdNPKHsrOblnjV6wd998vH8lKw2wNQKaWBuZ/90wQwk6rRJXktI4pCBnFSKyUf
c3lsIprL8QT+WjGgsbkoP/E4u3UpcXMIwdfKAipXeowVanqdpH9uefsAxIsCV9uj
G0jYGH2m+7sNIXNdF++PFYuQT8fDsidnWAU0/c4F2ycU6P/URd1UcAbSpxkQCRoZ
mBW0ASDwvS5DG5OOcVamo7mpY4lU5IkGjo9HmP8ggVTVuog2X/Pa9sKxPUw/retx
P8eR5w7hgA1OcnuKdK59NiDdST+sSWT8JMPZJPF81zyr0znOsK9AqXmwx13tvbas
TQ+BWSHXqyulB/b1L4svNUppNfu9UZOkpu7oq1AgLo2R6mIqIJLigYyyHb+rlCua
X6lBcwki8kkJrHX6ZBz9mkp4cqCGnjL1YODcmbw/vlfJX5tEFbrReXe+lggTM0iK
vAlFT8K46GRWmnJ54JB+I8DPyi1IF/C7klJO5Buc0b3RSzpY9tDdH+h1LmziBy6f
MtdwtTNqL8tFcj5jfW2NJyMsyoY90c0/ZC5pYoANkMyxRFUvHZtc6YxX6ksM3XdT
KoBTHfWlxxmEadCM5C2F4mcqJx+Iuo7NfhVkuTugYDDSqvCR2Jx79OrQ2tYQ0xzb
euf/X2udLAO/0zOsrJh+suWzx4Ph9Az/8MlNGcyiX1HLIzqJGwZp9SkCt+dJY6LR
dyViS5u6r8tE3LIbPAp1rEzn/n7LpgXnxsOS3mUpvfEzSkJZIVqMUSBtL8PclZf/
YUSf2dNskd9TKpIQZWTsU1OHG/tAhdq5pyBWQHUjXeqspDTdo+oldMTiH94iHaHR
X/hiTMJBURfzsCsylEiwBUc09GdvlKSLLvU2nyzYsnbmTQ8oSkJXXp8pQYb9I30j
+eUrtOnfb+SMtDwWRGjsPJctItY9c48udtRLIkNElx82OQcT7FlEK50WyVu6+jCz
l55ejhZ3r6++Q1h+fzCAS463kMcpkjyXK7WHkrf+SErYIYvsqTyCPMRPqRGPbeou
wUIGxiJca6l1Nb0EojG5Elf8LHKpvP0uowgXbiDNZkqrNUU4UvR9Ydxgy2FNIoXt
meqL5XLlWIx4hya9ABW4g2R3RS4MY7jjHokegO6CFRZTmGnxqFQHU6DWMUghOQ7a
jC2w4yC5TqsmUfvREeHGUX464l0ov545mVNr5EUQyqB1XBb2CGaxlQM7xbT3x9jL
6VXMtvzpTg9dq8OXflSh7l72qOjKI0nnyprMbY2spxDQMHuzTZB2+WLFrq+fOrm7
xJBhl6uyJ5EJNfT+QkJvceDlv0ATcSjBykSgJgDixfE+9SVW2N0WE6B2DAAZvl93
b/h+nF+Dbgh94SMQcYdx4BK9sQ/lahEURFAYPbZ5jBSIonEhABXGb1UaDStvYfhU
J3YRYIAw8MpAErMVgJ2rt8i5YXdphIqh5/MRnpYlKqXOWIJkiuvHw7O2UazfHD5m
lDpcNfwQ7ILpZpvC24/4nhkOm2y82gf7O+T+fRQDfvH+AK8OJBPKg/CNCugKM3Is
FDY0sDY5pxpUbLC9rm2giFr6UcQtmrznMjWV/D66cedk+Z63ga/m2779jkxlEUle
J1UMT0N0RVvDRojtByGg9WyeSPyiUY3118+Z5z/Y2le+g7WNNxpB8RVCzYNlvNbl
m/X9VZbsZw4B3fHc1a8JZFfYLVSXwymmuRvpgAqpOOYdVIUXb9vZ+o328O+/E34Z
2Mt/iAXuCBEK9cX36vahBKTbEr9Wy8c0m2XcXUcUc+G+K2/WF5hruXHqiSVcALhC
olSdFrG3lcFtQui8a270KYXv2fAVESPbezoHuAyYxyF8zXE5SvgiElGsg2W7tw3G
g75qedp+i8vqyYrI2TSK5IQ1sxwTuqKtJ6LwMefkbBYFUiWTGR5Tv77RddO7arX2
WBUhDVnoj6wy59sL/rHQ9NmHm9JX29aBi4cyjeoCHmdlPgG8fzPcpHOQGpZ0C2E5
qb/bUOVBL04w/0IMpwW0XzOSF1tvjm4S4BImwv89DUpt6TEB2We83syH/LZSYP1d
fTEmZTgNrGRLoJoxk/E0kKRWCwim6x2DSg/6Jmqv4cpgLzszsnSWGqy/mAtmaRm4
PI9+PTyESt8BzejvUB5AKoedQIRQR+fzQ1xVkfQI5siEHo0Z8jlaQ1zbCCaFHm6P
x3ezWJG5cj5jj60P8hDYwQ/i8BCcQC6x5RVDjhu6XqOwoUtp/BF8jJTA9cVMtZLT
r0T0kPsUX9X52uAzaV4bhy4UpFmbIX0yb0uWOgFvEe9urX+TGFos5WwNeSwUISmq
oYGRxfamEs7MugrmAUj10j6N9Lj2Fa8ona5FyPbdBLeodbzjWjK8NZhAt37T6frQ
+zJUJXR5qa7w/3Fw1J+CIQsM4PNzoChg6yEEvpktTlzaNDPNrSbBncLi/xB1HC6E
RYltlfHgHQ2m2twkCKn9fzOVnsTuvHPfAk18+GWeV3b/1dAXihMouWUoseEj122g
YkUJtFyWv36UOlJWUbE1YoASPtCmwYEzH7TmDXKV9JauskzAjLPu6xB7YF0j0UUa
Lr5O3Url3mzN5yi36gqPni2G2J92TRSXNYHSS1JBPRg+zrVEPPpJSEv6NlR/2U83
xJaeGhySEzZUtv9BrnvToSZrzoQ4Rp0ptD+uWnhARjc/xWdPpz2oIbOGzNG3D7j0
F6TTaLFi4xjQ5ynaZW1iJYpm7LRcF5dc3KXKvZlnsxpJSSDIFW9r8YrWA+NSL1jN
hUMmZWmr/DCQ6CNeCm5+R3yDHY/UOn2QTP5t9cWpBGaimEW2ftRWcASZ/DutQEah
lTIGfGgPY6dlxiF7DdbeRa0Ri69Q9WRL9VyI1MifiFsOLc25YE3Ji8hP0+KjmQPq
UdgK/xtjN8/mep2BHBaS99fMOi3ZCf9XxVeYZsBUuplytGSqJhD5MjvwZ2NbzDpZ
5jqayMSNQlihMCHwQLsAIHSpQ7805+40rsE3A2zEflgIJJT9R8ai9DfJ3brWa6WN
B9kTW+Nj7zXCX+fcNxiidikhDlbzGQEggN+8GNP5ooS+1aXCeESVzMPk7WqTfa6I
tmgPphpRXd0m87Q/zl/xWjWrhVqlVS4H+xAqceHcZjfpAEPSsaPj3yIMWj42Z/L/
hUCyGTYaI4McrfQnB0OODEmfExIIDc6yNdH8a4F3Ix4alhJOjbHnHt4WzHcyIEtp
++h6E9uOHNUIJSS2J9yOKu0BTTR50/oPentvlxJT17MAY/E93KZPn37Yz0BaEqQt
eamfuUAc4ya2/tI7OgPjKIqIkx4QlhO8JW9ZvxMW1HuelmT2Hv+8RaoNIyRvhFtC
BZ2JS9i/DtGDqyThvWAQOqibVRyTaDkakfTtU+2xLbXAJNphj1+CSdQk4Qcozce/
Nlp0HAugNJNlkZXOiusq/UgWWES4tVeP/AVXyfWWWe25zqgtCO7XLaPg+zDpi5tm
MWX5RT32GooPnLtzDjRKwlwhGJhfAjqVp6UxAH+OIRKbl0ygbHcdbTwJiHRva2Hs
dFLJfmcEJO7nbGID58N+1aH6o23YpXsNoc0mIkjdMRMHfR5GNrFjN0j40yD1kacf
XZOJRFpXm0QRHgIdzXM8IciapYceoO6ueV4wP8N/jUbitEgoljeh/X3ZKCshdooi
ECWLVsYxWcfnT3+E+OPyOWBrv340LKIOQn/aXqD9pdrw9TdFLhF29697AIWDwBcf
orO0IYVxoGdTlAkJZ8HUdAcfV7MGzlXAu1ZyNXredj/rwhWiIR3e8gznVZzS+ZC8
qJO/xKCaJAlVxgwoKLkOwSQ8gEd/hUU0DciGOOHGhlKJzJupDNMVzUV7736Yov/o
DC+rwzcHYa5qvwWfPt3TgQOknDvQYWtxBvPDxrlsUzo83OaANYz0aP/4WMpyZHcp
gzq8P066OCMhqlJOnSU/YOBrWr1Ku9+eHi7w8hgSQdtDv9YfAsWDDtzd33+T2N2h
tD1Zp6Qg9NOm+zzBaT1gaMMyowIaZc+RB0F72xXRGXcCcm7KBuqU+Xke3+gadO7E
3xmbPTr4/iualbtJZ6+A3XaXumQXwiQVjStJm49npiPKlpqekwwcOWZcy/HC/hjC
b2IYFr+0crc7irshEZk8y2+6F2XUn1T7OwGxb6dm6Ez2AlAJYdoPH/hzrjp09uJw
w/8zu1VWAg3rYWbezn5ZC18wFKpCwkjDqArcSnIbEiS9JBw/pm5kpFAFuIHn7vrS
dZ4f/DNua6SuQAoarDrBUECyqs7sRDe+X2/rRFV6DFrKlFgzotOt55KFMl/gAikv
zFVZHus3q4ryaCBEP0ariJEvdBXnJIxw0tu9JV1C8JPhDy1lhOdW+wNPr2g+DRvT
Ct0VZW27kiDn4pBjv0SIVdVWMn/Ge00kCGhtz/C/q5jSCrwEYoc9cl5WlwbVAkFD
lGhiBXlIU1Pw6vElIa5zGzt1mXjSneVdvUjFvSsYSX7SSsagt7nOOIdXfc0fkBmd
RKS3/BkkjB7EaTHME8ABTowb80PHj0SG8JJJigesJDcw8GdhABS4RsCn91jcSmPQ
Tt1qRVWRLseJ1PGDeyh/SpCaX0bOMAs19Vwq1jL3JNGuCnh1STmmE30PrentIGGl
xaGqRG1eSeCrnzoCEWGq8WrNgF6MB8F3NrkjDgWIG8Mz7mYIY6CLtZRQMoPYdFiz
vTwOPB+5zUNNbnx/TMC8sbwg7WOEu0rfq9sr9ZKYNhwniqQ0cv9HBbFIvWgV5mbH
nFz8J/oQNySzVUB2hK0kFpivugk1o43LOolVfJPF8b/3tWW8rybp5n0AVuh0WT6+
5b4sFRBJIH/fqvifiO4WdxI0cTTUXP7xSWO5aCgIqUorcchDMThllWGCag5ZQfAP
8qd9n/jTasyLKV5BBFRn11gSjYp+U7YRITebXZP5+ruRUJ/9FU6q1Igfif/FC09Z
2wI7r0OWIlAwnXeyq2mxhNgY8Ymxa7lu63Lsxwxr1a45C0MfZ3/iVRHOZedmBtHY
DNO9AhFG3vpfg12Ek1awbx3GV5zg7jfnexF/YMsjN5DSU666bHgTZQRbYcZ4XsN/
VzrI2b3EK30qpqXIm7/+vRbHYgkNoFqqGTs6Whb3wG6q/aS7RsyIg8zqkpQMSVfh
+XNW/TiNxVuO99xo8dQgvniaeP4ieej5ACo/Y0iGZnN7TNf+28XyX7PeJ4MK3L+J
6qN6gH13f58NXacO9NjfkBFyMIGkeuIo1LqbMSsTfRYeOQHtC3qeGc6uxf+KATsa
vNuR1PdZo7tWa01rvvCa6RCS6Ox5IJ1mhwMSIGgL3XlMXpIwPu8ep3nAzjHLjsLv
FNO53NTavLejycHRT1JDrcuf4AKsC/i6h1MY/QFPH/eduvBzPnAGWMh18ZTNVm9m
Dd4NsJYXdwMUTy2aUeL9rnsWdgG5gyan9i1DZkTjUD4HkY17vsBexeDcngjz6L63
lbALnqODEcdbO0zHCOcK9gN60WdIvfJ47fycEhBxpsQrM8dQvUkVTW90IH/uwXkC
wMb1DxU6vW5o4QgEm2yC/fTxDQHOidJId8Q3sbdV06zGuLNPa5PY6JFGxUZIW0+W
iY6Carrg9LZ7FQzMYShVb5WpC7qqjvNuiH/Wjq1lTF9jakePTuTegul4G16EZO5j
VwWbPoweVC9lqCyC1P5TnbyV6YL7aZfwRq+HTSBqN9NvXop56SIid8pH98Ida9GB
z+JubSt5uNCqD+EFwZwGoV4ENiYEipkVqiq3HUsjUgP9eHZKTpOy3SwD6UrBuZJA
aaJFgyaYmfHP2COjZP+YESX5ly4jwhzl/FNRBT4cKlMhdQhxVbd2atRw/eirAUnC
tv8W3WBNboJauW3ijftGKSIX9guGdcagkjqdbbQq1hEY6Oq9R0E2hWG389Fqga7n
GEx156AmcBSjn+FrEeuEEdaMsY0502g/uo4hC3z6FbH93LwmQwH0Cfl+gsQsQW7x
aQPFj3OSSvz9MUPHz/2rH3NZe7lAq2fv/LvUg/JPc9Xvjtxsqb/BwcEs08OkTZn6
JuEqpIRlKmU6st17BdliCFyqBVGyD0bsOq1EveWMeFFkgl60eZAPyX9CPxtroONj
5cmkbJ50e7pkB8uou2s5ujG2lo8yTOfbx/ADTbN2TjzsJRcU1mHTXcKKyPQMw82I
1qiv5b121Ja8Ebm1QRTbi5D+xxqNrfsfujCPdTLIQp7gWyWWJD23MlDJWt/X1kVk
rF9e80RiSbxzzhNH7nQwhkX5hgjlgovrkjlVhLQwFvgi1JZ4tiBonIyIIUhx0c8G
hJqzaQfEIwf2IH9pIJ+TibBnGHUzsCottfOsgghOdyCfMSDmoaQMXY1iKTS//i56
AD9dTYSSGWLATTFQfAHl7Sc+tKNIBeHjk2WPpWWtksp8+R/GiTE25wOsX3UJ1PdK
6v9+rADsBN+RkDABCDxK2d7xj+OnhOrpSOT07WWN8e81j1e+0frldS2aCgvOjWHa
VymdHVWJx3bprklsTnGXvhL73+5BAEMvOrLdY3zer4AirF596nmyrp7UGn5DFl4w
pbRotIntF2hvFlO5ZSfS3mto8vNHFRb0TP6c/Rzp/GFWdm7DgdK4unUW8b68im+V
kUi4oQQOs+TaW+lO/UC2Exo0HhVIYlKMi+PpENYl1VuZHvqFsBql9Gp96WhUdkIq
b6QelqT4DbzSJ7ej2QCV7MMlXotIRPGWVqWjiDofMHW++TRQZySm1WthMs8XOgyg
0cx4QcVJeSaI8nm6evClQ2dVvCSQTosyTS11P4TJE3Q2LForZvUQbyhze//fZYfJ
kk2I5KRxjPAF4XvMOvljQ69l6IPmg3z+k4WI1gkZlDN9K5/vK9YV/iXRZ9Zi1xaH
BrzJwmB0jTxiNlVT7GvRDhLbcxnkdUujIJ1Lhfe6jxAPrJIzyaEYIQgX08u78y78
AXW400Dr99/HcOZ6OJwWbD5nUjd9p4iEyoKmIagQ2vUrOBd2A6//TIAjsTHtz96n
gk/law3MzGO2I8Nm1+NREAtnXxgA703YeavitLSe720xS9OqChOuzDuS9kjPZpAh
9H/FlEqBaoLXkvusBGIjHvLR7LL+0oyUBB1AIc0bJ9tsu7HE7KWFBOwfamJWZC9S
Lk/vptYeDlkoWQNg7RZ3IUgyDFbrDIbVpybwGC1BGzpS4yMRhPQX9EThq92LZgW1
fHY3A06bfg4qUuJwzhHJQyHw3Y+y+NDV5XmSDVshc2u89Do/OzscpBEoAm+TYElM
kttlEDhl3N646ElXY5WJ7RqLqcA7oSGQncF8xDSUdt1Z4WP7+cHdP4qmBS8O8ZJK
XnpfCGviT8Kk8YFvF/1EMPq05H6/n2SEFDjGUGVTp+ubes/eaOc0FeMgdvQiMjbn
iyHbwChYTjZaRoCpqf3NhZWbxlgVWgiU6Yfzz8Ycezl54FKsZT5ac25Z0uTrdWRL
8AryDcKMVWN4CIu+alkv99E/wWiF7uvtL0X6ssZD5lyUwVPPdL3gccuUVPygD5A6
FmySq3vYKZuBMNhX2kjBrYQG57CkcZ6UUX3sUMiVCvWyWm8MND14YizEEQxPqIoE
WfZOdugUudoGyodYv26jNp4Qt10l5xZ02/iJmAuCgf384D7QMVFCkPmHHP8yAi1/
CuPu1ox89ohRedZuPC6n1TvaHJ1UHkGJNax0rHTnIh9bWXUDE4M+K0E2YNZt4o1U
70Uz5ujEz2BNhgycZGS5P6gq/zafZjj/N3bYDIEtqSKhxZsy2vWjspjGP1kIH6ZY
StwJBfgfH2lWrB+hTzLK7MMw4c+9hc3ZXlcaY4w9E3stW1trLCI3m68ao05GPIrN
P8XOpDZ+tXKtNfmCmPqexuPd7as12YdWq6isEhNxOfwXstp+usiU6l3WL0iqnX5G
THG+eRR/7ghv2wkmpWAGOcnhdbBJMwNSyyqK5uDnUTljD6UGVmGFoNkBvAHBMYFq
1uB3VUFNGenP1dXxKmtJ6yRVkKx8160oII3rxU8wsbm0Ados7T7e3Et3mj/T/ojY
id+/RmIYtecVcqqc0t9a9lNfGal8ZV+OvRSjGU90wbwRzNDS8g+bhUZQJ2y1OjAU
yzHVM8stJZmEP83xrOA/orMPvvMP1QRjLxYzaZLefXCpa1WMsOXH7t9AAHibpEyr
MdG3R7dirEFKMMp8H/mkgvcNXBMlGT+702UQAcsiB9G/leJDa+AwfWBVpuEau4ox
ll/GHiavPtBu5IICdr1b/92xtpf6Fitq2hrZtpdCfeEA0vP/VoSU6FTU6E4LgYBw
gCHJMAKBUwjYHTpY1Uae6SYSmSHi5XyaQQoGVAgnd7/ARTkk4Oi/Ip/lNyg7gqzi
9WUQMHRvyPOEHdmT9GjV0QAFR9PVmGC50NR3a1lL10H8VvxCSP0GbqwezOpNMca+
ShADAN59sv4IOMBZECo4GCLjDn5QmFftLJQ6Q+U49RH2dXLnB6z8t291RzTqcpUC
jyKL1WOBXA8n9PcxhG6UVaxw7VI3h7nb10fA8jh3HAOjUUG7rNlVu2aGPIe89SaI
+3fKE3GHSR/Nhu+4qvDg+/FjsB49q3gfgZZPkPtQhqkLJVsje5juMs9l7y2dWkZ0
HPNVmErFDTB3Z8QtEJBocP0hKdOZs+6v97qxUouumz2NE9pfdQ+1mpGpkjLtf/X+
8UAspaMgu+8uCJQjn1FYybv6SyKomsTtZnaFd8oegFLk5mEls5qZkk72kx264Ubp
3z81NYjy1l5x82xIaYzBscrk8ZyKDCQ1Y6fXfqeGwT1FPwEVUJ7uPZ67gSSK4C55
v73O8+5xxe/Of11P5mkfZBDu13WBPIZ+xJxgYpFbU1/v5GIUNoj4cSqviIDiVPZr
WgFJfdOeROBvow6THq7JJYFsnB0D8Bu5v4mdE5Ymfp4EPw4tEQuLS1IClCLQdcRA
8KFm7f+r6nvGYuBQ4byn4KZchf5hT/iKj8RmWpRAGqcGIg+gPYasffPR0ZmbBzyF
DMV8LUadTq/heVj/JzRn7AaqNUQd7E5ypklxn3vnzJvuuvbnL2cP5+Z0QMG7ieuv
D2KPxv5tol/Lmwp9SqX64Zl/9OfiH0vtzUQT/2in2gpti/oJNopDGOdC1R0F3L1M
GC+3CY2Q+9NDQJxUtARcrQutSt0fZudUUfhP5dG6KJB3zQAdJ+uEfa9WhR4/V4Ft
phIrX38VvAH5lUzPSghtIYu4GH4GnINNYsZX1vOBPvq5khSUoN7Dvd/Ifqul5onc
+Gzn/RWTGv3O2X05CaVWd9s34hgurUaT3exu5ydRdqbU0eqSpWvEK9XZI/pMzB2b
bUKH7aLhYT53KZ5VAgtDEBKn9hI3GUoYi+CojlFa/MZASD/laLVb5LNGXCOOWZ8X
s4qmVAYPgcXvhWKRs5c+gL3/4UvKRt7BfC5BRwPNboI/nHLn5YlUJ26S3H94cF1J
T6RWiy67ID/zfQ6U0cPQF1ft+TEFlmbTxIn9B1i5CKZRXSQq263AYrnts7YsQR9O
VapaG3OflQ+cyLAhJCRTw2wDweJgmjYM8TrvjXPtwGC6i0Q2j6jDDUXcT/9vTxhs
euGQQrjmHw6c+pvZ0fsd6lxX8fJAGTWjHlIoAc++CMr+C+FSumuoM1DhM2iNQZAg
4yH7J6XxrUrVxEbq3iufMKHdlwKdFtsEMxlpqUdMf/OrT4oHGuCCgxt/IJZBRzpY
adopr1Dg/Z+HiINk2KVG4wyJb2+hgmAAVFDK43aGc93cZpS107j59TI9DjudlmnR
rCTEdSmpyK7Bb4YTgL4MRPnRwNcBt09NxurulQ59pCZM4h1V0OIpWmopVhYtJPnP
6qi4twHf6k5+VtYB/SXPEsgrdX/j/XrobAtRXhKD+yWi5Dc/tDkTyDHVSXRPFRr/
/IybgLYI2kp/InJPAobcMS9tHGMXNd2DGHrsAiwFMYMm84d1Uch6GkX3CuvAB7EA
PMQZ3PrkzMdMlASoQnhULcZTfoy4niUBC9PuVM5TbSXdikRQeK8tqcG5gK5lhoS1
r82iPleqqnGz0U42n+HxlE+hy/Jf4haAFXWqL/yDD1xqDe6uP7mwqWaEdHZ3Avad
FZHd4QdQe+IFDhX1pASsdPXWGHInb4NF1Bet+gMJ+mOcS6sDX/04KlNq+vA4gFEh
TskCMo/EzPQ7lpPy7JIKHN/NNfv+oTnFO5nVum83NSVA1TMMBIua+5z96QrQsE5y
lJpwa6AYZxRuQqXhonQC/v3UBu+XplypPQjJi89wP2IjH3V3HnURkC+NGHWRZYbd
SHoiu/5QQcOL3Pjwtw070UrdX2XMqnhTPG7HyMDqb10qkQVqgy3tr/E3mTWb7xrj
7KxT4ckGz0yiQzn7sv2kVPgwaw10aYg8q+Q+y//nbmCCMXukuWleAGc+dnZyi+d2
rG/XhEkf9iMv/+E50gjEC9QD3f5613FJOw5DALfazb8UDG8fEh4yMALDrr8fCjLr
/QaEdCIX55WADECG2fkRiWU4+bei0yph3Z6FcosxNcZ4JcWMEbYzyENScOgdACZ8
ygzs84SCw1tMZN1ck/oewscdiNBQT1KrtM6Zd7mZ+xtuB1nUNInm726VSAToFxtP
RNHQDvMNK/BbRq5+zLmO6RdL+5Ocwp1fJ4a/hpOQRo6SdnJZTqV2RqjtrqYEfozg
mxXgNyU84QYs25iDCXAFJo6lqsUbfnDcEsf9LQTTQrN3NkL9x554+Wjy1idom+a9
kNhgl+O68vMTcWB2KfL8qaFqWGkzlGj8zYISrhprR4O3R0KjbD1IElpsSSjkzwLU
c4vCA0qRcahd0aKx+SdxUaEJ7S70lDRANRHkFLSkGo2cEhbIIHBxhvsm+VluXYPi
DKJLt5cCjVUuCXH1IOKpVRMjZVkSu7gB+esI/EAZ+xp5+IdqqFEc0jwsfFf7rujb
SDG24ljKA/uBGgx+FxKHEnNDUxMZRpTirQHc9lS8wFXJtMgX2dHBwd35rEPA8Kuz
L5m2OwTUYq0Rt5IUrYvtP9w2Ti3hzIs8kz9SzJe9b9g5OY22J7Y4PhVfaoZGF8x9
6VcHvMLGvkUtsQCBU6lxLpYHgW7JUbbOEM9BJ3qgX14esK5Np0rO0T25WaPxUafD
NzD0MjMRR9MP7gNHCklTzBgQYMGsIhLWr2onX7hVTC1pL7eAyyTgMgNcePrTOo56
yaEfvska8+UpKL4w6BBnyJYO//+xQvmmag6VVW7JegI=
`protect END_PROTECTED
