`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MqPoyU3fjB24rUgOvxFG+Po3pRdnfYUI5vz5+3snjZImO2bzkfPNBLPvqLXYkt8/
QmRjKjZU83Wc6SRbQHQjSVK9a2GhO0UjRyzjIe+1+nhTVu3LiwGOA9q6Bh/lajSG
4YxwyMeu6jrEGP0SQ5kkyuVfERGiu959XSvqZaUL2Ed2QraPgZp0V8h5jKTvV04I
AyAwG4Xnj0HEHiVsdQcbJC7IeqAsC9ta0xdFaMBlueBXkuBVvRYEiUihibv5IKzF
gpADl0c04w3/VmUUA3FU4BoU3/ScqUW2oPcf7tmBli3ccTr2kmx4g72YV1B9XczS
H0Gyr3/V2EELkn0i6S8otr2j1KVejDz1LAoaENlTQ03miRSy+nCexRhDYH+TclFG
He1ESKMbaRTGQ+wemFBaRR5T9tsy66udpJ8rz13LeA+2qqK2E6YxrGgS76o/gTA7
JhYm8aQ3Fwy3Fr+YZV0kBa2Ng/1s4Vw2D+I5ka4ftSv7wGt8PgIANg1J7T2s81+I
srE3LnYYP9bRFR963dOTzAl+uGDMnAx/sUH/adFM5aUzCypoMyxzzhMPf2Mlj5tb
ovEFXsAmqVqmynmWpALFRALwGxBZwk8mkfzl7GwSLeYEjAplrdMNfB5IeDWF5MBt
fS3QnqFLg4siC81Rlcqnaii5twM7vlYWNCuS98SIrgNEkPG7kPKqPUIBIzaoLKep
y/K3po4qNKYlQ3rRmps0CCB6p599snYynx8rO7sSiywym/jpSIJ09CwW3F6N+5ot
xu6dt2aMDRug2+2cmU37kK3UgNXj5egHC38KTgxieZqgEMNTmivWQZqGi0C2ed5F
AEuiWaxaN9/o55TX/il08wi9lmyYMlz5mrBhn/R67TVHBG5UdVueTewmSk032ncT
b6aAP1q3wzOx5S0HQK0R2rF8jO9y3rMbsj3vvaz1l2yhpH3tHaWevkxCHdCVVRHp
VDCFxV1bvZHmqBan/0jV0rxCYbMb0Q1TnH4hSYRmqaWRNghIOVJrD38jN5ZKcdCX
wl5fwdxbdtY1g8z+AH3DEFpzaWMFLmxqwm58B1eDRt1hCdQvZGx1IS7D7kvEjzx5
1LSsd4Eul0ipOfmEY+2Z8prlDjF/3gB7EfD9kI5dKdjZnps1xSkhnAVHPoUp3B0q
FpEQymZ+RMB9gdTiBOxrtrPhh95sVk3g1VvXd0gQBP4VNmReAhEGC8ayz3OON1Wi
QNiRTrbpr2DOco0KevQk3CgD7+vNbRH5j0oaJmn4ytgCxa47usF0/o0KAevGRkw2
oFyt7PEcltTivVHYzp9ksDGnxqdxdVWg+eGQ2W1X0i9wbTmLJmkQpMk2KVJKpgSf
QeUnktEq+d1Cpj1mBiVZ3haFqx3v3edCXa0h3j1J678=
`protect END_PROTECTED
