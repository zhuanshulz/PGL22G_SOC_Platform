`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tXmDpzgRo3wXBl+vQ5/aUmh9WokpDCXpZPpiqBsfmPOk08RHxMkmHQCTz5N7N4Vp
LHZd+QJBMVQVb7ylSCGJpHjKTAGvDLI1ISX/VsQEvLXhecKkVIhvf9i3ssB74Tgw
3bEDpHETWnQBEANMbZFw009Vp/KCe0hrxl5sMN1Il7hHpc7EmoMHkCF8+Fl5FKP8
lsV/SQZq3VK5oJ7ORqCz4/6+BbfDNMiq0S/BadANmMH/krt0dbhFHwGtUAQqJ+Qf
hE6OKaoiV0ZmjPdXzm9j4kpI8HkCs/b+5mFjnUubdWUiEG0IA05RZ1A4ixbFKvSh
roPsqH5MhEcmtcyfrKFpvlsHR9S/MYrodcBrO1SY89quudywALJK8Bous9mRvMGO
EcvhIuIOWjphlcRobf8BPOU+gGb6Qucqrj+ZMeFFhrlhYEAmV/hqBn/N+4jYIowz
CC78BAJI0twDK7dnjBaRissodHcK1fUON2kDmxHtrsYcPEKHFEVAxCx96CDi3aNB
JwhLQ64tW7LuPEHarU3aICrcFTNXRfMwd7MzURPZ3CA9uclEZymKTX8sNYPUOghy
Y51m+3LgaXB91e6Ss2oev9E/SIXsQm6m/xOUyT5/jvlEH2aDWQg4AU+EdLFlVgsn
hhGcRYj6GbaLE+/Wu1shbsQmIIs6bU3HgczWguiobIMITd+6Zf9zcCm/kuU7/ACn
opKuTQ2UMwNVfhaA9bHMiTMFEdlKKtIDqPyAfhzhO3A8XkenZsDvnLnJ4IDpvCyO
OI9x+LEIn0t48JV2IXMHukA5KHXFRp0fn7RWbKS6+98fv73RpRF2GT9CIBqcianA
q4UBCanJ8JskDkgyl7OHPkFakDgX2NMvPMbrZ1EW7zROHZ6OgcBeFuCGRlqNgvvQ
w+3LRWq0ucgrg9ovVvwu1B74gJjE1ceoLGuHoP1oH3nPyY4N4LuNfcVQsMuSBPDd
xkVX6KTDg1XLasISCFiJKmANGzwR4BjXlKcxM2Q/c+bXQRKgIkp9FOgfzbH5+pHT
+bTQnIaXNLwNKpxU06t+i/n2x+jMm/IEEihbrtVb0/JYA/QzbQbCTaHxvqEYm9Wb
LksTO3IqQ8CAJTQOsQ9rMMDdayGYNA0jiXQJUQr2+1bvj6i/aVXT/zAvS5I4+U4g
14gw9Egt46STf5OBoYg1CzpVAh9mgQllYjq3/HxNGUg/X2malcLTKZEjK1DohekU
jMAB6lhS1J0BhGYUFBmEMgEQOxKX1K6NDm0ED8DOyrX0P5fyKHPQjwu4e9iqc4YR
Gnmy/ma9gXFFD3+PP6CjS7DMrB9Qq2J7UVgXJueKhJ2u9piwVhJ479hT2eLg/FeS
CbGn2JMCgDkC4RNrGczK8LOB/KzYA1VJ9btEqhpM1o8TqtfAERD44YHHigaxjZL/
wnPQs26aIWUH1RbXVUMimk2t24M4YfIxtFzWJmKJAy4vAGma9lnV/Att7QBXo5bb
jAukIsOyxtNeqAG4WPWFc7EKy/vfRIlzP6eQnIsw6jr1UYr1/rQgqrWJS4JKAk2k
6u+MzxHPzRgZ+J9tJW2OgNPss+TbS27u2UGyV7U9Pixc9GKC1CuLzHB4cG6s5Qjw
QFX6EMr6twWVSJH2l/8+SXBRhI9ffawSHxE0JxFr9g3jQJvrM2Ku+MICzlePvfuZ
uokaOFReNv63C4GF03Cb5iIP2wu6raWOkl8VA38lk8kZWFCX2wCgNn3rWD2oIx/Q
+MJjOTafy2i4Y+0djcdPrAJFPhAYLAW6hGqB7DlucxcqpGWDFz7cj/OX3to4qDwK
Vw0V06vNqSd/6QLsFWCZhmzfxAXjBZ99V0WThBOsv2FO7FSuPxCGHaeupjG2eNRl
M/Twh36+ZAOb7sgnbk1YyFyu+IHCzoqIz+PscI6tzJkYwWvDgFp9TH06dFslwmOv
R7aPu56+T5MZWFFdiXZqKhr+nPv8nZAIrktBlp68cqD8ZWkLVkbI1csxwrOsuQTO
TBypmCABj61YUYpi+l9iGw==
`protect END_PROTECTED
