`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QyZRO1oP6+CQ7HxHzpsY5/tEcBioZGG+MPPR9Nuf5L+ZEW9nJRNeF3QTfR1c24Hg
kWxaBHgMnmUSSIkE0SvmewhVI03DL4mXc5q2iWjsrUooETG28rHhFSkRo69N+e8a
W6w+8zoca1flsWN4PmfGnVnrS4eO6O7SE6vM8Q5kG5rj8Q1wQY8dicfpSHlYK/JF
ocprKkSe7GPnZx0QVvDV1dRJz/t++IJlFPs+SpizMTnk3ejzg5wcDaCVO/iOpvNw
BTZKpdi2KYQJV/vZihoK7GNkihiPsrNUJWpO1IEnHCQlLd1UD1dXKhhB/UWHXa+1
J1weTICm6iPyb6MQdkwVd4VqGMmlVoO04rphVU/oI513jRf4Y7QNyeuzAwdrIpQ9
PTQ1nUNvYLr1YXukmxpJiA==
`protect END_PROTECTED
