`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nFu4KRTUcoKfpkqlmXXAf2ZDHKX9gXgEEyIQ/ChhOP1UGCvMd2aMWmleysOhWNV/
tc2GoXkxDUjgpyBsPY/1F76OHV25rWt7wuYXCzRxTpTiXOljkP6CmEzzMigVmXaH
3ST+menC3nJoIy+Kd6xgBK+6j5NfC1tCe24PXSt1cpUhz141SoQj7EQNJF1GxaVm
2VvT/6XuYfhUF/zsrjVuJ83WNFqfkRlecGAyd/V9YXFra9Hjq+qSp+Qa8Wxg3kCk
FJITNySLvjIysMkpc9C4u1YCSGU4xL8+g+FdIGJO2ZPrxHVlYRf+PLoZ3VyuVceV
0ck8kuTbinGbFK0ROwuOLWJxK5kK71toagnMbTUgNDjp1HHftDJ+B7LHfvLsaxGS
pl2o22a246j7kytUWAZW0qEpbU6N57MEyRLiF/pZZM+0QYl4api1RftG15tFRUrl
+SP0W4l1tppkRCzpFkco11fJG9+Ng5wftdOGWCL/nojQv4aegZQ7Vm6AFXFUSbz1
1icp2Vu210hIwmlwDhhqNK4XfNf3RIrvmOXbYKSH/eZROCWhmrdWabJZUYUng8pL
GMflBddJog0gb2dwvQ7nbJpBUBYYKaZ0usoO7N0mtouwvfABqWUFeUpFQlIE2nB+
RQ8pg+mGqI53eoNEtgR4aonRJtO5qlJniBoMSF1Pm30Wh+6CZgrV1SljfIvrdQV/
qWeAsG9W8KqeHk9Z8A7RqtHzmXc6DSwp+a+hEvkpQdzsRbXkAq4RTIZa5Wer54YW
Hi07HsdNCNNCjHMI0/xm0kYyDjbwcwGtcLPO4eZE7ed/KiCbRmh5g78scHDYn4fd
OWJKiUls78YCa+4qtA1idDfSyZTyXfLWTMqTcyPzlS30Ozqd+tpZF2ysWsz6zxGN
fwIYYurxygJZHSjCKiM/SyDiUuU/WKAimhL3iTuclXW71P8h0s3Emn5orukYgamy
DMFxUhuKQaEpOZ9VynLeyQ==
`protect END_PROTECTED
