`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J3OHTjhVNyVqexC1ehuiB5fTW26StdnwCMmhtMqfmp95H/1fT6bdsgjEKILUDfUI
aKC34SttHqRnrjbRWVogeXDgEXH446ECsFH/mvqJ6oeh0qWNajKDyyTXyrdXN/ZP
p+wDJmiZPGdJOTEutxnR4ncUgYwLDiGPM0EXKl90kNJUPwyD5a+B3g2Pdg3c5Qjh
v4GhKgduxBmGm38n66VMybDPsnvDzaPe14JqLtMZmwuCKtAyxscx8wZieFGw+wGJ
wuF2lvrJDd9PVztBdqhU9iPskCArLIquzXqDJOe4n/3MAy1TF0kSibLVazGs19Kc
V+NHFJJrQ5CZXZo8SKGf5AbglATwdHfJioG73nHHJDUPuLOhJi+1vCYVTZSkvtRI
MCn3YJ3gwupIELlP0tAfGrWKReYvd7nITv3Ogm+61v6VfmXi3WgSSiupoYVXY0IF
1DrT4UkVT42OLCig90xJzfALMWdz7uDoJIN66qY6wo/XWyZdYZwV8VCT4Eng2OBJ
xH7dUZfLEjyOJnW4CGV+oPwT+b9JyRuM2T5dEhboFTKjI3+rdEV6rwvOWDG+8ckE
aGXh/10G69pVRldGMDHzJuo7DwCAwcLKk9JVq5sA/sJSDfwwmbatt2k0myLE+w6m
o2mPEyuNiu9r6OaAfhHo6z1Wcsbb+SqSGtTbw96ZfNU0f85teo2xQs6/2ggAjWam
Ism5+hK+kTC6YK+bNRdKtiSUm1hrkUPqPS0bPXMaeBuM3giRZAXpZ1f3YI8wzTab
n9BbJ2yBJm4tGFL3R8pioqxESioyD1MOw8yh+YVKemWrG0RmJHtVXPwYysaez49Q
J5RijcFF3UEnqtgNMOjapPnVRsHgUzSCIursJfEwz8cY31IS7AhnwUgLFZOgjUE+
iHzzMcyczr2Rn8gaa9x9ZUtfEP3G8efCPV770H/gTyQLD0s8GQRcqRbnNfwnAqGW
SPVph/USFpPCLpUEaLJRC8NQXWv40iLdOPqcDr7OWXDj2eQOgi4ZzI/OfwlPCFLk
I0v2HSCc9WlP1/HlA8dlfUp5ISqjZGiWG0DfXjWA/VkeXC7MXsgHn61g2e0/fKla
coGVIVUtHR8u0rr5xRxLp0dLR1U8P6jPXbyHCHF81TVkeBP4Vo6hhvyFM6usGIJN
pmnyEn3BColGzJEmdFDgrWAC4hMj+4b/Ly8uPrPZfDVxM0oUR9C57DZ0CibSYYqv
qlqQiLS32Y2gHuQsmrGI0yKqxi5IN3tswZ7mI8dQBTXiVmw9V24r27uI3nQk0svW
9B0Q8NOyINtRdSBNClAcE2FZLtoNHbcAvQylMV3duP4=
`protect END_PROTECTED
