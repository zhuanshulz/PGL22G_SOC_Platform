`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W0qnTxcGXyAuWEXxGy+E8LpYYpcwCxZgjq+yyPSxmyTd1OnvFNfVo2LvkMeq7kPa
1W42BKxV4O1MX4dcCX93d1Cv1SaIIddQKxHsV16zzEuHYHls2Fva6awnsX7sgf0J
qPV3xIazwT4qAXqLBfWeCNz/QpfOlzWAQ23kQYCxeWJHJogm0vvRMStAAv/IjdsO
K/PH2movskiYYtMC4BBW5YmXqoAYQ8FfQaThxrJy1qdyhkH1sGBo9WPGJskuAVLb
rH/xo45gBYzsRBvljKz3jvJ39iFD6BGfZEwEc6rXyvCwekX9NLHCgRVGdBPW6cca
B5x7i0E5jsAgP9Pq/4k3X7XXsxTpA1MdRXLceVtBgc9GvcCJh6Eo2mmhNSiMZ0WK
+NW7ajAqIhlRDgrnrLEoCvQ5xOx2pn11K5KZvVFhca4ggMdChy9h6yssYXLdLa3o
P/yPkbeOzHcQYA8oFNJYZ8BDr0p0R8IC0OOSqAUzuTs48hR8DDSu9eSVgHcHEuKE
iwWpPJfamEcG4FHyQsXb6Dr2J9AOz0sjTw8RqFo69eV7eQPNfCsQubG9o6EFVsFc
m+KvnhaI7mkWLox37ctAmZon3rl2URTLplFZVH01ZGvYeFq13s7txL+Z8zN37BVf
niAxOFGMtXNZPuZIQF7pspgRNmFizIIKrI/DHkYj0r2UrK32j36fWNovGcZ7DZ86
j6ejLOeLJrvHt2LRw9LlBB84hHSRUsYATl0CxJWciQQ1r1uNJZHWxNTGcTa44Vzr
PFd/rFXhIyPqARCXSj8Wb+i7AZ2WjQ1PK2jxktcsmclb7oitBIqFW8iEHKUAuRB8
7hsuQCVqwMNpagTDXPWBig==
`protect END_PROTECTED
