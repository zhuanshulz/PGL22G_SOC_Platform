`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rAHA3XfTzVCY8C6QZNek1b1CdH6kJXbZTvQhIJtSMiXP8U5arZW3RT0vr+UL/D6U
jYIeyfvI4jaGlnCxg0sYlTOfVa4godkcYqejbBxdL0Zk1isj+UGgnLgAr+qZsONU
FI8p+xZmxeI6mfi/oMlJWNcpuk3ODKM+OLJVPtJHYTa2i+5bS8meEgLSHIXrzUiN
Qnve53lk/KZ06jD2VXyq2epAS/3KOVwY3VsSULfcpbuVUibfbCFspbVaDPLXFYoJ
kIJV59mUNR2cWjuaDU4RbhPiCMqftRXn/CnrA2wcZkHR7VS7OUVD0rDj6ODfYRAH
Pff6K90poZOAzXfmbhmGi20P+y2r2iBGDke0QWpJG/d0ypAUA2VltpnIZ4R7MC9d
pwjgtcPai9oSXQNaQc1zP5vCi5GP+UKwKSaMqy0kpWApy4lEho3RplKReN+EDArT
odszK4w23MEYKFisL8v7y8bnL50D+Yjjdgu9uEIMYGbDmbDPxfJej/ZA6LRrHC8Z
iyLcxmhe24DNZF+pDnjlqeAw72hSmDWIwBNc4rUB81EXxTL9wT26vTztfB3siHlH
xENWIj0xh+fTtQJzZs0P9FuKhiUwOayJ8F6qeZDrbVF1fBJS+Xseuqbsq/EQCcZR
ZXboTKL3BlmjPS3dW1o92MGF4XPNOrgHrUrDoS7MZUOB7ASoyKDAzDHWyd9zuIIF
Pm1b1q8r83ofLKvNp5FYJJsuoHvv0Nnpk9KV2dqmtVTPh7FnDk23x7YdxKNdmssS
+N1IaEBTXEoJqU44V/CnH05jlZD0dC8i8wZH65XT6Awor+xZMEMCYtEFzpT+X6mW
EjN31P3AGHEpczVhDxvEk0E84uj9X0sWIJIXcz0CeZo/isQOOMnoV/EqG0zyi7oa
uMYdGMXZOcy2eLI4lqWUbEmWbFPs1/EeqIlier4ieRjZcQgYnBTSR9/ea1GjxHH6
mtXP0hv2PjaVVLJ2b13aG2kQMA8dj12K/1vZTwPeWLQDQHTkhC0gByOWadwDSMLE
4s19GrF8MaUYv0RPCuJDnnS0CrxgS5ExzzgkMP13tKw7PVlInfKCPuu7yiNd53Bq
nbM51munycqoXf0uPb4bdPfdzj9IfUHbXAM2L4nB9MTgJ43mSzgfd/Y6F7ASRawI
pxodPIUPo6fm8lPU1nh99+R6YqK0/RSGwyhAU6p0U3IO/yrf4Eeda7s9bcf9tKSy
oPjh4kqXfZxoZOCQJmKUmpy/xspzch517oOV82d+VCc3U1DkafVcSlJutZ9d1PEh
+LIlnFsTGZXkjJ1/v+IpvE2/zO/U6Y9WugBbIdwtJnCCKgy/5x+B50BZfc1ghrob
QLObbzBsEnN7tLnRKgCMM8JDpSV9IqcY//OL+46SP1jmidPo+0mI+ONaotPLQrn8
HOF1ioqXY4fimSCzbWc4yF9zZKRSz2mGZNBfJzOf5/xpj/mBb/q8/ONWwJqXbp6j
v18Xh5vloP5IplLmchOO8GS9R+OsiNiLZ72D0FbCBv59PTnIJvUcNmNi8pTHNnIw
TtckSpWo24KgzKScKhuL2FNJ++USMIkqlfFIdOCjyeY19fYBCZD8/WdwBWL+iWJg
nWsTJDf5BWOb5zmzlrmP5CA8hSI60zsjujG6Lh3MuFuCW0Lgcu4YToZKQCvxg1nf
`protect END_PROTECTED
