`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
65ArhQ0/v6/8/VLy6jJsruyqQ2APdxcsdZGdU0CSK9C5uej7sl+l6ldcDELShAlX
PB8j05Q8KPMakFyT8gh1gmA8gWA0m1zYSVp87xNg6Wid+jXJ2vSRxgBd8J/zXrC2
7B7RrOUH/IMQyLOb7sUNk1u1mt4cMtYbC5Umau6xNJDcdK4frjaoYtyK22EQiGea
PM76blKz9oOxW/oDRkuaFeFjJEjp/SY4Mv8/GXkar6aWy4c7uFujH6x/dn5pwF4/
s0EtHHQXmgSXJ6ccOmmDxqSU9g/CIyrT54ixbxLsTqEZFdM9Wu3f4jtgMffNTbmQ
bbbhrfBkJLtEQ3jJ8DYicp8aqvj+MUXZUWgjo1A6v9ovjnZjP7BtMTiqfgARIKGo
jgmc7Zvng7m6IA4l2//24QvLxNLPJ9MWVTfuIx+LN10Li33QajiaN2kkZIIy6QYx
iZbX2bZqzcjwWC8pcT/+JxDAWm88EmlMWy+wLN1JP8PxyeCOi3sbFvMCO9cvar+8
l7P3QIqJxcOPVIiz5vUYzCx+wQXRYO4YbfJkqlx0SEFD03A6MmVivO0evYyOI2dA
1NgxpLQ+vWs5KSUcnbgu1m83m/dwAeoDoyAUL1LAJ8dodZTYgNUfL+d43eVnESsn
6ogyByKDqMt/7xf7De9aJZE6Kq2V5QdP4Ki5/T2qaJEUGuD2VsJz+Ak3PJwpTNeR
3LP08XWl5+8n3pLqOqkU8JtTvYUt0XDpGUbilqOEqEbOze2UB0puz82GJ8y9ah0O
JuoIeDPnY2sDMfFUFjhanRZuKYZ/73S/rXd+EX1URy6gsF75AAmHaiDO1tXbVqRQ
4THATcgvexKIYL5KlTiKLCQZrY8q4HDmg59NoqtqLj3b1mAsERNQd6vYBjZbOtYs
hH5PoPifeiu46vyuZSCmmmpTfSu7yg2erMM0/nCgrcp3IxkBx0Gg4uQMqhEltSus
3q6rL1zMxrwnDNEJl/7McHZqEXGvTfHu2kVbauIv4g4SzAPmPwcxW/FAa+WTUVb4
Y+zO2p77CgHPGmNY7+cqd9Qgfw9JfzjAAMzz/VAh/gseaLgtYFPBUdrMBfbpAH3X
ZRFYST9+0qr0Hhq3cbYL1CTUr37eItnla7UBGF7Ih5MCj7qWRLcfR0oNxnn5FU/f
V7jTGoyh80VgwRGJ00Fw8XnN8a9E9duAU4oWFY2SPGK4U8GQUSQMlNuNcuGn9eHV
wcvrdcg3TgwVfLVfkGoR0aFjXpyF8Uq6CwhJ234XF4jTbr0HD4+mh88WEwEMqosi
60xFGiTf3TyrovClABoBf8IhNJEFjjTK2COdLcDvKpPmT0V4qomfnfnk16/Sac5e
PLb6KDkicJ26KxdL+6KfvWHtOW5LqIwZC+6gZhDTo8MA04GFRKeLbdlRFrcCDqNz
0gDEG65GORLY0xjFzLBRTL3HTAjjMHiN+cCIApy+vTELxENbNdwO5DhrYrf4N9Ru
5QHQEBbtxBEtRMfeXCxL+mOCumyEwm5Ko9H/ppimp5lQf/2nEmZDqXzJT5jZmgFB
QCH4uqQ45xmbcL3TSfvYERb+wUPhOcvTr98ISpMLCiK9//OCobT09Eage6YxvXu/
2auwcK0Dtwpj1a1gCAUDS4Gmk1mu/bi2+HziXIrhmUahziY2r0j2+/V7uq01UQHJ
fMoTrITTbJKnIWiqMjwUpgBv3DM3xW2WZqe6Zyc09IZqaARW5iysWmG7uUbgR8ax
L8LxDJNJJqVIu0BXBsUukwowNKJhZzt01VYtcdD/ExwtvS8am5e+egI6/ZlxuEpb
DyRxmd/Pl1qTrX7AorObbO3/JIVlcaM+b1SalXx5m+kCotZ7NE4vuUcURxrJI5Q3
1gjWYbhVkX6f6uOwjZpEH7oncapeAjozSWdrA5Qk8Rc7U7qR7qZcXUqtOb7XcoB6
UcAaC1xp8TaSXFDw7EP6hZ5XjHqxwBKZ8K+G7Nfd8Lqd49wVjocJ83+cDFlMZWIw
7Kt3FUUI9BoyNTiCb3kFJL4iGtr6BGev/QO8bWvB5c4Il993KCp8wFjl70XFfrOa
w36o5mrdKWq2ZnOWPT63FcbLnIpM8hgDEXoAv0xjXYgaL5BSeu6eqFCWmiFSvmDA
+Oq4J4jeql9Fe7DXsDJzzwJ2acKHBKMXTTjDzpJ5JH+sEeTZv6bW6v4N7ec3tWup
m7Wsi1CwvmQfhmno32gGTvggd8mWweDubQ8wqoQuHtgjgI3cUAjYR9SIFEA+kRp0
6Zzw0/4M4r337zIlnZkEb7d1EvwaA1lz/vJ8OMPPc99TSfpQbeI8YDdmgb7BPeoN
i1D7LuUiN16FGegQFV8Ijo32foi5oJSEcCOYYORZiUC9TFr1kiVYAHQSyNMV60jq
DzzI/z/u1uHGQG1wn6LTpNU4jmTwOXCvDx+flBSExX+DFYgsQt5SFcKnZdGntZuP
KrR0oVcSrEezCy8dwnlUnwVxSTkxWgfwmyzm2a2R6RJJOcHp1q+T7KXRN5G3Q1NM
mU4oY8E2hhp/pbjIyoDHpu+92kRtooYTA9LAT1fhHVOrzpJjUYyrd2EDjD7TQ77+
xwXa5CwQL5h7aWb71y02zc+ubqFhfL2mw7B5tgqmk4yJDdYhhbS8RjqXeMuBj0Lg
KYTEgMms0U6TF07haYcsDfh8Wm0rCv9LW47EPSzSf/ccwprI8dKbdOwTmIKTH2Da
zZH5tPg3OZL+eYk9inpImUg+q6sS3/3xAyMPH03UNODHquKaMsIjMIJHOV55zH7Q
gnWgRyvGjqXV7a/6/EFVkVFpYMu56br3+VENMNoVdqfMQcyMJvfC9n7u+7bpf3Qi
gd+DcewtE4ftIZAG6kigqUW8YVv5aptk1dpO0YHVQQIwOv0WbMqB0k3f+oNU1yG6
3+WbHAXZd44CGMcuJmUGoi+UQaaNAfskxgUH0r013lGsvmtOaO2+ItShfCcBGc8m
4jZmvn+Q1Ay9DVNOJU8+TM5FjuYL6v/dQXXo0QDxHxvXrf+1w9goW0ngwZHt2KFf
6Ft2wdFQfDWv0cAFKvYEVTuqBiHZGmf6ewpD6KEZPorqlVyJAC2Dl/z43S/nbcmX
y/4iaEW2erjJgkgZxPNemwcqg0DJaKPpJnrEIVn3Fym43Jm8LHxM1oC9Qh7qNIg7
rer07y5rjvBzSd1jncm+4wDb2qgIAiGFQdBkxWCoWuulJAvXwWC54+QzW5VHVULw
MY+IF+p0GUy6uz3ydQmeT6eL4rHIizHVOwo+XH8sLpj39WqJjY76poSRddesb4no
VaUORYtyL1sO05FG9Jiw/p+kWYCCgN0hdfWcBXgVbBy/pTiTfzaxIpgR6lAe0x/O
lHy6CDXAe+X+I6tqog5QBluF0fd5iCpYjDdjNIuy3jufr5/pyirVanDTwKmjGHei
WLUbq0iWoYzibH5HN0ubATqImuqO/e+L0jRxcChiE/BPcZD5FKLQHkGKKxfGmz5r
8u+b245f7TdPgt58IXUc2KPDPAqOgUuW26wCLjk7yJb0+S5h0dpau7sPDaHMqCp7
fMcZKpiL2rZFLk8ftM/SxiU84uzftOOxHrif1C4ZquqexHao+DgosGuuXzCHFLwd
5TY/zkIO12lJVD/K7wYg0m5MmAcMPxEw9y4y/Jb0nxOC+14Dsmcog0XDaX23WYfg
gPDRvIvYkd0nWE6NQPbFlj7zGm4WAZRS8YDYpNQyLp/CToXt6R9e/6cnD/3YxgJV
ra8xpmjtR315gfYRLueIJEJQA2M5z1f3E7BGs4oPsa4INfPgG1jEo1Opi6B6Osml
j63ob/JiiXjmRxnmhZXwtTl85Fs2sZZry51nfSfPHzlCT9Y1PyBB8RXm+QawfV/2
k+DNPD+JT2T49qBhJi9mK2P4uy0SX3gKXcZbjqKJxaBwo4z2tnoVGD6qhCPAYeZ+
HjYQ8smMnkQg3UpIAdZoVRKhnSNIJYS04emhMunxQ4WX/PtqphuruiUb8mh2lKWV
K98P2gZ3v3vDoD+yMNFXMMYTtDnHDqz2lSL4xi3Im2j14h5sAXvoUxJ9+GHAJdX4
rN5knEuPxUnc3Xb+7RjCXVGjRBb/h5lE+tHIbe/PzLqcbfhUaoCe2Lq8uRwyoiL7
ZIC9RcgQngb9HowRM36ff9jHg+ntRVACMWLPPVncQZb1Qb4UYpZ/QyArfkMPlzdl
z4JslyAOqMADvfmLaqMBLapPs4t0LqRPilpUc/PwLqSkSpHT42SvPq8yHHd47C7a
DEFdnUP1AhR4mrLZWBhkfGQ3iD0i9t6PEMmxuJ0EFivkGdGei7sIM9NHAvxFC2sl
uvYG1qYeXbqfLh0VgVwHLwxsqzOCzYSCyjKMjmWz0LfDyE5+LfO1QZPv4o8FtQOA
cNY1w6KwAN17OWTJTe5QkunQRI2yuLUGTgahFSlr59MyDnEbMMM2t46b4ekf2E5v
3XAie9vlsg5A0Rmumci8tpQKxb9hhhb2/SkErf7tlgKJU83q1L/8Efd7msXsTziw
ka9xJRn6ES6g15q/JKFxLgiT2BjyFSSKEXgtpu5+tznncV5GuCNd+xLKlR0p7RLo
4+qKdiDXW8Jg7/05VfWvN04RFQ9AfYEMMriwvAgg2Elk3Ngy61KT7+BzzhSc8rgj
PBaXPz9DWZjPDLyImdh224marjz9FcKSbrE0JJPVrcRQGo9HZ+jUi4o2vPjVjwuh
9r3+8FoE3P90bsVVftJ0DjAM8So0oLYxwiP7I4c1lprR+uC/tSM05Rge3ZTqfqoa
yY82A+PvOa33OjACYgNtQ1X4SU3/eZXezgepYKNIPZxud43b2IdVYctbK02QXT7m
S5p7IOx4VSYSFmLKiXkrj14fXBOCA6TvlvyUhoiisai4INWaEpjj16QQ7V7glxiX
CJooGZ5grqiyaAVuPphPAIS02i+Gr1Tmt83ijgewc2j06Ejun93riO58Bzi0kOw8
LR8JvxJHBXg0uI6GuliO7dhYUOstKFMtVesqzFZMazdK6VGiwR/T0BZMTNfzuAO9
zSNPU6M/qgu2uvp+YXEZa+BfR8CtZGbZyv9W9anZsLdwcvq4fmcAeYK3PtMKVLb2
fJ7nRTbSisPXJfblTm+gTQ0KHR8VNr++KMMBa0UuP4qGPQrHQj0Fbk9F/kZW4C3F
biHP+YJSGHV/W013G0Wvrm8UgOY6U5oMbfc/BBLue/rXvMwyfYTlE6WpM27sU4bb
gupJdln//D3huWDhYTsXIQoHnFTz8NtvBxE6hxdoaNuUrGIgMbDb4cpXQyNHHfA9
xZvFYyWf0UCJGzobm2tUaED9FLQozfiOr+NgNzAewnxkLabRIfA/t9SqK7i7ycWN
V6MJMbexkFzSZchNu1EXGh5J7nrK0P+ogx+0lpHNw3edHxxVtRW2mMsAaZV/XX3r
4VB6ITusDIgGOdXWMRWY0bhXmxQ/gx14OD+ulA0YDJSwaWCb9Y8VgokEjSmjr9Hx
s5p0iebUshRDlyjzWrtxhS8NxJWW/WnZ9brEzKIJhuHqgqEqnRWITVbPD+TTdP7s
Q7cFAhr2C8kJBx96/+5T2sXN7TcrJ0Vq49sQMP54vOfn7yqmjqMkUmz39Til81HR
zGHT4+V01AUTv9/MZDCEYolWpL8vjTsrVHPKcazU0ADd1kMikf2//OCMfTBjHW5o
KAWaYKEXUFReb1lptVPo5QCYbRbu5lhkJwmVUe/sNaKCdqZ1VYio7whB3JQyuta8
+Rgl+WjMPNGeLZFbD+FMBP+KPW+jB6OlGRJJ99BTeqC9T9ywD2Yrl1czcajzHM67
faEJ9tNybkKdT6q/RGT5+2sqtNXrIIJuGdcZSvELqSlp0Qz6HuDi9NeFESQB2UoW
dtrhA94X64fcP/L2HDVMb0GgkMwFIhkS2MFd0mEyi6yeKBd5tSee8DexTNP5YeAI
RbdNugTUSlUzw9YLQkOPIUqOLlmwMpHMi9Y7htB6gCbDIGbAAKJ+K6Z/OGdgjXED
gv7D0vpMsdm3aV+63qtEGkJ+X+dybuftME5oFN3P94V2ERSVyDnAmfUBkgaJZWRf
5yEKQrb4OXFceZhUrk0fyhNfpdhNUNDAsM/JAiNJMx+uv+TzXWAvU2kRhEXnMLXT
OcmqtioZwVuUTkDZ59ZSpn1m8Phzr0JjogLAoXcLK/fHazdHAe+0xBMngGqMkmBT
FAgsZOTe8Ml/06+vHSYR8K9IZxezv55IcSXVVE4O8SQVUW7oAzaykoboNpE8XzzH
hKaY1+IxJdJH++Gto+crGTk3si6W3UM+XROWGs3k1czBARs9gbTEZS0SJnpCpbxb
2L2sucCIuDmium/ngGjqixg/w7+/d/0tw3cbTRxTZOWRSx5WV0UjTZx3+7YRpLmY
Z3VY3e8Ys896i9j2hLIyeCj+4lgRgbbN9uVeli6MO8gHSA45v7EpvRoHPMyr6Fgk
3RJFfCZ2CW1OzsDCseHeqyW05RcyIJlXzkiXkC74Gau9g92TMIT30fAaQgeypvj7
9W+4fEedQwBF0GjIyAlu0qHh6gkhPuy9oh8XEQFIdO0ip1oGbX7Sfbmq/ZAne08T
EN3QdG+5KYTs4Iml6aQG5jamvw95KxmUatuegYecWw8H80eaZ9Aq04Wq/y/MFpWe
fLqePPzw9dOPyxmDVdKVkbubOBW1uHiE6y+UDwaNAC5GC1x+ou0DTzpJW12tjImt
YyCGg+eUGGuW86F8dgcXADamu+4ItYnW5+wTbTJEUJq0YJGzrq8NAOljCu+WfROr
juFwWEtyQJfLg+HY9MVfed3maMY+oZp2mLdG0XQJXmnEgEwTEnvwgzNHBW9UdLWK
oWXP8vB+1fBDlLT2hbddEKGOnroAZKqwiomR8pyGukzH8Lbkhfa2FUEyKhVzOdrQ
mwdQMZ+Dpk79FjVFn51x+kl7WCUoUnaTHG2Tx/CFVzI7AFUzRQiqq9cJhA7TVbUn
Mw4Xk0FJK9gvVEH6HPEUg91zB9dPIfRVUE7HKQMB/hX/QHFtnl5+peC07A3RmS3o
19kQS9gL3jTRoQwvinwE8mIvn6PVlE5R0BhoaL0c9z7OiYOaYV7q9aL2yt52chBa
Nul/be9TtFmfGJ+1Ic09qlEVfquFP38g21x61Xi8+IeGIPQS5R0MDvFNmGHXDQxP
uSnTHVecrh3cFNuDu9VuN8quVtvKoKAxK867N7Q5ER4IrSE1CWVbm13S68Iv9rvV
FZOxV6gCUwU9gJxHwSRnKnakMoqjxnj/5YXgsdQLy1Meh55HAbfDWJ8V6GbrzS7D
wuLrqDS+bJqobhl5C4knYGGv2tn8CCl1NZT9IaJ+JvTJK3GLa+U0Cxmu94xeyc+2
MPTGI3xvvNm+ZHamhd7ccRCXy52K+WneYLpRqoyXYfEg+m3hw5ABchuRmp+lp1v3
dukt40F5lZ6VEzhyPI8V+meCfWfJoCIdk498pJZdx7Rj5Diz/Odl3emnBbLsTPLo
EVM8gRii/CLjpWss3Qmv65DL27M7ebwQPyA5ZDFLgCU3/gjU9Bf5ROhKAsVNT1NQ
ECzaUXTgJFmh6qeztGLZBS7c4QgJnnn2ciB97R5W4xeYKIlqFpGDYbtw9PNWZgHE
y7TZN2rW2Nm3AB83BLmEwHYe5KoHs47jHWPctwXOj3J3kTzPQyjwcIzVlU7eQOTM
vxuOQ3+fqOPhqUdjTfu0CaoulXH2LrR3o0175LHa+6/u3jXx6B1QLV7bXN7Gm9eP
1JQ8GYYm0jFiQzBhHgIcqr8uAgSpPH4Dhx1jYoe2+UPdGcXW/3lF/omlA/FOLpgx
GPbUvHu+r9BFSqMP6dOr6K7kHB6qVvJEwlrgUxRYwgYmPE0StBl6dvWYA3UhIM57
JonuMe0HsG3AiJu0LVFjNpMivJvBTZFbYAoUR5e/l8LESA7Fp/PECdSfT8JijTVx
pQHN/LxCRgfLmVXIk5qI0LtBF7TlipjHKcpGVge5I5DeaJR8n2Q1lEdTfbwYTTvG
LSmPfN7qXO6kOyCl4YU8JPHf0wfg34ZkNNFInQ2TxxgFZMH2qDAxx8iUmzR0i1s7
t4yoqCXgl8UsQKfoO6EnlbEXXPtVvLbMYD2jYqbTCWqFTKaNdlSQO2PqRW+QGU5N
uaee65KdG5GZ01e84mCNcRpyVsoqwvEPtDWlYCqif2W1vv4hinTDvVpqFqq1Cc7J
SaP7xDJ5FqjiUhH6IZWj9cvHnZ9SIBZtKZwh3QMkzIMXD3h4TynpHD0QpGcrnprw
6dGj4+yi14rD8gTFZksQQNSxrYfRqDkMl2p2sW+re3GY3E0z5NQUN0rjB+47K8EC
2vZ3uohV3A9ZpJ4mqcZUt4mVqimOspDStz7ULBvubcJ3oTP6/WxK/OV9dlywe2RA
iV8G5FAUB4VsVeown15SiA2apmrIHkB7dKsQZ1z5fgi2qBm/7eR58iHhtffJPxiy
9LWvpJ/e9amj3y96eULN1LpUNQJ+pyCTyT2qYnvIEpQY8NBOi9k/Vuyhk7K45o6F
WnD3zdS3LTad7/KSKUSjCj/UDvUDW+9yvpY/nQGYYTQ+cSmGxGitJI+7RDM+YHgZ
mcjgxo89/tM2hki4FT9fbMAOpzuIkVP9mh2JHFpdCALlCF5nEp3FzIWsjBa/SfXz
PuFrrsnWruMGbCV5wkiPq7XZ9eKX7bNd5uLuSbJlj5pVctGbimkBD4wI42BNdJib
9ePKmXkMOn2axpitAiODSQEIbImQTdGDBwXWrbRykihHheRpoyDKpMJQt4ve4437
ShJ9+qzY3QiwDC4B6DnBCcVGyW2G6+30o9IhJ/oisrlCwCvkQHcPlYskJ+SHpK2H
jb2warbZe6iNCU/YH7+ZedXkefPb6MIzysjM454JsJeU0stOdPLnPcjYEaWkU3gm
GYerrGdP1Cd9PF28+Lpn/D7W2Rr1eEgw2h/YfD664E/ZHkSP/5CVWe2BB/OAdGMy
Y/qt3zlVJzkzkuy7b5uyk07IM6Jo3txMf/3J9JaqfJ87rEqIqui8HERkJLEGIcjJ
G/ImfYVayQ20r0/3NTnJqDf26+2lNeh1NE4Y92GqFb7BI/6jMJ71rTRWN2c631Sp
58KvSUaurL3burrov9w3NLFBq0W6vtzPFC+N1txcxUy5YgAc/bV/2b/GNkxHv7q9
vyXGbWYedw73p9jY00x697vkzFDvEJk+TK65r/zipJsMo7abbuza8xTrBRfDzo21
+Lu52uOWt95gIs5LH+zXgYVLBMTG97HQy4nkKKNgqIs+WzWf76ifImqwmUz2W0Qu
ElsELWeQqSKyyhfMlS6fIPUjr0nAYHaLdtvwBnKgoWStBoD7ltxfuJwfD7kQ+FAR
n/WYnwGDdwhvUPGTwUlzKHnf6gk/kO7cSg+n2YkDtMvaWpUtRYnwQz0jWlmFWP1Z
K2ySQ9ObMS/n8lhBMf0yej8JQmO+e8sbJb0nAmKk/a88YHexh0XK/vXvW+A3yy4/
L9nPkEaFqY8WCCaU3bf62m6XKnDyRN9lXnN2qRYfRoaho2Fs2O06IIaa8kXKMUiH
OV559qfQRbu8ki9S6OCCHtwFCtw0Ea8wvNhAccJ6zJFYKLrC+jqJwnxrT7p6/yzN
WfHf3A2l5J/5isDK95vcjXgzdDtBDcjnOPLXJEMQNz6RjjrNoUuNyBUfFxXN6C6a
GGrdXQmvUCSRM6wnDGS70wJC3fHStiUs6GTJRlOwc8PYS+0reA2gJBJva5aPsqnx
KuRKwiByJ4/+n1GTaJb9UpW79j22KyiXTEgDZ11mkYBOYyMwW+N8GO2xQg3acTrQ
MHSYPedVfuctR3vUbFe0UzlnJu2gr9WKQi+VoghQDdWVmmFZnVKPEnhaIwGgD/+G
iEY0CtSnuiBp2oG6vrfZhIm1iOD5RhRdP4A5sP75IcN1RbOnt7so9hGuNZv/+Mcy
f4B28YAI35/T962hzwwA4OZInZlLRsVgUPHW8i6DJA8AvpZ5Tu6/BLOOr+cF74Tu
23bxvtu5yFC9WuUVa5OLCyc/viFwbi7W5iQyQvulR2AiQzMonlAVIkbP/R0mn1Cy
VLR3eunCgPFItDBFYSKXzP5gIFMEpprpPRYghfSoQ2ttFgLyNlNIPiob1pWs6bRr
rCEAOv3ZsZOA71U+mirj7HjtG1imkvhIkL0+D2rEGuttDPBfRwbd8W5qxqA9dfTX
7m37Ya4atrHQ6rMY73A/kyAN7gS3jvpmTKfKxzFTKm6vzYiWaNymHQbgwwXC+geX
RjJ5SRvvD2LxD325hzJilzQq+/Jnk0DgJmqqXLHsVsUqaTkPAJ+JoMr/sSFhm7PE
Jniu0StCBm8Yez6FeSA8Gcv6ZR0RyNQiDKr5TjRxLydvT+5OKZO28hZJCNsPesIU
bxBrPRdIqZ8Mt+9L009hHGbYXK72AatXexDpqO3p5EnF8aVy8hGeLHwQXmh2hozr
ez+Lxymnqkd5fHRzHOnN1SZPS0NjqM5HUyn5cglMaTy4+mQlwKSidsyku3UnOK/J
9qeAy2lrAdpUVJr7rOaAD/vp/WUpSfmmYV6AYhCS2iir8ErvEPchbRrxZFhI7ie2
sZ8WUfNdXAUUsTSnuyjZRoI98NSSMGZItKC2Y3hkS8q//59qlMfyKVARvZvbIpgP
DaxiErEt/nzq/ELw07Ci/FFLetzrP5FWB9G5MaaGrXy7J/EV2+fzXYB/6FHSW45i
UFA2saPm4EUR0QdIz3UbvtFvL1LurczDsKDziqDllfPwRDTkRJrKoHPzSivP+hJk
XZwwgpdQ9/2XTtC3hSgMlANfQVTpzEcy4Y3q/2HERaCzvm5wsXlBwWZJ9mghaaL3
x0lhuBQt7JOH6ZCA7GF6lwbJF9rj2Sb1hVAHUB+FbjCBo0q0sO9bKUEuBUnjpt+w
3zBDULZTbabjoULnSMS3+opCW+gJ8himPd7EwE9LpQ4QflWbMuLRgGu4IHd84Hvc
2X4y31LNnMcriSA4a2yqB73HUkG9wgBL7hx5WA/hmjf3cm284A+lpIUEc4XJ+MKn
7aWoIOOrXCP8CldDbETvqjYhsQEr6ktOPqMplGKUhbr1S/BaV1kySpeQT2UlzFbV
UFengF6ftGieyjW3bSAiB52AYOwGdBJAStGVLMjZ/42aiojYpFOjxE8OVigjyvR/
qR9e6nKOWdH7usIy8Y9fmqs4cMahZeN2XPL3oP7UPoX/9765ymDLaPU0KDWMKj87
e8PTrHd88krr9+UepHQPmtE/LU7R1MU9oZzXmp4ixRz1Xzo0SgeF5Lh4Txm5DAPG
bvFDP2nNYY8+xltaf3+Q10gzrvfnQFHnxkIWO5d8YIsWIkksxc+dk4QvVXE6XYnS
ndgcFo8Gm0lI/LvRX2IeyhQCdDZ25iapi+JylVohmkGI2/MDK9PKYc9BzglQUTJE
shCdHM6KGoxqIrQyoeRXDUaUgOG7Gemodn/tWqUwa0dn4TrUgWTNCGqlmh17t21Z
ILUngJJx33nC/wJpRWi7v/SfuMFBXFsM4QoxStZle8CdW5mEqVB0i4V2HbK24V6g
zHgqtcokgqoUGvgwON56/YQgz9DVA6Pw8dGdW3cx1QGCLnuNPivwnxkf4adsL/od
9FpFcq0icDBhmwqkWtS32R+evvQ5hndXin/nEAUQlv8eB/XDIb515V4tWVpQZOcT
fVRgy5yVMGKQMAbAgWZ2VZhOQ3ohS00G+FGtY3lBZ5vcDp7jAGVXqSVNpOxy2hxI
LxxNon31gOJVB/cjMpKENYaI3/bDRowW5bwr3HS0i+36ivmsXFkFa4Xs+SkjbNn2
LS3dr29zmGeGMD/uaEhLG3KJ6wAD46h0OluWcZlNqxY/SSpi/NBJFojWUwxugdY9
OisXDDZNi0/M6maygQ/dXf+pr7Tv2Fn8n3T4srTpTFiRno9XZ9jEIXAeP0WxdTln
Jk7KT/eiFqGoP5ZCsBsrIxaBCgoPhcoNYTxmykcr81R/i2O0eEX6wFX/NGoWZkU1
h1QnoJL7GbnnODIdrfPe5uAwDRCu+0sDl/preQsXroexraZ98ioiN9AZVNl5Dw1n
3BWeLV2XIMA+xil9jF3Ldg==
`protect END_PROTECTED
