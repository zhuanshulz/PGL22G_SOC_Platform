`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mh63dWC4pYAwyKW3Ga/Oys9dJ4VRrRmUK3vzz6M8sFfp0vqbH5JiRkQMOCVzLBCc
uT+P91o0kOgptqbDy4AgQbHLyqAMCIEqN45vdXv/I5KdoeXNIOwC5XSI1zmRR2OU
4DdcSXTZF78wRSrxwJAfNgXtCm2nrTMGITk6tLr2yRl3oYlF3MTMNoxNSSKqM8OW
HM17qcu3wx2XTlpTJFxPojR5vT9ewi4WHukqRT5Fsb1TFjaGxKkTvKmInbULjqNb
5DuyxkyplNeeQWruN483oQWQSkO4U7RYvHQmxFlHYeDssiWDeWbEfhHIiE0+KsUz
oDNrePmSSMhYuT+E/Um/VcPzjqZbzLgTDbdSdeMIz1tKz8GQAgQD6tsIyXN+Osef
7AbDsoVIyk4wMXYm4wvZk3X/cF+Jgd1/Mjm1IGLGhpB0tTM6WDcaCTSKt7S9x2Sw
ddyLrKMUupfQ3j7o1nkao6+GMo88MHEBJTtCBWZHVR2eMViiPFYjHs0/JhHd4KUL
IlLeYCz62y9f3lSkWAz8Ge8X0eSLvMzO6/zITX4niLI4WMLrW3HhurpW21TycnLH
DmidrTBf9E79/5Hs6t1IJawe/fEB3QuKRzMxsi3ya+PuQaMs5O09qCYzA31+HN13
Odpoil4eHewiOIhqJagLLMPoKwJHkIatjcIU1OO25IEUCTR03I4wSX5zan2jErd+
T5EItdw6vBnf8kIwCAosjBs+VtdbAMTOoYRPyxyyjKcldDwKmaGY6ElTmGOX09U6
oca29EtYVczunqOJR8NC3zJyRpB2aF2zG484U2OyF7O3Ya6mCxTkjEK0aCy217ma
orocA15MwKoOfvtyNZz7Eht7q7YrzZiA3ffuoTfLtx0i7g7U7SoibgtsNgYKHYSt
a7FeQ7/b4nKhwWZMQkVHzBAUVVbPWlnaOswbFYiWr2U5ZueuWYiSf1HUtHDvLGuu
VZZS6VjTMg5xDjMKefSS1ukKHDt2D7LneN6GgMN4/YYD9YnolaYUYXj5nlh7GE18
znch8kNrXoVkds5ys/9lnpycMZ8z5TGAR0+snr/Z5ZkfY3Xc1i+u0u4RTD6u2Iwa
y1QGyqQGwTFFklgsPu2gZ17IAcctJ7IEGpXgpgxGEcGEXgZvWz+fLee8Rcnz/Mpd
PEGmeSycuJ6hGd/P09wXk+XGUUVj9zJZWV3iueJcWKEjTy2jRilfd7pJK4013ofN
0mjy198Ji3Zy33o+U4vak+OIWe7snR6Jc1UVpvD3dTKuICRjoY4Jsog6FLRoKovY
6B5x+zIb+iJxWSk079wMREPMJaR2WZg0EcECUEP9wtuE8d9y4wPYTKcm6sK0kaNZ
3pvMqo+Mkuzf3OX3pNwQ+nXIZ8G9iBhhcrJhpLShsNMFsRkrbWrgjJugnhqTHJMp
LLQlmsORHwy3TiFe6LsSBVY0MsLlUn6PWQtHSCw7+uJo3PIACfWi/jjCDJ4VxvSp
UXMFl14lPFX3SLoYk2IJbIkneFSthGX/mauuZeIFxfpr85x3w2h1CPu7zwOoxrOi
ZZ1ynE9e/+zSmXuCPxxdewPdYnqwAmaO8FSiuBUm4rG7c96p8/vPFuBRJtFVg8Ev
ZfKmlMTjYwekNj2M/3FSE9vbu5mJJw91Lpz63mElQVBF+3VhMx9titjG3xpxYjd+
EdBtTjtnVoYOFBEEIq45PL8E+50SCo/fbg3mowpFtAOdL+ygESd20c+xzaC5TBts
JfHpji/Q2TZMvPnszIME8N6xHfm2af0aaFbShJOCLf0TG4AvaZaQlOF7sDkektEF
aNKs5z0+DuY85wlvx55LcrVjfZ2FNlUh3vljmIrZ5tEXb/TPzf27rO9T7q1HdofC
EDSPGGSOOE3dkHYXbzyir89QdA6mgMyZF9OWRTN/oTwaSmNyjNPFo+FAYBFD9pF9
WGzmMdNHlvCHArMIm8GMu1pJdIE7n2N5On6BG2mTQ91oQjcrgORrEUHydvQvOJa8
+ZHKCQDWBdfFsLQYdnGdEZvpJBF/O3NxePR/jzawyVL+Lro9xpqc0R0TzGYUmtbA
LCUqnEgWqV/gO8CQji1RW4SR94Pj7sUauNvIE07XPlyAWyRFmV94i+R9Xb9hjAEB
LY9I6cDkc9FhIKRf7tzj7TmH4UcgGDDQdfUaPNsrDoYRvJFCIB/mCPgf2MDwCLwm
gBP2niQ+cxypwgSC2OZehg1bK2dHZ0O0v+wWlaxUhae/NN3a8/lbaJLUVqK1FG95
6dkD6cQfFAtSwqYyuQq2t01nCjBBl6xduDv9dkNmBxn+xbBE0YWse/a058car8FJ
daCSn4+qF+ULwpVEBLdGNTm0LGFCRZaBynAAc6/S7FgVE4i8d/a+k756fGzkr0X6
qn5d3e9IigDwYqDEyksos5NOU72vbguNG9srPE7ruXJ0TQLzq83QwsPwKsYl1v59
AgnX/CI1jhBuzqzqDJd3PQcwhxkKdrzXdYEbKm6EXEqJYBJRwHJV7liqLjPc82ta
koUJ4r9/ueJSrVYAD/MWJ4J3d/8H3NgZgp9wNg+QOkf99x/lK/hqPjkSf3EMxjpk
jM5kKvxYvDzq8kh+KGimksSMN4yKXNGi/Nje7odoc9f5l0Ns+sVb4bhfV3ctBloE
`protect END_PROTECTED
