`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R629D+2ECd4FyCZ9iBOBc8VbV3k7WucQ0Vl6wFuivS7IURFtDSd4sicxbDX9EW5V
shWJs7oUHWWgeXV1BCVabj3RGO9+aC9cUS9cGFHBFAjoCpaLr90uYOi96W4mifcA
RasPP2LO5v9R0JqFO01ugC6H2CSdVA9gLYBzKTE8y7ISriU4Bh3YHmmPhEZmoxFH
1mmXUeBDCIo5ed7RoW61XgPSKcruY5mdLE7+vIbobvs3EtQDhZIkKJSM7r9twByL
bSNzLhfK8kMTCpVnlUwhxwgRv1RZ4zF+hCtqOZM1OvReiNnn7w2qDiNNG6VGA1Qj
ZmzIxMc+VbPmXqyaid1cGHEELGBkSH5IN57ItrHEJEvKEbGrLkNii6rJJ2Yn4QuL
/Zg6VUVriXmUaDOm/zqTv5DTBryoeojaT6qgI+V0fbuxT9I8xVsq5r7VIx93YDhC
G8hATwuj9BxQi0JzgRbxplji0ba9t4KvsqZiuLwzw8WcCHycB8eEr0gmzHL6fD5k
z+DT4o99An+S6fTMd4VjF5WFDjo+8ZuErPZRasI351pT2DKctsIQzkvwiu10KfwH
PiwjnSk6N1kcSvBGSF+yLCfHTA0Itf7IDSxrDp8g5TIvHxdMUWDn3XLaGiVSLOVG
s9Osh4wSeciTPesL16MfAIk9qtVgIea5Mi6GGOAVQkA+YDVOPJr489q1YBcV60Rh
2TMVNCJ8Y1guMbNt0kUD2ARziSpynAJHP1Byp1N2QMFaTWYsTADQKLqyDTGKeF+/
D5NHSiw2bM0wPWKBwVAd7AurcmsON3yU6W9LoWiPrJm+7sMriwqyaO5Fd8+ddzQm
N5M4sep4WafYtyp5mN/CkFgUGOOEJbR+WCf9Dpf9ipf/3HiPj2CjNMlq0avSMztN
jW+lG9b4rn/f6+QEoU2IugnYqflGFshv49cMove8G5ngO9wEMLsJMF8OnfyilZfC
G0Juqhjo8k8OupcQxjUYHNE/6nyr/fTVXNhoMjlC3g1xfxMJqX6SevbKmMDLY606
QHux3w0PkLJIfYznnRnsPNF+cEdzz4L2v1i1h3naAtfTRrxl8cE0hVlWksLcL4Dy
DlVvHMGJfHwQH8p9uMXbSevHAK+dq5fPC/Um5uIqBGV+nr8BKZDiXGFJNm/os2fh
9Q4yzOmLrIFWsxRMDKdymBMV0X9mu36xYl4t0sVSBVXAJrxzId1btE0dxr+ryGYc
sGKO54iE1Ia4hI/J8TO/ajlDxpl18DxZ4sMp6YDBiwnqlUHGEirWct9eu6XRlvvK
Yq++kt0o2sex4Ft1Arw9SnF2BUq6AFP8Xo423+R+yt2ZUZswVurOmo3W/8pH97jT
1f9it+VvMi1sMqBzjeC1RVLG8rFmS5kJZN7ycjE71QdisqUuBi+EBZI5pXqUxpMY
rPIKSrk8H05BZB1iq3jRJpsyrZztQobAG+qIGKlVhVN0ocnk9LLYBdIZ5yOxSTUi
vSDLJEZxloCRD7eLLu2E2TgR9+i1eQxg4o+yB5kcR0H74ULIPFoNqAaRlFG/rb3t
xRiO2tOrJFh96HK7YcJwwTexHJUKro0QqQY3/lb1ErXlNl9Cc06m51ZfsNR2zuKT
Y+4WlFUmBKpcNSFRWBGnL2QOS1KnzGqErlPlD2vzU4U9l/9sR2BSmDLJJf8qQ0Kb
tR7EzIj48TLC4vy4IWeYqp710lpnIkPkf5qOswR+xxrbdTar9kOQ3UtgCALHhxwT
J4HMv1HoV0XYxc6GiUnk95EjtAn3dRcJTY0x5A+HoWwFVy2eTRYPZdq4QjNaE/Gi
XOUAAl9HiQtsR8IQ3Vh+IZfaJEalD2xvjdDu2Zx1ou6Xz1WRjVFfPjTcpOS3dM3r
dw0BQDJ+J4r0rMELu+FKzOTOghYVJWqZ1Wp2WRlwpQwC0tntv2eolye7nD0WPyfR
0Fd+64E13o1ofGKNBznJef+q4cXU6pxVR2om3+uesyUNdzALh9XsFNIBc6iPjr1n
VLtnG9KnxFUlhyOUFVuuww+Ovt4IQm5c+PirWwZg5ln78EupkiTZPA+qSEPMefhm
JW34pzP9hh+IgKku9/wshSfMxtqQUEeRginLI3D3XrHAaevEgulXpAL42RydauZE
ULp8HIExUjlKYF89NAL/bZovuy76aikSz1pGhx3k5UUEYam8LDVd7Rxj5GdFd5AH
dP/NZpzOwlBBEJbN64CHEJPEwvEZuox307Rrl3bVLRvzFH4izVEaou7GSY3Sb9+q
37jkPqSnQxHdIsdBnvydkpYs18nMRAE9lFJGVriqWFOZ6q+5Z9QWY5yV2N2rHSkq
xaC+XZwt2a89+bpVjCEfh414m238nxgfm1ZrneuaytFQnr+UShpKPA26ZUsef5Bi
Hj9Q3t+bCA7EDTxgDyPMTUYktNpBRYQHUvTtoq9gK0TZxMnW1NxAjb9M2pEEkkR1
zqD3EEGFZ1RMiZmQg2jYFlw5nyq1wULAGtiWDd6Hm24nd5myoEZgBNUujvKkBbjI
p5YW2QoW1C0Dqn5iYMv3ZTNXRgN8HXg10J3+zPqI27dGBTm8dssL6ud72hPgYZH2
c/qLt1IY+3Gq578SjHaeoqMtBV0kIs32WwvAcG7nv/bfP5cwy1iJKR3wXWhWqAUE
3QX3CV50ZGhN3GkG+cu7LUYqJLQeXXcpgqYjCeq9UccmVXGXwdc0DyKoMJZZDr8R
W+qvKaO3YIquTFJGwsPl85bITvISHf+3JsJ9+302yrz+hpTUGkOFDRSta/KtAkqZ
/XhIuTsao5gGT0sHyR5uLk7vzMPSjxbKvOfMrwvP9MMDU+DI9btlYs7JxE9Eca+R
OUDROP5J0eZcM8KB1Q2d24L2by8j8oo5rIgcpRgahy7emJDCXM3q+nIYQL7QxJAO
eT4+J+3jNCfC9lBz3aYr8/feCqh1gb8uTNYoTaHGfSyy+g108uLul7aqtZfu9l30
7DPrfCt7kyjCN3DFmNIrR4ln4BDEVSFpqdDWL7aRsSt5S78AETktp9GH2ZEebHJ4
few762zkk2hGx9YZC8Lo50D8w2HWS6kqeHj285gA6b9by4pbF6mRCWN3QNGp50H7
0s1yMnX1DzEOoyt42ogvieNTKoisqhXrnjANCV56fk2Dz+jsnAilPoIHq3+W+GKk
yAT767/8DMLn8+7fdOrL9mgSlc+saB0VEDmL4mVkRHKJ1okUewC9EJVuCFXSRxNz
qf64D/iGRJZq2CZ8oG0frOpC0axk4My+z9sk7bR9XBWZzQPuFiNeXdMwAmQdgwZS
ZY2IFHIkjVYPDhpO6k7WVf19CSdJCfn3gAIx6ND0PrReoYwT/AeM/EZDSIotqz6Q
zETmMxQnx3hcpNYah0RcxWBez7MSGL2DLPXt21cDXtvkfxdfDUXjsIQ0yofl71Y+
kL5NF8cNTyGc6z8y+bIKUwamkinTnh1LHNXMgPak6Xyf4/Z5RH0JDqKzpmxY8ZZ4
LftFcjcmdZ6dtQksZgRFRDwApbEU+OJM9RvX2cGGoWef1GcB8l2Dz3yuey7OFQS+
0VeNz9SyzxSH6Q3Ok91M/TxdQlhCgx90BPVsfFr8pb3d3XfDnK/NuN6X9f9zpEms
EoZTndIA3ERA67O701EVYEWUFCFY0zjnYlKC0r5Yqh/wFCHPo2bMmsrVtX6lMZuZ
2AFhSt1/0d6jdGP/pMko66+ZaxHEnQEq2PN2EqS8uJ09C0RMxLGwqxVQr4yrPvaY
wu0jPoKH2NBLZ2W+9ZL/IbzIN0kJ+TJF5+GEcDQ/W0ymb9KBkxAOSbhnGN1kqzkI
2Hjj5OiA66rMJ8n8Ot3DsXrNFGJu2NEMHRXO6AoQOMaO4iOckU0q9kc50M/roarI
VoqW+UTJYuChsC2c4gt9WJOoRr8NjYn8cWK0DB7eTPgfyP3oQj7drgjmmqfuR+nP
Y9s5tCQcINx0lu8UGPtuED9j0bPUNwi+ODIA3zNSEZzucUxSmGzKPzUmTppORnvy
AiPebZasxnZvxLoqFGaLiBtFT7zb+rl3D6kBk7/662zlKmeJwn7GEO3+K514+YAo
YsLYDQ5Fz33GCpCF7u5qmBq0U07CGGCUqqHzfyg+tO//XS/WrFfAENljLX9kjGRe
N3bbUgZHS23HbNiRGoOrdcwbpxMe6TqpZE4D8Jj/DtNer1Onz2J/N8JygNqiAduo
LZk0ZXyvfutCW8WSSLnPM7GyW1WTJf68iO2xo/q465FRNZtv3tdqFse+b+mfiknl
AYTVJWxy5urGRH4RSTV+qQFuI0t8xlSbUuGFMbxVa7mG741mZyMd1xXwyFG9hjKg
OWpJmqfqRm4QgizC8xGHqf+AkxQ+63Cem57JSiA9uliClbxV0qjL4vJwVn7BadsF
et/5EfZ4YWDhCYgv8xSeBun2PWQGc+apn2RrrQapPFFbn4278QRrf5llAP1LBS6e
3LNzSu+Msq7XauOZHOjhErEhmqdx7FWsh0Fm6yoOLdKF8oTu1335azGFSD8bUSle
qOh8ITNfkZrcid3CqoxrMsrtQQka/IM33gLolXbkzjgDLLu1WeTHI6bMxb+cJ9LK
5wv69SsQCL2RznjSIZqH8SQNmmKfBZWgCogk5qijQFbagwzsMvsXWxwL56ppEPNd
6Whbndhd4TRb+jw0mjPPB+0zkDoOGiXeOx5SSxJSDPctGHmpQV5zoXnlhrB7B3+6
32YLKGcehqKoFzTY90pZQ6Gw8MNO/e7+oI5GTLAFcSoj0AIjjwUTXxFqf7buXxpI
l2+nDYDvtFKXX6b5nUxV2Z7px/XhwUC/oSfLmpl22iqoOwAH50SUpGIzSC7+SWeb
ZgHZHTH9DwMRSfOSwOjonAyxiN9C6fw1abK2pC+BVgDGPEWhyyspcnMJ6Iv36Pwa
hme0P1Vz+GqGiqMelvQV9htRHv1+2kqKoGS0Oe56r8k25C/XTDSNaK/rpJ+a5S6C
gNpc4R0meqODMYCh9TqGO/8GKk4yDJTuIUhSAFIy5P5BgmIJ+Wc5NZkomHyAPPOs
ChZoZvPbHiKR03eQ8QA/PKdNOKI0MY5zcsXvi2u0pQ2wO62KpFv1KI0u4/r9bLJp
59K2fZNASibLeO0FPgQKogtTTmpKC58ZSYzOL7a9bFHbr96ibVMa8PWpdwoltohd
qk//wZMnwKoYXWKoQBhs6bDAQ5qahY60s5FLoytzaIW062eXTvpYTWldxSqRIwiK
aG3xIq0b+NlW6k4933+EZBCDbw/OnGNzq8rbyAsQJlE2NFmmZXFHL59jnDHEAmyI
HZGKMT7nBjyhwKBbAFJ7j0xr7opGZfdR0Xm/kkFN6kmbZq0soVltSZQlLKbMTjlS
Zb5WFdo44ipL/YM7Ev+g5E4EMLLGvXmXkkLi2SmSPvj55Pm+/NyZD1FuLK9STVnM
PLQtaRu1gKDcqHNKA62vKpSk694i/zIcbanjsOnmarq487hWqulup578oN7rZH4/
989WrVzYem4jrlk3iOKYa0ZtbTUVN3PsDudaKzZ8UWurgrYTuiToVHD6fTIsDkgl
0lSEYG3DHtrMiPmStk9eW81SOAnJj1hXYwluoqYQ4qaWqj9hApHDIVayGjR+opkG
/AKIkZ18idEQd9JBul8+i/QyhSAv2yiKHmVTnlu3GX75aVNL7TiKp6CZq+Qt/1tf
FAJHghrOhuGpvVOQJOTWHqEbawMxS6ltTMgsBpDQBgNWXwtcP6jZ15/Nkmd4mSUE
`protect END_PROTECTED
