`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h2LBowmA3fYRobgrzShLdoDRx5i9NQuyVuKP5L2jNNHia358OacA7izLCdZ9x22U
kc+TTMIrb+wFlLCRKs6EbBNt9c+8w6CRcpa5nGYXIqfLeALsqlqvuoRfwq+7XBFn
Zvdghpd24aYRt3dkNPp7NsdiJffbAZoJNMvLB9hr/dqE9DHUFr3Ac+uRd7j7/h6L
5Qtgw77Ow+phwkHXaJz+NeWwZTBfX6AnfJBsZno5dOzawVoahADUrvoHZwpc2Jsa
/fhCtHfPM5bn8sAKEWVMdEdPDabLn2oklsWMz84r2Ud+Acd2IeQ391aIhqYMIUHg
ELqTnu4Sne4rILG42br6g5L494TkY+oaT9GveRpiEWfBdlkBsKQnbwAYDRDu0DY1
yVVWi1Y/vHIgJz2OEQUxLAqkCpSfcqZ9RvLoCXqyOy7e8RmFm0S09s4KMTWDN8cG
AN/nlrn3OrvFNsbFXSP01YQbrjNHIBn0ioDe3KKd1oKFiD2vQrI05zPphrpjouNk
bH9gXaoTB5gwn9eKR7s5ADCB+zLfxYyVUAm9LdVzylyxQKTTN95DMSAnJjQQD7BP
Kzq01c9Gg16L62r70wWhVE1PTXAJ2LGFeUF4eYu9mlRiquZ/min84UYH/VlNCcUD
hzIqJzwVPN9pwRgSmpHA9MNmpf588AIiPrBZZVGvdugHynqxDixY3l8IoygDScMK
xEH37cOoshS6WLhOchVPQhRBLElDpPqIUMPHO2kp1TnYXfbT0a1zLOSIFmyF2A7K
iZB3AZphmxo36SAC+mjSwnJzrk6dIGc5OH/rxrttvgTegMbZ8+lk+7TEWl4NP8pO
UXJh87ueLK3PWZ3FUJySC72HY+hFVQftBq0rkebKOJMusbpH0bzovsLCEfp5gA5c
HBzWHzdQ8/YHvLmEMyF2ZkEqAsme4WlGBJviuhYBVrgjAqvPeh1zXox8LjLgssPf
`protect END_PROTECTED
