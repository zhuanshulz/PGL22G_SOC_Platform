`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U42SAwcsnA41HhMRp36sI3cfSIE9G5CJVJTV/w1NzhzR7Hz2N5aLk6L+UahEs2Ka
sItJ85/3M+iXk7tH/JpkMQCLuYnra/X7XSe3BjrJHO8erTHELHJF/nnkIzDpZlPm
7Ki1/fzLvvgPJBdcpEQCuATbB7XJeYWX3Y67ZtfhYsxF8cGU+FwGTMH1x7+5YbcZ
NkpLaCjBIgHNAxa9nPTjMotRM0JoBnSKIvqfSMExFNj/ad1cwuWEaC5qn+4vW6Ec
phpdeEDOac9TJzvYbgj+YottOxk6Cf1F1aasg+N1GNQjzY4jzM2HURKDdZyvcsDQ
BfkhNqn1Uw4RgnnRv69KYcMwYg4/MN193hRid8hMiK53DA9ZLkM6RYHHiLIVTwdY
xFelxDs287NSXzS/XzPV8uE2CiznxI5qM1Bm6v/3nR0yR01U7EPtwz9wSHmpHN2u
JrIZFkP25nihfopAnGxUhIajc5Qi9JKC4Wfh/HaafOdXE/jcaSvkDjnEqNLFIuCT
4TrW7Y4H7igDD+Ab6ZBGSxqzqdM8aBAtUm+7jAVSDofBU3Ryn2KbnDQSTmxhso/q
SPFCzGtxJyzMXnG/dM5duFJkUR9hvaVW5bmLbfugRdwgHTboseGe1Nd2TwhLF9Ey
c9XTFc4VT+47TmclDRhuJfTrOEzCOC7Zeqvm9M4Ek2HaHOtWDPRW+0JgCPBg3hUT
GQ4ulHk2nppfb+UrtkrS1jJnXeyY1DMhwhhHxQ2yrx7B6/psDTbLyUfCM7Pa7/rd
lEOIjtpPm4rMhqOWA4dA42iKBLqFIj3rlLDmWuIlJsTrZiNqa7nf7SOWLMXhdL18
mmN2GfcUSVPMjUAGdl2Xk6v71PVMaZeGhKEbnuLeElivXoj+4UfcwK+GoSzcYcwi
S831R6o1KIIsU1dtFP+83D7G2SEYmMme0OvNIr54TRM9rQfQ+PMdLNg/kIk0b3RF
pAkQNaG6D90f9jsr+7LDyg==
`protect END_PROTECTED
