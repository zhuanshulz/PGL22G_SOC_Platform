`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vX65HG1N86hUTxFU/seOwTuX+UKLy2fSoO6S/2E5ABUBRqb/pzzKQjsYGLfyZv8e
lLxi6pqdB1iShtc7Hx8k1R3Bj2nlTc7XI92nYsxZ+fkwXlFJQ7aA9L72gqw4xmjQ
fExlstssqFyC2zwTo/PDVC+tVYqUO8rFrta1hstYG9k2DrJIke3qNUS7fazgExLn
Djyf9TyVKkZnBDK3aMfwrt6ncPvqUgF8UdxQcYxMdgT1F/grp/driipEfPgtz05X
HKJ/dNAB+lqAJ4B327xH00MAMGi525QRPNoCz/w8C32d+eUjn4d466kfxz20RU7k
LP4hgA9PHhMkyeRGr87RFC5uYu+O57geLvSiFAeElC4j9Zm9NA3rfC1RY3LJbddw
M59bDZPFJaD0ZhUt/zsbZwibM9J+2+iLs1kma6zpzPRdiduj2o6JkIVxiIChOx8y
mNaGs+JUL0g0u0fKen3bB1zpm+cPrGWxAM0cSbFGw0v1M9G8K892nzYmvoEDPGXx
51yCdmnd6bUl/C86aUJpuXk0tEjge6fsbcbRrEgFgSW0Z960/2c46Cdq58lLC0Ms
y1jCMJjKDieZoYDu+xIPyiqvRJdNctjktr3+WMBP3crbZ9TRiCNYYLAEG9n8gTn6
TCdXLTmrVfu70MU1gr1liJPDrYJNT3/yq3SO+jmvck6pDxQwxUI2YvrB4RzEyAu4
RzIA+tK2Gs7lCOcGeK2skXV33GaQocY7M1o+vP+ifCD8C0nIekqNpMFgnv6/XaE6
PIsAZ7hFDC9Sd8iCkP3S4H8i39bJrRdxptXv8IcrJo2NAURI+bUyWtUAr1Y4Xnr4
dkHJjEic3bOMwpeCbJkx7kqsgdVOxE/z57kaKS/ZKUAH9fposCs+hW1/uS+NJSFA
YbQsnTobmkXjfxVgz7tRqI5xluCes5U5shNd2PTknqpQqvJQBXhTjf8aOEGPEvde
QJjsvbTcvwAZMDL6BrFZN0rzMMCsMPstLWyT5ZtTSVfRVCrM9fff7hI7axGjufgv
sdXVUnaUen7GSVbhiVkX5Q2AtYtccpVSxr8+H2soUYVCa3Uy/l7+TtYSZOScikEx
hWCq6NgGl8rKE6LJzPdEYoI1WGdC9ckqOEkQoEN3h37WA2+xl1z99l9CFcPrR5R2
/A9CIn1LmB83NMY6pePGcwotjPttPv5aND1nGhpw28XM6FzdC7ejvBQTqPqhI0a6
dHpswc8gez75NWXs4QE3GbTuwNecTRanmexKbJWOGXs62K2kIBHvkgKMQQvSZGf1
eReCyP+P6Osv1phPrnz544hDNvfxm+qjNRCIrR9IEsmU5y6R4biKj4MVfeVLIdc+
juRcYgcYOp1cJYJVCHgbth2YpKyzv2FLQOiQaaaUFmhpPPnjfEg0ST+oEUwPuY76
z/vBPEvrpAsLdLKAfEAISe2KWbmpYX7CQBGoDgGEzksiP5kcMk43nrSZmdJHdfqH
4eZRVh1WFeCgUO/IP3KWkDWm++zB8sE1yCqmgS+/pdY9+BeiBKkB40Mj0Oe8Km5G
ia/0ibjg/5oCzPGshwYvha8j3mphvzh03nYuHqjwQAx8RkUBt+ynfVSc9JJSgIGG
5oApxqauAcXFx06UgOXez97cxTzFURpedgYXXGo6eZpJxCjuw9SeP1+jXKQDkqha
DMrEZqiqHjVyUNultZ6aWxC+r71HUbpdsR8SsCnIKpiuxnevNyO3dSGLewB1G7JD
CSMkhUXfSPGC+ljUjmNdexyN92yZ71HxOKDHrpr1A4rZGs9Giv9dD/5+/PoBjXvD
5Yb4EwWUlQq3OuS0yElwovI146a9bSbUIrjREEFmscfmQVNzzhMDNvLu/xyn9HY6
iOgrrpgqC7BTFnTp0ty6A+fWUEV/uR6AnkFSy4fyfsFEeccXCkXaerMuPZuLv9Mw
cvoQq9ZGSqAkedl/Lug3Gckq6udGfwFc1QGw2FDakXrdk0wJUzU3ZxieKOQ0OcMj
RTbD38h0MxKAjSXfhNqPJBgUNIoYLjBxw17GiACWySOzZkGjyYY48nanuBJkX+uE
5W7WTjAwrAw/I6WKeltE6rHzNbs+jNUZzwUeKVlhlfFa76A8h7ftG09RT3hVDVmp
338IiqaDeiducclaxADBpcsUwJDftKOmRymvM0bGjIFdsla0aGidrj4GonCkl6E6
20UAqXI9Thzxe+7NATMo8OIRK100jaogj3ToKzBevG3tpuayapoPJvHY0zGQgpD2
LKoTyUdy4dVKMHXzFgmk6w==
`protect END_PROTECTED
