`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Fmxgg6kDN4SnVXIKMSB3exMfIWsLO6rplBMPoxTSDqmypwLALMnTiNp40yUy7eKV
Ki5ThJqCTLaEYbWBjW8cYgbskBUbuE1CJ1jHWDECsbHY2s/dw+G1jTe3aGDb9vK3
0OrQyWBaA6sw9f6bnYbxeC7Q0NJMFap3+9sB2qYUE0AU5FgmbVkL1n1GVu/EQbum
wuo4wsXKliXsnXJASJZvTNcwTiTc4ZYzXSamLASOh352VTrfP3Z4jiSdYP5k9+8G
JYyewykNW/TlaILhtVrpJia/jYOVRbfgwyI/oWG/RkdVPW14mpdrWTA7/ng4qMDF
mQuTOG9KzLoQP3IT+BfN/485MJFLzzFahkK6IiBn4gXWFrMA5ldc2jmQAWfv2NhD
ROatVhlfF1oUt18Tt95zQVmiQ6jjD6uXA5iReEnYwwNoUaGuPYLnpm0mBldeFO/3
tL6FxfT5iinRLc267OHulq36SDCTxVubshWKUfUPlYX6iwIgqeYTuSxaizmxl4Cd
eamS6wk3gZ6T3F8LbHhaA77fMlZ3Nxhi7sE76GuwJV7Io04qwqstchpEa6jQUAMi
N3t6tAkSyBVxxjF8ia/KxuFqTt+gMXc3sZtonUyq6ivMQuz7yenHI7VnhxVpbYwC
rByo4+8gCQEr+Vo1z474TS+aIc596pS9+EGSQNXrKrHcA/yp09XhCiLmeR7jyWE/
fVGcx6zBjboQ4TA6oL2fWSuLwDYkdM49Gpvz0MQwSugZgoR5lLb8fBzQBlC16XBD
i2aRNiuw5DmC7y1BZxYapV6fsVLLddp2w9bqrAc7jj8YHHpl3Ot2ySeD6zI9mSU2
fa/T4XEXKZns7kx2Cck4lVnVvbCwYXMBoLgsZWRsPU9wus6f+GQFSKhFp1oDaJCe
xm425dch4+YIBGt8KhZUA6fBhGZkloj8TouQCZalg6konyCYmZx2Y0rBO+WfbbOX
xPZ8xSX5KwYyBBZEdtnKjhnpwECxcvfUX5ahk0W/T5P/wxzhI81zBaMJ6wkzC0jl
3xEI4DDMlIwaCg9/NPzkqfQG9bjPDTP01NAa1YjV5XUG94nSthIH8Tqp2gqlGbw6
PQ3YZ44RTF9iYX/4f9NNRBSdqzXDZONlvRhQuUzp+bIA6ZwEyHSi1XO9ZvyzpYi+
ravUXTzt4B7xtcDXcnaLOJFfAgmwe5CWq8fej7nKjPY=
`protect END_PROTECTED
