`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HixEVw+JTOKPiFS0wiMPF8wXQvR7WYJeYO6vGX6sE9vcAqpFGBd1bxO/APs/g5Q8
Zvn8DvMQ0PfdYgZeULYRz22G5oNmG3A9taPym04FExYTjmZO/dveqcXtYz/AmwNL
zkRm6Q1irqXD7v0jXqDoxifznljr+cPlzfgb7uUbE1uI7knBOQV03B0k9UY2ioyG
HWSBgYvGUe943JTBjmD1CCXlV174wGPtug4mxGynyVipBLKYKuSQaKZml5Js6Xw2
XfIxXoLhhA9Gt/cOIzrG+ZVYkAHmYjVZa0oNFpvH+WMKtJxBQKMnbRtxvZzniDBM
zOYwwoM1DAi005HiGscgGlmaIAFYK5wGfeuWAO1Xj46LkNtGrM3I8dR9WyXkSr9l
b85FZ7GuDA/sj8F7KNxA/V1DcyBqYmnFReO0ieRgjcirgc1fAZ9l/52pp5mRFHi9
zor2YlWEAci++atDL60kmuE9Kh0XyGpOOp+hgiJsgAOjYooZBpJgu8h7lIRurHl8
nFr8ydXuPKioecdbQ1W//sedZ6KJ/4eZMiLgw8u09tzBea8cx07hhoVyDA81mRWR
1rRAIX5EJ05K9CG7b8o5DAU5yw9qIasA6QN65gIh4W+5hVWutjUi8qVFayKe5o/E
1Ujfm/AanHSDLKPlYkXjQUHJGKR5Tl4xu8CVtfSsUheGLk1CyY295nsOhx1fYuT3
YyTmcyuDZupmho/wlwlyHYy1uJO2TYPj00zngjJaqNsadidJnlyl0cMTTvKNVfrE
A4Z+RSI5lzgw3uSb5twj1IQfa38cCO5x7ZAWLAhzpVPh1sVKvmrtEHDpn7ubsxC1
g6o6amacRiA7vgQEd0WUoznNUnUKgye2DveVDrCOsa6KEA1EKCuW3WcqKCGsKGJ1
uopQwRTC44TzfO3DzjXA8t+ldFLyxDbaOYLPVyWx3yPaDe9yu7LHxOWs3sxp9eJO
fn2rJojzosxWfoTkjhV1YTKsFu0BbIu2jzqMfzbn8xHwssOAZnhP3kyh84rf7UuP
zI0iseNnMwO8LmWYfuQxHNc46BKZo+Bd4BcXsR7b+QAHd/U+H17aWCPIoL6BkiQ1
jxejgqZx2WCyxmoeIu+5e0bKW8gNhb0WugHtVitE7SwkTgeCsNSu0QTeC2lSFvGI
HT0AeAe9uawMcMe3kHoQt4ZjMH6lMm6mQhJMIlCfcXk=
`protect END_PROTECTED
