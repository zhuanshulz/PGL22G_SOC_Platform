`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
upcNlKS3R3BNEoQ+7lSd18yLtwN/esvEsdgtmas+ng0sBfUcRT9Rt6T9TXCVUj9e
EKmG0Ahh3Tykem00xTeL8cdwzr8NkofOv29L5ZwP8GUNokq9ctzfeYeUMO0yHUNO
8Dvtdd3DK21ISfA4D0SvDPBEjdvF0GWDeRlAnZoAmlQoOO8HCKzfcR9TMe5X5sQu
UuuEDTXpJL8fLWXZvup08/7TtHKCfsWVo+bN4SY+4Of/sHNp7ltPvEeBx9WJ6y4v
mzunZ4wWKouDWlSMCERjrp+/+r2BsSoroHaZC30DTw9Q9qEGlEGW0iBpNS5bas+r
obC+P9Pg60J497KS0SE+29OPq0kr8l++g0jR4G09UkIypK/olkYzzbi2vv5fngLU
UKu5KLpNXMIXFYmoAJoJ+TbrVaNpIbo1woArGALa3wWsRCYxAz+cIq92Zfwo3DqH
QKTE+N0i/0BkqgLtx+z4iKeuUULW4dlY/x9v+lviqvkkPGeVBp/oW0ev0fYnWtB0
wGW6J/qfkY6z3l8/oNcfAXkUdP72WKcLA7bpuX1Zq8ghh76sxJWe8QxLdSeJJ7PF
g/J3vIPAireA/kWPXxf+3qbDVoL0EEjRH7hMZ1IPvX6qZvJ+nndaeUmtGdmctqY+
YHRSlgGENt8Mveu1KmtVbaGjI7LI6s84u76cemXY8orZXeD0aV2nKyG8o0PHuK4u
1QraACYGabjYJ5/fDKtTp2wPyG42vqhpn31HmYyh7GcJlF0WHUU+KSGyN4XjI+AQ
cIciChXHuF1t6Oh/H8Do4CZMNlAZ+7ZXNNmd9ponrkRpapF50CA12Oybvuf1ns44
GaRhy/eB5IbllcNxmVf/Mi6vyYoIVJuGY0pUrl9iiYmkPtsAeRgKIQrY8UN6cL6V
j6XXefBLJnEl0uvQos626bdIdWMYzPMj6YGB0dRzpohdbLzEZmyP1RE6oMeJX0RZ
yuv2DE0Q2Lk5RXQfgLqlTQ==
`protect END_PROTECTED
