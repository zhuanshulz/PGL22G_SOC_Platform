`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sawnhr5s7kyNDhieRyRkLrdKCtSdnhVOCwIygGBBM078ZQxc0DNxlyOtKa8qyfQn
4DYy03ULQbWxuSPyt2u2wLxf/K03iV/KuA3o+6kPUyz2l3jw4/ykpZqV605ugpSb
jlWgQv2YvoQ36PYnFXtzuCwUIyIIYS/0tWl/udJZwPrStIORXCViouIGoQxqW9TX
wCVK8Yerj69B7O3xk6LaWGknIYo31Ewh5qTEbOmSFBcYLYFxH/hUTI+kSqYyt+JQ
ysAucUyZeRt6aTZBt1Frv/e6fMj+76B6gGfH89jNIYF84fsj3VbYdEvlQrYGC71h
awA7rvC+kTN2x4wWqJoIlCTIMiFKkUgC8C6oJQhA4hgHGGydEw2GU3i4F7yCi6qL
wRAA/K6WTVa1KTkOpwUBVKByGu/Y4yz1JsBR4FFOvlcRLjw3gdb/DqgwI4BGXsM3
ITU9mPrP2kmVTz5ttS+xNNKRbBpCzJFBaDTJIKYpb0AW5JmOZuxuhAZNhVjDzxXx
flEAm0zxAyFIOr64yrKSB4Pt1trHAnubBCWMTteYjW8zq60utPCVzZVGLtPcAjbu
uwUGTou5mrjBsYRV4xR/9GGVwcSt8zHO3JDEaKYkcbRbV0eEgG89pYSSm8rhwDtX
Pok9aKvkLEn1zrj4EDCyszq+aMSNRjLob2ZMU+qZQW3uiLO6qH0kERctoOzRn7J5
+nu3XOW//ypvz6vCWsXoX5jkxsDPFzLp2AR3JuhOAor0iX76+nlN6mJ+QTB7/T++
ohAn5DHO12UV/7GJG/0Vt1ObV/sbet+wovbHJxfFANVjXtt94wlfy3cNl+D0yKWC
RcHDW5rwlHcA+tDfGxcv71pkxt9pd+Dr1ld+iqR/IMzaKY8htHzIDDn8BWySE/Mc
+ySTaXnBTTZt4952jQF48kCJoBe70Q9Fk+zGg8eu2HtBGowViJg3V7XZIwrIwn8Z
gSmINfipAbXzPRZUqB/k5MIIv+r/A9dpqbO9BYl5P0YjvW6okqAlMjES/aZh/30h
93xmfPmHggH7NwfU19tzpupBSkx4NeMpfCy2i2Eu1GxvUcknCViPF1gsWrSuXWtu
7LgtFEE628OIhfL0zuEUzLXSZy6OqczvfpA8uo50miAHFYpGFAqLc/2MuEQqV7E4
+gwmqNyLf+OW2LZs7efCfv/hwFIadpzRSqy9oHcDLnXZULA8NcT+W2kNY1Y7foWL
hu6nitIQWSAIpnCZSTxMJlvFHQI2mmfx/5XjuLX6j/Hq88nu+Yq56YPLApRqNdgD
pcOcju/TxvqXGK+eeEGkjqakFTAU0zOOA70959dsN66jc511GIJI+Ds4ZWo/xJWa
rtL7BVW2ARJjQUKrgDtiBfJupbO/24m5kPtUzBTB1W4WI8f9rKXl34SKFALpxn8D
MQPgrLlHmeDFitJCSZCtbYN4E0B+3H1Pb0a9lW9lgK+tUDiGppj6KpCge6OzgULq
rIx8MsBNt72eELIOkLNP610ebl6qZPL4UOHdVK+lblSNKAWO1VfoermJYVfUsiZt
WCeWiNY3mkWDO+bs67JUvmA5MI6psRgTz5txNvnZSoPwf+/UrC+A1VoJwn4JcM7d
WjlI8vkdiJr075m2aIBAaBQJZox0ED8g2qZTglma2LlBW14lBmx5jwmzZ+L2TwoO
Jq3Yt0nEQDMrYUMdFeHnvk+Y0folQfL0H+/typNppzoCopOPU4cgIznEyHaUP3j8
PMozJolaxjSzxqHms0sXEOLjBBO8N8WKh9Q51qZcn2G/LHHqpaGnR2xPn/0bOaPx
RI9+gmP7S1ChUEOiE6sNOaEN/tr9fNkShR3+lQ5UJc9oqJc+KaB9kmOd/VThnB+R
SD+OBf+3QphoptbGQvFZVA2Zuq5Me5W75x9lWek1kKIPzAeWp1DQlz3wpeTNfgSG
40BUg/Y8FCOnhDlRZak/1+fgeSSAto2CpWYjUxhrj4k=
`protect END_PROTECTED
