`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C5gkwLkibAEYif6hjshDOQgjL4UimOtBZ31jq88IVRP65nb+2zYDXy3HVwcjISZf
gYYb6YmteLQJUqSWs+LV3cMZy1uERSTCa2kxUkuxAGa18B7lWSTSpx4x/zH7qsbI
9N56ZpM+GzFa2sbXQuc6C5wXaaH5RTdCP1oHwMuQ094rMWHsqMk2QSCpnkpEXW8B
E4GVnkuYEq6WyBBEiThYUNNjBlL0l9CbsG9lBp/cXfqI4l5tOKz4jN9PoZZRUBEX
PM8L7sBbSCKJIWM4TdfiRbQ0Ui+QSKj+1rjfOEBAMYC1C1BCt3taIh25TEBf+2lO
Z+ooFkw1LY8Wj0onn+1PHt58k/awvVVQNYWXCpGfvJeuA9EN4B5u1ByySKjzLg4V
w3R6rX1y0erLv4wel2zZKTPaDMSpvjj1MRKWfcN436DmgmEzvi/f/IrYl6DfDLT3
jCxPuujHqaUyTyKo3EQroqPQRUJSUqWJt2qaBmtvlUegsPTCLwEVoPHc+B0U6EHX
ehU3oc0CsUkLWtrV2hdFt+dOthATz5UIyuvSrHlPuKCU3/WP9mnQkrNsBBMBzWUg
yXSXQz69k6h1lDXrmLJE5/WDm6n/SSk7FHq55dbifHUprfKzBy4blwJ/0KQHtZ5l
MkzBZ+0y7nXpwo8EGmnOMKqGpEk7uW+D74QvGsVOg4SjesQgeLmWAdRTYtKT9ALa
z1su5aedWJ4j5BT1prLBnFjDYXXQJgaO/TTklv3gE82YxgCiZ8msA+jI/zbxFdzb
IUuASLHZAcaQClQFuXEHYu8VKnQNS3HYZf98sEy5mmfzwPMrgWs82Aq5fo4uqgPM
dC0wIr0LTnFw2dS/PrK6n1oQo+9b/unLzG+RKyeCE5m6QvLnGP9NPrXLEdJt0EGJ
q5zoMCegjDsPU5EXgfUUFNCJcBtgWYzQ9EfiDaIF0cwopyaXgeQxe3kqHN6ql5E9
P+c0lv5gidLvI+2nNeHnS9ygWjeD87oqO7Hebmh8j/1E/Ezuk8V3p97UZN+jvuib
wgVHKZyvneqR3jTTtIEO3ClogtEF/wnXnI1UA3OZDor+AxyBEeP/7L5vGwukKRdE
RFTgK8own95FKKIupt89BuzyRcxIsEBvwORYGGg3p0svSG/6wFdyx6hTqGk1mpZx
7U1cWrlgz8tfd4kbw77T3VwJrqZixbdLiUB48qpXPc3uiQDto011+PxhlmXNhyAq
0NCPZUaEJn/8gNvAGHzKIHz50NWoXBd/Y0odDKJmtZu6c+alrhmWVqGZaOmPI5E+
Hq+UO/mCLfqfmgWt3iNHRP0ruQhDPESSVm4xRNdTfnj4Mm+S8lkcjMPK6BkDpJuh
C+rZNouq3OvgcEMGNTFB3DO/jMUUxF0jYfirgK5fw1yBqnoYdbNSdR8m1NHXcf4X
vgPakmLtbtI87o9+pLOFpM6Ox2CF2wdgK3MT4d3twi3zR4tMIl7lVCr2EZyjwE6L
lKrJx+o12BjKgMC0SKJPEQ1QUHwwk0zLRrsSsdHM7Vz/uoTk4JsDWToqcJ6xie/s
ZKWoex86iUpnb5p+wHb9W41fGcGS5E0SySQrV3+1pRWio9rrmyfTjwv12A66NGrr
tSu7YMHgQofTNLh8g9JJwHowIkjMcMHd4JMhGvNMc2RGkuMVVhDRQ6k643oYDd31
pOJAwfZkHvQfD9iUppJuU/D2J3j56rL3cdx1nDY2fZatGu1sw5YCMqg/wQWLUKJa
PYWhbkJ8faH9u+cy2eDB1m1f8ZWVDB2H4OsYpAM8SrrfxXgKDb1z+DVH5uZMBe4c
rt5tmkpso3BD15INx/ESy26lIv3/8cpzwP45KyDVB7m9ZYOt5ANUXQGnZLsx+gW2
jl2HV8VyQd63Uha9+rl7/9uoe8iCRyKBsHoF+8A4t+vejdE2Ur76UYs98UwhW7az
DDBQsR3Cz135cvANyw65rOngq6JIZYGEKpwLQ+ETsMqmU4oXOhXb1FooGeVNicM6
SYkQQuqGTHm4GE3Odeq4vU6M3VWMxCRCdcI1dE/sV7FbtgpjC4+c15xo/X/5WrIP
PIOeVJ+CqPWimsgAWtMNvQ==
`protect END_PROTECTED
