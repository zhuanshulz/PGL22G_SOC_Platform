`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I7HBDcsm79BjOEHmfuj695WKLsW78qrcwH5P6nTVBQopkIA9K4nI10cQhk76VgMo
GrRHRiSMmcmr8HmEQ6MGWnBU4QjWt41uKF1swfe8p2NuY6CGcaLtDrI/cjcOyZn7
Qt0eBpuB6vuSK06FF0PP4VFJgDM1Yx3tt8G/f7VJlfLHZZAtF8GON2rAj6R5ykNH
hFAh3FVh24sNTeRLM+APz6vuJC/7Q2jPkmpR8HeCp2Nlm4UakT13CsfdQBSCB7cm
JrfuZM2QeeCM9tkN1+2/8vVk7Uk0oTIQ8kwwJ0JHfKHLH3lj3OnjMaDZqa4McrP0
jTwF/Ya8gKB0ncR7B/LljgsgiXqBRLlBrN7dJdiXYsTULmvoyE/vHen66l/uRYsU
whRJF40ABy9v/GyCfXUxDllfZNK69ERdTH20ILv4mc2s+WXZlI+Aev88nP6Y5B8R
GFyOlt888hN5bBVcGP7D/0aUE8Spm53iwJCYYYdB+ooAjmbzuQWah7xwOQUUehuh
ISIXYJr0OtG9bffeOLYwaSGPu5dMPqlAgWy9EcsHb2JbA8snZpllZC/YOvwM5O6y
rJJQEmsjua1DuP6a4W/b8w==
`protect END_PROTECTED
