`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sYYglme9QZNR2FOlnwdvbc/X/X9ncWCcA1ZNOvVJ5djjmkEueLVAJ8cTmiV1C3AI
Zq3P9K0f9lHNqYOQG8X7h+AjSklzEjEWDn75RWNF/xt/r3glZMOvnGJJ8Hb57Tyg
klBb2xy/dV8AAdV+z8Kl/IP7Rjb1OAeteRgClmZzWyQxP53k2K7me68p7fVbxrx7
9V5AzO/IN1NI0g0/leIo+sql3tGhyNY89vKVhm8X9JZIo9ba4M+GEzaNo5puzVdK
acPVY8O0BWlge+L/FB/zeZPDYQ5mbF1Z5ltnF3Vktt8IpFonLkt3MRDfQeb7L7/X
inJ/RS9pUdMNxKgHySQ85+JVelek5/QlJcMxB5elzav/iSV84IiTDs2mgToqxjpW
FZwKx37HrbU5pu8GmIQ548T2AKTF6txuvI//3Qe40yLa3n12XBUhSOxmrParogwY
4qWVm/UpIAgNajeQ0ULmRVUavmtHsSrnTmY+p5ovC6+9IzMF5zNMZxOOBunKX9Pu
NMxbjzr/VmkvNiQZEG/IaZLQ1Fm9LdE4/xx9O3cjel7dWWJQ7IErizx/PrU/bGVl
Sw99CcrxlHi43gZt8cZnkQ==
`protect END_PROTECTED
