`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jL1Q3kaiOK5QBFY7nbKccgwwWGCPoWUR062UCgFzRLQwJ7h+RVg4/531LVLNsq13
Qg9qec3IX1Q76707KNzjHRDsdruFL/YihLQKc49MdNz30PoEnTecwjqNUiazyHd+
PRRofvs3DPX4E8u+XYu3X0hEuarhG1nnyLNz6Wy9oF89tNbG9+WCxipkUrUSHSN2
bIZZju2Ie64HDhl+nFFTsqXZlwjA6D6pFD2Aq2Xjd8hwcG6SXIMy/ksiDHvf9tg4
+EfO40jzri90vrQxV1afvwVp6KWwMD0ZUq8J1EJZXJZzu1Vyv0XW12Mh3tU2tYDc
Mi4w3IlK11FJXqxy25RWK/au/ZnPqoJphYpwE3ZPeFX4rRAY6W0ZtM4tiOlJjLAj
GTXQcsrH6V5Foibtm1xXVmVszL9NJ7q2Hm1/HMCyUIagsR4UuOtRNk2SUjinL1y7
gHeyGOdtDa50qr73/CFURbhN7O0meY1NRg77KllLTL2oXdgnFxmaaq4dkrisnTyS
obZMorLQqUtY8dOkJdUNIJFdxw+hx1CkoCR28LoeODhui5wL2IbKw/IjFe+kUQmc
Z7W4OmNL9rKcUx1tPBVHtyRWREO3uRZkBfjUVn+GGD6T5U96ABDxhZsyVd4PIVTl
e+ifyLwsVcJNod8p5GCYb5bHXjuKmdf4D5DZLUHfLdJUE7nOOX3zivXjt5aKi2Ax
myyTklLauluE3c7FvY35+aoNd6olBQ/nWZnep5JWRUodE9ACeOMTfFSn5T6u/TvM
4EVSm4njfvdKVnR2gJvTyAb2M5CBX+eWaReRJVAlUORvelzPPQFUpo4OIo8RHKnk
76vMvyB4jkNsbNErjOH6n2CU/MQzewB+Fs9mCYS6W+FJXM4ae42gzM+8zZqQQ6nm
DYnHe5K5c+cFYh5rOAMNUkPLmyo2Z3V4Hy/jNjDCqjpPO8YqVQ9UDSvECNO9xTlm
UGyDicjc6TN6rapuIPDrrJxHBbT9rWZseDVX8BhhgqmXL00vcHMUeMkGEPy8Zsvx
GSK4K9L8KPQM2BloQj+UNTkdvqxCXjJ9HEag0rakgHigIwtluGdm8qZuMG7fgXrQ
XtR2X5rr1HOxWEwlGboy7SaGZL7y9PHMk9zvhm28bB3ZWOoTMu/BoaasMYvJT3PQ
cqy7kcKdvrRHNPyZ79Pr8oPkXe538B2RyNum6Dxo4sCKB+JaQ+t+RnMaLOBPTsrp
rPVinHdOdIDhOMqVTL0pVpsgdXChv3DntHm4eEvLKrZwZkMQH2iGbe/KVFbSKnTD
Giq0YbwnH1p30rBaxxJjS9vyhubpK4eODLwbyyfqBcoxXCfjOixGBRUK2hky7+Dg
aIfMoBlCVfKqCPF5Xsy8IJ6sc+Nf9oDv8Isqojdx6MXFu4KzERnB6wVR/fkI3er+
LIHRzSwOIpRbt8us90niUI59UkfTRr9/KyyQrN0a6XiZCRBCPtpj4NAjM9OoxKr9
6e5vC3t8T//QRr1BMpwQariTcyS02oxjIIvog7cPzPiYURVg5TFIJzNQCnCK50Xa
gf/t53zpySfXp51SF2rHUlGayZmUmCq3HhoXS0BakXgzqK4EAD42qYe8j+S6v2DS
cq+LGSoMl0IZ0IWNAyNDF6B3B5CQyB/TN7RQp+u8C6ac6iHJT3BMI6B7pPUe8r+n
7+yXyYfEBXMzxUoqu5UklPeVzlrZTBg/WsNtmaloZ94OL3sj0OylKpApD6BAK6TH
UlX6k9xDLBTEzOepBCzbtuh1dD8JucnlXlZlK5ALT2RXlt7aTsApI+BwHzJwjw/C
tofLHj8ZadBW9fjJVko8+5GY9WguLudUlxUShyFGKiDUs9r08Ek9LIcRUqMhFvqZ
/N0mPcjGPpBOxgWpZOJBvcgqoqGJaC408xUoZ5YdJFNL4/LilXYLfsCFyIu7+2zC
kw6YYPu7qUy3vYGQDFPBDq8JWA98CDE7l0+gqMP2E7c4Pe5O4vdkTjehv2eIYoAK
RmGN/kpd3PCbN4N+Y9oPD8ybjBavHCmiENc0MKbthSmNE/xpyLr+7hbICmZpDnn7
aL8bLqtvwiVFosglOrt8dw==
`protect END_PROTECTED
