`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dHV1UZwKnXbQerXxTtl015/NW/pgd6wUQEq3XvxmgytXePTBK/0d1m6palmZceZz
KtuP4xJaf39dTssAPaXmRkvCHtuxTeK3LhFU6XwMBXGJQVSz2eKrofxCuJLjTNik
l+0WiPpYczIfDCksXK5TOsO+oKwXONxfedVHRjMAXJQfA4JD/f648KyXddBfG6iQ
MQu9DuE54sAOwPkaSRgn68olf5Epa56JHBOoHn6hY7kpDz3n/ErrebfVx9BQzCHy
8zYLiEWttaVkuXhoqwyM2oaNND9I71XVPz1h2Auyg/VLZLpRkjJ41bz/j2TZR8SN
SS1EkJUbH+nuNi9Om+7vdRMoP0A9UZPlaoYfFWADNP1kRTw7iHE4Z5s9ItR/wgnY
C5xJHGpMVDqJDYrh9axwdNutEJewuNcs6RknM7aFwDA3VII+RAIYTnWZVx+T8yj0
tI1lVWNLcnQ/mOFO7/VYRj55tNYcvAg4Ui5j1gLiJmM8z4KwomNq/vGA5VpUi0uF
IsRnhcaHj835OUNOmjCyOTBMN6AuIMdePhPPSPuBQekn1i6YvqxLcpFIHGRgT6aG
Bq1mZbx5U7y96FnaFAkYbPVqDSzfYxccoAB6uXY3lDnhGUR2gXaRGaowhcyGMAnC
V5uy66bcwhFT5Ccd3sFBxZeZLSv7F2AyWsgun3/qezKzUYRwertlNSXPi+1v0m0v
X9G5FORbUJng28wf9SJ2/MJTWkmggISWvTRXQad28GU=
`protect END_PROTECTED
