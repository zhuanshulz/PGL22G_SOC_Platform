`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kwfAUAbPu2ceK8WivAXY7X6aFPIBA4G3W1mIOM2cRbRiKY2S2smrG887n8jXGPs9
0aLNQMGX/iDdXdI7FRLrwun7yEAx2TR9j96NguDqWIFJwwz3PG8E8Jeazt7LS99u
wV3Qpwar7GIGvkAFOPfNnkOHpyjKeqtwalVBZRxekBp0EClAjkZVef7hqvJSgtC+
LV01/UMcCV7evZNbMTT6ETgB+MDGRSRgvqFXViC6hhdTEgOxKaOfCwPgNhLUq3Hg
925eisnqkRNGfqwcx8OtXOMDGpQYHrcABgppVdFzOvdbXtuCDr02yrFFiBuv8vLb
RNvXE6aWAiVlnQeuscIpOPgoFi5MB41ale3T9VucERo8DpNhR8Anlg1/9uQajum4
k32BoeoxKMja0Gv0tYWu2hndyA+doztptASewm+9N1xICbha8fI3M+K2LI0zK0NR
AvwSEJity6uVcab0tyzVrwP7cZd3tvFxLbPX5DLwF3vmVb0BbaD7jP7V8NUzzcG2
gDfjp0N8dYZLetwpIvQ5mohgYr+4S7tJadBznw2Ti4TIqagOcB2CX3mYcq+YJlAp
Zl4uYy4HqQoYpHfl4SmCEnIRv/astQzLeDFp4UR+99Ug3g4+cR/9X3r+tD9QS9oD
0jKCrp9hnDDiELW/HbWy9g==
`protect END_PROTECTED
