`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wSbTSW4X/++DdPgyOr7WYmuiJHulRfQJu5XRfQ7uQd7tqHpEOmc5jhrlN6srin69
DCCUFJ3pGX3a4V4KMohAEuNVdZIfqjgAuYRENXDDpuenh9biJU5tb7lJS1+Gg4by
PlNfVNcG/sw4KivYYxITAAvxVdNtE41+lYsGwncj4ZrFNM1FTB6NDnzNZDPpEO8l
NaHqoa4fNrVkhuY81gnuF3+iRoT0G5pELb7dLaUH1Mhm3hj74PhS0kSSMyGpnmuZ
hV8JrbN6lrlDEo3ZE5fja3ERajBXFBRZBg8BhbcPnzMbcNuRlxz18MZWtj5dNUNK
EHQkRIw303dY3YYoSlUKEhpoRjCSOacesFTOJphh4ipUY5q0sH6dVVXRcVN4Cjmv
SCwotmyEES1kkw/9W3R1r6NLaeia3FepNcV23hvM1zMdoz/KCtfe4vPVVWUL8Etf
/J6Y7lDIy+P2iZw7ofezZmgvCM9CgB/uzuyx8uygtxrT4jELHrVOJGBc3TF/4Z4z
E+fJsdp0tGy/sFEsmVNfjFT/a+3GT6AwFBIIUlm/LHIu6mLSfw+b6YFTh/0v8o1O
i0zdjXLE+EL2pNk88o/w/woaljDEKdsIb4ESWsaXArS0cHoM6Mk/Gz9uPicTtouR
MFYJSB6bf/KqRfWv5I60rsStjIm6LL9OIoDol9Oy+sgZWspr3mUKJQTI7eYfw314
XRgx9JOs9k4X0P5LI56+XWT4+r4oYXplBB40I/jbdJbuqCdDFmt+VKvSLXbzKRL8
/de7kEGoxwu3MDHjSLjGTyxtD/4AxYfh/WFuuuvHFxH5rivPvlNUZkqhNdSRaX1M
eMbWScm0Q7jWPvpeGEznGb4FE6gZpa7WY7Ei+qskzv8wSVeqKjcjK3b2wJyfXAJr
Nhqzg9yQ29tcnvDrfLvlZ4yz2UhqiQg2E8NpGq26C2IpfugPONqIO3BB8LFBTgKy
JgTsOl8FDEuUTBEbpFQc4vAoaWwlWXFW/nSbESudxJGlLB/N3e4JSaeBlf1eQ5j/
bLcwoDr4DczaLBIGvmr0YnRwnc3pKjwZwsyyL0Hf/fF9HLitqpzATbWxrorgQbz1
uZbOr1StY2hZOfl1IevLq1nohRkmDK2r/HK1SZI6Fp/kGhdwGRzTxr920Xz2/Lzw
+/CPQMOcimdpynee8InTUpnNasatHAirrjm++R1fZl3PGmfkOg6YQVgnzC8wlI5P
cHF2eBX7/xoGuP1l9sQuEOzGPztUgql0AZB4FOugKmEy9cASNpfk40lEDd1JTS5Q
1KuvkVMslDmPlYwPWjpXO7JlslIMDD0G4wxbs2RmRYmyBC9AL1Kbalv5PZkmcro1
YQqSGMyIJH2/wFjD8ujiIpAoaFfbXlF6xLxfRDujEkPn6S2bZMLxLGJyRrMTFJbn
jynDsjDwuuV0GsDuG4Lx1eJMziflztcfmtocxENQKy5rSTz35JTCj8eKeU4ydAEw
K9HKNHOzRjAipStxdfvbHXul1J2JT6kUnJQEECjKADvPNUEciQzqwZ6rEWSVsXv4
ZmJ/jtgQ51CmMPIVXZJyzJVpxZXn6VHkCoOAtqsxpRyPUDvMto7Y+jy/ZRWsAdtu
ibsAWgQbxIt0rA7NRaTitQzmAZqc6mXdyjUrPXtUVR7d2ZnoTE4Y68uNWrPuUn6Q
639lx08pZyDFzk7aWndDu4+03Q1cE2WDXYPhy0PaNa3I4eNJHHlZi2K7zYK19fc3
YZe4663OGpY9j2dDqRQjOlpEFtzK4G/JmxfAZOeUA+q0bwadzTFOX0ZOlAbG3459
ETYAuZFozrvzfheeDBAbG42RrbqhBcsQVqbomhWlhSgEMW+GBCgkJp7uPxX02LIt
LZSSy0oNpSqYZqkANkUBuUot4OyTW5oIfKZE6pBQHmyN926O/iEEY2ve2Qq18W7P
QaTloEKk8F2C1FsNw/q9SGF3hbohJ/P7+XVALAaWhO3Ig9UMEHGzuYhRLjId3ASg
eqEuglq25ymaIhMufXMlBbmleAOHQqhvGyyZSzrCcm92+yfJSircv4HvDEwW58ZM
Dii48uMHs1Cbr04scDmOGjEOfqdMA/yhfYs7zImL3quFGdaCQSRjnmaZgHBfRUxG
zRqIyjUjFuy2nMKZTNb6lczKRmNmhLHUmrRWyQJqOA6VFhy7ga6z2vHhxhGX9hpm
TXOl0F/baB567h02oQ0Dr4I3hwOSEwIOzBByZCmBk1qTxS5FaF/9keAbZP3/AEoP
rLtumZVEnVf4UVFsGKEJwmjxqMY3T8NAZ9zenmujmSZmsi5oPt1+MVkQvOlsVM8V
WsAIOwsPxoiyWsKg5+/V2P898T/r2g1T6G9Rm2Wiuik/i6jj4JQu7t7r1qeGl9r8
xe6H76tvRYL67eXjQ0sw3LQeIXSJvuWSjDu7UP1kVhvmWr07qxl8SRJMPfqremIP
Ol0IZXPVCeH520lv8qNJQ+7sUv2rqAhGTcWLa2mzTJYLX4mlSAEsxhD5t6DNISuO
2vEgqo3KvPBO+U7S5sL1VNnozeEv5OTbQktvSSzbaXb6z+q9vBm6rvw7UV3KWGV0
q33tCO/mvlXB/nW5P00g8aTihybQlfB8exvrmAzCGy4xmHvsRF0M2lMm5UHIzO57
J/j6MaxWmT3gFy93L7B207KGVioHxUaD2k8oTumFUsTX2GRJYyGdr/i82t5SLHgd
JCbzF8nICTDzz3Zapd0/wmkey5a0akHfe2wAZRsxzuzkwIhYiknI7AG3FwiiCpeV
RNNNHgqVu7VnVVBc1XLoEG8YWPmAM353hyEHu/qOfSdSjueB4WOhGxDeXqPiYO2c
e5pOsOd+0wXS79pNOIg5PGelGa8IckOu5niMUQSnPEWqwpoukec2YIdqZYKD4iBk
j7SvuevhDfjBEvYU8HNL8Ev0ip5kAPFO/jDE9AAD92HLLqoShsZkzhTU+evaqFpB
zG6NdQ8iysuQw7MEDIrroDGH/Kg3repz+6mkxTIBRrAENfMWvtP7bcbYzYPMY8jf
qjBABbbNpWOiRSouaSatdigPS4HEfwpFiZkXWvfhRqUzO+KYTT/stW/r33pFFtOx
PXhrZofevzMBOjGjeW2jAEXLm8fMonziub9i9qDKaau4xgzPCGoHwKzwy1PHZNNo
NFvqjNz+3IkqdoKKrhlk97Ri5s6iQE6SjL3tZHlXmDDa7wJA3E2zHrPSuuP1UziQ
rBk8iMqHYUQ5e9F1VoGYyzrc3GSg4Wl0X3CmZZpzauEfLFS7kMJlNy+e/mFxevkH
n5/D9bLi40FKmC8FLlVAAWHoAeYwkeV5kxWOGt+e8unmERcdooMOhnlmOwlH1KQ1
Q2A+ugn2fgPqXvani7BQXg==
`protect END_PROTECTED
