`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JKikBZW59XDvXivCuiTt8NS9sceMYHihakIuFlS6QSmZzebkOCulDW3fhmMtYUaX
61ZbZD2b6UXwnVITF9ypTdVITIopY37aKbgH1BWH+6p/TLNDuOK+xbCsBxagspSa
65mibwab+e9U7eD4c6qmFAHWtiov6vKcJ/plc0FNbDJqCp30uBTItifvjde+gdyL
HOYaxBpb7LA38Db7accdSzjZoUjwYeoOFjctR6zaxtBxvRkn6zHyGjdifguL7860
NKRYxGSNbvNiLFuyejzteYkH8ssxbCR4NsRoTSDNbgDHjqFyYkqJiz5gY0coLEFN
ctGfnF852usuiAKRyZv/jU8W3t6TiZG8QYeg2YAI7s9sY/nV/PQbqJvZ2lEQRcKl
qJiVQpZGvFW22a4Amk85YNOeu4Zz7UqHxkjkHataQDNLAoeBZQFbJJc34gNVljzF
ywZHmvRDRcyr5uniPENrONhFmzbkyWp5wTy2Uf13u6zqw8IoBaUisbTwNSbni+Rc
3tQznJG6jFXtzJknjs5b+F7MXSilJMNw9SmFCSbrjjV2u/y8dRpITOAq2xPm7Wy1
2URj2p++3nOQ/4OM2ZepB7WvCsIYNnDRObZuPGDR5rEPbLXTDbdmrC3gDaAvLU/+
WNJ8otSz+E+wX/Ug+JrcpsGy3gFgjrCKTjM6VFd1AmItjlRUHwlsso4WaHp8Wmz6
uqd74xEvEHHh2IlIz5Km4ZH7Yv7ac6eFrMuLo1zVLGA8DNMGr8CFlK18R6CSlR8t
E5cUzSpESUz50TDEcwqXq98e1OnKWWuHWO7r1ZyTYZUHL2tTnGD+bK/xQomUrVyq
TTR0eFP8G11nmeb5Rje9ArVZi0ectecVQRWkaXHpxUPs9JSxDaHSIOKcQcyuu5SX
rVvQYFbJbhIsrRt4NKyTZozf/jAlUaGJkRttTAgr0e8AxiezmNad2zBgRszpcba9
HtjNqkZboCYlWY4n0TnYQJ5FIUhGDAr5C/9uKIrTXJ8rMn6MiJT7dpCNXJbDjOof
6WOv2ZjatkHUv9jQqP2ISgDXhQgKqXJShUxhLF59ez9Dxi+lxH1Ui7zpaYLpNH3D
GmpG10vh+IQg63QJMvLH9vJl5fIlI55x++64CMOPnbUj+CJb3Mu+5iglnj3HZkqu
J1iS+hInx2fwN8bPY+XZwYdNds4UUdQVFSsBA2Ars7I3BGVodD9Imx3V4gNUr/CB
dDfyo3+2C8jGi1Cv7gBvQSb/NoHoc87MrFx8WpozdxjoKpfGBrVHzRZpzPFe2iX/
k+EYwovlBKv0nSi+zECH9ZgQNAhDGv2SugbmmYWCtXcdzoO0tXbzhVhVOR7uNVwY
JyJ1l4KVqZ8IyWS7oXzW2dtQI9wiI8MT9045d/MMjykl8+oyuqZkTbR+uIoFPbr3
ndKhidv9fOtjbHxBi81dz3hXnV1Rdl4qpU8897QPwv1yOZTguh5gvRQfDiMzQXy5
IUhuFr4Yb9wlz96/sbXWrafvdL7Yt6d+YoHtRzTWBkr0+FIJ4+LGaakbW43l3svq
6eXfBXEtyh2k+PUz8Lew/s+SU3+0NEXdq3oyNSG2G06inG09nFv+5qNcNBmPMIRX
SV6LV0UGcL5dOT7udVSwu91PM490CSTzfCFjcAzx6SEUs7aUUn+Q1w3zdDoIb7D7
bFKlA3Qt0tflkNydYoNEanbbhFKstTU3KrxCUZlm2Jy6CQ1qh7McCNPrg1RdoeMA
k4/QuKlVi/0eniqmFqoWci/jwViheLx/NxP+P5xSWNH2kmzTyOrG+2M41amHBLdz
HwKe3/B/kgirt538hqd+/RFX2LKPlVqz7r0VcO0FbfQv8OZFlryHnAWIyhniu77T
EbkGN5ONuYv4a/kpaxkznpWagjySxSd38Gal0FT19ih79levtt22mZonUvWEfxUC
CQWQ6Rsy9Iq2VzIcUlrNSVXO/Pm9wcLb7W2AtwXpaZuC4vXhIZ2UJzhlXuyzp0eU
XXUpnkmgMnNrManAQZ56SMVJVDo5O58vUGYTggkXDrO5YQ1bHkWRxMuT5QE9MYgV
evn5xasdFvGaVqojlRhcYM7v2lM+oWfC3RiGwO12wwze0gcQzId9OQMY6YPpkR48
oPHeR+iDjGfJUnOvq5dilQ9qaFurwzs6tQQI0lfUSdziizCeamWNUc7PcjsA6U7O
YMnPBPGaia/5LC3k7E5u8hPTWw03JoTEtq/31jofH60gcUEn9h5qTUsudlbojPmR
4grhGvqkRv7JyC6ZYWIjTUGLVXUCfIZiD+KmP4G2JMbETh+1hp+mHJaCU1Y00Dz6
Ae1V6kT69Vwq++wS5YLlqOUWdJya2cdk8D1VRdCE6zZOaQtlvuxMimK0YFW28kyq
MYtUDzev0wfzIz0sg476M5jYJXg8rKiOBcmaBdlbtdBrcm9VjaLdSGP16nLC5cPM
PD9hfuWHEiK3D1KRe8vROKqrhUpnUdT+5kZBNsoYIokilSP2orBfux7QILAxgIMi
Lxn7/KugkxIZ84v08UGB5E+pL17z0TDWuPQ9XpBn12No16VX8iOEWM5tFCuxt3Fn
uGLMpOHhbFpk5aikoHlOtRWAA/adZPdGHGAZB0Yxphvoy6i9200ZKByVV2wVAArT
s4wNWOsYjq0xkIS7rQ7PoximPocQm2JIXT3MBTUTUaXoO8uoAU8PB0MXNsfCSKHD
S+9x/ML4t93rnvlhNUPzHaL/zQ3fIUUKz2AQBpy8E1TceksBizJAjzkfY9ntXLJ0
g5S1Pq9h4jGXnAG6g9TIqq2z6O4H2uymVwvYJ5/2DuR5QbGIDwSBlJ+zMvV1dvkf
gt71smZO6vXeeK1dpr1P3yjmxTqjXxk030Ie9LFOL1y56FbgPb0ec0u/7mJacac8
D3RM9SEXzoL6omsek99jvr+k6zgtCcwBKSPF1QP9A6e1j5Wz5WYh6Wq+Fs/BYhhu
3KdOC2A9jSZdmBuV/61ZsNLEsMr02h+KQV9CSgJ6/sGIuo6Oo85bSCyoH8GlT4R6
l2nIRrVuAlvnN5S6zmFN/CtrdTe07VdMZttYAl+i1E15wOdm0XNExL7XPuOJ3cVp
dT5j0Tt4LDhGkrbwpEbGc93i46jzMOirpbKbDLUTrvv1ZzM0HjOnMQiyxXrf4jzu
2x+Ud8TsqN2DOr0topstHxj7shFs3HGXZFckIcHlT4JQnTrqSLLV6ztbfpvvaZ7o
otcGE0l8Pw9q2VVCtD7LyaszbJ4u+h5mJVCt6ecFuxNn9zkgx9YwbvYYq4xcaajZ
D35mPBXvnJNFS063UGk8lWsjUIfKOvj5F7YdsVde5NEFQoqrKZLb2fmBwHE6buoZ
bFlnXC9h70hqewFTvIw6UHa0WGi/nMFAaFeRUa8LDhwa8T4fAlK/xUL8ak0r9gHy
QY7ma7SGi9frOkqMqa/uhD8eKN5m/lUO+PczmqQsgW8d445hltwjQ8WUo5GEaF8Q
NZ+iQp4E1tcDQbAdAWg98kORm76l8mD4bYCC4FYLOhUBwE5ILUdhnUwZlpcaqdyN
5JKAnGnL6vIBsCSWfYvSDBx5HXycf1O0yqdF1VvdBDQrXQsOEC41fskkbf8579Vr
3h9ioNbbwqADNRc3rwefYCGajYg1ifAad7y7R/1Mv/MHuRoyeDBuA/mZfxjDXzT8
K2TVWc73YvApyBeGZKpdaMvPelOMaJ7rF5olZ4WF4Qak4PwF/vDrc0cwH5VWsabl
U+/qlCqg9+xNj0qniEZVVsxs8IgVK5Gt2PAJB29B1TWQGxTwX+O0keEPC5MW/P2D
CaD5MqYFvtSssIu+3Wgo5sGRKNSwHFfzIpumPiZnUFqc+/VRBF+HnmvZKTwk6UhK
hgKc2uLYlZSkDfctHgGj6djhqIao7kZZoVknEhotM0d5AMHyV7KuaqxzJE+Vzbdq
A+e36E/xIq+o9bz0GFigTej14T5W2fRkyb/JkJGPAk2S35ekPCe1PBiZwjX3iNYh
kWMNIwJ5JiXqV4fFkzMyFBBOBQxAdvvIUkT2zwXvY4luHNWECZKxCjwjHD5zRcvW
MvDCUmabKTXtb+vH7y9HVSGEBdWymbZyS0NVO67X1nL1iof+/qk5Wzu3tSjiAiVj
kkZ9OQDVrvkGpjSJHtmwpf+ToRC2K2cLlJbJuNyTiOok2OB9qAYUTTLPgrX7jBIn
k2U1XAPMJgSHpV9miQGyUKxiEstQMpD4XySScObFJjNjvuGFnemrB7q3OFW5O0Jf
QvZHhFamS0vUfu8KAQb79kUqH2OA3/TijvN8vrkgh89pgbla0p2Tnxk9oluPRXkj
bfAvtv0u73lwtYukfgacYZOFpKSC5EY/rpvOeky+eP1JpZGpr83omt9JPUJeIlap
AFqquDz2zMn8IwvDZolBd0F9GPS9zmkXrQUriBEXDLpuNEUiHDAR/FsJzU3syrY5
pFWek4Ze8M6bmeZtDAzyWG0+QwfvbH7ULqFzhy1kWkeRIaQ9wetK/xJevITpmXaZ
Ui9/kfOF3Bx6w+57t0Y9M7/V4p2AKGv/0jDrNJBqCvr+FihbFWC+18d6StgXeuW8
GawFoxIUTU3T5aedODDAXw1T8tH0gDvAxP7OZk4lhUr/KNwnHEwFpHQ+Vz439gvT
5/3qiWKXp/WIZfP81cDA+QzlPjTecuzQDxtAUs2DxLBFqmrppOJOxnK4DtD30CM+
D9SdXryqj7dKF0CSZoCD9jVMeMUmiF7+Nj8F7vbfSOKCSzThscrKGyaLXZDEJ0cm
thRNmx+MHwcJ1XVUNRcTvfykA4OxABymdxjGFvHAXK0yI15HNI0HCwdsS3ED06Fe
NRXxnXJOR36oxGhoMGZUrt4D08cF01DjhLp1BcXxVgR7w1vH0Fb2yGzqAAV9ExCR
Eayn/oAkETY2vd6SOhBpqMC3lp8VdNcW1RGcdTyZmrzSd0ynH9i3HHPpWIJEjEPm
nSxk48d/1p4vB562aCuq8VUxPMY3tFFJyIJOVCb5hcALRIIx0LkIGb9ZFJsXCl06
+MFxI7I3RiermNGCcQDNzzkohNpA3RiBIy8gb5/rqDzYWMI4T5XNb/0sHUhN37J9
rBA2jJfMrD1MQjIiDBB5qHzuVdTvA1MazhyhyutB1J1xSr2wW7owgXhpGlLdPSGu
ur7C7Rk2ctcJpEYYdS1XIozinw8diN7DWVpPXBUlVrADReVa3ah92N7qUn3wa+Kc
tqay7r1gvUeioVqYtqzGLtJjDHk9p6++jZ3wJ02A4j1BnXzg7eKi2qZ/q9T3s2sS
DAD4AVb9adej/p9+LSZpSYUfxKaWyqd1FwbyQ14Syxb2HTg/LiK2fNYsYvP+/bpz
7VSy7AQJsSHOMb4zSmj6rXdt1dpLe9aIakhZj5xoJ9X+EXplIT+qNgK+dGBhwM2h
KWpXEtFLu/QgpBEnc4K3yhh/QFVi3xi22ktOEWPftZibk/YCO70rFslmMsu4KJk9
G1erm4x1klwQgsbXIjf46kw4JWlihP/pGzELhjH/LZlufJNYW6m+fOvPsMIs6nL3
a1olwucDi4Lx8GLLn2OpcN7xzyA0TEQsZSLXHl1B1znYA4tcha3uEbrcp66cW83s
JmiRNfI5ZYZEutfh9o+YVqzXBPGHx/+TuA10m9Fj83+V/9zkDf3ZlCur99gJqXcn
6YqmDKI6LxDcnaRd4pNYDsFSV/ZX5p2OzRtoQtxWSxVpSimc1WzNP1AukFSf6QpA
hmRPBldoYfofVdhztSrVTqIeOHA3Xo09/p8ho0pbqjMec7rKh1Q0X8Ov6AjbKgG6
GwXzB0xDri6vCVG0gACwN/AzzhKV5pLAg/1XkGomWCPOHo4Fs29eLGWcxX7YVlch
+BL7YKUKmimGrid7g9M7040L3aYMPj/yPU6ShdViA4HrcZ8C2ijU7gUBPehpwRrg
tg1HmJhW8AEr2Jg1HImbEtHaZHpUCwSlGwKLsA0ByYVaSoWt/b1ngjncGOMGxVwG
p2n1TDbBoVc2XprFAJHAtp8xuK5GjTSBPUbVC1SIvx9ovRoMqLjUfUaMLrIxYErr
eXSfUkznGz8WaLq70lHgYpjwFITlttmbIVfKk2nDKMnV7uYn42lJG4KG6yITJBZc
E2dj82JMpOrIjt0wbvXykPjoAMDtiIrF8d8DMyc5ZxbKR67CIwzklDkiJTQL2h/F
cl9GMdXlaPkJzW3C1ZtIbAypm3rSBjiawR1d8XZoRz43cBVzeIiw/SYEsgOZyQfu
DupXfg8Ygwx/iO+KndHui5P370Wup7kLg1+MkQL+yYw40/fg7rIjOY4LqMc4N7Zw
N6BcL3ex5TgKUtjXNglTMqvrISyvFOks0dlIUVe3CRAaYj1jWjBgXFCNTnpKZ3bW
e6vXdsMG93pfxxgRO8z/fOXV+ufDJWjzUOOnvfOJ3ihdFGJkfLYhwR2ESoRxoKZd
azXZhude8Nsmcw2Co9K11QXnymdsadRsVEG0SD1w+galMb2dqEh/5S1O63LCR+Su
fbVnvpEl3A2h9NlgQy8ciVXPqYvpU6+mwHLuXklhEpPzB7TU2wYx5MG7WLvETyRK
+txFoO52/utyUe7tXZWMmKPQT+802geX5qyVDmACsPerFQqc08Mpi1r8wePP4tBA
5PECjFnE18KI4b48VZgFkV3w140K86wT0ZWquDMkRLGjelUb8xi+7uULFLWL9Z69
DbEQ1bGgMDfDTAr09aj2Z+97kJR4VkwY55++r28Z2aoQCHxjSnOb1bMUGUd7HVAX
ljHJJlyOFmdDaLPViEVQt2FWbi2OaJCSPITbdwdXgFjWFL91WSFhnc4yxv1iJXfV
g1L/p8rOoAcnYihkmt5YFRtPWPytddiTFQ9NqDQR3rW1IzTMzcgBF/jLjV3wNlex
L9YelGU/JfpTtkK6kM5ceWjpCMr5u598fqt3FYbSqA5CBWygIK6h8WHxEyJ3f1Y1
UmHTk1ShHaJjcBEhfOn8SwQVV8RoMgIGzrnKZRik9J1bpf6xdYAOZJ0Sxo5Wx1le
VHG34KAow1bFtTu65sElF5T07OT6Pay9opYQbmrdNocIMZ2MmGaP+wXFxtj6Cc8p
yxkKdIuWJzS3SSBkFSeuvxV/sCv4e8Cs3fCaDyVyQI8DD1iHSFyjljLx74SnVB4b
N9hMaXYZtVY5ujrxbD0RdZpupSYVmyj+qRSjlX4FrUYuQIeSRQUzM+HDSeYNU5Oc
dboZN8DgBqciReUzxwER3sDRS1ZUnxddzXDqDu2CeiEDPb3vBnPX8/51GXHSDFZ1
RnKvnx+xqa/0q6oLh7KpzqPw7EO25iRBEBItbf6im4D+Qag6PzB9CGRE3VpA3TAK
y/8QQuRe2Fo23B3w1ZQ0ZXWomSnBAp5wQDp+fT4wRZoDaIjMoYV+8U24t2O9Xvk3
gEKKBcP6bnFFFKjfmY3ZOgwUBRlbIX16VuIoYuu+2hmQO+y47PsxYKlEkylZqtXX
4RLfgoanIWBQ4ICHqVXJf4iw4+zN/l1pyWVpBMAxTV61laHX8MmW9LjpV22Oiqun
1zWqHhYehxlNB5+6+dE54XP5oMjkTg0/g70qXQYIVoMaWcCIF7BVuLNrKFlvMywi
44Yn34u246JdEvEv/MLVEU8Qaq/6bapeiMPDRVg+Do9Hdayb9uLQfzk3LNP4Ou+w
bfBBsdq8YM/cFBggoD/PTA501bZLwJLIH2T3id2Ga5GeGLznUQ0IPMVL5MhrDMje
yy8S3L2ofKIEQLNcuJFM54mrgrEsDlR2nDl7WZNHAOlVvrEpljaNUTcTBU4NEgrS
espdKQGBwRo5jpZ8PboGtYBtwd1jVULIMhYKWkduQrA8Avd4fi01asmUrpr3NWkl
VCwPJCRXGrlfsrSZ6g7Ko0XtKky5k2MUtfBP5ig5S2nGKvOnoCNlpokhFTTuKIW2
VqgWUbdNZQTGkfuVOlQHE5y2T7bw+ht6kU6wTuAXIzB1nIn0LsZr9yVrV2vDzFMl
+sVKwad6Nlh6DBq2dsQxqoBUizfo/ATrAZVrbe+f/dHYtUl/d2Scu6rZnZMgEMLY
m90VCZSGP7d27ikNzAxzBbLipmMAhqQxYZVCQiCj6aiv7RD84oOOtWmdcjOzLdNm
hX9xYnXApfrUimfaFOP8WjnOKEAiQejbl8Rs10lfCczgktnxMPz+vk8q9MqW2j3+
WmTLBa033K3PRD/EeD732ARLqqBTAlfz7/peQ85eOUc7uVfezOqljVDmpbhpJXHl
LgElRO1nRkwt/Jm0cNeZSuWlXAfcfsG4NbXrWp2eSKJu4vQOqdyCQYuJbN3WLS0W
gYF9Py+BSFhLFuSY6kMCQnrj3TP6M/zHyldC5+GyANV1uUkbx7WkEvBYmqKxub1w
PfWQ97oV7Y0DckEw+mg/p/gn2WlNeJxf06VksX4DKtwZCi4gziudM0wN7jMpBQyD
iaUfNGWvq6e77Xh9Kc8sJesJhyE8bCjARfSTU2DwXpv7J3xz3FPB+glzu5xrY2s9
owx0O5R2+T1oyuYL84JEEKjhVhfLgWgWntgMxR38JU3G3TSp0itNK1PmzmB/nECY
oTdq+092OLc1mI4uiU4YxMG7ESdx2wwmnesxxesHyPF4LeDeQ6YfcHYCWKkA6FSU
xYg5E6xhgogkgGyGGktJco40aXJjVypxRisjJ0qvBB5nw1Hp76LVq0bQMaKAC4v6
5XNuLPVefIsikB6Oer802e/5AKcbqc/rPgqJ2QUPiFuHicuKx2gpUMzNA6oKQkd8
vkWY15KdZwqzIRjDJs34Q+yYCCZk+B3r2LWPPr2ZLKq/kTVpSontM0W4SS+lKpKu
J/c253ycIs0xcOm7G1X/smgJrlQ0FCKGQsZBVAlvw+HtMAjOo5oxQ8I4f+Qt35eI
Wf30JtXlf4t9z/rhEoe9EZObFoSkjW7owEoowkBYGjOxlgxi74sF3/5M1MHdwRYP
QMECR7Jb/4OPdGqGqi11xUsqfjoT17rhWVs2eJekjrV3ZZC6EK0kepJk8N0F/RqW
WJSHQ+e0ieiStrjRk8J+OxC8ji6td+wkAkEIlq8npQJxSJEFzSfWtTuWVJG1IZiC
llr0SzQJXu93l5CePy8h1Ni7F2BkO6qdZYPgekQPlzjzV5u8psG4GGEo36Y2dFJI
48LgnjiaiZtsGKKWOvyteRHpXb8Otb06KOLK91IPaoBdoc0YiNgacMvfNSVn/k3Y
pp2utsGTI4aS3JsWm3usb3GUO8rMfcQQb2TnxgFpxRLeRhuR161Tlc5kxpcRao2t
ywRLR0o/dIEg502fxcaXe8+1wnMH3GTbwsk+EpAc8V2GSIsiaA+DdFo1pj30BRdD
Pz+xrMqDZL1cGioCBbCMqv4uw2vvTK0WczOnzHV/fiXWXS3acvDC8M9v6IrKsl8x
GK9ABZkqwtX1IgXBNL07+6iyPkexyBJQtOmjm7FFH4WAj4mYai/rUFdGqbG1irXq
JU5rMe8DDORcMWisQmjsmduSMAqkkpRuEP6UHw0lhcGdVpxoCdg4ISvuYECymUWj
gTjLIvTH/sN3mVI4NGRgbD3O4nXKHjn89PpOl3re2oBgztkHd2tqUF2sN7TncSMr
k5BIf4lLBh1SOaL6iGxjnDtMnlHzmoxGpGyk6BX0i9XrtXIhDt2E7yzPQVvo0vcD
1nh2YuvnQbjGxjwV5cb/vEv4rRN3PXV/UFVZWSO2GsAo9d5W8K2LbOLPdy37MiP6
OCHUaGHGRibCiN02oXEMVGO1RnpREyTpIuJ1bpqyWEXYzvwlaHN7uAj98QCaWwFy
bPjn+trL8IJ80Yoz0QQUbyFbQyP8MIu35iWQ8Fm0Y9WmIskRzVbCJ0dh3wI55/qc
VB4Ciq8JZbX14SnxS6o5XfU3wB1cg82tffj0J1BsrjFebI3OxCJUW03KgGMJQjAB
PMSrRJgo1AciSFbxIf4ZCKrehJCq5KgersqhOn5IE5RmpACZ+Qv1tXDPpyOfxvt7
mQD3/3Rinh+8tmsVAt0tc5yeTri6nIev1mKTtXlPHCok2ra4HmpHHYU2CYk2qXuL
G6Flcn7JUaROMTtoWLdX8w2dfj2BeHSSgKWm3KxElgCTQ3yZCPF5z8JHhCgQGVj1
JsiNag5Y7fcNAfqxteGFaUJrG5lDadFa642UmtBd7ZWCwrai40I+Urh5dFiHkPyk
sGwOm2r+H1jwdHuZ27ex9bJur3POHQ9J4VYfbCG36N8pfft1XRgYQJ9kV9lK7pAf
Ko8X3/bWAOox7YfXZKl28Yke6SGaTc06sRJQ1LTw6NDZchrcNaFxaI9l2TJBO4Jj
uPRjXXzfC2WUqMGxoxQTQJgmWROfJZHlrpIJewP0rvlZMDmrhcGG1SFMZolgmfEK
936u5gBRrLSSXDCHSlGm6MT5+IjpH2fnleayV2znPnHyHTZKIOSsjKffHvslPLUc
jswEU08vtn9KSyUHWKqj8RMMExAi90HOP4DXX/pmHCIOKiGcURAZUgahszm5IUO2
OnCHviYvAW259BWNv5FK2pFTU0SwDUeeEW+JTdZHLQsaylIAZapbL0yiTCQ9PpSL
1PDbwlE0h8yeycMAGkU7IogyGD3n1Iy0nvV1o2+czBmKcmb6T8Pw/gLbKh05I/j2
86IyqH0L/zROfCbyXGh5biWZPkxcMnbSqydeHWnDk9rBBeGoXQvxD0Hi9IrxVkSs
`protect END_PROTECTED
