`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
36saiiqH2snEgIeUZGD/K8F8zh8DmHKkbimA44gNdZ0j7pJ+NIlyxofkmmf7F3Kp
ntcC/bW+OyZ9+HVmo7P9vvi6kFb6sX9YSAyxLb4b/LdhAR8RVFSy+9WBzJMqwmBY
EWe6U1tgh/jgST7m+JhKpntOeUxL6fkGIp/Ys4Sgg3RKHAxGXIWctc+0G9X8qZDB
ADg+Z+R0lW8MZVbn0yF/zZBinpIW1vlbk+x+FSI8M8SDc72Md8HTy/4Vji95v0fv
e3WwvtjAo8AK6O/01TSbHXgyTK6v9e0+ef4+3nlAXq4XyDuQNTQABciVRRec91yq
9ecufrl66Tgcfpmja3aEyRDT7Rmo1U+FdEEMBu4vi/nSvuDyRv9UOmwxNS1ZdwNC
N5gKoZ/VkgvzJjBY4X9w3VWj1SUf3lGn2Y4i0011U5NqduUGE0Pn3uoUDL0P0P26
KaXuqO3SzvpjYcorCCOD55MQoBbNhVswS1g7dhQE/PEtDYVtLSGL5grGSXbsbIt8
+V04Cb9mhpRAnAxJfhwfwz2rFqhSjZtmw01UVOzcfF+CYf2/9+0SI4+tjTgNIJcb
xxntU/vjf8hi2zkZp5CU5jXwnFq4BDVyi3SLDG32wmueu4j+J2J9CK3dh+4cYTN7
ujgpQKmHbj39so3ghiQbwE4UZb4uT+he8nys4VqSbGqaKyj0XPZ+WBbac3KjuzPG
bsHhHaA22ygue083XaWR4A==
`protect END_PROTECTED
