`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bZ6o3ZK1v5hnuEZFASYfWPWIoohYDiLlj1Q2uHIEH08T4EfpVEGsH3MAu8hE+R8k
LJSNIEziFFmlOr7yMXIUbrBxVBljn5Ki7Rm0izzolbhqD+5R04oupLb3E8cDFvtQ
mC7RCBPjLRn4KMflyu0rTVWDBKz+C6Pzsmgn9tH1rAEfkx1iqnRBcIZPTmwWr8j1
fm/VMXUywggb+YoI76BDYjI4bXdcdtLjUN0+7Pt52yM+625dT1k1LEK6xQf+d3Ir
q3lgD588lhBDaZsp1oezzKGrdLn9z63X5NjM0hoh/LbTaOsZ2iNcSm8PczLWhRQ9
7pu5XgDO7Ff3l1o63bf42PhwTH2tGYOsdlf9rZWjJT6hLwJxO9EuMxWTq1zOYRCn
qp42T0pvcGLBAhY5pOtr9qDdqSS2VVoL4sqOc732Kx8j1ojQbTOZEcj43SGm04o5
49PscHpOgc99VwpGX4X63HcKN/81yWmhTJJXvdB1TtZUAdTfDhl7qrOrdh1tSwym
PCYyXnLuk9AZahcfNJgtzQz8tnAFHNk+RjHKQDyesM5yOb9NqOQt0QGgkV8PMlq8
H6uLetUVaiSLAoXEhKcCSV8+B1deco+kckvEui1u5fNw2vrR07fSHz7HHOjTMj4v
uteZ02SV2a3JNddDPBgXSw0ziYnQn6q8Ee0fnSAght8ySgOmOzfZCPkSbe1pqUWy
Q1EepNZl5vol7yBDA7CndoCb4igVheGrf0Fv3kHLkZ/4v1bvU3HjxJvQL6CnFdIM
`protect END_PROTECTED
