`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gpuCJ/mH6wMLclGkN5vbsuKCOTgUIy8fLSj+b0HMMp7dDdt7G2LVsS4UA95q7m8J
3Ya8eLbgsNHqQYuLc7pfR4MLA/6ttgwpdYf5UUKscPgPbVjWY7uGWqoI/sesMtc1
ojr3r8ZUeAKM+hP085n1KnDHtoX/Q/smscofiG6RkQHRTBiQpeqFZ1eEMmNreqcA
KhXkTEdZa5uwYqNDhgFHEGx0bfVOZhmRYFCyXLjb8wKL/Q4JiSWtY+iGCcDi+5pK
uLMJBh1Rv2qhGMopmaSP5tkO8328djXMM1iqWpAZjSoMECBMNumQc4lcxygp4SoE
V45281wAuwaPMFeuWqNDVbDlOvmWvhH0iM6KS1s9mRMASDbWDFjVWfB1P8F+Zl1v
uRrdonaXnDFFal394JF0eEuN/UEvJx4OIsGI0kA9LQmW10j8vHnb+MMLmikjXxxG
p8aK9dIIDuUTpR0RKcPynepuMzEMjaCdgje0AaUKbLhH94C5yNZ/PjDg6clTNoaP
pJqTRICikk/aE6iMrnNnYLt5Qq4UkgB/jH+iIOMWtY9d850FOoDZ/CX4V2EFpPR/
Po41VYlj1bA3KYEpha9exs1bYFMreV2H0+5xzt0XpVNm9H8DvH6JNcLAnIfkB5WR
a5A1c1v6tVHWt/aLubAEeIO2eTSUKz+J23qi3L6CGsYUkMzkXZUUx2/pJZJbUCwY
IhtLQAd5u27zv5xKQyClqEsmJL8YQxxYFHKVXhJagdlt1JEqYSPJYSl35aBphTA1
1HmOVW5gGItfVJUbIt5DwacOlzv3S0aj5zfvmvZb3L6wgh91WLtlDUS0/igpi/2t
8rgSqh5KJy6RhUm58SKMaNUZa3Nnt6r6inKimpli419rz6luc4LVPqtv86k1yFiE
WFtoa3gAPz2oc35xsdahMi50jHeQ22wY3O2gwqig/TdFcTPkrW2j/asodZBEPgyE
ABHfhLpFZcNkpCU2JPt6RtizW7oiG0Q8KNRRd3tjHNAFqE5xj3Q3CSK93393bWZ4
bzdglDVD5eP4o5ArhT6qtL0I9fA8e7QF6xeT1GRXzqojZLFfcy5vS5RW20P6LHNi
2fneJgckozRRo9BIeoUfa45m996Eb1JgN2YJCUvb1uZ7SJlykwfHr4R3eci2AJzY
bQXEAeOXw+NanC1x83MZakQZZcqOOIZe8zu1uu6YM1C9q3wyRe7Tijdi+9aMsGrp
XrEL7gdTIbK6pSORI9syohI5owhsmALZsp/AYiyTlbePwgKIt8tVTBrSEycnzG3b
jYtm7HdRzD/0S5JD7A9WhpT54jVz30eOMzbXkuPxZjfCI+fXgx2N5+41w2WQi6wB
mSvvyCMz/3IGy80cvIxE/o/NLDsXfciiKpLkpTH57xxbZ2z9J/yG7gOLk4G9drns
3Uv7iIcoLVmheMKxBjhBR1LFhfWSv3pCb8Ifnz2n83P2yQidvpLDprSWotFwfgag
IInXArfsLCu3mmO+q7242QvDKnEvioNu9Vhmgxg7mM3ChmndtRxSLFRzrS2Ff2eV
00wRtn+JQdGhQdtrfNep8Tq8y3r+c9BZ7TSEt7MW8BuXkzO9EFHV4qQZKi58SGF2
V/xcNCeUad878KEk/ydfX/K+gbvYRwo/XF0w3krSttchGPRvorEUzBoIry0u0PKZ
33tPBSz4z/6K4mbFECjJsAAV3lIsYdcUGCqn7fG8OUXj7Vi6tT0Vboq5V9DLFBoq
eEg5AEDUW05Y3FvmCGGKTVIQ15btKIBloIZ7p9jvZDjSubw19EqV+Tmf2hjuChWh
r8nZm/GtRmce3uux1ruUhy3s5mnN+V8DDuxiQnrXpIhH+2VAGM7AQbdXyhHfBIuC
96UYB6WMwVFTj8yKdGuFtc5EjyQNzEOH2tV2ROn7UvOK/6KR7XIA2cQCOEEJJM7C
KXPGg+oxAHPOfybrOsnOjDK8pStRGj9YoVWKZryXyFK+P/m6k3HaG6jQKoSvQpo+
jWUEoMKpL7FBd4ck41HgqGVVPw02jtOQHk4+jnDLowx8YxF5sgxCtsnBE2Du+16H
1+rr6nHSPkydrydriJmVRj7E6U5Ym/uvyf9CQSU9WteL/b16m/jwt3ZyZixcjOc2
An/F/qUyA+r/HtvVafm1SMUWettqwCnJQKQqy6wXZnPzrXVrC/Z5DZYhiDQQc04h
B8feyyaZd8+NVrcCy2RiaQiDjKIJ3o8G8O6tFMTh2LfNicTrGf19LzEtJWtz6dLE
JsB5MOHla/crjyF87SNZFcnQ2d6mleXIZ4wSbTP840IT1theQ/Ca3xjA72/LTfZg
HgG1VkzJ58cQoYgfV4lOXbmxWSv7rABerig8QgVMm3M6dxAwHrHin0mQCRlNVmil
o6lGSTKUDl6aErfzfkRKNnM2MXKSP/cvv+/iueS2QcdNfdyO9focoF/6POzYnbUy
DVeES9/C/wZQ6CiiiqQwWjjZrmT/6gABlFWv+d75jRG4Ibkf9+qNpg/lk3U0ilIb
YpOrq1FepnReKAKr/KR60+7PEkF+IQ6SHEOK0VpSQ5MEDwtgNouNHJIlSwbeZXBt
xPMCAECiMWmzTXDDxXBDbc/HoDaHflo5eu5oCaOv7AfhfgymzbQlXGsfH1OIvsfC
rCk/JITk3MwM83JXuUH+D56id3048oq3daVQSAuCfML5t/hCzC3b/20MTT0kSjbn
51DigaloAmjN2dZCeMPHl5Ez3y38z6n4UdClRtAkRf8XDsZQqcGs5KEezqlIB8p+
GvVjrv7sva7vl2GldqolCg==
`protect END_PROTECTED
