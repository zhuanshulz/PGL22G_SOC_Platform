`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BeURqf+gKPebQVZMtSpfQZk1dnw/z+ZWx6iHws4wR69DEkxB8I78Bfd7S8VwV5+o
u9Ij/ZcJletfNJ/J+eOAzof62AWXUGLWpgkdmsTlHVrE/UaEWm+7K7/GV+rAZtPi
WJc1QzUINlAq5uG6yIreUkYD6hbo3G3EYNKZ07kOWPcVtOGRPcvnPRJUyLuu3p97
XSWostf91dB64g3Zu4aEmxqVF8WnAM9A98IifJRIHr7IcfVW8QZnL6h8GK3H7p9Q
65e2PTc+JCQbaqdRBlRBxTbrlUrofJEbGoEfUQ6LLqwnFgEBCOeM7ygV5tjqhKi1
XykmY62dOSJIa/UQTDKKQ2T8Hhubp9+9SPiWONWQEe15J5HC94X5Y2DQ6YrB6ubc
GFa7jfl6J7lbPrJ4JGHkXxV6LOOeFknjFusUpuG6WFwDM/kB0WWGm1tnIkAms4GQ
88VoqTi5EvbPQXPAHvB2jhKAlCoEkJrW8ZfjXzr74TmobYsLG1flQ8wLi4CPZfOc
NFUP2JsJwCsIYHoS22hh/QpAzZ+3KB+4EHEpVjhetIgM0/Iv9JA44qzlbNiJfDHj
70RvTOaOx+e8W1YfDhpzMGAlSm2TG8n5zU96CfzvMAyTzvvvROGDHt4bRgU/W19i
pPKqLPYxwAdTH/vPOjKBswuDpJoJ90PyU5HVFpiPTqR12aT0FKcvh+7pxI10fC+2
XRQ95KbtRJOPdMzYI0EsT2ej/gkOWUg8A9OUxf2PMUdyXxXGfYcgzoAeVzvg833L
+4cNTVWXl6EikyC46m63bffYWKAkX4AJ4taLdyF8zCpEV6BXZQkIOe3eCCbaKtfI
CL0I7uotWJ6dJwxvxG8KxHHUgre7397TIMP1xCp63R5tjyNaLekQGr49n+K9gFbN
MfWwoIPraQR8dIMHglHQLNgBJ9EbABgyNkT1h/5PA9fKICQGWnRomSEKcx6ZPOXw
Nj85JA1uwB5wwB1/JtmNLE7yLA0bHASDHuZvz8HBWeMxF0oBUTMgrDMnts+Rnl4G
+c0nrE9g1SBgCOa91XE8+GTQbeq76aDlB7zZjjhdporqFLqR82goEfqG9HeN5n0z
F9PQ+8t0AqNcwy09ihs7mXYsoUwd56NsvGV9kpb8N2EJ3upl5yjouklCQVUbj/lQ
7/6CSCOYk1Khe8sZRUF3+X+c1pEuaf7ym8V8RZp9lMbEd5bCK7X3NYn3qB/jUObG
aGFfImctfhxOWiO6sb1hfFGUA09f+PvDLm4pIymekfvIbl0UkEV+9tqtCF8X60LP
ovOt55kMQC0Ydv3Dugo/tmA0YPlulmZ4XRgKtDND5L9fh8v2vON2bEeuhuaoHzjN
9eP0/69iDiS04Txt4n7R7PrkJerEZ5gBsALwiaFRM2SzrP9b3ie178WV0a1orlLo
I8/J7B8dWiaPb8/NT+u5ZYISEkgTzncDJcMXIyfU52urOAS5VtevuFOgAZIrmPOa
GBrbAo3fl08f+dQNEY9apnfbzpBVJqcmp5sll6UJd8TYRTT5dIOFDJMsSF2SZ70q
xjNRnhzGpGKpUxajlLfGXhMy/6SUuhv4Nvt3bVGvjQ8oVWgdBm/IG9nvrAVpBnOt
AT9pDJY3CQR+20mtYbXIDRjdU31wmOAQkF1Yjfr9aW5+UGAhSQFHvDHG3EbfhIqG
u3E5p+CmUuccsTxtbMtH/v2GEkBdoDR6IW67cf13vKfQTYq4bfQrzeXfG6hmYpkj
CN3bMVsPMxwzUyPkmuW2wAMDELhkIJzNo0eXn8hZniA4CxWo1EThVhUKCb6fuDzx
Me+Oc+zK1471eIVks3elFt2KkWwyM/KN4knll7tmigPm0UNiJwrxJghkJZrptf77
oDPUfVXhzPZXAKb/XdwE16rEpU4EIqG4nOS8BaGFxirZU5yO4L4n4tV/LQ94eX7q
JVdRDYJJxy64i9UK5YOVpxPaR5MMFZ2djTytUCFNGdoJuc70xOVICPZLViJlDzI1
sa9d6U2wVxtQXUldpvOiA4VuFG9rbVjo66eVUT9A1gF6l4lehG4ZIf13a6IxkHeV
erofnMw0ZReh8Rns+ChyJMWT1cL5CnemfljBsSMo39Q8Q4lSlkzFpM0sxfWc+Gpt
iAMSAKyJZBqmzhE9nbCK3QIXlyIUs5L5vwNVj52Exm+58qidsEqAaqC/hhz/LzJs
YEDtZdCF03zBfSt+ZwkZjxVrCj3whGxzx4ZViuhAPYug255pRpStPmY9DUIjmW5X
lZ8Fql2KjMLDvXVhV2IKpKbo8VivBdsj9j0BIoEJllUxbvVcRvpjXXyj73w62o4W
fAOxRA/g4UbOYSwnYIvY6RCYFxYnskQpy5x5ZNWEOqZ5gj9JQqZCjGlKerKdnfNB
VNyeidHusH2g8SmISzcYd/tTg7bMf8LD1pwQgxRIpBOL1gA3eA9bRPo/KogPOqOf
gooL4VSzOnGmqEaEI20RWxmRRwJClApyOw6IhJeueUlcoZqKQ8Hv2aPwe0Go35Cx
RrqrPuRPoupC5yZfhv5yP5rpPVaYvXqWcmZTB90jcoBrUIYaUni1qhAwSaEOiv+4
5NjCPcxB930zw7kSoFm7iZxqk60IuS8zrfOdbWlXb3KeiVcHMixDV52mFvf/e891
N5BxJaNgzDKKqty0SXUksTbl8o+h6sBy7TpD4Po10+TdkCrnE8fYKUQZAz05KS9F
90I3zBo83XiLwS6WGXM7HhIvVat9B8rmgO1iK7tnWFsGzOjCgsv/TU1+wfVD3uGe
rw3FZdWb4nTYz7M91a8KjyWcOgoiyUxC25WqBETT9wOfDXOKB8D5vvGlEnOFqul+
9xpCqYLtA+YWNE3IBgNhxZ7LDik80ECP5q4oxIOYjrUx751fpToGhWJnXdg4F5X2
9PaWqE0KZAEBsRHYEvHVbzMB+Ggc218W2G01MhEtPBzfv/RZCx23wSnoGmpWT1Ya
eCRpi9/wHlemoAJy0TF/j3bZdra0/FBvpNCfBA61Butvm0/ZqNrxvjP34pLUsu8/
EmyNrxeltGYiUAp0Frzs22pBkMb3GLKEkk8UW9XM5VHvKU1YQ65CxvB5uOM9Bxwu
g87H4VkYXv+V4zeU5UDZGhloKyPNIOi+qHvoN2VLIb4/32qNHzZIozxYt9tmLVyR
p7yXS1/GIcT/7TxTFNAjyXU2T8XK2ULKj5wcqmL0YJbObyjTlzWUSkXwzlKbYEpR
JgIk5MOM1rdHbVxmETGwxZ4vZ5AgQy1c8/oKN1smP69iCHXhodqTvH375uSkro2A
WgKVaNv/DCcgvaWE8DcpVvzDxfWAew1H/LiuhQySrtMlrYBItV+w9zkOEGZmToLa
D5/nOqZF4PUXsfkSGcIRDadBUtNPDGt90Idd90Q6Hqpv5X8lyQQF7zDxUmWyxczA
08EYE70nZ1n9bX4BeqQkRr1TwgYAy0wEqkFynP+P9JKudLnKMVmw79SToXj/8Bk5
zZ9Ky0+Niz3V5fZQjcvFkcri6+KJBadFB94ciPEezG/wBkW/PQbyhMl3zn4AYIgw
evNUgT3WVipcCjlogVr0w3w/JPydEPwXYkwvrsHm1e7Wdy5my7+36Uf3K0bhKnB/
Fn0tp/b9jYWis88iKQ5hQyFKQi40kiPEnBWsp0X4/K32vWUaeAORzd2eLnFQrpMZ
VyxZk9m3wMDWaqZqwaXwFYCo2+zXcrmCX+A0E8PrOt+0igFB+uBh5Ri2Tw/behRX
UPsT1Yjk8COdftQOb1uWUGi9xtbXUcnNoCC3J19iBsvy1iNKwpCq+snJmFDUEppT
qyNipJaAhjpA6ymKug+x6cFOMYFnzRJ4WRnKZ0cdS79NnrZQ5IctMvIb/cEkzKda
`protect END_PROTECTED
