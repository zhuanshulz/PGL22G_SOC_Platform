`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0c5zEoIAkinJINNNvxesEP9w2CbPFZxKK6mWUsxVQ8PfzfQClrJjNcyApMuru2Vq
vJbityckmgtz6p0S50UT+JHUXdD9bmHeOt8SZfA/YMy6LGiolW/O1JoA1C+BxRX5
9avvL+bz4SsCFh+mCTPESdTkUJUjxJINtrikPXZI2+omOg2A8CIRHMYozolR6fpM
5hlbDeJQ9hA2vt4paV0aZgldeKSS398Ntm9PT+hSfvbYUJbmMGtAgsNQRWy0ysqL
ZCxHl2HzOyjFE2ruyqVsjEkbpkuasnERtGFwflUMWbFp2xVF252E86xalBUfendt
KeiPje1YG867FNtZWCclC0GxslgYfgkgsIrfbJ0Aw7X+M4GcR4ZLpsQnERXWN+KJ
Bbh2J47m1UfUTU5/Sojb8WTyLjoYmTRNXY51Gk4DiTQqHW7p4nIQ+yv80GZpmgOg
SVM0tM9b84M3mUOnuB0RzBeSxFrgPAqgBZv4aAv1LwlGiWStSYU5LO6wpwMoj/Yt
Uuk4zecjXtNZBBLWy3L65e1qFJWIiWILX5yYKoi4rEuE6NqkBeCQ+JJ+cTlgCq6Y
OJqsfNRzZIPyzJWXaE+QWJvG3gjnQs9u9BBswWhrkOdoUhNRS0FJhwjP7PaHWJ7y
TxjU71pbFbET8bzDybzLaoKj5TH+wVw2BdqWx/vY7CsIfzOmDjVwgTjOvXam0gkv
Ajzsy815Bidmsa/H+hyfy3LwZ8QdkFD/73uInf6jZs0qII2yREGw4cxrn2nzrVy+
2rxik3iIT437PczqzvHLuxhL+v4KSxc8sFT52OHcXb/i85ZaWbls17HClQ9f351E
gjvttHfsUlupzVmHtqsBxWI6dPD36dKO+hMSlRaoZSWY3HV3++WPDtAUi+SZSQ1+
Q45iquU8jNT2PjMi9KqwpyVaZcmcGJofPkH8CiSjQ+Vo+zBHWcMid26V8p8FuJGT
`protect END_PROTECTED
