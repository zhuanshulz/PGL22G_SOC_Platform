`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HiQ1HuXpLl8Zv9cyOdAYdae3fFQ4OxWP8SlOKX2z8psiQYCJG3TnV9j/+3x+qp8R
dIQF76BoiPF3mapp2hUEOkOm5IrdpmTgEljDXsctYTLONUh+5EpQh9+26NBDUcPj
Z7efczteU2C4uRRJIha1ELdGEQXeEd1O8wv8u8FEWqNdyagIzZU4WXaHyhhZjcmx
dCytZh8jIKmRzotSVvOBFnQ1X8C2ACwq6XkWNpl9eAleyvHf6bMarh+foVxzL6av
YlQzrElKOrjtACf+Cx0MR2qkiubTUl9FDHyzyEVqgtF3cmaDpZl4sAx6rgWwkqYZ
3h+LyY5/yNmMPE3AvL1Tm3HQxBN8Cdl4bRuOeXQUTi4nTYEiyGiZyzt/1bftpLkA
1FImQmWT5okjmd8kWfhvZkLypo9Ny5k/MLbmVgUtKJxZNtuh6NUXlfA8kLHPFEJ6
jC37yn+Ql3ObVZ5SZLOyw9o55+SvzMsP3xepnw2Jd4+EJXf6ktdidmWAlFauw5BP
3FD+/ohbWxa7BQTK7HzaP+9pPBkWQ0/D+MFjE6je+kgVBbt9m56SEAyrsLieLXoJ
P/ltQAjvzZ74KpN7wlyLsjoHofGonnO0lp6yVPSaRPHR6dpulnEuZvSQKXsX1fBt
rQLpOWIUCCknscuUz10WJQ==
`protect END_PROTECTED
