`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x/xeLV3b4NSEDWMEv+TdDWU6fpfZkJ4NB5Yg0otbqS5tlrFT069m/glEAD+XLE8b
A0RFcE92H8kNEWE7atrC6mZJ5uFFtcvn0qvuC3ssATYAN5YamcgdXxdXee+V629E
HCuoe42XH7yxrz+sgw0acuoTZGk9zKxkMZeFhtDenTXSFUN8h1AhW6VEWdxCMz6a
VGtMSDdf1J1FC/Ez6GpMIPx+8aOXC/K/JY7ZfHkMr/opfnlOWzriljQa5XEWu5rO
hGinHUYRXiJTng84NBY75elhRFSgSg+U63Bc7ZLLlK2mC5NFbeAfLMWCQVaOzY/a
ocOGpbmRPd+8YCfRdMfqAvGSJYAicBdtNECsZGc0Are4yU20qbpd8aYTarhATgOD
QDefDeZSGZd0fOGkjHZ87knKY7R8yaS005zTIP4H2cn+NNGh8fyXO5icNLl2Bi0y
k/tc6eUHYrIUEsbICG9eTTMay+r2+jZSRhTJVquV4cnqtIPQ6JuI16KDr536LD4Q
smCAZ5yn3Jakj7Bq0m1ktfSKYRxsBGRteajfe0xxw5iXwJo92hFH6H3osnPUCBhI
4pVF3XYZGADlaVpWH2P5Eg3aRDeHvbqjJM/psbhsdohFr1donnqXCmTVs0M6Gqkw
osaMOsXeLlaIgvjk3/IIqeM6hsE/pTEEzUJRFcBRHi44+LxW4vcay19mtIJpI7LF
y80jZxnaqQy1G9Ks0q1fpyXR+K4SYMhyP3rh7e7bZoVQhE9zaFNi7RM7jk2u2oDM
fNptFl61n5sHqM7syQu5vf5G4KY0nE1s0ra+Y2TRbM0Jhx4/UHV9OIs+zTUpPNtg
UT3dl2TLZ+kyHF+8giGb0pc7WSd8dFzM/Wc/pgnGfETTm5WpWAe2j1CeEhtcc2DE
54I4nSUrBjeX3G1c8avmfnqEG0kMC5Ii7XukDXnyRH2Ag81VJgb/3SV75mLlM2rS
szNCeWYzk3/M6JQs72KS1B/pLGAEyh0Tv+pZ0VKvToNO2x1+Ou59ji+PJXjQzZom
fR4tf7EEeojzRW9hJ6QD6bERY/FkDLi+pEx0tOjcbaTrKbgDBaBYVZe1YbhETKoq
cIRcnQgCMZtJNtCHa+Pjihk/EaczzIOUM7r64u4f0mzHFijzxma+ru715yL0Qat2
E62axc0cq718+lGrfFqqratIDU6dX7IBGpdZlUFWGAI=
`protect END_PROTECTED
