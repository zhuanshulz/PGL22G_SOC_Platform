`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UxPzyTPM8sVJzU6WzoIVGbGzpSSyNUKTFjISIfjtGncA3w/CtHyp9QtuyJ/oBJPp
vufCdjFzNsvsETyBsJ1x4RHgqmEL+ejLkNTQmqxLzEZgjfwraiUD+ayS++NvUwKB
fYkA/8IHiPGgOPeDKZ19+4RMZnTkEqpbIMNp3iJAuhy0Dzf8fKaB5h9rd4JsAAp+
C23J/NSibE1skKOV1Qo9qUupnHfEr6VVJBc7Wt266X7r/7j6JU/tjZ9RY/yIx8Tg
HW3JZQhDpu5zYvmbu/6Q00Jhs9XAruyy/0dThRI8YBMbYqqcCCgnX9wCXDoLhBfl
On3C25dwbmCM1SDinME4w6i3qmKhrYX6DkGfWPssRy4zT+vWxwC3oAQ6Vdr3hp1W
Vav5yZB1j0+7Dub4rqRU+DdQHs9CppIQZ0mXhOnoJlukvjCvASNRmoG9TyGbc5Rh
8wa3zI/F5ZTFZ3XfwJ320mnGDuSydm1BxyXyFaTXfa1NvX7499pfpSkvjhU1x0zi
izIDfRl7+J4Kfaww7woJtbiPgxXmwMlLng/WEOxpwTLGBnyLMaDgzLp9gDjWwxWf
Ta4xCnfGzu2R14zJg8uYY8RXvpV2HbAsRShelr2ROHN0jFuswEpQW8BifPiog735
N2HqMlHP7LPsShecI/OnXuq+4Mb7S3gUqMeWpxpDmzrHDBgo2mdGFsxSxokDBtu9
RMxJMiODxjgSfvBQh3pQ0KwABnXw5DM4eb7/qp8wcU5x0wK05SczlNxJuWAtfBWd
7Z57pIFWZjCKYuySqT926l9inSqog96nJD1b9qp3GlkSPKdwhU42l/FO4CiEWwjU
HD1GfmHxY2LxTnbkf4cX+u5uEfcTbZOgzE1jv58ridnPWy8ddnr6m3whlB+43JOr
9s6jQN58TIx+uMJJIdFaUOi2JSg6+S1r3inrBiYBRhaHZ5OhlVJpMwFYXJWVZSJw
ZBQGEMBJXsaZQGSYhNv9yJnVplie4BysoDIqRi+ot0V2+W4SuLiDfkWnuo34yoNk
0kUgP0XeKjBSfa1hifBISxkn2VrvpAV4Xh9aVfM3/l5hrscTQB5wccEIi9RwAvBB
ZvvUBYhoSYPs5xeeWHMo37w+eL0Y7TgJcTvXZOd86JyH5uCN1138y82rSTrHL/r6
W84P1YVBpBw/+pVEEtbrJ8kLhAhrEBqShVhxw+qEJfchS+PnxmRINMtyKQT4ldNT
fEWE+nhrV0cDcSf4HRtZHxHwPe0NQWY7x6Jneb9jZWgK0/3BQ5Vcguc2Y3zunpXK
jjnENEUHQKF08f22Am7PYOwtJhcVijd4cTDdblJaXajihiqVQYVfGc2U/Aqbf0oY
Ek74fpqthbpJ88oK4eSHQ2W25roDOWXTG78JX/XIpPfch6CxQU/UAOl9QJxeqjJj
tRI9OCAENT9lbtRlBYP9YcbhP0wEHKT94ryv27WWMpnRKE4KOty/0cDZ7BMz4fW0
9JMUY0eskXRS22dsNEqXNDG2RZdcwM7TT44lq3GWmaaFTtEdcaBltgmOEhlbEJYt
XSCS8hrii9JUBFD6b3mJNzlwhx+iBxwejaaCHrSoQsr56X+L2HK93H7wwG0vrmfk
NP05h/xOIadLeVqWdG9YFwyWKmbHH2LUtSId4n+jI7ZmBwOneec+NqK9gXYXPdF3
fz+uUwtjkPhpnCJ9yuwzTCxyGtVIxZIeyG246BhLUXKzvAP82xXrzTrGAWIrH+7T
gzMhmNIt+WFECdY6isFinkMwU28RglWP2vNDL8jSWOTrWE5J5bt4MTo67XEkVgsN
uIIU+Q4PSu21yfHhK0lW3cdeahnzWfJt7lzSw595WobA09gDN+t9rY0KTbd+iuFM
zCba/e34l9XPrtu5GGsK3WCo+E8F7pbj1GgaeKBMUPXZwoIpX/erpAarBBWFbvpc
hvLoWKcMH9kWN2Lj+9VmZpyVO05JeECkfKGsHyaNauI72X+kQB9OiVDZ8+GgMB27
y9k0G46IhBK1aUDQKqgbGlUHRbBqkc0dzNiMZRbe6zbuvn8eKNdQU3PCbtPPU2Rb
EYKTxVOKLlhe3IfinK6R1OEOLRd9f0NWfR6cS7JdYqr8/ysaAxiOKyswymWnK3Ft
rIe071x/ePI/SMOERWWtwyfyzbV+AFUIx3ukhA3LLDESKlgclGx8YFTs/HbkTEOc
1JWDW3ccE7vhMX2F7BK1JozyiXN/01gDYPWkiDqVXad0L0VNsNduQ5SSpHS2KUvO
uVWC22ycoGXcNdj6MR9UPQajLrR4lIMLp9/5Ppw2lhpStbGXcYs8TF2fD7ztNyal
KSAKOOtUDGb7+ilimFt89tsowYro7VUlgvZGbntmd0rDY7FAFt7j7Snz607WuAIH
XZbnTeK51kvqnUgwEiqiU/v/9KwbY0fdrvTY9m4orhmOJLOM1aSmLfgehXM+XUy/
n7EcR97JCn8PmKjeUHDYbJv5cL7BRkFIrCn5DAvh2+1NeW0jieHA3xH8BVDKX0iu
0n07fts+7+/MbJgxZ54o+ijrJy+kMCzxp9b91G76PF+u7AjIMTK/5sHxxlcO1Gi5
hwW5rwh5l9W7lAXMiO8/F93hs/CJBHspybNdH/Fl60UlqyrrfDh5B/uSRrDJhAkl
vCYHgVsm8AudEk9gRNJxyjBvYPpn8o+1eNdz+52I7GVu/HPwr6XKiakhF9s4EU2V
PRzBljbO6IwVv3POE56MEheRgCX/FAPWTvp5HBDgwSgPWOvTHk7/esCHvpPXu6k1
409F5h2IsExAhEx2T8yYgZkHIqpXzItbbiuCWN8iqsjVvQNfC+WeOZ7k/37febRD
WWilzB4x8O9GoHgMebDvPycvFyVRnGo/lE+OlwH/KgSSsk//aIjO/OvrigKSCWlq
ed3Vr7KUwjRBDLxuILVmY4SbcDsXPJWMLUUYzNk5Etz8BV2O9RIBstJBU7Bpwcsm
GEnZuer3EgY5trfj21vQhMhP/iI2roUzZaCfJhg+JjAIGsb0bz17sAnJUc3TVMYq
f3I7rvWppbaqa3kQQhm6EGe0fkYaXycRO9Scm7PJSoiC64siwuTKmie0tOMX85NC
6WsJt1rJlwhed8eqbOcDW6L1gEWs/uzZW5QGmiWDPPpx1Cx2m463eyah104GAeUa
5kyctULZqsy7YEdDzt5AGNfofB/lHk3F669tyK3rkJUWVvHR1uQXsDouAl1nijCJ
IjNn6F/cFGbvkwUEB1zNn0dBjuOcvrPE8QEUP7m6Aj2U3YUZOTVwtKxn0jn2OV2p
PcKTCtcre0TXsab1oOgHpUCEOnqq+Avcs8TVnZzdlpsMT0zAR4QZBpFS1bXuI85Y
QqAz7WCelVhWYDZZqBesN8ItUykaGSsFZCzB9Gox/yY2EiGENK3tjOHfnPB7oXFd
ugb0cMApjPbbkMGUKvdh0G/EhdVTYZdZuXm4wusmoFPmD5p0yMpEwOwtEi4SoVw7
O34l6uUD/3w2ochYTFNTVhH/AbJPVZCnn542wEXL1KvJ8ZNLaW0fof4wdFgvnFGH
G0Gb0UQUxbkND7cp21mPMr1j4PP+qzohT2ZvmA7GYwOQTU+knN8F2hRBu5ySWmUB
yl57qy7b6fXEvH7E5fqTL/86EeSRMDjLagKFUbjEcLBB377VfqywmVUBfiS/Fj/U
8cSSNR50ozc3yfZT80n7qQKSu46mc3hVp9QnRlPm2ghES3Jt3Bn/e1yTD6ZVZmK4
j/+qTpSrd4aUWZL1QinzJbSiyysdFA+YRGcU09ix4XQJ+BePMJRWShif0Vlq3FhN
wy0O7Z+44K2WEZFiQJsv0qeyUl9uhQjr79PZ++AB9bWK8QXx5RRzueSGUlPjfqrQ
74peIu/ShQOJOnOqAYRYpyQT9hky8bQU0kAeMkWt4s1kzdBclsOxE1Inc/D4y3CI
YAJR/Gl/qXp3yJIOK+OUQMc4e0iOXgOXUZZ87O/hc0aP7bU3bqSKxb9phzNbbzNn
5/BD2nj5qu+9L1QeTbeZhsD/+Yho6HRSrsJ3MXf50PQyBdzc8F2zPqU6TONBTkIK
fhUAet2vyOh9gWnn+OsDdEfC3xlk8esgYegTXBD8mb5abJWwczFZsnIBeSwwW926
Pt7RnfrbZCq6hq3tDtwspF3TNmctl6zakSQ3GbvRsXz+4GjJ5b659u5yD/sk9hWV
pV+6X2oE8+iNR/r+dEDXG9n+zjAKsqlSFyYg9SQNT7WcDUlCtA7ezXs56o0okPnK
rNHZ3ncTR4isHn4mSgxSWacUcwTE1VDgMr4Wrj7w6k+DRNr/2UQDFUop91TATMez
mtCfrXdS1oXfiuygwtBQ7LaxAvE04tIp7MSS8uaCr5bCvj+Q7SkVTw/jpX+ix1EI
jNSu2OGvBAz/bcVqJIkrak+KOSUaPQ34jsZrZdYqXAHDH1hErxVruya5EbzwvuNF
61B1LxVZphJtjvzasXAj66SEaNkUZsZ7qaKgZsQcf7jjoiIbnd4m9tuDUZFlJJgz
MxmhJs3xgOuYKqDUPCkozLCINOnxRR+MtJlGSKH+CYZgiAY3Wg3Pl2zpEF2ymApC
22qVD/dV/5Rr/iPpLg3HHsZYAzvQoZL5w/OLlqUdBD1JTh3TXgED31LP9P+7gW67
p6GmPHZJzuSeXxpU0vxrij1g3ymkPfcDfVd8aL5qDDx+CnL8x/ML+oeQzo9ZIDEu
mk6r4tn75XFrQlzd1FBYjTo/7Fv7pYzg5CiJ5R7MrP2CFqCQ37VFs67zFEdPYriJ
ENSw4uAoJOcwZXjsnEv8ddW8NE8NmVJBopUteiKFCDgAv3LFvNStF7tJH+3150jG
yZ7tHX0LLEHqgsT0T1A/k3guqfi6sFeb3WGcjzIdKQoQc/LZKeoxzBKDSJnt/BQb
LkC2CAPcjXkp3Pxk0jxmLfhN6TF6qk4bWZu/rFy6LZw93WfNgT0V1SOhBKxTKmUi
15XheOlewjrXjxg7cyaVWI8ZQO5ByHGX1i5zWGBYTCFu4pyq4nMdi1iNDgvifYqy
5diWypFFbH+ra61vgFKOYP5S+EOK4Z0exTESaV+RrAqTEF9Lqa3t2200FwKfYwy5
StHI5afjVTm8WxdU25eXGm12q9mNAdTR2ZRHLpC3PIgyvq/nXVa4BNNoRVtHNeiQ
akcWqmwO4whIb+UwJrFO8Mmw0Xd8QXL9ltZ22Dns5MrueI95i8QbvB+AoNbeg8q7
v+tRI57fgwFpMqTI56/9RrYoUVIguN+cs4lHScH7cp/T8LJXZ0HoybEXVq/2fpqU
Slw2EP+zYZ4cNemsREJgXzYaFMTPgpZHLtk1RG7yPcdJiz4XimAkkpX//G+Lavwi
ZxPEH6uxnpkBGckazGdmFjGRsDy53sElOiX20mEsfG1W7umURXv9ALmi3IOI/RFG
M/w/SvS9x2bDOgq/p2T3Jj25+pXqd3o9RtHiF6augh13d11t0IV6MhJCUk2zxSx4
UKCcfjwKshPf+/66SqYchprFL5PWhBy5OXjKvrdZZZxTSvxLyEtwvHRD6SU6W5Nr
Dow5i73VZ6IFAhleZvpGPtlWgmZG6+1MKdOd6LFCqtfqZdpkcSCHNctoHcVn8SBF
S+WsqjTYW1wKU1eiC4YD2/5CsWL64H18Fgw4jFIQxO3jzO7ekbdT5G9gNzTSPNRr
MesBeVqvQ5JR6vOoyoc6W80fD+rh791UnQzKO1FZdoS7U2cGSy7qEjfMekMYF71w
PvXhjSueESh5CL/n//+TynrwKCn6OJNFTYMEIeQ331ZEpdjRv5xlMKjNB2jzCt36
RUZIhh/IVdNNt4XlmZ772SaKPyWn8lHPL7BUOtO6z+cDyyWC4DX3xuOSqCg1xn0a
naiQ0nRoxIGEUU9OqxNmR6vLGfcQ4TDtJSKLhmdRxVhg8EApmOrxLYBb+tmpthXf
wfctrvfHujTHIDyJhmJhyfbZradkZiTI2+PuTffJX1L4XHajbkeerWDm6K85uwnC
JeylxEw0J+JUXoXSAupXGeamkH7fknlNj+nTnEDC0J8H2hd2mQT6ul1BVGG6seU7
uHfWiStGl8KVh6SbcUFdaR58hGralrEbGGo60elBtHLgQP5iBIb88FOvLWhwndag
1uGOfGzLG7y4dePQ5VglyPR/tdyKFY2ECTdfAC211kEFjg26rp2Uoafx6xwsj9N5
hml8DEdprOG1R4y7+24NmiNVs/PmkjNSY7scpcNWR4ttEhHyNa/DAVk8YmoiequE
9tWuDi0KiIFzuyEO5w1femxe8PkOk2ZVXHALT1mvFVR/R3olKn3iYClEqtjNBr2G
cBK2e4tXdolkYvcIN3FkFto1CHGqruQjD4mQO9PtxIbrKekX0O7FwEhF95j8LYYL
itRsduTMq5mb2V4oDNS4ZC4zS5oOLwoukscOYpRKxWPyMHcFK61N3vDfIDVg5tgQ
T9fHYWWA+R5EuQiXO1KGubl3Bj+vg4ctaLl0J+kCl0+2GlRVQ6hxlk7QKvuX5w8/
E1qjEC/gDnd5M7LKTeA7VQynygXucnxmjtnFqHwk8FA0haDQOqvcuW2nopV+EE3T
XtFjWaubA1+74XOlMs/2dr5XiV7BZARgbrbWUO54zuP3g84rj+EM3Hd2TJPQP2sQ
e3WwDK7x+WQjwrFLCyrZlKPqFihEFZln14pQOVvr7j5sFaMOE/xfuqP+LqfIJ1fz
Z2AnVPZkYu7aRhF3s17DveP5lAIlqobNrkQp+jT9xYT9cX7+74vRKenRdcQOQJFB
3MZgXg88rzm/joaaBJMR1qV/Xg+KEpesksnRBYq89cRbDUayEQ6WVzrW3EsIAwVd
fxPud/zQdd8ZjgpBU/709VarD1kiDOyVQom7NwdcPujEkh/l2ulTC94+DbXkUiOR
nrYhmW4HbtercqDIBW6p++jjbiEn/zbJ1hJqc7wo4L5K1b8vk+Km7GEcSaaqvh4R
R5Osiuu2v+Ou3Q7ZPcoIzXix6r1tdiVpBAeGh9OOEVkR0pEC7TueU3h/994aAPA6
s6hvdFWjBCs2yDuBSjGsXPrJvzQnXvW2GZtQNGNvSmNjAenIj0E/J22bW2ElrLT9
AWEhLt42bh2oEdg4wFU9CFygr/UUyNeQgZVS1Oyw5VxotDXE7ZcYM38q3GlC7TMo
6MDh35YIzhbiOpWCGQxkXjnvmHMjKAi6JIbYaukD9YdwxueKhf4RcKNqYH57zDfu
Xx5DdlHB0n4aBzE5xWeyNoSVaaBqXdOkBAIhDdv/VCknAKK35gEj8flBaYySGnoC
I4N+4Ds8deHBRbCrDgI93Tu2jB4pJbAlm8V4jJiUgiLLpqRyv2Irr/wXJWiXmTuN
9rzpz7LJJfr0c/CQpoPSBKi/JKqkfQ5DA/aB73RNom+pjbtyol93tYJ4IFFBXGOM
8JbEQ1EljEUrT2kpGE1KCLLU0Ut9iGgJRRcZYVGpgIDFkSqLNgA5z2Cbmxxb0uwW
s5lbikfXl/ug+yulw7Nw5X/0ZVQTGLb28yYSE4pLS2p5M2/HSShhZir4UySEGBAF
9XK5qA2KP/TsMvjNqthauv3OpHEPziFQToMHURYNiYCh5xpdaGp2azPmCsfc8/GX
M0LFvnr3q1lIrY8Oe0xfiwGFZGRV5k4uKbeW8d5XQRPvjGCy3E+QTi/8y6x6IzeS
oYsErgtSQhJdLlNrjaB6YYV+pLVQNfhykGq7GWsvKRGl+coYYyqAK8r2My2rH4Z2
V3xrIJIXWJmuwy1T97LQ+hq9xVc9+4B0q7KkDZz613IjfdYKAakgEPnR+3ORP9Wy
PEiv3PNbHxBxVcLzU0u26F9xxIh+nZAiCS3J2ie7ChfsboSdwqfX6DTpVdQKTbar
gT7HP+GmwhWkIcmel01gK7DVszXxuECg6oC95EzuHBRlQiWaw+Be2nkxPNbwgvNB
VpM2L008QbnGrHGbOFnUCNZHf0jc5mzf6sfoaxrDawMYYhSvjOo9txdOQ0gs7Upk
17sbrVAvnYavQZ5/SpW70zUwrUGGAwEUBJag/Z5rOrBFjvaOR5ttEDKFAc5mUJgD
LyZOsAaiILgAKWOHtTzuZRKuaJeRgtMiww/0X4akotu/K024wgfr/rrnx7sjzOkd
y1ieb3wB6nLjPnq3KjTAie6s5KI0ZWSD4VUlm+rgeGYs4ZOGNWegUAPQv8RvssKW
dZUCD+NZLB/P8AIzNvIzdC4r3fUqfqcEi8Q72XazUsSVMyPbCSLTkvTGTf91ffXn
v2Vt5klpHCixIbI/smeQHQpBmlPFAajsn2QSljAR/6FzUp3bAqdEPDBigSt3yWqL
f4Jy0qsx2aVqHQkgQ1zbEcI+8LQ/0+Obb296p2KnIn2Tp+2+6WI55Ki2FHEwsq9t
d31AhQbEqRGQXPLPlWKTWK2WTZ0d5hv6AvIDP/xADYeCWkKFcRQ9Fugrlz7dJHTi
/c/XEjZydirxs3A8dStLkj/iQc8bAZ33THFqOzzx3X33FTZQlEKBUd9UdV9KHbW3
pLW66Yjul4Yz5D5OjjAOZYHpXKpn2HOYMiaxQzugLCzd5mT/zXlBp8o1u1M/Rr3u
2QaW0ftH14XWwlPeVPevfXliKfhXHKOgE9nX78wpv+zDWYhji4Z85vjdeIS3lZXT
TNx3xpttUyKSIQB/RpHkXbzD8DNB3MLowtPdl+kQSG68Os5SoIwVjdhLS9IY8a8B
KfyhR4tejwayF/rgPH56BD6qYpiuwcM/4PXOxYNeiJkZQCMvlYmySCS6uKj705uL
7u/2RrgJ79TywDnjStG02tVTOPkQ+gotyaWP7+MIy8D7vybL+XVo8TJvdeXmU1Ht
661uuuImTxe9CpuOiditEHcrgbMtC/zjuDE7yHr4/+1DPd/LdZiYlBgOwjUsa+wH
Yeu6VvV12kYuCDFWAyRlDaVlyZZRehqn4pic4mIzg0DjofecgopJT6cuSmnCgHY6
AoX7sLVyjmGNNL6iO5eRlzevLYvGYqfxoZI7ULmDEa3m/JHiuoll+E3cXLrNa/My
YoGyRs35EuZkx6ob/Jj5uON/rmyDDa3hmYzCPDaqsLJeIuzCzpzOkn3V8GFWBews
1I8JGQ+piXxA6pZQ7L0qKZyyOU4te7yeVGMHUd+pHH+lzOaY2dahpF7RafO1ox/Q
9/AR06uinPIycNLsWVrCh0n5Ekr6Js4u4/HBSpuasErtjdXl/HISEvTqM30A9zm9
hbQzlS1ylCYTatBytVXsKDpfgVFVVvGfi6pqkMqSwpXYKXN4mr8KwwYliqyc4eDS
xbSUS3Bcqydl7NIrqF36lA9G+oPZI51E2VjvuQHzZHgZUVh0Z7++7jMDh91S2m4I
BAaZkEnPs9Nq9QAve9ka0Or5OJPPchY3WMvQ0RebmRomVZR/1oCpWjOM8Razl8Qc
LMSsQQcmgrpr+jTb513n7FzHsWNOorU6IEGYjeCUniyd3aPidwzRWqrOlv11R90A
aNKlVuNp4b/YhvqtWC66UDDboApnVVDw/E9bpaNXOtZH9wkepzUU+N3vnr0JCH51
fHfzONcT9cdichfRGztFOVQJALl8Sou5z+d8nPAOLQRTOtAQ4aOdGzN64mvhmVgI
PCO7tje/e3WECBa2MIcuLX776/Hr70Rae4S7KSs2t1vils36LmBl0n1m+arfnvGD
RCjlwx83r2X7n9+WfNwI1CsHn8Ngrl+BvksphJ80yTCYs1MOCWVxORQacm8Lz88Z
AcZFYQ5VvzC3CDwZ+QR7c9m1SD53mDkYQrkIxs8Wr/hgLtTJQspNAhhjVy/xvpDe
1hW9FjfkZbMNkxgjJQ+51CbXcB7foldbgHbLW2+Wh2fUADDjzUbhQu0ZSHSYRAxB
gF+5sfZW/yBezRllvwb2ILDWeMNxl8eoadYZ7bNCdbe3VN3+UiqYq1It17UvGqAu
ejp5QVTEDxI8XCCJY5zUbF4WgQ2CSqS1kHe6eX3cfQ1Tha6QYSEbCqaZJvPBZ2mu
SV65glomHgFHvy/9uKry3A1WzxIPV+6FAaAH7uQU4uKiAIWR5rDc5gmOWaNznOim
1HFiQxvIVpi/H76EmZ5sXA==
`protect END_PROTECTED
