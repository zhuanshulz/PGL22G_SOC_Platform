`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JF1vgx1RngZ/3WNygIn+GfSwLhAWJXbDPVvNcF4agV9aPavrsuDhZFIy8fg560nQ
cLkKeF4jzPIS+LPLJnIPC+hmkDBYVS6p+BpnUNqLmgs6S4ltYMBGl21QP1aFPMJX
HErsW8RIaeASXsFRxzhybm66ItbOageOo7lN3Y3oktKD+cDOeHC6NqaQpcNIMoJQ
W+3fn/d4dwta9xOP1tubHiZvLbLAv2fj3b+F7Jsf4Em/o7uYwFJ27eZpByNAUYJf
FjmqXBgOcYRlFhTncHYIyjMexENKNwReGG8Ztwkx7mUWKZDaitQlHUGwXdAYwdQS
MKNve2yjMwgB0u6O5pfzyWETk09Y7BZ2n2OtENpP3OmBJ20uw6Q9xA3/942CREhP
sNLbrkPxStHB9LvtHYLEHSHhllEX2b1kmjj09YGO3c+t96UmO6B94Au6B56SBTbX
8Rn14iOP7KH7JYTkXuLuGg/fefCgZh2VmtErvg78ekbwLmhEAPeJl+qMkJu6AX7V
eKZC4y1dkcSf++s6Ejzvuyf8ebJskMHJ/hvPUa2CElBhke00E3hFj9tuiE9BPhHC
v0i1ZQoEh2DovhB6R/2zKIsJrM4ks0My4cU8FAhFLoX5iC3pdpgb9E85PtU9SACG
ZuBbBkhDEQ8Mi+FXISM9bOJhnVbLsNtsmxMTlVtWa8O/1Eiy3ESaqBY0iTVuHLG4
GEw/m5AqevAXFXUovDMg0SfK1J9U8cdK+ZNvOZ8wKy34OSYfihiG6ZRoM4KzX45R
oRwHnQZ45U/IFih7TjslK5PkQfMutGSpO3YJzKUQA5Zn/xTJ3yDs/jd4lyriGpQK
/QdJtquTJjnHUVy1H91ZzEHoxVMiuGuBQ/P7uKPVIZbF+beXaaz58XnfBWF49Ecf
yJg3es1wKKyP+Are3TMzk0EigGtzG9NqNSFVUa3nH/41bLs+BmAqLehvYAAUhmq2
ZbJqovvAQcXC1sLwdCw7O+wOpOVX/VvukQNGz6fVdTIKC22RNzJ2psVJDtStmyH/
XFH0vKethqqV3SOy34kDXrdlRFFbiHwBqCmEBgKNwZbvJ9v3AmoZTFpRw5TXkQ1d
zLYojkJkbwOnXG4gQKs3NDlsftq3MBcV/mmN6fVnsykFdif/NeXrcOlLv9vZnW81
HYIOjjct9rJct+j3ewMTRRz7zP0+c93W0A8UxE6nfgwGzW/PZiZQT0ydsnbb4HJy
jcoDr2dSeo6/9LhJrODH1yEJAUP3x84zlj1zBouxO81dX15U4/CIk5qmtcIsUn+d
kRcVj4fvgGH8y1+CNLLJNcI+oiSiKikJOvTLFByVa/uppV7uKbHlE+31gg2mobQ2
qhHmZc3oLPoVDfdu2a3SlOIHCdQklOl/Ut0hqmyHBqGg4wxlKnB9nhgEVNcbMdoQ
/TnuI4eILtViS8uUXYm+Hh1CnJa9OxDVTbQH1XKjnrogLfAB3mXPJXRFikBSVELP
TbTFby2No3/2sD2vV1VGzw2xPoPEZCYhfX7Ib145G+ekAzOs41wUU+0XnYdzGy6r
88Sy3MRuZsrw3CrZQ4NEFAglrAhCXnkDHeRuzOmJfimI7hnLm5qvSmyIPdngmg3m
MOE/5AwDIN3HDb5T+RgP9iqYpwyegy5sVdLh03yT3CeCVwI4AjSC0rgu9AO++zcq
IM1y1E+QRA74I+A+3qlHm/uYCSqI+Q+oYSNQ78UfiU6EUJZfno0qvnqdbbFtk8Up
i3r6YVkgW2f13s9tX+bL3br4XkudUSGCBJpAuUZh5VYsW+9TXwtdFtrVG+Khsq4V
78/MJjUo9D35fB6he7xFL0zltUjY0YzzdTJCRNLHYRPEdMzYFq6J14b9Jg6frJcw
VvchVenADpvXj8rZVfXaNgfvjQdncVDTP2KOTyWbHXZgcqzXtSZoQGvwsLzjKN3D
/ES8JQgwS49rOfDJ0WQ6yqoBVexhpgnuNd+RH3/5Wxq2yKHUP+jMLPBEE28WrCPW
7u4cO+Etmm7gBy0xUVAh7O7/nHLDjokjoxtQmv+q6ja2mijzPEdEVaGFnlydcNwj
/zVDWMQZtNHpyX4+svr79RrIGlJpFF9GZxiJeByXxqZ2FTVg4+GeCRima9QIBmHa
qgWCt6R5wfixCXa9IRPb8ZUvuTITHAutjsQVhZYL+MHETLPC0e86jmAaAFUgk/+u
ywafBQEpd/FTTfJKD4aOLIQ80sMr29NmGS8dXzgdl/Z1/m7fvIF8jptpEqfKlYUA
JXryBhtHGFbNViNr8+dv0ng+Hzlm8/7QHM9LPQJnT1Nz0iCRhxNJYf/r4C55dwQ3
kBBQH0IEVID83M338GBLRE2576BV6Nbo0W9usMDsYx+J7kWJh4Dk14HOml5mvErC
aB8ZtkW+/y9eSRRQaS4IyvAplzO65Ud318Y94TsppK2ptLOL8tMsVV/+k5e0KYkR
JDx5ZK3xgYY3h6Nw3lMup2dwnkuDYOD4QRavGDv4O8P2TSH7YBr/bCW5nsuGAOcz
OA+ekxDCu6zeKizEoXDz6P4YM4B4Iru99C4L8iRRXTrBIBDHuhuc/5UXKXbzFgge
VabMBUeFqLfGZ7wO91kYI3I2G3kZ996DQ1wRNKlXzzRd9d8g+lphGUJOB0tSDZ1t
ZrulklVOyebYGWsHekb1kXteIWkGxCZEH9065+lSWX4=
`protect END_PROTECTED
