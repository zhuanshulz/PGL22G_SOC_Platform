`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wBl8sx+gYAoV70hwNpymNExDTXJLmhZBSP2vmomO4NPK770JcVnzbuLWqJLpLQ7O
NKekz9nWPMFTPJtB7rtoRgi0biT8fyHTkdjJu03oHrMP6vUiLvuWUPiX1c5aJKoA
bNXtsNPT9a8I4tVxJBESGXx073yUAAbNOeGks8IgLij87GfyVLRXqzO92OlQVl5X
oqEKAEAE5c1OKxWT1Jl1DZOY8F9CHWGo++Y+ieYeut0t4NE3tkoLUYsCFZBHs3Qr
Zas32Ga8tQicadi9JO6mKLhlXAhDVo2jIN20hRh+9DFArgJQnCEXv5tjj/BZYIo1
DTxYzuBjlPHNBLjIYFwS82I4pkjaWC4h3OflMhi8QNCSiyXBM6Xx3HGtpg1wOjAh
rOZnSO2cJpNc9cPAUu0kW52tt+dVUCQHic9lY9yGyIpPD83vh8kblpzoJjdHz1ub
bD8YfX5gikCrzBe010Wmem0wpDXgRCq2OOeDTNQ+PnNnG84b1RlYIkk0rty7ZzXX
lCjZwBAzV/Q2B6v08lcOp8HwOnI6wgVEUuu7OxXjFH//LLQS0Cv1UN5lDBdwu82c
DHBi84Lzv1vynlxs3jHMlclziB0j1l2en3hovO0erym7n/rZS993UiBgfDwGP8PU
6nZRkpbBkfELtf5ZIQMadtLbA2T+dsTVdLUxJpQ19tXABat7JOSlgL6TCaYXv0XS
a48XUZcwJ8GtchGYBr/P4LYfoNhaxy/04fYfqqECjj/j+lPQQ5iDOmhE7EPMteTX
mG+A4I5L58ldny86No7RHyOpaavR8WCZVK8qKvnDgmah/13fvGA+waVmcVbTQ27p
cAn8mpgGs6LWtC0Z2ya9UcqfeZfoXYOWdI6R0An0RG9fYn8xuHT0+EmGLXzRCzA9
lUyERRjT5ODAXDhxEXu2Drl9kUAlVWBw5OdB3TB0IhMLw7cHHio3D9P71dwzzkdq
E9Ut6dfnuLtGHHvch7MHMwnvkwRRLu+TXo3YfYnLNNSe+/gZqkg6wsNFvmEwfSEb
pnlnw8y54GZ/Htno+hv7o7PJxOyXLQFeKDxh9fMJEFh17CiFmpteYeMpLRkoiVnU
vCJWQ+4QH+ErgF8lpkReNq7/RqLsABff42fAasMN+3leJLYGycBA7xVK3qQr5mmc
Hy3zH1vTGAK03zRFxSgbH0CB0tXBJ+Qw0xsXhMq2Ela3vwt40GFiyy5dssYKFfa9
eF+PbEwzMSsiXVbqysQzmYu1WMmM/yzQnvjy5K3ali9TZuYYetawh8hF+IUpGMUb
67jtBGzOakkvtSgJufOwzyUMjTFFJ50tmyvbvRIjRt8f6C1T9qAqC3hXUVQuH3Ip
0bYEgDodRws5ecfze1PwaBPVNUTlOu/sU+uiEQVFv6VuEY87tc3hdDwQ0LoYVcOM
UzKSms2BeU6vDaN8OK+d6y4vCbo70ZbEQjpAmTdDoTI+IN6xFFcxzwdg52w+Y2gn
elsKJTM+u+Sw/TOvxwMvJbMqZQh100dH/eLlDmdjdXB4Ts2RlsuY17XfQcTlyW8h
pchSRsNj13Rfct0kOz48tm2xnJWDemC/j8R1S9H+IUBNHjcZS/PkFJ8K/aFBpRv5
LZOmzxo4uPGFv4toqH6akER4eBRFfaCzWLqeKxYyK23/5/YwWbRCF/IW2IY0qVB3
BK5DmExah81poN9oSupIisJJjgcLLndZFeymPtkp8F5ai3QPCpKh5WypMtJGo/n+
Eb/8PRP3a2Bu7pImWzbL+OvaLvdRTitqvCpvqQBk+SoSC8nFbDfhz9nsl8FYefMF
T6bv0Pzw51CJ+5Jy9x1rzpFNq/4Wo+eU/DXcFBox8/C/YqONplkN8iAiympBS7Fw
GNu5PBvSWIXWwZ79CEb1h20MVDSiasF0CtUqX49wn/jpxA/m2KIFYNd/gzz0S7af
e/Dj3cCtX7HFmLxGby3AlZgbbKE8KAezp8Z+wj3yq979RF28BMDS92E+zv/OKqk2
ChEOz1qne6QWU0V6iyPphA==
`protect END_PROTECTED
