`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hRkxvz+XFR9L/uZ6SpIXHP0nHaYIyli7PY7XdN8UGLIsCZ16mebYDGQ0m2GaqcN0
m5bixykGWdTvva3Bv0dNWBfFgZGgdPsg59fdmfArOle0tieLmd7jr6otrKgzTLmg
aHtCp2i0QFJZ5NnaFWzE1uzR/KCMA2DbhTnYCckoAE5EX4hYsXQigizy4GbhVztd
BU73AhAs+k70ZH3BSja90uJi5X1mm/z2AcAFQHY+Vtc7Lz9RBMf8zQy5ULHfoZvD
zgQNhaRQ8cJS9AJTlEWEqw30orargIvVCSLrDTgf9KlDxzguifme+zJvxt/BKJCt
q4VfbICWeLuK5MK2pRCIfFafjiEEGmntshlMJZLOwrFCPaOStJ6L6Umho3ZUE6QM
zDzL3Ea1K5a0HZRLGa7mEw==
`protect END_PROTECTED
