`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X2PKAKb3M7Z8XasmS2xyBHHWFJHoHHvIwtmfWw596FOhB5qJP2tPFBkchf2vOmYm
gZJ5b389BIrGGnUmG/YFoPBlMxu6okB12BaAFOojKjgXpUUi7SiyzLHxJ1cvkeZ3
qVvwo2O4gZdbczMLJZW6Z0Ha+03IWRll6W+ISo3g/cFhXYhbgjEGqKa8e6rncbgM
H4APUfqDqHYk/ZrRMMbqOwA6BEdcvZejPTAx+oSMzBy39uSVA5fa8G3SitdHkf9o
FtcF5G6XHSewVqPw+tweqB1aSpkgSisU7Zq2ylUQVpfXApqWAOO9bOtQJCIs1oPX
m+M9FsOsJjopiG366NZQd1BlgJDVVoiKGPMOXBbcvMUKLEQSbwWtSRoEgkgwL3hR
H+UmnOQtJGnVoJqBiphvQ08xOHVMkGLaXX8Z9G9+EP7LZl0H52Zchn8walGa1pnC
/MvmBJjECoKhRH/EzctLZ6nLIzK+y9Vdd96kghhxL7eAIll0m6gzbyGqbC5Vkfhl
P/tbelBr4jnPI4T44NuJBK4VsKCitq2vul4awCz4zfVt7ZuUSTL41obce9QhFvnU
lGMludAj+nXRHo01pZ+cYHR5ArVGyZHdFeJ0vc8YIvie6km1ZgRv86y4v1GkqdGk
Y7VV8C+HfljdSqBhPBzBdHrp8i8ngfdNGVo3ry6VniUW7haoKsB0obZOz3cJqadP
ejgh/wvUsC3QfLTYpObLafs/W4x+s0ovt+TfjMzMveGCZazPeuLgN0UrRRbPXGTZ
wvZRioSPMgiK4JzYDPPD2wsvSo3vsHXBoZ9lZYxuoRBpEsfCzk5SNaEbSR/jWlmJ
/d/1ru9GfFngUjANdDzI3y0qQaHgzvD4NlfVtlFnVBxmVM+TOJd8UQK6Fvn3O1OZ
VZjZsv2uVa/BbfW6WoTGTwhBC8APmhFOn3TPbG6c6kpMlhBZqQC0J1JtPGtfAXyj
gBbzpN3lP2fuza15tXuM2HswITIKI++YjkQkHFxOI3lIKK3AVHy+lSdh9shoy0Zw
uEMbEeKVVhovwMceR/57LKRJf/nJkadXaldlSGoh8ZFREzjxvUluqrusDMxmNarz
IU0Ivf0EXkjDVkAEatDLO/tLgv7udL3deihRL0rbLLnIxx/yUTtZjaLvhm05N2U9
6Iy14r1wjljzccCh3oYVFPI5mhlidNUPcJmoQWJaAasOlklOcHF4PluRMUII6H6+
Mhyvil9seXyQQE8gIdMCXhQFyoUwAEN3LnFAW9SOftJk2YUV3SbJuBO7kk++L0Qd
axXHFH18KY/W2ZtOIou0n9ZnmJe7cslRZxnGI3CczxD6PMSrlCMGEAjrLIxU2i2S
OfAWd+h35ruE/tEarkTI/7chV2+ABbPq0tW7e7uxASWzIuzHVjzsWja6gPcKjDzR
AyO1AVYLBfcPRpMzMBSFWLNl3SSkCcaVEodHBg//31nJr6tPY/jwlhP7yjmC+j7y
AoQ2wU0YinRfQHbRMwwGzQ83XFSYrSAZjcn5B2tWVHo4+43AoaVsKqHmHwT7Y563
Azed125LnQyAd6dWDvHtjn9dIAX+dIn4t/Kw8lbnh+sg1YuKNzftHS2yeOCDHGzS
ZRCZsxUStYpLY0CZP635rLEMABs8/+CBsHGvzCOWwCSVLJFWidDWa52qOoH4RVFf
48NTWBZ6oHmcBiTgPzFw9GbIWMz8HEHaurwZiN0G8pbqm/cSfzkoL1lPrq4DLUaO
xi9FmrBEhC1g9ZG3eYpoJYG3tRQPnX0iUp0hB8k6VrKbu3WrAd+D7UvpDxY3/le8
7p+k2LW9O8FMqfBjns5fhW0p24hWr5aIZAWJ63QYwKfUGH7i2NjOl/UYmPkEYyQd
nnL8bf2EkLxixnYB3VVcy6gA0LGsVm746chBubcl7SXKMBVHynrvyzYbZ4jlj0p0
wc20yqFnDhbdRfajMI5wfDICyoSnJeH9VKmcwNeoKLs8g0VN5S4H2YxNBxTx2bqK
m09fhJWnIPI7+yjZXy+12g==
`protect END_PROTECTED
