`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bv86jdqOtSl6Ur85g1sIcGlfJz7riE3dccOK637prWRmEIJ2twXaWG4aezg/S9Qf
ZQLQa+H3yx589MUfLgLNZNKZBs/8KlpTBu0Rs8j7SdMqs4/V2bbuU9iMiygdJBix
gkyDqhLXpeyHzaZdEUypkj2ZVbX1kfPoK5XAP6SoSRU1YiHC4x+xlB2IF2mql1xY
Xid/ERPXbxCjm+OGhr3oRvir3Wg2D2AcpOPBWEHnJTuBNVglzb7HVzWSQiAYK3o3
mPO0aDKyNjj2/1Y9skqSHOFFNo8XwbIhzAs4pKgMr1t5HNYj7jUjPmdZFIqsn7V/
l+J3GEWwNLhH9TN+5GlsAW5u0PCtF7U6T+uXyI/Fo/5mCHvsdv65D8uvQtiPBwwk
iLwVOteFvhTTddnHDw89v26lltZmQwOikCRHjhRCGivd+IAb3H+dwNTFnZzzAdtE
UeQC6ekfla0FVHrYmRjMkIyTmyKnHdcGYJ8U4oQGZ25x1S3FFfaCCHUINAdIZq+4
6hnBuVrMXrxp2lCS79NDqdQd/W7opO8W+Hre7Fpmc8YRxzguxhXZeDoN7x9VKYFg
HYHjWcKWwQAixTPYMOEIJ88WnAHyu0OScfFo8/Y+SdGhmiPIz6sanQlRClj7iwqB
8HH0j81DFcWkVcxkPETKq3igFlDpntzsXrcS8KENwTEr5bpZQeqWKvt2CCacmVew
o9Q7fxS4ScvqKPLRGroQodsGZAm7MqlANzlAzSrxzZOO27sgpLMe+BXhdb9aC4Q6
kQGYsu4FsyxCefbriClu+/Xpx4jOrRFHEKWgs6etniZ9fUt334QvWMsHY+y0mT6+
jwLuClrCMoVcxLQzBGvStoWtyk3hQ1iFqc5gwxgLQQEJ1qaMzKLNbczHJYi9pmFD
YS+KhDhS7+u4LnsUT0DyMA+VjO80M4gnfyI6ltjdDft7VYu7DTaO99CVbUqCaROc
UuGg7xadf8ofVHTDqU9PTzRS4zZATahRPSTAgp+WvYmMbfVpGT8uvve7zf64716Z
zf/2sv/EF/4nJVnF9W7yC66gNXwe+6QbO9ytzCca66nNnV43JdyMWbvmPzs/YRYf
ZCf4m3OYgOD0HALQbBGVy8Nil3LRQRsD+yziFEqFRe17pdqseUBCOT05CgiY9MlR
k9SlWcoptbUPSJunUZm1ct9uI3XaXelobq6cesYijenNeNFPVCbMfGFaGETVyBSA
A2S7NgELsMkxv4miX/FWlV5jz0OmQhzisCVVlIVnm5DrXUnxsEOykcFM0cNOD1qI
KmvcjHTv8zorjsFoXidJKUd/e4FZBfYqZzeajfI97P1BSVmSjgYF/qFXTp240epK
6q8bui0Ub2BKUynQ+H3JKkDOkVjRuhjEt7mlUli1nGhe3sDccqw9+atL0lhhkZjY
YUSTbOdafuSjRet6YTUCDt1L3JDb1EYzexPfwqdzyRbPEiMubxRmkS2Pk1Oew9+1
bjG+pLHO3MhYFY0aYETqqkFJDEbKfL9BV5pUt1hKwk0p+L55Pkzv08MBsU+6KwQk
offMsMZMpPjDTcopaMRUuUUtQgQFr7FBrvKNYdteh2zZOhQu4taFZQHW5tOWmOBw
MAqwFwFCIfztuDBC8l3nGcuOjRAeLnikuX1sxLuupDZzjU3keveVV8US7moQH51F
7AxWEyWKfs14F1ijUtTVaTiv/WK+rEoSd4dwBnkHZZearaiKNtrfEVZN83CpYFQG
z9FW4FWQja6vdvaQntL5aChkHeAGPr7+0QmrYIc0GlGL1CWyAbTFHg+D8NZyayVN
T+JHkyjl8HF0+84oZVSMEnkK+mDlAs9jDLFSMU99NRubES7xEOCKapXeo2t0N8pv
llK9qzvxjhBKhJkLNUECGghnLmTuo+trcQQeiE+JrfG0Hz6+YpNd1fUZLuK1VYnu
zJA77KYAkUrWBsFIRju5Krz33bu9G14zQEkTGg0MrNMLeUZsu8RdR4tYhMeW+56b
URQvcNblrrnPIBA69MnIKuidG7i/gzP8jgjqX1YJG3Ih3WYobkSaWFNP/IUane1T
hKis9+jz8M9pIckHlQj+1bVrM3F5Feunxa9/xqEVvxQtEQ5SePE1MOR3aJWd9Fk1
t9WChntkQd0QP6JGsMe2M30HoCUG8UjTacFLSAORr+v39BNuqsVssel4IoNjuKa4
AYbKARFv4GmLVHFW317wR6Ycv3T2LFL+Q1LO5zYxRkYLsqxCU3+HQWg/jD8xTSS/
tCo6jaPWKIysgaQ3LZmTC0qgexaY+/aY9EXO0UJs2v6Qmf0A6NZKFGQsPzXFvM64
lLdarLzpcaZ7LrUh+Hnj2gY5f8u+5DLLNFSaDLml/c1dpMKxoZd1PHb0o5kO6oW7
q2FeMFaSp+x54Y7WluA3KhG8wwGtAuXZU6c5NjVwsGSZM2W15z9Hyv4JyG4G0EwG
KsGvVR5vltWReJC6NmhEHl47TFcQmIWZqHnQvRKYkoSR3TE3/TDC/DRxvETG/HIn
DKuabu2G2NuvLO9AH8fX9IxxxznBTVnypiVV5Us/V2HPxDLE/b5xU2Oguj6d781d
/wsq1TL5Bf0/FBniYTIkiNqRRFgZ7+VwCfcVJtnTDQIO2Sf1Hv5BxSlR7Qm9bE09
oFK1o7nhDqQBosQhzyCBynJTZhwVNeLz0EXnFDtAJiLjvcD31HPO8O+RX4jB0fui
ZSUqcwtdcsA+1334B2wNhqTDQUv/Phcp6+MRDqopWtFDttLqGSLGBdhofHS54kjv
JJA/Y24HhR6hlVPM400Pb8d6+R+VvQ1AnXP3mZ3OqeQ/uSty3EW8ctexMiZNjIWt
iS2mZiUu4e+L+pd+DG8w/VnjVl2WI2rvukdQlgw2U8MJPYo88xCscdEZF53p4vKC
sbK3ZKkWqus4pXwkUMRtdIVO/Ov4PHVv6NbSo8znXFs1Tix7z2BWLu9rcSy0UpID
NBiCFZksXACbFTF4CNJWmnhQa8UhrlgXTy9Kfvsil+Gr50Df4tg3Ud+bU2QtObRk
hOr3o6BOq1STt6Fhxb+ki9kjsYckPp38n6SST6fZGrwYXUlPqov8yi48cvzJGgLX
G/cLsftSIi+kOmjS8w6mqq70fT/Qm2fwF+E1gmCJaINmQ/ruS/ZChmgp8na5pNUD
pS7gR0jsqahrwI1qRMF7V2ueTthxYIwGo2LPWZjZhXz3Oh0CDCTwswiT2N/1uPeo
UdZtNdQEi0VLwKfWcsdaZB9qWCEy+vWoxVCMviR99rb+KHsgKjg84SPTsQE5cVTD
iX1U6XFlRtExsTiIz1DbrUsFGiFoQdgnmRrXxn/liShintr0ix2YUtY6ZzXJE46b
So7OBBo1n/iRoGToaClSN3+QY3rpOm79lwwadFOmJOW0bMdv3LJ5DbIYu7DetU0l
duVYFX8/bHVMjhBqF48HaeApP8SHp7JW/IQ/d5ny8hUxz0qim19HKiv1THGZaC2H
zafP3b2SXNthqdHZNvKT3yCbLfPPnvtIbiyv4QA+kQCnvGqJRIwus1TYt1ZaXR/D
WNkQ6Io0E3k4Tl6AzCWwL+BroND4Rc1xlBQVEScNsvNOYxgYJT56LGkZllkIB8TQ
s/9UWjY3A8B7AeUWAXsM/403rjEl2vYBMQJ3co6l7pAYZwzODYWGWKYVNV+FWJkN
OhVfmmBy7qg53aRWOcQZFG6+iy2USGlyfVYhifFReTvmhm6lBtmqbJQGUI4YzTi5
adsP6cLyjnRZXCH4g1vthPGmMrkNR+5lwN2KnqCwFr/QZ36CZcP6lOb5MOaEiO0h
FODHGpl2quS9ueRhtebzOIsqpR5F6ptHYPNZMW0Gz0jd/dgn4OtlEMPUsIBVb5wY
4zUC0wEtfhGmaNAU8THdkM5vrYWynYBnN6EkMFVBG8beroqKsrS4imNxH+iTDMV4
ILjie2mTedw/pjF6344uoxAQYXI4crmptvVv7aa3ASdbtEyTOmODl7/mfF8YYFCA
MqRW0YinapNlBfx56EI6mWuEgMRxY1LC/T+DqmITEbNHSTaUSF5eKz3YJADx2xpI
So2oxnzX6onAF10ZNCoMxy6ASoE6KXSZEwRhR3AndM/HgDy9Og06/nEhScjiOfzT
0a3PgnrcmAd9uDQd0XR+CjomUSCWX+YZ0RqOV6NrQJzwlnEqsOiWv0ynhbu3yuLK
Mx1R004pDvpddVTegy84QJNuF4wV+08gJSb0vErRYmHbXX7rEyDv/yWVtTzfoXYG
oZc6I3m7TKPn6FNn5BZXps6Q3DXKPkihu/kUSgStNaGFfZFGycfphbpMB3YLj0dX
wmR7QPxkDxxpM9SUYjWSk7J6MCRFhJMXIGySJQQ/K38JlD5PSFDhl5+gMevailxI
fDhF/HA8C7uD9O0OoieU3HMeZJBA7Ji8gRqokbBsEs+4iEsRuOjEoJbMkdkDqSDP
VD6i49pfjNM2SBldTEewAkuMQ0K6z786MfUB4tnNyJPZe96WqAG97ILPMCDIp/WL
TxjjB0uhQog4TddkCzhuJBsjE8UbuSSDixP5bK/ie+77AYwUfDlEnVXClMWbm2y6
Mn16UTSlBHNg7exnn79bGAsOsMBBVEAgd8ShAJNZYdRLsKze2iUV9FCF+enfHSqV
+fOWlis3b8HMO9JumjiUhKMFmARcGUFstUkc2Lx7XyxATEYIVQS2D8SiJ1/636j1
Rq+CQEfue1f+9KHZ0P8/zPYe+G906ovdCVueVBv8iIgmdOXmm6kx8vmVSEzIcJXg
I06DYziHfcDmFG8pqAmviyjqKnBJlLV2icVHQudhBSQjqJ6va090eMbOrv70w1X0
oX7SZfvTiC+PmNeix0rm4S8NbinTSb9xzEPCj+N86cuTKP4i8O/QGhA7SJc13LJf
ujcqwh8O2/lEwS1AtQkbs2qd019Xq17jTP2We8DGH66MrmblJ0gS9h3UDsnSJ6Mr
wc0mnYNBpMhWwHSyVCJU2B6roQChfzW2KZdCoon6NhJHK1ZlBajZpi4FuKTrPwNj
wVHTalJ2uZKlPWh0VGZ56J7jtFPalOjLAKaM1VIfqWzEee4N7s4KyxzHwu9m7oJv
ybiRRLKXc0ScQz1DnD03ufoTv7Ha4jD+o9cgdUjHLUNosSjO4wWjf7SB6hY7b/1u
Sz9SclKO4ae88ZrC75c4eSCXe3vsRNsn4y1wSQ93DuCDt0UzRwQfBOOgY2ENoG5F
O5Vb30aOAm7urDffTe5gYRa0FycX07W8S2Kslmn9y90ZAuxEn4s0u+IH+5v6yX9g
1Su4QFt+7czrnSPWjHpwV+mE1ravKVkBj7gaGPWNWdfrRRAyxxX+EuD9yb0YmyZk
Zc7c3UsWRCbitqxc/mfPNCaSfDpBKfJDOYBX+s4C+lghTD7IuROOlMoioDoeKq25
yaNh6jrZINj4j5LMME4EPmiI3RQ8K75wORdJrVrTI/nKdAr4LdoFJg5SSXOBXM/j
hbw9t2byD+roUyJatH76yMraEP9kPEw4jJekvW75lkZ0uVUkFzqkKyWV5CMFR+8h
tuJv8BbS4DItErEr8VM7TMv5e2BZ5rugVcoLbMKL0FjMpcsJF4IsEJv+IZWx5RMH
JP/iwFYicgXeOsNRBUjbZQRzBXAAtcT0G/rYkDFOCBhoheV+ExfM/ebcvZdZdUeD
EA30Wc0bK2qGNYYFcgx+23wLO/aaU1kK4+p8jmpJADGRSR9ZcTIDYaTSEgH5fLxC
g4xCQfnX5VBuGDPY+hjDEgc2hu2NvBSzm+uGBaNUPhpmXtanIdcoyAFPJi+wMaiU
L7NlyAcaWpxptMQxyFSsrUcXG+E5UkUixwee/Vu3JlqhZFDrsWrrPr8+8jpn560i
af8GKANxHiHj6nx/UWXLQygCb4AZ5l1PnrIz5zZFgq9GcU2/NOjZB/EnT05UNCPu
YSvyc8GP/HylV4mJOTiMwPP6y4vvp56de4xZ7+P45yt5652sNGBJnx4xUwVMVduL
MXMoljTXa6+ib8C5/ElQ6l60EXDSJeadSA0XjK1dfwffkt6P4nGkoVEuTHdBQ2EW
GQypAxHjOAeYeMsIa6CRDlOh7lEwYL0fBQhHK8J+CKxIjDQ5JOK+Om0QB8hVJ34v
n57tSGkOdD01Y+J60vj+pgNxvky1wQPCyv+Q4uNvnP+WdGj4JXIt5lbQ26b1qyef
vV1Ozwq/2j02xWFmRqNP0Re1x0thvjOpF+JrGoYEehA6dDeVhH9maIHOcLMlx08G
uf9GDl1lOm9GEOHlBzAUBoVmvbCmcLzpwfsgPoZbLSy3YeQhkDb7dvvvms1g3Ya9
EXmcLtvN/3nw4MNlZXdKlCkiXM4+N/Dxpcs+SrGBHustMYrRe6aO7ZFb1MviIso9
7PwJ6A/chPKYQ2C6RGkB3fe4qOdAy8G9tDfUjGH4bASdNgFtPFVuBWcaTnGXhzII
gQWvPL1qemIQ0LswdtKPexB8SRVmjq2+ysMxK2CbCKcO2Cwff68rscbSemcziQ/d
wL1SjEnNreFtKa21HzXat3XFc9s2HQ/icIio83HNRpizbZvdX6CxyaN4QKwShcSK
RVWa12Ra3/+9Mk8EWCcDqGGlDkJDXFZpspz+/+N4zGieqwqU8f7QxDRLBivJsVyH
hEwq7uNakhC/G9xizKr8ysDW7rCmvX/gY9cVp6Ao4pef5v7FKQMBuGCtv0h/Ym/w
UUyAOQWNqchOnMWj2Lk7Zj3IofY6yC+KmCkndEGUGk5svkEXtJT7EZ1yfuxd6SAM
tls53XDFvUM+iR3c8QF9C9hc0+q55zXfq222YCt+KVBrFknif8KtrwicVLVTtIYZ
kkyG/+QG7/ZPPqeztnLKbBSAOFldl5qgMkcz25vAsyKf8YKivSa0bHbX4jD6mIq+
RUqj4z4KXRI3/pjQcDhVe6t2kvRdWnG+eyD7hKVeaa9j3gJ1lZlDZ5iMGKDAF8sc
TxOxygODp3NVq/X4ENqHOY99Ymcx4aABEepuAqKugRFI1rZQB9u38L+I+lMP2h7O
wQOU4SjTspKClkj2e8hCSuEzPZ//jpom9QK8w44wMV0b8omQWSZvk1ys5hgAWYlh
b961UEou2dp8mRC5IH2wzNDL0lVBfcOIfTfBfsRC6BADNbquxsFVGrdkQtaca6sr
gRxXjBKrI76ZQqq/PPbdeEyMMBpWxgKkWQ8SGf81i6M9/TRus7vEwHWMebnWglKJ
`protect END_PROTECTED
