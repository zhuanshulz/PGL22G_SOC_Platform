`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LEwDQ8IaYuQdDc9ZQa2CbkkaQAtXiwbLkPOF1tFrBtZ5iLVkLLCq+sV2lcQiWGCI
e+uYnpe/uqaQSOHMrRJzW15B9Y+XIxCRkqaKOtxKyQyfLr3pBjgvL+TuUvH7nvKF
tFNczl8JooldW2HhR/5RY/Gd+QGTjTycYAOQMOoap5rwkjW0Pl3USMO2zRUHIv23
7H0xmVWspmrC5sXOFp75MdeOGP7TNx/lrQGJ42i1xNICUrjmgC40jzrTYqNmn/ge
9wzZfv8ZCb2Y3PU/vTchNm4su5mC0jHYTJPHaSF4oxuAnHiqpNd56meO16ilbdu0
EWoKFDZja5IQ51+skxUmrVCoRsoG2llEe+LUPxRPRdFG/cv+1UBD9x9wVBAl1Qm2
ACPsFT4AToJLzHW0Aj4MGhuzNdkM/jIBungH+hIe2YMulFHL9p0N32dNWOjvqya2
mzvwnybp+q1KdjeSmlx+sHIzFoq3AEWRkznXkVWn2gsCIk5BPa3+Wua1moQ4pMLM
jXme5uyWlDbKnVnzB1t6NypMpblRuBUI1pX/2yZMRUHOc8t71+k7evoUG88jWnJ5
+eZFQl+JIMg8puomIUtxD5mkcYWdTPv930qZkXCJ8QcZIQQNaJzCxvyYf7GnuOHn
HkibqpubVMc2qTTtx5ETOg3mnkKyesbMdldICQbp7rh1U4n51WHpsq28p1iZ/2oF
0DJPTGUhtTsKZURJ1aShn1lfgITob3oxRoBsk1drHMnZFqseLH/4GtRZxl73cZPt
afz/xx6q4sjpfphrW2PIjg4CH+QKkaCoefOWcjwhg/ouZkB7hZm+DOFWCwIQ91NZ
yOEkuJIoxVGNyrWXLIfTdUITV+JlpxwrC2a93QmfFk72jFkydy6Qb1ButgQc+AKX
9FGUZFdJjb6NF9q7nf5RPXhjqIaD2aWlH3yTZdUVr9mIxWeRTj0zSAjQg/+hDRKJ
wvjX9Tkm7ZXh7aH16qFUUpCQDJtlendYj/EKWupueFlgypmUyomo4+aS8KtRncQB
dKi4jNu7HJyRzYHRGzEaZK1RI0wkuHfr7Llbn07VbFMoMBxxai28Qw5AamhR+R4W
qtCWwSF2rBsJdEuNvdxxqhv9mhKiHUnN6VdUTc4nPc02ikhIj+EN2lZQEUx8DT67
85xOgSFo+9TmQAkg1KU3SwRHA8BFcxp4D2pofyzqsBCQGKUZ+ZJdGnVe0JOlgrun
9rrekOZYIvGbx1lNhr8cQJgts15Sh4v5DOtYaBBCNxrzolUnGEKnpX3QNNqqMGRr
89qjvFADKbJ0DmRhDDOKOrLFOPuehBT3KUDmwHvvbL7cNlpvw7pTYYne1kKGuo4H
zbiZd+2O+0OJktVF3267QkwGssGV7HIgXZIr4/v0Qa6Cm5FBuGIl+b5Z9kqAfafE
ekjK1zPRsLuxSEZevoVt4O6HDoyBE9ehN7jf3vnNjoQ7Wb+ViO0MIxQYruG0gV2B
Q+E5DGtVv2oQpRxeCx7gHxOu27OKehcXRthVaWHvGbZfLOfv9BK3J94L4Uy7jXzl
HP0Zxd5F1JInNrVCbVRUqD4fJ0KNoIShbBXtV1fGiOAOY2esEDDF3M26JiX9j6hU
F6PKlWKT+bd1TfHk20TXJy7O0fIspxadFTRVtOn8SN6935JmXDyYm/CgsAPNMT/K
IlImzMBcI9KFcUtpCFCgVinPrlCPOgRGoN5DBAEYp/Xpp4QxyG9hNk5NITqldG3a
85C2uXBBYvCCgsr16c6yPoNJx50Iw5QXZz84kRW3FkbMN8/isubH3XPca6p1WWO9
STPQpiTwW9k/OkZx+JmlpoxN4aE6mZ+sqCthpAlIURsgwmAxW/fn66ImTbOlGrhN
FWLOHEm8zzErMeHZQPOc5YAjVQFygfVBAR90+RNougYlol/YDkygPATjNg72phLf
RtPMUPeiInFY5gZtRUXi97Zlkz568yqtaJhiRzFo1cXRbipwsF3angzISqK4P/q+
TcSlSTWV6zykJWDINKbmzYTSDyXluEAe4b2NA36ehRdiIF79f20/2zXtue+3xHN6
sWTKOORJzJb8PltZc4r3slZd0BqYg1TTFdPtOT/2rIe84V02o7So5pDCvNmTvyVW
lKNJ2OOrF0Z9ujmdOaZv1MVnGeGZ2A1XdvECgpDrRmkmDApKiwt2i+pQwEJQo8og
fXSnlgqewxjUTsFSBvP20VJKtyCSfs855kMGi6SeULPHfhmSWLkSSARAUDdp092f
GjZrHvzzoK1qGIIaTGEnZeudepf4cLx++ylvqliNg1yO+k23RsI5W1n1QjyCHpyG
/Ha6umtrhRuq+sqzCuSI9BNfz/YkGwIt7QnZyRkc1t/QX69qbkk83XjPciJcsCuR
Xe2WXs/LJobJNUhFwZan6ObaexP4Tz7d+P4YF65ja8O01mrgnxdriumfKOxizbNo
5Ak9KOZjNzeeVxOLjiGssbBdxpvnH03DKRVsKeZNTticbrrWvvoMs1YFNj+Zf9IO
w0KP0mnWLqpvkpFjZev1cKAJjmhLjsYsDOQ/63BNEtbUGXEMqqcrW7cW7uiF87hA
nKIbrkUv6kYFSOq9+gvhEW4GdM+sS9ywahraBnyj6ID2PIzRFlNcVr/jg9oDGJPI
0hulMNIq7KtGtAi0P6vLqgyyZqPelfiXJVShsUac4a6yOZrcwhCgjcFxRgQfKrCb
VFataTDta4ycvsg+VtBJiT84pQycIiMT+YW014g7z5E7bx65zzWfofQYObEyjcga
ghV1Jh8XvRSHZIljlBC4RgAcuQ4XsPwc4gMZq/aXikD/ua9uJRCdGvH9g5ti49n2
bjffcurxNdp1SZwCIbkGnSAxkC4F6kA0JHUx6UyMEmMT9dvEGveJSWhgG9hHp/eo
`protect END_PROTECTED
