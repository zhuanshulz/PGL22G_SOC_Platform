`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dR7FovMulGa8ZAaYSISDssHLK3ycKZJXo9PnzpG5B8UXhUIHkz7wA+Q4+53awx6W
miyPwBtdVai6kwOGHc8T2t2wRHH+s8Yk8X69LYvhZpxu5hkqa0rAMIBccPLcYAOk
Z2/dq1WysuOYPsTLA0YF15HBSPGE25OPe2a2IH7V206QTsJX55SApabylPOT2jlV
30oMtiG44zw2+7/3HMNHDrtiPIxvXA9cTI7Xhu5OqZKxsyr6ylJvXGZae0l63UQe
q0C7PgY08lOR7CrrKfJURJmJqLyRw+mewFxCSo7h/dwxl1AB8OXyOB8OiqBAA18p
0/QjhgegPek4NgozAf32SFeQeMy5V6hZ8GWNsnjcJEI3JkHFkqjNPwxCDI474+9Q
GSJl26BEabAoNxiYC+K+cg9E6Rsjkf5R4egeMeJfM/S5HT1lpFC0bcSIix5fTU3Q
EOCwbx0fFv8pnqD20QWTXSkdAIuVKcdtekPnq9WSsbPLjsrTWRov+KL36JQEnNlg
J2iehyv+pSEQrUnIj1qo3hRRPf6Dh8mEIw8Zoq299blmR0plkcy3RRu1tSa5HAxg
+tm6jWV/m+p0n2zojgOtvwxMl6CHdO/Q4+rLxhjwPmtRwCRrkjwSsfiU5xYw0HrD
BTsFNo3AZ583QLg+aIQayE1UeJgVR5Q4awS9IF/Ah9HlTff60iHRbZZubhx86syu
`protect END_PROTECTED
