`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eVhxjg5MQ0zmxipNwn88d1VL6CdDWwh5VezsoXKzpRpV3zo5iNvWDF2hlPgUauJ9
2tZ0dLHB11nVj+zrJmzhtMdjWlv3HFhI33bfxrsoivFI3n4qO32WssTVWzSiR4Z8
EHhiTYRr9r9eefzE1rqL/dNSXf3YLteWuGQzzNawbKxXYwbhv7NpG2kU8pjKFVWD
rnZYkn21NwNvdFNDsc091pVeuQubkL4KrhKGDjB2M4C0qg68gnbCU46DxpSU4i97
OIY+45HuXB7RmMIM7VxIWfSxPkHSd9gsg6DM/kTzLY7LkmID3Je8xYYaSoAxXVaS
zMBIds8dab1Arv0yngHrQLpr5ecZ0uBlSvk8xm2swduRHUyb1fPhlvdpyoShWxIE
hN/IjZYBdg858nGukN9GRR/jfmD2dR7fA4h0SSWwqDWbFM1Lbt9JqGFk/VIlGrZ2
+H2um14v8P5L9AFKFV1PtZKgrQY413MlWg5EcVKL9jz7SXg0JyKs6UFCKrj9crxq
XkmkHHW6q9STCJBRoBn2gYEy5tVNKumYOVWS31hqhxuwQnHqk2AY1p5IUXldSmLJ
7LfYfXbL9ZlOgZKArZzBXALClMe3JoQp6sEkaDLrJiIOGdfWcWIO4ISmNQfydXfj
CY/cuJdOFTguc1uh7VVMDdsUXZ2rgVh0MhnebZS8UEFZcj6umsMNXN49WtfjI9BO
8bHy+D1WfNWGI989uyvvHL0KbPO/kUiBaJgT+R9ULkel7t1bFq3MEwDnVP6BgvmN
0eDq7PDwFyzYkncWHpM0T0bUrEDEw8M9QqTtFT933FDa8kVtC7B4WahpyQIIQIUB
9587pL5dKW2uOZVeGLg5rgGgkeGnvBVFmBGLTSsHXkwKrE2d9MVCySjN+DK/4gSg
JMoapQjxrLT0Y/UXtFtkb/VcMQGB8EPJkR8lw1E0X74azmN0FV++kaEHEGPde0Sl
mLLIbrFs2cItxkyLBM6Rui6+XlfqIIFb54IbOPy9bl2gr85cLz4OUVBkEy8+syjp
bnJ90v1olxaPXoDr6C4U/9t6rj/ZSSpiLpTmVnoUb573NVPnkV2o1uD/mI0N2n8k
TuU8uZDrwTs6l49cF1j8Tg9E5vuKOECMqiFopX4GK7TXEVxBVg52NpPIPpDoyOLf
Vt2TMh+o0VXwaD/+NW4OwAxW9Ey0TMbGSKHP1FbWG4vYkGIyqNoqesY+C8WoiFyA
Blw/zCKvpQPcmGUzCbCWXZ2oQ3/Z5TfylMIWKfCEwkVsaHydB9CLs19L9bKv+lEe
`protect END_PROTECTED
