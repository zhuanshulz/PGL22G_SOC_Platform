`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F1yxSRFhF93Ala75fXVlGplEgafnpLQ1j3uzEgDOfLWh/3yhHv7vX6QuoHkAwOhJ
EhX9c6TU5glp21J7HiWzdsr6/NKT2HH+Jv9FOiUAkBoE7v5QRglKPqHG+Xk2lNeJ
t/TnvuQ1LSynuPhHgSMKNMsWszWeMggRoloiFh4KhuiupQRXSN/KQzxL4Vv8PjzS
x6KPuWKRtYOBM9J24B4YkJkkpHWp6k3UIvgXDqdP/OAgO65V/JiK4qenvtVQvxya
MhqrUwZilaZhsHobEznl96ttqfxhNGFjM6EYYSUin+4DTkrtohC7UovX68ZIDH2N
9fGkipjhiqpyXpH6S2haVU2N0HRnWWis67+DGc9U0EgLV94ibB8dPGL1vw6J7lf6
vTD4XoVPvpqg25JLr7WR3s8eD2pwjGI40OrvUcQzGYdJhw7r/Ia1hfdyQUJ3N6FP
16ISp6YVh3UqkDpr1Z4zIKofT/8monibJYJtBtP+mn+H0fSZT9jxORCN5+nG6Foe
n/7AT0pAt4t7mW8enOZQCua1F7HDQ3taZInm3g6tcCgu5Zdd29ksooS4FeN4bms1
ksZz3zzKpIokcHSF4PqjetOeW3z6FOgR4S75c/tkWLI1OLUGPSp3uW/c/YYl3jz9
5XjIULWavKk7CMb/nqhrREVkryodmvbI1fxO1csehAgc11X1pdGe3jUdW/7d28jh
tEePZKzCaZJdjMosRNz5wcKzT4cGuRPT/ywHHNnusTaYIgGxcSwladTzIHmgeBKA
S+CoKg7FA6Sb/MJkS2Jt0bmBiRX6Bt6F62Ik42zjWnE3C2ZtIRL5ILWWcVmgVkLx
sh3821pn/isDNVX1Vv7stlHLg7b7P+ca/r0ZmiSkeX7V83D3TDQW/X4XgIVQTPAP
0m9abzjBRi0UVLlFIzLrkvgJU42n8WL0INrHeEyzcLUr9wZPr1EN6HG87580eput
/uZx6j6+YrMVNZk3MuQNCG0MKC71Secz9gOtDtiXzGMgDdGn0Xxqc11WsztlXBib
/iLbtxqqdWqnM1x/TuNewQV93FEWk6VsUKb2Us1hR9thwe1zUfLFwp8vLggR13u4
GVryuCYeSNwF6/gquUd4H28XzkJiWxYaxl8b2IxoRiH1ChWLxjbEZ+10OkfLtePn
LPJpCSlf4Wn5ZO7GTc7eOD/lHH1S/i04vkEpSTvni4LePiHxe/hi+DQ3TucV0Upy
4zDyxv9XEtOUFyBJnbpVMGyM0+o409XwK/VRLKruvVHQ95wETQPopKbAMiOerQN4
Qz67crqJJwIUXRbxeB9Xm6rNpFmOKBQax1KwrcKfGkoiWbP12vLLOloLG3sBARnL
W6+3s/pFStWHP0Jt6e5ijOrmTLEXp04Kkl/beIh0w60Sv25HGTbOH3FMHBINEl3O
Wa0MfNYacfqzZzA5Hh9tJH+G2/zdtr8S+CF0fNePUEdPcriinVnAydoJdQY8aH0W
QZtiNuGI1Lxx1sudTRmQiatw3yCL4bqWaxmUtRGJ2Vy0BrN3iXaYR4kJZaD38d0b
AtWyWTXnQZplzNNz0f4IdhgJpSkCqINOi0iRgjPIfDVw2PkkdeCgD0GuRvZm0aNp
zRKNORDkDE8vqVKAHOsl29kfhu1W5Xl2TUypHxCFkiyH2icVsrJZJtFF9qnySQVQ
zb51ft8UeCpK7KQq5mORMqkDMb+AKHVc57B6h+qCqNliJoGzxfReLEJ+lMMFK7sM
PfVMmCCVZ/9WpjuK+/2RaO3+82hlqofJb6HzNS5Li2Of8JG3vRxFWZ3Pjbth/rZ/
DfobxN7ywHfNQLqMungOLca93A0OyzDW5WSLtpsh7Y3r7wb3d5m82mRKVG5cgdM6
8HB+s53raZpfbWoPWg+Ggtw3Rrd7QNEqEgbXSGz5wrwdD46LOVs/pePwYVjNGU8s
JWiLSoz599m3MdZ9jJ0DBojSD2DWhn/SKBkB8Eg6KsoPF+wbRt+v2krrIE6Ouxw9
OUG4FGznhjmmtAaGkeCCwKS3xJPhwasSK9O2RhstL02DSbLi6XCxQCQq9yK3GzV4
YAOEiijqY3g76gMYPcL2DEzzGMg7sl3W7V+o6tKZ1fmq3oHZEuZq4FftnKOMApXR
HesazKnHGz1CEUU3UC0U/iIe+YTPbKY2l4NyMqAUaVlBzRjg/yd7F/cEVUBugj3+
dyn/s9Hh1s/nrTZyzLSAqFN06FMns2BfrznDBAhSlwoAZX+ooYZ+iuzpaL64VYEE
JyUn8M1/s9OmM9i6thfiIK270q7C71WSgCsXng4unrB7hgQt7bDEBnJBTwaK+kQs
DGN8zPpUYPOhfQRqwll9VaZgQaXnLtZK2VMgQj5aGmOKmkNaNvCt4pnRW34BYDgF
L5tJaC9NvUUS7hqLmewPpEcJYRkyw3mbSOvAWWpqw8D9DaHTsCYluJ6WKzDEJq/O
GcnRSDEH/GhkFGFWpn3/XFRGIo2Akb5fo58Cr9TWQO5u9DjppTanaXefZfV7r2ia
sLbvHpeL+mI34HZFdWOecFtJ6TmGoRst7YTAdWyV2Mki1l8JOThxlgX2DhxWtzFj
sphuLjET8mngSk/79c/hhH54XPLPEa68fC26cJcrSvxQGRPw2MIO4LTnJqh90FJ1
Q8ePc8fAXySL1iJ6V777aSItgL+ZYX3eVaa1NV4Jexff3ji17HHIg+qZ2y7TSfUE
An/oXw60hV+9c1VzCqv13B2ueTlR7ESodVo6gL7KZJ5jsKjvoO6idg6S1iOnsUR9
kh3J5Qv2i4toA49UVGgv8rXalhsROBLohPq5j0zF9uc1jKdhQdzhwCNEllt8Lzzu
ww+hfUvEfUB171LAneMd1IHiGGKBf+fEFKGTyFavHs3sLLhegstvCSy4b59leO+g
TZfEoPPjJmkrWd0OONDOjb4Mj7dY5pEiu6rsqTfarlhnDUdZPUlTtA4LoM3GesOi
2WmjolWFcv0Ot+Zk601wjIuFsRLZ50DzewMshF4KYqPwsldqnUm8zLk13i+uEfG7
HyU++7qwglZOb8bOVgfYwaMXNrQo1TZLI5lZE+U4uV5NX+INbfck43VurPtqfK9R
MZAtHGLcYmwDFrT5eetmI/Yc+idwWNkmiY0Sh9R+TL4C1xyo6vOhqkewzWuv82NG
jNfVimWb1X41wLLvqc7DO933lSbJlud2Hm6g68iH6SbOEQugevMT/lmE+TkHqYVz
jTupa518zK1rBQQG63FGrD/joKVzDixJPbVSrc8fCa3jYIEdmnepQ+4ODF+5EYzA
yjDuRLh0h92gInOKxzHjRskcub7MmtVy9HagYmXfR/7mR0ZeGrgqNyTzyqodiOhy
22R+gPEXAnmIvvI6oOKrGI1TffMGPW41Sq+hRh7dA6pI+LS8sjcTj+ZdeYFp7CbP
nV30cej95mC1MIhTaEI+JN1JUOUN1+bLWMM84zMmhYfTYP28mgpPjpMfUoLF943H
ObKSHoS6GYs2sL4iZDvoG8TOwmKBRvVm1LdEAzFJC0/UY8M1isEpgeC1sHkclk7f
82PyEDDmzfgj0pwHhwjC6bGFNXYed79iT91Hba+WvARmKaGuPeuvhf6tkA+uKUpm
zjsPFOa4tFaluQSdXdnKH6Bn8v88W7xh4TVL5dsUdIyvdMCvWCx8/VcYh0TpgOc3
WQ0fyPQMztetZRkFaUP/EXPGLfxvbE+6ReFhaVNg69cWEyIicp7//5kJMOrAzqEs
ND6W7jCj25iPcf+o4770E1rwWzN1EPtyNSZMBFYaYo+2+hwL0vy3ViY49vuAjMH4
D6faKSB8MJOj1d46Y7Rv+wVb+I054Znz0EX9gqVghUqa1cz7LgWYBVjyjHoHIQsX
tsQ9ozb5a9dP0nOJEvIJQ0D6jPopWxVyAtQmwzQ/tUrY3arRjyMGe0QL/ST/ITbs
Q+SFhl5T1cV1O1KLoejzW3r1uMkWTieCbZqbuce0Zl8rAFOwjX4n+jEhR/XadFzG
KloKfRzQEPTcncr3JpYis3auLWLG0U9btEncMR80vAnAMaKXFHVdosy/PLAR9mgG
UDNgnp4ezkHzbTH8Pehy8X2xjo46Gy5HjmNEZh3uMlv3MmH4QhiagOKS9cvc+Gnp
Gnu1kh60BSJxQr7GkzZ/JZ1eama19BEr9uePoSYSzktTXHXuPruwqltnvZD2UbeE
ABlPG8aFPT3VkNcCMnYLRYFwW+dSVfgxiNJCh3vu7K9MsD9e8A3wa7stRC1+ibJo
qiQWewdZ3UGg8SeMnp67/+uHPWVeyBA4KIubU+er8v1sU7+e5ZnS2mdd1FrhDVxE
BDDoxrXQB5Oq1zbdpjJj6UEK7TWpWjXR8AyABsRaf71dke8mmbUCYvfTg7VKkRc7
4+X4krO7v9cFIXbPRYZtD1cXmtJ1l5QxvPcZlsL17t5wBzsdHEbA7YClOVcIv1LF
Bh9jvjLQzKcuah3DDApZdKEryh9dIkiMcGFECFTgYawH/RXGg1gCSWJouBUxKsod
6qW/qTc9ydw04f0VD4MXIFlkxKkQopq0Flr0lp7wwj8ysgO00oSSNmCBuVzHiSuK
M/k7Oycr4F0I6vA4B8TCPdGES4AJ/iblRNqULrQ9621y3o2v1UnIFX/BGfmEKyl+
xejjyUA483gy73nxSOPsvHJSrFoWvDE/apXRR/Qr101Sq99dZEsaNAgEKilTnQ+Q
pcM/JQYoMsGYfGRqayOv9X6pbKuSYmo1lXBfTc5Tua/VBeBzbdT37IGZbiFh6zEu
fGqguXmYX41mk7Y6HbEYZSyBork7BrHdNyYOHVIUX1J73f7x1XnQ3PXjP5OfebHp
kQxKMjrWPTQs5iGLOxOz1eMaCXdazQu3jQ8IoCjmM88EZQDrY3C2SOe5aa03MhAc
PixTVJqap03GTEkoTssqaWdOpYTzDBuBAB/1kOctDnZ7dO5iyQS5XLaacIgKdMBX
tPjbRA+bsvVCX3mMPom+PXLr//Z9xy+ZdGgFNaj2x4Db8ERaHsfgXh8Q0fuVqzCt
b0URwBWBjJhxEY0QSsDDl+krcTSzmGOB8q84J1MMPtFltbzBAaZM8Oy3wEjnVBxo
OpS4ootcn7NEX8i0Rpi1KA==
`protect END_PROTECTED
