`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XmxTkLXsMVo9/ezOdYAizx2DOAAX6D82XGlpEKKAGItt2MwB4bfLoTDew82Mde7I
YdhkzoiLGiG38eIcKzQdQDB+y1lDUoF8ytJcGwGKnbQfLHKcn8wxRZdtV8Uf6krb
vIXFfbZ7LLpUX6ApyDwZkmC0zFZA7NIAoaHEP3mgdCu4IpClTkO5Vedvb7RlxOTG
UZRilRJUrgJK0Q8VkZtPDfNv/N1I78e7MtlbSVRiG5U7UlNnvh/wj2nzwXJYuSgE
x9HxIPIycN1U9139tjyARgk5oIKoCWEV67KGzOTHwvNUwhwEe+9dmTfny5Gh0iAT
gnhKQYrpvDdJ5YOJwMbcJW4Ts9Ph6C3zhiXP8Zb/gHavqAsL0hSldkQ0ejL2p3jh
gvVlX5O8WXsADobBC98w1Wz+0nQ+ZyqXnOtRjAgSziQUXjsLh3Oa0ERrnHch00NK
UlCWsPvq7jNerC1KehfE/VpLxFAa2DV4YgwqrSEEphSDfSW/IBFAPem/gEUSMVG5
zS4+6lspnNtQvFI9srDjVcynHwCSWLhlgwdkwvl2H8fnLJsCU7dudGx+l2xF/f6B
qxG/JsgII+awm9aJK7YdyVyIFu1OBNR/zCcJ+QIHfsvEHf9EUga0O/PaZspTmT9L
K8tuNRObVrEz4hZFAqVT+w==
`protect END_PROTECTED
