`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pGWL+7U9fjJV42qPhtA357h7NZtT+a6qu9iSdU/D+TOKETTx3dWnTAh0J6YBs+Pu
W/MLiPoj3bSASBY0cIBirbKGGTzmDJllK3cXa+Xu8vml0zRVn0y8lQdfRnt/qgPq
oq7pvoZvBwMQ75xiQvwlHxtNdhXF9syfHQxMv2dxr8gjCqVgY62EiY8Soe3alz/7
K6XNVfF878uWF/nTv45svarmmrKWf4FuMfYpFkwsOHFg4qKUtarMVDGiUf1lcHav
k8qfNvNUSzdaH8IQEiFDK/cp09psyTOGr+oTeWVYYdxr8Bzgtp4nBb/KEXgHiKM0
mZgJUq3IU6oaJvoUxXlHow==
`protect END_PROTECTED
