`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nF7ikvTK10xeVcVyoKHodF2x3obOP0Ew7TKxdjY+zqsBNKo7DErvHkXjGpOYtVIJ
5VDN37n3f1Y8d7ZSyXCQjOOY1kSX6jCfKZH6MW1sO8xhYLi6VXhiVIrzp0WSgh6v
N2sxG56z7rGPYBsBqXYU3111F/QHmGRLH6WeiXR0dLiK8wm8nyo1MvObIOiZeUrj
lw2oN+B1f/Wgy1cruBxeYaobc+Wd+asee4cmRXiTxIfcvnZbatBw9vChGVXY6459
uHZr0TsSEKzR4kzMwu/tP0FmLxOTwtkyrwow2McW6tKeCblYJmzN0Kq83NytHGA2
TJwLPkCJEqofYWid84/FeiSEg/nw0f/aFHSy0Hc1ckYqjzj6IoXxeWMkqTCGUTpp
YBfD/aCF3tDvVTciFuGYOT6FUMj89wpGX0MrkJmnaWXryRuA/Ej8xTwCM2DFtKNQ
h6wosDrmlGIlwPrwvREDBeUBVBTshkycXPq+A9EgcOKVqCIUE4O43Au5NaPZ5GZi
x73ZQ6FSndgyNiKIZ0BhoYSaZEJkmUXlZToS2aWjcqqS1B1DHwyG4aoHGvqIhTbt
SgsYBpRwvxVnwblooHawZkdQNCPhBivimwx/t1NU4/8DT2jI4qRmgRFY9XVE4tCX
GsDznOVz5T719+24TIG1O4TvKJ6MtCE57mfZFWkjCZE2uyQeK4tlGTVFCkACEaZ1
VyEN6yrUpP9QUndXifzbVMgVsAqj/5TCexp8QdDdyT5umtnztgik+oHtEe4RChB4
WbCllvSiMZjkJ4BrUt7JLkmZeeSpMWbc4EXaCfRsRk2DdaOay77p+FBhvKC4hPft
+ugPWKUBXWhmJZhGPsZiPrZruf+YMEKwva+fmbrsWNKF3tI2/F31oHodYXkCvXVD
UPO/bYSoAxL8Ddw8ryrss7xUAF4GispWsgTm5ObqoK2ig3ofgk60TZ/ZEDDxAZ1q
ZGG1BBe7DNlwIlsx92XKY1E/DSYwxiKOKm0N3URNalGOUhEyXjzARr39MAVt4FCt
5uPqxQCrw2fPTV8Z9BlJiVRvd2HYXrSFZLYvZlTu4BvAAHVdFGlVF8tFS2pKXgSW
DIfxHRSJjPBvvc9+mNVnb/8wTxw58j4Q3VfQfcQJhoHiUhg6inMpIRq8igVGWNdg
BZmpXTjvM7UhIAtKz/7goshzLB/FqkB/c6MElBy7KQ7PBAO0Z85QruJfw3kVRBmW
QmO45i/6srQ0QI7AQcmzgWZU2vEXJaMsTgf+jt79KYrpQsy047PXZHu2s4hxFI1U
+Ap3hi9vXFPqKDnokPHjyvVUJuL7zGX8uUagfdbXFB7DXSKi38UVcwCVUOY9Qow7
r6cbcFvXK0XwpaVVP0uDEmE8v9g0qaBZWDAie5N0XL48syoLljtr2qS1gZSwWaw/
EuXjNlsEMTCUyksy1nkWmsOj36rRDW6FcfPIImRl9Slq/NlUtTBaUwLX4IBvvBUW
TOm+46WuowlN6l44QlE1i0wr3rrbLC0GPSmHBNWK4mVTNRM5Rsh/qLnzNOG3vCcw
5EzoP5yxtPwGZKeqcSlXz+/Z4rL8Z2yTffeaqGjsa/RZ++22XWJ4MvPEPmdiU58E
WHZDjRypXtDy9Z1FTryjaKNHs2aGKg/5OxqAgn3Qt9YmwBcd83tnhROfPBy9zspG
VEdkWR9e5+dX3boCPqBqbheAqSuAfVmM7EGJ+9OanFF0D4QnS6jpim5O2C+pkLuI
yiIgY87IMQ4vwn/E5wsSx+C2XUcftTCCvtgBuwrDKrXPV5ILg/xlxQX+8MTOIjMp
6yzWHOrFqWrdLsofewwi9PesoIn9qJ0kldi/h+EiUJECeArbRds671SY/pRLsryG
jntRQEdN5jrvk8MBykX+5f+uhsxkxHRj/7aEsp/fykTHicj9q/1E7ehVji1ZoZZR
ti/s/zrj3amK7ueL+BqDNSIOYUR7vJNamEEsYhyDIhuUnjSivodhcOs+4ZoM5Nyu
mevTRBW4wpZODZWDG5fg5h4XfsPy12xjH5MtvQIg8DhQiov+35bC3DsDkPZxqs0a
nHYlWcPAf9N6yJUTmceRihbskKuBzGhWhxUbOJKlQgDgbyu+FsuZcZc6NACYFmb6
kqHkHX6Sl2LcJBIcWIPzUEXzIlMrFMBhzMSS1HY0Lzd3Saho6wm5CGJbHHYB8KGz
zytDjPrZygpaUe/GMZOeSnqdUbTwyZlUxxG/2j9lwKrgtbJ2qJGWbdYW9PmtT0Kv
vt5WyJMT+TrwXoeGLEDbYZ1XAHXxRVtdPFaZbXsz0iE9wxRqLKogF4sekMXDPPb/
Avizt/qIX1fXguaHBjB0Qku83YG45nu+BUMX/VBL/rVMBF0ieuKP+2cNY5t/uTMt
X/2ISPb80eaV8T9uzMNQL287Y0dqPpX4Le0W6q0OyXTkrqlp14wGBOMnJY3zuJpj
Wm1NcErNgurk3pWqesDZW2q3I5tKx0n97vIFzH7OHptQvB6I1qJ92KPphfgmmRPo
wbUN/r5vsrU8R7livupPhhunzsMITSJxU3aX7JqIeeLbvbaPWc1DDAtmo3HKXJhD
MP7uFKgOSe8moLW3roDA3KKdXZCsq57ZNmHXy9dQrgh06lhm5wtSnB6LNB7it7ta
2FrZUlSlTJY1Tdd0SBJwdx9bpDXIOrBRwZmgKKL9l96yVR6i8e3C75zViI5x3zh0
60b/CtrZ6mSfhHvEAQXzkEyu5GZsrcLAJJSaA+/isilsgjZh7ELejIM4CLUB6elJ
86g+RN6CvWXLBu49P8M49WfWH7siXd+laktuf1936NeAAu5gF1FQmQbUP0Ulv4Mj
xFoa87oxzsZMLpODPvTZ8oJ7Pl1aOJ4/Hz1Ndp2Qej5VRjusawlCtUr4fXF+Qhf2
jcnQ/rJ9p4PUjbDQG/6WDuqxYh9ohIgzKLy6N1p4kekOjcKy3rHRL4Dp1hOIBoEG
5uHQfibBUIZBNztz+WQBJFbS9BHqfddyFZDcdUav8SuArpfjP3k8U6zzpM5JZFUc
`protect END_PROTECTED
