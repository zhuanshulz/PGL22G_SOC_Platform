`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0VCnNNLA5flbY50Fjjp3L1wUFOgthGuVDZbIkO+IPfvco581zzWwn0l2MYmC/4YB
z1rBtKVKnXjJ7EbCOP4PlZQzqFBDEV4bk+0gwoeuFH2+9ukUvVGVp6jjZptbcgUc
FO9ouOwlU5v1QXfHYhlxlXi3Oubx40sZmYZb8qfFM4Snw5+zSvdm7ACACyGblDEd
1ea6kAoMSnksciSLZEpwC31yEoYV1KvsNq6ExsHYG3LdxD2k+5tobrxo8BGETDzj
rulF1ZKOLNvcwfqX3SVVzdhyJI4deb7ywHDubf+IV4gZRo6IpzxHbmxah90nFSnZ
dhr0QDYGRQLoeU0xBO778EgrF5PBAAxgZZGIu9QQGmSbC23rXO21+3A6j+5kszoU
7TFFfLKLVduXZXDxp0f6e1foesx96csZCffelSXOwRdXsVQvXEzxXGiP7P/Z+MIN
xe6WmX7dUWQ47rzBW4IkQqwAi/FGK0KLGV0KeAe2w2BEv9s/rXGHhjpwjFhBCCMh
pZ22MLL9l5zvDc45R1zRAMuEu1S5d5wwGTeZzST98v/kWN1vTdqsEIxwtpPUbNMb
42Wqucm1P02XDCfHmDH5hjgteW7yrosoUfYFH2PVix1W2+P2n9Cl91tyzl28nvrJ
FrnVtnzgRA2IA+ASJtlv0cIxIbXpbfQSaaguFDDyagMswjmkFlj6/BUHdHmut0vx
rKd9EhIUnt7tI5WanQJH6X5X8zZIYKOKEDfqlDuscIHSX8xov+PuwEJCrRFsI7GK
ZVf1m5ujpAMsnSwU8tNRMHE8Dh2xoknJBG8Fd4WT30ykOYYl2LyQmla+yD7Y4Foa
uC/8UYsNooPBaHRZDKwjcCG/Aw17Z8LwUa/kW/MF9k5NgcaWAJcY6i9I8ncqtoAb
Nc+qoFWKlqFRIFl8QCTbUA==
`protect END_PROTECTED
