`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0khySxJXRfXbc4Y7iDJea+qYRtZc34CcxTkSXUXiqDh7ktncm2r6kuoV2nEcg81h
XNuafLbyPX9ttDP9E9l2xbBg1vYB7rpt1sYUsdsw/54Pk4/G9EFrJKG+kujq9KdM
A8zCYobTxXIGmNHFx2z/W04ZM4epnrOeNQDbsp0Z+fEF7DBMwLbsAWwZs31BcQHu
67xkZPg8rvoo7PYl1bGTDgxJtg4Qjyi6JFsRhpvjGiwNwESdp9AxHdL0T5wM5lG/
22zscJkEQLGU/nbbCzNLs9tCAVAUrVeeL3cuCsJOBJ2XwkaD6CXKOZFoZkC+wloK
nNnxDalSLTyj1kJnHhO3sqEY0PTBkT7USL7AbQREyHpbYnpQu2D1GLLW80ERtCDq
g4ckvOfMYLgzlNjbV1EPqZz63gPvmrnGy39vw6p31WMvJf/CYYVix+SDXTYy28VP
wRkO4GgT8PcX5rIb4RpeeKc3xHEVC8M59/zq6lEYCZiECdh34EA0OjFdxw+OseZ6
UEPiDf32fdDFeCUjR3g82AeDN0YQoq8KfdKDFAev29OLcheCPiBZCQ7IZqjBCM82
0CaMAK7O9yj+7bSP7Wq3+lLoPaNh4T0RVgqkVXuF2vtoCucibEkYa+vVlAMPC5N1
UZutRPv6WaOvc55ziMpJ5cQj3OijIIsHuyXh8kUkkBVtmU+eYKyia4CA3bHH6/pN
hxLED8oPb0ojDxnuwQGRcg==
`protect END_PROTECTED
