`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lY4EUvbkAwmKApwkermk8fUq9+gNSOaj6ZWYgAhAn/uz3Xd1ssOvoQu7/Q2TR8Uk
nVlsQddm3Mdg11S4/6gZsZinpWs42HqL3hcIh//AfG3rFR7cDS9WrOjLp3H+Aq9c
IiQhRneYtda5gaU+UMSafl7Ci6LUdzX1bweKK03Ah/JynlDbvlVu1ukYEbMiIM1B
7cWZL955xQ/YnSmlbgviPxibxy2+HXWP/voj1/h38LRxEui01D/HX+TZGFTbYZak
gXFnLcm8SWBvEzVxa8omTVKlkVnwTHGjQSzqk8apT7BkMF4HZajHVqO0r3wzNo7U
gd9Ul0DVxaTWyi8vMiV+gBaoQE6QJg/HDFXgB/LI5ZKNo6F9RnlF2cQr6PNMEAHz
Xs56I9D25dVIBVxM7YFIqC+fafPx7RB9ILOOOkOMk/lQwjyQze7Y8iRZWAD8DEbZ
vhyyk6U8EPV0w6fmNuY+8kGD7GJ9SeOnxEaZhMMf+bXqFhqgocQgIWGWu/wmfBZj
kPD2AV+TCXSkPtGTC/R3HxpngSnUH6rYpuxZTpe6kAuAKZX7Suk5shGSMRRgoA0d
HSQBe5m/QjwerH95rLPxN/3KBR4PIxjc5Yqb/V5bcUT2e8RZXTWfeIGg2nHKDhq5
8tIoDFJ9Aa8PZW47xQ90rQFrJ/DKCjfdItlakUR1bZw5zACclFHeux1G7PAHplru
NKGKRf9UDuitspks0ITbndYLf+nXaiCVvjNUeMie3hZHVTNSCEesJpXzEesKlYPG
mnWwvFF4+AZOQ3lMkLKUx0XfZvQhQ6wIbZ8Fu6ltDDssQiw2E98cn/D+Ugu16+sF
uiwDoPktp7XLDWSXI0w7qVHW+mo2l834N5/aAyJ9TJ4Em8nUxjzqXQfvo0/U+kfR
AMp5nJiwKaPPVhnt87UfD9wK+m9ZebEbkFksJCXKrzsQEBI4ID/Y8IvbuCZABUFJ
5zO7uQYNNTaWt1XigrvBnHPom4tFuuS3el67N+XJyZ4jKrBCVLEZPTLgJtQStL21
vLQz/PM9yBbZdAxkDh7iLX129oCHqnYLL64qRI+fZ8FvZfGaIJuHLyVW4lGqN8kq
hwQWAm474dEb00hBke/dKQ==
`protect END_PROTECTED
