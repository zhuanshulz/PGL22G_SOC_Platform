`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o976vpZFhYobj0fEx0IUzA9e2NkD6Ewtd16Qm6I4U191sWBNAl2fWbW/N4531l9i
ZgMo3A4oELU2wg68iHkvYv24AwQCn3u4++m1FCEAuByn47BUWExNRGc3a+ub4CBA
MSV9I0MkBh3phQewKsPmWKCmAese1Ag+FT7KH5Y2b5RgRoHGhSAdtsCedt/hCwTa
QDq6NTg2nNFHuJ7js0cd81CjKJDlH76Iy/l0ZC9UAj7qvO7jAPt+1O9IGwJ8hQuU
qlw3W+g5yLCapjemeYuTA53/oOXFLN/gIiA3jRxo71jii383HO8wCYETh2EDLO7I
HvEzawZjZnUDbXP8+2trHYkFCtP4u82ARB2Wu7nSvQkGGgv5WeI+L7u2W88vnkM3
F7qfpeb/jaXkLNqTTZGThU6wzpr439fJDfEtQU6QDaTiI9W/85TCxq7bK9xCkWr1
IizgekV20W5Snj66yAv61Geh9/GIdfEPZSdV/nyO6wUcgdoO1C2mq14G8yIkMYAg
B5DPcY5CPgujFy6GJ7OsD2XcMUAwo6/OlZSwY4HRa/PMZkbblmbqV3Ti14gCX56K
BlM0ZXdKVgq9B+NFf7OulvQXKV17rCW45MAhOi7nv5SrMCi6Zyn+Y34/uUTdzrO1
8HXe89ONKi8cIfArp7h3YUDSN6bb5ZAmadbY6WT8j6lqUdYovUwmcLNqQw5/mBYn
MvZD2Xe1ns9Nj5cx88y8fYk2EbxEidX8JWILLEU9V4KBqCOKHZF7t8CMIXD3vkRR
PXlZENZy302Y6YyBSKKMVvZ1Fl297z6ySvJ8CHutaa8A+ySWLX1YiEHYJ1rHVWO7
UAPaLatDNNOOlcF4StceO717JRRCfp6x/WZEutO7ukvKixPp+6mURQ+nPSUyPElj
8jyFFZ//K2CTEWBj+hDdcExc+VQ4cNldJDbaC0Cnsd/OwBQE9xlpdFM9Ktd62ZDU
2niRIW9lpUo6yR3cKpkMUSj1q0XJHoiyOYjC4f9hL4sYggnIa4L/ZmOEeaveFDOp
tQTiG4AQG3iF2eq22kQT+Fkuts/EPgXc63fa/GS9lF/W5sqh6eJAv49RnPMTu5or
OuDGsfgNnaFRvj6vYBuQd/grXFzl5jmE7IoNd3hNUaRtWvvJ01LXZuAMOPpArfES
NKwfWFhqg+b71YWC/bgb2J+RZVDk4aE1HHptiGlfnsobDvkAl3OAQ6a/cd08fqCK
7/rMjgBkgVimHz7gaS8zAlMGTYA7fHgxBT0DYZeaY82VfssSLOjPYI5DJpfoqm3Y
Aeu8Isq1Z0pofjIHiDANsplQmLNKLoN00dwMhCancyddzx6tmOYUHIiMnwxYyVSB
qMcDyEmWb1+5EURjmMkzkboi5Xp1co7HhvFOQmbtvaCvVqrp6BhKT/WNrqkBe6Nw
GSimIT6YFJfby+K6Y6i5dMAVQKyCVYQ9UQvnX5w+kcAL0zL0tZeydUdqSWWO58ad
Lkmb61GxsHpoREHiDQgC536tsOYj6/L2A1W6+gr78/lSh/L2Er3zLJteC7Rag9x6
GzZ9EqNQj+gBDAk176FrbH/ImSG+2tg3iyR4TGQZhedikAjZTo7Lg9dqOlQzNgT5
Axa899B0Jn//ChIibv736QhnOtL96Q/FCMgGXiQ4exFtMqq1DblZ5bNGPWgrnuTq
zCwYq5orznx/Hu4lIdafSOUrPI8AwEmR/WIZwiC9eIwJb266f/RpVYccj+rOYHpq
td5qxMueqyeACPraKDaQYT28lTra2TMRRnW6WZY2f9thtMNCURbHdsbfdDUBxQPT
vHeqx5VPCLFbFCBVZ+GHyvo5mH9YeIP2YNVffgJn2v0gZxckW4VYuhGj0199FcCk
6WLH4N8tC9ZYx0lgjnU8ECpB1AOrOBBkSTo0WOO1+na8mX0rJLNKlpATrku6gNNG
6W3lVo6TU86MTEHULYPtR5+K3H946NOYtOzSE8ucSmfw/KsldCvW7cCKJ0ggFnvm
d02aPtLPq9M4lH+B3s18mAbRwiUfNBINGtqdXtf9mhPraPbOKNbFcQko6wQCE+KD
bKmqzC2bMIFQXq+2S7RSo00CuoJgUREyKsrs9onfLdZYkynvXiF+0lCsW5T7S4uk
U7b7fR5NX4zg6j91DNC25n7eSXfj+52/ymidXkO3pePNukU0PnvhGOcWPr0SIVSr
C5UUaSjTdH0b9LEkI7oa5/CJgTxp7f1bLRvryozOwhWUxKOOoBxnQpL78P77dIgU
lonDYy2pNokhSHsPcbRY5ECrzMJykkpPootpIi3tsDBl2j2MDdmH1cVmXbg/qBfb
flzHPK0KXb7fE9Ns0OiQFnfWktIgWyKXv/5cBLl6mWADokhhjE6Lu66rqzT7yTDp
6y0JPJKI88yADh8bUOFYuw6cUK5ZrF2KKp1SBh49tlEdB9RTwP9nDQm142MuZyyK
Kdt8eKFJPX8eyLlkFvEa1uDXx2ZymXGwq/0JKQ1GQLYK7t0cHdztBjoMSNcwhy3w
xkavKO8Lnm1XAM3V+BKE5OQgYsHyvcbQF07744aLuNJCrQKRqtFaWNhjTJzmFB+7
kFhyWd6creMDiIFIL82Igqt8dTBLXFrNtJmv5/cBNOD88fZSB6EgECwY7UmJKify
rv1oMCeDlrN/ay1PjzYi99B2ePDy8N795JaBZdXKX2KkoquzdvCJtcJfXwfqrWOm
U8LCZXlsHCLLnQkpNkYtp5NNYjmi9vnddfUknqYxlzUHUzvx29pP7nBHuRg4BPQt
ZAQRIaGHolzFqxwlCF//EsQpU0QEuwcMQjeZmA/rMTZKhNoGyyVtquojiNAKpAEx
wW7j8M1pK2CkvPymIcJrtCz3SV+rRkzZCldBa+DC0OK81zkoHvsCiqRwrAa8dJCe
2yruToixQwSE0W76hnGOcFYy7VJn1JOGulsNuUlb+OUHwpOMWxyBRvtgjBGUba/d
ROi25feIcleDJe8ZUATW0xtFHHhkv1s7dXrrQSnpOM6oEcXZdAiVthoR/oMaBT6S
jbIDU33Hi0gEttMxOyYY0L6qyuuP3XtCLsAaAxkFiwUE5aAShihTbLRe9PVnBAcD
YRGkFPAJC6etIbnS3CxC1OWU7RcIMtfpTlMeaWITyYxzh9UniILfWJuzeLJEYWjT
rlznjSKC5DC/7qLUVHL/CE7xWKyvPB7cc2TMLHddmjJ7FgK6DuG7p6R4CiUYCNuQ
BXIpNERoL4VThdnsr8voJpD2MyJ/Vz2Q3/qH/a/n03ZMDAlgbaK5vzHf1DrlTjwa
m/Z5V30gzt14gUecOUXCH49fDaDVo5uhvfLxJnndM7LLNg8QqEMNNS10rFOuRN/s
8wzfwLWIzhL/pJeut731wTz+wIsymreb49nSAbD3jK3aC1squ3P1yVh6ipYQfD3/
X36qXf/nJd83snWqCFq4MrybkMM08M3ut0enO11LggwwaayXjWhdb72ooJARxAjc
mAeINxAATDcL0ehaW44pkh0TQqaXZZc/+jlRCTFgBHQs0NO2xfZzqUBNJZV8cv2z
pC+6whDO8371HEZplYMsJi+ZTDgTqYweVBtJ6AHNORHzrVxhIbz0K0Essj34SQOS
SZR1ljn6BBuyE49TZWi55ukUkOpH4FBCLiSHv+TEi9ckg7emikJNWorre2mGXoL+
jDOfSGL7XmoCfS2UydGC3JekvX2jANDk17U2oCfurV7XNI+zHLQhOSaz4RUVufHj
Wm1X/BVbj6CNg6sJK84cLiBeprtv7/cChC5/IqLafWJ7cpEi1OmM0NaSAnr7NhhY
lRlgFnsr7xiixlT7WqRZvig2XwtN5AWx67YI3XZJt8c+jMg9oHeLyKzTY0wqhA4O
LGFXbZes370WZSRW36ISDkbUwWsbj6OORUZaULJJUc6QPejZ0iii3vWZdD410Fay
u7a1Dsmmj8q4NB0rF7H/oFZToBv3Ri+QDI2FenSoE2/1+/+X1sVlDA+PPx9em/K9
ufhGKfo8XrqQ852rdsd1rxhV5ljm8VLz+PZn0xztcwm7kIqyZ3EQAb75BxDKKsYi
Gm3lsTT5UROj2HgE/A0keGl/AuRfDVUgRRMSuGJ39HRRwuJHuVOByaDoQbjeiQgH
Y5L4uVxNeWr/p1JpMlYXBBVrNiwqU/UPHwjBLYfYN5yx7Vz2lfO7atdFtakyxAuh
A3J1BdAHUFqUt5MxZd+CUBNMitABpkxYzMwTkSrngCJ6LCzyPgVMvCCp3VPBfip8
Bzr2GtBUqxVTUDRS95wnAqCruY+rWucCNVICocw3XwlJJmtBq1Vb6XOffdPFvYwP
TbCHNON6Rg3EK3dxejD+WS3a/QnJ0MMFXMz+XL701XriPAkG9v8epalRa5pjuvLD
oeUY8iBbuc4AoWpISyQY1ZlzM+PYeRupYGv2wFfKMduDeHHK0reLggW/gWkwWhx9
c7Ui9JO3FojvYYnloeIKM+Dt9pXln6sjx/EyE/iA2NDWXr1eFuIgAo3app23lX5b
6mIXrO7cYVZmFH3KHxMQFsGl+iDPEayFUbv3pdraGsBNV8wX4otwtrt7k6y5EMEZ
O7oX8Ucif6N3z9ucKBoL3SyQjV7S40hCpYfDkrfk3Qa30HrkrgWnWJp7OWBG2Als
ipzRAd1M3qihFyG4/0KtBFs1HWaq43Zr07aL9adtIzDxT7EDw6aYG33Irf0yhI7K
HBP2744/Mrp/3IBQpWXPOT7/SX+tYlWSxnfmoWTwtnOXaGcteoL8aGrgOr9MKfV7
p8UUM1JuL1xudL9cgyB8cetuNlTcbCtbCQRk2P7zDy2/ADDC0BwLldiTNLHz6Xn5
eBUAEXDcdqwZ5ayjnQNZz/q0Kg3MLrYWScjVWeN3pw8uDrgSDZpZxkVg3xpuic4W
vnhjs6IpPdluhu35rV1D4e6M4NACE83BgQZw/DwAGLA64XcWjydmjORkU0tyH3Pe
iCiE3nETR7hB7Z9rn+NtnQWJWchOtI38Q31TpK522AtZl5EWd00ob2YNiCk2O35U
NtqaDVMNL09J3nuR2Kq/7gQzdoSWd1bUqnghxBEnKmH0y+L2fbuiiXcopoGmX+Iv
HrzZg7AAajpWmDIKewWeFAeZZDhQCUlR6Tld/EB//urbakj2KnoomGGvjQ/u0BUl
rHiHTQUqBRRdPnCc82XeUqxUTbgbfxip9Lj5WVHUmGwNIUst5OosGP6DyMDH7GXb
Q65Ae3ZuLqTg61Z+2FDmoUSUbdld3fDQLliQdeb0ch9yctRmKv5yU2/aH7GJJn/C
XNcKUUOV0x7fE1wioAIw4G5Ast3okjYfHWj/OM4yV4PlIC0X2QuptLi1v9LBa96/
5m/+rdkytpruXhwLVzqldDesUpIy211DhxyCecWDapeHwuUa2Uknfhm3ikzRb1C7
1XnTZ0sVZvg+UUYZ/5MKhufW1U/R7NA80zeiRe+TS0AKkNsnoZIS8h/ar7QijUh0
bi7i/fVQFg5orjn3gQ1Acrz0i8iXIkQTqu4/T3+pzV1A19sNXO+n7dlD/6Xt2TeX
L5WUw0HeKxqGr3bMEVSKaLDxH+tk7ZKdhB6qAQVQ163/EXO6yAuNXG4xST3H1pKf
MdgWqPkpL960A2vsB+x+R1hBBv2KusG0nwl4iZIecKHKeTEvvxQfRLeZH7ZEaJyX
Samx7hZ4nL31zWnmXABh0QSwD9Vst+pByylTR1Dxrqe49B5sN5KA/RGEoujtxvWs
gsxUEL1XHKbAFjY5v16sg05mTW3sJb6hx37cayKDzjLsKIT1iJx05G9nBoQey5uf
NKCHkv1L8x8jBnWlVf1INN0vvrFYziBv+DaA110myOERQt1qrUK8LfwxxVTyWzse
7I/2VmkogcNDtc0hZFS1+BzSBtmOsIc+UW+ptVb0dt3TaJHKPbOa29ojFDiROe6u
3OnIaU1dleNmUUcQp6R7lvOj7d4F3+04xABRsP72QsfbmNn6ohzk4mUv7EDLsGb6
XOza54ibB91ISA0iaVE+W+MFLY+gLLfs2jmt0SbK3WCW4k/5aBFjQIadwquz/uKR
h5UrivFodqW5qByrlak8UFCS1fxKPfygljPQWaX219OnAkDOzuJkVNYH//5l+Xdq
2RYSKoADUTQRzrho8JHtbPPcVAkb6k4iKYN/lc4KldbFcUnwNbrqY2+5i0THbnUP
z9dR6nylLcc/fW7Qs0L+LePqzEPUGreOjq+qX89BCvNk1XD7pBjLj7Bu3m6Q4gQv
q8EWSxIJGQysbe6ilmtthl7CgSA2gAFEQKgItnJAfU9LEDX8WjVqfS17IikrKHgU
wfP9TMnGIXxYVuzKDY7xzjEga+/gJBrfCYHR+Dxs37j1trRnTzEHnfB0a79jTCUe
IlUHAII+PIeosRPvc6nT7u3o/mLqD7tRgDluP/UE11DahA4GqkZwLgUfe7TsKVrG
fp9SEqrwsVqt1arkvs7Iq/kRI4cCbFfJUpW1flgFkjRtRulgF6nBBgO0nYMo1oFL
4t9ocLKoqv5/63hrCrq6yWfTgL2qouA0xGDUEn6PJFc31dVrImKRQc5hrfv7WJCZ
9GBXsrS6V4RN4tJ9ElYiAq8FyI1LVUFE8fo8IxqxY7eZAR2bSHgIjHpvW6wks2+C
lb6x1BWvxoNYNunUIdpWuKYEk40dV2SsACt0DA/jg1OPUCKoXy+tJXzoh04YGdul
M/LdBAvlili7fTm9jvQqjH06hCreDp6t7sWn7N5P8wap2i8eVZIzfhpIqRzHx7Qx
MXAEjkJs64y2tyJit5FLDn2FWsQCYQhvNEwqAh99jfEttabSbhnvIF+8AyZ1nZ18
xYQWYyUQjlaqlJpJgV9MeffHXvYDF616oxUxro0rwZJ8liUXm+XDZeKgAYnA2n4t
Bx0IHrANAf6/xhzMbBShyxkWcohZHPrDmwIHDOefhnNgtyH+5UKbyNiCgubtgku5
E29F8wq6UrhJmfepl6I83rF43HoD3uS7twGhUP7wd4HHe9bsPrWrNE4GsEpz0f6E
AzLMkoyDIdq1KQF+i9C3iMaZm2WB8PKmkPEdMsnBLmrvcdIzFP5JZTyiOhhBrA4O
VfTWWo5luDKaTpEVAE8CZvFGc6QgS1GJKUmYkyKokFYsRJTPLZ27/C2wX+feONfK
egN698gyil0mzDc1qk8Zj/BhinTwX90wMe3l2uv+4UzZ2Z4RImCk0RUkuJWNTBVZ
uRALJge0buSJm/GNRua9GoYHaTZpbU8Hml+rFqwG4iPs/U4AsU+bzVgMwrm6i08L
7DQhHCL65Ix2m3lIiWELnv5AgA0DSmPHL+qDNL9PxD9PsWpuO/Q2+KKHDKfkrje5
r21/F0hAwjM522486xo4YYGPic3UkBr1DEdM8kPXp7G5cJoNJp+vylw4x/9E2zh+
a+N1lGp3Dde9BopP/sPmByx2yAxDbamjl1kbWUobH1pRyvGfNcXQWkubRyW7xK1s
aQDwudHra6mDKkiwmZZWPBLWFUCggGkJvmF0QvZUAhjSc2cXSBNDvmaZDEG3cPmw
Hj8VkGNvXfBBUg5R3on2bMrdAOUp/SwXV9/LAZTXcpnN6I20yHIk7s8YW7k4kL1O
LcXmSK70sv8qL+f26knqDOPuksICQpA9ISudJj5/r//zn2Key/uPQ/WtlLgqDMAP
ztmjsPWHB4BdEKwinuN7A8/prp6VpljH5jbWctb16511ANrZ8iHwSJ+yCBkiEHHX
46zzT0tyJ02KnlS7EMr2uGaEFufVQLfY75xtKnsjpn2viqbHQN0LUA/hVO3ukgSp
FF64um+qtsfmax/c/Wpvjg==
`protect END_PROTECTED
