`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8fZmJc031Rv/+wh2gob3/45Ya7+WtSB517uWL0wq+IbtZXwJGa0cqtQfFf0ZdbJ5
J2KBkIsYO5nswVnLi6PycHHnIPipeLs0b0hPTfby0jE4Ps0l+SOzPDRdj60MYFsY
8/4JuK01roRhLlAxiQdlsA+1nBRMvbat8tk5C5FCToPd9vI/azmfoBBK5AF0qLd4
fJ4eGU4UatDqZxbQ/uP3wKGwEh/Dbzxoci0x32noUIZIeVCUcnBv+QFF95zLi4vL
CkKtqQNQwEw7G+QFW7woRf16iqSO4Hr7Ok3ZB1HQ0A6Jj/UPYH4Q0LsyhgHqOQrE
g402UrOAZ7uPdkIWeZcNGNFiA+3Vd4hogIoDTSFVaH6pT8ktH3NyE52SWd5zjt2U
CRss8A18SB5jfMOGLBgrk53y81nVRBivJEN6Kr5FMLxV2q5KQ4NAIDJWAeqPGKr1
BnJLajOCEssJbg6KF/PcLWBiAgd4QLkgu17/ZLC+e5expt0BNUEkV/ZpM6z4QUcH
GD9ccaIqEdaFIOqPnKjH8esp9deb1TnRMpx8f6YPidyme2MnaNdZWSFGc4gWQelj
MJJC3+sBy0LYKIg83ibijA==
`protect END_PROTECTED
