`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
90IfC4RdyO9Qw/RWHxHFqI9v3dY5F1ES+vxc0t76SrNNwQ6wCDp5PYLXlzQXB+p5
//uDiX/QgXR/Mx1+7499xoAuFPFvflxGBj9BQNEenRqS4Me6ACZXZqmcfjEhPZC5
aneoPbvqXHaqaJu66QO91E7B3Fd6RHVeFgH7sSCJegjXwjMR3VGO5DbfRWFU3w36
v0U+XtdExIY3xGsd6CbEUD7IMMzVytz2m6/IaNenp0vxLE3LKG6C9BeKcvPK7PhT
UuSfYYUqgviAoof4JyAP8gjzcd8JyYDy9vP8b0GyTN4R61SIuGRMe0do8eikbr+D
FUNkDSpOycT0E+zvIJD4h3kdAXuhSaSkml/XNYVM/CjA9M9oWDB0GA3TdEysMTHz
JKa9YDzBk34VT3vHuG5UbHO2AvYg+mmnaEwPtv4Gk6OAcEMRi33BFd+ve/CeuPzR
PuI9bjagS/raC1ejGU0/UH1O/XpVpvN2yaiAGZtx/Z9FXM4I20G1JsLzhCUTxfFN
fTu2Gf/4411pbBEt7atU5fZvyWHI3fQeNtvIC74S6CDePzHMhgGAqOvmhHm55fKT
GPR5Rs3SbE+XYv1F4p9YOfxK4RYLoiL9Ba3v2NjZejF4GVsmWdbNmyr0FXbzEwMl
DdvFXgaQIkJ3G+owtIFOWhIB6igEgwyNla7zkZTnD3x2P/0odTq0e8QqZ0O40FTk
ODl2Gdno/3Qr7o3JEbnhmonpKsC3nY2UgahmUodQkFY1R0nAKtC1UcRP88AeZ/v8
onVTWEQU3+CjLrr+j/yupUqXdqiiDAdmAsJosxopFq8DDknufptB1oM4WkKRa9Nh
n8UK0LiIWMPrDwaMaEqY+VMWz9p8/IzvaU7sJZpWlZ3TrRK0A4WcRaD7ccFnzDKp
7ShAjtOBNdCmF9z4okNYTJ/JRBrZjfWLKyzuGmOO3N7lDzYPOjJOsSopHNbMvQSl
fwAiPr15vPzSiCs5XItD1YX0Dtehm6qXqLcdCkT5La1aVu7xlwXoUnHPPIbzu8oy
J4dpsEZjkE4De6bj3TMLxuKDc2y4o90DstB5gRRq6Kb+dJtdXjfgBrev+Lx9LIhN
xunDLn8QqTXAxepFJpZIjvIF8EG/db59gtrzGEUBcPrObpetCHOMhWR1tC0OmDjV
bryT69cZsbMzuw2tplkMuOtK9GNQSh+hK84O2Vs6Q18WCbzvqxEi93GmJpvRu52u
35kVAbKJr22fGVCOegPeqrpWh8Lw9rAiUMvg3skPKKMD3sExEyKMQiwzy48Cl4Xw
z7oOQ8R3f4Cmz44ePiec+zaaeInqx6k4j6N39UhqnaHBU2M6hL3u6/qBty0eGVqo
8q292aeUDPkvRVDaMhbuENJYwTSgJaxk17t7n9cx0GZj2wroiJ9aHOb0bb2UzVuw
RfTf3KSXP/SrPE9+Ov2heg==
`protect END_PROTECTED
