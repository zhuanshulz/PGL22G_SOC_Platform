`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ms6n+bNH9YL6GDRf+A00z3sjxBCxCwlmxDBo+In73GxN4Q4b3Kk+/OVUf8mTeil+
tYUbvBD+g0m+fuZZ5AwgEPROc9ugN8pQO7R1GMQt4f+eCe/LMHmWcxBBE871l5Nl
bWsFGqISsej3Rb/tlEqkufQ2DKgT11H7dhcd/Isn6cYt4+Kzgxsp4SFCGsqKDKbM
PI3Q84bSy9d2r6GOtDR3YhU0SYuSyywuAPazwT/64ZrzVTg9QgCHZjw+flug3qra
GHeQQUYw+Y11S6K7QP9BjICRjLeZZNOxcNmXVruJIcqtzzdkK/fnZYHYcaSyfvNt
fV8822FOCMPN8UVjNwFxa90VViEjAs8bLDzss7nemnvssQdnTqfTHxkJgOYGDU1z
3r3hTv6BD9ljkGCattIlg0PepzocdN44S2W9IvpqUzJXy0wbBwwbSJZSU25DYEKM
oRQu+yTLbvMuxvBBSqP+4quKhfmekJ1ZszuyA1mkGTsH+6cUr0VR/43LPZuV3q4Y
6k9TkQAVOYbzurh9PbEBIuLAqVPmsORWWMdTOwQCGnjLJ7HhREUnTL79silcsQHu
8hxiAGmYRfS9Z9t/fHlFYd4pg1uPzHKv7+inLguCXqj2OLY6//dGZMmTcmOXiBhv
d6mSKAhvP+4XerE+7ZcjiciGuBkCNcOL6COfLlP8NgD07NAqzfrqc10HVoxk/xP2
t/Y3xPhCqX4cRyGFK4FA76f7M37EiCg9oQq0wbHQaFFcsoSnBsVdQcekCD+hnxeK
mINoZJ+fU6qwbm7DMcgClLEAMdOgRuudmlIoI3KTt6OC/F8DsFq2ZwUq5VXcBTAi
3mFng+ox474l+pxNsxBqSkJAigmr/fLBqrCVA22HIpSegLgYhRj+tOZCvF4KfHz2
5oQ0jJYLZwwBdDDKm02xCGKTkmYpeZ8NgLxNgGixGvL3sF0tFAYNgXv8qHl8syzY
8RiPv1WyUyukO2oqTpPmPFWztuuMGqTiw9sp4QLVWJrAiHVC9qFuJ04L8o87tdAS
vyB+vxaHszBuYmLdd4CZ8VkyXwpbU8xOMLDTV+FE4CQdIPSpYLaupVFZeh3IoVHe
/t1Gj5l8NTg5ZefMFvNuy4WOFEqNLlBTNYm5ExdtzOMc2F4RqoJKba0EWazoYxRC
iLRr7+6299REaEg+vtM1QEDx+CA4dRfyiwlhbnvQzsqB3IBRdo968XUmlyuxIpb8
KhXrklA0Havjxclqk9s09bjytjU3URbKf97a6/PyAL87bo/TaN/OlEzh3utaGd17
CQjlPfEpNYtnmmm5Pg9S9RE4FC4EQ0m6btMKRXcEXAOCHHAdZsBfp02ADlb1QcCE
PNegmOEqShsIwOqXUVICX0XwhCYscDa5+9/85KiXroFFQ4CNDVmlLLbpawTHOQw7
6i9c93yJqUh48DAfLfwWjJbbLeT44RezhsZgf7m35SMlrJfhLrUL2JlrnFJRacAG
uv/a+52KJxisdIX4ykSpGJpiEbGnsGfOoc6nNzMTd4WgQV/iBqMRBHgAald31n4G
aNGUltYNwV6TAS5x3QB5dUiBGfRm+6auV8LE9ZP3g6JXCXmoa1sTLT55dEnQTjXM
98misMkBTLOJbDZysu2+xfGxybqTrpjzLh1TpgCRMdzy1csd5E9W42+zqxvuR5JA
BI+uryYEMa11r3x6kuPLN+L1Dtoyvx2neLnylyBVX332uZBVb4MgWSyjVOQCgIoJ
/G/AR47VKG2ZDJamHcpF4c8UB1D+7jTaUfX89Fea7mCIjMROvYBpZHKEW9F+sLLP
9P70YvhBtFm8p399CfpwuCM38vc3l/jDuNGM0MKG/2OAk+Donq7DtzOc/Qlq3SZh
pqUe33dGLdeOK3IJrm9e78GA0CIfOYGspxDMb/ucJ/ORHrcpGhZAW9WSNHJj9ymy
ZhqsICTG6vXZv5GLbvbbPKvUusbLKdCct6bf6xr1oY9bW08qlVgbMdg98yq9zRYZ
udmLuVLf5vEh1Vqc+Y24VfgOMTaJ1khp5sbOd9xV/+qBP+mpt6DJm/pR+UKt6Sae
`protect END_PROTECTED
