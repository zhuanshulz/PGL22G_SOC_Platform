`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rsQiEHNYKcIiC5vJqH+s+2GE201PMxO8jYJQMcIbKFYvFoZdLxYmucLRaGZ7TQyY
35YKSWv99h+e5g9/xxg5FkzdiCLk8cpSw3pNALEec0bm43/c0Bcq/T4xo4XRCBxd
cq7327IB9KCAxShPEmkSN4yKMf9tyFP6K1zmNZRH1F0LayjdVHkYXk9c7Bx44Q4a
Tv7hb7pczxydwcr77MeFcz0MQ/BDWIK49eES/dGZYitxItQpsDjNovcwR3apnzl1
cNBPFHPbHIi0YqkurHfMR/Tat3aSQreDMgol6zktPERuxQPMhCycCyx5GJsWKHOX
S250go5YNCFSNE7yCxi+dD0yoXSGOvhHEv+AIgxyWcuKqY+0RiVOGi85/l5QeVeW
UcSqeq6Mes6F+XXlaTLO3PQkGU47gfkSJRGnhpYdr6kEe7aaRxPcc5IkBgqj9Hp1
cqz+c5xU6FY9pA2MDBZtRaOl5gri7Ruc38u4lsKuDU8VjbrXvfwUPjsczj4gP39z
QALI23YJDc3ItjHtUa/esx+8sJfKlGQnG+NDpVC1nidgi2BKch26AZL1+6FurCaA
m0bmOoM21kF+DGsbY61SiddpGY6xJEu16POIK1T7N1mg1sFmxzvfk/ztnAz2zNoO
juV4YjBkCHIZS2DngvW3/bZHcHl0eOBEXcQRDOFPwUhQE+648X02QgflhoPV7tfR
+EBsGOw8boiu5TqwiQtAbw50SCYWWELtSoYzFwNib2UhvXbg4Wcos89Ro8dyBKEN
UAMO40PgPFivtWgYWwA7gzAMHWEyhuxFp865EC4ZV09ntYwdpSLBUs2hR9tQ/hqy
T9WFTDRTn7pleDVdGa0NxVGe+MbFAbCQyrkOKUuNtH55+PD7MUvXU+h5gdmgDjRY
judSb+XqEndzIVKLKuiEEVAD75xDozcQx2dXpTrqR2dQGgxwm5EeX5iYj+M0XqV+
8MZvIlWL4pKIZDliLHhbZaVGHmFO6F1zNcgSGYJAHq3jopWSVHv9XPRICt7K3rN6
`protect END_PROTECTED
