`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9A+xiQscvjN/TgMzaaSPawpKvwYk3NcDxArFW10fSKoICVdQGCSFrpg9+k/tZjfE
aags66a65ZNkhoMCSZJ811cDzdQXRDlopTwcTnV1QpPptOTvpq9ey8wMsBpPFYZw
76+kQ3WL0fjRPhA3I3O7rcgPDHN4kWeKaVcfCrBrfjLSLg5exENZojA52V606RuB
+k3v64DMK9XhWeKe75/yNkB7/U2r126Yi0PXucAa/E+R+vFtp++HDNFD97gktxEb
zOvMKAFtik+h2NJxznvJQoJyOmqVu76MF5kF076/QKVKbY5wnSUColMwWgH/owZQ
wDDbaN2qs3B2Sv9YrCgXcAY2c8JY8NJ80Be7WDs3EnyzNr53plMFv4yfr8LjcDI9
SVfyFfhC5l5c2nYzo1XdXfAuESKwbC/pbgGDndXVHkn1gomOGKDof8WpI8lgolrv
7iRQNDEBxtVhHztydHdJluv14Erei/lRdby3WLgnUqhMatk6LPSN6yLfbfM4RUH+
r3i3u6lZYBenkOwsdAc0uWiK8WwcgXFcXtsyg+YxnhK1TcKDFCRmqc6EsIxQiDQf
W3Fmhg4DKK4EUvKOme6PdvS8uMbx4O4LAOZjMx6otB+OtPRzzfx67FZnqXv23MZG
JS1TX4VBW5yA5V0O2/wss6t0ROkSkP00SNCdY73lGTc6Eu2Xox6WPCelx2luNibt
FVD5w3i0iiKI/RKDCsye2fTx4KWMsaAXin8DPPYivsNPKJpyX5SXFXINXvZwCCRZ
8v8tI46pnr0PjCTQKeEhGNzGVZAlqQo2hezRNUA6oa/o+O3sOqHxXZjzHkm5qoix
ndCGoQdUiVbgyd18nB0SovZNdZvB2HoScccMy5uhk43ZsCaf4iuS2IJS6i3xV+9J
U6n3wo2CX0CkY3Eo0pFJiO7PqAxBBfaeeOq3BhT+9dv0iqfOq+Bp9VJ+Amo2lC9D
Q+qXHxjP3tFFcdusSETyjg7AJmjp/4KRILGGy+cB59pT/54vVgGRXUjwgkxbJrVz
NvvoEzJmy16kj0sNjAjl7FWJiCUec+xupFMt3huIeEOBz55DjRvjyw52ldgHEjQ1
MvdCl7eHFrbqRTOozrP3hk7FgQHIat37p7m2kqmK6RNVmQexwXXZ6dlYK+kWBtAk
uLVKrUYVi/sfu76tNOZLWZFNC/dzg/Nn4QsKlbcPO4e2489n9ChaLXPfPZLF5VQC
gwYXYczy04W7GXmIIX+hd/iEqET/NDyibh0xHfxkRedBiARWA3tLXpGMqghb3l9y
izFmEx1fDX7Dw/7ZUDPfTtY5WpXPuF3CTQv7n7dVE3mLIDLL8ncTtSyo4G2hYrom
7RZIsOeleIcOigz0fkRUXKI3Pu5nWqTK/28nYSGfJlwSHj1qWd5Pn4WlHwWzF0Hh
y/+gEIjybOU2xx+19vIaMavhf77SOPnPmGYEH8iuC0543Mu7HtOOQ5RGhtPdV/nl
QzQld8QEuNSYNzLw5/pRIKRSICEmS8DaSDpYscijlRDERIxdf+wqqzD6UilVWgCx
wU/0aso0K33fIMTyLmyBqaM1C/oFqom2KgkpLaQd+VZKIgAiGJM88IrFyqDOuZXH
hCxIyUXG2Wz1PIUs5jaGYXDHzJWhjhx4743kK+G199Hyk2qE9RfUjWxRXhzt+89o
C0ibIv2RgpXiHmuL3oTxc4vEeI1U9oGDeqdOft7SAZv1Z4fKwgYmt4ikiOE4qag5
0sP2X3gtOL+rHXHu5aT0x2ms6hRdKLhL6u/gCib/nkfPRQe+LeHWBi2B/tapuez8
t83iT384W8p3HAkcNIcJs4ylMLWECNbcjA/OYNGRRnjfhekBXK+zwYNDAnXm8WFJ
w6yVqTOu1nFLiTV9AuA/yxr+SAogvN0zop0j5nm4/FUDDmBuUKPa04d3ZFRYJ7y0
Lui/T/9NymWpLLRfavl1NA==
`protect END_PROTECTED
