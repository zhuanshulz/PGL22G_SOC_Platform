`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ywqfi5UT+L8GbPu3b/yZPlvCq8Pec1DMXm+N/d6xibg3ymdejYx/Aqts2j//pdC+
jKJ4cG5JLx/OwCAQksB927C0RKPT/14qa6A8LcQTCVOGd2Qlb/UnJ7OaumwwhR91
HarVqp8qhAZ4oW58sHHNn1Ihh96D4TvZL26/SCmMCvfC5LEjzoVg/kjNv5EznmjD
dLm1gNncCk5hy43IpcLHkecIb8POGStc3Zqb83tDHtW2/QSy4yuK6HW5WU1N96UZ
45YjiG+Y8W9+sKz2P5xx8PR8+tbCcIFOumqyZeJ2UFoNh2kMZeKOGfUfnS/OGZ6C
jJUte5CSf3qNNXTK1wA+z6i5Ks7zDUJluYAWRnEy+UiaK9j/h3pcTetyPXHxJepC
XYorgfLLAzf1cAYg24/XoY7auTO01miN4pZQ7kB81dzPdd1RpbjAHkCgzOxpdvD1
sNFldj1uc3og5AX4+yBqO2x8RxBFr/Y+qdSU0p2lG3eJM4EyPpL6g9vy0TrNxIP/
IQGm8mdrk6iZsMIR9P106jdCqOkvup6a9+zBHmTXrZhV2oyExJyljGh094m6UjES
K8gqYCdBZP0plMt/AxrP9mWIo70zmXCUuj9bkRdcZtKOlRK4M4dabJogbTt9igGS
SyyVB1UufyvynA6pSYcdjNbyoKhrwR63dcUJyJuAnIK3Ut0EupaeqERWOS7fHBW1
rxGU2L75QUkwpXE/5EREDx4pzq+OoTsLXVR7QFOvmepmLWJYuSj/i/L+T474n6Xq
ckw7Xio7YOJcc2bIelUQ9HOIrRfw/ooNSswkSJloWnAtdCzpF1HFppNdwHXyBK7q
P7yih6rNbufHoE+T0vfO4Gj0p1G8BWWhQBacJC6tG1gKYCxw3lowxBr5G79ON91X
l7KehTNoFzUhMcQiyLDg62wHJWaOOzTHaiqHVdMA5PeGENla0xAZRIZT3oVPRLXi
AAhUIsJvtd5A6SD/jKiTfzz+SSDuydHIuc0QqmatwDcTICvOx7yu1watBYAEN5pf
UNMLCJCj9HHXHuEwVOoOtbCfNkIEP3MzBaB/XHcWD9xEPqnz1HCVXV56EvvDEPmH
koMLUgJBFhzBrmFIrNS9RBZnoHcp7gOvxk+Ujs5aAb1Hp5yCn/qMEjT0Tyn/IAMa
u00RYlFufU6qRaKYUPtUR/7xwGz4TdU2pocSpZHRdHPr8VrHSh+u1mge1RaOU772
2cdLW5i31j+rULjEVsAaCCNa1vqx+k+mrzSBt5ktgqThNUjDWnLtjGl+AR6l/4Sz
heVEl1BLyBK2PVizsbOEHaHYq0wyb+5jj9s6JP4yPxD2+w5a2hqSKcOQoBlss5nh
e4k382kxwVAOUj0j7mih3pZYk5V7B1M89PwilW2uq3sDwE2cVv/6su7WYwojBCzE
/K9ExAp+S4IrrYwIyHlEssKGiPKVVRKIyG72bkkQJEN0tYuWtHTN6JoxtSYT/zFW
bLnyNXkM2AWy2Y7fQdHZk7LDTs9Ytj4lVS1qcVsEEacg9S/lMO9wu/s7582l/jnA
z1EOZLvA8kFupmIhV1QT/JSw3Pxjiwi6cwx5vsK7W3AKY2MVEK7mCd2AlD3W9dWQ
lu6yl9kHhSyyrIxAT9oPHhcBXcUEIgf/iaAf5Z2sSjzZ8c02X0OY8HRLGLdSmBn8
PyiyWpXIO0qIq7paNABfwZ1DUGJweolwFqUxFQikS5xs/iH/DabragyrHCL5u3f7
oSw70TKK9IY6+mGt+iVcS0u5EFcCphuNwYgOHGGBnP+M9/1dkYD2hGPfvNpS/977
0Sjgq9WMReNFtELYM6NxYX0K/oaTWwJk/KIPvlyEKPajZtbdmTFnUSxn3qqVq5iR
XvFkAdPRAdDL5tv2rjwgTrkDnV3xGXzuTjaxM/KjxEki0AV87sCoPHs7ZUqY7pZv
Wwzy27LdkwsUb+JuQU6ymaSy6+d8TkYlo2Uco0vBbfVENe5ywOV9JpbIL8d4Bz6d
dnJ8VV4wpa2AQysvRfje7jUwzffV6hoInIcFCix0F/2aOGPPjJ0QPY7sOkWfTcjl
HcNXn6LeAoIEftYBf83vE/YgJtFFmkIimpaeDFy4HSAreEFZASoS09b+mV28clvH
iUsj3lV2ptafVlKID4soEWFJSRbg20o1Grqo923u5wTsgAtKzMhv3JOMY7545Qdf
VNXB0apRA/tZEJXN1uWAFB632PKR6eWihuk3icMEc2u+H+ETEoQa14S2ZJ2Nxuwu
sc2PNkgYDcSG0Lx4PzCdb2363Wyt3UHFE68oOHmpL6WrWw/gzuRyENa6xQeM8+Rj
77zGFX6vLIieVrFtEaNgMZ4mMBA+TdUPDLGoAnJkvwNEsNLQaK511tAdKqA4jJkd
aTtD7QrjYIidFZqKAvtdia/YPGTZpYjBEPHnpcTVqESIDMCYhX8wlv/MOri0D7nH
cNX90IHwmFzYyieSwX9Y6+cBPyGG5wPm2Cr0vhqtbdvh2LcdUI0N74fkhdcx8t1M
hnFM4fHkfd1BrzgoCDEBH6uUuXOi8xm2JHmiubF3LYEdSePHuzE2qnRhk1HPtwQY
FDo7sVJgepxT5yy1lJylQqceHcVB1zUWZ/5NWc/qR3HdzlcggQYAdjuUZKOrHe31
El58mbm9qykdy+SlF8KGK/7YWkpyuv5zRG4AmCgX8sCEsO/c06BUdtBnOYzyQxMl
5iQQT6Fi6QVsVmR5p3mrYUmT81lHDpULgYCGXt7uVlFIhv96ntGI4p8uEZynSAgr
RuQbywlXTQQQwk+lCG0up09f0Ctjz3rNMcGbs4bYKh3sgo8tsGeCLPtYncApg/bX
pgbKU4ZSb6Rx5CybGp2ERH1tAneE6jVz4IafVHXmlqPJScOyqbQhNUJ2A9j0ZMDL
nybfmhCtUjMgSa5T9rsNdENKMe36faKg4uIN2+Xr9VkaiPhWb0EWzl5Kjew2cS+O
g314NgxhpTTPTOv3xpUO3Ee62sFU+NodMKO2+MXcJArmO7k7oIUfvbm7H+bgbDyS
zMKt66yBqorTXGj0Crym0CgE4yzkUt3ZVmovzJT3d+krVs71PyzX/Iw6VzINuxC0
XQD43belhaM3akO3BP05/YsZMZ1A5TyT33SL+hZfdLHcF+GCNFT9KGvTi2WrYTvR
w/CTh+oGlnzCsqTkw752hjTPcsZxhhmo40egiQoo4J0SrBhuiEsfXf3kahLnJjTm
/zwjB7rP3kn1KtzsGMzEr1gu3ItTVuZ2ZegXuwxLoU2Q6IpL967tJ6CNalD4R5KT
W+PQX81cLNQGIVU82R2Ol1aYTYfSvG+EvyNJ91XHPG+IyW3JDpbZpFLmd5lvtSGV
QvTC2q6Kv7mYLjqUXbRjVhAjhughFLCFLafyrLDiGNViNM+KKPrKPKLp/2W/fKim
Hb9owMIXwAnebmlVvYh4h/y+CJ+senM0/hLFsZkFiXBGuOqeBrAaZyAl1UELHOvP
6wV9aon+OGSbxRIGTRVvm84KELfR8IAyXuay/hAQR9dMNkEu+8bgvUxMGGdUvrmK
Ip4dHer1539hDIVbgPzl5fFZirtLTBLS+c+GvBPneE5IIyE35xwpWLGb0w0S/kJi
Gkp4/+yyb0FPnhA7nbYvxwGiUtPwY9BTl/A/sGjIcFeZFtyTP/ONTNuXkgl3xtFh
b/GmHPo0yHOs/KgHiziZACkXqgMMdtnl7JSCE0K9nZtpMioAG8ywYbKZuv5EuT6g
XINfGfn9OQd/8SML5ZQjEchCqlPX7n4TAEQ4zKlhKd1xEaDLeEXgJQPn+7CCKs0j
L8ND+TAFto2EuzHNXZ54CSX6nARwrda5AYxD4IbHRTdD5fLxsdDdyC0we6lWWQKf
+Mvk8Zj5JoB2EwyLWAS7MLtdv0B5EWk41woxLJ4U0+f0SQqP60j36p7wjjRgGBR9
gWxyyXYS4z+dm9zRWvhHjCqg4f9Y2lzMUFHCRzdmt3VYNBqeuZrX+26KVwwNzQPU
mqYvZL4u20Zef6DcR7mDjsVErbxwGyjwWckkyidaA3wxiqiGpBsAe0m0frojvR9l
XIYAdaAXmaAezlfzrGgUIwfzMSNOAdQ99VPthASzfQIxbBlQzB2aOSJDID+vxX0Y
ddnnXC8VB3hOrdLOovMmqNjySg3hQP77RUFRH/0YsHIinYfFgXObcGpehLW6GvUy
ATAIPNQcQmp2EVcpYydOvmfRNnY30TqHNMTxK5d+QveXQzI3FWnxy7BNOCu33r2O
Z1nwpLu0ntkG1+FM3n8hTVnBLMETNy/uKnd8HfKHCpHoFuF/X0MPVT/IGed/ZXhs
vHFzaDtX9qUu+3FVgNMoYcs5V4UIARq9O5SR4Pt0tQye+J34eH7qGmosgLLOJETD
nn2P5fqXenbS5BPIsJqnx0WO57mvggxlFUg9coK4iF6t0BzOOC82KBQlLGaGfNNq
6BN9EckTDWjIhNNK6p/Qko8xoPLnz6sBgYBbCxKizrUYNSIOR854cSC9Cwg1sk/4
6tRTK+pNWJSrv9Jp2uqW6ZtZt4e1AswI58ryimYqBBJ8EBkSzCjIZgurAwekWWVl
scU8xh2cG0sIefgG4Bsb0pHoQOx2/GpfsK1C0JA3jzMj/o6/B4D+WU9Ahlr9foiJ
4cLinSDm5s2yA5qfxWaOQhdzc4QwDyGpqXfNrW5xrt1ven4+4/xKMXa6jA74BtGL
SQaJ4qpVCDcPBs/m4qW5WhcFD9NtQZpuengHfgmUO4L2YaO5JFybHvvzkZikjav/
x3fSYl+PwGCJUO3PyUaT7kExZYYSp0s6Sea8TwexnvYHJP8DF3AFXIkl7O8A0nTu
2l3Ht9/yHJJ7+CO5QeJXncBAaaI2S75t3YVHGkBENlRt9hEo3V3RqH+ONxfeUe47
Yi8KtJJHpTsBviTpAD71jpXXAHUhe67YZ3hGFhof/zQrc/4Y8MjXHVNM2YjuTtPV
8wBs42L5na8+60VcyDcOJFxKOLdyO2kIejciJVwWB9Uo0VjKI7luaJbc2taXRLdg
6J/s2Dt3C4pZn8yKohKt/kDUaYt6Jze2/kFR9ahljEWUlu+g/eYRw92QCtxo+94m
8im0CCnWS1kegVR29Vb8hgtGy6E5uktRv+HTQ3iwHVACZQC9YzTjsQTpbnN7Yuqu
tdlk5FrmFN7F0LGlteIJKTNfzXrrMQo4SVvRSKxH8PeIYMjBGVQuCBWF4bkC8wiF
ip7h1F/OrXM+CDhUQRlPKjZ2sx5+qKT7tXAelJoQv+Q4mtsdQFOP77Qw4a2YFja9
lFwdiMc5OAbBGKEG3vFVNCvet8cBKdxX6AwhosL0pYvP8gFs8PBJYOqZt2NUi/33
ltFD0G6/QXe3QmF7C4IfH/yBqsjp+RCm8MdAN8UZs7mShMwh0SieQ+ULTPAmpGub
euzM95SdsB1lm8/g3kWeyjNYR3RX+SJvG1sHxO9uLXabB+78e16T8XWMGC4l5QVB
P9ZgiB1BruU5XcDxKxIerzRRmpcBa3IS0qD5OOmwLi72c61gGh65UCS6ChmgpObx
/jrilx5OIh6HX4IZMGJpcyGN9HJgUwYKOd8mrKfmjFrM3SS+EqpB/2vJmql4PnW5
jRchN45SyMzJ03OhMMtPD8uUMjUvUU21OxdfhCtncaycp6JJ09vo30i59eCndfF0
PbAUQaaHblB1Hif5D2YYA1TLC8IK49zRgP+RHWicIsVi8ZWnvpAoHZY5KJ64xTle
yCQ9QliqZxVjkwLpef1F3GZvz8ZIm7TiuLespSyJS/I1ZGuQyjFiHrL8ndIhfLWh
96WMqyODyRGfGHb/6xdvMkiJNvpdN8ZePe4CYsew1aeFGCyY2Ho5DTJUqh78BHZ/
Z4sspQzqd5am6hdaS5iFl3QvzOI7nzAEYJfnQ0aXnxljPzV0yFrl8YSvWN77IeFD
hgDi7vCHE3Iz6EbybEFsrCg4PMTmzG/O5rXfTwuZAQ733h1K0nips9i/24BUo+K3
CCVTAWTTsFaRqWjWrpohRi7DUM/fCffipiBdtcFSdUGnsBtTfdeLY3RAqBNefu9m
N0IUfnjx0HNJaA33Eyw88tMzXALFikz8qxmBn3ibo9eJcReuoRsD0KzHGyjFrSrT
ztUl62hqYoM9fdDp97+uFFWRVwFXnOePrn39ghvtaIRN5k6kGVCDhpExTNs5iw9j
hohiaGQCsSQokgbdqC7VktfNOha/k6fj4MAsldOaW6gP32AmFWXQk6QbvNT72WHF
nHgapFDL9lKliMSiXWYbPbxH/NDdGe0aNqTz9NmpR82udCVRWXZPFN9kdmV5MkEg
6cvLEF+mhwVPB7IHIUa3dB1sR6c+j/MNTQml/EXxt+AxNb1tU57E+DrfHIwt815L
F9maCgeSYVtiteI3uVInyA3mZrcAq5JLNd1sgRyPbsqBuCYPvp0s12ci8d6wUZcm
FztJ4YUwoj9dkLTCS+7aZ/AMf13XsSrBRyPvvrjxqwyrtDaeEGGT1GuSzcJ+UDwr
91MwhXGGBQK4N7rtJFLgD/Tp0AysFvvJ6BetyzSVtvM0kYyqF5ftcFB8ageKfXPR
Fsat00lJWOFoadlLhxSfXFyyCSnmkcMd4Ac6/8bYq+hownUvHhuVYhKsJiUmBlkm
TZ93oINGTnh+jR9DolkR66p81J1JGg9qwTpB8BPEQ8V5O/kjBnns76NIvM1onoTn
7TgDtJC0R1OzvgZ4IpKRS5tzO/VtYhjQAMQr8S8uU3vKc2SesIpakts58M0y9X/r
hOaP8DtLriXAG21cM6i31Z69mveAypCGaRWrTmeII+OEFGj3eGK57U69Jtp894zg
lmb/awJvscxICLL0UM+0JwHrB0E1FxmvcFs7XBZoEDCiPK/R+CdK1FQMNYZX/mNE
+CRzDDLgDdkbCWs4Tn2i/5Qrbnjj+81tdMuwTisJlFQ2cyBagoLvUMXeajmkGvqi
5wI6KcvjM6PgvUq5olxdqescqGIs88cthmgn8aJa9VAIak7csxHH/6IYWpnRI+jc
Gq079TPUni9icqu53TE+BjFqOpaASiMmAGk0P36QW6cVyA5B8XHiyRFmAX1mplKC
1VBQY5110MjePtJrYvhXy8e9eYx3k9wUx0Be6mV4BRi2MbGtTuF63sNWycBjXWf/
E17kmpmhqf1f/NnQtyIHmk6v/5bM/x/JCmjWrVjobKJHKgEE/uUzS4y2b7hYf+n3
Mkj7tauImX/48eTtS9BTGKn0Cw0hjRQo7zWfIH/20N8=
`protect END_PROTECTED
