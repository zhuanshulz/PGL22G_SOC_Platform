`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wTMKHPZWOnyLA8Lki+YcycQF2PuDEMZFw1SvvHbkOaK7nHJcGfESzhXCt9Q43iV8
WbqoIF6lEo8K767o1pDrxiqKnLmwJxCR7O73TZ4/sRecZIGER6Qq5HN7t9s8otFz
QUmz9j1CIpv6DSJY2bEhlYPTlJAUIhegrtBvElWvN0Rkpueq6HiVQKhH7eUTmkWu
tDrXl+r5bHqvVnnTkWAez2TKlP4k+NqbpAOpqXOqIvZnWOf0OukqT5p+hTRf0c2C
TZhx4LHjAENb+xV1yxlz7Wf5zS0t0YDR0zVuLcL/XWYAVuRlWVhe2pRcT3M4N8bh
k8QXOAFWkJz9HZhpSI9kKRLL+pE1YFvsu/WtJ4bXeivq0w53rN0DZ6PU3FUdnedf
5+Y+K2CeiOPI7p3DiRUEaXew2zt9eGQlVbebq9uMS79cZkU0KOQKDOPU3mqe4A6a
pk3oGpwBpoQuY4jBFnqMJZfuBTVxWiiIXxz1ac0AqgLqbpznD6bgZfVU0nU0JCgu
5IibMecC9kRJG8QmAh16c6nsgspSE5o21ki6yWAt5D7xZt3DTy0uok7/scu5/7Bg
/vam5thFcfHG2xv2GTwp43mOsc9DUZZxB5C2hxUnV9WMkC66AsptaMyNczNKT/5J
VvmX80TrU87ZYXPdN0C4X5uRetj5lXr4L4nHvRmogcl9W8Qv3NEldK37cHr2Z9se
QlspGwP00bAqSRo9TwEHcwpBnpqUsVB957amTSrpD5EXtp0eA5M1rNlAa3K3FGEA
hr9efIirl+kZOyRIyJnArKzvJDXltQBR2GhvZLpIZBIe8hQy/UWalQyiuaFO3ScG
Atl/N1UJgQGtWIuD81U1y/hBgeYVo65WXK1aEFZOelK9pws5rSc5EBl1shobEQ7X
z5D1j8O2S8bxfzGoZR6Lfjr5YxsyyEM3UWj51VmsH9PuOc439qT3guS3pUxHnQEd
NpIMISOUHEOBEOsMRmsRz/99hSB3kzsKhd6zgvJ+NqA=
`protect END_PROTECTED
