`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fw+L2EpV7hre+XyRZvB+Cx6FAa2UDYQHkL5GuORePZGu5dKrw+YmEO4L0y1MjZ1j
nEZIi3fZrabwTarsUsImQJH//Qm0hhzJqNLtdUHAs9aN7vUG4UUSxx/sxviJ5PpS
97OrCNQ6C1cBFwnHSCLJoghxrhxxPEJANI3QmhiJjdyl1kEeG4XiNhWCCkrPiJ/C
aiBvtyJn80I9hBP31PYSRHiKXj7MZFraeIK92Ujmp6l9COVDikeYvmWCQdvgyGTT
TLL/WV6xP2rAZPzIBTH3p8V/4UCDMhlONYfgcfb8HPhJtU19Z/LP9zJTBU1D3ACA
jcHFraWNfHPkD8ZwWADrKFLkciPz46EB7Wf5Y+C14vIc+Ogbs+GmWbR2Xu6zhVcW
7jaGggiKGG7wMJY/EoA6tE8cx1Uar/NOPF3kYadu1jfedGGMebMXWQvfNxGBuBE5
sGFE6XD51JNEqapy/KvSOECrIWxrRFX3bIVKx6xL6s+IvRPgQ5u8JdUwJE867H/n
FCqX8/2D7yrSguviYJBUeq/24KPuk+Ql3qUQyTTfZHPqvFkdxcDo866PpyTmI+ZV
MhVtKjp/VsHumhWf+aUmODM9livz127v4FkEVC//1iDd44k1U5niZnZiOYgVaXIt
ZgNO69DJnVaeJdx9aPwy/TWK1q3TSHldzQCbNxagN/S5PeiYmE9o8KNeAGrTiON9
8qnF+STYd9Lh+KerZrUhSlLiRBiow1Yl9XnYhdBScHV3UvS64zpuRgUZc+k8kkeY
gWbqOTduc+9gvmvZsSdltQok8k6tZ/F9EHtJrU8t13DEX6TuzIotje6XKqqz9pcU
e5+9NFFNT210kTpdrAQkjEzUeX36cpToQyArJTneI3xKKdDCntWNupGUFT/cDjbD
VCWmkOhG9N/AB39bFKvENGlCjlwjUAgEv8bL8RPjvEo4wvv3M5jeR5V/H/1FZu6n
tz7HfTm0RgVIn4qtNjcQKR+/gzrL0vOtE+YmUfm4lwXzIcuSmU2BkNgP9y9bmhXR
s2TlRD3cxZJbUT9KzC4HzJ860wzjXV9RwFoFPE4TR8Ra4aZiXJWRzr43WBQzWO4q
`protect END_PROTECTED
