`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kZ6h/24QxBexiWYOSfdgH0j+isTGfDB86mdWyJSqR3ZTn+aIhgGe4p7H8ahwNiGC
suDnOZM2KKH1/KUFmwUMF10wIP/cYixyKHP2ZLmZcFSAVnKXxUdCblzNB+SKqlmK
zbG4u9FMxPMmzWnxzDv5EcS4KzfitFlj9prWE5O9R2D4OcsoE3ZVMPAvvcPg+G+4
vIOVLTLJ0Wz7sBEjRvP+KQy2Czei0HVMhfE2AcPmNxxa41NFgnjLmeUgp7JEj2Lt
wFHllf/zKHSIrFYl4s+Pv96tjAEB42QXe8Tm+76mtRstaDNwStyDueeH77PAtGhH
gpuNhN7AcxW/pm21HxAAGQ==
`protect END_PROTECTED
