`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jgPn6Zsg2229/zhWFKFfignuGdcm+BmmEEVi/wVJbeCGNiqI87Ci1XdAEvDm2RHP
hXM6Mh91QjCUr/QLB72aUWT5RIdXwa5SPfkGAYEVGp9UecNSvWJqlqGxnZilCTwj
e83BB43Tx9yGziEo2oqICuVB3WL0egETpRbfaVANUIlZC+qgBKl56MyG0ViPPl0o
WWPRKWlVfVS38K6pWptwj9MUWOHctIkhGSEsIm/8zvY52++5fFZ387jDjsQ6cbTz
saLLdZukFBvPih+Xynd8Pv/LLSQf7RMkoyfXAqW49+8NJqs1M5dmsFJs+0X5I0HQ
p3VDpX4WxdDxsmxCTq60Ftej4uo01Rd2Vdznlu1ukS/4x8A63vrmW60T+Z4CyKRh
Gu2bCalHRuqX+1gUyJl78rgdi6fdAYI8/rXcf1H2Vx0ahfOAZFZAnWzCV3nwO7qU
1kBb+tSXHnKzi8pkRBilEFxuEFNLH0PiEeIK3lsl3VTIycq4rdR1L1JqnUNa0uVN
cV2x7m79B+Ljjw1+oJpLvkOrl8T0aVdZxEdvaRnjY16Gw7QiN30r/raDczAL0Qdb
rKRohDfRI/84TNhkZ10UNMrVaev3KKzBBeRVBkeNm8KbLj8RDEf2FZ9HaOi2z3Yr
WkP56iqrnViXLdSpHhxZO9zhmdWukthhcLiruSGjP86/lCOBq8vGvLuBgu/8R8zi
bNPUao29hdX1cv+gsca94mwFJKKZT9ln+aoML9+CNz042iEABB7muUzd5pVj/uQW
a5aD/ES7Vvv3xIIkunh+3jzBOB7jbzZc+xPwpqkSXMY1opea/qW74FRMXubl84ME
6l5TE+wnX2Jnssdp8b/I90FP6uG3FGv00xuPjPx2plyQJZ8UlmIqOdb3Scn1Xy50
VJujwwg0D69D3gCgsawXIqtB5oRFq/rHK9CocOH0JaGgyTJcF/W4kmPYGWahnOxp
r/k8oCMkqdgH3zdahf4LUzO40SnQq/O2GCcaEdtNAdSFoVc1x4Fh6QrkXHDw5dQo
w9deOCK6QV3k0mt1Bd6VgwimqcfCNNxKhkE3Of8IgyYW885P5KPYGn1emxYWtD9v
5f2abbBPlcyO6eMLTs4gWGDcXG9gunsg9/iyhrMMfyrIxlDgVXNa4w848KI55Q7w
iL1d+4O2IvSig988lx0GNIltTSEKK5wRY+OKRrDan4aI9rHduco1Le9ZtFcGeZgM
GXrhXixJJ57leS4Qj9m7ywg2WNWqDzF6uISG2ivBnIYV5PCE2iNYcmMYGmWrmbI7
V+OhMhzXasP4zo4nU1srSBpwNr2iW3fcBBXWGOXerD3wc0gO0yA4L6Qp206Vtaci
oDmpATWSyLn+Fujc3z+PNGNxERrAwWqVRasmpjPEZH5aw6LLYZlp+fyNO2qe2fEM
teZmysp30qwzmmqVsocJFlMMhAvHW5KKUZOE4oGsrpym2nSsuqvnl5Axq7MvkHHa
SwUKmjnquV/TU0CTtymYzm9wa67IU8fYcD2wTkPPSimh8XmIQIlo1C17Br0AjrLU
ZpqKvoztfO9JpaqXnYBn26HFQNjQCcShDxY2354Ync45bm3Tn8EPBDIP8aeC2ztr
LUCK9WCbT5JocA6hLY7khCctSPdIFbEMUeLLbAV2GzL9qmi1ENB4YI5PP+bWLqk0
QWAtH2fLacWuIJUcSWS/F2Cyhudb+fS3VEYYXY6Vh1uATh1/Tpg61c3uGCYLZma9
hbyVlmYpHFXQpTZQBT9eS/rLO39XWmZ4+V8X+aLC+dOm9iC5/ca5blYDwM7MZDSr
w/9A12lFalM92D+IvRo4gLFg2I1z2Gr7kscG0fPTlIh7GH0nWCgBuQIoiyBKQXrm
DPj9U3RLBDIKIDke3CKfUMWzPzm+na0s+S9n6z92NKDxVhj8NkzBEIvTPwn3yzl9
Qj5kizLldMjhvondkXXJYfHnwXJyVJ0CNtmrYTK2kRZ/MLe++PGYwJ2c53RFLHPH
Vs61/Dc2RcraSjHRy8XdjUoQ5+LSLIGgPKXcXx3PZwIHCdR8nkUk46S0HfwhTp1U
aVmqbExUCTqf19JSxCmWt0t//p8pnCJXJBdoSQAoXFgdparjH0Z15tzvgv8c7Waw
uaIWSLjsRtCvTorUlwk2BCgYaF9DxVqlFiKhAEOUVjCNqM4khx8PTJhGTlgrKh9v
7FhMyD+Ux8eK73R8Pi7CYB2N++9N/O026vspbPt+2itiDaIt8NpFRmpF42mjjzcB
sjdgtDVbmXbHg3Zz6RyntWI6L1qknf5olduMmkiJsMO4FeJsvbjOReUMs1ds6wO3
M80LFO+QSoliRD9K9aK/dhNwO6hgUERx5Qo49NCUAJzqN3GYPwRavlne0OBt6mZY
3D7iH57kjr30j9oOL0wT7eJNuH/nRbafDBpRmOV7upBXSlmlBN4reTexYrYG5TbT
u1tRjhMzD0Oawx5g8ym3RtPLQgheEzne2NsdRYWmx92dZwezELkNdV/AYUUtHxOa
A5OQ2mdX2H9jD/RLF7kT3i1q8KoGETW1Z+fGgPLxKPQANUmI+NZVVya3NUfaVYvu
kB+2ZosPWQshbMg1hVP4YZDcwX5v9J2wbgDNipdDs9E4b7sjxE2vZqzgX5pk2fSS
1My1XYOJI+iDv/RMwUtNvT92LMwwVb1AibrxJv/6pBST/VJtPgse38m/7fPg9WpF
K7YP7jGi8ayv4Z0d1oLdHM4XVR9WfX+/7+XO4IqyPFavEm6mDCl7JNQjD5pZbJzu
wuMZUTEWjk3lZNLaW8aZpe20SGciORlpidUAEsszEwm2G/GvI9M4Dy+xW9pmVQOV
bHP6NS8tf3qngtMI4Hw164wChy5FZ9gwXa76k5TyLGGyMHXbxq1UiyS9A2Uu3gT7
O/D9x1KKcsmdZOxmGKCJtM39OxmqNxdr1qKjPrv2IriUWnigHae0IW3rAuuyenAc
/4qGcfYOtUgfb2BeGZnrUYoHB65OkkQ3WupdmRP1zvbcBpuLp+ED5dIQVterXtQO
PKo54CESjcZ4NxpmMRMuGJAUf/CVBYYS9AEB2jFt9h7FumVBJ95rr3lVKOWduDuE
dH4IoC6Q1iEkRNg0cCzg/5kAt3lHRt0LVy3zTnQ0MZKedPrpR/jsFz7XDenPs5AJ
qTxkesQ0ojHC+WunOCsi0Q/nx8WZiBCL2j3JGgN0HwSr5jvJ1K9lVcjPXaXCUZ2V
fxadrW1mZAUjwpnHMp61R0s4nc+9c62Wpl806d4J4+32J22Bxzu1mUghJQD+MwS8
YAQWDYWi8HYHidCa8d9TeSfDP7jTOm4f5cXgmEMM40FJUtTsP0er0oDbRqEpimGT
45Y8EUHWdaZwm3FtBoByTfqXmmjBnOpHYWyneizMRR667izVqREhUUNRghhpDwG6
Zilgeri6O51qcDfeKqC+mAbb5ep9V7UjxzbkXOZ+vb3DZRPP9THRtF91SYyjiYuY
1bE5cO/6aUZeho/DOX9CLTi3T4TLwxMjpyXXGf0rQuysDfiieuXTYphNe0GlerFE
+fNinELLU/ZZiTpAMJlihJ5NS4eHKpCXeVUEMBQScYfsAuZcABcf9iTqs8Gt2v8+
KfEs8q4Xo2EYJNtwL+yztW6k92ihQnap8AyQrDlFLiLp0uVpvhSDvvxsLgvePMjf
nKFtr+lCZXLj25RSAdtevkSdAezaZJcPmIWmjDCdJCcDUVEvHOD+mgVExgeZy5wr
WXYWhTvtnAby4FkgqHjK0Uivbg4a6H2U6a8ym6fS/75wbxs1xEb23HldMcRyqn7P
dXCb+jEKYXeGBY+aG7Nz3djweYCqJTu51eHygRHP0o6Uaz8x4j9k0A17soeS/5cB
nKCMIZ6QlwXfxuC8z3+B+MejXFwV46Jen0EwGi7MF8Jzz1G0WlzhgUyLtAJ1K7nS
bsBV5UjyVQqTEeLnK+nozWGUoWuKuVBrtdkmTcbGtJ2TZvW8NmQFVdqLltVxfZqQ
3K28IqZCH+VxzfDy4oA5rESpLsXax3ILI8MjzHmR9Q+TL74p+1DQQnUivqKCD7lK
/nA1vGkCkRneWT1C9GCl7SD43qRA+MUs46dJOs7+PyYBt0BHU7DjDa1DEi5xWYxQ
pRuwIT30eVaTbHLuO2z6TDH1wkA7Jl84uFfKijE6lTjQb7TyAMY+zvhjjNHlNRcJ
KoNJkF93XxbuxVFIyeM2dpzZpvB2EeSKS8SKrw590OMist0EKsJ+HVdmzPxTEkKO
KHeK7afLo9hU36xd5uWaFORbisGDXDdSeSOElrVDq86uXsOSe7/PtdQohlmebcDv
kSOSEi6a4YGnWG7BGUuaistWWG57aCi67N26NWOCtYCCaiRurHA+lVBdyfrsERCp
IVKLFZCsWFixpa6wIkqVJ+enYoOu7DDLfH3PoIJ4r5VwWpzMaXw6NdV8UVEXep2w
3wd7kGCmsvZQ2MkY9Kv/DeQfOyQCeb4ScxZ0odIN17YzrFIpMkYE+ctARAKScF0u
AMSdqlsGvLkEiVqKTY6lqewadglJJCISNK2cyW5mhXuNNsnYl+WSwINcfKdOt1y0
EL8d7KVRJMkB2Ob6xZWFd7d8AY5G7mIDebZ7gwNLZ5LHdh2YldkkejhE1iM7QwHZ
+8vwqMwTlXalfzZKqkAssSQNUgN+Sei2zBjyLvqOBQO9KD/rdPQzWuUkRTqIjUhk
MmJejZNCodaEJy+sUiPOQgBkUhMsuNvZ6bSc0BBd4kCFcXLJzmF5Zr1p9hwZSlSk
FhhWYQ/brT3jVKAR2hRxYuh1cSadgY+2ATw2xl0UTnXjFN0pHv5KHfW22KgkOTAm
JhMfjvrjNYPkZzKB7TKrxmzjdFlMhuRR+nwpwSNMBvW5+p7PcXX2AtWYKQJrsIkx
ZYrRihWTGp1ZQmkfUh/QBJCRR9Mlaeho4XBHaFnE8dArxgx68zzvKNynD/atEL7w
FfpHne/91YiKZCNjhjsoCGvUgq0U+fyOjICY9PbggYsCeNa+0Yv1gqgh3OWhyr0h
qwgTU0l3nAxdZaqM7ok8hD5lR6n6QdHrg7BPheNifEdc46lVWc3K0VWtdByGWXMp
3kvfIwEt4ub4sfyNj9rALQ0YhfsHY/Gn7yuGklyRLvG7aymmam7XC3nJf3kk28Mq
B5gaVIRPZItx8OD9Bdy9jEjm54zOwrTQm8Y0n50gpee4XEbdXZEDZIkMk4BYy9Pj
geJpjm1cLW6nfnP5Rtw1Og==
`protect END_PROTECTED
