`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r8dT7VcxUKufeqLBzj3HBnrK8oytzePz7uKCFW0TwHMUmI0UgFjaJ/oBU9wfyBiD
E/kV26RDMOKA/uJWg5JOjd8xxm7LjXIoxEE7jAIapforlq+f4Yn6R+TMsnKWjsPX
wcezYiNg64exVE90wseDRW0Ze51M+4BfNqAd0Je180wg2SGQQR9lTSkM7GWNUCFg
Rmxt7tTJbML1QiPzvjR62vAbdAOcgEnhkv9FfCjfUuqmjyxoObWfNmltEJuPMG+G
aBLUoMubJLZWtI71vRll/o1jX4xdTfZy6ybfsDegwEuZss7Wt2ka9yNY6/Y2GmEC
2J3RwErjEWXlQaP2VgHtpkjOOLvjsDyYBgFhlcs7ccByfSrX4gOEX/KXNzd8DepJ
gtREQ2koWl41KdyNzzHBjiHwhnCv/hHm1+rKzEIEsQaIoP5HUMy+4mFNWuVzPh2v
LxOoyoMpMc5etFwxNvkCcPcuRgDJdCAj3HfK9Ii20xSMZJAwygGKokZG7u4NVt1E
dYSS0T4xf1J1Oa1XAzpCUSf+nX/M8LVrGwROXycRfkk21pOQvFxFCLjXai8JAm0A
DUUlmJSQhDgj36Tcq689rGPbH1DicP5IyClVfm3AVXoeFGzbJo2u+EhGdw+euifk
tNLib1DflFoBBACRFgfJHnuLxlL3idAXdROnIK6/lqwa4s8pI/Lvj3xzGYmEb1fr
trP8hVD+vfRBnk2byDj3YhW2j3w2Fk/RhJbMbthnWUdTt14S/RWwvAXd6ylFT1gf
Xslr4SfLDVHkoeK6vAK2kWFjpSIqciW46cFWuB6rBFUaozB6yrJcNTYTlOTMmnZ0
ul2n/L5DJvPezwZlWsKd0vlFnkQIZl4LTvzID+hylEt0+KcS6mMKiI45Ce2pMXnI
S58m7Btk2sEbOs8ej5ZeYIq7ybDCIK1S2K2Dd4MygyFtugL/vP1h/2MeVzrOqUG0
eGnZupMxaxmkdN1zSqBs394kwogdIk4y8zP1ob03n3dM+yJpXzD4LBvNnx3hypc7
M7BtDDUQ+bv99+lvag1Vql0a10Sgby4haTKUaFSENmaVWJxcVkGL/9okMRHgP6IF
TgaRC6ZFGENZJshTJpDlGM8VgP8GoHrF2NobFE2tyYygYofI3CIn90+UTcDWS0+N
eQaXYd03H96Bcy6DuukRQ0LOV6Saq5mqhIJ8rhy3UI/BOcfMCOhJoXFIKIE272p4
GSGvM+YcBJ1cRJoKmTKfE86y1w8IQE9AOf1YGqJuvBbCo2Y2r0u0lWgGVCg7Z+dO
KgqQUPpWJRwpgA+jeDCPyRsc3dqg/Z15mi0MoF2ssF4LiXnPkzD13sv64rQrYUMw
4fNRSIvAEG74RF4Q68B46DynB4GUcSvaX/tBK2G7MHSBPke/ysTuyDZ8dVS0LTQ6
PQYMZRLx0QyC5CsF5/6wrDxcKQcevw4VVlUW5XdCo7EyA6DOBMjfFkHOAo31VYgz
IZEycI8hX0/w+2xiq+sKlpSSLpScOyWhvQPSHqHfYTlav3d5SUA1PwxNS3GNwh+D
1w8lW4vqU49xXAv8LX52QRxRKZdbGlQ+yTEVaJc1QCDEUZGm18LHWPQW05z75r1d
+GhvMiZ0Mw0HkRmy5TMMmufR8sFyqujxuBGGwJpyk1xpJVWvvokgefSl8luwqtma
tDmjelhztN9fwx2QmxbhWST1GPqp4+sJAq+jV9PG52a98M8fsgRgYdFuqKMet7/d
dvdbzzYhU8fCI7fsyqS1exjjBhcrjF41b4uMmIPAew8AnlvH+h4UAprgknrMI7e4
N+4qnRPuqdS1d3kMilMhLWTuEkOw/jmjrV2qA+4kUmncr9kBEmw4RvcR7ZGwqV99
iMy7RI6E3IGEAmButf8gObMF80o/32BDvrR43seT66phKAsV+0XQlr5v/qmCBeaW
`protect END_PROTECTED
