`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uLcmFsAya/iT8EfRPR/51/2/Ptq6Abp73a/z5x/i5LO10Qmo+Qi6h7hWifpAbQyC
6/wT/CyYZBHMsTqzuY7OhcBD8FEY3eOo9i0TTKPKXjYxnzx3Jj829OOl8yh21gvS
xNDhXljcOPgG0f1jHfvtESp4su3tRVHYqVZmXQKdt3oo2U+v3JIVUcArE2ubFQoh
CXCc/r/OrWmvIJraXYiKmCln6AZ8WQu5DXkxarituS832IvsyLiNFaAk2/7snTAE
048QlYzeZBOx5mzVEUbH81Fl4XQKcQb6ecRdyu7f/lC9RR7DsP1lOA+6b0VC/xLT
oSWSAlsnjLteWkGfKvLm4fYNXgfqK5NV8dA4yLw7A2qJeTRTst54/c6gVB7EIgR0
SJ9TA+ei37J31evgtnA7DWJLA32yQt6GYi/U813kpFY0FuyhnsSSjqAAEnYeuL9I
zCUGbZRXIRO+Tv+SLNY4J2lV+XTqfWyDkeOWJJ2UcUf/ZBx/RwFpTGXW8/bodjIh
dJMIoia9wqyXY/2iJQ9IBP5bUZxbPWosgl4V6zlflMCaN7xYHyEPJK4hYG+75Vkm
BZb+g+/7gM+DpaMSC5xgrSr6GWDHjbxk32IcpTl36YmdyOhkhUESEvQiPlz4cCVU
oLPMvoXJ1hEotmPAmXUwclm6xKPJbxmHOoRyi30bG/9GMEIsctYk0HRjoW6SVcPC
kp4LN+5s1DFw5uiNGqj2Iyqb67mMUHMTimuVPa6iTNhXaJZmVC83ZH/gcPssfmNl
4U2RtrloIJQXtICBPeGCWK+wPvSsEHQssfwkhPuYfJw=
`protect END_PROTECTED
