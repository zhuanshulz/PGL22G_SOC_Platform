`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZQkzO/nR+otLtbxqHYdmMd63/gtMaypPHYqULHm5H1qPtSiwc813cHycMSnDW03U
KOnAkb0ka6Np/kUeyzFpTjB++uLnn5vDxN2UFBN+p93M5DZryGc+/Gg5HPNhSxId
ySZEqy6fgH870x3BgNyrcj+rSatqMxFeTOyk4vYCqSAArY+Ld8hGNXOpehMpWH1g
u944ma3zhInuGv2wqgAabbC3thg156E+RWknZVHLtmojeqB8lEcxnxLI09lxFLy4
JV6wMEix5djE5v/nt1lMiO+MNK3QusECWwyAy9g3JWAMZ/PuXpa8+1jF55JryL8j
54bR78W4wCNoEce20Q6beq26GjZvVjgNHyrsoNN2yQSZSps2wia/2RnFvtbkQo9w
oEte7LJPan9nO0iGHWci5SCvUzUJ8h7RX8pJP2qg3r9jkZffF0FTaXUChok/YiBv
o9PQvCfPxQk2aCvflJfDjtAdwaUeWsKeVowAP9AKO5vdydsF3d5BL4NfiMSd/LDq
IVpMfOhFUf3Fr9YlZLETIzbL4o69G/nvYCeGrcmySH5wBJoaSwVC9MzfjWNqEZyF
hrQghoP42YyEkdyLGMH/ob+xhQeaHnXJTrYgeE9CGi5chVcRUb/pjAhdDvt/jHuJ
g7zBh6qX7cu14Vl5Np1u8sJrvYbrvWQrGjJjP+296kdWY4HC4yqnsMYX1gWfsFkn
Cz1c8ddNpxUZsAw2nugU/ZmwDYEKO0tCx0z5nKCJ9Ma73KzLFCIdQTfEeKa+zV39
JtsMQkEpQTo1+stMVlQS3XCu+H8JLLOACsCXX7LEsevcW1AZ45jBWOJdswU0xt1/
o3N/D4O4OFWjnxR0NqxBdDud7BocPlo8vkQRyRhEKqLOR8uV7VIwKnjo8hgk2DCO
9feKJUY5BDCu5DgDV1++l3ddKXOXQYIolEipaD9GwDpT1w8E4Cd4NEfElRL4ygdj
uk84JcCkHKdJgcBZzQQbwF6NyjIY7oHNHMJ5Ecm9wX2LscEA5eFcvfDHez9gr8/M
C9s4aLdr0UI9RGvmJw9nYs2Ucigbx4h08/DVhRddlHeaQ+I2/aXfzhLgUED5BXVU
WP2KKl1FuTD0kZ1Q6bQ2Dg0gYrhZ0LJTL/tN0tPSqBdT9OuuYOSh8YabJGPcllvy
FFL0KpRW+dBATF20hPeC8zbb1MPY+QBEOEvNH6XESqVgDPm/N+JOMLiYhtp+wARo
H+2FQsax/3diMQkY/VxCprBGUxHdJ7uRCDqijme3w0Oe453s9vTdAq9XBYNn6oE7
xMzNGRwQP4Ftyi4XaP/UlGNpYwex6OLQ+29ql3V6zxUIcdw2K1p5etzxDdhv8e1I
+lwLoNoEnJO3FG3CnJGaPym4vNhuOOJWPJSUw7LrjUuxQF10h+nXHAXefxJBfIvz
jUhfZO1QNYNNqSG4LlV//npu2KVtBNHVEIsEgkcJrnnpXaO5uuhAt+9Co+tI6YUA
bHg5BfZQsuwQR4pagKUSUtbfX3PWFWMVIHsO370sO1h/7c6XRBbyRjDBUKSoDyYw
V6gl4nfElztHgR0lFy/P7Ts8BxriG04lqcwsfwD9YkrcKHUAaGEiIX4xsdB/97SO
Y7iUqGyg0CJ4OCUBOw6G1iMvNSMET33UX8Z3cUrMbPvGIb16Bck4dC9YY1Y7NUcs
PJrkT9cUYXkz5qdzR8FD6/OxNMmQ7rKwUZ8ZBBgEubFqmQpPHQwuLnNC3Dn3BzR1
10tmfIi0V5HchZv320OaUCcV8TkJNrl/XcbK0SxlHURLzkWl0I59VH5GJm0AHsaN
/jNeicxwuuK7S9g6h2wBA4wnYjxLuD8dm8rrnp9NDf29sznAJX5JRfLuu7hTMjXI
3mgyR9+hDR7JJSB943cCqFvNUMYuwpU17pUHs2bN5mM5CLvnuKyiYesGj55BR8EZ
6H2qnHnmHO9ZrGLYPCIBM+IWE/FgpYAcslDp3oWGjUUW/++hApISrLnwPWVC6NKY
XfMG9jgBIK1gKvUd+LBC524EdhyVkVz/MdVErHMEqPcIiMp4wqpGYhtW2Q9ct1fh
NKNZUSPC+pbqlkJhAq/mXViHOC0yuW1aDxLLrzmsKkM+hn3X38+chOEhZACDWgDK
bVDGWqcRQRSt8gdH87oDBKeLc0/wUrOZXrDz2llg6mlXo9iLDLmfIwKZvvleOO7E
Q/PAXQl3ROm97ybJ/FdaQKNEEJr4GsM8xB0gsitnczWhLbdFGNWg77q/v+UJxvWG
wtL9q40cxXxG+Xcew4cPwRUn97zHQ+g0OeVyC+vqXi/7dwbnhtR6aQv5zRmisYOh
3qurcyH72vXcYP98y1Oa/GJZoHcVhe8GDSoNxRs+toP0yfCpn8SluoFnF2dexqWH
1LrPaUWnndUrCtsAgjP/laPB63jgjjKlS1HOVdYO8DO3EGr7E9Fu+5TlV4iDc8eK
pFLmo6+cFIvgqJVCiLGWSJ/L2eXPJbcy5tGaes7ghiS3MTJ3GjSt7XwV6Zu4ap/N
VmSBOfTymmAKSXQhp28yS6c7SoGMWa7cqlRIGNnLHVKJTDei+g232ZjET764NzAT
TTcjzCwphRASM9cMld1vK4AK0XzNFw0cvBb/142TFCP9pirpP88qNG3jKSx3vFIC
7aBkf3AOELMrTS3VCmWdSZ51OssfTevrv8mb2eohGXU0kBla6aMR2W4LcMZWUU7G
4vGgS/gxt6DfagHZwXFRgKnuQTuFGjrroY1MXA0ZPKRw6T0HJ1cFBoTZz67Mk7hP
q0Ah9jbRFRtUs+kluaGccyD883SBzTigaMPvJgNgfI19BphCiBjjYrxOq0zYsrRf
pg6VAYsBD/EZ74Wbgt0KDKfdw5kztWkSh/AmqRCLPO3Gh0PeOM77pYtCLguHhZX8
T9PnZGJb+zmNzAeHjM7vD2PNkEU16aKRe/hRpGf4sFeYqs4zzVs3LRNcUBaYvb/s
teqxADDxGQ8AXUCBYzP2B1d0DO/dGM/X+igL/FsguDilM7WAIg2H+zfXNlj6VZLp
+VlMOgy6XTbIF3OucMdZ1NctivtWt17VmKeimT+oEkmlN2MWeVBFsQNQ7my/H8CB
TZMY5X7ZywyRBE3JWxl9Mq1Ju07lsOuImaRXTQ5iyY+wjiTNf9HevUBltCTTBbD1
3S7AwSA5ZDDGC4Gz11LrZ5JXHKSFISVqT1CYHjREoG+AGea+XxTJ9xlIsIvGG0TY
0F0YgoFME5XBImm39Ltcf27nDvX9eYt7SSxR5w3Bxfdyui5rZ/I+fg3AvNIdXcWW
bprnV2XM0/OO47CkYMRqJD56iQsaP/X+lFYaUsrTzkODwVCUhe5V1Gos3NG3eeoL
Y/juBzPR+39pEMDR4jc4dK1gPkzg1ufA3ovR2bnHy/YLvK9pnxT+JDSK8Z68cTOt
ob+DCAWgQMSXwJf54ow/B2fNSqi1h8IVoD55LCULikZaEH2rEii+P+XMkqZ1hREG
IrnQuPG/s25AQCfIDGpXxKQ0YU3yJUC69Kkqn5hgKUtgGcoNwBbvzApMma2xl2OU
fDnmLyFVN/Tvq32JbP3sqqFxS5bIonsrISfm49Ss7n3IXJz1AeHSsRm8Ae/o7wJH
KfcwJl9CZZ27iJqPKiCXo4kngJgJrmK6RJVjTJl8tCliAwik9nCy89Ze6xg8C5oK
PZtJCN8cOQGEUOG2e918Kfra61qMgZx5H59sWF0Qu41WWwBlL9GnecjkxQgBjiuk
Emhpfd47DQ+t957FjXF1nMKzTwZC4PyKfy9e3O+oS47bpJPufGDgbGTvOWsGmiJF
q8yglbgSq4h6LLW+6gnuqg==
`protect END_PROTECTED
