`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H4Ys4ZJE4uHk7OaeSCr824AjXtDygCX963JP8P6BKc8LdRarIfNkwjr0sU6Qp6se
JUggHhernUyS0MNJUISd5Dpy2VUDFo+gGArks738dxszJoHrOL+6HoZCNT6BZweR
5NHa+ZWeEyPAlV4cJOgTxumznDP376aO3eccyB2iBc6Vk83AHDSqInCFIRL6ijCy
HT9PX1Jkw/0v25i9rgzody2auz47FYSZqVfrxzxkguKUSRAdLOC+4h6W2ZbC/ySu
8t3Ighrh//julwyMlobFjIChci21adzL0YnRKA7FoanAdlrh6GWY65h/AoJdVTXZ
DR/67dBP7jxaYqfn4sCLToA+QlooV6Ag20MoEgCfosS4nJUHfaRpKCiH+8vcutqw
OAjik9sAqxakmq1eQIF5NnJOPnOJ0V6OUo3jrStNoC2sraAh03chQr9CAsBouVtw
n3dxrxtJgQh7vlHQKxdDlUQUq/3AYbUHfrL2eNZ94k6p/w//0MIGL+b1xpJBm65c
+ZKFndu1Eh/vCP2Ny5Zm1jnS2Xt3yobRn6Lalj7QbLDhsedHqa8BFAisTZNXdOet
1z0Qkq0sNNB57JnHzjujXf8eez/eoPQ9yzfy6DMx0uo=
`protect END_PROTECTED
