`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IHq0BKw7kUy1PaoA8CMqImboI5g674uVncgIEDSyUJhiedV30c+l9dMYgzvuunFe
UL3yNqVZom+NNqKLtEDapPSbl0/aZVBM4ws66iK3NRLaFCs8n2NoYV/rDXjAjG00
7pSnU4fB+dVmVPk15LewF34B+gZhTPtfqIy2T5yc+H94tisUnAT80vwzGU7B3jMD
XaYoJBJgOblUSRqdfdkQK1xuYCMSUUw4nJ2sS+lSgJSczRocmdKeS7SU6PSZPmzv
IdIOSXVdnjkvokJYs+++vhrjk1vo32n9AHNs0DxmHDOwKni2/N8Sdo2dojMN4h4v
Yw8QWK49hV9tx3Bq4ayIA7d9BAErTbGZBTaFeD+zP+AiU+HXpVWfXzTm5OzzCLLf
DFfxwJ5qUfVqBlmmbLlGdTfmhEixSo2inJYLbP1uBb0wfjDs9bBQP/kAFjtK80Or
GPh6lg/MLbOVYa+9T56ZsEr9J7+UmMiZY0zsFHat2jOwaHGGxgRFGibvy1L/rPCJ
zi/CQeVIJ2eES5vf0aHU8aK15znWe/ZnWtGqO77dw0x/yoxt4UyOTSH5lebhEQwq
4NSEtlHeTqbmKoTI8EhDB2geuH0aXl9nXRUfIQ8SQPSszen6/htlbAS3UyX24o7B
rTE34zx1A/nVmw2dSReKguwsO7Va5lehpM2HASdXqTxUcMALmWqZSxEuDY0nVFxe
g3bsDME29XgJVBKhEjOdQK5ykDb/TgaLzUXiguMQCJKCLzvnZoutqPGxH5XtjHf5
q+RKfs6O033oglc9/MXdPKjc0WkQEkZwKr4Z9AkyQ2nFm4j0Rx12CheJ2sdIyqsB
rJUUMRKEzxf6x5CIFZ/ycRkbvRrzWAU4VYR40WDYtmAA6jGRI5KwIei7n82T4XYP
mqcE+yqPUjklkSuOsDVGFyg7Ma8gvXjKjgqR/dS7QsrEQKpirnR5IgzdNxgFDI6J
KRQTgmDhbHQQZqhYMep2DGQYHlpVfkpKdLLZr2XYMi6pIlqFLjMlOIy4PtVm6H7H
mpLtc5a2tdnJqMvm3gmmnbFULRvRKdKSwEV2gjUC+rZS23XF4RLL3TIzPKr7wDzb
nhvR8TI4wuReXdAPrgtNnsue0FgUbcmNTXJjuAwY/JupM5MIxcOqT1Lm2Xh3DC7D
IigtsNSUGibwNX0Bt1jXRHXlWTgrzX2NudtD/tID75rlewe0gMkF84lUEDgWcgLr
Z/b27w+M3T3n//CBm0wIX4slSF62WU3L1NzC0ssI8AdN/9ZU0BiXUVC+T8TPSmWW
xUdChb20An3IB7qvBe0+j3y0umIP+Ju13ZJEKUP3K7/FEmNoaV0DtEUOkaiGVmeA
1OVtZa7AAlnhl2jRmRX/YiXPUjJqTPmB7fSYPSlasM0y7V69ZkBMAEh2V0m50nEc
PZYeBzW6RB9mkRQtNHB7JKT4CLWCzwk6ngCsUNTuGSB/zwV0ddzw9nKyod+6FzD3
7ZuLoCj41NU9L3lzMk1BDFC3QT8ZM26j5Z/U9WwZYHb5YTDidKtszwUH/yUeB2VT
y3EvNl0s8lTqDppATl2oi6H4tfMsUTJYFy08f/uk22TL3Or83HHlz8cf+lErS5xX
oKwNBiZxgUIM1O6H3nwBanpoy242rQ9uquUNZnYuHX7Bjrxs6kToxsyb7mylOVmf
8i4LbCFnmo07kKdTRVuu3j1zwdXg6zvMj2xwWTPb9Dwu8NQQ8dmnnfP1X6PJdRb/
PYu7h+vwFWxHDgt37xcOxgRUg2a6cGjewu7m1+6KPDwRzAVvUHFwNbVsIeUv/yHQ
SW41ZRNNbCu2GSDSdjpiAreeMHRo3ckEwRdGrfEb7mDm8hnul9rkmPzE2MMsav0U
w54f+Sx5Le3IdQVB6A021lP+ZemvAu/2lKnG4A4aHYquWL/ilDM6JM8pyWeeXty5
CxUJrNIxKw8qUX4rE0xT7VH3y6PqLwYXu9Gq/iM/J3OEoKOVnzTS2jX9OzO1xqwq
0ktAJKiM/75kyxK3XHF1dMH1fmYXA9rt3cqopLqSXlMqD5Vkz88qK8tCiG4G4+i1
TdPsQ9Uqv0+92yRDtOA9ib2DXQoJXh1PfWL2BkrZtUVwNYf5IjrRY56AeIRXR8x7
TO7axC6fnA+3SFLZH0iUN18nh1BandejGAszGLIyUDn4jXs8XygynleQEm4M3hbw
3Vi5AyV6xHkoacDDhzdZcivnEcXzp9K/lci0qO9ONpmJ59845c0aS4zIKMERQOAv
7YCk0k2tnP2YQqVlAonIR+IUhq1I2abFCMKnLKEbYVwn9AZSaCn2j3si8CiniVvo
i1IC1ER3lk2uqdPNS0SQyDzLqkdl9d5zqMR3rHH5HtTSBllrYXQgRH/uz1KJ/srB
Tzu8XyUUB8jRbnw69clmyG4X14jLqlzdW7HQXi6XFU+83Mpk4qCI/+VXAgWtESux
pyDpLPU63XXJ8tfS9/jrQMDIkTeI66mdGZTu2M4ldKH7npMgE2r75ci7bce+LIfN
Ovc4OlTpNz93mgvdWe0mh5BxMVMt6jdbQKUeK12sTm0lfFJ4hRyOW5r+hqVS78Kf
9mqwHysvxihqRpTaZ27oGdDIbWNbckiqV1+iWFa9Hfj412pziBXzZirzKN46woGe
TiL8cY+yWxf/6V94U2v6mwTt1vLV2ddRJtkMaRNN+6kDeKzpb6jSng/gg7AmvUyI
LgFC577UfJYba9MY+PaHrDemZvdXg6c27VqdvGEcKZkMtpInr5/wJp31ZOForwbl
i0vwhnLkVwimw4hvZzS4N15J/BXIYw8OXrV54USwk9/o+5V8EBpoxHINozT+AxAm
YAkl0oAnU/bkfknV5DyG6rGJD+i3TC8Pw+viQwX5+yr0K9V8Z+YuijFJJCbh76Pf
mC6h6423jYxm2ZZrMORyqD5SfXSaSteRnZ1b89e76ZLf/nHFYdvKhcVeM3XwuJbz
jGrOxO7cCF+cFbmQCN/DmXx4/zFA07M0fl6HMbqu6pjzBRjdlMoiIaLyIzm4CwzH
ZyTHii4ufjRfaT6Or5oXhITAwrOxauridx2mQYpH2V3mRvP7aA4f/o7Th25dYUd7
5ZMZNR9VAGg3S5oVnLkqe+mAS0dlqtbIwctp0jZZjKp8qkbP73R89I/bSl0FX0cO
Yk5CV4PKOh7WthMSMHpqcvsote0MXRBZmaFv0EwQaYYFnUyEzT46DY0OId1nQxK9
DCQKNFnuZT7pS+H0pVffxSWcH4LRr1y6Gvl0ueQs/uz8RE+Y2vUQjQK1m0ymhcW4
IZpYArg1Uw02CjP0M5/zAVfLV0eIncuFF2g1XtyRkSU1VnOjn5Z8eoQQIzJrQzkn
xV4wJZ0Bk8zJcOD3bEwbd28rfWwTpvIed+m5ZcUqhEFjjaq/D5sdQQtEKdqQXk0D
DjCuqFjmZCg99ymJASsOU3Tfw7QaxhNY72KUX4p3bUVxnKDX64G9QruAUlSKn9Ve
tVwKBupXSZy1tKJxW7LISVIkZ7CQSQ2xjc7lZZRcXdlxTDpfsASXqXVt1PZKOpxg
XgoMBv4nxQMpRhcM53RIQ1v6++5S5kdVYyzgdzLCdcHfRO/MIV5IrCTOiEwuDy5c
Ojf5srzyZX78KXPPGyvjrlulHRGrV3fJKi7nluCnGDtrxm6yrtuE8iqRGZjoU3lS
LtdV7TyX6v9DBjouyudQ6NRiMhw8wtNbT8Gsx2DahMCwC3rCgI1kORk8OmRMECZl
wELaOq4C+j3FhS2kCyG/34KAz1VVeKMUxIJG3LNJKmV7EW3PPGQX4dDo1OeenoFB
sJO8d9X0H4b6cJrt2hK9oS7Ph7lqRpIggr7uYVIteOe1PsSHvzG5s+i2gMZJRuFu
McEI8bBjpUkiaX+MewPyJn0fwwzsQ0ISyRWpKyEVj1tTPqanUOYLyg0ArgWOfGPW
6sLlXOgYiUDv5VzG5TyxxNPqz8vYr0tTj/sfoO8dNdCXgykEnU2ZB8LPnTB8s02B
1iO1MGpue1aoD4BFAvWfvv7F2U/+AHrgAna1TKykflk6r0pDyoNDxGoI0MZqUG99
zF05p+AgH+Pk2WCI3ntYVpGHQTIqH6kfKoPaS7g99RmEFnJJAmhNKFkprRjdoITa
Z/cBA6YCDOPLZmtbYyNbeHgAsDqk5XbOCiq4i5ToqRC6VIlz4TzMJq5Jtclcyuh5
Tp6vzfyezYMv5+ySfK+ylbu+N7xqNjh1Zxh8RGIo+Tm/20YHHWAgEXQFSf+WPydY
N9GsEtmsE+FPHT1GSQcQi84BW9R5TckGkPKETPST6jjHeT0r0ujmUWT0tehiZEd/
BCot4yHgBQhnl7tWWvOoUstoOUWBlTtOyNJEOxmofPQrcCiilMlLMU430xHw8EE7
dJSWNFRJmpdrfk0hZOnNCS5PJSJl74IRYI1Z6ubAXSBkdCzrrlVfVRYCA5il8qVk
GWP15zmYVdPSuniBgrBbkBwSkyz7mDBQ95Cq3bIoPUrBH5ZY0lLcPSfcUzWLSyD7
wWw6bAp1Gip2NDpaxayTSMX18xzJasvv+WJQ04PLZKEOk1Pg557kqdlygkcPULQE
o0Jt+Vc69MFWxfoYPfBD+zhhoSs/1QsKghmokPyU5ISvwaloXfKGmER/LD7AKfni
g0ob4T4ObPFjZmAx8M/R+RVKTk/9e/nTAYnUnDyC8zWuRCTRgwuEtN9xhrg04EcL
ovgEqeQ15z+cHeNp+JDgAhsQPpn5LVM6HQDNZj6wz45ciS8p7229o2YlW1cpQVY0
8oRYbSZDWN8cqOX8pj9Zg5Mm8wshKR7/yKgtkeIhJr5rBfCdW/dFg6z/q4pPGawn
6LR0M8EQF507s4xBelsStlYlRs2Eu+KgMROQMXA8YvTDHEdsUVHib3w1S8sAYU0o
iv4G2sMLyhFOyprHDMXHJMC5n5VQheISNIWWoWERUCeuBKLzSZjLQgeO7m8GGrQa
islCXGHC/e1ofmI1zx/6Ohuvs0qMVwpXqAIOF/x/415S/rVZNrzCNEoHKs4Tp+4O
aH8r8UJl/Fmkj/q2EPU9uwzcWxzaj+HHzywVll6u4dsYEdL2lLe8ai1lfyl6MK4j
bkepFXDYoWkAxHsyMvLxEP/Tg0Id80LKNCoDofIYWb9up6nHBlG5QE9/1dTq/2Dp
qHFNHPneMgR1uvTOahxAs9h2ZFiRjEe8/52LzSU7Z2lL0W/QSUaFHzhXTW5zLFE2
XJWoTkX0DFVAwriJZyHK7JpLeMTwNW9Mm6lZZpJMC27fOFsXPEkt8z3FOUkvToBa
B2NsVHTUdy+86Ai7WZ7uw3Fls+7YF9JSTpfkFucNFupO4QBT6s5NrKJ0tjwOMBtr
1xUwpxQq9mCLg6Olys8xWqDiVhUyYPW85zxYleM8N8HZgBHyLoLQIbogtuEE/6e3
mmQCii1l4fRf5t+9ly9+FLvd73hiwqP80vnEy7WMZnr4SzLylC0S3OPznT11PwQg
ylJdlE2h1OlrECmGYyGTB7Gq45HexNfaKBUisO53OTfi4XN0BeLDpj3WXsz62dkF
`protect END_PROTECTED
