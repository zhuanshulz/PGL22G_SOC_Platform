`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7/GyDK1P2u4aueCUmq2IDvsORwsNcYwPGknUb9AerxRW6CexalBSp54h1oQ46X/w
6rUYCX1dgCTi4ZEhl28jU6+/atnVO4nL2UKqa5wC8pHIU/Aej0AaPRJ7SuiC70wm
v9+Wy4+IrVgHtk4F+cK78wQXD0AsB/smVOjbmjXIRRKHOgi7BRrr7nFxc/RT2iZw
CkuQt8YBLspGq7VltjQuzY66zp5o8+lhauSv/YeOIN32PxZRcI6CcAwFCChNduYE
T5jKVm6e+YUxHC71hVyNG+J4MARUFZMxFE1cXTl/A72wpjqHPJoqDTGg+K3PuZ2e
buoyk+4RmbsRRQdOKL+qti+5u3CyBHsuDUiluBSirmVwTXXOszUT8yAUsIdg/lRV
PwDEr8PWcfabbxQrlwHH6qemDWI+AoPtRlfY1qaAB6r8lfTqe0FhMK8klFn21TuR
jrK0fk9eLs83Q3FGRszr6jOfRhBTSdhfGxHl68679qf2GOg2/Up9hmOPSaV75rBp
yit4n3PS5do18Gmtb7D8TCHApHHs3jlKpgky3v0V6ePvJHFaf6Eu+9FatRrFnyYl
OElXkt2CCmYR3GLfl42HVCfAqjkZY6YNlG+EaAzVpbEIjogT/0K5+rUEUG3aqXal
nLRyQZQieyBlA0jcIphU9wSx6WbaaQYpv+mvzlnobY5ALIBgllGGqy0M8rCkrQ1f
QH8ZpEHCknX2jXtyjw4gwa0DaV9ihWLsgHsoKzjEFaBWSjZDghiIq4X3iKbt7DQ0
VZ3rFF/ElPciEpvi2U+492+n9pW1pJAnu/7Pe4A4iZ5JGzxI5VrDzWl0JXj0klwW
ib5846KXIq+TwloztrkdVO4eff9qim2Hph/WUmWWMyU5kcr+i9PV7/hr64zljbTR
ikeizujzkGUIQOgOwM84l0v554zFgPMwr7UB+WrT9QjjDVVYcU1wXqef2iIW7Zdf
gstM9vGDUt7hge6qjCFi7YMedRmNz0YjLYm6THUoYIPxLrtaLT6U/d7VcjNQ+B7M
EZcK2AyRi/cFJmZ86PN5S2JTYc4hibFhCxj6hfpTVpYUxd5y2UnX6MnLWMWzGeB0
gXrwWKSfhMO+fh0xLngOMfvq0SMy3U1lsP7zhXyrgekpYhMGODesIwsFEtGoer9N
yr3ivxsXM7ZbLHQB+7k4flCsD/Cub6gYm0YH4Y/umLtF4ak9KpcPL4QBNlL55oUd
+E/PRlRyOUdvHcTYW7O/kQCgPR/RTfXhWqQk/4r0vG1omOUiugyFnT0+mPS+7OHj
GRJNfiMhNnhUH/fhs52kDBskpwh7Iq7f467XxamPoM1aol3Qz0hTn5zbGZhVBgZ1
Hpp3xXWoCEGn4aFH7KleGFT8yZCQC5r8nTcp0fPEwLx5P7Lk0F0H9GZrWbo25cWO
yhZKEMyOXPB8h3OaaF8DWmMTX7rG621uuVgZ4iuegeO3z0cUOStrZW49W6tv6a1m
9w98RcPebnmsX66Oz07nllQceMFngUHURcHbbNOohp1mOPmufwkhdsus8mApnf6u
rf3RN57vH0cU8uU5GS+4HNU0VIgKkI8T3gbZmg+FaOE5aCnkV0O5yxxWvsKHnZ3+
NQVAtC5GT2JvQmkK1buNskdz69wLpKdXDOGkFvDJeIE4YapMNhjGKARmGmldjuw5
wXFY72cbSQxVzEwinpNbE7FzxmZtmOiQu+xXXgY4HIeGqL3thxWQQys7FtSUb70v
4P1nhC63vJdS+PBKwLnfoBJrQNFLSnoCK1Lie465iLSoeUtwbmbeU3b2wQ/QqGZv
A+JzBJ+05XF+h9dKtuIIEnc4P6dbh3VTa1rBZ/VxH9A0zcs055VhvCCmhB/+ub82
jYMuB9cjM//2KI0wQXDtDdxjb3RS6h5CldpKdQDldIJZYDV/xH6Nj9MTWHZp9Jfw
IAapsLa5p9J6+p9UAYCLzkiE3zh6KQBaOLJNkqtEletzxPO3Z4KhJdKCiMocWX7+
Fn58OipoKVY3KE6xXGw9IjlUe90vWPCK6fwBYXzGwrrbjn58r+Z1bye+BVDuQ3Yf
+0COzEGLfgzNv5RA1nyI4snWNmBAlqrDYJgTcLniEPTu2N8ApAI9paVkyX56WEQj
8BkLcDDN13sojNwdOrLDOQ==
`protect END_PROTECTED
