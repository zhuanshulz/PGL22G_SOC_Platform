`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
itXVAyP9wQVP1AzXkJAF0gCZCWWqH69BFzV9J7Iyequ439ksgoSzm30pzYg9lnEW
7XDLtb3h6k8fqbup/b3bEUla51J9BXLxfKHYzOrUy8dqnZbMJUZlaXNvznh4cofO
K6TCL0ZShRUEtNY7K/EZVpKibIbDEeqUQY9pto7Ppsbamx+KNp3bO5X1RopWMIqG
GnESP+U5xN600F0OZDg1qj4UM4/2sf9A5EsoGn/j178mAN+SrXRWQJBjdlEgJJp1
XibNR6KJuqFp/MkE91BRh9XNd+Ap5/6RrLAQADhqW6YXe0KHtRGZa6hx7/97rrFJ
J3iX5vqmlWi9gniMgSyVs9VKGIUjL9dJldsjqX1gc8KiG2mSCNVzNcZa6bn1Vj5f
pmrYBPR4VQ35q8d0qvjm+GKkp2KGuzkhPpiDcZUbA8jnXMjnUvT6alFONDNnqO0g
06lhZC7r4saHboW8d5EhdS1Khxuu35T8YGz8S/je0XTz+VygelKtq9pJfnCrwyRC
jY1vT4ygOscJ3wD9bL2v41ZeXNa6lLlsiGgKPFGNG/D9Ro1WmQmCztHd9sFrPgcZ
BIJHtkMq51NO+VymdlcMVCKJQ/YwexCjnFEnojFOjNIzUGlUiwggC8cfBREu5+Eu
`protect END_PROTECTED
