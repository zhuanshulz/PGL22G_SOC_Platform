`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9H3qIKOZ8tPGhUJDgT7cei5P+sZCMmQfCVqgUysFCdS8G0xIRMYVSwxhd9syMxV+
a/F2StlSksGS+VuwZqXbnygK77J1Fnn1yNWwLhPwPCMfWIV1ax7fzCivj6DqqfEN
lLBPLQJ6x9YOrzD6vyZG/28BnACaUsSVYgxmoGeajI5Mu21qFw8auWZjBWGVUpuU
sQikJKvWcwZFNO4PHsQtd7LWXSMLOmDvj1iq0RvoGJKaohnIAG7pXh1TPapLOac7
4Orr0SpoVtrOyPScLiqXeR+eX6VFS100+MRR4dPTBqdmcsgTTraB5L0zGiENCQxh
q8KZ9nzPzzH8YEy+ceGwQn+UdgvN1iFF1BrJWQIe9/4RR6wIqlhBCK5nZHYml3UR
fPGjy52LDejedsKypH2utDbTHPCzr2M2fhoiQRR5aS2pd+0aCUPnJmwmUNh42ydm
0hrCRJ17gtk7QiqcQE4pfnanikock5RYsg5LE1UumgEjXPZHu8yoUUDVUJYDhNUW
7/SYa8kmJuXyBfRUOSpvWn+84sG86bgT8AAC1qU3wrYQHbRJyPPJ/Vu4eca4D9B4
t8VGQPn8V6UjEjPelhj/MF3k6j1ZNZJqiTv+JYm0oCuHinP/ryiq8pavXXREI1gO
95BdKKaL3Gdn2ANIPUeBZKcDpRPhVaSvniIM/JVhjT5s7uKZFlN/vVc8FYl1srHM
3A5p0LrWT9edIw1v9DwWikDnwPjxjJTIgQo+oNKO/Hr/nTY03y4r2y8GFeG5owAl
/+hQzTso6+st7Gf4ySAWwECr6Qjbym8/sexLArwVwtezghASH00MfsZY16GBkAjU
wMnaXf6BDD3iEtsXCrOqH997pJqJyURjcQ7FTG/Y8yrLn6AsLHegxIpLPOJpCXJ+
QZrCYDlIbHSQvWypxIvJfLJR5/zNanIjnH/XDDcukSoGMnFdiF5qX2VBspe0frX/
5sCXgHxd2/l1wpiTr3z7296ukK7PXEMQwhafXwURUjN4P6Enkl2xVhWg0QtKYXJS
`protect END_PROTECTED
