`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N30zIgZqMmZYZS1djGFalOJqNtKUwsF1WF2j3y+4spqNpT1qKrrkS/odHlH+fB+X
0LbIqY9avA+De+kqpzaEhw2rjj6CWOkCRm3EWezljUhtyQC+h7qe1h4BiWaxxMn3
fzk51OhKljjopU0tuPnjFkAFXnjNXZlAL3ZfUbbEbf1kJoMZCAn21nYb0Mqd+FbU
Uoa3bsGiyCgEUX1KKGnGYXuB4jJu91klsSXCmE9MObD94M6ifpJhwmE+5VMGYEFJ
UQXt9sr2t2GNOCgV7bcSdEL4OxVchIRxDIJt1SdbI0iN0Ks42KFHl+NLsha9HF6l
JMuyCR0phIIXtTHnJ/cJzQp9gWMgMbrkH4uWM6wGaH0WzdwsYdFdW+Bu0WCHyYjh
7ClQBuKl9LzsdxWenXe11GUu0+6r9yTfoUsPOqPPkgG2KcRQpJVlQDCvpgpj2vt/
i2BksViAHQgjzewepJ3oFe7KQlPBy9qB7+VwRf1yrAMQVmmIGrpqKjpgCeaK/K6l
QHrXCpmBmEC30wQjYmHHM4tY2fvkeLiY66+Hg0JnYs4rTOuZppqi8O0yLlc/UFzS
cgaQk+XoAEzYob6cwqBsbMiJvfp1n7GzY+0XiY9wcmm+8IJxmxpLzI1zFvssLr22
WpzeDbaRm88loqM4Kqp1PCc6hQhZXBPy+jnheY6+JATlBNh4CrmjctS0dQN1/jj/
BFaqqL3NNzrzjZ2M5v40/BPqjV6qPiBKXI8r6kIAPSdNNw6cP4aXgXcikc/oqz+x
nI17V1Ioxu7qdVCIc/w6vQ==
`protect END_PROTECTED
