`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JUPBNM1CEm29j9nJ7OLyjWPlngFM2YbdfIrUxeeSEQ6y/AePdIQ4wUs8m+ms+8pX
ohfTbd5qa74jEUZCwg61Uh4jgHLn9/cjI8V57lBW87dWgs0eY6G70HFuDhMLX6FS
gLbXjLb9xrNvdYI+FOD+HQE5Nz680bQLBJTuHYPW7QT0WOpXo0fArgqopEhHg3yT
Dxql5z8j5UyE5d5zg0AQES827XQ6blWCgYvB4xSJII+ymSAjf41DOwsNAssJ3erc
9SGx/vTHuKau0ZNzvJSFB2lWNWPGBekcctAZ6MOZGuFe1M+2U9etOiUDXoxSoHFY
KlZ2UVTIM4c4QCVKrGCFWuC9tbpcB2sXdvqMo7e99I/oKH/s1Iz5XT1Ot1FerDq8
lJJmhJaV8wMTedtxzdzVC1I0yg2Tfz6N+S2fNkPBwbY6acYOhuXffnF+Jndvp3et
JBNhVeSeH2Fht46fOhW0jcn5Wuj2yz08Ok1rg/P+GSs7L0iTRPv0DH94qYU+O5ga
FVQkTup1Lvi+IafW3dUCjqnx4kuQNIlxtDzSL3LZqwAwedff+px9jAzrTKvIv9Ry
n6Xol9D8fZHBJzcaojObGJmb60tEHGBfR9gnwYxuEwhoaCl1BZg/pVoaCzOCDgkN
+83hVw16ODee+MXorAzufaOakTYaKXWuAx2noKxekPpCr3aNI82Lu+bY0Jwr0sZc
Ia4laa2+sK+xjKJdnam9/OCnC2z3Ll/TUC5+mmm+5ICKttP7/EUURXhN65KhxUs4
EGxGukjgOOGqHSEvl5UBE93xFge+BnLJT4rOLOhG0LDK41FLYFYPzcH2PqhYm0J0
YLv2tMuReOLN0zcocT0tPri59qwWKMaUnPMEXQ2PEwJTdAQrUoFRAPZXv94Dv6T0
lxL0QgCVKkbiY1Lt3pxVCEF4+u+/SQ2cyBWOpPY7gBOOWFENifOGJYQEv3cdECAr
xgTx+d+FRwP6/etwKoE8TzrXfPUJgpQfeXPSaLO5gZj3AWE1NOr9bP8T9laPplNW
Dp83CFIHeHJ0mo/1iLyJJcXh+1YOjxP5Wj/ExXDmQJXAoFqzap7bz4hCuVaCTTYv
MSJTbPc2XctKE2Nx/weNQ4OERfY7wGKgVVYrCMxuY5gLZN6vRkLQM+43CjQgM7/Y
HajkY3W7KRU/zIqq9g3pBAoVgUSm3gjjGJkrYRQjKh88xtMsDbQZ6eqnDWG0HwOz
M/YEkHRfwImQrtPyQHmjyE7q8fHQVboPQ6w9a8h72a5JK71Tu5Z3Ca1CbhzKwGj+
Qvf9hNuOSMch8+kYb3vvJtl6W+c4vLwLVGLGAWh6Ag2lV+exReS5zMMjTSC5Lf6f
rCqn9+p853fkwGgJnHCRRD2U9ZqIWvM8SxkcBjkqF4nfQqz0rsUTzYeSPjXcUbGK
WU+RIVsfPkRQaroSiOJ2rUT38foprlHSNZDTiQVSCCOeTY8EAyHk4jp7Bs4zesR0
6np40Z9FKp9Z+HekapZJVP769Hisi2Ix5XeeYYFe0P4WZTa30R/JaA/C52I5sgaz
5ODZlG0ufYF6qD0QlYn0A173sIuQmWkz0cwtbIvSmQRCqXVQKeo+Fp76+ps3nyUX
K0beGHMFFIX7oQVCV3fnPbwUYnTX8514I9WECYktRQLTjouFZcE4TsMC4e3WKX6a
PUGilqE/NIhH9aEYcxFExnMQkpY11+E293GisezUcRLwhtd2AYFlDHX0/Y+hZl1v
MLKROpJcVOT7o3iVGZpGGtGRTQZbY2sIbAf2oUePB+mOhFGzkWOFNzGhXZMvu2Un
SupPgQe49Iyuk0oToZrr3Y/HRwy1ntF/rvVVOMbrKn+bZVIItFjmz00PFZqfJdjH
EPfaQwdz63aQzx0ITEZN9/WyJBNhpn+0ihcInYfZb1kc2TCXkzwxFmuAC2LuljfB
GmKLfR1/rp2zExIUYcryM1QzvD5dOv53PIrkBhlgsgQx/j7phZC5aDbh20PDg1df
+p52bf4s0Sb29OOM68KKmvFb44DL5XHphH/nwstmpgHTjvxhWeHH7vEf66r9ko+Q
iEnKXbwZs3WB0CNeaf3l63BKOv9MdwoOgh9NpTlL33QTFVaN6BplNpLMTPLeY+kJ
/cc/HJPfaWGIRP88g50qNYCq4KJba54xqOs14QZJLBdlG5eZ3wR2VB/KGng1nuwI
KiP+T0oddrfnuEUArjtpTgpqoJha4RPw4lqWWtfO/uTiqsqqGJosy4uG6vuaQ9tL
/RwGJ9FDfnC7DRNkSMXW0PhdZvsl+NZlR5ghIv/EN4NraAbLK0m4qYvNJYx6U11F
49aO2SdP9K7t9E4z1JmUekIcXDP73udc92kqEZ0qh7oiJSAtF4mZEyhZhcB/krYV
B0L3cseEjquN+4Jw0+fPqdbOJzTjiBk6z/IyGGgOp6AWi2tGhz7VfnVME39ZgD5/
tGheiIXWYL7AR8Fa/5nBQDd1x0FeHnA2o5kvGUwm9GZrfcwlF+5YwIf9IhA7UeeY
ajVaEqEsqMTp5ivBACScHqk0DSeHr2Kz3cx0HHRLZLos2IO6MoQYv2T3W3ijtUDI
L3cRLzyFEDcegNqJMb5aftWkujE8d2MvKm3qRjO/iSdvS3NrP3KJ4zG5fx6cm58b
WVitPav+G7zesQOUfdV3V+0VA7Mr2RjrEfcl+vPXe4EGwhPbvAVGRNKOyO2rAM2e
awUuwv4iTAE+/0PSBvm6ke747L+fPCq68ujsep78nzp1dMTg8R09hKGFoAsvCFMZ
0bk+Yg490rWl9KDVB2vaFfl1kgWAMpQGztJ4UKPFLXBIs9VJn9vQSLFI3Qx3usDO
SAD2qasS5gFvv/XZSFvwRhTumnF2s31Be2Rw0/fhTfjSLkgV1bEgBr/Xr7iRi2X1
hIYkzfgiR8aOsjS3OwvXVk+Ysov6dT5j/RC2kF6hWCt2v9tVS6AcDHbTcerjuXWF
AzX20SeYcSWgbIN4t09Of0e5bAQDRESwEIwKgZUomW80FjmyUUPgz1KBB0fKEHtK
j/SxwbmAGM2gRpB9PBYPrwmO5Les2UOZNAtt/uLzdVKnfpdLvtxiChpR1xEOAlDp
uh4BvE1sy9J75UBTxX30Q5dWF+VBJsxqlqIk8fC8HanS74B1okeGnqOKQvk9DLfg
Qe4w9bnM6TPawYYoo9pxo00E6W3N5VNruKvN5GR8IC73MQQmZW/I2MD5QyGp+U8a
OZaTGXQyYjbgLsRmZJBrfhLTU0UPwq9R6kJ/Y6tohwetTE8Lg1c4C4ewetSKEO/o
n5Q7QpyT6ecj89vvNeBBJdB/DmdPeyFvytCXJ1vVmCcijuNWccsRu2EuPE5KP2SQ
kxlJBRxNEABBdQwtesUofGrFjB3Au3laSRerVMh9sSVQ7se07qBIY8Ch8gtYcOim
951qea21z0AZTHr4t333Tj/TX9Xq60YnC0G0t6MhcYfGJrn8O3AVmcPfxceKZqSI
7Z8Bg/sIJKUJ149/YpwJrWkScT6ou5RxcpssfZr3ouF8mQRNhEOxbETUmGdE+AYu
LXr7e7kQTTk+Ybpb/8u17fGfUGEX2D44BWfpXfEn3w9ROym7765qN2E0IFU0RCrq
bt6RLPdSxpA1qOx6elhkoeSFlj58L/1if94Sgv+umpSOVIYF7XP65A3hASaKpIhb
iPLfXlB/A47ry9GdjaDMGrJAvBe8/xkuUlCPQFJr1EQyjwC9HUmfQqz5/4CaGBmE
1JozWCTIymgqCOcc5XQZDwaJmIzDGssNYWHVJM/lPSlqYJopHtykR05ZmgxYmOfL
AdFjZS40+H4SPO+nZICR7j3scwHjT9EgPnRC7wg/8Cu4l4/7HfrGz6do6f4zfE8i
ANz47Gig7hi2SM4UNwILWds10Yzm+6FF+z6UmMYfdmNgLjRIRl1kGI+n2XAI1GcO
q6t6/OhyQsPEDh8mclmlXuGgMs5xWAqNvbnn0ERO9ceCAsElrDiLfa5VUAKUWhKF
EbQtDAY+jrIx7JmEEmJjLKyeabvNhzF3SkhUOq1vpNeEoV1kSHEvlwgOieAup2MK
JzNTrsyxhd99zCRBos0Up40Pv4as9Dc7VTjEsmNn/TQ/sbRu3VUy9kyYb5IUc8WH
ekrZAJq3+7Sq9Nk9xzJQn7nQzba7txRtOalNrm90nfYLO2tzBuLe/0kRQeA9ciuV
taVRhqXNuPoFvjuP7eKo3h3Z9+LgA1Vkl7+/LMc/CSdGjegKFSJqSpvK1iCJM1hn
xl9jttQv3WOMSjS/+JH3I5JyDRwoQ2RzbeTLqh/BPV2HxMl2Ul1suZ2KXYiJayJM
UsOsbawOzZgLKnX68s8MS/Cah8OXYMGWh49n1p+4028Doic9liemjQCeYzfa/kG5
JfRLDCKQlypwys5gkHrxhew5sQtiI+RJZ5A2tKpMQHBNjPKQkPIHUDL1hlCAyw0a
eEnjXpxXd0J7fDAp82eIdVVkmPxuja3sQ8A02AWR//VkbgHaD6o7yXTv4QYoJvKy
o3nxxbm5lhqhhI/rXDfzXpGJL4eahuJb4qZp3qPknWlpvYreo2bY85T5LwJbAxbM
ierN6hJYlol2HrV/dpzz3Annol32hv/RYaNrL8qAIQDblvmuiA0+9gFm2DtNARGS
aH0WeaAB7jzJrZTYYYkj6iswTDtaSTIDOoYEFIQ90UnI4KoHHv+yCm369pa2uycX
u5MWXJbpLMG6NQFq7dTLdb1QW4Ld0Gn9scrxv7hIqptcJc2tDlW7b/C1N2p8VEcq
w5+obR9smxsDCbc7Un44ReA6HRW7y+3zRCnaD4WvT2aRSNXtjAElWGPCTy3PXdD8
zVdpJiIxeSTCQlsQ4wmJDnOVRqijWwuS/9dE8yOb5MrmhtjzHLiAtmmBg5XgiA1t
8hBQdyPfMVGaF7l6d64VuurOGbPeOEao53Yg3hw+lgmm8gaV3EbJVOeIIrxWPRvA
YPHl5ns25qX2goCMILxm01ewhhCIARVbPfrkCtyyDPJjchyGqGb/diWbCnZEkREB
KX8IG68S8dl3qZ5OvDMbAJ2pXa3XISgJExnEDHkFczPZapBwqXjFx3EqJlFDY2Ln
R4xgOzouR0N7ObmSXErw+/uJOlwxVSkNIwqYS7uHbaur0qlMQpg5ua5MwULHgt9F
qPxo9/s3tU/kwqV5LQMQF2GeZ4QGLcKm5ae+BcJ4qhHszcKhs35UHfs+2x2nqNLs
+/csif1i+5ul/zPRSHg/fw2hRl9GiQGTFsOWs969KUjAGnWTDx/S41HsKYnTkfGD
BG3R2oJaIEu2dLWVQEcXw7w+YG33QvOLWk82C5WgXXLSNtxfgC+Gh0o/ikDwaXpd
ODuAe7SW65xM7k+c2b5THhnWVGiW9ySTGW9Hj+7fVbAGxOGT48dbxPpcvoPeid9B
OWYedCbmYH/JP89FwXvd7ucDtrjJNvLqGP9nshJYAzjigyfm2AZJ58ax1KVqmSWF
eB0G4ogtBXJvqRqP03a+2xkHr6QmETje43DG1NawE1mcCRrAiZe7qf50cJ41cAbo
R1YoPLrIK0LM8uEPqrhB4SX9PFOPRFmxHTWz0LLeXRcKpEls3XS20gQ0qzm+jaxq
WmDmh2pe6qja/1GEW8VveLvLaUj8lQyMwJuHaOkT34pHGpAFZm5LL/TB2Qg6kOWJ
5SeKmHVcDqBp5hPArWtrk/jb36wz+vaE8vxwR9ddPu5iuFrTJg5QHfZMBsJvEl4v
8Htpl/PDQWHNVz+1tcnYNqUohUDD++jcp5GK7KciaPNpelxMwjTBKEzZZy5xuc4A
jHx3RsRlatIKImkast3iGgQRnemv3aoR1/fhy743xm6SCYXLoYTv3tT7TA3dOMDr
IhSTMtsxxpjPSlHfg0lEZtpX4eYYjA0DfRY1jHUp7fIJCEmMmPPeLgHIvtYaHOsM
C1j0nF+tiqShBXS1OYOZdiDMxmu8UCi+ioknDB0RT2mZth1SHqmgkhLIboA6jcGe
rgAKFEtM+ddk/ulKAv4gjEztzyXUar3M+bgv5nMyMgWDwGu+ny5/d6FOxIEExx4+
J6nKIvPCVMWMDpRT7EZyy2ThpY8YLrst2/K9EBGc4DaUixyXSyUfsYk9iSVvCsJ5
O+GJ9/sEvhXejkoyyZ97Qe8ncGAQr/DnPFz9ofv0oe2bn0Htbbwiqz3E7RFmrZWS
+Fwei5bTMxxB+Njnn1U5Uu7eRZatRmTl7fPpoHKtcYsZYYIFTWm1QEVKQJRrlYk5
Sd+yhgi40kO5iBfZVDVuxIawYsVZcPeBgUplDGC921EPMjMgI7+RlEm8OPBj80d8
Sp3pTqu3HQtFYv1RiOGnR02BEchVYA55BRQKAD7/BJX07M3e64MQebIg8ZARGWfe
7Wy14zcmZ1cG78nNoPnWk/dD10hv3mUwlGbSfjMsVsy210l7cSg6j11H9CLiE1ZH
k7f/tIZlTNb/Fzq0T638nANbhmVz2qC7yY3/0wpzUKWeQqKyIrKYbOncFb2+/3Tk
Sd89ZNnaFEh+60u8WKKPPT1nKiP84ahDjaHDVrjgcoRwerJWKSf3igipWGIUAmj9
uh4DuIcSD8y51CaNKWJX5dxwxGG2ibx/O0y3R1Vym72+KQ2E1b9Oce/j+Rr78xSD
R/OwUw1QQ2KNGCqBtPLMT10M/sd6ripRMb5NBbZmyHGDiSbslLpBWaahhjwfKLcO
91Zb7HsL09xIKtg3gTBpJYgtRYm4Cha1y7/5SMeZKlXrm9AcIg+yoKFwILxjJ4Hn
XfbOtTlDBR/sB7+aaCAOWmG80ej9B5IJp8uuMwanr2pEwI6vMzsLZEvBq5E1I27R
t6d6WcyAcaiibozYE8174myMPNXegct31yK72lR0XThxSmeaPTrALyJdFTN5Va/i
3zTVN5rdrHq+mSCLZM3rko9ZGrO77L9t62sgLoTGfwEzEZmdH2gmv+e8DngT3E/J
H6XVKKy99AIyR8VYYMV9SM6d2yAZ7mUO2UXD5/Eqk72NTZfS8VkIsYryn2/9s1HT
U6+NbePAm4U86qllAvGj+C01qHdKHXTnznZfA1S6ld/XJSd533/MfinCb9PWc7JJ
Dmb8ArXanliW6SZ4RtmUXKaN1OUyb5El+pwg4ICdUL7qFKPpheL2lJimY6O8xbrp
Fx4tnCzVdE2zZJLkNcxXQ/jVIHd3j9dKPorQk36cO+rg89k5cyTMMZ9g9P5NB7dk
qrvSgJtNowLBP55j1LNGrH/UgxY2+1euMz8WypLjXWVJ6GUYl3nCxMbDu7we6Sjq
p35+MQWjgc23GT34cDhqydif+yZ6f5PJtaQ+ZqSumZV4Y5D0mmB2KQHzk10MAPqu
kp+X+DaAv/czYDU+092Jx8A0+0HiMmWMbHmlgdiA2b3MpTRrzd0hBkuzR3LINlpp
ZiE81ttJ05dIhGTzlbmeberplSRbiXbYr8qRWITGWNDjMtiqSGVqYQl4qXXdLyqp
srZt+0yA04YsAuaVgw+AtbLAttP/WVUAwUyCCUJLhZWYgQ1nBQd0Mt5MfeARtIN3
OLjWa3/ard2EFXW4FePgKVPdomiEcNn5IBycpVhiBx0O5es/QcCj6RWJoNLYFqQs
iuMEP96o3fxYDW5p8gI1PP/EnNuE9PedIA5/eP5MRCJHWl1kcXjtJ3xu1BzQcoy7
YcHtS8897vQxdWpTx4jeD+mYrM6TG8Kl4xGAQzd23Od5IyR7Fzp0lmUg/ebHWipD
QOEVUgRM6uXnwcm43d43WXW8Hj6O81oajWcDvGF4evuygUOSI96971EkvVs/P3Yo
Ef62YWjnNTHkmaNFBRPHhSj4dwgSWiwNCjYDNPAzoFPBCF4l96YqiniZSreJfKT5
VXHnSp0Knxnud6G/a1oanGM9jPoaaovzrkJgOY7+NPkZHnVp0eqecqkccnpV5k2w
aJZIzw3H/tNHNiNNoLeJ3H+MNONI9riEaHx7HykfFrxb9HxTub90CTbFktcUrBj3
JaFc5Sg49GOD+ClLjTHx0tNWAfIad99v68qeOg4d/9oYC2DpnS1n8qRO2aaiJFMl
YD4pHgJwJuuIxi7CtuDQ0aJw0hF9NJ6b9Q1SMmJFId7QOe2GfkA7N2MIBiM5RBd1
+s03eZNfixoaYFEZc6maxrA/R2fz0EJIzK9FOFZXE+Y/BKvYcEZkYSvs5pJNHqzd
wKzBwPUbtWuKTGXPqs7ei3rQQ3LNYClGMHGjafuABFuuU5E4wbmjh6uJ8phpJzev
pvP48RNmcg4FDmYx6dGk9resssaqbTVUs6Dm3HmYNOjpzOyTx2ih2T3mFKNtfk3i
pYOdkYbg4vnMEMAgV9ESgABA5y3ySmxfhhCV0gdDPXHplSXJL4utfHmrvC+yfLGi
QegTmMk/TaAISRUVikCHCQk4i+uH+1ODHiofTnIDNxNbRkRxHIfo9fiKCkBti5rB
ogHJ2tE/nNXhllsq3ImPKuYvulfj9VwJq2OsAQmqPtjyS9LjU4M/zhCj4MaABmie
svz66rnagrevV6bsw0anfzTInr8z9rjdr+vFSJFrui3XEB0ZWy3kbMfnoPqWnzLx
IrfTr17ScSWbJJqzsVKpa4zRSc0VavlAjFMkr5DbHnt+fzFsCNQrhX+46DXUAaaZ
+LL/iOKKo8IocfsWA0KQRGxB3AERSFkwl2OQvWFdAQkDAomrNlomJQ7HPxt502++
ar/l4tBy6+V+U20qjdWNSNt3eWHh2ClcoZReUNdz23l3qgF5HZF9Bx6t3E2oMMsB
0L8C8mZqUde12Q4tIvK+Zni4sYGvmknefkzSNHxhQP8wDgC/dA+gc3UqfFjqnMBu
otcrGC14Kz2YTuHpBhFPuYUJ0Zp3ZqKrSCt+CVMQ7CMwsEYf9ufxGDfulWf0TIXd
ZN4Y/he0yQRwGAdojNSn/TF6q8Oz129Df4SUpPu/E3+xLRKP5VL7S+FW6+oeTbBd
M0XZcBYy+gHkA1qPTB4+7Xgm3QfxwBd0W6LWYE7p8pH+iU1D39xzw7qZ0CH/9WUt
aEAIv7rarNJBwyvTwhIjWabOkI5QLzkfvtB52PRjID8qU712GQVp20wGMBETGBaV
L5u8468b282x0sqDfIsBQi+a4/9U/sPSGXKPF39XNcew2uhf/bKHArVYV/xyPV49
7PCrH7xrRhcWn3hDvxw+/0CZI3my5Qj7TdOB+A1XVu6BlPGe9Be0sZ7KXXJ6y4lZ
iVAAFVb3GSUaaHgZb0NMF5qVrQhfHi6iNbdr1iVR3hRuIFj+6h+t3Ycoge7cfFAg
1SFOoeybhe3/aYV8qnarQqFTOHt4sbCPD61GpisvrXPxcn0HPeyu6aB40tAieQWv
eP/1GSqlJIDb9uCmOYNrx/3jK7unOtyowFMRjOXqV4zkj4QBnTuM9ZU70q7UN288
wkZO50fE7VaCXjWVoqD0mb/lF15y75Xat6dosX/BWLWUx7jc2+tJpo2SHUCXQF5o
kJ4StHDTUmgl1hggSL8Wq+lg0CmxqivIF3kEV4xBBuTagpIPC8rQUvedHKBR2EZm
eUKLLKi8Dl4vX6HRlU8XN8ckgCnMp7MW/aCak5d7pYo9AMM8dvbk4O2G6w/UvIa2
SxxNDNIULejn9klqkz/wxXOmbZ0spn2DJ2fFfqd0rrQZuBz6c41lVnGtIyXpdMXy
vaD77EUUswl/NN5PyZ0BMBAgIpjPW5a8rjvPhiCiDIm/hu+/98jhQvVkSdLZIcje
RfE16lI9qZ1ia/HOkMyFSFGDZKcYxwsZWCkat2YO6U5psMkChWDCCSq3zsMT/opt
GgJ6vvZ/m+v1zvIxevlOXxsCMuPrn8lbCHEdX3TbEX3LegCRP592Kk6Z2IRy1IAO
VI151b2pS5WaEN7SX5DKdM7C9l1r8MpTXDpY+yp4PTasmqNovOcoNyWw/+pBbPFT
i2Pk3z+cC+cMq0NAVTB7f06/2vUdv4ULHOuCmqQgwwJOLjOX+5WwVJAzLt/JT8S5
RLA+WRbU0hX1nG5QyObMGh3TyDjY9N3vaTEs55pvFYOGPsPmpQbINiuilaueWi4V
Xc6Uhp4wiWTXKA4k3kDGLgg8pyGPHSzjg6bW+k3hvWDjrcJQeVCvyiZ49UKRanrS
9H+Rx+sOUxWdlpy6svELSXF9EFw5FiomDFTWtx02Fxi4xSwZ+WNo8Y9Ra3MWwzuT
v/8wBFdDetL9IN8wcBATpBL0aRQJZo9ynTZizwyX0dTVPZ1CLdxatEytj60XZ3il
8Vk931C5/M/79C1wq4G33tUoya2S5W3/16P9alcLLYaQsGhDWnsZ1iA/VEMIJW32
8kcY5wX2vr1VFn0khsQLfnysQbWDIDbjGYeG0YK71Ife5u8MVWVx1KJtEQtwewpN
Rf9VGoPGc61oAJrYAoQCW/RJgXYGuTnJOFtMoyTraefP8AGIIfo4Xg7OTQRRvKVR
kLCj7m7asHRcI8oy4DnlCefDs4ZxDr2v12SOLe3r6THb7ELk04AOG/0/+xjJfvt1
tFm19i2KEBnOK8GiACLnzfFoLCgPJBj+7qq1WAnAVu5vO/0xRoMu9Crpk8AcWulQ
AbR/29CAxp+qU55BbD8kus/ovNSgb/ApqAjiOdbwcV8Uz6e+h18AclUxTzS3/Jfk
skHvfu1IJ1FeeCeHFr6il/U1WapH5/pGDl3c43F+U5p5gaWdP4tCkThLwdcogm1y
+CdUbQipFZe2BubCWRWjC77pdQvVYuk8OEF+B9wQmyxBe5c1hNms2HxI/uJrmvTO
iNFqIIQYtdEO9qzlNIo0hEQlmnztpmk1WRx4UxcDSmaKTsW1CPyd9YtbJH1F5lmH
GHqNr+3KW/Pf4KWKkNFgxzyK5UaPZRwqMYmBZN1ZHxV3LnBvu/LtHeTDi8wwQ0Mp
ycENTerSrC15XUGX+5/vNeGTpOAgPyMAo/2slwnws/icwxnPPoCNE8EC3FdoI1Uq
7A5HfyhZrI4U0lemIRpQPwV0MhsIE8qkgjXreOy9ZVoMRTPQ1rm8TgdJOrYzN6j2
rPEEEQIiOzfXieJNik5IZawcxpjqbNpabgUOfh0fHBjATBwfZIL2qCmCOVwtsvaf
EEZWi0RCNF1AsYYtcPUzZw1DlbmkXaTVBGdid/jO64FqRSbmL3ceQ/umg9kf1/t1
OW4soSv0wbLBiW27WRIG3Dx0CkrLRbedhf0zl+E0EuZ9aPHZufHYA7i5/5ZoLhkU
gthvh5d0EcDD9WBhrUse0n4Y2abVMo7XtLLSaj7UJKLrr642jR2/eiSp2/sCHbvB
srJZnXtnV3GOqzuC9f1sNR3xsvhFkhM/TJRGI3S00h7BD5//9zm1kC4Px+sSjJAr
vxdwxGXLCqQm0YThC5dVczyWGtqUtsdU0dUeQViWz6U9HhP9bq/Ef5vzudoUWXCA
ozcb2WZQ9Icl0J9y9eQ5CB/6Q1qzp0iU0AQXczpeAEqzME0IDzb3QxgStenu9H07
LJssdvsZzwCNvq0oubLUi6bQgfpp7vi8r+1N/Jl40TLUpzDS4OmERU+C0QcNeBzz
y8oGElMzgMMVv68UcOtEUwVGd/z3HQMTP0GaI8h25bNYcBcgokPm4VZJghjumw/1
atpM1nBCeH9xzLbDbnqj6Upp1iQm0lmouFH02ioYc4tBq6jPBzepg/hcLo3sNqda
UilK5m5uYgdWqKS4QcToYfa7azx86yjH/qCLCz3GmpeKvtTfatynL3crusE2zV3S
ps4/jjzSAMBOs6dYdfwHQtTySXIwVRLiD+z9ffF1niPqmj1KvC1JlwOwDQYYO5Os
cXNHUGVOPOksDzHGNWz87sj01u83FYf3AlKtTSbuzOSDH+eLpastc1ca0pb+woJv
b3Nb2zNcnts6Q3/TjddzLO3N6p7dap/668FEqyM/oDB+bW5T8LBZtM4f0ASd/Wwv
quR4+yh0afuoMtEYXVQklf4bjSFOus+lT0J3eVYK8Hd0N7v5tOmhVQEq2AnIatA7
W/zESZvLJe+SLsAe5V4EFilSE6HGJeozEBr7myB13G2ZfLTqSOfBvBDVnAh3jQ8l
W4aiLkpP8X58MGr/ARWX52xu4Uj/ercyPq4DHktBGZx3utmQbgBxKsaWfN6Dzfxt
vyzmZ0v8pbkt2j+5adh9OTlJqfgSkVjh66toli3JP1kYyRZY+kvqgbpNzhCltMLM
O43pxb3oaYHgv6ZH2Jo+ofxzbbKGGiu50Vld4dbS6wgAhjzrzBl6/KYbWOxbWWVP
AuAlB8zrnB5y+hfOS59MBqLaVy3dCRdnqBDrMLfsVH5Mw7GtZ5iTo9n5FZ7hjnLz
lgm2AxacLU7nlNUucpLdn9Gg98+fkHsU6xysJBSz/7NPZIGh1lYB5pEKwcVzmAT4
3qu097QYHelGGlAwOzVfjRYncECNDKRm/mGotE1RFTXjPKiZ8nWyMtFgKixEhBXL
dMPEVxqY4IknancPZQvssd4/j7/lIn/fVgu42tAQWLtZ7+aqHxc7bfXJ46DVZrAB
Ew2ESDpph2M7rSnRtgPR2edtWiMSj8HNGZuJC/Jxh938xcB1cyxELYxPthFnWgY0
aQza8pd6+lwb/ki6E3sGz1ZzzjSjoHAnTiKZN7exHGsQW5KvgeX8JX0wbBF22jbO
G+SkLevhsj0txoahdSWsEF9SnDsLpUxdpCb8JQpUPZLoX4svyEVIdBCmf2dIOWfK
3+6Nnh22jQ4AufMIQokkcO7bjflinTYfQl56+aT1yRga1SRycruvGAoIq2wb7vo1
oXM714xvF8+Qq08OpfZh5b1ZHxC/himOmov8cFNIWY7+bAY5I7PxCOZDvAZ6OWLI
Ic0qYbaQHhvoMGwXbVHm7Q6dd3drXtUU5WRSlxtFpmj59XftNtLxwIttORMZt2ec
JdtY9NuDSEFHuPSn04gYVz1O9ZBbXuDSAIS8qOYWWhhmex1rzihZdYG6GL/MyNAq
qWZQBHLewqcDS09neqHVg24+Tvb0MRMPqpOhg9DSwcyd6rUMIh4byaXAC6iO8eW3
x7DN3tO4ZI9dHpkFscKa6aK8Q+FDt4mLyXY1TzDb06MnhQBx8jIJkqCRaEYObvUb
zvqFdSpmHWfgnqbBKu7OopO+sIwhcHM2Q9a3bDl7E1X0ZbvXzxmZahohHAT80CBz
9so7AuyRhAdLZ7tjdHh6lLrZ4CZSnNrPI9kG3LWw9SjADBkgr0uVd5aBTHhDISam
9ZUR4x9MBNsLqkfHfXnii/tO4AmRGDoOJg2jJ2iADcoYma+CZEA7uJSTX4QMTglm
b4bH+hrvjjO3hAeKGDCfpt08tMS/w6JcyswHrPRur2G7xvXFbXPNbVF77YGiYKvB
Iv4zFOJLtVNm98l58baJt4e15o9tKy113c4NhmSH4WIS/3HmnzWMn2qKfMb4LD7j
BXvkcmbr+p5qQkMAu/cORFr6fvszvcTgjhHmzHPsY83jLBXj7lHkCPHMf8dZoEet
uOUqupN1jRx9JHx0nxos9Qb9HPHqtYTavtjlXl/TfsCiLgRbliq23LMEKZMTw3mP
i/UMRtVkcTX/7+Kl0r1fJUCviXxFX8lscBsaaJ7q0TPwL3tgDwixVRMuoBdi7kzf
nKgoSDhg2trUbSSD4+T15vL8LS6bVYQA4cmgf2ovb+I9yxhAG9TnieE4vQXtfgrN
A4pDl1UvJJwRWPiuXGxlpMvEVt8kY1cAw8Ih2iSQ6qiXelFmGxcypDnsFN+ALtvZ
IeWKqJkJg1dUCUV1+ivM9a2SXrAaMjDRYj3uBmcCe6RnzDC94xtxHRCpPWU9KEGw
o9To5CKxMwg8XRhHj+j5fRudtDEAaMXT0y9SkDnvWPDvpe6KB8iHD26afyBi34Mh
YzznDlY8WH+2qEsoUVKp0MZYQ7CH05ntMRSl6qjoaMXbtCCLAaNIFyPvpvKVuC7P
FSUclO6PM89sxBfgnRH2oWm2mJDhooA5RTgZ1XEwymxnwb+0uK9Fu7OeoGgPrtA9
yad9991QtTMqxNqsF+yTKhhuQr1nr89EVvajpHAaxWMeZekMUg05fAtuoP+LtlkV
BjiCT8Ysm7deERG1iH3T9lRFGzX634w8kZhAbc4s0mqQOXX2Ilsarb2yZyClzzaI
aWdTFDkFcIRQ2krpVdZuXEoNjp6Pwn1WWBiep/aXb7VQromE3iPo3wB91Qr7eh+t
USm9AEcqjMaXuLRYM6zPatGZtJ9krKo8nF5J23akBYdFCE2LBj/vk7maXez9mo+2
lRn0ZgC1STmNp7TD0eswmpBWKOS2Yvaqanp7GlyVPzFDK9aA185UhDPg+4SNBWL4
QoqsDgnrE9SoHKGrNSAGvdM1iLjccBTeIqRu6fdAdFrhiNIyNr5Z043rGQ9cDeDE
jQ6cYPRBjQu+bmqE5lMVtJr+IJMZiGRbxfCvmI5SWfXbVlg/zvsm3vXr8B3GXUcS
nCo+Oeq3+mlV+PqGZEdRKxXON4KQFMeZsiPZX97S0AYQlVz/z/ICUqkIEiHtJRN9
60zF0mm6UutUVgIOkouClmBkz1RNckGQ3O41ksrbhuOYF6nQu3a9xEy1WoP51xDX
/ITQsWSPkOq3GqN7K2ALbDnDAFDvdupDPAoKv8Pn4PjZ4Q9z8/sYKY6+uLCV4LsE
Htt+AjFH14G/+1j7A2kPnlDzTkihAdk1q7dp5LxhONH4DPBXY0L3rTHUImDLUv+4
tJDSjmiuuVIyvVegGlJs4NAM0kD6W+H9i2+XeBQlrL8WZZaQ2AzahSHxDFHwqsTK
0p9FaGFYWlXbCO8I/12h2zUJqM1QBpBVdtfJ7zaUoFAVGo+jRPN76ilsnf2Va29e
SBW1xv2R/Q2S4o9c+RMFSvLCeTKm83orPZ03DxFtsDxiSqVJJFAK52PT45/X60EB
CFOQj5bYY7y6+2jJKhetwCr3giCI0JICdAjF4B9t/zq1jEJPWyCcg/NfODb1e97Q
VWwvIV2xpfQBb6NfVODbvWXjdifIYaCfbO4uMDTisL5pO6vOdL22bBI2NSDkfzLa
1zfzieNQVdr6uhXNG4qowgarfW5f4VJSJS4U6SgVnLEZd+3rfxWS/Bywn5MejY9L
f8xO8nrzxcC6Gs6gZ9QbqfSbLbV4iqZiy3IScBFoT+cu0BYp0+J/TYufDWeA5gCO
KWDh2RhAzEdJDzLrafKW9kV+kKeyCmRrQH/9MS6TpnxmOKYvdif940dB6htfb16b
1dEzFBFA623wTQ6t+u0SX4LoFZo9ZecaAb/8A1NIcFuvz3+CkvXvLKS4jUprP3kP
EGdkyPJjDllroQQP9o8F+rRT/2TsRftFrUnDpSZhU1H2kg+oZuFAn7rLWEf+yii1
6jJjd6tm+y+4liB5QH7sO+IIE8LmjPGZl8sBOdDbW+XvUi/xr2E/6mfX2ookPxsw
MWkuGx+dEwhlrWPIKMgSjjFW/M9jRRz2KTprM9Ode66nRstgjBIE/5jmRfskBwyH
DM1nrdB01sKRPzOTF9FGw5ldhg/M7lv0X8nYIoarC6CjD+3AynTkISZ8rwaCLq4Q
M7/1Dpt5Qgo6dbQHKBspEqB/4/+gpZfluEgk+1FkL5M1i2I+iJ+4sO7/+jgnIZ0d
9m6XNejwGGW1ePN42gh1HSdK4HeYkzv3M0UuqcFr2CfGFH+vANG+aiwkSn6tVjfU
laT4SJZ2BjtsYhmP/my+XVTw2aFt2D6/onL6EPnAahCDqFkJ2Vl3JN7NlMK64+WZ
37TgI+IYWUa0omMFHyWiBfnjFvmRYfnEdGw2BSpipq6h17MVmPGZwZBrqGrOadyH
VYGedHLQKHxqhpnoJJQ1HwSR4xvekV0GAgajA1N+DwBk/c50qOTo812B0WeLkbmu
2JxE1oPsVvPr6j3Fn8yr6PbtbbXLuNwZ1dHgKEGJfCiGs0qKs9AmC7f5rzc3p1UM
by7X+oI1NAk51wd+4cf7emENKGsCMCucw7O6RcJU7Zuz9x1RYT6/91U+dS2rxs3o
MNfLd6OGk5ghL1ONJWKGPq/S52O3W6XMFnt9BjvYQn3I+2YhhiQsI/M+pC92M9dk
RqNJuGzytOfkp25GYwFpdIszfufOVoTvC5AUGEa9c03Mfx4PHsW7GLIZPczosTg1
JeIaR3O+M2uB78AWEkwRBjRvzIed3X5MOvBy98d2u5nDBD/lDdtGdB3JwTomjaAL
DIUBQt0wu9jCEhxcPfrPojzER1GcBGFF6w4SzkhgfD8FeQdbK1efXIpGGUrU+Utj
n1n6YIamNXQ6bvLv0fwdGZz0TV5Wcyzy1/YEFb12L9Sys7LVVDqSgYqJMfEoB36g
VcoVrok+GcpyT2p2HTSyju8V2pf4iJfXj9WJUQ2BK4gZtCBR5tiPFX8fUMthRAcm
+BuIIQAJgBGCLtkFR5hVSxgCi5XANyNgkkaFkzUzJ7eK9XBDgB0E/TOs0Mv0DhPQ
nvXgW+1tk4cZLbEs3nh5m7GLHb5n5WE/QJ6R9B32x3woGmLtp44qIM2kBaAg9hTG
TWE4RJxsPcx55xXCF87oIJ+VVtksbdUPdcJAh8TyNXgwsS5TCMHW9AMa/4Tkkv1Y
Vt2FuOidAUnEF1+B8Q7pL/YGqB3+GJCSdPsPZEC8+MfdVrsm+0qwKxQ+1mb82mzs
Mxfq3Qav4eRC2PEvm0Z3opD9217Pi0nLsHf9jMxy6/uqVCD8QFbZfWKBiPlXTxpn
Xr6cmZeggx+M/52Bwc3NWYI/IcbQDBeZup0c80xlo+m190Wl7t9zOgWauRx9hvRV
YYtKhrKFjoUCUoPkALcv6+zHbLsL32QFOFgJFt3KOaA3WXN4KRcC9F81cucO6Bde
0hZRvMA3MTCFlixZLLyaTWcXmPMlcffi5RXgHbdSX7kPXv+8x60mqu0h0Nc6cmEK
HgdLHVbVpD/uhHk3lIlySXVqwh534+r8Ymqrod5usjx8VcpRxdzb3Ua0vJ6EN8yq
rTVz127ITrf5o1sFdwe4jBuFiFZ+ekziaM5tuYRb0HWPbWe4x0kiz4PF/H1Y5Z3Y
wQuENcbwm9J5xvqrjQUbn2bF6YC+RNYWDz5zBUvTs6E/8HtRx7zeGGcRINn5ARFa
aPi0JZa8JncStQz1CIgCGLu6GAOWjCaevWaxrKNEXdFoXeKdGmBAFvZJVy1jX/XL
UToa0dDuKjFkiJ+EJ5mE6U3rmwK0f0rHCaAy6IEf2xZSiYnFD1g7OigZI+tCUk+V
jn0tvHoVfIuSzSd5jD9dxYlq1pdI+9JQBnE0sg8UfkVciJmPZ1B8PUWOcLi7oTRh
Fkn1qiJ16D2zlIHifoWDPOP+qLcXhK7yxv5hRlusZ7r5Lohr4JVXtX01bIZZftdk
ENIGMS0WoiFhc4wAwoPjAW+v24Lr2IfdPuTNV2xMt3qiFvQ6eB3QimlsFmMHWBlh
KW8OqGCHws6dj122wO2EB4cf9iOQW1c4MJucBZHSPzfk4HOM+gqMrgFhrPIediUl
shFR8Sk9kzeon/1Nw9wDIvxuvERVgDcs1Fu0Zal9CB64fJopk/MuNHrEvNWIFDKf
s8ZheahLmYCZzYhQ1ccEOruaLvld1V97MkKbu4/V1stVijDiS5AiaIOQ+w2oC+5+
88hbgPYeFruh9tD3XuKI+Bi6lDg4N4KVbjf9GdBmOe3lgkNsJ1q100wVhAflfEz5
0IuKv66rtkUs+erPo1Ks6TaffhADDviKHEy1qV+81Y8MIWjge/QkWTRndmSpTHAg
Z6rQ2apsDis0R8m5TFFOuGxUzOqdfTOykVUBGhgrNtkqohZ8FU8gEJJeepOUcnF4
gPiQr443VHoA9zx73ieDPX0FUtVkvtcHNrov+gbUnDuBkD2xepJb7+ypynCvfjR/
JXZW2JNCkGs73f7l00vDNvtT2O+QS2Q3LlVy5p7A9FQ1HMntsnyb7faEOaYXZAHx
TxU4Rqcf8Rj0OsPoUT/8bAuaUUuWqzR7TLwZhHzAW8NjsPK/2wVMPVo2nqRcN8nd
dsPe7EFr98PXdU96Ht0GrQQkiCDVkyriTxzmIG6tUZqEI/A5McM+1TEy4owDY0fC
6g8Bm0mlVUl443IuRTVUFVwhu4vHF2s3N1NL5GA/e5+XubMXBKAIw0qeaDTGDdUx
tzesQMokN3kMZozNjFaMtV838MN4zUiogq/qAuD5RLjch7BPGsl4JB2D7hgaU73h
rU81xNXxXvmq6cWU+hKfufmpTv4VaUI6+g+qqpw8v9zyOtcXrB6IQqTUNvhxrHO2
PaHNgHN6IXYqguw5Fx037vxuhXVm1Bc0RsvT6ef/Jkc5pIRBRRmQuplDM61KK5a4
eg3jlDSh9njKHJ6Evgb9qLP03UN/7bbn/uVg1mp7pJNgyRTtdVCm6VTN+USytPr8
Nnp3H8phvTdUXn3hEG86WB5zUATdoozxV3XLWFMn5hzOK4mBnctQefVIIvSBuLlv
cSSgMCqAjVjJoFxe1hn8fj+G8Mz5Mm99kDlqOygHSyDBLfMRnnnvGzUPbLccxv7v
gF7kuBw3bFDyhmRiKGuv58X8OFhGaNmGmcOhzfWPsTEzUGKGUAYoxAmftdpT99eD
VCUIXJbsWvXAqbo1pOe7X/jlwDj8bCW8Z7QhgTMv1gQhXkD2Qv1McxpVPEnOeZch
s+qPBb54RJeAmucJNeHrwhmzDvdDiTh/OlYjylzRwEcUxfr6vkkVuN66jn/578S9
tD2C/CD+Tz9EPp0KPNOCqS+iQhL57xuywl81kFmX3LG+juqb3DarX/RSjBtHJCHl
Lv/8J3JVnoY4f1tzj9XEPbjpW286uQHWfzsJzc7/XMO54WQp6AIjyPmd9RQnjtK/
3Xs9mn+XiFkPytDCdC6mNkonAy41kE4ssUPoXlhHZ7oWMrYROQRF6ArAX90G+5mZ
W9mw2LLCoyhG/RPb3qY23mXRmVD/DirH+uGdJjI2y6hKmTbF9JdOj6NBw0aDNDGU
wePRqCDLPgBq6cYa8zPARRxJ4lwphIgEFAsfG3+DHF6BFdBZK5tdhUyDe3NUQJgw
w1/UZuiGh/P0WOy3Rz1NyLucaLDPtVwRDvZMsUOVpkw+rhcugKaY+C8964W19BjV
pCa4TkIQee85v+57lahPbU5r9pGCBb14IScbm/8q5kogo9isnqXLu/5UjEgoGXKu
EY9lGo+tEWiYXC/5rVRbOafXk7+HzhVS4YKXyoKgZfOM8KbUQHonE9F+c1OcRWrP
HlTZJcSPwfQ+MF6Pz3gc++6mh/ifutBUpJiV+yZ8G8RCpQAPO7CXPLn7YgBjDLla
bfl5qBhxsaKaVcovMHthPyY3AcrqflPD3u5deCl3FSaLgeAt8CymGLA2Tof0cplz
8dfHOu7v7i71maCss0ZThyCKuguEFaIegSlZS/mcTwBgMyaNCl/MiK0J6cs1Y3wW
YV1ppUpifoLvmGZBTJ0gG1TmEk6VKHmnHJMLZ19sQ+9WxIAMGNJrpk6xJowoL01C
RdrWgVnQ+Gl5AIB8IDgxb4qqPkcm4QuXca6DfiKmylW+vz3X2rOsRBhAG6+GEVGT
GMbtyDw+ZkaC9HHeRpP4v7Ez9h1ZkKtqYn0emkgz/Sf73oMGjSNkkeYn/JisJBg8
wiBu0jYGHS+N/lKe0qoXYOEu8rtijkCTfxkBH2EH8hDZS6QIeaNt7G5VRmCgXP1c
gCS+90aH4i+jRQpsX5AVwzHlngDf+1RwJRZJml3PE6119i5gt9K3PcG+atMPQDg3
P1yeTnQ37rajspp03MP2CZoPhH+/Nz4KYmsC+1oP1CjYp65Dpbaihvh/yt6iL94p
BWtP1Po+glzsPvThMmKiMOJc0teyolCgwwr4uT2ApU61qDv+Sl4CVy3O5FN2PMFe
KEp9F+Nh6Y0j9slBGQ8M1Voc2j2+ica6OygTuVVbRS51Ahwtqd8XY+jIFVzQmcwI
UTKFB/pQRGvLw3bTwLFbIeogZYW0T8aPsBnB+4UwwnKHT//EYernkyCLo6YBM8Zw
64UStUlsGcBnUEEWdOKDSXjZPHg6uyF4J+wb114x6bxuTTkRLchrUuBenNNos8MQ
Ee0pboyESxZq/7/kp+HMZ7CZY1dLon7C6xljZij7MMeqtU6ndRzENZnAdb1Fa+MJ
n6PZiIjUDtqfAQDMgqZRnUsPVHoyVf9RpzGfNoHLCOfev2zlm48z5goYUJKTiFuX
1JSLX/M2v9cIfB5lJYJtX32Lt8ll4Up2D6SUAeNsUc1fglx3tAEKKf16g2yy+ocD
7QG0JoQ0zTrCOyhMNqP+xDPlR6has/DyUO7oiLmHnrA1/DSthE8REM1DQr64A6ej
JBPP66L8VDE4BDNIeTnUJZEAxzRP5QlsDon3s51oNFn4lkPC0Yxq53rlQrhR2Yfy
78tzysZqg1uLMI4iAxsXKzVk60EbczNjzoaX8dnUfjmG2KpU5i1fjaPvELKds+7k
qThYm5nsk9LZ2fh8dTF4nl4+osznIgVPOYVx7DXvpqVn0Ow+86mLodUSsYxaw7D1
/b5atHKRo7EIeyLHHrSkbcHAmygyfo2HHy9vWMCAR2SW3pLa8+aeA3uOuaCCjV7N
IDFdf9NTfs88ic8JRjUpgtwhqRpMe0wNeQCFVN2hdkPjb2lONp9Yp7hPR2U96abs
GZQQpSgJRdJwmNvVdr6C6N3lGZZ3LrlyKSQtU3LKrJJGMbJU7lNnSCDtlP1r5NDE
b1/bJ6PfmhI2iVJrBCbga+IGEAxb8nT23OsXdKXBe3RrnZWO2WS6zpTwICjOBJnm
uvjsKC6FMEoyhHfJiHiVkePCGoQcZuN165ArJfpBpLqc+KszQxyk2lG0vMdOBL3Q
2U5ndJZv1gvG25WhLpyfJJaZX+5vCW1FXQs2n2MpehOwNDta51FnTwob9EM/HAKa
RYbhEy3CF5L0s5G9Yi5r+vueKwsWpaKd38hMW2SHDwU43TOdrQx4Lm2Psvq2iC13
fCrqydKo5gVa7ZU9o99CQm87zU88Ou8NVKuKYxJI5JhLUc3gaG8EV62R6jVCiRFe
tInah3Ne8Ty48Gcwds9OLJnzpKF/xQW2+YZxn6EmwT1riffhFiazpEFkEDDCrSkq
MtdPGsHCDktcT3qYxM/OAVhcL57o9oHiVn7OMXWwPyEJuLd7QZu0yifPRartXqn3
FLq3CQbYgTLsmP9kGlzgQZw28sSCd4n9ETVwlHTe4f92hLTO2eebgr+MSPXsk96M
4D2b9RJefLthZ2AMS1zOnFbA/PYMStlC5TFx0oIw1EA7h14Kb3PlbuJGJ+KEN2ZW
gflyEa9IduBJLs9Vgy0UkXl65CiDBQCmOAPFJ/64le3FgzW6qttGSpw75RTsQKqE
Jj+QwxK8IRkH63iWsZ+5v9CzAYTwAJOJBtmQ6KxNVU2LHempQxvSZ2eNUhifxejQ
aNgkJ2wEl97FT/N5VWmKXAWENAnWXop28c7s8OQdA5rfU/c5+Iu7UcKgZfoJKf57
po8G1zXkYf9WzfzlrDQuPwsUN2Kjab1DBVmIA2/60KQVVQOhJt+IYewBwVG40CQ+
xDSR/gPb2p7ZwA5JA8NKj7qvjLmEODbmIZUrzQlDSx9SeCyymWU3HrMfaULnXNuI
8meG2T3YkKzqDSn3Hg6V/5stMIOGWETRaU9+rPXbpt9ft2+HaUHw59ev/Rc3iqF2
8scVkDSHvjPMbsqyDdR78UkZsHuBISQEADsbFBVtuGcwUFIIPCKSX1BQJX5hr3oG
NN4QmHyFpsnyOJ8kV54q8I2I7+f58OUlqA9zeuaPpVAme7B4BBp710JIhgfJIYN5
e0ro4f2OWu0E89ayUpY/T5Twp9OIM3wHjYbtx4IYlplJbmaWDQKUwyH1RNq55yHT
8cjIU7ST4NI/jzmt0Y/8sIJctJdGE+P+5mDqKudd9WzRH2eGTSMHruK09bOI4dx0
2Tr104fobYEYNKY/JLAUkSy/HMfts1/qbol0pHCrog6a8tN0HIGL8HGZnZPK6kmu
lu04OzId2CfKf/IBjDkZbuEKacSz+r8/4rD3Y7SaHDkkHZaP1/aGvGNh9sCklavV
eYpJpeFEc6Hl4sE5x3FX3hRgV6/LerWjqFFj+bttX3Tzt1fIXT3FyJrWRA7u/QaG
CbffNREX7YHtUCq0G4dkXDm23wPgCwASb0lOC5WTmcWskWmwTv1gA3Rj+R2tL5xH
tu/46K/6Fpulfok3AWZYHSpl8dFqQmI4Wj4SLn9dhM9He0oGza3zzVbDEjqt8e2t
3ZJk0yV/IkqaffIUHu1T5y1yW5A9sY1H/HLcT32AyNxMJkw7pcQ5sFYaFNxEEn3p
rlodDUxhVRjg1sB6/HyjykHfs8iCd1YFvBKI/aSl5ljBhE5nP1iYEfknCOX3F4eo
Mus0t+nTjTLTrzrh7hvYQEmxDhq/44EoUYTgGJw3crZIrxk0DgrwqSYbwPkDePgw
ur1wiFNFEc535Ih6DroyAYAyg2YBpYUBaSzd0nJzSD0vtu+g7bK7d+ra3JUBhQ6h
UpJZ8NcDo92q5AccwGrY7FelWn0PCcxogURmZlu5xO8MeIMxlRIMvwb87J7RcioC
DLjYyhbin+PSM93jvmhUR7Lt7gLxgzVHiP6E3GUzfjhMz8zYmWWeZDfPMHchBiBl
Yla+rSwx4z2hJECkc1jqghi7MMvPfxr0qVwfuafOc7pVsCvr8r17Rdt8IuLyAKUn
FzaNGOyOmHN6zUKM5SP3CSBwmWU5BZyAYC6dmPLrq6To/sXd2ltpPKtmOJMK7sZv
Y1L3xMEYvTJtJxM6m05fwsK3kNfNhqIvxw7ZVMcSEGdKEZtI5QrPqrmG0seiBhNl
ZLBzreDRN4BfsglWnAAx2cbuynh55HONppnYiVZYY1fwteWTn0OavIt5iXplo25t
R+PP/1vFGVcA11mOfWOzsYcgecWcUePygsz4LDwk9CA5kuVDXcLSAc0xJ3NDv1Sj
D8AvwqYxfcxkOHbuye6YD4N+OkYU0TEhzRptvDhfmmbQ8u6STsOlpqW2Yr+W1C7S
YdVULoQTOOb7egz5/a5DOLY4z39KzabL5Q44XOup3OkhRmV85hT9S1x7loFivMRH
FtpQj/Dq/p1Mm/Z3OvsXJrscnlx/NX5oSFtonzms/box/v44LQ/ekHpXfb4kOt93
z7wmwPnd0nmx3EZwkDp88BVnPY0G0MQmjJ1BGivGV6TRURkn46HWMcTwaR/YW/LD
X1MqA05tA3Bb6YCnv8IMJONzjR8pgRIDIStdiddfvhKDTkDWdg9JNT732PUbD/A2
O9+jjre1XYYIkB/Fm6eokewOEOGn+Sja9HWvXs6Lboxqn7geH31+fkojHrk90Ipc
Ig6sTQFaWMX3A60KDnQ0F6VOVTOJZGI3QJPlF69vWmJC/LW/8A6V2Kcgl6LRGPTu
hbARNMThX5JUlbVr24G9dmn73cRQTfZyYrEwgMD57AgQGC8UVK0jynoXIYREvdqj
HsYHmr9llNZ+E2H8Ql0O6hvRs67aTKugDx2rAQ/kn3WKaXfGdrclS5Qx7pW84sKw
CPMCD0re8cw4Mb6p7I2ZaW87OxIuvJEXzj9fCTEcHPa+RQYi1tKbKLNpDCGXL52t
swlwQKZO7p5m/kloRRILabccrQvoG39UYVtBkxBF2S5Avj2nFxLIUWb4E00bGc3x
/Xf/iLj2MmkWQqyLwN73JJh1zz6ihXSMaRvmX1gVy7AO/vP1i8ypxAEL9ObmGDHl
DIqjhAi5jfP5xZxJt6h9vcOT/F98DnLior+NSWNpKVMcBnV1UwJl1T6IxgNLkppI
weo5ImzP0FDgW38pR2LBObAA8YAEyyUlLzmAMehb8E5LPuXfWxADgfrHzxUZL5DT
fA5gOLEl51ZMBLPlxI66KNF8fxSS6CmkXjzadja3C1DESCd4zCjmCFVb6N0A6nFZ
q5nDay/KCMBZacgYAYJLAmapDxxioJoRbOjgrqiQYcxAKhGtzmPEur2eaoeO1CBg
lAPOSVZw6u85tKvIbrYEO+QL36Y7GrstxICcGY+RQEmxgcWXSsaaehYTs817R6+a
SMVH4DK33YBatepgfP0vNSU+FRB5a6lh7Ys8ry0mUhZrge3ZB5xK2MtxfOQzjZFr
bDAUFp0wmEHUJkZ9YYOQfosvbK15UVZ5jmb92KrElkNK6/479SH0hnQiHs5IV07r
v1fTOx47Jv+og3NGaHeh29P/4foUqOK/7s8ZvLnEqqfwULIw3j5xjFR2O6FhKSde
8GhyzwdIpUxaVEglT3Cfrp44cZOkZkxhU/HOFO54iw2bATvjDh5cd+v9iSQz5gvo
pkeIpnQjZY1eTmP/ixe9NlWpmummqlNz0qUBiHS+OcChH+wISj3CY2G3s5PL/bY4
qUITtjqIRZfCDLJB5fRDUljlrq7NorBNM7djcEX8U/weIoWrgxTU/72YQQgVWfnS
Z6nuprzw6uudrr9o8zBStY+iHVPvzP/VdpdDo82vKgewDToXYO3XxXsDmycP4QL/
mhvs0OzyIiMDZE78E54GL8WDXNPbueYBt/mxHrwRsAnKX1nx76MqVFnmVhbptkVb
7Dg9vPYdI5Q95BHSZmWJy9nm2XkWKhfwg4o7679ds+b+1a10g6osTShrKMjJxQi3
m0XxVvpjjEN0DVKh1KQj/6QZVwx44WcoDBwJN7Nyn2XvGX/exBcyobCN0+g50RiO
OQTCao6QaWNHOTqiCDdzaqHDoiRhUDt8hmNaoMxi7H2ZLUKjh1YfOCb1GMRg8hO5
bTJl4TFYxwsBSXaxJ0wIy4qESsOW+/GPb5//kEg/rgBOIqbqsjKQeNdMu/JeD9H5
c0K0onBZ6D+3x5M2Hqfi9Q6ihCKeoN2uWm6l3atDZLHDP/7fOyRaGOORBgMUCU6P
qAdB3Fx6wCxxHkl8jWXLDgWmtMOhvUjs2YqGQNoz7OZYrIFvt0qEifMb95DiLfUO
W0srPo2nxigWtNUQp/T4mt8CBvUn6c+KiNPU2pGkWmYcaBCQMA022MwbVYm6EFnB
TfGjjQ8o4Eq7TRbD3GEN8pzFZuf1AjM5K0/X6WlFH8hvR+wAolvGK9/LJIyvLH25
kRCsnH4VT+HmAXKvayOGfxWbBJuRI4FOSd/FPlokHy6PwmcROh0C0KDHfJCTxgNV
mmHITW+gmig2JSGtLmcI9ZqAb6xhowbAL9FQbslKziWSKqB1LgBgRaxtRkeHYgAJ
nlvnVaNOjAB2It1DxtqNpl5FFyGB3vcFs6HYmhnUp9zQXiYPjTeTKjlhJS19IK0E
TF9rzyfvzFp2YuRD6b9FrHYfyxxTjM9OTBnN06lBhUciTeDQOrym9gVTisKGYSIy
6VWSRLvQMqqaOodL9kMl4rJl+jBIlYsqbJyZY3E+ja55sim0qLf5reou2YnwItG2
/08gMZHRmbLf/klBJD/k8wuhoXr+L87ssuhpg0Hp0MVVBu/pDQ+Rcq89bMa5bqBq
5tU65E9Gj50ZYu0N/Xfbqnp2yKLvp5YZbvvKVPDF8c4LxikGFXwt6PZETsTcak2B
ptMxxi8Zh4uF41ZNkgOccdmw3WVoB/Cb3dKQPzNz2jGioORTboJAEG6Ums6VaME3
sIb8bBPwtTW8asu6Fs8JemV1y84tr3eMsc3JcSJVzIf2VTVYnICbMgJ6RCmOQAY3
E+GelMiHC0lpmysz+iP9NLVYLhRIJce92t7xahBJKzoxqVq0VBgunkuBE94qN1aK
YigXu1VFdeML7FS1Pjj10CdTOg4GsceWj0492k3dGLIv8l4dPHOujBTyW270qRP3
Xabe0j+LydpjLEHRJyK8lPyCNjFOurErsLO0OgWrQMXpn4HvAXyWQ6F54DrYHk+C
AwDDC4QBmZRzUzBD0UGzGsHku2VT9EeRMFbs2jGZcng9kxGMVemB1tnO8/Oo4XAv
GGNRw8YQHy3R5dHBWOMFFIVwzA8Br3tFwHiM3kqTTF1HJ6X7/cyuDZ0cM4yHv/W5
45/n7Y0BRHxL0dard1d9Es1hA05rfMgnBlHYLFMRhSFa8uRjtPfyJikGZxJfi+H9
8tk6kK96Y5oH3FgOQkURQtBWFFeqS9Yhdry1aQ3uC5kk2PO63DsSXAIWrudG41Ie
JyJGgAtigjg51mcFn5eIjpAOO8TzM3YroL7PyhAYy0BrWt0XKFK+T8OShW671JZv
9lERvePUK7xbudM01Bng7X1sKlnX0XJ+gybtmOruVaQEg0/BtTzZ8bUgr//Ml8TV
z3xPx4NbgjxivYg3Ag/2mQso3+Y64A7FRxJv8gUJgw3UZk06R2hkyiuiChLrdJnC
uBgQQ1YdiAJzje/Wvm0wK1X6Bt/ioOunVPDJ4ueTgT89WVUE1Z4W++W0sqq3JPlZ
kBfRK/4PAtcdY6GqQ/cJHAD97beekcIcLq0jaGDekisRI7BKzNvso+F41S+W7r/D
rXaEQLET360qzEO1/HHuw2AUK9mUDLswRaUoD4nJ4U/fn7xFlOwe+LpUCJhMn/UN
P2Alil9JtXh6YNveAwQC6dfKwj/S85UGi529+25EbX7ez8+6F3gjadnOgqQPo3Wn
AOETW9mtfaHLc9H5vmE3d99PuStzPnP1CvpNeDHGdq7ytxDaSuG5VzlMA8i7V6p2
3QFXzIT/oA4H0huRucG8+heTAcjV1qiusaZzFUjcIR83NS+JkvnJ7OVzoWx6ykKf
y5WN6vb5rnhgsM/CzqCyGBnC5mJDiu4EWQoNJdh5yTB/P4brCuV72XYeafhI9flh
fGsspUkGi6lBsG6RoSFFJWwnv5pJO/mbqi1DhUfg6vVq0f1zmW1ouaon08gd+XmT
+zdrVkIZkm+dYfD/xYQcYMNq5pyvZC64d2NRFW/FuO7RI2Xr1/USL0gX4I/8CYOo
3RHWDha/Cu6X3H5SOTLyGRwNmde9oRom69Ixh7yzGm+0lGGGaNVV8PXDSt14jFjo
UOfJ1+TUYLR5VMp+dsOa6ZihkpexcAu681jINrhuJlV26EZ+AYjU1ECNg4cB6jkG
h0oYxDLyoiGstIVUGBE/bW0wjT/azzLJN7cd/8YeURhXsml3YGrWv+mrIOfS7pva
N2oV9HuGvC1Ns/MPKkX7hmWANFufi5N1H2Zp9fYcD10q7Dbin1HegW556LkMmcqP
vmY/tUZQWARLz16oi7Uq4gucDRuxGvVBQlkMH0ahWgAuisBHsKtOpcRze2EAcL2a
cIvrq4K7g92VtLoz1EmqztUoCike9EELXlkUBQttLXN55lX9GpQxvmfkUVDpSF7C
b4NSItDIDi5Hz0ijYBAUgSm9EFzpsHaankMHyqKIeVEUs4B3UMw67dqAl0FaJUJk
WjeqytFMnhsMXU6Fi3mKDv23O6vAbG70rOYbzWATQU6ofAj+v4xcSXAt5E8oPe6Y
0wX7ODcJ9+3snaizyDulBtB5N7YRoag+Zvz+RyZLqftv0tQJBkRAI7spvRDfws+m
OVR8y5w7VhVLula8gB1PiE4Ngcfg46EB0gg6jNSw4GgneR/yoqysNbWb7rwq/MdI
4veq9xSKdtNs+x7R+auW+RusdGBVgr5FTttnyW+VDEvnFHQ99Ka4WNF7JZ6qEQhU
SMYfwUZ3W7kwaZOjNmvE9yFs8RAXSbVRThJTvQX517qmor7LvgLMmlCKrB/EREnI
VXXUwqOrKOntmQFDsVYjUJLhuW0aLDozvnUmFdSkG+nUFdsYIrw0DhdStv2vXJp+
pLFtJiNKDf/7Ynz2CoExSuejDdEpauLPRZeumXGuCXNy60mlBjVx6gspRqCNzK6t
Q9kI6Bx6+TgmyTYbNgtRvLHU5INb8Ldax5bsRIhWpniNRjyjyMEWzwfk1e0TBmW9
/xGbj8bcyQjrZQcmZyUvCdeg1eX8k56widA/Fu0RsuB1xnLytQS7fzE14tqN5CIF
Kc9fAI+rJgctuMi8rjecF+o6smo07sgSX6Vg2ZryrFyiwFxZla0v8GZiQuetfYZL
OVNbgboe1nvgfU2Ga3Fh+/Uf7Egdox5IyYGedwOCmo0vDoxA2rKjl5dSSAr2yvNp
iEwhgW7C/FS8W9DCcacCc9gf5GllDcM7kx/aQ1Slo1CtJ9IP1l3sxpJiYpx1JnIA
pR4aLIOdvqn+LjqBAXgi2K32T/Anrrz/neiOlnMgkCXuLN0HovJ0v2+S0HCNw5E0
9vzl9hYjPbdsYc7lvEtU9hRre5fLes88LlI3JpcqntD8S+X25s5QxNKqlxtXEj8A
/YgZN+kc88Bbl930S/DqrXkH5vsC3LG/UjiSAoljOjYp+OsZyXTaDuZvZI+W/0S/
WE/6XFqK/Lpx3VbkD1wgCsgPN6KdhAMg5BFrbfpGNbQU5+rEAQjs8wlNV4DIbKAC
TPZJIbbLwaxBaIVOwQM9xq8Y8HyDR4XLMKg41SOIBH4a+QcbbKM1YHI0BGTZHz7K
EklIgI2+inLcoI6Q3eIFOjqNa/5W/U1XfE3uHTaRLcCANgMLV3/eZIjxYuNfZAm4
3S6Tf8AL30voOeRq94LkT5S6vHp9F3YyNGxhLiDjr0cLZ34XmHm+zo9LeqNf9GVq
1ycnPgYR8Xoz0hm1veprxC+LFH6wRfNz60EY/Gh+6mS3JFpZJhkDQ5KA1DL7BepW
1s3vaGTSuXck2e7QHcfkVitm8HQHvbRXb/cJbLTNAWaQdW1jGL/ncDbn4XPHO6p2
Mvz0R3BgIoJgrZvtaNtjibnd/L1Fya5rlojJdxEJRY4y3rpuLtIkHemaPslKjmjL
fNGufgAveVNsnuZzv5xMs8VFBq5/Nrr906UVt4TaEoyYYXeM6pT2c8b9V9fxbSJ9
tlHG2Llfh0t4kA0LKxWzEu+bkR/BWc+bTksz4xl9vW77CArt+3hI0rwXvBwcUR88
wSV8RdKyIt1yOdvSKl99bAHuybqQEjsEC9Ey4hj+nS4Ys6kPSB72ABfdOGnPT6OI
tjYINyMvDonSxV4J+wIPziELUNaES3hr5pyooUqDtxEbqsk9w5uXXNtTXi1rYux0
QataWk0CyTJJr61cu4FCHau/vgj3Mm6CYxis+vU/nB/klkAd3RFFZUiftuXjhAUH
txiylN6I2CuL8fv6C4mAteOJzfdjLhKvIp6nfrpGkZHkojgc9oy+4HH0rP9le0Af
k88pQZdK8jhY6UkBIiCVNIuN2IDAiSv6VxaOPdWQo7O0Bu6pio4gHn6w9wFDR737
sQyFSZ7EFg1iiFBsvx0m/PDMHyZ9pMF/SECnNeQWr9GmTfc/B6fZ/fYZ6+qI09k7
WHtdey9scvIKs9300/VkOVD4a12ZjOJhU8co6Oi+uWi/ZzGtN3eGhI6CkLddG5sK
8FIURbyyaxf1rj5AY8np6QS5FrAH5sLgL2vBZbjQoidV6wEgmEa3NaMjz39HT3z9
PXsPf08nF8ztPIHpOz/tKkitGvBnCUwLxEQO9va97n4ADpV2gAojmPjOTK+M5RpF
N/TKPVOrucb37A75HNzrAQk00idtySwC4QGkFZx9XU42yh5rw3IdgyYtUrji55Xt
j5waY3wPi5DzRfRKA5E5OhHSjm80hUG0tx6DBonErqAuCq2CYZMXB0TFLkR9+RGF
nJJC74eJ3MXJI9b/sffREcNO+zjfWw0kQdSMqLo86Dt6F+vpCmyhYeitOvoe6l1r
oQ4GOac2sDg7ZajUsqorQz2m4KMbmnbc/3arB4AD/asHBtagTlul+VMee0amYvRU
6VubYwb6xYcfHeCLJ9+1aCq5oCiRSwZ5AtbS9S64Rq8dnA3HWEk25LIqaN3GooOC
kucvgiAjl2l+BPcZL61anKHrc3AyfIwfBgmaKegKD+9vNapvBlpRxhpecHhXD9Kr
qiIHoFkNNEjnZA1ri4GOtT9SQaVZ/JSVX/n9dB8XlUJIVyvOZnM/eS7iennuaAus
4FqYmt407RZ4JXvqCBXLk0OzUgBQtliEsevYFVkjdYR+uxVmZuBXFRup91JabnrP
ph2z0CyZ9Wt9C0BGi2ZrYo3surqlKqHefDYS+Nmu4e6y9/j3orVYSoo8IRJva5w3
ix2C1NQ6jZETqjRXNaxuG/BIJ+zXiEuTt5Den3z0tyUE26/NbbYR0+LqBbwpCsxf
+UD2jYP3YnC4GoerD927/Yjil3AGyJ2jTZSBBAtCBnxGfVlum0NZMMl0BK3hbjDO
DbydC+fQuQXkIg16gXBOfMhq+yrkhgewtUDL/QhV44fkbuJwge31sXva/69Axs5I
TGUiI5JN0emp//HPAfTA7CkLBCJbmSs72M43Q4l15BC85AM6Cb9HfDmx2cieIA/8
Nfx3TQmbqRQ/NI89kBwxJsHeLegvTyU5OZvoKg+JZYiLwM7xIipZ0iVarHVQsTg4
NyljzIek1Q5PSSr930UZP0D82Ujnteg4t076FGXz01pWz/8bQj6PEkALFl2d2u7V
PF2i5DKwDcXqK2RDEaFtDrRi6ORHYG0G+5UheTQL+BgmQgJTDSWnBdxy+5X0axt9
XJcVC6B5o8xkKmarnFeTeJAoO4HCIc7zPJs9k10LxndHiPRSpMTf77zPYRQgWf51
`protect END_PROTECTED
