`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A38JTV2yqP3WRZvp/NfytJL25FxQlNLSgRIjkgfYULIhEGDwzVsL1IpPNOA73UE1
QAHbePVBaJQ/TxdWkyyxZSGXNr5H75DoVb5Shb3y6/GvJNCapG6sUHca7SXr6H2O
qFQHR2r4tT67mCQK7Bcsnw/TFoJyeFWQgggLhQiu6YQpjEMmv6oI+OO9MbrgR6ar
v8xHBH+qGMttJbv6T8faBlz/cWbkZ87pU54NCfAselFR+O5oborUpGi76Ahd1PrD
rNyXxAvf1sEAPoG1+6+snuev4Ru/zh99ftXYC6/nd0UC5H5S/w9SlWQQi4fc7TkW
TZ7ZIFq7S5llWT67bwTRQFX/OMQAVJeWxpNumvJelS+0zH0y/jUHUf2W4NszQ4B7
OQRFzFRRiqB/gM7aeFRywWvxXXJq1Dp8++4PPkPjLgLWzsxHWtIFX5oObDUgvlPh
46dYDdya5KgOTgQAXbIDDFzt4KbAMqxtox57nRlZqFvoS2YbjL7pMOUPmVAt61cZ
6DRjQ/G4p2dy2plWCxojDZXaRP6gTHfqMWlSwyQnQNaMlxCw4KgMJt7htVUHspo1
SC5Jn3seMrZ7IZ9ego7Tk+vxckidUiS8zrKC6LfQZNj9XJU0pnwZmuBStNUYOPc8
AYnmIzFL5AOTKCcofzKKQ44mvmXLCn5OuBAHtjCzhijYqRQNsG2Z3ssJGuh8v9Mx
15IKElNSC0ri7sxCaL5CNWhMdYn13XoMdBYAsJRDkHgYnxCNpLWEcMSxGbFENViF
/An2wHhE4Le8zSdhHz09eX6LuNzOvdNztxvrD9ZnM2a5fBICpI9CWxNtJ2BXDv6v
OLMGXbvSDSkeJGLZE94thaJh67Gy3s88+dLhjjOo/++BMsSuGN6ZXp9BhCKJZrD2
cyDjtjgFUJIR/hxGAafcIsC/qJc6y0N+UjVp5KXyxAtvOoMAv7sVNXYKU7Rsnone
ycvEq6yAyV6dAjXDAg222ChOWulv95puGqiqrimKgb9xZrPg3WnkCE44F5DVpgpu
dQvSgphQav+VOQIgSgj8XEj0YzpMKEzFPrhyPG5V4Zk1w87heqNpKBecjaG9oi+e
qYNfJi8LzffYqOqLetayRnerEILONWaSK+WW19LTHGbD/0pEhKIK0wvf9Y4mJidk
cmJKxqXPYUxWM6JC3U+LstKAINAeBlli8JWF3mnNkc29NQUqf18J06mpRiUbPkNT
Co9YUrNEh4uDjNEpYdquWKaOPCkN69NOh0vdSYEsMprFrRsxssjj80fD7hupagpQ
9F6wotzWvEK0a406kdEuH48Wq4Qtelc9yYTD8vbWmBzc+v/YMWlc6FmRxBNQo5ho
mw2Gp++7Eu96NuiMZZ2RPCGkSlJ+hGaGnu+QStMEquKvig+uUEteBm4B+BLO2BPR
vIZJvdQvIuu46JL5cm2esACxWn8ZUuFRYeym8UVFNRqDlRaye5Uw0UIaefoN4atQ
CxoxbdSX8ACM9ouvMMHGQ/9mHy3O8cAN/0a1+JgLm7wQYpPv2oxQYnIQcg1Ii1I/
knQsU4DWvRFdoysQsPzOVKSxbxZXfjlOUJnvrfv7Gs+UzVQ8wIcpTh/RIDtbzFq2
domdZCF6mtiRk/yR2yDbJWNvVqF4d6T+jdr9MLa0D+L0jp1GcJWWKQrNnwg8Nzn4
UwczdPRWiPZhXIbBx++QaVgczP2Y7LiLHn8n56SCBb8uBfEqlEcpkg027MyNv1kX
`protect END_PROTECTED
