`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Sg53xO7Mt27JtCNqk5qCe4l9c6z0qc8f7iBg/Ta87ttgVPlgvKwA0THoKJUvlG9V
5fiyRuXgP6GIk1QXogdmZOvMnu45W2KFSYwnYPBkwNvYFrAQzmEr0NrIcvXVqZoE
bHEkMY90uVqIQw5pEzt/MsBu8VuRU0JF1B2nktFDemUl+cDgS4fDDIA63yowS2M3
qfusra02AI2Iq9rpUloo7IL+kDiB/HybCONgYkpB7QW0mTqQSw+Ql2SUaA4SbXnx
iLzPcYPYB1H1srgrXcUTZVgKULiCj8V8QsWypyhqp/MffNC+vP0iyST1u5BruY4g
rGcSInIBp0bRf4iX1/rTNRWRSnej4/+sW71IEcLyeV2pcbZJr9/uCe+jVa8G/uvn
OpHXtgY/am2iaS3vZPXoYoJx5uYSMRTn+3HRocWY8r8M0AeTRD0dRVyrETuKjwIa
hXCIcuWWbi2og8RlobGmJLk0iig2Cziv8KPfl0BBWUpEafOgRn2WpPQ35E2rwIrP
pTG7arao8BgkAZQ7bD0NhNVMII3jvRgCCgOPlZrCzjEwKINxEL87TVHKXC7YWWkr
vCATHtFAqSH6bjp59cFDCelBiz+N1XT3QHshN5KAU7hlFGQ2Lekp/qpKWm9+KQIl
35P3KBxUv09++uI7DSmM1Bxc9WnOHdiBQSqVAmATMg4Aed64jal+dF942RnfWcIk
+QoKN+Ge3dAWAMJrz0w1LBYSC0c7cBW2NGVSnQxOESLLjPpKySjbxCt780Enveam
7LlqaO3X8b94UtnGQWQ4RChCMwLMBbmPIZo+9KIqClIZCeJ93gKkma2WTGNP1RE1
7MnbaHPVM8MY3LOQDXvKNeCqZmJ9A3koS7M5d3BSJufUFgNO1+OnQv69BVoT7lYW
Sshc5OuHL+XFNz52VKSutsFmXjGUwmjmgJa3Ly4QBDX801lbrSnxvyir7qrki1bU
`protect END_PROTECTED
