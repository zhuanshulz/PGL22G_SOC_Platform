`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ljGeRGK4UjNEIaBX8AiD2qwQ8rgte8R8rr1OSqQjg3RA8uj9XQnVMCRuywKa2Hhz
sR/hDOQ1zLbqbJC3DX/hihbrBCpPqhy3fACUFml7YpcRV8FCnUsVUMlD0toCCEgn
uaoFpsnQLxWvsdgq5+7bmJLeKBru+DMo/T8GCIc+cvrrVFBV2kiMRUgp2P3XVMEg
tZ8sj/7kIJ2s3Rx++/1DYIcovb01zntNoiM/zYxYhE6FPE1lfnDCeXCkLNqhHm07
GYow01qyMQsi7n74Pek+je/BVaSihBCIVsLXeba+3H6VsUBL3Sj2ikyArYPrAwQt
Lv83y1kuNLdWnz7zHkDuaELHuZC7QyYa4z2tSWN74QTAKmfCJHtfZQ6MrgIk1CQT
1THIlafRsm0rKfRWGptNfQOykw+nhe4kYvO5bDLMNzWfuw8mZKWbrzdwSABsiTYg
+HI9p0c3RDueUxmH8wiAcs6jybYgn+iao5tKs6L8k0CYixSF+NtGpA6ya5im8IhQ
LHM0DlIooimqfadezTX2nT8U17kSkB2YM72K2wM+Vs1M4tBE/8Gx4O5pGjRHosSo
QGgjLNoQBn7yI36SeaiOf33ut4rv4fh5tbE0CqaG1mA+1k5EblM3Yqy+h/T6d3DM
NtLD16r4G3XwN2sg0NRfdovAsfbkepjNu1qhK94llIPQASlTPGnq6FXsco9x8DS9
LyeptRzdYvyZjT06eoJV+ZPNreGeKMxiA5vHry7FTNm7jR5JxMvtDvl7yh81avV7
nO7COZeturgQ/Q1Ou0tVFrzJzHJwRIfwPCKEWZI1eVU3YYzfDlk+WHq5CPVPILfR
cbkOsAnsAs/kFV+ZSuxG6i6TyvkEHYqVSCPOTedajok9L1SQi58d6FgwBeUZPwOx
XE4+Je60LK2z6kpWp0krfScohON4UwQN1R5g0+gPhbqlRdUssgG2RaoQy1vI5Yot
agqhJcc8dhZSukFAMozUoloObfhk/AWArSwQHgAfM5EJNKRTH7Qo1Xe0JSxQCZts
crkZzOEQwLUci4XcooHQvnhFVNRR/QEWmLAt7kb8kTYpRQR0WCtDVtOJrSx0VWIb
xdvTcQHoouP4xoVN86o/pP4/xJ5PIlevMPnO3oEbfGIPwjXPMi7M4sGd6TdTPpxE
h5G2tkGoIhQi0hm7xW3+mlD/pRJ0U03YJb7Caa6Znf5lyYx5Q/BsBKw+oklcVmP7
RiXQPfs6nW93KzG6tnMAfb0P7vruk8t06LZuPobdah0OEJUOr0HIpEdYXQ8VSVlo
uIopdNKjvNb3l5IujmjpmKUTshmanjL8kVh/KeGpbyMUjyODfYz8xA+b965KZ2GV
p1BnENEb1BHAiRRD8k7NJHJci9XaLhsYkveI9sYNlOcY8chNPKIa6cfQVVlFUh83
FZZnw6yaMHBYbyM+qK4EZ6wSwvd70ruYiqWmnRIHkOJ5ftMgP/znv0ySwtbvrmw6
ex+3g9VbNoxq3y2qvnlUWPAfIwKMGaojSwcsiguV5jxSLCs/zjnZaWToLJwcxdHL
lN7OfJwZu0qQM138zgqIsFQi9RdLy7kMUdpZ+2NwOqSMgz/mBdGeJGt9c96/Vr+B
LDgLhRVileD10u4rh2UnNFth8C+rBrrWCQ+lQnnxG5KSioQaNBLT1H3QWN1TFyKF
`protect END_PROTECTED
