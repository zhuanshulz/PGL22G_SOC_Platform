`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VY9TPWtk34OwRCi05oGClq3urNR2iFnFAIpC7IIr71a9XohJWxaHiK9RisTzQYB8
mLdGS2Yt+WX7NfW/jvVSAwdQ4mM/4jgr4I9bRt6gYsPRCfpj73G+IWDKtPP/GauF
epeo0QnZ2v1KdnEvBIgQOe2kjSqymc7ntkCga/tlWJ8p9jF2Jp7WraMi4TProkFS
vFWbebBi6lVxVgvSWR8H1MKDFHTsN6yut1PuVeY1z4txPsNdDueWkwWsLrixBKA/
Y/IHiOA0B46T0c8Q3wK4RilxV611Nv6uOGNWCh2I6vEJd7dgppOI66FQaot1P+ZB
iDb7lMzckmY6ZrFMP8XRdDHFTl1mYn2nEStQk/cqYUsTX1RZWzHinleEHfx9uZJQ
ZX4Xe9NJyZ31EKNV8/LqC99kygXBBC5jyUB9SFup8vw1CQ9F1QYgiRI2AQZpv66X
ND4HLH1YKX+ZlSIT++gK/dYCO3JJ+pjaWDaFIkD3b3544UXYOcQo4EAcVEHa594+
bwHw91IQnQtoQpoAjtpYu0AdMmNwcwg8E9/oJHM3vmejmeNlIsT20qK028Wb4/rf
LNABO5nIIBfmmrmMhJ6pS8Z0psrjJGyUfxZYUagtGeBYZPRUkdOwbDDRf8Q5lbbc
qdd4RiaWY/wuatBjwnnz2V9Ppkzxebf06ExEKwCuC7Wng9th6dGRDjoyGgrWF9+P
fUo2CHsYaw5EVTx14lx1PfZTXnTZRXd3hltAT0cdKNS7hlDcmB232g2PHgxg1OGy
T2rvptU5VRg7Kuzgi1rO0AHvXkTgp2ifoOG1UvtptfaWfnPG0aVB/oXuOqARw0/h
+UgK9JbzCHGEC2kDo3+imHi4Uqrbcmb95IAsG6jQfCAv1iF2JL3M6FEbeIYfA1Lc
d6Dlu6Q1OQUJBTD4QjAq+4i7gvSCXIHDeaKCHhk3R03oZCtCiV4LspXdNDWkrxdP
M/4ka+DbPgi7ydwKwXceBurgRzs0tp8p1N7W10Ntt32sx59MbILbYXc3I3qRsRNQ
8q/4sPd7nm4WKLi/vaii0TmtV7OWADoCbR2IZs3Vvs6vR/8U00Gf4gO1avLa97kw
MKqzDFyLSwHC9wQnzGCI6bfM44/FB0XO0Es5aBFmzS1L4WhpwWCvNfqA7ZiuOeIi
Mter8WjlxxlANMY0jbcwcpqaZch8lDbKC33mlSzpVEbGUfh18YygUWM781pC+6xQ
oDV68cGIpDDnKE1dgaqBLV2j+/auxtOt6ciJUIIo3Sp9DtEb5HDotfVCuBmsQl95
BwbgEgJP8EQQWkRGtC5y9yUWig/9Caa8/qcx3Zzgqc5YODgJGCELrxnNURrZPhDP
vvGgKVauTG3/QstdeZCz3SwI9UpaweI7Jiiqs0kxYJoyAdmJqRf/aGMv0mHrcWJe
FUywDow1RD82nRi4T+mXhWUgJvsojKlu4sD2tJ6ydXmNbcPb9J4wcIvtSVxPj0xH
GLM5JJpwu8r65nPbwOIy6VRxorMzJ9YbdLQvZXDcBmMvrCXTFS50L/6WXvBOhLwv
Zu48hLSVMTH/sdcsX3n3j5gVg5sXnRZux8Oh8DyHNbF9s9gZ+eYjqqdhq+aOZrcc
2HzfthRtq8yb66QjhAY0KVpW3nStehtPuVTMwcENJQUHpuySAH5lckMFkFOr2cpo
TyKBmY6PwexFFoXn2thu8a4vz2VHGO7CcH1N7p6ScqZ1jaxHmUHHWMiPZCyOXe2h
SkyuffM/WZao+p8rIsXLJ07dtHKH8bhDqD99AbXcevuytPlq+C5/O0TeccRhW0jd
TWyaE51iTyv8tC13YsdWg43Uku9pKY4N1GqPFCR0+FLedGio0rE4YsYTkRrICQM3
0xDOGAXay1MtYiUks32qcY5e/7nUePvMahfinUvAGiZvAFWC5eFFrNLZFKDyXHm3
6Ra9xsC0Uwrqtp2hASBtHRQ62pNP9f9tLRfRVWxUcjvc0QX0baZy0JumYtxNHYOI
rofpJT58ARrBRYJj+3OnxsDLuvkAlqG6sYbY7JEU5h+p+XU2GF7TfTpAOkw3UsDA
bZu72RDdFFaD7KKaylJ2igeYwFoeoHtNCNWdW8EcbHLTX3KZKuLjCcWDak8Mux4O
ok88DE/R/3LuywxFzAIyWwUHcmoFsbIZvy9sO1HbCVle6QBiLfUKrNmTpPdrPAvp
DxZtWqFDIV5A11hsI5OEOzQLsTr1uQQKf2vz6Jxm4cNLpTztprb7TOYLakKpm056
PYBGoPf3D+g8iRPCfSCX8FYAA4GvMQePW2tASvux+ek7K0xb5bDVnNGex1NLlL3L
9JgyEMVLR6b1D2e8ILcPQ5XJeBdlRy7Y81ML3H4VDgwzFkqFzcVjHMi7lYcNz0sD
5GQpxA1VSQoVDaeTegXFTOmUj+fQTGByiKe4RvCZHYaM4GchGW4cfnF+xsfkOJKA
yrAuKg+s4GqfmcfEldvhOzqhAv8mM13Ttmq3rSKzWOr5V/dkIy76PTxQcoEDHxsx
z1t2seWYR0o17llqvh5mEAVfTqJCYr3fmOTAJ8q9MNsxrga7wIEJZH5fVG6UYoja
pDiDHbf1d+otQyDoxtuXW0Z/RDcwONBhEwdKD4kjVaGM/YUNgzzVWXzVY2BWXwVv
KOUMkCnTs7tS6NkHEyxFCkI8EkeNQpuF+LDKd/FZBUq/hmOR+c4ucf0txa28momu
/2o2jRSEa4H4skyi20i89j3gde5CRfMxCUv8gIzWFTGbCF0oYD+srbe/ZB1m/MoG
t+4k2dt+MmhLj0NwrNVA4aOVbEnm61K+cYEvqDPXZVTXpvx9ZaMRcmQSzVSNMQ/X
Ytsr1Off2KqAO7n1JQ6AS4Ecm+yJio3p3o48UmK5gmOy4DLS9pyQnMsgEEiaeub3
xjnKjIELAKk2ymT0MwSAC5mwnFZXHAnlkykI2s0++JgENWEnDsggG6NE6OzKKiDL
zOQUyaRulekuNgNX3PCpFapAlSeR3A2NUOnWKefuU6DiCKnPyqLyGofnPmkcaXl9
SxTGYM6Ih8ysS/h2ziKVHcF0Qiwgxfog3LCWZxmMmaSCtdsrDE7CiyL/57s2sEht
J7jM96i4YZB0R6uCj4N3WUO1QA1W/RFRgXfp3Qt8OBbLYuqXEfJHQPdPoAjtbX1k
jEScWPtTvVdA/YWkzU+zaGX55hAZ7HbMYX7wlqTnlES/z9gT9dckXJBqCs/KzktL
Ylefd+AnvXtD4Y/Tm4i6B8NjLtqX7AQuvT+90pCXuFffqaVlYwlEIjdnamHvadpQ
+cicEU907XCo+H/KMMWZsk2Lw5tl9ftOqt7c0bqjWzybwbNA+6Y9ZqREMbOMBbQh
4CtVTVBSHnDEkGx2cMJnzICVV7FazsuMf6tD2devl3OovNHrPfSgOq8QhR6k8wXK
cuqN7+QerV3h0tlpn4QPDULiRzXXHI0VKDddXRIBmf3WQJe1IqpY24zl4okNVX5f
rCckcyKkNeQ+c47OLOEpLN/aspZh6gjsMxzwHD4rev5WPT6VtKfh+l8CcKE1en3l
OEKnZ8cGk7OXdL6GHj1+vh1v7T9Ry/bQQy+ayJQf/mFlAG4lYAqa+EK3xB0YM7IP
Fj8s+HOA8jx5uVmG5++l1w==
`protect END_PROTECTED
