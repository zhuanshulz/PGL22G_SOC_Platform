`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
izC4Vs3xCLMJd3gHsUFUtNk3MfHczP2TTNQQIljTIUpfF1Fcvfahj+wyMHtpIqz6
QfDVJ02M7iuq00geD0dzcUfKwb6O03mTnczOKxcbJ/qJiDSVyES3fDVSRctG3OPq
y39Lbodx6EkN0y3BPjGFRFUY5Dxe6ceXQ6GWHTkyQnAkP1apWmK363QdtmqGE9UQ
w5jvNONx+pHclF+R5fQMdrnFw/ttfmbU216Zbgoxgub+uP2aSmSrHPdL4AQmftFL
w6H6Ixxp7muK97ptX/g1O2VusMctsKpwcAKZtgmpSvcRfaFdqcA9u4j0jObH1N/c
ZclXcZp+YQtM/q+PuBXOEMFMs4POR5K483IVqKbC3gbcJCMof9jacBJT3FvbMKZ7
ACCgg2BA4FJFXcvHxsWOvywGN2mnOsCsVBFsN2R779V3oucAUXxFjEMTIDqGwv1R
EiUWv+MUxwi6jqpzSExesgHxaLJJfMG/fyftEccJh+3la85uhn7OYS09vm53VNDq
WNeu4yUtdaK4ommb+hcLceYrD0okCYCu0zG+vmW2Ul+0I9gdZtURmjnx0THzFVS1
n8HQISoDPnCV2YlVW7Wsv0VtYpCZ9BM4H+hiRdAh3rIrLjc2Lhw+Xl/Ilmlv2+rQ
AspJZm+0+a9L6P0uWs3wRvNQs56KF4HedJ0Hmo+rrEDc2A7kEbU1gGVj0hN4zGp1
wh26yDCh5/N68kKuOvOxbb5x+MlWoYGdWxfzLTdPZkPe15nYwpf/eunYtLYzWCmx
A7wKtD1batJS2wzmB8MNOLITY39TnXWXu3uvKgrpTZv7TIccPpsQ1hHFdlXMNX0K
CtsbB5/MbLSeqB+El1EfDUHIohDOx5j19GZZS9trA6gVXyQE0B/s2OAg7TCdTusp
O0iPC7mHVRkQafL8UewqAmBwnY8KEFb4qg9E1SYEz8q/d28XcXSJmcHWfUKHH/gH
bKRuWxn/uvLe1kZlqfzVeEdP6SIZz3W/VPPkgwNQBaODnloAga4PalBtSWdlRUzy
1JfF9fsuLGP0qFFyL4E+L/AfPJW2meofBnwAZlj8W6/312mZAVcj/xChxcT1AcUa
EHveN9617uPcCDC7ANzCAMeDMYZR/Jf7PNOF94CRVYLZCjBmzZKUvHcPi7YfKvLd
eHHIvcKHMHemPASUGL9vOr5asiBAkOww1N8eLCWZl40=
`protect END_PROTECTED
