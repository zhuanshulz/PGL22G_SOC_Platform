`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZHPMOpAs7cwmqPMEbRERg4NYqvP/VbkaxAQZ0ODbkWgGl2rN3+KfOgS01qHUya7S
c/8ZtY0te4u/0TOpAss8rGufQPuOSDzOsarv979wHzF2X3T3c87OV2MwHsV2JuB2
q7N6QfAT0KkWhjRIr3N/6+HQ4wJacMzRWoCrQAEYBj+6XmKotgy4LwSMkWP++7c5
QTTzZXogRD+faOj3Ih4jKL77alSPgBfLRvZsJSx87VpjmHaWq7bmKTL/oriScic/
fJlX58ewoDzmcXH8TeeByAsz/dZVQeeCfxn6mb0NeLFHjXOlPq0aaB+7hOcWTSuI
LSa/HZrsR+CO3ZexPy5PqqjPV7ygGpz1YwX1xu1OwC1NMKG8lJCNmHHIjYG/BJ24
0cyIEygJBexs6hkvE0Ri1bRIvXqkmU46foKLHgB4h1QLLgbGUOA6YgijTVtXd9B/
yFlZP7qF8XZq+c8xVZeR+FrxR/eaHzFTCjwPWTgktL7RlBrAqQttWaacIIm1fQHx
Uyu/ehFTZzAU2dMuk2V1nU+m9vc6Ca1jdHxBky4BSl+mG2AuLINAB2kAg2S/zRur
WNwoay2PPS6q+EY43Nww3VTOV7JCSwsyLziKClwAkjsjXipVgust9R0psnFwza1x
2mjAOy5nPtKY6nVtBlcpuhRn2KnlIy6DpqCNNX0qYsz5F3s+2wbqhfMejLNzeuyi
FeC5Jr+84BNRaflPYBvKoAM1cc2mnfokt9wzU9FgPq2ixa+EWvnVhcyLNoDQPOYU
DUYkfEZn9/POt0x4YJmZO/0zkJ8eX2LCySwlh3URLwG8g8fWsUM6gvAqAy1PzN+J
7kBqZJ6oNbzlYNPO4yaNvrLPeLxdoYjTmm6YyPiQCjj8k718KRHlb3DFZGS/dAsL
GvjtD5iReypyHG5zYzTvVJXvsTaci9HOePGwSKogHrnZxS07r1gbIQwMmRvoUe+s
D9VdL/bLwdABnzX7ZE4gEYhCPxluFu2PoQN0IvbHjGAspzmZuNr16b9tC4hl28ph
IXWjN55+eeaRxZi5DALuI0qvMz9S7lmZpDzjGsQxqdCFYN4lSmwJKjgGYe5R7k5l
d9e0jcgES5wjBaV4GfJuR3rGOo1RxXeeP51iViwG59LDQujBAY2xPbRt8LKEanNG
4aCLFg+GCuveL75lt5JaJ/NL9uOS4QV7X441nsEQNVeZOYlr0s/y7HCVhs8cQTG9
mTGbJ5kFhR3vmf4IJMns3EHF/37YYU+7TtEhZvnXdrorCJa2WaH1AQZQ1032QRkk
iL01TcloRrIqLgiTWPmeQuR9b8eDSj7x+B5diRzSYazj0z43+wl0Y+eOfshp4Zcq
zPY8U+1Lhhs7J5VKDlgdKciF7X7aoiOC0juCaJdxddiTaPXe1B5mBggLs+6BV7RV
u3v3sqO604hCfpZhFTxYD4y5OaWGpwuhNUMkxiPySpBwLMcZ9E2AjW+vyF1t0VuV
pMAFQheoklBTpyaxcP4AAHKoHjhS+7BH9odIfuGO9GLV+vUxPfLkMb8LFTumoe1b
OlUryg/GammQr1kR+eSyW+Yp0d6tPkVBzTZ+1E0Un0msNKbJIMPaN/cz5psBspqC
T0Ijou1+mvJ+AALjl/0b3cL28AUuuIMV9Z17WJVz/BzdaF7+ld3+4cr0YFiIdBuu
3arq8KPM8zdujHEU7E41XKrQDePXV3CYn7oLXQ+3TLNiPJEY3RVVhCWtjMWHHQnB
RDu+NtyzcPMkKh2u7HsOkZpDvRurS0fnLMVEzAPncGVWACo5koJQHAjRwvNFBZGe
TPN+Md6xAfIq1uKAl9qIEWdYAh6GPHCj+5BXq8Fuq0a5if8sGZGAyyLgCmGHMBv9
UgaqaARBbORsc3va8W5K/w==
`protect END_PROTECTED
