`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6FTD8YcXBFLHN2mMHS3oSEv/6I+fu0ITGa5+LIsy2dV3bRLWj3XhVaUCVAHLdVTo
doXpfixN9/asuRs7FcINeTcvlIUHo+FERlNKo4SRg377O+yl8n8yTmTA91XKmfy0
ghy56Jwho54hX/tCIWOOO3YYzdpyh3al7wTjGsJDh75BhWc/t2sTyb3BNTPE9OhZ
BxCVLziYnsLdmL+YrutFYsDTa3FuispO7WRYCScJCnAhgDHpRN6Cuwu0a4a2EPVK
R71dkz1nCzcrO+pIofrC7b0mPn8xHThUqZDQ/wppRRLQT2O5N1TAtylOT94zAzfR
IlqlKLSsvv8v1PaBU7Fvb3wTGbTCW7WacFu3HXM6oiL8A9x9TNxRyAr4zm+prDkR
hGVzuIufph9QyxEQyV7hSpn6X05ZQeVD2wY98eimn7ApJlhbLazwDXuSHKC8m5G0
a1XzVeO8rm9lA4cJiGpLzvngBMeYohEAtTVeq+zPY+4qRkreW/5Ll+hgiO9wH0Ls
LCLTuwyeRuflL2auGtKWigQ9KCb2zBA82OOUHaPfA9o=
`protect END_PROTECTED
