`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l7iU3WWH+heaOjNMBPuJwMsl/gg1f/Pf1TNNHUwutqRmjuQ0zstUZaPLv6X1eOrQ
SKnyq83nE5lnq2D1UvI/CXF0WkDu43EhKbYN/zlAFJNsBIexBfovfR/+bKO1GEMt
Q529sAhqXCaqyWP0r//CCLopzqZ2tpefkmiRQLK3aHnCg4WJ91dRdHURIVOpF0O2
lrV0Q9v6MqOG6kL+5xcpp3+HlycXJUdhlttLFEDtaynFgQBYO1XWJdmbJv4CuI7C
MuPn4eP3DPPxbk874yllTlIgVnttV0FTS78rIEuBETHHsANO5FoJogZm2Xht763A
7C6OI5eX4BGSUGZMw+w8nFzZ4X8S1xBBV43ocd+/WQsEJkgbdsObP+r9GHrB00rq
COxBE/XhQ0cHTK19r2EzZSyKvklEVnk9A2exPZfey8+t2zSKZFdL5Hl3KFh4XkDg
zInDU9pCTLPxE2TMJEJy45rP2ROLJ12UR+hzwOwRgotKSprKGGeJbxd8Fho83qXF
0Q9K624GuQ1x1c6gam1uePeblmaZfbEmk3TzyT1+vvbT/eaLCEz8cytjh+UpWnP9
T6WNvn9dqG6ZQYdtoVloao2BK/kKoY/Z6ghFGPapBKccagUk2VzPZh+5taZ/ydZh
Mrtpgbo7M+lAJNobPt7sEF9AgIVZU803DW+P2oP3cs2JmFMhnSlSOP0amY2kRGrf
WZQXN5oQ+OWd1SlSZ5hNkZkj85Z0vLPp0WHkJBGcHUZemlab9HR8sxhz1Yck92wp
FcJ3b4nMrjFyWxBTAq8Xt0G7lRdz19LMmUkE8vakSjp6hvJcJEPJOv2VJ54olYET
WRedbNxPgkd+Z5C9dqgdShbBAsrmHSSI9fgXZrNy1dWvoh+mPmUun7wMIkxYBpHI
`protect END_PROTECTED
