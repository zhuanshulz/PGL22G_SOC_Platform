`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8RL2jCA+S53+YOlOOrgeux7bcT+6Ufl1XxpZOsL79NFIpUc3fcMMXRSah6NmSVGg
0v4aT8WrWDuuTy/5/R5cu+D2wele5wstemqU5u0HbUPropL51lH1eQL5QT874Bpa
u4gZ7+oFYrISJ/abN5sc56T9H7JSFYYLRF0ndj5OW3/51z/ur2Arj7BKM+4bh7nb
XEDNKNLWs6WkS1WY2Und+dSM7tlWPaQtLVPdO3LoXpH+zxHIqf0K05p5qdTTWCXi
CmXSpJx0CtvfchYJKTmSkmvdrqAKakvvsRZeAov8ArcKSHUQh/OYRa56A/JZd5rd
KBW435rRePRsyqkz3ISrexmZCzy4zfL5m2bD2lUyG8ipci5reBh7mhlFR1MeQ+Um
n07krGxRksy8N4k5MXtpN6YALQip+GDyhzZ5G2ichTHnfg+DFBGgoZj42uPzVdO/
EjpkFz9sR9L1mF/IEsYRlT8ldyeWWlmpTHEGymcY04nta4MZASpxlIEnNMBb32MQ
`protect END_PROTECTED
