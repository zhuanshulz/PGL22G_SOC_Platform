`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QD01yDMmQ1oYGVWWt/YlACqQeS+/pK0Wyc6X0Zii399iqBA6CrO7/3bm248meImr
rueyjyO8ZNjxyrKRc/G22nviCTAgDf57PWeocMdiWislGGz8Phqa68FW2crZsG1F
Zkz8WXTjIflTA6mgpKlUC+emCYaxed7XQZ8Ak+lODHTap+n7/pys2ISVDaQQGg1V
Vt8Wt7HQ4jdn7WUpstza4lYXBnBBJ0ZfJ/SIMo8gqkKamCuFtpDpcWJCch1SG90W
NpmVQ3UGhtWDTNwTdWIQHNDrUUHmPIyq0cF5SVPQbYA777Mv+JUu74bAN+VGHHp0
lpAm3SHFUrSiXZt5oaqJqvYMrDG3wwa2LlLeOzBfQRzLAlNc9np4c2+dsw3Bwkzn
X0gsxTe3Oiy4+Sdp1nRKlDDypZiWovBGMKKrsINOP3oY0CCwgptfQivjUTLnUT8Y
M9VX0ulfwEgSGj6gU0GJvfh8qZisYs4adAJZXsu8M2ho9W3FBmXavOoJXU1iBlQ/
Le03RzIniNganjG7QK++TdodZthHuD6mbZ32lIi5gSTvI8pZobley4HWTYDvEkKH
+3CXarGzQ4Iuer/UtZHmCw5ey3BEfLgUUgrkTgckaZIEv2MP2aU3OWTPHVJpI1/e
8hKzfTpodOgsRexqE37yXZv4R6a25SRz1YBe/4m+Pmg4h4ljPnGQxZI6sQzILz9R
hJ3ow357Wa7zELvUNNgmwxjbYhFCHeiL7uOVMiKbFtRnOR9YnoO8XKlWl5UNMjIh
K3oFDjQ0UN7CtEg2h2XsoScXgbuBwx8z7J/yIOiXL6dOFs/FsYHuVuD1c+Rg8u25
cBu+iRQ2MVAQ1AbM99szhUCqujOuiss0EGmtXTVWq3wfvMoXVnOcG7m1M5DUZjpc
RmluU80wfSBmVjyrYeLNcMd/E/A8D05ZyaS/qN8EGuYaNH+AfGN0pIx+jVuI54K0
Cyh/kTGUtxw2OAySO7n2nLt9oTxX33jcmqa0D4Z41+Sci9C333MwlYPDxGn2b2Fv
`protect END_PROTECTED
