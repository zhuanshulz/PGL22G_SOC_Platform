`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hwWaSsrr7cxfsS6Tdo3Yy/2pf37cA2j2Bgsf70ARbc820+FOnjxOFb2Km0Pivrye
tdjcorB5yXWRatHCO1UqnnUC5JM0glda6xTvpv8Hp0A255USy5Lb/q2tyk1cNJJN
ndmFA1KJ1M/93QxPcMCWnksp1c5XDaB2MsJ8VPUy48lSPV+lv19uyd7ueqntDu//
J1Q/O17rTlF9QyihVM5RA7eiJSH4S4x+m4gq8n/pQ880KZwDNvQt+tqylrlNxURE
+rmxMdnek6qlVAzjhwwft2yUw9rt0+VW8jyvXUTzEllRPsx5x3glTdcGP5mWTH6Z
Tx6A99BV5HcBm89anKOqASu/K8GjqfNVxvT44HIA8Me4eWTXeTONp8Lt9aA+JHkQ
+cKMcstSFJhk+2Qkr7MGx3VcYyW7CguLLM9VRi1TUwrGeM+ahWTdyn2cmTbxguR7
yNMVPlGNZ5EbF0J6hmWZ/gxiRlUyaoPVXNvOO7hlrnsi0s2hg7rJtDslsWBxStmj
ioOKQJE82wQHLoJ+Weyik1DR5cdg7nCb1SvyirBowF4syMyZcSA9N8gGguqDRCBK
MRZfXgniWhQya1jaI/L1FhCCrdqPmc6vv0ZQe4O3WHZIHPuvu4K2DGK2Zm7vpMYl
ZufXRwJrBEpP2RC6lpHCTA==
`protect END_PROTECTED
