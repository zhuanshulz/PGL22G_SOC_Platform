`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ecjGTKceVlhM5R7RBUb1CCff+DCjRx+GjeAtAnyNsMOCmUOmIEad6h5ToTIzzv5a
7mogahpWAb31W3+4zSVwyqhmhs+3LWMI8Nx2+A+8nbexpeuCKSi71wqmz6dYn7RW
arQf2gvaccVAtgJALb/hmVYEdT8ccfzdKFNemcPLKdwl9I6PxToFxnk611SPGOTA
xh3bxiNuDaJJb/ALx13FX/JdfJbZ/HTwQLb5Mo6sL4LvX1HSsI41YKn+C+xBIt9J
zFP3BcRgPfmBdJvagKsuWNV5PVPAVdCDRPCo3TYgiB6QDu75/63j1Mg4bjonmZqe
RgwUDXAyvp6cSv0saAPpoIdkL1IUfs4FqDBn+If5nz+YfFb9qu4AKhVY9bGCCy6A
UVOi4KObL/Tpw9lhaZIDTbh3aLSUAh5UHAjA2LwgaAQn/86yW8oJCc/40D872ZCz
rxAYhbnL/fnVcLFAp1t/mbqATi/ypkPShz3BvOBTBR04A+zGdyXscNGuLHWAa6s0
t7qba7rt3OvQFOVY7Gxp+g==
`protect END_PROTECTED
