`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3vvSbSb4f9R1sFl2YqwR6ThdSf4iCWwhEXHDu4KWGBY9FHeCeuj1GHoGsTdd2LwD
yr2ohUzUGq5vzprPBN603kvDQ9bs18HVv3R67VgYqvLxRGh4HgdxZ/MKRN81TF7B
30M2jpCszbo1PdEpszee+4oOdovezXdJ+il+EcnweHVusGgfK2ferqwuXRTEWNjh
on3Q0cSZazjuHSPPReODqVss/+2ImSGzKAcKPd9W4hu68jMlVQOD+AsCn7dfp8Hr
b99yp+WgW+LmWETZMJZVQ5Hih+aYqDEodUjYa1GFrfVbM5XKfGLggAwf79KMgQP4
Sris6DomejHBIqQew9k5iriJJ9loyhilUxAD/VZoEOplytJiq/SIFA1aMAgJds/B
dDdC3MgIbH0UtxdTc+zS/qJIOLAN7E2Lpuv/ygUgrUMx0jgnCJGxD9q39tX0rdlo
`protect END_PROTECTED
