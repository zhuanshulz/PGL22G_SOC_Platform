`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wU27FZBSuFaXLWXBzkV2FCrJkjbmcK7SydLE81zal3+y2S2twoF28IoT0VPCbq+J
B4OtWGApUNrO07vEwsMqg1Q00FF189V6DHbuydjlTAmIonCyvyx8vSYf1PQ1yHYI
Ex2NOPRfxTSQMRu5ZLlhZDWWYX2v8fpyqjeuhi0qvcP8hKoeKGbxi13mMZJuCpSW
ppXUqoss8ILYktIkddjEnMv8yKdla2YygLPzw+3Wwg7UDy/PDm/kX1XmcpEKaVxq
YMEVUTAZ2kQUZIf7JRDYJj9OnPpEOlXYQzVuf15kDGaIVVjt+A306vHOe9+5JA/j
kKy0QbBwMrPhNsdw0kab9cUaOoP0r2HQ3NVpbcGQ+2XgC3/mbFCmf7AxMuvqnb8d
IcwjmrbAltt9ImTLfharHfcSMuso8JUXds9DtN2YycbTPd08ZPq047sk2sCziie1
nay8GzDquzFNl2LVaNFVDdr5Oo5mHqnwZAlLvQfS4qbdIoqnOjkYqHYMU847Nrzf
/j98tD98s9Ly67mtWSIyBCyxwlTBvmDrldASVfMOBx/XYQ02kYcAh4DL2rJCA6w+
xy69jnBd5U1GercD7SCRGfWT4C5mg8q0FodzQIH2mffFECcfFOIhXomi2acxd5q7
h0SNgu6jE8kRMjnvlgQbUew/UPKkRSacH/uEiruG88ClsciJwEgeLy7Ang/y1laB
peq2B0dNS7dvswc/3HSZClQhN/GOdoNpdLX3fJBJojuKTqyu57nCr7RnSppKA0mK
3Zm5Tn4pl4o5jHC1dDhYQhd6bXC/vaVX+FnYNvDngj1dVizl8/J/fMQxZApsiUOK
3R3zt7gAQkKvstYQtxa1xM1Z1wCSti6bv+kpgPrAj2y5qELBQ2Oc6UTQnV3a/Q7t
guGBdB/k9sizGYfhJ/KIOs0BGr+lbQvXUVhv3qkgBNPXFoBt5Zmow7Dyb5utiKMf
IKNBeibM0EOcAYa744QuECXg3rL/21OIqpGfjYpswZQ3WJ34OhC6wcpb+cgKzVgo
pZyGgmIWVgsHENE8sRHOvZogvsHdr5hGPBwFODa4TqPt0rrJRx4pB5JMRT2bdkZj
BQ7kuLuugBgGCVWLIJPyS2ToiKDeso0gIGrPtl301HqThq8k/eXjujQg3XUYTH3v
FXIagKdYfBz2a3F9O1d9EzLVGnS1lrfs9ZqYpggGWA09QFubiKOjMWxlFDhqXe7y
gjQg3vg/w/l/oQL11aDdneXc9GJOAsBVo3WYdhjaD3fGLLujkE5FuokPs0ZKRW+9
gI79a6SO8nvjaCYio8K1ok0Lia4GoOyhVPskP9Tc+aVPsV6SOJWtzs1KLsJ1D/Ne
SKiCkWffKRV8Lbkjd/dlDD7Qa3Bvxs8YQjmFfffGxFk0PzxTy1TIlWKNksu2zdfq
ENsIujPPgnnnqXc4I7biq1TfitpJez2vRV6cYswxMzwr9t4/by2/+ZjNeAu5XSWR
W73BNv7gYDIQfG19awEufNH+rzaNxD0y2bN7QJkmlth3tl0AsjGi1k2yAM/K/aj6
kDRQaNDvFTiXuJHtLda++azAKlOrQPdytBffKGT3Cu6FztaPVyBXfKUu3CjoPLdj
QYyVjBZft2NBd0LFdq+lM797M00jn4xSLh/l25MPcRrNTTyqHGDDZutsQHxV1yxU
4y8lfX/zHBdui65bVdDjS33ZGj2f/qBduLHrn8Ri2cubMIm1b/b/VbKiW+KVi7++
ubtzzTIzSC/i8o3heT6q3q9BfQjzUp6676Ezr9+uZ4oRCPYD90srSrZnzvkGYgfA
BhPApgs8vphVu5vna0D1CNlIvytYOzV005YUb+18flsGUlvRcFgSu2814QuQcigX
PL16pEFSFpAexaa6CUyp3IKvubO9VxMIdKs+JJYBOHtr8M5rS+KhcYxkfDIFPHEN
NXB7M/ljKcWWL3Qhh21WFj/UH6XVFvzRJvx1hs+bbSVwSIuvfJC1b+4G5eliqiOp
AfAP77vJeUTgDEMSwgDagWlLsrZx7gwthKmhK3gjGb1VK/AqtLqCZf/bFGADFEiY
EIr8T7JP0NcXz1AxoCe/OYVKFn2FdAMQqh9owrkEcHDHkxqfM5MpimuOiakSC5f7
ExFTAmIYGE58EeItiTXPiaUE66B+dUFmNU45kNwfTUf/6vt52Vlav0ivXOJcG8aE
4iw+fOgKg/vQQcBPJyUx2RVTN54B3jINzqivLFnEJf6AYSo010gCTtqUbf20r1em
Xl+IrC/GEMxCu2GGVpQudCITU8sNO9AMcoKtyreh3kAgdA1uONAZYZrAu/mNeGQI
TMV5GhXF3EPLMm46BAEAUAXg7KgqTzFMZrCX4e5Btvp/5m7Q6d7QyzRX6z7G89Ge
1CBYEEoKkOTwEDjM/v606i2XI4RBO+b64WV8CM3DPHWMMEPJPe1/Sk7wv1MwainA
v6msXZOk06yBfu0KwrIbRwO7hl9E2DzMzfF3+FOiT+Y3Egwd+v0gTKZRuvfwfe04
Y7Nk4IP4M/sjtKavaIqXcGzYFkLGeO8EWnm27WzUjwbozoaLVypJAl/plMeGwf9h
2nkf/7hOlYbEJvQRtgaX3Cg++Fhj9mGC7SRAQsYIlwM2zJCzF+5Lg3o5lMYJUiVO
KQbj9Tjwd/l1VfnBmlAX35YDsov/D+kJPAKgwanUBndJTzwyw8uRcEDNiTfArHCU
J9Cuo5Q2Y9E+WPhE7LaEq9Hydrg+I3bI/gIkRXTh9fs=
`protect END_PROTECTED
