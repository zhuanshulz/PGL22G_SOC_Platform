`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WRv1NIlyD04KTuliS8gKmDHS0cX/CoBx2rStkjKgd6m4SWp3CqvFiDGPe73O0ROK
4FQbCb+OCf+Q/BMBI6ej7qu9qHHqUJfrQBKCUiFsydUow0rnReIJFI9Bu7dhhItc
Qlcx+5c62vPzpTcuq7e/Kc4XnNvNCwXoY+t7QK6q0dtN3463q0L1TLdV7A5MTjRr
KNrNz81EZyKcdYJdpJbNtfRYoWs3aCsIcc+0wUKlxjvDuUFxBzKbcDrYH0DRYt/C
fYIhs2anFqRwCEH1FyS0NT73yfD15Dx7DhSzFbQvGBF7lw0FJRA7bPTOGBJD9Bgv
OZKQKVEwZq3eHkevfm04+c0QUi79txge0Ttp95b2TPm+uDYCd8MeL+K93Crw2d9i
`protect END_PROTECTED
