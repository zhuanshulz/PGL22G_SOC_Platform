`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XJkOs87AZMnrDFpYODt2Y+xzmCCjAzxPbBP7+i7MFJxaW8lutxEwqzPoqoTRkZ6B
WygcX87viy3nI5i3nOq6QdFbwekqV/K1PQhbhIbmeN6TOfOg9u4ZrSMjQnHZyPO/
97KfuwWdGo2aWWqldWc7blxxjfWorUzzp6+UwlegvX9+AzGjoE1Dzc4vrTXLDkj1
8x4ttaIvNSXOL43p/cwNVI03cJtWdG3bsBY4DdaNsEPiPvzIt/VZ7z8cNxMtJFh9
IYLFMvnREGcZBfnSI9v/L1EKTY6tsT1W0sJ1473tGRJ51VfzXm30GQDyFxJv2jt6
ZW01giwAZiFnSI51dnxtT77QEvqHQnThLDjYE1YmKP4cJ1FnKpkR1ItkPMOdfp0d
`protect END_PROTECTED
