`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tYtctCeom4gvsSjmkc0S5NqzfWsWLsy/LCEM0ixoDQGfYwnIhD7HgVPCOISS1BjQ
TAorcdBQMet9778pztqvOKWyrFgzsOfcYrF4rdfsT1/hdd+63a9f0xA5dvBVuKKs
OBhSbGQ2iDpZJWYY/knZfodsV56WplAHN1GTdptyI0SJYuS4OSm56CGjfyGMUUV4
p57Afj2W54m7iyB+g+FUA59HL/mnj/yBVwPYghpbIUs0AFkOwfv98dM3R3QrrF45
2a749Q+Ae990NiavfltpjDBy3ivtQbBIvwgNXir8QWPfweZlaSpi+ZslHE/3t5c3
IciZ/y6JbFSvnAQV90FGZvAFaaCSJX/cNhXYi6XZyYPzvwRWMY1bZckKeELxW6hP
UnKeMSytBIHEmsDi6Cdgk2yKt1nSGRgG0iF5ZpazNyChl+/3p3zxNqzLiWysl0HI
/lHcprQX1Agut6GYIfxbRAKjNVahOXq7VtekjrKBvHVX6idq5nL+bOWLPqe3YN8D
jk8b/ejrAmEmqMs7dn3sv0vxeNOqT87NMdKlzPX4o2W0mkA9lm3FkYIrCub4oCaa
U9Qn4I/TaUNBGv6L+SMKwjh1isb9vuYenF7n8g80MZ5Wqp38NBImPpheYCWXaWWU
`protect END_PROTECTED
