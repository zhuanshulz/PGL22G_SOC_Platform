`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aXmSMsbgwrdVZAdN9dSap5boNx9lQnDyWlEkzephiW/DMs52DjkO3n/bbat5j3r+
+hMX/IlVEQQ1rYvEck+TV8t72pfDx+S//cHDuuwB98fxdhWtWbagPN1ceSClimr9
RFHmumuO1oD+0bZ78HW/bcIkuw3rVPbREjBifSr0euxy/GF75aFJ7PmkdklE2aLa
IiDyZt0OCos7VWB1ZMEvmgVHZG5GNKby18IeaJubtL/goUKvah1bbqcHC4XrnI/W
17Rii/7IX/JOmk8M/TDOIhqnIMz21Yx2QhTFupnRS7Viu7+fSgPGJCZH0J25I9BM
cD6NsE5VszAuyYwWw1p6x0uBVavKCk4Otn/jtyUKZJuV10nj8Ygaqx83r6lz8rdk
M92F/e3nyiDzjrihCvgycsOuhymdr9FGsKPpVGkiN6U=
`protect END_PROTECTED
