`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RSKZcTKLTNn2ixxsSu8D9v0WlHqZbhz5DhlNpWtHW+vkvQNP1YO5AdMFILv/56Ce
4EzCAr3IYf0DNS00ayhzCV4Ic3BdFCAjxUwIdRjnZ2q2XdmwU8N1QGa/2glLMXtf
JH1T3aLCciShe7e+JcYwvjlRqx71qf35pz5QYJqP2pOAkroiojG1nVIv8Rs6FwZb
6RmV0W9qVVoiRMMcjg0Xi/umgLJQsVgyVZDyyNVwBNQ3sGBljtrEezwvwYFCz1lL
mFWPo/lUu47x+XVvtIihaqfTF/VzGGCBaDLU0qlrnWKx4UrshfId/BbcK80sXzCA
1WahYEdtd7xPifMZ3AKB4Xd+h7cjacNKPwy37Oavmzp0LXIzXQ0Oi5aE8i8I7z14
qSnOONN7ME2Pk+Xnv5mObd0b9Lc39CQLoSmfRALucG+y2bTcoKK84EUmr+2EdVBG
`protect END_PROTECTED
