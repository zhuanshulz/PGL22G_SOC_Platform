`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5FInPjI64He72TiN/qe6sMezeiJAjlvefLjvnRWTbf0cCSIS4QfPpyaAsAPhAtGu
00zP8W4dVznwH3SB+L/cHpLYlnYGEEqcjZQFMHV+8NSGXeX8B+ODIohiD2GfdYdL
8aTN4zwRcQavI+qLqFs4DjA41Myx94gLLrW3v+Qa1IiyyHXbv3pkUAmfCrv4R44w
Jbuy7/t/127gh+rs7nHx+toBcC9zIFLIx/sqw1M7utKL3Mr5KWNZbC7ZkcbJvEkq
Z4CBXt7cShCne5d4vIb2bcglwyPz7aJ93b90vC/H2ZYe+NijsDNd13DcSE5F1ubk
eRx81zEoACF+QxWDsBYMHAyNb9DLW4CtciZoe5wBWg+UdVIFpd4BKq8yADCHIG3J
CcF60gE6O/CqeFsTno8Ht35ruwzlCTFfx3E5tepd6OBsLozgztR0DndI7EnvGGsB
CEqlnKTyuhFZWq/ng3nlzSo6ruY2ZmsKPzxE0O+aMJaUTpSa4tI6Rf1CTPMOUgQy
oauclFSvWSRC4wSQpUeGgdJb7lq6umnsMfvbNWN1hDpBEkRF0tNEwG1xpjRv+3iX
wunn03GRmgqSHaEBufQzQ4potcfymYlw158B0uzL0V4S4a9iU0ts4Tijk59kak8L
JhN0HpAeYE6u+EkIU4/c5VJ12GDbnGFMieg6BuZX7110qTYW0blzuQJQRgGIK4xY
ARJStzrdCda5gJ3BosWGz3kTNQoE0Ed7KsplDbVkYa6hE6jOFLzUpLBFAplNVaZX
VGd4smacPIj1viHujvI4ULfra8j0zOwk34xywzfzxEvHtQVz4fgKi3wOB7om8xs9
nWruHLATT85L5gB0N6/x60FsEXxSn9VU4acql5AoheJV6wvv9Pttafbkd/gA2YDT
zsW6W5q+2/9W4adt4KVvnqU+2a/pLUo7DRlKc4fsNvdLR3AAknSnE+wUQV+g4p2e
15WtkTXRyoe5jVKSskAYrLDa9nl/Tox438z6B8sN9HccvsZfTo6DN3uW18shAgmg
Ox9jF38whrDwi+HeJuQD62skUoB8moXcO+nvqyUJCn+NFh1WeazT0Mg+u7cUKha3
2YoIz6jHwdnjw5mE0f5ebsYXw5/UdT5zHIUATTDpP/ZvvqHs35cTBg7C+vyy1hBI
LjP6RkXggUOc786ZX9qJxucgyJsPWwVWesLDVVWAMRLhWrIJ94cHF/zz/KPUf5Rn
fEYlqMJ2ZceE3rNqnWzCSLhJhwdpfP+/6YNABR9J/8uNQ4533JMHFCymTFwtZsP0
U7+simWrkONSjInXTwJCVx+d9SyIlgS662eg43IlQT1Se+3E7UwoTbOo7+YVZbSx
26PWx4omzEDXM7a/1sxBnHOKpJWVa3CzXxLmG4cAwa6LT2sG8YCzsM9e+RFUL2ZS
Aw4DyuffSt18kyGbD4WUZw==
`protect END_PROTECTED
