`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/E1YwRJKzB56CmuoZ2IT/gzwJCNSubpmhUgq0sdCJreI67DPnwiZiOTMMwatzXhn
j9+ar2LIbh+pOvRCmakf+8i5nC3gFJNVk5W01PpbOJt3g0cXEkxVekvKGI65uaCX
EbcLkl9gw+2pIoLC5ktARV0kZ8ZGe++8mwuERW6O1/zqiNVxhNAFNVyEuzI5hK+K
9Joh/fttnNXsS0+DDfTai1bOeLhtqiMFnNAb97i3DSz8ZCvQFs625YoRI+89K++w
5kecGpOSS3Fb24RzZ+44CmXvCKgq6iGhIPwkKIAFahdt3c2EZku91vF1ORoEUUNp
FDTyJxnAYIXV2HJxPbjQh9yQ1+xVtd39RtlU/7kQ0MFSUo8JI9yGOg11rmBDAqbF
UStRulSBIr3M1+iElXe/wdyH97Vduh6cCpD926DSuOE0bLDi5kNgzbsoTKIMfDGP
I52QBwpowkABd7OY0Bnyyfh33r2UmU27tm3+SOlutb100yNT7365kyY55LDAqmFx
ltOFGyo8TdHJYGsVFlVdNWwd7FypGU6wYJkZNIIScJpMpZlium6yImw6fSHOHU8g
c6Z6u6nCiyXKD4mnIiSu+xZZc9A+PUVZAlV7gppdsd9iwmZcleCdpeELyRLJqhV/
5ZqFlnAyDSzQ843ITFdOmkslYkC0yISobx3LpwwJsbZkyxvT3yKFNCvdkH82gXnP
APU50EpRUIup+7QxfbQiJqxU4L8KEKLRUkM+GCVvtpv3LQPEPPX4q1ZT0E2fdPMn
9DBM5JgBg9+AiKJ6nrsN1GxDGSJWMfc/GGfdW8hy/uQuxjskJp6ZuQUWaHzHUoYO
VR0eQg+r/tIkVNrGxOvCZ1lS6B0qn8qWhiNKUtPQBQppZH7DqmG/gQid0qcMgCua
YRdLKBLsxDQP60D7PTcTzreJQqF+kUOduGgzY3KYLZVvNEV9l7wmpmPas4m6WzMw
XvFVTLu0pjeaCI2W2YxjEuIAeL7Rz/J4qw286Slfo8UtcS4JEyqAJ9Kdw8jiwWrn
pDYhg9XLXhB6Miu5G2K7HFZmspIklhOaDtXrKHXVGi4P1Iy26czzH6MW7OrIKbP2
ZNgl7mUjxGyCUTRPEY7RI0lcOJhmdICa9fGUOKf4MQ7jrEawZP/D9h52RtJqWZJQ
u+c4QZGk3Pvm8yiNJd8hIQXkphrT+WQQ7+oPdyRJYkb8Hv6szj9bmKJJ9bvLNC+P
dtYMUoUXy6jwhmZULZDVW3t862CFuSAzQ/zpb512d6iA22EAzxHltx8zfdcUIftR
637XeFd2tI6whASWf1jaTQtBaMwno3Bd5dmCCEBjGuTcBYxDsXu1u89aujsC5DCF
pg1qFLmvlKAkWQBCkv3CK6mLviId6IYn7a8mLAr0wmsrdoD18F5d0uUN4ttsTyd4
2T8fbKlypWq3/Q8iVC58lwR4KoKEPu0tGz5PxlrSc5whOJas84Gmhf21Wykmuch+
1zLzj5D8yOOBDHmBJi0xKuGC935/05BU/dOjK2BXp6yMyLZ4CYuRPf5Z35lZ8YWh
Tk65yZcOHjFPdbm/no35oOFb7fMojDQw2UpijkARnPW82xWglSE2K9RnbwFtGILE
PXnyjm4G3c2suP838UgP8ZoiUqgXx0HiRAwDK4i7cjBmYpoqfkP5t6ImuBbuZvk2
PC8/gUE8lYeeTSHGQ6bLviI5Z4J4ICCboOf5NpR6g2ztMaz3vv/SkrV8D7RxdYEd
RoAyDWGhL/4siwg+PDmQZDJeRr/Mf+KtF6kRfQCX9gLf3cDAM1D+4iQMHP0AzuMy
pt3iIJgTZ9ejkg3Vo4X1G5ofsZOSFXKMMgUWX6RFY0SZwS0uX8JwXWtokx2oUxFj
i6Z7F75T76/h872V0D/EHWSc0TAq5gsj12sq/oMO3ownWJj9sI4LqstjjG/rT25j
DS6FUzHPwJXl2TGcImgl3qk/EYlYmWZvPb09/7VL+4PnYlmfFJRO8n73QsDbGmJl
`protect END_PROTECTED
