`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EkVviOww0tvjIR+Z7pVuoYMz2Th1trmRPfpf5ddnT7cmzu8BURWWo9IZLyVGwBB2
iF+fC9bQYF9Fhj6R6Xg5ZdhpsbtOch2cOqE4L4K5Qa1yk7iCwDvrUcBoMlNC8Nn4
w5W/Lrzb94BlEAWY4RBsgW9FVulQ0Va5OSN80vvT49Qe4V9Mz8CiUbQ2unELNyeX
bKgnsJ69rK7o2cmoNaK900xlcWBLTt8vCGdQWo38XEu04O/IfrqmJtMGcZABDhsF
8lWAhHJfMFLg9oFQcVyOOY5oB1obBM71CAU326453wnkX5VbiAA7mQ2hFYHud6Qq
GV0XM4LavzDJjKd6HlknEekAhusRv6qJKXqTwnmrHHokQEfTGNJDDGSeae7DUaTW
WnGt5DP4JTdD6kmX5k/GtD3kNNNc9OI8Mwmtao1KP9Vr45moVchbublJhu+YA/s6
wDlG97h3wTcq64Csf+D4pW3vnIIMvAcdXsLMw2vZx5EhL/CEkafmddtuiU+k9h93
3VJL37DGL0Lv8MX4UV0SpxbZQX7Up+JnF7Kq2EgkZ+TwMDxydTiw2lnAgq7AFkDC
AJaUyA96M092HUJn4fxeSYJ938hwwQuSH8jISWKbjPRJN7fNN1STIQWc2GQFpd9s
b1McVGbvKAYuidjg6DOs6WiYCZ5KT4BzmpDtx01dPuyUEYjXwAVHptEYYd9Bi0Hr
sFcjzOZUMx5W1H1nJucpR3WxK71OGJ8J/844vUdJTZpWz2/jvdMTR+WcqGupqoqE
mllLyUhMHBnf94Ve5DgLJr8WaXaD382Wlp1lbUseCrVPYq0+RAohir7DXA+8FIvr
Xm2Q6AmyDh76giybhiwY0wpk9mv5Bo3Tui/UWzGT5U0MHd9k/kQ17hNX9EcJmtFH
nTpDtEsI2q7xLDDqYbYTbcLtpVXz2+1giaIn7nDuknd4sJbsWJnatUDYqfSfUmly
VbW9VRTw7Zm44aEg6k7Ta8sNV/sOj2aoXR0IqP9BvgDmyPfnqlmK9qS1Aw72y5Lh
mrDJF3KCPbEqCqhOUf24+GH0B0II+VEkMxtWDkBF018RR28Wi8gegi+XychE3Urn
`protect END_PROTECTED
