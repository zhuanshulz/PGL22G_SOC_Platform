`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1LHHUvMOAHTFitI1Vfayr5kqcBOdGRX/JNhgnHPIwOuHqrbPsL8Y0W8DCpzDjOpR
9LaaoGgKUt8rRlDUulFf0HaETAVo4EgI5cL4Dmh3eM3nZCa/l9tS5KvolOgFdQiu
te+EabL+8c+xIE45rjvyYqY0zNhT4gR8dzUgOfvVwLkl+InTO6vQN/OqlS5xxlbu
Xg4Xy/8nQNEzcmW7tnujQh8B2pDjyakp3Db1fvb8Wsg8v3GMBgGEZ3softYCpBxg
OPG5QcuWh0jsecccZu8FsHG3RIDHBrBULp6NqM0mJZUmguHWg59oxQqeKZWzORAl
NeiT88wzoxOTtPDxPnO0ZhHMcgi3+TIik+tp20REMuOE+i9D4+HqcWAvtQwRBD62
xPmF6hargFVroPS/SxIDoDHl4d1VUITwzQe3L0AB33qhHB0NCv/Ph4LpCCue2VLs
doOsnlbRxQoLIIrFlHTUG3VB/T25qVR3aNYq0ymm7Qaz1E7jNTpJYEgJPSeH3Mxa
xQVq2lfVqX7SZkmsBt59ZwvL7OLHmO3TkPfYnlakHmgh1mzGlLuF5jt5z2jdWGHg
nbXTDCQqlj3im7TdRthySYCBFiy2AG94WGu+pAVOATVm8RBup5aX8aTLpNYNHY+p
`protect END_PROTECTED
