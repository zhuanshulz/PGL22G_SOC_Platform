`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gSm1/V44mutPaUtDQGpzUdDr6o7GfZu6LtjZA888uLyhyL8Zh+WUuHL7UtjNVMz3
kd2f3UJpbbEFtj2SDezOnt0zhpK6BWEvB4nwnLYD2OsX7iYJ5ZQ1+H1ewzrqBMss
OGdP4J+PzhNGUNOmmPTk7083+tzOyGYfSIJE7UAeRpVbFpSoDIpCooEhuKpRSDh5
NE0izSXlIguE/mhEVEmJQMa/P/F448Srzi93KOgeL8esB8ri0LoK1vxEEg1BJGrD
OZ6X2b8h4Km+cqrMqQAOicFkn8ciOizf4Fht1oeS/u3zojFQLqTOtbuT6UTLWjmu
r/MAAelJk70pLrgCh47WJW0KtUMhE0j2oBhmxnNvSOTtYShzlJja4DXzKxwvENdv
RbuEiI2al2wgMOD2thotBTSxuIpwhxGiWq2eArcj6OKfA+1Ki/1/8OF8VHOs+pYX
wGbjWN+xVBnbFZw7+43LvNdgIT9OsGjyqb0CXQct4965Z7IOEFE5weliNhS47YSb
dS18uXLqfaWNDjigLW1WOjdecKSNZK/NobUvQ2lqpnv2KwO+55UOhcOX4LjCLeHy
jl6wmqQ7R9s7BUkMGXqc3UTZ9Zob7OlHaE6o5ry0Al1h/tuTyBU7Oy5B8XGpRN77
jn8+Z8xzUu8yW0RfhAy4ia/fq1SL8zuqf0su7iMV+XMw0XSpPVVKHkuap/7ig3sA
g/sdoBEmI5gLbadsjGhD1DQATxcpIcoWD7L5/iigYnEjZYDRaGDeJdxA5ADFt3Bg
TFyTURY8OGgs/UB5xdxgCNhwMz8feHBRjgHoQyPazsNsG/XXNBY2ZbSpCTeF4tci
9q9IsjqbhiO7gjS6njsZPQk4VPXLQ9OgFIecVlHiwBWLQiT4Y4SJoPTp9PlJPNqc
uXrgt6s3rd5PWyFdSi2+5+6W96XZLfRdi4zf7WO0Zzwxays7YiXauu/8abf5vrj7
kpCI2VzSpqAasibkwj3SOOnCSD9qQfKRn/mw5ET2bvXN+S0sng2AMtMN3m+4/Q5q
E+eif/Z93YBffO6MIENnLugCPbY1qXHcTMV2gdFstLU=
`protect END_PROTECTED
