`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q38QJqW/S+RCsdIejhTv2DS20Of+ZrEQnPtHL2pEGFpc+SIr17zNRFGSX8sCNUBa
Y7XHLmmGPViT90XhCoPZCN0UXegvy6unP0RDAAGSEnAMZCa3H2wIr7GmsqFF+DV7
ejMWM1uNt+7DtDxCW6dah3fckkMBx1h+erV5+jX+BUFfX7bGULUUuoA/1ZGEhe84
Spzw0QNPdOYcWrPWrdmrVQQ5qQSnbCUA/G5HGXUyirpztezHOl0TOT5x1bOR1XDE
8dc1MecXl+ivx9WPHdlSg606pocEJPTadCvU31g3P67P1+HdrV6STVJw6C02xUNr
H0IKESQ3MUsLXCo0u4E78NiVgOupuy5zr3ZgRz0vvuV6omawZjyAQfMAduU+eLR7
WtNzNLEX3jNlPk1BhK5kXQkChJ164fAMocx6CdgDzODz8GMNAbnwl4JG/VyfcRtW
GBa7fjsyLaKqwb/M22siZjc1ZPZ4Fb6ummh5nTl5y4OXDhRY3vDRl/4uwAK+VUU2
jjWsidIwzmlfGxcw/lwDqU9rYAbBxVfLQhfFbadkkD8g5f9J9DwmE984UPaIg50C
Rj6Cqj870I+aJthFPvW+2Lmk5wBJ11ByZTFfSlrFfmB3HT4qQ2/AMkabAW6IwZyx
2xCQnIS0amoVnmEn/o0f6uAip15LHKIOlfaFiSo1SaJaZBEcqmedArv2h9+GFkX6
`protect END_PROTECTED
