`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Nk08Fru/MsGP4lcpLlkCWGMxPXyJSYBCZ2e7rIDmAW9Ef6mIUBa5YgWKgwuH7jot
wZxRBl09yUH5+omM7oAdsm7m/ZWEau0Mzba//3osHQPyDAtGM5oUfOCKAztJ2r6C
Ves/FMd+z+FIIouL1/Sdg6BlM5dozV54EsjYEwlk/h5a4Uatzeb4BPiaW5XeGUOk
oODDgjwbkqHARZG55QHJYxb11G5jf8AyB86J3cvTQ6ybbItuyJMZ1EHK3Tj5DDU+
zrprbnOyc6840NSDiRHMC1K/cmp+4l45d8xSjJI/jWpF1lq9+VXg0MZSCGxzpjN2
QGpBiidPEF8OP+gQQZHyneGS7R5I8FkPtTni2mjxHdSBFV3uprnWZQVTkdxbiKQ2
idflKyT0jyM7BWTuXnEvqmtB1lo4j1rheFFpIGly342pwRCDjjSPXnWovctRXZ03
`protect END_PROTECTED
