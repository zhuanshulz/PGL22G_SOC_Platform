`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D+iYp661vSPUldbuFIf0Xj+K0VPZG17WW3lt1PmlZF6lepDmzUzpw+iwpcOEOgKH
f/SRx+L+9taRAqfHXZyIJxG7BYmIK4N9XXOIjgWIQQeP5tQtehlWYdStLl1EYuEu
pktUj/oP133jKlz6DImHIzJKB3gVC0FxH57lu8Bc361Ebe3hl3sLeFgHv+Aj80W2
5ug5/z63QxJ5M2ld3SDXgfU8vh4fuVXA32mV0tZT/7GqjTvB/hUQyt+MvoWVS1ua
1rQrrNy2qamNJJ3+Swafyo6YoU/z89bY/Wu9kqsrBXEr4vbgXzECviHyEAW4f0/c
v3f4JsRKRwHCSq5QSpfSnYjO7KFgHgS5npz3GrMw1895v1xSm87FXS7ao9+vEcLM
zehagHXyHEgNhjhe3ot9W0LdTUqApAlBNl2NtYLnK7JHyvw2ytcHbfx14+pPXKkM
4zut0kwOBNXAFasES7O2+DNd6YMN9UlzgF5jpn8pIMuqFWyIRCaYfnbGnUnXqjlq
+kS3wWD6wZMEFCtP7q8IeEPK+WdWzizNjHM11G7t8RE2ckpInF4MkR4o7vvrt5KA
qnjKxtizTlvbKxyhEJ8wvQ==
`protect END_PROTECTED
