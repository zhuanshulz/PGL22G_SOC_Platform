`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nRvK5XGgCVQRVyqFCoOVLaD174sVLf/QM/as2531KsHrrPfFSKr2GAMaFE1tdeDU
ZzjBtztPcN8nBFe6PpBkHgtShDKEbrRLWVkc2V38b4bmII4LI33SttfymzWCijaV
d5oFA0rzzzU5Yu5icqubuxvY32t3jVxwDmIZ/TipQ0WmTpK3ieAPQHAMIIwi7Pem
IWAt7slH3GzVRP9Khy6dCZAsN/RqGzXQC/JhA4GWXkXa8Pe4KjcFZOz3oigE27hz
xmI75KZ78EHz40lQFw+4ER2qWESIBJ5YY2PDPAsdwWABcBgPTgdgP/K9RMy3FDG2
LOVs6Fynch+7wfSaLzqmIuB/mQlxAHVtOOOWRLxtx08DkngTUZNr+AugaCWw0mqq
q1XJW4r4HUO3u5qxAopI5FUnM3s5ZY65BNSehyehVbE3NcyuZbnkYFCdzl6G1V06
paJzqgOSIlKsRINy5GzI/6jgo2VkzFqc3fiK5fBqXYR3PQij28GeiHJO2g8u0PqY
Lrg0AZYW5um/E/GYPupqMb2jty7Qgn41yWLT6MnNSQiiI3i77Yp/bqxowFywrSm1
uG0YFOM3BwXZQtx6pkuls54SbyIs7ox6Dq5TT6B8mb1GmALuMNLkkr2SgRIfjmAb
n0AZ/WSHW+EoBOSOVTegag+c6i/m6PrPs5mCqLI7ub1pomWnEG4Dl4TiQ4yvoMTZ
E0tgnSnJAE/5CurE9hI3N0sHOlkNCx0lzw5FTczroJTnu3MY1G0PCP62wG8nT8/c
xM+4P/LSNddZP+USN/2U006qs1Xo6FPCBWfa/9ZqBVt6WRvdaHN0sHiUOLX5PDKD
8akQwrnMpNW7l5tG2MgO/dYjvl+3p3T9+yX9XdZ70pZgT9qEyInlc+hrCt47izde
sD7ljb8ApT4d3OMTqnJdWlGLAa9dyY0wnKgXlmEsNczPv+Y51jZPCkjilcL4Z4Fs
XFtCK+rY0gF4xO467WzkbrYqwAtuoky4e862SE0uz1G8fApj62p7la1mwjaSBMyD
kC+l47EHre/cGlJZHrQinjkNOPEjgL9GzBNKu3kcScJrVYU068IxBxaLpOhhAMT+
f/KeeSEoWvV4R6XR5QWv0w==
`protect END_PROTECTED
