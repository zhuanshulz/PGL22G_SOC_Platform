`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RfmJzcmaHAGOKF7vilqVH1Yr4+lf9cuWvx3y4QxumeWOqhyglnCarXSJw9GANyJI
L39v7ZPn/YTTLMB16boQHu4LAChWVHJoPJMu2ro8ug8AWyrjqfDn4h5vJ1yGE6I5
dQjnR/UXxO9Q1FANz1nKqnedVTy7tMsrR+iE+BUJsM85dE0Tvg78UGW0VeX62PWb
UuCV2EfRmfhwLdR4pTNPe+a02NNZ5CRD2LZdC+q0eNXIUPSjNkn5FG2VffqxOsAP
1xz2pyZwDyOXrQDIL3463KWs1mJ+49+4lZfYYqbtjg3orB0ute278xyVvuZ+rPVK
CBt7vHW68Ni/NyiRBghWy2O2ok4JN+yJK/sQvt+Gx8XOE6p+6kAfPcRpdV20HidA
cr/L0UaAnEI7jVE8PsFtgbdqFN5nJSt50ZDRlwYDjhdoTeONVuhWWJGws1mz0+zD
LdRgmUSlglS8Ty/+7tVpssJ+cW0lN6MJtjgXHO5leyhlLJ2x8gn1Svk8lQ82CPJ1
qJ2Yv4YUnMGUpa+M7HeZci1n87YDmW2cE3iHbF9NKHe8Kkt5jECOxE71vv9ymQRz
GWEJvhDBTFkaxgc7mJ2DpPhYshnZxbnxqkxzqRq7i4dYo3WBRsBwcurr+HmWOUWd
rIFlZvYaGzfWJBotN3nH6K0pI4EgQ6S/os5ebMYbg8T1kiGC9buVrIFTfHO3DDnQ
rjZQQNgxni42WiQOv4q6jlOYLWaMAIUMGwtswLK8I4LrydyruArwzXS50X+ZLeyE
N2xEJANaot5T0bmA81VuBk3G+5tM6eiL+Q/5jwhEBnWAVMr3ZpFl7ljXAuW6pPgA
Pnzews4/fkeDgh3IBbCSMzCJlNtw7Yyw+OC0ADTJvtnEQY7KBckmVzUTcg0Qoevy
rB7fnsAhT4VRAZrcnkCq9z5csM+dqUEo6OWypaapJvV0CUOgDZTyDcnXIilkWXAA
XNTdp4QDRMAg0VTeT38cGv6NUeRzhQglq/5kswKvWalSq1nOSs9lgQvszpwj/Oyu
MkzNchCTItBBcg+9t6crwbMmqGRU0n1BZv8Cvr6sYCexLGRnlh7Tp9fHBLrwbRHy
poU3fMG6OWndQxqBl/JKP9HJkStGxSiLrmPPGHlnyDDYR5IFIweO054tvn2D/uL/
DVo7tnbxrQyY53LuWjFwizDvCRFQ/CLSNZoN8uCSosFol7r59sfA1K2CwGtEBm7x
ymQIMLZhqSDg+zpYygTO5jJ7UTG7zFj4sVfeoQ0NnbKuHsvgpc3ADYaXa5oOuGk7
LrRsg/zY9WpQpfiUxHAaAvU+N8TeJwcM3g9/rr7wosoUVz3/gSP+fnsWOVVwrLyA
fSQvL8+SubUkESxv678i98890Bi+wUK4N/EhBw8Ist8oDoRYTNtMzph9BALJX4GF
WKMX8I1Mp1a8dE4sAI+xunDKGeB57BzPKIShmYeHrAlwOSDBA77mcnYfXn9bE1KW
r8LBaEi13XC/TZRga+PYYVk9JS5KsS889vguoW2wFZBqEszxuJ4TF0EtfbLYmacg
UCxYEOsKVTL8Rfo+AOKf4XiojvUp9XcgCx3AjH/JBxwjqg4RPkBu9trLGgE00OEW
ZAQA0TAVfwDsRZqZIj6vk2Mjq1Ny+h6larh/ZB5Yc5tTQNoURewE+2Ah/HfeF0Li
T/6mBRLojnjLnmdeU2RcwRGGrvmHynvNrJcH+DLvol0rj6gy8RIvjmy1zFcy+GV/
M3U+tWhVrp1nCptZdOXx6+igGwtxKc7k+RK68Fapru774/sJ08pq2L7K3XlSUNri
d7hroQRF0Mz95C2fb6al04qkwANyAZF898RUNsbm/xZC+C/wg9fySd8tfKhMLQD+
0M3SjA2MMfvYpbTxkKoHj9I9kJ29xIdJdxFsjsIMMmGKTvV2PiFbWSBXYgPrgFE2
+QH66wcjUq5cr+9nVuWjXiVAuL1VfgYpTkRHWUKBz5OulZOxHb0qJUhYql26eyq+
a9vOtSiWgchYmBLIESp+wtoGLQCzGXLFfLXmO2FiWjVRx7VuaFmanH6anfxsy2WL
bmIofSIZtffAjgxmGDhP8Y3rYryy/R5O4cuyL4DcRgDdIiX6olGoH7uax3Z92d7n
3WS6JzIVd1irWj5+qhgxpL8OZCkFJmlFVubDnCIMudrhVXo280AOtKoHbEfa6BDB
TE0nrP8KLGC6sGEJFRstNz8YWhnQZJbNjqVJckX/5y18D8bg3gqLLTnpH8SkF3Lh
Zhve6HwyATRtc8A08HHh1WM1nDKSQdMHJe7oYOa80M6+eJeWYikv6mV05tCkxhVq
4XpBoTCxNGFnUAMgxVhSldEfLw/TEDmgOOxxSHtcpMWdC0XVKq5517hbiWDFhNhZ
HC6b9tp3InGlEO76SPbqbauUVfPIVVqvdACDE2YXVAuyHAmnhlPAH7oEnH2eXp3w
`protect END_PROTECTED
