`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BC0fj++ut8Rm7+xHVFtew+ZaclAl72o6TksNVXeCcmcX4MaYrqqjn9IOAUyCACN/
1/0a/pn3RrzHQeWcX+1VkefLvX6ru5mKmXjcqmDX8goYTlL8DP8RRlwBZFuGxFIC
sCjI5cFUOcTg55CMZdEP8XXTXnzOkj83LW565ktE/eCGXKTH0ryatv9e/XE/1ZoG
zAL1U6LLI2ETMRdo/Gq+/WopQwZBhm5vWg6+MoOwGqks2TvPaatOzaqERCjRHG9X
f1+SK1S+sav6xuEel0HzZhbW7hxK97NCzlm/MlohW0PHJPjGhC9HgT1h0SmJkBSn
oX/wvcobmkC3TonbL+J/b4EEqz4G1kmbzwr90aip3gQYvlx1seHvay6cx4LA3O6t
iOsnskoyLyq0fAbOVMDHD40uosEKWUDztu9I4jDdJ1YupciiRmRfHccnJHDcQUDb
c5F785egp1TQ2Fcubq73pWVJxMBlQVvUSptHCWp73ibi2BlJzpsIHksATXx7nu9a
ddGdzmvMTtKSLbYkjKw/dvLhmHyq1AACzVpanpTt7NZVoGA/mKOzUXr5s4lxIji/
HFb4nh2AgC1cLFAfx2bD7wRlKGV+1+nzOt4jJJocA9HgW7s58zlKErPepqLbwFpd
W3tltlBb661UNmiyMxIDqh5pBA7OkgviRbg8lPQNAnm0H8oop1QLDcWV25WgiYbi
V4jhyNxAUYGXvznIhkPi1RT1MtlIFf9zpFWY4mIKDepuC6Ob+mmBtB6MUulDe6VM
C5gImtyfO2V24oK5+WDeVN1bLnQN0/miCNOOrclVmi3mbEpQMiitZ++M96loVfza
KA+yHqc6t/1i1p0lXKTmwQgZOaWRwbfjw6GtK03DOMSW+PwRrqxOZ6kFrli2mcvU
`protect END_PROTECTED
