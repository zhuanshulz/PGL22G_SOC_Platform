`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7NNaw1OpCKZgt0/SrCybV8iletnb2p5EtAVkDCWxtS+8fBr3Rqe4j9/AR1JKHPyO
d0reN1r0T/EyIO6JGebZJJfeyyka2whiDqJFvEN4VPgUmLm4QAPJ2gIDtk04GOG6
uWyYfqb/SHpHeXMdIWpAHLGnUPOyHODh5S49txGfJqlaU6BpsHNB+b8bft0pmOWk
u+MqA5KyEXQM6aMNn+iAi/5E8SIrUHNLgGdvo9AVzmZMooKWkD4HCYTLt4eswiq5
V0IyNjOWRekJ+U9LjkB4giCsi/IzkRydilfKgLiSwUq+ocey255wrdxPklZTxTY2
H4TFOTWmFaZ5AhXLEl1ETf8HMWdvP5CMIxXfiRnjrd9LCIbbsXKatfAyUve+G0LO
JD0QgxTZUpUn4MdzWheza4g1DEUWudtKLMgx9Ejj9Zq4VbZuIjuC5EarUFi/C2mN
PjRF5fZ3HLzPQGgRgqCxu6u1VZ+o8N+ZWuTVic9IAEvbEDxrunljYDqJ+qkpH4ZL
GHEhepUBPmqwGJPHpj335fa66F4zzZhgO5mlRE3idnxfkRGU7k6uVGCcqVL/72P4
FjKD0Bxy/N6pF6WW0nt1LTaleCoxxWAmGvtM3x/EpD9zAE6POXauHid1H+CdTH1p
rfBtKTned9vMjEpJvhLYM2tlIR5vrCwp9evoNrVMrFPz652/DI+ctjn7VVS3Hhdj
ewYfIPquFf8jZKZfyF601KhquVABKhnJtF6lr/bfJnfjGVQ8nvVQIKT/eCe3OGOr
/BjiL5LVNFipbjwO3Sj37RbpQrLuIjaMUQKs4RTd0kQLBF1TtR1SMNEEHvxGPDMq
e84LZMoayOLbb/lKXLu/t3uGcUdpHSiCK3a+bJQZA9kL/0i9p5VI+Lzq8P2yHYv6
rNOUmXimojkmM6bU6IrTqc//YxT60TiPwOGkE9S0oVfGQ1qBxMUrXVcZcZfXpnZG
+8w9TrfHruZMiZRXKly+Ta4jkYtyD+9Gd0CK1N+1w7O5uiVYtXrtAN01ws0ET5Z2
t1+6H3FKkEToi6+k6GlediYmzSeytKNtpUyaEQiZfGl6CqFqo0FoqeBrbKLqPFjn
8p1/Dq8dttigE6npZRQV2ZI60wYmm4k7OWYLzq83qcce3VWgbTcJpD6WX6OyhgX+
c0QZjWCo89De9w3W+nhv50WynPCf6uDh6hS2XSxElzgEExXBTwqUw1F5wOfOoiP6
BNS+39S9boe28peVnMkRnbPgw0WcKVbpW3eQpM+MwKyWWVwk+YWFirxiEUENVyi5
`protect END_PROTECTED
