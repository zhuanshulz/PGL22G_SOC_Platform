`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jvXRA4L3EVOUjrNbyEzLHXfcBcxgKFH4gPWePk7KdKBosYuI5wJCha7mKvDifkte
rrYTtQV51pJZ+wtw6nbYajMWqC7Rx+QZVbBwduxwON3u0xc/wcgGOxhiAcQ5ieCJ
kvfhWhMeXrILbeNER06pzjPy0Dy7PEap5ZrpQvivxAt/PFCGnl7OgBspV5+JcYD/
5oE9jwVESQnCAinrggJ8JOF1tMCcQ5XFlPG1ORIC1O3ikOzV0Ic1dPP1Epq26Yzd
PRcPZj9ysMEYqqKai46t49+XJ5rdi2S/oVQm5R+D9vRI3hiNIZ86LtmhIZLjvYQU
+v0W4C1KZvxcpJikN3e2y9RoMck6tGFmC9GpuQrfXvmGdKvHhU++WY8OMaVBUr5h
FHqsy/zrhcSNxq1XxYAWp0bSRKdsQ/7Rp6JV2ZfeHAJctMI87NPV50ysyfwkUs63
MKupUqoZfO/U8jQHpBoXVhZwjtkeWihzTMtjQbItk7GD95/SiwF3FV022EACDDzZ
VSE6S2C1p5P3XHLjPmosKzKxIxlOlEUjBIci5cM7m0uX+vOjJ0J4A2RjyogbJYqo
dH1K85wEbDK4RiriAUz7s5aApmqUAU9vEER6SYyWPHIkIzp25hPNkBdbf1XYxUxC
bw4ds00W/zTwF3IaUpbz6NuzaaSP3TZIz/ysUwM0s+WoGrpol2oy82nkzEe6+JL7
JzEim62aLIY7MCN2rBHvEDEcQV7uMLe5T5TWeSCfrt2G1VDKNfYAX6UbvqViQaN5
sn5F7ThKmAeKTGhM08JTEgGUnNE1TlSkGgs/4oC+XvvpGRvArhNQZZ8qvO9E7LGB
LdaG8AHU9c82V/Q93YRxAKVELYeSHIL9IGSzLnDGNOZME67Uq2/Qx4Gnxd0vvdpF
PkiMpXHsiF38Nm/6U6EdKYA0gIywyWrS5+LiB0gI8VcVNfkltJHgGavpU0tVCtvO
H9tm/0e6u3mQ2yBc8mJ3B2kQmTql7E4JUnp3JM05g3+QIx2hNg6B7V4GqUx0G49X
zyhEutkUZirXVhL5yy337NpzfNPMKNqVb7rOZIahoK40QmqsXORwIjEwXEkiJsS3
3R3mNm6lm8VbVpPnpL2+BVfe2WV8OYA8LB22YvQWk+xLQSlWXd6ggNNhYI5UFWUJ
OQ+ZoDiKRTgcFoe8ZPVfG9j4B/oKIiKOr9EdcR8uQsE/Fyu/Tt/Iav+zPRKgj5Wh
ooWbHv3uAE51dqGudE8o9pBdUj1BYNeuOENf56A6Lot/fdNI/ZtMKqgKSCBT4ONt
uy6r5RorGjWWJvcJ40w3CMvbCnsGmWd8oIxyRlx5HQQFnHuAzc5UcO+aWjMqlI2m
vaRUUeoMFMI+1azeIG+5oZzyDyj93CWgsZquhE3a5XrBfbNPLomLi5b044dBsACu
XvIIPAALRrJNqZrLzqtxuaZEyph0UVNIlmkMPTxQXkAeYfF/UmumTUrIA3oipZex
f8dzVg5t3d+IhTGMsvCBIPsM7KDe17d027KFwMGlSkw=
`protect END_PROTECTED
