`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PVN4W8EMJB4AQsOuu98lY26Frr+8YseMmfDEkD4dDjZx1A9U+mQY59Q9YozIXyT+
LKjAEhxW7q/jtNrGZEYgOTAKTu9js72gjebFonHpkEBK2b/1YlWcwGqeKlzTRlIi
iWvWmQoEyb8PZcPfNK2hYvRYFvfaSV18tkmjm/mmIuNyXvV8QMnGOojWWCP0+GU1
5tzAU+Z6dWxu3OxLCGU9JAdXU8vsbtJ8Ix+NdPLhm7MUZXY0aIAG3ZtHD5RtDKc0
VktKrsMhckMghbIMroXLvn1xn/FzXuBhgv8VDIJqL8eDTd9Dt8Mx8WOBTD0jRxxP
peN6rx76TNLt5XGlYZdJt7Qyvoo8uktTOPnlNGmwK6UveggKIhbuQU5Cr4HuDirn
Xl4kpQXZqSyOMMb3zwLd1ehVZDO5a46Xb0tTVx5tn5usX6Twf7qh8z/1gMleblUp
`protect END_PROTECTED
