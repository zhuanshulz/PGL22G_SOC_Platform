`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aKR7cp3ROs5mdYGQVt9afaBp9aX2YObGnfBwpCQRAEHHa6Mrkjm8IW9RMiMwFqKj
7OVqNs4IRTsrXPo9886ePPF+jUfb5d4OYGnYunHbqQMuYDeFlxsrCbCzyTq0fuOw
oE+cdVoM/7EaVz6Cw+J73hKHchRmRlBUEnjk77qSpx/8bcDWxyoAXNjbSXRu7g6/
nVuDRQN3zY+z0+sRYIhYTgI8BG0QBwGdmQ5hFKSZmHU/5ICTzZD2BV1K/cfK/MJw
NCJZRynVTMi6dFZvr5ZhDoomQiq/uunLUeXEGNYpOzX9pyBmKFa+L1QMl1DcXLb9
iI8U2x0DD1lyeNpENyiHLnwx+FngYfAJMjTMQdRTxuRankhvDGUs+EZKG6G/5Yqx
JOGvgsc3SuEORYMA6gZrPWUnD80gLAnfj3kJ/KKpk2aZus/EZIa4RywcvGjUeP5o
TIt42DcQIqT1LdgImWOTZts+kcn0lBpq7AespsliDPuI75xH7ZnLDUV6Mv0N89G0
iXR9LkDV6S/GGB83uilAC2Cr61CJYR/45gkh/rIRMCyVDRWXcu+3bwsfpkxtG6yC
7h6kMR1777M3+wWjrEVNwaKaVdXidkdU3RF4tTKUfeVqYN5bKzIt96aSMVLMs1oH
tNHgvbTCx4QfxPIo0b8mL5BHFB+8zzEIFHCM+oE1KdrIiE3gqKIQg7pwF346Ilce
gGfa2umJ2ImQwpInEqZv0QhckKwvTfzVtvV2EfxcA58=
`protect END_PROTECTED
