`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C+FNjz3DkmQC7wIoA2QAVOU9RV3cVan0rAIsx9iYshkY9SbbQ8MXp3LCwI/E0u7C
mXk8bI1/m3n5dPLCXpGGKYtfB1j/yWSlL/B/ehQLddX3Vow8LF8UYO7bkj9sXpqW
U/rvsfgVfXtp1aPaWw7LEgd3+edHWz/S7q1d1w/tCx5Dvh9LjXxka0zfQ6Kb2J5Q
MqkL5u0gmfhNqZzE43bKQCa9xvsqUfM5HTwsVfzsXvICoU0n7j73GNWZ/3LIP2I1
hyPtVAc3QAaRJWJSpUG3/55FP9j+tyzRKjNvmE+OuLiGw8nP52XX97Ld52D6vqkg
`protect END_PROTECTED
