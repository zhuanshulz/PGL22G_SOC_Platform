`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bDILYLcGCJUZwqI00R6bax4tPhkvHLertIY1zIVwlvSWPiWoegHy9MVol74EUfHu
zT3NGXmFb9xM7s0TfcQU5lNsZby1Gpy7xoDUNgGD/zbL1GNARGrDse/GwhosN3nJ
HEv5fKpD61v62PpH7Uyaz+T6jlTlUvU8gzkHpgK9toU5moOaLk21HqVZX54XXeUw
Xdr3sY29SK79zf5kHs1cX15wbJYnAyR3bdX1PvKyroiDvRNxcTTUaqLbzs33cguu
Z4r2qrCIaFf0FuK/FI4+N55h5L1A+Cq9FF3mmCRnx9uAmZWWqTX8mIHFDji+5wW5
RO3Tpm4CgJ2jCl3C07oaswc7PqSPj7/BB2NNgjdgCQawqHldGhqgf/EdXy/Py5R3
uTI6QkMv+8x7OBTyPT6xnnURfOEr9hDffuH1DgrF+v3HFObKaCNRdxiWAw34hL7a
hUTljKAuYbZB31jesUgoGR7XpA88fdSbIdoGwnudwVg7/qldQ+/yheZY0u+Z2X0F
GmjMDIgYeA6rZODuTgoE0RtQlL5pnikBVTXOHM5L7vChV1C6frMhnMDyQs3soCKJ
gwlmuTlXB5Hem89h1MHYMD1UuwM0yygwJKevi2Y2kcd+BLL2bTzDksIM6/3i0a8M
s8hrheP6SSmFMA59V60Z3V+NkdHjCt8p09KM+VT6KVkvIG4Kb3zRkwWEAQGixOia
7U21jFW3fljNWFW/EPOtwT/Vlt+JZEgAG7c6l5xJt49ICnQRhB3pva91jbuvuFnw
G6duT/qW8k/YVeof2yuExjT/DZLnE1CeJ3CW81gjMSxo9irvYG716HLUumG52NYS
onS1pRMSF+JAdUAhsKUAg5dv3eEMxN+eetTbYtCRQW19xULXTE5zxAYpSnC1Ftcq
re0onYb95vsw0ytjDlzJ7+MVSU3Cj0/pnTE6/0JEcL3bff0lCKngIbvV/yPLJwni
+gV4rOwNqYV4w7DNYqQQtmr38CniUZaoITsrtrOAujvxJQygxtFH2z8rJ05hq+6F
Od1hevoZ4JIAkCZ2htCxJtZGSPeRF6zKD5sGbrEgqjDl627x+oKu8igMLBnJQZYM
U1quV0Rx0k6WR1gAdlqgSxt+WWEOBGqhhFYFv1oMlvJC8Tl4OfL0CUcK21nvpmCL
2jOeVs4wGVAxpE2/u6AwUz3CyHWYhEAg1UTw9cbXAxxwKDbYZ6VS2JE7z56sVdYc
FI+3Ne4wkDHbNIpGGqDj1xpdXCAK657OkLMpJTFce6iVzcQ+IETqAaYsgMe3kUN7
sw/TQ9CM+KYGll4vWR3FXIQngu7yLScIGgmK/tZZ+SxIbYnbXhzAxJUffa6L9JfL
8WPaWryg6BP0GZCM4bipmMZG2eDA5hDy/Un/Ajyt+GRcY9ELI7MZfaUHrp6/G4LD
BQ/vIAXWaghEpqmp62bAzv55+1lQZeS8hzI+r67i2091x5W8u62rUJdbZpN7QXlK
UEvqWZ1N1QB8AO9es+iLsGEIv8qZIb33Ed8Fjg3nOBrnqM+kWZyLll8AHNGx4gMG
TZevpLNed2oIeSp7osoLxgCEhgWV2TJ6v2D9wmHT5INmXfQIqFkTd6A6SbTBSv0t
0DYKE8BUAmVOsM4p23YUAPw3yiHUAWjj+EIVvlDJYb28MNj3uvRdDeBaiL9+o/3F
r8ydZ5SctXl0dYDnSArAE30jNcjS3RIhJ5xDGc9hGsnFC1+IQTlNC8dR/wjuwlJK
WGclOEGJL7g0eh3+QFHTcKcIf1PpCk5/VVtR79jyfXlMS/QB7cUzkRYdtrG9sOuF
06d7EoaE8FFBdo0PxW3rWrqJGO1wH3RIl0XPdTD5i+qmcY0fwZdUzRL7hI37BsyJ
ByIblsoWh3YhqYchXURb38FS2Pz8HGJaBa2UxaVNa5hV1+tDBVsCBedbUVmdWHhF
5ffiNphc5Zj8GSLdyFfuqdFQvjMClOFwGMmSFwUX3QeE/Q9eFoOF4TrMEk2cUjBx
ZpSHteykbNfNmOji2QM608oyJIYxekT41OQYB7PBQhiCVF5RqaCgqnN0T+dUsB2l
JmqVFarxAuzrUPvH/VGlo9k8k/I7evFAmyWKHUunWvH0XH/Lxf/vMGI4rRBzO1eR
znga8ClcVDuq5Vvh89RoUhY1e+FSTIb7+yEJ1AVhhu6YaXm5GqorBBAyBUJW89vW
6dWUVKuOIohjdqvM6gpzhfHr5069BAe47XmJoei4W7luzCFTlaIIgocjOVsiMuZd
6uVJGAkFsi9Y2PaQr5tFig==
`protect END_PROTECTED
