`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MG7K5FSF+w+151hmzDX/zvSnup9n61cgtTf5FINLGHCnpqP/eb0rsDRsx47ufOTm
B4G/KJ1bqGmXLPTFIaBV8OeQAJGTY9hIAwqUHQ5zZJW0E2DQY+Fqb6NXCjWm0YKl
Gu2iQ7PNgRAT4kAoq+nsKKFx4onAe81d/R65tRUarhA3TzTrfAMp0+9aMyIlxpNP
5CjGml/ahlz7hj12jSP07oMu5bekhuJKGUbKVu2xZnEOU1c9MyKJwCqukioVcjdm
TPsqR+ivyT5psAa7CDweW2XlV6cCn+j8bKZ5yyWkKaruksdJo1CrXBhckzBNJDEK
bKhaSbWHV80/5eqnchz4pdoY0wiJfdWYoGyMDyzGDe4zx8VDAhmTSu7uIET8YreV
H37dpBvwVpOc/ydrbq4cjqxuR3GrIFb4XiA05m6YReGXwJVPJX/ATzrl/FLE3G9c
Rc4RXgBroFpC/jxAxhFE+/w5NPWUDsnH9qJk0gWHlVFn+Aaxkm+rt9/K81SzC5cA
S71FBt5LmQTmPfzfj7DSnw==
`protect END_PROTECTED
