`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uTDHO9ad+Omok6o+6z3sZEldryl7WZm9ZjAIAQDhVSVMHDznrhHWmH0hukJL1l/a
i3D0nWLNQ695JKN4gMkhVJLtqXCOvpJy9Pd2lUWzJCTWFxq+lSKO+PCbYqT8W+7C
gfNi3e50UjRSwFsKCzZPw31cUH4mtrz9KnmcK9KyQCxk2axjdIt3FRA4+XFXYaVQ
Zy9BZ8wovOCkPUqJcTvFAR5iC35+5xuUZ6Hxc/KeZLFlrqwe9ODlJZvJV2nQZdVO
zYNzWtQBveRijxtQPHQCKV7pCjG/Esg1qe4gOjE/6dHMMVCgoIW1fOi2xOQhnXDH
A0B70RTSYLaFMJ9HSUX4Qo/jX1sbZccelCIFP5AWthI71RteXD7Ry2y//9I1wbU2
qzSKJCcOWso3bR0G4YcWdyz4Xd5nISLXNbbdS8+oI9gkMmLtxRrGiP5k4v1u+tFV
YDa6Bv8oCeM5/Kqp3Nz0LIMMpE+uS2YZiHruWBKINLC0aduhA/TisLkREpgfbFFz
5BdnGqdiAfmA4v2ttzTGib+FGUyGK5nvpkIxRHaHvhncz0lf1da/V7IhjJKY7IB7
c87TKnuxCrekdWBJDge2c3AaVDHXpa4PAPoeiIoT+jUU1l9eNGarq2fMkcX2z8mG
Dn4FbOHT5x9ljJey0nhuMpufrlNkmLD9ykbgFsGR5XPUUeK6xaa4i/Q2YZ8ZwF4E
bt22kRPjlXNyDoGDM0TtbD5CsF6W2yGSJM/Ju3LqQjp8+khM4rSUC3KYn10S/DK5
l6ygJJbpGEET4Y+cH1sCq7GhB50tErgM+mymb7LMtEENDYtPYdc4lkrEdVri6XP+
L03z40iwFTqFcx6Njr6GQhoM+GZc0AiEBgDWWiF9nUxFqofalOYY/rLuDUdD4RqK
98X/QLQU1ZR97bzvr7M5Y+FtLoT9PRhqDRK+WjfocnCwrDx8iRVPMuxoiqrRgefm
B71h5L7ZgmlAyRDtBKHi3ieokea6B6XAs/hYiVSrOUo=
`protect END_PROTECTED
