`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
udQtOod4hEkhtoMzESrbvMFUNAinc962gclkueoRQenr5KKOpQosHXZ+tlWGNDsh
Y4zqCVWrD1oZxhCJ1Fy+FKQabRjam8pHPFKUM5ccDBchh0nqw6MJDj9AcTPXed4n
FFxBpzm/V0T6WUiV8+aye4O+jI8lMLlygFNDU5h2VWtvqX6J2iEr6KiX7D9u702D
1Zut5QrWisc9Hv175X7WAxjohZpqQnyGnvH1D7wAmi0fUccXOufGtsY0Gck37A7U
NLAbnt5174Kt422hBlAy87+S5EuBvrcH5drGTxzgSvPkWF5C+kmPmJLsMBn1VaCu
q5Ylv97GZfb+HxxYZAupkqJbudYgeptuKhRXxBiVuGfLniBJN2LjK+GRowMihpzn
VviM8Fid0rVK4w5T9y36t2zBS8p9BWrCaBbzPGmO530PgAQf0rJ2K1XwpN7VeQbZ
1xC4ZVEgGoKIEAt1KOoCKY0Sg0FjFsf//VY5Aw05a2IY1WK0WUEHdvtW1Glmuwtz
zaZSwgsCVpkYmxmE5as7vMEn3Xlg24nRbFHhozKZkL9D11u/Wb/IKHVgCX/Y4+E0
QmKT//ws7lyuCk7gF84uSCuSMhtyZfEWbODBDY2YgJxBFRtiDz9j75lJR931ylHj
qYdmaXZdGkcS+ch4qHEYWoZ8Mn30RKlfdH8Y25SiOL8Y4QngeJGFkqO71DATSQWg
Vq3x+aHiYtv/NAG5Vt4AmtVPx8ogCqAh/qPb6smY6g1Qct7uShgobakYUG3MPLkU
OPgHxuc+yy/xgFzKl7gVoMxBG9KjDguEDp50DmDPrkPmI/iU5Lcl1XNM9BpOq7S2
QiWrKgpa1aXPKZPxJhJ8nRiwJXZgZWDzk7bzQ9fTOYZkDZjKMKfhelw0/6RZ2DhP
btzR3OCMZeV2MV6HWqv0Y5WSWSN00ly+WiLCWz5QJ97KWfsQ79kQVp0dmM6bA91t
TIiiNgjt83BUIDsZcRZPJsmqndLUYFJsgWogQlFrCPjH18RXvcwwB9toM0lqdKrX
Z6eXcccBia9Q4W7LXjfD9FF/RKeQDV0q9gkWPlCi6UyNFHgahOgcaW+voCNii2gx
GqP5SZzgle4Y+bZwE/fqaVnHvKewil6357DdmGsMOOuFkx/VnWaFcl3/8zOvp86G
Vn0p6avyoxUS0TT5CREPGVRly+2wpCZr5ColywR9GTcKlu3A9cUuJj6TMwJc0+TT
krfe1/rwKSvJd56goLTGXmyY/ssAZirFslQx4Zrki+DIxwKZ8t9CT5BhBIFZzfHF
P5Qax0d6AA/ixDU4qC5J6ByvJvhO/xEfl/FOKtTGOc4PB8KBFwfhCdJcPjKXQPdM
WUnpx/qO5wXhE1SGQANLdX51XS5umQzeR+c1wFzGsZWVJzkaPdIjUqBN9qOh0Dt+
1ya55YUXfF1hUP4L0sAmHHZmgSNKYZinvRZBX2HJdTwBrQ3KUvkaW282oUFwyp/N
5p0ewhzC/JKBG0WOScMg9MZDcaOYGTRNK56sYM/7wu7/wGBZRDedLuONW3nXoMD0
VYXYMkLtV9hpeTCmRxp89p1T8aFkok6wJnk1iw0EoC03pTKDeORhKLlVhj1OFAV+
TQIDtfMtC095ed3NJJreWWWkgV/8e0Fbt8qm7XOUjdSJsHQo4JxwbeDYhvtX+nRy
EYt2WvnlF5rjX9HCpecDZONYViApeshB2G5c0BSiFK17HpAzKHOdVn0BQBu+vXU4
aPtol3by4q2O/oIZxG6GE4xSh6eDiNnZKkSYzEWUpgPfcfGd66XYNmmShk4464TJ
xnNi7tYsVRh9/Pr4pxiB1HQuxYEuCvoU2Cm5ic9hTHkf05e+qg7Q+UcgKMJ+Zh6W
g6YCOJWt/vVYhtvoM8q1spNsymOjXKSIXZnMngMnA6R2ebr/U32MtR5PkZz8CiX3
m6v1kc43hDVTtZjBrsoUy7TSgZ+efDS1yrYH3A1qwQrgiPoQmS4jHlxY7JzxQ7OX
alqFdkR5fwA1WBVbUeIQxmxFXj0Dm5bUNY3D1I4Dtry4HbDyi+y1rk1VnBrrkb8g
q1+Po3ciT7CY9MsZ5wRZzRD/P3s4vC7v+4okAUlIETp3PqAf+IVYMWmwq+CLSjN4
Vtny4kO/0amj3mR/HCoODAcm/HMjwAad29wG47dp3VqWN81oxjZpX/Nl1+SbX8uv
7lWTZIZS63XO3hDa1G4H2v0jC7oVIY30hgN33pyI2VJCrSxFZcb9bISiUL/JaJNO
Me3xhR02G1+9hz+BZF+tfqDwpzgrZx+id7mRr0DZyNUoALqXL9LtUMtaC8p3vHoY
/n4oWAfXaBew5BJe98esbnIrCDWNZgNGmJGSohMQF+HBeg/LNlnT1IZe+44I4rX4
PrgFzbwPE1rzbQ7ekB9id43rkXubD724hd/mCkQJaQ+/ZCbodwdLnIdmCTgxAnaw
Zu7yHboUyCIgR0nPhWuUZZDegIpnq1YCdy+KHX6jcm7oa+P+sxrC3l8KmWNXOM3J
vQeBD9i1GP3uv1Y7WB3iH9MhmIOsx+rFu/38GU9XMhWgYxUhcnuVtlbiz3cPk/6M
sKGzYmmkFAob2974TIr9bh4UqHF9MF4sbPF/4fgOzsx5fwegML1K2Pr5t3dltGfV
fL/8S0E2ZEtWiROkarkXkZeqwryCMzhP1RvFeSfcKRAPpVsn7FHQdx/Y51G2tiPn
1cZsxyyEEgpKxpjinjFwqYp4MfV6u3nDdyzeHOkCoFIV2xner38yybH5ckNTKpre
h/JmJUto64UUoYOgsinrHWwlBvrvwYYyOZQ5vN7zCwF8il11we9rHMOPQaEaSYZO
XbYUX2LU16DGdo4herAC6yD3okCUbK5Q9Kif+5NQwr12CqAJ73238izXAdF2ru4a
ZkE1RK3NX1UcYgNI1YF4Hp8I5GhrMSu3AZIboaNgl+SbjwnY0MWGSKwy1uEjful1
9ONEk6QG5WQDgTYZ3jshU83xMFqBBnjcsquZ/aQO2W8vEw2RLQ9CuCQgK2ONrJdK
bnmGMgk+pEHg6ta/eTlg98Q0Od4OK6mQz+PSYKZNnwXA49pB4uAy+u9MJRzE5SSi
NCdrjgJ2lRu1ykL/PAbkv4WrDJWZ8WMTK8WkWLAmgR9Rhp7Dp/iEGWilY+3UU/Vy
i01Ft6ImdL3gJnjc11YCtXBSkiPBJr1H2gTmaJzRvXIUkh9z914Qll7xLPgIsytm
dCV3DbBJeD96KMKo4CY37y3FhBwYdkZuCvPtrULHnC5UgREGUwvn4paWoLpsnQbW
KOXVuJH8sCMeksD6CwhDVwOWm9z+0TWv+ecTigWWzFlH/Y6i+bpVmliwqDh8AUw0
U2Y/4f6Op/xcnN6mlAG2kfqi2wmbznh2M9hSX1zUpNTS65fzP+is4l8opF2zfSdC
zhIW2fVVQEK3rIbGVd4T8tW7L34VKpqfYi9inTwjGXKF+fv9fuEtzWBndgisjJTp
/D8wQ9qVXcQlYzll8MtOmG1mIYA3Od8OUgV+Wtmotgku0x/fJuvhQHAe3MuFNYCF
7L1V9ZupPDUFoiBQD6gtie5SIpuFZT2f9AbmVunHxTXOvSnHd6AddOF5ViFs+stm
yaNrWALlR1+o6hNGjLvGfwM+Gu6+pbYMRhz5iafVwfrqryoze3uqDvoIFvWS/WdB
1bCFgvQ0AcOX6ScPTB7pXkaety+dTDn3qw1HC5uJYAKF9sxIHUeg2n8Rrd5e4c8B
Yi8m4yKURmBL7iRFREKGg5gii7S/4mzzgRH/7TTOWTLRx6IOuf2QqaYWGb3CvnKs
n0nS1bseQ1Q5cvz5rcrVKFsd2duRIXpRE6XdKYRNZu5kP/3IeVg9denW/6sSzop5
AaqdUxt7chlKEAyG2kPZIsn9P0Iv+iJg1ioFp7evPLt/Po7VqlM5NyMhnod7vUi7
b9b0j1eMtJ0Mpl53E3NCuawJIMjNtsOHtrK1HWkIuYNF02ReZvnx8JsQVCVFbAnK
PTAkh3A/AABoj1sGpK3rrBRc88mXPVlI+Ss1EbzCnYbV7zgm1oh05idYFa6jegBX
WUianCtdkLYXdpPvuUhAhDKUbG/6OSQi/Z439689ohlH/7OCsfP7SBoJ9uLEYDK+
6sAxQ3k6Rrrqtu0mv8Qj8SaIaciqvj/+Z2LF9JyKYMc4ek6aVruXafvXaCjf7il0
uuFlDs/B1fi6tKAdoIxvxy6anKCrbLntW8Ffr2J+daCpw9IE28m4Sonu7dKPEB1v
RNay6SnBbsS1XbNsyT5V9BB0i3ewtvPtUyLBpIcZqPwQFyf0v0XM7Da3WQogAwWP
naaz57nNXtoEoz/JHYgJWxZTdt5TzS+roFayuaYno7ZiXLHOSrel6Zgtji0yvlCL
o6PFz1gOAqYNNTHKZ9s54X+N1fhg4X/RuehkY6ZYxiQGGfu5UWmAWLqGRhk67qkr
fpRi4mJiClYVZiWge19Rl1X7+f0H/Hhju6exr1Krb9ke+l/TOBVw2oUqJxVrArq+
SMhpV5cnuRl7U2b/lp71hGx1LQzO3aci8a6jpj9KwXCZbfOngSoKDxFkxNcjY5hM
hi669o0H7hgbO4mktBOaDZU6RnranJnWkohTIAp8BcFb4hnJ86aDG3qxU/7oHaSQ
Cz+Ohc3u75Etjei/XEDVilG3DNLK//892OszUiNy2wCeJaoUEwrSmmRloifCXRu1
stwfQBsAgtfREHHUVo1Hw9pmZgy4lkGtwAg8XHLA20RS2xE6uCGojUYypTbrgZoH
E2bBwbgNkvKjX3nh2/HXt+ZFzsL4S+RalWV388y1O92yIWQT1UkHn8GpEp7cyBD2
AvdZeLWe+esIDlfautTn4wxTTBIWVG0Gu3TuHuQ6mnpXAdMohzuhFqD+vLzXAjwB
c1vR2uZ2/Ze4kiAsAbU5QPPk/ivxRRJrE7NrcAmnwi0RIrK7Kb3Cms2tp54LDCEu
Ncup8qNXqtO24+mB02l5PlZIQZt58RwOxO6LV2I8MF6DCeH81F45yCy7ENO3pL2V
ZG8vhtx3wwU11ZWGU3g1qAzVyGekQ7o6YnBwr7fB9o7zPgNkfy/vt1UCFll96d7z
RicG16Hk2EGubZnaZ3JWkNlbZNgsMXAvrwGsArwzxpPgY63rACUhboSI/Pvypwwn
MseNrYFt0v6wlitHNcIw2CaUG0pbsh/ilUkC4Sn8IYM5sDht8TS7//Ir3Ufhu0Vt
37o5lPZt/uzq05/HvpIjw/tL+C2N9oVtYbegmpgrje14Q1sKEpegMk9jqFm8fcwt
HN9YxopOKXYhKR4BySOlxRzk6ryYv2J22mjsWYAt1SLrtzm7zGSMU7JO9RCWl5+g
Yiac43NRcY/sjYumGjtFAIhvk/Jno6/9NQwuARBGNQFjmqcprzCueU12NmyF4mhy
eBqBywMGoXTaHO6uNrc9efgDGcIfQoNhjj36jbWcWVLk2z9Rwa2mifzWTIGszdNt
ijydRSC8cJN7QdUtAwTqNILkAfv6ZI9clq2qbyusYKrll1M/AfpZkmnWE3f4h8ad
ht3xKOXysPyzmrtUJTnXLHIBXzWa22W7uIKdXR4DFhdtYDBWCfjImJkDnaoGcYuu
IE2CkvOwjjZHlZFQXZ+8ST2NoQ3ATduSPyfCj+UoCL/SZb6jXgMSJf+RlbRm8/Po
lBwzeEu3z6gLSH1AP4XPh2CuJgZ+tOhMtjAg8XyJiQrfYhqirE4oP6KLcBc2/Fru
XIxlra4+mrh+woxR2P3wPTpieo+gR8k2yKx/6Ncdm3hBsI2j7fHe7IZkKtwRgUhN
gLYYNyuIRlSdpo5K/2uQUAZxvApnKrhXsh126xUpSzuKCMYJL4b3g5u5p4020szt
YgwHulWstA2hWZSvDRuU1mz3IIdccSjP0yRhawESd/fBD2ZqRLefqHqprxPqXfan
SGstuJx0sbM6d7HprGVMeQfHo36hI2Q6qscqBTlRDyK8FTPm9JCB8UQjsoBEeA7g
LoHRpRt0kHGNJIexdBSY56xFMxpFU1t5eGJ86Ijm61qBxVvK8gNokB+8Jsv5r46V
AdWBNxQc6woRHWBCRD1VmeNaaSVWbJRD/TeWG6EdXWMncDRbx927/KT8QsZOEKAx
jN66GwRXr+AhOfvvEdvq30BntZvh8m3krJsoimjN3g040CC+X7nVW0TJ2R/RKauC
m8zDSz2TKp66gaAeuRznX7vf6SAFOIn3CrVwdlyzjPYi+XDEq8dvXZUcLwTeHtPd
Jae4tOcPfuYOpd7v12yvApl47/Q0kkXkGmW/ClyzhzI3fCDrQuWOCou9kcgXqOOn
Qg9CBRYMZoKZWIB5+mOPQoXzrugQdUezN0i5yXemcpxNjl156flauEx6PquTdSxS
07Db56TR7v9zzN1PY7+MBs3TyJF0cQvw6QdfGT/E5WTVZ+VPv8CbQBVqyx0hhYu0
3TpVYEUFWY4iKTe67fBR0vtvPdte23Auv2AeoFgsex2aH+OKTMeCNBO6w4poLibt
Qw1sok6vg4XYupOCdfttu6MOIUUPYKG5bP2wgIO56wMenRwIODk/XLyptdg6ORvn
NxXieJZS3u7jLlwHwbNYQhg1aEA6pamf9ze7h2s++4rh0FAhyN4/VAqKspsCcBB1
mONHDEBUFeqWFFrd0y3QxfvBiSgtEODHRMYPCppIXsjs8UPQai+UCRAYqEvnNe9p
Uo0XvkX+/SaraCFWTjY1oB1Djbb+v98XLpoPZIYyig6V0GAT3uZudT0JcTY28XNL
IyrfM5omMvtfbd78RL3zbE8H8KdopgP+UDE6rGkqws2exwxZ/sKd6a33Pv63Memy
LcFebzd5UObwLqGlaGvXHA3r0GtNTvvDorgxx2VIcAhLI/doC84ydnXmb0XI78W0
OScQkl31p9whCAmjr6i4Cdt0laq/ffKvk0v+1FOLF8yxCj8wti12j7IDKAvMGQVr
Aci8Uskg8fHAIBphzj2khWqnIa3eGCVFtJBWeSyFWaxYpOFw02Ecuz8KcHyUJkDj
sIk906S/juQlkhYz5s0U9CdYQS1K+m/XuJQdRpYlK/CQ3WUYWSxMM6/ZBprE/SOA
87ARh79lpfx2uQiZInnUrkklfqsWpF+/lFo1cRzT+GIgTZ2TzGoJHej2k/RSHaTV
1AVGabn6NzUeWgEXn5vzZNE+sgN2osBScnksI9wDJkdH0TG+PufNh7daJQ6JOM3a
8UnivBpOwRdHSdO4BjpLPSIfn+e5WrDzGYVj7AGsvW3Cv/b4GCiCyLkj+4o73XPO
SrNWo5MnvuSNPYdnbUv0lefMOla7o0u2ZhVDGmeGiX4Le5rxGo15eibOIh+1MuzL
02B0fNDFrMv7gVuuewVEN8lSskwZAPbNnlLK58Cxdnj4vims8CTXvdoVVaGdAy84
0qW5OW6DC93ffpvRIxX7u8SFJPVvlKLRst+13MzeRqW6JHzi/tK9e+8OieSO4/MA
Bm5lpcTocu3cTWBRZyuZgTU9nBLjuWEVpKNaZjv55QS1/KW9nobENWy0NSl4a8CV
Z4pPGFfF4CH2Si/DmZSlf8klX2/8UCRnc8YWSO/ilzhHeQVlU4tb6UaYKH+dGkPD
SI/3sUip1OKZtfZdfK6wNNawkXd2U++mc1SsCBlCs0FGVzb+cqmQWNki+bo174F5
YjVy5/X8ab4HHlsiuSD4Ek6BW/98wTzucQLKqdiVb3q5APZW/Wp9GF//t8nUtWDk
9VFZi67uHopVSCv94LE+89Z86M4w4YWSMRAgkTW4ZMWzqVAb2hY6Lm6+6Mb2oPGH
x8yeDF3ABjnMp3Ll3fk6G3AsdZyQ9rIK937jrUgYFu4wFccUhIAvBdHY8XBQLYEo
nGQh04VPlf5fO+6GLCW77NcEh+b+PEgvTcINls+Ob2SOD+WTwbS0X4c/5n1rfrO5
ycbban7szDPvQ3s/mYD4er7zXU+HdLnU3DBHB/dcP0NzuPeE5bJ5kC9or1kvEX5J
NFLMkJsHdv5x5BPQWb4GTeiGEOJvY8LK2UpUncPkgw/xrf5mqh58UIOew4hKlsUH
Jxtbnguc6pLGlnmvxOsqzXPTc3CJsYvhFyWBrHnSdj311d7E/KIPjb3xfS0iXKmd
zlPgd6GMydTlR2zORSfuPkVkbS/U17c1vFh1+dQUOex0RSo1xqB7YfLPeqIBw2/N
ArV1B1PM5vCAjyr+FSY5KyimnOkUbv8Kli0OiYgoDN50NLlnbVFX12xuIUxY3B88
hUIkNb+JSbXSSuGeB+uEmEZkFGRjfJiHkpmEIIMr4vsL0lso4AyD42I451dBiaJm
v3Cs5/I7KZ+H43zLwJH+N4bZjriI58zGw2K4ExUW8hQ8wIJbNlnC5ERCzCoxPH7h
h85vAUgDJYtKGnraI3mEYxLrriiXyYIhWA9auiEOvNXAsyk5gZ1lcuY81BxoGdis
9m0/0buPRf9Ya2l+3XQDmOumX5URR8nLA68Y3au82MsDuuk0TjwnHBJXA8U9jZGy
D2frTB+Kstlo82oQ6Cln32QYVSc6yjLVhAp2STmOK8o1DXvV8YfM9kBmIZf8INac
oWxW6YGLJvDDbX8T/LpD2I4mZCikQWRCPw+5aVKyT+9sqbPPObHqTe/OO/2aZ+vo
v3CICLgkw2XaKfZTnPWToH5pyLZrlF6klvnzU7Ag9U/qO8DvbL7TV79KnERuPf79
38MONDDr3LRDbZdzzjXIbstZB9xChd1k1/QmbqxnKiyjK9pwq650rjZifErJj9yb
NjrCo6OC1r52lO0QQ3p3E2xo2ohNiWiXDplNJVMJ/iuFwyTC9gJtF9ooJSDgTyqZ
mrq9iAjCapW3WD88w+EgZeSK0RSSrcHqI2FqfoPiuNBEdT3CDmFJM4PTUWeiqLpG
muac291k8U83kA9cHuhcxO3LIRuYOqT6j5Ji7HqR1hg7eSxYwtKlXBxL2k/tGwLO
ZeYXTypPpMWcB7D77yeoZ8t0oJQknCNx9BuxmWn8STltpWwavCYvZclMU90TlmIB
6Wwks5oQyiVWzSwWEqW+3/qUAhMXlwt0q23tzADEaaurSo479ul0Mp+Uyrw/tynl
8KXyKq/EDcNzBBBcs0oGd2MqnQaRl36XTvDelXzFWfKYf3eMLq9i2s4P23B4f1pC
QLa8cfOyI5ZDR6Ww2yW5ZfhgU4qdJSLcljCPSaDxwiRkEx97+nnAJNK6Dn/3gI0+
CCgaC3wNjzE3ET+g2Njw3JsMMUWJdujDlKcBxlM4KpyEcKvWj5Q02cy8IXDulfB4
ZceJXOCuclp6CMl5bB1MAzoWgSwjNjTWCcjXubDudD79nV9YxOh0lIFo8HLJuO+e
EGQjRWZNXwg/nZ+iJhd2/VbU3lYJQ4UNrGwYDZ4RFo1i/S0Om9cvsriTuUWQ4dyS
plNfJgGwqrvYaqzPDsAByNDhFg/uY48tKi6PNkWyiLYlsOwejzIBZEQ91gxsS59u
QWVH4hZzUQJjRUTTiB/p8/Owj/ml1/TIuc+hjTlssBDRGSxk/kzgPQqUvV686AzV
mEY+XkdsoSu5VpHh6A1h+y3VJ57MiuRKURpOb0N1geMesR230FHyBqdTx2MjGydj
PoxPwACAopM5ooN+Vqc3Z1PA2E96WEkY0kTVvOrhXWik/HfXhkYyGa/pgjV+WolT
kcKcH/GmWm575Y991dXAWDhfZZrhkyYZ9n9FqcRRaZifa89380TumjDmTNG9flfZ
Svbutd+4r9rNhZRBqKv6iydNXHX7OprTZV0ZRa0uBqIZSuGtvih64dA6uFpQfZ4P
NWWvOyDGl7SSYm34PQcI1HLj1l9fPOVJjTaIupUHiTAO1YWEN27NuDgqr54aoFlX
NWaW0t3E+ArBKlPwHg4YpeoewOGopFXYBMc4/iurtKE/Ie1Mr4v43ByKOTvxOZNX
on8zUT3YMkBERMu2tQZFs1JXGrBDE7gjimx7+TZ+YtwCuCFCOp9GxboRkBRGCCan
zye3CrZD12YY/OzNDV3PGgw9uJghDzq2+GjWfmtSEozDhUHGrfBBLx0rpO6XSuFJ
mHrEHFB1uj1OhD0dua6AQ9DTsTaWR9U/wmgZ9T//fofrKjgkVajGE1YwXrWh/bzl
vyc08641NGbueRGqAlKyLfXcE1XV5/5v8kP1uRqzKsTZySH6WujzNxQL+nuzUhY8
fxosKAzSABm8iI6WS710X4bDmviIAhWisuF3WDG+Z2NBQH4+PeWt6CzWa+g0Xev6
KaqTsaodoWh7YM4AM+WES66JTTlwyCUfVXEsiV6TT+mlgw/gJO0ZspsDfrfhU7Lt
0QAbVin4cng2EHHyUB3kmQ+sqt1QOLy3GqwzCp5MGzxiqjTD9ebDmA7QmdZtr+9f
4xdnCMMnOejZomLXoKbKFErAwMFo8wibm6KDy64ArjeN1zAfHICjfS55uokZPP/a
ctsItdUPmmFhS9KhZfsXbIkX/EptEpD33/EznpHBbAgAjF74FKoV71Iyfoh0sl3K
ejbK3Ot8Dga8+MN0nXDpLKI4oPc6rcROkoj8p+IsnIJ0DWYzA3Mniy3jBTGgESVI
0fgg0RxwEBhkihqeIaazjEbVVf52PETF8rJXOGshpUNeONtNflbxAmuuM6dQEgws
HoNdYWIfSHw1R58EEqyb5dyCvfjqAy4/Xah3T1GRKfF5yRSgl/szDW+tmfvTFmB8
zj3srHf8PBXwTcAjEStCACqtbPZaZ/ud3rT3PrxBUhsMKaC2ODOwGhM50W1OPq1R
OYfFjkbMQKX2rmMb+P9POC4DwDT1j6w1UGcckNdRKg1qaTtErDWFaskr9MB/brcN
V8xpdPr5/F19z/b4yAC4cJnCxvxi9ptsJbpGmm9z0GaYRi+NUi3Jm2Y7A6qItl3p
2OtPk2WtxpwbSe0CAwESFTegK90ugGvPhguYijEKRIXAngrCDBkujKGHzvHuFXn0
Y6pl1B2JWR4vrXS9jOEfrxSyOyVMX33yizQ+Xi4HGnvs81j6YARGjh8e0zpkL70i
AgLQMbtWr8bi5Kfacc6MQavV7xSgzG8Cg+NZYZ5wTjQdUsmW/KYn2W/RLlUZ1v3P
xB99E6ysD9EZ8Q2rZbkvm7a2cQ0CtTb5UWMY/AXQRW7BDsFn8+qHxzLOiHQ/rTRW
D7BPNa9irbyAN0APZjOHrHo3keFDxz+YPQas+BA3MsFpyKw/6OnrPzueUYbl675b
FXt9ZQbEowRouRTxXVO20dkHSmNF8ys6GiZROaGAr8ey9Do8H2vWkn/ardQpQJ+P
H4p3DcOKv7BrjieNPzVPOu86wwdgQEKBYEV7+EYrE4hLnV4lt6moulDfWEk6wRZc
7Wllb7/GWBCkUqGCuUMVndQKI+iZWJPxjivoE761F5uTL6TKbXBf3i7iYPivVsVG
TAeDNrutsRpnGghVV8D2UW4s83nhSpTFoOFlN0NNtuLdr2L2jtn5kduWYf/2VobN
ufgp7MtxaPBlhkCGsTrXxSuu16L7VbSvZNpIng80hlpm3L3P2+NZRP7fYXXD4ykx
7Mv16wuTbPuDKiVGf5hVsiTzJMw/KCbhW+kE9T3lfY9oJ2hg+WEMrHP6ZKCkqZg9
2FAq2HAjQfo7exRO92l4Zjx+5f4OXXQ4PuLhQQ3bhuaalrB96OVG3zjPyETV7OF+
gTVcyOF0sReqyWywBuK3tYEhodx6XdstTPjH7Zz9lesXLZNuNfFoGULuK4KYpUN0
T8IsoPPGqsj5L4W/8oIDyM7Byi2/bpusrU1I+zGZlIYI0B+G8KuZMSAVMALUNeP9
2IKFlcY8CI8izF4qt0JJITIYHXoH2J5ZljxT5qEG4Q2phoF7jvzLxr2uhvLulgZw
PG+hPU4K/zjvvYZcSwzhIw8rYgb39ZxB7QvdY26MzZnbEfuG9m/OTpJw31dkpfWW
tzuQMY1Kp2WZ5Q9KUociKpjPvA/7jtlkZndSy7pxD70WbkecP3UkibXJ5a21rkHu
s1NXShcbrwtt2LRL5lpK1EATdGuX8ifv3s87ANg2RIi8odXwFW5OL4ZF4QEQINwR
uw2hYhpqXo+6lZMvLwWRSQIfHJxwIZ+B0k7uKLJNzwgsQWKsbHBOAkavG9AJHq7m
ULcUEdIGiMIcZlK3JE+IlJTCYEL/okoPX9UO3r6z5yLmcOG8GeYhyLHAv7OsTl4b
YOLoIS3IHxS4ymjFNsfwayxjuQy99hwUP55+88BBsAP+i9lSLvkUTj9qSSr/H+6i
mgrrCYJdyL77jir+hR5D52BIeGR6eVYWegzVwB2kPCl+WP5qMG1yayBA/eKg/JUe
kluFweWJFyoql0wa4ZfZN2DJNlinEkG/V1bPm/xnAtk6edz99KA9gAUbmGXHV6Db
h1S9C9zQjds2IxrYVFLtsqQkEphvge0CHmjt80a023bf7rqcdjjwsoz7eecYEFOo
LR2AguUiDnsiI0KFk5NuAbnTLWQTCqrwnqtc5RpobUKZkfYIcT5zwXaecPUs8m49
6UWFhESIiGAxjFImXDXPWGksgNrnBqUrt+fAQgswBFNnkNIBHYJjvaessBJUvLfe
VZS0dr+87sYStLkdqHjZwRh54Fo8qkDdbftto4mY/rOoMMyZTGb8AOSnC7A0Y7ur
GhoNeB6fDkYpz64aobqlE2v1me+LIepTkat8O+KdPCcasnr1rMsGHHhcNVoWUJmU
DBKrrDYhz0qMbVDOGF8IBJD0chKGWQuiXcMX9CuoZQKmBcZCCFKQVlYjWG8PWpKx
7zow2Mj3ZGEVHB90fOnpmFdMw0LhqOt+vmG0nONgVo+3JnJ9K52wFWrfi8soD7H5
ROwfIVnbn6bRv7H0/xv+zxnulEfyWDOM3oyD+8Nv+y6mcFcn+RlEcoOec4vicVPU
1z055XuMdCcFRnn/M3pnufJyCehZRf5rW4f+ifU2MRQqfYLChDqutA4BgzgBY616
/qaZMPcjljxMh9Qt9gXgIL52MtOowUwPV6HD0qfTmRx8RsBgL0Vvka1mqrECss1a
2uA63OmcY26dWeJ/QoXtqIaH7MXRIYJ3R/2yMtvqehjO5TFGGZmJV4AwZknHQ7ye
Q745BDe7EAAiGRSr/jkV5hNg1KRdzS2X9+kG1pyeQsshOC5T/kyiVPH2U+BRaiSG
heauX0iRYsp5bh8UWeoP4tT8PspYwdU5J3bys7GJiAQvX6nzL5ReuVIdcTo1DrHU
bHYbSvpUiH49A2YXhAK3WLhyrjPpiuXTQ2KMKmFMjxkBBLk5bgAbSWSehhPvH23t
f0llSkBxdcYnqZ6HhSHCjHvYrEm+JxOwh02D2COkIWYR6iXeEuTmAFMypnjrKZ/l
PwLTaWuvB3vb09RzasPavbyjPeuBqCnv0Qtv+NxPjShnU4y/7lpAA6aCHG95x8bV
B4zNphQI1dhgjGrh+QKBdH0s5Zdjo8ngdiO0dGg3bXWK0J46CIx+HR//WwecL5EU
H4qbKFOhLGFzGeZ9dWhLqM3SPFZi1lN4Ri2BIYUwGk14Rvw0BL4L+stw+XJf3i+q
hV9IQz/4iS6R4xsnmVdFeXsSHl6uU/ylPl8ux66EwzKdkNWHXPTe7H/IXrNmOGQ1
3Dmkb4ITXu76R5dKE7KZsof2rCe6cdPNGZQGx86sn7UFvBFGeOuqfQ6ZOAyngo/l
R/lwge9BVxlBteI4DHx2mnvMTDZDIrol2FUYw9pPF7VBdGeY6utUQRqP2pFudYJ2
mS9HCFAEY1LWGjhjf2cb1pFFN33QFpzBHcfCiw9zfbgz6q+2OR6epdT0pt14Oci9
20rJVfWNlJrFQs8CAjkWkhL1G+H9uQ3omQqEhrmNicJkNQG7Nj8wPo2Z2nc9gqDN
FxPJprlLEG3L2g7zhmuX6DI7UFvyd+3aAA8i5QczZoNYs86I0eQcAt/tpQuSgzkQ
xFPfQjEi1qisRkrGWIx00Pcmw+ek9RpmIIanJEShcaLYIsCg/AsXFLwNZ5cubP+T
PzR7mITzKYQ03GbVJwqYofDzDKvKx4L7HaIeo1h/qhlTRLct3MeyB1te6rIOFnMl
NI7137UuUzPpXbtYojZn3hu7JxGo/ocAf2G8ko/eMyi8haT15qGG9Gc7Vq7ni+IF
NKuW7GkOgQSf4Z77ZJY0qUCMvMJlxNBdtvEgCXyvbDCykeTMlqxmUfV6E15ZMQXP
pVUgt60FluOtvMM+HFWCrkZ8kte23DNqTdEyE9s6rwXBBO5s8hso5anQkt4AVdZu
rt4qLFvY9FEKZPZ82e7ssZ/OvDy4XjttPMjEuV9PrbwN7d0xJSyQ8GF4QxC3gB+r
E9dz09/8XNa5JRkvuBw7EEGdQNgDI0/uYNgt7HYZ5QqqY2cSrAHOJliO4OsWYxOe
FR/IWUtvLsINmmh7dzbsuOSG6/j9bmQ0viQ4g4RUdPu5NKUF91+zhsk+HbDMx9Or
wyr4JlAGtJ9Z4/SEMGr0zEIMIJUL+kqGPxCnMBT6keOik9fAb5goEksu4RtOKL5s
W0WTynR2R3u0IZELlq1fEiccwtYmo/ZAIpOIuECznlXMIi8SMyWNklcuBfZry0wl
sZeJLFn75svtSFozjPLy3Vq7slO3CFMslZ5g7+G7c6kT7o/AbUu8zlvwv8vuvxV9
mCHuOsbw/8MSq6nvAeGq+6R/lTORS9Tj92ixTdFbGMhCGX8Y6IpddgMFXjhWwd58
riQ6oO/KliPEltMEMG+C0+TIKus81KPmqI3iQoRPapU3oPslexWDIb/ReataIrFz
OtzMwHX3oZxhI6oqoarTAhgj9Xw9ZEFWljskycvq0Xh0zrQGNyRG2Nmig+ZhJ6nj
QMteVgwtm5JaY+RdtrlemyZmk/QEb4MSc8WZplWj06JeFaQYw0gwEU5+XYW92jTM
z8EKnyDxuCIrGm+gARQKEBbacGTMvgK0RSOsFHi8NGLVzTxYtuKQ90osbG3m+//G
du7VsN2djjxlrvsIHY5v9HsPC7jnwIz+BGPLA1XpxOl3/OaPa426kTgLxIGZN9sO
1p1glJUKpwZbfjblUB3wnMVzmWMoPXDE0lrUNVFblV04D1zvzkLfL+yf7iP9veDt
9fexXQVjQK5hK5yN14+x3w8EFmKdIl4jvpVtFgh64nGgYFUyL6IZf5BTVg1Ep7M0
UGPfW9dENb8q6ZgHAnFuqS1iNbzL2ZVu1lOTcNa/TKhfj+p2TC7J8j/NLANwsqsN
i46Nw/8rWHHNaRL5y/DqaJQJHJVTdzmajNqrllTik7jt8LV0qAUzpR7uOUkY5z0S
JeyI4SjjDDl5k91XOcPUhP1Dl8kO88wfiq/55MfSQXq6hGIl1EiIuPTq5aVOKEnw
/6jGkUheE49JXDDEy+Z+MjyjVaxa75J8o6k5X42FegCFo+YnGCU39uPgbtm5nHuQ
OUf/7qFeE6ZwHlduOCKX7PH+Z+0brauEw8JD50G4x3hVLaSwjJ3f+T1ioaPF97PF
FIOGgL+/A5DC0CUWeYqCEv01M4vFgRG4airdeGUTcG0JSvA1vqsVAqAPBqzV86IC
KWvb3zHDDjfvwGalINETyN+Z4AEgWKHsRAYJKEPVCiGs0tJ0gy2Yxq3qk7KCIPUz
qEgZtkItYpxFTCNxG0dsZbX6OjuuLjvPG1b4Cm6/GGlDEKvJBJhet0xrFyyMlTeT
PHNFQSVVCxKLoSzQeop5joaVcWEG4yFyFEgwHpKTX7HoFMYTvkcZHipWox3C+7ja
QsWDPr1/i9L7Bjh9tISa0uzdH6+3s6O4RXheR2+uTTtIlrgghQ8xYobUSjiO/68i
6aiOSdY4LRTYXwReCBY1d9QRgNrh49zVhWIgEhjwHeuQUfGo/XaF8VDBVVZ1560i
POgGHwWLT3JjOSjrDr67taIgSQn8wTkbt122J3DUFRRn18ykV9ZxB3bPnN+L7JZL
5n0hEwF5fHTmrTRTJS7IMSplg8qPu4NMwwDJKHIghLoSRtfkGIuxSOBl2wBFv87I
OWfdjlGh9ETAPSbIFcWhMnhaP6+lMY/dHGb8YZHVImTFjp3wWf2hIo5zgG3jzDr8
vIi/efLk2JZcbQ4yEFIgjMJlWdHfdnHqwhooc77g7pGJMNv5/L6E8npTAkU0VRZk
PeqeFMCth+atu6CZeUOE18vW0Hzl7De0zsOOyWOTeBp04T624htxr/h+pI2NMVEl
Dr0eIyX4U7bAkoLnhUThjVvDO/2kceXUfgFUp1aBHnb0ltB4/vLPS5qUPz7ACF85
PtYPAqFoBEBcvAO5R5AUF6/dKidxqH9T6AYQBgjV3cKRMEKUd7kLKkZ0NfgsssG8
j9RLdY8noMHn7KigggYrRbfg5ZwvPFf6CVMHF89GaydomwzGwMMimOU7kSGFapmU
kXJ1zyAMwh3D29bzmAvX/wx+0XMqePqyli7OKQlnQEVsQqyymQVOOdPRAcVRR7EJ
vO8JtWhmt2Oxt5EgvvRdBbwtPBCG+IaEW3daFokCYKpLViJfLWv/IcE7wFZ80Rzw
1SKEUwc1Jj6VJ2HWXd+52VQ8QmeeJMPDk2nSWMP32VLu1LLljuGj9wJG8uNZNhZv
qm+VsKDFvXGSiNGIljJE8NR1+gQvCIcuB21MEAYtoPMqW067JIkz2qI6d+6HbXvm
pSeOwv/EaAOw/JAlXEU+qWn2NT96g5F4DgljlMMD1IGANAXyEL7K5u89KS542RkE
TfisgrDM4kdo6L4C3csKHhxAMzCg/Ui4rHCqV7Wu7okv0Mi0YIwQc2hK5hOlrpIk
2tOokLt6klnexfET2LWbFjooPWe18GsghDbj8EhClrnWhmeNxxsqcBX5VB8ukEGr
ct92QjyNOyzdrmDBdeT9kvAo7DR0UIBtQTeQhu5Ql9JGia5RKFg89Rs3KegyFCbD
Ob6/3OL47gYqhfrsSw80dJo+a0gJqzoDDKRuazLfF+/Jd8z5PQz3p87lrQNN8qF/
gzdT8UN6uTf6KjxDCIoCToz13YB+iOOEPKVXN0R6sZ2PojB9/eC4oIEnu5oF8kKi
CoZWx33T6nv8yxe9u8654vB6LmNWiF9j0bIBFhiJy2QT0SxqJKRPikDRG3qawIDL
hgshf+ZiidXgnftvEw9IywsUh0avCK+PelL2cJra+IiyfoBVbyLB1C8EBaBz9VHe
ujg6bh2jA/Spf9z9RVjAlbymkUPN0Kt54gNSL8uhJqz4pSYofOIOzP94EykaqmWc
8cnyyUgfjqTFRtXewSUYvQ0pzyAvM3N4wbgvPcTlvqU0vgc03OJASAuGwsBDmeAW
RUVMQNUZeAxeDwn+O0RXQY2IaNU1UHjd6iwwzQoG5k2kJLxRvJPTraIwcetsMSgv
X1oQYB4/8yfPlju1LmxoZjYJFyUPbejiPpePGF9Yk2q39uLFCIIjR+S29LclsT9D
RI6rF0AHe5BEi4LH5gLpxp0FzeF+bOPSjXl6WZzYYtv83y+IlJsCOItQHOZCCcZE
qk9rnFmSiHkmUHAjz4VHefknh6xIxA8crSEYboAt3vqZNtyyhJkC6nXtd2Pz4K91
7Cmg8RWFqwC9Vu6JUcCys4HJimm3HBz/hFQfNM8oYG9j2ArZb5IsF7PlX7N4iTST
BctRpzt3KcGpyR/rdDqpBPE9vFhBvn56P2Yv4zdbB5JFH5LxGi9fOQhFzLren/+Q
o1BsOLdHLAkH7TkZanfUrJ/tgBWmGLMXiw+0IXrBhynvhqVGiMFm+x6ffS3NmHmS
vb6KfnO5lLuj7aUWtrLacU5803uHmfNIhPJeUW3NG+lfbRhCciUfaxh/fc3xhE+E
kym1IHXpYhKffaW7FtjC9EwMNLoJ/eBxVPkUEMZtv3IYWyxdwAto4Dh533qHrwTA
7y9KBQ+9MVGdxVdaqMlcttuSYtebbABDzR2jeTEM1rxOrp8GWK+aP97cYIX6o+OC
ne3b+IiWvL7353MDN9iTK4SlCfSOydMmE4DC6GxvCTzFKbU3NIy73gN/3DnvZ1qN
LFxT6tziCUTszh4qsrkQEBAYeaU59TDzn6lVT0AWkLEf1IywENwITVrZKY5WjWl7
60XYJo5MtdQsBoDcqzY889itKtY5ln5X3/6uyW9eOC1gRsG/kU9SkFkrCZQ2KYt9
oGr8e6ZMx7Sdbc3o5cNThTyWlszBPD+K9+uBXu6YBL0FpfZZYtdsA73wumJNz5Q7
pQPdW8/w4FwKZCffa/5lvqe43DyyD5oKBOBNTfxJ+pz5VhLLazlr2IUooklTU/Qn
U8zwnOBaIh0lp6piJnupm3lHYYZjB1kVKEJEg1RgTWzkdwgOmMjBYVnEvYT09W4A
EcsqEr+AIT/G/z+VHQ1SJbWJ/4O1Uj0GZZbrk+4WpGvTHcVjiI0tkChR7LaXhgiX
ROjBnVeKCtr2zPYhFte1NJzRgMO4Hi/7gTL7UemHryvsgBMe3r6klXlULR2KNEc5
CScHTREIwqnv0Ce8v+J1d9H6Pui3dNlenq3CubCTZpY8xDQDQ/6/H/G2HJOfYv5i
5+H7pdchAlG4s2uNFuBaoQvVA4c38TzLXA9LNyWfm2tdWrXdyeP7kQygR1yiSNLg
ZDStKO+n23byMJ3ZM0hm/3p9LJMa7gxbn4yfsjt0eCjGUtYi1qpPr7K2v6nb00dh
OrRqSZZpPQxMLqjDd3/p6/8M6FHNAJJKjREXjZvIK0M2vBuEVHUQWY8QbFVzo1dz
fGQDxfhO16YWNuUkK9Pobw/WQDMxpyMDejZM8WlxCBHKmzn04EmPO7GjQtTZ4hVj
Gc4B8nqp+JfHU8UMoYeQ+DFqW/tow+7+MKR6Z/8KUyRlEchprcBNOJUGRYMBofbO
N5IOgjE3M8DL8XXJJwop491fRKtYBLX+yzclLRBX3wa9DA41r9qw+xphT679JOZM
U+2u5m6LY0T3zRI+6s4mErA4n1LqhXpPhettEVfdrDbx/SyOJb9o6v1VEOym3zCx
aVpMQ1/GOsbrDJ1pQ6EDR87vfsJFk1g/9xnNEioGXRxCNSefBFL3Zogn3AJoNZdO
go4a3xVWYo8iK7zpqR78uuUchi9qcubTiS5wePVPVkBUlhm2Nnezd9ICSoKfRdlO
J8RqGTeZ18xBulSBywLNpoKf0xEgvVsRn7+b9UHajY2KDQlfFLhyfz5CEFK3SNzb
/OoQVzqI/BYKtDnTi/FxkhnYoVVn3vO0NKUUtS12OxiQDj9vNT3jxgy6nAB+r5L4
Hd5XuOuE3Mo6/QkwaF7MIK3af7J4IJ0kNKBYBxB/jM7nGc5fnKwcIVJ3x/vSw/E+
1bTqSc+pxSW26rc8Dr3ILhDj/yP5lUnXE22CPZiTxZAn4H5ux371nTIyIpoHUOPS
R8ynh4FtzSxLQRlIcpaES44fSniplK2MVkgPlwUXgADxcinr7U39d/C+B4H9G+54
UrfCKnmr56Ls/Hj/XCYkGXvjVGBvxlZ9II5p9UlG9HclPfqh7N/7Lbr9+kvCU2bX
EcKAr81Z9ZxQR0w8ZbYrcwd6DwfwswEmgzSVfdT/Z+73F4l+rmMppBV5k3z1aAev
IcsxD2yadvG4UFDpGHdcT3FBV2ZP4q6QX9CQhC488TAzCzphxtSOgrfCYOHZxJFB
iNTHv8iatvSbXJzKn3H1Hcgf7DgGSLoYsiWWCGa/pAihA/zOp7V7/y03zpY14mlO
mbl+Rjhui4YqISPFpo75B5O0UrfTuHcSinQikRm5VAZd5qxVJDUm4Eb95hzeUMpC
DwzapuRsz6f6mbgCS1En2KZRp7kYan5KNfKdaakD5WxEcuDKwr6dyWGCYCxCyVof
yafEY0CuNNtkP0ZTVOmtEMbf/y2OClR97FZfmY5QtKnvV+KFo6e09D3VkDfAUEuO
wpL0g/KxTul9KcIkpuJl7JidntuW3PleS3kdkz0A0b0lPx+gDkzkMHuqCQXMRt3O
FU8fDNFss5htvRHKkxB8qf1Z4xJ2o3YxKlgiZgch7y/5lI+/5RfIQP2aIg249Ork
qf+FdUjkCzvwJvlSolqkxPHLIf4bW2dHMbFnBdcUIwiErbYjpOU9W7L6+bs8WXTg
/0ZYq7zUCDCTdywN2rypcP72HYOB3ZfxcNz8gf0hrkgWOLBkxphMGMHUBa8/St11
n2IJ92JDSpWLWNZ6n+L0GlzCJ7ERDtHP98Gawj1j4dPkakcLXdOa8OT0lCRTdhZA
f4xNPics0Z7mcdsdn5/cT1l48bU0/w/kdnyWIvj/aDb5idvoz3zipDvTQunokYcs
DQn26wtvw70gmAJVpbaYU9bZNzdtqcB3n0Ygg1ZkKpFWMg7NGkIJEzrWD3MB5+KS
p7Eu8WKt1pgCxC4HOWM3JNspQhSr2aDXCBT8WpS5x0fGEtXXRFZMXCTV4KIysdkW
yA/F76pll3ehwB8lTY0GnBlEhzOzcxqopuEtDVxIK4y+haOWBIJIgFxIzJFXqOiV
r+gGu3EBhQ/MWCAKORB/EBnvTePvDCMAoSJ3tjiQ7cC84bUsEwzSdlnOyrwKGLJ7
U02YehEiFHO9clQIX9qZoee8vsnqDWJXCptkRQsTl0O4XTZKfLMkb8M8hW+NpdW1
NUyRbbCLXkr3TWx4JxWPWhc7Z84aFRAJj1XCFT4dnFp3SxbMq/FQPSh408oHBXx8
G7Q2yof7OqE3uPXywZ9JFp/q3IwnFuHsdcjLC5gh2Cm4mZYLuIjEsPCuEhj+UaPi
uL7+xhCnR0NaWMSwKrYP6Em+DKEN1MzFqsYrKVJpv+RK7HI9locOn66NPWTkgidg
5CoFRCHBjxp9J9NW6lvUZxOy4dTDhRJbWIAp1cnCmWYaWSGx2T5W30kzyNaqiG53
0ZBXZDIkH18NjVZ59eTmzb4WnQxWrCWr/Fda97ya+tsqYJettfnTKlEPHSuLYbwJ
Uf+Dcb2SSbNxWENeFLL3EhasbNtYG8P2lmkeoDK7+oz3YZ5kIzDOG3zzkdjmmjV8
YtaYUQCjTvcBoFoRFGhGC2ltXOriWrvXpynxiN6Pz6AMtDLizPPZK3iNzE3/ayZ1
NgPq1hXdZdjJFr44scXZOJIlJUUDP7oTQhK6W20XjFkVBuvzeCd+n0ZweIxqxDpA
FPWzdujMl7Cdr+yMRevWAxLQaRiXvizN3Tj5tfTKWMk8EVlDYss2YiQneKp2dawH
2c7O9qUUvTBKeUhIYrBfwC4Oz2XYCHQ1PnqxVW0b6roW9bpJmkSnf7HSPbpkjIBh
aK+lJ0lCGr3RIr89gg9iWKqWplmlJqaV7geFC2G8eQJ/kJowt7SigNOcGleQcKrA
vkB4Kg0mwggLw3B+QwgTlpcTTwkSr1irp2QQqYXzdDvhiPDnkb3MswJGFsG+dxxg
Hl0QVPjJoKxLrcJEWhRyZ3CrsCeJoCaccwyRbWVuqyFU2qCKsTlN1r7BJ7e2B6to
Vk5HJ58fKzoG6vQrB6srtHLq4jgEctQaU2z/kntz0ILQab0Tk5yyAyMtEhpdetQ0
eCmm7+mgpE3XAUlJ5fSAEQ6Vk9zAkO4GP7XSrKosca2OmZO11oiZLQQaJat2yAt4
9eGx2bPDgnKwNwFGVuxOhI2z9gRzIiQDZfpb5c3krZICfXUQSYHNT1Gd22Z0DPnO
wcinklpCufBE395vTAfRZ6tJWsJpFYZbLBi6LIpHsMvkW9+ZzxMHXRfjF05sTBeG
3k9QUngliQZLAbmI65wu7jh8MpnPlKM7Xg1SfMq5UXJQUYB/QoJv7MOKgNriSI4k
Wbi1Cgi2ja+6G+P/egFD7QQo1H+9xw7MO9yCyMyFO86zFnhFa4uxBybZkCD7ErvP
A8QBcALagYr1+3sZWRFOEoTEaZDr0Hf24v6JEUI3Y8gElyWyfZJgwmLrfWxHthar
P9eOqa3qqpipuzUrY7WTEU6LLUFgS+rCLgxfjemh9S1w46h0aTsvXRlZfokJ+OTG
WqemLumQZWluDR20gX2AlzleRKR5OJsAlHiDt1Z2wBS1mJeIKhmSbqMh4EEuT942
3OdHFHlMEfSBVjPzvJwiRJUbSKbXNgzkIYGsHchN9AU87xQ2pIv2KXrvzlJyBsEi
fD8cA1GGwg7owoH/TjWTGhMs+SJys/xxqgaTkCu9VTyRAE3QjlNZg9dP+H0aTyNl
jGKcMjQ4ptLDxoVnvh3CFH4k57WjpAytChrLVPp0MWeW3KTNb5WXsMGLqaxna1T9
MAL7prxldG2drUUzBPrmJNVVxTXhBx802f3wP0NCpeNLVfy+K6bLWr4kFsrXPT3C
/1juZXiHezCC6hgIkb1+de6FtpVNelRNvd0xOk86Yg/vc0cDTkjbnOBh96N8aY0Q
AORu2Py53jZrctOe+WHBoPU9B9Sqn6jlcUL+Impyd2+eZF/x5UMXMwPjC9LJ+IeH
44XEkMzBH/oihTRP0+JGgI3dKNlasfKYWsWuidjLHMu4F08yPB/EJXNr8rmv2c1x
9SOwX86NGA4hZw4oHPuaIW+7t7rvEqW/6yalLLL89TE2JSDOb6nTlf6QoVP5jwyZ
YCRTQ+j6Y9CsY5eCfmGLaL52kNSMqNvUlCHiZyV9XE4vHhFHZHuUDY3qnNn6dePR
UTvtDhjogyM61K6oyJ+8aAKd7NLPoXN7XBMGlmYRslJTppulF5gIoYnYCUr6MZ3n
/PnOcBdG1GG6ts5gag1v0tDvLNpQGLnAlZFyI1wxRoAUV7Oief/fAzrli6Bmy7gx
1EMym01SiWazHrAc/WiWRIp8nLAxi+ff1YJNKRNXhgEE4YuB1cpSBtIb4czxfxnH
RXaQaVwvcRv9oYrvl4e9ApC3FhiFakTGzYDDHZj9Y16h35of9JLgc+RCLZ8sBre9
glmDBc3GD8mW6Bv2eElt9ZgjrJ2bEh3a4kr+Ok7NRS6S5+djq7mSzDDhPH/hQDVL
FlXgCqfeKcxudwwtzehe74AX4XxL2+514HJjFJHxHo9r1lKzBZwVcQp8sD6DXXbM
FT6xNxJ3CzgwXIkLBbpIt1OFnRQbfHm2N9m2N6VkSktyKongfGCq5kUxRqaNwpO9
7Vgk9fJpO1VHPfc24H+eZeKMNEI0bJgG7883Np2GKYJxMnTCTNDofEoVNpDAkYqn
u4/6J+tWVWpj/eW7IKE60ddmnQIK4oTmrzxtYNZekhPCK7IncVYYkeOR3nAsa1PS
qArfiRP95sxqpCArLp+imV9rdyiACO8R2vRQIWn2WTpjqzWnA+U/zyoGwsTDAlf1
HJArJF4vVFqk0uncazdGMzry8fD2CQnj4ApW2nA5rZ39/Cjph3kruBgWoJEVvVDu
nvD8kyms4Z3WdvJele6CIBWYbOLJYN2ahUyrsUKeC+5dI+nhy/vksJr55Ey0NMpr
6c3WsfzmmQLGIrZfh0/CKpyoWPauyiVMv7oIargbet6JXfUgXVt6LXh6FOdi37Dg
r9qh4f+Jch1qormYj8FafH9ksg38J5AZuUEJixRkFhT/RmZbLnj2SyKHKQIEmXXA
8Utn9gPcC4m4wb5lOrBpgrXf/UEjTmpxVeNHdBQQh/j9A2wquIv7hIyEmh9FKgVV
qmp02g7VMkjOuxlj4HGC9zO987cWhFgBbxRexuvR6+nfAoNzkgzyAjV6iVhGVuft
3Mv5zeeT9O+xv6P5GNpzIQASgWY44N4oPELO7RdeyPf+xZX2qponE5Dwr5iE9yww
jdPOzLMozZThz6B/zNHDkhJJSbQclTaJtZ0islIKmQ+lbhI2MOPEEOlxR/RQkBNt
JcFkakmUCs1yFdKp3PsPH9vWrlRVQ5BFDZl1kGFTGesHIDcYanJ2muwch+ijcDNu
AY1drmHxJBJZsrlTju5YHNjZexxqpyfeNSl2u+eNGTzS//+tFxfhS3f/GHslLPom
GdciNDdjSMNQRN9K70wAJbygNCtVTv/JdcLXHVH19aFwuI4JYn91ku8qv0zeE4Mc
SReurKNc8gDamAexNbsFuIEDDhsOPYlZw6qqagH5Fhjtrv7CosoM6MtRvIhNw26k
jMnXS0x4BtFGSMSi/14CK9qpyz59njt8mTSRuv0Cv59S/yZ6/sXEv9CQIrzmjL+Q
FIiLYL0afCORt3OrZLFkbu9kPmlWUbLrpkTI7ZQSTUDkgnrP9LT5lUQFs6z/Q2ay
HIUPajO4AgImOHwQLmiM3DoHakr5I1YDqG83HDAOS/8KWCEO6CR5+imSFeAvzeif
aYxOGQ92u0ik/PcHQ4T8CoQQdGxU17s/jgw22Dmg/j/X3ag2eY56Mkt1wDs5zx08
NxGsDz8rERbzga0dBWaWJCF0wXa+KI5Fmlo4UcuQ81UwWa1HI2wDdPjFYXyHnCbr
t00PZRFOL7lCejmbjcjQF1fZTefJCU/3u7UuKaIvSvhDxVFSx8ik4hbo8A7mr8z9
ul4XI8SZZFAMrnqR9nw9E+3pdORQVycvZQgtX1ud/zpX23rMkM90vDu/ywmTvAly
lrllgwffHEqEsZd/a3gx8yQG+USQr8aBj3/10OvgufLbcBR8Uhj0j2/C5pq5PHz/
5QKQOF+pRDYJhr5hUxxzsAX8PgfW9ZCG94cdP9L0ecXwmhGk0dN4Ef8KstLwWjhG
o0mLfuCkkz92XeoLAEqEErLzWTbnnzxpDoW3iNP9TgEv9hl6WfNYNtQv/0ahikmj
rZBEicO7aVKAT1IjJplM/DR1hi/1pls7NtZkPyxCOz2QuPATYirpWhj7hyrXqQRS
TSLaZH7jYN22Fd7eLTxr1FR/GAS+wjKwRi2EOouV8ekvl4ih894/bD4LIpA9zaE+
JWGLuASda3+4JwtJTh+pustH2VMPLmXArcJP2/i9+lM5obWLWtUcMceGr5JoEynj
63aNeran0zk845gZ4MbGTC/opInr83sg9LQofMv6hEex/lA+8oZ+t5TtyyCuaX2g
m9ybsqQNGLP+zVU+HP//i4B58nOz3y4yrTuThDo7Q8jPXiA0Tzzp3CiB1/n0uG9I
2zxK2X7HMVuvw0IWaWXALcV2gAt/rBh1niXhVZGlU9zWgelEfHvsxXLcD5KHvCZp
ViBwtgM33bVk/KSVaFhDURV0Nrj6XerBsCLYLtSGQ/dBA0P7xoTCWMh2SSIe9WbX
+hNqYsWMJ/8HLcLWp0pTmoNjRg9iZH34OMPSgHAQlRxyIfHX7LRCNxhubYXkCvRB
Rr44h8paJrgU9e/OsuKgQnLURGadpqzb/2VetPjtH2EKocWRyuYWgbvfCRpCXuh8
ha5Uor5wYAe1njZ4mxCYvTLGuwYNaJdAazGdIc4/OjwzUaDTsgSPdlxYJk38O9wS
2SJ5+e/tM5ihhoPY+mblAqYOVW7I1DsjNpcrie6Kh3sDjBMp6tk2Hv8U5+3DwLXJ
jVtCdnfRXZhM9r5mdFM2JgEZkZ4AsoV/EDjqncf2bPe5RUvA8XSbvRsZJsPVr4vr
mvtpfN+dikEOuvULL/gIlGYUA1QaFxLkq8IwQ1wFIqVS2c004c5Pgd1x1GjUggnr
HyXisnyu3o0easv/SUz3hA1h1S3EtEUiQGXmPaZdYfXXjrg+9WRhMIy402LJSt2Q
INPAfQvIpXzQDC8NoHv0LUiajf22jTvR0IbOFLFEgVCKQALlRLUEcMkFJM4pfFIq
XrLjD/EW6+aXlEv4sF3mhEe/k5LJrdenduxSzF/9utWBYq2efg6kiHEfJAbhhtmN
+bsdXQzJAg6o84P33M+u08VfF0hdYZbv//HXfDnKmsZiLTv8sobJG8pokmx0SCJV
/mySM0hfsyWm1debgod56nFsnTP87tfvTWnhPj555E7gqGQKiAj8y/LlgU/fgoGx
DnDRpJXkPvIR6MvmPPfSJi5+39MKEPkhwTXJNYg1Sk10BI7mbx5tb2IHnKsGGeMj
U1jJ2FtpfQ45E6SE3B89l9zesy1sq5bWQ5/M2GheY4IiNKxqyLohEab99WzZjaey
pRTKb9Y0wxnl0q8spQgXTzlJJoflRVly64Dfs540NOo7QbZA0e4g1SJ73asrXKD0
A7UF0iuL5vySnXEGS7wDUl1lAz2gPanCKkLUOoQYmcs0MB3Ckd6a9JpczcCJr0t3
D0hQOTQ2oFG4T02o2OP74NenW6oBfSVk3XDGds2BYUgIx3NJM8hHdLddH3S46FhM
mtUW/HP5tR5Omh4VbiurC7GixBDkdcfejYiKnNVIO2c=
`protect END_PROTECTED
