`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IwFYRVuo5AQz7OrgZtGndtJMNJCRpjA3Ps3Lc74gQBp6gGJx7MS/7GLlHKGNqzHl
38od2KMpW3ShifFsFchS27ceW4ga4MfQGSxkURfj8YPd0E/D3sC1ds8KkywwIjyJ
30dqmQ8M3khcDSL82QY9KXiCO/KQvsA8VbFhveHpruqXnVCK/vrjeqK/ZlsGQF7b
e5y/jRzAW2PXMO6HyDyFnS6T5gaeEPiAzsIp/Tlz9pZ5Wb4sgG4/mrAJ6qVbSQgI
VkYEw0/OY4AhudS1ZBZn0w91GRwuAUMYhV1+/TwPxnwZO21Fhpno9SeOX9cr8SnU
sy1Z8ImsQT3PtuKFaJGvhn6M5xXLNr3dLg2ph6BWHuplk78/xkrWUvSRJzQihaBG
ytw5QiIfCocaVchY5nU26NwyzlJfmyDVvYwGC747M7wAZ/UGmVuON19k4dViMAT2
72KW61lOFKBUz3U1ITVw4eXfAxYopExqxU8DnF4uqPWkHilu7XPT1uCMEKzSl34B
wnzb8YAoSc5Cqq+/2FOhDs79uBzDOqv7N6DoWuBkk1H2XdI9j2baSZcd2BEqe7Yt
1iwNq7IJGUO06q/FumFWQQNm+QdJ26zcoB6l8UrN/5CDIkNGLRzfPWryp3AHtJvR
W8bNNnB67K9dTsyWBPh667cT/QEb5zV1nx9ePTzuy3tr6QEQ5vhrTwQRBKetQX6Z
DAJ5+D00WDqEQORt1nFj6t/8pP2rLds48ge5gIAkJLML7WRpp60uBP8IlXYVh+Yh
OYqOkflsfNUrMeG1BXm56A==
`protect END_PROTECTED
