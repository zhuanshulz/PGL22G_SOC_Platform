`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YOTFSkKatiOnydM8aTKvQJx6GHcaPUM5C1MNxE/jGN8X72ibLaCC1vxWO+Pm03Z2
Oto5mW6Uyf/2udWdrMJZp4APK11d0C2PSiIl79g23YZvjQmCd77vemLGR1nzQ+LR
ddRtUdO3mNYAqpr3oyX2ZWr+bzc6QqhsnzVlh4UUs78K5HVBiJIZolxwE8JuefWU
8tmyGOd6/qFUeI4qDiR8hMm9Ypt0SY2yregNrg1TJKAhsWw2bzQIMieHMo8tOfK6
AUn+kH6JgwjuDiPYIhA9vI3k+F1NDq3TqabypqBnS2ucBam0Yotk5ts7ngaVC10V
QIkXvUEORo2fjWMEWzo4CalosYoLPwHwAFNLMTHlLOW6Dgg5W7j6gMMWOJEaBFxc
x0ahhbqXxTwN6mYUiIYD6iobZ14mWmzFpag1EOo3X67fob5VAnpfhXYl5DJsM1Ek
0FjJsFzN4rmOBviSfdDNZBR9xTrqpG7Xu677PYThuLVyKuBlZXbQ+lwmlgmG7+BI
olWU6/DMrYa+r1j/ZQ+1yPz6/RUub9pAqrKQGBj0+95xOFAOZdWRGpP6yCq97bHI
+9qAsS4vdQu4vMDz+/yd22JvLgwGEF/2SqmQNcw1ZQdmX0wUfNTjvBATghFroOFa
I7v4AvDPyowKK4L1nUCGT3E+dQotIVONNvq0NiyPKHXhz7buJ+/iFHbl+I+bGqrU
i6QajE4R8cgnQlX+rgw1n5oojl9Xcb1sPzDki6UO9G5aReEqZ5iHLyGnuowXYheq
`protect END_PROTECTED
