`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8JBXvlx5mA+iaE7qtgFY8fbEvUyCamVBJjQE0HpuqOhk+zEwbxEvSqJ/Bmv6I+Gs
uQSSRdF6Cx7OGhB0TgXN3dp+Lh9LqbGDyIMd1F4pa6IQaH8vK/kgAp6qBhSqja3V
G92Szau2pSudXiOfPlI7fxOfxT8I0TBJJhETsGBWl7R7JELlTsnheq/4862J6t2T
/bfEKlr0ha1+3fWAjdPYpdc6CDtmBIEcLQ0yiY9xrlWRZUZFHaB9hISaxvZWi8mW
nvJO/YmUGNJ0/9QWHQHPUZGG7S0lawapxL0hIr/C8SYUeGj2G/qFn+wS6eb0wgPl
WiuUa2OVPtFxXh3Mz594IWA20m+VAc+9ICS7pNXBFyRBsubHYYmZyJBBQ1baAdMn
i/zYKjkQsbJF3ZGmmBKJ7DZV0+NKW0+/N/fRwG3je+Il9grHrZDay6xyVhykXjCO
FvblqniGdmqvKSBvvloHehoMtJn5g3l20NtVj5FdzBPIOZkNfSVsjUNV4+0lFn6L
CQ/p/HgQ1mUQLNxtnAFYLv6MqcVz0k8Vea6xumA9/QKalW0YF65hbff75AmgRx9n
ajxlZEMzMEyG3Ni0Bt3oAkfa1secRWjOr9rqqJjpd2p6gfBLhrtPZu6n1MKeprzA
fiBCm/LsDboNnV11qyMJdoGl8wWMnmtM+R5vq4NYOP36LAe/nuw423YJFnVhV0rX
6ZcmoHB63bYW7Uea1FbE1BJycGqmcyISgv4t5dwRx2E8dxvlpD03X6PA9LCb5y+H
D1Kub5PncOQMb8mPd/3EgsHrSsvcQ+iTZmgS/3VtYVnTAdhfKTYKbaLhxqbdRG28
GWPH11qHlQnHK4Pf3O7a790ihxvtFKMT3Mwf6jCePs/fhhQvyUmRAqfgktrb6iP2
HLdjok8bcxWs1vCeiOleunmxy7Q7lbT77N+MNyxTaBsUO4JpuktcPU23kWS1Nb7R
zH6+q/V9w2iXjgol9jcLUq9B0BFSAekg+r1ciEBO4WnlpPmyqWzatEyEqgMjFkMX
773MeR+YZ/lE2jE+0FWxzUNUey7vulpnjcnpJucrkP4=
`protect END_PROTECTED
