`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Lh7Qk+mPgGrkkL8bud2KVfhfJfV8EZCOz8Dr5tu1vaRA6OzgVwtjWX8afRYGa6iU
+Vmd5WnxR/c5iKI0dMw2a9VbfEkJv/1YMxn/HaXFHeWBm8o/1XtZWMQw6OZqeRvI
9UdCc+c+NNIjEueYUvHScg5ok/t+gxwH8SY8M6/tRlf+mfbr9ar8ZZ/VDP2FWxuy
Upu7fpy2MHN35PQzLEqFr+n1oiAmsv3Sqc5MSOdmp3+BJZeESs6kbUXWWQvkBeX2
ss9tQjzMNsJ1xvLj+srTwFHLpb/HQJtEKcxIES4uW13eTllyGbZ3JH/3uwwkftlS
yoFiM8P4Wij9okKc4fTHLkyNZ9xCiz/FejwWG3W0J0FPO16WJIsYGN48aXE6pzW3
aVYcQPoHX3oPgKhXHpe3kcs6txJiK1rBmUqEHMfkM0QZsywBetodcYDK2d/aRt0v
AHviPr2FcgUdY1DtEcVd3N+SOV80ATw4J+FtjpMEHsb9h3XnXfd+laZxqV6uQMQg
9aogNsyiFbBO+rdPKqlVoq7CERNxyfgmMo72gyR179RaZGH9rcFoCMdGmRqTlYU2
QgXtbuMjzzQCNpwPIzekUsU+z+01CINQzXFIsuX2KoX0jO/dzO1YOpR4OMsB6TMv
htLaGh/Q7nExQIaI1R0ezCdNzydR0S+22sG0l4ASIlFwsIcuOlePlDDwk6AxhUet
OIUNQnpYp7HQoHP40vQTcBnfOaLtXjh1UxTn+SKS9QgBAT6XIKOom7dqdUSlq85Q
WBGadVYhnz9oHQHnOzXvLBAt4tebJMhC9jW5SvDkWHL7UPvclviH0OQRVAslsSLK
zMk+cDP1USEYNa+KxcP3hnQXfAML3uD1AyixEo7gUE7sI0IZsBNPuLyl7ZHnDSwC
bw/cHwRk4W1mmZGzGJVX6H+JX+qiV+mbcSXDXYsgTIyKGjgpBilMkgEhZDBGXtPf
jVc30E/FOh55yNimffQVVg==
`protect END_PROTECTED
