`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wIZwYXqHuc0CvpDrEch4CUqPagcZ7gHYgdXUB0yyqTgg9DWS632DuKQJ6F2UwX8h
UvB4GroUG4ZzZrfIYCMKrcEG/x2zOUYzOGeeyRpHYz6wUqEIqxc14A7lYAtjXQNO
uuUwv3rJu0qNw7lWBQOmfVEGqXKTx3LVK1/cCpYuE3DQVaLSTtV0sLjlrtifTEPQ
YjyJQDxn0YFxclYNQl8RDjV7y3t0Untes0nnXcqcSZ3ow9y+97Nm3FVkA7ByQD6c
G+uUtp6SIXjkWkZVOOvR/6btnuf+euazgT1xrd2ttfGz/FgzYiafd2m+TVSBldVn
+TBzMGxHuO9+nQ+ThTJpOsyc8fCxcl5xRmMs9cAmYlwozFuI8BjXss6D0kPeQ1fa
SaMYKvNCV5WzIkSCXJLGU/PQFfXIrZz9yhxjTOIboI8=
`protect END_PROTECTED
