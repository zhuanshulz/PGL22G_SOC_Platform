`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3ecGCZyShrGISjoAcjOCqGyR0Ig1fjcO3wyAvzfR9Lq2eged11a1k2UB1EyxIfAy
UAWlX3IwxvRskTCoZfQZQwfJnmiJiB4K8V4GlG3htGAQOgmG319Nhflt9vpiKLWP
zCjAqGoftGE2zE3kC2gSMGXoB/zaH8aE1F+V8kOOkn7JUI8iHcBk1WD57Zezk3Df
Udwbw+7Ry+3llIDWm3Fcd5TsMltxLDnFarlQ2COySprF3xN96HIHVGMjwuJSCAfl
WVxREspHOo4efbjEz9IcN8C7oF5rc/XAuXnLaWZNrTGxdXpReh9eC+hkJY1W70q/
PhUGWCup+Pv5hH0t3zCFWa9S1um4A1gEkK5xg2fk2nFHCYhCWktoxdUOgJOEdWNi
TT/76ca6I0zdYjocw8IjmRSI8cDiziEhj6NWG5RE6CFx0mWAgMcLXCU2esrdY+IL
jPE3xIrkiWVm25q99co0cgmUHmJ6Oy/pjiGJIWlB8OmE8EwE30YYCUKyx/PsX0xm
naLLmdScAJCknSJnE0ZWag==
`protect END_PROTECTED
