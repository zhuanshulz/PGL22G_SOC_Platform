`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SixxJ3+9abprEUIwLxOQasQoeQiAo2EDGOA4o9+MgvlRq1Bf71rJUJQrsQkFwlI5
6G2IOTGfa7JU5QxOuadABxC8csTEmrVU1WmUcwU6y5iPjTxZKR0IK5viay4poCyn
nubpHAf/bxBKcpTZJADEu9uQ320h8m6uWYiZOOC4ZKOf/1IPi1jy2j4+SnKh5iil
ZS+bPpZ8jWoYp2URk53OpdYwK5qVuRNu4u0Cp4umgsFOqgsJzF5XZqefp/6q1y2Y
AA0DNQR6oQUfJFtlDe1EcTbTvKQM9RuF0W7pRdO/ds4en9YnidaGFbtQS4zZ/+qV
oXBk8uU6TpGdKJvqhHYZ4Orcthzkw1ihGsjknOkM+jxNuJ1xgVP3maYU4pZtLSr8
b1CrFzwfYzdhlt5Xu2+N24SQQ8rO9jPi417ny/24oBT/kFlvxVqT7AwzjvVuemNP
NraAfXql4g+rDrB/ZznpBxp5fafX2MkJ8mOQjQS5tf9zzTjyGPI2TQ/R4ORHqHGk
Nb3KdbpWjTCRnMsOUJzF0h1in3s3SP2qVILel1FtWbC0dQfqPsaV7C3qcD/YUhF1
SMz1Jc+ZS6hXDfCNC1LGwlEp/lWzaqvTP1tU3BAtXYK5Gg8NlxecJ5JydMvvCkLS
yNZ6qC//DDe3yLQIRDxhE5llAP4vmhK+a3b1C1Mw+634WGQS1A8vTeKFTHb1uSv7
sNOTWCycsby21Gr0r6Rk4INIM1s3+oUMEARGTOtVlJ8EZg5o1NGR9WxeVnZJwQVj
O6F0Pi0bx1q/VhFxN7LyROCwYCDmCzdvZpC1uxOw4dZw6pzCMp/70tja/HofgXIL
A6yw/VNYJJeM5FgES6wog8pz1BkWoksDI0JhaQ8u81w=
`protect END_PROTECTED
