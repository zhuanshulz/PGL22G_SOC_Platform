`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sWHjU/2uv+2oTTA2op5F9pu1u7+XN6QJsoy3dsvvph1AgHXLUhQVw0sIMWT5Gb3N
nbTHUhIqBJjjpkflKfkWzuXZZ3ZUaNd3WEIFJKf6Te5D2EinUNJ8J9Y8lk4XNjN8
b2G1N94lKITmkhqy5cCDx6jlRgQpJaDhERNeCCrsJJNYIPt/7wFDI/tuLadZmT3V
St9xfHwi2NAnhmPqrOjXz35RKJ42rEe8/VnRrlf7Ea8nTVMGEAWLkKhps82dt5mn
x7m9tLCbIeGY22BrqEcOIB8f9EjvInWFY32CZhyPl9wwdUt2O6JVAK6DKeOzBzhl
7Shx6DuAaGA2kTVARc+3/zPYVugj3nSLfqFGiLroQse/3/YLry/VdUOm4TZU//GP
JuYT/TzeY7C3QvufqVetr17XNx34r536pHAM89nPp+NgA4I07yJz1Gtd6WT7gg6P
Niyo96vNsJ/lRmYAgmwoLp4qTMyIG/PkfCiVsLHhW/Ras05WmXl6qn7bX0m2ALOv
q8bi2bElqv4D3dmOLp5zjz0QgvbDib5UCb3VWGPBjxh/Iqe+kxWexNZ/kAFIGCsa
98g99nqc5mwaCwaWg3Rb5uRouo6fLQeWjcuD+6lkBZWNq5ot50TI7QpOxr8v7WFa
WfwmCzVdToCKFW4cPEu16Q==
`protect END_PROTECTED
