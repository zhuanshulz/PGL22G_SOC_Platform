`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w03MG+OWIpxI5hn0/V/09lHk/Z+axJhrywjREJBkIjTOc8ctychK+u95vex4t+AJ
OBZz21frAibF194/u7IVRd20kVYl7Wnhk9iLL7SemCTSfWxU8X428/iQydzCtx5R
dLE+CE2e2/UrJaGuLBt/Lgj4xsiafcXSnuJnpQt1QXdk3eOsiHRUo22wkm4KO/Tp
DK98vbg3wm/aDyBtM78vwCn4ucWRD3Swyk60PHxZpYx/yKWYdiWKxuqORMdVLBzg
kbmiGhxvnP/OZO0g+80/z2puxOlQPjRyFnBn9009qhxZqEDG33VSWbUj7stlipcN
1Idj/Vpg/xintxJ4p6iITbunKxqni/uDR62VHi+ywUTX4wyJCCLJ7Vu4O54AvxQt
FuNBHMptE9R290j3NAMmG3UXzNYeau7kUKMeWVbylhFyFM8N6En4+/1L6dk83jx3
zh3Th6gnt2gdU9RIYcct7393tYHkW/Kn8pD9vzUjcyrt1ijQAY2vB2E91YLMg5k6
9twPnYUnCQ4DlQRB2bNTQzkT+0pW8bmvXR3C5S85TkOYoZgjTQtvtcMBQMAmEq7g
yJbJYH1HvtAa9XyYCAQeey9G2JqYUpnh/J84zA1LefXQcEnRpsQrLlI5pAFNlRSB
lsyNJNQFIZ5iMyTmVy2QGQuujj4U5EpYp+DD95IgKhiFRoBNeh5g5OwcfYniClfF
6g3ms1S1wHzngZyWU0zsyI488CUkZmIHziGvDJcyK1JQJ62QpUSeRQatF7zn1yOK
+wxUZAdg1mjoeiCZD0OBbeITjIxB4njKONdZsTW6SSlYYrONNwBS7W/xLKd3DFj1
xAmW6WOKYtDZS1p0c25TUblydfhxUnvVOCgSBhrnG22njyeXl3ydqVEm8i2KVnyu
TPeviWZgpQfG7bpEPRchyNsnrVc5kLTS96VzIH4x8y0Hdd1At5C4XCbqOmaYdGHB
4LCX7DsGQTOny1Ym9Y9PW+q/CrBGbfJTPAeCLV3UlQK4RgagU8qzMV3voBv4nvxC
jILZ/7zPIkJi2wEh1pg/NRqPX+oIZe+okDCK0rVCD7GCGS9v5zEfeJOzcMWWx4E+
b3hLRkuQ4RxFe6bd2OpPRnW0dNRe7OS3Om30L9ZkVqAGmy26OHepkFKgjHy2tGhf
/AhHCvpAp8gA3PaCy26vkd89plsrWA9D7ruj/iiva8PdEJMl9vYC9a97t4Ys1bWi
pzMc2fIgw0X0DVp+FRMf94p9Z/5uD23qqvD65Pf5cxn00LSyjzI3yZ1XhOPlLtNT
Zdm2o6fNWOopl255o8UOgJ0pHaU1PcCC1m1eJLShhgjk6G6dyDSnfWI/s3Kl897H
RqLlA93pqUVoLrSoSCpuZCLiagl8nmiRgq2byj6Ye/zK+AqUw4jkFPIXKkuubsnD
NuqiCQ2PyoqoTWxHlq/yWH3uBQ+cYJY+tGsSBKHYD8mn9kdFvSgs9gOdGY6KbObY
siTkVWa5DOD7jBk5TgmkrK3L1mdmRRSNPqlAZpqSwYQxbNqFOCuP9YRV3mIUo7m8
6kkijm9PAQpf9XBKKvszdDJmooxghz7d/hWdHm5Tl3mJuYVQydkzg+chRYEsJG9R
RiJ1Lpq+vO9Bxks1rk2yiPAmiPoz1OLQBT6Oh4LzKw1Ez1EgF/IivZ+PF7d/nBQ4
I3Ik2/u4R3RwgPvrukzg4xh9ZjpQiZXIBIm6BTuYAQf5sbaIwQriHYfGIGzH5y6R
ayr3C95xkctKr2G1qChi5IOxu7Y5hnM3oK/HtLoZ/yOS7osmlMawnvp3Q3HU7X1j
AjrXM3qwmijex3IQ64fY5OjDgBqNqDMdvKUTRaL0Ng5D45rtDP4ALkhfKC2sHDNZ
OLbsshzvY54mxv9kXqwwCuin+pirpwYFyTcXGpPwRAI8Ae9V9KThAFKagPCa/8Ou
Rs8ZMeVmv3hQn1rEvkCg3I6ujqcMcC/GSB8zzEDzTflChmm6AhaxG553BSOc057H
xZF9524cHXz2cDYcZr+rukz9rqbQYDc2mCxt2vMN5KMM5gmmlWEJtJVEtoUR049W
R0VZi/CRLEDncGNnxig87RQV7P4M/qgvqpl5/IGhA13MauoLhA5ByiPxbys5nfLc
ZVsrB8SgJUpYkCZ8NgcqZp/u5cFUHMPaxLkly2dtb76ubn4e8rgJWLZMCXon7KHh
GqvxLRPY+zsotwmuI9SiIsBbhATIOcM9LdqH41Rvj690GYY4KtznVL9d+OvguzLb
MTzP80Y8vwQMbl68pi5+nHkSiDXpkf+8QgX5xVqDLJlbxLXHqDMSSPK42/D2Bhm+
GKZ7BGPaq44s7ht++oA3ZgblGQ4b8Qpl7tFXbztWGVxBnCxT4xA7YLMQPDFZjNN9
qfCfNBtn7IrtGEiEV5g+v7EegIG+K5xx7XT/viA3aZy8vIT4KHFyTC9S640gB8Db
2w3b+T1ibeP8gnri1W3dt2NY3x7pIlxq8A9kBkawnrE8XdzieGZlfJ5ihI+ETGyz
iCHMjX/tKFxTcosAlCRwOGvfsN+Pp0cV+S1O1sTyet+mu4KIKQ3GpMvwwncMDD8f
hJ8vCfGsgtPOsJuxt45raNmaS1oTaStqRvmYr4y7w5oB7hWA4EO7EApQo7RSJWjL
sOZUbLWFoMb9TN7xTp9NF/nDLMmun8+QUGVY+Wm61+Vj/h9XDiUrj24/jDDJ+pV5
863bS8YojdWuFnYIJCRreol5rVhGiesMAjMUbLCOshp46rRHZ3Xlet3sudoYRiBT
ahznaO2CVcbAqouU/ctSkkc2ftfIYGsoQ7hSzrOvZdoJJm7ooPaY6T0gtur7z4gb
DMzWKemXvsRtrCN884q10l0uigFylZqrPy53z5gDVPhks4CjihyGCZRwEQhoQb2V
xXDYNtSOs1lOo0cBjlxcaQHG2mFTTgRtu52Ob6h+ivV0JbvErWuZ5hhw+8+LRLZj
E2jet4BxhtCPhC9/Z+SQXVC8jwbpARq1Q3YHnZgrFv6sbpp70olYNBtgY5fn49BM
AjOmhKmJT+vW5txYgVZtK3/okUrgHroHE0KQfu07gtXjrgVb9i8xQ0wQkLyIlH7e
cDNWBUdkE7ILwa9JWWOBqr8ZLoFrAyB3yhqpziFZ7qsda5sJ2BPMb3IsEktqrGGH
XFid8sQFtIfCzVJa7l1VivtJ61hASusR35W5lDnAz8L2NLFcXMtsLOMU9FokCQIb
yIziCafbKoScmOegXSK3qKoeUDnybRcOQPXTPkMgS7LvjqAJ3OSEFfb81RoLB/cb
5obgz8epAKQIMIs+47TDZ6gVRiaygrTctj+X48D6cr9Kh4EyfwpyXPLiAdJDd4cp
CZbBl6GpTdGe/Ywe/1Xgq+/fkBVOJPDzXJ3V/+XGPm1eDcsGHblMRXfQvW8FhCyz
kHcGUnBVCYayiEzx6Nulnv7LQXMbnLkS3B+27MG28zoJVHcINJ1RT6h6wqCdetlq
9ExisLLknt+q2u13e+y5kanAKUCW/yROTSJKJrWmxvEVeIdyKF2W3pgano5QInhP
KNhMhbdGF58sfLCrujwHh14zXvNhIVpCsoO2WqK0FHY=
`protect END_PROTECTED
