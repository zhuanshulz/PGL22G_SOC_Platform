`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rf6btJzwLQDdN3o8awLQW7y0/dNvzzlcMXXmHeO2y7GSyXMFNWks6/qgqV6hMMRN
jddhAOmqLThdcKd4BQciDsYecedmBaH9wxmX03R4WNRlgAwEGc6DQgPiF079cEsk
vxcmsC8Vv1BCt/TXE5ohfCEfLRKpVwU5JELDCKlYlDNm6kg3DQOlwoJ/x2znazfw
cFvQWYDXUGUcBxsUMFuKCrdxcPIqA7R6AJOjQXXQaXtGU2LpPJFSQ3VBew8oA5JK
87dYlP5b5+rWY/rmJRp1z/1nTZDF8Nku4zUxUH+ZK4/ZTQNyHExA5CLexBaGZw2w
sOPFkeaAIxbYIUU7l+ZsQ/HrK8RNJ0BTIfpNubWB4gtDuM1GHziFBckDq+T4PzwH
8/l9Rd233MiFv37UwhPzTtDGZpOxYZXCa8x5nO4Bvutb1MDq8tkgWC0bNMyec2JL
4iWznRfPInHQGAWxded8Pb8reJU5CkiLZv0MdesKYwaAQtQTYnV6gpxjYR+QFHnL
LH6mijfrSAG9SSC4zJP0ekn/56sDuNkao+zrzvbxnldfIcco1LkVX1AS09xJokEJ
PaX6AqMn2p5x4U4Zn0TC5fZ+7SppeKIDO9Xkn2VRgSiV7kgL36Mv6/OfRJLrKVYn
fC0jh2tdwOOeIli4tb2QHjoimbRLyz1gCxuSTejV7ZzjNe3yrIhzQuhajuWkq1Rd
grc+YfTXpMeEIr6mSApFjJ2rFY4O7V8ovI/UpAgsUKdrqIjG7G5yMmHjYlMAe6z/
wzV3rbMpR5Dw6yzlYF1ehVfcFbtpEI+6sNeZjMqjZzKgA+GI3AnC80XJ3LZqspht
+VsdgAmXyHJrm0Po5ISXh0O/yJWdYy3Xq3FaUWnH12V6mppEAFku9wjre1tJaGil
I/jOIWbTR1kEr+fFTzLEOYPrqs/r2eRs91f+zuP+L3Xh7ZKjRhek+C9Q/99lsRMF
GMXOqSDm1xzQp8Xx3wqiGeoYeBDZc8rKauoR9ZBKkqvqVJIoIoIf+fp83huEHet2
1FklTA9531K4FECYPyLq8kWALw2I7L9qP9TROxQdti80o2Y1ehNd+S0VddvNtr39
Hn4tT7jbU32OpVhqvs+UqS8lClmnBUKCachgl77DzjzQ51vHxm7pc8aMvoBUrgAW
0BOOjfgUmwBluYu6G6gnb2ydxJNuOhIMcP+h1KusyE9AWpA3IgpjEs0Q1Yp+SQUH
IMxak5p0/GUCelT5rjE6Ni2irixd4H3HzzX/2b06lsCserscobXPltIVGsUAPXjF
TyixzAN9hB/bz6h4IVfV0nJbXKaIhgCvKwSn2HVzK+8PgO/QLCh6LDHc2gdoBDLr
SaqHw0ipizSx6ZsYT9EDIZdj6GR/RXASYXrc2XJ0D7mk0+wE5Qd7Dd5vzmgiP3ap
VhEgHDuMcaPxMFoRiSNQvnZH6kanvhINTpYd39W6FzS/krEPkg2afLBaHKfW75jk
rCIZcRGci2q6DYz3uSQ3xkDo8cjT9fKHG250ZhcDNHO8QtCRN3CpdGxOf0sNbjSW
A86viZI0BRcMIducUkazUi5AU1XJno1JdvFwxCRafXvIg6b2lgT5jLyZCJpRshNM
L1EzBswGyI23OphLD8IdbSXKjRET+nDN5KFMpPj7zfng0CszqlzZHsarivK+Dc/j
LFa4aRVu40tiECaI2AksRNw3gsARmhw+xwfv9d4LMKhT03oqzUBgtejIej5oTxdi
JCbcljNoQssLXRYJQHdcuJmBhmmYIsvY8lkSuYmYfVVPQG+ZQGkPrvCOdz+4nLC0
eM8E3Yw+ADb7tTEU1Fnk2vINUQT8Hy5rt1zjB9QU1XnV2VkJRXCxH1b3t+2ml8ej
MjHVYiFI50zYjtnmPjJPSjZfWXy6ASEckdVQOJeZRB00ZbmfIRtG1h//CZnmHjTT
cwaRK2G2b5UfKDXjZS5FjFyDLC7GbvmLyzL0fbTs8iNYd41pED0iYbv+zgKFC/8v
fT2UfJJPzTepwoGdlxUa4Lw8/g6UV1ghGMZqIl3DUtfqgg38K1tJ6odMBsaXjG71
pZtnabHnoO7wstYPqqDqJwEAA3RmdwYRiLQzNGNEeqFOgpQ22mlv5e+jK1NoqTVa
FSyy1pDItu4GuMKUFMzjwBdEG97Tbs3bwjzE5kyDbsswtb4GqYkIJo8tQDec623L
5wJAOGqw9mzkg8K2LYvwlsVtuUze/lIT58KwqvVKROP8bYBo+4Lx85Rr2Na30N5Z
B32CgEApRESCuMjzjmJvUpLiNpOzemnCMXONHkAO3CyDh+hOd/wPvQRWzxnTZa6F
gJeK2mjFvbp3vW6mmt5FxrCaKXqJmX3fC2WHOHYliyqjc+k74G2b+Ae3IpKLK1Hc
IZG4L11G9gtV2YXn7rJ8updevDwK7jAb4in4MC8qBuGqFoseJ4rXKaH3H9XH9VNI
dwaIrWkMvAuiZUt26SNGxFSYHAhzujmaOl7cMO/YzV9KfKqP83se/bmgdOnkj3Nt
iREW8XwsQlafBmBiD0NYWXGlnl189ehH4sT4xIbfA7Q2umKVLCrXaS3/bTFIwl14
e1xYowYotICM7AuXI232y8JDGBCdNyNIp7oqVZ2KGzXM3A+VgCNysOHZoKCwujxi
XFekJqbUfDMYqHfQF30tCqOrdlG6gxWfu7yt0g3nraoyf8gvdWOFGYwro6YfXMRZ
IAF1LDEvGc/fXsU24zAbfwtRHlJCEHMyMS/yI3H2QMet93pIJEm5P974hy/4ugcD
Z7+LNN8EQRXdTkdMAgS07jquVeD55nY8uS7tJ/FUQZ0=
`protect END_PROTECTED
