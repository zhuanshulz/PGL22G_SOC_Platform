`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OCfjnvJIkqKDqOwda43BRJmDNSaMPck5gh1LOb67V/jnmKCWsd3FNK5pl7YghkPo
OIKk69IdZ8pakLn1lBshQYPwjuyeqqB6ZZSNty6jezHAL046hiD66RUx1YkniIM3
4XKMJ6IHrNgGpAEPS186msbORQ48M8qypl/pXgjhRpDvnLRYmznwSfYMC5ggZMu6
/Yt3FMvMANvumoQo1GGjD2G75OU2ORH1OaXAIIvk6CoBdSbX83OAvzlgJL8FOH3G
CSop36iYHJOuly1WkP+fnT6KDfvWy2d6DiyZpUXZK3q9YZaGauQrtcj8H4MXgkm7
ttnRIsRUEsdB06+HKQTtWk7FyHVbPZ2UCtnHyyUAPbl9gogEJS17eNvd+2kLfC1x
fM5LNDcQ5ZgZCp5pLtBOb9rOroCpJro3+wImmJHoaXQnfcNiaEw3Xe9NTMcF2J24
wGt/nTnBzOP0fRSBoCJM8/o5CFbsSe0ygrLzkVlPQZCu9I1gpYSqY+s80vcCqYEr
0/Ivzsuv3ISf7i0ItmrRHMN0oDy3DcckOeV5h9bvww/cx1WxGahsPr1AO3hfci0W
tgRLOpW5G7D1RpRrjdRYkdReR0X4NfA3Hp+uNKmbDdkSgbgnoDVbOi7wsozZEHwi
t+vey6Ujo5Zt/JCFSPPQLw==
`protect END_PROTECTED
