`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O4aNl05ixFBIAFfPK3Bz3AvCV19XlEAbuNtCNysU2YTrkHNaTidwnPLhZDVDhiyP
iiKpAoDOrRYXOkvz+XGXH/Giwh01IDf0lpmBbDOvx6CzRVqw4joFwhqiK71z1zmb
LyvvCT9ay/KHtsFoqy9VmCzcMP7qeZUJ38MNxNsbHiEPmRE9a5vYGfb37Vtm7HFT
IlRUHaN/jHul9KB93dgwTClHXsK8PmFvzJm//qkWtqpeA5tFx5n3R4MokHwInN4l
4Lad+w3WJjHIga8+DC5R+zHLOoGgAV+s766dM3Br56Kins09lF4uB9t42UTDYpY0
YDMP5mrZ4zEpz74FIY7k+sLIn+aNi9a617llzQuUGM6wSJ9gLQKoCZwO7B/LhoNW
EOorZVDV6E+zrMg7MQ8QaugXJUL4Uh8RHc3b9wg1x5SzrVmETcwYsP/N3dfRljxc
f+e1EgIdL2bXz1OgbahcAGsp6g5KjJotuGSa6Tr4LPw8X0i7s6p76O4SOJYqPMUj
ZgvZWpkqj4r+6o4rt0jzrqboXnbwMsX8GW7Tz+Y2Z8z+WLtsyk+1cUU9Gxir3XUp
FPBFmI3Yk8YFFS8r0JvaqxSvRm1GCVBNPYDIpbyVPPleuoJSCbvtS5B8/yrnNfAa
Hq+5Vti2VOzpOdFrnGLoKasoTPILHn0L+0iKbIWiH22iQpmUeuucJBmb6PObjgQe
`protect END_PROTECTED
