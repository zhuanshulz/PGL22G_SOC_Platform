`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hvmNQNQ9rM1zLD/TGAaHArE3ZW8zup1uGUCnYsbmR8ZIEkGIf0zSnYfRkVAKA9Ls
OoDaZq7gtI0sU4O0t8Uc5ko2poM8B8d6t7/uUQfLYEOUVPOBKjCKgMQMJ/f6K8a6
YwCrib58FNLGNK70skSk/GDEPEamdxketnT2rov7mhi+B3txEaV0pnK0Pe0bujas
GafJCYJc2chaxDVFBRZYXTVmOJnGBI/2qsQFfkGVMJqh5ewKep3vM534HcaELb2n
Re5puwKYi8yF5poaTLwi9OWOenHx+yetGiJkVWjbUKXCKCWk0SManutrITatK8t1
Abr8TdcKap3T1ue5dDsXYgCioT1dO20zEq7l6LObxTeNknhDmGzwCaagpnqUEdkx
lwWzQzDreYhrBIBeSyyz6RlcJQe7Tp0uttmR3lliImnbtqpsreOvfh3vbuu7Qiux
y0YpiwoRcBHRogD5hcT6bCBCy+NksgW8dG/sgsgxEwXNs21KfqGNmm7cV5IG4rTX
zAsS2/DVzohY6LFZxNl20zJxSQfb1mXQheM1SzHDJY3br/uAWaKQib0BNX06s58Y
n5tb+7aRBY2Yw3zcNINd15XK0qM+hUJKkiy9jkjUEz7/n07y9j8w5JTcHL7ZsqxS
`protect END_PROTECTED
