`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zTjU5Q3zBNG39t6c7bUpXFcGPdOIKmv4yfnOqMOjsn3mYTtL2WYAbzWxDnIop+Yx
Rk5pQr4Tm6iHq0JvUciXWbrdMuzLl9llTxQAWHqJadqqYImLOzoRY2n2MnnFTaGC
MUIP70ZhHynMCv/LfaSbd+4b0M0ZR+YeApyqzajggh1T+BBELK1yxmUCp8I2CSVC
GtJq3QoX3oJAfBlmWmPmtfTx3ZD05iLNcMJDatID9JHOOpHU/N9vB+9pC2NHN3e/
A0FKGDP8qt6ZfutnBHYg634SlFov6A13idPSVT3LtkveDq5nzyaiuavcNyNadEYg
TwzcJWSQmpJ/JFir8s3BGLBgU7Mg/MuqLAix/PYQXFoYk/aTiu9FQBbcLUzlEQG8
wwk+z3Lmjm2cvekKyPV8Nc7bitR0LSFlU3uq1qI6xTFhdWxMbUJJi/iFRSUeeYX6
EXNy4RCJTI+f7W2QTnXmjd+oYeXLQHEb7+0tq0/HeXOpSLoJ/TebvbQmWXxulR/0
GXAIOEjqdiviy16X1g3WBQ==
`protect END_PROTECTED
