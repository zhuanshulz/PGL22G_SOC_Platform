`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KAq/FXrogbFUq+tMMfsf55O/AJBcx/n2ReDAYbt8TRlSrI9Uhg5tnAQt9ayfusYx
zTPv/Ef+yldsRloY3FhfuC8YbOirYAcuQrBsN3E4YUN5zsQ9u4HdESd31vzCGj6l
Kagpr0N9sV5aw/O/pkIK+iTjD/rlZjDFyDL58lumEnz8VgC6xwGhS924crmUJjnI
7fzAwIZ5EugVprE1LP5G0DLBGKWFJNDSiiIXOkpFmFRARjToAPiJwyqT+1DgP1sG
AhtGgGFSUEiE3lD/8vNQKJ4iIqVdOQHqDICDT5e06Upcoi4c2r8f5kY8IP6S6BmV
EmtOwk+pSsCBE8RCiqJZH0faGAzDpXjClprwjeGKlozBWE46ScBaM1j/lDvpBFwc
bjYqH2dqY2WMOKVDwsZ7DFLBgPUZNCHyfTZNxmqmCZmUEsupDnb08feyEhUW8oOl
1x+JDMBgCMkTwjFE0o/g7qwh9YiZWrnTp2qXm1R0UGbmaVo0a/cFwpAqwWAVUXNx
UYEgbpWZ4kH3PjwPpEEA2ehZr9hPvmdoWrzwJc4UbmuegMn+mAx5Ch2/HxO9Xlgs
WnwTNwxjoIh4bh6KBPAnFxfPW7w20vgYz1oRaaukd4BEp/aEL8VxEa3QBMu+xRTu
ljVPHu7EEEjRJAVAIUIwrs1pWF/IRQ2Orh4tJ6oZmT3bwGFf/GCXxGMr9ZxID5vz
C14d2UeAwFOwZfsx5+VAkw741Lh67M9feg6FamINBY0G2xA5l+Gj+5ns4p6+alHR
OclIGLoTQOiJw7o07m3ovA695hLqcRNqhBo933Ah4rZbHODgIqo1aH5hzsoda9nn
bzZQjJ7jNB/stLZ32X07VIllFGln7OaYzSEgveW68AI=
`protect END_PROTECTED
