`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cM+FWQl26n2ZSAfC6QZPuLglgnbXlA57SI+8RBqiECKzdmzfOJsz1XenP+Mg9Uk1
y6n5tHymf39ljwJeJl3sHuvnl3QIiie1GGp88DZ3B+G2vPZ3Bfv4NJWguC0DV9wE
9xZNTRf8xGLbfz4nQB38+5sgEEPKIszzlyGlLd+J776bgmTfmpMvpwwRPPP6a769
UvLZn+4y74kP+TOo9XgyB91TaDKPGCSydom48yg+U0QoJElEQq/okrGuV4dTirtW
xOQpqFcpfpapTwdoJvLN1vJ3UytEisdzdOSlCkefZ9bf7EzeZdmG9OYKcHuZ4kdB
kC44wKY1C9KRDoZklGfEOt4XWyvSJmWaCjNBq81t5cIJ4nTtpzNzuMMCkrpMS/Ud
uJPU7jBwtURiPRStKomGbXyakdR3m7YKPsthzRzLdX8Qqjc8lDsaQm2Y57d1Hxfl
2hlVHB4PuObnBUFmvsWOGe1MCKwPm67HhMopPAtB5+z5kkZfV8YIzBSVGhRNsCME
NzMUhaXTx7y15KHGF8xpamYoZnFkSO/VN8MdXsZI3MvW4IKqlm+hdTcrrhEIZ+mB
MJSZuF4ep++h90VynSLMQBqixtu2pvXWkqJiprWpu9bRyOHXbrL2hittrG1zWE0s
rDK8VyZoqdpWp6zYX078NyGbX5LXFmeZtkUwxvB49v14T5FrcAhYvMMsvhSxwM1S
lpuSbOCXqLqWJFw85mZQN50QIkpFqSkrYagBKT3fmt2jr1lMJuOoac1wi3iHC04x
yOnMXiiVrQT9u5dx42X3b8lOfWMvwhNPp+4n4HBIFSsNJTgkU3s4X9cbHEmFrmeu
QS4zNl3mm0IScNIK0tDVirC3xxFbWYs4oLA8+7fjA4o=
`protect END_PROTECTED
