`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EZtOgx/kVgnJ7yRXUv6ARKP/PSbxrRCy35CsyMlOGACnH5pL2g+PqS23Y5XUBRM8
96FtKlZMN3nMyGhn+KpqTIH74v3FvzNXTw604RqYmwpqwcGVthhEikdeDhfiI93N
YjE6E5HrW2ze2cVzZkuOI0RYgOED99HwJRhJfnwZVap41Sl+rlL/HhCsBYfDbcyi
h1XqH5gCaXJWsRW6bx0eIShp7TuMg4g/i1BB/0mdGyMhmHvxkEXZL26aImFWz6a+
gJ02diQXUnE3ddn+YPwz8gTEUyFiu3SG2eKTMYyFW4hOLYXnqift1JYT0rz+mlLn
nOtk5EaTzZInL4MJCwV4PQS+/c0/HngK5rMxxunVJAx7MnrwEiEEBsXgDGR2zR0v
7+l3efzJ9Y+2N0hCi74LVBp9iE76dcK/IK8Zl5IJTIKZopiRjHsykSMaRyPkLd63
xVaD5sn/BpNbqSQOZwekUwIeuWdTJchtpuHwJ/SH0lXuMEHSAzWAEThfG+F+Dlcc
zjNANYxS0CQAYS4+IauN9qmUgY8jyrzpqlJFNPqf6tQyO2e9TX3VPSaOS2N2GlD2
JBU2sOXkBKmwHm3gNQwRA8Y0ymA+VJNiubiF+dk9LCemDloLrlhHNb1coV3SSBSY
7/ZhydtdVRAXXUcbeS7q6ItTpn6KXFV23g7ASU+Jp/T9hbRuIsIGNS6PLlE3omDL
q/VxYWDFtg19cMo1wBYkjtSh2xu5ddR09EwXSAyn8KuVMUcZaVctBCeKvxvALGr+
cWtQgpNX19eyb6xyLxDLs9Z/aLXY/Mzl+Pbet6ybIm/5sEwVtXryBuJin5gefD14
Tw4wixXJMmzwk89Lm9pMp7yS5AKfJigJYr7P4K3tbzBy9W1CuGoy/Tar7L3+rfmV
+3P020+4PnrLvdI9M/U+IfKwHBSO4PBCXo09EUSaBT03ZzFlU+e5cGGYUIHaTEwf
A9XVFvnjnw80iY8wpmkVzNA5IvjJqhmcGP80ihW5uAA9R81LChljCi6q7NFHVwTB
yemxHFObgP2e3Z6V4S7kmTGAuuOBtPwhLoEYR0u0rnAjBgFE9dmG+vkOPgQcKlQf
jZCQ08Rq6xs49X4TlvMyD3s/Tsu+fboVZZOT8Wbyym2S8654v6w84gsYctSVb6W4
1vjujtKiGetn/hbcxePN77gmZN+QnQgmDneO/RsJvZ0XQVmbk55GmkwO60RJGi6C
Due4YMvTqFSq1ll4QsQFriWsv0lC13eGoS5L+666reKeM5s/y5NpDoNsrQn8pt4M
LygE7ROA17L2YYA3mz2cFi5+gwNEXwT7W1yueluFrG38weFWpLS6Fyv51so7Wyr9
cSao2B5rTQZAZE0Xy6X+pzz+WRC84tJ+GmlOTBFZrWsUiktVQlWEC5JFaqeG5QaZ
ttax0iAyGIOspA/6DyawuVPaB9wHKkSeaIfsdR9tGgFNXpklNuqNtiAIzxtOrbCA
RBiNowZ1AexGmcBJPLNNIPhDj9SwdeDbmQlluNSpWjMK15/XXkdvsKGAOxev2RfV
XWCUP9UmzZeMBc9Ewb0lHgDLxoaXiISCN0gPRZA0H6aUskMcCdnGmDEmlBo7p12/
/w66zwSrmc7WRYCamMLOqd4dDBOCXwHF5qa74Ay9PGmC4+vHjjWQWdJAL6mOdRf0
CPOfTWs5TPT4WB9xGD/nBpK+OHTQDHTAOdvo8/t1iJ5bJbqTIo5UOu7xhXLkciLL
FqxgS1L10DrwHJKnP23yFwP0ztJ2c5P5Bg4BFxnbuV4YocSIvfJJg6H32b/DWP5e
Ltrw+qhAeH2hO1Uv9vT0FJwenpAGCHNa5GVnrBtX23P/f3bMLpuJtg8Yy0ATCr1A
pQxClrHSP1jx6kPyjs3NXg==
`protect END_PROTECTED
