`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nVJhmuYFF1Vw6Yo24scxDW1BQOqNVV/jh1FeN/lIuQ1ZdYjdfRqToU+uqZce5u/i
nl07cCvGYkSDUrGam2lNGozdY8zY6C6kwRhVIl6hVdR9ILFlnhhMbt80CJs5F6Lk
JnQbBPYEugiiQah6ZegYF9Rse76E5l6NUbSNbt74DQTjk3te6SS9VgvndLPTx9/D
UDA0iB2CtqJEg0HXFprlETgR0n0IZ3XxyYh7IAGa2RXOvc4f6jaRfI3xfT2mRQPu
Ht+K5po4x5wKIhFJO1MZpnfZa4qTljzflsJmGaPlBVo/lA3gEPFVkUXBvMuiB6gT
Kwi9xu4eFnAt8J9626gFrKNhalQIQXaZV5RwskHXuMGibDgM5liHWMVepS/s2YUe
X3xAFQkvjL4wHQWmnQrhyG43NdSVPQ14RTEkDGwkhBW/mcoJ2T8vTC7bIekeV0NK
whO8JPIYW4o3Et7I4+Ynvj+ENQfoKb5ESBtszhebpbEKiw+po8EBNS0xQTFbCY2F
m1EdPkpjMipWOmaW/Cw4itpGH5RRbeqwx6nFooxclEqvAgRU8rmJYLL1l+g3YpSG
OldaXph6pt/57VDGC/T6MKmWx5jJtD5g2B+T/HSecglS4KOcAhgCTrgiUjbggQFe
rCFlH5CdE1GvzmSziizX09VER0QlW7L44YFWZLEfwOdnLxH7Zm5ZSYcmZXiMi4nZ
ptWXdfYM/fKIaWWZWiFM3O4xVSyqvoRksJ0Ra9boosZH94p7AKfsnVHQ0BZDtmxx
WEkdZKIbQLcvjRdsrBFcJOfH6+sfCbaMt+BxejB/6+7iPqKqiCGaERlVPPu5Dy6J
7sagIEoQt43ipL54Gsri5PywQLyG1o33jTy/4/lKArI2Z3TgDU/MtmJL94pD9mCF
8QSWa18+EqSziYP+llvkbh/btz2R7b1VBZo8UtIaFwThCHu4x8YfYZ2Vxsj9wZ7K
x4pDKLeNtJAz0+ulUOjvGYDbQ9MzpR1PZWG3cgwUNOKGTUiflGj/93/4nA7ttk37
gzursj9gTruuoyZaxY8QJz8EwwZpxT0cByPL5zFErVmtwZa+kh8AMky1ievfdp3p
CeBmaFBgkg7YNmKzwA0m2QGY/RMWgTSenwCEu8Zo61iacD2JcRaAiGfMOqUppbMT
0MVhdHEthHiO3vbpjxNl8DHjL4WDMawkF36uo66HoHtdIJgmO4SLwd78jvF49R8o
B7KmMHyHVj2fQi09DjdW/E7JJOIvpv7IpdKRht0/JxWt3qdiW55dJJGJY/e6usvK
lDfkTrsEeC4vn5q16JVyDCVW1g+dX/ILb/oxoiXgkcMZkttS/nVtcdATqAAp59t9
tcaakBHEaHwmXs7MWq8DBs8FI5fvWh09c6Up5nTl33TRNjQYGlRDUyctMvztHXZ1
kxB+JFGWwTfOfYifdc8BUAJZZOdSfaN+4yEKat0pcT5ydpGsf4+YPnvAbwaa4PBi
alC7x7fKgZCVS4o4ITww66SVapEu387S04nRMvt5pER6KPUU1s9iPPniSPyFb7wI
bU2uoKcJ8H1nQPCrvJqZd86ekdvGz0U58sAux/3hOKd1vYScR0R/ZHOeyi0/oEwZ
3FgYHZp9z2SNh90qrnupx0UiiCaIU+saFlHCNxZXBM+0onzCP8YtxIEX67OO4lcI
kkZ9H7RUKCWFbOII8Idj2RW6bBHbDqgL2Uq6zoN171Lf+OEUhMnVR3iU9R8G6OLH
IbTPADKsjJHCbOY7UyzCXt9VjcDiH13JEI+w9ByY7DWYX6tWykavpFirqztUc7Gs
R+p0tJdLNPf0EGQICGhwAPhXuI6B7PTdtCU+p/i/cPcpNRMzJMlCAi24g342+v6V
0ReztLsM2pDKFRXhz+O1qQJJ2jekB4ocSVAhqAh7V3XnxQuiWqWXAZLyzvJ7aiBH
KYSVeHc2nmEfUjpWtwZyCB1fF9P4uGgbSxshM83a+hbUag3FmMrEa0EP27dzSYFv
VtqyUmZRapjHW7IOyx/36o1Bj9M+XD6MERXEuf92FOApSoiDYo46FDgDwctpsYyo
oIjTfWIN4o29KguLHEwB/jdbYhBV8xwdR1EbVd4P3I7E8dMtoRumS7m6D7HFkc8h
+7xgFrwGyJ1vPakhmjFuroOnhm4Ce7O3jJ4MO5Hzk+/ECsxBee93j+d9IqxdQVyJ
`protect END_PROTECTED
