`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
68b8Svwb0eyzgKAdmPrHVZ1y+MiApcBJgUkYRt+Zmo00UgR60LDRSIYLGywook/6
jJ0BvDS0b4cW0PERrPOrPExURf60H3l8uOntFBtxDhAVjfRU6YAPGrzFe9yGbB8+
eUdmiRZ4anrebzGiFoL9beF6DaF689Jdzu0oduAZ8OLgzMWtXrXbxO7AZTy5I9ug
iCSwJx+A3pnRKvafjtQxahKvzkomrywCoq0rwq/fk+V+UgNwJXR9V9FsIiUg3bjN
nMKoI3t+NNhJZYugaxS3C+pnX/BRjbrJlqQ6chlbqriXX3MkgyBR+kJCV8u3TGab
6TpM7Jlrt7l0tTdD2LcVWrbX+3EYFbqgiO8rRtEfPFussto6eg182jmA1z8D1qKf
e2+kIsfNsTNHNDzV4fva9PpJ9RxhoTYyFp13++pYQFb3YFLvU3nIVVDOJ88rTxSS
kjk2JIXPCAJktJq3EOK3lTiOzyUINlE88GEomTL/aPKdUXsh9C4DeC1hMmVfvPNM
X8ryKQhDee87+/8e35AjpNna4u2U5nPzNysr8YjCNBaNBkqzVXe76MJQvBKrrzXi
zVTahsvMBCc2ZA8NWdcQ+EMn98UK32wmnwcQcg8wHL1X05KsviJCmCpdy0v2ZcY0
VZjkrQWsKYwBd/Y5xuIdqXvjfIn6q9m/HpxLtyRyn1NKnD3bY754qbQsUF53diAd
q7HFxw8YnIqPYAHWiF37BpR54sYKVVc+627ceoZu/mrOELPhMM2wO8Acp0BpKX9F
higjmWNKXlHlnLspE/fwiclIg9J4AclyumrA5szE96wuPAordUwx9ZMnCMW3dnS7
ep+fLAkXeToLUY7VGuxx7tHjXXqBHivsUfNKktVjKRpsINRYgRkf+LX03EuGRRjJ
Y1Cjpi9CS1Ie+Kzxslgy6+aUZj1BwTlGmkWtEJeL0k9w4gZX/GkCGuXlV9KsjUmk
LhFFzqJ0uFzCH8HE+Ku1VbV7/dhX0nSxxaeE+WyRYQLFEFdqwEVborDWcWKJwr13
iw1bObh1xYNA0XjdB2+Tav0dhYLTwrMG2i53uf5nsNXij/gJNYUDMW71/mOEAKw+
0q1t50jVEiMwKkurDPDddTH/Yq50TZZ4tA2WnUSpeDlEwEQMKzC13S3iBkxPfKAQ
WHv5Tmhp66EPmRO5rYkW4NtjlTcMSSSWRVVTIBExLVZO43608CMlS507cm1dvMTw
bStgUbGzrTBUR68qp+ch7Yme7xyp67qTXUcp5jWwg4nyAoLUqUUUdTR2cKL6MavB
M3jLhBGH3+yTAdIRdkSDiqYmfsLtNqFKg6S/HCQeWBPtL9vZs/E71TbwWnq4uacY
aLdqorgMYM2fsmBkj7XXJnT025qFZfz7p2MxVOsIieIxYK3uCq1Nutzuh3K+LX4R
j0fIhX7ZcLPukWQDZtaZVwZMqmwWkJx2WoGVkevQU5JycG6KAyYOFmO/98OXzTZB
2YnXxHhOj3cMlgqxSGUm+jJBv3Ze7DJauGb4WdDZ6oBwdFLfwFZYBcQNqAQMZe6v
`protect END_PROTECTED
