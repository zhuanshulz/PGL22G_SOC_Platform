`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m+NOaIeDvQy/pt9HFXqOyDLXewHmVDc4IZtIMspuWWvQNSPPUNxk2ui0PomvdgPW
SwFBTK/ly5CwR9lGvpgRlWQX91Petf6uNNsPk4bsQbVXwGyD760oJAxpYdRqka4E
xHwShZZbA0F+iRf4uAH3eqm2xcUcaf7YoTD87MQUVoEOByraRkVjrMglfzuWkzQS
GaO9Kv+J3Wb6Iex8Vc7fWCm+UiX7mErZED68szgACVlPcJF5pRmGBkKg2xf93h7N
W88A3F7ZaRAumWnzlMZ9sSV8A3W30Df5Ggj/As2F1T+xhuzwEN1Dbm3+M9J2kTYF
i/50ZyGCyClqRTE7lJJ8qf0ngyg97hX0Tu8pu/WwD4DOsIj0CXLVjKGdP5l9Q7kT
hn9hTGGr3lA8rq+ieVUnNbD1X0jAg/3/1IGhMy9UHw7a1htSg50CNoQW7MKh2JiS
xzoYfpKoEWhVMuGVW0fK9g==
`protect END_PROTECTED
