`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6QhbqVN2m9a/c5B+//h4zaJHRpV95OxfGBI1aSsxVdcb8UNCGEZez5jrI+yOtrOv
ryaWGayQJ6j6aGJR6fDAoOD7qNNz50sTCXapT1XXVBgGpO5J2u2r2P41ouEYoGCs
MP6JgiK40tObBpCDKKD1oB9vYLSwXPco4XsJUAI3Kfj/PXoqRfHL+Orjjk495ABW
ifCBGrpkrzRRDKVw2Y6OV8PtuAxY3CIAMbH1UxtVzc4zrOC0p+jMzZrFXB/Hs640
CY7LlTKHCXUtt6aYf4/4Niydks2iXVrRR4lnNR9YHNIs/eHIzDj05GqfS0ZQBNux
4e+HZNi5qisG4NKRAZZuLB+sof91G8UNd2Zm/Q1/dJqZc59y715b6a/2nqL1K1HH
YM8loMxyeMZSa/xszUVP2hkVWHF+aVCUQ3b45QskuyJ2HcKGsQ7Xb3UQobh/ZZ7g
dxojGjals8cKYvAQswsqrwZFvqOvTuRmDO8Cau2koFK+2s5E1w9JmcLg1QMxCTbW
8vuJrNa4jZ3Y+dgrhDmE7XISmGi28IOnoYQuMVeaV87GT/uZRNhKIGPNr6EJ1hoJ
q059UZ1g9usWiNW/GjugLddEjQ/5OZidgqW7GQIonqWERO5XYtOxz9S1GchGAqeZ
jYKwf2GRLYj4aIRqXIMCcPgf5399dyPK4pXIoeydI2bxzEYglxQJgwSoIM43UNrs
IA7n/aNdpLmT1NzAZYpOiv5n18Wyw2AcXpWYWB1dNtDC4wO6qTNpSpzM3kc6/6RA
ALMq/PVmBDCd5l5aAeUdiVeS/d5s7k3LDT/Sn1gs+SNq74s6a2jLINVN2PWA662j
i2X1jBilHLEfsTPA0zLroglFXa+uPezDdpYS84ebnEwoMP72BLPiu1MBX20ItzYv
OM1p1EyTYzENvkg65dOyTTc9D4b66vMgpXJzgPQmJ3IXtPgiK69O5IPvrAQwZkx9
C7Y0XvXUcyOYgKjlcZJucU6kNm4BWl9/+KUg/OMd8pZTd5Sxg31gjBUC+sRJoSJL
ItABlV2toW54ptp/EmwJmhh7WzXDZ/iqipiBee3nfLphFQaXPgdehQdRylIiIS/U
T3a+fgpr46X1HaCbi5yNqw03Gl3F6J4SNe+01jLuUwN/GdNZikdqSdTQA4ALcO1V
LoCSZeLKyqYYSj8tGkr9Lg==
`protect END_PROTECTED
