`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZhJNlXQZMOopvPQrKbqhhzb7A7CP2ZQR4r1+aky2Fp9LHyssbamyT/Nw9GuM7Dff
+YmMs2QfiJthQaCYeMXcO6z87uvYZ9cKOgx9WYTrHr+2a6ttFLCWMIZHKoYoz0kZ
lthHZb3j2lcIDVqCY8uI/xxlAzIqvHGPaoWgIDPd2h6w4BXSVBlYu+D1dLuDM80u
SpV3PEnLessa/gzSaDx3NJk9Af3Qw0LvDYoDdAZRm9GPzgymRyUrHskwvdPdIhJF
8KVTq0hJaCCYXq8ZwKWcBD9myi/q8HvGEHrYJU0HoxuZcm5o+J6gZYMBJLmm4S4+
wC5Rhri3BJoTQxZ0vHdG+p40quAVnYTcj35+NYqpwlm0YUMlIGOsai6Bhf+JEv+7
RrfU7PK99LK1Cn1IPfR3d4dC5hJpxvF8BPOzrVNo3I9qk/aycZUJ1J3lUmr4QWbl
1brHtFIHXtd+bcxNIYsOh+8nnwMcxOX4iXSb1YRJ9s+g+oCFnVrUgVLMMMBA3X9b
0Q/VGW6dNlRPJjcDK9u/Epfm7cUVnysZsKbqBqud7tgUq/SRVAsRwJILrO1ZT2G4
eC8bXkOV3iphdmjioZaPldItqo63q40mfWIKnmIE1TQZn9R3o2N0VG7u9SqWfwOX
8/cY7OkSUmOV3roaZWAM612+Lb8gVo9WOlMViYjxUxse1xTXc6Xw9hguYnCjtMim
igdkOQBgiPeESOkHV8YOLoyaUGEyRdv/VtbhVcSpZsYslVhz09HuE2IT7rJV3IOG
/cKssDYDSBro4aw122W6a6qcs88hBlQttaGr4ISrg5Ykz4lOtw1mz3V1ohbUHPvA
wbKJ6QtsV6xLVt03aFbagL0WWVWcmTgHhDpLYeHBQIG4htEOy6rcGs0AEzkM1Woj
PiyPlhJqEElXUyzX5HX5SjcTAd1INSqZgX/9SK6dbqMII77pmX8FauNcQtDTZxmG
YDutvOCY2yolTL3JaLxOZf/8S5tqLyoya8Pg8Mt1SyZvlECxVVbBbhARZ9vG/OVb
IVo6D6C9Z5SfZw9GGksa0r8pVZW64vtjjF3foXJkoGZ45NvwR7YpcBK0/BYwa1L+
lIK7U+ib5hkEMuMEdIPgTjvyxZfMyl6s41chOn4hFvVxnUa3XKz6G2M+8m4QXpJj
eysU6flGKG9ha3x4kzsDaU3CD9Qi4euN0FhTtpz+o+irhixJqh2Xt9EowqbrFO64
4ki7LL07TAEmu1oYnVvkEG21IMmyFq8Vu9Cn+sAJH+88DX4Nl3tuU6Cy5evrKV/V
Mdn7ZBCTnSfFmpFIhLClVYd5gUYAN6i/H7HNACG+YADMlhbGse7shrWeJiw6EHJq
c5Z6gKmXGHokeTW5kbcWmecd3dVudjudC+jBCgLJtttP2W4dv+MneL7RJmVuwgqD
qujpQSYar6HsZ/m4aSUkujxCth3KFBmL9s5Q4auyWX40irpm/H7Hw0KvB2dvltZ7
wigORPn56nGVGCwJdNjelRcmltsGMk14cK+vi2vivBOGqT79OEjg8MesrKvWfZH+
hT+df2j91osZXju8IGecXrB42ca7g0Wbr6wIIdKw8cJMLYpsOCQElO3C7eLYPm4R
AA85hD95KfirZsRNZnR7WWbILNdEfEUv/Nwxk0fkQ4kHEnmMv8Z0es7/B7fj1NiL
pwbA79brsqWa02YD8TDxgsxo7YHYfGTb5stvbqXXiir2xXXV17UuRXYShvUm833p
FT5hQbAO4RxhiflK35Yk1eDKYW8AHC6haDOr0HRp+mNNLhbuMsbeyZufyICpaw4J
b3I+qiBIvIZfSfqcek/G927v+GYKxopL2kPf4xlELC6mEdUQNAfxxE4psGwmlU63
3t5DUPlsx/axJH/QZu0sO0zMAeIhimfkGNJIhijGWMBN6MnbKOONFKHQgMuNcMYP
xCRmCjsIfYfXY4yMgSy9oZNgnDNzG0SNYIxDPaAx5LeyFT9cEU6bzHsDgP0BAAz2
ypSrRt7idc73NRA5d6dtClTzAhN+sM9oa9/UShrKGX2JAEugriJh3YttRHUuR84v
kbjMvXMdmWPUy8sBZ80q3MB+he5G1+RWf/2TKy5E+YEgoiW4Ii/Cc4r40QAMC7G8
o+wWCE0GmsY5oLKRJarRg6ASg0lvQ3dixue/Y0MPGJDO+9kYwh+Is5+z+hIO4oI9
KLn2TsWQbRUrkxNo6uP8AuHoXUTtwdyhSFlqarOXDAnpPGuBUe+SLDnjs1yUMAl1
hPjfIAq9z084qA9YcJQScwCzu+cXEuRY+XD4Ms9hpzFoKyGI81k8oCdaV+oUhHvH
L1A6vYQheNZa7NSCDR5SpKIIsbxu8LaO9+doY+SDsrvQt65nTn27LxarRGpcA+RJ
btgyOAHHzA08+sFDvRzOkB2l8JjSPwd1zY1cPiEIuP88Do7UZFH8kBVi754us3F1
h9wYIbyvtfwbEe9cPypbJTDVp8bny1Zte7G6GLW+xlfnFZYaTMexmmyzfT/GOxjJ
SMau0Kx780BLItfWMlyfVsLqcnttnNS4UBKYjwrz6Nqn9a0g+1esWgXDOCTxN4ZA
0/7/yEdlBfb9G09FX/jHZcJlucdu+6849ECb49giBC7LhZ3OhEZzzNH9+fsmgq3z
dcJJo9bhOJzizhfPkGl6BK8+uOTp/FUXjqbQBaJ8VPcWpCOAj8w51gD/3GPG3cEW
rJdcy4khB+yHzVGpl4vW8FVsi/9f6VakJIb/CrKNKhyaYMy8/b60TGgIkESQEXXt
KyCRXqsKxH/E+C/dt/I5ONnM8Bnm4wuoPpeN0O1Zn8XKm4WBbRH6+BVm/2o+KpU6
m38Ipa20cFvF/3dp/Hr1LqXMLFxI6JTT0hnThwLFhhuLpiUaUNSksNl0FYQBVXFG
kJcsYwebB0mROReksc/o6xWptT8ztvMFDO8TyL/TD1PnGtZHrsUhHnVuwHSORNpl
QnVI4WiCvF+fVblRJ386d3/tqITdjFBpFF1CS59kWo4Yx1COxGsaftLkHpvthSUP
u72jDzW9MesQ666xTJS+sHUx61wnPMlHIak8RB2LBhaCMMU/DIxK6lHdTLmtHc2R
Tm0Br77Ax+1MlhR6DLJ8mP4G8jnx8Hpvg1MwQ6HsOHbQYVYCwxGv9bxjhUxxMjVn
mY8Kj+HZNrHClARUnVmC42uJQOrof4Bn7BIYKjWzC1++R0CXMlNSE4qbs2Uwf5qB
tA957cHzJcjlsHmrJtJmLziQQiniWNWhP+NMhVHboGj9VGJ+87dudz2r5f9j3rk1
ZhRREKMydOpiomviJvb7Qkc+B097hXcUxIZxdyu92RFX7qp52spSaBOJfF3YySVv
OK1RiJKoDwL4e10iFxU3D20gRyRMgPORn8gfwa/Z10GA1r6cP/ZFXfKmXOuD+3bs
TCIyVlpnP15ZjT7rq/KUu6IrBDk0+G/7sGWtkeNu8VcoksXPM46McRkRkRc9onxm
TlSznOj9v/r9cqLXSKDnK3nlKjT3y8+1A4uuHt8qp8cwHxGpkgRF5aQlNdwQdrut
6Tdw4VXH0nabLIbAKcq5NWZVqW7pcE0WrHIlJvg/QbBtkzDFSHKBBqBEDMigQnUV
gfvVoOO29ouBX5So9aFwz1OIj+HVS/ChY/cQoL3DrE6SDGdA+K8LWmKiOyPrMJm/
DXLMBGBPcV4IYpvTwCH/fnv/Do9QCqTnktBQsvLYJLcHVWelKIGu8kqqmJGjU7eg
KGhV915cmxj02AFa5nBD9xo7+SFA1s7jiDkPQEtONt6z6gjT6PXqHyKtMxhZtX6+
7ocryGjNUgG8q9A/QoidWlZhA4KBOVmDAuk8hWktYjLU773c61KFBuXnER8PfA42
Aw1TEvFxjaCXkw5Xs5cP+VXRTw9ddyM1aWHWPgT1yMtET9lcb15yRK/3BNte/P/J
4CoMotTZTjEatK8sIsuxworWinxW0P6BDT68BwmX3G1AutexjwTUnzrPV/9K7Cez
3W6Ran3c9ZOA+A5dpqwqYGAkpJbBAs/dUsKWDTJA9TAu1Ws1Q+0xIsOzmFvilUHe
CfBV26/AC9cjc6BmYDiVOOO0roYVxGA+rtRais6ebeumFOK+M55m/DRTasQM07yV
dVwnXs6shNiR7wcAj1TDsfeJF6kVQIlsMF2SDrNb2BI61AtO+AYYtU8ABmCB1CNX
Jld2MocqK/ZcRczLwqIo07p/2oN5iv/U9xuK/uFzH0gZUaY8dqvKcUd3Xb2vZ12B
bq9G5v2H00ePH5+SWSYMUNfKoZ2X1uqspaqlEHDfM9ZeHye89OXYiJWRCm0n3iCG
NS60omox4az0rmFLrPoq/40pZ1GhV7019pxWKSN6BRwde2fnNFqQBEgygoR/XEqH
08varif4XAJlyXaGp8EN4vbq61baFSZA6pkgLbCfCnCYZsTvfyIJfv9tZPu76yMc
LWt93nO6B/EkGkqH04SmITDdUnGexC5WQ108gAqIaprlFKrFXKTa6g4TYRTZPAhB
alvcuSb2IoSn4eFagUTdzCF98Z6UW9NmEFjyW5qaMMftY/K8UBxClAhm81paYhBY
Y/HbCmbzE4ZPx0Z5TxWSBFR+BtXJFxhO+iKEFCuLu1DfaJiFnZktBS39rRRWdCnz
SaG6s/p2C2BTKQhxJqs6hnshohzhiSfKh3pYDe6YMEvwhX23dXo7BTMtXLqSEEaF
yZBeJNEnDCSxGds0GxWS/tcMhWzri52D4bc6ce+pVjLFD5A4l+PhVfu2pHdE+r+N
lkLlNnq5hwML0ZV78yjh7hPhoaWkKeyjsXA6TnTX2TZy5rf5JtZRbW4YOU6KnpcX
PEKPFaOvCOotZHAXICmVpJfSDLii7To8El7fuFU9NX0uwBQqljpw9+BCrkPU27Za
V8B0k2+PaC+WTS2d5VDxMLGkaeGC3f/dLql8TzmYnTTVa/To5Mo5ByP+h1vnuRzu
SeqeRoOvFlG8Pm/BnC93L9TIAHIY8yHievKed6uQmvtOa0IA0ZhCGn56/fsHLBkp
Y+bJz+7kgcWeCcQ6187yaICnjTMChl9Zb3bdnsIdxpv2BGkn+3PMv0JXySaIgAj+
DVyRdnf2IMih42e+ASk/wdzkEFfnPM7Pd5sBJ/omWbrzQVdVFonG6Gn7GhYEWs7S
DXOFGGUkBpl2G5tUwSSY6vm9lhT//ORLTyLrK00VcSfUFnvLu//tPAPEwLbQWHUL
yH1/MU+i8sFMluZdqXoc0ieNYb/GydT0ytO6XEbejVJHGwk5BdbK9jzPDpa8BVjP
xktJqZzWdvXcDAlv974llkaHU2arH6DW/uJxDRDxMVIOUzUPriHQbSEH4gTaJSDF
qeM8G4LXzRYbU4xPxxf78UIESvn5cXr6+beFvObyf9q8WP1L2rBKFz3DDLESs4Vr
XTW3ot0yfdlXKwShMiqntGmAHYExvKj+OQqLa5TcL6ZeMlSj0S1fKPXYFluKPXRy
4+lok2FnoGeVWQElrZZYx01sYCyn/qyD3itDbWuCvE5LRNMlumbuHH5hjH6PXEaJ
fE0j06ud5xwFRdrEMXwG4Tahj6G221dX4umKmKG1hZVaTBvWa8J5k4qKoscuIPHg
Fx7442jM9oN/3jgA0CZZgCLT3kHs4iSOtmJHzYYUi/4dtUvk3ZN3LLhAqBFj5sEn
gbwchj9+42uAtI7MxgbqqQXLAZQp++MTSB/Li4O8WTIDjxlmmZBdrHFFwZPNQQmH
jawkcEXcVpBa40GlRplAbf4LS7zO73+54WK0jxYWVc9XNTe0msWh3IIYVAdYVW4W
b9UW+DzFkMTiEQu/Ia4I/UfA5qCl7twt3cdS9kwvfbbwDnFQ8tgIslZcRXP23VH4
DY6QJiDYGQWJ9IFkdLVMyShRyonslOb9gJdHwbQGwYwhafB7ENAGQaKo3p2YE3Vb
Q9a4pMJdh6jgCoLHJbSh1V+6CRBGY/EJTUoFPtpaHr8OD347r/ytDCVEiOkWDzHZ
b2WpUmRc3Xozm5MYwNWaEaxbJUy1C68caMzI/ccikKxd/gwa++SGeuPNFeeaHbMS
jMb2L3uNygU7XvcUGpM2f5uCCcCv67hPIAs1daErW74iuTltAbR01jONAtSd2y7w
yALMDO86zlQi8L62Em+2GMfCfjEYrRag8jWubK+L9KZY4SdK82T8S4d5KZNR18yU
rR8wmzYpC4M9GuNaVvzTpr45fQqnFfMt/df8Omfta7QM3hqdaJj47jGzJubRdyys
`protect END_PROTECTED
