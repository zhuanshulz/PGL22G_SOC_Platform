`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i4Kra+RSQ+WzgBVqjUWrWBU80UoG/Pm66m7Heed2uV0cobuVMHARGCaJALrAHoPN
W4eHCShQAPPZ7wy/64HDvpXom1p+MgZOgads11BGc4Lr1XhVSXs1x9P3MThF2ZYn
jDJzIvvevae9goJpKYdQDg/rOsDq8WsY9821p+PZJbGVehUCjrTQ0PBPgydnondS
y7lnn+c84u34hqBlTWqeryPj8WxmRBLPX3KB21VjL3gc8rPdWMJAgip4IzX9jTSc
584xfCFja0KJs0Fc1bohjA059ND9FUgec1e0m7t9xbnPxW5/pUCoIs+pLCCYXvds
uDlzTGMtJb8/iT0gC8rxXkP5zAeHhy75LjBaP7EcxN/mZG/LrUcS/GmzOoAt5ohg
Lx6ArgQ3UbDPszOncKDM7TRMYOjyl5o5hByePnQgEGhuxHzMKAZ2yiNpNTd3dsDM
fZkQoV7sdmNyS3SrjnH6pUemXenNlju9zipPnajDSLO7oB1e8aGO7XyK5L+fbpWo
feySY+yaEpF1jF34NCH2LJQSmaaiAtz4B36BJMoNyZc8eKShToTa4aHImrm5UUjN
Rq4LlzAc2d7nhvCB0hPg66tNJvUfScmhbLq+t4/c7Px07N07XksJdHEQlIQTFuqG
HXNg88QPt0gY+oXbE1xWc/0S0xT33q0tRgsWpEtB/nhM1QV+Iz2sIa1qSXsK3Ks4
7H/qwzOHlcUd5Be0wVZaVDU5mLWwmJ53TABvSb2RJas2hMTBEIladqhFnFL975o6
t/coztrLuZDkrAOKP2UQczCU0sEZaQYym0tmUImTqksnDJbc9WMZO1Xg85WHt/KN
abM0uD/ata+Nc9R2OKKEsTpdoEZJ/AeyUoDOZ4U47YSaKuE9AX2pPBO8G+wSVGm6
5ZQOWEsFgjWfHkCY6xzB6oNimuIALJ+OtdkVIl32R6ro5XQRo6qo3y9yZD5m2DkX
Uo27GYpikCBIlfkJ4Sg2nxT3oSZMnY2lQ5u9AmYdRugIDXti62zGLfu9/j3/eJ6B
JdYbqpY+bJsDs43xhyvrZQ==
`protect END_PROTECTED
