`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VR76LuAxPTdbdUKHvinu554u+kZHnfS7nAAxsOWKbkvVc8yLlqHdbeijjIHPAya+
QT/Rjb0JMRJ43Qx2ppz8/RYa+dyLP9j9s++Av7Bv36rNn8dQWJNjsXWThWYJ/bJE
4PEdKoBPyfsaU6Fz0uZnZefzMfxHCyvMU6ac7jVM67TizYGEdvSO1na+B1SRgvqG
p4NAqBv4IwiPelFWxCdW6XnZvQXKCDqlxaYvu8f3k234NUoKCNcQ7T01Q8EekIza
thcCym+ycrMsm0zOX8U4BsFltEAAkD4vjnkpl+2FznOPbfD2W8ZuzMeKiFzFkwDK
IOK5iPlSIIDM/hLqjagPKX3ZmtTZ/9BBfptOT8eDyuvm1veEVQM2TLK5/+Fg5QFq
Qj7XS0c78rPn14kMc9Sn/1T4QeJ1IXEB+W8wDKUyQ1NRuI95usKWk+sUILOJWjvH
VTskAcqxB0Y6ezGKLpEc0CyubZmysYREl8fUCGzXVtTa3iWjkcr/ubfW22QsOX94
DgluqJ8y7Ig222T78Mb3eQ8oiQXYp99ST/v3gembOtwsOE04E3Vy/IvYE94IL2eD
ZBUfCJyYKVYjgtYy7/olhhSaM4hW2idYVYYneKFITEZoC8DbeUOfnfVKXVj/6a3U
kJtw0wRVFHQtVG4pI7K45+iQfhRSRYf+McKsgR+TcJqSodQSBlbjIwh7oiZd0FI5
+upMLpeawVMwSAYEEWiahKiwzcZSeLHkBHl9qSpaR3WIGowppGdFLBbFpPIIwCBs
4NyxGoZmLMLXV+XgKxbr+Y9qNMLPBqyDVNYQQDdRnrxBk7+8TcGVaJBOrL8PJam2
NdiXmWVyItBc7FNa+KcGLa1s8cvBJ6Xxd5Ow7MswnJpJSyblsPI+g2lslWAzQwpJ
XsHFoQf5zoaKQrbgPeyDu2sD+CJyh3lOTWRE1b3b1bkav7OincCE6tMmy4/k0EoR
qSv6LYtDBRokZ+lnWNhYi8zdubXGg4ZnEPXyN0qrqR8UrAeO8avS8Fu6LLZlb98m
jqwDPj644el19R6NJy4FNnz9vGNk7nCiFSUfkLAg3+sEJ3xUjiWis+pU/VjPrhqN
vHbO9kl3QXl3ZPFEBSIkWiVlu0gMlSwafUfErIwl9tTAWvzYoWigZFxFB0S1RNzd
d5OH7JlINuZhOHvh7RTjQ1Z7zehUlg4VFvHyUTk7wdP/V8PD/T8Pe7AIvRGN+oWB
2Yg5ax29jrE4gmn9aYdJQPkfP7hUgg75mEhSQBjCEvKeFrh9iDZq1wtJIxYmOb8X
jYKfkseuC0E6bO+4Kth2cwPrF9LBzqg+tkEstKR50iboJO6fBIJ9CuQt8yAkbV/w
8Vv4K/165JMTw+X0YLo9whe+QMvjmAtR7k1CclSMkiPzvyJnPOzD6XZgO6kgHMfq
ao6zq31Q0lHJlUB/mFRrTdo4WG9IFN9TVv3iOp+tJsdpHC74CEGmqMOWxRyK7CW2
oT+I3KuXwRc7ZVbO86Sao9lPVgwhNLqvW9BNLAQ7biFdB5hHrzfxEZmu8waAT/dD
eChEBOsDFlGbP75FSDQcpdeEM6hyVvf9HcL9L6S8r/FFseox5uOOJW9lLMKlqaae
kVXjy+kcby3Rcg7tNjfUb3K7K2rP24WiZLPDR041P5pITYeaVWt6vDPK+YrvZxMX
bfl9IZLZ5EGF20gu7FvGJYyCBoEahXzmRP7u6etDzMwPO63P8XFxCdEeqhn0VvxS
pFE7BBCoMWt5hfK7q6olbeWwbTq8bNwNLvcTW2eIstKBePc/n8Hly6WuTOUp0NlK
gU6t9ma9LIs+KYnAgbJ4Xg==
`protect END_PROTECTED
