`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TPl8SGjBhb1n9WTCwwR4WqdMv4OQrW/0EkLnRox+hDYz3RjBn+7YQseKWF/JEjr8
Kf0raAYnCg9Onfz56uEQpuU4+FbbcRT7SbCmsKCikoisaYU/FjzLNgAtuLHSU12k
6nw0jzm6r9XyGRnW08ifVBaeKJrfjqr3OoECW8k3oI/jS1KzSuHEZfUkFDWjnxQA
zILrlpob/JV60ssWFEXp5LGf5R9e7dBG6MsvBSbB/TiieLLU5iT4+9XOlSPBO3zk
OTiLBZavGFZJjhgffI6cZ5+v2w03cRzlS6XaFq3ZZ3Y=
`protect END_PROTECTED
