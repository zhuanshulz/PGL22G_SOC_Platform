`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vMHLsOuKuEEEbvmiaDLfaca6QqD/FYCEm/ywYn6UfWG1A9hpdu9ZuY7N+OQ/inWN
+ZKj68grhRnviMowg1fpPE9Da1pK7SQCc9aVE16y01jdhmxIizeBz9eZciGEG8dA
tMnnV7DVIymqE3yVuKLsXX8LaTGbuPMbxUu2D4Cz+rCJPbAs7MmhrPWdNMdeYGay
xzYUVKsDYefYTRyvBawg/Fr3lwO3Na/cbZOzYe7ESqLi2vTtP4XREotV77DmY8zf
RabNn7ZWLVEHq6nxhPgnQcdX5x3yGOxeuwaP7CMW61yt6ZQcRjPYgU+/ZmPKApsI
ufOblQPEA0lMGJzSb8g6WBc2axv3K78dwj6A2trGYXrNbwL+UCeyMxyG3DGLocLL
nwrO+Bv96FK/ySTWLvT6aXUIDW4iHume4M1a7mDXMtYbDa/Km+1eRatapOxJZZR1
Ei+UXKBK87xn/4imgTEFEm84CW7yzIT7Rcpn5zWciHigxj1bowubQcSIkS5vYUgN
U2cpEExK3L14Jl9WiA3yNNjUXkUPSv9Ro0NQwXrcoqcRfC5uWnTE3UedzzTdcITS
Q9Vh3K52A4qWf+d37ac6bnpSC8yXJq7Y9TKXSPppoHBICXM0UtTOIGIqEaPSmEaQ
6ZANk1Ty2TTr+M1QfvaRa53YV+D5ot516zZDNyhLfb73lQbsk0racHYOVbIFamc3
VK26FAdu2jgYjQ7zw55EmaBYvzlfzJMQURyAImxIkJpVTljl+BwxaEU+6oPXwBUR
o/0hAhh8ljcfDyYKcE1SZV8KBksmp7A4fIOQgFqlnEQaeQfxgMCzeZnqZsrIAHKH
Ts0SEyKuzQdqThsgEp6dJVuxOql6w3KAaNkwp1U1odp5zBZWDMLua4/fpUe0uWH5
SO0jHi+ndF0qBqQRLC/rVGyaygl5VKpFfcITA3MCcgWZ+cG0rsoL9Y4YBoWpkU7f
knlBHbB45N32ZXEQWflrJSyDPKyGctgf6LyeyHjWgAL/Iil0BsLp8ZQ2jDi028tM
T/h6DB/4uomZ8Qe9SR2t0ygFbnWAqPX7cKQykTtxqEd7nhtBAsFeC5XEXSF0ssCu
ZHa17fL8gtioS7oBFhasmXaP9nVXDbrmy9M+ZKMlzCNdApysPryhW8OKb930ozbK
e8stxpr9i3vQP6Mfg/aFvuMwHYzHLiosggAvfBkMeswrOSaVvXgKabASEkcQW0le
mu26o94lQRA0++5E68O2TAFhkS2DMMiNCunAeebuzmh2iAJPh8dIrcKqABtXbHZy
9cPciuzzVZIIKsJFByZv0Tm1ec3e5z2FaFlVqUahSi1uqe+k/dl6lwxZHoigjRvV
ZdGWbZSSyRRk8TqvLbbwd+kgq9J8HJ+ahvwqM0NpRjEAbLdOlb5hKMYzxj96j1C3
xKjQ2CvUapv1A1nLcOxsdBtMvlfyqDWi8cnorLnWnLPocTp5joOZNfiLkdU74qG7
/1/vJKVwuzbP+JSqV+tExTwVK0QIlwqjswbqeoihrrMr1XfFV0uKNPvNDet4+8+S
SFxbqUYLLRzjbbtcm7hxux7w0E7MlFF1wA3YQcCGVc8Lu4OwGmdZjFFq0COz1z7J
NoNFWfe9bDlBseZ+eC2P43uBAY2Xp/s7tJv+R2OHb6sgwP+l92Vbk2e+A6UcknOI
TQwOljr8l54H04BFfhcH9RkI/KOdAvgKXqh6cNOuYkJZ6mAJ5nsNrWrOywucuXro
NhpOVbbBmU/eWuPZBrPCk73u2SrLscQv/O7Nn9M9cFJaChhKZnOnQxbTq/QsFjCz
FCPdczEY0tl6xlCSKgkLVsNPvan5zzCLh9nzanVuBGVUHBM7e5sGN9izsC5zxvmF
643EEWKHLWAU/Evg+PtlyuKQzaujv/r3xAk84dGMYq1ESsURD2IKy2qlIn4gWjTV
vBLhQAc19ejnqqhqlMKck0FK/DPLXUf/LIfmGIEiyr43MT9JPaDxyxyMHht5mzxD
1px5QOVvazhvkIqFenPWlafNNffx/+TU4RHoYI72ygwzhMJBtoxpsu97nOdIM+NX
S4yVAqs1THri3IhW3TR8ZkhYSy2GdIrpPf/lApX1/d6QhF5YFg9X6tPHkkIH4hY8
1tryBojYCXIVrezvxL/alRIrhW2LX9ho2curo+BfKroHD1wzzoJjjZBMb++zR+H7
lDvMvXdr940ZDAwwVPEHLgYnjSL0Uj1NVmde8M2jLPmzsCtVy5+Tkqs7AoEv9pp4
Zdt+bKWydSzLOkanWvSzCE1Itf9k8MWH+I2FIz3slgFJJxWOuXhvdqtoP3P/iW77
ha6QeMSxQ6kcR38q+v74vTgebA0BikeSxOi2qlIP2Qsfg6l9OP/IGaVhW7zQeIwr
oL152n+969GnbC8guKAK+8IRGtvfFP7DGyW8YeS3PR+QX6Up83fo+9RyGFCP1FzW
df0Jsjjfj/M8eKaKuaQzPGLq5fXxzNZL8Ud4dEG1p/S/oZF/TYomtUStWohaZTZU
FRaWlvfTC9Bx82eirr4jknew0ZcgFl6Qq9JreJ0qoNRZP/o1vwnKmDCHvyjGoFK4
ONa8kl0WZSjBjCzASRzJyEwILfWP/rZzO3bOHIA/jIHRBKChC+1LvI1NRllR9lcI
N3M9Snqze+mjroL0UExTBw01HDn1N2CM4tDL0UUydhpbvi+e53vGKnWqgoT9D5oD
J7dA4bWAFeXI/HUSkC8RuLkTcBO7MCXkKy3ADSkuJi8QhNYzVG3j0IBHGTTyRHLr
3dZqS7YcC4E/6KfjolwWef+MXoHzlmaFn4I5WGxYhqvmZYL52jqQwUlt4uEOjQzl
YfNFurtyWMA3G0XnfbrwtKVHTFEf6Uc3v+7PAZOKJ03JzBHwhTIPBGSsXiDg3GdR
mVk94KVVuQ2XisCdOvaRUmFzRI0JLlFWp91c0pwPW4B0Y3SJFqWbuH9esdiFoLYy
Yg/IEIpegxRkt/yJf/ye7LrCBqEHMyr24eFaA/RmLo7NdFpjwI25BImclqudgrAR
EN04QgqHoXc22rEis7yK07GzyJNy1LhbwSpz7uI2L8gs+pVrP2b3xvqMywLmXh8v
s/OikHLdBL0qhz39QQyDHtezMSMj454MKbSd08SrACXTgedvUVuBKaNyi4qNfDzi
pn/zsVgAflRKn1fryHULvB5TIEmcMGk2JZchXYBrztqn3pwjUsOHVsMhgPxJgC8E
rN7/w3u4HFdc1l+RV+Akshe7ybsAwq0AMOC7LYK761yyYKOpkv3Mkvfz1f7nQOOx
BWJGZHMT9dbFAqClf+YptDmCwJ7iMjUbrehfDj5IdW96IQ3w2U8b8y0QGOo+EKJQ
Th6xYSmJFUvRYLdIU/0tLmPwhjzw2fEODJjWxlgn9BPDRZXKLTH4zB5oClvtht4B
V/dDNN4/4bRAcE1Bzo4cWG1VBM7cQ3AggfCapxxBc+xhtAO4OMOlouAq+/JVqNcF
sJMF14/sN2qmobVEf/B900w2pg0XA2EYjm3/usBdenbSVdJDWL1u4Gy3vaf93TwS
FlfZ0vmu51d99xxM1t0/ij5BGEn/iJD3liPYsnHpBNnv7+h5l/MpZg8xL6E/INLr
Pn0CsPkOAAjb1+TOJVS0z95QFJoQwjLpinZdBRswb4pNR/cMr1IxwVOjHUaKFCw6
xSGql+D3tGNtu6U+Tlljbzz40yPvEZkgsPir/BXSQwiJ37QyWN12vEczfCtHCiOO
dKYRaSFH5EwNvOz/xqdg2kTFPT1fLfe8zIMT5ZVqm2Zkm1ZK4H3r/YHeaet56Z03
Ppgf4fU8xC8RqC2foUZ2tmbAshy1a6N5x0G7RhavCga2x2h5qsFoSRlaB9Ff7mym
N+sgTZ4S8Ove76pt3jR0eOMDV1h0U6PtD7EBVMMeXgZz4oGTZKTPdtkHHdXDR+xU
bB9YEWSJ/ecNHWDABVczICHSGgWpbtkxdUl/sfsZMvgNlU/nUEcYfrmTjpohRp5b
LodjhB+O3kA0qoJzqOiH9pNNybf5ebQFlt01zCM6XMe1O0Iy7c+1ifxO0u8HP+Ar
7ZzlzwAKxz2tLnjf1UyXO/5tmVwDaTvdQj2GrxoszpnMiE3jDI/vEBVTvjhb52xj
NlEmPiWDT+QjkPGMgOH56Mj08y9Fvut4HGKlg5C0l7Na2ioth0w3Sfex5GxNPUXM
Blk9iNxkZ4NeUvYy3POP467RXZ9RSUEf44+SUq0A4BolWSbQhNznZQZiQ9N9DRkc
UElV1ZpgGqAtIKjotbAdlJ1lu81Dr9jfjTNue0uFrOBhsIH7T0fwX/rBRVgiuzSd
hg4p40aqDcQdZv9hFhg5YOwNfB7kgclCQ+4Deyt/G+nzKHkP1fxmO9g+tJfDgR7M
2/+f6m0XDqpbW/eaZjXg7r07o52qiVACczoOppHeS0pcCVb9Do0KQMNGf8nv0S42
vsDOKPHJUXyB/XCw+CuKIEzvIeQLTETbzhD4v41Mj4Ghpeq4+7Oc+FN2UFfSABgl
uglCc9CM6UPP0Q+PLp5bYm2r0uGUhMVN9lWEgBJqzn+u1n86R8wF6e2T0Zz9+y+L
Q0v1dJmH6yGwxgQ66nakZqZykh3e6RIn8NCJtGVgYaGRYrlf3kTeYEEYW2yFLZOG
L2om1i4698aTAM5+wz0vREcjuOmuvEV9JwpFiU6PvRbWzZXvOgpOyWyU/fVXOIFQ
GB8eYQAmB0lXN2b/Y/o7TE7mQQvwEt/PvpQbjKyXW951YYeV5XEC41c1VE6oBB9o
ulDNlOYt7dlvuEQmmUSE7IMwIEhTZyNsvQgx0Z4684y+8WxXeNXuEzENqWvmA4Fl
4NCswlslEwRRMuZN+hM+RUa3vTV3BnoccMeL5OWURz4O9vj3eKtV5EwqGWBEhbRA
FJ3fBEI2E2ZSPbyFAGVcx0eMdarA912KlFdrCpa3DaptqMyeMMeg6ppKW33ufjes
BXGKrp1xmggRYx7gSu6l1RQIH+lt109HjAA5rEq2yR1VA4s0Oot3SczSwNb4JzGb
uBA9x/j7v5sT6m8w6WnvuQyRT22CjGTfhpe1zSMYz5w9JPaebC3AESLhQ4/9+Pze
49LIT24myO0GWBx0HjBPz70sbGG3jmLLjTcR34jaJxUjAcz+wbADx3ffXq9n4Yvz
rv+/GSuPPXFZa8vOkUywGg==
`protect END_PROTECTED
