`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6KcHkg9tD7E8i9+gRS4AgSfWkCE9jlk+0mRY2Cmzwe6YQQCy7GtBdDecbp07gW9s
nKbHHd0oI4Jd/zsgvTMN1sxEh484yV+rPYKh/nNQ0DJGgZhzjQ5mMUw341rsgBKx
p59MeusUC2JxB7MvwjYKJ1Y4GRBcT9D3LQ2ECpXJo6Y8OtB8MeuIKaZ21UOnqNq+
aNoe2JfGRj5C0/tHZidU7XCHDKk8qU64cPzDdyWh3405julaijn50GIbsyvn4pc4
JGBvab6IF6Qg1jBp13RnJnAdi1o7dxiSoxo7NvQXLDUv8fJjtS9pJBMifNnZT8R0
m4Cm4IB87bOSkAkmvLOfUhJtCgEjiX7fwhq7xQrooED4hZUbcU1jIlusltmB1DkL
5Hosn4G2uvJXS7RbqGvJO5K11xyRuMLDBkt5nymgKM06JVIimXZMFddfZKL5h6IN
hb5l4wT7YQneOi6WEvLArlZTiptGONZHPURMfsZyCHufy34h+BpdhCMq08wGOug+
l2fO/NKftGtNFbqmFZEvCjKaPL7BIvMAkMDcVQTH/oXEAB95b1gs8TSFlqd4jza6
7/mUKkqUBr/yOzooAuTUs5Ci+RxfA9/lGXRks3UybYXlW30OEMXetuv2OUKi8kRE
NWybsX1afxHHtttkHzFaZ1yKbV8KCH1xntwEIBuVuFQ6vjO73bLeURqB57rdfeCP
kRYK8GC6DyqPIqNcQaY3MQkcGrYlTI0Bmm8zoP54HnhLZD8MaSzUeXk6PIwjYodC
OmmJmD7VBnEcOuzSgsVAfWnm2q66CuvqjU9i+Fa2cPjg3li2N8U/1CBN/+ytkr7O
y6H7PHkUSy8g017WuqXW4C7HNSSbMBfSqLAspUSuowFCLpkTfNeenRT1AI9EC+aX
K3KfCnDu04DMSKaPNoP8L6a/ps4aCGp9f6b/o/FFDAaZZ/Hp/8nth9yh7TPXoUnQ
`protect END_PROTECTED
