`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J6dL8odnWPXnWa9Lk+BA+gkXjeYNnVkXN38gxTT/vPiqBDi6pfSl2XGxaYUWCP25
nFvN1Wph+k7JNWpAMGjJAjxH4fpDZ40VUj7pXnD5XKMbaIKaOyhYyg2mO4CkYhpo
cJm8xW9rWmMB8EBHdlxrhT6APNTjuiJZNkIunlEyoKD740ajlbIhNjOzTwi0W/e1
wY+W3AFbC/ZKPtbfrTUkkTuwA4iryZD0gXS36cv9JzYpT60px6duaA3PMDaCMK7n
Ti7aCH/nK+xhLfNPjrQxLe72Tz8sUtk8rYToN4xPDExEvGYOX/a7wM6h18vO/6Kl
1+Cb9ZIatj8EhcxCD46dUUoZT9EpVamTeI7roelgugo=
`protect END_PROTECTED
