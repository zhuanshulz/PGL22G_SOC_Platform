`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gt0q9Ro/1SagI+0UL0Tr+cpqIXElF0z4QQ6AYGpFRhP3/zZUwA5cBV8DXPje/K0p
p0v99CoxKTsJoKGcJvwQQBQtkhhPqv8IhFkUp4LZS+cRMdFDS37/wyIFS+eKrGJb
IeYkQrqOfq2quR9+ZIgMhtIGRcdnQ3YY4nWEb3KlEQ+RBM3mJAmQAQwYW4SMs9+r
EKLPXHQ0ARxjZ37BwZ3IjxznTvUBNhvR6steETnIsdbdisIpAiNuLxqTrxR065IR
hGM01m307XuyBwz25Sq0SutEj8ktDYl9IcIE/fp3FRekSzFsmLOp2SPIq2i7D5lx
/x/JLA1KaLo4n4VybL3UMA/qGQAHnD7kKdB3rD5KCJXfCkqFd3uKjds7FxxrqECP
45hu86mvZyhxVVK713/jcR7tLW5db8yYWBtzGzMDQznpc/NNaeHvdsFP2MIV0drk
YWGPhMKbzwNzdnpHidEztsxcA7HjJ3xZf0i4tzbKvZQng5QY+94q/uktC72XtMJ0
B0Oe7qHq/HHZc2lzr6DZeQpHvYeyqRRcZikjtw505wgFSePsdg3O9rahXqBrBR9d
HDKieDEg/z8+RLxPl4zIz4BETc5bIc5tipVkmHX82Pa+6Qq9mWJcRKcJRTkqVdSF
mSrwSGX2US85c2jvrWDijwotF9DEBFABOxdd8QzUNRbb4H8jKv1exnYNU5UTMNyT
EqCqDYNBlrc+sEpHzRWjxe1mpc5Rgt9m0hAoKrHoICUFstHFMtOf8w/EMfoQabUn
YjUYWgTpnUL+nHsfYKlNGB/TH7EXoKO3vHfwFiTMgEB0NOwIjT+uud057YwSEgky
T2kgxiNfRvWV1JorW6sFeQz8NE95CGMgMD3ZxoGjBpkOKJhv3XpO7y1lZmQIELEk
IOrTzLIfJmT1GR8fQk8IEelWExURhkBlxgMC3IeiJOJjJgPfXyr/IsW/4s+ZDJ08
QkiG4/83Pvw8/7N3o5/dSEa9xJNjixWh2t5sXCKhT+tafhyo7mHkEbICZYIjHz0P
O3KOQ6hqdPaP0zPv4TnC608tzhHijm904xSzkJZl4qXvLNHiHbUiuF0mOM0Mq/eY
zbgdiRZA5YtERQJJMJ5HR5TWDgFhFSDYPBR2q0gmXQ9b2C4cH2oiKEyV7zftZtdj
i5FkwY32dvrN5b6RGjvisvhFSLHGKEghospeTQzxl94lst2P6Wn9rHEFHv15hOOX
hLfOBiEI442pb2b78DbrvYVSktQ9y7imu2uSgX/cPjKgBaYUZYxTnbYH2Okyfoe/
fKycJU+7/TGXzUp9Q+JGZaR59shkIMpNMDnSpkIodgs2ZloCbaH+fr5yHh2UXQO0
E0DV5eq76rRWiqoreoL/SQWZTY/+x0JBjOwIh9TRJDNT+2HN0iFl4/3s+6MxYIIx
AFMtJUY2D6tp46Umj/wJb9f3e8I2Jm+5nCjNTnDfYWxsg2d8UQfexQMJcI2Jt9vo
9eJI+fpWl/jhaC1zIY2YGkMYohHjJK4KqvbgOrORQD8IxC7vViNbBPqgcV/T8jrU
S7Sw4h54yyTUobqwiCxadj8YK6i3NZlcR9FYpL7TQtphCSaXYTfM+CBUvcUzOvfS
fzdRt+rPkqti212gWLIARZrJd1qIyVXqovGItm4oaSWzeNYZjD3SBubT7qmILdRu
VPwRyq0yyTpMx66Rj49pax0E9CgFSVqz65jmV2OroFC1axwZxOa6ud1mHDaKfSNJ
KGSABC9VQyAtLxkYdZXtsSn7K4t+dLt4/k2wuNpBciZ1Grd8DqtQswzWxRZsjLJs
tJoatDeQ+dDjS24dfzijas9kZ/Gf8pwMu4sJ+2zyertE75Vqt+AuxA7t+3XMmoAf
sr3hOl6esKVfdgfNTHLw/frW7NBMVfeCQvLkuf1VcnNG64p75+C9LhAe6ESw6Jsj
xsCjsZ3KTxhfioX3nvG8jASXyhNmXFUcBhpePvK+KXqJc44UQT1tIUPTjvK3na40
Ia7dW2nZblESOAfqysmSWCoPu6rdIsbwc3bkHOPTHUgPiyy0mps9lhhTDOuRFOhr
W3DcwdPjrZ2mtKjht+ef7fA3ZyFaGP7Sdf9+bIYhxHwUK6xaeS3wNEtlecxTAEhp
eNMgFoelQXzMT79r75gWvCbE/3RHYo7K8LNUlLW5XayLffA+TuhnA2gSlZsNENu9
AH9hgUO2M0tXZigFfKCH/n51T7HKJJkRvEMWYEblijaoe79UFbxpzD0QJAZALliV
k1Qo9wz38GnQ1w3UoNR7DeY8HjkCLh4A+aUHNRveZQas/WdR8uzBkFiJeY9aDoDo
oOWZt82SfTzJnhHPZ98/9WoDuP/ivargrcP6Dtw0agEcYics25bsjetxMSHpdluc
t6meaFGxIfHXPEqWMhDVuzKZQiO3tSFg6htF6tKddLHP/sURHUt+3xqgXN2bD9aW
OWjWyKivMOC7aFljYm9UuP7kUBE/rL1ndi579E/AxRJ96+cBw+jDLXXAD4oArvfm
L+dW0CWim5Jy2vtCjn7qjFIn0EWFxHAeIPFgq254JN/CVryQWw9m+89Ym5wr8oPL
roCAC5/6tUBRadPHdBDCuTwZJNzhd1VNxzC7dz6XomBqRWSzhp/FcarsSJrN7Jac
t8kyYU7cbtowmsLQgtdEG4dw6Rr3qtdudhusHFm7uBAX1gXcorzzTfvZbgYu1kpW
8AstOe6bzJMqGMmrhRvz9vVK+Uwg4+nf0hoHfqidCYvuBLUCA8u5wm+YB3yATqCt
RIKcx62WdpQWhI7/sS8TVVRI3zWpEhbRwRdGxYqZMGLTCU4KZnfihCg8lSB6XR4y
Glu1nqbdScrW3c0N5P1A4x4F4t+HbI9VVYoETI1ZtA3eMQvBGCeAvzd8M6brxZDT
DweXdT41YoPp7yV+vgsfBoyyELYx6MHCtAab2FT6d8yZ6RvhI/GnNSfhL1BXFtvY
QxAxBG8yLD6uutFEg9bz1BbONRhtxi9lksiqVISggm2DMJmPRBiPUSsfCDyy5t0V
xbYYLmP+pKFeB1KfTGD8EDgHMwzqbp/HZwc4qqyfU1FLrBnTWymFU3XnB22HGluC
AKT0jKK/w/D7PEqGkvCdIXDAaMkiEn8ziLU+ToIuL2K4cqlyEVlUJj1bzVC0ppPd
l7HzAoqGJz9QkPA52TF1Pd9HXG5USo5tN1ogOMKVQwKCtlt/46xicNLA6FVm61zQ
K7+uYU5AmvutcNanDZl4kjz6+KaRhKvRTp+Ri+kSulmFuzhXsAWX8XwIszGXK/hh
Y+5xCR4p0zQiK7MyiayN3Sj9i8gMR0ZlnwVmuLIFAtjUEXWx5WPYJWe66z4SxNTV
5Vyjo019/Q8+D6moWrv8zCTOUmiy9cQ8CqEQT+ZxEqg12XjKWzImjNqQ69tkluI/
X+UrltRN/95udNzdB8cwlg49GRuYYt6ogO3/vXTVk3EyLdfwsws35lCgGleL7+ux
1+AWmGM44WYxXwPNVqvXYnkVcUPmClGxmYizMsIKN5CXzOI7d9u7746orLsrhT5t
V89T85zUkUi8uv87JVQmitiNAQ1MWD7l4uAt/PcQcqp5hgywern72t+jeQXm5vMy
iJSByFBwy4xuSDNx/RUGErRv0eYO+dLN56/4uOmPtnGN3Q1ig8mMuJc5qak9+LlG
3wTXGKk1asnpKbHEN10nqZLnHRPDP2KiKQZai7jKmtq7Aqzv+845PIygSeSs9lLq
Pc9852wn2PCW4KNtAZjiDgkYcbOGL03z4mHurLkLiCXExKpGdpZtE0ITNPfSM50O
mdbfDxCaHsX1UYplrtzL/QZe+cNG70j9xlhNoGdZe9svMoDBXKsKr7A1cuRUxqv4
0O1Jdv2LvYWgLG3Sca1Ulkb3C9mYzpW75I+Edls8Bxg1qoBEx9KLfWotcBO3wAVO
Qcbfih4jfKqTUqdAF9js/1qxmbgGFfAX0GwICievc2Mxx7sOvKNhVxwgE4SCJLd3
4xgHFOhiHYENJcXww7Am4mG4y2NmVLJD+apmJr+zvWFFnKZl6Gt93jzgT3DICDlQ
q4pq5BulsCsBLUVAI9C1QBiGmZiVGAOtDeyE0Qa6Tu/1kbDr5lvOgNVZ311Jrupi
SoJ+JA2vxZ+g5RnwxPxg+ij7mFnPF0hac4TfjgByLBRpM1Z1tNhBMarrlkcugA0p
JGj1H32qxrgwz9CkW+PpOPXuXC+Rko0a++TJ2mabrSHpJL0jcoMjDnYaN35AXEBg
kqMhLhYozM4roUsguqwoPPomm/OU1ziscGHY+jCRlj4/c9iqg4YtDwKp6u+fcLZ+
5joa9ErhpYhjPMhaWx1AVLRUSBv3TNZ9+Qq1qLYf0wpiBAgVpRRou3VQ5ldOSCci
bX2TaiC+y5axVQr0I3gabRbhgNw9EUpIBMefFamZUYFOYoKXDb8aQh+6susouxN6
blQNBGEQe8nBIPmxDD9Pz6mi20plKhoIlGlOHyY4nahhJZGEfnUt17DC2UiZzwXU
NvBqETMFhYHp2TmJSKnWCbN6F2VbiqA+9b2j23VOR5YtEcXRgzbbtCcYwtD4hLej
FuK7pg8yhIkMJPWg7FgPSh/VpsG1m1NKzpQaSviPSnGpNoNkNBJ0iwED9GCB4zQS
EahpK4PXUxtV2ehsIkhgcNyOCDkK0NoBPQ8JiRpysupFke6tVGT3Ue0Agn7UWqEr
cfMZxganVLkEDzC3hF5I5ixi6wWymjKCX0T81T8g9mTy6qKohhJrlq8sBt0gH6HJ
qnvoAz372GS2AVmz4Gg91CPj88OWJ4m69otJAcZRwI+HixpjaEvF/ItBx7s2v1iM
ZNNrBRBeOFLP4x8JS7YfHt+aMjhLIB128XnY6koKJ0YUWcUq7BKiKvAFvdezXAcb
KvG0LPhLmiyAfgsQUFA0h3hKpe1Kauf88ZNrRFg7BxsbV1JFulG20XCYhXAiEWqk
NRPuO2keswjwwwDqc1DMN86+XI7acDmO+YSKK6vsgpnanrwox+jSZaEo6McA3c4B
BjgBPFqRJVQn+oYirIqFlilcZOA1L+DGQtw+rNgJ/C0ugz+j9BtkdBV2xON/1GGP
KbUPbsVEmHcmG+kK3nR6nnVNkgJHMcBqbQMfoHaH4DVgRR5dQ5VMBCBMnVcAG5MZ
38EE0RK0yCDT5i2omMqdCj9fqKDe4rPx9KPXvBSaJOvzYef1PwtT5iMJInTkItJM
qewVQSKMcZHJYSpcxJGpPPwD5brLei/+MmMD/Jcgl1L11SKcjXmfNbabxnYMs/Lj
1TXsAQInasJHqAzXs89ugiwKd+9oLBc8UwxNofOkP2tp6dLAlJKMgnl57Celehrt
5leEjPIh9+APsjOLz8YxCFKXffsWGxINjrqiSgW5dotKqBGqEr2MHbEpV4BMvukD
YJ3iZJ9QEk2PfDdzx5WjTOP4C6Zz7RvGXM4Eit74PplHsuvd02idUJoin32D3cNG
CXPJDRtyl4gEjZkfPYamqz49YWgTxynzEe1i+PDgRJ0rN/w9jk6mGcGUGtpg1TFl
gEBZ2hMKDJ9cq2kIqgjl4iNmZYDZ2YxJugsQXVcgVt1McmRNDyoLqCFMWkr22Ofm
5A5z5pxC3nwUgFjpjdY23BQrizMWJZuoHIdIPToCVkX5W8x5VopQ9AOgBHf8aAPX
/Z4YbKKRwSvme10SUCI9O1hdXfwe3vKLOjTvDNdQv7yzlBvKW/TAFzK0UoqdhBmG
H5C37ToRbfe1CLWZILhi4g04wo1tteIpTwRhqeR1lB+IUJmIoPZBj09AZ84uhRl7
9e5MZhLWPFQBhx2C0zI69VH1vVeRwv+4dc9cON9ZG3eIlg/G7qlaEId4apft0+f4
JTsENbqK1BQ15wxskFPiNRz/1dNoQeozXyKqQ4SW8r5b0JHCNCYC5u9qj/EKFXa3
l0GCUMQbbeDmKRnlHi0inIasduo63q8xRr+OM51HKWdrNuHLyKWk0RUje4KFx9BF
JaxphTKlo/YG7gGWmXZ9FuQ+VXpdNTKNlYBwiV9Bg8ZHH/77sL8Xk+db7FCZl3yz
Vx2x/LSieIr4YoCqwefKs3LRMk2omSVBTKxZV9//KQlRZ8/jlepfjh5mUQ5pTU5A
pC5SvAFvLHB55rAX6hOeMu2NzSER1tN8A+iVj5pJjRG/xx0rUvT8SFdLWFuMcIyD
zdcjX/GP+yEA104pMZDkMUx04u7V4AEAEXUm3RtyB9nK10YYjI8mLQyuTCxlyjHB
FVPw1L9Yq50HtIxoC7QltuHPo2pXOHHJmUxNl+OVKZLiycaP6fbsLpAFLyg/PwYJ
iM1iGRq0PwOMePYizQ0ZVY6pu2SZ8Mld1s4B92qWtqKl2YhyVIqefO4WEREAMG9Z
zXspwDLWizaZwLE1AePRA98v29FJFozZrBWyy1xfbQN9xnLH4N+zpALH4srf+WOB
N1PKVA7de4qaurAaJdL0sn4df+XEVrBdzHK4kornp0vRLXcXeIXwWCsDtQF3XJdD
g0QbWkQtVCZDElHqzJ4rutaYclqrkaD1lZKJHJpDYjaJim0A411DJS7LovvjbB3v
m6xrSBFfmN0wzU8LU7tGcs9CSdw++ZIXlGtXRlCWXqGi8Ni33Y/iPVBX19Qcg7xR
2vDdlY9nwcICbo27FDK6uJjTl1xn/ja1Y2m40kPM9XVDNup8+hxFe5O+MxHtHY0y
HJP7iHrelQVUPr/5Kojgbr2d+3D7egSSEjFPX4SRtNWox92TrdQ07wCQRU1IRDFU
pdN2Iv0+nWLxgosmQUkSwOTuwtEkgVhSw/PbSap6zDHMFWDCC2zuyijMGjupRB3L
//IQGTtSU1FJqP67G2catopoJrsNgol67KLvoPwpVG7ysIIiSjIK524eZXr/7PPD
ZPu0rTHSDNjfJpVxf/erw11apW9GirepLwxxGzQ183qcLdn1tlbOsfCKvem0dENE
e4w6btJwCewOK9pFWbygp4XasA8nbdQy1QlNKr20THiq6sqja1+Tp6KxHdnYUbrb
O532mxEHMWkEtzUQ4EW87JC9aK4pqXc85SMNEU0G69xFRzFnibIW312jRKM23jHS
HoV/W99l2Wo9d6CmY8rJx5wMVgqRNmv7+aItBryhNMYGFvOyviyLwS9AJKuuzx0p
KMehxU9tYCZWoHd8Q76tFnLuaGLZvZBgxi6e0Osfhg7nDl+kj9Rkx8kbAF3YAPEh
rasLZwAIG4Uv/TDaImlhs4PT3EjcAIeOVNnUo9zdFkacIS/DWEDPvpE45WFwqXFo
58EcYoNjachfxsiyG1OtBH0aMCPiq0pn36h2H7bBnVqk9UVfXW0ZXBneH/1n0edj
Ts77wWDxDA73psYBz61REAwxPnZPYIa/a8wn8D7QzvQqQUUIICC4F0ke3NWBsoHx
CaUPLu2jREsrH++mi/52s/N4L30qAlxvtisUa5Gb2l4TwQz1Igz2/d917P+rEuPi
xjaY+Bj3a9AN2uNapC2Ddg1EgQ+c5NmNqId7HM2Yg5X9coITy1uihY6h3tGjBAT4
P57WAJ9Gly69iidhmLbiWvzNp84umzDHgFdwat275XThAV+2VM6wMDvu3NlgXyKl
Vdn6jY+HJFgOsj4V+FLQCm/TjPQF8l6uiPTl07HfZrz9m6ixLbLZr8s6SlBNIS+f
mSVP1VO9+BV4BTVEKUl/lQQ7XiFWO8HPzotfl0iLaiYkP7+Z3aQRkuZDxbmJBJIs
R7x73S7LJPPf/+Ti9Hr4Kaw91NSOP2UfIDMyRK9O6PACqevnlinyQSkEhxxpFUA7
kz2ll66QfCVZLdhTHAOo38opbViZp8jeDqCgIvijtk2Lor+Hgf5NDRU3s7oLw/iy
xvW5etns64FcX3zx9zhfJ6WwaiMdMe27KMcMsDv4cYtSSiWgoJ68rL0TXl7XY5Jr
yYtJRxRFLRiecBvVrKQdWGx4Tdi9wuVOsQJ6+nkDs8GR1aWocQcBVZZ9IXySq0uF
d7WQdGGjb2tgLa88Rc40kJ90hjii8yh/Q11B0ty5XUp1qs4mQl+ETqDEUfXTflIO
G2uZzlEsKKo0ZMsP/dYJbNQdzzLa59fBmvu8Ep1zYwLF1qrFPGsnpFwpplyvH342
n5Z3lrK6ly2HWvw3UFiYryzqDQHokY7UP10K8uAXxtGcIIN+h7Irhhs6VbdbBPOD
MTXbyWmzWAivUeUqX/WmgurxIGFjgWx3ejwjI46L8Y2HGpXgcfch3tqlvIC1BMCs
sK4kwZ4jmAlPnjbRKYmIwn4cuELBzVZU81j+WwXSktd1IFejTaKXc00esAS9KGfU
rU2YMaoRQHLQTee87J9daisReMkx6ye0JXtIeS9UvM3t6oXqrXDIm9jLCMUZ3CfR
r+fd6MYkjoH+IUny2Z7Vslwm+tcSCxczPB2oA95H5CA1jh++ePZZkBCtsQXWwQni
naqZfVITh8gvWWJTH66oFifzgk61ah976KxIai9y4FjXTvqw0hj8ZJF9tRKq9FDN
tWFHbqnNv5Y1/HffO/UNn/YWqzqWcuSl1u+2SfXndnuZu4HBWVUR7N6NQp6qZvBi
n1m9CTos1A499EVEFRc8WKxMFS068XgbDcy8maPR8U6AN6OWc40jduJRyTJcDhvN
uIQq/dhR6SHbt0TQD9habYYXoguSaowzyhjKtolIccRCMj1GJunbhYhDBdE3a7Xl
4YGc4c3csZdsJ1ztzyFV/XX0JMZ02uL4c/tpglJ+c0BjpcnptM3Kig75H2U+0FuV
i9WqXMGkCz+I5bLRlz+TlLIMyVJ9DAjN7tlKUCOWkcTNXkMxASW/ItEZ23ebwInL
JLtnV/vwF5YdhDWraHLWGcWV3pKz7ohM56WMzrEhZyF45kEpBZ0lv08V2yshBqaD
I3ozVuwao6Fe4VfLqZPs7sxC//Ool1gDmDoXByWijZb82bfhS0aYj7NA/RoxKnwY
nHMsMTRolGMPAivlUklmaPka0MaeF8l6KEldDsTBbLPZucKHJktgae8p/VVPSrxg
L+Q742X7FJDCC64FqcSKkX5HF88yAeIQQS8ke548ORCEe3xpNjRoWxQl0eEW3ege
Ri5yyiXPXv8wdhQzBhIsLOjLCNtQagChxuAts8mQR2cHfvMRakhHYLnNnRysWLmX
xFzIIw7nGLloHppVZ71x2VACIIDEJq7PYia1ok4xbUJs5m83SQHneAlxAHyvdmUg
WzaGM8UUbtKlg/qOBB1F/dA1L0drfFpP+4iihcOM8+F139m+LZWtVVFN5VuIR8Wj
D4bWCqXVQ+pa6mKPp3gkMD+HybmPcGUQ7/xZ2hlKXTmODJ6BxZtrdpmVFH0j1Ewl
oAseeIRe4MFYS1nZarz10OAPNW7n0movV17VTL6TqDKwDSih7ObzgiqxceSyEYIf
5z65tNJ2B8TWIYzjg5Rw1wc6T4cZurQqim3IYm30HO7joxhh8RnRdtWw6J9Pm/85
oQb0Hw+qVExpSIk1cO6U8SG1qs9g7+9/oed9olQi5hVw7YOAqNklJE3tj+z3xeNU
O+oJAxXLJiFd8NrWz9Uxnah7RR4oMIKHyT21U/sr8HBwCIQh5tqfNv1wye5630qN
ScizswBXjdh44CLHJPBK/OHRQ8tGLAPdVdQnN465eDejZfePiFg1ZAssWCVoFxt+
R1Fxz7VcITgM8ZAX4z95L923skk7+57HkI6w4yqIZV+0Nwi4n+xpMOYj2v6oN3fI
2m2WR+z7MoKT00uQxPTtWJvckvs1ENlZJtg5BFvVHFoaIYX/sD1ChF9i7E3pdeuH
gbAl/5upAuZZnJG36gErGr0D3sumCZ7LkTPJvgShrF666VKaFYxlspwKG6JNqxhW
B/pir5IH7QymhjVymsPHnkWcc/cdgYtbsRYP1CvnHqcgOo8rX792WmV6hh364Ni1
ABPdhvwzn9SYOmgFOiSoYhVNm2s8z9DLDgCwr0CO+GULialcpeclqIkjGwrJ02Ww
XA1X87q6Y/1lhXnSi0W3mWQDcnTquSXJUfrz9oatDTVguULIV25RQuVo0/atj80g
5RtGwyskLFP0+pu2GjBna7BOEldBHP9mKcKrK1lbW2+BGqBj6WOwKve3izGhI5hZ
gFxaJdIqR00WrF4Yy/Oaz+pyMXxSyxO6F29BhVSUWufnmd/9o9Axedr93buMRcwE
7CXN7PzY6YDTwx6zSMQrfxEbO5p0YzT43nXyNOb9ssfVf6ahD40eL6pye1fcjBiH
coY5Evmmoyi1NaoMQjFu0jjxtIAO0XtVNw8jVE+yrPc2nT4EBh50GOAdSt1r3Hs7
SxUIrEwYx0VdYf3uR/eld8k9EOrDbLuqClfp10e+nM4A0a4mdyoKmjr7MlpZ2UzS
ddkKAplFawhl1XbVGuyMZ/fy+wfOxlSy46rL3+syk+tHCWuJMA5cOUKLZz7cPhls
4cLLASTk12AAKz/jfboVch0aFsyl60CUSlGe+pid1Obi+WcTaZwVl1xldvfONp8d
sbsfA+Ia2+QOnjgQQwI3307nlScm8JC3lPMVI78pMyJRuplMMT/sN4hkSfLU707z
TgFEK8LJ09L24wi1hnsFQJ33zmAcZNp3qPnn/kvxHmQpNvH6lx+U+eApt4n4VXij
8SdhIbrxVTSLxcJMNI8Tf6NtcwOUJwLrV84pdODtz6ECGiRITfH06KhWIVKUPzpc
GY+NdCFsf3t/lpMdgtAoXx6KVEnNWva5W1eukWGVL2X0tM9xSyFoPHaOVAeIJ7KN
lNneoVcPFHUeQ6hzyHGk8u4J0Ubdo2DkVTDF+TxuXsbcyLTnk0F+Yj+Lj1bO+67I
5RFfz+YMjvY8GSS1QY7mNe+9C8mG3SOHbPfMDg/9TtWgsxDE39sgBG2Ah0Ertrih
maVlce0nkAz6/kfGM3rgHDDgVJfvTTggd94PelTtRbYGsGmF092RxpHpWSgvZ3bz
JEaEf3FoDzG84wNKcFthiJmAkBB1Hah0Ca1XaxFE85tgc4PM2UISU4XwBTAlEmjw
xl1bN+twsoWCDYIN7hTiRJ0YL4BiOgPPhMwemQ3Kqe6bd6o+B22NcwDgWz3gXeVI
Lm/9rLO2g/TMxsAqy+Mi9VRPFJ2tP6X7Q3PU+pD78g7M9kCrgD3Rdm5uVsVrwMXt
I7L3qHn/pEqeFinqx4CLlK8OOy82O8yDs3MF9zjSAtw6H2aR6y5tHjSQ6wgc2nn0
baATShv9oEotKl7yTPeFn1k+ctn0oSQaP7Yo2shz4Gmf60PQKRJ644KKlkz3xhEE
XiGwCmbOyhcw1H0sATkKIJDJoVkdTA4cuIQ3TICIXXmEUz9OlqY8VUpnYz2soCa/
seJ/2uISVOlQbQ8cL3guO1D0MvyDc6ykwWw8k+7PHUQ63gEyqYfy92JQJNBHFvc/
nzLXnIGpVeniWG4155zhBOXPhf2wI7VdSzZR3ZI1lIX4KURDMydU7BSLl0tvlqIK
zUkIZ6RzurPi9zO21RD6Lohicz867ZaT4E0fVjQSJQxfKUuDReMPN0/VVwEATIvn
nIWH/sz+SWKgblJiLD8Qie+i+ggbTqbKhEq0r/I+Pj2DTRLEckLB9wuuXyvnnW6E
Ev1YJm1WKqoyqpERlYnEls9PUeOaXUmCGho73D/BdhWKEiimrUfXCQJ2+RvOOaUq
PBE5FbSnq6brWYumQnLMRERnmhwQAl9XQK8P/BHRWNP3s5to23UTDqL0tcaigoNE
lFHacqt8XiRzadn0Pnpx/zb3kqmZCobz3qCrT1VMirWjzuQ6QM7/0Vt06mcnxUAb
qqMwUGgn57itCr2v3hSMaWo33VqgWvi+uvJg4pFQGYTnAPBuIv5Quk76m5htc/C2
CvZDG/xOCp8u5NrFPt/95Hva70pdbpXyiIRiJD5l7l9wKO6qRyl0v7+LEaggmJbs
IvfrJJU4Yj4riya82T8otG4HS2WoYvXEMAlb4rwct44U+L2j2HiF5FVhACO4c7k4
l8cgq7+uQenrug2K8iXCcu8qs9ZW6+1j0IbEyxOtjSzrGJKBU27rUBKlnNyu4XGl
bkMfYlq8qgchhcDwdvxUWo5bg+6FSQxZxhilAt92Lh92Pr78/0xfqin2gE0pc7JG
wSWyXe0Qf5SMgza5NksydP/xT8VwmE9LRCAavkeuuhg7ANVSDJcIRy3qPy/+YMsV
pqQLb6ybBa1nILwfOHm3R0k3EI7RXwJL6wN2CYrOJtK5z74SJDcsRwBLdW6qMGoc
Ima84+Q8AKwTljVW/+NWyMcX6Qwq20HVSpc0yeLvhB4a5QKTmz2ZK9XzGLfk08DC
2xZClFPq3HvmzcxUZiU0FP/ZP0Gv9kal2Q4uNO+ZHPzf2Ms+m+X+JRjHtm9vrmkW
6/FMSya6xjRVqnZTsGz/xAo6+y5mNjMoDKhEqYAWyfooIIvp72bCH+nEsXKrSBSi
JPuqhS18ODgJqlr5MYrmhGubQoWKGtUaEem7zda7BYplodi62USXn9kyWLf5qNqw
fP6y/HmcxEi8q6iOW7TWTkE/ZSVNKkudyNVSYp8d+/T9QRYjFBJYXh/DDSq6KkH7
HlxPRJRpfONciAojD5IX/trB7cfWuFOclBQuX0XRxSPo71Pgg+48S2fyYncaaPzR
vcQEE9rmQO4mQ787cyUTlC3KDECJEGPGUbyRBIrkBgEjpbPqCwU1elHJ408X2Fv/
sgL0zTIlpYxAKd4IjfFqaFhXv0Bx4poeoEofJBnP45Zzv7fYsXdfPfAQvsNqMJ1b
V4IlDFA7e+cJnbrUoi87VKIlpoyL1zp3kKFBj0Cd/aI18W1dL7zCGE3amAk058ps
Jt0inl7k2eWxf2oCHiJTI5690lnLLRFiiZRZucYR41d1iKwDJ325JRTdJY9ylFps
TCt6VXrlMar9z9++ruk+XUEpRsjWwGr94kmFvDoLpp+7HoP1JPVk14rOj71YcP5N
sx+xyIjB0IdD/Vt3BPtQqHDT/YN7EH2Yt3abusPupj4iYGbks2QwZ8YsgVcQQxUz
tK8rxgdxWrhbXT4LYFDg0C0tuxTs1m4w+oJZyfq8WPqf9REtRjCf119CDOS71lh1
trLM7TYHQZgKlwCedpXnOTMYtsycfKsBhGiuKq39fvFfpStB4Cjj6e4ZkgAFko9+
bpbhSArm4z0lkCTIWn37QqMwbuAkJRn7EVHuOoCngzbK782LIMbDgroKX+nFkn3Q
aQjqSbv/JlSRDICfMv9Aq4TIIvx8LJzsExlcY6K2dG8ECjpwyg/Tz9ocvJVPcMLn
e+9mCtGhb+51nVqqOc3BCajnX2VQmgE/2/WTFBlUvFY3gq0jqmajs3X4myD2pZyx
vzyQLup95QbVICqJcewK2Axn3hGRAPNgUBl6xAdvxfLc8mI+76bMPOprx6onLsLf
NVfjd9a5fF6JQ5nT5U/82+PDXa60HcQvFfYNqpty/Ui0QRkVRwyE6zATPfZhQ1T0
yHZnhq5TNY6mctlUidB5qCMdgUFmIpYz6Iz87K+8oH6bKTqlXegJv/GA8juQk2hT
Z4updKuaFURy5QiPr6Ukq7k9dgPbiW7Powv1oaiSzRVn6dG0M9Pr1y0Q0UbZRnHT
oNIpkNvGciveXh2nHpwKMfDKoZsv9w3sd0OtoQ8yT8ipVBdIUi+/5+sUWkOJ8SwL
Pp99RA4TIH2s6D9u7wJjB5uCevtLY5fBgbD9UMS8EnxqDAwdp9DlD4I50LR6CYi3
4ypAWpy7tpYMq6r/SAFryviaC3VN9hPp0hpA6Hc1ImTQyPTJkziPm2urr/U29Ogg
1Y9bH/1qNJfzg0cidU7xdZdluBj8X/Mbt+wp2Ysk2w6k86sn8XCO/EwEQaPpGzeg
NiBQralEhdrg2XnoRb6AhB9c56bDeX/GN34p4MKQD/f2w2Ksdfc3gRo80rhZYVoS
L/sxKMqYwd7Go/for+UBMk3eC48KDV85TyTBPxEa015CcghkiHSudGn2K21mhjyN
KGCC1bzatsRsRAGCvbnya+TX/ChwUnAZe3HYkky0y06deA6Z1OM85vPz31OzVWax
PlsEe25NyVi4OgAiK3A2nXtDTlHRVHg93GUzSzBkHtgmfyAOSmDiJ2g8ngRAnJ3L
CAiETxNnVmdLU9RcZcyb7ScHDh0May9hyKa2BlqBQpZ73mQA2LegVLHvKEpHkVk3
4Nqz//X/RsDBO3ErRXKzkxTBQa7n0nq0L50P0OrypcqlpsZOTfYdfnC+7Iref5DT
St3yDpijFPYtqBu2aCsHTAr3EeLetLCKmsw/henfrDlLlzLsKufAs1VcD6xypaHB
PuBjwfi8DeVdo+O1eACRO4pbUaExr+3VQOb1EC6khczHCGQE7UyeXGZaArbL0bcU
ohGx6r2/c7l0Bp5SivuViE49zcI9VZCaQLc5MjAGdmZRBoCO6STLZO7dfCoTa7kw
9Wtca36x/IpTjbK8v4gx8qHYmJKO9yVsC6rbpi6gEGFQVd3y3Wt+fosJ/NzauKZX
XJeghyNrz35Qd5wHWJOge3QtcOMrgFKzMXOYCa9pkSuORowb9tNE8JEBVYyz6khs
Iz0gC5Uc8rdAs3EFe7IIPao9itz4MvVkuEnMx+s8yOMkT7lbz4QLM3nmzPffgVLu
ll353Sm0hTdjTiLeep6YAzzCfxBBKPp5gnRwhwf+R1oCajy5l3wbNlu32FtkBgMv
6mXEI7Gye4iZanq+gmqDIE+JDbHzbT4NW9IGatpcH+E=
`protect END_PROTECTED
