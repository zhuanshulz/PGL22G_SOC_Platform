`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
va7Y2IZ4xJJAthStByp3JDwBMKdN2Z+BPxY1TZTa8on4u2odRiDaB+yExtAGCopo
3XPv76goVftI0gT63fqZHzpvAqycbqV23LW2nr4fKI7P9jV3vx2BDrXpKaHOIXsu
JLTDb+a3IfjyS/PzmyYTWJHaadcBWJy9pydXetihJ8rsTbUkKL6KlyexmgksL9Wh
uv1tg2crjmLTHNdFIROSh/W8Qo1W6kXmzvchPLNyBBdDPMlvJyKUAthoROqupVey
WYsQpNff4xhC9ruIdLtVZs5ykW4pQ/p4CQEXHq4tVjXU98jyxc0rfEWHh7CPWqGa
LPNiBsn7fGp/2WO5oLdxw/09GOUe/X2EmlPU8WjR6OTuBziqS7aUJ667i837bzAS
qeYZX8UcbuL4qasli+IZSPh0GNUqvIpojVBgjTN0O0/q/NPMtTJcl04L4MyezjiB
tiUuYQtGw0hhuUGPGFfjARorv+2PISQSvGEJMRywJdf8oh0qGcIDCRLfJJ174TiD
vcPk4XvfbuYeoi6QOgABTgZckTVzcH3ChF3cf3OhSLfmLRlqzsyRqQWLwEY4kGdE
puRe8WLS9/68nNQQjpRPXcPRkMe0QnXSEmiFnhX7eaYequUiROqK2IJYx7n+ms0m
KIgCCgfm7wZFcqTdICQkzVnJL5LX5cdylZ9P+3Itz5tMCiP8nWMqp+yJe6HN5gD9
9a0DgjDGXrjVg9qodd/HsyB49KFJoOmmfRjC0Hy0/vVjIutetLW+lMrzytwUpus7
zmQbfCiCWqryrTyeSIN1Dkq6mHg8xknQ1LvLVpo8m5CRGvLa9hc67j31DrSlDcA6
inSc/VnKo/z6SSjxriI3LDMRaEacwxnqPcXHh68TG1uyzMbGTTOvOZyZKK+dcDKW
GH1sQKe1Lwan1UFlXVbh7pm5+115gmEeo4XYA7PJq/h/EVBLFLFizcNO2U/c9fiV
Uhq8k4opdcRIYWq4qnUIhbbicxLi4ddWp9L+x2r6EKWJDB8+mQ+0/6s53fzvt/Jc
tJ0yevVcUwFDc+6+TA8RV84nb7gqXZ/JPYCyaVf8q3GxYES70NOwUrFhjOhddkFi
szz/7KPtqTPVH/OfUTnqYr6bN8DwozK9BNwDh95Smpx0QirvjqnogBZkYEmBb9oe
jHsCImWfrCR91wEcHT08sA==
`protect END_PROTECTED
