`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ydWla+hXfSmAQT78OODkEUty04+wknjFp2g8+Zs2Vpj4UwqbIbaMLAI8qb2uy7eg
CN2w5MHp2vsjBrvjOQPU3U+ppfMMnXUsrp//ia6F6IJHS4fwGTepm2zZ4OXkSOqJ
MNm5KRym0hMePjd3QLDCDK0tww9x6P1N44BVChRSGOhnD9zqvB8noAxjHFiiX2z1
5qJ7sJQIABgDbknQxZk9G9gmJ7e9whXw4MVag4f7QH/l5XzB3wA5S86FFV9ka0gp
`protect END_PROTECTED
