`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yb5CeKT6hKrtrCZVRU+djEvd2HIdaCPkgUk71ddmm/3Q7hRLTICYaRxQUFzaDzGO
CG/ckNPokX3XXEkGpu2UOn5p+TdULqHu3a/HE9T1In36SwB1QNM8OeTUdrJNbZfF
wJ4YHhYgVgmrtD+bOWBMR3Em+WD+0L2aLO3w1KuQQflWT3EhbfRjlGBOt6OwS0sa
cRTNV0yVsLRuwdQTBIwcGVbAWKkGmzrm4p2jq4PcAxK5qvuDg6JvA4Tf/ektIkVK
69A+2yPqcAqhzZdOwiOfFRp84UhQV0j0j+BAHsVFqf/grqfzWhjOCSwE93/IYhl+
K1V0WCc6BXEPJuL47uEcWQ7Bax1IIhCoHpbFuZz2LgLyX+QmLcpUxkVYhx0ZtAYK
OEDaQkIRE6sGAm3gSHwgq4A3zQjAv3C72FqvUsuvcytFiq27Xc//ZdB/cgfuiYi0
GVPIsnvvm7C+HnkSf/2Uv9ZRGBRLrCHGCv0SznlCCDKba702DhrL03FMLPU21COs
K9MTGydmNbWLw2+7QRlPcRSKwpfK7Gxz4OrJonDEky/Lyvs8t37Yy/j1r5XvfAke
8hPXb5KMbW6dkE4TJnYDE9O94MzpDzM90IF6N0/pH82EyCsCwTPHaxaboPR1QrkN
avqOBncNxpE24E9LxonWpFmsuOY9g7Fi1Y4+zw6RQ6Krz4PbkrH6PnqzKdIy6fFM
ZPha4KkLKEkjfcAVoRVn44qSBnf9E0SXVapKtTgzBTXrtrJ8nv8uRgTLHBoYzyKb
j5G67wY7qMSIvB+4MMhZZKoSW6B5Yq4YMOHG/k6vCSNWaepRkJpWWFN85SeSb4Uc
9N9Zb9pOKLgNBRb8ExOmBzhkE0IKf1tEuoOBFgKbiVIec94Wv8kjaIFYW3APn78j
CPk62KZH2A3mJCYNwOhlvLI/uPrOJiVcN5rX4/01NqmFJ+CVFCN7ytNjKGXgrQkT
d3tK8JychygHGNSOtoWeLaSWvi10RbPuRz7EFWpdkMAxtLdfop9B9gkveBmifadA
IX6OITdW18VwHwlMsdCPo+ljONwa8p1z9N3Pctn234EGcj8akyQJnN6pocgDmeHE
/SwlBFefqH6GxZod3nV1ixaZTe4x+9zYrO9bl+/uzDfLp32sxaInAjEZJ+YEjOlX
KmjM/oi0LrhTWtNFGEafWqyvIGT2U643mxF2XUQBqXs6iJeGpfGUnpV81OgvHnC3
EmEJI2M+fFPE44gujE58xQrlzJggaLOl84Zym2zxwzNDR9qSt1wmTs6SpcObxkfF
`protect END_PROTECTED
