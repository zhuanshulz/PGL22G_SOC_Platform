`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zyi7GP88AdgoNsVMxPZjPlR/Q6wn4tb+97+ok7pX9YZ+GmTa9u2JRmxaqCrCWy13
T+zn7Z0R8m9eu/b3putnq6FNLSWToaGXL1oxN9t1PFt2nprmuy4hyUTk+2BJqdYD
c/uGIYLDqCFxyGjSMwMNzigji47aeZiQK5c3llWU6FPpol/cYasxopowjITFZriY
x7dVnpUYEPTqKH4P3J0Gq2hRZa6lmBiZy03RJtcwbAU2rDf+o+54/x0w5yXt7xOR
ryH7sEBdfXL8MKupttTlbD45s9tPLS3bpw/KDtUFqxnir0EuShFmm1wWDS3cwsAh
BcC3OuZjKc6pqo3mR08CtcfGxx5Cnk9X6Ev1sEdyyUAAPPIIp3OUdn0PRlGY8gfp
WqUypYDXltoZq9nWKWiUbQ7hHCg1ScsotlGKOVGwRoIza6Ybnskhh52oKkubesXI
FqaX12bcRnqC+03uPC1e6VbpnmVZCOIQzuUuRqpRZVi90olWuQPs6gv6ZeGSqnpV
GCFhDkt6u+SASZENOQrytyDlH/XNQwUgt7yUmoK7lliYa2ccItq4fzqzakJkjp/o
lvEsNdcqbx1rlT00+qmP3evRt7dyFV/r7FSJREMoyyS7FfGI0Joy6EPMkRUB59Gl
SITzh83b0YmzwFg9hyCHXGi95KUpCtaS/9dT+7E+wJ4GQ+ywUTtirl0WqncPNkT5
cKA73azWlH9UJ/roX3SS1ZUHYHdj2XoeKhi1ZGq6eYg=
`protect END_PROTECTED
