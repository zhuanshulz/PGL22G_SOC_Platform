`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VOGsYQcFoma3wJDO9PRKta3JAw0UnkdhkMHBxhP39l4x9ps17Dwzdh5oLlKxfmvV
6dYkP53n8luziX29RGCaZVfnVZ7kweQ1bpYFGTt6XmS9VbauNKKciYgzYI8R3XI6
FxMd8Hoh992VhkGbqL92KRls9sd0V8aZ/LcHwohwSn6fTQVfDrvNFDix3TvMBM5q
C5pi/tb94qvLYJOp0yEzCmV2K2ZKU/gydIRODSqi3uMOYgQiMxeYCrhAklt5BbtF
ne9Ni0p4e1xFjAEOr75kvI0mmU2Trx3ylIBHMEEWmRCbC0zaK+ffpdzdqV16jO2s
T9vw2skMl23ktuN+8wb6FpcyM1c3QZXlZxbGgvxCpIn398buuXseQIbX2zrjQWMs
Eseia4AYcFIairAvlBiJhMNH7OHEvNm1LC8XLYeVV16WaxCQJXywa6Q3wwaLHhnZ
/pCGL1vc5fqasA4zdracWwUhccbpXf2At8TeSK0ybkUoTes9wACjqXmkYn69sTEi
rH7cdWDS+wKXfZZNj4xK8AohGFTlUvH0k7JE78QES9VQnytHn0F98UtFnjIJkSLk
dY7VIwSg6r3YB5hMjuvQSg3MLlkpH+FYiDeAp3t6galyhqwQJnJCjy0GEz65Ykza
R+868kFYS19wqvFYLnlfEdABa/44DQ1iGDivlJHk5r3c1KtDFyT+AAsxzgF3v3Ns
`protect END_PROTECTED
