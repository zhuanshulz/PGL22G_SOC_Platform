`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iR8LjYOZH0kKgUHCMQh6v1bMA4viDRhfH+/1JvJAGfFh9OR2iLClIkFoyW5cdsk3
HbjJdFyn7MdZM6hNVuCggimaNLVc2u35dLeh1CAQEFv3oFmIBH4Lclf1UEc3Jztj
pF+MQFsd/g/N0b3C9JyaoJoXK6Qzptkn1aDP3lUjuBdgihBnuS1r7jIaaYFWvOxA
720do53hjVKv6sSIGozUtSm9R+fbsURnyooCEfZA7ZbjMl2LlUJ8PvG9OLG1p1/o
1nbKf3Hq2q0Uy3hH2AvRnIU0zyL+7lVTRxhXEVrsOy9cDcJRrg9cOwJM+KXx3IeO
GgkBnCIY5qQZ00JE9BSul6o2ubeH+YGh3nfA58+YiWd4RueG2lgkI0JWdEQ02Hwj
r0hhuaB3D4bFZYUK2HYxCA01eFlbaPyVMmIvHZw91Tl4YLVziPY7axLWvPjpE5ID
Bl2HQVo8YtfWASYEFMpBD1PvnF+u1FGCzSsSYXKctolrlYEpmCtR3gGDjiad+Xqw
rdr27UKO3SoXA3JwdN/ZyT9BDW80cGZP4Od8O+VsqJ3mpeI5YSwS3VLhMPYHF1wb
Wg87h1ElFLHUkH15mle5a1POvQ3NjV9o4ByeS3JqJ5SXwKVCQZC+nkkwJoFldlyE
w9qPKaeRePVqNaXMPjmg0xMM8NbBJ+GgcPz8QLYXL0NfOTUlBhFXiHkqzMuc8Fud
eSF7fuZwFt7b0OnxQ0sMj+HWjyOaolwedDpnweavPKb8T+I7BRfIc9rx+56vqtlp
Io/qbOhnvnZpXDlJpwjVVhmbfgdI9Gj8DXaAULZdCWUgRfOqS85Qig3eypzsTFz3
kY55x8xQt7k1N/UKOQepHpLf2F38XX24Kn1yNfbcGqR7A2TbAMhCa2jfpBw8iYyt
xUKaW+InoV37l+X+9xl/YwU2PqUaCZDolAV4YiSHqhGOOWnCMaLqkIyBvvSbxvsm
f179MLW8rdC/GAGN9qef2HXKCyhORqliSzBXwRSV/HvI3c6iChXD9vl0GkJq+Pdl
ce2C+dRyMaHQa7uBvqi0se3vLuWFm8iXLRHJPzQpNW1y2EMrktdvgXRX3S9CKr+0
/iz3mxUM2j6ALXVPXn4uptKhmN5p5Bz9W0oslQAPjCKxAArQd1s1A7WDleQ11db7
B/wBgnnOZMshUKWDlfyNEyE9B2sCiHvQEa6yBDq0ff6jimbYgfmlnlXTaPjc/BSs
LEdg83Kb1lhy5YXETSJWEkEFCTTFSZBeAbRDQqmxZ1AiXJlS1WN7ppco/UeEMXZa
ZgPK4V2c9IZ+tMn0AO9sJQ0keXXkmB3xDSLsT57dn1osJyUZtPsmRJn4UXtN1gss
fmqFDBantbSWxUOGCqXd4oRVdcTmm4RbdFVveFTdwBc6JLOeHVEx8HxwzrV1UyFb
tK9PW72ohbvL5DSxkxcUg/2dOxaFoVZxtyw3w6VkghlrT1bMVxTu40FMVGgcGJhd
EMnK53qb/a1+jITAqdTPpVcX5xgSq7eEb/IiGYX85dQgEKKuI7OPyRY8mqHOt0vu
iTikzUlo3Bw9T50a/H2Cao3UPNNO1Lbe11svQWrjJxI2iqMEn29HAJUeGX9YFNZl
o+OhP0kR5I7+uHBkmiSCEEtb2xigRMDV2yxsp+M8gjI0a80fLacRB2gbZfUi2Z85
nj6wpavEF84A5C19lCcZ3fHDCG63AWbPKcKwnjqAPKIJVLrqEnqcCw/RR77lnVaa
EcWKYmTeuVFgb/R50GR7jXrbli8LjxJH8ZuguWuPkyziGL9gglXXygYNo986N3/L
RBhoCzjQicdJCL2j5Ov2SUnokujwQ0VyrVD6CCm+6M4HqegYWM32gHgooyJWqcxV
q7uSDU1uXTu72duPBLk+Wq3ecPjo5osMmz/Kje7KlMKfDiFj6seL901MkaxMdht4
HkKceZhaiT3Fqz1LEjtT3o6crPqJ6bTxIuOh+FUFNyHRkopppvewwG3MuZCSwOIB
Dij3XVU5abALeZ/86tnk2Y/D98ZhqDW4uQMbMY/ZXXx3Kn6ffeIVi74stGK0KlwV
4uqH/Ch1PBxoYggVYrhDUtFqTWI6o6rLSpShnBWQphWg2lWFxzmY85e0wePQYwRY
NykRqHhBKg0s188hZsBG8pfbFq5C4jnEXsRe3m1RTg2HlR/MUH33GxhjAYE+j1S2
ska+++fw7tLk7DuhnhkuLA6PC12UzEBSNuFFRc7h+F4q9dK2vs6Bj6zYBrfsPYRG
fYn5ckqsKH3/0eUbMUmBtSBKUCnJ9k+Z+hm7+SedNSy37SWzooMyScwx1/7cw1nl
gsJKggiaQy4860S5JBadpRZoBhTm/0AXVcxb4hFgIYGtUj1uaugfal/m3RrP6Aur
4CRQG/VeFvTjkh05BgC1Ry9sb9EneH/z115aInf4Zwhg8WGqwu6ymq8TUhCHiOET
zyFi9j/8+nvqpn/y30uzj5AHS0CyOra3f5iGB+feEWx5C0FoIoIDevrqx1/YjdxV
XC2DzC7xc+tzIxtIz/F5y25DiFcMem9n2OjUazjrcjh/tNUfKL9P8ra0bIpcV38w
+Unp2/M2ZEWJDBWedcqEHJnhP7lyJKH5T+MhB64w5cDYkO1Xv4MYqyA9oJ842d0U
EjpMzNZ4HmR5oYx5UwDVp7EVFzhfa7qQVgNLrCVaAKPF9eKnlzieFxynC4RJkXg0
nxD3+GT676uuY7Xucj0hpUNR1L16q9MnycRZa6pUYduWCLoJua37iVPTs3k8rBEu
KcBE0lm+lu1hXCQfJOvWhwdbCvxcD5eQZhFf1V+85+9xtyfY72DCJFyX83ofXOqC
+zf1jvStappKFI3VyycrYcvBwDZNsKO55P2AJKCqybgoP52h/y/S8N9uOlQxdqrd
5zUhklLRqTfTy84V2x33WdaEIJlpQG+EMNNxZKiNhiSeZK+XnXcodSdHbbG6MQDm
kP8L4pYdy155cuZTEqJ+NJAZnYaa9B6Azr8Zd45mJjo+rBuX7zxWMF8gUWB/Jrwf
hD8Wec9sijZLRmeL7JEVuS1720tMyZT51xMmdbXV2S5VYIr02uf6b2FeYLUVCQiL
6hogaVOiCV27v5f97moC1xFDbYmgNHRgwkOAEa6zmQcvHa2fGe/JFSJrakL7eHUl
7Hct9cCIUWHTZUDKvLiMJ2Pql2wqBpeGE0akAjBWZVldnOfMM6zjgFCGQV3NIQG4
ZuI/YtNAGOmOCdlCBmM4dmvItuNHFlPBt80mDnmLrg56nhOeFX3LZRtopHM8ocQj
Nk+NEF+siMunneHMdEnO9+8XbbKWPm1XAj2MS4g/3lfpiiTR1ho2b+Gzrx2ogtuO
jVDp5uU+rPn6I8Fu4cBOiV5E7PdoRCb3g91j0z1jmp535bZQXprzFsbw3mynyrOG
SHH7zy9y+K+54A2Us4bjRz7xlPboKv+XAvI2A0dEPkxcIxQnFpzVEyGuo6XSXuvz
vLNBQ1J4qFUHlxpxGPYi1Rn5z8DwNOo2zmp0uE98IZsPiPc2qrEOSTXXm/mSPpbM
t6cYDCCaBM9kXKb1DG/LkS58Gov0R6QlDQv09kc/tMoMFwGwCfaTPFpoBrMONSCu
qzVs6OrgwXODUlDAwohjCKUQ6FtZerATnb5pRKUfsiWB/+IMTfKDGq4qZGT0uUuy
/jq9fUVdOLj77+TtfbI6Xl0mlCgGzaErx5bSDt/iFacMqwvEtVCRgb7Ie02GQFkY
bNrQrPKoBcSOe+RZ4aayYMfhluKsFulK0InJJrCz4wyJJBNqFoyFBddo0hClPQ/Y
JoxOScT0pzakF85NVZvthig9IZooOTUu3qZjYO1as8/CKO6DBWPqsz9gBMf4X425
K6qyKEiZNgrHnCxrHyt632HuQyfBFz1cO3Kk0Kf/7mJ1jJSQ0SxC4j1i+QOJM4OV
U3gmAyASMRX5K2uIxUJp9Mm5MZfryV4FGa/iqdMiTFmgOzwo5R2PmkUQm0ST1Sxa
nmzX9AYP3VodyBf+eGGnYCC/c3bGe3cI7S/W4e9Qd9LEyu6zBlCRuVe5cL5p4XKE
SoqV5ljY6IC5DTPGN/HfaDKagB9hv60JdIYXy0o0SX7Yu8Wu+diohsE35RKBf01D
ptcgAR+OzEI/qDq75Qh/EtCU6zQy3a/bZT+cKwSmcDBDThM8+sJrMhL/RZPj//6b
sD0Tyvf1kSC5UltswSo/kTjDSGDtvF7EvsnipamRaCUWn3CpTZhbgpCLStF2n5y9
ZYEWAkeH5w1TqUzkyqn6PGGgQ1fY++KwmYRJ0PKpd7JpZURcAqWCQKo5/D4PEl65
sLMs3Kv0Ho6uiwlT3kLQJiRQMZNB/CJ8WacDshRnF5VgJ7Y1Drn6KKFdkqI0JaSq
M3OH/m6/QWhFQ0TLFiSHFN+tD6dKgYokbF0Rga5y6BqZBRq0me+qFh4SkxFImfQu
J895ikoKOlMDo1QSOukYPUcfCmt6XOwQ0vkBgxaUkdpOhIp25B6FPlGF/7Wqs9Uz
0kfi8m/AQ5aT2s1MwZVI32S0dLJecFG7n/nrsE92/96TK1zoF+Z7U0WJpSTuNP2Y
JvrSI7GcE/ZYreIOXmjZNh/3bTyXPsxqtPWOWwEtHXSBh/+uyyHzWeNaZIc+d3ik
PTEWj+Ms2kqQXyPyzAYKpWblBQM0BvDA8rByXddFJJfDYD6pEKM+1LAl9scQOdA6
4Zi/aJhwmcavlZrf9UPyetR+CH7LbMn67AS0h2u4LJaYaMn92xuQhK4cEVFOVT3F
xZWbE9UthWsg/dOFRIIH/nwknCqAdIdXwgQP8cz/58ayvSgCxAa8QUQ6u2+9p1Xm
jPy1xYsJIq9eVC+EXaTAYE/ZGtyn8h5FQj2+MoYuX87rddUO87MFJNv44wCwnpah
y6ROk0/ok6YGzk6eQO+U4mCpa6nqDnE7XEKzecxCI/WNK6dbsZXAlOgy65nb+l3G
pBSdWZ2eCvxkAmDdANI/5kOMJ0bDOdbnsNd6fjXqbtEHwTI8sganMpMQ7ht4Xz7g
12vGq6oG37TgqM0ofczvIdg88nX9v/g/3NcQKFV5I1goXALZZzMcPfOm21AtxZ76
hmMRcjizfoODX/aqTGjPDDxCmB3eGVqup0kOBAB9OArqK15gxbaw5PBqzoCaf7oz
j+4m4L5K5fnmODcRu7p06aOV5GFnC6CyHQOLFrFAUZMScY0eDs1TddVFR0QxRV7x
hnxX8ZV8gMQ09ufsi+3P6cvdu7teGv9dNyxCLlNyNcbyLMB13FTaZxHho7raFFHi
hhOdRmQe+ChctDU1MnX654Aas9+rVFyd4TDiyOoVB7jgB/Y1DlHQgIWcGfYcAgfm
MgboVzGD/3zIjrd8b3QSkrGAGOsNXsIyb6Grqg2ZWQxmFnCJ6JP0SDYtxp7XdwW+
jnhcW4yG0GVOPgEozXL/Of/uXkdmPuYV0uiboBi/ZTH2rrrOo0ITjKPTWKHCnnud
IzXI3QLJIfS2+vOwVf2xoPVw80k8pMnAw7rmC74M/gmCgNCoaHCK6h1r3ioDZfvB
cL+nHyLt1sM3MW2tScqVTVlWmzRTKA7codT0UHXVmGSxKZFR6WGFvNGJVXF4XmOf
ekvNSIIJMXmWQCQxTJED2y6VjLJ0q73KcmuEqLCN+7jmpCc+bxe8zwQNcVesxWqp
WWO4Sb9xbPWM6slX0iZwsQHSSd4W5CeGqfRnVxOX5abVd/2t6hCFHJhrEVKo3SIz
TASIAgKrKDAa/7w5sB3Qo3xG0UXS0YwCQpjMkQFObqgEw874THRHWGDHQBK3r/96
peMbfX5sP8e6lLQ3AMjhmdTPVxbuMoa3wEz9PZjDmCyiCjsv9M9ljpvxMpcUIvOs
QCGO0FVhxWRyJsuVcjVl+POEL+QVrBuT0Lv/G3Lqn/4oLNukEUJ+l76iRJYNlXVX
bAqoIptfrz1f99ApNdETPAD2VBKIRCf2t4r01k1o3Q1ShQ5iwu67txnMWJEsCm+g
6Dam6qBCQzBC25YZYKQu/ECia/kRn68Pyj7PaU0Bp0/37a4pBNtD0qU1qHJB0jP0
45rR52drGx/lkiiPFRLHPjXIS1DZSi+V3dk+5b7cHe6VEVz+Pe00G34qaAa8pJQV
WqtBi0FlaHw9qZMupYdqE5I2eB25UQBCZgrWAXCH1th0R2Rx+ThTJgwhgj27PBp7
b2AsQ7G4qL4O1HYSEQpIOKQsqWwAURVZTozElXA0MROamUSFWVU5oTYtR+iDDTrc
LAVEkGLRAqyLBQLpwVl6jEjC9k3xvJDI6B+7gXR8fz8IjJzoxooRzOVRTYbXRsXP
Cvd09SOenQy/kVYE8wdd1ONigv8D32b0yjAAFZ+3skyVAXURTXS+2el84q0kqVkE
uugJrtiZ6fsDmPSSh8M9DO+pwStw2Fk+pCdSRVTc3PtwnxNJNIzQWq7FwBRaJD32
VexS2nzdcWdKZFRrxcWkA+1dSUWffCOJiU6TqHedeYOME7CIUdFRN7fDc1o1w+E0
nWbLHN5BM6Y4J+PQnggNG+62q88/Ptfeh+dDAmrvr5C+SeKc9/IFWtAjDyN4Gbb9
949D+zGqNuhVWvSFE7d+k16x7wqXdv7t/Xx5yjZlb615NhFitBBWAf9jZuUYqZIv
jqERBwprUTyNlDSZCavKNOj84AWNm2pnBJSGbRK9bPigjlCpeFsR0myU/ZsVZnW+
DQPneTHvHqmFS1h4gyYfP1f+ar7rlwmF81Wx9pdAqOmfok2J6kfW3OkL5ooFXkNX
j4JObptMClYsLlGwUpLqKXnHsoPXigcLa4HZd5Eu8CyBfl3wCuZNBREuWkn/qCj9
YFLXWkrzvvyK10vJyHjHBkT0F94VqvRsJLPnlV77Y+LsCq3qvTbnfqZN6MrJ0VrB
xDdPyNkuZc7AQkwZiWWztflmID5eo5aZsqEQtirt/Vffx6Je4O4LGHTMoY9kMFkZ
qdp3yQYiBWj8P/VZNUPa4KS0RFd34CNCFiKOYF63N0iZ1IBIvLI62/EvnWSoTa+U
i9zSiFHkFhYkmR4Eg56dUy+cQOcYiuludPjzOndQ+lFMB7ccRmDFPkl5clDDeeo+
iTEHlzF5nhMtYvkOVSNgPX1obv7ztyq5G+nOezZIFbET+PnZnB4ZNOqxCe9HvSXJ
QRUIrbj63tORMMpcSW5hLFy3RPj1jtxuSB7v7zkf9Of/kUjQCzpdD7ng5m0eUXxy
aJaT79PGwb3k5qiwH2KHbIqQEDj8lqVYe2isbceEOSeIdhY1KtoEx5U4IYSldPRF
Psvi68rCQ/NIQFLMvUiYQuNKN3GFhaUrN+MAet9rlWaJyl2yPG4PvMoy4GSlWGNY
pFSotJ1W+/JV9kel9Jr71omdqZCFv1JYw5JEzgJpKh2Od4ICZPBxly0rUBjLxOkX
nCvpUqVrFzQ6OUvVq05DFAPBFnyxT/qFahKc1ncFwGSuimDqF0N/YDkRuAJWGdtR
J/39feSm/qpmYIKNTv7Es9Lo1+Ic0iCg8CALr90GAcCp0FBtjXaQB2CR0GnlUT1I
iDfXQrV7nYkRVXW54G57b3F+UbxEZ5pq7aS8+Afr36QQrDa3KQ/rfwLQ+4NDpqsn
Ywjsq6hV8Bz2gb909m5Nf7x+DXW9DC1yp+uvvFMNL2pjvLtNNN7OFjkKr/8GVzkO
/3IJ37feCXlxhBqmuxxoNgj6GCWHc+who91Bj6z0PiBo6NAU4qSwi6fLAepDvI+u
NJbmO1IdlxosNY741B+x+6ObEGkJSr8sKM2wUqSPz1cdZ8BlmGLlzitKXisd8AgI
owkt5+SP9F+EXG0W8EelqKoEcuturnINOWfFvVix6nuVosTuLqZzk/LjZlR2XEuR
FenV16WH0GyQnvKNbV3TbXgGyrzUF8ipfaMXU/C3bEpKKGetHKAJsyGV0Dac7kMW
pHemfbhujYXPQP+h8wl/oveedhqa28PnwhZHj5Upr2GOkZ2ccnZV7IArm722ahvk
BsdDEZZVpR1sNMAa6avjbGgK9PD2hnLphaExl+W6sbJH7ryEseUlvHn2rnWkdyQi
0DB+XBn2XZRzJXXvEt0dZzcNhZcQyBuOZmNzufm/Unh3K53qhUnvXSmJMcwYiMM5
xhjF1v1adn17uaiUUkQiKdOx//9S3KDr6c3xtU/3QcZmTVFeKCU9V26HKhnNR/qc
/H7MwXxdyfg4YazHVYxZvi8+HzNlz/tBXsBc1Atod5eoaaRSm5YiYObviu0dJCEC
W4TgduAq66tjaNTvjYpbkCilzwNZX3ciVVAtFDxaQG3/bdG2TeZR3uQlGbW3a9sh
KFnri+5kxcwZyVPpfdYiC2ij6Szd3XjV9RJaFkm8s9O3Inkn/Fbnae8iQZJBvvHl
7sWV294KLX4jv5ZTqiVxHNlL3fEYd4GFHcCZaSA5q0Kfkqw4hNUcS+3zSoSULolv
hLFy7hnL6+c5nhiFrvrENLCK27P29/GMT7mUVasYED0biO98Wxu7RD7zAUFclrhN
9KsNpNirapB/yuNkthP1GCvJxedzRFUCvxeSxF1+6vB3qbxqHAtO7hUoW+987maK
m08F4o5uRkjhzRmL++0sgon3+Tmgl2jS2GvA35jHDeDZl/qHAi+WGEqLf9tCxkdQ
0YlQWo8iaWRf4bon1tW6UIHwwgMftkDVGhX6zBoxmC396zdg7IhkcWpHs7pR1XaC
i9cnDCWRzY1WB6m4u6sLhGICC/f/J2typd4v7seF7glY94+CyRGTfGoVBFtef1GW
sRiSVOcLg4aKzu9J+yNhm7uzm1boQW0q5TEdwaiB8WU18k20JYJ/OMVJ85AWKMPf
R2bI3RryIK/eNBxHosZO4oku/L8jAH7BILNi3b4NodILXsw9VdUXLlgWRc9MClgo
t/gDS9F+Hm057TBqD7BvWBKWB2ZctqignMBWZ5hcqzoheRA1/lMJCjS72vsuejlS
dEFf1URLumfOtbeepcvOfm6LxUYHlMUBUEYKQVub1TmFbtQCAMPQ23xuEgcwAYju
A/IqsBw/rcve6sHbMChrqfaaVbsBHc9FzpFMhUWYTQFVACaKuEY+Jhpe7N0HPcTS
MJ1xl0uc3AsyY2Cb4fS78DO4pCRTuI50JTJNeCUcti1ctfmuiPek+tD5WMLm4vTY
9b0u7uHd6x4fe8sNBEf+Mv/c/dUY//cDvlR0c8vP5vcqfgskj69ZMqrggASbdJnU
IYWtxuQ9TM+YwwVj/DctmoDKENn+/YTpkCLi6lJtzwN9JYMlABA0UXAeYTXurrSg
OUZxTVBGxLm6qfxKKjrFQMuXhSqCFkpehThfqnC6FbHR2G/SrW7wezqz55GuNYsQ
UQAf19YRwtPvPuBlD7DVzXBWqJP2mabSPbj3iOXF4lHB3g7HWloDzWR5n+NSTife
UJ65O1tzAZGQbRQAsozsfoW+IX3MlZJbHzNYaed+gZsxBAIwud05IaVws1v+UH3v
jYmgBWH/SjIsV9NOkgyFlosAOpoJUz7ZtWINSuZaYnnW51v41jxlgVW+jpouPwbg
HPCqG51j0QPPRS0RLwQuTdTqYx6VRnGI92FGqHsp39BRnClW+EyCHPbWVx3M7R3z
MIzyRGDbvGG4MUl3neMFtJVd40fFdZmZOxrp/iXoiwZt+TjV48WrP7n0Cf0eg2pv
I0XAgerAdosHv4McQneq+ZoKKFIp1SEKgKA4qq+jjQ4n15xE2048+TSwraBoM0qD
Qct2wc8VSpj/kGyHn9AII/0Al9C9LDizZKA0PiDk7xZ5VXvrP6gDGcQhQcJce8XR
+Pg7d8S/szr/OHJFYhOX64IwvlrqGeFcDZZES7efHn+VhWFE+yyWTOnyW7fCdTDE
TzVgWl5YSMEI5uF4RYuZqmAYakD34WyvAgjSZJv7iteHvMcx/2fLaAAtmAuNvaDA
qLL+xri3RRrG1qgtvylS4gseyAyAzlSPa1B5iZUAHCoHTAC5JEgdzQD/nm6Gyalx
2TeLcWDGIVJk+SkMf3X34Ga3ThQOOh9/j4iWzdtX+GhLkTu1oQn/ACJVK9nPzCT8
r/mOXFSbfuBVQ2Z4NUnlBKeHo7uIOKVCDwMteNya4hkicOUXoqE0m4tHUTrjNGYR
A3VCj/xAgszy91pazmwACDP3SWYyNKvYXZ/vI7sayrzYlXqwiJWmPvke6kr/5b9j
7SbmiWIx9lAsBSgpOC6MAlr6KsfL+LQSTZD+5tSstkhp5wBKfbsrJPl1oH+DeAXW
3VB7Z5t3KdaWoWRuKmRmq9MYXgb9qfx0S8sG3jdEcHOwyTiVPdP+aY1QscycBt5w
TUTqLGMZLxe48/RFNoCauNPjbyJOOm7GzlHSQNsleRcY3g4Gzm17mamWE4UvqfDD
vFWQqPwKC8o7u84yyRjWbKd036S9XoJbBHnVc9oz+g1ewCh0jbGT91CjqRl9TxPS
FAnLAh8OgLwfL9LjRzioXmIMYaB8kcIeI38NZ+usiJnUgSEWh4PEtZCbZhYgKKpq
UwXYTZQFDbiSPKk4Ieju0vD12nnTbetu7zVx6MkXOCLiLNPYnODDN4s8GmNeW3Ya
+NpOIbDk837f7cdUIVufFnxdDSjDugEWzYfah8SCjVSBTPmxzOujW5eA+oIS/lul
HHuzaJXs0XUnYLefY46xjbDg97EC9pcQ6JhPRV+0PrdH9rpFBegBQPq5XTMPfb9u
29eGR5GywV2dZSQWxJ9FXglsj6Yuanyj8NsGeH4Gw2G5oTq+BXXFVrN7LqbkbnmI
lnznok6gSTK7ar5jepLe7xbkCifKd/nfYiCJPVZqjxHS+ghkm0mrLTvt//QHp3dP
ZHfiJBu6gAGQar+syWxthFqpevtDzO71ikCe8oCscDcoTFUIUfSWrjZNM5YFwBJf
0WAkcIVjATxzTTdeSkQ2hd1+VXdJmvWB1A0j/LQ0slFAslR1dlpoUgn7e8DLZg1n
/CyRds+KacoNGbvbnnzyxZVEQWCQOtxZb43rhTWZSiY2vULFx2e/faW0pLMzbe86
I4IXk2p2onnVeSEVOnM9O66YLRTznb3htPgOXShCtyGpVd4qkPlHl2f227Fsehli
1MxVcqo45dQwygQBZAp2ErmToIkP52IRpc56ozSeaAkFhQGp990bhHarnXd2noGx
DULcCWzChVXucKG8HbhMqys9KXSL77YkPBM1RZ/aEqKdvcC+lA5ZvbGguJQwKp2L
+s/N2x4jdfsjbI1e+fV1jaJVUqFYWMhoGufmGShvWUrKh9RuNFyLTNZDMB2li9gh
TEil/oRRs5sbVI/3/wycYSW+WQn0sEkBUkV8hxLiIqWrcifY6oLgGgHJXVeM10ey
HyWul1cfXFXa5EekoL+/YsdNdeVdTpJoIg/Vz/EYIh+QFcFGf0UONTsgSyusC13r
dUXICryors9CrivGFI2RScXxvdLHG+X14kLVHfdN2VlhrqYT5xhJN7sutwbuZbel
/rjjGxnem0asJj4YuJcEvA0oIIdkhJD0a2wMep2CybJRSwJPYQ3970YFHBphyDk/
Q2f6M+UtmmFQ4Toh13VuUTBiuoCl5ALHUpvKWlTi2KXp9aYwa8nanbnC5w1Ffetk
8sjHidjAAzINBpNLCNB8DgITw2jycOxvFtythc7SKnFbXPDXYCyJjL1o+IKX6tHb
CnaFVUheBfpAhKNVDualhpJJ3seXG3UfB9Fg8GpHyXz9f1+e0cE49El/HtuFBsXa
0okarhyWf/cl7vAmrhBPFgzr9GVSxNNzOPUCmJLfUiTa7LPWmr7100RKKspfG52N
cqI9DMbCCsIp49rB9G1qCvPmKChbHOjzuwpyzs+4YggCe9dkXLwMpUGAyU3kgXbF
6S1RKUz2RMvwZik7tA1z46U6XxICDP9LuZAOsTqXf5mJcjTku+WStnMBAXNbWBqF
HNy/1vzjX6ZTW0jT5i3BR6ThjujYvASgk+gTOiK5tDkEf48HdrkC1gqQAWqKYL0j
zQUubI8RYeNLzkakEXj8op4OsehSwL/3DbTLhpvM7PsHfmoc++sZTNUpqzNzcssM
mm7s2fwbS9ghatuf5FMsTbx8/OUEmqOOy6sxb9CmeKEH5VZlZti6mMh2ReuhSkzX
QeWpwtc0L8ZMDdovsZqkin+GZGwAeYavyjwp5Sk0GyMhY8RS4yBZnIbuMnqNUG3H
pprcuxWmZZ2G3frXp+KEbWa7amScpq5Y8qFq2I6Ir+SZzlq+AsiwW/UO9WHdS5kH
CfNgyBeTruJtfokN19II1ucFW1v5STWkRE0aE9FDF4g2QLJtokBLfKqy6GSqVu+m
gyfpHE0+ttRqwXLsJmz4nj3a+0+T3+EcExlO+7OCeuDXDgl+vJ8lT2nI6TQ9kF3y
3xqc0Pa3+z9Ca9cG6y4eVquTEXiViYY+BBdzCz7mgAKjKLpM67bwhSw2JkO+7P99
Q5EEji+jxzYIQeFXt2GrghMRZ2TVPiZeVkNIRTeKrhXkEj84Cj8hUi+sDTo15gI/
QxhfDimfM/ur7MsihyPUdrHz/hwiZ4U1c4RCuVZnXosfU6zlZUxdaEtZDgsCg802
gUbR/aG27oC+18gKZ9kn2WyZExwRr4BBeN2ldS8tmoXFSc6Wlsq8NJsEc0hnENhI
FANtx7FiRy5+Z6+Yijw/JTlL4tApRSWdStZ1oJq4swuZEGVhXaTVxe75nEXIyLfM
pYzTsKEx1DH/Qi4hXykdMh+YOzgxgu/JcnJ8GDFZdG3eztGVz82a2EXcbvoMYD4m
eHG8gL4PT24KzPNha9LLd8hZKjsYLwZwHq3/z9FhOhf4ZEtbx3OnK6qfG52bQVlV
prKLPUPkNMLbLunfB2JEwg+jc7nR1Jmmx+N4yooWNdClq9DHSwmaHPOcvfJzLeEE
x9DLOjHgVujBFF7S1xqbwhBXN1jxlUopO6ZML6EU084kD+ldVDCeg8z7h+dloNrU
GcR9/wKXU+l3gsLI5RwEE+4JqBFKDNZBoerWhpI2FgbmT/8mnvMZcUfN/bhO5tta
X4T+IVl9uBhZgZaAD8MIRhzmIqUNJvI51o4qI9nu54ifJjdGmta2XMrS7FQzyU8i
F/vj1Cfw7r2g6wbI0ijJVGk6/chTJwaSmMcpwOPWpa+20G1Jz/TXljB4McYslZaM
rndqKP1Eb+SHIsSiwAJtgfI+DTXwdC3YD1IY+YuFf6mnFrI85vVYiwghuQ9lrnvk
U0aQpLjEyD47HzPsvA3Rk30BOtVuOBdrElv7GJNN4xrXhN7d2euw/p3jH5n5tfmh
zbxsyhaEpHKTC2tvSOkHZDGqZC/CuPoYxEsgr1lwt1lfwzH9N/RnhRBP3EW7hADJ
Re+d6Sl6Rw9ST+B1QRtVBB0vy8iuV6aJIfl+pZLGRjHIe/FZwyYXbFLLviUI5BxC
F+sd/x4KgfoyhDuQ+bF22q3QaDc/4zwTOIyMGxbX7k4Td1+f/9KqPCNEZFLZD4pI
qshuiRqJb3eqF3jwPIiTIL3b3iVkTTgB11Tesip5D3KiFftVAcq08LF0KJUVZBBr
1BgnXLb7DRjC7Lq4nQ1AD1HQ6ypFEwpMKendk5MJnCxmM8O0DpBfRo8oLzNv0+FS
O+Qg7bv/7KTADvpZ3i6ozZ0sjfe7BupB7L87bbziLwjG8lIhZ0cBH3MrmQm9iBpF
+aJb1aVgQf7NKkVAQuhyQttLRNqN9ZaHZUoGRJDowDUHWhuytVuu10uKLjFS+7n8
3LI/9dgMj5V427H8iHXL8Iu1Bh6JRctX5sHSpjIaJdMapcenFAm4e+/MW9rY7RKf
ZWsSUs1q+uE16kntfqzI4a2humFSK5bdsLtbOiMJ9K+T2RLx+Pxtrm54D0klqzr+
SuH0ZXQwBm13S9z15Bhvv4zu/2FJDH0qPI4B51ypzGOcGYv8CWINvVz9DX/waHJw
T50XRmVwX06TNTt0kV97oPhFCHKoAeHEOPgP2rYSbqruuWk/qlzzqSn13Fu+uOfd
nCrShs71WF+hitd/KDQ77/L0XVpD7WxXfWTFxpWoKmWcKviivjyU8dPW+XZZwg04
dH9QQITF/EvMY3gMoTrkFgHyCeUGM+iUDzFVOWDpmbYuBFc3WJRyrlx4ecwPfdqy
vnI2NhjA9RYA9AOx6huviu6p9BdzM0UvFzzGB8dYKcGtxUVW/k3teoMVyHBRL906
oDz8usHXvJI+iCT714k5lcQiKqB9hsTzLZicpMpV0HYuFQiIOlmRtwyqd5ZwUb0+
k+7kS4EvH/YtCiwdYcMe84FSO1wCzVla+N/2FSIn0zSC9Pe0taTfZYm1uaBhSP2J
+Jc4/r1SfYiW1h3CysGz2Mr6WlMSeGH+WEDp9weCBMew7XmlDiruZTV0iNBe2DO0
FLk26Qf9u4l/jf1RbWIfe78QOJQsxXUumJGtNcFrcZy/n+5oKJLYELJjX/9yyMyp
3lSBcA301ARUf8gcQvNnRhSPVBDZLV3dBSYlQvfxkFtdZIMy6hD68SMEhK26BMRZ
2a2Pz6Eetq5FSLgJ177EWR4AyV09zFeY28s4dRyD+GIisAjFNV1gtzii2CIfFLU9
bBjk2I9wZRixea0NSAaWl/6YzH6EWQr/VEUUPs3XhSkoq4AbFfZ75nMPab2dJkv6
/f7IrI/2Qygw38AkhT2Pojtnre6TtLVuZiJQKjfOjIBFF4/pMJXyIxmVXE0LDbgo
ZhmD8e1v+bSmOTsEbcxYOp76INwbi3SU/Mt/UNMP/UemVnOSqnAx12Hlw4veErzS
1DflhOQ8n7iKjb/ROf+wtIavoQucZnUhujAWxXYAmtAbVBZHXhh9a39rbFWo3gh0
SUpKVD/5WsiV8EYhoOeaJl28aeuzAisT4ln7H/X1bzMoocvghnnMdMk4i702ZLnd
5/PfrBRGMAduXJBB7JOIOqg3mqxJHLvHYeRZ1KZVSTXGhGZtPvHxQIUfh0LruDRn
+hKpjbABQXVlgBi8wvToN0eOv7HusXerHZ/K4b6TOsSqgLmA5QZH4ZV6Heh11py5
z1k/ICiBRXlHexyiz8rw9pkcAzr4JiZS0OWBjp+9rgyjW490sqSCTQxnGQEME/sT
uGYpOrpVQrdvMzPe5naSC7wtb1zBs9CJyPtli0NRbWuOZBXDUOUtj0qk3HYfyOmK
grDi5vOGJFVV5Q0MlQC/onxdaJFAfHinZusLJz1m3x2PwRUT/Frms/jII1p0nz3S
AaUlbR4SjvvUobk4z4ReKWgqLv6TJLXl1UawEPVj3j7jhF/6AmsgU270cwLlE4Wl
KnHb6ChZ6vUF3qQpeI+HMDb15v3f9/AHuf7GmySwhv/c/akMjzPngJP4kuVqJjj6
Tt85/a3gkuluE8jntSEy6Sda5RBKkuXlY9yFzVAaFlcITOENqKC18gMcwvk21hV6
35bSxK9Ig9Bantv4VZnHZnfQp2zxBMnLlYTjlNEmdXdKWBiaGJZWYbeqeeUiR9L0
lBfR7I9EcQ9FZWpIA+5o6nnnxAllhuM+8GnK8b2uawhNN4m12tKcoU/LJG9LZcQM
9IRqdVtjHci55CuxaFiOHbt4hdAsZE1RTqOwlfWL4AKZxU7GhzWMWLmtjU+iSQnp
vkR6RnIp8I7kLJSTuOwW625ki6U02ov39CjDpjplzmgDduGIHKWfEeb4KS1WiD6k
PwyuTAnqYdz9dJEzO8gF9az2hUyiePuPczWyzKqxMPk5/4oYFeKjmgMk56WBTLDr
OyVzj04PiwUqp+IPpSHuGY4Sgw6j0Fb/YV+ue8tW4Y+l6WKT1n/NZ1Q+37wPvmfj
FDvYu7K1Yv7AXG21xHeODuv8DKTf5rBYYMfj0gQPLWFTTqPeeohychUo6XtGCqz9
Mhxsnl1t3qDibUnY4uJpUVCt8VFJAAgymO2tG8fHfqxGeGXdjbpB4VS89JrKOPU4
kEJx/AL9LzbeK3Cr17cCIyK/30eDtqx7XxplS9QcQADlSqKXyrsDQvrDhYhOPBg0
51Y6wm/1GD2CF9MNnxzP6R4UHKdN/gopD5/9JOX9cY6SNZKz3GP8k1BsA4U9JQkv
Mc4AVhhyzPE4CLZ0AN/eQ5FCwURAlw4pt7wQA3ZB4QCfSydZsclarY019W40IdUM
8aBrWjJdmyuWwnSm03xeg5LibbIY8p2XhcTM1YQz2E+/NIc5SPP+O5Tnrlv7bxWG
fS95j9G7f1zbbohsz52o3ME0cQpnY2a3DyryRYQcr12WHiDSCVqr+YLOpYBOmc9U
kKmM9CgoX1V8ZCakUkqOblGLlvUA5MvqatCwDFl/N6XmkyJbz4u90ODgFk0jXKI2
La7slik136wZE+jpqgGgxMWeAWFpEs17gFVehffaoRdBuUqi2AD9uPuJftQ/bGWh
iPS/9HR9v7ElCDV2NJeSYuIwMfMntPjTipww78hU6SREBQydhDWUeXOsYZNVEl+5
O2L0iMD17DSk++njnhXrE0/pJGmMvLLsHc8d+8Cq5w9k2SAQ3U0sLZFMs3/lIV42
puPkdqVCAyQ0zu8W6hK7I5u3Qy1G0DQtoe+P/ssvavE6d++zW6zAeBjkCzBa3Uwk
HCUBjOzW3hNkz37DvRxjq7mAsdGhOg94YsD29cdp/h4nRCKW19bDM5TmXW4uoTAg
8hmSX4bN2dpCdiHbEVAmEWmnwtZaatu2Sn7Sl5Z5H5MvY9pUCEBWvlheNlij0nJg
d0rGm6l7fBnodCsMv3xI2BlWTS7zPu+DKCkuX7Bw0mrlvYypY5yUZ+XiASVuOSsn
Mfu7tkSVT7GeWDsj5NqWC2pzXW/OgN3tNV798cpakB2hCg/xx699r6zKlqfh1gWX
FKVk1fRq0sa0e06+Wsy/6yenGbie5gELozOBywDOBROAppLt+ux4WrTUdYjjKbLC
D+s65cT5VJ9ZWCWUGCv0r6Inb5VGTjaQbAv2Gyz7ngNAfuB01BIrPeZxgOVbPb5/
KSX6g8uS4CwzTHXR3Ud4Dr7vAfNsvkpDwk0keLKkIpwz+1OuXfwxfBT9djQinF4I
VLigw2g5VLVA0pkwCL8tMc4tcnbssPS976hBRmR7uyHz0IX5QAxa27oMxt5147tl
YY0fXix1+aOWQj109tgXSi38MJf2iY4AbbKjwk6x8kYXz+BNEiSiONydvpDGMaW+
weuRZ4Kya/KU21WLlzWtYlqemoRGGYYbI214DRo/8oHhgfRuL5Y87e6r1sIZzC+f
I07fkgiccQ/DbCipLcyFPVpWshETN/I1LngSPuXpBoe6aBfhMwUiiY+bDMEJhixG
mETzkf9gV9YhfZ6HKe4oNrrr2IV/VsPdO1ppR+wClydpwVYzKy+VpChFHh614cmn
N/y4YR2u6DqvqXR6K9L0dJF1s33JM4X9kPyW8QFl0MmdFU5Prok1tgwx+vf5cSvY
sUQvTOvQJgdh61XSllEHsEKeAojrFvI2dGhUkfMMH9qmPXVjpz4RvjyXwEbMrZHM
I09IQ2boYOPx9Q9OF5tn3LqFunKjRD1P206qgLLhY8afg118M+aFhqgp2+Ochv3v
FROZhrrfQ0mBPImocGowKb0JxSNsXEo7NBJbxHwj4uibvjI5Iio7x03Wgn1dt8i5
gXyWnoKUuxf6cLdzPE+AzNWbcljr6juzpR4+iMtO5LesJf4uyJuuzP3Bo6USqI9C
XbgPLbRyCpHiE/ZRp5w9M2kiJOMTmxrw1bR4CJKK8Ej2IPK407gT/Xll0JhPxaBS
I+jDk461wYO/XmBfgY9RBw4SvGxJEz9HmLjG2kOJocGc2svwfUvLuGfUFci31l6y
prlcieMvm923EhtN/0MPV7/7qRdpgmyAxYKWSgaQnKispGNsvwv9YOKpeg4/FDp/
/lF0kkhQ2G/sxBcCw0lHDe/jgShIwikqhUMhfW5aGeJF0Mh9L50kOsHAxkunHSbg
h1Li8Jycw5nOJ50FQ1iQwHdkL3mT1lWJuGTi8s9y881hXtyS1H21pTkZfmUfSvnL
1nyVSJlUdYI5oIhEiXCQzbCYiHntaEbEkTq4QtD6oi+ksz7vO1hBM/Z5jzmOUMI5
O7Wx+zgWyZhtECKd6+pg81tco2m+uPLepQpm+7IVRBxQ10iqIz9PDsyGyG7EOh7M
Lu74jFS+/PuyAZfZXn39SSsjAVAU/vkfMF8eNyu6xFTFGBhmbbDjgZ0LGcUbmgo7
FmgcoOsPDhAReIONwXGnkEG3TEEclansJqewXSoXBBwueMA20Usjf2LyA7s/kz/K
4FedW6U6x34TCEcOf7HelLTIh3f+ZcjImjfqjrZHhHCAnC/ywd/HIKuMz4UY3y53
yNOkfVv0RmginAZONGc5WFrQ2Fayb56sIbGUdIpgmLeyrJ3/61iM9glfCH+sa/+h
B0I/y99H7DnVDjY16AFd/9Rua7w9ZSLbMrTkJYkmz4PDXguh1oL5acfgT8SiskCZ
UNJ59/zrK782n4IgPQYi4bZU+b4S2xkBTUaGW4EVSzTNQV/cz7L1GJSjz5gZPiTM
wQk5thDuAZ7shV0x7Yfn4EDJOJqMqtMsGAa1iB28xaoGic46Cvd6N8LzcA9BqJoK
JowxDvuPfW0zHDV0TH3VYcJmYIr3UhxUssypU9Gy4YhfFC0tENjQDpOR1f/FydPB
Qqe6YLyGAiRaWZEmP1yo24D9Y2rArcOo4ouRS0JnB7Z8nPTDmMxgaQ7WdubB2ETb
Bc0e2BOSpehCUbfAI5PF2mIqxYDdFr3Y5Ry5d8cj9Lmu9ovXJsPs/6xNNXJvhQ3K
dOpjmn4dl53eZta2ebVc1cQ1Xq+eu2/Y78gr0IvzvAFgImzHTukMaCldj8e7iUhz
Mj4PCl50hThccri7cmcbYJ7/py/F2vAZWtTS4huMOHw71YZPJnQTeCSgXYFZUbDW
XHhpzypbgQPGb6kL41n7adZZg1evvZSH5yiJFfeOFP4e4qxODlkDo7gDWOLPFa1I
GIyGgEL1z17LdhMafFLuMSiN/AWgtVeMJO+wxef8zMXd85afenVYNssmI8RMSuUV
VQ4jYa7H64jDbLJjLiLedFTVrpTKF2eOGC7Cm7KmSSaKRWJZCeZwZgq5sZTnBEtp
9Ejuf97g86ysr7STJemVH+gPJSBJrIUFwkfvnv+Gs55GWjR4UA+GDvo+xtno2uJ3
WlH0SzMznlxstOc3f8FX5R1G7XfAOonNxzPCatHDbLeiNTsa9Lj7U8Ohj2X4ybdM
jya9zdIABG68hMKSjHbywUniOMAvgO0M2D6TpasguP99KqW4NkGilGG76E/ihxqk
pyrieMbvkTfOwv5cBgWKlIVOlWmh9pMKcP+8oqm8S5TC8GJO4TIwb7eOW4SYCSm4
IYNWeZbL27D8Vm+yZe4nLH0h0m4Bx8l4qSNbpgF5m/G48fvN67tD4WtFFcAiu1BP
RBMmoHv6LWzLG39B48qMzZONvEZ6eOCOJ5wZ9i6qdj/gpeSU+egSlNlWelETv0lu
PZvqZyy1q33p3XJOXYqDPVy6kgbZTv+zhqONQlMnrEb77s0hgsI8vqKIkKGU+dSJ
LOBI8bjHOLPot4jjiE/5YUKL3EEY0SXs/z5YIptC7VuIczk3uMfnWCRLgmjvrZHB
1gUKjTVuZldtf17mhPWqR6L9rQuQd9+YXPlz2PMt/RE99MDpb9YCusslkeZbTNVy
81P7us3/o3V2OH3Bn3qJQ3Dw9CRevSApwc47qjBj5FfiazPKLQxsnfRmdE+UnZPh
ZtiqMCiHNkdgtO6ofMBPfL1iGJMAEtzfcmlHow4Qp5xWba5HbRR03g/F8lYP2t5T
QJrQCzD+wTPI9+oQ2ib/Kwk6oZKJiiTlRTg1uYnFbpGdORMfddloneYKMBvYzVmy
hNnxKu5HmCfko7BT5f7/dE5Xs0R+3AWz4rHwa9XYEQpAt6OxbdEKMkOuKAyzJAhV
hpVYEsg03ogiBD8Ivz07QTXkPuKTkqvk22P8Kb4ig8CHKQ73i/Z0DzlYD8uaVyER
EDykPnZiCog6od4GB+JJXy6SLxrtOOES5gHyjZkckJrVd1blmIchkRQ+S1DSSbGa
gnisK+AL4qVKKhLrRiwcPFskZjKF+/mWWDwTCJORINhRu84OYPquocsIR867cj93
e7uwn3si4AsFYhV93eugEPgqaXI8mLBTQ98R9n66FE/Je0idJE96AQliqsTTVeg3
gMlAWhOGtCngFFojUUeEerJQn3/foBRuEstdaO4+eOTGpMbGDikGae07kGqWmH9M
ngxFuB0k0xROz4zZ/m6G9poRfsE+41gYfETrQ4wrWoRM8+i1AsNbqLgOX3Z90Wne
vx3ekRwg4at+GwIO3osaFB9ll9IYU1bI4YUME/NH5JAdD0925wGLBSHY4QJ9qojg
fShlzdq3KcfruBnltjoN8n7BokJhbo6TsG9tXZ8IsqhAwNhTOstnunOT1ajfHRZF
BGX/GxLmxdDV4V0SOhi2LkJo6moT19DH3w/3q4QJVP405BehS0DE5T8nSC7JoB4T
aSBhu9VM/kOoDeZUTYKqmypfC0v60g3A84X+VNe/dMhQiprLj/64UmePX7XUa9+k
7mtZDwyS5yHg5knQ823UrprkQ6jvrP9f9EDyio3mAqg+zoeiGcH1Vz3nKkdB5UH/
ru23FfUfWUfrf1XA9eHZPrTejjtuf84ekE6yjNuYRySFofnnF0tom/1DPNvF76t0
F4RhpM4tK/7WkQD6TN17kpHJ1AJ3ltRzvfuP/YJ1CV9W359341Jwm/StFD6aBNit
Rm2dEUNmLyqdOoRVNb99ihXeJXOyOpjXVJpaotnhkVALlLkJWD6GmA5+p1On7V7W
EMHdOXikEwrRfEmOpyk5UHi/aC9aaI7pYBCbJ9uxw/t+pAHnsmlqvhr7PMNuAU+U
WK1KtUEoBEgkxZ54tTLnMJzETimOPNTxOw/t/vPImFBj29EcVimOYTeQWoRzOMc3
6ot4NotmA/WxNYcjV83p0+qTTMOQKjqIf+qWtFK5ouNZugXsCdf96cQ+0Z4BDXq6
hwi4pZGErgpOfcsaUQo1lgs0Q1bnc8GE/2ArdjN3Ch3Q6WE7KjBCy5djDJlr6u8g
faRYa3u+3G3MWp0g2Dsfrc6ebh2/h0ILSeRxpChQT7tNWNtITbUKw/ZjmDcysKY2
g/gdf4FDqMFCSQm1M35DQiVbPl7lVarBGhgYj5jNvD5GRbCrJPDP3gM2Km8URN78
ObhnkuyzvkgnCaSNGHQVyDjzeryP3MnDA/t0OvH544T3HqvRGriqxdrM77DDSArI
u5efJAICiMfCCq1Qxx3hqazfkkEHZid4yJK61bKc1J0EsspuO+D5VY6f5ZTcP/2U
BUZYi2U3JtwwLmxHvLJHRLDOCvvypTIoe80lmg8aZfpTEFi57nPlpCTqIupLHhx7
Aph6aqb4dOpocWcIqErKX13Fo+r/XJK9RuTv0EqO8si5QUDm1M2FMgwXU9smRWgi
ZRDJRvKdeNT0+GJQr6/N4fReLCRxbTK9UiQQc5uVYarDgmSm6DS0aK7i68dCP9aU
aD/TAew+GO6XBQGN/eNBbBkMxr1Jh7Ekcg4mB4IQFgQolZdrJIvMBU60cna8tmh/
P3W8VnqpCaS0h3isTjQW9bbXnuaRQtvslOWpgb7H7n1PCmj/eloZ+aBMOps63LBn
hZYU9b5t6wEo3reX6hMOGrZr5jKLFmLm6290P86SpGUzjogsRogvnMgKZT5RcxjD
M2SioU3qMvNRD+iAFAS78n5Bj97m/S3vaEJLN+3OFvsCVA7gYYT39xpfWs0teaM6
1pDBJIjSEx+jJX6mvcTHv5phCaDZZI2MgGEOnySNKEUwYwPn/KWpNGFlFmElnoJg
QVby7kbDnGQrNhUPnQuT7gTsAbkvnL+f2yQFJ1KDZjpiNYE41HVpXzslYEP3QOs/
Jrk3tn6prSKyMIj4NE9lBDYMOAyAT4D8ZB+SBxacplK1jeGxc2KA14lPrGHoxjM4
CzK5NgEAL3C6hn10PxPhtt+KHRL21OLr4HcqOfjBdkrfQrrsT+OeT1G2aspuNMQ4
IliIBkuDC1Ve5fkI7onJGbCbICxcZhNFyxpeqdTnCst1vJ6YY07bvhcuSzHW5SRm
063XkPWhoVXBJFH9fCQw0Xx1j0B5WtxseMoxyBicTd1SHhBskuzqFnGaDWlqRnR1
yAKAMoWZcVgOdb8UCU4xi43eOdQwVoEhoMwXOIwMhNzbYYL0znI47rbYKqnPrBCY
uFaKt6/9CvhI14glo59jowsXanHFMm4Fdc316JOpsBifahbPOjaSpyJg+8TsJfyc
IWDZ0oVogyzxnykWlO39dfsb6Pc81n276OPUbQEoJqMJU5xymJOKvXQIbgnlhd4r
TLE4bXlquPzTQucAEOj10H2YYFwxKscGoo/+pNFiY40KLxM8pqxxoOH+nBvlE7lV
N6egm9s/02VTD/210T1X58qK7Z8LzjX9bPvL6CX0JxuZtyKQGnbiMK1lSSvHdF7x
T/YDOxcD/ceAXG8N5KTWBcwIFWQe2rTnF+aS+HS+DuW7bkY9x1g7W/4nsc7wUppr
APqf6SlQjx8en/mR5qMq5xcTlY/t7p5P466SVKs8rwN1kPSGwiXaWq/CkMEY9kwS
C5zDos1aur/EF5E+hLaxDinGSCYhlDHP+VTMEHosUooxjvOA9ySO6L4hIpiWI87Z
ahAjtc77k2h8FZld3yM797HAGAVAyR662c5gbIAbllyYit9pISo2hu64F0XRMrtf
GB0EHzlswm5FlIgmGMPH4+nwLVSezVEGrMEGK7k1ORatNI0Ail+HxQ5T7ZOBdPlW
z3aa8ApZxujV4BAlir04OAwu9CHvpw12c1ZRQCH9hdWUobEV+aaqZcMCwk5csjDu
b41WRKpnTZzoPzdh/oQANyyFNkv7VsA0+XNd+r86x4Ybarlivf7qmvFIs6eHwdTA
Fg3WVR/QMjfd4vMz1H0prB+UnHMPQdv+t1TK6Aw+8ruEeR7Zx6hrZbupfSWIfd6R
Mkag+572EwlFEYR6S6niGfeo0w91TwvnFQ9jExVb46sx80qf4z4sJLMIO6hZafnv
LOcljjC4ocNSD50ykOtBcJ5UfcAKU5Gt2E/fnQvFHRSYCkq2t5MYa3GQBYt+iFmf
A6UwOCFShNEcdZ2JgqvtBRwl9qXe8ysq7h8TsW2KLoFMXsSD6Wa9RsWRoIJ1lb2s
5Tfpn40Bsowg2ZbnNJZxZDJgSi4QWbTnup9s63kzTwDftERsq6jZU5OyB6LXgO6c
eytksx/qkN80wpAqlKuz7AJbjTxH72mMFlMzDpewy7+DHS49ezJ0nWbqSalWsVs2
b7+2lGNPerOYCTZ7dL8C8Xdwv550aRZUo9JmIJXKhTTB3NeXrzj+3zYdw29Iv2nA
EOta60QKU/Os8nlJWlOgUMzQrd/M1KM1gMOvJdqY/lhSkkvs3oVdVh6WORfqX1CU
eqq/oAIfARmX9ZxwfVWAB9hLPcpIZ+wljfrCSp76U5JaIR1g5+CUCPjUrd7n6gS6
C8M/TXNXK6T9QtZxRDfb898lAw97+iPAxQlkKO40yTxJ6bL3BJ3nIRoHvTBAC1K8
XAby0WSmGEI9TpBdlUVI7TehvYdW9qoCo0CwdeP14dc7YdIzwzkzYwv1VWM1XmAu
kChLjgw8w4IhPtB2oB8Ai3zaGniLW+EMpOefiqIws+VbdWb/ThODeGkmmt0poH79
OJok72lha4oJSUeFkU85RSEUhBzHwF8xrSBggCpjq30B1NdVzRBhDpl/5I55WZtw
Dy1FrKjJiwZCiw36JPB/UXekIGybcIp4j7IlDiCcnMiUymmrGBYeuXcO7JddZdO7
6FDsM0pcrloBJ/Xr0gkX8fbADTh2w4Lf36jaJAoAywkX2lZdOZ3L1TUd5CH3pXUP
v4DFXsXaZr9DBQfKy/jBHpbe6e/tOOYBSh2+l3QmOOmVav0BK7zWUterThy0Qg7k
3N/CcUfJP5ZYTi4XR9LWbAgmOdt/2EIuB3vy7i5jTYLuOUOdO5pqqKgZfy4OjxeC
qdq1kz/XV2WaekYXgzL4E87K6tSch0pb98V/CngP/lMwIObzulVmnJ5wiA3hfnZO
H5nnYZec7B+3oGEAV3OieVtEbpv4BWCR8ueL2n1TLmVQbABCi89RM+fzvQc2hcoO
TJQImGnODL9oGm0Q2/47iPWPZ74Lah5M7O4LRe/TpPa+DnOPaAHpxWEa0R1F5QTD
iYDELgB7HWJA6j6nU2Kv7BQxy891JcLgZ9DfTyPPb6WQmBj76mhGUm6vulRI5ILb
mp3NZTl1LSszBjcK6+v5ZVgYdYewmiOBET5QJ5IZLJUYS5zoKLfnEZQQBaIOnt40
ZGT1gdSATrC5JTr8Ek6qACFR2803QuDVZxt54QNZspdzL7C6y3akkDCghwpiCM0B
xd4uUDPyLerXFqWe+iH7uGlo+ar0+HnFdfgelXGR5fFGrYvD4PJiNZgVDwQ3FpAX
0OMe3EI/94z3NwovgTv65luOHbGKiTvNA4Qr6V1f8SnSdsRJN/42xiErRJUNS6yo
n5GlSwpZlzPJGXWkNCiLJo6fPDFwRgs3iXJa/BcUK63jAb8YlyH6VGc3Dda/X4Ei
y1I6KyjL8JfkerghRl/T8ADVtTZY39JF3b6/ZBGKEQ2dOFUfx1WyaARpUEs5wxC2
sZAXgOWI3IN8BNKlWwYmSLPBYLvYbWDmGagQjAnbZQgtgWJ0q5ropxlAfor7xSpe
HWSzvNal8wwbqnWjb4rNOKDPKkKcZV2k2jERDPc4nNyy+X6T0KRH2HRBusS56IwW
+PQeSRKLTTWJL1mGfuapkxJoB7tSN5NV4R/Oo5LuUhsi8KqRfeo8dvvdk32dY56u
hZYOrTaSYny7lgqf4V5GK04s/8inBbV+6RMCI8qk8zINU9FI3ye7TxdAg/EBV2s5
MhcE1K/2tm4vsAFSMmc47Cb0p6fjOTiUQEsSgae3VIAYQm/yog6UFpHEb48TdO7I
n6OjRis7IM4Rqf7L1/mwLAGDCe0vXiQ1FOvgJNXrG4IHCzBVVyWXUawK9yEF6k7o
eGZM1NCTuBiAYk2Pm/Gu4wiHujqGh0OxLwddGBGZSNkBwuvkfDgojtcur1vKibxM
kz+6oJ/sosLonGTzxzWYchs/fAxWukKUy+5qQ87ADaW8hjwmnHGylfGn5Fw7Jn42
BqdPUB80Kify/JgoV9aOpwVxK+tqDxjjfweY+ku7fNGeQ10nzinpa3g8oVXpTYoK
6m9xfiRjSKhvyavrvMwTYMePbxvo3QuJDOiLi7vyk1Qz7ApPP8DVBoZxgdWSXzRk
01Sxy2NS6HihHNXWIhLFdTcnFrN/0/r9xOguMFuI1HAQKSAZoRRpkemg3Xtov/VI
8mLC4HccF2tmRRUxFjkSPUY9w6DkwzAw3WDFITgeTvf+TsbFI0Cseg76AYnLCld4
29Pt0mK6Wzn8eTd46Qnm8PH/3Eq96BYdJxvCm8qrZ69XlylJUPwu5q7Qw0pdP/Cl
9I0SSVMzxaSZLy7+l719WSKKCt1WY1elqrCmlmyL07hJVEyeW2DjGop7L493A7Nw
yWSW9CxLXOBQnCj3pYqVnyoGelOmbMKlmMroK0O0u3br2ACdVbliSPS9LQ59wpV6
Ohb8mJihS3IyEa/ZK0cNeu6BDLL3sR1mkujqf5Nfw5r3UvDtYUgnKz6uYgTa3FE5
m8SbtFwIWbNRnAub1Zf3hULqHJ2nERFVFHkADi1EyrN8WJcRyxwdAs3CTwF5vXbb
LiqF8y8pz8KskVVK3SjYOwLjmcaXusTFwEHHBPHTSdXoVRZW9PAqINEjOY8GIjCg
5WRnTKfnIr9p6wevZ0QVFItQyFt010HbxxUNQRUpQld2XNdQ3W+CCJGzHedGCCvX
q/vmlbhebYV56PyBQhHwXs+2mh3txTFR6OLQzrJPg82bBy96OdHPaMspkOw6tRaN
s63Z6Zby4y0LbDLRv+rbwDZkIVAdE9wJE9cUT4EWNHHSLCH4tBfBexZYNpZMNyPS
tONOxrXVn9L+HL2bJFDBtwrl5fod8J2DiA4/g1RXRVjQ3/nvQCiYYHmPgP8CcENV
pULJT5evrKSNdUFpQd5ZWX6o23P1b4q3iX/3PstuexJVlPnLPH0jWgHt9kqspCaM
wQPRmzx2kIdkxN7pMLzYXd10AdAba4lKNCmV2K4bVA1aFN78RoByMjmdUvp8F37z
juB2Wfjaws7YQEC41fq3NpZDgWmtI7bdgEJH/eHYDYEJWhNJwLyG2/ANPvb0Gcmp
a/1wedOsaRDONl9a7WifsyOsV2YutkcdNFvXXmuxiPPyRjyYfN7zTTbQKGiMcaFh
DNoCb91xWLHXcqjdUWqLjTBpNgcQLioCgpdR20JNBuoCDjxdaxQCWHCvAtcb9LFE
IcjHWuoOMIQhQfZ1DPMQ7Vh7b10+MzOMvwfAgmo0bIzulKfHMBvLh9Ol72gtLLDs
YB7DGZ9duZyE8p8IU4RuHbZPIvWbgBi4pc25Y9Rsfm63uZBPz0To8Yg6tNCY+75i
nIAJzz5CwXaOQcwPg5em25c/eqceQHpWOnFpiuBhyjkCtycGZfQuQ0XmUOzwOyYl
k+1V4PlVK8mXsh/qMSmuSteHqI4ZwWV7y/RVhxt8TccSqJkBCcsOXI9/GzecNQJL
/fWp+zEkO9bxW8VehK/qLvrWb0g+8uPoZSCxK5qHE4InXTcwGSKcnMspZcrMSmLE
c5nLdkyYT8f1vBZFo3pM2NEEU4o3ILYEFiL/KzJ6DqyUVScy25a7Wx/s3RoTszni
VRH182XeRpd1XXH68O/RUM0DIUJLxbuY3/8vTxZ8WtMw91wYG7DlhGUMeXw0iLaF
TbRO869FcTDnqxrzmL+WZh5h84JTh7B3fXErQCCp67bch9YKNYSUvKOeA5/6FF3y
wet0SMJ1t5XVr/DfLTPP/pdOJ+GdB2Pcq5wAVGaWpLEBqRtZq4puGcEGaWyIApDX
e1yNROWqwGzrbRaCW1UBwZgBGNrGQBeIJangiZ/x+Lb5Sfv232IhbgLmJjGxtfeU
du2wGUc4ZMBARbq61qKSmBXPbSZFX9MknsPB7I57KxryAgcc8R/PXLyGTCJPwrhu
N8bIlc2fUQbghwHjiwpmddKWKGqbPgtj2nCzuDoDeUB4BCUQbqwrj5DEWDBonKUo
8bQn21m1fBpSje73D/choswI13d6aGPouAhWXGRE0sHVaW2X3g+VG3meF25By10U
ibqKP86kTSKrFsWmB+qPsP6HroqdV9BO6YWXW3eThqopa82K9jvStbHPWDY2sQfq
KnQWGO0PyeMQlv+EfKHNRbGw1NCpaignRWVxJtNxS5i41O0A3iTMzh54b+/xwjN7
zwWXQ9H+1rga0vpIFRv70GZdt6O9itWPl7Cf9xHzMaxrLNHE72NSqFPi1/oViG04
61rDlxuDaRsSkVs/B9vmcj4OKxrsx60aTzMl1fWkZW6M0L+TkwmPsSz+uR1HHLW2
LDFsf7oPgBCgYwhyv2cesJwEiXR2jdj/8ZMmz/bzg9DZfWs18/QM6+VUhPywIJR2
gXDK5VLV4f6JwvgKixi4ZLI4W7QjN+vZtAaTuCzNFmGhAVNytfRmxpJGKOcyZujp
l3DaIn1wAslCdMmg+nV0MBl2RPtiEyz4Bmnm/HtfRU/4v3LM1XC0jjk/zv/tXeqF
gSg1vMRLbqdFUXBL8g4nKgRez5TsiqrU8Po+MGX6ZD0ICdoPPJgwHPejDQPD8pYY
6RV0kuxdcTUYY8eLpqUey8ZO/EQz35CBFqXWjQRMyrP6AamuP7Z/QYk6sopjOAcL
gLQOYAm13ry3uTYl18W73otHrqY0DLQX/JlXGbtSv+557X8e5yoQcJwwSoaZYRtG
CCu7qLK/3+wAZT7tluwZps38JWUpxxXUA0up2vKVPeHOuBHjn7450fK0nn0nhsu+
SOuYmQmo66AUuYPSjdNYc1uDiOktPmGqRJfKviknB949LWWEsMvbIZIe+POUcRdf
MaA6RDqVS64UcLVsFImojiOG7ty5YYmvJtKlQeaZlRGKrZJUTUvgmuglHM1GFv/U
heSEBWcPwC5JCaXiEH9OO9Lh1frzqStsJbNmSKv40KaLtepaQUfGuVHjvyQchhD2
r2HsgxFNNq3sGGy/YdkVwU6Qj1RTb1TeB3gRrOm0m/lBLcuzv09dY/8Ng4mR+ifb
X1Z1VluijWGoUMw+UvidJE1aBIKs6P1zvPI0eCD0OkQUgyTF+RBXVivXomXpUt8o
kq+BtJljLR7E+Z1/k0K6OGPEMCY7KEtTKs7MR9T5kArS4dSDNZ9HEiMATMF5SNtU
+ngb9a3ZLTxEN2E1eyPi9np23PjQowzmBGlA6g+WctnfpKKjuLv4ZdtTFkXFeY/f
Hmlsq70uFIdz9D6o1R2o+qRH6TS/a4YKMvh1OIjnmhsyB4/Ax4Ouve5yOtdyaAqu
uhKtT9AyV/lBn+PTWJ61cIq90TXQfDqeSoopwAafLVwFYCGHGqepzNvpncM4B5i1
jfgC8ocg7ORvj3wwh+Nwao4cI6Si5B27EupwWCD3+yVRG6JGK6+cBNojqdaA2x5p
sO35LnF5H9hDi3wAWY4YH8ohSwCkEt9eVtbWG1i/aBlPdXT7OGT3Uy1ziOOOfU8R
T/lIzMYAvZxE7VWVUo6oQk4mY76xugF1UwskdbwirEDsZcluGE1RPFfZtgpw1Vck
dbZZ+KgPR/3EAnKZyNzlc+5zMbJohNRznGr3z7bGwqSo9DF5S2ECRclIhc0XOD18
5aAORTM50uLohDTnH+UmeED2DnONuXgk2OIcz87UgEvDRqHHOQSh3erMP32PKdun
DmVYVV4Q5wlf4qPozYf99J4VviNngbsX5wo0HaZDQo5JZU1qNR56KgPU7F2icLyF
11vBtEI5Z0zJQG5M1XQxi8GW/M4Hq5VyIT7WJzRc/vdMEAVcVUNQMUlVMgpLph9K
AwNF9X2x++u+0JulzdsJHALyU//Q+AwxfrRYDMC5Qt9X+SA+cEyNKlmcVo9aTR/C
uzrjrISrhXerY1PlL0HNJuAug3YXi0zWi91SAL6A842jUg4/bYcQMURCbjC0yTSd
gwiEPZDSf+kC9aCn+JcJ8EX+fm4IBuvVsaGvnL6DIquS4yHK6AmOqYCMjVvGzruk
+QWVxm6svHvbamkV2rt8ZJOyLtcpYSJRNy5yGNJccg+q7vw9525Fj/hTtmlUqb9s
QQTQjh+Bz94kbE5d6DJkYQ/FxLcezfsj0/847raxEgQYF8qNIiVqyVpWUoeWDSQT
GCOC4ZdiSLl3vETw0F16iNQpG9ShE2OkasJ/Pc78zzTgAbRzveuz3rXKDbhYVBv/
LIU7+U8PwvooLEqYuFpLq3/dDomjnbw70Isi/+5MYMiNf0GS81+9Sk5t/G8un2tl
j2sQK/9Goyl6cWmQl0Cih3yIX0yk+zH2vidNwVvwoAAHocTaYDRHtTM9rAbOiwzG
Bi/qJqF2fpbal6HxrjaY/eFhrsRm5cW6ZXR1Ui41HtauttlNNZJKYb6WYtuOXnkx
9ozn2IU593cGUHH747Fi0dA+EkurdZP/C1dUj56LY/2QjsGyH2osEMVymgVN/KSl
Czl9ggdiTEDmnnxjQfY+D1Imcz0XrAlDlETO5cgQh9sFeRXUnB76IDUnoBzvHI8Y
v/TQ/4fxheB6c66y8EEvLCAs9latcAUEXfyvmGp02tV0vT3raGInxsFIlWu6+60K
vladjRvaNKE0l/MPqgKHDHCza7ftucYdXFn3yzefDEtu1tqzy61QitUb2qSEV7tH
bMBZvMEukgvh/N0qHXeoj7wk+Mf5ABZbX6LocFn2JEBERaFPCSv3uTPrN+qm4men
14oedATCgG7cFv/ZwTaazI+G6FYL4FQyH8AdJiZTETpuWdQnE7WuPgAuxrubpUU1
VN1tmIw0GtoHWjU255z1PrRjIPqKwX6PozzCl51Tra6dUsutz5Q2H+TxNXnqMxh4
y9Hnzkc8CWAjn23WQuNl9t46zmtS7sKRGW8QyupQaAwyzXjngOrZ6SmufVGb4AG0
CKDzf6E9T9jjKxe+AzpdrVYhJraa7lGlHli4cHzYdjLuadbdmX3CImVznIq0JhkM
52+Hu9M1Db29phcXTs+8feTBQzvymL2Qx8LERX06S0EGV1fnK7A69w7Rdf3mUjLo
sN9awVDsRPtLGNucR3j/egf2zQ3zTVlRj3BHNVc9wxR6fWD1HMuso2T6Uv3YWaUz
1sjIJnJL7TdTnPWv+go2tzUHWDyKJ0lfKHY+81x53uictcHdC84i/c8qor+6lQTr
T2oKc4Q40GAmYH9f5xveFA0KKtHB4by/TET9uPoJJG8ckIsoR4w5d6LuI8gERUnP
lS7jhPp5xbTdGqr6zCg2Em42pTP1BhoxNHM1SekuxKjTcSBOe+n8FPVU9u+CYlTf
UY2qQmcZsNDL5oQw36hMBmyoP3UnRLb0ICGvbaZ82TY8DiS80yY7wR0V4ZF64Jw/
NptfKoYFwY6XO/udnSWepADmMza3TyjcHAxLyFeimKA42ylNtK6encoHjJemzj+N
3myoO3SikIE2TjAAMc/PYzqheS1wcmj34H324aB9kGOuWmaRs9RjuHP0/4Bc0Tmx
CjT7E+GOMLmQpxmD3J+Y2UUhkkrSh7/BfWpy1qC7qIuhl9wgsDbg2cgTpOh7ndzF
uVjyK1GDVfA2vlHVY+d8ISrsxVbho8OHQpeMhy9y2d7WvWbRzg6I+59okgPXAJhZ
VEEoNzgnrvotpG8wiOJMg8uBfZ1SzX6vaz/1/+M90t2f50Vb7bHCRIeHCaUQdh8B
/1Fr2VOIjLUdNIld70Xl9PY0MGZ77lRLnydVAk+++WbqYqYKzrxVNCb5MQcqk8fq
khFSfGLajk4B5ovbhP36prAbLA6t7hIV2wr+2Jxl0B13cd9TBLmqw/6YnKlUYahi
IHEXUcTZLQSvLeWiJhHevxWZ4PM5rHtriAO+3uADtymX4wCJv3crj3s/jktsKawJ
1B0c6GhEPib9yIKCkQauaRhQdWyEbQFX7pW1TWj4L1rtaMJC9xewYv0TgX328fNZ
ptVA1/x75m7OEJSxjKkEzUB0hz9PxR4wm0Ne/oHbOX0GImq1TumzOjF3HW8HrCWU
Mt19idwvEFWvb7m5Lcr7myh/oOF7hgOQrTKxBt9JOcudsZGyb3T2UwYazsrVe1YC
/fXd1gXFwdqSBPVZeQieOWSvRdqczgbZenY7XxyXNN5HHsDJnUXhAv9I9VyFhHlp
eKx7nuCew0qka4WULI8YBZbsAwo7sX+J8RATYePUC12L5wDGtOBIBNCu97navv9q
VYMyoGPHpkQ6H5csO74uWu2GF7fozF+O3nOFGW+4IYeDAi7mcMbghYI40t/P6iMi
J1+Ja5GCOcofuFQgFlTHvCg/V/Jgdtg4ZsEpYxQuUD1BxHWVhcFJXGKl2PYFnbrC
7uIK0On7Gfsi+62fG2TCPlbHx89QLpqqVWRRY7bhK+MV1jHpXqLHKIxN1nZ85hyX
c2IUAUvYaO94S3fSB7ee0UeLXIoyQPDZHp8zFBFSMliytxuQdOg5ZxgZNTv5vyvp
5Y1OtiUozgTgSweCkUCyzB7z266VKh3Ggp2imHDH1NwuxF22POihTUMf8uiyS259
YoefCVAWbMiUq2KwqGiO+BFzB2nD7eSadI9k06L4tB//ep+qgWzRHQaI4folC4S+
Ris00RcFWb7VLKjVGcnPc2xn8tUHiFMXvIZiveDrl+qdD4anxZ1TkYeKTa1pif2f
M3Yxm9RqWYQmdYrYUCn/J9un1T1BI4RdSsLHX4jB2ymr6HhFtfJ1rGfbPoiQy3XO
iN+dSGMC0S5zAk4mRaGtGzV98P4yYwl52hBviJBfRLHYHHp9Wfm0BNdn8AD2UYvJ
FUU9mT0F6VjYMimX6B+Z6tjXE7B5sjaIkj8mE8lGS2zY5IpG1G04JZVpHC1SeZOc
wrqCiARUtAKiF797cNNDpLOD0lh7vhKwFPg9tAhMPsDm+g+8oVA9f1bA2G9jlltx
3++9hbth2XGsEwo9WYI0KovjFykchfnO0tqeCMPP/RWjwN68QY8KBajc5VILNFFd
TbpsKHQ6IKa1bUBMwOuOIp6io4/nif/s3kpTNhVun/fkC0H3WNDGqBVwUV+5svEJ
jHBXYp1R0eQu971PmdZ1nOc/6b5Hrb7v1e23rgRfU3BNMsBnpKMvzDJa4sCRM6bq
ju3ZYcX8TW8cDtGVQZioAlmhheh80/OzQCRFwUf6ztYBX+zuCGDLtSWwoLETQX7T
mgkUg+aixmByHV7ZiRf1Bn35Kl5geqyajeOp0465ieScvOkTvT1R02FkjnmPJ4Wq
Q3lBDs4gisf3YRgHoJoRyQ4Dr8DjcbvmlMM+MWtL3Jj+U5+tkcuoHzCI8/Oenqnd
o+Y4zYGpbQrgdWB8U0zLAJjZQfmHh0l+hvE8ZugaBYBL3Er9vJaG4/3ymRNSP+f/
rUvh1xnGyNVnV8AKpIuZovTCYOPn/5v1UjnfQJY0L7AWakyDFaDRuZrq8qq+KtFL
vagzmgCi7dNRUTZ0nw3BwRI53u5fDYq8KYEeB8RrVBCeIbA9q9CnDyxvpCwFcV8l
7xAuVMIsazJsafNjiDVzcHEznj9GNEDo7GTbtZCz2YyFrxsGt4J/mAmCrlw3GfFh
Ma30re0BomkNcFiasY4wzkFfbqL4ryDPIiNo/uG3OA9HamJnzG/oTyUDlu0VcMYP
39kDOlN9vqoJgyB9o8kieXkGrhUvSIkKskm9T6pt1DESfWm07A1NxbLWeb+aPAZf
e64fVOYftPMw6BBbxP1AII9kqBavwVU5ru4gsfvWumidPntOtddMO3dhpuUXuvgJ
lvowME6wr2vMXuRCG7s9yzNvIqvnABgokOrBbq9nEpk+Fd7sfVG1+Glfj/+y75vH
RxoSWI8/JgQfE92uyaWK+8dupQHl3gR3ZhDi7u7/gBHiIkAujNDKSrB587hkCaCE
JrfI0L/mSn4GP26uB7lPpeleodfPqexCEFxoYZvbF0qT8+P6THvnq/ytaxS6Vp5p
ICJuS1KgJYGEsWltfUBJ4i+79oM6TT0r5vWSjUGGwJsEwr/nGsJ2nT2PP90ZSPpq
aVA83cNLybKZVC/d46+NsHqMOhC0KK0aAFC47LoIu+XA4I1lQlY/qIz0VYgHc6In
eIXlPf92pBOrVs7Qv8fh7q1TetuqPcPGXwvLBBd9cgD+eyIw0IYwd6lDVCP/UKlC
kjRI+AuX/59LCjG3VAocV0B7VenXg+taVPGz8Ogc7bmFW0TSzUqOTAUuLjaheF22
9IJLA6zgCGT0O4Dkvx0RuUIweeXbXvKZwBRp94RpuknbuhGv2x0V1g2g5Vc+hbfc
B9I8xfjiAgPnM5t7JD9prUY46QdgI5uVzt2E6KTikuOVk9V2A7N/I6W9dtbPdpQY
esXLk6L8RnydrDzH/p4Y1o9VBgl5bFQka83s+u9B47GAddq1mUufTJxP1E+GKC16
Ui5g/R3ZjxRe8Y/NkFR0Tlo1rymj15ZBsTUSOfedZ9JWrsCovPpGyagWhhd6+Uon
PKOt9sk3eR4tGjJQiazHqxDCZNDrCrqGTmchLUkg9skCMQ93Ra/Pj5ZcDdf0gutb
G/uj44oJWDWi0XNGgDtzVqAz3pe+MSaJf1XXRVi1y2ebBx5qb/HuiHLoaXdu1YCi
ICb4zf96EN1q7udY6Lr/ybskwfTyzsBqyfXmgN0SWfmMJ9R6KWOhP8cCPR5+YUYH
/WhDcQ3/W2j5gzsIpnlyOqoFjse+QR2Z9NE/hB88GsZjseK3MAniOR8d6+MegyZy
JGqrW0ix8uvXkGcNG3BSTZCCQ4UUm0uTsbH2sam5y277Ti+iM8gC7l4JiVPh8pD4
U/ivw7Wn0D9VbhcnXU/sT6OlZ4USJD26BcpDgdBDmajPgegJtQlyqcFmNCEbrgyr
kaeAsU/fySRvdwOePqmuOcKvxmFL/lnx6UiYtnBDGOL2Swe6CwPCwSOUH3WP9ixy
KFQm41cnHZt45UyQFB6Z34DR2QZgXaf/A2t2K4iqhgWJyLrDkOOwebglYlrujZtn
//q4HObl6Nb5AJo+ShsitQgLP1aXvIlmJ91ml1IBWRQngwi7Tjwv9OH8hC5ZuNGn
HGnqakKRAbtg3NDQE28d860/R99O0BcXt+4Ny6rx/zVFZgEfaRhyJGu/F3peR8xm
tLEc9TNpMlsYkYhox+jBMX94STwYppEW2c/OfgePJU6DfnvaAl+VpNSTM+gdz1O6
HE4CaiT9nXhEO3vd2MzTkdyuOFHbOFlNjEbdUS7m1eBxkZMq3maWI0rmB54w/Mbv
R1Q4REvHJlk61Otp0lN4wsXIN81c0ADmYe0TVfiWITvFkYU+X+0c6cC2rZtAd3tU
BRGYPZtJGpIC2eXUSu/+Ov8KUmBDhU59oYCPh+kJxcb0bKweLov7q9Pb7wbNE0IS
7q6KwcezISB/98iq2G40ek0fQWHpIQqYbSuxm3AuGq0t9+dqa2Q4vyDwiuTw+4ni
5av/eu1ej8d/loCyVcra4hBaVB/B8qmYJu8XNkQWXDvQLP09kkFAOarWh690mj1o
pJil9dkC7NqmxuxZG51BS64Zd7iwxxaS0RjYn0o5CCX5JyzdPfqH0bA8onIHoXIO
gWy975whqH6cLaXywmASfmZrmD/EmGpb2bHMCqLJmYRuN+yfj9U6gvimu7OCuYp4
lM2dHrJLnBtF5eXyKRgUze6fxNHI9QLKNbqpHvmmq5Ycqu/MeWZJKTs5aTGl8/zN
Epn3YAY5jjZ0XPECJDARo3/o2KJ0V+yvht3geq1ren1I/Z1d9uEkZXncFonSiD9D
3ruu+77Dd8O5TYTp8jGaBno3O1ogUkCtjfNUbh3z4ZvA/dNtPTyODCPUdzp0Xy6r
4zV0697MkX8oU3MiDBVS+ptxyI2VNKBJsTtivfJaFrBMNF9IC2dRB86Ybcstj9WO
As5HtypSJzdomFscQ4juJ/RIJrSY3SgT8O4OCRFA2dd4/12mOoAs2y9cwSQDJISD
f0zE88j6hR9v7j4yNH7X8GVrEFg5FahcgEGsoY9LkUlyyX86J0MypAFtJ1bs3IjR
IsrIdPDhYD2wZyVtzZ2t/L+wlvLv/QClIsGUh1Y4eZiL4AljLHCPKeEuB9m5gYZP
95Jig+GPxXxm3kmC0kjdEektB32QxVPmWY7CwZU+CaatDKSqFopqd5m2WcJMfDKm
h7aYRp/Fc7scWK7TfqgMYy5OSXVySXDiu64E2h4funsUdt2NWuEqh1OXheolG4fO
cxZ54nwkYWEExq/H0Sykn8WjMxUBgVCRBUaEa7JJ/hMndXI0Wrorntk7+GurS8oT
1xMXESROdrwkBkAiiUBCUQtHGAPi4l8U0fgY8iHV4GytIIgOcPs8WgECZGqibjNv
GyYryPRnwAzuXugLeOnViQWZT8wQlT8xRACn1ODgu07lovPx9eo2Yu7gbA4tGNra
yYD54/KUkAHRN8JvfrIqHO+3rxTdLscUifpsNodQq+YbwkQ/kubccOzMQf0lkcRx
6NMX1QJKtR/Fxq2kGouX451p5AfsyvQFOFVi4Lv2ZhR21SOM0WZh6bTk/uDppgef
QU1ZS3MDZkW3R6b0d85FuaXASU9b0V6xkjWmroWEIijECWek2XT6/uU0JEXI0JKL
vx4fiDRT5+T0sbkOjYiSdLJWIfo63IRoYLezpkNKYbrmsAbrOKG8/p/OAZ4KM+tG
axo38wDnjVYj3hdYFyU1VQTBwFFTncXqaTqAFnUIdymRgBnyliZdbY2H/mQEuWnC
upUg6CuFBXtR+c2seVatTtGBGM6sHr3hybN9dKmvSCoKEJQXBeW8XjLXno4QKW+x
20kil5itrT6DABiR6gNam+H8YWg33JKMQ5mrOwnKYGp6Vrz78itjo9Cy7gLVSYtx
b2ESJXKKeEGlsBR8GRMDNZ7dQsPH5sI7yDwKfjrWmG1eGaoj2NRcGu74YstkaTdb
Vx1+t6sS6YX5j98ZJ0llEqbCLQYbvzaHLv+kjTp8FcGcPdkKTiwfSVtXeAoKok4x
POarSpfzWRPSCf5fEvColzmmHDnEg3YZ70dccl/vETzCt026ss/Vaz4KwzQj1DuI
GMdYL3beh3rjCr1Ir2FplIB++jSGtmVzEpSto3LYUgtfSPYxvsCdsTsbIOqDQgRY
PDbGSK7+ifV7bHASx8YMTIKN+B9kL0Z5mr01L/mFkpUYtPw00QvbvB0XaW9s1Hk8
Nh6znz3NmEZHp2DCOg4Djco7/LWpaIK5L2ekW3f2doTxwUy5ielAaiF+ZfZW7UZ1
pzY7ZsWwW3UKU3OTb1dYrQgsl08K+kyUVajSPaETAC9lA/rj5oFvpVBPo1DOZuqy
4VVzHXqP5U2vh3Yq8L73hRWxKKVSTOhPRWxsf3kxfYX7g9uhMhLagxPfVK/jxEfb
8Ct3iG9Vo8cCGF94zm1LRJpyp/Nb0m7KP+T75HD3JkqvmQbojjCdQGEa0xMVN0VF
c5j21JNNA5uxbR0MT30ADMbunjKHa2sK57cXPrp5YLbj7mn8kEAUwqbNddcTZzBV
anD0NNGSRaOgur2qa9vMrL7zgH9ByIi9oIn7Dmr3nzWp/S9YFF97DqZhW1BZTaFM
Bm4BmvFoPiyCdhWL4CFaJ6mpfFjE3DKMEh49cxytSuS8C0/rRHk+tJURLgnb+thr
20eh++VwiKoRlTax9K/BXiKvi/6qrs9TRj20foOfazp5b9cqjVQNgnuD4A6Afrn2
yDEgGTP9i1sEA9BsuwS9BkwOIbT+KDoDaFCeZTJhdqLOSnH6hdJ3/0gb5ABE6Dc6
ZncOLEp+gnVpepYGRQ4oP1QJvS52SoU08LNXjEz5SPAmzjsrDlur/SCcr5HIAkCT
izIopltKv5EZqnfJJWigVTev3uubiDBss4GebT0l2DPIty2dqyrCPnhit1Vkpush
fxHzNzdYM+XrVcZTyL9MoWf1fz3raL8CJRniR+JAjnfwECX60N4vnN/lrHwb5Ozl
mS93f4WAo6UQ9WW7nxuMrq0cKtadEXp+iWsrAhrWZKtb1VGoDaGhiikatm8MVYyn
oY46GUJcy3PNr5W6j31FikjLlOQfxQALiOO9cF+x/izwO6cji5DLJsBjUK4PacJA
lRoxEcX6ch5D+BL5ug7OmhpL/N5kOdNtTU8DZR4Uo3MS4fxHz8l1dlYZMCKm90Fl
TsW5sZWc6yz4De57LJl5KVFuokSXIAss9Wludz/GOS9RHOBbGUd2yaC2ycGoAKBY
4Z18rigdjxvmN2qw2O6Ybm8TxSqbeqbe78gc8DbeWutAvb3zgMH5etXz3z1tjDmC
wgW0n1nA/ML0sFEuqIKP9K7nj/dyDMr+QA1J9Igjn+7MwHuavwQRe+R2m1JB7qJZ
YVKezWeVL/IrPk5RirAo61q/JVs7j30j/Er0/zvdKqoRV4T9LRKdyInuclGbYlJV
VqHJz2vhfz30pzRPTiSQh2XSxHgbPzsZBh5lSMUBFgaWvpyq2rGeyA/7v3geoTa/
KsSA1jmCEmCQ13W6dxR1N0p4EPj9E3TIiJyrIPiz+nn/0PfmOU+tjQE4QgronpV4
u9f+q1nJlHL0uuRuiisXoBlNQHrKT4pXHeOkr+JcHORw29+lBDYiT3kAh1/+D81a
XOlELO5jEzmizNVM4Ld4W62he5mcKGGqMtqyAC4o21T5Kyl7SZi7mI5+0HgJkuBn
fRe2zFov18U61B9TC6eSRbERIIg+9O0BeBJkSaeIxcYeenD2w2hRlwixey2VSOi6
LmgAFwlw70W4rwzoVuZhu8ARPnXh5EfTLWzfuJSktJufVUFZTf1n5INZsD1qcTED
omDl4/G4wcSAm5Q5t0Pr9ETu9o57iuu4/4tj3A4evBTtPMbkPe6RIAAmJ9NZ8ILx
gl+1l9Rlu7J9XLnX1OqV5v+8FBIsSvlf6rJBtllMf4YzKHt+PgyAjNKiOaBWBtKy
CMcl7G1ettgyatrdyfaAku/TGkazUo0r+GJmx/ZtW3pDuZHNHdJqGVox+2HMzzDM
A0Oi5IC436SACmbOzFfUuBbjfleACJkOTZaD7a3NIn/33w8/6btyv5w1IbfzM0bw
hUHuPXNZdbKvWt45MWd19cAdLX+47rQglfiffFe/5DufVmrEW0C6Ipsc4Nnwq8lM
K6g/h9Bn4fbN77NkfLLXssYDdmgYSsESNtH7X0TqhfijuX3AUOpe6iCON25GWZpm
CQmQoxCnGb+LpSsizqTnfNAB63seBBP0wRcYC+i+X3IcgGVOQAe5SM6AcwgfTl48
AAse8Ytk8qvdpDQ7pdFrTW/M6QZczFAn4fQha1tXn8sqj2BE7POzUp3wrj6CdAPc
ur6yOunz9qsPZhoZKN8dP8xxjBiYU6qZDMCJXeOaRTnZKs28kKuJGT3yEFZ39vz4
WHcjdT08BN4Hb7m/wDUke8nSQScPel56PIitKwbYHh+ZOHB0UEv1x7MLHsy3vaQ+
mafziF751A+1/gNsF4eLcM3/QuCWgED5xBWIUMNlioF5hWPvnlAJaq3Pbao8l4y9
x/D3HdYIbTqQqOR/f6xni0Ukh3HWtVHLyQgY+gfWc2xj1ON4qYzqdNkb4jfstmfl
TCmuzIscv72G+DFiC0rcUhpgZvrlTsD+1XBcvwizfxDq1ylknuSy5e3tgOW8iNRM
n3o2CSo3t2e4EhoHfgdtdcBwKAqEFe/M8+Oe4DEEF7LT6jRz84eOYYvUbyhVv7ya
FoN1r0gTsSB6GFgXW+FwZ+ipgUDFdGyrFv1vITEOixILC4UChVA76P0/WF9mi4Rp
TlCvwRG3ncnXQsBGZ+EE+GWX6iQxyoc8xHTcNCB7RszAMLQhx3nM6JtL7ZU0iP6l
/YL7WApOdXCyQBsY88a2PiCGG7qXf27ZjvVlOEzAygplA+epk2vDQZKwNgqUG1WS
NBu5nsjUm+LGyy4HzhB8u5sxlpdYFrq9cT+Q8WD8+3rE4Pk1bUXoQ4OJybcP1ngn
yEAbNw1dplKqhYwXNuCGUoWXDNbLGNk2UYZsdUohV97rY4NpLH6/2h1ghJPGrFXy
tceme4gB4I7Nm5dmFlCXuDgjvfl8b3WZPYX6ecReQA9VLnhVPRDD3D2o+OppiMZG
OQ70dObrPeB7SLhTNV0u044AIXZMAkz2CUiZKKxTGCCsarJaIkWgqENpt42vFtpN
tw87iyFRJLhy/aNmhemApuzGJcskpUopp11PKaV/xnZIhNvDjIOHdXRZf9hR6DTV
rxMzuIjUsYmfpkL0Q69dOukMcvhDDKFv251fqHHtVqFPZi+EIqI5fJv9DDMoqzYl
DagDnqdW1jYj7+NSRp8B87YnVTCo79aG8l3WAcZPS+FDd0puI1mcct5wF0hBQIRi
o4yLYEAYNFB3vXN10IR4jRBynUu8ZYEry5HmZjD2hTSyGia5CSl+Vc8wve3QO7MB
gviseQypKEl/QboHP4d1HDgHLWGlbzpAUlObfuQjcvGhJ6MztDnotfNShWUaylmL
xoiQgYHPEQhtrhIDi1QwWyX45A1oMBNeju5pA9nuuOLeF8CSc7377rxzufbtKI2Y
OPt78cmqqtseX16ivw3Fc0iK5jAZ3QzSe8vvW3k103g7ieen3gDuKKbPMtYdZAnG
VEvd7532iZT781c8PrUqLY/roFyLOTEGJNCwRjTTosA9OuVGe75MLOxWxzwe4xli
4DKP8aw3juTk6vyAbP+tX7uzfB5p43yeOgBv0YQcGDVV2yuvdzak5teogTTx9RgM
0wJvXxCIEyagKci5Her/Vbn8A3DnY8JyRv/JjBwKGBDpOPfGx57xKc4JQ68PF78x
i74e3aaFjXclzLmX0Yot458SS2jggURY2z2fo4iVKGT0yiwEBa67xj8Bf5+++I5t
H83nOVvKhDSirDxEMTAG8cKYaRUnEOVC/GL/OicwPYu+wdFdDAf82UfbaB+7ExEC
dCsQ1KgVDxo51fL+jgSQ9yrK8TBxYAyq9vyQfQxqFhaQrho1N9DJDzaS2cCxKHzg
3BN10ekCG5afi1sXgsrSttzIV0uRY0ODxsFrKkTCSaTa853yzWDUYRS29rENLrV+
fguQwCa/ERgsSlqyOC5b/b1AhvVZmo/gPtQIYG8LhdKMSkM+2X30lEYWlPCw7wCx
Luj3CQgjABHdV40ltPAf2g7DZPd9yyStjnDzoUBKcDoHUk/bBU3kaQpZN5sq7Syn
D+S2aGqLhr233enid3FQ+pBd6poFNYP0WlWE+hZvoC/+pv9yf1idmjdDFHOwzbvk
mb0Dxh/TZ2Nq4fAiP7/+j9sjKEoiQA0LO7fvvLBAEDbHF1rQmn3Q+qhjrhIN8T/+
/Ift/eQbbWRC/YuGu0u0LnN39cm6PT/7PMDaNml6K3pzaQU5q7paT2IXt/u2qd7F
59rMxrhYJZGVjJHWZi/r1XIhkTev219j0Zq9RI3LzQ58uPSley6tD/0vKlxTKx05
61PKJqwvINt25OXdGigrFvUwLDLSxsXUgtC5ArJgyY+m9IoAs66AIhebW+4bWXo8
szFzpK96Ay7ka1tEJ3gZkhHYSaSY9Th2ssdp7P9r+ny7n6Zc8XJr7tEMQvSvVeVu
dgvq38VQQ6irNyWJHuAKBHQ5lAgNLAquAM+Fa0jff2NUUa9pqbQow2M7UQAAiKJp
NOVpdstWoM7AEsG57Wn1IzdGsEKbmbX/ScvtD6KOrpysR4fO89B3o5MR4tacnniE
7N5ITVPYDdnfCCaW+kToll4JAkPwGfgBYqlToUYL40Bq2cGOSFzhZYJbDmyEKXzH
BVPNZe2SmoNAnZ6VTyWV/whI+CqNzSl+qwec3spXK2byesfFnZr8CFDyuaxBMWmg
HjHngWajEqZGrclyhO436A50OOWpy72jK1uIEE218nxAnBTrmtv1uZX5gdKWj1vP
nWSsp4pbbvuED/BvAJTvg6oAbjsf2lJ9pEtFkjihlxVcs5egWmLs15uhu4fHKvt1
+HDDD2UfUlo8ZP/tRmFUdqBBpvMungs6hEApq2i2pXmrgJkJxXoX2n71l+8MzI+G
8eDfMPcWvEPj1nK+FlfKhC5BD4OyAygxYDfUzEKCXMFn0PJ2voWVVrY8YzjkhIjG
Mr/X67pUrEe421qKGW0U7UsQjvxj2KZu9Ws5AOJsx/JBMESiSqOpcPf0ctB7I0fX
RZm3jg2PBc9TKOrzGbNi2rqujkIhwZGU6A9ESEDxOjkA0+/dih17hSILmby/fwen
CWQLY33VJ5dJKeER4OvBhTn72m1wg2YPqjOnjzVK2wKmiz5gCQuCfRARkavWhojv
q5sKI7Qusj+c45LKTWAo0+F8XHmfjRe8hDagstqT9n1Dp8zis7BtRgrmcUAA/tlp
bThEsEnwQ7C560+2pnqrVkJOFLwNICgu+Dj/C5OmGq6RBKMSaoHoGBsHh4AcUQ+h
t4PcNufWhrqYOrYII38DIBgFt/RFSGk790MarG347km6F2jTQSyWoWQeD5a/35vm
i/lS+FOodOIVD8hE/9ZAsFhU1UDWQHNJmSuobmIYrWuR4DqDIi+Rr91JfCxvRhyU
F3IGK+evnn1ygaxurJgEkfbrzclBVnO2oXBAHDSKoOvY+iG2o8Avag0xmV57vfK7
2zjMNjkHesPgoQCeJSYXfw0A1WYW07hn6l3Mhtpg6LHtNJzEpzuKl7Jn4M5ngX1+
H36oE5PZ5Y2BSvxWFbWtzkUggMYHm2FqVQm+eSqXIkjz6zft4bcD0zaE+rUVPDIy
PfUWRQOS4eF76cFBVFNKzHyKDeJk2P4S9YzMVWZkjmNj0QfJItQ0da4LqCgRnqXg
M9AG13sXRIvGHnQqmHXXMHVCJ1nwIMifPioJga8IfIhD9gq4BArkyVX0dZObL8ky
J2T9Aq55ho1QTTKxr120iW7cI15TwzoSTM8Iab7ZrhzkUGUfHngXMwongDeIEkh/
coOAMQgv329Hyj0vJyAUh/N6zJB3tZRGOQBl3KeolMbiv91mydupIGiE4r5p8vaS
NQztHXOhs1fOatq/AqRwFBcj1tm5ONZgjfsTyBU4UT6tBc+/xqAvNkuGq38pXRGR
UuVhrBlQxBPwg+KRvh3mXD1KT2ddNluPjEdVXOwCf/bIvwrHuqIX55UF155Mw2Ci
sw+32GM5+oqtOAFqAHm5lRSGUcq8WXtHkWKtn89hYgwV2W7qCEVbXZWSQ67+JhYj
eEbCsbwT523BoqwZda5xeyEHiaaa8o6GRG9HwQkowizEbFZHWgE+6ymyvMVC4n8P
WKUED15BLzkexfhV2IWTUOzvmuM4iO4OMwYkYqn/OsjPH4VJy0qDugDzb7oANvgo
PVyHoR4q6WUPjcaQYLxTdH7u0pDsGByltFrVdemgwdym45Iv1OXSLU4QRYCSacop
I/NTM8KZ2UiKZgHVUwVEFPSz3sha93Zr1goQGhgX43n3hOBC53eMYlwtxmfRGHbW
7Uif/9nwf2MGe1RNS8nEpi9ZmYe2CgRRO7ozs5TBmwkthYp34ZeUmTliFPQ/w7ux
g+hO+0QFXSpn1vsD6rk3eKV22Db8Lw+ZYe8woj83YKFaqDb1DOAaJL6ayD5g3PSV
P6SW+dz5Q+8II4iUONUQus6Jm+tKJzpaAYIz867ko5Df61r/NN+9QF54/z7C1892
biKH0vYfTWs8CnuazBN1dhLRwOg+WiLplJmkGwZ+pvW//HcLLC7rpcI984+hmldv
dONTSLPLuP09FZOalX9nx9by1oiV35NN+AF8LjEZJrAqiy0yOswgCxF8UKYpqepl
5uzcv2r1vONa6TApib5XUhZXFgI9WcI7QlhtGBzISSaSYSgtzxtA16xpfl7gwvfI
07YwkiiCkAooaFEDlKKHgT4+nbAY8MFnJ4ty8IfFWY5R3GUsGfE4Z3Z/BsijMxWb
q8LPcqaLIwGypKdXEmia8M4gp9uw9hOhid6p/VC6D9iEuubEQHZA6GLSs/N0av24
MTud3kt0tq1yT+MKG+1XPi/I7uBahGvrEcACFOb5QVkgAXBb0w+NpnjB0qHKt+hN
VqpdBFXgStz5MOMIVQydgnC0Pgg0JkAqKb6GE2DHsh66AgjjV2MrilF5tv3yNOxp
eGDJ/4eofgfj109p6Of6JSTP8eK6SRI9PkkOUe3+RfWRjymretY/b2fYvZ0DHBfF
jxOLmytpG/FyuDSJ6uNoCIQk9YNBF9ZgXlY/8cMv3f4wb1uSsDCdYXV9WtzIosWt
qYCC0sUQVDblytQC4buM1wU4reVC3eBaLL6NjYfvuXetjxSp3yEhSrZBadr4oVJd
so+8oWML5oxwIBZ85q5+0jSS7OzgCkzVCa5ANBP3gxOSbveu6kt4cr4WT6fr2TGW
tJQqgYsPN079rrCw+6+LbuatRE0KR1h1jvBjnDXvGgiDwMxeeJTImioFhe9UQ+bE
vzq5FCFw6lTNeHtUdDwvonnM3BCsfg7GVLaoFuYOgjRE4sR/o8QzLThpd4RC08/G
42E4YKMtJ7DPF1jJ4sWAJx1PBBI6ll3INf5M07bLvY2N2AudaOpFtwufZKhceb8C
rukSrWgoNJ48M9paiiBVLQbwRdHYEe5mqLRxiUCZOpkKf0UOTzgV5VJsxtuNdPm9
94ZogWiYUT64udnRP45sk1NSEEQiUFFU8jvDy0DRdPM6etdgVdP/9do1tU5M1Lug
XEqhBZ3o+WteyTSJkUtxfHnSkRHd1UROvDY3LugUg7lnLIIVDXEQUeDhx+JIxYy3
Yt5BU8QfjNfYVjFvFW7jdj/gL2YynJaEAzD4IAA2uvDOTf4aq8w4EnPUSYO34zD6
GeAa4kD13/2zVrEyhRTegZ/r9Q5symwSOgFfyvPSxhZzSiEVPtdKeY5wRQAD7Z0W
ag8bMEt6NPuUwKcb9BuJez/laCR25SUb8mrBET1hCqWv8w+z1lUo9JpP8MSnP4ol
sSk4x2ME/MrMKbez3DPuY/0GhmdqdpnhE3nqUYMAmbxnzdG3AtfuNo6a72ZXG5iI
6yVJkxnycBVhz6U/Cd9qHEt5UTpiOYIDfJxVSsNOHDHMhmIYyM2ZSZhKfQKL8GzA
0rdAVDrDY6MviVYjY9DJYVJABTKs/zC9Tqwm6H7RnXqkzpmnHCt/IPSod+EOYGPn
fXc/E3/8vp6JPHTrsVWUEyb3UNWMw7AC3xqSnV6R/wYfVNaWLf+JtB0h5CBZa6Gr
seuSdy/TiL4QXVr5X+2v3SW2d6YsfsFDve7af4GfRNAvYfP0F25mBIKYe8PhhBDm
LnyfGPhv4FRz2OqQLQoTWfJrkwFjdvRtj1Emz/HGig+g/HS9h+JQw7XNbo+3fNgE
OnQOOQWLcCzeUg2Tmk9uSfc4KRxFOVpqAekrB1orRfqeaQh3ItdF9ekSgT3eAAUZ
Nc5jDA/O0aU77HFaBtPIx5qxw6G+1yLoF5JPxDduZfmpAFOWVbIOUgjMhS6Ia5F3
t6lQnlfIEQhRW1JXWgjjeXsEKMCoWOik7yEtdQfID1Gf97YEYEgi7WGqIAEEcAPl
WPpk2kU9MffEZ+xCmgdHn+izTzn6FS5A+X6SjV2WPZC/eSR3g1neL2Bmb32gC4hS
duH6rtesP417HwRZTJxzoyawttC/wU4raLi59xMdZ6PTHc9c5MJ6IDO9tXKCqHdK
dqvof0cMHoUVzGHsm5Px1PRpBHQt0CYqavxHPox+iVj0jvPURlEfGFm/Q2/zoEjJ
AtMrvVBYNnKJm1pwD4zBKHVywT6CI27MY4PCem6M9IDFCFjnc75Y7C3eXysqCzvD
PoesnBRQa8GKKEygRxeRdVu/KNyoUUwJjUJ1p1Aomq/ebgRDEqTNUFzTMtX5vJs9
h/eLumRjlHs5JyMlHlg8tjNJUz1VNM1PNuVJPwWt6yzksbL/NdZXxpVxPTKp7yBJ
uv0sFd2dTAsvXr/EYIwITxpWMABBDGgLecms3MFqiHgw+m4SZE8/Qdz+agf5mssx
TPZxSv75iInIv8Wlq0j+9CkKl/OF2VUR4gP6yv0RiqxfgvFV+RbHBBKu4/My+fO0
teXBiCv1zFWmEGTL2SvgYVlyEVHMqCrpsHx/9nFOoSZR7ffnaJNPm+XnDa9NB2Th
AjFS/1RxTUe/aNokjs9YboEhHT5DJDe7/+IYAulblLZJkFisibOEZU4iUfutwOsf
flL2W6zVI9Sjqsph5FLQmA4Ja3RuFtJ6eRBFLrRLvZjGP4TQywAXZEWgJnKZ0KrJ
P4SVARKxY9CBRr7jQzyP+Mb/Pq3IBKt4JjlUbxWFf+BqA+W6Q3RiXOCGp1TuadZN
vyauraNgxiCRsykgt0z8i/mfVDMWQVkKmMMGpW7x2QpIFxNZltjbamO2bq0lUqdf
0sC/Cc/UO1FFU4eKbuAG6bv4iFZKWakXgWbLC4HBJZayXDML6YYlhJ1RnooJbiiQ
UUQswKVWY6wh0kJ0pdsEJfZG2UVskA8hBtk0kxCQeOUpEONvaQikOLNyHxX/u0bw
3YYvsJggY8unhtwr3BcSm5X7oWZ6h+cwRZMezi+fOlBHR3jJMjKTxDpZtMBU8G1c
s2V3mUTtphY2ZClwDT+EJmV8h+oAVDLD+1sdYiZWS92Ofu2CW44qdJXQSdnlbkRo
JmUHPpwIwBB0QTGI4k6vRD4V2M2KB48qOgbwSYf9YQvSNyQ+JMC4q8rVoW9g0y3W
RxR4X5Ss+8vAjAwaYsGPnWG3U2AVtSp2lKs9qdxrQdMr85Rmhz4UmK80Am+NYMrY
hHUY626kxpMEub1m5DVwVpQH7JbbdhKSflhxv+OUMpxOwimuz1zazbpTXhOuNIyH
uaJvfHD0AkmpnGnZ7L6c8BaWV0kKieVqG90Lpx7+8MkRe9q0/EoucKYWdt7vTnnl
6UDubXyGUgplKkkCzbj1jATCuOPtbTtmwFhXEVmkrFrieRqDb/ZHMWnPvDn/Efsu
SVYiQ1kV0qTmlesQ9XskZ5fysni2Pbh5Ed+LLpeNoGoYhcAyU/Moi6/Shs/MBzvv
rI8GByA1KYKXBLNUAUK7wK3XkNCKSWGvymRvw19IF/kzLRNFWvSIbznineuoeJU6
DoDoka+9ubzy8T+hhZOToGmR5lRjD2jvgKofWwq6QOWA294G5Vu+39hLiTy+C4YD
4tWbeTEF68PtYmp2mm3QjCqF0jtpINOduYfco5xECDAAvzzexz72ioFhWmHX4JmB
sIeT+Gug5au02QXvtphWDFBVpbpKAWFYntywn6xvacefyUW2m2MzPdU7qsxBMy47
/CnZtCDpPcxnZ/atl20PeDVlQfrb+D51i8o9X/VlkKw7l2Nl1xxrkviuwMlVVjVW
7TNKT7Wb2Dh13DfMc/UHyr0fVbIkoUveHUtXjnI8yNcnIpEh2CIuwjcOAC0XQMc2
7ZibKu3ngCQGFXPYghy9AIa1+LD1oCmtl3R5L0Dlo0DPi+hnwb0Kz/xKmsh/eViL
y/lJAnL6QolRQ1/WH5levxS958/DlkHd/E6KyA1VYcC/6qIrhedAkup41mrjMIo9
wxqKdTStbQByzTp1HWzIYQb8ILqYLEXbeQaRH0uClEllo+h+uh3b24BQZNBqSXL8
9invEOJS3oqGw64yF5sA9BCck8KKn0qiAs87w1+DkuJjfrBjFK66UUyJwoiRhhBM
TPdO8LRTWL9Z+G4ohZjXF2QMvC5Ur3WmI2rfju2tM6s0sHkkn2jSsG0X1Uy4OLFr
BtqYheWO03rhtmHbrMqQF7qtVBBfjE/cPbPOruRESRQPlCL5JgfKTmvJSisJg9gj
wCccjHRrfhXpEY4+m1C2TV7RN0xyxgHPtZJsdrfMriHG7Dj4FfrPE+TQDABjmw9y
CrsHGEttPEX7xAvy18x9LmZhpVehmQVaMv2U54iCffpY2AOF/e2YWbYMqvi5Fd8n
5O98PwzWSz4xvSnXDkGxAHANPeOK2FH5yaw3hBt1CitDOyoFOJh1A/qFHWhSiVII
sbkZmrxcB+LQJJnyC/R3R5RpnlAuP+ZWzNm5uxQoYHDCr2mITelpyFB9uHeoI3sD
WxFi+8hxAZWoiET0dyjGLLq0c6VykWtZG7Q6vcCZFe/8Yx5o/acn4I6ihvGnnLwP
rzQFbwwAYHITuDJFNgSWpGZfFsyDudkMk5b99ZtcpuCWKgNuQ9Kzg4Eemo2UU+Vj
yZN7bWG2nqT6gi4b6X6HENGukJhFL+zrYSGqYVJTKraIBW14XdUSQ7m3DR2ypD/F
fYkWri9vOVONtellsZ0Xa9IyHN59V0bH5Qu6u4mWo3fC/VOerVzqI3NHRFr7ailB
vigiU8r1jh4Qy9X3aR8wqGPJOEmXh2P8cnkF0OImf/L6UaY4htneQqECuwu0i5aT
9r2E20dEXGlE6hlrOhDc/d7ESZ4Soue4xSHUN97IlYzqCWsXWn76VwoSMb1LwTGM
Hq76pDmBJ9Nx/+NoUMm+CAM/2R2fgIxfu+I88mJzATkFV6WVaI8/mZGxIntufBp+
94PCV4uPzRTtCB3c/gH5w7N3ASBHeofSNYf4i+rSyrWrosEpK0hlF+4oDY+C8pHw
4b7G/gDwhr+e7tjdYCQP0bLipCoXRFCGoQAr+XoRYp24hiOU7tZ9WOvV6JtatOaK
eJodR2P2uvZ7Tvsrpm3m3Sf77v7J/b6Z4YLk5sgLiCgHGBZuIjG5MD9GX1Onf89J
pIJc+4PrQJ1TRrFEvydqWZRokK38lMwvD8KQS2W6NE/9L65YEiKDJM5Cun5WF629
eFV5HCGYR3QYenU+m1irGYcGrr7XbUrU0WVkf12m4VhKSuVKS5BqxfPGrHixo5Z0
978Blm0G9xfP90Xke7OC6BiwZMonriOWr18KPZiuWVz6o7ns0Dm5kLnU6HkM3b1Z
ZpqsO5zlT89Bqn12poowSe9TCBtjwuMuh4QeI0f+p32692JjelMVLKchKKGyzl1q
44C5FH3JWz+TL9R/YhBlVyp43bAUMUSzOKTu1lvQbmMb/PvBmvOkj+zbdUQcVCzG
CVxzNZQl5AE2IV83sYTn/Yp+GxHZjIIOvEttM/Z3o8WVnbp3v2D6CTDOhd5HBwDk
PGkE4cZO+tDw3xLcAmiS6obLzOs3xt5RKQHkqeenX2+CcUCmeeaHejTYu9PLzT7E
soYTMzpW3XiedEZ7cTcXtgBhXXxTA1iuSkQAEuNr7EN+U7SEhLGeJ/xO4gCdNcKX
Py/b3mKn0/NJSqZKabLZxv2GPGL9SSyL1K9JCgP6WarGvAlilbzU5v+Gbzp8Kr8k
Ti+0IqfanpsnmRxUKYMiYPvlyVsdI6yXG0GCW6dG6HY/N0lqMssRlLUOVH6zdZ0l
ztu+xbMc54BbLksosjuurLJt+Xsdb5Z29sAgNQcEcgxLDt/8pHEoSh9aoFg9tXgO
mAuBKB/WgtyVxmKBhcvgXLkkphh+nt7rsmj5cWYzUqMalsoaQewjg/BpcboZEt1x
TZzOyySdO05rqmpaqDulzE1pfYJdw7XzJe6+tZmzDcYtoh+3HKH2k/MMY+ZRIu4l
bG53MakS3ZR3IKBpjmJaYVSmBJqA9YKthD2C5UHEEa3Ohxy45EqOtNswR9iLH/h+
kl29ZO3esQyTkVlgh6s0g4NKTbATGROEHvrt+pxDifmgY/kSyP2lJmsOtfUQDIYw
xCzJDrSvEt8lBT5NdX9kctWXNjPljQy1Oe0MVe0/yZknreTPjkPHVdqHO7Rci4AK
p2WBA+0HK7qvYRwGmzU7RDytrrlRDSAO8yrO59WZyWQk918q7dpbUEd2mOwEDNJh
zMnLESVTWrR7izDbNXdNvVzKaYna9I3dGB75QG0LDWHgLXsZiasPt4TO3tWA5wC7
funw5+4rGcuSbavFA5mQshaAMzu0dRhLtMd62JtcKNtaAj8d0CEgUVm/Ria4A+iW
8dWo4MVaTEXkVHCdH0Vv5xsiZ7hyCwy0N4YxrE3uM24YfZ+du1mKQ0k1/C4+6pdI
ABunLDxOsvrBf+5FoxIpp3WEJgXvWGZLi3JhpaB02PKYqEkGyesrb1SIWFvKfESF
DM9SPZkZCPSdEPmuJ+TANSNd2QQw6ViAXZat6xR2ZfHQkzFKYQ8BuZfkxIeSWOgk
Vhq558CBa+wmnoub7YmXsqvjzx8ezfxWKOToc/4eY/JScrA6MGOWwm0qYgYn83uO
pED7st5LQfY5RjEff43RY9ddgF3rrqqXzEbwIF86dmfywfXe58orzGkoc1tgfM23
MclvkAC6pgXAGdJ1e3aw/bpPLtVxE4xvnbeID5lpDBH8CacBkJ8oDaC228BKxN2h
iaFsikD8u0BLqs9LIZ/LLm1WH/rfKgqKqBTwMswe0K7NMaVOMz1avdqB/IRL04G/
yQr8lZaHZVEWGmeIEweTF5VZKC/BjUAxzLewmvFn+iO5j+0RarvmeO8sIWXu158N
2R3VT9iw+IUdbmWBgfYBR0SiJC5fiXY/jVARxs3OFv0FKA1jzlO3e5mJxBnAwVkt
pneaaYv3SgEkmvFpG0oBn1CdhAoe9ag5KzYZ3nL4q33R1JWVbrncTDcQVQ5g+YJy
2G7KpbTcv2rceRyrNNRtGkvqlGgIG02lsVdW0n18qkOULVYpgsWgQLpjsJVq42Mm
rQkcXzTkSJzprvfJaLUh794oXv0otzp9El0fOnfum1MqvEAAxppfkV1V2cznZ/sy
SMuuQ64a4DUahBfTwNcXuB01ug3+qd6kXvTJ7PLiSCllnn0Ke4KONrPZGiA3gmnJ
74A1WZGn78wlKtvZCtWV76pyyIM5af5u6STrVKuPwi+iD/ffo5j5h4FqEDd7cC4U
+33jJgPBwqgvWzTRgh4Ni7HoicYmRCPmrvCYvr0viEimUHUVlPSktEc7MUYmUawd
RvP0LhEHA9fXhKYr3ApVJWcJIYnd2I9apWNOwrdkToE1oFKD3+YrvhHSvFznp4QL
gXdxCiDbq21n+dudwpPisL1zUQdVgoesZqFm1BOWITM2cqCUE/nmRQcBUDex9li6
RfEPT5Am0tZ4L31vIjSEbY/DQuD74DmgNzvL07axSd8U4r1UHoVZENZ6WVQJDzXT
eC+3GYrSGVPTE/IIpi2bFruJfaT3fTPtCk13GeZeRsrhbvNlsuk2HtL6kxn1RILL
JIGDNtsb2IJk88PHqCqCUftSiUVfpiUMD5yQk8HNxaZl1Y8CETZ2G2lL3RdWUDyG
QOrA6pvJSkAPglmkwhByMtW7i4aOO3OL/STZd7bp0jcMbEu3BGz0KA4H/ODXrnMZ
RZXf2vUgaILPf7ssnUkhZEertPpuLDI6Ne9wjV94kDN8h8BF+aHUzgrVeANPNoYc
nE/ludkYmmk+wj47/Fp45xwSndt+cUQ6ykbpDibN3LG+y3i6/gCWRGoWLbMNSCwU
YSgA9xHPTJNNO1Qe2d68K99Wv9eGAUPz+xcGGNNrv2slmbPXVGBia5TXIc+Py96B
mgEyH0wKC8UK0ExJa9n5x8R6gi7W+gR/MXKOQQ2BHq7oFW+FwkoKPlbWMVXV/MxI
KFzPsQppP6tukoSfa7Uqmg/dRlxMQe6qNj/SMPUxs7pf+qF3OQiTVHkAbCuP3s9e
IOO7MSKw4I3NRbxSh+gRSFdQDUCNWjMxOuXVe9UojOhXxcsdtgzha+rVTHwa/IQN
NB30DjJPJK2IK3Sx/4p7Jm3zCOJ+i9VJytq0a3r4i7hYxhXrPuM1hk0AhNJafUy/
DvDMe8EyEHsAGBbrQzLDL3cK9r7tG/yIaKKT79A5IKNrwhSIlh1cpUVUemhIlDHb
mtaH87+8/pJ7/LerKtsbrTbFagm263DoNtGrw8psdR12whar+VNJTakLgTtQrGIT
ccSkJ/9h2BXOuZe60TFJzo1Sq4CNPTQPE3MvWHqKC0xUSPZ0aRPn+zyameBoOFVS
S6wbr0W4YQAyCa3lzzocGsB2X8ZNnYflWuP+HOU/LGNJGZqc49rny4Lz85Xd5L/A
m/9cxf3qqIWBY1Gjy3v86r77Xg4zWebpHWnq4g58JdttAdibrUQyHhI8VYircT1B
mIEMKZW++TEo2XZhP1oEUJyort22Y+3Xx9rN5UwXqYUt06W2WpOxBkN6wcwTOtzI
/y+K3ilwq+eVg5dlu8CIEcXaOQ7nh8tjG2bOHLASiLcEzFG8ZK4tjaMToiZrM/a8
0p3+FPlg74AyTtj8y+ao0sZp36RV8mTdqCE9lB/CNJ3TVRWFdaUF2kOTzJ6TPXI3
7hhsIjjehNlGHtGc+HtdRJW3Jdb3WZLqdq9RrP2AEwgrn9A4QCg7b5/dFP3Q4/t1
wqW6X8IyWqKwg5I2YS7iIOU3DDYygCS21cjdD4O0rQcLNdzSdm8MkJnIS1UD6NMS
b3espRvgnmMJckRLApkZS43n2WDHHBItVo1nXrT2eqDdRbadsgg/xp3XS2O152UX
oCac8vN495ki3ndhQ3LROW1rmgsklXL5EyNr9XXyn46XyD7y0EOeHNiZcNylIOTj
2zzthfQIxLYgDbtNP5hs6KOywIOY7C4BFhe1xnCQijXqJ8U+NyCHe6W0Tnfx/5D6
jE6axsqrEbjhNKnYnzTEN7t9fhDcVbXEBmSMAGvz0HJBjvzSZj65OLozJw5xFHr+
rMSsU+nTJSUJ7TMbOXlWtzhv6LS5lLxKRFsm0P7wQLzle7fMnitInOqE6SP7R3r9
OCtOQfrTLDJ+WyTSGm1vlX81Z5V8B0OQ4GxMPzoKVPie05HFvM5zOLZbApMX65ro
sshg0bjAFnjaZjID4KMIU5BO5BXFnI8wIJwC8MOXIliYyQZReyqkQ4F5zeDCpI8X
5ckths80P6WvQ+huPT3kgdlVchbqZCAeTODqo0d9i5FQXcKO+Q6r/1tTJJEc9GOD
F/yX4SraiGpL16QLvFc+YC94n4oQR+Ms3nJSP++I4ckNbWe4vmdth4v7q1V7b/1g
+e8q2ZhmJkQJ0jROodWN3UWzu/FLHY+vdO50zarSBnsf7OTNYBuxzu35MCJT1KP7
GahAMq3MQ84mQPPOxPniu+IiuSvLI4VX6ctg5K2DKPwCYJxPc1V0idUsaNfTU8d0
srAmhxdQFhIztkyq/BGV61hiNQkfzcChqxc5SSj1L/qBdrqzyQ3fBfgnlfPqArFC
zoOBPKpJubL7OxEOcDnPJvk5OX6O8iRDBuJNX4clAXSy+UnWKblSX8WjjUVTzXgc
8GNDFltjb8h8w3duVFs4jrrb9v1gZfoCBxaMjYl/fhgpFq2oV8SxzvQ2tWM8rDag
uVAc+u+r4S7BW4R/YON4r4QBH7mG5WU64rfrdE0EQjnghQfc+/+L/hhukkqCSkjo
h4q8oZMjUlcuB26jIczjOAkFNPsDSbkHpLNPcY9oCEpuifrrH9RMTX1iKBtJqgw/
yIVVghw0BPbCOazEYpNupDwHp/m9n92AAjbAAndlFfNQtLVAijWENQG+aEBKW57i
K6Kfa/trdWhWdpSV//agLmJj7DWORZ8k95X0VuwiOXSHBHjTEZrnokZhenV68S0X
e6sXjsONbg0yvMxmMlXdsy1FUGNohDqGvmCxg3r8xhXHdalD2B0TBLwnE15PT0bD
dwvZoP4Pt9YfROl9Pza5U3jWRPPRtSKl2TOy63GWx+vhHzLXIAPAnV1XUw9BF5z5
qwTpnkobaiTW333pF3Dbv0pMglhu5zx67V06NZ07lYqfC3PqD3Jmbi/g7sIXi7On
mtLWpuRihpgKJW5QKqhAEl7aF/EE+jwRqE8xh91OHjwLDlBcBTRpKDVmdiYryScK
84iwXHYjau0pWiUKd4xnUmdlGAfZ1ysIw1uAqeHzbkfBVGJ4WbOGl3iysDVBlp7S
Xa/hJUryqOxkCEcfJjA9+gAQCUGVUnCkWkD7mptiOGWoTVabaMD63gDFQqmvhLkR
Hp9aZPBvQDfbd6EQRpenPRwMSoqByYLDSHSS21DrMF8yDjkr3T6W+JpcDEHOzAfx
qehzUMQCIyBJzOeBhcGARKyI8WXQ2NxRRvl6gkmebVz5nCU0P68LCZF5JcoqTWtv
nJIp2Kq3w44WKJ0Vnb6R94yQQgJI13rMrqg8lDgibnZqY1/2dB0eJz8TIM7DrpxW
oRC7Nx5HhKizWrlishUqIoylVyXVWmiB+bsjejG/djJPfqiAerH8QaYoRZGHHFGy
JjdqZ3TFz0FQ3UpfMM11CZamvrEeKBnRSScO/VmfuH5z0sQJaZ5AhG34LwTYC3vc
a0d0nyHOo51t9vyGbsAbc9HIy2Q1EFEB5pxHj/Z0yk3k6UVyuBo5lsa7McXj/1dL
vQabckzF9xMRxCoMezrNnsbDMmb4aCyExvZsi87VswoY/2v19pkCstzA3P60DV/D
aV572hOeKGJ/99ocW0Anm3L54VFJb77ZnjnyhVXH3by/WBRou7rcHU4q7dh8CETK
ZdVRRbJ9G2nYy0DswpRmG6YNOhm0vP0S2JoUHoCuKGAaJnPdEgkUIKlA3/IowEps
39VJMu89xKoBHl9SDeTjptl6g5beyf2Eoko5DG+K3WTx06eb+Ex7jrFzGqpCe590
UDMcQpNiXFpRdPCtUOVJNlIDO1afrS0Sv1iLXB5GdhzcCLJucDld7syv6Wy2SdBz
Dz6zI3UofpO6pILPhiGd50iT9LCM6Js+3TGOfFGCT/JPAatM4ID1gU3hiIO2akDP
nacuUS0Y73XPAcyes3Ff5L0vftvIcAfaGPJtqTbNX5XKUDNLf6PL3ym0Qept8hmS
bnn/+FlX7s+amdH59oSzEQimUE4Ow/LjjMVYtJJom5HeBnS2FCgEhtocrVt3eo9n
E7qC8kH5NTKAmPe6PlJl880ME5wmqe9ZaXZO8ePueq2tKWxg1AlE5Cq/Zii89TwI
lBh5egYmhYnhiupTp7WZCTGvfZZZZpQzcHKhcvns5oWmZTBLfFAcIqiK+r1e0312
3BPoKguVEqCLYljKrzOUEmAcskGGZQyVXB0FVrIrlP8Dji4sKG0O/Ca1S3tDAbyA
bHFQ0u5Uni3gutYXL3zt2bWl1RviNVvJBR3+EczXJfxNa5wlJ32jYIgipK4MmqRT
gaKkR0mkBc7eIPFILmDGeWlxTZ1NL3aRwfpUisuVDxJMU62izA9O9zl2VkufSzoq
1LSdLlHfVd+Kr+UTTWeW9sRqOcMO54XmA4DlzO+gNDIG+FrM5izJCq3dSlwt2MrT
p3h3tWxSLdcdqDjbCQT7/xk/rO3ZmKKCTWN0XAq1/ft8EPsP7OKV8qxFhN7Kp5ri
Gz1w65/Z14SkE7BGGvksNhvKzVdzI2eVH75y7RY1kTs+dKIj2ktIUWgboSRtJKhL
I71imzCZpc8qWAs5UjT9k+4NTQuPY0hx72GFQm0sTkzZ+2oteuWv7jJnGRDErW7j
IgCZpO4V4IsUftwfVzAt7kAy2Dt0kHUIxLwXEHzxh/CUl5E9E44xpnRK7jMpRbQG
OcIw24Mk5fiB2Tg65j75q94/mBvagyZg3Bo69k3TCCJhdpKIQqphV39ypefT8gvo
JrHztghZm7cchIMO5dbC3H0DxAHv8oUUGhdfptIS1aqI2e4C0EE+5RCWifXgzjgf
bNz/DuvChSkP5gpKyeBf57akf+Z26CeFOYE55SZ/EXQnfum/GRsgJq3MHtOqNrxt
ZSCjzKQI5TMmDMRXzhwQGxeRg5pHP7vdu+hZNup5m9cH9RlFonH21sxI7asIlbKJ
GcesEesoDo3MnzxV16e+kPuPPS08vbrkA+GtmSPK1LSEIEkzIpwuC8wLc+9H6ZXE
W6ZqhR0v2KLtXslOJ9vNIci0ajzSkWyBtI2HJxVLdN/DpO/60rdEgBlZBRphxi0S
0z3O68aY9x6IkroVHtLjtzUmJrGOFe1VBSyMEwvCwJMJ7tOKM6Yi4XmUALbIwN5Z
5Vkf0qEoVbK6MjVtZ7a3F6RdIU+WFy9d5ShER39caKGAeVzlkkmwo2JZPDwnY7r2
KRaOAKRxCtBF9draw95SeR4eKjoCji5BuBXxLOS14X+b3LaN69M2yhLUAxzDxiaI
nmm33xnPnBKY9WPhgL3PwuIPPc0vcL5JtAn3ZjPb8LnWuPSrlIuRCeHBogvz1DVO
lnwk9L86WNF5Emi4eDwRYpnHVfAGOUMBykDURjDs1LRfZZyzRwN8nwnCzHnVCD/T
wlWB1MrebAUFxXDCwxxYzhKnQA40VAhHqzKdBm0XgDi6d3Z0iR7FTU6fOE5zQKNZ
+2zb22xfXByrEMnAtMQAo39d8cBxHNnqaC1RH586IrLr3p4W2etDZRnqO9z0AHnZ
Ocy16Cg+G/k4FECsJG27daVfusKCcEPDEKYX9NvfxCoJowwiygiUba8+X7pPcMHs
jEoUZXSQo9X2FKXP42kF+avXCW5Ixerpd+u0aUbjlvAZTFwknHHxewjFNXSlclel
fcsKvsUV5uq40z5lvVVpmH5kux7IsikXwxE0FCfplvUuNiVwZiMJkdywpHuuVldN
Cik8HlyxxfwLNl8hdEoURwIgrLdL2TbFW3sHNpsjOzDkDoWWU0eOiqIpmi+qsWXl
jMXuL30eekITi5WAq1HVqmUNuf7Cg3pIitBYAIVvZK1WqTuK870e7c8cAtZfOB3x
48PyppBwyhBSBFJARYjrlde8/ZYZo5RujWK5C1lXdDISrGuyQlueVDvi5P7irjS/
PI5AKAwXmQv2lnVzKyyX6EYND7R5/XjIbI5NAz+EgF2j3LgZiJKdRMVQ3fs0yGlR
iZqqokXDZ0UuAoSm/gpirp7g65ZLWpNgbJwgPm+mNJoKG/l4AndCHHnbjZkMITyU
k7tM740iXGWRBMxGDaprw1ApIcJWXb+Rs3TRp8q+29/JqG2VQ2HvNEpBHG9lF92J
+PaLYrLam+fsStqnA/6AImL0PPLQt+tY/PZ+Emr4XFUR/Yw2qNvune+23Attr/jk
T0FJTbgsaMPgywoo742Q6i8tBJYHhkfCrd0itndhVe8G0FG/B55D0OeQKh1yWU1S
IqP/0gTEIAtRd+25J00bMz2pb8YoGYU2CWfDPfTtj5n8SOzrbBoSEtFTX4/TfQSS
uNI1RObugI+7fnROlnrIdeQqetTawCOed3gfJ5yZa0ahigv/7gOPvwKbtH8yaJ9J
giWsaSpWZNv5tGoJMuH52DA0KHwpeLfPX5IMHK3Mw304NFAe5ii9wCN3dPq3K0Fp
00RZRQu0/VfWBB3j9NHkMf8t1CXaNAWgxisG58HMBFO8Iksjq++LuPXjGfb7AUGl
vgnHGViR8y06VgqbBGN2vEU6wTLc5zWzVJgnFQRD7MIi6ydfhFhk/cffpBZZAIU8
xK+QEHID+kRIY0MEUXd/L17IK9IPvUYU2V6emiPl/uRTewhtRI+5J2KxPtr3tWKb
sPfF4orvUnsL6xrt4d2NxbVxxSwsofdOz7RfVEZw8qnlv1/CKUNSnR2TN9gclsNg
J+IaB1hiUFTvKsjXpt/Gm/lJWOUmElTvDBXv1zi5ZLThfNrFd/axXlrJtTb7vIV0
8F2hx9CcAgAoAy7+Ot6eGcxtbS2ligUyEwNJeRFlDOp/5L5PYU5FV4U9y1+UoRkk
5YfXerbJnw/wSPKo4eovpMha2DvSKb+vzfKCkWgmno/k/7OdzYeKM+SSfMFXB1EC
qELFC7IS0COzvu11b3wArybSea5xBypioeEoReRTITYMhUumv1C8zNqO8paAvfyw
qPhY9dIYdpsUWDbeMdIZs0dDtLLXfmrVUHw3/Ev9CEojbosm8C8LNM79C+dkusPQ
3M3NBT9dKIE+AauBF2gJfFkmtIj/FXY2TPwGlJ9TqLc0Dve5/001JEbogVqMuJBW
OM4Zrhy1IN/bJ5JbOwMk2dd8Du1305RrE7L55kkm7jmdKuqOqHqNvo3xldlxSNjj
Jd6aPRNgcvVNXNSG5AkxZ4t5H/mB0MAjGEPrXNSE+t1XyPrS0Y002sjC3z7mizS+
8/ufVRxMijE3KHckbjlKRNS7jgp75PRdu3qZR5rZJrVTbF65B7ow00mhzKM5DVkX
mEqO9LgJDmDhUjlTnLSF7RGTFzKyl3a9CotHnEwbkrX33YjOYoV6XHr3iIInFhd6
woGFj7kqfmTjU+oZug/eI1YXtlA6DNMvIuVR7Wb1g5VRoL3+pSOYcwQxkXvrsiGJ
yQ0cuNN7zgqApraOZSLnLNY9eJoT63ZfUUiuXbfParyLyclNpduXkXWcPGbSLgf3
2m2tUEDlJ3ov0302hJruDXzKYDJ2VBeKz8oW36yPJdPwCzRM696PHwYLGZmEABW1
l2dny0SyVLirPpV2ENFw0kyHfxsNz5rhLlmp9seVsoDMcsJS523RlVkEnFi1I/uN
k+COr+SIZ+N6SL3wFekJA1n2SJQ9/uFaqx6VS3Wjc+Z2AfQuN5XnxqcVA6Xsk3fy
xoZFoh8eoKXYXbpO5eDKFQJF/hfXg8kpmxpA7l/cdV3RhU0oDdcrJoGmEZOX+tHG
Lf4mTShLqNgO1wkmtgViDK4hwCWSdu2m8UIsvTNNq50dhJtaErv3Xoh3K3oi3+zg
IPr8uNp+0Mat+RTgu9+OJNvQ2uruF55J6Y8m5poxevD5yne/N517LYEAn5g9Gzzx
0EA9VnIG4ZD5VYUl8UsMgnGnxhr4+VBI+BC3XNiek02L65tq12FDXAV8YIOJO/6P
34mYj5ZfafjeAfeJNBHOYwZPItv/YhTbcXA8X/pXPaabUPI4kLLapxf6lnCpbI+A
RCw1GI+6youo0nm8a9AnwMm+XKHh7V4q0oiTaKcXiegTKB9xqQyFaxqI0s9Oxcnn
po3RmeupeJnVqPBpl3blX3ZvDU6cXYajjuaX7Ra1BicvixcYAJCdt18tNYPSTP0t
fbOHpnBHxZShUlF+oWgx3LPXmr2JIGhz3iUNyu9KOAIXNz+Nbn1IhYJ9Bk/9OrkA
Hkhg7HLMBbUKm4h+EHovHl1ytSkZ2bmBScJVvRmx3It+SMmuFXnfMB2+hmQckXZo
Ihmtx6IwA9L0ba8kG5mex6sL69kkfFDG8niiIl+BDbnd2I6yertKFq/NiR+VyLQy
3xMaemH4Vs2TM9sAJRrvNza2PInNauGI0iWMKV/FIcy/XfBDFq17qzvXiAdyBFCD
FNCidHZEvL9rsgVu3BSYXzBH7K7JWPcWpsjPNqmOLXBlkpN4hogaAbnbcrVCL7qv
CA0nxzbuoN3r3V2KdmUiBdHytrover3GnxaYdDd6plnfJ+IkFWNw3c3nb2Waeis5
5HWkT/n/tf11dsvIHffR4w8Maobaz2/0dJ48dvHPpAmbjB8I2HsIMaHrS/6WTOL7
NAwhXZWrT5cOLVJDxgSOodhos9VQKjKgicq5Ga+vpFOjP27g5GPa1vfe/tNeoOdH
2sHjpyEiRProTu0cyEVUiQZUjlsCh/H6uZVGUQziadbNjPtMJinM1B0CV9nMkLg6
jXxulHmpxEtJg+mEsLT1ir6I/sl55JRJDNp9ny4kI3uZ2N9KY2DOaRvF+g7hiMRa
pnWSiZ9XPbOdZOs6nPI4hDlREnd7P3uZ+5xdX0rqlQfMN5zL2pixFwV+W3XmVZ92
4KFaQtwJ0ARrrxuvp2c7uYgd23hIM5ERtIfq7IAcGaoCuuuUxUVE0A9fPXl5raws
7vrb06Y+C66TP5kphP+maJA7W0M1ofD0ndRpU4m/LE2kCQNEnHMr9XgBJ5ubWCFp
KK1dTJdlXLJ4CNXQKT0W3kQeQUN96SQJrEh67Is+8wA8iu8rabY7zWNCX+RMBAL6
7TC0fq5dReuRJ1jZIIZxhN7O0og28ZxenjJXi+AJZPad0A1QtnTeGtu3DvwDJ+9E
M961hcKDUwFvjxCdI+oCrEvf4tPOzbzSu1y9HPEbsheh7HEfp3iJuSgIrM3Qh6g6
1YKRPGs2cx0n4CCFh9+IRef/Co2sox1Z9vyS7AbT1za7RU1diW4tnMg0uq3h6f+/
5fKYq32O/ztMnS3wfRQn3z/Ko7oHgxMZT3la9yCSDTcWS2vdQHi/pqbUDlA6p52c
h3zN8RmBwOWOqRE5tDVNxgbZfr1Z0kY87aEHlgUgdyPaqyRpkzA2PfSFrkfu6hVd
hfRlWiCKUUEDUz/BIXefdhGoTJr/4cPEvt7VJPqNXVqNHTuFch6LfZxsXVuiSiOJ
DnSUekXMMNWOoWLhvmUImmEq/4mcIkvL9mGMQoTZ67YlYBb5ljnIBDQ+0qmeIi2L
3lbB+BZb/TcXhaHWMS6Ei+nqHrj4pfv9V7BB3tnePr27O8bJoZ0MBW7IUbmlnuXo
Y1LeERQ6ff9QJ6UakV2cG17d2/gwhvq0KHxiPio++GI47P4WAyzpEPeX1qoQ6OGz
5T1W+gbAShq9WCfpS2bMkFSOfnVH3akmClyVqQxAiT7Rto+QKV17zmYvF+AOeNlZ
Fx3rHuFQQ2pTLo3K242E16rXiXMKUZo9PqU7wqyRmjIJLxv39yw47Y/fn311MY5S
aPT1TTkw9RfD72mLYwlbYNhyQ2np3odprM3BA9B+DvhV0McMQYZySY9DEC20soQD
7Y+TOePTiI4qsXvFeWm+dB9kzfgLfIMVGYur6G1eb6hSLx8hE1GwV+YNAV39QAfw
10208Fi/5Eh8a1RaZq8m0BDb2XjHSE9QTgXFZfEJgSYl15uRzUMokUbxg/faqmlS
dNWMFbeQlgVjZC0u4Tx9dLVzU2nXicGho/8KphVQS0oz8llW3gD+4GesM+y7Zz8F
Jyxk8kYHu6nmAQnMqs5PuOK9k9voTkFafqPnmsAVLGD101a1i8Z2u1PcilJWhFHV
IqJ72K1qjfZc9z0Dd8nlOqaVcpxgp8HQU6gzEQ/WoQDbnbUuQE18oS7K2Mar+3zj
kfmuUcJVTGAwK7Ldc40km7Aj2iOaHjdwaat7GQq9BAqvDmdyPlHj7SJi1I29HkG8
O3cEbGVvxyPAb0v4lSz4iD3wnbuEm6lwABypZj6lsYCArGHUOM2MDgXns4nd5gBB
jbQP/Cfmu1sAFaTIpME/Fp0TRv3LGvNvUkbOazCQnPCx2mgK9eO8I+Pyad9c28T8
cgpNnMMW5+vOPsAkCCVZV13yxnDMw67X8t/u0V/iSRwc/3VhaltuUY/IznQYwhLd
xw1q4BvZBzlG3wnL3mMTdZKq2qUNS20H5JYvgHDGP22eNWCFxXl3v/uuLEoEGSq1
aY8rSWXiheWAAKDSvYW5CDxXRNZqi7p4OGRFRZo1Ssj3Bgj2W3l05FiMK6m83KKq
nVBe/A32seeEOynQm974ryljcgNaOFcpwLrc3VLXAFj8hXL0aLanni11Rdmzx3ID
yDLt/HkA2KqbKvXGaeKke3lGYeGM8pLikflh3fSgl0p3ih3O+VBNKZ+lPukic1Ot
EtbPSV3db2daEcf0dAJOEr7SNVAwU2o52lXl7/CPP30MEqmye9p3eXhLt0SMc9yy
FVzm+BwSZ0bknSz/30qJIlJetS4liOPZV8aITpcPN6WJdW/TD7qKaMDxN43Aybyn
p0uTGZeD13TDzQBTHo8SMNEJ//Um1KjxVX0p4K7ONicULjBGcfv99lcC/HJaUiBK
uoHHZ0nv/LE7v+4XNKnAa1B2Uhw8dBYNDn33Twpj5bKkeacVD5Be3IjkXEA2i0QL
6z+JFLB+KB5jKNGf6AILuJu7jjWHs5NsEOTTMrAA7Sbv1x4VPGKYUYEokLvgSJiN
KpEXJmOYJp+0zuEmE2meDZ6PxgZZwBz8aunExI0GfmkUWrMLME60eOOMUcquWSdN
9ZXKbnbfI4ltknQC+J++kI72M3rd5JYsqth1SPvswFOt1ROXgt4V2emZLDfUMesW
dhYr+tQPonui67bbXarM5PoOsGkhyy2FCHywNBonSmqqWKhHlwZtyYZMr6IM/Peh
N9U1Nj5GBxeXJ8LN0OaQDemAPl6PyDhxoHp6YAee2QaCpcSMYequ8vrH16zI9E8j
JCZSDZOaJdjibF5hhibHxMKSPl8KXjItQYDSUO66Ju/SmlD54ADtHSS/BKUj3z0p
K8RaJOPmhuiFDUOeQ7EavRbZKjo33/YruME5IeI7aBWCw76pCwcp/56sa8V81orJ
tZpKjWw5MSv82FAvcgRrcwI6Ro8VFDkzP1is3XYar0iPQFSvM4VMfAZUPXGwP33s
FWuGNOTGd6kGFB33vMRFta8Y76J+UnL2rmZJFeccjmJS5nEZ2js/JyuFwMS3cmLl
iyfWxZTUfXp+U8t+JDqWM9nWGb7AD64FEq7TqhgTo3gkn4cuTZRdnTIJXS31OeCA
fMQ41vhnYpBCIgbV7KJxfh1RXEKyZKTd20vPVCG2Q3jXXtvIurYEQyt4dbRUvdaR
9dYsEY3vwOXvRAvj1Q8p9U7XU/8e2alfeZC8loGsNfr4+lGgPnr6wQ3omgOeYdzQ
5lZGfCyBwfTCxhuh4fLfeQQWej+NSy3aomzDi9yFuCp9X6uRm7EGmU36QP/Fa4FR
L1hck96tFje7sm6lPiMxIzmLpYldenN5oLixPCu7W6VgUjocn8vMw9kZXhvV+EOH
NbHmENEKKubXKcIsTsmsxgSEqcnl9uq67SjG3fe7rlK5i8/YxdPZiyUJR4zC6877
MXlQJjF1MPHVCXiR3sX5+GcqBigMTACdTN8J6UE4cGZ0CSHLgyooLAHl3tB4WqwR
22evyzgafS/HujgAUBxuYKLEipsImadzYgKpkthxC9HyVl9wqvRkOCtCaEOZlAXJ
TNIvSrKQ6t2jF7nnN0mZTzUxrO6+q6Ks2m461F4vzl2i8iK/tIg3O7dkousjMszu
Wdr6MkGtwAI6pDSXFxCOMKZclU9MIxICK7nSaGe/sg3ix2JbV/HBd8NepCX6Bh5K
0rX1pZg8HlbefY+nX/ehbJxeFmU/xnZsWWWL5ireDGde09l+kVJKHmNcFS64biD0
I4HrqXcHTvB80NdlD+G9lP40r27FlzfAVoqUm5qUfoDWfgpf42p72Smi3LrPAFD8
tShei3zYTSyBlMf8MaXsmv/hc70fR4SW/I6MYOhHn8mnj0ADsYGqVBIvrh8Ql0MX
Ve14tAofbGlH2Sr32E+oZCOEJ57d7tNvz5JT4QLAVxqHy2Ts41hBTdPzxz8aNB+R
2oTfYg/X+CIFeTWQ4d6DVAh9+Tw9JGp+v/jYZM69Wlr1thPjapVGuloD+BcWv4O2
0yOxqwe20oN48tK1dGn7H25pFbtJH5i1/2NzFU+Losv8rVdewI3ulKiegb0rXLEQ
7ae9JRRBGofLuSmrt5WDbdlrGiWF73XcL5X8OJnSpyW5/04HTZvfgkgQeD78WfEa
WHOP0SydFroDlnbjKZQxvc2Jk/qlwlLrQAz+3hY5YkR0bCocdSWkBHz6KHPU1jel
Bs/ARGi04yy+a5qpwu3JBl/JAPmgj1+gY4PlWx3ubJoN+WKsnNtSqhkRDQqddqgv
Uv4qcIEGdW3K2WCRTFwPpNvktkBYbJa6srqOK62uvQRztWxnCnfJbZoFZxlnCIiH
2+dvKJsrT4S1cJiM3fHYVeOADj0epwCCzuC95BD2xCKHzaN7VchPe28ql9uC47fQ
Cr7f9WOugYt12pt5+3CA78KHY/HtReO+n0RWqYc9KCj6zapk4Zzr9irgHkhbjNoE
nR02PwH+C6q4mpmXcMjTxeiflnm6+Fv4yojXrowi2JAHBAQrb2hvn4X+NMAenRq8
vwDwOSRCAQJ+hgiF4O1JXFArJlGnAR4LdElR9dUo3JVW+yDda8rgrFyO6Qf5Frqi
tMhTFvRfPXR+W+eSHpGedVT97X6/Two73drVyI5hgbjiNrW/lqMCh0Xd1ShFpPRV
8bwedJUYgGD8LmFiTzdiwVcZQXivknnI7XLiXwxmOg6ekYGkky0EqiXFbuWLaqcj
qhi46qOKDGT5+a2S1hf30Ea/9kl3HcuOoVzyRWuHrYxEerpPyXLuoLDacISGGhP1
WeYHsvmubKzcdF0pxU6hK95jq62JHchY6yIBvn5E6SnO2JWQXQLh8SbYVRgT8nVc
Ef1Ef5jB/O6oRt48QS7tGP/CdgumO3DSMdvvBDfl65NKt/1XLGr00s6If1B2eioL
kqodlUFP5fMsmBufJyegB/orHBq+Ni56Wz7EU4BZ7NciZhqLloWxnMGEfQLr8g54
/kpjOhrQiVfZvJ4JlxV/QyNcouKte9AWwZufRymfBJlGR5HSjtg0a51Wuri2ikUW
ETYvETiRp60ilTzdMxF7ASY8cfWMg6QEpk/Kj1CYGKps5N4AL52XAYfY79dNdk3U
pqo+dikTxIX9qSeREmQkQ/pdzv0suoMt51MExTBEAravj0y6qbCbHae5wYGxa4vC
+ZtOpzuFMQaylYWDE/wZhagB9jRdsx0+DtOmJ08hyOK8gmyjSYb9oJ2RjW+OJChp
5QVDP2hWuwvHtTDDHwyBId3fOOsehBwGqx5iFFd+KpVcTXB55hJdd7GDnp2LzW8/
30zHJmMFHg7A0wzpdjbhxXDdqH+mRTEH7HUxk0bQQM0l34a7cztLVEV567B5jmJy
0/PMdIG9ZYeL9xXXHitq69SCSyk67BZjvFAjht0EmGR7J6B2pJKrMyrUMYGOqoP/
qXCKfKZa+q1BMaCPQn2wgz1mjsvvXcajAK80Ij9JSgIKfoeUZQfXj6Uz1S+VD/x+
P9/nOeNU5dB6Z0HM6AJEcWslpmMaxyyohYe5qzCIIVpAQa5yxVNIgSEbhxIzkaob
LRIq6nIlQuVSIfXyUeHdS1/83eNedEAi6Vej3FcRZo+r5v2BaAYtj+zp1aWdd9wR
inhziTOXq/BMp5pwZuHHxuckJcQBB0WQVwFgpKXi7vmo6d3qiJpJ6OmhiFCw6EQ1
6IRgZMdX8722iuupyeomVh8OtsXXxg2sJHGMdNJcOl3tlURMQi0efV+0Hu1xAm72
UK+MtFm59m64wfhwTEAMlFa5KzpOgvteku03hVLmAFywlmEpOUjbvvQJwxwzRAtk
I10pv0acIksTauhl6bHFnMRcotYLpJy2BDxbJT4HRUqb72vwcc72bjTzjqWtDqxE
25ih1cenDK7RKaVPMKfvbgYlBbCWQG6CQrjhPkZw2V3xEn3i9oN3HCeJ8TlRP5BY
15lwwAI7FgYVGR/UjVCme1HpDS69SJutepSu0NSIpQBjIoKwuOfv74w4iKoWL0qc
CSnXE+rYrMIB3BEJy9+VvpPXSa+zGeqtuV5p0yO3n9ifxpslailIDTLOw6IfKydQ
VvacRNqS58w0Y56hhe+347KQ6VLT+G+GcyK8uTrZOfYeDXazeCMwLdvTV8c0T8Df
yPI1iD4Rcfr7d3EYY+wbPKMtljxlyNswKRTWucRc3SIIM9WZXJNqhZdOTZXn6n3C
Q6gYR8wFQnu9pyriu/8PfpnpsyhQ6z3Y/baKolY6QbpU3wN+t4OMEPzFY2Bs86Dc
1aLaQA9d5Zfa+nMiD1nwU+1vFm5X8mb08bbVGtmKrGjK/ciGLTCKpn/WILkIIo2q
2V6nVuKNgrNozldZSCP2s54gLNTWiCzrf5/0tU3dreedwp9TFfzt8B/ZgEWWNU8M
BD84Wliv5A4ruzlGN0tEgA813iFyRZlx8SFXHCeyhSsdLwSqzmBctbMl5XT/SVuA
dB2MdT9DcH0FggWfr5wUSZLkR08HJkBnKI/mXy5p6owG2yYjL5tBW/WtYwwg+LJa
hj7yLugFiLHGGiejDledXnlOur3B9KwLtSCzb7nt528MRUvBYVazf09yvCBU7TaN
9LzbPA4iz3bEz6ACyM0XsDsTkh0ZgV6tYjZlWj4bLXbx+DoDd3FJ0ZQb5/Mmin1k
VL02efBwT+rT7lRertBiX7XYSw3bHS6RLYKqmgF0q8kvL4RzX615RcON6hNh3wQl
hLlVuX2z+LXZ615Axsnex0nLzyVHSuwAaKLIpJ5fXZZO9VNjeituFxtHMI6bW5DM
mHEfkKLbbgMXy9IMQVSEF5rO+xmiJ9phvAroBsIA4Wm1YvdqMCosQpTPLfyybsgu
6FoFB4pYnO78x+zj1oEhc804Pe+3TKiNrtb9lIAWWo7wPNh1NsFrGVwRSYEEt041
bu/zDNCSyjmRo0ZUB9ooEeDiiDHk7Va42MvTtbnkN4yv3VNmDSsyc+lSw2NALmF2
FkUl8CCrYwF3X0dHa76INunkBNkyOP4MJ9TxXr4MbtXh6qMzmBFAh45PI0zJ5qeu
yX+rvHHn6tnWpNkV5a0Y/LafCerH0zweQaEwGftE/TMI0vNQWDbJg4HA+Fklm7fE
J4zrs0Bjlk13nlMmVoT+kakqHws9B+B3bZ/ouBkgW40cRrXHPGdIWpryon8NiHNf
qYf1dCWCzB+XzjOWv1vZseIjKP3rDvQG7Bqq3wEmQ8fn7gh6I31nwIG1lZ0ZQSHW
G9arGJRfGpHxHxvUK4S5nlcQl03n2w/V6pvkXMI/qFsJ4DO4vXA1CGINnqugYgZg
sbGSSpM8u9lpCBfNtc7fyzo/qYrO96bLwOB7ALgTAsPGhl/lHCwJEf/bO5lQ4lxo
XJhWbJzO7SRD7AAsl9S2VrWH63VeLR3EEx3F8PYFqhOxlFbeTTafl2Cy9g/EV/l4
J2cCyVLKs4MaKFRSvR5gBXiosYxh/SGJW+RLpOvxhKRzbifqgAVEcc3meDkze8Be
BEGJY+cHyveNtBzfVu4CQneP1lAi0/HfNqtW+GEMCzZJHEMD7zX3YRbu2HoPZuzp
WbzLcGR/yJ/RZYIGzN6dsmDgr5M7nB1243aiTZx4vHBhNveRjfu9VfNWxvUnz3cG
rrdS75vmYvQegyceKbr+B89LzPSY9fiFzROWutRuvW+/Kz+rsWiAmZAgx29U6RD6
Np5MKvUXqPQZI1IdvWEcYk1tz1wfiRhAOftMcVpMG4/1T3ycVRrXPolSLIA8oofA
UdTqmb8uTm0M2X01Fwa5wG4UskHk7rtXRQg5rMQjKLL878ZCG1ntiRzi4oprWndW
q8ZypOoKhPO/w2fpUSHnSGtk4HeYU0fGjxLWegUxQlfSmPmYV4kXPm+Cv7nD+6OF
VNr7cvVw8UZI316+XQ+1Xj/xbadbdhopMzD2oExzoPx5l9qW7RR9e5y+oazRKnKN
VmDh6uRN6F+4flF7S2znv9DSFIJMjWtd7xUkwsSQn7cIOceVdh3NLPSJtq1yELed
h9yKi+44RFLK4fEXo6tSgGJ6ddj4sX81hBmHoZ8GIlECZpEhuNFzGomfUfgS6Eui
N2yeW9Il/iNbyJGw4RZsTYSl3tzaok6hRm5udD4D4cA0QFwOE4M82l9NHTeXuCIu
TkG04KB26ukoPMwESgDYRu6qYZcVY2z/C9vFsgwJi6WU6i1z9t2z9mz890MCtia4
MydhoIFrmW1wThRRizmq7M2tMN7vUi3CXWCPxqe9cKRxvYyqqzzQ3qL8gEfKiR8t
9jH4ChdpJn5dDkfvd1xhoLsYaUk7PMfSVCCinMv/DDvbZvjVfq5/qvhx48L65dO5
pfqiWpJyJUj409KNUnZxx3MW88EgCzc5NSDz8TRZIES52nRuLC3wwdS2KPFUKG7N
N4jbh/WejNNpcCdnYuB3p/jiP6XAkPiZ6IlwXDxT4snhPMuA9+MMlpXa45c1by02
Prlr+ThbNX2G8G8RQL4l5Wdb9hw0tAsF+U8wmS8JVy3AyHHJ6g7HNKHzL7Qmbt7Y
Mlh86HUwRqESvUtd1QBfLq/XMX3xZuWge4bt7x+V1EoZ9LLxKXLk19RnnyzPfUvj
KEqfGQmuBREING8GWqiBsPaZb2qCMYeIbbN4t4JUYMmkCZN2HN6PBT1iZwF4yAhl
/+cgrkXKonf1NPB9tWE0PHeUOwhKWqW616DGFSOeFIdsaNuw7grKKZa+IbcYa1oO
42tH1rzQOdqeZ9aZo8DfCw4zg0ZoBPaTXMaXohQJDhpLa56wNFVnAyoezxrt1sWF
Yz3sgJCXmqKyvW1JA6mDO89dlHosKITZBqB0WPQwsIos5VKngv1CqZomX3oEqMZs
VOtm6K1rZpsAyZF9XzxwuzCaF7awRr54M6/yiF6JRcALzZnk9ClTdgGqB2cIt0gz
3OQ0YbsAuGVsyyCBXNTWqs2pkUqFez+i5Jz6d7M+0xVG+8kmaRdI/wjSRM0m6CNA
Uz5360aG4mzsuYhVBVtrXpdt8ARtIYqzXLc66QBlN+9L4f0gpSz/U5mtZBut8sEQ
DCX3MbR//u89bOaWh6K8SgeF0//7yilzhlR2uH4E9blPCCa4+MYofppp+wqtUwoo
C0ygbmF5jW5Or3AAkPEUIxQadkh/oXC8o7slILKYdqDM2c9IVQ8TAgjXZe3+jB1C
GNiAOXBGtwbZmtHiVNeOOh7ZC12QBzWR+Z39QRBlpx34PSqZ1v5tcNWotKc3tg67
+yENKXOflda2XcxoXf+bVyRxi46qxDZnldF5+PdXtod9fB9v9hBwX71t9eOJuc9r
HolMHzDMiznpHh2cR73acUZFT+j9lMhTpwhqOXrWjE9kp2uQBhymXa9xW5eX97x+
S/l6VgWvd008I2W3nam3Gd9u2SHVAeU0m43T+i7X69YTh198fXpy8SQ/PK37AXU1
6oQkddb+bmJZEpP4YkGLs2RgcibWyBmuNp4tGBH1venQiMYP+sW2SMS/pbRfQu3D
KEI0uE8/0eajefAKiAZIqSZon7oiQ+f4uAmxKCt4INijTNSNq1kq9B1SyATfR1Sp
XaFj4qjgnDVdVMszZXYqGVesTunU+HPfiOoQLk6CbJ1J+OCfLxA/832LEEEN9LJ0
ZeGuZZ10WarbgOzCPgjmJIbIvoHF/5uw6fQ3Hq1PfImx/voYxgoX0rs2UXLzRY7s
NzgbdNEhXLsd8V8sIwhvo/kYbBRanNIdRHYBSI6qIGOIEf+Bi9tKl0AX5nfuGZZF
Jv7kn0c/KldhArafwFwt1iJxEjrhytdsv80Wz16bwEXCRMDHkHrfJmSbnlECi1Xl
yLm3Kgo/sQOuLTGvYMUPAio+Ra6rmnue80WZRY+Pia+zOU4vSkMe8K11X7FFmTZ4
VqSkjXTje1dVPWGXXZUvzMoUIdY/+CMa+OdmZrs7G0oGFnX2VKIi+bpFD4NZgfg2
JDJ2t720wMRiVr5GrOkaGKF6USqlI7J7KH6fksTNde3k4SDBcI2lhLQJZnth5zhq
SKmuo6bGGIiSFKpt+BGD9yrjAX2jHB4Ai6BpurRqQv21h4wTOWL6XK4cQYkRAGry
+9mVqogZGLyKxaGQW6aeoF8Pd4p6D7q4cvet9z7JFHPjBzrpVcUsoLk9gH9+V5Dx
8GoDk48iCE+6gYfZCG7iGd6Bcj+wsvysmD0ONNMBVuxbq5kPiE3yrtg9moeT2kVp
dpo81kBWw//2T0W2Gq9Bd5IN2ufggQg2qpyolCYHU3I6pa9Cb8qekgAB5l8tKZpe
mFTQmxmoXZ/UWI3ELt2XiDqpXiH6qgzlsVLax5m2NV9THn1+5uERNclIraeM6+Ei
gJjgTrppapOavFb7UCBqs3WVxr2v4ZQ6CC+aRm3R8F1ghRg5TRgLgmBD044kPDnB
w5jJdTNyMxtNIds/N+5pFoX1zhLTEreoeC4/S6y0WcHgL++aKeZzwha4S2+PUBhd
RTcfLjNUYYZ7XCb0xjwXR3djbUvOIGXHnaopwXpP/L+WMSJZY7GWjbz7RtDQ4T/n
c4Q8bLbTdvxjA9WMhBjCMJE9VnXl4/JGmfvHDzeVyiTf5S580Gd+YafYinfP7dW5
NUVJgqULcIrRnvsGjhg7WAgUvb4ZA9D+lPHmDrco7GF1UZqHqoYXv26WxhoOgtTx
pt6SWbeXET3lZjDaGOIzW27Mey1hB8c3HDBxjMSUi3V+o1xosDGKVkbzFzcrnYrM
PCRUBmczj1i1OXccKDAQh5cEDPL7vPHy2uHwsduh7zrgrR+A5Apo69au/RxwgknW
1FtD2vYDAGweZCD/iMDWAGnrfL2QAKI6VsoC9de0wUeT1ps1Fs9AQFCJSGzROF/P
lK6uZunGp523fGkPltyVe3Picv2TmBj+RO8VsD6/LYI4zYC2Iu1vJIf6ib/7ZVQp
H7Gx44/v5UDGJ7hGQtWVLjaoT2X5cO09OBhpVp0KhIcyRHMfmyiJOB5H2XaB+zBg
KZMI7HC1E/fUCS/ypJGY4IXiJ8safxJZnGL6QPqsSE7Kpa4kgTbvoD8OAAgWVk/2
A43bzy9FYFgf6oObRDQNR9RTEE9IaX1lMBj3fXeZar9jbEpG2GvCMUwy+pgw9IaZ
oYN/I5bKISPiRmfuJYtOVg/keGtERNHr6smJ/nfJ+GXb81qCjXgrw3oQlxVxGFfD
OZeADa5mNP5oJQbVcIyejSIzPtfyAEur8dhy4kJ6QfpPFfkMS642giK0VdBOura6
KFryUsmN4aH2tuKLl0BP5qUuKu9OXnjaYIlNxtZxiRR7pzIEfY92bO52TIIgs9MA
AGdQNcDB/NEFPS5DAvteRzaa/cdePpF824GAuKZ5O1JQZRGV/5TKdnNS6bK5qXWE
ag0oEpHKLNcbM5DpfYdquL1HzGhTRMgEDcrr3xULP4YS7GgK+HdYV+tvy+Sdtlsh
eRtlAb7dt22VXfSDz2i0HGBWLDrIldVXkQ2MXGWQRYKJAjbYiNyiaAwdUfHN2XlK
p3cUdywIDeou6mQSDhwyAUI6fJ9XQngDTIN2H74DBInsO2xnTvcSi6CY2dBK4J5+
4F2661nDu+DbxJqXrSvrGX269GZaZesff3Wd9ka22yNuUNHItVGqDu58tzgOPtwj
A+jIFqLXB7sqLGsAHobTsBQKHVRy4ERzBGJ2D3pR0JAZRF8mkiojrrormDeUP8gj
cPJNdlVtTk9cZTlgnJWkJ894o0BUwKI/A0g/0F9hNvmW65AxkwAYSKg42bQOHLFc
vwFq/lHieCVV3O66SLeNRCWS3n14xkY6QH1n3XX53RWuCqdX4XU9/wI7Z1Uynpy4
szrF5KdKLWuZgEwSxns8Bq1c1uS6g2WGiZ8ErnFHErqZMDFzjTpa5QGeDO1f4Hw8
Hm3T202hc6M1vLiNnGfuqw5IKGHGMSltGoECenD0Nlj2rFpkrDymxmh8xMgdKUSt
DthS65wk7hS5tnembJQpzPls2SfVvfrItVdBkJdh3iiK35VjL8aygE7gDm5uvhRX
R7+8Os6kz7Pf1k8MM5QbNy123EFcJ5uUEK3gAJCaLGv6efsDqYbnUfSPOkpAJ5st
nDq4aO/l201aiDLzfGyaJBO4FPjV8K4UCC/LDA6g+B1jGEmlXxUbDAgXyZXpRxbo
ca3RHaMQSzsmo9xOh/XwpDKu4DZOZ87WvAZJFj3uR2luj9WDHZ4ic3vB7y3RI/hO
OSGBU9zgkkpiNCTiL2WsmUJi7WGat2h3h9zN7d6jff/+Z/T+w1nJMQ0CTulLdXgK
pVftO3QS9S3MFFdC/TcpBd98PAYAoFDzfdhUfz4y2nsECnxlU8qAcxnNHwq6Zb7V
MmgHgipHFRWCZMPz2Kenb7q8jjAs0L6yxTp3ARbJTentrPn+eRxL5ydWyKfxKymQ
xJfcw1HwvtnsCJV/mpW2Ak77r9DJdSnn6OaTLf2kvr/SPbkNOBBTEHnZOYMX+loP
Jek6mSzSCdP9Q+VjQbCi08Rtk4zBgoZmV6OhxmZgHEla4wayPwIBpkviKAB4JllU
9y17LS1A1D8sO4GBOhge2oYu2brYhX4V/YuLdd5ElHff0+kYcUtpb7Wci2cOUi7m
GA8b8QmbrBY+CaBxOoPYjptEkYPtpHO7t2VqjcpD+d3xWse/mJJUhtg9kapRkbUz
xwSOyu49LiotAeRBQvUYDN5UivRMo+5Zna2BPlECcrSA5Q0FkEvWM31rBC1IoPiF
7Vd76r7zZ1EvmBTf2CygLzf6fT0N2L80motQxWfstvkKJYN+J8wHadf5p1Oh9TWV
HR4A9d1XGGy4k3N8QkH8Qp9e8exzxf7/exd2H1mV2w/hszf/Fxn1WcWQHdLvA7u9
uLK53Ir7YKMO1YHTvKk+lxdbNhiivaGd90l4g3Wn4nvnUeHbvLlocnUm1VYHb7Py
UrW1+E6V2TReSrmaqlZ4+jkl0AQml6NTH4GFfZxcPUZqvW1R/cODHA3w6g3X1Q19
DJZnE/qINGzo1P+T+bpVNpi+bNWcDH3BgW7+uCYLJb8P97lXkD9Eo1+1gphLR8cu
+p8bYPqlOoCsk/KAQeVRk9FI9fSv2RBQ+ZmAN/q5nv+P8y1ajKNij3mDSlDn6HQ4
FFt4u7tUqPbT4QaELmlEXAAjagpSrstLWTHE4K840Z9RyLDNFn8mSkAiva0u1eXI
lEDu9kSE+tKPEofiNUAtsLywI1yqT9SC4aO4mJDV7O5DszIlv0HDtmFwDuKuGe+I
pm7ZDlEho/ZisztTHLgW7MbFssv3CsQHJDS5QnNPDPWzjGG4IWwxZw8oBQzxufNT
DiVbI75nyoD2ngzD2Jc0bO/oB9rR0+Ws0ZvHcXxAAOOakAJK7gpoHz4UAOBaiIYH
gmGLBpiBbj1M+KQzqIvC+pTWgtuMHRm+BI07bxTFUFB2dk1x2kYI8k/cFCYF0cwj
DD4cC4n00uyBGBznJK+AMfMnoN6oV44ydxVhW+uCP18wievZPD3SIy9JQ8R3Ob+8
JW+Ur4KQLsM15SbbcizEm9TTTndNBoTBOOR6E69Ad3HWDzPnu5ZMtZgBPm0M30eL
qfhh+dRGEV67ekz00Mu2P5Rnpt4xRf6IQyTsPZYCgRa+SO1DRhFbsCvedo3rlyBJ
NpPrYLiao8EjXEc1lbe0kMXuFVE/Tv5Nvph7kymOc9ile/tWGILWJloqZdnvS12g
DyDcTlPwSbKcdHRrHNL/IVhzcr9GJNbWN8pc2ponCTj7c/E9XJJEPe5A0V1DoQfE
YMtsYZ772eCZhnVFrdvec7oVrAZiTtypzoZncl5OsPLBG05xVun7cwcYIczigehj
bXjS2OdpVv5QiC3mOEk17ts+rPcCXta6oIZgvsmT9zPWPHoTuiYLNX/TAyoUhjTG
lhiy11H0Ck4BpJemR8UH9FiBYzXIi5F/jS6C0AJTfJ5BiBEFavyPu1IzBNze0dTp
aUw+pLOhGK6rhJ5I0lV8vk/mj0tExneZtM52yzTHOzhoY/hofPcftLTfpFesc4aM
O2xvgtr4J98Gkg8b+P+Y8HsZQ77YmuKa9xi9QJj0+XnY8w333TgdQilwbQFOfSH/
91woTuA+QzjVQh6ZHew0Lj4JdBELjYZ8e/7moZGGf2wys6eLTXEkba7QHofnFeah
cmfvg6H3E6qRTMotyUtZ6pvotnB9SRv1mv75lecICU9b32qKnPXw1L0LMPLmQKKA
VTlwCpOgoqxNj40tKOxzPrkNabgPkbvkOw/YLybOM/3QKvYRVkKLD9fc6L4m6h2v
2DRWcTxJ26+tRvEDBTFFi2djhmr9JehXySQTUtsky5TP9FGPC/4JN4F2JbXVdoUW
Xndi3wVB/j23g86lZu8Cvf312faYrk81r8PGmWrHIVvjhQ6Q706247vdBa2+2G9d
9x8iegzAWlY/cQMTP4fpqykGGcUuP+Us3RiVbte4JjygxOnxF3sLKW8MMnerop7Q
WwtWOMrbnbZE1rNiltvLf52uA/xQsnNPM0ime3AasnCoDR2iNJMYvvx0wGjt6THX
VmRUhdwN+ehxW04CyCkawHg31pBjqu8ftTNB8/fXMC5dCAl1pz8Uysg6dG0YBja/
DsrkqV6nKq2BTCZZUSx1PiuhlTrINT5+6CCfZ0dVuFF4Yt+0/WYNQ8wdVP8G4+jA
93E22KZk3Yx8iF8lqtvlxN9YwVfmC0IHxJUWR8UrWhdLVgkmYENJnhZCMNSBPtv9
B0mvzQFhOoDx80ZJ4NESbYMoxpk8gL6Mrwq8FwA2yC5ark0tQQhRdD1+QX3ir8ZN
fc3PMxL3d/19Cm+P7VdkU28jq5yOxVAa5ZxDv78oQYDpVE5bQkeix6WIwQlT+/WF
e75EyXI+LPTCTgQS2ykqUB4caY1ubkjrkSJtJBAB9J2V87LH3mVJsorls35/CEJD
JuhWcgYCJ3Ala8mkwPUW4wlafVBG0accMlkw7P2k08vYx6gCv9GzKuciAak+wGdz
Vgc7t/cEgjcfQ+iqZ6MRUoK9EbqkpJgnmDIAWAihjexvm9TnZYi4JNTrq5F6jKFC
C/SZbVN1Ug9ZE1xbdIFiJ7ut9cqux346yeZp318T6B8C5dsYA6sYuRRdjdFY/bS0
qq2mobKVgNJi9059j7e60uCWybhGF6/XIQ1zfl4ceW/fZXMEU5cl3VWXXks2ML5u
M2CpcxlMxaGrQHufJlIGTnfD92Di77J6vR2HZFeuq3rMR50ME6HMj4CK5Gn09ChA
IUzePZMUedqkzglbgGP+gtxXpmbS+G48elXat+ligKQQ8UVT8BxHojKhTwv6CXXZ
eyllioH5/skxr7vJDpf4DgGSLAbFoEBj2LkogUtL+TAjRuAH1CbMK9EDQ/GGznRw
23CsfczDRSmJFHa9O5EKXTxedbiCfC2GZJYQKi3coiv7l4znV402XTI4YYUujQhO
MQwhjQF9qino6TcyR5DZzolUwrnsLEw3w2K7dXIRCIXCOo9sBidVl+Lsc8wEcjo9
+YBmUvppjAIR+CzJzRKSg7+GyJZtiUse6PqKlaQcL2UYRUaoYCzD/boL897kY9to
sqnIHq9Q/muXe/EabUgVhrra5cYMatYE4KTRrtKXtXcqMoumoW9QbRMn2DbqaHaU
DDU7kVI7RfKePDkiTHeXVby9ja324VjNTWkfGfbMRnPwbfOftzHzhiaow/UaKtbZ
CbniL3mpSdg9GUjG2gOPnybuqs7FEt4GdIUbFdOanKbjicOajcqlPWom9im5xubm
dtDQQRXc4f1fgl/SzlmfVFVPdoOOT9SArfC75012UBmERX1/hTEBmmv9ASC/YR/k
LpuzOfxUL2N2DWCGfeXR3hi9dPcRHf7AIV644uo+n1Gzw9iulB0PvhwHp2sa1u2i
fNwIieFGhwTWzXcA957hUDddeJmHsYE3/cuMfSpsGQJtcQQMA20r4XjBVDQk9ozu
djFQMn0II24TViFTPiCBT5VcrZoc1ym9t0wD2QDpBLm328shLy1AV02FVJ+XUVcb
w6745VADYvy4VjKoP2LgBFjaz13ufUpZBK+dyVKWfiw82tWuUbXtepP5qW5VdIlP
1xAXdms2GQjZ5ME3HVtxA0Onw3Hupx9b9dib50Gjdx0f0vErH7l8FLrL62tKizYm
sRIWRo4h+hvuAComc7y2CVbChjUUSQQhpWKXDFcywN9KFYRZF6cUKMpTAfILN/6M
8NlauX9mDRMXf3ZoAzRi4WqmQJRUuQ14ei4nDnSaSeVrxKIbmIp/obkvaQqkz1j0
/B5Ep+dQovhcsEEHyLsFnjcnVzVekxBwnT1tdpvhVOtXSCQ+TrBXoy2drndvnuxo
4z9cOn5IoY9vyASbSl3+ZxrQ9401PSeVkWRMf/6FOgoZ9Q0MqH9zi9QLoxCsEt4w
IVkrj9vFLwnJ/wUj1FKyTFqIw/VBrI9iZABh+hcU5B5VzVef5zkWg47NS8U5qjT1
DwAZhvrTyIrTF2GoXIC9ZE80kHxSGppChIg2p+K6nCzwaD2oW/hdiKkrXIT8674b
lyz6E2pbqVhbe9+oIVHjfKiW2xurM+Ja1eXNlwpRTv0og7AcgekhbdQ7ZAr+BIUQ
P3+jADRwc7J9oU10KI09+K/9ea2NyrjC2VpTvKQBXAeeT2ev1ALi7BicW6B9KRPd
MkxSpm8+vaT/WWm9bVqbyf6xejNKi7Uu0Ca1f0bSxGQ3Xzp/uRrGFVgUuaDpc/mr
jqOJsW+djqLdFAxfMC4a1oY3sVlZL9TwDnFccMvOgfm6b+TEMtirNNvt2igXeuSj
/SGg3MOu6QZ+UeLTC1H0nUWg5lYHRsmx2pWt2vF8llKNwx/rdEnq4Xvhb7sDmDmW
HF873PdDp0VrVDFGY/IedN6gZ88D81eYMQomxOvgo1n3au11BTyZH/tA8DEwjdtT
Mgq5srlvjtrP7V9oBTyGubn9UMt4sVhTMWbLbhFZoKbhRccvk6UMvkTvIxTqBKh7
X/y1f+13Q0hLqA+C2RZEYY1fQ5axnauUYOaWsPEs5tMQO17JSrrPPUEYBHBzkrsh
JKyJfgWcgQaS131vdBboXoQUJXGN/Tw+HbKc8nbMByHbYf22e5xE0r6pi6aj3GDM
4C+Yx59riL+PfieKEJE+m0VMwY3M256u6hytsS3tmGE8EuAN+ddFxk0yabnh1z+c
gwJZRp71Bw/3OCVvmH65ieYJFB4og64tuOB58O04nLPenyyMho4K3M/hlMUshAts
JBeqT8DEU5RNuAP5Rzmy3hu9QuOpbd8GhwpTLc50TT5FbNbDPRYvUNd2GOmLXFBf
2rQP9J4/NwGqG7lllyXrNo615zQPUxnfT45jFjdJW3hfRglN1HtFNLFd8sGf/E/3
YR7C2nIGLZTGg4QAlMKYXqlIenemvAIGH/i+a3ld+SZoG2z4w0CTdVW/rytVq8M3
82TLkbi1ULBtW26TTZcnBXB55RjVbIoOrMyv3ntQbtl4QUYWg8HpXNgwdgkz5JR9
22lUX1vr9twnIuqxa22U7xunj3TAaIC8nxOrecUuUBu/eKmr3RFYFQoFk+kQR8vp
nusmZ/R+M9/d9jVApIiYNSUniCCmz5ybx19nFs1MQthxoXX4FpVBSpsRpa7TKSFY
A4gfWlwPzObPq1JS0/bCOrgkGhnPpcnd8MlunB7B1T2AsAC5s3v89jBm7YfcxqOd
mx8ZH/rnRp2qoDGZgttNvxiosSOiX1SPXEcLIwlSNgPhWCrua7g32IphxEZMQa0N
P0lP4RUIFquFeRD5C2n/v+DDc32Q36XBe2omPMdmjDk/kPoqy8BU09p7v0rVDsYv
lfqf2ewKBV5kp7kewaoUvsvCF8vSyspPPaBPt/UO0VKjEyO2z1OJNMPbIOoSG9XN
sMr/M6q21wKCp46mxs33PC3GyiRsoIlCzXARb61PznPAVbjLgJB3qsKzHzfD22Gi
vyut/dx+V3rdo/JfbdvpFlxT/zbdRudk6sEgiW1VqT0S2AMvTphsZHot15pWUH/Q
PJ0ISne9ZJdUJDFVyDkev6rviVs+yH/mAt5zUm+cU7NagFoTcDc3uf9n1vqmAp0l
rOVga8xdwjhVx+o4fCZxbv0LEvIV1rSfNZpqyGgjvfaWT4Xbv60QZ3JEWhpEst0v
/nBdjoUvmA1jxsEtt+tHzPGOG7fqQwPJCc5nMaEO0Jc7aQpJmk3ZEuABZJt6LWuF
lecQvMDp3E2/T3/rNXwSXE8tliDme6zYBOQ+tVOOM9t0mojFUTBDq5FG/E1NQXrA
JSBM2dQwaLtI4PqMsG98tS9UFRvF9+hxkuJikENs3ITNwKTeoh37yc+ygCaWG0QM
AM36RC9DCZ/ZDJuP+nA6Bwt5G1Y0r82W5BLoe3dBUcJZd61yk7tO7t4V1fyjTh0O
0VDaQdBtp+yoC5b5ROOrcSzPtDJIGecAIKD3pVywIJrlCOTNei7RGQ/GCTuo2cRz
qjlxeewMUQP/j3qN8HYkym9SqpWYyAggzVfrUb5hIzzIl8uKpXw79q7oAso1/hdZ
8bJ19ROf7qgVL7dzeJU7yVaIlanQxmvr79OAG3aI3cL+Z7Tb2cuJtfNHJNrBn2eQ
m3E8juWRWeNANyBL34vhS6gVC3oMWXI5qd4y4r2kr36M6Nelv1iBFl5z4I+xhnK7
vFtes2oLvLAPcc7AakiLdXFv6nX5e2dYRnq7Z3tl/VaxPxCIdScagLVN3ZwV5UDk
phWxKQokxrdOTto7mCy6oN6lYpH0w8Ems2V6mWWQ+4Lrqk0kyhapyqYLNwiLjTFt
X0n+gbZr47o4KNrwi+MhYvZDjLIefnJvIUEZU25qRFqTPPw1IbtKQLlihCep9SCy
p9jhxXdaqqu1RaHar2qd+aFZcezoOrOUI0KoD1oTStspxyTNljfBpynCpp2DaTjs
EjRWw8b25I4ErJf339tyMvg3h9Ru4FAXXTRRlWB9bzLU1kgiYRCqzaOp0xB6K6Ai
dRN9eEEhmCEBkahFlqwY90Yj6yQuUChhPY/HM3RROYr0zdCrwsqmtuzQWyOS/Q+v
CWpDQp/3OJEdjJCTytbKId0G5sbf+zcfqcdrEze+CmMAsqacPFl6BDhuu2nCypPc
gRBXdK7YOcnXGFPWGbVirFWamDYEeeJs7lth3Z36744TQY1bu2iOmTeEOh5eEFbZ
hbxtqActdtpMK8wxygiyVhchgRzSnMoaVmG5z8Yvt7/zd63Tlt9rN0suzXgm4bnE
+tSSxZkSpyy+c6KP5ZFS3sdvY6YqByouuKaZHPrTo+kJtBLfMi3o0MSibBPDynlg
cy0UemMlX4muzdd2ue6R4EDq3xielZoA8nzbCmHf4Qb+BQZj1hzgeAjMyLXhDuPQ
c6vCRdL4ywT4FmjBLkw31eSvFDytdOvvksnHBtB2uqEkxzeUaoHH/LWkcUHpsIZX
4SRuk2/U1TBItD/t20jmOqh08ssMmn8xQwB1sePJ6WsPzTXlD4bmQHYMoTMvXGoV
TOz+M5urSYujgW3dXupAARGSo5yKeJ9Ti5IewyyxmYhYP1We51SDbZTG6DGG8Lf/
k9W/gnKH9Sd69WNJngdw7THVz84nB5i/fTnTQO8Kzm+wti0tV9LG0RW//qgzbvu8
xstowS1sLHA3laOrnT8ZtvZ50y4kXAIFj7BHLUnTn7cmt4x+4nd2qGL32xX0phhj
yvHuJ8qonA59PaSNp63OEHIL/4h3v9dDt4+p5EW2NLlMEwSHAWItyVxouaiAwYvZ
hYvD+EAWw4cbmZ2Op9Mv/x6UM4M+fOo8Rlzz8FZ00D3ijD1VBHrJOzUebhB/wvNq
hLTb5/zEfIflUU1xlOzFE0rQXU07Y6vY0hjTm/VjpeG45nzvwSBTxr79ELwqEO43
lSbpIAMX3dhIjvp9lgZteOe1rlY6XroNWzmGke6KdOKCIM6FyW+Qu+D0oZl6hVzF
spMnD/WAd0T0vgF3vFm2o+IPDUfsWpNGuc5Kp2VWXkI3XSwljj3XMMUZjASuW9kH
7f7OiYGzkiuIpMfCf6RYMVb+RVMeHIFcuL1z9qR47jKKQLEwhzsvJE1HJxZe38uw
EusTZg8C6icO9oQ5yRTMdxpG2i67seB5pu2Jxs9DRWFsINROREf1zqp3N9fCBLWf
JFcVejwg3GWyPxKH5l7ls/xPPSkf5IQf4RRGE7YLob189F4gn/ehZJzrczFRa9mH
7M5UtvgVeA9KNFMFztdCMUhd7lpciScNuFc2mYiRqefK84nvDL4pkVrc+5f9k/wj
tnev92uQUx9jtsK+KH/YNPNXp+L2ZUQmYbk2eSxeWbb2ZtUV3x+hUKh2KzH/WxPW
wOxB8dNjZwdIeueRt/rP7pKiaXO3r+pOGDDKa9383GoUSB25j7xrMxdZpss1kc0j
QdUTmhBmu5TTxkh2n5VvnpoLOxlPS3XhWG9c6jVr6KMwLvPcNLm4CCaiePs/1MHb
sX35VMRcMbl/puOFCIjMyusRKY+C9gFhnBTLX4VfRmKPBIN/V4CHmuziIF54Echf
XXK685d4FeJKyMWvwlsdnzYU3U9P7erg1l/P2Ixuf/OHtCqD3q4DCd1wjLHTZhki
gRhp2slbhJjgEIMvyn6Mty2D1wzrfmjY9t0y7G+GB40/HnZoLskFzPcSIxQ2L8pv
jD5RX4is5Z7Owu6CsBQ7iWAJIwmBNLLVPyJTdkoFZ73gZI26HzOqFWPJLBQoTkXk
IhBGUSdD9IGqBOJejUFoOpmJuCFIPgiNl2WAUk8W/HMbAOuaCJR1/gYbPQ2uYT6C
fpqF5EMbMh372tPGvQMIh6zEIrbvVkKO6Jks6HPuq3GRBlkSf5tebQNqIo6nl6qm
WgJnxn3BZXs4m8FN/89MtTgyadEk+qIkIe61GGgt9dbA374x8tkPb7MPSiNHogFI
o+e1IT5VPkPajvrTLbMWXe3Jg3fVvksO1Xc7sgWj3oRcMq/Fa4tlvi0k8LN1lsz+
zgdn02K4ikPUgo9p9tN2l0QP8tC10orVsKr3YkJhAxmpZ9l4VK+mdQVFMtRz09Fh
7NAG3gxh3pJcpvN4pRqYY6sWik52wVRkf5Un40/aQSNXNHaKjJMVANoZDg7jihU5
UcMq3guU2/vIVw42iFyUskdZjf+646GsUYD9BufwlvfjRDrNx9DLxphHnW60uWiA
GgV4+WTOcJ1DIonmRFIUy4s2sDSCFefIrMDH4t0iw4hg9o1Aahic7xqjecfJbS+8
Rbk07D3YPJswjSghDtkED48vh4PwZc3xlTBm3O5KfA2MNofVMvH13BnQ2UFZD2JS
XB1/sLMmNB7DU6WoKIgYK7hZvKFzcHjkEjgv3yRqhnczWjZG3xfIV99D2zB2H/0W
HiyTdnvPd7dRYq1V19DuEWvduwlleo3VC4yIMBsZ0i95sGAQLGLyN17pzOcnjXbo
L/tiyJOjzkmfxnCjTJrr+QUmqmTiaMt9Y0199wWfkY+zJtxnHRNqSpY+wLgPYPpu
A/4WaEk1QeFXZsMCjO4SGBVSE4APNH9SNY6vdYrqT+1vwMb+dXXYs/eQJ/tNyTLY
Nav7Rtup6rZDbrkS1djP7KZOW6wY7VmHPVsOJXOLCfrE8eNxvv+i+ZdvjAXtbdKn
W2xHs/0ivkFG6UOx4qAr09SNiZC+erFIy2hu+Rvcaq26FjOUdIclh2+I9CnheIHy
yT0sKRP5icFPoJIAOKsL/9l6LMm/8qyG7AuWjOiCpoTEOQJu7NcqOLgq7sfRL5FF
FBXGOokzXuHDKiqXrWpeS1M3Lry8XZqqisR0qfppzQ+ESOtFSpL62NwEj8EhW7qz
pXpN63nkf4VxJGDBPlDsUtRLv50awXOPnYxWYPVzQqqgsi9SOfoKnYb8QGEhnqe1
CaX+EQilh5fyiCV7wGvOxGhR8zt1uL/CkArEXJ+FTFtIXB67MfML0vp/m6wtkRFX
emCL5pQgmk4ZtS5fhH63LavjBnCcCEGy1Qpl9uwAiuGDChM49NHT6nn+ypxJweYL
sZaMEXtJZ0C9x/ASaQFjdyBkb3fnAS1uC5QGf4u0TGm649ttVfZfndjjN/5hOp+n
iUb2URDnhYdWy6yT0wo72EUsfi/9xYQyycXa7HYppMjg2aGorP2iqLUuAo5g4Ej7
bEJR3dA0lQAcxTirbGHkh98dI6Z1INKNzyQamR5Fk1ZUtGUNHmZuSgcLitItXpok
uyLMjeqmxyZI/DfKtbZbK6Zx9ZB9pKfdQjtGmaFnygkP7LFNRGDmyy1zgnLjhKoe
wQJTQ8IeMBV4DeQ4giqtX64uBOOdaaNd//8w2fnQNadK8Fi8vnc2vAcrRECn/Ah9
/jnFPy74oHJxNw0DaT9XExvvi3YJENm7WEIaHOwmE8jA63dQmI37YtmtXtp82rv/
Acxyf8SUIOOoC5VX7Q8jclTWX3j/POYDrCClifr2QjRPH7HcuIIacl8YyhCLJQS+
BLd6Yl9xftEfaeJ2BoiiSzmIRAvvRR+SkTrjkjLFbKljUAQQnqpqWcWLCPnP+R8q
nlIePwBeA/n2PCaXg652K6F7ScvSDxr46vtWsY2WwkoyjuVAwL51wN8gYD/9epKW
Nt0pKlsP21rqMIgy2/gzz1BkpczecQOz2bEblIQJBfy7aKliYlDR0GFNRH+AbwzX
ourTMXWQx9CFR2JMcLDrEiQdT26IPinekaqghEM4FDbMRGLmBMPulgiAR7+VR8lk
leM2XppAB78nL1tw6h68VSQxp/JT0jmf/AhYZ8v3AzUyQR+BjzhMKqw5p08NaTUF
Gmt839bbs5jB/4wXjLBT+4R7+6eIV6l+mjLtCTxTeZoH8/kHQPrg7rJ4NBttdiIq
0PRO/S0gmtfxDBB0Ta6gvA9PRXkkBwvdN10Aaa+tYpGthBFZzHTI9R41pS4bqFyV
j+FXM+hCAxHWMPRFhMa3KeGoECsUhmDGoxBEc7elYK+MkP1P0Lj6pQgt85CDZm87
Ft2HnXyQSsDiMGGQ3dexHLcw4JDYdk1Nx2AOu53MicZY+FuNba4UuS9Es1QMahBJ
76x5IG1iqMw9RAmf1rCmaJyjSXNdt6Zqnyt864eCRvu/6pvBB2lO8fW75H8xCV5B
3dU/J5s9gVSE9lW5jE+ASV6iNTjoW+6V5Lya0Uj0hdAJxYo502XGHu2oIxyNgk+/
u4k9+af5F3ayZsF60NyXub5Kdln8w/Z2pn7Okww18qAN+JcClVLNN3tG9iTk3uyJ
IsuHvVkWDm6lYMK6aLTi9Z+bT23vCFKZkAtAscI3oeU6hhrgt4BiROicO0LhOLiO
gsWx5UpYCUnxP42zOQP57I+xD9YFqpmazw/vrZmiVIgHUtslKcZErymWZJh4bQrD
kivOoJ+tvDSDOUSjH5VyHX0mKWJKGr/XMK/pWfgfIhRYGTXX2hUsCjamGI+geIP1
SzrOi/lmSleZZF5U5JAOEq7e8yTudYOWv5mdk9u2RKWHFYeyvTGxjEpXWzUw6vHv
Z4RMOK2/BYWWv6kJgZrB7fGXcrBoMFlA+2jMK3MyImmUMyqDuDCPw45NWOg4H/SM
5PwekBqYTSVhqdp2l1n87lNuMZWnmX6W8jCDwvVxvcWsOTzJzJ8405rXkYXUeBv/
oqVgO218pAL4SM+hoYTqbDy240fIT6pJbsl8ows5CpYtKJxuRkY88ccV1wV1bvoW
QpE/uOV7QbtqQtGpSCuzzY1lq/NK/gQ7aA4A3Wv0EWUPsGc3cImm6Xi6z+ZDGcNF
s3P3NgA21Eekho8YbjNsAADQjROFFS/S5q+4KiuPQbeGsnfGqKogWWL7uE+oXWV5
c4XsPQZHTHpVfxjmQPBlTBmnP6UPaRQDvRLsdtSwa4x1K0zLloX/BkqmhmeJMVYQ
I1lODzargEQpViLnxpZAWJ4/T6qPfdRTERuOp0XOUJyRbLlEetM2VDgRZrdNJVFz
vSE3bSAe7aiXFpv5GRpjr3vpevmH6782DgwMuutbg5gIvNdQr7AvhkfUUtu9e/mD
Fmdw2tZoMR5GgFh3vHrMtQpZntp36lvf4Bch8rUz86P1FUkkAdGa2GmnJmS5VrBd
WLKAPWJopKFfOGbknUlma0lX7X7j0CilD2dfGfSJ5xu+//XoAn9jNS6E6f7yNM99
1oyH1cCAon40hQ3uQapL2veDWNIzY8A+2+6rHim/M9bCXlbiEEreXxcgdNd0tW2A
/RsxLkM1RZv9oxrqlxPGT2G//9kPgvy4ANG+jyruRt0/vDCSQ2SSY3GzeyV9Kj4E
1fgor4mfXGJbgodhbggI9ebe8kB6S7HosN0xYhtO9www76HiSRDjmEk0vWBOATvm
YZ4Fs85l+rjpFAg/onMyk6xawX4DeBz7MWHpPPsQxczARIdSaNtDYVg67VnEy4Rq
l8nIqxcLdIhCy5Mdpym2we0QbEUTHAtynxBqVdHEBHAz1zVyzmUzfJXVOWmx2xLF
Wp7lBZvqEo8HCIs8Bf7nI3NGBh8TUGDuxwF3g2Nu1YJUEgHP5MwP+VAqLzgO9YbD
xeNH0+N9z/L0GZbPDAZ3jq6A7Alis/xFj1IKqOSY7AGHojMQN1ktspVtedavJ4+K
5hxWzfOGR84rewK2YZJgPAJy+B1ho2Cc+WIIELeKTKXofpSrQ9SNrpAV79U7V9HS
SRkDY3JRBBuFW/74O5JTxgHQ6T1yOIzumrdDGChCfazZVAMA4lynSbB83mjeH8l8
jHwFvxuf++cS5e3NDGOtqYmcFoIxsbzIjFAC28ATCWU6G8jC9qpCztTgNLQ7WbY7
E0zIcl53jQNgQlmn5Xa72kFv6c47Cv00Y/3qzZNkhdChdzg3BnQeUKoys5hSX127
DsaezXbbkvQSyx6uBvaEBoQrikAZ5CJcU9H9U1bvH6tC6niKzSIzQHJrlLNpzbQ1
szJ9+7sqSYA6Sgv/p8HydqPfBskeBZ/za8twPt2FOF108zx3YXG2RUnaGfkJ+N1p
XrUBLzVjsXS7e8CdYLPrc+a9ezfBBpSEeIKDD3sVjI2x8oA3w+CnlwQVAngD3Pvt
aGLNewuEaLdRD2C6y007LFqyreOx94lyY56vQ1DX6jAiBItXIUJzkeWb614C5z4F
w4ut0P1Cuyy/oi0GTCOGYp14ukYwbz1bkntAU39iS6Pq+gsPSHBqdohgRZrDC43V
RZ6Re0D5AxatzWd6619fF7k8gQEjnej6xJkEHRo08Mw2YS+lQlDQb5mJtgeqw9cs
Q6tXkVnZyi3kZ80DJL+dSyOd/UmU4P71/N1/G7UKqXsp/PQonxyA8LU1UQXrKF1b
cXke6BpHA7Ip7rzPu6Xq2RCr99b1qDZKqVyj9uGOUDSk02R7KRPglzvBsGRfvySu
NX7IuRMPgvDuJqng3mVFH0jSiiBYZ77FlfW1uKIZheNDFJZ4FW2dikwrrekk6EzA
/DCbKUjE769cOj0lLwRoWX/Nihc08HAtG5x0vHTAl1Lz1GyoFQZkXEx/172vXKnA
PTaKum5OiWno8+KTXYR99j1BtCQvZQZU9dQUDJ8pUB/Fo+kglH4uaeZtWCZ2GXcZ
GlV1rgtUkkPjE0MhhwSVgGTS7VD9hJoP9PVA+yZBbqctnZDjH02Q9piUMQSvByqz
enu1CyoB1KKl8SpCIlVm/cuAPG2xcAfj4MYDG4fHiAL16+u+vKUirM4QaNGaUUb+
ISG2CRY3AarVEvAheRvOi5bM2Me1iQx6iR8Wz6IWhaOZnTwEDcW/kPGlSkGXTuNu
5TLZeEVxSMO83qhJ+kMkk1DFqGp3imL0znkg6+QpH0rywIof8z7aIObmS1M4Zg/s
zbaa3Ek2+ov+R8NkK11qZou6/DUjgTSqTX0v6+iVtkQ4gcj9QiL84w4kFwvDpHAy
i3HrEnS1xznx0sqbDjYh2NrXExdz5o96c+UFzKgcIyka5qgUXNkorU4N8jD1UnKa
gMkLsacd2GopCslwUsg6W4dhmw3GiQpMt0sxfd2WNw/T1tV0maaFbGpzjFciR+9A
3yCfh5kaIVGUGo/g5DPm8cSLvA4U7ivl0xGOEpfls6oPg6pHX383d6LBtKYcGAPk
GbZZ5pcsHHTjxuksTAq1jbB8Z4KCksesDKWqcDqJ/2a4yzUBHFVHbxd6h7DqZ/M5
pWfRxf61XZjF4w9Dt4IHNg0NynaPJ60t7Y0p7E+bQp5+HsX09cb3d2k1Tq3u6Huc
brt+kWay3+CqWqajMVb6xVQAXoifHzl+E+boXSTBVTrDFE43NltgpaJL+7NjtvB/
FTW/xeRpFcixMRwOkG7PK71ZjfGFPrbi5fRCT0vi9hKnwwhGIcgy4A6VtHw8YjSq
2M/3vL8cDvb0Y+Iu3IeVZ9P5mYAnbn5yhqV+U0RBjS6vwQysyZ7jM9WcE8rKrbJy
2olZqlRABSnWyru1TF9GUPpiBqndn07Ift05ju1NmyRpj5AO2IYbsEZHfgIKJHRm
PAc2I2tvArPSqIZi6ZPVeNrQMBNLCq3T14+9F3njxSir9QbqkMTlSaPTsVArkvOF
Vzxz0agrpfw5o9U7N2/GNL6j282YbbWnFg69QMCf5gntMhYphekdiTi+XKtOCOgZ
yB5J6zgmHS3xZbqVNni8SNCaOe+M7dnRgEOM77a4FwbKQf4AAjI9nGHhFxZ/osI7
mL0tciR7Y/A0Ck1iIqvnr8juRB91lBz1KrApVGpGSU0tT/sZRRnmJaLtYVzaw6l4
9TzUWr3Ec/j9Zs445Yvb2PPYv0JOc0frLR7WNXLZ/7OI258lAaoNCCwm80YI1dl3
9wH2LKdqyqJpgcH10pUYGylxCKKbvwLRHSbD5HAT0HOX/BbkjqC/Ottq1GxNkDnU
gdnAbi9glh9gF9bBBGdvrhBObQ8sNgfe0IeZDfiIpOooU2mKOps4J4+xKKbmHbXS
aXXR772O/E9Qi1f8S8JPe4Bnvb3MXL4kwgahTvxj8POfjSBWQ9+GJYDjPWTi8BKB
n/4Kpx9J21xpgOwISeoKw4jg6J+nEMTbqG6s9spk6CU8pwf/3+6I9Znuz6f6TiCz
ahg0/KHAZS8dvN8Z/zf7dKzlA6JJIyJgEQzHLgcBpmIFuf5U0jl7qubxc1DeTrMU
L7cmBoL+6Nx4rRQ74FQKXBPoA3Ttyf1hlUt83DGpfMhb4dWvgAsuPSLgFVbBKpxF
s1uv9KhjYVw3BxDL/6W7NHK10fVm/RUkWV8z1kA9x3HRpq9cTKHiFqJ8tYK2oHqB
PcrB1RTr059Iq4iO5Kaw5xtDqT2S0o5zf5zkU50xZ+SKHM03HtQLwIf80bcB2QxC
rUDRmd8jgSmJn2T7hI+54PtTtEMk0VmD9BlUfTO++7RHo24K6Q/VXpV8p+evlzOX
I280H8Ut0sD22uD4Uy3goSlMWhzFmuHh18UH19JCx2a8/xQoBeRXpB3Xf3bNez9v
6wXVtG3yQCWzy33D1TVDEMtiwWb78cb7nGOc70uOdZq/2oDhlYobED612yime/Zz
axozSDF6qoV21EGxE9FlIn7HHNfC12CIG5KUznqVTTAPeh/UJBbUT9zf/9rKijzi
pH4hhF3nHAAeQIWew/65kQXyfLYw0096IM397CwP5wpaOXmVhFt5H6OzDv/jSYT1
5Py8I5PJIAPLDb3X1QVS2yTjk3au+8m09xg0ZyM3pEZJpqBumpy/064b4mfiO/cF
w+PfURz1YZW4Q3tLSX7K0WCaVDfTSB3WTXrwVAAgf2LqSchYXFFSej659ksXvbnH
vPzKdk/66OYqNMRtrY0pi2cAezx8Tm9BlF5Va/7ZZ68UEJSpsZtB/1LdlKYfV4ZS
MTNql1rQqBomN+ACG+4aVckdGguBRvPYS+9QdFUlQQ1BH5+P9rbwMKnC61DlVtaO
SyAK0rLAJO9DYddlM4HhnmwkVxfu3ic9ellFUtoGHMYdFoX//qRAyYLrbczqISzv
pQnQlq/YqAm0595r2X7Ak3pA1pQf7vC9igegZ8uolmQDeIVys2mCb6B8XuZzOHhT
wPQfvbkiPVOr8rnyvbYd7KjiJZzBr0LhcJoR+CcpqxeAxo4A45oSXGBvtI1dx04f
pVtJGu7FPT6JZDWW9HC00gIsgXKx0Qi705XOeuQ3zUFxbzx3jnG+phIWySXQDIqZ
rfYSKwVTHm/hOqQkOhNZEOPK6ndhPk9m8II6Kk75FNdkLzzNNj7KdWz575w7lpQ1
2UGM53otJ060AfQc8aHhAgME0xWFxIalgb8qVRF5BNcGQ44QpsfL+juxgHJBwoqV
S0QFKEnBJsWTNS+nRMCaql9qTslx4rkuB6ZOOU5IkA+EaN1QXyrSqsavGttlrdZ/
dCGfM1PwvUBKcc35o/AOJut8WPY9Zt+Qebd8gXfzL02UB6ZxTUOrRUL2yxc6BnFT
E1YS40MtMOH92P3PUsbfoD7bMLtewn13vgcW2LqOAoxw3gPo6PNzlSI6GJ2bbny/
ieTH8zTioCkDFbDDBReq0T+S2Hw65cwShN8OLf7s0zXy594D3bCSESHhkV0xJ2+S
9h1yGhUoAkD7UTFjnfZYGlMPZqTphArcVpA2+1hIbx77Q9Jj6rTOiAVv1murmJID
i8EUIhzY2nloMAwuPplMW6WqpfULdewgG9PqMAmy+bdGdBeJ0b8W1TrDNESoPqnX
7urWtU7QF68TeN5QhmFKYn177RdsHfxKz9NQjiHaSfaGQoGr3XmEIZPBpquu4Lon
Qzg5/lYQwyEmkfaFFbb63chVRRUJ4hLzJsjJFKe53tAzuVL2h530spIPQkyga+09
U9O3s/bcFP9QrD1ZIl+MVEp3Jxbbk2oZHSeLS8eiHNt/Q20XZan9r3XMRAUHkGMU
9KsHAGPwFKrUVHITYVQ7WOw3xe15dFYm22g0odAwAIKGFliuNDSMFCTnsQ8XOKzX
53NZxO/Xvxx0rzJfMyJZqD0oYG7fCE2+TKJwSPBmICgqj+JBeKj2UK4QTP3i+PWr
X3sgWy1FfMOZKIWOTubdcGw6iBbBXqtcapcsO+34cveELXv5A37XQTVFgWowp5HE
g+DXC67V9j2fPoVS4quP/MiON2SyYGm0PSArJaPjwYCYZyBI75IFK1gznv+PH52s
RsFmPVmFio2nHkNh6DXNws0Um81p7Z/mdSEPFQHkXyqcMurDnTv+zrKiouojZvVI
0LGwz68jjQmhxv8Td54uYCi47d/X/MXSsFv+toA7pqJJG+GfOlqjbPkCLyXssaJ3
dtMNAf+3vYXJTNHRQBWMKRVGE9YExjuX57kHRzsq+47boZCuDX6SOvRX/kYioShB
M4L9pejiw60MIwIIVTf34UD0i2f7KAwr1IYpbzJmh7K+lR8/vixbqqIynSpxRpUd
HczecadoWElUWnjDwmDkZnU2vbf4OOOHJSBZalPNVzATTjuJzsVmWb5xlw0t6w65
Q3KDLRglDSqK32zmayVKjkFUdUmwcOrNY0MGf+l+tX2sfbVEEqvOuvHMgYvzJ/IN
NPvHCG+tvjcXXhdPLaJfmidmAyixYBETF0XfrRPCKDESfjC9NPZ1gwaOvlLplYeO
tvIpMlBbeEmKKMPyEL2OpnqpSkrfUd7KttDbcxb+Va2hqk+n0YLgPuve67BlY/AQ
PsS0UnqaxIJ88Fs4LMTGi2xD1no/GoPl/IlkD1fMAknrzKY903qw3+DI9cU73KHU
p8fro1cz+Hyq6HL9mQYQmBguu2hYsyOkXUrRL8usilMjFFVK/pPudW3sTAjJ6FK2
AlPw208m81vChdjdPQDfStIuWdrT2YCdRMniNBbVatVyssdVfKoAB1c73J3F38aP
ANrKGCz8zPZP8yPkX02aDCZeW+HZVIQsuAN4gJkncSU+uRBQsvLLHQIreVIn29xH
9uoOL45may4sESHSddyBhnyj0sqYuQzJ0kMp6ljJIHYXNTgRqvqpaHpkCWWNtpgV
B7ZWoJsS1K0G47HUQVve3y7UAsIir/oaLYLtEDVPGJvPGcU2/nVaLVmrdJFEVr1A
Dzdi2GzYXkqWtGyISZiLx5+/SX7Y5vEfJSH7GQy9wyiK81F+eu7QEp3wCCfy3u0i
kDB3smtsAkvdDWK34rms6fPprHIIeuNhkzdk20phXE8IQey6KMhJJZWeHBbPvA9J
VSfiWfxG/u/Sm0+oPUGW6YMkidMkPU7NOwfbte2Zf6/M0WIHn4bf3FBfKr1bFtdv
liDdFTnYuDf7sEwXNJ4E3OgqOn7AQJ+lAq9Ubs7xh6Cyn9s5spM12DKy1rUrU1o4
c7LwPompGbMJK8AxzaQaFCdYtNH+nNow9sqcqRSolgo1X59cD9VEhuHdEWO8rNjY
+1bSRL+AmlbuimzUNoiIkfqWgtiULyO8sWCBiFEAQfklrarXmi1IBDcBG3wNuOMq
YM0kukeqF4AJ8WD7KJYpKGPwLaYvC9qsdIlfwCvIV6f0VZImos7o5irc9FQ6kSaj
5IbSiFA+mfjXQkffrfe85UiqcOdpQ/2m3+GgKH3utld05/kIyHDrl9q4xb17fxVj
gmYSul84DEq1sfB3ql3j3sxM24W73WRnmW0DxVLIIGRAh5gF5xQtOigfJHM7qkLV
yztQRFxzhKSKwfv7r3YNhDZq0RRp0AW+NHo0FBH3rRAZ0pI+u9L4r3OMxqw0cHpr
5grdvWQ2a217GnqImSyWaAe33wXSobQtNUuUpcROAZLTCf3daeQ0wJDN9m5zv1S2
RGzygGHrqUFXIpR8cZ5ugd660gYN/P+l1r1GacdTuBMAzCZVal68xqLOQW4BDupX
hasYCozk4+5hylT+Fd9lcsTjmPV44oUxnrA7MRZhahuqMzVE2y5CX8ShQ/X/SG2w
+TZXCWA6q5z7npEs5DMhoX0NjpbQDxcDpSCrNJYH86Khk0+vDWBJBJRCZBgdkJky
pWPQ4IsHtDrLy6Zmwd6FTd/utwqeQ1oO5FHCVHpehkyub3xyACe9Fx9T5WjQxfBa
9p3kqQKylDEoAN2/hpk1tTFJsLEZhRFRvMngrr3Ie94/kD/O9eluS8SoR7MlAQmn
QFmRztwO8laG8vaSZ+EHayUIMbksqyEUANib5DTpS+IqM8JxB7mhrhU14CgCgB1o
aNAQKc/DyVn68SB+ntKrxAKRB+x7SsGEsriRNV0bPJjqotVT3XSqco7B7WH+324v
guqbwDiE0uPZB8ZkLyAHzvq2WK4BDrEOfMp7EOWXKJbBdxpRShCg4d4Y257aPMyW
3kEnmzpsWwaj9cvt5PBpu7Twuw48tm1f7hAkpa0E0PKb7E1inuI29un+T/DahrIN
GY5oAqPoe92wvuqcn5Sto+8VXfp+oN8/2vov5Jw6iutI4VkjH6bZ4L62ZqyDAmfQ
ze5QI6zLvqf+aBAYudPclfNXv3qN33IuxmjRm0x4nhLDgcF5oFtHpzMa8GVL1c8/
aDabycSOcqgtmbvHnXru41f/8ZOqxGzfUJNQmMMA6CWg9th/U91FS2lfiKAxgIwW
AbiB6ILw7yvvX4Oe4x5EeO3IlgN2NGD1Fyy6SEqRhteN61fUIDj/E0TgJ7MOyo3y
Mrz+yeNG6YxPc6Uab7LQFKeP11odqAIbkHxCideoGnDPwdLiCuNZsR2hw+KHfx/m
laAdZSQKUkPohwSGVVYwd1SIepT8aB8r9Ez/gAkv8OtMVACv5D8W03c3S8CPBhwR
89+XlTzH+wgsoy+i1IvYwXYpS7GSz7A6CO0fYXoEJdUoEjuJTuM6HD8iogeDNsVb
QyAU1MAX8vYy56xztGyP/EbQz8lcpsmbEx/E3xCX6C5Xe56LWRHz9XwtCoCmCLNU
PCHtYqmjUQpQgsgtZNrnUyHR0/KN5BinE1A4oNTqItc5e1xwUCGtDRXJOEN7Dhdp
310Tnq8F64XZjdQT8pKfOFaE+jIaJ1hX62vqw9AA1smoWTqKOGzgJNhwmOawPXyg
ypClZOkL3b7KgDymGco5USCqcfIBZR07GcqC/b8k84O7BcYjqOpteimeNwjzsy+E
wioefq+Dnwn0Z+3KOT3JBaRlmXEOulcUgBjrea+qIrw5LMa795wkQ9Wx80ZTTeXZ
8uPSO4B1v7bF5m5QaiE50jwjPouzBpEZVkSJSNZVEj9OzYT9weqg1nD4MQcDjm/1
/CcAhUXABiBaOaOuwPiM9QfJ+m264nNdj941XcmMcD8hJcqZo47qBBqa/wiX3nYz
tnFBmuyvyD5Du18UhCyWY9WY7nwhuiLGrwo58Ab5egNAd59JwyuBm6Ep1798A6L8
iqs89eaQVWMoQIRcKd1MTdsY/tqopOS70V5nyKtj6E5xrm+nv7+yfyHbZa0rNibd
Q+0s+66Bv5dc+cB3EDjOw4CrDFuWysC7BIxnDEJItZ2w/XDFxE9IFt1AxeIz5ccx
rkCdOsso9K0PP47MtgFo6sap7YkxYS5o6/AAc22uQNF8oIVBPvRk3c3T/DPb21ky
xwJI/0TChacbrQIvAA1yAbYCIoROVCxOYO7uo9/3RKC1rJb2YN6zK964oqA9kFYl
rxZv85po24eAg9LBuPwylqt4cApWTnouswOeVcSy4tS3ZLSc6iITfEOW8KDiCLS5
fEVet0B/yQuoh8VzegfC4tUEjNOwEFlbJ8a9wTLEXY5E+wUthYRx2LPeMmrLbz8n
F5uVBldh21Kk2w4JJPX1+3Xmvm7H4lyrFTEkkBbq3gC71wQBTlbSPxPBZMp8Ew5d
NV4Db/Ibg0evBJHoFvnjt4b0+OLKyZ0t+SpE/EW7WdwmErGwq5LnN3NH4oDRS23Y
4zMeWettHHmBZzuCX/CPIpdoNf/k9Ziw3nLqMFRokImrm3Qn0iHRr+Ulpy+4ZBYO
dHwBxiNWqj7EPPpUy/v7XDEl4o6bRHj2hNwVLAWBKQafCTEfmzK9zOJZDYOAVoKd
OW/O7ldlgY2/p/kN3jW9nqLvGNh25mSv7jMKpIs6DRfeLPBfPm9Ks9ynviwrKPZ5
/8x7CCyukY0kJR615EAgCeET0tYUEabNLEVN6PC4eopUH/nN/ZNIuK2BIPWDMWV4
7eBpDkGcZbJGBqfUjctTyQ91a0N7AG2yYSODb48FjvTzkU+ZvadksHxCPcVxcFdf
uLscSlYZ5ySUabRo1aXAKcme50fKpFFEU4whAIMdw0ycd6/apmV1ulU5zRF2iIBQ
sTB4e16pbGm/rlu8E92gwKeU6uQjL1je1qp/g4cnAyNPRePVe03qmcczdATlhenh
7TZI41/DABsePGjUIbA9XafX2H0F2+LEOpuJuuFvFvEB5nl6Dn3p0ZMJng8ZyEZ+
KOd0b34cMD1z4bYF4vooCY1E4Kh1opRfTdxz8gFlMwtJlDTXEIF3jmzJUHlPxztj
AbhHMCjE0o6TRGxKmWLHjO2UiD53Mohp9mIQ5g4v1l+Li0ltQvKZbHm0YCupKshT
gP8PqetSzwioHz6EfrUXpHRK0u8gx4iizc0tXzr8bHbw07uj9rgS9z4soWn4AlWy
w2Dhe5VOgUbQxJJeVHKjveffaSUBHPQiU4rlW7TMz9lDUZAtz9jdgfG7lO3me9bO
F7ysXU44FQFoaDszVBEsfxO9JI1yH0y/IpUfASHEDIRcpGl0Tlodf+04uMroGeKZ
YZ727VOJmjPEL8GcfYwY10KQUSmPseoOhhuSvIi1qUgIBBWpGGkXVlsIvMMfn9cm
hPK2N5Pv9Q56ZGooaBKuYUjhNFqGYIAqc3EGMOrCqVT7N7x0NoHqExu6xKGDh20S
WaJQfiG42Yc37tAo4+r5OMdXTM0+nkfo9c+eexu8osSeEq2jaxtPwcBzUGTow2Ks
TPd29UEMDxBcYC9O/C1BKp8ciBcPrF3cUPh9bZPxJU9YyvKIE+tpBnVHfd5voLrI
zVAVaDc+gv8TP+OlaEDX+W1+xFUyEPcpt4jgken/bRCsy42PmErjt8W4Is0Sc08C
TnV3pAHhs1eay5vfZQzuxiZR/zPt3c4PFeLHwelvF7zvXVYOYmCy6Qk5IiFiuGf1
+LUBFoavPTUJukbTE57rVdeaKif1SCOzbbwUTrIcRCP/wT+s1W5adfAJCPV6pSUI
C2bv1jJFR0ZOGv294YWyOFe/5Bl4lJtPkymwwNx5kg4WE13niqnBUIwH4E70kdx7
Aa3BYgoI0Wh7Z/F5Dw7Zy/9Fb9REs4RMlvHytGKaCen3qkYcs1s7xkCaWVvRnRG+
Rn/DOQsX6wW8I7orDuozILt0nQnMd75X9suTDU86/NUAk+NNV7yMfaq5vY5z2K68
FQ/uFvORPGh6d6DMngv6xKVAVREBmBip02xk5u1LmVcCF3opRYIBWJ+22tvy1dt0
vztRGnwNxHDf2NUZkZT4uZXH/CLjgud1eipJrYwtAuOYQv6e4er5cswBtXIawwqq
XjR5QoFzhONImOUyYE0mMY0jZA0pGpqOBbiLkn4om/v+k4iP0Dj5cTrPi7mGXF0z
VKxGMOBoHyB+xjLMhozkIOIlMhFePqUOKikGHmLDDNCp/kkRa2XLBrjf00zwIEPy
+b4y5/TjXjaSy3qWY5l7PeYKMbdVRiRL0P0hPP18Hd2kiHUneiaRu/jQax97OMcB
XZqs3PYlr5kZmY/d68jmKvnY1ZJCsU0g4el3zkaLhPVXBhEMk4M8xdiUIOKtQC1D
9vWmHASUlnqTALm4mUwjumMixjsGsXKR54u5Mxy00WMIf6vBpzVpftdW3Rll0N0B
b4PIDoRrMWLL/MofgN7Mg0h4UDxxB897OacqO7ocw/F8uNQHFaafHxKGUI4WTy27
yrz5xjC6JJ/PUKd7M09jk2mTdCF34/wn2P5lKQqU9zpUrwu8ZO+scYirSok+8FIG
+kyLQuLWouEESTZQSF/6srWmedf/YfUK4UhUDauQuHoOR8cY7ifIAoZGQsfuvzIo
8ohO9y5d+kB1BXOLKeZh+rmBSn44yIfiHtBYCFYgcapYVOdPObOxQIZ5l6hkqn3J
aQyRvJ9L/ZJporvZaDN8TZyoV3baRkc4VyWqQl0RqqAIoWUnDWF27A2rz2x9LBG4
Wvp/V2WaBUcGVdnPsKNNIMLFBLR7iQjppT5qecEuykVFFBo2/Jmi5ZTJNTlqs3Q3
HGhk4NrN00GGD/5ZSbh9moyGGpvBSPGidTcmvKHBM4NlXzXeMAQh2s8C44pybWcv
9LpULD7oObMoLoB7AKBQgNkkStSm0TrPNX8eXsF2Fu5H4tqTGsuoXt5Cr5xUzQmr
krEnecD7WIN9iHyqIYlQQjeNAaYSVmW+0jcdno6ALSwPDWJX68wZ31wFkFfOS1tj
t3YeLtNdLUaZs3hBFupweLgXek9nyzTBLh3iPsovngLkkApCXQDIvMfenwA+LIUE
+14oZJ+sa/1QV2uoz9klz0EnBNQ8jH1SSPUa6gFMs6V3NXFXQTNO9jrcCsaTymEz
HUGTtA1nmsFdNOk5kw+uFfBLPe3uAiX/XPKXBzG8A6A9FclSd0IilneKQUBtROvc
csNTp6L/hdky+eGcdu9rgF8nMjjXi+mxhXX1WETu4MJEmmqnP1K1N1FYq+c4WKMY
BTHEVLoTar0UfExHTBXJEog9aNYHSJmtGBF71nVBCJdny/M6Fg71W8Sv8VtuxcNy
c0zV2W53+V6a+JtFYJSI066iKjf3CpOyN2VKB5IIxhY0qYbIa7OS1A1ncU3Km2o5
UEGLeMrgxlAKlyZxgsOpLrXOov6se/3azU8BTCbA+g9DuXnWahL4h6SIw+tp+11H
dc0qrEj++RXjFV8TORG4IiXnVa0D0fzpCupTcOWLHlYck2jlH8mGWJEK+r/WeCcp
JIQF8wAN7DlI0bSXTSyP3pmS+QZ3kr1bOcSv5hvQQCKBcCzsn/E4jd2Ch7TTFnTp
/TzgDaIvHCZgG/ooJUDYjGlAJil07+RgKA4YNpHAs+x1dh+eJ6o6dp5O+YYjPepE
4xrlq6fP6uzU9cHfkP3dlzqFbNIdlll8WbNCqDHuBtJkOPWlSVU32zlb+oqmhAtZ
iCd+I7t94VDPQ0QZwM/iqAUmf2oGlA1aizj64laWWUav3jrxrH7RqYzQy3CURfsT
82VSzs3fW9t+mcxMjSDPopAm5kvj2ReJk189fMx29fliT8PFutYywcSjBbOubAZ1
95F+Tk6ghblNd9XM2ibN2D6DNkLs5F46/sCU+N6RIIh1r359EqN2raFSwBrvB+mD
KMBfmb+BVPscPomM+ORICC2vwHQRrUAOUuJzHvmcD9fLPkmM6iScimA7u2aLCHYi
/SaR2p4zHZvcyHOoZaC7+Py/ObKTaQGUo4apsfgleEong/WjVXrKkfUA/329x0EV
VCX68BMMU79PoDLUSKSxcfQYn6goKlmF2ll+sb7AI/IzRgFLdhpl6LPl8SkWEqCV
N325H8QwtLreZ6ZDX7l8NNuMESFFKAbDll0SIJzzj/T9W04Y/Y40EgCfIry8Ngkf
RVUsDORxYa0+lYb9EOnPUXgqp10xc4dX9ZUyL4cborwe6nRhbDbAVXEGVYjg+Dda
6dd6KnltIUBhXJpr66f9a7USLkx6++YT6+LV7L7r8iMdn3F28LFLb5YPcNXJ0Tkv
fuoka4XC+//+xSZHP7N9y6b0BcnJDALUgfeasEtY7ljbPH7FlXpMfciUl/Q3yDBU
MRy8L+R8POnWFYT/ji6NnQvpXD8+sQ9v6efX9t5nway8qxBXBJvNe3Q9yL9YTPwc
sPcZc69ZcApr++pfCateRsjr2Z8qogIo/lNTFRtSEkH1uz1ClsoEkBSTKRYACKOQ
ImClg/4AkYx3agXBtKSxd0yflZl24wVMmsdh4kJcFaOMBmet+9OjA+Z8+TcwL/1E
S1nxVkCmxJTXeIXp67rRYz2ZB36C+tylV2xv08pT6I208AvbPTroVNwFC48YdQ47
zfLbSHxiBR0Bjw4ecApRiAVum5QZj56zboqORAtot+/qMhwgwZyq8K9vB4kd4Mn7
V15BKZmRBBAt4Mhxc02DDJn36hSM79+/uI33x/dcHWrCX/NuKXlH6GP0vANrh0RA
qu4Da7d7zDmH2eRgps+TkuLbPJyFdGIN65VM6i/FXap1djsYLkctKaPxddLvQJ0+
hZWJXIWlk7lIWoCit9VPtUsINoZv0LsH36fUqoIp6a+uV5R817MlRC0v9fDblm/q
EuxDBNkewzSQGSsRtlSBPIbj7lCS4ZL91zCUoKQIAf8axMEOXHzVGFv9UDzRUIAU
MZs+xg7zzq3dWsYVM5q2Pn2s0wOhyf3UoLRkVktudUZVyI/dfiFDCkPPfHgyer5K
EVKbjFwfLP5XvSkpTQkXKH4xFZYHP6SanAWoYH8U79UEQbQJgWM1Rf4sfTTnm5uU
Gx3qIILBdp8LVrlB5VwyItHAMlxovNcav9vTvzmfFOLaJgz8T9yVTIxX8MUpeq7s
uyr+Viu7ryJG23tWz+ydXvdI+STFjG1C9hehpxNceyJq4OPNc/7viorQ4dP3Y3h6
wB1I6gsLB2+Bm2PxlT5xTneCqP44E8yTGRfq6LB0V1KGl58uFGASKkgm4vJbpDq3
qxM75gai+vRXzBRQUYiNG+USi7x6em/slNozNhJWtgB0w4SGwnpTkmpd1GepqH//
O8AqnJ++hm1HahtBdXey0Z2HiunkQiqM8iumHfrwMil9IJGRD3b6Ewsp505XZR//
EgptsdDkADaMNNIBQTG49oIlEhM/qfBC/ijW1p70bOUBCObfu8QfhBBl5fMM7l1U
XYT/eh8yvb1SQBgCDn5b3oPYb6riRLw2JhKmQ6hF4v85CRBE0AK34r3/gFiFskSb
13xWabP7JZRvs+UY8lSCmMXSM3QNHTFW/bykrPiyUmYw3bh2dJVqK6IqEB7V6Akx
r/LqF1S4kx6vEU3/PuDktzfkmD9ItH807WmOdrhXeiYtNZDdygCwFnIErUPQmDyB
lI35StsuC0OfUxEUJSIdBLZhr3nAX7Lg4PJVFNH7t99/QiOnjxt2sZOGpozrGmno
1nfQgP5Z/bygMMejpe1ojhVhf4PYx35Zr0YY8/gEMT9kPf2eGQ4hBKfNB9Bi01sk
mmwAJof75jB/FXLgsMZXNyDAUgoe6MQcH6cZaqxZVoTJp4g2/Uv1a7cEhjWdp+yB
0HvAuN0iOlzR9Ca9jAr/1zwIL4s1YAP/smy0ix/ZEmnXjtN2qYfxfHcHI13BlbDQ
AevnAg+QIO54kK9zDPc+8AXcqlqlVJ2V/spHcdSH3sFAWvdyh2Tq0TabHc8AscxO
IvDVcJ3ZjeLmnmuW7vtg7nk8OuVMd3ICXUjoi4drHZ89bOQT98F2yAoM5ukQDLaZ
bbAEv5+j0aqlTpwdfTLr+/xGJFN+L3F96ToIEGMZy446azti99KaoB1oxz2V2VGZ
Zj4o4Tmvb9Nb+1Rip+I43OPJP3zoekKtaJUGAxUP7EWmEu29/3q3rvTYE2bEZiuM
DY9WQogf6oCx0W8E31ZXOlfpVEYmdPJ5Drp4XZYtIKpMWKR+xsYXk3wkxjrI8mas
p33106IJD2syUrZdamdMUnt1XynklM2JjlRlU5VP3y1odgYK2W4WpOdxTzbFqaxA
UFeHUjaqlNrn9rY0iJqVbqHD+1VRIVFeWVH8XuimJj+eCyGBLJzeGjsitSHlljir
2Bd/qBje07U+pkmIsSmmZRHfC8GgFx+4kDzqq0Xj+K6MxdmgKLC2A5+KdlXmfLyy
yGQ9zE/7ZG1oO/WS+SPBZxH0s3MdjjMg5nJ/mWveoW8XxiJ3327ymGpwW7AwjSKQ
b11IWInehzp9jBJEQ8w7VAmitEtU/Y/g0qJm/6VfHK3BYgr8NiN9iFXIaCwhcr0d
i+b2EBsjk8drtprqj4qCFV2BTA354XcRO3Um9dKbCubkpdqAl16Jov471IUkXelC
NIBNjfvsS1oND2OHLX9Y7P9KwbI/6THB7Zmxn7UTLCCkxFAoxDHV4408TvywkNtu
vFVQ8sCYI9kGAB5aGEXq+i8XKk+Agi/pn0qXUWqQgFujZ/4nZe9UVy/aA3WtIsbL
6Y/wrLM7QQRkNy3qdotO8RyjVCRj3xO87Pa5KICCK8zryKOp9S1tCX+Aq/sPGBWY
O65VWQ2UiKpU/Q6iutCoHev8aQAq57yCEE4TTMnGbwgDq0iddkksPAno39QCoYut
8CNlt+NjmDJ/1blBA5sfww77SSxgD1YJnWf0jdzXUfX7FSb3LhQpV1GE4rIEHndW
5+8rbceCi7Ui0ATCVAt/ufGcm6S0AwlZLfyX4eXoI+Dv++mf5tMQuhNc0d6QDsxL
ndM2Voex8wrNnygO7sJyS9ru+B8ofGtRI8ruWYxQuNBj6hGxSjpoLwS12EDkqzPB
DwoxiWNiSMDpfCYzFSfZHD+IXDW0i4ESejw6Ou70oJL5XMXo3cGv+MSLlB53AkA8
PSnFvBBVak8LExNwOfCQzAEd/MO8iz2D2WgGve5JcvZ2JX5vZ9km2WIHC1s3t0wi
eTOjaIWT4yLO3yIFRF4CMQNBunCvpAs9zrqeuJz4vxIBh3AZOM2HjBmRYI+EXAm2
Z/FmUrfSM/hsP9ZOtqYPZkJobVyZOlC3d3yVQJ953a1hpDbksbbS+XkayWANtCdl
bu4i5mkP9B6DID6FZTYqZo8ClvE8WUU58gf1BYgrTtfNzze9AQd2OnJRXd6s6gD1
1/mD7a/pPnofGIq57IhTQnY2fwQhYxXTqztloTQ202Ja2SpuHggDp1Z/E3GhYk7a
YwiyYD5EdnWTvFpJQr/1EkRZ8b3EA0sNkEvV7ak8oXcG39gh5BtWgoKdMBuC6UoM
ejYUNUaKAR4pFV1onSgkkYNEHAjzeMciDAnuLhHlNZNQfZUaverXFvSwePTp20L5
Xq01iu1qA/IgtZuDoSnC5QykMBrXEgOuCNwY3Aj/V8b4NKox4JLAf6yef4vJSuuG
/kNsfjz/kCBL8MF1t+XhL/e5ndpb6oFsmFkm00KbGbGUGnKSnDqPyoyTUWoeHpoL
/cIaKswT+oyrnOGQ4frBiOmNTaf4YWa5PzInW0i897J0dx3Shu8ZtMYpv3mX7wW5
KXF5a9XE+tnZ5mQRfYqkVwDSp1wx5i6YEYUTBxR8q3f9j+w+SnV4KieyNePtwrQh
//BBf/2aSpzq0GgIGyScDumjQht+/ZFze31jol7gwbqNTtiqVrx6IkMmbF+6ytSa
dHBjYYd3OYrhAQ/sGlIl3ERyrJzqOHEyX1P5F+Rf5alny9jBMr7ctpUcWJbNwUd2
wRwrcoeSvKkjHXqJqjjvebs3dOxZkMQajEpkDPdHDdFnk9sya2D2L8PT08t+GSfK
ywSY6n64FiLll0VaXEFAnaAKbq2MtY+GrYbknY+/Cu6mhUYls30cIunZsWrfif1a
OmxhvXuZpAITxk9FpuQ/MosNlaclmH4jsu2l8DTL9EY5kUbFK+S09N8vCxH36XFK
B7H0s9FzOFQy/JXVyZQuoQYV4KE4Zmvo0vLPYcHND0OhupeGYINmLyG34vhJtWh8
gDT0esK0ifQfJnh4rjmQazAwJjXOCik5VEAIJ13F5/no2puS5mysEnqdG+U19s9D
DxATChnBYXz4NvB6t7/z6IJlEWi9/3ogPO7AobJ3Qy8bJ6X/ycu3GOYyBl8Ow01o
+iBrN70rfvXodr9eSxDyjZX78R6qHJRN7JYsV1+kZTuWlX74LxmvT2s7jX+OKmDR
KiGO2pt7aOwimo/KwQ22eiSEOu4OFsugRYXBOfH5+UIOPzaK7g7p8W6K/Kz+z/UX
PXtfoyNBrUNkweUFuiD0MP5zF+sUCZAYKQkpwiJCDa5urVgjcDjpeEqWPHrFAcPD
PnEQUBSyfaGUIPv+xJZR63A/KDn3u3tyRgQq7PCKS/nIWBpW7IlImulQDGSq8XdE
GgrQgCF6vqWn/bOfE0BYxuX6cYIGeFAAR7zNH8WpAm5dtHGPKuKrTJ6jU4fyGenv
Aipiah5WZreYlBTtNFrEG0YXyg4SSaIPay8jTprEWb5c7qeYbRalNVtp2g8QvGT7
fki5h0NqdW5JJAhDSV2eIRdu8Occ7HngQd+NGpKDRReDu8GZsSWhgELJrY2r2NgX
nF8r81BUQ5jLcxJmRZ8MRDrsv7gOEOgNrNddzBBSrnWddiacnCobczB0NCVp/Mh+
hNpLmXyK0RRc8iBBmafx7z6PrApyxQieLOMTzcaw6MmwBbo32WUkF8nNrZdUas5j
IEBweSDHFsFjKzoh43tyP5tj914MkUXoNdWWSpnk8TlclrfKUUCoW8rTr9rxKp4f
9tAdeKyQH/X84mDA/e4gQpz1dVrbz6WO+01bBBYjUgpe9MhjIyuYSeqpE5WI12aA
VUPJwh8Kx+cd68qxNOln8YoZfAnxk/LXX2YuLhIj6V5Kx5foqAHkqGDXqjNKfF6G
fu08ld69I9qy8qPwbUlWaOXptcJKVX/pQgWzw+mVB/7YcEvqX0kfAmpkJQUU0JwY
B/TKqGDdYj8b4o6sXO/5x3rVPkyv94plOdaBtuYRa5hBakNEKLbPSrvbGyS+gpk6
Yl5GXJ95tainIPO/FBw1SHg6WS2fVXdgfG3rm87D9C6tVN5TZ/hRzPhVFfFtwlng
jju0oMW6MDgOtempEa1gN6LcH0ZCpq1fJrxic8aLBc9gw4lI6Nlebd0VyoJWo9im
1wL3QgJdaj17Xzv3biVtXoAKq8URL344ZZgdKyLdw8jFiP3Oe9LHFZcZ+ojCaRYH
cvehZRxAf1bnKSNcyDszx5vg2oHqkOEqY6KOEApD5Yxq2gd9Lcoh7UPkMxlMNwiA
30L8zbb37nIwYHYURxSuMHRPTOU/KUXAKHeKo3auNwcDyjxbN5c1NHR/csX+jWTK
Kgm8SlnTzL21XfRB2mGe0oIHRtwmSwrvBf4A7Quix2ThSgp4UF3B/4fQDEkEkXFo
NjWfS5j6ETsCJHaJSQGrD0eDl+4i6G+EDf5I3jvahG7+GUWMOdg++I9lWaolrddF
v/Hb8q+R2zD6WPuP+WEVO0Q5v+dSVrwR42029gTL6Z/l3PSilQmchur9namwI8Q2
tYnTRpIvD6vesy7dJ448LKYrpCRN2GAKhMfdsM9L1/jT8Rnez/BEMTE60piDmMh6
CxhVDbK4ljeDYqCfUcPyppqaSVt0LTUz75YzHFW/4FE7o8bGotmXqCzSAzXuXSGB
hjuPFI5f92o67s4BtAIamCHSvBrhsMpuvoX5jiQ1My9ep2YUGdWH8nlKhOrhkYJk
yHG/tK4yxn7Vb9hwK8P25vR1LL1sHhpvX/sr0lzvf6TSkyJH6PiqhUCtYod8x/SH
963HSDRuBzOovq9RHWCqFq78maJ8jbMX/MskhGdK4mRHKrola0rAyqDcERtxR00s
C4S3zWTRKggl2r7y/JNu9l/HqASB9BZxcQ6KgEtmMcutY+Fgq0g2zSJreI88Y85J
BLfpc7/qVkXbefcSNHf41/1hR0zk6quh4TA7lTgGWk0i2mJsJTNITII4PXV4JJHa
aJLh3ti9e3vhI5fagPZLnmx2yeVxQMK6Rux4DdUspR50HXKJrZGD9Cum5nf6wjbc
4Aq40muc1uQasMiTwQyWp7jMNOc+lN9C5FbhBeTFJcshsS7by+GsLIP06gLh1YaK
ivDUFASSnwN9iimOlzcPZ0Hu5TNs+jkhXqqxmqixp0xDY/8awzB2vNhF8XCfDVSP
CqKBP9QD2j3oBP3oeDdwHXu38y9O1/C81AOkzc/NwrAJW/+pvqOt4uMzsnpRvVaV
DiHBNxT+TYku8rXShu86mI9U85y9tVJszaZbh96gYPFrxMYenaa1+yO0khj3BjJ9
7nd8Tisa44rQWM/+butltjbGz1NolGFF4MvClbUa2g7y0qwaV5HKpUB9WzbzeO3o
Rxo7K1Ydfq5p1uPaj3/wjPtO7ROuA8X/yoSjQG77bQh5VdZcJix5GTmxXsQ5BePB
4eC7VpQBa+7oaK4KGx0oSI9u6kzbuGjtvfOKQA1StTcOI1bnaY3VWBPCDmKRoZeR
FHFqi8+bvtOd0v3XAiwGDCjyanLt5+wxIP7L0xZSD7G99gX6MuXsjl8oYFubKUkT
0kGLiExK1PixMQ7MChENe4h4i2nISML37129o2/NgR9qwMxQFAbUsDnV8tZxf21g
gs9IVRDFxpK2m9MY/WQJlW6Ws7HIdjhwd5QDZjL3HF0pAEwYX+YBAmXlimX6EkFj
DKHsN0YOTKnigi2pfZHYhLvqz1nJ6wH/eBEmuV1PVHl2tlHpB2D2nIYbjbNoS24Q
RZisn3TeWvwVPze11TX3z52S+WhpgBCn5842ePtykgyxo4vM7MC/ZZuMVoNgUe23
dQHo8a/6z6+6Fik6I7INgg4jTCT8sknCKz7OOa3IYcZNElPbsjVSsYCCJWiXI4kz
0ahAVDfXE60pGatBS+3qq6bdsAMKZRCm1T++CAgkvDwCzNfgY6MkhvUNZ56BUwOT
iNNm3HjDcaobCrbi/5JNY/Fw05gVIIMlLNMd3Sh7z057a5GMZEzuYHF18j3dYNA3
GZVDtRDRLoUhbhq1esjjqUWDVadTjqH29WW+f7ouDW3L49+wgOhfpK+cF2nAtIb8
53PcZRHKrTwf2ibe3nNprRpRRE3yN8vkEkS9Q73nswbcJRbzFxm033ePX1d4SxfG
MmELP3ytf62CIwEaPQ6vo3Ao5d4GGuS66/iDeP+tIq9Ll5ocp3SMbVTuWKAOIvhh
Hsd8oH1OVvf+Wf7MAF9QbJNcIJbowaoMlsW+68GtOQlCR+20kmb0SZxRERHYIHCv
49mDsdFWQOsop4FBt9wenm/LETQzUarcVBaqSsadOlS+cQc8wWn9kxRyHONm2TFF
ZxskdA+0UG7e0/txAMeobeQymbQvZEjkSvQ5Sf0ediC8hAr9qiMdWyPsNSi+AwO5
83pJqhi7svO1nKfgtxt3VVb3cohiNf5vW0oE2A0L59IqIWBPyvl6/uQY076fkYPN
YfD4bfnMCOPY33LEabRUP8pQw5P7lS7Qf1bExAfLcckBkZ2/i4ReVUqH2qaGYk41
KZ4L83Mf409JvUm25xGHmPp3CH6y5R8do0R/9BqLWn56zYHRe5eUwVrNDANX7p1s
SmpRmGHy9DmHdO/yL/Vy7T4zQmcBqvNHyWEJkD3YS0Rl+1RLwav3qxynsGN2wvBF
u3X7WtzHPbF75PVDIfCRRde4YdMijrThLH/cmsbLORToC3r4lNYL4r8moc5adKW8
jM4UAU/GZzSv63tvlri+qb/CVrIgFXRmYXp57nrL7aZ2ee5AevbzFPGHjxKLuX74
oPNSoovvj0+tPoD++wkVIQ9FQIdDVw/GoQq8JsoIjT9DxNi8Ba/iuyPkAAKhMPSv
0aLcsGps3dlagnvOIOp1/rtQJJnHNMY/tOsDFTgVUfMAK60+r5MqEwgByOJtScj8
N9uu23jw8TRekO5n/IFhUY6ri4AyZkZRg6Wul8f2tSC3dimw5/AoE9kNewZsMA9R
Vq0+6YxipB2UpYqNmKhIaRbAudjMAiDuW2htHe7sn12VHCfMDSGaZZBks/iEH0Zi
sQyx7JaoMGBMY7vpSTlEtJRGq+lcgHVcHhqZSyrN/L3rb87RZY7jC11qk8T99cDK
Oqjp5sgrT1MwcVLp0w8GwLKU3XiaYmCj7SeohVs+7GTUBy6x0+aZ4vNXdQued3W9
p3yh3H4HZCCB6RXGe/w/7llIMcuHlT0XheCw5eTl9pnndlNeJip950q1ivAjPz15
g0ViQmbEcnnpy0glUTgCWbZjKz4DH1hNN65whZWm2F7Al+uXkDhQhFt1iyjSS3lq
+qGG/2Prx9jTXvbeKcMhce6axn/k/rKG+nuYcl57glt02uCKi4g/tw1qQUm8qJ2u
8cNPZueWde7FsFQKgezuqXiriQtuh+PXe154/gK6ZB29ucoAO/U2XjDixXVKYVXr
Np5YJR7IQOF5w6nRnaIwbrhQfm9X9tguwajzU5vhDPzESZJ/iVaaoq+h4tRSOo+r
kLggImRVXhy/Rxy0nkJ4uMVTsoN4pU/hovGtsN94p31h38GbemTQ1QfwZI4UE98G
qzPhWI3CL+LfiZeNNRHuxt6EP+1vwOnt+cP+H3Go7zlAU+XMK1Vl4SffuScxm3GT
xIG7zxKA7KKRKtKoYt55kGOjkOxFd3w/TcFiKosCrWDwTNAnjoNmmH0hHe5iw9iJ
c0kbRYKbViMQDDIho3S+3bZDiqmsvNGe34dK7DgfrJGZ7cENqFdAQlfLLxtoOydb
Y4BvObi3DWjrsxOXFFa9hPpyQMi+IjUxXrPTKu7jLMkMDpSHaQY7Y26ZWTTUPgkX
Tl5a1r95oSsbLqaTQJfxSsj5vmCcmj8hFSKu6X6WLqsrww4lN8p9/jDGM3UycmpV
+fyP+zNisz/fyjn6wECxW84zxWfDTAIPbQEKo/RajjOoCcKTVdpmaUDVEyu2Ejvf
gxNZebpaCilKDSBWOn12u41BkzsznpJ88vGzfhGN9bEcUtaWtc3H7SPakkh5KwHr
C58rSjmM83/IpuLUGHvYWIABF0GeZHVWGyVyeIlGN94OjL/KhJ96JYrwxKBW6XsS
/yi82oaWoqn+nK7Rlqu5TkIwUgu5oa5+mG2sqwrj7XQfuYD02PNzZMzsYfAjB3QX
D+kI40RP7/29lmlLOTTf2YKCWpx9I6I8wUWLGE+B3qEYFooZsvHS07luTMvp2dXO
Da0kfJn0XQ1+uod7dLB9dDeoDechm1a1P9r7QJZnu8Gg7Upb2y7lMV3rIunGT7RT
FQBdT+AB3XuHpJGf/ERQAIWd747nV4alVUg2zg0aQphcPZO59uh8um0faxVGwNl0
zvl3evT+Rf3vZ0guGsCr52NH5efCsDFr8jYXRd6wQ7jxSX1R2AkIvYv5vBoJHbDa
dofbIWiwBFdmcLbKo/AI2DCwT+bB0h/iYpfRWJyHz6GJn6LW5o/+T7v9LTEOEXmD
Jy1+BcbqLix/9vbMiPrecIFYrX+Oz6eH+B3cdYsOcLDSCH0j2pSQTp7WHBIgFJsY
Xd1BuJJedxw4y5cmAgmOQaOXELRk9zmN28/zaN4j/PZSv2j7yYIqN7TJwfIExFjv
6khv5hq4gQ/GbGzV2We3q9PM2GZuMO3/9GXhTaXS74fKpm32jzUPzFYagAo+HAYI
4zBnI6LRFclqhqs+ayNyQd9SbFcyvyaW6wFdD8+t84p7bvjxiQGLJALqxVB+MaK5
vIEWhP1qj3jhPTivJyMvaA0mZ8vzBu9Evu1UiSbJ3x1iwoJ6gjlrgNkcrliq4GK/
dkcD+IE5t0RDNEapYxbEwQ9lFYQ8YFo29ftP6xiJr9kAfJjYIccGE1x8w+LJ9vl6
mKN1Irp+5uLs7aBsOFkLopZXRc41pKQ6Gxc8dzABRs4+2eZp/HxxIlnP8+IqSH9q
8f5qr720l5UoNKWHsb2t8Nxjn1c73+Bv/Yojtic/jh4PpY6jdYTiXc6vfbXPDWTM
PAv3ceHRSoyS0zD3JHg7C5XNA3W1VlUkeKz96HxxTMTgqF2WY2PPQad061fXAQAH
Cq+6y+3nqvIQDu0Uo/kZiCRbIK79VAbYyF/Pc3ArMTAIg9Zr5C+9UVR2b2uEQh+4
6pMjwaD+TkC9Z6uHN/cDQNNaLvF6dQsctEXeoJhF5t6nJuriMpkWA8U4E3rw/WPb
dkjKzxBRe/aaFWgp3C1uLRuaSvaq8lIujptIqwvYUVYDRGpMxtl+LbXvy5RjA0r4
xhC2PWtQbvFDyGq21SpeNNwzMugRxnkGZMB1QxwGTGN4ApFn3TwzljfuVkXlHVfX
yVpqnPK/5Zv7UIZDUS9m2+bEWrbMywfOzoxT3tPql8lVvlWAlewbgzPjdDbMS9un
9FmXyS7AnvymHV1YVi4NUS5V48szHW7yP6dPZQ6wpzbGa9pKldj+7hDPqOr2YDCy
tXlDZeH3deAFYrQP/68xM+DznWqTSIlbzvCzFAFUdqAThvzpKVPb2sZMKexflclE
xRuodUyECsdwPkdf4EbbCQC0Eu6ON3vf5W6S4PQ9LIVGSQPR9KyMY1FcOuOtJvwO
SPWkgnHOwb7BLvgARodOvLGljGbTSCxH5CRjfW1+zM8ULJ2LUpYesImj1m/NFcDB
mBY0vIaOOnadsRms4fEUsvW5BATxTMqtZz/o5jRChGrYm3YleVzGx6iwe4Uq6wYk
cLr6WamMFE6mfhRECYZKPlzeZkVw19qiNW/fUSOqepbcHbrHPtAYERUpLjig2ynL
alME8IUp2Y/14UJ1m5j5XT7BvbEmDZyAvrDzbg325fJjexu9PjasGsoVYmcl9rzX
DNSdAs7KWI9SfzCYzWSPjNBlQAS6kudx5VNol2DwOugvgew0pJvD/E76du7N2xJd
ym9z+IW789jtkzV/ObU2SExHDHysh1euAMFOPenytbn+iDB19+A030uviW36a5Ot
82NrLOxC2km4F4bRmal8VU1GC9YFEAVLJG4QqIpS3y0l0V/Ga4MmPCgc/LYzQg5w
gwwlDFU2Wiod3j4JdCy16pLQIyX7Uj3wJZUF6o41flx9UKTlvYh7bnqCktClz71v
wbTGhvCX2zuV9r6+dfrULT5WwgBtLFBcp3wDNebLmOuOQ9I48HmSL4MjmMHNdifa
bPHo4/pScSODJwL3UyyPDLHtqsWdGgPABGRroMSNuabtwI9s0aW6upWwRLDt/lv7
VM/K9ZIjXJ6eykVqf89qdgpgegWlNCshYZhkTvt01ObCfo8MP59gFQrzacKcNs/M
JVWtv1mQJx2ZlPV6jQMFzgxjoGKqdurJ8qe7OVeK3VyksFEFiGwhur7C8z5/6oyf
e4XqOcM6Cfmy2xDXPr9aCKCg5Qb3tVfqKiaPvh2IcHde6NjVAmsqR2Ebrgi4fOQt
ALZRZc9f2pv+nl0wTUu1DRLZ/D/p7b7YpzoJCmmjS8dgn9JpZ++RqvGVQs+EA1by
JLRGuB+9rlLNcgUGimUydfa/xVqHLnuFWTOJ+Xy7uxVzaYspss68lfo5H/wxqYHK
OhTHkYFWjO8Oi3vZ+Vv2z5S094lHjN1vwtcuDW/1C/KPJ/GCvFdt1g39u7qKK2VV
3SaWEQOdWHK6Xs7qtW6WRbC9iyWzOkQCGjZIEh11G6NeUESsta70x0k43zRosNcu
xJcunErXJ+2LpxUalhvmTvZtQafLLyB2+DJBFB7vzqannmf/qd4SHJENpuzn2Utj
Lr916TGkGM6yvsbRvak1LzuPPm1vspZjTUeOo20c55TEEplKl+niE8EMwR6VnCy1
la/8h1VK4FUYQX5q2Q58ZhwLtFieJQHu3uOcUY710P+1IoOnfEuMCSvp7Zbvf/kb
TTBvOfspTYBbGRANgGT8QOUnUo56fjdok03xFzd42acyDm5C1mPaCC5eLIQF1xk/
bqZVPkXcypcUXxOakQuuetxUpltoPuxTVF//J8CQ+Ln1PFZsEhF7hbDsGe+C40P1
BrIX9Mek8U1QcxzKSz+t7v/t/6apxSJ4EBAHxeyRkRwLpU3sWVeKWggwZhZYZSQn
Bqo3huMKoM6nFRYxnn0Jcnva+pYREvx97kqrrGPpPWPSw9/QDBiL/iGrcGNsmL8m
9mRjKQO4ywQak/TI4k95woHw0J0Rx32HEghWzgWbskvErJ01ssBH0opK4eiL7vZR
LI2trjg8elruaiNMPiLNZcRdHeV6E0T6ny3OkOnOowx8DP5IKM207cGs3sGu4Ypu
K/Ee6BXkh4tSFF25PUOoPm1ppdyatpfmeQMjflxkTa10+aDwo+uatNsfVNCkwmKf
MZkkILPZkQPxtDCYUSJoCz9txkyNe0PWx4myqct4lvOiuCUIMsrsByd9a3CIhg5K
rPyspR6cqKiudltLkA27cxsvJ+llODtDe0qbwtOAJ30Xh4uggcbYKxKRhrzgx7Ri
Fc9LIGyczIeV8gFkgH8IYrqrdsFFgxBksiTnbx1T/71pqPfV18OSxuxCFwUXN0jV
lsM1aPN3WQl1NiuPY6way0zURuMcaSBZvflwx6W8L9Qf4ZnVf951YwfyXgdkx4yK
M/j/kGSwtrayeUoHtFm4Z0DWBO7D8e8s2+YfraM1sjoLjSEeIZSrmW0E6ZX/OJSw
PASGSY+IgFQzJtNu6kEbEllg8GFqXgRhJgsrzsZaKlLh2Dv6PQ06vVTCtIvXTuKk
BdQskXLygBZQiw+CzMPc6Fr/B1vlkJSTBoZfjR30v2O7aX6PnfyCF9UI1niQKo0o
k9yxL43fHZ7enlvd/Al3vrg4pUMuAD9K9qdbgTSTVHW3V4IKzuqjXjcXra47FhKf
ixW0hkzKbe8RYvfQ8QdWwap/PRjTkrF2r+rr5jwGSSIYR/BEQXlPp5CP96wb1GBJ
KQqOq7hOziBHccohXRh/fONcWuDLYWnvIzL6CicXwFVz88EaVM5sCWpIcGQJmVzC
C6eUlhYqHwOjBmfVI8eu3wCHQBD/cuiY0d5Y083dddLvxoWU5jqOiHtJpXbWqjyn
BZd+y1+rtWDhIMxsJtnAsRTGnnr1fHud5Wcsw6mgQpyxJrR6px+T5beraAEpjy8r
99b4dRS2kddkAguC73NcMuY7SQXd/X4E974Ex1JN4HCRIxEknEBqjQALXhdgzmNp
AWtN35X+5ibXlIUI3CRSTJaIaQaKp8LBGYhEy+V1KJC6BnS4wYF5RuZx5F6H0/I6
pPESCJgMLCnpRiNYZ3DWGT4MS/5KLrIaVLd2oJO+LJvllly/M85W3z7/hQnQJzhs
9U3vaImqcTHoiGTVpvpqk22cOuyLzaAxVjbQunjOZSZE/W9S45bBIUlF9M0eJo5v
RTjsIaCystl2vJN22FVGb0mLtHiIhZwySLaJyPoMh2EofBpOqu2cX+MPSehGxwVB
2yT7IVOtqjfK/bEcjyOLUAjXb66fAnqzbehFLp4Zu6i/2jNlFtYyVxsJ58/JiUjk
l729cVg8Uvh6Azf5cFpssaygPndrqcr4NyhN927ltqvVMg15CeBwNuzvYOWwDdca
Swhu7cNM5pKlMaZS2XoDZYHeXkLp3jaJlN/txpwCPb3V8OHf+fmvthAZtZ/vpI/E
ZiXu+9mX41Weo82OVbnBaXaixQtnQOsv0PvxTwXdqG7lDMWLX4Cv1hSGEk2Svk3W
XYcpJj162L45JtQ9E8dsmsVhOstlJAjbT2XR3irlb3YO8z32StezsDh/VsFLTnvZ
36FIOPUqnDnO5btRrG1R21ScEWVEuuffmrMTIjXYJG7a6uNqsnbUMd1V9ak+LbDG
g7tVHD5SkP++VU3USygvcxVVAgEVC2eW0MyP1zF9rDJkBIqy1YjLzJ5eqz93dYT5
h9yNp9A349twRiASmevQd3H2I3Z1+NG9dj3ji2m/Bnnjb4oyPXAalDnm4GIBMQMI
0dYzrO5Z8qvgdaUo+3rK8tqrSV+De2lc+qBvtexlfcFxlTJJhm+e9IfSBDX6H5a1
ew0kdFcCh+NkhrugAt3OqVM3HUOAzFZq+HmQxT0Yd8K5AHguB23Bp8CGUYwaQjKN
E+tnCeUelvOulod0tHu1tyDuRUQHzsFR8R3KZ5XebWWc7XZGq9qdtUlT18oyQwFx
igi0ZbtFoaqhDR3TX59LZe79ZJBgPbnJfQlJ3JUwRUTC9SOrnDXrmD4Wf4udYQVc
TUZm1SH3dzd1OCII+8So4+L/BDEbPHuaFFSDpR2CTiMk+dkOjJOb8NCk0Oywd82R
ENadE91Jje1Gpg4TC+oI2TthNcLFbaKNJilCCtMfvYJBL50MJIK4IY6ZberX4Xuc
BKQvW1AgWoWSMdwjUSv7zq8tX0IBeZyGCpqpBuO/gWNCjpUhyoatNchBSjpB6Ubx
2mJFJ6c+5NyMvJ90nCr1vlKOLUGWUJjdoZknEiJm3S8hSEpfrMlAvcMB/LN8DTQ7
BucZV8X+s4dcD88IOVYvTKlJHhEcMsgaC8I9JaBg8C1oazhBjtfDJvrpTMjYLUb2
1kNaih9uf/Y330Zz30i4vK/tRDS+PsjGCdotl//a5egsAAYuumeuyNzYl8z6ht7j
IG2u8QQL/6+kzSkfW2Ca7aOovjzsbyCA+qCGcYvo4GiNP4IbqIK3tLRbqDtySOXF
vw7mbI4QB7r3Meb9nEQLrKADA1YcGLIfz6W1xna8bUcOd5diMouw/4GBDH6/fHic
VJMqXOy7ZM2lA3ddKbCMMuY6ZzgGdUVM9fayb9ZJzlQzwAw8y6mmA+nRHStA9r2d
+EiQb6DVtgqDo/E5c/46erLnRmus3XDw6yzZ4ZauHJBEUpsrE1A7i5uHwZ9UZh9s
ogcD+gK580JGtXrhER3+mv5yAD4yOMdMXxtLMuZeoLdc38AUgC4VGcRvE664RCJn
ASfAFaLN+PK7/ToXdehbqRbLDFjvcOCOkRmzXQIpZBsSNPLmEvjwCwq6DTGws1Hv
ICZBS2mXxpUkErhxsPFkv9+aOg9S+1ls81LHwiSAwre4z9mC8BPi7k0m5vecZYNj
SX6dGWBhqyw9dpAr/Im4bNrXuJ7fagQYuNTQr/e4etYwmLGaMjPDv/v+uI+5w3DE
tuwRzJFEETQxjyyZRHfwPOoGX9N0QDOUwsMiblTb+lufpfT9QgmIGHDs/9utohuj
Iaw2csiehX1jjK8txGvJLI0v0sWqRp4nCj6hQwTH4pbnK5sA9apqR41o8s+Hm0cj
OEWMPfjB4h87Yvd1a4g84fh30NOSC+2tHiB8wRUaa/YJVFdqzyEzEHR1rqRHWqeF
cyV0s5hcaq7c8UqBAQ7qtuC0ry7AZ03K9Grwr5hUbUyETxBd5dwfKnHgknMlV+nW
s92Ct489vJofkZ6QcbeE3Sxdj8sTcYvvvoNIWQEOMKv/zk/fHb+B5Yi42fIVM9kw
9pyB/ruZkLLU0D9hmRAe75F5Ek00XjWFkcC8SQ9rlAqF8S4LUaMGBc/ExjhSK5vB
DqIMxU+FwLMQKOMvFJc+EJK4a5A0UWKtCdPCiQ2CswaYXbXl3uwBnAAPJOdxkRKA
Vjp8wYiJhUNtzlLWxm31mbh1vQ/gudtF8o6HcEC6nUWrIPQKBQ+hi+hV/hvbclCL
sH/GdcGS3p8blW5xZ7LjNcL9jFGnCaMqiQIzSpLdW+6qzc0S5bArABnM+LBivixi
SscvO0Gjx8QMCP+oMLVVTkHwbFYr9coFcncH/rSFKe3aj3DAsqmHVc7sIBuo4TU8
a2JVLdaYgq6ubBRwKAwjeB2nop6UK7nTbavP7+ToPonUv54S2clZ4ojtuQ08dtiW
u2nbNxm+UQyTuduKvE2x7oD8KEl/Qhm+R91b4UwiyP/H/fMCGz5Jv3djD9xDsLVe
cRHs/vdrDwL0XAVzS2nWEfshwmz64qLz4MHaFPze1o7TQVi3KDUDK9O+roXb08Px
R2zNCwy3oP7gU9BNjC9nDr29tmp8dxfpFJlwLp3PtjYAtMYz1r1CuhJv2xwbVqiI
xywr3GL35pnkCXNY+CyHM8nrxCOSxOQ+QdVD4UG3HLIS4G4MoSbT9DweWsAmVqjR
5rmqUsV2pb1UfEAbWdJ6EoyTpMuVTn4VCqcTOZTtyw496Ck3TjkaXjA47EO5OQWp
g1bbLsRJDwdjPPgd4BPC+sy4xrtFNILwTXf2o0N7Tn+0poJx90snOAXvLsG8hqJt
Cv6nU+eYXVU6sxUT+XC0hdWWe4T09BgbYGSssKQBGPRoDS7KsxlocBlASSVs3rrY
ArA13ccgAZI/9l5VKC76l8NK50C2I2QlQsNTSy/gLgo2qPBn9JM/DCLkMOHtC4JX
WEwE0aYcxTF47W7GB8CEZutHpDnNIP28EQ3g6qqXzhMjPJAFJLpf7l/ogXIv/C4t
Cz7G9bRk7bH9g9F0gS8gHINMbPYc4m9gbcuoDnsBX8BjNnwcmU6uSXUfy6rAlsSw
/auGvoP6VhtxyZqylSPMyRi2+L9YOQHU980mHgVLLaxy4lEIqHtqiuWxSrvOOGEI
41IB+BstujiiYz6YzGqMAYiWx+AfZwQ9DABoz057TngtSUMwSlqBRwQ1z3q5klFt
RRwkqZ+nAypb8kPpG0/PgCqjn6SRMEZctvR4J2Yj+uCY0EZaCB02KtrTykKiiwAF
gTACBJvLYkIzfUQYwEIzyY9WkiYN/NieLcQFxCFTxhlkBOELdq3ZuAmK4AO7H7Bx
vTXTbavgtlDmXRALlko9LEU4XkbljquHticjARKJkiDucnDQZvLUgPLMW46tunmP
gJC/a/8Zo1lUL8p53NdVkGuAusG7uS3Zps7vKipAYgaN9U5qAHivo8/Zd6Vow+Di
QFWIdtQJ9cFtil7vonZFnU+TLoa73Y1YEkCoS/OCke7Z7SrjQwpymCi8fKOKEVmo
B2Yv/G3GJm/IPehzBEWK485+UhMm+ipqW+iL2PflJdrlDQmg7xtbVUWuf0O3mIft
1HbSAXEGbxMte/ogHu/6lQfWf5z4VGERtVBfbqM6/ri8lYb9FYa0n8CUlMrr5kVa
5OM9JqlrmO6OxtHG1VvHAh8Hpi6G6VANxse5xbmbSyTqszPV6thtX/XVRzVxf216
UrCMAMskAlsvwHYACZUAkw1qE4ZwlCrKMRFk1ruoS/whxH1Q/jlay1Pdl9s8NQ+3
s/QqBXwkjizSmFxoyPgvqgN635yyFD92DqpidWVMeJGHwCO5dAVP/PkkxiidWXea
QT+hAGgxWvd1casRHzxil6WkL0I8ol62DkgvO1DUBrnh3/fkPcAShyum4DgVX+sv
q372YQlYj82l5UeprqznkKECnCdHisxLcaA5IP6zm5KTFTbS4E9fLXsTRao6c/EN
jfe86l8xx1o1cRtfaHM5ST8L1wXJuD1yoA2VZ08etfy0grRDbMMIqtCkQVLTInn8
6o+xJ84/k7xqFb4FOWPCwJGYwTdZ7NXkYt0p/oS/y4rwz8u2kezYtEYusTSLOD9w
FIgedKyLqQy/MpPSb/j44Qamth3Mqhr2Md/sTtyNyjtr/5l5WY7NZpd9/dHcQr6t
Fx7xF5wayRgw4djeArGod0F3y7r82dR3T+ff+NHFk7FePDDjewGawgpuj4xfYzFH
scpzzSy7tcTx45YKypogsiQCuJnC/KiwcmHCRAHyjYdNGc3JCFL7pbz93ffjFjua
XPMJYHudYkjJPtb1MatojC3fQM2FenTZ/Tr4yqi35VhFJWdNHqWP5AeknjYnXCDd
ms9MQ7zUKdLj8JadV8xOze61bAFeaDI0yyVPi/rHeRqPnBgJIYhb837C3evqFQRA
BA7c00LiIS8fFOr7K90B2S1b47PH+4KI6/WBpd7r2LoVwl1iYCkGlugtSZSxzsX1
wC6FmC/uaLJH3XQQ2dCgd+gamFHISOTL9R3sU/mynTerU/IxkiRyytBGyZf3odS0
hznxxbosFalhUZtyQaRrd5JSApkKuZhVITSLueXA1BpkmGAl4KDHOIZoa5YljdW0
8Nki8MKBsuRxPbi/ARgJ9XT+cCFujRWqHVXrHNUBjWKAVqZwz5fHZi4LbcptQsaP
VUwE2EYrp8Obp/kpmz1/TjLqq4b4fEvLIleqEMAXuqTSOU4F4uUlg7CmNCcci0El
e3/UyZ9y2zA0zo6aOvvYrvRz0AoFLcFlLMRv60cjVqIuzECeDpeJIloFF2wdUDYl
RX9IRdpmlI2OkCLVrvibscZisXrGdjKEpSy7iN9OjkS1CiMw4ERSWteGcNMbrt5T
031SpW7SmH5yQN78EqU8vJ4k0in0c512QkKFnwPJkfCUu8KcsEmH5Tf9ibYBUjsv
LcYvSviDu2f/irPbYrW41GeSR5Oayzd7+BqImVDGUZ7Kc96jvkkbsv8Czks157e8
E4AhCST2AErzkL0KQ3W2fZPf6sdAVMkG920ZFqM1H8ABq+IxLBwF7mFplDRDZxLK
EvjAHeB/+WAoB53cJ0b5FYd4MB2zfoCTYnOCS9KdHisn1+vGXm90rptbjAMM9rh1
fBEulmaNifUXbqnv19Oj8Jvvw/dEjVTMrpfFX/wkiTQlz2fLKuhH21Oz4Fgv49Uz
yCtGbvVZ2EBMsFmvLhTBMHhwMS0PqzWCer880zDiqAAXVHiD+EbQha7VzoZUaHM3
mblCfGhgmHfzOIj1AIc3s3fke7hH+OHd4h9+UdEwxt1L6/6N0XRXzzySZ3MAestY
CfGuQ765HyJzYPkef35NOR4mw6DrlBq9NW5fwmuiJ/pvSjaX0aOv0YCatBF85JVA
8TNNkctxP16BuYvK8aDLPgC8bsleaBZuvgvZq/W0eqO7LA6ueqc13xunZSVvl3Ue
XjegLRCERyWRXEDOgsWH+PoDLlsIbBESQ9Y7gBUJ5UbpT5+wt3fiU9wrfEduOODF
kTkmvgkdiNiWNhkBRjZN7xugsqeMd1JfNL56vfZPbI5cJxUrz0JuWNvEJWurkEve
+/eygPfYjEWUtlKyJZhGVVk5ccRRDnKPZHOdqneC76hFr1bChAtT6CkhK37u1Xwj
Zh8/iMTrBuyvAmHGx8vPZqbzv2NPcRmxndSYv0cWU86gG/wzKMSjfthEOxUoCtqA
RumGgeMuihZ+16kM0HpooIRbLo77KnQXhHQxpUr7rcBKMNoBfMzsBJnrVOCjOf5M
jvMJgUdOAJpFlhbnI2b7u4/9Z9+D7CwNIpRYEjv+wJyMtMn3j/CCGrovxXR6ztA1
GlMd4iy8jqGjetDm+vKgLlb72PTFrpu7/Azx1eyarDacQxzptouP0tBq3TyX9s3a
l5WRrZ7LtwTz9jIF16RrvONeobkoqB6j3HhwF8p/eh1aL7m3V6qczEXm55KcdDbK
c7WCAtOt998ykWKlpAhNyA0Bz/Fkcr+X8NveKURqmB33kagnCBRm8wyM3zzMaxHG
3yYXUIWzBrHnOJb4TJr/HCKgMLLTn+2O3wBWLk0rPSgzbFZjz6EdOLLVWJWSQdTG
1AobNQZhv/r5nrRvLkkQ5PyVBP59Orp9vNpcM9YpfxMvDwaipa+Qhom2vaeb7Y3Z
3PxX3F32AiatP0jQ5UeQR4JoVkrYE/HgEET3cMrN/UHqskVRBozRvIoABoD90IJb
b3M58ufXrSaF/x4XY1epgdbtyZDBcwW1sP1/xTCLt1s8MVvY89HWQDCt3kuQ4i72
pCWZCYicqOGDL3zTcu3thKkYzJYZ0t9SWpk+etzv5BvNMsNQzR5HXjslTGc8Udz8
qRTp9hoOhagmfylqjR80wFSAE6P9O8/hJpXZIIODoTUavf+HJC+s5694h8wAG94l
4yXQetJ+jz79LbpxlC9Dr9Nu+6ppN3HnjcJk6hixKa0KPpLO8GPm7Rcn1ofoAj8k
IdbhBCz8dTNJKoly0Zw1FKdLbqosodimwdYxMkOlVYIujIm4+LSMi8JVlyVViKK1
wnlQmzWxx+nf+G7+t4txni6rmGys7/pf5GVdCtkUDK1uwuLm9RByPkwD+Y4r+uDW
S4c+DxvbLUM5oEM21vrIBxN8o28U4SI+VhvuReF/Lm63S9zkT0lhSCr/venXejzl
dFjcGZzJ4Ooq5HtWrGjhJhiFt4iRRJegTLuzgh0+EHFUBaWLOoBFDz32kXZSy/9B
ev4jokDAJWiIsv+5/eBJMvMANTljowe0IqvY9w2JlkTl8D/AY5zC87IHjnGhdPtP
Spmdm+gpz6AFH1vTPf0qRCMjkORz7X7478bW0iTv1CKFG7lHEhI6cnlzLZluBqXc
+kZcSr8a4GWySRV/Dey/TW+QJLOAsLyLPHxmYvDts4PfvQqgQk4xxoBCh342kD2E
s2BdK897bx+mcNNjbgj6rlqnJg1+6lffPAg4SI7yGG7rajV5WKAsWTvBYj8KGQew
3+scIEl/ko4RKZu5+gN/4SVo4nJWfK2ytJqP2GryGoK8IKW2Z/AkbTNozR8Gs5+m
vMTlkl6btthhrCLQlsKqZ5lzOYcp0Q0FF2ofQdICwJE63Fmjvn1CxCxOXNsttsbr
QNbP66ts5n+CscoR8nsv5r/WfuEK/XY13CTVkkJmWvw5QH3VHHBnrdYfAFgn8vjU
FNZ1jv3Q89kIIUrlVo4eNR3KsBCEosw1aHv+SZxvdF7iMz8/r41slz86IsOxI0YV
ojxLUSQtvV53I3YjIOeIi2sghQ5CKFa174Y81wTFmAfzaYdNg1RbKFpTr1YndqTG
S2FMmkMOCh+UgXSFZ+KxS3WONlxMTJkSM1ZZ9UCbvJINRDggVMDOF/TvtqYKGTLb
RmAVb1ZaKxnewqBmdT0JlGVbbxRp4klIcXLPq6EiaedfpkOhcsY08TcLvktKOKyi
rYJcSaF16bB0VCn/97hK/GidTha6d0CT80G3bf2TpXm+c1B2wsfXfYB5yyOVv5tz
DD1QZlBOWamtPjTokz2sRGsufIE+W0y5DHpQHHX7mt5ZNV4TA6VxAxI2TAicTLbA
XHgkZQW6QC87Q0DgdBGCh/EqTdvq9HjPNFOrRof7xoM5awBzju2u0FiZJ1PwA0gA
uzTNL1lRqz6s4CMpsvj/1XML558gt3DTaEJkUHbJ9IjfNpwRGQNPO9MvExEm1wBr
ecCi1KAHcFob39mk7ZU6tqTKNjsDlUAIQFRmCvexrILrBaVDCygkM8XiZZw9hxxm
ZMSUgfdy6Bz9cMT+/U27RowgxdMfAEBrqZgauSByUmDkNtt8Gmve72/A+MNg6iyV
Z8TNTt51qYc6ywMbu7oLvY9blGASuvGa+hHJZvIoM3bRG6mWOXvA54RU/bX2c3ty
+rCLtGd0rjR79sBjnlMe06yFHrjZ5Qb2wncsfeDz7104i3YvSIjAy+KZY95iqGrA
k5yFintY8dsJiOz3TNwQKaxSY9ffxOiESUaRscptI++/PViE/fbXr7aFDPy2Av8w
+dS7g3YfHSgB4/x+P5rWdUjir4s9FTXQJZcl2I0zdOhp34TnBzI1/Lf+Z3Pow4A7
2t1KvGG2tIiWMFwKfmmXLuyDJOV1vyANP4iwKgzuEdqM0dT9V4olLXZod4PVUt3t
JSAfe4OcltWOo9zpcrWLaUsSwwQ+jbrkWmG3Yw804maqHMna1cZMK1ngqgRFswTe
oIAevacAS8B3cv/G3613aeQVfs0ighkUyYeXXozm9+/IdN5VguzJjCqyrU+k+4dX
43hb9mYWSCojLTHxS/2PiSkAhMvQXLP9cTekIP7gdtzeTU1vXR13BM1JA0DH8Sk3
2QI/8u7g1Lg2dP6sSOls1jq+f33k131Js2GXK/lEup9WiIFen6c6hh/MFin0i6N3
WgPJ3YCUYTTkz9K0NdS8RuueKCZB9qo9tGgd0U1xpIbls4gew3+NdQV84FYPWEGo
KQ80CgYbtMkgVjpRHGUEJURN0aIDd81BWWtuwo6PZxfpu2CXgj6EGEj+WMZFmRml
uUivSLpUeJNVq5ZZmG3aCoCQFFRwjoc0+doTk2ukd61JBt9s2od5ZFUGkvsX5Fgv
tN+2yiGTfwySd3Iz1BbmKkTMUY9S4YlUyLmLzI/gJJAKh/1kqIVm9VCsjj2t1381
7mai6sPQzaDH46myz/hpWdSiRmMIUZwskSj44aR/FyycflLm6MrmOtKhji6LPY+l
M5BQTDJZP5ZayLPeec1wBd05ryp66jlNzCMd+jypOvULav+5s6i5ltoViuf6g/6o
r+hCMla0+c4qrZvpBOI0sk/1N9zToQRcve0fvMn2AMt3ss1aOaiUQfQDCDvX8YVV
B/Akx2p/EroMZMR4yCyca135mfekm/RCSCAT9510L97qC6HAPg7a8xx1RuGXSHnj
wmeHknIZ001Y8XKzjq4MFB5HpoEIM6bTsZRYQ02Fsgdv+7qiszKNEjKwa9HDGygx
Tp0P1bqS2g4E8dH9Df7d2nVtODUb8173O23ZfJdAwl2UdQ1wP7Vn7fgHmx2JKLyv
d2qwZgDgceEXw07zCFNNHwFKbXnLqnYOtINvX5hMSKmwRNoVNPEItO466zP7/C/g
fFecYSuf2GQrgUUiZ8lOq9DqshcPUDf76f6/Q/6fr8DpVossacjSHy4VkluGPnmO
gwV6RZHpOOLRKOqe1sqmOFUfNJo0Uf7hJGCco2Lkcwr+UESxtj+VedByzpN5EWdR
9+WxqEO8cCJh3vEnxfcGgwMva133r0Szr5pEK18+P6JCVGsHkVWaokeB8sC7qpbq
OhbzjaZUxLdvyP3UI2VaCjTqzmosQpNReFIZfbLyjrZ0XkYpa2SbYqVkTB+8lvDb
UGxRMIk50ThYeR68x/YiJHBsQx1InEdtzo+gt7u9a2UUiBV6suqTwcfY0vWf4uWW
VUvvGI4/rNFsxw9e273O93R2vT/EeOQ5t04tgGpq7BTjg7c8QEs2/rCYNgRAD5G/
AhZlF00vlVYmehn2n5p/WSpSfWcZcgDb3/ajk7fTStiQpRQ7hysPb4bKrhd5OMFm
Ynq2jmDlAjuAsuJdlgYz+SFroMhxwa7jQSkiTZsIPATKgmddTJpoEdk1L6nAkPqz
Keq5aiOUHQrSpnxk6hRpR0VAmHbOf2xBSIJ+PJDOqnIUE5wYNv5l+7reYbYjl8FY
lyEYnS3y1wriTKLM5yjbRWRNYyRRcihzs3zBXg8UarAOkCAtMmw4Oql9q6BIv/O+
QJWSPGHHADezLe6sDOEsdQSmMG0lBjlN5bE4TqJ0B8QaGrvka0i1M/M5WqtShWmI
qsY09uJ1mMLa6z4ellf0KIiiXFn0obp1H3N+SfrKLYoTX6tHptoCp/hariwBn8xM
WN1y57pL0HQ84GvBfb/i+j+fyQaDFmT5rxRA8w/4h1ilnFWiPyOlAHxwenEKsNnw
Y7EZAcJCJITAGDohM4mCnVt1HKutY8xjPA9dwLxNoBraMvu9DQvorgdv50+7Nb4V
7a14lsAPYg8e2AIgnGHoYiHgc4rC+txtYlfw417QGfAl4YgUK5ihGLDh6pYEhx58
3tr1x3YeJZmjfwfamjaVGRkCiG7ygK5uoqZRfdIkOsyZoHPlpnHxMwWsQiReMWKt
3xoNsrDNUZAyYluD3hByr/+uLbKoFxQhiC98igAdSjKbLrJkdHl+2xHAxCWwRYOr
tT6dhaJuw7JNjTptBgNdT9AC9SI1PYzBhvyBByQ0CcPtgUhHtkx50C4GUTRvjYZF
AR7rvpGA+DVQ0UntD1CzXZyyTugWyiKgt9HGlscq2hU4Y96YQV1mEpopGoYQSDx6
7XuqZA7Y4qhdaR+aWW8gEfoTdN662eaCZVp91YMJg6CLGLuuQei+9tLIKqDKIav4
F1lQ1siKRlQhBgREfub75ErsNk1fGbh0zN8LxG8VCEZSAOteFWNjMBB5qkEKVj1W
/Jwn3U5yAW2GhWBc/7YzGGEffzQZc0f7J1ooXf5E10CKhnX8mJ55CE7KkYvdNoye
EE3RwSXHevsflw/E3t2xtu9g//3RQfoPFpahgX4YXxqq9tojaQl2/PCJnZcKRw2F
Ve7YUf1GTI8bL0+CdeiVTleGTtcScNVPhzEtNpMi3/ed5JS3TxUW1PXtu34kJXf1
mtuRINjbxTz3YthKIZSy1WoWn35LKKilLUe9KQ9lDZ4peGQP+P4nvKBAlJ8g268q
Yncb8n+1auHEgCCQcwFc6YQDbvLd5sk1elhS/kCzSNZFUfC1JO3MLHQf/DwbSBtb
HnPit34JkcS5pUad13kAVHjsWIhAAWFMW+ChM/z/mXLKKAAWwx1RVJAKaQ1ux9Gq
ky8vcfNYnCdrVDPfl3M5AsFEKZ1QJSH2JAvZ4e8WDsyfIEcPDbi2jqDSiietligr
n7HN60xh87Ug28H+FTX5XvKpcB7PDlWUs2kAuUB+0zHvxQruykSoMVnRTsPtqnn1
sQI/aHhA8N3oGA6zIMpKWIvnZ/F6JiFt4cShjRzx8YisEtnt64nXVRdHpWCWmjHW
ef0y/OOWFGB8/peI6vtOOr9r4dQIAR/NhHQE9I+VnE0Pbgk8mJRM9yNJxnU1OH7T
4jpAegxcYCD2HGHnsNLPh0fnYSlzH8r7lnFbwpWFW1yLYp71Sxz2NNDeGAVHGcdF
Qx59Rq9UkxMHLtqCOAXz9675DBg7f7iOE1NcnlUF3Z142jTgcwyC62sJZAPXyAj4
kQVhIXiTw/ImJ/AjsbvDkx2ZCTl39voxyCs+36ehz2pkhqaislFp8BtjOlAXFhMU
rkEEtigcsMUL3AV2InWMHJl9gCP4NvO1K2SHHFibmf6OXISetbed21DUI2LIUTbz
Iur97B8EZKtc5Gob6Oo5139UL5L2VHiUsN1G2UhkWpqRNg0oVswwXLM4MujBrgHE
AvuZlt71P+LcCv3N71YJEBwTLV76fG0HW7nHbon0NQTtSSJ5V2aT7dqbGonugu4r
R6i3O8b5DDCtjQZNdlwATp+3NGosG908GTN69KsKMuDdJwFvlp5dahnactVD0Sab
itwSzhjNTJb1xlPF/Im0HtwTKm8cZawzyn1HbMcVFJKIoV+vg/NS6eGq1slkRsBe
iNznjgkSKO6n/pGpbQnJZi0SOMz3P9tHg51JHs+/zBYiPO04oGj6bHCUTWz21MhC
awwX7vJ0DSYNGc0SbO9r6Segs/A2wrbDLEk5a8/64Ks4UeWSaSvqxx4sz298UhHp
EbM0HFxBCPnCvYxKG8Euoe8RqUXyPSrbkb+TgdRGpAca3HDgusj8liIrnmct2jpa
HSO8O3+hCZ8FgnvK5Pvqw8/tcb5yqHH94hqwnZ7HWZ9iLEJfY136tjm0DpZbcRYr
lavMwy6lcDTeCX9kR/MJVAv43vv8PkS55Twl6AfRJ3zPGwuyECNgxbnLr+/W89hC
S3OMyLvrmRgZksQP3Boc5jB4TDgYxGDaKlpi9LxVZT2z5HZulyFwZwayLLLfZ2tL
kJtCsYve42XNN+7W8iivKIh+HK70wgOk4XfndsjCXxkQB31BS8KwL6MQa+xpV12R
DYBdAjzwMW0QFh1/4b5H1r/TwJ3b5zJqxDjKzPmhtiKSVe+DsTil8S3gr+WMqxw9
BmMZ3Iq/VJy1WLvHKIHYdyv7/AVnS2Lrs1Uj53AJ3Js6uyJF5kysizjB36XP5Hbl
D85QGqPQjTVXMD6R9H0ZC9vT8FeCjv97YbbjzvII/mnUbv+u4QYKjCveci8hBVUy
FCasU4kgvXHHuSsagXNrU2tRlMHl1uMJywV6aRZlN0BKJw4T/73b+Fl2zbBsHteX
NMopaMKHqajepDlps5w3hBuLZRRng07CTSii6dNC+WJohP0Bd9Vg7mh85fE6Nvtn
RBw8uU6tm/j7Uqkg2Jh7kcHiWdGWk7eHposzRvVxZHlJYFnAUXDyejRs26JGy63X
Qlq7NehcVy6HhMMZExrMVFd2TFTzqfc4KnOghfzEC8RfeHwTAAbw36xxrrgTo51i
gbM0kcflCtMtAC5bE0tazIAlD4ihCO6j7+ddzRMyZr39736B0E6XocsNtRRvzSEP
VZRetDu6QQOM7zJJfXOSIhv5eBEf9j2nr13IWmiscDWle93ByFHu4urJKmuO1+ap
uy1QnCDfPU+bLv7OBOQUgxssJnabGjUR6lTFkb/G9Ku8BtKbyJsap14qnuUoME9Q
hhsONzhnr+C3q3nwikKdpvryVS8X/KOZFYPx9hUj6pwBYDYZiNK8No9GBxHbOnbx
u+NLYnWRk3R7PG16l/unVBiLvtk1+LaUlLXarixjjpPWj9UsIErrHk5jPrXfRd4w
6HeQ+6ieLXrk/yHgVrpgDXrmpdunvVuhTwrBNnj5RfGopv0yw0Cz1S9XX82/XtwC
kT/ALtwKaN29dQjMms6j9YPVGQyYo5EgDaGM23yk9wetKvoBx5JOQYO7kegNADIJ
qU7rKHKe+Qbpvt2o+U5fYLjS7Zuz+rr8Gv1MGOpdrhPWA+J9HTJyYmi73U0YxUiy
KgMRKOnmHIQIhcIGb3Kj38z9I0CQZY7L/kac01916RG5w4VHrPNN/GtVJjzBveQF
TZleGWPlUe2m7Kt7S2jw1cOVgnyZNrJ7EruJvms0rNJGKoG6aI4NpVfuGA8LocVp
iBCzeKJF5FZsjtaTw1balZIAams+BO3V3TelMT6eqB0dPNS1Zv1d/a7R8kxoHLZ0
NxPaxtygeIfLUfEySDsJklhbosf1+7FU3YtHJT/zcpoz9Uk7ar13Mq9Y5d2B5zrl
UWJ/BqRTVUPK3Sq2FelIQdh7u1VpVcJ0cgQHVVBMiOkdZyADK7EICRdeLzKwRp7/
B2Igzxqdk3wdyrJt3mKpKIS5f3az2iHLhKX5K0q5y5p2uw9fgVczE2m+USdG6zZW
qRO/7bl5wJsksBSSr6Fzkfp2DEWCPIGL6gKTZXokNMPNmHo6Y0VRcohvENRxndZI
aDpzCD2lSq6JOzo5Fhhh96auqKYQuQs1QeQVqrP5ylbCHwwlFCvVwzqjKbhLZkz3
ZtEK2ZyyX9OizZ2O1V3f24rhwjb2UUrQSPTc/WjC6HmoJP7HvShzryDCfeCsgDxL
KhGTEPPRyYuH7Ei6FGx2GfxUeYvfLoHDFottr52n733QqN18y3230IFErcxJsG5t
vo0GImSeo5S9dwoIs/lQW+PfVkZjAAbGUyyende4O9Bndxw+iipxgU6yAOtmSYCM
dQaQlkwm61NyMrdgAoU7dwD7UUnwwVMT/wnC9+1LGKwUbP8YF5by3mvvw0knTU6n
zYQkwSXc8sdd8UQTdw6EjbJtb1rXVU/J9WrAqMs6onPApXgcjkywhzOS9WWm/tPk
ED40cvstxorpDEiAXa6l1crdTi5FeLMVVn5jUjBljeT8Nj9T0TkvBMvxzgO9LHeI
yS5VLNcnt6lCuk2X/BKsMegZhGDbOK4slgmjzOawdrbr82zYR6S+BRTa74JDXyAS
L96Xas+gx6mHtK16BGoUci0qNp7URzBluagYsIPSxwTdxHnjYyZBTh+XhWcfutdI
AYAY1USihW1Skjc5XS6ZP7YcxD0wAMPRR0XNG6mu8lWLkRsh3/UJ/3s82tEQ1pi1
YQJr76pUTHByqnc2sEHVONhBoxEUw3qFFTimnZ1+LhC4k8dJbrppoDWNL2Mbusbv
vhF61P3zdZG2QTTqzEisUrWm9GI9AB5oEhy/LiHfuxfUGku8tYIAO9fEkdupSwfs
Z6WmFze01OP0nW23pf46D1GqkDw9/dBPXGp3Cyzp+DO7kSRa385aU+Ot4jbJEmnN
CshJ03IpUCokfQ1iWYsFdye4QW8Si/LSEXTC+NDEhUvcMkHmPQpe0bNmJmUJIXGj
tOqBdKd67VMxwe79sqyTqlhvtVJ4YySdDbO0pPse9P0mu+doUd6jvwmXqqhWr0QC
xa0FTQXrMVCcUpTLam3Jf4kY7m8iJ/5h8KRkEYyiASMG7/FJssk5OjeHf9+ml1+f
kJfUJQQ/dQD0dLZ3Nb7k9IIC2UtI/t1hiTG70oOuZmp2CLjnhfMleGrXSvxHs7Ju
Fg1oScOLNgozoenzMXrOe3n/lfHtLedGxBZ7ApAaofzZaWTLisQESC0xxKl9OzcD
KbIdOrWwLBSLc6rIzkLB+WiybDr+n2NhiNV0UXg05+HfpXpTxu6C4TCMOuq/j95G
0/3uwaLpAgUCzZ33MWp3L8K95fPG5t09Zs5rqU/6FjBRoRB+YT35DOtJYPzHFVpp
tmai9NGqgW9488f8Lal1pQMwfRIP1OBOR3RERl+kIqk9FzdfdrDGKBK1P6fMEV9f
YaWIqVtC0cSbgmC4VfeoR6G89REQS8IRPK5e5WPN9KCq757qyC8hjTX5DHED0wjF
ik9kRCx+/O7niVI1fP4kTeJ4Jg+MlXFezM67fcfW8Z9UV6bXhbkT1M6qyqaThQSE
zgc2GOXZNu/KS8jAywJj2v/6p241IbovjxNxUWCK9I+sEemzG3O4+t41HDvCugjI
Zy+o2FpgadxuyP1US4Mr6D+aCDSIwbXqHrR4XN6XZ0J7kdzTZ0Bmd+OAVXuA+RkG
QdDy/7P6yIu5DUc1o38Mo+weQThCzOiqouielDt9S3owdazPAWCOisCxPavyoA8b
6HWMP1cWAxHmlbmKNiUKmxGVBjDVOZhb6gPVd5bGcyxGh0NijtoHhr8TojgxlLnM
PQt5gUemP8I/7qzrnZ6r3NC0eAWNSjQio9Qchu8Z4pnKFXwQRTs2LJPDAFqx/KM9
gg5/NzfpK/4xMevPMa0qyBRyAbWINqZpSY4xhKV5upCpHLRL9ju4B5zV/Ty544h+
V3jqq/6V2CBqEf3bRdLI6qKO08GKBYmllx4rVF8K6a2nhrfaij4qxaIU9zf5WtiE
8LmtK0/jqGAnD5SrKB9SUIp9CJMxPsjIBp2Y0LTWQMI7PNwOgRFbq6UDa6sI9wd8
GPgpoCxNTzOo2RGBhiCEIIb+rarnPiCOdebNceELSZ2LA/GC0YKavipdyDujio6z
ePRiy3x2l4QZRD3Sz1YQvCqiFErnBh2BXiCT05RCNQs+KR+jFH4xQ2CvJuXgIAzz
XOruBk8dit1xkXNVcA8JcjoB6k8G9iMEie4YOIwkJhSppIpCKp0JzzQqTI6BVy0+
861FkeNBAfLGaVQJMi5FVRnK2iMOspKG7uW3Xi54glFKIkWmbXvu2F8kSs9MLCxq
VbBcE7if+B4p3c0+tb/ea93iPu8PedQMKx626L7mhiYStLVtwQ9BVepR4wYtU3qq
dsPjFmFqP82+byTdxgQruubtClnqxoUQTnKoZ2yd4hD4qmlmxjJsjqtyy2KQnyY9
PZczcIgF/kE6oPs3iO1ofINebVQnjOB+Ffe27/3iycCZhXiqrkJf6dHM1PystkRb
hcEpskFl7Ye6Cy42fTUsA7cxCNtAAr74NtWIvizgWqeojp0C1D+YNE5EWDiRtAPY
GHDNjXzpkEScUYiSH4iDNDKzdvn6MvvxPeQLa4uli3JJPY03u8GOzc4nUkF6mRNF
J5SMegSdU1NGGlZ2DTzzX0W8r6G8YwrOckH8hJKCmNfPcj6eTf/kRIUd/PLGdTfb
hwPWiIrFj7b4rFzuvsiyA++jXVWDm535LjlmBSxeOT8WKNCus0H5NQXei44UTWnh
FMtHY0lsRW11ZSIJbxnsF39t/RDuK1fVwTj+ueh8XbdmaRFFqSkehgcrJeiwb7Ur
iIq4kGiJyfA2ofcrJ328B1fIah4Eh6+QATNflDMxnaqmSB5LJ6cMcd6ba6r9tQyM
S1FINNoYcDDFwzOx1eaoJQJ51wsG5dm4Q127fIkgmilJjiAbANFl4TFD8TGXvNrL
/FBOC7UO2glWv4m48BRG9jCVrNp4xjlULJMJZup70BpmROMAju3ZY8J63jfdA6Er
J9nLli/hE50WU0Fq/JFlLJuxrRZmbCQb5Tjyrco6bNn+va6+qnuL91e5EJbRe2LR
mintdDmvj27a5k5FmHuMWt1J2L88+c1A4MUpic9Eo8PqtCBbqe1ul9xY9WpSIJqo
WY9MhXX0BOCkskRLbwVuPL8n4P5i0Sx36Yi1H5JSwEP7JyDwZJXTloGpsXPbMOgC
8iB9LIant64CGh9tkgDZyAkrq9Tv3VTecp+xR0Kri1aOGq7BZMQ8Uziv8X40ACJg
b3s+gBQQjzUsoJ5w4+QIp3UjD6XFI2EUZN6Htnmi5GpsCVRnCkYkjCwZLH2spXLs
teEDR64poaZYRqGJ5xQeRTZHt4IVKdcJh6uAxMLn+McQaYOPFxk5RROX3FVy2RWy
bAWNVN+jL5jh7aOdpzZ+GrO2n6XcQ7yDkP8cDznljD6EFTDozGYQP2FUopSHahSw
dKDzLJ5XvcTy8UtnlRNSQhFcxCP3K+O3+JzVbPMos+C/hDi3RRe94eFyYwh5G9Qk
wWMAIxsU1d0OQ4QiAZ4wG+jgL28ljrV8P1DlHKoBhDENJW4F+00KQkply3PGFJ7t
O5hRzYA0hLuIWvO1bBB5sSDU2IoMTlVnCzeNngYIUCMb3JrXOcwHSTG9r9CaQZpZ
mfvOyki/T5S5lEUTIOXo5GEIspoRTmFxUBbNVUkQzEkB1LOTZJFLKqOPDio9H39O
KoA7+CsNtdrU5EG0jyeehhU6AWBTWK3psqrxYxz7lBw4o5/K0zeQ7i4TP0cpJp1D
FHkHPIi54eUJ0hChIfvouRCDUy+9hdNQCvD6M34Ys6TcckLbkyYw58mizeTzLihR
qwNLoF9frPPfqXMxPVSbOzw+6qnbYfRcJG/5ni+6Gq5xpt3YDJ3MUFJzBO/iBEpR
izxpxFr8Nfvk6Eeg+VS8TccZCOM0e5VkABcTSkH7wKindPO2ZPZZU3d4jpSUwGOF
7MBJTiwJmxpAn10BvSW4RqD6+tMcAiObEwMmeSV32X7kzjodz4nOGzR08Jn64sUG
QwEo/eqxUOhqDE9b50uSMNwpN6UBezMgSwbIIFEP3qoGMpSFkJqkf9+yXpAK9iKu
RTekpHckLuxRiOdc9ckiTIn7KsGAfMEywuBu/OkGlm1EJyiXN2g69Doy2yeMh0r7
aFCtj2o6LFzKhYOVb4TSX6aRaNhSc6cSu0CYQ13elnLMw5o4eigi0qsPkyk2t43S
GI4Q5PsoE5fTtRl/iYn1gXzNdt9ObjBhNruvx8A7yn7fRCDE8ki4p3AAb9bbonZ/
PsAIFBpmUkDc2Wu1rzp88RGu3h/xkFudSzg2dKdSAVtv7dhi3nIAydLi2ue0L9v+
BV3aC1M5kR1gM0yz9hFtzcc6FStbIROVGXl3YObzPPNgF4Xjx+7mwFzrx4C7xI+l
qJFC0VLtAewmbxpBzpR77dUOlvndgV3gv+7f50NsgcwLbWAHtSD+3/V9JMlFwqz+
OJMi2NxDOxwrFXyCK28mXo78kcnnsxIWwF7Y6rOYmWXX9h+oZI7ZzosOKP7r2Xm3
kt47YOr5Tp2hBAgtQPtM1yYZWXIipMKOjqm4iIZjkDehH6YeMsq88Q58LDLFbJT5
RBq0O8TIBix8J0s7WkPFuELe5iGIZKlnjsX63emw1vz7wErSo+qwzoKzSQBG2tj9
X8ASZ5fJyyYVfSpohkF1OKkFm7INyok8lAjJwpJOhVPV2kyDMKjOvu02lfHBIGT3
qPypGHfO+akYtprVdHzlTtQIfpJdjZqME4+gni7LMz+Gb/Bw5ldLA7MZC1Vn8rQV
FhggdNQfO4VA+tcephPTBvdTQs39GX9WLKgxRdig1ZvyclCF/Uu3IfiKQaR93njz
/HBoOGYUBjNYC18+TcJFX7qP3kWUESlll7zaOWzPT/9aVRSFJvOuolrUtJc5rSoF
8mIaetMASuBDWy9VkQpLbXHgkBsyGrAii1EpiGYvTBVgB4WwjG0tvCEvJcbNWf64
2aaCIvqox/AgrDKMCanLS8wkT3GphIVIFzPKhXHr0q54V58uKNAgNgW3A5j78x6V
IqsvbPbdmgBnPz0ysEKC0jB4KFR430rZedIR0KIVccQ6nazjRjUDGlg5UXJJfESD
VXVKva9a8HEFd1UqWieJT9GPpIZh6r+j5u6SloF9BVxuLxFrvpAONgiLapRy1gPo
4Y7cBvnTt+mNIczSOeMKtkOrCB2jbzjX0DCq9bfAJu2G+GRmXcS4ii2MRucctdqy
B8UhNsjCkrHbU7DAy7bUYGJegdIklbYNCT8yH9JzTPKn16pgFcHcuZj2DzzhwCt6
r48GWQKWUcBmlNg+zLu/ZNSvt679Xsp9ZN8pRwhmYTM6sZtM6AYR52eHyACOkzEt
qdzNqhL/lHR0Giibn+riJyXPTgTCC5fjVxeiY7HY3AZ5blElVG3VxQooa4KjNMVT
/9gSzk96FbZ3VSBcLPcXoDsNqfM9VrDb/MGCCzQNpM/x/1KYKct+OQcl0OWv0LDQ
H6Erwwm4jasgik8n2Bd7JiqxxH1Oonkyf85BAKMtHHSi2i7SNtgby2uhCOUM8qsB
ghtJywIDSQCabF/HexfcJoRHyStbAp7DUtZpLwL9IDLQb6OOmwku1+J0//L5la1b
o6tEBZTbca8rFquLQpxf6DqPBUZ5WYdkY+3W/WO3NH31GpBJQzwy3HdAyy86Byf8
u6Pro1QzGz/1G4E4XksuBrSpqxRWZrsBLOKO++zZBkvSuM/vfLlVYoZInwjKXXZs
zjyM4sB40shH0+TLRWoe6IlN8O1vGkHqXukwdA+WKpIYSWj/Nq4lKlp9CzxI+HS5
bvQYiJKSeL0R0yWufqhvXu5cCVAYxtEKL4yV5q6mdrjTTH8hshCCPL1gD5ev/9Tw
35Ltb2fUcfMZN5Z5xSOTChdatehJSQdkQ4k9hwVb+/dMhqws6cGDGMx3km1nZON1
uOM89QUe5zdWEWDjRWgQ6uCmiPcxijIV6kTRKkqT3jPzWiEcD9WuXA4xNbvXPzbQ
1G2h1ihvclgEAwNaONCWGdpd9INrWBnJgZhmnLW+wDzvTLndssGVfxEcBSLxm+5f
O8EwGcza8k7ibLDWbZ8VnYu/Dq2VCLY9n+Grs+ooucuwnK1T6ebjVZjs/Z/2PnO6
ozG6IgP6Hi/1GN5acwWd1ya8hDFoy2WMxcle5E1vdB9h9O7NlKdfCwBm7nJYra1R
en2TWTBDdwJsNfjHRQjgJmUy6SHQRt9AsTz3YK6vzHPFzHw+fzhAt6eJ06TdSZ9u
0cuHvDtn9uSKa7pUzhGy/NX1IkGYJuH31COHS18AR/ZIZs93OecoLGc0ukBYOJ7Z
dpgNWWwaF2bR9r1r1lnbynfCefCeldtkZFYmwg3urKwdoCz8M5pouLy6w1dZ/eYS
F76Y/fQpb+sBDu32sMNkebR14rpNdIzv7WNB8kCOy8l1NTMiy7XTG5vjauhfHx2/
T+l+RdHKdPwI9n1BZBxxcok68jGEGBcQDBi0YcHVCbazOeKMsQekWOk8gcBZQ1QJ
4szFuxwzXDjAfUUzQiPvx8RoAsZcx/DH7/h72uEbmVUctdUIQ3s/UqccdL/VNfIg
F4gqH7DOusCx6U4WS99OcsM+CmQkI80gJe9+CxjJJf8XXoq44Kk4rVnxzPmljqR/
4qQ2xSAifRuUtoJQmqKP6eXyog6UHegi7NTh4fYwwWhyNQ0ovvmbwjRiJ8dAszG+
XMJFXpVxAHY+K3jm+mb4bg/N9GIkHoKEQv2hVC+tQ6oNAHD5MDHKQ3hs5FIYOnxY
U8IJACrSLEnNnuzN9BKhNLFe1Hr5Q1thlEMnc7XQZ4aBPX5bEqoUij9Z5bhdvkNb
u16nasxidtSx1puHCCQAaKmsgH2uEbLtC9Mr8Luh/vWmFEz2JCn7YTL5Fr9P41r8
ymmtvfoaOjpGMcVzqg6M0xvd2Z91wFLVUD79jEEWgbDCdKM9j2bWbKabl6Q0mV34
EoB7OmitDHir46C2JXDPDDjJqGpg0nfz/hx1T6UDcablSKBpDCRNabMjlL4EP67D
nSN68myOWcF1sswEbhmX0TRiekbWUlx65e9wL+xvd61LTIdV9BkPaGgv8Weqh2M3
CHg5FL03KpsQjb5626SUXcFpxlX423d+6R7yJjnCzluQfjCCT0rjJPMH4+EUr5wy
HjUh4Fm7Yk6uT/sgffElFF3drhwn3L3VEI/jIclcRKkelNMKmgvfYWXyAB+0VoyQ
E2ZjXkZlF21m2J2+lKCI02aeB1WlY7PvJcTAE1wLUufu8wb1YLGB58kkHgSIVHso
HKRbAMGFsTvcBROZOtMWUx5/WDHbW66tr3eezqGHWDv/xmFFqVr1JGw2tgyWnxWT
mWk/gEDqrYFVw9xPti57sbHkFyS4NJmXGXrqyKquoxOgChYugMNW5COSulMQzKoQ
uh+5AvR+4Kr3LBRETi0uCTYfizIdM5QDpFLNzTTQQZ6L+XqlpNONK/RpN+6y04Pf
i40pe2gHuu+qyoTQceY7ufM+oAGL3mZPWmwBS9zAa9L1KkEYdDCaSoC4hiIMiZH7
B/pPs9vPn0ew2HwWUrueIAnaKA2ZoIJY8s7lbbDNStuEwVzHZm/Gwn1SAS26Qks0
O41tyKFLE5MnbzCej2JD7j8oYzAO8yhfZQpEAdn4VvOPH4FUGW165rNUbyPUJ9If
rZxhZJuHjS0jx8dDzhhKTrHJdaAl6zjCd55grtROzFJ+VnLbqsqOvpqWBeTpnoBV
zPmYBQI9ApQmaZqQRiiAodGxmgZn+aPgeFHgALEfTcBd8hv6L6wG35C+0WLqaT6O
a8JssyXYx/IKwxw3tV2uvzr2e+vXNqqaOfUij9c0jjl6Z60ea5+BZVFh/KKhRtm6
a7EjFksi96li+WGWgLCDIU+NEB3htXJ1/TamXeZQ10ce0aEpFN/+BsTBIzsx3uMu
TbfZe3YU3qjARHsA74RcmvcYty0pc4uRsWRspH6yIk2IO7nrdLvaqB0Btl8wJdl6
e333okwWCy5tpE8TkyeQdFxTOAS5w/u6kXvjh7aVTnQdd5SfBxwn2g1Ooyn8D+ne
5GAWfHoe2LxZs9daNrBDvIxygFm7f7z1WVtNAYNE18XoStH4yfWHWBR5nDbIPyO7
LXc+hCRcV/sxo898OqOF0iBzGOKGiEzfaNfbrUiFu+yGJKu258H2Lwz7fEvjiFoL
ALbFvbEIw5DRPG9dnj0gkKWOgc/bCyss0XYbX2qOSBDYDOTjSVK2kNt3OJbZ/Asi
ab4rllvUydeHtFCTxko2eu3isNszLFoLR9jepDhzBXextUKMWuKGY1R/efxhhpJ1
BoFoFpS0hpBgFQtdZPmturd4oO6e0f/LugKRHpKueTlukOAPm4hFqyQcwLjMSmwm
fT/BXlTx9vrPKma4nLUILHWXDo5xpZE4C91iwMM4b5Tyyv9vVbEl3hJCFHcYZKDa
Ucyg9mMSzR96aqbq13WOxlGqsR9pd6GNIWH62cumWh6Mg2rUnHJRalueX5CUyWPg
HxeRWkagtQyCCJN/7PoBcg/MJWPlFZx7cpLYZ4UMwSJFU8lEGX8AekJO2kvbiAkI
FVI05xlSGgnI1ks+LpcTKrqia2Xo4g2dMMNRw83kB/30JtIhtSHvw3NXdWflPayi
X52RjF9+98lQ0VcBYAdMsx6IDjRbE9zOaEBh9OCIcdLaP9AkS/LIr/h+wJDoW5Z6
AtS4OIcGzHokZBg/J62DBoYScNxEUudBAL8qNhtzfrVy7d1SqTcUtwRsRYPdvWqZ
VsEyAmFOFOzXK4e3T5zvQNFyxCHKJEvMZ1WYJaJmNa/lN1XrX8kc23/iZgZsxtkL
pOv0uzOHD0J9L9/LWobj4r7ZFMB4YJKoExOmIYVHYp33Rmk4RD8OkPYRaGe8YVds
DHFUQZaDjFxNF9XAGhy7si/NEfMujquWNFnOCcKDMbxR9TzB5u9VZjPs5sOVOr1K
KtZlvj55gGVIZNr48NDO6QJqT07qspg9NWAhHRKMP2SbVikDNJ/G3g2hGlqoGTBz
mMtA+tl9P6PYnm2I9Lyi41Fc7fIz6tV6W9ApLz9DIpjgrjtLAS0JwA0RqgQru6oL
4LDSCuz6jEcM3Lfm/8ItMGQtCCR25HpJRTONuWPv6rgyfjrC+2gKCtMrYZq2ZfQc
6rHnUUTSlvJ0VtJYRkE8uqeFY9UY/M6paElnmSCFpYfWgT5i/J7ZZ4x2wA90x6zv
A24Ei6UqLOQKnDx0ergjFWnF59QX+r3uA1vZu0qN0nfJMnM3IA/d+47eSiwZxk5B
y+T2DoBdhuvUWao3zQhMLFAzWFmhgpvJWg34Zn++39ExCQUit0VDSgXQICE9aqa7
2OGv7kdNA3vAfjeh/grAPvZ8I6/7DlqBx4BApilptMwW9oqN23UXv9+5hV/O2w1z
Ep1Uch9OIPnMeblY0NKx9IzH3Z9i09EPxFwK5q7f8Brs74oO/25wR75Uwiyuu0sh
IMDflvehhygl8pARZd8T+tZyGZCKuYiDiYFKCY+GERpqG7rXo33SaESuZGT72u8r
UwARX+PmgC54p0j2j1RoU+XpC+tHGh6sE5PYwz9dQnQDjXlblzH7g4d4AbXo5HQz
DeaFeNzDzHckpTbhuhdaiRxFKeHFMxC0MrBxE6STRWn5I+vGIthOW5VLLy23Wter
zMcSzlRZc5JqlVuXiasmKnBeepvrrqw1L0C0/Miyw3BY7kekZ84cMWlqBzvRGgR5
WyheWPYIK0FlEKnNF+JuJZl1nSeMiaFvMLtQcn46nWWPrD3IsE0V+gvhKPnXepFG
LoWEXnxUUnJ6z1H46zA/Z7ZMDeSsEwmKdc1HG/juI3nTDUtBIVe4PJjIufmzJ34I
johegTJJiY86GKVqj5FfAm02yan3YzbAZPV0wLsAN3nuEF5jH/jRJ9S27X4XF7K7
rk/RKb7Vd/EkDDbZ+XaAah5Q1yQyneoKqiJNeiJjoYHSuu5mEZWO/qJ01b+Ea6RR
oIBYMhzuIq9iGCz6QsdbvjTdHzXMPcgenfjPXvxVPUabDBIqWs6gAJ3V/etH2voC
AEiqR7sIX6licKMQRKyd1q4+p0bCoudNR8xi1mnflSWeyU+E03EVolb30q/ZPF3z
3piONWLhJCCjx6Pc+mWykc3IHPDPuP6x2xLwTLl30/275zVsK2O6wJ4Ni+AzrfDP
fhIidd1YXPzo+JlPqiTUbrBQFu/pKKo5+AVIejLZZiQBZW4TJ3QMWIISQG+O++Qa
jqSR5UEGGj7WKzTJXe3T7PeWFdM8Yq1yrdNoIaVfVFqn1HIri4NBuhkkv9iQqw5B
U1DhwVxmg6dD78C6UdKEjnKOYjxAv5lRb6CZ7nPlLrMmx2lGFuFxYtV14nfsQvgZ
RwMR3NxLHa3f+H+tRyOhA4zO5vsOcERcnpYS+9P9yjmBFqQI0GS0GX2eGcPyy0EW
EfqUaQMCRb93Nb8BqSCOroGeA56oa3tF8FSEUFqL0PAO2D5uiFXRgeBLJ4+oVeuH
4PVM8g7jx7ndZnPMp3gg5gt3RWL9F2rO2FL4Gqf5AEODsFou7mozy+d6AjDnbXFa
uu6mnYxXSxpsSG9KqhUJ9TgrV8oE4p+O4r0M0gAWXAx/92qkgfQElpTEtMrXMfWs
ruE5M3R4+frkAfo+jpzaisY1eQ5K/CyXigEedkiA7Z402kM19Hg148KHJBSpnICl
8mVeAU2vaCfmkcA8h7gixhp0147zY/5UbJRI3qkNWx6TvM6MGOxc07OotSEOrCx5
CfIdF6AS7I62YUMk/dnyxtbFb8BvI1L2OHXmB7cmhwqxeacrB5phZlxSdstL/vOs
1TezSoKM/WOjHGdSRSjKFoRsLAVfAVMfyJ9e6VngnPXqz0v+aAQ69iOU1NSDQgpw
g1PU34FBcDr77p5VSCWKODEgutDRbZQ+S5coPbuoVHTGIHLPNWq8OA3z5jT3Bpf0
n+JSEAnCzT0uoh/O+N99cyL/aPEEzHf3yBlDtU7BI9IcIOTDfA5nLK5S1muasZtf
71TkxAi1/GEXm7DCjFXzOav2vuelJushQVNc/NsCBR5FX/F4LhEZh5ZL1ydPfkjZ
IgLDCgMutcd3leBoUFcvtz3w1lIhO+0kK9NfGSX5lojrdjS/3dfWffw8hHXXPHam
zPpB1+AOHA9erKEjAMEDRskq1DwBHHeCatJLo/2Qs3rVpmz9KyP0uwOGIc//fFi0
H1/dKeYWtzns2BPD2KWVxR73ZaQUBiuuCtHRSCuGr9a2jpbiek2XERxhu/M0X7dt
z9JEUcEpvRrt83mPxhEG3v0I87rU5khsVwRmB3vCt0Dd1AogO1wmXMl6UO0oMRaR
b319biBPsl6BusacVwTLA0vGjJYigA0glIfwbYf558UnW29lhdGoxjb2CRq4HjZu
dRQ5P+0GT2d3zdpE2p5jrc8xi9iOjg6ieIyqf6sDo+ef/rViMYh1ZdM/1mHIo198
q5uWpTzj/CEUmxbaGKyw/wXF4ZFBkpnSnNn8KLuM1k9MlY+nzn+BJJbho3DhI57K
i5jfIrXZBDn2JyiwImvd2GhfK4nPHNMw7O/fqwRR5K0aunFTzzRwr2zyVBGayf0v
NxdwDmHL+PTgJEFpq3IOqYWK68EthJ251+XinQc1+BPDgrMv5aTMkXwB/bj8GPrk
kvQ58ImalTZNo0xugpyQNfcT1m/U7TUa/dRGgbC8F7F8YedlYTRu/cAgcorhupUs
r9DoItJmud8qRP6Nq418gfrW+TFuKuNwYPJ7Gp5jNsf2Awx0C5ZWIbE6ZhlwjtU8
QbYMy3aZcd1LqFtooD35z/Gdr126aoYSPGp1nTZBr4RJtl2UYBrSAlaE8hMLprWs
FJImF7jb+kn4lFQ29QGuUava32/68TA9Hh9aeu2G+eCybHF+ADFJHIvw3zGGTZDX
/wiZQH4UfTiCqgGh43YPs24sUjO/ckQX4QL5z9e1oi7yGHFS8w+EXBDmqiqC1h7L
6TmKKzeQ/8h/n8VPGHa8mcP7YWmrQZhJFzRE2g6rauck86Tx8dYLJkWTNqY0akHp
j2Hb8/pB5MaBzTxha8vgyiPEm8NjzWBCLVFpY/ZcjhTDS5JdH4iCqhdgI0RMUmJR
vfbPZ9KH9uNm/4QeodXyDmD0Z5trlKN0LF6jOlCsbhW8WNk/G49S0IIPjogoZ6EX
DOzxveZ3HYBLcCvJJH5/MVGf0scL5tTvQk2WlrSE9E3w2EMip2O3p3K7UpBaETss
/Li1KL4/jAvo22zXu7L/NDWAwQueiqVJ9JLGJ0yUrL7DcVA9UbMqrmjbsjuZkxsC
CnNXJ+vKm5mMZD8AJgti8vC23kBERh+LNOg6hG37IXxTOVk9ikl9GjbjVnK9LJGG
uFIT8vB7//wN0kpZeNBJjKCVvpl2CZBfivaRcdvU+AWvmJFpn+JlIEeJUqtkBkuM
r2+NnH4/5W23hmssRILKzdxH6U/9nJJ0WwVGa/mQpt3WkrhA4eXRI3YuBKL+Krs4
umaNhm5mlBG9ubxKg3gDJouS/QoKFtcnZyJA69GVroPYYLnOD/gm/7qvJeqRF+Ae
DzGZ+cz1W1I1bpF/wZZe5dh1OKkvgm9lMR6o1HHExrtulBHDejG3XiVve5+ToxxN
UnILN4GgMITqX8malPyxvin+8xeeSzEDn9nBPWCSxuJjT0zVr3uMbU9myB4Sz+Cg
UD1HQgF6CoF1naOgr08JOEAVxalQ+J0GBU9d4JXUJLAdu9yx/1CGI2zfeR5qKiOh
ws8K4myVZKB1Q4+AabL27iGZnEI3Bf2o0DlrWRjrA8uwM5zR1yQGBcDlN376p3qj
x3H0yioXA7wFaNqt1rJvsxVHBEV8f2wYTHHpcrC7kpAqCVUwXm0tuO4hQMKbr1Ue
p7HIVCqDNARGwhAs3ZibifuZiqrW9yxE3WdJJOz160GaKRPKd440a30jLDjkt957
21Tl+STbwh8JexN63x7G7+98EaEbO+WWefAlAKNOCY2hqUAznq3tPnDFYZaMwT51
0zoADBbucN0WwDs+T50sz8STRYjcEc0ZxG6s6zVMhUcbSa6QTg7h/gqpZXxdz0CI
+m+DpeGWXbmIplIFGMOItLGC18reCjxDhb/87ovQvhoOa3m9kwj6zoc/kq2n7L+7
AUegCff5DgH3qD2KO3WRQPPyUazoBQlI5i33FlpHJI7G+tsaysEufzSdnb7pW3Y8
Q/LArvoqbPY9VicfOMYTFHaYXf8in1VW/0jgdkGb6OGqx9sf/R9jFW7B7ejOQeAy
2+35JU4ziQZ/7Ee+tJSeqscvQiKuO1KrJyi5BU0w3IYObeUR6iE8AqCL8MYIsXbl
apqLXXHyO6cAK6aswijDAtzm7HFNzPfF6yeuWyeC25OBlUbh2QaNclyOBIfxLG/O
Kf0pU6LOoxRZ3BecAPtu9MplWvE8b1QIUjcQIHNbYxAYcMQNf/b8mEMfS2Zbbhsn
IcjemOftGO46sD4emgYUwsGu3CnpEn3xNZMlNJ42Uf8JfdfWpoJ9yvDDPBCtZvZa
xlWJgXwHIWhtYhy0JkL5Vv9kFhB/H28o5upj9kBp7XCdIpzOHFW+Sb32G2774M4g
ik3zVe9GldPlGjS3CZr/r0dBeqTQOmCodn+7h8EAAAPRWCJauxnOcLOkUd3hsIb8
RnUjXubM1TNoN/EkmP5M31iYDp6NCm5P/sfEAQIn671t04NRUxQDqUg8Lc4hKRYY
BH7Puiv8mYG9kPNLmo6dsIxgPNdqE1MGvJEKRLiPucJGcskXAcTD17WgIUpSfq28
yipFczmu2j053EOWYB4kp+2GFAUC6Ls7jTDvJWtZge3vfPG5R1PwSYWy9MXJDBw1
I4oXhEP3ZG8dnIA6GsDCFXg8zBygIXLvJzrD7XYGNH1XJxrH5htvMw4zZ1aMA6e+
uAqCxW/Hm62AMzShmRm3dEXygm5IO53TtuBk8ZU81WM9iMHXWrTuYeeHg70rn2PI
vgHvr69MMcLqcjGXHIG9FT678KyutmfWTRtIAmd2qX/oHLuwp07B4HyD3BaRBlh7
0yZmFXbyhRqp+d2v/RrtxDoXu4D4fPoxVYKxwmj9r10fttSqILyeKFNIQfKXI1hc
iCNIUgTspJzmvpRm9DMhNXmibDSb2hyNLeQ7QTiuOTKar+VCL5wEJ7iTyvDvcPsV
AD289QRe469VvOMxTS6Xkbq5NXcb8vM9z7+P/p6YbIi4KJEq5emEQ/PBRvE51Zoz
cTT/st4erX5JViagzmXWPpMR44m9Hf/yovLl2dxWB//beUQF8chEvprYjPL+yPCx
jlcNL0YCrh3xKtCytHlmdZ6l7a0SGtr3yB17ouCFipRm0ZK2HGPBb5lRSIhfui9i
gtp7HT1Fo50hGgeu0C7ugxcNWmrZZ8JgAxNrYFbAuB+z8D6PigXsT4RYupDE5ydg
bXsTzVScmAOFRhSkaG/1Gw1IX7NNIGWWMAwL7RZVTZOFXj+lG4FPMP2bLHdKU4Dm
/Tx+IuFMuZBK57vKo21+/esWHUNAnwhxVFbn12iP5TiTwUKqsfLDlliUU+3VLW68
jGGTLhe3LCW/FinNfTkHkXmfdmRY0WJh6Bra75f3i30V6HECzubTSV22M/bxY8ba
XbMKxtAedSwzYCS+2SzoET0UyCq+RtPrOBBr4UrsEZH+LkjFRVKJKc5mjk/LroTA
TretSP7ruQAIks8HRriHP9zCfNGTJCmXtJVmEHY2Yn6NBSpQ3yUBTxncA0ZzVgbw
jpFVi5FLeG09bT7q/XaqHYbCcJQNqy7KOV2eLdmfWTStE8ItxeW9bmMeojMwv/IW
25uZGW7IBK+tQWeNTokbe50YLg3tBUbE8hium3nhboqP/9vAnRSC0E48UL8IegDl
rorVtZ5EJevpNEJS3Wm2Cy7v96RomGPDrEu4YW5//iD0ST/U3iG2WpUE1iL0t48M
TQp1ap5nHbrP7akvq0JIv8Z8UDAKMiAnQDUAl5x7g97oGOZ3IqCtkAU7FIGuR8oN
QVnCj24TBA4pAs7C6J0ozCtZ6//t+MHVj1EVHHHMoyzSy1LpbHHFcC0w+l7GQ/UD
NKuvkn31iSOavjsa5pLd3xiQqvs6Iq9BuiFuyfZaYzSFmvE7XVCelcFLkDhf37Z5
SVDczr/G3awgHZdB8LwEcUzt3clotil01EUk3myPCStwrATx/qxVrLpK5dYjs2Wl
DrtKlpg/JNAth1euPjuCciWCVhjVY0mS19SXpz0DhtnGvOfIyPftIIhYmJgTsB4V
JqOAZZkNERMHYDm6d37jkSCFcRUw6TDCZAMGbzWk+Piq/3ODwmbtOxAYO+vZPZcY
m2j3MIF7jiiWvEXCgkC3JbLM8Pi/ROKGXImpWxsKmVgUBOMXUhZp1wxepHFENkBw
vYXD0CaPQAO6R2uJycIvWRl9hRiEEvD3PhaDt2i0QrqWIva1u/PY5NbWqguPTfGS
qEfH1wEI/wDV21ZIxT1PR0xKmiql7W8uDE0a6oOmpJvKW6LaEXr+OxRPK6E99I88
rxkRUCU6KF5pzgjNoKbtFbjn/xOdfoM+3/7NGhKeEcusebVCqrvVFr7DkxNsCgCK
ojtfuAzecHAScJa8NBYvHAhaL5+toy6AkXVSGp2Qmp/XLS52jWzZw/HvYhg+bjVH
+2SotFiR/W3EAoBeGipORkysBlS8c123ODXlvyK2DbN0cU1jM9CUXF0fu2imqxNL
1BGfZbicXFhu8VSNSewyc5dOn+DPKBAMfgl3o1I+2QdUvUtvZb2o7xus+cC63PwU
whJNO99gHbEk9d5Xk3Uqlegwt6ekhAmILt8xoCuNvFsBA9EacfYIorb1bxbgbD/I
q6KKq7sriFJtlQP2rL7uIj34PPtkDchSPCh+6yDrPvFFbTiHpwlsseL8F33ACGhe
uCs9jAtFBWoWLOYPq7VsRaDZuzgPzFw9ZiC5ADiTmbZd7IMNnE3p7VW3A+SyNVYn
yEw6OvKQ5a8OYgmtcDa+PhwldiCGrzKIcL67CSoWqk8NyW+SriSiyPfFz70QvTXa
s6fbUILSGmBixYeRJ5XIuf/h58pOxTXEthmEK8apuazosP0b1tF7hzpVE6wRIoRj
DF9c/4ikys8jW8FpA9e5J04JywrO4EpSjUBZ201yf1vVIWpidQrxSDTH+cNzr2uv
2frY0LTyPoI9p71QdACvaK/WHZgDAL6h6DCYWOyzYSptWCQqhYki5DL9/u3ITGS6
biY355awZ+WzVhmYGI8+5RgL6tzrmld861ITR6VftrteA8yz7bE6bbDz9HwhWxqt
N8EsWRB71NhAglPH1e1YjKIosSHI8mhHctPuo1/uVYE25MfStI5dJL/OKoYeX9wD
z9+iYcYCAC8itaUaObunUaPNUBWYTeAk/FFjto6PryP7cDam+J0lV692Fp7151yA
dUH/iKZPc+u0YFwDl92xsXkbd/pwvv6T4JEUxP/o5vOwRCdaTMXMMO1EA/ryfq+r
mMqncCbz1iQyopXLiH+B7t9eag/60YjIm7APKbzT1S1sh0CMtKupPUp/u17La0L8
3fhiNaoQi82Bz5lZaCaNwHk4Ih4DmJmozVBuCXd/ohltHJAIth72lgNrykSZm5R2
B+HMYm8uGSuhF5oZ9FFlZQ+Tw+L6YzdtJnJ2p2d4IOjx7L1kr9Cxze40GJhwhSxS
orV7D1X0ZEu9dU6pk//3bu6T6enmVakaIS0wBNJDQ2/peB1Lk3fakJwk0pG1rDpb
hdjOeax2oCuEiFidH9NKtx6hxiehN6cYYFyJo93Jq0ia0FhPF8FZebMzsDDYnkBl
+MP4ocD2wWvvFBhORaXNMnzFe/c1sYHV92Xq3G9HlE9bb2wnQQCFOMVfwKwmGeW+
f7pCLQGqcdA/Wsc85Opp9cO/GISsz75drL2lk+xVp60X7/51ooN9I6J/DtKC9U1y
Ed8WiJzUqSInGijB66WAOwBkG/gWAKxjemtU0Q1dKw0T4tWyGA8DSYArgqruUY7G
CFNWM25spddKk3jP7p8+m7Ev3GMriDhlByrPeJ6WqF7rONPO87eDBv/Az+PCqGKO
BWHT3ClAtJP4f06SIQ7tG51iVTA6eNJrpJQQ8qEaE8T3G+llsUbuIfkKTYBD2DCw
xOzCYFt1FqzUmt90qnPEhM1/hSo/JqqUmihtFKaZQ+zY/ftKVHFxNrOKR8o3psy6
euilWyq2ELL3//Wh+r3TDz+AJI8Zic18pE+uW5eIsFPli2t0HSXtY28QcsyZuVZX
G2suraNhZrlKg8C6MiyOceB0OIhJ9U5ZskkVYzLl1HRqIdcghhyUsMRbHexwlDpw
ZbCHke1ih7v+IdHLDX3HvnpCYxoX5CwE6jvMEZwSMRNi0mljx3iFiJ9OoDF74T7T
HhF9FDaIfStdp1Ejac1sE8dBd+HIbwPTUPISMJjDxabERYwEgmF+j6PU27TfyrMb
nx2eTWcVvL5ePMncwrkkphtU9v6HqzEg/wAGNml4ZgqdKXHYQND3bHvLjNjjmbeY
QO3IG7tQEzLzsVfD9IOpV0HPnka0Hgzy8qydjVtGfBqZKKeX4cPCVyJsjj3kBleL
beyENEMSQOPEYaO9ABBuTH+KiljKNvzC7wv7r/qSg7twHR89amVyzWkivUDKxsIC
LvM1jwALGlk6zze5eXsGORj+SjIsnXiaGvNFFZ7a4Jjj1+zAQqMz3RnAaZq2QcgX
r7obpNh2LAIXSrDs0F2y04lCAb7FUFBT3+CSfJPEWACutyY/wRqEKIRuWRsUs313
5HRaqVoAcrUZG7pAIOSl+Aj49kHGXaVE2BGxLAtMHYl+UlYA+oKNJ5E/i2B74S27
xN1p6R77LLfEkG+TkH6Od5SXevFrzjMb/vJbXAFFYtGRKx4oQb1+FFc3oT4sIqZ6
cQYlHnIN1pHT7Ft2H971aOmXOOB6Wei2rrn1NkkgbCukZlGXph3CBxVdpSW1yD8v
NgERXLEE8jn0JZMopMlnew9u0vRPeOs/5m5tLxz4EFoj3gZaMgZagL+Y5wJ1pLV0
lG0awysd1SynmNwNujiMMIYXjBI80W3SwqC03NbTTBH8dmCeMpXZPQm4R8lyUf6t
C2Ig/MaXC5hr5/6zrwi/WW9hBtBzdIb+t3qjzeBZWac56vp8C0GBBWPoTZio+lDA
IV7iMo2IUGwDOSZND3s+NAlTq0g5vGLWMQp9gfE5hQ7YSCbeVCLshceVHuHBhLae
tNzwP9E2YgZZv0r8gCzZ72UZaC8QcfzIYDoKwFp/YdxUxoBYORLFxutMOy3Db93n
OVlmETPjJE8U46Z1P3EmZny3pRT+Y59e3e0jkkA6660f6xMAyg9TF6c12JkUWo/l
1Bc3B2yJ/UmkxCI14uiCsOuaq6LX++0MmnzadzEh6g9cojEokj3fVb3kO27+RiAW
hRurf4HFhkVk9/ncAHTYosr4gNrOP0/eqLZ2BOA7Q0QJfpXkNnFc6VvoiJvVeTJF
1rI2mFI7NcXnJt75OkNtfrVNSJqIIAcpQhjfS9+dF2J2ZDapkp9A0g51iIVN0JeE
b5s8SnbykrK6GqEw9MP0Kv/0nsK4E5o834+xqe2KFGHNzMYZX10JeoMjXg38FRN2
GqAZu7LbLtshN9XQfc0Lnn46i+zmdN41kHS0Ry1Mb+G2X7//OmzyCyE8DQQxDQ8X
560PswKF6D5spVsH+3ii4FKnL9++YGgfmurIVOOPvK3KmUNNzsvXWn2X4FU0QYhQ
zdq9WrYsJrLmnkIZDAu6S9WpWACHYXJJ/+NJmIab/3lB65d5rUhMUBTw11qkHGAJ
vkC8wb8cJX7wG3zabmbl2d2pjg8t9cViBfVFvWMprHV+jNOf5uN02YIxwuseLbfh
dafBO3VAOBFf9UjpCDMzfLFwaOzwXl3duv9Rns7yA4TarYn5OthTuv3Yb40c9xh0
AD72ehdghj5URl5YwFL6+vNher6TdDiqKm8B+eYw05hfubx/04A8kLhLLi9qWdFm
ix3AY09oQKcverlihxJzSAofKSjn1EeANkuCZUOWUAUazaZcdwNhOQedZ/LI0YPJ
0OqOYCrxprKSJxipV30ROxVz5CDDSB7VJVJI+eI2A/qmT5fWyM8qKkRQbi8xKxqw
s/cbGaagRFIUbNfqFy9GySqPCV1+TuR9TH/89AF06ZqosVGgvqdBPO1v/7CEP8v9
2UD56idW9r66smJIGy/mAnmlTNmz6cnUuKiI8Oeyfqf1ntanvJchv0c8RuLnvnia
ECERoSFXNT953mChzSdFiEbQH7kfB1Du6T6xC0qsfFia6N2mwU54G8vsONpTAJ/p
XwJfenJti0LZohMEmJTh9jhUErA2CzED8xF4YJVTViA8WHTNZg6mhCtmFjOrxM6L
zWhZEnHyICteVqneEo2ax3U8qMA9WTZg2pl49iyYerc/i7jtNPm+b8FICOv2QtOO
5jVwqlmik7RcgDAi8/3rWR4Y1bq3KupMxay9401n0s39uuPkEYW41Xn9DrxAR4OH
xTFWOEgcM6Ymo/QjkjtB0oMIixIN54yX5xTQOKOyLjotOhblutMe4cnjN0NjpkR4
yOr6EjFlcO+plzsQ98c8Y6eQekJMYinAGVeHGJsT/LXYADqOcSl3Ff/RXIdK55ii
imwK4tboa0H6iPOOyvuQBuFVWW9wXzwAngqKPPNLA14oIjFm+H9oqoXpKjRhmhih
4gcnXc3xE4481AxywsbchdOYtauoUZtHdUGJi8M+atrHIp7EyI9d+BJLrnYh+F+5
RBUTK1APUCXmR318I/NyRCSFFWnD7Kuh1D7zT4bn6LYmsWyNQETk1+0jUMnpOUn+
wL1QefPOP6za7OFexD3xdx/vAkvp4X1MuYLLFDwydMhPuN0ZcRJ8tBdsnDMxQ/kw
rJD23hcZZAMUfc2XIshX/kdultGBqd5tG+MmO2UA9gjiomtlm3z1fDHMuq6cdcpp
ghlUEstdQh/urQZZwZZjmZCm3lwAfCKMOBrZS/61mx5EQNBwnrDrpxepP2UGW2UA
KvYT94EteieAvomnjw89c9PNz1b7BXsW86nLFpPpnCQnGkRCzhOCkLVGjPj+dOBS
AxKtzBjaaoLEyPQAzDhVXKUgB0XnPE+kGmOtO4qY4iTfIMSr/QrE4KKRQ6hwpVuK
4DQdw4jHJH1Dal3B6iufBevIDo1SFqB7cxjrHwiBywR/pSqRFHUYneGwtlmoNZYE
7qaADMElkeRiorZWRDOkQTF0Pt6/DMH02Gb8sjn7dyC7wqic2lKWLmDkDW5Ms/Dt
NzDRoTF4ocHVVHE42dnkqkoLFCYk/7m2VdVQSsY1SFba2GFiGlm+L772tALCx347
nwyIJPLurykC4kpHGMk/TuqzQcTpietjJ/G+oBNH4bWfLnsAuCA9L/Rp8luU56CF
9AACCB0bmVIHhk6m3Q7cgonGd4vK7pMCthUFRsljCGk1Uq2WmtyZkgdmYYoAAnqs
/CZh252aMxjVkXpvDYac4j/6Xc1aAsF22pANFjOR8G0GbavBK8M0PQseF8j384vr
FD7YND3x+ePbtXUQxLwLAwXBFw/OPtmsOhoua93JZk/5plfOiXRpTCZB1SNIXwR4
7PEv8Rv3Mudiikr5MIcakfDrV+HD6/eSe/dE0WicnHOOJ1u5S0hb5nkR0BoOpGty
41+I9IcapzrgAqHCRKTsgbUkte72/ss2fhqd7BKdh5853wB2+twLXmhx8Xv/J9b2
ZKxma/qb+K2xNoxI9zrLyoNQr6HGjkPg/DcgL+4UWyNeUNoNTbCNnhFdyDYZudZt
p+RM7sGPzgKLZBA6tYizbC/IrhCM3+nPb4N29apOvne70HzGiSf4c0xTf62gQsQG
9PyCoXXNJ5qY+ZjAEWSunV3U5DsNTKV5VmjkgFKiPSe+YXJqFRjlg0i5b5auYEeg
eKbo+BdiJRl+Oi+ZwyVykXkPUQxNAu0l7mv/6cLzxZkrFkfZqtlHV6nu+pjDPias
NOyZcrpJi+ZZNfLfTR+ayiiSS1heJOk5IJRPlacg9IqDDxgaXI741FsnJtDOs7HI
9CSOVBgvfUuopkm/PV0TgtSr8TXh0UBrORnyezpk269Uv5rGtuZP0Am7qZpZnBJs
OAaEjurYMlXtfpNAeuZ2adi0F2Ln3+ocwSeJns0s4q00/gOBuxZ8812yDRVowkhm
SmXZ+WYjFXyLPJj0YkM+po2xLNnc85GM6W6smhosNC1NBVq4quh+LelkBWxNWkvw
W5DoCFy0j1jdjIn/b5sbZHnOY1eRwbUX1hrfd9cbmJEiehP1/T/G3rk/fTNgFhPq
j4BzS4jHBfU6gOnOZi3guPy3KfkhPP2qOmXkqmod+wyduVqfgbdyLWSKtePK6IgG
aJdKjktUBeSUcikVwywyeqoInaMPWRhruhhE71d+g4z9+eQksEzI4pyEsoTII4u8
uMpoEjCe5OfTMAu+XoqHaGgUT0Nc7vSUXBOKrGz7kA0OIqCWa3HtFh/MZmuSFMLw
DZBMvXZRpbimNhyZWh2+7NcObvF+h8hwapxpzysGt23Y1LfcAxX7I/WLUXM8jydm
rJ3hQBE9xEmHxO6X09hytSsXdGeBJ+v2SFvSNhqLN5O6pTvzSPRLgg081HYFsgrd
3ZMGS1nhRc4r/1LUBQ7TpnRTPzwd7Zrpm3BYNXnCHb/EBRRJFDScwNFqFnObfg0R
3vfyWSBilzdegujAxoJh0vJMJehttpt4LQSPcQfQHw/VibnFduvY1PekAWHy9ONc
l7b41LoFQWkP0DBzopnkGgYuOLh/W/K3uhRjfMhs1TlmGv5l3Fp0xzuk65NrR+v1
R+Z6soUOpsQ/8s/GKykX4d0o4gw7MaRsKmj4EwRlCfUX0IY95K/C8+l3PItmQV/0
olUh4fxapXCpMB2z+V8yk87HS/kw0e0zgskFJU16gY1h/4NwkCKPVLZmvvMq+48x
SOUCA4nOhs2WtIOq+6C1l4jX06R2DffoBzgu9r0Xd67/abIxXJ7IzNGQqc4F5OiB
iZhrrUiBWWgMCAkV/4WgY4CrFnADg5/JRjdhQimSQhUCFQvNLbBhoKOyBGr1giHq
siH+Zc3maLyj6I4aLLSQaRPHaRqcLjH6/T6OVmdhs72o/tPLbqnDtMNgkG/zJZaR
ERQlVDVmm5ej/LfzFz4Wkh0JMC7lnPPNtaqSoRum8PMBnh15yqutdYytv9JrvLgh
sWVqhFclzt+YsFpg2biyvHJrYvh0JR51YFcpmn3on58jyy7xmjj/Rr3RU9liX/qE
v5zBmfGW7YCKWI5SOJGXIPFVlGqJjPZdc56cX04I7/FQ7zKvSyIl6XFRbEWp6BqI
RMNGW1zibcvml0gc5p5roM8d4kKBSgPcF2U27OtfCZqUo8qEKknUwJTIJALlSqq5
V/9qjisbhsNygTypJU/atkOV9eAcYv2uuvclYn61SqsJFxR1oGyPU+c2Phil7/He
oerS59SdWI8WuFGUWLW0mYdMFesq+9iwOszkUG4KHspjPLXQjkj3XE3rDDwLbtnb
A9V7CmN9iS5/OdVnVpoyifvnoAXFuBO4KMmfC+rDEigQCsY0oLahM9QwSKU4Gsn0
CazAsK37slkZ5g+vOUStNzjZmXyKahPc5ASEG02EnVlUU4eKVAeNr0F/4YgTdvds
vH3uBflb8o2KJEAcIRi88H/9M4kYo6AYvUELw4N26IBMieu1dg9eJfXAysnN/B0b
hqqWVjBP2oMrzjXIkAf+b4xXf6ADLUJxm1PnM5M9cRSsvGH4mcjDaLopX4mM9psf
KWmA2Tr2AT4C/bAnxRDi3T427uXP3WKMurCzVo7QyjrUHjE7WZEbvorAe1/C4KPn
mJC1JZYBV/lilkqMv/IvjEKwLbuVCUP1f8fapKFTBFPvHetLos8pidi0IBY/Pj6I
qnxTwzr47ajrzxtuq9Vs2mfAKKn9PxfHczLs7hqpgUGeeoGEd+B/mavR5uCzqkr+
jyPqryarufrR/avChKidf27IiN4PW6tTMMTPNFM6H2LlWiBb2G+lfD6EUsPccDTz
CmAWi5/LkBDIHj+RCO3FznZzSYaOoVCrOAqzWc08gEEUiFRN6a/3rv19DiY8PSMw
uZKQ9oE8AAh/lW3ucBtwjd8v5lLn1Cf9FHqXTW+a++Z85lXcEMtLZZ+ppVhoHwue
hIVMrs1izIQy+dxrB2VNCQnk6waNwZyG8+6Iw/WpXiGFdXnFWXQRsC+thjaNyeCe
jdf0GS5GFYv6Z51Dh91dSprhKpuFCYxA7U3XalzDJlwHYQ3YsVGAldvIdWpQLv5/
dlzUsNJb03SNilBGAbWzx3QvgqlKGzbDOCwqjDu5L41r161pAiKqTOFWxCehmwon
pD0/rqVkOzb84mf0w9cam6pKUxoki4RD6f3IBijhrgaH0+YsCSjGDZcT1iExMcO4
aWwUJqPgO7hfeOuwa95hOI94oeadUp6NDUJwJzmfpsgszEY/o9HOdg7NYGVNL6xM
w53eYch7JEyDn3J1GjBbiRR+WU9Mun90Kl/Iw0ZM7VngxciUR0QptlYf5hNJJoNa
ORrabUSBo09u+da/pjFUKPt6lz4FJzQNjHeEuA2wnTI4B3iW7px43sigRR9xOfK7
3MkX8K7JSB60VmItQOqLOpGCpD52VE7eFTMTW2ThJYcJolMn3WJKQir54suzmQ+9
IpJJJoREh5zs82fKyiaPEKsyZ1pJ6cKCwVqlVB6Fs5eX8QNKvdDeGapANftBjAkL
EkY87otmZl9aoNWXtuHrcrEMvuSu1xus+Y0ykbuRr2FQTEmZlt2kgx6LZaGSxcP6
QwYllm+j2PgecxXmx+qm7dF/OyioeE3sIt9BSrnl+Zw34Mp1Ic+e0uQFTkgOm4Ef
2wi1cUwP16NqswT/i/V9rzYFyO8KQB+noJm/dwmPwnKO1BkadAl0oe1XqXsa1yAE
grMvMsT7V2hzANBvqgqZS8Cy273WqzCpWhBQcrCfA6jqXh03RwTExP9k+23ouSG+
qhtLaX8uTvjZNMCuviwVqtwf+1dDvSemmvq0AU7Zn7wZQ86bJzKMvwg9MrAKFF/+
ScHe/sGZjJXqehBxri6TBGqUMnfSaZg+DYTa1fkYqMQo7sWrSCjkrmN07ZLaRRfi
Q6YHNyBKqsW/BSXbrtSXb1DZwIXyTWVyZrT+VHWgKLTavdKqpdyvFchC4EBRr3XG
4yU1gEYKdENa4D3MuOAmLX3auPq4imZVGoqm9olUqe6cQg+DTqUsyB217zarzRNB
QGJE1yzxbKUo0oKlQnRfQ1T/ggjDugys7x7GgAa798FQcoUSvHbuyFBsN46Wd4Tj
6KbEJzu11N3LOUgIG4e0W7HxSLOfmxlyE2CCx2DHHU5PNxXiqRsLZQrJSvZGwwD2
MpSM8/AUXCsi8afUqF9++BdyzutgGJnkVcoyVTsbJpZ/F/+S67Xgq2pxaeMjV3MA
8lVjGtvLrUiDDwkbIYbRr2OZtCr39ohfapmwquJFoqflvXWLbGaJDIE9kFO4LdRX
Bmp0Ko3pFJmNDAJscgm/SH1xFfS/eQK0zLsRJqt4jQiIWzMjxQoiF9kux+ZguGgc
zYe0QJjCb0tVH/xgJY3QZt9y0mfQAjRj5MGRd0XzEEIyD0jEg2tcHSYg5zGjTXbq
5cWDgWIxyj6fzuJMrkZbENmzEbgKp/Ox5UC9hR/Gr/awbk/9NPKT3McyUab9MRWT
7uVMWkR1TYW57EGa7D1Ij+rpffS1qyvoM+gQkui934sA4+ouytgL8efSqVfcZGAs
hYZcfcZEvPqPojXXcZc5bZoBnnTheRlaaLhPwrGU/HZaIDWVDATMxrvFuav2u/Bk
+9Kw8NIoaPNv94kuM8Gna1hRksDYTmp7Xvn85kxS6nwOHoY1GLlFoyWSfUh2LLDy
76ACoM+GPuNYLDey7npS8gvWijTBbBHByZTRWDyd/x0Cu1vnfHrWkVComGLMUsRX
f3VzMbpHd3sKA6jHdMUji8fJIOfjhYZM7sHYfbMDMUz/9wT3ekzYOOZyG/1oZdJy
YenVRWCEvpMNjvwo0lwWZ1q57vp8kca/+ngbEkxbk5pjr4cDo3swB3q8cTMVUjj3
0WjO1TfTmGh092LlomPi6P75b3slJCn/Sz4n6/VMH7T4UI8IecdREGpaYGv9gnsP
WAKeziP5M2+r8M9ww8+L54M+0Dj7YjdyUDWr9l1rhIJ8ueN2/YNc9v4bAWWiFil1
ZJcICG4tIHe+GitDjk5SI+pv35/PhsJ29CF8yt4Ctfo33NQ7MaiROHGpZmfL+tgo
bJRSD+jWzffKat4kJpewdl3OWQ3uf0IAO9zyoHtPvGvTOKWjHYGPsPAs8QKrQCRX
TCGTlGRaZSyAyh9xcq+xYDxvoRTCaAXlsy+haV5nPBbKvyvmTa/CeLgqXYv1x4/c
FeD8X2Qa0LAx8v/BJa5sFhx+TGCGhdQ/BcOJgFUg2wP4fN/QZZMEMwnmjVCNKdSm
vt8T7M4HBuM9Q3BYffC6DUXGtdn44GDpQHhGwGX6n00JaeOV74RlO55pu4Om93uI
fweBXW9BuUwsOlY7LlR/SVJi7kDAH6OYA/sf3RMMGhQUIn0zvCMbcAhOaeaZUYoF
cg5yEJKplzNtE1IaSs3DojCi/jj3Q0yE4e5cdvRXb0wbbw5yr93QquWAKdp0SuQp
iY5QXHB/rVZ2HwB9X6H+26fH2/fbO1MNYJhDhsloGIq0G+eKXYkWEN44HpEwasRq
gIfzcyvuN9WdKYESvqMrCnQEhA4kuctIV9E6H4+L2CClqaZDPEXs/huvdq8pncH1
QdWmhJnhFO655YRwwDoqAcNdNDWV2epE25SfOoEQy2ML1ZR5NF5oxucc0xw9C88H
XHH2hzQ0oLW47MkGUlMTiCZLVbMu2Tfmp7dNQl3umVVP3fFDes4F6LWgyKxM7Cwq
19vBBd0uJm7PCYLqd2L28tGSsh4HFLZCxLda/bkcfMi2BC2SCP5PZ5KOX93TD6Vx
0bn2VNhneKEvPlhXZdnlIIoMnHnrlL38+nbZAJDu5NMs4Ayqlt7PtszoUsI3E4Y2
ITn6A6dKl0dbfW9q4pp1aapOKJhPWfCuDD0IHzkeMhP6hmMcP6PFzXVz2GgPLYNa
LHQ3QjfYCNjxBnrl4Dpg/Cjk/1xfqAkzqK7sB6Cyx+YBNZSq/eho4i4z+5gRog4K
G2EAvFiwg5I04i15lfe5N7khTm/2nKuADKognC/pVCF0sfkmgylRSFFWjyGGXP7r
rxaUoK97xBs08aUAvgeSvu1xJWfAQka/X5iOL2ZPP08TYCtoH6EOTjefNicsHV3Q
qqaPuZvYDOUX57vmyA52uGK7I8tt4hkgV51ZS0gxwaW6nq+VYF5wNdCP/YdZ0Hvx
hpTVWT4C/OydM00CS06S+9MYZilkf9eDgLnoqFBMRgdB+1Xxs4DYfFS5Qk+jykkd
5BjXexB+v/uPTQ8wj5kPGIVk/VLjuAh4AP/hJa+T2OiHNOKs0CYxy4wzA1WKz1a8
XQAuV2CSQPKjsN4319Z0Z1TQVRXIKD9NbCHodSKf+FgHqG41jwOJ+4iUTb3/EWRs
BZL8XlRsUOB+t/CdW6hWJ4OUy+1VogHO+kj2WTRD2v7Ch02W5zvbWMHq9MJS2Ijh
E4G+qTQviVAMzKqi7yafayJJ639Gl8/cRGpS6bxT+BwysYPaoKJN3Uy3mHmrO6k6
C39sZygkpC/FFxLvjq2+XRirTaoUoM8MqEmC2SmEIjtiBJUVvnPX0xcACSzxcA6K
iRQZP1DcLOIbF78P4oKkbf1uP4/By/AIip1/eLWW8iM7hO28x1/7GuZNHsnvAdwZ
vy1AHmtjOOmDUGckesz0prEwt0hjHqY5Sj6idDpXzzH9vFVmTueMwiWR/ooxGdBL
FFBwjSwWW2BBZ7oO6+yvxEOX/16N0N3GT6uiu57q693JDzfmRJPaKwHlrSXs2S9J
6H9JXTyaBlhrtMhfGY2tPolnkPMEZ5gkZxmwqgmG43YfZRsEM3w8zimvXD5YS6xY
RONQ0FVqNCtiaJ+t/oHAQf2WZqDchiHZiOgkfhUI7uvWkifQP+LFCgIM9xAmYfvh
fmiZSgaWya66wS+e40Tw24dLPnGLV2jg/Usme2hJNchkQp+WypbzqJcBI2ceSOc8
wDMcRNQXx5fKARsmsYzj+b4irNZbbmxt9lPmigh63a7+3IEhRtuzIoSpSWLqxXtN
X1bogyoD9Acg5TCX9mbk1wni0/hLLTMWCHZ5clrub+IjDwL2gsZgjsl6WD55cf8n
B0vhBAoxM4Z7ciQ45s8vmMP5Qrn7POvebqzPnyjmnTXrc1RJkHJEXFhO/Vdnepho
0wWlwSg1jtj5p2xgVtVAp5yKrDv3v++m5KC7w5LHqMRx8sMLzrqZfhALlUtvnAp6
x72ixMKH9WVwUZKqsW/rIbAP9XTX6FWgWfbq3iWQmt51oAGjd2DRh+cnUQjH9d5q
OTaSMs4n3j2ACLB+XndIk27j/qyBuF32PwSWKRaDkPuJOoEcmmOJOl9lVgCSsrRc
lAtZgx7dKeRI4JzDCJeSYyBu8CbBLq1zKorktyYcTGXplwdZTflMEttJ+iwReOb2
nVy1ecG8PYt8yDjUgsgYjT46VZOO1edHGPGxOZbFNySY9FHTxGfs0dl++vPN0ZvA
fmLUEx8ssG0hVSl+SDDudpOihoz0d7rJ3AyDNNmkJD0IkYCMxp1iM550nJgNEWdT
XEKsLjnaNpwYgDo2rkRnJKZGCxkv4p6m6Dm3Wq6R3eACjtDzB/ezZCBaRMC2OGQV
XREbXLP86A+0vbrhz+/LvRRdySTnQvy5EMfLy0oghHQzyoakys/PoutQfl+nWevF
pJCie043zFqDXvuySWYt/G1QktddbVYm/mhntfKjMvSEhYHFNG6VbHjfFJL2g4hK
H2hKudN/xEX3Ph+PNcJPInIjoHJbN+krFIV1t50pwg2EUYXVR3/8ztukPWgI3RW2
M67fRtpQp4cg8lTSfmNMw7+5GKHz4dcNkEJoCVxGH7ZT3fI61/D3tlDmnogvHedL
g+S1ChuTl54i4ufqkEHFFkxbfkNoJYg3ByRxHWVAkM0nNBCMvIcEj3+ajATZ/gpE
JUv/8JCLOHcPVwIkFH97glGy6EykXV6hgPnO1Nb0O8IdUMUr7eRnIwQCsFRtOlNz
CMhXQeoWxMDlk/UuyotC7CCF7vWy44R92EA+iDGRn6UNfdGxYS4jPPTO7r8q7iyu
Odb0PJnTVAo9UG2wDd7KHbTPRFmvpSmgAaAc09P+L8gf4xPYnjAWVSOzbovKs98C
fd8kmPqtUZwGpbLqlPrCNLqENcIV4wx/1nU/lRyL3W/5pjEQTGTGafIRWvflG7JC
vP0Am5SU3BkgS+1KuoEkDb7srblBy6vwI16Hq2x+liF6AthFL7ASZIUaSthvG8ns
v1ZXFDIeBy3QkonP2C8io++V41XlC+rfLTqRJOC73uGYP3MKpVYvYWU/2/0Yvomd
Vqh7qu0a5E/Ot8nBRfZGIGq96UaXFV2+RQL7OeuYP+meUa/DlWJaPlxkXFWPRrgW
iKfZ0lw0XHaDrxQBobTI++QtHTZbTOePzixc/Vv7QvNtIAcf1qo2gPbUcCgI3htu
YyrY+c4JrRc3411DPo+d+Iz5JrCq/3D/734NoxsgOjimxS25pcMJs5Lw31CF9GAv
XXGU7BWPt967HZBrjubgDgYkiVUZwd3ct9qKAxCGbGHpcNBrjVfmQR23tXfTAMrT
5iKFtZsLSuu+8ZBsUFETrRv0o58bV05ys64naEqDrDtlH4VuLtnp4sgVozj9PFvU
uV35G69lrWdGfM0WvutzktPpZPsTfEirNvOsywnsWOtaEbR5sMfRe11JgDhYlgkh
Hz3p/kHMMPnn376u66mCczm+xg8vxph+rGjnWlYoCZSTUafuRe+zThMgroZB6Kcz
iHyyfHZcO0+GVtRIDrk0JUehqYoBf5YYtBBLq79O3j/WKTrc4L9/HCPn45+8I+O3
jQaHirygR22FOO7Ryuuwsd17mcSXw4axT8DsIvdqhbyS+zPhXTDmEhUn4epswi5u
RbmTgCHpDIhm7ga7+yF3s0QEkUGOmfmNpRoSvZasku6HlOLsDRU5wxJIMK9YujNS
vg89gB9HiMYhXc6S0UQdR2csFvxgsRWQwH3zbVh/fXcokWEyDFbDcHDSsO2ob3qZ
o+OsG/y0RY4TSTHqBtO5rmTwmvSG7SSsxHhm59FgFFeGvFzPygIPOBvl14TZxhjx
YCOrr5GiWrl9vaAChnckrZtHDIRDV1SfUCbx+exTqvpdZeKTnLsfJlaRpYaVhyQh
St9jNqb+Y7EQG11F/I0kei8tSXc40rdyf/s5xkuvL26LrBzEwWUtQHw+PUbIAikR
3cIt49wtDXuEI2KxT9S61Jhd7eNbgJZ3DGXc9EBFLgsOj3BghozGV5VeTHNEG9wr
inLm2tD38AXYQtBq5aaCZbut7hkG9RXXN6BWDbPfmbx5sUrINb6hwslXLCFusfcV
oRRpEp3tBMzdp4hqJ7ahkuHufSFUheXD3j7RAQJ2pUmfzcNUQpPQ1aUy0QumEe5k
i+oh9QnHo+T74ZweDMEFywL+c5hn+SvWiSyIr1TWgynXhiZDr2EEiC8+4B0j+DYp
bMga4Qs8QrXWDW3Kf+VmGBtIuW7yCepmrLEWSzEO6Aer96LBwQbb4Xq3fLnxm40H
UpiK5wqPg+czal6rXK3IhCF3AAv3SbJhQJlYUZNAtaQhe3RNSsqOWviySDWtXr+s
TsyzQBj28oHv9rOhMgT5kNLr71SceQhqAlKNC5WAitEsy0k1c0vdOkBGDSFde83F
vFPvElKFZqZmhJz+2OJwKTsqh7F02rg86GuNvbd4lnZ0ZWiEVUSp/E3wDPDKclJy
vQMAMwmDxWoXe47kEloSiGUKZ7cx9/hgs4TLUajytdvbddcbtbgLjmmaHaCLJX4C
2p23bSRce4HV1lbqzDDO9ZKCjsLKLhjgsn/ZpSGHPjZiY6uRn3N4jQ+ctAGfxkYM
FXjP6GITGAJTdRLaVD8NuvRtzRsTh8pXNB4r+n5gwvpNXXwJBv2DbVkf0XlFgARc
E6Yv8vH5g88j8pCYDVmirHUjxz/D2nbsv+mbJzNX12gC3QmWDwHNxNKltfA4npGT
npMkvVJrjCdHP1D2RmoXruSQI6QTV8MfQM+3jZHBEVe4h2GMVdH8mPWpKX0IRCgl
zfXZa66p3KfNctoRDwfdwrku8ZGmZe+Om/NQsiR991cSM8ebtsH4wHPGoud4Sm51
tVpXMyzvD2CBFiUbdHwihwiMhXMJjSIUSWxoUj7ZcsUBjtvDxTNCxgs54Hu2LetW
NQS8KE0k1Y5IPTG4Ru6XrXf0VrCdp6rKr2ax8knR6O4a2sz2EBegqnFfFOVGPeMg
7rf9vnXvQcR2OdLJgxgA5W3AKRoTJp1K7Wuz8GavPVZPYhIF1iUQ/bkygAxOyEkE
b+K5nh7IdJKZ+0RBd02MaQiqJFC5XIPnudX1sH9/OY+nAS06zyNqdDaHDiG9QOOi
AKvcfQ8izmBCFnsyOWi7KkuwpPp+t1hvkeDblfKDqTczhP61SnVpn4GYiuPA3rZj
4Axv/H+PPYjmyGK1yMHc11Ugye09n39mjZTxLYhc+59lZ8ct3s7iuaEHxZeclFor
N6AlPASTlRreXGs2Po4hSChvvhe43OyWRSm2rQiscG67GAiHqI6zP18R1V56mzuC
SgpKCOz70xXUc26fZGPzsNV+An4ZwQ1SWncOKQmq/g+jJq1WM/K118eK0OJaLcqr
23SAl8WhQV+ZK5Tb0FSeCrZ9KSCkevChjHfmMwLhA+x4ZN75RaK+Wr/ZXXB63tR7
8FawL53NT/aiqSbdY+xu+4uPizUu+a7Gs2TbOFqt73gL8zz2h63gTz3WheOn3P7l
U9nlUNhRbr/tSvYp5MjNxxOnHRAPsGGkDVBEytyqQPiaFyeIpyEHsEQGATxN7fJx
NZyQLmIDEzcfrjbhD3N/+ietc0pIdbZwfvofwf37uwx0XreCCJR0FZ+oDr65huzJ
C8e2+4QoM9DMNY2fJdZ5nTK2AkwmRGj7agHgdmFk0Y4XNCU3A3WuB8eb9Uy+JmO8
4jfQsXNvQ8J43sX4UF6PweLaI+iCiWKZlMTGye3xQiG5Ef2Ph4TK2tYytg00+cbh
gv+tNEU/azZAcJLI6Pv+xZT4eEP/mnkZR9iro5B2BNkndOk9EnQ64SkKhhaK9opN
SDHqiTKDNtBnFXMj8yTidwruHePRJOO0u0L8y3wp2dQPGst2ZvxrdK+UdY0U+Zxk
Wfvic8GeAweROuA0iRx4XUPU58xGNwf0kMXPyvFJ/kKIIehkvN88FtzXRKAOA+zg
w1UKRybMWHBWPCt6UOU1Pv/WNXOtIyBTSxb3av38d7EhVK8bw+XhVDf1ZKXapu/C
xwqwfeltl3146qV7L8xyOotRBzNjmaombrPt5nar8PIyE9fsEcBcHed4BXqYGWyE
MOR8jfawEW1Xu7LdnWNS9kf17bHPsZxSiM79SxU2UZa3AtRpfmHWVubGU7gTh2aX
+z5ZpBXkcPQd1ptbDmo8HuEsAedyeMJ45iPM5mZkVFOHDPFbTu+pWy6r9YbWeM0u
BsphYP+SU96SFLKnjJOaiVl0xnc59otdk4kV/Yec/PsnJa73VZrVbHGY1cTjjTOC
nyYvghYUo4sBQZfKFPZfWt15G/leGevTlYzHLYSlD+NKZDHKXr2MrR3Pgfyp7w5I
dV6Dn6nkhUV0S2zcMerMpp6lx5mvVmFnTpAsO4TsPX/dsmRrPWo3jcUA9gcQhDfC
RULK6Etgcn4oc1nK3oevKDCuf2fIE0FtZXqPS/ysVej05MudHqHSUT0MCZjZKjSi
WRgV5sMfqGwJS5OXbnwKe4QdrmXjRRb3xZEOeEDdix3Ka/qNJr6/oZmBJvSyiw3i
At4DTAQ2Mmz6h4kmekbOPI7mUtEvhpsOqjtcgKgu5ztKj2HL/9b2aYp4XDgTteSu
2SsPneh0c52j4ZG7CcLwB0tRxI2IjDIq0nsOpcZ9Xx+Vu6aUg81y871VDmxOSIpe
7USJRrenh51cmxqUJ8g+w4HKm5RMKEpUjOIYC7Gr5Arlk5HwASZec9o0vCgUfTFH
U7B2KkbHPhZiYO6dsnjkCbqm8ODCfRuquGE1NR8A9c7RnJ05ek/NQjZL6xEkMPDd
Dz65QSJy0cxQu/I0E+RBFUa+STZ8QiG0PC/gwIASiri9/BJuNnXdYpDFemH2KuN9
Fk6aE9V6cf9nJVWZ8gjh6TMeHHnDG7ul5SlWd0wmxY3+LAeBV5kImhBE9hvF3cbd
4arprDnV8uto6XBfVL2Tm5hl55WD71pNAaGM4cAvOSoViQzsv5UUikZ36G78SxpT
Tz0ykuvBe1LsQDrD0FIxtX9zDoww+PlrfEPpvtg1HzvxYqL5Mq18OPi2axDBd1FN
p+2CMbM6YltPiEEsSWVodV2eQ66wsb7q6jYBhFCoTtPvn86VakrkL5tZ37NEkRUC
agJN+VvSUq/2VPAKJqG0i00Z7U78tWy1/7DFvR6/ySzcaLHYBzRwaFal/DD6sXnH
job0UqI5dQbmzUhx2aBbf87mfvQRH++SseZUkistSb5HXBZUY+bwaKrq8QpGyh0r
8Fqoy7i/BXuu072QTjIdbHp7/RL6sK4wtoiGdsMYQ+s+SCOnWDGa5rrR7lty9eG+
EoyKRLSKUC9fPnzb423vGzsGsXhuQS1Pq09dyH0rEit+Z+IRVhMqzjXpU/vn5vMg
r7r0Jmnn2W2jIgz/l9anuKko8kucZghoaq4q95fnMNxs/GC3g6Ngv5kliTArKMB8
c865PR85wZSzBQW89LsLvSzeCWubxJYTrO31znDnM0y9R052vy1egFFG+eEchR2k
GFYWETCxuljjTFYFIcOaCxEiEIk/WVNiO5ajTiChUT4kvj5rOqeKThrJs4weU5e8
dWTatDDljpEoQSJATMLbJDZZm2v8afwSBbIgWMWv7IkSMjdOO56vt3g10K6moclj
uox5iMcjakFiGqbbClMDTVn48uoeLpMmHYaI9+s8CDlSoOmQhAbRUxCQVCpyAkFH
q//tHvBm4v3csmDJV+9+kmS+U4aHAXIehysGZIzO4Rs3dsQxmfx+fONmZikPMJFv
VGkgBn+osflO0Jux/X3HGxFnkeTT+X9gfeEKqqb8coinUVnZYLcCJztoy0hJqrtP
HDlraU6rqEqbAicqNRU/CgXlZbttvtTMY25LQK2AW1pj9mN8lmyoZBHnMr8o9jXl
qIIpctBAemXgY2Q8yV34mVWaWLuFd2KJlnF1XpPwEUiby1/BudYsKqepThwr+P7t
250rJsa/oI3WO0kK/5mL20AxfSn2nIaCM8CozSWePmyEmzg1WEBli8bj2biLKaB2
+PAgZUg5LzXDBRccDDeP/4FYgyCsqZZW2kpfT+RnyTzYrXOAR29rkBgu82dnHJ7H
J+gsfIDwOVAB5G5QKTo2cHzZMcC0R24g4kZyuPNvs+GFuKH2MVSLcCWjQ2XQlTtU
pV26i2EdFEMO8b3UPv33J4V970mGisU5jVD4MSUE28DHNC8Iz7HlwdO8DeqTyPFx
rcmdZ/gydoCgFppmslXiBTYVm5ISm9IV5Pja/wPxDeQRAwl/MDaufIufkvbihHVa
rnQnfLkIpNuPkkjiTMAELMnNpSTryJd28J/oxnX7K8r6/XGJkn3K+LZeYdycWvat
krL5MEVLjBaqGayfp1rk6+Jsnf2gewoNgcyeWpGZDADauq8py0/ISmWW175bv2hv
iZ28N2NvJm0DSZqiLHIsE6vYwOHEg030MbOUdjhvrLpa+rybA4vyXmMl5hjzPVfo
xP7B65LRwFx+LDvksaBxHILSSUZQRugkDCBj3OMZzmYH+xdNukHvFx2HkIUxxX0L
2iAgt+zjT42h+DmR/At6CKPOb3JXzfYqcMdALJv3KkKnYr0s+aa027oTXI9vwoyT
phGatXOALKYP2KcvhTUrT14ikIr6gLf/fDUOmvug+onBtYs8nOZ272PczqlLJuL6
H38A0GGHhaeGxzwXlPOraQAxvTkDlSVFO9laZPUT7L/Brd6pRgYjqKLmZSr38+8+
zXbDZQKH+r+4rjtSGxbm+vG57fmpVLRqgDeRX+f0JnCZHnMosYzH7m9WCfxhGJjo
iTET7Tm6o3U6njiTJnDzihewd8LQZiIjEiiL7t3NbLbLolvEiErgHAP+tK3og536
rhnYhac9DDGQM5vvPh9LDiGxJI5tqdd3RKdSJSRB1ZciCDoZCkGyIrfRJoBQYxLt
A4ZTG6uAfIuNiBo4yIiuxmBuvPc+4Ynj7TvS79ZYbbKYh5l3ST1Hqu2QM9o5Njqp
XaQYMEEuqh/c9ypbKkX4yOR34h50FLhbmx3i2ZDLJB5k3rnctrzATjvj/YsXq2LQ
mzpX4RYFksNgxLfvj4gj4UDNHBkh1kCoLkTQehCzIgIEDH+Iv/kquHTX9o50vH7L
EFhe5T8N+u7AbXfCGLxN7bE8FcVf1GNeW2/EriE2JUQ5SJ5CM0uW03jjZdq3MN6Y
C2vbBBT+AyQXktNAG/4vclNzV8tgpj0OBiHL3RZV4UYI8QQfC6sSsuuMVuhQxoV0
VGFXNKabvzWRJ70sk2s+TCvB2UestekEyO8NyWvzhL/YVgpSTGsZODH67KTHGhbz
aUJ1jr/eSnkRFtErxsmLqjJbpm74yn8mwOgMCB0o5hsc0CGm252eLy1+opD+QuDK
53/rWQIGE35WQDreh8LXj6NfetAKF1uuPeQpWNY8gjhN2Pgj0QPxaoia18MClTPB
+gDiTY7Hq8WaYkAhdAnG0bSWiGNsKsQJ9zvH/PJ+5X5riHrqFrpRuSv4hxwZH4yO
Iea+KBitHisqWe5fHqJe4u0X+kmdDfliAOhcnIuYolOoqPRgJ8XnmhJDjr5C/xOz
+6Q7EI7F2g1ZJNlHCSNHO8LrKg8BbfGT//RTz3hJ7zz1AxEX24UzewYROktTK27B
BFlydQR772YDWDOHvV9GP8NGRxu5/8OsTYHVnjNg4vlL0iVoz8WDFz2ZbAjzpbE9
wtqQh9Fp59dQ92n4NeJWTmGCfTgeAmCe8dl/cIXB3P4JzTrBTuPFztXWz0htFZ1s
F6+efhXg+XG8CQmU6Uo32eXibWTihv8epC2X43tSHszkW/b/Sut4TC6Yf3bKCINe
W5PeRUZwnOfmtbj9aLFQ0SROxWPd6ZXh7QuJAJtarfKAtGhFB/oq0mkFNKddge8F
4eeJ8HWCOBzx6snaPXlHZg+PkpEK4/b6KclVY7bmPKQ975BH7C5AWlcbx3lfF9+c
VXXIaLPA7IQ86/+oCTiDl40wa1sSf5LnzibVyNJ70zluXqFixP+I5FO+VhAEF0XF
NhTgj/fqd99zV5OSK7Ra4+dbBLAh2DOhAJifj26QPOKgPZi7hLC9rDPjtH3d8pCo
kPO3Poj+O3a66vZqteri3+u5JJbfRwMDWQFJiLXlCnZkBZCjrXvF9kmlHKlk1+bR
ouY338DjsuOwt4jSemlgliy2rwSd21HiZUxBGAM7mRLMFOaLsqObNTN4qSOMdQYO
N6jrlL6qFUyfD6Z3D3xgQQWcWKsPAvbXHEW8lb5SWwtubyllXaU58IkiFrxMHJ2j
0yMCNRabX+Vyni53ayT+CcP+JH8+aSsp9oImJkoHSTmnarXsYafMS1xyGUPso5i6
9dXvWhxkwzjvDSOm81+O+2A2QYWCMioHCrjUjU0GSXlkzTORMN9cUIJAbxSI1hEh
SZ7ciSyKuD7Qq2DD7i8lhWrhHg+xivTVpddPUbR/EKFAJkoQc0p467sHcmIFWmhK
nr5hohynvLrlgk8NqTWyX9cCpL8gUstVw4XGgE2ljWCa6GH4LJSpntHvbzXuai0U
LDmMwTO55vxhLIAgTdi3hxc9KdKKVWanVOeKGHDWIrO10SpS+8rsjhr/WuPLlHRh
XoSQhhl4955M8oXbs5y/f+4mj7CeSuW/nLWx6nJaap8gH2G3YD2J3ow/640mbaM8
8y/1kMnIW0IOn8VqaLiHkE8n8Y0xrjKct7poXLfqM4VECvsDDr7zZP0pSSFIChVZ
/GCFHHoIUHnGnKZToQ8tS/wUFZfMHGINmHghjM17+FCx1FtdgzryrkJHHlVERRtw
evbbVzhOPAtuRXiPhVlBcqvAyQ+eBbyDOXis9GvovUuhlxnlBbJVHX5/aBIpfd2f
qRaKWgZm+5WbjcTOyE2q0QCCmTPnMH8fempKJ9C1fydcZEascV2+yzV5F87gQywD
qdCr86DVB6gGjJQJJN4ONuR5yUV8hPgYIyHjgdEvlLpfYsY9iGHPMDj1zk2YnpY5
ie/T3fDSG8DdovFmcWq4Q6ltEynnc5CU9EKRROJ6x4oy/vMpdhgJQ8yp1pNLlFDe
36D2KFacvwQNNEVxeFdfbFpwlDx75zl1zNadoFxzGLeeT7N8AKqA5ZnIxVm9XctF
dGY447GTKXZHzrtTt4+cMY786fkRa9f51cjZKXr2B86q1cAjgGeWXGtxYue3FPER
oA5U/1wVIE6yn3GMJyU3Xm1+skpoNfYbfAd4RZQ15yRolbEckA2TJ0DyPNua3owt
D6Rt3aK3ha0bqdiTxjIsatVgelO+i2nnqccb4XVUtl7kIx3fwQZ7GaBezVe1IYjo
0ZK2cD4AarJfFi5hYxGjHXQl09xD3CFUfKEZddjDDdnY1HSUtOp63uDzGzlH+hwg
2l+ld6cpYhvjmoKQ2dPo4U3ARhT+dKhyYSjW3TUXCFN6IAZKp5lAuOpXmlXAgoL1
Upl4+JAfBymK0TB6bSJGuiXKZ/QbqQjYDQQDsxQE/9nTN3Y1YwvwTU9g6q8GKSPh
YoLCN9nd+PE7BPFDzgwdbJ3wTkAdP1a5d/04CgcesID9K6udqKfqRG96bLIBZ+08
Y4fh/hYxWKpBPHr9PFY+zL9HWhf0j2rXyoya88WErN2cQktkCbnoao3gytfrPcf6
wTkhUJnObTV0DfnsbOkj3SAJweSDXVKRtifUViOhTtJPmWc05Da1OWdFeeyXBqxT
nNGhUo5YxY6DT1uPGmDxefY4ZJX8OlcKxt2pUPtUXUV/RyMmDjGMOSy72BVXQEI7
YN3DxaNmvQ/yq0ND2WOvT8aMpT95iV6bN+grAYNDhYGfWUHK2k6PgV0Ey6mcFBMA
+2TaX0jDv6bWf76V2MIFmKJtA4YBKXunLkS2A14lCjiKzJ5Ku2fc4rKLcvIeQBiJ
f5RXnhL9Uq96+t7ndA2LNZ0A6DHQlZYwW6YitOqEGR/mj/ELDvJrGLK/oUjuVO+N
fBF2tjWSybsoy82OYSgRG5+m1kIyqq+7QZwW+T5pn/7k8mU74D3MITuUBhiX+J2b
OASO9cWu96+NPmBExObgf1/oKN7M8KSRTRIKTHgqXJ8yaN4vLoGONOHkYwqNpvWU
w2asmUsSPpTGfxnkQPaQDINJNKWie9dLeuFauc2BTqjrhiSf3zG/U+hVJq+5QusO
RohLW+opoU25C3SPcFhet5OASZ9kPxeacmvJRk6bW/XOSJikyPmMnGFQBPuleAjz
fW8bjWjIcbNEgZRLwZSC3rEZmcl1LZbI0oEv6p0hKRtetXTM4Ym456bAc1pSQOKm
28SYQSAGPNOyrldQJgCfEHE7nv0xBjouCiCcFC/1Lu02uDrGkYbIWDNhlhgejQ53
3t5if5cM1FfmwmXe3TEjRBayAYsJ/JSC5G03SvFyI7GsuTzoX2c5c0rh1EIwEkcy
p6U9XXD1Lp8vdMQBQoGBEW8tDLCBcBajPCKHmmgpkaBqEB89j8+3HhFFCR855gNL
lZbrwYAkxSVVcP2ddcyBilB6ufkm9IUOd17iRIKkSQI+Ou+y9fNB54uODuafO2Ei
QPOHfVSZKsFIzt9t4dw3yU8GOY0g8QDAAfePJRWE2eZNc0m/gVxs6KvRPEWWUswb
SjkVoULfvbIzcxzAveQut70PC4ZFEFUAZYAU5ut5p5AS74/wJMkTwilCdnp+v3u4
3AL2uyZPBHYQcLhRu/zacxpylnnTUnKxj2eGW76cr9jiuH1RZ6NefXgQRD0NiPR/
G/veHxlHCQSCpV1aAe15L5za9abbX6CYXfZ0rxGqCqWa4slrJdqvPjSBy620J8p8
aWNhgF9rDOF1AxaUX3JMHP36/TEb0UNxJ5BYRj9j3RLIGy26yyQoRX23glKsrmay
SvedhD3Qhi03LpBJEJZeZ9jvJe5vPDZwVdVrl6kExPynLhdDNrCs8vMgymBd76xw
r/7CyulIE3f5AxKbQghcFGWoWtJun9wsgGlwdAh6dU1rs6+1pA57dFqav+PdSVV9
6+u3bd9FssHn0Hjtu6JdPQc8EpTs6Y4l3K+3jfwBXbzgoKWEIWsu1yNIeHhizmvY
bqECRRpuNsf8b5zAqkosZryTpoQ9OagHrQhjhxVAI6KgHvOGHdhvcPZzOpfaVA8M
QQkjsX+l5+rv6T6eDQUQn2BskT0sI+n7KrE9lE3BEkMircMg0iZ5JH1OP5Dtt9ec
Q8Oavx4m3g4+1bWrsRK/QZMPpNaf68u0T6huB9D6ICJ8+D+wMylHALz5MivRPesu
5uesCTL5KouXIx6eSCviwx+MRTY4L7Boe7/Og5D204nIJZXQbADZDzS7sD+YDMap
ao5pF4O8nBI8I0yKnp+Wwt4TrF2wqmIIS2fnY8fo53bA/oq34VdEjBpHT9ZbZLjQ
M3urbAASkHXwyEMEdR6SypF8Wx7WNKMRiW3H+GlMmGm/1H6/ZYb7mEzlsUhersPc
b+Ygrn11C3qHDX5vpXWVgE2Tik+PyXUZwrSzuCexMJ8w2K4tJ4a6Zxygg/QWv6fk
LPtq1AqMy6da36caxvHwDgdjCLxKTcbBeP7oJ2SxXWrKmaOGOzYQYVu67T/4rOxi
9igIHvIZSvsFPTDaNgr91C5rK/cUol24ChcSaZsx2rNd5t6pmatZ2RLHvP0gJ6tA
5wmQ/tYpvWDJS0UWzylkeuvuyX9ixrXIfzqtYvGgsgzcw6KJskrgaC6tl2FrTd39
z/RjtvxNSbT6VPag57wHIdFrvAoz6chWQlyHG4wNLIbnA/NoCpufpZ/fVdWhoAlS
09s1OuXhtRkn+NPKtOizN58/4yLhQc5Kam0cpF7IaQU5yVSTjtKcimod2PgP52hh
kuWXzwkmIa2IUBe4IxswWlijiqop/V0BozF2ir3xAxj7RZrf2/CL0dhdVhJJbBCO
iG+d0JsI1g0b1afbRWK2nuxCfa1OlxkiBBO0tt5GfyH1w/bkPedOF7fDqINW361v
vzi9DVVoQheu3T4hgLMLgyfAR3qA0CnsMz319nn4bsu8dmevgkOn+T5gi6EoggQj
2MfmQ11HsFcy16T7ihSzpn+XKI2Mnfy3FcWd10NLJiUsbwsLMYHKh7UNtVz7nH/0
JIVgHn99QJuYoG/JctLhLy+zsEa83mIZ5IRMj2sYlTVu05fRo04l6J+xSlV8KMn9
NpkVJ/WQxwdiEuoFaxaGCVMTrlYufEokJYCoHyYNfG+8bcEMphpMlX/osOHtrYPr
flKqKyGahaL9aiSC/R4e5SQM7s4HpfdX8cxxitsVfd6Gd1oJeVX+F+LGw4cvlmUT
UWtyuRbvouFZUbjq5NFVV8e+yUEbI/6DzQrC+FXIl7oatm6oLubvF2nzBL/9yXFP
wegQIo1m27H+PeTcxS/F/RHifRrdhDpHL6UyFaDoD+8vpa6SGcmT5dEZ4/Q15uFy
KMb0XrVNckwtb5tXy2eGGayNskx4Sr42yLAcY7TuESHX3MHjBViDtTUn2F++i2jw
LgvO4N3MKr0KZcN2NXTcCZSISB1PrJMh2APLAroWz0e8r6+uOqZGfLF/bIIwLZVY
MMmqP75hoxRVkMw8x/82KhNDadXU9gPn1lpf8ZRoYGRfCUSpToIhuDKn5sDyHZCq
A2DA8TWq+RUcUfw/TvNk5Tg6G3boHJagjHyBnhYYJviJevuHovp7Ou/LYE+dtgit
rya9Y5pMH4CzElZqGfy525IB0nR/imyWFgjNxCYw3xITxEkGu/nwjJ2gX05LdO0z
loD8+cGetO5RvZwbP654PJEQYeajzGIQmSJtqeH0VHZPEFP3lBMWpKBu6aXWdmwS
+LeK3Ui3C314v/jFIdVOahI6MxjTXDMo43Bu4GME+nLNwL7KrCnd8EiGEh+SoGZp
7oFDn5SiJ0GbTY1oKeFhr5axd9mGopAKLl+40tI/1lxoeDDtHxIgRnDQ7/66fX7N
t8f2iLzn6d7plLbFDt3zpktihQEoB2lBOWWOW9W7wWVUkOlgFEdthsAoG67KnxKU
RV+3Gy8J6paJ8hIQY42W2aP0X2c7o4hZvJFmdxkixu3+ILZTuBjabPaDkMm3pcuz
8RzzuZfBaDx1qugsjM9aOdrmqtkwLMRrUsBmEF+amUAVDNU4RvBitaZuTgnNMmGi
ZEn/hlDJkuMUbqczzR/9suxgz9xalbtrEvq0Xk8WGc3ct3FG5IGS28B1mlbxIuKX
LZWF0xEC/0LOSOVBFr+iEVNhvaTBlfgDxjnhGBW9v5vIJFcHd/2u8Vp4cCsl/5vW
oOLwIHcw3Oq25BMrH4gJ1DxzNodjNsgCkCZrVEv31FOzqrd9DzSRjTKi9mMiz98+
U8yGU3knw+YQOJbNDbBdEWuc41/enOMYHV9054LtBsyWecCLYnbUdHumPaW3esQC
15kWcTa+cnxsvkGNBbUR9CBXQHh5VCj7q3dlEBdb0J00eONHgMWl0ia6/VKD/jM1
HskRvPIrFOMSYTatxag0UrhKzHfjLMmT6luF/P2Vk6MyxJbQd91T4goPrqakSb8u
tbh2G2HwsuuwSCo8tGi9ANZTJH86P7jESPdb+j+bEsWUA31QUTFL1/wf7AlqNYa6
fuei8915biS64Q1fyBI2rOSCHXi/eO59mmwH5UixWctUcq3NnLvhqjiYwcyeRp12
rQ+UrbmsNlNNiVDja1uy3tGxLUcL2X/T4Y2JK2IjloReJfvYJjX/L4AgZJ7yxJ2t
AhnN8aBA1gbv7NN3JnyVue6BYOVuOO1DcbMaB4DPiMqFDG+1urfVKNMF36Or3Q8K
I9Rhvs4e9owbQPWYNlZpU1U1AA75bR9MaPdpMUUToT0Hm0j+mq2TW2wCjIMF/hf6
c2TK1i8XpiyWaBAO+KY7KtekA2pBPIyGmKemtetTiF6vB4CcmxEfFkYeKvnzu0FW
mX5pZnyD+DwbRNqGmiAcPmEv5EcC41iQEVnZDm6NYXl++hfKYw4SWrzO5SEKwQQu
AEJaSIvJabBA0z5Be6DHvK91c75xxLfLGFIXYbc24+RMfeJYXU2VuO6sCkcDTKOv
eqpL1OX2BL/EWfTvYWIRbLFkqgVpRIxhKgf3xDeAVEtmXSvOBPcWzX+r7RDj8n0J
BbB5IfK6ZuRhxiAMdcpgjIG5MeWWWGRwMO2XbkyyAfGk/aG2cnHwfZoiWD5AbLLK
FYpmlIoGw8b77CIaAgfVEaJeXC6fMMW5BligNshAevewtBxTqN+9N8Zkt1AmoZgc
XxdVzFfdakJMGbEAYFmb4X3OI1k7kSnPxQlA5M0zt9fdpk+k5kXjx2RGTwjaLzxr
lfA13Ih+1ftNtkPjH8h4mxeo1AFH3noN8JRj/cTb7aq5FI+Q2OFh8U9B4Z6APLva
Z8MEqqo7UrCyq/0MhaQVHJry1O12MRvQdkJKGaHGnM0O/heIoTvMZ+N5XolJPqoc
0tpGHdl7kGOj5c8PnNfU2xI/s1hFjxXMokPaUIJPsk/1RG4q34exGMiEhH8qN/5W
EgDWr86PwNsl6SA1oYfmJe7Fp4JivQyADFPe7O+cSyWlbO5OsgkrTMcfzOZbiD+L
0y8rqCdpWJ4pQOshDktT4Q8epJOVYdd0pjH8tlM24WjknApkm42nlKoChAnCwIFH
+zKREMYAYUS5wf5bQ/MtTzy/zAkHEcUNB++S4G064lFXSFMAhC2Luo/tPETsVYt5
Gd5m4jC4tzVAso48lZXDbRv23fKRgWu/vaOhIQ1I5GXfCgIJ6Ymf90mSflA+deJ0
yQ6/JXojXO/rc7UjAWC1NFVtgz4j1gY4WYCyAXjXg/jP5HZ+FyvqCfxEwsV7a3mV
dUX7/N6FOZKHrthOx2RhclkKkohrkGxufrTMvRpcZOvX4wBED8lTZVjX8bx6MhA4
7znsYVCoqhXz/O4xMHVwTjGTlbcYCSEW5tO3THpvv9rGhU5j8DDBpgUQwnfcHZlo
D3/EPOH3zjIwkFGXLlA4TL6X+x1YNf40/QbABnbGrL2cWhE0jdCNjZMwDB76SrqO
yDqHmxS1irK0zDtXaraYipNC2WbL1GgXXln7k4leIhngkt2DETkhFspAE1VuG6o1
R2P3em1OJxayimF6dxMG5WeokizgE0ttwiKjgw0LeqQlmuI3dGDvL5Ka1rzgQHgb
LcvhYSMfIeTCSW4a51ziFccZ5VVW4Z6NxXXyHU3a/syGqSw25klU0i+Ps4KX5XnV
abygJmdLosiX8pTcN0xGJR9r5OGqGusAQ8XpUaTzSfAiwrkCe5ycjEDFQOawJ0Qs
3h8WadoI4XzNgkI0/yCji0iu/c+UlyHxvyuK826s0dUpGTSMMsUpcZHBHk7tUvoe
eKhRVxE9rkxuRfwNO0F+yp9ZuG475DCS+YYbD0nafD22LaMYGxK/P2WTMAht6F6X
JLmAnQ8FE2VqCVyRVThfPdJjttRRwr3iwBEQMoMKN/r1IcACcRygJ6H+fqZVNlj5
aDHuyFPYNJYoK4pgHxKsKPLi811DhCxIQLy/ht56uXasKT3RR3FmNqEQeTkVqYY4
NS+AKZ51amabEoUWYaz0RTrcdTbB93VgBtnP8O9TMbAyNfvjY6euNxpAbCqFiI7M
OzKlHQt5rfLowTdoCgCixyZIjBlFesJR72ca0SDhANoQfHWb86EZlRbBUCtuQxys
ciSJNchJR2ebyGkPk/Hv4iASf6e8dO6e6p69N3QS4+Ok7fpJfi219I6JVLPK90Cr
XKGiHzrlrr8+HT5I8zlK8L1M2Td9XUiWB5i+E2bT/L5g9KZrQZTQwaKjWLMpLBnf
fMakUREc4zl9VP6TeLaC5Qvwe2yIU4Z6M+Mucui8f2ampGMIBNG3QFkfIjo+V6xa
ZE1mOlWv1A2tjZeynJmOWMiqT0Z7EwwxCEk3igSK+yL0wpXQvigpwjHsWkzVcrTU
R9p1MYxSpxXSqZNCht6hnULJlm/uvfsq0BiAVWzN3LMrm/O/40+2DHxnwrWzrA+W
6TffxidxH/OZ0FvKg1b52KxSEQ6Ryy377ZsRNwirSgI06V63Z7P0EVpxh1KYxGio
E6vWeMVbBbNrSItcft9Enta2p3C3z2mubIqmweYzIjwWRw6WuA0omt9ZrerQgJQ6
JinY27b6S2to6YPLz7ex3TEm3Dm0zYE6UjGhjPjU6dvvZzttMOPBsnfhd+N5r8kG
muqgZnhJVhLHiNGeYdT9kfke3eh8PJlsdoNTX8eY9+Nyi0x4Yh5r6+C7tjJnXFGr
9KE+cWIJZjq9eL0j81z+142W617KFRTnq02OBPFr2NKqa7Ltc7dh2084PJYgApkv
Gj1Sk2Olaz8MT0aWlX1UtR0K/hocqtNv6YIVd3lgMm9tPP47EbOCPObwpM5PvFfB
JQ0mmazv/8IML/UO9gvY26juOTs8aPAi1+UNlBU9irdFlBF+nzb08FKzlcl2VJQr
uk3965uFTytghkz0sNcGzWusGWFZ57pdwteWXHbH/C9S3syfBbwJevtVSZlFa9zY
ulhX/PHbi22axTbSnJ4RdilsvzUg750ey2fNbWSYBOB0kVm3YriuaT8nyQoATi78
C683QRkPmnriByZ9cyucAbQytdWeSQw+4c73awwFNJ+pqNl06GHXJsYcop51nkxv
72KQZ5yqfWIfiIbGtPx6eZBVN5JRRM6GJO2jyRuUTB3hQEgM/9VFjy1dPabM6rMt
DDJKMLrW9Wi/KOWlj90Va7/zS/nFGUP86Vn4Vhwh+9GZ5DM3nqGBF3m+LyXSzFGG
9y9G8VsGDx+10xq4oGFXqht/U0jpbHHQVuSD4LEqAXZswxK9LyajyrpV6wjVnokQ
jkIOELBl6mNZfCADV42X8HvmY8UOBMjR+QjC9FGlDna2x2fpoKN4J1fQvHurcGtm
82RNDX+z1jpMjNA1YaNB1KVFiXv0YTjx70E5OJX1NGkEUlPskzHJpBnrCKwFvIch
d3H80Tj5mLc8JDiqB/8XMqkFj/uKpcqVz0k1gqLdQiTJB6N9dgyR//Roq+o8dkO1
ZOWxMvfukf45qKo3/lNGJwPM8iioPvKJ5VqxVWdb5Ab34IQHw70fylSFbQEhJiYm
ySawmtWGTdWAb/8hrcw9jVRl4bEZBXdQv+KEbdqOQYpRxh9GBIKXU0m7N8cnSgKz
MHkypDZGOFLirJkUiOwYl7XmKiNtFhxCeCgaFTU1iL0fZA7AAM++M68cRXMk4ALb
R6xsldr4roVSQStl3viyzil6IinUCnL80SX7PL6TQCibPOQaMs1AEa6rt1xlpF0m
POPFFoNuwfbnYK5Fue/h28sLO4SuzflQjGSRDN2ZqkhuGblLSX5i2ocXaGsTwmzW
dNFLJQkwWcejUgS6ikFQYuzwjJUaKoPiIQGIgxjvptZbjz/L+bIVN7HlY83K80kg
sIyoIBpNWcigeBdpUSgqdmhcPlJqKKLlmQQwDYj7SIeLnTRKdog7RuLI3HzcXOX5
Pso8R77CGjjgyIATFlBoVha9H7ExnVbuR0TnxmyJWzKuEDNKg1Wczqy6sp3FFdWJ
UfKJ4h0bXuERqZekJ/tCCvj1u7++rXtjuY/d/exZxs9OhH0mTZAQQMcxGL6qdbo/
cUSIC8HSycc5KitpgL2P2HYx5awMmlQOMfycP5lHV/I0640dT8OPPTTeRT5d0h+Z
1BbIFE+rMfyoLWH2mYBC03BtYiJaDpij3YNmkhxLADc8ByJVBknroLlZvcLn2f09
5IZl0FVjTO8Ohv/Ot6DUrvFdfZdMY2hDSkoPa1FYWY5VvRDCJsOwaEauYO9g56L0
/HpnhS3YrK0NN0Pa2t1SxaOXJqlR72HiiAP+Q84Yx89LUXn7BS53QKJFPBrhlxEm
x5+41yQCGSIg73gdhFLZiy4Pi6pMV7W/pnzvR/JMUiBUy4Izrr1zT+fSR5azwFED
7Oxrcp+WZ7VCsdB/f2DFuTvOBgF/sWLLqGz6vkLYe/OIryPZcqrq+njrg6UCYBhm
qvt7IqSXKaXxnyaNa8sY08Fv1zUehixVLwhR+I1+x5I8tPq1v3EDeFuFSwj4U1ou
NqdOZyaYwjl7dU0CNX1UL7W2KR2ZrH83XsHGN2h9PmNfj6bt43pvVcV4OJvrc9Rd
0sx7Pq+xSbvkz172Au7Zr8o+ZVDh0QHSBBUlTSYWQizTNt/+wZTVs8YN68q9TIdb
WhwVwdLNDaQl/8mfcqnpaF3VHjHqJXsXbulYCg/0Y7DpVvMZ0ujVLsNwVAE1fPi2
zn3fJ+NYEXWqn+GFwjyn4ZmwuLdlUNZZ/fg/wHMLPgcbayGTIaPFXODBTqlGs4hY
Vq3IzVex9PheR/BzngK9rmVilU/6Fvu3he5k/N4kkPKBAbijp02DIAJaSfBPZHY1
ju6SpG8oqJIwRk2QNozxR7U1+iQs46h7nWvblcpTCk3KrmuaFuXif0iNS5k7D/r7
wqN8QUJCtGnV+wCzNxyRN5a5ynyBpF141j4LCTO11H6S19ma87fj5XTYsN9GHCIr
khYksIK/uhFUZw0R3jTOgWVFHgBFaDMgF9n+RBti/vxXMxo6w8CcyOTFnO6a6GEk
UUEBSfvVEG0rLvWaqcDX0lfH9tp96etMUlgO354RnlbjmK2vVaUaTM43Fb0kq2ji
hW1tM1NbRveW2xQYnOXqLqaVpiFoyFqi/gz9Pg00hCousd/zSib6yVUt2yivZjmx
7abGhnfJ8fDW+MBiAR0xJyXDEO9WByvLq1GLs4rogjNomFHZGev9QVGhk/GpetNP
k51S9Xdn1YpRNsSFbmu9F2/ZCr48ONskcCkcoHZ4UbVL3bLVAiXR0YGZP6kzykN1
dGI5OlPCrxQg8+jSxzlRuV9acNXRyDUDCO5eT/EZn/PJvKIdcujxPOmLrAgDQkMi
2OjsHAEG/O9YKJkE+tbb71dOJnvDysSSy7cOagOV1Maor0JK2ifreSJM/iMw8kA/
cUIccG+jHQst53Ao9OKWTlq4+ywXFIAMFYMPz8VTIQD8AWkBh2o9UAR2I/rt4llf
mrCHMIDBeOG/3VypTTWjpQeJtqbvTon/fFxL7VAohPCDMHIQmA3yBRmDKOPMSxWd
IES4l32kLI4QgDzFOOXDeYz+Q89Kv/WoK5v3Ah7/ifGNv/3bLqo9f8WEo7QxKGON
vIw367tx2/Uo026IIKmH+nPcNAsW8IGrgtUf1dXvqF0vCqaF32F3E48BskxK4nLF
hRvvo6te7kjkg3Zb6bbCOPua+VP3u+pPfRxv6uPHgtsP4ZA9/wrdCa0n9sdSCOuF
fw38xSkyY9Q6YKAcN1AcN6aHYmeSTQPAm4hfQxQ4uBwJHjY9vGsha2jCMuQWhVAt
d/KWINqIuraq6IrvLvZVxNCzrxb6RbFzRxl325KtLYSVHFIG/5bw7kLA6xhdEY49
V1K/Idd/orCUvlvTWK82fgvcsXbD47e5pijRu4lhVt672LCThzeTDwQLW+kA+HmM
EK/LA9nmWwmA6r37u63Umb1rVsh3Fs/sNmbnQGLFQNWMETaTNA4FWTvCVxrWSnr4
BLvEqrV4is/F4YMB5eImVhIh5m3C8ghKode0XjY4LFA85iLBPIhEXoBtzopJyLa2
X3OTV0GPowJCmqAKRCMXIOSoOjnBkiXVB+JJtf8wBwnSve8kci2gGkumZG8RwBpZ
7MCb6sKtZ07WuL+YXN5tubqNg5Wte0obCnEHRcbbYkyt7CWXbQMA1XcBNanmp8QC
wThr3c42DXasB/LQYbg4zFfCqUiyQyIJxqI7Wzz8NG8DYDLtbF+AedfaBshDNsex
iLMB7X2bE2S80M3mBIm+K9asxiuc89oaXRpQV7ZdEnVewqpGzeLIfKdFWH6fyndO
KqW3pwCVYMjqa0i+c5+J+S8dsMT/KP8zbmoF4abkagcz+NWADOtSZoP+/V0ql25q
tnM/bUuZr70dqXzkreP9eHj7SL8MWoEgf6fZEgT5Xvyn/Oc4RB0XrfQ7VATpWgw4
sgBh2J6V19f4DYaHR29f4Z2ufyAw5OhNRpy9KLJqkXn/xiyO3tUFBN1gd3wx8l51
P6T57DYmB54prN6faosqDynCYCBK1xsqJ3B7wLgR7ttwWNYSo5tJpWclIZ9rmSLR
y2AbdmLBFkYVgkToNX3uTdO0dermsAE/C8FJNfxXxiZDbOSJwFpOwlXbEJOrk3Jw
Fk+p/Kihqe/z6pBAYhlXLuprax76qGHbWhjAelLcVAQArSH1QYzud9sDjO/pSSlZ
MLlTzPYKwV5iV46DBfYtxOTGVj+Adtn0RyeDPwNAT6wvLSnYXb6Sq6u2A2gTe41s
8mb48hRVQBgsjxmt3TCot7EuOj0E4pQw5Kz2GXgaT9dCgJPa79+ey/We8nunK1Qv
Zezfm4MnoLo+zqm4hmm1ox1tLFvc2lP/GvQu7/hq7PdXItQleItqyfnUH8LBrtkF
X/LhNKksezZFFmgxZ4LhgnFPQDuMExQMnFD0F1+TzvCnj+2g6I7WSo/iAyweExZO
aSvYI+FiJa2Dbx5Gc3EYWmiWC03ofgMheIdMq3wRNVPkQfXJbvwloqZHqHxNomqQ
/ctM76ZCqNIztJGkk70nJVdzuT8lNsBUjyuDr0v1Xtw1COoH816gHhCKCpAB+VQT
r/jqNSZ5qBdsU2VIMT+x4zGkWEYPm+yvtE351r057xWXVyuvkt+aFLUn5kVR4133
kdLcowEdk6qmKnpeBFZJPkY3Uw2eyqhP7SsAIp48xTdHuQUcYBFVU71A4DE0gn/c
qDhm3F0iNn3q5zanqZbnBDTsBPbaKSjE3Tx+GMHkIwxxtF0CnxE6Nn7ytMDqbJSC
CO15eBO/njmnecjGUbtvW/41MJTXKU7jx+enEAv9frVOYgBhHRZx04QOvtJl6rbl
zPJgRJiEmyFkopTIhuWZNA2yK5GMOxD2R5TgjNeCoBbjShH3QpfsFfHFtkzYM2ZR
4dq5sXHDh73To2kU7VASby0JlkPyEU9K4hadKjy0kiWcPvgD13oi0O71munjCSTr
K5VJXDeKMpbWhHtQuNnwkpvTg6pMyj6hCmYFKqsJEmSrTl+Xyw1ok2ebiLrhk0CD
8isKsE6s6YfP/7s/p2QkQg3x9qGsy1fcu5AQ6g4LYryjZTEXRR0KHngjD8ZMdJUn
zORGBaxfbBGwMq7vg+RHyUc+kncxbg1HMU8GWd3YBVnVXbQDW8ztTQIzRZu9thgH
lQG7+pT1hVmgrxCSsPUzZXVA+XiZwE9tFet8i3q2UvUpIQ/FNtZQnXAL10cObGrs
5nSfKGvNsc7USBsRfviYw8et7kNU5b5oXbZfxivHju49+MWb09jnN5aBy7oU7LNU
VOo0KgF2nPdfFL5qYnF/dZc83bE+PfsmWWCwaFPb3m2sM+pYCyDnHLZ8jTi0TxzP
0tsN1IqudCeW6G+yXKSzO3gJ5pu3UeVeb6ZC8wd9K6xCZ83xvgwZ1CorSmnP6DtR
rDdD4Rk8YysbFOotPLyMbMln3Iljre4f7rys/u5ny5SVsmRkI4AS+BBMtSOCqhM3
wB+xutFrUro9vFmNAUHAimFH+3SxD39V85CYy7RVnEb15Oz58IKLbxBOn9aktzzd
d62CQLMAEZqtSx31bAjRPGsr203yRvSau5FhxPocCUjEShJ1E3l4CY/c3PPdZQOw
1TL1sBaQyquZsqtUg0BwvJIgJMHbHi6eU3iVMl8qa039A8DQuxEzKR62etfibzFG
MPyBmkCRO8rF3iIlhMzBt6oiAp7VDk8aBpz87zFIYHvXuVsLXqC8Phr17PvkzzQO
bDTmqbO8om2HyCbMwVq+gX+pxjekmhTg1vMkuHapk67wNAmMtiSJWMXOtiEbey2A
ipXOVDY5X169SstiWIJzANrCDHt8KJH1B+MIH3QCuCJA6uY6iIuYiRoNIzch0doH
DHT9Z2mUHkJ1j+aSikS+wcFJeuWCV2U6++HA00qyU8ZDlA9cSI41bgguC9aSklEQ
3XYbcR7BmZeUId9A+50kk1H8btTbA6lNC90zIQMd3/GWPAIOFCXaRumxwlBymveX
Bj4sbvc2YrnIfPAm8rySBJmXtUhu0Pp/fxx6+NYDKgGKaaR8R/9++8tJavO4wy9b
Dr09h1xjTPkFcUZP6MZ9cUR3/OoUiSsGs6PHUUmLiIK7kSq4ezbTPwquq/7S7rbl
IxjlhxFXG/cEjne0zGJ8pN+xtXoLj7RcbOGLng+FvT3Xrcx7Y5/zlLzHwPkxttsK
Kl/HCSJ0gkCny6byPzNT3lZ3fPSuuiocc6P16k1InRdw4rBfjL+muju/Qqely11k
oVlXPaKRQpvVZC4YVR8b8c4IIi86yV02NXM1SRE4ykzN4g98fykL7QlcCxUT8fCC
ITEuPJtsENdOmtPYZu7JzQt9dvzfCLDJxc2jEps8cKlcOn0diXBAH1tixnhvLCps
kmSpdIQRvGDR9v3Ap1a/qdhjtPUxUCPnhD2gIjIhop8xkE8TP2qxzOMqJSirH0ah
/F6SiM9xwqoJskKNJwsVYT5VA750xve2E5WwOxmuBe3poGMD5ig+vE6Sbic6fG8I
5PjCoNUXrwh0p5uBdaihXgzOdn5qCyKQtgX/X8fUtOv3i0hTBjkC2lB/Mx7I4ETR
WUmG9Gn8fCnjMrl9igbeAfFvhuIK5pst5MBSuQuUo+rTvpZA2MY3Ytf0U7ktSUEl
fX5xwpFsEvF948B93WaxqSVY1VzUMs/7s4Y0lxrEhDlqvesdZhMinnY/Nw65OYEz
Nyulv4a3YkD9YFSALRM2wZxz5FS5Y9KRhlZo/gq1FH9ILS2CU5HtlySW36p2F6r3
3trUVhXXB9uGWneY1CSVypXba3tNKzIoS4RbhpzmFLxNOPfajOcPqfXq249aWcp8
GGC2464zfcjoFKqHywCj5dY8kzgs3em3LTWGtmztcRKvESsNl+KUaxfP5eFK1PPm
Ui9CJQv4X3JfhXXmH04/XLkEZK9iMBjQJFa9fVWcJjWlj/3VmMdK8esQRlmhZejK
w70zmAfNl0HeMAbXmjyvMBOR6eU+lR8Oq2iVHjHoWRSU9Ir1tjlcQ3jyWiqt/SfN
2Rq4uJlzupdX1H2z1KG8Gc1SUNBcBNmpBpdFSpvp1yVBA+X9IJQP5m1wimX87tV2
Z/5L34y75jJGxpciu6cIho0/D6sCMqRP+xwiHp58CXp9iLU6X4XreZ07iz36ZI3R
pp7WCI/VAYZ23B+qCPbdjytNoXUplGyp9HIcVcCDU0MLoDi4Kn9LUAuq7WXM6SFL
oF7zM+a2To3ITbBdq/SNywJaWepwEXeY3WbB3qvePHgdaL08BzAz8XoF6v4a9Fe7
ZsMHAfJWxP2QE6Dyg3jIoUR2hLAIByiX94PbtK9f/yPrm8EniH1HDQLpju4VGr2V
0uMY63U/zrLG6VWQ9fP6qAYP6XS9rr+BNbus6P3OHQDj4ig89fM3ueXioG6hyqtL
9QMz8FH/wMYQLxDL3j5uAz71L2LpXQ5YaXmRbSJUZNBFiZVaQM6lKOdh7rWnLC4i
wVood5oUh04TOUAj32T9qtldHwrfZhjWt8BYU4CWqKY4oRo3A+i677SafcITAlCM
3cy4Z4dzriRVVnSbgzc/LB2rwT+ILlCuGwsnF0/92lAq5XWmyBf/ZsMrJZAcVAuu
mKdqTZ9Fm9pTaELn2EGH24cK4gv5boPhewa/hhJw/rhMcfW2dPMrMk+pdq2HS2/n
gvrY0Y1ZxfskZEcLyZvWdvrpE0tAvNvaak7zxH7FmzqdmrP15nxRmcoO3hM65lA2
h2oGsRG2RdIym9fhdklq1g0mfB4pSrqurcs88pQfxDQa2IhWrMGKlHF/o4yPHCQj
NJiNa+4oLkebZowg9rTu/XTCu72G7ZTdpY14fK92MOc5v4cccpbpQtLldnJLXkFV
XmB50KEtAAUSyZE6GgC3JLOOXBabCCIwC25M3smhLnhCIOLVRgGmton1ROWqw2pp
3Fq+1F0MXPJhNUW1uK0w92Kk9m6dKYIbaSnTEvGv+CySsYh+rJauFa6tkmVXX8Gl
aRqGerdWSHoWJVSPo23CUyru4hxUWWzN6bOmHEwRGhOgE+HAKMzT3Sp/1YgfoBiG
xg8XWM6E2bD4MrAU6e6dquK9pmAoihvPzSj+5XYnTlXOMey/ENy5GXPpO0FEguc2
NlU18usWvLmp+B6YFMhiJT7yThOz/wRy8HmE/xkzuoaLwVyoNtZ/bYew5+HCLBJh
vYWncjbbXHSQPCi1PauYgO10ubFRJTPPQd9N+ova1uf1PshWVr6vvVh52ncFuhMS
B4vEhftkcpLZ6sBiyQTB6clhRtMf5oN/PRXdJdZFiwSHgQGuMN86RNO3oG9Dm+u9
9nKYKIdTnoI+N44HdJiGNb90R8P43fgEprPUCZQ1vzloQxSf4Kiau17bygoDgB7S
542Bkzo3pzAN5Qjhmcu04S9UOSRdQkeMjUeqh/POFSLtBA5jusXw1jaNrh6jyYZq
mjETIZexHwbGJzElTu7QzPsdyomPZaBz4gRn1+dTtwMXkPoJvruO5oBxa1OTVVyh
cJVz+TymqdQ5FKSPgRc3Ep7DBa9q9ZarKMg57n0kzRevRv14gN/mOE73PM0eG2dD
gV7zt7F0ZRN1/Q3gZTXXoQFYhl8c/qlPn3xu6FXsOpsKVB7oMhX/Dxy2AjsXXR8G
LerZU1DmBAVhzidrRql7+OnPlSk+wxNivGxkWRmhqSbxffwLi+YbZ1BX+4cq6Yuw
6ffaqH/vL3pstDEGf1Vb/TDVzXKGY0Y3PvIYg4x5UtHx1zffwYKBV4i4QCqpF6uj
SptwQDSMTFeextBuV5Wp5RpQWxouZf7pcSJC+Yz5qALDR9+FtH8AhW5A725Tkt/a
2/Z7UjsbJTJCX1Y7bagee7dKnaI2Oj8S2RtEPVfIJMOlHiOzZMGmrntG53jL5HVs
LrO07nZOzYzRTJfieevG8gRbI0bzt/SOwEcdtpjYSO4iYYRqB/X7tWzb2v8v8ToR
dRmp+g0OVG/+mexVn6x1ESKZqAulg5GPtiEd0MX03c6HhGGTsRpKD+/2QnGb+JHd
ezz8Y6rDUTK7VkKXuamhJJyMJi1pSSPPUO2/vIcibmCY3a+Z1NJrDt3q2ZTlqAwP
BVx/RjGJiC40JzyrT6hRvol6e0M3dvrPXoNImdeDh+ujY3qOryj6KUlhX/yR/x99
PpdpTroNxQ52hUeNTO0wYphwIEV1QI0G3X2qconLBcosT/lutx/Xr+3k/QfsN3Iy
ALZcQi7AwgHqpS4uQUqqbYk7AuHu5mOWlTxbbz4zAFutPkZIkWXonxWEQU8lJ+5p
6FczH6wCbbZSpGA0GPzVbSWzv+fgxLSCe+3e5rIZdC8mQcLl7qe54okYxzE4UqRu
Xm+tdD0fcq9L7whbT7gKu9iYtXkJ9Gx4fV5ic6t94pvnZpnHST4qPVr1Jy9O5D6J
YkJD/FPLlI0qKEwrlm3PPfcUPHWgZ+bxfhfmPEb8qhNLae9UhCdPCul5MFBw69sj
t76ITaD0otFyceLZ5ie6oiNU+XYAoOmHmhgSNtouNBaaQ8vkaacck1aO+vqNoHVe
FgEeiHhUQqeRcd4ThS/oVAYFu/qYMdwBMMlFVt8nvLWT1Trk9UHdSXRM+AyZGgCJ
/HyS9EkGtPUxaMHJ4OU3WWVj+MacbKUNTXv/b11P/JbdKp8uqn4rSwnqhb9f2RdZ
EZ9W9ImSMAukjn2TPpYdaHzOxeT1ipO0ac8uz/D6DVOqbfWUiekU2R0eW/v7d4qp
5XYCRpMuN1KZ1u/qvLwF+f4rGBzS7QqXAYFeESqhErFQGR8jDiyA+I09mWLlAjwY
/NZEyIBPkiILbElet1OD0NPdQXXj2UEwD0I79mdtMr37jBtpeIyIDQEFhkRAiSFJ
kgtulCATvQ+W7Zi27aGOxp/mHKt+bMULkQbQ+pHzQ+08YUM3gxWhGY/HcP9Ws8Ai
Lem9mm+ocr2zMlFjIxGn7iUGkv+A9OEteHOEXxYWV3IpSaz6pGy90r3JZHXxgjFk
RjOvww4yLEDYDy+/2m1quY314rKus5pvwqcq81XyCBFxAUmCCfZPtimVLUQ72FVR
dydQYQzNe7od/CEGgyBg6jBylSqbhi2kJYmp7Qo3edLZNbMYzB6vJMnidb1+CBLp
9fYo6GYgCuTgDSXoGh9o7hvrga+s39/Bn3lrMjyoOcT/lOMF0FscVNFVwcZK+dxZ
xlkQRJBmku2GfYC34COi7MiMoPJBo8v7NGe7H+opnYOZOctNM67nNoQL+LbqobCh
zZOIGQxXz+kb1pIHFYWVKZ2K0aNdVO1HIOxr799sLPa9TXnD6dmVS889sXkXRsp7
EIAijYNNj29pZIX5sQp4lAjyZlPNVGW8zjx+FvYxZboEItP7vJuR2uoXZwfz1f/G
M1qlS5yqCVxtBKN+DDWgZfrqYxA6FlekjjO6z+SEY0Sh6XFuqhKYwU1ENMcragSa
dZ7Uip7Y4l0PQisq8zGblVzD9Oc4MOTr7H4pkq3QsdhKgGbZUbnf710rmm22J9/r
U3a/rge/WT7HMvbGBOpOWNviqmfNb+/paORwsVuecUOxRs2Nf8gHV+u09l3iDSf3
lMjyQOd37VrO2NijcX2ZJR6ChN+SOjlAXJHC1Dvot1kc1zQWWJpnjuik8WWIjx10
HKGrjHW7vb73QfKXLeMkm1vQXeF+HXPrBuvFd/znOHhKu6INs0T4FACypyBXUgpp
LZI515mfwgb8AZ4mvUE8qW6XXQi05oRjpbu70MxrOAExIrOn+LENrFS9QCnQ+Bec
DbchfXmpK3SXFHvHkqYqLuT+mPPOPNgXQKqUxEbNhoSFxKWBm4dM7sMRZd2DDNcd
gmWhxnsOdvwHR4jxfICegbxBpJwwNTR3yQNz/OtVr/6Xek+8XPZq1DkJKknC2Jhy
f0Mq1hnUSCif5diWDt4W26cw5ab1zM0Dcz3KmG6qLGKPf21ZfHH5RWKSuiqHMd/n
vxx9omcT1ZFFNtUA7KtZ0J1rILA23lLIO+cynQVoROz3fkVhFH4tE65vHflA4FBm
BxGFfeeV+8RUkTWEvyn0Dvz51mSY4jItXJ2FUJhMxByDezgLs3M2gq4xCX3AK1M5
ai4tIgyDxgPLwDYI9slE+9EEDP+PtC/HJfy5mo4gd6feoBGA51UMjiZ6wbGeRsMx
AhrGrMU+cty0QsLPH3Ze9wLG3V9E8/YZYTuH7+3nqQVtsc8zjC1x4d+GS0sdXPAp
BP12myxz7q1ECejDwl7Lgx4flf8VDD/m0GJzul7Nm7CR/zzdxfEjBM5hGZ7R1VLd
FKiv02ek7T6aOFmhCXXZxD0eXb7VgiTKDpi5dA1WN97njg1HEM7uO7Qg7qAQF2l0
UV3xZ/D/CJHchq0jsC6PrSrbehgsMPCsSYRNaYsyQHyk63ENl9GiuZCiI1eO4tLs
y3SBGUtenjMaB+8DbP2pF+zxDZ4ESmtDfTzmILIIgGg7B/kAdFMRU8hmlH1mbhcw
FCD1v7ZpZ45NYBnIvvVCUiVp88/Mj9DuZsnzAa8F+f2IlPRUYsdDevfD1bp7Lrhb
p6hdlmC5Q5t6DN28Gh+yE4cgz86u2huLJXORIRi1DvkgsiEaXt+w1gdcnpVW3N4N
tc2oXBttcJ2GZgl3mbz5+wWXLq0fbQHFJBXokgncEg9w9XI+ewOVRMTIcamXdGHy
R2ETJpp3ekZaRAvZJZZl63ea1U514nti8oN9oPw8/bZ2tDPWxS5yB+7rdh4Qrcc/
AgSe9/EnXJMks9rHZhFFJVqdz/KJ1e3Nc7/ZMz1P3gFsiYGU46VzaLpxFi62PX64
mBGHMFoRkSza6/fAAHLRPNWESVOwo/n/Nqy2NlkNxwYn2c06h/z241wgtMC648g9
4STwoeIMM+hf1OW8MVtg+HlDO4EwW0tLOoa8wgWVbOugVGIEn6iGBgqwe4HVPUXo
nQnBxmWhsEPr7YeVelNVJZgoupFT/2d/rs/IWx6ifTAWw36sWtK5lEU9oQBzT6QS
quO/+gzf1Z+l/ABHsYJKUigdv4+0iPZ8AasyStCgMfyLmA4uwKxo6HuuB9Ouxw5U
rrnGo0GgAwwY8vRs4TH1s7M578zuwsNDuB0pKVXPJU+815A6CSMJgE5zq5UgzNLN
h093fm08chHlPudpaLdK7pQByQWDN7Ff1XYbxtZXVgtevf7DgnNmrJ4N+I7KR6R4
ltSvbUszoxY/GbAiKX3x+/leFo1B5OBdBbNuQh3RZhL9IbybkX2fLnk5ksRBSCtQ
IhzqmUto6pi8uicU/Q4vFBcy6EIwKUUPLp4ZqwtYF2M2ILCcDbHNGedXf388Fe3o
g6PS2OBzC2zeX/xIxlS+ll/ay1y9qqEWRt+Y4IFrPDcoJuFpYj9uGiw3dgPb9Gnj
14MAHz6pfpGYaFsQz8R+xnJLLKveEQtiBpTx0RYL6ZStB/aPE7KW7fmtIfnMSxKF
+uEjZ7zmIfMpBhYIyFlaBMlolvdwiq7toit7UZ0ZPuanNYNZXo5YGIQMk9PwLrp9
EaxJJvzuhBSwZ8tUKYzOaboBwt0WUU2jobBZp8N7XiwKpU3cpB44XCaJI7gP03C3
QGpHAOx2P+Tbdib30LUW70da4ml3GGCJpqW7h7SPdtzlBPqsRUk/2HntwQ5ca+u8
ywrFyd8kiSzsq9QWoceJT4/LEABhgou6T4Qgetn1+Qy7Lr+h+pyPeotnwqqYRqw1
0oDtHvkNspQzk5ZRHWjvknIWp3bTRrW3TRw1UaPlBGbZ/4aU8fui2iBIBmGUOyrI
k9q980+PF5qlTqJOGZA9Mv2dlOP5Sor7JkvJN+SlSzxTW3pcjbAyFnyJ9hOx9BHv
pXQYsZnOpCmlURvwgvnwNYEBKiprf448S3PIMNln6vERhkEQcDjhf5gW2LzV7yRY
nlu1ruaYdC/iu9XNCBGR5/G70kIdkGOvy9cUuKc0BF5ZwtipcrX+S2F2U8mdVRGp
CzJPeQ5HwoYj3duyg/rkmxPCREGd0YME8///RcqxP26HfJFzZpEtzCisZAmDI0sv
HWS/9zpabX2tIShCilJEyKLQ383PFWrT4vulYq7ZBn6BPkhXxlEn4eFoKHf5imlS
aKLfflTMNSOAzvPe6SaAB34CyNjSQbpU5q6dqSXGKliJJdq4XtN00S3X1Ha86YDq
H/Cnng561ZBacRpNFcROF+I9njsZsnYvUHsz4DzsMIcGoEuT1js0auIqJn6tSZ0J
2MnoqBNaj016aJ2LXICKTbxXuU9sI4m4+pvjosh0vHQqPnZrGKeKM/2LJwRYN/Iy
Nw6cFInRitmjSiXkooTacDTIFGewFwqCVyFItocpgLCcc6fl5r3zxSUFezyXI5Yw
9H+gSoGyeW9jaVP2VdDSGFU6kGWpsUddj4H2ZiesVSe63y0elOx+S7/sjhzbaRV8
pdygUyF36jlbSKHv7++yPxokS26uOOTOetIncdjZEzS2hC7TptbAl2GwjPSf2O83
0vo8dJVzVvTZxyhAn2E/gEwSiKrE+b9XLsCgB+M7N5hQUVd2nIyIoJOoGWHH4KSW
Endk28blNuXPLu9pmQ7j2EjPBJCu3+jHKW7JRzHf8EPq7xTkgV57Gy1aJh6sbDFa
tS3imdOVAOabAPQ3M3UL5Qz4Jc6bdS7LEhK4tP8pJZo42MhJRq/BH6tG2qW4EKF9
vd5EcwD/8W86VrSZg3/jaOgaJk8/OHN6yXZxYJQSuQ6iw89Z9k+/iLeXmhp5RaBu
dnWG3kSrbDpKTgwcldA6Ip9Dd5xkJf/sNjtNbVES9Vtm09pz64JLHSPu+uJlFBqq
zYlOdbbQ3O0oI5bK/64JjHuFcW2W4gpuKILOBWX5BZUD2SGD+prpJPpjIkhHBjHv
ozcwN9QXUIV5VBnlRQAmzbHjrXp6g/CU/uYrI45o+bIEs3v8HLO55ecL/t75sKDo
ziyqsZmMcxKtnwMEw1koP9krN8JZcohc4yaGgeCDO0986FI8PMdwyPVJ0DkmJmbv
5uPWX/vN1P/+hDQlZbbzfMC5GtqiUoGvCOVr2IvTlG2uKWtHkgaHKd8GnpHU9Xhs
qpGi38ZdQ5XcmC3QnmQxETYkjA9bcZ0YR40TVLnhk1wtdX93lqwUE1ljebhVKIhV
/xpZBoDBJXGEvq0XrO7QgFY8Y8uKzwhCW47/hJZNGSgkHifCTlrmJCHJwjmWbLJA
Ns8mAm4EVyZi9Q1L/rufh1X69aJu+frSjoc+TLNoqKQqO3540UfWemA1PfR8aros
Upz2WlV/p9HrvhuGUSLwNLPWS89/H/xc/SHrWQe1MSUmfNv8DjjATG2Mtcsjo3wh
uxL4Tj8EOoNbPUoGHj71CCKyFOlC5YS+cFcolI7QQE/3h8hFE7f61dvjENyEJNi7
a7jX+av7a7+4zqgR/1PYnvHuBlaTdqQKM+HB4DCQVec76kG+GvdN8TJJr81HZPQK
61oNtZkJ8lzJPOmo5VbpRRO5FN1qVZ3DiWQS894EDwyPKu38vzEWUnIzxqMkBpzA
DoLlvbtuujwyaUYRBVGSJbiXj65JAveYSkJYi1p7tSrEKTZRwHw+T8Jb/G2tgyaG
vaaO3hvHnyVbrzfab59J5pB5H2SVADFrlYki0x9JwnY/AONREhqOloD8iRLxuiT5
qyjz3aKUYhR2Ng077AeJhBBi0ZIgtcGtTr8neTquIgsCb5zGuNyGBtttx6X6P7qj
eXmRa/GAQm/cXtGLf2ey8J1O3DjAkUyIgt+P38EgYunGKkrxFPA3DcEcpo0xSfYi
WMNOgymCa0BSWYunO8caqnOXErFZEywPAli8NTuNe1P2Nkk8l4/3TOauYeA+NJk2
mSwDo6M+VkJap7qDiUU8Dwr0riqxUrqfUfr+pQqOZJqls9Jzfrxj3q56mgtLsqKE
rjOli9dpe4spV+5wEUZxVxeI0Ode1VWu+Zh/eF7JZiVY6eB+L9ekx6hLC69T37Qn
7RcRVi76DL4Pn1LzuYNt7YknSV6+EGYsX7Sn9031L5wqmUqYZQNwAlTE2UuRRHK8
T/hk+2Q+1hg2T0jyCuhD351T4+g46+UdcUdWT+ltrpE=
`protect END_PROTECTED
