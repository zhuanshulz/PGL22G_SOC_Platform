`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
22WnXC9M0M7H+dRBGdCLexZRr7RyhlJzXEY+OZneSrhQetMLZTd6ReMuFs6NF34p
xQMk/kdX7I9Sa0dkr4qzbYelOuciqt7lLwlcMXfWQn2IgYsgf2HL3bqrwq7gBGrl
2+ZiIZ6USCGVAqydSitLecPmOpFC3ICqRmK2J7hZmRJp8I60eJI2dyO61MBLHtcB
udgNV8APBBO6qwywVDGjPj+42ImTycXH7Jr63i/Em8KDXJ6SRnv5cR+hsSX4pr+v
E0ABil4lq1g/Xj/VsjG8MNzmcqbeZnvFPqFZR0bDWLKpv0WL+Kf8Aj+LlG/r0MhL
IjcZe2bCR9B9RsvAWz37WxxQ617AwlW81VVOtOWwq3WzIuF0f22XpYE1D43YuQla
314kHh7CYPSOPGF6iFAapfgf3dbxRmNvDWvk8h+39xnsSQL+BYuuMA/aRzqf1rD0
rmjiTnjq0UhuiHtaDbaExsdFYaDyYaKNi4m5axoPrIP8k9nfbE2eADVd/IzSKlU6
L5dVv9nzlI8yC9QTnj3ItF55lOG25Vk6PYrcsQwp/EOo6CNEROyvtQdSw7JZkvli
z5YCVCByomq9fKX1TLC1xk46MgRNdNXPApDj3hH9lNZ3FEuIgpZAWoDMY2tiPY0D
uNlFyg10Re9dl3R7XydOiKjGouc1H3f1XJunEyMANz2vn3Ncd8rXIe/ZZ5H0oIof
kkngoJ2Z2CkkF/OfjLrrW4la7nR2asGpOcOkDrYtZ8c=
`protect END_PROTECTED
