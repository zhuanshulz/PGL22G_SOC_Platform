`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3M9B2Xy5tk16+jJvi7MmRx+7d0ViMwzEPTpcLSQtZtQyrYF2E7YWMcC75MRw0Z69
E9X29C6BF0tB8+jQOLJjdegt3Q1lCnUn91kTb0oymJtjDyJrFC73I4jxyolTWFXz
oUwgtjtfPHzYXw5c59JUd8sdhtUqWqWtp/HGczsCKXblmDtXG3IDJcEaT2EhXLrW
ZtzexufjnXrX4K0mu1m18DqoFt8h0qPfyx01ZqzYv9ZpcV66pEy+aXflXuNahdE2
C7jGD4WtBfAD4PBgtkt3Nl7FiBcrSMJfE4tIKlgS6819RGqaEYnvFtzRUucZDJHo
VPmCoAXqRgu0smkfLFJk1sm8lIt6i+RS0CLydKHGZeHIJBjl9raK9/x4ZgXExYj6
LPGYMLRxgGBUIsN77KNYqG/U3CYtPM2YAM5Qxpv0PqonyBiBgN5FurDmYXmN5gjx
RNFtnF8OgQ9kCQyIgLCuUcknFVvigzzaoHv31DOwueXKgU3RBXU3ZsLXQ+cJKRrg
ey1V6S0Qq+VBy/IQyE244ZYdb6TAsEu4sRMztwr6Q+MJVBudf5Sr0BLeLnpaTISk
9tFD4Sb4NtIhEfy40DwEku2FSb80nBW2FcEW16MXzC72Za25iqaryRnKua0ulMGB
MnIHSgQAMgZz1cX86tOvIhdTnHtwd0ikIpX1IM7PWDoCnzwYD6UiTqQjIXC72t28
C6HGizv5dCmpMsDGkBXRSjKWrtYKFUzTWPHTPbq+Qi0KdCE2U86tTutyuqGI8Juc
xsuOsGO28MbQET4CnV9hHvrYPctUQkfGrwmMdy6d1eURFgi1iGE+Q0c+8VZosnXg
OAsAArPIzGU6TfDJvaDrzbERBfnbJVHdMCBRBIHnhVw02Zxy7S09pQW6Ds9nrg5I
R8evOM2jYsp8MfBXGnLnu02hEH1ZBbdTevxzyuRWuWPnElI6rjI1sK3+D8pdly//
gm8Uc0ycaGvkXe0MwcxEJIG5GYlF7KLWjVvsGE605Hp4iwehaxYuJZ87/IMdnIR+
D1tD7ZP4r6PJgesJUox9UoUQamW1NJmlPkI33rkY3TpugzO5KDIwF5f8U1k9LlfH
yc2JrX1CyqRBonZzCyI/43EOdMMaj6+03rhTC+331iPdSCjE9jDbD1Q1Fk5pocjP
e1qSlL7li8aCZH7B9//pcXARyPgD/YErZffv5w9lxoKdpGFxOkz8sfIrH7wl7bEA
NPTLBh1UAwg47i9A4guYM3cXj7nhV84Un8rLgIVM3Jie0ixfbbGWyRumQ9xizU0b
+CyI30CEIWaruKWPuWrpzHzcLVJqcnX2PhS1xrtGuyGiywLjOaWVmIK+VJLsXMck
D1CmVDZDgsxDqD/SXoOuag==
`protect END_PROTECTED
