`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5dCT2xkDahD/9zPM9JP4rJ/i8Ni1Q61ArG105boAgovMBbsdgT5Td0mqRs6RYzA1
4fuUg2d3LrCwy/cw7UEOBkEp2X1BuXtAFKEX3Q7VBn5Y09Ygrf9J/bFDMbSFM2Jy
k5fWUuZg/N9jISbiTbrS7V8OHnQjlgBksx1YyLwRmEWWQmXQKwB346Lr+HfrFmJt
eba9OWfU9ck8KRGCcxjf4frwgtoSjPBvgELU6zpEkMuZRihQ//M0QNBc67JfN+xG
b/6ytIAiTh25FcaaCiPX030StZql13bquGs6TliLJEdiW5piK2iwPAZ+MtInG8yx
QK8y1IqY8a9rClBNp5O2Vsa5q0VvtUd+wYOPAnDTo1uB3wMoOf36/n2kZH+ljYj+
GFwEhscID1h4B/Ry0jfWdmSAuP0xwUuORthahEgIfK86OsNHoa3qzvn1iN3WNZwi
UAH+3R0ecozE+6sclOsktsCWG6f4j9WAQoCO/lbmQLFxp8T6dzIc2bJEHWeAB/R8
PwFVgg21J37RpxuYshvvMI9XjkT3EyO5zU8kmfWjEw4Hrl8jXWx/g7sMbgB22oIQ
OjgP3QInNJJ7g1tvfvsMBZqWxq+owVsHwYOJk1IC2aRElwx+BOn7OntOo4vtcYs3
bXxrEdGG50WZl+RTUTOLqkSNprGC8kpok74ey2kWphu9bSoWIgVt6howRVD3p/OA
6CnLB88Nzf77dSDDBFvqhRXjHQnBeBNoFsUu+3OyBv941yG2UU1xqWKYISYif1x8
+a/46uHXausQByo61oogG/bazlZoC2E6mNXEBc8PdjZiGAcNjEWzvgryrEy44JTz
Xd7KYsAlXJZO7OJDaCE2V49svIsd0ZVX9x+h6ZV62uULI2O73BJjNlYAnOlv6V1M
Cd6uMPRScbcJJKhEw0lUdjtBOysYxTpMUFPBVTzNknu8ho0VSyyKHxYykWm/IbEi
RK3DDfhtrZYYL+MxdEgk2yWcVosOtnD774cEOnhEcUbeAJZh9uL3Qz0TokzUaxPT
z8EySy7Sgu5lpdpnBZ9D45JLu8pwJKr0awP3oZKUhcb8jQIi4/kuDhHK9tMxRqOx
LEfDXQXdEZtLMPDogtt39I0p8aWxK71bZplcNJ9mUtHPbn6TDHoqvLzQSrocA33v
I5pb9uY6BkDNRk1H5S0wjjfHsdYV/+CwAUrOHbtMQ0W0W5izvVHjSCV4JRR6+uPW
usgyEslF2xrM5cjTIVeIskIsPVf20nettjf8RoAqGLzt9UpHSRqXcqmg6MCC+lgV
T90ur0q/OTAesCNRtusJR3bnttAKAldk5EX+DdVD6+1MdOc4gKFfheSRD0foR9Rj
BeMbzUP3Inm7QESP3lMuHfsj+U0TCKcsB2azbZAgK29hLVWpJTcV8aGd4mGReJAf
RQZU+3T99gBLEXb95qZnAlJN3J9I07dsARRG470pofcKzo4bxukkzvFYVhm/q8nF
T/DOmQ4ceMRg2w2tPSh7LWOSR3POwUhAcKyjweMt1NuW9RnXXbtBq31g4cDKozt1
l450kaxy4Ym6yiBTvmud3JcEp0maVsRwVzGeg51b6m+f7q3u5ZtmbruVn5pRrkJw
MApLsVCUgstS1xCT25d+trCxtaxHVfQZ4gYvcsWbkBorkaqIi8zS8iW+piPoP+L1
VgO83fsYdVpmj6UDlZIws0ffinsm9+lp4+5WXmh9Slbin+A/CQzEtHVWgy02BkT5
Ac8lI+7Vfa58wuhZaLE4LCinwxIG6iR4wiiWFYL3jLfQFXqzqU/faXkff5Qbb+Vg
VdnmXEGMZEqUQFepOgK8cXfFSX6vMnTXPu1eWF7XpvfLfFJ7kSJ7WRGHQeapAi7O
M/HmpdzEMVyHgTNOuGse88UOUDtMzckEpPNajZdDNrvVXfYx8h5829U4EYruzmlF
4BQiCn2ynXsZwPtBIBKrYYuy95HFBkooO+evyIu5l7FoKa4C8Z9AeBRMBHvTdHeh
GAs9ZDgnyVJWQkJ3q4wsUSgYWzFwv1EZEqb4txnSd1AKAIjmS6usRORBCbHSsRGB
HhCYFSdu+fIY7q5Fsiq/uDPbspB909YJ1Fwpg08f3R4eRH6FnDhGAQxFDJ4bV7Je
KEoNenjpVtcfU/8VQ/oA9MboydzQMEyWwILHC0b4FlZFg1CaO2JK5Vvu78P7LEBC
G6NmAJTR6N+yH4PMyVI6f/cexxqb86u6ED6dlkTq+V7StUrrxA3cjTLXY+XqP+0o
dmKG/m2JZqxrN/yicChG0DIIvi9kEBgYB4RGBcSWNY9RDSbKThET56EAE6k9OXaC
9qnFDnEy0ktwOEyZswtUNrmntguoMG4Jcn5Am+Y9QiMmusxumE6o2AoqZi5KnTnK
EiKbHkuoPkiYNs2HWN077jyIS9viXYNBH+tivUWd+qUsV86UJ6Rjobw/JeUUDNRb
b2AtK4AhcMw1peMisWyem0Y06Ad2myKS7gcNHKu13vjh6A6Cmyb9R03TMFM4N6Jt
m8kjNI4PsjgHSC/KsDsZbcc3hDPUibCiidBx9kqYsWxHNcaFhmA96utEa7umGfuS
uXyf+5X6H04FTnH7BDqz2TM2Le2MVsgnhDTHJOeunuSA9JqsnoStQBXf15mW/958
wvhSESovX7hPxAavwlnRJeGNBNTuIUBbOqFsYPPkTmIKGOZ4KZ1V7TtkYEjLu6Lk
S/6S0b2BhhvzYIvB2BGSXxLO7rDPSj9pdRUjsKX7DbHUStuHluN9f5pmYcNDVBRm
5aQguodGYUvupHee4tsqINKyAAXX0ktZX1V3yPvO0af0jgWgqC+9upqfkpyWN0/e
f5AB2UlwMGPFtZPLSL6YsNUnE4SutE6fhHpsUMKxnMn5hJpe9bo8e9mCEC2gU5rQ
lDDzTcgj56m3sce3Z4x9HDTVDqaV9uGpeRnmj3BqOZaZNpmTMKu7rfQnjrGjMeFh
bERE/SBO9AuJRB8iybifuB4zmTpZmtFHd2995Y/3hhuJJNowC6yJGTXrTGK2tE4Z
OiAQ2W2532VC4P/EwaiOOowK5LXDK9Nb2yxXAbDmORRydvwWmJF2QOlFVmTHo+bc
kFMFsU4bwjioCN+grxSKlzoSLjkmWyM5C8kHBtjLbCOnUE8ka6CBuaL3hvaKZ37R
Ar2T2wRYSSEjXOt3LvCtdKvY9XQDQNin6Zs4791MsyM5hs0ueD5pdqVXdRn0+5/b
B4YKMLbiB23652zIwlEECxemtpBSs+hrFM8JrndAahvc+QSiOtPe/d1ILeJN7tMu
ahIulYG0cZIKsFVyZ2HSgnvAWvaXLuPWM5HnhH4o35Jwk8EYtTjmzrtOUxS249nE
Apoc8eVGzjR9HVZ7mpCjZPyFMyZtxB0K7VZS2NkDrO2B6z/oDv66LPQhNDMnrNWh
qIvrxHyA9iGUzZGbQ9FR8MiVM6rsidmav/hIH6nQTUmCwhSzZZPiwM2qGOY7IECv
qOYSND91QwVN89q3aBbP3y1MsGAb4RoRiwF0202TXwl8RPvx7BViHdehAExbaPGg
sPruMv1T10okHB9EKzNTpMq92BMU4eoCgZVW8OnX2p0ADAU2UWOiKGeenYCDgjqG
5iZ3iJ75il6LdiUp/tZbEw9MNITaggdRtIYeTOl7rNOBtr63DoB/IXOxQirFEuMM
rQ6v872SPMhQ9m4IjCs1MkYm5DeBB5tuUFqsD+jW5NvrWahh6Bd7mehRzQ2lo/sk
6N3QobxFNJIIEzBDmKI+KMtBJNzn1ZpWLHAqns4zbJBq3WadYdX4fHESvPr1Hvpf
+lKMzYwACfgfg9/1HIlkhCmGcqifE3A7xnF1QK4xVC1/O4HqK/3Fxs7NOBSlhyAE
YAkzXCBKltRooWlgNmnkiOJS3VALn6jxF4yCHoK2NaQPvpl77qAiuTxOtX5u7lEu
lnItRPhsWycMF0htO1MUvwX1p3qVZRseEIsZT3DP9Uow+yPAApuCfqwq4NGHRuok
5plO9kQ7C33/fvYwj7V05at2j102bwP2vby7+S07ZXEhQREPaBSkE4QbbY4dL7am
ZFTKO3S35jmvt5u7wr2Bj5OIAh5SOsO977fccPMhL/vVOmHt/LKnRcq9gCYeBSKR
Q1Os3uY8s8zDI8NwWJEkW1ZErt9uKMZN2TZAOIDIqRiPRei3ssY26b7GXksSMG5c
hkVE76QI4yiQwidNqlGOSXFYxlCIka+O0whx2FoB2ks1LWZTyAtR3X2CWsBCvZtX
6DyKGjbjuXDvf/Hf+NUXcHZBaF/KAZubjcIUpfs4M4dXAnVRnqluz1fafRim5Wpu
UGEXv7yJh1gNodTndaTgscmJTovOPlEiW+GjB2wsmzx5sG2Hx5oEx1whLhy763UL
GqnUQBQ5E2luwun/R+//Jh5V5i/KScNVNqGdHddMs6gWt8ov+R8GULLvdE9TlP8i
5Sy9mQVBXwW2z5FFSSIl1itUlprj3gQ0fZV0k8NqpK4KMSrtqvVwAVtGmEC/tNnv
zC8Je4P8udPS7nG5BsN2N+oxrpZJ2Vx2VqKHYM1DHNVG/HiFh3QKtGYuk03OpI7A
LHv2iEccAEby/Pz1T1t8DIv1bI2J40zKOXaFRFaf4XMKl6SXwOUyfI5WF+ptiFRu
nNPWNygDwJ2ic+7JiXiN39rdfkFHJpfVcXprT+mL/kRLFCyTDH6dSncFXn5MhUXV
c9LRpuV2dWdN77tQmGwSljGMUK/7DGc3998158Ul+NJmCE47i8ji29ounksWfLc9
LHttj/P00FcSK4uX9nIZLhUXdcTBImNAOC1Al5MGhc3NE7/l/yJDUGMzYHpS/8F4
8OReXU5zF0uKKkUIJheA86czCkbvcdIOT3NOiofWwiNPwX+hjkO8CYz4AVmpSQfw
I5js1/Nz6LIm0cwEEvW1gWlI1OwyZoDb+XSgXH/cBGmTFmijfnoPnIuurpj4riFk
fJrm3TTHX0snfaNAYwF1pUDFa7ggLcwyEHrtySluRMCL9DODXqtu1W/3obqHQ/7j
V3RVQQvGYby7+66vW+WEAYP9xzffIm/11fce+VJRfPf0nD210bxVTF22umzy7HJo
ay16a0SJqJ7IfU1064HS7O+l+za0x0/r5knJ3dhho0O72+Mp/s6WejwN5PyiInTM
91Xe9q7H7kHp1/m3xhKuNQ4BRIO7HqgYsjFB/ai3nbLApe5RLN+9hCa+wRlHEGKN
dg8cONb7oP03zRDzztc5HjWBf3A18w6ErZKQja1n6vqDfsC4b+SAn/48AIa0IOlI
X1aRrWTCIPSyp0UaWjFvyWrByuGiIeOU80DEChcevvohJsB0WadxG4UFnpcD+jaP
0j03340c5McxgQKJ8ZcdI4Qxnfsx9OodmOsWgNNd6UjjK//EZsCtmSxw/V7FQ5vt
cQ1zLOC3ir3LAE7jY8bfAw5JvfITEz8aQKyBBotkCXqlacOGxUHOvagUsu4pYTvx
/Tv65q6jdJ+7HWJeUAKwvEUUasDGCEPhVvwvng8x7nl7D4ntqFRbp9REmwNAmZWg
sgeJD3tttr6Dxu3FU4jbroHgv5QGSL8geruk999RhkfuTp51KlEPXs7ugLgBmDbC
yIzzVblUquqPHcrQpZ66fCmHbAqRBkRW19ydgUoTFuCkGM5QC2NAVNH8ak5PvwdC
22TqguCOR3jHpMcJ8/O2SjSWV0riROiVcUGWmuTG5vwweWY+LdhZ7b2ym9Hoth8Y
mP6mqCEWng4zUD1oXXOlYbrjj0Lbxb7u67EPKzLTIsLiQYO3d3mTHllYKl1P8wxC
/pKS/c3UO4v4rMY4xNGIJl2YEZmcTh1edccXL4T0Jz6O6bDxXlZv5KFFyNs3V3cP
4I3Y53lWLVrkdKhQ+e/LqYHzewLpUqyV13sK2ln/SPfDS321+O9uEy+zC8GPUYgv
FVIcjKaYAQzMZNXPzy8hMTtIq+NpWTboZZs80zAPR1544PJin+hOR+r+KT6WE0Lk
FIGmail+M5x3DEqC0qsQzXK/UI96lAjjj4uwGm6vPU50mIWOTZZ0AURTY664ILa6
fE1WUemCau7xdyXgQXUwz0M48xw2pDSQOLZeoVYrM2EjHEjjbo6043BDelRddlHr
odrvEYILWMmnVUHxj3u9D5WzdQDs+qGufuoNiioAqOEvP3+9araBb+iWOtCB4Ljl
ZaU2WhrjDE8Eino5D3+ij7bDM6p+h4WueOYJ9YymBqPnJ2tc4+zX7M7WJN1uSAAd
b8EdD07ngDiAoHWHbGRRLG5hLN3B0D6HgPxy99s7VgPlDNZMAxelTH/fIvhJ0RVY
d0rFeyAh5DW6NbR5np7Fyj2Ie/oQHnARbbCp4FJvPOyNPQJbcHV8TJRvH3BgB+JG
qsj7x9q26yZAMsMn62O4O2Haa4AZQlEmKYe6QbY5dGBDacIfRsfRYj+CyUROTwOu
x7t3hMVZDHc8DI84pkSmHgXfOp8w8AEOrOmeb1BHwaEJ4i0q/sqPMqFPuNf53VvZ
Vzs+7OWVxDWCLwHmI5j4ZeURc1Vv8bE0bkbBVADHLgm2J2Y9W3uo5WwpzyqpIBIQ
/NBuYA7AR25W8j19opGp4ZvgNUQVQHu9j7bqPfnjo8U6ba8cLS4DZm7k+Ocw0x2n
S2h+AgR5E5U45ajHf0uFLphf2IAqCX5t2QMfpgMgsOnNV5+Mh6aV9p3gqk+ApWo4
MdLvUs9MH8LffEaolhRMyhpB10U3OdtdCtQEbg6ZsxbUWOe87t9C65STFRJzDOWb
WbQr6DygDmx+5kF/sTu82u+G+5teiMntArWgQ6rhjERYezZSrxUCktPFTeIL+HHh
tuJoFttEmeGK8HdBjvIFoilGlrZvhP/DEXx7ktjapgMGDdUiWD9kZvMQHeRd1fWf
ypWo9itMALL85YM4X1zxSfdVIxnzIn1WYG4i7VpAG3Y+cqfnKJ//fxaJ6oz88R5m
7gOxRRZKb1Do/Zj7UZMYNS3fsxNtcUE1XoX61Ts0YJ1oemmDXjP6n2PPiqgGuOP9
B9M82H5/3MEGuwRqw3IKPhY/k/ab9NORWFC7qUwaH8UM33EdJMoICrA7cwx4RmWh
XQpWeaKaZTv+la6gZYHZU0wwG/XvKh5G4Td3vfEVzzuQ4alx6aHqHc3v3PLEOCmL
QXJzN2ejHgLVY2xzp+1kA0kCk3eEd1rY4LVLH+wd7HSOEVpaHrJugc3d2RDoBfQ2
X6gu3N/6op0zO7DJsZV2oebKzWLQnzgOLt4eiH7BgCwKzbNjQHK06f0RE9fWMjRG
63kIoaqSJQ+JzjSQVnXmpr93gc+JErBcKeHrP0n0evAi6j9+R75fkNnvJL2QBEON
JKcCoChj5NieNhLKO4eD8W5asr4Eg2O9WVdsMOuDJNbGn6NadFaASkLxPEZrMoS3
qVjuUaEMCTS0eiRM5AvCUMhGNwHRCYu8eTle3ZqsLJIOJuj5WOTT3Qk0UHPcOgrL
biuXRoVrRTeLj4nXb++JCsWFrM/YqYL3ANwQIV/oyaEKmCtupfIwwHCaS7XY2Ss5
sZ8xhvXBei7T7sUWGb9ckqCsXCa8HFYc3f/WSJwus5pyidqArKmxOPMsqEJoNjob
qJwlYX+6VjH+b6NyVmj3kkAJnSBmGAq6h63LU2KXY5AwriWF9vs47TcMoWoSwrG4
Ljh48RS/yv9F39tBLvWG6PVIpF4aj2niK/XFDdzzSDiwpSTslUT304cCBE8ipI3T
gG0FudRGq3eK75SOqH0X4k1V1STfStidTH8K/pYGoSXniaURAwKc+IA8OjUKNY8A
6oCQ+zJNwqEjgyqewAqIFoi1d/LFIJrBiwWp/siJCML/LNOK/dFe5sLUi7g/qAK/
IbJMlW9WJ/lysh/TvS+Y3/8w/Omsd8ii7hVZhnUCS11/1t/KMKl+h/4dXM/keacU
8EDCQXmOA2zlbJYfnA/clgZXX2n1ioQd+u26O28BV/dbAMwjocQC5qXk/3p23fKL
BntZE/Hz3mfketJAKHy/xWF7p5I0+7vGIHNhZk7feKoCBoYEufPjJOLbYIY1lj/2
JQjiuEhNrm0Pldz1+1yq7+b6ALaNrgYb6xQ7qfXH1ycxXMZHQi4eIHV+0+Fa/+MS
Hp+tDC7vFTZ9lk+wkO12aMb42IIE9K1foYm41PvxBOZRXnm5SJmQ9GEmc/dytiYT
pli6Y1Git645q+GxBaJ8XukZUH/XCJd3TIo1IIAur1ZezIqTplbkUwj6SS8Pxa6e
5r5x9VJlq7o4JGp2HnlU9lnD3c/Xj7DAaM7+fDd4x75PvLpgOKjMqppwhiz/WYXF
6klC14xxpsAkgQ4SyyJp2A9K+LSijY+AAk+NtXW5EXh9qsij+QEy0iH7/iQteLPV
hPvzQsdnQaHU4rAky5AO1snF1VjkVuyApUSFcmfu2y2gCW3qiMoeygxbayeY3mUN
aS1kBKmD+BHQ22hae3qIAUmhJluTPphcCSFeKctaCTcG2O1uzXs4MKTMMkZVLx1Z
q/xmxKLmS6vyJmt5TmjQtdtIJvRweYuRLkLnN3+qrH5oSc+t8AJ2Pladh9OdKc71
uD3KJtLEURfVXf7z9oxftddLOMSjjrXsjVE9u9hz4og=
`protect END_PROTECTED
