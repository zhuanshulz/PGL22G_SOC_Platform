`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fq+MX90bq9ewpqysENHQLQum49CvMmbO9zMVMK4lbnYXC6dopk/zhQEU9i4wNOw6
tJA2fz44TxMqxlWqo0eaguf1plI56ZoZFFKqwg2pH5HNlGO8czeQmu8YWNKEcZRR
t7lMmMaGKkWKsEi0amo/w9ydYWuVqCZWi1EMfnPIlDFYnNf8wjDZHjOa+FxiD/xZ
qSLuLLpe8f91zmHyWnfFCU/yWq2eVmZlvMlfbfi0W+/jTXXj14nXsYrPAxjrDnHD
rlpC4uXCCujfudh3l44dbNhPCqbsiHixNb3kJMR2MC1JOAFKKe1qt803mpZ36xSt
wNnluSAx7E4PaSfLgfQK2DTmWeQGAy+aFx0/T8XFFco+DUarA50HJl5WusN++R/c
HBJl3Hgs2ueDUbY8HHD4iWAmUgDyYZWhwq3tbvhdPfvAhFHCIsIoDW6ONIDJNFFo
B8yAv7QHi7ZAiBqafZvcm5kXQfzGklhz+P8w9z42H4vBo9OXeYdC5iMjNX+aqXtH
jsCA1/Wr/C/da3LfBxmuRgbtJERo8PUvFdml6uAB8ctJk2anKxH8jqXh5s7ZoIax
ktdKUSfzcwcQwJkRG//uH/mY3ACqWzKYTrXdiVHmZpaZw7t7IXsWFfp7zYRTIQJv
bo3qFwaaBbsz8bvmh+tw0k7VM+wjwNCiVtWhk9TNY/ycmjNbXY7fuHJDYviuvCuD
sbAbBiq7rlMll2ABHX6+WbBh11q9GRitPyN0wbTtWkt2QC2VT17mEe5OxLssNKQJ
q9dTPh6UVKmssq2+Nn/VwRXdXiIWVHglkI3N4joxRAty3lsGPYpaSI3icXtLZ/xD
IOt8/xtIiGFmGUpdVkJov75bJVrbpD4pb+iYaRa29nJJP4hMy2j4F7qTKIWBkOFK
cvJmUarXUXoVRyLOzBYsDxQM+70BkDEc98NDH9OP8WsKaILA8TiMDoTTjKvcSpcr
M3tewXLn/HbsCGaIiWZGn7U3CUn7l7GRavo5TUlhC9KKgqKAxm+CSB5IrtlcYiDW
uMrx0EIO/xdEpBo1nla5yja2fGu1Rc7pK0zi5aAOhN+zn4HcaCmrbTnUOKj+76zQ
jZnqyqArXxbnC9mFbebjfi7liQlWIVRxXtBNozn+JsAPiMJCh1iRVAtw52asCgAV
/RVA2MpnHRDf/5ZJJemYKVwPBQ5cAv4Xj5AcJiG6ieXLYBj9FYpICCFKqmeUwoWb
ou37uKJwmB6Q7aYUe6QOwV3XnXjLsFHRmyHHf9CYCwY+s4z25exdQr5XpSx5/UW+
zDLOxiHaOkg7UDK0L+vYjErZv4NSh7jrm9wBg6D5quCEmDSVEvFqKgMvkufmU/TH
QnvklDIjrGM9HIz39FCvSWhlmolNw2iFtdvOuCVsGWpz74gMZclAuE93sx/vK4W6
TmR//SqYqln7FTKloHPvN8VYCqfobeqSDrI0OeGtX6wASyaLYtQ+r9fBiJARNiCX
x2cnT4kkW9UP+B9pTySdS7/k1XPLSVSNaFVBvLYiTNRZQRwTGieb3HQ9hwxqCenN
34NktStBCKlHpoOrp8tLe6lte9CFBiUBJ0ahhf5nmSk4b0t6JwltDTsPkOEhHSYQ
IFdHNEt5T+HEcLMRbxMYGLsaqgew23dY60r2e5OTroT2WT3tE7Jj87cJnt94myFd
fSdBtycnvtqHYBSoXF8lPmaOfgiTZp14HdG2PM4VutN+HKW5q49lJyERqHc2uvOI
zwIvsq+qiqyh5TZ/cDCD7tNcg1N6d39jYCAwwFwsHBKgs3vnNldu2eP4TpXhYBUx
UN/d2ERbVO3yuNyUoW0PhtkLddQ5HnVKKGiho/Pv2W3zvLCt2864J1sfofTtPiqc
S1dtM/hycnSka+4dgrQ3W6ARDbcITfVfo4WRAXvxAWw9b/CYKvEWemwyunPMmZlC
WFDE71ac9imbGp+RH1QSy4tZ5Xo5VPuhi2BkcGaonesTM+32CoJRgV43lFk2QC6M
GjAAV+7vDRmKjqrw+BBVmZcfXrmxATjNXUlULxmpnqREMK/gSG8GEKIIpW+HExEX
0DQghkoYF3PK2UHjm/EYM/8eU/K/pXHWlZYnGUT2ALz0c5PP3Bdu/DmEryxuX70m
8LGxAjL01t/lyVDI2SdFg1L9Bx03dnyXqxauLA4FRDAvP5bwBW997lT+24Q1e1uc
HvMHQ6jtKmavpLUy8MLaTIjX4+7d3Q4i4/6g7jGESg5YrtkXOKgZBVq3cuNA5YFL
efR+cvzqEQ8BO+vY6Dkiqg==
`protect END_PROTECTED
