`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TTJlkkqZdHph+weNU2Y19exzjDQoyQ18aadgAhLvFJJOi+EGzM+WvAgUA22bUa+O
Uj8q4Po8Ao/f7E0tNsq/KwsM0iT59p0g6S62EQD2oR+3Z6u/MrCTyJLW9f0U9fAN
R6WT71dt6cBETqnLAgnQac7EP/sNpFkkNFS2RHc27HPHYhsNXsxwdLLQzMqoOesf
AjZTzlbFIn24eOf1OLuQwbxhlXor8AFvseYgLwMeo6XFx1JjxgrcpyTjDVquOHgr
CcapKj1qwy6nMzJKOSOE3trEVpsNce6PUPLZui/NfhWtuvWd7wEWQUA0a1I3eswM
SvkJoQ4m9DuhChlitZPWyngl/1G9GzYopdVlduQVhh2M8hsS4VJQ4/T+I+enbEPq
X1VwsmcoRSZRxgORXrxMyZrYtV3kLh1rfZAtGwBb439SfUFgQmtdKPYUZ0DJficF
eQLNnWhrRPbkwf3kaqX7KWGD7ByZ7Nncpz/4DWBKE9lWFYbyo8tw1UXalb/nCoJl
hO7NGB7S6rIgpufV386hOVg3pz2DVyLqv1DvE41KKAdCXwhjAcfy9OAJnLZiv3wJ
aIcfhkjrcnoiYyo9g/IsqGOjASAeQbROuc6raBNdUp1EqYX6ihyDzbKzfAbooS7e
DbHFYnTzz5J2i2Q1aAJydJ6UnF6qZQ7hanmpZd3xaAXlVvy+n9yPURBz1rZmgHAz
FTKzkwsg2UxCRZAq+N0/GCZH0+pRPenU2f14SdXtiOqUTIiskiogbJh+llV+aXyK
TFetVUSwC5ZUuPP7OMwcIC020Q2nom+0D4xD4jO9ci063/L/lt70GXhNivE4PBap
sFgBYZAfUeieYIL4vECDzT/SQKZsA9E8NFGH5cGd3mTAZ0WMehSWY//0lh0QBV1n
69lLhBM2OMFiyxkBObl/FrXODEEdBRAUWqBu9VxpqxSkOy/RZf1ZMOhhs4FgTvkg
`protect END_PROTECTED
