`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hHW2A0b4QOFE6EYl9LCXf4Dxqto7jx5XiIKGu5kS8+/vSFsPikWri6up+N4q7+ZH
VLFPNsdN378xLU5Jy50yy1m0cX5WjX7HNd4dwr6kMJSiOiG7iPj1rFlvITLFki7c
4gF2Ltdyb4eh5Ovfgr0cMRUE0FE+AY9OVL9stM/BvsVUvpbQHqMgJA5ZnoWJqmjZ
8q4gjyrgH/LcxWxm2yrid23mkTKWC9POuDe1pN92CtjuvTRZckjQsC1w1Sjyqbou
s+zJ6zbae+2L+1wgffjMtQ==
`protect END_PROTECTED
