`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t+gemOw1rdTael0nUTu5HfU/Qo1vi84RiAAaBS//y4H6BNCFj/82dmICnMaKvjiD
rzunhUa7POacrsWaFE7uDFje+UEayVMSf3cSENKwUPtKm2RCf8tHzuMGqdoGPpIG
X+/P2g5q6kkwcxytEFtLJIYFuAJJBucy2m140Uaemkq+tcJSLj2JlQ9mWuAvZqka
VKTw6jARhIEG3N347FyMnVVqKwZGaQZS4wwrOnPbT6+lkBNpnb0XfaV4QSs/H8fJ
HEM1yl+8DlUUFTBMmiw5XHbpdY/HOqrYZVf11oewhr17DlMwM4WLKXhc5gqSpHV5
W2y/t49ZSu/LKLQgO9xW13ls7IURDdads8MKBkJoMPc9Ol1hJbovAq4psquSVFcf
bI1NAABj+V7cnw44PYET6vtBh/ySE/Kq0CFzx5iE/30mMvOfU9aqBuDcbNODJFWR
1e+xBG0w/Ld+lbsekJEAGv118LhN5kJeHzV9ve6xYnG6gLrl5DqHoWHpweB11isd
O7iuVO2epa9T1OA3sgxOnrk19jBFYtyrIx2FR4uat8ugc/CwOjA0EDz6prkO3K4C
BLsDXn4p10+E1MeBPmrAuytp1hxTyBWQjq6/qKwcmgR5L2FR4OICAYtPpKMS8iBl
+tKwCxwH9v9FQ6cyS4i7a4M4dCa9vOW5AoDnuKkVQVTh7YZhUkye+XqnQ7RPMP5c
Q87sCv/Paeb115rH7G+lw4vrzr2zJdAbdfsx4rFFyCSsia3Q8F9FQInVwC6/88hX
jLFUnFZsFhXw9UXAyrPt/M+kH/ttAou/VeLbqnLjGysGB119TOvwLNLjx/CAoI2j
BglIUGTc8f+yq7/PJAl1+VBvAUwAm3hp1zCyrq9R/gXYdl1z2xqacG2Ay+reX/o0
NlfYIhiOSnPfijMqYcPA8D6+xyIWzirvPPlCghNMBjBsCQmPi3TDDDWVKifclWA6
JdHXkFR0VUTzGGcTWnNTPN0doigT6dEZVPBCEv4NIintuG5SAuZhY6ZcYtKNQF+g
WdEaNor3VvgEJdweorz7c+R/JpwPumT/vcdQfoJy69sIytfpJ1J3DxYAZ//2zGlF
j1P56OJoIuSVUSJcwRgaLCwaX67W0Sne8NxXhWW4NyNjGV96kVFs0tMqSToRPtjF
9E85cA4AHLGXNBrnezg7uvGRzLddQlZcNYAbqLwxqsDHUzOr+9QvfI6Yq/dDZICw
teD7p9eLU57N2SNREypzikEITkGvO43rCMcWL80V6cdbBOjbffgD5gnowv4mQKur
tXasZfMS5zi5xUOMtpwPhIAivR1EOVBmFbKD3kph4x5RVvUswEHnCb4NHHM63Lro
54b+6RGqEpq5uzEO9PfjlbzFNIsvSGN1VopKGtnZQsqKO6LBjJeS2B7SxOWegHOT
JLcGHENlzoetDBVccMLFQA==
`protect END_PROTECTED
