`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L1jsyV0Oaz2HE/B9xp7ULLvuUWP5l5p4cRjWDjpgzhFNzxalHfhJHtTTiRMVS7qE
uBFOx8glWn+Cc1oNEPQsCdntOSou+X1AFGq0x6J5VcX2bgkIjgyTayfxDjIifCSg
nNctDDYRUE4HqfXAktiKnLK8ommYAipVuxT3vgVvpOTCFpoLt+M5N8Z3jtY3XnHJ
dIbUSkConqOgMPsMCuBiKTDa2dHXVqmJfx+kE4av2NZlOsc3YAoGooyiT1ExUw/O
eHC+Buz+Arm6Q357AF3+VL41o85WKustmh1+1YsjFDnLm6pSaM0MPu80bEuq20R/
kvh2GhOnFUZg6lR/1kYIHl5+pBpFTxD8DpAlmHB61O53erySGzqz6ggbz1S/R8mA
j0m0IIOS4lhpg7C8M2yWFUDcwEcMX9F3I+PirCwj54z/TBF1w7IvCFRL1pvuLycU
6DoibVzzoO+TVrUm3S3YisQBDXUp3VgakfCteiD76cdp2x2PICMEh/X3md8Uk0EJ
987SNfSgKHBelmDRAf8ViFUXpaWSLkvJNSCtO5UpOrqGhMKahP5JBA3Ty6SGFOYa
reiabFpHMC1l+4pwFluoPPHOIk/igXtBPhb9omI8yFT4V3FlF78x5fpKlyFCLaPH
2P/AgGQXSKNgVUO+NGC7ndIisvtPVpTjviT8BUyDcoSsWAB8xx1QYEspV4L0P4QF
BBG4CHtff1FCs1gFEEsnXriIpqv6DIMGc0PKstybKp2bCqxO42soStNzfF+aC3JK
0Ajxtdq8fqaoXesuZHwmEISFjs33L7WC9vDdclAOajQSrf5CGfooPL45VdzrP5vi
48Rbzx15iKxsfBhoRtQAjiwsGEJV0xqJngkTAS1lbHWTo2gZvWzAoKzd07VcM8+E
nNzNIBBndwYH5G0148DFrUjmDZN6oqOwD61nb668KdHksMglXoHZVWqLJOVpkOUN
pghNYRWRg67YI3MOn7Cq7REWSRnpaSZ+WgZu+4zbvpnUzh/QPC99wDYMCJRgD23Y
cowgGN7SidJaXtOaHV3wuVxMYbz83uNhP3Iwxhl0TAywhtdkPFncAsmcJiDfikgO
jDsqDin9zqXGuGkRDnNYdgkgJlMs0ip15vhCNPVIjONRNLfQbsMZZDJvZz59HW7W
ayGb1a8ALDoNebcChBCpatBC5iM/kg6GNImZ54yg+UExfTaNBQMtaNEiC82OCd0Z
IXvvDu0GuzyRQoJB1ZBtNNUAAFyYsulGO9KJvZe91oPlBzk1Rv08YpS1ssXhi2b3
O2tUP4hqHNF3MV4ZHj96ePrq+x1j37WEgpIY9frxRBAPdh838Oub767YJbZTbZr/
GqR2yRTY9zSDwQQHfa8tHm+zzrX8iF60w4KinWyVeFuhDMXEShefkzc0AhOD8X1U
2Tr6y3RWfagseenBKPqxb0O59Up3NDoOELaI0+u4Ga0kHVcrWt2NWMZJdNJZv3L3
a2dnpcPjKS5uSHa9eGklHuz3l/4Xjgk/0NNJ6TQxeVTYxy8YOzLfPF2D9EuMTcGi
wGZkTTvEYj5dbRP5e2te2GuRuCYscir3MSc4kMaTlBxEAaNVozagjs+yLVvW5FSQ
0S+yRl2DpV25oj6UwARcNsfp57YRNpFGLaCOEzj1v+jyCd/jUReWEmzpFNECleqi
9vFkWBo0hzpO5dU0VBFGCUJ8kaNMzY0ZF7qOGQrMrFoJtpIzVc1HhsRFy63hMJt5
u4ZMMwTtWfi0DMWiMSWPMYsR5CHkXQK0XolXoVNLaVoZ4TCpf/Gqhm4sFftQdhZK
0q8l44SxHbXjQvBBoGTziiQb2nSS/q1AcPPJkPMPGdq7F4288vIkhnwDQvwlp9+5
RT7wNRxLcs3P82XOgd/lhf/Q7vWxb3325/apYCGqMiiNigd7UJ4mYYvlS/xPBjRZ
CZqib5tBZqaO0Q/nVVwO1oMA83yrnrTpp1uTZQFnEsUq4SVvqVk4fmRTXfQyMQyI
W9cDlBXl43fedsJSFrTzwrOQJerjYonzsZ440xs2Fb90QTrnrSA+umxoh179XF27
0iy6GDrl0Jp5w+qUTV/UfDbS0LNiG49zRZpMJxhkeQeee/Lkvl5hDfnzaVVqanAY
zb5E042Dz1+/sEKVFRIjGVID6IrB8I22i6tU+TK81n3akG6yz2c9tjwC/vslat2+
pezzg3wxxyYS7zQJ+RBbf/uK7gNrj9rK8d6/FXbo3y8=
`protect END_PROTECTED
