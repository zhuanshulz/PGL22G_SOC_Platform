`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O6gLZ2LqMp4q2NZIt9chdNQvm3pyIsFIoPk6Xo2jm5lPKEJU19iE/27n8OkZYhTD
aPaBcPu8K3AH/hfRfcqThsIw8Agp/vutZwhv8nbqAGk85+SptA4eIp8Lwt7AfRdk
bxdgJbKEVLGH4/XyTg2GYhptTCCz5e5+qFdX85NG75qeGDHzONMSdddNYPLSc0HM
OWAwbw/7s2FqtvG/JNS0HzMLUnDwttW+ksUZsEbkVlzKCBSBpk0gMzEzh9fONXP7
4jJKRK6sCKW3Lca+RJRaA1pO/kyVQYte8oq03K4X2vpjOhxxpL8XrmKPKisJBbgs
0M/xwbK+A/GECN3GuUB/IDzRKPYc78rh7acnKpdJfRonl023QyshGHWNaisajAC8
26SmRq2gFddKylKbUt6S+MaR7F8bDkScy+X5Vjrq5qkXj4GgXolsquhv67rC0CpD
miPUQYbC53rXSQn15S2fFCo01dZQXFzaFFE6nGQJTafFK29aK3q+8Qe9QEQq2sNH
HU89ROTbQGi2o1aJz/I6ptmuyi+1V9OQvASQ4XdnT4YaHqcX7njZQ9pS/xIRQDYn
u52v5nrPJAAaFUpFH7sfcXZdqfavL+7zPwSn6LM8WY78s0lqnaTGRDKbx7WofMPl
t6/stB8R/GNcqNwEH/7HjZo+G2cqs9+mtG6q4Bu1HmXhbRxBa01b7+YtVA1BCIFT
9EnDfPNb+h9VmDDJtMCdcmzcIqWEmJwBrP8ebxbGFd4x16QzP7zW7tCGLpyTInjS
Hy1CDPofFgnag5xeIsPKki4UpbydKXIWs8qs/kLNteZsz55R5DiDJVK9o9gJfvi+
bIMolPLzhC8JHfxwuV+lKzpfFrBBkqpX5dcJbCxtpSmkD6rxI4GFyjdgAEUN7BbI
prKdsKvf57+CSnLisTT1FfeGxYddCCZl/W1vKI54gb3P2YIg7+BoQBTq00Srhv86
skxaiZ9fZ8kChXUmzy6SrDQMMr68WoIll7A/x8IxnfRdfTyMZ23iu6N0wmTh0zI9
sxjk9DqxWvmuDPWvNh1KbUS+crxJsmqynsxRFyL65EUprkxdT9hNbjWJg3bt+/eE
TqfosPNnE/NZSvHxt71s8FtUzAFEah1Gl0SdwTGeO/r5evloB74AbqgQjxHRoEWn
tx1LlBGjTrlpXBFLr0rjbXahQAZFfY261qpelGgFaWlGIHxwz4Kg2sgaShZiO8HU
yusdUQJKuSa0H6WH+8PTeWFJ1o02oWPC6p6u5ZzwZd1DM8mbEr0ALorLbzH1sHdN
TAMH02Z7jhZ6ZmQef7fSzfnGlT7cYQzmQLPrOog+0e8ndfFPw/tn4R79SuEABhw4
effWuvuHGdSryYIUViqhFRSLiYqcHxKccDAyWrsLvx/xJXBkxUg1w6v8Qq5v2Qh9
j4TyzXc8VM0rGA1Dvf7w5S3FnF6jJVyfZHynmdVLAa2kiwl8C/ws4oH0GZtSUP3i
5dWPWcpnTbzYOWMGAFFREG1pUSahSi8+yTRC9AAdYTvfWVxioNehKQXiQESTKbRM
y8L/p+Ucx4U/C53PbI4TLIa4rYp0CXExXlTIcWH6t1oD4VJl+oIkk7UYq/cL5PPd
lVICn5xRB/3idlD3TYxVsVTPYsLov5XvC7v8VQEeymd0ih21vIuR+NTvswrtp1kT
BxEiGaOJyeFfekiecxBy59OrLA+xgnZOaFVelQ1UehhVV4qR7gXuB7nq/8dAeVbB
gVsOMPr2wE2goPod046ZIc7ii74Ti7lgyZygFofeowyw5kOjEP89KBpwocjm6MKA
QHVr5FcFmFrTCJy20G7zCE3tExViiCpcB0uziTzHVqPvsstTrSA2wiGXtWWRY1cw
6o1AFHSTaTz2K74XlM0cLCOZW1NnVg2djDPYoNgGzHOnVG0vyQQMigG7OG2zX84X
0znZmmH8CYWtsO2L8P6xqB//a6BE1D8HRpwB3BR+0TiGTIwtZCX/ordMpORmCBCy
6qpM/x0tk0lwSIpfAwJmHfUCtVWjy3yGSDrB3varWrmq8jAyOYHYmIUB/wbF58MQ
NNeur4RxXW5pbV0C0yrE6Likrzubfssz/aKT5/wTRVSA25D+6AiaIH3ZpUd2R1CX
yrrbgO7mxJju6MGipa/A6wna7Iay61AkRCCsnQED2pD93TVnsc5d3xxsgc1KAc4R
wLk5x2ZkgTAoqpa+G0Hi470EKHyc56deN1akleyxKNFxJcsdezbXqefftoMada/m
Dn7XHhnzxKAuHSEAoEzZRn8f8Supfeow5RNV5rGNELFK3+BqBfjj+8IG1eyTjA3m
U/aJ1hwWuYm6bYVSWqAWWRLVX/7lyCwYMU1DY0rlTyl4/Zt3Q1js2JsIdz+JlYQP
PxR0OWmOayblkTMvCA/pPy1pGANVXUO2w8OZ4jb3AzCWbUQkueUAMTWvsK3eR/fF
l4d9uj+lmTkJh8ERicjmMieOAo9uQXOc15au4BE0dv4gYAuX+Iq4oeW9sKY5oXBJ
lw865HSryk/aYBZsH94WxbqaSN8KCyTq+9fNMdAT0P071IHbPQurEngc/K3CVlJD
4UEe5AzccSRX/1V4F8gh5WagKn0sQ0KyD0h8cJdL154DpLUgUrq5Zv7yH6gsOVRy
HLPqV1kxSS4t7NPcyHzNlXImOnTeWbv51ZXeGGTuCt0MKiROP/coOtDK6MbhxDEN
/Mc3sfSgZ7b7L/tSAo5V0z49356GRmVou66HhYH39t3vsk1BNi1kh7ZTDJ1Jv9id
fGcLjq6jJXKJuOPtjF1/jVw0TD+CJwk5Xq0/611tpV1h4+nya04e4HPaisVKHS7t
JNuvu3opr1WF5uOi9tFVA2LsGh/fkZ3PLoZ+thQh16gE1Z7MeOXfjHroysyh86BI
8fed+HI4kPzsgZSFGLRKkeqcaqdRUR1Uzr829g+GszQPoL4u9N4Jrh7Gj34Xo0bp
4/ROZWT2MEx4ewubLONQmCOAVtRP7ln8cUNt3VMeI3fQXhdBkgoabEWHifwJc/p2
QmmRvOKxihOQg9Khj1zrd9jpLqsI1vD/DZoHw+f9hRJC0gI++ylnmyL8QQDA6PKm
xz2OmZgHJFFHct1eGBjXFR/HJgeY9ER9mPb+Iqa4yce5DC86bmXbrcUkja2W3vcO
OauRE3jUctVL4Yo3gp85cfDR2zpKhhCnEKOepR9YJnaL67RbEZoWUOGNcm1fqaV0
16y3vZY+V9/UnE4p/Xe6/t3Rzt+AFnd9XOiC5NH1eCTpFv3Ky5kjb2NE1fONq8Cz
pWWkZEDq8a9J4wgN1x7beHHW5eSRb3hnekpzJ6UlWiA0BRFkHpy/rpawnazn5l23
9leCzO8Xz8kXyhG++CPS+KDlJsZ/1kKmMQG/W0kPbzgeVbjL/0WlTDYUdDu6g965
YpeeNmvD30rzD9iIdz49WzLvbDd0zKa5kOwINSoM6Pt5C0FQN/PMabObSDz7+M1N
/7+XEHnE+CcaPU/JU69miE51LCS2sDW/srGooS2XNcsCx/n6XvUTmDWzpMrryrd8
643D6xUIs0NM6NGZJiMM9LyHCNgP0Y2ZS03zrjEKCjYladzbjeHfnGWVTUoUDT0+
VabOChmO0u+994EOA7EgZd1SMuJRPanFvJsvISklaOYrSVaUeBe5XJtqa1ShlHzu
KHWyFVWIk+Bj+W1DsP3VmsdrzFbNY5axe5bQ/NAG0RYjDJTvTTFLFGOnTaOi7wD7
25gRtJniYVUPijvi0H5nmkX3yZs7IL4+5y2cixS2zKzVwGwch98fzmbON5NsPAHf
EFpGwxzHAaDN77uMoKpC00raPD3CsdzRvKxREpjOTwz5lhrd1BEqdJnJCekMTu7z
wvXk91lZE4wmsSU0lKxVcc9EP33mFA3GYJJJOdMSehDhAt/m5+BFag1TSaIsHl8Y
tFgSE2Frgqdv4j/yT1YPHSi2DLEeAgjUB7rtXakxBFKcyN4OImRyj2gNagh+J7Ev
GYzV7HPC2p9q156F9yiLPFJyuQS9hQkOr6/yrfq5tJMWe7f1P/JvVmi4PV3d/9Mz
Qh0xPEDFveIeIpY+bSaQurRlwZknprz/8XcMZG+R4sJQmhGxCf7MTAHDRpXQVzK+
1h0BhS5Lb1OjhWtc7BhjUjQd2HPPaW5+jFvl0qIGoZFB3l4TYwZeXXnNDcSv5hmg
b8ByR+VGJ7Jks52L+kj1lcNH2O0X5IwCWZzMWdnKUK58vFQSGKeHFlV86Sw8Occb
3pYs2IAYIP/fLZ/JttI5M0sXhzMex7DETruzyhzHxlh6A6Xb1TdRvb+hWLxMlENi
LaBbpNolZthAFe9A2CuzPjUC0YNx5IL7s3da0Tq622FKBOYUyWdxupYw27Z6yRyf
FVn8PqEpsUUE5B3AaH1UB0NFwqmVmy/HVHDS7kz3lmgpDN0caUIsr0K8jEioFPNM
U/SpEE6V0XYN8Gg3ag/N+syhD+W/rEQl8QZ3SGVVFn6HPPDcjYSIgnGSmBrFFl4i
X9eGmS9HYkkER+mTHiAI64wYbE6fPBRe+ZS+lHAbHZuaPKVDMu/AKgQzkQ4stEtS
vGotqmaQql2Z2sx+ZVXn02c8FcxtMUB6oK6WsTJs0l65a2NohKx4P1ti86HTFeBQ
QdhbnwZ1Ioh6D88UYngKmfhoH3GrRVnCOgFh+mpl9ts4LQpPBDYkHpJAQBNPE0fQ
Rs7KU4X+65IVi4djifFNUFXUl2ilNaZ899asYCN0cWnjEAXUZ9WMTUSifctRHhbh
ZqtXwP/SsriGnEVn0iUHpeRcINtgbbZicsCZFrfFySOHBdxsk8qrjOuW1wNAWATt
yH/pzfG8XMoWQEnwvDSddACqn0zKCzq1wMVieyMNgIRQmKlnoaGTq5dxcRXpGFd4
x31N6d6NHHaGZOYlYFbnVp40vrTYwmTdT2/nS7bj/SkuXGGiY1ziTgXneheGbeoF
fIKHZ5wm1QD1022B7WAkGyxGSzB5GqhS0kKGFnjxfiqoFjp2/KYs7jeNpH9D7Cm2
7643+XyBf9/623SJeWFeMKoNt6V6JzGkiEFCEmv3wYYVhXx3sD+7LiDSC5xWZTf7
/si5fXx1S9cr+T8sta98nZCLEcXhQrCY9/M8HDmNXPka99tW6OkTW6gG8jCAJ1Hj
MwnTupDgBGKwd7jNWjn8aAELeB6jDU9Cl6VHW/xsXb/RETFCFtviohpsqFxCSyoh
+BDVFAeAWeGostiH3h+QwlASocobifJLJtqtwpmJZ19BHi8JmC1c0eyqxR8LHNAL
pkiwW064AY7OORXn55EIInW/N5ylb3psW8PBRmzXtU3e90Ufq1hi8N0qOF97GnVQ
N8EAs//aPE9ceyEgOqzgWXaperGqylEK4WE3kwarUuDFzVLrKzZ169pzixNzlLOZ
UsYODWs9pHN4Vy2HGX7k0zLN+ToV7YH+uceuH5rNgq51Zj8Nd4Y80QssryTtN6jr
3+D/VYM5Qli0uqi4/St6tiMT83L2e0pxmylmSo4ICf7WmkPQLh7yOn0kAK2lJJ/W
Q5W/FJjOHoX4puc9T0fOg2aMfptFNu5KHpobb7LtumCEL6DtjIgQR3P1tMNiSmFW
77ihHcoPsKZqXPslxQRG5L2TBZOYz++Ao9wOLylZqSbZLfLpo1wlWbSlAYk7lTbW
YwMVvDycH1kYCE+WZgJpVc2hx184j9lO3CKLKv/AABaEbCmetR/awVAMvgjnDRyG
p/VpMDgALt0LbSNxolxwa/c2UUblW0H8vT+Kp6+I/wj0LZFFxjU1WgHF01uUdYSe
z6OotI0tupy2wdZPv7wjl3s5N47FyG8NImjP0E13JTPEs/cZj+UdwkiLkR3209qm
D5WDeXCYyRJRktxHWuYFMmFt7PIiNlw6C0mskIUP9eKyvv7WdWfm4shosT4AV8sC
Iat3Ssj6r76EumQRBlUwfF33/6W1UPYzT/PD0yuv2lDgGdkRDS8HJo1odIs2ViLm
Ja/JUJyfGn09bXgTGpL3AT8VaZVLjgQP5NRUKraFrUaD2hjUrJ4NoNckmDAr/y51
stztQ2PJgw4iwDL/q172owxHhVfVp+0thTo7PWt3xdOfhenT4hiWFrQ8BXRW9OU9
DUg0xWIyVRFRwLht87LEWtPxzkgVvO+11XRGl9IvXoqmLWCyiDOhmldxavAQpoBT
c7cdpN4sArU1yre5Ty4r/a4zWr7VsiWfcRKJ3UTc/wSrIBy4TnvdIa6aredaBmGk
DfRnwkYpi8XfabtVX/iGU66XPkUaA2vgTmLps47c5Rq155B420SLmwJheclJydSC
UoqE6NGAMO3v9ckftSDG4QA2/wTSFNqUakAtsNPC5cmn6HQ5CY7QXzVivNgGXpGF
e4wCPtJ4xUaV8iBQjDFJdBda0WceKDi43ieVQOlHVm5InS7NrcfpxF8ojWfhZuB9
o7qCdrJVCf6jeEn1kJHQ+RlQ61qL6xXcHf45CHfsGQ/yWP1hE0hAnIOPS9XdyZ3W
7aDxaqEY9YQy2ADmbie2XIwYAAJtYhK4IEGMffmsb30a7xGyw1pc4LrJHCg23g97
oU/aUf+9e6A1awa1qf7aGQsc5AuN0MCPGgVPlYAvJAK8GFrsGi+tDoB89k/OjdPn
IN+OblgAEaTIw8DxGUvjykDqQm1SD177t4qJxvbHdvwVSNYZ88mvRxFfhPX7w+pU
ZywLI0lJVJQI2OorjV/4JROyAWYeeKSsydTrejIDsoKDxPc7l2WCDXNYb7fLYjAT
0UYdGL0ZESpqWOpjQ/JRGALwWdCSuoFiF7UEWJKd0QWHLnp6vm43ZwEraR5rJL2s
7WcIxHDjB7WIWTrKgCaRohefjiIUSGsWepOlQRv8VwuH/lzw7OcPmG7G75cOOPTg
QyTRmAvOu/YYjDD3sZ+hLmswovUP1fCGEZSW2y9EU0LVziy0ll3MfO+ZTcpynscG
ohPglHO5P4YlPZJDDcsZxXIOiWZEH4L8u5Bc3SA7EbyRYvVBzrxOQAh5U8c3zeHQ
M4dHa70ba5QmmVYgL7ZCStkNS49dm+MEs0O9tN6kBvmwL3aAvQfJoOTRP8tuAmbo
df297h2AYAlU3iiK5HZpL5s9XDhT/p6EuC02Y0P7vETBU6d/sTvems7B3JF89UuJ
7Cb7PE+D7yH45h0/N29R4hfZMNstqp/6cPkiqwCj8l66CDEae/HE0WCCfMfOAuk0
b2HVtZfZJBJP3TaEb00pEaKkqBTu0cT1LMQg3d4Qbgvsn+msaj7LsVGYVQ9ZNU+4
1nPpJseMGcvNm4p+AUxn/nzDih2Kda23PVfSAo9IEjQpuqnj/U2oKRTQBEtO32MA
gy2Gr8W8UyhKD9jdkFagCuSjAQv/0mdSKjBoxsB9fhSAbiv7tSX3h+5r9Xa7PisL
FPnbmD6hRMMVmf9SqqKpQUcfPSuwcqr7We9iaLn9/jrfsC3Ou2UNf5vRyqgSIHFD
cDTpR5AGXlwZnEfJkSWl8QJsLVg3lxdec0sIrvzwmGzWn2dGSTdbCsaJ+mkbQvN+
/mf0AUW2y8pCyf8G1jd/csYWcaSxXJNaiRdhylcGIbXpx+1vyaSsubdZv9Bf0pzx
X2jS1JK5JRHavcmS0SSotkWfHTbJG9lhejzNar8XX3hRNcgCf6xzlnUGm83kimEb
72V5IZGllTS+/gNeqmNti00SMxKEkxWYE9r21O+K5GYmkJ+waNGnKUlAMWoRZ8xZ
SkFqCejgYZkT/14KTuDC6Q1OmmkwqkGIa2t8LxTr9dUIPSKOc0p6hrx8onWzPnK6
zRo2ela+g20Tc57Qi3DfXrimYSiYxhIQScCzy91vdAL88K1MchpSU/58HjK87yb8
HaAbiG6M4b1KlvnvPRJWh3IiO0CukTMq09LG0Nl2f3sardCIVfIgjDdALR0VPZ5S
V6h+HEQFPCp6VwxLQ0eGFhJ+rEXyVOVw3AE5QXyXJA8xBVGwlziWL5SzfPG9YWv1
iglw8NyYoPec9lWn1LgFhuTvP0yS2VhjbEgGMc8ICQuvmERHJjODFeuyBtACooXi
jl95oAfmzITIrkYgEMDK9MJgRvcg7PBRbO29YSppPh+XklOohwI0NZINd9bn+GlE
G3Bsq0nXugZ4bGF5jEICajxRWiR0wuUzPBCKx+ONwJm8tz97BQuRaE6Ko7aUEnXB
A+tCH2oSjGfQwEOQTNr4ojV91DpVgOL7ezA7w/FrRvPrkDNE66s4+TApBmn4JNEl
s5vDXGSoVVJ5dPDV2kGVSK2jUi6imzQ/9+qelRcp41OrX1hF65RKm3VBjFHEXn/C
tisiWrYa6yPhw2YJceN2F0oJIlLDwW/ITOYFdySMC4keQ4SYL4WbPNd5m7ZWwuws
8FzrLDhacerCXup+XDIOI9KFB0/SNeuqbTSSkGDFdvIPM6ipJhsoeeyxGbERJQrL
P90lotvlmxuCzJt3nI+zt/Wg75oY+rAMPASzfR5fXHs8uUqDy6vDpZ559gPk0Ygo
/KwVk2DGgQJ24xucPJ4mX8whDaf1VTXJUPHVhLZfEpxm51W6Bj7qmzwaY2iROuLE
d1fVurUVVv8bwvjsZq4JgwCNIEHNKtbW1KvgLBYxbXqo+ZyfwA6uM30ONdLrQZFj
tVXCIcHcMvfCyXWjh50DNU6uHAyxbBWwMEDLt1IFWbG5A/n5C5Tf6QR68LQj8o+V
JwUr0lOVqgZ5DcaOCuCnIs/vX6FhMd8FjgT4JIpspTFSLz1h4AyH3li4H8U62+ab
Q07a8OhwAlIQ43d2n1Gn8JjuWR//V6RkPaAC30a7UxGWryuDUjMzABq2pF2eGmUV
VbUu7tdpULIa308Z2T3AJjxfNR9KjY+GUG9m7eJzBZNbdjQ22hYESY63KwKflJon
mc4jp4GLwTwH1V87E0PNKGmcu/39J4OjWRt9lV95dWZtjGhQR7oJuxsFGhRGzAwx
GjgWnam4xz4pMARH+cv1CksQmO1sFK7CX4JXZyq2iEudzBqPJhhpOTyDfY0U2pJb
rbuAk2D61205b3t83K38BS8GpcPjmonmPj/r0dAA+iFD1CmkJJvDVJ/0D5jVWN5t
dPuHvly68502JXOx+Tu3JdTAFskgCHiBfsSXnba6ba9LESBGsq/kWNp33SiM31dz
PjfhYh66VSINtNU8tY5LnG1HBrUf4WZW1iFMDXTxC9Ti6iR4mIWZgyBcR4X4KUtp
3wWXU8/Ipyly5DTwxon5xN9fvstQOvI2Aq4UtMebbYQ05izqTmBLLIpeCC8nkI3e
+6lBAZDwzQYVlC5Ne0sg3dn0m1i2dxEaxQkvkWjKBTUBTvfZlhIfmdaGbrB8/J49
OxpYjzTAWI3ZBaw3xFUHH44kkCsHXjcLEqeunMF7to7RAvqlwqzKm8b2K5OOS0EL
4JhRX7xR6YoyzxNNSTCW4+cm7+SCuXA2Zqvs825uflXs2eV5xiga8E5/W3irwLrq
r5V+Kz0SxxgNZbAj/k0WZil9X0GZaK64QQ73auVRLKwrZgUhtSdoZAt6GhVgJOCI
xPpqPQhcfGiRHMnCDWIxFaCeS6S5y/FDmGQqZ9c5TSD5yPSTHev4Xl/eva6aJylF
NEB/L/Mm55wuCUhGgiOgbfpLSlFXWi8j0AvciOdYl29fUBN4xYFc5sH37DMFnsYb
z3E4MInlSa1XCtukdm9Y32Vgi1B0cI4zrtJ6iyX2shfyz4g3b3pK22A4/Fc3VQiZ
DQbg084rJ1X4vrN+rp+pwvwJnu8HkTT3OnvKMUgrd8LSatWlPxtdcLIPAxiiGrqX
5KAih34UvhNFuCM41JVLvk/T0Hvfg3EbXqYL8nd+AbWyQQmlTlIxvze+pzDdY9u5
6ZMOsaUCb26z9atSZMCcxrbt8BTe5jB2gAJsXAgqkUVJbJtIQL8nWHxEMdxJKqPv
lyQkAQO9TPAUM5jR0+vg8lMmub7vURQUOMAZEfU4ZoHU/mqS4q4PCaCYOBZDOLdX
2F6N2pFdPQxruqQFyCbOyvSj3zhZPbffQpiHIgbFmw3YGcxvpsVKSROfcVs0cyxt
GFr1JSDgnA76PF2QHk+dJ8bO+fFm3TreUjeNDj0yaQrTOaASizoKHqNFwt/VSxlT
+4WU1g6kbWi5FL5Djo03Wl/Uh4nyS/KohkaMUyV8fkRWmDEZJqXsfAZJ71lyb1Ir
Mhu6wchZPkkaG0b9ZpGDTTnJzCuSfPyDvaMwOUGw7AHSiob0yEwA4rbAclxVECDy
+iLY17H2peBl4dfySz+5wh2gbx6SbdGbBIY+N7PKM6CsKCDJdWbkJm2WvZX1y/NF
rL3fgEiN7QIYUoPMnSt39Jhlz9JY4mXpU5omtT3Jt7da+iFqQdOzeV0yfV82u0ca
W9S33qlXdup9frd/WK9Ilc7K84hWaWxCA1ZyaYVomzarupnQQHC54FRGJqmSWcs1
cWzixB2IoDivlyx3CZZtq+keZReJnB34QFOwd27bbhk0Se+Dj57qln+Wl+kJHQMR
dAO0YMEiuWCPr7Q6RWdvCbbiKUV4S02S8XjFjm9Q8KOYkMbO2FueG3ip6TiwJzX7
hACKAjbCLLdEOHHUBlmddxksIIEmAw3UjKFTvfYuEO0WhC1s8W7mgfFd1p4tRJhr
bxJ2TZEA/eEtkTHQzFsm6+VBwpO7mFl29R7Cg9SDZgRqaUSmNKJ1LEfIJiOBVzAP
CL6XQoFeFGJCVXPrrWtr7KbBLWOHoAHUTs3/Sz2LdfuKyuW/RvK/5IWcFfE44r9O
ybu35ZMDyRBUClL2EXiv9y6twTzdfu+DrXA99lfNgal+AkeDTPVYIrSmi7nSbP3A
5EsesQon7bqK0R6Wjgg1QFUdUAWMeD++WqwLtN3MkZuuX5RBXNZBMpZJpawiSHLS
uQsDuh+RRtNmw9cZomPatls2s4xJoEwK8ukFkS1jrtfYW3SGDM8e2ueL4EWvEyCF
wnUcA5w0QO7v+7WebxIpXAowGu+VVEFc9EMt0gUWmTMqDVexam0pjZiW74alkdJY
1mbziwx1xWgi8i1UtnY6K5EtE2/owV57b76qWsG6MJJXRQAcl2ey2jgPyHBVpjqj
ZHVA2IUTW4+qJPIh5VIgosXjRHSyOCcuFQ+0uX0TyTrSr0i4G5ODHgr8neB84kGG
09pdowwQ6DU/fsT2S/6sBLG8IKPCQm/9sUrgLb4kkfJjQhy4xCjZF6+psgmyKVBr
j6fd9mblvSklbMU9hC7Rn2lo+h7a7V2MSFEwL8SYUAdCc+D/1BqMSovT16bO6ok5
w0YcRKaNTV/4TyCr/UntoeNKSnFGhZ/2D+SSdViZyy/2dByWKAX5hKQ0wpGa3Ay9
a8r1mKUJB/sxafG7d2iUU0xu2I+21LLKm+aOO64dmB+wF4W/J/fG8RaqEVEliYgD
H1UKOBKR2uJh7WdVh0urOePqPic6YsMyN9eqWx1huS4pDAQJMUhSwn20eCUIQ1rB
PSlVva/qJneoKe9ygWPmbrjS8NqzTK3tw9xeKg8Q+hHYa5vwD1kvOKHe5u7rwG4Z
/YxrHWe+LD8uyrxI3zKAtOY7FwmT7mQ/oA4ACZEd7VFvkVRM5vU90QA2c7X++0fJ
FGtDPxqcXr5c+eHM9Q+btC2iqH37pyl+fWrG8IUrXk23m8pNLlZdplqWmlaBQnnZ
YeescYv7DJ+VZF7USdfRpLQYabNUprIeVNowbguD/pCqL71QsHuFDUc4O5v73p3I
nbPn6GVoO2z1JxAhGVOsan4uUNO7BbYUwVou2e/hJw6gH1mPJ0sj1FHDad7NCzIZ
2FaycgxkR4iuGKy8nYEDMtsAQ1UY/cE4YBABT0cvZxjFhVF9zo8ZWCG8KF7MOmLC
QUydc9135iV2XyeQh9UGBaeWgVTlXfSuOiyZnwAaX3el1CUQSLB19LuP1585HfqN
s+ZlWudNgDKrqimT5FB5Sm0z3+v/XkZwqmhhJq0imJuy20jOnH6jd1eNRjaE3l9L
`protect END_PROTECTED
