`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8fXRpWC0dnL+As/zcsolVbBp9T1TT4LvgJn1IyO8eXlMnBtu90Pi2ic8SS9ERJ5z
LOUOts1pNGbuxZRuQcGZUGfNE7m7YDzqIFuc6AOBErchY3+cKEjrlxShYeJ3R1lO
JGGVBJlzqGtBuLFItTD0VwtS7qIqwREkF1gC5gW9i2mpZQVEYwCOuNE/TRpM7Jm1
4lmDgCDNZLevTwo6Wmj6OuAbJHowAHyEj2N5FSvMEQMctWhrvlmerCaGVOcN7qAR
qEoKjFehdT46leAtljyF5oueZ+gDcEy36NGVjOOBVp4SlKV17aOFvGSlggNslzez
qWgzGzfya6Dy6CpPLHruFpaGujze00aNOJ2ji2AgK4uZnVuKZ/5v2e1cFCnphfWf
zoWUjDvJISRI9gNq2QTQFKmu8owOtvJTaYIZxP7nQ5UoDNG3uf6j1C7eKfcfYZyU
Pukcxt99T09zQ+2SBGZs/w91yoKzjCydKuaisCq5Dez00iz5hQmWeGd6RzrUuwdI
Ded/woj/GBT+d4frmyiN8SSzj5YI3pSpnibEVral8GI=
`protect END_PROTECTED
