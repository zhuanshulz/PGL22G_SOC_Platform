`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g9aFe2vhrKIOAs/PczLGwyQLoZ4YgYftNMMKroFx9gYTw+PEh4u0Lw6Da1FXbGBq
M7mMzwnR7tJkAoiwNCHIwfypBQ+GAbA5lhuJTyJcx8/eGTw1em1ALF8EQEm50bWo
uXw4dXFsaDaXQp+S8vxeqvLEGCrJ/4M4KAKDZcG1b+1xSxkneYdhq1LZz6Wm4wx9
dM8yeVryfDRuRuOLuPHrbsjtTfSSj1eqYf7Yd8bij5QERemFnTkNW0tU1XPDBEn+
9Zbb8A3aLRyUxJH2FBJlfrWCu5uteaP3BIwTAkN8bXY+DicP/1oc1I17bGrRphNc
pEhN1cLzwRplBCzuwadaQWKu2oWgSijK+LtAYLe+kx9B9KlgIY71aOBPCH9DgIpS
dWG7KdQXGnwPWtc85InoruZSciPyfwKUYrF/AIhKJ/x5rCTtPa4aCFb5SYKCoh4f
+mT73y1wmy/+2bCCt4HHsLE+Vk2I3sBhN1rIX+rJ58Gc/SSiczVoW98UEU5LV9Me
fekhzJm6MG1VhfVJ5J6DrLNRzJMbDAahMtQTLHpIAvEBHseYc3G5Iy+tk63ZNh3E
eNHWp2NCwnrgZiZIqWmr3oW4rsv0dRTWbixU4UGN4xY0WnR741jEhOGMT5Ny10Lk
cJV6ycDVKZcsPqoY6dJ8X4cJLeNZDNHsar/VqW3LT+ycEP9E5VumiFCE8hrkHj1w
EJ3KMgVPlXakKg5Md+p/Eysok8L09a4o5qZ/asrqXszE8S+ox4Wn7wKFIakUIHdj
5PatD8jDP8e8FoMx9uQY4dBBnybRyEeG+ZJSA6TAErHSWdiyFmwzO8Lxq53t9D2J
/lDMY6FM6vGEx6C6kVQOGEHCBU9beCXqDM+MFF1yupf3lEFRYQP3dIykbCqRoQSu
kZ+UFd8XqSRZlG/GemulBoEWoDts16Dv8l6sh9oFHeWS2fTbSUyL7p15dVJzwo/7
A0mMW/7GcUq+x1AXlqq/p+6rR1jqfZpJO8hndbsKNZBte1S3KDnCq2a1+AXaCCOU
DTS7SVTBpjOwbYEXzvVGMgs8jwwVquaYv0l1/xg/wkCDOxdPR3fUQ7//lgwdYede
EojbrKUhSwuhTIAR7tt2LvHhxNsMO66s2LuewzxslCn1VJN1wtRNT+XXBWJRexQ+
4OWKTHkcRZZwP/TILFLnrUOeTWMbRppp2A3ONmH0D5WH3ScZT7429sFGDBI37yHk
avfb2FIjtiZPErfxqLvDHZBwtC/BJ/RptF/gfLRd8rzcV5QnfLST0hvjJSXeFwKB
oqw1lawNUY6tJD2DZaj6MZ8/kbfBB7tYDkW0J39orzRnbrSuQZcTXWEOwdbaFU7X
he/JanJV0H0gyABn8EhPSI9d2iGyPTpNYIjdEmNL4PPsId2O0ujO8KfiNCtWI6Y5
cUgEeGcH4maCEV/iEyXqH4lSajoH6jkA1RlY1nLEJTJNyO4b41NTnVez7XXdLxQb
VhYr9qOyDq2eqYirqAYjkfOB1YZpRBbOZpJuxhgyJzlSN7KbIua7/pnVdqvXHIKU
fNO0bIOeF/9A8DWh/0Jwsh4oMvnib+7779jqu9Q0aMjtmEed2W2yonZStDCRxikV
VnUfzDuYIPFyOd67BW5u4LcOs8Q5SKRu3Sexby9GmT6u6q3g1ua8ORICjpe5GiTE
hyNSGQULEILwWf8XHsG6plWBJ42ACHVbzsrBtIRKGB1slikMirRIEkb/mrkQiA+B
H8biYgzBRhiwZezDRU6+wv8yVWRm/EERn0Wq6RC14I4UcEi+AWkWo8OQ2j0Lu+sS
Z/GLReAGqcszNnXXkhRR2wyNhkwjwz32nLwNhI//zvaJ9wm5haBNE3YZlgjCxj/8
OSNBk7wHGm0RuHPWCOGu5dJ0L5OJrRAhCjxXCJGvICPUK/jJz4KmBiUMIf+gi0kF
KPITFA9iAsFasDKDldxoFEFUBFxHOVPQIjX/dVuGL159xJDUozqo8oMGtQVQb5ZC
Wo2M/W79Ss+VbfKJ7e1G7wNtuHIN8NwYA+dWuwahu3Us9XPKfSrRYc6Iid6p51MV
a3moKBdENxDrv2YErX73mg/aKuilm2mM9+sqvpZRjJRjjbCO5FR/0gI87nKrsYXM
a0EDzaKePoqsZ1/aO970nPcGmP6oGC/z6/422T57kSM4Pvsh+LT3PoP0NAPe8XHk
DhwA22RCQoyJk9wp50qBNgKV4gKM2GSOUXrezhzCc1OQa/Slo/OAVrccmmj9f3Jb
Tbe8WeceGb+HVj3Wp3ad1mZohGDs8SyrhNBDOHfKz7/hONhwHlUGFHxRYGk9UCNU
Y9+WGEeOrbXi/XzHQBDjrcZuZwkGyRn6Cic1PutEew1ManWVNbW0PeJ0FZ1lfmEY
`protect END_PROTECTED
