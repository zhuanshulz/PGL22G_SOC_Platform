`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ak4+pZbqiZxZH4bn6DVf9flUPqed6E/RsmcnmmadCPEySqJg7XoDEDB4HlDr+Fe+
09qZeY1ViMc1r0q6Hpo/cTcgcSNNX5q7sJ/Q8hIplx4Cf6cUxAQHaZnTJ6+ac0Rx
c5pepd/0OAZkicyY4WTKYzQOtbec+qFlJzCxima5pXJ1s9BnnP48IDY9EeX8MHxM
b3yDRAKz8c7kg6VPFNIw0hfPM1S8clRiZb6RrElXwlZ9TCZqU7Y6Om765bWJTT3e
+V17+PEKetF5f8oOjuduTfiev1oCcTSdUtJoBu2SpvpsBqCPe3/1pMLddvAw8t8h
B8do7lHTsfJcQQdEXDA6TUXD0oYmpGfgIouLvZPZWs3UDciYiiFw2xS6gfCeEjzE
dHXhyhH6hgY2s1PIe69Pb58ysSyMact5Xd352SVSafB6GsKwJOmWpmHGQq1abh9j
jF3oz2SWSKAmYJoTzDoEy1xevfnYFMGokTOKyJjwmZU65QODxmi2Wbgqb5uxFjlo
uwK2oorEdwk0dZPyD9PMHX8ROdDrd7377UkngCS+1vWGa0/l8ocxmq+dLI9ACrU0
xmByTqUMcWTW2R5WXpqf1A==
`protect END_PROTECTED
