`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d4dW2Oro1E3CCa8HoGBqsC+c5bA4nvAgh4HKYu4QNaWiU9KZFarqwHaj77+cFPpr
r4VXY820ecIH7TeDmEeJgoPdRKnBEXQQGm099Zzf5W90bRHWc0OyM8S8Vc0vaqge
5xd1RT1AkW4CclwbQdXArV8YKnksOKfTvewBdCwil8WnzoK52FvTvyALWq3VI2lG
Bj1UFqMe9myTjZU5yjBPWNFD9gOviPgdltmmMf+p9U8BJRPS5w8eEQzBk8F8W15A
j0tcJbntzY+/FNMPdIYhBGi9IRdQuEtq6JIecMgSYKhhrISIoyAQ5o8YugA4gBs2
h8/f2GzVOJv0AxrsBzHAmmGZ4VTa89DgavcSgTluLaa7eVtUOcG4VlsDxEF7elkp
2Bpou2BuQkwgLER+zYzWpm28yV9LNQqWCwzM9ChQvkZayHK+Jx+8MGoX/YxzWVT/
V3HbcbylBUpT0Gx5lqjBYynoawrC4whhyDykUnOkcCeHDWQyX9hIw2eAUUDw7rhm
+xv4zogUhHnzHhbtGv9pWsaoBN9g1zIoJBlfT7iDm7edsKi1ZRMYx35RbMsJkr/7
FwWki5nCsKWkYX4OhLYFEC1aMLCcz0xvqYq9itnSMZpAxVj5ypA94itNyrQtmJAv
MosY5yknzQ6ZqsL5ZP9lEMz7Q3yb63RGfjY9QE0sXLOejqLEsPWOrgHdRt95kKm7
5ecIS93Z5vw2rphLFPZ/nzTfM80NuK0jTqSsF/a74xa0TUOiofXBD9P1KuYPsGnJ
7aTGLb9FDqfV41SaOTXZHA==
`protect END_PROTECTED
