`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O71BOw0i88KIGSTlyB5+N85pw/F5VHe8D2hc/nme0wNlt2UiyKlXCoScnbvUP6fp
i7EsMP+9zY9Jt9q4BbGumvhIlBVIAuidx7DtBhx70MnyI2cNRqejdUVshHM2FUef
u3eDTpSfvb8gpdxEAYBlF2p5ivtODsQ4YHgWRwCiXq8W9hlihXTu8QOk6e5pZOiP
wSIE6ld+0fp74U8PBCLlks1+sN0350eIAxgAmiI7qmJmuvJhtX96NbryoauXMLEk
N9i0/9EgSNjhsnlCqbCTS4suwTVEQWbm+jR5HxD8Yk66g268q7VsIHCzyzLC/csi
DgEeHINl8eeiCosruBlH1uQISmuxsChgyFytn3mGw20Tue0KO6tSmKLSY496aDPA
/xB2MAcH2capFzOg6cQb9IVyyQ7KsQaA/P16Y4PzNuqnrNP0o1JYmdlat3WR7EqT
HftNY8LMWlC+en1KTKfLzKZ8q7D0c/yjLRzYEL6LCFPs+g03vnFlKWk9nl2GDmUe
DdQHLyC/hwCydC/TrILIXc244AZWuM8GxcPccqvwQb+vky28civw2qWz8vYbYPSH
kZQDGBIN8rt5bvTAeNYrefwEl/rgd6x8d4Z+ngULga84XlLhv4J2w9cee14ilQUg
Jf2R+3i1//vjFg6FqwWVsAJwzs0spPHKWJjmF3gWWBbqt3cMZ8UoZcdDGiueWCui
RwjoSEIru0XeQqMmk/3C6RXAEs1Kn15sc9WRFD3QahRMooTyRQSQh7MshNyP0N1Z
yeUtf6FqwN2+1TibmQWhCHjyNfqQlcXC4oa7/HLt0ggXp+Ko7xC3b8Dm0Y5WVnlb
pw55mDEv4HZmagiVEOI8fStqw5u6VORDhdz2Tn9jg3xwfpcexcGlKxHocqAiHCwD
r/QKFgH2H7uLI7iccLysuZmcHJ/6sFvUN4/4vKEGZe735wf+JoRa96zMf5yno7Fo
0xVeFqlevGD3a3wJElgmBvJvonY37m+iTpQjPxdMewT46ZCBqoUlcO2d+JVEKGPE
uG8+wld8RyB8/J9kryS1q46CJ+s0lalG0zin9dFSLTQzq/T9BcnilmCiNEL9tVuk
`protect END_PROTECTED
