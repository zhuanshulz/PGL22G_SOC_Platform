`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/vtRVZIDj/No0AOQWeFe6ZID9VxefcVLmn08IirycvBtOE4DBZgDw+zy8IIipJJt
qvP6EdxGiTRPTPTjSj4n82C8kWRLwdonteC40etCeAHkTLvi38k6gOhJLDCekNWs
B9UZF+1PpmME8fjguVoN01YOBIBDWaLewQOrfwipCNDjyTC+R6ln9rLcuNCg7b6C
AxKgdvaPJvLbB/88HCb4zhAaOqvut53aFAaeFH1GZMQIxAWkOLYIBpRmdvP7JLNi
ILEbsy4cn2du7W5ri8VScjcuU919DHphxsBT8EdClVUR1otE9v8TtkSPiry+OmWM
ZWw8ziGhBv6VF1wYbIMNSA9jONoo9J6RhYUEQZW/8oeGtwJFAD/9z+dtWo+LSLJv
aU1O1k8PP0/LSFeb/D5monx2O097DWdPqkoQhxRu9b+aeQOd9uZSWBVtOsuArJsC
iuC7RAPzWjYhRmuWp6VgB4kvsXKStjGUjT37CE89Fvdrmxz38Jg9rLtHQYyauq6V
+RRwf4gG8HoftYA0fFNYt/kerWmTb9cl3r4I23gyCBr/0SAGt220ZxPMudINICAy
v52NjT+WpVyrb4NVZnOpq5ITDy8rS+ZW42A5DrgJYKuxlhsXiR4zwHNZlqfebSzo
BXfw/rrCScgLxYVm67MBKecX32ZTzCiz0rbBmIvG3nwaFiGfnw+0uG5X9rHGF0ig
6/hFRhB7bxRkuSNvD00K0oRugJbSgP+BgT/6p5iTf87961tiyaL1r2LFb4kOE1vr
PW7J6/rvXsemxFgKBPwbXvj/6DVy9fpdg+bFIKOPvqYZl0eeURxvncVM+y6/1DeU
Y60wh7q+zXW3gcpH/gtVvCAt9y22a8DyGd7vnnJWLuMNmNoMIl33J167Zxy2wnSy
oa0/8zgs9/XlnkRVGcLcDCmJ0/N7ha0279nLU2KJX/kSk0FB+I214WloYa2boBIJ
QDK6iFzfFpPeAOLZUahEoxBnvD3WyHi4r4n7YB7Hd6vfBqTpCYRC+C+1bLV/U9HY
R5wvKkcLQNeRlBha/CT/01BB/3zUTuANedwdkB0FVwy/wNOgsjXwq7t4zUPA9mNV
IfG4DtSDeT6212ACIBRSi/G8kH/ULwe4s09S7o4ctlA3TjQ87kghvayyCh1LhtHr
E2l8sVKjNeIHEzXiOfeiU9u/rnNzgIHRFAudKL4QbbQDbe7KyzqfgH705OlhfCbl
Yo8KIJCc6tEFa5QOTz7s1TiiO2BXu9dzIvyaVmzH4CDF/LRFcyJzgxFQ79Nt4c+g
XKIe2KVVV46ElhYr4HFmWjh2EcSK6Epqd7JmNhngENod69yKjudmjG/QKMAUGhd6
7W2HT2wlCVRUZuPeVUQ9RMQYGEqxAGS4k4/r19YhLUR6ku/029GLnqMQ5/F70XSz
2Aowkj4jGL8qtIrYOKOlGI/HvtjgqmlrjsO1Mgxk0ynjcqfRjRUtOMdkhdcYDfKP
v8IQkz3fQoe0qhyY1KFHL4EVMtrV/iTQRbA+xOKAKRPqOjCkgiWMkceyOjHu5lKo
yHZseBO6AHZObfPgANnodEp+ne4iL28pCf30AhZfV9YxefyCI+BUv1HGEutVpuEu
COabLSS2TrxkVF0NoBbuIJda2puqtwCeeyRRRtJ6pHOiLahr07oaLln1V4Mk2Jgw
kl4bM4/49kV3iE7lcL58MPxg6GDueqjh7GRTzzcm2ZpPz38a1X08YQSnWlikW4OA
5mDW8dX85gLJxZrWOKlBV9rGC4MIvLadnfkPZhi03mpGkQ8WD1BWERvGaEOB/y/e
J9ZfmstiwqdDXI2/U1aJrtcLP8i8deVNfXbR1n3A+FwjbWheHcfzFM2MqdMQL08Y
ApBRYcJTpZk7ZMYfIH0qb7Gi/+wyUc/z6P7UwnXYtIt5LUQExGyXyMB+u8nFVwhU
wP00vs195O0kObPMdIOGcgr9ElbwflAS4qrYT1Be2x/HzdU+6uuwIgbQnCCkuqvu
aCyJjk5mQFE62A9LpsQXM9/9+oO+mOdcLd+ppYT5Etu4RMmU3hRJaKdQAcvm7c3H
x/OikfaQb1EHnJjJPstkbaxCtT7DYNhTA0aaUzUIhs3hKerTyVx99KtFG1s+bROy
/JPZQ2ev2XQQHdA/hvSBCYO0VDBxfWNGVM9udt67I7ZGEuzcG7XuGiUCjjUE2anY
vVL5yfBOBERX9j17uBs7tWZa6orrkDa/1V/BKgbIQVMjaiCoRn1I69r9DrNHvlpP
VhJI8YbaXokFjzffHYgujGiXyv6jeLM+PnR1yXTPG+9YeglB26uVAdBhX09DNaID
ZcM5cBItEtITLVnB4L/kY/f9WIglJBpOwjEe4qrXjPJPVgiJOy1eEwXIBeaKhmN/
zu+LYjQRlqiCZKapFFkDDh1yd+lZ34FgJ5ILYDqYJTvGw6qhbsaZYKTxAmqgKEiX
7heQxFhIm26RBHYkr/N1M/7rSjh7kyfPbUK+RSQWunmrHt5esLTki0jJL0XV/Gza
Kwhi5zBoFLphIZot/PgIduW9lo1ejGfdRK0JYOQoE0cEtaciSArjWKD1ap596UN9
XylvOrQTT1nYHDOckk/uoBDYJBibv80Pq4ZonWrALmTC2aBf0Hkbnl+EetOcizLH
pcVa4iRqCoOVJbmftBeATXe9ugS399fxxk2JARo8oCajqOHPTOcEZNksTJeyqyFI
h0qxpqdXS1Qp5wjWWlAxPRLvstZvs3JEEAMxvJlwnYVPInvXmT0uEt2u17lqdgPv
QqHQpQ7PmFV5ZmguWPoKmC1HDvXFotf1sJQzUy/dUFPP/VEsVXkE48rkTEH7ZIW8
wgplYm0/3wsvvwMn9QVonJQQUy1Jsxc2sZVd9SVO35vkGcI5+g6Yhum74pylg93T
DuAw9CHgJ/O5FTOpGDhKSFeYehmmfj0ypKvpmGJ5PDI5YkiKe95PIugnyFX5lTNo
PhXuWyEeNisnCp9NBWQdZ+OFe8St0oI8BglxXfS5PVFqoO5oSgwhpFr6/+4YeRvm
7xUQy9oUlmLiKl07bVCv/8c3H/V9KMl1wwPojSO3AD2MYz3O0IYqLUU7VBisGV0J
VbGzAKb+YCF2eVqMvFC35AsG+Lr18w9oSQ370vkKfkI0xjfp+9vRlhtLsDy53ZzO
2FWofJv2cJwGZVJgbI04fM/MIYT89dGsutqOcoXYVfg5M4tlBM5ufKdzZ3qTZ4Vq
+OREBx3GygbNYwcjv4Ei4xcDmodd7nIqJ5JS+TZ/ZbprQv578oyMm32UBA2M4o8r
mTX6gzzyRUKRz9AMxc+ogN9mnbLphMzfmzZN5LN8Ujmrg4Tmw/4luRMRdAGo3UDb
i80Cy4P7F4JK7Iyx1IxfNY2X9cPUJZhk60S7dE4koDq1MM0A8uvMnFoH86SNsoDi
7E9PpgGf4WS5Fu/LPqoqMjmxiZRfV4P2t25Z0eXnJUgHmB6VLoYn5fRnnlGI2/W7
kpkzfrXGoV+fk92lFRDsMJ8BZNBqoY+pjfi0OsfdXViKr7+Wt4yYOEQimVgDdnJH
oMWxNANOPWqQM7CB8GT8m9NmDvngh6YiKv12ShY8RkSQX/4mzgL17HP6ReRntn9G
dyXlHT7lAXCerIl0ZG+OJpw3vOt0xFya/PSjWJgVQIR9uBCj72tatX8MdUCt23qD
TJu61V6s2PWgvPKsKFvKRITMNUQr8Bdbix18yc6DtJd9IOUxeR4Fttkri/3YYKWj
6yczCoLFgE9gB4n8VtoqRP9uETIg8Y99/TX8IeCn7V8sVMyOR7TBty8qF9O48njm
ZLBXwaGqj0EtZw5qOF0UPHHbKa6ogzOCCgI48LN1lpR9ILWm12TmnTHaTGZMOJZf
+sNvmxhW0vsu+skSx/MRngvyFEUHfp0KjvUus6cCqY0ne/yvpBzAsEBTops+gChk
hZFZCSBSr2ZWE5N5NTLHU+z4gg3qvVLTUa2B49NdKrzIfnEdGubZeiZOvvbp8YXx
/P894bbsTmZuCi/6OW1/xKxesV4MnPR+cV3Xi6zG1rQ0rgeTRuEd640VAhQrHT/3
gMVr4dw+mmblNMZ8TsnQWSOj0Byr4H+A5aATGaNiapaPhgMOcAJYIkGj6/2gmwlq
X6H9zXofjCH50hEXo4xHFtqbCkRamIaqqNYl0P7B5/eC90Q3T4NbSisHPZnSCbBP
sttA3rqC/tlzUSVexQZK9BTD3/PljB0y9dZWwRqWwLJTyDZzyPieYVtpHZxJHV0A
NigtZUOrWk1inVsROexo/yaL6KemcL5j6TFdo096+6W7itWRQw5G60wDdD8lQZVW
hFUpTZgFH+wmn05xG3lFBxguTJxlpVo5YWSNBsi5u+HmykytGcnuGkw9qOV8I8t/
GWTtyPNmWjGIahYEg71WHdmu10ZVLBuazpyFFm8PJOlhrAt90SC5IvYF5yhJR3se
W5WTApmOiqmqQgQiI4nORlrDwL6mSwAdT7S83Vo1pUEAQqbAO8fAVhEippnczcvu
RE0BLfktd90IivF6iHW1Hf7+w8LuBdLenIxuE8if7kb5aq3ifl1Nx4uTf4GiqTY8
19fyoOwrOOtMdw32Woc8CRJmlWstMnyLRm+7s67vUWAVEe/TfN5TJ5eRAoOqNSTU
3ewVpdbcOmDeVJ1s1U+MX9HHQ52eSyuu8R2103P11UQBLgfkoAO58EhpUmHY6op6
ibVipOfrr8Zo1gvBJaDR441UH2tqN52ggk9YbloxHdIQj3gvqSVaY4JnV19Po1iD
yijNP+WhKf3Keeui556JtsyfDBKZYFdqnNcTgAh1kDMGvcpo/bXLl77A8r50yhad
DW3Nfg6Xj0L9AjVxX++mMRUDR6g+821RNCb6dq35ripfsLoPp3iAVTMCOiS6Ymix
lgNRCMcB+ELzL7ahumRYP4qK/HeVePSfCK22+ELAqt9TZkGO6GP41eUq9twzlJqz
dV5anMJWWO6+yyXd4KUXAyKXpEupZg9msXU5dL11Ft+jjlho1aJogFFmQTNzof7I
VctgTbyNe+qZnfRjoDXh3i0WKuhasWb/hird1WSO9hXOdrVg2hi5ThtqpAWT7QOl
mk5mcnMgTaP0dx6jTINEnm7TGp4AFPm/7rCqqRZJWuYKUsoHHjfW79hJDCgUsTpq
pbF9G+nz5R6x3XZoe5mXPy114EXzyNE+/3Yh6Fdz60HBwpLmgK7HyoSSnWQM4g6f
ZV3Sw/FXHAo2auFT3PAfrv8FWGzbkAOmjNCkj61oxt9eTEG2NxlGwsbZrso1sTme
PioC9ngj5rp7kLm22rCN5GzY24W2wXN0Ir5Plr/qgmgjJ6XdUAELiP4Jg32xIX4j
xs8SdHHiM7UqykftEmxn3yXLRTAa8CsJShAci8Va3hLNKKWT9ao8Cpib/iQZja/3
ET01lR+zyzbXfUhBN9SxAvYiqBLgw2rN+L2ox5Sl/CF2tzPc+DiATHvhXicW0d0m
Kv8wdcCqq6gXJR4VEzM/oeWO0qekc22JFf8EBHtb4B5yY6Pq5uYIeqdXw6+2xjX3
dSpdGk0jPn3QvZ4RgvxKJFbfP6u6/ihWhjXz2PFQHVaIor7jYabsoFxJ9tevSF2H
+MIDwZB6bf4+zOgGJaOL5aUZRgmk4HIthFQcN9zkQadnD9QxSGSuydgAxnvS8OkJ
RnGCnQEyQScHepTkTlHt7He2HbrDDdFzR6rERdeoBXY1ozOz4zSIFwRtD5VWRYry
75htI3smgAhMwK6AZsoNmVmntjEzGSLWNaE5d/m9cxauKjbrgncrCWTNefUPwO8a
UmIJOs4tEqusshBTuJqY7FJ3CvxgPkdlnJy87SrtgLCW9CVHETf59OGA/v94mVRn
trQPC1UlMAG4+PmF/qoDG9W16AeIJMtbbVeNpmbxF2IQcHjbOHpwz93AyDmns+sP
bOkl56HUfU6Rxhil4ymw7nq31Xu8n3ydV1HfE33vHJWALOvO4CzHhFtObtKSgP+r
47CmViXJttqrEqtZb1wm0ZMCdykDtkg5NyZWcdSO8u1mJg6NAHDhlNR2jIsCMuAo
a73dRBzzW/1DDmLRHDiRPcsnqRjbxt7NpU79rI7Ysqe4XkBdBTOYxNQi01uEy40J
qTKgYMQowyoMe+OkB2LEfpoovAs60pwLFMTib7kj3ouo2l8+iWqVEVNRnmJB1d9O
MpDe0m5RNOpQpTUgNOEbosjWjZZDKKmY7QVXdHjJSoP15m5PqnvmPFJmgrGE7GPy
LUL/PdnM/2nYUhCLsEHpdS40IYKXSKQ6SgzmgV4GeT9btq2zCn3xK8uG5YyISixp
Pw0jiME1kmRoBjym+ItJxxN8GBtgyN8w9JZVjki+rcd9SuupLS+5YtCcmsc/+046
v0RatfKgdwnRZWKOMQ916nvBNaBp9cUBCe78nqKJyVhquije7LOTVlkiezvkGi/t
Ysv+TNoTbBilMVwR+CTNXmdQMyJHW6LWC99y29Y/7K70e81uIgNe0qJgzsyKEQyH
6p5W1qQ2ayHYRzKuWgzT39tVOeZgZAYDBTZv/SPI215W/VxGItpJgmhppXKSvWpq
PHYhaB1duWXjV72sh2cbUcV+ZqisN8zmZvYUQSzfwfwOep1zYApQ4ESPaFlsPVyj
fQIdIptAFkXVSlN+p2pefOcQxOMmdIGVzpiPt6yEyIml3uNWmW+u17odM9sgZs24
gxHn/NP8ttbMc/MXni+xpyhS+qFtK4yTaXsujHPJwyZ7nPllMDIUlRdRPLEq+NTh
Bfoz2JTgPJB2AFEy0q8/mG8CjMNZMWugWhMc4ZXvAjz0NTpiGpkfAnpx4qduSRzH
wNvLSkscad9up7f64UIo/CXSMTQd3IQLp9/SNXTAhBVP23e0SM239Vnf/+Cr/rXC
t0wLD88yTdH4yZNbcpbmI34JgMBW8yJszyg98TkaF/N1ejlBJ7UT5Css0H25EfFc
xYZ2w28A1wAI2eHl6/4z48vweAZSxiXSv51BjiThtYIzDUpWW750xz7n5uVhUGme
CCkQCWAKfW8bXXjqrHvJp5PuWEd9OTkdnTxXNhWrQAuPyqVEIYcbIrnNSveOOS7M
KnE1thjUHCjOhoxFFTet6u8l3O+lkJiVTv9V/4zeYXt7IRuddGvFwAglFWq/AG6W
wbUwhjv0VZ3pCJiQm1t7PHnk6lD45NAJbUl9CR8gwNsUH/63DFh4lA/ci8bP5cBI
5xqbp0+RiAwDZB1nuYbClKyUBYiAYxBErgCbHNNcZ4jRcDYJjICthF8hz7aaCZNz
ieBYzclDkPQij7CRu1bD5dBtCA8XcG0Mgw9vqJzFAaWiT+lY5e7EgmK0UOcobbuq
2lqIfXLWn4Jum/iCKeWMNSevyz1zrDrx4cEJwThyqrEQKiTD4MUEWY+3Dzbia3NA
BUOjJg7+KMWXpz3LPzuclM1VM21htkAMyo3m/OTC6LhFHc/U49E37XhB6dG3q/Sh
p9JZOZJuX6mZkfXpDTit5O2M/y4Y9WlqGdH4lKQYD3QANdnyWG6uqCQyjCO8USNF
aqd4BFIqjHFZGlpLin3G12qBMYf3/x/yAidTzuPn31E61lC9i5UWplrVYuyfq41j
tecn5Zo9WVXf+7sQvqWijc1i8PKqJeo/O3L9TEFdIy9qwJLuj7SDJcwZQOf8nHjY
FblN3/wjnWPl3+b7a1zg++25JM4r8WX0juSTPlrOVQsQzH/cCeSr9LszlrKuCRQt
+I9Kc8FQK0fbS/n0sqE7oeF9Ojae7wLvaTX6Pl9Qsd4AptFMI2/XVZZahK8OQEZW
QGRPIjSLrFhGyV2u8aQhWz/1JgFqrrWmEsaHm7/ibiKDAUDrucV0zxVs0iYWQ39c
u0Z/w//6V5qXN2JitJDtSvSHnJpZ1YaUQtjoWcW3P0fkhml2V/Jx1Zd+V7qKHpt5
7E26L1lUMkK5/7jkewCU1w8gZD8rMuIyWh0Y8zVCHAH4CvkX5C6gBxBc3gvwIfDs
5QScJsEIPwEElPhYIJ1UcqKoM8qDk18me0C6GxZ72GtCnpMMcYL0KY7hyEo1wSPO
cNbPn0sV+SJuRPZRPpxBcqn2UH3gltYYBGYi1pitSXAow8k4JjrHE733DkADnvjH
lZhhHYSW57NINXd+KJcMvInPa2ZquZp5jSdiOfSfCjA5PKHovt3oZ01Vf6pqIYnp
87necyg0ZEJHOUlfHVlKI+F6qOloN8+TR3ZzHh3isedRMOOyQvMjw5QT5l5BlXIX
E6k/rVKykyemE0urWVwxrcDUA+db+Td+CI0juL0/QOyHUS5KAE7+qfzEE4Jn1qe4
jcuYEnL4qBupcJ+4r9c/r9U11yjh28M3IFLm88LBWc+lCpEd2SW7Ol2Tw9bXR8CE
6F3bpOZQYSDE9cpo8LSxz9wHDcYMw0bISve/luLhpPMpPn9ZNH2kxu8DbbEr8Jxo
eufrDWsr70XaiJTm9GPRDgFs45q5Buox4N56up8R/d0jIfIcNlBTMoaEUu51dgkL
Q7+4MRVb/eExlaavKhYIhDVPe+FRF58UKOcF64S3r72H1MpGZchhTBN2YO02krIZ
Xa9vJev3chONZvUrnajrcJjWThQ0QCQV6i74QyMIGRd8CsVXryN5whVgG6JJt9LB
VXcjFrPBOQ6LoAYZNWs527hwG2dcnZ3OsxoODmTTJiPPkxCvs4v9DP83Mihg7rH0
rFS8uYV1ngZBR3hHcVP71ZyGgpNg4EmpYOHp9+aigrNHbnZZeODby9vzpwvDctQ3
w/dK59DENlBCrV4AZ+Inv029YxDViSQHUfico8ElRr2JgJEdczXx5XmoAyn3wxje
MLtIgCi757vK+oKEHqM7Z5yeewXl2scPX0kJxPXwfBbQXbbvFl8inSpAyxUTTtw7
ZAojmAf+BxhFGsPK9TN3sybSI1ZhiVgOx85uoB2DoVDmrbb7f1pYpadtNyPITEvJ
iiY41V7to0jA6FiViIsjpVMvqdPp/v+mYk/zgIOGYLode7eEW+qJ/Dpl9OjWkGpF
U/C6UsMgig/LnaFRUHz3QvUeLyNE9bRr9homKSljsBK0/L6G0wUG/u+tPM8MdNRg
VjFAPjXSDJz960OpgQ+jJh2FQRCmQp1zgy2YWP5B77WCCbr5mkQteCSB/L1n2kZ5
Wt0YxVRVNr63N+W2T5vynfYsyJcEVYCrJ0zCu/PQpHvWwN6buiAxgQGV9m8oMbnD
4QihBkds9Ri3fs+knjBKpKZdjeDYiDmclDaZF3dhKycTkBij2XS16NCDtJvcPKsX
XFbk2CQA7pbusTfuNHiS6wIPtYgGS4BAGk6T3BDwOXmIpmAarI1vAnpk4vrFmpva
JOkHGZcZnEQZ1oz5xe00AZH7PTGXrV85CivA5/t3BztTfAytIkWyerNojWFT28FI
IdKtguHvzNpQfMQc51AIHQtHBfNXqIX0Of21EFpxOzYmZI6AtsgfUapAnfoiAQGq
zB0qZslSbNLYGuL0qnDgOWX2Qo4QYKAdiKo0x0+y/Op6fOF1IJV0ciCbmNIiGx2M
4IXi0GWtx/KjbYqFDlsD5jzC8CNrs1JnrHlw+eZ5N1WWfhUhJivwZJOyy6Q5LMgu
hjyYHl0a41Qz+ahbIIBXg5Zzp2ZhPRcxArw4/48mXYIwaj6lOZik5WU/IcvckXJt
kky01oLuvBhCZ77H1j8Uv56TIuLeTKs21tdL/zBWUvliW7rpp2SGZhg05guanTqY
E6Vs2hL+a8lyQZOv+F0+qkUb2UiXcfB04rFN5eJz0UdZgMkwIdalFLXe31GqJPav
Cyz+UIsqueLvm0DG+Yta+scxh0T8cTK/oiAQ2/nYlffBSTc2/U9VXHFV0NqjoH/2
ik6tKMVeHAwCNE23tYbgsTdasVJV5E8WKFY8VH1H1be9W6P8KZIbjQsmNO9r3B9U
/yyHCtyyDH+jyceW9g2vhPHPN/5JJ7+wlAESTGuWfB8DyFLduP4W6X6qZN6EF7BY
Pp4xUiCKXs7Mpo3LLG8SzqDvbNWzXnsc1slSy04m7jcEAk79amxxrdTDHCSc1oAx
hdCRrr5fElEY4NtMOc2ethUc/aIqCN6/CV8fjPss0y/sHSD6Zf6uYgkurTApl30p
54EeEvLAaw8cQJRN+zk8+IszWzq2I7Ap/sDSjXfDxmpsKIc2CKSuX0GzLlnf1xHz
ny2fAAVTjdVlPi0K2qaW05wLmhmh0YUCdrJVuy0ewdSJ9Wbmy7paCsotp/0FmLRh
MVxoU51+k91kqCW5XdMm3GvVn1zoO9qtjMsDz4gdLleyhLwFrEFT5FxlIs40Njgd
m6mKmAzg+9G4NpCsf6h6/6f3Vwr0f2kO5Idb3PDq6OpjnmlmZHGT3MuK1L38EEQu
zEzeJkuBPrJREL+vt0EtdzeKhJYdhjyPYXehECKOxVawqq/UYMES+GmY6zC8xJ/Y
gmb1xGElTQ06p2KlpcYhdQzyFheDkTTGBzZ9aQNXHEYg95Q7PLr/Gn6P6CxDzGf1
BEj9gs+Achmr43/lkfxR+XK7dBMmKPvHj9OwT5raF/HVQl+ZPRc+eb8K3j8zXhlq
lF3sHPF7L1/v3WlWo++ZtrudgfuvKRW7N4hu8Q4VXAJDg0AlSCgqXWD2pVcgNHx3
aeBF6qb5AUEHF4hjrCHUtHOuE3LReG2oM4MX73yezIt1uA4ayZygnC+jy00M2Xr8
CUQEaprXI0JkwV1rlZjLaughX18CdnJEhr/2C7AEjQpEGIu6fY07HQilYrHOAyfA
W1IlUxcg8uW4JCPXhmEwxKE9e2q6tsWBJK30j3Hh9beu8JuFcQkAF+iOs3T5g/Gq
dmbhc9aApuHDicrpRw13kJDfzL53l72+wlyiIwTcoUi1cyAYZFvrIDfUENZuOFZY
PQldjI0fpRf9ZYnnRTtZ9E+zwOm4q2Fz3uvLEQGvk9/+j3e11gyKUNYQC0Cl9ifv
4kd/yUMjAgOD86GUuiTNd95Oq6gtegxDD/qK7Sh344K4MPb23yUcZetKw1pfESD8
K25li9i6Q8WJUgvD2wQMgccnsVsN3sinXiKrAjmthyBRW558zGISOJxAfx/pehW3
f8bZGm1crVF10I1otafCD5fOfuQbStUzl/l2YMSz7X3s3dGMnBsDJZ0SzP9x/71c
myMZ9udjj1eVDn0MMF0z8jXRaoGLNnqpdj9nCR4MVfkfqRUd7n+gEBIfdoKcaK0h
onTDjLoCiir6j17W7xZ+cPeQ0Hj2OlnCsKgQ6wfk0fCl17PJMabAcQbpBKK/Yhqk
L0JnG9FvYOqK7+VBx0PLL1tzAQ7+rHjbgO2lStZX94QDiKB61AmAOgyZYl8XoB0P
IKS7J2WzP1+T5cNJHk98XvvDX5WBtRHe3/fQ9ungV2KFX95qVV18W41EdH4s/UFt
8ed4qtFTo2TjDKczSTIDd/E+1i18UgVrNLqzzILWFFYQJ51AAl7gWek8TNeEkdec
2MG8qXRcpMjtmaSSjykW6bGLJdByj6A1tyyVjtOgIMx65DvsllEomwkFnYRBLMsL
FX29YwdYQV5OrF083K4QzweTYn2LBNzaIS90fR0LSA45nGNVwRwszOAMB28gxZmm
T/vtazcKf7sfemNghF46RAR84i/wQF7ZWI7FfGDlF5QpNANELpKjUgmlBJ659APU
cD+u7KsYU6cXpydQ09jFN2qlAjIc0qxv3Gqtkmja+JTPfhRufHZzIIfYcZPGxmdb
CbJ6JQN/z34VTxo0XraK0i11JBJeB2Cqgb3nm9JL3sETyqZpCqP5hqHiEv3++KDP
xnWq6Rzxo4VeDtOlUQmtP2J4UScSWqtZthi2DIxm0Cc3KcpQ0S8Gb7RWEzSdvzFs
+KNW33Mg/L4rz2chKBQOXC02jRq2BtzA54L6d5NFD2+a7jrOPlokBcPHvOhApCAL
bs3jWOebGXlfoXjIoLS/OYWnJAflTR+fflFjokkObT7sIUUIHBZI7myu3FVpyWf2
bjquiwfuYCXJ/2+6lBC+O9CDmhnFl/JMB+q4WbWC7hDrVCFSckwRlLBHd2ZeMWv6
J+8l2hIiFqXaUKpwIN2xZg7tPoOJEP0OEXR9aicS0erh7i/NSY+rqTYu3f2fFHAI
GJgP3/WabvFUyO9zuy31970y24YEVfbXZy/MFz2dQAPmJJil/2vF8OkaQ0/rRM+f
QUpA+n25/0PymrArwSqOtvdBNPJfQkFJ+FiND2xKTQemd3qyeTeLmaJQsZklajnI
gPEaRp0ad74CF0PVBsZx25PPufDVYVe9ksWEwTVQS5tjtSywqup8d2yv9pEO/mbG
iZiEZLo0fhCywm+AQRezmOCTwDkpw5oPYuq6ICrxifL+YypktDs15Xerw2zu6qvs
0uCB+lEi8vpvUK4URfO6w9I647zUsvWEwlW6EuQ7lpa79l4u4dllgn0couc6L+Lk
fOu79RTN+KWvZHPFXxGCLMTLkfzvnJqFdZMY2bZFJlo++FSNu7UZ7sv8EnP4o1+C
Ag1Wo+Bqswyb00dsZGUvzId/osHJbvMZBWSznfdAJdcjEtF/7IPPKqB+7Ku5cbmv
k1a5LNaZRwtr/SUuTZIlU6cIPrtHe5pszEXcH7s1JbRNtxYfk6A+C7Ft8UB8LNSd
h51rWzCpY5MNtMV0Jq/tOw==
`protect END_PROTECTED
