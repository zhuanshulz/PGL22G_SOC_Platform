`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JehUIJnozz4f3AGknNgxoW+5PLxe1s9j8TMIXV1vC9+CXjSetDV+ivT0Cx6XFyfy
Z3AlRkauTvkuIzNgCXUNvdPFxjvhdXKwyrTB79wCQt/9IEkse/8U6GbhR/AouX49
qkRAcL+4HXJzodGsBTB6QoU/sNq15e5Rn/v2T2MZ4Xe1udbjnv8OZ0GxVN8Z6v9+
fiWOlICgr4Y2/e8anrAy2lpdctdu+ikVPNK7h2MNOBM7td3LkrI1tLHLZ7U/0OID
fIAPmQBVvj7BtXxBycUpEV7GvoejSUMxIyN6yoFWi3J33Kukq7T/Kg80hc7ivfrA
cA1d0joUXvKO1GEPojPg/w==
`protect END_PROTECTED
