`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o+24uwPRvn70Zi9jwFmFmAoSihULux/pk7b5fyHfVCT7gnx/SXYfDPkloetea5R+
BGOHw3nQ+ws1GjXxSpsZrQBEnVuNTRm+NIyUqHrglutULnjiUcT4o0M3pKEu83uL
VIAs2zPd0iOQ5o3eBDLY06A3Jd5D7PzYt5izf8RO3LSjw/DBc+ZRQeB41BLe4O0h
hxldYLOPJKcCy1UqpT73NwS/W/CtniFfbXFjCliixZTwzhz+YvjsXJPDj4Mq5Paq
FBW42cYlNR/il3RXCFBtac1V6h37Yphrc8pHrdqWYjqSm+jJHd7KlH2oUbE/fsdC
OZtvt8ftW4TfWX8Wic2nCf3jqQGUmmkYvM8qyuqlhSNH4kzig4/wb6oyexE1ZOsa
9bV/VKs+0fNJ9Mehxbuj4ujJHxK9MNU159GeM890eeMJWlTqXNEyk5c1ZJ7NyMQZ
H39QEg5UDQs+SwGpePWx1VG08i/6o0pWc1l5YnhkFyf9fytfTOWoXOk0A+CWAeiG
1BjS04OUi31h2+/m1AGtbsiLEWdTi1UwQNQ/jJZh47VF7OALnNV4d9nDOczsxcgM
Rbc84cUrHVlqbC2zmWwdkIhoCxZgriDewpRt/AoS3AIwxguArF3D8z0MjhRa/WfX
l4aHKiJKTvxGxZ4KSCLiEISVxZCUmz5jDH/Ft5Aywhi+LiYCDkOCZXtjHrFO9UEo
q3BM4fhbxh3fdkTuTEGHn78BviM0tJjXAle0SIKM1m0W167zmu8tiTSnWtYVCvrG
YgmWYimrg6LNgrxc6UhFonKsZBSFP1UU10gR+aS2z4LrDYLxifKkv1airy6ICzd+
mF7LZ2iZ4VS9YEwYJ/Jzrdd5lQi4ikKhbFhIf21Q6VzQtPthzViUFv8q8PF96P2b
EJFTVGcAhfqNJScTGnI9n3UG6zn2B2w71YgUd+a99K9jssKUOiK/6kIU4vxaGD+T
JCgojIp3OMRoqabrEnVxYBHmpFobQr6lx/ze1EaPOAxLPq7pdL+ZLalcO/Jv8sTv
wMzBaitaMRUP/4vECNG12yU11GKhUUM6BjT9g+C1iLw61QSkyEPjG5eMZevDzPcM
zf1QQSL86T+wEbavJMhVufrZif5HecgSMFPbi0BaI9D7Ji2VPDw9bi+jCKu38jFa
D98l2/mwfjqWsKn7gJsM0kRUdtaHplHSRHdwT5iKfyddIxpD8oPjYCyA4dO+3L6I
70//7SSSgsMNJRm2b9Edof4fKoxU7EIKcAWUinp4kdUN2fWzGGkKjPs94z3sO4BV
kRXeIhoAkR7ZrDez0zX+VQewNAshI8tS4ulytISPwwLTE+jMnc72Afe8GcLApRCH
8bdEbvcBqkiIKhAPaDsmjjHLxZ1nmREDDk0CizCZMZZPNPSTNQ+eln1LMtAq+NLL
blI+eZvfgycRNfx/kpRyKYYQoxUK0I/kaAwRwirAr1ezHJqVcLlDuUakrl5l11Q4
yBGpbtJqyFkflrhd+KH5t4hpG+bLIIswZ7ItNk5BNp9kGITVUvF2qi+2P4dDndBv
4v19Hmd31lHSUvwe7jkBQV8/mYeprt0DYtWR8kqR6POfb9Uluin3PpuWeM91XwJ7
C+gxGjT9MAbYLU15IZCFM/LOzdTf7DSZGT2oC4H5M01AopRPpDHtEBe7G5OT6/X3
cpGe/YSRv275PrFeWDp6A4CuHWRvJsBqbVtCHkqmu2v2/wPRZjBexenIXpMqND1B
ZbDTkIRQzX44DbdwmKInKb1WV74BtTnOo8rAoCZawdM36yfhESaFfKLiSajojMld
q3ghErW3XKv5RTwSHJObBOb1FEUEwepAHgPmDTDRSjhmQibei5HFdEpUusr0cMMd
yaQ+IIEVolorbe39/roAwOEtHULPgR8I7hIccvAb9blTZtn9YFQmteHx0bk+Mkux
de4nfk3RzClgo5RqNFSeQif3MN3AASwh213WXGYKBMeDPCjlnSkmQnpiyobaw7Ce
LNCVvhlbA9FhLRm8G3Zlype5WBme6daoQ1T1e2k5yFdDVrMHw6rEe5aTfNhLbrl7
roXC9X4xws6u4vnVzrOslsIK+w43q8IWe+dPTKSNMlftuiCsXUYN2Rl9TJBHu2FU
/O+CnOxpTZ9F9vcIoe4na9xIb3VKytT5TVBjj4JQQwK0lrB/9t1Vgi9cQTBY3BUP
599KOFAXsC7687q50hwlWb32E6lR+B+LRKvD8X3hk78=
`protect END_PROTECTED
