`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qqRVcI5VPE8Yt9sZJmHmvLnQzUcgAwcJFpbXZw/cHq+lVvOHQBP+/Dsa7sjfVY+s
Zf0LukKkFNGHgxaZy/0HLN6az1qVCP7HFba8KXheu+qHYHHt9yy5C44VW/l3GU5+
MKvZNPzXxZ793IoptQwhrdKq9lMa7aSI9AsBrzpx5KtyiLIiCtFS9lQXfI2573Wb
OOELLx5Hw+Hc253OPB+iEcCBXdKwul4Xg64dr61205gMiFPDJVN21svX9Dh4+7dm
bnOfTG7hF0WRIGKT2bQPmaUu978BTiT0IGn4K78RQ0TAQS3gfvPDu9Rg2SEBZvkv
CyYgGzrNQFYIICgOWKTL/NuS+UAo7XGg7j5QMjLNJDclH1+mnKPu7XWfxNoJyEyj
vehKVCXBE+kVF+Q7x0rwJ7KebXEc8qLCNkgaE2dPwJrE37GDXEcr/QWeu3Osxr3J
NTcha5if9M/df3mmwHuU/zEozYN7GDRzAOrCl2vNg3RDALJ2eswYGW0GtSxbwG1W
8Z4/RUtfE/z+H6fuSx3cn+z0Oj5EWeoMP6+jgR7JtXlDTXVx3aBk6BjpjH2W1eVB
MZ+Gkbb02qRfz+PhgzKrra7d22IdIVYrfK/gpmqmh/ZAqUJEORIlSXUF9QtyHXUF
Cdt//h8pf65PAK4Bbx7+YUprFhg7ak+zni8/YmTxiC3tB6eYXF3uCRt3u6rSti5P
P0C7PKYQbVrDrDwKHJbdExw188bU3UVKWNns3i24SzpTk1GhoIiRfO7zGpQ0tWfv
mXRx4++rVQXE/UJffB6XmNu45Enzzpg5bK2il5fOoUWi9+RuxKADm9fz7Wd6UzFK
Mm4QHTgSjucWcwBF91Cgui3+V9gidgdABxtLS1LMcvxSpHnIZdgvwAyEUnZ71ANg
gr0SjPqgo9GAw+gJUwuZcbWdsCHQFD2ltZG8fWYDXr1mg9B82AJ76yDgSU6noutn
5kW8iK6SAWzzDHbxeXstR4ZKmY3SxIJUv5sRg8LjI/oNivOsYqq61O49cij6WEtg
O8VpVyU4SQo8mvUu1K8PMghhHCGwllYC/Lt8BHuSE5dwX6QL/E4TmOOTSG9YgT9Q
`protect END_PROTECTED
