`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
feIPd1UHp8U/8NhSD6XV0yldMDqe7Ienx4EnTAEkLfR5k9bbPaVIo2+7ozUpyKfV
g3OyhBcQ2GYdgwv6gA3XTWKwKh+hky4Hyg6k1WWAe8eG3owR9qAp81UtN1xMeDmh
J3xFivAjMpPVMRXizoKvo0eaVfU6gyrNay6ZBoW8u/I6lLVpa4j6Soho9+sDaMEA
6LUZ6UP3lzdA7bvpHMMXcYT0fRu6wHQSK3zWipt4mKgbQCU6wvbUTVUAUfI/TntX
6nPYq4Of7t7vYcmCeGZkmcoWUtM/ad+msPC1JtNHSrI=
`protect END_PROTECTED
