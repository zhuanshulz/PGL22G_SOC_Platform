`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KGOQeJofl9W+oHplMnSSyjjQAsNUWJ4XQpxQOuwFnGAEyObVSnJCUKy6y/TytXK8
Zf21KbF4rjNOON4ytq9Kqo9yxQaBgJpK83/EP1NesLegRNzvTAwwpEFFVP+bpxP5
u7RsJYReMAw/+MpuU9arH6BiAJj5lNjK5iaNfHYgx3n/jKbHD96uShpS2PKwN+zV
eIMpb2rmX5rTuXH17evjpKbX9urYdkOpGVO8yibsjZbKv8gDz05lUi9hQPFmHx9W
VLpZKBn+lvJGesbIn56C3n/75TAkrQOhELbylajLMFjlIThE1IVnZ82efLL9fJxy
0xly2iMVKPkm1hYD0gEFTZXG8Vzs2tkIIzNlH2otq0PbA7ULYB9/OSHMrdGSgPNL
Nn1Sr87M7v3HdhXMxLFg6nrNtebZAvsbHUaL+bzQ31u9nM45IYGWFxZXI335vY84
oZG7/XTsiBwsUIIzh+UqhSbrRGEp+ml++dcjn70Esv3HCTchAdB6cWqX+z+qybAT
olja9c5ioqIiTbhSx+qzzTiHI114JdGpKVbl2kiy6UMqv4uXFoOl96tyGi30CW0y
HoEWy8JfgURow4MdWdQV+wbiaYFtsQRgurx4FbT4lDtRQ1xb1KjwRsYFQYKALdjK
I8DMm22bN/kb45nu2lQTPxK2A+cV9WHTyWwUr0gJ/g8ru+i495Kl4El/UnzkaUcS
`protect END_PROTECTED
