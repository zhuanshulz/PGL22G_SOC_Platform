`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nQFWLLvdtEVjGoWxAdCR9J2bsYEgyxTT3E+G0Xd4Ggd79+O4hM9MQo07liyO8kNN
n29JQtFKMGM64WWLhg44TnWPQZBf6OlipIHK6GSqvE+OGc6uceH9xf782HKcNDcG
R05K4g62odO5/f9N95GMnMaxZyKswKjBOaY6QRTaa0twRnVfEOd0BO4QzQiUNdQL
5ndhEKBtrb4SGPNjyCzIFEMgPAJdXXEf0gpiUsBb1xU21TV+8QWdDuleuxYUXGFz
Br6hlzD1RuzDzxHRCnsNgHQL8RJwO4vZVHFoAEI9M55M67FpuvUHrXjsmGw3uCSS
pihuBjfMsMLP967kiO7Lft2oS/D9n8c/p27fdWy0IVFWWdFGOMBPbFW8jK92C7Dv
DbX48Hw7qRrqbZrOCsxYOr6UEYdERW3ZN4aDAw7TKR5vjP16lcXC2yAicrBMH/xB
+tq+rLc7RgfrnvF9gY10+gYzD5TAAh7qaUGms5uZ+FqHS++8drbHehrlgrMpQQYm
crtGmmsynAjiIIVBgL8BkSxjNYUNrxUSyqwI7OhOJTkP1hsANteDFpk2fJDIo+XK
nVjIDiDYFKwXBeXAzvKcMktMXSYoyxzaiP2a0zCtDyE//bEUByfinn4iiNEjtP6C
SFiBkf69zZuvfmSgJdnc7dQStlyqfViFCOzwULvjsniw7r9cl5UC0S3Ghaxq+ROU
NH6DhDbSD0kHr7B06cVEviFEpVPDSUYfD3MZYv2xomHNO7eQP/nzkStN2cQy+FR6
ghyI4H/AKGY0p5GWiMfsPdUs2qAiNiqhHqKrQc3Gk1frkj2g1bIuNBjMpSEow6SC
YcI8Y5Ol16S5N3y9PrwEZVL9eIgmFxFbYgaNBJ3RycrHGeBtBml+KD7qj+wT+pQw
rocJQyK0LCe+AdHSc3UVfIj3uJi6A7v5Yeop4qaZGBSlp9JsollqYilTW4uuPI9c
TwKO28jejMfBtkx1WlPjTSCLF7/W53SJB0eeNJuntM5bp7XW4Fjj998JnuHXWNN2
BR+s5nU3aU0LywJ0r4J0uxhCNum4x5QF0wv94bzAkO0sK70ErZ2YDPPvEnO6Nzk1
pPyx6S5yDlLl6vx7JutxO9s5YM5RtjKaP6wiJ8E+nSM+ftvfW8QFqTqHirnhcXOv
dZOoAtjEgrkVYgsWy8lmvk3UJe4hZxR/WLsZlcaRQRU8CvNdIgBQW0fkhfS7UCHg
6vQSxpJc7LnIxuJ1z9qmNZZ/6w6zRcMubkAK3/87ItuJtLkOwIPdc6EO+bLtTFPr
v64fElMV3cNl8GlVBxS9X2vC31ZMxvUuK/kdQBmcy4c1RTXKH1iLYFr0SlkvW6kS
y9vodzKmdHc8+hPgPFbokC+lWNKSkphDYLIw7EPiaQ1B1fQmFUAiR5n1DMilGK3C
KW3KBOz8B9FkoLGIGq1ruVYaYtSRhyXnySxxR1LnHBpD+gzaw0DqZZTTx34lzUN1
rYjVxt2C1o/bdGZqoa87GB7vjVbSzPkwQXSNiyQ8iliwGyYMG/js9KnA30emtb2+
W1aaFFGqNvpcVB4P8wZTuCDgio9U0LW8duDkVJUW5ip1sUrYQZjc1mDCy/lcZDf5
e/jvxRb/61tk2Ph/xGSIqqpRnaQnvEFxp5sVpbgPLQNbLeVUBAh6lbzdeHZg4UMF
V7AO0u95CJDKTRsATkdyjCxAKA4d6o50SnTfjeeBxF75eWWbD79WLDrCfG5Fzoev
+GkCGmzzCPCfFtSmxARHAqDxXC+KBUyohl5T6hrFKLQVt550NLNudP5xFEwJlFL2
cwl3MtI0BKPDIOF/h6NdWGZe1vn+SYRxNWHyyep/vzzvdoiu/xJk/N/RJika8oeX
lnAsdWhoyu3y+ag0LSXZxvayXszYe6EuB5bLNittJJ5rp/bwMuynsC/4uprnVc7j
VVAm9ELi92FCtlRJy7G9r5mQsTCaKWPsgOO6XuvSJyFAcru5gJWTBeXgHE0QiJFw
06GQWNjO5p2W5s4zWF06KXQN8nEAuaXFAGJBTDuxKobWx38W9MsT/N4XBmKpbq4Z
gwawPfqXF0yyQhKGxROFoQEsDj/Aa9clYQauEV/NYZtJjxOebAd6lQsNJSr/S8S7
S7Jb0EkQcaLrDdGeIFAKDiF1PmWR+XqYo83PxtE76gMyu57/sXofyYDJz4t7U2VS
JJf970S07ir/b8DlOrdjPO1OWDRImct0yVMwHHh9DfisZpTZASmoFWBlo+NrnD2o
uSbaJZw9ff/M0OO7pSkUpeh/P3xmg71xxrFSxfJ2zUqUj79Vlcvy4oraOdqkc+pO
2JA3Ph0WBpYcsUQpY6mc4WAB6fRV7Q8XthVFQh9xppMgoFkQTl6A7TpFQZ4d1AcU
1GRr9vCRtWvt7BisXhLkJ3D36GkjmIotMdmQHOY4e0/yBUEVy9IXthtJLIaneDdr
uHs4EcH4UBj5DE91TV0X8E2N9sc8cPzjYQlji7BkGWl08R7XgrEeO3gHMKMfZRxM
/mWzXuyPmpFWo0/zk5UOLn+yPKpyibLj9vFul/eAni9l4dQwTJSKfW2a9+zjubC6
DPHuXkL+PaJXlHoM+Q6znOGdIBw32N5K1Xvmk5fmMNkfQxkNntaBFlYHJu9KyROP
VI019IxdUlChvjRrJ8DA0C1njZsGsZPwfvopJKqpEHw0pUnoshg5lMT7EHiTeY4L
ytgQN5xTgePm7LYrzzq8lHg+0tdKOAkMAahI6w1ZA50OWCBFS7nYTNTVszn0Sjok
nStKXxobMirij0bt1gVhcts20QYN+88DEqPnfsi5MdlyF0YQFTqJb25sDRaIHZWD
fuVeQhZPcPzqVGSDML2KFq25NzifXmGr/E+5qFrtF2of5JmD9JSfK2meqFtVHodJ
WtU5Hx/NQs4iMbd8IjuvzqZUFKM0AUoLPDjZMtA2wQKuqZ0aoGZ0k2brRw03yqJn
qia4IGvo6PUTHYAT5yUHgnJRXdEFrGLAnGWA/FwnedI3T3tjeN2UH6mYZqNJ4Jq2
qSx78+Bi9ll7xKn6SSHCTn3BFuFLITN4YzCPCZvQFBLjn7O7m86WQVW/vRCk6t1u
BpJJevwtzBUDAKbuheGnY8P44vECagpQjPm5TgCBrUNEVXKkJcmX1h/HDCgdvc3B
qcMByNsyxE3InjYLDLZsgcYxnIIr83mprR5DthKU5djGwENuk/X996ZzHFLKIaLj
631qe83621AB15Orenf+fc4OAUaNtb5RQ2XCMqgGXLaKhS9Y8pfCx2s/2zEMD61F
6zuqwS6xFB3MxUgBNQiA9joYIA6IEGw3auBcj4Y+gJ8BXWKpHDEq1zZ6FsHvbM3O
FvWtXcFu7MBX8r7b2RMKi/TIV5Q+mkeVyfOujOrHCyGUzWPH8QKCMYFM46Tv7oOW
Z48v7AtI+XD6CgiIm4vnYswLkLZHarfcsEzKrHfmSbtMvH53xEjW4xrnmCfhNggh
3V0Exx8LPw41Ru1TuldWNdX+bE/vD5PQX4H9p49bn9Ja5M+VxLXngQxOrzmdW571
Gu9NDLI5Lhx9T2eBbTREluXz2+7UIJei+wAmK0Kw6TvlZt41OB2Xkl3hgIgFd4LI
XPBe0UVfQjAooAIrC/lTEqgVbI4eaNXvZbaeVE/ew/CbYHjOcL1Hm5BcXFYwlOfO
WNBJqwMg3RpPFJAxw1e7QQJF2cWejOH5t1rx5cRkJiSawij2JDR1JUgfNT3EfvRB
zE9aURkOILxS/sp+ZEETKH55Feek64gd3APy1LQW6bwzY53+lu7mCzE/7OkeL+MJ
CUBv/LS3SV8jFfjhL25ayfEBSX3J2eNhekvhF1zoImPonW9LU3myK4xML2XAaVGE
fPJxXMX92A40AfGsrAM0vJnOXdpC00i+bin5xKXZVDE8RSmBRkXF0J0wHYcYem3X
xnku+Tll+jfqLWS39I30D9nbc5ULR5swPvanD/Bd+BW8N7Wvy2lIdZ1DdVLGuTPb
Ma36PRkS6AOE9gXrCikh2fhGaeCTIRdUDhGJPhNzGTFiIE8+w1LZUmDhWjUFQeDz
AGsvOBFy2EF2DsiSAw70LALS21Y3zSsmvJbtJOV36IZ/rYozSvUvwPlhKo3t0zmm
OEYVpCUL9Wf7N3mRAvPyljfcaDeaeXEZvIcR6hiCEeS98PXBgrEqA/+Ok0hEQksU
ej8WvggzhNk6YZPKmnxlYR87lWJDt12VcouH9/sORxBs1j4TNeUDvR1IS2zReex7
QIKxNmjPufmsircqtUkP50uWYMyyxdPOLlM5dCAZHUNiPYUiai7fx+IIoRumfDjt
`protect END_PROTECTED
