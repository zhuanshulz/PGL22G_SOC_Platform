`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BbOPXcM0iBMuFoZIu52e9Bs83wNyK3CjJWNiBpBEa9yVs8r6ozDDO8B8QWYcYQ47
gopGJ5Ud12SA0imuKFKbVW5GWzqQuKJDXSIqlBzvVkRhsj5zJ/5OGXZ7FCP8jmJJ
9Qs+JUH+S2Nv5afnsuojAJ5DVm0z4C6XMPlUkR0Wv7wBwNvY3CKmfoI3xss5inzD
WHiZDcs/JAemV1mm+JGxyD6g1dvqOy0uchhwO3AmOlKdA4J93/KsjmZOC0v+vVx4
UXrA9ORU5EahVXjHUlNNJk4dVDVT1VSQD61bToofVw0VPCY8RtPEosF6fj0sTqSb
569plbVOnBeczN7ZssDt0gwZS2U4IyqKo+iihVazw2F2zblN9WBIP8ZGqZJAit3v
4H0vtRWUBUYCYD3c0tS5YHFTzBZbdVVss9YKyHQgQnJEN0ndcWF2Qplg68kV/gPy
CXdRGlRcIkPDY0Selr0gfRcbLC6KsiDovp0UDev3g21Z8ygzYakgff3BgXJ9njJy
AOZQOLT/GnHmfcfpRw35J1nEtpiFKoWJWWZwC/ki5lBdE9VOmAJkNgv1LQezCotP
WFHn4JonZtHLAVt8yYD79SQFFzfSO5Sghkzoyo1lKxYgI3tEH7uuKfzjXg84c07h
Bitv6639ddOIIiIB50gsOL2bwJzGhH1NV+/N1rh3lC+yjmHA/yBlvtFgsa8jwJma
cn1pA5IelNNl6x39Km5wVrXIrTTHZ84TvQPE5JllLOJ5h/ohWAcyOTn/pfdyR0RK
qXEgqlw9kJDVNLdQWz6cSHepZrC6Vjm9jJ3q0GkihkSW2RoMKm9MwMLfqXr4i3J6
VfEfD9U0RmgmVIr2JH3MgV3y2DDNXjcl74wFbiwOiO2q034fgkLytv3ykn+OIbvV
gZjEQ0+s8WKfy8Dy37ZxjQ8moTK3kMHpJXMAmNOb+ZsPw0gZVy+6TQJaVe11ak9x
feHb/n1uQHUSTumC2Qr/4vUCQflhMyXkpMovfdtfMYnQLrtfCvLajkFEYgijuwcF
Ojp/tv7bKUpZBO5hDVGNx08h8fBQ658aWsSWW7ZNLDqeyt4bb3Qbu0ncGL6rHPKq
w87M0nGHaB4qXMfcmt9sXg==
`protect END_PROTECTED
