`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XEOo4Rn8ItOW1ucvBSAQhOxh5xekt1g03183fRJ6g1cw/z8IeLwvurGrscTTxIpw
46r020qAG3NyUr0DSpD/arXJkT3yV219WhFiYPT9St8N/dq1+qyzsBdG08B/+9qd
JYTtDHhGCE/+pXi4rMaYjHtkrnTy1tvpYgdyEnIQQHo4O2gQDRM/apzVVROCo8l6
zzUZOmfqPULNGuZN9nK+yUL3OHTBdzBKYZp7Y5t0pu8DjIjC8QWvxAiJLoze9DKY
2VvbJBpEKn2r2yT3Mjmif6NvdYW875SSKl6Kpr3rAKQP/rW8hCNMPPEP5XDn9HrP
B8wrFsCxmY4xld0mclWCzIf106NJ/9vOnYH72BwQOcg5elmTODdGk3ACwtl+4LPf
PNl0qi6zC9S4IrEvwOhJieyUho83NXppBkoMUdMKSw4NCQkLx4MsvhYF9kwJVxmy
teDwCUyQ3m6N0Qrq/46Y/0SXhGvJW7a/5c2NAEXwaEjhVfjhqHrNAAfwHTA59Zt/
x6qrjUX7uyiKYcC+FaXnZ0wSnt/XjEdcM1/LAKUz+hfXZhns/He2Br5n50mqXhHO
mJylzohMdZX+ZFRyb7NX1duq923L/48s4nq1Dxwkgo2Z2yN+9fP6p0YUEYZvGKS4
HsHITrqhLVzarkjJsjBkmXW+wjWUK92KmjXRSucxY0FdgIoSdJ3mrNQKZIcOiZCW
1A1QBCnELfNcDHeJ8tb9041zr6VKLgj9uZnekpYA8lv6lAcFCOxOdV0n1RweKQMf
CPS15l7xIvAms7PsCu0EgA5WDwndtEfS9lu1NJFXwG0=
`protect END_PROTECTED
