`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8GbJCHBfl2QqaJ3nIwcdDSAhKDdt7PZduUI7cmY/POdYJWGrOspb8ZHJSeTYbgyl
IfElIH8l1QguiIjL4KIo0oh7Ii9uo32Q6gc4lZ5tTY2o8luA0NHMVamUeRdaCAKg
Ff//uPGon4X5pJcbjs0IEMzI+70yeQKAwSCw9DsaJstdlXtaIBjl4Es0nReriknn
7fwcqrrifRpy4jpdky2JkfNy/b2jYXHwLSwRImht6fAmyiAx2A/nv/YNHv8ZBElF
hDYelT6p7sf10vaspMbdB0VHWNEC/vLAxF3pz36dpH15oBgN1rmzi9o7Zg4tglb1
E5J8aGj5Slk2FvQqc9mGah2F18lDISQCB7ZgPoS0BZpCZu9fJemEyQHwwEAwiMIi
xLDlPcHvKJpwfL/T3OfhFoYUC4aXLg+nptnU4d/5o4NK/mmuXWB0olKQJ/DwN7DV
`protect END_PROTECTED
