`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ax8VF0bg/hV/uMhRUwXzU68rkdym0FGixSkZ3EbMWqhrSZtq+CkRXCjXNsfkvmG5
MBJyFpxGaFu5ULsHdHmwdBZdReVwQJDtkdwaveDPHCRXyUWGZND49vZwH6/Gi6N5
4wETsyHqYFKVfEu4ANJtuHsPDVLwfR4LFgUWnWWNAtX/8nJWijoyurtwWZ1iUAyy
bSuxO2ziRksRIQWH7r3p+/FnaPVIJPB8We8Go50IG11eRTycJURmT9v9c+lAK7/W
KfO0DmX9u3Dl8X5b8TtcSb/Z1K6Qrr7yOSAUVJPPMrWf1EUTGpr9NJKMqw5vC99u
n9+04qG5nWvC5ml7eVEreX1ZskaQAtZpzDKXYqjLuJ1ORA9a59LIqQKNJQm+KZCw
mQtIAF3ShcR0xSIsBSC31ifsEUQTIKNeFGzAxbeK6J0gpEbYdPvCdOtkquLuaAv3
BzB5BnytvXeBXwKd+7b/1VNqa0Yoy2YH5H5TXzjqhwydHwmOINzGCiTEw9RZDlub
`protect END_PROTECTED
