`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bLv/1bV+vYgwRA0oYHTsLigPl6K3Iwz1pRf1zSG+saY5ZZ3ILP2x7qIoYencAl5c
FoShgbBMgu0umXCH4t8z/oN8h1UVPf9nzb7k6BrT9u5Ztl20+0T+QS5/3fqQ0AGj
8wG6A/f1tk8K9BeW9tnYBdtPb+Kj+S95VSXP7yZRGmRwc1HNJye/EMVFueClvizh
qaHsGFEQvyTbMwaxqk/W7f8zxjy6+O7LqK4tox3Mv87MThF1Z0ZUCkYqv0myFjh0
1KYwlzU9TsntE5KkGFznguZ5HaIje7AbgsRXxpp2FXCOtF/ntqbRgrqRZmZMy+y+
GrlHvVlph2z0IQdTHOS4n+YzTQkpGlzwYXkpeP1p2+iaS7pTI3MELi1MPqmM0Gqv
8y5p3Lo2jrFiGxcCGp8WMT+BE4OUfZ3JKPq7yPpasqDhtkGpxViMdUsKnTfAbQsy
pVoweDMFQdVvktH6gh/svD7UHKTly+J7jBNmf7ThlV/5uQUnYhY6uMYjv1oNe40A
/HSLEtZSRIUlretm/11dFDW/3MSHUU8/Orig8PTnEDJSucwZbE0gWBMdsRQnl+rA
bSY+hFwDm7K15xbG/07ENI15f9TSIcFm598SuBtWq7d3X1Jv0zIblJHX7dnfmCN2
MysDO6sBYf1KMSHM1DcfDmueAMXjd2i6xGhMA2FMX+a3EzZGYlHwswPBQv6oWawg
6nYWBgyHHrAVADsf5BfRC+TdJUZDVsHGPtZieSM/+SDc2ZkkQSj+kaCCXlTA02Fb
m/oZwid3JVDDTiKo5d1Sc7KGloYACDQ5u0ywvVygZlqj0bfzjwrj3e2nH+6C5Vib
FoEapfSMTrv8MosWg0k2m9gYMpUomu8Ba7uwTDHByVdo+N/zBUMwLrCQsseYpfd4
ToU6ypm963g/AxHiEd3ilWHi+kVtCyTu+x0F+bCzIiG7z4KpxgRHzMj8zUlLzGq+
xXta4pOETumF0hVDkj87MKaoVx9G3pIfMzpjN3r5x4H32jrBq9109yYxHkivn9b+
O0u+3WVar6IfDtt5oE6lZpWLf/4u0CWYoLLTlePHBUICzPsW+Zac/aM29dzP0zps
nFYY5TWPQZAY22jrTHxOTaMnnTJmvdeZgkD0DbmIJv/+SlcSqdWCtH13OC+U9+VR
7c54hT0yqGno7I92WY4RYbq5/4WpXTCNkifU5PkBXda4Djchq4mIeeBKW3crhpM9
J5rqjGFv2fS9LyPiMNZ/mG1m2jj2s0no1LPlj3ac7lvugmqP3Izt0aS5y8ei9Xdf
UZAirFw/YxNG+lKRn5Ku73yMxD61+cTB0NYPgyKwV9Y7Bxt55q1O3uqULtpD2ouW
FC5PsGuzVJPI1j+lh4YJXH4MdI8ST2mpAofPAfZOrEPCGtaohxxnYXc9lSyaF+Gq
mC8lpH2k2YexBrhMsrXWhSMfrz3p1MwrU0tG80phnWouIPAN310WOhpMNOcjB9lz
BhDyb3+9oQ8eFCCkxPFTF7ep5WJneiUFDeSs1AswLapYU/ykeVFyxLaGfD5kDqMx
Rh+ZhKKGE7zpdW18ReptVacNmboX5nP8x5f0nOE5x4mnoZgzZYLCxt23SDm9DkPU
Bo9gWJT5lDpjgj8Hh6Vz1HsVnStnagViwFAto1I8RwMoEgDGuptOeZ8NCfzKB5G0
Ze43LhRizhnKBSCRHJs7aAn1OMg8N6cDchh6dWSeoT5verd7CvTOn90rM5NqggMP
s+bs0cozyY04LQfOG3Dn56ukXE/tCBq0zHiJLM2Vakk8C2+bXM5G0Cz0EwA2Q42U
QhlLpA6+qNNcTEELlZxmMmFtTihM9qbDzMgmSxkDzhbyjuKg6QZdzmwo+Mj5juBq
6+02Rpu3paqEPqThj9m1SIkGFqzDez6icFPD/LQqr+BF6ngpvNqjrzjf7IhybIST
KJPPTx60+2cHOwIlAHXzk/qs1HTklLNYfcduhL/FvCDxNK2uOW6Y9lj2TYDF2XW6
DwTy14fbdpXMgHpJhZ667iVGVpCT55wrhONsCycIA65KoC13Owln8dEqwNcCGepr
`protect END_PROTECTED
