`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8Ox/e5jmMHYfmmJ4VXkfjO3p/kzDtP+BPIHjEcpVJEPCCVQDaEuZzvCpuqgkkvFs
V+PHtbxvdw6ZVyqY/COnJT8oosTvWjHnaOXLMVs60G3ML4Zt5XHWu5n4AVOT4dyo
x95oVFZuo6JrwBzyHBODHncJzoLO2J2DDkUg+Od5DR+p8bE4Vek7GRmHd6d1/EJL
CiNsttWMY0fkprgCUk/+mdw3zXiSxBh2ahR/2D9U4Tyhq7jEMgAHZ8GtogRr0nUm
06/gGzksSDtPybmQmtyrzckJbYahZKdTVdCI2wBjaeXFNE6r+DsyZx11iZ4gcBeQ
E+Tmmum2otLTCOUPSlfq/tp4kliW4Mn5P8UT1NHChccMIn2FqihXgLZOEQMXtAyb
Ya+JiI7fxeQj1ZhGAlTeN5W4s67QbnzZYBHtoYg1mA2g7Qfiax9Q9rjITaRcAnU0
iaaV4QdvFHQN5plIAo8APbLZTjAFwRFXrbAYk9e/fRyCLABEZfXVtIYNG4sXATiY
Gdp0xhNtGgdnDlHBqy4N8LCjSeEsJ4mKmuDb+I8EJxd2wefnDePaQHrJ2F9KX5G8
Wzfqugg17E0epFuYdhP/YIwqZg1o4ItxZdS/jzAOlbMZNQa4ZsvqInKTfMn+vMdS
cIje/BxEWqDQ6yETz/oRoR4J8U8PikO7wOIES3VmbAJj1AoLFUa4d2njgEubEKAP
NZjwUMNYTz8ty9v/Uywoxcg6tssO6C1xrpsXxiJCc4Mz/m4V27CrERM9g2Vc3JBt
dH38iyxmQCez7938+Er1vSuvgua2JDcgaZ7ocrJOENwTi8PkQ3Mb8lwGMBmhT8Ox
93+6S7bkD5FSbTRLJoMSR32lgWyZsg1ylO5zI43ZUsie7Hy3f8xq0zcTdKgEE+Ms
RPjgJ6jN0+nM40GRhZEA8HQloSEquvS0DUa4g2sQFFdYBKm1cWh2OSKaNwSLjH5e
RBrreoS+2fWdGA3O56mnU7fBw/dZNQJkfk1bGlSUdaPwqGIqt9Y9mHmVR7YBDC/n
Brv3dteDtNs822BoYpwU1SOPRg/vIFNh3EHkbIHnPTUZIBJKNEphcke195eNUnsc
s+2rP3vaVZ6BruzljpugI/vLtNS/C2rpQKUJ7IhW3Tb0AWWNV0FrfHlaBW8dBwYC
5tAMr6Pw0+SwtEEo5zKY6cLGht7kYASsM7Hwir56ioLUxW8zK6zY74GFtZHYTyAj
c/byImPDa4Lpu+KeoNu0u9/s6v29+ZcLXWQC3BzNgNdP3P8XXtc7Pij0APcLoSna
xrsGJ/Nd/EV4qx3xO7aCYQNGVXfPC7EOPhNKVzItO9fM9hEmOqWmRGKfU0bqHJdQ
qV50lOEp8oRa8VpJrAJlhm5+nkYTVtZWYCQ5LO0A8a+Yhkp5MAASLHkPIE4MyQRj
FJvuq0ZtolxRhEHfVnRmQW3QUNJOSL4L1hUwznN6ncu99W8avICIRxXQJLSEBTBq
IV61OsvXxRIQTdK43cazjcJ5djopNL0m7gR6ZGMd65bTZNtv12CCmklPksyFWWk7
REUPYBnBpO665R5NgauhjhtEhFlscnqSS3ig65mbKLQK8YFB8img/ITplnV+DY3l
EkKr7YCxScl9MuoB/a0Q3mqD08q9LNsWhUl5hzCUVBgVA3swC+HFOQQj4pG+AaD0
/c59oq1KnEQgP2WgM1pBsZtBL4I76LIe49R6t53mwG/fNyNuxKec8srOLH0X2LiT
9kfSjsDgItoYMm3MnDJQu3GHLOe51i9yb3/rjuWi+ve+EQrzSS4OOS2a00K/wQpx
uEaYDngOh/BwOuh02eAq8cBk6DIkrEoTBUOiCuaoZSWkzpPS2QcXzQv2d10fU81J
67TAO/A3Wf9mRZlt1dDYBqrnM4gUYfUzBaRh8A9aNcM6027vE/ZvG9uHy0P90Fdp
qe8Uv2TttfgJkWOm0nNlqyNP1J10wWfK5cQJamBJgLMFHxlZowpibdpDLKns0Fyv
GfOWvtPR68VrJZuUNhFcsniykgzeYQPxV5NT5LNNNo+JD+h4ncEaa9wrjGKpjKtg
cmka4Q+G/FUmL5jr0UbAThxtZtO8woGtYRLaUdu6wG4Rv9kDzv64TfdW87deAk1Y
B2Q/BcLioAr/gI6iz8TkzzoxLDi8+fmxiFD+KWszvspUXPkM76Fa5zjvxBpG7t8c
eACz/9LanmXDfHgg9UrPYx7sXvHsaPVOQQ+F47aZzGg5hBqNN796PlUcILv6MbWs
6K5fhZ9uF3SUQu9wQmEc3pAkAkjQk88mNuHb8V3tMLd108f3A+GEv9+bHtqHKDTT
TQBC5SStcAem03WW1zT427htjJUv/0LMXR4+OeRAVlRys5ioShQpMkj1KP/3ncVb
Mcfi8jWB3uIyoFUejry7aTRwnsT9YTC4MsLt+V8EuTSgB39B8M6eLhA58wtASCvj
vtBvK7lrZv7OJmrhdYHQckCpZJhTfsdCAvwdI9bkM3/FFPDxIEGZPfunFSlGOeVQ
gyAUbeBviofaNR6o3sTwT1/8vAS2pXfPIlKd89IArydD8qDOSt29opG3p7BqsOux
xOK/eYIKMvGkPoa+J1kevMjwM16+s+LOSPAl+LtlId1yKgdF0N26H3lRGvO/0CoW
XLFuCW9MAQRvOZ08wuQofacYifRewGY6NmMxyMNXhNmwWi/fdIVtFVnxTg1QoGOk
jf6xZB9qURo6X58ch2NQaiUg3/jtWty1oG0sJjbzd2JxSwWtEHe2nQUwirrQwcJl
roRenEb5ML3JJnG7uY/a7LoYsHHn37bT92W0PvBDIxHXxEy7Eo3kbVM74XR3Irr0
J5l+JdH0hTwSI3yu+FWaH/N3oclrmYhI/ZRk+LVSNYnXyxcBDMzavJa+Dn0uuzg5
wgHQZkSSE1n3yhTfGDSfVBpjymdjbKCDEoqNLvjUqrrj3AWquR8jQXWYx0/MJAvX
6jpol3gXw3y/3WxrRLL4if0oot7bQKMQ0EMjzGjl85DHXAaKrFoXi/Dsct47SDaV
WSbHI3bH3tY7nmNg8fNWfo5hYL9WLdVj23nCxbphmVXIYwxkmFPUZT+Fd/L0hp2j
ryw0hdUM+KTGem64zJ34ygi7eNtEj0v7YBOq5oMeRCUU8SaJnN962GxdU4JdznKh
L+9DYTrJFxIQIpw5mL1z+nZyZnmWsMEb2OD3Rs0uyIy3khz+6eMsUOgOfyY7Q2a6
9tdyJ35vzSFQBf40qwhHaQ4UVx4oitz+MkVVu3XuVmY1EnZK2OwO5t043ysrpwIM
y/xLR93ZuG77f3TTRJBapr5L2dIaaYdOHnVXkO88+sDgbC9YxEl2Z5x7TYlwlKBt
NZ6LQeWktdySzfrHFpW/DM66lZzADhdnxiLf8YWZlogZh7tQZdiDYGJUNNq35D0d
JaNdg/9Bem/IBeIVAv2f7qd1wqLqcdnKr5Daf1FwOwHsnpcczYHnYThaAXRBr4cm
gfQVjpoHLYqq2YzJmRSNtbeD8zHL2y5QbEzXynQUC9ToqAEH7eqOqislqTaL6Jzy
YJNZQq38VL9vm0xBKi1t6Bq/Lal8L6iQmRypl/c4zchW7doQlgRFWevnc8bDHEOT
zXfW5uYFJqoVKbtMZsqBNzCXcvdvKP3t08vXFqopN8YxxM7M/UJH/6z1uKBQsmEj
c3ZyJ+T/QyYTZuPDOhDkaF6zqoK46Wl/3wA5jvclsEWzte5j7+pjnAlZVwQVIBkM
WtBsY/0DjQ96ToPphVufQgZOfRf2Db/5FcnDH6HhF2W7ivbSAUdi5IWU2GiAXalr
lh4nYhvLc7jINzWPFXs6nKJyjWVAzZVwiVzsLgo33OFtgx8L01M2Btr/CwmC0PkV
r7RlF8TssItUnce29zvQa6KTMgpZ3trPczeKkl9aI8YUBcGFHrc7Dt17Hu7i5OOV
ASBuDCx2FyYSpwsBtyYxyqtHljUq2KC7R/27WzXeM1k3Z6/Fw50tbIVzuCsVndYs
zWihHFVADKWnpiI2WrldODIR9LvwMeStTCEu7UX5QIozRfWaXebemzIkoV0hedGr
JocDSkGhc1hwiBdX/6Zb4sVQvOK39ohUBs8fii5S3zK6HFWE0plnS68lhnXSKGEX
m/HvpUTeUHbH7yUFcWo6F0Dr9EDvPYPds1+NZ8iY5z3tVTmB4zW71EeqWXs0a9lZ
5JUAxEo3IObB7KFA4F7IOLR6y37syDY4WJ4ZwndEUCTnErb6P4Wy0ywg9H+FxBLh
NCjNgJejZmzJXukMcQwxUwGG6hrPZD0ZqUu0zsPMBXxZ/Kybi6OgXwlclnVwKu84
eHRUyPSUefdow/rGVUYo5pgtgK/DSe5SeyhyzJmD8biDZ1Qc3d6Gce46qo7LQ4+f
nHJxP0UcgvSlwlV03/NT3Lm/XNraMGcsO77j6JSEgRMPJJ3iI8NO8Nj3/q7wgB+u
WAQIuUtfXMSUFQwiDpjP9ZTWPQX1BnDQHKVSPS86PYgnohW6YKX13scOgQzAYVua
R/F3igpnqHyk7GPHbiGULMPZCvpWIarU3vR/nDxvr3JA9XdAoku/PnYqffAa2PMT
vsQy9tXqkROJ6X/Hyyh89fKDt9gdm/LMUtcfOIbNhJgrfE3K4cTD/G3iNPUfAJ2J
Vf4ZrzjVwd0lSzsOFGfXMfyus9qV0tLMzXyqqmEq13bgl1dmzE7TMS2Rv4UotMtv
T680rIgRUDUFQFf++xWnL7kxOD3vucJy0dKgJ7IXJbxFxod9sjv0Y2rJVOAmUAI+
W9XPI+PJbg6ZnSJsvQGbZ7+nU/lmY+87aT5hoZOrcRo3K1LHHhG1OBulGwbACV3X
njoCIkb3ZN+aSxZHCDZ5gjKJBAcbVCSEZzuC8C6NbnWq1rKmrjxYkkQHF6eF2LP7
e1V2unaL46W1PFot/KRfSTnhfDxINyAfD6z6M8xx6DgTmxfPiLRGPN+TzGx3IS0N
TFrywlItoYwKzD3B9/di0dPnF/WOhTSa4cnCz/WfmLAWjlgXWVBMbB3okSiQzWBN
YH5OHjOQ/GMm37aHS0OwOxhlxUiGx2ivg5ldlGWIl6dDFOvcVIm0eza9xVxUe69h
uZkqZkufU5x1zZvHDByuqMivfl0q42MDCzHo17jWTt1FchsS30Agqu2X7b/31rVB
XEX87qBxwCWnwAZ4TI57NLBeGhIcXLaU938XR61Amh8Of6BDK5PcynN0qheEfwxC
5wHXD5BHXSg31eG6jIOk3jxh5BAGt+8lWfEe3Ur9y5uA+k6v9x7UFZNs3Ka+18D6
avr71eI616I4SW1d+PR2PRmSbw3sp4z8sJv6vV/7XehSnDyHSM3jsypPJBGfkLqn
7WOSy1j3BlmiaEPe+ELM0kegUtKs5q+6rz0K0Dp4vy4dKHfeDmpgO3bhO0q4BaYF
ANZ7DHhGQkmFQNI7F+ae5AZ3qXumRE4LJbsW1snws5ewFisNf2fFj3m0CKZTsyKq
m2kIFO7eIYIxAhZ6YUOK18t3uamZzBf2iTNYtRWMaxsGTfuBWW7dYI/U/uR6W4TJ
0MrIH4MYnv2ZFJtghziOYvnv35A/tWNQkFtaC0M/izsSUwK5GbKrqO68BonnMS8I
FXUgdFXlJdryTGUiUlJcKIaGZ/ntEGelSCFCNIqrVuvx9cjlmEa66Wm+bg2CSsmo
w54wGdsph7+lyzC076XQk5RgCM62B8U/c5VVgfGgBawuF7HFwg3hQgnDGSTOjXD1
N9MLvT2ps1vmfjSCeiN+Iw13gVJgbFyi16FBHEyhB0iOGa5WdeUH8UCd2hNeyivo
vPyLuD/HTxduHN3pIrkDBnjYDa71kLoFGgPk9C7uwAFjHV8yjrdGNBaE7S3GagJT
5aQTFK5p9qqkhS3hbeRSVy+KY1B2yW3amLRE/n84lifdTjP/0frAcc5kYacpAqip
j+QVIFzEs4eYw1ks9UQE3BtNougNldXeyB0AgzrulHwAWUKjHh+1zrQFR/hs31Ow
ZIKpzJWoll5PLloTf6pPuX2PPYjBqp03mU7VY6/5+C3p5RIeeg27QHYCC1cJs0SQ
dw8AoBShkajcDoz0IkYJ4R2jGii/7/iCpAUbwJHlUakB+WDN0ZGcHI4frNA+4Hj2
NRnk+whuYCCYrmWiXo2bBDDOCX/pwhWqhmx13hJH3W9VPth92+HEkIImeJgR+idl
nmhPpCjvGVNeMSdoLnXBwMqXnvHWujgpClSWkSgE88tbDKF2XMU2dusRXCiXuXBh
AUS4qxF8zxOc2+pvgpesPY8lIF6ZWgbS+6CsplwRqL+Mh2q43e2ckE+yMv226gBl
TVnxsz/QOBNlGC7mLP+D70SzsuB7N0D5WA4UIBEIDDs7e5YumxO1DfWu1H9Vn2kW
ptzTXAVhl1Sc38KIFKs+cm9nD8dY35bI1mtHcd65IqRaApXFDotxIE1CzkY9xvSf
SPcCtYO3+dbUmHCzj6WHGpq6LTuwtJ79YsbNYFfdrByN9iIn2kJhubbDRYkw63KC
KFvUXukpBrxSXWO+a1QeTFZRKGljUNZcQQIPvTfv4Y6fGuqy0okMMQZUN8/fIZUr
sfM7r3/VSXMNmNaRinLW6+dQQ/SZVr7zlusumiFjhb5S5eulCBvceBqOWbltneKY
0DOObih77ndNvO/2w3SSYvX/WEXZGm1uR9YXWOOU/UnkgbEdiuDyx+TwiLgyZ21u
N8wYKD6Hj3JvgnwcBwjPtwKwYI8mpI9Wtz58d9PTONgKT+zha5twepM+Xbium2tB
D3ZYOmY3FZNhJSOH3br3VThdDcP1lPiMqOCwSEmH8De3OUcIJANjZg8P3PP0NP5p
5nUbJMrcOamOQQw6gn/lnGVuGkx8mNuo6S8VXIV769BF2oR3L0UtinPNPuJWtyst
H3X5i7lnMOxSBCtk2o6iXwgXstngCUJsm4YLv1ER74y/7TqxhCOY6x/U24PK9DL5
0USQYk18uX0ZSOkW7ZI5rKDknRkro4PbrfSxTuVQH+QycecPjWnsjqVPOdPEDT5I
S8yl1/W1qInKSiPJdXc2KslGa2HS+QBcafC0ARugMtzTt3LdUOuBxpewpWh6vrU5
0Y+GSTTzFviR50L890rwJQDWQrStH/JGoj7sEHIHB9HaJBSCG4R1GGc0FnfwM0dB
HoIbb+klAFRx9nfnPEZ0Fqpo7ifOP9eQIiN30V8mIakAP3BZxjxgZc2WuaIZfEoh
kYFrDYV7aQ53qOqc3BHPiRj/rb35Xg38ICfyRnzfpdagIqLjJquoyKUHIaBrcJ6R
eTvloZMhDVUmUVaDBL4Wg5l6VIvdpwVxSC2RjXAOGt91c8uJMN0B2G4kxjsptTGj
gBafybHj6GAEiw6Da5OU3bmUzi9vNff5mxv36AReqOap4UzQPAWzQBOOIYZZ7aCT
Hw0txT0bhiglRr2iVumG+gNHFivLAml7FTvoiCOivQfmKj/CWeEB6jl5+/CkdmQ6
cDWJhQFtmxDEWn6UlcNNEKEdHmMNH9df7bxYRjoS14QbiaKr/33rTNxvCcKeuCAM
oqUQO6uxxg6BrQqa7k5Rx1jaITVx4ShESTYtMFRS07aU7wNK49/88bi8+4bYh0Uo
uVb2S9q7XVh/Ybkmx2rrEXvN/e162gH82D3bC8i1+jv+HtKsZM3nqNB374UR/aNE
jaYXRWbNy4mP1r8BY5q2PdcufyuoNFpgJZzI7VLc0e4utNyJuXTXRRSqtNq7J4se
tfm3uZtaaZ7+/OOfFxuvxnKx6Bo2uUO9qpriI0MBbC6F323aCuobfR6Hz1d5gnzf
HubVqs4Ub8DULkLjBrOR4vj6vsMEOyyhFjydqXfk4SQNixAn88vcfNR8JKK97PJ6
RKllIFbMFHHxLYTQ5IQwaWF/fHHXx0QWwJLRQynp1VXrZBF8GUQLhICywFcJUPzc
aBmWSlJ8g6JveTL8Tg9+lpEMkcfpoQvYk3Pc/KSmnuc/2vON7nkkW5uJ9Y1VRJNn
kzkVJ8uwxrHoelEa+niLQJt3aKDXuUMboDiRizDIhEfN+Yz1OGA4qjjl2qkWf7rm
6PE6uwSLV7ygEQf8AxT3ELj3+c4fBjpZXChzyFdAJQaVGdgZ4r8iRElKbboa2y9B
XkSdAIwBuHm5CX6k7yFGIBO3Cg7kRLJxolt9l/WqsLj1w4R0uPt3PF8XbTSjKBr4
yRmx3WaZ/XExZ3i+VaX5M79aZ/PJfltyfTM615bWg2P3gJXpOGGeDVFcl0SPWcSr
k5VudmKJIzgUCDjT7xWu1Os76uNYrkNXs7w/vbbUvDxI97R5Vn5cV8/C8zotiLks
/CHZk2RG+Z5FNVsqXWLpXszh9to+O1HRq11uhlQHSaq1/S2PGu2OFSs7VQWeNRES
EWE9rxEEb08KMN0ewEcA/saE7KWrLmEpZIEOSHcy4rGIYYesHeYtmhQWMZtShkQU
f6lpMfnDyh30cvjKUyXHYLpyFZ/SRqe4WwR1bSUtv13YSXpZObkFA/My7JAW6O6N
J1II8xTdeauPQ1e2Vh9tkCxJRPAbSNppJbJDheWvwYxsnCgBJFq41V8+87KxyoYD
hbx/kjuRdNoOifuRDf8iFpcOjUxZJ4xkmTAVvYi+hURb6+/Jb9xoJ3wLMf61+Mdr
L1RpfdmGALmIcpAC8eoqUIUDERyCvFVuDvMw8PEDG74mvG13o4MRpmZuVVkO4Xuu
h1ybJNTSwm+6WX1yc2PtgXuFmPybyp8CMW51KDDFTE/rN8yiErG5Gdoondmsx5eQ
OymPh8my4hW144u9+QOgrhcN4NqzyfHcbbDLRIeOsFipak8NdtjLq54VCh22uTys
viFSsKMWAmLEyz9pjo+Xq3gMQuzso4tmUPC6p/wE/V1o/nMAJ3sFmFOpThDecc/2
zQZlSdSKLusfVrw/K4JUHo8g67x14WkKkkEVR1L14S5ffmoAqkaYgK9frZDGeXXx
/xfLkE7PrCf+GXTIzMDewg0O1vA81QJIJqAvkKkTJ8UP9CriDXedhtYJKa16zeth
rKp1uWWxbDxPfjSvbTwa47x1mYCLqq8foiVi6rA1PRr17A2c0gYdWdHoEJfiv7//
Ra44KQ7L68ls9xOmtRVo1N9HRVEuXxqMwC4hkioolETzeg9WV9SEdziHiZRCBhln
BPAW2ItEEt7PJ5kOIGK7kT8r10/V8Yq8wUknjkJRBbD/mbPPjODkTf7t/xHSeCL+
YL2+FHb5bnrYfCYQ+dJ7odvDAxxAN3kYJT5vSpb7pQeYrdyZbVDkTIaHb9wJDcOg
FuhMCCw1oQxmpfrrA1QQYqva64ky5yjMDAW2LTzxRTDqSfOw5yZFzsWnbBahCjnL
l2fUYX+s5zCBOybUp6L6j9d1eE77OrJwwop0NnI84Zxz+4ZvwpAC0zVrWb3euG4p
bpGNVFKOwJCoTyqft3FnMW+X2tM5B1T6gVabUARwyMHa+8DCme5w4rB8dZY3DB7l
cYpGT6cSdHbItajAwyM60ED7aylo6zXdVFCpOnbPu/86avMbRUo9fRzfTLkCJ6Sq
omuzqb8NcNBcrnrq3TpYVevxuX7zOxaEB7vP8QFBF5p/xyk/jXPad5vu2zfXYxgL
wMfkWLIA+a0Wne33cGY/+ppIhDZfN3weCGKk/N7US/pakCEOA4dMKEr/79MWbSOM
xk0U3nohKBBgMv2C5pC0gf4xthDKjYPgK1ouI7Zxvo33yEef9M7n1bmSizjm6vON
vmnjqxVwi4Bh7lLX0q+vlGRVh25iDjoU3/wFjtbQsHdjdIQGEFbjZcVc8ZXK5En4
zXaJ3KqFb0xhGh3UIskuq/a5Ru0ky13ZbnDrIsDd1z9rlqLrO8B0+iu3XKaFRZCB
2w0049svPFqfoQxBqGKkY/PnzQ927v9dJYoWK2NhY2BCSlBwgqEzCqAsCvBgvkha
VigoMMOm9065rj3DW4MjsuksnDob88uqm/2YrjJTJ9z1c93DsvX1lw6PK5LOnt1W
ziSyTbcp6o5rQf56W7+49ywKqdTjsgYTzBg0Xow5YvcQUUzk72SN9Z1iqssr5Xyc
8xlfgXnxfOAc2c+ijf66SSWH4HM0Jy2rWI4vm3alIsRURW9iAbUwoL6M99sxQ2Zo
C1IjRoyM0K32I2Zu4fFhqQT9HQOpUHhFcI8cibnxCb998/+7/YeSa4bVd8HuvCzy
PoWQzmeuLp3shLMfY5E0yFVbVzVTyyUvnLT12WKiLSj28YqIbDQMDY/sB58+J8UZ
f8GUJQKOaKKrQvzgGQCjM0uKr//ynQ4xUKfBG/aJDYDzq4O9yqaA66kxlUYLK64R
pCosf27HOIQDzJKz7bHiqZ35qwGNM/u2ypZhbZUJL6krY93QeYfSHB8hu1O+2FPX
QfmZF0npramte8g2Ups9cmCeumV+Nnexo0BjtIZa4FRSHgR6fFXUcNDqmP27BmSn
eNLREd9V03ibrkgd/6uRH8VN+c9TkD3wAmUa7uBw6e2mnxSzUqNxuduk+feak5Y1
nWZX4irIY5QP+9n+EcMnpHD6YBouvFbAPDgRqVfWlT7a3FJrf3iEBztzW49CDzuh
Vhsp7dAJpILi2PhK/PTTOMDsiQzdC6NePiAF13uMYq8jra230S4bFVqMpwXmOqei
ZJ45XJmG8UzcKEkd/RW4ucC1UgHDwauFH4/KFzpp1F5qKfwApnJ3tMhNn8w+CF7V
Jkm9J41g/3smwzTeMK85+qSs9rRsmvzgvL6bHwgtczHYCWvOBZiC67qySbSG3vg8
DGHZUxXw68m/OO2EJV6xCiWD+sQdQGzfhC7RjLO673mK+rXuTaBGjn5jTX2jJXk8
ns4mg7GSRTGKpfB+hiUlGXAtRxa3ofRjj5whMEu/IFgbv/sL4uLfF9bmDEHp4005
j72S/VqaXua2HO9W62jgo6ALeNaPpYl/4JvJqjN4Xd+ez+EtuGTJBxopDIpe4bSB
l/nXKybrabkDC5wcbdzC5BKJspwOfqrWkFNUsKao7GZrRSWDOX39SriEYD9GiO50
MFIIpgnqNxyBIUF+fD1Q+X7VWksEAe0EYVnzebdWGPU94BloDfny4ipkguMqIIe3
g1+IoX/aqL3FiW6rov10CSd+B4xGRO7GlKONULEt44rVucNTf9Fw6trI2eUvLePg
sonQ3Jolqw/QDFTP9TxckQ/T0PXbUnRejHYfPTjp9plv8x9wJvXrg4k5nO4jdrjK
97tYWcclGlKS1RV2XQT1BvcutvAPkOUg2um0/avdB0AzKL4bWgSNQLP1TK3PvNaO
WksmJbCKUjoSSF95GvvwjrkhKS12tgLjscMzUxR3Of7l5WJcIn5vwcxaX6W9+ptg
f7ag5lQWhlZSRcPD0JLmQAxqbufJkOREfY78MSeNA9tDVahLuD3HSQW5oGNce9CQ
iel8S4f/G7JdwADw20gmGhHMchbLLkR21fPLNU04qxP5VL9yv558CR7USkT5+f5H
n9+8hv37Rk1vRvbRPYiIQb/+3uaWM0t19fo1g3YOLtn8TZy7zgzYn+Lg6zyyLDRM
ulOVoVw+xExKN37IblXWjQkCL1v77UR0Xc0G2zjV529TvxTOGRWSBP8SURfPkOoI
uMv4w8XpoWTYjtV5p2+q6IJGIZEZxh/unB9Jbw67y5C764EMrPzIlLvSfciV/a+p
R9JIR6VFsPeitikqDKH0kT/Tc7yN0aecPK5CqYkEDy/EGU5AUTgfb6mrDroF3DOj
HN7/8vYlPCmeZ9mwP5k2Eunb8riDj0q9tbiPCTIibNPS40gPNL9aEpQJQHezDjiu
t5p2D0gUPYb9IgWWaL7faQ6SSqnadWJTpV2bK3w/zGMzu/jWFs4uATrl1iInJeQg
jVRcsS6NUYN8LRdnK91Odry97nULmfjLqqwWC1giJULZoEk3Gwvw2W7TLjafoyZN
8mh0q/sA5UK32zR3ddXiv7DII0v9pbDmpbmSxUQTD3b8e59tlchgNtoGEeAhA5RG
7UsIoGUY7KdL+hAtGWCbO0hFcTeTdU+Jpzkj2hut3dj/ODN7sQeRkw9Fv8aUjqHO
SuUj5ZnlCdbxaHfe0UxEed/ez7cnG6rXLwiUOlewgjxxqogfIhOUVTmW4cURbZhD
58NjGBof1ThgDcfao+9T6eyv+u9bktiajKmfA5anGKRhBPKUmfM8mVAPTkRWQzwI
TVCd12CsR0KdaeHCEi5/R9+LJRoh3j5/z+LbCX8xAVf213ymwUdG44KtZotTst7L
F9xx6mParlfIu2ETUEpdq95I/TTpJxEOG4QXvJyjQQCPEuYO5VV7z56OFLLkCU4e
Bs89wesYJ02kZUsU0vQGFQFTgQ88T8Dc+nY+ZDnLBEaGau2j57dz8kdeNe4+FtPH
3tNCSqn0M4ryMv4qoxh+MnPygSFLw4orTg8QY8Z0iMWUsxxMmQ2GkW1QllWWX1l0
Ure4G9qbZXWI4cN4l6ofaW9MhNylVkyqIEVI8N284tJCkP+AhVHaI10HTfbHTBks
CzBw+0CbXEBXWx0U3Git/Gt1txabP332D7KCemgBfI/M4W12ncsNxTU6f9uKgwgT
9mGDKPJoV0IlRhRUcTpI4SGFEQkkuW9VbFVIiFJZVvOqOQTaMdb+9V4rrmy/OsG3
xqr7k3EvxBqIBdB3BjnnUozXPE+N4/oyf5aXbmAH2cJB/amAsYbUqau2Ue38h8ac
ONDx4v3NM8/7erfHLPYZIiqN4mnVAlOy1QgineUKwcysgGATioShXEd2xYk5PEKz
sSJqiUESJ03BNeiWbkW74t8b6ObU8yA2Glsg8llvtGsDEuxCNTrlG4OmLP6eBI/u
bYaTUk+eA41DMH5v1VmdcF/Kr7Hu+xr74dQEsA7awcAFqeCPdkBtJwpheALci9ki
Nsn6mLQSYwH377qdWI2kBX2tENq/UVfogTXl0xT3Y32PYNVdPVT72LzhBL8llc1u
Fel5EZE/4NXndH+D0sB8JEMivxUn0sQC2euamYXSkDPoK6NRQwOVEDQwUtot3pb+
lqnjWP3ovz+yCC/s/P7SQgRx7uJdcxghmL57G26n0278NE68cMcbG6gC055DWSAQ
ef5wqyl6ShXIaufmjIuorK/IW2rApF/u8KdqiwNSDopn6Ynj4AYXzKE+eraux2On
izhNN0kdQOYFBNFSxrS2PnOEbC8D/BTf6gW7nN8q7yND02KQqNufIZzydGJwVMt7
DzI8gsc1jLfrJZBbMryeXhAEV5rDVgkawnoZ7jvpk8PTans/p8N607I7/h9RUCPt
OVXgmHi8pt09NeXgLLLFr8xd4QOdSJZPhWIHuWKifsozlZeXDmmxnEDER8baTbTc
2y/EXMQDBa4eRiTmGBqn1I00ZrTxt+8+UqpYAQxGvyNtPC8TricfZy25tpOF9Qyx
paHSDsT8aS0L+Y/poK8yMbsUUoaN5zDI/Lx0mfdjWMdZoPXpXEQyX997yrPU3GGQ
St/KnFqA/lOABF/EBVUDJeYyZcp2B7EXM4uFAJH8cDEdw5Ef+3I60uw7iA/ujk4L
/IvFmRH40NPPENSw/n1nXBBPmLj6XPCoA9tFgCgkDc4LPwuGv3z/G74X14GPuZGp
2KhUt5WlkqcCTIvtQIljJe4+5nk0QJDgxjGWeFAMkBbk3QG/fgqOM1wDIXtMkphF
DvNe6zX3Jd+qwgDvJYXbuPUqkVPgzY9n4lwB5GBqWZ3A6xKweYSueyp6wtUIvv//
ZsprEIYGmajcmNGJOrOx7psTPV4auJ2F2wxtufp654X2XIeYSG8tUVEwrSwElfU8
CnHHYVWZixw+n/S5I6QIMJX0rMY23Gvn1j1OuqCrzM/3Q1VVq6BVFwLuCIpC9azg
kgx3P4GwXj9pVMjdMANhjyPvuzH3TIQZOXx9T5P1WSwloTt9OpRTwXd2z+/0dh2X
DCw7ODTkOTXtdamNANtmRSVd4O85gGymsRZ0iYIvzUlKDiSkRfqFEtYNUwbEzATq
1qTAgwamLF0ClGB7i8LqyQmWyFjQyYWxTfGRRfLptamesomILS/LvovbWvYt4iU+
WhA9tzOTFLo1H+1CXCjdN4UbDPNwxcyqDOPA8G3GKc3/f8XHfL9/QZhLHlXkadAQ
VrBIkL7/Y8Ab0k5496Ud3Ju2kVTX69/XdGv3utzXYmoH+5+e1m/BHltnyIcBsNXN
kG8u/rA+t/miy5HiGfIvLuwFQv4hZfE31MYh80PXZcjMkrngXL25qZckvD8GkWDB
NVWFhf7+G+gxFTq7yiCWpEskf6dSBZ5WKckA4czQNwLsTf233Rgj7biogPYikLDH
U3Kc6Ts5AlqhlVh8TofFIVDLuz/jxCArc3mJwSC6rZ0muDpXbhr4fOtDWcn986K+
8IPEMMBmWlAavckk89yBmwGJo8AlG5eQGbpPo2Kk0Ed3r8ZLKcJqrS7jw6BCAzfy
zBZNhHLqGDXn1nPxK4YdaTFTSCsUxZNaiujrsn7KpI3oUMYPmp9RHqWuZgU8pRoY
iFCyNGnGgXfLHbzA3kvPkD7GASZfgk4cPBzCgxSPMlFBfAWSDuSDRLHNr/VZkbWL
7bMJBSz322DF1Ys/E6lDyN8sXhy9sCuodSGsuY09MYyBi1rVv1mJcFbGjbl+go9T
OW2dcVGJRX77mD0NEYy4F+7Nk9EWx656JJPvWAw4cJ1J6yLKDmFlv3gZTYT5DLvW
T4XduJgLoEFB5GArSWygHQP7IHNfs9lGZr8BuKkVGeZde+fuTr2SEaq/fwLC+OBS
Lm1mupvJP5kY1Q4rslerlYq3h8aRMbjloBenESfYEqOWmBzII7frtIgEND+VhoiS
sU5J4GW8gBpluFPfH2G2vhUlYFnps9S48G6KdGZLk0ygKrewZjKZr39GIK2BIFbX
1/6ApRMs0J2LjpMVw2viCCqMtEOaLckgy6OZglSzGx9HuUa6LDUzgakaw9M2xm0c
iTNvuTJWD57gJOwFPFtPwxvo4BNVCsd11t4TjdFzaJx2/zwjH59pW/+FTrCwWjF1
2yd+MZaHbggoe9vqcJIaOCxULw2bhHAg3VWUq4lR73UhjZAomZFOl/h54+MubaGz
T+NnQ1kVU47z7jryfnYyByefN8sv1ygJVGJA15lbQW8OM8kW7fucnTEJeBDOxKUq
Y5v2O9Z6WjMW2k3REe2CoQF8AqrsDdT3iwoH2w4LykB61dyTMxf8Fk7cpn2nhxSk
0yGqBUGM/qkF27Rf/8RoMg4rOkg4M6HBelfkwRehrep/WpvBWchK4EkiTRaBcMGb
CUQm9jrbrnhpygUhoUCjvsbMpmcLeqzrKbCU61wVl/yidhdiQ8uNOXUyZ7bngi83
7VokKv/1apBWtBgl1gSfUW4r9avGnPA2ou6M21PpMpEHl53cls07y8bUfA8riuwG
LsNyAYe4Bei+Xr4jy9mJ1h4fyT9D151xZ+Zso0hajZkkgAsiTbE9CLY01NeNrIwT
JFRQlDoRzSMpv4aGD6DSEitMvfzVhSFyOzME1PRvKemW8KspNv/16pmnOvBQP0Uo
LiaqQA6t2mW9AuNYhaAuqDK7A8QSkfO6cPNUq3+G97g8UiIURPVOqVubCXYBp/BG
fNbw9ZN2P9dOiydxAtQuZ4o6AYE23ZLKo3yDTvDegrEa9UGsIt8bntOEN/1gvYMt
PNP9+J+DOaH+w+lcB1S+kMqIgIf3nlQrEmiXX1D+25pQ5/XD0q7FyBfudyINmM6f
Iza2QVSZlpNziKlBYvvDObaDgWSBWobCjrkQTxCrxVM3D667gfe2uknDBvs6yLZz
O1hx0QylxNH04gf2gq4Zi9tkXOjJAIVStNknJ2a+nLsRxbOQfkIzrZTSEerlz/jG
zA/oD4v6O39oAdD+s07lCj3EPvsr/5eKEDHimLhsnf3LO5FrqjHau2aZ0ZzsR1Qa
5vfj2Td4VfrAaKWmIXS/knD8Y2aGDNJCpsB3VxWgmy9aNxjLDDImZD7RSu8cvJcK
S52GYqZKC09mSOaiBnXgfmwk2GQDx5uw79GAOXTkk1CsyxspeIlMet6lmBMiXeQQ
upDyO6NKXIa2SHth1iVHgui/V+N2ykw90bd+UnVk0Eyz49opWCS2Ww/o+N3vNjKA
dvpDbtzxv2VM4jNurYO7XaoYpjdWQWa13UyACIwTC30CqYfJhJbpWAt+vAF6qqR5
xrHPj8S5jDbt6hCnRRJwyfMAf+pGJ5ipfxzwZS+kOgjKZaKXpTEb3sqVjaefqYqR
7W+UFRw5krmFCqlzQAuFYeaYoHBhMVC4Ls5iHKphFKAe3tQGhRojqBIct+0CVYB7
OPkNiv0YljaAeh+5+huoOH5MP3OZrhSdrkIASJ05YvGc7E/69MF3qCYZ71sswc+D
4ZHRpxFzx8+BBK31z4uXfUcedBHSH7aNzQL403VFRv1ypo9pcArV/6ODYZXDcJ7x
5w9/tw35quQDXrg8zrBtGqn8IzWRMMazCem+pcGLMEuWRPcn4uFZC7fehwDNPm8D
GukTI01AqeHN5lRgF0ULXen/0q51RkGf437Q91PQovUDRPEPPsmrp5QRs7jx0vsR
RVFaTOVsFOrF3Qj7Drb6rOszS2ssvmEl3EKg9JchvAZ50eCK1zRIDb1viUkx4PUh
7zUfWGqraJTxJHmYmPfGkHts2+rvp5npyqOuPuMLnaKSqD1bu2HnG2rQt7s1g+PO
D5gr30KRKyyaaXgIRWmSggGgGxjzL+Ra3sN6qFY6uZFT6D//kdboskNQR6tQcma+
v/QSxX2duzfIYIT2tYK3//bT9G0onA3Xb/9WVbMIu1a0YugprEzCok+6hYrkn5a7
D4s40B4tS0H5Ej4/h7T+pAOcaXZdeQE6USn73Zb1rWAiQcmng4SoeHhnjuYDtQ0b
TchFkNFr03z2eEDq1Et1jw==
`protect END_PROTECTED
