`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h6IoRKOHdoHkl3Rxsc/uYcERQIdOPSzK9wjqHf9mV+UlRimqJV7sTGxxsRdGpiXS
K2dLNyePjTEKX+LFaboTN+WgbHa2zKHzVhdWTqLCVT/RQ6/FFEO2ypLSRk/O4u8Q
AreqstfURu8bBHPTpsqtf+VozvPJQYR5OBiRXV7PxDAUrJqZU5xDaiiaVNDok0SH
Ww5fVr7stXU5iJIKP63zJpAp/UxcJ25Oq1FAz98LYE3amQBYatLiAC0uke6J9P3O
UbOJeXoYIC7wZdUsWWw3norfaRWVuSmXQA+TozHM9FYTgYBonyPisjsxmpxpd852
fQYSK506dg12W75LTC1qZY8db4Z8/81jTPtrghRrZh8KPeJ7A471yrIaqxEGkYIq
DFoQ2c32hR766R5V9LC1Iipu9ItqDtJtgygXdKVKTDJq/0BnaN/+G4xdhc1EYvS3
ZgXNdHB4bhS6Za9rIaIIq6lpMhhqaZIc9bwzK0UwYV69AmpzchH4eq/PfyoAFwiU
h1/PO92LGaLyVhK190db9NLa0EFKtS5UnxIRVMNxZzkpheLM64GmkTtpaix4Kl4I
0/brkNleImQVzzont9s8spONGyhOIHu67WVNvnFYzMTXlIg0uXnfpTJH9iS500yM
QDZGWF8esVwMy0PMt7xrqP1W1/+Rv4RrEg4mu5zHqQJY+9zIiPl8s5xSC617J8N2
28odp6n+q2MXrIsonePbOaJuvnfaUEbXuKEj+uSf2ie+2/RM7935MHvxZ9wLr1hI
3riVb5s4OP5F3Ww1rc/Wq3/NTidrrAOhT4VS8rRd2lscgpU2vexrxTSDs85Wor+9
QEoezWCJeshf06c/JlTXuHjR9mnbjF45OG0ggfss9aGcUA+MkDxrOa+qNH578LRk
D92g41+renud0fJwjpGc55rWzVZUAjE9l5o3BYYpMMBROTzmESu3Iq1qDZOx5SMG
vhGgiwFMhdT2h+0iCHZdSdhzkACimRC7M8SAuZqLoKQys7RYZ9Ne/2a5cL/ly2zA
SqyfgtG+CM+tJxfffj2+v+BS9hsQBjmwYBX1cye4bDwPNgZQuyDH8m/A4bZHXsVX
254ffm5ufbMHFrZIQvzxNdncPlYPtZfwts7KgWvAAOJy4aPKaFKytjvcZfJgOjpt
THyKc0QiH9BopjL8x6RxHaePHwXMsDUwifcBGaWUVX4b+gy406A2f7NQ+W9469uB
F3qaXtSQaWfRroyJfWtPptja465foP3gpLbfVpSiYZhVFS807dgEwjqD0s9Zoa2T
AtUxdX9I3+sx4zVAPGWbyvmqwx8kyjT3jD6iD1IruMN1NvDJbNVi9hp7wb6Cgu2i
KavzIcE+CAAsMg4Wa8gAAyloqM1p0rRNwI0Jih0YHEO1NKWLEAyc1nIUVcRtLyCS
XJ+thp4To1tUn/vxrQ8n1jYH84vXnyNpOi8AYng2hC6IsWogWL4GRXVclH6WSwFC
+su1R32BUTb35LQULmfdJ5vIviIPeL0VvQ3QZgaVCl9kDYl6y0AbgWnSq81qHOXe
TdF2KxrfQjFvPnl6L2FF8U83bDnm7MQGJ+028Jyq+vCsyh600EqbHyTgUSOd3vKP
MzrElxkehZ7mdNj7LpCoddT477GPGjGun4AZikEDnUTNMMUHofSKWkO8N5nBL6UQ
C9zHwbeegekiGqjc/Gp3F+wnpgxaUJgujDmNtZkcDVMhryyobjoHInpURbU31nEj
l6LR6Lo7Pb4WMqHWTCiYXyDCJNN2rw9zw/j4WxEfhk3NTMytYtEu6wx4EC6m8UpF
EBRSueq33UsuNd4SNAi/R+fuBgbPiAGKKrLZbjP5/IDvvtK7liMGJEcvmyRC0m6X
xcLNgNAcEvNcPTaeCpdlE4nX/t45VLfrYUTOHlroLengppnh2TdrYc5OCpqbZe2q
Q8wj/wQ+mkAARpeChG0l3t6iXeUBoEVIBADUj8dsj3FRLkcGSwHEYC9CGC2HAUMy
g7MjXcjM8hSjgZhJswvb1P4wl1NYlxhfUt9R12MHpugumtqZcRmbmb9IV/S0RpeI
nwwT07olVjiPe4KI0E0vAQIbgWBu1GYCrI+HExh/dGb4CoPxH20M7MmFVXfzHj+8
vamAv9Sh6IcmBjqrzK4BW3ugYM0gYr/W2Hya7yJ5cAEJxihQwmjMW3q5RK1OqxIc
prudJIK2Zl+VtgTINinKIQwnxCXaFJVQhGvlQdWmud05mQzuNcul7hg98iKQnfYY
/aysnTlHD6WTZSh4kDv/KgeuLfB5ETOCgSAW49tOlaVokdA5oyeJqsYOGZjmGFnp
9RRkIGfOnLjDByH5fBTeVHpGPjYppoGL/nsGrn+JSxmFTtQBUoUZifVLxrb0TTBs
Ml7atzYfG3o4enJ6e7enHdSVdgvrTZ7luiYKFaCZV+7BRmsCNIVM7ezdDOsgGCOc
57ENIMpi9EgbwN3ndO9KNrz1MowAF9bFZIbRJJ5vBQ2c2wFIF/82bk/6lnEtVGUD
Y44nhHEqKlW8UlK/evHcstyd1gS+cqqtKkpOWf1XQPMv95S+Pw/b8AhI/T+MtlPq
sadyy09z2rrvxc7B8DDi0EpsSKmLPaWxK7sEFwsfe+newbdvkrQ5uK5cS7D5jiiE
0P0p1SfLPlFSdQpYoAvBvTOUE4oLQCe69gs615ZHUs576noazF4mLVBLOuw7J3vo
/c0FX7zvu5UhFuqMxvVD+i52B3sIoJ3Aw5JbuFZ6MIKxymkXBuN/zJMKyFmPuxS3
KlGmksr7N5PAZjIYyZkKfp1q3r58TIj+/zyw8ROsPSB1Ywj6jnBcwPWYTRzhr/k4
rj4gE78SKWt8L3Qx3FYho6hWlzl6pN9vZpMyguOR24B/+AE1LhTZjwRRVgn9w6fo
Pq1AoFLGkUuEKpoAwlWLyFQKwQ3WZrXLTSjKsc9RrulDjfwcJ3VCji7KkdSRwqHs
TMAuys+TW8Jk428AdHTuo7aXWBAfZpg9qnyFVX8PgGe0cmc3srhLoqmY6q4neveA
iyqtEmYSkjmXIj4g5FM+Zvkic+37pvvYGYIv6c24BM8kBQZA0bQ73OgsDpFuDFTe
f7QBnxffC0C6Xso9euK6NUHQsxHW0yVqMOkKP0+KXu5ta4O2pmy7AeFWvHnEPOS3
lvDnNZC34PPuW2UM4qWZ/H9SypYfYy/ij1DrTGH5XR0YDmpueWB7SiVLjQ5WLb9H
R0A+OI3XgXyRclL16pjBvaursiP4HOMRrtkltySQULD/Bn9lJ2iJqu83Q/HI9+Zi
qMSZkxvLzGkBePF2iEzeO2v6bvL7pDnmRMw5YbmQRRsSAzhpOFcaLBG3AWWG9j7D
67yolRKSwRZudMhdT5cCSh5oLlcD65vFTeLp9GgoHiZK5cEgGNsl/DObTdyBHXqa
GlxZJlj/8wb9Ky0RAAuM7aaLISezerivXHtiXnE6XPDRTmOObFUJZ9JD/7xHA0p/
+q02+CFTuNSVPLorcSSmIJqdirXQkto1eIByFVn7gol31Ai7YPDACITItKx4+eCm
xNPDMeT8IokTMpeEMnrcDlKpTCp2rxn7V9jm3Qh03g79atAXjBUVqLrE1pWi27xJ
Q2IhCkQI02y5a2mmQE6fayzpq9I9KiXUqCuYpSkUvcgClo/FEhIMr5qEy+m4sPL5
4f7iA+0VvWmkr6CNcjxZeswbDvDKe2pRHjAXM6TMmEUZkwT/oCS2SdxFYq8kSWOm
+oPn9VudqQTuTQXjaLTJIWvmAOkAreoyDEBums0H2Xy6d/bI8oPkFy2FwlS8vtpa
opwWrDYlclO+QNyuXcRsjl+mibuLjLm+2XtoAed3FJDKCFACPRdB37pemU0xbHsY
mE++C0NdTWVRj6KYLqmE61hbSpGaPDPVY/IsRx+n/87eydaHjU8crEuZU+uiNJX9
OQSd7nXMt1wDD/nQ4g+el1ZRy8tgbZ9iBGgD0VctYC9RbZcJ1vJ83AG30vYHzu3L
WHicGpDYirQFgxGV9qzLojxv90eVbikrilELdlDhEXOAXMCAXeTIOtr+EwWw+y7q
t6rMdl7rl5nOQJQA1UO5iy40XncW08Gsdv3JZb6RjItZK3lSNe94ngHT7ZVwkbVJ
E65bb6yONNQ/+HdLjR7Q3iFmBTZ81jm9b0vFhedkUibAhYLLKJwciuIsKJTWGbuE
yD2p3HVR/0x6v0fZXGRJCR7OZROpdy0PwOk5Oj8U4IDBWEYUVR0vxkog6Kj7kJQP
lnjSOuhv71ES2C42eO3d2yXLipe2MZd7U0cSc1/An5EUUHBUDcTFK4rgfJgLpGG2
WzEGXgivzXz3Bmq059DAmbPjKuTPDdWneIGdmF1BEGe89N9O6ltWCKRCGc6s9LbF
trR46daOoInhSZxwDQd7xovpYvv7DnUxsg8Fvt2SXELhCGTh0I2UhPcCgpEeq9gj
2LGSq0xgeXutqvw0hU5bxu1p1x7QqTUGqCid7iioaiwcEAr4UEvk4MrmsYHWseWw
g0/hmhWExM4kRSNoz2qolWIvJqqTz74NrR+jeptPokLDuf+hEMwyBle0E1P/pjaU
oKy4pbvTA5QHv0T9fJR1g62QtBKu/oWu5wkJ5UQf8yb5SRGU8Z9Mirh6SiCtUBiM
OZx4VVLAgXdP1GZaQ4/vV7Ev8DnraD8ng/LUVMxdxJYo5CcoFSAfY2kzYFQ428TX
V3OLynMPxsV7G0MbgFTVxMW2fvFJxXNHjdzlS9FRlMN9KuKbLuiawercNJLm9Ab6
jzJmy2L50cGCOUg6SjABHQ==
`protect END_PROTECTED
