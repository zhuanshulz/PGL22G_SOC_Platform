`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WD/iPnJhHp+TC5Z3TA9ys9Okweojc9PWObKuySw4Fmpv7wgMtqTe5QKXV/AWeTwq
Be+l1wdZgmxOtjWdDXEy1RDUJ2JCXjD/XktFyk2MuTb6A0KYDA7By6G4UzFCCZuL
H5Hfh8eWF4aa1G3Gfb6o7+KCVOHRao090p29BT/6eD9WQqZJN5/f+h/4bCjqbxI/
tWP8eHD5df6qAJ6PcIjVCAMkTJ7AeLmYk+NeB5knX8xpbO/pUZ5pubDjNrqPN70j
N462aAwZ+H49soFGwvWlZlY8z0Eks4b8uYLQgL6YMeD+6RS4mizQOd+FZBT9igxm
Urk/YptfT5I1T1/7elh0pzORi8u0dKBTTAfV/vxVc6W51Qznfw7y9c93P1yMXyx4
+62T90sgrqEh7tiZ0ML2vQ==
`protect END_PROTECTED
