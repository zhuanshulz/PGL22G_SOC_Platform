`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jJZNDaio3c5ZKXnCLGQQyj7fw/J7ULIkz5nMn96daNvcVgDK31lzOctpEkjY3BjA
SXrBHNt7viXjNGpMa0sh7wOLx3tSFf8XWAt3IIWvhZC3WM/d6ElZhuHWJEPgBq6c
qWJKBp4Nn9tbmI96Sw2LRJfiPqVJMlHyf4S1AxxvDfjPX+YdcBeKKM7WuvPWq+en
fg8ZI6AfsnobDlmlhbguAS4TykrgeO25Oufxxuuqquib3uGK4QaGWVSsXg8gFCGx
IG4UKNpQX1CKR7q+eT+SuE+HxuQK/lxq+jST7WENejtM38APf7qMk7/4/eeAd4j/
wKQ1dHs+MYhRojCxnm5UkjOLExUsG3+piUPs9FGktiho+BUar84n7dwhei7OPWTT
KJlZOyBdabiygbX3l2WrjELLoF/k2/gX56FUpicU8rPh8KNyv+pShC/z1LTqBT7k
fhVToXtR29BiGLT2HWxvw2RhJsvttvd0uctmgdlpTYCGZchdtsqLYlr3VhriI+bK
RTR4JvcsOa9UQ4KA6qrSULX8NymAo74d99T7l30eYZ5i/qSSDIPJUM0HXzIZg37C
8dW40BmmAgjbVKUcC1NnWQxtekJxawPfjfSgQ3rPjSLQBzqYueJi5uGlik9xhwyW
oXRYpDO+MiBlyU0ayOpz20HUDQ4QHuTl33prngSoMZryKRXfEw4GdNyfPLv7Ujx/
s78+d83pTYJnLgUHBEBnwbxMyZ/STZAs42l+XqiIM5TJBnIb7Q/v7Sl6ct13M0oc
D4Eah/SLJf3UlDbpKy5epdyS6jwekoQiB2KBRG7/F8Ik/j3pGKRHSLzGu11sXXVw
+O5a2M77HiZRlaPfIZx4WVjEuBEPY+lWAgw7hXZ+LkZHZasxjMwkkJLQt0ENmjn/
wHB6/K+VRWNF0D8jpKBkwxxL6MJML9ZZSeqmyejHMSFwjSDqKSW9BK5Yh/r1gOrJ
6pFSHwP/PMjfboXAiKvDJb1ORjuUOk5nT3IzQUCZuudPL1SzU89wUF9j2spliul0
ZnGBxA6z3sNKGbL/QmTH9w0VyLDIiinm3dyh5grNusf0m0ZiPI7SjgA4T9Ascfq8
XgqAwYLOmrTz5QTRXK9ficQmP1VHNfQuevqx8IRczrrgt25B5pU6gNvZoPJkx1YZ
72gL8csR2MQSvSt6S+cBn61PZsKHGikufK3R/QEnNbNMpIrPolLv0bd7YFOcKrCZ
o0Nzs6O9JfUgxU+D6PQQTxznxVdXaAdSylccrMsLfSm+Yuy8/Sm3qmtMhAEc0NE6
Y5tWdr7pW37ZGHiAzTsu9s7UJYDqXJoIM51mHmICxmyyYLEK4HQaGYYuVjyWGR0u
f3kFDSTaWUHWpLGShR8fGcf3eK2a9NxSmcdtGtezm3z4xtaYgYsS2bifPbHc6Ech
LJy+GDVELSMnIV0serPicoCN5sOlSIMjLO4am7YHwzInUte7os5fedw188M8Wg7J
Nk59L55JfgzIVraMPI5neq54NoN7U6y5lc+ZGtYLMTVUfnrLbNe5cmJ0oojx1jSb
ac1wutjC2iZtWYU9syUAUcCZIH2HeurhvrjwwGeFBNgDf7WTJiLuYDbr/HUbwmVs
gXatXjCHGNobtdeevMcU/d+1E6rOkqhQVtmtaNwohm4953jhQvcrEg5f76ZzfRYi
kQPnYZ57u1O9lsIos3gTGcB775Y/gzBeFD6eSqexW8f8jbpUY17hnaUAmf29htZh
qkf1Uql8ja2d7X4EZ4DSlVYpSYiWmbEWtwvmTzsXJSqnBcCK6qRtT8jgAc7fSw5+
jXNVVpVcuv8wPRXFGSZQlPjBL6uqDjX4q9GpOnW1rhp/X5gm9PAZGz94uqyJzZg+
0rqL2WbAnv8RulmmjO+4mhzsPp2LgCiXfjZmcXpKX5NinEYfDTn0KTim8owfW4n/
/VxJf5xvknWfcyYbRNHD8Xvv7BgpH612mVOKbwO/IdI/MDa7mZZAVoHhceXkxrcV
UB+32nH7zYVw+j99k+l06XxjXHYPtZoF/ZMAXUnsDoo19vwne2H6qIyqXjf4MU2+
VXwJI1mGHLCwACRzv/X6FDwI6lanOnr/nc46DXGqZGgIM3tS0Nlt3HjVqyk9O8tO
DZHmzTQbWjTdEm66tjC+Fk/1CKGGHUrFNmeTLKvDEdG4+7Z/fOr/NQpEooSvfbi+
6cLVxUdMPPipIpj9mf7uVWtn9LQWw1L8dAfLAzwDJKY=
`protect END_PROTECTED
