`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
byul4wbk3UV2YDchpbUEggdBfMxX83B+qG4WubW9YNS6ESnNZdITJKbeIpu0us8Y
qWTDFVBc/UJVlFfmhXkKa0QDKoPSA77RYbHaH4dI4cpw+jCUFVi/xzNEefp+lt/8
t+rXkx2nXrfTo1XMlOrfwvon+mbOdhKfFdDVbmaMHj/FBoygLoBnzayQ3xiIJrkJ
edfYAT/oYl7wi5DJdrvfbADJGFRfIDEDgXd4G0qlhtMIfviet0H0puBAFFudfSQi
5tn1UIrAv2jiitip4vUXmwJdAX95e5hlKGcKPj/Ct6DrhJkly5nU9prYYH6VclgM
gZhbx3uFK5ozEmvx+RBJYfjom2ANVQEiNDXzhSNLHLZWRRiISeuebufyMroSob2V
dLj/DbXTb979ywEMfrB1uED+3yg1dvrTTGTbuxqqf1hDKel28yyigLLWcHyAnPlQ
lxEqEVUFT5iP3ZCycwSZNRJ6WRhek9gQqbsunWcRWg4MK53uyntBk8W++l22wrlr
kJEbjw4Ck1t/3CRSMJjQg0IDCUP2Zz6KVCnLpwGVzaUwp4MyBHMy1hHw1uw3a8xd
pTgay1AJKaNuF97QUdlenuBGA3GctB165sf7k5ruI2mr4Qx1TNKyALDGW318aDOY
3d/n8F6aexceINvWPLIzWTbHmQjj074q6hoM6CSILM9bWVt7DxKYPRm82Qj9ePsu
rKZmoc567vJc7P7ADJy28MI9Qn9ijg6CwLhV6BwOXyL8cAWCWbO+x9V6HoFYeZYI
VqydWp6Xcx2kSeaLbljnhhkYb8dCD2fkUrnsnSudaIpQqejtF/bRFJdCdC38qfp8
Qn2B8HoIy5+lK735Bhg0Ohb33jovEQezfRcK6Gs3GljqN8urhdsdAsziqUbfmsF1
wlrP4otPQPBsmV7Do3X1IE3rJusM2PgAouAUvLuYmEXSOLtvL0h441PdVkE6PxRw
qygCEc529CzrDUSNVzxf3T7KsyGYE8v8wMnGR4sI84qG3e4IelyY6lIYaJl0rQS+
YU9ZPPw+lrd8C67wejZhDTNfswyvCRsIs/he5QIsKqwUNY3HIcv+5lZmNFhI7duP
X3Q15k8l9hnDwhlc26eF218kb0ysJ1F6pZU6op2j1Q99z9sVTLLwTQxPiHZtdFyb
`protect END_PROTECTED
