`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gM/4R+gxNjZGFcTpR/IrPsMSzErBtlEZWltMmVa20dh44F7pV86xJWZhj0hV/hDF
MdFwET+m1fiOWOHwOnPgwigG2FNrHiay3aOOyHG4MA0nP/Xs+3moSy/SXCZEbt83
kTIkprS8fJfG9Ds8B2XV9vqmdE3bupYjjKqx5mrjgAersFuV2AtIfddcjHATbUXw
SY3HM8vSPLB48MILr7T9xb7UjtNMgf8asi09PKnjTjlppI3wuDZS0WyKl3Rhy1GK
F2f/MCarHgp5rZdV2PQgU1o9tu2zCLOmPbDBeMjXwORP0/5O4GeQdhfK7hxOI2YL
jLqrxlfl5hX4Q4qQMWJ0bnpO8LJr6zlezvmupnogjG6dGCN7uJeY/0qu8YxwjpJe
XGUOkWVKwOuOvhORiP+OCqKxzAr5slBHfBntn5FGvR8wom5nHuNt9Qn+lm7xKPJ2
6mK3KuvLldy6O/sz3c0gfUo8RWkxgB68oVbupEv/PsaP+ogiWIJjtaLOeKaVK3aI
`protect END_PROTECTED
