`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sI05yb53Rtyzh2hu3IQAAsL8HU5l1zEFb7VKlcZex8/KZ9TOOWevwsqS683xIvWi
ydP0tEdkNZ67l/TwQp2rpxY7ujq992P7dwk7/4Rodov4wbxTVuuB41UyaRMhrKUr
SKIhxc8ZFsdrpMQ4uC4Ek5yeKgtDyadeDuusdeTUneYZdHfFN6jX6uki0uvxM+2N
7UkZosFTTw6dFPBGv7ENx+9KMTs5Jt6fo0calr+kjweehJP6JfAjI4T4tfdzIAGL
tPgH/uZlR7EPI2u9bSzjT2/oLctueUI0mM5iX7DDPjgD0hTu6ZjuiUmKLJrNaC2H
wBkDsn02utnq+c3mMFcdokOsn1aunpmmeBtejEN9iD4vxp4S/VGOUEoyiAlqxcva
Iptiq3MUau4r6dPx8oBa4cv43oMPH6LX5OhMcaJLnsXRbId5RhYNlxEPRIZHJMg3
jMV0YOSYLtApFJx9ZVMVtbBvhwecK1koGJr2HZR3KMi4NQX7PEcGRXsliG0YVezU
FNkK3xUXwhWyVd1jv+iFSKs2jc8OW07hlbzW9zzRkDTG7hiQ/dpA59uSOMnMzSmY
sSxETilyELDq6e/iieadO637U1NcJtRkT/gSKjyM4nou5isRi1m4m4wkP7JQiKH8
0m9GPVMzMQM08U06yoM1L+WoK9SC5JKNqTCW+cgYdKBkWvAqEI55JYHHXNtCGX2U
I8iWyg5uTqog321s1WZ0Wo8q58AbI/Hxx2ifROUgQcFQX4j8zVYUERuJ+xUyH7cS
SXVGcEBpGxmQI63bkPbVLDe4trT1O2J/hZq9nxRBKqMLH0Bz2f2XwazNyHhIYUkK
02MhhEBu3T6eZwfJAQcMqoHrFPolMnb/oCn4jrjUTUUK0c7qsgicvC0llK8Eeckg
1r86DwIopUoK11SRMiRZV2p6I2fAtZW9zDpvaLXeNb3YWFdD1ihUGTjEfn78nsRu
jp6xrJ+YoYKiNQHkFDexaGNthzMnrbmu9Wg3J908xicJsVxABk5f4azz1ep5408C
8bCaDMSUB5s2L9kn5mvVKBSk6dKWl+9JWdiAas3KM0tXVgofVy+koUUr0FlwtU+C
blr/iMu8T8Vv49aYwrnCq83jJSCyhunOX4igaqQATeP0MDQey5L53AUDwOGXxMnI
ILgtabdXeqYH+oJ3woTzZcGW/MLBysuDYpIxtOZfFYrkCZeOMkM6hSWkZML3uzPQ
JPrTe7lpHVD9VHAZBDz3K7QEgm0KHSXhjgZ6hxzS75d1i3iGDgSjTJF1J2YWNvyp
iNMHkGJroxjxiqOSc9sAejaffxKFWAx7DVQ2Esh3FxP54++6DvnHPmRSmlwE8OGM
QvhcxWCrRmxxdYmema6ly+LW64UvrRcbqHaIJyHstn5QgqLHW3S9Kg1RDy8NKqvB
OrhW1Iw6bdd7TsbEGiAPZkyF9p+/kKn/SL6V1mpsKLuy1YJASYhlrsxHnTnk2HJi
+kcmuI+3q2ViIgYQhNzQibszZd4T0lwuw8log6mpk677i8rHI968eiWL2QvaEuCc
vwPD/8X7ZC5y1TqtTf5UL8iA5tyeBJEeaImqA5RF8Otu8JCpJgvorSwJSDpB+OxC
WBZTSQKBHKO0sxlNtDgR4UiBAjgBh/i6ILrV+/CX5D9A3aWZ6bgR04u3y5OWyG/l
JYEOZCubo8oMsfxWajbZIa8MI5J1vVH/FkqNrtTkkE9dfONygW0IvjgpT5HC8zbP
FF5jCXhcc8zTIu1kxDj9fJlCEKfr2R9WmuUisOOc3Dmgmwa1/SHZPVyDFy+sbvt3
0gmKOjKfkooqHE6nAV2m+p3URfMcl5+bfEEhC+bq39tEAjt60arTNCkWoB/qiZMW
tEGRpqsfCtB19a0QQam3AkF+sx1PaB3rKRs8BJKWSsqrgiaNPbmjP165XtcdLyz7
EDr7XFTADmGhG95sQEuKhF9YzebV4qoPiCfeSVYABmYwBQzu1xyxzux/AIQsgtA6
jjiyfV+TpTHrxkSQRiUyqGbNtweg6OUctbRToH7OywWk2zVk1jvdl2Viz1ZgD1KH
v9AA37d7q/vEBZiYudvzT2UCP7Vc5qvR+NZjt5oaN92dysqVaLQpQHJkutpzma00
tcgtnV9t48B6vqgHe8ui2J/0b7tOxA1VgpXlGnPM/XREYkRNXEZKiwx6fo63P8Cv
fH6e/33KLCkP+yubvjylqwwiCo5Ir8fTSqiXnPP6Ruqb5BMUe89REtvxdJHXsSU+
U4NQENNxJsz8ehPUfGOkKag7LMY0O9FyKhEKS+1tKtQNQPEC1dExnAoRajulBhJh
J+vlxw6Euxnstt+L5KoSsqyXns8hJ8qjyWxMjPtNeiniLYLjzQ1lpkhIdbLLnX8z
mWnWKc85iLQE8Fga4Yes7l7XbbLElSAs5BHduPYktqiJLAATNXg9+njnppQz0dD0
z19KMsEiDyBqs/FLTWfk1zNUeuK6DvhBbm4TJKlckOdOO+wbr59l4pO9MYAXmSkB
h9NC9t8xdIWcnsTd4GYv3or9uXGy/2z0MPKfvR6QMZJ7SyEbEJC6JW4alynKZB42
54gZE/+jhpQrxuF/eQFHp6ENdE7wySg/rbRPCKbSCMYKxbe7FcKkAkQ8rB9z/Mo6
uLMCi8k4cIeDYlZLZfRBMPlsd9YpIYkUOha4iw+WsubgABijvlZ03tfrqebWHyYE
zxCUgk5rnGe6drWtF55pkosq1zXS1Ny4NBmH7XhxD/oRLkkI5hkHUeDwnkjWgfK+
PTRfBvY3lVMNG9Ly8TJxe2MYhVWlJWNsvjmHPQH/cRM5r2HFycBUYt2JQqQhpNyR
7JImjMtuEzIkoHZZAcz6qsW5RK8PBmv6Buczrb4mKy/waL4rg7VX8wEDHJSXZpbv
afTvsnqtqjjSUpVLIAW8hYho5gd0/O3d87j/Ff4O4G5BTusChPi45wq+q01JRZOa
bEV9nInKyLLDbf+R6Qae3yO2dwsKOlkTbzcoQepMQldLIpUebebq0qqfJ/EMPxwh
oPoIOIn+M9iaO82izF5sxzj86yKRZ4pa3vmRZXHssKlikW0j5CiaGzmmJ1xA7LLc
h1Y9C4qL/Dm6+VqJk0rx7aIG1uDsqmeZzghuoPZaD9aaa8N5NL0LgqMmNzU3uoAV
wg1o+GF0CTf5eXbbjZKjnu7OeKOboGL5B/Ib4Dyy/JotbP6RieNbNdpi+l2QShQi
mlpGDOzz4NypgWZ3mZGqvRYPZGB/dpTu9dPEtLpsOsLnZP159rEtoGE5hvuttJeO
FrVTLm5nG93mbnzDDb+RRzCC5MUY5/HKkU7b49S93YFBloUKMYlLSihm82mWWVwM
751M5WPvSzqz/hpjxVci5JyXQ6WX6YrZW0PbM2uWlSLZHhQygA6CzlyP1ZbhKo/T
qqRZ6qL2PpLPV/yJi5sAjxCzN3W/uFsXxDsMjYkRXaz3iFQni0+94KNNsV6QWz7D
IxFDZUncJWxesxNFCefem3x+RNTqubKystcjMPZPEqcyZyLqYXMvAgIhF2+1PJes
khZWVaFLYJhBw1Fub57UkLzu0uNTGGNLcKk9T8p5lr1cnihnPmy3yjAbS8xMEuC8
DNs/vkm8FCBsw0QmTK4Y2IkU7Nn1fj7ke1kzBYEKY3Ht7HCuWWNWydQvclHhqlKh
z8I8Lp7tdNgc540/VHjriCcxPqDkHJQDOEswVFmdCGxzTGoKk61TsxfVpA+SSau+
8kU456y8vxQ5uDzYSeRm0PRs37vDF9qkrxXbzzLR247KvmsDLlDWtQUQ8GIdhND+
2wCYfhj0Ja4RJ+XU0cfeEA1V+xTf4oUy9nUQhl3/Kg9A5b8W2DkYcE9sYCrhA7Nm
tjEdG+qFOrz/ZWM6uF0Ivo3lPzt7/2HkiOMw1zIAOVKzfdamVaKMxRmXgGKXoVZD
R4XCBSpFlfTXz1im+HaNYJY5SjWl8Li5ABhYb0pARPj1wIE/iUhSxGOEWEkOMlMZ
t6JBpco8/o4se+YyXKJ61jtkUi7ygqzj8zTg+sL6YhXUYiCgbKZx2LxCp3+ZKBrO
24yrCvU7frcGQ/xHfCdCQQl5YXzVaUDtGzQFC5stymV+7Kn/yQTRKwU3Xn99dFb6
Fdt/6CUOzbSgQBOBT90cbN2R+WWyme3LjqnuLuokuD9ZhA2jO8XolE36wSkBXyM7
iR0alKvU/ce+m8oLcctxNKzC4SCd86OjeXQMNjgVev8luu7oKMDwqyTQN8hAHD4H
TvadEVjv/Z6yS0jarNokNXBcWTpWXGtWTGS0uZ6ilolgvmjXcK58bSjXEKhw39Wp
w99nywla+mOqbhAy/lvAGvj4+5bgd9qaoA/A/TV2z9eJ+fft54E1kjLmRvJ92RGg
xbmHDAMRjjF4a+eWbNhmY1GzHjncVkV9HqvOEKDgGX9Lqs8kmjTvyYlBqqHr5kBW
PJgFiNuCjSDRaFjh2VeNCR8drNO/98vbYcBMek9wQF/wpl1hJD8stynFQ7Kmnq6M
LtA3KWOu82GGofLoJ96y84kyL16jAUPToWIwaBJlKiulH3pHNJ9nH+JA21170JpP
DI6V5JwhwMGcHk/AHagrGcrotxcqOWmajzhvyK8RNv4b0J5eC++m7sPwByiKnRCF
ZLbTEtgMd7sUAHoh5IbQx1BhczPxnaYR92C+kVNTov8cV+w/ucZlrpeSsLndCDiF
bQxzXkQ0wQA8bup12RIuT151/QNERwsgkmxP/bFhXEzmaSPg2vxwejFsGnk0oiQg
JucpymhtTL2N1jMi27wnlb714rkOaxIfHJ0litN0vWpQptBJQBAcDIy3l2n4Cx2C
8DaDVOuZnGWxnAdSW5U34EVmpUC6RYGorozPm+AILyZUfvlYLpHU/rlgb3TixRK0
M/C7HVMmwal7CNzChFnv84TJmwGIiyZ9wBuFe1X1S+uRnYB2Hv+tvV+XNLBu/oYK
DsRFURKGm2wwzgHMVlvWYDaH+Zr7H15ON4cwiQLCxjwOO7iamOGUTXYkfpq1sL3I
1OmI/fZVsf1Ae3NQmchW/6YsfEBWbd1iAhPJ5CcI8tCx9+CsHkd29xCpuxAPRk/o
05WYnm/428U24fJ/hu/3GCt13cI1YQtldHBfGqlK5WJrLUlOy1X/oDmNSr4dR5nw
otWta02Os5y3zpfieVnXXdJDU79dssgucjczTy39LJ88Xy0yjEyCzdbOpvSJMQFc
qi0ATRrU4Oh2X2QuIkb1l94jKRJ8M23MeGZYnGPihepvu2MOkiKE8ekeHjQeBE56
Ucf8mhK5Hnf2OvJM2gsAgqEw+bGa/4SkLKehelxcwCjRm1VjC2BGhauq68HQaDfb
NUBwzudpLDnmhtlM2ES3ENQk0fAo+Oh/0dG9nFQ4eCMsAUpj9VJGcoijEXGeiV3B
nZytKtGD1SUmpyVgAHY7V9dAzU/tlWQRbzUGycc9JD6dmrjfMxp3CDIat9eNLtr5
PbOyp+v3/IVBOCxX8YwpQYpox14wjrl1BOFMhDT/JQXVM9oPOcJc6zJSpcqR1dea
TozlcyQaSKmIoudcyFSW4ZsbvXhpmgRMvYBJ0sh8FvI/WmRe7HOdOkQ1O13JV2a3
NIL8yxpu7Ak/irp5XHPR4zvLav4CpHv2xtF9F7JaUvA8/+GS+qV9CSSL3zs5QIiv
LCi06NFdP7kTuqY8tLQM4YMT9MS/SEyO2ZgihBUKF0R/rGdNzAXHkXWWIv3uKLkB
1sLsr4Irx9B5VPhaHk475pi2lCt7jXE8oSNKpTJIdGBRv5e5WJ1KonI40dTZ93zm
wzbiInOzd+cPoawwllLjeECdjkK81BWg/hKqXlslKs6ean1AHABKOVZp9CHgpQR2
TcWexuyWKtklU36CHnBGrBMoKXmvVWM4rB94vWl2vfEfViz9nlhMAqrXLzgpX2c4
2hRNr+r0PIRf330ALdE3TUTI3eknKwAc3mhpc0xtatOnKh1o2TzptiPghPuR+XsZ
wUSKf3uxtXckQtF9ryeDsFA1mYd4YsfXc0Y82Schyy12XF1FrUcPso79GuYc5yY8
KjYuEXw+avfigur2cOIitxkZbvpcI9rwdPDbo1gCznDKLIez6WQPjKKCYLZ+4kEI
N9Fe26oWmVbrMDDUPD3Ieqwp4oD0fEOjwvyuw0zytjRFJHz0guIP8fiOg8oPffsz
zf5Dsytyl93ZSWPw2eO/3/uoufSK+tlEddqfUNLZWpCpkv2/WEBoPgHF90jTVtzZ
VnxjgyN3qlP6wgTbzCMQqL4eTopFpb2NPmUIuMNmpsnXUGlq4UYWYc2VyFyrSUXA
3quvJOWAU5GoCq97AdrlF1TmCyh3yqFslaw2Zz7yND5MIrvFicn72vpw7jfV5FxF
CkqZpx0kEP11nCqLt6s3Su8ESYb8OKRok4SbW8L4PNG22nP9BDP0e032vh/8C9g4
`protect END_PROTECTED
