`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IhQLHrtbAJEJCcjMPWKwzpE8wagXsRCi718gmBKiDFLWAW1pTzV7NqjpC8f5CAXK
zjCtx32fJvFhczrkqXydv+X5sp7jWoxD58YPbyznHHUziPZO0eCo+79YQB03ba1u
auTga0yKGHN1CljgAMTaN0zjkHB1sn8fR1tFxwvpjjtJ9oVOrn27VZWTmPj2+n2k
CWiqCbJEZ1uP9ReeliHJHY2EQ5gTyD3jZRcpLcgX0fX2sX5HyD3s9COAqTuLu4fx
vl66plbmArCD/aR4RnrBDZcAIEP/lAVdzWaxJxudqBlGfbbS9xFjyUI06nJVX/3n
o4NXWiMM3dGpaDXRKrg6hQOEj7dlcvZWJ8vRFBXCqLaOWC0+2mBZGdusImt/oHB9
8BcE0XoZfhYlzbDW1eSidPlDNZkKXnQKhhbB2SAIfZMXtnqLMXfGjyq4bRmIfsvM
AehOkmWDz61042r2GJplGruQzr74uE1TnxDTfdIUEOiJDBpiHyD2GUYU8rPuLZZt
hBV6LdWFmyFqo2KpVt4XlaHEXibJpGc7uwHaJuP+m5nv+vfdCJnYXmZQZH2zQOAz
v7oup9jqxgKZaMypQ4ysPNnH+FjGBDpTha9mqBaEO1kXzf4MzEaLGYG2xoVHFKvs
VdIIe5VLBpOFaPrWSIxtZktMEAy3+y1Bt+fQFt6SM9CeY59FQdrz/FJb3g/lJ5S2
oKGJcdDzxu0keVG46Ep/eCREP4uGbZoFhzxxayMXPX5XAs0p9w9DmMksGCdURMbr
hw2mJmHPCeZH/kafMVXNNUIU7XSVIGrTRvLaIl8VbW451LwU+CUDUUT3O4SgnlJ7
mJOdQDen5anSpx7b0SmKkz9Vkzl4PxYDLvgbU1Etyz3hx0zDfWNTHb+i9dh1vGiL
Ur9T8epniY7RmZSKJNxK6PbJFZ2Rxr5VpDLnMZkiI56V2z04TooA+kOiwA8PYx/8
UFzTKh9eDRSEXz+ovz/ZcktY1JTAdLYAKJOL1R6C2EKHkQ8J8+t0UdA4BUGgo+FH
EAjjimIH95k75+l8gPmMHeOFP5XalTVoB7k+1yHbLAudZmKCYT5xV5+NDDFAU61V
IVNrhVp/zcCmgOI2qg+ob9FgDTrSH4m2aOJZaRZ1GAhxaAQ9tH9PNFiP/uTVNGIw
HhcdjApeTcVmFVmpfSMATD2GYumI7VE/1JDsiYPpfh+G8C7ztPlUIi24svamuQEc
lx0x8Uq4yqzYTI+KcBpisz4PxXTITCOGxFk6TnATAjxp3N413HnUV1+neWQ3syuH
s44hyBMsZchHD2n3cuhKvswctNMFfenJCMFqAe/A1DM2WMw6k4+VnSdW5m+5Sq98
EKNEjQDM1i3OO3r8njX/8mh4QwxiJJ+QXUoeNzaVq4PVbXKOkqxrLlobJvX4y5Vk
1CSO3MI2+2S23TMrYMl3DdpYk9Dh151jmg9ABDHMmcHfLBqOiRVUYqYlRYh+kQ6d
Io1/oxt3frBbNAidwRbf2a5QoQvS38CDEp2QD5b9qDGM3f6QWS7fB0wheu8VVOFC
fiW95SznhMw6EIsGYQLuCXROXaU3Vy13texVrX5SwSpIV+8AWQmMk2LINsL+4GDD
uTmkRP147BN6KOX0BZHRBSa7TcxL7KNshynYYT7hvc8UKYQ7qT2UxKI8VMEAb/HU
R903AxL8TvF0j6v7gbi/cdYiQnBMipyNUkDyctO1lNK1Ued9gVFcupmfneWwig8b
Z/jIcwVjgqqTfmN3bBMgSIxP0Ng2k5h/I8SsUzV6Yk31yuj0GW8DdBa7sVutZ+xp
pUo/4OKdeKWRwERgX7LA+wHftqDYvoqfHqSIFaWUsG8pgCmRdUyvFW0AXUIPQSWs
hoxHmkX5KlU1mBRKESp0Jy85VAqBWifBexaxKqMtKGBt6ZipdAasNfjJfltc9aa6
0jjzAea9rpL7JwGhrWu0vw5UYsIW6WhcO7fGQoWbCr6S7qrgwp8/Sg0Ax8KmA3/4
7bvLI7Gg8ezuLja0wbI9JF46A4hfvZVVIATScdK8xXyaEKO/auNT9eiYZCbls7hz
K8HClEFexKGf8dI2Rv65wMXtvBXwtDpmd5rovLZSqQxgTNlntE7eCnSNb6jTrTqH
1wUjLBRAoPBXv6SjMXr8q0N+pLS922WycpU2es1tq2N8ci8AYx/cfDcBE3WyDTCr
Q40tI+jSNEwkcsOzabx19RybOHq3tG28FAVBIzRGNSYXRzzZ6qjlEW2niQ2lThmH
+IOuj7WQxRuVvI66OoBKA/RLvxoHco9vWrKpXazRB6eOGrQtaF5DmBfEejhc24mS
g2O9oCxOjCZI1c5UnhC9wsBrHPsQTym0xLCxFjAkIuMFyc36AcEtWppU8ZNHLvcH
bTrHJFIpH4g3HnpBM7AqyP8RhlkFG+jRRZz2SK7mVn16dHDsqvakFCnPoLxo5HAQ
JmZRSFmW5naI6mz4XiCB0SNIJ1VTRLVj6yVELqg16vm76ENJfGgpVC/vloDf6QIE
OdEkJRFXMZ4kEjlZhB5dQYl5D39Ax4O8juhx0incogJ9SoLzSaeNWZ7k40S6pdl0
vRVsCnt6W+9NF0PDlqfyciwJFFT6lgIFWrG/wO0gCnFsMzi4lGW67X/Adriq/24n
vaVCZyiXGV2Y8quMpO/jrBxOtPRWjKYP3UC81Dxbtd/4YAKrsu6xIBjEptI22N6G
B+WtuBZh0UZJ6t7L/h102ejHOM2qltaL8Tu5EaWP87LTv/2TbAHBWr+6/oFxiO0L
+ezIVK0QdhhlwAbZ7408ZbyQy9+P57nZEtZ4ONehQeMOzHSveHSMyOs4zS91dk0c
P2510JH6ZSxiT1vGm30szvFZDg/8d0E9lhu2eWsRiO6eqI8aUCCUfKBj7GhSiF3T
DDU5RHckph8EcknYuwX2aYesNszdQ4QuSsORWmYXqL4D9bOGvGlR+W9UvZH1x7Nk
26F5xFOTe76jfMIgOLEyqwwb0rxDVjtTLhhB46znqDfR89mN5mWLZxw9Z75wY+wF
XdQKCvs23eXQ0Epj5syPw1ychs7oMbpD9SqbpDk0fiid6zEQm2PoYzMuw6G1sElB
x0ycGjwYIA+r2twinUGoZmofRrJZrgJSd83N0cYFSWCPnJl2dHA8FXVR83gFscqm
HHYZxg2C5DD3EWd0FMWeCSCrFjv44ovFswVuf+Pwv4w4ad3cNiDYOjrF9r50TWMG
pgSaVM7w7060er9m8eALF/hJ18HkY4eL1QIqefChuTU4kVI/QwOXVMtmKZG3eYds
8SEzMItVeop9vwOwR6oiTkUXtKqTJV89+31iavqLByNJ7slDmDY4fBfVek7LlaHH
0OWsqsYbefvY8d59RZtmu2EAPebRdvL7KzIYZk+W24bgI2x5mzTjwx5ve3XW42mV
3/0qBgN7LRSI37sGwEgAcgBVNBwNJkmDPac3/0e7eyXN05N66BjTPdJ133jhlkGy
tuXAPefeaPeMIg5aDitSOQLSrSOZyIXlvuJzsnZD8RuKxzPO76i1psNAXDo2YPZW
laiodPTIETi+97XACJOIwQrneRj0JBB4dnAEgB5XTYGjjZyjL2kP8GOD097ZNaPo
WpbJyyRQ49qyyoueniJH1XyldisJ7y/5K4NM+UciAfiR7TikrA/Z/FXhklHeA48D
VKcxPdVoxK8wNo23skKXnKRajFfCc42bbRVccjEBHI+mvaVEhYECWOJhiFiBJEeu
Il4Z/HO0c3BqdxbHBwi15au+qXXHkPgoya7z4tyHYdH8VQTdmyg0We+Rq7+P4eQX
i+x2Fp7hh1dHpXPt3RMVX+IlXiBxBSpzMEC3pQko0zMvbXT2YfwRrJxOxunHfDjk
ruYpXJv6QdgZy7eKnMb4maf1lUZ8ZstfRa+afakxnfv2HsJNID/nBAlfQgfzgWLi
nHhgCz1bZH81NK7/0holOrlWabyuClbxDFsXIsGgYSds8qj4X767+sleiUH64VbE
+30hXSBzoZE7+Td0oMEAohVjO3ZCi3V9gLUjpGYfmm9kUm6xIUoJj8nYPPglifVr
qP/v+qS83iwuHsaN9izLkpiiJIyR5YIce7IsfdhpGXjDyTZUfZxwc1aFf4P0fHVi
Z7SWPF1DLt5oWI/M8eBxUdPZ3NKglPZoZqpYTf4XIORxuRO5gcqSlUuk+MXX9zPX
8UuAN2uqjFqC/8cSZgSRKrY7IBJXSg4qmrp2QnGNuU0cLqrkqoujqTrbgA+9Uvf/
4yNphXvkiVZEBXygsa12p5lKeaHv2R9dkY8vhJK9IYLqnP0rnlWPss8B9SWWEGZ8
gIVXfuW8CMmrae28q2C0Y99RVEllqdSVXAVy+HAJQJRwQXZtn2sdiQzICVFc3yQQ
hu4B67IjTVBnpZnlKkOxkupUruFFdfVShAwBe1w/a9pqstASf8f0CFDX8tzeo4I1
dGVIjv/Pk7v37nG80POtsIu6TL2+iIOsL74skqdrqlfBJ094Lru6jB6seVu29b3A
yy++xsFUsJNMBNw/qrjgUQGZCe7+WV3l3diEEIGa3TR7T3Phq1LFHTPCTj6K8HDs
ZqLBRwaA9v0ym/E3hDlcMlUgb7b9BxD/Okv1gb1WF56vKQc6nAwTrHN9J2vt7awa
in5cAeYAleFpKq73UF7fMjKyW5nHOh+TQoGriMfSlAOPnxEex6Wf9aEqgIY+EBLD
QfexyLE28dderQmb1c8EDjk2dzp+QX9+BSpwwunwY4x3ZM6xVihbeLbjjpdZzeIb
/o1nsCZHIVZDZO4mYLesEPR3RtL9AZ3fQZBZjsgvnXYNd+VxCgavaVWEm4T67TNK
F+TT1QcuDAm9vsT6417eKJI9EerrprqVHMZtfttbN5Lkpqsh/+mjUx5MSSd55dHp
I3jO8qYje2pdCflBzNUPH1I4zCy+D1Rb4vTkblikFyqVJ+TUcLin41VSw6r0MvXo
TB51ydVdC94S+IkMHBy0ewWYFnjC8ZWMxo5pXXBoynnXvKGS4mXitkK1ulFtRBw5
xB/v1mhYpkx225K8iHHYSyVHMG9aLukcoUAQ6TS9dGAJD15q41E33YVsTrsRHSVZ
6G0iC9AEQ/2juyJ0E3To4RNMGP9hLYCEEqXY85kGVojVf5ZEyugExd1duqZ+1Dqe
prxYJO8U6XqXNrOXFUqSoW5ApHIlLTKuv9fqci14C+sGCO6HFKuhLZRHT8fxuh0a
UyRAmS4PM8lKVAa/kCk4TC+fwx69G/UIM/GjtW0E15s+lyjnFVF0uc7aNcFbVbD7
l6Hbw7YBUEhTivVHiMaMKqALLRAAv2L9ZbWlfvWeeAHuExeQXAMAcF+QqsMcDVwJ
iwg/Wss1xhvXUmCZqgeTVqGB7Am3dKX6fVfcxupemBIsoT5suFr1pfUPen9Xp1+P
vJ4adMp8Zl6U/nSFGPLc+ENzcxOrSeIgKKFyMu0UmZEA6fTDtzrCG4Ut/FPuyhPm
3nQVb3R7HQCf1Xl1gDEsTbM+INfL+BEwto6MozfMz5b+8LNwGv7XJguTZoOcfwqG
huxO2qLzq4QY+9zS+4L2S4FBEwLVgbT2L3VS/NBfKv8DUR4Xoo7ui+LV2THEXgFO
U91ICzplQnj4zlhgfoYahO5sDSb5P+EQ2FJLGKEtQ0xjaLi2xtao8kZN8rejEALr
qCeF66LKVMUsyLsT0/ztqAtT3RxQDLK4qpTg5dHczK1uK3kRjH/8phnOnDes86ia
/o4LaY6HAKsaXssIN4VFemsQ6xq01aPF8Q++QmN4EVWykM/MFA2bWecN2CxPm03W
rKka1Ak3ITs/is9/o6EvzYcKvpS1394pJYtoSuolqVx3iJl4WImLHP1KN60iN4j6
8AA0+ASJrhR/71XKSZpD5+i8Izb+qQ6qXfrnD/b7gIshQRU8QaMrKHMWqkYAT5uv
oMl1afSLOaC4lAAwANyEKm4gd4S0yWCmGrsEzb4PTAEokz3Yd8+4Qa2A68KiKo0a
2uCW+O01Ub7aOOeg7ygS9mOznCflVe0jReE2zcxd6a1oMVxJBhWi6d2fpLSROilL
h60VTv7j2QiCiU2vyoyKmI6oAVzZdei9e1xGHgkmLcomdIj76Ujh9GB/4Y0R3avB
+sY7ObSbgkAp5FDCS/m4kg1N6w0zDXBuKnnUQcRCyBTRwDx1VLD+eHmAD8G2llv9
pApsQENRyDXyNbbP6cFeCaLStCLLilv7TUlW/KSi3dCKhJ/2dGf/aL5wi5FlNO/1
hyqZrR57mUw5bqQaO6JuA3XdZIHk0annPUvZk49039hVuY7fLolDEKyoNVDWCLlY
ekzuqwm2Oifp3Jsu1Mwc9VHNdU4npurHLwu/s+wXpfUOZqXDbibh4VpBaAA+i0H0
jEt8roXSNvMUb0SV0p6yEaP8/mODUMR++hiwCt+AISCw7O1ApGbaLb6fMZqORPge
g/RZ0puz3NIMDY6wj0fquV9u50otw9lUMTSBmqaMsuj4GfWL4KPbqyOFYoUi1awB
JdLuoabEerrdaZBknIxUamYzGeGQJJmJQU1hYXwiNNoQAJe7qbXHJYMw3pxztomu
cwvd6ZRKhs1+1G8hx5ODkwOiaUjdzSZSH3zZjbsYvj0YPhZ7avelXHnDm/PyUHiv
lTBd117xwbAN71zOfAjcwnSK5ybKpmlSWGLVdsI27FSYqe01Xw5Ir+lsNmkg72eN
5UBYHbf2NAGrkP2gENjm2X8FFSEqKWSDC3BxbzFGmvGHIQCGnAdIbqoz066XH2gJ
oQ3GDIbk7yqW1D/NhGiV0/4ccVrFjHvHE0vH2H2nP1YXBINVyaoAE5YXnr7UiBFv
DPccgnrBFaFd6jys7LmIKlWEfAE++BMjdVZWXjerJsFXBsg2u4CKTAaqd5mbOipy
l3zdGOTOOk9vfx4vTogBqd4Vk548Z9hBdnqiW7DkJIZd3pckzxBtNdr+N8Q4KtD8
w/cEFyIt0K959+Bt9mI4Sj4QfMwiQ96EVJJMm08KtpDifb+mNhmATjgO+QEazyCZ
LxsH0xeYrcH8otCooE7D1iRkIoryvTyiIXxl33xpnfhSRwNKBk0DNBulD4Spq3d5
/lMoS5LjnseXd7+iaNBFceQM/S7x/PIa+BJL2nn+ZOHQbqe9MnC2zEnqTICOyN4o
f5nuaEARoAoLqCouvdoHGD1cK8FKgvCauIrwZI1ZIRMedi90XZgw3C3rojyge8bX
N80mA53oZfVq/C3ipY8CHUUKwg3qW1pMLMxdCQlFGwyIziQ7xiVTvULFNO5NwamP
7W/f3NxBkGJfZzPFTqGMSVcwqelHBjJt7wdnlmcb5zGU+B5L9SZGsBeTq2DDRaA+
9KBrTTOuCuwVrsU02Tj6XNgJH21TWz2XeuwjKetSoh7WAdKbp9C4uFOkfbB1XtmD
qb9NetR818NaRRvhR31Ip9u3OClZgT6s/FlRMLsy17nZVeoKlnBr2MFmS7qDWbEs
ku3BHUWHTcK+pDVJwhApsjkk6gwhRQj3wT0+YYpamhA9imYOEz9Q3kg1dElAcByY
f5E7NBDJURERlArazm5Wx87/1hrXZK36Sa32W1lprox68WMZQJmw4qqDpMWNYZX1
1bRfRUD5XE3e7A8w7n2r6ie20tGOQYO7Setu6hb8z3CcCcmvvnaCGIsY4mrugJE5
pR9KwUD3TatNmldt09utifVNX3djjVydiPH2eZE0hP3RlnOwYVsCaYRv68TQUohv
5jOJmLEiqPbhC4NPak/HYQsSHT8ty+M3kbxYGJmEc/FSTsAO78wrhTqzHJx8tD+1
ohCjpdbhwxW7qKUoWF1XbQt3GC4eNbQXixTFwhW7d12SKY31KehK55DYT5Th2MMB
FVPI2xIg4sCzjh0NebTlk2Pybhh5NK3dwoZUYrwyd60RSc75wy5drRqAtKElv1XH
krPvAZGNbVDFpgQSQL7gRsxCVIMTtSjNtcDvGyTQ+LAwGIFIyWzSJ9kLtt8a3Cfi
RcEUVgB6Mnd8Ib7At8L6Uf5nAaSdXluNqyynnndn6A70501woxqj5MteeDs25coI
cnS/eA4qsBALk+DedzM6ZOSau7mteGKi2dLtZd0s58FBAF8eITEWMDMQVvm/VQ/b
eSwFC089odp4Opa70JRsaNw6ig2NWPVQXY3hygqfmnHhbtiAq9rd+YPbdfbWj+03
cN5c8/RJrDFOZL6oNk2XmaihUNBgO6LHbPsawGgppYNexaI/iJ0OQxywbRo5Y2dv
Mtymx3rwBCyXJQJUIiJWmTN/x/CJndDIuO9uuLmP0vLuyUN+tePvJlKKjZMBVQwu
0Euj46LcmZI8IMWGzoAkmfMdKp2s7jBaP3tkda6VpTS5IoYQPF3ermX+4J6XG7bA
TrNhBDNcJtI+s+rYnOg1jiGP2XqZMMJna3J1pbvkxZ5WfLaC+mxBxN8bOCRrVtAE
q51EGHIEk1jfVNhlQAF9HXlDeZGzQfga4vtW3mdZ/c87kYmaTQdvKIM+W86NuiP8
3RT01prZa0yAfRDTXI+l+G/oHCNaFlPlNHmOadGPOEKyxzXsSlJkhE9t4LHIPrQH
7UbHtQ2znVFTsWWM7y3lzpyVC5Du5UitvnxaaxtUMDl5DdKzYy95vzjY7NinElik
9h3IgO/+hgrdHKvq4salJGpcV5EH49lH+GoqaA9aYmJNRs+80iAKboSGnRKFE8y0
e9CVev/rh9Fdv9VQ5hrNV4WM/fiP+Sa/ydflZb7ocGIXbiaB1CWYNoDg07YjyDCq
VYhDi7giUcG+giIfXJI2pxEbLTZO6kWAbYBwhiIJvDhOYqBqcr1gxwLOavo8UKzs
TCq9W1TWeqqrn8/zuoURvqCK5LEhGFYWFXyIvQZwdFSi590girMLmVMF82+XLamZ
RHj9TJJdLt+2ZPBVokWi8hQIFHsi5AD9l4VZj/25rvByLGmd8D8zXe6y0qC7Ypzh
eavlvljt2MTMz3zBu+l9n0OmhtP2zQ87wOFvUw3OKTY0iCKVIWgFNh5FZizPhhFi
XBG7G5HE3fs80+IuuwD+clwtWPqlfZqaO/01nTGnR8oVRaRRZSDrKMK+Z9W2c4Av
YkFGXkijzGE8WbnhXxvi6IGIpQiPFZghqZCS89UR13Sy1g50oKrg9sGkNOKkTrUs
eQeFqVuzfzoSKGYUb78ESQ==
`protect END_PROTECTED
