`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OoDV/BRcsgtDSM8NQMUkQAwI2IoFBghlJgAzjfy47D9Th19rONwI/nodj6IcEHkL
lsUvq5ZMmT100gVHSGxNcc1Z7/VGON0VM3UayxAF1Vp5au9dj3Qej51po8w4aHCb
f5ZaaBN9rCyMeJe8JA+y4qhpJ31Kr5+oh1AqleYVwDk2JVIrslpE8yl3V5Iz38Ad
khxAikya5f3Ag/3qq75xZkWpeZPt8f9FETB+1nlKaMmoehUEGXUc1O0Rr579VMms
23AHSiAcx0MREUgI7qemJJCC0CADayqnl2Jpv1Vrw3NDnCVfkwDJes+CNLCJ7sOm
T2641fjB5edHKVS49v3LskUK2mhFeDZHjwrvSaCMqGrg5HWpIv5ivyTS5AmU103G
yiIgeyRq+pxC++QdSnraTQ==
`protect END_PROTECTED
