`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ggx3mdfOGCHWJx8FooB1u1rSOiGGDH6AykllI6XGsBl34WOYlIpz+am7gSDyFI2w
xDOIqPAD8nIp72LqZ6Zef5kCIRuFmM71kqm3c1qbbPPShsC9II4Qwuz6eX7CMvRP
qxFVPOHL6+xjcv5v64oBRZyIjNaFZl5O96y39voCIgpssJ3lJYGpIQFYmztwdDnb
N8GYeBjyAA7hMLp8DdFfhHQ+m9yriEUvub4IjU7mJaBusuY6tW01CXZW4gvnGRw+
XCJh8WMFN6xOMEU/q7ksXHAy6ti7eXrC23UcvD3K+rRbq/k73kMJVvYrWTTOead/
3NHYkW1/emIGnAbyjFUfgA==
`protect END_PROTECTED
