`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3zuO6pv4oIOGzhB+d/SRF/PjyzuSN4k/wzWntjPjrmH8hKzP8cItHflqgEra5FQO
JlZf3HFlBcDhg5Gc4OA70P4qO823TMvInvsNLXnNWMqOhBERsvvmknuZ2pF1OFXI
UXCN7lKdDGu4vchiCsBwsQKP8P7Ojl+a7zD1MtO7jEf13sburF+jYR4pBIkKm1Yt
mp8swrFTKQ4pbIywFWgjJqrjsq2vmE3eno7R1hwdyMwIGAKbmHDkXY2sOFt+EvAU
lIVv1frLfFQeXE2YHY7PZycAUM//bMJtyJ7zRIyFRiNP8mcE3tYjIN+TyY3VbcJM
IR3UQeCrAU5ROfZWZ0bEv/Du/cYqhoa8lByqChCwfbbvr6XHrtcV//8qG9VC+UaH
KDNHicc6CPsv5n7gPdrNhw==
`protect END_PROTECTED
