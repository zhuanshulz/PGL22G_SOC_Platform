`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kzWF08iOUCEIc3yMDoKUOtDzORRGdsGC8Zqd2QJ1bvK9vpJC9i46DZBvwiqP7WZC
7S8vRaVVEQLRmJluxZ4TTVDxJbtEnhgo+jbY8RgWIBxazTuSWtHnSZM8ARQa+3c6
Xsv1MaZyxXJ9CGUjwTXeU4y4ZmEng0pniYAWt0hO/5fk7gIKFAQqRuTP41zfVAbG
fJ+5EFjjM1nocZCXRx1wFanKt+15yVECZYCYIG/CZzqVQ8LMUYYFpc08FhKScqlS
7FAkQfNa9FQDzwvDOxg7D7+fCSBkX68aUtj6DfFiI/KbZw/LfWmy9Q+zAl8R4bXv
LsnKWviJnCEl1UQAJxjCQxIOa4Tge4D75j3qLUjrQ7KtfPjo80Y0fhu9DKDOkVA/
xHMx3jWphWoEEftFtFxsVTB0QTyVxhh4DeuS5UAHZ3uDnn3b5LJqYYgOOrUIwS4W
Pxbwp1KxQwxpx5/oUhCy/wXoKErv1yTOVokprO3DR2iZ4x9L/501+1TArM6amcBP
GMqIL3dX2sE29LfvgSjWzYmqepSOY/B4sV4d9l+iY8ZVQZj8BR8NQDU5yaTpYpPx
Ql8V9MR7tLTHvZE+KNzhXcrVVOU0IDLmiEAmNp+NJqhWHB4b7ftcZUKrsknRPSnm
NVTqws77ZNuSvGtd4XUmkWXvmn65AojT2sQ/NZhUIWO7tUMJ+zT/90Y0npijrKHD
IjsyemUwN2pNFFOFgiu+ehgsof4ojEfC1lh8+aAra3znkt+OTyJlU5+C8KsPu8lZ
dHXn2EqpbYUn4f2vHc/qaYXwC7F9QM0KB2SqSSHJ0pZ3S4sibrAs7qCWSnnP+ar7
uYxYWyrZDIk+2LBVdDM3jsPTXVkcQNpzWbJwdUmWnIsbXH4BzLJvqAkxUGf9gvDw
cTUfWmafVjggCfy56zf0qnAspFFDrxYcFLWOci3r23AmT1ASxW0Gu0JApQF7Rk+z
Pqw3ZrLhTBG5uSmhu2wStj8xB1a/Tq9pxUrvQV5YL3JIcEC78hxHhdd0H1UkshKn
B4IE2V3Y5ojWUiUagT6qWud4lSxZ58FFbUkyqT8XZUbD82SpvWdPOpxktsa0Twen
mzYoVWxVP6/j+NfmRDIBok+qZ1YSR4Dofq1qku2o9wc4jqODZS0VOs3h63b9Ijt9
S9eQUZV4VCOIQOK+jFw3/Z/wQosvrS1VqRewQVvCe1fm+wxnR2vZNSGqpxx3VsmC
R6lE8P2uxGtDP04O51Kk2CPkuAdsCdOoUCNiS5L/krequO7QnNTqdqqiXu1lOh0P
YMjHDxVArNy0nYl24r6BW8jiVTE9OI9pE+7sn9fj1IZFD+600G9htgo8n9hxXkO/
TbFIyYooqdX74r7Xuimer8a7Tkz3dQXwwwgNUURgI3s=
`protect END_PROTECTED
