`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7vVaMmyB4ojFEUSWpAqbCsz2MxrN2U5xDWKMJEXVUKhMrl+CiZwIOCg5Zuaxhg1w
g51/uLIzkg0z2GuZgJ2+KjPOe39aM/Xp22xIFG6xi5vLyRXacxxDGSk2sE+PmByH
W3oG2lqWRVgCBNBkAJnhpT9ngoXvbxvBd8ZfQMqd6Gj2dxQCyszR1QOvq6uFAdDU
SMSg+qHJHUarGWG+neaScRK4iuLtwV1h+aFNBzUzPsl4HDaU662agrUTAgIN712m
H3DgT10SY0L4aWwHtDy3MXvv80RmJZPbHvgZ7tSqPhRi54NB4qRA0MVHTCmBriZe
9HwCoMbf7X/OEHFulg1TTLGzZF18OnT20Zai/L+mC9cpEuA76rGCM5iQJ8F8CpUG
37mpcnphSiQs8k1TIHhu/znJlplD+70ZqzaUYp+pFDDdPPcjpN8DffEuiJHWlDpt
42g5Nqk6bLoXJjaF+WgMlbfK1ZgFcsJHuGILQn2IEuGmj9mMRCdjtwYmIfDhERen
MlxXYHdd/li1fC7ozwEq0wskyj/DAR65m1dZIAEmcD4jYKff8mT/pnubFMZgceW+
JUwFbAmE4WQphwbPU0HJEyt1xSLbm/WElScS6aHKuLHgBvvfdyxQkuxDLbzXDYPz
GLaKrKe0Cqlg91bqdgK4zKcGILTjJ3pKDvitJlg+2yHpKtLZ1vCOw0nr6RJ7cfjs
WSAhGGJZDDd7YcHEMABH/2/0ULazu/tligSuRuSPgxGZtZQJNFQJaMoXEe2qsJqT
ByHaoMkcusp4mJ5O4taBoZcxKfG17WMQZ6mZewkw1ouUscyaA/MBchAOQGJVVr/s
5HqcizZAIYFnfcrhLX2qHv+mn1qUZnm8/gWuNWz7B3g4fYvwFu4FoDAzZgTpuVKc
+jF3dHscZZ9QnO7rwT46NRlAh4LwJoezkEUIHE/55z/iOjtF4OpTGtUUQ2Pgde+a
fb2odtpKWPX94Ag8s53ERHX3QmXyA9e/h6Vism/XohMAXjfyNKuBhaOhtddvEdY+
FMkn87TuUDIxAIHfSoBHxk2jcfmQbH6UNnYk7ooeHPqbbAhurr72tyybwhFBVWdj
Hxe+L5rRdw8KcRUeDSRQ6zyCj0OT8FwGGDdvqyzAjfU2HdFKryQR+tjTdrjOWNmr
h5hujshIld2HXirhe68A0Sc66+jM/JKlM+hvsWwzx7tQVKEtLU7dEo/JnLymuWwc
aKdhp/uzb6QwitQZy5j3AuAUGLnS/UnFOQi0+7u3fP0FzGldL8y8rkJpj0dwDgV9
8VWQL03Lk4qC+LM8XjKZIdcMBHIlSeLpZ7YuXEnd0AQots9HNMKga7P4kTR1fKAo
6UZjmKR5pAQk5k6Z5YXgzkR4M0A5ySfHcZq1yCMyMuVXa5NVkagfFlryUWVFad1X
Kfmp7rjRkEFFisB9bWRB8o4UIm1BGbJ1KfjLEqH1L6A6Yhzhsiy+UTEb+96gQwvs
ZBYKR4Gijgz+ow+pa31ZFWFy9FquKDCqqsTs34Vd+NzUQivWMC/ykDDdLfWUMpHM
fmFFLB9O0MVoPX4FXuig5dS8VWYiQvDmSS8RaepUD5OjUN9tilNFmDjBLOdSXvC+
fxNlEt55/wb8J0LzHzbXQab1mAMT7YRUG/T8JRpwwIENPrDFp5ypTBlc9ZBpd6JI
5ZaRbE13PTigiu58JeuMJ5SBAwI2ZE/FvQShDDG9b4Rski1yhZjP99zTKyy7Fmcj
mhAPk3neWQPXEs3GCFZT+SZbAH81+xcuW/outooE3Vk4Rpu/CnfJGSi/f4F8zynd
hvpEbyhkNsozcj5lgorDA/tO+izxc4hjimdTYPXKwsW/7DVCCTfDL9uwqN060xnZ
g5ycBbUebyPHIBfEB7FDfuCEllyHXHb3+LWSmJmoTTDFLvCGVcYDbJ0ySWJjDIa1
yDEvWVy4NCCjWaZtyjQ3X5cC69oTp1PWdng0+IMU5mb5SJXoqUXDaABwn5WOX3Bv
Jb2K2EuOJIVMTOsdGYGOvKxY/V3h35qs6rLuiR1F37EPZ/jMFhBm87AK+B9iaKBO
VL8WMG9yrFFVvHaorxFiTkD6jwN0HoT7t+LhxoQwTaZ15TazB3Dt3hY/2wy5m0rP
CWrcqvBe5eoClzkCg0rhPI+cZYBJQ05FdT0+/HY8xyJ6Xt5qH3tmBkmMmNL0H/LD
zMV3RbLAtlPuiFwRnuGZJ2zY8yemBHT5ebZNU5PBqjHM8D+0nj3SGNb57MUtcfSs
vt4j4+gOOgZLjh8RwH3nZ4cRLNHg0+D+utRfa5bmQ08wGxfLn/0OOKhI0mhqle+q
339m0s98pDyX1bcrAs3nTila+UK6EdPi+7ghOl2T89X/6I0JqRFSF0/1AYi5GEEe
7lGyPSlmj4xWxzjR3TyMIDUrc0z5+BWCkyiXgLT8wwa0mKH7FBYahWjllRlaz9/4
83Zt+IWZ/QRUN2poSeoR3wshr0g0qs/KoptIoXhzhcQpB+Y3SW54N9j8FhFdzERI
g6DyFojrbR3sabWXYsqlzILzivAU0qGnuZRCNwHM7zQWiWp5cdNeqjepOEvVsgt5
/HqPQ4sSnap79DXOt+u7gXJKk42+yZGEaeT6BpKf2VsMkRN1XbCzeRlByzlsfQih
TPlJcMPT1hViwN/h9P//EwiYpiEXucl3FQCf9lGA4FRzPuMl8rvmNPKALH+ZroZg
K9UUm8fu8epUyE3Dh4/ECBqAe/EWgVRSPywhA95LbVoNUTTTniXG5Fttz1gPugHw
VCmXPa6X2ylyTiSbaYgcAI4LpdyyPhkcvgFBpCAuLnHh7R6noWvg1NFYx+h7WLXs
rpVyuI7b81z4vatyKtP4XQf2/KEjEtz8dNXxeMWsSLJxPZTYoQdq6p+HeasL5PBj
eDuiu3oZmWLnSFB1dz9Pb5WzS5lYunBG7hVYDC9CAv9FFdhr6xyedY7phuGbBhyk
RC7fwJfEYBXI9xRrF9+lpENLYuOLBbZJNGVBUtczbU8HP2bMFib72QvASRs1SKdV
58ztMrWynm4Ee40UqtTbrKIOVkFeSUtVt69VZn8FnxiAKCOeAVyAbHgcNMozdocY
ZNc9AsV7CjZ8jhNyt5hEFazoTkSATnNG89VuhJxKxm+ZFWzESWLIzZmF/jKjY5Hr
JduDPjyK0saV0UBryvwJegL/4BlRsozCQ2NTdh7UjmVa4uWkipVhcX0O82xnEXVC
pp3b/Oj1TObLvuby8/Kf/RGJfW/jGK0iL02zqMv8W1XocX5GahjzXCHn4b7HwXeO
yPETHLiTL7puXptVOI85gT2tvqT77gTYRHgQyMcM2Yv5N1pEoMG0ifHYeVyZh5Om
zeiNLjNsdKklGCqHOGHB68wmzhQvijkvGgm6O5uV3UTWdb8HrtUtqH7Og1Qlnpy+
ZkiQfqXqxT3GnGnPhtpOpzqkgvc7SaA9NzzlFZpZmXuy/vTQamDZm0fEVyzMLfA6
UW589DaKX2OLngrCPHBLfJc3v6MvuQK0x+mD8IjSkxOokKuLG2XNNV9AfC/uGq3W
0jAU6DB+8i/K1RCdapg6lvdAvjdHYmGlKHlA8hX8CAuJzw6H/prosAW5oAY5ZeiA
9pxEvKcdO+QsZRgdVeRfgUy8vcwadaD8I4C+dr0n0JnlmaKkRfpRoWb7/Nq74ifl
bMcLeEEDKeeSu00WrrxPT2KlQ8hM7ianHgVgU/pyGCdoL4aSRRrILi76JKvJ2pAj
tCufvVULsCc2EwKx5mray+0XDZ67S007ivKXaVWFe8WnbiPMKmgxSyCKCrqIkVEn
v/EONwIupvjI/w5OqyOmJSojBIRJPvvvNpAy7oqkO0z9VsbvfXuFlL1R9L8tDUe6
XDXnV0Tdl3IQFZG10cLG5hjKENPDlQH0mocxInPQbgnJuYYCTthh3TPvvseH+J8j
ZEhCsRTOaUCaPNaNsH2LpIDRtEkXBxWHRhuOKXGoKFSKjc3dLbdGcsYrmNdqXpLG
vMKt0Cp+yk2N89udXmFy8zZ6BFsp8T3WD1RpdzB6OetZ5vADkO++b/VwwDIlEB65
j0tPp+M1OAasxp/N+OvKfsABaocAvQLz5LjrC1aXCOnijykHwraJz1H/Ph/q7S7l
OkQXHZ/aViBAxFtOwDoxv2ouvVaWQfvQY4lcvCoCd8jX0nNtgbptQhaFMUGMRPFX
141i2WjDLYN/S3Wr9qn9VflmnzsCc4sG8AkJ08bGw+v2YT/l/qJRk9tBUAkiLCGJ
T1MO83gHJALkWntk44/w8ger28+zvipd65dGKn9cHG6tbJZNCbXr3ZTDqxE0154U
afarkUd/eHEnPQLDf/agvRKmBcej6hzu6D0a6IQXo5PqA6broKecBfuPeIfz2ezH
zLDFlrche3J9YZStrlua+sax5JqnZq7gMzL3qcY/lH6yE6N21tSoVjWjFFal8vPp
T/CY2oPRIGY28V+BFPtLsQpYe+CM8pbRNyoErRahukKTU8Jj+PSmc/YEXNZoJIKY
Q4VZm4E8mu2pD4zGusAAxcaiRsEhTI3GKEmUf9mm0HGRq0nCf/U6IHm3GCS77eq0
mwJmt1r+QCrEgsLK820IqrVHF59dL1MqH1wWNiskXacClQdkAldADLwuYwIfpHNe
gwScQsj6L/6HlpBqY2ZkmNTOdvNGCbaKhzqx8MhWREYV2DY0pyR/jPDMZ+NXpSL4
yNxSGwlF7hCfIIKpmvduQOT8fZmS7vtD1t5p5vwT3WUmn27LkDrHXPZU/5pxp1Go
QcExsCoUjc2+ZW4+rCBl4nTiTh7fjIRUoFIK8iYDgWvIwoIRd/HJhZgsLsgDNW1O
ENA7Dq89YLuhVKvGHK9HVSkR44gNHmx86TuEOzzy893/nh3G8+1ARa5O9OoIGTOA
1yEOk4OjJIuh1ZQStoY+hnRIsoVJgQdEw5WjOwr6THAVhi7xtVMIAjW0K65lXj+7
EDe7EihFr5eLCxKqJHEoEGT7hbF9EGJWefm73HRdq78e/11T3asIdU0fxOZQcLV8
SNwUEaWee+tIBqOTxBLMIBSMIg9j1W+tjqUepLChUzTzVfMheBZPVrpEc33bETP4
fPA+beHJNLb/TU0UdVWnrNOmziARNaVnt9/adwittDjfCMFcw4r14JOPs2HdvZrU
WgozkV+V+IhPyMHuyLEPiui3105NtgyiMI7Ib0LcBiVYEMKsmkz/M+cLm1OwUBXG
d5RLsrba+dwRDeI+plJp10ovmk5I3yCT+TRsYS44d1v7gjmd70ufS6+lNXijQlCx
ghhuAKbMyoIPMNqzD2qfoS+lbfWIN7ZUHuGS46I+1/GzrIZ67+nJmdL7JTOg0+Uv
0cpf09yIMiVkRBDiQDgwjIS4CtHLojLvnayPcZP7YeuQ1/uoadIlOzbzHu6qh6RB
wk1EN+Wc5i8Z2yHbhvuNfmqcFmQTo9UP2spaqlAkyjB2q0ZspVFw46NqHHyaNURJ
HM646YfUD3LuR/Ep1LdcoDRvys9kVmSI1sKxHK+GEW7QhPaNSAohtgL15L9iHO4m
hbmqvEBL01dz/FckA/mkgF2OaDC0vaLS/TWiJi9whRg5f0K2PKVJbw6hNLbnVG4a
qvz7hf01j1ztsIj8+DCsWqQTZIGAYflK2Pid2veWJltUh3bA0Wh4hvYYftO5QO58
gZH3qbTCWjcasVZz9GyO6XuTFU295R7RvKO1axFBacnz6UdFSNm83cF4lTsjEBml
rkCEAWckPhwpxHW6OKivAQ7izcyXKDtbrWuqv8cs9gt+Ali67K84hH197PycE0/p
h85Zsgj4oiIb2K/mGH4yY97NVrlK+r3GrF7Oa4aZJ/5SWmc2bns31DHXlEZv4x9l
fJggAYZzjmMlzQC6maM7cEAxATWXrTRYRNZVicbIEOhVMdGvwUcHyQd67IFpLyEt
kEKZyof3XMGfaZ/j5BiDXLcHZJHPE4nlc7qFj15xfre3gDcMgK2+/jnRWjzF5VcZ
vs2RW7ZUvsKKTLWM3SGvtCm+lOhBSK8TuK4QuSeVMMy6fI/jFpe3R6+RhZEv/biE
oC/8Mr/BqegaUdqMU5FcQvN2Nj8ZRpoQ/Mm4wFMDXt/y3l5iM2BIjLtON/APLCjA
klM+wuKdhdOPlUU3nfMG42pgFwkWYxnLyFs2ccYHW7wgZCNOE0uHTZ1IepOuZDeb
YMTUkFfyZRHbuPUx6qahbTsiC8K49avnijcZqgTvCDjXtC3b7Fb6D7ZBt86jGnYl
oB+kHPkXInsuEG6ReZgGC/JVQAX8tVS/iHJjcKkEaMzPulEBYkpZVX87aFraTyCH
IBMfHKPqGw0j1VD9mQewT8GvpouF5oYZfrpfOxKTyLZRYGAO1cyPpRZ+//lLbMne
8bRj3tGY2DF7dGIxS15bjbcqUt40WYIAB0md2fzvPT2FjnYY+LAdXVpreMWSDL7q
WCrTXigplwbsvYlolPqb58Fs3V/4PSJFcAR5g2SSVnagiP1pvf+Tvp71v1z5rD9i
813U6HFUQhT2FIxuGqd/rAzrUYyNoWlwKvoDccbJdsyoUenZUguXxRo7U0p7TRHB
tC13FSw4BfuGvMhH1EYuxcKx0hQxREGpXIf2ApTb63b6rI73oi4qbaUEeH9sIIlH
SsO9ul51zaVIb1xmsLevsxlr7gcocqAXpJYxh0pL42zlTr9IL72Ra+a054Pg05IS
Wa/2sloSCRPbXluDxxWcrt84Sd2qrsgrdEpQIegrVP//dbJkGmPasSXnduPfs0bb
Y9niIgAQowibcF4eejFWlBaAWQcSVkv8SM65IRB6Dw+E7mgfw54sfdNBXi5pyVnG
IprwMSVtkW+KdbI3oUcDTfqZOGMJP8ECGghAAAFv+cgwCmfBn8iIRdqcjzSMyPas
EGQMUe3AG05HREHuakvZ5OAhRA+JOoq8vnoUDRIz08CGgoXZouYmkw0aoVN2eaCC
qZ0v8RhZ+tCJWJDEsdh7JsgJqrSIT5+vPsYbWVWHSdjOkG2Wlv507Pzux04GJTlW
Ed9FDB0rMlocjavL55OzK9HVl3m66tHHwcjT5ZIW2hzwl80FQPVOrpq5gykHgBOz
SSYFsbW3cuW6RPWSMQTIQ7HeBS6eEwi4fkDkBIgJhQple8B5xx3pC7SFI5tWpLx1
PLX7ihPy9z0nWrrSrJecZoMpfoOrlR4UdsrM6JdXCndTvr4ys4iBoVtX6Of9E9LB
nltnEw8T66R6vXerTlhmK5SGCA/Iumkk9kVks5ZHHlF1caeNjcW5syoQwaxzxRSF
EwRZRHkNyhCITfQoKvXmx++aDSWf1Fbdz1vgiQSVNx7EMUVcm/vcyZyg6nUlWrwc
ZSk+dPX6DHVVHnH+EYLHQccOPUgAkadjzEAm/anGt3qQ15+GepmElRbjDIVKzV6+
9PyxdfsREffSco40ZEHCSOHY8DNdAI0AdFsp/D2AYnlCGc8g1PYLWliGtOVpVw+d
C3+MEnwpPeLErLaxAvgPEnS6X098MosPK/Cb353Oe5uV2MigBr7Z9joU/W9SNdiI
pdGMerFuzkX9jVgYbQM9kL27QgjvroVU1vOaur4h1hUqnRU+qsevfEtxvA5Ql3it
08lAwCu8FNpPyAu9yjkJqh1hj4RcXOq/QC3qmFr3exOIEhPnB/92u7/frqH1kjmI
rNwg2FiLyxLYyHChuQ/D4YZbm611kDS5RvVjLqFaoe1rHkiECbXiH3AGL29SDTUD
vWN1UuXiK8avaeniNM6I8n/PXXkvUjOks5CRqS2m82UaZtyMMc8v28ECufSND/Dk
RbCI/uXIYG/38M3YEmvzL+55u98C/kN03MR5NuhTx1oPX82NWEl5a+7eJMStRAX5
ellxIAS+YhYp6ViAwFyZxbTJkIb7MjgBpzrGOs4kcJ2scCJqP8wg0i4sEOto1TnG
d5ZImroly/1i13ypABPYZAKfnY5qYHgd9ng78zx4H6nXGSk02OxI4Wpv8Xe5v9G1
u2aOtwAjylqHnopNWKfvchzpOx5Aj7H0IBoGiVMaN/K+PoGhB0MvHiy1m/wbpN8M
z+DlYAKmhWjuFFe8ZlqKa8US9fPx3SF+msw0oF0uGG6jEZHT/3apTYJ/o14aGKt0
9gboL51Hs78xjvKtR9H1yl1ceMO2eDGINaSXHUQm4/tXS+RJo/jvjgSdg8b4Znoy
k4yL+xKwEjYE1TJQHVs5Z9k5OT1AUQlUhu63iweYj/QEiNt1yheoolV7/KN/VeA5
9icaQgfaVrr/MiQqziNrvjE6ZsauNUXad+1kjDt0AXuJFajY8lzp7WDxL+PaTpdS
C/N5BkNXLRGHVMDKXBGzy4Hnevnk5KePlEALZPawqc9ETo9O4Ho7S430qvpGuvI6
cXToWN2Zwozv/yE3S5sYd1bh0ba6fIkHXOyK0FgI6bxQ4ZNIA8mfI/URjU5NuGRZ
6GBejFYK3d2efqK6lmiz7t4cP5kImBNFoP7ZE5CK5bCRo+Xr/FG+FnUP9sGJfddW
u0zo9G3F1zG0TbjRnpLLdYrl34TpiEk81Kpl5ld9icyvsLBPCNybg11y4WBznCHs
UbtrXAaqu+Mqx2dDIWyG2ujn2BQIFI+oLfpgAzOxj32tB8uGBwdIVY3LprQmhKQt
2UgjHCF0XE9iVpNq5D1OVM+O4Bq9WOV1nfio23R+fQta/9Dy1U3naCQqtMA6U5sp
0TLH/OotMYBUheQRKe4RrAlIOnpyx3//j80Tnrx26Kmq+zOmTSJf8GPcyPrxyWKn
bIDTswwX/oXqwsjToPU/Y4ZPbs2aBQ2GyWA77ITayJUYE+5lQGFVRIhSVv2nJBzu
45g1dOmn2eHeX5IjIrshyeh5AE4B5g9ZZD+l9gHhF5J9+1wF3OLHY1H4+VzEe62+
plV11yF/9MyEhU6gKGpqmIMY8pjLMOIcuHMqusBkDZOtorglOVYPUspPFfUuJhRH
9EPyIV+Jymmzkwotua2aIudaKFdtDZ/35JXWURmTwebrAdk1VsRqS4wKynCSZ/BC
pBLScYIyQJvB27EPhz9TZZOk3N/TUacYsubhyWmnl7dzn04pUc7hv/ZuX6bbdj0t
6uav4iB0zSs9fWnHVX/iiYBY6V2KxaTwlZRncfHGP0x3cC8Lk8szuzCDXslDc9I2
TAv49K41q+SvcKPi2UFoGCMndt1JRi5qOAO6XNrM08Q1r5D6fd/xePbwC0PtdPEf
Q8kbS5GWI+W0aMs9FjR66pXzNX3ToXmR2I/um4GwbfBpYNlwPXbtoraRvrExFflU
gDwa7K/Ee6AZBGs39rlBrQfGbpXKb+ZZeoKncEviRcG91U2CppYERTdzG3yvtTAE
uoamVUWXnZniREimxramyNA9SlOOyaQf8z0LRg+q5t5gQKo5+SxyxD1hSYqttjno
1XCzJI9FOxxYAYt/Gz7jJN3fj+JkXUt6+Z/kF6VNKXbYF5N+jgtZbHEqRNvKco5C
ggjbSzQ43qqBye2Hszmelyn/q3EjtXQ9+Xx8LDaZ8wyGCB8x0V/ewlBmESRYCEvP
bo87NcTwT3y0pj3/tJsRBT+MIMlaa9XhRbDJq+qZ2PKh9ok+2fpYNcnVL2dMSpVy
VIuc0XNdciakK1S7vFfpcF00Qre9mxyIEfCW/9ECPvoMptMVhDYchEjBBRs47VPF
4gpBG9SfGcBmixAeC2xav8kvdNG4wSYo7qycWYeLj7yqOcuEoX/LAg1i9HhFP5Iz
profUw6fF8V8r8GKsE1XDOMrdtm0W9fO50Ow8Fvp3JsD2xEaTVKuBRRJIDqRM7OR
Zo4tTYS5+soCIERCytHzcBb7U56fFoSNppJyf9LgEyf7VtneBN0D+MKi53Buov4U
yxeJycG00wq4tbxYs6tHjpQT84BoH1nmI57cEOy/XxK+v4oHToFcsNsID5gj4Wf2
Xvwq45uU0HqkznucD42B2WsbLRPpASvOAswMgerTe9haFUMPV0kzsWCbdyauNLUy
puOagTOLvmQ2EG9+pYStdIKMmYk8SmJR1koMnFzq1G9Ssan5pi/fK2sA+1gqfXRJ
rLMJJIX9ZBfV7VzoBnBEWVtFl/dfvorDLjbI4kLGgPnWKkQF+yuv8YZ0+y11SIKe
zLSiqJ+XGAeJ4bQzeGG31D0gAuF6xdcMEW6n6MGtJu4uBMDtDuRsuFj79TbdBdNp
kLxhlqXF1CHdufEokMXccgz1TmQ1fzft9yUVJHNzKiQ0GkGNPHa3ehkIzmEZoEbs
6VFOpWULy41XQWw6doRR6ntjHlad5FZEfEPPLwygRSefhIythv1CseXDkeqsA1yC
G5nqUDY7sLeOPaNyq4hHw6Qdf7hStFyegTSKcPw/j2C+XP4RdzO0d784hu/lRQk0
yyEoZ5moVKSXjom8v3ucNSCCxmLywHWlwNgl5wFZG2Fhu1w9yVvx9pp/HeiMitGA
ovE2Vx0qUe8B63+2VsZOUZ2aTbEfZnATL3IVwF3jXw6AAvdHXYSU9pKIe80VJAmB
MLO7sm7UeP2C1lr490aPl8xkKT4Ant/bdkZlYAbEMhxYCDbrhpHnexRXJp5o/jeM
qaq3xxISvaZIo0zFdH/hZbsTK64jEWq1xCtRDr2Cmghi7E/GS8KcpPm9cllLWqgN
xWIyx0MzQFdK6lFOUYRbmLpB9tKVD6FGIVHIjeTvrvlOcB/oBB+gNuZH3YwUv8n2
tJI4T2UfuPOAE/cP22zd0MUKGEL5m4muEwTsxjUgAwEeATReGHZysk/7FTzt2Kmf
dajdqRxthGZch5xZVr4B/4xQUNEQ2ecE3xs6IsVPiUGj4YrSXVgJF5M+gnp6sVAk
RxHND01mvkZqoQqsZjMlOYy8XHyyOVWHa9y3/2Q0gci3xXXmijIWx/i3GheYEZi+
0EdipVpBpFv2N+FmrjLbL6P/bbszRLdzXZzCaVOXmAU2FbNzODUZpYPRSfQiueQH
Z4oEcmJF19SEVm6x/4V+tgWh0w02kvAgq7o6PHzwUhkBklQKSsZj4SqVB46Nk38C
LQYkrTQJR9IItYRhHs8Rqtm/J7NCp12n7FTEAz9EFTkiGuKcdksZWHmblQkvJfXj
DJa+SU20dqqBZA9oFEDJv1OrlAT6QR5CxuglBZVkfMPDqV10cDFUY2K0dRwOoGpY
j4AAg6LWTlDPF5COsYXpCff/8RmwyS/+x765s7GxQ29nJSAEsCVap9Ehj1qdo2Qy
Xhn68ibx4R3R8DTiI7jEbnF2HH1rZTuIotmRk2o/VKxttV7mLiWYUjB4IJM88Bsj
M97nGHujo2WzFD0sPO5Dqdz/4AH4IDPRZ7FYEf3sdBN+zzJat1YQ7ZYXVohxtTvK
pi9E46cZztU64SlW/cblwpWlMn7h2PvpEKV9hVfft+mEjCDbS1wN5jeCUK9NhYGo
N25ghA4qxoz7mSsHfBUtZXoKRZ/RGvzEoH2Kb3hGT4vXb7zsPApZLEvNf7fsyjtP
NvLiBKh6gmj+DlxCuIBgk3tV3u+/zWK84hP8bIx/F9RTMjTaQ4q8IWAUZij0jlda
m7oJT7lQmNnoYHtd8tuHwBvAm0vnSO/UwjnEH2MpiWUsio6+6lOFHA7HnCv1UZrO
+BLG4jhD/TfZ9m5uG79Wq9VsmYbwzX+7TDkk6P9R2voojZc1YFAsN/Und1KO4GDN
IXyDHi3QuO8b76R2jflYkIGG/sR0NReJn5XSJyyo6/0X7iBBTLer/zGwomMJ2qd9
UhkhplWtD30CKvgufmAQNYP2D7B8H68WnX/2UQ+5UOt0+0zH12ZUCUhE3LeTswJb
L2uIh53TmLXTigh9fSEugIVXlGO0EeIfn/giL6CY2u4rtayWhgqqgZDzaxTvoMIP
jpdHG+opPBOned3G/Ql5YT4TY7JmDB0qvOCJpRmBuvtZ9tH4ZPIDA1D+ub3ovy4d
ksmQq/pC9xgazpdqAawHL96N2RSZ5YuqboHp0VArvTPOZG7q+Oinl4SzX5uhj1JY
eYOTHvVspaJDKsCAAK14Rijuylvr0YtkwnuYBnLR27rVDoo+Jn3E0TsNdJjm9/xi
WBSpfg4bZ+ukFl7I/O7vjab88PXccQtbSGewJo1nhkOgHKgrpmm26TbzmnWTqvPc
VVfdGs/PTRw0Ns9c0SQZjIqOyT6TAqzQ6P2IUKh13nhKY5ucpc6djEXZ+1MLc/IX
0IwUZVeGcwScKINeJtm44X3Y9QBy6EopeMKBt1nSLCS58SRVW0yhV0gAhNUEmNPJ
513xqax3mcAyYHv41+b9GEk5g/qFSPEl2hOIb8i6bxPCltaU21w763vHsaSpg9xA
daSfSNkFzDSdWH0+znVzezNJHVl2DUrBeqRjhWCEDyL+DUKKBTlvmqzLA9gArAYP
MzTi2URdTh/KTATTKWE9N6qFjRh/Pe3GBGAkAfSkq5JPHFGhr3O3ldAtEq8KKeVV
VrldmWj9WybV8JHaXBWrf+RPnI0nB6SMDVXWku1wDJXOrPLKO7ZQRCTER1AZU9n+
ampFAOd2EpNLXMGilgyAe8YITSwBBxjS1uINNcv5UjRUPnYX82QzZsLWUdN0R/zE
fwtEpFncfsmJ59evgerldc7FD9x09iHWHp6roDf3kTvF+TXEGQOMiF/5DTNAWwvy
OTTmdPL8bVtQeTmK5syxx6g56HZjNRXetEaWgeolYIY19a3s+w2VRJfai3ZP5QG9
us+SwUO8D/eCTJJlPUYGKQBKVeSrs0YLXJVT73W/jWDndH4qWmR0NLlOq46l26ds
JMBvBU7yzMlTkxnQRJMIjt3Mv+0JIv8zDdgjbd9GgO0A8zxwQjC63+SIoTNXUEs0
TVRf/Y65/Ofufw1q22lVKJowLIJE0nvZFOpGLjrtryH9vj3R8ed1wCv6zlJgLTis
fLNOLDZRXUp1yJy6uHZqXNAovU8DlE+TtuVpXfJP4HSYTn724QtqBJZQe8hqtfmb
AAtMLHN30MyMJ2YUFN6yt4IOO4iVp3kMMQLd513M0HT/VofN9vNz+u9x102JO4zN
bCgmeAOsnMGzWxYh1+hJpgIgYAmHuflXlU0XJj4TO0W2Zdx3As4pQ7hxh7cQIuHo
FluxRfD1CPocuIPzhvoCl/RkLc2BdWaGcbgcJa5w0Uiffj6QyfDw5iOa+z/KjbVx
VtTl++ZnKCeWwuJXuosLM0U6lgxUx986+wZ2lHkva2zqqpmlL6n600TbyrWjuu40
tSmKCZnZ41rgBaXwoUyiP7Rb+0AJfTGcrWBN1eg4LbraIFH2X47XHh8RMbVCO21X
ymNTL5dgXMgrgu4iM7JSCGWoRzg2sTZ0lptgHUpad4GQTwisFpbUegpHCziVkwpG
uhKTvVYAdCfpoy5C86SVPG/hI4V2eOs/66pCZl/EhY2rKuQS8Q6Ni1HzGLnwGltL
T3VFddG89Dpi9RKyEY1i8r/fxvwmyhkeEnwm1dNOhNhP4HHc5P8No+U2PjDYCxct
RWIeDSJrTtX9GXHTt9IBh1z7eqtORhOE5iRYIdjfzmAgUAGroJhQYCeq4spMfbyh
dzcVWaOZVZfltWJGqmKPqkxrXI3Iv/lOanoSlAIvD4d7B4ozTRCm+rNXAJUiQYZX
81ABW9dnyJYwBg1WI16uJET8YyUCDhSGyJcsC9okpDCu9FJrjQpN3l8HlMD+AdPk
NgTWwU3Zvyr0aPyglyQ4gBDciowNuirZs1L0cLNdMSfZjdwO3hfEEe9RbU7B9pOp
GK7udRP8MfKnYIdbnA/cyf4LsY+DE2P5bE96iaSpQXp8QD0ycE44Ep3RmlIla5hS
M2xvFtaryF0WTbci5pg5OCOzfy0PjhWCn+vYKn8GwgErMVtsKuscqB96Y/w7QL53
1cgcgmerOm9bMnGRZ3DU8WnP2GPd7xWF3jjPE5dkFzhjBsXDVqsquABgRvHdXU6y
fwDOfNRMsXsXjPZGh4MMC3iAwSOUFBKLJJlLNGSsU8aft7kSqACzpWUjLvIFc81l
TNZBbg+HQJ9UEZ5Ny8SWVxvnbNtY4Cwx+bCAdRVzemgW+pzXLH6iiL2y69hBRX6l
C5eDXkg+A/N+oOT794poiSU6h+WTA8UD8n4mUC9G0CJdl+tcXPg6FIIZ/i0sz7yg
fTsNWwLxxSmdB9BikWSK+sJ/uvS9SWVVI3g7dHswtS2IV47ldj4OzZyXNBeE41vc
Ek8PQqopdDS+x5Zf/u/1GxvI00XGKgJdzCqB7+SOd8i0nBtQ43ydWor0z15HR+Db
Iy4e3vLr9jCei48/HhDXKNxvH/LF7JpynK4nWQTQgJnhXsqdz8gYBEk1S/dJGNMP
iIpYA5L+MZMAeB2SWmkgx1ZGeMAMgxbHIE8w4D+HJ0jitmhFohsc8iqeBR6fHeOy
Hrq5AsKwogzTExZMorVC8xtpTxSdOcD+38+sQkbf4+yrMow55T86F4wR6TOhqnxr
F/SP0XTN7A8/tzf2V/UQuifXQvlKIAvRD/7915sZBcz7LJ4Z/HFiQ0WT+6WRfFQl
WSCbhr6WnkjvtuASYFBa21FXnXrRS62RXNCgvaruoszfc4D9rDNGTNYcRFXxHwRY
X9KhDIPpHUoi4RlyTKJbpKXkWi8BA0l8WKlCP5tlZjrSD3pvbUOuV8SKbCXCHSED
hb8WZ5T7LpEKEuohGKjPuCUXmAxz7qpExeL3wsSEgWukXn18h8ZpDKAjF+/Ai9WA
lMSpoF855NU+BJlYE42hcskbOum+dQwdr5cL/ZbFKqsTx0krvqiMsQmqoLLUXrl2
3GgyByGQhGomcVX8yqUhkW3cIg+lfxrQBi7L5Lo367eqf8YzEf79VXnAUyYztL0s
z2Y2dZQ3i7JtxHEgUQ5bJ1DFKiu5mECKcO7GvIIxCSqo4CsPFiB6oR4dIIiAo/7d
NP2q9YJ3Tr/Fgp4HmFhtnIU/AELopzZNv3FPEtQPRre2p7R30osYjF+uKruW3ixX
d4ZWge4aDjcKFGsRlxewzeY8DcgS7rFRGCvFncaYIhrNuYILAlOoSOioWrtk0xC2
TMOYSbWe8fQPB08xy047ulW3jLBiQt5w5DTb7mYusuej1qfwrCcPixhfcv8FjviR
j9WFXUdnQVbaHi8zAsN2JYGzQi/ln/J+tPwPloS0nfBq3WedepK0DSYb8wnzXOdc
eHXYA+9iejVKhlf0JvDP+SKeiuhqdaVJngi6Td6isgbSQkqMa4HkwCjr2Hv8iELq
yfISw3dlnikoF9FrbyLqU5pTVXm3xMHuO5qR5Gd/UQ7TQEdPkvrpe8OfO3XgQHS8
Yq6JpVNjaJI7ScDRtWV9wyAW5LLypV2IEr7/G3PmXm4RY+Pthk9hvtxvJqnpaitr
Pv1FRLyViCoNuqDo0rXKbHbLc0SNeSzxp7pIDgOdcx4+h8wCpbC7mpuUZCVVfDWA
HTs2xHAECSAq5WP9Ea2n4iS5/fHG36CxDjCZ+2YzN3kEsHjZ9I2zD/63iySUZv2P
aoRyr2Q60bsTPTSwOzjlohBURVL2a4shRdNeko+5lHn4GPBsfYAW61qJr/4HcTO1
UJk9fEMnTyUtQYgluATO3mPNBVkzy7u1f4vV4O8aCKt7RTDFIVmR/pscAAkbh2Xc
JO6SSHM6bRQ8SpFaa5dwKXDhtsxUMkajFJ55w2gbNAYjWAl4Qa5aiOS6hlJGDWSG
bk9WAn4aUF+EhlaVDisRt+QBEwgWCf3xpcdHZMNojvfHFprp235IA78jZ56GPmIV
hfTQtIhLALRWd+Cuc6xYqcHQ5XYCzmxivCjq27HAVFWSnurRvUyK5hRf6GrCUo/O
LSw5j7GYzoqP/O7aJWITLYIJYaB+KgPExW7aNstw24Gl7cJf865s0MwuCXp9h0sF
qp6aLw9l8PgjFGpM23226cKSd1EMfAR/2AhJrSxm4GeMvYAAv9UBtEd3lAS1UguO
AIaHOHJObSUtlWqkCtY8U7IKaUI+OxCneK/TQZ4Bj2iTkkffCAzDKAN+kqDbXXTH
QtddStnOoHogntsDX3Fh3wjmevaLg9S/VD3ckTb9TZ1CC0qgUUzYjL2d1xMBpf4g
rRNvXltqfTyomGXpaEXmDp2+Kc/ndcVO+UpQfMtAzEc86TvL0uUfgPlWKlIrOQhP
5WSIcn/JF29U9DDtbZK7j9NwLgy/lHQ9kZXFVhisxXoKLGP/+lVJEhvziz3QH00C
PmAKvbg7ANxLcESQ9E8F4OgeYFuQcVWrIYN1MO9QKqywRnTdSNfCnBpViSkGjJ4J
iyHsjbo+kTNxW/HgZHhJIFSHIRtMSDAWKxFd88KRwzF5pOX7CsKdfn73EdRMaehC
/P6aR9gprdIDmfQz3RCq2KOCi6JQLw1RaiD2ho/laGfLxCFY/li/yZrwuu84zxKh
EYGtG+qiYd1vBN2zCoEzVkoxd9WOnFOeJj3OxeC4/ttAD2r1v/mxxtYljWVulF0A
yjVIkllhazcZIJ9oXwfs/Oo66Hzvu2H2Hndk75NyLGqNRtzFi6nzyGqGL1w/cHfp
v+eHspwuhj3V7LRse3Onkq/i1/GmjCOkeHjkHSwpblqcUnosNF7MmK72vnOpCbRp
9EY9wniS8vHdsS7jSNPqCLLwvYt4PgvHa3kr67ZUgfjHrs98uQa/Ku2sOLH4XEkq
va1cAARsP9ELyFiYc4BJKGkJjUB5FbyfSalTYYCnwaGDXOH2STqa672VHY0tkfx6
KpJDQaTgeIxIELdPgVc3Ksjh0VgJj6A9McuR1FUu4AkvA8S1HdVtzAVvwmaisEH2
UVpkbAI6ArANM1HN/km37Msp+CsThGR3MH2IuWCUf1oeEwvXuetn2KC4kqIX6o8h
bdxt+oqq5F5FoyMUY1Q6sC3plK1HjSYPSBb1kxVGDlzxS8Y89jbXvCywd6MggyKz
EXCU9YBPgmBeKwsNN8lt0Q8q6MKT8w6lbiD3P/Zgif/oe3XZg73uxA/asZ98WnvE
7LJD8M+Ok3JJaCvoyVwRWUkJTKGfsGwdeYNwUTWyWu35ym0132fSLP+sJxnJRgjC
kx8XAKAxU5iONih71f5f/U25O9j5CoT+Zs+oRPN6Ywnz2RkdPq+2wYWke5oD+8vg
UFj2ugeiBtna/14COsWRJ0SWVnUbD2C8JvSkuz+erV0OoJDFKZr1vq+o3+cOFWeP
WuPbybQkRyfCEkk/c1obME6GhKmCGwiPaQkEuxZvqmsGCNoUuiHZOHmDkSkSpPQw
E3VCaBMWbfoXH5Ie2LvisRgJVHp5imrslMpRaUBww/wu7Rnmcf4Y0mzDWkbk/rHW
KPB41/+KGiIjmqobi+wfQdzPwJ4Jb8O0QgBJ2a7dRR7wXqAYvqVGnzg/iv63d692
UwWKeki+muI1LVB6sy1pakhoiyKClCv+bxXoDJHVn7LrhDn9MtMPtzOOd/sfQJVO
fZXQ1TyJQzLsBz+dKQglRvCeIC9mWaSOcUTeIwYEV5yPWPEu+AMk6UdHVwai7+39
uPUQVo6gs1T1mjmwk6miUv3P76tLe2ldPucAO5l6Op6noEx8AMZKIIOztrtbT8qy
oAwtk6PnN0MHLwo2A0Ynd3H3EgoyojBIgto924jVhah4YqP1JNGtz/1PGZLzNZVQ
kmCJ+bGY2PqtJRRDMjPjLqRRD2jK0B/0V58p/aTw0Y4d9Bv4J8UV4NMQq9fX06HM
mJtK1DTMrgVV2OCGqAbN57x+x2PAmEEIkJ5plIakB6ZaoLBJq9CtsnpW9SZL+hWJ
CSMC4kiG/fUNZHAJhK9WvUnLIyUw6eoguZBO8Q9ocjPWO98d9UTrGe5OmLxVKlsu
jIq9cXPtwqZFw2rbeadG1ln3Mbr36IuzU/Nbg+4ni4LEERKeVrZpwyVfQA2wSgS7
63XTgMmVv8MX0TcTFMtIOLo6u9gZ3hGBz7QXCOr1q4hRKBsDQ7O2plezklN4nhqn
A/ZZOKjT6SXVS7UVypELiY5ypRYWTYon0gST/hykcygJnJX9OaNgUHmjYZZOT84n
M6JtXMh+A7GnwKfB58eF19pqvp1xaBWB6JccgKKTBAsYr1Gl5Wg1RGAFXemR7kaz
uYbkW1DknLtIDjYNLlR1CcU+1HehUXinsFbBoK7H1jmDW/4DdtbwExnTzA3y4ba3
KQH53wQwCKncw0aVL/JIC5k1Gbaj/uX8qHA9tWXj0eaIX2HL7NzN660HW8KM23yV
PYraEjqRIUI5UUA85U55/x1FzIN4mQzvrglPL1jY5DMkY6Bz6ux8NQ4qeUmUcWQ7
4crt3i4hJ926uMLuOJXaPPKP94ujvAru3r3tSwO4xIzxjeI0YSXKbiUHpOt9hJPA
g6iNGLQwguB9hN1gCZ7Z+ub9idzzEwUKaTbWVFA8x+qWod1jrOlP7yAEpULOZ1eb
kMEShxcbSiXT0OMsOfEz1gRIGM41dSaqNTA8ELwzWzoC+ci3bKCWyT6kclyXV7cu
qMGRKd/wsn1P9eGXK8cJ0+CZ1ehLxxpmxw/V8WqPUNr8hk8mqxL8Ph1cILqTMXQK
uWBP9bJLgbhcHUtfSd8WM4n/xrTS+2EbmjGioMtoD6MbStSQORAVdtayhHZKXEh9
JJB1q4AvINWkveK4vCS3+Xtl7jt6iSj6ClnZTU24qZaRmBclpqCebZjJB3NkMcmC
bqhmEabVs0dO7/NNJZt8cLGtz6CXpYLP5rfsQOi0SZruedgQzJy/xcXozjxcGo0E
TAtfjB1HrGPrrQ/sDSMb5HPXLrEIJQKrxBpqQD731L0Ba/X+1FBZhvww5XXkhNYj
amV5ZfeOSjfUlXglojDPJ+70SSONuLno/y25+7wZTx880urLcJvVjVrUMneM1V0a
wFoLbkIUzNTkW1lJRH1E42ClmZ1qP4eSKqrzGYnmjE5KetZixBtscf3B5Wc/aNQD
T+STtPzbiP1jv2hE+T252CKE9ZwTJVw9cQdgUawBsCwEvbVgvSzhRQypsaa05DuR
F9j3dTRYKIhOE7KVwppAF7mdZb9UPrfC2KRHXDWILO1QEcWD5IW9MBoiQb5/W3vV
mlktgQFTgLyyEhxvQRVUR9gWWFumBB4lsqvBpQVgRa1dq2QEwt375AbckKTQnVnP
OUhxTeb09jw8/T7LJwXQEZIt8ijG3awtK2xoZlFN7uXh+PyG3XXgGn1/ZA4gJM8Z
1xjRJ5hDhGz8KSFzF+dFTY1eBlPd6t09Le5l8sKFMPb02yYxPhYh0fMWlVDEuYkT
3nI4HEjw2Q1iazqIUPxfbRuKG4YY7O53RhIMeUwIZ68PFrsXEQ7zjcBcnYocTzCV
1lGlpYlB97BKdFkYW17Cu3xfR6oJmAJLc7zh79BGLIgt9UarqnalG0BoBfv+ay/J
YZcmt2lgN1xixFMwAAlG8mVN4l+ajCn7fiTAmFofmyXMY4t8iOcHbE1tqkkYmcAS
D72a3Z0xnA6jivbwGEfCVN3+NNrTAJpAqkwf6XiNZjGqZ452s3ipBiW/lP6rtZuX
Js+nCO/YLnDGw2Aq56HSH8PaaQ/Z2dxNM5Q9Nw9qVW0YXXWHyfKmmJydgQiFy8oL
ZFyqDtNogPm3y5GDOgfn5ZSYT2ILOksj73xjaij+DRHdhTTNoYVU/3pE0IjtMHmW
XdknNGcuaKBTDpmdW/J4qx7WzfX44VW5pXiImLiCBBQn0NM69bT2Emm4N/jGuOkZ
2Wek8y40htDQrNWtw8X4JkaNkHPFWa/fZZ/Ikkc/xvGJBtbBJwxjQslAdvyye9iA
yYm+HcNtEzHmou40cjMQB3w2yQgqWfut3RE3w9sByMwp4EsX2SrCvLMjhKZCHviZ
/uqrkhSC/at1I+bDV3ss19Zu6upHKanBBpfNIs9ZJOzUgMkVcO0VC5nNOELtBy2+
0i902RTuRC3ugDmtGvK4h2gQJ5PSKhqY6hy6iYPEy3wo5KZLR5a2fh4vvwfI5jqg
7L+2esvwCXUNrqfUzsL37/AoaipAtmuug77aDrSbjq1yEb87TgQwq9rBTFGQNjho
QAlzvkm4yFrAmezlQJ/5qA+qWdp/1V3fuiYAY7e59afrlXfjSi0Vg8P0A+ml0nid
Gd/zyPeTSix0uazaDiTX98BNIwc3RRnG3eXRPA7JIGNXKjnqKHHhoISP0AwGwGo6
7TzhoiDubl9m43ZOoPouC7GTZeljzG0128tmeQZjc5xcphgr/LT7MoaDQOcq7UDI
HL1ZBxkgOCjvs8cXjYbXIzwLl+37tfbldfSI5br+bSn8Ab9LmkB0lH9YJiurr4et
F8lFkUaqU+X5lTCl0sd0jJzYruUYPOOGaqsyxBkU7UWIdAzVPN3yGxo+a7puLHoH
3GChv1RmkWYqVDVSNe+iWKKhzOBW3ZqW0zsvQfyyIkxsYlZdyceN191szbkPO0c4
p4nG4Y3wUb7EjT+IVdUGxyZSyf03n9GxthsrkcXDckbhL90w6CFY0J/omGI0n78h
GoQBkKDIGHqlRJTu5JpyoT2S60voA24V/edHnAmSGDp07n27Dh/OoGnuunZeZHED
JD6sQeHC5yjAySgpel/C1aYxKgiOY88KWV9WKB/ioN994advmaWZdlVOkK2S8+a6
04vzBp5ibPJr9jeUGQBJuSijLzSPQsmyUWdYkijLJ1soxLeQhNnTcz8dQomzO7QJ
e4twRLeH0MpTs76xnx9DJWPfm/dSb+gGogPI4YNp5F3CNRr5CENgqmdnD+guEIV0
UfURn7tQSKOrxpEJP+IQlK0f8QVm3QlHZiAnUD0nqAxmNCpbEd1Ok/os4jjU/lWL
+w1yPmcGD5Kx+U9/yPrnPn1TEne6njdrr+OyWPGb6xrRCfExO7oqYcZv2XpN4wpY
ukdeA0inXHjYW1v1Eu7lxBW2rU74gjnLbUTqdg+H2PcfytvD+1xK5a0upaaddF82
Kg1vF3K+IFKScJkmJhzMZbQ8h018YHyP+fc3AC4Bug+su7BSnGaKBCTWOSVBKr2+
CAlVMR2ml0Jg9EcMoGUFbknrwhJrKhm/5IlgUgdjtPEEWCyliqvxSuuhFk7esF58
V253fJ4fbbOabuxM299hpRavLmEutWnLC48KwIQL16S7EhEtVlqcmQuMBnjpmbC3
bA+OrrPxtnTuHbG6pVzpHbo2VRTAs7eykY68C9wxm88NCXzh3O8/4CkgTAfsBuYb
XWN64ht8oFylg2robbE5tFC2O1aNiz1vDgJJxO9iqbpdTMn1NxISm1spU1PCoNa7
6i2DQvijJPvwduFuQ1JLnaubOcduYv7yUBfYBs8tpj6a/MFF3/yQT0xSt7EZa6IL
OG/dDjzWoavA8UPZpbjKefP3NNCECyj2KJCfKYv8EwAXU1B+/o1fmQdlNXn4/N3W
28riEEbEPYFlwmKJ50rmcvDaz6TYJKz8eyKVq8VqxuuGDu2YJdcBizRZQs9XiwSG
1CQDeLXZR/YfIy3IWr3SlCMkeQauX2l3QPDhspEaV9Mcikbx76Z9tEEeFz36JViB
QaSstxCMYUZyc+pgylJr1cT7EOVj76TXcAq9ioKGNbqeCssajfbHdNxNXgAoew6I
hK76gyRugJxwexRH1O6XeFCs70jQHZEyAsGD/xwgerHFGo/BrWyKg5Pc+VmvSjsh
zBPvHycBdepLw/r4Ambvun5bF5Jk4XaZT97Hka05ByKWkGuxAy2vV1HSYvtPsRpi
zGIT0NqT0LVVsRiO9Gwe/Ea49r9zqE3OIgSOsI79iozIf29ro0clBrzXCc519Vhb
mPxotLdU2Yn9vx0IU9Vq9WoeVcpGvPd7EuVe4bR1RmbK/6sjjFgRoN16gqEC5nRM
WU0y3P3TZ4i3I6jfwq04P2abCDhD+dZnDpPsAi3Q0cLrcFAlZRQFe0FJtsXUGAO9
gDJW3ORcZJeklILyF/2l7j/sGDILAw7/F3KXwOGHd0Cn40mCGuHB2xT5SEI1agBE
UMdVaGIm1AJKrkxrCt60FXpDwTMIcvYpIoZgDWwekARka5iQ89dADbMf+jopr5MA
Jmchb/kwiLRjHV39gRZjVy8SAJz6aj2csczTqY0xQJUp7pOSh7E1dyqisVNnf0QF
Fx4KBaD5OP2+SuBpQ6R0T+vFQpzK0Q7fgUFituiuke88cBtTa+T86Q5tRy/fRWCC
dGc2P24FLN2iSr3D6RcgSSkLRFIUAbULFTdBN4w3Hc8L8RcbRLwJurxNIx9+Xo41
nY3lnxXS3SokOJ17lZVaBZ3bqIiJ6tWlcSn2NGildgFKIrWJF1f5UCGjyxgpljoa
F62TDuRBtKKmGAYcWL0JULGu9y6W/e1egTPlxzWf5FeieBxLWGkwwuo+NsHDE2JC
juK93aX+ebckGiSgM5/Hd1WQbzBQ3ocvGvivzscngxdQ8igtCHzDTdo68K8Vrwsv
y5z7ZyPLIG/GUX6b4V7SjdEQ6z7lhTQcQc6dE8TQf8by3+b+o7BNqRTAXFWeglU7
kNzTXa+LNrYsCJIn204w2Q9fHTrCANJ5Tbdm+wIm4S7XnCVPgWcaxx/gO1hbP8D/
rjLeqhSLlm3PKe0KOpRI5vDFc6Jr1MugZNjJOyc5yjj3U7BlHfa7DwPmd3HVogHb
emxb4dZwae88u1yh6Q2mB3E4eG2IBAh9rnk4Ha2LM+WR93vleNIq39f1Q23rsQIm
Wp+Gld3x8JJWu3F24ZWPhSkF/cvCC7wM4ewjHKLD0XUeFuNythIOIQcGH61drH6o
yS5adOuybgBL9ZccTy3S5N6LdNjaP5jxw9RZSH+0t999yCXyVYUYJFA2ewFYlOWi
LHimg5KBB8nhL6XNGYgiHYFX9QCU7nb21RXykR7ZTOz3Y+ZTLfHbEQHOFJMuaiap
86pG40an7FR82EKNLeWO39OjpSkemjJuZMPMvwEKjmOD2y4W88bTaRiOScvrXqSi
aHb6PdCEmeScOuOB+8ratyeYfvkCjfOINxp/8nlf72ZXgAUagHHAd69Kz0lkM7+/
PM5Ph0le26gFIuKdCK4y05zsyHE8ZjO/87gOIyaXyM7Pnu8FZASizo51j9ijIcbN
bQR03CtqPOcBghP4O0KMYnzaSNwB9BCTyCWOUgVvGEU2hHu2gzmas0EZyLbUtU10
9BeEMuQ1f824Hv/1bZ3SJ5yOsn0rgd3vbv2MDicNT5iV4iwH2q7JQ6tnT8Sx5e20
tEbpw+YG9LVDWzVMIghgI65FbjGNbjbsem89OshTe7+Mt9Mz5JlNXfZE2dLlOo8r
zggd40UanHOHT5t0znxifMeT1DiaE8fBUoYMUFnNHj4aeYQ7KwNhX9idaSpBXn87
zdir6FCYgiYt/0i1L5CIufS4tGPareNfuiPIX07tTi7esaX7q3zB0I4VbcCkw5sB
B5CoeRztKthdcBdqZCEEu8YbC9sZjxLoZNLGY6n2UdJNsPeJk/536SXzZOK31bdg
fi4eCGm3p/Tmc0ZEmMWPXbof7Ix/ZH9LbjpvPz8CDcJRkvcf5v1NFeQ/vhw+SEAE
IJ6XgSbppry1tYqVFOO5SAxV0Hm5rJgOfCjmxnJhEpIUTh+92p6ozZenSc+UJQPV
TGiL7LC0TllA/um9R9kqrYHZXk7zXlRtdBAFMM8fBr3Z/xqbLEFPyCDxcp8+Gvl6
vQL6TvpWBYUiKF+2AkI7wqtS63LGFa18jD5SI5+x7jjtZi7UC/IyX7KhaEp6lgjk
HmKCNSPREnSmqrXf6jGbzP+j8XcMXvjPRbGexl4KNsnVINTKpsuUnY2zJ2gG1NuU
gqF1BW83I2Wo9mPiRBuvu7Gwk4D2m9WBejX/qmc/rhZqiEoFI5Dx+JcHBVXvO0i9
H8qev7yg83HfOYcL7rrAgj1kZZwSKy+Tf19cPYdrEDcwKpyzqRC3m/ZW7oz98Elk
ct/rD8VOqZQWOAEg+4qwBCo0Yd5+CN6HdAm06cjm6suLuszsMen4EAzKcMtXqvQv
UU+m/KzenaV1A4glQrjcXGFExZr+6j5g7nS9q9SqrUkTlEipjxiSdvuQEtvbYAYW
SiOUEEfJq+oqDYjbDrVzolhNKWeKgryS5xt3rNKxqJxL6nFhF58S/olGZ7nTz7VU
hkmIwpg8xDW2cFBxzzRZQ4kbLd9hmqLS2VW+GTNHSWTMMRCQybTIifoKiVBTLYGW
oGbekYylP7Mn50tLJOLlPtOxjJSgPKPRctHyb4T0erYhfV2RtU95yhOOh4JWscMi
ne22zfSsNpU1LUB+TDjyTMw4RWgriasLi89om2ktGgzAuOkxtCBQp1JMvLT+Ulm9
Qt3+eQJTLfix2U0Jlfyw4P6gR5NQfwXUMick7jCW4fItah2eZuHfkTwX8/RyEhQG
fMsnrWaZb5jS7IYLooamxJcZNKYlGoJ5SVwOzbEjr3/IYp8XuIw2HwDQNPPvhbJC
bZmSI0PauN/pkDpzLS1j6ivcZC/+YJZuCmDC+rQ2KqssBT8FxA5OI39C4HfG3NMA
weFtuQYKbAOfZKr/3c90j3TVBHfCW8zC5V/plvgDzcOVeeXmM7JxRCSirrPkDNhk
Ro8w8W/Idv0f1TySKicqsb3cQxzgeQSS5wqARWQ3cUrsWCVhiQpZZsdLBJQRk/qf
TK/SRIo5wJQhK+WVrAv8Awg0tR/QwdZhUEkuQWjqwNroyqI6oPazguRGO4EHRNbQ
7cqlBO1HgvQ7a7KA9PSRZl7KU6BZKsSeMdCEtqBxizFvXd8c/n9imQafdWC3LrRh
7cCBmnuWhXLISCmcgqKsmx1HlLmgtQa+yLgb708PIY1xH1Hjr2QGixqhvVPK5y4b
4zdaD/O6/ps03aQmEbwtoqwuCBfkXEhIQbxN4IQGFVHXsyHymGeUp2RPMfhyaGFX
kQwyrv9pVF5mRKWv6CUEP4PfGkaSAN4x6GAO3PF/LT3auhW8FMAyw/x/Y04ntGj1
OoJOZSd2/DC3E62eKnu97hHdcQflsAZWE4N8bWmogdTozbtODFirRqcrQHz3r2ZN
1DmdZeJAm3Qjh0e7U3niZ+cVFrFU1cZ9gWl76eqN8CLGiZyjuIn5WjPpYF9JT5Hl
P6lTAswVVi6wXWcOIG7KfGsjJKzSUwB596v+GjloVUnchCCJ7E+gDspSV7VKADnh
oYd714qYFXeczO1igP0XrMAj4yn44NJGBa4wKu0Fy/VDFHGtHjziUPU+benKlar2
RFiIWLmj9mXTauOsys0uAs4xB9dIV2CNGpsicsIQ7ea9d313yi9vHY78or5AHY0i
DP364G6GyNbnNkWOySLNfQXmKIt8p3VNAp5JZHKCLXJuRNRPH1yQaVMcA+2qB0QD
EdkqYYLL7MIkStFrqbw8rgttbkdhF/vZZ8XXfLNkZhUJ9BP9nrxe3FYfM4tdC3Vu
dXLlEVRI2xAHxDzbMtYIGgjXECo8JHNqKaCkwojN9Um+cCC8fl8O42LZOly4DH7y
F/DR6+SAMw1iixHBSXjtiOmTIRwTUI29Dgl+qfU8BCVaAObiBB7bEzhEJESry7PJ
LRU/Bsg/7vhZlvxNa1e2sOdDZWio1PbO+Zn77td2dZ/AtFbgPDC613UKZgKExTHd
+GSt5oJeooq5ZMbo+chnOT3L9VVsAACXmX3g8zt/OXUjbCApKi/QgNUc2Dq7XGTR
XKWLz9YPHJZ9KOgVbkpmAL3YczYdN4glqc5wkutbR41kWcpnrEp2twzKRheUE2wV
ZfbO9vPS8XsCLKzNNCcQryKYDAe+7NBZ0qDyKGWMgEQW7/MyKkgKvQZtLosCIXEe
UG5+gMyPRhg+oSkqc4zTF4jK3I9vMoiqwqJ4gZG+ZCfv9xhSK3y8rxo6Z+kvAYhy
sdtD0q22kF5rlxHbUK0HS0SVmMk8rrdCaOMG5pSDM+bZwDH8kQ6pFej4rMa+Zp2A
GWnaZOLa0F1oGAqQEkcewbvDEqwqLwer/8PSRi7ttn5NRErgJSwSp5ZuqiB8gIfp
9DuYzRtd4zgB+2/Bx8PQ2IKkVGwGaWpT2dqE1fYK2IhaqNTBltQ6fGGXgDa+k13m
wwYxJiUJFVLQFErAaX5H3qf3xRmIeC2Beg7/QlRNsUt8ZBHinKGgzpz+b+fYe3my
jdYSfcAPF/BNppLa7os8xl4AiI2nn+IsUNfXsd9vRGjr7/mVV0bX8/OhdMd3sa7d
Y5mOfpsez0L/U7Jl8qZw0Nllt8ABlzXMblHm4g+Py/i9NgIB3hc1CGO1K6rj3qT3
f8w7TvPavRj7nHUEeIC/HXKcuUtMgss7Jy78uzKbrveQvsQryDPew2uScgRe3V1f
kW9v7eMRvsEtzbsmaZZMOZ812/r28w2jbw/0wIUEltNAFOZ037AxoCj2cvBgf0aA
v+lA9RPFHcqKRlcOi1OBb5l/y88BTX9EoEMrL+xa5qO0nPw7cL2ttmFtHceMDnxu
FUYY/lScQFRtVQvsbC6rQrF8b6fypBv0g5JEMXc03nFQi+6KAJUyMg2joLTdDP0S
TD5VvqKS0fppxIsVOE936oWhZ9vzhSIbVND55zFH8lFqFkb0FUdZVpEbK1y+fttX
6u7pCzk/bXtVvNWzsTybl4QNFQ2ZIs/NJZUe/kMmVIhiW8zW+WfKQS3jn65caE3J
ihYhWL2Wy15FwUaO2KdOsFFHkQwIf2oDcVrMcpo1dxPcPWwRWGT1BAU5UT6XoVPt
08RMmNix9EWjYrv7JNcw8Y0a1C+rGg79sZTOTiiJlNGIOxWIt0E8vRs76bR3GKYx
qJxJU5iyda4/5eJt2+UbWStzeH6nr2Cw7/gGD4kaIFXh2j9YqfGrmwsx0ScDX/vh
EDjQna+TeghuMg/gR9iwv+ky8/sTH8tnFQRH3Jr2PWtqBv/6scli2r7/s+tgJs/R
jB+vlUYlTZK3soQNv5Uq+pbFT86/8javGyE4XNb95TDKdyCJjSwpavetmiAspEMu
BjtAbcPWtgxO6KOIiaX8hhpebMkL+rGXZqy4+9lWLDyteCaXN3VlmtqVCYVSGf7H
zb0+BIYO2l9oRWCspD4+tR6QWkQ2vKUu0F4dR4+l2S9zi8+B+4z4JSU0at1xXM80
Pnz2tYE7u4OtjerOPztl3rzI1Te4sYGpqlpzaxGxHeaGl1jdVimBR6MPZNy/fQ3T
rKaVLuCWjQ8L4xXt+6ICTYvk3Ld7cujjbuMWdID+AZTntw7Oxn5haw5MGc0daj8R
8t6lVT2/yjLLJZCHVVIRF9gZI5xwABds0Gvo0y+7vn9yEzHHV26kFBKTYDdJVdkJ
itFueMvIsn+AYUnKqqHW0NJb3vW/854nznCLFGPO422pn1KjcG9d4ihaQyXaZ6BO
i4RZqQnMxsVcEvpMk7teb0AJq8vTP/UIMm8U8IoXmR7TjAhZH8D5VBzLzaK9pIzX
u6QCUnSIDzPqAHQ4fb9gF9Cs2IybmJKoDBE1f6Bg4hVOWGht39KrQx73qjPMokT6
XsTcDNFUkmA5wCwUvsM7rmZ6S7iwYFdpGFDb/iIQR62ui8ZmBw7zx9PNCwfwKyh0
AaKl4f209PCnqedWr5C3oRO0C8G8rYmRca063xxknP3xqPhI0tjxGi4Y9tdnzKLy
wSbeY4rOUChLTvlqpwl8lmlewbJhCE/JInRAra2MOaj2Xdch30ddMHJgEgYvDVCM
UHYC8HIFw4filAGNejcBsALJtPUEXJIbsF/o3bNqRC3ft/3nEOsjWSsbm/fBjmRQ
0jilfuRE1fxKGfsAGQA0GIYIo5g2ZrMrpQRCpuzYWJWIOPlE1+9F4Pgjq5l692ja
uWbQBe0jjuiijMLZks0v5IzPMggHk876Un7k6tRj1Zf2Iv5ZmPvp6EUo3oE+wxNr
XZ3mdGNv/Kf5Cwxgp/bCgkMiZcCRukxRexDL1OjaTli0YxP2HbLtD/LY3d06BGRX
u79S/Ewm+YVsRIEjL6l4gj0933cdVghqNR4uF+SChDPX4tR35WogH60JyqXokDbD
QCviTNdu4ucAi5Zy+T7YrvZyBCgZNzZwEKX50bK8cG/PVYlUtnzDEysvWwsOBuKP
PyaSqmTWpvpUbsbxj/NKtrl8I25FwKvvERoBJ/ubIFQz/RmtNtVGP4PrscSy3zXN
Y7cjdLj3Zh65mHdjz8r7lEo0Gj2+hnrjNLWhFoN898Uqelhx2XTQKTfG6+OJy586
wKODSMZtB2f341B+mAlmrrbQCjZf4qNsD5N26TlszOvfZrEqe4C8/tJ+PgJLmN5c
L5UDVh7IF5WFiCILCIOTGboIo7OAwrqNcvhgd3cU0zZuSm8lw6ZxwWwENijTEjpQ
ByDB1x6BxvNU+oqWnHMITH/Cvv3JH3QeZ8Tr9X4j6zdBIz4xY35sCaR6P1RWY1+G
IRMx7tgvwXPvPnqbSuTY6DDCWNLEEwItaILWMOJH+0kfepnv1gsHwKeaM3U0V+P5
PFfsexxWeL4jgv2HOBKQ8KNeSj45Ej+b/IKCIWjppOX0eGIb/TS0zVrrniOtA2ld
APYqbI0FtTZeXKVcZRMCjbUeniAT+v6jEHvN10FJw4E+WhQuyYIKGIlGQI0WAH/W
LVa6lgK3R+mcFLo4dr9aKLfpSChuHd1Gyzc3ngzt0Lrr3UdNE5Y+dU6+kDBXi82y
70GEjCZzmLQEYxtBmTuWadXgPoZWRM+8sLdOa8QS5dZSSTsNLpeLfEDoO1JTTbQM
I37/d5t4HZ5+RvK56k7N6l+cyQS9L1EvcnZSzcT0uRHs/vJBupld1DARqGyoA08H
D64zgMUCr8L6AMPXZM8WDLjKuJmV7vdhUoVcnPQzf0JGXDxG5JmHGtd0mCuYq2TH
jE4TNx6Gj6wxDxd5Ie7/ZzzYMu+OkY0GP6nr2UmteM8ldwbYDhm4IuLvh5gbrDGh
UEsDzB6cMEkOd3WtIxVcRBf0NbzeR2mPfEM5ZNgOCFWB9zrYl0YetxSQ5whTYNT1
XdkZM7ZdP0UlAPKUe3alP7eVdlEci8s8fdGKUHBJTRvxmMJ1Gc50QNHQSDBkS9an
ufEy8Ukf9EoMigW7HCJJ0rIsiL7ItJ3oDLM2aSjZGl0bKQ1Am59nOtGjx2deoqt2
D8VCx48Q0wQ6YM2Rp6nIRo946gAAZR3IRlL8CkcZ+f7lPrgfHl7jC48/tPG43/nh
7KMJQ77JmzVV3TJKrI3nIr+egyTitiW5Tpj6Rkt7/5breCnFpfWcrWs/zH+QEDj6
mUJw2hRC74fGnzXxURiR2dsg423RqBYTZYdrxvAuO2ocElm+EzbpI8INd9tjuMWb
Q53+UYxFvgfDK/gvh84qNYX0wBl+zrBcbDaQXy/ubTXbuW6tDikJfHXHPqh86EhA
4FqLpiXY/gH9qvcgtohegpfZmea7HbcAu3SEJMUqAqQMijuD4r/Up/yA4cc6FsBC
Wmlz1C2tuoc5M52EMmrTcdVXvLOiFFYx+Nj5O5Kz7rTv+98tr/8rJ2K2QGm6KC3L
QoIcpXn84pPBhEQu4W2At0/pWUaJcAcqUa/fPLs+hVKhDtQx4gzFyEE3RxTQ0FFX
6IXlcPSn0yvIZWVDtpauFjVUVGqEzCmaWeIcPcVGeRmB+CDDXD0Kkw3tmXyz9owE
l/K0ZSNuQE61kwnAFJOE3TGTZdvDr8zcV/ftK7L9ycdh7sru3dEEJYPVoLo0qVn6
xNuVCAFp+c4OqpHVbLMM3VyQshIWziSvHDAetduqewA3xXuzqdvG5yoahBiwgarR
vk30v7VmCAt/pqMdgSyge59Qj2oY5cSrKP00I7N5au63wQYL50nU+PmIJ7V4/kuk
doX7gV8yICBXmww6vrfFPMDi2TIbK6SP54k08+9218pNQQpA9N4/J11gmOYrAI97
26aLd2eSyfjAIeZcAk8gS3hOCoQ+MhEqRDk1N9j0ugcgC1sVUFeLV+9OWHj3mBHQ
ErRXr0mYbPAEPLmmWqXGEEoI485j1KCvVToZdOmhuzxA66rfyhe0F1H5OpDGBFhx
/BeMZZY1IcQ6ccsAgKBEhJgvYmB2BRORItwEiGKT/7k3iSLc8ujlAX1V5DQEn1Sk
Yor6lCcbd/bhfXC1PHHnrU9FFbt22/x4dU/imrlhYiFRIFOWd04gscb8OsLH43mp
mDQNiGlk6m3HUtTo5es5wecVugjoKzDmsV8epV4joQfa/5t60utII226EjqIjbzP
2iN5W61QQorIkB0CfPlG7fB28gXkj/YDXS+AcJmHWh4q8KSRbEtjyLUHUjej3Whz
iYoXrRBItysmB0u3SEip02aDYwbj61qrnZQVpQ8G0Nhf92yf4Ni/WLbm1p/wHTvk
AYRz3JjlG/M+3aRRUHQJHfzVXab9mPyTwSBfHfMK2sEcglVWfPP7aUrH6olmzNn+
bu10Z5lCip6FHmSH1L4D43LH0Ypam7AO9r9x7PLDZqE1hX6yDGnbrdwl3JQ7D+MO
NpKbSgEN7SX+qIhRPmZfDHO43pWaOevMHfca79c7kLsgjIhOP5wGQwcLwX+ugPBy
pzVFlBIL9QHYUfqInRdR9M/VMiOiTwpRwezg7QxS1/JIfHF5TlChJq9ZP+FfwTOt
2OOA8OmnB8geLGH1FtIh9nephLMhiWCZE5E++OLZX443RJ7vNiuazequn/sazdum
HpYaxkObjkCtzX+HkD81/E3Uupdi9qmXXvZ4u7i42ZLC4aJpXgJiT87uTYF153z3
8dswo2LAPuPF9oh11SMT2zWIf8KMcv8wVRDSfNW+ezrnZHeSc1bgr4+AD0bLUpJL
tGZVHSNDqocrXXk9+ZI7NC/AEumWxMf/O6+vuCajS82bCE0KK2pQJNgrktX6m9Rj
rgirIv5AdSvbhiPeATFs/6QRaucQl4aTgJjojtTqXabUHFgggUMy6kyyOk3HW7dw
J/XM5I8tZNtfH3VFG0qWAaSzHn30XJ+Yz1M/0zpGMAhdB2dm9Sj4NdhmXFy74ki/
u6XJooBMhcnA3Q9Hzl3mB0NRQy8o43hLLJy20jHlbiUzx5VPGRgIXnx6QpYJj51x
PYLzUWc1X0OLhzs2aVFQoDXpcoqU24eg3hCOstdaRfmzYQArl72Sk9M2sz3ei0k9
yEps7OxKQBMJ0LCDpkGyMsXrR5xpnSthC+4YXYfR0wpsdFUFsxvqj3bwKrkiuK4D
0Ms/tX+6zUbDQxdR0SOVwYFY7ok6BWUXsIID83nxThdaTYL4RmVY+5rxR0+I89Dz
3JNHGwOmnfR/o9rf6WTaHmnGinJkoBMQGhQ3NTQYyet9eJjih1GeUZl1tIj7+294
CHQohHYDFhuMyQ+YXNlfjObxuK2HkI1YgxOCQvcMUPjTa9l/zJOEZ14RbghQW8kc
5bjCKYnK+1PvRO1IymLmrdWSjjScs48f3TBrPOPlOun39ZjhwY/8O7+VUIS8rBRL
dm3f+Kygq4cTTCpRF6UrwcE73XgBTLyWZD8O5R/LPvyKQzb4DUw3eIVoCheFF2sH
03RHe9CIcfxmfQ0oX04AQcz24gbX/AA7KTW5qvPfxOiw50MuCZIRmR0Akr9Sai3b
sEFbEJbmzPxt/M2X6tqToBdDHc9vqZcZyT3K8z8BLAMn/CfSKtBKEsNuzymLm7rA
h/9TJ9z47P2RNu4vfKkjjor2mKNl2GxbU1EKkcY5IBBKGsdXC04ZogLTqM/2OBVK
iUtqLEnMWpviOetQLlnf1WwOSttJQlAg+j7QCA/GvpctnOfEaz5LkdPgF72+oZnE
SGtDyGCH28tZky2JS824d6ABkQuCLC6h5C3bAfnzBx5XZr+cEbFcnmXQ7uGGio8I
PfCLWd11SDBYyXc+S/OZ9jXSXJuGJxab/V+fLUjhSzvDyV09P273lJAtDrlpQrA4
D0x8tHHzfQStHGopaIZpbYpXq0/pmmzwuaWYUVXer1hT5it6irIP4B5q0DvBNPlc
7B9dUkk77LCRdLFJ5cq00R0Ak2iY3mLpfbQi2kBvE4RBaRQpHB62xJSyt88ZhD40
7Y38AIwGMf2KvvF0DBfubtK35+6/NJ78tfBbIgVoIXQR7R0JzVC5mikWiBcXEFJV
LwJCGOxkhEPFhrqOnlDvbwquqNj2fLl6kubozBEMsRdgvwQ1NVE1fxxKCQ1YBsji
fpMAjA5Dmnvv2g7oj2CXfpiTvxy7pE7TLUmO9lR2rxFqR5aN0B6jE2RhYa93gbBD
difvNYeeu0cZyQEsYTUaGkUmOIFFez7wp04XblYKqtnK1p2iNeSPWGf+gZ31gItp
UCn4SGnQm7DJ9V/psMYFyPo/tUZJbHWQnYHzq8m3Y3Iqb+7JGRbiHhJ7dhU5Ih8K
rrs8p6wQfvKP0OLu4k/eceB40+47JSAj54USjh2jTmrsIfANHolhO0MzKI9GtwGv
xyMPogb994B/J6h8Z/DbotnFVOrn6gnyrOYMH8xAtTJgMelM+Cg9fKRTphMKQe9B
9UrMUns/qWA5t/0KEc2PtiVexkpNGfgvCVYiNbLmzeuF6qa6IJvxgSM3EtqxMF3t
pYPtbe63JvggiNvQi54jFmIKbX829kaXsZfT7lUBAftt5vBevLiJZwS5tPCU4oGb
96/MDgfMk6DqtW7npuDHbXE5HoD9hO0XqTL7TRF2wyoD2ph0LJnoHb2uD587WoAg
PULZgCTM7FY7jYCpTOlPt/4L/6sXSxuFKEgGQk+kQuzzwLacnnKJvuz1Xg+9DUJ9
3heEz+ayf/GWU+2FOTbWEvN+Alr8Ny8M7mo2QER2inys0lFvzowEZF8YdXXoOUYX
Nh4IX8GdVNdxx7RAbiOuYlx5p9+1Qk2Qo+pmx6Vq6fvhPSATVQvp3rFITJkOECjz
7OT0pcKuIK5cFmGgkVRtdW2H2eeoHb9RKhzZELAGmZ4N6k0l0SM1w2wHxAXw5hCt
5gzg6B/w/DkbCYN4XUKjy1Fx/cYlnw8NBq214A8vN1B2SclkfSEhVpNOKM6/k46D
zvTeUv5e4XO7c/579mtqIXD9FYz1c3WLKVui54/qfNpYEEF6cwHTkU3clJYp+Mcd
5in/PlGOXTuH4hacvPpOtFMs/0GXT0dV9JAUkzombiJ44plJabnh71LvKUgqqAeS
48joALQZrEeiPTHmDuQbbjgHFJZb+I/uKTRSvD6XD0JJbKEaQFS7NRnHKMLO+tzd
W2W1B/V8cp7HXbTSAZ6VKs9dBrF4+dcrkIo1kdaVUwZ2TCqydf0neyBzRYqpeUpW
hSs/hrM0w14kf768aZqJUqXCcynLrs4poIGfFIX4yHs/RghxbYXAi3YlYDi6/We0
0fL5ANxOY+yERRT4YSl/LFbqszquJs4CW54vfRVcR2ONK40eQlON5NLlHzPg3v7s
3CuV1aoUoHjACZsoOhKrPNpbXX+VgIfNaKLpGI7gMI2Pg83eJ5j0Q+fNW1nQ9ruC
5CEUpIRQVjacxjBky8coPGQWTbxIAO+iVcLPs5uUKhwZ8sPGHuR/TPoqmh0zSbX3
qCs0San2V1rKKy5z/3Z1veVruy6yEb40K3yYRbb7rhobNL85lCRWfKolb2MoTgwz
5sTHOcJirVXf4vGLytBf0f16fW/CFIvTP6QkrolGLKi4zytTK+sCkskuWWVhvc+2
uHIGL5bLGCWIMGzRWt+npICNCAVUSTzsknavuRcQHedpBWwxXYvh7qQvv9cfFkp+
5o2UX17y0M+JuLNCSTigzfrKM4Boh6Iq4qEljga2wwNaH78AnQfTTuqY0klR/VmB
0JnHBMb7x4iKBdsh6uRp5Vavg0J4OQW/0z7zCKjRP8/lHawH6/Ekwu2Et3Kl2K3Z
cpo/ENqxEhx768anxgss65kwFgMawEXS+67M9PbcRh31B6agbLJ9DbbO1fhxl4gr
AWHLhhAbczysJVr8izLbcl4dBtNkJyxZT334yrxygZYiQ+6DYyAb67QFLxjc/9Sx
kZ1iMN8blFh/hW2BnVYv6AXgqS7J4nYu490DbP/AJxHWaWBxgtxBqaoWgKcgiKkW
cYZNTlv/w3eaA42wfdAx5K6emhmTvQhnjwOT70tjPGsOQYQ7SYvoyIm/9ABrLL9+
c0u4hgB8RCWvF22mMdxzpiQYh+C3R9gibx1t2iN5CEsP4iPfVG+CTXK9LfnrJW/S
xbKR0cvgLZ3QydtdVGoM7gcIGAoPY1RsHgLn6mI03eXKjHk//x93N9VzgGuxL3+a
MoiA1tYqwZqplsR9ckSctJTgk89/6WH+q6N187cEq7WV/IdcMlv0z83zj1F1wwm1
7N0VYHiMvYnB7djtnHdQVdBsh3tZ8OpIvNcnRHcNzj012WgiiRxUnLaJ6MwAj5x6
3UlSC77QH6r+gTiRyZVlQIMe7vGNU0Ab9r12DTVzhYhZlyg0Oxfb94e4GHqjKCfS
JnoLd5xIQt010iE+rNhXqHVThPlGjIAgg3vWlUlQ7OWS8N0MSl+uTqwMIKcTT9Gv
3ERkCaV3vXezMfU6Vd0iNpWKWpMh28g6daVYV5OChRSHP7yTBYl+SDJLkDMq2Xrd
Kb4yyL9VUy+g1hw2mF1/mO7stklWvnuMRk4JVF1xOfgsTEMfXjYSQv15JCjiCwmx
z0yXDWb7tn3RRNIWCRk61MTKVQg10PgML5lkKY2MkOMyC3CXvWRuEhuVLVryiAOj
zQIaJF4CMPblWz2IXGWR+vlsr9pGqlsakroBNogeDvDugXfdmoL29KxQTuuf0U0E
PZjZfa5zmsZM4/MiIQSk853f9dhcmCBM0PSEQ8KtDrbVo25BYMt+bvTi8Izr30c1
8jlt5bnC/g2zmJYAqj6YSAdAkzoefPYMjK4D0K95c5C18cBjBwvnuUy9S5laJby+
T+zgf2fQFW6llDUzkKztQ0+utbADncjBjTN/pMxCGQWpH555FdyZ6++c5/Hqycvs
4MTb2xqe2CKAbrZmlHl2883JX9D6a1jE1iP2oWEOQipuPYt2qnq8Fw68mjOWScc1
`protect END_PROTECTED
