`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Nh/6RYsvJU6cxSuj8O0C+D6QbXIV4aBpdZQmRpaua2zx4/H1TGqrSnhzRQZ9Q5oZ
rVifSkxEEHtXQOPTBlHZmimzcPmcbPEQAPIz77VD/QOKUDE58p4S+hhWoy4iEWKi
6pgOTF5DGMS+dZRoHJq/+FbRMHzgGTr+yjVCpLj/CGObFkwVrMKlYdwNXn7pa3L2
XcYbWOCVOXvfx29wpWgagE7Hp8EehHb6sd+ayn0BA3v4pURoV6Ic2EZlfegp9mYB
8BY9uaAFQ88jRYPSZo7W4X9NpJ4YZ4Gyxf2GK1m3p9boRLU6usN/tXZ4N7H1jlYK
kjoFku0fiwHA5s6bsgGQMt9dl+i/urh4xXDph8uTyX1w+e5QKl2WXFOWfT7d0Got
mpJqb95vC06uDIJbDi6Mxo9t4A/v9Z4dL0TZfvzI6Mlo+vfaw9iQOZBrNs45bb6M
v+BzoZVFjsbBhtoApuZN6Tkpl1A1kevtzCq1vNC6MJa2JxjyxyzezwWq+tehB3W4
3NUv/7W6Levqn9UEZLx6Dg==
`protect END_PROTECTED
