`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KFEUlhlNRxYe5PXpfFMHoDVPcvGK2FNsEeqHL5/ulce9v8EwYcHtDKhsJM6KXiZl
UxhnYM8e9ieaB6hXka6DyrlbbBZ6ahl4qS1S57JeaYR9uyOKSgZRTAMDA8zFGemR
tKVrVRLVkIaJjXi2nVaGS8JitjESIgA7qSTK8gSdcGP4E62AhLR8ntZ53rrE9XBz
USwoFSAV35SFOuhrHf2TsfY+BG+3Fqsgc6heDXAS1KRaMhQ01C/mlvC1l0INHYJZ
tkmZprhRM8NyNF+x5LrwyL7NExO0jnET4rsdKlZEJVlJmbrZ1suEpmi/g3mjPgb3
9FDPBISo/omlMm0Skpy4hgna17aVbFJ7891kXpzWp1KHlTLSmXE6tExdETAgQ1zv
7Ni43TxpuKmI5iMCAku0U/UeNIG/bJQlkvyBa05IMgY6y0tAlg6lhdvkKPOxnjWS
zClVRjv93xWYLcR2XRpLm4iQBhdMxOAk4GHXK+3u4rKqYUm0hOGdz8Ta9mlE8XCZ
7NiA2Vbt6a8HdmrZwVmaHQgbZTabUaDFscDGlJDNng82FzwO8RwF6KiR/qqwqxKO
5Eu8dsdoRjlR7Q8SZEkdluvJTatzTZ4D3zOLKzRrCOr8zeKixJ6C8gl8hk/NM1bF
dhzPKXxD7aeMMTzLFoMx9WQOt9kxgAPzfDfBM8FrcD2N07SH0uyyH0RIbhR0Luns
gBSxN5VxbB2bfbws37voAn3QsskriG0QdpqJWQKvUiSAw6CBwiCm0uHwDXYwGkxL
5qi021/Bk1cHOE+VgrVLf7KxLDU+CTus0ZNEtpHFl8/8OEXQpYG7l35hMntMRLOK
Vbr97jinYaIJhEyskn/66y+c1d+61YGp1mCFChvoK1RgZIwgvq4o45TklFwGDL8L
/EN2uYaEDvkNlvJaCY063oieteb0BG34QqOAQ/mZUfnlW2zCJDq8yTOdccg0mxh1
q7QlykskAdBTwOEfhxEgW5LJ4XneHhCgPqrFIFiEM2Cb3vhRYsqOGLN2uDnjoNeG
nvqncNmmwsT7Tx7999lGRPr4WqXN3q2jQyZ4ZxM00uaUREr6fmLM0W/vWn5y34Bw
xh/JVVQ5D/CiYU6hRnS+kBYVXjiod3YdmVxbQmDJbsXeEhWlHWSxN5ULrD8rDAYd
zC4vdKkG5yqKhkydQvPNABbjM9kz3Omc4mEdazi+ghPTSVovnCn7hy7UcJySqwY8
SIRRJNKWqW31++e3TgMbCykaAEGOljc/BUwD1VQTEc2xf53nN3pChTbBrofxhxyY
TP8ERxKHmstDQtjf96fYVsARYcJWxnKirjGX4u+RFMIxwEf+OVRW6vmdOR1XMpPD
/5RLsi4fFHOqncvCVuU/+f5teo8i6Pol12GP53o0xDiF6dw2FEdJ+4l9BrB7lZSH
zX6tosz7R5+kG6/XVGrwg7wEn8ILM2tASnRkEaGrvOZb0CWIsT7rM2Drzw6WkhTL
IbTOeVbOHr9xaDrUIZROe+h1IDOloFw+BOUuRHaZqScFxamm6HtRZmBJbysj2UKU
vaMSQ+7ItMiKnDnYjFyKWe9vTeoRsdjsYphYQ9+KuHC7cBqpAyTO33/sHo3Q4W1S
IesxTHIXY6TvCmO+R+3ITJ/jj8A5Ii87aI2xlskSeoWZRP7fSlEZON9V9KFwYMUv
PudTxHRsSU37CClMX2GUwgQmj2mEH1c0G91DciYdjryu0rGd6xnu5RAYfaGX1DAN
DvI+MRI4gQYR6xGIzUQ4k0x1M10HuA/qd2ckB8RSDn3GT5BpDQimA+eRvfzoarZ+
SYOdlb+RpKkMDKdw8rNIIVH4ZJ+rRu4JH4rw4C1INoUCPHRK+dZA/hoOdJZZb4wX
xUHVX1wQUTnMohAsZFRbcEXi1v75YRRpii1XffkSxkDyzDEi17WL0KfpZZ8tdmvW
UDc+xEg+ER/Cd5ZiT0xdXEaMXRa+wAEcXjppZ+lOAMymCvGPRJEPv7o7LPAwnCHI
tkVS9lsNYQi0G2IXJeMNDbkGjVeW3dW8CF4pwlZGpZMotWvwDQEq1/DKeDy33wvU
PX3RnQ9Nl4hW6JDTQaNMo3Zd4Dz4SJPdXUI4TfRB7jwGXzwfeFuzvB6nekp3xVNW
4NHI5cgMgr+ObcohkSwRb4wUiu2fW83BUEemYfYHuPOe3Uf8cQ4szLzz2JV7NDW6
Ba5eKtIupSSIGUfp7Zehlf4dxl/mhqTih1epOTSiJr24+E6+5iUCa+mlSlnuQxRP
LnOzNxCYNYVI2eBlzKBQ7WVuRuplscjM/l6cmD2qxiwHPSLc3SLsq8DXb4952+aw
DILIpx94MC+qFr8HGhQrH/KhMRnHi6cnjjP3gOTP91hjQQb/gP5dMC7XDT7UCT1y
VIF3S7TvtxVCzugkfOgdVPv/z3KKe8UbIHu6tqRebV5lZDIosxoA8k4hmwMkGyFc
Clz1T+ZkaV7Zs+mmbtE9R7gqilsYkHwPzJawT57vaYJ/kasuUuePza9JNDA8w2nn
Xcc+U8Z2vAnPdN4T7Hm92l+HnCoCnc6fWizC682QQ7Fz4JMOvNH0YSb3LnqhZwNI
lmbf8kp05gWCgI9ZeyB+KvPtXA96TAMPs9y53SZdApGZIPwhSnTDvoq3NppvF1+/
IlE1VAKQ40TGHZft60Oq3As41eswBT8F9E2GV9J02ilkLLzbC+4v64p/xczx7mKV
wLwEaiF0n4BqD8iZW1vCRajTs5upM5L4NVhXBw+cikP9E42y0WWscejdstcyLjeQ
WYtTd6qsyZlujEM1ohnSEwGXm6Lce0lSWC6iWHpWYYuULF5Xp8s21u1SOWUF3E86
L9PRhTURU6kg+q7wo1Sr8B45lVx8J9+AA089+LFbFFxWxKGfcDlmlUU3R4R2/GXr
4PsRs8wTdZiSLyvjmg0oOoJYZMqlgLfM1X85xE657fVP76QDw5wyPg+R+myo70C8
JCwaR7uvJOkz8Xk5Caks5Gnn2Y18Gv7vx6NAnMBM8bAA+eaVJgMZksKmFqzHX+Ky
TR5YtYVh+yd4tPbqt10PkX/MWKcFhbl2fffdzIq9VNHu2uIMAqTFbeFgqBL0gfL6
K3Qx4PWgu7zwGHiXHEosSEoEXPtW5OYtJ7BMXcfenfOKo+PAglrpEXv394RR+2yx
kvupm5cpYplNXzEL3fQ4g8Io8Cfa+t9mxbhoaFkepldATHWVe9F80nW1DRjU8Ncn
O8ra7EqQNvPal93rRXQRd2oUd/l7d8ZjB0etvozzmekjXcRGUE/vRkPVRHbAlg8R
eu1L/wThN+yFzt0/aQRPgP0o7QGIl2oN49gP2TCoVjGf3SRAAYgtGNb04Lv9eBud
WuDJZ+346GXqAMjuj94kVW1UtUhrGSBptoncIdJ8FF5nU35PT9EDP6njeObqoZXB
+myTeGmec/z6uc+7q9NTRJdJKQ8e9gJM1QrMZVMu2J4qpUC4LN8W4MyPiYTSGk1x
uGWdOimNMxZ/dQzLHXKbLzMoDqPt4BYCWwLOXLKbUWfAP4CTKbwoP8FpX6xIFPFg
FtSmweqNRDKlXas/UaIQ2bUsIDPBSgtT69DgX8OI/shS/yRYC3imCjlZ3nG9sPO2
BHaOnBAOP+h38foixAsZpfn+6KBOU2oVpyb48vF1weJPx7wlpsW2FfRlO1GjFLKX
qU3g9hr2J9XoE064AUlD+Big9Xa0RWvbE5iHNSTTbleukGRI4m5IiR2Y/f3ln6L4
cbjUMEtNANxONsGDUe4hbOeqyHtaMvdKI7BLONz5RPXy5oIdgFbyhIms/uDjZ/0c
uAEx/9zIBc8bebv1OoSYqC0/3tQMDUFp9bi5eXZXxIhF98YxbFrGaGb+9p5jPylJ
vSfjasiEVd7j2ZMPEL+xjAVftqqXef5mcX7LDSkoEzm6vyWjAIJ1lwPi8WY0H5NK
XF26jZ4iFT9TlJHvBdqe+AXGNP6Vf1Sk6x89IL9L664WzSkvnoStL+co2bni1Wp3
rssobwEcGrtJaOfVJziTJ3Dn+qnXTmoQnKFDvvvwPSH8G/1Cxfr6/rDvw6vuXw1q
CMqN2HC+rNgpNTClfZqE6MWTlX+s2xaeRQ7oZS6zwcejY1edDlgx+aAWw8XWBurV
0m3ut0uXprSRRIKJqwIxLthMnNlL4Ww7tdxUX5EjSFgedhlGmrcxDy1vXf1CNhxy
Sy1MzDNDhNX7Rf+F8ZEjQ/UcrG9In4/r2LMDN5eSrvYpxehRqd0Jjr0oWyYtXHh7
G69y/t/GRN9DQ7W+DQYuchuPXAVWbrMjxFbCqObzkxxvfZ3nKoF2nfKTLeT5qVeM
N9B4e81RE/12uH5ljagZRCaar5jKwiqdrjRflechX4lR27Gal5Qnj3Aaq6qvW6U3
3Ojly5YI+hBivaC4fM9A8FI04r99bWWfCDEYuoZLcrVvzotA+iIVsc9cWDGZiYwj
pRg5JGVGkE6SxybuvVL3/IwpKju4UCO9iOSEyYUtsmr57iDdL2i/MeLT/QHU3a+r
5ZQQBo4lJ8vzRs0xJiSugWmr4RkgbGPzVCTWDwvqAEBz8JGaaIvoDuHKF1bxXbH/
/z3bDWbp4L3q20mFl9AgvDxNiYKgff7mocYD4nzZ7SXdQ0PkyJGMVe7Eb4qEPpgX
RiWKkLHuYiMl3UmsBJViwwGuHnAsudxSGGa9uPqXuX2ZidNMwyO5ObFGPKQYlBhM
GR2HI5GOl+MpQrsVpUgkJ28CUS3ENajdM5GW04paRSZhY8WwUv6y6sHgrc8HX7i1
HhKJmXE/kGyUsyot/btTmvcx/CEzJLE2DxK33p+FEFEp4EEeSON1mw+CGMpbgwi0
F1qL0urIRFw/FO7i0g/NS03q7eiZS9/PE/tqm4QPShTJhgLKV1te/uzGGJuCyek4
c1Mmx2k4CYJi8IFv8RQ55D7j8gr0pyMf0nIFvuw+OauJ+hRL1PgedqPig4Qmisqc
KxcejX6QglCVpn0Iv1ooCgo+AfCAewmi6a4KEwe9K3jap0viZW9z4Ekvi3mPte30
65cAuf5+qtb80CPyGKEUik5ng4gXv0pM10fKzSv3YHX2dI12ky1ijfDNosspOfQw
0r25N+OWKUuQ2rLPd7td/WdSuU9BZMhfGdgAg+sWPy3vQrVG/zm1764ydTR57nSq
90XpmRhDPMuEOpe1f59CLcqqzr05AHn0o+pQkLgzzZ+wHPWK46KFpPyQ/xbcuCoQ
qOQ78B/dBx4uHSvv1PRz3xiXWBHgEg+Wp5+RYvXPdWdH7sGj6S41ct4+O6tvsI3y
ZwWd56Qd3VqqK+O3NC1abGSiMZhaOoHe7Eo47miayn0OD+bHW8/sOuTVJ6YvnaMp
UuHxsnFSNcQsuigO4aBLVbmA3EII2xKWMLEFPMwEnoDV0bLp0XOAqMCa2JnngOKY
NeH3sEZpJmhE/GxtdUx0imsbOJe7XEH+8gO0lbThquIUxbrfIN6ZgXS3AZjZEWur
7huUKIfOe+pe1Ood7sZlRQ==
`protect END_PROTECTED
