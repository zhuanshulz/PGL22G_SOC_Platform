`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q6Tkuei1fVMOlB1SDn3OrrJR3jfm3+4IkNjlwJZjXYQhjApKFKqdZ4XmfAl/eebl
wDM0J0jd793gt1FsG5i7wLJ0HryXDmtesKt9yVNg9yqadB4B/6qIxPSusPAdJ1fm
Hw/bv+oyxThwX5um6pcB0OI2wAZMmGIfpB+O19F6zvC4hofvONMqowK9LZhl5DWF
0Rv/oca4pq/Gw0qdR/bWSlKRTH2kUQ+w5bsLmh9qZAVgol7ZUQO823Um82CQy7gY
Api3r3+Dqgj4t4iFx1XSOOFEBzFk44V9t6yinnlI0sf0HDJDf3kffeXSyEhBc0Lj
OdabcYIImXgnC1N69OPsrngJQQ81tM4/Ta4dkCbMoztRcpWrFluPjsnKD2GuTtT9
iGft1VkQ9G+ja0thv4jqt4MWIt7ff34/u3vzGc9YSGE+D3wbDCx9fr3wB/41lBeq
RclFu+P0ZcLX32/Jp60z5gdRyBc4fP0KWMF6SGLg5OllBaAzT+7JrbsLcej3N7fn
QQVU1zrK+wq8sDTGMSoNI5GI1Brjbe6wmy2vPtvvzBDjeGUGBeJq479GPVYPxDrj
OegpewO25PoH7EiFz1ls2WIQ8rW4dBOMRRhlj0K+t0pTUSndKevtjb7FKGLk5b5R
PZCN4VMBSHnz1T2IpLjhshJH/CjPr00PtmeyKP2cg2nAb0Nr+PIWbHFoVY7zPOC2
8E26gQsOivPAPtsZkhKIyU4osKELHmRsAyCZX7AywinDVslVDEl4t5TGrcS1Wx7X
bQz2/Goj/lGhxoUvpS2oBppzLg5bAEpuAiKJ48XBkOUv9syVOT/rzmwZZ3eoRpZd
0haRCDvVZDSwOj+in0ik+ZltFVVHUs1Tv3k43TnViOTY5DzBw1VKHXwtG8Tivr+N
/ZItmY4NgNyO/6CcpG++6uU2OXu9rX/bNKpSqPwF/aLg/sP4p3hp+cLZjHl+kULA
61HUjFWR3kHfWpVQKQL9ZuQPZzswXUSx2P8cw/Sh++pMHTZd3P1cyJsqaL1i7jBi
e0zDnH/qgPpmlohlBlKbXltJZSKzgUOTNlA8/jsUqrWITwUR2wXviPZtthf9pJGp
CH/bb4pA4wxPeQ0qTnk5SmfUTSNUgIEdGR0vNdbBYCjaBFzikhvoVL3sF2eqhJHs
JtlbrpbXlGksCEIXhm2I6nr2iEQVv1qC3knFd2Md2+vd/o0kwKZBjk3b68SYvC2z
ue0KVIlLwUm0q9uNR3sn7+4weqjAGLo+WCqf8uGhRp0l2YDkU0uAFDiAWyz2bQpt
JLz9/RPmbncai2JorON7cAjrNumJsWdDRC1CxAJMNe6jsSeHGbOhZEwwgBdk2OVy
lP+Ud1/5SQfsvnfdSkuylREvGo9dIDNv6QmRUSCmicHofi++LzbuFONFVkeZZOMB
C0tBeymH41dt+JHWykDh/wN58FSzef7Ezxg9PVfQRpMrNeT2pCV63TAnNSvbIa3j
E1DLrMLS1f18DGHT/0RIP/B7xNUHX98QdWTzXuO8KUgyoZKiUuy54OgOBjYYI21C
QPJ/Ay3NKM7M9YScaD5mep7MdJbDHGgR0t+Jg76OxjTSBA6bmz+/Rmc4CApHU3hk
2LK96l5Ek4QPBzGXLh4qBcWtUyFsULyCJL/nF67rsWgBOKlZ+djqExhvHx3tLdv/
kAh0oRu/ZD5+XfVmy814ZBgmCAzBYeAkcr/ENPP18CWmezHkPSADesGnssrsibH0
fjEkW2kNARAoRfRzi504yzE67FE/8ygHFuc0WibumrKea26mv1RapeLWKchbixum
MQNL+yIkO+2Lc3osWW14ZCGHcqJgrNIm54vXLyuZ3AhaUAidY4coVIl6gpzARtrG
q1QvDoiJSQqOGtVWwxCb6uGJ8/GAR951azd/MiaZNn8hbn9FemvpKqTLggBrdOrd
mw4/GH1W6JZMK82Cf9shaGHhspnr4BcI/KXibknLUi4Kd5VbuH2qO1TXr3l4LVEW
6QmRJqc1FI4x+mfR1tTc+hyc3XNA+dsgPEbpWgn8/LPdkuK5Nqzq+0aT9K+m9rCQ
ZBFIh7yeqFeqLGS24bvIvt6NmCjqYsX9Dd5MsCoJiZNm6sOzuHq8Bu9Ou5J5c8eC
4lsyUU1YKz9M5q+VVCzbC3X5DgDJNHbKbNWVpHG2ppErteE+W52BLJaoHtuk8xHh
YczI9l5F/p6uF0InNqFP/jv8vZ9rRqwsWXOmc93bPZZHKf7zMHR7W4Y63RILoGjl
M8z/u/3Py5vKOcPji0Dws7WsjDiHfjYZTp1lf4+bBDJhoozo2bNVa+zp424OMp2f
Vqs4zrJE4y2R/dEFLSv/ff3ZC0hBQTyA1B/YR35OUFtFBQvSWYExHgmU2VcrZ+L/
euTGTMaMC8tMmgrSEuC758W2dq/nbTabTesgfqzgdTL4uR9jqnrK9Z89ZkNUUn/5
DLohmcUPpBYDInpVwFQ0j27v2O86T/iepl7/A3AHLy0JrT4WFGpW3eXKOlBkTfdV
mKabFG+d7unaFsMWBy6wwpGpZ/3H7dDFkRhVSxzG5S4DdrD0xp9/L9LhGt74X+Vl
GxpBrTdO04Klf0ZDkAi3k+9/8sDjWalvupIQLUOz6yCOQQTEA6pF4UafrmXhBjKV
Xm4AuIJdwmUO0ejok1+vULQfWneN3Q4K2ycuHxfcDB21E484wf0pLgXvKuwJd1ss
hHClBGReFXHocbtfuuYTRMl2g97hK19VnrcifdxZ17jcJAyOXpRo6/e0vuY04VJ0
UgxQpo0D/0rf5AkgpYlbgxlObQYVis52O6F1yEIQLIJvwuYPcc1m8VMQLnIOb754
fCdYLb6d/PNfy42dESuDik8cFDB82mRqrbKgONUaRoXks853Srnb9DBO7UtJbi3k
RRHWwEeud3egLRJlolwT8g8nbrBDDYMXlgtnSAMittYA8a2zyXMi+3AcVd+DeqVp
7pXoDk1AknRaJSYJQ3zfsC630+5kUlz8RMWJ4iX/slQEZ0cIqZGVNA8Tjub5WCdq
eP3mKeKSgwE1j4raTlWK1itfaQ/TMSTkm/BBOjkMCIoA2EKTOq7z1j4eCemAvHo5
XyryMD62xrEwgzYJZVLZ9Jau1t+fi9WMIeoSaTOo2hUlKCGss3cfX7/84ATdwx3S
PGfEJ0fjw/JhX8jMriblHjbbTy5TKpwfwyZsFBpiLf2SKJaR00rZC+DnP/vMHO7b
VaEHgHJHfiriK4rpezzKyCznW+US/VNDsBC6ZPFjFeEHCd3DGNmecxzKVhck/b/n
ALtMGUr86DWfHOWqBAKzunsxC5XljJ9ZB9V8f6FjFVTd0Bko865HQYIsHs0b48ne
zH0X1beatCAskKWOxLdDVvejQX8r7jeFqCbYYOkZ2Tef2WWC0VXIjY7xfltbDJuQ
elkn/C7faFOcZmZJ4wLREoUVgn+zIfqilsD2bYG9fOmx+2VyJyV1nMdhWySnavqP
wOsyNuyJZOZ5LHKhED9G4bdfQMLn/hA5UQ1CoVFDbbuQ2YxlaXB7Kam25P9M2LMk
w9jpWI/QzXbj4cJjlCG1tlNsfSiiL/J6mPTKIv5vdRw=
`protect END_PROTECTED
