`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2hOGaxuvlq/GDSIcDhUOL0EkAprO/t65N6jAa3AUboFIdDGmU7+3jE61G1eoUjcC
9wE5DhTBbgFwo62vM26RITov8ucSoxS/koYaPA4M8Du4K9C59T12LPhH7qL3koZ/
OFR2QgBMDJkmbRDSWvAGtnUSoWw3MQuqCAZGMEccl2+XcndLfZG/HgnGQSTPhGb/
K/V0WXJd8H43+HnVHWWW6j3n6KuGwW1IR0r6EF1dCm1ab2JPKtfia3XMeeHh7oul
TySqmgVnLoygz6aiWan1sYnQH9JwQEmaiXfTy7CYgd/UxwIxtGWdetYP8YkvbRsB
iaHPrCwO6KFpAa5YCUs4UjQveFZ3dGWVqXj73CFDS+WU0fraD5iALi+zBRfwtLS+
JK4JGn8iRtapXVw5+qQElcE5S8vIia6h8zuCwTShUofOcryy4DxHRM2E2JDjrRVZ
45/9C3+W+mbnZkNXF+IohSKkw9sqZTzqEwaBwIJGtKjQwskGgfDBukOctn4WnmCX
Lter6MvoHS9FPHiZ4GBRjs5zLq9Bg/LFXvCRKEGaIj913kcXZDC29jJjBCLih1lk
9bIsZsmaoDHLMpeO/xTt7w==
`protect END_PROTECTED
