`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wCiX8btTpMWksEy0Aw5du1S6OXP7V2jx04yWXt74SccjfoGf3+AfHCZz/QnGRWeR
Ocu7pLSPYNQmABW35B2l1c6V3AbVbDAitDMvRx/GNS1nkAumOUD6wrK67ka933wI
/4RhyBmjXMae9V+AV6RY32R9TXnHeH/DvM80618U6JYWUBkUOiSlJ+if4WkKQNh8
tnlHrqu4GUDIOsw5e3YhvmfxCndVYTJaXNF7uhOdrmKqNQWy71HBE2I4zZ6s26al
XgQjC0ZSY8t9fh53VLyGl65XDELWs6H6/fT4Yd54crH2WksXUrB7bu5fTZGon4vL
F1626aZ+pnRiI09OrJ8CpJZxDhJe+IwneBLVFz3VhhjIEE7Q3ZkfA0zz7H9q0NBJ
bNtKwANBT8p1jv5hDRSvdVXXSmSV5nmYm8m/ThHR6cM7v53xI9f5K9/8Tb68Q2U3
O0en0vsPHToJ0xU2xjGpSwwhZZhHExwPwzWvgxGZKZtsVt/jVN03HkNASFSRygYw
Y+BeOgPZj37/pVoMxHHZZHi3ay7Fbmtwx1935Hcs6S5tapYXeGgDz3pV6BLr9yGx
alEyt2+GY5riHzHUfA+pN/3AB8nhLE+erbg2a7Ccjyqvb5B/y8DVesQwSeZbHHhX
63NdU3BkWwWtbOYEg3GDk2cUSv8wNpD+TWHw8Vda2h2VpxPyP+2nbqSN/Tp/Q6TR
pLXFeH6NqI0fw5cGZOGrO88pNrXgnJCbkoHdhzasDUUut+vl1zxFhAHGzrSk0N/m
WYV0z7Zurz/zOhL+UaIAXwth1UrutFFhwcqDsqE0M4LfaUiB2fLpHJsSXQ1t9erR
m35TH03xEABuoNCqSzscNwVePc+fCJh/lqI7AMUhBv5E3cIhuI+3UVg4jFdg1yng
khnYBGstc1mSQ9B+MQdfzkffSmJULURlfCzjd3cev3gb+gfCmWjc9CTBEvssyBAC
yqJYW7IrgClxUBTmnArBNmMxGzHOgsApylt1pZSRlRfmCeJl+ZDuMOjMl3LEwpt4
Pn/lT/wiS/ZWnFu6VTwgLZS8jQI5ozf9FBzigc8+OcmoXTfudvz/m9u/FTMmc2Bk
FlD4AlMC0TXnCYY/le4MM6OFKMv/YJ9Ae/HJvq236qMhuBv8VETgYjTy/3Fl1fdI
+fJsn/s9p2XiatStZZsx6ldBPlXYhf84CitM2xefiE6NyuAwRfCr7tV85MSvkm2G
6IJu2z42w31AreawVrYilmFm2JEXRFage92I9dCZ3k7dHk9eVMMoKsga7XBy1OKi
A7J+SFLcRhzq6WTQBRZAGV83WhVDL32qk0UlvxDVIkgKiC6A/5TE7/KeQKeAq4TT
YatXgNdILqukLRE+jVJdt5IQ5dYuZw/GRcrqmfDzLgFZsmLr4wGtx5UOHZhRt9j5
KJf3E9ha9ccqNb9WWRwEffXxq/ZlxSaQvAqF8P80bbf66tKlbFvMUGagJqIFV8jy
UTGVGoIFhoGrLPqJSefotsFuDbuWLlRuD+L1jMhfhM8RzJD0dt6CxWhYAsArG97O
/9UmljeQqTS5xxskjpmg0ZB+LRAv9g4LuEwgxQ4D2nsxm3zwjRWS3faNZEHDUVu5
30gldjHT9fWcSikYfyYC3D16P9AhwQ5PBUP6uS3NJFkUOjPCiZvz9xcngA3dx7YL
6ehXEmzDZep3dGo9xL7IUE1IIeAzMsCWlf94Eps3gS1SxMyr/Lh16IljruLsZbLK
loxCxPyU5sId8j13bTCfDWEoT68AMdinprrkDCm807FjvVzV/8Mg7EHm66j62n/q
LCo82y0U/K2+yCa8g9NvvuHvTq12jSovQ/QGbYKpbCbl802ymRbHMfwM1x/fRDb1
CGUD5N6LgWkbDCy40HM088jIOEPgXCPTSaMFEYTHwCK94R5yAfNzIP4Zk4KWRUo+
iubSv+x2pd11RDtXFKjBV3EUyBCloz66F+H2m9FkTU8POgZxDP5h16H9P3+JmkRf
1rBrCVEBEE1IYOz/DDhvVdvecWsEER+fgVo4jZr9LNzujyvDeexxtayrZquiPn4p
k35LjM2D1FE0jK/PJHAHira6w9IUJ9xKun7/XIafN75bTqNgF7Oki/A4Yht4RI1t
iw/eH3Phw0adbjZcWu4tE5ytasucTVUCC5myeelsyWCVwk3mOaZaS0+irJV6La7P
Xc8OX71jKtVyGpO79ybnYZtJNEXz+YF32j3p2o6ianSyr1N1n8WlIKgpbAQxeMEh
EFxZAxJA04vmaPqHQKN5Z919PgmWeVMu1B/GMa2KycY=
`protect END_PROTECTED
