`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
udIEsw7a9OTmJyMQ0ataBMOiK87yLFQ0zp7QpDPi6LIHW7st0TwU+Uoaj6nT7qyf
2n4mPdTOxPKZHsJba8RmA5zPgREXrN3RI9VQEefqJhV07fjuz8dbdSXjw4U8sSU2
8OuTwyvnC2/vBG8UTT0rX1rakNQJAhn+RRbKteeqOW9ZqRt5VJWtdf5TZMJqBL5b
H0jSS2WkvXSdWA9Kc/63zbBUkoTqLyhCW2+kwBtHEznp3Qu5Lzka43jgTOXyZ2hD
GolGxr1D8T/x769Q3GcDMM471dDwNTtnQNI5wzqe1Hre/ukDVxWV5IQDjlZvjji4
yUviAodXsUABdPEgtLzGfijFRJukfaHEo8Gelgm/te9oYvYlcrLG+6wYzt/7m9eY
erjFVifcCqLurxEyl6KzTlfKGv6SV/32SpIEqJSYeq6q/oJ0OW7ChxDR5XQZgSjW
`protect END_PROTECTED
