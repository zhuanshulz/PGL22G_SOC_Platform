`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I10fqunOzj+QqDyNcyC9/NKkY9LhcdwJk5YfceORqOj2i+0hehl6CZSEiNf51KsN
7nZVNOB8FBVBCQDUfq78do3SZ8YtObm2vTCFfqMUqpk7URd+ua4+HN8Elk2BpVp/
qyZYqDQvg9EeaqkJTZ5xXMjn/HpVJdv8N9jRwK4iYZX79Yt2RVf4+9FN8YGFKNyv
dbjaBi2yFPnxaQI43Zf+diljwI0UMAKCq6JsO6mwHKRqoWX8glSel2LLP1XEMQap
/flpyxRVur2Qxeymj3xxZN9SfkIiT1dIZiZBzuHy24UpU+4rqIN2aEQLfMozHvg0
+aRjB9o62dO6GuhIBk4GjHhn0x+Z2iQgA/FBJNZahN+sB3VFz9brTGJYtFaJkU1N
FnxoEkIqH6GKP5qhta63raPpN3Spk9wkauTcjacB9QxH4U5Pj6O4+YW6FnXokvZm
ewkHRQLrfHJMWniu2WbBL14/BFbHhpZNZUzfYQlYKi4ShjbAwepl6/15CsG6+vU2
a0IlwAhm1GligmeWCYnurNM6//C9QMbSTaz4rFhE1MO8IjOJyhrPIJCB9G+T1oHy
aIEgAbBsWHFe8WoYa1OL7Zg5B29lztouL/W7V9h/JB/GXQt+YNzDW6f34EdP1d80
y8+vT2dw+FfE9R7Rsn9e1NmDi9WmMaAkBdU74h7EQqmJrFWCnwTBeiGfaTrQOiFe
fhlD7JHZ1mMAXN7CDMgr0C+bR5g2EkDWZuY1WC2aZJFLuTHSc9gWDeHwCT9/E0WA
cbhRxNLLsVgtevu4bbLAt5cFEkROdAszq+PFdjSFIMmq27f2LJo6DI68SPvmqehp
WCgafllTbKfnR6kApTAvKKLZL/4gtF7svkcw2yi9sLhwzCcVSTIJjVMMd+Cg+r85
UIzpQ76TJUjqGrePVfqRI4OrBqelz61FgglfPTmZXx+C1dSFVvC82zpwjK3i3ARe
JJgPDYCDhaqTdds9kTJiF/XQ8/GJWVciFDIgy6o1NnhonT1qABFZe0hzZQYg4xzF
DAPdCwb59rsnr8wmLgLBAzAYbnYMYnpzp2L0LxShLGCKybxdEevnTZcs3whukZYK
7/5yJt4kXhgTmuHzUb+jKDBLk/+qW9TbySSMe35DlyhHMxO5/UCBwvtsuS3jKiL2
OBAG/1RJwp87ezE19O4kWqcws/nMu0vms2QC9N7hj17XX/lLeUE2bnnLJeAU0N+P
0LHZ3myOjaHCqfdRKBgvDXYP0mDjRkCPFWDr5LyGodNRRj87upDU5AQQdr8owBay
eOW0Vs8lVD/vSzWV42e55M1a7tmcC+CiCE4StkBmLod8hXEr7BkmbkOvYcdaqx/j
YKkhSxaldulAawiPTcgDCgUBAD1GNR3hH0mSJaZaAlG2tlwkrd8gvhXSWk5QqQEq
q5OJw+odKqH7ylBATjTCeQ==
`protect END_PROTECTED
