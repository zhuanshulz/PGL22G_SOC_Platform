`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MY+16EejO9iDMnTvp85Nt+4ZSK6C6o+Jrq0BrZERJaV9nd284rHdqLh4lAcXv1Xj
KsqBW45UXoNqiaLZjySC12d1v+g9UAqA963GnD1iZQH3FdQ6Fq+lFsb2XNiPMEDi
JZVB1v1g8UCUgqC3PgUdcWM7wUrPaeUrb1PEytFG/z6YpWDNPP8xVQum0iJD9H6m
1zTkiPz7CEFbXwn2YUcZSQ06MbXK0E6/pIz2XQNbTj5rwOdNflf3C1uxy/+haHrI
QuS+9eHNu5HXFSrLxUKOgXKudNAmueiCX8QASrxfh4YYxrvC52mX3bYtXiaJyj1i
Cg8kLWQLVkDTWrnGjMJVi+WFN21GP2sFMACidIqSuU7yWbEFuV+8gggaLwz3tZCk
O+c6A5PF3TbTT7yewinDFvJQGgFpV1ftGHiot09NLPOCnhyHZl4JEdYYpr4JWz1z
K55v+6TOS5gB8x8cMLcgrVlo3CdhWwEGRT3qxFnWVyHvD6WhGTPP1cdEuMv53fPJ
/PR4YIjtVP2Z1mD7sLxrnkuwzyIGIYk72S4ky6QkHj0UFxnjzzb1cOQDZJquCYFC
plLOfezcFHjzdDTR+Sefxfcp9F6jSoA9rZNwUfUoR4H8vOZQgCNzDO529igHzndA
B0VGr+y2BRfi8tw4+Y7yni+w52c673ihjrWJfYiU5xLipzkDnUVETJqN/fvia6sc
H45bHIds0y5hZRplNJdrhf0QniBOKVa6J/W+HDpqnExZOEUi3aqCfEmo/JU2wVgT
FvW3lE/K6pQQ9dtJ7dC3auINFGMbB1mf7T8ggfiI1fFfWuH2nmkJNhtKiEwUa8hh
0c0823H/M8VgzutzYcPOUOJvK8fLPEBX9TrNZZB9Rox1S2iM1/DeospoLt8RliqT
89xZn3WQj5PLQzgViwXPnVBWb/iClcXccM1+TMVlkrg9rkcWFwkWsdXDbMMRoFa2
bhWtcMK4PJJequzz9M0f6C5Radj4qekpV+BWdnXmbIQ7LG/B/tVznhK5lKmqRaAu
eGGWMOpxnIOVXlWLw/jVqjP6otccR26KoXCL3Oy3E4R30PoSTuehBokhWYk+EDg6
1YdFzt/mV4jVJFOwNcaDYbnprwKarv3PhyhngZlfFuM9ep0H3bm/8IHj7QYphMcs
z0KVp9vRsBT5n6TfeDJvgOFTxXTGk+FPLBQBKndKJ9mSZbNaz3Cb3K33qqH/w1j5
pjQ8ukLQFoYqQ1+MCPA/XE3s1O69D6ugM2mmFST7phFqhBl0PIQdwRjF81SEHao7
yEB28gEZZbbQREcFLgTPlVA81mZEFhq+eDgKfCAVnm0rWIpsKvwtDC1nmxBLOELr
Tqap2mI7gl3wa49GyXVX8U8ZVN0pqgKRIMgtpG31ZzXeCSbB59ZeQ1mmAe1zDM8E
8Te0b1FkDLPqbM75e25M9Ku3/gPNbiLxK+1qEUxD7MU6Z61A9donXheYQNZkcRz3
SORClTQJgYV+xqEzHiu/Jh047GYjKefvFP0EuXCuSXj4BQzgCNBHR7fNs6rC4+JB
ocn4ABzQ3HurzTrWCbKTQOZzugjiqIGM+XiDlju4RRC9C1WXeRow8CU7+RWuzqW1
Wg+Vh1aSybFCr5ioPEsGbfExsXnSQtWTmklW7gZQlAAzgO4X6iu+iZwZHYDxCbf+
XToMQEnLo0fRJwDvJhTpmN6mO+zqocBIYKXCUZvo/44M8orZvqkyMWSeSWT7v2uv
BtgI1lmxbAsPDAnZhYpqvqp94IKQPlC0ErO8vQxgq8QpxZN7ym0kBpkIaIkHG7RB
hfrI1EubDzTkj66s+XL+Y6mbAEjKGIDacriqgE3azYhcUL0/LGLQ0zyyqG1ttFsx
8m0EANvUHD2Rg4Tgkwe3AIUJmCsIdPRr5QnxLo42F65wJOAzfrlAGLchsAFsTmux
z7V3i+llHpmOQWEzxvpiSlXZPA6HW2dhzWZOV72GDvSK+er1Yqo58S1P2KPnScL/
EMrrZ03Ccp4oGu9LBg9q1qqyIGkGSyJHQJvWhCE7xSafFAqcOLDA5HlELhi+QF0G
ASC82ffcdj7wTHOY2JaMdBLYQk4la1gN3WrQ4Wxqi2tBxKHEgIG3HwE/4nikvg0J
HksMTx0MFMPd+Vdj8BGlRJNeTy2LEcHs6zRYhCZRdWeIYTnlMDbeEx7PGF8GYxjD
OR8CrD6FmShlhUTKmV7w4h98vJa5d0LkkNhtaY6J19FUhMYq/O2g2LGaCtJyswNd
4KuWz/77NKSaznLvMaQbmErvqXrw/8WZ9/7vb2fkHjWF0msd4Jt9NbptGFnYaIxr
uIZN9qPW6heaNTAF6rBUTyfdKhIKLezKe8ElzVjRRh5JDOKy4dKTdeYJZTCrKjmU
/yJIoJ8R9r3nzMBQWOO35MOtpHCCWYPsbaaI3Jr7ZzxwprZPhjRWs8VnNOVJy+8m
ZStNSXLOryng1Z60SGt+XlPgMdlIz9xww/PHNPQkKzqKDGQumzZT8CFPUB29NxYT
earPZfJBRPQzmXtc/smzr/TwebgJQGP65tE6rm0BhY2ITNjcEhPQBPNTImRfAIaI
jKsaGqqSH77pyqqnEOFKbIZzVZPJBSIaWX0H9d2gxbf7/604GBR6i0O5ECWPHBqg
ZditqT1fCLiMppA+XoZnmJT6JRRFS7b4I3Kt3nx1PHuBar1IGwngH0DqJsAaySdD
oXcuJDwcIIanEkmeio8dH3nA82b8JWSY2yXyQyoAkvPofoOgS/7ljPs/ex0DrFQt
dfiL6vRoYi6YldUMTYe35FvwUx3nfESFw0giw2+IIUoahgAjwXp9a5uED67FNgBs
hjDRfNyHpCItC/ZSOAL4CanLa6wPNJMs0TNJo8CYgPyBMViFpsn8PHsosP40q9T1
dkit6OtlHI/WqqYhY4od+D1AGsFfE4020jsFqTSO0kmmTPBOeELH+5smF1TBCTot
ywmQ2d0GgPvtAMWOXYwZAPC8JN7nU2asX+MT/bqHI769YMw0Y2X8+GuXfFDoNWgu
l3L/NrnMq150/rxdGo7u+yx4yX7qKMsubuX5pzHRt+s7RmJ+dgp4t0DlwskSxZ60
f2YOk2mkiO+dq9dkPOx2JYTohYQ7U3vaDs8omvUmAqP8xVx+p5prxUKYTQxNRpLB
VMNe89+ojHFApyK7/UaKpFKkKHD5sTZRV59TQjdNEXQKQEvqpCYkZP5uEkIzqrAY
LrW/hZhsb+Kud6QRdpB39Ea634HPix2ozHJdUMYFY1HDF8RPg1FaG1ckNO5cmnAM
KpYCYAjroQ2skqPn1xbIYWK2suorsJjXBsq/j/TTGbkA1op0fQeQsvWkfRHD7G+J
aO2C1lvVaAr8rrecpA2QsWND8rb44fOsyr0nDfgUaF03WIXiUGW3eKrnG/ClktGx
U7PKx/XdZR98TR8PdXUj1eW1G0ZRCPMln2yNtgPonPVXXBO7tMwvBHtv2wuRDAar
bSr44cYtDJSnzxlsLz5WB59CSlGlvty4rc6KNEdoktyLliE1mUeKbJ3/U5YOjnXs
onhNZRyn4IBz0azneBiHQ27JmM1f1z0rN1PpBUibyCY6AklQNcjeKd3eXII7AE5z
ytij7j96blSIjhaANeX7xMJlmpuraGWSefBABf6Hv7W5VQs1Xo3JZrYeEUARbIRm
qKVBAei+RhrBgVe7t3o1LuOUZBdThvQTm8xCW6+SEBJfEsRIKvRqP+zn9YgOoXeE
VUftAuu1TuccaLe/73nNqsIWzXuIkZtk84bV/YxGCHGeV3sTkiz5iqa39y9QFKMZ
HPQkaBM88TD5zZRIlj7fdoCkuKIwb6eY5TaCScYfFp+Ae7TL4JoS12qspgORdjR7
FKt2/t1Adk2zxJ1GciuJ2/3EYUnAKHV2II6clibXPMBGc0QNn3643m30ma/08mAe
Ej+KsCOLh7py1r8+zQGQmFytwoodRTjikzN7hnQC+AaNLpPRaK5voLSqVsK0HLt/
VFy+LJr3C7LYLfr4mHYBySyjx/rvGPT6ZGPQbJ3T4cV1mcdRHr/NOikYQHeRdKw0
2GlSm0Tg3uVXSaOqJyrSn1dkcxbXY282D3GrR3LqN7PfQ06JnTbCCleBb3i4yMx9
jHt6Bfrh6VqD83sgEqDxDUEfZPZHGeO8slFj+VEWGEFJwXD5pF6gbHh1m6I7RhPw
L6a6lGRzvTCLl5+aiynDJNjmEYdtlqOdAG/utZYVJU8ptg1lojUTtQtpaPwU3Adb
+VL10vXeiOcUMZxbRaohcNSFi0q/4Rt36iZY/xETzBLLMpFjPACAWSjFc4d7o6SU
3iP5dkhgXaUyQEXwludegvbdrw2U6UbFZP6e8wGuz3qQQg2HlTZTWU4oVaam59mv
x1krlqTivJf8RTj1tzivWnLVyzrxjMq8NABoJ4FEwIlQ2OSFM2Yx+M951qrJbuJJ
jLxC4s/2Hg7MbC54H/lBPlJHuKPPkENiBpTQPMDn2UoVUeA9BeeuGV4OhzVOqawg
TPnIpPX+JMxjjk2XU2eJn95sns06MZzTZmoKrZF32+vl0CdCkUojDO4MvUhjZJeE
Haf5Thn/TnWPUh9GJwVVE7CH9HMLduEYKUx0zkG46fZkDbY+MJfkyyXTYGv1njWU
ODfOT133m2XWtn741pTIPLZGFQ5sDAIkpMeWTwbUa6Cv5spGU92gQtZXDmZ6SlVE
fIz4eJKljryqVHK4Wjv/bNsMntsUzGoE6pXSq1unlW7URsP1MSA+P8sYUcEBR5+r
1/4n4/QVoWxC8dHYzTrVXsZbfybSlmvNp7S+APzoBYEHJHIXCzDcDRfvb7u3BnEO
Nl9r1FAd8gztWxMumghxg3iL8xdxtZxWUfgP6YD/RwPJY4K5oty2mUGePNfL/pPI
CkG60g1p+YnMqs0h6hG6YLqg7E6ycr61JzFchr29skxK7iq3Tmx3CVtIgJZebZ0E
jOj07/yH1AWdLU2PNpjS5zmisnAUWU7iH9Y6UNoXG0tz4GehS0f56H9a6qbITsg9
gAcA5iQtTl3NzLjmmGq0uPFY4y9os2vnECJCUwSz+mVWBo9NwZz+COcSUF9RBLvZ
wyLdm7WrAx1YKWlI0Vh2z2NxlT8GOeYLJSRB2Yzr2zUCp8C4wICKcvHGnBtfee9H
qNVQm085+dI81wP53aSL519Ct+21nA0VKIPODp3iREKrJC8pcrMlQV1NU2wYVEZM
WRnizjLasphzBeS0CZCpg5goPyEJkK6/dmYm6A64w/EltAPxFvwpBGg85gaQ3R3j
ndeSsOFLrtnzhEqeyG2DMcNdLkGtwU2SGXKvP9Gawq2lZS6or/GNko6hBssge2Ga
U5WN1oPiXp0Vv5B7WKsxC+XiEmdAHwp9WJCGplEhvBB7IiHCLPqyfwqho9WNvoFp
hC/yDDWG2LCmEBb7kFgtg6ORrxaTxvtuc53Ijv7e/i4TwDlcbamocQr//acL1HWu
5px3mQ9/lEsUmr2bO4YqYgOT3Zpq5Oabqa4LTgzAHdmoj4YA16w+Qz3up1ONwkZB
5FqK/kiiI1zWn8nsFh1Nu+oqarUca9d97U2Cb4jii45175EovX3OjqK7n8nXlzGP
zskcmIvAqESrlzN0aNcFNjT+OPYEhi6KLqbimVBi781hvrrHhtRWlSfC1++GsXYl
MT2mXJvHxiX/BLaamTVaO71lXXmtjcc9/pPOIMLwXIdmoKEfer1JBxAYDureO2mj
q0zXgLTwuGeR4P8OiYDZJe60Z5tKWysiUQm4xXUy9Wsl2SVRldOcvIt8zj6JHle9
x7oEtzIi8cMJYnb2Hh9y4kZD4WUhy0Dh143PUQ0b3sErVj30kMP6BPapi/YyWxuU
LYVfkd7sWopDzhoPeUtCS1re7dKsj5da4dzopOr+COCrkVACbBt5d02mNbyqRRAB
57V28OgBBVivnRVohJ7YSR+FNIR9kKCOIb/gg+joX0DquRBW4xxXlrzKhiXyT65C
7erjHkRdxwQgG/UPwD5GeoYj95phd1ZUOZm/irHrljUuMpzTh/I/G5F+xi20pffF
paNop3MvlKJAH90Zd+G/eFIj9MplLINfO18P1/6KSExwY4/IQX6UtgiYG8iUuT0y
GE52MihP3VYye4R537VJGXxYKOKmtLRaJt8Osbe0us+ApbKZxrjPd2taqSve/9hD
ZyC0ClnvI9+ZBfOuwLDt/7Ux4ne/LCKBZQ0vLMG6bR3L07nxK5bRftgVs9LLY4Um
h/NlrhRmdb6J9Yh+aiFSSMF9ZM5qYq75Fx/wot4lo7mTnMNqPoJBMkW2OcKcaL3U
l2hd04MmaxQQW8O7ZMuAn7dccVZ6ipsiXjolAUFIVg7i4tEYzH3fbeZ0v4a6xx2T
8/n4g2cLC2N9W1cWQlmnViS+5OmJXw/brIgACoTQXWXhVMp/XlDgUaKwtK7fqrTu
eCfm+yoac9cfWmPcWc5IgeBzGYqeaF26SLBtiYBQ4PIakqOTg6iovmSmQb+RQU5f
ARD+xbQAiRBFGTv4OGv7CA1Og+qUAigTHcgpD3It6Rp0ZWM09rO0AgqRHl4cXXhV
UJX1TxdT9wDphubzDa76Yq5VKvhCADSguIWAYSgvzTJqcIkUrN67rdRrw3KQwdyI
WCgDoVX+dx0K++MwolqsQhmWRZ6Wj4yvVTPoNTeTCPbpGa+a/+utIzzjxs1SYxvD
iadRDq/El+TbLk92VjFzEy0vlZkSqFvB2BX2bwe322c7mlRmuDkSjykmu0KD/UW9
EuDwS1k0WY9N7QotwCKzOFwN/Jr4po4zhWhPuFxGnwQdEzpwSaPSScl9+RD7uBnS
KTx4oVaJLEnry5r8majXUA==
`protect END_PROTECTED
