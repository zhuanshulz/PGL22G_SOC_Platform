`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tD2qICwXyjL1f656jOtORZjkq8ApauYp5MbjEpuVt0ty5wJKgE3WkILqLgKY9beO
NECB/O2/eOeCu2eh36/NzsbmLuPEOQt7asuTKvCdEr9DksF+7uk+ksZT8xMa/ha7
bYJOtjMzy0PFEp7YbADbofvLHYFDr5FNZumMapV5QD7R80d2qdI/a19K0fYWMW7j
FKdKUSiwsoyHA4NV6GQ4J9pcRXVl0cPQOz+Jmp8YJ+OmWLw19pOSwhCL5NFdB0SP
5NlI90/V+YYYokJFTNRQDDULuh5HMBQRMgFuTVf5GMPlQQkh9vYrmb6b0QsNKbJ3
TkLEyVuCFs/EoKEI72B5iaLDiZYT7jUDArIuyJoRF6l3ELrh8x8aXYWoXxCq686p
rYV3gmAxifgKDCsoF2vBwXGKgNGaO+V9Z1KtGBlu2fKtQHvpqD02K4jOtToJyUdc
iP0UB/EapbQxqmeTVgyUTSEPmbvDnuSxPnPW/9xOsJI057c2RD8pLkVDGdzmdLKx
SSFGrfZiGJ5zYUq1jTIDxaFFJrjsaiDP2FmLyPStNSxGF9yrm+8iQai+nwN59kD1
XuwARoVrLlS6aHhK2D1/CCutwZPxmS59/VND9j2J39mqTlPqtL2NAhXhhUwucYc7
SkVsTEZcaz4KRfU7YEX+7+4DYHHLYJaP8vLluwkD/+McholQOkZs377qbtQtFx9D
/i3UQzjdCWxQ68tc9PXVL6rVN5BaISUg/av6nUrl95H7XCk0GUYusSLaJOeWf6yc
6spnl/UVoTVk1ng7OvmeLaOIEGxQTA50ct3cCjhs178INsRvWFS9QOXuo4cboeGE
MAbApikvFnNDNIicWwQppdW3ZEruRccHnPTtC3It+Z5XMDNebY/kimWaK4GAh/Br
iB4EfkXZ9SLn110y7EMddM+Qq+UKGIo+fAg84SmNsaXFyMUJbqdepI6PmVUZWrLH
eBUEqDm3Tcp00R7rl8XsNJrG67tzZOPucCqYWYx512rsxDc/I+ACJDlObPB5+pqT
UdTBasSf2BNHigMwW+WZSrrBZYqFvik8N1SXZq4+hS3Gw9Ga26Qr7LASuh+ANroV
67bCwde+iHNbFWT15P/fw+DZiFCLb4JBMyfpEG/YQ4OQTelLQpHkavaRv8xGYiFS
BhgqvkkfD7JtgrnH7RDuy9gTwonulE9ZsTN6gseHr0TQ81Yu7RFrGu9ZOqPhFeJR
auhq1HbDdBwnnWgFLgfhSYv6oQvrO3apEH33Gs8lX8dn1GTHGf77RzkL0pCLnHtp
8CYJE9TIBhl+V2k6mO6W6srihl8PmvLCysNHPdLonZOhxUO87+TMucWc9pCYNO5B
yrqOAgDIfHYxNkmps7f94YszGL2fgjt7oQdskQOG4rLxG7q9U1Aq/V57M5tnILkU
2OfIbKlUvBwLgN5Tij+t+gRp7SWe25b2TjaIyeGrW3JrC1AfBFQoLni5gNk2LH7b
oWsN3BIgntaRSquSmmpl/+WTAAogZrnNbLR8KbqFrGMwL9EoLTCXg32nqqNJtKie
FfmypOw9w1LRvbp/7BmIonaeRQp0YNAuFImVTgBepbrHKR/294nHPbzcWb4HZAHu
kMPwo8j/oG8MRxQVsvHbhSv8oLLPKVPipd7WnuHpYDKZkxa7MhiSE0kKmVSBAkGn
j3Uqm6LLDGLRpP5swDcD3oLn+UbEmRHXQvybDfDt2nP1GjT9sK14HetZmESQrE1s
6CXpCFKVUfGaxD+ydSEmBRdw17WWIatccLuth8OX2s0rZI+tBwaImY/28BCPn5bQ
OdzHy1NUtyQ8yF+av08xb/TKLHX7ajSCxdEzHWi3zH/+C/aqjobyxuJUlwCy2wzM
QBEi3C+88MR+EyHVjKRx5KjD0eKfXnBi0Cvjhqbb/XekkPCQjfuuLVy+FA8SZl0D
d2vT3HEu488576KbcclVkcFDOzwy/xb1arWuEzpE1NvkHS/LX/t9EqotWgbeX4OX
rllStZX3FXKZqy7EfL/qSw1GOaxmbpryGlXt7/aJBSBdlotHSWX8n57tWHRHx5S/
/4xL7CR16Un4ku3NYrqCWIIMp3aYyM80/rkBBp04xVoa7HQFiep68PkXlHFwjtqK
mgRt/uqJ7ulnI7dphSzQR4ncnv0INyQYm7YMhi/xoovfiSFfOm0Op4Kl6w1Icpxm
jC0X5TBwjVuydkDgB0t1z3+JVF4F7iIdG7zwVmYS0khaTe6fR6tp/OGkoqJlAe67
tfWRAB3Blv+EjmbTSs9q2onUiaMsMRFkSrYnvk7uVkkrHIQpAlBRJCkSDVxW8Ued
tebEz5FJ0TGz6G3nHaACykcT1lEoqWW/lLdN+XVlprrqCmbdu7vnJ/+BSpJjJ9Vp
70OzltIn4ldaPEQ/CeafjPU3k622H2U0KjgEYvysBczpdr9xIngkfTPJlKONb5lo
e/PFCw3hjyyDdMr+XJ+RsVADeVyCTrNnIA/tAhzC7cgZ6g3DhigGR3oFKJcB7TJ0
8QKkEl4w9oXZs49x+jraF0lNBknAR9baL7LpibZ7nrIDI8BkG1cV4Qoy+YIIQljb
rfWwSfSJbDi8JtfollAxVz0DEmtif2+3uGADSuybDKETm5HMziJXQr6qtc1dMViP
QlP6CRK1Q8rF5NPOro51w0rYRiLlAtltLIdLYsEcb4/0iEz9B6q0j+bDtV1o8e1U
mDhGgUJddBYFAEJLy6MA6oqvBJvwM5J9wF0df7s7UghKJi4bT5b5Fszs0oO9d/mJ
7+8dIHtSbLUeXDgjZWXgPIpBFR7yb4bw9gsrzYmBRh5l0eBbGL3vTBjL2pYWQToQ
N9MqMBaIIHrSUqZ8dbaHxSLQ0HJvgLyZaQa+qzopFxwILt/oQpS33V+YrrNoijuN
8CyIGhlwhVhH9AYne9yuyHMmpMixCOJnV18DgV4hwe1vS3DOy3n0Q+97kdtOlaMp
qH6c1rzXjLPepzXtw77j3tJ7JoVtu20r4N/jO/hIVM7Aau+Q2+bbgUPngu0gK8BK
ANrVKdgipRO4+gtuMNvcHlu2COsE0B6fzJgir2tG3dNWRDTqdAwhmO2cgoRuJgtk
R6SUzfV3B5H88oMaSzFTo3BelE2aKOIKXYc/ccwmlndBuwrRGUVBaKp+fMK70Q/Z
rBy8GI3mmVyVLUbhFK1sk/DR3Exn8RQvparc1ZcjQvjR/D5Swgn7zsqk3iIy0zXH
Q2/OFqdoiJ8Z96NqXy88DZ/PyeKXlhRMPo9/RIlFkyVHb/Ls5vxCx+dNH862fRTH
clP+Kf0cgBl2o7g1qevPqdbJnxQXkQqkjIjHYoECS3U8xHX+KHGe1tjbdX5PU1JS
JGNVRN5UstCl9BhF8Go6ERzRCDXBKCNOGWfLznnbb3ts54GT59zC7cR/2X+daP4y
+f+XCgwEKjO/JK89HW0SgluYj13XyMP7VlCgecDrDrcmqQzniNjD4jGLb837Q93c
mmDBxWHwJ0AVLuRe/xXPu0z+labm519uiSY4pxKo1PHA7nXnQd7v/YOmIeb/50dP
/eWCC4HJM7EDNWVW6rfoD9Sn/tLPhoInHQr1XrHWIIJKl/E+Wme1gkvTS/vSjff9
NmRlhSsEyWWA3687LqUmMbSbC3O7Il0DQJBVANkRqlErH+5Ev4RDXvLiUqA8iP1p
5nlCu9fa3zBN5tZCdyw/B7c1+nMZtxtUbis0crkvXqBLA0B1oXtvgkgPVr32GFhe
USY+nTqQVGPMtmu71k1G/AkzmleyibLg1t7OnGHR9+jTray+NgXn3g1G92EIaLPQ
/w+4XHGLEVTZlU3eXujHjVf7GmyJbOrpRCQ7EbAZ2GnduMFowe4ZGWrj0M+yFbCL
jaxLQlEXrHCpo07/Yfym3Hmz5qs8XI9k3y9I7R7Y7iwo5zgWR8luzAYWI3LCnCZk
vD02O6N5Mw4BC4t6b8cRJ942PVGGdUO8NJmfALPhG++lYb+3Aakd8qlSuFKFG0Op
4rRgKaDaz505Zx/yKAgvSy96mNZkUpKKwOqIQIQrZmxRzvydZ1j3tUkhSkdDRlrm
2lNwRl4MD3EXpI/IJZitDUTKeyvX86nx7dQx01NE6E2MEdQ75+0lJ7a+hNGmsgp6
a93XS1KR0c5nYq9saIloeGepOn6Bsri1GpPlsA03pfQLIdl/3MxItFdOGuXYomJ0
gW7aD9cCGY/Egl80hjya8iR+/gQAHfVW1jvVTSe8sq6HAufnWm/Erjb7qBZ78umG
MS4p9Dx8JbGcyE3BpcnLFrqk3XSoB3lO5hCFmzS2ELPXn8EpCUSvCTDaIT+ZxgFF
EvmLIm6vzGcSD5dTq4LYiP6tRKGWcVWxF0QCWmSX1L/LS/PYiVpL2E2xO2Hl8dB3
9QB9pPIUBLcB9q7d95nlIGoK4optWP6Aad4voAvjADXXsbNSQwrkwmTQoXhRF1Lj
F4hMe6uAPn3V54juNUudqI4WwcCLIu8ohDvvodFlOcyLIHRjPqkOZBBjRJ74e0gW
ek0kaxc0f1FRpmcCrqesI23DfLZeZA6w2+v58U1dHSOjXaT1nk8x81s8pLPXJ2PV
lu/f5DhjeB5wrt5Q2ciPgjW1U1gECC6gx84M/TtmLZLalyzs3IqhU8917OJq3h7y
c0iFdevKWZmXvqUDRapqKxF9jZRPLyhHzPovZWJRyzRX2UMNXpzMI0LF0P+SFXHz
dionEqJ0PbZBhmXv0SKM+Qrb3T9oxgwZDJ6ziB5lWpvzdLUGYNhs3gw9kWL+px8G
c3OFXw2NNovGoMYSNLWwDTDi4AXZQm3a7tIbey1mNPtAXltSjc4nkLYpeLotPPeZ
U484f69Ef631dA4by68hSvdvs5PE4Fj8z/i73VNdkpJ/exUvJuTg+O7H+84cYf2A
wbRawib+k3U/V+VE+nm99Hy4ZKOJO2myxyX8kQ5QhFxanMGik9MxqKr7dq0IOccv
UHFvouoCg2UsUi+Te1KgORfWw/cawTnq1Z+zpuhBGl7O2huhsMD1X8iUNg/pAAnh
6aBlLfCuTpDXqJcNBjj99s9lOwtt0+EkHaQ4sB6aAIl9B/hOjEx/GFp3PVp5Fz0d
DmG3jbRWKn09lt7JspxZV7HHxGaTLA+f3insTfnEOoMtzagtW+b+cVj4MFhXNcYu
wnyd30a/kM5ZD8jaMEfJ9AMyQy0suFhlLmy2mhe2KMpX1Jc84qW/xQoMb1aifT1f
EB7HnuJLvMapoNbVlcs2ihuug2DeRccVw9znj0c1GGNNmbawUoOBv9NFWrGXWL2F
yQ/bOfeLBonXf9Qv6oZgy53eFACNjwyuOZUF/ft+jLttle/m5kT1jgQNOAe0+UkJ
pyswI8MJ4hnifcEV8g4ec5YvJGvqxUh93b3MqmINolyKWsd8kg1c2leM+j9RAQ39
9dyrN9O7dK4ejzhGAPBx4JDq4W9NLabVTEaKkntdKze1ulTIxizPXZ1CyFJ0xR6A
cR2b2e1GFt1+5II/5X2maqUQaGtQ0ESf2VPAOTvyRnCLNDMCcKKUOk88mgZ2MOFV
qiXhLJK9KfizRMoxfRc0jmEd0QKi21R+Sv7Ys/ylVEzX+SAQCkVjqg84H7o2hpEJ
5UaowAG6CPxbvnCNeQMhRIJRUoML4ZKvkojHH/Zf6C1I0ovCtbpN6ypwb5SQ/DoL
KQNygljAQk8PfpmUnMbqT1KRedzljo3exSKIiL+8r1PLWF1mfC91d6PX+hIs70CA
KuPHCtgAc8blLd/nDjvLcTPUSkweUVJxiE/GHxQ2f5K5izv8PWkjHt6RI98+MLsI
C2KFUct7VeZ+N5Gom9tJNUz/AZD+Ov5ANhxhbHNCLNpp02IBInNCqbb6rdyUg/US
EgGP/c1I6SGYWaCtz1uqCtSmpldCcsO1z/KipRroeoBLsG7IYRwXlceEQJuoRWD+
`protect END_PROTECTED
