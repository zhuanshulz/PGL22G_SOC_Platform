`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DLmoeyu5KiScC7Hv0A574IpC4xOulEOpR1jJXmhwUeoYiE3szWzILJyqjr/qin6d
ynorkuJ5ebImW3hjAoxOxBEOT/KHEdxM2uNMLhojcab619R68WUb7zxfGSpc/C7o
s78x9aS6r9PKGQzkUXC6RwhCMh+1BBf+LX3RPqGuyb+2Y30o5nQV0+71Aj668Cb2
REf+oaWknPOsIHOm21QKkp4rLYycRrrVj4d6Gp7mJStyyK/HPSamYUGPdIQ+llNH
h51tHKA42H6wQ5UDp7M8xwVJHKemY9AYnMppelK+K2bKrkKHEiQ35ndt1MeEDdt5
+3aiFasq8bFkn1pNsurBPsxP0H79Hzqm3Aa1AgWs3UHtgwLAJLJ7domOya4n4/3M
UrecTo4eb4iUS43JXSl5dr68CMl7T/Sdz0wIXXH4h4Jqg15PQPfPbjThAwJSqHeJ
D+Liw98OUnvssBh6SY1XzHSVOJ1cb7t3jnrM5Dq91hUZ3SaLnkClslTALhynFppv
dA9nS0OJ7mGKu2hQ3B3qvTiXlS6piBbIIs6FKaD7tDCqKAB3zBNvZpZTdqPIkwYw
KpVA15FEw2b5ZWZ1gBtfIc3qy+Z7FR64MqFsW+i0qeLYxoXXrnyIDBJrdpHqGLls
yGCX/I3sjXz7DSVVxCiAVNzDAUXY/60UTtLea1Yh41u51oXJOoh++mlhVe9Ufh6+
+byNKqK7Rli2mR2b5GQZgRCJZUJTwqFkeTAS5qjxN8HicTDa1inDfoxoJSFt4aNy
S1qKSWEdvpvSKJW7m1SNnexpCRcS8huMBbAUw/2+rmaJAxZeCJTCg4wt24jhbdsa
1rCz3zTEktZxgg9h+zfSTqkbCQCUIJuvKcD4cPfirmPKUvedg0nvie13WlXbJ9Ah
b+Wh3emoRSu8iu7hYoo07A==
`protect END_PROTECTED
