`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KVt+uciLueiDP6d5CPrvezjZEEo26E5p+6Ek/yIoXkkVJxN+HZIFBj5ZkezN8nR4
LGhDn/luywArieVgiOFrkcKmqlUaTJR1pIEckCplc3zazNOlljoNnc3XJvCRTMEx
4u6di1YNNa+3FUMZ4yXFQ8kR9G0zHTuz4pgg6dQZjRHw5YWpdZ0tfmZx3RBinamW
8uRLX6hUVfgJiLzuBASIRNeSjGGCk+ZfvMBXluzjXo7Wledbi8/yoPMHSbDK4L1X
14kRr1DrpfOkUbUH4hwQVWZh1E4AEispQMbreHWt6E+w0vhRN6NJbw0lzlNdo9Bw
aTj9Ami8/lR3Jt2NOah0YOizVbLETdG+IDXpxYIV6orHE32W9ESzL7SSJp089Whb
+VCuNhX5z2NPhmLwhhYWT9unn4GHT6k0bWIGyWXQDroXSGJpeErfoYAnTgMVw3nx
giMGC2mADjVu0Ny9gaCTi2IPUpQYJY9BrZjH9/a77wWScWcMiIIlkkReSBui3MAs
bJwZ5UZqRx2Tk+/djOBZp4cJu+S9afH4v3EPI2xMh4aqGMyvIxnJ80ySjhGVxcBR
euX7H0+L5OE9ZQd00QRC+zEJSaIyqv5f78RzZk1A8C3fEl8WtKnFXxYVpC/BQUxx
9PshprBOAzVhFvj1chj6r5s0i6NvD9gNJYJE1/KlYdr/n/vej/VMktu9+GkQBXwL
SpfC81H/38qqSyR6eONhcHpllxjYvGoa549465u1qwkUfD0FwhgTmTBUVznP7sCR
daWIILQVRP29RJwkOiXdRvZexvBRDa+ObTbysRVoA5WC1Q3Lk3SOUE8fhbUQIgGS
6Qa9+lBrnGrJ6VttscHAVEWWvh+Wdf563njJ6hrba2E65gpad8dYmrdCe2ih1qul
8mm77Z0j9Hu/XzDhLm5aUPqKo5LCv0zJqq9nraZs5GYi/dkT/hQQoFB3BNWEEq9X
76szcZw2I2w9xZqAx9gy4ACVAm9gtrgDeI8r3MHS2zg4wHCrcqwTAapCM/O1GTst
SDxC0QBiQh9vDUZUHFkVlJKRofRQ2MhlcYY7iGNamn5KQ2zE+bnyx4lfrV+AFLlV
i3MplC8f0rkP7MsKLi37VvoKoSD8iYGYaSLXs3gJc1FkX7cQ1aqxMJ2BwRa4VnHY
xS7RDMUZYEBmWtNZSQ1n8PhhXDh406km4aVnyWvEB8cps56qF5lYytbZsKH5e5bb
9rB41dsvjdY04RQuO/UbOG+dFbgLrrLBAGw9OzWF+OucYjieVnZFpILHthKWxI2o
Qx6te8d24RBNo8ejARYVMZv001F+CFGxOjVnG/pTesEJFbKFNprcTeHHeYBoBSyr
hmPquqSl8/BRkfLbgVUvMFbiQYJaoez0DdwaJCLEE+H5qi/hT4C7yqXyH0JaXLNj
R6ku6nSvFlvvobSiC6tSbyf18ToPSNi/TuFSCUtt7dwLE4ovuFI1uZCdJ+o6InIE
vbRALhS8lQUWoPa3O1a8Miu5kUCeBQ2vESIl4FJ0Ot4aIqnbES5q+MGpdRWKunqT
mRPglcrPgh1qTrBekDFQlj6/9BGwu9VNYdD+R9KxYqz5jde65PnIC+Dbp+TwMrnT
b2XVJcQJlXuNkdRrlQQCcfO64rpmO1jbBsUS+zjNf1DSB7SNQOMDzcWL59rXO8jN
OV8HOOQ3yp1Uj3tRJ3qaT7IGf1PJRrE8f+MKr3uUREO4X0GZ8mfuXtN+jLtUXhwR
cU8NOLh+bS0UOc3Rh1V9HhvlAj5W5JJjsYGsV7FY0lNyF545/A/6em52mRuzAJBt
GHwIYNbc7BDshdZyqsirs/WJ5Oi4AfSxjmYSEUP+3HLXTzlyFMAjZi4vHzHE4FPM
RUbdie40yE++Wv+FkUYnmYGWXFaApPVqW7d2nWAJJxFcbvbR/a5VDuwHgZh6ACB7
8kZDicDbOPoCbtXPh/W3tnUnS1w+AmADPWWNqHGExeAbHFqOPKLUYxt5NGR63Tpv
g7QgyLhF+uj7hvjjxfQO5F2uOTfBTp4dJY6jtcLaURZyxgshlp4PTm/2cdDmT3Gt
Q0EGJDDYP3lNYa43DJSoaTCV/ko9sBtII4JR6NysuX5SajtY51rONGig/goEerMT
8ywPZaJEsKXCaBRG+CkzUyt7g4m63zZFPMHbiRiw27CZYYEW5EuFx3v99g3Tl/xi
1Qa9X4sdfpDAlbkHOSZg4rrHQI+0dt+XExaptTiUf4M8TjNpT990KDmcegVNPo7b
4LT4SKI2jX9b/E/6p/9C0iyeyFPKmW8FI1JtYHjU1QTCFORFNyXhAKdiMmvTW7jh
UP+M9U9JhV0tW+br71YvbApiMuubf+qPBZB4iZLkBQrKGRskcBPeQ7wDymqPvqEr
nbtOBYfSh22p/PgGxwtXutGbaMYoBV8BDEIaJRnj1QnkM13r0zLxvrBVas7Z6ANi
b/lxvv7D8kXP1TQ44oim+/xvmvBiw5oB8A3T9dpiCXFo/hy17DLfCiYbQEF4WkOL
tci8g8ymEClFFctqvzRTUR3nFQ24b1ferGuRi3vqXKsU4QL5uYI3RCqP9/2cgXgL
5JYssSXtSZgph55CMwmR9aAxdobIq0EUWvprjTXuP5J6YyjrY9ES2y5ZEe4gCR/M
PE9eFF4XFGS9++Mt9BvoUS1OyViSYBtZxLqZmgtWn8Jb5W+9n3yK/c4/X6WTTKmd
Yk+mS5+pz/Dj60HqbAf6lN+JT87KJrgYmF9SKdiDt/sTvrO6wYe0TPqp99+S5DE4
pBVF1eDt9E9HqdRf3vhnr/pr52iOAFoWAUr8FJzrJ5BVmq7aF18gUDY0tHLVj/O1
2tc9TcbZz/co4wvoplOq7O5lPSrT73t6nCmMMzLWA83rqHmppDGKv6IH7JH0N4n9
`protect END_PROTECTED
