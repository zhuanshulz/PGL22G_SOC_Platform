`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8HffOxJUkCgfaUqFQLEWPZKfjdElI1ckwz+7rggnFfiTBM8NVcPlsn8yG0a5jlBY
FxJ80ErQfEOlnnG6u6Lcha4ct7fr9hit649OfcLlLQ1faJQ+oHITEDDAqQ4ssTUE
U6qvA3EeyTckkgyvmCGetrm0AaDkiuw+efeFV6aw23Qu4M+o/73/+jVGgUy1rKCu
2GOQdMF6t/ZngqonBfSlHGAvM+IoH46M9RTu98FKC9owCekvHIZ1UIPoZu2REm8A
a6LH1V/ksJrxq2Lo/s+pot4w5XAIA2J68scAuSAEDutkBbbnh2M4YgDwzO1Ds8fS
ROsN5IzNs+Wt8vTOyNICSDyfLCSjfnjOvg5dSmY2UgMPgHQBslZv1g6DQt5ppAT0
5MAIvDbtk1FgNb6p77j1IAd6ht59W/oxoIbVS2ai7GkyXuayO/fz4j1hyyAF8alR
98fKqwfLZSHwh0VL1JaT52vTOZ/oS8IWNrN/YIhYclBMqnEUwI6dnyvxcwVWIHXb
4e00DHMRRhWBjmbKLy4043hwPglHGSfyyo3cYNXOyA0UZnRfi7XRhChe6+BQvn9I
n1zP6Zr88GT8e3OQmuKisvx08h9oDMuv3EClyXr7oPvG7U/FJpr0Wm+8c08sCl5U
kBdv1pJrJPKsTswPVCfFP2JGVFYi/VvCZpb7HEZD7dPDDzdVcgxhJ3dMyd+fgCpG
zJPr+7FjWf/KbJrxDGSm01AKUBn/YnpWqj9ED2ivS5pIVBTTc6Wm5BfiD16fVDIk
8iddHAkVXuNLnX0cD5mjVk1OF89PdC3PkGLlnSCPAOUFlcS0+KvvXiYdS8xrqEOX
t4+wHB4eHi8uy/oFgQ3KXUNCzVC28r21K9xLDkbKWrkZ0ecZlwhqOjZDUt75LwaA
hbna2vSLW03NnrDOhGKdkhBJK4vL/sLy9f03wKyZpp9WLSmVb/CSqayHVf/QGyON
o+r8MFUxnIBV28//pWdOtsInmqv95c72Os8Sdr/UJQOGk4TyOXfqQPI8hSoA2hat
ar1Tlyhn2zlfo1w2vVZEJafQUrzBDcU4zqqrM6WobaKsBw/ZSbdWi9Nj10XDMotH
ZzgiJJHOlomP5aWSkXys8j+kLc1+Ng3S/doskJjbu0VFqXNjMZ181+reHWBTjq3j
8MGNiF6R6un+9BAqSs2j5Yd0QMwAakCXHr24nrXesa2RmzvEqRrSzeMt1URBQ8/H
psHA85Nau4FUOY0TFZncV7Bki2L4Eh9I2cOdbPedISqLhiKzUQJOgc/PjqFvthtB
7hkuuBUncOl1zMjgaYRWGq5UEYQwgSRPuJMo1vU9jrz2Bf2jjKBLHOUzterWsmC3
NbVCkbli/izr9p/GxCGYhd1edw09nTSbVkunzYhzQzSnf5omHKhqpbM4EBNGyNKO
fRfAT6mB+kF0op8P/CBneA==
`protect END_PROTECTED
