`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
of6c3GyCmQk1yKjhPQpHtyDjTpSPDO4W21hNVXs9gjPOsd9P4syOkjiBoM+8ujMU
t/yMMjl9j+voSccvLxuGivZgOSwNlJE2ds3gyYM2nVYhb78DBm16tVPEC9VEM7n5
rq5s8HWpig9kj5PKMnoBs6GZVH5s+RmKFArsdJ7wArQ3Gz30RZuw+FBvm9IfgtkN
fOfcUfvu4KNCPKiTpg9Xc8Ounbs+PZMVDg3zvYXtRiqCz188O/fPqBIYvBTd9ByH
QbDlIZ/5i6LziSnFi1jLTc1m5E53Cun73fIVWwSQOrejQuMf9x7luvGL/nA8yM6a
eUFRaQOq3GdPx+S9wTvOuK0ioS6ajOrnjfyMKF28pyh4j/odR5oGgQzQzkwYBoo9
9jmSsqm395IgsM8T+2VQUAaTwcXzB64qXi6gbR1fGUEZmUZzFU0ZPG+2gN/eesTO
O4qPpjBr5/+riKfZVWWKBZUmYC6ho0b0UltFwSvIkn8eI5efG4NS+h9LjBiYUcZ6
4Li80teAXH3M2aA9lt4Ik0mr/i+q8WhUhtuzLUcXm+CajjeoS+63ugwPKZXIQFCA
OEZhhDeP71DBXYAmOlRDq9q6xSmL7bG6tDBPRCwXqfRnlpB+N5c+czLsXGOaBN4E
RZNf3xQkGdEi43/alYNYvPDOB7wCGtRkX1crTTLV8WDEy+h+e8QUqcGDyzPicyjJ
Y1SqFqa8MAfUNFcTYjrIoxTNv5KBbGAvDrWOwYBWo4yUypeCobPAVWGHX2uWbfWU
pLyKb88OJoZaSOFoQ9QLcG36ZaZV+tBZqPYX6kPefGphVEh4TgP2gnmL2rK3UZN6
W2uJoxON4R+qrc5tym4vpv3OnT2jBzDNRKhRU8UKRBrAe+z3IVdDdviJqozoFyXC
xQygvk8eMA19rAHQK9cK/Ss/qUYp229Ef1tj+Kc8i6MF6DE6ryiabD7zx9bzAF6r
3lZW16MWJtErBU9mK+MZv1qaUe5OsxPJWgVkpj5ovvFmhOpiEAbxD+fV0HXZMfQu
9Wsoqb/Hw0Tmf/nFZvXp8U0+E/23qYDE/vsT0B8enhjteH8i81cHcrgmeRhOEV1b
BUxVkauxpEssAq1IEqycK4Kw7BqC1V0uZ5tczvuakjKcHJr5u9grEtKCdNC3zCAj
pUnuSz7BN/9MOC6nbhzq9VSkQHCVWjaPeZPtk6BWK890b6Aw2kKFR75y6LJYEMiP
9W/eQ4dMZuwIzG3msDTPXJA9EJyF+Tjr9GUlFuL7YqjizZ3OTUzbMJuk/xky+pSi
IiK9LEmhmLZu0W27ixaJDWEYeXdZQAnjszYipsPm64ygiSfiMlEPGRZ/MxymxyuE
R1KBgJsr4Bs7yJjxOJDYADwTFr/6dyAEo9Gy42qMk/tk/B13mPW124QnI4uycCNT
1aGJm4QPkdeJWkXlOnGvzYlA5w4tSnHMRTJAgx43GCqttZjbFFae1tupt5LkQtZL
j+C6EYr6MN+btfulOZulhOi6/BUHhTkzbzIMOe+ChCDVaKDXsMi+gh14H6QnR0hM
aGHUaGNLI2msBYA8Q+DSYTtUU9nHPvvkOFOrY73ooj+p14txKgshNLDO1Zju2lca
+bDZ0DH8PDAF/MfwuIRNfTLaVIgvyaUP863QAFxENoJvIy/ruh9xYhvmmAcA7uiz
DPGLsJLEhPnsBc+2lI+dPzW0tIvOVHLMJ88P0JL8pUAjAHu7APK14sjxCM7A6UIi
S2dkavhsaQxa6FneFXwGQHVJ0srj1EKt3AMbS2U5gXIPxjy4B+x4c4ZNsHwRDjuC
b8y3Wit6D74GKh04m7HgozCRL2Aw8Zd2KJMVrEI7yS8WgrZXOVmdtisK3lASoPE4
sbDSGEhPJJ0y6ICJnmZ/NBtw2WksjkC7ZelG6rKzzwa6M+dswOMZ0mpifdjVhvPC
wEebjqmaTGZaOqpb5LwP1g+bHP5QoOhWU3CBbtdYTHUVUukap9X08IB/yf+XgGP9
TkRZlMFPjXcVWvOjGGNCMlA76rrypkHW32v5F0BlN1I7iNTL4Cf6rKv6JEPwYhB7
BAxNsfZ1rNWKJTqyUFitU+Es4VyX7/ZJp/MLTHsmRDMypKdu/kddEpgbceRSGs0u
sF+RBYx5BL21y3lcTMfZ8Gq/RxXvIDPLMUXpK46dLZGCQoCG1t6ttHMBJn8Umn2O
iP8NRaAVZ2QgS9wVMN6kYmGb+lrpWBwpcnjG0kHWfZm/2WIiM1/bJ1HiROLbcGQv
1EqWSFxW48HJjKbOmlIJaXN2CQrtvZy8ZpcpOwFj1VOIL7nYn9UwT0ZWIc+dAxrV
1HPzSaCVI5Jioll3RgfBEGvJGaSfwXvUJh6NNE6AoF3e8Ku9lZCIIVinu3hJt1Wn
V9RPX+vTpVRXvFDDTAiDXEon0DudVyHOB5OsP/WPgTokO2IasxYcfYtHYbuqWWsL
raRGuFQ9AC4/Hm2lEqinSdbVFKOzLMpLWvXY08hmUYp5y+zoCyOK6du5wQ1OS8er
zuxirn/GV+pK8Bb/o1zrqWYmVYvNGAwENvIzge76vx2bGEMkfc1RWf3CBKM8dEIO
WsYCeV27KmXfN0/V4GfR1w==
`protect END_PROTECTED
