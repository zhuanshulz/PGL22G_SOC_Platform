`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+QLDT0hdpNpexFfXgeKjZ9TJ07zv55uSBuyM5rlPrUvV+dw3yGW43qtBg356BqLB
Maxjc6YLzMaP8X8svDPGAZM/C4VC+MTPutgvRVdObrl+VIHjEuN9l8CB/pIEUWuY
3XIEnu2E5IAeKQ2j4wN+/Oq4mxDbhLKFYX2NK62l1S9JgCyowpj2EO5rPWcOH0n8
uWS5E+6EqGLY3JrXcn87Jh8nN/VFB4RNOpE1w4ANuWtKZYF5b4vDjC5Q0gCnWiAh
Trdmrl77uCUVUlVSDZ5MqC7N4apu3BanhvH4FHFq0nAlH1xO8H6Go6wK7B6lhRzJ
AZOtcuIcmDX6djOo/5bdXd4dDNf8zVdAK0N0NN018DAuvosNlOwd6psWgNEBmHz1
34lEYTSqYfWQk5JL1RgTIe0MAjU/APjyA0YNMm2a8UeY3eoP36yfsEPZP29EgkPC
kyTiqjjK2j6H0PyS3OF9+rQobHfGxGd9KAh51gF02nhi0HN+FmyM4EDr4gFlCAFf
VpzqnpuGS8PZLauFR2VALS2k/XWJQATfIp6W2IYrQHSZql1sblZoeBBrHJsc6h05
AAbdnqamhjmwT5NqkAfGjzNL0ZFBOcUlqByiluXNALV2jCPrkIZksZiarb61DmC/
UDOWSiFP5RL8eUdSfPARuT84/VTCiBq3z9U94Z9wq2O9ftB2XW+GcBjmDg7LoVcf
DR29sTTNElZuATNBYeyG+EWCrEwn3020TyVfh6BnHGoVSdD3mgDyl7n7N5rNl4HC
6Rmq8WTS1oWa56Nup2Ngi2KWGiNNv6tkgUN0rrUZpvXNF2VDgb3R97PWcS+DcnPv
xd0GrVPA8Nl0asWD6D5Biif599bKrsBMYV1IDPcmh0pwesQajYMNzuFWC+Lh3Q+6
FPnk+AFFlOS13tIS111eauEVCFr5xiq6HhGwzAqKeahvlfH1EaMZOIQbhr55PVuR
9OFEUovCzlPhB1MQTQfOSecbabXXl3MofLhDqOkYso5o3vchjX5oYWzTg4GggpDM
zpL0B2Pjzt0iUwlztMLfKecHQkXfplDJ8TSagMsEEVzqoG1auT2IhVWh0E/1NHPk
mvHumrcoH2FC8M097f2qqZLQO1zU1rpPRNY8JvqYbtJw2jnCh45M8E41PWsShRck
yCCkvnHe6i83bTOzpmEJtp+LS6BWgAHbH1BzBhtiRJFVdESp63VsS6sb206sUB3O
/FL7TWhLyYNtX+dG67NciLQS/UVBKS1nClXJ6NV8Qti+MRoihmoYL0OQ0Ts94HxK
uxyzc392qyAfWfk98l3ylso2UhmDhk3x0sW3sACT/NzTh4lc1Uwye/cY0l7Q2YGu
aDdvvRxgo3tpcDRYXTahbGteJbiK6sf/yQk0WP0+k7nLssMu5omBPx87W6Nk29It
O3IGAh/yVd6mb9r8tyTL9bTi5uuQK+uOei81RE3EBq5qib3+hYrJsM4ksz/q7T4Q
aWP9/bvOdOQG6Hla32FkmT+r3Zw0yR/E61jIPOW+DsL5eW1JMSHM8oIb36534uuE
xEjE87Gqds5YNZMuYzA/q9/M5bwvMZdFJbpUQ+I9ytpxhuhWrHzVcOwjGSdFJzhZ
8A9YahGx86DjiL0zRgOMYSJEF7xggKOxfh/oQcSnR8AUDTdQ0zIh1VnGxu7RrV9n
y+fd4Nsq+AF8z+05wGMABuktR1qtj39y2y1mDXDa+R81mEBQWoyP2rpeX3ckGP5Q
LSiTMxHAGYn/QjUqwXrvlO5L8G7VnPpLFA5pYBZrQKL4Zi3R0l/lSAKefFTlrnGV
nt8oB7PFIaI5wWA8sx2tj6dS0d1HBJNsF/ApFFTTTs4zx2+va4GNT27dIinG8Rm5
T2SSBblw3+j4wSMlFc/xykbaOn2NEff294LhkE+cKa8d0PZI0s02l14cPKuaa9f3
3ZMGFq/jFC8bBgn2yXrZVRWHGSELQV7+qhHu0/SSCic=
`protect END_PROTECTED
