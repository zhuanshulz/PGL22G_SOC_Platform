`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XKk0oUufrLIIq3J36nTdVRRXydZI7hza6uJbS6p2h276MAMIB1BCvMQ7+wXN4h2q
MjglBm6qpwASE4csxk9tP0+n2MX42GZ2GmqHydqWFoG1QpKap76e59StM+buAZMk
XXVq7oyawUNfEBwYkChegxWcx6gmjae6eM+XMGF7+mnktpVQs1335Fa7BDtCh1gq
t/s/IkbpiCHElJ8MYOqZH+fRY4+ZUj89lHJZimp1+vlZ1EqjK92m2TJKRjUkjI8d
rFFULl10v1riggwbYfib6RldPbtTOiSBzmMSzss5Y1kdtqo6c5CCjzYbtwNjuwQ2
UYcpXTqrgn+1vnQYpVYspuar4D6ndJeo8TXb2vk8H3tEfweL0xmCAguwS8TpRsaq
1SinWSb0Mljeoxm74CwJfphoL85U6f/eqoB3ZDERbXprQkSYqryVEsTa5JpoJwFt
nDCtzmwqG4gy2QyB0cYoYw==
`protect END_PROTECTED
