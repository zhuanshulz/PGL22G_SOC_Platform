`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u5Iri5iCFB5ikj92fWnmYFujAdFeKmzYANr5C2jxVO/yRBjImrv281ZuGs+OdK19
1XJf/hbnRMZ5JDsfqj9r2xIuycQn3yNDtOWVYau+aRa7p02pQGXKLY44qRoH22MR
CGW1zvkLzYkm8FhnUvoSx8XY/5mTNTH3feIHBzgkH1Sd+NE9ZYkHyk/cjDCtvDju
sDaHYGQaAPjIvE3jYVytn1iCqb0k9Mrwr4GTM/Uqx91oktBBCspdfXQeScyjjBWk
X3fyPQ0yXdp1xvSS4ptNZo1EHSr5jJBKkiT/WlAdRHvNYv+zCC08CH/ncXkamGAF
fJcjKeLYDKwcZKkSIe8ZQtlmrbsaEyl4oy7YP9WSdzu4NlYy6PQOpwfH9EbLXZAW
sgp8ZrlVaW8r71i8c5rgIeB415FiIYwR7je4loohsTNvhFJiUDMDhZ2NsdvWWxPH
f+bP0aFHxCNzRKKtZpg130YAYNDYwa1quaMgRbU3MN5U8WTOXevimDVjo4ick+u3
VY2fu9eN9B2LNBo8m0D6LMP4ZpWLsMJoSAttLbpPj8rZCPwHj2tVOu6PopZ7+qWa
4kNOWzk9zweiGFXLWXnUzpBfvzc3D55P3OsYF1Lid9X5IwCgrHpKIBUM9R9cevtB
sh+Qas0hsSfK8hK1ZK4v7HbRE5GGNoSOBVA29L0rikIEE0Z99YaAl8xiZYRqD5Ag
lD4Jfk6kAyBUqD5AjL/tLGpjB2PIqMwt+sTH4+f8FIWAjKHVrT089Rpn4Hm6ycUw
9QEeDPRkHA1sFZFp7pR9vIUqbjDpsNUssvwHDuHX/Ynm6OE5HUVoOijaGOqyfok1
LrxqMdc005kNi/xI+qS1G6tQgf8/CR4MlZ4wqgPp1kKMSTqGl/5ZV9FUgaHTNgvv
st89bcZJb3bjc+Qm4m3VyP6+3cwBc9rLMw9r91NWW1TXZ/P34FjC4MCFtESA3vbG
RcUF/ffebthxtpCrCBWb3w==
`protect END_PROTECTED
