`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DUyw+KCDNvW53r9amyLT3eWRkRRyNkh0FCDf2yINRCd2yAKJEjeDI5CmWSxM3NIQ
vsRlz90oknaftE1KX8ebXeWraPm1qbP80chGzR98+QHp8zRHS5gt1v2+p6k1OJvJ
yS3Ybes9zrcNAkeF1ECDdcTVLO/E2SgUDysxDKHnu33sUqFD7Pijlce/xwl5H+jP
fMrALTUZDW78nEsEDvlm6+zRqzyc/FrkdeO3Mim+7ARRpKdIhhW1GOlRECTpnKvN
RytZqOiHvo4DyzooOW03T+a7UwtpviamVQy7BvOfoEc=
`protect END_PROTECTED
