`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EbSPrPipG9eGDS05Dz4CRKTgktxswzQhcQxKPuLJKFnzY3OmaBZWXJUsv6gZ5eCi
qu2/JpFXcTGNACYsI2aRETb5++t0g+mmv0wbRM/8GK+E1X3qdJ9d/Pt4MXfmYSIU
uGqssPMOlXmcvIu9wDY5+mIks7lWhw4330kjj2iFupi4t9SKrr3LdPaPv1ibDUlV
Vw+T6NQhtETVb0kTOH3aJV6uP5uyjbzDEdKG7Bi2g5pdKAS4um9acw9AdbZAJTkO
V8mZgF0pCCO8SwTAdGlEQ+2Ju2ek++Fq/HafNvKL7taB03ACXSeHW8QYkeNF480g
48PxwiLV5AlawgQSf7rSINZGKnP1Z3Q1R9tFU7hp6kQGnOCvByUxJGB/jkmfZ4GN
ThfjuOiwiE3pk037GBWuILcbYAn7qABUIg39qwGLG64oMSzsGRRvIFESDn1TJcxo
dGNZ2wDZyk2sfiwFxh3TMOgkNVHLNSFFKVSr627UCJqz/cFqbYCWUmpeinS8oqGr
COGsMXpK8WwZDs3MDjKeAjnE75Np2BeVBUsgEAdp4MvxbHC1fBFbsM2h1I1JrLGN
sFt1UkTnDnmUU0cAwswq0MBLbIx1SkRNCi/laB3oe0ijAIaf8t3YMzypNB3S7hkq
usdQAhvsB/wo6QqnSJct98CsA9kRq78fAfjuucgozSpoiLT8CAeXX/o7+ZHCuyGH
VCdiD1btcLKVtBJYXxM2IBNoOC9I7jbIxIwD54WUeGbhgVAfA8IpES4OjZ/jVaRk
It4/tWopwTibQCCM/c1glcszpUm5JxNQVl5rY2XIGcb5uCKxSFr448fHl8JDHhsW
n6O+FY6OWbDVJIFUeT7e8+51BNeOM/xeG4DQ59Z+PW20zSbyOKNr8WTSUzq3EvVN
aearJ9eJfBFNQ9txCT6n6QwALwRKfvblMSnxFEAdiBc9ZI4D/FAYWyzYUkcAqH8a
dsBq0UsiM6XjuMn/SEHqdJEzJQO1C08UtW43w5v8cTZ6t/zbuZtfs/0FI+t2Y33f
dGQaJQGz44psvRyaHBLh3Da2rVfx0bhhDk680Ye5p1RycXkAyZOIq1Bqtu7DcJno
7a/L51Hdu+V8j/GxCm49ubagDPGrrlRdb9i3xaVgF1JnQHxcy93eAQEA1GGY9Nrn
Vn8FCWd3mo6YwpSKkcUPEw==
`protect END_PROTECTED
