`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H3wP04lgXNlbJX6m6AYe8LGPdZ6O4+T9E8HQmb7R4VOuj1avOSjabcj3UV8Qajq4
Klx7x6E8qRoPfXq3qkv+L5/gcZNxF1eQQbnbaKJ7lDiXNm5C47uE5TQoWJHUh2xE
o9ewHZ3JjTbYqETEZAqDKouDgGFcglGCF8MPe6VsWVkHqpyver5wO5Nw/7pt52fb
pHXQDsFC0vHKDXDKmElG5xYQX78+Cbm6WGuYZavDWR5Uk6IXp7cnepb+9BJG8DIq
09mfD0iLNeQhCWkCrLlhxGzhZxKkHiMy+0mXYBRE4OBiGah7bCsBmpIqJA76Zml7
7IW8nPdDLSx5VCbODH21OOPb2ExCmhiyrJJTSAnT48M6lG7Mnz89/VexShniz2OL
TY/xSeL1NxLsL0iOmdUWXOVOPIfDlubf3ljGgRGZXNCSs1llAPcRtgk9Hp7IQy3U
WQbjh/gZyXEODL7QHsD5hCknVCs+lPu7KzSer5YLUD94F3nMA53Ox6LM35V586mA
klw6qWcogF5H5Z8UVuQvSNb75SV2WBFxUCd/KSJqEZo9ruOX+6XOO93FPyTlFb0+
4aCJmkxVmlJGQDxncsMonORIP0U7qCG94SNFSpJ4SQBu14GK23JTyeDciwHqFUJh
znq+wgW5ToqfPgFjRX5mxTPYN5kreIYMJwX8FmG/ltABEBSwYHbEq+SyrCleQrMs
zPuDdZmJuWLD9w0AYXmBdZykADpyIk+OZIxzGaLM7/x7a5GQzzJJhs5b/o9lm0DI
oGpSE2FKEsM5KwfwT3h54XWk2cUB4xeToES6lvHhp6QzXDlFDI0wt8pvHNC82n5n
oL6dWJP24cguAlTJ9ne0qOp04covlBY1oTk9GReqWn5fFVvC/YmufAlE7WxRpNEh
fZqPKiktqTVWzwWJ7YzsPh7hQCI1NT4mb2v6I92XLQRmsjDKWLIU5yFT43yowbmD
97nLZLoJBMU9Y6qLy2h//qlwCmSypNdGseeXwpqft4uQE22QX4Rx0yLNjeemAJ5X
WiQhO/4zArcCwrv/VJoouDmACaHq3ffMHRV8vQcsInoyUp9EBWMewIbEV6IKLp2L
gfwH/jqsjak4QWB+V9b6BA8zsq09OcE9hc1lCRlJ1C9zFVSNA9r0EG2OovvSmF7k
UfUj8TrGSi9L44xCo2ja0wi7WcGiohqDH+ztO/brisRtQQtGfZ+z7aRK0ySH1zYm
NNELtU2riZwOVz/UEZilCLxkEiG21WwYuGXUEHAo8N0e5/+t4odOdxR8jgEFyZo0
YDHxAMMPDBP7lxTsr4YikuMLrAzC5NAgZtQ/0gQ6kzk8mkfFlDTqeJIo1+Hn4zTv
efUAwWLjITkUyt1FJQtFUmQ0IeiVBIuBESqOGQy8SbPRw6bUe92Ibo6xw14lcukT
pWAzQYqJpoTOwlhE5VBVNwv2sw9UdYQEz6twh1YQ1cgeLoGnjBpvwojJobcOaMYK
Q18SrxyBkOqSEFomg/iMC9mLL5/G/Q37zegP0g+9lJzB/pI1mwNm5mFHyAmAdeE3
nm4eBcxYlGW/NrVdbFo2VNbDY6dlugiZagHv6Q9fohZjdlcMajtxdhC4hYxoFUeX
AMG4eqZhupaGDtKHkAg+vAyBTWkxpSc44jVEa4E6XrPc5B1m+aSreCzCYM2RJtlJ
qzAhtNI8s07etOO6GGQhzXYh/PR27iaxkOhBmF3KCee4CVOFOQUd7y+vj0i/XQfa
vmDA+Hbi0whVwwDd0UpHyjcrJX/8YORMhkv+8FZdoBxITh8/g90GQUWwfGpmDwzt
49hZu1GvvCHyugKw609U2wQl7b7g8RP3hIE+xlQJKxZH7NyX7hoPRWKbGxuxVbRF
q0kgw+1pKduUAEea60g0lXr7Wr6Y3dQtQ5+Oz6bVzsEgHvF75EGj3GSSpcJwvrMV
ZGCN7m03MHQ2pKGfag1MGkwBSHz9gTL4T9VBA1NeBpoaNLqazNsFU2SP/FKaEIc5
GXhuUGOQZMmWuje1Pxju+0epja6UfB+hNx52W43iLLgx/jZBmalN/7E9HptpyWVE
hI0KyG9ReLkZNWtwwOGyIzxIyLzP1BkQj+/70O54pdv8Mti30VxSWt1fQoommLDY
V/NVRzhX8IgLHyRpP3+7BbWDXNxdJHLto6yNp0D+cXN1nNcRxn6J6KXmt2zvNfld
Jv2yYbi1hPPgBqjQ/hjgHD90E4X8hTZ+XHNwLhAo3nm33PnJOBfsNlJNlG8axbn+
wtzEhb/Zz7B27d0JgJqR2THquYLr4YAttcdlTGKTfsHvPQ/Y/+f+/njeR+fT7ROo
Z5dEEtoKt6bi9Y51yGJ2VDlZqR/+HP2Mh5cdM5PRs7N0r5zp7wRQwNDSV2P41c4G
gd5t1u+fAKX8Ep++oyU4AMSkH3OyYs0ykCZfADX/bq8yK+5dHjbI+1EoOw8heS9y
VzBcQtRjUx8OopmyNuzpLrpulQOCgyGhbvNrbB7/AMiWNLViMbzQzxhYytIknSCv
ByJeYZDb8lnvAHazqnWYgLEVcIZm0r3o1AHHQxAdMUz5faWpVwnOdpfIHSHDZIrD
MXE3McuS26Szamyn4og0Wbqurz/e36NsbUbqAxwnY6okNn4CF8O619BBypPk9gPd
JC9JZeZUr5D5FHQTblZihIUlzD51QmcTlkzxELUfF5Nzx5woFVoBimgZt5kNdvAy
mxGGzMQVEk3DRGmILC1TXrnOfN9wCbNpFSESFmboLYX/tqMMdvcpSYuUrXnKz7cU
BiTnq0NFF85feef2eXXO+aeys9D8weOzrtVjTNUh93H9sMYliriicFBoLeJP1FlM
IGULA6dKZ8LTMTUHLBVzg8e7fU8Ck6Xs+139It1hRNgkoEzqrZlbHNneYBZfxTM+
5fyxoOYUuEC9D4cKJvZNsX//zUjeUeft2Ne//odgLMznKGa+lnTLU4CIHmOvtq/W
yBrv8yMVIpkXY7P6LCE0X9kAruBFd6Ppl9vO+ORfigrzRxPdvsCU1C4DyF5PTEmc
C0pPup+4wnfWtBFxhy/MApijLLfYpwYNBOhD5J39h34tkZMVg4WiyzY28wK4mYgS
mBjiXh59MJ3FCuzG50/uDiiSBY4XVIokir2kgzcFXroe90+QtH0IUsrYQP07SIGZ
Ajyuq5opaQyQyT6xCXM4UWrjGooLUvFTreudU/IK8pLraUVM8UygbeFUc5Ouy5C7
TEST3pCl+bYv1VVLrb3pt2jU3kxnRbyDa/T9woZ5CNfSnKdtdA1En9EzsLuphS6k
bpgZGl7b4YRB5LCK5fu6zqM8mc5KdF1mwPioUsGDBVngi3LpwTc1bSnSktkTSqjC
qhfnaSAfDnqg7C0zALSGidho0SMhw6q7klEvSuyZc1dX4So99ipH/khEmbyn0HAz
sWXSNrY5E6jl+hLOOFbW1cQN4GS0FJy96VWkDQp4Cahs+vn5WJLJQvh0YO26Jxqe
22EC+dAkiliskz5cYSmmU3ztiUWwBDvsX+DCXcnuopiU0knFOMR/xbtvJvIYLlU7
U9ebHJJys3huiEVNi/rTKff3ZLj0vieBXZU2/+X2/ttsRjwx9aeCAEsZzAr6tMng
9CJZM82ysQKV5PJrSOnr985aDxSZen7hs5S5UqowuxzDlu2YszzswkgGmPw8isBH
Ms+Vegbv6WzNEg/1APqX1vH3GwFMqGpX9m6mv2jpacduJpC/fzkQ4X3wT6CwinRj
YRAsccC42oHXzVV+d2kf9NkB/+egUFFRykmXtIY3BQ5DW7Wxj/WrrUf4D8OAe0u3
uEQDeLRgxf4UscAbawsAd2z913GHsC9PfXjt+rLGjqhSnRU79KPcwXJQRfhsU2nk
DdFpwYCzKEc1nIhDSjyvLM6yJhNwX3IhVzt+hiA1hwq82e6PkM0GQAXDFziaUR96
CnHy90sNQPe4kko30+ISVa7xxszO55sNnR4C7P6uAmrJkmLm/jdtIqXcZltPmn8V
rwkZ769JMvcMiqyBZZGmDMyvA/ARnbXcMEFeMDL9dMDIVOW3hlrvoX1L4jCoGMui
L1dgc9X3Neul0BjE32gAsldX6p2wVZ1gvmHeEKe1c+u1xCWdhrs3rOH0fAwkf5HL
GZ4G6FZxH9mg8Ed67YTkY20xwVWc0C1LeYt7/J1FuqDVWzLsdraLLdVH4+dTUbIE
hj8T/tdKStWLa6q6NOEECnIW3z2DEZXM3C6VGDRw8DulKiB82Slc81x/zWjjPQdW
SGKEfP6zEMI5SX5uruXhK2wrZOHtWA6RvdSj0eTXNhv5Juk9rjp2cSteE5rwO0r9
PTrE+rLpieRDoo2PuFSyoNLZuTOsOhTo26TNWphP+WqN2fqfTgFB+ekepYR7d6FV
tGHGD7HNpKjXAHiN/qj6O8QOfY6uzuTKfPHURta5yFxgmcoed9+ghevZ87I+9s+I
yqWzgFUZQ08+tDcq0HMpx8qowdH4zAHX03ufY9qimvb+vhdO4IGIEK/sHnfO9bwX
0FCTVGFaShOC59LiZ7l8ZGnPSwEJP0JTr8nj2JXJxies8eIXjTsmCv9mMIBWZkjf
bhMIFAoNahzQmu/PPlYPIWxY9//YWgnZf8oU1cHSGllakfnuj/Y2xIECM8wkULCG
G9A1hrExyMdC9cFi0n9l5M8x3u3HdHbpEiHRCWxTcDvwIkEF53om5p19dhtFb1zB
xOco8VbRxmHeQ416ZSIRgl4RgCYMpCSTTWRO4Zv66uk6m/xAxYZX3GFwfGVMmatK
BdOo2CPuNtVB0oJQ5LrosxoCijIeU1/w8ff88qBdE0EymELjoh7PA5hW+/Ja5U/G
mUP7zSvSFQ9vkeDwRQhl7tj0FyzLDudZiaWtCagLzOYUGjypwvYCbLAamCBWqJhK
DG9XVxAC2EAQ2zkJFQ/yLmH8pJg2CkpoHZC16uNSZPNferMEgJGI5YsrwwjZivc8
XW0bePpPwqVC/pQrd0Hc+eCdIWHpeiBni0EOY8VECqdp2s+dbe33eoffUsrY7Spn
cDfuiFup3wXVd4PwYetIlUfAI4uZ++0qWzpcnYkOmDVkyzwXLl6V9Jv/j2+14Evp
Y98uwu1jpqvgQcwyfPgruM1Mv7HeTXZFBJJupgze7c8V8fEDEkKv9C6DjM/ArB4T
pYIYgtls68nSge00R5WWGTwSmQiIOg9G3Af/m5EPEEV/VO7KAkr/Dy7Bx9Sndn9Z
lDRln59qiGdjfOPrTOxkaiOXxcbPm0nBU5+dKP2X3XGGueWhVKdQ8VzixptnfMQv
0V0QR8jrVNZI6D2S4EjA8f3cM9dAg6aMdWbfj4foTM8zrOs1zgDDfIsmUK/PnxWN
g1oCRJDAjrkV24aIKjDDgQqkYp8Pp7hlRX8TEAv8qVdl4wGzAw2UMo/NZBnEwGf+
eJtYn/ybqFJ582iVBiNXnzpjCB/5LIn5Vi9hQ/iDVi0H4R8HgLqOLhEq4gLOWRep
dwmqa8uvjUd3v28RwlfaTTih80poiQlc2xPlRR5PEItlAQkv6tkKvcsN2kpVAA6b
RItWqRqhG0wThEJ5bZPhNXi1K/TUJLs0Os2+8zQuRZ7J5Xm2XawObR/q30AGEb2o
By0wii4JCYOOEKRm3plB4CP877Jf8x+jKWpKjzS/zhdTvU/WK02ArSX54aLQ+61D
LIc8LPGO4pK+xCBYYdY8Unt2oBQpF6OL4fgPlZhQh3ej0K9jlY8mfR9ED4EaRNuD
zE0nNo2yByA1yblHzjYwKMbRO14GpLW/ow5lmOvHiqHiZGrry90X25+4q4rIrGYX
gMKM1D1HfbXaa/6h7X8ruggTOwBlrSY/ydp0Ul8mlQf4mt9HQsmANyBOR9yvZNtl
RR+Hsud3Y1sIpd6tR905NSb67S/GbfAPwQ0RujxPkdy6yDACjBhHfhFN45PcyGSM
/HnuVtDPMKSvW81btCNR2bPfB3j+zWteOOFUgctZ2n8=
`protect END_PROTECTED
