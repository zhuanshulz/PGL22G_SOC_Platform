`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e7t+3B3+V4SUNjyyBDYN5ukMeLPZe+IGMk7aQri5/j/4a1Y9YUfUrpFZ+wJ8WskA
NwRjzIdN4EJKSiVnvS1l5vrd8LM7i0ETjoqPawi8RqxUEprz7LdWN1piyri6mYFc
5ivcS/LdrDjLofDJYFs7LXGYvW8Onhv9tsi392XlDOi/PeFUiYzvCDmkBvKKejrw
PzwktIEkyFWogwXlfbPTsODP+Fe15k+00hHxB0CBnSpMIUDazms5FaZqDbxmILAo
v+grhAp6YtsF98IreQ33g6z9rPOxWgddjm1vJXsogstlcDJCPewtXibfmQnj6+GC
2KHAl0wBMQJ3Uy68cImOzcTZukWE9L0yetHxYOg1vXACjJfBbzrA594tWOdilx35
eO3N/VKR0YQPrg6Ph1WQB5K07YQZD2bw4BYxnzFzUPgHdlwkuDURaF8AJdeeSVwf
8U1xUZUx+q0e/27VJ6Oqus8ZibnrPhUzsGxXFAuxJorjAgjO08U5/Lr7QOhj6VwH
X0PEwV0S303w4vJSRS+yI3c/gHdVBKz/KfQnt6be3ecrbTTrQCtgpsHWDbDuZmtZ
Aroc2s5/P5LU0LlkWThr6c78+U0gUoKesEHak85PCjo5o1V2LlhRbpgBEMB44rcm
kMzMbo2eqZKg5PzMAEkoCT+ELnoJZE+c3gHmucxUYVlJ6bM2zrQXL+MJ51w2vc42
VQly0x7EeFZcWco1mblziyTiHJbfHgLDACsY48E11SFoY8OAObz0WP1iYR6Ahu+R
+GMbi2wz9U50QoNzZGH8RqSiBbskGS2+/6w4D7Bwy7i9xB3k/MSLrSUE0XS9Nxin
e0afbCKeiZ9Zs0aLvvSHstXui56eC+PSkI9/VmLiqSy9A5DzTckTwnjZds8+9uYs
`protect END_PROTECTED
