`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3eXv70ldG9/gKYdYHLl/s5EKku4drj7gXFQAJxXhEQpaCN1Y9kJTsLF2U+eKDgqP
szMNBkcjHvS0OFM0am67OhXlNaDCs9ReIh4nC1+sFscyYX7Gqo3nzYTT9Tr9nnL9
io1ToXfQLyIY+Nln0ezPxpB5v7rqlSyLaSVCcyGmKjEFia7vu29HTf9BtQG3c5Wr
vyOCrre1luRhpaAQavyzdFJXAQgHMweTisEjiqh63hUwyk9wbFQXTOi6+wNW0pIG
ODWtbO+UPSqnLvvaPQKNP4o0Hri1n1E5sUBRrBudvLcQLEDR09Uv8dYZjJX2V3sH
sxuTsmXVn7gmpjhsTS5Ggay7iK68UlXtRKdl6JQ9oEfzDfbk/PIYXbFsX4gvUg2X
H6WannlqdTDOAsEfE/b7vexUWVpUU3kkXFooH1GEU1KEmw3fjTKqSWGYb+lC4RqQ
ZTGcFU2yEheEN8uGfO4ps1gOtvZ1yzjjApLFa2wUVhuvKl17vp1gH3bwAHsQtUFD
FcFIfAPb90RL7wzhp8+CCtS4cx81de/oLyKorinSaFRFd2P3BIrYy9XfdZskombB
myhVCxIIFWmXyLdDCc06PoI6+K+09NK3VlfIh9edahMNNK8LiCkC5IPQS2u+Uiio
LgqSXn7L+bjx07pIstFUnWIYmg0X0gVf4CCJFfPcajpza8N+lF4PP8MWiUJEaz0R
ur1YJYgiUlQx5Os8a5WfpZtQv5g7Beuri9Aw1Ig6K4FHeZIGeu3JN3d1/xjmkEgm
1Bbu7wLZtXvpM5DtqoGlJ5qg3kXtQ1+SYJtG9H1igOYA5JRlJggaRRsRleMpZ3hC
dctTIoZJkhQ7XgKa16iRlBb21fCxa3/z/PhCD3SGPcVudg3TNgOpOMieYuGzVkwI
Aia8mgrBobzanMu94kJdQ5ERIO5pPL4/6yMhvrdV0B/7Zy58bsYKOl1thv2Gq+gM
mOb116BynyEO05D5QmTI/jzjANJbKa51OEd8opx6n0prF+kJa3gacQxq2CndeOiI
+sT/QNzjKbUoAmS0b72H2CDatOGNAviZoxH9gASZLX9xnc/oOvYDyE1W11tsNeml
Wp09sw2dVTcubpfGxJlnjnNVwk9fVSaUv01HHDoAj0ulclVOE/vQiTYsNrQIHFdR
SRJaxjJ2OoNADZg4DtaIPK9n4HwlO0vCkbnAbkpyDYgU1e3QNk03dOSOdpn1KBGO
wqxv9MJCJY9OM1JVwPeRx+jr5KEUvhyfD1z/0vphq6edHSpLH93FRik201/JU/jr
OzhdTR7IZVKGF8E1szCTu8FeTy9yFTYUO/G1J+Rp3pMfVdD4ljJx/+zQl+CFLEnI
6uUFe02yiNkiaawDL9H2llQs7zp7rL33id6STl2qMMczMfa4w6OJkLnq6k0S+g65
1Rh3kGT2HwEgaRGmQ+D+3fvO+bUYge89HNpvxsZCA72RArmd/4SMtc2fu2Y8f71W
dTGBtDLWTMd8CIyyXk/2drg7Kf9J0NYAYRS4soi4Xrd2kEkNBDBWC/bqBcDqE5vL
9MDUnZoGzXANtzTHXod+hrqJK6FDRKNguLoBvsB+m88iWBenkERMmTCR/9KYI9+J
AcwlNihkWP91b4QA2UbJnU/zjtyqmamSmwHWntkxeeKXRjKIKnl7Hmj86vo9jRKc
HrHQXpgUfzYOEiuMTxswhGTTwOwjywN+KndnlSVJartKO4muitSICVXT+sN4iFX6
JnzejamnM/HvvvBk3hT6QZmu0JltMUOF2Nh6dQcT5msW5DmIldzJKwulq4pw86qL
6+wfj8s2YZzFhUYPra1OIU+91OSZhLSEEaVzoxN0At4DXPd5a2FlKJnp9nTHvdoJ
KGSG0y1iWAuJrA3cED5FpwmOBnZDDEUnipFYRksveX+QdzgwNT0hlly0y81/ZZiL
Q6GGK59pL3bbsYgsVC/BBJsideliPewsWfchScROzUDHCC6AHHw8p7zF9Wo8Ikxp
w3tPzdXJRA84hEF4m2bCoyZTHEW0Lqz1biOgbeXt30vZw/6yhFef5WS3DeCzlrRS
I4tIwcv/StfR2aaoH3p8Y46HrlrQit/ZrIFOa5qfx/SgZtyfMCeV+iO0VOfNZB+Q
AIFGJ4WByrhc/rNaSI5jbEtS7jZKKa+5tjt3Y3AepuMciswUJg/Rt8V8Y1+a/UAy
1clOKwDHeO+fR5FSaogCg/eXGAa3+23vDV3sVjjGAWXy+K2irBTE40m7rBJaRBrI
9ADj/ERvE1yGT5p5x8fC8o8ngrNkFq9BE49BckV2PPH+qviJ2HumWLw50/ww0v32
Ntiauxj+BveP9kUh2d5azG4EV3E7lnLAqJv3xPdG7IqwUwKnPApNDhlbbXAVbqxg
MHt6YAFBJxQ/g+FAMRdxG+q8vaLnhdWJR98SgAAZRpp1ikWw1Lpb1onIOb0xGpm8
sXhQ+HKaIEOT5Ovl/0b9cUqsHZYKbvS5JLDGITObJjBfxLqHMuUg+4CTT2trr7fC
GdyQ0qUpGiJTgxHihZ8WQsyBDlquJ1TOwIn53fgzfG/YM2wKLl0U/1Ajtix0SnRp
VGi6WibpPCzcOehIeSVFyAdNf64H1nQqo3237SVH7Dxh3YPEMrFf7iHBk4vzAQar
8Qn6EULekeiLS6TMoW94fHWrYpJHvIoX2msRpCym4O1JkQfqu6fDpEnri9eOlu7/
NwXCEQPqvfriH5oJRjMaR62IvLyK5uuWH0Kq57AEApL2XQFjXQDpHiOANhgqk9OJ
4mSnBetpHSJP9iuA2dFyFiJUXwham7Uzz7msYMvL/HM0nyxh9l+ArIjHxXJwREQr
xo6IpzzufIQhUWYSFfwrvFahVk9qkNkYebBhmm+Z9p6DzeYhqJcngLwmKEB6MKCZ
/KOHq65XbUghPHXgiGJ1i0yDmSN2gvMNYcJdkiwAkbof3XLMcpF1UGWG4fbjf/4p
hHfNkFBK+jUrgNDVmBmzq88vahnilnvT8YfJ2doB56VKPNEQRtg/MQY7bknF80B0
GKkfpmE7rmDBAlgt9sEd4YVaLLMo5W6CniforC06jiqKMrKGxcSju2ANlGF96Vyz
zpMQsrfJvB2feNPPsg1ushSR/cwZ4yx37CKqmNNUtfEuFkErJRVW2QABcxTlDqF7
Qj8SxErwrmNakUZCUwD+Xkqp+b3QD9Us1B1Px9CXSUSxQwoG19gk6iuzzhAsRh1c
k8WVMqvPW22GNI4qQ2PgnOdidpngvb+ivLYR1bDboRIVJ333zyN2X7KksJmoJZ8a
K0xpJgbOyfdkvHD2bxziwBe88F37xn281ytnguDGm0P8qVzhKEG8DXEFHLDlNm8x
2DT9TjOTPyjECo5mLaRBOPSkHjrRwDV9Hi718CppJZWJN1A0YNJbStD4RD0MlaH2
iWUBewOf2SLCvOXIzlUrg+/7Yp/L+2XChJomK+K17+O8tADgUiMCjXXyxRSLf7NL
8QTlWNLK60ONBC/dZK/M4r/DQCDUhZ7hThs4Z2ez0doe7Yhlm0XLZKVd+cO7rIaK
YPEgAx7UwE9JYiPV2xhqvXOx1f4q4cLM8MHflAwW4sToj77tJ+yvBiFCVpRbLIoW
1IfNGKfVf+hybcjYstst0dIV7WQ/9DJYCXPBpJJRrLrWb3eYibwAnxTGaxfhbuNF
38E5mFnV/LLR72oyuYst1IwRDB8ePKIjhOm68+tjnLGXHkpKy3jU3+vUAHGhhNW4
aX3DecYn9o4cIITGbtbFAkf3xhDXNm5hLQSB965IgeLcCIJ/mFpeNPUg5pWW7BKP
S7k7u4bFWJZWKpvI8KYM9DR+fymY1cTzUrJ5DxskCXRIoROHTD9fTa8nrVfYo6Gw
D2BHyb9Y8mPY37hCLeimaUQECZ5SmyANiGVc3EOoYV4GV01ZJ1cUQ8OuRZ/E7w+k
EsRR5drreDtKIc2NOrLk/bSk/mS0yZWaBLJ1aoqQj3APsLZsReMK93mDR2b/lY2s
X6JHHohyXyLLuP1qpBVsRu9HhPdSwH8sXUBBf61YBjj6KI0vHIpKj3d1X08605oC
GaxEqs907KX5ASOosAa3L+ErSX2tiQfXN4/e6RkzXjTKuz5Rj3ehb0+7aDOKM8Yd
krhz7vcSO6c/XCQaKYxoApmmuZ3ghaLVGFJdkrWa+Hh1Ca9A5xCkQDeSfHq+mD8S
hyrMoOEq81Y1PVEWh5evF+pjXeSOn1OR7dmlzdP5r+2dum4TQGjxqIe6WsjlxVTY
+64d248uMrpgsDxEPvPSWpqbLIPWWeFDJHuXMndzSk7g68/jcjsRrloVBXnE2I85
yyM2BNwVE07OfvTYHiWH14SYzSD3X7Vts3dHTkiZzCjdOFzkKi51Hg+BnDEQWwCI
Lg8182IgKnBI4yDXWcGqMzfCA57qg4VAUwmGymvS5rdA9fYwRuhiK+tTHSOMnvEu
ETp21MuskUxhqWjvYLBX+TFsi3BiSBms+rbJrfgBm42pF0koWvjVfjrY9AOHhWPD
4WnIhD30/vw5WMsez0nkyWl+rH5Xds0v9TyLhbSrc6BoeS/Pabu5/l2W18OIG9ir
qLDzPIMWskB7FwQEKbjsXA==
`protect END_PROTECTED
