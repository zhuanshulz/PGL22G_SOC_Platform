`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MI8MzW2RNy8VOo0slXiIDH8e7Xx8WxgbcYOLUoCb1IGPveDyh3A+2H/pG5ilT2RO
UvbmcGKsbjqiVFCidKqEbPcTvM0vhi4MjLb9VlHCk95V4Nk5Qq/6fWloBrm3Daft
Iy1rUbSgVb6IyEE+mSGot9LsaW7Ud8Jk9NeglhHz8RtoR+qHXjF3m4eP83EqJpqJ
avByM3Upsp1X9OD2BMGADEL09kNDCl5ljxM1EJMCfLOBMz7oQ7abUk+/fEuAdr2Z
lFNBMnk8KELNYNYpKtSTBlasTyK+NheCservJSXo6gOK1hY8zAt9Zw0ZQLVZaeNz
jzqqDuSUHXXpRS6maiNBH4lPcWUyomf24LiEEB6ZjVrakTRO7Ea0TqvVeEX4SSMb
VtfunoylrUSOryXGGA2z+jLj1V2ZZIgOPFJI3V2MGU3AioUoYng3949dFILSu6s9
guF9B0I3G80V3D5P/MDayj0TxkcmjbQG0KG9hlITRkxTBETnlhJFVjMZIXxV7cKK
y2pGJp9oYIe+UrJM8b0KJQLXNJaAb2YggPdhCVnlYHpwdWWOn4TBe0xza5WIdEkE
+aZJOK+b/MNSS0Wcmb2SqhwEMSKa5VssL5K8gWKFh4n1RTuHLBiAvYZXVtJCn1s9
5u1qc4SzVdWLlylNaIt7bYAzo4Gd3vR65fxIE5INPUHcmcaiEar0BoABBnpyixG+
ImKt980RanO+uFVCaUuhaq8MidYRFr8FQ+MU7CtFzwlxmY6iKjiIgg/AUOu/7hoe
Kkx173fJzfsQ9Ei6A3mGCX9lDxUs3PHdZXwaVY8U9GKmQfVxwZ8ajjz5rKrycDiP
Q42/GGBay9Qdo8QLQBw5OhC+6b2GKieGT955gmTPMfnxP96E3E94wo/V6s+lkAWY
z7sBESo4FLU+SLkTI+WtZs0hZfY9qFVpgElAhfxmauVVwwsX3dQpomuOUawS5lLj
I1luN5TaVcwZ4omFii6ULVzXo1KXTva4PtVVvXIA/zIC0O82j4bPONwUvDFrL+7l
Gsz3gQi56OfTEKakMDPUkWrXydMqdmZKTqsDsjSHi1MrJlXN4zqCrvz3x8SCsoJk
Bxj6G7jgkh51x6HiqGi9I1Ubt7Pp0eSSDvrurfjIMHTayJgau1T3RlEUcR7QIKOg
ojBxmvZBGVXTBW82jorY3S4yZkJiUsGms6fJgJLrkzFB3Y2YDMVPDkuQt/RqmvNl
q+Vv3oyzFazcRzo5dDIowv+2Tcln80WVkFg0Q18UDhXtgObXKG8A71LAm8cYGSlu
/xq+kRohFgrYunqk+vH/b4dyrqKIaqp/f8zMRDNQ8wm30BLARlRKc88bQZWJvitl
JgMTtg4Wbb4+14T7PEUG/DyYT4NnVVkrgXrCtTFzBgJIrMuHFmAtQf9WKcDvNFdV
jqoinvYdwXbngSLdWXlsqxBw4iQQPyRtJKJgtZCRNn++BmEz6BBL1k/NShZBxhfK
HnXxhhyve6gGN5nlW6IRr4SZaRkr4gmfrV/wl7LDi6x56igCUgyu6+CazPl3KWBy
eYgNpdf7APUUGSMbWLk8SbO9zWc/jrMdcBrHR+bKOgTQpeojXwxN/yLzIuB0W630
wp84ugT+b3ADKAY+Su59ocdIyeUJFLNlWbf+XpRFyktK0Otp2b4D0h9v/vC4VAq8
+G1VRnHxmeIrvyqkbd/RTKnc2dFXviqSdxESG40bLuzAVyNbVMXpgKaDbcY30QPe
0wQGHQ7RTTZAkK9K3tVobaswHGDrHxPG5LyMNWnRn49/GGdg4jcD4/gnem6jpSX7
9i3kEJEBb3IzQXFjbMyeIpCnUNCVpUwryFu4T8t6Xi0LtkN8joA9/SlqqIZO1YoN
RSx+sCkjKeM2/MxrbkKblbGl9aZGA6+cv56WeAMiYQllQ8P/HAWwXqGF0vPqBI56
U108uc4jVLnAWm1pisHmOgkZAEMdrwb2Kvzfqejg4MNwvBbBIERRN4anHHPbHDko
rXjnYfvbbS3AtbXRnAKVg1MnMMmRGTMVCutAnneG2F1l/Q8MWIAzWfOoWo0O0LqI
Ze9kmDGhI4UzRkkvoNMHQcc+QFjPAJSkG//4UXPvnS+6Ss1nAZPSLNhsmPwekeyb
kD5ZQtIjl/gZQAa+VW42KX/72U62pIhfgeVgPgNb1G7acLkTAg2tlR58VqJ9jb6f
AUbBMghfLuYRo1WVhAXdRYtUbLqti2iXNUq62dv/rN4ttJr8+sSz+BGvOoAVEYLP
yMonQk8L5EINqedg4/yotG5ynQ7VAPHHP4bxybcbhGfbuk63sl2K1kodqj+665zf
Mu5mnjcNBhQH/nIyHO8pM92J1QooGmLVI7s96PStN9cBhT+0nuDsj7K25m+tm4G1
f9C5oc33AE0cznHb9UuwAcYCd5SoAjmLG74IVTVkIEQwMfAwrGhyxWezYo3TdEBa
4P5K9fAPymPESR4NsDNQ42B2TjUq56StRN4z6wNn0QhoR1vv9wIfGCurp5VaYVHj
GN8mvciIFQEoLfrAVE6jq0xagP3KpnQ4C2yfvV0HPR9AvIRqqr9MgO/mu2Mhk869
jSENTIjKbIK5fjgXdyB3hxePpYPDpnU+tOUVltEkA8HgECWJH0/f3gljjr8yhnm+
gaBmgnEr7gOpchwC+xoaOUleim/5ZpuYn2+KF8MccL5UgWZY8W1oDSzNoj2or/CB
J9zUj45MqZ+Pp4IWwK7za0tSOdIw33GWL7Y+QE/NKUMrA8jKIv4bviiEjRfGNgR8
YD9GoGbu9r2VFBdOvxzqpL+I305R/iuSaw5Nd47zqcC0BhQQoh3KnzJibfKsR2c4
PecnS9pODsolbYXrhYv13afPynpJtRinwZyX5jP+H9d1i+GXqrMyO9qOtYJceBCe
H/Eni6dnas0hKJC47lcA6iJNiIvAfBJQsL+fEk4P2Gfc8gkTHuTx3f767MKztddE
hf1ezcFTozhh4FRAG24ltcEPgAd5O2rFF2VZtbVZFE5P+XA4KegUTcED/X2NDFY8
yy4sOd2cQPYhpGG/Affc4AZAbMJb2WPgs18VuH3SAOC6Hrq/HYIMD5omcewqzzdt
s2k6TcwD3zesasr/0ObEyN4sjOad6p0HZjmoG2UC3jM9XFdRU1dUo+4eHv6Pkc22
V5hatetNgq4KUU5cDteSa0mapq6ykVQRv0dCgJfWMZ0I//WVoL5rDVQmPd5wIpKR
ibqFGWnQI9fbr/Moeey2Z7CEOO6CGV6+IgFiKcgVlTqnv5Xds1M4PCpyw6Gmwn6S
QjnvVRyLknEGpbT7rNJ5MzRoxLbxP8WVc/bd0Sw4zWUtEeOcckfgTVtn3CTZLHTr
sTGu+GfDqcqujyBOcvTN9yaX+nGxu0wLqEu2BiWRAbAXi1DROGS0YhwyYboR5D4+
dTaKswe6HPW2JGfMmZOBna8FYjRvbZnBJqnqlyy1NBQ8UU6FRqJc+HfOIHX3rV/N
slXAkHDxa2L2Vd+ouGVB//8QiaQ5rEq+AZB08LpsJ+GxOcDddqEnq4WaKWHFl4LI
SCQseljWvPLlMNbJ51zYQwrhQ/24JrYcsE0KBJg7yvsYuZjYWY8x6/AnLZXDxpP/
kwNPHACeXFJiTXdixE3lbkOci+I29f4fYLKwVPrCU9tdHwCRq5gyC3H/+MGlpQU1
jK4Ipvw3iFejazKTK32g1gFxHy9baRbR6TFdGp0U7/XHCNHOMz+dI50WL72EvpCx
VO8earH8sTTVOPJbj4RgzJpK25dA+QiIfZe0cjNRvwt4pFInl3W09uRu7H5eXJpV
urk3jLnA0FrmWaZn6hldIs4Fjq6m0R20FV3O4COBjJrZoPXAsmWZ7s+6OzX1p/wD
59X0xVes9DWGrkAwdXoXHbuESUtclcWr++Fl1204MgKZMciEfr5YxCw48lB0gJRy
+uOFNjZcW08poBD/yB/98gvtijLSp835Bm9SjorbyAkcjC6netOZfy5NweTvycHc
yecIl2IiDC5giErkrKUkzaL7O+vxnHANx95TEHQRoZjF8TKR0ijwPlzZmsbp+urG
XjnX0fzTzvkLwFjDt40dEgpTXU2nv/JJ9loFNDiGQnBOz8VFrRii/w9/HqqJ8Hw2
ebIJdylv2TN3nkBlTM+HJIIxpqSUCWMPFoSSlIOCm4XEPt3pwYVBZp76jGp56aMG
F7JyEnJ8EQITRuu9cdZZZpHrFAlq56QPZASm6vOvK4JDBLwlnOO+OHpQMYkhhcRR
HwPlMCNf7CGNPFMWG5KNGQMg1R7DHkuW9ElYGi+bRvu/xUeev9r6KxNdflQPYhhO
jrbwO6U+Dt3I/j8TNjN+GeaONJkWSbRLHUxR1ZorDSDtD876ucikGWrRAj1UgDuo
HOqacx+hczms5V+Y1T2C2g==
`protect END_PROTECTED
