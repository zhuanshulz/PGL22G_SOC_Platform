`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zY1/rCjMN6fcPlsZORqicT49LANkuq3ItSSAM79394lBn0uCcrPE8t94vdzTDxht
ATSZjL5KXZFhFC07wgsiCp8wf/SdZbvP8yyRYbojItG94bbMaZjcF6OLJcMy2Fw5
7txywd5CfZtc0T+2IREdi6jB8x0x+x/s/Jxf6y3sk/e9CLymxiziTtKMKDTh9C2B
kS8te1PeOFHcXPtqD+drnxfLIJk72Y5cHPMrFLuzQTOOIpJCQb5uHFa4vyPFv6V9
ykQ985PmPmQsp0xBW13bNTX1uAQXbqmw+XH0zCuzkY6aW7w61ovJg06GjiRU4ufz
WZDO3u/Jemm6ZfMHfNK/5r3hU9/gu02kXbo7IRWdA0KSGv2JH08ClQIo0kU4nzeR
xkTrHDlqsYmeyoNrMGM62c3r+VMMOlTIDVkNL16/M48cQTA1vcVXZ+PTPAJzb/cG
wgAPI7yDiavFhCwITKYg1s8kqMoXQnBLwAwhWosHZHS5TvVFysBf1XxFdoXrHRoh
1+r1PvWj/8QEAykL34bwHged0VQFo0jFnt8n8kCXai8RF8sTdzcTxnXqb6LvcMuq
2SxKSoG5YC2mf6TI8+8ugg==
`protect END_PROTECTED
