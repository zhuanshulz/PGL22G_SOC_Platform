`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NP32UNG0t87YXNAXXKKILheJ9amuHl5++JvolI5+G6xObnp6LUsvTZRkAs6C/QVA
1e7ubNxFzpmfD++ReDPiA5ex4SvAR4fD8aZ5T+kCDRhEo3icTFzQm5y47JI533JV
f0XHV9IKHTpJRaniMN2eyuQXLmAIGMEQJ855r2kaQeAERsIxKDaGLl+Gkk/jVNXM
BEZcGbQuff9riG9x0pMWjjCuiYCEUXfhKkcRR9cYjLjzhWK7NZqM3It2MsmwWkGe
p0k1nyR2XOvnikp2LDVUWAg0PNQCYszJthz2nUbSsXCONK76q+7KZ/Zez2eViBZx
tgGVMAjRXGYcmTblNTXB6wczsrJAVE/cUVccCFL30EVrSHA+tbKmoym1DHCBnMcD
taGR1KO2mATxqmFnOReZioVR+GB1/IopYqFE99cAUtJmHk035M8srXTwsTOC55Na
aQ4vhdHWOu7wSjtsyYSfNaXer5KoHyBThPFYu/NOHZY8d4l9kux6GhK2zZOZFv2d
q9E6tHOuq567rh9g5h0TiEmc575shS2usdlA2hChNVSNyInapPnCSOa+6HgYb80Q
uPMe6oY+wK++9Og403CSRimXhwTZKeiasHZ295iYyuDfctc2lVMhBo8ZP0LdeH2J
J3Y6oiAgEtHETWGOEK0BLk38R8wKFL7fpC+ta8MEwETHcesTkRIsqSoUQlEMAYvH
0wW5ognBLnAVf+69rFJmLRTCj6nwgb+WsQ7G49VmIqA=
`protect END_PROTECTED
