`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b/QqhgfzdWWxec/yM0cpAnSTK6/33IBsNsQc/oBfvJOrCDzjckCJLd2uG4Gg/Prw
Kj25jfY45y5kHuWcZw4THNOqcM7uUggnIcUni4qZZJqYGalL6K0Qfw54gdoWyT72
J2VuOeX7HzuCisyp6a43jK8ZCcPHWaYbK4G84xylkRTV78RUlwlSDcoOCBfZwPA7
77sErJ2pOzp6s+Y0H877kenWteHyLkOI7BVEDpmsmbPLUgLP+8Y7zTvF9FHOmZ2i
d73OIdYqRDsYc25EDBKRHMqBfx9weRBJ55j4bfzFCWjMO5amZUb3lMUVy/S23d48
gyIB0JcX8nDiTO7RVUcLu1AnDarKQzSaDa/ZQYBNa3gPxakny63mX3VUTot50gbT
U4YIQ286+1dMMYDAq7pijfPvL1NyVXebHzdrUFr1TrVyl8aFp/qO4X4+THZh8rEJ
7ungSZaaFm9FRDY2PD4jQ7o974PVDjimbEBHUeBf4nyWkUTxA1z4fBSBryCpD90W
0bonqzTrkTAflwH58r9jlYJh+IfD5Qq3EHtbtd0EpZhhQyJSHLp0Y+scvJYGgd1f
GEGtZOlvmvU6tMczmnvvv29QuSRhtA+PXrOLaVhEKukZzAKTMRjA4lJ6scI/Iuss
tv/6CM1mPl1+7vBrTLCRTIivZsS+sKvTo6Yt8VJxh65NA6ZP2CSksJiLbSsqW/QN
E1It0H3rAjB52deleiEKNvcvcOCrUTFq2BJsL7APJ08lGmMwHrdj4PDkCfnv2wNg
uK8y4cNDLd51DM68su9mAI2uCaJzNKrRefGBcVGFJANxftcSJHBb12rnGUhLUJpQ
5ew/fPy1EEpT5Kl3pXRxwA==
`protect END_PROTECTED
