`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
niT9J3E5+Waf/PlNcKWIotOli5MZTKkeG6BlKGIfCt0aB+Efx9ibnpXECHos1dOe
gqVpzIGINkHmj2B/DRQKFs1Pl/JCqZsCY2DeuDBEUKDejJ0Cy868M9hZcrFkOvCq
oEfQeNN2YFIHaessyjdXcwfRFiAcu2ZXdPVA1GacRXUePB+fM8L5K9H+4kRFpnr6
kWExecdquHxqIYoH6AY8LJUhrefy4qHIr4MCDTpp//pgBVeD5qqKV6NnZ4VefJKw
reovrORFz5m/RZjwP7HSxi4QQG6jPwgww/uhrO7BMHjS/3HlqlYDFL6euPsIuEKQ
UcjehHvXqNe6yyuRYvBQk7XXhZMjp3GsCYWr4XWU+IJhy0A4jNIhFc39qtAMRJlA
vr0DeFjAQuSqf7t6DSJaJWiRwSyCL/iMPL90Mx4VNP/ovujFdmulRmRI5dBeN9+a
QHrzDSZ7zK0EL08MFKkasulq6HYBPyY9JBldoCZ7SuQSdSQnDf38LclYPhx71sVJ
YIDHQKBUrnTctbsRorXdIItJbEZ8DNtSHPT2LpruUIiNDrjwdIyMqez+wN2o2vlX
iPd4frb1yAgYCYuwzalZwUgpEN4VMRmxIVVANmaOvXmjNy0fltVNRa/yuTBHbWsk
9kMiEOtWbA1sgtDc843ENUjszN2svHuX42L7NZx4qf6aubXwCn9JbawNrE0CzYb/
rOB6p/fF1yFbOBllspRPHNs50PQZwB2/G+AdlysHBhUYNFsq8Ig1G9O7M042vsQf
RmNAlByJKaaq93mNnAa74Q==
`protect END_PROTECTED
