`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K11SEGymcCOMT30SIJL3eLmmBBovk0Iizal1A5IG7L0gS2uTwtjSI7qMWn15mM5J
/hMfnoabiae8HTJeaRxCOi8F5AT4p4w146M7+eyfWplFeOleaNSAzJzMgGCJ9bG5
UnyrBMVTyoY5/6gthTvHVjXcnZX0e7ZpbOWaKmpW/W1bgQODGLsZD0vTk4VqhQS9
9hNuDaI38Ng2Eudnk8gKOLgRtYo5MKlrGeGjlb+mPnlehJBTjEGDY6/yvx+i4VqM
d7rea+cPTcuXYOmVzuWZEhylI09jDv3gJH+9BUcs1pFnucUft2lT3BxQyJpF1K/Y
yOYgvG956uq68G9KwVoKXSIntll92GMv5JuzW5XuR4R2ksWGTmmTwP3ouTseKkoH
m85r0FmJvCK6IayyYr0cccD9usFdrFRYQTENZ6iUVnDLdYgbW+wyx2+0Z9DLMTxd
bBs93HEc8Q2rAF7omN0NXFCM9SmPvpEK8HILgLx1j3GxmXCHfEvaWrdNc6DF3fSK
mj8/Nxoc3yLzDXI783lC/dGK6Eb/X6WJQgIsHsEMLQUwrNdE2JlfJ6gJ4S0szq5d
xLt3ubskEkrBcTpcG+ofF25/DpZMEND2Vu/xlcObGiEeIBB5c3EyY7xva7LWawQD
ILRxhB8Zk+FwXYHdhdDY2FyuEHZj23/RucZXOLh2Olt9Bx42jZHPyXHsrxDCLSqT
iXMXu8MtpVosNzYs8nkiwxLsMS4p6yHpib1fYCxP1UCTlIKlB9himg1oTJYNR7dM
qOReQ5v7tIczFibcnb0TcGJvQ4mOkf8F9avbFhDGTVFRktxxaXBYiocfo2qLNDvT
mJar48Ozvie1/cFH7uRreFBmiuYFCLA1G+gCzT57FL7LTJZ2w2c4xnc73Vwai8ue
wp0hcY5DlzdvwPDHcAPcXk2p1jJIOSk/AsFLq+YvMDqnseeqsBoIySQpfSUZwUaB
qg3bYa1IE1t5D/HGYYBJin0HF+SegFRbStpYUqhO6uX2nZEr1wdYOgV+nO9t4ScI
ZXZn65t/Umsg+4HD3vNoINJQNdSw4l0G34MTD3m3gMKyXWCrn1/ia5QfogH2F/WI
MlEXAgbfBNtoeCXd2A5RHxjbZqKysnAqZ0LP+Ukpa3hHYJ1d1RoZ3tuNgbPthflq
z6TogR8JzPFdEXMkXT7B+aJ1AccYyeLb+v9p9XmNCF3aTEnkPcDl7BFGdKujMN02
lvJyyyqJYjdXHc/qNrbvWXgP/TpayvS/dTiKvb8jGIsiurgqaQkjY2qVzNNzblnS
W0NnnCB3N+mw9VJVaKDaKIcLOndn/Ki9Zfot+ElQz4wvMJAVEWp4I1zSmqbeztme
Jd4FC5VDFjGdPvZE+3QUoi3/ZxL+8FJhqKohF2DOYMNWf7G7XzKsjv2aF+4kHlr6
KoEulYdYlXjYPKxEDpdjixS5B0BkeIDTqe93/gnXTU7/j2lOav9kRyOfix+IHjyj
FSWd8tVlxq4ZKpR+ZdeacWJzdEkp5lU+1r4v8Gw7J2w=
`protect END_PROTECTED
