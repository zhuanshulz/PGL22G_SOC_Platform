`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ntw24JukDr5ReXcOeWkfISoCM07EaYVR+LeolXcMCc0RVEwB0Z7TbwXYsE4fbd35
f0WKO9511hcknnOdyVHfCEOLl6wJQ/XwL5BkMjjri/JAk5TMRJcX594wCDcSEjaK
GAwdzmXu6MBC9X59s6ZZ48GDbcGPKBm1XFAdz+JgqwGMEYp6ffSXkRVgijZGhJz3
DMdedbdyvStGPCSkCLlJ2M9/p3DTA5fLP2W0mgZk/0BElqvBLZJO9pgCkkkBVI8V
w6eNipHPDsw7x3jp+jR/teNwjf/ep96G0NkuS8Cu5swFgYRCugvvPLLJHl3V6gRd
UIZtsg4FGT2TDX60/h2KArSG3G/PK2/QT5vxoGpDjXts0V81OKFeoAOKMcZzMyFI
9aKL7GewlYaGNIuvYm0uIxNdctUCW9gAqNHLbSIEF/Kyx1IxYskWjGuKKG/ZvGOI
X++t1CKpF/cA71GHMMY3wqjTsvk58xdpwBPV9ZjJUkSJvfoUnG7ljSjcp7yrqxBr
i6tg+YW5NB3DXb0NRlanwSPw0vWAYIgnsm1MBNHt/0aZqgMS2luR2zRtRHHFhxdP
BDyXe1MYi29GGui5jurPLJBRK0urqv3yuNdP6+bqdBt6kTMZaBFlfa9eF91oxn7h
pFGsfMprWeVValtYoLtycSDoW1W9ifk9I9s2jBQ5CNPie3smCXKHA2UI9iSi9S3T
CrbHEMSSe3S4Z2xWdkeKlD/xdnau5cyewFjSlPHBf1H/G16nGBxoP3RC+ed7BDQQ
jqq2r3S6lMfTHlfDeYhk2EMipVKm9bTJdgFFw1mJs9vF8munfzh/3gAkPAOokJEJ
49dn6R11/UBi4Kf+D77+p0QSQBNEXjz9CTQnAemzSSi3LDO52D972GZKlBwl5iiP
jmhBriqpoylSg1u0sdZ99klZYQDemMalO6VTiW2GEOk9m5YMqBqnrn85UCf6dDLI
49dxRotpKfzPhYbdmKN/GqqDl93lYwYKCXC+MBOcQwiFxxeh1eTf5vXJTBR7AQMv
xS2cUeVrh0m/goz0KILdItwAtck03egpYcqlLlIYXpH77xyUdkag5gmQXpZkr+Bq
Q7fVa2rc0l+1azCTsFQH/5vd7bNozg4svzZvIkjgOMz1x8ii+mYTlJ8+qAjCZD1O
nUNVG9Nv3ghKzTJFUrN7OCkr4w24E/Cco6g6zsu/OCOhki7JMeRtxYZgHhLrFBvN
CFofPi91rTx+FQbSDGp8yRQQBY2l+YJLJrHrGsfGxccoJ2mZJxO4/Z4zOfPFYtVN
eHNgyIjQOHVx9k08ofsqtNpjfWuEYGz4owQV/ZpCUSmp+g+TwUK1NXOU7crVI6ZX
5/3bzGh7b0F9Um5dFhPup+Nj9xhcE1H7C3fpnRz8MLUYbCCF+3CD5j9sA9/WobSO
al1JlQtz27WKKdIeAKG9JJ6Bya78m/XY5llEkXQh75I6aabICu/+k5TToTjpHQO7
btdcmp6IjbPE9x4wkMA+dLTndjrfSe/VW1/p9Rdu/aAjMOCkfhkkL9mAJTqbdvtP
MHIln+ecIvEBvzymrmcIOgjX0ZLbgYouYjTuu4hac0s0nLT0XVqqPqT+lAjAHVjF
81McZqYLr1Wz60ByGlRYUBSF/MhEE20EHZ9BbKx/7A5aVSbkiDg99yEK3yvrGsFu
CB8Wk/YRCJdYL2VA9HxPChj+9xq1cB1rIMlFfAC7zIiiNejdbDknZ4GkkZETyTB8
tuO/poxTlMP4L4v5lQGExb0QSRzlJ+6N1p63A0FMtv+X14DsR6YPkHaFDi2MNymS
hPSJrwU/N7ULbzk95EOPqeZK/x/i6jxwUx/6hh95mKFrW9OFJqm2PdIBSrnhwTek
LktyzjOAPbpWcKtp3/fNAgyq2Ln5XJJWLeX67/SckCQcjrzTaikyisMQeOsGCxH8
fTso7lwYM/PLpsbPfBD9DrYYpnE0ti+ZSSsaF7s2tk0AOdGF9CL9iFUz4lc2xBe1
/AsorpDsNBPgjkjR3Ydb0470dK5KrEeuAxjfHNxPUXIXtcvlo5c6dyZxMSfGW542
emd2yuTZP4zH5DbZnLApIu3QItqxbnK5hmQhrtDicFQ4OjoNF9jXlvhCt5xclgU8
eBJ/jviwFfDQgxWKQ52NPOiVFZXG9/yuzJnXJlu6yrdA0TbQGJRV1NBJKz5iDUaH
y0rjSy1L8UjzQUMN0a7zg77q1iAc7PYg+aLh76/l2LgvLmZ1/pnIEyzNBjTQbrn2
hX7yjQCFFREphHTB3FqF73Ea1iOECuJdFCQtTq93/C3AFxG2wa6MECERsW8aX5Wm
OTAD4x/teRq4pVK+SLT2BNHxJls5+/vll307pfHiBdUXcLHaSG1fZG14hVg5ol/r
ynCzUgtldQuWTYy7rzzNaQ==
`protect END_PROTECTED
