`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UQkxgBM/TLImHj9oc2N00BH3BSq7CZTTErDSwWS8yEs88f9AOpr+zmwOSY6YaAn1
QgdUEVzGFjPJrywO6gAfJydbOAd5BSkG1gbxQsGryT+tMpJYRF/748gAjtAGzNY5
n6x/aS9Q1Le+KB1SwnNQdAEUMRBpmwnlqxCOwaxWYbPx4sIMd3/Txd+GY9r3EKxE
+3IzSEcOZMJW3jg2uKZqiS8MhygxrpN2N/XzBhqEEayox8FOsAyvpGDoLxDgHXZd
HViYTrCQhRKVdwsHFqZtVCrCorybVnVNYZsG8jyYrzjM2Ag3WlDwGsvEGdZa613m
yXAAe8cD0dQdZkAu3VFkzJAD7vfnSU554lOiwhfN531O+MmICsLHOI4IlLgSZkNw
EH40UY7rcPsKraSfm/FWdaIXY2ca7W/352WHozvEK+3cakLvk+T8giwbE06SQTl4
cyO6sN8wMqU8VQhcx5zEYolVK2BvX9kYr5a62XDHs5Tg97DfpepV+9jxBpnpz4it
CsYzvbwc7Gx7KyJ9aK3RtA==
`protect END_PROTECTED
