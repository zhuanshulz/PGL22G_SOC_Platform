`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iAcCg1ljPqmqe58DnpKpURa10hKin9AtiKOVjRAnOxGUBfYk+n8MJwlXGdy1KdGv
V+fhLsaRYpcCK40XRjAIOZRWbJZ6hRzJ+FZjYdlvdd38hrE7aZAW4yjEIEX8diaq
pGJlkQxPB3PbJsIY9b/zz3DjUDDaicT/V288ed1M27jXEoxIkekSlxS/aYJilNkF
4mt43oI20QO8OdAAWw60DDEjQLnge/tPSkkUXWfL1ufkdiqBjQqXtD7vxgReSe28
Ewz5e27SlqqJwY2GygpY11HCMTGpcyXETkbv1W4KAIQS5V6iIQBQhCqqLRYp9Poj
Iiwr3Oqs10yc9SweFdRYdkNx5C9ZjfHGspWyT/7y5xuhHdFpYBpFNGsi/lC7jrOE
PNzlp8ByRhbjgZQg8cu0BuHisVsBaWtgqf343wHpLgn9SrHVSsHnik5Ks19nbrfS
`protect END_PROTECTED
