`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/4/xFrM4VJ8B0FnwjrMVGAbwUjYUdK7XaM50UjnSc/JFGlaeOz2/HA8ZChoBkBgu
e8s6grhd0zXFCMjlD6d0FRWNnFoR19cKh4xO0mz+jGfHrp/9q/5B17mKCt5w1SkU
MBX3uHUztNXJwdc1aH1GM9GpQc7SSCMO9NY1H9/5DIDH/gP0q9aRQJOJeBJYx8v1
5d7fmG2+w2L5G6+xtQDLz7s3NA/tZO77TcU0JI6piRfvwo3zPm6148fF4gyNZXSa
FC6xxg7gxXMZWTgtQlrbxipx/6UXhVuqJu/v6JmF5fkIlSb06Vl+vXlsN4AaLvEv
sI1rBxGQf9h0mgK9I1TLB4xLI+Bhac8mhPwoOrajAkPtgHUJUkpbS/owZZcbY2KW
USh/ZfShjqbMi/6wtOGvsAeibGCapy1uKQUTUYhjqlsmWK91K7Ok9j1dSs6e8cyh
3HfTkaE08LxfWZ8GATnZ8PG0y1HbZb3WKimvwE8LilDaaE7/Hun+K0YMaULLWBt3
Pzlg9O1leAQvxSalSEYioon0kNH13X61OaC0tnPykcybyvppZeYcV5eWZvd62M53
C5nPk0QTmt0rlvOmk0ZCELfExI4dWaIltluMPsqtDRsmYDMJYVmuRA2DEgyqz0xf
lXMl+I14uFHEFBN6pu6ALsl6DoUw3NzchZ488mXlJR7LP4VKeJP6Aa61CnwN0LCZ
+atxPIB0R46akWdekMXdZrVFUL5M3Rw8GPq0C6g2jVe6DUYcy2sZChcErZ/fwEvw
1yMm7k+F2wWfIHPEznYFzgU0z2ecU0OK/F7uJaVWj0AMb/GN79ve4tbIVFHVUtkt
nfHnsWWAXARqQLH0eXJRmXxPW8Hly63R6KMkUjcAulI7FDeW+p1DbCNi3FSWw3tF
CBT0KCPPvow701/UFUM1C7a7u9Hr6XmpqzW1CypCmdJtiuvODJ62Mash+wTNSUW0
eWtV6fK1GaDvWlZuHL86Uh9IuiIcywUG9HbivPCFUSU9a7WHuMHmoc0mI4eoUmB6
mTRqg/TO/9OFlZOqH+Lne1cK/0BNgJxtYOsp/vOVNZF8q9f8eFgDqZPC6cONYnq2
4KMTp7PyVFjrsru95EGbasqXe/yh+Ho+pcbC3cF6UK0L+ISOJ+W+q6I648GjEQFw
Vq1OvSb7evm23MQr6cvlPw==
`protect END_PROTECTED
