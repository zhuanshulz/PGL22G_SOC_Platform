`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CGFFAfqboc4ckD5uwhXpw5JoMViyvfmaaF/iY8Q6JHD0MggIMoAw23eq/XNvAXaX
i4yY4JQNG7SXIKOiswgy8Hy6lnFO8xkG5fYKOqZcfbyapo0wLPm7n66+iHnFlZgX
EllfoaDA2XCKrTu6nNqJ70+r10oEH8et4Rfni/x9xNpDFOIpLlGg1SQGHGT3R24t
7ZBU+LzpODDt9Lr/1cbNOFN98zrJ6u5mWCnJTxOurGrKEVmhc28Opnk2ukcijH/v
IuZytmcgpfimoG995k/4uK0Vxe0sDVltE7XXExarrDmbFAuRyziFAWfrNGl5axWv
ZnYCupbNTvb4sBNJie0QvaaUAlNJ5mT89ygve4YeMpStI2YhJSNliIoLWBTrXyg5
Mtl+vzpnA7T1PS5jEzSJvpRzqibDFJBDEWgob9UfEDTaeGWGHbwszTKsCcv/GeSS
ibImXV6tXTkb9VIq/22o2IphLh9VeEpJUHfFiOh5JYQrb/4BbcwzZzGbTDi4GS7L
lF2rr3xrCOccAAI4H20lIJB+xbMBxx3EpRIVwLQVfqsYAqAY2wssFqmvLhPP1iGG
cqCGDv6B0xDLv4M7GGmDke7D6BlItw0oNvSZwO6ds8y3gn3qMW2b/IXy/nbJpgGp
oDjkvhpZ8h+sp/TQYUKQc9kd9GabIIp9ZiOpC1vYB2rW3tYjZn+ih7Ry9eS6n5hz
CqcndfpquMiS8lTkqvgEPHLx/9GhLIMOceuOBbtseEgnsqMnon0EzW0AkhISSY5q
HdOX+Qk50VM6lFG3OHKN5iJv1gAXdmCaAvFCncsw/G4arxygGV3lN981ipkfydiD
ZoKd7LhacdsZMJBcQXnAnWqV0HVJfvZMnziplUwESDciPhCoFn+k/NJilto7AVh2
YhZFJ/RB1j8V+WBQ4O5pUHOQTlhXYyaKDQWRuErEx0wAtyMycv55JptZQbVOyXhv
iwlpWt+3IKfNXzDThN8QSUtoLRtyikgld279uKnur3RuM0nA56QybPU7qjgfYYjt
V4GqWdu8fp0YPe+PjyirJ2qqOpDm+MCtr3XMI3K8wzeoPpHLtNKBpHDzDhgPBux9
0rPsk9xxpl1rD4oX7sfv2tyJzN3o4SgMPZjd8Pkij4DcKkIut+WRP8U28zzIcvyW
c2JSaAJ8tUZoJUpm5UusoBaxC3VUqiKQaXv7UIh0LcBxs0NM+b6pNnq7dzNk34Dn
H0qUcKc2g4jFUNcNFove0ppHxuDIWTmjQ3RNxQ8uKZysGSIuBa828w8rzvF6oQI7
9JPDFbON3QLUlIJ7oSArww9TfC3dLIEXPKg+2nZh1VT1dUNcfIZvsFRKPVFOjkx8
eNSyQ9Kp6TVbH7JXE/otSLBcvV1qIz1L3pRbxv6k+c8OYcGh40cqglVh16Vbej4q
QRLyCHaMJb4Ykpa9UGWe3nhy1XAXrTOUcL48GKKbxskh9Z2M5Ss023KxX6A9zQFT
UgCpyCaQl/OWS5ayiy0J0xqTbRsfxNIw8zuv1vrRZzQmvuR4nBAoGj6xAeACzDgy
YkEThH+u1MQY6P/BpXT3kepICnJqS+7ZOdVb3TqiVXHxHA+7hLiHlvqChbdgFQNK
+oT/3IwhUfTY2Wpib/GaMKrAvTlT8QiJHRlfdTwyi7d12PZRIO/S5cgKn4MN0Cjf
fhhyfCgirzm8E2P/EHdSOgmIUs+/sLPuvWjd+blmjwv8qrOyj3qd2SJ3UlraHCGC
gcAQN56Oo+Iab3y3CaA5Q/la29O3NUS3r6mSixITmt4hUl92NoA6DQIh94Z//qob
UfibySL7//IoUEZwKzbIhBxRdUlPDOmyjQWqNj8mm00Nfuc7cvQdqcHaI51pemX+
SPwaIMRn/tnDvcEImkBIX4hRk9q+gE08kFQcVrWPTQzCgyr4WHtX8zv9VMU+dAnS
TO3N+J9lrzp9A4U+4VOcCA0mPcQ18j0qOoYLHfRr5qeVY7XIHxyTY3z0rW1ofbvO
Ll2KPWJxbk3D0kCha720coR2odbcUrrjeVgM9plnxmxO0wjc+aP89F6agiF5lEwb
mIEcNJMkOT2RZ7HONk5uznoyt+LTVE3v65BeK5gUvwZ3j4o4cOROoe8DaUIfdNvn
mRp1IYmeB/sI7cur5UDHcXzvZp2dM2mjNkV0ktuQzhxkOkiTNSUGWrdgHcPJX+FM
zIy7+5cXXCG4KvHdBCpzG7PzBjrY20i+HVf3PWgtVO6aQC/SKYOwh519n8OPHWec
g/QkSZxwEBmXURrJbnGuHtz7YyYicQwv+0l0ZcUoGddDvGkVvKWLGQ/zCfCU4Mpp
k90Tjo5DMX/ZFC948z4zNXp9P9cmxaj8ACEQfbQpkMLTAXy3Q89btwTvSsTBV5dB
Wc3DvydpgEVIDUSva6O6frLOWOT7A/hYBpzo0q2XSTdg0FuwgdFp5IyAWIME9RcM
3iLA3pJJ37F3n5bQYJcW9fk+Xv1Fl+/zHQ2et3AN5KwwLM6ofbh9S9PMZHWBTsj0
HO0Aq8ovW9f0I3+uMtS1nidxIzoyOZ3uCCRckl/cKtqApDiTNryfGZLCdnhLwpZe
/p9PLBDqXGbWmHz6Oq/oT256xyRONCVlvpKZymT1eJlRl3TzjNoxokkNyfx7N9Vd
6o0ZVvrs0g0xfWcjK3PBtk41FZGD9K2V38h4GQRm2PTgc/RwbycFFfbOw66Du3NZ
DwR1j4Wwup2eSjLt90Bptp1cfXkYhIk3MA+BKpcKMlrGQNQF7l7hSKDJL6heUIKU
RPfSqEBk6JDoDdN55jJNbwpsXdB6qdqVxGE7ANkcX6SLWyf2fTAR18V0cN5rXCIF
hRkoP3s5Ne2GnEhUnX3XbEvYvNyWHt/7rOIS7E0fjzZLLG3Y4eKF34slv3mIOT4d
gMcV7gTb8QLyfwqdyRBHZ5ZEq1C7dwNKzUcvEoLO7GJtnPeSI7JG09TMJ+bUpluX
KsPHU11HfKroLVP1Ps3obdtZOurM2ZwI4Sc9/3xD9Pps6GcM7pkgi+ESUq5PyUAM
6tm2CkQ0C4rb90MjbNl3nzi05el3Pwo0z8/+kDTgrt7T5kqrtGD0X7CLd9LK9Poq
BJV1xulsoml5hcboOQd0lvV7V/wLDEpivVSqILo/EBXj+83Ll70p6no3GuWGiinF
SNXOhe6pBg9vc09VquPvUmlsOo3khFoefG0uhE5LLrJGCZyjIzP6sFsZNScwsDkp
wa0mErMK/c0KJX9gh1bawOY2+7VLGnTVpMKBFV9xm+nAntuYQ3pvNpevMm/8K859
NNws61NBwhCpXa3sQ16KNY9Q/c2WyzYWkl4U8F/gxnPQ6dc6FK42I844vAWHX5gE
pVhXrjfP7P3JeqomFhOFXYzA3cLxcOKMMRHyPs2F+JCNM+SU2yPGGoGX6aqKCVYj
B8Z+xp81ihYkMzTPZTkPX4j+orlEgBo2wQE2cjjbz9aG4gF5J1ADpa9oVU1e0Jfd
CEiXoGzvCrpzhejPAicJJtOIONTsjojjsY051JdijWB9nSOEw2xGDr+FaAwhIs3M
+GpBOVulfxJaCH5YPIpd88jUuv5eEjG2JLRrMwDRBs22z+kSQ4j3swZiZihCK0ck
d8quqwBG1M8iju9AsCQ+RL9JSU46QkOookLfrPt0UUfagbioZHzA4JxP5If9xAal
3RjQOj49Rkx4WDGS7dZi0kvwA3fUTqrS9BkGlXVHm//VNnF+mdJYm/EztXt07Urr
HqU7/rAbt2zvtAuF5De08TemLIj5PvpDKyh3uPkcLwXN9CJU68c840PQ7c9QOZk+
86BRmvqfBCEvuenitGpeU1CL/8t4Bpx1KE9Dd9DoLxOAZIfUj5QhX5ApjBQHY5ye
30NtL9r8OibZyAhhNWxv9SQtM2gw46AnZJAWO3lskt657DxnSkw66kLEMNbfZcd1
df+dbfdBsA3xxhBwpwgMwcTfDmVQiXucixSGiVKo1ddGalVbUU04s13gdIup77Ii
AUhXHxRdZTjuLCIGt96EsmiWAB02Ty9KXGJsu2K7j6ZuBHyijg0NCi7BwIgob87Y
oUd64Ljje1krMCHADmajHUSqNUda3ZDSqubpuPO/6JeyZB+9xZt+pAfMlr4K4Zda
LJ9AcQNFFYBol5FEVS/f0feZ0VpG4aMfTP1AOYLcEi2JVhzWcoZqwVfBMyrar+Xz
RcXh0lOy97FO0cbPVBRtB+elu6tdAAdzHX46K+oQzSbW6iy5F4zVtD5EfbX74EGc
/MebrdpEVhm5k7t3hBC9Z3QmmehtbiRFthEJwIqqGOBJHNv6d6dLEBepUn2b0iFL
Fq2PJdaoUkSAsPtf2iMY7ZdJ1KxjkTpkJlaBqLGQ2ALl8w2xRHiKW/Te7HjQHlcq
S1XJLmp+UMYy3bW5L8YkEKAs6claw8akZ3/ePAtP1Fgx/wmNMrVw1Zk0JqIH+QZR
VQI/CNdPx4fxMQSvsnASwOyDKIcs101RMCpwqhacE4BXDtYnncXhYf1idr+ldLqj
64tTn6jdnjsVrC1npzONB+rMTFsYSyKO74oSYq7LGfJDpEqDQEMV47JcZSqvGr7a
M3rp+Mz77lDCRtgj7pOhlbtX5V4Dna3KV+Lge5CviFRaPC0zymn0JTQAgFNjp+Q9
3tifurnMn2npmUGhMqf85UKtg/Ot5P8LUaIkPZ1jtxc5D6HOdcG8d7IabKXKKHTo
A6xPOxL3LjigZveQ2BG8XVEgBizlBfz/MVGwCobrmQVgoyFF9QkJer5wd3hVLNnZ
ObDLIhBAmbvXvcXhy4B4DOjiqTEKzUlda80O5vNJ2PwFmsQU8QZJPLCoQiHQPZKz
f8L7nff+JlvPKlZJpxM2d83EapkpbXXRemh2EIEaNnZ+eFTIf8xyqCf9Rl/ZEzyM
RsZAgtw8/XEB4+JTA2rFndgtJv9JQMp5l/fUByS9escEMjkhW4MuHYZ+vuMYAop6
7d/7D/SwPLClvGvUY480CeSQNeXrGOJrF8MMpdbsohE=
`protect END_PROTECTED
