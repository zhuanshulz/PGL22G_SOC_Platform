`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+DUizP7Hu/07FoRO4PX1OWGr92IALO5Lp5xoneNjen7vlMTkF1Bmmcm/u614jzEE
HQS5KIFAQgZb76vEdGzlvN1u4M0r/4L+qH9jUFW4zLfR9dsHnHm01xdfsuy772KJ
LcszMY1xqHizO6M6YhgHoWIovEvj0arLQItExdBh1M5ONIOFM4Z2nxJo+lS2KqN2
TlOZL4uGavWHJemwLCuBWma/YQC4uY9g6xOFamGhq6kYSLFOgqb+p5stcNtPLKK/
U8zMK6msJvR0WWYTz34O+vAW3hPfawWvvHEwlnaRcNXqx2eAeeBn8VhzHB409jDW
NP5MBj6OdIRISpTEtKDts7CF0zMak/vQpRiS5snJm9yVBXMjSDdVy5HFZ+gc439F
hmf8tQJtZvuzLVfMxMpVOXV05Qd90P6X+cf2CXtZYm6xFYLFew2x0xHKmvbtzf1v
q3yZeJtk2rV0ANyHticScpDzdGtGq7D+CBalTpEjvg56Ocr/WS8qvxlWzpCTL2GC
nrGrUEfdKBXv+wV+1XzU1UYnYpInDHKiusn/MxQtBfRWvddJf6L7uYY+z5Ws6uom
8/l2XrGtpBtS75yIdgnkXPy3I9osf62oRqRGhdmOHf0grekuyzt9f5SRx8ovR1KZ
9WllfPDei8uXIMqKzDKPiSqtTBGGiabtI81KuEbIX9V86vw5M1WAMn7d+fFauq3N
oZKkOka6Lh4PC9OWUtmR3mBJ4TiOlBVoLtoQc3YJf8HW7cf1vEYbWmd5ZbCwlQpM
3heaq/W+axAPNAbAjPYgBPRbayI6uW9YBbPImMRyu6GF5W0OrUP8ZM7vayRKWo9G
fulSikOpPvDWsjoph5YI68gWv8UZu9MnC38OvBbxtEKUZ3MBJaDzt8UavZS3hYS6
X21QhutzF04vX0Rp8xrIwJFgm4TZni5bcFTfVQFDDnUIHCQT+ZuKTTQY8A4abIgx
ZYaxeWy/neVWV8r7jbsgWPkeWiaJToCEZuB37+IlTbuVyjRXKTi4xaDr0/pOlZXV
E34KwsX4VPwVbj10QJtPAdkuwFmr9/zu5NADGh+tBtM=
`protect END_PROTECTED
