`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a+VFH1OiK3+cKPzkYO2Ktj/Kd7RIVLzm4EMTvAcAjYNltw+WYUcTduWHz2FEDCNe
f5HKTIeseT41xZkoMYbXbOVAmO0NglflwzTsXxISyDDu/vs6nbtolttLr2utDqfZ
SYQMeTnD+k7t8zrRkV/RT0IAjJE6oGaYvAPzT58Xy8ujOO319xsCZ4NB8R/P7WD4
7ALXoQQnvRFAsQmG760v2hyr6GN2mSKOo0DqrDU2YMaM/MpGY6JbO2JIq++HQkhH
PO1EnQiyyULIRxqoa/hbDqjHLoG7iggPLkPV0wfDbynyN/t8parKwGYRUoFx9BfL
k5dx4JbUuU8HpPSl2gX1PxcwNWAFq4IlifoSZHmXxFer7wznjTFXm6zjtqbzphMt
g3/Kf5JS9zpjToqKHKqdn6H/05xqLLYQ5opoDuB/XWtjjc6HaE7x16Y7H9rcQemq
l590Nejbfv9n7NFYBx4Feu4NGbrlRGk6881W7Tvo2EQLis15u9DjHan7OttWiz3K
iBotkG/H16nMJfpFP16U/6jP6pydZy9HKu5VNtKgBJg=
`protect END_PROTECTED
