`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aL3UwySihBXkz++gAaRHB5XB3fGjPUUEOEI9yftRgMqFaoQpCjCRbweGdlMAkWe0
sz0Y8UUXks1qMdvOygjfKdRLcCr1zY8kHdRpliMDjFdxq/C0kLj4VzrMjaKPMO9v
Tiz7gW4+2kDW9VKVnRkEBob16sCpvDyTlwHN/c+0lTt49Mejq6Oc3OpcxGK7KcX/
uYdcuGpbtNhld3yc1c914F4aqdpaDeosqIkPWTQA1q40o0A9xQd1dVmIDpSLWXZA
gG96Ccco6f4/wTUDLHfnClRIp542Ee3OA3W4Y+EGZWP5G7s3QVQNeJF+ShooRD2v
rjWCcw3zm+qj/RaMvzd0IK/1g1n60jBUjvt51/wS5vApyDFc6LDuB8KqoW1MEFq4
pJSK+E/CxaEIjdUJkYIguWlUEaueJK8nnD3whsinJx7AxqkaYpL0O9FQR1BFvX0T
p5KqG5B/Ekes7dAS3Es2vYaXyU1Wv0tp9L2tHekRHH0XEQ0prnHp34ChgIS1b65E
VYjf0r+8vI6rT70l0Xh4WnZt7Qk+vBqpJTNfviT4HZ9c48B7UyyLMqnpPhbj81aE
lxJQV1eFpzKSf2MhK+pCxM2yqdCAZd1RwbVTeIk/OH4sRQpGbDntYhCIf/rIKJyf
jshHNV/ungdS2zjKolnc+QEkwB1XLKXNdzhUa3i0ACIfR+745RoweYggujyOUqig
3jqa2mGbNTG/ywJtpNxeFeRh12nDQobdWL2mnpm+Dy+lxH7NXkiX3DlVf3MyA7vZ
/lK0tFek9Fgjsf1DAQMg++hlnbSXuQzi6gEzcRAh3pp04W0p79kCp7Oah5ApSd6E
yXNRIlfZyvRU8Smjz/1aTOZWrVWMK3KnWzOuMBtkxed7yd8QCGsr4OeSO1ZqJ6MS
8yuVdkYsFni3leQEI32lSt4lOSSlTR3T/Aiv1k+Bfu5wcb7WGY7r2CDTd3LReyiC
dM53+K2aSHgv/x4TyeIUXcFYbg6jPsOEqip3eDq3cQOxtbN+rpE2D9BzEkFaI/he
nFT6lMLIfMlGvZV2lRJ74fofmBhg7pACY+9uuO7EG/qus8GuEM4UfMbP8rateb2w
bEtNBBlWVdPv6e7Zw6NAN1/nDzTGu/6/M1d7JErK8gPNla1HnNX6Ba2cgpY6/wum
ucTfNJ7clDNHMtyLBCsMno/zs7TV2rvY/1Fu9Id97g05wLoDj8SZvnKMBLnOMWX6
8TDZS8+AGswKb0N8YsSAStI9KA9kta5/9L0WZua+TVToXF7SMQE6jQsVQXsScQ06
XWJBCXHpmp/KQIFgHhvgeCuRl5gfR9lwrkJOYzLl4Dtc3GGu/tBLcrfjOlbB4zZr
KzS2YNPwHs+sJXub7pkYVv7idd7BVBg6eM44PfjpbF3SMASlJ9jXZU6e8Ic0eR5/
0Y/72YDGZFIJF1ynU45v1DCxuzCWj2WxNsg3t8FJh5Bj+NjvCSi3z43CUQG2k3z0
AGCr8KzOEPK4//EtlbO/rwJzTq4H6IrXwvvq7WOE3RheTMqcDI6spGoE09WWVp00
3mxYu8uT6c0KJoaDdCKJZzyieHvY/8rsasJGcHzSDnZgnjDY7LzAFqkJWciU4ds2
LumPJhiFbHrOusJW0NV5MA+GqSYplhPAv/en72JXz+RHwr2mWICmsuMIbKMuhTHi
0AzjdVoa19j4dFLZXHd08V3DNnMrTiPFn7X8/oInMLcRArXGlHO7/k8ZMxHNWBGm
emKwXHvK1ilArQGKYbH8DazFfq5je7sXFUzRmr/mmB7kDiIV1zdsCHHNWPHkKkpH
pEuiOIsaHCWlnjqSfX3gPGAOR2pxqsEu1gJeKD3IuEMrMu71D6fAnE9p1fUGB29k
CcZtgoydIW9F4LLTyiG7GWFIF8CnneFiKESkWCRDPN08D2IoxwBItaSIAXMGuKZo
P/ZSFt6CDUcU32rJ+QdUQ8JOymlek6pRa5/xNv2U3G8IBY+yzdLNRQyH5muV7mds
uOmWlHPiXHPVi/JEplOcr4+py5OWG4tIVfrH8DNyzT6WSwMisZ6qm6XIvSlLzqUU
rnVmT7cfZ42cNjLOqy7Hsdqw6v5EQ3rXluXsa9BhbwpbvBJMATDaXoWmZRlLYxrx
8w6172mHExJWuqzOSJb5y8FjWihPtSvrRnxqhgYz/qhI70sVf/eeyV/wcF2NY5J0
fzMH0SseXE/CmF3X/jMEiY082uwzNSvPwUo+5bc6eSo3Bs7nUr2MstVbLT2NKoxx
leqRABRDbvOUHOVBUFPYemxWMrB4qwYZfxh1DKkB0vmhWoYqjG0NHw6jQYY/HwF8
fMRLTZxBqbgHT/6lKYei3xmN4nFRhB8DbGV0yLUbOuZt/5/lyKHUX4YPPs37Xutu
TlqtZjw1It6YQs1kw6HBZIYQ2xPj5nXepvUHqwT95wPkMfausxIAzu+F0TQLOU2W
y2wE1crasCg/oCcy+UIQCZtV25HdB7mcVhd2bcJabvUEB0y89Zx2Cg0uvMrCAf7K
0uBmXIZg+NJAnH0YqBQ0oTrfdYVplCbpuybQMq2JIfKiWfr7Tsstks6iyE7vWD6X
hm9x+HDGsLcPWsRxIb9MJFku1TIxo4eEeLK7+8BANImotCVnoraRXj3uJtudYlVM
n87yyrkoTG5Ce0V2IZT01Eqmtj6EJqBazre7kKDV0ZlxcoK9g9tUw8hPgS68kOYs
B5H2zUGAx1BUpoOhfGhErGH9USUsku59fV2vA5CPbKZMVIrHVJOlH7TmyX5nHq6s
9rMl5scPD8tXNzjCMb8WZuP3z+EZHM8TAkEfnKlqYrs1jw45OCTFV/HeBSjKXBd0
8nvCoQXLhsQofTNh9KT32Sw+2IhUyaTTY14kfXUuopyx/Je0RC9FT4Jb5BgrdkeQ
CQIH1ggBqz5CugjbSgPAHJx5DSbtyD7AIjJ1Ppz481D8rW9NXT+NZItV3ImvUFNI
L6lrjNzK4FW67uObFUYkGdvAF4DTZO/NUcAUYwCPdZEKnhRLMna1n+HKqWXvm0jS
tbdgZbO1uo9R2DnUA341rPSNA5tE6Q4kp6EObiR2WxT3MhPatJMifjDhZbnn1QP2
v0SxkvOBa3vtpuKuggEWi8ZT2+Uy0+vQ/+UQegWnuVxxniQk24k0X07LokAHY02H
tUmtdVaqUGqZZ6f2l/YBNsCd33fxF9M8olR0pSnXAa3+Ci1GzCf2gdVqdPm7MD+s
0MYwe2lrOxjcGY1NCdi5qiQj232Xq66N4FkJM/4cQxl/ZJR1Ww/SVCVmcnlyq92W
Q64XrzyZBG4lqvgQnBggAWJ+CxSA4VPJ2eaWllp+LLO/3RCn9lvXb/56xrZatdBq
+Osc/zIS535QoikAV1G7DXhlklcdaiNuZk69NVPDyEhXf+59ZFUaY/H2UyejZWSw
ty0PIYXxWQHg69F5kgzFICTeOTNpzUkbfJZ1kcCyMbW041pGdiwQFEomKKl6p1+/
8cztesrTi0FqYRfSX3FT8NYAfU8YyYJ7Zi32aYHAo22lgHOCCxoHDrrOPibGX0SH
RTO+PGnIT5NHZF0WwKjeIeNofsA87En/gD6G/ROt9bGLZBAgYrCGqsXKK7uOdIwn
PbIwqzdASQuTCeeLJZd2yqpEdLlkcI6kvRS4j5CjYXlELk0AE0LRN5n/okWeQCWV
VP5wUONkd9r22EPucIEpbREkYrTpeYjFVeEix8BJqlIFWzZq7qyvMNjAoB8iDKK5
AEJWJvOwe2UhICk+csKT1YeuwTbLPx7mr4wazX+o3sJ2i/GRtcHu/yXttw0AE2Nx
r3YMMg3hsVDXeY8EFjBeXMlo9x6fC3WIYsuh65t79OqcKQVd0LeByx/zQmrnuhmm
ATKTUVjBpu2fLOZTRkF0md1FXezKke6l5b1K/u13CKWGFBca6QnXMKGzT+77HAW+
ARaPcfK+Lciok24p3XYR+Fz87ITdRemdwLqxtr8h1Qz6/3c3IXI4EnlXXQbeALkn
rfCr2Hqyy1HN9YbTO2/UseKs8mGNTyzQCuLDkOJX2eIL7digRNqKRBV3UX4cuKNQ
5bSf+LfNN/FgJ3qnzRTSbT2TeAyPtsjuOhyD6X8LTbHi6U8/1sa7ymIsqAUgL08s
u0pHq0w07KjqA6YezEkYwWAkl48WM8gmFMlc0DSCKXM5kdGND9zoQuO1ix2JHtGG
lqGoDJ7xRRIyFXpt3EqvL8gPh3+jodm4jSsyIudz2/KBJojKfx23u8bQ3DhRyl7w
Ub3+huR16UNXWYHILO3b/ngMmDbvOHSkEo+9sXnoJyEFk8t9UPJZ9tOjAvcjAJHx
SZbQuBkUwxwGrFkpMBIQRKkH24NxetZO3LPNLsOAUfQ3fTh0ePMdZrpwpwBvYePa
q5mlhlBHKEi/L+a27k5RiNu/4TrlnRKywY2AYjRa78Wnxj/z6+JPAmCLZs4hkh5l
ALzxoDze2HA7hs1u7nvBQpdSUIACjDTs9+fpLBt1XDAZybxP+k9KnfvQkKAvxhwN
/E19z6wXrLmaNSt8xv1sF/otsX0MrZ7dMDcdwFgmfmNS9l32HmfMxefbuVmgcTbx
c5IwVcgWu+FJ7xen6/B8vL+Y5DxYh2Xk6IH5ioPgkSQyJtrrCxxM5wzluoSga3Bu
jhYXCIn87+gr+fwRBlp2vNLmcq9tm6jeobGqDkwvEUcoItJakFQ0DwvNEWtZc3it
OT2nij1gfwx4ItaE0IM3klooPUdqBqMDuA9oepttUaoXRtNySi6tcBcA/j/S98Ul
evQRqBc40ce9YlgCOo5lDRH7jisarNigvxlKtrrvCdP+Aujeose0HNAoQs3gPt9L
2vg3q1gOl11TFc9blxUvJIit1KE276m2rjAmwaGfTejA8UZzcLK3ogYhMx7+19Fm
quAnlh0ZHFt0NLzBmX2+3DTeZ7IKonHBHnUw01qxIuoZXCmfEIHc4G7n1BkvClLr
mt31CPZ3O2w/iVc5uY5lwdv94PvWqLLQLivTjPcigzuFjONPhFU6Bfjwwe1ODUEh
YqjeWlag9VSKhWedK0bfzgR7yFLhfl+vw4tDkQi4yN7qovk6L7OnT+bBHnU8PS3Q
DIgMbJRbe/xR28FWNzQ8T02r0upXUepspEyNvr/+o32kNZFI8GgR5vphhwbVDtfi
C7Ho5NYUUG9H4x56uo2q11wtmSdNtF5Ud5k1Tr7lb2ZZtrG3J8pkNvqqo8d3CKTU
uzEu8BIMofvcvMvn5tR2/yXoRzGVXOs5y0R/2dUmhrpjSRTN/4iA2VDLHMujD/gW
vy5BjoidH1WSWAOM/7LTJ5Vpw7gK++ACnLnWWJ2RcNnbBDq2ObWp27OFr6m8Iy+a
KN96J8G2+ILm1j/iqO7r9vVVT0QWM8rmYYRSJvxD4rKcee/9iYN3AmCG4pxj6ol+
Hhmd/+/r0VjvZuF0aihQeKqTsoPhjroCJbvWs3tZjRtzB2sMA/M6pNyL3sjw8x25
0aOaHVDnc+z9ZJeSZzKJC7xe7sfQXmPy3vcb6DAgc/Umbj1sqcce5DoBYWDjlyWK
yznJ+DzbYwqVi+3ZnmOMVx0Zd3nVQ1ht/Nk00t8JX0c825fy6naHDL6r2cw1vvhN
qmB6+lvZtyphEXGeiVEg2TxczRD8gBHcKJnQW3E6jDc6F1sYC01L95172w2PaAyD
GjgClAYonSV66pbs4pod/A/1zFp8+E+lmoQoSdP2nwoRUQbjYg0QsKx2ShtKBvkX
rxzo+giujpIF9wyQnGWKddhVYCVmF5HSxcn3kRXI4IIT7KUtfHNf5hFix9MzmP93
5hZcbaO6aQrbNF/bKswTUIj5mACXlFWDWGu+slUQPcZGp7Old87TvwCWVlusM/Rr
0yEFFWpCbnjoH3i7WhyaMtUlGkFK76PHaQLZhAme5WivHvwPWzzy8PeIBbRkigN2
Sdnm34iyJum9PlGjo5SBRCJnAnBLYVWvAMnMFTTODa2jpqa2692CYWtRH8WHm1rT
Y496HhcFudXBqwA/ZuxqWhwCZwA4pCy+O9hi/RIa+PNd5/Z/q5giJuMilk/J5SPX
mx+QAhdhM/Skn/Cpt1z1kCVz2frgz2hdO5vBktoQA5BN1J1v0/d9EGNT70S0Eena
mQnTH4s+n7MgTT1yhx5quQv/mRUyC3gu4vMoxvo/WS6Gqt/oS9J1wF5dpZXV7wE0
FnR0Fq1fIEMZZYJfV+kyHxeaZstg9FOQTP8lhQYQW035HbWz/U8ES7H/uCTEYCj1
8JJH1HDqO5CaND37VODbq+aDFQ1Nkb545uGA6LCElk7ZhTRAx1GWXHA5Hwt/1buw
HVrmlrOCzBk92hLpWPt2LP5xzq0tZrHH3BHZT8jGOa5mA07TLbi+FnjTPhWSgAAa
opmX8rOcPmiPmdn/XxvvANAecdELPxZcranur+nKu9GkSg1t0eYvt0W8W3iyf7cg
/CMK3vQjpJA8lgcqntIfLibT6K7t+4NtS2ontxsoorBWCdb11zf5JfgNxDoX9odO
+6FFM23NQOJn10q/Pw0Z+n3/Nw+FIDZZAHKLigyjSk1bKojhqnwzoHkHmdeF/z2y
qGp3I99UfqsaX0PXsbg60nQc/nSp0Keh5TuSv4S4E7vLkY91ehvHEFfDsdN88vGl
9myvohpVwFyKXOYtnEUyGmQykLjgCUHeCChjvyCLT5pgFzsDo2U/hLEQNcTWhc8k
AgX85KDk13zU3cuMjgycUF3LvA+UM0Y9FqK8BRYJv8PxtgXUWT7DF0Xs56oetrUu
Jp8PvewFn8MuL6YpZTxCuNryRo4C7J8245WSM0cjHI5L2TR1C54Qp3KurQjPCZ2N
2RdA2XReb9JsBfOGTZhIqFEEiN6SgpcM4M8xHQZ70bab18MCfnTGIdfHpCQcVmO+
3ndg4c+M/VLBNfr+Hl+5/4catWGgg+FQHF+A+L7g/0mfVEHTslWZXNFiK7K9rWDH
qRaOc4ON5XsHsKHLL2Xrecfpz1k4/otvMWGgPnX0PNZGLrynXvGyG99OSFA3h0at
yBLvVbRyLpQljcxKfzCR/AZy2WMN0e7LErqC3Y2Xaqp6T8vzwvPEeP+dwwBOncfE
sSvyHoczKqzGDaqj7aqSrZqb63cl0NLWbFlskNWnqrQIK/HpCTwqDuxjjuwaT8dQ
aBPRpgy1dpXTeyo8N2hdFw6dwzIjWw/gJ7+2xcQ185SeOodid21mSzihK0K8F6Cp
HYyRRZdRyXkpyMmdvqQCz63aKJTK0N/ytbozzsg3kOSV6WpwIt9bKVXRkkyRhM2l
7yZeVHOd3xmU+0ElfKo3xpQpO4tjqFgwofgRLmb1aOsC9V7WGc4Vnxg8l/wx9Gut
ULWeqB1rPluvBfaQJI3kF0/Su2RrzXQ47rNk3c48SRwG/DUOKl3rrzonckTrv+BO
9v9Ffuf3knGKkk7YG2cE61r+ovX6sAxAzL+uXQYvDhKcNentkvagEWP0o97ZETYI
f5PBdcsQ/qPKq72s2T8ASHz5UmiPG5grEQje/y6hq6DcH2tJYVKdBiV0+kOpfO0O
WmhMJwniMonfTDLNpXBzmRZJKjJegK0xXOxuAxNPYvk7xw0+8V5zSmKhWuCaqggZ
6ZzkT38Wlv2PfK0KLJ8L7rag4SpTILF9ChhXD5cTA1GcFsI+2cX0sKbUDwW1P3Py
vIhcEhwoiX767E0Tkyx6IOVWEvmrUvyIYSx5wrMqYzUGYAlWsG+ci04/Xc9qOiso
1twWVfAEgdhnrEQQl3xbjTHE4WfAN1+Uxdxp+lJRQiw9Ffkmqy2w5BaXWBnK9QgJ
1AYxpgwwGPWdJJSRsJbz/g5sy35Ciug5ch+XG/srtZG8An2Iklr/oTkeRQkGcSTr
q9DxPeHm7tZZZSoNfHjtnNFlwSsvWRM/pmBP3ciaVbCOCRn/N1OT1e8BwvpI/U9r
SpwyFpSDObhSMZUt3d0vcU3gYLE1l31PbFlRfvmFuzu2ReaCfv7mOD97+Krcw0Mf
ez7TjcD6GpbFTwSD7pwQRneHecGKM6QUeCzUsnkw4FD+frxD14kthX0bMdiGQfCo
eW7Ow2ESj3IizecQWHt0Yp4rjdB3eD2UGdNtcImRV9rI9a9UnJBma/1K2mshax4z
umQ0uFhTobSFcEpvYqzeRxGGubh7OyhJdEQI2ISJWfkYXvRt7C1Adj5L37tE7V/Z
732A21xR5C0EHRw+OfAOE1sTTYJcPPShclvcErXp73gXRWFN6yrpM0aUFPGCJcmz
Q6B4DLGu1kI3JgqflWuLMs+96gku7Gds4SE37TO0tZFQltUtjogJQqZZUQL5hZmY
wQ93N2c15ZBCkBXi0o2cJC+cmwG5a+8V50c4ev9JOKLDDcSccaNcE+0Z8mesjzyX
8RY5P+I/QRPgVa07g9ISDimlmuQ+oFaPEth0AKTcdV+Qa0pXR1o5Yx+HG2PuhDWz
OH+9UL16vIBAIx5t8DcfEZxUqu9CsFiRX/ubZ6/uJdiklfe/hPNnP31P0R1f3b1r
Q7dvZH8eMdWB4J58Y+vTDm6L5WuzbO9izymn7L5LPSh51i/sa4AN0qSHyVueHCFE
dEKeqDFKCM0PCzWW/m4zP9MQKnzEmpJRgv/jtTYSuO6UNSLOt70FCWqvqho0CatN
AK4hFqpf9fUsSCvXuDuAkH6VSVJ3EgRr9nL9aifbKCXcxLSKpV57j6cL6AaqG2Tg
xVZJiG6XiTjH6ENlml3ti/LtwMuTq+48uLaqyI+8FBw09mKxQBmEqEPSA+vFkn+T
G+PD1nE2O1R1NHufrjTH4aZ4VqJ1ZLzTCtUFz/o8an8pYDIAjhmqCKviUHVPqGJv
QcEhPbkrxNvOce2EGQQpP7hs0ni2muoAo43APUA3EEShc5nudyyIbuFQNMiCz0io
KK9rmMD7xGpzohgUdBkFn39A+ALIzuqIvNCBgSlMs3cqzx+VSfIf9wK076Q7WZ2a
s42mGjApifErTc7P1td86WAWo08QODlXc2vZn28JXzRLDcd6V3xiPuZHad0zEPRV
lPr3HzT/gfj8m/liStq7PgAS5bJWj/F88LBQcYuTc/WWmcvPlxtnza9++hao1FgJ
ZwVrz5QISu6Kv2iXci6iI6a11FxJsA3KCM+go/Boidx1RSd+vUKDDbl1eRwHAXN3
HpciTbEmea3cD3ZqTqGqQKH6xeqHMTqLyrl8/AtO4X+EfzAdeMZllzIq+/PmAN/J
kfe4z/LdE06LUX4ajloMeNM9UNddhFHQ1yjwOAHpXZenFq11WVqyXIjH7cKwRXST
HzZ4NtRvxyVDz0cVL1aTQxU7p//oQc3QrFhzrRCQRKaSrgpiun8fF70pqYoxEIiS
J4oXCB/7sKlKV1TiS9ff5jgQzRRmXzH5CMzp3sSFYMjfCBPyALo2E2VprSpRBNMR
6uJWHBMwPD7NfGbwsl3LHqb2EfcDSdR7rAYit3tqKybuqVWfsSCEsnXYL0DeVTeu
pnAoYEUyg9t9pm+n5O6AktD+Hct5FUno/pUPbFm2LOBdyqT2M67aqPe99zp/LaGN
w/L+8cAPj+K+u16BySMwjZ/905PngMcDzEJY9hZ+mvVZLiQTxaHuFqMsPsI/fGb+
qAOUc0dnX7PVrY97BncxzG9v1qVBlOMWNT5EEm3Nry7hzqJZ5Knoexoj3gUMrg6N
YP8G2lkBmtU5ythUg6mo0g09TaoKYWx2VCE/Efj1LvLZCJ3CcYgDOJ1z8DRVVjF5
FeNmqUVEcEhrgp+Sam6WqPHlp+73zfIpv5J0SZIJG0wikl2CzFx0NAkLO4ICBaHx
6POpPD5buJiJcZOJbKFd2L4q6+J2yfG0oPaE2N+3u0e1dOHR4iXwnurqgvzGF/DQ
gvM6RkJE2reA2nbYuSFVp6r+2kWVddS8FEZ5aNtwlDn5mgOExWFa19+LBug3D8py
SvZwe3CLfP/8Lh3sJoq9EL20osP3AFoNRWgrKqgkdLRoB0mfCmWGYo5DOghkixQb
w3Ht/EeisFkaZd8HDNgmmJAdtg957NjuBEZYeJabLb0cWRlZufJ6WFyXNaJDu3Nw
V4izbLKXWjL68B/eZE+WtHOa3Np2KP9ulQoKGXrs7CDvvNww1uGRClohJ7D+Nm0X
5LQWOy09ZNDlPY5PoxepXfeyrDZLEucCZXsNKJlTUjeq0GrUzxpbK1Tfd+Et0D20
CJPwc6o0OqJ36H12paR5moTb++v1lv+Ihfr3WDOHgt8LBnY7J5Hr0IuIHfFqpj0+
mrtccM/6Fq9ivV4JRI3p6UF+0JezmvvK9eQ8XiELw+N18+eGWjpafpU0cR5npA7t
4Bzz9d2SvV+wDr3jW16gsdT+n4AkdxClahunjqiZqgHqjOlyjUL8E/l7oEXIywCo
M6tt1VUOdR0YIINbd9Ik61zVL6CjjJAD/5BkJUtyHQcaXiK20OjlBgIxOi2t/HeL
2nsYRUkI0ihGBkl4wY8dyUjvkCPmPmhrdwRnoprJW9li8d0WH3aGRhU3vQIjavDM
m0Q62EzGYldiwz6RaPOlaFj9u8Pdv8M5dfB8fEonBB2RSIEYyqfZEbwL1b93Lva2
Q2NLIwflI0kNCqNTqWBF8zbaVn3PrdEdOcXuv3hwFKndTMx8/Fn4sMqEtFcMRXIo
aisUrZs5fZxCR/Noqm1eP48r0mlwo3GvParxaiuwSFSmHub8PjpAQTT4W9rTjnEW
OxylOsl98XzD7g3HOuIw4PYTNDZqKwA6x5YmS3RV0JIso1/KaHzctF6poc9my6o+
R50XkF9Vn2BFjatC03ZapB2loVzFUPFvqXASZcWwv4GAowIr4U5hpuADepQFs9IO
FwGU6HFmas9bQTJm0Z36WbMA8cmatoR1PVNV02eu4iyjip2EksOvfYEPTgCXQN9P
vrAP+UC0dTR4Efzd7fchDFsCg22h/MDFLufa8B7RnT3scKFLFCM/l6KheRwNbUYL
cmHUUa2SEy+sWSt34VSyrIaHeJudg75fuANltdP330Qi0KU0f1gg36iLHE6dg1wn
cK46pq2FYSzrneq0+1D4li3XSiT/CYO8NXIMeWSQgOx+WWFh4vS84rpJ0qcbn6OI
hTfK1LXdjQECTDdyv5qQJ6ufUg4Ttq6uom6Y3BHx5iQzoPK82c9REJFGlYfz4CCt
zvfzZVvZEvIAbyIFsfEY1cCrku+1qR5972TQLSYNeQkTNHQKBGC/3wHTQIQbIJT5
86Txzj0gjRUE10jkZhQ/Yt7cjUJaqyfGsQRuD7g9aepkMdF5hpvXq4elVQ7hg7q1
IXRHfmghC49MStjSVY+ovvd6YVTvou9Y0KhGHR1R+1/1AVLKwEck/FuFWjxnSbky
ccAfIxch2aESZUbqmqXoC5Fmx3+Ej9EKgv3lrcP1Jnzf9pKa/r4RQqA14bmjpck2
l/DeIO6WbJiAugQiB6Tyz89RI7upW8+K7N7bhswkcvWoo+r+g4dFfdjJMcsrXgS5
56YERi2DPuY8Gp3OgzCn5qV09nC3DHYzizKEKzmjFKUwgFZ3RX6+WCKStv1pC/xG
MvsDhn2sLaO9xK7twnoT4Yj3SJ/SwwsdX8i88FOq5Ohmmq+6q55N/mGyZWuIcTom
WyUL8Bw7OTU6bvCJFwoobPUwPoMqt3HlCSaxJSH+INofeor0iCvBirP9Fd5WjivP
5OBtaEDzRsHLVHD7kV8OEgPkpZ9bOWMh/CWFvfraPmw/NQWLVvBsmpCOl7em47qI
PG64e58OyShScyQg+L1NDk+vEZGJr1pNEHu0IUjcJjom3tYx2EEcsmzD+X3+uH9p
NDNtZ7XivA2VjbHJmy8/54qToXRxrfjODF53lQjvIezNwZKgHaKDT+V8l51Pv4Hu
pG6qfZ8gtSqNEIhGBOxymy1qfGTUr4jYeFrhXttGuS//tk9vtkb06pwOnDpMqGq4
0ip6Uf1+vNIc0TbK5Z3ng1gndIa1erEXALM6kNDSJPFqJqt88yL4U630sqJdKnYt
ELKEb1Htjwc8OaJoRFYg2+LJr3DnmW7oXbc4F+90NdKogsLhH7ll+pyUT/ncpqQa
CEI2moPz9AeOXqNmBRRz3maKbsploSNuhZ+AqbaypqS1WjGMbFYt1/dKPXftBG5g
r/PPv0hp+gfpSbrlJ48re67pAo6XStUvobE8V+hklWM7w80L1ltHO50stuCAKB3z
xnYaY9egDBvs/ZguaeXUk1gRPJKxYAQoW6Abwuz4z5ko3QIyz9UpO468vAQjr5Jp
IT/MrywXhKRwqp5tLll8T1qbgZ+1zbExqd015HkssUMaCu1v8cAXzK+yX4k6DtZh
B5mQGGo7XxksoEu8F2BvzLaQSy/GVG8kgH0z+phqGjNWPRmkgXH9JHoZdX5jgwud
zQfzH51PCRFr9UV05Ao+7rSgcPBmYpoCqw+aM4Zbgzg8eYVnyDZprrC2CQ9k8f0r
8fX09nEVlXG3r1AwvViYMT6lqsvAUBK6Ajo1HKh+2wxhkPO1dziIrcNIqwrkAE+o
ve2xjUyIsCwSSq+lg+7HS1s0FtXIZRwy8nAV1lfNBif6K1UzTfBLGgzRm8dmXwLh
dw2Ai4qv5+nFdDZKB3hMRvsbA5qfP2/piUjDMLzu98Kp85U2XJP4pWTtiE0DpMya
V+kwLM+rYdZmGzxZBjprCxK+tmRI5XwgDuI1GKRt5n23N15rFhuuyRzIKYfjxiKQ
7sdrNMeFO2rGCDlmkVLkFeWw0/VWohw1cgdX/qVeB8iMkDpE+9hNkEOphVap2X6l
eO1P4cXlK+pU4xOgZD4BSlury70nQ2rEO2Gzmx4RPlD/r1lS/0XL9ecphc2S89mQ
Y8mog8yIxTa8DbrVxPd8+9K+ahEY1nr2ygsjCH9SYxVeax7vqx9rB/L5u978YcjS
FstRGh6uMf3MdboQ0YMwo4In88rDM2QR42GQidJsZdP7oonIlgYFVpm2plQbeWXA
RsFChs/HN4kWAN+mJyaGV50WDLyySSA66Obj80TSjRpAipzyXlwGmoe5RBdmS03w
/TZinSmMGl//Iy4xxJ6Q/B0b7IxYoc6DAsft2/gt0StE0VuFIVD54AaVfkCsBJlb
TsTWd2K+CCaJKPdsz9xiRoTOSPXv8aujh4flRNBUQBIjXUg52bu6jb590pqjDt9Z
WjjOJJm/ELozO7kT9WNe4XK00DMFPSaQopHUtnRhaekiMNGb+oX78xh4UjUnsnBk
ijLNWxX95ZN22bUWPe19HQ8S+chUsBp61Vj+m0soleFsdUR4cCNZxrsr6aXpBUy7
/Pg07tdkW/3cqUVobvDjhdHx0x7JdN4skeEDv51z77kAfn4AfQVvCNS8IAE8/qAB
0ZKuGBK+n7F/wj4DM8DaNC/uSCPlcX5TUDlkisBCbHHa9uiMgULnVlYvvnpmfHPc
mHc8zErW2IKfGjZen1jFeW8vfnsmlj0vPh8pY6hGWghpFauhM+a/K7Od+IjsXi18
iGzMKMyBCGBw6m9GluU198gQ0e1uDSfdASJ3QEY5o9w3aFAcDtpFwQ1zelMd4TL3
B+B0IHNetQOAiw25ri1oHzfGFHYJvSylyoozh4NLrAsfImokVhCeYWbtYArbymlU
HNwG3mZ9OzlyUdPJHOdW2M/jk/rpD7oTp/QX5cqF+O7k6Rg0wynvdl5KBxOtVRwe
e9GPVkGPqVCt4aaQ3EKHg5girnisk4oimn7lg62d85vOfO3WYQq5zhUt898YRyu0
uVRo+MA45C4C1R/q6nDX6XWB5OsvxE2dLYFCXJqnqIh/Jp/M1zQpgmn4UUnddVpq
fmlK7km1/lD4eFoE50arST2PI8hxsRB/WJtTNMkn8WEHPsCIzs+9ZHakexGdtjLd
2X93W49slvvAyuO+QRGs7TIKNH6kx4OJO3UFlJlhhpaJObWsEVQfMrYNq4b2XdFh
rHAq3DOlDjjXik+BL6xG8tEA8xuMNlmOwnp8OtwIJAYVkWohye8x/VSA7+LeBk5p
/gogV7zjNvVpCGvYRpjtw7SJN7nQTjZrNOx11GTbnwLHfnw17VwKX9MZeapKs3nl
a3E4BLEilOWp2o230vNbPGo5F0wItYjuuDajhaRyyEdwe+J0W/Ptb1yS9KaQRMNi
d9C4JJTgzdAIQUcV0rpAumCk6Bgwrj1SCqEo/e1+kNu8ZgvPsHFcbxvBegGMc0yV
4oMT6VxPTFJNToeq9Mc4YYidTTEQq3pw0IGy4KTxisy+gkAxcZkvI4CtTkSu9kCE
a/bxJcg4XVt7RWaAOGF6xA==
`protect END_PROTECTED
