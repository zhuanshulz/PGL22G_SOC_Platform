library verilog;
use verilog.vl_types.all;
entity GTP_KEYRAM is
    port(
        ERASE_KEY_N     : in     vl_logic
    );
end GTP_KEYRAM;
