`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CpV2+Lp3j6a1seDGlf49PGRpRwJ4nCNYobdkvvavXi5yHqWHv0EF3z5kdKsCJcHJ
SZhq6Q4UHPZhByNpgVluiP1EhA5eVFZYuWLbKGv67lU5iDRt6LRn6ILPiRQVasEp
Pt9gJnfhZyvY82LSIl4EVP5ivqZLoz4exirezzTuFYBugYnYLxAKNlUh6QdEpNo9
Xl32XDIZMVgTLvvR6115nIu0d36lWAhT1KjiwJPdkq1Xpo7mRurIWiTNRIeMFkOH
ojf7oNqFiULLNkph1kxXbtQvgLYArt8f817+8v6KaFkhpHXvV0fqCckKkPZFEjRW
26zn77hvGV1Yyi9apoejyh4ZeW74SUwrO6Js9pfUTyQX4FL2gon8TKT6meF639Sc
L+AIVbM0R26JDOoU3j2x2IMgawNF74mWg07YxuJJ6RpdG6J3I1V2OLMGxFc2Qwmf
6gxSx6VdH0H/yMC0mDvleCwcCikJ9zpgULUISKD6Di8I7dl7cm/IL8/pKRw9CVrW
Gibv6OYRquBp2Gj4jbW+CXtSf2LqR7hIz43i7b7Y0ozJG+ffIUdQna5gV0rawSGk
XMRjIZZDKp1p2WhuidwUp1lAFme9W+k3rHsY8VTVg/c65CRhqZhOWxOuA+zb5W6+
k+1PXDwWWLeLE21F5Zven2q3yiEP1JSwF2GmxtaYApCeG6jB+JOu1TlUahj4r7tw
bYetuRBR5yBP/3g6DAh3uFOwaOoTS4hN9bzCNhGoaRLqQoFdpdAqtaDjNGv/s8aD
nODyHuUH13pRRwqM/POCnUJNtvGV07vNEQQxc6wolps/UlqqRBkEbVMNNIoEJjV6
03Ro2zv4zpjbqfZ4NXxAwvydN74M6LuyXH5vpidB9YvCeux+q9WCCTxDijZEWS6A
xaQ6Y03Q5uG9nYPHBqSA2av/QwBiV8JQK8VmqWAYCLa8IHDRuzGqtLgtVLh7fSOg
B+PFj/RUH6qz3KAx7gPMQxwx/DevlOPddnO8Ri+FNas8aQZmqsKc46h708hVnQMI
fMf58TTc+1F4Ux3y0tqkukLH8qRJJa1+jDZDXrsB/7LBU6kApl9PyH0wmRYruxhk
IJwx1tYG2PHcHVB4e/TejOyu+pZ3+f8CBZjBuHUYt4sR8BvllX5Idk/DMhRl5i7/
azjx6FMQmxpyclQSCe55RmZF4d87g44RVJHwXg5bE3kBcIOqaAwyrVvzx0kiVU6F
zq4rYMdyxYlLiSYc0dYS9KxSJNE5KQ6IjljROnR6Tndu4EWS3bGYFGSlJ03AdqV7
UOfwXimpjBBKkJsy13A5EW5B2nxyX77MVYzV8cVveLBmMkCPKS1FMxPh1WaQKtT4
4vOlMyOUvY1cFTsmcjPJWKr5e1qAt7cub/10GnTcvbDl6NMBFJlgiDud9f4tgA7z
X0TIKqvSd7VA4hMuimuTClUO7cGPEbN2KgfNwQxPZ5SinJtJoQhEc7JDwffsuyGW
CSMb5EMBmSzVc41fgU7T3Vojv6fOQxWn2xkiJk4wik549bTgRirkBpExQaSIqvuH
oof3jcx3ghhyiXXEyg6rz72ZCRSefkLQMFtVDYOC69kkui+IYGImhtWONo1MBR8v
EZR7vAHo3hacsUS4j/J0dmbITQqHSBOXw8RK5zY12WSgF1dTrMYZzHTVkPCly/Dr
3xE/t6X56MglNLDrcXUXKRtJ3Kfn1ugo5H0BXxNxAwXLNwCiZqnKQMsD9DsfvpZk
hvBiTTe9e5W0bj6gv0NaM06mZUmz8qsSO/MrbSsyfwRRqIVeoT030qnvQctPQzsX
qn+H/2QO99VkXp8w7K5QgfS4l7nqP8vblUtnWbqmcqOlGFX/uiN6YbhstfABgEXx
mXcnEEhZpB6IRjeU+7CDSnShkhqR6hukzjH2YwjCmTKFVFwhxNQQjDAufNOPus0o
waRC56xe9dG6whdsN93NePea/WyleX821rHflFsF70oLPAbnT3waWrNrfKGqfkYg
E4qK6sCoGDLeBnz6lNuJOFOnfvbgaMN67PuKQgeiybmk5tUbDNjPYTZqRnf7191w
L48XNvbHBtK8WpZYX4Aeq4ln581fg5Q4uH+bXIlCE/YGU79i/vPCMr8vMKi+11Bt
PqvTfUvZwNEXmB/DefGZophgrgbjk17s7+LFQpRRhqLkVvcUp/ncvr/c0Ygzowrv
8drFiluVw6LrdnQv4+SwNeFPtZbglqifQR2+HU/MWWAFESxKRsXN2Dc1FMchjdQT
3YdUq/a+grk3cuLtUcOWFBhnbOz7XZRwAZy9Iuy1OGFM21MUoGZzwu0oOjOku28a
Wsqy/CiVmdHk2FAnQpsTzZ9eX57IoA7hIW+oPtDVGll00xbCrGWHxQwlQqlP98ub
qXUblUNELD33Ajv9iQYrhVKpjvF8bgWETKzlFvfCgV1CIx7I7yaLPm8fBVf3t9KB
BDxeONe8qUwNNvwVJuHx9g7sm2Ec7Lsls4YkEHM8R6EdGQLQ0L916xzlvUVClmzm
0nYmwr7TseJWII8+20jcwIhvT3fSWUhl8ium+X/ALO9P+33aQLlfZXJ8NwCTF7ui
HYTsYUZhLFUw17CiYbCuev7NQ7yRN+LcoSerBGahJKFmI00c4x6QJfZo0Kf5Thnr
52EwAUjO18Ce4XuffOG1e7fsq6ua0cGuiNy/Ngi3IvhY5WN1FXp4sEQWI8ZNdICl
5/IEPJsjz1kY742P1NQqqI9I/fpOCJdKyQ5BxFhBUTjGd/0ous2ZB/OP4nr+ewiy
tfRCkPOYJ/zNX/V8UVKhQjKreF6P4sdIQ26wPYEJvAytG+KRShIwiAZ184sLyto+
+93esYyCi1bsjDZRJr7i5Rjm+rBL4tGub3TXhk6vJ+CtMGJkQ0XSNAsiyj/1fKPx
rN2oqqjssQkGkH1YkwjMZcFU474wZXU5TOAsv2gmYorL2z/Jvbcuffvcgej31AaX
uLDotmLbDNZ9L88HIRN7dogiSNSD5fwdbO2/FVQRY9nm+MELCxfLc72uyY1y03ok
KEYmfIKh4UnGCxNFY/9OQ7OyFbmBEKv+E/i8qyhkm12HDCqoaHT6YLmGa4N0Oe13
lPhFFCZ8NIkLddSmH0QoaW3ns9rvPvHbbUoZZjuuUNi7y0s77a8f9SIt7VIIgO7C
j8L6ukTdCTXNZQu+yI9D2yn3romT3aQxthsts9dar9ioHDDb0fxHJxv7HajbX90T
010phhF6waivXzfNnEB6GHyhWSGRF3wdNDDYnhoj8nN0nAAU4sEV1QVOTupNt/l1
n02T6wsie6L4R6Ut1z67/q/ZiwywMPNaUJQS4tqrRlaUtxyTPWRaTR/MnvW2RSvw
84TtqVl3G/NXiUb4kRWR598Kw6/h6+n+IEv0Noho/BdSrJwRS9mnQzCq83UY23Vv
6WNfWGcnysqbTTbPErajDDkbeMDo8gVt8T0QX6t1NFpK0QF6mjZ4MBvyLMaJGPVL
UEZGiIhoMkEuJ1V4Jj+73OjPxqCM68TPxbSe0jxiz38JQ3VSLaeSM0LbOcHmtGsH
V4T5vfz4qC5g2n+atEMfaD8JRyfGxkWhxMnBOqSupRjhMa0fLnDi50eQe4+YWyGl
f1KCcJaFlV2+p4tWcXNbcgPdD6213BFuaajun07QoMxKD14K9dei56Rqo4t/AwYj
T4HPPZ+DMXbIUCbOJVhXbCAtB08pTADwmjgbFGQjPMh0dFzIqPwmOYL82KW6Ueui
Vm3I/GT6yB+R0XT7g/HYDNMGs7Yeqqd6jiCU5e2QDX1LIqgfMR1/Jjhrspfurg8U
K+pqf1Pzfl4vsWoB8UQ6xnRqAtrWa47aKrTK392z2NvZRFGWfZvbPkdpbnLjmWBE
mx7Mbsm2cXWxcewhickr1sTFqegjSock9Sho0hJPA8X0BGJi6SukLr93ujN4SrTc
wLq8qF7DpkEwtkMfqA+lGoT7aN5aBpyspgt1BlQZscE7Q03vuWu+8hEe7NMhHRol
wiWqkREO5aAcTvOFHxOz8OWQ1vw2V1ETX6Q9kSrwT/9ycmncMzHvEftkOuY5Z81g
pajAoSmoCNfIlMjfARjf052kO/z3YW2Eqn+gH83oskhfLsCoQU4GaI5DRCYG+m92
MgKzhil+cRbY9mW05raXNgaTiJUBhqGBpxam01ET6b7ma+HzrDtp/2+vp8hS/x/P
C128Dh8xDE5k5NF+dX7ssCJdcSmkqddXYu1AWhG6oECDZ9A3URCE7Uc14Oo0hTRj
7O590NU/GZ+9gRgAt+QsIMIDs4p300A0EbpGs6Q7bUrzLiRoSJ4/LxXhvuSvM+k2
AEYmXO5jS7DOuRRh2QgPSd8fbcbRFGi3aAuGgSdDtyXirBp3MNQrfR2LSm+BFA6k
M/bWHQEvpjq1JDQDhaO9euauSxv+M63MQ/c3WnzY07tZEWWOtq6wEOdIuxH1QkwU
F0UqIDK88yyXHy3tGRyPl37C++P1gx9myVauMlPaGAOi7Rpinr/ARlu1NU1C8KkN
vlCOkIP5TYFA6G/79JMWw59PW6CIzdchclAbOu6JcHP5Iugxkc+jwkNAPeeldkSK
BNVwSSgkTW3Vm8hxxpGWBVcpnL+fKjEov7UIAhh2D/MCIol5sG/2AzG1j07NDaG0
at9HQo+VrRDshcN0S8QpMyk1fhaVrpDLZIjoVaIgBjHu4NayXhUZgj4OU2OoVi7E
ygYnsAVTNEUGt22aYAvGR/iVSpr0xcfHbyzFbdFMaODBg7RUiUHZYekTft8r9wXu
bxpzSDFbrpx2WEvn9SpVwjpmLnNEZrurIg/WbNaWU4m2kg1aJ/yGfPl7qe0+jxZW
bxoTkzRq/CoebqU5WMyh1fuOFYCUigNQ6ys0v2pJNG9UBvixQlQgWX5zQvbdIMnE
u3j/XZhJzAPpOg240ehMconqqX4kNno1N7N/BdhGolUaKN1CykId2iM8EsjHxiyg
faOsVfreCGJvAeI5Hfb1MOBkkF5lNarHRXH0VswHdvXYU1FTcV9hyHWG2ivy9oGI
Ftmz7FogqS2INLK5cDmUjm9Dsm2Az7nsJbXyc3tvVz0Ml+3TgRJ5dHybE+n02ah8
L4qflNvErJ+GRhxjkiSFFw3npPbyrPeSivvu/F5UHWmK3udRoSRan46YV2Mj++ut
PqTFm/VF0hnY6Bq/fXs3r5Dd6MojlpiH65mWi+LI4QQgS+nmoXdMfED7Pc7OuWG8
xd2TISy4z1e0R+nGgvhG3qWdZHD68NfyoskwIB/GB80fjiTsx2WEVbFV0hitrjN3
CbcBi8SUasIkv9VX7lotH7cIXsxDlcK88ICvxNPEGXPCKR0eq5ENmtwoFgfxScvV
b3+bl+mTAl68J4Rlnc9wMLIg7W9kMbKtBCQu+YIzpAJq7FTrlHyTou+ms2UiJpl5
XK2e3bbAB8BqPrNu4kXBAoLqRotiqB3y5JEaq2/vpPK6bE2lHHkIDXGLjOX0XQgh
I+8ea3z4pU+LePiNt0TNXSaz5TUXrryUfAWIreVmqOLD+eks9HS6MCHC8QPqtZPu
CGeYWARcjohd1falm0dCLfhk/YyXtL73WRPQ48BM2IZYKYV45n+KHhk+QzUhVG1F
g81ywJZP9HIFChfqFZl3pr9SdAsPbxKRD+eA3ScT4qRgqfpRr//zuDxF+hMdEIRk
FVwkEHDqn5PmHbUBp/Jior1gSPJuVMTRUMRzQwv7IuavyMowuuPRAVOYVEqYqQkP
GO7SLKrRtrjuG6peaHNRaAR65K+cxw12AH4/dRE5K/tJhUSo3PRbzyuogp/8S4NL
k8yMqMhNE7ya/xDN6j4s2FF7B9wsIdWpKp+3plwePxM07gNzsjVvcYcOlMLkOdP8
ePXyWhdoyJs/ug/KtRr5G1bYtbexfBvioBoQDULlHVAiEkrWdeQHtPLdkabrQ6bk
FhMNxSi189XBXP2h++YvTyLCWbZU/+Pu10D/ZCxFVLoYsZCqm88sxOw29OPV3XXX
4MgAcsfve4nVM8Urjz70zVPmuH32JCoU83T8V66aBBvSzBVHpUMZZtxPy+1d6LV6
xCFURnnForq/uHHCNe3lTi38u5sVQ0CpP8cfQ1zQG9gDSh/ogy/ALS9Z8h4xHTJj
BDNmxyBdMrvPeu2rlor4YiWroqo47gVXQSUZk1ooUpJLhDUeetMkptNasqu3tdYK
jkc1Ms0WAWQLEBOyCeyiVsY+nOQMmNSFhtNCAqLupB+YroQI7jpoIQEOC/qb+VTX
7jKYURN3GQ/hJ78I0buPpMhKh4yuUfLJLs15aUS6sW20+W7QVsJtmPjAvaM4mvgZ
5cfQS+Adqu6QXyqETr6ScD5RrSB02ubS8EJtAQfIttkZxb/TEiAfmWeVBlrnGC+9
vKddRZEHx3bb5koSsZKWL09erb+0NRrlvqQE8/8yIVdFB/qh4OPFLzLP5BbuWyOj
1y8WImSoj3tOjn7BzECaWLHx8em4towy4506JijEKZGYfpW1SjGqqnpVtcK9fRPw
Ib47t5sTIpo5Vacz2bgFaNY8ZaIBkLprfIOhHKTHFkGZ/CvBOvwD0V0PngeBcxJ9
V37IduylkJoeM5KBQIdwCzg4psb7vGtm5JnmwHDPLHqxyBo/Fk6B1TvwK34geUM1
18V+HponWvMtlEhFZN4FFppZHkQyk0YRXec8kxzeyurY3p1mH/5tyCyQF4e/X32Y
4Mn6P8zG/0R368pdEHZQggtuj4Rr/+eOrO2AZc8ArgXIKwthu6FkcIzltkRJB5xt
HkXayFeBD9N6ceKLdDOwDZFb+/yTHZm4cAVsgQIkrWdr4DCXv+wBh1KVsckNqkM3
7OFkWjNsIO8e5Cla8smRhmwIOZ0gYSj5VBXIb6aazRrNVl0hhK3kHef8NeAoqxP2
6tLf0AH8mBB9F8hUTJB0TJA7dhZRIMpKzl0VK3AkTRrmFDiyEwB0Ah2a7ylHf4Mn
aRHt36+EjRrs0+TBOoDyq7G99bHmcZPmiFtpC//FYDveOQOyvwhigyoE3OpDHB56
YioFw54OcwddaSf0sWKABFKSIIbG4KM5ovFJZzHJ3Fod9GIfbIgmvBNJay7wqwoq
1g5WyA7d/DHQCM8Qp9oRqXRbkS70Yx6SNyCjOxisgzpuu48gAq4PVqSejDUZV20K
nTB/rcXUqN6vze2YzmH3Z6QukGj2IaenvdEfd3yN1ztYOhN5zR9+j6ui/+YTks58
KP2owPWqGcckyHx2UJsP/nh48hCz+h4lkVUY+wXIikRr/HMhuWjLl1wdK7x5PD2A
2hfCQlcTv7+V4AEI5ALN6/6F+ah31WZYY1ciTlELY2N7ouChDIyL+gzj9X4FMRXX
BmodIm6nYLN0veB+GJCx4lOakWOcj77pPKN9v+Dvhq4YYcTavjp6PgRmIzBx70/c
+7uwf5CzDpwblZxlH7H4igUYArwuVzfal1nh1ELhpgMYXMXWGgGy1RID9oTe6Y1n
gkWO2gP1D1iFoeTkiARI4tTUNwJgQj5Zq+JyC5Dv7BdLX4s3rTVDH5Tfjs6I4hSw
M+CkFSSpKWgoK+qBpU9rSXtIeqLZcJ9M3M6xOS4nZzXUI37dW7iJ4J7KbP4H4N8r
4VvCbFi0Uenwne9xXFSgIWKOAyBEroNxv5w+/qVr9E9IvnUiMVjCTcSWHtO8Bibl
FFnCDEm7ow2VXFhCIH0cLWlyrNCZcaHfkKnwB7cb2jULWICeSImH/na9BnDyBadK
TyOU5vFxrkWGbm1HAs5TyjrFR4BU+OfWJrFKy/HM8xkv3prJcWGUVpzgeId8go6I
zq7nqxlY5/4mUAdarAG/qH5dylJuEs8z1eXiR0sTGX4swEWRaI9FwIKztWrurVPt
CfvSX8PGtbSVVXJaJtpm3o4bcnkFj6B/5Km5BlXqDab+IoABQgOzBjJ9iD0Qsi2L
EuqbNan7722/G+4jVtwG8Afkb14anhpwpVQY1PmDxOolEL/LmgdsIqcyuR9pNUDJ
Sa4tkoRxqM0keLtDrTFM2dc6oc739NJ+PCoiA61hWuhfK1e5EW9efY7/VOfDBfkI
4asdjXE5lx296C1JhvlAFkqv7XgnnnEbXLWCYYuuPiJ1QI1BkeLClFW8U/3op3C8
Zm3xXkgPwYrWyH3E1fk4pS0GbGKH+UyhwVXxLyDPSJX4BTWrVi8swjDZlI+NISDI
K7DBCK1Mhrk1Kb+Zanrylf0q0H6sEhBrMSk0XiYA69IZnX0K8S2WQBbSVxXfb+As
y+/0VDcz9gyZWOS7ujTvjoQdh4Gd+WXFnymetqde14kIMgM8+XXrBska1ULOD/Pd
MTUgp8v+cEVCDm/CPJnqngkmu1G7Q7iYNK6VsmuJo83ukvAd4RcA6Q2OI2ICMNGW
Rys53LNg2oAVP25k0JAcp7SMvLBGyktT+O6tlWb3YLcCmpdd0+jqJ3wkE5hag/Qd
sXuBF9m1V2qEbpeHq7ybSxUm9TZgZEsHhJicKWgS0++7QnWMeP18FXwzj+xHs2Uw
X5cA/cTZGiO7y7LyBqg9Ce41HNIP3whzEZJi6o44Nq3Eiz4SsQRZiZUfSrSLHQyi
OfesXU6qnMfOzr1k/EnJPoO9w1UV03yN9FfB3yO7+c8zjtmtcRP9/YRoTUIHtt8k
P9YXuARDcnoOccGkFf7HkktGg7kq0iFipqSyBK232Dlh1J/jBrPDdZZDsqcluwZn
ykSGmpCgRW59hwy/joHOSJweRinTk6jWZbUs84/LA3FmcG6sHXZSzBhP7g5evWwy
SpdqDCO1by7QseMq8FTFwAle7IPjXMd05LoqICkRsuCtEe2BHWh3e0qki+avS+O4
fijONpxAP4CYWBre2gfG2MJn6NUKhgU7l9FxX427T5W0cJk/f+BO8hdMchOzCx/T
UBiKCg/Tl0HSn4ujWWvDYSM/alCljXEjg91E5x/fXwqZR8tKjzgC4+e1Ndc4ahqB
+XsPP+E5hVlffiJB6PhkiKCSTFoob2BBr7EHMYSkQ/c2K5iClmIwVgLJiVz/0ofV
NN2yaX3oEidud9gCAAY56V51WK3biP1QarJsttNBCvpjd8FQU/4YSVnqmFvvrumm
ZG7IB5uJbX7CG940u7PWEMz6DiwHVTAGa1obyA6YBOMgR6A3UQB1soJB3lMpupLf
D4ToPjUvnSSxnuEvkDy0Ld6ka8G1X+ljJrvhz5/1Y/VTIIH6Otz/tPv09RI8KrR4
0GPH0g6ZFqArRjtHf6VSBEhBD3nYiv6p7LmMcMpyMd78/2zqwleJBhP8TuVkN4Qw
60Jp6x4BDanpUVPLxvlaGU1FnlmoZ63OmTpQiDzIREROyGU4RB2izqdpSnizd3wo
NMxsyHUaomotOmOIO5QuhA/a4miaGy1iJD9a/jSCqHUwPLzhuiuL5OL/UUse6IXk
XCBsHlYkaK5Uhh0Kx/2e/0M4nM18PWr1AC4eXefHkJP1Y9pzsr7/kjhUX3lXeoGL
AVLnJ3gl/VFEk67bcXZq1ny9L2/byBH4Z7sLfGRlPY1jUY3jr1V59hmE38obT8LI
6F6zWELMRDegsagud0pImyut9khbpcWX0La7uIgwGxhLNN4baNcRpsiPh/UZakzf
fwFklFwSfQqisjRCza+Pv2tyBDpEUOqVNKbLIthWXJivdA6KvVbuEJGoUoZJ9yni
Yqpj59RWCIQ16Y5UFK9zYG6+nyZ86VIoqmdRGYXWYB7BYOwtQ9O369DtefKvV4Nk
LUfQQ8cTn46aKp80uhdyEiupk45nZyvlrbUvHfiYlvA7y9oeiR/sKvy6oME8xNQP
0mtXRA4F4V06vmnBbAhil0pY1iEcl8/DeiRWrS9wwoA/r+HgM4n8ysM0n+xr3gWF
dw0NU70JoceR4ZWEvRwfNxsVypO4z/cVXx+P3BjwRv117AY2jb4f6OUfc8ckvybB
7iM5bfn2WaG4o/jJcB1wWgQaUvAN80fmCPN+nncXVQ19BA5oDM0sE/2kNtw15tfg
WF+WE4nwYIgnx7DF7+5wanmEzEADvwTOsNPy+up6BwwgIr639y/EGUK8zXBUh+/r
siZR/zgz/fFr20rgdbu9johFobjVcPR764gBMtDt6WFSyGfOi2unRcElxcupWUaH
uMQ9EHbZyl4lQNtVgmPqgOb4jgaaQp1PNaizL9+mLtwh6SgOs/+eQFawmlke7lRo
gEDnwuupg7wgm00wSr/dvwiCzoBjCRk/ziESHWJFnfYvMBEAzSYc8XhOyVKHLI1K
0T++eX8ylhntV4vXcIedPosB3+cGp8XbjikZDb7m7dcwXNlRIB9hcoUSD0IKnhH+
Si/8w69grv+qza+RDNsgRFm0CDCowpXesybNnNNq/+MB6554t2KeMzf5Spj/ex8I
dlwGwua4+5EnItA3zlcdY7UHnl0bdnBPqlUyGHEKZMJSdci4H9NDm/coExbVwdZm
NXi4NBDEpItBGJGMdqHC7palLRVVw0vG1NJUS4yZF7vLBA8t1vkdzhC5X4n0DlXW
TAv3VtfvybWGVz6FOYjV/b5/U3Kvr6qyrCiXI3S9gdmD7iWoTflM4zVuMVEV51q3
Majkn1RgJymp8DuOS2Bi4a13VQKeehgqLB8+q05G40ZspG/YB6FP2jM1Zi418Gnt
fJWaBgD9RRMjmDdazcKzqWQLQvWAl2959vNkWyoactFf0gQBGeV3DKT/QVqQZ7rT
ZUbmuEGXYlzP+DWK60uFpto7QaoKNy2UzGDZBupYp8/Vb68ZuHA/Z92eV9UzU2Zt
JBGoUSjaNRbAY4NmsxkcaYm7kD/gNSyX1ZSZVZrQCwSAZbcLIxEqYO1I/HTqDXG8
k2BhLJQ1jcK012/Fh+VbDScvf7zgZR+QUGhUyYYb0YcPPcFIxw3dg+fL3n5CmRK6
90bVb4PBFAPNp56bF7c3+Pts/HDXJdYrHXHz1qAyYuV0H1CyYkPD4lCNyaRzQ7NJ
DHyh9OdX9uZkljuR2D77PKo+DmLU63fWuwYGjfoeFn/AufOShI0wE2hOu/TlwIHV
xn+Fd2CyNefcyUdGFeTZlEyibJd9f3cAwpMMOGKbWSWKOnhRCsbqP0aYvkVolsX5
5avQHtuMm7C6CsKZJOkRr9I8/y/OiQMOA96fL5Yf/UZ9acA6MP4WVXixa//a2kY1
vrqYBv7DBiSJ15T4QimfWYHjX5twI0Kbu/DLkh5npN4=
`protect END_PROTECTED
