`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9T6UhPpqmy7SXw1uOEvXkPsM/Nc+2dOHrM5QCbO4tKX3h8uQCYdXCpQ/x1ZWRVkT
CSoZhtrapD5ytHgqdmjRp2tYlcJaNbrEc4XFqB6aBYEcwLljBaW7JtIwCuFdLr+H
zBMLH7PTpB0WBVVEJ8i2Myljz1z+8WHo9xczcGvdq4lDXvoh35bBEBZqcYBJqF+Q
szsCf+EV+aJzfpP7qo/1ty1RFeUlWjfLm8Xq3Az5rE7laklJ4g6PcjBQbaJ2sw2P
eVnldh14jxKspgccNyATA2tUXKnw+Gd0lcuP8B1QKvxdLtrPVp1AMVuFe3Qus6o/
ww3ATTVl/54Yf9U0gFv2v1/du+mz5MiVheAYJQxY/m85FzCbstcpiAYgDJd/piAb
eoy/BulH++GQ8bFp10W0KgkN0kA/ZFI0kSVQF2fH5sA6/KJHEOB0jqbSwXX3Otmf
ZlB+ONafrPZcl/xVVmDBGU68znJOqzFYSdiz+2rnb1sEFBd15bDwEJzwwAXkwFfg
/bSHaPAx0kP9K0H9uhTlww==
`protect END_PROTECTED
