`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QayOJDE8rhwUv6kLz0m0NnOhB/LBE0wKWeCa8AVZJgoHvaeqDrpPU4kZLQTwTZPQ
wkQ1HFbubWg2baNbCnaMgMNB0zQE7nLjKSPv0Sqi9B3XjDTusIGyoZymHqBUGG4x
XgolCY90U82f1Hgf+V7sEQOk9vno6kXxkF9kwY9+y8h+C/9A7glojwyJL07xA7Lz
I6lwZC0Er3x50cQqOO13VICoZWgqzxi6J4RoCBYmEgOJn0xwAWa4Gi3lxgjSc+jg
Ik+HyDlzx8+yBiVo/qOXsg01fqoii+js8RWHmxtx+heFqpPTUWkZYKsiF+e96yPi
tOKdcMhM+0+tTBGtf+xoBxQZv/FNh8FM4Mck0B1F/lhy+sFqX4VdYfTcldoCumQc
wvu/z1z+PdYjRQRe+rwyoG1wcpLxsamTAJWMb6+Yc3SWRVoiUgwPjUTXrz4hlNaU
fPLIREKoXn9NGUn6ANtUKC/6lMj9fKk8yf+9aXBai6O0gq9EToFOrOlF7AniB97d
g/uMPBqowSKd1G7lbsTc4FGXZ5RU1+VjPu6La/O+eZcxu43toGWAze9ADcnXX4O3
BQE0nolp3ePkQ5QTyWIpdHtCvu52q8bgesNMfsuVWrpEqPb2dq0Dv8aIClVLiWz7
lAWdNM+ctV49oN4rEzs1aSKgu7/VHrSrBsQq7ueMOBCyfLU0v6eCeauwKsSb9x0w
N4v7WSesRHv23D48WHSKTYSWPiS13JGcfyHpfB/aLfmEua+u/sFHyEXlBMKF2oTt
AQIPzoB91pMS8iGwPL0bhwwUrOgJ3JppOPAMORfIdnsx3R0IXcOE74/ZRiEU7eqJ
mQ2adOJD57C8TUrDXbEKrCdTBUKHnJSA3TSqTddd5GpiQhFMmIk73kd905ww0KO6
3qWZZZyZiWeFijXI8D2ciZ7ca7J4b3qcrR3ODmlJybs18Fgu0KhffFRY8qZzNNG1
UE6xKdEhqkQNzoS0IYAanCxI0rQj3c7fnkjan0mGC44OoNkgtdsn7VVYNe81Nj9+
rwsTT/62hCSeWs4n5ymp79psL9kd9+8oa2qIk9gmYwzTrTJjRRODuIFT5asal6EI
t9yKfAH78PWQ89JncVPyu/fSAe4wQcBCDhNdpNc5B+somQSw6UMUykcLG0qvCHUR
fgNrweNM5z87/gP6EVOwu5/6KwEKwORjp0oOhAE9y6Rztuz1xJIYlqI/nbVzl0CV
upz8bpRZ0aZAj/khdikCevAfTHs94M0G0B504AsHsJZtVnlUPYvlfKHdTtbwNfYt
fd/04dCpWwlFnaI3jbP5Eh2UBmZGIOgg6QuySAyPs4ATUfMh0KvCblKEfV0ABP8Z
RBrHJBWVSHBNkd/igI2cJm5pxNJKAwT7lH5figdxcmd3sapSK7SqBshcMwszjAbL
8NNcOJwG/7kjYneLaNbZKCpIKIJP/O+TNXixHekHinnaaNK/r0NKHds2of6aD3LG
V05jcWoRPm5FoMhYxK6ypYSSbA2AXyg7o/o0/nxku25v5LUl5e2NJHqA74VtNuLW
TzzE481hcMrhLFLTNt9ZhY5KLQy53I9SKFUcVkZnK9vx0dAs7PeA8rvrG5EL3400
POfV/bAZ+rRukr7Xxn+dQZCmJSll7h1NBO0RCEWA+7sJEhNyCDMCp0PhDyUyiXu7
QTeVrWSX9HV9Q/qi3GnnXq7F+/1dGgb4BJJ6Xlc3JpArAv1hoGrNs+HM/HWq2cdJ
z/eB5Pk1V3xt4sMkoxx4Ig1Jk8EpgKyn8wID4imwjP7/V4bpBuK8BE2OWUWbTJC3
fiq/Wpc8d2ba/d2B9LcyNDIaBYfhkn5GtnV4xc5uHoEjXi3tKnu7GrBuVkM+GT71
9rZWnHfiwgPqVlgCgie7wHcP7AdtR9nadulfGdLt1vpS5uaHUCotXUgmIcx+XI3i
8Y+mvqvzhSn71z7K5/tcceD0ihTKEUYQvCZ1WOZVFIdF9sZUvwLrPPQOO4qlycw3
Q1YgUSeD0cBGnO+gvOcnfgbsUrWrlR5gwIyd2wUnwU+KAet91pYyXUW0uVzMM9mt
dQ9xsXSjmYk0jd3PcWVjP6ewJxeW7b2YDy383x7ir32CVlpeht58VLD2m3kdF/3W
zZzzAaVHAu0nkwY1QN1xV4+C99gGbxGwOz+hHuL+DgMOPZEkBxFW7JyQ8fPJmlDC
2KBYCUyTxeUaE5Xz+LNvtQ1piVFKDJf5WXm04GnnNs71riFb+Usci19yTmacWhya
ZGoZtaT74pG8cQtkepXBEe0rFaz1qq9ZYOC4IqhA02Ro5hgI+WffHiHEnpc5pXFm
1OOmrhNGR169VTutfS344HEZvafoUmTWDV5Hs+ZN3BOly8yaveXtDSBSOJvCHaMo
JYS9Tu4sdyYcRno+JBFTezVNR9QA3uFyW0c/bCjoxz7zo/x/Vk53o3EUfM3iv87Y
UNUzRomZWbmiUyFQjEjAsjqAv+etJUL3CX48EKl/VdCmCaNh+98oJ52oa+g2rKeZ
0cXqhQqwt16p87DjBSMiUjIXsFQVxVKvcAUCav8UGQjNMtupFwVp9jlheqeIURQG
vAyYDlBaPE5+Nl625GLjUxvMI7J28MZtU6W55PstfKi2FpeXnVrxgXkKFh+35P64
1sdhm4J+rN8aXK9Cxlk290OL8AzEjBPUpIteNXR/cA2Zi1Wwwco46jzN8ZXF3sY4
h4Zf9tMOddfol9GRArFatrdvboc0LbX+K+LfVcVRnTPixuD5qaJOpfn8Q4Sn7f3m
werlrl54UtZ+9ybLfZOihSoCIJ+P6LVFHiLBgfIgmDmXLb43l/3kkXdgPtCpIE5V
aQJ3H0yjGo0xkG43md272VuEw9BMiaH62Tltc+dyB4Nuuw+PijUXD7Eycqx1YBU5
77l8uphZZlEHnhRaKXftkTaOmtYcGok/RnW2A4G5oQNjPaGvKyYliz4uQ5QZrdeP
tzGQmsFPBqpnGkHpLj6ZLz30uqn6bS+ftIRoRA8IFkuSxpj1GowqbQaU+GUThkyB
rNNui8VVuZymYifkuUqSp9A5lidlyBwZM9OoJzzUdg0KGsATEPKr2pckevY0BZSB
JurFTJTa/D6c/926AtRNz5SfGeQJd9digVMkkfTgAq2P0oxU38LAMn+ZkLAu1LGh
i7bc43Jokcs8TeEWJEyixj90HOOhzEA9gsJn1MqwPYDZ705sl0VH5GnyGOkrY9zg
AU349NdQPP3P9+5HHtRgtF1j/SHH34hp0ZpoUawfab9s0mCoawuhG3ZhbWNmbJo5
lZyx+hrWp3FJanQk4bTAfVk8iInOQ8CoHRS/mQpXywq6jvg2dlmQJjRhFv/4ZW70
AqIU2jLOJDWtEbZ5wVxxkeE6XED6HVwi/rxWi9lTjqWiKR6kYZkOxhsyKSpYOqVX
MJu7gpbqjUDkyB6i7eCzw5nWEDKVRFvMJQqGZbsgokjbdvf86jy6VfWYG5TQP7gk
v7ZS2ioOMvW3B7eQ4ny5ex2z/wZle9Io9e8aS6zWKRejdL5k4tFRkh7TuKgIxHdZ
ovTBmW+5ZMAxq8in0O1nJEu+dVD+X/u1oaXBSXRJx5k1yJWaZ99p+sfU2Okk3YWW
fEhPegO6COnKeL+W1gt7HjM97x99RdwS8uCEwTv21s61/SGHJE58Egfmcrk6xdi5
LCxWlcNNohUSbUyBRX+6Y+ZAAPqfKwvCJOTvMpeRRMfIejaPlMmsLbca8aTOVtTd
/zLC4lYaXFNPykh4RQt4MakT5TvKyuBb3ZgHov3wPpum9S2A8Qwa7MrLO0GkuEih
RMAi4F55ginDhYbGG+yoxeOJ4fyP0MCwfII5JGc/beORAAATeSkBkjytoEbn+C0P
oyA36osWiuo6xZj3uzbBUFTolk/K+GMQ2b6GMlpNUt06c/dBSNg3dz+Alim0NUhQ
kL5xLZjRF5f68eMi/eTMB38sE4wGo1r9p/nFLgFSGV15JdZ7b378miwQfuXFTCi/
t+bi8yX9zJuyuWr9bcmi4RdeJYNWmsmJDin5AfdT7w9m6LubeYqDd2yWfOqysvLU
DfCQKuPBXCUsStX1KJ/ZdNr/GmeZrHoqAOSBZ1vNZRmRGBs066Rr8coPI+D07Jdb
dMVGEX+8JysAvHhepMbzhC86yQvmZO1vbsTf0SICtJnvAsuORFQ/tR9qfND653IE
nYeH2BVybZOXujyMnzZRBd442HxIf9pmmjEOfC+hCz+y6mVosP6kFWhdBX7KKTFV
CfTs6jcJAwLYhlVBz9ia+3D67Rzb4GdUU0PSKfMYNUfmQ83pwKncnEqEtKyusOIZ
biWrDmB1iECMbgJKvkC67nBNpJYobKbuaec7QtiaFD1Z5EuevFjhGb/78tuHVtUH
3wjuO92hi5tkOhClBuS1rRYv567FROFEkIAefc5PG7s50lrUi39OmVNOvO8ImXkd
DAdJeZZeGu8tKn9JhzP3WfXLrJfbATkiOUIlIPdLQBXATGow0uyWOi9To7iJcl3s
a0ISjmocfakjgTt/is7OKVKNtsbXXtwi3O9E0+ouwG1/uxPeXbMcA4STgYt/yvrl
DwaUTxIgi7TUyA95QuysG0DJE7nIXf6TMIiPWORSK2zXKZjyKjKFdiyi/OWgK+ay
eZOoRSckin2HeUe+wnnZEBLFCgrXtU6IVR8lwBZ5FgLGsYXquYHW9dNt+9pQKPYQ
4MFUSZSzxyBKkWQ1dwYs9CH6iPQwS9Tcd0Nk3foEY+dSJzMTWPQLplL9z7b9LO1l
8GHdn6+V+SUq+0cO2AErJoebhS5Xan4ZdL3sEusllKuZdVQi7kuo9/Hy1d9SUK2O
uH6ZoklB+ACKHSksO4jcI/vQBm24wVpSyeBmcDTYCwIiF9QyRdlCHt7VYvqbUEjf
wVpwzPHUpdZ9JSM8hpLFFYeaEES2EQcRp5pzTV+Tvu0=
`protect END_PROTECTED
