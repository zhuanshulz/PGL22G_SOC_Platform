`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nUgY6ATPbLPC/AQr/LADERRsaBuwGOxXFenicxIgEqvSUFvEfJjC/ts283FjjB+O
JJ9UIc2rS1y/UDdnSpK+wxPjgfNmGLbjYtGrsaJm9438E/2ZEq6GL7hfQqDM/seV
slvnLLY64YbPyg8kpcaKH8YmcsFBuN/QH2V15CaMHuea9OuJ4wyHMbaiWGPaPxuY
HtT6CHXKbKLEpHfIek0Goj7L3OrWS69c+Jtid/Ug0HC+Zd9P+/GT+J45cGc5VYFy
CRSCb3q/x52aTaT4/G5h7loeSDVD+70POyOkGvQvjsYrEEnQWLfa4eLDa6IbfZX5
yCJ7wqgj4TgKCkdtjQTgBr5OVOM4P2WK8FjSW1QeBHdMgUnat7hWCWiyH0Dg8AvW
kbc2mGJfrlsouHkuBZNzxg6BdUkI60PNrI6U463XgMMfIGohy0kxrICdl6sJyOPX
zlK6eEKcJrn9E0XKNOzv9ZZBsK5It4880gJFuZyPVrc1Y9mrvmOXQCznXfHqDq1V
lbp9R03KeeW9UCnjT5wI59kFfnBhG6En0AvseTXUqorMb4luH4iA4PcIx+VgLZsT
E4MPi2/U31leHUyMjrWp0fgKYzQb8+7m4Iw5rP6tZT6AO6KwRYNLFXtd0UGE2AVz
t7OsloiXrpBMzC7faLdHq8agSpeh92AtmIWY5lFJAC+9b1KyE5O7m0+UG5ilPgx3
dLmksFaJ9y8wwrtTSevbzS8KK+dcyoIooumeaeCN7Jq7OLyMsB+zQimm6zlyDUdu
v3yn/JWhdB4S/S9//nuD+uDUTUOrM4hgyCjU/r+D0Yemc3PpLZRhO5M3m+igJQj7
IRxzr9nreQT19aKTwOf/V5gochWQWawDYxCcdBKHrzVSGQR7JkY1RcVIoNSArNEM
0zouM6B8Ub6za8GYsE1f2npZCnt0CVr0yrwBbl32fjXhwhfbkCBLvEBUVr9e6eAh
cKPZ5oSBKlb/QCayRYt+szw7VvcGyJvlLEtlzDinhRB1UG+WNALgcNvCNPISOOEJ
wtqcye2ptv/XihBS6wyX6aCx5SRl666ziHuD9owWI2xog40vaBfl85jZ1SPskpmF
u7j2+Hso09NlKT5XfDkeyBYJa4Z8i0tD59uzrZJfk7aQrgFDdiI1RZAgT8wWY8uB
rKqjCeHHiV+h0q/fybCfk92HCtAmDJucCKje5CeahJNMPU+pmvnx3kY10hl+RIOd
oigiQ9R1PNcrJtNZsSGXuECzGo1iskJrYD2atNMHJLFLTJMfdKEPmolgYxrOM3br
wAmYqf4P+ZdjEv7vHVUJgityefwEK5XkLJuwg/L/4bGZJ1Pw1317yJ8KZpowqRw3
JlEsy/zeN+KmixrKpBRY12jAGAAlPh8UKi7OLpk8Xy+Cj1DnQ/pW1G7YtvMiwdrD
/V4L+YcVJsY8Pz2wr3nUc6/kWNt0ZpOPjxvK11qAw9u8/sPlw1j/nIXB4dwegYMR
Zux81ilT8TAphzJhzQpC0QWZOI2UR+xzM2S5B61WGrewCXeMkUr9TIRKAMSBDn8L
y03955OA1O9r1+0sfEJEFQ9zNA0FT92yr+cF0dysorIPvIGXMFTIxLXGXhBhfg3W
2XWYN3gEfwZJsIla3EXWwH7ZY0bv0gNYMGIAq8Y699ZYcLZYQu0Jk/w/EdMdxPOA
MQZwEk6zYn2Q3Ab60Q99lTjmIHDgQzC5EwxM+RQucd7uhabPa6AUwGkjWFfB/DmS
iPVkfgQm0qUjsUx51jBCCPSfnyqjJyVcf0G6rZN1AtZxoNrsZ83Q5N1YEd30UnvP
vDJOiCGvWpMEBcwv2LiXBdPPXBVkopQRP1VsSbIGELfClg/EMfu394qkb9+R7fH/
3xGbeT/kTVdlksKZgoYnvjM5gaDvlKRXDfSNoJYf/dAE2bpDLQgZfuLL9YqCnmLN
7VgcVeqnd9yPLyXkAQr00gtrgMu3Epqo1p1qe5rs4oRYTOlWIy7amiFhdQgUtveV
uSAMX3a1c/AOta979YB2EMyycFvI8mYI+kwkRw8MYJ1ukfjBuHmLvuNzJrmZ8QMv
aaUy2lE55wytgcSCgcagLDl+lEixCh4311r5eUlMI1xb5XQW/mLyK1SHQtFhd34X
kn7XZ0xCrV720cRfE3LIcvJ27Lw1eCXX+1rwTJgj2RPWOFEUSmXy8hfcP6EMeyTB
sMkG92X+jAVkeiTSt6tGFKLOQWmvYN7vVY7dGvIjOmtsEPNqru1mwruqDq3MKGTW
c7ZrzM9TCpcMqsmmCV2D8GHeSIGTZxUPAl8cOW5jIezNAq1Lt18aO2epPJ8RVMcA
eJmuogXeayTRoGHAE5n36UXeAKAr6A39Aky29emGXw1YVr0jNN8E/eQmuOMOajK5
pRJFKwtC22NO3x1xFcAMjB1bpxZUziGN8XayrG+AeGdr9zbhqW3scwEZ+aJc5hON
AUGMcVVcvRB9yc38S+XkjcVjoAPEjQ4NeclecqjC7+E9DZiR8KBU9iwvOMrYSqyi
ts+pyC1eu6ttAm6UMON+mEVUZJEDB5NRZmhbPHsfS7A7pr7CAnWu8AKRQEaNNzr9
DtpA2hNSfkOG20j7hy0LnLMTW2VV03ik6kGY9bbnWPQgPUZfIq17f4WNWMwZn0L8
vt0VNb8WrXFpUcxvMS7jUhvyDhD86vYAGLUuxYgdXq0Op7cOxOVVyaM70vzZhk+8
Ml8Ww8ZjdyfmK0JHbnsLM0QodO+uOjS0ec9NSQYGhi6nR+KLzHZuaxJSUkGxtsQp
uacvQ4R5f+3fsNZ7YOrpOn+wFb7FuzRmaEE8PkC6sE8apLNz99wcZAAiwtAo0zir
LCuwfTrpBxIkoFeQB3Tjmr0ZJFKzclwAw3xfBwU18aSlSFiFaslajbhduO6A8Los
DsNjplIVVrKNxepvZaeciQP6A2fHGkSqm2W7Ztt6spIRqRRxGqWQQnsI9jU1uIby
BXwjDFPPPVuWTCmf/4oGp7F1EPCRI7Z0XlELW6HHME5nkt7lRKiqgWXRsS4g3ISs
MnSYz4cjUWqpbF1RYthCGBdhrL5H3YLREdwLSAdW53H/Xyh79lb+9Jttben+MbS/
XqTnkRrpQ6E+25QoiDwh2oedspldg39t1z/VvZ61iVJMjACBvYp6qcZlgEiC/ViS
qHyUPs/FkgjD3q6GnbGjMBzokU8vOK3LwM11+zfzquv4j9LUdYJv2VtKD+OG1ir4
OYuDiHnelTyCdb/rPc5+llEsUqFfWGe9pfnEAUCspGNFOhoTPCkXjU8kKmOeLT4T
DAKsGHcGaDkDU8FPOyytivwgxeCnthYEO9EuV+rbBqb1+XhaHwf8YQZ8rDujOqMX
bQAW0CUtGKGAbGPfUYh2XeWaGGVUns+/l06Pmb6OsZvd9VVsF+kS3fTtRMmkuO+B
puayt+T8ZN7Mwy2TcO+2d1KIX73Cjc4YGvstiKjcQlYJMIalkUtoRHd9/u0F6jq7
wBP3hIxnj2HzV5IZ6vZjmcgoGeTqnOmnPzA0rhCcs+ZL961Q4H+99kpffu+Yi5LS
gCkQ1s/8mG3DlZqCiFB1ObNGB095WDV7jA3ELutGvNH45XVcz5gzMGRELm8nQbrz
xH6Ogc5EIF7dPHlMC3qIG1M7GuyKUiR/hzKO/DCWShVWBwq40kYPv4GH6tkOYYhI
AGVVZbnifoNHRmjsf3LKKjH7GOK5a0+Zbwb0h/9siYR5hnEClNk9fGlPTLnJU5yq
iFnjxfddpnoAF+6QP3yIM4+OpYS4EkXJnHTfNU5Ojti/PkQmRzybqF2c4GQakkp/
N0iGyM2OElziir96gi/z75l4HCa9UghMLgxxb15KtOGHmu6ZnBu2Q5kbf890Ahb1
pC7jdItzw7y2x7K+tcTkuBmEltjQ1Sob8G4b9LTARo/rKEyukbWvsbrC0AoPwu/+
P7FlpWxqvHYF6BbzSJWQjDGGla5XgN1hPG1Xc82AcCAitr7SnFmHMctG2/dw9RkF
TyCsNE9rtQxBzg2USp8ctT1qPbr9yYPXIc9g9hmZ+s/yF4CoRFnIPBqaEMqt6Wpc
H6ZydWB7/jAjRaRe5df06Q==
`protect END_PROTECTED
