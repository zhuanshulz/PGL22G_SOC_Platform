`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3ry/MvX56izTyC4gmcfSaRty1I8RmDN11+pzP9xm9vr2gJJR9QW3zkPzUbUojXqv
4tNCImpW/c+iUhmvt+geGhtF4YqqNgqxCvGQ0oFhaUeHdoC/n5wQxmlIoaTR8BwL
IAnpyP8E2MxCjA4hV+5oxqPdY7XzFRmg0ZHtGEj5aYNLmgYMids0++MVbTyYoRi/
csEEUdZAwsgbpLQQNWwzM89VfeTuqIAikfDSVqTnNURBg7yHooSdsyJ2BDyOjYl0
Qk2ljTWC66FM6Ws0q06CsTQYXAqJT80hgbvW7zzGYLJhUL9gqhTysza/277f7tLh
U/7aaoQRP/5loSuwKNyU08Yejs0KtHnxkpqINGijIsOug9kNhsW5lTqGIYIeYJiq
c2mdZOPhogFWJ3AzWQWV8ciyFQNo38yeVfJdL7I+9nXyaYNZH4Tpnl15ZjTx528d
0mY5t1vbyobz8CE+bwILxQYBoXG/lmxUbs6yXZFh2ek=
`protect END_PROTECTED
