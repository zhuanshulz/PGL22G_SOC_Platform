`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S5xEI/aV+XthF9uUAV9cdNOvnVB4nJGjVllVctvkldu7OqCel4E6BtwInECcZVYi
KoVdHnZ/OnliyLrGrkRJq+ZwTw5nnar3GNq8SJKtMI1m3ZBEWjvoIi4QymJVgVTj
ML5GFMqFT6iIBa+jeEfTKMZ54q7R+8JFrrVAmIRogDVy8K8sSHxVsCldzmbzCZ2a
WhEOzML7n+fmJkFAq5ib8OeqQQ7lc9Kzila/UtbCh4pjkS33y+wmfFbZhh/GCvnb
7pY48kkNzznailBRZYCYo6Iq8Gb3VGxeA/ekD3LEUoWFdBrk4UAHEYpCVetgxect
dsUmGTXFQWedskBpxkrhapNEgF9pkz0OrBPkLX8AjwKCpAFtWnKfDLt+4VHVzHcc
2DXXFU1SJfYRW161eOH4OvUSpKS8bvNRMxEVGLdrLHIWwMywJD1GBDtx742+Q0Rt
tdITtMC+aCTDMXZ7wahP+eGTtflig67AZVhQIrTb/zI92EB5fFOh5RF5oqjs2v85
5cox3TKjo3c+vfE34zQDLJYVFMEM2ziN8fH2EqF5N3K5PjhI1BjxRLXn+aJ73ooC
92pWIhJz6gI/hK21iwIO4Urv2F77YzCTSiMQubKxX1j+zfOuyCuBQlmpu4IKfKE9
/54MiREthAKbY1VAHxsfdge6ofA5Ov7W7d1I1UuNqxgxi1Ue+DQ46J26rpWIExwI
lCtI10lsPGFElnmVAY5KvsOXxLy8UtUEXB+gBbAvDvlXQKmy/aRCBl9PPs94xPa7
Mp9WC15ZqDkv7OxrYquUoTVYMbG4xB6iOyeotSwCvpJU2g7NEIsQSDk7yb0JMNLk
bphhyO2rHl4PNgGVX7jaYIOg1nkxZ/ptu4Yz8ZaVVacZgOBntcKXJSVNcZR+q9sE
GkY1r+kn2bWOw8l77cMPqcHYoeVL9Il+YyytWNCJY5tyGy4EVv195XuO58xg5GN/
iRG0+s/QsYT5btGqNfgP4S2iTJxX/cP5EcjeriU21NZxj7cfBc7gUEllUWWTR4jG
rCh1yltnb/+lx2oT5TfuWyE8yJOYdJnNt2Mt4uCGX/F69vRInwXcEF/7vC0mZB3O
MYc63F5+W1c6Qq/DkLA4+ZzrO/pbEOsn2/2g70Qbd6/juEDgGf222zHUMzdpo3Lr
4d1aUNLe31VJG9D7xVP9s29puEmHILeOR4nrY9vXAoIaSdITcUMjGOpEIlsbMLsf
MMKttPdnZ5ya/P8alAFo1d0VHahoTAaqybvdQs3Q7tSRkb/Edi9VrBsxlSUqmtvV
CLAsDpsMcu3Z+yoKnqjSFwkl3PthdoTVqy+OpRZLTV74UVcM6zgai2sd3wZavUwJ
mVkdxdydquqoNY62pPBHnJLnKso0/RbZyb9a/j5i0h+6POUunGZduS2P7kCSrHaC
NhPGQ2IEYD0pcu5DtvTKHdCKVgeeCpOtiV15SNlx7mE3HrH8HYm1+yJ6IaH3etPp
mXYY9kOXmHPC2qlabB/kDk1YIZ5/9uz6QgS/aUUgKAg=
`protect END_PROTECTED
