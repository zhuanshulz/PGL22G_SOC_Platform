`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0W7bdNhCKeFipSrw135gxluwxfAgL2NQrMXpf96+W222cnS5dMB+tToX/Gja4o0F
o9Z9xD0zRC53Yr3rPdY31IS4acS6wgFb89P6OsMB0QeXp5KwpG2XkmoBcgXR7cTr
JvK47BqufXAiUkpnCdw7kXxn2Q/g5elQWE14dg2Zd3V/B9jdTP5SNlZBnvnhNn3V
CBlw3uba2BaWHlJNfiR75zWH4JcrIOymFmz50rXQ6Pfn7JAbTNTyPQC89Qun4tey
Iy32lhzp+RxkYChN2K91vaH6F52+GtcKfEvsy1ndbNa6+ttsm4qTiCLyGNRhfSMC
/NulNZXUD8wtJJwcTzPWoICPQfRhFJn8glPSsgkkem94FQ+caixq2nRJrmBB4iHL
hWI4s8USr7z/9n/gEcVoRQBgzVZhi5VXTAWIwXL1Yhnd6+ijjymgcg0Yv/XOExWj
bg+MkChSoK6pYqOG6YM7qsOP2OOMcdSqQcMqX8SljSQ1yXcUoQalQMd8JnIhqSfL
yZcaNIqhInflxj76nCOQM8OVBdFuv16aAN1TeJN/D0H0I7zCoSM6A2wnnp8MtkZB
LQ+3MOT7vqffiQtr1qGKbg==
`protect END_PROTECTED
