`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZLStunOaFcgzRqG43osrqiptdBXZ4ekytAXSXNSorvo0wgYCw9S2WMkls/rpzRDv
nbYeEZomP2PN2Vq4CKHoSQfkfFev3vEEDZZSQcozXNj9s78zU2qWBgCQ5xB+xxnl
H9mkSy6Dj03ODx6U/u/Yt2bK+NOKBUFmjXxfFVrHQwQJyzIi+7J28hOt8JSXF8mi
QQUqmRYm6TE+aXGxRYgqUi/XV5gUM+5WSO83gZX5JYdqDoNzDv86DvNmn8sQZtVM
4lr9OqLGYnUCy9joNSZmk5OZZ/zy7JaNYyg5adZceIBDIFpplInmg61mcC9vo7ZC
FmEWeWc9uJNqOVsQAIhbq1eEz4VEcUzlJ3w2hvYwZJHR0L1SbKwS6W3J8cO/fV8H
gvDIg4Q41/Pp5VLEg1TedSIk/SdXpXHR4xy4i65lwTTyy7sAtAYsj6nvsgg38dEJ
lrAjYcYV5ZevVBpP0awkd5Zw4ba2gc1iOzaOfHJRltLIxxELBXpvul+r298ao3Sv
Rz+eOziLfLmkXKzSilH2+Tk3A0SZ31o92Ujao1NoOce2xjjaU3Wz67hc6e/bcTbS
g3bc2dzkE4QkIQOBcw7hI7sBE25Z9NHaVJWRvchfPUQv6ChJi6YsEvKrHUyBftQQ
o4zi0Cvm1N9liQ3So8dug66mQ5da/ym9cZkZ59hrqpjy+oIYY3Xb4RkbBaDSGOFd
mYUEjyYiHFScFlrmhazi2ASuqEVix+YT+ROudDfFuLmGU1L8b1yevRzIFlUs8CTN
/rOlnfP1eOQTEjuS/KfB2Q==
`protect END_PROTECTED
