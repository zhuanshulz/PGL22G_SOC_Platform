`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cYZbRDp2M1uZVzFt3qw6UuM1hKdsIUsaVyXcMytgMNq1LHOcGGng9uwFEXpHyfpl
dRenHBZI8XTsxdthPk0lPACyNDoQ5P3+KJnAzQd1xrSazZz9f6MwrLv984LUQT37
BFHp6qwmNMf2Vw1z+x67wHpdW0wUX6enJ4MlenTu+Q9FysyG69lRohwhk5Uu+qo7
IuN2Ff4Qn12OoUKuqBifUN5bbjV8CL8KMJTgY2q0nRIkSHKj410D+L7bXRzKh+8p
vURGkotR5HrhSlak6X9R9jzabcw3ZfU5d8uexzc/LERyvbGoiqPnHnehChzvQJRu
pdyRjhUti0Uqg1aS9hg+sOqIT2ut3whTERsfa8F+ixZ6v/Oj6HjfR3HwhaglzIOA
0LRBb11egHhGn62uYQ+j/OMNu6/K4RofAOdI4x2Z1G27esAG3eQCwi1uoQ6GSjS7
MoHPbUgudZndNXvyplxm6ZnUiy2GXU2Rijse0ue8RlsYoVu0XYzwbF0O35kkm35/
jBv8xeWZTBA7Ntmv9fwOHFjFMEJRsmPhlh1dnd05p9nTMUfn0hhtfqICnwu/JJgS
z7uO5hz7+xcLFfFbjXPeVoYOE0Je0ithtSYgrB5C7sUit+05hEgFhXrTJY9m7z2l
6GoR5wEu/UBLPjxX56AFOaD+c0YMR+PHcJnhquuVEhBxcoMG6zz0R4jLUBDjznY6
yjbMcJckCdiUFv9pJ5RrXAeKcUsA5N9/pphQlReT4m+BIAiEAZghJjai5ASOEP2B
`protect END_PROTECTED
