`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Dg/TRYDYiV5vEkBq/M4kHIpYKwhZE2SWseLAU2+Gob2T0n8D7V6Qeid7SbqX8iTZ
NWnsM1+czrNPedfP9GIM2AHDbdShqKBoyye1JAjWO0JbVfnAaO5fWmT2iUjtMaq6
IN85tA8bbfg3CKRFu7xDxseas13zuJcndglJyfMallOcnIju396Ub3PzpkGA+ZZE
7uo3zRDDzYG2ce3FZyfHyLmqpKjVF6VtFIrjX7rLyYrvhkPqsYnwzhkkhYBH1bU3
ai1VTdONAub97X37jo5JXQTKf4hKrQn0XPMfkpuB+NG+1yu+oMY+VluXP7qMYrbo
PMJSr9mzJShnTBH+p6lHHB+QebFqFYOxkiFy35ZQV1sI0Sa7oRATBj3g2jAFIooz
iL6RySy2looiHfx/6oSofSyfX8tV6ZZPR2Cbk1ZA12p2aSn12oeAjNxCO5xsQumw
np6dvcq3S6QlRZQ8BK5dCNQd4T7im7Deitisy1MwjbBrq6UG3KVyo/ZrgF6W1x5a
PgJvzmry2mHWqbmFV7xG0QbIjxrMMF3Q+ycAeUjLX1n90mnZPl7QKjfJBdp48xyN
Y03rFhpkGJLLJwuD1Hwho+ubC+EvnJS89wksctack+NT9CFxmBon25qLquLaHd1/
BpRpF6kjAeqPbWD5qmJyCCOWJhuzzIXgnVWmwS9mPxfzdQVXat5LXaJk5EhFi2Gi
vB4J3K0iKOjrUs8WcfmbgKkI6wFC32PAkxp6jQD4ptx0cUNXM2ba3xYz2HE1xFob
8nknHLqiFj05uuD0lY0G7sTPv0WIGQA6eiY4PvrnpDv20tmVIYdqk2IWjzLZCM3Z
EnDydFfTru/8FoVx6OSaxHcqUSDdRjHVRvwkjjSnReuUcTIWzBAEVc0nOJo11OlP
wvFsxD3bUfLF3qy4SR7wfIlqmLAM91OxxZpRcqk7J9CCrkvUu7MceWOi2//j4Wza
WQqsnhsabFyigguDfvfU3kL+kGaFZwrw4YyPuIGeH0lYa405cAFKgszpY8sieR6H
4sMWNR2zFIilL/IvD6XvzkruJXHjxOEeATInfTw6wAMyS+C5jDRJERKRUH4sarzS
NHnGl9cwfN64lz5El02MmWlC3B2MCQ2Zguxdr/HQhiyx/RNQ48WIp+KZixIcp/+u
SixfMG6akto4PRcz/xUYguIltHouVpyRsDlIYEclrnIdK9r5LVoWYW19TRHer/wO
GCo/XlKtu4zzRxcpPurFnJc2bPeaVL+eNJ4YJVwQJ0ZJIByLuNdDOqkfiQvMmh8U
RhurmGlZLXG3LjHTWhugecM0dYYuM72SeqsclZs7XBI=
`protect END_PROTECTED
