`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VsfGHHBeCSmvJW8lVUvr27MROvIaoTthPwkWzVLhmZPynJb+zVJ32WxipluRJG2h
yQXDSorhhVLiPahKkwCbkkKAC6T0zfs4HAzJ3r7o1KREtC4jjXVQAR9EVMFn4tGt
Ri5arvMkA2vlTK/06XEmBTsSHLFftvY+Z4FbZszgnzSEN7f28ikRehaBrm9F4Fxu
uKkWbgNVenWtsET0ly1vpRgmJbm+Ltj04488fu2U9HvdH+J4vYefcre7KBFFgFfj
FT7aO/UB1+XSEWCXBo97TefHq5sMsMdnbTvUS8hQiznyiIKlpVH2IikPCvrJvR77
WuEGKt1gHjtBie/mvWa2CHCizGLTYJLLxk0RZarSadYCYytijO2+rg2VOxf7hxk2
s0qX1wm04hmLGpu0TgAxDWeUkmXZbvxNO6ZmPjPl9Ry6I5TtYJ2aW0vL2bM7IUA4
IQ/gvcwEeNqF09Q6uUjwZsXTvj/pp6gYYdQ1vZKhD5gnW223czWxPUQtvCYlglvG
Y4VIt8Fi6kpPm6Th3mZT0sytRhYzNdP7Ko2+KCmHCZLwcviOf3rcZYpQ0QJERzu/
WsSOX2nH9K5aqZqevBvMYU0eQtHY8GIes5ayK4T6PV7SMfZ6Sg/ts64PmgROphOm
Vij1MQQ3LGoXeo1U+ClfrkmLkGJKWASn7ZPMgaKMdEaWuudad38cAuRugcRPaj/0
wSdnxwHGi1RWN/Sc6CFxUDCRW7XYPPXGxoh2NbH646b4fmIyOPWIFHh0gFHdIxJQ
iLnRqWjezbvtof2PT/esJdJfMC2QmPp1gVHRYJlueoJZDiIbFpZWkstoDkq2SurU
YGFKNgfxHBGGWlk17EJpZknQrxRH7SDedbxXEGVios06sffSVSmvRFMEXTu4Tdb8
87mfFmxhecsUycCwvJ+tBS3AQ0JK4C+lafO0GMqDF3TNgVcLFIY3IHS22W6RSUYz
qXOGp9Bn/DUsaOS7lmGj6Nj29y4p4iuMDn0XbUiFHOzK3K5OgFxanrLJUZve0o4g
+QfCWcDQhoa6Sre9sDDBDj0QsycpQmSkhKZ9uUrAOALXyjk4zQg9Qs6VmDJzuynB
6g6zXt1EkC3Xv2Q2vOV7bQ6utTagDkVEi8lnZGFe1HYolI+93J0XqA9FLwCQYSj0
aqzz0DTkGGrgC0ZYr/WDVo4kGw+MssYUBWqTW4rcqgsEwK84rvYeLbKY3BOzli28
D1H9FQZK+Nw1BHbWCFvUHKs2AHiI1pY3AA0IlbkwKF2KPNR5irzt/6nckGqNCnUY
gBt5kPhKOn5amIy4jTAU/oMjrla5cbKCOGgPNl9U1QCbPWlFZOrBJAlcJCaTwD1I
JIl1wERNazpViMmXmiSA3wMvOB2oDP9r+w/m1egHOe9pwDreD3WySXTSJUFXJFTB
iPaC3czc7zg2aoYwh9rmmoCi+jI8pf7IV0wMOnYRCE9sxvP1SUsGMJ2b0moMoTK+
DBOjF5WUxFOHnf7swiU8JoCpUFy4FqACFfUTYgnMfWH+7x2HSSa3eJoY6eZltFbN
mRCWOLbyPFZwHWLO90fyts2R/ACeS3fdoNS4DrIPJEoDZBQSk1sRdpDUDV8m0Fk+
WUxfJhe4y0TwpXtNgmGvJsG7e1bQKRxZVNvu2Yg7ufPbiitYnv1/JN6jWN4mMWgE
q2E3C68F4jsSUIRvzkS1rKy9J2VB1yhWZLWxU3cOAkEjv9s73EthbX893BTaHX3Y
P848EoGWg9OIZFibIwNBrp85ZVjzClgu2bdgb415lI31hcBuhIa4Q/7xz1DDp8zd
agsh8d65LgWAKB7fiYxflmdWr4i0AGDJDY28EaRFiBiee9h+AhiJxOT6seVKoR+y
priXlg+d2X7I7g8npDRwNN0J2XLYmws2lZyXAf9RtB+RL3O5Kpbch9pFLbcRhzeU
Ke2GUC7dy7kXDhdONNK1fydub5w7ZBMQmcGyBvYkZt0O8nB3KukFhbhleKgA0kMX
XwhXb9wOfrjKDOKNH64fJnHq6GJacW9qMH+QdXka3UAU9jylJWXwoQBy9V+FtVat
SXShbshViLiypoeMr4tBa+s7jUrHENYtYtSyd1fvbwNwycYw1ZY3VpI6gnvOO789
GZHOA6Nm0E0yoFbazs+J30wWR6PH7o4Y9VUmmCj5jELaILbsCGHa7lDu8cuo9JQ8
0J3uF+G6SmZnH34jc/oyifaJ2LgeneIKb2EfogR7XuQMDQWuDhMiBUs3lpg3MIvu
r/v2ibUsJw8FuVWgq9cC70A9CoZ4R1kYeSNukmD7nlHtyPDY1nRJwR2OTwgdo4CR
EuuKGOOhBlfDd6fxHcfSQdqNKdOZHdpSzeg1ihkAWeZsMkpd3tKQe7x1BJeZ/+UM
UpL9gs0T///+tzoR77FdvALXwqXl7Tck0jOexrqR7dJNziUXoCaEnm3kuiSdVjzO
/kb9jLN4uCDAzOVi0TaQW2fKsRYZrjW0I94CUQYeX/ef2XBf3l8w9Mbgg4LIaWLN
ZmF8rU2yyNavwpPNAo0vWog7cGviW1dUXbECniqa2v7xh8xqt+HWsMl7pdLy69HF
AN+JRM1fNtT2ZFREwda22uC+8Zv29Fnwxi3YAJZsr17Xe1WZLaciwXBm64RWUpJg
UBraUhDmKoxtLD2/KcRxq0vdJ26Nc8maKISokRdNjRlFp9C+MErJ12l+/MwhQohm
xiQ2DQlqNWFsJ/VK+20U2SpH99G7tCtg4TemL+VptTEVkzmBxS6Kze1GhXocvdFJ
CF4gnd5G5Kf5uER6EjD5kdYTUOVKytP0Z9hx40rtec26kOvKKdAgZcDZ+r1LquQf
7ESsJqBxZJZ5iWB82vyg5dgOekkmiQzgHi/eCvSBZu2onuVJPpvAIiqSCJV7eyGe
fDpfbRWAuV9kvtNG6ox/7PyYKh1Kc5wvqtyHROXVAMuXJQu8VveojokBrL/9uuo0
aa5gZaVqJx1JijOseX/OoLJ/KS041wQcsINZp3767HZZLKlNtoEHlQsG1MMZrG+Z
Ma8j6NmZSmHy4icbo+3wSTfzF1triUYKeqJ2FR3HBtuh7RVpCOzNxz344UM+3/Lu
lNMrLaIc2hjQW4A3irEBwlaNAuYXgAi+nBrb3Duc5Ve0CqR8vHW7AjqQs3/CiOuq
aTyY6trHyEsgfrTpTOlo3KF/Qz/OZ4DkCM8JsZTCXT9EtdEYuv2YN+s8gwIBRFbM
pVe2C3YxVLBIFMAeYkuRqnmmydkDON8Jumb2xmgp4TgsNNJgnu4nyt6rMXdIM2L1
8IzA6b0+z2fN9AC6AWBcs/03zHAPI9Q4sNGOLcTs9OLf3Fr8DVKWtVQCUpglaoV1
AxDNSIzrTGI+CtT8BXKtlOHYuhhgTC7JoKqfMz7y0pfB12PNzQnrqNJBKmbJgyBs
EDnRtI/ici8Ox+WMMg4CisiLonGKKyGmtz65dS8WOa3eoCYsVRzs5LKvRmKRgT9k
MkV+KBtt633klsDsT1uYmdsG3BHAikLIRg5p2h49IxEOedyXiCSRN7rEVGLaZLGt
naNLpr9eJC5RlaL7aq6WclCW/iuEGoaySVyfO1XZsEFozT4WBnSK0OsxVmaPrGTn
MACHCJ9rz/YB2QVC5eHcN8NwTp4BWZ/jlqICzlDXdwfHrsueDBDFezOSDyk88+re
qKPjZ9e5fQUY/6eu7R6jxXv4d6UjdLjfynLysCOjDQYvmbng2upr9BnM5P/3OPLy
RQD6mM2wEt044YN6XzxMsyyBXbiHUyfjmomKZ8zOyd1TWB9QEaQEgnakYVtWj2N6
tQirjaQ0ZjG4qAnXsXu9qUVamsH77B75UCMAryf87RXWfMidMX2RCwpgb0pJiRuY
L+S2MajUbbBkQGZXTkn03CJ33qwPZnPK7N24x8WYVOB5A64Amo4Pb5q/tcRx8nV4
9/4lAvpz/wOSiMslLiYMmhqnOAG46Xf+GOfs1qcZfw2GEoiuB+p18Y6Qd1KszIZq
K7Ta8JMFuGUYlYxmfCXPv3JaxYN1AukoJ6VXFNbQXmQfxQ1JpTFPmCWRNV2L0xNI
m0hg88LkorOr0g+uCp9uUuXuM4IM1y+6lecShdAKxb4wa1stAhSWfwf0Uo3kGssE
PyM6ddvU2FEz4hWZWHH1ZJe0zRIwbKdR3XQ36OrkkvpMre8gjRaSYf4qnAn+SN30
oXhzVQCEocNVsJ19pp4MrZ/r4748ekx8w6746Lw0VEmct2x1MJX+jT3sQHp16Rid
LEcbpNRTvHmawjUqlyF0S6UDMDlvNo6A8eLSYkHVeASNcu79G3ynqabLQSgsBgoh
7RXtxSI2OqNMO2XHwh9hAyfzLl5KhE5vmbYOxt3esDz7WwD55IuGljzbnTovJywE
ax4HnD1RfsxsxuX8ad/NGGOHwlK3u9YBfsrEkYVrl86Pg4cDIn7evchNn/Thq/X3
iW+I3gg72Ix8G5dXMYgIm2oT/jpTHCo79r8mnDszRNdxXK3hAAeVm5b+ptzTooWz
eyO3rmuuzm6tccMr4wh6QtsmJs95V6ha16gn7IY/6yhM9Y8/QgzAexF77glbJ3hv
moAyTUZVkMhNfmD+9vgwPr6Yr8P/KqsHOI2TfhRQS6RRst7P+0wStnYgqFLqsCYP
YUUtnX0sVq7jL9noeHvpa13xD/yk2dxqN5VFTtnvczbXRTFpUwYWwAodvw4fjRbV
CkX49ezmG/9UEEvArnjVilyMBGxRynsdRzr7LNev6ETbYDfGFc8L0qIdV47Xb+8S
l6UDttwlSRuk1Guo+RH0cOla1JY07e1WdKMDOvfOGLrDnkSpBt0pfDp5ndYG2xaG
RTX/VIBUzVxpl2rejoO0/WPTWRlZ1OppUYHjZJq4ulnbAtgC08pRH5mmrzeHd+gB
L089lX3VbQdsQgbAdSCdIvPguz7aoof+REfn0/agRFjN5UirSP7mBI6A6Ww2/+p9
wPgfRPLC+rxftR0apRnOVGUqSAlnM9lq3Vlf5fkxmRn0CCCFRzb2F9Je8pUgB9up
B8Ui/PjYOGqT8Hi1Ahwl/BlQbucHRtfjIy5VPLGyuslRD5HVKu/vH55Sb2mdb79t
`protect END_PROTECTED
