`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EOSiEyQ0vOJPiKQXvW7YdK0x4mECo4/DxRZsXsNB/+bDBcaAfHGbPhsUGwDlfesJ
MyuOfwXZkUmppq9eVA+6VENDTKzOJJrbqvuaCie99ToqcUhe5mWUrCP1uDvUU9sP
oS0c20hPuoc+n33+savl9XLUNzOGS2/MHkRasK8crQBrESVYT8ns+K2rb+wS88vp
1KNqFAavPkF7acuYaIWjTRmwOdMbO5GRu9Wb5vJo7I0fAVrLC4COE8Su4SXFkFdW
W7kK+GurB9XiHn7yZDakztAevtlgfOJhpa1R9F1Pev+GQXl5Z8haZaib4MaFKeuw
gj9hgMJGygWHuHLTCmaV18cHi3DGerAzp6NXbaHKJJ5nT8oUkf2LCxdhHtemCekT
m2ZaEfPrDqJPpQ37uQ3pSadvUufs3mij0TuGvJV42ZDJUtgi1L6EHFlBM4eTudiu
tA5ez8VanO6o7DEUC8hBpjoRsgeGWGOjAd1eH3f8q74kPcH4jCzh/yFfpsTlIA7p
06Y5Qrz+YrMTEl8KXQm1Vu9zzzx1rnVKSw4fvxXlw+PThh4ULPl9ZcBP9EsMn6WU
pvWVApOqZnH6XV5NGuw6Ges14/1MbY7yigu2Ylj7zMd752JSt9SO12eYsf/6xz0K
o2RQzykg/FejyClAR/QVDv4mgJXsq73hkhe1G4U6qwMRNZdZHyvDV2rHh5MSNjlk
ZZnKPDdIyrl6IhQj+t3K4iUe9+XeK1OqLKAtFWltjrV5RVh3PJzJf4RqUdYK/bGK
`protect END_PROTECTED
