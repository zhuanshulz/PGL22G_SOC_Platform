`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T4jNFCTXW5AbyOctrBCteJ3P4a7LowguHgPTHFZlOY1Dj4lcOEzPuOy6qK5edZXx
/jBD9qilniN6uraFGET7Pr8T2gY8Ay+y025UCtjt/0u3UeM4ygcZCgXMSO1wzhTB
70f/EyuMc9vWgV92F9SIPybBZwAnpjYDgjvp4gY1e0fz14JnTsiGQnoUaXKRN7uY
HoxMahLVN163HJhnsKrEZoGOUHNErbPAFqCK/fFMuNkhU0/ujLEj1ozDPtGDVe6y
g8XLG4c5QTI3U8+U+yTvsw74nETHfe9XQmkPaSlTsBEExTKLsLr37xqBwosFEBto
OM1iLDYqn/0G3xyIWQ7mo4HbPHKPleKeGB71QqcThrZOuBblRtU/2UoSfd/eUwE2
mkUMJjhLZRZLwDnssHYtdbwD2B9jcU6nxnTrCQg9dyuFx0gt38Xa3YTDWJbnBwu/
uVvpfdsJbF3YGX42DOy8NLSp1XhWke7lpcAl+o/CRQLhKbzLlwWRnTmdBXQfTlaM
eZq334t9mfzgUAkBk4p0N3pL0ooZDKhUHYsXRoA/LEqG3CcK3IJvj96P/ElsV/vv
gLSUO4XYsDHcl4uGhHdDSl2ik9svpirIK0DHy2QHdAhyijEWmTTUll+XIbL4XdwL
8fCM4Ey4h70lbAOng4+ITQLvr1kcL6eWUBquuJ2Dzv2s/Zyoif+ZWbyA7jeow0/y
AVelTcpD5RNJOJD88ipcTkh70uSnFYKskRRbjDy5AtIb/185KvI4WL/Fjh+qJR5s
Mv5NFUEJG9tmFe8uY3CgXO78qLxHNfRRVh4l62gpiQO/h0LUWWb5tCrGcLOQpuOo
4jxKdVQcRdEzFN5nbm8h1x+SnMaBEd9vO0+ZD9kYOAggqoAC+51BKSlvHts5EvOE
L0B2Iw6IOQUJSHMBekQ0jLMIYeYkGB+HdtKiS+g2pmBTmaSXGL6nYTv2c8y91JKI
EjSMILWn6kdNcUw9zL0RerarJH0O//0kGo1nGxr7gzr5vTu1Bls9Bzn6GY5iuAri
A73238MxzZrGVqSVyqVBU0huNqcAL4hzJ9sCMaNBIQ9Mx9B86Srx3Fb7PvAdoue5
RhkDa1sS+KosD2dehCm1mJRRpyvA74dGKfI2SyGP6YxmBOPKEzo2sEWs4F4SmQZG
faUi/TlY8ejnoy8XtGDi+pv/4LCpcY2122dtk/doWkBPvX7ErAPkNzl8tD5xMSL7
bfoZRaOd0uhUmCCAf5TG0Ngl+uPvwDrGTH/2XIWxvvbQ/ZiDdMznsoi6BmYQQyr5
OcoRBFMMp3fxyjqGshIPjmEK35yMAGgW7vu82m8h8Xwf3bdJaOScglBl/J/L9CoM
UnH/VxLmQyjHTkXtgbHTWxViLQs5GDdO8C3wwZ9IcyIk6jjwabMc4EsYGsh2Pjzj
T5gj5+Sb6EF+rN36kyWZC4cplSRbSAs417dRb8iaYLsOMvxmRGmg4wTVs8RNKqU4
gosNlYhE7U8zr7o9AgjsHg3+McaV1AiSMx5q9B9e7VyjPKiSLpD/NV6mG4xjDGwB
F0LCocPWWuyVvxrDB/5M8mt7J7N7idwOxfOMvU/AI8B9I6coXhO5U6F82C/q0kE4
VwNJqHUmi8CA2gCBRpveDh53pZUUpjjLVY3yHVPrE7HbP7iAwSr1428eTFdhGYUB
oJDnpBmNZpL3FDRn+8x2vPAAzxhDEZvkioFvOA7hz+k0x4tGU3Ds2qh4/MaahJt5
1CeYBnsVAFhJdmcS/8tESUkdX95cj7XHpy22+2czkMrMOrkcSSoy245xHYaAF/38
6r1c43tfEHMb8p4m3uOGcPZRSypaDDAF149yympnPHtxLklJo6yQskwkR8U9QR4l
lWLhT17T1C/I005U7hBQvDGQ1xYEJQYj6I+g3V3Cgbw+Mx/GA0uqnqbj5aCUo6e8
P740D0e2AfvZGmJ95VSZL0NRh3Xv7d0jn2aDgIfuJQXMcpj5C5XXxGKBwwlpFRT2
lpXBCsLZc14PefUSm2QDHE1IPoqTjVCXjLn/9ljC+6MyzN+nlULX9E6mK0kNuC5E
v6UM8oNYnFORiTYV9HWAU4twOshuaEBsasRZL6tlbRSTnKlZBZkqvpjcRP1jePRT
qTG7GtmGj6MARNHnaJ1h3vEeoteIlOxbGQv64u9eq5aIfopsRGOxTL14gOdUMPvM
8uKFqI6Q/3vj/GwVugP5NevZaTdGD+CzngwRI5hEgHm0haHE+81Dwa3VHQUaztFR
ogF8gXMShqiTeJZlI+b0kUi/UGr/8JfFIsRsldHrzNT5HWMNEAWTwhJLcZI3jdvR
omY0mcQbD2DgNbfsCXXfLOcGgITSGULw6ThO2xopSdrG4duCMoL0tG8ixKKbchBV
SctRlb+thHE4OPR56Sd70MCpImazLI0ATwnb5kC1tkU6xT0jPodJHfHoTRuWQiQ0
GP7qzwzLvvBVEiqrPgZVX67uFVCV9S8SoiT0v94g2DA87WxccsKehtYNro1o3egx
X8DkH2gc+fbxYyaDZhAMoLGcJXhMzfoM7bF/ckNuFwZGYLY8zgozNSAxYpZqNAX4
AyIAX7255xdFKOw/QHt4UD2wraLJFrHVEnQmm/JsD9XbNp9GUdkO75S9UtRKFHtl
OVFuBO7FLQFm8tA4SvQeZCYZ0bvjz6jAbDGjI0EO0TcIbnxRo5PKW+3IUH3y9ywu
x8X2IdX4U8YmsmLRNlTIemPvS42SBulgOs4FQZ7XUaB+Vj54cY5POtUbFyR2MEvJ
7Z/FroGWHA+HLLxR0iorpzraPPVDXp3VTft70kVeQLmuv3JWwqtcaN3pzmcxigUQ
y++tFWyPwvcWIuFEKKhYckgvxShVTgjcDkQy71WDlx4/D02AyhU7ilB1xqrA6cOh
0Aqm4SARCaOg71putmh90E15D0VPMpv9Km2/c1g286AaOm2zYRrBEUdvTBWN4T+i
f3A9KOGQd/QXprN/vTZHkPJjgMah/AFxhTbb1srK4cYV7RONtJ9x++S472/bakhE
sKGwQB+xPQdTjv6skscXsW2Cmm5JsQ40EJDfha+UZLm79n9/zFgLWD+QdqB/Lx4g
uDP5/IdSuYnnnNvfscCArI88yK0wy1DKZAKQH+4oulCKEWza/AXNhlRMnt8M4rEH
3AdLEm1qkM2oy4OV/0qEbl9M0iM0dHALQOAxxyimHv92rf5g+oblABjMqVOJMvIN
RzNR9p+gAPWhLWvYQ3+xQCD5Ndb5Ipw+6zSHV2Xp1qP6eLj9BqE7w+CzBQmqzTcj
R3QeLMqKK8+vR9TNZr78x3v6MZrVXUaRoJb1raPFUuqI3BVWM5+vJuVWLu+ledvA
ME9J8HGizrnAHFu4CaAIe3hewGb/UFchYIK3AeVMfDNQz5CoIjaNhxEmfRr570LF
ulN3W97wZcV9Zplsw98Hssachg+VW7r3wsIHoLuexJ/kiia4ZPekj0+6XVmguG74
uEFpMLKMFmVMQSyWcEmH3cRoAGrJdIwwnKCAVMandvfqywtZEHlmCXe4uqH7awW+
Sd08vuQP/x5OSDOHiMNpsRv8rT+BL/jdLGE9yk8yMHM0oeqHLl8LG5WR1Yahubb8
Ht6lBKRt4LiUK2d7zsTojC1e2gvbpTuKPM3BEkIKbhYR/Hq+VTdrv1Ux4nRo//WW
yxUloB7IuwnRJisVBe9QZAyNYygG7pcnd/xYG4QD/GtQdKaauD5AqLqk5QCso+34
NEMSNmvZaL+vDetQOpb2mYW5OjFKJjjRKCiDGnStSEaFA53IJkgBP6fTpJMfubR2
qa/ldYaTo0FfzlgNTByjMawOl5EGVULSiQtUG21BcdCcSJCe0/34KINnU9dsz9do
mFPIGJilD8vP3IeB6UZXKXR1mYI93z00KDc2tQS4oTNXDkaOOW30TA8K/Tl57O2v
4J7QxM+jbD+WuwgA9iZmrc4ATfbmLfOBwy06vSTvTPmo/kLiVRoU7f5ioGYkdZs+
xcMOsaw5GcsvNgqAkrGYgLsTw0t/K5VyKHE3Xz+gqX9+TRHSsrnqh3JfdFA3PMAy
TUz33hLszhIMMd/IVvzNEDBdynY0DM/ihWP92CcrWxBUnICttjXp21SebE4tnEeJ
vfJNRSLQAJhiKv9urcDRSbKSwfXVXspKXGkpREZGRqodtNSsiq2Y5/OfPR8rLsrl
l6NtC8V17HDUaaAj1mTQ/Z0XaqBLOy5qjNyj91RYgIhQ3vzPU4oZDZrsFNO8k8XJ
P0+ki9XgkZRjFXMYhnue1AvSkCqU8Td6OkJmvFcJ+rIQY54lVCeGtKGUWjtDXUlg
K6613Q0meGp/RH5jm5x0VBdwWOcHW4ng6mDGzxmJiy45MA3DHkr07dLoKtUagXHF
aFTdANUZqTj9NPyP8puqsQpbRpHVDNQG0n+WdrYJ8dQ0XcIV+rAVG7Jt0Nu99RQQ
W4rDg/RmiJt1ioDr1ixQxgrdbAuj1YslQj9qheu2e+iNLhUxS675fsQxrpn8gvgR
ElXRxYRYNuWg9Q3I3E32NxewfdP9DKMz7zmKg9+kdqMaEmNshRc7p461gPnk7TUC
itPq4K7SsJaFgqqPnDcINoDV9nAJFJrsmWUIvhDGHScFP3IZ8rEM1MCCI+3mUu10
4bmetd8RofiYoOlcjAQQ2HVPeCAJCGJd7UT3Q26MQvQToVwHwJ+UlQ4BEwCWubRt
FYDzNPfZ890Nf2zseyG0PzzkW/WdVOFmPS2tljyuHY5u2sCo6qsYikqj1gfB9GTE
FLWusPRFw8nfWFPBtvItRz7j/aRQ3FQZX3EzAiV6uesPQufOVy6cBCJV5Iq34iWk
rdFkzMPl/dPLytZfTET/EY8Y7ibmq5VEIaoJ1xz/T8DkOYQfiDCdYg5WcOGymlDt
LM7OlOwL0hU6P7sDprMtUFO/6XbBAWHqYQZqaB5BbOOL1RAfnmbECcAeptuDB0d0
JZw4N4Z7gf3ikOpARW2fElRb7ORNgFkwR4CDCDEWzK7SKRjSBtWKPhYAZKKkAc6I
1AcMvSPgx6TbRMF+NDlU3rQ/EXFd27STKMWoesoEP033E90y1Cg8Z4sFLA8LN/NO
FJJzJBuT0HkXbrQNOYx6aRyDyhOAIrf48aRZKZGuLbvRotXooRAa1TCd6FGR0u12
m8koww4knCu07YuRlZlFvaLY9sALtox+pTLKgrxA5BHdY9X/TLySEhk6LDETelKI
bv3+KLTxrQZ8drkOBrTRHbH3aMpdavog31vSrgASiVQD+8zVJPBpM9Szc7pi7vYu
vEht7zJ0uzjMFI9c66PoeW02+JGm17jX8OyGSBQHGCLKqqEfnTfQ7DcL9L3GA1GV
MB0GjoBCo/vsOZt+WqjtY96oQEz9sJPlANBVympsJMoF8zV8ndyJrK0Gp9ofyuu0
sBdGZwlJ5lf/iljhPKj9nKz0GzoCupiFordziEYrqhSWX/aCX0OW68Qld5Rvv1Ah
9NAcih2UqfEHS+LXy5tVsmNxeXRG+ZH+u5MJO3XNQGZ32Tvf762pfVUmf7nApcAe
EGNc/3mZ43EF3Zxpgbn5w39bvXJmKv3k1ALtb4Uq6UHIjoYWsccOxxUJ4Vnq6GoJ
4URRzDKuwty/HdMLtoJuJ1wbgPOk0I+Fb+WkhHGZxM2PWbzGhgZV+95BtveWggf9
GbThi2ZiqT/QtzMuyyft+t48Z+XfFdYJouTW2Jt0UoE76qC/YbGNjxA7s7vsY9/z
ned1qLPZhX5YAK4dDtFeL/f596+qq1Yi5pe0QdJ5XPsbvhRUE+w2gOhKdAKYgsnR
DscKIvksJf6I4WP2Paz3L3TKy2xzNU7lOI/6aHzt1+VafEW8Uw9g1NQQN/kUOlS4
cdu6orvvI0n4LMJIoVq90/x3KdpHdj/uWTS+4OgSL+RoYUHh6+0s8paejWz2MLf4
hAeDdhOcs8WSIYhPh5v97QY5LWRc6jRmWfn52Znvv9OA0+1ZnqbwesdPGnV+sBZK
4u1bo+XtbM9DAX8LDbikotcQ+PIZP71JOtEBE95EOTnu8LDqMx1E5KRAAtgzdOwK
zBU5vqOk4tMpSB1uRPDAJMXX7AGs35o33tMgxIhHkVj3cZ41i3qT6tv0s2hKA/nR
sPRb/hwtinOIbYDnh2N5cwixbtBpnvBNyAXDx/K1TiZ0IXi7Gs/xAKFb6/HaBNsU
cG1Dkjo4IMJpVECu0nxuQhA0ZR52zWtYm30FP1dTBC3iQcCYE9lZF5jUwphtSPth
JMaBhYgJztI/CcOqka7hNFftWxJ2sDbqbB8YmJp6KnQq4nAGkt1Kj/r6L5Csd93q
FIEaK+pM533+HkEWWr2/oh8CHtbleAXPsR9V7+Vw4nx7XGw2N/sJ4fq2lMbzYELB
Fo4g4v82E5unokaaXUFk6MadyZY1/1iXCavnuo+zyb0XcNhvIce7ys04Tbv/LCZq
32m03FkLjpKpGehmgVTkIlg62tUSoJ8azRgjE6drxSN4Ml3GIpI1UpqeZ7YGmwc2
A4ktCcuGd7dujCVCHwAhxZpJ3U3t16bCSpIQ1dTO+jVczIjFJU4WIUTeLWPwaZRo
RvX3ux15WDNGY8Sf9N93gzxkWUKn7F/HaYYpGrDDOJqPtKAzog/qX6ys/rrHik/T
DQrGJ36CqewbfgO3niC8xYLFndnZpyx6OlJRJ4GwGIKEq5fazdxz+RaGM8IPjtJm
RiTyTUlobzg/IJSo+ObPFKrmhUvVhGPVn1EjuXUAKM7aZYvU1/7bXtNPr/vdVvDa
ZZAglQkre+CzKh/92G93oTBUzWmB/r8QSbiouU8hOIt9ZGUnAK5kULXpskL9yWHl
0j7Q4ddSO63zfqMfjq+WQZ77VGmlxLfD6/37frmrHl2+M8b1+5Q3Gab0H6ScLlyP
GU1L7X8deqr3FNaMt9QTUTnIDkaQTp6bvjB3sAgiiucbKRajs5rC5wGfr7vWGCho
36m7z1aiEz/GFNV8x4vvDUID+axmg+GPOamdivNTMBkKw8mBkcQiNdOxwoU3RZ4Z
x5SbCOnE0TQI/wteklphO9zBshbpXRzjQ33+WVMrC5SPEauwMPzuhnSfkxJbqrUq
F9H77UWNF7wCXHCdBs9k0T6Xjdmwqh8tlzl2XJt6awmCBCpk1F5I1ZbTxBo9Yiyx
9o80UvNBBrdxEcPbSRnOON+RykSOxEasyQjZBQNvV5KouzADbM1/8rOIkKDRrKrv
JOxGFo2igFc+Qx6v1I2CmnCvGm+HqlFDuOfrugQOL/8n76i27JroV735mSnCboCr
leXSQcfg5KweSiBOU4qN2zp1YTuveYXGPskX4bS2aesE+DVVBewlDOrMjcUV1JYX
LUEFD1cOiEw6VzYjprf4UxPoBI6GoLl3YaTHB46iS+afe7t3ZX0gCt0H2zvns+Mc
tLiaViwqBfRB6L0HB8YJiao2ooWEvnRUPhfCpI3NJeZQ9EjnDI0t+sX4YQQ8WIl2
EM4MjX2JoKB7+uz54bvAcNiC+YKtrvz5Kt1GUKJiG9KQsG2G5y/FkBiUtHYEHNcD
BF0HYXtsMuH4t9+c9KJaAQBUdRxTTGhVZS011iBLMvJGLeFz9cRlVMt0WCjKof/p
sWQlu41JQlOpd3tLul3egRtgOQXnEnGLZsWOIM6MDphAYj8NZAAX5vidLUAImDHQ
rfr/i7SZvUSy+LzraoPB3jIG+G2OG5C69PmsjOA+2avv8bLHonO0XnA49T3vGIxj
NbczMqVASBbBHmKmWMyXD9t+R1k1X0NqPXOy0vG8SNiUkI1vbQ5bJtNvKkRrr9rm
o12F2UNwfuLnYcArdXsBrjjJ7+FxWURwIeapK7n4Un2OTsCeUrolkqRibUi24tKW
Vk0AxNJflnylmTbRAOx6tMz5oOQqZNLaCVtdkeUCRZgubaxLhUFdujuVUJrcd/8S
hMxxO+eERrcOxYaAXFkPr/EqELDR0MdUwNllU9bUiW4IYjLLfceM2uzbuoBA82Pv
SqEniwl/UF+2lzF0xLQiAwZQ6dtvqaBGK6tQ96POgDqQiIaHO3eoNL9rcGUKSqBe
5OyeVezWz5X+LtaPytj7OBbf/x+SpplhikQNBFB8x97Y023+hTX5qt6D/5LpTkrJ
pV4Ay2UoBTEnWN9XXR7/K9r2stWbC+Mo9MS0ga+MMZN0RiBcQo3ZzACIngvPyY5e
BRnSbdgoDe4sxu50oSV3OhaoPK61UYskpNE54Nc7GJ25jIS14QMwiJqZ4b8kNN74
PQwMirtNQh+SEKZSFPdbn6S5cBGj4I8/9I39qXDHGWd6XA3BfZG1WxfD92+tVNdR
AOBx9eGd6+CeJx6dSKNllzH6XbEqu+tYbCYKPWzd6K6mtj6KfGsuT/PTh/DCZfUF
iUvf5imB3XhXXOMc6yw2Vmadk4XTlgcnqSLj6qMa/Y5gslL7HfDNGVKqrpOzyyLp
Oa3VfBtlYJ6Je4BRze7ai8rS3s0I1zJFHCTS9f1Ilfdj/ajz6NZC6/dnwSeC4vPI
ykGqF4T8eRA60iocykUCbnBV6hPmrs575hWfakUvA2MuPOmFpAbejzVODsD0p8nt
UmGqjqkNrJdrItHadZk9xpbBqAYbF63nuDobhcF5Wdap4MH5B1udsYh3sUFQ1Ibt
ww/LTuCkPrm7UsbCvNtODnDuBBazNE1MMEuOGdFBY7L4lkhx/NSdu4XTaUUylYSD
vwyynqx3ATqm+2VtrCoMPZEXBStAuKz+JphtTQlXyFbCph8ehjVMQOgc3P3conJJ
lipkDWibFL2uo7dFJ2v5EOEwX6FFlNi7ChvryQSiBAUF6A3L2QBMpjVm+++Z6L3c
HvmyEBbo80FnuA4U0cuGcthLwWB33sGJZ2OxtpbHI38hteuDydzyxRSSnlCUV5Ge
CmyiBUdt5lTt8x/mtoQcbyMqH5drDg4vVvfD0cEHdXQIVmoYyokMpuHREr5R67vp
ayqyoRsqNBfUyqKgS2n7j8Zo+LU/UAUzDnrH5J7Aol161ZvV66VbR1ponjf8xN5P
yB7wMWS1p7MOBrVDQVuaNtg14pU+GZvL5L8gK6OZ3uQFAD5gTStzRQWc4zUQ8yDT
JabDLOL0lQ8F10xT7zRdSwRROz5hBxDwqG/NenoU9n0crGVZylrnm+WmgaUafT51
QYNPYEPnyI8rxyF5otf3ge/Mw6PlvzfnwPoLVLhDlGXFK03XFL2zpS07hAOH05Ed
k1fxR1o/uu7oob4u8oBxytAEzqc1eIydpwQEDEFFmTGdlKa2AXYyEPOS7XwNm8FV
TPFc5qXVJ6MMFImSMPwIWQELuFU/e8+AtS7REWAkZHTltYP7/oy2l+GPqBVzPFuR
XiQEaWzSJ8wSq/yM7cVZNBgCU9ircmlQM6OznEtx5FyJuojTv/kkLcT0/msQR2Rb
xi9mKSt4mCWFlFxcNEiyy9YhAPuYzhRvNvBPGkhCFDa5SEUUCj61r8HpaL6Cg+U4
Nqtj3esELRYtYOTB2cerIUHdDdYVFksD8IbOME2PdnxtSaI3nO9R/+WuuveOBHHZ
bsspu/9QJobApLfsuQsmv2TI0uQ4tcZVIDUM8FAXmmo32uu2xRBL0JiDVuFIBfRB
5LtomLpWsi3OjT74REB1lPZbnW2MUXj6QWlhSB1HhKY3jYGorZOvsPIrFB8RYsIp
i2fhJYw1hvJh+7IA1ATeFrYTbl5yqGImPqWa/frNpPPiG8aRKB31wm0w6ZzjvMye
HXr2DklEa2xZFOadtrxxt0U5+LmdELn4Vn3qip2TPxlQDfBoSoGdCoOmGPgaL+WC
Jve4loyPPuq72vxVRYPMVT3qQPH/CY3/YheCgbWDLC2iAm92ttrL7RUyXjX0cISF
jvFnhZweiG/kT1ZERcgvFdTOyU1X9n8a57SFETCKpvmukC1niJPW5efhVI14+Aym
Xe0FFdIrjTRSqDYlveTtml9C7WJuOt9Z+xUwSfJKWv4naZT2MAvi3WLqhR4c4wxr
p5OmjdXXrEBuJPl/wEpSMmhdq7Lu0cGFIkTAbTCIr7wP7icgxdoU6uazpPzHVZJN
dme8hF7aXZVQuhE5w1c/EplCr/INDNTLDUezoCohxjyaMY7OSjcih7aBK283+l4F
yp5FvnFpiQ10jd0/yRMn/i9/And/LWBEj4ntXh7ZLpDSHVfuUQF9sn/c/snPeqeG
j+DnpUF5lb1JQXh/VtqIXUNgsb11J6vINGUBiFp7XuNY5z4riGM7lnb4ossIRA4i
VEKtmlrpfHTvqKgdfmG9WoMG6jpruJTdnEmNb2jomZgID13CmCIAKfcV7taxYHPX
5fpgP/CTyqlpqy8zurKVyKpo1cPx8Tk7F4XHEtxIudLX8P5kzKJi3OgDa0lZyVp/
/QxbgBZNwp1ubska4Z4RMNnJP3/zUsBOIkKYFDd+rGrFycYMROpNEFr8VOGFOT0G
175ilofPGiv15CYK3Lc3FjLo2KNY0rH8bZhYXD+lxywwOUsn5I0I/UKXSClpoWPz
ppyXadlRoNuzYiBhPpN/jGdkMG43ot8sQVAgXmG0Ft6I/oXaF+0mubNbOI+Trovl
Bi8f1kzhY52bGCMdjhXY6eN+awKyp9KQQM64E5vjBaITzRdL5We18Erwl/6tT82M
Fu9PxLJCWhA8/ajt6cyVER+yFwer2WHoLwHNfCo2PKKDWlg632AYpGkZlyJWU7HU
6koxqFhxDB7cj9hIr2uZ/708QEl6AtHVn3TvH1yuIhCj70E6Dp1yo9J77r1SHBgO
JsYrYI+Db0bjfi8QK9a1qY1l+CLkJBJhhJt1UbvT1oESX6R99OW0L2u0Xz/JqjTu
uJ/ur3TaHNdkNXg+iXSuQ2CZduyfSwbAWnYt1YZ7XAWbAPtO1xd5S8mAS7fIpjo4
CKC60uLacN+LMVTiDqQMi7zDZqZAm1PcP061l23SXHxnmq8DzxDSRe5uloskJDe2
yxwdj2v1RdrHMb11pSZIs8XqdL3xEtOj5flk+UQXAJZg8RDU8MTTRtjB2+e8Ca2u
slZ8o3wd4Qoit5i/xF9LKNC4QuVBukx+h855UCgGKJtH0ZI0kz6QiKVmnqEvxpF4
5S/3h2oIlKrl+yqqugR92d9WV2sG4rXQCzv3jOQ0o54Zx0w3GWGZwpyaLyaA9D6L
vB/Q2cefDJ/2gw0LnLYcLgFmsQOW/vzGZcdOziKimJCVfNI1VwB/DjCFsmAQXciE
R5TAu/Gue1r08lh17sdi0fAlCsp1y+88XZNEf6tu0ZHvIFYSZMQ4KC/zLwbX8NDY
ZVut6BN7ZLyXvErFqxrU7kxwCjPO2edRXVowbwCVBWW+cXuNLmHzmTYI+Hkvvb2f
P9OncGdnabV02CamjYYDJ8T+wVOpJOs2XPaw6hmHzKNfUgm+JATbqpepQXGWDd0h
V1xbxKCI9OYan5nKBQH16yp9qzFNH1FRy+9qYyYyU6R5aDv6ZdwAcHTKWArdsyou
zNoHlbkoCFOaSmP6CFtvJy7oQgx+UaEj21l4F6vG+5JL5Ew3k9Rvjar5HG/77VT3
8SrTdhewWD9WH+e1z7P1fGPh9Yat2Z7rFjI5Rt5muDvk7vZ/XhKRytCCcPnBpkMj
P5B/5XeJ3cfrDeuPU7tfA7n4H4P3YxoFE9+J4KEWqtzFtxsfTNI3lY4S98p9K8UT
Gy1E+lqJXlrwAaV7ifTnWqxD359IPLCcy8GjcT6cYITToFERp6a4zJXsKb9X/lt6
e3wW/4tqI0HGQOvoo4rtLCaTMP8ukGIuyp8OEiofeVg53VIUTjVUoKpIJgzZe3B2
voAzk8GHAZwCclqCjzUNbdtNDv/Klq8t51pbDBTGo+bwhOeaOyW1tOmP3eEOtBhb
oOdE5fzdb91e6ij178pREDJ9IWyY3smV7yo6dlI+c7qmMEAijFaUfwk/asla1L7p
lSfKckV/CW5cq8cet5vpTvbkIRDFX8K/5/kZlZoedVgLtii/4eCFZCfmYIdkwFhS
pjR7o3yz2BUopmMKMENXV8ooBtSMY52e5RkXwHfso8rcEAk308ZnxdWDNFcVRX4R
Gy+0bl9g16ho+8vKcmLLhLyYpn25aoGL0zHxXLI+rdixBr9IPiYvcfH/xx1ws+Qd
foSmQ6Ahq5yNIx6n1w6nO7twZtax/5DsUVhlvhM5TFStgXgE1ycHQusAmScomEWv
k+yVUUXKTr7H4kpSuSBnXcEew6seQGUXPoKATc5tByzag6iqHU1bLECC/XUX1ndX
Vs0QaIqn+Xj2RS1ebX+o051jA1HZpVydhegwL5TnKdHdTtZGvJpPnIDyeN5YnSGw
8auw+xTlJ9s7w0LTsgBaeIG9RNT9adXOP9VguUMAidK3+S9lygEZEMu9gNhq06Yu
qyr62To2kcksDylYkhZljYU0kprtnUiSP+wY9noijf2XsYxu61wXjb3WA3g0o+C4
8BQ8CczTkxifOb8EbXLxqFQsJqg5ykIXJzu99iqny/pxf/vnWtoUkSZKAefX25h9
dSLeEcfSnpaNDvnGg3n104Yh+9ge9k82FaPLO+bFCzxdzwwASFBBoUtBHJ2TYART
d2LBaEUguToyKCCBtdZsRyVnobypzYkXf7ZRLcoM+fJMjxEy7QpzD1K4EoxW6kdK
otvylY1YRHjQSYmgprF89xYSzFMP1IFfl7qoBsYCgjEAuQsA7qUMsxUe+jnnlhap
HKzaivjN0QvU5LeE3YPOmRKYu5cRCObnhuygelvh/03Yip0e6v08rnGJf5MdxtrS
BWK9RqTP4oPKzBzfBa9Dohl9hi3zSR0gvs+rQ9DsNuqBJdkHxLyCFqPd2pYLIzXp
5f+iug9oLKrkEwZxVDnQnWuetOvNmQwLQUGi3BiKzmOC6rJr1+UU0J09ryTrhoYx
tAX+VFo1Uh9aqc1vLhND5JTEjK39ZHPWcTKagILIOLCqXtGPhH95YnIQwzcnCa2a
4TQ9xYGMXuGjfPnVgEjwvHVASYihxpXa9KIXd5Dk6JvGRgaRvLc3uEcwFbgiZ3b6
H6SDXsxFNP/wPdx77VAUQfBDrIuieiNba2VaXNZ7PVzZrHxEFkbpcfYkZRjCt0nN
l2u6uL6mba1bWxVbKKw6OcW4+fr61N6boabNsuY1rtKTpqa4EWSiLUqK59mU1LzF
bli6zncgvDVnf6DEMXzeldl805Lf6e8AvlX9fCENuUeKByl7K00cX3MaJYnvg55M
AqD+GSgrG+n/edEDi+mJOPqD7InVK3AO900lAyVMMMCgpwU7U3enaL5bF6RcyGnO
kp2hIxe2InTw52BoD5VwkGJa3K0ypxsm4rZAMXqdRiuM2VGiokJZI8ryfX5OaB54
5PBgY2NOka6wEaZ/UYQog9yLD43Fa5mwHtwaIsMgzUqrrl9DEhHkp4tsNS4vZGhR
+NIzZbX+NY2p/eXfoMfyeCW9vEj2sU6wVhcvydM4GyWBFEQFvLK0wVZKNylgGV/R
bKSkPtt/BMvn9vpFzRxz26GOJQ3AS0azYfPg1hekJhvGUu7Jgd8L2Z8qCpOfviaM
hNcXgJfgdr2xudIH3RAkrzN6NfLjTLIsmk/3Ewi3FHqABSlKwXp0S0olc/4AWZ3i
UaSPo+2WQ9Aa4Re5XjuzABu90NR2KBZ7Ftw7Ldxk38I7v85wYbVTsGV2y4ATWWSH
38LcnD3qHmi2IpIcATL/QSmv88RD3F53gmTbxx2d11tB8rv87PDi6fsplNMbVF/r
tp8SvNn/2mFIQH2hPzUClvVVHKAVWeYl98DuE+cyS30oWKV60ptNpbXg/qe8/egE
eY63r3xoBBCl0/JQE8gwfl//iHA5tTIWIa2uU+FegDuAwTx9RHOdEUnKi1FJiUNm
djcQ0YKkbFNIbn7AivRvxiHynRdV75tbKjm+H59s5bYScdfJwfRoYa6v1CjZatjI
f3zNOiOFziQuCYf/zPzVOSkVAGUCmJ0+dtnmBP8VpciI+sFXzdXTgouHVO4cGRWz
oimHvnkTCNLjfWXV3BycdaZeYQIy1f20N6aNedH1eddSEaip4+DCjUMl+VYGmVYd
H1un/z7OEb4pp3r/1J2Qb3X4BHh4diVNljfIakTzFEAcYI3N7J/oHSjOMvv1LDVr
6KfGxcqjq+8wIjXkRp+67O7jjWpA4ZITgLnAea+a04hRNTt3WEWY7OCbRZB7UTd4
C0RlGkVFNc7lo8nPKuv8EM8iReNAgU+TyGkWVUtjvABaDVJJ7coc83Ixah3eTAra
oULs1bFnCAdugH5e828NwCl4Zx2YAMCEkBq2LrapPMaaf60jb1t1kzUDg6w0IhUT
HYpjHI1DqUZZ1JCf3tRUdvuXpt8cU9X2wUtIv2oBzQkmAVJo6Xlhm+xA42b6J57H
6VB82n/YzbYX+BXB9W0OtzHyrOgpIZ2AZBn5wFJ7ojI0rEK2SsbJuM6ApIKWNQQO
JgAxGsE54BeoK3q70elU1y1tVPx9iiD4nskMwrJFv0k7pGIzz0krmfwkOCssX7VX
pZYF6BC4OVqTKGyh4d+/F7khI60PKYhafZjWUs/MB8U1UQt71pXannr0hDMxNCL1
wXgEzdr3+3fWMqRc8Nu2KRdCnYArZPaTZCEkm9nR4BUBLF62ocde81mmMwlvaAiV
31cH6NCadZpKhjBixeIB1AGEjaADqWAwHej3oyh3hz6w3+2GFQigh9I0/3oYvZaL
mZvBSRpBfEJcnyv60WBLvkeJMpmN189OMqttbM/zfWi/mUbwXZ4bRUbpuQZ24c5T
Gnhob2n70DEff7Ot2Ej/Ea8+6OPxxunCR9JVdwT3PNMX8PPz8Jl/RvaHMoT96+pk
mPlF0hVAvNQPnxEFKxg51UOa4sBvogS8lRc+Vc9Eitcqxvc5M83Wj0a/vWQtNj+j
LBqiD8ZtnJM/aDJON6oiO9pGULLuNXZh3dOrh5xQ72V+0YpR8scVSefXp0q5qFa7
OWse7LBtTFY/1ZqulZqtAegPgsg/cdrPczA4x7Vmv1Y+uTERaNsr2IFedscpsXN6
RtdVU2Ye/7pylCnj8Fg9W86XrxIZJczyohq7nKtCq0HHjPpYljTL7JQ7Zc3gRHTZ
cVCRtYmwotDLk9U5ReafItpNyRAgai6C+FwR9wZAEPUtDkgv0v3wmjugkRpQ0IEe
+gDaQk9nEjLEVz4CS69pjWnDWdOxBiUal7CsloKmaNNT5TvMsmOSDE1X/oGYjuUF
QHFlAYGaXkOBmPDuGfk2UVnoQVHh5CXb/LRP7motjI8JOdmiVWWSR0SOHurnb+LC
M4p+VdvoJ08OhXyKVXXVP41eV2AljB8SxDErna85rd1q/VrlzlxE5SkgbiuW6SbD
YPLiyLbAbKR//K+wIlM8QLzoi/j3N1FaCmVqGu/9oTDLUpC4wVRI0GNKuG8QJRqd
H9O7RMwDt2XF1n4B8Oo18q5IwesYorpedfURtaPluGz9t//hbU9FmIk4pTAmYzAp
3MzKtY6po6oDRsO+GkNMvSAhN/3zBcW8Xe0rPiD7k6mpMe/Le2jP8Wjh4Hommb2H
4PB7CTfhyYVXTfD9WQAjek7MLQrhdMyk3Z9ZnQFFuS4e3T9jx705cSltUDUlxQQ5
NIF7MeFwgcB88oyKb/M5ps+eFGzBDAxdp8bsgu+NF1+jjYMnIBqUfbLH2V5h0oZR
XNof1HNdK2vz6VKeBOjS/Cz/AaTukbS1420t3iFZOXSsPHWqi4yBzEN8Lzam5Yru
oEVdCgWN/zE12LRI+6GdNwBXPimz6fA8ceZ3Xy6AlcTsx4i3lQO+DcxbNjJ5gXjp
lJ0B9Nlzk276IBt7MhifPC4LoMhK9Lkh3XTlywOf7letnKtdSVrsMQnMPvg2srb6
EEdqFUjMD1BylZn8wwTunFS88UPKWSZRwUjlhnT0UJzH+RE1HcLiS5xlXSg9U0qM
2iC6b5eBa3iW0fSlbiwkNZfJFBgGlcTdH8s0kB4VtrYCK3EqV+iyCAfWxMBtjI9r
f39qjVTrmM3XGYYRaEsxFAkM4PWy+ByVqd2asg7z9za1CeF1G/dVBEki9oPbd/cw
T6NNJFoKME/0LHGI9htEt3Zve5r54ZN6QuYBIggdOQy/BuwL2g6Zh1x4T+PpHgLj
zhG7ftcB+HjJu+5akKyY420kJyouAAvJ+4+3wIf8EQlm+Cs1YU/LUI3fEW6BPZOn
8AXrAROsp0selAm7ykBiruf1JS/V7nQjwciUI4CYhoZ7e+/JBrCKaLVPVoEQMkna
AEKlk0UKKH81z1BP7HSoi1gDwB1tZJuFbtkdw7mLXkFNSkPGL/VkSczkjijB17xM
HV8LbBx2qq9ovwpJiZ2U1WcYiPrwHWXqKHe0su2I6zVo4qid0vcOs/Wsxkkorlq7
MVMz9j0AMRc3BWVCc0HiMkfupbl4uSXZRlRdXT6s29y9yX7qR5TVYm7iJd6vCar3
J5cAGWHv9aH5Uz8DlDoQWqiPfBAfnFGwpTLNbHHHNOu4HjI0oPFiNe0ftT15G7z3
PGybX8jdSZpdYCKaFGtK+Aaxrhvs4jWlyZCe5ZSn4KUqBiJGiJu/6tzqshSbYbvY
fi53qMniY+6yLbZVsh6OiU8M6TfijzfMdBia7LsCCZwIZPZaPEXrcQ8LMRujMsV6
16oaDWri/dYiqKuGV9g4iZDyWtt9CYTjmRpIytorW9CF8W+k1B2zv8b2Yl8dOzDp
dwS7Tf8NJESNa/L2mh+bZ9v4ggu6iCM/hzgp49d3AIP8iM2B9ldZqL06Zf57lPh0
7Awl8x4WTfdFn33wVjQ2hwoQrSB3RPYqA091pXcqHrtS9E8sRuKuR7OiVVWJ08OH
bTMFBCVDbFX4EBSaZ2nnr8pOUmkZ8GYzN+jZVWrh1WmAfxwe2njaXYTgyg38EMiO
SMXYI54m6HF0HuBWqnGOXA==
`protect END_PROTECTED
