`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cSnUtimq4RSlOVoMxS3Q2G9EP7AdnHfsoYoq7P3dHau9+cTD9lVnOhlWNseT9zKD
oBz6R5gWyhyzeMhkLwPJVpc5WztMQGDXM/qz2zRbh99LL60ZiZxrpoZlYKJ5/aUx
rws+ajFEREK7qod8HSLQJuy17B5nVlUQZg7z+OjQjfDMlmrRiRHe6IHSkD3ovXJO
+WOZEdgrlfrssqLMFcwiQokQA+6r77ZG1A+o7IoGuLEO+f8jATTx3id2EsP5Cb5K
qdSjivF7hIWzWqxsiw9ooMSirmQ19i/1IB30VXiHf1YwM3oWyaU2B3GKdT7aF1v3
cPsT1LmaENJgCmsZ3RydSoWtYd5orgUqdIGNOcqF7RD01aPrKoHF7Q7glQd99YEF
FanDp8rEiJ4euw5zlrYO5PWiI+rEe4o3caUwRP3a92uoguB8JLtYRolAczTDU3EK
E26gRYLYp47Or8sfKA8wUeUpPp/Byqahp+mleRHlWQ5rx6zRcq2xBYYU+HWT7dvw
uDVXlnJUnxrrcGuLUCYaKNq+8DccMOoRrRniRXiu3ikCTnTamJsoHAPFZwL+7RKB
s+CNYBlZgsKXrZKHSBG2dgIOC6HL0rGqmQNozy61RfXeM3CVntSKLk5Xn+nA2xUJ
HiTXkNF5H2ez9h2elMXxdRuxg7J1v4o6xr1hIvI1tTked9tmK5ZFd8pZprNkS4ip
x8Wno+U+IDxjT08Wxt1iDKWYrEek1Yb0FdnW9U4M6N6if4hWhuxFSaUfeELslXUP
/A+aZwFT5wW+TpNP/+ftbNmEM5KZqJGx6rdUKSYhK6JX2D5N203LElPK+mTHbMVh
D+c9CsGCw70JZTDMboIZREL0ADCKA2BiZVK9zqvnY/TLlT5WhDedHFPY88SFaPw/
wkVK2PrdoaCfbMPoTGl3fIUzE99SJ1rMNfWWaP9NjQ/ZRgPPDwFrl2sPXExjmjwD
z20ilW/OL31xsb7Y5TmIEC+G2Nyox4Zc0llOAVUnnJ6E8ukuVK+neykgJEawVNIs
r4mp2q/bePp9BTnSJUbuYhrLG6ucFjTjpepLQADHRoGRNgqc7o+NswqJ6m+6ALIg
fIVA+p0/TLpPGcVhHDDfgNInnrmGWxy9/Bt53KGxMdXA1pa0tFSAYdLtlj8cuN8P
lOdKmcLgA7c9alyXg9VKoBLMz5mi+lfXYt4Xid+neKhiTgGPnMddqReHthAUYWla
ZFqBFid+slwnanWEcGu/Xpr0gbmkosy4JCBXdZGiLVzm4+OUjlgZTzZfvUHZfZFx
st8geJ0c8JObnVOTaDZJlzqfG1wHaVWOeS8kdLmMR/AqbSZQERURhuD8ZD23iw2S
A+h3qrnL7q3S5a46UBVa/losYWkbDU56FR9f6oE1RepQ9vg4w/VjQoW2qBV3kQwp
JLMZ1XJdY4G+p8SBPCgUAprcPK9gasUzJdQov7COU1M8WGxcAJbBfB1z8G4yWPXW
fDJxZpLJKu2Waf/+99J8Cfo1kbbWcfCviUJceIt78ia+UZprl/GnKnzCImMyM5ui
Y+Sm8wya8zoH9O8c+zglzzSZ6pqbR4lwIPDlf86sFC818duSy8XuUevhCyAVzcCD
Jz0CS9lHdgrTw7fMRmqCMbyFFuHGPXYCT8xSrsEOfJ+xUewJScohJw7e6FNYMHrb
141JB9L1SdMJqbfQaIEFVwBgnB6jpoplNRXT8f+hAbw+F8b0IIv9QNcWlZvT8efu
Q2ZqC0XlcR7wuf8AaQuujx2P5OZA6WiTxstGMb/VMOuQerY+dm1SIWbZt7pku3w1
Lv/jSWsSRO3/sPk322mQCPL9rV4m5d6vjxi6UToV3XdXG2n6CFH0YdHBfhSS0bcK
Eatp/3ejR+BotOERXCZkAQtgseq9kK/B/4y2xdZSQo7Rcwa33J6HvoWEbZU3q+Xi
94gFlNTjb53wiy9eU2cz/MyCW+KnO8zk1JMVoya3n4EPlPMRTHwqDvS/ks3pRXlu
AMKGSCuYA6Q9CS9BvB2bixpZaJm1WUh9c6Vv61OQNocyi15joo1Z8GtGuQocU31e
VrZy7NKplP3CFb2KOuKGgJFLxjHxZ2Pv0Ncw3p+qyycdM3+IBgr/AYObPik/304K
17dHz7dcjwYgby1PqBpilNxEXcdlgNz3HYwU0k/iZRc9Au9zUAP7fbj0SGiOzcXJ
93dDGHyA9a4wgpR0wBcW9lvn8X1C2GZE9n3FBHJr3VLloynX+rTaYcZN+jZa86ar
MOo/q9Dr1SXenid2o0XPf30dGDANI9yXRSteSsAEtYrru4J4zMqUTOWvOLkDqpa0
nJScQZTa3v+I/4u7jlBDd64umFwr6k17GOg04gq+Kv0Ofbbh4YDHhO19MF3sFD8w
OmcsD0SEytfk0LJk8cTaj/xd/VARy8e4S6YvelOvKYOnOAnrS+unFZNmT99x2i8r
UAu6qFtZiD8RrujLtGn4ae/0TflkkJeM3Rs1AJWU3Wxb4mRBN9tjpHesmHP+3hGT
9NheHOZ+Ej0fywqi3mJaTQaIti54ma0eSG6mtyJ9IvtVS+jqNb/O+i95eWdiw2OM
q3dYOEgi+O5HK0sRkt4q/AcqHfVLMvl1oYZ7E2FyFCwfocOlSqodaJcWH0W2MbMp
jIvCj3hCTf8dqq2G4vgRiLil1++oKaYn5xqyLVXVhvNjvq567S4VJmglnFCy+USN
2HqIXYspZnGz4DP4GncGgHxvSv+3bAX93ktjt/fvFYz+L/UbvR+efh/U/LH7X4ix
5Cd/n5CXJoXsErojsu2aBLIQ2ZX+BwYP0TnCf67EW5Ll0+aJAbvX2zbjESy4y/D1
LOw0wuG3cVWcuCo38cvcqj4Ve3zbLI0u65Uctl9himkhMJfKh/Ji7qQvx9EXLEh0
FI2FMRYWaYukU82BCE8bbyxaqtKeMGZQcvW+Jb18x47epAULefRZHQg/93V9nNqN
hynDBISX9859mll4MsK4ZipLeSGOBWMzdnWpbSCsnPuZlNvhEpap3lgxztvEw9wG
Op5ab1Z68MW60dJ50bk+Yrl4P9p/z0eqPazltJ+YuBOHHnYs9c3kADiBTQUkkmTr
MhsFFEYwQWl5qwEhVufwKcQd/Q6ezMUfL90vKCQgx1gSFmBYrfLNqdg1Olm6cnF2
UTdO4Dba151CxH73L5ZHQAXQ8Kzxpagw04qlyn82uM31fXWySkT2Mbugb4mL73pw
ecHrzt9cflgUlb+MbCqDGhVBjMlIsuHxDm0Xb5dVLah2BV46VWD1fz87BbP+R0xM
6GiehemKmSrdqOTasKd8YpJBtB7sPHKY/0MmtBkRSK1i5ouO6e6NiaG8ktEGGT3l
gp7HvUF+M/iIgNY6TteKJF/LUdZeELoUcSMw8QEovAtqs8xYWhmbOf/6VwSGD0er
X6GIdrBVpI2x/VYSZvQ7DH5ys6MFtQl+DP4sBimcJzak3O+U2d4f507rWLUgiF4L
BPxXWiosKat17WQLRQ3u7ztR9qh0qvvQqiSX3D9+bk0wFPzeSsiJAmER38vW6mh5
fMuZrTi0eSCgkuJDpL1fSKc5VQRtZsovG4Ra3ZiodAC7SgQQ7s/3idQnHn62MAPU
gXViacpgz7NsI01uO+xtOBXYFoUu4NxDMVa/S0WmPnQI6ciI8nkYypQCXynEpcUH
2U+NAABq6pnK1tk3t73aPCb67nof0I4hdjOtwG4FwDQMPIfDBxjrSZqHy5A8YJK3
vSLAYunJGsDfuOkr2XIql9KCo8gYL7+ksiXGj+sS1UwYU5vm6yZc35XMJo62Y3Ky
2CAvQUOuCLAgrxHmLYrcoFRhQIqrCl/OFM9CDHwnMm5IdYaLlFOMWRxfu9wEIDGg
x5WMdjuWRCYiI4m0DcuGWaqz9PoPyJXHEurS8j+bQJail0wIXL/93ErVETSIRlSE
m6K/fRuVfAK40cssBTAKU5SIAZ0ihum4gmBf1hxfiYIA/QVEAKPsxy8GpC+TO1Gb
bXX78Ny6YC4uYY7nkqRvoxNqDDzIrXfjR/jUeInKqxvr/heyXu+tVeU3ZIU/Pxla
jFg4kX0pF1Mal9bklXgvGrFBFltKGKr9LvHc4/K68N2ZR/KXbUoQyLz401TMavcf
Xpw6La3MLTYOQM9oE4n8DcPZMDBbsXXNHY9DSL6DPbTqipAgPwUGltpQjCObCJ05
C0iDUzjjaP8Zh0agXH5o8pVeVod9E75BZCwxle5el73WK1srPt/qCqm5tpKo8MW0
GGzrMrax3tLfNkLfR1JdRbvnX5Fyu7xnlCzc9EWAgMvePmL2Bu584BMbHB/xPrvI
K3b8yUEvDRjIta06zxQ/4vKz9WMox4JODpUm386C33tI1yNRYEs8yLLr4T9xFQx0
c0jr91R2lC+cEP31vUe7cWsGiRKerrsN7SbYzka8vXh/Se8H1jabTiOMIMXeFcXe
4/DtV7yJSrmH+rTPN1XCmlzA/5wcPk65+bc0paMFzqh9T1ZbMIaalZggTS6DDess
tCGP1LY0T+HykDh3d96f9CgKY5wMRgF0Rz/x6Cyv9Qm/M+q1wH3ahLiiDdqxtYX8
baoYqVeEsQg4t7GQ1/ycZS0Ez+zjQDg1wQklGO/cyXXR9BbY7sUd3hKL6XA3m8+I
P8bArM3Lzpa9tQa9fxhUdMAcxAR14xqR5+erWGHbz+W5OEYNWILXxxns1hmaxIBh
DP2OnfbypDuTl4sYc2EUzGELq2qq9iUq5aNPwGivdfonXgRhjbl+y+e5GQxSzjRS
yvfbKTq/k8lv0DfyBljcNpW37fmxrhsh9UdvF9b/lDg0sV/6BubEhgXiBXovr89y
9JeSEAi1kMSg6XikOLoxeivndhXfQs6/Rw8UyLwHmCDvL+wjpNiER+K3OpxloCUH
iNEoJcOkKZmstJj5+gIYLRv6+D5iL3QU+6jhVQXOav+R4hm+UOhM4186ojTaWOtj
84zA0ATXwQJRCBaeC3LRD/otoNHFVjhcw3pYf+TYHgXpPp+l1FtGnhbN3NxCO9gK
3Wfsz7gZh84AQPlmpZ6kfmcscUF5T34KURasEpnXx1fJ/Lj73n2fW01uSUGuc3u4
ey7Ap3EFqA7Ho2vrkaEmwzj3Mj7cUn9yF2Fn5uQiXn5boefMBJ4r3JuLPUaW9CuK
8xiHQRhqgaxenhHR522EjygfHkvVrrRP/4Zdv8Rqe9IIl+Qe2TdRax3LMGwgP/6a
HCrVGb8TpAHsKkQx7HXcIItI5mWoac3teFUHoSZib62U/PG46N1SUaaVfvhyPFrA
tRRG0IyrUFtXWz4Q6KDXZ/yoUYdmSTuTr+viiBi4y0ZaIy3/X7O7QtcQaM7RU4rm
+DHjNsbgovrG01Zc2WEwFTGGP6mLPiQn2jlZejBL6ghaBDT18q93w4MvxOpTBnLw
p511Pawu871BW/0uGAhcavBgqc1y8gQus4jwGxg+9ev/akh2bb9nPkvUqUoIv/Fq
uZeaSqcyGlO5pTOq/hvTdAEUArNQzzyrQnTH16a026k7pQY76RktluTRw5A0btEm
FpXGx9GmT+/QzrMGwh5Li4PdNSM2zPf+YTYzW6gIr4nZXBIKB2D1KqleReLyJjAP
WY/7aPD2tLCm/Px6u3r1VmZsTAuTM1iY9E8FdunKJJAHvqG12kRm+GDrSpGYprQI
hmtXQyKbjJdx0sMBk/ucPIq22wYbG35gZ1NnEfzW5aOssJ2Y6dZz2H79n13I1zez
ulOSu4Mhy/6nusrYWSxa+AlHna8VsqJcV9JY3Y6f+L0IP3Q1IVtdzQ0jzM2+mnH6
NElJ9nZh9ppqPqTBQugMNVBlevqzwQaWLtH1LtOgPPFwjs/xYL1YDdvOwN6DEo3e
K1WwSMtuybbNrs6t8ihIRFpVzd6j3DBDQtcZ4YcEZOkcJ08L0qqIsLkutTUQDIFl
5ozdJDc8yOPtBWniIMWSEOx6Z9ORxv+PI7L2R6538+uKkHVrxWfTL+zfPAkVvAbQ
Ogh66AeSlu0546gU+HYHD+TPzKxBYo5xAVX5NQVzEfW4oJIYPmB5l1/X9Hd1bc9f
KlL13ax/mqmMxnA2/kAeOFQw0ODU/oGMY3ZEyAheFRkrlrrXWAFv1KDLS24F09jJ
ppFIy+xJKcLmBPeSu+EQlHCBPln7xgsrncyFiWtgmRYahm0DkJo0l7Zt/J6yaM6C
84/qrkYp9DPFj8GkvKPNc93W2DgB0YleJMYbo4BDrN1mVHZy/++qn31jM/sMJvSv
wYHkc5pVD8B3i0tvBlvYCwQuuDH0hA9GxEx0X4dLCxxXNX/geA+JdwxJz4uWEYu+
cawNJ9hXD3233R3+HAWMNUVeigpUyUKtu1nHqChlNp/mBhEGIr5fgN9fTXVDVK3h
Ktr/WKBVuh+CTzHJlkEph0/hMsPECx4MRReTA81oHoWlRtSXh9bdEKHPIS4gavid
QOeKzmCEPFdyI+Dq2Iq90BELVBN0fhXmp96bbZbDaxvBwdtzGkDR/+mKpN8jcPfL
sGReIsxSnHB0OZZWUQuph1D+jBVuqTnR08xpBT+73SHijDsIeXcQLukP1Jbb4UYd
VTHScN5P/a8aZ//iXgVCBtySSC5OYxQ9xGqnGRfblrXVSO32jVTTueF99hO/nyTT
QdSDhPmYZDYZdH1JHvgt8syAHrxMlTBbwME/ivGE5quOW66lbB6tjf9+6Ir/q4vO
qTeAXp/wHF8xLUF9+c3Mehce+aa+gEJyEcwTWGwhCB3SXRUL8tda2oHALRXXaJ+u
eNyrMlslAi9Z2dTkdkGm4M7IvOirO2Iw1x9umY+34nZwNmFbrGjfz10sjkN/+llx
TnJYA2BHe+RY9gQDcQIIY77Vb7rqZBufa97lO6IgCkb88FwXawyjYC4V4BuCSLLP
FvR/jcbsyc0LPqsTR8yPjDjf/uEnc1algv9WBMX/9mxLQ14VdhA/SHPQ0X2WSNc4
TzWlD7h31QAG9lMrM8IR9safbP9+1SQjG2hR7OfqdWHb9scdw191ZAJMGnzTR03n
F325Tw0hTl3rzOvy9HI8Z29i98Wg5x813ffKgB2d6rq4YxZ44JWbbwYNZt98oTlX
L8SGzN+XPsU7CcojNQU6Aiw1huVjWTWssr7DIXPGxZqJgPdOlb50lEgRVFoTOLHl
Dy6UYN1niw+KCSNUYNaXQfcIXeGu061uPuuFWLW7rpJLUXrtttWERiIJlnsemPEe
OFbIbp0mmHeFdWMDJYSyhfH/Iu3ErH80+uFSgtP+l7T4NvvfFlop5v+TvP+zSokG
xoYEKywsvJba8R+kzLsZMS/owV17lb8Cpq2E7Z7q6ziIVgLWI6FDRvWVWnESMjPo
Ms67G9Hj3awVn+RXzIBT0Azwvvkmn14du/8j2/M6nqnv+iyHyi7ft2kdlzDtqNMn
WZ2GdpT2p4JEqQ1w0Mg6Fig/T5+nozbbCV9rX5D0bmtYo86w5oYLT85XRltotNzx
9dsLjsK4ljnyvS6prNnhV9Mxdv7sSZQcG43WMXmdV8IET/O0BrT1O0rcyicvHCaS
6jLi7637xVOKrV5s8ZeleJ51J+fFx2mHXy+jhlbUgvBeoACHKgNWCNxnXphkbHPS
Qi8TGD4QZ9t6V1t/FcxABGGxKNMRAmKKsqL7BrvGOFV/vlDt2xoKNPECSWB5Zmv+
94IL/7NrvlVU09q5Y4DCiy4Quqvu/p8gT5LYNOABCUalc5Qjknt4SfiI4yyUlJqT
baWn8KxACxq4HEcmo+q3KoOup+dKtq8MHfb0ONzlbZXflLOac60Q+0zSngmnhgKV
VndAcSGJV2PTEygNlRGGXwkiZg4dz9Mu1WFhSa9JcQVlmGVDl1PNeKc8qjx0zFEr
sscHG5FHkIRoHsTloS9LEn6TDmo4/S0IzBss0IKieHezSBkvOHYF3GOSC7tkvI+K
DB9+vZjloqIK0rI2gZbog2FDdGLPhu0FEo8GOw/romR2cUJVWnLR0gg1srDtbZoL
7pDDR2HO68JAPCQagsu/LIapgEUz+CFOCLHhNhSNg9J5cN1jVDT5EjhWC6lueQXb
DtOecqopPT8mhXplu7MtWMrAyJnvYFnWhkAQjMYcv3SABPyPSFvHMs4CrxYHnVOr
nL9JA0ehLqZ0jgOw1EL3s6wuwFsbBy1N4SuT9+GpHyGVUgHphf7txa5jDK+wLx1D
m34d7sGV1eHP5GEr9PCPNgcAr7VIhO3+WckCyRI0+ExzdIMF6wPX37uH8cLX/xDz
dfvmQzgE0ffjD8EwWX3ZHRmOys0dOShoe2Dzl0VKL4OIYhzT/LcoXcn2+qBvacSb
sMujyIMU2y4w2z7Ye4U9WqNeNcC8mj5QT1Klhnz1ln+qqLsQZ5MGqbEtc8t801CT
EbMe0EHAzGILCo634hKrHZzpkhcHbPq1jV1tNgSsqi7tZqeSPFIkujDCN5p8kH8N
1D2KgPq0OrIcGBHuhKf7+OC8hZHfRryY/oi/Z4S9kcJ8uMj88cAmgH0LByy+Y3jj
2MDrT+17cW9Zp4uJby+di3vy2UdnDERDRLs2zE0dQw3ReQh59BLJwgTjrDQ5uTE8
Jy1jRXfNyizKIZb6G+BjCH+Duu/6kLw3O//CIb5AC1j74EzbnSwYGSMi1oKIKMbi
6fjvB3zw+bOEAUKX6L14RJP7ll38XaK6yv2qx1mZDjYOrk2E8nPgAjR7M6QMLRo7
8LwxNXejfGfvM38dsMMKLcZ6+q7rMcQ9l2w4wz5tEcLcFAx3BbQtOrEtHJnFL10f
pz9Es0LHWsN0y8YuRQYnPoCz9uu9UiceVzHUoVosHDL8XFgi4275LVZiKw5Q5BYg
CBDfGdzPcqWXWDczNfDLu+EBb85QzgD0EBYrDHb8xp7AOJ9n763v8eFO5UGnRwHK
F2+gkIYeJsmOLoKSvDBLkPxN3roIysBpGPEoPGLqFXSIs5K44+240K1ThfZiST8y
e2F+uv2esjFCC1rjs2lVvPFdqXp7DGsl71EUH/eaiuUF8xCWbCWFviecRU624wcD
D0N+wQdenxNwh+SnXCYos+JGc4qV01SSsFu9WeBg9SSX/prbb3gcrtm0uCT2YW+A
IjW4hdvo6Ldd/6A3AWfGDlksqwnS2nfhcTxBmWUEmmMiZ/x+6k77kKEmoKxf8jMe
FMsQyJV39moktEq5lsFjSf6HDsjCMdQJD4hGMVo1ufozY8+eu9LC4bzpCvYbhwuN
UFWg2ae+FWVitXcG8sMfCKZgNvyuJdU3bUGn/EPWYQ3g/rGQ+J3JCY4VK6K2SvSY
G3G/pHJK7Of+mNQMVuX55Oxm2vexLf3zgySbK0HyHMl5WwtzRku8tvr1q0Ownyt/
CIdIuEn0E5L62lFHiCH/IesRN2UB6L49yy9l6bHawjsoLWA19WfDIyMY8GnwNh/5
OlnfITwi/wAq8N37oUziuURQ5KTGKYvnGstTHXvwjVfqyyFMznyjP0S2LiI95d4H
1D6+Iiw3g1V8CWsyXLHMLzm7tTtQm+m0dqgqKFpA2dxeQKcRLT5AvFKlbhzhatNR
7JXuHlHKUtzJd2spdUkIgkEDpG0Z/8tWpdVV8KW43fQCtmPKZAMWrgfHaOwitbuA
VFKu9WU6xxbVn/5NY4DJNFHfzQ7AO+gMimFDG6BQGAs/t2VqyKXhw+nhBzZo4OHb
yYsYNRv1ZoX7GJBcR2USv8puGVbCf6BJbZxP8z+obgDpilVAPrSeW4beLXnOmJCR
JDzHFICUqzNmPCMiw288NQ/RuFUxX1qJHgK6TIoFRqX7PCVy9kIommCurUJAwg5Q
B7zRieeR/UVT1TLrr6wCgCJRrByCkQjv+FyCzFCeJT3Wy3nKVvZR3+9M9vZzkcC1
th+0qrh9x2P4JipiLxNyYEHIEtKCSXwKMoN5X6s61/0tL6bszKHIUqiEnwigiXOe
oyzXXyD4xI8lb/2xnK/7m9iHZl0lrQf8C2DTsxod06I2yEn+T+idCIRf4pk85SfN
6lVSmy7ti9/48puN0X9Fjdgml8PCjHlxT/olEJY9+2q3iIvLMX/tfrXKUXYXqoKu
1ydV+/U2yNEOablzhFNrLTEhCRh01qZyp7szdYMOQCYdRsRY8cp1bSJpjn1Z2772
ZWYJTGhw4Vz6rgaJwiiBFT4Qc3Z7ZPw7TWIbEEw9P+X7G8zWn+55gZlilAVzP3b0
wFPewWX0thC2rWzuvBGfdMR8snKzgOG6EfQZrkmbydE0x0zz6jL62+7lBRR6bmZo
boAY7Tr1LmO32yerzunP3X9RJCDxDX0jF48W1NfUo7ypPFsc0qFVToojxjp7Fuoo
XzZSNzGAufD1bUDa3iXXxAqGErqP0rDxhTPMHWf7ht/MPYgQo+QIQS34k2GoSo9j
caaRVk9cba8G3G8u5+scDGDXnl61OvAMDx9X9Htygd13i7yfKUBF7Gd4PgCWroQd
2AAeZRldxchIT6KFZ/qrINzy5UyPNAJ/OYLDtUQIQho5MJviS4HGFo5KZj31Hc8t
83w26qJ90DWzmt4kGvy6skl/+M6c+QuoivHIsY1myqY/Qlyli9YcLLKhoKGun4/B
TUjIbZ0HI3wMtAvF3pYdFgN39feCs0FgbS6pzhGwq23/Ae2pfBKYUdlP9CM3/ykL
lDFvOVqZPwOLZnVqKGpoRFabyBok1QHWvCM3DDU0LNcPKONfi6hiKzcdsHV0bPI+
UjNedrgpKpH6OKLwq9E53MYVvpXXFNxHpUS9GNK6S2OBMXFFqVc+5sp26Lw4x7Sn
31qoUQwtKR5Xm2KQmFPLFugFyKf/83dsBgBziSqyIT2/NIkZAqEzhbdXeHaCKbay
Y27yy2ZzG9Hx19tJeptHDxpM8XS1s+y4z5fRNGnhVjxun8DrlTpGKiFXwDmOqVxB
ScI4RwBVSgyz9FleV6fsWyXmJY0BxveVDzIkc2SV/Q8OTEv/ZxtIoDRXx82LKQ5I
q+jXbHqOlEx2xsJZxs9+Uw9WIb+CpGRczWr+PMyVqZGuNAE62eNDOFLZ1uFrpG+P
3tlUoxwjQgcHk8heNeJ81grdmvCgL6EuMQApnzYlhh1ONR4T5c/g3CPIVidNSWE8
4OZp07mglZdqeOgHBfaY+P1lty/YEX6pwZlgRc2I5J7zKrN+gmNu2f0YLhd/qOR7
xKyPosxhAX8gBq0cFTm4HPfahDzbbeL0Au97LBQSQAClc2XboxWXQaZB3Y66cfjQ
SJ1hAF56dyNx0oJuWtmva+x2E8e1vEROymZg4rrZsCLV+pyNyR2cF3fQ2Rl2U0tp
ZuV/UFhFAi1ZYS9IBIBnJGDSrezflVV9Q4c7RurU4/7M+a1Kymbnz1AuHqAa8Nwb
btE3Lg18OtXD4AgcnxybykU9bg1rEzEYE6qWR6AVYMpMgklyfd3fCowH7E0aa5vO
HXJXrHn3jRTreZZ/E/EWar0wRRGxALTQ3BrULbFo+k3T9q0KzRpqFL6jIJJ7ZZtX
PTAwSTi4YL1+adehoCcM51fT0x0Nc1dm4n+Y9xuLMFzML6BB37+CdJWS9g/K/FeO
xQpdquCRzOdGYfz6RK9UgRQ1x696gTuIlZlYeJGEu5MJ/zfZxhHg+8Z4SJp8oEnR
B/qpZkBm9GAik9YnwtyhjNulSlZVy+VQ/F3/HetR4dkSPVRvzzTclsD+JzNyouZa
YmJmKAFfIV4xQhQxuinyeF4rmay8/NyEVWEL1ue9I0a7P8XJ9j6GeMupe0ZRpL6M
ve0Xg98XUGqUEQSSXdTIPBvzmCxJ9moIDaDzeTyL6pUVwlJ207hy6TFB+9RrL29Y
DpnXazStHQBPovA8MPYgK4dbKbOc/Twr4ziuCLI175qEuRWfLayDAGfi/Qxk87iE
bAV/jgG8ZeDCaGoq2Mu2pKjN59e2rwWV8vkvNwLqsGo4+yC1KJqAStbd0e8a9OyV
8YKvvW6/W7klC6t1pnND5eHhLd05pBzad4wJM3+3Ke/03VggiyWFpIgOnPTzS1RP
eMn2f0sxmsdSRtRchuPLkmR2YVl3jxwMNkYqw4B7jHrhXZd1RPwsu8U9izYFFFWc
EZRB9rXNqZGvvyYL84CXnd4jDXybSduDGZiDWNylQkb2AxTxvjWjR7aEAN7nw5za
pdsdXknCrMC8S3oUY7Z36B+XUvbXuJ2wuQ52E42ooiCaWY6tDjEU9toODTcRK8qZ
1zrHz9NeoiPNAFsA4/bx51bailhwIac0xkDK9s6rwwCL93XLv2OLOBQ+UmjWceyv
t7SXd8pOrajECgNyAO3ZyXNxSBGelWWITAyus2XZoUBHv7C/AJLRvzr8OnEp4PsG
BEDsLw0Bgjwo34MziJfBiuAFzpiJc4LUsxeU3jAYW+fH0vOWBdeeAeN0qwIWN3mU
pjJpucN2GrOcyIQkO5VdE/HstfIsg2eAbsDTGGgJ5HkWxYE1zasNTxyWjYlQpSjl
6gB642sGGu3LUBDloqsHlHVdSk8RkQSrmaOAwlsSN3CFO+pDzCWbBqOaeDuqMZsK
Sa2ePJVg9rIUSL2sHIJsM3qG6LZrZx+/qH9pLHuz2uPcfKApM/13XbC3T+WEHUan
1RpnkmJCDkqNHUVhVfUY3zzq3kyI+STPeDV9l/Oh3OTGZJMZ4y9Ua6E0lIjCEG1s
RSoadsAU/jSaIZnFhTKY7RwCjdQ8oMwVe27M9I4NXmSozp3jXx8FBSzkjjI48f+0
SEyYxZ58/TRpRyQe8kNvfUYyOcJx0IBdwR+nHSE+ZhPXWyvLMyJN+uIPdEal9LUv
+YslJT6hA/9ozhkJD36TfZcNkB3iPZJEzv4O6TGvFDLKRJLiyOiM5FaZKCR5bxMU
RvaEErVs/DGrF6Qng2/rpX6Xde1QLfuivIshQWartEvUfbwdxVdQboCkl6Hv3bxx
xO3khmREBa7d4TemJW+kY1a+h/gxDFauDe+0F4wBTRdNbB+sAJn8H6foLxYi4p9L
ZH+zZ9uWEVYAtMqqG98/Paob2isF9gV/Ei12s7gEWXKRehclmiPxyWXSMMtaT4Ac
7vT9vipbgVvGE1ATVj1yreeVmgKiSlqQOX1xd3i1OeT9njZsvoj/g8SyWMs2VfUg
i8L6MThM4Lb7ePPpqJaBRo3Y7kR/qWXnClzYgMkfp1IkFaGCWrLebiUY/l/YdGHz
79A2nBhr2SeNCrP+JxnNuVEJBIyrnSAksmhSEJi/NCi+CtzWwy+3oM9CZ22xCo5+
4W9y4REU/J+s1A+F/YsN4BU7ckQMkM7hdMlHHS+ahRr3Btz4qFgL1Cs+BeAOEqq+
///4u1N4VhfGpI6RHQ68tMzu2UohQWTFJgmiMc7HlgR7VmfhHSm+p0vNRkkVQcLl
t9LhdBSLOLbOvq4PXdQEvbdR32+mOaAR3GVuJEX/GxE5s4WzE3N3u4pdf/zf5Qnm
KwOdewsOGZBmpy6Gs+hc95cKt6O6btree4HOX9BQt5lPa4wTFL1cgPfidsTOCT2d
g/R4UU9b1O83xw9Fg4FvrGOxD6SdO/8c4tijABFv3c+nemjXfXg8zLRDsyec8IMi
jlp49HllWpgtmUlTP3cHeoKK9Go7nNOnjHCaVLIUBKnmv3wiZpfUD09ed0lP4Yze
Q7FcXdvRgTGcdiUAoDpXc94aKrLMzJ3pIqt14nmrXjbajD5JFiO+s0Gmp0HK06Zu
rHW6nvUj+ljEx+ykNODSrU4hT9lHxE35+Jsqw4Os74m2Vlk3qganWneUNAk+3pfc
CdG/Go94/rlGnSO+pILktfcMrEBuuyI5UcTV4rKgBA0P9xbcGbHV53YOnpTb/7pq
TDvS0pGLGaFKyuLfaK5fsHVvrlAUB5Hwrka8pK8yV3S2lw+OJdq9PVNHJatFDe7U
xI1/OAzbl3OZqaw8ho0FLykWy7hhsmFiNRAtMiVg0L2YhLrRuT4BwazdBBLF+2Dv
xJFMcMMhU8OzNK6UkC1+WBsItyanaIQRUA/uNqTrwwJGOweK9jr5pTzBmIYavOqm
OH7Mdbs8peIrt4s5KLO4ULxzuxNzcSFXDL5CupJWsWKjBwHROPxUtgj+Gz+uCVpQ
gSd8MoNmftwUPv1zDVWoWgUiAuFgSYbbbe9cR5tRfy3X/fNn0A/g+TGE5hHf3Bjw
3OaNrPuRYxLhDmTZkhA6h9+Vyt45SAZEus49XqK0UOOxhMfxoV7qN06EHyaYP9Rk
Pif5HBO6m8c48rQA3oCy05mfStV1tHYtmz5DUvrJueJDMGx8iAZM2Ndo+b0Kcg7+
gUIf6PF0KJfSGg4M/VrG8xlH35wTSR/9M5w4kXaz0i2PhKfIpQ37P3VYwvDapb+r
kvZQ7U9L4CAVCezKWlI4HKJLDJ8V7PV97uc158enjpUGjRtA8TBZtV7zXbNuudRR
uIsl/a6F81FzqbY29+QV0WlHW+HL2SpEgA67UZnjZ6IoElHRsgMUXDlcwleSzAQF
j7yXbOaRBT+CziNhCp5kcucvUU+jOoNbLAsEyHtReovEkTpm2rNjwG0GfMOF2uYy
BhzlQs5SRMwacEFAMFuaxunr3XGljjthesMhB3tPGzM4oOiGAjAyH6iTeSxHnWXb
rmhgOeQb+jpfpT7ruTYSARWv8mLrMDqcnoxfgB2psbst3I0/dn13SoU8Bw4pUE/d
akBYxsVQ3cVgt69n1yiY17a4nYJnLhgFUiyMnc8P7b7ScCVPalPnTI9liu0nIUgB
07HwREIAVsLQFqfPru7sBIXJHUzfwwWX6UiZN7zfRcbbAP8ECUGOXiByXjDTh68z
L5A5ntZKLR4HCOd5AWtc6FJ7XGIlltkhWgsACiZN1jgGoA2qcuJAaxCE76TjKlVY
NbkXjvokFAYye2svSYRF0b9J1C+fFU4fgmE8Cyw5uZKfv/PpwJtT7C3whUVdML+e
+EYbr2HbynMcssO4NCQiiYIjBNXGV1xk7l6a3rOmk5Si7/6TcA7htzzHxd8Yqa8G
DfgNZhQ1dBW7BH89L9O4S5H0k6RIXui79rFK4EJ+64rnZxXM4LB3iqVJFMDl0gUx
oI+0kEyKpxKWqNW1+MNsdzxbgDiIIB5f2ZVuUm8ipq1W8rEpWpJgBSyrMtGNJzzx
bmdA2meae8KXYcpN7OQUF1A7Ozj2lCqn0O4D/jFB8Pxm++q5gNLcYSQ0MkpBxADE
9sxhETKNTZPv66oLeMXx7VcCcIMhT2/aep43K+OWS4dFNBzKIf/I9EqiZRBp9Ft9
Ld53razUH0JHd5sdUOIo2wOD/sUBiscqrU1AYdprVTUg7Tnq+WxGvQVIP1ozuhis
WJfUpSDW57A6ZZ/LSGYDJa0LyUtWZYc+OsZ/Dt84fDY20dqmL2T87Fgw2YNwkuu/
w7XD9NuLvnRibSXA9YbDW9PrRi0hzAWrb1x/QjSOLe6vHZS2vbFA2e49VFdpj+4d
8+0nwVlHwgALk6ofQF3phUO8qyzIjJyFueewGEmTOlVaxPIihlTlmGo4Q6Tey/IZ
dBLOVOZse4RjmMWcR9sawcNy7zOiRRFeUzo6RFRUi+FcsrtKk0mM6i+23FdQFshl
YJqr4/sq7QEECuXiCTP5iVsNVJJNDbPXK5VGRLyZbfK83OsZrTplGOOlYobP8Wfl
nsq3kaR70bKo7QKuxNcfrp9lvu+I1Ckuf0yruw9e90jL3QGqhWl9hNJwwd9Z5WUX
/5fmQTrOrbs4zogUNdFBcHoyUhQ0WaVZTdmXQnAZYR5rI6n/LQkRa12L9mtnH4b5
HL2gIRtOCt1uhUwLWymCgkSvzU/6gVSnooGHr7r4Exo1H6D2FHrxKIiiwaCcAYI0
i4PRjtVa4l2cA6Ba8EXQTCuG6GWZ75cyLwan/5VXu7J+fHIXqVJfN7Uw0seWG372
r6JMDgeoiCGAUyvRgx5dqU9NqdQwn/GAEYeDvS58K9u1fFdu0BoI0N2nJtCSs8sX
X1+gv3ptlluiGzhHfQmeF1tQJEw+awD6ppYBxrPYg1AS32RtDn+NtJVwi23l2vfU
5ScBLkUojbkG6Q9PN4IuYPeytyNz/0exTaovtMwhvd7pDyUlO8SjFhJ7BS43WUS4
V2SBvK1Gilqlf+uhHo+oAih50Td98cTmddRoG8QOQ4bfXSyWIpNVCxNqR6OQeOFw
5s6uETcuGMlM4fLo+y523+Fgm93i2EDwf+h6Fn5/+5NSKeYK/+3ZdKXm1Cve6FrV
lhTEotwlx4wCpWUPFVkfSGYwD4K4GOE/ifkP3Fn2hOaQa6dSwsRgAl1zgMl8/oLz
7gpzuqfFmcuPO7EzRdSIRm5+lbPmkGOqtQe1oF0XuMLnKHRjQwNtI5ZgeVtQnk4k
JYGDxT+lXPIu4/0XTL93u9OqQ17ufsbc5MpPFj3aziMrq6KdY9qa6QWPv/px6FwM
+Ezj35ZNEBKbhAk5cmcMRCAp6LPyoKmHp4mD+QVMcbV9+ouI/OWJAWc68TsddsJe
RLa/a22ZVcfiFeINBXvk0+edTOxY8kNKDpJzDmHtXUA54nSGe1LQOsFB5rBeuxdd
rS8/DxdMB54ucaK63nhFjwUGxmGaJ+T1rN1/1/iNcsDwgzHa9iG48Py+6ms7JnCR
a3ZHDCSDEt1SVFhl/4wePi/gsiaQRzJ3/7Dfb3+DOaGsUaY9Q+JVG8xMMZWgbVLB
32KMWJJeOA4LuyAcoaQigw4X/BhYsChdaOklILzw+jJmvVAMSjUgHD3raSwmH22C
e1GaSF1Y/fxAZYsCdkvPzGVQSvCx7in1AFXO2GTrKsYMdpRT47IUPFYAKMCVL4/E
6bKJ5nNclRKbTmCH7kSDeYDYe68t6p7xpIjeCYLG1WklLREXJMXM7CeAWzP/dUxN
ZA02OcL1KjmWXBvw8EcsySpN+oWaRWRmUUSbJRu2D2ZoG0FWRZFjpYkfFDuCP/Rn
SQVNv8ocBB+daKhLfbi+xOeod7d9ZwxvSX+7YXB7rkxQnv0pGzJaB3av0bUkgj/D
olkXE1O4HQtbswvyKz4n0QOYWNZ6dM5JTY0SONvgHyN2LIjGCE2OTmh+lvHDew56
3ZzPBhL2DuaIJDCABEhljXWhwHHFGRsojqI6E/iQ0ot1kbCv+m5IgaAe63eH5vuO
PTV8Br+B76j04dO+UqnGGP66c0c8JSMRlmXn4kTfaE/zrkLZvCJKBoord/xI1BRL
mwfjryeC5tIAWZ11Et8yf1YMNzlwG56qvdFQFKx04FyA7sQQol1Z6JkgyKfKHY23
q2BRf2SGMk9MK+NW6PQV8qi4eoe69090u2VCf+rHwD0wjIGqOCOqvTcXEmGx1LGM
LHXuCQsyx6+BVh5uMKKjezETrtGeDUXSE3aKIvi4OMLUX90PHvTuKPuwJTtsVNG/
RR0x4SVRSDbh85rn0V1IUsR0qA1tUjl1aSbPIrZCiFhw8/D8496l/KKikG5zw7BY
n6nBcXNmNrpJ0p292F29fggMSK1+QbH04rq2c1T/z9pW0h1eDH+V3iYm9bBO9S6T
2QUDtKlaZPdvA/UNoIHr8wvcQLIFM6zld2fb4LmO/R4xUFuDmOrutJjcxhVK8VJZ
vCbmLti5vGlJ2fLRwmEauzttJDVor7VQUlPD/YaaSiPWj98yIYjrgIsmqRCBcPTA
KAPM+rgYlbzw98YM9pC2cB55M30SE/ys+5FXjsokXp3sQ9lC5KHZslg353r9OOT+
GSISP/3M/gR4cwBWOeavcFtQMM7uMEcz99xZ8dTx85nteWeGcvzMyePq1Q2PEqWh
ovwWiX+YwdLAFXU5FWbbyXR0GkPwSyhXEhVy1gEg+qQ/cHXJhbszdCgn7GKQh82S
bwPwHJykKHUg9kzxaR6Zlt/WQBg7zgi2ye/3UcVH4npY0waX7cj9A5wPZ/I78K50
IOChtDKXmFW83sdyQ/AVs5Sxa1g4rHhYE7UutLL3DScIIwxu8wvYZJXIf6iyorMM
Lg8IsQp96dHYaLLvimPpZqc8rE6JtrVs52k8w6BqNJd4yE9nH4Jo/Sv71gEX5qQt
wYPHXt3asNNNPHx4Q5k9LrN43Kbmrf+9wsx+90rwqT/VtMM622DsGi4YUo8d0ggy
ugo8l58eZBH0+xDbZOAHdumT7Kswy8hWYKLKH+mRy5Ap8tHnL4atmchyF9VLRpxC
Fw4BRUIu72wo8xa8CMzfG8PUkDBKnb7LjhFwSliOOmqPCWaSgH2gTu9qW4L3GBZe
4zagwR8bou7bva8uqxdIffPkK+yY8ETz46yC7vMfh7pv89qZ4IBcPYQTPeaPn1IK
8C9ebssniMD1m4UIoqJKRWMtkLwSwrVCfWX97D5YTZizuapReG58P8bbz9b4Qbkt
ovdn1FZ8oevpMl2RCtu9EqdYUOg3jebxDvfgWG0AfoVzHZLUSzWAGKgNGY6hROBu
sO5ZlFDcbM37mumThFGvPDGC7u8WQnLNLEIiaaVBKBJpGmKM361fRU4KwjA8F3VO
zfv0ZM66gZt6zFIbXiAC1ftLhw2Fnyyp9bw60w6OokFzaaKQauEP9qR8W8m5JD2o
vZB7lwuAxjUNmYzO3iWiQpKyylHSFpmldxPyAH0g2UZbapwBDaQpd93+1OjLey9p
zZpoifAXWnImqPSB9sRh2KZwcPgVnTsLs+mK6Q9DLk8YVgyluG/SK/PccYGUe2Mv
MfVVaQHSMi7pP+ljhYP2f/nFWZ/MBrurnFHR7Kq/LrZw2BfdzZo6bCY3j2yhoiPj
RC04f7M6s5bHMqAjxj9LbwGMRwA0UuVHWnVUIqSJ2nWIfCUR3vByzPMrnzA1IOCR
myAIk/lld5aQL7/8xiVx/k809TsEmkKZsAf/h/MfWOH9GY88pYN7mMArXlz6pvkP
JQWG7jKRk63PRhMHPzW+TmietxIsSqAu1W6RSmzMTPsm+GHd+So/g2is5HefWSNA
WKlVHHTkcIVDspTvp8S3e0rshnJLNwNB1NHNVTXJVJBZdhi8H3yI6BkpdICN6iQA
oa7gqo1zX4sUousUlaDRxkeuxz6InRJ3K+9qAc+PgTp7i04yABOgUByBa0/slnCz
9EQEkqc4zh+46HGCkzzNt8RTYk/QWraEGGFmrfmSQAVrmUetEFZ39FFeNFuU7gv8
lQm4gGw7iug+Wwln2mlXF4ZFm0jCQwUvNkdVpkI0ln1ECK1arg60ZxCHpnB0FLcx
p4IwpYFFC96KgbhjwNSYORcikpb2p35oqgQiXVfCk6WtRoQwF4pDV0Q6HGf33mDq
tRjaPxZkZ5KJOP5EUhsSqDid55Fi0F6WbDj9G95IpLPQTrFJ0sfCAcMEUffUAPdP
YnNNk+wS/tbkJhoqU2GNRejrTiG0BaKGDQXZcpYHQlX4cAW02nTb1UwRTuunxtzU
jxqadbeMjX1+o18zg7VRFNNauiqSZ3uc46hjPrWO49oLgHOHe3VtElj6vFZpcWk0
OOsz62Z/ESojyndtTODcXUUqDlsr0EcO4776AfnuKmIuLUl4urRbyWWoTJ8YzpeX
9PqAnhRBnj2SwQe947Yn72fKPHINj2ocWiD5vZ0+Bs1L2TxYpwkpBLiAcuog27zt
t6WHW9piy3mt5FdLXorfNklqgwrrNh0GwumpfTSWj7aQ8odDLy/tLRPXgDY+C79n
zJye4tlBhiW8WTFfVPHlcT9xycu2qn0mPISaUicCaABrHACAtnXA8U1MTwvyqixG
VyxKl4rx1SQWbQ8d8TIViGs4Ym+29unzzzImkkmCcRcf6PplWmy23VYVPJ9AvHou
VY5GlmG6Uf9wJqMDX/CU5dKLTZXQFfl79J/78TPYo7tzdFPhDrbCnyvyExYS/WqU
G4LECvtbgM7jpVfBDk25rcELocO7tNYsRE04zPYZyDr99P0vgSnQXnJFMWgqGAGd
f6JpnD5Zv8psKOBPJOfTTwJFgC/INJhyLhDIrHQ7NqY0h0d7yTjNQZ1YudYpDt4P
dDtNtBs2cCe5kYlt6yu59gh2iPWawsQ7uKrT/B8wxA2UTQtTGjD14dzC8coCc7N0
3ZrpXcNrlURfVEgqRrCoDDJFHQNJQyiinOfpjRq0b/y2KVWYQTMzwS4O7m4N8aKR
nhj4xWejAlO2W8Oo5+jS5LLjiHNnk1XDdM1SZAh5wRDxjzHB6thBYnQWxAncC8PE
mDrSFtygHNHt6qEn1nIoM3Y0lli7YUKw3ah0lfOp0UgD2O69VLSNjWykpu99oVMg
b347X4HoXCVWWqXzbuxgz7a/D7O9BrFrU7X6HOMVmUglKQT9WI1crenjUnt+X3qD
5ZNOqlUQPH3YL+zHyf1F4+jDNFLP+dJnG3tBph0+9Iz6qPDpeDUQhdzUyx+ppqo5
8yQylWQhQW5CRPlqR+ylEmEOIup5ppJoZeIIcn+fAkYRoeFHrIkw3LNU3iuc23hr
tocE1/WsgXCTTcj99KyCJpuZRr+VIzGTXKTJFy6OYGtxLGlTtMFbrpM9bE6YFqrR
LxkHMAIsGfX5lR18YulVh9PmkmuVZXlAWmGOcSMANRG8/gXs2jtXHOtW8RgrEPbd
ATwq8McJbqptsOM0NqvakooPwoLZr0tCAPYAUagndH2VQT+fhzUKEiJnRA9dAcxA
tPOMR5awdD6dOO7U+5i4N+EY1Gro1FzGTmMPMNBMvXWG5izSzjOKa9YKs+ae4Xl4
9XfnZQeAmJTCgYa2hNNNqs1DvtC8qudwwEMqT9cNXnKLsr/dTIEyrvyR01k/Ia2h
3+zI4UX+RkF/E6Z/+1BgGqG/LPiEmfJXs/+WRsO+CNLy+lz/wtLLrpLDs3Lwc7JN
uKkvHM+l9GyTYxi9lb+l5DWjZGDTfASk0FxYRLJbKzDrSIX0NyPpew+EN3Yrsmki
pXD1qhrDhda5DQrCozAnVbToEzQLXPT7oDlZkkfNegm3vQW68ySXOsvvFDC9SZNO
GLKJchCC6OI8646fiCw/XslWzjsHMuvLUWIGEmTQd0mX1zFH/ykeXmXX8OMpVX1N
WMak01DIeE34uDw0IW01pX6L3tzpvMqqMxV2RXlUCmF7oI+XSi/uJGgXcolzkPEA
EVgCdWfTlXWQtAMOEqe3TKR6tnYrdxTdmhVQeZ09YCFUGQoEc9rTKUjuH0imCr6x
KZqFuE9kLI1MbYyBXqZmvs5LAN1dCjt+qOUTH+qv/kWmdcEA3dNRtH3tT//Uhz+x
a76svHdSiGEC2vqr+D8bZsUVR7DxziGpWDqrnCfGZ5hC59F+9UrXwg5YdgJdS1AD
jUP13zjGU0C4J+OiM7SaxnxFy0rSs39J7meI21x6lDobvd9YE7R8NdeFVyYFHsTw
2RVSxIOg1QLxv83saM2y9gA/m6LT2rSsKE+k4U/GJTMPjM3AgiPT+Dwsb0A5+Nac
bVoIISJjwn4bGiJrfKBBrnAaFLSQs5WdEo9J4ZWiFjDmgHunPWxP0vWLtJqPjjno
esVaG+2dwKhPfSBVg4/ZpU3MSCEJsOQNrFna+hW9g9b8rbtMzRQR4+YkTyc00xNC
urZxwDADUOF93frWMD+4lKoAh5iihfy2BEMMT+cZriSD9oFhbrpCZdRI7Dg5V9mI
Glgix71d/CrHsUsKp6yDuGfeURgkYDgSZe2vR9y1jzIOjxQ3BhZNfg5PpkfCDvde
OUieKPOmYVgNOacbmka6O0EFanIGu/z81kq0AOjioFREjbpzftSVOPZVdw66cY9Y
1NtUmj0Pbdd3bEJv42/9NmxBNnP/63csPeOWxn4Gg+yfJMNaY4/q191zxpvNDzMl
rRrJ+PmhQ/L8E3dU05MNmk5vS7ppiBBwq0+N5weAke0qvMYYpU+1gX6RnVnKqrLz
kgOBvqcYzJWppdzR+PnxvgYrrlpX8v+S8lm5DjmWL8Y4pFR/vuNtDhARdM6JFucN
ynh+znzG08YxIOOjhkQ8Lqyk8ed+6YmsocSHUQBGpFvifTNUGqYdSS3n3IyZI8/o
mzQiW8Pa2uZQB2Xgh4L57N7CFJmBsUJMHoJZOvIHwYay4gpdFbMav6b80VF5oAd6
hAfVRdWZ3isTonzJIX3/0Uzie379kJT6zUIVw0LR8rh77ttzFm9SLaFojxSQ408c
4SkQ2J4Tz5eqaTS2clncw62/6YpRQEHDRQIgsnI1hYfP2BS7kQTeSNcPPvL7ZwS1
pWRiMMhb15SjwSdMoADAEOy1Z/wK0KRWnKl65yktgyma/9L5WUsqMwxTKtSuWD8b
TsSYzVHzlCyfOXIFWmO3GBXT/B4zBa56xaD9PwwhnYDWYZqaDUz1WfeGuU1Vku7i
5rq/ePvF/z+tU0xFWiPfk8mJzWUTt5dldLyxfCp+ziIux7GTv984By+acuPz1kT9
+4sX2vvJxSOXBM6fj6/1SswdO3lGHOzjMd3snBtzfpqkbXLNEj5JDnI6z4rvWyqL
DW6ePCjqHsJyPheAGfLTPLO8t1pLM2Lo0VCNchroikdLVbrqRb7ocJD301OR7SNr
ZuvucJ+F1kDjsf05Pn1GuiHUEKBY4CqAruRzU9DBm5nuCcEdrQDzYnYIcw2ririQ
on1ypUQNsApUwOap4gHS/WrRkifJxxYGl2BKlXGIi3t1u2qjLYt3QOfRjllgo8ZD
ahtTYFU5cjgWvsdgBOgCvheA+sb4GK3LQLmNKNrRw218vAxlX90xlpWyolZ7DZ9R
ltS6NMlTdjLZM5RXg1fnE8YDcHCMhIR18mHyJFww3M4j7opDTDlLbOwujI8afd38
KVrsGhozLH9l9q6VHLLNZ8KjbmkFpCpGcyVymi3G/tFkxcW7nHnobCswy4V7o70l
XjhSW8kgv5Fsg8zD+aGFag0hCKY2hx8JRoZ8RDceJqpoyeOZHMAbdSFT6ioRw7fU
8aJmSeI/1fEdgTP3M/kFJ4pun76utnA7EKZyklahPL9Ms6wgVdxrwdnOKEzsiomH
uOFpNxnfMsuaCMhA+E32SWoog+xFE8c5IrZXKzMLusehAd2FP1VnJrq56j7I5j5J
IUzQ6mybmj8TVulJTeNkqbR4l0xbEv+FEPG3AmvB9+BudKfymNrz9QJXVBrEGXvU
eybN3N565plpIrp7AIKw6cJVlw53EAxY5zC1A3gBesHA2gjAI+dYJ8iWxdqm0g5p
9T9EkVUkQNwxiY0uqkYJvCa11GXphTAREL1R8vALwobwrN0if4uKVjvfW3rTTpcA
2Ia8Dbhy7iisrItroS/l27aIeWR/FldLFhc27XsU3y/nXeQdyFIy0pQj3hJpcpj5
HHGkIEgT3dnSPCy79uc5LaoVxVW8TW1gwBUxc0e2hWjQTLSs/O0/LeGjZTTJo0C1
RBIgoEgJB6mps3wBQL0RCmf5N6GnbYF4LBTp5AB0ZLsmc2sZoybgumbvOM9ZLAoH
F8mUBtxfhdxOPx21HpNP8VTUX/1YhCMd4vh+ciKNXfeoDFzg3aeY/s1zx+tFVZuQ
9Q42drpnEHPKT96fLy+YWJMWWS62RdqLUKcHHd8nowR6SaV9zXy67WX5gEoGqRZS
1ej0+kjg91CNCULbLE06hGg3nnj8iubSn69ew+Ug5W4lAukR7heqbkfHZKOKFWog
KunXUYMPMjS3SBl/fAIIDHRuEuDTrDanJpg+RrF7alCcZYAxGl/aBQk1R3vyEWTL
koYFoO2OUnCEB8RVcw0FgB3nvkBSD7n7FTg4DUcpTbfn8YdJdX5w9fZQxi0FYt+z
dm6OfsAfxA+KlgilpbpdWBHW3hlrPyVEHO9YkUALRyvPBLA7IcFdZC3TwJyPBgqf
9zTMjZ0sXzL8IFA+JLF0OjeJr5hw6bOny7YeU8DcpZciDZwkTRcDNTaRePxw38Kb
GOLPcs0QX3wTXii8ZPSJFO/bSquKXO3WqjrD+JDlhljdU2b1MTuMUyZrffz6nBGZ
rg08PUJbPnPWQYaq+WGcYMxQLpEjlAcXs9XloYX2qtDLEAt3VpI3UnTDYWawz4KW
sCg4dCGkLHTUlDR/xGT2DvMyuO7tHMeCaaLnz+hJCD5M3jhl9BGkGOfF7AxoPdi7
hq8cvRyDtt+X51vTeZStvBkSOTV8u1QCDI9z1C68nibakmJMt0l+qee+oNyBUXIS
9veqC3KhFGz2AHKOC7iHg6Hi/p99byGQUGJ1TYghN/oIW6n124vkassRJ4e2CHdV
NRo2VgyDQw3vcpGDS8TBkVaMOqzP83cqx2jW1sSpaWRSncYe3vMTiqtGn+rXnPcv
EMIC3J4Z8Q0DBLaa1gNroqf0EvKqNpIeT/VAwcMuPwKTM3D5VA+00xxknAhv1Yx5
b4d3P4Rw7mj+xCeiMQTDcAf/61X+tT3126iKjUysW+3IZYTxLwd7Pox7wVfJBE+9
booCS/Vc2cuAC0+o+dPxRRrpcO1Z5XaHULHfPSyWtsl8vAYZJ4NdPt7R7pjXHPBF
uPCCjB9i+tBjHB+nGtfraQFckXkZR8EGbt8Jr0NZtJchy/1VaSDZPqhQtEMv64vu
6rY/UDhDHdJjeXb17vw5kvxzFme7azea01r7doC/n3U2Zn4n9X0Bzc2Gd5+8vhu2
Pw4jvgq9QitlW0gfy2fR8K10hrTP8DcGgHh6vVJEyHYwWISWlIsMi4OIEylmk8jl
fH44iky7MXPYGup9T2ITMveahw/Cdgd4CV2cBPJ9E7KRevZdMSbgG3URoI03Bmno
1k0tUyOeA9ytXHzvAqusEBTosw1Wk9dONeUPIpBRdMDKZJVQoxLaGFsVA0ZB2drr
K5uuZVRuU9D9lP3JU7apgO7JGlcJirGMU0vfKjAeQL66F5107N2RUbdO4pjrg/pj
GBq54QlBo63oqR8I7Hpd6SqN3LOCm+X8C8w2tz+WrSkfcNVEGH49PCz0GM1k/S4N
Km5c696KhZ5xaOiZ93lqFA9DEvYUyO1lHBIfO/+DEHEcp/FLXRU8uJXDN4tBJ8nd
mnBLG5pwx5Vua5llc8nGuCUxcjytMgEJvMa4j2jn8ye0oUSTKsOW0H5byNU/Haiu
oJBlJwQqPhGhfXiZWnnraBecy6W/RnyzN/UXXo5MSfVGT+Vm71pv8uQPslD78lNI
NHJ9O9YncqNQyOYmA0MEqIzHsH6xTIMbx4xd6yRvnfYIId1TEdEMXGDivKXC/xgB
jFDnXadvUqdEo+5EM4UCm7sp4/OK76nE5V8omsxK9VvapVwskQiD6tKpiAiegucN
EOiUNJaS3DofpBSmC+ZNsAzVewFM4JMbYlyu/zngOYGzmMk3LH3sWdWjRtjDtjaG
HcBsLOqlzNZJRi0cvNoWX63dvkEH77XZRR+utm8GofFtcJq9SALdM2DofCPTHcoW
gnPELuauyvhc2LJ4S5EkzBhzkieNUN/pSxK1zkT2d4S+A/RyBTkYitfdV/ARHxBh
2cmNqMECcXs0jc78yQ4F4SJeuRAuhqty1fRrZbs+yEEyhigYSLqyGDIY6vHq9g0t
0G5MPTE2KY1v3WLSxDuQEiu2l00qavnCY1EG4rMAC9S3VKiQ7ni9Vcl+WFjkRGqG
63F4a51TlglwfnYIg5OMuvviCtn8iG7MOtTrlXhtXcvYsJSozdMljl72g8nnjQur
fj9k507dLB5jr+TC1S0R/l6OhhQGAmm/BnoSBpJq1LT7ewtJEsMHmDJ3yvE2SaDi
wnFnVo+vD6833PPrBoSk9ty6NOzS+CVB2wOH0pMw5gViM/iv22Q1/fb3dm5Oe9c5
Iyh/lMEtnGE5VLz25wX7UGK9j6/WMKTymPLiq0oU3VJ8L2lNvmpDNQj5p6W7AJEM
g7bj10ObuPJ+hVuSl3XC2T4lkfh20bRIcfFB19PJU1gzcdCoz0uoKh07nx9qu9Nk
tEs5Usv+dCFV2K4mV6G8UlssJksC0rkJe1CsanXfPUQ84qGy6U+yoCRmXgHOo7WU
/0CCXnhl87B/4qZnzwT5McGDZQ/UprCw3BIfqUgDdweBGIjRNSMe3hPf80dPplJ7
rBk/LyFuXTDd/i9o9gaH5+kkH+MVpy6/7rkziKdnb3FWnVIZ8759w0dVhLXgpxB/
Bvww2GOdboy1KsjeMAeYqiClaWio0XW8foTC4tXiN8j8zTmNh7gNxqXMX763xAxe
G9F0RtQ81M5i5sU4ew8+0E3uE+3aPKsHhSTz9LcC1OW0pdezbiNR7qmWIhR1pTsE
nc8N4AeLtwgARL24pF4eM6LgySoSHJIOkgYcloqWBnc=
`protect END_PROTECTED
