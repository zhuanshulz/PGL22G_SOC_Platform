`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E/0UvFun2yALtCGLXyh3H705nHew7iu/BvuJk8LFsFj853iuq54SGoa9wVRAVpbd
NO7POHRhVaqK67KGaUR1RcQT0REpB7BIrb+Mnkxi6KAPOW0wcnrQs9b2kDUEptGA
EbQhMT7zbqw5oWKoM0w53z47sW8/wWDKsuuuxg5GpVQVyxT/pjhhVR9gH557SLtd
Bnr5zTmK9xU2mKOfaErUUOpKRZiZ9SQELQQFxN08wyD4OJLCxEaSWuJ6HONHDsPd
N6i9QG16iUvrdKwrPhqzDc40yvna0k8Fbk4YG0i4wZRxVzrS/HFp3+Thay/jyvJb
ZRc93Ye4naN0SIMQ9qFWdhtR1oWf5iOkEKCQpnb2ofv3QCGtxff/h9wgRitf8hTY
B+LVqqTk3rx5PPUe0QM/kbk41pKi5uvxvbm3qKfZzu60Y1IYcfKeR+Nf8DgLtueS
K23LV6AOiqI6ChO3pFmF1/I+av/tCDaD3QTM3jtoA3F2bJAzaYdeTgPNdxndMiAB
KnuMvgzIvkqCc076Bb72nRkGgjck9+iLoxBMt+Q7S2AjXzZ2BbxH1jf6gpenkMyL
xI9C1+tUucAPl6DQe97NgNIk/llKl9eSflcJ5QVjhEjKrjfNK/MJ3nQnRNBI8B02
/e/yCZ3OrZ/Qm7pvfmwuWeiRh3KLRCuIzrLJJJIKPMSreSfcCq+aRoR1f0bRP2FU
wb6yx6RQIBqZQRI/T26KWOF/1Qt3xHJy+aBLTGyw2gdqktNIZRDVh+l3gwse4+JT
pvfXt16wz5KScmlmvhjKrwZeNDDyLtuWJN45rg0xw/3I6tp/Mj9VjWGgxxWXqpLl
LVyhvMbSHIWLQ7VDBXG3fux6lQS0P4Z0lXn6vo+fV/opSamoByGx3Ah2vq3mV2tX
`protect END_PROTECTED
