`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WOPN0ruFdFpM3ykUqP8+mD3TvN+/mtkdTZ023jvH4RjQJ/baVEiNE+WQv8BBoKk6
RQkGidiTZ75O0wu0SSzHpBkoXjAUT+e+0CMUi41y0LWoDgKVoaMgDVWHGGiQbe7e
+RemfAGYosq+rOUuiLMaaZrA5VVD4l4/egL9gcpnBlfRAtPTIZTsVBceaw9aXlkE
MQkHT4ZACSpPUhd4lPaU65MLKaRrYg2/zLZU9xJxvEHJZrLl4jujpREwRjDqGXi3
zQY/hrQz8JJSRWNA+zAwvxrkTgxwI3Kohn/0B/UwABCEExqC+8EBQKxAiHovC+W8
KMD0bBsQs6/ftAc5N5YXkMAoDm5jEyeRXIybMFFzYqUe8MTmZl90Tvs4P2Y0vjqo
S9eiJSSH9VuQavGP7lWymTjIhsQgX7xQGP5yeslcjdQOu2/kZfxBMNdi0xgx3uhe
AABcxZX4bYa8CUO9Jh9lbwfSYneUvi5l+BL8DQMwkUDVHDb0bmAklpdRMybxjB5x
atgLucUgMuu4KnxUv20J7NumTd6M8gN7RSQu4P1aVZJUITsU4INrUSeIkb5mYuHD
NAz0s/lVqfYiSUOCEZm1ix6h5aVVPrVZBuMV4aStRfwU83Fj5m3aj/LNCvkYJr+i
VDd73MloFAukyjGv+B6szgcn2qdu0u7vWWYZsGOgmz2uXnOMAC5ZZgDllpGtEmLL
IifkzwCemM1ZbJdtlA3I0gkszqlqN1AVjLPygvBMU5+xkPFyR91RoOrF+sJmsF0s
OxaEqHYkJBMHTZELwJz2elRDwnCN6UMRCrlpiBn9LLDRQ071XjpI3Tcq3iDgWsQA
7HZi5B16nQPlAR4iTIDB9jFHQza3OOk5+pNCxaKP3Ecgou4H4R01fvaxR6sR0tNi
k5TVl6RHn289VjyYoR9lyy/DTVcgMUyB6P7o1abrw7IEw0wprZPP3c6s2X4WLD8z
Etz6utSM9fRmVqGy9Xu8YimMs1A+yyJshk0Z4g6gTxBngUl/WCs6AJunHcLKoOOy
7/N05a52ciNOqGXLW+vYH42riGV5fc/zUQt6sKYj1IzDxKilGjtGb39GO1ONPA9l
ywDe/Bd/oLAYvKp5RE2TdIobo24RkRl0VUsEB6U7UWXNTTvPLYeXcSPYCU67qQ5/
gmoWMl2zlVqA82Ku2Z6ByCRousRMFv6m31IAgTdqKfSgKwkWxWxUJIYNHiNBI7hi
GSrhM3CsA5cfOGKkPOvUQoD1a6dRNKFY8Gf1+qxNDtw=
`protect END_PROTECTED
