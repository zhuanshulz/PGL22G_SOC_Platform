`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j5yz3vbpKFEOtkcKbXokdRriIWZrmDzPnS+gJSMuFKym6QLi4xg5Q/6DdVbDtCyD
y2d2nCC+gGMGtIULSBwEC+wzEYuozBSMHtNbBr6PS7bU81H1J3tBZxZ5Dn2UibCM
sT5gMPSDcearREb/raPM6LHGun0zHs5HyfppnHJtalQJbChFBRvKyAVCHKTVno7B
mP2Xkdq4J3M9ZvtcbgOuM1v+kmsDrAidBwH4/4Shm3f6P7vZVLj8qWudyjbRigxF
dwSZ3c4pPnrJRgfw50XJZE37ZR1hhOhzGG92kKk+hAFFeJbYJu93LO5SyoXt7QtU
QLYFTKGHd+nRF44qVqzv6W9MlmfTqEy/2C5RTjCtwG0P0AcrqGqONZ/+1SbJG6y0
2Cwi91TD3aMJZL5ln7lZmxJxBT8g0e4NjwvyQyBWp5pW8shkktPDkma0RLiDX3E+
54mPt3j1z9OSJNIGW2SSt0jTiG6bf+/kxmLeLA5IkJBLCTBoXuJ6ki+5EcO6LOhS
NGao4P1F2dTi+1J65Ym+LD4exwxKBihGlcK/DHjBrhnCJ4wurTr5g3QqUep14DGH
s94VnOD3QlbAHnxWutphZGTREKOxUa0qyCvaghpYCnCbXt28FUbUVOX2Y0V+EtPw
+8Fh3jDAJqoAqnv6v6/BqQ==
`protect END_PROTECTED
