`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L7Kuuwzuzr/8lnw+cPSc/FXlnx23W7teAn7TfUxgPT1YdC7/QZaztB4/36ptPAeO
5bTLmjspGU4tAkpSY4T1BdtSTglY1lKacYim+XkXaqdG7QB4zhvBl70VugRKOuvG
CBT+MR6y1DDXUTg4c8N73GlzDUtwBaL/A1ZPYPzkuxnZaUhvfGokCXC67BSyDtaA
CyWVffzojpLmw9V3HeMa+qHsiEv+7TW+0q1xSCtvOkcECxOzBOm4bEWJfweUuTJ6
IftTSkUbzncaBpxhZiQMjO60oBYMMfjNwXnGO6scxH8gp+ty5BjaZulc8zR0jGnS
wR+kATf6TwEJazFqezTx7t7Ci1jNdtyAdmN5sulKzwfl1c5P/0o8eCnj2dKu/f50
rMFU0H/vseiLSzJpBMOg/cQpCbFM6V4lHanhf8xE04GaZ+iYBYj+qNGjyK3oOb4E
CryYRBYUIqVV1QdQwuGlN3JIB1kUtug9cD2SIlNoTFsYCT4Ym6a3t9vXJHDaAv9L
Af1I4iNQuIlsyLlDQlnVymKKCN86ldz2LduLiUHVcdiRRphX7uzhkYaP8YKI1wyC
5iuIvLdmKqYvpNjDWYZZVpTrrGRtlXq5ifq0aiHnraQguyAlVAKgN3sFTJFmRXHZ
Yd8RkZaLEvNZSZYu+akicDoiJjjeSziePgyCpNajuI71McBHMemwoSWxM9Z0JzTP
vxE6VN6AJ/AA0BYeL2/LXfOYVwV9gpHGOrOqoV6zVIh0QBuG014Cp/7ymrbkq5/F
s6J2sxQI6uu3XzrRV7AV0Q0Xx1Zo/FQKR21gmMZhsNgSNsK2Mh/2Z29lKpTEdccL
JiKjOV5kxE/4pQjlQ/KYQVNPryt0YSvhJA1t6b1nd/qENwxSK/9492jDYGWLfjVX
/J0b1zhN9lZIcC0/o63H0WVZTuRjqJD1Dzw5HJ9m84fSno80bFyr0jB7ZqL4j4XE
9VMca46vgAyZNS1ZlwZ0I1fR+R0uRou1YqkJFUdsH7j3Izgd2eTDJDwedHec2xp9
pEq7yYl83tq94/+Yp3JVzm2rl0ya8HtfgNbhjncGpN0Ov/2j/1vzMuji5fQbISea
Vivl3q8kedYk9y7+ZHTntUOG7MHMSB5emNk/cZIjeecTR/Y9Tag+528reZkccWJH
HRghLJLxU6RFBKPqxxmDxzxdASKOepNExDwATpy4pzFZngdSZf90kQOY4Al3gOL2
mCRAfg7kawQn/EUulen5p19b6nMDajEDGWceaXVOUxqUyY15JRPuoOB5SYxIFu3C
jj7Ad4e2lpLIRyYUPBofCe6CWtU6uT1/GhIattAPD0PHjJZLieSXi9nNcuwGtpmK
RwHjD0I/DTmbS1SCG8jh/ulUw0zaQv0cotAND5k6mpODwcq2SZUFylKni7YVGjSQ
bILIun0ynm3X8XJIzQLAJyRGPgIicCKDMi6DSTvxBoHILCfZO2MAZ3oW1zhnheOb
PBQhzq7csH01XEHfJuni3imH6TL/jBqiSQkM09pLpanW7mdkl+fM4i9wo/088Qg5
2YQdwaXCguGrjfDzYBO6KaPO0GB7TQYg6GBkPqEW1F/phbFNb9uYxqTmA1z2BPh9
fqI7mcDaiOoDFSmmXOgaeoSRe+s+BQIDD32ZQtHzCIlou56yEUiMr20MZVqXc4xy
URiZG0OyL5onwEBkuq/Ke5CX+8/CA8SSTWDx17gWZKgD2pJi7nzfIjrivD53Tliq
CCAj7lOqFpR5rwelfDSJKVMzpnnZrxf3d+oGTLM+3bGvy4wil4n2QZ3KhJAzQ91p
xm/f58HpkV9IzbpDXBUIyARkP1LS3/g6TsxOTYyNRcwCFEdZtv4vGan3K8SubZhd
4MVYDslZZ1mByRz5mg+QdPW0dlOieoDndI+3cGvLVIdmBjoDJeQrkEPXFRKbTiFL
w8pHw4ZeE1r6MBcttzY4knmOq68Q9d9uU/WwNwD77tf40E0PzJ8EkwstOMkgtcI4
GUSKBS28BqbRMvd7ez9RcvQ/g7Y2MqeL2ucLKCS9RCRm4iaW+G6d+Mx/fJJlqIFi
YAbTFqYtxDoVpf6LnIONnzwQ/1eohdW5ubgBgQfVwy3c+8RGM1j+M557EYWxw3RE
SOJPPeiHw/HRMZ3FnYKDZVO75i+HRcsH2CbrMubjXvdSoK0KsD0R2NGdBRrMNvAB
LFARk3INIFjtrA/2d11OFlnkfXKEcY6H8aPWAecPBNJpGBlqxpzhEwUs0BIxOD1o
APsXYWJwsqLALYnShoKw3l0oBT+PZ5VbfrBpe9kfH8D6gdkKmRymquvQIbekB+aw
qi0nsOL3ENi7k9725ZkKeE4U/XqIUZCJY5TK9LLcRtM2OKV9D1aQh0t9jB94ek8Y
FgAjTKlJWtmfZtn+XimvW0a72eT/xzsE2zwygAU87+NqfRkERC8/uV4Cr8l/9Y5k
PRUxsVCkki3Gzkv5PTW3/e++d3jsbib+iEFIvkuer67YBuJWaYqfxtZZhGKeN4fO
MPryu7i00o+fVIOhZCvj0I+qTcvmdAQ9/1bRCPLXGK3F5SmKun2es9fO2P1nDlpi
kVGBXBFjLirYleY0GBthxrxyM+XjmyRxKCmIcaf90v7sjjq7UM7IrNJL/MV0nPct
rmg4gx2OAt/97xnLYi9xR0zQsHauXODF+v9yGdDPtKv/7uTHqAsGf+qOja5qMKYc
NJ1/Zem8PBA/tYCI77g4gLFKYlMOmLTIYzs0r4h/rpyGTp7Fp5beeoTLyWi4iwnD
gyVn48l3/30INh7CxsGARdvCnP5cLmNXjUrvjAmU/gYW64beswLsaBXsAiLlAw8N
yS+9gGHY2iaHBsmnaW91iWhIPRnJjgsE2NqZNlU4ADlDjmfxhFzbWvOeGGvNuZfb
fKca4xhRQcuTPAkayPPRG2uEHAF0bqodxYeUA+MhRF4O63PvqjqHjf1HVuwdnPyl
bO+lJU3tf79ok9ZnLwLt7aQVs3gl5SIqvbS0W2B7zkXBbClP7IpD8XdsQIe0HKVe
9Ls+Ruz/qOKlv8J6iJfVBJadKkwXeL+B1JDnzL+vWbsSRWEv8qIlHU5jNtuPp4RR
BH1k9/7wlFkZbt1iBeGluH5Hix/2AgH2Uyq89K1TfqCuzo6w0tTAIFgcB09JUVQt
qo9OojAkDwXejvGpQHbjRuU2JAWUvj6DcKGLjMHfWfKbT09EpBYDHASpvsR7Bo1h
OoMNjauKSUB8M9eZQWcewS/wTw46R5rGGdkm9vFvq7OCjSu1NzJlgG/ei+PjrhZR
MxmRcO5dwQ0glTN11rwnHWzdwoETL6RNinSdaP2hi0yJDLcto8EItpu2UD82InJv
enrzH1ZjGp9yt2c+xBBN7VgjuNaFsC+cfrd2ln7lJnraVPuM1wbaJoM8y1d4X4EI
C7UvvFGIMbbcZw9Oa39oMZz/C95M0Ad2XaH7PoSevkuiGceF3TyCI5jCGBfrcT1X
sduMf8pp6AR7wXawV4HiOVSH8xiomlNll0TkRLScMj5LNvJrcLrwgTnWdChJD/qQ
2PHxJUR55xw8a2VDj1okUM5HuVTsLkOfSHJTf7QnkJBMPuYjaiJQKbGAjG/w/ZcU
+BFgvWlmLj5p8OMQTk8kSf+BlEwSUknEVJg201h/yYXR6nALwRhD4qR5eKsrGn0G
i+uClLwJmjSmFos2x3e+H4pBrjESQBxOXlSlvQyK1gywIchS2hF2wQ5fFxT1drT9
kRdwgorqARNByHNSdNt5rg+YxxONq6RICD18sWlSLMZUPhPt0QlKXC+TRVhD0scz
foqj1odnUJhDY3/ayDObLdEJY5LKoZujhJAvVpH9gijWcwYJOfukLJz6oVCvO7o+
++FuSVo9NITDo2oipIRdTymv2XLbSD+FFp9LTqRxYx5SEFhcCdjsKx5cAWuUsvrl
YO2s7GMrUd1xf++Kb0FBC2G7UH++wMOlG7hvCKWcw2Hvz9alpkmzdml4J700X+ko
HKYUhokyONQKzB/DcWN9p6g4b2ASHRKrs6mArIMloJb9wM4zYL/FjCkJp5sTK4r2
WK0vW0B6eXQSYnPGdzd1xiO9v8Daz+gcVn9og35nFyGTTh6qL8bnSTEYEg8Ix80p
ZfekRn9CCWTAmcxtxzdxtXZzQFqd8kDh0AeMEr1JMg/y0Ny41tViZCON7cJGvdE7
3VjMoW/Z6P45EDVXjNfb4kmS7UqKe+F8peQsKpMvbUP+4eupfnIH1B4zdD0Ku/2B
uy8Jxpffs5fLDxMx9p+dNr203RMCiSWnz5eGbGAXSWxD/TDRYq1rWzlIEzzVGaNq
zQBnMHa8PB/A4RTO/5BjfCKgielp01H9/kvOrA8y5jUaDUSltSJa/DiUed0rcm6D
Ij7CgIbyq1YqD5yhpzZeRA90USI8ecs2zWDXZTT5piJBXN5MUv+BUqd6Tu1OBdj0
xLnwwLWVpPJGI1KzLNZBFoiJ5bZW/LHVGmXQ45EQdgnsZJI2EWIJOpe58vHj2DuS
tpFs4BfsJzb0a9rAwviLAgpiTVEyPV8BH4ax5RXqzUAtNXMmGA2+jxIsKc2S8+Ku
VjCi5R6rrycJm25UhoWgEu6dnl3lIUuDUjjMN/bfTxrQ1Nx0pKrZCgKAETIzaw8I
/7MKuWPDI6yiwRWZ9Dtw9VJLuz6zbO9JzZG9epVhqhj1sOJtklH3ZirQeaXT+/Mw
nYC1ZExQQE9phpPq5xqzUViCzvxJepKexYUt427etUjke5Ls9sUaH6UJzqBuyv1O
Qz+TdYy3FuxbvNK7dvqeXc5yZsdeqAW9LJCZS7+KeUOwy9PmMVkPO11LphcOouuN
TPHFS/oa7xggGxXYQp9yuNk0e8Xp4c6rLFSfdUn45K0ycIiY1ITQD3JADRa7/C/k
QbYlLI/dj/aOfw7/Ovv6g5SemLaC9VPKlFrH21vC+lJe/yXsOQNmZ6z4WSacDTYU
DBcK1JoWq1da2Bq9NmTuwW5XbioBDIw9ezvDHSNxiT25ARKg4vTKkIvcEWM4G+0g
KV3CNchqT8UKhVJcBgG8h+Q7dvQWNpb7VRWkw0Z3bV8SpkfpXtwQu5y4J+aDpmF9
iuMYhWYdHRV21Y7dVa1kUqEyA1MjxlpOubq/HLfxNLNycGKJ38HFjQ+Cg2UEeWkk
eGDthID00QB8AJSJJYFXSqNHwr0I7dZZqdvNxd/ReD0X58LIDrGLdsXvOMqgWZ9m
YNPFk6yvQ2qbHj1YBgvImM7QE9azfZRXFqAVTt/bydvwr4BP+p6E2EoBrCHf0dr7
wvJc5YH+Y5XXn8npMxXqAqVQQFCaccomOg46cBvNSMVJktFAvM9LcT/EqQmyfPnq
dCG8wmnCNDtp4w6W/PiJfsytgO+sLg/qz3sVZFOW2ehwU6XH1Q888n6x+byhgSkc
tz7MeQj/eArgNbmbPrf9gVL4h41DQ/u0dfBfrONVx/OjpqkhsJ5D7DKL6p8CiHN1
vDkhqPMSLxlIPC4OXTylK7fVJB+tNwe1Q5ya8nt3vH+mYPTAEI5ITq+sjP161Ly2
ki8RnB/aLbteO4UkYzMCVODH/mXutQBVmq9hzxNrw2hbgsx7GM+GAPz92Q/RzlCl
WWbcDS6T2SddgM7LuZWP/KTk7vgVBLZKqe818n0nKSO+OqadosaaHVcsQyttNb9M
jIiCLmpffcP6RtGZS4E7zFGsEhODLrGJKSs9Y5NtqlA2eHbZt+CoixOiUP5/X6Rd
aFS0NN8s0V42Xupy7a/H5/TXIwkG6iPWgPsZr8Z36J0V/VzgyHvFPPI/aSML537v
FpFjFAG+vEsUEC8QI2lDe07OvqaLY73Pt/Jo74L7/mNhxohzdmflOMjWROb2RIM+
iUHExOzM1HHhvIsRYqVOrf8k9ogc5LZi9oqr7BGKrJgpelfQlVVS+uiX3rMsZhFN
+3ZZJltXARPifyVWB+RcjvTUEMafFaUU9JKh+8+uhIZh3qjGB988Y+ygPdpPmNgm
eNjmDDTy+oF18YEvgaGN+soEXvS5m93kXMimO8Xu5IZqlXUCf8Qhye4UHkARFdDU
bd4P98502Mzf45Mztl3nc+yrhLgA8db5py5BAvlsgepiYBd0R+DfOyhd6asXgPvl
0NTIpq3Nthnhv3hfORWAe5AQiVMK8Kq4gW5Bn2zhZL/JBNpc+XTVpDu/+ev1F7hI
zp/dBuXLl97aB7F51CR6DMWbDKnKPwvTIG+URYK7pzGdzZNuDtXJXAMu3KYenQn+
1ynOODgHjyOXe1rZ3NYrjs24Ny6yHP5fgwFhwlwpcb+KAx/e5/qRQErs1N7AgPoS
nYDEWkHo90pOvUU9guJojG01AasSBAdNXwjbkE2uve9nN3pdp1cYww9iMgq8tVBC
f9fwjNvOppZVjgUQd+6+ZchhCtsKCjZrH+peAGDDZVvDJ1XlPYccxFx1hTqlbxW3
hPVNObK5JXXuUvbuoPwbZ3QfDOzuXzw86ckW2KGlFkW6AywXvGyhBWJPoJmi1AX4
rjgCqALKovROsSxriWq0rj+EZq2de0wMWDroMP+FsW5FS9CXne10y2u5wOF6+LlL
fC4760h7YJGDMiIhjywT+uMG9VfeKqPOpACfqUquobFIpZFLs7yQOXbq79siSX00
FhGhYVqPS1/OaSrGp2VUvToaoATCciS52774nhZ9AQs5bkNixvBsS7eXwyfpVb9g
AX3fNN7NTFjI5eILqp1LbTj+067OGgDFVopJ02PoMj49WHuI7C8WJVlpcX8N84Jj
JDu6/sVizMFIhG1gUS8kvzA5UTDns8A8+fIKpSIm+2bcUBp1g6oOCJe7kpPp26Ax
lCFOu3q74HBzcZ9Ks2aO5uvv/8ej5x5NDEsUtGDDUowXnwvRZSt3GwZBxOpIroH+
9hQTVX8FokGF3ktFGy/rRligazYjAsaJpQ2Vy/4oKEhblUqVvkgYqRlidX/98n12
aImTti6Da9YvEiBxhua8ptcuf6jlSC4gPCwBQ+rrPLcD68nfhDQuZ/V3y7nb7XGI
wBpzDJ1TYXTLTdpnn2EPe7ATl6Ykogimajfm2D77S8uvxiANl338ersVfNYcZGWk
RwjBuONDDl4uF3bvYTceNU09lSOtTxu8vhU8DJn4hG3ZavuG3shMqNQ5uYrd+/8z
IgJIxE1ipU9yJZO9AHHpdxTi+mQSLzS6oT2riSTBUye0MlJM45L24iAbMl5XIsd4
EHcmgGXBItwNCh8PR6Y3hr8Tfma4n4JRp107vjF+0jQ46fhvwJRNkAJmLHWd5Wej
fKktMGahAGZ/tJHZI2A27mhCLf3ain+NI/pCs7zKkNo0b8L5S3YRA4J5YRAy6GOv
1uA8+mKAffN9V5FMZ5p/D+QtgS/GtLc3Hpb4r3VW7PyBBWrZVXh1qdMYj1MVp3mC
SOU/smvs1OYyKulygWnnVtePz8yGAZh0x2Cbb8r49QkInKZxxJYWw+47FztE+l4Z
sDCIsEPJ3nCC6l0dhj3bHqp5st+NcNnk+ZiIwn8V8IvL5rxV2Wqm0r9T6xzKuFm9
Y1+rTKX8MGCP4lb8eYdHJq1Jt5DvSdh0aEcgJlN534uu9buSu1xly0wIvLlvF5nX
algQuEvTKXejkr+WwVf2V9fFdpm6/qnNH2Npvr6g2LzhojHL4yuxAzOOfVY7MGHd
qBqX1TSuiu2KniPngAGkEUP5U2Bcts/b/GKJZ+PQ3DB9yxl0LYU6j6LQwVJ6iqqa
NsoS3UxUMkGDJ/gege39GtHcun/SWGbsaFGNCfYN9Vi8LGcV1vTlT7QhcW9Zq+B7
MacCxXD2FM5Aaew17xTlV2B6XlVgm/DgohRJeUZqOaSMp2HpWCdfcKQSodNoXPdO
CfWeGOdN8FMWbQx8g0HDvyekQbb41E0mCOlqjbPjWCxkTUa5JNtBe7yIZOi+ti9/
z+6iYaICFeWzccuamHpnJlIbk0YziML+x/VrWWXLdF9O4VfHDyRiw3B9GnICKhpR
mulJW0PiEFhZ6HhX68DdfeYa0zQpYXRO8rwriTLhrVR2l45DaWadEpZZoN2UdLSw
bn7w+WSReCKs4jycmcOl0gs7Zk54T51RUwDsPY6bQ1iXrT2KLSuIKC0EcOARqtw8
Kg6wz69SZT7EolUNWLNer1T2qQ7C9EcHEqF2MXENg/qIBVNox7wXQ2jyxda6oQp0
Dz4wixe+cS2U35bmqITBwffQfc/Rcx49wibV/wYfzPsesC067ZCzN6lY5JJy0IBC
NugDx2ekv4BVTb+KExD2Mu2ZHNgLQ7uYAsx3ux3HYI8z9xXyHHQ4PPsiN3Jf8Ghr
1k43kBgMYLKTQe6upcDgRJT1iz36rTTwKhWPAlAaqYtjVZruKGuT9AInRqvgIQtc
g/k5yswBqESwEbYTBJoi1U5sdovlJQTgbl05Hc08QMx1WM9b2BPVhVAG4aW8h6Kq
sr88/EGzAWnHHjEmtRjejgUxS8fK54ZdhE+kKYLwW6Mq4/qmZem26QeK+yEk+ZST
S1vIhtJU8ihxmqA0VZktT9J5uAKSi9OCrjAY3BmvYkB5NCNKjauX24bekBObdwMF
T4pmi6gVgYsOn0195NLdpvgcCSuQKuRP2M2Ff/856TRvgmhCFiSwhBsXyQyfJYjW
K11r47oTnhn9whnqxWylO1FV+h00ltfXp7KCsvsGToeWHE+EcqkUEGRDQt6X3lq/
HJ0Vrjm07DyZHiV6H/pyz33OHhdD/cWXZo8hAo+Q4AArz4Wgt0DB0SixV3rm9HxZ
Zxkwh7yc3YILqg5EXqairRJprUu2FBR9MuTokE8Ms4BT9BszlXOSqgkX0sGkYDxW
BqwTer3Wle6X7wc1mc5Ku6Z7w+KQUtugb10EyvE/O2XH8vbm+APH9u+BH49lbzkS
7m8fNnoaeK1Fg3BCkMs9NnIOBnHEAgSQaBqK4pMHbcmo2pqC+rclLxITXLidL8PA
pV/ou3pVGb+mw57ytUupA9umIHAABVoA3JnTwSfnrfyUeGtShW6Fsl3iWOLQp1XF
KjXA/gZBkolWd/HK+/vvvWku1Eckt3u9VvVmj7wOqhbUA4Tb74EMATLpoqso0xE8
MMKXivs/vO3XHx1wZUPDRocya0hUKGR3l/GUba36ne3wQeOwrNv94FeXcngP/d2L
G1sHq8794ZtdicmlnLtjsmM9pP7Zvy/jAdBjgxH+YRhiJH12ix7LjX+LDGpQxx/K
7tA/DSaS265PR3FB77lMBk0Eq3+w23KAoqczC3qIDLlo895+6pnH8H8e6vHfZANh
5Xaw8fD4DzRvivCt8EksATFVvYIly2bUTzibMa/k4hIVFUHVYKTcN9Cg9gqBHgJu
Y2WYXb4HPM/ER+4HWE21pRCx9KA5pT1U03WBqCCBzAW3oxPSPDx528vxs6M0A+wJ
kHkWhgeaGVLnsrenmcEhysEX9vPW+/Guhneq93oQhPmz1c+EyqUo4pre8JXcr4G2
`protect END_PROTECTED
