`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zZC6bft1tPgXthTRz3Nv0llbd2Pa8fFh27rYXLzU7E9J/pq1hlWQSKZeFq+nSkqE
ecHPOGiFqht05toEZt4S8owlDuuuZh1Ul5OLdiXvUSP8+pALCcjOqMAFhMtb1AR3
38niexn/mK7OiX0SVzhu2/y3N15bsu2BiJN+v4JYsHvC+Zi5kTIN/ucoNF/jsH8G
MtBW1B+4TP3/Co312fMYzTM2F2ZKZqDFEN7EB094UTVKUE4J/BC7N/gkekAeEBiQ
Qb+Q/WfDZv2bUf9eCy7byYgKYaIlb7IvMneQlacvZoSNUoA8mbIHbwwEk0W5uAD3
5CPmPXCiJbibkpIcGpq1Q2291F4zEW/r1KvQDC9w5uRaIFghDRkq+9ueT4BKCngJ
QCx2m/+OQiXWreYC5XIgxRk3Dq9b0g1LxZ9v3J067ipKAVtN7wfUqZH18cWh9vOD
Y7+r4ISvOAeeaXNMbQsuVXLOK+aUOcqaLb+cZVi+Uk0irJ66lmTBBish0HwJzHN+
QS2ZsSufUBSEkNNDRvCRG2kTxjDi0PMVvlwz7QU1ea1g825julII77606aJbtLuN
K0y7/ozGN24zB4kSU2VoGgByjEc2zRlLt9Yet0htEbAxgul3Xaq3wXXTWSOhW45I
oYuhHQvrfGq6+u/dc+77QSG7vS9yKyAlq1URA7/kw3w8+CTmspKY2IGgub1831Wb
LBxha9Hqlf23sLoI4aCx8M5fupyTrpwiTJF+xKjiVH4LjY4lctv23J9ceFmjezPz
RUqKkfgAVMOIpOe9GWA0BOCMAGLU6Od2as1o3nyztpo0RBbfOUf5YW4xnQjYan5Q
OpXvt2kmVFEWo5Gi/vbMcWC/ZOqrHOuYWCN/UZTWY72kJucKVfE46JDHdbkbr7u1
x2eZXvdSMWwZEBBB13iV816e4EqwEWDzu0xIsqBqazJcIbg/YUpAZW6rF3hVBDX+
9hH5V1u0J0nEP/sHajGTCUven+g+5UWGylAqAuCBdRpclF7fAXuP6S5GzriH1Aa/
aAzEeWyfU2+2sg0m0vS/R5PyruH8wLpFFEATkGk2Y4kX9wGCFeEn6n/ychV3sJSS
8qVPlgqeQnyog1lbWHaGKCG90Ey65K9Qi6ZNuCdIm8Q6S9rSYetZw/EKjdtg2JoC
sjJmM2giMTgq6oaoWu6vOAwXt9Y1tbgPVQNnRDYYjDpFyAL+0ksK6FppL6QbX2le
wOx223J6siwHeW4bkkavzSa8aaF5P4Ec0aqdHukF9yb4KsVBGXsoj8InB7y1cvya
MOusUFezNMbWP91PnTO82zkhCes/D9ADybBytpH0PXMvYCr7Vv+tq3e3bwkmfS+J
vOt7w55XWpBtBhNO6NeGaBNww14njhlRWW0gR0uj/tLeyyRu7fKvaUxCW2PW80wy
5vTKvl833mnLc/jL6BfHdZe1PyDjwYLFzeP9Qqq/V3Bmak5pcG5NQ9+JQBtNpNPO
lmee4l0ebdbIAppmJ82AWENrdWvVeTKwYtGvHAxLMFBAc+55O5L2cb38shDpZc9j
l+wN0Ljd0LKf5Vta6L1rXbUZABDX1A5FEQKNJcSmgZIbxNzvpKxZhfqyf7/vSVvv
P9rWSI1A7vjAGDZqub4jgpGvzRy90sLhTfA4nY6U1OrIzSix8FM/oKWniMLf9zQl
3dCmUOfaQZCt86/xCsQPT6nmQFT3bSpbR1pp63eDvxvT8fqk7J2e/cPQYh/77rHK
oSmIATWT56gCNGiuqiI/AuF+SB8hvafmL+XxvgFDkPuYtTgA+y/Mor2DkOs8yoLN
NOgGAldRIy4Yba6HovsFkTVYhg82Hgfv5PE9rDGynDxQekmCTUSxIZBv/MTWaMka
t+jvdGoT5OPbfxtf/tTF/NIYI5Xi/HgPf3zexI3Cfxq5BL7HOsk88jDiydBaEqpi
IMNSSfpdmTDJe0HsCTA+ugo9+q6yweKWaifmmidsrboLr3/H/6qkQsHP3gNHHKWd
Kc1pyBsRaECiOCinlcgJDvZ8hn+IZOrrxbHXCNCOPjUOw5rPBwpG1uCnnI52L4Eu
BMZ8L/2bKBdrjEKdvByJ+uFuQ6aIvaWcNQsL3uVh2Y1ZmZ9krHVIC3V1HCpkVf2j
i0mcnNxbiW2VWLDc60LHkSiW1SzRm/hYU1GE7eezXfj8ZgYqlfZGkHdHP0wDn+T6
6rh2ChemyhkVJUX++jBAGxstrW4j9+grnDtDLJngHfITNr9a5xtJa1lsh+A/9NVF
7gkjlInQFHMdeMCrOKGoPe3heP9ouXT0z/MnIL3cAuBIEr9Mp+kolmCyGGrWZV6H
vuOUXo1Ik4RU/rEDukJqSP3uik/0bh2gnlyzIFsRCAFTJzyJ9lPGe1ZaPaRS8hL8
c9lHzAYsZmnZAiWg6WsSN0PfFLaZ+nfxUWnAA8hEGbtsWenUGhTi+wyhDGD2Fnlo
fxngFu/FlXoG8fYp6eMXJhcXCWTR32rerE6igH4TEiAqoZuQL2qXfOaeX/pTsPh/
QNA6tEqeNitm4XIu1jgTGBCr3D7FzmLKSu1O9ZOLZztuTW9Lz2D9wEQSbSG8nMjT
KEH3uN3jY3YA4oDl0JRUnVfV8eFztLCOx5uxth6fnp2BpKPVw0di5OjettJsPIuZ
CFN6rh4YzLxiJp3SuAi1ufPovY54OL1qScxa/x2AkxuCiVy94U8IGiXSF87vjta3
tWeBajuZ8bQ44hD1rW2opRJLkef5ICsr6/Q3uO7W8iH2vpwbYAXdBbq0p0d8hVE2
3OlIBIHLibNlR13jt/Oog9fWh18EWKYl+x1NyJjm9qw5yZqdg0iF/HkfukRzNVJH
N70zUJG3XQjBEzOZ4b7bqnUG6vfNUr0Y/NzrAxQoOerhzbGJDghQp9nK7sWzBrx9
hYNPDm7V17b2jrg5ahXBYphV6JWZDaSMZb05IPUAqc5OapCTQnSWZixwuZxgfzvU
2fAt14kgsLAQkTlknrDpBqvZKxURF3pOB06slXBg7COtJTEvGVbGvC0Ru2vTftZ3
02g5bg8eMOwfz0tdFnXRNrHwWkOLzWX+yD7mhmodqBLkI71pPfW7lVutW+SSds83
5mepvRe0rv/5WLr7oArp2ymkmJowpeXnJqowD/KC8/BQcGkDznjmCiFfCTxesMb8
S9dilexGL0keGTPGsWkCuZBcRIAeBYTgj6+rV+015NSYGE09nq+qn/+Ld0ejQDhS
FHsMk0D0wtUjtiCJPYSP+tew/92MNQ3sFWgYBGr+iOB2ADd3DWUzjqo3kfU2pO3l
hGS6aGcYqEXSRliB9ApH87qBUtYNWs/mIh2CFzbTDfmdjLGNxsqsms/lhSOnfL32
7R856H9tkIYiZ/ZdUp9AogKZ0pjhUs0mJnlqcNadDF43/jN+zxnm1TQlmQ2aMvOP
hq3h3aj4o3LUJ2ofodhPWCMt/0cYIco5PNqZ2E6Y58bwWeyyJshLrNrTcDT7v9Cj
p07/4TzerWNkU8G0K/kASEk+9QlwKqmq9iayohrX8oeycpljIHdWcE75WH6p1GsA
6INLp6NDQlmCYo8wi7zWT+oTxBG64Xh+U4QDUxTClzv6hIC9WMpDLP5DBf0hZLvQ
/MVc6ooGA02isCUixPDkuRjdTltCTts2py7RPBSOlup/ZRndbKzyq6/AwzbXt+9q
SlXRpfbssh32iBlhJCYcOUqJJWp1vQ2J6J3vzPnsNk7k8H50fOP3qhGB7/8L6QgC
pfgADPdWcG52tUxZ0w1YH02odGNf30LD76GWItu+gv+S9fJajqJbFOO3veCJQL69
Zm0zfJVF5wLXGOFoo337loRO6aJxIb/oalGyuMoIhvrkal+vx3YNrimVtTbqWzxQ
DeHqT3ELVKjpQh/vLzbWoCY19i8IVCeiEbBKb/lYqVCG2TIrPXWbExsB2CIoMyWV
p8urcWvo8rEEDdAAeTNPWFUJ3VleX5DHAPwnOGzEeD+KGX0N0zvzYj3Us2lcgHg8
Zo1M6Khouz4O2eyZN0obnPibZxQeAqYmD/gF45D8dZ0wnX+4dCQlwkZ0gHgHn4f9
Hrn4KcGMABa7zDL7f0X7AujryuYk+8CjF+502jKXR3A6Unl6G7S0hqZpEimK82rr
d+weI/atLlnO564CKhAuHnD13u/+8vv0Ruu8CrANdsysuo70o5MM0mThWlGxzmwj
gkAr/7MoaOXC+wQ9Vlf2LTbHBVIDzNx5JgD1Mzpr9llNDzznSQmperwlWuoDlIVp
A4Pr+rkKplr/fPMBzNeWhHluRbySoT0go4ysYjvEqjFiSoaz+418kKxqkhLQUXN6
ttMt96nqm3FvY7SmlMXhn9MzyiVk0e8UzKuXxITim8z+Pmf2Gxgl2gDFm8d3s8Tm
25bMOMr+8oUYFlZCXscGGSQsIxDkNQcCIczlfDqYMpLisA6yZ0Rfwi2TmuzjN0jc
DxkqhTS7lqmcfMfcooE+yCOQHILCVhXd+CaUHNqEaZXrtRCBZhz8KL32NklyhdTu
3ySy8+Pzl0n4MoKtw8M8qqiFllpRRS29Z25MKYq0My8qxWl9tzCQvtyi8r0UoKeb
DRJ2fA+xMYBp6MP0F8s5f4Lwp48t2AJK6F7sCG83B76fjVSHzzEG/PfM8EosR8L3
9OFDSQRuvljfGf3X13nTIg8V5hansf3sfJc8Gf9f4AA5rRZhhZGXDeNA9t3p83um
eVJ4Z0hjwwk1F+ACktWiksHkNfOz9XVbKGJsw3TghfSbS6B0p1zS2vzJyr/H8h1p
No6suFvFlxcGPC1nOpkAh8YDwWKk+X8SQVAlMuqbsXZ6qQUtyFVnDwPwNXREF32u
jPT7dD5B59zpUwv5GUrv0oI4BbtP644+8gEMA7dGXcsgsj+wBcMlfy67e3C6Nn0o
TaDN21cEEHudUsX2t8f6Vr7vu922OcXfVOXr/lfcKcRLD/MhZYKTPHu3kpSDAOYA
AVmbuBVOkd29kmJ8dCeKl6peuYFKkJkkTZiwHOHMY69c+O6OjXTYKw+/7Jyzj4q7
yc3RGepIlD2+2NGrUrAabaufSJf6rSD2qZQBRrVt6mbjwZvakzuv7at+MFie1ORo
PvmmImcFANeeus045RqzqrOlhn1yz9ixBbWaJX7ZFlokiAKfyvONhVwLcra+K8QP
HhR5B/iKguSchKMLxfzhlwAEHrmOP+7uvGxOy9fG6G2Qw8kqYegepBvI/GHlFC+o
2weijhSr6P4wLPADJlSx7srY85Pb8E6yKY41EfPnnVk6CmsvxUBYRk2IIYbm3CYP
Ac/KussBDF6JAu4DiD6BiyWXQzZANOvUpa3xEj+hpCHRHpXQbtGHqqk6iZf5V38M
yz5auG55ETpV40yvcLWBpTQSZfbvuWMKrxMS0KFfjj70DpHqtefaHMdzcJUsGeS6
qnFoVcwNHkjWqx0WJsfDw00F423F8EfOtHehOFKhrKaX2iICKx3BovnTrtJ77qjh
jat62bUVxiCnq5IZ/vxhREmk2L6C4Fgjq2WdLcUhYVZCeYstoDMdfwRNRgKm8Uhh
itwQUByQUYYsSH8wSgC0ek9WUnmslY0S4DuPhsD4+6RXobgMUB2Hn5rgQltG6wZm
Q4JJbZTsagNqeG5NT4KNuXiqnfklnxur6oQR7orDPn7od4C7EmGsNK4Z7RjJgEIV
rXW1sywRanLBWgMJ2D2L4TGg/QZi/Af59MIHQQfkZX81ek3kb0/Rz8AoOty0OhBp
S3V6Kq1wZGuOKXNif3L5czqJWXR2SKbUrQyficVm/JsOWqY7Ads7vQsCg3PpCTFa
5kyhyDpnspZ3MqOOghbwiD/kX5Q2uasM68Cwg4+xQN+UOpA0SfcIHN8v6fBhaRum
KNgSXYS1WsjKDUB74N6r6SNQAHWPAbxgQleDNSD97IhjAgaHXUfRbv6csVmKGBs3
1Tq+3kbBRIBXHRkXAAfI4sM/RWQg31m4EExfq1b6cBzfsH1ShU9GAuSRFSBbuoPQ
PC7fUhiwN28LpAImqsxSLgQNorfGFfCAAqsEvHlwE3vvKvmUGN5h9e6XDTsFtiSG
M2YHnEcJr3b9S10hqproZlPRcrn9lBWwQSbjFSm2TWryYf5sHrC+VC/AokYwO3Oj
1u/3z+g+OnItw52WOCyN1lkilUjSWNHZ2uFtehFKFwb/JmHr6S6G0/TyWExLljlX
vGzpR5SaoSUYUkEDRFvTrbQlmvBX+UDNU+aqMl6D+tJw2QhhjzlaEML5e4izM4kT
jWwB/PqBloWcfmj3xb2hcbVdpSSfRpfJz2+s6Z50XJWi4s5tqVldw8WmJhoglEcp
qb6SNv+hsXdnQWI3+n0q8uz/EVJy9jylqf/1lwJNHNKQZq0GaBwVaJTh/YVzX9Yx
9SJlaV5Hy500z1/ndE+hx+d1UTMeDP0d2yasrQ6kIIWtg8nkZKUrJHWLEZDQF780
FG1fNHWzwMsEhxj1KBvGmZshwCjRAoXPXsHbrrioxoK5O9dHEjYr3OqSsggPU/QS
4tVEXUUc7bl38pPfjYtPmSZjokcrb2dRNs4Dc8xq+mNCJfoC3+BZzq2pPKUeFn7j
p1QyevuqrJRkr8sqjnn19QGuRSUlsAaaLGrqqOp4CFLImvLrBFgwXSBUi+465g+t
V+Pc5072mp+WIlexU9Z9Zv0PzHdpa01YUVqjh3vx9L/NSCiciz7/0vpuO1eE/l0e
HbEqgDY7bJiG/pS9EiJLR1BzSFOzgYHraZxinWKTNblStr2CRStZOrdo1OGpmiw+
GJsTeIUBWI+g1yVXtYN2/CIW34WDbu/kxt9Pglq37Q+WvI5dk+yl07QUtfdubqT4
PpbEu4QDV0Od5c/tKBzI+gKLoNaQqQr3yDLerGEDZ7KX5DPNAYz0otwLi7y01Gw5
y6kBwVM4b+Aqz6YDgSoaQNuLnfee6Eryhp9z0MN/HIdrGOXxB6Fg2RJltKL+dAY3
Cy1Lh2xdLPbwvJn4FvSyAyLnuVJuBobFdT4Q/xEA3M0aAJ526Ef604msIC3+HeOj
gz28VYW7ffYMHNCHoql79lt8+IKGLfizzQkIDwft0zltAUvmSrjThmSRREp1ofZc
ATFJcF3QcTErlBYfdnyc9l5BdenHzo9X7kg+kjdk/kR5n98juyONCAWJSfjk4WfM
xZ3YvgxeLMb4fAD1wPQPBTZvFXPSHmPQfRsbJLKoFcyyR1tAdKkkT6nww3V58XDw
53UttiLPjBtlJ2rThsW98asizNGgzhKPF/cYVQI5i6VCwd8ZOR0DBgO4xN9TRMpi
2AfwYrbYUPNunQBgbsR0S/pz92nUwdxzbBxt26kA54D03sm03ETj+OjJuNFiDcfO
IuASKX7NemaPspT6XTWOVVZW1c1/ltShCsUWwHOAr1ewDeb8W3YYjD5KVUj4o2Kv
krw5H+r3xFEET10CS/g4XOVIfhLLCdbKqpfoUWk3Tjt0PVnmjwOV8IGT2ZheoRxA
gNBuZ3Va2h/UHg/KX7i3bUIhaDssKgUuzv4q+a0fq/Ri8ddx0EQq9j686Srl+oID
DH/Z1tw/e5CeOTLpwYQqkkwV1l/FXAj2XE3xIMdyidWbo1/fEBADO5FIvxkz57H5
DzuE3Bf75LT4c5+fJMMXaWurz96blkGWUa0saM9I+zLqiokaQuU+CzRzgho7zkKo
gvY6M0nQmCq8s7yMEPqj/a1N3mgCka/9z8iUHFM4FtBSQ/u2WWvPY2zWqMc8dlNe
svoKvsI/20SRBKE89Wt4eExQdw8n/dWBUxpzGksP0bm28OvVp9yDlqvKZzRCUVpX
mJP/UIth1DFUfYsufRk+T3PH2EO3lEi6LtOvbVCG7GaSB3AXsJC/MCujBXBheFiK
N/3HFhd0VtftJTpmPGW9FrScJ1vE4ovtZ5a5pZ78kI0MAp8jhV+w7+uDv4sgVOgx
cp0rp9m47EIFyjP94IGAeHBF/9SXnYsKlX8YkZspKnjziAxgxePx7juJ8rpM4yGh
FsgfDOTkckXWqAjEeUbt5CdXh8ms9A3eofjnOC+sPeWSmVl9znw+6z50uf1KUK3M
7ADS+KAVAcdT99F3qHpItxWi6vTW6Y2j744KLZubl6ptVL8b+NN2Im2WCNA4CdAE
lH5TA2uGS8KZePRfIRBQEfCdDlBXTbZBs3IHZaT5PRKpO1GO6vDO75djt3mlizzL
B++CTUJd2JjUWUlHI7HrpjGRM/iYJjGgenkQJT/ecUoo8H+bnbtx0gXrnM24VKqI
Oj31WSa2g0z5a4MbKVK0h7YSABhtE8jGRGh4BRZwSu3GOitr2dS5KIanT3PRJF+Q
2cjf0Fi3SbLgXii79rFsMHWD487hZpeZD10WLVfy3FHOhhlgfMVZVxmhluGDAMRs
1yjcnN9hgi7eTub4MYehXdQjM/TlAfay/5ZdX5DHxLj9MEh+XiBeKNAWNEH8sl+X
GlyK5QKLxHqW9zRXp3ZJLOO2BswpHr57eqA3YioZo1kdNdK1VOUvXOhL/0R7VaIO
0gZeNJQ1cK/xZ0yhsQ/HkZKVnr816tcyeWnOjuQJhAkF3PGFbbvfAv+VB9nWiPov
HusBx7zTa0zDfMPDurKviTM8JZjKZYe5R9qYO7zChRkPmMopmKAbckJz85epXurO
m6j12kzAmtDLd0WJCa/llm0Q0SnYiKWld5BwsY6qzAa988YDyInXx86XHmFwQv/7
8z+TiDoZgy6LuyrclsBnhFVPYxIeJNrWVwJX28jthnBG++0Dl/NKQdjgOZhTT1eo
pfRkmvVZEKCXjGC2muN+Qr6w/Nk8sz+fRSbEqSMQspRtCIOsDSD33rlYxXXEI2xV
GhJhcQZ7RDL8ETdLbzIN2uzvrlywwXlO+9LazwKuyPRdJSPGCIDJJZ4g+8RiDi1x
DdFqF0xIo/IuULg674XI4PAnnWdMlW0QrENmDueoKvIws+sWCwARZSyvlT5TPeAL
UvpOsVKD8z6vhWk7buNYvd+PPRZYD3K6cYCtslIgiIcNdI84fg6gOxk7Xl6S75ow
CnoIZPuzXeaHdabxG9cDwj6SypRK7fymaRXqZEpcHhhiuzkr+KXw4KhHR13vwauo
s9KcITeNnMAZgxY+8tu8CpK/RksIRPVqBeerkZHbQq5LHVwEcflGr0DJNiH/1pI6
JqcZF/hkSmmL9ecyOq4wFTS7oXTxx9w5TMRcaNy6FHVhJrov4EnxW795N6SDJ8Az
3p13MdAU9z/NWH9w+iJUeL2ozIz5mWNC9WgMqh4saO3PsYUMcZPQYRnkrr/usVg1
wEFMZu5WHwl6Qrcokq6ddTP0K6wplcHj7AY8/B8TgL+2EQ9KphiMA+5h2hn9u2MM
TXYlQ+whBSyv7fykfIoJzoVdqVVrAlYd8Ec9GbA7OzIZbbkJkypOLvKTt72jEgC5
bH56EwuK0EZyOwxmb3p37EjuHEEXxpFPY2wOup9XQ+AaqRSq+NKT26BYwMavAIOC
iusvRcPVRWQmJ+vCydUa9ZVUxISQPOod/SJ0Xw4ODhJcvXmdEgIvhxDf/X6Riqnw
hCsOsPcEsODpYGkEflQD5VM1Mulhl46R7u9ZW3dRKVEh8o7pWXEXzafsqQNZtGyu
EeJatcU3rgKiZVGzAI1dSbWWcd8RZBS2NW2+2qWoN/xFoqvzReQQ7EBvQNakss1c
31G6OnTAaCM7aeWBS5aGFtY/TlaDbpVVgdtM3OkZeaouPA1aQSHmZwUMeCl3E9ZK
wsPQ95mpwZDs7Q3npN5+YaOjng0xhMctPNIfBjc5TvtF3Ow/J/XTMVE65Vk7DrKx
BARmJLTt36ZniM6kgC1m3prbUrpmbTTfOrIzhr2aZJO6iVSygcPMk2QzKi1rRvw0
cnLaqmdvRksa6z/wSni3saAgV27XqyRTIVounJk+hS7ZF/wiFWdzZMZlMAxfn8Bl
aoNcoKqPbrCQoX1FObZuixvr/LP2ZBFDIw+2hGKjdXH3fa++4gkNXogoCCmGRorl
pKX2UuMsyG27jgG2lM0R9dv/u1/XxqevF9V7kksxyJV8BwAkcD5BW01SSEi6hYm6
S5AoSQcmFAv0il5T/P/jVz8N19ZZpqpZ/qiixxcefMWg8wi8Jhbe18xFz1m1LBEz
9T24hRUa7Wvo0aJJNbdAMdFIckJeUprAj/8nj8h1wqyWeYW+BclMRZl0OLQqK3UP
E0IBXMSzwIrvhGv8+HWVz7pTeIs7LcOkmF3wy82TyEw+MfHgO8PVvB7sWiB9E5Uz
gyO+k4XS1+yrgauXmpfWX55KWMV1jYnr/4Pd66Y0Gk3218NPZinDVtH3kGiTDLid
tGMs4jn0rk3NY/1LEEvY+PvD4Tc19Wb71UVhJyMsGmebYonAs7sbuDVNpIQGUtVp
DVE9u75OW2C/wXkuNrYooq7lzRblBLbNwtu/+1UpQLUV+KquJoq5Bax1J19mFpnL
WW40inmXT5jpv1a02Ziz0EP2vl9/he0ZcJjhMMi/KpBCdNFGSBGmES9YdMQZ/dR9
KqYFYsB1xXfdlpCUZQGWsOcFRB29NJrs5AxfQI5veMKRN2wx2JyLwqhpZMIg5//D
u6HNxHOwqcpvQNxpQLkPGPIl8rpVZKdGvj7/6a25/xrltOZvhA6qi1VuFkehTq3g
Db0njEnps4vw10Vj0gUE81ejnc9iSO2TCIvqi5vFXTWocyNs62Hh6eMjeUvMjOa8
okdH/nJVl+7E1JyYPfXQsYkasbW5MjvIm5SFKCT30GubmlzjJQz1xwe50J1U3cB8
cMeZgIxkjysdCDzeUbvvdAM52XbzvIY/v+3HPoLwqyYzNfFxfA4OaTqATkQdmiJk
KVLjSilN52KorS0wxLF9TcE8bx0TJZ4/2nZxJhoC4IerCPVtBtbRpMx7OL2VCE3A
opc5QZ4VrALwHMUoNBcN2SEv4wSGSHcg2vffhn0uBzuVg1xoqvRT9BY7rr5opBv8
R/ktQozNLxqIhnQCqPVtGVeT5NeGMV7ieMYVajnCViSzMT4ukM73ybsVN1YCz+Wo
YjXX1QlNQ2I4GWPxNgcW4zXLS3GK5gJMF3RazmQhX++K9bpHe3RnpBb4SMDQ/RbR
k+0MSLc+PaYH/7DX8ArYHeVzyFOVoUxwMD2y0TogjFduBdoZ/ibMCHG8TnwgMOcp
hcdbq35uXUpPXBvJPIu8zgc0FiCNUFySyRuSvGFma3NSxUXyjZSfytfvzjdnV65p
kRM27FfnAT+aBBp+xk/usdyGtc9fIZDtszyYFs/tMUQ/eu1OkTTv3MEsNOD9wvuc
hpoTS+JKe5RR1Y5Q3Ix1/yq4ThL71UBI7MCI3jm8gvuf3RGoJiYJtg8B3lLj5YOX
FaPNaNK71KTrKKymtdOi+oFE2AXRzYNit+e9rrqzRqOS0DCMB7ahTwkb3nOTPI4e
gZs30NOYrrSzP9hsZRHhFXXj8rOt3o0Ec8/C6nbrT34uI5KstL0jdf5W084WQUC+
QxxUNEo8iUvWRH6uC8ukyTwU+anCnLypv6NYjm4Ezi+s9nLw0KZuEa2QgxRPoxmw
MG33EtXfW0jpY8V92p8T57DVzSgHAI7gvCuWajW5xwiuhdDleltZpFiZzABbeast
TPS8gS+LTurVVhYGjifk/El4HRMFBWo50t2xU2SifSAX5gmBr3IDZcOrn+5s242m
OJMjasCj0kqCVg/NOlfxdM/WfC1vV6KqbV06J5D+5iVEHq6aYfN4htJHJiRTBH7J
euG3KPvyGhtTChr5pcI6QKF3AnFfBSzL7uLdKDE3Flmxx02I7mSXhdTkpTFFpISd
Waix4qCUpONr9qbZ/uTZ0JuetDyI6pNXCtYKgxKQsFuPFwcVLWTtFtHzjs7pV0TA
WUCdl6ojU9G1CDOChUQCximqI4FDdsIjvipRJoYi1by4teUMuZkxnr+Q3rzK3nMf
neWLLmcKBrSrIp/msvaY2AmjO1mSupBZ3ExZLRukbeBlwzmQrN29CBOSQvocF5C1
1HTcPHJot5FQaJ/+8hmyTkFAsFzke2SvEtwvF9IDU7Dw61t/z6/p0GEkv2FgFURs
QXa9xjsJh+cSNp4sMxaG0A06YLlMbHDdI/OGl6TGSSe8gh2xxKhCRTvWUgeraGHi
+5mwTLn7dzU5w1ATsTbOCV+Ebal5cUslNlX/Wf1TfYIFxBMNcZtzGE3UB0/S5IAe
i/zBsPp9ABgCF3oQ/V9teFPhS18eaTeA+b98IzkTBqd4Osmb9feE44EcpxZq/z/C
3a9Pz1FyJE40mVdYYZCuqmIcPWp/8q8B5C9rSpjcFUMy+/7jefwMGgKIlVRsA4NM
jVuE1pl2LWWtGMSqoNS67YeTU7FNy9JViTpIPMq73UhqtjTUR0E74S+AJfzLSZqB
tv3YzeEfH1UbOWb38K9lINQfRqpsg+rGj1dt5oWyUIjqtaYHrtbKU08NpSUJXnpG
DZp9lWffdFLnUn6QNkFf7/45AMPhSojCKVNPNJ0ZeNodrZlGq8Oxy59AhJokLEih
zUEQrR0YURDbZUJ6ZmXJLvW468xGaS4jLQHsnA7SY5S58KkM3KR+hjI9KImETcwM
W15fixEbUXeToX7toPEnJFVXnvAMLXcJoRls4g3jlnoBvcxj+4uaLpBgDeLHjp4R
U/pbaHvaKrVyFYxGINFqZsTSYIrGJiiH9sj2s9qDzLAHgpX+P+bqDWqODhZwOGW8
MkciYrAJ/VEsbIuv56kfmLSITgtFX6xFAAS7CTFelc99pR10l4FPY9gAjdf1cB/q
Uzn2p1I4s9qzT3e1h/FWmcEmrsPYLYLXqC/x8XhWFQq5aTxaOwr5fctOu8yU5Jce
8c00HjiVWJ1h6iRUxKyhuqrTR7yKHPfRX1dWvtur8cvWanI8mZwKbGoDXG4ZpeKV
r2ZyNkDDfsDhdahBxJEd6ketm1C9q65ivuqYn6AtWokfL8eUhWDP8Spp6dHdFX3a
taSu6cCSJbDXUlpwjoVNmVE7kr0T49YS56UEA087Q8lDolCeTWxLKAiZCzsP9tLG
S3ma1MG0oCdSms+QDaXpfy3XUe10SjU93ZJBqUwQF/r2c8NbFztX5rEimd3ci6tY
BRlqV9Ty9y+BHEX3XkpyDjWu+5xfqyfGXUmNBWXZedGI/t1WabJoLb2NK+z+psYK
eumkNA4AkP5DeJTu6ze1HlM++tmaQuj0xmj9jXi62NdtIwoeIO4E9gtys56RJb3y
HvSWXHObXkyNtwWlHfmq841IdUFlsikyC37mV/twrbZrxkGrzvFFLDyy/GEgMz8d
C1PsCJStHGa6eO/HDkI+VS3a8pPUnNkJgr+hX9bM48KReXrIGZH32MuB0ASGG72n
tXMmE0TozByB+wBe1P+4BrWhSABi6bGvw0eIt9OzYLtJikZcVBmWjuFhk5ftuzck
gAMiB0PXBqCXj/VdR8floyiunpl2EL6mGrnn1NWlwQOhFTfT1on3YIpssfhjxSs9
gTiL3J8r5BP8X5KodLUY7RuopW0PiJO0TvK0kyz3rHt/GAmhxWmu5oGWZ9F/mrc4
MnLrjRA96uYYWv0g30CiA0uDPQLPh/EiDU0i2rBLhi9q24C4MW+lUpiOAH0H7tii
GzYgxLkHzFqag/CwIM4YAqGLXP8LDU2I3uxZLPw/lrPT3VFRfK54N7rLtN/rCR7v
bCOf50Qi5337xEfDSb5Qmvfn08eEBslCfN5xUzwHdzBykCL400xUhC4rc8lhLpm3
foxRYRvsEBMlAM/n0ov/izhwW9kqCzSMt+9C16L5ZM8MjW0gTm4MmffjFX6s0JIH
I8BGsUy/+m8R7D1ZenHB4UipTT4LBKiw05Eerr6x3n65CIxraW52jBf/IOgnTj3o
2APWsDF2O2elj0nLAvPGQfEqS3w01hB0sJnCwyOUkKc/qVenGSYTUyp82xXHAtTN
kyAoJFqrKNJuNM8nOodgeR14pfwjycArDrtZFoaC3lIGf/kyR3sF/dbgo/SjsK3/
xBZNYwPa2eNf9fFqVzGQ9WP4crHpp+03eAb3r4CvXhAKsOu8oUQTMQ5SOSouDtbc
6U55jthhJCRkAL0p5aNAk//TfiUPk5DU/Y4cBnMm7JbmR9zzCPngzSMpRmuze8XQ
Fd03U9HN0fE0K/uroq2wjkfzwco2z1wy+l5AhoFz6dINgGT3B18XOkheTujYzBuf
DihLxXCFpKOPltNi3hv/CLH2XdugomCnFsiYeUNLNQcKur1ZVw2R+19PD6TwSDxH
GC0xIM8PTzczQL4k1ZFsYPPM65Dy3+hyrJ+MkVzqTrEOaueUrmatdUA+t4RPphxr
ZLuPcqqNFK1odUTkb0mmZZqI/BB+Gg1yeloErzxzGkAtP7rQtBiE0q1L/0mf0J7t
oNmd20wzCM780TyeGmiA0c7whARRRYiK6PhUdoZezhykls2ny0SugzWyc7gW4Sin
s5ouKaD6B5tPRKsPWrVXyFidCucbEQnVKh/rXqnysRCAJm+zBoIGBhCif6nir6KB
yDBH0pSAj8JF/qs/i9MQG7eCGpty5CukIEwcyYlUAK0S1TzeHlqpnXurVXX6q/WL
N5ss/6QevHqcIFkX9GrgsqWmhcx2RiJVwijxGeGjApI3mZRHNY78cVvo62wjlro9
KteRW9fr2IXzvL6qVNvMzehMAiEbC+KLJM/9FYC+sPFHckoSG7vjzorqQMBdP/9T
XIEvaC5RAFW9gcQ4fYF5fKzcBI0OnFIRCrauqoziT7kDc2FFDDuL0J6S/r8oDMyz
AP/sM7zqCPT4UDM6Bgm0LcvrT0FQoClGFnhglwpsJlESh462Uirj6IvMf/soVmUH
1bewhkYZW/gRGHV/XPTwbHxdKQvUydEQ6bvFNUDgFsmP8lhH9hpc5Att6NHz6aSV
phhwompWqk4uDS0dPXc/7P4EOEq3zr7pOo42bMxmSYA0QO4rLbxYumOFEvCo4x6k
y0j3sFBqpY+gup2rb6T4cagWAnBnE5CzIrJOvNWcEa8w99SdGRY+7mJcxFBeN2Fo
UtKTinOIic61G6RpKCr2JUJwydm6wUXUgvGa9k8ek87nXpPNP/TEwVh9QFnZCwQH
JKkKLkxO3nmLmfFF6o108n4C+TNaM608RrS3Mw/u+hH0bBZi36O+LLSWoPb97bmS
tEfrlotNKEeynNtzICR7p9oCWiHd5krEjaz1ZXZQ602kvtjjEi7TZeRcSO/pLZA9
TmjYl7b9vN8pJD4WQcI2coLgfuAiYElqmeCQy6nOLDqhCEI3t0L6pUGVhe6lLgG5
SIFAJd3rmkvN0rByycjlT2whJsLTDuCtBzQChI81a4tqZIq3HbKXwLxk9oLMGmrp
IaSnV/y+gsCLgQfsh0sdnoTIzsNwYIfMnhwhmMs7TvNRTNVof1aqGof12mdV0jpe
izwTtbXphYsJnQO9hbSD+IKLnAqYOeNXi1WloMcDmrPIjJsZzLOzBH0W4YK+QB66
wWjla/bEhnMJRZh/shB2F0yBRArPFCi3+zp2VaqIm6a+SBtv3GbestROXhrVHS68
WR9jtHK5DGjsnU918QrRGJZLqAY094EhITg5si4wOtR2tqG4rbjS/o/T4v54IOcv
3i1gdSbWiI4Ae3w/wMmly4+Xvu+OpeMCWVql8WM98BjU07KmRmbOBiNKHwlJkP+6
XMfl3y8m5tNU8rfpgiEhcYi2c09C1cm4Tcx1w9YsJj9SYb5IJfrzIgkFdxSySuzI
VGZx/lwkQ8m6KutvcnkscGtNNs6D+JYKRYlUnFosonPdfzE19NTJPuNDfnBfLfWP
IG5vOtradPiirEFbxFmiT+GgENP5v2hjEMfbsyuFWKU3p0PTpYiadAB4+YxHOXPH
ERfqyLgePChC1T7zDTSVubSiQhLDdNndFJJyzUAXPVzkJai9CoAr05Z9amD5DhEp
0wvXGgGMDXwqriIF6N1IADucYljfjHK7BptyO1vF56aynfgXBuUcKFwHzosyLDos
psm41gNnDR/cMgwFcemXLkDyUjT/vgG/k6dUrcuvZ6GWhpxm0Ok8/ZiWqR+W9jFp
+/wlhVcgx5ujyVgzlZYU/W2AQa7g9crqqQZ6tdfMG6ceVodI/5OApQZwho9M+SQJ
C2+wVsRIHjhq3Z15mLOvvdLahdSeQGRSv9ytKixlnmu5Tqmnb/4IGlur39DR4PvF
6iJDPg6lEKr2qnNTpQ3vRoA1t2dKGwBl/xwALZ1yepwebtpL9qebAjdiofsh0ccB
wn32OwaNuaT1hia2olceS3lCieY0avHBfRVfMvEFn1dCDnUZgTKy3c9FifiDcf7z
AvpxiT8qwGPLywSMwrAYom/oiZzWTQkc3gQj+FyPnIhlbzyyO24Y2Onfr3yPYhnt
duUfEXFeuRLZLnG2LETPN9aT8Gh1YlHCG3QP5zaj79dGU5Ht3c89o8qAIldjYOJO
5z+CsvekcCLdmSIhzLQiaK8epwhilXCayjJAz6EN2RZO+zOU1CEGzWxbXaJM4kX7
/e3kJsPh8/Xom+pQ2p3LgAikiNL9KQj4FXajlXheYLR081XYmzdPOnxSnj3nrDHI
vwSFzbyWONOTJz/j6S7lA8CUgY32RdCMioJvrkBSDjteJDRFM8lFsvcx532z3iCN
/e21vsXVLNBrindsZoRzbo1MItAQnqxvsMq9RSgzm9yoiQha3iBZlGmkhE5nFWrn
lPsG2eYtZGLRAK9CnAlUTtaKjG+j8fQMhCYm5Qk71Ogty6lXgzgHE/wZPpd4w/AN
9n/bbQyoddFfm2OqCtOkr9ZkmAWSkurbZ7kj72ov1k/6KIjlPLOa5MBGx4GQjXd8
dXVKQrY7iJJ3b88HdBlXMcMQfCMjqM6nImk2x/xLiK3C/WOX+1IpzyylQYPZU7pf
kNlrwmb6MwhZg4WmoBcN4Q5maYMh502xajdGQs87vZkHVEGQfBbkn4xi2x2d9CmR
poaq1TKwqqIBEiUX6/c/EZiOdBbMZxe1itmn71nLB9fYHrDKyrYPoS42+F6wAMQH
rWyoM2xepB7OBCJb2fac3fvTwcyqX8H8CTz9p3KUvrebDOoPV1AFdItPKKWxjtqb
KjFh5NVFJ+sK/7+XQwnc1DgbLsZ4acJh3TlvxMHVIuwmpTXSBzqcsYgb02maJ3ds
Nz5jY79IWJEVbYiJd04npAGL6tw9dhjXSebqgj2d3VJom/99QpdHvCOEyEJ+I3pp
waBQ3IK7YrpPWSZcMQgRNX55t27oorNYeMH/z5FfJPexO8kZdp3GR43NtcHI9h6n
l2Nr7/qAuHQDD67AG0ndVn1ED5CEq/cLUsofztjv0eghn8AXwzUXNeLZTRFhE1ss
AK9cSJLvSWkCmbxGE1+J/bSbw3ccM6wak4gZ/F6wvMUN38ee7jFaNl97F4veLqop
gqKPWF5Lxom0IPyf/h8NnpkyN+s2EEJ8GoNarfOMDm+Gyf8STsGiXEAOdUMhOi1j
9f/XaeQDBSzFWDJ5X5AkIaJPmAUFCeOsQIgJMBtzqgOQbSDPwJvLShbfLsgdUjoa
KduwOzn+ueeWhKgidmKBZ+Xtd9M3g4nj+SY3YSyU5bnOFXbYNgLTYOpxvLUDgR4f
NGwjpYQsQM1vuxzEYMSXBRaN6Tm/GpEdQsP8nGOk5oYxQ2TCtfOnU9EC1gjmPG5I
d3ndQ5vCUBNjMaBLH+6BBzu01fGamIibZ0P1Srsj4U0GawBUcAFbAKC1CEE/0EAn
psx9AZTUqSfJjO9PRQLbsS3mF3Xqjw4lLDV7SgUVoOsUI8SVWOxggkWAuyM8Xe5i
0dtNny+wkWm9o1HuhqfKlH7bRU/gbLZtbv6CxayE9AVvSA2GX4xFdBlOWKNzLLwA
HSJF6Bt4409VvsKWzQsvfkRkAhmtu43915dHvZHJvY8d9Z0YTn4H/dub1aFMcVQ3
rdL4QDInBfSSzY/Wya34OVBnzrouoruBt6N/9iNZpCnDtZAFTby6sPGw9kto2w/F
WACMTUHYPlNhRFeI+8VC8DX0/WpjzIPjmfEkRDLFZgRi9hp+ayWJ0knsga6urm1Y
fSlvJPBYh8v1rJdyT4I6hE9pOjgYv9DkIsxoEK3CwWTLHqH+JOHKhQUkAjAS7nms
4YFU3RQkb4Ee8WGTVQlZ8Fe18EIEazku27cZhnUbP6Bhng1Z90tuFUei/NVZxhVf
3ay4Eiaqn3Cdv4Vtqx1hz8de8+xi5hlncE1XLmIxd+p5zYWOF0Phqm9e2ymYt9aG
sqkzqP/dKEA0Wvpks5xgiJF2v1/8gicuqb0DQXCoBI/iWqiG7LEJ8wxCz8W0YSMn
M3GqQTvpplqS829oK+LrqgIprdp+RBEBCx7kVzx+a5q8QNPXhJNvWuacGI38ONw9
k30Ich6h7sxLmmnCBKjcWdVenjQTYd4o4kO3Mrevm+4dxoYdEG1V1ozjNjWAoTEk
w2ouQ6nwC4odDL5u9ybb4+Dm6oF+KKwvrk4cRIs0kKsPdyNSa9ev1tNi13AQ6vTe
0NthPmyqTfqQXE/OkrVNdfP2nw/0dw/B4sgBXiRetsGN+hdZokosFaoCTtdxoO6y
wN8aUHxrMojwddxdLEkbNkCJar9guAKo6sH2MvVQw8P8R2FuwHDHeY2HIOz1YUof
u2lri7PLvmm92xsV2Zb+8kpsbdenv9j3sVJ4sE8GnsQ0Wl+SzncGgp0JrQd1zGLk
W10VvY7nOlBehss8ozZ/L50+8pNPXlQbDznxZsSgNZF6ISZABBCx3Fr7FnwaU2UX
krLMsJ0Nc3kGIdfBBWgamQETpNOxXajA3fmgF0TSZCjgiuI8topyRjCwF/Y/kAok
HMJ9efsi60NUVZEsbDH6nqVpx8IkYs9gDxOytIXEykmqUHJYt/TIg2TJ4nLEzzKA
BcSNYSb4UabujXEEdrZH0016SoNUGEW/9ocEKIeIMlGCEPGvX4GRacHTSqgtSnuV
bpgnNDTIkIneAWeV28Ya8R9ocTo4I64PwbDuC0/CWaUaui7mZ+EVzTHwqnDCz5lO
CD9ZgqCVZTDxaVNbpDpesZJbI64v9OZ7tAqteKVscM3EjnG9x3+LV5uhzfcY0NsV
IQncUXfSdYKIceFaEPANo98CoTGZ/tbAERNATTnk8yozbuvbreA1U90k5I79a0nx
+qWSYhq5V+x3ntFaLxm+TYWz0d8JRrRT6Ff6MVgu3CBuBdC2YN+Ypo0zhzhRfjiA
0jTjH9UaqEbC5P1LcHlMmMTedOplnuChln8dLsSCDTto4IcCm4ly43mIPD30LgWo
JWED8t2Cqtum4JEPB10hKqzZr8ap8vtmO+IMTGSTt1I3NYmc4mFz7qPEDR0rkjbX
qQcgnOHi55v7Z6uG4fWQfmSKgiu7quiewKLPNcPNdeBv3RN7QK8of7Lp8RXSY8vf
U/WcikE7AgEx0ToY/f3pg0OyZvtIgWptlsLqUzJ5O4nIcUMSRaYGTlbLkEKZRcAH
gn5gQ666zeAsuCtTur9qDWwV+z53n799s+GQ9UI9ijO1UcoPDCPNr68+OsQHqvyZ
SpL+8i5o4SkrTzX8QB7RbNpFqEWNCpYN0frCJiND0YsA1GALwwajjWQRiodPVYzk
bOFCJeDBBxfJwD7Qhx9vmn4BYinlTHWx/9aLltUC6eDDr7tKOxyYUKPyIm9KEwvd
mgepWfpGKqbxM5wZwhkkcRaUj1LNFKeDMYQEzGOw0s/xdFEXxobS3FbSJjxgDinS
cYdDE3RyVLxfuCl03UimRuvzXgfax6Nm2QfjsZBNiyZMmXMnCj6XYyB1PqpR8TJi
i4sPJdJmyz+Wb3N15thKoa6wwEPUj2Ba391LIc597z9CAPwfLNspNLWMaK1Zi/pn
vCXUtFZyrdRWslSd+qTf+GMhESt11QMNnmKvzG6ogRhx80fPucIlyKMBn5NqPpYR
hWJMMI09zUeh+X1tMGDx497oyRXZMdHHhq+aEFFk5w7bPGTvqmuobT81n4JzRIUt
MDqnHWy8/JpsMtJk4gnIV2LhShx8FEIM/Y0T4sa+u7Kg5XoKLyepzXL048qfYhdN
63/vYNNOlQ1eapF+1eAV2RjHi5ADt61Llrzo2aY7MnOUWEFRgE3sHn9VuCiDSFIs
Zntz1ITb6DBYpw7CnIKiMNZAPdaby8pJxGZoOEEU17w/+qHDHyjXJHr1iRjFkxmO
kOUS5nt5q5N2vrIBJs8mVyasMg5wNe2AFLSZ/6BgORbtG9Q8VG06a9PHs9h4YnRs
arvPfW9cu/+ovgMvXWe+CjWRjdLgWP/g97uHMMnZ5yh7L6GR4DBjfrstTME/+YAp
lcblrCbXyaWz6pluFi6UjisJNXG6zD0yHaagcEhyLtI+dApi0fURigNjvauZ8GHP
bOpSXoRXD6GU0rUXmZ3siYCYDT4/Z8V8P6S3bCnuOZgBvUz7oJ+0hWpF8EWqN/i0
nxB2Mlfg9VUNjJlVBRyf57IRHE1NR8DUxpYwk91G1CXwdnEK1Tv9lcgM3AX5oriu
j/4F7PiM9Tc4hL7TafsTUNpbmWY2R3dBS8CjKKONnYYSdx+sIiq/ZqlheTNd3CRz
5nvb079T2e2glojZLxWClp3uRw2iBLS6aXaEy0GEZfuEa8N/H0bnbUloHugTcl78
rclVFIxYfCl09TpglE7GRG1PjdeABTnPZAweEE9J72gHr7dWA6FR4Y8QhtVADMYM
vdi4cBmgT9e6olHGXC8F9Y8IbCqUaEejNLSFQOAXe7yGWG1fa/7un/YR/myOWxwd
NMW6UD2+2P/kpiSuACjLI506WjwMmfkZLGdBGuG4lNXnmhpB/8WAuL/drEw3nfCU
K7D7EOra1xX+XQ7WhrgoDdwMUJ+4G8tNFyZ7XAycpNIWeUdfiJDnubpPJDPA0aNr
BIAkAIqD7SSPB8C9DqVVGAAu+Zj1TcYWATyMi4Y7THi9I+tWGM9daj1kdn8Kn60N
sEfN5R799z5aG1ZbF1UZc115oe164U9ysZ3O6e8dlbCntyLyV2sPfYGWHZYsCg54
vqo6wPlQASb1cYjZLwj7tnxOQAtvVicfZ4sfDqGudngCERHLbUElGKVaAuFRM5nu
sD5Y9ZKFODfxOBxo66KdDKSqdsRVtnHq7Bv0brqUsDzfyFS52Lm3vfY9RvIvPZlF
qPZK1+K6tvDmU6/NYXXNRI7yV5/PtdmHXpoI2fNl8RRVF4vIYSrcbRKc9lI1GE7M
h9dwMYaGmdpvePpwe6NF2OlhOE438eO0x42ZTG8KAl52HPl299MmtNj0IAC/SKPt
moJdMztR1DsXMN7Sh1u+rMZ/hPuMkZcTdm7C847lBOHzToMJSMDoF6uWdwTdve0F
cVCu8aSOtWhy/5KpfK3mWdxJ5qLYwzjr8IoxQq5Ttza0HQdHFBfnA0EsEJP9G61c
nVBNzI/uNbrTjWijyMi/NazSKto1mWIkSfJslgjM1id4aEghmOv4QTtJyFaSEHTQ
wtGXxyRLToMWT1HZKbXEOSyzAS5BgHDH/hqydiYLgu8JSAxjrzNWoR26rq1xh38n
RfIabVgiK+mNmYjfvECJRO5ZpMIkWEnS6JUoDOIT66uZNthG2t7+5s4DLgx/LZrg
nSJHySvlC27JFIYqgvvUG6fZZnPMR98N/wni+nY9fC61xN/3Mgk067gKYET9ZMZd
oDrvmPzVroRJnSDqmxvgtoiUq5C8hBjBOXdIXzTMsaUUcKKQA7pCcEiBrDKLe9rR
ZF94PkvjZXaKd0wMZMyz1Os7O/a2SxiC6Gr1lZb4gohOZLJOfEYfWYZp1rt4UXQK
0yVc1hmQVrtN/I6tfnwxW493xcZa2n9lM7vsl1+KvjGr486j+/DfTu+50PUCv5yS
2oENCgJY5lvnFsvcE3fZi/LPyxa8eqsm085TtoHN8mcN5c2zrKPzIDmdrphEHJDO
XcMH27TPhK0deUIXRN7PihEd7MYbhly8oDIJogjuO+gjG5t17CwwWYcLSs+Hd9Mb
0Jv0Sfr1AWdsfAuioKz6EGPQpkd6Se2takV/ExYvnHXmsZT2HvtjepkMngEcQazm
iO94yNUpuyTFgnB0SHI5cQ9NNegVvYgSK2fEu2G+XdDIXrF1VRsBMykFARRLTMZq
OBD5S4I7ZFQHXv6Mcqya1xOJ3UURy3MgbsMxwrn4IF8VgM5CPe3j7zDCoa8P58FR
zFhVbS7RQ+L5mFzWbBEJuZ6ox6RQXfTWKbaaPopXnMzXgWg1pLmR5fgJVgwMvRM2
F/csym7bYKf6qQTFztGRbE9j95cVEdq81iCU50CYs1U9aEj/Z7ZXXFJnh6xziIj7
4+ARKfbzh5fL2OWn5PiJiNIutfscKlgWRVp9lIfEi2WOTxweBUxOrfjD3sN1kY0Q
YTVLmsc6Pn4K4c+3xTL46QPlNAwAtow20xH/3KO3trm0KbC4RmOOkBDnCAiFZq7r
tDd50x/ZzzXgIvfe7itQ860hqkTUjM5soW+pePz9lJ6AxkURBN5ceJS5LW4VlrKr
anoFC4rAd8hqlCXO1dn0fk48DTrYMa0X1EuObNcNGxKOr8sWSb4LJQ1TmDNf3Mz3
spb8blwuzRhCwhvosdVAUKV+SQw+VOzpISTKZp+sAiSOy7wilf5jhpflZCIHAkkl
gA5D49yR1dNbzWgiHd9/U7h/ZGHvsjMhPDMztqz1D+/dDEgWIJd828TDZw3XNv5W
dQ5TVwmICg0jSg1YovbdVm9SJjtMdFNghJHpW5Ucv7sp2i6GU/IM18Ai8TejLXoH
evD6sLgDT90qIYjj+RfohF127X29GDQZrNc1r/Nq8iEY2/fDJjbD809QY8hmD62T
vBQeJY1KHC9Tgy1WvniFGA9PA5H1nDNAnOU9N490/oKgHOkfB+O0GDYb/ucLSIt4
qQLX9nHq6i5oh6Ez7N2w4RtQmPFW3eqJsVW7xJFanUzxeAKknCPqq5tF4WBikcVd
VjHZz1eNboBp83/ZRZZXNd+9osaBBBDyhLtrHPhlqw+oc2DpT59hKo3fwX9oVVJc
2TEEgWFd0EpieWZDujNRxn32ZtqwXEnBJ126++ixCBxQtG/+jYrwIMkEUbBTSh4K
OzAm6aVu/1cC+Ivf+4zTczIMbuJF2E42209boMfBNaHRHCfufk84g2m1pUZpukEU
2WodWt04VY4pPUVcqRssPW6u95sdcqchJFA7wCA7t34ZDaHipaAyJJmhmsP9H00N
67McpfHO4phLll0PU9cc8rtRQQwDqvI/9RaBlFsv2PKXFV02v2isaIHqC15/QnaU
MvI6q3U3UQgNrBXb8BV9oMACnzV+XJk6fE5ziZg/k6WPC58Mq734mmoUW35FH6VM
/Ni2wOw/Wqzqz+C6EmuymoNoEUGzpxUanNxWDkDeQyqM+J6IFY647b2S78/88w7m
2h3oRVKTX3iydfjBBYSzsDKvfgZ/7iw28P+2gcJDwogIQupUUiiBwoRBIcRIaZ0H
ZJGGE5QHIecKp9KmZDKWBMXmuQQ4jh+M69nqvtN7s0qv+ynXYd6c7vIpp0bC63v0
prZPqwwpqu9B/bw0OFUfYeKasZ1jgcf10SPNGy8VXiFxsaenvJ1MhUNNfA2sus5z
bih97sV3v2y4eJH1e0KlgLDeScZ5MXlC2SmXJMYqyFx+ue2B/zyI7XiJ38rjC+Pj
dTn+3bdOcXC76UIrJSJBKLnf091HtgOHamMMUAbb+Cr3Bz9aKxbMzOwRWThKvyKE
0lMX8aX7N2UBtvaOvRJPsVbLEhukxvkNV/qevHJukKoKmYgfnNT98Mefe5mkGMVu
/o1wZl6h5rTbDuo7PhMrTHxTt4eTD+d4c8/j1p/jGlc40F3+SOoDL/Ba17BVuCIm
69YLuhSAZyYLzWVj+G9FGtVWUE7DeukH7iQRlfnEqbJZX4ZHlBgI+2PN2VeoXAwr
os8+uTvtrvVai3L0v318+0lTcIHO2v78wT2wKP7qH82mVzrG0FT86RJ6T/FIMqjc
+On67LLRH/oKuFBXTX8MKzQr95Rj+1YE0TZqTRCkIiFI1TyRuWpTwykGULUuVOs3
EWGaL/7/QmM5Hpxmx8BFzudsq1T3vmKgpNr1TkAIFORJhMzUJjasyCGww4uzRpiY
fUylIhd9ookU90yD9xs69uMh+3GpxrU7HO962bsmCrQ7RYMleLYH+RqXbh3vr0iY
J/6i1CEGzpZfYMYu9a2CchbZw5Oh0+LMWt11cDv619gAs16dI6gJjjd1IszhFRHI
xyD0S+3zeaxZSVi8ePnXyGAqG19TLfteu1d11uxrAkjSJ+Kf7CJ3pqYVZV+qtmKj
/A05IdXRhq0AMuZSNVyB2sx5izo7DQ12hd/xlI/z8Tz9ArZxcZeIP47XtI2BZCBM
sIz4ePGrrNy4PiC6lQdpCZauB5qjlUd4MG4YoPQT3NUWCitn3mo4aHL/MdM/v0A5
THq4m0vlx9JgGV1aXgnwTmBHkC+1FSuDAlwkdRB6adQoRnNY5rDQEbj/x8B4Yb1Y
Ah3SLySBO9HJk9QC7l/nJLhNm80EHRy/GegYyzCg2PzawYfEZt4MYO25wOxaW0AK
eVcm/RWodP6a9AOWe9kLaPgJr4E0Omwl+Oed27S+EBvoheIsMMNZXWgzB4WqqDxe
u4QzdlFk/BREDAGlwHP0yJ+pdzW1bT1pUfHwN4ewqa4GK3DTmk/XnmirekSnETNw
IPhaMnQHyq7+YSmeOFB9iTfHLjQJ4zrOkj41MmB+1NPERU69baOufw29KA1chkjs
0nESOLKw2tMIClvO6OKUKZ6YLky6KKRFaTEke8g/6YiecqEgHu/Vnl1oRAgccEou
g+R1IWJW4oJMEBnYDvFg6RIcDwDT/akTFs2IpOokzFqw1KR7pKyvNvJnyg56sC6M
maWYrexkaCbvXw4MaIUyHlT6M1QqOXQ/4v6kCbT9j49et54dV2hgIt2RL9SVWxY2
vGscepD1QdOuLgSrO6KycgNsYRSrz1Wy8ZFmIaxp7dCeDuYfBYQUGpiDg1NwSjgq
bIMlDUoUn42NU8WsnfRFcoB0NAzNWHPTY5HJXMOxb/ro5NssPLLwLosQwHjlEB6E
6AX320qsMg2pLooa8pTFi8XmLzNNwxpxe4Z9ESEk9bn+AH+UpVnqZtg2OMRZciLM
jkwFBQmxZe/9qtUhV/kGO756zvbn12kPFYmux98QifvhnwmeDpQpwdpxWlPX9dzC
j265NEXaq4ohAY+s6mYgZRvAUxOjIGagBOg4WeaKoBvI7/OBEPhfktNz14EF6xdd
MMqPJJDUnpbWI92zpcZqEAObwf4aSDF336Q8XqcWtko9wlk0gYr4fT6BeTGJ6GJx
zETMZ7seE1dXaulTmu2eSHQV/weA+Zax3Ht5J03JnSEMXvLd65YLIY/0RPDLPYEJ
V4CArS5rcWDFslyUZrtMZi2sPz9yMR15ny1ykayhXzXHd3xQXl1eCB9xlV8r4lEb
mWGJ1vRyfd6Jzn1D1QuISgzQqvmKpvH2DOWebI/8iNffGLg2J32sLnZKm/0edMHW
y4TFpOhabn/rTT1WlBdnI9G1qnc1nVOm6Sa4wkuEiQoLyTZyWLIThy0rk72x/o1Z
k9G3cXJwQM2KgJb8ZdKSJUJHF2WaR+GqtLEDaK5jtXb2JBmEYyksXdjYUvFAZNTK
qWeCkgzW007Oq6xVQE1RFsLnWvky+ygwVDeTr3kJSkBOKC732B/yOoSlr+7HRKsu
P6CFnuhisw4tQTVHBHh5kbcmxSKJIGY1jDNQYrf1gCigwmC10QY8vU/QFT1o99z5
Elry7g+Ft+d5WTp+Cn5LzFjZdZByWht5Y+ffTpoEySGcx3n+yZQDKCn7+CWAJfad
Br9XfzXSeJGxw1bhl885q/ARFWi3w/V/tx7Db8zJOfyeaobUHDmA0EpDLNe6p5Sf
Pv0MkiHnn51o4wwQ2wdsl0fQVnIZMKQnLasuhF5Pv/V01yrrEPJl+dieai4k/vD+
zcsJcO7J7qtuO37QnUV3rA+HXmLjK+hrY2pL94g3wPOmRgrUqK1NtQ84QZmJJdns
ifEgnnUgkbnHhqxbn0G/qioj3957Fjqap1WrxSJnyYDuHfXfNMQLJ2gMy+9WutBf
O1koUQQRMXMqK+zU9DerBjgJANSMyw4yjkXfdOLqQK/R/vvLR9oJErAv1ki7b0Ca
DhDxqTv6/48SiZCMG3Qv4HfsfnMDiFVFLkS3ixOCGQTdQbOPyBZUJIxoprOpOYQK
iDUlgyF9JrJ2qKDyYJi55C8fwnmd/nBr57LRjAW75HC+9Lbt/2mjHRmiD12t/WBX
gxMaiukllvPO0QlBcwnS8qWxqyRvk93mgEQwTSt45qlCyrB8o/Ks2N1FSroPsD3d
xYEK9jqaKe0G8ObPuT9omrgktSxlFyyvj3CFohJXIp38jQ57rVJz/g0V2ZfJLaJe
9sxgv+9kVqa4N9cAD2lck52A0eknOH88KXhnKWVIT3kL8f8nRHo5XhOvZjVtO7Xy
CAjK1xzcBKzR9ejyrLMbGWCq7M85iKw0wlPkXKOxkTq2z8K5nxpzpjVgFhp4wIwr
+s/uINLXbhwTvG0w1e9NJ+6oBMNkI2P8ljBWsv7OXtabk3V58pH80x5tZGulSQY2
/4bPi3rHsAdvP06En0fhvGLJunATFw1wJY3yT7VN20s+l4+9pVfgg5JX0szVaHEt
b23klvNSSe/+2IeZHu3OhsfMqtCuS33Poun80HGeXbfBjORdLZzdeV2MItXwlTnf
Pu7AXRJTIoVJDr+lwNoj9bEw9D3NzAtph3NxWkSZgos4e280kB751pJBDa3ExniI
G86mTPgUG9xBYHetSyZKw/CcZBqkh7v+ttq5horMoupmnmKjev18ccoF5qiofau/
sxHp+bbtRlug3ty098j5O+zJRG4w084jPUL/ILGisGezPL6bser0qY87f2P+SPuJ
WSc+OhWDXpFSgE/k0s0pX/5PqywQQIu3pQ32KQ3QuQ4HaUq6CG93cE46n7+se179
wAN54iSl+yIhhxoVFV2KdhkVbXoWbJg9lItgMKfBdJpxjfqK8B9bmcKC2ZZjefYB
6smj6ri5mqsf18QLwAgTT12PlRBMKn3oGHS0eNfkXcgFIIDBw9FBc47XDWaPbZUG
MuByDBzmyUcypfUkL8y7YiNOxfiIgKH7P80WxAz8+XM68Znk2a1BLCq3ogr0Yr55
8yxUBQyFr1TQpH6EE6nyKnSSCAuczY0ViueXnMUVhYnjSS4SX6g6km5fjsHVeTrw
Ik6uG0Od8Ymr1o0sdXBTKgK88fProLX9TLYuhOXPWLj5R0ejdWKV86+zcQvYoIKN
7SNoRKGHhMraoJpukPcb5jYGem6wONLAqt02NgxbRH5AonpNZdDDiuuW8tzG+X6k
TDhTZvVJaG2DMAU1/PetGIqZGTVNJ6ZpDP5776CnL4V5/7nai05zLTPODX+uIaQA
IA9W+o6j7L3sqkCIOdBU+01yLls7GKwy18QTu8BAbHsRsd2X5xh2Naf2/ly5Q3zd
ECAtkW8slup7IWQ81GTSUFPy+IRf/GNPIj7IGsiqxAQZpjQY+1am7gmtpK20CbYz
XOsuIAGXWqF2RGxt0ZqdPvOMppOdlWWMDXAgep16mpYOHiv14dyjbg88e1T/pK77
xYSlRWSpmNgtxxJdv2oZH+5/iD32D8Kjy5b4CmxuUkcRBVSwuowzX+Jj/T4JkyvO
2EhjEBF97FdIih2A0i6e9Drb+woDU48L19zx0gAb1bTwMhl8PAgCsLdHtUsG+ZwU
rb29I1ImxCR7HRv2eb6S3eikEb3kbykPIli+Rn/A8zP9m7qmbL9GNwGxl1RUj9C6
f09JhMXxB08rxR3MH3MPovUJ0p8oEMbgWsF/FK2G/0J6uH9SDqcMmfgF76DMK+IP
rBVj5v7orkOcT61cTtNzo2tQpxMA2R3cgJUD3YJGsOKVDThby493JfEF+0yG5mOj
sbMHbLOQHhMxUjfGfwoeYUGGfUqGh7y5Fat5aoMfKYYHzXf+Dlzi4gndbIAUHniN
vbRVE4lOu/FjCHEvXNYvV4PqckQBZFP/Yd5KWRkgutpztnQM6zZp7vrJWqErSA/n
25ycLy58JIz6ORCIN3kuXzFQEa4CtHd5oueluiNCS1L/x8PgZ+kN0Zeln4tRUhoG
But7tIf8kujcbllXkXRpZtEzcfjVsZBgkuTyHfXs/trBP+Pp6hyrEc/J3n7x+WgQ
Q78VUncK5Z2T8o3QXzQsklegYmKCMFNBJS5bj1OnEOnpF6Z12LLnTq36/dICpt/3
l53cFBSfXVoiV5yt753d6S4DpzFWbiCHSwHdIJHLnyvn5f/x7Bj8bn/XTuv7dO5P
Nt/Lbm9uxOK9ZC/hJurQ20wnyq9eJpiikFXtQ0vdTTn9bVqjbXV1s0yZyGpKoNLg
WyfpINnZhk+zgPIW6RiQHD48tn6Ay4fVf2aXgTb4PmmVj0qvzQ8LO+9K7Tsp8Rm2
oMUppbHKlbGPJcIT0benOCss9WfSAVcpE0aH55FCHvTC2af4ImQRBXDNzkSjluCJ
XtlMSGl35iqkzLsmLnMz1PlYU7+kAFs7bcNw7G314Vzc4SaGMLeR3JKNp7tMRgHU
ZbhvwZFmJEUy6glejsLvYcp90ArYQt5as24T079bHMB5uMXpNBXI8ldrDP8RwVN6
di0Qh77RfAwyIYFtL+ZfUJXW6Vu7vOgOBv2k24MZJmcNEXY1nDgB1frGLx1GEJdy
ee+jZ/GLJFGhonn+hS8DeLOeWFme35eD+pD1pfhFPDH63fQttYqayQBPEL9yzKD4
jJkagy55Ab1sDHMHXexLl2XHt2mAttlVEx18AYLflUSCTcd/Q4ndL7XQLc7iSnbE
tEUkg250VCgW/SASYpDX48MzNU/f+zE8TBNEjTqZB5Q4/X5Cl5O9X5kWk43fY31J
RmxhhDDNmGmGtLIXXizA3NUk7z8CRMbMl3BvNu1kAR5btJAV2StfTJQhtf6i2I2f
7spxen5zMLt0F39jp/3xiRx1yQfCKkpy44IaQIfCadZzBjr+jFiX/yla+4Yr//X0
Cc5tXNHJrSrRi40KcEljhXD5vC1o08Hp9fgVqZXsqb9psnqerEhITnzXHtM0csl6
maRjw+85iDIeKgvbvGUe19xKkYXMKCdkXyzrA/CEdE2yPGPBE4GAh9rXdRb23+2z
jyd8UkHADTpXd7+nQCgvuQpuA5hkQAOv65elL+6O5qUyOnBP1vmWg+bKzMA52l/N
Gs2rjYC7LleqlX8KnxN0qipGrtBaXjbZqfmqv+La9PUT5u/wNA7MvQDxsDsDEV+r
r7jrzhxJQOJtCZpiQxqF7GkAuYroeRthrRn9aNrkZFGu6SVAsbkqyHN31K4XULY3
WYUwIRhZ/SOB3TSDWCTkg2upz7sxjssGLFqpU4Pq+ZwMErwMOfP1NOEHJqKAplPw
L3HmcY16sko60mkBvnS3uHI8kY6YoxjABjHYXgeMcuuGOrgLdKmSYLIGHLUMvzfl
lt8J8VE8Cq8yz67BTvJXXph7gV0RA/ev+CM+0rMsNNhCXqSz1gj2nPQ4PxIImqrw
GGMXBiVadwUC/NfOBDVzV8RSAEvlrdNr1jM1ExnnrAJsYUNvu6M6Hz2TKzx8GpGs
Ss/j7FnXowIhpLvyjho1mIaWf+7ff2CkSzdZGD3RxLYfBVr2Vv9likU9pgz8HsVN
71BUT6cMt9prpFQrSp6QotPFEwaHgQ16cvRZcgYq4zjsaf1cuBJx29sHa/DF3t73
//H3HJpXknmEdzy4vmL1HhJukRtzF+IZ9jDBJJHPCnBwGdcKXqLNcv2FgiJyrnle
Le64rp7NH3X8pVhLuFWOUyZmdoSk7TbgZ2+xB0ITK6S84bVIIipoeTR1RhYiRbhc
jfrU61ZM8ckL7GZfKqKTRdreZcgWmIcrNrvGSqZRMKnxj9FtHX3cS8t1rjJubyhp
jNcu1dmJpBNLuDDOQ2g0zn9YLhH7giS2z68acJkGySTD/8pwuDlqoi1/0eLliN7N
Iz8cohUmIwCWc42dahKpBah9UfbqawPYU9vXcq0UE3YP2hLuZot71TZzdAUwsldX
o2kwUmyv6v0xKDB9W2+NQg6M8H9Vrc4kExP0Jjd3uwQHB49D2THnesHKANJ/lIeh
X0BBeA3Juug2M1YCkS+vPgQ9Aq0O/JZVOA+wbgDgQDD9s6uWvQhfvceABo9eiikh
hn3CZCQMd9b042PfWaryILO8D8fvQVMn+XigGrPgH8vz2UwBD1HQjs4EvG5XQmFk
aYXSBuWyszqd9cZQn16mgsu5ib+Lb8ZLEwCvdzGAKr47q/d1zt/aGMMoTJj663TC
urRumqtfVu+0S00PrT9PsAv6wyfkn5gRLMDY5wPEHY6Qz+pZeGMoNJ6AvDEW7wGp
gWAACRymq17EN5BvbygxI0LjW7xvvt+uuttUJRB5bGtQ2818ucTzglVY6dxalMZA
3pi4tOYrncu798yOqTLSVu2PlhuCbyosf/adfNABPAUhMxgJAneu1Pz6kX5G8Vnm
8F8gKQiXGmOcFUixSJ1w2Qrs7kaDaW9RCJVhlsSYMdYWUqK08IrOP6GS0uYVRuTU
je/q+V7GkvJi5p7UKsHaqp/mRHotF+1rDjUNTvzBC4JL/wTn6WgSFehHEtQdw9bK
Hicr3vPAA9vWmElUnVI1L8PZ1BnscFwYG9Y1d/1iYWe0fjWkzF7qGQi4cjwAdQP/
Hh8LDTaavpovBDysW6vRCBYLeRKDuHXv4i+0JrRqZ9SfvWPDSeuHug6Rna27EeF1
PUKWkjL4JUg6feXrLScCVrCqOY/7cLMvZUhAkDeDFDUePBXma3uZaeXfVUzvMQvT
lmuRA//p6zKtD8Rc/syCFvtyFLitbthZLvLhHgD1k9f9nR+pxnotxZl7P0mC84Do
8dGp7JMcSvYSXDM0qZsNrsJIiL5hynfXmS2NqPWamctpNfDJIt2QZu3i4rr8utLe
WrCz6ZZSEE6qrFDepmUGsYyOAe5A/Lfrf0194fW6rdvVTR5+8Onk8ShyZLWK8px1
FZCeHlzlvfC8rAYbaqm3F1e3F1d7EhjS8lYJ5982kWOsIhUGjb/iQTYLOWVcquD1
Nguf4Ott1XhWezmM+Evmm4iQDP0biwasB9ouUjUGcioxBfQkx9dAsTWQrwElFPtu
i3Zcw/zeVZ+hcMcIT1Wt5q9+QSa5cpxkP9sz1Z9S7dLny2hsPPVYSO6UHh8nokL9
Hf9NcqToAS528ojteIPLAXnDTcC3xoqos5i4dooocFdVTHMITJ/bvfWLbez/cIX+
YDEd58F0TXIIZw0VucCYX0pWM6G+S4y2jYS56ymHGeF60lZJL0qnJLyUIh/2mhc7
M9hB/laD0OFOu5hs7uDrFbZMHGnCCTu+geU0c8qbHfy0Iu7t0cyHEUZw/JqE4QVw
fv2owmcAZxhqcFDOnmJRMT6seUuMrVme5/Az7gYhJlrZAz+8jz63m6gtpgnJ2p5e
BLUJtyhnJYv2hd32KmDKbvccJyI9JdeVPPaSnUF2s5vPgFszxZXEBTKLmaAsxQuI
zchmuaKMN4JIxUuMceJQTnkZYyuBaoKDMXSEt14lCoAIwkw6qPaunnr/091tC4KJ
/EMpN2LLdg+4OXf9Z7FEh39Z7erLGyAAtrN9B4Y3qkm0kxr7WnqP+5L6iFjBvrzD
oWzxx5BR7BAnIaauzJr8yzORp7e6hi5vB5thZfLoly5JgPa/mLT81CrMgoPfowDp
LQB59fXQubQPK+uJd9EPUk7L1z9SkbU2k3PclDpzvlm+NKzNlsmITFD4Ek62hE8D
KmAiUM1GnseAGf5TUxi7K/ZKiTAz+v7n940V4fOuSxKwqWgwfOkhExZQ8kGu0pNc
X1rarjcxgJgoQQ+0P/BAf+OYkxnWlpUvJYmkU7UzEKR8vjN77GSdVANMn6tH7EJJ
LMXuj4yzLxRtZp3UuZzhPIIpFDshAbbR+eGNRjKsLPiamg4BW05LYbTbLlouwiP6
L5MIproxWcd/cbhqZWxUmkXJBGR63KUcINt7E4MGo9ZT3rdI1UXePPlAMK1RSofQ
FoFD6Dnvw9dPp40LFsXIImWuGdJ563XIUn3bh5m3zvwpwFVcjlQqYMcM5PRCVuD6
K7FMJCL+tfRVJpgzqDlYFkQfWXwIFeDW26xPogoJIm3heHM/A7giUyNmJA28eoWB
HtYvuFSYZZCV0a/3kuvfiRYpfKKsPWwlIQCySj1S+7rYkQ2dFRJPxxGcNCv5cEPn
yYDqJiaRaNHrYMIId4GTLfY3BX6aeNyPrJRjGbNjbqmztDARhgpFf184/4stlUC5
DMZRuXm/sjLU5+pxXywDMIT5qhCJqBIW1MIVQC24i9XJ/Ea/RQTgxF60zjecTqdS
H/cDnF/kK7Xf/Ai+ieLQzjee2t8uzk2DNqdYDvs2s2acglLCxZfcThslk/2fobN1
Wrv2p5fsC/ecmoSOTiiv/NiVxCB5PV1i6SMyjxvralQ3mog9FIYrkJ2ia2kfDqLQ
+eUdANVX+xA5etei94sudTq0YtIIzLKDJgm7JRqi20OeWVmHGPTTjQ4wq7OWtWIU
S2HmIACYAx6FdeI21sDRwk4eTMz5CzJPo+gwUzZ7pfJYgASm13H2H+6TX079JHQF
3PCp+4eVzyjACfq+pX6k3dFc4byxtdQR5g6N81eK6l2Vn6VQZLbXMUYcOWXweUXL
4Ji2GDJc4TvHWvOnvlPAdeflWxhmn2WEEbtl9yKvLKn7nKGrHKs3xQCqHlcIolMm
KBrbC7I4ZBz9/+FmcKt0uXWOnEIaI49yzsDbGAFuTpochxgaKPoZw+N/5ifbxgnt
ZJnMlD8PrhOxLXqRJyt6c1IWsgaUoando+4irUbbYVQXlrDo1zk4z9rUMBZ1O8wy
4vJ+Wy4DfpFI0c5LJQrHHOWVt2sGJUz7wLDVe3Hd7eJqqFNbQLlvf4ea9lfV2w/c
YIEhWy9vNl9fouNGRU6cJBwKTVSkC4H4wzW3/hWh9TKFnCbPguHuxCfk21cofsYW
oLEx2/JzRs5qFVhER9ms3tfJUiY0ih2pIIquwwZQSgo43uV1a9JY/xy9LNA5uwcE
p2tsDKMMAlMr2/xasGiEHnvzez3i32YYVbAFAckSTfTI1gz61p5FWGMBroBUIzHB
dVwnDnOf7+n98U/QCvzgQ/zUYQV83REZ7L6g/LzAZbETi8g5kec03cKMAiRH+YzJ
gbroJwkhBj6DgJOY5y9YFoN8tBDiGFGJkTpq/2VUY5+3TXje4Vi+0Ii8cG+ZtLER
PI1wXIE2pn4R9WPKKLAQSvk+YAib0Aj0Fk6iDfkuc8MgP/aMNyokm7t1XTiahDBR
RXZtwMPFWlEF1zpAP3/h4KeEmwzg32GIirB1Z5xPvyeni8/yWEg+Nobfc8mRIKW6
WBYyeEi7MakmoN1iKGsWYue5lss5cdNfbpvVkWRAJawFjoqfEqiAQQWPIc/+DyWr
cchRBl1j4cPinL6hE39SmpT8fPqIo2/FthjMlU0w2ZIBpcCALn4wQlDEUCPofL/D
7bRd9HK7V/Vf3sECeUa2zwRf25C+fsBOreuwpNEVabw4eVBvNxqPJ1PNAd0r0hu0
CmcXNoptv2AoSpqtQyu96OE57qaZAZmnCd7YqnKn29pJqDvHbXDnLwAiipMPaYdF
EVgg7FbRIa7atQbKyyoqP4gAhUxMnKxxwQjMlYuMPwda0lSN624Ya2fV2UV+p04a
fUO1QKXcFN/wx9JdIQz/WJgqlA0e1IYALIqSa/3hpZN+fAV3NKcQLJfIgzt3Fkhi
e6uOPYbg2mEGYTeovzTV4VOd45621RedP7V+6xY4Vd/LKCI8FFqsBNm+DA0oOEXw
4w3FRgotX8cteMRTkLOKrAixjNMp1tpIFkrC9UtTx3fI2XDkXucBSTG0AtxlGYux
2rZI9Rs8RQIjdsS4niKBkxbd3hy9Om5OakSKkgb8HP9f7llcBYylIP0yAdFV02gg
xI1AdoTHcSrsNTC7GIDySVwiPymYgRzrslr8GGTLmmJoE4e8Xr6I02f2uMW2E4VM
2HjXqTTWAfhQ8aQ5/7b7+2pt2NgSIxv7CZBFRAw/WTDWszac40RIbpn0BWciTDVh
AzA248vaMQpPxhoUuvg1moGntXwS457/l3Eo9UAnU9CnklUYpDaXiJEMWRNZGizJ
ePflI2cOktpLSBt4bvyvV7v1Sey/NApzJx2zikOQPCkQC0KNcXfov340IX9B3i0u
5zcElmzM3q4ZPoAh6zteQj1PQSHZpJSaC25bu9pwuSMCeHlK2sxlobO6HD66qOcu
sT/fvBDUbfHNfcDLlnjakr4zcOoBw+EKYfKj1GXgdF7wYS8wpKHOm9CzSQxzsAoo
TGem1F6vp711PadGVb2MSGZRFiJc2tjsKBl2AhtkDsB6wBFnUrcj6EcjTE6rz/eZ
WCi1bD9v5HcouezQ7vhYpsrykCxeiE0rC3BIF8URVLp5sUBufyFfSZf3xTPUnJkx
ozUC/xTCbEw1JS+O4BjgaweSvOT1CyziS6acOEyq0sQ8A5psTxhqDtUbvqVFfTGn
nEeVSgcY7qwRDGdvdYr9v2nYCrdsLppRMlAk1F61TlulOXRBQZNzJEhWhYHl43s6
nDwQ2vWRZgkoAA9N38acDNTmS/RY+Tv898Tqgb8CkcPIW/kuzhrl0Iflejm8hlnE
aso+X6KwTVCLR9du4B6Z1gSQrmNAy5VNuwdnZ2iVzzKKjlTUYSX7VVlwhQT1OQ4A
CRKQqRS4VbLmpB8V86jc5vT96FpVMt6V0mEPF8ONcVQ1132JGensaw1yqnJWHGfb
+Ca8E8I6qjLMUk04PbE32q6g0+e3CuO82h20c1/V88f6FAYFkJIkpOC+pq7Fy06o
ZPg+3uK/Z6xppjr068wpm4Ggf6V2hQ0DzHHs8lEetSwbJWTFpdXi3n6vyvFeGRRi
/mter2syFMo80vRO4tC3vZMBCvPA8YCiMnmnbhH+gtepp9NlS8BVaXgzLtdUSROP
t4XO+I6j7+hwhQvvAIii+S+gdx9D1edJ9CGd1Et7rs9EPT6clmTUj7xuLIQx1Azy
btYyVrGu3DfYyBxBlbJmH1vEpVXR4xLYh4AVvxRmB9m+zomnc3Utt4Ea0NQPCFPF
hVR0XcBF/nAvfcvhz2g96cD/Pxe3lWPfhzzez19ISHiBY+WPCGK9Ohn3ITMf8glD
iFRQRIF3wUGUxcDIrBgrphfcIBvDUYAEfa+mw0fbXr+v2VCiBbS2TUN3rxLPET7t
SHo/KOYvurKAtsLN24k8H+IEs/lLvHOSsXzMJGMaWFSWd1veRTy+hXPV5NHZLeqw
HnUaZNMpyZFs/F8FNBekAOVo7T7ATIYYoCd8JKd19SzKPZ0toCcSvh/ft7ZmfVCc
pmx8am4XJjeT5sL1YbTXjyvtdQ6vbXGH1XIspO3hljeweIJvmKqgqx821y5iPiQR
WldHunsb/uNOKqBUdfbm8wxOfYj/jOX1ALh2Lxyw2YV6qWz9w4t6yIocozJ2Ej/w
v6kLxG04QnUq9wNVWvwPpGgKZCIddXVxOvUAZO1WHebTgo70wwRhzi9GgR9OxpNa
jJJNneWKADidJjUek8wu5zhiM+D+zSWmVVdiGBvuhyOwNsgYeMjoYnHl44uRzgaT
dWakqQ6Cm5u/fCLe8l4LxHiNV71E2BzNmqmTI+wz7g05Umz3P+RdtKdIYbHYawJC
1e3K01bhMSDOtrrmqcbRF98JTCv8Q2jBetHs6yUTsJyP5fqlHo7jQ1NlXS+z6M32
lK+sT2hHQxXMhu3YVEPJ6kP6hZpvQl0/byICO44fskM7KAZKC9WBqKtqMwYajIn3
8JYQhYftwnGBMdFWthLfLfpbWcSE31xwfONBQVfjY3e3R25mFXiwuat1ha1V9U3q
bAF2BnBmy0LUKwUdvpxuHtEuil8NSegJYC6wT5yCJCKVlIRlkHLysu584GHxYMg2
BgQDP9MeL1yA3wOe4KjI7EZef2rV5PkhSFWtyKjZqecdsA2SSj/PVhLOLtvvZddp
ZCfV3lk9GGcfDDE0DLQMLbr67PBPMwbO0uLrkuUl2CZeFmYdEPrmoHTjoK0Z6e0v
l8JUBsZEpPYoZ88sa7L85+pup3cMj0dZ0QApBKHzp7+J3UeMAfyZ2Pr7zchMSN6L
PwGxqfOUOrJJSs126pJRvwteJtHSuH/5lMAgNBZc38a/kIDHTf0kRoc6WEP5GhBO
hZx4jWbc2nQYHy+CXw739gcS0ujsx7GaZ+zrIKX6QkL0hqqjCwCAIlxXpks601Ik
fxpTXrr7yF+1tLPQrWhjopsNSjwARcfPKZIDk9jAgZevSqgvGRwlIV6sAwbvMgpn
vetPm+h/4C72RUx1K+n83Q/dRTJrBJgDFBOJai9alMOCc1iEZk9gRIvrZ/Wa03YW
hN8QdtZXNf/zhNvlzzoFHpvqTuUUue60wrebswNw1dClNFZy70rbLnw6yt0Zg4PF
qSOwr8QPEVx7Zzttz8+yzcvi4XkzbSzPUeUFOJgq048P6fg2GGPfFVtSl2cIhKCJ
iWQSH822KqqubRCEININmVWZE0LZgxzd94yiVzc2BicLnle6ZTiEGvZheAbHHEjS
V1cefxX1d3dKaGj8LfdAUyx71ImFxIDhh53AKUCWFmDxmUP7iC0JTmsq/9QWm3zD
b+xj41Hp3VVNpw8cbwXFnR4n8vVtkZzot04O5ckNo3z2fYEKZ6dNfjE6N5Q+Owr9
KhIHlN04Z5lDDW/ARSuisqm4rAnU0rW8gd81KOBR2ZdCkzlZWMQC/mSuejM33D4K
AMoU3NyVe9ptUrqd+GL48l1NE+4HntYyP9uEhqC6QWc/QQFDzw8m61vxr1uLtWK/
tLY/gx5o2jSRP6Ii+jrcFCTok3LGw4rr9pxQz3YgKNr+mSgWGWMmv3dopqWWntFD
janRBMtzrB9IfIB4d0MsZjxZxV/xrWqpzAEd+zeW5mS3SG2QIEY9bUHiET+0HB9N
boQtojgFgEawEi1bPd6exuU2RwzcO2m2UiwQ4eXQcOtDbBdgznCS9oJvEj0cO1aE
Nc62Uh9H6MwNTyA9iFytVIRJnRoeKtuwhrwKgf1Ud2cFndRSOtGBnrZqcZgyzwH6
g52R35Qj3p/QPwTj6hVvMMoIqDmuSkOV8hVAFQlFvsJuGODsbKr/ng4pZ6+Sy2Al
ZjzyB0l5VeKz9Bf4XbOszaRrIu1aNvdnX6bKZZsMrPOXoh4kCTDLblvyJvqnbiXt
a6AK3KJtrH8gaj5FdHu456Dy2X/A7jt1MECKnJzoRX3oJ8c4i+zwfT2GV/UWy4Vl
hIt4o/eaKrzmiGpVaSSE9nLtCNNh1QP2F2TZkfgPYWSPgLo2kKcR8eIBBLzycKwI
pPWoUprpVjQYQXjiyd3Lbi9pEQFuiKwnhTnwfFCgCDBdCNCQUcLl9AdnYTFzQwE/
XElCpNifT40R4P973AAMOrZILaoJnFh8heLq/cDF5CmUS2O5YIG0pMq+ODanlae/
2Lx4iVYG2qZ9Nxo5nAUOz1cmL/qvu6uzcPrMTY+/cl4irtUkUkUDEkFneVGoO2Xh
xaXztrSCoGVHJjk9lAmCL/hurOfPeyJv4ZCG8WFCbyWz/vqSxhw8PNdd2Tu8vMxv
uOZcrrJUibgh5qYPOkzkJQTdqPOI5c3GKbTrNt8c5WOcGM5HKPym2P9g0/XmRJql
fgnKo4l7Sog1LtuA5UcDVKgjFgoHU4u9jZDPlNlf/R/+6CdRm0n9+pmQ0ntZzSbi
N/MJJzknKJ2qJoa/itnV74h55qOD/BQaPgEiD9fNt2YvCkFDvPfePb/W/2IQUajz
9i7r7wxp+Z3B+12Xc7T1mqQdsL88kb4bIrEVsq0HRBbt6Hkd4xmq2iyvh+0jPvd5
NANoVaJ/I0fH22cSDr2KW4+L6la8KsutEqRcMCpwU65C4s3+LjGgPrGcHa3oZ8/G
6Xrw8ZIYXo5grCWdQbKSkywDQlqViQuTJq/BefNfafNZnOazVfOB/DF13abCP/Nd
6brVSqRRsYNKpw2sXBa3sy7nnfEXfsrOEYifKYY5McGawZ+mO1HhqaTOWCyM3kpM
GpHwb0qg1bzKaYI+lZ4pC6rsL+r22PUD12c6AdCz7v6drJ9T+nOV/TBD0DDun8ca
+6+rWxcutepD3Lig4h0gDg+MArHJFMnn+fcsbOVqBvH+fs+C5ZARye1hqIV7MWvW
EyAL/bDAaoasCyFFG8l/ZamnSV6a52Hpt5qUlkgeGSOlmY5HtOvnQw4droQpFs9I
hLM3dJpRkNWSQSPw7uuy3uV6G9ZjrSloY1ZfcEEP15WttUfknGdoYjekgDza8idy
qBphYlrd4Wpik5vMvSzK6QSqszv4pcmHVYUPpkUPVf1QYnm3e6A5WsUbBpQr/GcU
TGwkGFHJu2YyZf6PcAE3nUd7eeP1k98yKyGdSJm3Z92B5AfygHhV3SWiztAvrSfT
y9WQja73EC2foQbYVDGW07/vmMhDWE0aq2U+WmyRWhJ40BRxb+9/16xBTlNSP1mV
mrrxgIwdupM+fpAlY/B6hXniDCgx22Swf+1iNNc9seQqedpXYbUD37xLWmKwk5Ly
+UQCPeKLNVaE1vt0jP7mfxFeccdipIoIeE75pXbgCGCeLiY9TujywBKkktvCTDLe
0eE/tO6zWcpR2SpIPSh8L4KTP4qryoip1bp1htFin/0wE2aRGLXpCx0Yzm9k5VCB
YfvNdIQOEIrnkba1zEHMM6KzPnm5vtUNHBc/ZpEcWl6g+Yk7/VmaNizV9QVvB4v4
8X6L3D/XqD9ClwRA588qb8h3OkK5UEiP6czpqHHXHGyEsqlHK+3T8LkbMSJSZE5M
I+zGEQAv0nq20vZad7GABQ27OEJMn5s9JleD94nA9PNDUVi3+C8tdZzDO1OlbzU3
WXpQGW4EvaN8jfrqC7u29C6iBbuH+e0FZnQkO7gcCyt0kJfuacXTWRYAx9L3Y9Jy
tf48eVyzbeEexW09bJxKSwSOGqddbl6nIuvqzOYj1sO76S86QUOiqDV8Ldg/K7ZP
1ENYgH449T3HmZey7GJ/7+7hdSrrA8qsFye8wGCEQNC8WjovO3bMk0Bdh2oKhdUi
EqOvic3YCr4y7O1gHYOAlJh61Azz6W02bzd3qX6q6S5fspWTEjBjv8K+AR/y7U07
qkj9uK21JzEECrwX3DhS/wn1gTeDUxEqlK0NuwjcGYjsGPZ0+iZl8G1qxSkSvuAC
y89f+RucgLj78Dy68ENaJ+FIblQ1WneasekTaFM7JwItGFg+2FNmy7G7OJAcSM2p
2h1VPsVf/hOE94XCKcHvlbwTu1mGvtI0C7epVtyXCvDKJ0oZo8usHuaozW0NJmb8
2Nf7qA9z+Bn3LKHKHDxOUu6yc3gOemrpg2PkNJQ8cfQMSOUHOJu8ZhREAC6LFsuf
w5wdMtqRpI/cZ56qFaiwbob/1iajy6utw6BNPEdaGAhHLCs4GTx9STQhzg/pyhqd
MYDyxr+5+Rc8rmwuM/m1C8v4v+8DXVY5PouxYtxqg7o68eUixBfsJS2HP0yNd9LD
ZW1nhXDQuRme0NlMo8oFsB2iEgnykmD+wce0g33+lYqHid/A1PO0SNSC3FMqtYNd
BzjtcXv0V94jvuvRQsZ7CEmAEBxzZ93UhF55A0H1OqAhAyA5e29055KB0NvgOtpE
Eb+bEEetb0w6P32ySxjIR2wUJhFfvk5wSyFbtFdXOIJYKMc/CQ89jqPNF/RaoI9M
fdG7eRi2MrgzU3GowZ59AkMJ9WCJvVMxaUZx5r46oByZ5jSQGpGblGAitA1um3nK
m1sA13358TPksHJ55PQbrabfJ00Q+1OhXbgachtGuU1K2Vrf1PCzTLu1eqsRbxNF
tggs2tECvdIzZr+ZX5H7iuzxpWAk9nGrfnjs4qEPQ3RqJ2q69Id8tMLu2GAGWi4e
Pq5fskuBX09FAFNmLkO/hvixI9pqDjp60E2MoRVzhNptumUFblKt4aJ8ymhG0eNj
2N6dq8GGffLc+F2b8d3KgFBPY7gjh6aODYuEaIfHgNqsgkBeLQmJQKhIgCuH1FfN
NECEkC4/GccezfodM5l9axHWTljplk00RX/04dLStVTHXHkwh2/RnXvJwqYb2aH0
QzxIigAQv8MUeHQhiHURRd9eX5fEkIMfmTkUudEphqjdLah+2uMZHkkoGWFwIVqa
FLgUdl6xy++73jMohSyo89GXL8JGYJM4RQHP6ydpdA7BTycVsayOY0GQXuI8V0dV
2NrVi0Zdu9GFIWn4LX81GR2SduwwxnBWUpLfM7gj3ajL/jMTUh2xI6UYspKtF/g3
dsfhJxoq8XjarkKAFKtL4hVzntsRzDV20OVtqzMEAcLG1UgaSfcs/H0634cXV40w
ys4Qt9iy3ClozG51X4xmvhTZVLIZ4c2/oZ6RRd3HDlFQfCAXjw8ZPwtLEOtZxfWD
EVQkRyu9MphIeuPHYAFgcdoyaNSScmpim8nMFsbue0k0tv9rbqHzC8GlZCFBlzDE
38ip3P0EglUIAcoIYTOKLWV4fn4D/K2dSH8+eW+zTYjVpgVXaPpnbs74pGcWkEk5
MspSR3DUySzCh3PwuIia/TN/kMJ5Kg3C+7cJwx6zHSRj+2SlVc1bX93Gqw91/oNF
Il0dep5gm4SdcnHawAJBNRUXwwoSOXKt756lZKrKx2agFP1/eEa9nTpPhoQYOttB
nZvORF/a7jiVbdN68h/LMJXi476cxji9yaq2jJpbCgfQKu3BXa32l0I1BlWQb2KF
D1N5/KbjhmM7BX2gM3SW/k3Nqp/XN7x70ErxTj9vYkdMMlE8pWVmSZlniY0l13fA
eY6DeGtyYw7jBUJtjacfsMu8nFqnTS1vlWSImYnG9ZjBfIeQkeKSp8rbHbdZKu2l
BHl1jPS6prifZuVsdvTWlc2wt07sqPVNIKkfVMYGVzOUEBgrKO0Qg1uhvhkL6TAO
8TCi3SbbndX4HEPLW2FaYxun33GSzC1HSXEeRrzocwWq3BxICHfaNs7F32v5fE15
WM7vnPeEOdJWpRpJJW8B+dwoklr5xXPkjQcjT/WldBY4QlI6gjS29H/IcQaJGOiO
RstHnqJfaWGwWRm4pnXOQH7Rb2QUsHPpszZOoLwdcH5yS2QSYrH0RZT1QZzM85cr
h1s/+cRFMvGAvbIx0MZAIWiDjNsMX3mTQUUIHSHpQsIeKUjN+uCGBSZcI7W9w8yZ
nHBmXj8oNCqZhEJYJCO96abODb0FGFYPtn9WKFVk6BW+NBk0LK98uKLNvOb5M5DP
jY4T8HyEovrikpmv4fjal1om/rUuBlQAmQSYPnbv8z/MC2RZy7wJLxzYCuEiFIFc
ADii8fxUBaeGR0PqdVw0Q6jTXQXqj8AzW2KVFqKu8WS05H2wCY1HiyGC6N/tfISe
qbWs9obT85YrlmXaWLz443Q+1Pk5gj6rxA9q3ZjfAmvRD1ZPu1eJB4C/N9P9lfD2
w3ANCC3oNIysnFQ4P03HlASAQlWCB5RxsIKEf65NYV7Xa7DbqLJJTWk+parHdMOR
qrS5I+IvCOhprPl3Ih+iqSa3ElT+F+PtfKOQsgerlThbyHCPZR/O93V61YSU3nmW
kkyFn955Zo2G2Yx0vvFw74+VYv0k5FlSDXg6w2EN4yfY6M02vdGVe83YAtjibJfK
vlV/ntp9N8xx184TueMTmb/rVcGS4F0J53WMPzn/vXVELr8MdBPAlaICL7zGwJtZ
57Doezp0IBssQN8c5OtEhiwXO+j1qMhZnyTQ7gChsSAxYpuIBa5YyY97qbKLhqr2
f9/YfFdeK2DulSbO/N9pJdZ+6Kk1QS93z4GI4mZAao9vshLyVc5/HzDfO51VuAY/
wgWwyEhDXOYq57cIinWpIQeVLYaao8FiwamYfqJ1MuCHWnokPI1d43MSYX1e4DQs
y+pbNIp2f3kZuS0L6CmIIzGlTgjavlkzWU31ErK17yRb8dGKhQ9009GPyFI+CkZ+
EU6IWF+jNQzeNN+G/y1OrAhiJbe9HSH/lTdjdiNmuMtRU8BLH5HKjqEfkgk+G2Yj
VK65WW3v5XkQvlCvPFsbhd/vgwy7DR95uDe2OqOjttlYZep8axHb9rZHZr8cduFe
mmQy/H0XVxb2I9nnkEiz2qoH91e/C6pbqwAwZAqjICEwfOjPEZVxrRWOT+Y+biQE
0fBx4kM9AZzflfIMThi8t2f7N6dTIGpwfteFpMi7hzh7wopjTTULVpPGzS2m4HYu
IirbS/pMtik1ZHFx7LphWc5iUgG1EPIveW7rF/dAHwPNk/i8L97mzvkDgOM1oVkF
PPZ2k6WRckfkuJ64hPM3ZltkcpQtacYa9vNsU+6l7wOOsNnRiSdRzMTqrmw3nHy3
80RnR0/jdTsZiaMdP5DKPyffESgIyCzRuf8B8h//RueEIktpElMR1ZvSnFBOwf/j
5VSWxxxmMYDKyaX/4/uMCe/zQJP1D0DxvWaEwNGucLoSsFYZRM6nRy1iYwIg5KfA
NDO0scj8+15fJG+Fq8wfMUsD1Hpy2S0BNnsS7R3YurVlpGVXKzgmOc0KteUMqwhW
KrEGefoBaPvPJK8vA5CG7MPO0BTUmBv7vEEY/4N+psN4kuQ+BkPaNSuspZQxdY3N
OetdNVTeJcF1GFcdgskANOedYg76c1TDeGFmz/W/hxXM+IRuLQuXyLQeKoGc8WRC
3YH2NgtxMzrjjQNEN1c+OUhLlnfkyIk6PwbS/VTT0kJGFtFiUEXpde5BGKS1eoVQ
gVSLh59SdjwGNcTRasMj0ShMTzpzchz/FjYZOA/cCwqYaCWB6vv/lYHsx2dNgCGa
zc79elJ52aq/IRA5JaTf3EN4Pr4vZztm47j2+ATkd0eu7Y5WIzMoRp0NZT+JXYBB
6DEfkTSGUG7n1d5v2PX1JVYWjUC3Ekb0q/oWqLpyYw7lswCUqI1+OuoXvd0BBDK6
fHFPTcAjQ46AR2+fb36M+EuADvGQHHjtxB+Aa4b9nGY4ugwAxJ/Lpmv0wdFJlAut
HqPhlAznYVWrMrphtGrrkyED1uYDeDYGXVqEyvGdTYtBYDHNnJtKtRsipWLkFtqu
wcOpjux9LzTuWax5dGIm/pRhWS+1ubbwJO6YKUG2cZOpqYbZ5Gpi1+CB1aAf5anX
FA+MJyHWn35CEuFPaU8b4zAPFssax5Abokc5Nr3NT9VPt5QEfRM1OSrGBlAz8R0F
FPiWFD1LsqTmJsJGM63Ccxrk20LxxvXvezTqq49ocrqpmL1l0jI40upYBRMBjEZm
X9JpPr7hfL5OhyeUypZ4vF/VS4rlKVkRr6yn4BJPoi6X/BUjn3P1wwCOh68dwjOS
QBS3n/K0J1mF/8SyQXMTkjSl4FxYrOo2xRSWpC2dfgXggN2M7U9HhLvo/+RZgVaU
3fbuIIVxjI3dcTvFxdahXOvQU3QB6DJjysHJtuNkZ4tH9L9kl8pgt5Ah9dH+mqyX
R17dQRlAHcpAZN4qX4RBtl/c0qa+Z8aP+wa+o8iTOjMcDOdf6yTnyO8lg2alPJic
ZVnW2LR1EQruKxTra7L9DIzz8PHZIOLArBzp7RZ5Bm586A/YxIEH5HNmJADLaJyI
GFa6t5C2/caP68jxzGtH1O365y5mpO2P/c07SCI2hXDUY9XJeaHaE3/g5bEmflsH
lDSLskkgdVjGtrfBhjz9h7LbL7xOxGBcIfLaZm47jMTPNGFvsGLNHBzbGkvV3v7x
ABtC3rnVlGx1bKSZIr4ZA2hO7Gg3otwZ8jkWwvJLk49TuzGiOiTWBz7ua8dSBKUs
Ebvw9Y0EINgXIO/Jb3jPAtutfbNWPlk2K0+dnkU32ddL6Jws4WCxBQiy2j6Sedat
vwpLk+fNnoWlIxA9NmHD1m3X2eIdfAQmqtS8VR5OtJ2Ky2P21sckgq7FCCuY517O
FLHbjaJP15yLdcicSROCfyEcpzDS2sSUxoyHvqsI0ldmgxmV9073zBHplV03q1EX
ahPmL7AruwicDs7OU4Wsjz8wY5MggYYpRJIZU64ZSz3OKpDLBOGT49FX3eK8A2HY
YccDA4340EIE3PoI7s+biCfh16xmMUcsIKsbnOF1PEwocICvn5zsfILig/NrUxPA
4PldcrxOJmSupQ1xD/FhWhqkPBOxoeU6KzyLKbtZl8YQEbjFy24ilRiYetGUl6cn
hRRjK6QIOSwV2vSzTHYdEei1BEcGrd7551b0SPk2oCcduGlO1Zj3FKPKF04VsXfu
ptvpXKf5zHoPt94vYrat+92p2Jc+8WsWNcOIWJKwYxiZc/LMH0WNUBoTs5ieMwSu
pM0v28qPTWngWM4VoQfMFB2xv8fa/t8o5FvPJh27abX1QkoFKUkoL/7ZIObTm13X
p7Wzv6wp3vgSVo+KYjVzUeho6rl8t3XuKPHbMeyVDkTraaZ6K+ySLpooIiDzVacm
Gt2lMRM6bQDfpBqqRracnw0IR7ARh6ujzwt7wVNdDA1GF9FErl1+nY13O2bnrwEX
+mzl6GpSF8s+krKJ9W8cpZEi//44P/eg/k5xnVh3Kd8pQL4n2225o72aVRG3khAd
ZAVh4qDZj3ItiRu27zj5tIdntaOdM4oiRxidqeq4YA6vo+pgY6QySJrn99MQBBVI
zGFnd6nHWugJNAATfF2k9FFkrHyqpMAcq3C78kr4jGM8D15l5FBQCaue6XfRLM4Q
q37j9OnG+nRp1Ye6hEnQjursZCclJeriAt7IJtyU8txq/gCwwm+ug+SBODwGQOnZ
S0iHhFLhpwlU/nBPN87orvqV1KmoPZ3kG0AqDdQ3HvllD0DknumxznnwmNonqMei
9PnAPdpL/Oybu8ZhvFukxFPU4UtFU6e6vMibVrrOwrqF8g14uqVBWJWc6vHP3jUI
5hrPGgup6/aTwLxPENqRYUMIW36wpgo7qli+q2w7KHzrul/sjJ28b8A9ZLcv0pG0
k7WWdCil/S3cQvoL/Ce5+rQJP7/qacQIRNM/g0wC+721gYamaHfuWSar2SB/fz7e
nGQKqF2IVjYBpizx5+ohUwP/GGNUtdKulJcs5UoidTXpM4j1u5saAmFzRAWP28n9
iCRZA9KlDgMPOK0HZyLbTjdh1+a39wmIJyYnAr08r5U6wJxsjwQuqTK5GWTJaN5Y
Y3DketlSSgZFsENJqkMPpebwvPya2s8Uj9mELrb4GLYEjijFGxtDUyfkHeYDNJm/
Xupw59qzMuHALdzQcqy6kv/t5HcSe8ZYgFb57qVnShT18glcjsM3Gs1LMvi1ym3y
9hjIPPRGgtHt9qfFSEPYg/cnC28R0lJRq7wiwjE9A/NBjPbN/oT4YqEGe/c5jEuW
oXbmP9thn/taJ3sAkxM0GOn/LHa7fM3E8oymXlch7NsyoMAFkCz72PpEvWy780Jo
je/IrHRY1UATNYOlsqHTcOzVuaL6TtUh/FAOOjTxFXBf197tOV7FFUsG1ovBkhGe
1fkQQKHETrKv5jlC+DrxYgNZfaf5TkbizwCFL+kYTybdzpE1nq3L1paFsG59XxMA
NCkxTMnrlmCHo7vp1/q5tkmsFXHz8wo+grQiHjvTCnabfo804KIeLQJdXtWuIKll
aDNAsfSmdgN8bCrU/UL7enUiByCXr9do+sJrUqO5T3GXQgmwlauYTvF6QGKbysc3
TU+t1aJU6pL+crTOLZvpeg2uDF6gWyXnxrS9D7yqwruW70Jn6Qrz0yls1sHuPfPo
bFd1IOYdHeuEwNy0I8E0RAmndFNDjd3wThw+Yk7wDxy3N9Ad46L8vWAaTn9298rO
iLPrZYOllU29XD4MJww3tSoEczLgT401ebakzEOSqmBW1w6GZ6H+Q1qmUoO/qnsY
2YgTAt/kIOpHt5PgIdQ0groN9Q3CmINr9TI2kHeqCM1EwPbGGM8Fswg1bsqcN2XC
qMRwYAXClPpjLwErhnvgxTwtfyKkckFYBjYrelTlTwoW8PX4h2ABjt33htPBYd9J
gO+A209OsgOpTdLNqSvWHAAIepjJqJI7ydWM2N529be4hVHlQ5zNd4fEGpZgBM5+
5S4t8KGc4+dEqi7BWUsG8ijsXqDeOY0pO3WgV45MVo+kwezJuhmFqm/+hhwd1Dcx
O0qqhSjU3QKRSFNGtMQJLkFtlbx3rqcZCUCcyAYjMA8eL/wJWkrKXUN7SEX3MnOH
5LoDOvTOTFAzwSYwuNdp3XmDd5FrCX7rT72waf7hXIvKqXNM6yXaBco0zhZ2M9nG
XgF39XBqEmmCfu0j+xebefXib0rXjXlIL+zjja5YqzlgjiebhhK/llKRPqByZlGD
p+31ICsPtRcgYNKIdPvUApNTsQpLlcaiy4g57Yjs7d3Wtzb+UjN69X/GVxRFtEn9
hHlUfAEz5H8XGHo27xmt9pymqLgZ+E3OrNDGaN+o8inFhNblT03oCwusc4PaliA7
IDhPZw15lPOIUd5niqa15/4k2txwZeutezAucOCdFYKo98uQ+wv59w79G0N8wheR
INA4fZR90qvaAEHEpKQ0/2gH87R3NcoT/sGGOqcdlB9rP98PX4h1XiFEW2SwOHAD
StjNASf7nzPqEXEAbtNcIJeBveZE8i+BRmJcPIG5Cz3mXW87bdvbrn0oe0zhMmjm
eiNBuTjPT8Cq6N10VS0pGr5WQ83eLz8ANHCpQMHDvsoV3LWBRV1V6p4tAt7MEH0M
ZR48JC6gdFUijsqLC6PGrP9scSs5UUEzB08tPEUqa628QYduwrgN2A1bksokP2Qy
/7IAstN4e+7LM1YTHqAYe8kA+4DxZ8u84pj/RBm5mnHMuNj9b+2GFRZeWlkP1GKN
hKUer4TGEmyRWj7J+ND7rg6h4UGY70+IiGTeRdLl/2BA8P/cHcmnrauCHX/EvuRi
r3OSVJB2D9vnkEHonJScqAUW3SdoLWF9357JNU3hpR6nQyuwp6kjZHVSeA6vLNnq
Fpe5RNCEddrDB7winPHgR241F19bTVvIrwT5YdTovZR0mrPW8D1joWUTpagIdVZo
RP5n+IwUPwV4EgFtr/miUQ9G/69pVpEvL4gmAMgFSTIY0zj0yZVqUNbnmGSxZ24N
VdzDWNdA9KkNBERuMGU1HITkiWlJijJvwJDHd5wjuVl7qly0JbGoNsMComOumkl7
DNrOJaC1vlYlPxnDnbiqDHF1keKhE+eRmeXP6fxpjux+JsR3FwQclhl69ZIgUJpU
Dxwf150bN/SyYtkw6HsGqaXe0bG5SMU00OWKwxYkBeiihBkc4xlKEWSLHttA8ujD
xbMod57kIm2gvnmeA38fSRGCfHpa0vvx7GGNA45bCsvJoZceyVp9xU0tut4zItpV
kbZ+FmJzCBut5zPySTItWnu/DIwbFEr2MvuDG9FLfaiOC9j9IJ34gQjt7T2XpcSV
KGvrTbsiIR7rc1Ck+/z0WxmYODQ6y4mIkSira+/spmAnapnRmf+IpWxDgSEPXr+K
fLkmOZ5eWPrhWrAqzRuQEH1NmUjQic2QT26Bl5ny2tgnoFwR/ccxMd6q47S/cbAq
Ue8zsw0niy/d2NZZ7iKXfXEtjqqDrZwZcJ8nVCtDRTQzWJ7ix1catnwtcCO3tLuz
cW57/TdgMZDbPHpUQtCt+T2JvU4Y7AqMrbKD8jN6+oViJrxSJyds3jRy/Pi2E5rH
M9AwDLuxGxylwezV+XcqM+Vr/UKh9dbmk9DEXKl7CRlAiVIlCugfrj0w46n1M435
fzRSTZY57NhZNJpAqpNL+VWGsxDrvj3YW8AolabysGrDA/Ul89iZurhjD1wgZVnH
/Db517pWEWVXdgvV18XCVvOTBfqFZnmMPDKcWTs3JHI6uQzV/P5Lj6ghjdXtKF52
ItR4j6XCWxmGFlc/7vSruoKeBnQiYVqfSprZsd0pJa1gbgctwJQS7ZYY6NrqPwwC
DWmg2EjVQJBTOzCoZP/pAQSvhxxDIwt1vBPnGJqJ9PF98MlN3O8RXVCK5E3M50Z/
yEgQDBwJLFnYFKs2vtXJ8dvAX2BMraxrRnJ6tLSHyX0eq1OQR7srXTpwMKVOJK1K
VrDUqZ1EA9umc387sFIwOEh+ZIVKuww/nMvv0o4SMJr5bWUAxMD01u7IG+KMYMcH
KhgaRjtzWgsyaqZ/PlakPf1FykgMtjk4J/5yogAddMupDy0UMUwycgjvdorXyquM
IBMOEpcaEd8vh3IhzFLokdlOgViz4Ex3/OgiaP6kpG+fs7S+HiswB/uZqWcGfMBA
m159h9LNCHjinPEIiSLM+2Yj+X4QlGcJGpLqYdK5TZ4H/ylW0BDCE9qUrvWBy6KB
49Aho45Cc5Sq7KVOWB1PEPTYwQ75MZr8BvWq3DZNI/vsfHiwWsqLkV3IPkILc746
wdl2lF8jpGtSpKOKid8Pwq7mgb6yDu6G3t0wCYLHM58Y1RAoKRzPJi2qIHL+n6D3
59Z2xdI04Dm5i8HuZUzS6LDuPOfo20LSShI+cKO1vpd2cD7HdbDaA+niv7WSKyff
OlzVr9CYpAWaSUQ72LoPTPqZwqVj8EgbA6dtNC/z47wLCx94/cMSZKjs+zYP9Zrk
Tm0r9Ehh1swEvhL+jt6nFZv4kBag9C+wYgTS7pv+J6tqqAqI1YUqhWarjgd+aiFY
kCqa8wa1PTmLzdA913YPtz/H9KCLvES/IX7g3E39ufB4TQsa+Ly6ksZgVvInfPiE
pAkOLIWSBJM35ND95UurRILH5S7kCHmGZo4aBnt62NFFxwX5T0NkdKLGTUw39CT6
LCtpXPesPxM1bISvUJyfuJspb1slKtWLls01hrBWo2742CxgxNQvRtfkXTz75OBt
VszcZO9FOxcqSgS3JdxqTCqqNbnYuO0ehW7KYL5S9t57saLp1cLe4Gn8hI+WMBGi
IRmmIVNOXMuO7bRGCEausZNM3TnqzwGV1Txu1tlOsoa6DnYxzB0JdBDc/Gv50DmH
A59MW91b8Y1HVUMeTbuKnIBHP31ZKKmTK4P0fcizCIdX+gAdHf/BAoe+eGa9AP0Y
LuXSRuJdjlHvII521r4vuJhQdT0XjTt5zCaJnM0k/dNpElZEl0E9Eo7Nu/jiHobY
Cy9IewIffbVGsGdHOSpLypRGCrP58qCnZoi6e7mm0uMyzwKsEiik/VJs5lEWIL4Y
KZ+nBPGbYCYhIuLvEcjzQvUmwT3FLvzbbbKztqHowIY596yMhElR/DG2FDkPmVWB
T1bnowSqCiXzvkbjcFIoVJ7UcZTKCKbcfRo05BbdS6lEXOH4qssipze9z8qgWp+2
Hy6kdcJsoaRBAVfw2JxH4OuERtTkF621aWIgpyIw7XACRbQn/VgEIjQTWSt4YCuL
RQp7r7qxK9SMZI5sBBKx3IordsjD2+gfOQtfuwMFW2DknUbsvUxQZ8RQiZ+kzk5W
ImU/PckFlUVc6XEOnUCZoJ7u+fCoNIK2jAVtF2B0GROfi2TVwkwRhNFFIwb6BVEK
ITpUTWN8Y9+YZVBsDawnJxb0vXKJMJtADsCnG/EhJB1p75HYAjzcFXRR66LP1NcM
v0aFXEVyF2xY7hHYZ1PmWqvgxgd+5fQKStYnG+fAV4SBOsyiqIHfGnKJzG9c1bFv
aukGIZe5OiX2f3/il0iAqesmjmrhXZ06lygSbdq9cnKddETdkstMVDJDFcG60Svf
9Z7tAUwubDOEYmnTQAnSOJljDmFwdItLxx/D5rv6zuIqzg0tZxkzbvRgkwde/foJ
GfonJo41d0Ctbb06n7zUhRf7Dd4zTb0vSNjokEB5fj1ea9SHgbP1txPHY/xctZhv
JIjN0omb+HBQhaHg5Y+mJpFNT0KfAB1GGYnjQqJIwjR4+WwzLj89XDxF/NKXUUeL
4g1ytkrgAK1Fcn8Dx0aKFEgqF8LJ0NJ/v0t7sgyjr9+VrAO8hylZ2tSOKGzOjeu1
XW+Uhdnc5zik/eJXCorKgwOz7ECDkdPDrszSzeLFgYeRHS6KE7m2MnQ1NgUCWPTB
FIa+RJYhcL2JqZtaHz+blCS7ZURbRuDZSFAGogBmfwbBoWQ/n1KUmhgxyfMUZCaw
6ypv0Npu9mxpfPzGLhhUCw0dVsN3zowwYXxO/2Q9OnbTOsgWVosfqD0ZpQpQVNVG
2uFzZC8Z+FNqM48pvqpk5vkMR2gzqP4KCwxEzADAlYffiIAAscbJqxOtc7luO0zv
Enxa3VB9ct0/IvLK2vYObAHwcJl03gDpBR6aJ17Kt/UsvmYyLRVRjBvWGaM0fcK5
cOm7EkE9avPBGHL2I84Wc+E+gPZnzfGIO+4jDnGSZbfJba8iV80TjLlFf1dYvuFz
qsSSoL03PICwBBUnXqrLHUlqkvX6CoFcmFSxoFFMoQmYgwNreHex5gqkVFPJzaj2
z8K7X5R94X3Ji6FlsYqvm2sKoq9TCRqvDYoYL1mb9l3JG3CdllJE245u/H4FSmc2
QFR4Tc4ngSWarHPr7v7aDDk30Inl7Ks9Bfh637NT1AL79BCCjvVV4ZHtEDmrLlGp
Qt/7O8baQKiRUMuAv8khrlRPXyTYMHoZ3FSDD2NSZ4r/nRUq03U3NVuxqSD9YlL6
xryczgjnB8B0B7bYIodrYINhG2D8Cf2yBRmgh5Gm406LnRAyRPDdInTc6CNYLG2y
MYhI2MxOocd2cS6xMNBHYwT5nwN210dnDFVPpalEQdzSAQbaBkoSG2C9fM86lmWH
KKMSo+/gMV5vZX4+ZeUOCjWxfpvXuZiLA7SDF8gNwYa6sG+5lFk/JN26qAK8hR0K
pbytLEKqu0HegQbqRrL1ben1N1Mztj3VX9P0Lwo3vuxTRXESsFvD8arH4Tyvgr63
ndHFFAxTm+aRj/Mwo22lMALxJS8DlPLXk2lDpoMhX8H5ZAKjlaKUPvuaPRoLcMiF
P3OyIisQ/TchKSG80PVsMQrVpJ5fMi6tUU9wy0yVcCU92oQbpDWgBfgVrmHnyU6F
Wdx0PcESaO7wkYM0YPM7QvwWv9w10+sN3TpYPusgDBB2Qo6QGFyqjzimOSEs/WO3
S05b2u2fpcl32IMX4RHrtGo42WjbNx6n0D3I7Umb6gXh0B4F+K5x2fkAnFk0iryl
mFlcjd43yBlcIwuX1T4JKgL/jaTDl1D0XvNDg4QWwDg67MgDr/6aqwkb7XXYlV5y
J/TL8i12exyWctCMEH7dezOtRCG+UGnePNRRhYBnUOH4HQ/ZzAiqGxTOaBB1IZyI
/chXBX4wt/cH/xaNVCZExu3eJaXi6FvCQE0BGiEqrwbILI+twAthWH/RYGOKO0Y+
EcWQRnBpPlYurq082n3hsr/G/7SNxshe/DNm03hMsCDh2pY0iCgyx51wr/V9scz3
EAm38AA0gHycTjS3wlsf7cxClZaHYeZ2z0ONvZWg4HPSTVsfhzHc08Ok2tx4C4tV
sqFlz5vPGU+3EJrG+vAG7rbfw3LCyapR3T8amKUqUwpQEf3C4IsFYBVcDdddb+oH
diAZfbS9xhixcwJ4AR0CHvxS4dMZ/ou7EvuStaP+DzaHEHr98Wq7DOEOjHPeLT4r
1+MZq5gqpe9VcyIF0jUsFtWAWTEh7d/OGBtvosPx4b7VbFFgsTnf4frlYsaE7qCW
J9rY+/r8fgInDD4R8GdnkEF5GogZFJqvEWQ87yUl35YWHpsZLoHpPjRWInrfQQUH
XHXDEY69JYusRpS8KXVrxRMVKscMHDaF4C6KT3hLEdxdX7iEGGqbKN3lbONYG8eI
E8VEVXHd9v2tUS3kSyEJLGSQ9yuEDHRXb6821NzS/dzJOl4WFkZjDL3xNVc3N16B
Nvk1i9k7GDSkkdudws83bhhlJkTAIDYI5PxnkMijPNNhMY4zoXGmMs3aku2D4SaB
GOs56WmZqmH2mwvJdt006Uw2pa4Nn1nd47OgbX4FuS4lUeMSYBueR/7SAfzay8fL
FxHRXKTdArz0cm4SeoSCkwACkojY7pRTod5pxcNMQcIm720S4KoTLVh0LPNABBbF
KFZWzNLwJ7ZXRBP207Scbr0cXMMyPdGsdj6wxgJ9ppcp6mhzifoAtfjyybdOSSU7
WgUAQglVrZbKl+bYt1FROh4ffPtvcEl66vfou94VLhEHAS+gBNG3fG+ShMlKGq/D
xios3onTAv/CIHQzeIhZxgRAkfWYjKWOngNMp+ssUUpP/UyKwaMxNQJX/fbOdL+/
guBTDiKYeVh7+0lL/GAfYnMcw9DwRgWpU5s6BoNcZeEGi1rvvrdF/N5KhYJ83t1i
pOg1/d431wScFfNOA8TwGVyeZAkuG+2RNRddv410YwZTdWTX4slKBhMAv+9TlGBO
ZobltOjV1QNZsMPxCa2qi33w+63ngj/C38CQCn0R6n+Hc/QmfakXdPvvdO1FQ16F
R8vD+xBB0fFYSzsPud5mYN2X2Ep8kh6hparpO50THNdlgYUx85H0ncaP8o7nM4Il
WeaSwti66MjsNmjxbH2XAxvMI4zvIH7BQkbPs7tevUMxnmLHBWFntNbDHx+w9+4o
2k2yS4bH33X56YHiO/hpIyY/tXjHYRlCyhVuudG7fzYom6pf8/HnDOcWLyhsXwOk
uee4sJZPNR1tTw/P/88Km9hGgeBdyV8NKDThfbP1zVmf+s864iukay5fnpZp+xnM
NAfCpbXbqZ2YGARKPAqlSjlIRES2dfww3T5JgtcsfUz82lwSs1WI0i2fWOOe1UbI
crwQ4jk+fpjaeRYUM9XTcI6F5m7Jd/N5n8+c8U4Hn0r94ZrG70mEDohOuJSbS8op
EqVlyyCceNyqxxrYtDlzPGjIGClUGPF9LykTM0YptGxDCGfH0X4uoJpH9kbURMm0
ldozKTU/r3vqG0qYTLGjPY4K72sUz2kvvMH/Enw/Y4u4ojbWYAjdZYU4QJBMZQEU
YLg20aazaaM772nSJ7fwTLz4Oc8zYQ9FbRIEoXCo52EjCtA+m5Uo39qW6RWOw7vq
vWVMQx7mlRCqW4esZnzaSnvfA8901xXQs/RA69zVW3+O/jT0EGQwBQSKiXu3g9c4
TM3+8TtjHEx3OCIEEJLjzd4R17lJtbxWz6jMBySXNkkO7VYlYPh1CJgObOeTlC+5
5PlO+ZvmAwEO3L+MuHKH4gJaNjSTabxr11dDgp4uR86NBMGKYe0gcUc0Qfcjbxd+
0FCwS3E488xTrSMEk+XuKW8/XN7aeaCxZGgQl+yWHcRW/51kxiNoXmAr7YXOGQSY
KSOrKRpgG4cAR72dkz9ffnjDUQrOTAjQFtiX7RaO+KR02EucTIfStVFaccVFPFoU
BSl8P1sM/wr+29bkXtgwFy7TGmO7fB6QNKGUOKaqj+S+tmgb+8EnhrqvAEDqVqGf
2u92C7vh9O+4VVbhyv4Cf46pYhHXWf02bSw8pd2ecCox7ecbXAZu8JI7Z+eXZisL
0FB4b+EtZOiL9rJitNQdeAfRnOkyoz0zdq4IERY3J/SBNazaRxrkFwGitXeQF9ed
4Px9lMo+YefCrBo68Z52x5dAa9wQlrwHhmbwXxnL9Fc8dGVVJ37Xr8A6j3Ppun5i
7w9Jg4ialDXo1qlRRM1dI1w5xgITutZcIM4sZoH6JuHybyhA9zYFKjLv8EL5AVQX
sInfcAeIm0aj9IJpujPtNf4UDRL6kH4VIgNQ6XjFohARHfZPGNhOmHOpcEI/nWBn
NBz6bLCk9LMcUXMIGMkLwvDrgaykLvHfDHl5k0ULRE2yrfsOfY5UiqhM5xnACpir
DEZo3/BxpGINZxX0eAgHMJD9x1Vnp62mm+pXgmmJcRZdo2XTjJUbVC1e2tHGHxrh
pI3ytt3Ub8lOL3xyn16XGo4GDCjGvuSErasFRVSYHjAXrTrS78WFERQAKsu89ZRo
Bm8JH5PYMAJLZnaypIIfF9LSWI1nLexqzeQSn8qymeRvpcgdtU4ZWE0QUokaP6Oa
Gy30evBO68tyFgcpdWNsmialv8YdZ7yijUpIymuhovbcEmYe2Vxeijkt3tNsvylT
Io5P0tqSaJyIPaVS3LbuOxXXCWI5aAv9RFpKP0MwwnzVTY05WGGfHpPVejb84/o/
TgSLdBN86qjEdW5ascvWtOQTnZ6YCzomNWcw3kQ58wn1nceMNJzzOBm9XoSnhYbi
rx/8VbLaO40ZP7ee+f/CxgJA2+aY7A2lB1vuyTtmdMWY0aLK+40GTDgIkFRY7gWQ
+4QMPknTIsHFtSvcKY22ExcXz4BPnav8PBDi0MaglAyg56xD8Zq8ubzoddT+oveO
7OeCJg2JhZTAlNOeX2DfGdw6lYlKW7ZzEf0yaFKWe/G5Ogetq065Z32HeYULBFWB
P1pB2sNKJSvgC16dS0Ivqw7k3v0qgRfUEA/rFx163m1QevEpC+dU4x53aljTjnLG
dJDgDQ+LikQHmMHZwV+LMONn1KOYLA5SjfWC4XYb0IsqxrVVNv6JIGlRBWeat65w
sRtvLuGVorXvxWlgcFrPEvtqwkMLr6X+0kmE9E7ZYO5OaAPPjZ7hqnO9UAjnmopi
txKpb1XLsTLBwK+tNh+THk7rImdYc2123bkCqhU7nGEcXvNgKUqrn3r1/jjbNZdx
urRWStgLVFTeki64f8pfFSIHdVoMUkXCQnYfKFdwPKODK66c012RzZgp7LHYCdsJ
5PEST9L6gfxTsJUgtil8Ek2CtrSYb29xPWBqTgpeqJk48dHWbFuqIfuwq7rA72d9
0B1mqcfTEJZdisVoBJKCBqf/IXLSVJmxpNCmb/6q3LBgG1JJo+o5phsztLglaimd
SXvsZcY5udOmJZ7iue2X3BuNOr+zkIgFd3tNO4Hds5VE7e1N8bGNmJY+V3feyL9p
A+fZAGNxsG0B7x7VkKDOqRL8vDqredsxBBb10YCUXJ0xtLmK7LQJLCcxHSGUPrMK
ZEqxHxPOQnyFhJGofIyqxFQPp4SAUAjjG8uX82p9fp8HHFeBDbhQYZxwxyzTz3Ef
u7dFLHhXGWWZtollkpu4xcd8bMrZVhsPG7HxTh91MDMYdwa7eGElpw343Hx3gS2J
ZleM1xxOe/sYMaRAK9t3aeWbr+JWjkzVud9ooRJx9z4GHguNTXAxd5vhmS9ojEp3
ZlT+vU7zLo5EKuG8PDgIt8Hpljeq1Px63e5ucVQ7MKSgjKk8Txylg0+s5zPPPSjc
jp8Uk5ba3LlyVzl9qQooBo80pWjHJW1rPbp+rsdRiHl4wfm5cCuld9EqThO3Y4nX
IRo4YmEFDi1+u21l5y9JwGu+H5fqOk+UQUMFG3UFGnZblZrwOPqKscFFq8G5ziKw
ARjbakBUTz0nbl+77xZW/Boh3LXkFzgF+3uBpal/MjSDOgdb1/v0r5rDA2C8diNx
yZfLYkqykzPCMAeXImaircKNbaPXxI2Ac3LyNY39YHCHPPGFd9Iw7QU8m5bXz/W4
Zx04DcjerJmuuf1KiG+qHujYNaPTfIX7Ub+niAv0biwsq7L4G3JluiZFRs8RDN9z
yDRol+DKmH46uN5kzGWN43vcu5yZI1R/rm5hjIf/AoRHS9qNJ56dbDhVh486ai3P
qH+iEk78FTaTY+3uSC5//PgJ0NnyvoMnSmhVt4e+KFvCTFSQY/ZhVmzy2IrHNBC7
VQMDWi6ktuqQmWpjFVmwVVKUR8PQj9tMoStWOpjVieDepGcLB+fe4BxCGztshG+j
DyIQS84naLM68Q1Mp30RSuSI6+h6fTpAIGfujQNFlALEyd4cgUg8SqtvXWQHx839
Wa+xg5hIixc32PPxhAx9jWZRlBBrZn6Mx1hTmMQEak8d1cn2uopSNR3/xULh+uCP
JMtwAFL811FaMR8k+FYNM7VfuGheYcRWg2xQk75AT11QQ3yWFDP+StRnVG2bHmku
E/nAYJGuX1BvUCzeNfG3tHBvYij3W02pQj3LBioRWSz9Rp7AYibIg4//k5tLNa5j
DlWjh4Q2TsWyBoVqxaRpp3g1hJwfKGYmJaZVv3w4fd7gcSz4KVNWwj9C+lBoEqFE
JaXkbJpo3xW3u8VCyArUAB05tLlPsH56DyxByGnx1k4P598h3qrQFsC42A8HhQbd
DnY2fu4ljKcvuWB1Y69yRB8Y5C/z0oMymhIkmgWFFigkVubjOjqvmWctwnGwaGwj
wYyDP1gNp+vuqCy1LB9XFAhZHpKF3qdwrOR8NQ7ijCtfJO3HU7BgXr4YkFX8GLIF
qeRWJVrThmXBN7CcH+pChCAtear8X37TsRUOzrHFJSH09QFF+FJjM3KiVq05IvqK
9ksVmtkAO/SauV7mq+X/Oc5GPcIycYraanjUSz+jOWuRbH/5upy3y+cD4wkORPWL
1wdL3MYtOlQOhvRPAoCrqflbYG3cR6pOQff5LUeHAuVc3EiuZhcnrXgxNKzvLpMG
4MosnXY8hbK//wdOn/1kyFeghZlt/yf4eGazuBvq6FIIVL85Ki6xtbiTWmFQAw5O
Q7RKBsLK+/Sd1RNrxwC6YZ46mrrnPnrM0hMkXq5BncrVLM0dgZoMtXma/QB+Mcrk
p0y/lDm6RRMWC8U1mwfS6+nOGejqIYorN54QuGCMC2OWp1VAQ0PoNbf6O54DdK9H
nCet0BhmrNaZnbDyIvhwE2aWr0qLT+nAIXydw2a3vVPzj6KObm1C3KMZv7QHUhot
z1dOXDv3SJLA6kEqB8VD+uygCmYSItPUk4oR5+MG0ecYuNCH2BOst8zZgdZrQWjM
tX26JHsJbn9KMssNo0Czom5RF/RwMGxQ6DTSbBeFeig8dN+YqV61qKjtsQeONLkm
haK2Upu6ija2o234IWf36mZ6L0ur/TQlf+j4Ns2di2q9eu3x9i2LO2u/xCIPT+Vy
VJC8PBF1NqiVnZq/IG2cNuTeqSyZxHsuWYq3UVkoAfxl8nILA8OR74kZ7DdBehGf
8OfeZ4XgR3pfNDDkpgL/hzsSTe63J2tOo4x0lGHYREY2uHENFe9kioU0hZ7LxjWg
ZjD/520Ya98f8Z2cIV40n14s+lzSFigeAAU4V9s1Q3ot+P/v0WlPhKivWQ0EfdpL
JHaMk7/5DLcE+QfbgsPowlUqbq3V+wb0qKHVUvhdwjVraSYEUvaQKs/blyT0DOEn
0rEJQYwEHUxZPb5W0SvcuG8R1C91KlP5isNwQCMVuyG+0lT1IfiL0Tzm7o+DqaHt
cN/DTICB2veoP1mGaR4S5TvhfsUEynFE4m57xBlGKH/DDG66xnRg8TPX5m0ay8dG
1/rAw47s5LTDgCPmv8KVz8bzFPql02Sp4oi6aJz/6WDeyzjiuhNdDNLPxBb0Fcww
21a3Q+p50XpZ10H3w7wnamFMa5t/fvbpcfQuDXkAHEaXlbBA2UNPW03Dw15q+xNp
gkwXrx44W7lsjZuJsaZ9wTwfo7QLkRfEFN85hmmyg86vzqa5B6N1oWd7CzZVFppi
QaOMzmoW2vvt8zcBEGS1ZEZTU/XpxD5jYc48KrPEgobA+5mrPSIaLZvMarQUQE5/
bjauSlvE05qD5f5l8WOMRwrcjUJMP3GZuYOtv2VWrgRvj/AnJYSXx8A32J6eVgUS
N4v0Xl3gwmkqYrPyFi6aIuwoLhNjRr8I7n6em1wketyV0VKzG0IW6i3fFrDoqwrB
cAF8vXkIpP3rPIw6zMLE6nckSCclvB+S16A6+PEc/W+bEdqTyg28b9THaf6IRoHv
UboETB1UE+vvGryG9ckPKlo7tmu8meuigjTj5uS4rYcDFlwsr19gZjB92bdQexrh
44eM8clyJsvBN4Uggz4ELn+Z/4Tp4zP7Dw4RViBhgWUia2bEAARGEbFEa1of+dSQ
Vs1nrFcPYg1SVtjrG6sg5ZiXFBfUNfAnhcUHZ+hWqqVtLjyIfM9FaU8GbFPwR+uc
4VHHP6glUB/6GrS33WUFeTAldKpe/npxdo0ySpchr4iGpPX5sTMFFaA6aQtvCMw2
Wo5ciS7xlAKCtQvoa1N9ZjH4IPUW/bszTYGLdablDtxPY2le1+USwcNIZCVXfepB
WAHhRYWMyEHRUC8gikFsVy4AqtJfnL0LNTDGLIaZK8VUsHHBHZjGj6DZwNn0T23R
mhpoKCMte2EnedJazyH6bMWO1u8ud5G8NA5DeSz7Ts1DHR6E2H4Qp6+1O/BcAsUg
B54miRV6pd7vbF0wcDiDN5t/Hv+SQrNU/VMIU3+qdz0gFnQLAF+tss6Qc4jpSksV
DHFyCpXUMeLSV3Ae6+U/uxsng89mwCVgSbUu6DFhw9JfPTIkHXCdkUov0nSFACSJ
lVn2pi7JBHhLelqof5OdBg192WiEkFIsIon2LgDn+rbLav0E6xzEiWouAZnqrQSY
K5tC5M/D6fw5qAXTNUCa9M0kVGMrP+x2M6+0TVoxCeQzX89e6yxsl0Jy302djnnU
pjYPZfIrl57K/rtEWoPInsSs3k5OIHai+QFNsXDdYPn3Gf1x+WqNn6Y1IpfHP1KC
YkYSDuJT4/oCt2ArCwx6WqDyM5IHErEOlRgSIgz3KvdTA/5OZY/jcj2Q+bSFqT+x
PHzNUNcStKcL5xGjkSx7ckIp5/NQRUIpyU9MtLYYjIhMUsOstRkfb15ARBtG0M4l
R7UfGe6vdcxDN93IsR1E1ex9Y0NPgDoKPDxZaLfDldTPo5XvySw+OfbPuToEGoXT
xxJ1tNDaISyY7QZ0ju7Q6dy9Z0GMGURvxuGjcao8rubG95CZzK3FR9CLl5P6G+TZ
4U84wJltE+HIIoQ76GZz3DhqFCoJ4rrIn0uBi3jRyV30Uz6Ak2Jegcr0BknzPB4o
Cf9nFDZ6PKWeAz2DY1lWaMWiVVpRuopYCDM+/9VXQJh/LdQXNQTf1ggz8uWD6JH6
5l6/sy+AHlgx6GpGX5qHPp555aHzKwdf5fWSvyGIvySWHyANfFBiNJ4RmI2Qunws
LoTVCqVu+zIMF+/oTTRUy67vBoqE6k6ygPrBNwSrH+PnG8FvdxFmSRqpIcxEB98q
uyYWlvcp1gEuMauZD0n8YgiDAOEuG94joyvg7AYE7BCEkeioj6nw5SQGfUn7OUUD
6EwByKRn11Puhl1lCIwOknpPpTRe9JDb+KP0ia5BQjMOgcZgIuKhF0x7XfFl8eSK
7AfolheHnkHElujc35qPsYVmLigag5o+AvTtxZFTjmNxM8ElsxW9b0bBvwJyuZiJ
tUj0iCpCLqDRVIhcqM8rQs5PjqBAQY0VUnbGRAPnct8xrzxJqlLf0dqdc5J+1hdC
EN3mZd+lTbqTp7fPQKWY4bQbc45t1L8tudN++JOPkZrcH44e2EMwCnXjt3oCLSKW
1IcgksWJhTcdwhv2vy1Ju8B7+z3SulbE4S9wjo92pkJXIUn+6wHbGo0xRtGCcr7n
HRu0YgZct9jyvJNzcmkoGPks0ZOOBeq3Ej+gmLojvqpKTmO2BWx61uxSchiWIMRS
qiBuZvcwNVPL0X/F043oFyYZ6VowMICzNS5d2x9tIxMNTX1e0rg3zLIU59SWBwic
5BEgHuZC4JI+GJWs/xRJ0snNmc5m/QrBNbY8Ca4NXD5KhfROzcCXbSs5EztlOogL
Gsrvyu42ym9t5QFDrhtQDH/fYRiQJailSnkIjox7BkE4nmC/QvFQR/p+dNuOhxy1
aNue6UJMPT6RqWoO9aVWlR6xoxS7Hev+sTZYN6YDBh+uHgC25fkOwA1FUpUEjfiO
5kEP1vLE7+0Yr/FFZnC5uMwEtI8ckRFJe5jeB9pHcj/XGvkEAQCMqTSyrWvmvzFI
Ehv0Ko/HrLoDq0vHZWW8P27MQJNswKFw/PZpdac+Q7HjzCU0NHfyhMNlGvMpnxqd
w1HDOrcCfGl82LOJHCmY50trOBkQoqSCAY7swEsJrb1CqYXSWrgM4ZHr0TqkqW9V
b5nx0EWO7lu9H56DTa1BKmxEhMGOyoL1+/o0wdzztVqaLK0J+3tJKcgX8ciHowN+
AlMdwgUUfpsDq3eCrsWpUMI8s4S2zN23fs1U0SWCkYOw1nQqOhuJKnX1W569jE0Q
OGfNRkZMayFw/5CgSY3+5pUmvIPuvRy1OXC2t+MVWLNo2ZvzqsxSp7IPZfFeHVZd
EniLPiRSRMJO5MPmiTa7hdA1Uxqggmt4D7kVyve/wx/RXQBzzcDq3uWEov/Fc+/i
wwnKfBy7w+hJmjYnnZLqAQOJx7or7fwiuYhU9fzM+MyR0WHDC32nrwT3H5R4U57a
pSCkOe/sduzSYAWbzNmqqsqCtPlfblK7MG6qhhWPih4yoQ2pZlOGn4Mqjq6shWMP
Rdu8WMJG43W5FG/zXTV3jWjrScUq5dRuXwG/cExTHZPbbt6Go/Y7ecJCGxjf+UeW
IB3YxKfcfL+xaydaO+B7sCnE6ZWnt0cPrFjef56NEN/tTd+AxRd+aygs0v8kPOFQ
6GYjMEmXBrzdlXCbPWjeSUEfuKk/anseeR5KZLuVyq4J9iwa6D1/hKJCr1gJnKDq
4TXjlDxopz3xkSrwQ2iLHpnld8MMgeZ/7fnBNLvlkvnHtrum//ZjtexRJfBTqj+D
gFtmoQvABdd7Q0Om3Nu0Vi1JAhNAVKawGG06m/1y3etwod4rTIrKUhuBlyJEnKr5
Ml+vBsn/rR/DKUKppm8DPDBfTCI8K7dUCr+5Hw8HkRngUlxx6BfqFl7aX3pKFSBT
QKPpVfS1QjeRomSqmPje2nd3XIi23rZXZ7SDTMFiPaD+jegwi6k+j/N4RjB/Mmrr
xZs2wnHSQ6w8xvHCGAfiaEVO1LMh/xynZ+glFLUfhM0JPVd47i4OAMtG8D7fTilc
DBlq44q+7nEarDhGmmqXt2ZhtBhFdPdoWyW0CO6p7XgC4pqexfAZpjq3mJsU04UT
SUBfn8iKTYo9+1JGijhgstLi6x76Ec5fL9uyyuTnZTmdhPEhelzW7Q6WWsnRsLQ3
yGCQQBQV+3ABiVZjG36YzAh3gCsfJ5+u0xPeUDLAPiIA9IjufkllRnYp6MzyjGW0
kKAJM3CWv5fx5OKCrY9G1GO/BvdhtFZ+2Dd187GyGU4iyUSygSdTXKCYVGux7Nrp
9tWBsTNsZQcYTS7QZbEGQBqGUHNThTn8SqfXNvrAcieVRyfBtfmiXMJ6Ps4K3O9s
pru5Z/YbSAF+562cAcKg/zy+jcEr9eSI1Q9kgTn8jo7zVH0PzDrajYxNtAsA46te
mlQ0t/eLtFJlqhNH4fEoZ/lHyWx/AJfRXpSeCR6pZjjai4eHaJ+wcMpXEql5hdnb
8MiRs4XH1gJS9D8RPPYGPXyYvtyEJEcLalAmhZqkJ+WEBIYPYwCeK8vgNFSPBq25
VHJBydopmB8fDcizOWZOF8nqM2CrWSqpPdSrTZfaAc1Ma76qNfeid3IvsyV+VlKc
CPtzqSAXDzkiaD+vvltwvdiF47cTMhLHK+hAhPbv3709QPyZP1IrG0AfTiWBr5h+
xpnlzl2J6bnx0WmxyIX/L19oXT0IUKuteYdAWvmhHVlkaW2PIVoI4btDHbMY8+z4
eFxxwwL324lAHK8IZI/cREK9naq7CJfJmQ/WNhwXD5RfqmLWFFIzTadLkchbXveq
jZ1A23aFnHtMG4edTFD9YOTAtKMDGzASQxvM7JwQ2mU5YAEg8ByvELvUFWNjgvTu
EtU7CSDqx9g665CSia3MvCT0ozvulQr2SPidavmkA748SgyH14qeMMSzAeP88W/I
33Ac5zm4vs7VmNlKUEuZA0nTUUrDmOgAnqOi4xfEjbQgxD8ve6fFE+DggLGF4vlr
0elpeMaQq0TWrcLQt6Ee0HcHBgbW5fk3MjFuQoII1VKB3qps4Bae4ryQJ3MeYWGU
BTINJ2rY1xwEANCt4MkAMMzHOUvlJ8jshn3dcyFuC8dtKSDCMCHzH9B04zdjCaNg
zNcbEn5VoF1lfBmPOQkDqQI8D3i/zzXoRSnCHYiEJgYmlAvcGDBeueO/xK5K4PNs
Obv6Vt/okU7P27ojQcDXs7z0QON6NBUhQkb4NxSv8as/hbObPVMFt3qYhueK/ZQO
wb9xih4Hz5dlkPriSYrowSZ/dH5fkIVrNqDIYF1YSeuAEclcw9GeZ9qfJL9zTpfL
ItNtx3kNbSlfT6W4et2ypkaJpfcz9sbbVVmwH5gzzTdwBNt81Flbp/+fdV6sS5a6
KQzlnlfbWy+PSJsPAsY82RPptrBrVzHu4QzN/FxB/QdwsUW92jabFWyqpfhIlpI6
QfK+tE2U6xWc5m7x7NPGp35nAl6LmZyMhEbnq3xt6zlnpJBe9tW5B8M7LM0szJ17
qTSUSRSOLjlL7rs0Fih/UG+xKmFfjReKZQQeax3lMR8Bi6xxS17Z831ViJtNmRHn
Tdg+FjAVewddoxxfPDBLLogGAGs4cmMgvnTlHodSx0rINIypvybXjuMpZDqz4suP
2+CvsIqaO/49+FcvRauMArqnAFEau5DR0lE595sNr62c1pcicg+r9nWK2b5mSkRK
wIX/G4CdfrzegaApxuV8wVP+JzTW+QNiockujyD392N0hpAxrk2rSOc1Uv1TOAfA
e439l0SmXg75HE/YnaRsbsZ598qt5R+xwnVevYZDOjAs80UbPrk6etHj96zApywQ
vp7ppgmn0DqHDJb25e7Pvf05fCTIwpw5qkuXyqTtIyyKlLRwwKU+txJIVSsgtIgQ
zUZD2Mxqr+lSfiFpUDyf/WZwGgQmtrFaRmuY7ycA4c04ZJVD0BnhwDOkd5NrlO1V
wQctxdRq9ki+2A0azleko3DjgptyWuz8vtU421CGanV8Uh5DMcZjW2P1NSUWRdhE
pnnDizOF7/rdPNSMCzFvluCzPvb7ol2LBrXXJMppMpOdPVKAxpxIJ3D/izJf57ll
wGDrXToLmKipRAzq5gDhgRHIjEzFbud2tnZvA34HblKe/oMhZbS/knHy1wnr5mRf
qSTDrptCXMLlaV4shRkiWIU0ZEm9UgMF2I9IB7iOeg7ovQDH3OF1tIMpOk1C3b0t
35MMJBS+qHT3hJtQKjhg0b7WdVeXLyI2eiHa/KYyVu5B+zcZ7TZNaWJXJhpL2qzv
6mkfB/ngaU4OyzvWTEJgJzTqCk8xLgpc24mTHI1oMXQ3qQQoXwr0PVda4ZdbhlYs
/X7yamYmasSSsuHLpbZlDlHtWnpN2QHM1wqUq6dYfC5jME+iD82hRQgFumLdbFRF
5yHv+NWBeMgfQYThMxLG1uNXChoDTYPd/lDMdy3WMnFgl509TS5XlFOo4/IkFDuK
97Plan+4f468DOqDGzb6ltV1iv7Qyn0i8BvjLqLhV5dHIAjjhE4y9221ybeEkz12
pNifucUboZ8fOvFM7lz3s36yDvE6b8PU3JVbWMQJaoDP9bG5ciZtxW2hI+kta2+4
Xjl0IGruP1iKVAVck0ENlRGmCwKNpqwn1BB7pS9hptMhfkWEWYS+MD0gdSZHvzTH
I3IOHa4vOzZoKVTOuGE7y60m2ninH6qtWAAqHS3TABfOPhrjhZFVUTSWljbrVY1/
uD8n9yaZbgedktKErSv2/tIGBX5ZxMAVAnbqzS/lVbRIY6gDm93Vy9tlR22tjypg
HYQ1yesUI6D5k30UouwmFcwtOe3s56mpf83qfV2vhkkCPqpBB3QTPmTVvTTYjeM5
Ak2Nv5w+mAQfhtYBRVrT4I73akifXv4SXDQLrQFcxwuSE8Ydb9Y+IP8puKu8und6
5E0rw4A8ogsiXMLhTD34Zb9rVv7fx8JFGEpe+mpwRFJ2p5PYlYwVY0LRmjfYfsWb
lrFGM2VIIbj08bYjtH9aVAKJw3ev3xYJoykV8ARDwkjgnavYN7LSrCH9mBb6loFY
9DwBQvNZgJxXlm5JlgcwyBsA5Xlq2FpwBbl8lWhcU6seCT8cMsWGohVFd6uVGbsa
I+3Wpf5+xjlq6dLOzSmO+oZBDtccSw5jmLobIZ/BAYTGkmyZw6D1vTvUjZSiKsH5
LpYoWm8hu+S+VFUKhNwa6iTngTY0rQ9eUab+8B0h+tPgbW194s4CfFdWF3ua5Ol2
SySZG/YKn3L45dvVbzlAoJhl3vSH9ycwz4dowZvyLstqfz5+0//fIj+JFwWm2+H9
X/b9z2UWH6MOYf8gS3TuO/P3lZjYuRCOdo8r5X/6Ho7U3OhxLk4Sj3rPWElCb8jz
FmxV9mMiYKd9e5h8XFcMuKJm7S3/uuxBSPebW+u5G3px+LZ/PAc9yLEe7oI/nfoS
fQJtiiT6N7lmd4fNua+kbOVYggO0kdlUiupqYnwcPIx07uv2o1+KFUxz+lF46l4F
Ob8Wqoh3+X+csvrUVseiGzBo/lvtiRAcVrYypyJ0hQD23ZIOkIuNZNrMJzN78KH1
omAcBzFhB91JOpijxvrfFqE62NStYA9giyF12o0YvKsV9WBZ26FPVGK0I2BGUlcA
UnW5oFfr/qVTPEdTuKHzS1SEDn64F+95jdbVvtmow0I8YRdHFXUKmErM6twvM+fW
FlXFV7NT5ufPLFK7LJKF+zmXB5miLQ97bS8MB4tdY3heiNzxu/+klbkQO/uKOOn6
VBr/yYT/y/5udTSjNINtWRXynaBr9ipbXOFOTCwr4d2xx2WOogO/tlE3Av9Fwp1t
ZlsvYKq6qzR6z4j7fLax1DQ1FReFBZ04762kRHmwXCTJhmeZW6gCWpA5VtV59Blf
2th3Rs/BrJ0WoMeguCR3F4xRw2p3jYgxD9kZtZUl/Ms26DsiiGTVAw2vyzQ5Zf5d
03MKzMw+D2qRSlW0yTNR85ONkzyUxncaI8WE3FadI8n9RiSY7+qXc6d8QAytPHa+
H5ffoSXJDRXtRxeGd0PXCyX92ohulRMC9YqLf1Vfasg/iC+EQXwAnhP3uRRqc2E1
bJKi1VUHZrERxRNC/KnUKHSylIWThPLEGNdVSxRD3dMZCcFlvAwNeUfJMlbuOMMD
kDdBEq1tihlP4vmwOjdYI4J3r2n3nQRDjeLkf7ZXsYWYKCW6O69gi8rRS3x1Ebj7
YaEJsKqhWd6v6XPmdE+/iR1s5+HKgJPlxi333zptpYyOkyHwDlqfVv8enjC8qX+x
FIJSgknBtM4MlalTCLqZVo4VhYujWHG0Z4Vm3ml4xQqOh0KQBOFi1Vd5ePqiUb9P
2tmH2w5eFhRUmMi8E5nMWYPHq3B1c5NWK14nIveWkxaUuTdymLzg4pvppf2z7PqC
fv7IbhXtMh4liQwIvJnaKq0ltnr+KcnxUcRtgrXJB4OgVZFbdhAYhHZ/kB5z2YWZ
Wh5j7Nz4J/EiNro3xZ7ONCS1HpeI+1mugm0e2VZn74jf3/zADSE1oxPOqBSs4uj3
/7U9Mfj00y28m+Xx+Fj1Qsis2+Lb6lDVTdpgeBYE79qADLrcVU4iFS/HKS9lSqqb
n2KdWFldBgKZOPP3ETUbwF1w8iuycSjlhP5bD6crYpkpYtC2Z4cbdLjFJiBZPMCp
7OSIREv4JD7X67jJ1hMfiQfpMIvsaZ6ZmNaLSa/IA9NemqUAoYr2V4RJlcPtZv1H
7swJ7FXSWu1HJZyuNzoWJ/xTmpmUeG270bbsQfCpYCL72CwlJM41vJHV0fAJV2XT
gvFQkjqMhfhCyRJmKtXGfB62If2oFTmRIgzUoQ+J08cwVWg4Iuz4g12ThcXYUZ/L
o2ku0W/kK2gGDhd+CjKN6SSd5yo1lyLaPkJqxgigcuNxeWoVP94+KWDVxbUjcivA
tTj2PMevzrFJoqJpR+q3NngOGHFkT1begrRarvL6mXwnGvWAQFe+ViKiYxkCybx3
SB18y16oMcOTNpTod7tkvDn5XUrL9qp8ibkrZroNA0xqn1QJQGpsdaLuQp7y63cB
xV7pB7ZJ7nCXfHgKvLsmshfSLSbto8E2rcI42YEfdeArni7HqGUYHn9h1fiIcqJ8
3hbJ0b0jYtNI/qMXgsPgqO6C9DQfPgwQ8fTHzbKiyDn60hG3ngrxmRImaWEX5Pjx
Qh+RJs8zliy8OEtImOW4xTmo91aOBeB34o7JULKqQhrp36nxGifGkF4i1AntKS9D
5ZE6qSQH33HzESP6v/noYFOUcnGfFm/jEmcEm5wejwxB4sIypmaitVncLc7Y7DUt
0V83KbIu4jMsT6RiPXV4nU0+QQoXEUIU9OXgapHTB+w3oa2aXmI/ifL23yoAhdNp
M+11rw11Q9AJe/NvuL0ejhBOAGKfXQkff7B0SRvyWiHL02Z6RTY7sLEwYDctpSp4
zhJkwSyr2saT0ymdowIb6eFGguhAxg4OZzmasmFG0mkjdlweOA+T10f+nCLimss4
DJoonGCsQNK3eRcUCNhkVqhzfWY4M00OfFHXv2woElKHMHG+bQNS5ysmoj8gzxs8
F6tnXgjpaj2i1wKmWOzYVdgrAEOnj1wkzsSDFSGWHioG+xpOeFZbVqqXhtsUiTDA
yieEYHHZXs/nVmQVpXck3wNNHd/Zcgt6mRz4u0L1l+tGtWXHAIVt4l4D4GoTCMI0
VDIhbkQE8JPr74bxlipgSzb328m6UdMXV9+NpPZOLkypHSxkVz90XaNHut2k67UQ
PT/YSnvyTDeN/A4RmsVQuxKNTseQGn8vJt6iPUtJtcqWIgy3DiJG0nSQdwf1p8nm
eDBJLdq/tcDXlU00b/ECThrsjaD9fIOwPWlyqPl43y6Y0zcQmc+UT0lyKOI2TEFv
nqhi9L+dBr1WMAoke//BP2qWwSdzY9JnMnqCy0hGOYA6Vc2fEdSB5c7218vUL8K4
Kj+Cg7IbQqCaO7TITSasvlKX6sBg4vnQoOFdK2+zn5T3XxrRqj8HvMYF2Fy+mBfO
cnIxFbniiAUb/U5IIyjN14cvEx/mlIm1wtB6Pgf0FPCZqSch8lbubJB8zuD1W4Uo
fXdD6xprV6fBQNSFH3I2W3xpf0h0I+izD9NT3cbahxxSjPwthKz9xSr6PAZO9fpc
ZCQ2YJbOatSPYktWuAm8L9UBs+xTIOh8OpZO1WSc7leGehpjJAQxDCikNrnigTNm
P8d6cXv/ejj9MldcBSX3/nPjTral1So0uU4w/eIXshe0PdaxyCYkHzjiDxdMaA9a
vWRBs51X4I4hLBLNjbF5MuvGGfRLC+kwv+Vq0URSWSENPLwwB32Z8on53h96GDLj
RC5I305mmHPY972VHQQYzOB+OUQsB1BUqFKJTSJ+g/NCQjVK8pQL/VjMHEMlxD+U
tWn4eHKlC5L0MqofNbKJzMEXgkiWhbX/BfoJbVQ9wb5LB+d+8gfOSYZCzCj9isW7
29qJ9yYBKrSUNSagqppZMymMtk2li0i1qNjQsIsMuzd7V0piSZTKV6m+d/atPX9S
mlKXXrks4PAWdDKzMtBY/cayYNHGGXoNSWJC9zZalag9/f9VtJuI+I2xQCnB/YM2
TUHPiFlGlmpFmwO0g9IQMoqOUAJfZ1WvgKwbaDzVmB5hYYUnM4CodvxU+M4S6ouT
+THiaoKQS43t7vzNcaSCpGrKDto+KA4XvZi8KwosLWHN8zP1ZSFX6GEIPIOSzBUX
L6dsaFRiFr3N9ui3O5twr3DqVRT4rqjt8iAW56w3UN5UKHe/eHuzl+s1l16EdYcO
IutjmurlN5J1opdb1mW4mYAmeuLNx+EOYTIkINVTgu2ws2z7zGeJWyR6c4517zNb
jvaN4qRvsWBFXEAIr3MYTHJ14gvZABtELRATCdXVdd7jZTX7lMYFZ8gRJpMTzVbt
/y4pqyKWJSatKlNY1XSvjNjUFeuoTsm1/+hVIvMmGZEMxzd40b8Lcu27Qx/dYxk6
KWh3NnwsRDcYLsv35TuxzmwhovNFQB/+x2Qq3HtCW/IgL0OXd5+tPevDwjArkQTV
FXqVXXxXKIXhNmtGyMGvWwAY5sWFkQ2A6vTulT43QWukn7Zjwaw8c6i8zdojMYRe
oQpE85sbV8jih12yx6sOIq+Ql8YgOlGlWOs5kklUAc70TbtV/TGYUmZJpqEP56YC
GD5IAebeFV+N6jDFwa9c1OCiDjEOzHEFd07ghRHdMzxBVRkg1pyTGbxh2oPFlZ6n
agwG7SoHGVdaBLXNMddrxcksuE/TXvinA/GXXYkDYRXWGTXy4d81FKde4+h/vhC6
dbt9Ge9EyYdw43EZC3tAkp9JLfxfLArxp+dCqU1Unzna25N1p9PKNsFUFyv6jV0E
xpq/9lDfSyRdHhW7L6ANSgTkw2ufN2YI7kJ1YUZVN3Dfqm+4BBRQ3jxAFxZdbnyX
rr0Iss0EjnMy24NIMYR6e4k9qgCSW8y74mvaIhNx/2ICg1xjQxCZNN6NiZpKdnjk
us7+piV6oeAGO17wrNnbCFGB2AW9rGQmGcjhMus97PDdON4pNKTRISJu1sI8qIAQ
HFjExruw9iPxvytH28KW3LqzkUTKwr1OgvP1dMFeuMJVuXQq2/01NwC4BE9bQE3a
bm75UWgKSB7hEfjEBhWzHcQahbBVGqFO8fIf7F5+C1xHDs9wawYYUmlpooSpWzVg
DUl/cZUCsgMZIxPoNCsi/lrVgVlBjDwf1vl4i/5/qzKCgrwYnbh4BIBDRX3Y49Sj
hIVGWpz6qdemARUm0z1iJNbGoxCBtkHyukOmZbR9eBmpiCMwmXcfuoyk3SqT66Sa
gAKuaqujBA4u02IoLvbyOYwj9WfEGTTeHNLM4xj/apAwITaoaWD/njBMKzFtcDQ+
n5hJwn19ifDRCcDrRA8tg/Jf624PN/3oBQJKQL2PiF5M3C6ZAy8R6TVyCmuaFOWt
43jWOzkn+39QlWmynN4RpHMnFK8xl8WmNYlrOMCHjTZ54uSUR3csTF9WLxV2J+rE
AijoM91aG12eVSI/l/tRUFB9sJ9GoM2DQNObZWPIEfYsogY1YyvyYKNgbWtqDKuK
ceD6a2FOQOI9UUbZAZ3FO2t4sOiXOEG+KQw0EWsVqKJRafZlvd4dT7vKBZMLJv/k
E/jduMht2U4A9g7HMX/SV0ZrbdkJCgoprwTijc01AFNeIy5wpy/LgfJMVZx3mCc2
F+QyzWZwqz0IznZJZdYUW0120s0bMg3Dt7XMW6q6FI/b1+Yw2YaVKnMTMgwzJnfR
yyY2uXPrfGyYviMfzkDUe2zQzypjjjRXbQ7fNX976x83R3Nq6LEs2ck6W69r8oRA
TuiJjcVASpqyq1TgBFEgxdaQWDrxF3CEKd2U/QCKOL31lfHSIAwmyGLZC5Ej2Yli
R5OLl2GNqXaKJtqMkBHnpzH1y3RuYgtk5xsOTkPB36CbtH0SEUUQy5keNhUF5qez
kn60hDXfmn8qDh9VuY84/+skyxfHZLMs97r0AXFCWm1fCf48MOmA6WRxJ0Lr0a2p
M0gQxZhiuu0HvlIF5Z7aVTaKkkgCI20477o0dmyftNW0Iq/DYp/Woa4ZbjC/4F4B
p69MEEbmZT33YTXBEkUMyS/vMUaBTh/9NYBc0obHuamauzfN27PKGs7Kjmv7vEsu
Qs23zAz2nptfF1SPg61ti7ZJmyeZ12o5qVRrNwZJreAdiuhCp9iNDt3FbA7bjIxq
91xvCQo4if/V+v9ewIAFX+JhfqNQoEz5lUcPtLXWTcxMb0DEReJwBOTGmYt2/TkK
ecvr4D0neh42d9QcdaS+U771bNlC3CNfKgjVGVu2wn9qz2vk+hQWG/pDpia+NS62
w4L2B6ou/cVQQB94XaL4zkX5pivrCLd9qyUBWVT4FZz5e39BJYiztqJw/vEUFoV+
TjQpBPJhRQsU0lyohcCvg3D0ajNa4okzUJn3P+zejmndgEpZ1EfpOHWzAYxwKcPX
K/gDcK7mjg43JIcsbGFv3pShJn0G8uXHgragePnS/aPe9k7s2VGX/VGFzda2oG0f
CyXyH6XMsd+YflO50+6UM7bSNG2PbiFemWCoNNwOdpD2vDB0QtpF+3YD48i/Ba+C
+ZToo8ZdfH6mAQwD1h4Qj+WPZzKxpMl5Rp5vCkHGDWfQ/DGprj8FM7EMt1F2am0B
Kd82Q9ueS1vwHlpCrLZ/9ZI0BEqFEsu1hPh6YSXsm3j9LjfD5b6PmVmeVfF/OLaE
QhnAOdyNrHGy1sklhI60NZM2vfhTmuU9Z3BaXsW/R1EiYb8OyEqTm9ZLAJ3ueVOE
+AO1R1Ki9CDhbQvg15yzM7KwskLwLjEhZXVqMSSXpky8K6jlmbnXJK5VFoHpI4QI
h5DN9nhKxp2IUB0YGi42C6LPCwpYDfFCTDkegaMKBI6784dca0wjlvpWqtJKAxGj
Xm5Kxw3NmqXv2y3dY059jO82urBchSFq838q8pULStyPfGl61FrjlrXC5dpq3IAq
WmjhPfHEzGOQFZ+mBxTvPhzCpUuZk2ao3eIryFl9J5l3vEXdZNAlJsNmZG+KteDM
BspxSoXhAtbQ3z7bG6Y0xueXFg3c4VvhOZpeb6YLWCc09pOBrx1O0BLyneS9C5jw
LIMx402vDhRvMpjBpSsQ+K+9r79ASp4018BjdzipuyEBo+WRTLFFgENV7X5M4tBO
ISk1y5tIZYNn0qk7eZi5cor2Gp/rSHPBhys7gNUmDFi/QKlKM+eM/ab8+MdR5O0n
xZ4Lc5mxgpM3OBSNfAOwa8toZAg5k2yPt138NWalG8czMJHMyL8DrBbvlqheNTrB
O7r1H+uJ65U/7GkQJc7i/iqqoXlcNnpKxSWJBamY6FOzucA9S/fX1IlX8nCyyxHS
PKiavH0G0dicI9TO374a/kTpB65Gtqhes5bfT+zJncLJvkrvVj+kK1gbEPuPOlr0
Zw+y+Sgb7Fomc2ht7Ese97340bXIUdllY/VO6Mn/IkaTSc79N16ByIoLN3Cjk8N5
40nm3XDNU2sNUOmmjEqspIYxJXyvmZKQs3S/Nk8vjTeldz2aucpi0A3ROGhs1NZu
Qk1p55KfvrAU84CJFuWdfgQLdPt4a22comoWGFUcadE3Bo5T3JwMoHTM4L9CRy3z
YQGB7EA9nknk8qM+pRuPbFIdXb9TjRGcZWLRqLRF1b+6vYKQUBy5YD8MulzEpbhB
OLDoEzW2OITK8MN7fhBeP5dh/pK2CPBUPrnbzsZnzb1IDFI8F09JwEB3mWyCIZ+8
iV7biMuZz9qgrcv4zWo4IfkZtQovA+dtb71rJmXIZYGHdbee236MwuIjheMRttwP
3o0cp/r81a4H8/smxgqzl/yxYABzHwh4tGw7zUQAMSUO8tnpAxG2/9XENAtsnbuu
77xbzcn+zXEuDbdJbwllmQQwAV1pJObuqegz1iUf5axcXttLr4v4FC5dXSZZNRHX
Ao68lAQVB87pwYise/pNC3LbNYur9sZ39visFOCId2kKOm2M8OG/HouBIiOa9h6c
ZPI4A0Rok+YddPoqhQJtTAcUPWSlzsGIzBrty7b5tBFiCricb9DIpnphU1x21dXm
J8cS7PLGHcnFdMm7OdxmF2vGTXlfTEovI42qR7wZ9CMISxY1BLZXottmoyeYUpTM
Y6mDr9DSkyUvsdCPsEPmRKKGhKQaGc06gUCVs1UYqEd+gEZ0yUZMWWO8lVtywNaV
MjxGVq66F98PKhq2g/04wBDShHyolcXvpXJH1uqaQ8o88ClzsDbqyKJ6U8/3CxXk
U8uXKfYAPjvL8p8Kz1vfyK87yeV2931+4YFFrPoxl5Gp9bjoEg+6r4LQYptv29Hu
7l9KxsXj2PiXw2GJO70B6FDDbw7p4QeH4SLpaIHQyA7FrV68gqClOi13DrAXYcPT
uwjClV+jOp0pRx3dXVMy/KNdC5/4NN4d/a+ExkU4NZjKkz9MNzR2VY5fVV3YK7W8
lnw2L6kTFVYQ+5gc6xnVf1uRX4kansB+tXe72LOaQi9rZG+uh4V2DipcpH5+Yaqs
GFUdcsRxr0GCHADs+u3Y+26abDttCsP91YDQXc/EN4NwPFqeWwCys9vOTQV+1nN4
Tg4pKQmKE3D5krKzM1T/yyoAxH0P7foiZTitiwnXWw/FApIJc3gds3vYsGzLBy/Y
275ImPTji4oGuCYASOWmBvwc66nTrzHopv2fYmrBzADMLXo8C4f7MW+qDHUEFPMC
yvY4ZYsZIjJWvpF0yhZER+gB0vfmS68lprj5v4YbP0NOzH4zIxR1KBH0KU6LvkLY
q8xI4eS0YeUMeRkuiRBuk8XTFrueLm1BlxLaFGs738HVClYEm3WU4tY9CHLQ948l
aHudGrDMEWDCAAwlkFtFI432kFWUZWTtIu87oGZV0KLTjBSDTSNYcVARgJfhrkg9
8U5ktos+osJuSqQZhqdafQnlnonwl17IG5JYxlh8vQDLfnEhk2GsSLxIXULvoM2J
WzrJ8Tyf2Rg8mRckCbL70Pkd0xye8DjAhePSahk67UB0uvck80ncsPsjavV2qpsr
JGTk9ie9z1yJO+gAvwIXYH87+dQHZXOgx9lT5nIxgQvdkN17HurSXALcqd1BfMn3
9rJCLGnydU7JW4NtDy4seKSjCZTM68MJ4tcrX74cmHVQF2gLYQIz7vf8ydVGWBcd
lYTpHRO1LCC4Bu+2zPYp0kxNU9nzuZc0hGW9biQBmIzPfVuAyuX43dzcEZ28o5ks
EXk7pOU6sP4AaO1ilkDCXEJ2O75kTH0Nn0HVNAYKZC+Qf8eIH7SajSl0x+7aJzoa
riLiS5eHaejwFxIKVoTfv4S7ybPcvsuRyY0KvXn8WkogpCk2afiVFu+KUnOQyiTr
rxg/jzgC36C/7oMCuBOYnNpBrgkX9rsiVAkiODPXOPdvlbQBGYgVD9cbm9tL18NN
MWfMJhMXt7BqN05yh5Jk8b27Wh0tPKCyhBg4oc4qDd+1E11pbUxIydbkwrNuAsRZ
ZfczL/5wVeKeCl1sgyOg7ShnYb1ne3hg7XIV+RLflZHmoDQ3Fl7b/6/i2EAP2SNN
wJ/juoZZA4qB07f9m7k4emsdOQN1pvUaCvklOb/pM8tk5pashhghFqCcF+6LGuTq
hAcXJBO6sl7nTGc4an5ai0wAV7VG5iCFelJNxEvowJvkkz/hU01+tCJ1ULmSjRJn
+ZFugHSX5j45cddnMA5ZsC5KpVd6uxSyzpDJkYPwubpg4aECnx6vyvdND18w7hPf
rPjmujrzkOoLgf6cgsnz3jCrkUxOZrkYgn2s05H0hoFPLVbYO3o1YcH/uBHWpIga
scmf5hDv/Our/IMnH7GW8LObBh/Z6T5/iSw4LM4kMW/JWn/rpjS/4Jy5Vge7JgHA
PQMS+fDWMU6S6IZjG56qfIqlizVflHpRNiL5XxS+fwpc23O0xu0oSshEQj2hS4Jw
Py9S6JmwxBvnW2pILzc9v2w8wPXAfEznIkMln4OcgChNzMzGfrJW47PFu+7Ic4KO
SJrwsJy56m/nH8KC7ncwSjarWmLnZJXMmJa2hsE5N5SBbNmNynuHePJ7Lca0lPzZ
7AtOMkPz5apnlYt/fb78MA7t4g4UzjOsKMZpZy/3EhkPulM0KmGWptah/4kMsbEU
YckArRmVCAghhoiHjq0FR070rQU5g2G50Ybg2Y/Nsd4+NKaTfgmCDUJILI8skGCh
vlUFim3X5dOo0hco+kerU3sRDErWNl3d8ZKz8TQkmbWMGmOK9wjMhEXuV0lNU/VW
M1NL/Y3PF11TB0ycpmTYKzQSaJY4AkRb/piSuohEsj79COkIR2kfhQLQOOjrbYAA
IpKLtwECvn/h1VAqpRtKV7oyRfGqkzd1cpFUEvZeXEA7Idk5X50PKJFrxCpPlq5z
O2Oy14y8MyM0cdQSPun6JSpte6HIPsVAkUONBwn9aV40UW58TQ930B0PUC2OVqma
u4EPBuFWD79NUh9jD5D446pNVeIIvVdZ8cxk6X8TjEPLntrfPXZj56jOCFp3cpCX
Rw7/XIgZUPNW0sm6D23wn8nuLBbZx3qXF76Cc2V51SPiTZcHF01VzgL8ccJownOi
g7VS5CzJbhlxPns0q7D9KQUYqAX3MlH3HKToYOx0KE191ZbZ22slhD8+D6QfM8Bt
C+wTBxUujkPipND/PuTv/kXtCGo+ghIEwvww7dRjWYCMPoxvkwpor6QrhPwdnoMg
wKLWkh7KaASPdLnINefzkSCNM48af68EK6htsNWrNBt6VcAL8/hWEz/8b2fshuW4
ZeTEoN7j8bdl3xJWiDhm638F9nyLVLx9YhsWcRze9QA1mVjkI48AocDoteJPb7mB
mjW2m3Ra3EMa9Z19XN6MJ37W0TBNNVkYgPwsxnQ0M6RBh55ea57O3AwmwZRHwpIk
l8PruGZ+h8YEzWNiDUAAGAlNmwdOogYwsDMfOiCltv5ZLig6GogrrXl7cyO5CBtt
N5h/4Hyn6fbGl/wbdMT6vXbuE2Ppd+GfoNzJYkLkh2uvnbL4qix4QYIDGnA6cKRf
fT0rGNcGg3XZKikPDvY80dak3vyzkIJ8wzEAwOtMnPvtEsDgja4xB3h24kuJ9dUK
0bYnKNLpMtHZglo2qVOAOUpGdcxt2PFAWjd094HNr5uC7AhaaSA/PVAnyNrHaPqF
cqt+AHu+0sRXaGiz0B6YUx7Otb4i30yNbHOYYTytYrHPbMay3A299+lcLurPLN/v
gfQ7nGuS1hkMng2HrhYKRBcirnTGFXgETeoJ9IpHpJWJ7FPKnSUiulMMygmLeFeD
MpXipQJ+F0p8GDZKhevG2NzTJ/oyRskANiduRdF/CthwqRjXBXvd26Z+V2ve+UUu
cqBJjIKAMB7yceLmcjuseqmWRJUd0nX8fuWRiLqXjNVzR7EwZ7X3edCVPql7NfWp
BuG5v6KBEiaMEdwx24K2VQ3dH7h1ehl1XJDxQSLCYn0q/uIdT6sCsnga0Q0RFrZ7
cRhR8hbaGVj+i1NapJtGpYVFA5sQtOPfL9rDCMlgymx0hp+51nGOeVCP663jcr2D
htT4RZ9STCcUbbtGTda6LBSSm6qmnJZ77TR8gclDv3C67vOwYEmVkgR5t7KWOQuz
+v4vR/oWzEVkJY5JBvJgdumFY83ZKM1rDkDIytxmrzVOCQw937V6FOJiCvGoWdBR
MuOkCNC/RpCEIi5pV8vU15dbTGZG8ukbNZe7UTUS2oq6XmZ6rIeYfWclfNR9iL3y
qY2tWxLqJ7Yy/7diLHcQKXBDWb/bXx6HnYfSYrexZ7r6MaK6dTvra2K6juIHYdLx
2QA30vsx52/YMJ+S8v9idaUK4gzkJgsvQI4k90kKbbREWazu8ZBZBYY8LJbj17S1
7hms4onfcZhpHUEeh7JsfHjsk4ukIWKKDY6aGF8MPAaM/XOI+MCUGVXijCl8FyJx
UCFTls9cMK++2tqeWf6LGVfVKwnqPn/meYoY5E2j2lX0D8i9GbqQUgj/1o/W/miG
hQxTt7Lnp6fjT57pcf5P4VR1eVSATbn/7am/5XQsd5RpYacp7bxtEH7xLscT/+DH
0IjV0zzWkjLpIXzbkxk8nPACZUkFYSJPvBg6pXm569EDTrQN6kBdOY85WhuknQud
3j/gfhBUn8pe80WQwbAiXUzovmDJAWnBG3uvcSKq6d4oFHEWi9bbVbrdDFFWe0bM
iNaCE9DsoDQEOZpBnpPUrawP+gqFcY92ZX808ESxb/jXC+LYT4hiLDqpVkMa/6P0
Ddq8DXNdDnsFT+6OAQ2u8qmWpV0gkqT0Pr89sFeWmboe7eCZ3vK5SVryLpIg6Qd3
nlHlPIioXDPuI6kMKLEFealWXF6D7ZoKovyQvBStZelh4iPCZad1kAjfjrVoy6rU
c/+ik9+Rkiw4g/8EwAz9Tx2G8AgBvX+HU+S9A1+IGOmofKC/FZVeNWPTVoQaDp5z
HivIXbYEbZ+i5/LUf3goWJ1hNXL6h2QNjsqDdd0YhuBD2Ls95NqnuIkrCU//XpQg
EVvatEmAkhjkrc4wU3RY2xT10wRy86S3otyerNmGm8c3Wo1DdVetC/LaO7Jf6Nai
9F+w8xAuSvhjQ1uxQ99usQx8tBVY0mxR5BalJhXlGKYHBg75GpP29yvFcOKBs3sZ
rUgw0WcNsN3aT64V1fLYiq5X4Sk1QpeZaEmnfplMrQ8B5vH+auaDLwKrMNoBsl90
ilD8rUnCN8WmezpCdM8cgdIZtW11yEnYrwoYnNOWODrvZjbsAhDPSK4/IXK4vmYP
AKr4duhmWTjCxbRbT/J6bACqy7OBZv9HkiwfqShczzd8CaIxcWazn0a8mKefTiNX
fXg+Z06zYog1pFLW04vPbpLrp4Igrqe4Z2xePtIdFOn25AQSmOkA1fNB9OWCA2Q+
PBVBaEq1bRPhADDAIf+sGbwgNjbRR7q7HcOvNcphcRk/XUJf+X8XK87fFpX5BN2i
2m6zIIX8CtGCDsMA0Icj156bZ7aNHmbPn9XoUH7CUYttRY5MJR5XndLDWbKACptx
mXDWpbqpBf3i1xBFTAUH+p3jJ5ISfjEbWq1ruJxwhjhvCM2MdfCLVbU9hZbx8+Ho
Ivw+qxGDcJ+4mfMhJiN98ecG61oOfH/68vIRKQ8hGl8sztddh70fWy95W9qXzcx8
gy0Qmhq8EIT3YsqKJAoSKMaYDP2kbT0drXUGvZQib2NQ4o2yAVoHWU33wdKwdXR8
NM8nFlqo99JtoI0uIRULj8HyaxRrsEebw5A+GyXlKuFImSXDhOWAHsaS0iMn1WTt
Gsu+QqKwQw+CKpouUzQ9P8vCNcNDTatxaWM1gMpIBcU7NnFU6PFwKn3KSsYKEBPP
bOec5+/UrvxjJbP/bYaS66h9xZOG7mv9+3da90QgX+P/hh7pbXnkkO1efdfG4NF7
fS/4Ub9aybfZbahDtKIhH/QqMYnNNRp+1zTi/usr1uROTdr0mtxX2qRoZ5zJav7/
geZq97YIRCJjkwvu5u/3I0pPo/34yW+pmaFJhwJrzWHnTZNTftJKQ06EGFf+ym+H
vKyvPpqjkKnYCoNmeSS/Mftx4BWNY78DYm75xWJQcgJH0hJzuBj8nd/2vHZ8FhDV
mXKX4geALdEjNQqgYa8JL/8FL0nC3imYyCPc3ynRkAGpvaXzsNNAzcZOO7WF7rkm
m5w3OzikuB08bjFN4eVnEp/vvBhNSh0J8NxIoI5G7bO8T4g01fcW6A0CAGI8x5ly
ADO8q04wU7tQV3CFI0Rc6UNo71NsiK17l400rMqVNCgUuQRDnx6v2cDjy1llHxzO
0a2RVAdoudCDxnSc7x26bLprNhrUx83CMPlCKmKt8iHqH+xhMWTYS0T1yAh9rWP9
9hxQ+rKNL34rgYkM9xj7KMCpjpO+kjmJPBiIc4ZKHDZ3rNtZGPO18z5LEcjN0ooU
0avHwlNvy7VRkpfmGFgM26i8q5HmtHa1NmuzEob7AdF2tvwpfv+kSC9/7a1+6jiV
4pWS9OdMxds5bbr2JVyCLju5EldVyfFl08lMlEo80+U+r5ptBD/pA6eoNjX3x2ar
KkYdIwvldCApIUxoukPxmCdK/pMXMk3XjHBD4l+eSq+kxrxx42C27nLe7C4+0cTP
Kk85sHWZx5MpwjJ/n/ZehJUp42K/M5u6qu+d6gk5nDTKtaiYYiAm7o350qHq/6ZL
Z5zYCwUFQm2wmT3mefU4yZx17tx1dRvI9ji6huqK2vBIRZIATbGY89L70ynw4B7Y
Q/YX4FtVDAIdu+Y56ppkUPlrmbh0y6WOTTsOqhwamp9qHvctil164/qj0Cf+5EFI
rIX0WtNCJwtzW9hBVj/2xYZCJ/5mTYLZiWGaC6lORXzOcLXW3d9BCD2fxoIeW9p+
0qTF6CF1DbNLqjErral1td4lXQZob6eeWjdbijWMAawqZkMBuIEsNU9ZIGLD/RgC
r5doCv0VmsEdQXi2XzdUgJnBaigkxYTKBp6u7A2/QzXaMKm+sL7N/beVdx+moVev
sAvUynYN+OeJ7N9+4WD2LI/VaT/Bl+At1dZYzRk6K6YaPgA1g97nvnzu8k6Dvujj
BbfjSWtXa8x7QUp9J3YtZbM2aDv9/Yeugx2DlONI6uF/oey9PW1JpfpYUijQSLny
rm3rpXND0tt+RXLn8pi3j4GL4XkJFv3+cKuqXmhzZWvfMMCbeZQ3eETcS7tIZ/mq
H0DQKSGliWwmPGrg9ldVisx7/lTRiZO9N+rl3PQ2vxjhN6vvUciHxJ9NKiw74Hbr
/SiGnc2nQ4jVp7CrFCF/pviBpl981TUa0jONUB5FKYtCcYWY/c45l+NHk9Jr7pAb
hXqBvICMK1YGSqW3U2flZfvYY4h6q/k287ESPgQQ5Avd5dwNhkWOoL7mOKfOFXD8
KO+VNvWP4dcs9y1nr8N5WbIYf8QYDhe0W672j3QvlWIrbuQHOgstelN4FrcaMTpd
agOCpklgL0Fa7S6SPs1bw3gD1dVeuIycYz4uz4YDqhG5jmFmtVdmEGhwiBGxKUjy
DkDZu2FZJMoyz7DTFyY7vudfkrmT4zyshM6OsmvIjfFWduEEjti+OsWaYC/cPDNS
3lw9sMl6MbEOwxDDL40ZgI/M31KrbfS/cObocQCU2ZJ6P2UcCWuy0BVRE5LyVULG
8EDDLhOPdDdTOKCrpKrxWFgkrTEuEIpuHD1nTF4VY6eWIKmQTcl2AGvDn93qRzcC
QWwb8lr3m2x2+xWyEF8KVNveiXVIK11jKtufJc+OvVwUItqY1QpJeLsTcpMaNlxW
NL+oyPy4FzBWjNl+zWnlK+4C6ORCQ161WXdEQCZ+qyVwJ/Mczyexeb0tFvIH8TCJ
6vVSdL1JJrXVIBB5NSzw9E2qzEX9Ka4kSjSUGdNErppYZ50zxX+fYbl/vf/gYb5l
Cpve2vruH7Z9dG6vVLngkenXUak5ze0MnMLIraCyBVvE7k+QYu6fLX30RWBOjYHQ
gAFzuk+R8NqRd3L3kylsbA7DiWrt7wOfkVIlTNe0VYr69/wFCr68XuMBZQOXEnsE
Eb2/Hq9gO/1NO++8y9F6BI0ZTArbYNrQRSZ0Sr/UCqmUYuMHu3lPY2EFGMMcjPQe
5WSiFrARuMW+T1zTYzsMnI8ANOLuj7LLCJKCeSZOnly7evoIwkEd0e6YeNOcF3gl
MUDONSOhx3p2kCn+iKa5pG/CaJjfaCZJfQks9UMsUW68fEJX7LsmV3KU2SButrYc
CKf5ujTDmiH3OzAfJCEuvqKsMkhQVMXM4pSv5VBA6SalpfELJEIohsacwukpQYdo
y5m7KCS2OzD+Vlc2Sxloh3iCkT4XVhVKfeoEDAZZn38c/tpd+ZFz/rOg5b+6qE+g
KEP1NngbmsMAHM0miIMujrLdGk57GjJRfj4+gyyTqIQHBFbbJ8yfem+dpFuUVd99
wCLHOi66MsXCgmDYcB3uD93nhQpmt2xGK28PUEpNF+o1+98XyK6xnqAGkL0gk3uo
3EX1fIvDxGKwlxF5AiYNK9TnFnYQXBxlisyz6x5Dr1fpk6hiLXLuEVGKjN6DSQ5Z
Ntolwtm2BLXlndsXcL/KKpVyMDagbDGl9W0OCqfUwNSvHF+yUEaNpyEwzEaZ8RUV
bV92MGALq4ye2tCmkm2eR0KiFk3boUb4Jas2pUpiKermhOgDPFMseWQUavlnBq3B
9LRdrIf9l07RLebPqtig1vM7qsYfY42Iql9NUMntQnxSwjxgHuLmyE84KcQiTmlW
afXUFqBtOXhd7JWnWemVcIzXOdgILnACT096rbGsoWYMMiUdfccv1rdEQgYCNvGr
mRGlUOM8NcSERdR+7W8jT7cPe/sz0Y3SIVuaaGDjvQtNZJYTipe1QFt9VFItJ3A8
OeX4HwcaC1ZJANLw3ExEuBXh7XwS5poVJfJ74lLN0LKse/Ji9T7snUJX/pGR8dZP
EqYepL0awGg51weplK4gN/vTvTEYGgcHcTbsKelHyhUv48TMkH/lrHD8WiOdH3Ow
UWDmm3h4IqGNtohrYjh21tbtqU85fG4MzetHXDnm4MkuZl0iAxYXc1nqFHEMFNVF
rCaAsefzleR6WKvfFIyG5wMzfudn7WU1b/dvufvpKs3DvRZ+UNzWzcxq9YuKi4kO
D0317bTdrzIJ1KCPGvosuc2tKt9otX6yMdMSUaCZme4TTPbsXAO7mB0ObUKJLThF
4EnJ+5mAEcxvhmZ8X/vp0bHFAK5TaCOET1UQ8wAila8PSvb+Lw29sCIcrLc2ktCI
zVSJmYBgpdRnsCpjuaeyaWUHu64wGlFJJostM/rHOBOlDH0zZRKzkdu2wz7W1yAL
z8HnInhZlkuiYvxeYllSOJAAI3ecBtxNsUlQ2mmO/120IyvrECtnNgqCu0i/IfjW
s6hBnRhV4InQ3Fga9nHyh1Qy1Jq+nqfQAy2TL6ujFS2j5eA9PRTrjZYNflqeap69
gZRTnKFkci+rgGzhpamOnkFDCPbxeNVPTtzQOCFgK1vzAYClR6hBACcLsL7Nqlnn
sgwxHjlcQ8fbz7AMKaPuR3qaSlNH9l6gTqbSxcNsgX15hsIESQfsBSMfowyNZTD1
CcZivgXB3YyUZUxjKTUU8jzmY8HxmLE1mvAlaKAjnKSuecE5jFb/BLjNr4/MeEO4
lYN4q+fQDMO+Yf7MqxYxTmbC1s78pNI8zkSz2rErkLAPd4DKq7Lnp7wAclsD/0Kd
cbMZRpP0FBMcZ/C/JJuCtClhPaeg5XeWUKu7b+RY5JHYfdZjQU5WUJxctNaMIwHu
Lwjo2CIT9PZDRvp42IQyypeK848KAOLzFbtfaHCeAf/ckWqMqgKHKNC07XQbauDr
l+hF5fsNTQuMRV7OO/lY63A5T6nUI84komFI3qQKvcBw8tz2Ojh1Z55npTKrwJRl
HKjY546QewSzkbt8reNJrP9HOgufe3ATyrPJw00qwK5FZDc9Fgu/miwTaAAxH8cd
+KCSCkrOKl9RtxLoB0v47lk5gTIrKzb25n6Smrogx3tQqa+L/Qw+1twqjeLCf58t
osOpipCHsU0OsdN+2l+kS+d4inWp/gyq/ycc+CZCaYwvuNpsYy1dRaOm2ukTKDmX
WAAFKKQP/lIaaj/nny1rl8OcaQj1arsWhQWDUOuD5Qs9NRm+q0QVSUMBy+rez2fb
O5d+ll8yREkMN+o+9OKNGTug1lVsNFZyI5v1RXz3WIJu1mDX+k4PhdAd7Uhj+Rbc
8Ha7XCaRY+NRDeOTkTx7dNF4GOfLbH7JrDpm/OS7CAdRUzMHajIvBNvlCn3JR5bl
mBQ0nG24NX6KcGQvE04uL9wpQU89QcB6x58ISElfG4JGlg/WBYkWy7llOgdfw13H
IVelfvGDHeXfaHz2XOjVTl3mhDEUKs7m4yinkZ3/gi3nNTrsZoH3+FiFLDQzhP2l
VkGdLK0f/JGqwzJlNY9/sQNZMcJ+0vWdm35XpxNa8PJ+vYi7+Y16sMCsO5mAyTWQ
eWLn87ZzgiQccRMVVxo8OOFNAx3IoSf/9A0OQjmJFNwE9ZByhmZb9iJvS9hF7hPG
6gwyYVysGyGoUcmsuDcpxP7Kr/877bXEhMgjpeLu5Nj5Syz7sg9qNZ3/hGkOX9yr
XLilztTdG1wl5GdmsliQuSitKGQ0vyzpQrqt0PQF/GNcwmLVsskp7zE2SkBEY3me
mY4SVPhXuwHvegwDSlygGLKdLja7Ijh3pn1erRsxdl7LcrTkH5RndaJC93oY/AOQ
yU7DwynAdhf8xvX9GrYzfOCcqpTSf2a8gZcNKd8ihDrFi3nwsgmCkQZqnmK7P3jA
LgGhJ+481c8O9noH+Fg0uDEhDNaVaoGaJ05tfGU/vOpJ/C62DgwUqbEUOBoi0Mwd
r0eg7xjqVfwUK9ffnDyL4915JBzeFndy3DgWT3HNG1vQVWoemjLYJ2at8M6Be0sf
Og3jDOpw49SRqq05AteSho4MeYC2pI2pX9qIJhLpSB+GsdtUfC1cjC4shd5+vssQ
FmQwgilhcjp5wr+DjRmTPeJhHQFjPQa2LQaclU7w4MZ5IclXYF4AQ6T/qjDA8gzs
BpjpHum1H3sGlkyG3LQLhvPXkR0DX46s08aH8Q82IkEHFW7poJa/mGxR/k/JBoIm
IOnNOlt1c+k65BK8wa9Bi6k+hhvhbYkbH3Zh9bn899EnX2oqrsz+bymHIHvV+yG8
InH52Bvi2AmMEo3r5WiYiUk4nT4Veos1l5ML1s5J5FAiDDWQ0v/xPglBfI8LztqM
omC2GruuaU9jLnCgLo58sCFwwW6XJAnOdvhH2OUuSnHbxgGmJEufmNxa1XZ9FUcL
43FBhC0NILz4KBUEs8fPQSKJYVvUo1JocY8pys9PiCfw969BzCpFjF8mNTDcneSQ
EMmfALs+zeUOrNCYajdfvb7M2wrkLjmIyrcpZgfe5IEx9bKmdqi98CgmkS3PZTOO
J5XPFNbK2/pZX/ySJDI+9piyDip4CloSEaDiPrQ57aK2JtgLs+oTVCvzIxn45fH9
8Qevx4QXJU2hHBBUxxVXBAjjYm4x5m7MR2QqcTjpde9CfLL8aEJ6OYC22zmbSGXg
GDIW5Gbqn6ljrW2XSTgzQP9ZtKh7yn5SedOuzbuKACsjIlbEM3yd1O79VTlAIttB
JsXEn1/7hoobF5AAp8XA8ne/GHpppmauI3fy3EZSswOEl41bV9zW+0O4UdBszcqy
zHtTdxppSz4PXHEezJL+SDYMXWyyXza6FbW2zKPD4dyaixJyH1pbuz1sMpFODjNY
KWgBIcF2oPQH5C6d86CIuILyuJgQpBnwywEybMuYwvoVbHLISAs+zLWPu6QRQGNr
xkJFGrOKXCjmC/4/5IfOxEHLMBZvUzxhOnyEnUhf8GgUSARt8+dwzIn7iF8SIt5a
JdjQyP3TGdaZtAOdK1PgGAIg4ZKX1CpwR7heLvxLojgZNCsDhSND/W8GHryuh0AT
gJilkOOgy6YlH6u73bNrNbJh9QRwc8z+qwLoBxY/UmkMPWne15Wkz+mMW6RtnQ0l
aKkh2wv3wmnLnEbhY5HcTkTr4r2Li/S5T0i3IKKtp+YUe0PIUSCZP7bGLX7oW71U
10CZXX739hgq9SZMEyU/VNyuyP1kYU1AiiqzYa4hb9RtYwFlEYksjLrP9VKsQZE5
OqP/ZaapY/BNXMvgiujLUn12AP3c4Mc0vzelExY1JOpVjhIDoPDuT2di9/XTnQeX
5siUSfV2+X6h3Nb2JDIXyMUVGmxURxEf8TOaN66SDpQYhw4RJxE7/pGPFXN1Bjna
nWFnUYYEpe8oyqbFYLzdELzovzNfai/Hn4GyYtF/s3O3BblU0g1VyH4279nV5618
CIih9h6qNX9i/t/NHoqL6l+RX8bYSopUlvmg3uOHK6BR2cFP44MPeodH7nvNVVgk
c6i8mj/l3R2xqf9bdvmCATEMoD2fI+dx03BAA1Xp6rf5KX/yvS32GmV5YOgPrULB
tIiqTtF8NnwnaaIQgn/QOhOgoKHQq+ZLq1DagALQMaxUsOjg8xqbwNHd3Qfkd7H3
UKIidRLPJVrLj81kc1T9swlWy8FP4lBo8n5obMIjbnCQk6X2wC4IrwqPpqTzx/ga
3ea3XTNet1bT9tb7tGHFFqvyDgvZDVFGnh7mO2lJGPvUeaJUryjE1Q6j8apsV0Ad
cbzBOr67QSWDQhMveJjzVbdMQ9wmYHYidL7Q+qc4aUScaQamOTixi5tPc7auoIQo
rEX8/KVZ1SQS0pNvsPvT+d2Xprfa4Yr3GkDLQxT5ddzpQyhsiq/6LAV/BnMI5Rtj
Qa650PIDj9PIBQVXEWdXlrdTo/sEta26GWn+XJRsIo4QNQyr9pV1yRuWcNn8SgAA
jSECDqebdKVjcnCPOkBVEhc/HBwZB9EjypBXlB/Osy6GMGbXyZ+od1d8gsfPXB6H
ewX5CtwpkQKuwXH1JtQrWzaeQdoc95+b8w+0sfu2x++Mf/E0RXiRAz1cBsGdfpeM
fYW0o4sfM/uXgHAlZVCM9ZSPzVLLMOsow3l0jygTR1l49Lz7bNnggdlNUZIhirpX
GRBxaFbvVn3UVp6fORWwA3FEOrdSxD64WS14kT64ipMEqIwMRWYXrF7CcWHW5+WO
XuuBDRYn5DJHcNwx6Q+6RBw7BL5UICA8/4R7zj5apRNwKPKm6eUaRzIuAiATyDOu
cAmUkH/CVlybCalkV84eRIs5KQ8hnzVcCCjz7q5sRdwy22naq+//vfdV/O23Do7J
CWXE+NaJ59YiI5tThUC1MC0qbBuG1SviQXhw+fG1/XcpA9Uih64FGSBbQGNHyrXO
QZxFwFZtNcub+QJt5DvWeUjnp6diVfBqs7tpuBGXnAB3Q1ktKFC6Rtms7kd+LMTX
GInuTRcwAJELeWeFUy82PlcHLFA6+xM/C7WFAICg7EBXUcl8QK4X2iDKYbL49IZI
7O3f+IAF6oa5iOuVCB9Pi4hmEblk0nT54Mi6xOT+ywRBL/hPFvloEi5lg93jFSD4
7+e0peDE12C/f5uUOj4traLVbYns4aQrBSi1fk8UuPRftL/ymuok+6jr2iIYl0DS
0Ym2AQHM/8WFux5xYAfMh+Q+APOo8Oy6+bhvVkh2gMlmGk7hsYi75OEnZ3p+QM39
HI4JE9zXvI+3WhPy1BpNLebzf+oip9pJko64qZtgD2/R1z5Y8vedNfQOivXLIr1i
gif1F7oz9wInfR6jHAdG4znh0FDZKwnr17FqsxqqmsXQkWdzirN5f1rLWYK9GkMr
6nSR/Nh3vVUpWaD1L2/nHfsWMVupVuq8r1RH4wEFIzM6frtWPtne3brQbCeskYof
XzEiXX5pB+Fwxkp12mzBz2bxJjn75agxh+hCCOpIi8WOkiKbeGuHAhRj1/zl3kRA
dQgky50GyzuO83qmLuYHUbidPz1FPh8AM9p9wjFkvujuM3HNh3FTanK0qxfNb2hd
LsbtN6+PvaH4V6Iu7PKVzBgN4z9j6K8Vlms+DUfzOvIWTRnaIbYT4+AtOYvY/TmB
m5PKefkLg5a0ojeD+AG3T8N/PYE4khdbKf//vhlbqWYDKsHfJ0fHMez+OBK/xMyv
4RYyBxwvff+r1mFsVzyxF4bmLjczELJXN4Rbal8lf1nsd8hVeSarjKWw6GMGE8dn
J3knj6eHTarS3Kef28nZQNHPtf9Qg07qMsLm9CRbBy6J3jpXU52L89vLn90M1h0J
AyO6KRGet2JWcMlW9L6kXaFYi5MwZk2T7Ibp1L5PRNkPOmvQvhFAXp/3hYNJcMmA
PKJ8tUB1NS2v8NUEDH+YddgfS1WX7YXNfMt6QyE0k7Qn9ojfvSNoqEhHqlaD1gxN
1gLpbdk1Nn3JZY4bekscX46AF0SLltJcbqHqdGYdCgYM6ZUUAp2BXw7PqXn9Q8vv
N1ffXc8wDlsv0ZNPshmz7aF377tv2TKsT4+ESIanVJaO1a3Wpna4uWW8SBtm4HFf
NVkffsQeTu9VfWHAp0bfOnQw2QPlqYXVWHk8EOsw+2YXDTw7vfI3PqL8cglOvTqV
ylfhwoxPQj1/6k26YrVX43MUbaN4JXgmW89FHBDQf9u4ZMGz20hH68dm2ZbLYBbh
IlGAexOECSQtvYXIv+bAxpSyxNZUog4oILLOXNtsX1KFviHanwcKAU9ULT7CkfZ5
YBwUqKQUpgcRGjp3UMmQv3r7lHdFCRPp/7h/10HNnAcvA8NIIAm4MR5xXbEawKlC
YUbmZpLJinE4jUc7jHBJ1sqF4A3diTdnDNJ7QZTiJtftvc2ZsVQbytAJQq++31nB
pzpTINUN98+cSbcC2ktpVnwr1lyfB5pw/oEMLVc3zQohmKo9np9w2zJSdhyomqYh
qvR+LDL2Z8f/XQB2Sy0jyFw1iTX8ZRlhRWCJMIU/52gHd+sE4s2YbYZRCmnOE1zI
JoOn/JD0/38sGxxF+8Cv7QsLakpi/0s+KdWloAvmdr68hUfbvYPiLVy/0+AMacxz
r/fQ6zSGjIn1LAeYEwRU1GgFpZTUOBgGQfZv00jwoj6rARsd0JYSsr8Q7sgp1Dnp
OPWiLh6sR3oUoJ/FeGC3t6Ylm4VjRkGbBFwGAI1marbE2HJfbpLR5TFQKrrx96R8
y8J4Nl7vcyIjdc7clRxlIfv745xSorjuICfQKoGuhnhhJscycD7uXef9rPeE4DDe
H+K7gWqliRdu8KxGylsXHaqc5ze0/B0LYbcTe4qwfSPjyAxDiM73RURmLrMczFrM
Xr0mJHobq9ySoSFmep1zQ4MGMvCLP7vXBeqkG7OMybOXahIfNHGcTynRWPjlg0c4
b9NDYyWMMu7+zw3BYH0SI0FhltuHtuk3Wp0cOd9Kvyg6Ao6lXuL3EecC85vVubp3
8aByQsNeAsmkFOkT4w/GooIKxkOzRRSjkfDZ++oHWcpa4PDVc6q+Gf1BGM5+kSW5
kj41UnTk+t4y7JcB5G8glkrro6BBlV8NmyWYgvmQU8XHCwh3XWdMmeD6vB2T43X9
wjh6qJVrVUtszurP0kQiwbbU5Qqe7tUZ3gjuDYHs2MgEBnEBn5UJR2qY0nUd1hUL
dqbI2V5zmXoaS3qjH2Q0QDiNuxpTaNZ5YYN+Gf0XCVwiaVAB5qZtvBrTkrASsR2o
/gPEs6dY4wjK5NEL6ivNW54uyYd57aNJ8aSZVn2pjh/+ZwXjziLJaSGjLVrWp4jA
CK5X0zkxmMapwNAT1WIr+d94p4pvUJlLwVUbya1XrhRw9fS4tLIuvRfunfq7RmPQ
+EpRCy2OUzGmFoQcygmxWokA6CCnzOuZnjnt+xsmO0hfu2yjkVdj9G/beeUzAcNG
0iYR+68PUwDeW5pUvxQxqjY06ENGTUZ3jgr8XQUg9TvZeDZIWv7T0zx4of5wS9Xk
NhaWJwVZM2llYzo1nUQ1xq5iy3F+pef4XOcmX7PYAGFDu/RhTLv4fTkQkkg+HLK6
O6l1IPebmNXPvhfKtiVWmyl85AipAs2WKdhKZLnmFnnVJwcQIl1q7baPe1gutIiU
9h4iEgOXKo4kQBwZ9u3RypuXRIzjOMbf+2WIN0k/FIi2vOvJ9LFVMPiX02axoTp2
kyR+GYu8X4b5142x41somUfeg7xq0HQgDUWCHztWA0SDm51rf/9l2fivQIGvvk3C
nt4pHHmWA/LNma+RUXcLFfy+vCOs+IkS+KIW2I4jjQvgMWsdvYS7TmB8VSLtvGBB
qGvTr+lYUdV8X6tmOl1kqpbWGchQoojcL5Dnotvs8l+2NQkc97RyXWxYTi/l2XUM
Iofn8RY4j/1YenFk4caAyttL17SBptVOf3u47utuyWhwAllUPwENr2q2ctTEoAnt
/RPdSrF9ewNX4Mbjsp/E7VXhXzl0OzbRguO/OysGzFWb4grdTZ396cY9tuoKdp9y
P0p3ZeZ2A11Negb0wZvjkGIENHLEYziC1Ek08Y6UvxuGwZP6/t4VasuXdrfsJ/oC
IgaL+hghjMWLLfogAxy1cCzQqyL4zgyx+4R20To3WuzLHzjAWn2LdlzXM4s/utOs
8D2Pf6QRgzMrowT3qackBun/hRAai5JWitxAKPi3T6DfGV1+lBAao5Ki2sUudgxi
GJIRE+iJFE+AV4WwHcStN43c0kfTjLAC0kXVo0gH1OzmzsH1VBPXnZwngIRAl+MO
v8LNf6L6AYZnUoQ9iK3LmSYics6QFId8gPfBrIYCaln3QUrqFaxiC+ZGyEtGDdul
pJdBZJxMq8L/f4Q+ykcRK9PshMy3XX07QodWg+MYBsrF1tg+W3upGyfIpuBzwfKv
z4aPKGNbW/pGLU2Mztuz6XM4d0v4lkZKe+cVyHw/dLS5MG7aUXVhW7yNSzBy0D6q
RGz6G2Ifi/atdvw6CpdEJuTKNI6JWhZsXy0WdSOjV7pSMyDbqx5LssElNTJ9UOK1
RycQWelbjgpAeRUCCaRKjiEzMKQNHlzxTCKlVKaN7zuWgQGUcl6FjbNx1wWDtWHm
k+cNbxV14KE/9lRHKu/BSd45JEAMdp7zkwrJoegoyu79tja9vQ+E+wDVu82YtBLs
d8AkFqg9vbHA8McKZTGQpHDgS22MMSiuaF6fm0xPzybkMMY+gAsJnQTBw196+KD7
wbZQLnJqDcZ4+xoJSsDyVSKUtUBY00jH9WdhRuDpFcNSWBJ9Rfr/ZHmOd7NhlcH0
NvFDyoi3xaIBtmb9MhyUEeQYlAEdV/ZOik3B8mfbMXi/EErSB8n2J2A1oFXRw3bw
k7+sbdfpNt/oZKPJAfq06J4BGcQEyg2Pvjndkehk3lBi7DMKtm/ksX7LG0QgoURv
Aasg2nsoggcRUOtfd+TKJyI2CCohyqJlECqvqOg8XHNqQ5crrhmYygaerTrVPECF
JpODmtiB9uzTLhQAa6ha5T4/95jFwWFhrawahsw2ROuX0jxy7DQbsb1p0s/Bd6m4
zzuvpmHD/Damc8+Leaq3K++QVzqmuxYRxK9oOFQX3Lr9j42tDyUY+Gzg79rD2AGK
awisYmm1DE2FOxLxfvklpatsh742frmoquUqvewJVDdx5JURVDFjDas+R1OmTcsQ
WBc0I49fXw1xF+Z30OSihUnERMEn4Wyz1mw1AKBFDCuwH1xim1NkVBvIKRPQu+S0
0T12+S82Ty+v+HKPTKMHaf5jL3iyn/PndoXGI4LjCOGSFpBPB5zbx9dCcrXkw+xU
P+eRdo0yxebuhIDeZoik5CqTGVxX3iRQPzsPE5s2FFcKEi9GcCwbS2kNRllNn3AN
p226uRqC5eNy/EctZ5RzFmXCLmu5LnObeM4sBGILifAsMuxP7IJnY3RK3heOAnDz
mpDakkw+i5kFXzqOAyncFPyWUgo7jIGb2VwmVj+rrfxt4vsLOS8957d92fIUIIzH
OV1MH9N0yrupcGUP1Bep+2L1UmEYRapeu5B1zblIjj3rBnp4XMyP/JWOA/DKYpBW
MYUHsJbXh7JKDQIctTTMYN64l5jqJVR/6J6P5YHwh9TiSHopS0VBNXtOrxCs6yj7
7xwsqlDL9hpnxfyJF7kNVip5FmQYUnrp65Wd8DJWem3wO704cJfnSAbkHvwO0fqp
4EPj1cuZYiXWfBcGrx7uQQM0kBfPxB8oi22Q1TS3fugtvNDcwbF58nMwyf9G1Rrb
/L05DCPdT969Je/giV3EPate8ovHqHqAWOgPU9dYFHo+ln/6pvFRBdEijrHTB/Aj
pjYVoVHOSXIVNxF7VhrSJgXiZgsm9rs1C6Ove/+xakfUkqxcXIahY5yGj+TVX9ov
Qiiob9JrG7cwjqnuiAmSzElZd+mtGW5riOd3SwLXIKWvMZNZ5cex7qMlQb65ctlx
zL3s50XnNVTK97X98wAqlrsYFhQL2qLEtXiSCJlJ8joSCcrtM4LCkyewv6qiC493
V9CazU+5zMBQpDqaTMZYhNElmEzU3q8a8aPwXijSu83sX4dnLoKOVln0goZZ+Oay
HNRNmgygG5v24KorA2UCWyxMqlMQavWJ5rA1dvreJcB8t16X+jBA0CkQkdoVVLct
OIfHeFMoIBhuKV2WGW7Ezm2JeQmiEQNaqTQ9+/GVdEAs1prk4H4/76mxqA3p7p36
FpstyoIzr8kLnPCZ95CbSt8eHj1xJHMuTkHJSU3VgewYbYB4LJBHyK+Imeps/5Pv
SYT132LrKOu2ju9rNLGZzzDAS/J3tbfdEBg4zGBajMi4zrycAnDnV0mr2tRUdMs9
v4GfINnDjqb/prGyTuwzX0RUeD8WY6mF2Vtan732YuGMSVjVgQFFEL9SD1847fr3
/qTNCNKCqdkOTg5dLNK9fwwJEmumOTxoCltcqboCRXdW18I3MAOawnAklN1fGPfQ
PEGN16r4DVjpl8QyQNsuEoAT7qzpsarGvjnJB+oD+gy1oLEgOy+OV8uW+VyzJ7Wq
4JU9F4zVyXly/9jBaqhF8B1yuI8bG+by55TFFk9I5lEfZH9Q7j/RRoJFNo8CIozx
kCQ14IU602p9C55KIfwpK+lzp3fSRNtS7nl33SVSibgsBq9tH9VGCnUQ55VBdsxx
/Bk0XW8uWn+2UQxbzVannXxRy19OwXM5izuR2bI8EJ88VJ/ta9C2YZ1mGBbUUPou
mbJzopxVbVTHCfqVQ95DnPM90JhhxZesm+ECC76US2nBlmcZwFIE2wlb5mtf0oS2
qTM8lDzwWbmQqGYhbVq6VEyrTKbZf//y396R3Q5TeIBYZWMoT8gCHrBdFF4y6iiN
fG8+HIkwSn4SnDCWdfIUr3a36NxKuwst4FhBP9RvEH0ItcSQ8vRWp5NeR/gSMnBm
uOYzBeWtxnUfvI4z0ST1KriEYUAsh/95RwCIN6A4yKpa2dPF32zC+TSU8ypv+Wey
j/9oNVWRFM1EhYKvv+ClhiFHQaNFmVxTJQx1eVDmi8Pgdxa+bp2r9bf+WJzKlEYc
BUASQIgWj8+gN0P6kWqfW1nU51jR8f5EcKWh1/4xolZ7o/BIBXzYDaq5P1pTq/jR
Sm1JOcD+x7TC5EXhai5x0u4EmglOTwvT4ebDtPo0ABpaKDeldtuMs4q8C9VBAqy4
JCjwFzcNUYqCEXSyiVmYyrUMORv2dcD+7v74wcsN1t2jo9q5A/Mfea6dbP01b0Vk
mgHY0kT7AJ4EWOafJIl/xJUigAOad8JMYNCVR3xg2380sF6uQG1+VSUM5RugIM8g
dqeocEQmnZz8Jh+fohvgjIKYW1rlTBfu8VhnCy5XKBy6gas8VQtP2ct2++2+yUwS
Oe6KRi6g5Od5D/i5d4e9V8Stj1aYfDyZtoXNb7MjtaFGx48YaAKI4BHTmG3vM5Li
WmhoCGko4erpmKQDJfrJmD1XVuFY/5e7S6QyMR4fW3K95MXAZ2/CtRBelv/6Qyqq
OfWjCFO+uPNHEsZouFxlEjB/n9Lgf8TGFelG0gafk40HNt7Wq1jOVJGNwciZOOXo
1wBrn1JguG9bI7rZ+i/ilZOVcLqzYFO4w5gxicwyvXv5OkYSHyweqpvc9GzWjjqP
VKUFDSBv9SuANWpFFVIFyxX8Xhbq4nQWO/YNMmYlPxN2L8oDcOdZmPd0W0uT0hfE
zK/nzw4rsnuNVFcz/gZcFJldwibVEFP2fsXGB1gW+6baxhPMDOlbTV1B0uKIDHee
PHxCcKRRhDUCCNcMf7Uc69hTS61VXftQHBkkejM+iOIC6RpISYO2i0A7Q9DblU6C
uxxYxVTTQD8uHVPIiqzpazEPOfljtNolKJvf7lutqbxOiFWVp586PAU5LsQITkbe
m8UeNQGNPCeZostg7hTqYLDuhjACYiDQd2NhF9BpI//FqevK4J8daek9kxKGDDqo
yWwx2tT4gv9vOLg12aRr01LAFydWVINwNsFFF+vpEEoOGHz9ClipFqWV76Km8rYT
orugKauBiwdih2XAwTtYg2TneWkPPcnvJ3TNowSPAmgA8cONzGWW4FMWgBtFxaBS
PhJLsgvq89RXwR8Yby0ZqYP8VhS37lAlInKCSaVo65jifIPYfOLcGJUI5mJtoqde
xxSI0gIOr0rC8FHjkfUBNRfyc/hNH7YYMjCdvPyhy06EhNTg7mS4c8Np//bVm8iB
dJygoSIBlK1KjhkebxwjeXm/KuBNRPLVDUsW3B+/bss/7ZdxOPoBhZJS1mTU22yU
2KyyotHgT3bkrjKpQC4mO9wwy6KAA8EkZnSEO9rb1trlnKP1x2Dcv14bxWyrrdRX
my23BjsrPgN2CBOrOx7BEqilbxKDy02Vv1Hs4jWWlmHrb0AMrDdGXZ7mr65eyQRM
8VpSJPIB2EZxnrqV8MlpyuQumA6ZtlvN2mCzrmoNSmnQp8wn8/C0Ct2r8dOf992Y
DSKO7v0tjyAa9n3strREoU4EH32jJ6vv8oLnIaJrzX1xQ+n71m9n/G6AWgdxuEjU
JKLRXWVTovE1kimmicL0Lmjn0Ssc00Dj50QIByfiy4cywckzFdRldIjbDCaDzTBo
XAUGDp9NU4sl4kxk8LO51WE6OXDvVjlTX0QHjpzS0rdxaoN6n5Ytq+EAWMVtCjJM
g7/VGqPiVF9ZPzLV+zOJ36HHvBLkezvqeJ0bm0rYaRzNsCIlA53wgbMEJgwb4huH
39QEKT2bsxJ4za+smXXVIqGWZh+xBOBe68N1OUxuyzhqpA0OPs+zojq86fAvGWK5
EWnhP7Zz3VZIaMg/53LN0plLnSjc0yYTm4KccuRPeLtWK8LL4LU16pFWdNrqqIoV
7q02Z8AM4ugVgIVKahKZL0UGkMUAW+tTGoz8npavTi/oIs9FmL5slVVE77aVN2uN
jqmyapB2mgP4lhlcPXVq+rGWFDMGg42kQiP4Ek2kRNqm+ShQyZfFm8Ld9oy7xabw
SiOYcbeTyATVkQ/+rdPPn2ROS6DvzvRW0o59L3BEdJb05gb4TIqqRDpPPD07NQiR
pkf4efK20c6ooVC7bGEFZs2SnRZDxIVdop98z3PgkrQMMr+B61jps5cKFYl7ttE8
ROb+Q80ED55YPeTRGK27Z716mZD8yZi5ZPM+t8VQ2v6dSrN0jXRPzg4bYOpswSQH
aZh7uiKkV5qyQ/ek9WrgGPOUpE58dZkZlV5DaPPzzPRUjHi4nbpfNRsyRt2eTdh6
HGfVfHdR+O1dbEBEYWs2v+oYahA2DWEYTAd5GiiGBKVVYi5EPMBA07xwZ0z1dZte
V2rssCcnz0VQVeNyHkm9PzaPXgCF4uaNAARwqKjxt7NE3WmUFZvr7GAdvOywVMhe
N3c4G2qyVKX4A6y5meDGRL+NR0YnhFyzuMqAcNsOQDmGblj6C7Dts+db17N5RnJ3
Eisg9nK1TO/b6MCOI5GMx/4UjWOQwgKupnvBXTGYDIW3OLFjlqAuauBKP9bUoRB1
n8D02h66atCpoE+ckBR44TE3pKj8HGBdroE6jG9Ly6Q6v+OzXMInMw2x+XWv0q6R
l+2/L/BhsvAElPNaJJPgkf//xfJ9TE/1kcOoC+fpPlj9K/SwhnBgJjTr5s7HPO/W
aT0xGsPnRbkMdC10pQE5LGtnGpkGee+8dWcpKPxBD9Vayz6jSCoaAii7RU71wj1u
++0mWNh9TQlUReu/cbePk37IiOsr93/BqdcRWvo52vJ9nAMH8K3CCczduBl14c+C
4xhShqdnb1kxSF0jOnlqs6cn9foz9CLVv4E+xge4sNEkbPXtyCVslSS/JYhWZID8
+8/Tzo3iLZQtiIRWgfIpYd30G3Y92TEaq5GyLq4oylKdFw7LcGp3UIYiGwKOph62
1+vTyh9VMCllgSqVvvmuUg+YgpqPen5RGGYE+d8SJPh49+2GFZ783kgr8QJphxzb
QZ+KLQBDaTtY14LlIq8TBVx11JaobPc4L9N/UJxSbSPOyXMyOpi5o5owL2DY8TXq
96XB7uf7zRTDSw8dQS2KcI2fr8sX83mbXIXdCxoUXelizNAFxGGYyew59raYN/JU
GIagdKjbO2k5pCtu+2wXTf2IuHpwEimiS3xv8c6MaNBGlGAQOQFxGo4gbR9jB96/
IdaR5n8zafUA2OCUu/b0cNtLcdX4dDwdS/a+K2RKmhA1VJAXqnVdCAGr3Vcf4nEp
+cRC+zrmULHR8En0LLDLeCoVCx0GWn/r4ZJMDLf5SIZf07yfo8joUPxRYpNmb5CI
fttBCnJJsf30gPUQdACrCes2wQYLVRCo1oZz++WKMH4YWPwcgRpBqZ6tbiwdKNrK
5f3oQ23/LtyCE/n3Z2b+7Yc2dKKHRSxy3m2XR78X6wpzWNnkHs2P2o9SvjvTXcvv
HFKOnXqPIRKmZmO0sneWOxWpqOxFf04DICjFQY7gnuf+ZNAvkhXMzfCY2eubeNhG
gIiY/jajDQHqDCw6nXJ4PglVxBOrunBGS5hQkGjIn+uH3aHEyATwb+g6gOm/M8f9
xo/cLvT3uIoocMpBx+M6UYQlicVxTMPRC3MBQOCtBNUvzTG0Ds3/tHR0jbPsJMN/
K2pdiXH57GKvEGh6j92e/sNDeyIS+qi5LJUwajAjvBjetzSlfxwVO1BQ5pfNU7UA
DYHjaIG15S/S0aEi/+YuE2llsCcwaVB9HI/Luxy+Ghw3y77xgrCRezkhZevMxFm1
e2igqLgYQyEZNNOMesGWl8klGjSmbuNl33DBaQ68BLv4CzPp+P3Puiy1jGJ4BCoc
WhZ5GNy3lUTwhNAXHXv0mcCmfsG/kV5hMwtkaapeN//aaAe8ZCqN9lcgG6NZ+dL+
7SFJadOVqjcje2m+nLtl8f63rdzBa6hl7/ZFJXM3MG573LemfQ7GuuyjUmUmyJXx
0v3GdepcI9AEJLqJ4ZDhixX0qIhSeP2M2XUmEdqg5klwD5oNrJGuaeoigGNbT+f/
Fn3jbjV0w1srnddZnmZr/JJcX1TZ9BjpCL7Uza1aF9+i/8UfY4Rp3xQ+7dG5V3gP
oPDdHqN2umthNfjVweoLxOjgzg7sDp0tCpYTKDP36p2uCUOPSsDQJqCYq1zY94km
siIR5yZBCS0HiQrJ4UxFb+VsJ6UyMAOBqxWfcP83oDfe0KGRvXTHajAR7GY99prM
Wne6lccuc7fexJpeIkxPejcKHnfosAeg5mjMAZZ3UlXm/yf/wPBcb0tUNZx2u25y
G5WTsR0UGUIAv6E9rTSduuPbOCNdT/A8XFvuy3yxJa7ECSrKtpdkIZZdFG27qpIR
V+kPJ2LHHHzESSVwA3yrLfjFKA3viCRS6rdDWR5Ha9F4jaKBWcQQ3VMomgbZ7eRZ
5pSzzvdDRGT22EYljFy9ERc+v3TbzYGPqfp+pS7QEsPf0Oi6gqGaMeqhAYRk79Sk
`protect END_PROTECTED
