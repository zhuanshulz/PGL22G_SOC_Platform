`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dAEt/XxfZ+fjhx4i3qzduBkamRxKA29pW3T6FlRNHTSBiXU/qhZocAYAJn3RlIv/
s94VTNlXGQt1ScpAugOM5Iecuc9OQYNdlB1Q1oubSh30CO1AADfFfHleeP2J8laI
Gm8EHVJ77d5W53CIXYJaB9qPE9kAjxUbSpb67PwBSfRw7ARdPE6T4V3Nk5tV2taU
kZefD7Cr/PqQLmGyRaFHsn2AI7YdlKUhtgg1pTIT55xuCOMH9jDgTacy9GcUpwHk
mB120Rq0eBCt6CfQXgrx+5J2B6EB/oHZCAaLZnu13oChCV6JtSouAt5NN2Rn5KQZ
WS+xi/lCRe7Ff2lme9b/hILPQGsUIxwWFg7Q3ds4elHTjOIv3JufQlF6JyX09Bij
hCncHavH7vkkFb7FYbmCDDBPZ1pghaYwRtd5vu5+gww=
`protect END_PROTECTED
