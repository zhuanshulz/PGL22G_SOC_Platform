`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yXdOkdf+r83H/oKjj4Nt4yZFAKftaCdqx8lH5HCiprekYIMeoXLQTE4RCKH0be/Q
SlBAz8V4w295GxJVGxwAAiRcTDaAiLDADkxWZi/U7eb4rb1qLRBYE6fWbpMwoPcI
uXbkhdfv1ae6RVcm9+mi8CxeOg20qe6MOSJlaqXs7maopefRSnJBbUf0XJn4uDHP
aN7kq4HZrtjCthZ1EMlWX8iWRbGBeOvJ8j3tSQwin1ClNLVxS0WwSH26kdyYfkwv
ytsEemRSgk5SMDi24b3m5i6NSLo13/pOw+oFs/kCb/ZsU9LRbSAnOVcqodJJdAFm
zwdetuuxZTELDrICFEImVk+lRyTV52jeHjqKwBrbMLAc7VgjnLsVx2THsSS9pIh/
p5eVp7nSTE6OL2Is+vwlIEd036TGR/pUkz1eEQwgBbKkGxNzYUh4uJmtlgRdSV40
SbEUBpjSI9WAgq5mOiGorsQbNpxxJ4I2jxg2d1IRzVO30p5686EXgp2YDkXEMIor
rMrNr25hNnC42M7xwqVlZI4LZYHjO/I7/3RawZkTcScH8ERC4vIuXH07BFLV18kN
SiK8kuCwToKgi5+MtYvTBhkmpKrYzlK+IH2F4TRYiNKTnzUWi42t60NfTM28kncK
JsXl4V2QLT5uWd4aoJaf5W9RjRZK2/Kr5EWhBGDVUhspz39tWw/ntbZfll2ayKyl
oyn01vf8ORgg6kqOB5C9kzkajKnhWblrI5nGKTTtsOfNnpwA9IlUHd2XXJ77CHcy
YcQ6IIb6NYgVQlryCu6RVEfxgdxzb5etuvZI2DEWFNGqV2JIRcECzLAzvDjjUD+M
MWoALi1zdxMVatql/ESpeR1e0T9etHiFMo1DaN+3e47Y9wCTKzJMU9uNmKWMDuWx
ZjNuBn4ZcUZwhXZePbJxsgxrQO9icYn+RafobCT65mvWTwIOAQI2G6wuUMONfjfc
fq2lSMx5J3OkQbLG4qTsWY0fOT2AzznXfC+HObsCw2VTDRTSZqxt00UbSY0N/+HD
9R+aHWfSpfNZ0Y+Sfaxzbv7s7RbiHhx68AMBOJqVcz1H++5jFJYFJzDG97hiDrxD
kC5GU0QaVb1sEctYD0cOy2WU6/uEgyikIG0XSxGPSZimstHfDRWhwQLgc00cpxID
n4A1jIp3X6Em/lTdR91yOlw31eYVpwfAWAOhNGfCK0bQBjVy7h00QR+85krcOymn
nz0CS1vShscjy6Sp98fQf/NeiEBeya2a5lYjkbGdHCtu4SZzboslLWLgU0+mCTVr
lZSJ4gAjsGXFBIZj1+6AJyLHxgsGxnYvmtg1iyn6gSyyNx6aoYGVgqbIIatDqaSc
R5IwuZpj90VEFHKCMaLjJMWXuwxPfkcJuc0TCRuv3keXHvugMstIuqwL5zzjcluX
DBr373TH3md2DfQXIOcKf6eALr87zqJC/+7gdw4ZNQSZrs60TfLi2lCyiz1QnRnE
aLIBpKJ5N69YFFg3oXzT9Ph2QSp7VPJru5ql2GZu0SzBLSuJYzhR4MtQkrro3ecv
u0UjdGLgbiCzdDTsERkRs+jWQp77zZh2CvFSU4c+sK8TNY7D6qiOnO62SmmFjFC6
9yZK0DbAFEXWepWr25883dDps2b4PrXvXSq8nXDn6qcIlCveg0zEXlvr1RsvKf10
sNuC6+2A+Tnt/zM8PZpR/sKHfafDMIHFNmR6dsLAssZy5QHnwh9hv+s8S9qrtRVb
VFovfYymkJTQZJNhdO4dn/BMJdFCmkv8dKX0z2cxFOG7RtwfO+KP9xxtYsH1YK7p
qebFfaBv3tc33ffZKvZljpaekURXWjfMEQUbrykYc7B9HAJeOGK1nfnYGGEisGpR
SvLBAGnnTOU4+leXrVguvg9d7QJ2QLsd7ZPyN2mBCn0Y+qdX18BeaDMnleVcip6K
byfKJuXVScYoSz3UEPJjYK2VfT3oFj0JM9JF2fmSTRqbUtjP3koukAR+gbW8c64w
y9ddKY+UVjK8yPlPqw69Mi9v/+G97X+vQ+orxLVrr3XWypQou2oera1hO2qYsV3s
YohzUFHe6ltxn61ya1MtCGX+3Pu3of4cAr6MAMkHVTLDDt5hpMnDz8J+WUfjNiUH
fDJHWKlEQRUgzEw2dUNd/Z8etsE9ZwMXoFjAJQeEBgG9FI/oAV3/kJ32TaxX8RO8
RDR7zbytpfFD0lMuctxh7JAo9LMGv791sgm0mbkiMbqvVp6nuqmqW6Rw1o25h0UM
gR17jwfxF5reh9P0QrnY/wV53JNOlEtLnkmXKpMVeqwqGzSE9wFh/mXhoN73MIRb
6p7nPmVWvX8SgA6cWrEmQiSKRCMv/hnT7t83usRg2/Upny02WQGlrm3UlgPO2YJ8
N9Jpt8fHhEvrLHL0YaVgVoJEXTH3JiC74mKHXuurKzAmE+RvX10qFLmidBO/MS2H
oY64XkC2KFJVPGP9QxVsDvV+jjygcY3alGN5vTzc8S98wrQuNPsSETRcsOuok+is
aHk5WqsuSVn/VbBR/mmGIfEHQeeRuyn2AOBCAdILJmmEKH3BvbTkJf9MG8SqIukf
p0TdQTzLy0emmYo4uov4eOnui1fRngXhu7ezp4KwQOoYZqV04JwMrtoWj8ZzTmdg
8mEXA4ZeaJNNeqJh6BYSM8PVaf/K4xrdDm9JXGRe43uvy5gWgg7POQcSDuTkg53J
FFPnnWKzjbWYx72v4qVDwhjfqaKsQp2fwcsgpi9vo5L7+IQyzbz8MfRuL7pqJ7WB
pLck/Bghq46USRPiR2v6KA3OM7ht5b7S9csbKmt0/geYoR7SSiVOTNBB1o8ff5fB
ym0+F7OerCPP64OoOMSkmU9Exmjs5gyNnc3ZYcUKqPE6EIFwsXLbnlE6RL8bdb/O
PYJ+L8NR8bEBJm6s95sLxAUblAGYYjnAMxtwpAx+0GBogXknaCRNTHk3rjzXE/4h
cg8QFtGOza+I8YQ3RMQqZqhSq0EimuShRVnQ+1Z5vp0wRfF7ERKQe/hF8zGOoiAo
JFzg/RKn43leUTHQUdEgrcaYQ+FIOIGpNVA3wsvDlsF3tbzujfjCWVuICeQjMX6W
v9yIJkKJESYuvF7nohG0+45kT2yAN54o9ojHSCJYKDDDNOESY+eYThVmUlACMD53
UlSCYJUHURZqhyzaDZIBH4RnYJxSGhCac2VCjVPVkO/jrZ5T50JBB03ew+WhbTJv
+8FA3+rYxjbpk9PngYcY7Ldpu3bWm7MrTGDcpYlP8qeD7aMs2bMm5HtknpVbqecG
QU5eL8ej5xAgjGNuIPWKIg==
`protect END_PROTECTED
