`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b5Fvvd1FynoS080UwsdBiNx2DMrTdWC8gJl3zGeXBKDSmFpJpNkGHDQgAAGTb1Rz
BIfog4xUw8f3SHpwR/pzW74jagd9SaH9OIN1AF/XzWJ2m6U0J1tblSSeOUleW7bc
QjSBIhb3swe1NlTU3MJgjT6X4Xav2Zwc00nSHbSmyyUihkjnDqviimHVgrYRg3Om
GZMDLMhPRKw24cqb0D22dtJSReTFDKI86wUgs4MrO+Zt8dBn+wsYBIw01jB/8lAr
1lVlcxFkEdXOn7gHrXFh1D9Q7Q429Dgl4akjCL4XSyLcfVNIUE0nhcCgkIe3dx1U
0Heq/SeEHv4kH8hBZKwQH/FpXISS0gfStWLFgQzs/M/z2V+gN1TOIhKrOV94QH+3
RLZdkQI2IPaNnW+ai0AN7jFTlUvI0/IoptzY31Yz/O2megR2RYLBLPzNKo+/vYiy
gAbrkPE6wIFOZyg5HSdF18/i2gtsE4mmgxxAQCTgfY8=
`protect END_PROTECTED
