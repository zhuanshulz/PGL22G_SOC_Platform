`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KxevWG/hHJtSayuU6MaaGo7IgZEBm4j/epYLg5q6L6NcWjV3zDt1x2eLiJf1y7vQ
MX/ih/ipzPngQ6sN0H0Tu9R/VgkGk1FdlDBTUpWyeW7kX8blJB2RiVaLpdT3JIVC
Jd+vqDWlD10KKa6HkoIOkYNlJamyyVK90tjOz43Hll+zce+wiTYv4xftrIv1Uxa3
NIIeza6g/O9VD+LuJyiFZtzZvATm7haAYnkvxSJbrBVOiBzUwcvMT0gLdfCdg9wK
kJFlcNOEEnewSoxcAhQ620+CxDJTS9qOUn0i6VS0yg2+L9G1BbPJkwLaa6huMTe2
IgcSLZVCHtenrAVy7B9SiFrGn/jXy8k4xfCVUyIoRZd5AuNb6NRAzRmQ5R2J4mk8
fXMRBvmQH7ou4d/WTPUZNRfMTWW3sMgSCkjGZiFrjh6r1ockaI+8RKz6ZLIeGIFo
CPjAX/cD+/VUk1nAGRfwPNIiWsRJsHAckKAbL6UFt8oy5ksXDBQBxItKSspB0I/6
U+1o1qlyWzGHr9NPVRLg0ABlAGkNLSFwSdtcYqzR4dCBsC+wxvlVvsERDy8XoG1M
bfkp9nA+SVZc+9pBcNXQof9szC0164Q02d5t544bq82ig9lzGOYJiERMMdTyD9sx
TeUmZynwuWy4GY3sPtwSHZt+Ms4c4hkjZ4RDsH14LFE=
`protect END_PROTECTED
