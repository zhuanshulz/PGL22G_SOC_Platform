`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
94dwHr/HU7iL0AjcSV8BdVML4J19uJTbHz02GXAWIBuVdwQSu8lDhb/cezEC7BrH
RgXDxGij0ns5T9SF/vAVeO+y2HbuMNOvu7k3lG7dikdNbzZwpBkwFyauPbP6IZ7f
HTgrC8MadxjHPtPtSj/pO+iPCTKr7p/K2/DgWrEeLxCM63o3x7nRzzxYw9b8UNSe
eZKn5C1emVWKx2Tkvd9o3UwUeZOAp/R2fqm2Vvm5qMbEdm4bmOk1+6NCgTwxCudH
YTSOIpMqEqAZiIC5N8hrHfgOKwdRQfkBBlniV9Canaz9fCW/x2hkMieXjeYUL+Rc
vdEnHfp2TiQ6ta3/F+/St43hoOYmRWMqhw0hqvfmWlqr3KUzhLzwHvbQaYftnaAa
ScggZ1BWQUdPmFC3IE93dLfO76e22EZI14YXmJT8PcTGSRw7nxHj2gF3UASR1p4+
u8GxEvEGE7n/UVmaaakTHaeU9SwLKYuCIXoEsYKB3c3K0ESZm6TnGsAObs1gzIfQ
1lJByx3fx27POl1IV4w2Zg==
`protect END_PROTECTED
