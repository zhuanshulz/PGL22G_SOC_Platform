`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mz0/JFfMRZSu5sSGct5/s/zW2uP5haBM7rANqmRDBT4M0zhoNHjUvpbghgPAZIeP
/r2sITqaeHAYDiI/eHuKRzKxOP532ZNg0F9G5IIdYuQgKHEp4dtntRcr/vlwiIAH
GpAOMSWjvbakqRf1E2u9lAdq/J5xIH1fgBFl+FpRUfNsOTdmXhkpwcjNi2tNMKJz
XbNXVmDjfuI0g2x3uWwszFYHhZ7sqCuRAMPO7U1G4TPQr+ODBjU5RzEvQ1cWU47i
aBUZ6N2+zVZFlw1qEoIwPJV05aT46z5JccDL1xvSVk0NADGwhPwgUQMF0tateGSg
hyHk3t6E9XXjVWvMN6eoTk7Tf7FpVSI1mgJ1lgnQa1Rne9yeZAHuRyCFnQGOu3Ir
ccFapkv17+ozSMIs+FkGupX4+Wuq0IzWcXwxu/ecvkUh8PUT05F4uEaifh/6+IEr
eJYXkNJOJupfLOj9PXsMIN+CThagz9IYI0zt0SybBa7DzQy+2Kp+iIul8WCbUfSs
lS6yieSrvEz3I4tNC/IG1juRNJvUsfXSK/B/njHDu9+2AzlmQGMWD1xMcGW8pjN7
g0YkyS1naeaKgMTK/jumgv38bCACRFJ+BBfdZOtO7c2IACTYBia8t7OyIVzv6vfn
CDQ+eSqYWKF52ltoon2QAqRkqdCzWc0yP43Wqpe9F3V2iwzGCiyRBTsw7b75f1dF
FDg50jfb6VpIIPqwme7JTSQw+cGXgUDw7mHVN3C4cl3hnku6BWRxUqv9QRNH6cAD
1FolnXFAtIWuIui7Uw9xMdhTXdPqtvXJePpOMBzIiqH67Lnm/WR7I9rSW5NYONvn
nZ3o/vfqv2gwUX8qHQK5UFiAO67pFlfZWAPR4jFny1IfqOI9r89kumdXP3NbPl/H
3mJ34KsJoWz4zEqEV0LLY5Lrgi5KOpY3iF4eM1Wut6wuuyyOASk7Br+sMNHGUkhF
wc0LvNL7DQ+mZ63ti20QvRQeqP3rhUGH+WT281k045tjtxS0ETzGys2H3kDTUzXK
0mTD0LLCT8jtKu6pHZKgUhLiwORBirU/bgQjZwGXAadDcUz296dJeTbEx8TrBi/X
Z0TWw4y3uo8n3PtH+mQkeN2PMtuBkVWp1TSuzt3GoeTa4ga4bS558SNkIY9sFd3z
pxc2PLJWGak2u4xYebUSb1GUcO32ZhLAscm7ABSOYoSPks9T1T3dN0Pe44JdrYTg
9R5DA8SvJBxfCqSHTU24IVGnDsJuXNqTnRgsneAesyzEpJzCjAX86g7ROrzHe8jP
8u0L75/kARCdmuOrA3JXtCvKYJKKmqEFUyBXcH3zSFhLj6yUdp6C/YofrCOY4x1z
ljW6NOqOmlijXQ8nLLJKhF9TuRi9Z3V9YDvsLI1Q9vtjOCvtUCsKRCQMWe/8Re70
lQ53m4pNfux1MzkNtxHklpfRYKDXEGlrT8lTzHXLAVJsbFNLHOSM5QqoTFoN47PH
B/9zeHA8SBjfP04u3owvKPpopJKRn87edmQt9BTW4OtchdKeGVo2qQm3xA4qtPBN
FoYhM1M5YyDintiniddo7heQLiC1ZyHbf7OlJEGVa6VYUcH8NkA+g8uQG2aO+a66
kosvoQHwKyAuDviHJkc/XWTOj3t2qKHqZDCnqyFJkKcEhHVZyzA5fwYmaPZlmEJQ
sWRQ9t4JLy2bf+6wWo661GfmpXqr/T6kqPQEajNoopbTWSk0t11FRjqQrIv5zbod
waIGk/UOKbwYk2wVmJNxYPDM+OkIVUXHXSmg7JvJFO9L6kSnvpr6/BazKx5P3VBH
wapH3dORR2fHf5PL/wXE5KPRyN7S2Xcg4sDqef0p4WXf0amRvt+qKzgcm9L/oTB/
phpSrCqbW1CNLOfk7nwfEQytIAM494g9Q0Nka83JaytOkuqC18LeOLnaJvv3YRxz
69FT1ieMz1/82ZHMesVgKFSwc2tmFJ63ERqYMB06VDU=
`protect END_PROTECTED
