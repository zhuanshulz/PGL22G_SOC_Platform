`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MdPwViooBQmGjbmFmOD1ciW7HyWTj8B2KR808X15hsE6sQv/ObttWjNzGgl2VBLd
gs7ml0j4VGk2PznUK6phrgLgHLIitOGUGh6IiGZPyA7zYVt+5/wzi7hhRgYl8NKm
Xca7aMPIKCzlf6oKw176lmUuq4eSj88iHobcZfCWzqWErG7kPRWIGBNV/H7EciK2
p4uB4ctli3ILuGGRKJRNCMVcnETpJQOjmujhkLtGvEvI8u9BHI64WC9el7Exd7/l
AxbdfRY4HxLXkNxbwFfgvzqI9vbqiU1ihWjK1WxTdaa6i+2GVYq7ZZEiy8MJpddQ
yO4TdAwUewSXyzmWN7pGFY7N3qBN9cu+p3mv4hqk8m7N/kGmULGvRFVcJeAOLjx1
ZhO3XuFCOPlglZ290N51OuMV5b49SQ0X1XmDNukECRCuuWN4WKRLuFdfUvXVT1FN
tkCQY7S8rs775V+K8cHgu33+KR9nX/NhmuRdsIcV3Y71j7eb88WFsslSYYHtJ5Ta
Tg3iCaYmuTHvocbySGucu7Uh9A+CIPJwKS4XA+zIIQqtrm3OISNpaWlJ7HsTC6vW
ev7jm3+ZhL4FXcUKSDKMiW8d7nDYUkwW37gM/Cd27wgsk//E6Z6e5bjy42uIhuwg
rGGHoQTEZa8sIGBB3CrJtx+Ge0EKPEj6PZUC9eHiujgt2Bptv5hXz2GhBU0q8RLK
J56VegX4JYwL3v8WsbbvUzmF42YzwT4BBrgXsR+b9ayShEVrcdRtgFianjPMOers
COCko3loBEMqJf+4p2jA3GSolep2RD5Y2ljOW6naP1FPg8XtSX2fNBMCMdEvy8Uo
LRBhRZK2gKXC7t+9IA66WpXVZq2hA0IFiGD7aj9M88dWVeFPv4/NVVFBRhQNvWxY
/+/sgq+DFi5nE3OanuP3qegAYaZRBGw0GKzZNF3ibm79KiQvS5FL0hFsbR3jh1BO
9zrO1vTZQPl3r+F9UlbTA/6gZJOMj0XbX3tmd7rzvQvZTTytLKnUcDfVQQzrFwJj
cBlgovVnJ1ym513+T7Nv/AnmN568ewsYFWawvraDNRU3PYdN74rZUe8AYp2mVV6N
OB1hlR8b8dXE9P+P3+/fiP/sdqDfSbGStsBKnSgPZVjfZMPI3yDONcwBoe9woLzd
bnWvF3M0DCWt7+rh7avfewtKaTU3CZpJD4GK1o15N+Gzdez2dY3yf4OqYuOl4s6Q
HF7dcP7s2DgnOodXGZ056gnTNDPijbGKnVS5Jbl9Q2POrk/DwfYuSqx4wKuZh59/
TzoIP+UMU1u08IjyTawquMm/wz5RvhlnvxpIMBmKQRDC2378FlAtyc9/b+thY1N2
0i0U0CvfgadRFM9pCyWlAklE5THByafHkK0BwiV/LckJV31RTd+xc8dAlkrxqui7
mjHV6Vp30aMvHgL7xhLXRfID8pMg+J3JN+ob1AX9ly/5TpUo55kXEPoUFvIoF1rm
K9Z/TsC6QdxqBC5xaIknxcehz//RpTnf+IDESRVHM1Sm90REVkjxogQSsbPpVeXH
fWqAAAqIWcLeZaMFqkVY5hJtzeHBDPQIKZj62M5gr15A3LqEmKWGo7+mVWc+1Cf6
ApU8HX4iP91axYkQOT/EToP/ZCORX4QC3SXJgQIZQYwGf4vZjnV7R1jyRX/J0/dL
puGGdWmnH/FJ09xxjTafAUKsCBIQFh0VywjRbOT9JMlp7FlXry3oeGXDbpfqvzK4
q2nqOWwmIVHV48EeoPWnu3T0t1+/A8p3yTebNdYL7fuW/fhg0IZfldBkC0XEv29d
u9/1cU/D763cQ7AB6OlV2bYs07BrGTlsUILqm5GOAIFY5pFnf3u60MqIoncT8yHg
t1oEzIRZevwscq4W0dl+sYvRapl0BJrMEejPjj8LA7XEwfZes/OKj/Uezj+QJpc/
7++7GxF7DF+8+U/iUeWPccHpj53lzwAO1QxCL+fUX5iOkhOou2xp5pyuMGnzRZtT
2JZ4CS1n0jXCd3qwksk36X2CRwBQL49piR9N6jZKLW3qmlcn49U8SCBf+a5sxece
3Rbgr68rZenxJ8lmhZJPtkTaK2PzoVOwtu92aKmEUY1wkKGe8lghczZ/vbEg8/F8
hV+k11FEtVT4X4UuSDuRS0QGYc1c0Ycs9KbOV32dXfw0/E/oJEIb7zTTx2QvKpcg
bKKBtD2QDhgkdrHoNqfjPwJIwuhzeOH0wKfRogjYV/JbV6A55CEd5YrJH6WYekLT
RpDVBem9mY7B4Y/5K/j69wkhFTEw8/NIZkDY/KlO83XzL+Fh5s3TMHGqD7QBeFdm
ktR+yM4F+fgJrhldACsqdxRHhLUhKdunZYd/ByiD9/hA3LcEuqo9aj/raXpNjqsY
e4K3XAIN1rAAB+bNYpzVtZg+XzfTgdBNF7GIalUsSz0oqOtbmm7AcxngIsJGh5dM
9CsdCpsZFIaUvPLtEoJ7Plqogm3zhQCyFJUYV2wvIJ3wW7RtHpQUbQ4hTOrRexOn
wkC8wyPesjrk3RSCV5GJKPdEH64UxW0rOL5PWmuv1PTtHWa0SVD3riNsiAhE1nUs
Khq0y5SJ4Pr3lobX9sxPveClAxj2o8zI7Ze1qbR3qFH4x/iWUgKg9x5XQe8GLhMk
Y4kFyDqso/dZZOBEAJe30bOsYhCzcCNFy8c/9BcHDOmxDexPyI7XxmdorIXP1V7m
THrHYuii44sMCIIq4m4l1jrbVvP0XRmKxsUrr6qWo7POqyS3OV0nAABZ4lJDLXwZ
rz59w5ZFKwtaRSNIAI1jRc3m3H13E8FKeSN6/XX/BGBYBj7bs3DWUEquWs0FdKyW
2wy2xX3XcxlZ6POF8WaKVJC6JwM7VpefA4K5czif6YqXNoJ/SVYYUJhIJvBaeARH
Dm4qDlG1PIPzAjQ5oLuHiPrdi3BUl2ZdPDrtzXIfsFWU+O4SE8+lTZwOVmdvNpUa
SkNJ9toaJCvr3Ja7kAygWnvv863CR2nE5IQ0M7ot8qDZBr8NIRcZ4dCu24+CJd2G
64f8ZMkF+wdTqC/b7x1xEdVhxzRkhkO0ckXc7FGSSHjT3d9Mhfyf3GMGp8J6ls8N
ggD+Ujwya1e5Uzse3P7fIkVnrLQuSxfCSlrTCqcMZ4+X8+iboTnUtoiDgUir1SG1
btzFAuihCcazwDRU4eM/kVkenLARxDM+lKlr5y0bSWWPt13bw8cOdAUvp7+l2Dvx
5Xq4jXYt/0/WDZlny/hQU1yVlHQ6PuPjsddAw2czmjAnJEMPqndW9hBdcuIZKXjr
BgzmcwmwIq/DoU3qth9PwgDIZTiltruGD5VYuuZfqYT+Tzda1aShsCPO+jC3oVA/
euQmhXW3y2MqXeX+wfzUaKn8wzfqaaeRDDpW551lpIEZLEQ9Qz2Bzi2NQPiJVou4
glv78veykcMzdrhn3ZnZt6puC/NVAv6o4pVvFbTS2iW356pQL+wGAUdWtXshGhFG
BcOlw5PF16OEnO/EOyZP0GvrZIM/bCiQTXWn6bwx3ibmhBZ4OmD1hHOA0ej0DNPH
r4HnCX6t8rHHfSnwWacqrmDlA0U2STR04pVrfy7I7Yx5+LsGsJl3oy8JJGVe/AOc
YjLXDsxGZHQ8G9Hqjt+9wGCJ2e4prxL3TNy+aGbTmRYs5dd9y0/yHj2zjxMjJX92
y0ldt7Ftuk2PtTm+6ziT4EoDeWtyG/7hnDqP6vlXJWNpUB9pZ94HDWcI/1I1zmjE
PZyFVRZvZEhW2Gh4D04Q/vgmgzcZmlY3AiHHuT10URBwj3KK3tPdCab+xyUM56AP
pNfQCL4rbIJIhvLgxYW99r5US9hgsP6vBVdhLG9P516/wYH2wwyYOozKlhNNaai9
TRaRcrRZaVR0lveUAyoEYZkncJqE+k9WhrtrTf1lbAYVc3H0enxVBYQ4RX4zBe1S
4JINVRvw/HxXGnQE/ewxBULdlackcscZjnBK32r7CnLTSWn96HuWYCZz5lhZOVte
0HduGzj9LtP8t6qw1CsCXyjFLeBm/b/1DWEuSkUBANmwH+5MAy4NrXkhmvfWD4Sq
6V8X97wn5+pHejTfWqPQ/8h10ztbMb8/5iCJLRH3TwZNLEjW/+jOlKvx2Tl8APiQ
eunpCLoyNwtYdFIc1TN4Zu4IdBJrqitc3LVzNU/ZrX8+fV+A4JsnROwF5ha2R4i3
/tmncXJJIu82GgINNTu6+yIUdZA5T4k4ZUod5mCkekk8BveI0AwvBnsQGSQrY9Jk
2auhxJpueBW8QBUhGC7fr2x1qpESYNz7ZxiReZEkzH3+FFByO3Umjtr44IUm5eDW
jyEuRE0zTn7FMo7SU0HjUwDBVAeLZYiYvRit+KGXNHMuGT+DqF4zt24JIN0D1cVw
EefHUmS7Sa3Fw6MVhz9xwmyPdNU+x40jhMyN8oEaw5P6kwBOs5kP7ACBSz41l2Oz
OPZRovdAzdzp2uE1IbLxUq6oQCcUWPG4mXozpUOC1zzUUdvgyPOVbOWhJP6lEq2z
IyIototOs27cErDtgWlD8IFuINDmpkhngj930r+20r6vSrxjSgDMzj7eOugWK+sk
vOGay00Fy30y0QMXDEPAlqr34BWEevF9CXEEgZtReGvcUAF37mU1snqxQQloJcWL
LZ+vVWAMblZ6NXoGKjrJOQqYFhQTHdoKscWpZvIU2OXB8RT2kcEAPIeJuhXAD0Cb
rWj1uChM6MVPiXsBhz3/mSsz7m9wVE82M9GcZZX01qN9vKTIUW1RLdrFbwYaa2U7
l/TdQU16B8Jaq223KWzP307HhMJDeuC/qJKq8ibcIE9UDRlXGL1KkAP5PXFE4iRy
6g+c2bBLnlwiagNBjabqozEs3ALqQ6UPIu2wy1/GMw9odEGm1jpnOYK8L9smG0bC
Q5dyD/ZqydqY9yOBFrYO3dvZ5kQBeW0hk3OshKj2lW0YBfkU8LOip4nDo3rs4GZY
kpPuRmYmB15jGABtQhZxYLw0cAsuE8FpnDExgTMvhX7ug5H4Mr2W5aha5/xldEFw
nLVgyVSLYGWnmI7OblbRlYJ1KHtU7LsMMvKK0IF6/wMNpg7AG0Xmm9V20XGPUR0m
QotThOo8mpfhGz78ITBU3Pk3PiMlXDVHzdbQ/7N0EkBp8zJOeOtQxnq0HrD4F0ke
0r8e+OHwaMR9Cl1oonT244WN8dIoGTWGKgrisztPSqBspF4O16tgdG4tRDqhOl2c
o21SYSEfXUGNwRwKWdL/TmA24F1lDHFRrR836Que5DWUlus45hnYD5KFwvKQwbAu
HMgfXC/c6eyjh1EYNnKA7vNLukjRACTAyGzl6vpOcw7DGlVmFC9hACWpHjKCMS0e
Srl/hBqvwcgTvLN2nyZ8qcQl2RsT5O0CGbZCP+YtFqB7liMYzcysqNzWN912KuYl
y92wxrMhKe0if7GwenyFNN9L54Gl0mlp4ttWg2mDowYYmpU0OO5wi8/QPTokpH6W
XYX9K1GcCnuDd7bDEuA6VG9eP8icSKgvmU7/MxywPfyjBDG1FXPFw6iplDlmq4Yy
U1MrRl8QEHOgCyOE8srDVBvqNEPUrzH3uPEaeIi2bgbw5Rt3Wt3LSIUDY7dtAT6w
fpKIY0DKkEKXWVuwYd8MBZ1DjvnreVZuF52h7CHQ2a5ppppO26av8xIiChlkHukC
7DgzMe/35gzPZX6dbA98YF/nHIeL1dmAAayfv6n7gINvDxEF88eXv4iKVPSpWBIt
/xMxLIGQ2eZhh67X7hyvGy0/uxeYrGo6Shxa/5l9niqWeQNh0YEhTsmSxA5KRT2t
yFjXhW8OiykNJ0gcoZQlq+e6OyFm8xKdNGQt4p7CBaoWVvhvxc+VdO5+kdh+Z7Oo
V/Z7g/TskDMXqCkOiPlaUgaa/YuoLIc8eCbZrBz/VZZJRkBhbVgb5WiXVP7QFoi3
y/OGc+iFOMNQOEIBIuMtvwRU932gwbohEr0llJqIwom4gLN1rDEHWy+/iva8d8yq
Qd7ZDQ58mrnXt2B8n4Y8i1AO7B4WWAnLegJuhMMD+VR/8h5DYiSsKVKaGdI3C4mb
NCFDbCatFsl3DmeDeeaRHQFGH5mvw2v+cN6a8ATdvYdI28G6YsOEMpVZ+9UcGmog
Qqk1yHgVq0NM8Ti+b/hy1A93otVX9Kr9VHk2Yy9Kt4wsgDsFRynyeTZX/5d74LkT
kerCGDisP3hjOVJOfEPk8hLctDMfR72O44v2lYnw3aD/Ts8KwN6g/p4gm4UWFsws
C8Oi7XiMZSsda7VZGvpDE8RaVQgrbay3xBaus6au26ENHWzVyn2+dlCap2Miq/BF
vOm3xWAO6NVbyroZjku62Hg6o82KwKDWKC2ZgGoqJFSviD9NvonoxvIdgyr4Fdgc
UdRQSK7Uwe1iHv6uNpTbeV17u90jNf9jIb5/WjBMGEgMvkiOw/151zA6hIErFCAu
tsFcBoVDNM3Qt/yEgL6h97ChTHxEMhT5+EGJjT3ZCGp9cyi7AyVX6TTe+Lgj5/GA
1R/iJEpO+juaw2pvHkjBCnsaQXZ0BSMf2QhQEOzOqqh30oGUwY877QZvL2/n3r3t
y48+yMggUAIy93mZaEFDLLIDcTX6RBjVXKQV2KB2tEZEDhXpvXcGFBWcgGQcxuiM
6CAt46YHaIyMIHNpvVnzAOWnnNYhY1ADAnWW2BZ8n8NJsdyZYXdZABie7S9Gn10V
vNJbuwSOCuT+7CKrlJnsseI02qA1rLjY+yBzmNLxol6LPZMKvGIJ//Om6ZvGO8ir
V3wS3pCX7TsJpx4DicktnnARIWOHHoxMPEhi4+cryJ6igJ1kjELzE1C/X3tA1m0F
wVTVqDAFyFdeqxr0fgdkbcSfWMOGsAGvXwuN7GXdoE9kff89pTltvBe3IpRcNH5J
9b25ftGYZzrZ7iEVt3+iE8HCvk/CKxi7Sy53XGE7SHUi+j/BdvK+0tLatLgxrxFU
hVUJ7UeeCl0Df0/BBHPEvFVdBkg6mQl+o1j9Jqwka3T0jS3BYI1rYO470Vn/THmJ
fBR8+jFPXG7WWAADZyccZeFffnuc/ODU1sUhaFZaVJ42/6KTRP9Ae30utlEammC8
MrZjv7jihZJnOSK/8TKLdFI/q2hBjMIwUsiBKoX/rLDbSu8gZ/xwlnRJZVxt2ANQ
6VRNyZ46gXp6N3Zm4e2a1CxwCWXyTM1+XRAeOCvLjC2+5J8CD8cEwoCz+ZlGAiP8
pzWmPuU64P67fiW9zuIVAcqXjvGumvMustbrSw/NXp+lwyTKwbL3niA0DsAHXXWo
7hebsVDN6qfqTpil1IMa11ckelwBiJxsMhECUm+HRS9sNcmjmP5iqH9ytGCs8Kxh
OMwRPUZ1FIV0JqHKkfVVPcg4/gvpJudJbs8aOGrrk3fMNd+48hErQP0Ndh6tX2c9
xwmt1hSYF9Pc0z2nVZdL8dkoalvJmSrc5VrI0wYghQZEZFNBjAozanv45hti6zE9
t3I9OiDF8z0eAkVYMllyjMWu1nmbg+zykov5M0XsQQB351Nars93Ck3u62SnK9Ux
oBrAPkxdfoHK7lJCb8J41GC6z7J8n7IEKtFCOv3mUDmUYNrADlBFfIx1EZUMzCzA
LzoeUPxYm80Z1rqi5D05bVcGFGSTaALTd9q3L6bqcvtvfKkNY+U02YlMGv9EdY7N
rqa6iC/U9Sl1mVXq6b+ijBwedAukFTsEqcUfKyD5Xs6mqEsHCV7ftQOvO6Vn5DaJ
9JrCOcVAryGlVwJis/eLFz2licEWyuHV/+a0VocCdU9oFUPr7ueqZKWKxA9AwQ3i
nI34Igo0s8sj4W8kTj6SKg==
`protect END_PROTECTED
