library verilog;
use verilog.vl_types.all;
entity sd_card_cmd is
    generic(
        S_IDLE          : integer := 0;
        S_WAIT          : integer := 1;
        S_INIT          : integer := 2;
        S_CMD_PRE       : integer := 3;
        S_CMD           : integer := 4;
        S_CMD_DATA      : integer := 5;
        S_READ_WAIT     : integer := 6;
        S_READ          : integer := 7;
        S_READ_ACK      : integer := 8;
        S_WRITE_TOKEN   : integer := 9;
        S_WRITE_DATA_0  : integer := 10;
        S_WRITE_DATA_1  : integer := 11;
        S_WRITE_CRC     : integer := 12;
        S_WRITE_SUC     : integer := 13;
        S_WRITE_BUSY    : integer := 14;
        S_WRITE_ACK     : integer := 15;
        S_ERR           : integer := 16;
        S_END           : integer := 17;
        S_WRITE_DATA_2  : integer := 18;
        S_WRITE_DATA_3  : integer := 19
    );
    port(
        sys_clk         : in     vl_logic;
        rst             : in     vl_logic;
        spi_clk_div     : in     vl_logic_vector(15 downto 0);
        cmd_req         : in     vl_logic;
        cmd_req_ack     : out    vl_logic;
        cmd_req_error   : out    vl_logic;
        cmd             : in     vl_logic_vector(47 downto 0);
        cmd_r1          : in     vl_logic_vector(7 downto 0);
        cmd_data_len    : in     vl_logic_vector(15 downto 0);
        block_read_req  : in     vl_logic;
        block_read_valid: out    vl_logic;
        block_read_data : out    vl_logic_vector(7 downto 0);
        block_read_req_ack: out    vl_logic;
        block_write_req : in     vl_logic;
        block_write_data: in     vl_logic_vector(31 downto 0);
        block_write_data_rd: out    vl_logic;
        block_write_req_ack: out    vl_logic;
        nCS_ctrl        : out    vl_logic;
        clk_div         : out    vl_logic_vector(15 downto 0);
        spi_wr_req      : out    vl_logic;
        spi_wr_ack      : in     vl_logic;
        spi_data_in     : out    vl_logic_vector(7 downto 0);
        spi_data_out    : in     vl_logic_vector(7 downto 0);
        byte_valid      : out    vl_logic;
        wr_data_cnt     : out    vl_logic_vector(9 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of S_IDLE : constant is 1;
    attribute mti_svvh_generic_type of S_WAIT : constant is 1;
    attribute mti_svvh_generic_type of S_INIT : constant is 1;
    attribute mti_svvh_generic_type of S_CMD_PRE : constant is 1;
    attribute mti_svvh_generic_type of S_CMD : constant is 1;
    attribute mti_svvh_generic_type of S_CMD_DATA : constant is 1;
    attribute mti_svvh_generic_type of S_READ_WAIT : constant is 1;
    attribute mti_svvh_generic_type of S_READ : constant is 1;
    attribute mti_svvh_generic_type of S_READ_ACK : constant is 1;
    attribute mti_svvh_generic_type of S_WRITE_TOKEN : constant is 1;
    attribute mti_svvh_generic_type of S_WRITE_DATA_0 : constant is 1;
    attribute mti_svvh_generic_type of S_WRITE_DATA_1 : constant is 1;
    attribute mti_svvh_generic_type of S_WRITE_CRC : constant is 1;
    attribute mti_svvh_generic_type of S_WRITE_SUC : constant is 1;
    attribute mti_svvh_generic_type of S_WRITE_BUSY : constant is 1;
    attribute mti_svvh_generic_type of S_WRITE_ACK : constant is 1;
    attribute mti_svvh_generic_type of S_ERR : constant is 1;
    attribute mti_svvh_generic_type of S_END : constant is 1;
    attribute mti_svvh_generic_type of S_WRITE_DATA_2 : constant is 1;
    attribute mti_svvh_generic_type of S_WRITE_DATA_3 : constant is 1;
end sd_card_cmd;
