`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vBEoczmjf+cv/Dho21aPAetV+xVPVEI9FETTdocN/WDYBM2+hSBSozC8khnl76Bl
jFKA8wRJfxDoAW8BmBF1o6Z5FZXT9oFDUY1SttjFxgGlOwKo9DRTg4P8GBD4snQ/
yjTTDHmEq6yx8J4CI+mG/GAkdO5fRMfE3+Fp3Z+4+nfDo8+FooLkAaq2OKuvmurj
3e85ykN0PzfNaHOE/l7TAchMEdWTkeU9QsoORfFf/W2JAswFmaTvsXQ8V+MQVcBi
yPMPHz4XrK1vR0t3vdopXodebsl4ao+4X3RB2lhy+FK8uH4MNjLPj0vLL6ovQiPY
AWv3fmzkoTwGPTci+Q5b7ZBy2emuwJQbkq5on2xhuoposmpY4L5y9f7ZHYOR6azL
ytZ8vTk7M5qK0Pr4r/Kj8/Iine3Wi2uEVU8BlT5gmLxjPGS//GZuME1hMiFV3LBg
+kpWLk8Yyl90/fRY8rTWdt42atvIEQBnweUEoGerV82C/yAIABPxwGfpwR7C2MbT
6hoJ3/9W4y6RmdsJzANZhv9GQ6hs5F12mvybNvJH/KT4aWPGNo5myUSSGzJhq4go
yKoMl9HEmaUCZwhEKRmwydg7riZhozAmKP2Tt97FVxxRhL5Vq64iG7BbIMRHaKnW
yks2sCP5Hnm+7nU759QTtI8SMGYi+TxPOLI1ZVe2oC+bpcwa1/NFxgtHdrZq/aN5
RSzVlPmTVhRf15oNMZ12Gpy25iqoRnMEDFGIEbh5YDA5GRJaGIofzH44hHYia120
BTgVcHAc8Bz0IHyVpSWjpAzQfWhO7cGGYsghh14xugG41klZNSxa2BTmYjMCI/0s
2qWPJnEUzMlu2ESmddeX+5iwm27yuJ+TvCbSkjYF+QQLBGwwid7zVlvWodgl2mV3
gX3yHj6n0xOx7n5gtnrjTISseEirnOmZjWaGYPTLAo+B2e54s3mLfeWvGDNUEa3D
mv3UNvEZpQB3NbQJEmkBEi/ussZota6urxwNob+mPwGIib9+vrwwn4ELocglU3/+
Cbe+MTaHj5st5mwpTm7Qy3ljVrqnZKJSGuO5KlB0cP3RN6KiyVWx/mJYWMaRs/Y/
hSYuMz23Ks3P5Y33qW0apGf1p5fEiPfLlPZY0z6ht0rhszYEjdSCL+qeI0xrLDYp
E5QIQjfM614ku22Oun/dbKVQTaYOZNrGH36lvdoasCjtq2lF6yNL0mDigEhytBxA
JX6AGewqxptbUV4vO1S8SNVKe/tEKOQjjTN+l9HWduMOGBEDBaZgJhhY5H9irxWz
ubQ5AWetx3dcrpzMDlgEG8Q9B1smDx6tI6axCdNd42G3EzkPHZCjxSquY5VCa1ie
TLZPHi5a1/YtJp9LTyEC76CX77+qt0+Vt4spXw91gyZSgi9xMa2Aiyw2QIoulKcv
6oAPL0BcUNzuO9hL8ljT4vLpbi4U6Nq+DHmfjfJqSeyuYLWVBBSqu+8RK1una3OA
1g5My9u/GEb39BnAe/eYo/aJDY5azNwb1+S8dCUxw+Yy7jmHsLZql7Is/9kd4Zp1
3zBXkEB11+G0Q68yJ2gVCz7GEN/g2/0moMTOOgefAEUKvJt/lVzma+IW84amuMZx
fPaRULyxYCfQTOw+KVItNUV9YiWn0G4TbC5o9rJ6q93dkLzfL3KmhOqJcch6ykUU
sROAgc5w2tOKcsPhERbe9PtUSPiBB+qg1svI+HKD3LjV2tnjvhN+hcVaM2zvN96u
BfgOaLS3Tbx6+nEwNbULwvLKTYT43JIHmKgqUfFeT8y+sSWqDZkrO4zDOcBhqOZz
HA1obaVe4epfwvOUP32N2b/SGuXhKx2L3F9rozvnprDH7E1RHTOeFsGtMo4Xrz10
MRB74NiyDZSlmsklhvbeJhVVs0V2f5W6OoEEA8NaRlkoQGLCM+fe/CfX8n+tbA+T
tEVduvTMnh/A9/FkA0RRKND12L1t8zp/pZ9pTcBaV2XX8QcrGz0BeGiuTQLwj0px
4HkM28nlXJcpO4bzC1Jl4sW1OPK8xAg95iMH2qZye0cMCBjM6amlGox6WDI9VByp
D7AUVbtYQ6AU9Y530ETMd0MBlK4dvdkP6EyBB8AFx+upF8Jznsc34nfa1MjjgK5F
CzV2IT2YOhto/YkXL5Xr6BBr7muF0l42nWGnSuPC0UNgnlJdrHRVmC1vQX3PjBdj
5xkah7AtEs96nKI1M5CQzYJMtlcmeUOtn+sypwf0AYDrm3MAIiYaAl2Iq2Cxc5ex
IVTMWqPllZBMOhnIEYO3S592RcgGzduYnU72m3SuJfn883D1FSE7tjDPbi2FZxUr
ZGxXwSKH9Nm3/PbfPD4jB8JgCys5k2nam3fqS1d/DJtvr3DEu3pdO35kgfqMUlXV
EYEN8j1mKVfXaDjfWkCjntW35k2MpfN6hflsOm5lrWUkKovE2hJUkJiyhSzFAgv1
Qd9Ej9XpluykcpCXYM6mG1k+RtvUhb0FUAEGvlbyZkZG99/drFQnaVMgXp0ut4x8
eiwsAwQ4t6tdFYxeFJLbkSHz5thqFnuzAMvaXgV+25xAJooOl/8ozuVha7jbz3Nl
qboSoecaZyjPtX20RjzCNuxWUU68hGJNzEQEc8KyGYfTLZCMNk8ueNtwRTSeEGC5
ngk2GHk3+tWhiOvl1HX/B1iDZLsSFIjJm7vG213mUkQxw3FQ60WzIjo2QGGm5e7R
BqIxeIGR3dfusD0/gkyjp6WLuary6K573uNs+oWmsgf2oaPQj0p8g8mhOVwcxcVV
QVGrcyGuzD2OR15oKPd+z9QHh69UgWqm0hw+jVm6aHkrESdjrreAZ2Z0ScJSOR6A
HmCyOEKrnBVYfztNhBADv/jvoGz8uBPKBxTNPKB/2vl1rivdFKiZA5G3t8fayG0U
Gs7Xe/d6tugERa4VqxuoGJdDYf5oRomHYnPbvvfUgQ8m5nl6B/y+pxIIgdubpWLq
m2HePAi7hkqFrlhSZ5hyuP9DoN8AKmk1ESp9mbUSxX/5ZUbfd0ykxPMdb1IPcM8S
bKh1hLZwON3FKVlgxt/rFWCdlqxAnwu1f/UApi0UiHUbnYahgTBrDh3AAVZrxwXX
imFbj2h6iaiflzKxgi0tKNs8FUvB70cMVx1PToGn3pOpO5JGM3DCj8OGHl/huHmj
4EK5OTnOSQm56z33Qf6EhDXX2dIZ7MoiWRbxJ6vslGjuXjN7gWaKJ0EY0a0qATwC
OgbTz00jz8/Yk+fVRDx9ck9uaWCP3/20YDGR2kvq5UEqz46JquqTDpmXypw6bxXo
2ysSe9UqSVbbh5J3aAN5wJ6KUmI7YRiszMOzckO1j4EzZwt9lI7M5OuWglUws8Ol
uSfu+gMrcauFRBR1J+/5By68NbUpk2HngIdJWT1AlLyqH0bwpnkSIRyLOtYsH8ic
ShS9//k3r2XYGyK7GLNq4X+AvxrXAjyR/ocT6kcY2Xw+MrlGscBdqTFze5vqtNmD
H35Ff5lJEDXIHnS9BTxUHLJAdSZ0RaoeOXCQGQKe4WXmJgVxqibtzg352XJ/oPIP
B+Ewz7QVCyZsjbphOhtzzGjBtYW1J3r/6PrqaZLGMwN1gSmfGIfrM3wd+IXe1toU
CgMHENTkLex+k6/LVPxJoTCVJjSGy0YcTS8saoE7BTzjdgWvUTTHWkkrE8yY4Z4v
cCVp9hugsQaJnddXLyIAF3mElOYwRgDg5qROLankahHmgmQCyl30GNoSZ62B6aqw
XtHhKI7UpX7eqpJWM9UbWrLlTn9dK84h80b+lKqoLpdCxWWyl+aJ1piStEhuiP+X
kCD8RRiZyyELrqpxcGvGHVufLCuAqBT8ui2zNqrpwBtrrt6+H0Iisn/xoKOZgoBd
9BEUZ/uPeOyYbIYRdvP3grUvS1BR4kj7pw7z7YX55lhJaWU3TheHdwC5xJSduvKt
FJCY9W7QVmSknzzPSejp4jUUG5dqn3pLIJlwCsP+Q4fFr07KxUka6bDFvYiodt//
0FPHq0A/pZEP3Ktinof5STqtSpQYJDjvprPOVfTimAvYY2eVAd5UfKBa0dneMDCS
p78cNZ6CQEbWvHQ4HIv2RpevzvUNqc0MQQYHc83VsyKxcPC9MYQB6MjR2/jyjxqG
lkzMBfBZoZPU83ClErv0ZDVRF1rZbyTMhQN0eObr6Bx9fFrF1bgCpZjqiKKw1wTZ
9gGsI0aQsLPlocMdXSac+7wZXtU5/Vio/zIH7nhCGHrtI7e/b4Q+5p/7MHhUNe7c
48+as2mMUsYlYVyNsY/Hzak6lgF6YlxApHubSZbk//GvdZH7Wxs2L4rvhIZbr5Ec
k25N5M9kL+afYZcGjKZlSaUbSgwptLUE7zIPPaDLrGlfEYBC40d0VI5bvmbWavQG
/OgcNmpFyGUt0ByETHJyU62dduLkj8s1vlqHMD7ODZ3cqPNqdjgoLu3GSfyG73Ui
mFDoW+7q42OKqkwq9AZxMDVotEacFTO1S6Gi0dsoGoJRHKTHAAJMf3y11ykW/RfW
lptTnkS39ltL3S8liJT9+vltu7Tp0N7ZZIRdrXTywNenQ6S5Zf3waUnuvI6afZd0
OVIDxhKgz0DaBhsF369Ir9BHMo3/NhB3zM+1fvGGbvATiSbXrNaxg3jRIEqkEIej
CZKANHskwoONMpJ5ifBi/oK80pCg1kCdqKS0GJzKr82xyJACOFNAaqnCYKlDpuEK
sG0kntuzS0y7Ea0uJpl4IySCiBZRnLsLq4aKXfaRpOquEpL/ByNkK6UwIeqCaBuO
oyLuhq9nko8zZE0kmm3iKWBEsUK3HBfDlMqVbJ7GOSmG2ePY00u3C2Ltbdzy3z+4
URX+7DmZgGuqOxwE6Ouk6ertcgUHxFE37s0/m06rjoo6wj3yidplae+gzX+aq2lj
BlLnRD+LoreQAK1Q2GPWtdF4ObeQA88sQqvvaK7crc+rCgBTeLhHW8Dy6lZAgCxC
JnGEI2QgpDZgxPWzgOzAX8xXu3HPcS7/zbWj1dimO/YmC80XRt7wBeU27y+hz8Wp
j/IRhyNSUB3y9uDGIM8nF7AdOHynbs713e9bNEykILETpxevNsOQR1LnKEC8jf0a
sseUYyEzeh3PorwU7Vx5KVpLmLR4beHSGxcP13eERRmeJVVgXGQUFjmsLCpsJFW7
HV6Ztfu2j72oqhdhVt79IhnOydrIvOgXQFJDqV4gXfvED7cF+34e71DZZg6mPIQ7
bKdI3VpHLODs++cFu7WvoGf4PTERRUDcs5wKL7nj48MxVwN7MG7fDhGKsb5sHXK5
fx0TM7kZKfR7rxpnvHluhMIT9HZHoJQO5asJ/L/EmHdrbll+dyE65y9hHQg7T4XQ
sqheexNDXYeRsoe3955jQCRwIm4WDvReNmQbviG5TUUuSFEfUQpA2CVKllynzmeO
5vg0hS1cgsaTbewDN64ag8d8GqjsnjRKpWcabTQMW/BHeNub8Suy/+EHn6m+eh0w
R6p+wT0xOko03iAZP6ZXUca2V+mfQe0A3wVHKRJpWSgvIivY0ZCzJHMpishEdoN+
xgbRRmp7uycDBaUsSx0obgyLicQ24GE0j3FI+xUFhJkFAIHrbeUB/xmlG4sEMiIu
iKjOQ88wKWjM/C7xy0vzi3BHctGfQoHt0QozLV33OpCLzLvCCVEN27T3zFYfUmeh
zuZXQsiweuz9T7O/s1PFUzAZPU9bM6DLxrOzBBkbLlqpm1eYtU47fLQRwaSRhuqE
JpQd0RdYAPW6cgHKq7qbmd6CISJsAwNuNRrtrRLPPRs45NRfRlGkqZ3oYhy419Pz
rzpoF1LMW7IVRwfzYIJ+bmPJMheXGQHcgpySgB4GNaVUVtRx+weTPDg94CODDMvr
FfSJFO3NxOSRhkFZ1Mfp+E24k6sq3h5RYTDutI3+CdPpcptYSDWVCq8/wgpcDd5t
fPdbBMoykKmZSU2h//XWR8soLGace/Sw4YXDhqfB1HLNUI/7m9fl60SxjPp1NXGO
Na639kHEOxs3ZBLwLUqymLuE6U5OuqNI+sWhFEne/GDbHuykiwCtMTK81ZydoMJ1
K3AprcXNpqey2ZjZkLM2rmjQRdmaI/3ng1Gh2L8B6PgPkdkK/MR/E474sGZkwvuV
Iby5xwjo6bDI5hdCgMacCT6bUNDJqaGp5p18sAUzvsg7bYr1WIltI74hOJSnJ1kM
jF3wrItfRjnArJLrIz93jYXofLuQzXOmG0hUOnUmWX+LzIjQN0rhTCvx1w3oCh7Z
3OHe9Vh2wvG7CJnxNq6miVHeLryhvP/qwCNy2V/3DHZEWIkyBTIKAO6weB7WVxIg
S3jr3+CmMVDuVygTEJmq/vPRI6YHMACccj45/C8N0/RZF5P9zCH9TP6Gvvr9y1Ew
f5cXdBnbWGVwBN2sOBYpqSl7NFgWBQyucYYgPmWqciLRg4GU4tSurduHBVE3+/a+
IsZLmem1QnOZ4J4Wbw+xMBxhRds0bjJ1XObyP2Ek6g+Y0HKpl2+lhR5B0xVkeK0j
mgX8VMV0C+QHzI7/s3kBz1+hM7Y133Pakxq4Q9jlmjvAqmjaQDCc2a3/tm9P4pOt
BcR1QDDgEnhrYyg4Pm+f/bi03QLigWggXj2vjjQZsDpvf+vd/kbSR7YTSwHng88t
G/G4Jk7ZANv9b6eBhfgsNXqQkXDRBHjA6X4FT+pgu/LKVqUDpEpZGkPD3hXC9SjN
xwRmcUsGxiI65CModUhJsaVOerBogi7rbgQGSOKqXU/Y18qllC6u2cmhgD6LcioX
XlfrEAL7/yTbZTCQORnGyfQvDzsJn2/LWj9TlsD834o2o1Nqh2cs4jBw7SUeNegl
hEQ60jtjqO8k87lyKJ6t8fA+FWp84Tz7ZlwyRmMxfhVmIi93CmEYnrtBN2PMVsq8
yH6Vb41+nk+OoXoYXdQ+UDYxki15UY5jnQjc8buA97l1GMRDRYQPCjRgO9OpMMN6
Sofm3EkHdBQgNlzV7nHA3TnAF0Ctme3jtfMCs9i/zxULDkqNZfoUp3di2iOcmUUH
cliv060xBBP/TWNp8ux7vzSgx8IuxIkXfSaolLEF/sTV1i4Ge8FjBgcpZae9hElJ
WZphB8F2uM0ykDkIybkfUZ65sjqCGjs01IpDCVIHXOYEb0j9VuFig4wDt8IEk0ID
Sogo1OR1w2GYTVSNXT5NgIaIO1KmLqtFm4gL7jL6/U6ejlyNPsHmw+aMjvy5sKPZ
c+OgMHWnwO5MuvEUmUzDQIVqGQ4tgetGzjI2Fzye+tZ7GymLWZPNV14OiQtqLxah
zOzxJ2l+EvBjAveTaXqs/7L3m64ht3aoLdmDA6SP0QOO+NHEvhzi6fadD72Bc6NC
/vD5gt+FLotWPoVIC2vXetxgQVVp7eg3SpRH6TfMZQr7cIsdpmPfPk/2ovTpiJGd
vwkZ10Lv0uAG79fQA6IEw8w+A6sTPBZgtz0fQ+wNQFx/th9jky+0mGQe5DSFIa92
oAjEl4U8BW4lykc0pxrZ31tuzrfcbijnd9zCGoFI9w9hCRhkbN1rzbHOtPkLQ5ln
CO21ho1RiTRiocEunP+jJvZy6B5JGWLx/6VqiTqu2U26L+V9iCt/30js4e/3MeR2
9aiQvxP/RQgPjdJKkHkOIkYw758VsKlVPAOys1BeZkL2gNrRqNA82xtCAjaurO1u
FJ6+3fIIy1spw9gqpQWGkl2oWzYTRaN7hqs3vYgRzBbtXtAA7hbhTlMmZ0q5q+Ar
jFbal0cprM3+hU49dQR5ecknTUOXI37KAcNn9KhCUpUV3Hj8/cJtFxer/TAz6rGi
eZEsCbzXdhIWyjYoZazJfbfDdozCfwN8Ru4MyHQveY31aUIk5Bu5feoe8xz3KYGF
G+ELMFNu3XdJT9eC0qhgjJOznt64mD0YgHBSskvekaNletCmnUgyKSaDD1QxyWN/
achsgwcELBePmFIK2Nv5FSkZk7DK5TgVlsBpb2r4YTBOr3yEL4h0JZD397bbWUpP
6LMHWHQAo4sasGy5+LPXKso2zdyMh79T2nRJGmPcGapERFXwdNJ2tdkTcHCPOW4A
MERTKogxBg7cSFx7W8h+Otz+i5BGnTGBTFNt8t51vBZI+xKR55LBi6LY3JU/anQm
E5Cy5+g996ixckEkkU3e55nvMQ/gcxrijTGIxlYMfJV5ect1lPMqqOiSclDYdOeK
WdHZPrwCVgyR5cFsLiMqTE/ZGbkf6phbHYcgyJbhaJZMyXjs2P3kFkN4XYv+HNe1
TbEtlYPWba2M/z7RAyLjxRuHCB+38D3hW0uvvfdhaD74xLmgaZOXWBOFLdRad9Tu
XCR2GdjBy+aVewo8w6A7qA==
`protect END_PROTECTED
