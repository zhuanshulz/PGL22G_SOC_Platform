`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ALJG2/mo/HKJZfpPk9IGzzqY/6Y7d9V9T68bJbp/YQ561qRgELznoQsd/px0N6z/
5MtxrVcgLz7tknodPl3j2UV9J2F0BBVg2PBRhm3d6EcJ1c8zW06BKGLnS2xJFQWX
1qtyDYRouBMUWR8bb7ws/m4qvQY9EpLvbYHOlLpqzaCA69XoYo610JcVRXDtY68A
LuXhWOijNuqehe5M5X1bOFLR2G6C6jJufSuJlcue8Dmlgmr+wvT5hD5IjPkWkaCG
XSr58PQ4i4iVJMfsawlxFlRK0spT5w8G8WYw9lRK9unmmnC0sRY6+u/y3w8nWfFZ
Sinh5/+zALkPbELjYCPxSYa1Q5nTcsrGQjgNgsybz20ARKB3sR/2bdmDWSwpa0uH
4xl12P0LwVlAnFzj6Lky6YSQwlw/ORkXycNc4o7QDY7imQYNxMzA+fQiWtkSfi+F
G1VnGTiP84+ewqEHuLyFPShm2FzU+tDvQExsu6osEiV+5iULMlx77t3VAGv7HzLP
Tvj9/wmPbJAm5yYGvn+SSUCwoYvyae04s3cl8fZUDPSvtIEwNud6pjrIwMduwcQl
uE/2IBTSYytUghzg5Fcl7JSUg3pwgowkRMAw7XVy6b6IhK9xd7DYSB2D7BkL18O1
Q2Dcr4IAKQ4BXt9vqbPSpVmbj2VTIbkjLACzivxNOvDlQFb7IrnVs9Zxu+Dpe0j7
GfRCpy9tq7UJl+GW8wdu6zFV3/O53guU9JcOMDoJ91CfyHJygF0SNegPsX63qEbd
XXMI78hZJt51f8/DCBm9k9VLv37U3rWE7DpJPZ1Fj4M2Lk9Vf/gPXX50/iQwSx8x
4wHG9rAWhJlFiTCamNEQc0vdg0lAGzFvWibUDfoKpulhQIWxfBa4NRF6nSviz0eF
aCjhKwAWLcRZyl8VTxC2cQ==
`protect END_PROTECTED
