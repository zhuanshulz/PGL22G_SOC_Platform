`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tsvUu7HdljcdBqGECJQd0hoR8aG0DuCy6I2pb0GjVinxYe1Mapa4Q0IEpdlS5V0J
vm1LdMK0SaoHvR7nKa/iCMQ5e42NKOS38i/d/Yf+ODpppnaQJAYAN02Z09kcPJen
1CCJ5z98nzmeUuxZn89EgI3TLKoMjCbQTLrWheQ/NZfeG9oNJjW2UBE19msJE/w2
YN+YnAGUDSpJXTvz9WHAJNWzSzZzhEk54Wk2Pc2k6ny6IwwxFdVV2Bm1LGzX0qqG
okHCZHyjWs+gnEOB1ky367YfRTBm8umrKNKJnaE4xGOMBh9BU/ozMwxfS3J3mBoc
kQQ/W85gdvcaiHUOjA+rU0Irg+iGfYAJSDZdg4G1cY5IsdAywD8KhcWUqyWUtQAF
ZLzCs3b/NWyQTN88NFeqCV7VPNS0UDxxnjGYdae/M79ZxsSr3KC0OAHP84jpyA0z
7BrgwxB5KdLKeNbafZsJ5S7gPDn5ex0sCh7utYyc9bmCHm8YZLzpTStU9hr7Sx5V
TRWeroRUoF5DgoLsNAy1xx4NwHYFsl30AE6EXhHMjDbiM8IT+w7IpKc51Dru13+H
LGLgOeNGGI8JcBhNenT4D1m8x1/MhkpnAmpYMt5Goo7eX+NSufILif4eGarjGMoj
UIcvqGlk1/5RqVqRZTNlQFaBrwjeYL49o22trPW0Z/Is7fPCn3v3dVi6yuVvRMak
0BwLO8Kie8L/dv7nPmqLZyLG86MKJ/mhcNtVN39gOk6gTJ5O2hLFQBaacGANLb3f
zE3/10fXCPjMPSKKb3dneaGmlf+5f9WJK0bIvTG+ouNq8MbR41RJd0gyEcxl74rH
xUb/uutgreoe4XjiYUemhaytdEMHjCMasEIPywx4tfA2gqEHNdRThEVhlY55athB
cjwJfpB7gy7EVbDOFAn9Dj6NIxqGOmL82YfIvTIVln0gsZ1BM1yVkMBTB5jvXVap
XUbPrX4hQK4b/2hZ0UcNuv8/relbdBX5InCzKNagMQWmKE+AB2ynHvfXmKMlGZ+E
22LYMLNXtaX0yMU5SfLDg+6O46nYTz+ZP7QJfDP9rj2Idksmyz6JU3bCyHv+wpPB
vo3NBA82STQAeHYkgvwFJtR8jh59NvuH+7BUQMQEhimMidsddO7bMouaIw7XI+ZC
DTjjrCY8k3cpoJe/a5H8kPx4QTvZWvq92zBERea1fLemeRUniYu5/aezfKx1tFLC
Yy/zENCLefYyXo/T6/VLHtiERPMyiuzfxtm8v02ueuKLgpspgQVb5uu6uRNo75Aq
LJYcO7lF7g6rUsNR3ZVOYmItGYuckoKj0p9qjuPvHFhbYRlnKb2K+Muh7NvAnSlj
OGdT0m1xJP68SZqxduBkmoeccZbXDC12EpIANOx6STdatyRbY+dWbKRYAMpy17NX
bHihOD9xZ6pLyeLLP6IGEHsRbhWEaSNXVw53DG2Q/q8=
`protect END_PROTECTED
