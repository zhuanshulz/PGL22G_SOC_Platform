`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UPtj7mlMEw5PhGxwWZrLIygWK0CZs6Q888zMq/0i60WW4NEfdOou0T5lCPJopnma
kI5ezKhPi2wdbJNNHA8LBtUakD+j3Cg07pZjdMYRPBNr57ZMlou1b4ngqoxLTq05
z+/yyhGUCkFrYR6KfBY0rJ2bP0ZQSrmeD6Z2qpnjjQiBvFxYdBZHkzgH53czBrLA
Io8s6uriKGqnPe22RbEW/k7JQVaBif5Uy1e0DdOpHN6bk8xoMa3PZMqfUyayzIxw
OVA12CufkKQcPmSjiNsKhxihpto9UYDdo0pt3EwELwUIf0LqCLGSFsgq/9ROrzmL
xmz89aj3826VZCr/By/hKniF9ljxMVVVqSMFsjNY/QyJHDuPNepbZKMO0oIAQfqO
3oLYCiD6fBZiQasOy0SUxG2UX1eH8GmqDjXdRuVHuiPFmTagmUtGPmL2RvPz/BG+
VaaR5AywRWZirQ5vCzp41QHKKLRYlr0xlCynodVn6NCUg4be4QUGu4Dw9JqTjwtN
wUao9akF2ZyZltpbaYoIpE8h6tKPi7m8FBsqfKCt1ml4VJSKAzSK747DQI4Kh0+A
we9ZxXhbM1JH81gXbIYg9p+aFGyVoIGV25t56FhChXVEHlBNTM06xTvdQF4Ln2LO
FqdAv3WyXbkl+lCKUnW8rze3OgQuBXtCQm/hCR44kU6zgPZaFaldtLIo6OFgjYUW
jrH/cG8YnT/wBnU9oKJjb4mgNWGcYpfcHPiazQt9FUHqFUfBZcZDqKmi/vPEG468
8dfEHoTAN/giIz15MHEBgg14myGXFU6y7qI7NiBatVmqtlOthQkX6kivKObfnFXX
afbgOm2qEHzj+NzLJRotOZgO9ySjERE+9hdImPsayRV4lUxCsJjVa5zA69ic9i73
se0mzLOqnCITkqunWChjL2bjQ9/AsftHMQU6YdK0S5TihjMK9Tm6NsBhpQmeGAWy
T7gMXlLjzOSmmKWXkJGcd79BEVbmzlvVpYHPXwJlFkn7U//nu/6/u58N3yLCKEfX
uUvU3YoaVJf8kO/qw/aObFnGfQu1/SoBAr2Ps6x7GtDer/qFJd7VPimXAXiu0r9E
86aPttjvdy2SJ8+3slPjGjHV5zp+EL/V8evqat8TTjMooUmRD7Z1YeKJ85lNrxWs
0KmhBAJ91Fyi/Emt5uzndp9FgDwzS25l4Ha1Gu1V6tTz3DeJRX4b2i83pCXc7pT/
z+pkRlu0Tg5rMsn7hxuAOx0083GVbdRJJR6Z4IbXklh/0GsPlWGX4TnBdpbnp6IV
x04MYxbgjMxVVhGcA4Zpm1LV9W+kfRfqc4JnGp6BXIXSaQuZhaFsi0aylEWwELKo
4jdQMa2oVV0mCuHnsHAD7ktQ0mkAa7vTM9+vt/VJ6+0JN9/aY874kabKSxQzg1HF
ZL/kS5NRkxmTHUA93SneZL6zvuO9ShlHOnp+oW+KJLrpMHxu+iJ+4PUmxmwH2z81
/HVHQe6WYYn5VAsP1yEEWUmrsCuS+YfgCEVCop3AmrvIDpeYMs1Zx9IqwVkDej+C
11v5t/eDkw9huFNdi41+Ga7SqoLtgYYfcP13XRfkbe1YL6WSlAoE6Tm+Ue0aGsbb
CPpgGuhdtUgJYYRdlvcreDzD3n39g9ho/N04Ls39V0YNzHGrtg0IO2qciWJl+n6p
yM8zDToWKNmHXn7SlSs7yA/0B3Cj5veUPejRBwMzmbEJNtvKxT1m4ibfwV5uEu/b
twZ8iQ3caOMk03QP5DatRFF9KKQRzFbqPBwZUMCXyKb6OucCW9xzlWzYXRmhsLdt
d0ag7k7KjYlpSebn9uK/lLwl+WuMVjiWexqRFOrYjIXTpX7eEf76zX9Kpp5BRHOe
q6/POyGjDSxzqXNtKIbCWTTg9Xiuuoo4uls0ah5EMBNW1JZ+zjaVXah5np7iwf/P
bIz/LjVEUEHrtZZduOQzdlLqmLibbUMpeFeozT+K7Q0NxW21KiV31rVf/Yl9Sll7
cfbJpZH9S6I87Rm3YPeWs+sC4H6/Z8gQT2sq3U6ULDevvz9fD0G5GLUn5JggvTHH
zjSpx0/7posogAVerCMvnM9uKNA+DwF2ILHLKjTmEC339bqHjm0IXexpQRC94Bi4
HJIYik7zUXoCWi85NiUFSbxqBmV72M9EmsJcoksexN2+mxZ5FNjDeDc3z8nBtcP8
9Q8fFY5rdoa191XsG58336yyB1OghyLZ1QrTGhodKRr6rKZcJhfQw2hgxgq8lIxk
JMp6j2AY5+26XagLVJve/Xz1U5KEn+oUvdsYunTmbPcyMwVsbkWRM3pQgLqdklvu
SLd2r1onTT4TCzSho32VdJqDxuWbNShYQ9l78zSLk0+XrtJK89lcZtBnqmMQ+T9c
hWi3LY98vLZ9edvap30swLDEhjHA80Jsr9x5bbYHxFXcJAuKa+xeiMu41cHQtymm
OuTEpj4/WJ9uJDJYrXpto8qoJskT4lHcLzbYi1kdv+qsVhqtH1Dmxo7GJXKw8sbQ
wGZdVnSK7SST7xhd1YfQjVeB4wTKTAJRlGyAXgU6WSGqIxLqkCXNnRADlNNQpAmV
ZfI7+wysxmvp7ZDscOPkYZ9ApAzm/mxCgIDoQeaOmV5QQTWX154vBu2rwuRYc7B6
pBAeMz3HNo3M4oFkYTGhiyM6e/G8xCKVzbjgYedvaEYjqP2M2fmr3iT/U7MMG9xb
qJoHG7jx/QpUfN29s9uVsIDFFuDdEH4opMtZhG0rUYRjnTh7A5TREPRKbgsl49j3
LYpyoSYivLCfbAQpCAMNFUOSB63cBj77nEQ/vFmCRoXZpmwjpYB0LuHOU2ihWQfU
U/XjE/1/TceA53umQ9KHwyblKgqlLagnbRlUi9Ll7Q3cfEwtckUB2xZIEmXSyWM6
TjODcCAtLKnCLr6ekeQflMDVNpDDG0bKU4S1qf0jkW2i1uYMK/yqLNH115jrXJTj
AmcIMDZivwPbhxW1HPLwLIPBA5Pt1kIChaYTm+NxTIsgrY4xHWIYHzV6LdSMWfFx
iSGUVHS7cNs5uNv6YVqoFlIWRv72Wo22fM9jyH62z3Rk4fYmTfH6QvTFD469Wbqm
y1Mu9ECmptqeDCq3T1sCvQeJvsM6V6r2ajWQsCXMhZelxoS0mJm2vlIqE4teNwBu
kufuR0MZMSKDylaI8xz8NK0pto4pKqIMavY28DKGkSzDdXG240hchcpBqFSebcNp
QAWE3rVHR7PGAQvOuMi3XNgZUWya0saEW6wEMY68/VehlZ1mf80kBfyxKcPighua
JVNNkogZEPKE/7kThsAHRhxe6aP1wul2M0jK3QqlBE0Hwp5RkiS8jZvCXLYzVHxe
paa66DpHadX/u2WgNu/8BsUJ6nqDVZ7ft1uSNTIXpTC3AfU+qtC72X0nQw9OUDcS
ruEnUvkjQTuEDSRx6YumI1v6eQESISd7bxPxTzxC9rPQ0OEK9I7nE9J8cfoY1K3l
S6vcQMhrEcN+Xi0dgXojJXJMCd5IsSq+3CikOSpfliThx3Oq+EgO/XTST39DiDP3
x4v1NAughZn/VfqbdNMrimEBNM7nM4TxeLqrfIUvIan5z6ZzrqJp1IGg7ZUQlSs8
XKoWb4ydCFAQFcEGdyncJO4pEO+QHqWMn3WcMIFfDVUo21H+6UHZOSn5Wcc8hlG2
gT3Dkz/qPjzoNvkj1flkDmYM9AOPDEnys+HW9Ois5ZlL0ggQ92XLHnqNVW8rL/mY
vsWZd4mv0e1sVXVDmmFb1cRdZM1yCek25IXSTfqNWqz4MhJGd99YWaVQb9V70e0B
DoZeWsA+QcybjIWYduCfNNA9kdigNzUI2TUgkw1734ColuEkP1rlZQvyeE/ls5X0
AgCf4SGTXVww0Mrq+l2aq0JdMW/BRVgOYTyR6KD1NpH+ICkIB6z46qYoHGXiEVfn
PVlTXb7XfsxW2V4LbzDuj2aD/aUdJ2zU4WpSD16scqHYkmZpYVzSgChmMBGtP1oC
jH9/g3sSwAM1Rzpi4vhW1nBJpzBq/F5us7i6NncvNpeZNGzZbIBz0dHvRgSdvJPp
3dPqcRAPwfGSy3ef4Ip9P9sxkvA2eSz59VmNsMh2smjkvyPBM6rzsvfhjFDMu3NF
f6ls01BgD0TQKR63gucRY7vcTwamfO2HQfEiELdQhcI/zz9t66K30PRremB9VuHR
SPynvBifNi1BuJTv0uToniywsR+Y1x+yPAQVLhHvLKSs0Rke4zxHQHAPCrnsSvEE
6ervPcuEnwdz6DJ19ty4qHhrwjv91qswfEGux4KEbfLFZKhiWL+iIes3WsjBsWkm
izOmJwClYdIM0JcJErotJFh2KF0JRk9mO6w8j2/vAVnizq0AiT8qv/To+ENeduEp
/+d6OwzPU2P1BqPl1d3hCcxTrFIyeaJUyzdjC4nbRU5COu8h9g0fU8che6kYXDZA
ZVNkhpbmtyoZhD1D4MJQ7oN1IxHRu7nA+wp3PH7bE4QdtAHGdVVJ41sdamcYPIUy
qZQum+MvEPHV1/81U9XUr94Ztf7kpNkJtrrCHooAYRM6+ZwIn6YYLimYWvUWEBWi
UcgZs6vtQbkonrP3CPxAnTsGGCt1DxhTHLGoEFIj60H05PnpHeCKqTSRq5Pd80+S
/TDC8S846EIwfXk13KBP3n2t0U/8pizueVsHbLM+sAj6wwA//qwUVAD+BDLVSjKs
`protect END_PROTECTED
