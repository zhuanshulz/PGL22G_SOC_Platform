`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jh4eoFHFzsFVr+FsF5Ek9sDuZ0KtKDyngRZC/cOyjYm71VDvVj9mRHCw0Y+zCAQX
A/ybzNOZS5ByFsg+PapZGhtRpY00xK1+GZRkPGqrSoz9ta76RdgRCDOGd1E0B0VR
wko5bpZc0bUwUuH95H/ZMWtgAhS47hyMz5NOlq9qz1rupgPFGjn3uEWa71xFlp+O
60TUuwsgwwhlSkGAlJ1/DIKUSj1TskLWwKRRzkdp4PAHbvNlfIJMF7u40O1x6G6W
ZUtcZJDCIHPo+OGfLXpvzjrHPmhNGL5WM/CdlMR0Nxw1EhsZqerowPfKxtWbyLIL
nUa09SDmLGN3SrtLtpO+CXRXGqbS93rpih0yHMz+hsZP0ybyYReuQqNxf2eFioqi
/OKeQpFr0tOxD3c+p+Wsq7zHe0X8b93ziFmf6fGEKATuvsWvPhsDE9UzOGEYJWb3
HRSfmzdyYMRJXRHaeXw4p9SFMSam+yKyVaC8Rz02Lim5egQnB22ZT6m7EYKRayBg
JvcCTUfVVc3LCdY/60kasK1Zcuz2ZWLpCv6QOd+tVDRtEK3vO6mx++IjTQ3HC39S
acSw3l+Q0DE5HRxuMy4ZmMhpu8X383CnmvYWkx7Us4hsnBc/NkpP19BKxLKRCxpO
Gip2+uX61D3xHkmDz6WXdw==
`protect END_PROTECTED
