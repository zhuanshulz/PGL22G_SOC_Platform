`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GM1Nz2L6WElpzg0ZEUbZP+hqNGFBVFYmxqw4ofW1k1zJ9iDmUDn5z3xFCiLXudAG
9BNFNqpO66SLJov3v+O3QMUawOex7FV1IT6PbEnG6TTllKSZjRM2BHYW+mH/Ww95
HRlRl1XJZorJhjTPhNHPUbAU9bjG9qetJq1QLODyYNlUzyeV5sQZAx8EAucNRGRh
UfSaPsJBGOK0S08Svrgp7A7/jWtbpXyGrRAXeNOKWXXe2AZRI+oYlDMdGye1KSps
SLd/J/FengIn+CA766b4Iupw9DWj3LJXO0ZSV4wN8YBxjnuCw/+Suz9nCTq3Jc5K
HIWkVI/YCqHkeq5WsRd3Or1Td0z4B3QwJk1EmQQ0apbI3MTX3asLZ5nb8zkqLPwP
4VcGjYQVNS2xLBD6PxPtSyfy+gTs/iZr+xB2VzRFoxTHNLGM0r+fQNo1DS04Ja+L
+chkgVLe6uSh25uyGfspBQolqI2Or++EBQ32MHzOZ/tA3S4Si4U/BQ6XKLdJ1OFB
zcCEM0SWrpHu6q6I0zdOEr0TX/6WRLxVkt03IdJbz6v/CStM7FG6OZxOnHn9pUWp
crYOBi/aqM17Ey8GlJ3wlXgzsY6mxFULLAo8U1dqTop0n0u2JQgvRGwvz6xb+fEW
`protect END_PROTECTED
