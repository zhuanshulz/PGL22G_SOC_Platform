`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+1oUmpIdXJT9dFERBbZ5oz7XQ5XcUTh3sjZxk1p3lAhbuuxLhe9iTyAcRMJuSUX4
aJpgVzggipHJfbzWVw7N41kSodXQGYCR6MYTJWQlE3bF+RKZ+jvUMW79JCVvyWpl
dzQgdjA6GKMpdx/P10uES5d1Nf6FQumPzfwsc+0SEGF5fu0cY1EscpQ/CbWrXeJ5
5B4AKLCMMT6M7Nw2nFQ6kvek4orQEdt1xWtJwqnID3nSa9oVsaF8wzPyw7NQe21x
`protect END_PROTECTED
