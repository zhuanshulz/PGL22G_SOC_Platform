`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vtn6lra+MaTEMf5j1UJ/9xyin9kj+FrFObfOXS3/wwOU9x+cq37WP0MZReMx2l8s
q+ZE2oNyHS8KLi3yY/aPSKEiU8Mudtm/ZJTbd9w5c2kh6QjJg0a+Nwi95iu9evSW
kEsAZ1Ssw63PgwU6bc0gjuxWKpwLaKomY6a7rFAJ4wTO+zDE8hI1Hx8HcoNV7ch+
uFNXWO5fsD3hz0c9t1+fWx5qUk4xbu5PTkk75A0Ky0ftv/wR20Uo0i1D1+/eo7fw
dLmSS9GMpzU3aZj4r9NF4JUdSxupzETqvz2QTyCJRI+xzvJs0/SMty57FfZe9zwX
hUcFZ3EN5qzU3j8CTIAzdbycl9Z9YqkGJNZbLNRluZmXbthc1UFbFDaErxvHTS7p
rBOSjvONIRmXIP99G99CwK/5OdyAqWBqJ4rkchpR/QZt2WRyiavbUlh1k73dHW1x
ohtpZm2cB0saM7u5d+KXEGavYGfDUtJ5w4d9fnmPXY67x3v9JarFlpenJxmN7eXP
nycWTh5iuu+Lnj4hiLokLIwOXN8p1WZGkVJDNSotgnvj+ChVCaYKMzVs6kxk6lgL
qcYXB/MdZz0pl9gTdTLmbikL1hhDp+U37IkSZinHjclOx12VCBYDNLquqPXVXN2t
U1CMp9E8WrCSCUeW7d9P2X2cnwlco+oKDndi0Uezl4T1i8mirGLUGBgbGm6Xd5a+
fgEuQj0eQ0tjC7zLpuJjFni/ZpO59fILwJ0YwC6ATsC3RDdSVaF5unj1ycrRAjs0
6ALufOUlzl33Ggh9Gq6pQMR4gK3sAWl/tKltWDgAxbdFa0437cRRNEsCsdDeerG8
LyBf056enU6V9VoMBq7WCZSINcjPEQ93IwF4dQVu9sFoyDzFIZRHnQnEuw67PHTW
E2/TqS+/WkJ3Ps2JipSwSQ==
`protect END_PROTECTED
