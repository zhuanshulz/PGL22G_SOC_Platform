`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xKWVYksf6mg9Rn7r0U1J1hmuX1kcwLl/5EhjRCUjjIeIWrlNEb1nDGqqfYZUBRGy
9+NO50UkMApOpVxf1qKM5qPNrpBA9p/tidDZAAvHAzv9mrVxHKtIvaF2buy0K4c1
f/LteCw3t9OTjmaq4BZhF0zqZdq5u2IxAYL5OMF9Ddsp6o5vWFFOK+KKkGUqyqm/
cjiDa2VG7Xi362ofWYILXAQFiYdjevlCFqgduk6TliOA9ZetZRjx7aBHd39Yphqf
v5IGI16Qf8vn+Rr0pyx0trrrfTgMSdtP1MCpXM1MKsMTVTa4dtu200k2wVG0ti+l
oWRWcz4bCv7jn5URJGPfHdc2WfGuzyE3M8yJ6DvU57f0RCEtvEssMF2WoI18iw+d
nmpsDyfOCgvhTmGCwSdjiKWZ5bSf/l433a2ttJcqPbF/zcss37OFK4kIcb7bU81U
UrUXC/3DjxDrDZn1cPhXvlE/EAT777t6FVttLqWAE/g5WndOvrt9LL9tuAmqy29X
qOTOcObrWye09Zc9hXaSOA==
`protect END_PROTECTED
