`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vtHXdSqVZwuciQnYTAC6P8eMUTzeqlHTzlne9O0q5ZnAyqRcIp7mhkFEIAWujB/c
8a0hH/rC/Zq/g+lik02k7r8pkP2Pdc93/vmEcqxNPJ40WnweoxZaciCKIce0oKoP
HM35ybvY8i16qNE1jimjctFST76FeTlS0bPj9lLw6QLsfvvVQ3gZGZREJ9URYmr2
+7mi7ylQwZq7jd4sezu2u7bOhnCBHrnR1N2shKwbTbAc5zhMZcIkHgmfMQOYUMZJ
Bv/RE8AX5Q2ba9l9X/mjSksd320k4L+LCjJR/hIRtPNo04ixd11d8qTThY1/aEQ/
zbM1/97zqf0t+sFBGFPZnUqIEEzOxBCO1Ee8DqKKSIhv+fMiN47CBkwgN5ieTQIW
uk+rtdry87E5dsfZC72mWGfAAceL+hURQ5l+YtLgC7L6SWa6/FkheV2NbMu4cR1e
JlgwX2H/+UJcDGjLIC5jR7doWzpUdU99N95VLGqfLS8zrddh8Uk6jSuva7vK6ZjT
eHZuGIu19Oy8bW+50JfOO45bLDBq2iMFfFJ2l/AP0Kxzkiz5WMPjDVwDf6HeSGQ4
/7D81xgPmmYsxkfZzdahE3CJJMHlMcKnn5ZOOqsRhAtLttHJlpvidCWN9qKPkFm3
rxXYj+DRSCOMkr5/dtq9RQF5qCxhnZ+PKVr9TjkuS0lmOn0tNaPQpmF8+RrVwZcg
hhGZBRT7w9R8zp3B10rqgOj4BZ0Y+KA2MmCBg35SCWWeOkwkCYmuacfGc5VbCQ5/
z+RZQh7RR3YEUiq4FSEIeJWAJWQtBs31wdVuwsxbjAoVXjLjpZtTLd8rHNbgHDW9
JYFVQ/w56D1vN/By4WOwJHajxxFMV67rPu32cZcLxHZYuORwsvQpNQ479vszMomQ
yjg5h/BMfnlkDaNrGRpnRdiF/YGKtmYHwXiNylJHFZ2TeEInOgM6uJ+ykjw3vQ4w
rv1LbxAyH7Ula7aoFoSPMPiQEcoUpzEQhAaRQ972qirY9nVBl47l4CRKnb7MGixQ
fdguvOzZEHg1KgX/akNbFy5y6KAoKXm8Cup/lg5UC7gxih58BWr0gjPUH68ULouf
cQJtvVjqvYkC+uBRQmtteLMM8wJYV2tIW4CczG/967XByHeU7eIQ14X8BF1Rul3T
Uxp40P8pZgZMzXGck2cRYt9NpSZ/u1981y2WAYHY0693YUS8yseoP81pKZiXUSgY
Gl3KQ3tflaVjO+GejF07q0Q2n7I5c0cD466shVLJ/XyiI3hGh5xYbcE8PQnUsFuS
n6cRtvXKJuNasjFBDyBt1v9oYWtRFx3WN4pKYrTv7FchNQCsltgBuKnKoCtk13xu
wXpdes1X72rOr1cnvXQU8uK3cHHUpkCMjYMnc9oUtIDX7kZdL1TUAi7ktdm7AeHz
An/9gE0GnUYT4Cp4xYFxKBIM8+hF6XD+ysT94euzJnd65Y5FGClZ268phw/u2zG5
P4ITkXL7vMt0d3vzna/K95qjT9Eo5SR5FA9GjYANLH6jb293UpYi7EhdKRq0Tbc6
Rp7mJN8LsceD1KIoAbW9bEDyBwoFbHZHNCPfklMcdIs3CE7TehiquCr3IVcnIj8+
KdMlHm/mWffQ4RBRchV0++aIjrY9yhq6oJBcEmuC0hsrYHXnfbJBJubxxbxQyuHV
4IqipQKy3YMlzwvnRGaAkZUCPDjoar1EaGsrRqvc9X7MWtDa3K+Sr999dOOFruME
rquFDdFcgoW5cDO0D4SHwQc6IA+m9rjzHmw2+HuJBZuMXinLXUhBi67sVo8cfQX0
7wv1/AXwLZeqLW9APR4lXmog40Gw0Uz0WE5Yp2D+yiBFh4b2ep6usM2czWGnORxB
Crk2zi4vMWyS4j+ZCBYrcMo8uf+g+3gOYN1t422UlsYQCSiqeVmfw4XmxRAq0FIU
hTE4nVn8xHQvnyEax4+VpyV7L56ndGOqVrYCB6okbf/sUQyc/MNDWIREyAY68y4q
bQRhSlXqaPWQPWeRIGvzDAqkPjt4TW+kWi/Yx6EGz0iCK854n237+u+ilk9Oq/K+
Be8ze0c3NK7e2sKvun3PFWUTaMmofcomcK4b7VIhit3RGR52HC+GbhEZCtHsP9WE
SBB9VO8ia2qIPNDLkTengJJ7qdUqPn+zcu7dRybZHTwfR6AbDKFZDpV1dcq/iZxd
8AiRTLt2s9GYvA67Py0drhOKii8sVoGOwrQnzFCocMCLdYA0sWb31yaWbtiDvNim
Ja4ZVC3IqrNryaRHaBQlsm3C1zXtCLSKMT3zpz5ddGugaEkigjf8hJdeIRqcnGSV
7mx3x2lpoKHvSu51V5exaUrBK8+PuzEmvKbkyVEF0av2iG0SvHE5qAGLcDpU1/Zc
bZMpto76vAi1bZY8T5DzHGxrH23AAcahYr8npAbxeUMJt+rTUTzrqY43ns76ujdy
/BDMVJIfVHoHv4f1NjM8odEYqOmc5n+ERogvZ68PtAmIqxTChJ2/3/7agHnglX66
ZR8+jgcDIMQ9/yMEXlSOem/OYMe+2QCNdhZiQqyAANHgRf6kc2r/88tK5PmuGTVC
td0zfLRk8sl5kbVs1ySzj4+wmbASB8pmJzY4X5GXESb92QQdBHCRW2nFOunzlyCf
q051D0nLHSZdY1ZDQbgBLTxKOI3j9Qm9JZvY6FLKgrZDto4ChGUGi/VHT2gsHu9q
4cGHxCPu3kDEsSp3m6Ym0PPLItZKkr7wkQgi1oTi8ti4n3BMpyTvr5eZQejUXaSK
gRmPlKt0PK1RY6DP8SZ+QFYeuhddqwc4heIiJ3dH4RNkdUlBdlHY8cwPjQH783NW
UIODy4zCcF3a1sTHQE9HVUg5pyHC/uR/SUf04xAIFk6hCksqYW+6VlwU4slVj5xf
tiUu6JQAYLEhFjFAp2Dy2DSHaLtI/OOYCeXweCiXknObmbWNUJWqnVjwk47hLgVH
8w+Qa5jpfTFofL0OSxUKTw==
`protect END_PROTECTED
