`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MkW/d09CFe6/vsmSR/OKehP1NvT3LETxV4YiAhDqHmn+vakx0l2p+zgTvD2G70dG
KdTL+U8MxEhEx5LxPM+6hqQoGpVjjNSbyoR5L+2i4OYwEu1KDr2MThd+aWMG97aZ
8VvBAz3RMX0tRsSULgX8zMt/R1yNtmnGwLH7RG5rvzU4Z261qfReYz9WNPeeyglO
U4J2pyFORGRvbcIPnFH0L0DgQ45hU3q3ZoF1dvOu41jj7RrleKU2vvSmGSH4+EmE
CxU7Jboyk/qD+1SNE+B0cXTTkmZyRW3BinGXx1Kn3gDX9BW2b+kG7H2fwHdt8ds1
s6xHakQ7F0rkZbqk2reHRna9260GOUtlxh0hC5zAQy31My2THAU2iBgBvH8cSCUk
Fy7UgHbXFuASyrwgyrKOCJryEWzaHykrLSPp5B+mqa8rQlrUHBjrPXx2AhLE1JXe
b1+eO/WUvc6mOYTMi8TfCr8wK14EtL+ZoViU8CXI2lq//tfJxNaToXK3LBSVwCnE
7NWUtLkW/qh/9O89+/gUws6CTCgU/zlcmlPy7xYYPAmi66jRsaOkjV+bi85LtBuN
jdzU0Ni3//wjCTgu8ZQK82ADZSmK5kWavBEytZIyrtKIa64/XWcg70ytaknlFDzJ
I3Qpt84ftQgzh0YnM5BdpplGErfygV8NQ32+HOSHQ0BnM/GowUt0JrAyosAw33Y2
iWVQGENNne5g6eytfKpXnaG/+1lhAdJ0Ovlx/QpE7Rfiyaw/9bdbQ4+XrrbhBjEI
nJGsqGz4psN0hmociYqRa9ilyaPCFUHKTL6zMge7B2c7RwJrarRKnUCm3jumMqgw
OpZRDGcVlLCAnPFLvDL7QNHyWgI3InuiI+JaTV2GlmzH3yNMamApbCYQbTomskCh
IOBEj4GjGIDAic0IVtHrCicR3jq6rCcEd4ebzPXSj65lu712XQDpgqsmo0xxTlfo
ujcQ48bWHX6OLkl/K43tmR1A2IObSPMxMjfcgHYIJ2GVUEa32gtZR8RIfeTMWA0N
og2HGy8h6Jh9GOzni8JFel4Fk+fzt8ADHuAzfpg0nKSutzfM+ZAX78AVZEVef7Sg
KuwWkdq22ZdqobDuowryIc3Gtyh/Y8rdXsIaqF5VuRvjfmgqIeN2L7LFQnbcqG8G
fJsOCbRyVyBiMVB+fyn+COs+Sb852MTVDmNC6BXocIyGKJpmSZ1zD0ALlG7VxLKH
NE17f1IRxWbJnwUAy9Hu0JfBgL93atdXouHJUdLSY7aoNPSgTq1PBwFkVSJqnq2F
60a7ittjUhq5KIXvTfwMdBtCPt8/c99I01pvsSHVJNK4+EAlWdoE9CX3zTZd9cw2
xx2+Mvolk2deJAMovlFUgYa2feR6j9KFwEvn1QO/u3wYYh/Kq8evYyrUO7bLG2D2
75ZEXEioJ18CK6D4dbir7FOLiDXb63y6LXpHc0gMtHQESwLJ1PodlOIt03PDgwgm
evZgKoDqIVy+iemwCXnrTLnA+DLuJhFISrbJkIchr3R70fc9tcFpEMavSK5xbqzP
atncvehMUTGvMczkBPxtlcNZxpBM5X8M/TdNhXBM/CJnpq8wulQTnVs2oaKA+IAg
Zii2hrUqCu89oY2056nRjHzQlx8ZKRiHEBHE2h8RIWi6UFp178f0QCHT9IR0lnI/
cTrIzoXIi5zylAF/JyF5Fpy8NUws06W63kVK0gwIDEkMBWHB0lRYZi2VbN/iifvS
m8zfn+z4KQgDZJs2EwsM1Ynw4HKk9p7ZNqNyGqvemfTL6vN80Qm/vTcSXdf+iJY0
2x/qnhaIADvgUmASLTFoMfUeWiNCNk/e0ODCyfWeSb0rd8ZhyJkIJYgGW+6Ux+YU
SOXs+d/xgFGtPL4k766J0VDOlSl0Nyqh1/FXLgZMCYqHX5oXXazHnkyXJKsbeAHH
PI6nKkHzicDC2i5QzjhTLoTXtvUQinxTLlZonRFaxNEKigY3s9ILKlVQ2fTyfvxO
IerJFuhhMTrnMqIBDP8uHA==
`protect END_PROTECTED
