`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C8EVoNbaOE/59tuk+ILkREhENLmt+XFKCi9LV853QK+IhGXV4nflDEGWOet5lBtn
bRyNo3mBoB0ylKPT4pwjih3kWGnnr6N+1ptikiqEsG8jnkgo6uEDF88uI5Uil2er
B7KJ7p0HJiqS7ARNgALuozjJRe8Cga77dDkp0n4U4PQ3GpcgbCYvaqpth0EV9AkJ
9s1wmUNbuWzl/iTOd6c1chn2xjQmEjo/L5juStPoxTE2yGeiVpd2aJ2LXIHGGsNs
VbGWDZnAewRZ209KIUGiDdEbXp2lS5Crx57lrsw1c74JexyFwB6DeLyTL7oc3jel
8ha/Ru2gl3KAWv1THCFNI1oLbzt5DhLOgGGrxWU6cUXTgQu48jwVtdfLjio7csm0
26xp3ngmoCclraxCxowYpIi79OvJiXCQrge9496TOq106py0mG92ZKYJfxYS81nK
ANU4DQtd0rpU/knessdtyFNQzYGfzDMthBuAxv8+tZECZTknjVp0vX6b748f9k7B
K57WIjCNrGFv5O2pfP8YjOrk7C/N5vHOcRgQoksZ1GzerDCMahkxAp1/9a10yyvu
oTMTlsd4FRDvmSzyL8wfj0QRsavBf+gaYcIjMbaHZBXXq2KXNHq31XHuIaMumVdc
aoKn3lZ4gYivd2Bdo7IyaWKI1PU9rlalY+Dl9/FrwAOMRy73IP6YDGbmbo5mXaiA
Q7EiIaZbG3Hmrb+T+x/OqLxlJoWPk9kMU4YpfjA8W69a4/nZyb+Ay5XnPYbN5XGR
cxOuTzQ/aRo7FGIpzROZ8w==
`protect END_PROTECTED
