`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
76G5Wamd2f4WdSGH5VVYSUG9kMTsKeCw0W5dSxS+PaUu8qdFHs+u7CdPGZEX2yNf
7ynQ0Xa3N6ZuJeZNRWYwEvor5+RBmjinkj/hZDiL9LShFmYMnXDcpiITjy4im7NJ
sC3pbmw1IdSW/Z3HpvWFcF5Dn21T8LjaATuPtklJA24XKqjiFWBbu5v9LWhlv6Tt
S3+2Mtg8p8cyFg8xbMJyiqnWzuOM07KfD7lEV/O7rmukhYJFfLK5UFc2D9eGsylW
16r9wzJGJfjsDflKCHXkTWBxGvza528we8GKvInZ0su6tgzj5pTHyPzQ+EtLr0gC
Rj5OUd+0ELOAtx3BFDWjCTtdzrktO5rljvBoxEgjZGiYZfwhwoHVF98ieEhXXXc2
Lz6jcgpntqfO9zTdLhhXGqpSsEik3LSy395k1a9pWv94mw8aG4FfloJYnnP5N7qr
O+Pbakaol5ILTY6D1xLiap9SnFdqeO50efIRuyk+WiUMOnjYjrezb/Zj0Ri2m+dz
4wf3V/sueak+I2+Oz7oKyg==
`protect END_PROTECTED
