`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vdUfJu+t5qOHEyIJo8/zNxpJSO4+XWWgQQM08elAJtNVR5gPLTrasVWmyOLXCA1Z
JIX53KcZT/0HM6aYw6OPa9M/Z7Pc1ylaJrtXn1HbprWZn/9nhg8BW0lnEAkl63ir
o2n4nu9r14r9C7QD2DJcuQcqjD80fA+ZRy5x+mc+yLcc4Yu5333c4IwKoH+xoBQx
GCk9MCsvsmDCxKN3UCtSe+Kn02ry4JvrN9QSSF2mEmlsU4CLBsvyZXTz0oS5WMNw
FvdzBa0X0qAFMrygmHQpLVbspxru6X+hZpUFCnIBo+hgMt0YRxIjtur40UG3s6GS
s/mKeS5c3Oao4q6YLiRddw1TOG/fYgVwrfL/PmjCLeJ+zflTOvZD00bO2bg76OE1
s3M4SmzUiPRjIX05kbPMToABP8CBqqZv1wpU6PZtPhZVmAPnOINGOnG0Tj+f2xJs
v7OQU/nY+o4B8YwEczEGi04HZ3MkcyEf7g6arYcrcOtyGwpTGONJ5FM+bC5zILNE
H3oKkvVqRx5oalRTa4HOdKXoGYiHZlrGUkyng+1J3CX7sPHWRDztakUr5MvdWm0t
uHu5+OdtjtmAcqfZ/y4oj5H08GLwcebY/4yXvCCbv07efO77eth8OAfuW6X75ref
LuRtbyIs58kOf5SUBvkuSZV1IgoLGY0o020nD6X7CoP2s8Iz5/69wvEqQChSJdS8
+2WoVjf+X7vS/IgvAuhiaJ/H3iCcLzi7JM6EaP4Qxpz6qBGUdkXcMcSTnpholPoW
dGH1DQMe4Rn2XNMhgFJ6cQxoMNVrlNl17YE04iy/491ZF+xyrtyHn0WUlSUIX+9Q
mzL2LjPfLsOeIzJl5z14lJsweBYT7r+qOytosGYZbM2g0f6sBuAXfkjiRbOOZT59
Ym/RiSb6/UWOVgA0A497uRhnAuvlNrwdmSEFb61KX1dc+ofZnQTbKFrXR3S/Dwsa
/NKyLV+VVWRmp4pyAegDeVE2/z/I512ag0umXmlRD6g0Jj0sQ9BP/zEM4pDbKg0C
A6eScWMj5CLvvQ2wW3Fv/UEBQzjbZhsIHEqum7DT8ZRW6HoXLbwgSeBffSPMdUBg
sa22owpGOHEdAY7C60ZMkmWIRZhmnNQigEgXuwcAhGRu56Fv251OOQ1ZMaJX2F3T
4E5ctKXLVsAU2/QxPCxTF0wIZxWhz9gkXJ5PJQs32FbcbS8mHerOK++Ey4TLoU7E
FzmHMF50kaoFtYUMDINvaEmCmoUoNOFM26zl4OUDH3QLaab5Vhq+hVMtzyP1cif3
8ehad1ksYfTv3nD60L0KHE5Wg5v69ho+UyVMdFkZwlH1dTdfs/Jxmr61h4u9Dh0N
Eib4m7zDbtGl5WrQD6cPmGbL8DWP+seCiiG5LWpbl9+IPOxDmR07kzE96KrgqBq1
r3z4EZDvPn7uNsvfir8aahgRqV5gBJn+kKk/6nDk6guHqDkwV9aoQZezq7kN25VS
zsNqn/6M03sO+6WnxILo4PzcWKyWjAYOuZyhuF9zCG1jAnl2cJMHlPXRtJgZvMli
iahvxm7f37atHuPE+g+koQpSKUvGNlQpQ7GELCNPLelta6IfVfF3jxPGjeW46mIC
no3hZambQEXnH8FkkjnQJzDEceokB0Y8Q44NVXSKGlYl6Ez27CbZ8W0eNWaIngIZ
/aJReQQ7k2jmpVkj7e+29fqt0CTlLq1meyK8wvmT+oqihYFHhd1sLIMNm5G5aZna
Ma4qhlcdn6w5HWzRM2DKzZ5nSKb3Dx6m/D4yMfVyIjaG9QiUiZOH0k7XRHAoB0x+
OaOfc7WuVE7a9aHF1WtOxPEWy8e+GEMXjx1no4nHSjDqtrHqBZTmXFiIIEbcMf31
ynVrnUX8I3l3et9zduS1jFj0xbh1WTZ7JwlCVmxgx3k0zpBmsRxABk1pOOb/UBnu
r5Tadz76F2RILm9djHcbDOxhp7B3MBJEGVzUcjVTKqLxtp1/suPBAfnDOmXt4umQ
e6LjElGFK4/ELqK03MtecLcWK0sCUOjZP8IBIsC/snOkfN3woTZNbbEi3sTiF5bK
EkHEsV/ZU1dEslTimmGsRun211HqU+nURFPHNxs04EWmpIBBpf3Wkbld/g2bN7Nl
YBZXl6rmDph1zUoFpmcfQ0QL6WSSs+wqz633bHYhTbkffa3zihjiR64xYNtqMote
4KP1iFObMuy796Zp0Wp996VC9l5f+OiO1UBe0AxFhO8a5Wr1ZGt4EmT8NIxWN2VY
VS0rVlxfNMuvkQiRv3NY3hJgwxYJsx3mTdJ709wIFKi+fnXA9d47xWHmBQbdfOUB
S45yIMMuB8gnNBjqovCkEZ2BmAKTHh5ebWsVexU3st1vWN5kYpUWsi0RSVKxlKeA
ZS8a2PY8J7hdXUIfhXd3cQeq68ynVhnRxrG3yUCzAOXG1hRJ3e6rNrDeNbAwoHJt
uH5WIEkeDYOxuMvuLctoLJAPhyBxDqirjb1Pw6z3IaItyde7NUZTc2TXU8CphvYw
knoEE+Z+nJrIaUUnyxS8eKTcNm1hr5gdlowwf4ohF5A4agM5/TReXQElsO9DMMOs
FCYAOZqc7t97ctxUtyuVDzj+IPK9RIXlveCXb8fFyH3bpdrbmaL2YISXnpRqvoeI
aVUevOp0hPfETplmvzpLhJ8Ml4E7vKkvOooTx5IlDUdkOUP9KUBy2oa91UEF0ugw
TUET95YXWMUFN5hsm68r9MPgfDg3qqXPrhTab/+RaN6RLVWS27JrraCytt0TirpO
s6j6/4focf+b9tbbgfA3IOcU7SmbvzNuEi8UaAuA8gm47dBB+SOffPpaWyHNCSRM
Cp1QDZHJ2R7iv/0GPcyGmz2X9UaFN4I4Rki5gs3I5yBEF6WoGa8WTg5OR7o8sf5a
HtMXoQ2rEtzS3yJBpsM587aBnWH7cstlSwhTcluqYV4na7VfNo13BBms7KU7D/Pi
cpzCVDc2Qxj8Uwml4gHulQccb8InqaE0ARQIpVBrh4GXuNmRH+8qgv9PXko8F4x2
OmnUTYz3PjgEcZCHOzJcpmyT78Fu/2j/b2pmI/TxuQn2mzoP6Gh9HQy2JBRT7CEU
v2iiLjG7IBzCbPUJt2vDgIidlT1ZLMntI61mCUqaLXiUOtoyg2hiX6S3lmmgkVRM
BOaODDjAQzC9Ndji49Y6cKxTyE00XHmIR/IDjCGejTCiRhBO6JjMYpwjhba5oqVi
0NZ9SAiBBIisK136jqsrFR8eOfKgOb140Dlc/KBeOwUzIgrZ25sVcUxjW0exlFl3
nXa4Z33O3d/rsrZhay5TTR4IBsXlfYBWnQ/t1NDN9a1kE7O32Qb3ew5dwl4aAHNV
Gf3tatf+baQt8+lRW/7XuXF3FZkQ1oW5T1R5TNNTUeXhl0Eyyjjga4EidzjpszMU
ZjJfoiDIj/2zoLd6qpwS5NGGgaQ6cbHzJ++U4Sa6f/4izsFKpfuHegbZZhcOVBaI
3BdPYTNM1mTQLhA4dxQedBwmXc0Z+Ks7sKu4WhmmmS3egyAH057K77ERZ30tG12b
dA4NYv5tiNky7DRW5AfsA9FpSmA95/lY9WE8WeRSsfvSBvVnnmIvZeulLQBIiyTa
uCVs1ocm672awbjaIuREJKqpijhUxjtvy7CrwgKsudngTo/HTOPR0g1VrTTarywX
UtVJ4WIQRj/C/dfsYWK/g0bvPVqgn7bMMawb55DzWfTfStFRmnTL8Oc2XIc1GvHZ
5jc78CyZLSe8dxPj7OjbmVP7EITAF93jRf4OyKJZ1/9HCFze4c3Vu2FFqgGQRwHE
dYbhlosI9R/iTbbEYa3FFrdHqATItt1Kv6ptCEW/KaedznbTFvhvkxF4xk7/zMRU
XU6fSfw/vw2PX1n6xBxuIIZzBQDNMnVNPny3p/Kew60nx40LfA1Rxi9fpEGsm7DN
1aNwZ0WD18279TLoXC0MmhvlYTwVsX8bUw3qpzud1A+HtUHFGy0IER8ymJmVFygb
du1DbQqoAW+bU2B/QWqt4O2enFQLJVMnE3KjQ28/TDIUBdW7p1NUHGhKMh3vc6TZ
1sVQustJhvrQYPIr7yW/iV01lfvRcvT59Qr1dwmFlnBPi8NkpRhfOn86e37at/Ng
aI92Jsx47hmpgrsxRosGBZ6bHoVKxbJrHZhBrDCFPlZxnsactQkDwkmPQ7nbiZLQ
7iAYOc6PnsPwPRD0YqnWGgPV+cT/t1+7C9mO4DriuwgqEQtfdUz5OGYHHw5n4CeR
MIpClN+QhDymyyNYyLI1WHmMb3wDUHccw++VG5Yy4+DxqbB1Lj3GdcM3eZQzj2iC
RVIOVPTKlZ/PwvCFG+uU1qXO5Wf/HW7gPNk9o65WIcAHiVie/ctafmfi34Zdiw7j
FYCk7+x9yd5Jf3XKBtr/3lftyJwGVShi7OojS4ryTYhBNC0QvB70GLiYesDC9aua
rRHUlNbpcCymyitW/gpZWNuJZHrLaLFfCUzESFtZe8s+fUue4gjhWrP75pugPIEc
XSc3c109qlZq3ZPgdHNjbt7PBlxpoblFt4V63hnDiwDCdIeqxDog6gkONQcszxNs
XPMrSc1ODy0FfWFZ5yppZ9uUJbMIM2oiqAeKLE8fNNv81tfmSgXySbv1tEgi2niS
OMKbBKdwry93OsOJg/o0j0NRYem6AlvjuH7OEAJwx3I6c0ki2jHybW90h4M85NU7
xf/pdpy33h4BtdmohfCoYO5/SoPq7tJZVnLNoRXcVaJIZYpJHkIG24Pjp+4Dqq0Z
6g97UHMhZvpYkLifiUetJOhlBf0X2EUfoSMlSWGV/NBKg3QSBaPLlK72tO0hwsmM
ioeZG6XPft0z9qoMM2A0MdO6Bx0TZg7mevlnIrS7ZLu62VlIGZu+LGtR2arhGBa9
MT3AIOfzkzk2/eQQM3ZTofzB2CW/FVdhGJ+bN/SNTikyRmmxGn2y8xEINoWP6Z69
kVAyO7/Jswsxj6DRuT4AhJ5VRDNxW0s9O98NAKwk/5LuiTSxbmlq7g5BX7DRF28P
LFvLNgXhK4/aRVl/nR1BcsTDC++5IanR+7yxcF3VMQY7IEWEtvgu5B0QR6FlFE/0
gqKpx413dV6X7cr7NeCErHO2vmpHrWGIKuEWWJuHdgc7XprDBzRQt1ZMFYeVtip5
At8c3hdwhkbVfN38ISj8nRPf+Q2eFf62LSKKyp5AScaQRnnT2rKBpzfGhkxjM2t+
qe4vyNSLwYbAoeFhCAtrhD9XxjO9Q4RL/8wsrRSVpCn9x5Mq6/JRDKvpcCTlLOdE
JusroIrzekZRSO/AIuVnYcdLDplKpRS13Xqu/EEsNy9DJUMSChv2sTb7Yiv1Qhy2
ICgjUmBzNpRXn0yTQCMO61nLrehFil2bXms37dne2ZQ16IlGZ51RhqjuTvY9ZWZe
iqj/FCrwjEOyrD1eMs60uoX+zBBHP/z0/62y63yDRSv70oHygmk2Eia8b6bcE/ut
8qoWQQrSQQX+XK9rugU2U8bqO2EF+YfYHtgsacjzQURCmmGO42fgHDyO/+YarSg8
t9Ac7VuK9hdHyDad+pklDJ6Tt9F9ILDqn7xf7DDjuEjtEWFGbH1q/9+RxuirUH+a
pj0T49ec7b021ZnXgXI503NHBpW7wwYHzlZPShVSq4wm1Zmln3yZv6Gtx/uDIsHu
+bAHe/RogE2hyk3Ge0yj9ZnLObJvqBDB7N23anuqmig4S2539pEdxPoDp/Uo/YYn
x8KpHQP7fkJKXEL2WL0wp5hi1yis1m4nlJo5hfDj1qkj2xqKD48fX09jZu4ppHbE
UpeYwMk/L574qjVZdG5J17aeP4YuY6DE1OghsrQlADusnZB8eHqd6+F/ZwVAK8AK
ZjBv3Prn+4s1gAxqbZJYo6q9CANtojtHUZGpvi7ULhXEWGLwAcuebYkghCR+gfaP
hXQ/OQRoDRdOJoqIAUghpk0DOTUvDaXcLhR3IYcUUi3EaQBodGh/7oHMLfOLpiuY
rl2Vx2BFJpW1VgNG6of7izxBWnH7ncSC8NpvcNObpOrXD7Sk2D8McYmkLSXHABMp
vh1bkgH8B0jKKrtPyFCxgeEN8GfG/Q4u5Yj5QqYTg37rygujPjzo8Fw1nwD5+iWq
dFDPRuKBQH2M89ys/efb7UOGiFu8wnd613y752DbgtKBvPlLYE+J9UvsNEKZOqmX
iWggmIl7x1lnpymiSk4QHvM7aNsNKQBypB4qEIg3QRe9F4Zm8yeHgJpqi3BQtl+H
ixSuD90Z4fZ4VS7OFldK8RngrRO7XZtwAAThpP84+pT2uj0vpBO2PrGGKXMxvMxS
0cQo13TGGdzqNQCB1Zr7Du4e6oEQNsBhWUybNcrTH+wz0TFln98MXfogWMi1MOib
KTb29ACjrP3MH9YaITmLuw4D4MKHxeDXY/PrDRZskG5b9vjQz8S7eJjoUslbOfiQ
iniiE4KRwZ5lZph5Xxsnk5E+TuJyJZZLSiT1CxY+FKLoD43Gdjo/eYGi+Ni0vjEo
zsTpmrcimpjoVTqhgi8h4TFNQW+Ric/neXfzkFo5065yMR/o3fWXVxE55EFOKIj6
h/CaXGU29yCndnSh3PYffuo2+cgk7Nv3ddFbys6xiTeLKYcBcNvrUM/dQ3KIZWmK
qEorSrMdo8smhWptdNQcAIbvA9c+MC+yNvXEXDpRIlW8OdftAQK+JDwFH8sev4Kv
Pjony8T4QiJYqeSOZ6kAXqry+hQl4cpq5SpCl1O1a58fmOeVk7y3+8m/nz+39OgS
ataIRP4NoFTkAfAV+z4q3PknP4j2ELQeP5Gpmxraj+wZWEnCbyxBpa6YVazUnZM6
a/UX1npjwIX9uT6+fr/6vm9s5jz/OO+KGAOp/WQKEziOhrPv7jmvkVQedJL0KeHu
QseWyqQpXQ4I+fdYcz+6MTxSWhTep9JyJpAbNqUI/dundVPoCtkGhUDRMseDTiq7
naYlsLojEniwASc5ZSK4e6RyIH8ulyzKoXTEf2IrMku85WesRNq2KgN6pJynnR/i
W/lBCkBgUo9kH6+7mcgvTAfBHNtBfXfBQVGcXPgS7F94ntRLPxVYYkkAm4wlAnJo
Zud3E7aVQ0X/GzgeKWmY+Z9NpmWDpnOVTMumN9ri/jvLnseyzeCYOnSc2FmLnBzt
PglmYBpGUWgTNoxHO1NcyGoa8yG4ZnnVw/JJfN+ghzDBfvnRveaqhvEGTzLQazgH
Pz31cPNjcVOr+s+32maisusTwlZAy4Q83ngljYZU8syMZGVJkVrvzdnHgyw/4BeL
lgQhEO4tdCdHHGdGVovjOp/tuL8MXfFMP5C0/q63egmr5R56Qk6/y60Y+RN7jVRy
v5PKYQWJkQ1KK1V4drTJq7aZ3zuyaUoQcxArF1RJcvfAtW/bWFTn/eSFliSgotUL
KU+A56d7PepSpO2DUISvfKxPHTiTVJf/PcyFdVUhT3sLtjT95zKiuDFG1erkXGUK
jt7CPOLT3h0EsFX6CjvCsS2TFRJxBmaz5omimNLIp55HtwMzsrMzRRHocy3fYc6E
yFQ/9T3c/W8dYN6AdqeqKMp5/3Lizql0UMpu/+eHtVbXiQ7cGav/nOTipHJWagd2
KRwkcMLlXBUwL2YdCmb+2XNUqqBhtEfJsAZxf5l0VNw2E+bxA4kFb9FngzXpm1U2
mADrZYwPP8hxiI7B0wmhW9xpZ4CUzg3qJ93TMWa0kITlBP3sa8tWIaB2YwyhQks+
fCr3a48/3W2NXa3s/90tL2lQxvgS64BPfZP7EX0nCokCHBfHVFyo9M0fxR6uQtbe
bxv+JHvto1K56VQCQ6X+iGFZR5hFxpTvfVIkdHr9S7XMrGWyj2ECBA/GigAokK/K
0skte4gZpcdJWy1CPaPjmrgqEDUAs+Gkn7fVXz0D8z52j3Jw2jnC5v8doNi1tffs
E5f99X7pqoYLbYgp9C9wnKE4tuXEV+G9cRxwdAD2/lOxtU3XLqXE/omiRA2MIzfl
fZR2GxGGC1XOUa9I0C8P3Kwoga66mJUPKF080UoWYYe8KlEgMP6DydQbN8JUYBgA
L81f54lyYr+gqfu4HcBoUU7uxpWdCXLr8ZpZItnp0V+0lxrBd1j+9Fh8YMSs7TNV
mDYAsV4kXDL0IE5BiLdYMyObRrEUGA1XIEYVbTmupTOrp3vvQKjndXD9qcR3I0Y/
js7Tapw/oVZF7K8hxZlj63KIByWjBwwgTJUxGYfI/l0xXm4dI7lYU0N/wQYxjq7K
0/bx84iEuClB79DeO4P5aJRy5QUAbVqxPt9UYJf/1WTeaoZ4mZIywcBr7KcQ27UR
iUsqPsvI1jb+H6sHKZjqoMg2UW4YxpgBKL20LT7xJXXjBEQ1UbtIpPXtIHY9m4ot
fkpIc9hA7gctVQffD/fWaS6Br5aHeYiorsd4/17jpMoLLnZ2Jek1Ni4yCxAqRgGe
xztJxwNoxcJFTfXdOhdxA2pf8ys0PYcyiVumeh35kSg6ICL6Z9VnEe8EtNdAcMwr
SKredjbk/w08bER/zbo+NeUZwcpCBRk6FyjFsE713LMzN1Hsao74awHbyKmmZowr
TWCCpPANKlcOYYBL00cPndwDSpH6H/c0xPO3HcIrJWtPXaZmO1L0O85beJglqYAQ
ZBWlzXiMwG3cwAKDag5RVnDn/kT3muMqdkKR9AfH5pSxFSsY3xP1j1+EpHnW7WVE
qwNbfFF8ylNVQU1ShIYxt7dBA9cQ50aPX6cXlaAd1Mz3hoIpqnkt1kVoF2CG7bTo
nPPbpCZyp337C5zCuyc+FsucY0YF5k8QimPOPt4SNDUItGxaFA87E4llFbK6d2Cm
Vp3zyPFv6aUWfV3AbVqhz7g3nSry9G366GWPBpFGupdXco2ZHN/x2zj6x03MB9KG
9Xa1LGa4clZ4dv30qhis73SumvXknCEF2tewirvCcWeGVWbBH82nJA5nAFbWYOMq
3YMAFaj4M6G5nePei1GYvlqhWNw5pH+8EBGaR0zTm+qWf8gpZ2ioqhqQI28e2JOt
s8UXGRQwOncwX/Oy+lwTLtBoKUDcJ0sVRx399nRn/GM/t2Wd9ae3oq0q5lmrAUIj
KNZxM/uVG/Pn55EmpJ5OJnfIyYeuUhvH2TPdfP9+bhE2iXml+Sthk1JIf0Q7XVj6
KaOiMn/HCXEJbMQ/RTnAD8yv9yqzglBDnFAg9MEr5S7DsvWRvrhijCxjMrdBOCZ4
H40T2p1yGnRV22SZrYfSjhSu47QQB5cSae2LJN5pkIC4YgVyY7OWFo8pdsKfhLcw
Eaoor0BbFb9LjFTTa9EkGE8hJSxP/10OLzElj3yRSgYJff6G6xKsvQ14Ras8ia/2
0HaOi9W2aA3lC2QCEUd4Oo0t4SYzwqAdZRFdVT7ua4Yg1kK4RnNhF0ekAlgrr5OP
97Ve4gKWvD1x7EuhPlKFW/X1SNJufI58AqFEMDAvOmWNXvuJtWSSeLdbUSqDqPkw
b28cSq32NOoOfUCM40PCQe30Nv6ZpSPSqi3cRrEQOnIpwP+WuLHOyu9tFk1sRJ+l
fbvCUBumWiHcHDqnj6LXM+IvjOW0698huMbvTDbv4FPn68STFRD1V/dITfLzUKJp
DXtlQ9SPB6gtBQyv+b4ANxDQcSpF4ffqld1mXWNDORSE+5KE4B2eXBDERiB2rRnB
bmHnxKI98Epi0CRbnvjiMEurFZSI65B4Az4cWDrR368QEWtaGKQ5nR5cKMjqiRw5
s40OYnd1LN6ExIIAk4Sp/KBPf6wWfu/b/gCWjLjDTj5KI5yGBGIuvcTQ5hAqM8ma
VoWRA0G6s2lXVFpG7kwVYF3OscQvwnj3pgyFgXb2WZuhXgLNNe3wOsD6JVrgxI3g
x2gnZEee86HJlhfzFIernGbM2EO6Dx2eYY5w8qYbth+0El2e5bIwEAOs8TqxIBYn
wECXEtiLOUGoSUzE5qBmPWsSENSWqUKOw+eeM+fq/sKrdX8qLtdN8g++GWOxQRTV
khaqDTgB8vOKr2V7OHQiLAiF7zWQOVINolzT71iF/fiWQULQpyEYxdqY5IYsE33R
W6TB2m2tUWazaC/QDs5GjIucAx8HAy26Yfwfwl2axu6fCnf95li248HAIm924DBJ
u/MLaWaaScOKtOHGLBoXY7nVi4rWif03NtuCr8re7Ky1I1U5Pcu0hcrAAVJFWvWi
lEMfoTrF5KvPQkUwdtMQcTy7+cc3gAb6j8qQy/gcih78M6Ifg4cJIrUK8YlWRxX2
8R63btPOvY/Cdc2aeTbnbxdm9fvWLGcECWOuo0+39MRoFqLOxoqpzV5vrCxTzNRA
sZndhvxQ0+2TLjCSVRH2EmlgQvk6cUog27Tiz9Yxf56NsC7aQvwmy/OH/WnGwbH9
stnvsMtsqt27hqm0iogJ2pmBbxoKl208doV6XhcwpTtNdUcPf/rEllDP2cQZeVCA
NSTvr7iX/P38uaGbDIgGYP7T1witZRMAvhn7MVvmJu+du62IqI1NYJx61peQ04eu
gY06pvbkBTLWTL1a7jVpKuKSDUtbwOmoZiOtD54KhRSG3eeX9Cq1OU9FW+7GpROj
9f/0b1we02ZdjTqIiDhBAheFsM51ifbAtsZyl5hKf7yCEFdAu6cYF8/6lD9atZaz
`protect END_PROTECTED
