`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/+KIrCXPwsw9w4UeNO7dE+bShhupCINLq8EMNH8XpmjbqjjprQiDUSVr+jAJfgEI
5bdYvrpYErIaVizxSKzXKzmqncDsQ9F2GLXPsL3/EP5YxunvwTsbWnhG0D9TBekg
dTscXvYDoetcAjKjVcMDJNNJ/JjeJSNnGhedm+KGaEkWBl+3Dv8vHIYLcTTBH7JH
/rNlqV15gz0Vqt9Lqo7qY4nmSffGcZMolB14NIsClONz3RhETz95kt8cjM9PTB8U
V2QQod/H1f4jHYGd3DW949jC13fc3zZkH6JZk24HK7W+pjol1B8yjVKRJ5FyzYYi
VAoPvgRX5+ag2f8DKdLXOeCwz7jpmS+2EFX+5W5sJdgdk2X6krtZs26o6kgxSBvO
HJ9mW4zzs6U83cLh7vb7aM1cY0N7w7jaB/INEHj3mhParB65Z3LykzzLTnlRzLH3
6DH+xo59/jC4jXR4oeeIL7EDATbXY+AaCdr9BICxpHjXSSQozEV2J62vlktl+vja
yH7J/6ggqTA/u4znWpDdwz5e10Otq6i5hMB461hBz8BvHikOJ/K5AMtbs94K7/1r
fMNY79eo2DNnz0G2FJIVPMiZpvPaF5XHfAFE0+tOFCNgNwnp12YEXIQ125Qx3hjS
3cet7N1l8WtfOq9fYjFZWGlaGMfJuL3SuqRDJ0+bm0wo8mKkPrBejwR4yOoKRNCk
UeC/ZkPnbNGEgHs98HKqjkXq6tbu3SuqANpIoQ0OZdXU7GAm2AyC8xdqFfBT0Kah
we8YW+BrAO8Zdbmhdva70AnLxD2AsZ2DR/XRSmiU03SWBVbr6bYhnIHFc0e7HJ8P
GHcqdMDNcwyV91/82NxFRKrjTkwx1NJ6yZgoYOTcLy41TmnptnsllzeUk/l12YWa
8jTjGo86+jbKPe4nUeHljnwuamVlyvxskpLXZ5C8z1TIzyaZOdtYtJY+nbiXUgWa
8+7Z7gaQNn7GwzanmYqL/YHcTbQ80gsKUiEdR0ZxcmUcdT6g78SItdR77ihJ4/Fo
NKPeJ3YagvTMfaSTOocaBCQU7BNedc9UeEAC0GpajIUyndjOywh5oqC7puC5zqj+
kh5jGqQM9d8/WRKZlxHSTigP3C0PA8HfA8FEGgD0hlA5j/nhVKkD8hrAff3JqkLF
T6OT6fMIndV2V7xV0SiLqmrzPmKG099LCWUHeqCVzI95suyGxQACR+RIimGyCNDF
Ua3PZD7Isl7FXPFT2FlZ1Pe222fv7XJ21g+5eIQubtHygraMI9f8zlId7iU1Ylta
vAB8U9dVcNTG/iEV0BruFTpBTVINc0AHvyOg8SX9a2624XsnqqdwbBiFJTgwfS14
5K+i0186H3/0ylPURUIDozKjcIfrmehW3o88WWMVlE72RACK1u4ydUP1/oJcUS8C
22dpGx0UnUKYZvHd+OJeeAnAW56KksxKu8rMaXtYpqOtVFxtdEmAZfGZXg59+vNA
HPPGyA+/nNRFfFZUu3ssfPVbq+700WkZy5eY3to4p1zUfHXwyFTvWBBB/ZD7yF99
jwSzKU4R3e2sQFp6ZmrhYtVomOHY+CBimEzdU7l7uBYxRcv4MDMyRo3lsQoeTt0f
VujA6+86z8JW37gwtg/MAT8VvSspjOdmMyEfEkANRJunp+F/DEPtXMCCaR+iugg9
7K7QrWa5Zhl+G/BIRc6iLmBRvY4iu6+zE4m+on/zXkYDG5NhqlmjM6QZECzBpc9P
3gBFsnIeE4M0UiQEB4tES3UDEkfTG8Pm5D42aB1QDvawf2OCMAF1I6fOvtRiyF6w
dC/PehAOxdPxKF0yl+8hmHXB4fOqxbs/DsPCqInQoYnFMNSZTs8WneSj1vqJ+d2x
PVL1RZQYP2eJ658Hd+91qjgZ544OyrZBVpCwcBwW5i21OJt/UKbQu69tIu6UzhJF
ismPS41boQbB1qlQN+uLyFINJeUMupJdtDSOG1ThqEt74vhcEEVKO9xGAXzvQuqq
t3jBOs6NdnoBuudg3CKzSYS/kZX3EViPkegS7B+jSfbFQcQAPReF/TI3SRJmOXiw
wtPfiiX7bS1vscJxtXa43ULnMGAy5whI6qaquELe/hv7eKYgRicgvB2NZOwrvDFN
DfYwQGtUCqlAmN48SioiEaltwi8CWJVVXSxdOjMC5QpQFMzNAwhPfI/OcCwDzzkh
UbxPHHrXtqdFoj7cdij/QNoxZAOHpYCN2lywiIBwiWvAkNBoSATgUbvRLsshXq30
Z7BLXkleG9ZqRcyHj+pRwrpkcY3aGrGz8QvhytGZXpoy9t7D99SSohM24DUkns34
/yhQ5pSiaytU33x579h/tz7cl8cnOSIgvnel7g1IUCH+/flXJf74VeL3K8DxMt2e
JBTVS1CnuEHfACs9VARqYj6WintKxQJUd3VJ7ryZ61+L4lIyqvyCUVypOxbfiI1v
QncOM2tDmGdrx1z4xSm3oAEwbi1Q2FMt9pHiN4p2xfFmtRDhhb3hJCzuQUxFMW6q
GhDI4k6VRLgrYww78T4Yom5f0GiD2KyFsvJqJ3vU+4sXZUzAPw7EWuNEUN+DwIaS
ASHswZS8LuL3jFJdnquVcz0GwLSbtFGLT/6TVwpTKcrA2tnnNaKOSXqQZsVPWJx9
dSlniy8/wW6AluaiGCuwyGzs2rdFom0bwPLNKzViiPZ/BTo6lw1LD049MWBG/u5t
y52JedaxqY7UCxin2S8mABjkuAPiBMIPtIbaNl17Qce9+cBIzBFevunhQa3iS5Vj
QyNjx8gvPW/NsYerAwCrdQlejwyfWap6kH2f7cH1H5+yd6qTvq0qdUfPbzBVGTZQ
6aD05e2KhDG6hBYSYoxlVd8j+1XXc/6pUSwIwCKxpfy53ygUcSv65rBYm1vc9IrZ
AeVbuEiB9i+WCj4qO7O/Tb5u5sXzJTfliKOVjFVSb3WCv+RYFDjpL5W1T8CqcdQX
hxT9ONxBx639GmMAjyQEq/Qha+igKEIund0i55cePs8nr2D7fG2/EV/rJ3WiItUw
ZcPNIAbpRhmmV5OwUZFWJOjEVLjjgfzvFbIWg2uKRkcPopOyL8ugeXBitPVXARhJ
i9XOgbnscGIfuBB0H1UyzY3qaQl6z/jABgUXsEikT4MzKIqaoHhCNYtZQlOe+IEb
av7/MYSEwsxIvAFPO55nT2wwaxyWbnHwncgdRwD2EA5/zDSFEckvRGd7WyLPAoVf
QVmoX+ZSOL64FaqRAhVXkE0A8RQsPgEJTjuLph4QKT8xNnxmm+yLiTRgHT/dN/dk
XESir/UrwvIOb+a5E3+rJISyRswu+hzzT0T6McJCB6g4tJJN+vE9oPqyQfz46jET
38OxcRdEXHCKL/457L/b6P3BEpNCpvYSvDdAVKdYjXC7y0Cg5YUgKjRzchAxQVz5
eq0iS8AGP6g7+2F04p26OP6jilkqUYiOSKN4nHI/KX8=
`protect END_PROTECTED
