`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4qAB4TVxRwL68AnEAdM5tpeCtf+tjMuMQkX4jNwzWpZfHHjhkEZ8nptfAhDct/CX
IxdISWgPrCFxHUcKWOthCq0nmzaSlqeem0IMz6z+zZHRvzRFDMW9WEc8lOb6Yb27
3HcK2DO1hWxedC3pZoz9YrxztRTvM0vF4kGSx+VUWybEKNxo2/2WYaT+KFG/boww
fJ29huJGEsTar+8CQEedKB/SoxquXSg1i+2Ew/H3+dh6lHmm1w/dZit9eTbKNtvE
RGR8YjNB87KYA27lwPb3pYqZB/pSEENU9Qc+gvSzjZr+YlY0mw3f/PY4mTHNPIpb
TKi1VmPiEgD2gdQzLB5mq4IdZK8Fa+B34oua8uQMioqpLacylkLUJ+6eGFtVgTZF
FRGn6U6MdASRpJ0kDpDJJ6HBaTMIBOdd78aKBG7Z4aUB67cNbcZ+9yrAgxn//WRw
r+22H23muN67eBJBkyYr2JexKRbWNptTSqSILMcfYWlYpRoLCOa+SlUDZJXblC7A
lylYl6buCO0o4zApOTq7zG3x1ogYSwFFxShniAsxOQ3DuzwkJVgvRLs+FaSL6K3w
eCy1HCMDCZCbbqvR5+gMyd6ELfCR5qsAJQSf5TlyXnpnSCDZnznWEr3BYv5WywRu
Yjtgl4mPSgG6nsk6jEUcEpwGUCug2m4NPTJ+3P7QRloDwEt0O6T6dpmLhjg+MWeZ
Ya4RoHlFaKTPnINyGgFjCSvghiCsBRi0pF5Eokzdi8U=
`protect END_PROTECTED
