`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
840uagVzA36V6IkJY/k/2i12wNzBRlrwTvxbbehmV/URk2AeWtkbNydiKHTEb248
Xk+LAdo+h5KMqWgQMPIYsoLwAPe/kn4InsZn8slNb/RpRXt7Hn/YWtSA4397BGhs
70e27E5ySdcMH0aX+bKpKe0QHPdwysmck/YGMTN85G1hbvv+BK8HQLqedW+hKydz
LbWfqHcLwMHwH3fZbV4uRcUZy4mbAUIwf1L7g98KE0OrnBn6pK9CqzsE23aCG8oA
gEe5gs7jS2WhelZD+W+yUhkgcFdacDEIfAfknL0qDF2zmA/gDdQ7LAoDSn28Z6Ik
5csejbMUBMxb7mFbVCGOdQtvRyQRQNiWvs5NjVh6fzT9cA16T4uMhwCTfFM+Yo79
nUyvWfQhWGXuCfJLSFboTuo08k0nGmwPfo2khXbrsdMmGT67mUgOa6ys03fv7bUs
DhdDfrcWhdpBb2/UYwlddGYHT0pumXbvI/MKoO4TgQ8jrF2xrw77HkO2yFPG2UJ/
1G4Q63t8o2LrR2EOkLDEiipsj7GcvaTqsmyMksPT+JyoBc5L+2h+j3RHwGSVt4Ja
a4S7SanaFZfIQRPiBpz87yXVAlQwKqXKTVifixRUCh+lN1Z8oZXIrNXy/vRMJgnC
nkhVSKJAEa0pJFia7XdUYL02ojewbCkWzDQepHYHbt+yFMiNcg0fVhojXie9nf2c
xZVd8ZKCpVvwkAJ4SAYJgnQwHMYtvGPtEJGVPLCjg0Pl8RSu+BzDKFPMk7HavXo+
Ryzo69DH9do3iK/0rPxdMUJxuzAhRuVYSUXBC8tyOmmgLcIK3SaLoKruyBniiRR7
ytHJC5bDsX4PE/oTLO257/VTON+6RXvIvfGmEe1xhA8wjUIL4QzGdCqL3FgwHjP5
zOZb3Z7cwkbwjlal25MkxKhXmzIf0CEgS0PaDoinG9snx9VJylc7TzfecnJjdfLU
Nm1S4Y5gePoaKZze0UZXT8ckGaUJEXXJNRQN0j2PLKmw3OGU2+nEq4XdCnSU8+MR
q4dEAuup4GGIKOaI8GVCMOvNT//0t2pk7m/LKXTkHz5/y78kVEijDYhQCJFQmsmS
mmf1m5Lp6gvkiYmf3tlxwpLTE1S1RTFkBclKuL2qd0k8hCHer9LalQceXtcp9ZRi
CZziaUlz35rgOUYzCu8jJrBOu6WftuIDK8kMG0vNHwGTZSw8ArmdiM/jFTQFj8Hd
z1X3TpiusYAYAQ/uLVm3seZqNcFVbyFhUK1hbdOCn04oOTicY0SmzHd/jNuI/YIx
gJUSJTsVty9VvqZdckfRmkHHqgnKsB7n8ilZYB0hbw/GY6ZcJgTQHpRL0CnNi9sw
E2BCLabu8x/e2JY1maP+iMnh3wxKX+t/5Jj32wnsy4CPA0YIrGrHoBE+QEHGZGe9
IgeKCJYIrDONd0phs3tQJagDcYzTOdtAjkDwO6leq1M5BodqoNWJbbJTfR/qeFVP
YXm43rw541MlNfuJ/74WpZjcgk92L1kktucU54ATuj3i7gIgBlEu2ESLezip9J5e
UTqP1eqQ3jcdJQYuXuOpH9mGk3K4sr8U4lawiIM6g2jmfm1F/SszExDuzDzrv6gH
NXNBvad/Ebl60WS+eT9EQMq/waoU0WcLxIPQtjFOdfgQRIeE3sYJ+EmaiGOLWXdP
UZbfc1Y+0MIpA5TDME19Mm041uQpD2OqhhKFCszutL+ViaBJ9D2I0/bSgBhsqYhj
/o+uOQDFhj7CK6NlHJoVOd7Cfr0RBFtnbigDqCX0apY=
`protect END_PROTECTED
