`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iywGc0e6Lui3TnI+uCZe9pEDp+8cl6cD+H9suVWNsdwTJJQjC+V06wUBwqNu9vMS
1ED6TTFQ80o8ZsuzeH+tKZignSX+b6w0Qi7fn5ODDy7mA4LNye/H5ylhZMsAu/Mc
/NMlRNAmHc4zPwU8FVqRST3lDjVNs8Y9B0fEPlOEjycM92NvRqQwTWarSO99psYE
mSsX0LBgALCX4cGzq4/RbdAsEgANLK5Zp8zMTcbIhNA4wJ5ZIb4ErQfix0mMNXv/
0pNpXM8ehi12zDC2oosa7Z1N4e4IxGDe42bXBEyiGInECpIcpydsElxnsOx52eAZ
DEeymzR/VlbkoBt054GagSK55mTuiOhEV3lIFSC2Q5PPaYp2LLWZKZgmD07NntYG
NXLYTniebPu34Yb8QBDWagcoxLQUQB7a/6z8NiRyeGxIUJFKSzFd8FKM6ex7Jh6C
IaEhPoVpay9d+bG+FAHGVYvcjHLuHUiNsrVhhAJCYbJpwO32RdEKRmyOZWGpEkj8
g3SKNNWkPpVlyyYcYrLyXgX9vEMMqu14nuSG7+BwU1y8fP0Ux+ajufvJEmkNDWeB
VlOBv5k8Ol5R2BhTLpR/SFiHWrbNaQP+JPVUVE6WiRPM1FlABjdxTS+e9Eb68vO5
L7w0GukQz4ES4wmUUjrOWKXRCuIJpT/aZqwpHtxo9hjXNl74AnPJWgjZ6vstHobT
NCGzbxddjEuFQijVUPlpIZnJGxhy5OmwT0AnX8Fq+7B0REtGV9c9ttAPOhZiqR81
QUxO8FaEIijCq3xYsLihHScp9chPAU/IS9VnwaY4T2Xy7jxmSPV6EGTj+B251xt4
vZEE9jS/Ch99QK0cC4KSEZxP6X9KmTfYt8VWiqMdNhTk+6TE8cdETIgW09DI6ckc
uxqRdg50FuAB9xwPF5pCSQFLntxlCmb2IpKgmsFyhzcfe+DawgjkCNkmYFNSaVHX
apiyI7zvAk5xqG1jtmfbxRmpw8T1HSkfC6+6VMwjkZZ9y6XDb5r/geu3erJfn6IV
pUCSAJf3Gp+nSj853cYuREvTkZ8V4FEF6iG5gaAXUNAStiSFZZCx2jA7m/cpA+xZ
0SRwm2vZZAUqqdkFpoL1b6FX7cuo4LJKVTEJPY8kuyMP0YgrkH05iRVsIAmiV1Wh
MDaLPnU/vJ6k/G/IlGQHOWUwH9dm9B1p42RqCYvA+N9+rZJX6vZfDIro5AWvDKQM
15zQxUr2makbCOfIdv/4ngRPycCJdagZmdtlgXzassYXUn2jyTjem/IjBFCXCmkw
Cn1/glB9qEkw5TM7gnc7bd/yqxbcYcA08+voot7yWpECwruW6JIjyoMlTmKClbun
6xC3L5C8TMFp3of2aSMbOgZmZw69uDPBJVRQxCl9XzY=
`protect END_PROTECTED
