`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nEFA1kutueKWZBTt8P8LtQIyTuBh4r0cuja7VOzbz9CP8a7X+EtvfcaEDTELwAh8
hsa28Oupk04vMv9C1Q61C/vME5Brq9vuyCI5PrmHz99tpsMRsQPHo30mNAY5jecA
oO7VyKXYBBgKjAyoQX9HctzrYBXV9CRJ4gKK6RbcCDC0Rp95t5zvRp4Zha86t8X/
ZyrVNcll+Cb1uJugCurAanc+9I8Gl4X6FrgpVk+81Ltw4gIim/3h54rHN7yCFgF6
QV6rbhjXVy3xYuredZCQLdYcQtrp1U7QrTn9JDMYWcv3G3rCCTfBRXDaGhkYHkK4
gCn7h7EGd7c4xhJE2OVbwWXJsx4UE81KTIj+Yw9seeIHixw8az9g+LI4KnEN2TsF
SeP/0XYPTEgF9EC2x0xzggMA5n/PQJ10XTCvUnS7nGBnp0nSWXr882qLNv3miA/P
a3BWy+aMAs4fvuoLS81UH7S5K5AKDoC5B4o+6qC3wyLO5bbg56hnmsobAysE9F66
bx+BvpX5fNtuF9EEEhx/eA==
`protect END_PROTECTED
