`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H6c9zdkODi+b2L+wHGIRrmLuvGSf/jal52TsEp8KPOLbJ4z+w2ACcBmE3/AY6ghQ
L5S4tkppAFitvs315XdH4Zb0uoFuC1uNOPXkqI//q+822JROQGsGU5IoCn182Slm
j8GxBfOQIKctxCHCT3XeWJ96xLP6zRnCBsibGt6xCEO6YcXVOZC3pABZvKxjHc0W
X1yLoW6282RF/USUvM+wKhX1mMjwuyBAq5IfwkPQWNz1QNMC6/WFjuO/IOYiMMlT
zHvhcG/Xvm4gxNuWYTDYO179zuLDyZWtns2leghs2++s6Mv2IDHp0fMZWVP1RNLj
HfuYpBnCzVYwRxte1ZmRTOhwt8OD6CN6xAjAQhvIpvun1lOYuIyj6/rhoBs+ZaOt
gzA2pbL0rxu5txCKvkBnc+SBJuQE542DLmmgoJQkGmRYrxgT64/OW0CMkRLchS19
2C7KKDtgNbwsYnPRkqnwbYRYDMMqxm+yhlfoCvwV0NgeCsGGweTYm5vTZ2ma1c7+
NTQBH1hojNoLgfnMQShq4H2AimqG0W1wtBF654xh5kgiBlOfbmUB48UgPQwbcUHu
0N0cOb1A+xCudG1iSPrcyXG+bV5oLuDHP8GwOFjgq96y74AG2aw1u1D7G1H5jait
WtXZ8AIZR/fdzVlin9XFvaYWqiKU/KM6JjaR0cxUdp6RKqFCKN8XV0UPcS+KeNyC
Mtazk1l94POVmAAl6Gb8sekgtQMKUxibM7kC951HblYQvs8kpQZPy5yn/lO0h1+c
GeJUULf1oeriFc5UmPDc9ASKQKVBCKGAMeH4aW7SAqwpekpPWYuzBmg0BojJMw5H
bocE7386myblzZV4AZJzLqk9n3yFQ+BK/fZIMrJt4ljqNHZ7swgeXquBoK+77YqK
L1taK5pp4Q779fij7VjzfnITAio+VkfE6VmV9qOUondmWQaOKE+jHs5M8amHiACh
ajxbX06QkczVes5KVuwPlZKnSZ0IWnq18NgnzI/lbyum09IAcH/sOxbxyxDP/WtX
iMPqzAWRK7C11p4/Pp1cwMLRph8FcCA+NCLO5afqqv7R0s4Ze3NB3BiIB+mZko+D
+pddpgoYIVhIumW/35Yh6DuzQ3Vj5MWWhruVJtWC3ezs7s9fuSvZ5xberwA1AaAO
xCxudJWeGnwOzVBe+j22Phf2X4QvoV2p3EBV84EjOJk4qnf6lnqyAWn6soBdStzn
7Ky9OCKeWhUxDZwzNbBJdDtgINddpVzBsZXJ5RgNbem9HDgBwlKUaFjqIyx8ZPOq
b0yjeqnXROgih9ksWQFqzSyzpZQwHfYkpHYssaknf7R4YYIaUJtoQ02v979kSGe7
3R82IMJF2er0lAyHvmhnzEIiKp8feeq20ulef7Pq8XLn2v5rHBZyN5YENRhELrfD
zKw+O7OAg8gCJlcdnW2fHd9SmfcqZLQxTqoimkNh8ElzbW9Z/wygcIeZX+7MWXKr
znEK6UJIUloOr3ViWPDbqP5KOp101A3SEnij39h8/tFWftEbwxXW1T4MYDrFgIxR
40NSm6QI0WvtuA4q+Y8JKuka2qcJWr7liGDsDJ7QdQEWW4GeV+T3X4j1T3+2c28q
LwT2gWNJ9lytBYnN+hs49dgYKZKmInerZ//5kUmntAHfWRlRG5nmIneJJffxgmGg
6abUtP3cDX4MAU79mMnFi+wWpGSGN/cE9aiLGEtyVl9y4M4V0xL1f5kzz5vIKTg5
DztaZxIggp8vIKYvD3MdFnfBh4agj+Ma3PadUkwIyFfngPRp68QmBPOz5AaY897B
5h+PGv4RbhoFQEYws9f8Ep7IKeVUt4zPtg+xJ/UzdnNhw2mZq3AWpbYQyLODO1jp
faaZxbnGZqTBl7WL+BNCAAbf5oW8H3K3aFHSFiglJCRMVaOmNLfk6MUeR3f/jajA
KCRkUEcvYpzbWdHfB/AhByEex98q30YExrh7NrnqwgyGckrzf5/1LfjekJyqInmU
+c76h0SZ6RSOz7B0VMyDDk/Ps2ZsJoO5pbB6gsj8jEYgOTFTB5EN3i7gttNCY64/
J0Z6FTdgqDImOm2j629vfDQGX/0ZA56CFVmfUaoTYCLQu6aJL7V7vaGeE8N7yb1F
FccS9Opyx3q600m4oqD0+Gig6siKvdM4DQy3is/KvEWy2zsIdxaBWt4OVI5+13ZK
D8ljrrTJreLgAniO2d+is1t01tIZE6x6qHa/XN8CXqtVf/spBTVXbY6VGoFMoJiS
IlqiwkuBBcXi3ggotUoDphWiT/ND0I5v5XcecuDFnE9fYWRAt3Y6vPVaJp/5LIRA
8WJmp503yZBEyvRd7amXL+7cWFS/kPojeSHbvoOTLPf7j2eGjefb0SFloAW59oXL
sutoBaF184qDPZaQdPEjLpFA2xkaZKNmaOBhPTztm1tkT1A7DWbVZ+lTDvLJP6j3
pRnFs3ESSojkH/IA5yYOk4xb8HVai5H8YfXW/BNahO63C8srcHm7Cdgw9V6U4ECU
fAGWzrbxzXw8VKwp7NJRFZyHTJcTh7Gs1VKMxyOh+gqOh0GWqtJqK+CZB0ONS43G
/NfEe4abxnpNL7l4Zl0zhmQZ5dDyGF4fp/BZsC8Axj2osWLSK2RiFR5aqyZU8Y1l
uWzxSE6do9uELZI8nA6GlUQGp85XAarDUEd1mS45aLKrhx3JK9UuMhneK7Y5qSSC
F9xVKXxcS8Z1ZsS23u00swRpNw9Mb9zUodLL979ZVxDpUxMUs/+siHHMzPsMxigU
ehUTNuNhcRySQus+fw5yQwMEP1L/qkwPPzComf/u6Bt/G2ixkAA3EqdySJX447rq
bCMXyG6+Cc6iF/NHmEJRG6ItXLQsSX1IjuBhxj8kdQvhJCaYVzH6ggAUiCrtCX2n
9B0S7BEvFJF4s0zZaJ984sxIWquO0iV1MlsL8xg9aJi3ZUkALq6CKGmmBI47sb2b
+AIZiR5ZRyK598dbvM0/GRSpT8IgKNsS6X6KIoeSaxlz0l6lx0UHiZCDNbPuh5vP
5tj3k3PlGr+421dbqL79E1MLHck0iywzU+Bz2e0Cz33aVFSwC7J1BRtIWp7T2IC7
GHL8BDir5u70/SLttVffZs7ssc9uHjL8NMPDNzAoS99ZssYcof4WvjjLpyfZ4oeD
CuHqxKVMatPJM0v6T0V3ml9GXIHc/OW4n+9T7ObbwB+K4JuPn02fJKoMh33BQBwv
SXY5MfY6Z14C3YeKXcj7XkS3XcKmurMpOxVPq9rOOVwq4sRenmUeWUyjXeHknmH2
Mg4/muM9p/ihH5BWJ0EDfRMy/OiNnInsfN3+UQ0A1Nkf11thDf4LeUDvXdJnYKuI
`protect END_PROTECTED
