`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FZPUmzWLlf5CB6NW87kowfY2qsbiqf1t1Fe8rYnJVsA/cAB+t3WCpseSSFiB9xtK
z+nikXIcD20h/MCN0hLjR548Go6SPJOxyot5UD2P4+0/pynNvt1cP0XnRortviAM
azdTtWHfuYGwoJ6AIMPGFc8yZOlZYjl9l5ENHhYV9CC1HEsdzVoSdxP2xsGYRvrO
qr6gNiODpTB1Bcp1t0fLQ0iqVFT91DQeq0fu/Y3FFMrWl9ZkN2YS/nxgnUqalFj+
jqCRve789G1GhF/7yWtvcmpZ1mlbP/jfy6iNUUTe+uJEmUxRN4mAzfdCE/SeFm5I
zE5IOi3inCBLqcakbM7TQyIoVZQT12Mjmku0IaM4RoCjnyQIFjS0KOzt/IjDx45X
OXT/InDInLDWF3kzRJ2ukcLk5lABgwpGe26ULgEoszJCz7w8JMS8mqc8QGSBakln
zmxw7DsFBlksnS659P/HBpBfTJXpsIv7BHa5YVAE8//E9D84dnmItTtG/EGOsc3y
zEPv2fH6tNDcLBOhFj7cDkjBtSnJggsyO6dj+DLXmAI/PTIlcXtN4rCkS8P3ahWr
wd30kR3gCzlW6PBgeHJGsVDPNDssC/tuJp8BobnTI2FaNk1RCQoAbJK75k/1muO1
Vbz9NqEWgYvjKPZGNiRxh6bcfbGUM1kYaedMnBorsKQ=
`protect END_PROTECTED
