`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lciwNXLw+0ReylP/qswSFBsOTc3W6qc1jS24m+WqwFJYO2yFIP7bblp6fupPJWgr
eeYvDbEolO3n0lWP+qtSoQQggHimgnyY2qUzYCic9fxbgQxliOyWsdPPUmmZXTAx
NphCALg4mTUiBU3AdmnXLbmIEFDdfSqtUb2hK/Ijz+szemS2jKCwBe/+2TTIWtqe
TSophM5/DSgc05IkocPw4Lr5K+CBpl8Kz3bBmCA8/PLJ3Ik7EYhroqDzoTOT5A2m
CJgj8dDqHf+MmQ4MsS3z/0FpZED36JadZsYXCwnE4rjNKUzNqKtP158EUthtR3Rz
XMvkt4SNvcalnuwTet7Tr1QkZj5mv74QSnVvLcDnlDt1TfIqvQrPSTe+DKV2mDyc
FqYcUJn8A6d+JREJOEYJhHtAnVI/5PY7zpnZ31ImrZk1jtr543v87UhxK9Jtd+x3
A7M4Yfwj0XhfOVkeIomNIQHb2hc37K6GUSv5ROrCWRoA++uAtK2Vu6u4/32Ev1lg
xQNu1D9ZbRRc5RNrX9N2oTo5vnfboqmZP+HgyrEzLdBkMnPuzpCrw2xbkQEM0UGf
TLWX0+3peWEaSe2j8JITvTqM2pJ8b4qu8Zz7ESzbTA7GOPxw1iBHtkkZ8+KY2h1s
bB8WfafvM867MXaKeuIjf0X4SM3vvMBCYq+g6pcxmEXUJJnNA4EeYeFJmBC4YLUe
UJEHHiM5IX83huI+9bmjnZEiWmGcgSi6ppZ8sG2vxN/VQuR2Vw96f7SUV2bvU4Dt
MeOwa8Nxsu3C7xeAFtYeVADcy+Da3HfuH6XfDQ/G6w7gd9ahd3ou5ub2e91l9UWP
2tAHmLBvk1n2dogdhQc1rCKxIUzEEMHsGewX/QzaFzJkDo2N03QvA9zn9Z5WGPqp
Krzj9p6doZ2707RiRY2ieYUBioJqL9dn+CLyAeDvRy9gWRs/NQRrLwDrHFFr3I1P
FLSUTXDj/QcDaRWkE5TMFQVS0ijLOL0A/09IgmhrZ2eSwUeRGLNdJPi00+ptzey7
0Mc0CVfREESVmhOUWPwfUcYnAcM8loP4RPWebFPtIrFfmVfcykvFkksh2b10A0WY
wm6xJwXjnAZqDMioJ2ghoGqZRS0bGixiSP8hZ7dHVufT3Qm/kKQootsOLCeL4khV
4qaGwCOtC7s8mfaiWfI+3gVnRAevprukD+7vKo/n+2Y7iFXuw3poY2hYani3YoLU
Hzwby/yCVK9Os/k1kGINsZ4iQkghzYduqyMGjgDsUg04KD6z2DfhriUKJPUgG3pF
kpGcdEzjg29Izk/A3KgdgL937/NTG1sXdHJIrwZSQI9bn1TT1IaokNYQNsjL3J0+
S9bUNg5yJKXFlHgt+h8kgfjdQZFe81DBw0z5fay5mXnSwPm8JQcMM8WBa47lVffN
KHRkEYE8elTObzOnjvTW9JlyKbMCAx77bQcCeFGoYov6whw/EKGZTfX/KxseeHa8
hdfXLyK40vHae/SRPNgMJGshfMkehFGgKkEGfk31eohbNK28t/0RaG15AegTXGi9
8/wiAZJXSloMRRMJ0TnyJgnntlTG51YG7st89qQojIDFX1rmcGRTz3p6XuXy8C+2
oaYfmExFs4XWXfJ1b1c6nnOPTqIwo2mmzp69fhSCdWI0P8sbdVSIvjW01hb2/yya
ebEYeloLzuZigE9f7rb7GbIZUp3/HpEmtR6hq9tcZYouGcO6NDtOsW0iRqAWM2B9
uuuim4ZbKKG5TSOprNWDrRAs4oNDjoeTlDWI6IibgUoTr9sqWWc4dSJt2Si/iqtu
WwAt618cqoqaXvEzmYUVsgJ3f11azfc68dN14zspAWi8fPx0eR8O1g1oTwkpCXBY
t5LA5+yw3KLSlAz+TrHBpKTiXPbpRu+BqBQ5Z7Fi5nM1hjqrj8Apict7LwOhUsfH
iOi2U7J10EtY+bjTg2RHbTGGOHm/sxsX10TrUh7el6K0J8KtImLaNlkzKJnMRWzU
Hj0EayLmYxKguSohm/ebqUd8cGf91ZE2LT26iLDE2VNYWu2xBLHHJlQV75sdzeHw
uOHW3Ork8gAPEnYq86tD5a3/Wz4ajwNhZ86Ii78LhA3F1DC3cpHEAs+r8/2lwRBT
0H6b1iEULDynQMdPZfRyuLecqDfpbl/pfdrqgbNCxePmzOK9bcFWXnLFHkiDhQ/X
4wAvph+87WKhtPJmiTR9m3YJHeXEE3qwx/d8dYXATgZdQruGb1Uo24S4U8etBdAW
onmavKQZyNtU78YtKMZMDgydBLLKBOrlHTyvNcDJr8IPszYJUYepHC5m6cQm7Hul
ew0K+uRsAGoZQygmKXaXeoi7hq6yrcdC9q2QT+mgYJlLDwB7pyY3wAckeqfVEroO
xYqTXepAxSSr26QmgH00Fo2WaYs0+WDNYLpxjaRdWk1960aTTbYlOtn8j9UHpgSW
vb++/7MOR6nC5AQXhaqyLyI5J9G8xQr8VLe25V5grtPX+O4nInItcbGu/nIuqgtv
HTk1ZXP1asi8aMrOpao108Wdsc1gXq6pj3Nf0pDGRLAyvpxWPDIOCqKqwRp4+JgM
5minqFH6oXjZEBeoUPQH1LeMtN3gKwCznjj84j4WEkM3Jt8HPOZBvcOYzf4G0S+G
xp7Q+ugwn3WhxZDzPwrJ5+rAlCopQBYwrkTkHhsPzi4iSSCqafBp1lE3Qi/cP4TW
dTH+wosUw8PWi9khsrnDX4Roz/HnbCQ7AdrCbsLqJVCXXB/gZBybJANG/unGcnSq
NXwiM/fO6UbRiExdbMyrPLd53N/EEQYT9fPEz+SBRJenloP3gYh4ph79WtagdagW
acE30Myw6/LUrC971Q8hO3deqfFNy4ajQ6WS3Pak+20ke2r1JnskHnhQdS2iWthL
9xi1KEMXLInyYTkVXaurCBLvgWRaAiUgqTTgAeI0X4GvlsaN18dbb+jIzvCPozFp
bO148twRN+NucTab4s8nPcElaVPzpWfEym+uNiFvKc/oxMHo34seghYDohkb09Fi
CnMMFfK3JKAivu6GA5d/yGwzwZv73MUFgTgBjp2hm269HQHQ1Plqat2Ax/JryjYQ
vAOoZ38Qzb6aftB2MXdTrVTWhSW6wmOFy40Jz6SA2jANuSkmp2pSCPBStfBjPrXc
yaa7wKo4ghf5PNVFHWkjDF6Gf0xpXYHQ4NHresbkozun7V29+fIxysly8rCIHHm+
uqhJnt/K7Il9Aob3rVejOZMOhwez7QfoH1sIYTzSDiiMoxFekO0F2kRhaiidNR/i
40Hp4Q80LZcceMNkxl7TSuWYwDfkFkuC9e9qOXtnIdGdIBga1SRrD2uyyBYeaG56
/Pu8tyaLlkEHiVi5iDloQOM5tb3aYNOlEcfqoly0S92baTo1jV8F6YY5CZy509nM
DxWpcSH7f4egrvft0T76K7r6B7Cr6FuWtnuk5cB84eQ0u8PQM4l1QmxQBGQHKTIT
ZFdWK3dKkQy5uBDlxKENRGAt3OmABQdd/8PjBGR3iShKiv+fiwMkW3y2rcR5QDp+
3dSQwB8VfkDyzz1zPTNMRBU1O9401zvxBUuRvYZo7dMCratspMpiYSiJzlq/24a5
PekPpi7gyL63CQi/XMTei+9KNW2/a7MxnNnrtoTgwRu/CeoDe5P1lXW/6B1l+iXW
d2FPtPby6k2LCsGQ99Kx6ppC5AXeCLfW9xsc0jSxv6pdbqhrozeoSXjCjqFY4k+B
RQpyCRDBpo2wR4gIWeN5/iXtKhofkr+Uoqf5qytj3QXAL4XoZF78iYSlCoAkP8pP
6vPSBXAmvDytSubXZdEBnz1WEs+SGwpADUbQCChgH7X/ivTnjkKrLmbGqMf/C6ud
DtM1xq5S6k/fA2S39ME9OvuzpJnZkZ+4LykSI5aNMEF25cD4fHQIwbMOKibcHQuZ
CutqlAQvr7y86k+l81NR+D7wd+a3MViil0hoMmy4SnHz9Zai6fKYyAj2tTvwctQW
7l7byexKqm6QYtSOKN+xSvOeXSM0UmuJT07bAEZgmsLd/SCQ2kfpxp54NnklXY7P
KQg9ErAWgd0RQQNYDzTwmgR4TIJt+qsHU1iz4sydHa2uL09WpcCVb7RZSFUf6MFn
Bv8Y0t90WXoIcGqnqumbvjv0j3DPgUOP3xhv4CepjyvEmY1pIzaooTZpm7X/gidQ
AiFXIyIF7fqXv5059vR3eC8gh29ogWBmNGUAeaFOK0imoAWAgkRK6ylkPqUKK76P
gShtC3v2WcYHwR1RA/r820jrTR17UdHul8BcIHHfIOiBDQp+lPl7oTf3rjZu6yEx
l7FL2gaskTRGZ0vcJI7zzpb+fBv878v7/Q8CGOsUStzH4wbzzADXWIyrBvsdfOWF
WXxH687NFYbj80VnsaeMkq6Biidrw9q9YIBmz1OhAmnnXbCNflXHyGE9pyJZKVx7
67Lj+TRA4e0cdjRighDPvlVe9ol501SH7Pxhk1cbVlHE6iJpfSIUOYHo8gobY6u2
4Gr8XVjf6uF6MV83Vgjz18A+8HFzbXxnZ5fZpA7D/IePPPwMjb1Lnc9JYnYdleqP
RKIabn4AptIujlou4EYSM9Ij4EN5jc9/E4s1TY7clAAhYEt4okPi6fztj19V1SNz
JTsEkrQRn2/b7kHkXsnqaOFHi+tO9L38bDzseSTcw/dqgsufLSMo5c7dgV8NZqmr
j4Dfgq/K+voqhDurilutJQid4ew2TlsvP5GdemSAKPo3UeHHX+hNfW99wBVvLQgj
+MwhpeDbomcQx8+NX5miYoj75CZjQg2S5gFj9iR/y/CNu5IXSvNJqGE5evM2Xgna
9YnJWLcZi7zIAb28sHDDrpdH6AJrod3UP3IoRPpcAFNFqfECRL9+5GePWEp5mC9P
vJ5qhHIDbcfHHX7XyYMx06oijvnqIGW4KLtXQL87VghjUVm5ETl8cNJC6qe6ryz3
F8mobnxUpEGBXY+X3T2lP8TaJ4vE0URizuKPJFLexfwhSZx7/ptN83izCmz5Gm59
BIMPFGmWHsY7GVwiLtf2ZRVECCdfYkulrinA/5QcNw8H1Z04d96ZJ38OvU0JzVE5
AUaJ1GFCR66BbGn4P9d1QJnorNuU7ybTSizVk6WLtihv+mDDY4haenwsvKqWl+hW
dXyCVzOBTBtVUm6CPJRvc0Ntia4d1EEsGD6x2uD/1QPQoSCRyWnucXOm9WdBgvs5
9VF6LD75JomsyUNLsPoPhrkbomfMxs3TLt3KSijtM2lPvXg9VfXwiCv4Qh+lHMp2
VvL+Es5pY/o9uXqQLL/3xCQ3ohb28ZrCN3YzXcvpYMawnNXGt2Eyk3hiJufC7mU/
86iw8S7bW4M92hr8Pscx6/ZVZ6AgvGM5WMvMPUbvUPe0C7Np+V1bLspnip8AAf/h
7vPhRfXZFGuHc/2Y0Q3Vos0fOE7y7z4GkUQ9P0tAL06aRxSEe/drAXN9RPRroOsm
x/DrAfiWShrRQOSeaNI4ya5LjqO+XVkZfeCCIdEs1yAqO3WMJQI/zrc60P2PJa+k
9cjsVJeEAtFQO1HlLtnptf+ABQE/dpZjiISZGTtOYuQhw+SkN/S/lZ7I3VwyWXaq
wt1nHIwDJYI0VbtHpG8dUTWmn1FL5ScEO+Noamb/Je3Ksv0z17Zaqf2oV1DaGkKR
Zq+F3BQeqoNFh82GP52dQPcaiTZQ46Fj+bVavPHBrzBAFvaZc6mSFkO/kAqDsJRe
B4NhACm2Y1Y1kf+9A+2rnBt9p4BsriwXRuhSfmrxzylrMq+vG7WpD2wpV1PU6kxT
am6r134Ew+sV55Jn4B7QIgZ0KyG1oNRu6+r8/Q/PfKuYrjh3BR2V9lFNzYSoMZ+S
OqYekwOWqpk46T4UhG7VMsUODfWqq3+jJwhskt0ohdPLClFw7QMkbQqW5JMKpsaR
PmsTVOgdNUBgWoIiYx+kJYzxCUxYslDgjosJZm2IhuNSxbSGLVXJFIpXMh0ppPEa
MXS6IaTIyD5O/4QNmTwxljMzsK03JLvsxXtCD7vxhalmLbgjxzBNmKoCtNln/nXh
6LK641PiTarW8P7I3jlTcggTg+vIGi6LRMZOFNefLtQ2j1d5TYxRQyR+aXVNWei/
4n7lFTPHcH5y9vSOsxU44oDJUM0NfIENF+nk7FiernsgdCTzlfnbrFn3eNAaYuFD
zAtuubDNW0mj1GyuQ5acY+E9IR9CD8xXZ+5BgLTzPh5Of7z8mRSFa0zR12IY9ngx
tgL20KmGzb65bv4KQdsnSDJeJQTnS7cKBHuHKSPRWPBg7lG0njBZTLA8Niz0DW4D
SC9rGimldGtVdAeGM9LyqthPNMGiz2ljM4HILR9iwsnN+sReRnCleR7ocw9Ekty/
Xfbt6Nzz93rTtQ04qPQK9oZtSRynNWC5BGjcRoVFYvk2MTGCNuosJVv2Q6sCCvqj
KBZTL6/rLgLuB6IEX7yncdyUvQsuLO/GiBfOH1v25egpuGx4Fmdn/Sk/jBa+bCot
hExuDuzMJn+64/701Dj1+nxd46qXIIdnsOzZjrSZKoei1CLySO18uSXaRBltD4Qw
IO+9gCkCRDormgAWUfNm5FQrvGZslAmyqDqV7J1n+wnNiS3Bbe1SS90uDr8+/f24
Wnjo3MoHVIyORUa4oliZZIiFqxkZYVqllbdUGkkTVKn+AQjSlODFIkURAtZBw7l2
SwoA5yXOzDGZ0Vo/T/ZYMmWz6l0c08tMHMf9ZV7hHPUbGX5dkQEa+ymCMGmHo8S2
Q6VWqhCVGhOiuNVQmD0/r+sjGChjBhwpPB6mRJ7akfJndisHUNpkINjS2M85rXpM
+fPYrRf+WmVLIQ2HUKJqYs3uKhUSVQKaFI40rmf94WPOG/HBRqMdsxGGt02bcazZ
AKgLQqMGwJAnGhYhjnatyY/hFWomdCJl3ByOwsgII/P4CeCJp9gt7mqbDAV1tHjZ
0EDRa8Y2v4Uis9M76SWdMs4XgBZkZD90yZCVy2n0nwzM/wYpbOZJ2VzmxFuYMlVC
azxGuA6qAqA5CoVIQjGAgfuOuY9VfSH37pWBun+WgoAdcStp9Xazm7yq6ALNu5n0
UeqDN48YBnUo93JcqM5sZYCYXKG43x9bToSQveUAawT4TS1OnwNStTe1FwjJpe0m
ejpBekycaJD6gcbFOHFdJvNXrRkDHE220nEqZB5ao6U1PS38Znt1E5ZanuVxDyzi
5RyPNchxQa3Wn0sMBy3kCWD32IZBcxTrM91uP0iBkbynW+tW15VYjhoxvo+G3Y5k
giS4qRHgmhwtshbqjOnucGX3KTX4+qksTimNMNVFPYx1GSdIjBydvgn/hRnwtw9I
EXWPUQIETOFcF9eah3ju+S6s5IIQxsMsi3+EZpz2KPcGx7LHE08BfHY1ykiIcuYH
xLwl9Kq8FdAFdWfFNBMNwXCSaJ6o3hQs4TRGZUBeQ0gHZTH560VDWRgu8URmhz88
xLbE/v9E5YJWYOcDmYGMI7F3/0g3IiaVtKNNiAZUydb1kOOYiFdoEH4jnl03HrfT
m9RnzJWSwJorXLv7vXbE5gogbtJfCExqwgciG475cV63M2XNL2eJ2SnpvAXxL/ZF
AlIgSakf2Qsow0WNM6cwXpLvfegZqvyZMFvwIqugFL/pyKdtWjFe8eRrCiCwHBQz
AJh1ASc52jXNZ62JU73hlqyP/2/01VtEqmt9mkgSOfCdDOvuAMqMg7mz1hRkRDL7
yuepmJluWsCd9DGqJuY7PbExOeCJHrwygIaLp32pJ7igiF7wkKtcFBRe5oBBVd1H
L1T1PQ3Jp6Wz+eyxZzmkILDelUTfALzDkC/aR6BvneAiripMJZsfX4h6PV5P+sLQ
drV7eOmHNGFmfJAknh2QPSjQ5yjU73MTzY0fw56eQ/lDDIZppeNZgG1BQEdgbjzY
A1iTpgFemuyldWdrWymEyRL5zCS+yibHaqCtMYMw+/PYDK/6Pebep8vl+Ze3utTU
hoyKbrFfUDU4AfjSAZEtsbafX6TgWQoqENUZg28TIWF4sHj3jMxIOGkz29nPA/Lo
HSSdLosspTIJuV0PQoco1hSicDOaMk2upy8ccrNtjMXZpMbI5+UdVIHOuiHJH5Hf
UBDWoxt2QpPFMHZdYWkL3FvrZfkDJ5AyNm8W4mh0x7nqEzyqhYsiskgMJcbvHq3j
1ZmtJpmjuQc4frG0w5jtpRy2oktQ9tthCerro5vHsz0QcYpXr235CrEk6tlzTIU2
wmBsXnpLTRnsRFMWKgeomEPuuEoOEo2AQdo/kMtlYUmyZ6GH+dCLEXgX6NWheSVb
+yPLbW+7D1WCDtLsCDybnC2NYbvTP/A7umbnrebHs1Zas/uqKtA5p6i7+tj1yn/p
ZJMRdv4HTgiIc5Q2mv0uaole1Pv9Qq/GLn53GyoZG6yLWo7VJL6UpR8VmmyMclYf
LpZ/27wZYTPBX1v4jDhPCONacxl2qEvSoXtfo+5YTUWgSIXRy3ygknov8CPfuVIP
EbSbuyLlr9JklwthFim6PsnpoDiCDn+PT7s7HNaRYnO/h+LeL/BqlSdQZNGL5So6
mODwVIeKX3oLMfTAmtAI6vbwgtzXNswpOnEuOwvDxtAbjkgyhJ0ANqhZufuCg8kv
ypKVA6AdwsugUxWSItUlPROf3TEOZEEN59/ehuZI181ldBWmqFLxbbT2piEVC6bW
G8hoHaZCyJkfRMnLGxZ/2CAuU0B+03BunTBuIqwNu5VLR05513P0miJjtlfUudwi
QUZI+sW9jbm78OT7orPsFPjMO02/2EcRwFIFqwalgUB4kG2vRyXea8qxl9+DzTo9
eG4wY1KgAONVfrD2KXE5ivIDZMrI1R50WgXQtMCq2+nG/anDyPmPQzf+Bc93Ci0o
+SmY7/RhW90Hz70DUtGUBwYheQt5hAs0gIeL9TlLTBBoHrrAcPzqUpinjR/09bDp
Hv0CUIkpIFAJMFVwpiZaZoNAVQgwUafnG09/KL2Hpnm5B6SOJ4hDfFqytrE3B6Lp
lfTW35btsi+S1msEIj9t7xrQtd7GTr+JYogy04+uu/yq2vWYV4vvv7JXgIVxAlhe
VkUTDZ2okFMKbT+8OL9Lw0pZxNmdZ9+KlUKiGwN4psEOZQXVaIdAqW4hPS+e48JD
k0+1lG9oaWtWhxRoWR2Ryut0fVrM1fArNkBvShP6t/GHWAmWU3o+SGJ8gulK9m5G
lCG5XlK0yqidE98Cn+nmxRWktkZUywahEm2GK/S2X7KH9xJ4sGsvtLgTtmNwNhqr
JilJFB3gWPXKBJMiIE/7GilKaayvtP/kO11AvJM0ii8qr+kk7Xv6szwy/XfLChV4
GZA2Es36yXZu1xvE7TMVXBYL7xzTKDQJtxvbBU/T/EaS6nnr0Z/nHjeY7E+AHi1j
YmFsJ320nbfhy1v0SKw4ngHyGds4auRtEaZUQ/aP60m3au4skA57PIV99+xvwK7y
h5p4kl2kDwJRD65jb1tmwvbdq85cquCSO91/rMPdUt6Qguh/gMf5hHk1L4NhdIMw
CcTaFuSSHsp45Hne5aebXDwh74QDvqa5VeDXf7u2A7Br8JUjT3Dc5QGgRdMXTIpg
eKllAJvSPXeyvrlP/a+7ERQhyYkMmU6Vo/Iw2WDqrwETkymjKmzRWoBP1FLbwTCH
5suZW5IaBRO1lPOzcrwTDgNN2gVCh5wtGR0b6uqDaRmIlnZrC1O6cpFNeFoEyIxM
kqQzWGRglbg+Yd5u74MbkqYXlwNLTSi45M504PbNeo7npE4Wxo81lVaYBNln1+v0
hb1n4YMxkiA85BApeJUdLMTwH8dDoeKbuhx1aWJncoURqnM0IIphBpDbjJr+V3/x
x1wXuYl/Q/HBn9+O4gn1Pss2Ybft3TqvBbMLeGxe22QabqnWv0ba/rpwkpoypnRA
swB1oXfZN7Jbvk1IEZFChh+QfD7/yo/2Z9WPAcHz56yowbG19C2qlGW7mEsLAwcL
Ld5UGr+Wq2yEuka8mM9Lqm5zvBJWJ63oBeWOs26bHWn2xE7eseEGylVuOqt4THv0
4Bn6HbJ1DSqT5AMCRVE9vmv878NVQX5hhnYxqGUaWDFJLLWvX9GNYexs2FIOTwAR
2Yc2x7SQVBp/JT4HRFH913e8ofw7OO1xKlMHlOoxsXwGO94SRHNplrBxXLVKadKZ
0AI0eFulgw9NOPtrHA1ajeHdkbg7e+KKVwBhzBOsNFA+rw2659NU8JpvRFhZNN9O
cfM0TMmQDtuJDBrTlPIcmbQa2sjnRqAJzGksxBMPkR2Q8mu+C6CVqOfcerjEt8Nr
//s8UXUiG/kmCaNpnnRGT6WYxOWYj0IgrGZLqMgo3/NovKyIUNTW7RpVU/PsGjlz
KOgYA7zyOJ+TOGcKaN9b0NQVrPm96C7raheSBC7xdHrinSKXwJjVuAtc183OCKiC
E/UslIVzKEd595Znh9g9VKWrkw3Pa0Os4W9ItLPmECCbVIHjVP6nAC10XBQHB7wH
gOzN0izl/xkuGicG6Q8ZGOerDxgXKNl0gVprlJlgi5/Jrn/m3sjj1Vaf5DnzkghD
5IVLrwWCqc2iTVtwFlmjs3srefUFOK1qGyomvvSTOdL9ERD+UItwXDWqb2hHPbWZ
GCs1ObB6PJMqnJrNaLhY53ApBrYoXhPeDVCOvyXjSqihPadkArHInGOt46sf+s7g
yCb90b3rR1qZ3joc3JcwmL+kcS9I7EvwNQynIUsn4wWqTHNf/FNbtXTqtDiKgU+W
uhxRAqCdX+sapujbTZ+opZdryTONYCSuWnZv0MzHNJBzgBVTR2vLQrR7nFe+ZYmx
MY09wvSMMS+cqJqTrQLYCzmmBYvmPktgNYrCLHOAw1fDyeQEMRrCCr+bctAoydjX
aO6wAuv0SVkt+Pczlljv9K9lIeZDParbWjrZRzGMPSra9bKH/bXrBEji8nWVKkBx
VXDGZxYyQkCFpWY9mhQH32sJEU8PTT2vClD2R4bqiEbdU7Wlb6eTIrYdvK1I8IOh
CpxGSKjNi7Gn00Hl5OpR0ryNSPtxLmZUwhROL2I9hOgs+tabUUWZZ5MMQmNeEqFQ
3HLeIvM3PJTNmmu+QB7TipGQJ03ur3/nTMhqcMbaWTD9cVoTzFtqaREU5r2mSJ7D
eYCMLTBY9pneRlg5ZrKRO9JESgq3lFt7+tGAeUeXdURxp2BAOnsO9q3sPbDwi9/M
YUWzKPrjTJzkGvwO0riKlZ2PY2OWA7o1HopS99jgN6sOejwit6pJSciYCYRTDUJW
P3m3WQLndp0NEs5U6NI8cyhmKSdoaDMnZ9uWPmUsuJmQtUv0Kns2iYrrbwTeXPaV
CCtdzWnsoJE1aGameAQC5TBdCeg51fKgWWodRWjzlczbcswnspanZvi2tNwn+0Ug
x61MskweKf8FKRIj49hTXKh7bQS2CG76RX08ghV21NvAXJI1gDi7sTcq+1SXFuZU
53yeygnBiysz7HHZmgvFdZLy3MTf99lXvAzj2swIuMSg5ByivlAA4RSZiHM7alCk
xSaEXFq+jje1KpzF374EBwX2QRuobPQ0mpDC5aApNT8XOv2RFeXgk1EnNuYFsyiJ
Xd6jCQO0BFXXFx/WGBHl84H6gd7BsDQsiAM0LNto4fffHKshpf5MvGRnYzFvk5a5
IfNtFrWhuyFMOiFmTvMpxdYNsNtFmroOdmNxYhGEO0lVHCrazx34cpfVbHphci89
ddbBN8U9LBlOapMt33IcjFmV9EqQ2ddCb2kvMDmXKzQDVhfo+CYkajQv4+ami8as
LXrQHTyp03ZSaJLsk5bYs9TqTvMQOvXd/z1NkIXHNN+rjFgStbJzUNuZ8PtUkZfn
J6DjZWmSoFLrtsvMgbWp31yhwuU4ngJVozG74/RXmDbrJ1qerkKMb47PusBtZse7
jfZIrxCqwhg+M7vUzUghcj18ApQ82CY/bFQws2Fv0MIVY1MNLUZTDKioSndhPprC
xJsT0ur9q/TYm6rONXuYhypJAB0RVu8xgGyOoR2ygDf3bavu3rAFIDBxWvA6lmkK
vNKoL4qboAGm1qCxuIafmRwdvjPTrUSrYwNUQng+E67dLnzSB6NSo4q394KzK+L5
6/2mYjKmq2WBARSlX+eHuttuSvlaiMRJM1nNlNJhTs5FCodPvWXtLpT8tgz7GTKh
NoH+X4gSMMiDyJTxv2YTY+iMBc1NEVM+TkmTD+g1hUDw1CotBNDLsYnA+T+57nbp
EVJ9LNfxWPXVcJ1hDmac+VIloFpkq2mZ6QIpJ/Bo+K0UqSh6J85Zkj6Zquw3gmOV
vAZJQxyNhOZwp5lAzre+zHjCo/vhAHLuXjhY9+CnCWitBwzMYnOsSaChDNlSEljY
oGDz42IhBH1StwQ2OTITOJWmCGHNvKZyVqRGQ9WhpM6WWBMdWB8oEaxUBKl7SA+I
HCpRgNIfK5PZcfffySKFNiQlgGQ+mKB8m1YqNZszgBwIlBfzHbOUfgMjrFH7RqdD
25iINBtSE5eUfKS08OtTroxH0ABlTf7CWEb74nTCkZXKhPAUD/NKr5N8kbJd/RwR
UDYB2h2utyvd9/RFWX25PXBiPl0bRtyPHD6N3ESO4Bb2SvLtFqJeLXnNrvxdzFcT
cvxNIh0mTxe9Le+M6Vkv4NvPOk9EAOfy7+Mffoj3OoTqysU3m5TfgLVYr7y1T6Z4
gmelDo1nVMRhJqLkmcH59mC9fcsOcD0a3To9PGfAdhRREpAyxZlt62Cj8pvFv1Fy
KhFeKTWmouprltaP5bEGCv46VdAA+Lne0og1+BtelEU7svBn4W0Mf9NY+wV5Dqrv
XTgP4kZuJA1z6od4UD+bEfevKrdlV2Bzai++waNWdRqt7IgqGxQdoV1/nL7KQB1S
X78TZbtVz810PhEH0nUb/DWRfcrLt5+lEL4bG7WPje41sEaRtBVTHBzzGI9xhaDk
PRFkt+8flz08NhNvogTgQ8/NTDwzRzUI9Bm0SBjgakd+aOXCc/q7nGAGZf6q9rrB
3oLB0MKjmTRUg241DjnN7FxTQ5biYAghIoYyVA8Xer1PpTr/0OabawJ9osuk6WxZ
hE/TFgrfBwQbECfUnqZpUMiLgqZvkuhzEZAa1Rsp+liAeoxFJ6OBkBRaHhm/EIcs
ZPBEuGohsA049zb202nXeJR469NHtUM7OrxOQl71qA+904Wxli/P6BL2VpmbJmKf
eF6PscN50jvcVlMeTsQxFFV+OZWQINHn9RY2fxdVyvth6uF4KvBPOHSGrlsaEoy1
yNr0tdid5+BEvElIgv3MqSMxSocXk9llxhXRsstHWGc8aKS2DksBIQTBCOidXkVP
Vd7ydmkC6E8gv9VpIr5v5roWXwUB0Xhbfjh1iNoC4hZ3lKXApIQoTSPsA4UUMc41
QCikR1Bwtjx2T31s722YT2sD5+ZLp3nM2yydWeZl5GgrzYj/RKpdgW10g+kXaWlC
2mryjYvF3Kb1Q/D2PPfOIUZVcB9dfeXba2pzQ/oVyzX0qXtxlRuFwI1N+MQeDm8x
2Sniiy52EIOADVSec3AXQKYPicVuDIqvFFQLfNc9KF842cSPx156lrTjG1VMrr/n
vqf/UST2heiQiDEYiubno3kQNevGdLFqaD749JJSDZu7IRsT998zYEhDos4BM9zr
wEkAznQhjt2R823q19oANROU1O67W2VmFvfmxq+rvoQ0y1g7FPDfa2vlX4p0fOyI
1AuKzuNcUEJNyqnovF5M9lKBZJVfcQm4MeQFE/FXP7tGfrw2mueMzNP1rftkbQzL
yD60rPzDWxBHedA1dBPNZJ/0h+EyH79O4PSMsd+0BlvaliXKQfR73hSScOwLPXAb
24bA5inG0eNOSgM/6EThAsr1deIFlfiiNLvy6cY/pHg1llaNC4lfONmD8EXFuwGn
7HFvwLremkDnloKiS7Z5M2I7gF8TdHK3qM7GGAtVpublorttVTYnslZNX4QTvfEu
m4OvfB8/glngfbAl+zDjKWBgzSCXIwpYh+r2LK5T8egq+x6O3Zjyj8ILiDrvWEcz
nfvMmJ/9P4NEbQgUGhNCKHIrEJcUV/+91ifD1hinRm9eTsSybGBaFjBOcU3sVodC
2Xqy1oUIyK8Wr2akXqJEMdVPcE03fTTQWBvZk2Q6iTl5kztbb6SDqcuGdrZiwFs9
5VwE+lga9m8Y8vfM/PsMrAwIVM/Pe89cEHxf65mst9t2x/Kf5Umn5qRlx/pdfLcY
P4VkfQHXtT8DoZeCvezwmUmpYlCuR2lsr66IOE8ovYeoYoZiwlQux8WPFhWN6QPP
PQaMQcXiPI/yS9RC4xd55e3EZLuhap7v9nPbnqz+mJu3zpa53SuCg03j8/nMRM0S
T4ExUzOjEwFLC5T9LOh2ECpUojvBQ/vGn1mEFFmHpXTSNhw3dAYs7xmy+//WIccE
0eRBJNT6uN6G293mm26x/LuUXqQCLSTokEVvLoNSMOpcGuSHv93jfvk3T+zg78xQ
It7qrbeDxCPJRuk/d7nWT0nln1X/YylZI45d48OotDl+6ruE//dwwzNRcCKK5za/
Vmpz2pwQwc//cEbQYKCLMJqtB9U4u516vYpct3xuO7G3NergfE980Ijzaw6Hq4NS
Rf4GEhkpF/WrTMTO/7tSeaoKy/QuRtCgt4eMjsdb3x22I1PsojtWRd+LPHufmLQH
BHS7Y0gbZzYJk1kRczkhCVktNImejCmVcXrlBnEOIdZteCG+vdFK18SZLvgNNWKi
SncNWXzfmFI1PXkZ/2VEFdDZLQ/JJkCJV6FWD9Wh4C8YWPrQnM7Cye36/tRCio/s
v+JhUu+neOKtdXActGNU7nKGdBfP2sCK5938pXnupL2Cpk+i+fLSnKuOe3eQTlHI
6eDYplNgKa8KjgcJVGzw7ViIcStSrZIBbf2ShmTqsXZZpawNzVGcxkVKuH+kq2PF
B35pmJQdehub4ZZO+Q3ikhltA/8W42229BfSbrGR1SS7ph8xU0EqcpNU91dV1jpx
zaOU4TRO0QWgkyJZkNhgpAMDj42SYCN+sbDz7N65jso2CmdXS0fec0BCwTEJjz1I
lZHX0m6pUM9vsA2u8MgJMxzGctxlZabQlhlK+hK5rgcNvD3ZiTN6k+jSRAX/n/wL
IVhwA2KkTGH2b3K4ks8+U2TaM4w1/Qjzncq5NzB+5OqnGc5CJFBib6wkTFv6q8tW
U4E6B0X8gdAIlkEhYF0brJf+gN9v7jwjoVsqL/YOx7cDtm/RyHL1eDtmKubb32Nz
9keBiU3TalKimFfaPQIvjuJVlI6U1Ft2nB+1eE5iWaS2+4S1dCRxUD7tjVAx3But
TwNUseQ9Zrj27Q+u48y4UEEwbVAxaFrfSvd5JUBJ38ZQ2CBpRT3X9xh+KpQaA4Ao
lWLcVCvTMlNEBSO0JGuxazq74DEe6FKJBlij32bF2qxetdQPEQHW69+v5K+isq+W
HhfrrhYUBF2Lps5s5VS9FJSigCcHEs8cFJyzieOT03XagecC28sW8NIpqEYWZR4I
JGLutqFkHugbkzjn41HLqoyZFvYuWPxS0LQOdxW0UsAKzSm38LXjNK+pmPY0EoUV
RljIc/GfNBSoPDndSsLXi76v/Z3+UFL/O4iqdyLB7dsdZNY1KAbBwMjiTPJav0Ia
x8zzT3rePlVzAKqTY88VTLloKCau0BTMm4er9NUPaL969L7UyVpBGZA7M/8NTwbx
nZ2IYG+bz44RIAeHjq9M8rYRApp+cSf0gi+Ewz0dcV5JdwvyZpEbqz+KdAa4n7Iq
Fg+akLpQAYbUyoREF9OpdJenHOIwHnsG2qHKNi4WKsthEIi7Laij6+aIMMYgnPKB
HFeZqBcFHFSbSlnERBVNv8dkv83XmvCJc6Fg0cMUyx0NGsYVRhK0EBHVnLfwZU6e
Bp64GvdPLH2iHMWZKiFdoJbi9ZTn8i5CSw8HZuqpARbAATp3e60yGWwH4IZYQ02C
rXbaM9+Z2rehnmd4Oy1tLinJ460y3OOE9gntOSO+87DmsooQHH+WU4hKUW8fFOUi
t1rRW7LeFKtP5DjfL2mYYxQXonOojwnrKizUF0ar5EW8PjVOYg/1dd/KE7GDaKWo
vB3/ZBoIDp/e9OYYXg5youHGcnpJldyFbujCeKO4l0V7sdGqk1M9gDnO5dMIKAa/
ngYrZrWXbry68jgBuwhDik6ALCSiHSpDiEzGNvoGtERIIXxWrvisq5MuZ+yxz8jf
7EaXv0UytbotXN+HmcHPAdL4+jPg4FMEbqOzVy/Yr/nS7ea8n+OmRj82VKBo9d+C
62wzoWxGeFuncMIVr5uUIDjsnsD7Z86RToCnipfGc1P+/JeBAY0EBupFQ11aGvw6
HZv1vsK2Jy5wRKCOxqcPCbL/op7nQLfYLKwgIjQ24QQ2g/BIxK/PJjOs7S5yF9wN
jaaTYQdI7mdc9PyfjdnJQCBk2DY2Gr01X+OLIDPxPI6RoJ7RzgXE3GXiwlf9u42N
DBPIzYBLSd7bKB93tQweUm2Inbxp544OUXsSqexmt/fBPrUAP3HhX8V1xM4aYFzn
MxODfhn0pNvjw7IpMyP+JH3KdC4OXxsDAF6unxyOUhwfJ++8SkXF1DRuYPNggDNr
eqAaPDKTDQ4zWYBE8GS7B9BXtvkTUP9JGrFZWCjykbPD4UIg+IB39OSu6v0M4lBB
grRXfMClpllQRTAJET76xq9oerVB0c8QHUCwF7T2BqKBFeHvPdSXXnxNsAfZYA/w
Xy0lDjHYDAhyZv+RIIRO1oUUS0Kt4kzorXX/eNgKTVdTc97MTns8J8Xew6g8+LWK
96rpLeAZJOIRtMyLej25whOvTZojNsrb0MK1JgNE/feDJruZyyMI3u3feehrKKn/
Lm+bVJ7qqCqszopGL+8zjrP9Z+/L/T2APdjFPRpYKn6aoaQGFiws4OLjb9wHEHtZ
YafkzDj5rOFRtkuo5/BGcEmkI8hQCwFw+LVzN2umJ3tOZw21lPKgJyp180Mf5bB5
4XtK6IoWWfBWxsy+H/rTXQ7Pa/Q9Dapf4ps1WwI4Vyw7jB75R4ne6PsBGXrofZXD
bDuKNLLUv8KflBZ+L0IIzb6mNpht2ZdvF+gtyHqHatx/nacB2uwo34CPWTje/u1L
6PbwLabh/1/dljYoPPweagFqfnpv95ba/M92B7Bc+fcPlkzXgFFSECOJztGoeJJ9
xZOK7mEgwgd4ZzO8HLZLZdTFL6dAVZrqrt/u5bzNsnHdbenehoPJ9o3BUW3RA3vw
RYGJhetZrjDPB/+e/JNHdmHkylV/23lnCol0APPGQYouGzEmcdNyFKgH3Qm27YcQ
WYkz58aWokCFhxeUPyAQtMuouEusE37RXjM2BDGdVPPORZv6bkQA1kKUk5HxvXaV
HficoH8s8LKQYcVYz6OVcLntPHlnzMo2PbFqXUVnPi84KkIBmKuAovFZ1onZc2L4
pk325ZzyPF+oJdma1ITB/t0UvQ5JHiqC55txmA9UetywRTq8f4ppdaLh5zep6EVa
R3UDuPyo1KFGIYXsNjA6MKjvhTxwxAraY7AInIivh+OOPYBJGCKMNfb/RnrGI1wC
WGg9hL1sfoA8HbNwPWHDWyLkWuQxBKADNdsGOcY77/elnCmGj8mGEShyHSDgmqlX
y66ZPLBOAHLHNCJOEkg5Zi1LrhUCj9y8CLiiOoIsup1VgBI2i07yZ40T89QSbEqp
YvhPC8smN8Zgz6lPMqDkVcPHp6Nq2bJi1IPYo4bbCRIrxKkmnWPkeZM3JAPNibJ5
clXhHRviZjkLnlCVZIiFzZkvjyxzQu7i51km9zTNK5a2sG8pqhBExeurSrXAe5g4
5/jUCqaG0pknP60rHzTdcQyyIu59PIb72M4C6f4+wMhmCKsawxpiu18yMBCeL33c
2Igva+7FeydKMJye7OrrgvtxroUi3g/6l1skyw87oBZhl/rEcMY+MTaaI16/svuk
476dsvO6X0xQJjTDYG/9/rv5f9qpJfVx+K6Vo2wIUQk6Y5JVuQiwwFydUqccr1PV
4V6sJ19+SWNQJJFOp8DgsjEJXKPErcWm9Isylga72EzzbzLVf77qoE/Wyiad069x
1eSHo3huip1hQL/mBHeUFCNpo1QzeyL+tVpHa7tHNAPlWERxhuMvAV1fVyfaexsl
JggIT0VvtAhqpHAqK+C8xC95VSP/q2xvw7H2nIUIMwwxITcjLZNQuYeYZ8dGyjHu
TmScocMVF9MEiZfIzdBarv3K9eLm+A8sHFP/SvWmVsjNdWw+6wFsFaI0e9S4sWoO
CVOnkV6mQDkW18nHsgdzApAv7L9nK/9X1IjC+F13XffRV7bgVkKq//8kVMDGr98R
i0qY32F235XgR1LEWMjJY8SoccB6Pwf6oUIROn0Xia8whtui3CGb7luPZrY7xJJc
xveF/lO+netDahQLy4XUG3mWHznv7csfWoQhNVYsx3uP+MoA6ngW9l/wN+HeWIWV
bSSLRjhCrEzg/RPrHbiygW9rXpv3KGYlS5lxp9oD8IZNIVBaGIXraxJgZp+9jGUg
sCXjgkNRe2ToXYW8HxLxDxgOfKuhhcdtx3GZ2CyXoV0Rl2g3c7eV8Ib+DtTFSFcE
1Jk6UhWd1CslJH+tJG/ysJONWQIZGhhTn+bODNfPcG+ANilxJQ4Ag1I7VRCtN1mT
6a0tN6zWFVYciLU8X9O3/gphKbhp8eIeK+R8CeyosOWmQD36qvVW1B0lnN9xzc9y
RGXN0E/sTi2v2Qznz9zrcGsqZdC2ROH/Csg4i+DWOIuTH44NndvjftGN7a9CvXnI
PiNGADWbHgjkNvMz1nIFozeKDa7GNGrHG7TnLHbQ2ktz2ESX9jfGkZx0NG02/eZ1
JFEa0+T5+2bbLO4s7LENe20QLs2f+w1FdfCJclRQE0gJw/FhOJRfoATQRfrty2EB
tbkTdKS8Elnaph0dGSI4MAPLj5mJWmM2CyNOK0ir+1PvjhiUokbQNjWQ9UrNMFyd
8oo1km8yxQPo6pliQMdj9xa3izl8Ji1szN6uNZckOKdVYLn5MWlJAvha7Vr2KqJq
4mEr6IcdDELQUpl3VfP3bK3y4S5kaax5CMo3WuuNpp0c17kZvypfYxbXIXHUbUcj
XMlDqYRyDR140nlR/EjEEx+wqHQR0Ne8jvLCwFNHoGOdNFhO5q9SdFt9wcJwaYkl
Pw1bEFGLIduXlfbX1LAbRsK/LZN7bF4WKKkxCaEkEckKagdXmPkEe7KwaTclQ7/j
yN9zWksfeUd7ZPT/ifJS/SkUK7kI1rJTs2Ym4O2xHo78fonmuM5V57/Mszgztd/n
oGD7eZr4xVJal+Pi9BkdaFms9oCuj0z+StVUCORsMBUJ4ursBt3jKoJ22XJg01fi
8Sm4VFfbSYTGS4oyqfXbtls1zGNloW+1E0K4Mp8Kj8oHrbwTfus+hKe1kh8ftGRh
/8KScZmYLYA+hlUqd3jzo4AKwL06/VCXWJC7E6FCvHMnthuYHX4Vs5m4c1fZx2UI
c+CADTuAsnzdb85vN6Cu+L0/ZklBWW3PVl4hYNLW8auqGQS7Qn+3TzPMRtIJzTb3
l6WquNsputAcPlPMlpKLNeXR5Bq/YsgFkFMfAPRoAq/ryl3Q4NOiuRajQh/olGFU
43M3q03gro7MUvb+FoHJ66hsYYh7HciKvwBLqXz7OCuh6fWfHJKN6qTEJAGSQcC2
rTktAjrZ2fbQoQLQR8ucuCi8ntHJNWq8T0bhuTN/yPXFMyvQkIJ2keXq0l7eD6qr
ZasIWrkOv45edDo0+6lHhc607YCNa+Fmuhd8ORGLTclm6+0hGa/ZDuULcMgjNDBS
2fmG0adfpB666/DF2lzMosJGusYziFR1Stx6QrTdhAyjgGltqyFVZaqsR3mE6aaE
qhtCMm5BT9AirIUszZX9TVw391fxSu0ZH2KHfplSAxB6VBv/vdKcwcPGAnHvK21c
tXEHtEH4ICh3vDl7LT8IZ9nz5bHe2X9loofhHNIUd/mAzo+L9cpSCyrVn7jxKYfY
OlMOZb6zAAxmP1tXSmCk9HJNfr+NHLXOTO6HfOv7o6mtk3a67FM/QPfdkuoJc9cD
/spwB9fc82tDHQxzEglSgktoQwF8ZaU2NyqfcttkuZuc/gXltXoXPuVtvgIpb77v
94fVpnkThEA88Op2rQFxWq2nMzkjLn9jSNJArpSPzREHmXgc+C3ELf8MqfI++8iZ
jR3Hr/zEQY6oZQJvWfYkq0XnG/ROgSJVs0atmRs/DniaeGqqd6Gvsl2bNtYHrUxF
0ZoiAdCJgkeGOlUgruP8oFvNC3cdxfZrJceHR10bl27u6xP6YjBzNOHe8p2zIO4N
xo875UZPiAMe9MPJtJJLBcKGZEDN83zEr6tj8Uq9vzAmlmH15NgqIv+7edeajQ2O
a12DJ+UZcU0B/FE3LM5b+H+WIC5KJ17e/1V51E57hZTnJJehAhCcTMTetLq+Gymt
52im7ZHGKJs9Uj0MThSerpf2P8l35IWk67Zc9XZVwff+0+jOG/oV3TwQhefy7mkY
H6LhVRHtqk6Okm3rCNgQI2R2JPJrTF1vIioNZEZlZQ+MQUP6t9HZLaprSf73mFAP
1bnX8CP3d+9ZLSXtbM1VLyiJM+4ZKhRTPGkfoRXbENT6baF0n48EKWpQv53XB0Rm
ZxBmqF2jKcG4WoOUSAzqKbQ+XNmqgVq7j3A/lLVX9UJ/KgUUUjtuNcx67hfVud0d
Lp3EuiWfH7EyNd7ucisbrrJ8BhFEm62W0wPkIx++8d3ln9MXxaN9DQxZ41iRTRlX
3wllsS2cHl9LvNqGhZwVWcUuStLi00fIE2MGZyP+hXdi3Kp/uwH6lA05515uBllR
2RGNx+FEZuS/AowDxNrNuuWTqRv6ucsjBaYoS/fUqu+HpZH9GfeQ0MObbTMhO3x/
FEUcMqc/TV0JUtYEKlzxE6PKgfbQYvLx8tVgrv3KLTz/ClqYP7humHUpCJpwouvR
qYyWYCUWx6LzA8wffTorjReC3RqmHHhcqMSe3oxvnw571JgSxmTXJpp01VbwuBni
5ta+640TRfSFc7eV7l5xEez9//4kDAoHhYOfHRZ8T3vEVPFYMcEa8WAbWdkl93Cl
8EpD/SGqoTEqqjdheUrwlwsYw5w+Px+3f+6wfF9b53rnrVHvs6Ed6YbccrnCcI8E
DwxylXraBLdScpkVDcWvb183gzJkZ4oURN5P/X9HoU0Md7jz+mUkP17VqkY0Vsoy
7ilpCxinmU2GdTwmBliblQUx98y27tSSJdYqw8FcWehvy/J+PrfHWF+C0hh+VSXV
+IPzbn0eGpWztGl+mA/v7BS9A8U1Lrw6vQlgyl4la/rNS4V6qa5QDrDRFXqySb9f
bhmwvoJhYbHeAvSTYlFvAEkVGF72x5X/0uvrRLBqcE2+ha7MUDqZXUyBKtubbOGT
5KweBbqE/hUEFWxaKeu1MiuYu5mRcGbgWsGBE6LQpWxMDNHsrYq2evbe+jP1WLvb
0ork6Y8rSM1zqIQe6lTLb0/rvar/VwAhTy+DdZimvvQ/CzIEchigIwMB8kt79l/x
ZTzng/ANFGViGMSrqckzJ59e4mu5bZqDwYOkPH1Q5k9pcRe5/OdRp+wGI69PV3gL
64AcZZU06MCk67t8oHIGkypTXMbbBbXDW0cFwHis3BSCpYoV2wYxOaVC7r9dJHrv
01MW2kEvpYhCAO97Lr0ohR70hnD2IKrFvT7zHigfDSQDUBimq3psGRRt44cgkm6P
Zvg5x1r6JLfvo7HDFb6JeUj9H4Vb1cgBNTc8pG2AwNJ0RrlqrfM8c10Eb4je3mYz
d9BOptorSmguOQt+NSvFD7ueGOB7a+q6Mj00q50BNGY8Df3G5/IfMfXngyW6hpms
9rb4ewDsSweZb3H4FcMmvB5kLTopaVsfiz42LX2r80IXWK1Mzq6HAkNgCnllx/61
MW6AUddT/QW9Yiva0Qpnt0qU/xbrJER/sFiJglQT/qYZE277NTIE0ngTTov9vonG
9q+W2G8PCA03rwLoeCfBx3Yb+xyy9GdeLCMDZQZ2akOwo7oods6hzHHoqW1/YX57
76rEu9vKyeY9zixRogim+jSKq0TEmBkYMLmlUkQw3H57Va2n4y3p/XxMEgA2hORW
0QmLr0vEHRchuVifn6AoGc/S+o6N+pMi5d9LNf1nOA6z3Vz2bU6byGErJo5hjyJB
TKnZeuCSyByZaS77mI3/k9mjUDqTygJ2MDFSw19pHWR6Up0RPT7Ul66I/5F/mLX+
pALB3azT8vyKHnqodF9sB4adDKStvol3GJQhCQNcNmsdFInda2YSMT3zGE2o640s
n5pf/VKRavO2GfC3ORZdqllCKNFavU+tEWoT1YqRsYJWTUdscBe1UwWp3QlooJW8
F6cc/3KKkVZEVv/Z547qfyzii+8SL1NhI8eyZT0USIp1PBUGXGkONMFLEScEa1DP
lN7bFqffVFJDn5j+JUMLqExkT/Npz3v4vmsXIY77Op7p/+6VE2Gs7fYMpxyM8YCQ
7K4I4AZbrd/Y1xS3R/NEviV05Ff4UJabJPP0RIxfpTJPPL/shOvakZyGXr2FEj2V
ljrE3HFxfEoP17of6mdgkGzaaixh7xfdmLCFVN6GuEkTmqNuC9x/eiAE32gRjxRS
t02vDiqAaVsm3Jzv1SiAYtHVXrR1SLwQuuwFlpEdxabyIsyvO/rv6KG118kD6rKl
MQq35y9Y8BaIYF6nE2bIQqNG3UdWOC2JsTi2LEq8lfuPRC+qn5i5FIJUl1WhzAjA
OH85voMzoX8NDLX1ILiw9JwxLbOydECXJ2RrbJAA/eTlPTXNdoU9fouIahMdwECY
EKxR/5w/LH3VuquN4BHrunohwUqzXq0BgLtgmo+erE7kktPccIvmwvSDzXk+3CD5
g+ZIIR1gzm9+xHwtlXouz0G66Dn8RjWjNZhZrQR3amEej+EroaasWn6wFovshN6x
kIcXYQ8OnknQ2/s0BAJLKJb8BTHJoeZH98kf2FIFpsBqYETydnS82O/22GqVrXH4
tAA7wyd5cxJlglcyOpf/QF1kYk2IbkrsBGDuN1zKguw4ldM/9IELd8DslDKA/OGO
W9h5ZoBEwALH9Fcw+YaEk8DuyPcTHEPjikLZMi5QFdOr3+3HjQnMsk/OFoOYquC5
P4i7EkxTQXBR9ZFo6gH+LjxyX+EDZ9pk+75tR2pE3urB9g0AU8+h7mbtgiIBh9oL
RmSvvdcSyu19swEP4O9bJSZ9drfGoZiJMNwFaNBYcHft67zjPac2C+MVaynK+IfT
HTYmLV5rjAmz19YTPCTO1+T/1ho6nKnetYCL4a3RCwYAkmPujY/uHXCoLs9wlOo2
2yM73r+5lWJTGd0K0txEj3dVLUp3H+gxttp4LryCmqis6qws0qUvW4o7Qf7vVT4f
/+cWAzvXlzkdrF/zlVFg8qDtpnxu7ICOQqjCc0oHrSw30r8Rpj65aC1f40QGkTmK
pyzG5z1ghlUBCa9pWaGXJIOZflSmTIg9aCCmvjTlNHfb7pkYTVRoXesANC7MlnCK
alnmIH6gSeVdGbw7gqLYR4v+JQeC9HCmWFjkMPLtnvgR2Ho3EOZOOklEB7MqbgTJ
AuhxId17ieZhZR+I9/U6j01YQzV5USm3H8sVpcmCKHaaX2CX/FtgtYXweyfK3Iq2
hvP1deL0XQe3hQcNSIyKP7IM8fiC2gUlwk9+hYuu5Ld6aZl1dgByEgD/L/g4YXyW
SZgDzcutdulTCqcSzMCqNzj0A1kjnTuGAa9foHff0239oj5uRfnuwc4EqC3nhgrR
T8v/zQaVgvKzNUsWzdlOAdCB3OX2EH8rgA1jQO2kuqrUb80sok6FhRbqsByvHj+R
R4/3Za6VBMo9S4dy5x9M/f3fn4XtkxyT8mIJopn8kxZxStVtzuEjZi4e04Fy0lxk
jfU/6aS8Iym79VCU9FcaPJmajyZprc6Ux77zqwk8//xaqztsxluJ4tRIsyj5qjlO
MDwr75CrrxJkveK9mDG1Nm0OyXLaqC6zmLqZyTU71nIAivf4vQAOzbdK9Cb3077b
VGbyH/WWm+EwecDeR8PC0zcd0GznUJ2iMKLmBEFTn+ArHaOHXl7JrbwnMAq8Kkqb
yyT0asIKhLVuUdhPYGPe7UXdY913Q7uWfsVjAzZDGl8vw4D4+hpZgoJz7ohUfvcC
sJs/rlneqc0C6yuw4sfiM5FOYpsfW0AwFT302hrcIEb0o4XRFUQ/G1ETGQirPxBH
/AecqjX2AxtMEPfI8OBf5SrbkSA8H8fEgkLhS6DTWdVDBOsCf5Nnt5Hqy8Obo0E8
+ALjrkcZob5QyraFoiwFb9QYGlTefKQvs8/t0uZDMFYVVJWm3gowYHh8ssWV264p
uCHerl6L+s1RmSMOq2Z9yzvtvCmzOqQX55m5AQdcYlftFLc1Cy0F9kq3t8RItViF
svyBvv7rYCmjnKjfn1W98AxObxOP4aIECVUFrmvQ9Rseotp4T+WGoc5LBlnxFjcn
UU4nloPwBkGbT1vuC+4K2vMTTdp6ikFoZzGfkxoux132WN/mPTA4AC6yArSAZL5K
XkE3i7RnRKQbGGyr0Ont0swpymfbSA0A619k56Xi5ATiPXZ1JZxzr25SBE65eAe+
YFLwvIHkcBjkHCgoPYUJlrc8S9VAxyWaowr4JAOkLGJmWJXQ2qFBd+zqxgwWjmyc
ISrEpr9qe+k/rWQZTGKksTnXGk+erP+33eNGiGYyXVelURHODOwjdK8V55cIcFAr
MCCf7gHAbWTtUfP8I1VIJhDZbQgOF9uJO4cZ7eLgpHJjLLklwXQMMxEl7DPVZ33y
da4g3O1bjwkDMDlRRDPwYJmJ0B7SL+7s+rYyWmDDN8L3UmPIUaInFsG20DO71KlR
5o9o0xjClqnMkEK71MB/jcb3n6qq5+VctBrxQiXCQxp2hPT3qMoyBg57Mc3ovpiq
kZpT6Hw2Opcw96YCTiqMZDdQECVSDXvjgFPcfTMOhExq1KTI4qOY284IB1lBk4+k
eSZsJ10D8ivXB4xQzt1ZCCFkIGKAnUwd7FCTSsES+IYOKcavGSdb7/7910ZRpR2U
HdJekQjhq0P/orj3f3nILss4PKZFP/sNFZok6uzcSwr63Ve0SAV3wep+dNAiyfyn
uEEWW/hZn9eMnWuIudDty5riXQcm7w5E4N9jCqGF9NLwb8/YPtjAXdsd1UaHj/Oi
wqg6wmf3hibm1FkjTEpPSyit5kDgqTrx8PzXundv4KnF1w/3EUlRXekDCal50clj
LbBfu5lmn0ZTEhgQ8Cyfpf4lKs0WC8qWMqmlHwh3CSoEeQspthRmfMPNUfCd9Eff
tPwEPalvw9p7D8Mh4FtNIaRsriq1fsv5m1GPncD2jEW63DUAbPVd78LrtnY3YWcX
cU8DbUyog2OLwCvDqHhR3nMPXPvEhRf5TtljK63EwAljOH505qk+V44ClPqgseMh
rmxoPpOitWPUUPvoI43oJCu2Q0JpzqmmytZ7ilWjSqTqmv0kEY96yDnZP6iX5RxV
6FBa9d2GI2JXvT90ji59wWyO/5G4Pwf4UpCOHyw4Dru/kmqfxWv9jTrlVYE+Ri8q
CxodToBnZZX0Wfq0iEecQVsRpOmnNWv7kWiBFUm5jQPlcVWvVRrTX+YtwVi3LLT2
N3EIQA/6eeb33PTMnuHSShI4w5gg/lG4NntcTRLhCTu+7FtawU92soLpViqaUrs+
fmznxzzQNFK/VxgkhTa20eqhrEs5RM+Vr+NZea4MbxFQNS2GnHCCoUgZsyIat+Vb
+wPjsuP9r/UpRVz+pzp08kLYEdb8uLShhaeIn0F3RJN3Olt+xS8q05n1kWrjWQaD
VFegkSre2FptgN3q+4mvxbSP2RjIVnbqvEUQbpIUoC8F09Jz5LpA70HY/1VEGz1a
NAMjRV45VLgSzR2t9zaWu6rPexRGaQ/tuic32exXh+v9HwTsm5SmtLNBJp1NCxso
fO/Hm5dz9sEMswubwad6bFtMRxwp1Wxg36IBhTb2t45WDjf85eBV7JpITa5R/eMb
YyGLA4IifGzc1HgGWxxH6HVzm5xHcdA37oGYyzWyQP2WGcv9ch5CYol6JvqK279z
xYq0uM9DVwniJr4r59fH5mAOc3yd2hPCRmiSvkjLfpGia62QZdXibLtcU//Cv2OF
Lx2VKoc1pIJD7g8Wi45jomAGvNWag4C0LcWhIf5bcFp/6USfgg26pv+LYQ65/DXX
GaNAuMLhxfOHjs0VDC14qhrTHbQYrKcdG5/gODEfTsGE071LzZpPrqLeClVvhDtL
tomrXDShkzFEJPNmCE5N0BTQBFZ8dqaLW0ZcoUSoJdj3JxKQs2bhmuffj8PCBdJi
GNCt3IZ1zqyvwUJLN9qewdOK/4teoVogKqz1ZxKcoMmbgZVUf0VwJ9lpeauGralf
EppLBPQ2eYy8z8nqw4xLDk8pTaloEkNYV1mjoYWYUjJJZdH63+o/mmFbkDiJ1xID
JKLlQuM+PU1FU5o4ETtYaU9j247Y6VwZfsT/MgeH0ftXSqyu85czqL+40SBlQo3L
Zn0VU35end8E+OGyAajw4a6bIzwCmckC25a7C/F01mw34/QuiYfQi89GJHj9mF9w
wepwk8TBbSLZVZan5jzYY/JBuwMw1/7mCqt+Bv5pmiX8P6IGyPO5AabpCEdxXE56
Bh06mwMHO45utTh2Ac8/OxR57do+bdw4FUXKKalVVUE1LyAlIwMENRdQENcK5IqT
14q52ll6/8toKINr8vcDTbqZBxMvvxum6ZqkMQu8B0Ep449EBcSQXCsNeQPK55rT
UjznXl6CY+63CfWVeYoThoqzcRt3OL9drGuKU+KjNgbfNKH0yBQfqFDLQs2D5Vr7
KsRXa8gYyGcfYOJ1O1K+OcknYYL55O7lrF3uhm85WtnLoK/hffsHwSg48XPZ+WPT
UM1jtEPc4WWQspRJXPG+VKok33rrNTXNXsposlFnrJgfK24IQgMe9g1lHSopK/ZF
dY1LDu18kfi6P9gEDvOY2FZtzEc1BEoppP8QQcFaSwhIWmjfxW+IPGNF/41ACdUW
w7PsNbg9qVP9r49DZKhObA+SkklA779VNFKo2RVAee6wqE/OLcNAnAN2oa/7uPcN
g+qo0ZucZb48sIhsHZt7+mW9TyNGXUiZkeKAZ22ytkwgSSxartHgWfWFY0Gisbl8
B/nXAxAQkvMG1YGv0KyujRhGuDsNpIPs4vXE4Jzv3Jz9yphxf9B840pfX3uEy5Sz
/2cAfoQQ6TgvHi1JZAw2lVA6hQ5xJbM6RealYLg5QpNSknK+St1FePYLSi1IyReN
yjyNslOIeBOTeMyqKEXkzTet+38pFHw9141Fgkrto+xQhA1JEUyRtQvBRVtxx+gY
pVwuvOljGiqpRsfeCzbh7c5dppc8x1+j4tMeP5/f26f4TEPao+cbzDKGWHf4T3Pw
bUIb7EM1ICwypKhivrSV3zIheFNm49+kHAdyoOtPQdsjQ4bJGovbCGzhz8bRnJsJ
EnEryt3JsViC6q9jOUSsTthTrOfYadN3VIfjrUNiFDOuGxHqlXsFsaGT9Y8mbvXS
KpDPv/SL8pmUaFOzRk05mcxjU2EnD/6QVhWTzG7+sRIhr3OEpOzItJBUxexvpvJK
mztusfJeJMh0tnnodDuhbfMjfn6ZU9qkI23jme6ATdfFFjmAlgM4BvJgIA19qVCs
zMUIx0cep2c4Y7WeUSSD8t+GvyJldniBqJ43mK+IKJVTPGqy0D+mVOlkFidwIwo9
XUBFYPKkf8bCU9tqILAqU0v50DCiGD+2oHdk8PYIDxbQtLuX510rxR2mjw2leYLu
PArsSDwqtYVfLYEiTb2FbWzZBkPkFOH4M9HOn2Lhbl5+Ca0xQIkgBOd92NIDNf5D
Eoer324gDlZVNNe6SLRh3A/0zC2JVOdaKHgbE9Hmq02Gv5D/MW80mcxZBEjOR4TH
aXSSyh08DJLOIQbQeRUDMHxkPx2LMe/QTOr1LE020gifvbWSjW0G+hj+tbiT8DKo
mxjXjCGIQ0UuhkdYVYUr3bP8zxT/rMF1OaDwi3zPm4x3AQEfrV8ncwmYh6XKkgWd
abZqBSkAsNQAAzL66wpo+jX3n/GPKTNK6hPJeyjS1tpmbA3Pjp3Uyto4KWQUD+8z
bttJKTOlIPEOv9IJUvkZlf2xnarzAQjlwAqfSqEf6GhyW0mikMl2Xml0HSFG5sHv
Djl+cVVT294FIJ1EWV8oBit5eGM/x716y6x2bk8FMnMl/JognbXKEFswxmWDNvxX
kpPsL23afZMCxN0WxLp9660i9g34zYUNtT0xh6dP1sC6pSoYvxB/xFUrTzq+JM8V
gBb05u3O2PylGZhtyNtWxdxa9X1Ee2aqzx/nRrQb1Xxv/Nl+9qdiVyQygAaoPnJl
Z6LIZd/l1HO2o6nCjdTvycfOfDPhjrYxB378PIEwHk3aIHf7BnAekPnQJ0EZNxj4
KSMdk1ZtoiA+GktdnnH/m5X6O92UeCpMhv5mjP0OJrgIgBFU8/P0U9ziwPht3DKY
w0sgYlHrVw2++fjaZ5Rn8NBFWFXHT25AiJymAkS06CUVGxy0tiMTT4kP4oFohMXI
iLzIh/ExStQ+9vh0y2wxFJxoDJeZ+eF8ugCPjrN2w9AjXcH3Lhn8MAWKb8YUb7/D
wuuEPFhseVTXzlZZh1hgkVb/BrmrPd0tQJfE78Cpam82nIT6ksHGpRDxbrhh0nT0
YiXyGfvw5swx+qODJpl5Ty2WNhrmp9IpCeXHH90Nvn13sJ6pwgx50YdVMSAC+qs1
8L018Z+a36VNOoDEKLjCFSveXqamGyUCMod2cCDlbXNHDS4CziOk8cvzXDtWqe39
6X0I6vcYEoyI2vNYYs2o9iSI6WBYNlhbYcBUmAzleLClMJghfFVCDDMcbVffISGr
uz/DS1gZEren3JUPzyfTU++xv1n7m+vt3mfWNekX4Ff4+nBq7pRV+SSF+lE9Y5iV
uaDXZD+Ye7nXM/O1XSdiT85Kpz8AwCS0fq67U4+0zZOtgQRcZF0T/uuVa5Y4x6zh
KkSps5/gTAtOZX0EbxEnP1GU6uS+DlUCgO08+3WjAzlSSXtxJWt2aWaOixMvt7zH
cYY0ikcwfLlyPoP4TAH4bfefUWBEWzyUtDwj0IXFH8/dF2bLM5zh2OrGb87dQq0/
zPmJnHm1iAqVMRbHOUwGddi381R0mJEAa0pgYhU/UJzoa+fj+qJYCfYawafoljFu
cxjMbgMzUYNNPQYRWg9AFMbCVA2aUa3KzHKm1y3DJpICkTOq7tZAQ4GO+B6WzB4s
4VxAUTz4lmP0/fnepqmKF/aszCnkeF7tJnxazJ/ZIlR77uJ0droukEjpP5U7X2P0
NOVYUB/VUi1V1qHKghQInC2zYBpQGBJJiCeloJGOzQKsDCbuVBazQN58T7YfORbS
M5CC8Fk7xqO0Pv9LGkBBLrduD+1iCQdbwxa0Dn23tr0K0bwjirs1lrEn2TUsgw2q
CPctJdDAYVu2Zk4IaPkbYbafzaWXPR8/n9c+wHvRZ4mnIP6w8ldRTHVvrGbyFT9x
6zthMeer5/2pwsaF3oCL2Q+pVlIYb0RhGbdYnhzsdsdvEOlLjfeQ86YD38MyfGE1
hgakV4iDEFVXe1Leu9D/cD5Wi5miLjQBQAILub5LNboKvAktke5CcfBZH9+zaHU7
2qD1yh138WXDJ9vhAEagBuqaHYB0105/pPzbngNWtxRvR95AK2G50dj37894RCyP
Ve5IIidG1703nhUQ5502ygt83OtF2gPkRDe0B1yDrPS69v1GWuNn3iiTEXoOoaOz
S4i6+A4xjb5KWKITu3HAyKuWxSad349Bz6t0i9rMpMGRM7iyj406aW2oTFWvlaQx
v/Oslfxu5QvkmvxDTu0pkcfWWJoS0910QFJKKltcTZwXmlWu/R+kAtSfijqEnVqq
BaKM+KfwvNC6Qxy9wuW3O4/szqi1m9p2MEed306sh0GXhxLUBv/3lJzLxWOzVah7
exG9knj170C/GO/ZXcEHCs0BEI6udyIIjQymWCFjeSliiUxgzSCw5OKC0HbQLjIR
wM8nW5rumAV+ksGYMXbIyE8xexK1ZSvhxevkahifAqgV0LZEtHca8YLPb5IfP27u
kg2OSyLQVZcxiIbldCR9UBAILXc6A6RkaWWUZayBAcJyZJeVBzBw964r1hcF/BBx
0ETFBdVlWhqfhBkTSb4AaHAeH3CsgwLfx+brDjFyBB2NSh/86a+H5jjxQgxZHERK
fcn6np9Eq0Hvreklbzlj9iWB1qUaJhON3a24IAH05vb/dwXlzMg8Exy6lGl5ZvCX
jUEVjhMcVAo5P+FYcGbU8TBXAbXXkHSKmYmOdfR3xxS+GbG8pVG7cVUFdbKaB5ir
NAaZTvweySccf46gON6NHz6zBBQX9DKDVpaxLsxTSV9Uob4fGa01/GDskhAzBe+W
uSXISAQK17knLh2JpSEho8XgUQ6zUVMMBOCcKTqU+L96TEFHd1ALtdaZLyWAVipr
HhIb5M8dksGA2hNzvjDGodZOZnlg0tmWWJ5DlHmXhegEaxwb4+aU0cDQDLYrJgax
ImXu9+qqTal6plZemPqVMk98SnpP0gkoEohIY2vh47a6pj6FXdrFDOnjR/eRvcBs
s+A0JYSfY+m5GRMi9ofeuha3Jekc6V1Vg7f9XqZpi+Swhp3xwkclLZQFM8aN5lh2
qF/0EvkoEUP79pjzaEdYhdTYKUzt1Mi5Xefbmo+D4/qFamhNa2JFGK4Jc6ETaxC9
HZC9Qa858qlVX6lrn28dZStRnysQzMyH5U9vJxB85tqwZszxkXAiZIYIoOGYprEX
I7GHzVp1Jy9kl1eXCm9Zb9kBZU5ZB6Ae8L8nepvZp2LN5yhC6SQkEml2XBPQfwZp
+glydbLo6wvyS8VyLV53Wi6OF6Yyt6juaHidKE04eAkOPqe59FGrNzGXfddIEZOX
GbCo6B5nLohwUyNUp2mPEvbPtTXTLMmV6RL9ILXACjkKKBgKzfDqeZVUPX7MNOys
+jU1b7oDIuJcR1KuUDg7BFXXGH/dnW+T7+M+38iA0DTQosfUo1df+C72UyexvkD3
5MkrwayS6UCRNcTP98PHIk6pexAG5KkY2pGYanTT3v8dVbACxP4y8zC/wmv0KZ1y
WtSuJnzuzcYjCsVCTZ6vLYRm3IqcgJlF001Rssd4YOxmhKeFeakQIIhfl5vE+hyp
4vmip8EgO4pWeLD5YTqVVPcS9/9c2TN7spy6G1iQ1gciLuzsYyI4+En/0wiD7sy0
359rH8Qi5xzbM2rfXmfD19fPKAYyxR77t0s1nudvAhC9jjNz2QurPeClzByjQYD8
mkXytiv46CmgeR5zwgv8KJI+8tkKi5So5BczGg6NkMp1jHBimS+/WYVcushUxISU
I9G39kmQsGbHjrgcAKvD+yXuXyIpzCIvDIA3i7w0i6DA3M1KKHpKGWk9ADgLpmHi
7ud24hB3XWq/zume/SRRafpQLLOhCWlIMFJpuOQneHSIMvP885Np1bOV6x7zIvzF
WmUpB1ZIz7uA+1WUVymvrEXTSkK1kBDmIPUKIxTAhEmcN2GHLHAjDclnSjnvt/L5
v0UP7F/cooqPLxTfnId4+PIlW34QD/z+NqMo6X6zOfqSfBHXubU5pDC9t6kjFnaQ
HrCDhL6RDVM/VmBq1f6lXt7TqNg+6cE9niEgFg/pXbpqRFnjdzl9fa1IG/S5jdU/
8adL/8djifCZ6bKtNC+ZXNOCyt77uhQwk6T6RHQ/gnJWUh1siEukMVx0pDeEw0+A
yxoBmUCSIMsqmobfHlGEePhXO+vbfCQ2EotqGPOlJ8pOJEFMLSU41xbKXOPiqYnB
ewFJLI6dvu9psbLE8xOkzCM9l8ilCKapg5HgOlC8jM23XQniYi4Nda8WkLDXjn/c
zufogVxz2vgr4WHVksYYbYqw84ZdsDjf9zQsqnhSHFFCxiF0K3ci9mm/xF6xmUjQ
dx0HsU4pd89eLb5R9MDNCO5OIn3M4MIq0dkydHZePO5E+JYO98PHIlX1TmzxWFjK
S86ATixlUux1pR/nZ/bCWC47T50E+Ngiw1Yfx1PT9a5n3zOrHbv+mFwVvJjPbEz+
YDCFQGf0ZwxSN+huIdFdJ/J6Erjki3ol5+imZvg411wfUEzMjFfjqrIJ3Poo8Fdw
hOGsnOnRcI1SL2wz704old2zjmYYVNJKMuuVBJ28RNIZYr2qMC5HDk3EeKlb9K6X
O3z+dhJBA/mx64dtP9n3HEg38XlTnlH5PNW9Km+6JaqSe9tPm8rb10+CZit3MT+A
6RPqGDfbyfRkhTlqdpJ+Hvr98Z+VbhSafCzQj6+6e3+BXE1RFGXAyuHb5H1FEoA+
`protect END_PROTECTED
