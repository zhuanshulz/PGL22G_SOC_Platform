`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jgLw7kNToK8W7QAyQZEsZe17f1AcUusjKyggUFubCSg1w+NA2MY4ZQcV+CFiy/v/
PNIiBtew/zeHVRdA42AOD+bC2+wY1Dny3yOeSgFOVj7bPT+A++ohMKNQVmyM8mWh
EU3cCC0jO02ZvPBxPTjI7GUxP9RezYBc3I/ARAOAmsjg8ZBAfZu1wCaGMl76T5du
PpKxizQvKpjor1HM4maoEHgIrVFzP34FbiVdFglEXZJ+vH4fsvzPB9xCQfmeBrsv
Uw3GnHtUiS4GKt1J4w4qRg==
`protect END_PROTECTED
