`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1VIfQrg8vuz/k4nqgItW8GeCeE7sOAYvRJ2NBnqmW+J8LV9xZThWjHScEYRyBPec
Qsugiq4Wy4zuOroQtEpRs1QS9z2gH1aueTClDtgU/zTqwik56cWn5A14lDOVNH9D
uND7mnGlTmoFQnzCobORVU3UugHKpKHK7XHgLMQJxg000zIxiX9rp3I5c5ml7bwE
wfCLYMmG3bEkk7P1ZugojMiwsXAzxGHedzn2ktzsL6HppZc2WMd5j+vHZ5jrKZMp
BGpxjxBOS351Ws/9ZFfWxfwwHZpmWs6jQY1aZIpiQZyBcEkKiAfAiS1T19jUxmVN
yIkJmOMz+3Kzvosn9vEGdF/qZbISc+uN3lCm48bHnt/rKgeLRnobAeEnJbY3/A59
PE59TzhgpD4FWaey4iDVZu8eNll9R6nTeRTY8AMwa878SYrWZ+BlHlSLGMRoyNSo
l4aOe8yWQ0Jx2BVE1cpQorBrZ6TVXIJV6PvG4bKqXBHjr0ahuC5kBRC6XjE7+ZMm
AaUbiFPzSndUKEzgUrQXxKQRGR3wK12gKeDk6MZ69tc=
`protect END_PROTECTED
