`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cFPiXDgwKy+w/Mw2d4nHKeBEivU3W4Il94Q/rnTu7TAvS3+2ISznnV0x2sO+wnlX
MozzZ/ReY0wKALrHTrDzcw4hmUGHgdf9maKj6gvJk/kwVN4JrxUsyfZZtvvMAMoT
WGmY6VnBuEE7fPs7Yel8GsO0YHMcQ4fWXQ3bO34SAzyRSP551R8y92SEAx7t1EwB
IA2u7owvVBB9CpnxaIJO7Pad7fX6Wq/Nx6y0HyweW2a0fgQDRmqO1T9YepOUGs6/
5CQAu+odGV5AiaxkwbS3I/O2Tzt9lmDGjVramBpQNsup9+UHEnoox0prSUK/Shft
qyv41i8q/eXsDPrE+Xr8rsyocxPsnMUX9lGhOhZTCvYGFKWKgpC6mcYy1lEoj6Ph
zSg/GUWQy04mK68SY8qRzanhgrLwK500/vumbCl2BPojOzY+I1yB5Z9grGmGjLZZ
`protect END_PROTECTED
