`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tx0TeZdOXqxS8Sd6qRQFtW0gGp+QTs4ylL4oCkbKcnIH0FS/I6z6Fsrm7+1eX3if
w3m39KK38aYfJDliu4YxTQtUj9t7pYtAkc+Wf5PX5Ya9EVxvDQB9hLwgFdjNOsij
JWX/O1jeCcW8mG3qwmQr0o3e8/hw/A50ze1XGPF2vNU12jGEfTDwYj8YMT46hy9C
2q17gDXlPysK1GaECALApxc3yp+xHY/SsV3wxMQ/D4bq3VaM7bgOZa5Kzec+Lryf
tkrZHdkDTdU0bzHbBCd8ASqhPPSNg6Tlf3NRMVDCEfDxZbHL0FsO/v6aPF8B8KYP
RvFtC7upQbnI3uQfT0WImjQMtrlUAf7FxJV/kJFPPAi9GA6jwt/7T+HFS28Fg6G3
/Fdg2CuWuutDo+uc/psoj9y186GvB26gqoWYeCk+d1MZPwrQs9MzOHOh4KtIu8Xp
JDlE1HzBdRcJhkZh5EbGl/9MEm+MkafoxAvd1UwwrUYXYXz/BtMMVf1E/BzRiXac
5TafKBpfZILUrQTTplNsR22f4z4Gq3u+oBquEY7uoNjR+IG8n7ZgddLa+LQp4gUq
HouNW4+UG0msTdxmTnFdQiNHQIBE9WiA4t7V+Pr2mhnfnYLs4WhMwgxdL9uL2UmX
K8jS2JiElEDkTZQvo+svADB1ID1OscHuBFfX8chLlvp6c2s6L9dhy3LKgPNfwFt9
dXiiEO/x/hTSn06hOAkJOe+1Hig7Aaflw68iAodVfEmsE5h1WAaSdfC22vi2uxvU
yCbTozCmoZ2UesAfcrCX2xcsAbQ2dAN8xwJhwPVNAqMdJ66vCobeOTSJNc5Kf3uM
`protect END_PROTECTED
