`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qjQBN+CnJlYQR2G5NipB/6kykffo4HsehGrEFcIRv3g+Gz2G0Eu/K9O5a8byH8FN
TN9+bXxaNZOXcB8x2bA7o3NZ5bVfigZ5r9T06L6rDfRTFTYenjfF1KZwPirHULVZ
xZAb/STkaSpxSlTR7vACLnglg/NXF6Hx9A/Y1xTsSc+ebCHdTsDCb7zunsNkaemi
0EuHoDwbBqL9qLdijqGr+9wZPG20Z6ijxm9dvSLgbvCylrkf9ncWpzmbG8Np0B2k
4UVxFZSplKUagNS3kYuR1dUkDwVSQEtxaZN8/lNetk4g5jy02lixVlDo32PSVKhm
RBy8SyfV6EAH2ghkLnc7WONFzbq6jdiV4KflWXyeh7JnHcemp2NZs0Sv9SBXVl0+
2v18sgrDfNMsqgKC+HXHg+uS4N3SyJa9n27TqkPkvdXW0ltvXX7c9ZrKTn8Jof0h
0zt2fz3V8lwBj4nFo43pJgiPL2QJ0oNyyFBjn1N2yYKPssTAXeXSfEzkeTyMu4hp
FgH1V4PTlPozSX41ZTlFyrT+ON8JODvAmXylxG+d2WAaJmP/jVhA6oNKXUtoNtOw
Atc8KIdKcRAciz/3TBgCqrfSxWFTPSITMQ/WK3y2f+OvPQGawQ3eGy2QZjAFM1wr
7tyFCwtvsBf9fJKAQDOXX7nHUNIyLwRR3U+fdCWI8FBhLjBYsI7hZgRODsQX0uv3
aZbWgs3OApq6MfMuVSaS3d6/87iH9EunRRSi5rRtYUDUbH5dMt9R/tPRyhUKvAP6
X/QHj7YjTwGo1I7t3P/on3bBAHpCFNXBnYEKB2tQINYp8rJp0mf8Tg2GultghyVA
abmzxSrPe7CeeZED//5EXbDOi4qME/J/nLuJyKfcgcapmQ9rLhiV+MqYIxAqQx3F
uHkARI/wayr0pe7w3UxUjxB/cabJAtcSiP2hhtwWteetRztyA8Ebn7d0Mj10I3DA
m7eZ0cxLUCA8lLLt0noeubk8g9S7ZF+ZDCV96IZtWqw=
`protect END_PROTECTED
