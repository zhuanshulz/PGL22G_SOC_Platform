`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
REVigoRNSRAQkTi1s4YdCOxRG2jgh2gxefnxRclvXtHe0Replhox9p/zlx5wtcqU
NUCu352ahiD3c8BQFzGfyh1NbLTeJvOVhDKueJ7snC2mrgl4rM6b+eV9l8DhXl6V
F0kvHdnuKRF2PVr25K8Me2caJGF4Fw6mwZr3fGw4ELmdQxuuAeM/NBIKBUHBRqvP
k8fLrQqwCM/YISHbt4dJQHX5gTNdFsqzdD7C+bQ7DDXQm4gvQ8HRZPyRlFcIuQTL
6AoqvrI3KkqlZb2piTHf51c8VppesILRQouy/Sd1ekxGlZyIQZVHJ1eK9m3zzq0X
jWNCxWZZlWyuxaM8W9LedRX/vFs4hS6uTH12aEoZQDbJqgbq24Tqra5sR4iLzEzU
AGe5kD0glNm5FtbcT00Qc2cgIM+wE4uj7FAIdDO8UCx9be0mqlks8QjzaYR5gg3w
HLwSe4w2yegF6EwMHB6xT9oSm+yK+bC6OvkF0Jky/QDq17OtoWv1TeAEiDcJikc6
him4PU3kvqSmNhABCRdMb4uqd461wGxZ9mqBmeWtmpUE93k2xbeZDLB5Kbqady7z
6Y+uWYI/LjoS6iWV0bgz8ntkdY3+WLxYl9EkWjgBNbdO1r4W567cH25YaQHRsQAi
32mtIaOcXF59ihV++xUCrYhddqY6eALW/WO8DZzgPGCnTwNOtf+v2I0nRMimUQo9
fld/7kTwR58MsDnKaW+yS/Sq7PMAFNAIJCZjY7pZIXDTrY4jmeguPEUUx8h2/wHX
dfSBgq7KtQ32B/2x4Me3gDCBWvlvQft9wkHtQ6Ah7GLbU9Qwb8l+H6TXqNAf+am4
mNSdRU8NowdRdu//uV53j08Pjg2YzDmUh/t/HNPUn6YWDTVCuPsbyF7jpr0c4UCl
ZgqjHsfXHJknOb6z1ko2Dt/JUDEq9yModTkv2OiumDRwGBnjnzzX/ZuMrQmJOsbM
pvy32ocYToEQLyDuQZ2Ey3d+6cc41KF8iffo73nVHlKfHx0BgEwA/0/zQzp0lFve
gyAUCrzEcYa1SLoCqKJhySbYfitjli1ow5q4bbtTjf14VHPUJZTS5KGO7pTqBXXQ
h+LePrXENxWaqPDa6r7TTu198c1GR1YfatcAlNJ24kKYN1cseI18wugF7tN108oa
WNg5tQW+42gQ9ZsoYgRg2G5Q9TJKTo8yM6AWoNyhysVfRpYqiO4AoRzVV1AA61Qe
KhC1NOG56iMlJsEWCtC50w==
`protect END_PROTECTED
