`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YRgfmPtsBLKz6ZWRjJg4/7x35oOBFqwwTt0vgFB5VSk7DSqG+XVoEUobafwB2889
4rsdF6BLRN8GVMI2ADGWt24ZT4EfwFlltqQFZ2ydsklcSVxqPWqe7fHBHx5q+EK1
1tMNBBft355DqSK/Rjm44xrjtKktoAQGEWk8Rxt6WSNOGful7FdZCAsNYLoJxn8J
DLM3+0ToptTrmrxg+NeAY4vLNvozUNyRLgfTwJKDXQuAX4Z4MxntcOfFtUJ08SRy
T4ZlTGBtkAMO+bcaL0iN8YskqmWZWSwUE/iCxzKWVQlaGwOd3faTnd3EijIKN6z0
7gjMrLN4O2xw/0okj97zp5ayhwOyM4TqCGYEOo7cwwlRwFov7rTDwFX7jXCJRNXe
3ocjgVDzughkJ7qcjwXqQA97xDpgs493zAQuL+lfo+9i2zTC9Qkk1Cp1E+Ykkfdt
2BcGZwxRXUxu21DOqZ1wcgz0VDYyhPtDZ986213X21Zi4XkYq0lZGhflf4Alm5qB
L73M/lX+IKtg4O5AsK9f1X/ExFq7rVYr4wXUs0ntffYDXV9gD+9qI1idGhVKX2lV
oMkgpjr9jd3/Ne2XxNF2+g66YDv/6RLkaWoRrQmy3DhDVeadX9N8OQmxuOuP2x/W
9wOqOqHEz7WPJrPiw4xCiByuMYtPbzAkPCgOG5eztwkDyEujxXtzLWN/u5Z75is9
TgN/5riaIbzpUKYyNvOgIUlcmWUo+YOw87OqiSXxBzwwEN/G4u3F80KLxN6i5udh
ztBeOu84YYHR0raNi+Q2SjPexWYgVImhqVJhu2n2m0VdMJ+7BlUex6XRguVHmK/N
/ImVkwTpBdOgN+Nc/ognhkuLTvzFHTyEnvoYmDljkcSA1QzkGUZXZeJEbel8dzcb
nzIikEuCbxqgXPffqRmNHmXW6HGwXq2bVT4wdjIS/b2wcah6y41/XyNl/2gw5H3x
x8Kt5VMVkl+KwJ1xIrysOAuCNJumFkvnEXeg819NMHHB23o0QgFRj/U7KMUWw1nF
E6DczjMTC4P7z/BtSZNO9eLB26Gu9TgEDlGavY9WNJxeBazLtlSgQsza0yxiAlXb
aeMvZD2/pSEGry/3YtvtuU+WMMZRnCG3mANRaj4uhJZ3w5u+waSy9KYLHQ0ihN1T
l95JgJmeKLBb5TXHjqGB3u2B7viQAatbP3NmQ/otyNLv6c2v7YWl9fqlla89Ozpi
eJ4n+ZZlRetEjLXDi6+IlNI1rQ1gZjnV5exLuJ4PQJmeSqPkxPqaQVWTAUTb2isw
EGlRe/5089tR3DQQj05aZCaJa6jaWTN/Ic3ntkt7s0V0YgAoCh01YPRXwi1w2P36
KyCRnsWFf4gulhILOnKtVzIZ4WbfRsLAh+ovbBYyZXfsnUVu+V2lJuNdMEr59Qjv
l8/yZ8J7lq6jNuWc81jenl7mMpYnP98SIQXXv/GkS6xpqdAOVSyeXmK9TJ1H96Su
7qHTPQ+pZIGxOaChI6pfqCnyAFxY+NY8M4B5y1+O2xsKFrBxlg8+y7yf9ywDtlNJ
vBqebZxtqRDnCi9PtajmKqQ2SleRLYiBVh+BP6jdvsJBM0FVrG73C9ie3yCx02/R
unPS3dOiGpthMH+iV3xtzQLMMQG6/3QLsgSgNv4za43b5lF9NEn2QU24NMjC8jcU
LZpSHSZ68H0JsdCaJD7QtiqYe1F5iwViu9cxz5Hz6mJgIPk1xUHnAmzqZITGjKNc
Naq0sE+e7pGHJ+bbQrxhXVrYKawkf0VufxfAFtinp6xIFEbsPHE9nYkZswtHbp2R
uJcxljJ7jXpNAPPXxyMDqU+oQR2rTkK8DS5i3OdDflCXN1BJxikZdpjIVb9cDA48
41d9v69nia0J4BUJ2R2prmIMXgCZwW4mcemZwwM5i6Su49dfTWjlTpQ0rCGK6UFf
XBpus0YkN1EfPWusZjnF8O064YJr52J5FRp47L3HGhVhDpu60VDlLVJcQPPm9lbL
4LU88Uqr4kHTrx1e3g+Rt2iNDLzPsQtFVE+ZMX81ppL9IhmkSUAmkroJz1+iohOJ
zbQKhifTYYTFuQYT5QbbxKVhp0m2XiUNEGO72YuF6GO//iknWIIhJ0UTxPNfzuVb
G5un25qxOOYBAo6w7pahFAEvPXHcGOGiPzbgwTsFTYV3WOEg2eJ51cQEtddZrpNX
It7VqrG0Kj6p7iu0IPxe5GzwuNJdnVrQMJrsGXC3/fQ6fDM7qANXeSv5o/iDkw75
iQ+FLMRqluMVntDyNlvvOamCfaUPW/a/j2jYLkgnusSL1HUJRl8eGm5Uzx5s4RYa
aPIFP7yFje2i7nw0aQHQgvNIRCWpM/a2I5Izqv6tTLtGS8ytBmUtD8FJFnl4QgzE
fM/k62BS3rQQ5VvpqDB9CkRdcmxT6FOZbcphv6iOfnESBTjFsUJGJsheH6MUUAxp
ncfeEPihKjm2X7KPyW7W5iCnCJgIicjagPwRrpR493YJ4tXz7ndGNcF97eCLhVgg
ROm8RrKS3QOhEW4loL/Jn/GiJ6FjcZQphc1862IP0i+ACXUK8yHHPWF6xpoPOigi
3r6u8gXegyheqDkCaZsDhw==
`protect END_PROTECTED
