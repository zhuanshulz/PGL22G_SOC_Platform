`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GxXbU9IZ4nO0xDNgo9j0FgzDqVtKaCVfG+IvzDoL1kk3mrTsXjttobjvfJYMUCZv
/+s6kinwWyNnhbLgBHDa8ouO/yYKVoJhRN5CbfLO0F3l77tbK3KM4gs9s2KU8QlC
UfUl4pVz4ipi8RQFri8gkdlRBrOVH7OYUlqVyjxd0QxCnNAgVpMt1CfMUoXqAe0v
jVjONEly5D+lAgGok/iP/yOgyEb8surdzDfThA0Qf4VX+M96WtVsaNcEmimGBpCB
SNxL+RrT7Wo5QReMkNwICGLGXOFgcHfRsYcx79Jq5sii4cUr0F9BxofRwmZh+9d+
X8xcVXOJ6Xev0lpm4IqsWLY4Y7UV1HkKVX1QnxJFVkxZn2q4bHyOs8ZgQs7z653C
nnKxgWW62EO7c+YDNPCN1rNTKnnCxb78OPc6phaHi1oI16zfi0OzTiZXJuf/d/2z
GpvaxlU0D6iMU2emwxK8r/S1F5ZSgd55crzJiB1D8qIwDZbYOZKPJjcfePGCFjJo
5w7lBpgbXbBjhXB+JZqhQGNzoLX1rWyf9kxXgWNH3k/jYUhZlWzIV+lyJn8W1Rz1
5LftfKtV2NlR8hhAzThg6UPygXjLy7qTNNenYlYDBG6V0USzvU3abZK+Q8lFnJN8
UUzZl3zWnX3Pze6qGqC+Gt5PulZBab+XwmU6EIjQLdwrBfkKWulAKW1+EhIJTIq2
NJb+RvIACqCB+MOqC2RcCWYfDVVvkZjEMJoYUiws7yf+d/7cf/Paf65enWEzBjTV
D0CQkUK/qJMbd6N/COoaPQ6Q+bGB8pf0auxsYOR3Y7X7h5HEHfYf60nKVekoX/UP
Z0h2McXafQjQnXipLGPQgmjbOVdgQ2cQUByd+GJE9NqFhtVem8Ud/AYmQ1IKTEuU
BJXnGfl+tNykgfy5bQIqsRMksPnuJ2FQPRNuFg/IqBLChPxKS4Hioxn/bR1tyQR+
7OaXTsAQDC813PM/hBRkwAaOnJLKDw6MkRm9y6NqboV6B6sm31xt7FNfCx7YwLsW
/5cQgNnleBYjNt4JTvVLsEck5Ncxmw8+aeEYJNeE9oyyxRkwqb7hN2wFfazSoulH
5Vk/LTmgLQOwxlm5EnC7R8f9RdypF3QosE9+dkJL9AwTjDNpvVUBohUtF/tQmCgs
h2I+tK7a6+b8uoZb26eJcCf7uID92C1Xuo7bMmsojOndsDpK5mK+Cb1wpj8po1eh
Mo89Qc79O1OuJOg7FhsZLNKV0DjOsQAk1/2HolPtg8phm3x8QQq61B3GWg3McpID
S3m6dHb/j8Boh2r+/7HiT1uxazYMF7CmeQXEIA1N8gecXKFO9sQF1F+G3lJkRoVe
lblQDlrqZAn6bNA7lsM+InawiSEPrdGIj+pP641t0rkAvoFhu2aWmsGoBEBYQ9fe
juGZks3yJQByl3fjUOj7H0UAiVaWQToDy6DvLu5PaxXVZz2B+aNlFr9qmKJvuw8P
wdlejaCs1kx4k4ObupW74jFOSSTXeh3YTiOhm8scK3hy7m5eINlkBojcii4KusZL
84PNuYA3JRDWsJopFj3VzI41NIWuJDjtJX3iuPWjaSvLCyXOA3PEwX3ztSPjXDm7
1G+tugmECmNCtYpU/ZaIhqTPuDmh1O1o+BhO3l9LGMOewT5kdjEBn+4F3oxPk9iX
S9jaim/2aoXP8UPka6foodZK2zRRPTBi42jtKu6dU290qArw7TubjFSDQPLQ9qN3
vbib/wZMxupe8JXiP629LSXAicUK2WTYpn/YNLhDBPY105l7+CPxC+s4k0SSlCkk
Xku5jGvZpGUaRglf/7flbwXPkBOeBrjFPQhaz0iZ/L6WmgdUWFFL4YxUl4lUeV9G
YRbIfYk8YdZ3ICkhCBFcDNkSYlFw7POM1sanaVkhSugAylqoC+Kvt3HgkBv7ouPM
kfAR8RATgOzBdM50S6FPnOKbNLiRavmTR0X7ycaZ+TRE3iDgaV87hioY7oSIWUOv
`protect END_PROTECTED
