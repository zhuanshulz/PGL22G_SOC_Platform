`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xBeOrPnrNwf/KkNhc/QO7NdSbQPWGEli5C2hmbqLTYzico0iIHrFzGIuwv5z7vVD
CKegidEDpSIFsTadEjYk7GEvNSGIVexJp6VdwV25DXLJMg4md4k9wFjH9O7Qtp3I
cabQz3FVrJWEDlTbtOehQmrKf/OHolg51PCYp6KeUy/sk/w79xbTvaboxAjqsUT1
gQ8rSshnPqmMhFKgINSiVg9dfxK3Ow4dsfrJApIG2r5+4uUiWNF3l3nYKhK7hYuU
zckcsJO17fAUa+dBDPnUPQggFCXC0HeXwWWAMA5ZXrDPSoeZxKNnjJpFSD9xnzkp
bdojtd0+mmqNhEbuFuq/4mAI/1Abv7r15VFVDtrILftyPEXVmRrc/C3awUjo4fMq
x9ObvpmQcDU0S+4x/nzxYm5CD+1PZfNOda0vs+SA4ecmQMf0eCvxtn3BYGWJINUC
KRmdweSYwqwGmWvFD2dvi4IJ+YcfiU3GRG04q+wmfV/wg7btyyw4fTGFNcX//WW3
luaewa5bTmcqMp0Ao4uD3yei6HDa5oxSccxqEjw7vvlxE5g4mVLCgfEZ7ceKw1kK
JB92hyRjr1ZmMwSprAuT1s3HLcdIEr/xS6oqhBfgV7Kl+1EGl1xhTH+63Tq/kVBZ
zvYcbSqg2ujNq7lO9T108iE+Myl39AwTbuIRdcKxblZpj8OZXIJEdWvHY/rFD/sA
51wtIbw30ls6sFP5tjGYudZeQqPrDeN/IaFcz9qmJEsjeKkZ4sEqsCO53BtpDpcQ
IVkpogOd4DEaql7zRtgi/+gZpQglT5qOXEQidBn3k91EpWodBOyp52SKw/N9Zui9
zIdzDEADbSoNor43HYAd/OTaaj/aY3nidYYf1rMt1dGBv8Ul3NVKJowOpalBv6SA
X1IapTzjvKtWu7bcbQc24xLs0GUZErprg0MDMcv7OCMbe4wBQcQVq8e/4dmU3inA
TUn/5ZFY0cFgci0Xn0l5lT0DbZTTv5dWI7VASKbqDrXUQiS8CJ5qIeYwCfK2i/JQ
V//oZyV8/QXeNcOhW1VtglxSwSyCCcLCW+C7aUeQ6v/YSjGdEqIvJPt2Ze7eeOjW
KgjSGloKPOGuuwBKXtQIO+u8+B4quFnUAiDp05IIXAIYezIUFcqA+qZaNOb/W6gf
/946hzKtLdVyI+0zkqAmzQ+cEjgbj9cBmj/ouVivFem/0JUqZPpa6s+MkSAdKPmF
anYD4+Xgn/R7JsOg41jHDjxec2V/YUpujXuY0wbU8yOKzgX++QIaAuL9IP7BvqwP
Da7Jqxz1iNFfWtTK9vyVhUdFuvTbsiTAIxUHVBj3EahJwaJEg3RKulmv4eEWj+h0
VL8S4oxJSito0YqxbGLoGR0Ca+/2cp2ODuKFminSBetcUErZnRFpbRoaN2uxjhI2
kbHDO17WCObV53y5eQ7TU3hQE4C5t6RefId75PQJu5ivCWH5C+QU+eSM+imlnjh0
vLaC9uy6wLzf/T+Uctkqwj5WKcqYIReDXs4TvSb794MKWgWbeln0lvvVN6ua3i6Z
NjXJj0YM68mB6eA6HoM5kHCSFUDNgTgeJZaRGJ1EqxFRxi5PJbLIeUFMrEh2u+Ve
FKsmhMkK0JOa8VIzG2SQpv4swaMUeuxfKeUhpgr6FPGOTy9GWl0TcIewa4kXHvgj
XywCiv/ezliow/ty+WVsdPBU1Iil7sYKJ1jl79HmuN6FoHukkJ7hBvUsHOks3cMc
VFS8+mUXfOLmRNHlx8u/4zclO6pqcfCXnFIwvkVyDlPPPBkVw6Kn6KvF1EGAkj2n
BFTKmLrDAyrK4ZVPKQeiDmdXHqucO5TdTbliljFaZQpbdCj1jpWCDHWr0Wpchfab
QUhP8qTWBv+gNiet5oeLlMJm6RKPiqRJBjaZXscgbrci/yqjk1nayDjcNkcrZSLn
Z+FaefCGC5dmlkSzcsbqyW1lNJfXPrlsDQyKk/7byuJgipMZheO0VoobMU+EmcYY
QZ75xGWd2tnaoUjhZ+xmvhmIxI8hS1lnIP2Gw4b5AyyGVUGsy0cSS2eH0dSMho0N
TiPtzEAVvW+VGnZXfiwts1xg1dOKlkrn2GRq809d9Rn6b4flhrzLLHj9+Qg54TOz
Qs+4unP114r+M8m7oRTAiqvUiRM4qGTlklcw0VIU26H/kafX16Xxx00rz9Q9d8nH
SSda8Hx8yRaLdk1B7GFTgMeHmRwdafVAftdb2J+XXYLscRbEmR7BOFdRrOKE+ChR
DP5kppSr5tkR/wZ7l4Vvyx35GqLTVOkhSvVSrzlVJT/m8SwJT1MBrx5SC3aWKuGE
A4ohiOaZyLhG1+FLVjQ5bkBBAYL41pFSD62vOxy3iO15AxBUfGm/p8CJAePpNKk2
0GhDYXE5/uJYOHDdcyQF9Trsfa1wVsxpyiUfuAGAi6WHL7BU6YnjD7HJY/RKzlLl
zWPAV6y/Vn3hgsor0/h1pSmf0pioHod+++Jx0Nd3ZErRWf5WZiC5nddP/K1r/0Jy
IFptT3yxbG5bMMeiKeE3SSpfQbLazQJOT6SdDRuBth+B9p2Boi6QIICDl+3ckxD2
fVhv7sPE9R/1Vd53Jjw22aFFjJ1rCobsNRqZXXGMSod90s+Fz07Oq5sXGWgyUIzs
jsUQVBtE2tPEvSuubi+c8IeWH8lgmNfo5dsZnkD+nOfr6hF7xOCdLd1B/RiXl24Z
hQRGLs64owj8HNefnGJiG0TK+pESCh61GqqhBcNM+k+C75XDJmc5iRzFBMgGeh7+
ItKNcJHOCg3Tvk4jVFqIvqVJiql29c5NZJqSEY6PihJoZ5R1DE+caGhPIsZ2t1gB
ZfIAu+9OryTM0TCDq00zi3REqubHbe0c8LG0UrMcA6WhCWvkXO6VdXfF55KuO/ZD
kU/jPnZ6aFpCAYz6V2s6HbZgLBM3MhaINncfaFwPSFYISj8codSxBBIMb1EhajS1
gH9qTu/mE/f3AUd/DHPHDNbv0iZkKSfYsR/Wf8q+YCuoIhjQMb+7ZmXwvLXPqafD
TBGYKHbR0WPkchRSpBEjK9opfdyRbF+mHpE0Gtnsk+tNKjfr7kgr/HtU7ntnEB6E
80G6V4xQ6FxQKZn1APzCJVijnXiM7SvRSc2b7ihvKebqaDOMAv4q73W5oqCaxlo6
1Ym5VMA+jaHCd5XXCb6Yrz24R5nXq8eM4JMxafdwlu18Bs2Zvy3p7iZncboKZUCD
fRg5w6eD8OHmpBFduJyZVmWb2LB9pCx7rXh7WudGIYfPvEtbTBgogFl4t+xb3cB7
`protect END_PROTECTED
