`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JKCDazluxbcskljKFPuF6l3UacY3s5B5Y0ujOFRqANN6kPNUGnjWWl7unFg+o+qa
y+JK4i9AxAjWJdK/5HtEbGyoYb/Sag8pMsHYb5ETWXbL3qWYXS2X5FUajx4G/nRo
mMoAjq9fGH3kRqiZ1KceL891s3RrIgZvSuSGCta4cfXVqxLMCmZC/2o30nz9BXXM
eZRSJueTxm0umsyj4vqpXbjksGpG0UnKbhclYCFAI/e9yGu6RZe+49PP5yBFzcHc
xk7NIHUpcCIjCA03kl7ba1Kmxd+NzXVLA1eAHKb7S2+6YwhS3Gx6q3E8mgzhH1LF
VgqwJVbaPV2rRR8w0GcEtomc4ognkgPS+fxNqjbm+zCvo1A3bjGUp2hPYkS5JXSQ
Z+Q7+DhFeWREYTqHmMVaL3HDk07A1EWqYf7NxHFByvRxgI3WSXs4bYFTpsiL9yQI
BRP4R+3UT0YbHh8y9tbJnkmDZrRL3Zbhrpz5uckHcHwItHyLB8zX78Nc18eryFp4
mnSn661S/waqzM01SrMR175ygQluXArsv8vt2aOkJSE+Hel6uvN/u9ACTHZGjL7Y
mMLFJljSfsW9kQbhTMds4M6RPpaAngSx8ULloIKXqTgtu56Dw2LBTtnuPtjd2mI/
SzvDSHTxXZzkFAiAqiAlJRy4ibCJby9/NZzK4sYMy+GnQnlmiSwhMh+W3514lKMM
ShsQqhC7prZAtR6fxc3hMA==
`protect END_PROTECTED
