`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aoP0AJA9+L0t2H4AIIA+qmUvWp6wrqnAhSC2SHAA8jwEzKsnbCV3JSR3p/PnK0T3
8DcIlYxCp9rvVS5f4cztjSyOuKNP41Ky9nRTKQ01QoXICVUTRK+bILodfka+VEiw
waaxbSUfkFfTcrYqXSMQcZXYO1SVGqsG3ySAnqOAGJY6hRvI3l0VyQIsbUaWkef9
P2gTH69umBDF+wjWgCIIPa9G+WzWZJauRds03ZBb7y+OnxlKLrfO0Sum0eYjc6c8
sl/vJMhOUMgaZqDmZu8ASQ==
`protect END_PROTECTED
