`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j+sYdAwJLN40G6JF4zTfcpaoK6T4PtDZSfWam0yqRsdEt9akvTXxFC5VXFL4s1CD
ygKOFiaFEkQlaKlEBW3ZGNak0MNZNrDGjRPoa0uisVZL2nOXaV0XyQEDit1B1Rfh
CH8gJpB28RMtYit5lKzePJEWuYrUYGx1wQRA7iBjUUMR8XDFYXwdwz2spY/IWEUA
qxmi/L8K7d1ZJlqArR6UR6ObGl4O8TdSr7Wh7IWna6zRRg342JlMNjcBBjf0TLcY
YmDcl2Gx2c6L507gQFCnhKQiNQ/de/tk86fxfBzkRrTGj4NNaOSVPiQSj3wCtoyk
F5/dSMwDEx3QPORDQ8l1RM5dx+CUEyneaA6ZnW35Kp9r79DY5hl1/xMU/OXhhIgY
lREGyobI1nGSvTuqmIwfsN5xJjkoLNzVs545jR991Lx6vEeSE2EsC1b+kRYo2dQU
O2YexON9R5bS46MOCbyhM/rPYqACn5RiSfQZpECgLKXVz0Luig0IkTLKKj1zWVWT
hDRXXjclQYKl6U76I8Evyd/lAFA4zcKnxWsUCjOkRDQRlxYOFpMOxj2rQsyUV7Bk
basK1SCbxZk2W8iFR/8yAlvkAVw38ClQ813+gFXKGTe4qUdgBR1DZs/qr0mAgk1m
By1caTmDr54XZ/eoyF5COA==
`protect END_PROTECTED
