`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IjNEIjSC7nPNsQx2z7+saxV7EdSI55+x86IMvlBYDvwgP91xmnrblJSMxoFKOcD8
gO0sIoWcIY4vcZTUbt7ydc9igJBSmvXl7kyqsiGao6a64VgFAqvVc6IHGdp31UjO
Ey+xtbPxjWws+IFlnL8yHHueCnsHo7Trp6LViteKUw+jsereVcWNbDemyKVj9jbu
5YVLnf6KxZBrFiwF22dwoz7KoEzh1o5vXJbW6FiNWB/JWVq5TspT3qE26yx4+fLI
0ds28qd5JC1V1fnucv6+BwXwGbyqbXkZKBtuTf5nz/xfLxXAThe242O3DWgu6feW
eDKSEnRgKYNEz+RUuj0QtkSYQnNuKb+83xDxzDTzZAoFuXW2DdgHOjBguUAeuZcK
e+DAoIdB5Fw+ZGAfptp937jrDSlswmOX7ctPBcozkC/koaQdCwAu2e1vWNk+Dmc7
tV2PDGdT4yrK9ymXIRGtobhwXUME+YLK3tGTCJ2rkNdm9KZxyXcT9pLVgPMX5mgj
zoj0Zc/eP1Rft5lor58Z1FEB1o8V44PDhym/crwfTo/lpwmyxNyhzrSbE0f4fkC4
/HF8vffq9Mz2No8pxXB5IAlhhaNI7ykh9xUOLqy7dcOuwycfoqQnTT0I+x7ujAGt
jm4+taCnng1GetuohMIMPshP8pu+io0UypmRYJDeoMVwpLAa4HO8u0YB68LEzoIe
kc6fX/32FFjbbYSH6bE6XAmQG39R3sBc3mwZwqqex8ctwAA9JMBXFXGoUFOLq7Dl
3UXEJirstwJI0NMuqALGb/tYMOuFpdutVcArz8aSVlIafEwCQrMM+g7CuBL+M7we
QYKjqPWGatn78HlpyyLRQLr7LcrSiMXVqyq8qHcB4/tR834EJDt21zOqVl0k0tfJ
qWzUT9AhbGQM86BnaOE70U0pEyWgWiWweDWRNU/2mAwetfJxgg7unWcqFFdkLR1P
Rx/cH5yIJyNqfj2mjgUwXlqRTT+1aGXBGdxiPNINGWmIw1FqpUb6hQ6gGwQms0hn
hpDVNrVgPwRmgvywZ90eB3DwWxSrki/IobvIEgnCrj4D+SrelQaV04hdSq6G06lP
OBWLy93NsptaVUzxd5VeSu0v+YN+OjfD6lhLR0bdMWxsU9w7RuMNzT/cOHNDMJFi
WMoSjUv2dk6wF7IDtugvYcX95cU8WYl5z+x8GraTIbbwoxMpG7Eug47RbHdGe0CH
QUI/u2xNsI65r4qqkg1uhHcXkqsJDr7PsKhrPpF5AjStrgYG7QY/HfWHtp/6e49k
b0w7F8KaIXUvgf4cKBwm7kWv2bLtD2eOoZD9X9qmALgl2huXglp4BciiyuIInPW9
9d1FUWMh5rpRDzd+iFiz/tJMpxa/LH4ruyREqlVsQWbcC8G2SCSynPffT81DPYpY
lm3AutfMpYQvk9fBPNdufNkwXDu1Ntf5DtEaLRGNvsCNZ2JORWkQhrva9/snedKs
omEbN8HeQR5mS3QFftE6zlUnRiWesTMwakf4PUIT0fB1Wq+pe0V9Gvcg9iUo0gS1
NqJ/mDI+xFo9PULJhGeZpiU6kLM7YU6EdbgBC0UgwKWwqJVaisBSqJbJ6yeKI04R
3V2tJ6IMj4JboHkrn+IdSD9SeU3KnUGwlZt9JZr6/tiRT6ZS0O2ZV/Udv3+MO6ac
mZUJGuc4le7gdUxtJ44g5BW4VIREFH8gyv7+5eOmMHz1TmVNBURELalJhSM+ZLxO
NKoN/fLBMbX7JdLA04DaGG6EczRE6i92rEYf9017U1VVn4EZpxmn9xeKA5boIOsA
IdOSh3YQCv2CviCdt9kqEHikMALfCNoeUSepKWDhpc8I3uYeheN2/m936XOKFdE7
bF/VVRc8pDCb4jhxcHuV25vXxTsp3nX3eLp2+Kyfhax0JKbYieyybAgGIEB+bNGX
M+jukReFyVD9UcZCOSD73Xnd8ry1AfocrqQZIJ8PVz1y5fWJgCWJXJ/VKLVSZBE/
wyUqgqBfU9GXojfTVNDMyioiBgfkg+zmdlVu62W3QTVvqUdQviXyZu48qW3La0Jq
ACg658zln6MJzVwwGWiXmtz2dgkjmD6OEEWA+sdJFgC8kHsbDYRo52DpoyVC+TvS
67TGIIUBjgjMWiOnsAsX1g==
`protect END_PROTECTED
