`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B8ly2+6MHEt6VnW9hs0dk1dY4x4aFxeUu13rtqme7M92Pt0whfV1g83FxMKq3fEP
ss5sEQ2Sl14aZ6TEOz2USii3ejzwcPF5tnfYudF0wcfuGayqie3ebm4ZnlPZ9uH7
IzHiLQ9HeyyDpHJ8miJJA3EDlcKkzyJxklazASBPWZVO3lr7CzqxexaBMiyvPMZm
RSAse/ymPLW151cZZcvccoMb6AW5FuVe9HspIxjKh8lqVyR8j3oMQhgwd0pbRQkJ
xAVcVzhZHWTu5pme+Nca8y61JKPWE+YW0a+iSf1QNvipfKObn4FfaxP7fKcYz9/B
92gs6APOxCIxIarPpEwvG7D6bGw0lqxMfAPbTh8fs1g2WxiYpSrYBUdhIdGgRhBW
/7Hli5VSMLCixZoPTztessvjN4bsiEYt93QuRQf2dDqw9x8Rtz73B+JAUnhqLSZN
RBkEScJH8DQy2/w0YugLUjdYGSPF1arhmIA7/dqa+xtEST1i8LyMZoY11uu9eo3O
Dz7QrPeWZd6eziXJrcRsk0Vly9dds7kdEAHw8k10DYZJ2Bw7Ywp1HFoYlrbsa7aG
s7lZ5aFAmS/hFdw6faTjjBwfMGlas8m0REX/cnFit9EQymFjNx4GMk8mjpc13oWW
jvRSZY++tHSmfk4qKn4NyxLUjIm515aAQD39nXuiZqEhw5erqWkrPioRA2VQ0tgN
R6GQQaKTs3AF5kmp94vCGf+r8VeHBYfwHiK6XXIeqCexzd/LNlrwa3wXRLN4t+O1
f7XRq/iEnVYuqpvJIwZehl77AWI3WKd+mSzUr0DYknGYcSdtqY+1CvRzI4slXNsC
e0mVsZBbJjWzwOGqA89DjFo68SlVRUYsOd36T3hvIpNqDtdSmF5HdRjcN7LqE9tg
xcAWyoDQTGH6qj0uJurhYdXOjGCXAAhq9InqbAvIom50ST+U+M/NPuS58OHluxOr
gBplc41Keu3YIsYVJK1yAgKH/IKi033ppQ4KpDz0PJ4R3Sze8R9WkDt1Zrpzk1Lu
cY5avhNPAAWZtcTOcRoaMS6Qegzom97jzSzy+SkuWUBdAmPUDsHJkjYZPyqx6/rO
N5sDpMj3xWUwoMPc3au4VvjH4rQ2Zl6rCyGuLGi4UnmUJX4VNE90VgJGBhDdJE52
mdfbCxLDclmPc1HEngi99vuChrf89VjO2VqLnFI1sp9Xu907lW6lQ7E3JkJSm9JW
TqDnxF5BVPTByhIOKGL5iPeC6dpdnWGv2wjBMBJUPxrnhF/aWSYkeaWsDg1K8Fqt
7ET/92D6we70KdSccgeyVW3O0XDdUhL/TIC/f8Sc+f4=
`protect END_PROTECTED
