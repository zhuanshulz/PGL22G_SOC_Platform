`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WA+IPtRzjx9p1vdi5vyq/Jy+AMdIGhJgNY2lmcRhR0Pt8UvEojDJdWzRQSEszbu7
9wLERFDRkIz4MZYcgO8rRebXR5d4rjj/K8Kn9Zsc8NEDMurXXsi2SbDHwHZ9WseR
hDAwPrc4YQMRrfZ8kGCepjs/vEjwhN0wU/QuYKYrp79t2QvM2hZdDs2Ft05dMU5a
HKZ0iJPioKLtMcjHFkdcx9KsmimfksnYtU0zf2LBmXUxMuqUMZMKh9cQLgVDJBs6
b7rYNMLmHe8LvewjovPK9HhcdqYPPFOY9VSb+ubTAcsnCxNQYAeWjywGzOgA80/b
R2tZdUsdUxVuQ2VK3OTT5rmBlLAzB1JDuyCzsPgAXlEr2KxIsvO4hb74MakbD/CY
TXf0Qc5BcIrBlcWNZhO0b4OeEPFJQsZti1HDtjttAFztcCibIXvjZyPGfQAW6Le2
eODXmSSdGrZhJitrkI+kLc/JwY8rBknppSVp4rqTl8YF2qtliMEVmQL9UgnpQCNo
6apcVd8MaLk5BVMNeIySrUmzvgh8FOSwbAEyKMtzrKnDJHLOYYpfhUGW1rlx4H6J
2p+3dGZTGTa2yl7hr6Hu6TPapdB30xYDZOE0aTqPecpyGSV90JTEs0piPhframuV
HEqZOIk/Da2w6E9jBYI4E4FQenzR3sydQ6Bxp+qE3VFlvKarA96lJHyR5WvNFJ1r
JuF8xJDUPIjnEHna5r0s9KVijFqKh9rP0CYCUozkm1Ar7gQbZo8oAmz6n1/GnG4Y
wxAfkLcvmcUFIwzPOAauc2YNOTf+XL2k/NEQEw/idQJ5j4ooNFK6JgJ1A7EVe+jv
xoM43YmYSL1+O6Te8pi0N8qM9fCL3MhZbSjvoTh9MTyAtG1mkav47cTMOe8fKis4
uontmSbvp260YjGW+zHUHVwpQOad2RjFcRzdCYEZQ6xiJUIcO+0wr3G2HU/QLaGs
rQY0gkjQRkkAV7EpRXlw73hCvM5o1ExFHvRrF3wkwKYL7qGY+kbpEHwNVtPXtmC3
NoMNtvOCUcDccIO6OSE2zVJTN4KZa9tgjdqSIgFbk0Qwss0FveZM6BpFZbeXBseq
VKOvSbk+F2+TOKq3hABTQW9kuarWPn2X0lUHsqdM0757+p5VorQmoGntEnNg9qmg
Lc/Qh3d8sxt674Cel/EMEAuK8FeA3/+GaC5PfVb4h3NtvoTNvh9PyLWHBHb6keSS
+NdeX0Rtv1gdI0iA2zI7E1F9Hy197CWDIsNMvpgBly9Q5yFIiF9RROPouWxp+c1q
tqnBNodkhyYpPiyZdg+frXssERlNbTE9kTWUDlBYPI482IsedIB/na7t3hU5NuXb
FDrqQKfwzoof0oenxb+hpokMdeQdop+1YRu11SrrntQpky0zjXoV3pUc1+F5P2gE
19llPSjvwWXXKLRH0bEfSF7vLpeR406WFOXW/SWrSkR2UlaeFzUf3W42UCtJ6mmY
bk30NBXqhM2/c06R1+PDY24UyJWz4+uiqG12UHFo/AgshWCY3F3PLya2P+SLHo0N
AMrW+g8LLXgNCYqXRGXUor92it4nDzyMTkA/a+0k3l4uDGWNdyAAh8q/JAl04t7S
2aFZuVC4PfC8xAIhUvmrOGmoOtiR7APRGRmhtQP1bAcfO6DcA1n5s66vukCZ9MKi
rsaI8UffIMBMGLEyEvOJNjHlEsQtqh2i64gEcN07QN6DGAsDgv0T8qzg+RP71UwV
qXy8/Byo9H7iEZGEwXl2Qd5j+laGFOHy3cNkxCn6mzOA8d8CI2Bncz7YLnQ5P2bt
T+0uznLr/v82rITCqwRHPBue1JYS+nu2aZlyrfvRN29ComGt0QTG+Cfwi+NzEepY
g4kZDGW9Mwiwld6M540YbgdG1/lA16u2wdUj+ZrcUFKwS2y2jrAuVp6tI7RdGAaI
X+GeU+EJco3LXjbv9rrjQggmGld3JX6Hc6lXM4KPFTsQRHOSeeyBwiIO2pnuEc5p
OfykLPRzHgwMdjTgjI0VKGPL6KAGNVRHDHHb6JsXghnXPX56XinMW/00PHukdeFl
V1KLvlwzEt1P3PaM1d0oyv0afsEO/CcjHOYMhzkBovfib3ShlO4Y82ewUDp1+GAE
TeDKXargCz7g9ycjkrG7O34pc4HHJZm3NPGv6nKSeyNyGj2P8bkpc7+OfdjMH5S3
LelAvnmY080OJ5bsGJKaErpQhMXfKN3+NocXl7ZROm4ajL6h1o2v0981Q3FPuQ9e
tEife+Ep1I2ekdTvT9SWs2hbGGhmJmC6HliyfTE+9YbBbtuYLEMe1XU+RNcnx+Zi
JGT7Fm48uIGMANWH9ZTwDMTsAq1DJPT28jWDB8XCjZVxJA/5lBiH8R9faAOMpuvs
WaERj2xaeeQoTwIQ43zeZ8zhNOFxVJDK2a1Sr7akdaPiwYQgMIkMd4mkbV+Zh15q
TEDO6CvqAF029Ap6GqE3hHS1EQY52QtBrraEkRpIz4qnxae4wBMfB69kumC4Rg1a
TkBbQBX639joUYWLUkHuRgT4wbQLJpVTqnaiTCgOxCsycCMXVfDD/g0DU14Ipcep
e1eI4Ru68SsSkieU+28INWBoWTrZPfPuOl/FV2I32V3uO/zcyZsXMpPOKVwh18IS
tRs8hvKqQJoNoXDHCdzZLLt/IHECxgAZqJpB07orYixZC13A3mN09r4zG2AuTvUH
LYaX4ChuF4kEara26pNbryNpa328NhP8ORHyFKL4KmurNdNNmTYct5ING7Ff60u5
fFBb/1wuz5+6hdt83njjTetit2tiY7GGaV/bx1Rm/M6p675Gz6A4nR3wFkQ4QYqU
EK2W1L7xbro0hmnXeXaAHqD/TxsK4roXDpvg2PY99JvqpdVZYwU0YbdI2IGTpD/J
lQMH6VmOZqqqAhko1V04ZWiyPKupoLLfVOtBuHTB86NeVO2OqYOM/oxWtf2vtLVV
IB4+FoCaGALG0Yq/6QCxxkymgFgmwlCuPcXAcAAudKeMoORLULFIvGWJIUsz3yk0
yG91nKKXiOOAgWZ/gqPJiEOj/CYd77xEq525rfFVdjavUM2Jgd2qBTJ/wgUHtfBp
dEfVmWC5Au4XxKfUwF+4UYPfNoTeZBmvXZTORcKvVQXLcnbx8FEcQroMJPVd1pqR
V2WQ4S5KH3YWMnp3QeqbPa6AwyVmY/+NUWD52hSQk3ku1CfU1A+b0WQO+S6tnYnS
Mk85Ozan+5PYu5clj/2St9z1Odn69Bnf3himkNza7sY=
`protect END_PROTECTED
