`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RQYWupDlExhcXoubmlv8qRSPqnpPotMUBbvMd7y3RqW4AffaC6TDWLsoG5Mlu6wt
hdGsKQEgtwMFAg8mhiS5yllhC9BC7r6kJHZDx9VuXrPtXgqcut27FMuQVAHOfF4x
YXu8wc4ZKFyIcswBlFNIk8AaZyABYFTyOg5aCwrCobT/4HaRivK57Uv1rbA+qLF9
t7JFzTpGuqffoquRN4ffGZOvZNjC2oZjNa4oOWfVhsj0BDFNyV1B6e0rglkG7n/i
b7PbPlzqY3Fpdoa3eqIsKv2QteO0MhJl1VgG8LVSr27DJK1vNraNqgN4Fhy/tdrv
he/KZk4y2N3Ne36KLrekXPmYy3vELLheuNzk/sDGeRkyNJdE6RwvibhwUUw/XJ8W
wlsBptDA8v44OeD8TJvQgvo/oeI1ilnUXXnbUF7BRUn5FzNA7gL9aZBU9qEfBZi+
8aTa4KpCd+NHUVNOcSxJAXz7XnNWrKTQXmyON4uEQluP+A3fb4wg6wPTgZIUNma6
ZLgyBuQe3TYYUqkDJ2DslAZ+LGC+gm6/JqS/HWB1G5lcb+LhAk3JsFeLZNm11GBl
8LrklPQ3kXdgTV3hUoPcfA==
`protect END_PROTECTED
