`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KEPLKUsrtf1Waf4yih71Sp5+fwzYbOz52I1fai6WHZ63tHqpGr8VZgl4/WrzsWK/
MGmsulbU70q1lr3zvzD72o7nHbVjguNyFRn3oJpGxkLa/e8WgyAJBZS//Mmnp7e7
fXj4U7+mHRYqHQAJXXGM1N2BDSCjxlepnWCaJQOr3IC5eAGACtIbQA21B+NeEChV
Ihbh73UtoM5VVR3v+uuXKNNjDbsuf4v0nrCb+sTHMKojnNGsVOTHScYYS9SRRGGh
bYsVNqgd/EC152odnd981g==
`protect END_PROTECTED
