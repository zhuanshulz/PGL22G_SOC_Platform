`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dJCcS5mEoyjr11ZYCqUw45IUrZ4AOyzZwaFpfLo3dj2KyACPomvat4dcmOTTiuZg
HlR502pEfkggrNcyl4nkGwxX1P/ook7LeYHjZA44Z4iNnnNXHsOZqwbgTr40dG8t
DrEdckOHzBhHe/gJSU1aaddPOsBCrTSnn+Kxrio1pccl3LdLFhPmSmyKkvk3BoA0
6OjerNkQTgs5OwGydhf9fja4yCaRpxahNi8l1uY/bf7tu3MacWV18xbgaY69wT1y
lWCdqx37lsxWyjdpGk55hK2e59MDGvTHj2syzi6fkc7PefzSJAT6cPYkwhivyczy
D+8uc4Y0OOx3C2gHm/AAhFaPkRhLoxg1Sd0nDpgVA+UEFOhfYPsFDv7qyP66UFHJ
M/a7L2GGAtI64oB8m8o65YuVVuS7wnY6NDZygy591R8NwFr0jDn+juiWyaRIRgZ7
c85zMTmClcztyz60bQtXSCK48yZenisfumrnkkolek7y5uHaGTzx3lwl3tVisVZa
rvk6HHMSGJR1F7UA5e3kZ+tCcwdv+sviLb65s9Z+8YKBn1zBAFZQcerwwMRrThQp
jlua/sveJ8k6G465aYmfYnyynFz14xdntRH1IRBAu9FGTwKy5YRlQBbsBQuanKgX
I4O1ZsD6k9Fmlk9bTXmoRJOmG74A714HhbsgGGyHbl1tZnmOizdaDqRkMGRsoc+N
+wkmxHuMU9GJry1SvSEWBCOvA0tAxkOUiBGGMHzMsDIe4cUAR4alsWecoRiDHxEp
dW2enqme2acP8jSWvt18uAvEnKiNuys8Yj9JyU2pQVVDvt0XlkwO8Jwda2iicth1
93SkA6z3A1OLnIqPCjvNUhzqUZg2rot6AkubSveUDNI=
`protect END_PROTECTED
