`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oTddy2MIYgktREprJdfRx2/gHAY9ZeeZeGVLWEWg1bjBtcSnU2J8ZhiU/AXZX6Nu
NiLJ0GciViKdP7mhXuqnGRXPmO27xyAI/p7S/ndPlUWmAQakDU+qyRFqoQnMWe/r
p/wPndO7ypWf8sPWir761Ek0CK6DAVOTGaqmGSixmEDpT1+yoZYmfyngFuHGeQB0
qufp72icjRRLAF+xL3guP5/rSvMKvFU3Zg6GoVd0k2LyJ2DlsgpE2DcmvEzuBbXi
RQrH3sQGZTTiB9rNDdIRtTZzqzwYH5wLxj/YeQsRg40sf0WI5X57uoAU1mFEKvOT
aM49e0NSAayU+45TuHMTZFj5BDsAR77lKYziZMdwJ+ru2Fr6p6ePno3f7YC0tWLB
CWp20sf/HpTqPJB4z5BunnPF+8+sdarigX0F88Fc7BD7lMbQMII0wsVuxlLmpuso
S1sRZaKl7iJg6rU3GJwbcm+j9Pm/3UPQyk6apMrjQKTv6/HCMwNeLzPv0pq/WrOn
B2vZL/RHXTV81M02SCgspKJLWhVJd2TdS8qWavjdt17cR4B78T0xeHd8Jvy4e+vO
UQWoXR1vPUSQl57vUZUnNeheLqZnseVfzXBdapq7u2lCu+kBJ/0da3J/zresUJCM
ixIWrrbSVAcWJqXKwoLrJfSdKmOKEFuAKEhkkv1OuoSJTHDgXeCVXpzqeVh2Qq3h
`protect END_PROTECTED
