`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8igcVMG0McEM6SqMLMOYJzklXDTFGAYheqRMK8Z0YkKFHyuYbokmO7rWJ8zp3XjU
wxUwyJlhncvuBpDB2d8+eYe4gbgoUoHnoG+VH4iLtdauaIvEL6PKwBxUz+ntv76H
attPkxUyPaOOs5f+sbpojNd7x4KtQ8IXJBqliJv6nURMEEies7YQoKiC75DqsEDY
UhD6QVbSpivdZDErh8HDjWVhoZOtHlLsT5lUrSvGot/2zDEWqQBlA+2qQV0J8Nmo
n/7qcxXBX9bAMa+OCUMaZJqER9tQCVbcnyCAiEykqss=
`protect END_PROTECTED
