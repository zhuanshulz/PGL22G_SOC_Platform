`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b9JmCZJN37vY/wREyuffM1gLUXpdI0Zt4ZG35jvGjhkIa17a8PybpUFmzjbG0UuV
tKRZLCxTmKObMOGxo4X5Xixt8zb5jKb0sOBdyLA7ygDHJ9+ZfSOEPpVvo5QBZsoK
V43Ok6XHm1PvyftCAgO2ga54YlNkLGz3x7lnCiqi9bAtbSndcP9RnUdC5F8WlCnj
3WZiSZZ6mJNiSJ9GEQtZbYBEuLCMZH4Hd/iGwwPdvhIth74GtcqKtEfsdDsLeaJ6
NWyWv2wAYcx+kiHQ1Ei5l3nkAhUZf3b+XDHboMVQmJIG+KvRsx227ZdR+d2HxvJr
W8stAwWR+jsOLN+P1xfH9huZQqocswbZeLbVb/88EwUSLh6U8/G1y683TNDqCHSb
dAOatLHusulhVoiUUSLD1zOweD+ta/hXx3tuleZdQivrvm0qRelCi5oqBHYvoP8c
ISGitbeuSO/HS41D07YTt43tRkwaPNIHVkPSX8WNQTMOogvPGarz8JjjS2HVi+XD
BEOrDifsEqsAU7x8Z/MEBMiP8cczwmWVJ215bJDGP1kGKFuvVkYVoK6/ps36ZDDG
vt6a+U27Wg7W6fQjN+XJBlBdvY32W6xGg7TqNZvkgZ4fzEjbjTat7vr7Idt+MzsF
Y+vxKIbdvrfOVQHRZohF2TnOA9UJfP4qceGjgQZ7YDRarQFiax67+jwMeipJ8bVz
FmBbFtm42JZbcC0ZifuLwD/DbhKJtwrnH1Im1DQZqJELdOzu1Lst670qheRJOZQm
bXvlYyQIwqjnAFv95VPED2bZqiplxswAcZWKk5/J49mWyt5YH+4skX0Kl/dferdp
frG5jLw+IxTaO6IVCnTWNvD9zLHOsmBT/Hflx8jFqi82A4Inr0Lno9/es8O+EFBo
d5PbWlHzBa+yfhgJcOU9MY4xWyhJlWY9Lq97x/mU4xaDxVINY6qcqPtp3Y/wBvpp
jaoRv7TfonrVGyvBQiKOI5BOU5+Z4x9wll3KBk/LF+vALjyKuULZ1WswBXUhVYea
WZn8jBPp8pIg/wCErR/YVYVeoUFzAi0agc+mIFNrX3/IsG0gSdA+XZZSzzC2Gf+B
c/ksI8NkjPTF/nzonTSW/ucnErgbReKz21PjyfQgp9811E4waJxz4er7HkDvGlFE
LE2bi3P5vhMQ1vNtPIo0pR/7oZAW+yGqoASFneXKkH/8Y58M2DW0Ds1IVedlHysT
aTTPGqMXdPt/UDk4/fXQ9t11u2M/czBQdJ63n2EimhyPVLST8yvHShNytP+mGKtP
zyfKbQ8g0XWpM3JZvhI1dNTtk7ipsEbTJK/Xt2cK3W+DA3iPc56RV5cS5Bpt0MrL
JTCuDdMizmx0uLqBWQVSU6jqj30tSMShzc7nRm09jkmVaVHhAbFxWBZ+0JfDLMWK
kO7kI83/LpgYOynBZ4Swfqc5WY6EMkcUGIztwxl9uj3gpI7xPXVPeNuI6b7OKKzG
cYzHLXy1KlqbI+QeDKszwkENG1dSFQ93QUFuB9ZEqyqVjQ4SuIAUR90Y4D2jiEac
t84f/Hr6wfmcgYhopT9xWbZIi98w3GgX4VJ+3+DjwqRVOIPxo3i4xo38EJuYg/lB
Y+QXm87jboCllVS9wsFYkgCJSnShS/dvhdaE2xRGzP+u2qQ0usXdxfwr6f6KECGg
Sfs5ov9+27tAeEGqL8qpB2nqNMzOsOsjoS9JL9cTCe50h+rTS1iWB97tE79yxa5n
iwdBloAMRCoCXp7QzEXD7cKVJEtCY9O3DrE9Hbr2DYGGOF7mMtq3jZbkGKRCmCUx
s7rC3lvOHJsI9U1yYF/GLqmj/vx2YriGzz13OKCOId+kFcvLSsc0EFhqGEX7PhkB
YaO8Wiyu3z/rJe7r6R2GaycuLFeb7pk36BUxuBtZZx9Wy4gM+oyaKLK2UdJ66xUj
ciyszh/IQU1El6N9LwCTIMRgLEq2iWRrwf4YEosb77YrSCzhpf1GMCmbSDkKJpLe
YkO3DxfgQDnBQSa07OzuMuHQk3Hy6hRRuiAQ/F/vsyMaFAJGU5Nr3Ju2TvNdeDON
kfHXDk5TUB6e8x2u008pVo0ZYnWBXbSC7/awTRNYsLwGyBtuePRad89M8qZxw1sz
8AAtjPwYP/sBpJzUKZAy1NTXbZp05T9QFaCLqu6/AJY/a78yEzLvUZusEy3t/gjC
uSpJBzwKa2v5vFNL82kjdh9PhD2EolyKi+uMrz48PRMKcMwMZCjmdPWdZZ5EgKPA
XTZTcmw+SnD9ZhFttennEyiN0ODBc/NCMCQNppRvrs00JXS5uQGbvAhpXI8o/pTo
JX9LJQExeBfhQTkotYww98zS+zsrEf6wfjzBtsrxhRJoP3VPUr+s+d716MLdI4Jk
NPeunnep19fNm8UogwpDgoiDdWeeF4x+esSRIuW4lu+zd0sl/3mvLhOz7PGIaLXc
5oawWASGJlZg4vxvysEDx+VEVCZtVD9pKIe5eqbl8Jm5CuGTnaL7/x9QH88H7Cua
P+0mSQljECHVrA4bA5oDZ1gfNb35zr3lmOJAdHw7z5Y2JRTA/JQ8E6Tq5jEu+fIo
cUDjw5EwNTPFi628PPWMHBJNhG7MBTW0/+fa1kMt2cjlvvD7lhCjcfvTWkm71swz
xBJPiaDe6zYJj975pRKnV1r4y/+RRZ9pvOImlVwxMvP5U0ztGJq4OX2IungRvJuf
R9TaC4+XjnfUjHKB/EGxYm09w3eKOiINFBWrqeZmDdIrYz1iu1QBW4f0phUN7v9q
/6BiejWTupa1oqJTqdZc+4CZ+NUgWzyXH++wIZD2sUywYpjSfjL3CHViLv4I6U+I
NaV/49XW5eL+RzUz9D4NBld73Ho/aPO6uCZapdO2k8rdETmnzN1HFE43h6qwtiFw
7Nmmr3unqpB8AvPDm7S5s8CnbrusGXm1OxGHTLixaFcmsCZcAa9EdhLIJ2fmiB+P
0QaHAdGTsF/6HLIcWQLeG0dlRJQJPSAf5B1xXUK/2xxHZiYFLy/wNkInXntWXyuz
il3mFviexcjIjKSSsyaKQGI4dYfQcNjY5uwqr7+qDXpq73pEFMAIUpZz71kfF1FC
uU6IO4Ci/23zpHYjLzn16kcXJgj6lZiPBn6Uex7yR74tbQXYeR1/Qoil4CGoQJeK
3arrDcWE7C4KYhpXQATU/LcrWOlkrHyMu9crVXbT2jR0cwlTID3h0Q9Y8bigpuu+
0ZnasUME+FjHXa/hEXPKpnkvAHP6oSsX/yjQF5pCZVCF8ZvjK+OyEpZPIN4azfWz
t7eZci2GnykRzA/fEWC4g7cLF3O2n1wvP+n7N+C2OoUoSNc55trn53sK/FPMhBA2
fabY8CdVRudVbpxPzuUHGf4TCw0iV7KISzLtgdNfeBRR8Yomepxt6VSJUM39ldh8
UhOrj7zk8HhlP5u5J5F8KLR3a6aG+BJfDTICnC0LmbhyUNFRAxAbl0rLHijGD8AY
F87T5BI11FpLhJXNG7o0/TUhGF4MNZHL6xgz4+Ld+iaXI1apsm6Wf0IlVFJmcEsR
g6jcjnpLNr+nmdLpA40LAcT4NI+wZUGrrHEiHsa4ywCmuoIJdLejtyd4trYuQbB/
g33RRPGCr3zEADsko+7UKzOC5Vdkj0yTyz+OSXcA6dwNZyU4U6tZh3A5tibdvIVJ
UjH9s15vlmPHvAuMfmOEanhtFh1kzWaYTPYlIdZrjGEegyktUhPSCiy68JNzGUjX
I5Hjo/SbhrxV7vaTLIS0V/CrE3fBnf5kBq5hevccCz3rOnM15jELH0xl86Aqs0T9
WYbqYEc8TiQU8+KZdlIk3ljBxYWiV2d0de2PaBpdMTUYWpnaSL3OHqTHWg7l4nPF
FhNBsSMOn5mf/HXxguSxUIrS02rso0M+7a6fHzUWAA077f6ghaU8LbrI6Byyiz5A
bRajpTOpzMYoFFz1o0s6eA2QNFDzxE3mQhdw8OXwMhrNAH+yNEbIgftyLPabtRW5
uNtBROETIMV0k5zJxxdAUAkR24FBKe8BxLQ3/6+7Puv/HqE1YDGSpPdE0gz1aSOt
qjCo+s9ZM1ARz5qsNWvvCtYkKUofPIbflP+xSBU531pfUcmzsVOEsJ4+gyt1RhW4
d+vE1xud/J+gjeQN/EqbFjw5c4ynURrWkevAmR/PTNM+ttNdrzewoM2dST1E1NEo
P5ksrtY4xUNRIjg7Gf3vR0Gs1SXh/Yfs01SNjtn+3CipA2CmIInBY4z+hn5vrECr
5vu/DqD/BylMnNZbH0pFqOIZGpGpqM9sWxoHIZyvdq+eAKGqLjwq068nP9Um1mg8
ZeHQUx2jKPuBNUReO/ymIWLQ7CU3gFk7f0bYNKWRjVsVio7dg2Ji5gl1opslra5K
4acL9gll5f1GTt0jUO2mobnSCTD3lL1uPfbR3mvYlpJxuWAQRMvR971N2BbUFbxf
9PABxqd1HaUBpE2Wl+N5Wk0PbEws7i0+qw5QcilE+ZUBS0HdOy7frQhzkWNs7iwz
CnLYZneyvbh9xXZYa5QAicquC3t3bidKil/jpSaoKuw9u10yMvI7Dl1TkBAwvT+v
C4XtaBBk7HUCae3fD56qxGkkA4w+YW4iGd/W4ATlj5XKFXaDDA5SSDZJvqRcpDiA
Qmiph7B2fqkWquw+m4u7UjKUJdjk29xLf0Q+pQkRkjftfKXJeMd67DRs3tCCDaOs
V35DCBAEg06aCtOxS0/Nhiep3NnV/H+YJguMqL5K14rDtgM+XEgPtsCF78StcEqU
rPpAaE7ZjYszWhW4arS6VOG1nH97Y6nnELXcbrZF4DTgB8UgEIWfwp/upo3LDMxo
sb2sbxKREn7+kupOBlICDnZ7G1e0NgF5gYwl4cWsv9UQ66LqH+TdK52L1i401vGE
N7S4iKa/gaKSysMBqrdnpG30FCX24Wz2RG4PnqXCjXI7he5CSM/E+YtWqOqV3jU7
YKHNFY3C4pg537PyO1U+eXPGufAzV+Zffw7K659a4OyjanRZLkQ+ao1UvEth8i57
KzQfUi2KoGRMo3wLLf31j7rH54a43c/VfcZtUuJu/I4REy5olANoSyeOStZLP6X7
mZOdYJgAQvK7KptBc062TtoOZL7pi/jUNfaxPBjOsztWcR1HoTdoi35Ckl7xDC3t
PrXzwNjcGhS/EV1C4/FqlAt/ZWxC3QurBk6jtExLK90A1alUkCHEB32uusm2R/JU
bK/hdMOx8WLRjcP2M9Z3sB1zyRD/QMk8L6qdK7TtQ88xtS+G1edjLrIz13ZWBRQx
GX1kctrQpEPg9CXSNFX5baTOmYCln9jiwAVtJREI4RlXWUktdRx+bxcoWBPEF5OL
ka7QWfLHDbVimrCubAOSLMoDMDsRw1ZUmpn13W8RigezhnJ3D+q3f+cqPGEAydGG
2N017MXjGiDnmyrrtz+s8X3O0wF5z96G3jbbXcqgaml3I4rbr5GN5sIPBmdcRNIQ
R5eJp5A0zLumg2uYqlAJKeQzjTVrqT4FEn0dvy40JEs4cG5tAtSp17stcuFMSJpB
2oi5suQcz0Ap7enDYXDFr7sk7Z1ftPg7kO3DlXym0Fo8Pvy8keoufwgeYsAqVWdG
4cdQxglE8E8kUygKZN1Iyx3EAlmuJo9xW8cIvuKoVNF6GUj5VhT4qaQXkOuRDR6u
kJLwsMTdL1HvlEcdUjE5ZKqF50/rPYEj24U+KKxaXda7Jnxg64jJ6HNneCvPEakl
1rwH4C3UvhUMFMR3OtjUl8oMzZt/O5kgK3No8eTGxRewHsWKCSZOuo94m8Fpkya+
FK4JOQppxgQf2/mjHQAvTY/UIfKiWKnyXShoUZ7/JSk+H4ghUHCeLNgE+Lkkeasj
JK+eUWqf6Rk2NAko44cphPevqLEeotBf77uXpB/0QtAD2gSVWNbv37+R0NLsLIhu
GhNu3REJykenqoL4fBOxDvjLmG6N8hiK2wQnpEjF2Zr/JGkonHQqK/MKBERPK9wT
tiilOgIr/G24k1+vyQTXwaub0zcMG7ahL7JNhC/ZNzurB6AnHd72vUmt1IeT92Jp
I9eiX40UuM4oyPh9020bW0RKxhn3npRX9bHBrfd5eHnyIbtBYypL4BD1UEcyIvdp
WcQR/L48OsSyzzANaIpXDYbLVdX15meBMQEno+xyKjP9X5gacYOIpShvxYjj3/CB
TDsAuSuPdqBmK3A/7r6phUn/dRTIfJkUuOjO5nKTFe1fcWE42ctl0Zk4Nh1HOhj7
igOf9ry/abKfg/RFQpS1up38NoLjVebN5elDdRi4CZAE8uu7fn1oGpPjRcRx7yii
obwdQa3GpmA/Jj2ySjPKapP21D+Two09Hy0QgYJEj1Hy7vBXTIEhdQnAXcBerwy2
KFVkliK2lPH0NcXUmToGDObqgiY8VrhTvK1+PPdvs6IuIGUdrLs1LDC9CLmfFs5+
yLYQzdzqiNrZ7I4wV3AzgT6oXmBh759nLt7LfY9JowcMFTbSGhI7629oor8LvNWl
Wwp8GUAk1Iy8ycril3Y2urRDBd514eOOMXTrXRu6eJoIrTdbfMQR9Be8Zi0Xoc2q
MrNI9+zrqvvDiJIZogrNf3U+SOiEKk3RKFwh9gwdFHJV/NWT7tPr0EB8expyquU2
3Pth0g7ntv78tXKzQkTmMbCo5XyHCWV/IO8FAuUec8eLmJzdOHVwWxeAYfQ/hQ7o
PgohLuyICzXDMnsXDdqor7XPN6ErSO9JKoMZ9qQrF3Tj/JD7NarBceN3FwKl7HtQ
9dm1vdEY4I4jW47MJKD2dmOmRon6zbL6bP9AUTOqRev+h44AwPzfTXvSkV3vL/b9
VS9qAqZczIs7hHPLwc+iCuAdefvFf6UQe+unornsoTI3Vi4Qs6UrzY7gFgZ9KLEA
Hpi6xEFYWrcX2hz+MnqG9UNIW3rR6PmvB67uuuBbKfVOmEp3ucxaWqHjDZLW9k5g
gdslwpLGQy2cRJlakqprJ011WdlSeO4xBRcV8Q1fTm2hZF09rsvhPGWidwMXF6HA
iOm7oC/3Lgk9Ntfipvze7Fmm0VciBhzcok/9+K1zFX/Pncajos2T3nUFXqxi3R5H
LUZOVRTg54WnbmlEDV59PnrSA/oE4Q0pXL6h6OLrocx352t1ivi3qnEqoVcfJ5Jz
V3nqyu3X70vDf87VeTyFdEM2naMXFHcDBfLzgaw+K5hWs8Zt7pANGhTdqQhb1kbI
S0d3VHkblxv2aiayUoXp1IkEMjGE/GPjFAlNCMgQI3wBXYF+hX6E9BQBXzvvBi+b
0G+QHeVMkjNfZ3AjJarkCO/KGxWeSaq/elp9KHflO745DgI50Xz9yPo64ijt4PpP
AY3JD8PoIlqUO0ygigOZ8UXa2sDMAkLnBZ+ddfWjrNiq/bN6mo2KjTPqPyTfeyUV
3m1GXAuxzxvvKL8vFSUb1jVGuuXpR2INBCXEuvo6WvR650UwK7GV4EO8iKeCEJTy
6z5LdKoLxkNJJq4OasfO3KNPtAlu1PqfTnA522gU/tmPq/W3sbmMtogwox6z4g+v
jigP1m0rfMbwGxX0osQ/RxR5cT7Y9kxTQ+yIL+2BXaa9qjXlkzeEc7/bmmLVP5Pr
9nmJ/CaGB0uFFiPUenHdvXwc4n27oLDq5Gj2Iavc4oEMBRmR+L0xm/XAfdXoRM9P
thapR4xID4ZKeryvgmqkXpDUPmvhMnpBgUUrJ/fRiuRFfDd33xkcXhj6zjRI1DfJ
YiEkFQXtooeOJCsA+Qb3Yj1CosYR6miMWohDNQbdVCDmizENzmUFraJSDMFUfALM
ymRCOZtS2b2CWoQ5eFhkdeBF9FQS9XTkLjIyZy+xoZkdobkdMOahXagR8ZIDoFun
44wYETPqfS6XWcbY3QoT83/H7SFKJXKSizWg763mT+PEj48Yvowock7Bo9qCrO5U
0JdyM+kRwzFD02ItbRcXf2oHe1VcsVs+tqiZO4sZ9zEDwGEKBP8EBuQsffvKAOdp
9vtxC+LDZ8A9EUXwEK0McH1fJ+auTCcG8UXSaacciXlGBo9Ju3CCgWqNhcZqIUEv
YE3s0iWQafbBy2ALZhklhvxa4Botb/BB6HdMxDY9gcjwAKLSylfwQfvnr95artmf
mplDuf9vG1D+aHLI/uuE2z0KHzm74C50f9EL1okIMo6F0YSq2VKhWM/ZQszKcTeH
QbUfbbjWVDDyE4wM3dhlszawor0Kcs4LpP2cQY68i6Woxuq1Y9YvJtZqJocxnkD3
9Zy5/XkjX+REk0bdgicRUZFnfZQ4RCS8jLbVtP87UTutyN7GEOebiHpsBNgM9P1I
LaCjG5Ie3yo53yWnu7+plr6zwt/2VfPyCIVeBUrvFSBMZQ3n3pMGqednFwSDlPt8
QK8FJO6Ku92+9K40BiEOQluP/liF+yRXps51BNU1utFfn3sEBbYLyz3UcATIMPmt
DcN2D02JGMVSaw9ajKRGcWYOpr11Cmf6NriZLWUfSENzR5aO0yWANz2jtMGzyhIC
3B6uzzUQMNuvPKmRu4o0Jd55eQbycuXKhyUwTQLqAoniYQft6G58sWW3VYFeh//F
Z6LtPKdsoDaR0n2Z3/+RfnCkXgRhD4dWAZMIIlCGIaX9URD4fAYCUn72cGggIgSl
dND1VkwKvcw3QqwXIb7moi1xyyfASRoyV1gmxksFwiJHlwDt/j+jrIOz19sLFVRs
t5Q6r/5ZldJPOZ+9O/bHpSiHrMDPXmB1XaGO3uWfzrBgekJXvnUUmZU+D8Ac4qo4
eJLi4FpDA/1YPcNg6Bw3J9QwTojQ4b2gjZmIR3vHRsVUvbHXlN1tQgzD4wXgbrdP
H2349kp0gAF+cWcLfUAgbdOtlQ5sPTkLseX+PG2WqdUbG1x723ADi2RL4ZHgCUug
r6Dc9hn6fMEImc6TmL+hEjElSeZwsvygzcAZoIn6ays956y43WpUwD/TJG6AYv8j
nKNnXIbIaJzG1EtccdEnFqa/FQPhxM+Wi4uvd8fGUlwkOuSEJ6sE+todpPdni8gf
qWbKEPZz6jZanOk4XJaeHQt9pfLbPhcZFPQrNpHiyDDZO4aXTwi0kOnB2sJwT/QZ
izd0/JwIrc3zn1q0uXax49NweplKWCaPU3Fvx0KIGsC2YSOZWxpjvKJWQYF05wEm
SAVqGT/MUZyqAux9mbwQYTSLuSuv9JYtbrmiwD6ZwbfWqBKtQeV47CEvV3VAD8pi
kSpcnB0YsAL3mJ4iVR2kNwbNwDUmWAURAFc29CNJCYIVCsK/eYXv4pXf+td1EGMU
M2rhQjFE89W+dqa2i5mDh91eyujBjy1dPYZHAN1oi6JMFiumhVDPF6vn/AZh0QVN
OxlQAvkhibHoiEpDQS70+Hg1nz64HFqDkUXXQBz/CyGo8ZP+w1Qgoz7kY3FF6k5y
l1bvR3wxGbmYwJSKJNWcrNYizlsyn2Usc2uJWto+mDlK7+1SlG/YaXWtPjGUXVAv
ZH+KY1p+Y+P5k7ZNn1GoY4rIhLj7OsJ5V8x1I6sqj2yvjHMy0HpDvFCumNVWLUJy
FNtDUOHv32g7t716GQeu0WymEarNBj8DblciIn1qruFZBbp800+9U5RjnFHdmO5X
iWT8lRqn1WuASmju60prYuWNN9+SYPqAsyuoKmWM603CMJ8ylCfuVE/L2pMPRMjC
H2WZIs2+fY8sePCDywOd+NaJok/i9i2oD/YC37K9VdoHBgPuNhYYtIbT7dCN5FqM
q8mv4NI9OooUqP80Cyls1GBuDjNYCF3eQyLcD/tKwCyjjZfUcF3NRQTTQaIym2P7
jFq2PMSdxLvRxQtQ+I6d06TrNeirSuSfbn6ZxP8wBFWeqT3EpbyQJkoCzYZGpJYB
gQJL97YNMu7I95OfGfvn+XYa/c2DpQgRcaYYRvENeF+lj+MC8ISP2zP6t0Q4nYYv
ktTsIbgrG2FRIVQBQL+yUuqlWQevkHtfOeDpB7POm0x5svXAGkpJUota31GD+5jp
842SEPLuw1VW88NWNLbNH2L61VEMVxGiBHTlRXk0Xfx7XcA5kPkBRl53OW7LXeEh
mtXsRFoEmG74vSL51tJgf/Xx9lHzC3/vRCj9/PDQfSGzzXIoJqkj1WtxftFt+KAp
aOyYi+/tarIjYfXeGFtn8UQ9ukvognUAksTZRTmuoSjFjdGCDzw4ilv9gMrz2qvO
Ls8V22Mtfwnpy7xvCKcqqOh4KnvmcUboNQjCRBn9Dh0L2qHBFPn8/1QBYaJ/EX/z
wjekH3cmulO53JbZWbsbMRBQ3ydaY5jR0+WWFbqvMpjYxUAragbukCN3ADj7asUQ
8XakY01zRNGdtFN0qgO8HQkg2lKKVAzdt2ySES+sVkBRxraLgJgMDTKtvp6TVcSj
ijcEGm1ClgpXLfTqgrMvT25W5qRbjiAg9ojAuI5V7p9LKUJdz2rugfNMb0Ovvlfq
W/hjzKWi8KHplTWY3L5C+5jJCUfi2kdfj1g0B7j8tS49X3JAkiiHZkdIKAPjw5W0
tkGkleQ9JLmg4PMRSKi+NJWxJunZ1Dd8DyW6HfYyNbQV8Pe7lN5uBGvU2n9gDl/u
MJckIFBKjuUh8L4pnq70vUcfvQYKQK49d9FawZ09d5K57A8aZzTRTMuEULbFU7p3
GpPpcRyQje0LmoO14PtqQvMsXqcx4VK5yQwVwty7XVcFoEHlYUtLHo5pR4IOLYEq
hBgRyhp74jbWLBlHnDyDuipFvOUqt2qvI4WLZ1Ca8gfOA6TOLRZ3NF3+hhLI4VQR
/RAyzp+e+4UAOWzAeqeNb5eoECu99az5CAdErFp4IbcE2dr4JNVYHG2/CfwFiYpU
8PoJKdg6Ft2rtCKlzcIG+fHIP5baqv6ZeSbhX3ae2n6SBsuUdvO9qt30aiAXPf62
gPDo9m8J4k6ObVzqV1zphbJ1cW85ojc9hKkN9W0DJ8sSD9njkVdz4BtELUg78mBQ
Xq36T7f+Bd4mfKNnA0T2ClSfw7B+I2Qpw/8ycJD7dAsdszp2XAkhG4F6jNaqYUTC
2GVrvf0SGHeJFFUIGwkpZe0Ol3Jrte91baiRK8zZlItsY0Y2adi7zSIBySBwnSDg
jOB4bdE2I5DkJSEwGIHSswAc6WdnMW2XySbHu5/sFVOPVaNiTDowJQarXs/P4q3u
A05GvZfrEWJpkM3mD1N9I7H0rvqMAXTe+qFPbZ9LFguE2yzMIqyIs74L5rEiw1Uj
wdsZxUJLipDPOHJnScOkCSmc7FN/sjrG0VUpL1C9tD+YHsocP39bZQrVsaEBnFUi
yg+YzhieTRaSzxNEkq4uLmE9gvqOEEOMdL2HHCjvfLH+iC8jQCHfV+fFmfSsGMZx
wCF2YpwALCphqg4oXKY8iVO3L+KBlPGGrr5LNykzTjpbJZwXrC1Cg7BdwVbKj7IF
wtntx954+AG7Xwdw3iXFWnw557+9tGQtw4ewd0ThxPJ1Rs1dhkUiuAb5zIji0Ewv
jbWxATATxZRaX7uF8nwiKVYgTtUEnizxq4OqGwkTGtGfsZ1GNxtLsmxb3w9LMfy3
oWvmD2JIcwZED4wHJ4sedZ6hI3OSWtib4VcZ483pYksUYzXNp78V+YyNdVAYeKOm
+PNtNRiLwziABvM2e9m3Ubhfygoi3sah5mx0Ubi+nNeomCeK8vRSDf2Jw9x0UrPU
V/Rtc4A+qJA9lQm+W2PEfaT52KijmYj0p05J+D94/S14MQ0aHsVWpvKJ+iY2M2h8
sfFDCoGXYZy2ZQA07IQ1RROfns7/l6p0Y9CEb2HsRKOxAqwCnUxd3fcfDqGix2Ga
AvBuO/WmhoWAuP6XjuzfWJWPPuRZzM/0lpEoQB6vQ7GxhBueHr7eCDLcBgXHXleA
nY0Y1bRKWx4dT5er7gRwzZgh6Cbd587rJF1meNccKoyLxvCFXxTwoGb/hY+4PJJh
totoOu9Xtmx4fbSlHtVyiaboeZ86ppSwb4swUsgqC/5cEo9VqnVKynz7USp6CmLh
YfMqEw/EP3v2f82LUQUcjr4EipW8B067Phqr3kqV4DF2ORwSI0/U745SW3IIDEXv
lgNd5w5iKvHBvymCyPeU/vK/mNZOcgLqhiagzIr6GS+qFfXIBZJOAIkgCHG2cbi2
EsJ7Mn9WvGEMZCw0Ra49Z1X+NUBa+dI0CQjIKBdhNPU9Vc15nZrzX9HmT0XqpFsf
sQqLktsV2e1YmXgPpIn6UA7b0Vc6p+5XHZtazSr2KWw/VmWWczWGMTTDsBnPdgnD
OYVcPSNsl3fm3bQCgDqJNPv09NmszC6pCmlYTsqNAAn3nVoiyzC0a5EOazedtOcq
bPHSIOMPszDUSbXKkLR3nUTrC/Bm2MKaOB0N2M3ycP2hZJWAIdL5+zBN/YpdqiNR
fF8Oy1Hv3apzsBTJ9Ig/k8BFja64cY4YZUvmvmTC6Yn0Fvfm4Uou22W3D0ruOW0O
h8dOQVJc4PEy4zatMWm74RRwFD3UE5PQmw2Q9hJt5TS5i6lCzHF3xIla602aAklG
/Jg6iR/hRpVm/yxwqeTrq2SzZ5LXcJhDtnQfuaTyrdxZoBAlQvTyCGza+mYZEgW/
7Z7inxJp4ZyarEVT3Bj/ujtW1KUIqyoUlkKajXhEPfJNtnLBG6vJzdfMfwgE6r2t
CZNCnPlYR/Zd5K8ipUaOr0sq1LxDGtnAS4VVBhUp+KdY5GhDsXGyv0wPDUmrZ8AC
A5IrvPne+wyJX9g6xDbV2eZhEeTp6l96UIo3RUgZAilb+r/HV4pjIQky6947yQqz
rzNhT8Yf+QDhgGt3Z/9ZPaEACuNEyWciCt6D3Y3u/LBqVGMKRi5FyHFFPbFg7NnM
LzVAhtKq6sXemg++nOsOUbFMEAGqo3TNpEDaDujsPvxE1zGVc+snfngsNduHsdf7
Awc7ahwZqbhm0LwAB6LWz7TYo2dPXFQyz08RtmfuSbLuE5tWYLhwrfDdGvdohGtz
c5sXA5aULj/dOv/+qdQVTRYz/ewSIqiJdyY6C2WcBQ+EkCgXZ5CtXJpo4RqrlMLi
zjaf8WG++aQrP77GtEnknhUmodIIggI65CzsVoSg9gydwZDkMG+lmt/rV8CFex/d
u/74uxlq8h/VNAWxuj1lQHFCxDfX63/mdDVaGqz4BQj10pTkZq/EJ/if7EqDOHiR
H4v9drNkIBq69bGoTy8YZdfJDaaCJ69MJ7cJ7FBfykNWVcJoxfalTJ1zZgtdV9pe
3UQdUZxrQGf7bwmD26P8Ctmja1FiHGBt6rX/WflXjO3YPKW+qzTQ9TF3q8jSqfP1
BIz07KAbrg4CUMJBWoTYElvL9CmLydMyCQ2MrEz+zRW1RnJzp1H/KBWzTV/i4d8X
0iDf0qvSkSewzUuPDqbElbZOA+NrIcYz0/uqtf9gNQ18XrEUWe82ExHnIImTCzma
tQTK0bxc47YF98TVgqp5EvnKIJm2gp8HzgAE8If2jCUu70A0TZMqT34fQw54c87N
tfEgyA+Fo+nbZc6otrSK2qMB8y/GSgm5q59niR/xCNqblocb5gtBN9PC8albsc+k
FJxOEDb8CiSoaMnn/IqvDjJhhAKtVJyNye9hjQ7xOQpfc4FxfOJcFLkoLdiWUW23
qC5iXprxFQBXL5HIT6Ni3M7bO9lrl//6kC4rGaM8DZQ/zi6RjztNTqtZYs2dnQ1t
yEk/56KJ/TxuczhfhsTT3Ez4+UCQl6e6RbF7QUWiotKXQmBDA1cBK1uDLTTLo94N
N2A1hWa7wX9MCebLqcLz89uarG3kEFhCmJERI+xJjkNVqPlXK0KGwqbyHQVq7nNw
YhDbwNsMU/ccQWmtm9O8emME6c12IEJLfgZBrS3S/N7MymMABsPlvM7hYzdrRdCc
lPHKdomraQToYRuRY+K5jFIR1PpFgMo5+nwIGLFFY5Kq5hd1YSW76S8IGUnaF3R9
uThOioLA7B+Tkpixf0/V3EEb3n5dFjGRTXU0Gz+87kmTpQsNY+VlV6F8thgEaI83
dhpBxGIn6xCPMK/KRWMCWtkB5QIxJwNAYmnhLit1utQAhXdHxoHOLhMkK5ptVTvs
bIdDbDNRjLYJolkA8pJD2KXgG+D+5CJYaJLxNarwjdSE3JpynW/WZ1P6lYCc8/0B
Rgk3GHKzEI+an7tpXteMvzplKsFqyLS+c2nDmC55m0P+aeUpGG1bo4xShdQ4a4b9
PiBDhi+wABjqTYIoCBPM5vuN3qdEziX3PifJVS2u5L8BidzGjOdmdRwnAi814box
dRicyCb1Nz1eU/b1aQL3nR4PV4rseHwkVWpGZnHW7o5qtMc4O7eyolSURhX23zkX
DkCkbtvOr0l8sZ4A2Q8X/rFZWTWMpvPUp1cNn+EtPaIwcf8Q+KdDpVHeu9jZeNjm
4WuG3401UCdIOAGj3o7qAjwjOfKxvnRRQ3Ldxkikx1vuPas1FpMM1bfkp+q9Xabs
cnsOKOq3QZskQz9Vl7RvH2LNQKOlrQAbuhgWyvXvup/Y629D5IOdIAMc27KbNtaz
/1rIxfRNjAyq44tVoaO+jWWnSbpdEJq4gWT4+gr8OpGrPKjsTNm+SXPTV386kSMq
y+LvIB9yuR3sR9SPq+wuPA4a6245/9/Ym6YwyvRH+qeDpgazl9++Q5EIBUAQg1h1
OxWqNAw0SoYsRP+cT+F4jZXAIB4J6QCH5tUwVBIxNOy+/eAQzYTD/Zr0ny1A4ZyL
8JEaAu/TiYRJlYc5vaDkFMmlujyleokXHpdSaCx2IWnujqub3goRtTe2u7NTeGgN
0yKdxbtazpZDu/rz3VjjkGkeXbQrvwdj1fe/8ybQEQClLZnGiZSajxGD7IBHWTK7
vuUyE4xar8fgJN2SkvxC2pCRcdlEPyXpdgzV32XwR1b4MJAY9Mcd6Wg7iB9x+jED
1HM1jobFqZxeTtZ0Oq8ij9WPpLZpRRMeWxakaZuwGEAJD+H6g7weONpzqE/1125C
so/sGpQ88xF2ORc7r7zAWOMqwc7uXNBCaIVveXeLqa+mdjljes+C5YCsW88HGmSd
CPui9r+llDkMCXUjAFNxL/W0TfuX6ZSnPgIGr/5/v3xF9UQVn07bvFEPsGipBvAb
U7QWyGYfQ4ZujQPs1evxWMasVFefwA/OQgFfSCscNYejOrK9i///sngpLP3ODj6v
TPX7xbS3W4NoiFPcmoDfthC8nGXrHccfTi+rNnFJDhpuvaWeeiKSyl/NLtxgX+0K
wCJ2WrK1df5sNR6UjAdeJ3RO+CpXLk6yv/OOg0iXqTEvNjvcDCMSuOr+P2nnVEyW
puHlfk2uRkrvk70IYHrMcj9m27NceFv4TJGN4B1TFPNOjnllxxyLN5OswKij9ooY
HZ1+t+NQJ/I5t+Cj46KTFx3aAa5aZKWJ1iwCzqIvyKFCE1UWsoYBpTDHZqH/f7Sy
t0ej9mY2XkRTSTmUHYadJ3rvEkMgsZ8vDnq+XOHNzBOIrcTpNLfuVXG6h9OFHLZf
OvNkokXO8/fTrwCjqDcn3oQEcxldvLpq6uWa37JG56S5VP/oLUd5JdPfOl+S6NxP
o2upHeEeP+TyUoA05zm7vz5QRJmXcOsQ39kFGJ5QLRb4Y5w0jXriFIpPV0DCyAYO
ks9Ht7+3R0EZnjhpPPgASEZXj7wOXSm/7xJv7zJs4zSWAvihXg+2msSFg2+ezw2e
9zqUqLQ1nI1QaQM339LpdL2V9tlzMvUWblqtlzQa2XRxXKj+cF38/n6pkNZDHRA+
GeMvvtLXgDgfuMmZX3vrZ5ahgu6vvkOnUJJmKXIg/AnyQjGTtTPkRJW4pLHo7L8/
tTG81pQV+F+fck+/qLNBOMUy0rzYL5hrGfMxfa0UiuhijuKYCX9vwvnQttQ/7gdA
gtob/WWh3Nc6u6lFNZOAy6Gr1HasbnM99+gIu2zzpkOOwMiFMQYk6SNPFvbl4gMr
1qzlXHuD1/e08bKFvMoK3tmvJJy6EhL332IeQxFmykG+FM3kRQ+pk85QdXArxZss
hnQqpwzpmu4Xuqvl9aVxEts467m48T5ZksTTT44wuAozqqcBEP47KCI5maLSv6/9
qF4aiZcwDOvLY2T35mb17l8p1CEn3yLSSJhwq3+rgdR1fpjMBnw3ML9hlJTJAc+B
5RR3ISle025mnOHCKhJRk7rHcDKrwu2cjzSFvWtstqSjBuS9erWd7ZPk70Xia0p9
2x6k7SNaJuhL+zbwx7ekxa2JBbwnbPyZ/scZ8WlhJ0hMdPIsO5++CaYooRvF0yqy
rHKXTzmkU0OJO6W9OuVdB26vWHHJrNAdpCIovIjH2VOJ9rty3vsa5Y17FhYjgKFs
emni1p7CHlEn+S/zWc2HpNIVKYp6Ow2Hu2RUvv6L7wq/HmsotxnEAzQDSN9ftN/i
zBr8FIJLJfG5MWlYp1c2uaXlmxBmlKsCrIZG0o9SD3no1WOYiavWG4N6ws2epOW3
KrvvxetQ0a1R/mLSvDUuSCMsx3TKj+0c+w6j7Rhp5Xeh5RhpFsyySbH3sGkEGxkl
JxbTOhuw695IwhRD1+wgpI3dxBPVCYxdgjInkZUBEZty47VcT6kX9Oi0QGATpjnp
E0bS4v5h/ceqzryizxTioA==
`protect END_PROTECTED
