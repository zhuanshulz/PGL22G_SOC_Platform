`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Pwauk+jfONmzPPzq1CMiUEGx/+wZbTT4nl5T191t/l3byJ2TGnj9uy6pLIaESjlv
X9JdpgeSB2Ug36JDv4YUkb3j2IFAOwFd4QVH5KSJONb1F0eVQGwY4WVRck03iOCB
dftE+CIeDLs4UevbBTGz9um9PQ2FrpQzTYNFOYnvhhsRFPXV1I+Urr2/YyLny0TB
ZM+I+7aX3rvSYqLN3mWXexodUChMk7rGBc4jb2CMmBtdtjdtdvkuxYclZWv4X+CB
0Fzw1kZ5f3fouyaB/bVV/vqnwjpIMiCYtOfXowdTxw8Pa1jnD8FVICsLwggc6Mku
z+pmXtD3Fw7baqepvMfWO2OdrNOfh2BehrIBQYDVqCNkVUg8YrpXLYcHfe+Vq53r
ldYJOu0kjglnnJcTJL2BGc/blgg1sotRoyw/Dj6Ns8r6s4CIpenqmAnxr6rzmWSO
7zsfsALm8zZTnnqqTEDxmS3UycshmcXPec57H/hCLf6jqa8HUd9hdwmxs6aKXF9T
H4rwJhPfEub8kfmIffXc3skiAq9IplQeYHA3l9WrFYqlxLigWnIYE3SSEbBDQ4+m
UycaX5fH2+lFk+hv7xdpOPB+bZQ26MchNjv9I2QmwAj4ZUby8zkswzgdRiwNW9wA
Yj5bsOlDz7YhjcgxZLM9XTO/sOJGNmLAqAPm7Fe6APHRCglEU87qmCl2TvvS9d8F
hNIlCB9cN+gYOU7l8tI6CTjkBIeeHDVpRwTyOkKtQetWZ9Qfx9gcmLv9eSI+zFQ8
cocyVxfkJvaYhROHP6bcPZo17rqlLiqna+LBtjWcyH/bBQOvDQiRsP+iaPb5GRYn
9mBhPk++qm/KPXveuehPSf0VrTPJKtdPR2mNVwpIa5g=
`protect END_PROTECTED
