`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y880y/hGYruKqj++vEJA01jOQRVH38p4VdsdL0pxQatlC8yGcOKn/T1iP5Ouv5hn
DPr43sEPiF0VWP0juyY9c0AWeSxt1xftq2b+JU6fediHWpDDtp6LtVAfG26pI3uO
guzaR6PP5Cyhr8MRe9uzR6b+4Sjaj3bgBaFmfRC2N2/k8WJnsBTr9o/XElKp5vVY
dqITN+viiREmrcZz6/nfDQNDH3v11Z5tuKxdTgMVUxUAd5j7a18nte+ijaMWivBn
/EKj00Q+oIjciluoQiV/upUjr/YCORoOnMFkwWpN9O+qrIZbAaZiOsEAzbLpudgb
4CkBZeQHepoxP13GS95xqsBLRk+4j+FOCaLaqKmZoXEaNai7BOcPhBcJNc0tHPm8
Nsc42fvbcS+DotKlCFGmoy3vJsWu2zynMDjXzU6pSwpCRbUrByciAbF4WfIlLoL9
iMC8G1B90/oauECM38RMvPddPa7vpEy/LxnuT7qf/AectPcAzDaTt+HW4udOpmV+
Dn556OiOOMvD1hriAfXv5qhpOJXkhgWZV/OV8AJTRM9gI8kGDezHQM+j5myvQ2WT
ut/rIgknjQ29Ov7hnSuOSgKWYLYNvbG9Ds2XFEDUibeLZKRD6LmdJ2FIsdvgWQOl
1HbBeHHR0BAlsfuVHsBsZ1/kXKPLBCnNyv8w8VXBaZzhh+F4JkUFYlLOQIDbfrTg
0/Mw5anybo1q4g1Y9dSG6jEI0MDB6dGlj8pprncH1/O30Ts3bgdMZrDF7jeZRJnQ
XChH5r41srI08wsOLH4deR0GwFLYdsHoa8PeeC4KT9MN1K6S+u9BDg5xPp1KaNT4
lAt0M1CBLCMR7U4KbBQnenpIvRkOgPFDoUBiB7P2lB876pXzvi5lKjcrcwVS67WH
kSTRdcgURGzh6NBZl/K9oAU5dVQ2MLt7rozWnq8wfpy+JJ2/z6aXCm06qjI8opPU
cKqBw4KcN9MMXizaHlnKoVESdX30mZjng691zuGWdH4o38YZ4VJzi6i2ZvZoGesg
hB3PTs2giZi99eoJ3hr3+w==
`protect END_PROTECTED
