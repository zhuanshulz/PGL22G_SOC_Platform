`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bQdavCBDnDWoCxDo8mdyn9PsOWqsAGLVcglPlLV2GNkIvbd4UFhXLJ8ZyANXfo5X
PJ9Yns6gGnmZ5beU/4Ez+l/11d04otvWCtyLC+1RU9j+kIct73OgVcnFvVzsOwdZ
64fema4poq/NaJNhXrMpSJgPSWLJ5NXfYlKQeXLcyVhGAGvCBZUe0VEjonHVz541
g6fu2S1A3L6+6SnWI3npRVixb/0IjG7kAKFma2JT09XUWty/9O0qSCXs76vg1MV6
E0LLPTU0dMANmUBRIeVZba9jQ0oTIU8L/n8IxtVdrKSi8fl41bFnMsxpYYraM7FF
4GUI5NIfWhfbucTXCddP8qp+XPOQlfKaEyFQcBebUqp/DTu3aSaGfGp8czAMVdvy
wD46VXnieWxEdljUA9KVYqSnd9YmBN4Gr++ExhR6Z5vd/qiJEr0z5MWIH/AgxBus
MrhUC7Gj4TQUytRy7UJg0MBwv9vSsqJBlV9YzAutq3+qTGJ72IfHgAfY7eQG7XXk
k5x8cbhE1+Il1gM6XsnBXWNwbmxh/e1GLjOBHWkpb7uPhmqvgsGebhxzEQhltyJR
Ei+8HhJgB8cx/e14b9qyzntpDGwper4DgPfwq+yCqlVZjV5rvlpusggoIGA0GwkP
lZ1GETFCg+NqWYD7FRUVhXG5i7UXzEDTVnO7eUOGX8zgeudGQl1xUsiXTq0MAZdJ
Z7jguqzbu/CiIaCjlVFuVnYOBHzIp0PodomJsgLttL0C/q/daluRMvO7xcNRytrh
pRVoYzgrs1gSDWJKsFvz5BdmWLGEhKXB61VZ+Mp+friR1dobOI1hlUtwSsL+Q+1m
wnM6ggF6Ntc0xawskkCNGU1qfcVkwiEU+BbpszTNBoasT8HdziwqqDqpPD2aO3Jc
XBbdf9rr7p7ymb8a9JyVghvuCK0l4If3Ku9IWmV4QKx50Dfk51/XBIcj44XefjJ6
224vny/Ht7APO++mzG/uhZBYdH+spmAcC3Aq7vq+ERcuOBxSvKbktm3qF4M0vG57
ML7iD8qgAp1etkFm5A0+OqFFvudvzyYAThvs12z8VwQ=
`protect END_PROTECTED
