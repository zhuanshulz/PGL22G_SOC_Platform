`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZzgxhhDg9y9X3FBeItojOKuDsdqs1FTBEsrsMQI4nExOsO1FFkBbQT4X3zSVKbgM
vCm0P4c+PzqihzKCRYfc6ELZv71xWxhocdESboUi18k1bCuMyUgMUeqoSCUnRYM+
JxF5RtZbi6EMZC4j05m0FyGilyOKCr9kxhkSJ/vLYEEQCpUBiyv0AloHLy7vYUa3
yJv43bHrygttlDuZCi/oX6MoOq7Qxf+6d+1cFntXUoHVm5Sn3s0+b//aNCjM2pgm
y4ANzBqmlrdkJWdn0QfDhWyFNr1tmbIcRB3/6mgL9W8ViwIJUqhARZoXAucB3Hpz
Qn/atzjtz661Ybano0UXVdii0hZ5sKNS0GLkNvvuhWp7fInl3lu5ztxvCGWjkVOL
slPRHA5wN1NhxA9srJ3Ef/MaSh4O0Fy5XXvY0BrtC6OcJedSzvDZnPqBJoFy1RM0
DcqlhGAbsttH3r2HJopC3oSMK3WDIdqcMLEZwX8OmrgF8dytJyksyF+XyaFDkJXH
I1+bbqM5wxEjvrcDPJuFi9vytn8CiZvQ2GwZA9s17r2+Gsh72wKKzu4/PqQ3d8tF
uEOJIcVLYLcA4kWjxaBDnFXvzvyMGkJF4n5oDh9N3/Ojz3kE6CXHWesX3v6rMr55
zRY4BhMCMFSn1AEbs8PRbdX6N7Zyky8ttAv62rL9syxyc0OQ+8euZRPYMP4xkkLq
2tbZ4HEH0dCs+jQDLvr+Rg1nUp0sVrURhanOFpJHjlwKBwPMLPAi9OkD0bYzSxAU
GFqpMBY7Jdi0SHGoEh6aBBeZecHOCGFd2WZCj0iI8jRHEg2yM9cY2HAlh8hOYz8+
mB58xADuguGc/lNKmmqhnOz2C++rl0skP+HVaPA/vPWlYKSn999g1ti8iHNTE38F
gfSdj5sz4b27M66Qlr7NMfXUNYJT6Xo7NZ1QPW6mVLaGzqf0lglcTpTLJqWFpOai
42wVoxOnSWYF/8cOoq0lpdx7eDtV3QnWNRo6L5zy66JJRhyhOF21nKfAzpNLk4c/
BrHTOKrtsj8jMZNS3gEGk7lNp/0T80irvt+TOBP6xHQBcnvLGcThsuWDTaYZDs1i
Fhy5weM/Yg/NT8If2owZ9a04kRzDikzsco1DSZdq+ryRF0VeL/s2Evc+qNYVq+qR
+313oSwTqiHdQXcFrFPg9wBerMmSCwcCR4AMQjxQERYjwUpR6yb7VddH3pT8IhvZ
MbGmho+SeWxN0jybtY+Rk32SFj3oPy9L8REBKXsQv0BHW5SRTQtqYeWkHJXBfgXF
5P8yT/EVHjD9y/SnkM241ES3JE2DagYLa3Taii2Q9ZrRWy7ttTaFh7nG0QzAEVK4
xkdSRFNNOXbEnu3vejXUNYQUklwps4dVY7RPiNvF+gXz6m9FbhKeqPRMAb4b30+b
5MnhJeIbcBNXYQ3WURtVb936KxH9wnNmQl5yysdwOe1HV7A6FLVUb7BL2HduJc+w
mIx0e9ZBqDvnS5yAD162OiMEkWPCAIibJrigDhjtrdBoWMFwiCuC7yX4314E84x1
x+yozsn9vZfWyzDoT8Bp/l+/O5SaKWh2e7kMcDuwvoT8g2FnvjvOS76Z/4CQ7+Xc
PUELdjVv87YPvR1YfZoTtbAPBp5msBFOs1NusMGIsX8OgCq/2N9FAw4NXTeeBIX6
GcBiz8HSZG54YS1ip1siWyoLqTF06YZ6MGcg16CzuE2alvmaRtnyVKthceYw1PSO
8yb4TxTAvD2VGa3gjPBVSoGmsoiO+GfB4AIXYSrMVHtcax0X5+iNSK1BdCIMXrxk
Q9TKocb2Vt2ePNAITI7/CQ==
`protect END_PROTECTED
