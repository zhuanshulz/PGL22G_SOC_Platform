`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Cn3JN7JM9XgNQbiEk70XwWjF5gzuCBFCy23BTj6RQ1r23V308o5u740OUvpMwocd
kC1aS2g0AGcqNR7MLJ+96Z+9lq7WeaSFVOMlhptZUq90Gf4YVArowwr6kpv5vSdw
0/xX5sKxGyCV/Yene35jnKcMSqDocR+MHSuHbJibDFh1pP4J/hbBkNXMKdmSzOdV
BjroDnQgxQ9n2ghHHNykOS5Nnal9JpVTiDXL7n1EH1WVKvUjTMblAy4IST/CIRaU
eyFLXyaWtKkjTvOr+AWrHgPQUznoreY9Hzd2X/fdWWuqm4tboTlmEyaMZSEjzz1e
Tm7bmR4OQu0iIakajKSzryiXtjC1839mI4dC7G2VMwQhRf6KSZvenpZbEr3bcjfD
Rpc7fFX7PvQAqBs1Zu53oNr2g9h8CqBR+XsxnroKuq4emlxBysmHhtBKplqSQ/a0
cxQOM/8SnQnxIZ4ZRUpujsFVW//yo/w5fXoc3bwvbPeLIM1oAge3Ls2CWngL3AM8
g9Q32wu1j9TZe3hmKuinATSVQMByeMR94GR6Y2w9nWfZ/IJ44w8lVleNYyVrZ+Y8
v8nXeUzMZRG31CGWO84HqOOfJ9dJ5U9GEWEL3B/znrJ7z3ag0xuWvpDrqYKNeENR
XXPo7EAjW71RkAH5Qio4KKJ8WMPL36mmDc+kOAzhnG+HNT5gXdrdzhBrkCuLxSD4
DQkrYK6K1plInpkrX4CxoM7jgUCDGMnA2xYGRbmZI2hSh0Jhr0Bz8hjcTWKsvXzn
gjfsAFrpHGBcTQpjW4okHw==
`protect END_PROTECTED
