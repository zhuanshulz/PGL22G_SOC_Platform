`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BNffuUoRMR/DV4XF+msbayiXE+lTe5kXzMU88USOE3Z3/sPxlQVLF3PNjKdDFLF1
FLg9Hksf2hq2qmAs6oVUVeuXKx+A7rg1c+Gx6DRchn6rptWsFMEvR+vI1bMr8YLE
9qgjsuVWn1rVG7mkgBh3pGMjOzVtgSYJPvbdTr9iNM7Ug3nM9D87Kr8vxBfA+UOp
Cqloj7AtTQzVI3H8B9pxNj08aUP7bUPyYyXeoK21cFB8qa9fm6QZPGi96JceckL8
6YlCVFFI1iwKy+8m9GX10ex8F8nl7xlZvWQsDbd8crk5oWHnAREakOicgl7kumXU
R1EieiI4hsQPnGT7Xl+8UlfIkJkuOxTnj08wxrVA7sgt69z6IIgjkRyekzjVOsys
fzEA2mroyAtKY9hLy88Pczr5U0+GHcPT7PA89mhHyWALfRHgNHQ6ty9h6/VLmhos
tOP5QyWOlkGmL/BzTZ/bC51Px5Y1AlNetMeE8UzIS1AYnKv4JecIaaYSGzIo9A9O
sts6UcTN8d0l6Om0KubT9S+muHhuVgt0p2bOzDTgGhqSkeEwCOebzvWLLUIb9nel
An82JjxQmPUWVx4ad2sn4NFCQpbUrqYW2HX624TeVFzjXqy1u4m0YCzlDWLVLNes
FQkXC4xXUZ3T98Y6RcZVlVxab9RmWXaeAQ2rgzXEofJtv5JGmw2s2zZoPTCrIi5P
4t3z28wU7WZNQq0rUhGIQQimILQRD3t7go0xHOIvnQQVHta1xEDzDn1eV+Vyiecn
1fi/oJ857cqUBC/mHyhFndu5vkLqy0QLWuLx1w14B/PQdGggiAfdut4+zaJP3Ffj
xXjImeV30smdBJueO3sab4dPerHCsAvlqlRwwXxF2Psk1+c1fGX8yM14B78pj3q6
5xNWSIpEtTNUQ9vfeR6+RE50wWOcvPBKTMCWEaqG5Xy4UvWQWmRg2UyNpm8lINOK
4gzTLGBSv8p2Y2MuHC7Q+5Y0P9WNx8924CQGYNlAq6aWTNXXg2oIkA+KxWTOkdYU
FE9hMOYpSWydoVZLtfuRBHSJYhlQdOHxZbJXWQtBx2JxljhwvoY8lSS7aGmgTmh1
kBB9VeYgN6StN72RNfTs4kDyMwBaLCt7ICDmIc8kcTNq0R2x5fKsqjKrvNsvq4EI
wcpdesbjSwp1M9806sjhKlxQkDnusy+FpFlzmAv+jTLpO6/1LE2UbVJF5BVDk3yg
Xp40t2wPaflwgU4lIuVnEnmjKt28HyO7nKxhL99pB2owvcm7Fom8L51ROIFMOUlw
+DeMSWZHMpev8UBhKJ097N9WU85MtSxT8D1gnMB/oz5yChHHqro8Iwm/1e0U8XyL
eCklVmYyE7zrrCNSJIIgd5wlQmTrS6VqD+gRhNtQVyAz956XwLBTyTvvrwZPLKcq
zmEAh+J6Dj2kbE3B0nQmWNh4xMURON3AeQ8nyr3xYXzUDv3gt5YkkC2gZsYDTW7U
ewFVyVMWcXPIXFucdzRsTGjxGclaUAv0pJT5Cyb5rJZlTDU6cdoVjSLjxnEFTypv
L+qGL90Ent5H5eyg61LOTtdK1AuqTc/rTNRkAUE06McW5CyjbZhLhRlfPtPUQkq0
tuAzSYG1VZs/LC55s6EYhEU+0+tnTrZMfC001aRZh7USpLdGIFN9UBW8mSWrocCf
6Un+ToNDy/5rA95QJ07tLzbnwDA42xixtNV9Bs/uaf+D3XZvvoaGY9N5lh1BflGm
p+6ZqKKVqRwxeXgwzXyIxUeeoSugD0c3WaOCCXTauYHJdvuBoYOzKHfCZLPQJKeq
V5jZ4/sex9PaV4CFs0bilMz/xoOnyfW61EzvWLMuzv1OsqOX1IR98uL6Ivxw7Czx
J5lsdz+FSk5FG7rohLD4ilsuott+26MBx/bysfmn7kA8TazZnE7V0i9QoLkGguMK
Qq29ig4x2q5iJYuPEzkFddJR0eI7FE7KM+IRrLVGP3WOGRyEEt2F8Q9w0tflXLQe
dk2nPoaq5WEY4AJolO0cacwzkoa7Z8WGbdpmWDR8qUhhApYSm50u2Wa0cjICEbfy
ypCUuvmypjRF9mJEPslE4he0u0tlCN7Dh21eSkKJRxvJna+DGc7RTpVbr4uYbbeb
NRMXHUa0rp6Jr2Igf0rNiKMYbqmKbuszlNd/gMvxo3tb5mnCdQSU2/PW7aUH5vTn
PLkG1p76IwzqNJqVbMRpDE+6LfDEA5ikvmR1RfQQAU/pWA0HKEKu2sWrbiU+z4PH
aZdpUbBF3UGKtfdhvJatJZJFkRW0k6PUWQLKsTXgjB2o7Kyk4+xaAapZzWWRltVM
6yqMhWDlGcdI60bXxSzkf9Ey2/JFAYbNBI+QOJECDziTLG8JlbQC0PvojHmpMDeE
JUppjiLJMtU8BNoiQIYu+BEgCkVMyLJrwxGLIzURwMXmNAItnGIapX3toIkFvJgr
vfLOCatVkR2/4fKMhSrB6VSACtuTkgzDWl9iskaC2F5VRbMpvuKr8X84IKzE6pFb
vGk2MVAnZ63aUb5lHKlXWeRkNRq6tmYhHa+Ut09p2krwxm47P8eil6TNAPWpXuAg
Q0MQ2/zwAHFmecdozKLW4JPC1kmPngXcbG96Kh5C+EdeSJmlmlxtx1m4Y7+NTC40
5ZxZkDuA8WCvoXHidC7lXg==
`protect END_PROTECTED
