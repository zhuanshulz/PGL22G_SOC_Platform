`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8jBJehZ0SH6YDXQ498XOd2pNXHON3sakmf6v9MLGAeo89PJ4oh3MVhtBo4ltW4rw
/JLMhNaon3lvXQedcfzxrTvjyb115kUqQRmRgqw/UvRS2cCvtlwHjwD2tkKR6I/e
dVUPVr/s7uUtHWYu4Dfw4Z8XWx/f1XnJU5ATcauZTRFQXYe2+Wxhn2JW3jO3WVmk
ux3b4sRlrvn4wqDKMOtx3kARRRkaJc5EgcJ4UXPYIn6IqqE+lkat5mg6buRJ7Ocq
xepRInwBMvKtvnR9140X4RxahvqpDk0NUPyN2/T+BPGln7I19soSElCxcfxVFuwS
q/aTdecIbgk5ImhFs5eboOFlrYuNyukC7N5RtgiGLcTDD/ULAfxYu6Wv+82B3+gq
qMtM9K6M8MgTHNGgH7frZtfoIIaPG7kHATzgfbWiE4amEbLnp26yeJHqtKddjRzU
lD3JRVPa7NcXH3XIWk3R4XKQEbqv8kt4oplFPriDRzXsvBpiZxO3OBC7AOLEcqHI
dsncfcPHzEn8WpSmqgfNNobkHAMtcbps/lJ76dTNy/IqDFm1Ml3EYN4T8B9vN568
PEixiJpO0ersuan8I3pP1sMwWKaN795z8C91eVhmGkpPormBCITNFVsUW8H0kC6g
eAQ88VfPv193eHzwe8wwS99atTs5CULEUiBgxj4jXJ7tLH7u0Nv/6WXPD7JBOvOH
2X2rDDoi4a4LUYh33ScpitJPVEKpx2bEio57m0/V5dD7h7W4DzKTm9+0mUskEr9f
YRk/f8HmVW0GWq37YdkUTDUebEYZUFu1FAtLLFXdBWSPl+HvmuKr1i+r0A4/znfw
RxllfpI8YDIDB2lMwNjchpNACpwkinTipmYLElu04pW/wYvhDa4Y07uokgZPoHNo
vean1qBI1KZBq1ua0FsQGZJdJq8nfwQeYY3iZneo3bA+Ylp6OHgD5k1kRM+3criF
9sBYfcTZDNG2xMI9FGj2p41ZplrHhfeCaQOgOPDpql60imOD5yFIOXZhSyiKPGHJ
IXyT/iqRffVmyJmdZRdnH9khB4YFD63e4rvbR1gkndih3VgeT7pshKyG9hOJ0haB
4/a9Ezar0rjbv4fVTfOX1iOA0iqTscje/MPnfuLKOB1ksJIGT8lhSdYNdgVq2udY
ZdDsE8OQdh3BV4+sVxPOS2CmgrvgcWl4I/mDxqOvjjz9k7+z6OltrrXReNfxMlI5
`protect END_PROTECTED
