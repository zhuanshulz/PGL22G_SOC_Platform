`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RbZWInFmNLHBWR9pUwGtoqggewco33MUCzSmY3Nj3RfryoTVaPgk3FyE3f+9RhvE
paCFE1jy/VrAmynUnNuKAvH4AmPzx7MH80T7HgqKCAVEGEtRtXXBVbKQ/U2Ok5s4
9iYshpue89abjR5XtoamlbZID8m4yE/Rky8vz9fCrg7dwhtvpXJcypYOsum+hfOs
HkQmC7Wvlq5byiuAJVCBSPUiAMyRvkZL2zBExSCs3WAExALFU5O1aX7fUAfMBFBS
zYzXeXyhJWoEuzLJEwEoaxS6fV8Rt8HQLY6Wtz99kq4ZcC7KTdcm65cep+e6HiB7
1NNcU3iEaVf0/hm1pH6Sa750bdhiIqah0S8ONt8c8WqQoJla9GSoERG7VKJeDj0z
gqHnMgKr1qh34AVJiTHSo+ekCrVhcB3bIr5Pr55FM+PQPRm+4m4WDp0kowbf+0Y2
Cku4ZvYbFjJD5c4ivsRbBzYTuJ1fERZ0A9dImyWfZZRWPjB1e+sZW6pNzPUglgj0
bWOuUVoprkcIQQ1clTvaUEzq60Oy4h0thJvurjwjKG+LR9tFMrt6qQHxU6JuKVrm
pioHbe3GOnVl8TiXFM5hF5yc0XU2LaaTNugbHT81CH8eZQZ/sW3igDs9P5UbPjzG
bvO7qA3ifjg8xw4YkKxYKIjF2JaSHY1IgNIRGdf0GArMhGuE93KUkVccFIGs673q
/mys5FMrDIx4vyIGKm5a9BI73JJqwtrmu4iP8gjGcOOC+zijlhRp3uMA15D1I/4o
ty5c7Kdi5p1wCYisB0jXOim6zK3yrHgpLugYXvqJRq/eh40oSZJHN6r9Izt1uLJn
a04eCLwZ8gvYMAIu5EKVYe8SCPeJiAzppZA66o+nVjL5aOG3VG02Yl1aEYrrLKL5
a1uwATBTDGRpOTK04IV94NWBpiHWMH0XkGDIfJCTNBHxZxH4RlLp2cGy6WNdS1Dq
Mn8Vbyz4PJR9j61btC8k+f6gNFXoYLs+k+CUhrVeOI/2xQoQ/p8UO7saVapQxIvZ
h28nIt7kYY0wQXsH2Ybw6o32A4lE6wKgmijpFQKfbiTmgk5kjTpXHV/9qpzb0S5r
d9mXZLzZtcr9P00pE/etbcnmAzbXvhnUOMHLasB6zX3LDwLHwxPo6zqJrWmpWRZp
b+DpQinGBTMwT9UkSaxOrqX8XrbKGro1nixrisiLoRD0grJ0UIpCyBkIbAhsPvj1
XgxAtuJvnnEn/xz3mepYGQ==
`protect END_PROTECTED
