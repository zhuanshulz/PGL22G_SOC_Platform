`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FtCGEKmit6GdULPpwp4qFSG6BZTkXVZ3p1O+S8cMpLL+tmVBrjKssMMBzgCcWrIL
XhtJsGOW3izaywiSLpbgtl7OIf6vXWJcvUuMetAfbDlerB19T1lkd1lUxMaFZ6X8
4mnjaLyOAuDR86pRSkjdESGme8+cJX6vaMM6LEHdbYOpP2SA4T/8NN5C+4jZuFLU
Is9hafeA9uEvhf7ToW4s23EeW4VrcDDVuGB9IHknmPFpIyU4VjZq5vzPB9xYAJti
OcEJ1TUYGmMxKT+WOuaSJuzmd+3BODFJeHuuZIgZoHu3loduqrcy1xJydXTAL6rp
CGmay6RiXQWEiGWl3ptwNe5uPoGNHk/WTI5K/0DFt+Ox10qpgQiOkZ70F7Quvmuf
JWokvdn5g1j9Usa4+vmdcxvgUFXg8dEYJjMTlxikXrVK2OcTsCOzI48n5vY8WcRH
3MBNG4tY0ikE17DnlUzPaG4lzDJUijAcBI06Q24bor39UO6Q3ZSFMnnxihDcL+jP
o2XJefBf3UNUPEn3hhrPyITiC4ZEf5aYdE6HR3ZFh+bK2q+RiJzMkfl5tLSd9pHU
w9xaozT/p0x1HW6dr/lxkFHOAH8IkuXekjxNxnN3aAfVTnGwgXpvuQlzTszpJM/E
s1O1wU+ab/OnBA74iWWNIhvtHphRMpakWmeCdjYfrkvVvB5BxAF18t0oCw3brcOn
Rv1G/TLKZRJDD1VloCvu1uyNs5tgR7oTQuSgrn4jZH/4DuxheAtIR4przpc2SV5P
3X0jibGf2+H5CR8bo17htPa4pEgBJHW9JhAGjQrAim874EMmeDaUyNyGlMGkrynp
TMUOVxcVfatySCxEW0G7aQw3PG0Rwu5oZ6q8zwA6fNJ1Bsprwxcl5lKzrFBU8qyR
eQJHqarT3xi21odLL4YQEb3Xq+B51VLnkHMZhTBFb/i/bE8UkzmQuqiWSteTp8/G
mawgZym3ErfpXWf3q8og/3JAN6aOvLfeSg54MOfU91IRjDDgxxWIDqedjle4je2C
5h0EHkJyp2K0zGqN4tXdpIhE82Ah7nzXO5BwvGfUwmc+VAWLYTvcZKdHm+ObCavo
mI40WmcdQwMlTl6o/Yd7yYd/Zkadl9iFWcqMeTQopdd6XdlCnDkXJUh3B8XPemO7
yZml4AvCrRi3kEzya+j7Vw==
`protect END_PROTECTED
