`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7WRwBUPFic0W+m5L6jJQVSrD9kOU2eJ8LpthxN3i0i5BscM0hGxU15w6b5lvVaRx
1EMSwCLl/Uy0CZiEnvGUxIAY3CX2ckg3y2Hh+HsgoIea48+s2WTY9l4ODGgTf3Ns
PxH7/+TldqKq6Hi8Z5F56hUJgUQ0BNkYmwn+4ssRVuqP9kbBM4UlQawa5hWyyYVJ
25Ol8dmyZT45MK/idUdZasrGx2Dlo1nrxf76i9y7wtBSkzh+9k0sA+XFvRhHSrEt
Apjw50r7tqzbFMGuVZi+lMuPMRAZgdFe9CM1m3kR7YLSpoR3z31rFjsFC/Coghn8
vyDBSuM8NwHMonnw+uW7PTdX5I5pVFdlJLqSgiFKhg50ZPRWOMLQgaw62zScIHo6
8PLUEzOCeK/qovnndmFx1MfkItA3KJjg/a7RgAqHeAu3OnkTskchL6+ZBulrJw/Q
MUey7L0YfLtqwZoiADEvM/+iNNamiXnhj8lw2csxn311TffTPHb6YWzrjMao5qHe
vQS9vTPVWpQRBHwhhJIia9/4KJlPhjVVL+EKC9vMQ3Nq8GLVP7GwzIH7i/oUeu3S
3nLagAs6swXbxmIDxwlUD6fKij07sardXh97ZEUFd/eJraeDoSsDVQiuJOF/9UqS
ibbb+IPA5+HdfN6o7Mng0kn0JggFDQ5e8pDem+eoGNG/9VXLR5NKvvbJhcdM3OpM
DJpmWfl7/GB7O1hKg55eTKRjxiniICC4yAEo1zXeqZsfxGjWoso768ZRJDpRLL70
TaJOIHPEsdI+8bUepE4QZL+3WGu0XIQmt7c5Ax8ZwBZxGXMWpWLPIbVgpM2w2m21
YZOLwYv6anxg4BRsaxDMWGWOiDiRsPsQmQn41GRWBn+L7dgAuLF7htGzNZ8nIRoL
gEF9clSB7N0fd4rMynBICptsWijsBM82PjoTsPehd9ZaJZz3a7wMzx8I6VDwRXuU
dU7FYulOMazRGEh9oc5yvuJRpFAoBJvq8VmWMdQLGwI8KKktsMBlCwRNcs1g0iiT
ocSQEkWuMBfhZzkJovukxzVMVtIcZZUZQHQrQb+ILGztm80pgEDqYL37t8GWkIlx
iChLgXTT+8ChgtWainGzfYJMsSceX+M9/XCj89IVebhXSZwOxJciYQa+304jiruy
M2jkdjUq/93KH6RSac0u0TIp2S2w4ztTZZAN2uMXyO04OK4moypno1rzifkAA8/D
D+QgPn/inrwqH70cHjYoMNPgDolhc+U9pHgwmCTQnS5bGH47F1o3BBtDJX688vmJ
tiR6ZuO7yJyf/ezTIDkCEG5kiptAeGyO2JceQUPDxKbwRxwzbXIZ88eWv3vyoz/r
y0wmqFf1o1Iy6c5zeIJhkPSZJAC6humVwUJkQY9nD6lk9TofmW20S03SOIXvOLv4
7sKrwWFgwgeCrGVLqlh6ei841WRfgF1yC0gaks6ilTGYStpWCvnGhqzK3Nr4Wc0e
8RkA/k/SO1Ql8GN4yJmtuUbksnPVGVNN7EwvTxbm0tKpSwVxPqLx6PXkVYkta9Qj
bhtNIT+DLBS9F8WHRNqcItrVeysIptEgD+uSJlcYRKG25QNwe/y2HZR2bLbgcZmr
/nNhzzZlfiLX0xTsFoPXKRkI7OiztGkNKM0zrIV4pxZXPpJ1JCl/J/BWFCHnGfml
3fJb/VYmCgVCD4+CKxY+PkFIOMfnS4aUKTgNatgzt8NGvpTi9x9D2LcgZZ15h6Ga
WKYyjO7iQXpdGEuRt9WxYzl2FAjQkdLiqhDeGQByPusrSljwoUQaP6QVtGhGyIEF
hfpOxNlzBOqIV0cuHnc4PAly2OByUeCa7dzeHQ9kWj3znVoduf70Ghm2pBGTgVQ1
weTuOMUsHCvmQr3Wn9q1c1swpmLOa4pRPdUKnkT0cP5ps85jkMAsz08RVr3qwkSw
VwhVfVlbZN9/sEp0FwO9Qec62yEZWbtSFoK6YWigMVLH6IQMuluGb4nKnocVXVOP
sXGjs5YiPSPxQ8Dpvw9iLKHQ79TOy/n2C9VWKcPBRcqv+PLoia0S9Ao/mRku5dD+
BtQzxFboAXJkWz3kwPy5xrZeMtyc+LZgCda7uYo0Q//o8TW4dYN+dy1ZAHrhGfGi
updQQHTpYSJg6ELWGmvJ8h3e9kmMkU3lL/yeS3wo+hO67CtoHDoflAQ6r490MOQF
w0cqDwQDyanMBN2q5vacxRhj1cDK3/ThRtBi2Zi/Xcb+iuO5LgQAyn9zb47NnRy7
6O6wYEf5eM4bUJDzXfYvm7baVYSpPPQ6ODG/gffIdlhW/t/voaFz8C0wq7fH1H4s
eRkRkBUziiT7Tl8uVQpH0B32ifvym+BU3dwkb9G54TqsrWvdO5QeYtojkz09f4+d
umgD4ksa5L6bCXbMMiAkNXK8vyXHvWeCj1FkcWUhbz5UEubIFHuHsg7jJ+/qmJic
BwXNq2Ez9QmV47S7A6NpZAilfQRz+TxPEnVdRZEJFSv2nkE1tC71Ol1d6ZCQDw/9
c4GAdGLD3h8UWdPc1/YLFpvwmInkr+76IqfDV7SNp+jvj1tvE77e5tL2WtA33yLH
aqNGDrNM1Nehvqy9t4mPqKuAnSkZ185C0hE6ZGe7+vq8+XnshpAEQCdkXAoX6Gvy
TnBBqSlQ6DgCp770pY3QctxGm3HLKSvHvGHHZA4lc9+YvLzT71/Zl1d18x+UWiHm
7bjfIOKwvi63oPq6LQCOS8lC6bd55qmvibdm0+kic34Tnlov0UFFyVJmDoanK857
uFbqJo4j5hzaefudA6yGMQY/gTBhjwtf0+EySEZMDq32kWut3LYaYwoB1qVpz9B0
xQ5nG+J6ev281t/sKXXHpOCJQCI7giPdVgBp0rtnX0+7UD+YUDLs1lUwqWj7XE+t
g6Sy6nk+tgkcMUThq0uxVb4zUMOxVirU8TesawLMCZE/SWVJ4+YQocerqMD37O96
IeyIqxzP314V605J0rN8iJyMkYcesd9cXVV6ksiBuAqrn4+jVXvsdrlBOV59FD4/
DRuSWu0OdaTqfLsFOKtYSEFqRmg88fmbt8el4jyPWFrRuLGnt0EBaCQqqHcdKHyY
M/7k5ypL9DKrx5JZQwOYch8Z32nopje1ISIfAnVWhYAVFYs5cJEvx0ULARCqfkV5
AO79qYl/nGCp/eQ8c5n+VHrt52/aEB3AYHEEO4+gZf1eZbbIFTlb+4Z7hChgCY5o
Af8ME/MXKQUieJ9PnLhxYUFZqmNZU7s4b3wxAbfDq0rd5SgHhLOW2e/NrYE2hUjm
gfq1KPgmkpwAiCQS45k9BcU/xyhqmPINERb0hnTiJjH7YRf0fqyCriHc/C7tTy7e
aDZYjGHmDuwABytxS8EPOg==
`protect END_PROTECTED
