`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c0rpPhZtluLpCE0+/iHXlq7MeyJBiWFVnNUkPf6F8/zsBTHRadCjYDCy/ZYCK0Bc
AdVAX4iXlIKSDlkIUdAVF9qvXfSk7o5gCX2hVmBfxhCXm5MJcaRumFqPe+If2LYz
mKpz2Euf8RVU6dche85CiEsNZu+zXOcma3aKd//5Hep9rCa1GtnSFMUuD1C6eS6l
t7FJBg41m5obyaimba6q7nnd+9bgaHHHlJPN7S5ClIQIOzIDspvEmvZH4WJr6gvk
x847frOlF68+aMtHmGGmJeDq947YCs4cq3Ru1ZvWJxJygBIU7LgKUFxc8zrn9Oqm
prT8quAv4XgXPMrFF92DD+ti6X4hpAwI4omIlIyU0Q95lD0qi7q+7jyduae/20YT
n/rEkUNHKY2bppUQyWz7iFWzg6R4AaFHrikSun6qnuyEOI3r0cfuR4B6jK3Ie04Z
smPrigXa/wmcl6aiO5FxzDl30O2WDBnUCXJ6L+ZIsKbwFx0z4tw9eg2Ko3TqNqiV
Nq8No6uCLVVpMtkN+OGB0zuEekf39W9PbYT1EE60jqBMWJ6UUh1IJKu7yaukafJn
`protect END_PROTECTED
