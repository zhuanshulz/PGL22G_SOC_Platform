`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eL30dH/AHGRIAi7LJprX/090xcKrbZNhz6bHpboJ6Yi6BB2g7/s44Kk5ylD+OcSs
Vaj71ekn7Yl0J4T0jdobs+elwUy4evbrzhi08xvIjlNbQbvv+zBD3j1Nv3pdJpna
kADXce1tu0FQQFzgIc2PgZaFJPwzOrp6WfvBDhpZsmZi21/29XgeIOPtqoYTcYYf
FIEoe8sNCJ07w4u2SUgu++UA+yrLV3xXHacLVck8gs4AEP8hRXjfgN2q0ICljdIJ
6StqVr2ASoV6fFfzcMMrLX2bxlyyrEeTQxiBEn01Znm9B49WtIY24GadjJycsajd
McLmM1c+P0geovZewll6Mr/n7VM/Clng72ernxHdbUpSUV0Z8hQ0DLV0390Nr3hS
gN3CfyZMAX1nXvLC2+ESRpqjcezwUNg4MPu07UkduiluZ2R/FSLIPT2Ayndc2ewU
PssYleyjSTiTcS10Sdr6uudPSXXgca1d1PwCSZY0k+Cg7/RJUEsHxvaZSk5VbZ2V
Wd60xXH6L3MNdiSjprB6FAdF2Pt1mStQ55uCVJZbRMziPqw2UdZZEFp8DRj48DEa
p2rgDffQIkhCq4ZvJMOEh4xtg060SkmT2kbmHXutzvnDt1gFabVOsa0fA89mL/6D
ak6K7Z63YE+DgB2OhGSywT11MuSOUqYKxwjjU0nPWxk+oKC4g7FwnAulI+hEvwD/
eqV8OniZUKCWCLhrxKRHAfdJW1BXH6bhZah+U+8gafFEHnnxHCHnJXfMO9kP/r3v
gM4LNtBC2ilnvY1FMd8zmuiaq6ZGY/Ackvmhq//py3FUruqbIHyzE434hmtSGsyw
F0bZpNEz1h2l7a9O253XDGGttbX1QZBLeT/pKBnQ6EFal4525VcdercHnS+Oj1XA
apjP1C/tvPS8LlbJ9hW7/mNCwvB/NsPIdrUSn3MzLsAjSszSQQb7lr/cHo4Ikoau
AEc+/nn+AZ48e7HXtlbxEEFX1H251T8fxIw5rSl0foGIRUzzctWEIq25MiFeUzyo
0j/9ZLb7mQRYVf29Hn/9Dpkb9oVEHi77CmELVq+A7uh+mKW/aeWB0125jCRUb93O
YqOqz5+LTqXlI6jcAXE/uvUEW0AD2YbYpz5SgEBs+hPMT+a/YW7n4QPrFmP4Q+WG
RAPsu6kjpaS76t/c6CHdtJKH1m8ltpC4nm5vgQ6A2ugyVRwFWHipWeHXvtUbLLu+
0YSoXzQ5N7CximjXwq9FTPM+UYMWImVXVmcf1CLN2owmYcuRqOFa2LWkymGzFvbQ
7hr+DGswSr7zw0VJA5d/t+zdqG0FgSOvxInbUFL8P68vN4EW49F7TBR6EC/3f5v3
lnYBrojunJPoA4a0TyV6XcgTPVu8ZBzZb0rnnu94cOLFAMHMddWHoYFmotnDbiFd
fJCHYMCtEDvqkf/XZ60/hkycndGdT5DWd9JE1VmDQ5XpHpGxuNnQSilbV3342N2z
IsJoJZ9kdkhRF6AL9QE6ynz+pdquZmLXot2S/s4WBYH0sReOhpV7E4WLne7UyoqQ
HSipbgsMkvbxxLxESECLL6tqkj78ZmMZJPEGPjHKWbCqNzpwh3MHI+5oa4iY9q+K
P/qhDlHrNcBuS9eMmDFL3QjejBFbLve7T7ceezXsssl8QrB72G0GmN5G+1pbwmid
DeXkf3tJQqXKAY+20/Egye3lB7LgsmDTpJ9DahT0/CSGwYABLklQv5NcC4aA7x9b
K5gGoNeeFqythRP0DpCHoIIe42JxTs9AUkgslkTexhkrj2wP5TUFh4INplRKpKcz
lIeYxT46wBrBf3I+z9vm0mgMHy29THEAxX+jhMauDy61ustYbucxSwX7C/8HshjV
2PpZ4pTRsv6qB/rGfsPRyWxafk1/wk9DL/UIr9rh9An0zWi76yycGHjh+2YChjBF
9srQPO3wuCV3eB8BKI35rdC5jJ//VmcFW9XSSry+TsZj+Q7pZEnJn6PbPg5V3Oqj
+IlknbegbSCTYCxX2o3mrBP8ZoMG9U9dKwTRKfpIeOkpAHASNIgx3r+gZe9K8Hm5
G9JawM4Bwe0e36rfFudirGIso4RdOJvoZCj2gmd/tmgef+Ec2hlNPPIYUgB3fLrN
NB9xeK+fcCZbbG43Zy55HFuF4EP27chxIyKJjF5WXJIqygduAHJkp6zccW+4yxDZ
ko2G38NLSyrcmxF03nVZzWSUuInChgYIra9U9SpQ1mLFs1n7MXKR1RcRnQZRr6RN
UZSv1IRLxlXEl/3DDha/UfnidTN9DjFyLNHpsS6r2Na+sTHmkW8ZMuoQ+KVYUw1m
hOzqNF6TExMvqSr+7xlTXa2OPPgyNfcoUWQ8erosFVCpmWTWoytmgk6Pf42xo/uv
3+M/VOt5JvM2v1mVzdCu5enaJDJsSVftTkU6AaRtBhp5rVTHOQt4thVhC2Qsgdjp
8F1SH9fKJWgYvIckg5vdLncssm9rC7jEbDBKUh24mqd7pUsvzL3ppcnJv64QIS6z
LzxK/iQhCYI0hQs9Ul97zQjfMG+Gcd/PX2/3UUi2BzXvH3Ht1xRY0ZQX/kB9jQNo
M8mUik7ISLNQCcg3/PQXT7Stgk3DFR493z2r3F6Frai4/9Ffxa3hHkH/b10KDwFR
54g89PLS82f/thS5g43h22jjjW5axXuJiKAtWGE9VMfAHk9AtcElVKTZ9MYRgztd
elqhcKcOOUwu2gvmnE7DkMmmnwjAXEk4GIFFYav64jfq9ypQIVB/wUK0ZHfnKNtm
Od7fkJhjoH9RDKpmq4H7+qQw8T3qI2r055+2p/xcj1L9LAd9K7SdRo7Y4O/ASlKG
FMH9UNPMcByrmS4ZKFoJK+QrOz6Lic1oaBGWF9SuQ+YtQTRd3KFiw4YzBrRSonpW
l8ixuQhk24CHCnmT/LiNn9XIDH9QMGRRqO2loq5CPiQs7qnChaBTfdpecZeYIXMJ
SKet9287QIGF72NrNrpFLv0B06DgGr6XDBi5U77DFD+z4RXIBA6yX9Kk1rFBRReM
aCeEw2JBYP9xhOmI4hpF41ZPUM9gphlsw5eogjAm5EjjbQL4LBNjYIbdP/B8xoqu
7RZOEPaZ2aq6rL+rUbPCm6JTJ8Mv9M46dBQgNK1ICmvc/TwEzgDTGQC7Wz4+EBdu
AZta+ydnXeXntRYvzvnFCSJtl9tIp2qA8iznFCJx+sxVT6WhTOncaAd0m382AWaG
kchiwu79CxqooClWAEGkFtz9GaqqrG2pd3aUv1VyZu8zjCUBC06Yae+enr2cSLGe
1E2Uq0wfO5jzqtwEf3Zt85dLuYhUMi+TUe6dmNX8yLHX1gT//RZNFG7kYHN5CI3R
XEeKqlt2a2FvUD4Z6RAdyoVW2RAuifAOeKFE/8ZNZK26S33Ql9fJ4KBlhD1kpT53
jFns3Zhk8rYgjo43ueH/+KlSI7f1QEqCHe+VN+Nu6lCKkNUBq7bP3HOR8U5ZncrM
PvOmBiNwZ2rC2iCuaQyj83wvqnHYoXxwr65QDy4S/yMN0YUgEgmSKf0YvGqR9Ttr
djSKoR9+KQn44DmieKYHMoV9LZnLF2aHmchLl1MxEKMAo2j3g0HaywCXh4hvc6fX
5lKfjn4wR0SW8VA3v2Y30RUm21CMU8ewzaZp5hitA5F402uhr010GkXsPUj31tQg
AmWTHdKVjfN85y1W/LL4UUDEyjpr9oj4TsUa/izJA7RjbNE3ZWCKPmIDWMiJeAop
ZeDIz6dDr85QNpWoyaJ6USYml941/Z01J4zd6Y6SmxOnvm/KuJCGrWwjm8EEi+Sp
b6OovV2YTDxWPXl2vAHGrCU1YImmb68lABNKTKHckVKNm37py9eAt9ON1dWGuNMk
QkNWn8+8nulfWwHb8qywMfj6l968ozYQxh5ZAzlJRbXZChC+T7zc+N9slpufnz36
MgMrHvPJOA4RQVfVc9fHcFtt1yUDW+SodqHjk627gNasxR0F1w+8W98l6tqRv6kw
VmSLxj3ee2rlim/bRoGuwZ+GkYeKgpMi9k0ONHmSspYdTzNrrgUMAWisR9CpwCuN
j3o/2dpWV5f5tOmKG3Q1LUtoT3Bkz/H8CB4ARh/bzxSeY+BFGyzttpvFbyY0/aY6
WO2/dkWEm1pMxNvZoqOyZ+uZEC4QvQkTl1cSqB/aouVfnEdTE979jQBWomeh+WbW
kQ3SD22mP+j8wfCbFrO9s7PPsQ5b9KeHet0lKmOuVm+xN2e5vkB4K0MWplaMloWt
xOKDo13BK3wu/L1PPRevZgmOL6q9BxmfPAN329m7WtLia/c6CYmjvqXz7goHBRm7
17V4tM5EkmghgB7lHdJOExdt0/+kSw5Z9TCYd1P7kdAZfkZ3txdMuYcZTdIYRL5w
kdZ29tEkqAwRXwEKquZnnpaqHOXDRiaDCnKnuRlknxqFGkVJdkYCT/ag8sMyA7yZ
3j29Zr3j7GswXIwyyGHggRvTGgWwFQ655j0VNGaQTkwEj64HU8bC/NXZ4aXTgsI0
oK8pxwSYVWJPFsDbhqJPvqHEo6AZAAhBl3M8hCbnXW0S4qPdb0AItTVjpN4po5W0
700galTN0rGnQgHy0wT7px1TpH5urVRH7UvJJ/qvD1QFZUEIqaJ92UOFH1vkan1c
WOj8GBbZb9cS9KTFua8jbqxrzWB+0XHY7n3ZTu7efJLosTT4/RnQM/3+8g2iOdYP
w7UoqYZDlKR7g4enmxoLxhvARmgFyVC/BK9If2qXGUSqQ7wDIUEzHNjL0ldI23n5
eUYepB9g04iWSzsf3eBLAyS+a/0dRVCIRmRfildcd75GY6QJ87wlL0VN7dBNaHtu
DIYTra5cowQEfPVv0hU213sB9PYvKbKqitF5RbANUyX8oO3St58YzhjdyJnXUBSE
y+qXzTRWXLh3TQSF9ISzFG3ysov40VBDV38R4JN16f7FNEceTWg/9X2TE/PkvGDi
ZOsr5EKQUa1aASqaUkYlOC1jJrjpClt97Sfvj2k4cLWUyfoVbS4aXpnMBgPdaKQW
sGFe8A5pkj12R80sVneWCLrvwlVlxQRGpGIBoVvq0TtknxU/DGD1Xpc5dX74SmMs
SQXlmEuRaPMV5AJTp17JbQf2CFXsx/ZdLvxR0C4geyOuyM5UvzwCIjtO02blXa0v
KREFcp5hgYf+gPYmFiiUgY52lKoOhnNfbUSvFMl8VS2FvQOV/mxK0fIOlniZdLFe
J0BNxEMcvuqZVtvC0YN7NussmOMg/91bVM4WRK5w90RvmllSmu1NOg29twpUofyg
v/7pgk3HBg8TKJlkuKZ8QUeIKamHUoxSs/49nFhfarzyTZq6k6bSvBqRBQWWJoci
gJ/R4vUpLDjY/nqyGeZESt3k5/UBGiAxDhADLSXC3509M4QiP35oPz26CcRBOLKh
yI+ZV4IF9LPTxgIMKiopQhs2skA76xCutxGrEjgVp0vwlIJwfxJkel72/piburhf
YO3NzNW7bc+aQWR5o8A8P3JnEy1m50+F7r5wfSRn1i8ddQA7eD3/cVA+yyAbcosH
Bh0cU9DDagUygNiXcxZepI5Oo3q1zVfs1B3POo6Z/rKBPH87Pmm9cZtc19hqUaDU
DVS+lno/3cSP8+XokD+7TzKqwJTWJZHV+0bHSfdLUPQE4MJmgItiD+UjE+JCv/Pq
N+dOL+HbP6NBvgJNOInrLuZHvtTZQnOFoF88q+zBIPJ9ErMpAkYCcY5Hg3QmIBtp
8M0RTxI0fYKez/JRVaOuyzkfEbQAQdVP6K+ieLBFTg7yl0LKQn5pELmID4yEn4sT
twoyiSgzj8K55fMAriVwjVtyYAApobeBnBEyxi0TFuFZIpbGtvXPOorYk5+6wfb4
1LpSBkbOpj2U6VzdBeM7VSMBrM7xJ+TsmyMkc6iKNBK9pSnQjRHUEGUzxZR/v2LS
ZaPmZT/Zv5zkk9tKJ5x7sKUZTe6n9qYMs8qoQukVJed6L+Xp++hdgljd0n1s/0J3
UjdVCa6afIWC5pDY6H2PVzx8NwrFyK2TZnabGZ6eoy4KIRKueAjecM2H1umjsxsV
YDD9C7bmaWL75ChOB3XNxOtSfrRsdnZyIYnbEFBSnmYG1sLAS8RLdDvnx3TD1Laq
9QerdWNoaYKHnU/JZtvaLGY/YHG7DowU/5OT1muIniMWNdgn8E0IfF5bPAJal6GP
tShFi9s6WEfvY/f+OR6hVnb+9cazmCiLV54sxTtgxqLhgl6FnaOfSU8u+/njkHow
9hItiElhP4SowZl9etsPGqheZO5x37E9/FmL4aOVlFDggwu87LY6k68zuHQGUto6
Uw0vbgZEoygWcUxV1eTM6xuOFKSmATN6/tmD1ZpLTpASzoG+TTyDCwWSMT0iUCXL
VGuQgeAWLCtWz4tt7PrcSfkiusdqQeADB/RFzuznuY1GFg6I9N9bmTs2TQEx9K5m
2m/I7NoU3oAxl3uzeda6M0M9w5RrahhI/7tXn2sALC6DoYYysQt398n3k2L0dqd5
r6SnkBnKtkreoZpcMOQXvm+xHj+C0VRXqDuporkzPELeBYQnlG+rNEVK1rGBAJj3
uMn9XjgRnR5t4e+PwdDl5M8B3SXAxV+d9heD074OEWTGtzGbuRIx3/EaCFvT8Qf8
7KrSiz2ZciQjnF1MPMF8n3O3Tud2VLOZfOd/AfOKJMgpuHoyGOB/ffNiOkdO8c93
32tB9MP45SldC2o/gtOlYuYvqZLHm3hDP+Uf0j86fvy28NCUlYlxGbB5f8xRLqdQ
Wo7GlKFUabVhPLDyV0maIzwjbrbscCJhmOUR3USCQaW3AoOBOyQJXirLHGhDaWOa
Re72hWhCtfyZfN/KTdnreHc+QwIJX6VvjJWeCFZV4kauMs/RlZXl6qGrI5X/Q6bg
fXwqSIlFnqLjGls7dKzwSsAh3Zyq3WsQHMaGRaKrJZYSGM6TwM7TyTuzTv1tshGM
90ck9P3Ysj60nasVCO07QaayTlsNkvMxgK1SacrQfHE+6HEP25wjMYmR+omzjO+W
vZNQQqf88vS1XCWgih63CdwTzxsot1gvVKoE8TYG+kkxCXHsshmU41+KdmgsKHJR
hGkrIKerI7q+lXpnqKUTfWyT0k+6zlTjhTmr/Xtlw75gOeBCCscz33qFRF/rymLc
OP7krDC2btTJXMRxeLmZVQKLY6Bg9s/Ks4Y1dc1K53bCfFFLGsNo2JQtrR/I8GW+
5gJDKsn5Pme7Cs25pIdWWAkr0Kv0lG1NlYdYACVrFWAxTxbfEnbzBqcA4GRwDnqW
3v+N/LN0Gze3T0fe+GArCXhPiOpIspRu9RCvVHz9RcMxZVCV6XNV4lTPgXJmldmQ
mHvIlNI6fjhkDHhVnlth45US8vfEeUmwenw6gf/5rc/owGLSPJ5xnncEYpWwfe+J
2/3v1BsEZzPx7yE1s9LK/qna9XZovIvncGWWzALpEKGm9aHm4FAB2N1wY8u9oUpV
cPUvT86VvmhPl34KmfoGYoO6nLMrXJvQU+vzp8UQdDu2ZoaPGVjq+vSSCg5I4afO
vIZMirMEdFCRrxL43dzhl3bO1ovGElIM/mcvwkiV/vN/7e8cZ2gXYBqDi7EItqvb
+S4H73CQLjFOxsRm12IzmfhxpNXVggEDD63TC/krNQZFIc8sqHVHxDLcNUWhVfPl
aUg2HaVJWhL7H7SmrYahfpY5gLOkQI82YiY0JFgcSCMuVlDP3L5yRwH/8Kr4Sb+O
35w/Zx3yAr62JYlkMA6+P/5mWDu9hfV5yHclPavwwpuEV6ZO7WgrdtoAkzrgbZ7O
iAzbbuPaMl7OW+7RI0EL2VXxCrpIiFAlu4S3/rbkMfNJ1ZJqwZB6ZMEVFvr6CiiC
9fmdQAjtbeOo3W3xxs918sh2e+A9cWDOGx9pbgmijXHfd8L2ruleS22krJdExYxM
5eIryVju+nvxpYZX896pNJ4owLY6qZNzW78YmzFas+ucz0DKZacdOnJ+n+zUtou/
OaPrRcH28goFuly8tMv+yaw1Vk1zH/t2aHJhNfMI6Rxd9v7koMmN/sKR8KcZFpAx
sKHZBCD9FFXTWke4P2oSeTEkt1PFHlFx7EaozxfpD1sXgzt2OUgy9TBPmpMp+0Z7
+GfuS+GoljFEfKV411G0BxmykPP5JgUbDHOVafZFTgBKyJ+c/S7HaIvBnHVz8RS9
FyYyxJeGH/1brDcA0ZpMLR6MsHCOKVQjxe5CyaIQkcetP4xwO6xeqvmGFSFQfRnY
cOAxM3qbMlYH7dPIIDFRkVyBnB3gyKRex5DbvRKP14aOfA4CgIdTKfZaonsGU/gI
PxcafNu2GBPt5UrOxwZcSR2EBnR5bRRSXwifaAbqsuH+EMVXc/nuFHMhTKGqVJS3
pgQrWJgpCfxLBWXnfSPstg3yZu1A8KrHSnfctw99Cg/ciPGXgdK8esxAPxhV8a+U
O3rPLnX4r7Kw+TYtdFRi0mRgFCNJdqYCM0pPMCtwsCYq+l28OTnrppmx3MyoswR7
W1jI0VZWVtJYHtB9206pbsi8YI7oNOjtp+o7KATNOpCtqYRDvcC4HtB7KlCXEt2e
IGlHhD/PxeWwfSYNlBlPvkVXutgCVuhTTOhwfjyE3cthRia5vYb1HxhdtAPcFv59
p5D5MINU/vNOTb2aPmaCPh3pxQTN46RGhcE3FfzKBoZvC/n4ekphgIRuA6GLCp2v
uSj8Dzoq/mwTpDB99k4PfZ2ipgPQjLZ7166/zDr5INWSgP4DmDrsTgVOYb+mLUo3
smWkPAW6rN6coUtqn/fzYochByaFKBlrJy+X3SwR3qcRnfJq9NImUn0omVjmiS3A
HjBNbnMEPyppFiKiT41VFdPjfBNYIgq3pKLYWFtYjO96VQG5JInv4Y4k6EnAjGT8
WdoyylmjrvGrUsJ2YPM/HhnZ53r30BSWiMQtEL13RtZBpWrC8VrwNE5wCF8yYYEM
Z26YP5MFKZCBApKLfmRJ2Ciq3PIALoRmVCltJMPABxfobGRwkpEMJdzyPaHTAEWB
6d7skk0LAgMhPWdmYnWTJ9jPMm/loWQndi20qFravKA2JQEQO9P5kcWNp+dj2SpC
+FXOVYmvMwtahI6Ll1EGoBUoViDXDvM+zoxpQzI/aWVi1L6/bzYmRcZAP5fQColc
yLEaENqRQHbov82q3pNzbjJgkUsRokdN8MSjCZhU4gM4cmrrzlfNPoSuS5k7LqfM
/u4rjbvgNoePEswAWhTRiqfmRFGgSxMNq2B875LDlBrD5JRku0zfo8dnUCYNESjv
x7YeZ9Pe/8MiIwCSLO7GdNC+V325R4WYImJfJZNmNMEXXgHacWmdN3lYSfFCYwpw
U84fijlbCTR+8St/JxA9Wk8l3UidNfK9qQN4Bl27r3NORB+pbZj0YhfqYhGSPUW+
vlXdEEPLDi+IyRriLQ+/69PuE7BFE6OnBuwj1YxuiAhoftKkK0O0aWk/vsaQpjyV
fXIMMJ2njB6Iaje8h/YMlrO9+x/LHif6i3UEmnGP2mJMqf0LAxJQh1OrHXAcy5pc
iGA4fVRLswmrcyaE0aDI4Ag4WMiyUaAmrE5Pj7zgzqwlmEqTBBiFNM9Zr5C2vUeS
Fs5/6veNXW86FAYTWkZIMRJRdCl4fce12euwC9YFbLvFfZXpIhzpppcBDhvyr0UV
sXdc4/+Ln4mQyw5EILSGBpUSwrW3fXXrQ9ujWBbezZaCCDIG10Gfv3aYj4/V2K8c
`protect END_PROTECTED
