`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A5TryJpFUKEFxroMia2jJf88qoaJLg1WVSpJ3EEROnrS+l/TcG/XbOeMdDNfUJF4
BbBcU3c0/nuXl8QsWt1rxhWhmq1MnMqqnvLWshDmtJv7QnRkGIgTVktUtXMqRxIW
7CObf6PLN3EXUbJgmHjh6epCq8W/zzGK1tyPFnOWB29Hnh0DRfirpTyXltEppV2T
51D4mwTFIkw6HbjH7tdMDQq7IRsUaH2erAMkWljoVSm77YawJTogtqON8kTYVIoo
Tj6ykUWje84kQYUhfv+PJe6J0BHvgZcq6Q+KdbmE1gcoEnyOlDnbHh5BNoFnLnRc
nKcrmH7HbtUyiMOs6/JkYnEJazCBgiHBpnK6NDsJkhQskH/y8n4iXy8yi31sanRb
p1ah1Bna9BnuRqmhgrAfpC316NoMePzOAR3HofkfPD7+MhkuJV1ySQMpAWka+uJr
9JHpvJydfaPMhwMovF67AMCbKGg9MZYGezH8R1uaCgYQkXfj8Jz/JW7KTR2xhsn3
dnQk2pifk8glddTPulILuJPdqzCgGgSloS1buOktkLJTkkYdsKOxZ1I5aZHg3/7r
7h+zbMhUIFPjW300Plbf4CC2YJgtw+RNAwNvwKR795yVt5AzHcKt+hC82M2cerpS
B7ZBlwqC6AWJ2+xLvU42siFqLPUB3cCYnE1dlvEtFppSjojU/do0ALLwY48yevkU
`protect END_PROTECTED
