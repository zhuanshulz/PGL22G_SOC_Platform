`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SnySOT59l5nGF96IAdhk1x2YkBs4ioqwvhFGhHR/f7a81TsqjVV/pas3BR9Ebhq2
a2/pT+j9ynVixR3488fwnXVdyZ1IG3eTWwz6c1hVVwFfEuM/prnrYym37cH/kOOp
oaxrrRzr3Aka7RX8vs6jDR62lBcZnUl3xdpGtO0X+YDV0nt+lN3hc89pul0QAPV0
zVHU8AmsPG+2ungOU1YUtupW7/pGLpf86fbGWNdpHCU5OoKnfyaL9zPzTSnKASvi
6ajaLtLeozU38T9433nEPLUUnto9Sf5QG8EcWK46XtRLl2yZvrk6CcwKHplYyxeU
j4/R1lmgKqitlHcI10Quoy7Akabr6eHwFKX/Q/sZZOIjy/ue7BiXt0QXzZTBdpiH
iBZOQW5uuCopvzVqJQxaowTZ8XbMwgm/x/FNJcYuFjUM4wlnr9kju9b69LsdqFBf
mk055VOVudtU+FbvOgSyip9KKr7LHG76vsCC1iuWq29Xrxnmc/IssBIFV6osCcli
LJ8X192kcxE7PgWHzFX+6keoufWHfZehi1aq/LozQtdKU8X1/GkOj4KjRSAx8cYh
l0WB5E16khupF8pWtRxkDq9t+0h3t9HYJXP5qgiAff+ks99rfILcz3jhDLJOZg0B
KzXVGMRTKNoZP+OYtjMzT8Z1Q7QVv20EIrI8avlZ05y232le662en6qZRjoMbr2S
BADvVa8f7E4hZZelOB8kCtOY5/shhnfEzcA97d2sDhqvEEpoCgpb1pnpeFy78dNn
Vjy/9sPta+zWYeEoBNI3M26p9sfMsSH98vMeKCBho2vM1ofUKN4gb5yS8qsDhqJk
gNWdnD9Z0Qn2URwRwTCTeaqFtjoG8hqTF2bomseirUHezXBLviXfDoAFjGVB6/Oc
yYD5YkYjM9AVsasGScOmZ97OvM5wINg3hlUS+TQP5k4hU8M6xIOCaUti7bOkYvni
kV0wNyPBX+2HAr4dE/C30n6MB5S8W4ug2NpcFSXCEErGsNY1yjPkd9nq1AVEnGwG
4q5KdKv6kWFlMzduVnfeqMLb0DdV/xRh9KKrhsncMgkuy8Qzw9ddTgGQkoCWlQQc
ykJ3V8zULbls0RCr696rrEZTG9UBN7aSDMGr86xTjDzsNg2iN6aGQf8udLXCqnJn
Gy9jtOSoxxY9Z/4Sp59nYSmnvHNJMLujauvfMo44kK+UDCKWStWqkMfKuHxwvt+w
MVADWrkv/8uJMTthcG8Sdl+oLosqILd4bRWicLy93oHXnz2PI9gnaby4aXhnU4oI
6aFzIsy3GP7uCWDoLfwANL3dP5iLmY9eRcYTz7LsObm9EKyZ0tAowpfqgQAVw9d6
s7rq6jxBi4Q5vjXRrkPyP881Alt09JSYP+/H7oNNThwvA4iMZF/lelsXfECVrwQL
FqmM2hETpQKrX9ynqIFt7Z5RjT0BkUcjxkv7Y4iCCzFksHmESVDL6jx6xPpIB7bV
lkHBsQmbCcLj5fAlfAp3aVURY9e+H/8ck24zRVbfpY4lDo3A3i3LEkdig4QBMhEm
gFXhkFZFNPfv7mb+nKOh6uJ09YAL+6udmmUcYZFFZyLrX1/yEoVrOPkIhwZniVsa
oUXmll+FFnQ4R1nLBLkgTME+FttCIxfPP295AjgufMSGvQm2fgjnZz0J+5z0427s
E8YATQc8UhuY5Kv0lC973WvRczTqQ35H5FujXRHeVqE3BjBBFi9uiR7a3HpGAcX6
49tjyjg0T7CaTqyefzqBDG40VVx9Sj8nb+lRR2feRP+fQiwR9O10H7BGx1b1qWpi
GLRoeQQkq5heQAiHk85/3RJNFsBBxu4QcsfuA2ao1mDKy3VM8YlO6GvzDEkQ0vmX
Amjm74JhjlHW/U6nfD0Ie4zX8q8mnsC1UmHxzTGiLK59cQAmd2NuPnt6aw/5D3tv
w7hGuP+aCJdm64roETF208AezB4GqD3I921gLxMxLG5dMlpC05vhDRKtWoyyevUr
Ybr1Mu6b6T5wnQUfCCKyB5ItkDLONxso0/jH1j7ZyIyXbFM5B+SW7fOnfkOWTecx
SzKER6TRtnPYbS8sG6NCF1jIidDmXVTnwkgRxinsFXB0VB7ttUdtMgi3JAWEJVZY
ZLYsaM1Q/vQXNo19Hsci/zfa+bZ9b0LS5ymRWMpujYLlcIFHzgL6nuVVDYTCOTnF
m/tehztJbRwKQtLb5OCacwHd1hHzuurIwgN5f6Zw+6JeJ4mOrRsBRnsvm2ROQEna
2qVbaH5ipH1B0hrfdFMK5HLwDi5jS01a3Wu2uhnAB+x7tKmbi6b6tDe4rVN+xmJ+
bZgqHRwjsnST5NsvX00S0N/KPdSsGAKV6W6yyZt3jSftc78gXVm/4Nd73JvOuMQ+
vcz8rnG8hB8ngiFnnTyLcJ9o8uPLKK7c0bMn80nTzxTCqAbgdX/SfhKJcYxKuFOR
2BUt/X2mocZtB6BhHWaTk0o2duUx/NKPnpHm8RfvBuk9c6b1O9qn0Sdr1i22z7c9
xIcsbxj1OB9T+TrbQIWVgUoXUKgkbXDq3b7AiZX/MQ7efobUngPSzodqSJARWJ+v
UYXjOobvbsRwW+aQjmh9JxbQK4vd1ZSMcsPe5g4M/o8woUahnydk3ImmtCLHzfzI
XwJS+St/YNZbR9IDnMiAbO+SWK+Te4Z6S2kI3ncKw1hXVbAplNTNSMwR9tidkGr6
cwJXLj8XNLUOQU2boyvc/dfj312ZWidBpbD3P2GI/AjNSQ6eKot17q11fOEnCjva
8hJOK8tKt1OhCnzn1rRjMivKAV6pxRDXg4pqddtpaJ7P2q+iz27W593upm2mzOfs
FcnCPcaYjHCmx5rz0Dctx090WLedY8Aq+8hVB1xgF9LpXv/cKP6u870Ytdn2aQTr
7yuY/WuzfxqE1bGg6U3AZ+BZgi14Pd+vgDhyklb5OIaHaK2F1PVrA0X3eGJgqaHo
KtXRlVEgavtWfH8dDsHTTfvsguv9QzJ4R/wwfozaiADrjZ7z62diFFJlS6AVKP8G
PWW8WW8aIK97qs8LTXyFua42sjb6q1mXqN4cif7pndIXkvIIZRG/cAWrRMabijMv
otzx7gceveaHvmk0dpLCOAV0k50NDuoHhId3KRjoz/MD6q4KSm+e7ANU9rMu1qFx
IQy+bc2NXNCOpv2urx4YIHfGwvLsk0RD7ieU7oJ5SrgoyVweZGa/yYR39rOEz3yK
zV4soy2ZYvnjJ/t5DCx1alBUerEw68rwrVr8tiabh0RhJUbRHiTtZy82nuvDd1Gb
ThLeP3lwX+PGJ3icxBVsKoxQQZjP3+rofpXBY0H9JlnvOhP22a8JWKv4mNnORq7S
`protect END_PROTECTED
