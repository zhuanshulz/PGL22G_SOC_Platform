`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+IAY2xs7iAVlcQ7Z80npCfaSfiYtcQww6L80eV3VeB+7l97g2LHrT7oHTsTDJiZ0
LD+p6cf9/wu0vk+dWodo3mQDsEUnOvznUczDN1IzDieiju8edK6sfKXCFJUiybgZ
8XOcUJaHFXwm6Wdx4vid7EPsCjiHWtImYd+nJhouGXAC4wpxA79tVT5ieIViBtZz
vyEfmma/ac3A0KMrSn/ASLc913B+eHvwz43FpBINMS5AuhJ9tbiFfihehz43g3Eo
wecgiGZuwHKFFyn0lM5hCoOZ9b1IeDfBqC5rqzz1dtSD4hELIqS+jZuaiLCBHKcN
NyW4qGnSQAAJ2FCh/M3/bqHeASBUXxnDIHhjQllLf5EXTO/4W9tkdyqxXsE2ai87
WT83nMWhKTz12DoVv2s6sFDyhUgNHAM3IOJmRnNKrQcDU5fvakjF/4CpHjP61WCz
/2tje42dWY1rCylnVADWXp2j5sUQef22HW7E6/B2TuV1rGfTh1/2syijt0lpfCc5
YCcSjDGwL1sZEyov5QfLNByGo+/+5zPx7Xq83WQhAgTWql1ihJBMISrstU4jogq8
ksViTVlruUC2w068sjhziCcnJyaIXO83z8L0eUI3FBMsttzis1I1BrEIk+DlW1rr
hWU8mlIz/3xwGI+lEqHtNFoTtUt56IuQgEB9qPHTt89cGpKtD8g5VrrWx2X5Zh+9
UH/+sIO4TKoJxBnsQr5kkxfDO6V+X0FMY3vGRpoFCsr6qLZHxN47pS962vgTakKq
ZqxKOyzzp4pAK125UGJISntFqr/+2lDc70LFFJEDHN/FndkrMDnW3DIX5ElSuyLg
lFZSPbHQKpxUUJLsKKRwDnKwLFD7nLrI5F4YL8Ckn+y6gFGYMfgyGB8dimVc+JBj
7VmYSRq5Fuqgq63FxuYGQAVi0Zatr1AbQrvzAqOi8YbLmZ2v7etHHAsNMsjj2Th+
3fix/GN/m3LNLuayIf8OwM5XI8sJPzQRXByRlEjAo8t17kjIC49MKxTq1EIwCFVY
TP7jDPQ95TnoyXzuxznwSPCt3qp8P1JdTYZ7J4yJce3LL5jlSRXY18kndk7tVXe/
p3TsCFyZ4u57aZscngCXCKW9kTgx5Q35mBTOo0UzrDS2gKn/mpDSag9YJKmWhQ6Y
yxb98IJJRKLKLWvWJvb5Z2UgHn3RjhMYhkCi/x2JGFjMgKjC1DTYnFWLIQr55QCP
dxh/5TC61U1YpJztg+Yn0S4t0uDm9Lu+8G3iPMy87Pqj7APKXm4gmmS1uv74gGUR
9SVK7qk8/B3+cU7AeB/TG13hPUiY1n2t3HcLJ8GHn5qD4gb6TAjljkqPGuxxfGOY
OLfLdH59Q/0J8mTXnMC3TvwbMMwXt9H9i8BP+j0xW7QDf93bOhbw38NCUmhUudrU
EaVqpzvjNLH6wGfhqd3Io6JEaz0Cn8jNuJ4CTLcj+rRQ946qVwFLGvbv3OapC2ZL
b2FyMuS6jcvpVjx0ZZmDcMBzhPACecTZK8nQ0EDfrOKQ7DJjy+vwo4hBxD2gdzEH
yWMkQwk09OnILR4snH0OA6Q5IiRymq23h1mPZoIEwGzHqzpTj1ST8EvKZJlMXRWT
T/lVV57LVRNkbmYbCCDFb69xUbBeB4Yze61qoU+ImQkZ0E0cDUNEBWPowrivCn5p
xprOhEk9dZk0KBhuG1R1+71oGoewIxUJlrcswY/ztLdvwKXQPT3KRk/TS8BhFKLv
D7+cxIYgfxfCEPLKEA0vFqCRwx6MoW5Qnu1TrWlAJlQTwuoUnAQDzTbVVOqBrV61
3XWMFPxi2fdt1lNWEX6uci1TQSExCc1KEjK1CnCiuQdNOtgOMRTtquxsUPey3fkm
BtnA/7Az+q3AAgXYAaLA8lS9orODTRuq9HUnDycvlK1/ZwZsbDC59rePF+sZiKCq
8FYkDCGgoMq2ZbH5+pkTjzF8uhoWppy4RgKRElzx5RosagWz14ucXdaaWRyB/prl
W56M5qapPrGxne0Pp6OIcNWZ9uIHEUyd8dmuir+ClOP9UQP3tnLrcX1mZoLx8GT0
b9uehZVqoyGGCVS+EUatdBtNsLpl91Yu5st04dk7STGoNDMWM//b+KQ1x3spua0n
aib4J76tsrmdCQSSS3rOF1QFuWUxKXdy1/WEbRvYPzQ8nXyuvyaolB6UhEl+5eK1
7AKZn7fmUtIITMoZOH387XLpnLZHif4TRITKAekkXaZyC2hPWA3Lf+JER0jLZQTh
EG0o+YDG+/Em46kNqaYdcRkSG/R2kkx4fuWJ7Sm7r+eyS2s17tF8iUWwcpKjuZ3Y
vedmbM0oYPaCRm2x33i+PyW51xJwjGCeBCaz4vchqPHHwV2rjybkfLlwkSo4NesG
Dv5rpXC006hsPwJeCVk7kZxnaDTZPd0o6syT+XK4TUNS5usA/PDrEJAcU31Hb05t
cLxOdVJ2GtgO9pVqyLmIDeaMi2i8nBd10umTjCSjshZ8tGwLk5b/12CskwRFdWmQ
YqyAwWWjSUStgtbcRnCHH9kE8aoPQvaCGcFvp0SGWGIeVB2oxYpdEq8DgX9cjSsd
Lh/OANDSPkX3QTnoAwGICvrDxHOOhJZmdX18Gq8XCmBm02XbLFPd+hPRKk+lq17K
FlTs8XviRgwcb9Le29cHBwMU4B1aN6MHpxBwKBzZIOpJJRUQcKQITTYAiCrSaJAN
ZTwNyOjJe4wqfatpQEX9OiIqYP1/tKSOpm22XxIisENqB9C755Wuf8UO3A3Gqe+H
920FMUhEuIGQQmGpRotBDeD03GfWbszudrr7IJ7eosuUfk80pbtyqwmIaTFk30+T
/UTEMrgCs3eXKZM1R8ltUmUgGxErPjtc/Jx1zyJFCv/SB4FrRsa1E9GZodTXYyJY
DS+OGSyrBBpiOCB+Gd18AAF3TF85BQ0aWc9F5JROXde794Cyy+AxvyxLtSxZoZjn
flQPqLwcDJ2AZfxGI05STq37pxnG+oyiCT4OR9zscAq/D2RJxd9xe2byRkmyuJFy
lPspvRxNS5E2Mem19Yq4/BTPcNlWh9xiOlRAXvOxl67KGHT+mJb7uUUmaXLut/7T
q96lQTl57hHpgiRvO+FpONU4ODb7r7DwYSvaP5Wzt+Hf7phxLb+4eb53iAiZy7by
YhdtHBGFC3iw/NcDHVcUadPLMrtjJE2DDM0CB8ijN8uwLmJwEenWhri+noCSrW9J
yHtbccIvwhSTEGh3ugc4L0c/ybNw+CKVPADbdzymlSVMAf7/Cc6uCrs3H2t4eXEO
d09cPsO4mLjvchk8JcSwAGGu3kIaSZVBAc5r6Mv1uEtwi079WRDXKylzpgFFfvBO
SDrutP78AN7HetMqOVi+tKDwNTgmFeY6JPSBPPnKitQt1BZqHBbJJOZuRTiqMK5w
mP+zQaBCUkLdA4rU85cXvuPzEuFMa/UTC+9jU47wUALygqcFNJvfoAyqQr9B9VZL
MDvBPP014SCW2LzEHfHIrLizXa59nvR4VTz1VxC6RSU7haKeBl3PkKy2GvFVoEn4
BiH23GucZrUgl/wRxzJ+JciJFnLFQxIwMGbb7Yq2YCyUGFAoZTid2/nCkkGZu+56
YNkvzy992EXthRvFTsIuHiRH4VK88mE13Ro2lln7UuZ0VMgM3VdASFZKA/WonHDc
U9zTY5UIn14Yf/rB//pNhtwdNVo8WHzQiHBMuLDIS7OCMGxtcMK3enrjtt/84Efs
1OGc9LVC11uPJbTmyN22Wia/fjgPUHDoXvcypezemxYefzB6hnmsabWw8ACR2qJP
UqIX+ljrUR3YMbhN9yN/dJfQjI6h5GJLRunx1pMjufDEKrUJ/wneq8lhkrpsrU0S
tE8i7VBBJx+n2sJhlFO/BycKz9jCxhYSP+KxcVNbmWtIwftkY+AaBVvzWMjJikQq
4IQg3kRVQDLrAE4uQ6hS7FWpEExpgKyWMOjpO9IHpEEHWzefv4JyP8MeNAhSC5rd
8R+KZboL4A3phg04RYuGni+Rm28PR3e/eYuQkcaIsrPXS+ugVJKpJv+9hY2M60LX
mWYcYH2lQDLjV7jR9/0NXQZXkLuJldDvgWnkv5ClKY6C46hGF+xLfTd6fTC+BW+1
s5Wyo2nHKWF4FbQXveTDHIzpC3s+bPnjMzx1+rhinGNoO7oB8lcqOzU4cq3onIgp
BsPuYI4aY1q3mjZRgCpfFK8gxaZN5gU7UwcZE43s/WOZ6UT3EIhl88LYSHTpogLm
lqZrpY+nG/y4lZR5NeOLRQK98s+hnZ7S/Uun5kmQBDYNlZcONFClNwhRb+mQOBvd
nyQMn1uy3aaVSJz1jB/mR2r9l+mBYFSiOkmh79LT+aZvcdN8QUVr5A3jpOp137kz
HZNqg/yc4kJu8ex1rEgo4Gf1VC6ReD9/cmKCax088fVikQ2N+PQlNQttA4gFBHCT
PpqSsbPjrG6Bcq4qUlr7JySVPjr6WYkD138orKIOP/501Zx+53mX1AuLgqIQ7WbF
ij0BMy7s6w+asQ6hHKdiHGNEoHoX2SaCi5C0Sc8dGixFpG+RbJ9LbrttcMApTIWX
y7WaGW9lC9CMU/3ApBRh6STa8my4xCiUJA3XL5FGefqeSor1rwY6iskA9niqd44U
14ZhKn7MUPe8E5FLP3xeZs/vXSGbhv4O8X2ft5UQIcCaQTxHaMj492gUDON+uXOd
uRqKCDtZ+H1d1hQZZSOwqwycdC+YJuIxtqJElD/MnEvu+sl3unfXqF7BNEsmrKDs
9UL0TznDRVeZeOFUBEiCY2AWgHw9ED2GWeggiu9pC+Mgh8V1QzlKQUCfax/sxg3Q
oOegYml0M6NNck4hxjB++s7BV/vii71Gc+79JMjylxsbT6mkN1iGAr/d1XS2mlSV
9gJZuKay2R9npkrceKznyEGcx4HsqYZ7Ye8tyRNliWuOS/4gc5aOa8wWm+bbBOro
dJUQ6g9DIst2VPCONskbcVhND4Hcd5gvpQ9m+IoaKwxwgXuDIDs2Z8Q91NM19WX0
HkAXXz5SwVy5o6unD/pW5yM+6LfWl/jmHxhzSfPfhnRDidrGFvXUEZ9gDc0bgI4s
ynzJjHeu/GR4kp+Rmo7CQHJa2477lrT1fo8Jk+XFezcq92wow4/dBgvIwUI4OcFi
KCJQzGxcG7g0sNV40+u1muP1LD3DIGS59JCM2GC/h5JXA9s9/Ec9NYH1eyexuxiE
W4XrVH6YCIgk+6OiNnJS5XiwT5kex55eU/0xt1py1B5N9R+6WkSCC+DTRVK02CCP
jJtW6cbGg25KqYN2ta56k1rhwOpE8csQygmyQBZpoqHly/mpiWeV0Oz64H7jtaAo
KWKDg24VPmBUIuJhAhpbstfFBAT6Hz9MDtrrSk8rMrXQ/yjtcVHmrJlIkAP/EBar
ajk/VsMfvgqOnzJ1glEmBmTpuQeDYxeTyMfDSZMgzde3JSNjB5WQ5M2FtG5alOCh
G8AxG4tkPOubrV/YbDHRTJOpSKzJX0maKY4D8VgwYR1/toS3RPHHiuo+DUlGvWmO
2JepBkOC+WZ7qHnBnG2QmUZ9qfaimNx28otqSz1YjN2tbyBTiBaLVA/MtNt52wjA
AtNGPbp8/3Rf4hxZr1O08fRcfMFZvprPWUu0frf8IHqd975sNnZ23VGiByYr+1Zy
uTfg+MKnJgLC/U4sJw6VOhOAr2dwZmZDnxRw1xdeqcJENTCDsbZSZQA3LpXWz68Q
7VkTWcV3mcb0ReEVK+tHfFDz2/N61umu/9X6cmyyUQ/PAv6k6iQHC7D4/pv61CBZ
bAAKo9TRNyA3uoXbMY04ceNXL1lQzVo7s4nHbe36gwmWPkcJPTOwXixJI0iUXaHt
R6kEaDG9FbNvxEgD8D/vPMIanHbq4Ia3CsnWt6skbHU55Ud/E9KQiUxuNqtGxsEg
JvLk+329tVD8TE+N4VO4B7trpOjKZaoLdYeThw7NpaSBqNNag5Ox2aA9TgGt/cKZ
FsE0Ih5l7KASGtKpAhTr7j9FWaQ2VM76nz3qbRLPrYD5QV0v7s4agEZEdBYAKPUq
YGPGHIYvJeb4BozFgYqTzq5XlRwk0IghgDoMRgoedbig6bcLPmKlCykpcQKbgvVV
7sGLNxor8JJQ3315Wil+hH7zsY47SYmqyf0jIDokg8LC3u3J4ab/7ak9cY1Fm+b/
0M6FVIzlD0Xa2ThLBSquvukK9BKM7pBN+cRrD2cavhP0+AkEDnjp9NCpmXuJsRhi
1Cego+N1KgZmDk8cfDuU8k8828MjIpAWh3ZadEZ8QHSVW3vxs7XKd9XnmzO5+198
DlD7B2UrMMWoct+vU/xRKsGx7KWKf5TZE9mgOcGY3gwcBiRsZMPqSPUGsXpMoQ8l
DvqVN3iy+HVNzA39HazoMR6l8Vh7muMc1bGGldxfPVnlV4xYBpHCKiojmheoT9dM
zdgdRfFMCRGlmT/9dwLoRsiSxSN4b3zlmyWfiVLDDjxWl/hNvpHbG3VBOu/z76+B
jaKRooQAyMQ1pHzjQL+UO8LAvR+m9OKYs7fXXdE9OZsIbV/pN3lHSK3Dy/PfJcjq
VSKwQr9VnLFbZcop6w41mgopRIxgRILEUKQbLP4UixnJpuYiuuniicKTF7d0qZP/
LR/No5HcbaH3VF6ssIui3EB2dSuTEhnEXB56SIDAur5Burbqf/7x67n7jsX5roWy
VQlxcE75PLcQDtrvIBybQB/cdCmK399UjehaVuOBu5xSCFYXM3ylbfdGwi5yO4OQ
+Bl7Eo4buiLncsQ4SNuSKRudvmFRfdZoTkWWx1VKfXnVdB/jHNCl329XBq4UkOsn
5UIXGPIK3QB6UF4nuzhr6pM1zhfzQiKsJC4PmDytX5i+QCaU/pZgAzqoN1ZPlsk1
HNL4r6YuA664ISvF+0lFmLhpsDmDBX0W6NN0P2rpW9O+PGqRj6QSP/kkbeKwFnRe
+JIOpH4lCXGANMDq06zmJXCE/MiPZrI98TvJknzH1Y1si44JMWN7Er8ygsHu92Yc
aJQkcgDw/5bfGIWrs9xG5n/TCUs1degiggJQRTfrEusH55Qh7Nr+4vygdqRlZ+rG
GFw6+Pdj/Na4dGWVOItx3T4rgAp/r4c127MWu9bz2Br3i1Er6od6VJuOySPMVR+F
q4xEMUa2NtHDl0PnLSWrpYb+9dHixG892yrnEjqDGdT3LgEQfT4i3a3dqwMwgV2y
oRx9dMIkxCjc6Wi7AGlmy7MiUc13xmQt2rsq4CLnnrWiD5+vcj4UATAzrrqNe/JF
Ro50geWpeS8EkLs+MJoGUKXcu1QR8wSQQoxgUvyaIfvdVPlqLKPefPzapvIfY/Rl
FqRuh3hRbFz/Syt8W/jYgeprsCcBbRanGbTw+mvY99ET9LcYsYGHm/qhIcbIvF1Q
IBe4UQCLnglIG60R95Rizek59PBLl9rRRcT2EqPHNkazS/FCbllZGL8LqiCC/ZEo
rHv7wN3XP5JAbQS/2fcp1tGMlb3TMrY0Xrfzs8OnWOnSze2vIAg4sySToVZwAzNu
Jr/dmgVQ4F5Q62p5aNnJ2W59WmrgNJkvcL5Z/6sdliQFnDy7xSjVHvHbcgif/wKE
DGtliH2irQc/lxFPtEdUnCxJW1f6dka8XRNHNQtkip77O3r5gX53ojiLvTUMjYRb
CnybYOxLnuA3uA+a3hyHHmdeNSCesTvqf9I9+xKgT5WugR3QfsEVL4M1ar/H+uBj
/cdiGAe1pBq+qOCcY0cHybn7obFVgwufeCJZhBto2Thb7nuWGtIOuH9pe5dWnqPr
G1PlWuWTqUMpJicb52tMdjvcqGZmlHcd0bbAfNU4W30Vk3VrndWmXrZvfYMWURNG
pkFFyb4ChfSk93AGykImtLWWbkLFzpxdBTmwSX3GI6m86y4h3qZNiHTl0jrLbhw+
NJ4Dx7AmaT4Lcv9ClDaR1rvmZ/t1Qkr8FUdRGPwSChYpzPsEnaUVMP/7KC89OMXL
iizjpXYOmdIh+XyY6vEC2uEVR/oe8XikY4yGjGrKd886Pei+BrJyOOi1aFe2yW1m
2Cx7oP7t1pL6z8AwXhBlaUj2ETqJ/RxpxzkD2yYObhxPjc6rr3AI2vhZxG0w1hdn
WJ4YgVkJQDO94o2EtoiFnp6IC0acoUnIrW64qbXpWhm7OtE6eT8hUpaVeeyGbEiX
Uksc9r/TVQ6fQ9fOpFWImEhiv6D3+/yPp2K/4ZCH3mI=
`protect END_PROTECTED
