`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N9Vsrk4JKjMc7UcFs0YAGLdckFIgakuusAwAIQm5VC9PuEBjDmYrH9nFciftlmVy
GJeSjpiDr/vMY+i8VSj6WRehUXmc+w33IEXdGtgzlowhi77dEB+mWl9izhzhG+Jc
I0HyLu5r6WOS9Pk83Eu7moYjJmPiidpMSIWBsdkVm3I0Pv2WnlDljxGUgHZQoRao
ysO6W4UNvi7UsVY67WHJUm7KOxI57xefK6YiAhZZdC/7HDP+ckuIU1Pc7I/1PrH2
28mdLXi68AbuUt2RF98pqGaN4jKem7glaICePv6duPjIBB1EhRFef3qB2GbmvXZi
CuIlCqst3XQW6CyYk0knXJNE9qGTo2ypJrp9jUstruge2FFnbR/lkxN0VB9JZD9P
EaiSrgOp5SssfZ1Mva2ssu6oCR5XxQJSpDykWmP6PHahqShjOSVLYzjIy2tcyBDS
Rj3COJQIAHBHXPrKkMzZFXFBd7GaKx7sUCCl2rwMH2Tka0HgPvSlc6+Z5UhEnQnl
J9xb2goiI23ukfWBUDnj7VfUU64U9OVo6WYNWOoezQhPD5ZW2Tshf6rndcBqaYbE
gDVqTSDb/yvTW5nUSA8mGua3952AkeiabPlyHiXpK+rtB5r0re8C2uDeVUYjl2qz
nHIbSM7fhsn08ZeCoYP93zxlf5wJUt3ormzsUEbRfn+SGbEHRp13txp0ixlBlyRc
8RgJuagQLvvCrPta31qGcIVUVSlLPiDau6Xslp1i/Ah0xPu6ssdfO8NRIRo5F90S
0ELecgkN2W/1x9glL9lFZj0MKpVbeU34YOavUzjYuTFwwBzxX7xChCh0LBZ1T3/K
xO3qDslKxhIUui1AK2DyP7oLDaYVTzAI0FOvMHJQOPT1sKFL80jJXAIZHblKN01o
1Gz5eKaLkz47Udlbibk/gqOB4K5KmhXm+F4LD9OvfWM=
`protect END_PROTECTED
