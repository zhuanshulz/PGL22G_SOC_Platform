`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ovUMHiYqdpS4Y8NvQ9Z9TIO7WrVI+EPZLJynjv7oU/3sscMu+ovr00nr3Zg5zryr
SRmPxHRjjfGy2Wbxgo2NMJz6a3BagdqYMVPMT42S8iJG9zHuHgYkoaRwcxsJYqhJ
dlGEKTNipo7NVQr+rUZxepBs/ihdKLELS3vAB23hfuXfjuHbjjXGerDwd5mDu9R/
gD+g1/JahU+N3QR1PQ+QrA9fp5JVkNcAHY5qzx9/3BH7ko987rKfDvSx9/nZ2DfW
BY0s+NpeW3ZlsKt3k9Rj0YDw2Th80PG4zkNGhxmOmD48v3pbK7irmcKZiy/WAk1e
u1yIVogR3iSaR40oglh4NVnH8LCJ/FAatFwvQN9PBeP+Tbhbz4Z/CVig1n0WGlvP
kJnWOWDq66XC/8HJATiIOJpZwwtl2y2lOc96C+EYq2UXmbUjIJxtCsLg7z9N5Uvd
8XztGcpxfkQvfPM/+dYQ9V28qFm8bbHVLEwpogBVkoBHdp7G0ksVPjF6v7FHXnjg
aFFSkxhEPntZLeBCg08qsLjwtRAJ7+U/q+euPu/vlmNIEKk7S7e2DY/bvgr4W85/
F/6wvtyA6eZZreJRfdQ4rrTnGXWP0f5UjkCefoJjANwES1YydfcobWuFYqBCLId0
6+6Q6GeDn6wA8pYiL7Y1ZdjXkKesshiZ9yFW8VfAJ3MfaC+ET52dJSWPYPsS1gpv
AfzMWfk6+A4IqCdN3CkYmexg0L7txfpNh4XfoBHRblYKIybl5UgiW7INBckqyZYf
Rd7obDtf23nSMXgfOyqGyJFyylCWDoRDOF+j4UR59tyC+6zaYDYYSEnte3DE+RBg
Jm6SVEI5Iboyw/iJFXom8soD4blCdVak8sS/xTyv7FDjxxmuY1REPLT1jSeQ5mYi
LkHD+0rdLWfDiCMYWqcKhlNL8Qcq/jJSVDZ6Nts8UsAZH6j86VNirrLJXyURq0rY
gbmY5rZcB5xCGvj+00wBMzb/glEUR/O5N1BzmZg5yZauiUNFMSeG2pNzZdwlUSgJ
vCt+5uD/1rwkWLVskI1h3FtFVlIDW1il5cs0tZpmWEnfMgSZzLkD8RSf0F2WVrEh
AVLy1LesAptJvCI7oGxwAjE92W2M4QOT3oQiOFi4tZw+lXUlUzzEkYRallaMPlLl
uljNaVukEC9ygvzLxNanuA1OXsFEaswm+SLuA2eE9y0JCvH8C6hJ7FVfDvj8IpmP
n9KSBq7PBoH6Yy9u8W5PW3Tl95JutsGffyXuwtw1LKncj0m0v/CrfiZUYOfnZC+3
v1TrsQZnzqsF2Wqh+PDY66kjXe9c6sFhmrKOLn763qyjqR95BdIZ3LdORMNVZ2lv
DpfEirlQhoLnYWUpLUPgz6zZQwO1yutr/xSV9/UD7vSP6ZFtkYNUu8d4K/d/J1Y7
xrbpQfROEWyhPq5tLCTfHxXb67JR7alFxDgOV0+AFZPql0oizAfO5afDIAiOzzbm
eFKllIvWt03kj4/7JQd6/oStO2zVtrcVgHe8DDTkyM1QGO8j8iMLOyHti0VxpYMI
xpvOdOmviupsnWcNzdqZdqm7EPgt1TwW9GzgB2GYmMxvms/oR8eB8DsqtocieRNJ
RhELCx0+c2qeUdEZsAiTnAgJLBKEbfAK/DQGqJiYSqJTGpMFjn70OWugilt5vH7h
tw2e+1SBsKT/7TmqHL4P+pdV1TxggNDSW1NFG2+hylkzIKQ1PHgfwS7EA2YfayOc
ohR3KnShRS1lMvFCMZFdmS9zUeOiAyIKEJ4lrcMbdN+BAbVoOu+0II8qTBa9xNhH
zBbxRqX7oFcrVlkl6mbb9RCCQahF+2dkwfUEiSrts8c6bY6PjcV46MB3VU1dc6wM
t4J58TyBz4cji8EYIZyuM8GWZDDYcJ/R6W4XwFM4NrsgW6I3315hA3jdKwEPiGsv
gEiae7IuxU8caEA1gqnWYhHx9YhdigTRQ8s1/j726p9GnGGQ4Kmg/khe1+IUbJ6/
BJviAI0T2/Zm4PWNkGiZ3zmOCwSi1GSzdlyyBIldt0Q0t/vt2ppHCLEXoBmQNqAB
eCCfHeAqo2codebwgkNeDpO0fCGNbng9RAHNqwfojTJbBtlSrk4EU6Do0oBhqtwS
i1SprhAo8pmfboF9cbyKug+Jre8IkLYf6F1m3RLo67jrC4pvQRZC3xn9nzX8Yy54
JUet0zhCHPA1K5wffooh/1tX2hVf+RYzru4ODwpFhM/Ll8cbeKSZ0lAamXMFyENR
GXjqAnY/qForWL3ExfGa2zs5z0E/OTaSo3HEpObeyEhDix9jpva6/0CEv5RO7FYD
T3Dl0I6J8ciUf8MM8FQfNurAGZCy2qjJH9l6fzZOOCTvt6uPX2OtBM7/8SVykIme
zcIyhfJMYP+U5ZT+/kPTsdfUOVCA5R6zuTk9Vztmzggjp4z3qd2NQeiiD9uh8eOJ
CX9wHePNA/eFP6ZRqRXbHTDGV13akLJq8FM4PD8pvPT/GHqR9HMmfswo+fdPD9+S
`protect END_PROTECTED
