`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9yc0DNalyed4xAFzVXQKVctR7E/H1bGpCwbr30xg7e15Qqp9ksfuFWK3w5RV7zwj
yDT324q4WmH1t/H/rHmKb2Mdojemi0wzEHmwO2NGmeb8sSlk5oFCf1ZfP+JdlwH4
hCO5STRdyMkhI3GnFtTtNcHO6BYRUBvg/9ShQ2WIfO6VkRAyx7y+xTvRd46mBkT4
2fqyT6cMjQMNeIHK2EHcjlqCMWs8Gr12Q8Fv1o6Ivp7DprlUK0h+/gDG2uToYkiE
PFlbF1tL0AoCb2ZHrlUJrNMkt/STQaGA1akDPIcYlfZClUJOdGyq+rLrF+Swx4q7
qCK0hMNrqm5Wm/f5ejO2/+Xf3CbZ+6E6K8hnPW7SLP0kpM3dF+/yIsKLmtqYjGWy
X0NOTa/yyfkDRtHprrIGD+rNiPX/HXVJyXWBs2ugZbKU8R+0DUpPRkXUWtaN/tYZ
wn13wWgVUnbC5wiOqzvKePSTASn4yOdJUU3ifzmtFEVVlfL3OlM3FLoXQJ0QGUUT
IbXe536x84sei7gDdliaVKW0Xn4Xa3mW3e9QdmFteAWPwOCgLSqR3djr23u+kIHo
hvssKXwI6yHi2K7LYBnfQEd2YM9BgwlZiHQ7uRCSdCPiPiRPyH8eMcOM88GBXqZK
glgdTwUgyIfs7sVAegs1vpOxJeML6zUxpk5d5mL2DN4bwjzR9fOGa2H2bQPKT8Gr
Xc4ZVHQWO6wuk99SRvA9tYtx3gmirXuIOM6BRLQvaEgZSnTm+8ri/AIZFgtO5iHE
A1kTpykJbsCnjKQ42WbJQWPYxW7qOw5m95+BShaoZz3bDDtJtulfYs3OwmrPtkEU
GYqJuxmREbnncfIknMkoWnArKFsDiE2hpRk0WE5nJmwOmNaf0kp0z6oGttQaqKLz
ohkD2SEL9GcsTQ8bUYy2OfhwlMV4zz0G4r+41lIo/yIar7FZhHE8UbO23yIE+1+W
7fCxmI8gEXEyH6DEPi//EJlozXI+BWYdMEmRKXKcRwshCu+nzUB52d0y6Ae60B/N
GwR3ms64i3PHr5zHNNMocWoaOn8mTVhF/fdoiJQI4PnlEpnQYfQ85EYhgPgtHdSm
yMjJ02RcZUm+mSknABahrixQfofjsfu/JoEE0JKVS+Sm5mJCpuds/Zx0R8JP8/rM
/F1HqsIX3ph2JCHsGS279ytDZYCIjkquschFv1dEqOppPGi8pTZOKIYiUPWXAC0x
FH5K1mxg30TWcJLqc/XxtXceXhxCkSVG6pRcBWFDM4ygEOkpMJ0TgRjE3C2kN1aq
1MU6u9l5J/H+CT+7M38sntjmRCFZMJlAIckwQaknBwFEoakdj7chfazzIA8kHYV1
Ny0AB8vKiS1qod/9M/zcrWkFZgdq+IU8fdgXvhwILXCTsEfAF8bzeowDyBS6pBdd
teVuj2HzRWu2j7pKq1/ePsnZvFcAe/GanJ8KeJslpUlcKG3Vz7QeJbuP/KPs+MR5
XmNS6p7I76rTAbk5jtwCxmBOttGfro2JT2RZcshVC1IPT9y3hYO5O/yVD3Z6P4zl
DpLxpOtCsKznEENNxR8OtWmA8v4kbEZ+sule9unoNaRk2N72jtfW5uuAQJeYFljA
FIl1TGQnV6sDY9wHr+vdO3Jm5HH9yv/h+/hVXg/nwKaO2WSDH6CkmDg1DPM3s7za
QZhm3rqSzgefCHZBqZ4uG0kz+RpA+xn5MX+mCiP7mnF2j0VjCEPbaZsPB3Gn+l2w
zAVrcAhrx7z2LV8FyQAPVyxW7eqc5YdUNnSkvicHhlTFoFix3NFyxermgtv3MDh8
BkiAvABW2MnJ2UOp/DD7dCUw4qOJnjZ+liL53G2JkZotzlJjJnqwi2zKQdW4eHf5
DVE9IZlj983A396M9d6eZfQFmH+xtfXhi1rl1PAoUV4MPb+QHw901wxXsc4LyH05
huPTpno3Zvca57cHY47Y8+b/nlE4ZVNTd2Gz6p7g+ubI6lBfylZzofSnolrX7F5x
+Cshiz+hzCSEeBE3xTBz1Aic24HfDPQ7yBXily/qYiMmcSja29liLOf3ojt2S7vp
vBaRkNticKu/jD5DCYQta+2hrsyTu40SLtuxSIrYZnpEhDj5RVE+Zr95jg5dbPUl
4UxnSv11vtozepka9o10+jI7k+4tRJWiNyDCrEDhkHtYaZVopvcrYEE6DXxx6tUg
VRUUitDZRfWbkwTRTHOcBVRufJqPZiQ22MhitoqqM2mBwJ0+3c+gSgquDrQFAAsT
WepVQSJfHGLHEuGj+k/+0l5/GgNb9Olyb6v4DlWWK9ovj2+dZGHp9CrTsYDIlKaP
ls85F3V9inA0IdcLglHD1552fkZcogwnCxNjl1ZddRNOCGM8qux0o2XZ6IHHMh/7
rxZMbFcTwxJuBybSGVQZgQW7pVyxSO06p+bwW6S8JjMNE7vjFyk1uz4WA4OGwDm/
Pa5b8fvtujaY1gUT1mAOh00keoBU9ysDnxoGtXPpnp4Pqp/1h19RjO/KYztE5zW5
lp6zClm671CbHYU0lv4s70WtyYrWAHQaEss2QvHInot2ocZQCXxnsvgVrjyEyB9u
IW+KqsiEByFmSSPOvoalH0W+RB8akSJk/MHpzPMSP8GDsuEctNAe/ElWgBtKvuaO
smoBATxIcwM3PzKPGBeMwvQwbcaw09SkZqpIiQVswvJDIXskAumkFPG8ZXZ5/x/c
Q5ChHUimUV5b/JX07fx6CtbtRuopW6rmuB5DZPFWqCvtR//X8D/U54lS03nFpfnf
Jn49Om9MjQrNxrgYUkqpupORp81B/0Uv8FU/pFcEigkWqUGBuzbjdPoFeQ+VfAtA
yBiOA9fabnLqvGgLCoQR3K5GsoIoshuTfFSdyeEhCQSaa8UN2Ikjx2dRNXadrCB2
LRIJSqxgDsE+WGtZZuCdXC512+QHex2vbgNfaUoC3XBqnNuG5I1/s3S2I2vuU402
y1AkQobx1HXCqUouI7YlDfiZtbAyJLctzbp20f/zcDKBFm0BjG96LkK5Qw2qV+Zs
7x+sicQ8LjttcT+yylfJ39f+vKrKHYlsTEio+e1FffeO+yfXJsX5OAERC8h4QdKf
5akdV33MKRVh3NDHUBsITxUEvg0t0G3yU7Dq60sp94qvzEH4f8w8oOFMsdU83ZRN
HlQw6xDmu24Hv1/bGqWxRFdWSyEPoyzejg83EYugqJNa8hPjDQhhphvohmTrZqla
kYNwlcIsAVwNsc0rRGBNBPSz9B81zlAU+YSeF+yn8J82B/Abs82HXK6moD8vCIPD
JBxivxRYxYw9PfM055IuWr1tPsxO87AfbZxvJg3hcbkQ3PDnEIwwUfdRA3QWjMte
e9kckM1v/mHHc4lx+6hQEJXINAMJqdYONhFUyOFYPoUjSIoRnhF9XxTAi8ZdpZCF
fsS+X+VsS52Grhy3L83+PDnMIkaWkRRbL+cMSWEEBB3JW+KYdAdbGS/ON36Fp18+
RY4MjaOWAFcX2ZI1OvCkDc73QtOUp1XqcXBPqQngYVzVb7oAoqNWi+2a8h4Bm6XL
MgIe36s7ZcdN+1saDT33GXkfjMKrjSZzejAaiHB4Fp1W4VHqur9QAMOxOTrCn1e0
xQ5qFhYw3IB2wzoyBX+rInOwRZUBlu8KpqHH3P5FDWmyiByYK3pxf1U1ZFK9KJMK
KuYJlPCeQpv6KbMghgNPtT+6YZptwxAFogrKn5UYwxx52t3ptXhob5Jh1OTG1+yo
//We4ovccQwm2yZDYdIyQgYQYBhgPzrCcvKZxOIun2CyLYrR8AmSfO7SQwD+p79D
cT/NIMu+lpp8fhWUZQNoyDDr3y3Gxmh+dY6QPyCPWKSqs8Gl73xkxoDDkWWtTNl1
uSbA703muFo89KF8biaZabPIYVzOX9ZwwEfJXkqUcnqsBhTXY7444yrYw76bYlq7
sWKnJWSifMHzTEkgElwWcMtbEY9hM3GH6kD4pTNbmFwCGgwapYoPILBCac7ss1Qs
XuXDoofy3sXzA8AKvglWnD08NByxmdVufcq/d+jzUYi+Mj2LKKfy1rOytd0ynrjT
7Ag8BmqYL5/f6T8ESVcrpNRNj25NlnnMDVCPpC5MGgC97ueGiC5M4AhiFQjuIQW2
bO2YaqMqDk88zXtjC9Oy6Ln3D3//FLfqdolDz6ntg33PFkMaloPZ6hTYVVA6tlKV
1wVexM6dEG58zHzQ73SwQJQUpaMA9JFOz+/lmFJmfbYGFbNHBz7hBN0cgokW3T6C
sdiieWY7iG2Zw0ghjSVA987uoa+0bzZGfRfp+OwWOmnBgfRAlWbfiSXPThz0duL9
LyRO7JscD2htXPKYoDqu6i/aKvYzEO5futEDDl5ZaKKG9Hne+qcpch1kuWfVVtz8
VSQGYeYIZsXlGs86RFQzMTylDh1Lekebvs644PR/IrCUoz/gld/GDTQSf2AijK3W
LfaFKnv/C1pRCr2hcxJPBy/ovJxckUOMWRX4T9rsl6bzWILw3pAkYNQhAwl9ozMR
HCLPbcPVQOV+EbXPkNe15FTiieqMIp4tqsRo0skKbYZJGrQMYAknURTfrHJs+akk
3jVPVGMf+2ndGBw7QJQBWE7mnjbOo1PKzUqz30AJPFEU5/fxUyW8ZOWB6SHcwJke
8sNV4Wl+8qUznKVWHm3pWf12j0wqAD9rwDXzKlmICuqf8PsyzGPYWZVItxBYaxht
5vKj1PmtIfAHqLjGyid5nSEqrkMZQzIpHr8ZV0zeewwpF12usTGk+HKVvdvJRniU
npvQjWU6eZwob1AME4QGOq3lOLwAfZRmP7ndyqJhBI68OyzXAKQwyIAovcILgpjt
+qyAUC1WMWTMQOgDMJ6m37poY+E3FIU2TzmUQEHxml+bmaIppIBIjQKWbtB+rFId
XL97NY3W2VbulsGiKnlkMVR68CrKV1u3MZ60+UhI12ATr9rd0yxNtqCcLgZ6S7KC
iXFbwtOT4R4yo/RxZDyWvyYegugd4LRVBkN8jyMUBxKBCgI8DZwrfvpKfCs1H4bF
SB1kLriBsl+6BejY+67lneJum8DS/5L59zrJOABJM1cI2TFBpqx6hIoeV7yqvgdO
YZHyjKZzQ4v0Jlnm8hqAh54MRv4M9eBraqReBWRuzQuNlz5S6moDKWVzE4KHhjZ6
ipr0TmSkpGHsGdizVA1OtJmOlL8XhG1NQ88Iyc5qWEdAcwofhsiWOvSjqBfyi1Vk
iE0PY3JS23Vn9DR2337zd9qVdBxL0O90IH1dVim9rLDewZLXrEeFlst0MbK47TgN
YVimli+zuvE0GN1ypgxkfq5d0+KQMWlISub3RsgvPivVoJGc6jy9QVWWdCMc6tnR
0A7ck+8ZLR7BHtpTbzurWAzaHid5527KpO2zKvKVQVZJouVyZ+8iDyiiggyNtt5j
gZ6MoN4USFge8K+orIVVPwWTry9ey1Dn/4R6gqWVkevnZ5kF4MK+AmpmRD3OkjCp
v9K07DrWfggg8HLPb3zvAmfJjuUIm2HuL7k6HmWZRl9P8dNV6SFzjmxvikghp7oz
B4lMIUgm982XvLZ34QG6YdilAnHyXx8tU0MMYBzbqWXFHv2+c/COQeoVBaXpO9HW
mI71zVq9DMxV+lyJjvW/eM/y+wUINN2qbaAc4Xv9/dgZba1oaMBNaIWwXMouJBtF
qZ38F1f6tPAZ+YTdwxYAfj0rXuMtllhCmxislZWQDOeFym48zN+iT3e871ccJHEE
4rJBWJVnm7cdhkYQkXb2yEFLCX0DIRVTihYmXurhiESiGF05vuq7287NVToYDhZe
0j3xv3rLC3cmwk2pIjpQfzx2RRr264yiLU6wB93j6BcXUlp0WYI9zG520Cx6tv6h
iOFSDAljg8C9Zkg2r3uVMcsEBarNsSN1igdTxXv7yHrbAiW2jsal5xVnGPPBV5hA
jc+JXGU9qn6DJ4TH5eQ+LE1pOUev9utCloEPfP1ogZoaNaHjDpmmxSOENxQDa+oi
qAaTqKCknhBurAwi739ueqfhVZIlGfuPKqZAqrEgifUubdveeJySYIOXflXuyw5b
iRFFzXnENMTj6GzOpsPD+Ov0KMmL3ct3NS5MiSzHaxoqnlW8TVn3u/C6jZHPh+pP
IHVFy7dVukxQiiWFREEYj3QZ/axyKEglW12xOjX268HAKM0Mj1PHWkA5Cqkr4XRu
wPoMZmCRKEtEz6QB6qYm8sQaK2spNGbOsx2jbZRIx28U++GTiPsxmTQP7wGtCQqd
/t3i6tf0Ud9ZMb5hCSsK6FJ7L/enNXJO9hs3bF/ecwO7bOjsotMjaQVDfWlwBu89
ePJJTGlmoao15Zc033QWVgkwxqsZWqZzVd8T5gchw8B4Lk1aoLOOzER3cDTzrb5/
nLfo/bzTwHjrQ23+T6IlARZlvjsDu33XijC41Rj0zuo00Uf0G2wp8p1/Vd4zKWJi
ob2n5mlmN51NIWdru8vails6BVbduOUTQ2fb08v5jOzvS+ixtfl5cxHuEaz53z1u
MTqFRgTpSzqo9/g7cUBVRUSrvV4yUDWWmKUgXaRelteR55Jk9/zNdTJDORzQPSTJ
lhZS6GDDLpGDw2LGSViX2pXNSIpe7MfVK+2m6rVjjFMLIRq5xENlAfaASCGHEEGd
eLDPCMfP51dKt4O+dz3lqoC5LEHGAEHl1qiFu0xoVVPHRNWuONIpw73bJT379Qq6
amL7fTbgZf+1IZH6FNqwz3YoWY8k86fSV3fuB1Lbk6z7eRIqwgMvlrTtuMa+AvvV
+I1hhAvOaskkYPdXJTCCXM6WHNm9IZIlXAyq8BD6nrAI9k34t1i1piZXqz2W7Bh0
HbGlkl15EvZBh3peBJwuYN+jlOcpYlWEQax3YWcE6DQlgY14sKAwToXCPY4MLaHY
EHrrxfYd/Fq2nzTK8ix+3U1IuWwEG7Pe90tMomFqupwPem2jhvv9/IKrW2Dk8tlg
jESQwJIFEMidwbMwBaTbRulZv0iYGQpVtkAiRhGTUQjeA9AwW8S2vLBO78tSSNNt
Hox4FLsZam0QFSyHohomvyTc/R/oQfJXtzaaAy/l31URNH/m4uX4LpzYvC/6H7LG
rTTU1PvBiItP2FkTPL2WqWqm5/yggI3yE2dWKg9eak8zyt29jFbdrZ+WzWvSDWCt
6Byk2jw8+oyYdym8J6T8XMuqWsv6EVl9YWICEM+zueYzo6yhbjXj81MZCepYzK9J
Xlq3fy0mpZ1HIxyFCsiO8M3zm/HtREUiyq3xXJHU0N35dJpsTx645x3D9QO/G1aJ
Red+btDz5p8BbhQPezkWZkKTsXJqCwu7iXHgEycKareHUz+UAe3ugncLar09+ZqZ
h/f/Gvb1YWSzKFcifTwVIfihG3nrqhhWtC6TxzGJDt29sUtlyVEWsU3bgQppAVFe
BrbOgrSbhBfm8NeZzI/RMwghbCg91yX93axwpEVnJH47FMWdd68BbGOLAyEECRKo
dXYR9ptwLRZoz7UQLVWo+bA6bC91ETuJJojlgLcOLNUz9KFY2/Rh08EV+PsL4qrA
I0nD9yz1QupsqMhp8PIoDq49GYp7P10JZ8prYkLISIMVafPBtkT617gyrpTAQzep
e/8t9C5+vT+5M7ha54NcIi6xzJTcsHNtEuniLDDFLq3t8ve6lmiUCVkfp4MtYZqm
WE/Pu5QWiXyqfFvP8Dt/oqtcA2ly2jkZyqMDHH6P7+JzHSbEw6loSANjM/AARrml
G3zrfYaS0LTYO7I7MVowYx3G0p0cLWarD/PkkViUwLUuvRxmhSb7lVow+apdQcER
VWATcDQZnMh2tRfCbUcYFhPKFFVvbElsNXPmurX04YmuKPdAFUWMnw9xXC4VUAhA
dEQ0M35vJT1aM+5g+oManCcqhS482fMujgUaCpnSmaxe4Glk7xSSS4NUWcFZViP5
Tqoju26+tPuGdK8vvzMvFwrRlL7mWbOOgxg4L40RNXYrRVj8XbcyJxtJJX7MXcUJ
zrqXB8sZ8thb+EzdbkomyPrSOa5I3zYT/5ymj/kHRgYEBHcdI6HdZCG3FmsJObt6
pAk2ATJ3x61YAslULPI6KIH6vhNs2zPalMh5BVVxmajexLsi/z8OgyuHreVs/Gvb
1uBkxfM40mwCoIqOQakqCM5iIcMfwI+57mjY7SYzeLSKSmfPvSi8POKtT9XoNoeV
emsL0EvRA8lDQilpyNHbxWIISiVQlbOJ0IcOKpnl08H1DfzkBxRQDnuWnK4h3Jok
u3S/7F+cVOFDHwvwDH0sI39JGDUm2ZsyIqqvJiGh7uTbxTN+blnijXxnYdW8NQKe
u2UOHA36YK42vHHbMVWMoLHZCKycb0tNPEHo5I+oXw3H8mZjJj4zJCFIe6xLXvR9
sxdlaKjHDAqk3lN+CElGASHkTJTZ2d77u2z2ChfKJWQSPqwhPNJBwy/RUBlG40kK
Y4JVkqjDB6sU5QP13TJ7eF9I7LZ2HJ8zpnMjuiwYo/UNtXQg5hJWUsCaEzvda3NG
5x9FFqMie7IIwjo9D8e6s1G2wJjEOfCudgguWEJFpGNO+EJlMRO72kyzqxrz3EQ4
36EqrPqwOYUrKKo6KUyw0CjpV+hjiH9mGWDShgHQChtcOyQuqliFSmx81sC71EXf
Sct7S4bWPc84f2vBPkfoJr4l6JXLuIbjReUtKZZuU4GM22SHdLj/m+2Ugr0k6nAy
ORUK04cxn8316b1MC7ulmSUGgsm+56YTaHdjiokFjfMnuOuQtA1AZg8LTcrLAujb
cB9GDqhzKVg1+RwusL3icjUFhLRVlyk4QHOXtMPxbcpAW0ZZHErOtC2Mh44M/8sa
jW5LPn5sJQwU7kdQmuID+9Kxmpl4C3WNxTzQU6uSTlZ0YmNrWrlJH/ZFI/wuVu7v
kj+bVLDsuWptrYG3R/xqVHcsP3tHRq2J/2xk13lRlcpGd6BkuVncdDfJUVd85C+I
U5NHejftIaZmJISWumvkFPkNQG19Dn1LVpgF9gZ0mza4mQC+1N/IpjrZ6t1HnVud
qPn3sDL8FxBu93BXlWgcYcLEJV3LuU3hcO74dhtYxZe2NBkLsHUliHmBzDDtFHxf
hcL2gHaiuJ32X0c2NYdyA0Hdy1mWrRtZ8l4fVLu802Fl+7JwweYLzoUyJZuX8/lf
W3m31i7XxRbivtJI/fipkuV9rzZJcGoMe020tt4cDlgaR8yXZxHSbNgIo3LUMR01
tlWH17Mn1UTTCsrAxhVRo54ccGVH2i2S677NH3xwDjJu9BdAW4c6Q1yoqp4Jifak
KJivdURdZ3w1bB53vXVICagN23sQPlWrZZOJgqMC7CQK8XpoaI2MF6jotW2otgzO
xzlkCnDwf4myPl7UOarMYwFWCWXppACwKsthSous/FRAikDmBoHt/wGahu2yzuav
4ErA4BakREpu0jBG2RuJvzAjQ5QHwmT1PtMV0vTpBwySgxIcuJUa93xv5DvHsVUo
uHInJ+22KgD4gHPvIaNNIdkQVq9QWwPVrWtVlzHge+e3abb4jvVWJIuFuulIeF1O
e/gahp6nUNQ+3K6s28ztML/i54v4G9cMpG86q+uWqMUR/SHVt8ifYpWa+eT9tkdg
taip/P56V/iKVk50mHNj4pfhf37Bb0Jv7WFNvu+7RUrIOKENtGXnEa7ZQBjZ5K1x
8s0DYd8a7uT4NPrX7edQStv/cdX5akRHQof6cyq4/Bmym7lZD8icQWRyLQ7Y4Juy
qsawYJdvAml5XoMAF9wA2MngJrxe8ajMsL3xsLlWS2FhUPNlAistIahm6HtSRncZ
YBjxw8ytyXO7LI75KD+VWc2zrIqGUeRBjwBhMvU9iivixMRXI0IagtGO/4vVzrpx
v3orM4PgMNbQR31+T8OPKw2W7Jdf4XpgkDYIejc5zftyRVgwc7wyDZ29p2OqQqkA
V6dJeAK5Alpv6TQw8hGpY9jXDaXshSumVtKEalnZIiBgsNSH8plS31reZI+slBNh
jQK0HvlOBg2gewfRgG8RnP3UfA2/odrXnQHsYZ6laUNYEVUNlbfU/J5O1P+pHEx9
y34LIpbeCX6a2oBrNJdmcaHKL/aZSR33Id4PTZIM/bbsLozs2IagngzgTlM/ir/5
uEk5aEFogeErS9pEG6WfBp+SXawwjDrHjFmby6lNKAgzwkDRsvlzqOLVjk+2366A
Kv9dl7S7/FF2WYN13hhwJ/3G8YtIqOfOC/goGnhyzZ6ZktqISaUcWtb2UeveE56u
MAY9kfUdBBainPjtIVK5w3x5s/fn5GdqGF2u6McB+zjvpWvQ3jypNWebIDeeMML/
PDdggCYBF0Mt7pj8rIGBPOVcpPQuCSQzRIvKGQ2e+mhb2CxK5Lf6qeD5W7JC9SMa
2tD0Zk/+qDzbYNl4gilNATnjmljn/Dbk841HJOhjDYfBESZjurOOasYv4xKcnN4/
oOkpe9RJqsifSBs9HKzCdpu1W4qCnYYhmauMhhwrNSOz4xzZX0sKFq7x88qWhQ2y
4YZrdjf8G2l/UcaEE8WPFgYewnNN9kfV9kt5Pi3kS6oHnKxEQIVv3jkgYjDn7WX2
mnqoEVgxy7gzNqoy2rJbUDDdBx9tuTUnpMKlI5AAl61+TW961PwkG9VfkZYWqgl5
GQmmdgXosq1nrbYHrQjth/WzCBQBtQUWY4eTDtNeQYEaaKRDDtlUuOINeOGxDA6U
KnOtpAbOac8xgttt4P1PrtrJ1dE5fJdp9YSj3Wuggx9rBY2DfsVitfAWgqCo311x
wg03g2CZAOeWm7hNWs8BRa6+2LlJ+eygNgmQfFSlQV4ha5EKea7vp68w7ZD/87Z2
kAw3b/8JGb2MbEcKk6i+FWWx9mEA1gxjCQypX5b1PlDXI9CSWJAAN87fIeDw+1eH
SJGC2+ifjg8RjdsSgiTMJgIhiAK7dbJ8OCRhd25QE7o8W5KbI5aEBuYf+SAMJa7L
8cwaDO6kWWrc5+NO4SwwSrEprXd3DUr+6yjIav0RelqxC+FitrmQ4dVfpuqdrTCi
A7rJRvfhg4+dQFR9QFNowpfcS3oaw4ZAkhT0QP2bpMwvh9Xw+uYCOQ3nhAaXvzWp
Kme78xiBlJh4LPapxbB8q7PCj/gRn+R5jWaZQJ+qz/IqgQzYd2AWe7Q3qJkeDGfX
4tcV320crM7YVY8Cu3RaWN2U0ME4gbda1ADFu130qf8G30AS3dgVBWF5f+Lt9Jtj
3nJdFSjiDPqpWQ+PHnXvoFRvHR9Z4T3Ct0xTUNN2yTvRY+UrFT1AE68k1EI/GzwF
IDczRkEkqNWoa10pMzMcfFKrNbnT1IkhcV8203Yfzjm6P9bV5NClS6wNuoW9XgLf
XuxXUxKKnPMbUXfGIWd+ovK9Bd9QInvixOYA0UMw+BvhIwjzjL/IJdkRs4lnhDf+
s/yhgRDdX5vTz6SV0qNinzJYuGsYD/+DtZLn2OKo9ZLkwaAE+NvNR5norm43N244
f6CwTFzYjIk2u4J1YNyOahD4YkDQNcfTs+8y+kXTUR6w+Sa9BR3OZK9TeH9NiLUz
XVUGBWOsAuxCztdziOAi+guKzJCXnTY6d1aixUk6yGiS8Fc6RoywMWogDAB/wd2Q
ICCRzDqCUhb8Fx8rK3dBtmzu62PqMB1tWgbV5abJ4zoJqSE2fHspbex1j0wV2TZb
DD5lcGSVp3nGTD7ivRsTI0B+COgcJmevmGx4DmQKJ4EQ53Y6CoPKdQBATAwXihpV
NRcm/m9k8Rj9DsQnhvSgpVYre7sY8TvWQeuTpABOr6OvSj4EJgjyh9TdPc8T8sdY
rs48BMmrKiYqNI76egJz7Yf40sCVpkxiDlP4IzAPko7HXWszLCTc1Grs9bwsBWGO
F4zuwIsNkCxb8O5zwcYRnXAslo+PzAvIgU5nErnCP2ElCRZ3M82U7WlNwCk+dt5x
PeECv2kgKSVGv6KwZ7Ei7hXf5+H7KEqlG0KBQVW+1AEWG8+g5l6crnU8rvMJ1b26
77MO//D8bvgf/pcjXGEAobLNEoYRgY0gma0pUzENKGVTuKtBG9XUfDJA6g0GObGF
NVGuuhaNhMoVfW5Epm/lvqsd9lg0EmxmvcfmEutjbq+FJwpE5g2uHzXI7kKQ6coI
XHEivJkXguxjNbWY/cy5FGDrr18Uo5O4IyyoZBExUrU1x/KDLqb0SekEPpDj6ReY
eGpIMy8EyksK8CTsqzvgWng1nXXnidI3CP2EHYtZOH7S0IaI55hQK+ORqqzuuul+
zTyJEEUd9Vr3M+DtRLbgNDcBVe/VitOngEV1kW2wwJzqVg3e2bdyPpKOhBfNWiB3
j8klYoUnooNBXKHPCtZgiYcfM9Ck/HDWg2RcqbTs47CFsj7jByrpT4AYZDumbQSz
PMo3fvNeRMZr2tOtghYQgE2gP1kL38BUIGL/y8/8PxF4NBI1koLiVFkfJqJ+nzKg
69GURSkd2kphRNwcZ+/X+Z25MLiyxJUiuLQBV5XPJiJ2yb7nxQFx1wUajv9aKPhN
MENFzr6VN+9yP02Sy9WnJNhDNPUBD2SMWd6rXgnQmKeXtwxHux0QZyLEkU2qwbNx
muKH9efgUNxcDLVX3pk3vXB21skRMv3kYT7kKqRdrN0ik+mJYMeBdNch3uIiI35q
sEeN3n23y8HthCcA6sBNAXCFB2tnGeuV4Iyd6rf4vFtHpnJqCS8d9BJqbxtjW2DK
ZVRhXCY7BYLPIFde3qGfxpy8cpI8qk7zH0jxyz0sArE2PNimpH5liiP4a2W/HvS9
HtVxceB4Gq+Gg4ym9h4ariDxFJFLhNTbbLmAiKRdBSOECV+2ACmrStl6wuNjWa1y
75v5j0q3hq5GG9JWP5DX8lEd9YQxTSEtKW9TnUNPGM7ap8rEUDopixQpi7eelxSG
toNS32i4NnsTDH0NKO+iOPKntXivYhLnxSxiVMeoSUbc4MQc7UejN2KMnb5GOT4/
K0qGluEnCDRe9zLjsnGBi+JjBSM2WEem26NASXHYEOu1R2os/XIeTS33ju++Ow6m
84c/BLx2KqiYN47Un18n6JlWBWTrdcAHUHE//R4pt4SBWmSnSmWy5iH1uQwnFMgL
0VX6AoEph++zzgmz2RMoSd6CJeEWnZXhCJKAJ9UrWvwS7pwiu8Psnd/g8UNqZPPA
//xj0VT3EUXTRkApcYsoOm9wEB6TPjtNcjb9Cz1UDk5qLQRPHDrseiRmmqkC9aG7
GCFd987fcaYmJcCLOC4pNKRqtr4pm4yfc8jiV0+n+9UUB2ZbBoaKZWuR+n/+9vt9
4HlLCA7l5f7dRIY3NnMImjRom3vbK2pGBSpj4XsEwnWd1GsxXbzD7kN3Ut/dOhqR
g4kcGIhAH3wm1sdpu4AISawaV+758hGfbTiuf70S+V0Uqts6f3Ybvvy5RwKitNP7
yV3zcmf7jodDA06QICHkukI93VvyNk9yDPWm61EvgffQRBwGUhvAxwmXSNYUfpf8
K9jhl2UHb9Jput0V83LWiUoXGyTaQT3OamXXr0ATovDx1RFFsCbSHe5ZgMoNJXfY
wV0LDtgDAXzFgsE91GtFT3sqe/+TBNFhemdXcrr6WYkKN9uRL2Cat5RLeS2GVrr5
kg/EwINGOq4UvMzmIOu2znshIAQyF9VbmQy5PdGexeBXIhs8Xp03tiTjZTEOiJ7g
FFNwcZ1AvgpyOmvjpI8CawoG6s4MRTFuIGTIwCF8Z/QTxucZiwxBAOVOHlDt7dU6
qsnf459eyGQLQSp4qckGpeHCF/+mul4l78BJ4QK+ypU5x0S6dzR6uRaI3pRNhdX7
5e4SpOs08oZOPHj1C2NL96wYuEuFpNU3IAtAPv24/ghJ6IEbfQrpOG3rxe/ZVbHJ
LbuIxmABiPdSxA5WA2sLiR+BmGvirwlvTgTtoI68in+pnrb7mLzTKLdbhIfm4Upr
PE6hRVHGe8W/s2zYO5cd0ZAf5Dl6fn9igDzKbiTtt6OZdjv+DwEIjOIezWo8KLKR
HMkqfXs36qpkIC9Cfs1PXltQ6m1S5fefwp+OBaDf38aI857FOoJ6TdM2w0wyL7Mu
W8GrH09epc7L2k95VXylNe0qFmGbWERvvRMmTklVFQwqMBKTYBezt7W3g1jjKw6Q
xovHhW+/FFtKKNMi46+ReAfK+oi0PKf1mhdIs6lhUEMomspXDfRBxa+5uwwXhCcf
OsWtp+Gk21MmiWpwb99gxhYqdQIhPQEURGveEKy010oAAb5ia2+fB2Yy+Rb6Qnyq
fMB/QOHsv1WnvfCeWvc1fD9Lm+aRZqysaVzUxzIrEVH67JoEy9EvWe/kWZqjS2di
xT2E5fBVNeu6EKjggF3UtXyshHp8pphBHqCo72/dQiXF6RUrpo7Q8ObHWbOtbAiy
GAGUball4bff6laZO/sViUYLt1knxDotZzcqk2yf1vReWqU0yGGI/dnwuIQ5jA83
dwk6HrMJ48CKHTo+HIOG81OyBFNOrI4uRhV6fxy+LKw8k+eGe4lLET9g5J5VJP3G
tilLlk4uCho3nxZ4EqT4054R3mUpYHBOUQ93CDt+RE9ZMCm/k0slIAWyXOQynMBZ
K0ueVYuV+04tMnnWhuvaaFLMTp1MQliWhkGblGhv83Oa4GHOrAvjgNGxg0e3/WmL
VONH426El84DZZ746vIk96eOHIa7N7jDxdiAIhAA6qmgWh+p5D9Lk8Cm3aDZ/wCY
UiJ5ksVKPZa3blnvpBgoOiK9Rzqko+MeDtg6HPJwcMs51L85N+49Tn5+muZNVHcE
dPB5e1LB/E+yrCrW1xswyNIX4mXJ03TetkleGOlHk+FCbcfZrP8ZBTMf8a+tPtG4
KWiZorV0RzucEfthZDLOc8zgut3IoH1SxqyxQT2ZGjIjUni/77cellBAYiGPWIVS
tuEEBZTNVmckdkd7DQG9WZg/S+ObPoxl4cihQxKE910qaYGwlmGw+7WSN802I28H
kTokfauwoSDwhj2ofr685vMqjuYfrpqyr1DWGS8OxIthZx5N28FU8iY74sqcXaTx
XvAd1CdQhqBdGT5B7nOBRdjc9l3e69ZfLTmcja/gAiwLv9LNXcuz6w2+yrTdpCQf
BMhOO9N55HPFRM84wSCNuJItfiXCORA3iqVofS56olN9hToBzshwyeO1b1UrT2n1
6beuq1Vl9GJeGX4KL1HXW9GB67bMZYVhusHLugIf1IAVdHOajogy5LQbYzGxz5Nq
y3PFE8bc/FXq+ynwQMRzuIZT1Gc5PmoEs0yRIdPyJy25Ltnb36DgS/zS7+rw79QC
Mp7v+9RwDGc3Zsownvf4BoHY2vzBFsnYO2hTZYIDzDBEz4kxoYjKHbfEBN+C12Z5
dPqJPB26ZvUgpeFehC1An3S5i3KPDM8rPvuzwl3+C7t36i7bVtmcoBsED5j7MZov
koPv5cL47EccKeb7KQt7ObpJQ5xEHWtkIkmEncUTmBxc9T9Xr1N4S0LwkCr7hDnG
8+gkyxvtU+tGZVOMe3U3TCpnqDtJUTHjFOUttcLYgijS0aJCnxknKFZNpNTvc1KJ
+WdI7FHJxCCWz8OcBWUJIrb+MYowONawt1k2pGFqcs2OvTcYqrZLwF4zAnAyV03e
RzWNWhiPgHe3mOESRU/BoJp5MLDWDtwGpjbIdG4XNXGmYztXtyzlrJiffQb9yH+a
0+mjuqijSrchpx2ALKHFqGMwysE/xQs3JvzWqRTMl7bbg4BOlFIIaJK2t9c6VZb5
kS/KYzfSp3PVUrIXsybGYhCTWz1AbBXCWSk8Xrs7jWoeJ2JurptV37MCJr7tcFS+
kMAtNxYqGF/S/bxgImU5uxkdqbVxyFtEENJsupeoSaMR7U+KKBNr5m7pPXMUk58y
3/r2pr/orqpcEJOrDQlvXMrMIihpmIV1drXExq8Rk5oqt/VsuB9D1DeAqk6k0J9K
sBbA731wBsEQEzyRB0fvm1Ha6Jcyi3C/SNHnrpzww5sHxRqKPd0qHlHK84QDEUlb
WjV4f6igrH6rmrUc6l9xGmVOb5pqvrivFh6bQjZgd3AzyQu0COUp4U5lZZxhvu+N
ov9FUXZUarBdmPcFldmw1KVCFBWQlerDKYZXZoPdypcMIBpUx6q4Zsjxd2cfnHpI
RrkEbLtA9nAMhlMH9y3yTVeDgB7BWlPStzrz8YOGE2SV55lwtH0/o8GfKlEAa6Mh
zbNWgpOwIzesYPO6P2lCOTsHhYN+4BU7HL1WPOa37hACL+HNQq/r/T0HkiyjleoD
b/vzKcZtVBmkTsfyoYvGymXJ1H1YKvHdAmdEzRdS19gv0mO8Zms6OtD0bq2zwBrg
3n6kA0csLoApgT4rN8FUYdqy+vcgj+jVH9+AGXxKmJtl8mt20ruGYHNewBSSiGPY
6AhI9HHRTaXDHizksH2SARFbeno9KJMrKMOoSkjhzTrjM8Po+O2DEuRktC0idaNW
FXq3eLf0HBhgDDCVfrtxWExIkMubpkxG89XapNtp0uTVS7YfEqu+cRRRiSMPXGE4
4hwCFvC32nZ8+5LAibHtI1JhA9YERUo+lMBlZBnkHFD9Akngp+jARsj1lchiwbq/
CfNpjpPBU+QesvcHGzREZkQXLxbWtjsVEO5u2XFmaLZUb7tPMfCVUGfjbUVTlnZ9
`protect END_PROTECTED
