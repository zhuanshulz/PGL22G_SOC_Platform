`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M9JukC/kDqTBVM/4We41UXE84recxG61vuaMjtSD8Y9pwebwdvYFwa4QhdF8NwgP
OQMTvmdT9NgmGqiPHc9u8NuCUy2d3BvxM4FxLOfYaX7B9JgHqSMyd5v14zAqeu3J
wo1QLvpP473Q5iGr2E9GtoLFynG4bGratxJsB0ZFPJEvNitJILiX5gpKNbyrlyNV
1CZW25KIFKUhE5MnLkmA0uZiBGPFDcFA9/5RgymtYWiEoEskFGOwezcoD4YoW8Z2
xpHGE0Fr3SCm8ej5e5P4oEs/656t545OF3xc5TKn01a16sFKbUnHkYHSfNuNu2Jz
yhNF2PEyn3RbsDNjSrs2W3FgQx8Rn/twx42NbYl4yW2MHknmUkNwrI4y+nWzHN6T
d5SUjICJExdvycpF7NQK/5uLyYI0bV3fNkkxHOKwvt9RVoEmZhFejdTFUh2Tuehu
m/ElJ9/UcVZv3KBqRUNaIUYVIRvCDYcKrzoJlajzBEvi2D8N96HWhQJuMPf91U2E
86Ft94ruAg9yeLvpSviUf2AUZlasid9rREBzm8P2jX0yH9J6gSJSHFPzSSc6/UF3
zfQkw1eYI+mHL4F7pDT4pEJhWpgIzO6MZkzBzbaO9A+6Xwa8t8Oc29beRDGWKgqA
gywy5IGZMgdp+bI3HPYm21Su75vYdhe2NZM0pnzzSc8=
`protect END_PROTECTED
