`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vXlxHf3bfBs7q7/l2QH17SIGsWkEq0E1hdXYEMBYEq2237quXKomIVu4Fkk09iOf
zWsNBCgtwEL6T2PWwhdlJh0/wwMf2hWf2B11UAPW/H/El2y82ljW8cqxi0Z6WnPu
W0NzsFXky0nE1f8hT4dhdmIXLnD4/Gf1BzUSnpFx9fKb5qGEQMOJLQpxl8ltTYg2
Cjf3VK7FWvdi5kLSpX1v/mT8c/hUDwwSBB4YQkXG+RhuYJYkC9wMS+2334rOYA2M
M2Pk6W/JetFREZgcXqBk94ZsEqa01SVYydryLn7uf2y5KNZPlSnrtXdpTsLLIvlm
LygGlzl/4Tm5sd1HmNMWcAJluW6bx7Xo2AOXCJiZlwejvLhqPgpTOvfbBYRsDL4L
ojrridOxqjVctwfFP1oOkf7dokMR56OgKkBHTFixRtjZE0RyhYdYw1Woi09ikMb9
piiQLc+oRD0Br2uilpQsozfAwUZ2MwjIWXla3Xo3zInM6N00n9tmel32HbtzDG5F
ZdSwvSIPqufQicoB/zNG5unULgupBdv67RDpBgdhZ/9xQEzvZu6kwdiENBf457kA
4dbBPHgDBm18o6DZR8IqVaOYHP3TO9vt+I6JjH4pV6f2mT0hP5YQ3zOsNTvdoZ02
s8YS9Vpy0I/EOL+LpmKcDHoP+olVABF/VQYApm0r06TQJNlqHTPdr6oBNdPGANF3
/xPzxLRq8kQbw9k7VRCBu5MI57bzt7VNEVHVgRW728pn95xBjq0BVUqdcTzy0Nd4
zJxn7nxD5ObO6kTUBEnwZ2rQ0jshHNdrZV5OBAMqAGQj5z+nvR83YnVLqqp6Vsdf
G+th+UFxDwhJigmxzq2NYk3GxJ3x5iqN7/3k28+DeAL7Q0XjqncTKVzRUn7eD2Kw
Q0jrMDnj4ImT7OjUko4ViQ==
`protect END_PROTECTED
