`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xwGTfEaTLTyGg3R1z9ymiAuAyF0iAHAdt4ehsdt5no3vvzkkoi5km3yFf1mERIme
ioqU8MN28+GiDY7YvlL7w+nmiVQiCCC/ZsMzP61Y8yCX8or5XCvtAlGThxrJ/54G
BeYCGiJz1sPjQW5BmqwWaNvQBzUTQOj8BFptJKla/Og1aE+6l9Vs/wBcRS4jKarR
MFnvN+qVIVvRT4AWRztGsK1zkmFa75brOpcXax5XwfhnzfTfMzagxd2ZD8uTYJuX
PMgHekpj+SJihTXJKokITrKBi6+Yi4t0xRqazs0KK16BQFYfJmEztwM5VXrGV5N9
qEj+BpZa/C4zxIArr05CL1j0s+07uIASSDVZjlH+RTSdUAy+Et51vs2TK8jNhSK3
ZEVsvr0GQZ8muqphgqWcImRFO1xOUMM1oO4xEvmJybpth9O/Zw4u4JPhIpZYj7HK
4OI8ViTEP+bVSYwgSme57dmyb7rohi5o9HCfBu+6wH1K4Bd7N3oLO7SHil11yaJD
dUsV1VCByzAc6MSKPwZKd+pdkUhUFZ4N2QRKphbVMyYKugqnhFj5VbAThqaZodJC
aHN0VuAFE8JdxGNiZ+E3YpDZ0nE+USKduYmqBZpEqe+EyU/KglGAIS2lGxKYCYX3
0khzfcNm9hM7HIq+zxJzgc7WUE+NPXM0bZC2qDwR+Y26PO3w5Z+NXakvijdaw26E
E++UDY8zTdWVjFCLbtquiKIlRkW62T5h5eBdVl+KAPdMHzfA1Ie1G7roTV3cY+wP
Y+DNZEbYJYggNZWhB+2mq9apTQasrgmBNd+Ittv8wr3h6RhfD+pCgA6BtkjZP54c
NT/tNL4e+xazVuUxddIlKuezbb61mA065maKUvteHuA6uKuDga1xPwzqsg+8m97T
gqEvo0FpSnqo+lEW1zoNS3mhjhhaaBgoaxSDMDGwpdhLIZkwmikdsiDZLHrXX2Kb
umuxVaI3CDDM/jAOzpWsuwgQsLkC5Khl7e3b99AZoO4HL42E6Jw7eAsxmc02vI01
ahVhISNp1AKXkZVIu9rVmGjnV+aRVCyajT3tT8ijv+eLQ0OtidkB2d7L6mxP5M9n
ifcClo4bznLQ6JfBcbg3WA8oRERkHq9+ey75YJjKOqF/UcaBbRG/dx3YNQjprAoD
csVxoSpiVXLjJwLT+DqhpnXRzD5lfwPmu8zDvgtWcCbpnVbCDunixdQ/D7RnMRE0
r+vgnPfTU99m4zSQApPdgsDnNfljiv0pNtdmV35aAeOFw97Z3kz2HpX04vhLq53/
KGjgsr+RIigG83JSxno5mNbPSq1lQ1D8S/juDrcyTHEayHsXtRY5rGb7OYELoQ5V
XIe/fg0ZYOaa+KtHI6A+xqliHEpFKrXV2qYQA+7aECOthR1aC5+zx9ACNTK16TXT
Z0JdNswQCfzazr7yp3FqohWEsTf1m6BaHniq+ruazDw9jRrlcoURoSbGtgCl2RD6
fEX15HRO5MPRl9aypIQT5/lW/vkQQkEUaNIQglXej2i74AABPjb5uNAQ8NOdzRF+
jKZGOymvQakQzcyVtDZ416joFeZ5NdaVqPmXiuN6C+s=
`protect END_PROTECTED
