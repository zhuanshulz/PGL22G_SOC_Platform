`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cj+pMTsO1LgGCluJtR2lRQ896udIzrjBAjppdQdkiJDTkmxpBhKFpBaMZAXYs90g
EHCcLt0EqZ3lY1fm2UjYLABkMLtgWPJPF8mVvYLo9mxSjUW4Wxllk2F5RLSVmMkT
3iPg9+/+PpzwPtZW8s1RQPr2CXkA4wFeCOkBb6JRD6RI13KxcQM4PTXOHV9Xjc0U
EYr3jdQ6mDgfKyIhdtTf1vT4mEMLquy/KKLw53W15wF2NuOXPWbw6TKXlicq3luj
OxRr5OWo34VA9jDpVvZTvkXRK3b71eduKzysdrAuI4DC8riIhm56WLoIBc6s3yM4
k1yPNkKxvumwV17N6q7Qv8NDsXAEWwoubUAuhlWikajIoSYL2xQWKp1V+ZlFQtvP
YPbubzfThqlzhF2xCvPj7nos7x9h+DoNdI7YhiSBH/kvkG/6dDDFG2XqxIdUxwRq
BCU5WPz233/Jbbx9E8swWq16neoaHpTVQcbopbPhiaCynX98H+NvA77acx8ol4oC
1zC9iReZz1woEH+q7mPRgp06Wj7t8ci756fn6I+bG0Z8+Y9QrENrf0Wb59gzPR1u
ZEum93sBkccgTgcEd4CjrgckpLMZA9k8u5o/OEpd+iF2otrPYoAUagola5u1HqVj
Q/7oJE15fRnpNRdpcPvh3IsrFkvX5fRx1fjcowzRbHA=
`protect END_PROTECTED
