`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AroDhw1FLx9rv9R0BHOHsNCiUm3O6/VQMggpnj6FDAide/R0gzVP73aB6hQM4IL1
/0rpn98RqbaA6gZvuJZHVROWt4R7CO6R6tPKO0HmS9GJHzyOblDArv6A2CMZA1jT
I2CFm3bau+libsgjnwwuORyCuvvwHY04HIKoeyZAmRjV1FaL2NrAajeGre78qQGW
eICnPBpOyP4GFx2sEJoPaNZjj6fkC2HwtzaFMtv2tszez0U8Q0/j5EG10La6D349
f7OQAAyZ/Zc5hIouf3aPsitNm5r4dvdXm9YmyMlLXaDu8QgC/bDtN/iyzeHmb/nK
PX+4DnkIoeQnv/7aEpjIeFD11Z2otXqLFBuB2ip2KnbXwPuYNGzyURdo49N1uPsn
OqBJIYZ7BGblwmuI6hfzftgz/tCdlIXd/YQWSs0hHM6Cq2mdY//305H4QI+wLnkt
SZ9QbNSOGnhYppKf1JhH9nMKqtUeFfFLO55WlhrvnQHR6FeZU0wmLhWxIcFouQCa
XA+d3obVkK3RL3JbCjRQzI+gfOO7/36mwJTUFwLe9nULIrhXy7HvWNxUe4PlfiYK
D4mpxsnSzM8OXAvULNn8P/pSXSFHva9WGKODP8qqUBpC8U3JYHw6NNEeZBrgxQIL
gWGuEZm+ooBnFoI8DwGjjwr6bGeYfxH1LdRDL6DOQ4mD4SBfO7FM+NMEwN5cE7/x
rgGlh+zVCReEWGN4AG7IDwLzvfLlqUdt6+CsS/W+K6MtTLgC6/MD6jt0jBMPyqgH
jkqwG+3ApT7P5X4wNtB+ItOaM5NRVXmpfe0gJ3Tz8I818ToTZLFFe/qOdgrDG7CQ
AC0pJLX6Njbl5l/EadvgvXwHV4w+O+o6VJScGq58YfCu39MHzdo2ZIzQRfNv+cw7
1GxSJ0zizyWvlhVrqZKRKv0dwX+5V7wPTkhWhUMyh/f46lMXAQ9u8BAbRae4fKGP
oirLQexd3MYWqclWRvd0tc1DbXA+gCdoImtBPAIyBCWYDecV4sOVes8JG3wCUESF
AKNPiCtIov7fcwQQ4b/xNBx6ecG/dyDWXu8P7LmsKxVAeYPHKO+TitElfguxBZGD
bzmi72Ud10Ox6ICAXeHHNgrsV4H2Y5bqLockFUYTRgXVuK1UxSK2XHEkEZOe0h6e
sJaguN0mak1LHROc8WhX8AveXVrzp/Hlzcyg5wQeqUhrRDQfg/F/nWlo8qn9xwFK
i0rEkufvDOtRJvYfkhbbKm4hFJdmLcTv2hMQ3+MXsAkT8ltAEVikFVi2g7Cln6/y
+S0tU2FRdM9qDCfkdjyEVpeWvvFUVV8TzKdTjzrb7oJskQiqJtXUcFjegtS2J4pO
/ugWN3DLlkDWIDVKXUBEQRPNiMfcJz2pLNy2uKzmLzaKuK/aRuOZa3aFaLj63uMP
9sbPMfyl1V5nLKx4JyHyo7/OVVsB01j4oORyPJSDicuGxCkWJkkLCP4LAhm7amsG
iGe7bPSy1lcpAVruynm2nlxgMhQJvoH03YZ4A2/b6fl2IVM9GaJR7gakMjYpngNF
L4ZU2iLZnDC8VcNxOEC5xRtaIbghUdOOhEHX0hu1XxwZiImbgmHnPwn4MRBytIfJ
zusbDFAYU2jBhFICkJnW6KzscKyEVm/XXmFHLBf6XxIjSLvFwIMMbAXxpKY+vluW
UB5PnhWfeLusLFZnlnJioBUCG+MK919ZlKGTtO3Atlj82kC5N1uSwDvsCvjAXKYD
nojwK7AJrFox2fbc6SOjAyf55tbHMd/hmOAMACAafjFIm9KkqghX9L4IKQMOSVfM
qd89AdFNsT1PcJ9ayIwK3tzqDYJsl/wKbT9PMxKVvl9UI70LIyI8PB7L7gNNkpYT
9P7abPURgOuLXeEa4U30749kaTH3DItgaDzv6IlWZuwJFdGc7L2BUa3Y5sfVFyNU
uE9p761UWTwxAI5jSbUluVUnPpc658ooF5Xf+k0TcIy9UowVDy1BJ76ScIK8UTAu
gEHgefsTLbUrxgyW7yXT6ovRVBD32naxQwUV87gP231Ub7oKEk1pQAxPRGDmc8zS
HlFXw1aJyqzlIRU/mzsOo2UI0sQnooXEQ8uzl3BLi4GPd9HjC09FNqHb4NoOx/PJ
sWeXq3ilQ6uOx8LYMGaY4NmBIFDvzaXfYUJc5c55PMfg/qC75VFsiPeu7bo6STXV
NvbizgufXAq8YTbNUn9hzX5Qo94x859+Q0gBfa1BcgIY5Aujn1mLcG6+z9YN75r3
R76KGOfX0B4KKxpE8RSGeOGYKPmCK4hLUNmAvnLi5b1xuLJ5IGaXD2CuB7w1oOWA
pc5A3u7HzdsAWC9MJfhZGIZ0/LXW6JItexsGpYUNCCnR7ZaYIbsNLeWYldEcXvEc
xRjLjDUetJDJ8zrOOmUh1gJbiB6D2FP9yY7ZUMG9wMe+bAp3o0DWnDwtN3Jq5b74
wba6mSaPDmRxSXvNRMN3Qf4BmX4pAy7Lu2LUSVKcxVO7uWKDFE33fAZrkthAiT3I
VGNRcKUm0v+jYCsOEr8jZLHuSbdD5MrfHtdGXjBiTSTiPL5/ML0pzfy9He5CPunt
fzLexSHgccmDNpUTZA7Xe6vRDXeytBx5TyciXneEkfXHTCmjEw9C2jtVhV3elLf0
F7heUaOrbfHpzqjwA3a8LLHc/Qi80gxDReugUlV9awJ2zv4+PYgA4KUb4rreB+qh
sqVYFULdHBujWjcjEf2xQTw/KonVruQrcUbqPCswlbmf83IHMnUbDl3EXR0Py+w9
oeX6AXZR17euhG8BTMqjjoysp+FU+erI5VhSfsN/w7+RgFenj/V3Dr+PcdAqi3WP
h92Eds5jxUGh5r3EhhOEY8nphTzxOlR8zUOY7tN66qxGX/SnWwZwG2tkz64PL/9E
PhbxkRN5e96d3jTFhqMQdIC92whatgAwYCnUF6KzczmalvVPT59lGDavfCo/IHH9
+kIRLRTJKNLY3Gnvcea/sqEFOaes2JGeGcVydPbNnpEI1nz3ufrVaFp7POU6FNaw
f0H98QRnJ0VN4xiDI2Qvu20Tp5mwLizmkF9BmEUbSbN3R1Xux8vW5YVk076hJK7D
6DtaF0xuUhuWQjtWJISZenlotwVv+vXG4SciX4BBcGbyyUuFa4wYF82k3KE+l7UK
JCqKv3QU08afZ5EOiy5CWR1WhnJZxeWj5QOWK0MIquMRsie8Z2cGKm6EmK1OnTVj
7a15r2NWOZxeZSOjuSbZe/xrkstJwthTVqY1GS6q2duYZhEYsNjmPBWZnCRDF9d6
exB1/N/LDo+Su+0UXWvHYIbj2U0J0WEajooVhvE+3sOeymEQmqKd055keu6rSX5R
u33xIqIecxuIgp1LG3tNKhNPHFcuFlR9DK1gKtBS3XAaWZReC9QM3CHD1JLJ117/
kYtCgDl3tWUm4/pv+GGDYhJ1DBVS/HvVWcFluXR1yElllnASJdDOH8y2qRMDmtWK
ITgQ9tV4+UNGY7cW7l54jMXqlU34dMdxwXhK1zFa90imuP8V9vJLeectX9XYzzyO
HZLZGYjbLnfveS4jRzk1A484ML5a0RS55FAJHMYX3s84hk2rJ29cnjAqIoPf2VXT
IA0ndCnNeryBX8FL18fyDg==
`protect END_PROTECTED
