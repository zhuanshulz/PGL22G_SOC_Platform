`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WFUEs8SCqKlaDma7ZGJzC3n2CvvZij4g21rMyW7YuZx/IK+ArHWx+iWC7RqGmTc1
hChWp0Ltq5jql/tlmEOQNMoj3UDp+38E6Cw77IBTsqRvnfu0SLiqUp4wudj9WA3k
WBig9fGMh+dXKKMLQcShgUcR7hgC+uVS5kE4o0nE9cKXT40kRvVo/8ToKO1iC2Lw
uCwgGWs6HU+vRMJFeENfgqzpIdIWLHxJPPwR9g5W+W4TeIKYQ+b0FZuzWZ5lq+/H
p1RV2gwuKGN3iI+9vrTMGlOoMzf6I8DnylYDJulfQAIw2EdXe+vfm+AjbFmcIhqJ
1VVacXK9EPdCaKGJ5o+8ce2O9SigOLXC7ti9NwftCTmsCHJEc9AKsklPyluJpJTl
/ftt/pL4UAMH4KdwSn3a8GkOk1KtpgSHs7Epa+eFr+11dewNC8yPQHFkIosIiUgQ
Blw07ia63sRZiDj5ZZ0Fh5AqN0yHvQH972BrG8mjuL6pDqJymXNW/9U1kfHS15o7
CPhOsspCMigg13oWXLbpzgAMGofahFwRwK3YEnv/xzvbHq17oMUz7z+BWdjwMgXj
QpzGQ3ckqc0Yxk1WjOQ4O6vXyZw5nhwy0bEQfZWwZ3EtEGe2rgGCpj6bJWUUVPSP
m+5MIuv5tlIyy9vIyeFAHUu1AVYwsOmAzP0bRC0y8uYiliezxdE8fc1XaYpwy98z
Tp6FFy3XXndSN8XhQJuNvKX7GBpawOjfl/xmVhNAkVvH1xdHGtyeq9TixGlmbVPu
6sIciY+V7tHFWMnP9kSxboWIwC3SuNhzCG/xSdrtKQ/aWX5QJi29IPPgl6uhdQv0
0zv7FCPgpZEDvjdsIxffePuI3/ZAQaBQV3vA4uFtKy8ydLCYaotEtXoY1l2MWTON
GuyeroJVWY55BiPJ3VkIM/+rjE8VIk9e/QTUpQvW5aSBlOKQ12IjIFYChXW/22EB
gyYdU0Eo8vKGxAd+pFOcMoYkCqPCSkamn3+R7v5ly+5p18Jnm3MnaQoNpDlWzwkn
uubb33sjUb6ufFq0DtmWbodfBZ8ohh8TOSC3GIW431480+PhapffR2eoGrvvYQvs
0AphQllYBN4Qi8Jmv2QHAwq4Q6IB/dQWsbTZLs5YDdrkoNkv84WbG/W8MqWdMWvE
q5tWuAd8Wi0L+7obT8Gz3zK8a6w4IF2zW+SAbbYKxt4/GPgHj0mbhqXxV13ihKsT
OksB3PnPVXlnQHPspOetmuBOmk4lf7oFgpO5lBcTwYm0THeW9rvkQOXyDi+bu2ZX
R1DfFpte7CeZVZilKM/KsZF3+HigbfbIMzetYKFFsK4+s3vVnXeHpxgSguyNk1aC
oHr0CdZsG7EZFEuPUt5Aak/6wHByhAwWCTsRp6EzmJk+0LLEAAPWzxEo35tPvjdX
STqnBebAvYfxzpz4TobKJDm13pZkzY/mg68XrVxjKdbWQ+OYgaHQiCKVkRpFK1qT
vRV+b3Lu8CMb0tH01TRpngiDBzaruSMvGzxnukUbomKFMihi4BTD5doy9J7RHpYa
qz1Jnl+DxhYSeY7jxan1wErUPPeRYnHstOiIfi77FY4tN4Kaj38/n1UNa6zFXm+W
AeJ8AmEqDPB5X4Ggx3i505dMFxkPmW583seQKyEAR74751WxuMk340Jqdch/yPgT
+eG1+lJokQ4AK95/AYDqJf+kCpa7aTahMza7MHYdh5LuBB9aj0MQ34ccc7hjzP/5
2GyjHm5/Jhe9+N/XAQIWssGEqBqINl7NE6AJE5XLR95ALA+xI8ZKM52r+xfZTXt0
HO1vc/BTnyqfUYyljQXw7yF1VIyBgOb+ohSV+iTvJ16ZwBw7bQcjlGwUkWBD2uYB
ZmSYRmx9P2HzCQihlMHjZuJ0tRyVL7KIcHCfqh8caHcNt6JJj0MZk9evpEg+39Nl
IkBNyp2/HL5j1jPak5iVvRauuxhDv42ugYOPVP4KtsJZSD+xWWmVbVD3s0xxidgk
mnyKEe0T56A7QT/YW7G6vXM4SRnxZ2Yi7FajjzO561/KLlkFuw9gXZFGnn0p0L7J
N0tH9baj+EAUr4qzwmlyhstDbcT/sl79PAhHY19r9ktS34e1GETPqzjaDUhtRFYv
uNWU1F5RfBxTGCXkegITayzVdb0Jx9oEy1uoqn6VuRjNSUP0mxDE4c856UjRhAQk
ptQUoWMOvQNlb9zHsnSrJ6S3i/8SMdtDwBnubf3HJde8WcViZmMwUgXZMZviX7MN
/wiUQ7d2kXC6euwG2N5BJVqKmfZZGdTDJONBytdVC5E7iGkCGrzb5MMDUesFnIvN
Mt2YD7InvMt5zPVC457zveygg0v3geQjB4ytwnFQ5YLUnh7NsGbgPV1EJ9OoWWMO
`protect END_PROTECTED
