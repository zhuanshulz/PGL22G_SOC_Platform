`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q9L6C1uuuF3DhYEVyinTKs5Aiocvc1UvCHz/k5t4EcbN5sSJXF+1Dku61k8Wy1Te
3GxqgtvRfqz/dcdYtpn5IemOXobb/a1TmMHGRDGxP5TlzykehWNx13TQ/B/wT/dr
hcKcoCLs/6EgKNS/bItLpZvaRqtD33irjkmpWn9b5D5gVPIlLjIZIDxgdM71pYhS
k+qxZ8Tn9x/xpFaRyZXe585VjWtvBcvf3wrEglVZNZMDu/IXLTx8nUqeTHGj7bj4
PaH2K7fJZq4VYSpeHn69QDed46puhNWcjqCLvuutAM/AHlizL5jiwhdwmKYHuD2O
o9NLD359HyC8PWsvs9FV2UqRiniFWRHzCm6lB3DoX/0SiRmOvBE54kL/11l+L74h
whF5PLdhMQfkPha2ZmeqvMhluFDc6auXipaCoOK7iIE3YvbpU2ovCtoTaUDGakGR
wo4QyXJITIUQ+PP9p2125n0KjEpzgJf3q16YKracaNoNzniDXcEhRIfO2pGoM5B/
AeLU/Z/yBA4n55cFUBGDueLFXTLZG1qczoBUY69zi5FowjeL4spBNy1cegqtx249
KDS+rBMqMnbav3t90mP5kVNJjK2qcmVwzN9Q3KI5DYmWkq2FoLNJKzut9UmqX/Ny
9zcN0heqjLKCJuhZeDC0+ewLtMnqVhWMS9VECLnqei35Zj5CKbNDryUy2fTd/xoF
kc7upHxpqLDgiMoXr8+K6jatNsUkMcW6IBe0lq/PygO+Vf5b8rDpF1UWioJsfEmV
CDrDSuhagYt7P22MvdY7H5T6DW7U7BumqIe9y8lg20lEjVzoiFEKlMGUblZeBnIF
`protect END_PROTECTED
