`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OAnzmGq3Clh0nKiwKqzKvKMDSYKUxCr7potK0nY3eQkTRuGVjXWogwzrt629whiW
yDyIz/wiEcK9oAJ/77/FjTzLbynddSBPmn3qx8C4dUusbiZGVYxKPLqwrah3vZfy
ksgenNkxLwpRjntaaifilqe+jbHbDz5EOyLrbeZeT91iR+AellJMjq10cEBrO7Sd
UMAOqT6QwKChd6cYzbxEMybUC+k5N09FgDg2Ja+Ua5PT+nO+XnbNtO3skKglxu9T
O5rosod3Jhf6IRQdFiDLVC6Xm+c+YtilXzLNEFqkhQCbYzTvF/yeWlwEeJP6CY7e
N+MyA+9/2Q0HrcK95owR8hvehbbGG+A9hyh7jOc4P52ShK9vQ7FnEGx4k6eG58SN
q/2n1fI3A9tVY1pFBeGo9Kus/nBc4UtCvwxuRQ4bfN+KQIR1OOMV4cA3aU8uvW9D
cqHnW0tzXRhceLjpFAUrKs5M5GEycQEltu019hZZv36IrnjoxGPuwUewnWUH0pbs
EabIz6IEiuM4tj1nIrk9W/59qMaBD+65WJUWzzKUvn7B9iuvVsWawAaVP80aN73T
QqKXif+I7cr/tFcRiqTgm2vdxADjik0Uh8+QNGHt7s9FvJsSooJMeyLlnoGUOlbm
6jCX1N1qNMNT2InXfYpl5ZPttornakKTy0yIoOSnpiBuV8Er+aBRf4LmR+XL7vbj
twwZt4EoP9fNJo7cxJ1QLQjOCcMSZb6C+TcQq18X5Gql/edo4HTlhhHpHzYTNpXi
whzNono24DebW8k+um+/8I7PXpynGeLfN7dpH/eadqZ/Q3jhzWHFpXZfrBujL5hk
2J4XSHmgh87KKfYuOPsTVyImfPbvDKPh13RBpVMnf5kpB4P/QGiC+06jFTjmOX3P
zRUBefXAh6KNjZzjYIEvrwBSRkAxNG6Txxbf46Zw/JIDPtxuPIOnSFzH5cwufgff
Tg8m8lfTgzcIJfaNHb80/uIOrGWQF5Y+VJLqXxLf1ZzueGQwI4i1Ou2equZTV6O8
st35baGt9WrnAp1WvcDgJ6YlBfjjtsH/8qjm+Psb4YCNLwCWXGRJbpgUKBBAoe0I
wR0G8UCL8a+S01OtEwNK9CGVSaolN9IQAOfdrx8dq9njOkkdQ3uQgwU4kVA7+3rC
iLebZn8sTIeicP098nq/+++rGMp87qss9riaBAz9Waf2VyuZWEB/ffX+JoLrsOfl
ZZ84v3vgzu1buquTTxNUgeSCNbRoACCrwhUbNq/gMXYvKsR9fDChFCmgMITEpxKR
J3KjcyR0GETSClYyvTF9qcvxXGOlAc4TQZkhZckVm3omGbeY8JQo1orr4g7R47WX
CiYlCuYzQCvmGh/4BMEFvm/SpfXxXvfU8AmrpRY8asqg85JeixPdCzYzUt65H/hd
2mEt2K0TnO114RzoFujMsLUu+pELEEvIQ1Zn+s84xLg5U3RJxSBG8ZOe4XfVPTG1
XOYyF6qwugDVLvQa2W2eWg7lODC1FvuTIMXiVMtjtveL5oKpCySHPpCjpq15eAqJ
6MNsG3xLIkEMpaOb8ZC3p77RcyJIj/Uv2Z5VNHxEyZOBHzH8YzM+5q4OD/sb8NGP
LP+XaE7gpErb5/UJEJdbbtg5l5k931Mx9BjAy7jHzA5CNiR2hhbXhtXN4FtPqFgm
Q6/El5LmlvHzz0Ju8lLAtKsXQnCySlhpQ5UieM0AVo0oAgONgmGcm7oTgUT6ge7r
STl2Ke5rirXjvHJmeompRbPr195+o5vMrNb98ZoQfIgcVvL98Dv2sxfMUGEYgBye
ag//c3F8lrHozUp2KPkOZPfG7hXffIve8TmCvOqdpPClHkVBNkJ5WYiLoBn9MMe3
Tha7F5DTP+/fll5qKwCpXeD0IgJ0qCmUDgGxnRXorBu6bzvUqrmCJWduT8c3VdZR
0oQPjlmqiHDs8TZ7A5G0GcKAxErs4FG5TdnVFDNHnwjACuGm+c2Xr/C5w/dw6Vfy
aGRidMwPB4J4v30bUVrO3eVhNOOm3/qQ0PwTb0f3TR+lBOWQDa2GwoCVi/vAsQTb
9glaWoJmldLHDmz6mSaUxs3qJpNDMgre8TV0hrLqgxB4egSkz8KT3wYkI9tSti/L
NwgEyMHVPabve7euk9t54WUfs/Wcs1NCUTGnRSvPp9ddqus2H/eNKNG9CLSVZonw
ogE6chC2xsUn10JxfdTKBg8+x3w9SqSxn/21oM/y8dwbVkXQncTKYLRT5i//Isft
KShfWzlhODhUiG1VX83t6TGjmASJD9LkWXuUnQ8Bs506ZMdgyc7TpMIaNpE1IAYI
jSxyU4SpU42FUfr6gjHU5hGG5tjzrhxdyDoiGtWA7I5CsWZjGm93ecizmtMDm+l5
PCFUk3NlkTxV2gu2WCs7jbp4SaEK1ZdwSPjF7NSU2L58Yh75IagepToYN/OS2l9W
RafTuAnp6mjLsJ9cBAaKj/L9u3ebad7fcyn5FME1xMM8DDyiRDLW5CeQ/9Zexq6I
3XLRhGVP7k/frbsBaPYEGHxrC+GKS1KHA5W2uIv7oiYSpGmXUw4KZxSNUiwWrDG/
PUG/dNLY09w6+aIQ420gKd7lLlrwbKK9+Jk7PHlTcoS7J8HekUaB3qt1aSXga3/m
D6g2SKgbq9KEhFT1JVRDjyQ/ROhtCwl08ZS6P14SZU0RXg5V/tZmXiHZg4jz/Pif
Y3AJ2eNGCy1zxJICaP4RezwaOT+Tzh5hnTcUQGPaE1PFNXzX0TvqV4HyyeJJGNq2
IlrcwXyQy8Z01GsB2a04EVNvOp5WbvU+D/qwTmsLrfiGrgqCNDy72pJI8cgkGwaA
qypJVvlh3m/mZdv+NbpcaGebCvwWIjtVsDdMCAIUVzxpSATjoTCCteb35AEAM0DH
FScJf41kajJUXGNi4YzpDbPz2Owi56HBj5F1vFLmwaqWESkrePdtyT04Je0tlR2o
mYVp2SZaPZADAWKdfXhg84lTN5RgDGWYlmHdXCtqrOYY3bzj1pwwKr8ezpP/2l7H
GyqBs3oPvO//1GmIRApetvTH4X7cgOde1sGMucCHax5ACN45KlVMs4PxRpf4iY7U
8uR/NU2KXxxapK1A8k14LUjjBPbkHy+7Hiy6i2DaPckXchY0BryeJp4ta5aq/dmT
qt1Cv5sgnTBfUUAP/S9CLpOnttEfdHsiXAIl98nk3+bsP+/nUDx9jmHG5wdZ+B8G
RqD3tWi5SrKaTCC4qc5aMSqMyLDUywYghAqk7UWY9l7zudeHKOmyIAudO7Loz6OT
PZ1Fp3mUNHZefWqA0fxk72L5OwG9lhI+C/dJ7tpYSgKpzFd00OEgGSeAbPOkU/9C
rcNWj+TW4qHmQdGh1aEz0wfIBqcqtvSsR/0ivRxc43oUQRfHCzKqUFUtCbLJbc1L
cs0zHeX6MZQDkqrZkaLlyiIur1hhBxqkcaFGsmQ6r4N19OI6IPh2TrVJmWLlWunf
Cxm6k5LNfYEPHs3Lwvw1mJfNTGYtVGD1K+bBEL9YPG0xNygh9hdVx/6OVLPNUQMA
lskCu3DSgHwJjz8q7uLp1EX6kuev8ndY+sSNjftd4qhak8X7jPjhFhI5BYY2prvr
b8FzY4ne+I9UE64wc6nxOZFK8MqRC0ESLnO0TXPoJXDqKJrKphoZZDE5tWFinIQr
Hvp8F5+bUU9tLqEHvP4dl3VEplUkF9QiQqu13l2nOHd09ZYIJsjEnx4DGD9Pnx8l
4Pobk3thsZTynIb9aq5lK10ZFpQIi2JW5wfHwFvQh8Kb6cd68Vh2L0dft+D8G9gP
oqPWRZCSInIQr0xTMizgcwWPXVCowWnqTDG+hookgr7oVHwp4N98rdFzxnFwDRK6
ppYVDjGzqnGieQDV5idYvs1IJe84/sq6Up/VYvoKV8jS3rm1SCpImQEYh3fLbOHa
BUuO+z9//heUIcw+Jew5Dqlit9ffuIjdTD2ftZS3HtkslkRA9RY7zPQAWjP5Z2aZ
/H+KH6g9nm5wMmt9wekDIL2np6j+MKIx9WkECkepSluLl+ovfuGhE/8CRjw1lzfw
OUDhIbKTI+jkJbaxwfIdqmhQ3qMwQhlFmZy28o6AfIEzBeWDt9nvobVfRRpYXuzJ
TjWzto5R1LFLdo/ywq0F5UenwjmJuG3rYFLFSV2XsZ4dero+1WDGaoPAdapcI0VU
i0t00xW14nFPDgjk7D9lTw5cbNwIBzfdbk8c5IVkPC2skNpKjHC37s84VE347SeI
mC7yoqAeAV1hfhrV3qbXWi8HvVIhNI4LEVs5JBWnSZ4crhV3X8BdKncS6jONblnU
NuSGrKFozsE0YZnGAaVcUySEQm/RMZ17T6UcmYVRAoroxH/U0akJLRsYBZ0kJsQW
f2bgWXy4JxBV7jOmBy+3Xn19rQ5c3+/i89BO1/scGNmHPBE/FvgdH0CRJhRU8Mum
T82t39zM2ICCDVfMdZcWsGKY5U8G/9mrbn6GukdQ2dUQ0Z4cp23AbxBZNY2jcKUQ
U2WXjxJkr3gp3N5NOoGNPjnf+TEeDEmmy5YVbHrwcN11IvuUlHf/ee2g+KUmfkuw
423XrTdhvalZVc6/Y9Q1vOomyfo4vgtQ+dH+/inPYYZGSmuedO2nmMCaw1C/T/R+
1qLEopSF/1ay55X1wEpaP4FUItJprUIZFGp6uqjkZhY5/BMytjD8fu9ZYlUFWVWv
rdjLjfzMI2S30PvUUQGOubXCzvFzDZLx76rqjHGEy9FjU7eH/i9orj6Yt/DTcvX/
I8OXnUiH1uZH95T9tJqgBI+B5BAEeusK0EtvSVQGfkohQonfS4gjGsjNUslZ10Ja
GQyO8VITRjFCy5ceyMGsjelEBIJv3UCYvyYRen4tPf/ZFD5tnhj+v/LLDG7vENXH
jiwynKNTa20cpBHw8otBbDCEte4/1YIwtHTL7fn2gziiA3YBgc/MMULZgLB7jvIp
XSrdk3Io3Anrii0KY0mAeEXzGVKSSmxjpz3EhJtkGzOWT9zWAGKWjnoBSyYA3XJy
wNNgC69d0rUIc/Ww3g07xN4ORl2cZ6iWzjigOzh1NQ4SeljACLbUWvejJMz35X7z
5r6/E7gjL6Fq3umNWssp/jO2nz3ZOofdUFqQx7jzBE2dMqDodfVQYFT7f+mXoqoL
LfidLu7IEA81HTCmAm/KlIkbP5XWvJzCjqXbM6PybKh0kjrbOEq54V0JjcMT4M60
tIz94B9+peP2OWokQsWWuDSm12ytEv6qmmmxSzPcPzdRQVp9DWvIIo9UyWSkmTRr
AjQ+j+D/pQizjdxo7c2PQjdt4vk5o4+3HcV/38EbxdXgEyx0eEORlp8vSU8tb7+/
kWJMOaNzcSjuvEO627kO9bNobQ9OnNQDUcutv4WCTL7nGFMqCa6rhHiVZWwMgfmQ
3cuVeGsahPeehiIGB/lLWb2NEi0bUwAss+qOVJHwxb/SXdgpHsxWBDlE1vgQtP+u
1+nsjkM6Sh91PLonXhnGNp0aVddotUe2YN1T40nagfG8NqUvg+Gi5z33pAREIk0p
jG4FwT8tWIVgbN1Uq+XiEjQRxaa7pJrzd2qFCbtDXuDvplSc2OKgczkQG0GFi/2u
PLJ4BY6QVzthq70WgdL8R+kIrJDVec4icOSry6miAKw2ICxUhHUN+6AmXhQUY2y+
nTKxnLFateXz3coIijem8QZzDXj1DtBAR7MaTfp1TfPtX2o9M8N4oAeCEtw5jwcV
OKgY20EuNS+Q5pl6RxIovdbT2bfg/zsbEaYbRZ/VvQtb10iUqoq2lKh3ONiPOwni
qP7s/c3jhA4FLjlCys3+iRpFS+RPe9fgWqVAXmQIZT+o5gaDyel++1N8N1Sd3WIw
PqMKEnKx2+BXYdnMHJFAfmhUunsMrv7GmzpULXB7AijW8CYiBQgRtrIuuYL6JRKo
XDZOXp7IzH2685v2LBJFqreNeL5TDv0cEHuNtVmgQacndQzZYzeT+vLF7groANku
zSZvW6c8IV8oR6oYIdHYwChLOMF3A2CAMEjnATBe8sumAbbyekEI2jOgxlkhlxQE
qHV1QY3kh8ygwD+Pc0r/g6rpZXzdY1ogFjrbQnQBCpCB0DK4ne7KSpSCBL6AAQtS
36U3lShNRzy6lHfEqxk+nFnA/gtS/MTntsYWFmPMu0t+vXQ/D2nnUWXwLUc4dcbK
F8GO1wIwpGEz65oahEvtngrcd33vaHAZX75VA1Sj0/Yi9wM6+S5JY5bR0XZZgjjH
n+Xmy5btFkD2BiVWmybE5x+7jDNy04GL/kdrNZf/4VNcjcByslQSkudNyCf5zfm8
t+sDovaMov/U1MjRRmYJN5rUuebVnMygZIZif1/NQcZS7ZHygaq4ZwwQGcMJi0nF
IpBewvLpoUMa4rKFWxMEp/Xod7L4JuzluG+VAunCjSO4g2IMc7zKYciJ89dfVxi+
gQWvvLm5WzoM+A/mbIm/ru59AQqifcZ6R92ecLse0BdOz/FsMxfE6akiwRbdrHIA
Lfm5C8tKhtZOz8rjrTnAkWoYzzTdjn9QVMJDlYZENubAie63vJ4Ig0EDO84w8rhf
PU73ZKbJ/zoJNs/u1DUa1LytBmeREuobQCMT3nYUVCk8orNmdO+YFhBxZe3wV1tX
TU6sxnCMO/IFosftbNWRPMmqf0OwdLx2ULYGG8s2z9E5ZzKpaaw/Fr0GsVnqIAh2
CUjhFygtGcYqsIEQodAir7g60/nvTs2W5aI5qV5tOnU+genXtwey15L6ToKHFtZo
VOG+/Wkj1OPXnGm3KYrlBdT5hngWvNsw1YDAQ55V8zhKJtvRO7bCpXHRXHqHDJ5m
GlPon+W4TXzHmq0ipZH+Vf9E6w27nWh8zeujkexNHQMzsBF9uu5BodUmFkhuMqSZ
eSkqlw5JEEXSkIhYM76jvBzWzuK4owOnI2gENixHtP66IzOCEpbyyfgXtxwO6+gY
VdWxgmq6G6nH1VNEVmJ0hegiEyynuyamwoCxgDOPVB8kXs96amEjRRMF/HDFHnih
jsBP6quba3RlKhA5q1Fa8KFTbzIodcvY3TrsXPJSLwuxTxSUGYwtT4ktUNJ9tzwe
BqVaCiUHkQnTRPja4V4DdefSTYMbJa5sMVTy3LAaawUAAJnSuPJCIFo7KG3tGiAj
4hMP4f6As3be87dw6EEnv8TglKoKgjhKLqK5Z9771Bv8huBlnlBuCShmzopk69hu
3G+6+lWYtNhv+oYanh26KRFRsiGFMNlJDN+A7S/4WSK8VyQoLMhq5yZCBL+1d1pM
c9mUyn3MWrM0ufvRwpvvAHTPibt1Iae4LvvzuthMJ17WuHKUR9kPnJx92KIvuh6P
GOJN/0FiUiZf/60+D+asYzfVF0gQPViUKNx0uCXlyu84U98HAw3WIF5MKiVtZr6f
rSTwCyBQjyro7jueWC2fdc92UDa+lLzFvCVNUDriPlLL2QLI02oNjzGD0WBHWQh5
Q1CsGrGFzk12+b71ZRLZt4liMfoBn0WO/ZNXtTUU0r9EU1OE22GuGIpl2aJ7udJg
9MBOlGDqix/rtkhs+l8rdxqM45WTOfmnqWeQ8UwUMI2msz7Bn4M/aHnIEfGfLNf0
6S3ACbhaEknjRRsTEfU3uOnxfMsZUnu5X5zffLY8RU8MY7bASSCN9csORyJxpSDt
k0phbLt+lRB8C6zoAw5U+AL0wOwOIMJDU549wAxRiFk2/lx8GwcM2FIzz+yYXdpi
f3+33WExyiXn1I17PB0JYcBJ2HsaSiXgFnFlp/tmArFZwCrbrp1xB3nOzvFQg/q4
aQQ69RChhjLbIUg8wIBgJuVBUy43tQlcsN8SKbhb4k6YaIN1u3lvd6oFItr1IzfR
FntqHIW4R3cVYTJmPi+F4EkN855SfLW9Uq3UXCtbF4z92goxCXZWUIuic57HAwnw
LNQO/q7hqu/u9vrBmr2A7Lw90zL/Yu+VwttfcwzXbENNaQXm5s1NGcc/WjdqIIP+
VeukA9wqUGiTGShWcj5w+ZtSbyhvOFijjNtddCiMDC5q+LrCrDO/Z0A31l8W7i3v
fPKQZWizbYa3FLq8azz6wpLu4syiyaIm49OclSD069lCoSpw6oKekSZE3SBwxRha
QznAr3GnvtSXPkxCfNJaYkUdpM+9pgm/E0RMzzQdnKGYb+OVosirLERe2b+W2ZkL
Zt92h8nPJWlqsXR63iNvOJyS3qr2hBsM6ZjT2wrc83O2k4uqGnvJ5Gi7jsq3qthZ
7WxdxYasvbYDyKiYzeiF1yHvY8fReqtO/zAqIrFw/x46aNqlTf7XYju1FyEbpZR3
/5k5WgQDyl0C4fNMSYqMjtitvRcdQ81gXvE0nS99G3ecqSbsIHTQniJMjE4JwQN9
prwUteg/7+AM1nKvXzBEotAXpmLnYBbk24srj1jwJqeDmGqFsNI//p7tGJdaRLiJ
a9vcQZP7wuXWJZD436LJEBjWZqlo27vfwf6v5i9ZxjaC4QITzJorlGeurwmhfwDo
uTkc4QyIec5KlOm9HzyFnHZFbGZl5hzq8kDqCT6+szfT9Q2ak8fbEQrnPjTsXhEW
++v6NBO7NTsHs7rXwlC5lijfTqWklfKjywbXaKMpYwZ8Nyzc1fqv8ScVIW1rqznz
XOESVshDfhJFONl7z/r4ghsBgHJwfjGjv4d8e0M2GpjOWQoJAf3nLDh1y8Ui2mwi
eh9SVCNHh9tyYeIhpYYXqZmH9N64y7tZ0w/7WKcJQBsvd2kz+lLkNGlPeUd5Erik
twApHYd8TdJvBtOFlBQx4aLktG5QWXfRDFLVvR/w2OmyYEw/rHk3j+gdFw/49Gsj
hJomrWiX8EVpi0IwByj1saUO3xg+MdkSb3vyt74a3Xj60CXxmKEyL4VqTln/fy3z
HTMT+00o9sXwhtSfq/P3xDXUjj+2QuSPuliOcnu8WBJ5GyVKF0LyW+jpUEZdYHfY
r22hlEnUUabXkDSr7U7he/7GaImVKc3COh682DZCsY4L/ZdAb1gJ5y5/9lDTIXsd
hx250aR2DVpjgWznio/OfVCvrmtDQeDSwkXQBYy/zmkXRHe7TxJz4e3LRgVDTZ+a
7Yk2wsnUmvVCPQ7Cvw2YFZkbi7lshHufRqqZ0dVg6tAITxhGztvSlYuIuHUT9TAI
bcI31Z1nYqiE3FyMQok1dd99ES8M0vme1msyN9P0v4O62FqFpqT6BdrOBY6LKTIu
SEXMbL5jrZ0hIoEaaEdHsB/gu4+bSsSR4I5wt0vRoICz23qEVv2kbELWIvu7sPNo
T/CuZSBo1MFwW/AFuI1dqwTeyXxx/zwgCVfV/YnJiN8VTKSPmhrLlP1wpdAEvIY+
WA5kN2rQtdokI7Tm0Jzug3g1mHVOp9JiQtrcH2uQBqaPZZESXBcwTBBQ+urEcBVX
FJapo3E9tpMm3Dzet01IvE1DBf/WOp+WaYAh84Jdr+anU4erItlPSswU1k9HGVY5
3cBUNt6jEa8nrPOA2+prBCPX7lQeVKYdvyJSm0YALjAZG/awUVWVYnOCCORNqilg
Z4WJ/tx0rCfgmPHpqyR6/luEx3b9ZGePZDOHUlsUVft1CkU+lMzjgIdGeCRwKPeI
kv+PQjVBvqQEshH64VbmiYqyGL16S64mfYKzxSK5512ELb0d8v5BpS1VSFsCznKQ
2wa5WobT7JecJADMkx0QpCnnzoTQPt95FkHxOEIvXFCndWhOVcr7r/2Yb6wm/M7B
foP2Vak2Jb87JSltXxMMHytPP+pd/mxl8IrBrBrcTec+D5xY5fjLFgzu65GcxJnG
50nf41GF5qQtESPIMC2tJs7Rvl2Nm5S6TsFWlaW1TbvZYaZb7WR+/kd+NuExeezf
ziNX5odnbM3CCHvzZNdxQAd8kLnF+jOvxWgg4giNIUotyLnt04yP7TIAyfaf1L7Y
glxzLTJ7L7pN+wdfIY4btq+3kXhUvBxIrzBL233vmL9oT/JO7h5ak6GI6WBUUKMC
vFenYbVni6rBDN9AxGerS0UBQIxp9hQRSNcmVwO6jj7Rjoe4+cv+vhd7zoJkLufP
3VkVbXQw19ScSYQYz5AeCtcecEo8FQqUA3HdQvYxzXUbBXhFK0y2dccX547MV7y7
lnESI6zTyayzeKSpIXPXYPjjK52Kn10z//Dzdk1Vu9j6w3jGYJ9AeXmA9PNTbyWB
Q45Tz7/8+u2WdnYYv9GRsR2uAOb0k5foTEaTo6ZgN3y2is33iDGVjUFJACq95i82
KG02BIbgjuLkRmwTSfHjqp8wub6LrTNKCPNzgUNCdpG2fYxJIw5leS8e6Rs7xlGO
/cLGC8127dT+tmBae4m/VBqcLpUZCirP6MF1utdLdTy6vgl1ESFZoyViIoR2bMMZ
9pqj2EjjMeABPkXD1u/AUHRMvL4XDqFfH6b1Bok11Hwuyrb/q92p5rwaxK/ZWEIV
4wfRqjS6+v8yUiJUYLMBifoN44xKS+HAnE/JzNn1crrUZle4EFoI4wfByPaKfJnu
Mu00SxApVsEa1hnGF+0KVlFlibm8PeKzy/J9+e7FPXRNwrmFjLRUM/qblMBQOLVW
tUAKNZ/tCbqTY5J9kXpxNBtEVZXOAqrmZLMwz6XK1EcOOIt+Z9h7D3Hco/DawCAe
Xh1S4J3Rk4J6o3tbSAoNArKcjcCyTB40goEQmc19tHOiRJF9Kba18GsfbAchbhOp
brUFIkAEdIuQsksnHcpxQORJll156av5ymGl6mKN1aMojgZ/7kPFI0PeihMoJx0x
5wiTbHULzm7OVUNPdP3KqkQsN/JGLrrqo97eS7YLG6GQy3g24O4t45nWM6ir7AuL
DIeEL2OT6yBZgAOKr15n+JmYCZEl2ivwrgrNZqKufbi9QY5gVauKgqn2YJpeC3CZ
JMpxEArvr28oNVWuPK4eQYe4rB4TgdNiODDF5OqIvWceXvCgALHUODhTx/0EDp2C
z8IMhn30/7MnX3OaucNBoWh0goZZ+gb4F0UmNUx99w/NBMtcmi5Wht7Qd3n1Qy86
LfvHYFOEsX+gP69UDIqvD12T35mNevsHyLhvV2Ccqvzkaf50rqyd3clI5MfvHGBm
Bb3edqTKkBS2dyyhYd/YKvEgKMDbvFjUmKA+OoYFPokIVqQKRiN5XpYF4B/l/MWn
TuXphymFMx2rrWDsiPX5wqPTxou8kX1ZZ4pWWdgkOXM9UIEEeDjls3q7w/qMsMQD
Ns66F/dDVjy41/etxMivhiRsOupg95hTpMhW8tXfM0giuPeKJ2q534twFnhY90LX
KjzM3pwCryYEUJB3Xh80cAwbBj1hDRrqJKPdMcuFvW+3kZeBJD2HL3G3cEnSMhWe
ylXMOgKUdbGivQmlFq4TV2IfzsYVt8KVrYgoMqtkFGBiixEKfOcLsdxdq+xUazeV
PhKKwnQFS9fFbxXEXot2/PtFku84tsxliRQecP0W8pyFuuUjbb/9URHWFLjIbYKG
dDm4tC5P1JxwulH72xDtpM543F/91bgDCgDTkVo2Z6dwMrxzrCpTrVnUkLQSFxqq
ABR/rOds9H+uEJKOGSUn3taLIOiWw5jzZteN+FzovDlt58exxIoHwewBYuRs2k44
8BlEzx88ctK4toxssAfGlOIKC6akbaTYpb2L1UbPlm7AEX4+Sn+6fOICu6Db8qfT
VeqrXy/tbF4EqkyvrAGtrBOQVmrGeMBpdUY74y0lBA71/0wP8gptxs5gpRuLaqHU
VO2oha1Uj7OYpPEroshm2DP5ewHEPZWzuIiz737oMhtmFbgx2piqopwe8t/jisnG
5ZmoVG97rfiVf+QRcYmy4559wfpOzvHUTepb3e+1LV4ehFHhmJFUpntYpUJmSZHa
Si30K8zbbD0sTS2zF35sRtIbV3Xep2UD5a/Ve1l4TM+/YGFCiv73S+cxKif2Ui3z
UFEFdrCt4i3xUGdjYMjrr0o5Ic2h+bvSLo9A29aNu5zrNIzSG0/hbBeS4ybvZ2M6
z8CYKzLTCmIR70s8e/Cqsw16NHHaVIDHIXOmYOYxaDb2Xbo2YNIsE7dC2mWU6fc9
PKoYV6mhptq110h4Yb4V01lNTbMFn7TrpUMj+6ALS2SYn0rW4b7LDmWXc+wzeQL0
BgKwLULd9MO6EvMkgpIXLdFUOUSJ2i7YtV0avrOp8otQAsYmr4veBJe1sUDk8u9C
AujlEazV9eCLD/iwAKHBRO5M/ApCunkU5ZayVZEt0qb2m3/ZiX9h0lgPcxFwsRHr
G+R/nlSf8qpFwAuQDI8jp8i+MznDXursQJLjHemq4NDLeI4JRv4g/4jbXs0FINMU
czVa8g4EfdF4PMN05Sb3JndgoKHI5Voubb0o/ZGbxPcmwbcdwUYERASE0/ydop+R
cBTNoGhPH4abe0RTsgq+mnHc5ev4eF3oLQ9wLWc5YyjppNbFLXoNXEpNW7Vg/ui+
ckXMOf/ZxE9ZQ7aEo/e10fZx7LgNih579Ni60LHUikNf8pZUN5SwpfGYtSrFdnN7
RMkhEK0hjMMY08rILF5AT8ccem1q5E7ez8z/2kjA2C4Llc4LPrfHhBya7xW6TfJm
lMjWOsUJ//l9R6CrQBR2NCiCH9oabagtX9AlqWhsB/UWRdNcdwGSHYJe8hb1LLJe
JGwhIX15wNMdFoAI5zbFimIyEn0kghVgIhWtRSwQUDkb9Cax0Q7Hawb75xNZvsDF
BAJ3p/0+bMqIl51vtq2qinWKx8C6/Yugy31nvjIN1OPZaOWFoFBeX/MggPCLZ37k
`protect END_PROTECTED
