`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0c72E4FWQDBWMct6OQvKJ0LAJ719fnOZ4oQLv1yvvh49DxsF/WoBN7YQanQLNbW7
n7V+0lcSk13siPrCbxcud52R6DPiUBnOM5XpOx6hHgEsbX5+4nDFE4+czwXL9eND
YMVANwYeARk5ThITzjfTxKWGewyU64VKj8sWS26df5uDliNZX3/pIYWa7Ug3/8QX
+cs3kCVALAqrjZlZrDzEBsV1TilLO9Rqqnwo1ko0ha8tNN/Hr7AFp+Re+j+PbS04
dOIryGoEii5ThVTFRZFcNLoOStO5BuxYVce4S0zVa8ufAzxX+Lq5p1pcQw06gvgT
DnGonbNaHz7vkNrcfOXv8G3TxsojbUgyTu7SWZ1sHS9EzQs17VV8FGZmBI2tJ/Bj
3lgIfoGEkAZuBk60qze0Rh6qFA8XzSR9RwM1lSfB/2vxPByrBcb+V2K/snaZjd8+
Jy82lLpRJBk6LPfLIZI9ZTwiiInK2zMIy6sdf7DSMGQkudDIXJgvOMoD/jte5mhx
ETOUp1l8pt0NAIjj377ZqILQm+F/rOF+qwuhluaIWhEoWz+qxMv9vhIndcqY3zFU
B85dLxiRVanKsUjWJBeOsRxL7DMmuArhbOFG80UvIamIttzu4fdd8O16HX7pI+oy
kkSrY4p8ZrX2c19ZKpnLFd588v73OczF76VBy2DpUDd3zvNg/3+K/r3FfzWYYKu5
xPoPiFhyMhLc9ilif3DP3JCseJCdS9pSyp4re6DK1DFax5LDOBkKZWqW87mCYXRB
XqtZ7fOlxu4PP8HOlr6+3AA0l5CVD9HFbYOznSl7oSg5zUIgEesjPS+YTSqPujS0
GCXfES9G6DTK7X0wkjFs7rB4gcWsj6oObaQ014pPslgY93Gwh7RxwxXJuurl3z7+
OI5Dd0vrVBDYoPKu/fO+lyXKt+8a5Hc2Ka//8k+0+y4oU9GBhjgW2Z3Yr+WA1dO+
Y6N6q2vzqmZ4O6CK+djeFz8xy3UZSpCJsG4fiB9B8L8UT+ZWPuSorHVtge/ACJ4T
ROKL/uzRJsDsDK7JKnfI9TVTwG9AyYCYEY5KKWZvAqnB9zqdT/fKrsXAVzFO75GM
R/M3/8/xPWEikqeeKknYHVRRRnderPZPOtE5GnXDF4Qspdey/QyG/cPmGTQEazz9
vaobJz2HQHNKFVCZkVO6zTkeQryQOelxHvS1Mncug1ay8AF8syVXFb8UtOtKaKEn
5KApNu0b58B3DW8rbto+NMm6gxZ5nRs0RDhBdGSQnbngh9GUKkS/9bQ5pXuj3X97
LVOixfyEHraphUUfC2/3Y0NWmaIjXMisCrcYzICmdkuxI44gdZ46m8MLTVD6E80O
4uaRxOwHH1PaRXc3i1prrrdTlrI7Ym7z8dERbVCUa9t9aFU7IYiJ/zcbGQuNfpu9
0aL2SZV0c3ni3fu/Bf7iRr7imof1UQDA10+GwXCwm1TOlLGCW+seMdRflxJEx0qN
RgkJSPMepR1870scmJSs/xr6utU/JLXeBXuRGwb6EaDofoA+I3DKBEWrydE/nskv
a4E78S56OT86/qH8KV4Z79gtFtkCRUstkl6v94hExDN5FwOQE0YpZpHY/VeqAvn7
8XyFGSNbB4IKaePs3rjSkccCrSbslqlYtOv70HRAuq9xktEauzmequnjc79gAOSW
r9C/MyFVgzOYCZmyve5fp49o5GjYbY6QOisIyehtqNBx2X+wPgFcRwputqk8YcWz
EI+Eh+vNRzUYyiQKZCPqFbcoeMjP9QorIWtUdUFnGA039w0OXzMB0D6PZDJWas0C
eHEf9zFWi5QTVWqveCP3MbZApfd4j17usAAlPYvocpy5lCUSBmuUO07uz05oLWtb
QMoEHvtaSwNm6fW/nmc2MA==
`protect END_PROTECTED
