`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
unsE4yPxd8dR4sY1H3afD+958/tSEZsAL4309t/Os6LQeRxuEV7ZEf0ifG25uDtE
ust5aZeb6sBIijui8DDDE2p0uL8FjAQZrdOn0aEop3UD992C7JfpJ4B/ZaV+Sl/4
XkM6B9RIuj+WRcsxvwbVtDAjSajhkwzYXEgEjNEBjpjeM/IkUORfdalkgsmhLN9z
sHls0ZgHJa1sA2T61IF3zWqhbhfuq+Kx8ZyYhczo99S/5YTydduqi618rh7UuhN+
8diupPeMsBc3vbyi5hKlA1ifrITJe70DMv6zwU6W7Qra7G0twCTZCFMePuH3WcK2
cJzrlYIOHQd7JrpHbh2cFaGh57o9xqG0bV+15pV6xVz6DCt0qMmxO9P6SLHpSipI
RXW/ys+Lk5gxAraXOF5bzKrQIeDVrPJQS9xeX1Wg7M58VFIH7xr7lBYnI6TWsqVe
pnvkEdnmCKPJyHnP0UBm7831tg+IMOeRFyJTNviphfsHQAeAqYSrVXxS7X/zZOY+
BJ3KRiwnU3yHzFarPrH59dVUJzSlpyHb9niVD6MdwU0Ht2S0GOrOHYTK1TbgEU30
BPmZsVINF9Yk7dbdAtGYgbgmd5Ddnnq9YaoI3DKcwOFaKOLTGn/hoFUN5XVW28ep
71I9mNReNKvoft/iJBTbhHlecLbOqdQxjblq6Lr/2SofshRhCvWQtlvB8v4tNwM6
wMJURPGhc2Xd8rqtPzmmnr3ETxbP/jRs1E/wrKKCqFvLfItjxBQB4qnHLuyfOt+y
WFhRHgmAy2yuk4dAZkhV7uItYxniRrAxA6WJhvQTdRPzsFkqew4uzcD8q1zdDiV5
YOwq7BOyna3LyhJ/Y6SpkQRvXeidCs434iPpGOkEIt6wFOwCK4/HoDbFiCHtGw8n
K6EHt/poZSC2fKkQcVQ7wLrva3cXfAJcODoryAOq8aTY8IZcBH2V2B06//YySDD8
CmKQ81KR5Vadn3VuWUIBMyRUw06N23waVTiMYx77pRCF2puk3dgcl1mfTefpg05e
XyW/UTw6ZFywnvSAfmNtfAHA0BVzmO4veYUYYuemK4NPNBV+52jwP62nKNKLmJYL
ORd6xrDhBgEnnyvN/8BKJCdyWRw7T44H2OH60A746kxDMk8AKe02f5SLXcwS5cch
vTfqJrvVZ9oU0JLxIPknrH6gG29SP9FS/grNGrNDIIUSYI5fmeUjwsLDsAYVWwIl
E3q65nivDzBWZJsdXhTM9Y1j0vZP+ZxNB5r4ZCLkNsB8c1lMQugeQnbR1SgOp+/+
ZGAI2aD+kdP5CL8isMTA3K52p5Is7xgtrp4Kywj492Y63aYnAY1fD6rApmktjgPq
vO2ubMz+G1KKFPiDet5IuWzKX/PB+LnTzihevsa8HEM6OAXIPtCq9sDI+ygBMW/h
lSP7KjcdxWumDFeichfwosBz2uSIkqtichRiHoBpIVsrI+l+i3USAWeDIqIPg6Tb
Rd9oXWWb7ybylKpRNMuk6IALNagK4d8hAPR3pLMnloNGL3/Hc9C2xggLLbgOkiaX
Wgp88XXmAb/847t2zhHgPbqCgi9Mt//4xMewAfHHzeWAX/oQbSevFNNSMzK7soRX
LSfvyEZZ9ehIeoP4ZfXjWMXLR0+VpECJ2Ee0/QUtPImtV6xYbu7/P6Yi08QBVB70
f+jna4Pu2Pg0sHj2iOKsiai+abkeMF1SC6Yhnr3ClG4pzaer+7UYBvl1IJrmbz8D
FS9FkidBmDtcvhkJFkNxzZF/0iwPGmNhjH/LBFAxCEvg9yBmEIsNFvQmCyX/j81m
UtqQewgAVGrNxgm52EiGWsq9W8LMBjeD9Z0lYiO76wzRxuhcNnH/gkaV0kVWZgt9
MXya5GgnrLyobEZimq0W81/OxPlfFsEzk8xnJQmPjNZf6Mhdz+p/eMOMVzRYO8TJ
uMhv/MpHDgwJjkQWJoEIbT4Rbj2nsSS6My5TssSVgGU81AXnKzwNqbim5asU0Enw
lZwY4rIu9NOjliUJS77AZBmlDYg9O7RdQRCP8jQLS8D4O8kTSAuPx30CfD121ZsO
1LWMBxqgyMqIBdQMNltLeK+mQASfhv22S/z8aeUS6cLF1ruvGHirS3V6BMXrUoax
iDxBwliyTEO/0mVmRskj41Y1LhON7zU9lugPFDNfIE0D3NFEH9UxbkjNE95nAzXA
A3a6OF055ju4lT3IXOkq90naW6PxD2sug3q7trXJ7RFCjSqex4r8lII0BqSSUrad
uUGdccHRjgnKQqyMlJuH9Wea4keRbhwWD2P7MQZ01Y3zB1B1qZ3k13sfjYKHdJNh
2tY1NcqJHYl36y5ugkNUT8av0EwVbRDRTMh+Gv9BdEJQG4NcRZRuQaNKNBZgsHBt
bKPxD6VTp6S5au56Rc0zeZSC2xFqfrmPWY1phPU0H0mZMX2/RX4XBVJsGjYGcyHc
3hNO7KeJo5rXn+QtQp4gQgpO47pd4e/uDQYZOt/6/uUwdZzAVHeCgYZq7nQbNnEH
6uu4p3w2p1ihUL/x+dbhwgwfEfptqgfQXpuxGMKq9DKVLfNX161PBOOk0MRPRI8K
/OIcJ3wbavhRsH+uGXPLDLxoLi1p6uTo35M73LG4lG3J/hlXBjUnw7J9bU50BqwO
q3ex8GBEhuVOaybjh5JbxLWXGNDeAP9qN4oUcVrkISBAmss/8j7NQZTcnTXPWOVV
+HbExztNONskI3g8RTv77avhEI/uWdOqVUbBVr9iRxt2xOTPNPSaMRFhYMzML7Bb
A91m698ctC5xEPzVWIEgsxqOMNsPDchMVulPg42cmS8RofzQSSPxWkQnAW2UNlTS
Wip5oCTZI7YQrUcYR9WGj/rNPeYLzYNlxU8s03AyXl5CC5g+BAv+2624xfyxtr+J
ml9CegTNAlMz7JsYjknU5guwGKasfTCFpwL9KGZTBb/8r00SfbrB4Bnvb8WWNDdl
0wquA0dpwR+krnDy/7n7Brlvkt0SavhrdEeHkdWHw0KPlDJi8OyqAhQIE/cj3ZOF
9Ya4uIGya/iY32YU8+AnKZJ1y1oiIarQoRYOnlsuMgeVHBRVBZLYUdTDBn2IOcLn
p0+nETJVsqOt+YGkPbKNrUk+pbJjrDSgVcjvd08KF2DCQ7fcl/HERon/2Awoh+yW
LGZ8ha4ys2H+s3e6cW7LRY4KyF32UrIXCGqySM7Rxjh+BowgM6k4u44v4O9LBOfR
n+SkaGaadyPI8ei2KBOPIs0i7dMrfSbTWxdH5eFzT0T7z7kmcxn3q1Eh3FyKrVFg
bWd0iukgEmU3Ok9o7sTZuNC5oP6551nTz8QpHSCAYCqqlel3y8uBBGBKd71esa5M
fUxld2P2of9jchKu8U3GASef95zGRnB/NclCSn+ZEDGu+mAjVa8VJK4CyQMfleSD
LRgdMlPlBvA3ZQ5vGat7XZOa2Fhf+HgQooR6ZR5MYCdXk+p8QZYyBbpMUx7DHYns
wHA7gmW4n8ODBTk8CGmulLbRlobXByhFgncpMZQObtqDBk+t/+To12F2XGzM4aMJ
ClCflGniGB618fRm5ViKmgrch8sQuqH2tegmaZKbfbEzswpVW39w7uHxvGWw7S33
uCGvxpisbdSRavUj2MbPM9PaDHROPwKwneR87LS6pTpg+52Jn5r0m6M9VBfw8PLi
JaSQUDvG6y+3mP8OHrkp2dRocQX7ZLDStpbTyhRAqD1zMP1QTt3AOwftySV7tz/K
u5Cyq3Ojh2Q7V+qVQdFKvNTvupCRAiWlovutSHyzHBFSMWMA7g4IDAXXOhbWFtz/
Yu9JsKynYf/NvkzuDsbofC7l1Lw0/ZLkORk1VgmGe4AY6pvKnxU/EqvL7/fM7+MA
DoHIh3+8/RXt1AmpIXmuDcTSI8kwhTQSNwNW0vGEnqws6Gplw+tJhlOebLSeHDbW
o1bhgD3YIatpVCbXk3qn9sm/3rohu8uc9lRJ7AkZwnR1T+sQPyam37SHRnuO7fWr
ZbnlHxCf2K97GrYoF0kOerlko6SNXlKOe9s502FYpFDVDQE//O7gMdGufdNlXzxV
t6ASolU6Yx+EwWVEk6y6/YBhf+AFQL0cTVhUwPfowcOHYN+BufLbEyhSgnREhGRO
FR+sZhDbDpcJVE+NcosgpP6ho0FPv20x3hND4auug9X2ymFOrLxXDlqI7mebAPMV
Q99ycSPKcF73f5wbIJCZ0e1AS0l5AxSI6itfqssRsDimJGYqYAw3Mt87Gsk7d6Fr
8X8Vp/wvMvf7RHZD13cQxPMZklzIZhEWif5fi/uuOS8SlJkoKBTORBIU8sSVtEnJ
zzmFKrTVN3vdXqaM31NR3wkjqjasVvRAKmb1w8ANrvfyZv1C+xsWhzbzhCxgNdHR
djtsA+8RYztuucKRYk9d53bCRAKk3ZGw4n/RwLWwdU72GChnfRJsvdM4S/NuKuEe
sTZrmH35HUhwfA+ceaVeu3VYUDntTn/x7MuTU1ggBqrw551FOQ9iZsqWFWMGp8/j
XFvIjaZUtcjYOzLC/qSIUbakjjEyE6rRJ/ieC7i6UdEHsqmj/i0vFwj89LGlyexW
GJ2PDAuOf0C+hDjXOFtvZYCTCdJP9lhihbvsQihTDc8loDl7K7OXp9tWcvZvvEDN
ezMhkBNzn5pBX3sgMc3vh1mcT39RDw6RVeg9EvKwyNLOJbBBJbbs7kpjjF2NK9e0
Yge9ffbfAWf3gDmQ2HIi3928Z3pNz+yu+cyXpR2XPhLzerVFuSMLN1rEhKt+vJHy
4cCToklzzZwlGNvEh7ln3hG0FuN+PZ+NYAZeB1iT9zZ9qLcHIL8H9hmYcBNsjHQE
x6ZQf0hlrDpYL5hcjnxDp/YDNVYAtHWcrVpLG4bxrXrE2YpF7N3KSLXLGtybRaEo
PlA5cNSjRn9BNyagMhSGUSrz2aRZOH3Hc1RP3yFMESQDEVlWSDa9PiL1HkXVUubS
SecgI/bduJfOZxlm/2hBcw1WwDJ5xYo6pc4OPCsyme5CmoBvfDKVW7ri0vgV33DW
aS+r9ybyRCVAYiuNenX9QM2Mk5L2zCCBVwg6JHNVwZ4ZURZpXFU6ygXU1w8GxCbD
cRWTVBqhqT75NGO5vSr8BP7WrZc3du5dmQOAuNICs5xLRgEA2D1k1boAyXrL0CP0
aRU5gNKkwTBqV9GZcriNwf4BZ0ic/2QRW0rAtAHW+Tpuov5mDA8T51kodM4mB18U
VCNmOGLAudSRI5W3uj0niZb213rFVxbYp7dDzdr3qsDEerUmQX7Er6bTSqL8zOk3
KcTjyOFaGMGIpd3k1dV96owASAfb1uKjkafgi5t02AwkbpGsQe5ctyhPgOHeQc+f
Wca/IUJpzRGvQWpoxRpv1VHlLR7ge7cww5HFmQCgn1v01kcO2hWChYri8i844sNm
BtfnLLZ5kQcMkDuxbXvCAnJKSKsWxFKZOIg9glcBI3s=
`protect END_PROTECTED
