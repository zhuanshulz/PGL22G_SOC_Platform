`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cBcut+N8Sd6Kbuo8sGfeW7mJVDEp8BA7BhXvPI3mV8+0QKsB0B4poA+t6ZU9cYi8
huWCTJINMER/c6sTrz3XbNYksjfuPic81dFoojw8finPbPY/mTooqge7JWPrt90x
lac2gpF5L7If2Go1b4Vqnb8R6p2OArVquvTe0rgxWgf6ctp2G9Or1r64LjTGx2Mm
CORrpn3aWcAqHbxp2tbTOw7rFlic4q4zZ4wQObHVfVe4NURnLO/yhvg37vOgmTVR
3QmT9hLD9pOrxsoRZnmW7X91WKxb8sMW1zhRahAPUj6p1ySjQ7LA4de7wt4qkHBa
avREqCt56slQQCv1hti/XCQq5ZMApYLC/QTEOXkyWafVfok3qeZB5seZCO2C2iUb
a+swxXM3nn8ZluRjyBFFUuTKAbqsgb1vDgFiCT3GW71fv64yAIff//bBbyQJtraQ
3bX3928ef8F0Ft9jvrgHip7lv+UNs8o+am8akPEcBQj/udZ9CnbSHxzgM3yrTv9A
7VulSA+hvI0teYWtcV/W9NzU5bgKTxoIkKJINSPqVjAwcfK0qhRrbj1O6Ny8OMEE
6s+Cs2upFbngCuwmZRhWpEI9A0XX7L+iKemPiTXgjXByfSSO6KOQnL/dCaLz5pgK
OnSWVp4V0ErZkPf5SXv8HPqPIFHLjgf0RmF4mMWOwbm/1M/3CF7Guisr+ix2TlTk
GV1Ydt9eKz7ClxDpUk/wOh/ivvEWRRAHGiJBZXFiHkFS3FjlpSkKXrCf8L9F6Zjt
NhB+KRt6R+stsmPmo3cZ1kMSfwU8iCUvOH1U63DkjFoGOOvseTOCYn69t/HRtSLl
lmI3zhhR4f7+4TrEs35LRxiBGPbZl/92M8rEJ99k9v24GlbbB9x+P+VZwz5wpGn6
rRFhFi43jGysdBckQhueA977l9hyLNBOxa++NADaceE8jWxbnXGKKnYZodKC6Q+2
Tugk6ZJVRfhHYGKzt4ieD3Uh86C67WDAti93VQnjsrs+N8LC5MCZR6UkRLi2B1Zt
LZfBc3SJd84CBOlNOnpBjXG7Rk2jH/QA1OulJcbMPx2PeoqxIoJpEONCLYY+TOyP
Elof5AsElAnnHbwqqw8qBKLmwrx4PQMiXB/M5qD//7NyQ8BXoPv5k+agfNP+yYN2
masLwuDeGxquSPsNE/8AOdWWQoROurYtnCS4EtgLHe3vFP14abKs4GWdI/u8f0Mw
QxEKBJo96RmuZMgTVwbOa46YPfWKsxwlndEuJy1uy4PJiVE0I3AAro3+cFizbH76
38nyz9XzaPc+9+/DWHCTcUZ4q1fZX57HmpZsmZFoHuSeDmy7iTct9xZclplkyMU9
+2iV9aq3KEL+PtZCY0N6OQ8GZtpRO+Fy1iq/Ylcjkyr02dcm2NwKVcv8Gq1ExSBQ
IEnO9i3Sy27L2neFjQytdXdH+RjOkZHWKO21cdYjJX78z0bKPvlMMywJ/bKcHGh2
26nh2jp2wRKeO2nAzXJ1bBe5Ew6WgrtiGi0OFF+D/24=
`protect END_PROTECTED
