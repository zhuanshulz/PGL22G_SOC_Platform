`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8lHqZUB2J6ZokmGc+oiON1gl3cyOOZfRPL5s2JBAkUrOn5SVvexwnS2+HwrVGpSG
kZlgD00f3l6nZ5zIKEX0ikA018tmdxlmC3pf6xwnv88TdrVZcoaIbjQF2F6JKxQ1
yfQ6v4zIynRYeNy6c5NBPKQ2vf9TDNtfIFkVEcC1mC06VleDuA+d3K2W76rkhSKd
gFan3glovisGLyBKWaUTboycXnq/F/sEJE/gGUSdwi4t4xyYfXtF6FUx90XZ/e4P
eJz66DZJ1o08BYCH+xSba3revOPY7GSSHx4OsXr0kO4b66WQQcRWLDONXqCGdAGe
1RUXUNtZWiz2JyaiqfwhHNla0EaYB8Ds6lnJ09J8wP/W07qx8dePy2kkHfN/HL9z
JvX24NDiWaQKtKFbG/Fxl0sUs9kurbfWwW4dIcuT4vGTp7RLu/qg+BD+1uqJdwgF
`protect END_PROTECTED
