`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9hDBz3UWttm+wy59Yjc1I5xcm72OXwoiFD01Nn0ACMQrdVqudpufoVWekUMFF8CG
qIhnk3vG9nWDqErgTwvaWxya82JJFDJ+R0gcWoMnOeKueB69+hTWi8z/ASwUK0zC
WlScr0cdfTB0YY965if/WpAkrhKPmTkEqEw3HJL7jljiV1jRzUzqr8VLQwfQwWrN
FphxFO+MPbhxlSGJWIihTw/Y5NIuCKsb7rFkgRqaGZV3FoAddyo0o6EXpFY/M3LT
5SrIgJ2Co9Xu9ZbOS9OvkMxos1V1RTTD3kxz4vQghMtCNZl2B4Kp0uQ2van2Rq9z
SwAHXEQqOihTs+2u6AXg7FYWShpgtJA7MzBe/4OyQF17Ummna/PNN0wsmQAk+c/9
nhLNGmsJMAFBnSfegRNWE15BMIuWIZHeljOb797jCAaX2wsZ91I9jSXKkmKb3Bcq
`protect END_PROTECTED
