`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EZ+sxFfwVusRmcXUyxjIxJ9zEK7kaYhhSyAZBWhd+K5y+O46QBpi+4lGUNjBxs7f
5vEYbzVjHMGUSsOMNrHtCeWD1+tRfkOWWFBmVSj/WmuZ3iZ8AYVdBH40TVWLzwxJ
whjZZeEnMJJtSJjWM9ofHpOBVP89CmAvcQ18QLffvvIIaYv/KA6c7kp3UP84vDtu
1DUJK4MDHfCShM8GMo+I3zp8YlOgwvq+jwrmvu6mk9oIdYoT3S7yrU8U37vi/5+I
2EOvomiEdTg8leCp3XjyvgiSC025JewycBZp5TSuspeipWc/zdzQIj7qFFB1HGoL
H6Zo5RhCHTirDpE9ylUrkcB/h8L0rd4zcAIMo3pciovW4/ZewgklUJlCBu6f8X09
ueyU7AelrtmA9rAO8A6lFVz6Q/CLFkNXSMDK5cFbP9hhF5RHJn77tE/UN2bunQ+N
itCzXiobxx3wilcZaaagEr7WIzmOiytrm0GO8dRM3hi3qRbMY2nABBz8oYGZTqFm
gHxd15XgjJNNa/40r/OOWuFMMj9bk+8RY77/axD01FCjTiUOZmLCnpQlTlzRsiQ8
yf/6gVfysW8JTrd+OEJpFcyMWlkzUjCElm/1cgLhIDqXjIolBlk5URE+RGGJd7+K
vxXm5sRGIut9KxKtCxXjwA==
`protect END_PROTECTED
