`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oXHqRD67kQZBu2/yX3yNenTFO7PnuAQnHdzRaUKwag0SCwVlJmYhyWEQfNcAV+pO
w+z2XI0eWuM22XCNdP8ghScRzr5sw8ejDRZSR+ZJoRH6t3PKQpZJY6dm9uVSeq2T
/UbLCOqb1qWd9c8xOh0mQm+aHhTjYjHNUXvtzMfC/ME1+71wf0O0pbuoEaEqI6C1
saRswW6XafOMBFVtD528VG1BpYCR8No7TrGQ7EeADfiExMF8zFscC6eucJb9b/uy
KfioSNjSKy9SDJEMGxR3X2uvF8HYy6a1ihBvs8t/+/dObEnTkjcBhtuFrTaERKd2
8OJ8szJzksuMQl5jF/USBOwf8oGIze16Cgx8ivXY7150+EjPeITHRka+Q9ZjiXUI
YiOUY56YwdhF2aks0zY9oBEHAAjxpzXtdYNguQdRehJ/gs4dsX0fFIHAAqBZjiZ5
53JZMAHqrhM/KDCTXj3kptVOASdMqk1uw5sTfB22oRCf4Zd8K17nn9OzUUPL9yyk
+CV8J2+rB53gQ5X6hIVzIbNnVE+BHfbLYrBp0kr3sIej7QBUKJPDZoS5QEXGRKv3
bBHMT5CxQPExaMD6fLfhecQtLneiJbeRh1lb8qmj6IwaIMHBkpj8HtDsup+f/KUp
cSTM4X1RK97bkk+uD3LeQb/SNU5jECxoX3g7AveHfW+yXipYsWBPE1c4Q8zP457/
BNUQUFWdFQljAFU64UH7Ath7FqvOmaI/TiBgU8jiJbXQINXMOPutOQr0HnFBYFvo
EQm552G+9hASl+pmQgqb31jnEYmodP/oLn3rpcJraFh33Sw11v2EmABSGLROAt6B
lTGKELx1tKA9nQM6Kj5TNbcpv+LPxzzj+hCV8Cls2PxL1AUl3cT3+1DzJ+N9Cg6x
O0MZIS9MxQM8IlbuFuGAdGLW8ojeqor8/cmxtVo14Cx0bki5SDYq14kZPO9rOoVQ
8ziEket5tOSkRg+Sji4mRs/a8LU0TlGBLEUVlc7CYroiH74kUv7r3Yrup00QBXoP
hzlhjYvB91lid2GTrjhz7e0eGNOXkoDHbXhy/38r7uWI2ivlNEor8QbNr9hNVTtH
ZYHVW44fm9UNf1hQSZhCHrwREtVj4Ks/q9dOxwi3wDaVr0cLEeMyt0rzJXg7tPN6
Rd6JhE0jPtvjtPQ5L6b28xtn+4BQttdwxeCirKxnFFpoVrLKwOf0U5iCIqdljyds
TAcBfp27M2K320wF/Cz3VA8BiJ+3aSj0WWzmz75rEPllyXdpTekRVU43/oNjUnlZ
uE6jRkPi4PB9h029/IP1GOitNduo63REZRpHqNI4VksJ5PT5JS6SYMCa7JL6fEHN
b3GzvfQLCXGFKLE0FTMLShFZX3QrGC7OFLM+f9Tn1KL8NB3lt88SSOymHfQL9nfw
MbGbzy26RVIyepTW2WomeDsAWhVTF/9VCuFUrIjXEKGrk1bLzsn+Lp+VpVglaETg
X90K36l2m73cHsOsMtBnwM7iBznS2afnMYmRFUsk9VzqPyO3jVJ9yXW/Hg1gsvrz
vaBQuUARJjd7dcTowNOflBuWzFScOGBnVjxzB3pnlJIq9AMJnLULL6faTKGpOoj8
vYpFcaZNGhEJN5A1HUguw/r7TKCTmkJn54Ke5cxiwnbPiuLdQZPhcPHyPGZBaG2y
anyeWVKvuIfFV26aocezDdtsRYxZ9x7Od+H2SXaqE4kMQ3z5uoBnajZonus4KJWr
TyjH/boCTEPh8QISjXF2iqL5Aur75E/4N1gBIwxs8KqKCuEAPRmVeL5Q6dYn4KHu
Tw1XTMNlgJEf/wrkgtOT1W8Si7io330NDaFiIZVO35Md9+c/57ICeP8oIVdZ/LPX
ZUmq75Rb8Zr8hAy4XvAwGdmx89Mdy8Tmizcbp1jmHREzyuYl9RmswqHi09KguA99
wiF99+IV6aTf1UIuxtzLt2aySXZbqWQaT7YhsP6YeKNQndHtzQIY2icBE28i9lOa
29iavEJzYaX5lOXrg8BYuNPDW2CAsiYKnaPKt8SutRZPL2wJblTT7aWZM/HepsJ3
lSOAwxY8zZXD/kOmkQEBVbJptQRplXUWCLo/oct1oJHpCZjMVorbOzlVfbHvty6O
ghI96CFqp+L2XLgyLprzl/8ya8+Clg0/uPFWDJ6ESVqkws+qcVZ4RlZPEl7RJ87Y
8bP+YP7fYKVatqydLFpTwWOjzFJuR+Io4LcF1AJH4bzpfqAXdgXWM9jpbLuHTtXE
kkMWK/JSTnvbeZLiHU0xKWXrXt6N/OwvoVg7QLCKzH65BPS8DIPKW/9zMCPy1uG3
rHSnXn1SQ1rJtrG8WHGAmzNLLjZgfunOujj+5vJoD7exYNtL5BA+pA7TQwwhhABY
s/CESuTMgrAEQJhsUCXCMY5IV/8IF+jJx/RPI5/Bh3iR14wEmBECXJYsSDx6f1Hp
Jg38zqrYbsEwBKfFU9zVLjzhQ6BbUlB9dDf5H+ALu/32f06hddD2urQEGs9qXEBS
bDeaxWTMYrbN4txU2yCukDgJnkQw2+mOsV8nqh/3WYC08lv3545QJYse3DI1kv++
YA5Ve2eAeC/P2TNaAmmFZrXr4rx87eXrW/LdTr3dxSnPN3B5Lw+N92tpYMn9U/md
awOirnX1helaq8EgsMg995DOSqL0VjE5pAXrmm5jW+wmWyGy236mK3xQdF69c+Wp
PQeD1KI8bI7z09Jb532RiEHPmZg5QFatEAnDc/gXN270g5NX21EnVO7diXVXMUsI
N54QvGzeGS2rtvtpPiD64mvbjyNIjMlzN1AdOGZnwb6EPVyBWcs3hJTLH0FN8/QB
rjJN1djSZRgt+EMenOR/ZgibWjSt/p/W41Y1bpiDk9rHgvOBU6A/vE68MQ0bYLr6
FreYjuP8mFhNFonxJAkMEUt7rS9o8t7SRZV6jepixHQjaG+XqW+Ud+VP/F++3IxP
jCkHGFVeFxW7wGKa5gUNKKKG0N4eCO0mFDGWixAyYZRnbsN6vtKL1XEu1txtgwGt
bNBHQ6H23KkhajfVeOz8dM4sq9dO0MiU2xc+lk5EMu4rYF9l8YQWyHhC5APuvnNh
+jdc4u/c66lGt5H7M/Vl5iMjmWOl7V0MidYP5hYchnHvLmoNyylvdlZe5GCUzvIG
pmyE0osWUW5VYOtUMDbaxdNN99wg5MKieQ6ByA1FNJGEH31fjnm36aHvEkLjSpZf
0ViYL8e8HyAhFfjR0P9ppoAiUZ8UhlI4qIhusMMmxUy1XJ5+DN18Es3CLCFNqrjM
7jAMwtsYMb2eFU9oVtCmUqY99GXxkg2ZxKSfAblRgqVKbKWb6LgwUTd1MzuZS7w6
UmpCk+RVh76ZlJR7Gi2IMLT3NtLLIVyIuCs77T9dBURE/XCH8U+ASBediTKZ+80a
LJyUm6wg4O9aecspWu7exZjzLtP0/O+elk/4MAEKc9HCYr4i5vfnbzTh1Ak1WxkN
eF19r+4xEsd4hGlz41G3DbWwEskmasQgM6U6jGI8aopB4fNmK71/TmsRvZhQAHF6
zvtOqJ9TNuyQ35/4mkTMf1tyQ7ubvGn4bUeVqTV/0dbXcHawaDi3DBj9k+IaQ41a
2mrOYWr0kwh8MdKJhs4uYH59nm0lOLG5bIJy5lxzyL46cF6ZwJU3b9FPzbEU8Qgg
2mPnwP2XLXhA0ot3zLZpVYFAke1FpTePrbQVp/Hyx6m2UiHPhnjNmafdf9cudVqo
VALZNAQ4vYYlnsT2LVJchClt3TlPwD9wIMgiFbbeFFepds/DT4DRTT6QX81urGDw
W1ITGEbSjcTASomE+NvxzjoO9WnPO4b5+m82V70wGqpLYy36YjBSlNO5xAcTgyHB
NZFX67VY5vH2gkAH5NpVchiEpayQ7b1+eHUV7qZHwJR3OiZBXgqUT40z3TjyYCbm
qW8np7UzsWFTmq2cwBjcFJVS8KmFft5PgWq2F+Vd+TxssZXKrC003VhjZPtzVD2F
p2Iw1psmYXIQXWK0hGVtrnsgOZ16ngyxpAc3XXYEn/InH75uwaCt3+F3m7ipNgmc
qo4k35tBnYFwvCUO80tRhvtennQlZ9r0DEQC7eRf9DdOUS/kvKO9A3rl93cPVQc+
3Ok3MPPCYdxbQVVPaMvikWeFQTCozh7LpusaO7oBCXgQwMudsbJ+wdeowPPoDEk7
AifpO1gmi0hLtD3JH1ooxi9clq5ne7bD+ixoa3Z/tnI/0QOVCaIWsciiyONW3ZaJ
wZdx6fLJURffqcQNGKmId8s5r1NjjlE7I4mhz8Ve0IVU6dEA76N3l/CxL9x7dnk5
JoDJHQBIMlo5AXxoeFUPg83mnKpj8Ly7hJZrd+6SMTvMQ+jsT8OcvJ1bxFxj6HDR
+MhdSgT9xPurPw60Pau3oU4MqOQBnZsRE7R+RxeJObJDsOD0ZGqlEdeWuXX7XoO0
beuZbZ2epeQAFb/UY0Tk4KU10FUsJQQlwUCCVb5MWtziRWNSZuLTjMWfld5E/9/L
zzbbpPjMqqnnA/VW3GoC5s6QsU/SEF/1tb0aSN31P+mOXDvM/ScVDWm3Ln/dqaHX
xYf23l0gZiVKMHjcmJlIfFGOdwoJEsSV26SIa10FCMMAHLYpLgtQJA7Q7mo6wGH8
adFc9zgHxNKGkFyehcGysI7Lk1DHs85Y541XQlzLQ3NkpGLu3Vx9oSMwPIYp3EET
UIRsmgxCAuM6zQDVaKPf5ZHt42VrcNlnnC/X5VnuKs/LNF15xlvJ3Xkoup04+2V2
sWW2JGDP2Y0LGWkN4/ztr3TuVtGsaIsjue/0bph2itwhYlXVhTj61gJyAMGiFhJB
q6ub3N1ocAaUeR7dtsuAEr+zcj7HU6PhzcnWpD4u7a2jvy2v7rTX26bt2w2/3hW6
19a7c0P9IIXcPoCUix1+ST/zNOESbqgWBYd+vyBQTNQai6V8dEuscYHAOZcaWVNW
+JoBZca+uRskMcrd5PTJ4D9n8ym+0SQGFeGYjckjwdOTvTkA+zVbuOhmXUGPZkEo
jb1Zzmrwl2F5W4td17SbTeZOLWzMOMCSxW2ryrAXYT65POecqZqqv1tw+QH2CFmc
bgFMPaY4RbkXJcaLeQSYGkXyni8uiK6mzrzxIhjBpGKKXVGqyenhlleRhPxGUmPu
A/XajSnV2EDGw668Y/EzF4Mu7jBtVv+epob2ACdNEyUcO4HuGhXyIfMXfVlwShUl
QG9O1YdPaVzig9T2/CFIbE/JrzmAXBO4cJXd+3RqANmWtfBIdRFAP0qalY0yUcJQ
1uXQrf0cPquVie6w1L71bGhYQnBc8uHvZx5LOa2aWckvjKhuYpMUzKem4XLCzzJk
UqerW4Xi5ng23STnOw8U9bARCWFPq9IqZCQGdp2YYwZJMnDJY9rmrvdi6Ei9tpCP
1Pd0NvKJGsDo72FRIjBGmW/O05ZNynl9kJxZRAXTRNK4t9soWY/tmJFKGsGrBTrB
yaEGQQ0eNhYc2cLeQvXfI2i6vf+jLAVLxEMvSR2+OvdSE5zw1+nSx8bbdvnLte9m
tNKYp+COM3g+otw79+LSKWeggoudGUIH9hybBxIk5HewlhpMm72XJ4t2YyTfXzPT
+Jb6zd7xJMDrIWMrqbEX19AlrlMf2AOeZmqwWB2PvClhE3ub4n0xx8X4I8AgH+Dl
o7cOS3Nc+b5OOKJYosz82fzSC1zNhEn9MwGfJWhma8FSCL6wToX0xmrpoaZrzRt+
FjsU+teuA7bowTCSUypaMhh1cXYJmuW0MsYsgS63x4UHPvaI9XH+0iA4fObmP4ju
mIwQrv+rZMbWUj6DnJezSmzKEXtk100kz/g8VbI7pxSxOTYJ8a0CCdiHDCk6po0n
Tpdj7W3OSgTzz/O1CzJ/YNiyTVLLbhcJVmQuzcurWNnPhM0s6CISh+JRv+OhDRLG
hV37LdhYUOh79csRANggJJPVDuUjjFxLuOaUrVK0uE5tCHQHWOXXCgG1Mz2yVLoZ
3TEnU5pgOsqRSipO+Z6H5LC6KU8n4nKA1bUyqzxhe0yzNdyqcpn/7U7A7Y6LM5II
ijsbLmd5E7aigILrG2FYwzNwthjIX/p3ngUZDemIjeF/Fq7kH2gBmuihw66P8XnM
kLTyGeqzeN/RBGYQMMzgYNV+j2mFO3WGdFinGSWZg6q1sQ7eMGdJDo26dJ4FFudN
P9BC3+q02CrpqIdnh845JHcHjBTEOhxtRPSvRWbSwHMcFqyT4m0DiEdXqZMmbZYU
elnJsXIevlYks31pJ9dN9kHtiWT8OAd4/dPgeu1vZTyUL1jtzssBSHGdAV/RfQDP
s3fSFqvyJqjP35HkiXAcsyI2XjeX63cLw4qcGxfdClsx+V8igSdqcdI565cGIQaS
NI8hX4gh3waKoG7cp153ReY3/+d1bA9DhIrssoSdXX0Xm747Hdlnps9lzvL4LfHR
1hstUt/txaLvTIjMaSPNkZ9WFYmH6hu3Y9gS54LgCwgY7ZZsnnVMU5y+TYQOiUFp
nqcqAJmyYo5WRPFO4ZcQlEQq3rozsjWdOioJw9/U7BfIk++uruAndxTdqN7CGw8f
OvkfYBFaHJIZMr8eCLrmc9FBnpzmWl9QAkZJ3y9icvEMfiMTFYmQ3ymUwRGsaG87
q/c8ucoYRlb2zJaFpxQnJ2FUh1Yd83zAxUbaaIefFOplEjRkA32gFmNEEagGsjiG
R+P74MYoKYDegqywvXgjFc1Uz3Nt8JfIf9fFgrK8iWzTOmWz7KUPo1PFf0mx0ynX
+oJ5bCUYOaHnSauPXDKohHr8pN0jz56ZNXHBHhCUF1m4DLgL+sFm5E2Y7kjyhBMQ
mB39WtKPSQDJ8M2zwCw6kPKpVPXpAk9gZxgprgRWHxb/Vb1J8DdcbKOufwbjIRew
zDTXceY+/b/x7U/caiSadP/jnyn/zzKG3H/Hj7C/i9vBUU601Kpag1e7YmNnqpAU
eFutvwYAaT60z5MK3ge4oeLb92q/wAplAUvs/fg5NKtIAqGW5TEMOOYxDz9yt/Bt
uS3zWaqjI1D7p+SzkNCVhkH0JoQWsN9rbCRxiPDBMq9J7ATi/is/xjoCxMdCvQyo
0g5LBxHpk+pBzGa6DW12vJJXd6A65w9eU8O1R/BQWGWomK7oDFWJP1Dk7tSfHScU
AdUk8XZF9ZiGoBSwZi+ikKzldR0QDK5spoLiC7VnFpDchxeB7WG+ZpMxAfpIHwp6
un1hulk8HMkANX2iV3+xCC4k6IOinFW7ZagTuaM4W7memORQFG2L9TqXktVTjxfN
V2MWtXgyEaBFxNw1aRkgHHHb6y2ZNCf4y3tnz2Stcm+OXDjm8dmzped3r7I/zD4V
W0beIecC0Q/gDbEGFQbN8DOYU/nVq4RTsRauMs6FpA2Nk5GJMRlEcPn10//Cfvxd
/WN8gWldjYId0LDZMgq+mDwih8b5bBNNc7QPgrUOaZGIQ1Y5vhyumIlBL+O65kQ2
7n1MrvrnQo5keuI3B+JLK226TB3sNkRwWkReLT/jvK/3Eg9hr30ASrt3ELjeGf+D
Qqc0KA60LuZG0mxdzmJsNRBW10DJRsi6szIg6sMuJoN2mkOFVAXYxFhmySjaZpRN
n1jLRECDBicc4MhpSvXj7e00JE+eoaWFZcY18/A57pvNHAVv2HAO2kTunWCCgzcZ
Sfeb4U7YDXQraWRZrC51eK58KinVDwC4qQMhERFoeJdO76kbU+Saxezk1xk3jYD2
e3uKSEmjRvDScjREnvG4AyCSxwZyXDee3eCYWEy3n+zemasjT5JDReEF6WIxxvc/
/ngFx9NMvzFLVvFWI4HN1YFyyvt0YQ53+XcS+KVk6tTuLJjUp/vjr4gPtHmcEb/Y
4p10UJzkQ4QzVF2grAhtkJ3ShCA1YcjWEMGXSC+WUJD1JbbeRKhnl8W8jbD/txP5
uN+zu3/+gaxhFMPLxJBVnkHDfAfPvULW3b3fv7xK/1aIrJiVUGAjtWNyIBCOKkkU
ixRrc8jmgdwzyFMwseT6SQ==
`protect END_PROTECTED
