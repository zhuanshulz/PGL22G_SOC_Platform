`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bh9fNCqN/GE8joKNCuaLDAw96vTonsXq+T2MidUOv5phddHOalg75MreSND/UQdK
0PKvHAhFz5Te/2FR9Wl32+dbdSYK0Yfb5UrJbTIcekkhfNcv0gOyPkfKnQN1pIwQ
wJhuKQpQgKrNzS8fJQ68fbrGIpwf5zn5Auigjq8d3XmkH4l2z1C7oHxOHC1WkA7+
YJi34SkJHr+urqzWW6nX01NcVDsc37HrvcqCMmiiCn9yd+3cRD7YHzAIHj/y/lWi
ou7YPDGd3cJPAHv5XP1wUhoFcvWQawKmpta5BOibXFMzNXORwgd5dmr2Z668Uydc
1yAf/Cgw3xWr0SbA5PEd4CytR+tjCoJfrevQL+vO01IvqYPy5cfDxMtFOYYZCGgh
fmtdPmfTW9jqmxuyrcjmvmZMff43mbfTKYUhGjcGhgeVdFwoahO+9Z1JZmoWlA12
Nfl45xkY8vVFS1DqQ84DIYuIXRnu4uOjO5J9+mx1RGHiz68bdJXBlelW/fxd765F
WdcZ4ycnhTy5v/5UNhc0dL+Hg11ILMcUOEZe+JVtbB55GUglaihzuAU7dr4MsiIq
rH0l23iMIwX+u/fHSVCzclpIY0pmrBm4yUjw/FzlxLeBpWFdXTyXMegBJLqtfZdM
RXT8SDgjO7UkqeXs9ukVn2hVvHDGLmRmkM8jwlNjROWNiqQHGvCaNsvZHjgFMJpp
`protect END_PROTECTED
