`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Cp+/ri/Zevakkaimtc6FhK0XQwZMOg6pilX/NOwfex+KEbTkptHacyFbU2s453Aj
U8ELWtH3G+qaSwhdumWoG07PO0Vy146/XBSWoAU8x1fkbgEL9qAz6N8t2WDleT9i
q5NFe/JjCTS1MRnOe3siwn7ZOmVPJOwKr/ORULeyCV7/Y8fpr0ZLjInY0x2sYNcl
mM/PPT4UDHLDcK0KMONasneuz2V/5thmf4xfs2sGPgsYZRG/IPoWs63l02ExDkVm
YUDcmIndo4G59/XEBMqmRUAKvG5Ece1Q+Bfpqb/Qhpl4+IMQ1oXZ97dML8CHoVmi
naC5LtYFkppP2FfuW2ewUmb4TQdf+N7W0hTj92/kZwFg/6ipP/dTl2GyegC6trOO
`protect END_PROTECTED
