`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9ND0qRrvLioV446He/1ZPI0y//sHQxMqCb8bg+Z+ekuFd0LrqDlIJjfs1+jZe2Zg
+8HZxi21H0P7QaycnxRngGqFxpWRBXhtBzLWjkr/gIn8pLL3M2aOZ9cq3Ywn1DlM
peoW9YGFVT2VCY+c5p8sX6orTLN8ZSQY0PJIVKkLBkJC6hoE06bbR7GgQu5S2j40
ThRpcmyf+P59NUyTO5MatP+cvOYwOaLQvYuP1wpRo1dxuPWmuAwV05Azfv7gfbQp
gfen6JqxbL4gz+/JLEkDIdTzJoAw9KuoyE/R+22xByU/AOu42Ome7hDllBMMaTho
2EmNUZlvUA6ksyGpW0+UaIwE7a2/SoH2tdf0DczmDpprTqvegLFWZVDFqVHjKiBx
6aeJrdhwruXTyYiZExtKtRFmoQ6tlUTeDItHEtuCjDL60KYdUgx3hbzHdIEbfD9o
qusyqxfShcgO3yvf+d7S7pUVguePy1dJvevnDYpNkUndI9/oyv8bBMFKLkoLxAxS
1+aOYui+jX1w1cgBZQAmuvY6vf2kx8NuHOXlQF8xKTUSzlAz2QcztcNcycphDWCu
eTiDWLGhJd0t74EIo4PsqCvxDdbIr8eh5Nx9abaG3N74O45kSgqCJJFj8PoL5cjM
cBTo0i2GIqIEXwzOxlf6hcT18Vdvu4OIOp2WBhrmK13dZ7yrN9LtHfEptfVQ0cNV
fuHj/tpNKctCxzXi3+TRO7qfxEEIJPXPQngOh4hbMaaCebzqUqDrXFUx0hULoGQk
ql2VJI30XXDGrM1/bfUpvf1la0qWu1yrBAVAbKZ2TK4p8wb+StkeueWhVtRUR0O9
svTcGrcYQfChNtA5vYGJ9omsIhqoi0BZms0TBYDZpMnCK07j7B3RaSdvTxUKCvoD
ufbDnwn9cvc5ToYM6hPk8NTRPaSaJkjeYCSoWmXNC7ZJEytLuF2ltRTkSQGyOhPu
mgkGETnzc1EHWtg6h84hNS53V4paGwiTzuNcSSScNAZ6ZrWgHXtaEUjSA69q4Vfu
zr5lbubvxbxjopFj+1mZjM1/6Z8AiNrdTm2yNu1gWQMYKNxFQ6rTQOrlgzbKCQTW
E5STZ1KNNetVzgJqRrPxjogNQEGvnrkJV9vG9ugtfy2E38QfECwjH/A0WzO6+6c8
lLpAh/+NIW2EjaY74bcCxZNqWY3py3JCPubhtxJzPVUcMr1oYzQq8yFBvZ4yq4d3
vIFBWwvj9KoKgRiv1ze9W150Lfc1wfl9DGxznIjuYrHYLMOqWicvI3U8L1FlDICo
/xXzPrCvZ0aI2t38IGJ6nHWA4d3OOKtYeexDk8S91lE3+LXX838ZKP910uqv1y4O
hpTf2XGi7+SO4vI8kavE20xl7jO3CKDHieU2fSvn4WQRC56m+lcDaq0ndFkyf7G1
Mq9nm7aYzWwMyk66/Dx5+6E7liKxstMG/bqQ8VKhf8qyMqh7k+1I5oJIVAxlp15+
sC/XjgECIXjySTw+aXunwWJihSo0Vp7qnGZoJor92v1Cx7R+jOycLy6Ir5Oholn6
WlUROEmbfFPnjcWnCcylzGgLhOzIpdjpQCwfVMhYXQefEz3xfePJx1Rn19CLkMdl
73Vvh2gpbGkA/dqgezWwvUMT3prXXdx9AAeYS0kxlKpBcypQJ9VSrgnAReoxTcBp
V17KPbAt7UEM1oBc8ZqBa+SMmsZX+8/lx3AashMM/1gSc0OB8om1Q2VwrUgzx1v6
C93Z7gBMel8JxK5XXOKUskjewapvdr1LvvUihsw/HHvR+bTJwB3PPMvtaGF3XJWA
6T/sTmFYXJoc+aUhdQkmNh2ZvF/jGkZM91botaJuPIm5OQCJXXx9uCuG42aRWL/C
DMts9ewhjy6vAfvMiwh094dd+410OJN+P7jQV5COnm6OEpeUCoBuVGpxJN06jEVi
OhFz2a+bl67/ILI0+aD5eoc1xsvkttee9Qgjt7aqabTzjB2Q4Lux/cY08J+PeVxi
Hmy9zNGt0iALZDa2ge3enuyfVYFrfWiEDC5qW9BaYKQERqR4+lYwC5uoQgOC+W+A
xSTDuon0DCjo0dlfaQ5fWxV8vjvPRvVNL0BcgiAvhg5um7j1+XvucL5JFxnxQ0qG
g/jt+rfP4T0an8byuSTCjonEbjbThVWWZ/kYcYJVz6H49o4r6yo94Tx7rYAaDpuw
ALeI2lsB7BfMLWRPuYZv7XGkNSgvUSB/x+tkU4vNrMYEfBxm9ZahDIR3kzHIjsQt
Bh0RyNyQPB2ctYDZsJVasb22oZBIJClF4hsYKAf6NVqYDATZres1a/TfnrdX7Z8F
L758NmB0pOb2ddxJUwmpxdtXacdgx6qUVT8toeZjQcfk+jKLWwFF8KwGp/sy9PiH
xOIx0JWs0VPSbR5oTeRrNqd1XqHi7qR/ZH4NqLlmY/NRv0ergamuyfImZjJskAv0
su1X7GVzZhTWeNP/xNhNaaaz36dHPlbvNshLmNWfXX0rkLCsJrRPpKxN9oGC1MVs
atFa4Fbs6eFaXBzkSo/aMXMigkZUrz/UdD69TymrYRKIO3hBreoVSDY3vwiuYSMl
EpIGSxSqEwLkk0dh6+fICoWBcGHxRiUmY5C74Kt7Bw5myk8u247/bBCx+ArjZKLB
wwQe87L4n+TBXL59aA9gOEB366gwmjM6xXa518Pn2zMCrLQ1Go9FcEEG6/GMtXkz
f9e0SwJgf+bT9Vkj+OLBNUgHYEWahTJgAB/o6IPPHszVDMjJEqMgrWLwzYo2Phyf
yOjcWI/qDPJpWAAjUbEtDTxsu0eeR/vF/J1OwxVf/GpDOUs8ImDVBHF7iG3W0wgt
zk6sGPDHgLK4iz2k6coZ5EIjzwkkPHS/79779s7LDcr/ln8v24RBGPRb5ZJv8s3v
tLN749rMHuu6iVajnW/9Cb4NIhcH4wFed2NMUcxhRQNVkQ0QRtZogtEOaERj0gKp
y35953+d5SbjK0Xbz0NL8UbTbdQ4sTOu+tSHFipNzqLAjStvOzyTT74GKbvgJCdy
Ut/iLaW+VfA5NQYq1VAs1lECqa+aQZjUaRs4Fjptt75Wyw+dlUbkImElkdazRMWS
lhrjtx//sMO2KcacOpMBDYDC58LQYceRtzLmtwOk6+33UhpsVmiPxZgSuHDUszep
6gfMQfuKahYe0e2QT2I7OOUkDKrz3gIRVYI8NtrpOrzCV/iq6Iiv4mB0qx/mE1xr
o2XJfvB0tiz0mWDab4nDPSrxk2O92nhgXzVYsVZnPixFmmq7WxjvvL9HqYiWzms8
s50HfzfwdVTGYUoRrHU5xFcdZ3wDA7wtVuj9c9L2bSQD6tgDHbxtvYeto3mNMTMa
OvBCxKCXJ2rmlzCn/n+E1mPk/BAUJhBLNfBtGrkV/5U6/UnHTgHh5rOChK24geyA
96EmrNFFOs7IQAMY6yRTZ/nWzqTJecrIUojYAjJyLr04mOZzs/tmm/Khbv9QPIR/
mDcuNB4QsTUzlzXILCLx8NUkPN/3rFO0ZmX7HANsQ6k/GcGztQMxVjvAY8GDuFIL
lG+2ENh31kLdzH28FCPOGWk41HQOjlwksDO1CuXj5N7/kOnCf9lkSloGJ6z5ce/L
F4Q1AEFNDCZrZIG3QmQRQWuIsDb9zsDzv6mXqPeGUL0CLN36RW3I+tQi/H1fYTN/
BvojwoV/Icy5BuMcdA3pH6S1LLATUW7lH7b+3l9+1El6jnlHu67Ny/dqF6GUk3Ns
`protect END_PROTECTED
