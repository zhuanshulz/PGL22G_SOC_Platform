`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SeFafex5or9ubmQ/U2B4GBN0VqQFk+ffO3oou5quFxIfrZG8LlyTbfppANUp3LYb
3sJTW2Zip+LbUbUR2r4IOdib11P1/kA6ThSmUoq5Lm/dEsqAWUhQHdfFzM3epwfy
8helcLAfTb3GIHdvO/ovFnXMacJLDHj8ox3MVpX2EN77vUlV4r11Cy67BRgB5Kyi
HozEBJ3gEkiOLhzrMubTxzw7Oy7EV2bz4gXV008A2booVFXh4kkRzDi+xWebX7cq
iydrBYm9x1qH6abHB+dV25RueAAHp/ImSRCNY+9MISV0xB4yPDjWkJIVTCKBefWm
56XrGBS+7unzb9Uuth1ZVF9q8uu/gQ9M/lQGKbNl77CQ1+1YQN6Pe7KT2ijCn9mM
0GjmdodITQ/LtD8WZ05lsA==
`protect END_PROTECTED
