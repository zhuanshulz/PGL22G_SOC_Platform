`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ji7lakjmGYWKkpWZihHc001nS8Xay70t+CgnwdiE5Zbl916QGuObvWb3OIO8rRrB
xGeKKB/G7Z0fCVAMtrfx0hkQhv7k/LJv4nAGLBTJk38+PKtaIE4tBgKQKiGti1TF
FLR60fl0CzZEQdyGkkj6ECiR3uHjgzmkQna5+SoY3m6nVTloT1XPTX0xOqHHT2sF
wzW5NtAlLBn4OuqbaIHogDgrR9xrUOpkZ2Ue39nNv/SyLwdOGN6P5NWIaAc1Z3Jd
ccIX+gOZG8B9C07cHn9l+hA+TSW2ZeQOemgHCO/eWbWMjtwO1S0s21ufyGAwdjBN
CYIbr7VPc4a1zXhwyTBbhxISztuqpqKpFtnlgWeYrxN7uN58DHqkn9psrc+xsI3W
o7eR9+a8vInsoTgKkuheyA==
`protect END_PROTECTED
