`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bu7WESdCrNeGAXOs8kCLh3/9OOjElpinXSmEuo7RWUqH4B04V0GYITKO6vSdeYw1
4lvc9YEbi+8K0ExcKSeTaME3mMpeeCTZlxt6/6QSlr3Pjq5U4wxoCZWxvTluxMs2
icgonBI/i279VZAyjIKNSkC1P/xZEcsnveLbQ7QIde4cQtcO8qWXlNQgKcmAdsCd
x/El2MTP4S6TQrlFaKggPOYGkcaht1bMYDQ59g1XsBjMwuAqxETdi+Pj0AWnbftL
20XcNiOKA+R5nM7HK4uRZW9BPLh3JUloQRF8gH7z6iMyS45N4EyJeOjHZ96APnX9
PGjxMq5e9r4tXDgI5Uu2iccLZPzKWVYshn6eYo8u0ltjSg/RvcUhHY7DQSFQ/b36
tWgvl2ImAzcj1nflC4KcI34islnIpf8HCHFfLDdoQ7KIzKUhfD3/98F0XxN79/bN
4F4fbzSYVqFXdXt6T/+YZHIfttl2m5MgvVqLi/UjkKY77+GcRG04elj8pgvVM0h0
hPincpOW+YQwYI4KXTjwXVnEOXZ0PEuhXhAs0GP8x8R8FpqkqNquWO/95kX6IYNZ
igXI0gWicnwLX8I3l8n9knLGFJkJRgr9hfSdjkR4h28uSn897VCld1209OSikthZ
/AVbPPdCuSHXm9tUPJ7IHTgoSxAbdsZoYTmyoOPQwKnuhuy/lRONGmTPkACgZ7wZ
JlBrmQC0bZw30yr9/ht4KbPgrJrJozRCUv01MXDsXoqNLg4Mg2noKbPKlYLRZCxi
6uqZnbA6ZbwPVjzLP9ces1tYl6ly+GSKfDryPT34OcVuLPmG5wAAgERdax46q1z4
JHocrz+UcgGN1IZVh+vDcTRFV3+269eE9bnpANU0N5tONweg5kT+KluSIiwAg+cr
ruu0mU5HP6xT279mxCkkw/i9g2wGtAR1nxI2or03S4i54Xh3Q3TZi5uJMbix1Zuq
lkqqWhVgzVI51Wwcb7rla0VBc6LqAHamYHvp5DnE5YCTW8BMi61Ox2jILaxjfSc3
nsCyZ8V7gkSR6EVsYaczp01KsyruLnTmXwkwYazSSe87cPUsjKLP/2QaczStLEmE
Z77X2sckfPpnp52yyYzWQiUq8/KQSsuPp8lUwzt2ITeGmGqVxmHzajo/BtYif/dj
Iam5LKRCnW9kPsewrVBed4z+QI8hmYG4xlDZLDKPR9rEUHdi9kIiJOhX5086QQqB
Hs83Czw8dZ9w54578cgPtWdcSANHkwf91ToJwZP/eAfhyOfhqE/L2E2Iy5q2336/
xxxCeF207FDBcxnj1N2qwvFp6Mj59fOd7i4cfGQZSXRAAh/iFfmS+OVkxKC8Wkle
ilxtN0CUhlwsenwDgdPHWsoCd2FKdcg5YoKwW14LQ9w=
`protect END_PROTECTED
