`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fdW1E6fTA/WxYzW43TmdMWENB0MOxOWkMjPvTcs2mn2jgDCYzeO8RIYWYE8OwHGx
d1Z62vVWCzgtcRvwrHm7bV3FyiGV7Agqysq+LU2odJs+2JG+BWq4S3p2k/cILbXL
hh/2yvzlI20hwkcWlpeoVJNuElSbojhKpxZLJX/5VFNJQESi4duDq8VmuXItX/Sc
Ihja1OoTk6eApy2reAfTP2hL7g6gaKVyAymolhVDWWbdJTiHVMawwURe6UXzNFGD
4993RRiEnXPRY8vHflRXbQ8A56Zb26NL/NkDCivhRevjLDZ/cYpWx1cOZZda6Tft
NHImZpDJbmEYwMUtjA69moOuKduVP7eCDEWxyqYMVvb5PN6gWZ0mj1y+4YOi5jgQ
BdBUo0MyNawIEZjS9HBuDfaVMzSYVS1W090/ehBQS6PEkp4aYJ4VBGyXaqx9SgPD
2GMiiEW8A3UubvBOWkkMcrHyYIUWFoghjAx2Q4IwIFvp633N/EvFls3THI1Lh7yr
Njhy40AG4ZOlcYHjzw3QoUMVQZueJR2SUCJZB5fnNG5k80jXiFYgDTxKid6SEuER
wKix2gE0ZtRPbN8bFPCFSsR7CKjLX5QquLP4Iq3Rjm0C5qSz72KdmUzWJNdXc2Ux
zk9uTnX16VVlDk0YLThaG6JBpw8TNvv4+szV5V4gu6+H+yilHNCoXHPNiE0TAlNd
W95MWjv81RC7qBLXKWOFkKxc17rKvp2ZhsZ+3gcq1SbODFnp4Hhrgm5evOLMPEbF
23nWCYd57lNVCD7X4pTOLqb2/kBSaHApvpU+W8xpk6UUTuot+2D30gr68sEP0uH0
NvQgRbpqKSnqwkutjTK6f32+WtzOcOCwJiGBiiQUfZKMuFLpY/wx1Gx3THE7yAT0
p+ZuPcxE4eLBNlE5AnRuwblTxfljpXCnwM2BjL21/4sr5NUvJdkLFI93RZ9oiRHl
OQP6WlULX4pGGAhmHcpRB+QeCepwKBgNAFaXdO7bbNwTscfhZeuRs8Y7y9Tj+Wsi
m4Gi7ByQt3RlfvgO+HZIjVI3u1s7O75rieZX/9pZYOkqWVpnLURzcPXmQ5Ky+JcM
ojwS3f0/s+EZUmxPPdGK81XXnp2+pywr36ZG2qJan4jNdre/oPjTTgI7UKsQkLGR
MoxjGgtMQiDUz+8A9qylMY/1UahSkOLGLJAJyudLcvqDuq0zhreXxfjDJ10dCQi1
IEvAyt39jq54SdRwTSUveqaEkYVZOb4v+oSxB4CNSOCQNkQVSBmzWn5rU8kaeQek
F0jFekuTYdTDhQErSZL8CxFZgCLf0GXBkjrMRtfb6roUojGr4cpLDIAvg0wYQrcZ
MOUTsIawtSXthwsD9MAeYPGBuHTwnEl0FjIrfs+7S6keYUCfNaUXYONnIGAKx27S
ik84wvl0WgKn7sHZZLf6k3URiHxLe7QYpMmAqu4WkN2a8tbmWY7+yQDi0O+LrEbP
8hHGsluWCCBdqtzA1Y4Ap6qTcJ8Auo/G7Mqk5yxSYCDVJE0Ny8hRBN5He+BctIL6
LppHrIs2M8gZzhgU/E1Qh1K5q8lkMCePUEmkYZ8YBbWCyt9J5sT8WoSsAq6XfWLj
QbBa1HR99HokqUS5EnNo8ffo+6e9nOBmPksRq9G4A2ZNXzJUCMRceSrW/nvlvjdP
62QMYjmJkRKbKY9q6SQeIpCbgsfJR2tRq41spAbPaFeZur9E0/wLwEZOcSQF4kjr
hCvngLFCae6n0ZUEzulyqgNv4HfW3gMJzfxBHvUm/Rms84geOaSkaN5P9SwkvaOc
ZilDyBiHBqBQ0NnvxupM1UsAapRMk+SFvKnV07FUpuclNTB/ysBwP+Z7eaMlx9vS
FcbRyhrWZlsdb+I7VfkKJH58v+Pc16HYj4HU2SgoyczpYWZCfoLlKu9pXdHXYk7S
yxUgmUY3K1gJPaghTBV5bAQIJtQBhky2HGtLmW/+C76PcgzgXbuTU+yuK1EZ1JOi
sl3tvRIRPVftfJyuQfwFAUapA1qQ69wZjpynd5W3ZQbW63+/guOoOMt2NLYodFgJ
LyYtjEzB8dTDGzKoPpr4irMmfGmbfFhj12LjT9nT5b5FY5FxLZYQGVUG2OnyUorb
JZpnGXVRr9U2zsNa2NtoO//GkqFfpccUeRBViPPPWmFztouLeXzc4ozrv22bf5KC
qjY2SV/Xd21gG9vvO7uwFPIOrMZw0DGagrRBJ2V9/bHUgMw4bmywqEAyGwY3tCj+
ozyzMmKvUgJdPKKxKz48UnfQygdQ6xPHiRNf7SbgHERzQvQq1/i/tAvvcWPCLwBj
e5YVXTFqMMDeId3I1norTIrz3J980BlkHEBO8CXC2NhkbLuRBaqQpkwqZX3rtmFQ
jXKoxw2F98DHpe87N1JaJyPHJ8wG1irEEjJQpYMuc4ag8yZSLSJEAddpUrZpIK5b
etLVixfyFEa8VPQO8X1DnN0UELm/z1ArGy1vQv5xJ+nhl6xrqoOpulN629usKdqE
SK71huU6NGa2KNi4px+IglZjArFpn6j5fN2sM/3AOCmCTfH94hYp5gB67P2GfiKP
e+kvDahMe3AtdDJI2tNQ9tS87AF3gUjDH8GP/sBoVA3ddIBc0FbnaQrVaKu00YAU
ir5S4tK/+crJ0iMluZhl0hjC6FkfvayOvUqwyE3M6XCZWCt9FxNbJJjVJAtla4Se
73hBQ++Uvyl0l2yoIlctSRxr75mBWnG7MicT+2OUBOGx3S9fzgsTEkK414IXq/8y
/3UlUJvhxAbuupKfl5bOYyd5Y7E5+o39q+7WPy0AWDViUKWrsp8iFc9GfN54ca2k
peBsiMhuYZop4mLAIGZd8zYg5lGdtdLsSASgJ+8NtadkIarb9KvpwD1CQJX4wM/8
mFioZuOBLqNFkuAgxTayayUlghF4vVnR5d0XJq2UyT7i6n9e0clWBHxMa63ChZ1E
X8A9qsaNiXukdw0+xS0iIoXjW7XTkGsoElbe4WSKgQry7PW6qzuyORPSHVL8gY0y
tfKcR0n8nID3wWWQUyWI9eSlCChEb0tRgDP6CIu7HyeAyN5I1oSTkM1eWO6FcQv1
9lA3Jjalxnvy6aKZMlKSUMQD1KHGthqDT6QUWiOa7hPDfHSwP/jH4mbVM8vRCNC8
CGK4EcB0Eh0hmM/oiV5sK5WqDqJEk0ui+avLIFJoYuITl61/uCynf64VDR+9HgeS
/FlYOwebUh/gGWNheIZV3xuEcwaS6llj89MZQXf0/ygb/mNgpwgckMWPOco1GkGy
E0wytqRBazx1MqnUtOHUvh3S+FbwP0GA4busM0arwj5OwxQubXPNj38ZyTZG/uLy
IA5EY0wnYgvcZ5tIV+vxapK5t5fCl8km8bhNa7yNMDKRftn1b8KDhfy3czsO9CK5
ENHdxfZ1EoINkQq6Il7zUTjXGknp88djIX5gs0uuaEDjqH/eUKE5J/MB2r8Z1tdX
Y+CIc9ppNT9tp9K7U9a63nYgPRMNRkj6NQxJdqoILV34s+1F4FVUOaJxPtJy+n48
GV1OHKsU1h7odnyj8O9HEUQSjM6eXN5Ngvr7wuuQdZbgbBlE6A1m9HIjjpqh1zGb
Mz+WuOoYk8Zo/LU634e1mn8Vjlx1t16+xEcu0kQceAL2r9MRbWmTvQLPCNcffHEr
yZsj7dh+lyVw/hRNn0vZhTkuh1Lmegu2/uxRbW8676zrwdrgNlqO9RgW8IdNG8ho
/jztUMrU+KHV2VZxETWQSpFjwgfTZqRPnETfA0vdF9ASMv+PFDRtwksF+z3kAOrS
QcF27BUPsw8ff4kj/IwaRyHxJ0es+6mj3Y6vIVGjKBrI/v0T9WWAV3vrWfwFyNG9
74/mhsROTwmdTqBtOHXDPO7DeFMhC2DdPF77r2/4wkyFMZBFMf8dw22ov6gxuCsR
+xgXFEs4iKSC1n4kNXmiGI+AGv6g8pitEcI0Y8ekxzRlDsGd5j09uBOQzmP8eZEN
zUjKrin9JiMxm2Bnex3Qa3TB0YTuzH0MqeIbTkQ+z5zaFKKpgmKCjEGCtYgUEUSJ
9RbPDI6TX2EU6PKuGYI6/nfN4CsnLGKHAbzFm2vpd8unY4Q8oOoLpKyHfARiPhxX
txdlUV+puX2Y7AU13l3bWO/JH+b6U6GEgotYjkckWvYc7N1ZrlvJk6klEx5DqXTE
V7UYNMVOopD5v+lpsARELtyAdQTBH2Blbg0eJ0e6Av9SmmpL1WxLumLvZy7x1Cmp
3xFHe4PJPgKkJmUlTtHzWw==
`protect END_PROTECTED
