`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7zcwkWKGWm+s4t05tzu16v5DGIcSkN7mYsl+JPdo9iv0VN0X/+HUzXMPGIlt9i8I
9zcOk7KK1ee45Pj6M0gNcJbmuxw1BfHklqzbXhEzq6PUvMhHC2DjvEa+oPRBwVC0
elKCRuTKN5e8S6LeAerb26ua2ot5/TYRJbXdD+zn3FQZJTzxHcO5V4n6wzVAvn1f
0X7Xb0V82OG/G29Pic4in1ebEIzUmGOKVl+dpTSJmy50yBHBp88d76GNVon160oD
OM3VQtQ6xTljP1YmEO7iR6I7PRO1GkYxeixGyZ+9TLXDOvWk446my09TsPajfuGA
yBdZ9zqlZmbFK4wXyg0OobIWHAMtIomZMfRGGvyQ7zL64U7XauQDm1IZJB2ENd7T
SFykn/1q/NPkinM1iAAsZ1XypnDLh2s7N3ppK5S3YZbPQoOzN9se5eGq9hwfRe2A
JZUv8QBx+eyyNZHMAo+S3SQXyaWYv4dWO+4rCKs1NUtnJiAEqba6UYOor3O6+W8+
3tbvkYobbCFR5REmgOxKV5cMIVE+o4/4J26V23Po4js4bWIXlS9HlCAPnDVYvNed
fTSEHz53V0IoWRQ7vnGFVw+KG7xunSVZdS3l7agM+QAag2BKz6Kc5CDn0913bBUY
jgrNCupsNnY30GEQQpiK6wWl2JNhNWpI0tfdQxVyQqECWSHaYAz+N10RLCdOjr3V
4Hd0Vdqzzrxh5LVozCasQDyW0s8JytyuW1WK//Hbd9eQjLv9JL3aVWxEyDXTey6D
gjyfgQGi76v3hWAvzcY6lkrbpO7bU5Id/a4uFvmCdqSbghZLHgnbU7EyAW0J11b0
RACPKzE7TFtJMsozXnab+KfTVdeoBAupL+EJ/BJ1O5WJXIspHZTqfN6cRIwR4/Vg
CvpGdHN6UTZFx6XrYqjvZQlIJ3VQX/9w0GX8gW1yX9z7aqFA0Ap4lzlQKNwzQryM
2zxvU6nc5rqKbij2M1oOMaYcCZ4x/F2dFxzeFkgtlJN2ObsaMNhikh7Cu2XD3LKM
oYFlTX41lXoxfxBC75voqbwYdmq8Nh1HjAv3IKdXPKFlSVLLU4Ra9mq90OrYbQJn
S1GL1cJTwa/WPwdI0RGlL7rEVXYoCr6139aXhic+8SS/uUE0Xjnu9+toI3Op0+pS
VWX4hn/0VB4SmafmflO4Z7LsJ+hRBhw8PXY4kkT0ktfhrc00IjM8dg9FeLDFAwxx
2dwE2bQ9UuHUFKytJKnxLWu1vUnoLQfVqSxBlNxFrORSn8niRN/Djmz01ZTQ3EbM
lBAZsoRYaX+zKh9RegPlEcGy1d2vKOgs6T4RSig1Hegtu+kLXIPbiSP/5lunUT2Q
GYuwJh/MiwwMkAByL30aYRuRoD7YdVRd2s5rTNNql8jIZMvrwdqmWG/r7ir3MRvM
7A544uDNZJTey9KcnY/8kJRdAQna09N10xbjJA7bCtYXIJ7QqXBsFdtCqEN2lBhZ
xG9YRp8joqGFPpc3oLgkVDwVcIUdGLyvo5wcZ40TwoPXl1Rh8frx4rRIRpZVuvmA
gExaSVy7ViPrzymVMuZVzoPLzZ1kOB8DEUYCPYj+M880GusoNLTlEpJkjXhED5jy
tv5E9D36ZEXGRWT2/usPBk1Z+xOUjQy7KxBDaF6/JEdDuQVg6uJ1zO6+nV4XfgMD
RBm4lG/4jD30RQ3Oef0JrKhRcOmn/kY6IofdSDLGo+rzPtXG8Ek+RvaVzo+Axp9e
42BENzuucS5i7cjrMpV5QcS8oUWYwjkX6Z99PMm+FA1fdPA/f3GF3tak74PYBmgE
YwumpdU9u/hNXM/GcJ+kySN+YG5vm1JWv0nIgx70rgEEHiSurzG3DVdgcNW1OOm3
DPvf84A01lPRuaDxa/Cc1fZk1g05WZZ4VzWFXArdLbOYU0TfGeZGsDOzfLD6QQsD
wa8U6NlHnc8G9x+8K7Z83laf8zIkw5F6Dv8gPpUsLNeb18NyXJ/MhFgEiwXEmIqo
FWf4lmpSv3HF1BEBYerSz+lEzVb/X1pX0KcBmhmwnlopLGieQC1RKNGJRrnW+J8I
LOs0OAhsGmY77PiFr2KGZijYwu2cjhWlizKkvYqZ7bHsUhBBcwTA+L0/6jhj5g93
ah27wYzdxASMlqLEWdTWM9bZj+J7ZhymlDRun6g7R6jGQqZFufKsmhy2SrbIYxd8
W1nwjm1XeNW0VwWd+0cI9nFR9IRSbDuwn0n1d+If5k+3qSfhV95zPW3iXuRPJzXo
hkTuBgqj7OpDKyadyGOfGeQgkvg0LX0OPnWVXF7MOAJqjQEpLQRb1Wwh0X4S6cF/
pWLf5OOExbscus9VNRltCOuDSlJn0fF1rf/dA6OYWaSbeR1O3FCtzPzDhysPLF3j
8dP2WEnGfe+7QO7X4Z8R8L+WaFGID2RBKaUaf+YOGykheHuC7Lg7Fj3GnFazRFws
Rd4r/2IWvE4MdlSNKxdSYK1mlCPrPACE0uYbCt3ElFbJNkQn9EI4rpVrB8lkoCtA
f8yYkrE9uhJaxFRFrdY3hGFf057DTKfomKoRK4h+wbkwbm0DDKfAszL1zWjpOB7N
qKPRfDLTXMddPQ2/0LuEaSivI9sFQyHBvG1duYKHY4DwhE3CIpBOAivMjuSJegV1
+S4ZRO0J+Kbaf8/ITV/c2kVhIO5ZI23VYx+wrzfW38zpNrHnGfZjsKDEYmGBiCJw
mvndsnTRoIwx6Pw1bE43jo6vGpsF1QXfBYz1xKoeOJ7CkU2c8cqeUCYZUk+rCWik
3aOGm3dfg+NIc4qpHVaZnVJ1/8MftEJ/1U/FVmunIIfG4B6kZ4tZeGyZV+9duEhx
BVtZx23soMoy0v2wxNoPYagyeaKVChUtWPyqL2jdX8Z+s6ER2igV6lPUoEAJQOYe
eMAQWShgHM1FfeDUX+EEpFNzGHLzcN1pFPAWzO+arJeCGs1gXRYbOAcvYnUCc62u
MWv8jzmTxwHUsKletFobbf+ZtHPr0q+LLNuaKclI2VJQNdp/xun/T5iPEeh9rdIu
KFAnsxY4hgZDfnVjdf1833FsfuF0nShJPgryL+UNT9ZkBQDC3utLv2lzS4RmqJwu
thDijaO15YMcBXHYFcoEmavCSDlXSVnNY0MmBgZrv+KNx3hN/9EYCWYMt7CU3uCD
/61J50W2tRmlStUi0kNXUmd8AU1UyLr0ZIQtz1iqdn+VDHFEguVnaS72wmKXu2oD
MCKkkLdOanQLBIDbuFN6SgfzZhasBe8DzaSmAR2meqAOBgD592Qx9P/pPTigjAgu
coAj+5HzEyZFpg+Gt8rib3d+kWXhRqSSx8OZ9QCyPgG4sfPBoGnbogGTXppZC0yW
4doos2MYc63zCT81GmMVH/BC/b+JwPjLlr8eiKca51lwmWbkQazY2P11YmrqHHxz
fBE9uciPFAOpTpGqxM2F3mJfSnLmnMRWnJmjVOvclAh9KPSX0cVNoDRFeHVeBtX0
s77ziUJ+Ba452Qcox/EZmDAWJV5LyaYayRDrxuZLpVwAm/BAxWHlRSFKkdwsEGgV
2Ui3P8jYFn4z80PI8LjVXGdUkF8mGMGamc7w1qdwTo1P7jrlT0A38ofn4Vv+CkuK
+2oZ2WKz+l6Q6tU1E0UeaEIzzKjdhZw3Q9y2zkVBSF6+S8rQ2/8r6eYkMGNAUCrp
+t/w24eiHwuwa0PJfkV2avs8XXLSI7r+eidWuABDcrVeCxOtPhiqLOg2rw1KLVEU
7YnmjDuUhrSfOJVDbT9p28AlX/naFo2I8U2Pa7xg1AP5DXSVz55Pt8g2UObTZitf
vV04DTPj6UBYUPVBTSZBayMIgJSbyAi7o4zLZbFLy6CEj4Skff7ELmaWZlcs6jh/
ebTQa0ufwN7RRDWf3LdZHGgsjwR7dCFTBI35/K9XaVnWLSLEi1IYh9auLtgy6MEy
HfkmSxDQpxzDD2Itsll69Q==
`protect END_PROTECTED
