`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R88X5ApY7/yvsxnba0hZ7PZfgFSreq5or4n3D4zDgziT1jxdwjhsNHlBXrVzzXYI
lGg/j9KHqiOTptBNZc4wacvtMovCGpO+/rKt274YQzX24lUattjAi7yGxNBYYAqI
McL+mCOCazIMP/UMQD0ruyKD67guPM3kEQ5BnXFrj7dVuVGBctt/L8ens9EDJLcm
3bFX5FpxrvlEFuP9gefxnov2k8WNK/lJunoAe0YUqeqU2lpqsOTNENMx7nSvzwq+
DgKH0YNqueaCzq6T8gVtg/unFR1VKeSAMsoY5w27/HmP9dyZ7W1dpuirwhgCe/Q3
QVLu4PsDKSqU901SBr7xveoJCBRso7Qgwpzg+XEPYmdjWFhkatQKhSz4bmxx5XvU
4gRJ1lbrlXgagPaSRaOz+68L2r2B2wEY9kabfcKQgSM9JCVvKe3jD0RFOrocVVDr
4KpAiUcODxJbnMAtUnEtC00BmyoR+xd7Mfh5hHcNv8XTbFS2Rg3x+0w4vI+onWK/
HPSW669QO3vXLilwATrKlKh3sTDFBgyz2tTYlUtC6jHyyHikMzjUOh23b83IpqFa
pHsp0Hdt3nCjCAAqDd9nBV+BEo2dEekJpO3z65MGnAblrkEVwn4YYXLfSxiEDq1e
WEjDL8kPL1ctrtfZcwtf08N9nAsOMPVi/YGY+psIyBRAT1Upmj1/9bvJ3g+ich1N
3W+Pk92zKAmRYm5ds4yRoTlRpAq4JyYe1yhrwEO54A8LKm45rvkM0xJn8rFhCSZS
8D+h43XGjmxYbSBACwKPx48p2yY8Fgs3X6BF+iG+xugWjr2iJyIgpRCrS7pJ6AzS
14VGUG/m5pZN3VcaJbDsOgZ60iAiCcBr5rKgJSxTrbA2R/49CXPUfYASyIhaQpOf
dsxSElAkQ9jl8xZKvkEiNkHkDbLa1QErZKlIsfJRldEousoj8YFAkh9bRmLrfOM+
iGVZDUoj2I9dZSv4m5FQAt3j9VhahCrKWte/G7MmtWJYNO21ZO+A1zjYSUKpMfp0
pAXmrZC4JUkYiaJ1fiV7csyE9yMJuyxz+rN2cVJXe4X7/0Pw8Y+qAmnulMMFLw1G
UPoIKDzEkp+IcoopamaykjXW206DMAazc8rhigcMDi4c4JlBL2gHelJL24kTXgYc
`protect END_PROTECTED
