`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JD8+gyYy7F+c05QUTbSZtZUK7sYjxZOwHZNHdQcfH45gmtkusplW6oc8hB78mWJi
b9mAOW6IYmywIGE2BoztreRsTGdUqS/93AVmUyFkPjMK8ij0rW311nacGjqpsKRE
P6/AjJHP/a54peOspsdCpoCt0njqKrszAgEh/SlAXbsc48HoVCf+uZMDad1Q9E9k
dLRvick2f8bKQ8NUOgeuaEN4AXOMf45+3QADK7+bccIYPR/4J7b5ggXgu+Uiltx1
kNQ5AkM07ul53/hCQnn3jGNiL8WS9sFgW3X3VYMvwO+MykPa4FQsJUWOhSPFohgB
uWyTQSH9eu/0dcQEOmWrax2LYDoJdwIa2sLd/BzrIok4x8Kp0l/6a1ISiZgch3zK
yrPh3WhgZEvcmMiDtmGIItzXMZuHt17gaV2Z/cIfJKoUJRegqAmk7BdZSl9UpokZ
oo81jpV4zToAX2x1j/StqhKh9FZ9FrNMEoLQVL9f9I+54pXYl3hhNFc+jV86CBDd
jfBdXcA860+9haVTxAsFflpqxXwqg53GtljSkIDolesHrJ8Mem8GdFteFRNu7AaY
AYEtddVFK7tH86Rl16fqGr4FycIvACFavsGAxCji9vpUnI9dgNqjg8om+xVhNOHA
i6Myu9+rm56ewm0gVRyvsc+PrzednshRE4dyxY5R0z4gi+Sbp76YYQDUZcpXnIib
IoJoSx5DkYVYO1Q9cdLStC1D7EPG9TrRxS6G/6mouuUy8pk7jFXHlfVt8W+spynH
o1TEW1siBE1+qKRWkXmLZuKl/Y2sM82AfFF4f8JBL8NhuiMXHRYckpdV8da2ZPI4
+Y2qdmmK8TAfmFBuRyoGRLEiwVdLDs6N6N6//Kz1z3D2fxeCXmPlXxg9JXL/nqcy
iSK83NWkKsdEvKt35ydtunbKC24oyDFVYDW2zdgtCC3DnTm8fcJ95yRFFp7ece/A
ft4DWXUHrimtbwyzqKsJxoMtY9aIX6AUDaegiGepVsGmP3rSYUqjCgA/ZFTVWS4P
n09EunDm/pikbNQG7LbO0i/liAlmURdbB2JbMylv4DxnTID9c3OcAD/OMaulXQ4s
Wbf2ewEIpdE9P9cOKgDF4N50rYZGwQdJN1PwK1i6VKckFNLZnuvMyTddqSbSmnED
MrtaABLbs7r5eC8EDn1qevVjur5S7vcLHAyxhygrz7XDyaVD2xjbjDFKYNdTt7gk
RqQbX2guR3OUpBMo0qD/LTtnrqS6vZsPtM/J4QyC9ijWBiS1q7i+GjsNu6Bp1EKA
BdmFN3itdff18lFsDXniEFVlBzgA4F4dhMxDV1S2blKhlwcE5yb5oon7hVr0OPFd
hkthFNkEQqrOtE7QAbhBbI8/N5OHA/LxCMoTAEN8z58SjC/ht0mlvnhczWkxospf
xFsIlUTdwyjZvrRGaSISzUFm4tmgNHxtGbaSglMeObj/BlcjvfWyYGD5Tyk8ZXFI
teEnhY5b+oCiGgygwdq30amLDkQHUVVp8c/6PFt9/Tx2hIpdbj4S7N/112f2//oP
+yqrmiVY7pP9zlkY1zZVg3TiRTUoCMxCsJbA04NqZZUUD8z72y0aJvQFuwojpIZy
2D7c7/T6wlH2PTtFRJDZre9diaMykm3OY5XHV1BXQZKLWLiVWoF/K//QYfbOJuc7
wDtDYFPM/OqsA2snYVF9gFeuIYDwP8kZYRRWDfxg7e//R83pG1Civ4Pd+AIkk7vS
4KWv9hInz4sZHBMaXgzYY0vhg/x7gjbFi6RXWUMybQFvPWx7qTMcjM77qH6XhYWF
d4roV3I+OYZU/pllesLr7r7fWETUVBZiIqFULXIhNqbpmEz+dpgrXc/+hjFXUjQR
MoNxPMYEc2NjBxUT5VvckgXVMlikxeUMrSwvJ4z+p3gxHTvP4hF17lKS1V4PvNqN
wrO1gALLRLEH1onQO3qJM0tzylAtdoXlTkqooBs9G/bPmrSIEy8XhXKQwnj5sICg
xtLR5rmVv3S68IccE5yh/IOYpMO/aj7gmjD7WC39MRN9UAoWvfvRfZ7dfXPaheyS
I8wH6YwStlfoWc0u9NiMtQbkbziIYA7CdfouSvpkrbwMuKMWuypRxjdFekj/eePr
3o0D90DK5LC9FTY1N9dnZ+K6rHQpUzt7XgusgxZbKbe5s2pvtb/laoZI/x0gGCAu
T2eL6ND4v5AgWzueJd9G4bpoHGQuWDEjoZBtDlA1TB5aIfSYRXCupJU2L0ommn1r
reJvfA7JeNPI2ULL1VMvsyfWrQjBqU3lb/BtAyhNdoH5pP7Tns2RiPNCKiEEblcz
kht5xhL3ynLD3GsIvjjIuQvFXkOGqmMSewui8jyL8FFN2721OYftX7C16IksH6i3
lz8EMd2/SfU1tzyzqHAw1n4Ux/oTzRtJfYeOyw4zKpTqgyJ2gzGqoAtnm/nUw6HM
CqILUQlPJgaFFOkcg64tQLVWHp57thpnAi7PchpzWc9qQr4iOaS4oZe/YZzfNE3+
etjeIthieFgsU0Y/j7DB6Q==
`protect END_PROTECTED
