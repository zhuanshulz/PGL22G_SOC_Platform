`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WY8EEDgxxGEbhWMyXbcRx9Ugy2181c+4mVToPcyellb10I/dtXm5KqfwE94c2DDO
jcamMXdb2aRxbyWDRZa2Pufy7/VOvEHCJfhm6U0LPbj/CkSHz7dTKu2d+kKD9q3z
HHnIz+RoaZeqA8DTzwfLF0nr3kl0Z1VTBwLnBdITJ9+NxYm3o5KVh0R6tghPMuod
kb4NRAuatKIf2DQG/f4fbIfuY0ArvDcJReOveJx1FwT056bUcNj9t8S78VB2luCV
JqNC/9qcD10GQXU2voDqBOBcdFROk/oQpD7AQZwzGCorV0kG4SNbO0GwCh/dLaV8
mNZnJQxrSfoRUWf/UGS4C5QLhPKm00oGVb9TgZQ3jjNpIFeyh1yk7aOxe0q/6Kt5
Vg79qTcNd87XkZH7wnB+jHdabFAfZiX1A02ivEdiRfLAej4VFnW0zjAqtF/VSCzj
nO0dumpJDOUMeTb3lSiwoTnNN61dikz+6Q0hITQNYUO4S5G8gkFhIAeE50iisMbl
qWfQhRuJGn7u5B3WVOh5CGIjdqYUVI6AzwfZM1e3lsBmjcd6ws93gJMYKrKT3uQW
2WGzQ/S7AqDc38VUc2ZaEVL9f5t6Y+ZYSjdx/DjYaIV3i7N44h79lhDBQ09zp7QC
MpKH/bMlT2bZXQR8X+gtmzMXzghwRP65dR34yttDHF9IUMYRT9NtCD25LIcwpJ55
DtLxRMOXD+MyRrbhJpj8N2cuZ1j4/UFJMPXFKIHGnFA+u0o6KUNtn2lJvfuJqvB1
6Va9GMYnSvOPrVX54g8fZp6kl5wrqVqtoWnkTNljwIhWm/PydKcTSRMXnjjK01rr
O1GT97FCY5hNEM9rx9Zc8JlSifQIYOR6l/nwOHpbNRu4K4IlFQXAJhYhcqrrVdvp
TOxw/JkuI3eleZKg+FTq7PNJWZwGTtHCIRwlCyxoitNhhule3SsYm15Yn4qof0Zf
vCLpX2koDG1D6XOYhpKintuDrT+GHCmXdklxF9y9uPnJwHpFeXC9hb+EfMR+Y/BV
AHzbOSmIevBfbxHsvEHnPm5qXXDmsBCP60QwjEZ8/NE=
`protect END_PROTECTED
