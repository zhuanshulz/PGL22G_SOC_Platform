`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h2JF0Wj0k5PYv+pC2aQT8VSG/rUVA9JnCcpWgMc+RAj1GrMDqNiQjEF0r6H5abv+
svqQCzxL+B+IYtfYCo25FKr0reD9tLjJE3Y+rXlwkz2cl7XrwmpUAsUKJbqGGPEu
IX4uYtSqotdAqZF5Ea0dIXUCU/lK+fB7RQv/sEJd9gL5dHv8Lxg1qGlLiS9qfO+u
AMTQZZcyXGQpb8+/igBsb6Nb6z3YZ4l0e8mpO3WTlFJyuIjQY2KXZaMCbHVzg6s2
Ikw8uE371rsdEoF+i8Pz8At1Dj+VGZYAkfYk6M+CB5p884zrAtttP3jctTpGjEtc
Ulch4ymbmCiEezFFdE7qBPHKJmw7FdVjtwf+5kKdB5gQfQXEfeLu2dWiJd6sVThT
2+Xi5ujMOimroYiEmGP1kHcTYFvz4/N9y9pOkh/Yrmdpt1BSYR/qzQ6RQyVx7c6B
z6lKuQClkqFsjmEWj1fEJtQkEN89Q5C+ndduoQM3P7FVmqvM+eE1Mg7o7xBM7Byz
3NYrlFxKFFOuiIQMmktNy7ohu2fNiR8w0L5pp+9Zhq3V5EO4vN/ZigEeRboD5m/+
FnElbcr8lg4dq8CQdF7pxoAOsW7u2HoEPAUYgvP0jl93RQcxm3ynS8Dm4h6auvNZ
8MPaQqiQtintLNjm4DHg2FFZtGJnHFJyL/YaBEr2HpxksVtmx8SaDgy3NrcOlCD7
/lHCZEKP5ALenFP/XTCd1fUtRc/mEuyl+vqOpMDTYmqu2XTIC8qlo1PJr2Wk8HZ9
g2N/E3edMkbosUlKNGjANQtA3OppOwoOacSpBVmwg4XB7lndqRI0hSSDr0XCtBmL
/0BHi6qWZzecoABeZpd8mg8t3xIIR+83AE8pKNzfT9LJ4b+qfHgm7Y+BVYkUX/qe
LWbhLp0o/uR65p8Wbjt1B2GkKfsXMuSt2TefoQ+oNkVALfTwMFwedipsAzZkHtcu
37qcHi8Jf3QmeJ30E8zlox5jASYIXzxgSFCTp7JShSzf/Ry02ca+V3Bx/gKxEGt6
1MYeko642hRhi+q2dx6ees5VvjQqwK6BRxHC3iJPmSiQOSnjHMwykDCXXxSHMvRa
djeiydkpNa57aRf6qN6DvvwUEaOW2msImLsRvZWA1RdXR5JIHabQvnDa0VPEu6b+
voYb1veHN4y+eN4ZQq0YmljcQhUwLDenCVxSagImhncpyOi7CwE7efXzOJ1hOPHD
g1pgSrMI1sptMYJbPdY0GQY/MfVPJf5f0c39UKYxQd8DPyaOPcoGflrap+pztG3t
icVallmQSaB14k2GJX69aSuPV5AZ1PWLN5pTmbuyDDMSOBe3RckpQyN4JArjfDdO
CZwVTEFoQrK0v+V897iUmro0iOuVqhmTf8IE8y2tN1XZaiUkP6sVJ27MVFmsH1h9
muu6PxeGzt37o18XdN6KvDyxp4d2FKsgMOFGW3JyXe+8mRDjoddvn9q4Y1SUlhg0
Jiuv/+0N1e5nifXN72nWBKzRmDb/izKP2h0+LoSVK3wewU0LuLx/A8BSnSR0K/wD
i+NF5dAipmyMgIbXh6QquyeHD4c+wUwz0OAvqEgJKvQGVPqZzvEo6PnyZepPSgr+
IgTgZ2UwLC1trRM7yPBn7O61aM1s9F1ITo1eEQuBPILEFtpzhBUEKwfHibF4S50q
niSy0oOgKI5VaYQnFzEvapHbWxqPMF7Xc4ORuhssuBs=
`protect END_PROTECTED
