`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0Hkxx2sEseQ4heAWD8aEV0zibVyjeMpwEzz+vkmU9nZ2vQR3F70YM9GmVYfhX6lL
giuOZqCwup2SpHK3oUUT0Ve+p7cGli616z8pHF7sWKxa2LZQWmXDr1k4hE+mA22f
LT3tlABb7PyUip13g5WGzSPsdeJqEO9ztWSWN1s02/FAWBiZ9CiRmoQbsQAkehiy
tRyrFOb+ttR798/48CLbfPmRA1NxAYvH4gj7ozn2VtXE4C2Oz0fYDkENAftp9cFn
tKgjabJWuinQy48wDrKBOaQtKrbmSJ6XSBP3AK6EjNNoinzVzoiGdme6oqdtKM9I
mGuotqd9hgo5liP9divloNQIsLcc3jfi0DM4fQrN2QVXqH8ZEE/RUBdtLv1pl+rZ
2CIjgeikTV3WMiu0XeX4+g==
`protect END_PROTECTED
