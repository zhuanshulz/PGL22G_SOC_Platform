`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L6cD8ve2TDbgy3T5vsS7cI7PWEIMJx9E3LvJY5/KHc2sDh//RxVlQ2wUDG9XqPmT
eTwmi299a1HwfhSm1w/0FiTIC8eQAWDTm76EtIUdb+8Eu6Od2W/9dTb+1N0cHqst
BoM+89uXsKbuvAOFnqq8k3azV4rnxco7d3wqSO1mN93WYUizkMsgKw618UBcgFLv
j1xgQc1vkL+UoXtO0jU6CDk44J8OaDQxcfHEoCLrBmITeFxd2+cmH1ByLzMhQ3YM
cPIRDIW1MlBnySdmQO2v1ZpK907qrB+2SGfBG+fZXiWEFsO2+X7rPxR/+9LYvvYr
TPe5ZMGr400s8rFq/QER82cjPw3tWBRdAJfVGCocLWyGbgeeewLMQ8ggvT0y9bwf
pmi5FjTgXgRkl7kSNiApyamIqki+vRf4dqz8CqUKGfEkYC6+4kYAzd7seOIXK9QX
IKUffXtedQGtKvK+Xmgqiw5rwn7UhV/PMP4EkWJC4vjHa6Xety7zUQ7s2DbHtVnD
w3aNnJ23FPC2tyUVrgZ1XWPEM/PLTLTYPttE+QnnJKee9zeQfgZmFiWEgPK/bvaz
/XiotbqYHpQxLNrPBxiTuuGyi1aBDcSgt9lSsS3d/HVjpO7twqbh1jVudsG0q3O+
8qsIGn2OJbuJR97t8YrDN9zflAREOjShd2QFSbQmLOLp9l0Gbehl9ATLnA8IL7Gj
oVvkiOPnvRjohAvun2+ytyn5FfrqRXcAJ8kon6xfnlyUgbwdunLduogjz+8GKZUH
q64eBUBc9yO7biEqclye5lgqyLHxy3eqxJOGettomVSEDnbdQO4KK2++o+px7dRE
Mu77MqzPA3g7CXAJKjLZ8wKzP2D4J7jiNXY7JeUb5TUVudOsC9hK7E63nA+b8bMq
eWErnpi77DCaPcE8nQxh5L0vGP+ywkNJL9NAN9Zd7NmJka1vN3stxXryZFoKiGsa
VkhvIP221vOV7eMPhnb0DFmd9ugfGCTV13JbE/TuE94nVpxhfqri76RJn6bIY85b
uqzXrQ9Py+Nz/Nh0xZVkhZWZ7Vlg6yKLl3e+bkMYBao=
`protect END_PROTECTED
