`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fWfJaT6ZWEKMiAUM6uqlk2rimkdayi86bwOpcEDFGsM4AsUoDKSe3qh8BCOJz6uu
6kIW8QPHINOJHQBX2bq4p7Re4YswG7g157KBZ/3RoZMHhGGhqchRmlVNzYr/mnP4
8Oy5X/gdjK1E2cJaakcOrKvE5XnWHr/BJP3gyb6TgECgX5caZ2ntUC734EE8wXED
m6eArCxfy61PXA7YuSeqKANCZnr/J92gvNq07AdBJ0s0Uae+ljqp5YVljkrdA7zi
gwLNWRT/F3KLcsEAbKt0tUpuIEZgo2lrM2L6AOJWfGuicdUaMePfLhxP1NHPgily
tbZuc2644BkPfYV7iy3wmZsO2mTu1paFGCyGIG9qM71u9sQy+Hnf6Eadgt1PHocG
ntQuK4u1oKAtOOqsur0EvrsYONyo3jHYIP8+XtjGh/hCa3QM0oUUUOLYs8HamcLb
TvdTvQMgh64YjoZ3vUVZeA==
`protect END_PROTECTED
