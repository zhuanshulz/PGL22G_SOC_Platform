`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tNdKdWRy8a0sORvhNfndu1fotIF6NBiJuEk1Kg+KhSP8S2V01DPG61T5Ywb4OIW6
k8ViTdiLiBbNxHGZFk/eWaami/BVt8V65k73PxdXvRSinzAGqMLXeBVLrpxzQpoD
yWqgGbeo077xHEODkV7iyxj6AzU8m3igDyul/PsU7HzZw8KUdB0DeBib3ygOimEn
atkYee0bC2UBkWqbI1HiCPVv12KO0mR2UZtmt7L3kyGcRhG+g0sjY6eMfPJbGOih
ljPgRB+4ybAnWAWFdJ4hbr+2VMphGSBy1Mol2GJLQ6v92VbMZ8trUpFmGAfP9NUr
F7VqTbeOXyS7TQhwbi7HPSRxNxea9LilYUryXkl+hSLLWJAfI59zveEy6XECoy0H
sJfnS0h0kY69ngzWtlDWvg==
`protect END_PROTECTED
