`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lGxZkvXbW4r0Hv7EwjnewcgfFj7WbtHU+SASk94rK2IdlZna6QoaY64YT004eq+D
CMTv7D1hmUIBUNKHmdrCfHxY0PAp0X+l9P67IXVRdKIVGC+aHTv+vIAzfuU2dIWa
3yv3vOAbpot/AoLn5PA+0449OW60HPwW3PtN2fxDeSMawqwHjxbKncnblOnfHkfk
r+LC4p4dJNwg/MNyX+237W0Um5LsOSMRAwL34U5NnFs3BFt/0s/jMfTNWJRxHfsx
P0N9SFZlR02OuGESBb7ZevggLBixBf4obWfAh4Wl4tWKgxsgTBE9/f/XvRA30por
Ufafm3hBH/diLGF0jfvlDN9oqy7dbia0FLsxZ5dXdMcOihcp60T+LH/Mz98biW0K
nS9EIc5fx5doPQP4SdG8gt+rtJqqy1Qr7RxBKC/nWKMabQVF16peBHqMtixXGenW
fTOKvviZrNgsCMVE1uMURBrYn70C+BqCi2hWNm0fPf2u2inPEdhKFjuF08wPpPUV
vz2zFRlHEjXb0jLkeeUKEe84WA3nM0b8VTyU8dHaZPfl5HupLbmBua1IDsI1YXJG
AhGySItZ+/jLitlOoUsJi0YtdfpmOLYttcfSI+sjM+qZtQjncb0N1I/BGXr51lh0
bTWzjsrw55r46EAGYai9vD5Ktz+TAqUetQS+shbIxCnig0jOsCuYM2KeTLh/3skK
w3oOGcll7WX5yIr5F1sUvp3XZmXHe2P+6gSMCc3GLIOyqf/FcBWb9QEJkNONJiU3
0+Jz+DmMxfyGIe5t2GiENqp/Omur2TWtCak4F1CcB1NhWQ8ZPGmUbHOPGM936Lyz
04AHmN2w7YRNJZiD2MEBskVYmGstsJuQ40ZS9W6RVfawutEYrNI0ESQBcLh+F18N
/aowRSSMPU7n49+R1A2YO4Qgx1JTEN3htD9J38rh0ZCxKa9hOralLjoRXuL6LzPv
NuSzj1ew186A5ctfhQXAzKM0lYKyY7h9mDnfOILq4Ydj8dpDxnOR2vqQvBtMW9/b
8KRZBq7sEMYkW5ggaEQ9qUaef/cSFAmwIDl78DCroP0E/tdjqMMYHuXrtFCZfJyz
TafRFX4OKLu8b66Bes3+328XPLXMb04ks3UbTPjLxxpdey+6Y1fyKmQOitdcm5vH
1peHsnsHM9w9Cx3n/ufre8CPBNtvTd7BSIlP4Jz3nqajfJeVDY8EnjF84TzspB3l
dkyoNj+h7RMnNYTGTyScVuIYjBZyBQujD+fXBrd6nTe45WwBI480INzWDwZ3SMKC
`protect END_PROTECTED
