`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7KUHnAYzmEcIwWcPagAIJgph1z+cf0ixAOtjL4PSF2bIc31ASL8vvMq1KkBgq70+
slWsEcf3dKpmls05mpfvgri/LUXOl+5edowyUWAY0hg/kHasSu3hOMQkd0W2i+uK
k3TLvj4QrTvaPS1KYXpmdFt04MZOUOZc/ZI2Tfxd18YlaLgb2ri9JnWqfC5lmRA4
GJaN9HF4MmdKu4JKk4rGS3WYU+5Cz/Cq2pc8EQIyMjcfWzCt6YnfM60h88aeFSaP
Deq7vuRKurtxJtk4NYQTclZ1YdpzF62eW/2H/eWa8YHIl8uOAhrBd9j0QGd8oFHa
z0y7k2FKGPp3wfr4rHelZA==
`protect END_PROTECTED
