`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oG0Vx8MXJzCjeFKpB8v8Ygx9QLrC8F6kta4DfGUDP0jaJ7pagLHT2jH5mcI60iFz
D4LCRliJRrElv3VXso0Geu1JOBP7JsJWBsmLRfp/3OwR2GFrbp1XkPrEhHifAj/6
bEUuzBd+DCfS7OWbz9CiUNxl1yXmvSh2bCkBiNDcI4402B69uJjx8UILFQs4qjqT
BNrHZMHH7xcZbUvdbmSOUjbwEezuon2mnN4CYO+/A6cnBXdCQwzyklrMdnzTf3h7
Hm9kCRrRshC/GlU+K4ymcLMlxcs8IK0DDYlxPNRv+iZDr8l1XpnfCYxs0cUibYOw
flTomfcw4CtllfsOJ91jVHKP9h0oe+jXnTKJhdjgz+1vMsZ0Kcb6F5kUH+K9Dg00
9rUNvR9w700wMIIgbzCsnSpPKgiPLbf820lz26YkVcXAtlhEDokDCl7LzXgfqYxI
uKCIBp+PKEqSZCQcQcfo9mU2DTzTAgtUtOZL+cd0BvQq/EE0OnrI+ztFvyh0c+Ej
WTsbGdetlLUZ5kyYfrlMyM8vrq781F21EIUQ8UGrJJJgFM3z0TzPPPqLG7GmDJbu
LRRFYdgwYswgPVv66MwzgsiBiQBgxfAQ1x9WdgLDRiibmdONtQIw8gZS2MSbMXfv
9UNlXjuembYro4hH47BwQvppXFTrzPtIc7RVP80EErFJylz/uNu0w0Q8iSi/SgYW
R14VplGoiE8Oj1SgRtwtf0zLou4CpjyV+36gKvEdCrSWBN5eF5VmF7UfUeIFZQ7I
KTpHk7PFGfUXkxLXR56IKM2j25ln3zhIkLfml6vn0Vc=
`protect END_PROTECTED
