`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/95mWNN8Glz3zqT/j2ehbBGOXRGWEJcThCsciqniC5xO5piY8E57vgC6gRuLNbA7
G/GkJkqJrx7ZGRljkjSU937yNAeiJm7cU08JQmLzg+R0bkZRximEDZZjUVW+d6qx
4RsypYO8OnGZKpkhw6Colf+mMxrSHbofLWUWCe1jNLPurGUVeG0j9Flb7kswJtTQ
NZO5xroEideUgIbI0+rMsR05WtSe12v+a1b3aExAugyvf1CLiRBt1M8FJs+1kL16
AoYcxWN4K9CbD4MGibilEuNSGEU7hF7Zh9xtZuFQvthVuMs0njRKiyPgIKDP8bIA
o66e6TvvPPjQhdItMNotUiXo9HAjZKNe4EpF7EGWGJelmtlzaeEcW0eXTIvMIyO0
+cxcudYv+XHHJ8CHfZTksqKUOJ3nwwOIZjTiD4XKoFJ7OAhUduiVrdmHFfc1ESDu
DIKutMNYvVVG/0ICsNfXaeQsF8q6rWr2KtX5SuOZmINuph3rOMti241Bo7FaUPiq
1RDYzjZdRyTWdjR2wGIyftASg2y3+LhP+84TqQL1i2UCEIrty03oaAPOfKdojpZA
146CCQzs/bz8mBEx6ezPNDWDNrAW1anvtVD2mNrrFwKXFDkhUfAiWp0/UME+jEHc
qS40PT3vkzl3tvi20Q7Dt7p6FTb0ocYY1xb3aV6kqaBawO5QaPC6le8EAjjyEaz0
u6rNVRe6gVxbqmPcmL1MfBbYUoD6l4EGiu/zTh8ZL4BRNRoRgDEyNTD+fn3gYjEc
DbNUYOiGU+aCSqq2TkYoWpVUEapv7u8QkTDg8hGePso3wrDQLL9bChhnFddB/4pF
Y3YC2SZ4f+TQ74YStKzn+B+X37WUeqMenU+L6QoRA2SBuG4VfcngOxfiDNk+2kyO
oz98WgTJVbBFfK2eMX450wcR7oAYg2/WXFRjonPRuh7l9mbg3kJ4z7FA+76bjfSY
a81Sh1BgkZR8IgjZ1j3s7fh5RiVtr8k1axcdX9v1o//I8Nc47S3yt9kzweYfL+BT
ZfQjveUYoTEpokyyfu1V5GvfWun3fwV8RGb/d+bUO+h1v77jgDUegyKp70JePcp7
pSEdLv/nDdX1Tb67rRpBQSIxsxSY/kno0vTBzeKe6/Vv0SWL0e9lTKdBQAXjCRVJ
MBzx3tEpK0HBvtnwOjLM31V6mePw/Qw/ovyCH61z/BRBUCmwVSIbP6qDAzId3Pxq
qrkWm4bkRblswaLV0ckELDc1LdztFjWbN5o8+c6SRwDbrmE1APlFPteThl7VlQWr
iyCgfoU46CeRo7XfOjxB0ACrqYD/2udeathyOZOeFw0yXwbo2hYCXG+OaOBFf+zz
HZFHYM2irRQ2gz26++kpz0T2HF+LohjGKtPfng0bfjTwH+rKgESeqEWHcogl2A82
vVTv3cEmEevvAWy+BXNMjW6TcS7SBvK+fMo66nYYHF5P29a6NRTFEWMxgOLt662J
w8N9/6+XXQANQquhcC3faePEthBxcT9n9/pkcThas1TsY2VLaXjFiD/x/b0ta7bL
GkwE3zH5ol45s+A58zKmpLux+MHxcKWxdvPIAHQ5ELMHzXaUGoKPdFT7g/PI59sk
W36h8ZhfsTYaRep1BO4FjnjlsPetyInFAwhRa7ksNWQpSWu0gCrAFj9r1lPR8wqs
lulq6ZnTy7gQaDGrvr7lscIdBc8scML7oFcsi9/GdSkjTNUlglLT2hZxASqpYFxI
yDY8cRxwtQFb6y826c3vPyW03GhjkhKYFTf5uxEarE6P5wzhJ+XzILMYS0v3C68o
WtKsR2xLJwAI/lHGvVnTYchtR2zoWgu/cmjTQu1CuriyK176s3kyc8oRL35YH+R7
te6QZZS2nWIp+LlQkZUyHDhhUa3M0im6gP0mGRkedqsMKvL/RwPzmWeYHmgN2+s6
c93WhC3I1s3k4kdHWCtckQCnLSUe6/5c/3qWIgcyFsw=
`protect END_PROTECTED
