`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
moIpMDjNYhEyucnjYSpaP9lkAn3t0LLQizaRWnpgfaQ1jpKbIhjJCODs8pYAyIbz
ykacIA2gcGDfgMhYljVvdxhQ2s9e9ERaxTcPoL7N+yfHbl2KoaEhaSCY5s5usa0I
EnYiMO589JTVigt8hmwY9lbu7WWhjKGJFzPEwVJtshnhLZyNOdvlz4wa0Z208DeJ
e33YXatAHk+pI9yNYZa4DrSs3qPE9sQr98ftYo3j9HsHoVEmjrp9Zqo+oAoVdLrP
FdKczR4sbh7Nps94zElRFMxWxoXTZzY6fbbHWN+WCjTgkfGzS7gsb35epC2341r7
eiRwA1USSBfq+yMNSsKibaxgfb1mBOeEKLRj5TLVdGLkRaztrFxJTGr4jZ7d/mRc
E5btIXvzqsc+95jaX/DajjlfqlV2yBaMY4VDjtqEQyH1QbrSaazBoptOttOCB4px
xaOVNOKHZMOxJkrqyZ2xI0GXt9MXSmPbmYR/61y6LZS3Nuy4fUUNLMfcg4HN4Zrq
nitb04ruMtDl7hMJ0+gJYGs3GOHlURXbMDAUU4fj7eLhsyVJ2psEvN7aAGQmgBa6
zOF574SyiIR0vvYo15k5es5s0OqHijzvfyXh67RC/D2v2YokDWsqrnLBo2/ERn24
aSuzDdQRlgeT5aT76UCQH4mR0+VQtpKxsKXg/Kh1Ck28h6if4MahS09dOTgfzK7e
QPYY7j5oiZKX6FMllHni8Yd+vi45uEoVpsSPG4iJY1DJlKGyWtkzX6UpbNlqX3SQ
2PIuYqtJJTvchzjOSs+VC5jJjQZOoHq81yB7mD7p+7alAdSpffyIKpJMhciQRNwm
z/VAAjlGdDwK3RhBX+olH2O15Biz6dJfW81DMfk7NcG5GW0MhbDgzYdpHjCbmM54
TmPdvVKO1orcpi70vNwLRcNE/c5R4jCiFq85xskfazpr7So9RwrOXFxsQSw16zOq
M1KTtEV+v/Q7VdcoC/CFWj21j1UOQ+4Qpvhhbldpm+jeiXPFn+wiQkYGB+eOmFnU
J4leekfnULc5Cz7HYoJjmHubWrnuMsMSB8SkuskNOEbZynnEdBaqSeTt8ZiP2QPo
/xF0YH5cwJzq/cMhSGneF5BOsirKdxWFKT3ZkLsehIXILUxRdu0yRStfqrn5xuEL
sp0/IH4pqFJwKUigP3a0TZckhWQqyMTGjdYWCHt6sja0ceyrnLYXeN3Auz7evgUd
iYgUx5914GDD0OBqdXEoZDeXYq9JLG12OvL8L8HTNVHEZsgzgQDSCZ6dwYmFdN4h
zfcPlwwBSMR7oiPJxLOpwd+BuRzY8IwpUepOKR4xNOPyC11XichieRw0SS125uMl
mgUP+Q9ff6QYkjtAasnM0pzZntioc7BfUnKdGZ6XEabQqu6DOuavKl0jWs8V/3Ta
IgMEEZj6BklyEiGAhWCttbBb9cqINhtFW7jYnvvqka2uODSyFaNm9rwzRX8fU0Op
a+adA/ThQTGbg26b9aSUHxlLBeB28Ix+lclu8e2YK3+2nICINBcWhUpxwdMCHxCi
2mbQROYaVMR/7C9XfelB+oYmQSa7jzPU896k8Gke3XCkL2yX+CeLuuMfPXmdvEwP
gVdnuMQiP95hYWbAg6vQWe6hm1bsQLm1YaMu129B8YuT3teF+8i8czgBOSq2Hsju
Cuke3WAYe9YrNrCZ0ZHcywckGjxaMmQweewNQ6TNZ4WdU/S3ZbHV7V0QMiOFRC/a
eRmcy8PZepOR19xbZwKzjFn2bBjAlGEVyujY+N5YesNObOdB/llS/G8070zQ/Q13
kJXZCnAib9NHgSwJNuGTsPT7Uz8uYBRJdbf6GpsLJcv1fMgx91ThEzhSkgehjHhd
05THGHJ2aTet7CkegZz2LIQaSznEUzIzV3KxTQS+iRjBpM671WUlt+qet7cwILw5
puFWeRpW56kPmbEYN8ROqNlnFBfcMfPNk+LshxhakVsEBItWiPyDnFC0woV/cBGy
Uoc3XhhSUV2PgiDzFaXXZOoNgzty2PQY+mGoOLSZfi+D0IYqId9o4+OIaKfpbseW
/Dbr9jKG3NW7Zxepm0WbiyN/noRYtNJXI8eXCAvsLsefZNCaOuu14AuIxtHiIWPT
8EOJx50ZAzFtRrYx4ARS2If0dvspex4tfGXhD5C0etfnxqYGYT271YzZDXXOC8Bz
L6A7aaOGQSYlPYG+7ZoWhLnChvTeu6txYHp0ZhhkFF8xaEXDMbi+5j2TOe9IFpUc
LjPpfcO0rqCU233r9qTOrTr8UNc3cc+8U6RyrxDHC3c=
`protect END_PROTECTED
