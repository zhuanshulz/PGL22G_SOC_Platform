`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5MMn49Q4W+iTjmXDXTpBgdYpBolAE9YiRe+MjAK3nQbsfE7bfBNtq8xq4U3eBwhN
19FbtBtNXzrhfUCbpqokR+dMjBInxjaIro3SeUbwQHIuXYjA33OT9Nx1IeLSbj2l
GxlQ7EDaWq6gB03WhLW6WbvaTkEJwSR28ch8NqZ/11CsW/vq8pKVJEOx7BwTbIpY
exxWZiUpl8hQRW1YRzYf0a/OXcoNcTIV1gcTE8tx3hDJdvvznt5nCd8GxwdI4M6M
9wO2j8DAAmIBnu9s+q/xcPAOT6esRas+HkfS3ycpLDKTyu5gvvw8U9Q3cKyFiIQm
XbqQjS6Ld7bxpMChwk3+Ltm7LSCMExATBVmBmxPd4FbFX4wjUQ0eYrNw3MHJkrYw
5y2cHbSF4rb5M+BJ8ApTH6ziKBQ0gk5C+drlt/fnZPz1KgDOkB27mFpEk5TznO7J
/MNsRrT97glMhLelrOa9QZDMrCX3ReiR2LOr1mkgJ+uFV1O7l/k7Aog+2aHTrgXP
P87hf8BzafFFDx8nCsdAFxR4WQkEbO5jvBRthxAajHV+NU0wGNsSkuIunhM0W8Ic
rkJyo+UHe9rg0tLzVjCtXBzDd/vjxFlgknl/hex8g/46q4GfpZYIs2RyCL6OFmjg
V+PIFk4vN2MSY7R4cDnOHRBQbu1SjuNEWQtIgGrDhan9mGMK7/rAraM7H+czBnI2
QeUeUnxv4lrD4pCSr8r+wDvN8ohKAIEc0i1W84RVyAG5gsDVuXrY1pZ3/xwsBL9j
qyaCy3xbG+FavYmGAksCFnKkkigCusR5zjNLlbvsfcAhMH2wWw6JFzZZD8wXAZqL
HmRyZRP7x5xFmKo3rDZ4ffPde23d6IWWE81T7e+c4m5Y2jvODxkOaXqRuNj4FmLV
1w13c923OWWXXPYyzk0Oz2aE6Ldnl7ybKNqW+EHqlzgANkYzDe31OheelVLyduH2
igLFmsVTHEOa+DaD/SGJRmmdGn1/BEMmVweFH/6Rje+boTFwry34+dHXDn3r2iWH
BQYja7vG/wvPM6yQ5ldgV6NF/DVCKPv26ltRVI1enVbHtXuax+7LPJZZyymhHpiW
Ch/ZG5JDfcFeZthjDTrj8T6D/V4fj1I8FhPjV1l0OpXmz64qLskoGgvqzxj61Itl
89KBDR7X0TUDXOAqhG1qCdZOM6HfgLciasORnlpFIzi+bRb2MRgtXD57xjWXnYGm
yjiE1pEgQV6ZmBD7G33e4FZVEBZOCfHQp936JyX23zFZ6aukTF99fNBlV5jvttu0
evslLDcK7y3P594nl0c+0jPR5tQl9Jp783h6vdKRElDbXhmMz36SrAZ5lnb33mkC
rkl25ljOMkz+NgRYHMndmaXQqbBKG7RPhh+r9+f7g89n0Ll6aCyC40QczqTLhyZ0
mqYSWOHDmYxHPwSoDe1bu59ubuDBwq4XvsazQFXxNGPJAnNNqXpEKV4bPHQXFkhJ
lJ4DrkITwS3hCFEhl3FcXVUq78xRlXeIz3iNHHNMIIaADVrSgtH6ibScCds94txK
hPUsN4KqinoPHucXvpbPXmn2JWzrcXwR6y65aPZLz4zOpg3l1VyqjEAoAj5h9TFd
n0uRfAsbiYperks+enXuOBfua2C9DCUTCGrVs5d6Xp5Hpflcz+BBOawSPJ4HyVaj
MhpiWQu0CDAlYYdOaTq3WpyixXjmuYhiAuO/GxNKqzp7HjaSuDcegg9uus2b8VFJ
Kw3uUSZfArID32B3Y59P4Nji/gN5HNBqPf7xT7tpuJirtf4KxZPP+Gc555QqO7B+
p84WxaeS4MQ/b/DsN052S46TUq6vf80vp+Q9qOnzGwmTxXD1GogiglJOdXA7vZpv
igQoDH1zkJ7IZrav5M/yYEEW96mMssCNh/CC8b4oHiKgdrGhdhBXYn26Xi4pvAPr
YsDnQ5pRjZ1xym1fphA37lxXNcm/lAd9YPbZeQmx4z0cJ4yKve+kLoVmvQku6EV8
zLGxwTQgIPBP5Un6pQVT2XimDxE4abGVZKtAFg/U/y7JL84ZF7gbe+L9ZCIdWOSP
VqIut1sA37B70H8QpeBzihvdSqofrCvuAksdt6jkcjhzig69BHZdmfP1KTBnn7mI
Ip0qK8FsZdyFP/faIaGr6ajdWG+BccXIs6aV4jUB3XWebbdK3krKRt7O09UDfu0h
MAcynyYtuElnycHwI+m9tlrvbd8d1ZkJNwqBpX0wZOUUPeJCPAm5lSgdEte92pDn
g67Vu738YZSRXkM/nfcYforlNp85iDi5RDIqo2Uc3mXhW1diUWUIekCW1lYqAsu5
PhB09A1kL9+/SNmm2CklQI5XkG2qEWj1gaTEejacFYYrbvPTR/kxVBnaAQGsKvDb
+giLco0SaqqyRWDQ982YykzBozdywe/FMKWY2uLS/EOpdJDEcKFE1Uq8EM/ozCQN
zw9wthTGIHL5Yq9F8SLUQdX6X5gucoMOU6xNa508dv1m/OX4oqj4U2+Vy+hidF56
iXCcTqSFvsEE7A6r3Ml/FWxIemz4Qi++s24XMDRs+vrYIt1Gx+X4QNImVwdli7Vd
dm40oRwYkYGS9OQXmsNXKEIkbiy1/QVnDrd4v10Jjzw7edCLBK0JX1AIEpHgFk69
iW3KqZ9kYIB/YEV8WKqYuUh5HBg0+PO8b84GEKTdgQPXPnBWNtpEUXU6h5D6O265
/qKEmhKlO68M1f3C2fer8+j97Xap91so14t7h3qxtWjXvOhbybNHzWCJ00aH7dEP
AK0dqG0leGICWbO1Q2OLHVuwwWR6b26nPHjtyP9ikDBQrLFtvr2wqvmHTwweemkP
vOww331qEPb66G3E3MM/3CHU5tDVQ2355XXeXP9WKjUkGWYHf7nZ8GhbTxmn4KJT
FAUG7TuZRA57iIBo2ZRvc9gXQO5Nu3Rn79Hd4GZYQrUhWOYawSQSzU7kd3OEAsdJ
0cYG4yDXj1V7uwGrWFDs0BWOxngVyd50XLgg6f4DaGSpoIyADNEAq2wgiix18yLK
NDVbZyDj81CGTeu7ldNp4DfI+PRoE1gtBprtEX/+r9Cnfcfo84TzDUP9s9AIBd7M
BPSyeLTqSJgTXBqb9yEGIaYIZ8NHURkANEv9aeh/NkH4CwBR7SO/Y7ZpO3chGM2k
SPp2jJZ602MkIIXP0WoWG0L1KPEuUpTm0UF/ZpJ/MCeiJgsRQQIX5aUNwm4I77oV
lyEc8KqTrSmdA7IQQCtLRnMCU4ghA9hMgVm9h5FGVLOq1y3725s3WZuQBzK++FPX
B4Sjo5uBedorccfychSk2vSkq/T+mpB0Y0FuxgZzkdsjEdW5cYT/Jm7+5pCGFNk6
YOTKKyVg83FegeSbxMHN455zxNrEZ9v6/S7QAWlMLW5A8Pgqru8oY/Mzb2ZuD271
Y9w/k9m+Dty8Np1mkJ2gv59d3gJ17HlpOb3/iJHdKX99rgmwirG0Winfk36eZX5Q
RVdNhzzP7HUiC1b04v6cJhP6i+wOLgFKgXahsGWQJcH8AZAnHyjLwNBij0bfs+df
xR/v0W8n+BuQJZFOX3sjHQhTdu+FtxdqsvFvDF8A304tZpkCCtulEqqcWN448prH
q+JwpusSVUvvMF8bcg8rVeuww65DiGHrswwu9BMjtInyg7zolNZtbmMUUjgKcSpZ
GxPmOwDs35ry7JLIP8FO06IhedzOvEw0LIoGa2imWCtXdhCB2FlYren9Y/VIvfwB
XvFCSXLwbmnQCludtFSsEfSTGOTklK/vkA5usRY9wrNuZ4C492wBUg3h1wuSD/LC
9vuUq3Z27i1CB7yxZmKZ7jfhOKBMqNpjqLzcdgrE8ALnoPvksYK/UQ9o3yv+qZ2p
kzpB1CsFNYJ7l30sM8dEIpwLcGdZTWvCXl3uKeHPf9tu8lCC0NltYtmY7GvZFMzC
BES41qjL+jiFTWHj9LxAzhxoHoTy/ouoKfzuTJkWNjyZLkpDnUf4Em7lsBrdD8Kj
gfuT4SggT9Y9ZKea8+zFHnno+NWyLuRsFEOTmb+BDSaboStcS1qd7nrdLZy9lxLb
B2CtQcBG9w63x4XwYRliu+kv09sjgdO4lXQ3GX6DCl3jibRbyxsqqXftJMCx1URU
YCSv4rY4ofgh0O4AZj2xCgmt3co2yui2EyJ+OtICu706fgOoTVTv6M3hsPtVLM3t
Cqr2pQsXoQF74fbcyGp4nwSx1D8Y1WKq6+WiuzKfakAYbZx0QxpO56r86ucg4c2x
v+WigqkOPA03kD9x+whh13V9x1ZS50+5/lc64o1Qqy63gQl49To7svugTQdItzEL
oVu5NHP2WiG34GeLHGFB/IfJ50eSz193D1f/Nm80FL+4FlTmeDRF0qcoeRWJH56T
7SVOSOwOH9ulX/vdA6Gt2Dj8BpA2frSZRmPWP6MuHSVa/41gSVtp1sbBByLpdP9n
KXxlM5O5A3LLP+8/tZLi7a7jhOTcxi5i+c72PXC3IdlP8ZrgN1ji7FtZfjDw21E7
M77+eihfFGkW6dbbtgoWFcgyNU1R4i7scRMbpKvoQvL/M2T4X4kaQn5ydaU5wZVw
zV2zV3FxO5mL77mlZ8Q5oo7UR8Frg9UEYVtaBKNyI8T92N+z52GchCjAukb0/OYS
vMquZHyOf9VlfMbzvv/dseF++Xd8z746HcFIOtbv8pVmB0Madv3gGAl9mnCjfpcL
w50gBHMce59vratPY5ELuc5Ohn+EmAocKSYNKP5JJ65HP5Pkmx3toY0lth2l+dZv
LbXMJmWHyz/gVdayV92l5j2vjnLgYRrCPLNqD4eZVHVnf/FgMsk5MWKttS36KoQm
9YoUvkJUXUGUTMZRqYkmPmV3hFIISImsELsLE9+w8VJ/KSPkYIdFSU20Rf7uFRH1
x+sZwAfoF4E+BAPGpdx7exdLBCoAGBj3JOFaY0FrHSNP6wLW8oZqoN1Ui2SGEoVx
3AhRzSRCsaOO60eFOfeOSfmK7TGzhpo+v2YRmXb+2K+wz3243LzYTrfhLNJw7my/
vM0gYjeH1iVCwyM7OxLNLET2xNQEoKvMQyldHcLMfMwYyW9i0w9BFVLAFz384tMc
jQKLw9fZJnmTLS6SZKr4J1ZA/7XSBRSLxZKcdMvcD6rWvSWBt25mJ6DLsuMqPRnt
bEomMREv+7o9PVyeE2VK22uucj+1KlBen6nZdb0gLBN0JQ0LdsKEcfxGOJuv13Ge
uKE2V71WZjiLnw111qzK7kdMzXv1d5milmzvd3x+9PipGSMKDwXUIvxgfH+LleqH
DDHareQQ67Zu+47UUAh1xfnEd7XK0/i7ij22ujNmI16vg/8RZAB/Ia/0l8CerR/O
ljCv8KX+8P/oWwa5rxW5qXUx3NvwIQcJXHuAebRUjJlpLma+Ybvr/bidCveZG5c0
XsJEgUx6VhOVgQQX7JRkhokFTRh/FR/KIu1vLfovcP9NbKcbPwnj2Il9FkruftbN
0ffelCGbygXt5kxB1J/paqnxl55vqKSyPk0BmrtaP6TJEbwmoT942JiLNU6EOCR8
/vwGc48CHNra9oTeBWPHToG5HXoVOvLnpwJUXdfbbl/9yGv9MQZXM1cL1bnzkrXR
eABvxgeEdGLPwYgwXZq+Z6h/ndTU1WI77tpUXmQ8ilRtqi1DDsmxlGoYc8trh2r4
8Z5D2G5wV/ugv5k7UnkvDKJqhmU+P/Te182uRRysFvnggrVoJewMa/a8TcN7ilMV
oSvIXRxz0LmwpFjherc7sls8IUbFgSgDgRUg7mB4TK8UzlpzojMcf4Tsgy6Ru3bS
0Q+VDLk+mrCZbfVkCNB4yRZhBla3ybZsNGus5PJmT0aXenRFCyp72D1SpGDrMN90
+yLDFiFvc/VGh+m7E4kKCJ5x2ylbBBYWl79DMVuIYUmtfPE5u1mdYNZ4+PFeUqee
xsIqU/jwO9RwAQaT/j4VvZqHOMDOb/T0GK5H4nrW7Ulvr3wYAj2Uh9cvL3ixTYRC
0jGcVcpEfcjbCfzksNarCCuZNI7i1nYiqKR6YilJvpMYr7xWulHg7IlwxK8mSG1i
uMEdnpRoRLYrZNP5pYh1Pz0MJmyYdvtGL3qmkllOkc1nB88bRYE+52rk8Y1FfOwS
J2OrCAu8fGj1fgktc3BHQKUymr4obajeSJHdDc5ZRhAG0xfyaYbJoVBwyARgMdQ4
6Y/CQKrhBjydmp79U002XAzqW/pzlyHbFwWOcIdiTX1qBW+LtB6DoM1G+AMRKu4e
Ncx+QsNJAm2ACpgEu1vgd+bqVNj2coG4kGJzdfh3Fpplj6+m4Uvrh4fBOz74YGqB
fR3/A8j1tyIUcPU31aoSubfWDwA0K8eGhev0jLLq+4GQCPBfnW/nvc+NLOX5mojv
BNgoTGrMcCNc+VONN5jxolI6+mryfPM5y5q4BZG0UM7vOJuA6+JoXkrxCwc+gY2H
KyQkGd/QcDvV9LhaOtiTBxQ4/CW6D4YlEcb7bmcsquQ+oayZavFH7mFeLRs3h4Vi
FSMmFyziz5QMb9GF1jkGdTp20mqAgRGKNzaBTJas3b/CdmW36azuie1VkEbe3/Dv
P2OK8K0GlBCNgBLQcjM6Qhn1bCJcS7jNWOOgMeKHRJJm6IfbSKACf1QJTtXDsUZt
MiTzYUc2pJLwlLrhSKlfnYEkkE318JU2yBfTQvWtltLCfS7IeFhqPfEU9t/f+p7X
SqhXYGaiGbFcY4uVCPiS/y0WjJlKc5v4fzglvboRtXifWzqJsIQkfAKiJ90u0bFN
I1PIuuS6/9DdE03vKiOzSUkAdr8LVQyyU9kElkSbZZNSJRpWIHOhBKNmJElzkkld
C1BFbG/eanlG69QAg9l6JOQlnTLeHASdXwzOi3XneKf2dXUuATVozg44YVL2i2uv
7nQHkicJsKJc6yGF18WIdCPPwTsFBlGMx/ACmRAr+w2aKSTDsFiB8b2Nhh4W+ehv
w83UTerkwQ2znSOWXsVT8KGP6o/9WADpqVlad/bnH5ppZUTfw+gam1O+sw55kBai
XHw/+S3+NbR2QzF+rQNpOTA71YLXiEWkwwW3ZylRgaxsJKE2cojFh3Mz9IhSmWyV
r4tug2HVLVMLsVk9RYiOT10OjQLY3KCXtVxiKUAPzrhH8TJ9Ox0GJ+74KbMCnOdV
zgwhlDwQrFJPaJtG2PERrcGbrepZmKfzd5jYyqUpxfPwm+dRxVQV0NC6EYXIeSC6
Jcw6AZhcOBrlpvt6XqipfGS8CtN6YUfodQeYgTMPuUuisvZz6hqnCyZXNTnMltEJ
ZdGM5IZ4nF5LRxxPxGiZwTeQufbGmcRvnbcZOxxgWg3yG3aSFcJFh+JDhnl+0IxW
S54ANxR4d6SvxBKsZWOjxm1Gmo9V/cGUweu1yVnRNCYQ24KrEDOH2ov0/HleMjg+
d/xPcSrSXVmM0vW3YNCJXogDuFU9t5BDP7giRsrxVzZPY4cCMYX1SqLSwUlAkJXR
E0RXAt4PTCUZzLATkwpkfe/qup9RqGquImwJttQilgpWFbz3QwTOvk74T+bQHLXM
2ANkFDZ1gWW3FUnydyarCQPQpGcRjYuWkRgdQBDCxDuPQUNcRdRgcfuiymWEM532
4BChdC101TalORIy6qShFArJUD/QzeEfFDv0m6HyD9nPCBkCoSGRhWuJkrbfMgYW
4HZtWcRY4q4Ky+km3KR2FPRPBTSzNZwq3pc0FghMzKVMU5lBT4xaLNhrDURi8mYI
34cSAO053UKuREW0UEJY9+yiFqwGSKUdUzCCA/6ya2P4IGHCgCmznev8oo50nzq4
TU3zs4v3g7bO13HvcypzFosD0sma9bytVSVw5qy+ro4thcPhyenRRC9DklQc8Rey
H9kYDNodj3cHI6H8EBNtXSWGO+7l42x2d91kbTX18IWwl1v80rnNwZJcD6GzxMci
69M87JjC22H+51zAgmkI52WGWglq5L4m/EFVXVGDKb5ICTrogniRgV5+L2FnPiy1
bsXHnP8g+q6szsp5CAMdRMtRmtBD2NYRmLBuMPTrNWtrFSy2jWM6cgJrscp/Y7ry
GWaSNezm2sVkLTc1TZmop1SGSY8W3MM2vp00PlASa2H1h1yIKleIqhmVrolrRvbU
MOKEmNJsdrZx9JeKNuFnk5ULp89Vp6gYlJhjPx6BTl/1uv/pwLQgO8gwBf44oLng
FyguURH0Q2Ens4S7O1IeWilPf4QFahLVO04wEw4w9Rjpyns+L9Mvqz9KgrnqRfW/
4tyJv1RUgryoUN68N8amcVppOUMBZFjq/0pJJzUiBfR3c0ehG7rII8VbC6fIqS6D
IhyNe6ABbre6DHwIlfVZ5P+W1QblNF8GBq58QLG1ZoHw6aLLXqfEr9bHbMoMQ3fs
BGK4dewSOPbpmrAwHj9qGy8VdIryNJJ30QY2V+CtVZ4HQ2RZo7xO6J0SjcL7X3iY
BNxsWHL56cYIYokZe2dUCg6yk3e2pSLgLeI6o8bmtHlyKGYvoFvo0JuvtoaEhi79
ga24NOzyqSpAbZv7YwnLQhJ4TPg6ugACHZdsNJPTWL2Ui+aTGImpKc70f9eh9kzD
U0hbM306iz4+0CnQeR7+uXSklZlJjf1hZkyq2ykjnfyxm4xN6hbjjiJnnr9tOS70
B9d4wVTIKpb5aPLiHJlqoa+j3dMuT+lSvGK7xLxPAZW4p8CycruIrBD3ccGhhLBI
beZMhUGFRhunKSyvIjTu21+H3DQE9RKk0ZBjYBcAdTO60cBL6fyalaSJZ9uQSfQM
D/sh6q1WHJCt+YmY+3nn/CoOm2+NCrt1DD95caeP4DVQQ7dM8Uz3GslKLqw4r8XC
i0/NJjCgGsDZbUT0SiWom7NfveHbhZqK78ki862WlBvXJ74PSzk0ZT6xJQDkObD2
/5TNpEgdiuicdPWe94rDy/QRxrdoUiCj9niGwcF9L+0Wyvy8CxDYXQHjzHegswv3
+ZfwNT+h6scpKgP/73M0xxR/UPHvQVW9gvtloRODlPrMTEqVN61IvWOjhEOit6Xg
oLlq5LV6FNF2NfZJCkWNsIA3f6q/LZhRc6iqHLUiMcQ5Qc27L5gnv48Inz8OyISV
f6PyBRslZr82GYhTZiAWxHtxwDhcTQ00nvHQFvMXxVdeeh9sDOXBgfIpXMuJR3AP
9tcmrrBFUXDt8ZL0zxJQJBp77qrtmcCt1tE2CcHxc/EiInO7npNVJFzNBPCVMMjN
5MUWdni7JHWap9hcCmJ9SpsIdQ/zOTF6b7uQViD06FzfGJ1k8Mf6k41fmSsMKr5r
55pd7VVhEGaqr67Cu5TWSqMfW+uBhDViAi3N1qpp6asiKg29XJqdo4y8of1Td9ZP
vW6ByAyKgsCI+cqNJiTy81Z5BncgFCubOz6lY6HYlh6e6dZoIrNt9ErO8Q3C4++d
WS7bqbmGVHWouxCwxr38K/irG+Obfvf9Vn6AIc3S1DZBEYINza9CiBdlUWvgGySn
QCR7amqGo5t0aoV3aEUBBm4L3qGPFAryRojjNxLBH7pzK+kf099rsB4TLrmdcTnN
HuV+NBkeMS1X2SRybT6m5v024M8UuMUJirNVnp+nz4qBaadUbtE1zVGdte4t3kNf
kyUK66kVIjWf+TfcSPN636Iw1M0xsxk7wBeVOwN1Yw5XZj8lGqgQ0Ro8O56Ejr2i
k12HICIGeFsMTMPFVbTcOd6TLYyJZKcVQV/K5veYN1VZOuh6LZRor9n50dNbE1zy
bmryO/nEhUDmS1BKqvMyL8OzZr/6lGpeQf7ROOQ4udPIyXOzzd6GUH/QCM9Ww0AJ
aCaWnDPSBsl5AmGwrmrCoeNAWA3Vs5aO+0LsMBgYl06YpLWXiqWqZ0X2AGdrIuul
ksxQFZuixlVxdKHNtnEWuYjVvA+s/8hqLYbAAmvEJC8+/K42q2t/e0dOWhSaWjpv
vbj+rY3hSWCQMZS2TXZcfSX24HSnuT0SrWlHCd8CASdOO4jQXhSjF7tqP61QP1PV
a3EElnEDt8kCd+CJw8uoUYBECel7quaGYrSUFm1jj/MEDX5oDdNUSYvbXn1vCVP1
78dh9wkWYgGU73oFZdaQSTwFpilWRNdj2iNHt1geo1Q43N3tXw64P3EX9INee+R1
gzjylKoRjRl3PAno2Uo8YsN7OofDdVwJditWuwlkbFqGASNIm4NqR0tT6Duz86xd
oNwBGIi2cq6E2j0PcqkXfQ7ry3HtzAk4rQHV+NVBf37g8UAgFK1axVZ1x0biKFfq
Kd7Zy2NAopHC55eFjRKBMOP0MihqSDxDTyRh1JBiS2Fi9OQNZsEmb/uqupX8XtiW
JWBgGrZQab/zIBhL5WIx5uVhq2GMeObTTB+ztgBqYXibsoeNV83M6Ub82lDdokof
ZZTTgWGU2HjDScbXxRn1TNw2fB18j1I0SdjzUiJUM5wHjFEdVHB62lO4b/RcWOIF
+zjeEjnd58Gjbtd3D6m5S1KAuWvUnZZ1VlvXcOzo3sjtbIlCmqxIUh71/fS2Qla/
0z2LKJojbbfq78rpCPDUc1Ugbz2/3LCYw3XDaQRW6PE5MOqUyw5bKqlElp/Wao1B
FybXdYoGHjKsYrVUlT8XyygT89jEr+zf8xTx0ST3ia6M6R9G2pvqloUDMqAju1vI
ZGB2F0ZvfYZ9nNpqE9BNzGqGtOCRvMYQgzgGjWMFWOzP6FGQNCHuldDpUzkxf0KS
TRGAYkcYhUd1h5KDKBv+U9NVTsRuXpogOl5GZMbjoSHrs9YUBXtfxEx+KlRXykd3
QJLI5Tz8ZHWTzwGaIWVuNlcdtNTyTSX1fjWAOuKkabrzNcNRSAugx3vEjA+3uIs1
4lt9d0FoFrpo6WQ2NWOfmlGUJckRQof6bnV5qxt4VMnXa7MSXCGAwxYsOCZMMCmY
T5t3fzqy9vjESuIZpgGoP4LkfZQ26ROo5QeLGLZfLuRDPB5m0fNfqxWTxUIJ5HV3
LyWrmJIWAx3rK/E4H9Zg5og1jTHk7Llk9LUvtFswhd1BlHPGyS/RzV8Xg6H/3azT
XJyf9q14xAyvofnNmuX9ipmbGsV6rsAI8pKBAGXw4Ey9uRg1cZ3UAJYXhypLWg5G
MVZaxYgbzEOOKhdUeV5/j1cETncI1KVu3DYJsRg641i1GweRhECGVtkP+VAtc303
tbUnAZ6l21IHroIAYCS+vYm2TAVFu9ZDUY3ahuh2ZW6B7/ogsY7+dF0l1B7z+xf/
68j+a5dUgpJj4VE6eu7N2X2ZFU7kcjTAcS5ApszZJXXH2BdEUCkHoNlIssFuqYEY
zq8TQOBjZJtwd7i3JTsp0tIbFtvDd/YJ0JoO6j9xp7D3DeArnC4ozxBJ5jlcLfQT
MnZ9+rF1GS78Qv9/jknlQ0CUHySIcCmYNQbbvszgkhv7ep/LDJdRk4vHIvS2PvGR
xk3nkTxtYOvFmiGdxlw+xWsPEjXoeyQcFUgto5TmXv5BuWZVAr36HACtQAW7OX+z
vw6KHat1N/sLNqE6jfkBEjkhyQvF/A4QFQzM6IjdEdKesIMnwDxA7Y8d05vINhU2
T+Bl+NzlkCB+xnJHARdFqvTllURLj9gVQbMc0N+GwnOMDWo5BRXI7B9Hz+7ci7cG
ELefkXqLDKKYGxr99kahfZxZewHqomqD7AWvPaDRkPuE6flZ0yxMrosYfRO/E75M
G07n9vJxwbAqruAuwhDrgRCDMkSceo1SmaMihDTu0P3oocBgBERaP0BPngpTvYzK
xWIptxFydZVPhxWDHgeRJpZ6vNcQFwmf6zNTKZHCQPlFhvVjvhW+ZKe1V+M01Qdu
cRGHjd0CTtVkNLpN3UzK6O2HNHNzzgkXsj2MM3UrgKXNNL6P0kZUhjcd3t/j/ORn
AEXYjg+7M4yQuqpPz/RRUCrvqvGemQkuTtT53pu9TGBoQQneAxI0K7Mg+PYKXhtp
Inf6A5QcBlSxKuk6svdbw2aX+xeV6racys0TJF/cI/3CG5EBbMUHPoCyqUzAGeri
oH7lkx5UPm/yfiODnS6VxthfL1WbjWD78wVnU8PQ5t6b5ccMWkSjw8relWe1XY2n
mXhS42VO6ywcFE1AN88uBA//1mrQ6Jq3oI4qHPqxiphg8er2JpjybZk2pJYxJ/6F
Lxz30Ye5aYji8Ni8VhujaDfdLJp6b6eZAjWpDTrl866/cUxgJ29YPci2XsSodfCT
xvl/zx8p12/nuG9LEwjqVjpgz3IRjMYyKO8sXVQ2/86Z4lwUb5nySZQam11oBuzu
TX3IoiD2AgHWXzZ/s8kUwmXBcbQbxhiA2jwcdCyNV7c3SHwzD57TRxZR0bsqGyD4
jZ95lebR/7SRm9Whg/JVIBE5WNXpKrVX6JT+eizXZ5mxOTQtAOaaaGZ+jhzToF+W
yy/cojZQmlvyWGIVFhgTMAOpursDZS2s5peJgffOCG8rWPh+gt3UE57bW4ur8Eyr
WJjEA8audUjObM0rye2mLlEeiiEUdo6obod4qnPDvKCtpAUZH40RfVIOEhWUY5lF
rdaxgDz1DI8i39Gbfj2GGjl1cpSgWiQYFH1UqqwCsc4zePA0oqkogHz8J0Xi1T1O
baF8Ce3b0OlE9wxBYmKax/OsJb2LKRG5zu+qhhPFt2R2AgsAvunKDeILzBTf/FyR
izCFUBc/xJoH+otRGZuE86UBYYlCYUquSlb6ETAeVaoXzdEw8C7VIUt9XG4Gl988
BXojOyRVk0B3Nuinpe7ovxiFLIZQc9A8uUi63zOXvgeSaQatHhcSZrVSFK3aVMIq
HpUXvSgNhA3mGGpuv4mCwCWrgzVGhJiP9gh6vk91tVlWHA9KaKF6uNrGWbJ+Uv4O
JMMeeEkOgcmFlkq6e0ZyxCSj0if3pYBJDScaliGXAjEiOS5TEDMFZKZZHuWjSiRy
dwCMWBMh4OM3mbNCiN1u2KfIAVoR78Y4weQCAEJnjc8XrIyIOjXuo5cnuMNsCCSN
T1IgbkUn9sy/lV7bMSgCbDJce9b7cm4bUvLQxcwo+WnzNmc2Ott5hF9LMg+EueKr
DTV8ejE5xjjUpsXIQev/PX0F97orhssxADimkSq8yrlSLMCgHan6l3q5WFy0UpuX
xOHyQN7pqVECXrZvkeHlQ0mOu6hxxks7eLpSjcnlq9sN4IYWniJK7AiRtt8i+AJa
ziTv3XwH7Xh7lRLSelL9O7HR0+5WsL9Y0tCiiw1Is3s+0trZJT6XfG8D0a/DHuPg
eWqRFz/aZq2R/tuCVfUrw+IvCfIuxKRZ7rukEaGUYg/8aJbUI49X/MizzHDEK+gT
Ef/Tc8++rQ6ALX4TR9ppduqrL4QELXcT3IyyE1N/pOuLLWKBHsAnqmo0Aa/wg4mJ
N2zelWnF95+1yvo+zd15FE9paash1DQ71DjidUXCnRjn0fmMck0oH3+LZvoxWlPz
YWhvlAZooGcEULoE4YTMgVSrnU40sD3AEa/nE7Bfa3Ej3N1ELmHmIgyAfl+3OyDl
x5+94g1hJjmnRNn+6hvK09GXNFMwZkoA/VaNfevMJPIL/G4RDmeEK98VdzhCc5Gd
cxBTviayKJbcaXUJp22NHUUy9TD5+d2XweJKV3Zu0VCbVQoPhUbfQJbIHQUKiSvB
3gv6TJI4ffGFOEkW/c8hA642vD49DfidSCVOCNy+mea8U8ZpJ86dabqoVUF0QpfV
DNq+dNrA+FzvHwkDYIGJhPNMOmMFHzHk+ol28hI+BoNU+MmwTar9JZG4sa5sV4ct
Syl07l5NCn27yYN7tjuXmwS0w2kIWW/oz6V6lRsjhESVfxTU3N90/3xJYPW7X11+
nnA9VUbWEM0/jtYitptbGFson2kpxJRE1J4AJHa4UOgh4lCr6+P1D4uTkijG4SfE
EJF0wYB3Mwm7cXZQe+OebD/4K3izgXxocIwkldGOe/ZN0BL7avcwLRGz2HwQ2iJa
3pWZKdkC6ipFj9SJgzewcUPPxc84x86m5Hh+TupDDGcoha0rHzU4tNlpRi2/lb3P
K2vtC9T58g77b1IUs+8dH/xpKIgcqXxOZ8JEEwcPQxUaaaJqBy2ZS9C0vePkFJFe
1T76r2S+xF7HsAOKh4dC4INl7Z6HkHeTBvVpr8bQ7SeKJoUGe4Gb3IyEM4puleqp
4X1/qUpSCdpvBq0DinHePfBdGIB3ybExU4da+niJKtaUhM4qsQTr9ijYE/xyzoWU
O/F22yGneAJtnIzODBb7lPx+pL6bUbuYsYNS4MjxIn3jDft+EnmVW/fjJQOfYIdo
nWxCv+Zhbz0ZNMVywhcgHBNu4rg39vJfaGZoF15U7YcGjABf/YGoY0RERuaXLtTH
vW1y8z4xzjI3U1bJ5wi352N8imNKW5fxZr94T3nsZ3Cig6V3FhdKLCCZXgm1+FYi
ix3itocKf6jFYcggBAWyu/aymq2SfwVhdbaXbz+LIpet9BLt11N8j7RYzDWejQoM
GTOVePZIJGLr4kreNdXVNmUQFhwwweNXsPRXco+MvcB/NfKBT1NGtE4NT3XxLggg
8IJXJUOwSmXYl+pbb6joMzsSrYZPRy4sxFk/3fN0xWP+Pz5V8IjvjLjmll/MY1Ob
mIW5Wy3Cnt16TH6fxbp2r8+NMkMQeb1Qd+30CyT+yy0111s3/iVDIE72n/vqWMDx
AXvFIuy3wFA+Ybr1it3Y/FSVG3kRor7HjvcvK16Sj4EQPVQ7jpBrLYcjRKcl42Xh
W84PM1sz9y/fzRTX3fBaoMdo2UwklpJDu+LBAjKGGyibmEacz1JBTHEnG/MjwH1s
u4H2WWTD09ou7xf1pbQzfpWOZV/MPo/wxKnypGsrlxGODOCEIjbB/ontGbhADAOF
6yq7wtrFnC0/NjD/PLLYhJblKDnMh9DkGaTVn21KnFwXGQvJgoste6KDhwp/rZhz
bpeQMX0aAmqxEpEhKFH+gkCOuI1lFc9ZdFKlAnKG6iqxniPWyM0HTx5VfGZgJsdu
fD5BYHhYy77a/21KLv6JSjxKS4BhT++WMdiqh3etgyur0obLkYa03EVHM8c8phpI
XMa0ujQCwFtsqdr47QKZxZ1wUS3/yBr0KTbOuW/OWLFy1TQoyOxJ4269dsRaMzVZ
L5u9qFhIpwmqDwqfHRx+b99aVp+cljA21D3Ysrvp2y55PzNp5Cj6hBm2sUgWP03u
x8R8m1Co9CluMPkyDp2ytmwZ/p/cqIba+dMFSFzo030sna244heDONCkQg06mFa8
pf/YUQb0UEA4SqSdjq53VWN+xxZd8vU4X191nWrpGr7ZIOVsV0vReXRLSzM6hb8A
fXe9EBRjtC47krW4xsyKDBkoFMBfk5yJBxOSDbbqqygyeKOFHgzI8B93KJDWFAaT
VHIHueLn98Pd3M0DdMxYAqu2XwtnfJO2kMJAS35d0DamfbkuQGnJf20WQ74C26Zl
hO2YH6TUl+h3zqf2c5+DyZk9UUe3Dq4gWulxu6iJm9MoYz8LpnO42uTxyDvFpHkC
OGdJrTcYF0OocxmfQ3Hg3ljt1kn9pepoQWgidu3YWOlYgyyMNSOUe4RwPRUNvzs2
h9TzwS9iRc+0ye6hrAYB50e8BQtoc60OKdjlxS7FunNYzb1QzFuJ5qPBeI+LemCs
mwNBEbS4Nufa0l6Uaa/iQzYBN8uoLcMTD91RmIX1WNpimVqKYRXuXqo5hKdQR8i4
YpNaNOefOb8CYKW1lMirVN+O5S8hoYxw8ULmOx+BFX7CzhVXXwW5bxNaA9OEWmXH
aeZrA0LseK7khKfuU7wxeZgNBXRGIS2uFpjJSSjT5SzpufA9jlsOhSi7YIAq0gqj
41iSGcaTa7ilpC3am0fneKzpdAOpGHBzV75Jp3A0xS3PxGLAd9aWziwgYLEjUUXj
GQ1U7gpReM+TZmDpNzJbSN1GtxP4ymH2B8yjvKXAHYdJsjxNNIjxfBVAAah29KFA
L9+pyYAe6IySyG/QO8qu2BhXYM+js9eBWe0ozkMn3/SkEjZEEQbKM+Bn6eLYOIr5
hz5uQGgYFF3IJ7l2s0sRRnDl6DZbVNWx38ziWbkC7CnBKle5ux0aQUN3VNjnDTlX
kF/wKQ5XzvYe1jTAZO9vF0LMubCSm7h6JcHLFf7XPzUAoQh8S+Gb+ozCZj0jU9l3
daKkt/0qKiS8lCf3q6P1+oiGjjVrv76RCwrTNtd/6prCIxIqColrDww+PuwXo+tI
0frk1K3Hs7IdbRGwRvXFJ747UC0qRy6E4YGZJ0fUTOSt8f1Ws88tf9htGg84tzG0
sQfO9NUsh5vR7SUoSw8m/mm0yoW5CL2WiBIE1ZrHOil1u61JsNId0m0EKW1mTYmS
7oC1Hz7cJWnQHR4sfVrzqA4/E3iXGr4MunxbbyVQgfqn7Ac2/7F3B5uwE+KjJvbc
R6UCdfaKf4GK0qGOGzBb4VNjCMiqjSRoacAzkbn7NYAvR4KIdw3GA9PRm6LpW4oz
NHjKZIUC1cjEtPcw/pdhyaqA0+mgs9/YyKmbKRyJqM1YjM0CTkwHIScEtd0ACwg9
M9+W+NcxNMGWUki6syzWBm0M/1cnAXYn5cJFRhpYs04UR68yo3kOUi9mZ/MqeuIz
hjeZDF33cRE9GxQwPWECbxtvsJkyekHu8wwqT8WHfny2fBjcq3qOK6fwtH6I/FaE
Gm+RXcAifyFHCwvpTnnedVswk+D04RZwsm0xxFk3Oe5VSHZZyOA8mxrjM6lVqsVC
LI0i+fR/OicBgDn3E0sZGH+VavlUwEp/ScCkoDbH1OdlvR36r8IAM/zOyrPYGjt2
1bvd4iwefzZmEf8GBQYksNemoh8fQDyk3ChWy0TBnUKjvVzieRB3YTt1AKafFOG7
aoORtTaCqVPUJMStMv3L1LxpgvD/W/rav7qvspS2jN5XoGgIuzvioLOOfbuHJOTt
8CkrkfT+/WjjqGICrBBfL8A4q6F4rL2rxxYu4UDDgwv2lBjT8NApldPoVmARnLL3
YbRJ8Dr9KZNWeRWqCnueYtoo8F3+u5CIJDgVYaAIbA2pFxWsZaneRik/lAMZq3Sl
RFxaA6mNiTOXHDosEoZYYKO7AKF7ogtKbyjDHqBScHZ+E+Wj2cNmw4oDxmEfth9t
6zp/tucuKDF/H7RElAV1BU6T/ZOkvSZ57knuiXuLObcTHmHm+b4yLPiIp9YbUAgr
IpLYSG1TM4cMqtS10M8V+XYbOHjfW8P7mprj7zraWDY0CUNC3sOJtCPGLgRMJvTH
SudaImaECXWO2y7XzJ5Pd6LIjEgn2eIXSiNzOFefAC7ANsLm6s44KWrHlyj3bj7Y
aqlAtZQxe+yyr9jmlgnjXZgTuaPE0x6wzLpj6T3oby7AgXFe8d2OoZ4XNwo4XPJR
O5D/KnzhVax+s+JWJdIG/K/CVvFefcqij1zqnLQXqmkk0a3p8y7N+rqUenivmkAS
y5S2yj2zeTONupVwX2KtIw6SbuK4ta/PriG+gFkHZSjwwlbIzB7amj0dy+SBlAlg
f5ORjfp97zOaiPIzrzP3PDyzzKB5ly4HsMSathk856MNconV168LwK7vGaVcJtlk
qk45b3ozX1+HYAYPgym43dxb2BgtyQdplG26bEhY3NaKF+boSk79LkrPL6/LWqnI
YHnjaBxQ4ycB+B3RFWv6xsx1pzc61Q61GksQJB3hSElY/F8I5wXzhTED8mrGKgzN
AndgcBETFV8qOxH4SzwdfQBBGGEcg/7aoqa4HUbEbrnNuYPGJetSijo6aO2tWRY5
qqFKBTw9jo6lx298CFNIHMumCqQCthnUksMAKdnrjQSU9pGQ8PEtNKBg7PbXFBuC
9TxuWPbsgus73KUd3Q5GblBmaqLXkintB22f5hoyJ7jegVS7pXRIP9v647tPqyBI
PsRIdk3ujGp4MZR+GEQwzXTV8vfRP28rHP0newtEogVq14tWfwSjcpUD/bFniPT+
u2rKfqxbbavQvg0bq6bA64eUhzO7MvQCuRJ//PwUO4cHJzGETbQxMzZovOVEyB44
JcZvZkcHaijkhlgr5eU9B8DmL/yQdQPrWRkLaDxqN46bjJEcxM7bvEz2STu9EYV9
0AlcDk95P3saqCP3w1fFIeLHh5bd/eUoBJt63ERSkQLhpQ7cvwjcflNc04dSd1FV
f3ueOzUx++IsPwHPLeBa/BC0CHYZV1QlKSs7qELhZdKmfjy6gcoeFjBs7bQ2zDJb
axlFf32op9zA1XoQ7XAaaWJ9nvH6paf3tgmQKMOCKjD+1aZGDU13EJ8U9Vw37/6f
i4ZeIyIdCQ9G0AhQU85X2sA0rHEeMatrk5FTV3Oe88sG62Qv1NrqKV8M7XFPVasL
vYVPR6TkPsJ0CPjYUB7DJYgbeSQQW0NW2/Dmp9sF4RANcz3r2rAoVzUg3hkHwYZl
vrURnykY1Zg64k1yxVVk60B3Rxa1jI2EP6BLKlTvqWcT6K58WKMCEt3/v9xoQICf
mAKmv7gySzRimiWsHO794fKk7jJvSoOYfluxTwUA/6juCPVJg6CWqKq6Wrr+oM0O
WnRb2Xa3gu18BMWNGS9KYlxwy347Q+S0L4C+1GcE8umQQ7o1YN931ve4EB+aOwsd
fB61RKM9mfGVwSkkI1VnLnI+Uk3xmt4BvCuVpG5P9P3tyWlIlayI7JhVSlRG/d9N
VqEiWOGKgwK+JZEWKweztYmrN3TJJgglultKBOdIHm1DkgCNTogTKHxNAdEgC1W2
GWF5E0KntBvX2CxP+j4Y0GsG2pq1Y9ZrxAthbzEAhrUDMd9woMcFtzdoTuOaYVh7
BaZPg8gGHuTkvzNO0avJEqNH+rJ2xWsOqnjnq9mAA5oAkTBmmrHqoorVTGtITVJd
J0sVXESILdTM/xuGZykr+tAgB8AHDyXLWavGQUOJRvcWzvHX5YzkTtpAWujtz0m+
pr8aibwIZsDsYU7cjdupwNwtLGhMYckYGPv5mPDt7W0lpgAOmoS5D3qs1M//M+bB
YA6Rqtdj4z3hPIHyt97Kn0NqFsp0P0Q1apzq5KfZTAC+Z18t44MxQTznOdUwxZ55
ruuI6MCx5LDHGVB87W+GvoYdk/9wYUqnOmlMjObmyQqa3Zd8r2TYQkhHGq6PgiwV
Mvw8eQB4HUa2tV6QOLSIQLCbmg++1QoOgp+CEF7vHWqU3N9hlEiWX9d5eMvNzFRf
sr3XeIfenZUY420D6Pn/xsvIiuN3HecqfZj8YQrKbt0AsQQLCDNK44U49Wezustt
a6WF3OzOJW4ghySgJ8yuzXW3C8lwxu3YJD69OZloJ/qhISK4M9hcJCScQHHWbvQG
croBt+6MIG1cvmBt70iFD7CirLDVvNMTX16yfpRKyrME86tLmFnG8LuZu4DpIwvJ
Vx/IXd9g69oxH9LM8u6v2WRC0jRCE7nKbZgfdyhznfiua5hU044hVvu3VhXKNKz7
9BBdPz6Bj9Cnjzd/vMN3Oke5d8SoGdrCQmQXWoZeVOqX+7DzMh+vySNumTc+NimT
dAfur+ybd0AQeXf+wZ1q31P8ShcfZ1KLOWCGFS5HnPj7iKyPpul96q8o+OZn6P2q
iyKPIfdXGQ7AAdfnfNdpNoeV8bC/7oIpN99bG83hCaTfbZPNwGDXddDTp8cR/0FW
u1ZftV+Wblc+VcbXYtnHvaDT5oDae2ndHuGXuuSrTNmMqgffYKrCX1/STTaSMXhE
POBQHnHzmnO4Ntfhj0SCnk8htiOGEYiFVzCTAlUjPYKANsNLlmQrW9jCd4lBeU9p
fD3ziky3YyEoKX6bG84UyV0FPt/lgvwwtj4gcLwqOZM/0Tm5YnIXCVK/TqkWjgPD
PafoKZ+E7p9RiZ28KZMVP1rbnIE11ktLvrs75/22hj7xFPNGXHkGmEmMO4d02NdA
Kmtjuu/lw8FcKtcilykh9VbB9wDKFfRBHCkfWZflM05sTaqqfABFADELmunAbejm
tExi/o7yjD3faJxD9KhWpzqpLjXOzMGmwJkkxJVTKi+hmTr8A7aI3KlbSl4aQsEK
KNsp7NNPhuIJgxu5SnofOaOpi11hf61hCuWMTeXnl1dIYFtpZGEAsd8u/wzSUgYq
VWEeCwPl44rO0X771twBUlpzDa++l/+u1W6Dj3d0fC3BEJQrWS2CQ5DNM13ImeXT
ZgZHHnUmZrji3rimOuvUEOrhDioMUkX5GWu6CS8gd5pYDIceeX6CqI/iQKlyFwRU
SDvp4UZsfquYlTTiqwhhYAHDJYPvTuyAyz0Tb34BSK/Q0aTowd0EFwsniqt0cFgJ
y3MItwst0mtoHQ1c0wf/ygTSKs9lXj4GG3qVR50yWsxq/PvCIng1XTO4c7wonrgk
FyHZd1uN+5Ki2Pw+Yw1fFYbp4hiDHawoY2bkc/bXaZuOTlGJ7iYr/ynC9CVEGcwy
oQyrtPH8T8bVkc8hJviO3BeLU/qAgGy8455NesnSWvKWkCBHz40Vx3NIu12vJlWo
xO0Uzm/uRsFwBM6mWW5mQg1eBvSwnuertnupZfXON5M48MdBL8MVyoadVphHHOgT
zEtWp6yhBh2x4GWz/OlzI9zdS/uQXGgCnMllc3X4xT1UunRv9x531o+rDhGMN6hs
RR4HXwvL1bYoQ2LSqp0GsXBYnomkOjpoLuPlE8tcmXe4KjwMgrJHosDSXIM6SPBy
I06dIcxiTIWzk/cDLd1atfhNUvrETvYF03qOxm8OFgHpU6Hqex3Ct3jnUx/bmfef
oHjIaeUkRA8P06t4NURG7UeF/4BvbGhAolzTR/1qaofBDWrlwKVSbxNtLtsu+izT
IH6ldOIfVJlbnHIbYUJ+P+vtay35Av51zt3Kxbgi3RC4H7a1nEjM8kZkVJV6vj+I
CHFOTjf5pmqrmbs3e7iT4dtl7zlU5OWDx1Q/P0wobVfu9D1z7VQ7nAKtQgXOuph2
KkrnODLWjHGda1EZVsoQfDQ4PXE6s0qCtkqUC4jFWhd0W5Cpcem6kNpi9ut/tlat
wUTRK8gi0StBAXOESHqiD+x6cSm+7JFZVduyx7xX0iHx7JZxZ9XNGhRYP8mLBDHv
ecabutzxPUkM3NdONah6o+T4ibrNq1ewz4qM0basbQoWylXH5zA486MaEGWnPMhm
i9y2OlbC7XOlx9ZK8ujAX5WKDsQsUFacvPxWUMuwwE8Dq5l+GYI0sb0wQuL3HMqa
5sTBrQZC0vsGwRENwieL0DBy0ZrWspKLw0+HZjY0CeiZDw2LFw80fHX8PSbeDuPb
TT63h7zW7nJhBIbL7JbY+Z/4s/XwgD+d/B7R88ARcjCq7MJGL5trMiD7BPu+NF65
mw5u3cYu9rsn86tuwU5mxPlLKmOykvVCJzH4cV7NTrU/KwOvsysIAktvbR5JzCFe
IbPIldxodZJW8FV/mudW09Djbsp/F73B10ApVVf/2hZDQb23DsKyJA64U4rhCLmx
ZNpdA82NgsEDvFzmKVBqCLyDfSaucvz9Z2aueN2bMKDXMw/DSVupDVyUsP9JXi87
S0gBC49na6DZ70Tp3e1K7DyfS43sLy1mJmMZQ3bdNm5b3NfkrmWdMSucw2RR0hPO
k1jQxvNfdCj8uaAIEHXZc2yB0CzU80Aa3yAjNw4ocVapx4BUPKTT18fXEHfeFVMY
DpvkKhJ0YGH/gZ/PbmTPEy3eyePXbYgbq4aXQ4CAhD4xig+821QVnY/L0OszrWLz
ZHaV/2lRiaTsguy2q6wwnYAdsZxlQqYxGJTbKMNpdiAzAf+dhKvs4rfkt4NuSg7H
ANbNIy3lpTMKXaem4vtR6GGWweEwV6FNpbDu+UquyTgOczOZSr186emunJLhumL/
gVhkc8QBqa7IPv26oJsJBhGigocsroe4OfZuJGUn0OFQxexFZtFaj/MMZYT31VyZ
pXcGZlfb86CrINY6J6UkCfaQOkY9dv8sRpO20CeZmXHj/BZLbal384sWEoxp45Nz
QvNRqGBACdHoo61Wwj5Q5F0eBgeetTBVvBLD+pL7KOkR6ObP2y/NX6R+ba2cSghn
AIL026CDumbB/nkh79YixmuXF19VPshTDv/Yw2ksh+v6BSNQNZEloQBBW2dNpORI
cNxBaRt8tCvpKPIXTQi6nJ+jTbaqoWJgvZolMajrzugxQn0jN/HGB1spW4DLvUhl
WHGMlTrAvtGFS80DdtuSgZEOkkzqyybh1rzXoD4fR9ktqGVshxH/mGuNzW0iowk+
7Oph7Ud4RMpHzzLO4ivz/pvK90i2pAAWs3vWh6Ud0VPgrm2CoNsFBUhETyh9tGSM
EPpA+ULccjGZZEn1Kl1PzXUoBcBq827g0CVxRB4NcZ7NTUPMK+Amb4xjiB4aVtl1
vXq8d/hKGIoOfeC6bgChL922qOkXEssVTD8XaN5BT8uucixoZYcqYcRirm1aOqe0
BuDM3k4kLXcJi9IdCAdXjFme4cAnSYaIjg83CrSt81xE+hpcW1f+D4UxMYLA3yK9
Sc0BW9UHTGhDPGul2Qhz+MpFS3Eq5hxWY3b0cs8fJlmh2Iltn9jImO1HsJYJLrhf
nwcbs68Iw5U3yJEm/hl8D/Nw881ypI9WzlWEZ0Oj0GgiyfJdBW8ICuss+QdyQusM
Yvm+pl77Ii4V2nwSzwUfVi10EBPnM9XRpMbnbW0/hyq0YJj0kqoD2hMsW9UBKJ1c
absm41S+hliPFoRPyyUOftc54zntoIc6x738Tfpig6nRK7NqiZUOQtlJweYQIzTS
fVRRYIMgzujbsJGsbry29FRVicuLtiUcAwcUuEX1K6Cmby7tCnLRU7c+svquvMOW
LHwCXk5t9z8MThc1SwXwkALd/JVHWkI1H1vRcVhfqXMu9IVgfNXNFLx+Htd/L9Ub
vTldaLbDQ0SiI/OAmtmAlBi0vpAc6jB2dCBTkk+U13HmpeLv5Jp2Y2djvAuO9IMe
Epr98IpTvCjAven2kF8IZNNfQ1m4n4MNZvbOKVt/aunDsWcL+iz1S3NnAkvzuMp/
q1Ufd6l7x46xH9fmAPpdiIyT+tEUGA1yhU1ZUocSX/eYbuc+ADIPVF1Y37asEz1u
AQ3v0ewfZOgDsCIUphvYk/g2dS6ecXNnQKVm4Omqa9P0sfeg6bocoJf2GSUu6ciq
M32TxnExR2eGDAW0d+JTZQppBoscaKQHnnRm3FgoIMVSSc8UjFt4E8lu7aqFPw3c
kHq/eW3COmB2H5I0ISXdhU6AOrv2r4Tm+F5RmK8AwYjB49Zati2HPPhgv9wZrHnQ
fkrGG2Kbe8D730UxcuWMD2GprNey39LDxurYiUEs6fGot1pFXzycW8QK06uDLiCL
vcmGcu/nhx9QDhJtT9DN6Q1eSE9To9eyPGIXGYwbuebplySbwsrGwSHrXxU6Ovza
7/07aypytQuikd4XH4je7XKQwfIPqTJRy1V4ADWNCtlUYIhJWGU1aZ6DE4Q2+6JG
1WXit3NenhcSZ/R66AEc9rNX/qi25EjMKe+wD2+cBNDYYMX4j4thqg92klgufre9
s6zR81VcinDMIy79kqvYq0aepIlInZY/wEiHoKPzlQTI56rK74SS34el743qfa3J
mrU9m3yd+x4ORHbELmJ2x00dVavaPjpO3zhirG5SScZhmnY5PEVq1rWdLye1Jr5X
7b2cSBnhgdMvirY8rEbUVdFz2tEdaGPozqsB5cRpkipQdewGZrUdu2LpQm0fDaVZ
xyKKYn3FgAukdje6QkcGVT7Rjfvv5HUDQFCBaSodTBz+LihiN+XsF+nUW16PNj6s
dR8mMPI/K5qx+48TMdkGQG/HW/qswH1GKvqwiBmzeLvg5cWIagL9OUY0Lqk9DioM
nMpA2GiGCHS4HYb5x9KqyWJKzjsGoOzFfC36AZyh30qqQwS0jwOFoN/tfnQ9hVST
q2D2Cdj8FmxFGI0CRIUOMDSV5eBTwkRR/OZkfMOoIPQnY/q1gZjYJf8qxNDe0HDX
DZVIN74TKyOcOppeIvq1DhAFG8LN4u+bAh7AmliVm8dR89sMM7HozAAlLOEL3/0C
UTJgbumc1SeT/HdSEoMBlKXjDq1NKrMk8NZ6CLAV88C8tp5Xb6iD9Lx45SGfbsuw
AQPw1dXzNDcKtJ68D0YlpoTonqCU5wOW9ksR4M12geJWaiStmXQLo5WyA920h8p3
LCOsLZV24j2QSVEciysuXlNHUXj+o6uNucipdApFxUIRUBNyTPTG3nbBpSv1cb21
UtP2C+ubz94z455mXdbJfJiXVuqUzNj6/0v6ZS0396AubQFBYDnXuera+Ye+XOe2
F1tlJxgGFquwGYtO9p2ACdRc0vx9Uk0BULOKsbto0FFit4NZfi+XCaOEDlYIuhB3
cy7HdQ/vFaul/8DlB7rEI6VU8PaIUpI1z83EFW27ucVDQwuccnPcTCM+FfVuFwqw
TGbF95XJHP8CY8CR5CPF/v73063DrhNTA0tOgQpMTGhHA276up9NhVhVW8jNqGhX
4DZb7WoYQsT3jcD7264QzKFmsQzdE58OHqkxhSVpgDd1RpiJWPaxiZZkHtzN+VB3
XH/h25LABGLGJ7sRWB3tqJyoxQ1lMQY0ojjd03/1sxjlCGo8KGYcJwitIIDUJn54
SJnWJAqD5ELqrfBNWhs40GXDllHOVQrNvxQxe6lWLu5aYCr5fWvAI+UnesHBLMiH
fF6BGq7mncJ6pdNgRNSewxPsc3AudgMxS2ju6pRwA+wGUBdUg4khsV9Ry7r+PdyO
DCwb6bMnU5X20KwJQDSo2yf1mUO97KHH9m9Xy02ZEJA+wSdODmzsrnRorngAZh7n
vCn7ohgU7KajdFJmkcHVmaFF4QIHAQAkpIoMVLtivRIFAPhgFQS13qoB9bs+RBqQ
wsDBqIkCR5CnObdDbaunJ9Si8URUyZH/jIOkp8iSAxN1LvvBj4Ok55xPwg6tMUMk
`protect END_PROTECTED
