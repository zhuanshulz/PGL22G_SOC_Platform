`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X+WefHn69jqWXIjf08mwwOriPESr5s8eBiuhSkEjuOsYzUcv7b2uGw72ilvb4f9i
Phj9of9x3uGpRUzn0gozUMFOx4cGufcduAi4k7WSSdgZ0HiZNCAtfyvwtMMYOweW
6rEhgrcTer3aK+fzjg/8pTdCNGjhLCyr+iHpmgzeI5MWjagCnkQmXOdN/MZReten
qxfrwibgpLD1Ydg2eeh4L5a2IDgKM9/Mdq1hWIdURtzguidT1qHy2rcC532nkk2+
ROJ6hyu8l10kcYPx40g7FpQ+APu/aU11KT0rIiaC80t+8qL5CSB+murzioBSMIUB
ZxppwV0OJZjpeESfLEVxFTkPxFfQP8W+aLrhJAhJxPKmr99/GOa+rqCHNuZjDqKp
S8JLm2qU0KSeTmhewqxD4xLOiZBpv72wIvO509v/r/n4wdrg0MCnjoq5ZIArmkV+
Ezo1+ZmEtpihA8EoeO4QPfSYdV8luew+ygrsnGt9+2gp1yUKifw7yTzdtHzRh79t
brHdyPb31Egab+SDixjWoiJ08DpHuFubpMi6uREHtDHYzGSN2IRqhtzVcoiO7lsk
khGwjTl1HxLFuAwG44/Ac03DwI67j/PPf20pkB2caiiYzBGhepvm3gE3fgGg2DTu
vEiTPEqNmhtpTxCPYWG5jmOlIxawQjb1VKJZ6LmfnJbdHwpHcMQV9wa1nPTFkQcj
zOuAHjMHBw7+rrTzZpBNUXXr7PiT7lIbqOiFkuMIDqQH50VGqGrKzUg7JrQN9nf4
YRSDf7wl0u4/jP5jwXUdauGtctY+iiffYhtlCWwoRx6yLzjsmQZ9ldQqC8qsbOC4
gA4q4jOkVC1Y5KpUbu0zkpXg/VRDKh/qbLzd/C9TPTrOYNhepCpoyuUEpgz3FYZf
Sk+HPuhaMnd/vZfuuA5N735MR3tsxc/qkozxoqOg5jCk5LJQm4hZo54ShyXikunn
89oA7KdmEdodZhVacAFvp0XU/5WFdPzyupLW7jj+12qY5SN5iLeVv30d9MpLtpLt
bd1Gq3x9SiQbMEXDOqjbnN+pdMqifPJ1WDyAvcdVwAzjTN+BEUTPjSa5sNpPFGRr
Bhhzh2vp4aGYO5O5wKQp/a2D0omGflPpT1m+4GmJ2E1gJfboGfL9ZsT084udO7jv
7plXe26hqh6DaIPwoJtKsPgSoQOeqMRgWz3OKlz5WfnoFQPncalb72twJ81D+H9w
MTIWpa54U/bkFik3N9D0zxJarLJmNDuR9nfgKBxIMtXvyUZ6X7v5kvmQ1HcawAlB
+7qyq8LeUMe8uXgofvHFks1OGaFpZlEH72AIs/wcoW8/SAKWbcWlUpcVUwiWq6TE
k0/tSKUv7oQwn/HManAh7aLHbxZTWhYWg165Yze47nv+UcHTSlLAIwGh1aDbNOPr
Ds2fib7PD4Pen7zgYm+7NUWNF12YubBD5W3OyLtAMwhwm+oQeSZhpMTJqeSSpmze
ocUbrEo1c3mFHHCXG6e+HeYH4U9KcYIqHL23tQtHOk3Fd17FFKsZQYBIdrKS2THA
ckDbp1jAifhDQBkJeVHC1BZC78RJ5CkT7VHSrT9iJ+t646gi3jHRjCdPavSTSzyo
aMhLjuf3UeVnwxacEjWwnukR8e07cze4lW+iPognlsK2Prr1q5wXUKb9QAM/eTLD
KESGmp29DX3qr+j2kJDzKUhK044IrTUQU1mevxH1fXjJNTyEwiNci1fflw9efaaa
LtbUDC7D2ZT7QKqMIQJpgpTU49x5vwES5qKntyD7qhSAXf7V7zEgytEgiBwkv7iN
SNlDdsY9qSTzsvuchyUw7OeVqSEdQ2X3J989yEGTlQxq3TmMUfRQoYmBsxQHt9Ox
9UXoNXGPfe/8252N0D6IJPEUO2haRQ3kspw/9sVjMKKGrxUdeRqKk/XPKHzicfou
oufD47mby+MkeaJ1rEP63qGxihCCCVcRh2xX6YttYJilntFx29FZ/aH1m2ydgCSZ
y+Ok355G4q5/H/LTcgYJYj87MJWxnjbAo0N3cOtJtaSgMOMjsJjmZMyzWBN/ucKE
w6ObBALE9GUo8wDWIgpZ64VuPsnq/hB0+JQg87kSwu9IkV0K04pet2kc1PGBFFAp
IngP4vRsa1PA5MAYNf2uUyo8CKy1q0XOb727477DIuYtPM1HUVfkYEFL/KWi5ytv
9xP19yw4i+OcRS2BV3fLhm61p0WXl15CLl+lpV01rp7Q1cdmmMMKW49I+WltVCd+
Q3LNINxjdcyf2KO2kJ2RZ/0N3fGBYEu2BZzjDKfuGKQHXIYUHVBfU9kK7yrDMipc
b3yDVh5qosI1bubw0xW8AHI92pgQmFv6D3c4pHhF/nV7p3pijUWZKzBZSTGg34E3
IedN/1omuLv3IWEIhYse45NyLkbhZZd+2cl8UmbNKEF3LafX+WmZpWG430JUbkvI
moErU22elJA2FuTPiwXhcZm8tj98t9g6MzXpZp0uyLNmzlNjc2zuzaEGy1JRYfrG
k3y6M4uvsDwXTzI6wDFA1yEZnd7jM5g1SeTZOJuGFtgZKxXaQOg0zbE0D6NmmjMo
nasqAWEEzIfxI25LX21W+JYD2XeDSQHWdKEtE8O1WUsvqi2sNvk1JhwZ/TRxfmby
DoskJ4GzPIfO/b/it8+5cJW057V5r18VSOrOWRChfbg2U8558Vz+mOT++8UeGUD0
DPILYpP+EFpj4d4+lSSQfoDEZv6v/+wRB1dDiyMKRZMg2k6nXoRnsDP6Onp5CqsT
N7XCaxnjrTtSlnmjm5k9m54brmP0ezjuoecuo0kbSsVbHKf6pMwI1hdg05fEJBhN
a0zbjnI0/7YiLSYbI21NX1G6LcCK21uwC756YJ1eeqkKHscQ6vxXh9ErVT/TFRbs
u/7N789b8h5NkKRedXYShoFxxMKEftTFRzGWlma8jN5A+ivSQY+TgM7nPceXzQMI
`protect END_PROTECTED
