`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+W/3UCX02hNls4727nftzs67rwLPk7Z+BKQ1tFVkRD7YJVkaVhRgOnLK7dG2GSSY
JmKzAsn8W5FJWzu/EzefthRsDoV+AQ0vAw0BZhHU4xmcLDjtH0+HogUtXtBBPAzR
ZbtyO26AZNx0GfCosNyrdl22RS/YddZ/FwcPAtIzEibI9+rd+fiFOELZ+GRC2fh7
siowNCIZDDJFyT0PtqTo66lG9giFzHLtYazCAyR1gxywv2MiLLLaHVNgMDp1mEBq
GQGs0l0/hCPCIc9wwrzuuhPR5q2s0yXTp6PMTQ8tG/OafllIajRSC7LiJcmHe5Fx
297ekz0KSK9/wP8Li51QGniY8UiZbQfLpsTBJQZFzywnehyKS1Aapenty5s6TdS/
Cz2SwdFMa/aL9TVKbZFJJxk26wWQPxmqxH4VVJ+HeCIDEaSy/VrAF5AO7MQ5rsQl
u1+E03iMYYtZ+5xX2czwFbip+H++89ou/+tvTsJq+FQ2khDqkQBB9mV10Duu3yqJ
TRbrGysJzwbfe6YQdHBwbXhIWZkvCUugHNe49wXhErTqLYIlWwQMW95RBePiNi0K
Lc/NaA7o7wvZQBfM8WQXFEOEBIuLrUR6Z/dHKbNU9Cii+1Rc2totIjsQZtWvW/PH
m3M4jPjuX2mIS0YxWjb5nA==
`protect END_PROTECTED
