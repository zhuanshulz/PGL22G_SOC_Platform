`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TvTj8HZG+5tg3buwzLRHkSXULeLvHow9iZdOrD61L5q1QtmfcTp6JpTH0b7GAyuH
Nfv35VPyh2Q+ptCJvweBUGMO+RPlZboTtRxNUD4cF3UBs+iYKZ+zh+XIQRBh8ZK8
uKcD3mENYGCCe+Y+3iBLpwYi/t8ABMjXmb3CjSLQYb1VL+mUboywA+GDZU6ETnmq
MU6H10R4VTQkGJ1v2btL1PulajYyiQHGinDsrXIiQsJM4Bat/LfShD7HbcuKRLq1
vnc2q9ToGXPBx5KXYsWrkWIZLYlufUcik4wbPtED10kTWKGwjpxf5w3WExG+1xm4
n0VXZNMbYGK4nBMtcqudYEI2qW56CR5/1N1gWAQJnB9Ny79iKemIQDd/R9phRcGT
aPDm3UbyLmFZXnV/fwGQAYNTE6q6wBhGJ5tAQHnBrlMtN2S1QF1bvGXX8ZCaItOg
uhN1GL1gkzxjf31zcm5pZG4SO1TYIMTobWTf9nZO5vf+NM5z2PotqjWydm8j3GBS
FKE4UPgOw9v8b03IIUfcXt0I1BWXoBKnTwjaFLix1J9P+LzM0KkhaKc8k+KxMQLZ
EaEccRFYkx22ZTAFGuqFFZW8XN6/3/IGfmPrnsVWfUpHHSBbWmI98qQP4fTvYqX2
oFu7ZHvpStnziRngeDCQ+spUIj/sBNmf8/19cjZhKjIOGgw4g8RwsEgkAMQvxVrH
ntYqd7d00fyQLvami5z5KUS4/DYD739NygB/7lDUmyhHMH3nKjzAFIKsdSfrUzXR
YTLa3v9s9Xz8GBlig/W1erQiiQzYcT/IC609Bp64Bw9Kg5dHydpxrlYra7EGKGBi
c5NEFrEvmbiMAkIDbiitlc7vDHbhgURBz+3PCwhINjUw5LUZ+neW///Hwy8888on
WQacG1tKbLjk1IHIl7P4hO9a5raOdWh0dKyEqMueDioBStm4xJ3pmI/50Vr3cgL3
emI35aV/3RnAvdXCWcU3yEQ2ofDkfz3Gqiz2VOXOhC9czWNNE6dGS/TRGOhotlVc
c5IvSb/guunjxu6fkRqJ50fQ5PpCaDug7EpzNtnGauwr+DoD6Ws0yNWTh4rFbr+z
8Rpy8dgUPuB1deTHvfH5rinXjDe2YWV2hzEU6/yWumw3fOuDsUCp65Q6XjK5AuAY
vUDOCXJKU7/bLWULsUTYSDWJyz4LzwIv7Y2iXUv5XZY5TFz0nyEBRC2ATaLeO1J5
1QpB0jskUsCRzu0hyboNMxCQ5b2nuK/iN0tI5WOhuJ+llwNtOMCHlzN6doUrVDbS
9O3p9+xvzsDx81nWcQo599pdoENs+3mDnJb7V5Y+YEaq0Yr8lO+yXRztv3W0o8fz
csdt7+ztwZi/cw26NJujDbc5X2PedKj9MHbLhSXEPr7SWodS/Bd2lgYZM1MkOK5e
G1ZAvWYVZArxbhAOHvD0dPQf341ka6m9Fr7I7KDeyXi62c4HTc+uhfDamCjs9P+5
utm6oFa8NWaNcLDtwpcmVrzDMKXj6BTdIxs6LkJsOLOjqD2von4ZfuRz9K59YluR
nQYuSHt+I5EGjkC0WprAOQcRjhuVD/CMQTipI1/4hnBJPryTUQCqOhbsdAhsuV0M
telDbnGqrz4F2AwDqi0QzpDHUt1DXH61XdgLGvDMKP5tEbEC3xo5TQb0pK+K0hS9
YVsRlhfelECIMm9plBfMXGdaejoqKTnh2eE2EBuTP2C/o3Hp8CcnfUnLyv7sgv2c
YL7HnTt3YiWoHHOeRTnV+Frcay/d4L8I1uAppXIHbhxtYa9/mgm2yKM1dwqRhV+1
dDIt+5uUgr3N7lpq5QG4lOPqthwuzwAxnAx6L8QjFQxzZRLYd04yzchU7qFWhcFt
6i3LrXA2N6pUXMg0pnev7+omSryMaYrUmyaygytdVmaycPzvDwE08wHqDqB9fw+0
j6cgnYFSCZm2zacEuM2m++VxvkeBh8U5bRJSESqvcbZxVXGlXtmuI1/XbkbKBllN
sp5yzARiP8hTGmD8MwK1FpO4/p+H3JbOkYxAgrymx+bC4djDmVSSTdc6S7tq1oPq
Z8Fh3SuDd8N9ZEnqU0pc71lGKMf8a7mHg2y5REvR4n/q5QhjZ6vAcm34HKdlCgzV
WpEb9vmoyNDEry+kOfYUSO459oRRorO6qPDRv9h4kJIlHV84CBvk1/qpgM9wLUbn
pGWzn/AxTqBxAWMbUZNixq3y8D+EkLPcDZm1RL4Bg3H9MGDCd/lVs+nTg8FmFb8D
qjfw4+aANZQJ2gkjsq+fDoPiUIXrss/43cQtqkzLJvJye/+miUuhviHrefa9A1N6
pCyxIOWWFIBDZeviMFw5HgKNCVb0t8MLNYQcSBDSaXjX4IlnxNtOYCTF7sm4NjUb
MB0OMbsZM1MNuxnZ/ZST+xzwCdpay5B3BOWinCFOD/85gAe4K2OcLltoOuv4mjT8
5hk3amngEdmAYoX/uu+HCbxT/jamsXZj6CrrNxgQrfOLgEQmt57EU+OZDmO/Mx3G
HvfVVeSLOA+0EzZRpKBnK44Omtt5nI0IjxQeT+L1b0jzOb5AplivkfvdvujXL2f0
x3aivSWY39KIIPIk7GOZiw==
`protect END_PROTECTED
