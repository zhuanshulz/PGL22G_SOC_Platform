`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gc92K99v7HeO6PDEgjbmkLLHX41SMmsCyfzqo+cwdsGMLsXsb+50GTV0g9wZkkXH
WjFzQIagiGbgfuJz7UwNTclLdL3XjKGI8NvPuv8sqrGtJkV7zZs72naJIOvFdlWV
AfwameXqUhrj03HPH2FlsAGQ7il3RroCcGZcs+5c1RXhMtawxCWq/aYu1SIcCG7s
6JsAIzmBomXQnVDDUSWOcjqI+tguhDix7xPjxv02OjnoJArBs5Z6RhUCoo609WLp
h7cr9yd+IyTbD2DnH8QblSP8wSiPvzP6TQ6iMeQ8UbjF4pKMpxEGlr1e1QZVVpGw
lzuB50uRgEVINJ1tUvAvSoXXU3GiuSyjFr/3RpVdWqhfv/R27GhiYl8XWOwL06or
ZdXIKbHtNHEZAf6y1sziocsF9DlwNyDvUXk8dhEMyMio6J55szPEavJj3HjVfIPu
CUhRu0vvOwOsGUkNGOlETVlmRMbONaHNoiCsQ+ZWmPDDKj1R5YUoghdVw2YGg/5k
EBi/QvPjRjvIJIbVOTEiT+V41Jf0I4m3LnVwITSd7E2laZJSThacngUZCBr/d5+2
Em0sp4cBP4spCK5znuRFiSbXbgTXgQlJ8EP2EhQ2Vf0=
`protect END_PROTECTED
