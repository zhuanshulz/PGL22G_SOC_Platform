`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gbbteuEt5+tiBHuTipPUhbGD55nq7+hjyd2VKUBtyel4aBmijHVziiiHFB1W08oB
VDzSsKJhwcyuXvDzD2zcIx1aEvKibelyJG+C4UgaehXSzoUKiYELYR5Ta9KKHi+z
Mtm2RMASMb3HN2SJDXpaxtYA0C+ZLpdNKEPDxTcLwTwWVdhPTkfhbOXAvmWUI002
HMMguisJdIZqecWBkp39f1EQIYaIBbqaRe+RJlUzOfLeqJSdubfHDG31vfTlzwl1
Hkd2ujaCWwBGYgI248OVHmRZ+9XJUGUrNQtkyzV4tm0BJzKpYRgNd0t8Bj1HWsjP
TimcoxhnfvwCtI+76sTrQtqqTcrwgjMu9jkJigT/eHuaaFQqQZz5y4yrbVFNo3rE
FsDPvSw4aE8ooEbW+96ixeAPnepRmSUv/d0FtDHw3ZSZHEb2w2LVnkTYmninmafl
by858xfXC/WeYF7zYYBvCwqGYpqWCVjsFj+ta4yJWCRyspbvmtW4HjdHRgHl0kBC
3JJgYZ7mn9D1yvmKDgz5KTES0z4rRTjEOggXAiZgB5iPAzp/tQuTKj/VXVkGSBdd
pxicYpuEGhG3kEIYE3KScuBMDtjST6uQzL6cXFLZO1CyUBHn9K8J/bb83qkDpXwE
6OFjsvoeoGQ+iO+IKN2esyOZYO3PmCM31L6rBY24fxUp7sRau2HfbR/pLhwnxJIm
keiugJoOW4JUVlcfbArwqU1sonzT4vgnfUNZDP5jG5SW2eHDWGQBht3LNQDU9AJP
qpB+9JYi7NPu6ZQCYeeTkBi4GI04tc64sG3LQ27TXkvH/+PopF0bkBFnlkgX3eWY
/PTEDl4pfDdoYP1j/qq+hpsqd15I3F5PzDKUDCFGVBRbTP5CZd0Kwb4JyDZMxbs5
DGF/datkNH05351ODsO7N4/fRj+x0ASb5uAZv5O0jrxbd6Aawe7384Ak0bAvfNmn
il7T6wv9FYvIZobg3wbJfkCVzMsiS1T+BeT/LsD6boWp+VD1sG4igagGYS24reQ5
EfcE4ZG/i2uwX9NuCgos5cnvidFGKBLRdpBR359HhSWWtXIAuDq9fU5U4NdbvW7I
pkBMVtZ9LhLeeNIFAx34TeWOtkxoj3hzhqUqrEYjqTBqQJIOtqP2bbe1lowUGgkX
c9U+mxHmVeWEXdmj6/hoIDrltTk/0IqBtCNRRKeHew2ocV7RE49D2td99bwap8my
rWfXgLIydd02Xnt1ezxDH1I5ROFrRDtnTJCfxUstDCoYYjy+ZyS/6RyHhD71HTu4
xQwRJOcX1el2abh3pBcc6eNNlk/bPTPgN6fbWIa/uSkrgiqw3n6WxM6CuxEbPY/t
jqwaCWwrObVdBvlSLJLelktpgd2ewl/ZGx89cGiiwa7FyDy45jPkmCJImEzXi+VW
VdYBy2j33whE6J6rH4IbKd8BqdU3yXj3vKz7a8ouNfm9iX8tYMnQvFTG2kk5A5fC
NS4Pl6WpZeCQeRkmv/pa1x4bM3asSlX1MMhoaO/q9dBQv0cwJBzaThtMyCUs1CnJ
Xn1v+UTma/vHaKLC8LHKsjMfM9zwUVeGPr//Jj+OKsycIAHQWWQuSlcEeC0Ekj0M
ev8X2F5NQah90qGRQmewX7qIndu1nF6lRmc0/IQsvwVlnKH/vPkl/O5wHaj1hLJf
YqT9BroFyLCJTDeR/VAbmUgAH19AFkFYtMzUi8XP/ZdQyIHrtzS5nQbM8bdbZw10
QvMmeWYpdAdeoTAFhdfkcuMABl41E6vvgZCSAAh1fVPoPWv5PgJ9z5tg0jMLZs7A
RUzKE2jTHgKu/l3Ip9bYuojCfWp7O/XM2Tp9UO/T32m77VHnPtzVTD7z18W8Zke3
NBYdqtT0V2BXgQWsNBWr7zI68Hr0Ii+OKOI30mChGjE9AJSXZeh3Zmq7ZwrMS2Nl
be8dLu/77p2/wesOZ1/RyFQ9uJhz3CuVQSasRpXBam6jHE6rQarieTiJF+T095OX
DMLtxChur0uiIlfKOHoqQypiVkiYfb057lnQTKSzabpVf6C42iLild9mNeESUebg
LAXA12KnrywS6o6rjllEXQnJITTN6vekXru2L9+PvRwGC6LR8BV2YV5p9lXDj9XO
eppCvJ989r5XTLVDltONToHfPweZFo4yVPrbd5LKy+KyQcyb/PWfymWSzvttIyOp
lQY8SvaUh97q1ojBdoXcVTQoVHYJbXnAZt2p+6WjOOQLhc2ohjbbbjSb6c+j0B2H
b6awdmJnSA2+92oN5wmNrxyawfrgWmWsrWdsOmxcDSOYw0AddfX1dsSZu6msa+On
QdiYOE+8b0DGi82qEk6dHTTAk4OP6jIdRXLYmSaiBKestgL4Wo2cbmSI/IdrYYHe
sYy9LeeqTGjtkZUkk0WZvjMmBN+lEdLuQaf7ErNdAquVwQy47ejNZf4ucN+3CL/C
Z3BVrqz2pvqPLJ63MXtAXyMBGZdankxqI9dylr821/UfW1/5zWajdlgdvqgwJVC+
4XUV3PBUHUsmqvmzTQqdn1QrelbrTMlmJjpozQA+vPbmFzzO69Xq9ytiyLWL66Fv
LW2I9mTIEeA4KB/4XPv5ybB783bgZWzeM7CKxb+vslAegZIo10wAGLtGg6RHTeIo
t7SLeycYhcNVUZNLs4EXDfASonGRrAwyFvfNbY+eeofGi352ALvA7sayAsK1Gmx2
kbs7dSvfFdPohw/ma03wi5PNNP3oZnoKfljUYYoJp9UgYxv/2uB+vpAk6t7kWlhl
RUvOmF6JbM+MD8k7V+fs40oeB6m7I+kERtSqRCsBN7shJNZc+DUWKKa60V1LGR5x
IL1dcQ7BoPRDoA7aN52V2osI/I5xDaVh9ogLTHpN8/b1PtuQ3Fx/Hpc12qiSNSFK
`protect END_PROTECTED
