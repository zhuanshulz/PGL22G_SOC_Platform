`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EI0emquegnyuAXC3RZ6EaO9ezFUBNaYWMk8LIA93Xtbx1KsU9vclz7QqZkpRh8G6
/r24hxBy2YvZtiVSteph3d1V8f3RTgiEHi8Teiw7SDUKogd4l6+dPvNp/XvNKtSV
q09x35NshqKf/k/KPyBr58rQx/cstU8yztLjf2AxjQa+byef8qwiKpn5VSGEhs8C
q1GnJlDoTUCAv3S51ttGb9V9LuZKOK/PRlGA5+lr4bYkYE63KpJqFlQjs5RT8h9M
CPsgsf6CdrnmsXEMMU+SenQ35zjBm92TiD6yppFyuRAx41tN1bOC4RDDhX/A0DWF
42xutzIhSkpG/KN+Mt/5PbL7jqXpFIOWTccep7mveBoCqPaYm7y9BnnoNgw9HPw7
HCMHvcTlsG4TNH/7dR2Un0gsyNU6Hh98entKu8eFyidQPeHFoVCMdDUAsFbsDnOj
vH7U/G5PvgfTD9X79WH+3LFzhLSjtBegm8CavJwwiOUyyvui3mTSvZC2k0SgHYql
aV50Prh//iAVpNlIxdFJTxPSm8YJ8b4ThR8pt9J+8XoTQ5YqaJMOzQBqmxbGjfHI
E+2AyOdet2vaPqFigR+zlzOPnUX0wSbjcy7b5k4inyu6oTBnuoHz0IeG3tlJea1r
fBCZAAbWJTLKLFQM0ZoOo1va8NsuQaMonft8fKOewZHGZkH1oZRDjQ1PzMwjsVDp
QOC2Zx3wLxDdrFEZ1qiY0FTMoiVI2INny6YV708h/zsCSybxztIZnrY5rW8E9IBR
/qFRcXMQLZIUb/k/GZkIccxa/8bqX5wgyQanfBpI6C8u7xC04cu4fiDvwbo7UAwk
vNGeW85ro1rwL//u5sVuO5kAC7b69ghv2C3GCVJLLIA/rOxIwZwaYIByn2riVvHE
k7RmqJBy7EgDa1zmaPjke1PgDhlAoH2fQ7POFe+Jw9U=
`protect END_PROTECTED
