`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5Tn09HzKNLTmfantL/E7vlN3rDYPqrjlGqn5ARqp602Vfj62+P1R19IKSeOwLhx2
TZsZbaOz/pJ2GEQo0dngvYS4qmiTcM0I0fUiNG286TaJLfkY5kfeHRdDDvg7Qm4+
Zo2tnOt99onGuksvXiwnjPV6xKvleHZKcVNyI/b5vq5jovnl6tzGbjliULF67FgP
xRf+vWgVRggIij4BlJ3WG35pL7XjooAgYsL3fL3qy+2C4raidvfWQT7UajIkdzY3
RVi3AWuaPKS5WTUZ/u564a1GXr6oVedrx3RXvmelA2vbueAJ6RfCOMdibpZZsdYy
XYLYx4ZVmHU61BJUMWKF9j820NeJOEd4AKPeoW2jliK/quPVKBBv4v9UN+lQNtyS
bHsDomws0nfJ2wX2t8fQl9ZpSm/I4pb2skQmnUk5oNs=
`protect END_PROTECTED
