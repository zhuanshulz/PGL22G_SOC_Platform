`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kR3fPdM5i5ig6DMxTj7v42GFd5LGtt+UWy2qIoptquZhFx/zMycjJm4hOQwQyh2L
vCgNdL6VyZYPz2Su9n6JtncjXT/6qjUQy0bpIeZ4zw4Wi695EiTW/y4wdGqpBdOK
5SPjhyNYdRD04fbV6a51gFemwJYfHliIK5JVkDw7Dlp5XCOrpCMuavxUEapv3vm7
CF127cdqmsy7F7GXOmO7tMS5LMhoRSYut6s8IX0kxSin5UCr+dpBgqDY8T60YbBm
rCi2ObjikyIObTb+xLfQTUy2XCPZLOJvs3RAkH2pv9CyAoM6W6U+oj0D4tX4rLCE
vxM9Z7UkYEOXYb14NU4cQv7ELnm2cwxcshKX3M6uYjHv6lqrUfGHjs8yX9ubA3RT
a/kHWry+NGDbxzqsSxCb5gm/zHj5D19t/PxLA0if5nvC2mA8hUs/gKngqhq7AUH9
D9QQ1wguOm7oldqWOgREIoRgXqXebuASxdavvmsT1zmDQH9ipUy51Jym3EtteMWa
xTAR9RZWmf5FDCCppb/z6MlXwtvoECiiPWiI3wAYLHu/G9sDM0Pnhjj/o8FCJq44
GZvSChi/H0WZkRsbmim6oTqa+GP8at+T1xpBZavmJFRWZy0XgP+5Yjra23jT8zjo
ctWCJydiGWXQkozFkEkY8rLVpFDRZfo68womdTDrESWbb/jNFj7a6zHxBGkjqzm8
K14dClngIYl3SYxmho0ZXwp1K5KwbjPj+nBdyB+q2ZfLccL3cl/EEviXf8eBCAyX
OakOCB2cMRrE+3lw/lFzuATlUfPZ5Iin3E1zBxwj2I38FjT+C4YmLqwQZeWnwtvs
TM36akfKeu8gwRVSbkjhnNClRa9+eXYcU0d5GJ29tN7a4h9/lnOCHzZeuFvA9U1g
LvSqsU21hu6MawWjseX8kQRGFkQJHcpnsdy7/1i3XL3l3Oc2a/okmdhPbK2YbEAc
Ih4pVz341LtJEZo5yuNa6tmkrqTgYpZoVm9odG+BMkZfN6X9umiDo+zCUxiCWcqH
hwe5zjqOJQXWtxuGEYqqOurcXt9l89DmmjEFh54Fv3eHld6iTQkvEOXnGZWZtjWb
A/YimanWeWFLcuc5os6hGfAIKJYq3FySGEPUAb/yd6b3mF1yuxLRX7lQJd8ZK2yw
uF+kVIysXKER12b/InzjMZnQzjCEgFVNNm6HQH7qxs5JUT68qri1Fm/Lh5jvPnYj
rhLGc4yZzhNzsXGsrHkAg2I+kQPKXtlnujIdfK8Qj3C6wVnv4YApudagpeX7bDeB
`protect END_PROTECTED
