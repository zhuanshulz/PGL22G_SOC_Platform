`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1IWTT91NyK8C3q+8J9EGU9kImt+saB8nSbjGwrRqKAXDJAZugsW/p8ng+dn/HCLV
y3hC/dtVx8px/4Rkg2YgIsZ4da/zASKMWpjXDcjmu6qfp+f1+j8B7qY6K8xl87yp
05H/BDKbAg9WyqlTM1tEpOaaSROZ8km/xynvkWZweVuemK7SZ8nJjIIR3S+jfkNX
lMucczGAZT0b0EZc15wg3XxE+kEz0GlUYtfzs648M6v30zWXgW7q0Dksj7rP/xR+
GORkYTxaI3mh+MI6EpfAoCy3xYiQc5xlRuBhMwVWHhjBHeNpq0ao8857aurSKmMy
v/uy8F2JKsnl0BUCWrEIA/MUjfzLFMV51J41iH267HvjQN05K3mHnhZMzUJvnsdW
RHvMehAsmVblAHHUGFr5FDl1RUCJDX5/TCg+dN2L1WKYwBJVEVNciDUqoRY8Vr7c
rQ+BAkCge37YcTqBfjx1xeajRIdrFNVSGFKhEZrmn9xaRpQMw8pRKrgv4ZqByKjk
HGVPusRohdFbBxFwEUH3VsEqLg1e8HYGAzCJ6wViVgFvmVdLY6qWDZv4QGLqoLy1
Xg4UCX04wVfdXR5VvyiyRxeabkoY0RDN1ZUujbEZSHjNeoy7bntVyW2R2k8yJ5Mq
WmDA3MdwO/DsFXuEdCwmeyh8UMGetHJf7mhL5jZxaLd1kjWEX36xsHq2Lp37kT0/
HmWj350JvgjRuMoIb/za7ddsrN+sAefVEbdWXZLd4FUy/U3yLhRnPhzuuUtb6+pW
JhwmwuFjlcrhw2alYP9kJvNlsnGStEf7ZLorHMDzFRc0RLsoGTl2A9q2lwLKxPyn
YrCNDKo7/Dnsen0ZOh5shw4blyCt+CIe7LT5n4INc3kjG3IIrC6Sf6BMbnfDWTxb
RaBC2OfWw1UrnyZjcRGfxpj1xsPGSG4Q218vN7XFbXs=
`protect END_PROTECTED
