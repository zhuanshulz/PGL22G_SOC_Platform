`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ur3gbCHUfgkxfkhBMJgcDpwAYAOl+5g4N5fv+DTAIqqDkTU3CgaYyuAFNv611tRH
OmaXj0Q9BXU4SNLVjOwNKqHa0gCOsEZyFQmgpZ0I4lFLK0UsJ5u9qBjtCUfm4w+w
YrHQiiXqFyIYldbQ4KIEFoy/E0bwsgN9qRwWPNlS2WQypxRi6uWaeoQyuokmdX+q
hhON316exmOcH5veO7zvte4aDQIwR0bGvm1i12dV35Yij0eFKA2O8CzbvA2lQ3UK
baq+JO1HrQqV8WV0mQH8fURVUjTuM9Zl5+y7OikJOqY43NRYdCY7Vmr+UDlejNYm
GlNAdM0IeZnKyLrY3A0IsPXhAy8Sk/neaCrlXlh5O+R7JPGy0NVHVQFtw5x7GC3T
AxLwn8rP4DBc/Xh8zPJdzrg1ThFPvqha1SBS0Wc4SCFwfaPrH4gI4CLtMTimcclH
RhE+nF6X7tljagdJ5xFoonvqZM3gIs7PuQalo18aCtOxM/m5vmX2PyXNsfE83Ahe
GQeZGFZu/rNh2PYZgSVxf7pnVdkn2WM2DrryRcIJpjYUr6YGwmXe09xM1TA4XSjz
eERGEmQzWjgzSup+IfnR0lvinbXvp5NIDfTMpFse74n+B22kUaebPxjp783NZLyH
GVJH6G+okfwFA8dXmwuvJzDKvcvbFudV+nQqOkj47eff0ATTdBcCLDlD8TSy3NUh
+H+krtTZ1fJ2BvbRGpz1XR7Lw4GE2CHNyyGZMLMgj0SLT6XsluztpwA1y04rUlnQ
U3KXIJTwVm6dwN48WhkGr/2Eq1pCc18qnFTtYvnwu//vkrDRbQxPKAPynkgH1itX
gCjdQIByjdax8iCt2V7gwt4ZFl2h/OBaxpp8xSjsStlIAnNTWrrHS0U1v8dr+ijP
BNORzWZ4e3KommAvkX4pxdYka6AY3jkegHl0T/XfnbXwmU2tzg1XrRky8gzQhMJj
j8rJo/etZBkgxviZqjGZXC4Sv4kgFjTl2Zggd0eykFMa5FXQXICTC8dILaaHN8mz
K3qlw8rm705NRnd/e2hdbIp9GQIPxmFC4KUTtU6KPqfsPvppJkIPJ9ofDiWgo+o+
FpF4SQfxKB9Oa7VxZZVb68Q/vm8AZhzI/juAnJ+aJXnJoE4Js/hLYLhv5G7ZL31n
F+Wc1/K+BTf+815kiRL6xyxML9qyG/c3QvkBv1i1aCJUWlOP+uixOMKeKECzvPIH
K0bE6AnW8Tnv6yiQ0+S+vJiBKUg822u7NlB9q6IxS6czxLBJHSY5X8ipTmZ+FHkl
1Ccx6SM53klBGXE1xllZp9mxas9BNqhWmSGUK/ikOuTRfpB8KSHnEQpxPvTjwyov
YiD3Teqa4Wi21ECzJyTefSej/pFLA7Nak3AoQcuU47CP6Mnf7vzZFO+Zo7BCMZ15
sCIOv8WmbU9WIcpzruwf1AyKqPlkuM4LZN0Mdb310Ji5WR7rNz7TmK0DXjN4nRWH
FrRuka41JmuS7zA6zrcghqC13TevvzNo28iMpyzEZJ1YaJkTYtL5c4xax1PRZtM9
wvVBxY0qr2m6TlOdy0yhS59/ncDaDikvPEsI/RkXqflB+jdmfpUNwr5OD4/6t3md
arJLRGsjCuLhnvAFXVrEHNv8HxPiCcv+E70tyu/UGIrmAzGHchyFV8qljkP0mDNC
ne5yBlSBzMsT9Ndo9WkQ5pco2qp9qejzYnNomMu8wFOHHkI5fSrS6JtaoBSgxMKQ
Jk5XxiOSTxpEwuJ8eBg44ONHRddPgT3i7urbLjh0SjV4AcTFJzNK1RYs4p3jj1tv
cLHzoJ6TmcDcQK/V9vBqUi5h45FJIVWVM1sP4R+XOVaf6VgrEGcl3x7AxcssO1Au
1SRI87GfGUyhPnscdEQFJNbHMXiN2YCEBacx/W0Rw0GIoEHbtOWfMxi/zDFwOfAd
4aeW37hTmr2vd/PDlRfgm8HrsPKFWdXBft8jLkk9XhxYbM9Hi/BJ2rW1Zs1sy9Md
MYbiMYdRtIQTsJ24hhSGE3ro1vmNpJvUlCcmJU2h4nRfnBNp3tXXvdfjR/4mj3q3
NGWmx9TPqWM+1ju/3/KQfdNfBCoKR1eXMA6e+OBRWWGTMgTQliv/zL8/foV9EzPd
CPtfRZtutluMHOfXqrNskgOngYyaCV5y6KEwKc2VnMuR++mwhDVvP6Bw9KTXXyW7
kmjJcTNMEnfNkzcZW4E8pC4JdSas1/wZlrs8emr6KwXs1mDiNqyIQGTyVvxS0EDq
yp06fj2GN5ZhwPHaKfAvciVJoKhxtgpCCnquFNMA2tUfm85thj66On0hb8u7yfn0
f1n8GBbmtbN2KMCYFZcuyKJ1c86S/+sYm6keSAf5+8X2LnpIajh7DS20k15mwfcH
Ou27Xv/ewD6/kQ/pWDYiCzos6MdKLcky+OIu5ciQBs9f/cqOLC1yKqRLauSigvSg
Phn5+Dy1EPBuIS+N0QLHvfiSoziZR5B822rq0HvJFeVuWCYaEuR1gXMz5PmZISnm
X0MQu+8p0CNLtO6/sALXfqt7fQZgCkMdSOo+4VlPN4YL8c75ZVPPbrJecPiit5U/
Xx8R0AHEN4iycZPxHGspwBQP8gBUVSV9dErTrPYnME+N6teV5XA0nMMQey2WIHV+
88i83M3Pe2D5S1jYflFV+m9WxP0jsNS7+AtL5Ef8iUJh4jMgvuLAJXzj0PRVeOnS
ar/uetG4f2Ouw11nrzXJUMq6w7QycEfs/0XO3VeVzaEDNRihxQu17vijnihmvvZG
uzyl2Y31z3pGXsH6SberbrAp+YGBAVLRAjeVUrYTXCPjA1S0AgnSA0GjMc4h0o0b
OAoP89rSP5YAcMqC0pLsxCaTF0OugY4fsPIPyZitJyrJspzk5Qhs90TSxIIDij1C
IjUSQYVrVQVyRV22lReJyM+yLBzePQYtbex/zukbsX4fo/WlEhTYTgklOCAf+gjF
tfrWJoH+h8E7AmRaUlfB2MZZAeY69KwxLCGjLoGFl7TALr9r+2q8k5CarsuvYwnr
FkjzsYmKtWFXiofeaAkwUSm2N5rXretn5QWBMXeOhCCvG+JnmKFyIUl1SlUsOOHH
57wb3BNLobTjzEYaS6nAZln1a37HFoZtlyx+OtPf3SnBdRDZYmp08MfzwoY0vfrp
XVTJFDWAiVFzoscxgiKs5FDyOkXpQ1Pf5aM+IEAtc55bUlHuJRAnTj9BB7iZH/xp
z2YOK1IF4ygcOdn6QpsLinfzzteJwMzMJLtsmdCHlmrh+fUy+9c5MTaOunTY4/8H
5raZJCrjvKEs51EJDVEDiDWKZuBOUFZ0a7ENle/wy6Lc9GqHbEb/uTMD1SKSbnZJ
63unTbIQj4e1IFcmX8zt56ocZyV+igiL2ImHGCFV1B8RQd68EeuZY0MTaUHI3TRU
fENbwvjo88kKENSo7sd9PU8tSTcvESfP05v4xAWYgEtSOWADC/tiITcLD6BDSvz3
bL3PE6Tpq/xtwP7Jlu0uEG0Rp68aRbYlrPKe20fDQnvOtG1cNkCKp0TmjoymW06D
YTVUuoZThDggIHo1Tfg1I3eklVbsiSM4rDaqsmOF1dz+/4bsRHbMmQ8NfcbzL2JX
jNlgTLPOTxIOseBno8cJh49JlAPCwchBTJfBYcpmCLqmBSKNFERuOXOvJVuyp3EH
X4fxWEcjCqfHZH5dt4/kNsUonaQebT4qQWCj011cUo5ydq4CJbUXIaL2Yes7mDXs
FzK7Oj7UxnzDWA3QwYlg5tBgeup5OvHcsVJdJqUZUEa+9rXHPm6HLT4lIDCiOeKS
HnObX++wMvYItMyvtMTG2SDkVnIoPQqph/inBwrxgTSx6uOrvx5GGgM3qqFtHVKP
DbPCTV/3mrZhUd4As6qEllSCVYu+4epV1wdspk2aiI4qAHfqNJUOOhYyXFbFOAWO
spwtg/V8Q2rAx8peG61wxcJTCCLJZ101ZJKRTEcCo3DY9UkexsDXZjg0JCnQ8SpK
LLb3GiwBmJ6kgAJhFGZI7cqfwaYNU2LnuAwcqMqBR7F/Ba/nM8IKYdMGyhuh6uro
+z/e3+90T9cpfk/656cmOAEWTgLo3scUcxT33ND4Oj/4HlDISk98y1M4LzF88lTQ
LFMaKHRCQfUpl3TnOsbjVXomRmPQ60vwTsUTb4YgDYopX/v68fZORF0QWnm4fsrT
SGURSEYxKjnb9slnO7ki7hETQYHd4+wBYi9koN3N7+H5qt8+fW44nHWAaD5IdIxf
roV8/90Knnk5I3nAtOSAREaqLXModlJkAD05NMS0bdiWjk9QOe9Dj/gT5r6DJDDv
l5PDZ3TjZUkz27Zmcrxtu6O/uCYYG6LdhctHJOc4k92GRWr1PRu0Toft+bvLznjo
xYgsP00afjGAj1JA4nbl7iwCAF21E7I2GeqdBjWdppqiPYh0IdliPZb2SuSVcLie
UXeoLD2CmBKTg0gWq1bG0W8RJirCewFJog/sqYSU9XFTw1hMJ6VnOYDCfCSO/LIs
Ek85wqnMl+Obo90xxmQYSGugPixfTcucL5nsFOfXCMgBIBuwtGw87bHEYoPS7IOC
vm40hwN72JSfKzl/drxzAAaSFGUGIAXiwbS5QhqRxXxf+vXNaGnOn5QhVkRsIhq4
o/Ysud+RHR8y2QJxzwtol19qzRFm+ph9XQVv/CpireRjVmz3l8PMNUev8ZcvB3Ih
50ool2RSvW0iGLjkE/5mklZcke/idi61gNO/IuOGpo2zLhVQztr1rj6bFB9scKOx
JUh5TWaKrXFUNFW24XiNwUvzbjHskd5dFLD4zdi2xPiWfbhCzJQPa3ElVh+WVSKD
GDYALLxvCgs+ItobfugVzJ+KrAyU28doae4IeZjEQ7GFrlMdHGNyslKZeIjdwKK/
77qwxM8wXdcVqXYL8ibF6g/4ivTnWAKrlecAxEBVkeHky1wJtBKBnIN2cjcLrGEI
8G2Ta2/pTor9v+9pKIl/y8naV/XouySf3teGFdLD9qHC/ssdkNdgvVLMpK9z5Q2m
VMHBfeNCIoPyWDFddBa8xkLIjTEhHfBtl2sd3FnZVqTV89VDsLpLgVoVzjcjYo8Y
LPIKODgOk6bos2G/SOhpXuOTUOfNrMg/52ebfiBnj5MU1X1RHbtB9vp38Y+0B/ju
khzmpIrXWhQLKhldJ1P5QbPBAmObuCPe3iJ4NbttGaybhahnkTzZ80BdnYKS78BP
WWdZJ48da62CjmaGJEOvrFqakeWAmXbw1RjL6e0aIFwJqJjbDmAobQf4qWK4NY6J
0hw8yV1qfXBVBgNfY6jWHD5JGg4rAP5n3ca4RBmSndxx9G5teAi7SHv0xiTuxd5Y
FjobAN/69sF5yROS9eI0/6Z8CxPTnT4fZrq+3+1tM4Eee2ZErWT9mHX3VKhMAHHn
N3oTbToMZw944NxqpIAeZttxhx003u9EwX4RmwLqm0vdwia6tV2dPr6T2D2hLE5H
vC+SDfoRGGcCZIJA5WjiV7sLHirrrlu1S+aZRv1J/Kx35VnZPxuxH/vMP23f30xz
so2jcFNFn9eTObyy9Xg7akI8iNGKZVX0K9R/zPgV1FIe4JHaaC518YtLF2ZNGdfn
6AwCpFCRygIOQ7Ot0OaWcG3gOzDgJtCEstAXv9dPDY/xG8fOxjsT6iYwOds4zNpi
TZ7KXQUCj/iDQ7ctiukbVH+aqCNeQ+beMUEdgjJ/DH5ws0Qnr5WBk2BAJoYJKoPw
tSL87/M3aduXHAa5vmvdWApqoGLGhl1pGMhbFgzT9HwHWj2saHFAWOEwAsdkmqgo
oD6llwVWqA4NXeWY9rLke/J3LqEGs1SO+jFE4pNXTuzP9bTUJY1hJdeLdFSwnOht
1ct9jwOH0F4UjfLvdW/I12Q6sBW/l0XKf7lDSRkB7vnyaeFtj+zNphaa3Au+X2Mw
g7V/Sv2UmjTmB6flJd8jBx09MT7AeViuelhwzrfJ6DDJhdbwYfUnjXmTCCOx/vnX
jXkswh48kzdqyfSaPJ2lOaitPSITHLJCt81Qw3BqH3EHi1GriNjETTkD99IjkB3c
s72u0Dne47NTBD/c9txOf1uKFNPPuW+VDiJIZy2lJn6etMlAFqKEdhuTpRnX95O3
Xg2u9sJxj0kN/Jb0Kf/aj5hXnTGq3kuQIaAfO09vvo4BT7brEy4aqUa3K49aa3S7
A9SZKyqetgwrDbMRb0cireFXoZ63HbNVAhJyFZ2b1d7zglYZvPbKENQR1Wrus5VO
e4OtcOew7SeaALA49/STQ4yoVJu+pWt7uXVpK11ViGqpmsBEqZRSTxnqQtJX7BNH
NCLGrA/VqLywcs5F388AJj7SARIsdUSoQpf91pWT1g0IQ+7HVFLRCv8o5Gi60yYw
ZYW3468MfiAu/pWwxzUHsqxgxbBoBJ2QnCky3CcEZYxeEg5Xxlcf1D1ktROWLXqe
SJVzCEcNmJG93deJAPabSL7NmnLvPn8QfXanNYuWS0p9yq1nhES36R8mEKGnlFTm
3uXvg10GsecFz7PEyDwV6A1L337lODeNPbqDbeWWl9YOnzPOP8N32gmKDtnOv40M
GhVRD1oo+V572vq58+5KHWVr0Sl3LbpEl42JhND+NtxA4xCmpUWZV7Jdq+FeGsPu
Pfnq9/AEFpJnIeDjWT1Zpb/KIoW7FiNPZ/P6kepNTsWhPrgJHM9Svsrf5hm1JXNu
i/9qrKqzjHyY6YIQsCKAAEiI5mkyRA3AduABgQUG/BLQbFP6QFL0XgJNhbiDgHRg
FkEOGH3b3j8/YUTJGbLWX/uBHIEgo2p4FhvOMuzT2Vv+AXrMktFY8PCwcpwB/vXE
SRrEe3VuUmhcpXDcN7024TtkKyG9W/jCdJaq0+Fg7bYlX0NsPa8GaTKjwIyYlwsK
iV6yrFnNGGE6jubZWAS8nj/YJGjW8XbADlNzlWQLxxrdmSl83folKZJbtsNLR+EA
tH0H0iJS2mkIssaDNe5aP1Zrgeirrtk0X5AhHjRFVGm0H/yCseI89W/4+d3mNhSt
KYbOma9gz21m/fwXmRWTtAuomF5w8BKd0WAnH/nKBysFSsgbD95Focz8SC6Ri2Nf
7H3LII1yQhr5OToPKvJeqWaS9CCyS/DgveXsJCTyWJtaM0OY0vP2F2XpLiXGftAP
Hd7f5PEGEI/RKTUjQb8sWgWCzvFYD/d0W9YF3wAk/Hdc+F1F9Qw94vzprKBkJ4VZ
YB6sx/ZvK1dgXqkD9H73vCgpvuvT9531t187OeRDcTs7iCzBBwYTdEzesDmiZPEJ
Tl/Xr9N5GVxW/62EbYeENrlj8WVl+4UeqB9yPPW/TS2+FPqzw1pkDLtWbYy1SD0V
HU8swyZNQYTDI2KbxF2CAiskuDKAgwlgDlHYihnsCIm5PeAIzPWsOG4iMeqVMRCp
Lg+CdKI4F55c+znFhzg2Wse7kzbq7x1XYpU5+n7ThCmC3pjSNdhpdd4gEO78DCUq
7UjgkeNJjoMS5lSXIQhd9yCjybHgLOm2W2CovYZliHgpOFUhm7qYYPmTUMNOrzmM
wdi/y7/91jMb90VN6BiarwDyUKuZHZijzs5j8MkkYvtkQouWaHCFp+T9GYcMeEGO
0lPmvCY+ofCmwNMBuCV9KtPQb5jpfmHLxQXOEZLoC9Nn4pTDfstAV9765sMaAtUU
aKdfOU5/1TUrst6crHIQ7Q4KXEUV2ftkAYu/WdfvWUzVnscvbXPekFk6QKJS50Aj
9GNABPxUn3nNene+bfB/MeJiXSx70Ccb0nlboTILWuI2xCf0et8TWB8PHOCyAubm
ZwyoKVGn3A+cipvZ+QHvqE31A3NJ6GC7WOv4UKFNz0lGcRCfHafxx4wd0FXfRClk
XEwiDvfRN1CGRFk0iI6mvBWmm11GORtA7uXM/b6YDIFe2u4J0zJgmVz0G8aLfn6Q
H8juZTSefo+sbkOxI7QFnJ2SaRm6qOhDR+8T+03f+GQk1vu4r0YOUMS71fELb+B2
vvo59frbmP5G3aHMW9asgyrwVoAg4lfxh7ZHLeT6m7jCVEGC6ruXrt3WSIprUtXZ
kcoo1zLwl7kJiU+G5WGEPKWk5rnaKqCi8nMmkFT+S0V3Rq6O/UPHCKOOHUQ9TaIJ
lBDDWQCUQHBO6O2nQVekVee4lMFugLMOEhJnLetperOIBAwrDmy9N7t9KixufAuD
yFRGWgyC1/vHCkVZBhrmXqgNuZ8vFa8pZHnGBdM8Z+rYzda2b+eNLfL7VyQZ00LI
hOnnbrUQCYfzO5/oRUXuf6lEb1rdb6ZNxN7VNP16QbFbwb7XUGB8of4ia1FhUEut
qBPBgYeqhTeYUhlLkFtpG0jb50rj5XYZ0n04c73EAsPaQ+33W4jlGfC26CZyzhdD
5o8It6Ao3bXw8GSYSLg9FOmTMT3r4bJQfcsOGoIj9H2LwX0KLnN52To28YeFKdNX
GaLEFvqDgSfG+6ZsvBsV9yE9ql4iOGG2K1vq+ta3g1z/xdAH2torfa4DHFtieIx5
ibh/BDEHHd6w0fViayJCU6Zx4DVnTc5stHhuO6D2nI7YtBZabQ2sYpWGu4z2ugoW
uTz8yg3ySoRMfsvr4OcdMlAW7LajR1/yLxS6FajfGTTYCVt+zgBF/igUoowF3U2L
idEARR/JePE46x2vtgz6xaNpyOWLWYlf6nFm4b5HrXwOhe6y0WWlwDX81Q8+7gT/
vx4PQSEIvSfHC7jeGdHtGD5RIm9/H5b9tkoloEK3dH3xcywd2v+DrEchrYcxwg4e
eHmpThR8hz50Y+F9KX8NVuTI9OpQNTtyYTGfPVo5iH0PpidM3MhOfhKNk1LlNBd4
JSzX+esl2aMeA+cwuubyKjRGsMculU5c0xm+Vbgut2pkYXcqEfBX5NWiIHWFbZjM
hz/D2fOUbSk3uV9hOk8gac/w9FLQzn/EirIM4pqbopT4ruHi9glu5k+6KIcNljTx
74WBN2ocudIvRg2xLJ4t5IbMw1stb2az0ZeRkQXlXtUWtgvtHBiNO0aQURGPjpg0
A7kyod7XK9wDFH1SnslIvmi6Fy2RkhUrLmqJrHIaicXTOG+Z9D5V+Da9q03ANKMO
riAsafv6fMKkhYwLgN7HT3v1jUpvEMOCnpYkIKqxcjqy8neCz+wjagdZbi50DOIV
QEKJ8LHdnHCSAe6c8EK9aE01CnpvFKkgRAnDMacSTUebaJfMSM7dfs4vy6qTd89R
C7/8QzPALTx1+NBokR3SGeNx68ddE3dQDlGrDQVLL6ovN9M6VqVjp/gq0ojVAGk5
rF37s7M7CXH8iTieRkVMmYJSj0510QwdqxUuuuovhzv5JTtR5K6FLBEdSL3I5pmX
vjJCaCP3Ht1Z0cyomFMt1eJ2pFGTbty9RyC9IF1W8aMbiX64YVci1FAvRfP9YnAi
1yTH4y5dfTILwqlM8rs4nBB18/AQAZ8LvtRJDlFm3MKNMj2R9KbuSVsSs6TNTkOV
kKAaVtN0fshEMcaQ7EDSH0bkvpvE8ESkM1VpzCgbLVLfDNXeEB2knNEHC5CVqJ8d
cvWM5XpKQARRQbiINRQoWAG3VCldxabxHMiaUm7jyV7UD/8W5xRC45BsyUapOypz
QLtd7YnKYgVGetUnJ3uk6oV+3MI1yu2Iw2+Fn4Ja6vonSJnNgQjhoBfReTGliAlY
5mwtE6VpQRdNJNKMrI9K0OhuvaUMSzyx7hR4GZYyO2uXvkN0vb7XMJT4YuRFW0b3
ou2HunhpxjVTwgomfQ9aOgJEcxJ+fU4pd+UcNu2G7DsuAmElimhX/M/njs1e8TDr
tBdeI/J2WqDHWUx0gpatAhWTrd44nIMP+iy6q+QPWiG01/cr/SU75YpeCpvipRjd
czbauiP3WOYqhAexFTaxZEbYFF4z3cTgYAB47HJXG74QCi/7xiFEyuVT8C3iTbog
4P5pmktu5qpRR9dZrMKV7osgEAKZhDUoUJrKwuCL/ZSdD8fXbCZZlupM3olgSZsK
nhi94/SmkKTeDQUCmcLVY4iZ6796MSVno7YFTDT9TzRj9fprel8RE1jmDYE8D9Fw
x3OENQFjSpRyt5tUdeZSWIuKP72eqSveVCxEJoAzXyc8ZnkiveE+7wad052TWHid
8ZMfqqTnwl7kQn6NY8BbT7pxMMACx4yyyjw3TL0WU5Na+j8Pl8y3EdyfL7pl+8ZE
5HChK2STJqqUH0CRBOE5jV5P+K821L8BPTRNetX4DEO1+z0iv9iagm1AmSfL+66A
LC4xVK3qQPlZugV0ivFIdbQC/BFoa4n2U+YBqLRkOIWeUsBpUdbQDh3m3GCwbtVH
/QIRrCHgTEMauTxuXIeSdj9Lu+5W24Pb2HDZaoTvDi7rxJ8BAGqNwHalyybyEIKA
ddA4sxCdw9x9SS6HLxrR/Pfq0C7bPDOHHfnoVzb7tD8m5dQvHl+gNLN2tPq3xHpO
iDxu+mI/nn418ciFEQlEzEvSrHtB0VxbCE+R15zsnzF69lhQPPS6sNKcJOyZsn7V
kw9kJ0f2xjAm93bVLtfjqXVFCcutpSdzbkyPajs81lmUPR2SmfePilidn7XFg7C+
VglWtRJqXldcUtqnT8gTrld+53YQ3Je3zs3/2/Qllpshh7gyng/jIh2J8HXBkrcV
labWrYrNFBdOkhO3AHKKCroslbwAvriTEHmY8jrO3B09wnh1laukQqAxVe9i+yVX
aXAzVOpvwpnRCDtrSboIXH4TTQfe2+owiXT4WGGEkUpqtKtweu6jFUX+ZnTuQBll
IYFsJudpYG3gwJY39sDa/qKOMxi3gEn3FxXl8wUOMOEWjiHny9CKHN6AnkUdQmws
whTNp/X9RMEpRWnlH30QcJc4kjZzMmQvX1nVbtK3fBLkyfYoK4SZk9aqBxECCj9S
QAzIP9sdySHQrworVpcRU2q/Z4L97wMd3tXXzT6C+wcnBxod5yqSgU2icP31j7kr
33tELkhiPjR/aOBbqtsHtt3aHDpNbt9Sh3VedDKPtoJ/+4zXExm4dxKIfkV5+Lay
0bJzbUDzFXVNYuIOzRHZchZJNjFTXjyQWk1w+VvVetkt4BPt1GMsFf2QJR8Parke
3PnoPA+PEI22jaAtV/FoWlvLrVvpLR5hs5mg8tEBP8bjkC8ofWpEe/QMTQ1EajX6
43MoJ41C4a0ICMKsMcO+ex16ZB9SlpQm+3tz6LN+AUwEGHC+9pDP3Jx7rkZZBe9c
HylGPt179MI4SmmLpnJJ88Xi/xNSB9PxCRKfwzqds7jU8qPIYb/th2CW3Yd9DdzK
jrP+nSxHxfZo8Zjzi2FTaxWuzJ2To8q5xu4QrU9nbcHA1nTDP60MAVIQuVgtkaC/
DcFxeUdpc7XG4LSirG4Uft4XPjfIdsrrGErlRMeKJGC2L/jF3gYOo0FeaOTmOWdp
bpRibf1L9nuzW5ffTfb06T7Z/Urs/cWAA1H9GTNyaC8tWJuPfavuRKXqInqIuJZV
pTwu0aK5g+2tYXlTNfZN+e7Lz+Zk7u1+ht4p2agVcx4kUZCwWKcIN1gniFeNIkqV
8toH6TnlbzC2Orj+0g6BFJcRImZhkY+jMamZNLsVxuxYCKNNQhqDJcD562B7fpLm
bFtzGRhDDhLhV1LCgW2kiyeZmzoH8FIb5k2RYPc+fXSlhF8y8wM05GR7vSEm0ujr
WFzg+mrIui0o9vNO3nFuzylQBMTGhFqEm/85yFbMWEN/iehKpQ5HghWcpqt1VLa+
BQz9oO36C/BUNCm8qWB7LSnahE8SpIHs9mVpOagwNh72S8BKF5hEeI62hpezes4S
qh3+/UHpzy1rsZgXZ53J7NjT11CX+dYytdRXXSf1K7YQQTswqiI6Zg+d9rR4cySP
driaanx0gDB4CZqpWQ5a0KB4cycIzCRCHIipHFQAddtKtpEiE5NoLXQlrz6RhjRz
j69KJ10mREkp0NROwDK8qnT6aYUXfjMKhAub/MCxJo4NflVdjcLUQ3YRn712HhWz
kRk6YiVcvfGh8NiBwqfG0Qw/JtDC8mhnw7Rda20xvo/BKME02nBgHw7q5R+cH5Q2
SYeZTCmSsyhncarq8BirNnmB84IJv7d2UeEPhUB6RUKajzbieSkar1b6Pr9UZJ/F
uz01JucdqWeJSFmbSAvq5zfgs6d1oQ5M0dPa4KflWw7uhwAvgdhzm3B9Zr/aScSk
bGfT3jnq1oolrMnzjSnQ8YkikMuvd5WXRdzvcO1dZRpB/AxJgTIOvR3h07GFLzWp
TikzGsj3V36RRsOi7wUAGyKtsT92EDfJV9uk8ROjGBNMEUmtIKGdVMyJ0yoysavW
dCKgEGlCleAvs3V5ODuB2+6t7EYeUco0AB/kFi2f6rJcDrl9gvMRFuHBXQrDFrt6
PXWvDEg0f1vdQ8UkrQ1HThNHaBJ7sDBYRkiDaF+W+wRTyAVqxDmKnAcdiQyjlFx8
L/viwDuGYJzDtVRjAag2W49E2erZGsUbKg8ulVev3+MmcRiO/W+cHEpVqvlKWPHo
ldEIGxeuvg1fzg3w3QZHN8WzQUhRV32tcbvKsj0QW3kR+fubJ4I1B8xb9sxV753r
6ns+KTvCTNGbctyNUaifCSs/ctfrvdhkF3j3a72HHjBzJVbzxJpu+1r2GijXCpQl
`protect END_PROTECTED
