`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AStyuKUX6mdApBsOsra5IaVIlOGlCFDh66QZsOn9eY/qEaxgMN7uyNJVpP++gtJm
HuTYPzN8qhKNI43BizKJ9gLTNVVYsNGGzpS3rqZFj8KRXkSULF69ZfX1rIyPMNBv
l2/vQu16JmqOVI95eC9eBUWjky96JSSLb5+fbivnpkXwdCCmiYhDPzsfuzHpe8eZ
flh/OwRZnmIOBAgZM46rX7dbZFIuuxqtuQZfEQyB4q0NDouPCkEa7U5Exeqhcjcr
X3h1zxm+cBLs3l4+qOYDc1rfvh+IxuDozzkn6YU98ZIS+gS7ABVG0rulnOkk580x
Nt2whS8RSrwKICQWsiefC4ObBQSWv/9dQgEy2pky1RbdZf1IfplQ2kqPGwP2k8p7
ev0sP5VGjfctTC9Iq1N1SgUXZTNtVfu3JAyD4nJhNhy4dfIxxMtgE77X97Cx2F9g
A9mbbKKezp2blxcqOKlB63R/FcwBLA1SIFrnNrYfpmJ1KnEhM5QGHw9V9jf9VAZo
sGcDcYzwVtUNMJjzjMI51sGOkwrZJyortoWWab0HSVt8n8dcIwUzFX5Nw/WWTRk4
nD4WGLGmpazxC+L0/fYSu79bqEicYsZQ7SlH9tAbiMSq1qODMiw9xjz+PJ+GJ+G3
+QQyisJsv6lOlczW6+uCs1amEHemgMNWAvsM26A9b6ZxPeN3OEmX1LWt33Di30TO
tJXMp9XMYCaa1/YuVI2nQQ/HxwbgItWSq8/5qJZdNMdlZy3QSS+r9clDMtsmgzGX
lZuVD5DqZ0p8/BrDDppNGncqF/COs06eTZ4tuqk2SEVBRSSZutftdVb9MfmKXOUO
u34wqMsWu6QyE7UGS3ylifp3FtcdZmRwkrfjZRwFuDGaGXeCFVMTvoNK2Og6/Mn7
bQzjLsuHU/jHeH+fawzxudj+pSkoNLmARmrjOEDhexg=
`protect END_PROTECTED
