library verilog;
use verilog.vl_types.all;
entity V_HSSTLP_LANE is
    generic(
        MUX_BIAS        : integer := 2;
        PD_CLK          : integer := 0;
        REG_SYNC        : integer := 0;
        REG_SYNC_OW     : integer := 0;
        PLL_LOCK_OW     : integer := 0;
        PLL_LOCK_OW_EN  : integer := 0;
        PCS_SLAVE       : integer := 0;
        PCS_BYPASS_WORD_ALIGN: string  := "FALSE";
        PCS_BYPASS_DENC : string  := "FALSE";
        PCS_BYPASS_BONDING: string  := "FALSE";
        PCS_BYPASS_CTC  : string  := "FALSE";
        PCS_BYPASS_GEAR : string  := "FALSE";
        PCS_BYPASS_BRIDGE: string  := "FALSE";
        PCS_BYPASS_BRIDGE_FIFO: string  := "FALSE";
        PCS_DATA_MODE   : string  := "X8";
        PCS_RX_POLARITY_INV: string  := "DELAY";
        PCS_ALIGN_MODE  : string  := "1GB";
        PCS_SAMP_16B    : string  := "X20";
        PCS_FARLP_PWR_REDUCTION: string  := "FALSE";
        PCS_COMMA_REG0  : integer := 0;
        PCS_COMMA_MASK  : integer := 0;
        PCS_CEB_MODE    : string  := "10GB";
        PCS_CTC_MODE    : string  := "1SKIP";
        PCS_A_REG       : integer := 0;
        PCS_GE_AUTO_EN  : string  := "FALSE";
        PCS_SKIP_REG0   : integer := 0;
        PCS_SKIP_REG1   : integer := 0;
        PCS_SKIP_REG2   : integer := 0;
        PCS_SKIP_REG3   : integer := 0;
        PCS_DEC_DUAL    : string  := "FALSE";
        PCS_SPLIT       : string  := "FALSE";
        PCS_FIFOFLAG_CTC: string  := "FALSE";
        PCS_COMMA_DET_MODE: string  := "COMMA_PATTERN";
        PCS_ERRDETECT_SILENCE: string  := "FALSE";
        PCS_PMA_RCLK_POLINV: string  := "PMA_RCLK";
        PCS_PCS_RCLK_SEL: string  := "PMA_RCLK";
        PCS_CB_RCLK_SEL : string  := "PMA_RCLK";
        PCS_AFTER_CTC_RCLK_SEL: string  := "PMA_RCLK";
        PCS_RCLK_POLINV : string  := "RCLK";
        PCS_BRIDGE_RCLK_SEL: string  := "PMA_RCLK";
        PCS_PCS_RCLK_EN : string  := "FALSE";
        PCS_CB_RCLK_EN  : string  := "FALSE";
        PCS_AFTER_CTC_RCLK_EN: string  := "FALSE";
        PCS_AFTER_CTC_RCLK_EN_GB: string  := "FALSE";
        PCS_PCS_RX_RSTN : string  := "FALSE";
        PCS_PCIE_SLAVE  : string  := "MASTER";
        PCS_RX_64B66B_67B: string  := "NORMAL";
        PCS_RX_BRIDGE_CLK_POLINV: string  := "RX_BRIDGE_CLK";
        PCS_PCS_CB_RSTN : string  := "FALSE";
        PCS_TX_BRIDGE_GEAR_SEL: string  := "FALSE";
        PCS_TX_BYPASS_BRIDGE_UINT: string  := "FALSE";
        PCS_TX_BYPASS_BRIDGE_FIFO: string  := "FALSE";
        PCS_TX_BYPASS_GEAR: string  := "FALSE";
        PCS_TX_BYPASS_ENC: string  := "FALSE";
        PCS_TX_BYPASS_BIT_SLIP: string  := "FALSE";
        PCS_TX_GEAR_SPLIT: string  := "FALSE";
        PCS_TX_DRIVE_REG_MODE: string  := "NO_CHANGE";
        PCS_TX_BIT_SLIP_CYCLES: integer := 0;
        PCS_INT_TX_MASK_0: string  := "FALSE";
        PCS_INT_TX_MASK_1: string  := "FALSE";
        PCS_INT_TX_MASK_2: string  := "FALSE";
        PCS_INT_TX_CLR_0: string  := "FALSE";
        PCS_INT_TX_CLR_1: string  := "FALSE";
        PCS_INT_TX_CLR_2: string  := "FALSE";
        PCS_TX_PMA_TCLK_POLINV: string  := "PMA_TCLK";
        PCS_TX_PCS_CLK_EN_SEL: string  := "FALSE";
        PCS_TX_BRIDGE_TCLK_SEL: string  := "TCLK";
        PCS_TX_TCLK_POLINV: string  := "TCLK";
        PCS_PCS_TCLK_SEL: string  := "PMA_TCLK";
        PCS_TX_PCS_TX_RSTN: string  := "FALSE";
        PCS_TX_SLAVE    : string  := "MASTER";
        PCS_TX_GEAR_CLK_EN_SEL: string  := "FALSE";
        PCS_DATA_WIDTH_MODE: string  := "X20";
        PCS_TX_64B66B_67B: string  := "NORMAL";
        PCS_GEAR_TCLK_SEL: string  := "PMA_TCLK";
        PCS_TX_TCLK2FABRIC_SEL: string  := "FALSE";
        PCS_TX_OUTZZ    : string  := "FALSE";
        PCS_ENC_DUAL    : string  := "FALSE";
        PCS_TX_BITSLIP_DATA_MODE: string  := "X10";
        PCS_TX_BRIDGE_CLK_POLINV: string  := "TX_BRIDGE_CLK";
        PCS_COMMA_REG1  : integer := 0;
        PCS_RAPID_IMAX  : integer := 0;
        PCS_RAPID_VMIN_1: integer := 0;
        PCS_RAPID_VMIN_2: integer := 0;
        PCS_RX_PRBS_MODE: string  := "DISABLE";
        PCS_RX_ERRCNT_CLR: string  := "FALSE";
        PCS_PRBS_ERR_LPBK: string  := "FALSE";
        PCS_TX_PRBS_MODE: string  := "DISABLE";
        PCS_TX_INSERT_ER: string  := "FALSE";
        PCS_ENABLE_PRBS_GEN: string  := "FALSE";
        PCS_DEFAULT_RADDR: integer := 0;
        PCS_MASTER_CHECK_OFFSET: integer := 0;
        PCS_DELAY_SET   : integer := 0;
        PCS_SEACH_OFFSET: string  := "20BIT";
        PCS_CEB_RAPIDLS_MMAX: integer := 0;
        PCS_CTC_AFULL   : integer := 20;
        PCS_CTC_AEMPTY  : integer := 12;
        PCS_CTC_CONTI_SKP_SET: integer := 0;
        PCS_FAR_LOOP    : string  := "FALSE";
        PCS_NEAR_LOOP   : string  := "FALSE";
        PCS_PMA_TX2RX_PLOOP_EN: string  := "FALSE";
        PCS_PMA_TX2RX_SLOOP_EN: string  := "FALSE";
        PCS_PMA_RX2TX_PLOOP_EN: string  := "FALSE";
        PCS_INT_RX_MASK_0: string  := "FALSE";
        PCS_INT_RX_MASK_1: string  := "FALSE";
        PCS_INT_RX_MASK_2: string  := "FALSE";
        PCS_INT_RX_MASK_3: string  := "FALSE";
        PCS_INT_RX_MASK_4: string  := "FALSE";
        PCS_INT_RX_MASK_5: string  := "FALSE";
        PCS_INT_RX_MASK_6: string  := "FALSE";
        PCS_INT_RX_MASK_7: string  := "FALSE";
        PCS_INT_RX_CLR_0: string  := "FALSE";
        PCS_INT_RX_CLR_1: string  := "FALSE";
        PCS_INT_RX_CLR_2: string  := "FALSE";
        PCS_INT_RX_CLR_3: string  := "FALSE";
        PCS_INT_RX_CLR_4: string  := "FALSE";
        PCS_INT_RX_CLR_5: string  := "FALSE";
        PCS_INT_RX_CLR_6: string  := "FALSE";
        PCS_INT_RX_CLR_7: string  := "FALSE";
        PCS_CA_RSTN_RX  : string  := "FALSE";
        PCS_CA_DYN_DLY_EN_RX: string  := "FALSE";
        PCS_CA_DYN_DLY_SEL_RX: string  := "FALSE";
        PCS_CA_RX       : integer := 0;
        PCS_CA_RSTN_TX  : string  := "FALSE";
        PCS_CA_DYN_DLY_EN_TX: string  := "FALSE";
        PCS_CA_DYN_DLY_SEL_TX: string  := "FALSE";
        PCS_CA_TX       : integer := 0;
        PCS_RXPRBS_PWR_REDUCTION: string  := "NORMAL";
        PCS_WDALIGN_PWR_REDUCTION: string  := "NORMAL";
        PCS_RXDEC_PWR_REDUCTION: string  := "NORMAL";
        PCS_RXCB_PWR_REDUCTION: string  := "NORMAL";
        PCS_RXCTC_PWR_REDUCTION: string  := "NORMAL";
        PCS_RXGEAR_PWR_REDUCTION: string  := "NORMAL";
        PCS_RXBRG_PWR_REDUCTION: string  := "NORMAL";
        PCS_RXTEST_PWR_REDUCTION: string  := "NORMAL";
        PCS_TXBRG_PWR_REDUCTION: string  := "NORMAL";
        PCS_TXGEAR_PWR_REDUCTION: string  := "NORMAL";
        PCS_TXENC_PWR_REDUCTION: string  := "NORMAL";
        PCS_TXBSLP_PWR_REDUCTION: string  := "NORMAL";
        PCS_TXPRBS_PWR_REDUCTION: string  := "NORMAL";
        PMA_REG_RX_PD   : string  := "ON";
        PMA_REG_RX_PD_EN: string  := "FALSE";
        PMA_REG_RX_RESERVED_2: string  := "FALSE";
        PMA_REG_RX_RESERVED_3: string  := "FALSE";
        PMA_REG_RX_DATAPATH_PD: string  := "ON";
        PMA_REG_RX_DATAPATH_PD_EN: string  := "FALSE";
        PMA_REG_RX_SIGDET_PD: string  := "ON";
        PMA_REG_RX_SIGDET_PD_EN: string  := "FALSE";
        PMA_REG_RX_DCC_RST_N: string  := "TRUE";
        PMA_REG_RX_DCC_RST_N_EN: string  := "FALSE";
        PMA_REG_RX_CDR_RST_N: string  := "TRUE";
        PMA_REG_RX_CDR_RST_N_EN: string  := "FALSE";
        PMA_REG_RX_SIGDET_RST_N: string  := "TRUE";
        PMA_REG_RX_SIGDET_RST_N_EN: string  := "FALSE";
        PMA_REG_RXPCLK_SLIP: string  := "FALSE";
        PMA_REG_RXPCLK_SLIP_OW: string  := "FALSE";
        PMA_REG_RX_PCLKSWITCH_RST_N: string  := "TRUE";
        PMA_REG_RX_PCLKSWITCH_RST_N_EN: string  := "FALSE";
        PMA_REG_RX_PCLKSWITCH: string  := "FALSE";
        PMA_REG_RX_PCLKSWITCH_EN: string  := "FALSE";
        PMA_REG_RX_HIGHZ: string  := "FALSE";
        PMA_REG_RX_HIGHZ_EN: string  := "FALSE";
        PMA_REG_RX_SIGDET_CLK_WINDOW: string  := "FALSE";
        PMA_REG_RX_SIGDET_CLK_WINDOW_OW: string  := "FALSE";
        PMA_REG_RX_PD_BIAS_RX: string  := "FALSE";
        PMA_REG_RX_PD_BIAS_RX_OW: string  := "FALSE";
        PMA_REG_RX_RESET_N: string  := "FALSE";
        PMA_REG_RX_RESET_N_OW: string  := "FALSE";
        PMA_REG_RX_RESERVED_29_28: integer := 0;
        PMA_REG_RX_BUSWIDTH: string  := "20BIT";
        PMA_REG_RX_BUSWIDTH_EN: string  := "FALSE";
        PMA_REG_RX_RATE : string  := "DIV1";
        PMA_REG_RX_RESERVED_36: string  := "FALSE";
        PMA_REG_RX_RATE_EN: string  := "FALSE";
        PMA_REG_RX_RES_TRIM: integer := 46;
        PMA_REG_RX_RESERVED_44: string  := "FALSE";
        PMA_REG_RX_RESERVED_45: string  := "FALSE";
        PMA_REG_RX_SIGDET_STATUS_EN: string  := "FALSE";
        PMA_REG_RX_RESERVED_48_47: integer := 0;
        PMA_REG_RX_ICTRL_SIGDET: integer := 5;
        PMA_REG_CDR_READY_THD: integer := 2734;
        PMA_REG_RX_RESERVED_65: string  := "FALSE";
        PMA_REG_RX_PCLK_EDGE_SEL: string  := "POS_EDGE";
        PMA_REG_RX_PIBUF_IC: integer := 1;
        PMA_REG_RX_RESERVED_69: string  := "FALSE";
        PMA_REG_RX_DCC_IC_RX: integer := 1;
        PMA_REG_CDR_READY_CHECK_CTRL: integer := 0;
        PMA_REG_RX_ICTRL_TRX: string  := "100PCT";
        PMA_REG_RX_RESERVED_77_76: integer := 0;
        PMA_REG_RX_RESERVED_79_78: integer := 1;
        PMA_REG_RX_RESERVED_81_80: integer := 1;
        PMA_REG_RX_ICTRL_PIBUF: string  := "100PCT";
        PMA_REG_RX_ICTRL_PI: string  := "100PCT";
        PMA_REG_RX_ICTRL_DCC: string  := "100PCT";
        PMA_REG_RX_RESERVED_89_88: integer := 1;
        PMA_REG_TX_RATE : string  := "DIV1";
        PMA_REG_RX_RESERVED_92: string  := "FALSE";
        PMA_REG_TX_RATE_EN: string  := "FALSE";
        PMA_REG_RX_TX2RX_PLPBK_RST_N: string  := "TRUE";
        PMA_REG_RX_TX2RX_PLPBK_RST_N_EN: string  := "FALSE";
        PMA_REG_RX_TX2RX_PLPBK_EN: string  := "FALSE";
        PMA_REG_TXCLK_SEL: string  := "PLL";
        PMA_REG_RX_DATA_POLARITY: string  := "NORMAL";
        PMA_REG_RX_ERR_INSERT: string  := "FALSE";
        PMA_REG_UDP_CHK_EN: string  := "FALSE";
        PMA_REG_PRBS_SEL: string  := "PRBS7";
        PMA_REG_PRBS_CHK_EN: string  := "FALSE";
        PMA_REG_PRBS_CHK_WIDTH_SEL: string  := "20BIT";
        PMA_REG_BIST_CHK_PAT_SEL: string  := "PRBS";
        PMA_REG_LOAD_ERR_CNT: string  := "FALSE";
        PMA_REG_CHK_COUNTER_EN: string  := "FALSE";
        PMA_REG_CDR_PROP_GAIN: integer := 7;
        PMA_REG_CDR_PROP_TURBO_GAIN: integer := 5;
        PMA_REG_CDR_INT_GAIN: integer := 7;
        PMA_REG_CDR_INT_TURBO_GAIN: integer := 5;
        PMA_REG_CDR_INT_SAT_MAX: integer := 768;
        PMA_REG_CDR_INT_SAT_MIN: integer := 255;
        PMA_REG_CDR_INT_RST: string  := "FALSE";
        PMA_REG_CDR_INT_RST_OW: string  := "FALSE";
        PMA_REG_CDR_PROP_RST: string  := "FALSE";
        PMA_REG_CDR_PROP_RST_OW: string  := "FALSE";
        PMA_REG_CDR_LOCK_RST: string  := "FALSE";
        PMA_REG_CDR_LOCK_RST_OW: string  := "FALSE";
        PMA_REG_CDR_RX_PI_FORCE_SEL: integer := 0;
        PMA_REG_CDR_RX_PI_FORCE_D: integer := 0;
        PMA_REG_CDR_LOCK_TIMER: string  := "1_2U";
        PMA_REG_CDR_TURBO_MODE_TIMER: integer := 1;
        PMA_REG_CDR_LOCK_VAL: string  := "FALSE";
        PMA_REG_CDR_LOCK_OW: string  := "FALSE";
        PMA_REG_CDR_INT_SAT_DET_EN: string  := "TRUE";
        PMA_REG_CDR_SAT_AUTO_DIS: string  := "TRUE";
        PMA_REG_CDR_GAIN_AUTO: string  := "FALSE";
        PMA_REG_CDR_TURBO_GAIN_AUTO: string  := "FALSE";
        PMA_REG_RX_RESERVED_171_167: integer := 0;
        PMA_REG_RX_RESERVED_175_172: integer := 0;
        PMA_REG_CDR_SAT_DET_STATUS_EN: string  := "FALSE";
        PMA_REG_CDR_SAT_DET_STATUS_RESET_EN: string  := "FALSE";
        PMA_REG_CDR_PI_CTRL_RST: string  := "FALSE";
        PMA_REG_CDR_PI_CTRL_RST_OW: string  := "FALSE";
        PMA_REG_CDR_SAT_DET_RST: string  := "FALSE";
        PMA_REG_CDR_SAT_DET_RST_OW: string  := "FALSE";
        PMA_REG_CDR_SAT_DET_STICKY_RST: string  := "FALSE";
        PMA_REG_CDR_SAT_DET_STICKY_RST_OW: string  := "FALSE";
        PMA_REG_CDR_SIGDET_STATUS_DIS: string  := "FALSE";
        PMA_REG_CDR_SAT_DET_TIMER: integer := 2;
        PMA_REG_CDR_SAT_DET_STATUS_VAL: string  := "FALSE";
        PMA_REG_CDR_SAT_DET_STATUS_OW: string  := "FALSE";
        PMA_REG_CDR_TURBO_MODE_EN: string  := "TRUE";
        PMA_REG_RX_RESERVED_190: string  := "FALSE";
        PMA_REG_RX_RESERVED_193_191: integer := 0;
        PMA_REG_CDR_STATUS_FIFO_EN: string  := "TRUE";
        PMA_REG_PMA_TEST_SEL: integer := 0;
        PMA_REG_OOB_COMWAKE_GAP_MIN: integer := 3;
        PMA_REG_OOB_COMWAKE_GAP_MAX: integer := 11;
        PMA_REG_OOB_COMINIT_GAP_MIN: integer := 15;
        PMA_REG_OOB_COMINIT_GAP_MAX: integer := 35;
        PMA_REG_RX_RESERVED_227_226: integer := 1;
        PMA_REG_COMWAKE_STATUS_CLEAR: integer := 0;
        PMA_REG_COMINIT_STATUS_CLEAR: integer := 0;
        PMA_REG_RX_SYNC_RST_N_EN: string  := "FALSE";
        PMA_REG_RX_SYNC_RST_N: string  := "TRUE";
        PMA_REG_RX_RESERVED_233_232: integer := 0;
        PMA_REG_RX_RESERVED_235_234: integer := 0;
        PMA_REG_RX_SATA_COMINIT_OW: string  := "FALSE";
        PMA_REG_RX_SATA_COMINIT: string  := "FALSE";
        PMA_REG_RX_SATA_COMWAKE_OW: string  := "FALSE";
        PMA_REG_RX_SATA_COMWAKE: string  := "FALSE";
        PMA_REG_RX_RESERVED_241_240: integer := 0;
        PMA_REG_RX_DCC_DISABLE: string  := "FALSE";
        PMA_REG_RX_RESERVED_243: string  := "FALSE";
        PMA_REG_RX_SLIP_SEL_EN: string  := "FALSE";
        PMA_REG_RX_SLIP_SEL: integer := 0;
        PMA_REG_RX_SLIP_EN: string  := "FALSE";
        PMA_REG_RX_SIGDET_STATUS_SEL: integer := 5;
        PMA_REG_RX_SIGDET_FSM_RST_N: string  := "TRUE";
        PMA_REG_RX_RESERVED_254: string  := "FALSE";
        PMA_REG_RX_SIGDET_STATUS: string  := "FALSE";
        PMA_REG_RX_SIGDET_VTH: string  := "27MV";
        PMA_REG_RX_SIGDET_GRM: integer := 0;
        PMA_REG_RX_SIGDET_PULSE_EXT: string  := "FALSE";
        PMA_REG_RX_SIGDET_CH2_SEL: integer := 0;
        PMA_REG_RX_SIGDET_CH2_CHK_WINDOW: integer := 3;
        PMA_REG_RX_SIGDET_CHK_WINDOW_EN: string  := "TRUE";
        PMA_REG_RX_SIGDET_NOSIG_COUNT_SETTING: integer := 4;
        PMA_REG_SLIP_FIFO_INV_EN: string  := "FALSE";
        PMA_REG_SLIP_FIFO_INV: string  := "POS_EDGE";
        PMA_REG_RX_SIGDET_OOB_DET_COUNT_VAL: integer := 0;
        PMA_REG_RX_SIGDET_4OOB_DET_SEL: integer := 7;
        PMA_REG_RX_RESERVED_285_283: integer := 0;
        PMA_REG_RX_RESERVED_286: string  := "FALSE";
        PMA_REG_RX_SIGDET_IC_I: integer := 10;
        PMA_REG_RX_OOB_DETECTOR_RESET_N_OW: string  := "FALSE";
        PMA_REG_RX_OOB_DETECTOR_RESET_N: string  := "FALSE";
        PMA_REG_RX_OOB_DETECTOR_PD_OW: string  := "FALSE";
        PMA_REG_RX_OOB_DETECTOR_PD: string  := "ON";
        PMA_REG_RX_LS_MODE_EN: string  := "FALSE";
        PMA_REG_ANA_RX_EQ1_R_SET_FB_O_SEL: string  := "FALSE";
        PMA_REG_ANA_RX_EQ2_R_SET_FB_O_SEL: string  := "FALSE";
        PMA_REG_RX_EQ1_R_SET_TOP: integer := 0;
        PMA_REG_RX_EQ1_R_SET_FB: integer := 0;
        PMA_REG_RX_EQ1_C_SET_FB: integer := 0;
        PMA_REG_RX_EQ1_OFF: string  := "FALSE";
        PMA_REG_RX_EQ2_R_SET_TOP: integer := 0;
        PMA_REG_RX_EQ2_R_SET_FB: integer := 0;
        PMA_REG_RX_EQ2_C_SET_FB: integer := 0;
        PMA_REG_RX_EQ2_OFF: string  := "FALSE";
        PMA_REG_EQ_DAC  : integer := 0;
        PMA_REG_RX_ICTRL_EQ: integer := 2;
        PMA_REG_EQ_DC_CALIB_EN: string  := "FALSE";
        PMA_REG_EQ_DC_CALIB_SEL: string  := "FALSE";
        PMA_REG_RX_RESERVED_337_330: integer := 0;
        PMA_REG_RX_RESERVED_345_338: integer := 0;
        PMA_REG_RX_RESERVED_353_346: integer := 0;
        PMA_REG_RX_RESERVED_361_354: integer := 0;
        PMA_CTLE_CTRL_REG_I: integer := 0;
        PMA_CTLE_REG_FORCE_SEL_I: string  := "FALSE";
        PMA_CTLE_REG_HOLD_I: string  := "FALSE";
        PMA_CTLE_REG_INIT_DAC_I: integer := 0;
        PMA_CTLE_REG_POLARITY_I: string  := "FALSE";
        PMA_CTLE_REG_SHIFTER_GAIN_I: integer := 0;
        PMA_CTLE_REG_THRESHOLD_I: integer := 0;
        PMA_REG_RX_RES_TRIM_EN: string  := "FALSE";
        PMA_REG_RX_RESERVED_393_389: integer := 0;
        PMA_CFG_RX_LANE_POWERUP: string  := "OFF";
        PMA_CFG_RX_PMA_RSTN: string  := "FALSE";
        PMA_INT_PMA_RX_MASK_0: string  := "FALSE";
        PMA_INT_PMA_RX_CLR_0: string  := "FALSE";
        PMA_CFG_CTLE_ADP_RSTN: string  := "TRUE";
        PMA_REG_TX_PD   : string  := "ON";
        PMA_REG_TX_PD_OW: string  := "TRUE";
        PMA_REG_TX_MAIN_PRE_Z: string  := "FALSE";
        PMA_REG_TX_MAIN_PRE_Z_OW: string  := "FALSE";
        PMA_REG_TX_BEACON_TIMER_SEL: integer := 0;
        PMA_REG_TX_RXDET_REQ_OW: string  := "FALSE";
        PMA_REG_TX_RXDET_REQ: string  := "FALSE";
        PMA_REG_TX_BEACON_EN_OW: string  := "FALSE";
        PMA_REG_TX_BEACON_EN: string  := "FALSE";
        PMA_REG_TX_EI_EN_OW: string  := "FALSE";
        PMA_REG_TX_EI_EN: string  := "FALSE";
        PMA_REG_TX_BIT_CONV: string  := "FALSE";
        PMA_REG_TX_RES_CAL: integer := 50;
        PMA_REG_TX_RESERVED_19: string  := "FALSE";
        PMA_REG_TX_RESERVED_25_20: integer := 32;
        PMA_REG_TX_RESERVED_33_26: integer := 0;
        PMA_REG_TX_RESERVED_41_34: integer := 0;
        PMA_REG_TX_RESERVED_49_42: integer := 0;
        PMA_REG_TX_RESERVED_57_50: integer := 0;
        PMA_REG_TX_SYNC_OW: string  := "FALSE";
        PMA_REG_TX_SYNC : string  := "FALSE";
        PMA_REG_TX_PD_POST: string  := "OFF";
        PMA_REG_TX_PD_POST_OW: string  := "TRUE";
        PMA_REG_TX_RESET_N_OW: string  := "FALSE";
        PMA_REG_TX_RESET_N: string  := "TRUE";
        PMA_REG_TX_RESERVED_64: string  := "FALSE";
        PMA_REG_TX_RESERVED_65: string  := "TRUE";
        PMA_REG_TX_BUSWIDTH_OW: string  := "FALSE";
        PMA_REG_TX_BUSWIDTH: string  := "20BIT";
        PMA_REG_PLL_READY_OW: string  := "FALSE";
        PMA_REG_PLL_READY: string  := "TRUE";
        PMA_REG_TX_RESERVED_72: string  := "FALSE";
        PMA_REG_TX_RESERVED_73: string  := "FALSE";
        PMA_REG_TX_RESERVED_74: string  := "FALSE";
        PMA_REG_EI_PCLK_DELAY_SEL: integer := 0;
        PMA_REG_TX_RESERVED_77: string  := "FALSE";
        PMA_REG_TX_RESERVED_83_78: integer := 0;
        PMA_REG_TX_RESERVED_89_84: integer := 0;
        PMA_REG_TX_RESERVED_95_90: integer := 0;
        PMA_REG_TX_RESERVED_101_96: integer := 0;
        PMA_REG_TX_RESERVED_107_102: integer := 0;
        PMA_REG_TX_RESERVED_113_108: integer := 0;
        PMA_REG_TX_AMP_DAC0: integer := 25;
        PMA_REG_TX_AMP_DAC1: integer := 19;
        PMA_REG_TX_AMP_DAC2: integer := 14;
        PMA_REG_TX_AMP_DAC3: integer := 9;
        PMA_REG_TX_RESERVED_143_138: integer := 5;
        PMA_REG_TX_MARGIN: integer := 0;
        PMA_REG_TX_MARGIN_OW: string  := "FALSE";
        PMA_REG_TX_RESERVED_149_148: integer := 0;
        PMA_REG_TX_RESERVED_150: string  := "FALSE";
        PMA_REG_TX_SWING: string  := "FALSE";
        PMA_REG_TX_SWING_OW: string  := "FALSE";
        PMA_REG_TX_RESERVED_153: string  := "FALSE";
        PMA_REG_TX_RXDET_THRESHOLD: string  := "84MV";
        PMA_REG_TX_RESERVED_157_156: integer := 0;
        PMA_REG_TX_BEACON_OSC_CTRL: string  := "FALSE";
        PMA_REG_TX_RESERVED_160_159: integer := 0;
        PMA_REG_TX_RESERVED_162_161: integer := 0;
        PMA_REG_TX_TX2RX_SLPBACK_EN: string  := "FALSE";
        PMA_REG_TX_PCLK_EDGE_SEL: string  := "FALSE";
        PMA_REG_TX_RXDET_STATUS_OW: string  := "FALSE";
        PMA_REG_TX_RXDET_STATUS: string  := "TRUE";
        PMA_REG_TX_PRBS_GEN_EN: string  := "FALSE";
        PMA_REG_TX_PRBS_GEN_WIDTH_SEL: string  := "20BIT";
        PMA_REG_TX_PRBS_SEL: string  := "PRBS7";
        PMA_REG_TX_UDP_DATA_7_TO_0: integer := 5;
        PMA_REG_TX_UDP_DATA_15_TO_8: integer := 235;
        PMA_REG_TX_UDP_DATA_19_TO_16: integer := 3;
        PMA_REG_TX_RESERVED_192: string  := "FALSE";
        PMA_REG_TX_FIFO_WP_CTRL: integer := 4;
        PMA_REG_TX_FIFO_EN: string  := "FALSE";
        PMA_REG_TX_DATA_MUX_SEL: integer := 0;
        PMA_REG_TX_ERR_INSERT: string  := "FALSE";
        PMA_REG_TX_RESERVED_203_200: integer := 0;
        PMA_REG_TX_RESERVED_204: string  := "FALSE";
        PMA_REG_TX_SATA_EN: string  := "FALSE";
        PMA_REG_TX_RESERVED_207_206: integer := 0;
        PMA_REG_RATE_CHANGE_TXPCLK_ON_OW: string  := "FALSE";
        PMA_REG_RATE_CHANGE_TXPCLK_ON: string  := "TRUE";
        PMA_REG_TX_CFG_POST1: integer := 0;
        PMA_REG_TX_CFG_POST2: integer := 0;
        PMA_REG_TX_DEEMP: integer := 0;
        PMA_REG_TX_DEEMP_OW: string  := "FALSE";
        PMA_REG_TX_RESERVED_224_223: integer := 0;
        PMA_REG_TX_RESERVED_225: string  := "FALSE";
        PMA_REG_TX_RESERVED_229_226: integer := 0;
        PMA_REG_TX_OOB_DELAY_SEL: integer := 0;
        PMA_REG_TX_POLARITY: string  := "NORMAL";
        PMA_REG_ANA_TX_JTAG_DATA_O_SEL: string  := "FALSE";
        PMA_REG_TX_RESERVED_236: string  := "FALSE";
        PMA_REG_TX_LS_MODE_EN: string  := "FALSE";
        PMA_REG_TX_JTAG_MODE_EN_OW: string  := "FALSE";
        PMA_REG_TX_JTAG_MODE_EN: string  := "FALSE";
        PMA_REG_RX_JTAG_MODE_EN_OW: string  := "FALSE";
        PMA_REG_RX_JTAG_MODE_EN: string  := "FALSE";
        PMA_REG_RX_JTAG_OE: string  := "TRUE";
        PMA_REG_RX_ACJTAG_VHYSTSEL: integer := 0;
        PMA_REG_TX_RES_CAL_EN: string  := "FALSE";
        PMA_REG_RX_TERM_MODE_CTRL: integer := 4;
        PMA_REG_TX_RESERVED_251_250: integer := 0;
        PMA_REG_PLPBK_TXPCLK_EN: string  := "FALSE";
        PMA_REG_TX_RESERVED_253: string  := "FALSE";
        PMA_REG_TX_RESERVED_254: string  := "FALSE";
        PMA_REG_TX_RESERVED_255: string  := "FALSE";
        PMA_REG_TX_RESERVED_256: string  := "FALSE";
        PMA_REG_TX_RESERVED_257: string  := "FALSE";
        PMA_REG_TX_PH_SEL: integer := 1;
        PMA_REG_TX_CFG_PRE: integer := 0;
        PMA_REG_TX_CFG_MAIN: integer := 0;
        PMA_REG_CFG_POST: integer := 0;
        PMA_REG_PD_MAIN : string  := "TRUE";
        PMA_REG_PD_PRE  : string  := "TRUE";
        PMA_REG_TX_LS_DATA: string  := "FALSE";
        PMA_REG_TX_DCC_BUF_SZ_SEL: integer := 0;
        PMA_REG_TX_DCC_CAL_CUR_TUNE: integer := 0;
        PMA_REG_TX_DCC_CAL_EN: string  := "FALSE";
        PMA_REG_TX_DCC_CUR_SS: integer := 0;
        PMA_REG_TX_DCC_FA_CTRL: string  := "FALSE";
        PMA_REG_TX_DCC_RI_CTRL: string  := "FALSE";
        PMA_REG_ATB_SEL_2_TO_0: integer := 0;
        PMA_REG_ATB_SEL_9_TO_3: integer := 0;
        PMA_REG_TX_CFG_7_TO_0: integer := 0;
        PMA_REG_TX_CFG_15_TO_8: integer := 0;
        PMA_REG_TX_CFG_23_TO_16: integer := 0;
        PMA_REG_TX_CFG_31_TO_24: integer := 0;
        PMA_REG_TX_OOB_EI_EN: string  := "FALSE";
        PMA_REG_TX_OOB_EI_EN_OW: string  := "FALSE";
        PMA_REG_TX_BEACON_EN_DELAYED: string  := "FALSE";
        PMA_REG_TX_BEACON_EN_DELAYED_OW: string  := "FALSE";
        PMA_REG_TX_JTAG_DATA: string  := "FALSE";
        PMA_REG_TX_RXDET_TIMER_SEL: integer := 87;
        PMA_REG_TX_CFG1_7_0: integer := 0;
        PMA_REG_TX_CFG1_15_8: integer := 0;
        PMA_REG_TX_CFG1_23_16: integer := 0;
        PMA_REG_TX_CFG1_31_24: integer := 0;
        PMA_REG_CFG_LANE_POWERUP: string  := "OFF";
        PMA_REG_CFG_TX_LANE_POWERUP_CLKPATH: string  := "FALSE";
        PMA_REG_CFG_TX_LANE_POWERUP_PISO: string  := "FALSE";
        PMA_REG_CFG_TX_LANE_POWERUP_DRIVER: string  := "FALSE"
    );
    port(
        P_TX_SDN        : out    vl_logic;
        P_TX_SDP        : out    vl_logic;
        P_PCS_RX_MCB_STATUS: out    vl_logic;
        P_PCS_LSM_SYNCED: out    vl_logic;
        P_CFG_READY     : out    vl_logic;
        P_CFG_RDATA     : out    vl_logic_vector(7 downto 0);
        P_CFG_INT       : out    vl_logic;
        P_RDATA         : out    vl_logic_vector(46 downto 0);
        P_RCLK2FABRIC   : out    vl_logic;
        P_TCLK2FABRIC   : out    vl_logic;
        P_RX_SIGDET_STATUS: out    vl_logic;
        P_RX_SATA_COMINIT: out    vl_logic;
        P_RX_SATA_COMWAKE: out    vl_logic;
        P_RX_LS_DATA    : out    vl_logic;
        P_RX_READY      : out    vl_logic;
        P_TEST_STATUS   : out    vl_logic_vector(19 downto 0);
        P_TX_RXDET_STATUS: out    vl_logic;
        P_CA_ALIGN_RX   : out    vl_logic;
        P_CA_ALIGN_TX   : out    vl_logic;
        P_TEST_SO0      : out    vl_logic;
        P_TEST_SO1      : out    vl_logic;
        P_TEST_SO2      : out    vl_logic;
        P_TEST_SO3      : out    vl_logic;
        P_TEST_SO4      : out    vl_logic;
        P_FOR_PMA_TEST_SO: out    vl_logic_vector(1 downto 0);
        PMA_RCLK        : out    vl_logic;
        LANE_COUT_BUS_FORWARD: out    vl_logic_vector(18 downto 0);
        APATTERN_STATUS_COUT: out    vl_logic;
        TXPCLK_PLL      : out    vl_logic;
        P_RX_SDN        : in     vl_logic;
        P_RX_SDP        : in     vl_logic;
        P_RX_CLK_FR_CORE: in     vl_logic;
        P_RCLK2_FR_CORE : in     vl_logic;
        P_TX_CLK_FR_CORE: in     vl_logic;
        P_TCLK2_FR_CORE : in     vl_logic;
        P_PCS_TX_RST    : in     vl_logic;
        P_PCS_RX_RST    : in     vl_logic;
        P_PCS_CB_RST    : in     vl_logic;
        P_RXGEAR_SLIP   : in     vl_logic;
        P_CFG_CLK       : in     vl_logic;
        P_CFG_RST       : in     vl_logic;
        P_CFG_PSEL      : in     vl_logic;
        P_CFG_ENABLE    : in     vl_logic;
        P_CFG_WRITE     : in     vl_logic;
        P_CFG_ADDR      : in     vl_logic_vector(11 downto 0);
        P_CFG_WDATA     : in     vl_logic_vector(7 downto 0);
        P_TDATA         : in     vl_logic_vector(45 downto 0);
        P_PCS_WORD_ALIGN_EN: in     vl_logic;
        P_RX_POLARITY_INVERT: in     vl_logic;
        P_CEB_ADETECT_EN: in     vl_logic;
        P_PCS_MCB_EXT_EN: in     vl_logic;
        P_PCS_NEAREND_LOOP: in     vl_logic;
        P_PCS_FAREND_LOOP: in     vl_logic;
        P_PMA_NEAREND_PLOOP: in     vl_logic;
        P_PMA_NEAREND_SLOOP: in     vl_logic;
        P_PMA_FAREND_PLOOP: in     vl_logic;
        P_LANE_PD       : in     vl_logic;
        P_LANE_RST      : in     vl_logic;
        P_RX_LANE_PD    : in     vl_logic;
        P_RX_PMA_RST    : in     vl_logic;
        P_CTLE_ADP_RST  : in     vl_logic;
        P_TX_DEEMP      : in     vl_logic_vector(1 downto 0);
        P_TX_LS_DATA    : in     vl_logic;
        P_TX_BEACON_EN  : in     vl_logic;
        P_TX_SWING      : in     vl_logic;
        P_TX_RXDET_REQ  : in     vl_logic;
        P_TX_RATE       : in     vl_logic_vector(2 downto 0);
        P_TX_BUSWIDTH   : in     vl_logic_vector(2 downto 0);
        P_TX_MARGIN     : in     vl_logic_vector(2 downto 0);
        P_TX_PMA_RST    : in     vl_logic;
        P_TX_LANE_PD_CLKPATH: in     vl_logic;
        P_TX_LANE_PD_PISO: in     vl_logic;
        P_TX_LANE_PD_DRIVER: in     vl_logic;
        P_RX_RATE       : in     vl_logic_vector(2 downto 0);
        P_RX_BUSWIDTH   : in     vl_logic_vector(2 downto 0);
        P_RX_HIGHZ      : in     vl_logic;
        P_CIM_CLK_ALIGNER_RX: in     vl_logic_vector(7 downto 0);
        P_CIM_CLK_ALIGNER_TX: in     vl_logic_vector(7 downto 0);
        P_CIM_DYN_DLY_SEL_RX: in     vl_logic;
        P_CIM_DYN_DLY_SEL_TX: in     vl_logic;
        P_CIM_START_ALIGN_RX: in     vl_logic;
        P_CIM_START_ALIGN_TX: in     vl_logic;
        P_TEST_SE_N     : in     vl_logic;
        P_TEST_MODE_N   : in     vl_logic;
        P_TEST_RSTN     : in     vl_logic;
        P_TEST_SI0      : in     vl_logic;
        P_TEST_SI1      : in     vl_logic;
        P_TEST_SI2      : in     vl_logic;
        P_TEST_SI3      : in     vl_logic;
        P_TEST_SI4      : in     vl_logic;
        P_FOR_PMA_TEST_MODE_N: in     vl_logic;
        P_FOR_PMA_TEST_SE_N: in     vl_logic_vector(1 downto 0);
        P_FOR_PMA_TEST_CLK: in     vl_logic_vector(1 downto 0);
        P_FOR_PMA_TEST_RSTN: in     vl_logic_vector(1 downto 0);
        P_FOR_PMA_TEST_SI: in     vl_logic_vector(1 downto 0);
        MCB_RCLK        : in     vl_logic;
        SYNC            : in     vl_logic;
        RATE_CHANGE     : in     vl_logic;
        PLL_LOCK_SEL    : in     vl_logic;
        LANE_CIN_BUS_FORWARD: in     vl_logic_vector(18 downto 0);
        APATTERN_STATUS_CIN: in     vl_logic;
        CLK_TXP         : in     vl_logic;
        CLK_TXN         : in     vl_logic;
        CLK_RX0         : in     vl_logic;
        CLK_RX90        : in     vl_logic;
        CLK_RX180       : in     vl_logic;
        CLK_RX270       : in     vl_logic;
        PLL_PD_I        : in     vl_logic;
        PLL_RESET_I     : in     vl_logic;
        PLL_REFCLK_I    : in     vl_logic;
        PLL_RES_TRIM_I  : in     vl_logic_vector(5 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of MUX_BIAS : constant is 2;
    attribute mti_svvh_generic_type of PD_CLK : constant is 2;
    attribute mti_svvh_generic_type of REG_SYNC : constant is 2;
    attribute mti_svvh_generic_type of REG_SYNC_OW : constant is 2;
    attribute mti_svvh_generic_type of PLL_LOCK_OW : constant is 2;
    attribute mti_svvh_generic_type of PLL_LOCK_OW_EN : constant is 2;
    attribute mti_svvh_generic_type of PCS_SLAVE : constant is 2;
    attribute mti_svvh_generic_type of PCS_BYPASS_WORD_ALIGN : constant is 1;
    attribute mti_svvh_generic_type of PCS_BYPASS_DENC : constant is 1;
    attribute mti_svvh_generic_type of PCS_BYPASS_BONDING : constant is 1;
    attribute mti_svvh_generic_type of PCS_BYPASS_CTC : constant is 1;
    attribute mti_svvh_generic_type of PCS_BYPASS_GEAR : constant is 1;
    attribute mti_svvh_generic_type of PCS_BYPASS_BRIDGE : constant is 1;
    attribute mti_svvh_generic_type of PCS_BYPASS_BRIDGE_FIFO : constant is 1;
    attribute mti_svvh_generic_type of PCS_DATA_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_RX_POLARITY_INV : constant is 1;
    attribute mti_svvh_generic_type of PCS_ALIGN_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_SAMP_16B : constant is 1;
    attribute mti_svvh_generic_type of PCS_FARLP_PWR_REDUCTION : constant is 1;
    attribute mti_svvh_generic_type of PCS_COMMA_REG0 : constant is 2;
    attribute mti_svvh_generic_type of PCS_COMMA_MASK : constant is 2;
    attribute mti_svvh_generic_type of PCS_CEB_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CTC_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_A_REG : constant is 2;
    attribute mti_svvh_generic_type of PCS_GE_AUTO_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_SKIP_REG0 : constant is 2;
    attribute mti_svvh_generic_type of PCS_SKIP_REG1 : constant is 2;
    attribute mti_svvh_generic_type of PCS_SKIP_REG2 : constant is 2;
    attribute mti_svvh_generic_type of PCS_SKIP_REG3 : constant is 2;
    attribute mti_svvh_generic_type of PCS_DEC_DUAL : constant is 1;
    attribute mti_svvh_generic_type of PCS_SPLIT : constant is 1;
    attribute mti_svvh_generic_type of PCS_FIFOFLAG_CTC : constant is 1;
    attribute mti_svvh_generic_type of PCS_COMMA_DET_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_ERRDETECT_SILENCE : constant is 1;
    attribute mti_svvh_generic_type of PCS_PMA_RCLK_POLINV : constant is 1;
    attribute mti_svvh_generic_type of PCS_PCS_RCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CB_RCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_AFTER_CTC_RCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_RCLK_POLINV : constant is 1;
    attribute mti_svvh_generic_type of PCS_BRIDGE_RCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_PCS_RCLK_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CB_RCLK_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_AFTER_CTC_RCLK_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_AFTER_CTC_RCLK_EN_GB : constant is 1;
    attribute mti_svvh_generic_type of PCS_PCS_RX_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PCS_PCIE_SLAVE : constant is 1;
    attribute mti_svvh_generic_type of PCS_RX_64B66B_67B : constant is 1;
    attribute mti_svvh_generic_type of PCS_RX_BRIDGE_CLK_POLINV : constant is 1;
    attribute mti_svvh_generic_type of PCS_PCS_CB_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PCS_TX_BRIDGE_GEAR_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_TX_BYPASS_BRIDGE_UINT : constant is 1;
    attribute mti_svvh_generic_type of PCS_TX_BYPASS_BRIDGE_FIFO : constant is 1;
    attribute mti_svvh_generic_type of PCS_TX_BYPASS_GEAR : constant is 1;
    attribute mti_svvh_generic_type of PCS_TX_BYPASS_ENC : constant is 1;
    attribute mti_svvh_generic_type of PCS_TX_BYPASS_BIT_SLIP : constant is 1;
    attribute mti_svvh_generic_type of PCS_TX_GEAR_SPLIT : constant is 1;
    attribute mti_svvh_generic_type of PCS_TX_DRIVE_REG_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_TX_BIT_SLIP_CYCLES : constant is 2;
    attribute mti_svvh_generic_type of PCS_INT_TX_MASK_0 : constant is 1;
    attribute mti_svvh_generic_type of PCS_INT_TX_MASK_1 : constant is 1;
    attribute mti_svvh_generic_type of PCS_INT_TX_MASK_2 : constant is 1;
    attribute mti_svvh_generic_type of PCS_INT_TX_CLR_0 : constant is 1;
    attribute mti_svvh_generic_type of PCS_INT_TX_CLR_1 : constant is 1;
    attribute mti_svvh_generic_type of PCS_INT_TX_CLR_2 : constant is 1;
    attribute mti_svvh_generic_type of PCS_TX_PMA_TCLK_POLINV : constant is 1;
    attribute mti_svvh_generic_type of PCS_TX_PCS_CLK_EN_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_TX_BRIDGE_TCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_TX_TCLK_POLINV : constant is 1;
    attribute mti_svvh_generic_type of PCS_PCS_TCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_TX_PCS_TX_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PCS_TX_SLAVE : constant is 1;
    attribute mti_svvh_generic_type of PCS_TX_GEAR_CLK_EN_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_DATA_WIDTH_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_TX_64B66B_67B : constant is 1;
    attribute mti_svvh_generic_type of PCS_GEAR_TCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_TX_TCLK2FABRIC_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_TX_OUTZZ : constant is 1;
    attribute mti_svvh_generic_type of PCS_ENC_DUAL : constant is 1;
    attribute mti_svvh_generic_type of PCS_TX_BITSLIP_DATA_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_TX_BRIDGE_CLK_POLINV : constant is 1;
    attribute mti_svvh_generic_type of PCS_COMMA_REG1 : constant is 2;
    attribute mti_svvh_generic_type of PCS_RAPID_IMAX : constant is 2;
    attribute mti_svvh_generic_type of PCS_RAPID_VMIN_1 : constant is 2;
    attribute mti_svvh_generic_type of PCS_RAPID_VMIN_2 : constant is 2;
    attribute mti_svvh_generic_type of PCS_RX_PRBS_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_RX_ERRCNT_CLR : constant is 1;
    attribute mti_svvh_generic_type of PCS_PRBS_ERR_LPBK : constant is 1;
    attribute mti_svvh_generic_type of PCS_TX_PRBS_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_TX_INSERT_ER : constant is 1;
    attribute mti_svvh_generic_type of PCS_ENABLE_PRBS_GEN : constant is 1;
    attribute mti_svvh_generic_type of PCS_DEFAULT_RADDR : constant is 2;
    attribute mti_svvh_generic_type of PCS_MASTER_CHECK_OFFSET : constant is 2;
    attribute mti_svvh_generic_type of PCS_DELAY_SET : constant is 2;
    attribute mti_svvh_generic_type of PCS_SEACH_OFFSET : constant is 1;
    attribute mti_svvh_generic_type of PCS_CEB_RAPIDLS_MMAX : constant is 2;
    attribute mti_svvh_generic_type of PCS_CTC_AFULL : constant is 2;
    attribute mti_svvh_generic_type of PCS_CTC_AEMPTY : constant is 2;
    attribute mti_svvh_generic_type of PCS_CTC_CONTI_SKP_SET : constant is 2;
    attribute mti_svvh_generic_type of PCS_FAR_LOOP : constant is 1;
    attribute mti_svvh_generic_type of PCS_NEAR_LOOP : constant is 1;
    attribute mti_svvh_generic_type of PCS_PMA_TX2RX_PLOOP_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_PMA_TX2RX_SLOOP_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_PMA_RX2TX_PLOOP_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_INT_RX_MASK_0 : constant is 1;
    attribute mti_svvh_generic_type of PCS_INT_RX_MASK_1 : constant is 1;
    attribute mti_svvh_generic_type of PCS_INT_RX_MASK_2 : constant is 1;
    attribute mti_svvh_generic_type of PCS_INT_RX_MASK_3 : constant is 1;
    attribute mti_svvh_generic_type of PCS_INT_RX_MASK_4 : constant is 1;
    attribute mti_svvh_generic_type of PCS_INT_RX_MASK_5 : constant is 1;
    attribute mti_svvh_generic_type of PCS_INT_RX_MASK_6 : constant is 1;
    attribute mti_svvh_generic_type of PCS_INT_RX_MASK_7 : constant is 1;
    attribute mti_svvh_generic_type of PCS_INT_RX_CLR_0 : constant is 1;
    attribute mti_svvh_generic_type of PCS_INT_RX_CLR_1 : constant is 1;
    attribute mti_svvh_generic_type of PCS_INT_RX_CLR_2 : constant is 1;
    attribute mti_svvh_generic_type of PCS_INT_RX_CLR_3 : constant is 1;
    attribute mti_svvh_generic_type of PCS_INT_RX_CLR_4 : constant is 1;
    attribute mti_svvh_generic_type of PCS_INT_RX_CLR_5 : constant is 1;
    attribute mti_svvh_generic_type of PCS_INT_RX_CLR_6 : constant is 1;
    attribute mti_svvh_generic_type of PCS_INT_RX_CLR_7 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CA_RSTN_RX : constant is 1;
    attribute mti_svvh_generic_type of PCS_CA_DYN_DLY_EN_RX : constant is 1;
    attribute mti_svvh_generic_type of PCS_CA_DYN_DLY_SEL_RX : constant is 1;
    attribute mti_svvh_generic_type of PCS_CA_RX : constant is 2;
    attribute mti_svvh_generic_type of PCS_CA_RSTN_TX : constant is 1;
    attribute mti_svvh_generic_type of PCS_CA_DYN_DLY_EN_TX : constant is 1;
    attribute mti_svvh_generic_type of PCS_CA_DYN_DLY_SEL_TX : constant is 1;
    attribute mti_svvh_generic_type of PCS_CA_TX : constant is 2;
    attribute mti_svvh_generic_type of PCS_RXPRBS_PWR_REDUCTION : constant is 1;
    attribute mti_svvh_generic_type of PCS_WDALIGN_PWR_REDUCTION : constant is 1;
    attribute mti_svvh_generic_type of PCS_RXDEC_PWR_REDUCTION : constant is 1;
    attribute mti_svvh_generic_type of PCS_RXCB_PWR_REDUCTION : constant is 1;
    attribute mti_svvh_generic_type of PCS_RXCTC_PWR_REDUCTION : constant is 1;
    attribute mti_svvh_generic_type of PCS_RXGEAR_PWR_REDUCTION : constant is 1;
    attribute mti_svvh_generic_type of PCS_RXBRG_PWR_REDUCTION : constant is 1;
    attribute mti_svvh_generic_type of PCS_RXTEST_PWR_REDUCTION : constant is 1;
    attribute mti_svvh_generic_type of PCS_TXBRG_PWR_REDUCTION : constant is 1;
    attribute mti_svvh_generic_type of PCS_TXGEAR_PWR_REDUCTION : constant is 1;
    attribute mti_svvh_generic_type of PCS_TXENC_PWR_REDUCTION : constant is 1;
    attribute mti_svvh_generic_type of PCS_TXBSLP_PWR_REDUCTION : constant is 1;
    attribute mti_svvh_generic_type of PCS_TXPRBS_PWR_REDUCTION : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_PD : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_PD_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_RESERVED_2 : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_RESERVED_3 : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_DATAPATH_PD : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_DATAPATH_PD_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_SIGDET_PD : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_SIGDET_PD_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_DCC_RST_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_DCC_RST_N_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_CDR_RST_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_CDR_RST_N_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_SIGDET_RST_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_SIGDET_RST_N_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RXPCLK_SLIP : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RXPCLK_SLIP_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_PCLKSWITCH_RST_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_PCLKSWITCH_RST_N_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_PCLKSWITCH : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_PCLKSWITCH_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_HIGHZ : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_HIGHZ_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_SIGDET_CLK_WINDOW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_SIGDET_CLK_WINDOW_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_PD_BIAS_RX : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_PD_BIAS_RX_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_RESET_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_RESET_N_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_RESERVED_29_28 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RX_BUSWIDTH : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_BUSWIDTH_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_RATE : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_RESERVED_36 : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_RATE_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_RES_TRIM : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RX_RESERVED_44 : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_RESERVED_45 : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_SIGDET_STATUS_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_RESERVED_48_47 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RX_ICTRL_SIGDET : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_CDR_READY_THD : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RX_RESERVED_65 : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_PCLK_EDGE_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_PIBUF_IC : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RX_RESERVED_69 : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_DCC_IC_RX : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_CDR_READY_CHECK_CTRL : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RX_ICTRL_TRX : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_RESERVED_77_76 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RX_RESERVED_79_78 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RX_RESERVED_81_80 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RX_ICTRL_PIBUF : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_ICTRL_PI : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_ICTRL_DCC : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_RESERVED_89_88 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_RATE : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_RESERVED_92 : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_RATE_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_TX2RX_PLPBK_RST_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_TX2RX_PLPBK_RST_N_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_TX2RX_PLPBK_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TXCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_DATA_POLARITY : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_ERR_INSERT : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_UDP_CHK_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_PRBS_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_PRBS_CHK_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_PRBS_CHK_WIDTH_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_BIST_CHK_PAT_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_LOAD_ERR_CNT : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_CHK_COUNTER_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_CDR_PROP_GAIN : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_CDR_PROP_TURBO_GAIN : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_CDR_INT_GAIN : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_CDR_INT_TURBO_GAIN : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_CDR_INT_SAT_MAX : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_CDR_INT_SAT_MIN : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_CDR_INT_RST : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_CDR_INT_RST_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_CDR_PROP_RST : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_CDR_PROP_RST_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_CDR_LOCK_RST : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_CDR_LOCK_RST_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_CDR_RX_PI_FORCE_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_CDR_RX_PI_FORCE_D : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_CDR_LOCK_TIMER : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_CDR_TURBO_MODE_TIMER : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_CDR_LOCK_VAL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_CDR_LOCK_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_CDR_INT_SAT_DET_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_CDR_SAT_AUTO_DIS : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_CDR_GAIN_AUTO : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_CDR_TURBO_GAIN_AUTO : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_RESERVED_171_167 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RX_RESERVED_175_172 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_CDR_SAT_DET_STATUS_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_CDR_SAT_DET_STATUS_RESET_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_CDR_PI_CTRL_RST : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_CDR_PI_CTRL_RST_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_CDR_SAT_DET_RST : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_CDR_SAT_DET_RST_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_CDR_SAT_DET_STICKY_RST : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_CDR_SAT_DET_STICKY_RST_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_CDR_SIGDET_STATUS_DIS : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_CDR_SAT_DET_TIMER : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_CDR_SAT_DET_STATUS_VAL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_CDR_SAT_DET_STATUS_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_CDR_TURBO_MODE_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_RESERVED_190 : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_RESERVED_193_191 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_CDR_STATUS_FIFO_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_PMA_TEST_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_OOB_COMWAKE_GAP_MIN : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_OOB_COMWAKE_GAP_MAX : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_OOB_COMINIT_GAP_MIN : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_OOB_COMINIT_GAP_MAX : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RX_RESERVED_227_226 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_COMWAKE_STATUS_CLEAR : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_COMINIT_STATUS_CLEAR : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RX_SYNC_RST_N_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_SYNC_RST_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_RESERVED_233_232 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RX_RESERVED_235_234 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RX_SATA_COMINIT_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_SATA_COMINIT : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_SATA_COMWAKE_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_SATA_COMWAKE : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_RESERVED_241_240 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RX_DCC_DISABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_RESERVED_243 : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_SLIP_SEL_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_SLIP_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RX_SLIP_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_SIGDET_STATUS_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RX_SIGDET_FSM_RST_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_RESERVED_254 : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_SIGDET_STATUS : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_SIGDET_VTH : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_SIGDET_GRM : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RX_SIGDET_PULSE_EXT : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_SIGDET_CH2_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RX_SIGDET_CH2_CHK_WINDOW : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RX_SIGDET_CHK_WINDOW_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_SIGDET_NOSIG_COUNT_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_SLIP_FIFO_INV_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_SLIP_FIFO_INV : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_SIGDET_OOB_DET_COUNT_VAL : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RX_SIGDET_4OOB_DET_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RX_RESERVED_285_283 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RX_RESERVED_286 : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_SIGDET_IC_I : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RX_OOB_DETECTOR_RESET_N_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_OOB_DETECTOR_RESET_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_OOB_DETECTOR_PD_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_OOB_DETECTOR_PD : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_LS_MODE_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ANA_RX_EQ1_R_SET_FB_O_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ANA_RX_EQ2_R_SET_FB_O_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_EQ1_R_SET_TOP : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RX_EQ1_R_SET_FB : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RX_EQ1_C_SET_FB : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RX_EQ1_OFF : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_EQ2_R_SET_TOP : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RX_EQ2_R_SET_FB : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RX_EQ2_C_SET_FB : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RX_EQ2_OFF : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_EQ_DAC : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RX_ICTRL_EQ : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_EQ_DC_CALIB_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_EQ_DC_CALIB_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_RESERVED_337_330 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RX_RESERVED_345_338 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RX_RESERVED_353_346 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RX_RESERVED_361_354 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CTLE_CTRL_REG_I : constant is 2;
    attribute mti_svvh_generic_type of PMA_CTLE_REG_FORCE_SEL_I : constant is 1;
    attribute mti_svvh_generic_type of PMA_CTLE_REG_HOLD_I : constant is 1;
    attribute mti_svvh_generic_type of PMA_CTLE_REG_INIT_DAC_I : constant is 2;
    attribute mti_svvh_generic_type of PMA_CTLE_REG_POLARITY_I : constant is 1;
    attribute mti_svvh_generic_type of PMA_CTLE_REG_SHIFTER_GAIN_I : constant is 2;
    attribute mti_svvh_generic_type of PMA_CTLE_REG_THRESHOLD_I : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RX_RES_TRIM_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_RESERVED_393_389 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CFG_RX_LANE_POWERUP : constant is 1;
    attribute mti_svvh_generic_type of PMA_CFG_RX_PMA_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PMA_INT_PMA_RX_MASK_0 : constant is 1;
    attribute mti_svvh_generic_type of PMA_INT_PMA_RX_CLR_0 : constant is 1;
    attribute mti_svvh_generic_type of PMA_CFG_CTLE_ADP_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_PD : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_PD_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_MAIN_PRE_Z : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_MAIN_PRE_Z_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_BEACON_TIMER_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_RXDET_REQ_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_RXDET_REQ : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_BEACON_EN_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_BEACON_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_EI_EN_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_EI_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_BIT_CONV : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_RES_CAL : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_RESERVED_19 : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_RESERVED_25_20 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_RESERVED_33_26 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_RESERVED_41_34 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_RESERVED_49_42 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_RESERVED_57_50 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_SYNC_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_SYNC : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_PD_POST : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_PD_POST_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_RESET_N_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_RESET_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_RESERVED_64 : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_RESERVED_65 : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_BUSWIDTH_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_BUSWIDTH : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_PLL_READY_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_PLL_READY : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_RESERVED_72 : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_RESERVED_73 : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_RESERVED_74 : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_EI_PCLK_DELAY_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_RESERVED_77 : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_RESERVED_83_78 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_RESERVED_89_84 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_RESERVED_95_90 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_RESERVED_101_96 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_RESERVED_107_102 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_RESERVED_113_108 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_AMP_DAC0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_AMP_DAC1 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_AMP_DAC2 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_AMP_DAC3 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_RESERVED_143_138 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_MARGIN : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_MARGIN_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_RESERVED_149_148 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_RESERVED_150 : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_SWING : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_SWING_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_RESERVED_153 : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_RXDET_THRESHOLD : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_RESERVED_157_156 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_BEACON_OSC_CTRL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_RESERVED_160_159 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_RESERVED_162_161 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_TX2RX_SLPBACK_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_PCLK_EDGE_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_RXDET_STATUS_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_RXDET_STATUS : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_PRBS_GEN_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_PRBS_GEN_WIDTH_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_PRBS_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_UDP_DATA_7_TO_0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_UDP_DATA_15_TO_8 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_UDP_DATA_19_TO_16 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_RESERVED_192 : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_FIFO_WP_CTRL : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_FIFO_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_DATA_MUX_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_ERR_INSERT : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_RESERVED_203_200 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_RESERVED_204 : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_SATA_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_RESERVED_207_206 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RATE_CHANGE_TXPCLK_ON_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RATE_CHANGE_TXPCLK_ON : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_CFG_POST1 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_CFG_POST2 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_DEEMP : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_DEEMP_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_RESERVED_224_223 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_RESERVED_225 : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_RESERVED_229_226 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_OOB_DELAY_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_POLARITY : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ANA_TX_JTAG_DATA_O_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_RESERVED_236 : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_LS_MODE_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_JTAG_MODE_EN_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_JTAG_MODE_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_JTAG_MODE_EN_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_JTAG_MODE_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_JTAG_OE : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_ACJTAG_VHYSTSEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_RES_CAL_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_TERM_MODE_CTRL : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_RESERVED_251_250 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_PLPBK_TXPCLK_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_RESERVED_253 : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_RESERVED_254 : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_RESERVED_255 : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_RESERVED_256 : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_RESERVED_257 : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_PH_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_CFG_PRE : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_CFG_MAIN : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_CFG_POST : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_PD_MAIN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_PD_PRE : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_LS_DATA : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_DCC_BUF_SZ_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_DCC_CAL_CUR_TUNE : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_DCC_CAL_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_DCC_CUR_SS : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_DCC_FA_CTRL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_DCC_RI_CTRL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ATB_SEL_2_TO_0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ATB_SEL_9_TO_3 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_CFG_7_TO_0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_CFG_15_TO_8 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_CFG_23_TO_16 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_CFG_31_TO_24 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_OOB_EI_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_OOB_EI_EN_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_BEACON_EN_DELAYED : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_BEACON_EN_DELAYED_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_JTAG_DATA : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_RXDET_TIMER_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_CFG1_7_0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_CFG1_15_8 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_CFG1_23_16 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_CFG1_31_24 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_CFG_LANE_POWERUP : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_CFG_TX_LANE_POWERUP_CLKPATH : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_CFG_TX_LANE_POWERUP_PISO : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_CFG_TX_LANE_POWERUP_DRIVER : constant is 1;
end V_HSSTLP_LANE;
