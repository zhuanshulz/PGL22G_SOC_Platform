`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WIKd07v6PTymAKva8LCV90sv0LWB9mYetDu52euXtZ9cOSu+GVHz4qqbpHwy0CA1
eYfAw83VU0lEq7VoQndTYEDN6RL5St8YrAqf9GATLr4TJB+IoT8WHHBAWCKUmJzA
vQW2wr8383nhuUTbeeOFH8/QVBTqIJefDLHWA78OIy5L+bfy2GiELeVrhiNzPKkz
l9Dvpw4fYVqcrYIUfi23VnywBqJ044hRtPnhogJHrHBPzwFipj1dK1UzCyOXdUOe
qvFfcIBc6V8xL8WOaVjsMr5kEHOc9iRXFu6Cje6gBE6XsZbmufu02C/taFK3Tb+6
twYttXkIoHf9UVn5dmWF4o7B36+vY4h5wHp1JOEpTUD94AEqZJT1IgdbZYubE9D+
yArlqilFxsrsMFCR8ESAsvAsWEyWcAG1ZkW90Rm5hOj1sCBUAPprpPp8tOoLmHHx
pGSp71BnZHA0cj4HNIkpmWDlh7drGT9PWm3Zv1HbR8DLLx0j7jCaVeGtKVLtruOx
38hDi+B/009Z7dqE7FySdwkFSdOO2RMNcyhVoK5UzQqtcospp8GmEmlyICUZa2UM
j7ifREXSjN+7CWMEkssDtKOE0r98IABw+FpTHcb0s3HF+CFoRa3qa9Oxq96+AbTy
IUiSUoWakTTG2d0L973LmVaP+FRRcaBZclIgwgF8n4MOxIhMuF9futOO/3NwIbLj
K9iB7nJG+28nePIbRBi0z6fHjBu7HBtHe1Vh2uOVoezAbLDdaeRtKcbcIwgy01Pj
72lLZ2/DaWO7BKmV7FpkA8Cm9Agd6yy/MQoMLXI5RZOtFgagYXizhFVUlnOlh9Gk
LrSIMsLh2iIw2hWFDyW0wC/bOIuC5TaSoUDA3B1YvIJdDnXsuTPbcT+o584rmRqx
AhOddWtYJUQWz3FVWgrbYQY/Kw5ljrcFAB6828R6IRurMkKlnLhhzlaVmNRyLB1K
SLj1/vbm+NmR4eLoXcc3KxYD74EKJYn52hiBQgPTZVmO2Ol/pemsx6qagQjLr8ik
kV5JpmCLsDqB79yEAPrpr3gvbe3kwwqK7nwJ3t99CnWh/ZEhDD897NtpzRTaYoGw
tsTZMceTwq20WAF3feiszp8SmMHxEyirFRFMi8fJ/Z7KhdMPTaFwfoH6ZHWbzGnw
w6sIYqAf8l3r9b/VqzR7X3HHhxtcF85p56owF+T23DkJs28pnbYQ3QifZC0sPBnS
LbrxteV3YFUTnawXuD3RGvzYbF2x04glEHH/jflo9FoVsmDTHdTnhn9kdujWOMdG
+dvIE31m0rZRg33g2xQs6+4TzTe0OMqEN+70LAej+CTsu0XCzf6h3klyZCAah4Qj
z6Kw9HxQnhtxWw6TFIitFYRN3BhHRwh/KpXfL6/aHwT4VSEqSlQ4Y6UBV7r/nzjl
12+pRwz+u48vqaOJOXVv4vvFU+tc+vyU+o2asp2wQbmF637MeaUwbg4piNlKwpv8
s0XI3crJfWuGOVPw4hoR1MwIq/wU9KLNQBedqDse7wqKCO0c+MlHk+naK9kX3kxX
zfdBodvQhMmmrZqHtZHkCrXIqUr2wzVQCGqJf3cb7vhw/nMjOcCqfAaNPKwX1N4E
zVNn6Kld8OwI59+hQgk2BQRahNVMFIqO4bioViVQu+bvD4mPx9Uttc5kbAUSOTqe
vlex+lail82sOkC0EmTuYHriMQghwpWwaUwQ4/2EbPmmoNuNQ+xanksHp/jKFf/T
wMKUq7Du1ZE53COMdELpmrJR5CNPfaEzU16yv09ruOjRa0Fvlb7R77m9/DCUjvwD
dIH4esAekvkky5C4F0YNPXusrruIYLI6Pqay+wMh0GREv4LmnIRo+KsV39NfwCXO
ZpziGRdcj5tCTb+M+IYYk1gFsFYx6PIymAv/EVVt0CIZ50878fIaeImHTZ7Bdojq
NWU9679TXF6w9AnEbybC92Kkn7TvSiTucXSCTG/n8r0dI/RfFTdusywvU+VB04+v
zeRv4ocL5OUByJ7iP2kzc8HoqyBb7NDlb5SNqQiVNsotKiRrdMXhq1QiGbnJ4bAT
ej8Gjg2A9P1wj3xN+pbxEH513ndex4edkkvP6riFMvFGIY4HCIoHomCsYB/iONkk
tUZlEqwX3gu48z74MCKCA0qZNL2+yZYth4lyRuWGKsDg4ziRuGdhuS1KWB6ZFhjb
t1SwY6kQlmNlPXefX4w1TNIvTRAms66A9FHzG1OEadQH8ceydRDzqBL3W+kvJrfu
Ad6uyrRtx8ixz0RJP12d2ZfBbACAh5weyk83KJN+XzsO3W3NIdhX9RcpwIDlNO9A
wFfhEz23i07cUiqvMzA6Zkbpmv2BK5+mz5vxf8dnog4QAwRWv5xZU69V6+kO2SF7
Ma7pxroNwwYEH7ulx9kqaZm6A82b/ObXcqjXMFCV6TaMNwOiYu6xcSrPNvNabX/k
CaTIffHCh/Q8bhSLu7GnDAHde2Lgyz7y3u3Awjv24W/YxDmleXiGrefXq66oyomV
zXYAyqrw7hTr8doSRelpNQ==
`protect END_PROTECTED
