`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5fKyRkXbIpit0LaZvMoPBYuq7PMxdKCIhyGYpE8rckZwVsklYqMuoJqE2SFxq0Lm
r51iAc6OjwpjaZI1lLfvK+W7Ot5H3GpT9K6eMN5sKmlSrgkpLmW7ZgEARYrPQJ6L
WUxiFNCkJGPt0SV7BbNGT+3WiOpjfcAbXsnlHubMvFrlbKn8YidD2ITRydUaIZWF
t5GzK9jKjWhoZ0l3eWvulwfeeRtywfuhknD29NyVSbMmBBELtFyFfh423qtaPqhL
Di6uF424kSfdb0AaAsgf/kSOAEjA+5SwEyQboKd2UAgVUwnaVq6E+SHHoKecsyur
b75v2mPWbLc/aWEXqQ4yzzMOWxle3KC4o4y8Pns9JFz4H8342N7vjJj58jHWYJtr
sIJ3G9jauwOfXYFyES0273dXw4KCR7onpL8UWz/+1FrGWRlswJnjg0eNvfxumK3L
HO7nmgqxHgBgxJ7o9GWCJbE0QC2+U0ou5wQ8s5nD0alURkpOtgaJ4BxqALn2XJBu
Y3ClAzNXFU0H99d3aN7boCpiZOeJq76i1/DO+EtgP0b78dHL6+ff2PQj3p1VNAYP
/fIW1g8x8thRNZ0OG+RiK3kvGL7XfoYD3YWAwyTC+tX+8jIm8ij5MKT0R6hJ9Jf/
jiOzvXDFuVm5fkXEN17lr7nrjzXJ3Q/3ARxFG+V3f2EVaeluwm/M5RCyKJFKU+9g
8ifSO293axuI+8WuzL8fYVxVkCWd9VQ9KHi7Xyg36VnR8MI+lwuNOv/oTE2z9tcv
Not0L+xi3N31cMMc3VNAUX9qznhJz1fiIvpcfAoqAg3gCaUiEgB9u2+VuxMeMEwJ
Q3Y3g9uWIs8Sq1qCGKYX/in5pcrE+xdyvTFiKpIVKynPOicyXyK1l3yh9/5zPxf7
Zmkby5sVc83LVAZYfCMS4Mp/qXSrSp7HxzCjJuKNBnIakz7dLcZnQnIuGR1ut8HX
vpPGtAUK0gx53Bve1mvbJH4vJDdkxabkRQ+AJ2erNmk2ePNiLKlSr71dN8Y1NsCj
qL1xlvAWnsSP1ktbEFiY6mYJ3IVH3B3xpHKfYZCHauzcGlvvZv7/7ZgVrh4VJWUL
8bpKcbJobEApWOkY+FVCuf71ivVCKsbOJeJ3R3P/FMhl3RSDW7dUbuoW0B7Rl91a
xTQuOEAGpt1NjBd4Dx/mUizzXRWPQwEdbmEpmwyqOYJe56Xe0yD+D72tZsqd38WO
WWib2V8699WaHRHbCCEcVZ0yNyLD1/99GdFQpoIj5kVPlOmcsyxamy5Kb9jPBvl0
Bvg/ZCxzVUsD8yaibQxXLXfX830n6Td4K05eiitaTFoJ6ApyLRQIgmtlXgOJZ18i
LYWDlU/IF2L7E8Vd/qsEEeXMhSd2xIlWBeKug7m3feOMy5eBEboXnvl2DgvjCd4r
8uAUoLRZAH16NRa7EW9EVg==
`protect END_PROTECTED
