`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uMGtOmbIsi34CdTbOHKm0XHZMC5LBC4COyKXYhpGzB3VByR/SpPNkglyQ9hLmY3i
wzPxADXwUV/yIDkSNcw2acD3RnNJnGSCOoVqVaRsyDMmQegIjogrFTUjd9TDboM7
HDw0FTlOnOX1S2dMm7Gyf5rKcDMIiRHCw0OQ9itIovOGkFdRrwPRXUCY5BNNyVmb
uNNNiWPdb4BNnWOYa6SpxiA+QRoyo4t/ApI71FTUFnSQUy9ILw0yNiLCzKral9Xe
8B5BrE/uT1DmHokR3BgBSubhliM6ilYw7/J3ApVvOpJJVbG/GZTyUrZQnG4ui6R0
xngREJhz3F3UHhHEVxYlw7SyxdWqNXC3Q2gijjZB3csY20q6PYRRzh3rYwb01a2s
zon+S27r8upguI9Gdm1/EbgBAow8jaan0pUfUTfDsiOXcfuGaR2Ipj7GN31jvCI0
VcIDqBeMUKjAXTabYIB+d6ZhEJRyiF3gcXMF9SdBylZNxadO34WebJK2/gW7UhDD
t1VrxalhckeHYrEC6fJXn23gVxa30kGQakVegma8f+tgYpOveQaweRZxhX1/dMCV
cyKDGJPC7bNS5fF7fqWIELZb3K6RH2qMh55syMYR4gE=
`protect END_PROTECTED
