`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+eNoKdDpwEHBO5r73obdcYEQW15VKIfFNTErOB8Gg5apFj/Q7ThL7e6gH65eOXby
uYtmoIbzDaA0DW5wPuzPfcjOvJIHPF6PMxuND6JvViJBzgY28ob+eqYnBrBNLX7B
TqxkR+YsHd2zKssWVWAVYc69700WsRjWgAXYMhqF35lXdjjEiscW9M2qxy16r2ja
PcBxKVucCwUWT306qa+Rn5Vjw+6kuuQ1keYG1G+hAkPT9f5dbqdJ0JrKJ6kqmJ+B
pjwUdqE5n7wO/1599XsSa7a5LJQojYDoL26MEhBDvY6lzqojS226wl8WTJkQuZkl
QHtB6BYjSYkj6z99YrqRkpKuAlUORPC82Roy/q8HtxiRLsY+RDis8hm7HHXpUBcu
k+h722GybALJknqndv0xVrSYaFV5uRvf8SFozEcyHbJ8uNfS/DxeygHDeFxl0hPb
nNjSwtbNW+mOgGY2BENLcvEBKyfUYLKNLhpJHMvH1KefkadYhjRelQkBxXlGB433
H/PUThoSsNlimNId16aoWSNhmsWo1UmSCOuJZfvjPGANc3jdDUf7FqZIoD+6U59S
IJeeFeCEhpR+iCvpuN5JDld/WRCkQMhVYwaozi6EcaY=
`protect END_PROTECTED
