`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OPifvf2E46cPp+9NOFHx0lwFc1kGWhERQEICYxcN+m3itjRpUV+yp/REDwiryD6B
m8Tbirgb6FTGlN0UZ1XicJC8ETwAC02K1Vf3zerSRBt6fUct1g/XoMVGlS9fKMzE
n4+PsSF5Rvg7iNh5iwbcNLyWrnw6GqwjvTuzM0kBA2evX5t0YTp0fb+LTKszH0gG
KK+ogfTo3yRr6BdFR9RZ3rCs2DxwKytW74v6XetlH5dKW1qqvXHQKT1OJ9+yTN0+
nAYoAwZ2jo9fOx+5OLmS+AOMOwHMWOxxtLXKJpPomoF4S2TNw11YAQEpUh5ZKpup
kMOwVzoveOtqDeM4+4A5hWxMVvsrZvizlAp82z8FjH6bNLVNUFtFPm7XPcw5MvVY
N+AOmOURDzmQwyfhp6w9mR1GORyTUdveTvYBCuO3b3kQlOmbosGQOc6DFukqKnJe
s6YjdES1ZozNr2BkhOsVTpux9Mpxa5A7apihmdfZgLVyI1vI5aT57OB7H/gWhomj
pvfGhjhLSefESIRhYr6lqc+33Vlvj9drwlSA/Rno0qDrjr5RXBbq+9voQBC/CLJt
rvpftYOgi/ANoJmH91At6TjdZrhyX+mDXn5aQH24GNu3BzshjryQvwxplB6U4DwR
ye4Y9IIpdVcFPDLDeH1Xa0byeH4UAnTwQqfSUzisgSABG14Pgj35jaKkq3AlU68C
58k5DMefqjZJ0EGzGipdwGOJsoMnZkwO/CRxSTl9k/EqaYMVq0vMAV85vQOsFZFS
CmEeU1BtGxWPeb8k24JVOqKh00Ic2tbN/+A6aleYOFxCcx6O30uDj2neZT6QsjKu
OPelx9LJUGme1AB4mwkVX53SqomWS72L5z9nHR8jbOq1111oe9c02lrCCmibZrHy
v4EtPT27DnXjOYzyRHAWOaAPIEgKH5G8GT693g8Mc6zZT4dRKBwmsRwZ8CraJB6L
hQvzrccCvb+L4n1ba7UbVRMnprkSnTDu/G9jaF1kymozHySVEzLzknDVjkxQ7wYa
2Tg9jwwP0O0whZcXru2WEopXn3D3azYJUsmJKMyIJ2MKQgKzDnrqNazFrWlsC01O
AoMiMQhdH5304ZWer5GjhCM9Uq84lHgKIiZbsaBJFKxVRHWo4jTIlOrzG59oGMwU
8nJeFVrpvNkc0+wLNUeEVgmm4+f6KfdGYovloUebQXd0+qrt1XwJunfq8FD6KlCF
aaqXRwepB1hEy+6h94KEOWQRoQ34pEN3h14FHO47Wptb/4IK89d9aljQW7mhcnVP
LgvoIuqCRJykd+ix5WsR7Wrk3XfkCs70iKHW1ZdQTEuC1wygYW0xJkUqR799PB7i
crAYbKJsC7ZVGy+m+kYAugdnQgxp74c40iAaWjVx4oA0Ug3bjJMRY0unbmqv3ibT
x5jK+PrCqV3oEpllmU99H8mat/1T+hUs7bbP+Nd0vApB6BlFJeOClRlk0nvPkFXR
EqeAwDroTdq5yt19jyN4m5ZDbz7k74BU5wZiPi1cQKjnipEfkjKok7g4pqHQpp93
eJxi5Q44N/EB/eImZLzqOyY3Lcm2T3Z3Lt5QIerlOrc949cGcGa6v6pjc9KHOzLH
U37fwHwSaZnfE2SqZqrnulrUrw0kmvUnEFW8BAA6msXRtoRNKw26+KCcuwmjysX7
DPIofQCy8I5hyB2pgDjAJZNfIlpEg3EgnvvK6qhIxUp8hrx85jui3zWdV+q9t/e6
TPukcOYBt1yb4Q3Y09BHTKsXl+dg/3hh943TxX1ipBqkwAmk/uzkpgy8S2FVpyZ0
6ERroKniqxL378MvxGgdlu5oxQlyub4jDTi6TiGCqPuKASuHtra/D9Soa6JlBsOX
zc8lWBiCXoOhkJSmkWzESYUp14y/f4hBj72js70hO0gDOAqsjtCmv/Q5SOS/CIE2
Z7IhszWhmPIH5DcGf9bu1T2jLxHPP6wjZxQVyuMvfFgG8CfLG7fA4mNK0EMomwag
2jE/7hcGWTvb/ZcOLwA1uMKt3U/hWYxsojTX3p/q1Dw+BFcKLIwAgmWUkKimpDwR
ss35AFVlUNQm6YBGAczj2TJvS8vZ8tkzf8F30wdXb4vOADbL0qh1/NDD0LF99RcY
TAJ9fEhdfhpRoET8cM0DaULkK+Wf0b3wEmVBYwrT9sk=
`protect END_PROTECTED
