`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D/x5HJs5bkKsLd164Ryskk8lCy1zSjx+yC3uhznrxGE9H61jJD/47ngNDOg9S8xY
T3Dqw3vMBrM/TJqnI7l+aYOERt0IFAULDlyQb2ESoKvb/0S0ZLF+vPIYm/Ljg7zR
2nB+wq91Tcm6mWSNNpfeARqoSukExdioKI/9nPdDXug5hhizFFXmJNpT5cMW5gLy
pF+Sj9QCOinzOc7+w9OpSmDM8ehaApUL6lGv/GvtKD02xnsknRENqabgM6SQAH2o
XIPc+Il5AxxWE6vH9bu/Lh3oYAzEnjCog8x3n1ogmhFHOxaTS/0G4lu5Do3hh7oR
uP2czjEn6Ck5bt5fA/Ixh1EIEDIRQ2L2vt8kDm1r+qLU2oRcu9YFOGQKi81JZeKl
cob2Rh1oe/cMbrtliZNJxP6C6U2RVJfy1kc1dlMWCmZ1sbp8YDcpb++66+hlaAjV
nQmmYiY67lTaqCZOXqdyZnBPwnJhSgTAcz3D1DrGWVnW/ulo0LF4AH4blfwjtZOY
z4l8gymSL9bf9H6gQ1OTcYapzS2/85laVy27mr3fwh81zXJEqZNBx62PRGjcsLKm
KrCnMMSHyUJ0B77jNi2M+yezlEzSfS5mpvGL7QOgc5w=
`protect END_PROTECTED
