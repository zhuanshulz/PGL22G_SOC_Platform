`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IORQ7KfNzB54rhNu1tXnVhkFrW4K+emahrWmGduZ8HbCm6vh3l9PpHnRlv7IG7jV
GpGG95iB3/qY5NOiRwo3aDKTJGkFIgjZwue+pT42Eqp5vfAl7P867tZKtcLVbP3V
ipPPYAPEILn2x2M4FG8mIcmOb5LyDh/mVx1PqQspScWBlmgfFI+G/xGCi//sTOiX
FPjZvLWDZzMhAOzMx+AvkE84uTudgigfsuAKs5FsDUkSEW/1jhURSh2gbVlrkI09
fzI4uWmCEeSZB3cBQFmGO59aVGXpkrmIk1KsAHAoqT786zb4Q308uGh/U442NxPi
Ubz135RnHJEKegTCOdRPwHP90g1XYTNueu67DxTHgZbV0/r2N3UvREt4zSrVcJlC
35f0r/lCQRfS2aNjomHGqRRqs27Fpia0+eRYaILIhWWnkaiUzENgH488IE7e1izF
Jh/bZUz6MN0ZBBkbevA7byOsqFfl/dBYHDI8xDuOnaTW7+xHQKXk+sll/24v6Jzv
RN6gzHMlCQZAWn+GUb3tgnL8NbfZ6gHSmUE+tjDqPyNULl15crhyYDMcHBedyjAw
At9+cr2xrCYJkJ+6C5mJV5LQ0DlFM3q1xq5RbwGsdIsn3cd3qd1D4R+tDFnFJYPb
SPw8BCuy2Kcb5+rQ2chVATvurSv320K1MILa3D5Xajfe2yLlPhxo5tKcf1HVooFi
7wlFC7P959JkXRlDMhmBFEWLsnF0Ip1MfjObIDXFdk2GvA6xxjP24+1zPz4lzPXC
8gOC7Fi1SPPhN09bwgFCJCuIOuhBzy3sxNZPCXZQKv5PFZ0iVcxAwjn5WRi9xSOo
y2SWtZakpBFM4+QDTUe2GMJshcIlD7XbGxClUgj6j6DkHmgq/bBwYJS4Mhj8aevs
pl/5LrzIrO+eBLoiILO1s755CRrMqLolVwy0s7AwcVGgo/oylGNEADaaRwUPd5Ge
ZCL5Dnyw2iSMPD/EgzBd3vfo70s266fvv8dWhVJ8dqrnJSqsN9+L0v3QD9xZPaE9
7Xmv+qMegpJO3r0e81uzvUWra3AbtkLjagWRLSDae9jfyxbOgI7+yu0OCC7grnm0
AX0+fHun79MuJaTbrqgBBm6ZUunKNElDSnQvc5YwYbWggBAUEbC5pBVXEWyNtDn6
55ev+CoT3bgDzgkcrgrwTKWiWydLToFwds+pT/tAmp1tE/CGTyqFxWF18jM3J1EZ
im4vmfJnu8/G4kHfbHnO93ownA1u8uNuJFtF06/uKNCJJVsP2VFbaPb4U5ICrWGy
/j420LRV6KBbuRP5eC1fSyWqoMCDvKkvqD5wCvFIL8fMZh1V2570L7Hm4o6M9ZsE
lNDt0U9jFm2mEb47U6tYGLcKX55avWFVqto6fBAPY6LnCdssTrj0O/ragRvCePvR
Ndf51YqsdPlVMIbIjPZxpFKCuolwfg/x21tG+DhEzJa96BjJ+MXsN6St+ui4SFMj
coUcypQac2EBskUGVjiu9eTlXQ5Yg7hoUg9xqhis11j9jWhcZmAYhZEqfX9rBi6w
K9ARY6Aa+XkVsQjABWFJVYKK0zYTlZPMTkr6qGPeAEcg9O87lfSOZNFqOHu+Hs+v
i1TlztxzDor1D7FmSr0HmrO9hvs+sTbgCLmu+mlTBhd61xK8qYPSeek3dd+CGAP4
dfdMCjNxp6p/e33soxUJm4uzf2/7xN/VwiGHNxwv21xXyXRE1CcCHbtso4gHkC9L
ziZ82KTgFBFwc2jm8yk1uJWEPScEuN9VyS0/axmSLITIEFRupM30/MhGoBri8y09
bR6dvRFwn4u6QlaNEOt+Js9scl8UsSgOHYTACWhFjFpSBFHRMn7cV4qO9l3Dc2Pb
8c7xkXQ2dVBqTxOTPSOi/uhgKRdcRc79r0THOZYGfLBQgKRMEKY3XUqkf9/qkEB5
/qhY6HPOMDA6i5IqD5rWB9cawEgqOpmhYlBqbhDy4Znk77UCLwg7aASz78moG3VI
O+SpBuLgiaoXm1DtKf407Zw5UnAcze6D0hAcdiIjqbY6VLtRpBkx/E1Ji5FHG8/e
0VS0p2WNuBMix3jftlcT0tFOzYE6d7Fp/f2ZzmJbIi+/XEyCwlqFQoy0rjwCLoQe
xiuQawgj3BM/8g+gmVLU5iC1LmjDDVnOaPFGmhiDMrga8RQbasupt6Vmh0cB9Yx3
ezY5VIAIwmhyOVuDwkwM+q4EcAJlru30M1jVvSEYMuNnEENXmbWz6bNaXaBdhq2X
5xN3T8OKOSLIpAJzO/+Ac8IqymI7Fl4yPog5PQ4jXvHnH520k0oKad/7AjXvjMgP
fu+CJjXT3aoE2LrdIErEtBuXkMf4mqFf9PQHhvHqMu9+kVRx1EPBiO4wYv2JU5iA
xz1egxeclGm363OlCYI2PNXumLiKufkJiQN4rs/icZ+/7Gmj+cNhIgrju7KVCN7D
3EQ4AZAQSL6NcYelUWY5tyXrDM+cbZPTmpPPsQnWT0mPvpB6Cd0gsN4ZWZUA3xu/
+5DGrfU8JbFskWqMIx6rmZnvLk+4xUK+tx5j61rtPkDYMRJte2OZCEp1w2o9cbCE
2Pb0g70ZxnaY9mqJgGLWSv3VVMj6APHkoVFV1hcNfzVZgtQF6cM3+89u9nv2ni9H
VF8hqcflCkKlGyUZKHdHCtwt40C0w+UtV7gHONBnnc6ZYtmQDv6X4hub03RglUiV
uySbwKTP3RBv/nzX3d5N6ctnWkvix2rgDIqemvg/7qEsN5mb3pZYhF1qM3iqgQFv
0VNPxecz+DjjbEWEWBBiuacO0I9oreOuPqnTSws/8RflqXcSTNBJTL/r0hGyYDUO
uO1XZDWk+vC++zLTNJ89TAR91umdo2KJEK7twPdAMXB0Kmlvo59GKTuKw6PDYNlU
GnB3qSJScz7jUhRVK7MezubQU5eeqs6xUQAzl5fAJJVHyREVyj0Ig1g1jv6tZygH
XyvuugriQDusBl0ARvK+cpol5CGMchx6SD1tkJ3zB0RZVlNTlPUvNiCwBZeFXs9u
297GQh4jv/Z3aedPEg5gkfgMlF23M1JFb/5XWjaYfZaUP/j31WbWLnypEvvYmlz1
yUA4fYpuQfHsVub4yRVucxE8MFsoRIj43e5LH9h+OkRfzXmbJvwVnsTqtZjq9OLE
NXbTvgBGKVVViNqqiFbgckZDXTenPz/UhGDHjoBgRdBnVbt2/71uOkKIYFenY704
rER/qk3ergIu9bqvcdU4/E9E+Jq+74ufn0zr17MmtD0TpAOGrPyzjpTRYPpAIZNe
uuS+Zn8ckgZYtPgwwvwj4zIMoF6dxSImX5s5wP/p37zWDgB7k+GEzzEmU5qizI7w
sDes/a9vWobi87vQwMFe0HTZIUtCU2ZCXkYsGE67aPMkx3ZaQUpLZLjHWsBum0QB
9fBMeonnXJo0lBYuVS2rCAtT/ZukZ6rObsXZrXhBzOOcicjHF/gWdTU8rluPssL3
9adSgAdwgQfDpWX8Pi7V+ZhDaEQjPBiohqjooTGB0wZK5S4ENsrzxpHhRjlHvVo8
kN+C6APjZnb84eFILuKlki2FBJXje/SV1JPlGtu4+IysEuWR4SeP44TBmrcDDe4W
29gIQyUzYaN0OEEUG0ceuo3Y+tT//V70q5Wf1uMmW9/fn7hIGM2gnXDtiT5q3lfC
Fc4JHz2SNm9TLUJkJxFd7eLv1UK6hY07Pb2aimuBnOAIV8e3i2Y+yFUgzWMQ3l9w
ngToIqh5V2OqjWxlIkwIsBbg81QxDNumFu9+gfL2Tblt5cFB9EBCoPWkEewoSwi5
Ji5IfUEHgeKDJzKJqPT6QKf8QxhrIuQ6ElfGAo7yI+56vhEBAhMxjwBYYniaySp7
WZ3EKVF3dActLtDYmzuWHZePWUvqnzuWzzcE/tn3NWc5FzcK1rHVygGIDK641C4F
XE80Sg4kOSRrXC4GUPBWuDDrIM8FiRjydfDtxN3WNK6u95FrN9x4yHIFgdMElnei
hJZtNJhmG8ObORvJQbnA6dYAGqlEJ9PipWc6LKUpUGOhjb18DHTkB72buanhTU38
0E4gmUJgsqq+xzbdy/UuozqoSYgG2baFncs3YF0PuaT3wiy+FCp0D3GvQ/Pzbla9
vVrhmXC+ojm7cJS+7Jb3hjdTGCrGiv+n3w6fIIbNG69AA3wJxYufzJJ04MYRvNMH
k+E2IsSfbCVf2ZuZOLY6s3s6FNqaBLcCZpCCGuUDomo1G/tpZiJTrqpT/OTQicid
+qKT5ALSwsFkN/AqP0Wiae721jvIP0Fv3LxbvmGTDtz4GoTwAnVkZlTcE0mVAgpP
jk3Gbn8mA6gDlLtIDfoQRDR+cVifuJ0wkvTP1aigFmGGCEgqDGw86e+oxod5EiQ2
XklY4MbQAUgljCPGpATrwO7XSfZxwQSwHwORfL3PTfZNWbOg1diGLBsVRLsygLPu
BOYwRUxXVZpKeF/zQBKT6Y9iRxrTr6vgkKtEBaZsyVEbCUODGHYOa6x+5NqrQaFb
kJBen/yylYMkifJ4YrRnlmxIdr7YhjncRItryhapJjRALTmHqPsfy2UAQjufkF5G
jeNISjfpkEOGuWAmDWZ6M6+Tct+ydNmnLMrAA9aLLvvimALtgMAn2dbgH7Y0oCxZ
e1d+4Bzwz161pZLJ4qho7S3SsdXG6dg4MxG4qsJdNQA4Q84+r4qUAEJ3NHVTHEeE
JXhMwZ8AwJVfvT8hpYtRLYKhIapscqtXaUa923mv0Nf+aNGFK5GbAsS8xSb0i1ui
BN3h5N4u7bW7Io1zQ+E1IUIg/X66xnVXp6TUTVYIuywOP8V9a3xAxcNu/SnuVwP7
atQDm+3++kBsJ6su+QYgmXJ7SaAUkdOfs8nwNMrAbl0do/kRykidR8p2a7b/uaHq
rzqSihvCOe+fowX2RJMg6NBWQ6sMEqMrJ0H7eNRCp4bRJJcba4U7stIWyVe7Uo8T
9vUskXJFoU8lxLQ4wUzDiYbrAW3ikhjoGngI7t9Wus+XRi7+LLgS8FEDdSkyQNFs
l2KLIOUKjtOChwovUTxAaYzOEwvPANI49TW0X2Ut+MEUMYsaElFv8URUnRee0LUI
AfzcZYKKRHcWCmm1NkkRoF4vIgmQ+iYvwmuMM2rrkSxpHxI/Htjj6IF6cDGlyGOA
sKYHJV568gyTTQ65TxXzpr9wL2PxCrZk0JW6kWgOhpasPCL2cTo/J4TtPDWr96dS
1KSqvm3DbsPu0bktC3ag6RBTNRbVMeQYrBLhmaI+Qakv+nwngMx3gX6LZ4DgW8EK
dtxN+7Zy6OBy6k5vAAqlffYEVH8fmNib/OPm70Jw/qBnsp+k7/ci7hPkV8nr/QrR
WcEVrE5cYTANaSpchYlqXZcIFodKDz4TgUadI+uxBC8ZYXUKwkrwtWeszWGj//yH
7SGCqPpwfy2V9gSZmYxmC029JBJfLyRPfpEcPc94VLNKAjAZ47XWtqfg2a91cl8I
E1gILOLDE5xUCBIe9jPL8kOohWllgMRvxi25muQ4odUvn/LK94q2Sn+OiUA/vdt3
LJigfeip13sfjEv+D1ziG4SlWz8IUtYAvl/RVwIJS5MEqG1I67vvDnK+mWnGmO3Z
wP9UoaWmQCGSnYYPDDova0gK8apcR+QviSeE1/cloDKgy1HOOmLg+fDYpP96rQ20
i/AEqM9vzXQIhs4XYGt0w/IzyGHDZmk3Ed5xZsxID3EInIml9MmJ3nOT2wjkdnav
6cTNrwfAVd3pJleGddq2XsN4Ce/cEZ69Nwru448HtAcjVa/3eqPuTo5gJo7zK+MO
wEQaR11KUstcz+kJHRP5ppY4MZv9uvQ8trB2sQx1Seh8rGk0b9qG4n5ueLnkuMnD
snA1OK1rYMYW4jRd26ipwhjT+scicBUu/dGa1en4nv1SLmCVIzPNHosiOOmiYEuY
OzmEdlDsRi5ZBatIfcFVR3ozyEE/9AXpzsOscmhKeS/UrKFUscMq93l2otRoZfHC
rBicHnaRtdNTVIh1alCqBhEj3lTK478laYQLLxXxr1qNKgmcMrU4RPQfc4xqpI0w
8nDTw6/PYTKXJSI5QacwKTgvtXRf7YUadiphcf8JpDcuOJB/sMeXTA3Ol5jqpgnS
m7EPR0X2a/gaFLbDPNlh3C8p6DGMkhYf2Pbrn55paHEzX89SKS2+F/r0uBGCNC6i
nM5/UPtXyNQTuyyf1QEB03Tsy3H9CrgYmBFKJtpt6wPmuiXIvOj+GF5rIhAS9FQC
w+Jp487Zj6hX7uOk403vdZvfwOj7W6dtmR320V9aOcW6yVJQ23ko9r3Fd2w1zi3l
1Lv9KzNPw/v3AKB7sfkxNV3IlNhzFnyj74KKIDQG/50/NHQ/mBuHdBnyBWPfRDsw
IRYK10hfG6iIF9w3MmfDCzAkTICCwpzoqrYpvdrkkA1Z1IxjnHBUyScghPeF/98y
5qSA0vm5Lse9XLTUYimE+6ITrkFkqxwXt73ilnhPsyD293HcuecmPTSPvT8M8N9l
vh2R8VADFRzLpdOzljSkUobfqfqSWl8HhqFUbT4GpkwM5wSePS56fPZUZQV9K70r
Wc0h9eqgdJ5gpnh9/326F3qtw3WvjvfJNQNISdfw/Zutlp3FG2Cw+jyRqLbgbhHj
Th+L4+rGZd3S2EBm91qCi4bKLs75+pcI6OCGgKknV3KTfjO9M0KRNe4JOSprCvci
57fx6UkYF/CLfIbHFuLx3UL6d939O68EzKpCWDndkOWs5XtLYadK7kMTt10GJQ8B
M3jAIPF+iyk1TDG69zDDqM7VvjCf7dgFaeLSOkBscbsaXN5gsNd95j8WEUgSYgmK
0y5tcMoTdvRhi6DCRTUTLHfGN2Q64rIrCva3I4zNdxphlwHIWqk6dw7AaTxh/qM9
cTpYL0qP2YV8Wbhq9DhD/nEpXv80ec1JjxD6TyBf8NyjGeE/KuL5CSe6AzlZhPx8
W/M/4Q/5tXfth1rKYbJkwmLChaXW1soQSUMXZOnqL+KuIvsidSIGoK5yMENFHwYm
azW97C/MZoQf2Isv3rQRRNJCB9Xun1joS2rPxuZzT67oB+pWg9HD6+kzdajdoYH0
ycr0b3jTN1gB52VmnLsaIWzXlkcbKYJlMxZUcrZoBYu9+k8ISWS9gmWOFHBwTm8B
KSrdwTwgCwMXbrIgzrNVhO+Ol9euoc7BmvNKRnj3Ue13oaa+1iFDSgBETrgHBzKp
hOfqgSmJiLmSfWL0XmuUPhcNGnkJWGuPvc/Y4jNtgdiaCAJqXdzt3AbBxP3eDLlj
QXKqpNe9Txn/oBT+n0cxMLH0jee4sbqfiMLFjWNaOvzvBHP/mjnptGZ+EJQIiS+D
k1SRXLWQhJX1ueE2WLHRn4EZTeMLYaD65/36Ble+LsmP/Y2pKAortSmXirkuarMg
LtEippTKl6xqZSLrIipvoA7uE7sX4Pcf2NGtyR2eoUqRIPgyL8HvlEVHlwtTm0j8
bCcWUqvI22YffNSheXRSKr96takFiGLEiOW/Xgb82S6lfalnElX/BJNId7NfzSeN
SWXoJI6w3KW13R99cOF6ZYHHR7aaVjVW2AWa2glzmFQGASO0m0PWcjoTKVeZ73aC
anbtxvZT4d4uoVUXLwmljnsHNtqjjRCO/L0DxbRH8Xq+YzugzTARsF9AYJB3e/oq
6ysXQpznEWJh1ENiuK/oheC3rNAUBKtwMGr3hdtofjlxDDcqELjyrcJ6iVqoJYqy
ECwPz/7woEdxJoc6UBTr6iRXiCgu0+nzVR5pwqyCO8xhp/XEkeANz6iE2TLjLU72
YW8HMNkZurwvw0YTWlNuwGAfRADbDA65Ctk2rOyUM1F6RPlyBQMoywh29bqS1yzT
iRo8/blOhjwFkS5OunV+9An8NSHMwMibqjbe1s69g2u3idzXs6GLrXrG9Wg9QGaP
96+yRa3fq3nt1U9IXF463TfEUI13DVz6N3BAWp2CWOLQ6kZCeVcaqxOsY+Z7hU2E
Jqc5jeEoKtF2WB2wXRgfsZqx9NTA4Z4dzNP3unT8fWPpYoSe2ot58twO3dTEJK73
iTmsoFaLWcBwwF15mdQCsjpV+Ah1Fp7MpmW4a56GFcyMalx+kPkXzf5eBbth/RWg
/dxskxpYysoqxWKYyn1MgSprDESNRIA4D9rDOMhvtXPe+3RljaA/rRDxKphblIxM
/P6eaqZCU13yHqdVNz8j7JT0e7hFKA7lkSl9EOfy7cgwL1W00CdF6teozIQAboZK
HZL8ih/et/CQMYQ7XuF88dQut3YPQdYsxmjQEE+zHGrwbiU3H9lSwv9wMyVHJGUw
4OON1AmRQpsGwfyNOYj0kdbUkYM1ms50YbKHU9OZvbxWGA2c5SXfAqvpmf9i4QjS
80pZZln1FcCeoNvUhL4a6XDCJriHf4pMcrPRHIAHx6ijx6xR3VIjFE9cAChVhs5+
hxpEKbafzjL36F+uMEtOtrnPlKqcdPQcQKqTChRkaStFvrn214C32g0BV8gFe6mz
j0LeoW3upq5RidPtM9K18k/UNB5zdc+2+5RKU2Vm5jdLaUMQ85GaBtbV9aqkoMrU
u/elsE+mx0U9rlh3Qdc8dbXifqYxalGiVN8okm9xn3j+7vlm/boGHtBA3KkWbTIo
usoqp0pOMSNapB1Ygb+2vFoqxRn9dzHvWXfNLsZ5VpbAADUn5klPFyBcUkS3glUB
uJUth/RtNtMOlYZjp8QuqJ7zQI748D1HttkAFE/l426evwfRp0GrPnZMzUO3IDyh
uMPbN41sxCeUYmsFLXraZbbVvBTxLsEjmYReF235MyfOdyVgRewS+8nyoIJPWi6r
DXF7HvaQZ2mBlprSWaMshfx455HLUqypEg4doCCYRrGRxUReaDVIWAwqEOfs8IZ9
WtM5TMuCAN9xKbQTS5Gp56GOCaHcCsavhJ/Xsf0v7rJ6zEBGnnSDJ6riyyuNU3py
baifUKC0+rIq9TIpgWKNfHK3yVa3gfmYOjs236PO67IdEtG0xLguAoI/u5rMdzGQ
18YX3JDqzRVkZ7VP7S7c3yiRIxLGVP/dQV0UkPUd5F82O8Mn/e4krFmoauACoqAx
7azZbeV8t4vteR5n7TRqIXn2il9FRkCKm5ghXtymhCwb3ag/wJWl4XIwg3JMjzms
VTBKJR0RY1HyBIf0Xh+e4boPycQXUzFEkRLbV1hzGqNpwWeltjsZ4v+UJKOVXiFn
+Q87ULeKV+KIjmph2PjoYojzLhyJrjZIkMR+Awd44NR7RIhaKpbksWjJTIiZtnGU
zdU+wr2mzySfv6e25mrmWE/b2POYObloGzrNdPKVIDmpeBwXxWCUvf+0bJTQjxKS
QpkD4ClGZEvClvmGasDCM5iMLTJMX/D0ljc8wny0XphOVEqALwHJIgef6VCaD5jM
K62EKzsenhNj8lIUA2nfbQhA39PNY5lxcxoxttow478Nmy8nCegqXWf1f7fvQCs3
tI76DxtS9ZVYb1X0HoXrApA4mABNoOXwDxq5s/V1n/uwYTWDCrxVuETcKx85tZ73
mxZQTy/LEbT/fsC/d/sJugB3B4NT974I0GJdVcJuA4MGp9tXsEc6IDXhyRYD8WGI
1s4Fau+qqAMeKFvuhSUvGXbCIdvo6BkP8fGrgoNZ5GlUNBNtfy8cG0/r6WgpIDia
OyphL7j4Ep0Npmw1WqESPc+OMzTE5VNHlrUX+hqxHS1SbS5EfH/gm0H+W8AeHMk4
QmfF1rjLMTmsIIz+CxhTLL/4ds19Y1WTWb5KcAaDapXaDxYrZQCJEG06H7TdS7aH
V8AJpXdC/KOLHycwVQ1IGd9o6teqWhk2D+u/dAyMHSidRmgx5Vx+T4o3YIIb+Nrq
jcaAg8htutWAnDQpy6sBYJq5LVvgE6Wr6Rh+DDXM8yqUtz/6qJ0gICYE6sS7cs7o
LOvjwY9L+eRVCUQBWk+5mb2/rup/thsRpQ9Dol4Y0XkJcvWKe1ALpWY1VYemVf3J
gqpGuLQr+SxPmXUtt20xtRnSJ6ey6bW1RH0AFmlsuD2zsxsqHpdc4wHxqIe+3Y2e
NXkBy0M94jGsJcej2Bop6oImcNm3epkuPpAo398fLOCokZ3ux5UJLGcjlbptzPjs
xEj+wLcJW8D6CMnDrFOStCq4W1Fu1S3oHuztbI+uZZ1lsa24kM+y/b63rX7llVkL
qefsyyxzkU0+tICAe64dv9KvSfsTx02oszR1pE5Z0YyxHGnHFKLkLR8upGNLgWJ+
DYAggAUvS7leh9G2CQkJS0pDEoQbhvEPb524p6P+2LEsENG9GdXr/qp0RCA3GNhZ
rEGjlviu5ha5FH68K85/OS0gwvESyaayd8s5EQr4wwgQk6qmtkymnYEKEvILULEV
nO8XGD0zDxyZGuIFNsrwuPDWD8klzdHpadCm6aBp2UrGpQ4kMW7N4A+ppnhudWfa
RAGovdpRd702XQNLxlPlBbfxG52zLhIk/3RbAqtk+uYsRnQfxmUZlDgrUhuny+dN
V9FpEZYr9ZRkbXiLJ8x+InoGAWUQczbvTc26XsXgkNfoai56fgTJ1FTYH2kcr/uo
IIpWn4zHiDC+HOf70uF+LymipApau+9UTKguvDP2lhNtbCUaTSxNkl9aIEV9m83s
u1WBVPYtjq44zr6Cpu62unb2ay4mLhFgpDnM/UyxBGfAWlckorogKM+ep5uDTYEL
F3RKkaXQ34Dvh4fH7or8r15FyWmS4B8VJo4Buh8mxpcRN+MNclb0w3LGeqSQYupb
WVAC4IETzR9TG9z0KymuELEiXM0kzyXJ2y1Q8/3HCRSjljrkzVie9XAQIUbtxZRx
YvpseHO+YRxTcXFVrczcOPEl1S6eA6bSsTu9f6pdlbY8YMI7s36nw6xy5pjiQ0tN
CkmNp2GVvlYNvlSw8Vnpx4GpARqhev4eUxV+7v2D1RVyO4Mm5fOO2c3bNxWPfBla
ln+c0hGH7GEOCTLvU2tjwiRZWEPb4EXZbfoXTgMtMCTMQAP75Qc62DENP4YMft3M
kiegKuDxO9iH4dlpNMhrxQNKocFzcuzvV6zY6HcU30znTwkOU85F0KVyGIsAKAXx
5sL55+1O6uoNU59tYkCSBlRYPXBX6DFPDz5Z9BlIIrvES5uKBWbZELCOo3M0Gspe
y5DFSwfrg+uYWQxCSOvPdS054TAZejSYMPehX9ziJ7NaTZy0WIA2ICCw9qF/5TTs
hkfIqsBjZ29zEMfhGQZ6TZeHjrh0dj4f2N1yJBytOpVV7tGcfhSiH/AasJ42TRHN
W0x/eiK1xkvMiGd0y2C+Tb4J97jdqhbA9sRCWiFXFtyTjVgII/ubHzirPWu9rR6l
DZdVQaROjimiSR0Er9BKo8rs46GZkfr4NrFX1retpvERrpFFJ/1NaOnOOcs43RRr
ar7TeREbWbc0/DDlgWRYUJUBSTf5r/we1cyQTBodMTPeEVHeTkF6dF756DoiWXue
2PfEEsz7OXB2eDMaSs/OotZE8ai6haOF+4WPiRNw5vvpA6xG5zPxECZJ5CQA0SBl
OrGvqkCMomKu8ecejoB9x/4fHQY6SUvSpXxtTDMMEIc6iUTjBS17GzMI4O0vUnpc
W5jeo1Ply17GKduD7IUkoJyZb/tkO7cznM391Mn6U+EtMkZAA0iI2LdK6PlVYsNV
8vkHOdBVanjn94R8rqYNfzXLlTbxc3gukzznxxiswE1Xnvf7E4ZJ+79Utzm3XfJR
6yYyKucu5mQyBs+Vyj0UzuqMcolO8zALCdSM0X4CkRLeJoWaYuv0ybrJadOkGBXA
AjSxkhyAPWeSetUn3MCVB21PYpxWp1tqrCeNuAqdrc5oG3iKw6B9IbkReB1hBKGD
+FI1TUzEwbL4HyYiqkmILr8F4Hbnzf4tzx9Mu0m8Rtj+gS21kZbo/dTeMKDrQdVB
P3lELEgUGeUtbNcOQeh9xPls6Kb1Ym0IOT5HryEKUWyEzz5Ek+pydSNI/K2KVkey
i6IGUfjc7J241avSXIrI6wMXB5IQakL+wYwxEqME5W8DMmNzf+ciMcRz5G/8olxB
bWZd4cvz1OgB96VQqEENJZT5PxUdEHcVyjIadqsQVTEg8WP0lHjtzpL4YwEc8/WG
fzrQKPvYvRTVVAfg4DzDNTRP18kSggqYFC1p1o4yNiZs0ZWS8vSI8kKj1t9qdMDb
gbNIJRX+lbqSWkbKKiyLG0q26QZhcqUOutYO8VAslXeNZs+UctgmoF1T4OCgRFGS
Xu+hsv8R5TFqYlqKF+W8F0qitolbRb/eyEW/bmZiVFhTqlhXvqn0qSVKNZHC/VxK
fl5lLM+jsN+rxDTCCcx8bwyFrlqmreJjfJ5h8vjlGb1TMzEwAfpIz7PXN9CfrUtI
Jx+pQFxKxFAdogSTwJ1grqE3TXYbdgWxcXOvSN6agPJrOtcG7QN9UbiMjeEdijE8
GDNpneJmW/3Ab6QxQsmbZDqcx54kilD4WL5pF/TY6mtScA/0qr2qOrGKDRnGfOHe
ot24Wls8iZbISp6gaTygHEeojxNTTalPa8YIpKppHLpT1ZohbxdzBT2T0XfC/dtf
lvBzr2Jl2HMO8dX3JNUAPz6ZHStXD8ugC1k8tHgxAxuI6EIJeg1jucJXIJ4R+obm
g+OTL0FlzQHKdsvHUBXG3XEch2kLsJwrMesNEX2VWW/6ML2PNVsqaRkMfm7bmfBj
jM+SQvgQxzec0VmvPoUnpI9sRz4qN2jirtQWX437hVxj8wAZWytkM5ZCvWWKFjsb
+cK9b+fxrhgYEOJXnko4nCCz0bu18fqFjNU+h1PsjrXkk+az+vbe/vM7XCemNIqQ
9TETQKgUQHhPOO/3+nlDL+mVzHN7q3ygdD95J22QWKp5eyY1JOwNcrX4uSyEqk+e
x2mRD6fgotdsehsLsMdIKOXte6Hq7yw1+B6CTU4gjLDvKcCMWGgPhBjpcy2MtPx0
PPza6PrVz1Oorie7PfUT3t570/qcCdAl3NRsPHQukz4drrGNUJRTELiU2AL2QCF+
wVMvVDOfTbFvYXVWcUm5gmbNSCbqWHwKVuPxm9DSKRcGCgvzxcHzsUS/mUo++U+H
hoFmFPSyAr+Rtk75Iu7rQ8YPg2HgAw/+QYLPGUlycdMC9gdV/5OL4RMWJnZ4+QeT
F8P2zjQp22G7xO3B0VqJ/FRuWx1zeSMHBJgKZgdhItZfEUnnb/vlZcMnXugbnMKM
PdyPZN3CVNO44LEHCFpNjt/rygh7J7qWK67msQLeTO5ciIU74k0g3yZYP2dzPINc
B8/HQJxl/rwFozClWFYjzL2WCtlVmoqEUI57Oxx5KomBGW94D8VBLtXngubqoEmt
UEnfgD9gdbIBv+1AChqMeeuVLDdQpHEp6KlqzHOydCdSsmNJxnUQZ867vwmfOh7Y
9+YWFj4Em3fsW2U3brFo/IjHiPGRZ+MNbfvi70A+Q0MwVbCgP6e9Cjwu+ODLH2nz
976fLQJ3UgiR4VuyT4ETdrDgCsyrDn/LTIgIgdDNFLXTFuc7gqHzU1nF4OZWxHAF
pWXDtI5Wyrj8QwGcUOYphdk9zwRUAGgiJUethHdPJASSgWJNv/JRKF/YIFqr7AIo
ngq7J6SCxLlfnoVJhdkuI2rNKvkKr23/730TrxNSt56hqvv4no5IY0zwquuyqyQC
nDR9AeeQuAYorMPiX5nxQKroA+Gh9C9U93Uw0iZxuId8HNvGDhtpehQ6fWEoKCDV
uEk5uxAEADVq/gTxh+fn0mmU8lkCVKxwHXJiBh08pkizWc2Gc1DAzMevUD9bhIEM
jpo0krp6tAR1UTuMR31r63toDFwR+dlwFOOu15Lak3qT8BNCKfBs6cx89cKIc0R7
lDrehY1VcLxV8oqCK1ZYdjCMSakB3zsGxgR1fei3e+OZZzZqYLjxD5oYJHapugAv
2UGxSxLJOWsifXeoYAjKBW70d2Gu4vGpc7MHjYAHU1UCTMFoU8FbPlODLkJyM1eK
lBL6wDdZ62hb1tC0HC9O7/gKcG1V4lyNreEo5f3WMV7QoVUwAi8G2az67y6XIDSx
D1XD50B/QMAJiX0Jd5zarvswbi1MFbFJBXc9A5n2nRA4KZDtRxRTzuP1sKnBrMem
Q2bRIDcCukb3HNLF68Eq3GmdkrGHf/M0dlkEGql3ohYZLwo+XzoTh+zxfD+Lhow9
iKZ8OxTaaJrvpLzKYpLfdUdv1GK9FZc2u93IdtqKKAQ41ihx+XxelvAoviNed1H3
E26/0Dc8P/qsdwnERyJ5XP/8bloiL2Z7GYaDfbnRTu+aiHmyrXOI2U2D4T+Mhwfa
9B/87C7ADyo+lZlitrFzyARtvmvBo0HuOVPQ9/imEjJyc1Envpp9/cNH9uRoNw0a
nin4+JXWVz9fDqtjlKGgBKH4DvpvL7pKHzsN9dSTGspxSY6ij9kyX/0yjjJ4Y5Gs
WW3WF+716/Ts8mm+Po1KritsBq4n8FPBYDWuoIP52X19FpJI6ywhTZ6qJvp5kz44
+HuYscp+kJ1FXBvIXUVH/XNBGCFxNGBk7pcES8rX5AlDKiFcO6IXEWZ9E6A0U3ci
EAcFFN0NJQ8WNUhxgH26vO0yl3hd5PXx3Zvt1ID0Q8KbYRuQmYOr0CsdDpoBmtDB
sHJGQu7wTbiSWb4RNldCl2XvORpDjSRlU/BYSbgOtOO0KzVBM5CJ9sz2k+wRBLJu
AxvbQeqOFjwBQiIslgykVCsWzDi26FCkrfSQE1t3YOSU81/Tzb9dnrjYmpyfSpDC
ow8D+eHmcw3qhaSyA3OU7N1xYQhQZCcgxge9ZE/ZSwJUZ9ivra0gEcsrEDdMRJEr
qN772affYJMYJ3lS+8fFl3ifD3DSWBqKk79WyAlTALx4dSaQ64WKfjhDtInQWPlH
MjjgR8l1WODookrVUVnLqjLIWW0sJbCSILNiu1h0m9DeLWP1aWzTfU9vapCrhZr/
nLB2ACRM0f8XWKq1lLI8apIHph2Yruu3OL5Jbw+AIL3edzQuoVdAGRxxaRVvSbvq
WiZLYfhRsaYzxfzRg/zzRT9w4crxtkn46sZNblKdYtvt6dqsrCBkxxgnq1EFtzUY
cY8rPDBRl1qaR/iI1MpQGITWHxYJ9BRoqoeXplUiftSVB3MDKbmvDCBq6KSBuTzd
Q2EK1jqdZxAPPby+u3zShm0lVcKZL7RBYNsy8Ps65mUAMimGgu4/5zFwAkQGwoQA
Dh+xPn0KUC0AjoF5pLdH3019MHJzr3K3bH9WrSENAB/zw4mFRsJSk8li8aH8peOd
O1ZvlcwUQnX7clcOxMLMP/9A7h+MWKH+NMCXD5mfGmEXwCeRU8EUcfTuU5MsF15L
k8acoE65rynl+G5fQNLYNts4kiIgb/Ob/F5iDS/AAuOMJd1iDy6f+Me+JY3iO/DH
UfAaritpDO7aLeq1hDDhXsE3MO54n0bNM5Dp+W/UxzEDvqIWwyGsuQN+GD0fqgje
2Fad+NfNXtwZGUZqJyBZOSckqMJLw7z7I1+TfKGNUN+VuEOnb/SrDcDY0nS+TKkE
TB44QxS43Ik74svgmaC5rEpcJRrqkFzdXqFv2yeq1ammwlEhIQ9wowtt88xBx6CM
rfz2ECNTx3HhrArDOYBwYKE2R1siqjFFWR3nMRBQaCtvTLzPnIMppjDkUuMYpxvA
BPWSNFAAO9AXAunIndpjJ0rCnZpsLmnJb1YMvsnxcmqbR5eC8Iw9sihctKvGQr1r
i4wItZq4j76UEd1+e1lBB7oZIDJe2acHlbXLWLDc1ofzDA9P59t2izi7I66kLi5+
qI5dkNCwf8YmtXCqnmYjyiTRgbVdi80mMZBh5VsOCFkfwmFi8M9z9jpHaD5BRA7k
+cLHN/eBQcwx2mTzCJbCVsS/Zuah3j75JuR0ilLJVeOguFSutmUhMv1MFHQ2ZFWp
2pT+/tbtENGCIOPWHWExvjCzyrs4HCKZriuAWaUcq3kkWzEy4GKQOQyRoUe7lkIq
Z/9gCHZk8gK6IO04kHPUyKhyJnGSrhRUGLKS4dJEY8feRIA1tRwbsjAv4RSeKkrc
HPjLizM4jT1s8bAZvyX9uOe3+V+yONQetwp/4vx4xXxSN7g8/8mwhzMRHJFVrjKd
VhwS4ap/4ZoEh+8DgZ6GXUVkmKYH5krCFSueVOg+K4h/0luhrG/ftaalyh/LbiXc
8u0p1hWS6kx9kPogj46YOuxeb+XYpPDIngOkQNGePzPBFoPZqygGM/DtXDzOsEpj
vueQ9Wk8OoG73mWxjSxZnNuthVRZMoVP83qAp9ju/ZhsYfnPVI8MguZLGFMSeyP8
rC5caGzxycGLMgkxHzVXXjB+VhRjxUgeTqTGOr6DAzBa8ZWWAtqrTDqds6Xtnt2T
TmpCKDCzb1jiQxxW6mtX21ZLMms022EDtHx2xPkQFbkfDUi/duoSIlyCemcSQ1Xj
C2ua01b19GwQ9MQqQsLreG/4CSUj/wiL/k5Vo4OdHF58hvot+/Hrbzmeguk5f/z6
SZbtU55ep9DBMuJptJhPaZKhELB+sr8GO/YR3w2PK4ZZLaqaveuCVX6kGmsM+IZQ
E1SduzftzCESv61vme9ycROCgHkx3IaJclrWGUOhKZhVTRFZRDGoZwpoVng31otv
`protect END_PROTECTED
