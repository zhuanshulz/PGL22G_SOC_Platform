`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FNMIFW5mevd8RmSdME8ozWSV7ql+jpyGX8Q2Ra3SvBulD3jAAyNvW0773aoEGjQF
h+aN8p0yGZInk497Ai22EPg1aIvLA406urSEKc2/S9SK/cpmk9VfiPY6UjZ0eH3v
yE+O9adzlkLfVjmvkskm8IOsT45A0IfotGkr3qCjwjbPFKFse0w++r4zplf5p+8S
vz35DZJMaO32gwc/xyYn8tmRdQGRu2hUgnwiGRhTkvq0cEYcG2uT7GK1/yGek0PJ
DM+H99K21KdJ0tfB6Qq5juAQfb2SvgvfQ+Yrrvu+roZiDE0bAcVCNemTmW4gIUdl
sQ0xWEVYymVdVY3BIhAyL7Xa/wwUIh+3Ul8LxlKAVyM1UlJ+cp44MXDBZB+Lq8gP
nHi5DCoX9nI7PKdd55J/rfz3cRlKeCG25ibeilyjLBkqn5Ik3n+A39ilvnN2Svv5
kbRCT53eXzJiMuG/6lvb44jSLb3jxyjUE7QdJ3bdEqKzhN8yAoPxCkykcQxEQ4EL
N9/sKRXtMXoIY/v/WvEb9kxrJOjXNtfeKuHMpNvYJaV645lO7gxa0f4EXx0uySfP
yUWRK1HC4/DKAvn/ZHMQTrH4WG4bDCgwhTlPB5ek1mA=
`protect END_PROTECTED
