`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bb48eCDuqk6u/B9e4OVQW9ZDms9zDFA0+KnO7BrB613dJTX8ARcTF1BEkU3/vGPk
9/98hwA/Zy4EMuvEBLyc6NwXE0ZK56FU9Aeou1fnhyNBbTH6S9XZREmrYdTm8TGU
tXrmcSTh8wG2IJVJCJLgyhf1Tz6+tDUQHCmxJueHaC8Ge5q9UJrZm/El4MhN/UyT
+OJUVZYs7Ejfv/xaiRZLTJhCnyKNjbPBH4AeoL/WG2Rr/Iq7LLG8bX4YgaH+ImsH
+kB8p8VdrIymB744DnH5honKjZPh72ytlghRpc9QdwcF6IW+22UEjCUZtavbGPFt
CNkl04WUM8lmkzQ7Zh1P73ZVFnYvJI+SK8WWPqs6pi6PP5CgnMBDkXCROfKknFgQ
`protect END_PROTECTED
