`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q27u7M0vxuR9AncxzlpVP/WRKrehJzBuNmbgR6So6m8uxUuA6Jdr07KCq1mBzLjL
p98iI0fEDt2qfgYRgZi6GQQG/zHfwk4FXz8PvUaFarsr/DzRfoUMt45VjuaOEuj5
VuW62TDrRZGUdcesOwAeCzSpR3ma1QJd9XhvFIC3zjDZhlPWQbgSxog9IBJmPONh
ncB7Vp5cchFuEgHZ2fldxPWEfGD6ZCFn6OHkyYaxtn5rj+gwWoojUYZRS42QROvi
NbgNRQWrO+nG2zNDiwDT6yzzgC3PS0AG9CJWgVH2g11HG2lhJz33dNYQ+2u7oTdH
rPDP9uXSFDcb8Pu+njIWneVIYxR2hMwOlw/OL+fMFvyLBkTiDRiCsd/ZFj2HHUje
M8HiBNzJZ2KsHqKCWf0SnN7TUe5uf3MtrDWAaW5YuBV2rDyrrSAKxADekGm2PbKE
7SZ8Lap+yxeK2BuvVnD0m038lDAapbLFrW5hQ+SmPTW2Jb2d6ldnC4HZHriW+inf
H3FOuYAk0yrxuqH0yJwB9i2vGGkCoVZqi7Hqixm7YvT0DUKtI48UlT5NRJHSvtyQ
4IccBYNv4Zp8IfY6tJ1navm1lAo26/As4fI3MwuhhzDwXnjlVi0zJXLzTAfDPcPt
JvfOAr195OiBh8VmlLGO5e8RXOyisNdpLED9ekJ7yy/hYarDCyHWhA9+U3h+ap6e
WQ9lSCrPmokr3KscWswG5WvxgJF5Aa91CdmuGWvexxCXFzqBKTa1/doax2zlqm+1
fYl/4xcFAK9EH75BHrJnxLtf/gL+gXTFaud9X/oB17Op81hP07lR/dMaVTyfNi7+
CGMCh6kVZFwsuUwD07L+JZQrV8jFIJmTIQTtZ/vMtUVYr/8TgAXVH+40tp93+P6b
T4SaKJiUYqexDBf46jFryxCVK7QhUTb/oKhVl57ysRz++xlNPmeuhwR0cQ0TwMOD
X2ZCDC/QPA96xUd5LtHMnrjgVs+iY44ISg0wOVqOUwsrce0Gu+fL+15AdRrArKQH
wUTTdEFowlXp+QhEhrfgSd0bKpVs/dy2BZUL5PT7mbRQoDGUd1BOa2xwj34b7ZR8
ksL616a2NdLBFiD08jKJM/5jJsL+j7iBgvDuIfjB49IhNoMoLkbiH7tbwhV2glzb
gZ04NCzFp6sclk9v6AhPvDk+vMA+iQR28XpAOyRobnXPQbBfxTlHQ/1T3e/uqq9B
ltXN7KHc1AIaR63ba3jJpKm0Pso0riMcNOzkI7SK84k=
`protect END_PROTECTED
