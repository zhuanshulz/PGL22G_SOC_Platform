`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xKVny+R2uE1i7CS8Bm4f9pLOgjwBnJYtmff7ZsbD+bsMvG/wUuoXj9QllV1IDeEW
6xLOraCi5NEN5weBX/5j3/gKQut0qAISJ2orpnVp4umsmNdP/EJ1HbNVCcd5uSAO
jrKe8VpQ97nYCThjT5jRJd8b0Sp2+r+7uwSDM6KXPkd40Onm40e3e+WnsArZUhED
7fP51N+VG5FEWx2s3nrdoawfSTozDQqmj32CCSlkFmvTCQlUmXjfYo1tPxkZoZYx
a0ar1dMRhZsnZlDyYCnR5fMNlc4TrbHUuthqC5OT4VSG9u7HV4l2zOpiyH1eZ3fX
af5RlNH+UdZImFYQmL2vaAgknSZlOUJ2XT8SzBzoF/1u9lrJ1NnrQRpFenVpE0d4
zyWM3OSZVmVUuQOtvq4BNjrtxRERGJnhwSMfBtD7DqkouBw+7YA4HXztknEJres8
nAPGTzSANiR9nLyQznXrHHnnLO/KjzeAoOfETrak985/xZ/A0YYDZ8CZqSKGdDOr
hnmzbDPO/FV/MAYdML66wsZj/gl2DQ6CfJppbt1kuXJ3vQUh6wYdlSHAPlQylcn+
/dIcG1z7pQD1IwTk5zIR+ZS6oV0er/jbAzpjuFgP9Aued1f4UQUzipM9l0l1kZ3p
7nh2epQZUe1ptdAjFK+URCSXZ/ued5UALgQyAZDDltb5oej/wtKpKrkZ172+qkIk
rqJv/3LPVcLWB6gKZS8yqj85KCDfNnQpE8l8bDcxhFc5X2g1Ir8Qb0joCAwt++cs
oBkX3XRF+4L94JEBzQTLCVbs43+NRksqo8V7dFj8s8LcKi9fKafZ5CXE52Hg/1PY
wY1VGeKBoitgRCSh6Rrll0fGEwBJLyDhO+q9LBOOeVpxIIrZtIH9rBtfcyeX+AoK
ltm99UuX3A53MIIgxtdy9kNNJhrw2Z/loDJgvdSZ1DWtLXVoc0aZ88X6iypvj+Dt
K043vvW15vyX/CRCUlhCOTtjB5HvB/PjpCoreQJ6TGLJE77WutnDSi43PldvLOYI
VibZcTnYBX4FFllchOVnKdhr6zhIzH0Hes5np88XfLp9DEoKDtJ46qBzlX8SQgmc
Fp7Z0AdQ/+wwpOIUjhDlqMWjiHCENKjBnI1Dj/zpuwu3WLjKGBdwy1d2utElbA3e
nw71frX43YnyYtbaOS7aQhVNHoWddtE6DN1g4aAD4nDm4VCnPubmLMbaF4faDyUc
kZXgejdTqT9mUYhF6ItSTekJk2PLSUp6IJ8OQiRdaBqY7wlLgw5S5PUC++ug/BWH
YVqSBQ9g2Ux4/A9xMMdnyJCNb2tvLJCmiCeHcKjnYx65ecNBb2AN5zZa/e+rLw2c
NmarU9OSAThtitUZfMfA/Yn3TPtWOEXpGCF3rVrFnamz7upTyx9BzCedlg8Cmlbl
izaE0L3eJYvZYuuDoB/vm1bJcP8xyPE/JqPsrhMlEuqQ2LHCXD2YzajiGfubvWPt
nmfqD4l2e0aomi3DQdJsKobwRoi8e1NSHdsDi0KSFgoJ1BJ96em55tbkry8B8+Kn
vr1fzvImFl9A1bKYugdbrKnv/eGQ4bEtRXZQ4hykeLmIqE8YTb2syhC3AOacnY61
htGlcy7x/c8Jnc+AJeAiVdU18KWvnajm92ONofo8EclF465L+X+rQD3X4zHI8279
M3E/RH/1+5ebj4VU4uUJ1799rw+Hyy8Q7UdZzH7STJXytuCLduqqlt+dVASkIxnP
qAgZr8pivUXP0x+JsxyDzPx0w2jNLmQsJMdTmolETx4f9WpeOUlvREJgUnrF4eE9
JSNI+W3FolaxFWmJnXz6sjUVLd6I5HDV92l2mW5Ncck7clFCbDp3+EcRio77xGYp
pOmAWmosCV2+g7ryElqlRuKcX0SC0LldtyzEDfZQP5nskhhrVlS/B8zmfBXYt+S8
G5SZBw+omHrYNaOWW4aQKdajjvS/zmjVPZdZ4ln6Gjo8F3cIbcRdljx61xs+FIj3
FluRaPqTi6ZNqR5z3eypQegZJkCBrQehw5Xu5CDvjIE2W0ToIxCpA9bQBFuH6j8e
wrKkE7rfn2GMLPKG/4ay9DTLvja0eQjW8zJMWZUB6jd4WL8pLAiBTgszULwdbKkH
ua4J3sUICAU/JRjKfjvDEoy6kWjcTORKzOPM28K76pQ3Ac/SuQgMsFeupHV9DvHy
twJTnsezUZyqdQsiIC+FTO1eJ9yGOyX7tHZPTRQ1KtasxE4B/xeItoBEvBUbWRPW
6gggfeUwLMU4N8lGLjjp7YIUO2htATWAU/Del7QlSDj1MxuQ5DhcVLpKG/tdxVXf
tp5GVW+sYtg2KfMfkz450a37j2w9dWzBUiGKNILG3nUtwRbIDJZMTjUr2Jb5G1q8
kmtxnrUpQ+62q4mxWPPuD8SU85RU/b4tyKJzk9GAR34c1Spn5NI3iM36zqwckGSZ
g39Kz4X2DE3+eLW67Y7EgRCeaQ0NFOgOcSanxeCsmvWt6IBUT0CZzkM/MbEBmGLT
y4Si9YYzcWdH6pmG0cbR4CR9DORsduzxW4FLfLzB6YBJgCfFOzlc+DD8hyz6sVln
+XcnSvadrqdUUwJc6gHU8oLYqpmvJzh+TLLcQNpWUNpLzNTTrM/uMkvf1Ped2r7k
t2EuUutdhTLyo80XK+68vnh3W8ik1lVesdr2Gmz9ZInMqiuMKm57PAmG9O7iwNcN
mex/Nc9+fTeAIAOzhl/82AiTUO2Ry7zWLTyeJgkTy5owXM/nGZ/F5COxBQPvd05R
TonCDQgWB9PgcYDPHwefDO3BBl9T5No0LaUVjcKcZME/62e5jACGwKeNNqX6yyL5
9tlVQvPSwf/voWAJESMjWHpB/3E71H9FixvzefP85ugE2PNv/YZ+T81KctKLmXIr
RXxXpFuQsrwmOuJkxAA6WnBcjcOEfCxkLXQyM5kjgXc+50o0/8+EPz6l+VfvJGv6
yYrYQKwFJprn05qO24RluheRP2PWJpVHLW9X9rD4FdJU4n2vaiy688PFNjgfusMF
vcRqEwSpSa4YVTddyLogAfN+7pXhWY6xm2+58OfrGsR9AGEUH8y5jNrfCN7H+4Gr
3S3mdrxGHpVhOhoRM9FOYj7ywjwmUKNosnGnMKokbrFYBNzunj/ch2InwXm6Wdul
kJNJDe/8oHU75PE/XrecCPljosHjn7c1RhHMmlB3VcxxX1VjA69KY3oAweOYvcxI
Ui6GTttijoaxXjOCRr2Mqzuigx+diy94FpJgEEudhEeBf1op0U6osXJ18+GI7vxR
yXMds5c/eSeVZKpi9Xq/qcgydPJt/8qcpOyrEK+NylwehlJI0uGhayXpZNy/tpsV
NEba+dGVzEpre1IQRnz6IIIyrT9TLPDxrqtOg66zrZkziOjXpZp3UXW5/R1QwF+C
zyNrNnhS+CXqXDCQt6G+MWOohqdhczIq3P2mSC7ZgnDWB+Q2zo4vKnee8rtPoJqd
HaVZ/xNbLc3jhwR7mgl6lKzZaRbG73VkRlURoQEFf6yhxx11Z6fng71DQmuOWPdx
qOi3GCslM9mpo/pQ61vaYGWhYtmbDJk1GAk81m2Mo6PksvydZUI1koyecqkhgSga
iAiZHV2bV1AEsLbCOf9KdQmlT1jYX50Voi6f/+IHQmjfbJzSV5LrSX6bNMmb40kG
QxY+YnicE1XUM5Fp+Y5VNAtSoec2vi4S4r3OuJhxUZZbK9CgL0kIOvPk4lQgMI5u
bE0j+e6Pq5nhvJAvwoZnIjrdmSSm7nyXMZZSRdVoeAkKjydpW6Gb/lDSE9aAJtyg
q6bCkcyyWZr9j6duwHMeps3vV9YlbJ9Pbgw44Etm3VSl2lnsGobIgxDxiVI7wVcy
BCn2Vp43a/lnrq2zRoeqE187Bz1E44+JLBCEdnW6ujO/hxGWAJbrvxrigK89W39b
hEAYRNtbyR3o310IaeXQwCq8ExaWiyVwEXD+0NP0CSnQs7V4t5yV+cxdjmt16IOD
BxXHf80fe4MNAKbx4I0jAPcs3yGiGM6cNRmGJHbuLXyVfTPHhseCjtTu9qLjqnl8
`protect END_PROTECTED
