`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xxDKgWcxuwUWy4rLEu6o9Oot5zeKllVA1Zy98kh/orpzeOW0fRFI/KMcDBeEvxAU
M9GDy4J3DNoJojxHwp1Gp42hx8U+jCBxF1BTnVRYWQxRMVdWCJ+v4EXGOXXDsDnA
3w8YVWYksmIKb0fS+32ioLd+qH6yvq7JcxbZyPPAkUDPCDET24nFSN2uJAscBIYs
pTzqRsZonHIQiiYx57FZciIGTBBV+MLi6hIOQM0fI+/FDOR5G+DxsJD+xdHyEg74
KW+nvsVgOb4XYP4r8Me/8tJUu7/aXjZ3eJNB5hYLrt0G2lpkC15kreIdJnP8Sm9v
9soEZ9f9tFhziWWfjksjvOJBsJp+QRhXUnYcJNfMHtpiV3hIJUM1Oo24rlWfWMjz
tF1nDl6mUZkNBe7Es3a2cWzA5MlX8q1bedkq0iJQFSm5bw/tbdBTyCih2RPAByRA
i8eE8DIUydbF7BcubFXRotHnhPLoK25QfQv14lTnjKzFwM657vdviJwRGAuQbzX/
P5xqPeiM1fHTVRrWCrBCDn5n5ttFzTN0SRWpxrvM2QwAMiYbPFrdNwx4TFRUchRs
yfIhwLABJJ9nV33mz1pLHf7mZLAtLkrstxinNrqryHoQ99aMqeHt4PXh3IBrVp9x
to663i2regbLysTaYPoqCcBqtS8RgMkU/AQoSK2OvqyJW4gSKf744wmcppnpO8CV
wgv16835T2Ji5Of5j0EPZHAyYFFrOsvQ1ROrwUFj9mwJy3Q8B7e+SM7ckf1A1Bv9
/+wEJ+YaU1o9tUUkjI25hC0enQ3hxhp3MrVUl1Qu0RgHswGniK9Cqoc6cWdosI4a
H0+wjRuseBFV+gQeoLAPScQ90/Jonfemz6+5e52nysMAgfJ36CCj3S1FzFG7h3x7
JMkzT3NWPyiux7Ycq5wCJRxoHsE4+90wFlM8ocuH95wwLmuJalD/FzHQxN72aYVb
DwCz0Cy3hMMg996fEPjcNALey2PLTAratOBwpF6r8iDJTaVduTZLI+RCNzLylWo3
HoQwPfkNStr7mWnF+shoIGXK72Eus6dtUU/ekZDOL2H3Fx/Us5bqOrzwtL+A0A1/
s3xs+St0lV3N2siuYeYODDpTwz01iL54ZxVDWN2DeGgswuZn5+WT1axpdsTsbrW2
7Oo2DES4ZmfQJ4fVbD7D3OS1W9zwSZ1e1EGdLKFEbFKYR9zU3JejRMKM51LocTIs
jpZNZKQfrivvzERy21Pf8cVqL7alnKsXDM4OOc3OwwvQCquZZGJP96Hp2tfqrXcj
ASprcNvt63XA1XxnC4igoirBE2U3KdtPl8XQWLiys9ZhL2hrbkrpqkMgLC1+M1Ii
xOM7vGqaH8OmmQ9XVhqlPPGi1oo1pC8UtEE4NxAH7Agnb6c8lXwB9qka5N3z7lcZ
l0Dqh8QsymoU0Iv5BgHcngV2piQ8rhxKADB4vvIBBOssZAdXxaPRlMt64h5d5sc6
IlAek3gGV3cFC2R1KAAO8okgIy8ENtumFW8JQUC/mLhcmMgP1TvYxx16Yes+SrlC
6MxyLlnvBF2cYGIFb+03U6A9p6L/1J8HK1h+L6jOAZ3fDqqwFN98rZL9iA/XEiK0
rZyLuExuBx+SMOFyg4PqO9hE1dI1OETPBylr7+UJ6dlYJSw3rZGsBwdfphqbGyiC
3B93w2zGAMfNZrnaVRPOd5MYDrXbb7CA7HtJIjDZ+EH3+N++4++6LrrvDliZZEz0
1GgeCjfz0SiICb7EEGvV7goO3TrMaC1lsZ8VXziyiHCijWgyGfAKhWrGvKNy2n84
vBgsBNDYbI/XFHwpQqb3GFvGPqckQz/dNhqA1SeqWurbfuW9pIOTFKcqoIEbsvA2
qEwm01tyuFpPQ3feNoCiPXCDkQBCOEufLFhaQh5AeRTELmD8a7QNysHJkFaEJy8T
FYScw0Gz8FLkxGVaaP3LPHQG3H57vTQv2K1rPjhidhlQb6iCiNH1QVEbDQh9HCNd
XCBMrLecQ0Jxb2HvlL78rl5t+qGgtxpunGrTUtNNZgplNn4qh7ihJcSHewyVwBvm
8s15sc+8wRrObzd5IHK8niagiAMB6LBguhvlNHIOBUBhpeiQcXIJBZsVfFnOhlfv
0ip+oOd2oni2M9lRe1vWxx4ghhJrLSB/hfilJrA4Qf04LWA/VO5Fu8legNqV9fsm
qSoWgN9mS4GRwtQMnqvv1Q4DzU/nHP+DvFKxGJ+SBaGQV1J7suxYVLFucks+tXaS
MyiIFtE4qE/7LB3rDx5sEqq8qPCwXdIiqB3E0lfNI7iXvEaZEaqfDg+9LWn+MJ1r
624RtEszTD6Af6uD5R7sq+HKRURmlQMkgTjxFQeWyD4jez3oFa0gK3jmGpwWddMT
enbmF2daa5IMpB5OVjm60uWZAFXfAsWZUn14rj9U97adkzk1btcIZz9LHyJeN2X1
SWBb26wdgpRXgfKj5pyqwvrGDiRc3KrdcxWEaDWurgOF+biA2bBospvvrVZagurl
oghaCEg8ngk8+6ZRbjB33R2Vi9jCbU2b9e+motixhH2aIH0HDg5Ie9CfIwa8HPyW
het3Gs7fp/HhC19dgBsjx/nHas/Lp/FQWAdFL8xKCtmQp+o5WmuHMB+k4tFHh8QZ
o8IijJgvhY0lrgNwErMSqo455M6ZAph7Xk1WNJl9HPUEbWPjnTUcAQo5mYvNZ4l/
sND4nzXZJurHLw/Jrqp2IX8GbtAGhKU8nXPNfm/GHRkwlBEtFlEJ6uH1DMUDdnIX
v2sWnlWuFyNbQG7G82Aurgnc2gffOJWkqYOvnlkwNMRTI+g06wtYv6dO/cSmrAmh
Zl7qjSomhE68ns5pkfAAMSwvsBDIgBGKYL/oLfxDA1EsWF9LB9UEEvti34IsHYNG
QBz599Wss0fGRuXS9P9AWXMiatpBmTBHLQiz6xCE3KXQII2O2kZckFptxbd7aads
XRNe29vMiyODNqio3/+fce7v1zAid8dkAKKbptCdTT6qQSFPtiiI3LzJfXOdTy+W
6hTmYUMwCA7TDE0cD3L5IWPmkRhETnAUungcFJR5xooniRHXyIksYlxvt5jd6J9p
q9IdfNIsQISHVR8nFYAAyA8kLsOIpPldKWSfEXfyeyquoNYIDn4T6ovUsq8+0h1U
jo2WBig5FWHZDsTVjDGlPVq3bIAhdHRL46BwtMWx9xil4aeHZ8XOi73+S9ahvEpU
t5x2NqMkoMKVSJUgADn4vGV2gqkLvszRD9tehCD2SCT/nfytfErUX/B033ghDJYe
7IeHm4mVgswFy/LCnDo0Gr8SoiIhqVJ2JtknDg5s336PS62cmzpb1ZjTu+U4AEFJ
oA4xImINqSrWUtU6m6CkQib/wocs+g3gaOB17qFKIWjTqGwV7sEzu8XOONxX4R0R
tTAzsnLoRh4/xrRqTEB1Dy+2CRVCg2Vu0UJyg9RCczG4v9jyjDQca06K71KeCoFT
I6audlI6sp5HRc26oq6/OWsIcxsJ7dJoBLxxn7eA1yuCOtOz36AbSgycK2emeb+y
2e8RPK1Uiv6/NguEjEanejl8Ic3sOfWvK31BnEcO6o6VxdAqk3NsGS5oUsOcR1k8
Efiqt9XZ06unC70cTxchmK/QU95CcNAboJ34EuY8iEygkYNWZz9qmFAuh8cuAGF/
UlTp3hSWf9JTtAspjasB6rx/EisuJQwvAk00pDfYgC5JIv6g/zTGjPNs1cuwV0rE
QA6Ne9zgi0feZ/xR5imxVmqst8BkflQENHIyvZ97Ys8gh9QGoRIaS6d987Q4FPNV
IWNwdsHFzcX57WTGVNRH5EyDpOODhoRTU3aPpFbgJY0Xwtke4ib1lFbTFEQ38HYB
/JLbfJK7Bj26XB/oXPJSfKr62wF0dhH2q8X1n5r5H9eWccznQrNGNPO/lWPdI4a+
658Tc0tLpUiJLpmNaqPEK9WC4Pe2hIOWj3h3kqpogzWttBaoRd75XcMu4amJuCDp
cMqHY24E4nLR7X+4r6TB61ZgcdT7Fsg2EMd777ZOQe49uTJBFUfT/9lbbXVDkLZY
nZnrAo15BamaITDdljUVdDddtKPNSDKnSdxRbGTkxHFYU61TAGltReI1f3r3LpR1
kP8M4O0Hg0hgKGj64m7c0UqZIorEC74+lpYa6ESwziGHoRuNOuk+lvgyA2trOeFc
pvplT5V0EtdmUbU5JamQIXxTzWcfCPUUv7LzHjoai4sVg5w8G6OyijGRpTDu5ujT
cd1C2g+kCSQq1+wLZGR7W9ZgBQ4+Ddp8oqX9nT901CxObIbItkGJ684bTT0IULKH
I1MUWWj7Cdr3sy+n8A1YsAIoTq3CY8piSejEteTwdkFpMopXN7Tqdilm01dBO+EP
my3YbJMecforc+Du4JrpjiUO92XaIptzCteJsGY3rmO4nVzNBbVE+BSlV+cfVwF9
uibdEXIoPxFtVU5zqTSlZngfQFOHnAGPDM4lihx8MEWW/BFau7QvjLeLKKCDhPjI
nC5GlS3s/YX93f+XjTJzo+lXr5ajtPJsE8hvjBga68bTE0Aa3haC0acnlkNNV2TI
GPqjdnnFYg1tNhD13sybyjek9VIomh5QykH89pZYLM81auIwQWI4kVPu+FS6f0e7
/MK8LFan689af5xR5P/FLMSptMURP2J3cBKc8qLW3KKcKLTQPlHcUlUkDt63EEoa
UOMy1E5dNqIQyRLTskW6rxPPoKlIeK/RgtkoG7yGCtK4BOrRmD4UZiT013uLQTQz
1qFCD5rnISESti7fnZYoYaIMidbp3grb/7tKIOWuNSjWIV1E5bhdfCd3tQse5o4h
sRlBhq+nDJ7ZfBavVrzRqOgzBWza7mvs0EYinF3HAq5geLNaQ50o/JHdA0bNAjOr
/vMFBWZIFLRsQlG5bLxo9imzhVnvbT41+N83QzUBuJCFoWrpFj6oXXGRN9DbxsV7
S86XhH8n7NL9FFY03wKDEhWnAtizBT9OU1C2ZKYn0U0DA0VgN45m3DD+xek389Ll
Hix3f2CD7JMRa9TRx0TZI68P7kTs/EX/QNt1R5sEgQKzs/tXqtUxE1DGcQooHIdK
WzShYniGJhmFs3+oXCJmbjgAy99oSbiGgM/EWs99M/wf1nCE/ndOd/ZNwnrX+12j
TnCrtmRliHeN6ARmC/jtNW5V5JZ+FsR3rHOzM6qEYEmfOHSovBw/wNUm+Eb/d1nG
QN8m7f/AXjm/X7djz7Eo9TsETIED80jUJdcrJH952v7xSsmoIjQsLdejMI/Ah90R
zTbUgBQUUcn/gqtIT+4HBSqsTqeU4TfOWojqLAh1uEdb14F3v9eU7k2HzZyw4fR/
xH7akV0LO5M3y2YBaoD2VJB905A7/fNR1p7sZkQFmQWZUAHSNznLTxekSGz4uQak
p/DitBrfxyhkAQAG0Ct0OJ0LG73ItTuipDFRBk/MBiet2mpFyvlnHrpDBzYNrrGK
hKDmSNpQqtU7rLTXK1kJov3B4k7DGzoQ2bqHq+ljDFe34ZCBzriqkBnmmAAxOGlo
vxC0OYu1xcBXU39TwLuZzEfFLEySB2hfkI/m66mDgZEGev9S6+K7DcLSq8J3ySpx
G5Hasz/jdepqlHHx39qH3LNTU91g7IeFylAouRGpvRC4mLMD00YSS/Pd9RVZR9U7
Q+GVWjm/B23T2JICLThz6g9WZDye2pDR3UwWWGjnTJzbAKkjwGKXvflFO93C5gX1
emYhTP+3uDgw9Xa6/v3sENNim79681j3I80pqxkYjaynHCILXOGR8e9Ltd0JfJ7B
cwpr7jxedwgldLkRPgAbeI0fw0e/cQCSf+wpata42rs9hs5bquCH2awsd/fyjAZG
0i3JRkL7/jGQrNROJ/vtFX22hMFpfnhe8zQJ5yvFb/m51psTixBaYOjaqAsbBg3t
cewIO4CGGRn6L9L/0gPrwqyXr9Etvk7qxHlNsUwZwAeXSg48h5beLkTK3yVRsyi2
bjM5C8/Q4Z/juD0XmQp0Nzx4PBDeVEw+UMmLbqtwf2/VfaDbv8pU1Qtp1AxWblVM
2H/Ow0uvJJIzHzWwpbM0cenanNb66BJrJtp2FldC3gqAaEvZtn0O6Muq/Ts5SG2n
HC529JdwTDlaL8sWQ7pCNKwpNBuuFvNpW4QxfmwNIZn2aGH6WHUIkCVLXo8JTzcZ
YeXp2ZikNhsSLFdW76AaIj8gktBpSM/d2Ce4Ht54Rz27VucWli+10W1VNffgtc4b
AoErMycPdGZhBsGEYnGNsekaKhMtnPLd5ddzBGywtUXXvxota5CfgRN1o+oSsBYC
mnOQh5agW5lSPGfRkLONoMyq6Jgz4ynx6AFDwOic6DC1pKUV12dRXcMiPLSM6ZQZ
KARW3LegwfTaLIplcoAx6folcCn/pryCZVdSzyW3sDDN/r29Ch2AUAwUcEEAbdk3
NA1L/ahQl4W4+qyqkVofCS6gDg/GjE7ExszOCOaXSBUsUBSH8cbCq3iDroTI+H9n
+bL3ydnU7WkKRrhIjjct4MBY+rRQPTijuq6mQ2UgZm5szaXAR3YrTPAO5RuSK3Ec
V4qFQMKpelRdH+Fj0GiXSnd5xGkngH9dALn+LMSAKFlnmozgG9mRpUPoC2jrH1ZX
9tG0w7KQzq66IJY9ByfsoZHZgX1+CwmzsvUmohd1XO2doWU3DyOnUNljBLC1fnDK
sRrvxCF9KIxmyfE6IIrzJkxj02o3eOkhbu39npyjEPlN/YrMO3Jp6jILFyrVLfxZ
C2UQO/c7VgZGwrwO//q5gry9BLcuZGs0VLkvQcFLmY7CwE5Jq84SoeCNPP6fmzC5
LB+jnlYYJ4KhNCH0Whpe7ZD3ya2/eHb8Isi7w2T8dfqEGAU6KNiG/7z4DxzL9Gw1
3rWUgY4fKiRSjc5wap7BVzYNAbwo0d/NFIm2/SjyzyV432jfOpg7NqhamIhpbsGo
EXcy/MXwFuZwnQ/JK6dIIdcFipI9awt0rnXMiToZldWlWRmvro41w7lOaI9cGWZU
GcqPxqW/dIZ6LxDi/s5sxyJR5Wbbb+4O6xchGEDZlYM9xDHvBcM7dMfSlMIC9Zwa
3Mgj9txGh6PnbsIy0VE6G/pwFazjiB4SHCtvVouTD14HSBl3RpLlT2TtDMc+Pm7B
VIFjzDrfigXnzUa5ONGjjoBwkPFc0G9+pIhOS9npdlKo6Aazwp9i9/NzIlXL7vHF
zKXsD6tnm32sd4atmV1V786Vllkv1hYNbkauWgsKnNFyK22Xy8nmakJYqGRkD5qs
iKwA6IlFOzLeokVAXTYz0Wm3DWqbJUH61JxXrjv3ZZ/iOZrYFOujE7FbRBMWizRI
Uo6y1Vhv9I57K6e6zsKFyvIaIcAbwDXBIe2fu50kknxWrcYAGWHGAXMzMv/zt9FS
P1o1dCwL2eZGV8p6lbqtvPIDVayrGcIVS9RSr9rr0Zklt4v3AapZpX1wNa+AbHHE
qoTm1yeAsyOy2EENF8ly0F1NbyAKgiyJKNtcH5q3qddAVr9eiO8vedohYz2m3Twi
e+XAr5vKZ1NaxYcrOAawG6Qvc2mgcmR6RHG1dt+Jl+al3V/l9fQa+9XGPaX7CVJ/
ZeqFmuw+NSfpE+GLXF37b7h5CzoSw3y063nePqm5zzAjbTbjWtoAItyVlwAXBUkX
srsgj0ULylJ7EGpJ9LvofKQI2DZhJxaLj4+UYd2d/zxphoz1myiiIDvgPb9z4hI7
N0/U5pUgKfiQB18liIBzr0CkjxjgHBkRbZFRUtMycVtNvb+dvGX+ep01oas7p+rs
t5dEoQQ5xoWeon3HGJWTsv8fsNAzw80S0oni8+hvRmqfUF497vvhJ8HU+BBC+5xW
6VKu8fyThNZPHg+b95qMAkQrkTReAfu7TEIw7nlXPZLEb5EGi/AFOi9/vvJkOrVU
c+NArxEMvwDQlshX3AtI5F8kqbXpwfDnmVyzA3FOou1jezSNDXMw0e74eB0thtg/
oS3ycRJ5FKukL7lrcOeCn7S6BR8zAwquow11KuOgfe4meu//5AYdgwDIxJ5pQYjL
Pip1cIIGvnh1+B8NnEI+S7GlDjrEqE+GvYpDCn85cer40fEznklhK8NLGiit3hGU
7TxldoePdK21AGqEun+bEuh1KLwiNQ/lQmw1cpRd/yMhhkFgFG2PjH0ImalIGI4J
pYyZ2vYOLRtiOzd+9M8tatwgwiUsX4iHrWq+F1B2XSQ/GqxyBlPc7UglYAhXUNUi
PqCYMafo6i6t1mP/p0yN7l5MzBmmkpQ7v0+FafpP7jrdoxYECsDbuFEABPbQdDai
QmYVP3fjf8xL5hKmAf3GabiGGHqoZXB56ewNbxQUVOqjrVcGlPv7gmTPKB0SJBht
MLRRC+esz8hkvQ90UUpJtZ4P8V3mUdI44IEB+ARq5hbvyxuTNYc0RAmw2LiPSoCx
GxLwsTjruyKgsZa64UM+N2Rc3ztU1h40mms7FD5U7fWG2k4qF0pvpuem3RZBO/nP
rA6QiFzf1OayogDEiWZOEkLsXdKNkGztTRLm8srY5PJHE33tlov6gtYgEU7G4Uq0
oollRw2FJ9tk7xx68PCbPvxegWsfuXqpCNq/4aMBu1DyAo8Hm1gHhvl2rz9pE88H
wFcKqij0sUJGyBGGeHfAFSf1gw7yBiVlJAAY77SwP8D9vDDFy12pQjldpv+f5m/D
ONVDWQq9d2r+uLbmX5Q1Ab1cIH9QssFhwY9ADNUbdUk/mZxx7/lYWZqVm+pJ17ax
RHln2XWky5foilZiy+C3QjZ/NcNWM/DuPX7TBlB/Sv49lnN8ooKN4Wh6rpqpsz9G
RTNv/ShLcJx3kuW2saGCIHG0BVmT01k2Q3XXoa81rZw=
`protect END_PROTECTED
