`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0EXxrcZE2hxpmS9QwHShsovbgA0eXdukoxGqGkvM2YlcPAMVOQk+hEOlYxmex99n
w60alF9SUDhlopwOn0any6CylPFpxyRYbdOSAt67TYl72apv4R7M9Z+9lZFayH80
7iS2uwGAucEpySySarlCBZ5UBQR4L+NWAYVCnjffMugdqBFKqgAh6+NkjojLlCBx
XheP6TbXdAhnxOwYvNwPYhuo3+8sNss00uheP8gs+3uxh9mswHUzJOvP/D5XreLx
4vmjSA8Srq+8glmw9NQxDzMFO2ErBUFCL+hTReQx0OzAT+n0OuuXyBd+rLVYcdoF
30InZfSWxW/UvGTFwqL0dtqo0ydnnFG3RW0yKP3R6xtLkr2gmN61amBCbuHB3WXs
ewdpZUHhLqcny1meyUjyHP40TF4IqXMR/JpUctNh3zeFc7bxEW27QxHXxD7oE6Pj
Q+Byz4U21J96B25KNgKQFTpIMiE1BX/il/LAhi1+ruyONQSKNIeUrPQD9wQvBOKn
7vlmZWa2Lg0juX9Ftr2NEamheDYjvkYxEt2ogSZ5ail9rQMh5U3+rB0Zy2aJHbS+
8uy+OaBPEGQQqfdsuB4p2H5MXPYnQVGb+2GrAx5EEPrv4TRIW442Zz7rC4U+bs53
7lnlxFkdi8f/TXYanKk5jKJRoCPDx2t1JsYHwfuJZoaISUvR6eLH2J4O1Oh9+kYd
9JG0DAgIcv68h+0aV23g7YOQR9/zg3qdjStkrpxTqLZYSKoPj31c8OEOPsynZPWU
9IzsMiYj/UCNwI+mJTjBRaImBqGwg62eMm9io0ORWT1GuveBxzib05lTZ4xb5WN4
48yRQGaqjXkwS3GZ4LVjWgYsCb6f2UJaM1k2Lciec3ECv48ZJv8jp0AAaaqEgpcb
gKO2GymbD1XCEewIRMibiyZ5rMOfs9QavlaAm/o5Zc6bzhZuSRcHzKyTKn7G6oYc
jtCT4MBX9iI+TcIR4eHVZNN5ulcR3iVGKpXj7sG8hDnd7rkeHEFwvpm5DTA014uW
8iacGneBzhAEEUdtqM6MALeAmDHnrvEvRJtNsDu3UQ/moSvIo8GP0yWtaj6xK/dN
7ejbQ4NV74oaxEmF6cBh/v7cUb6clnQ2pW2jFdQZTnpw1JbTD0mPKl9iH1UE4q7y
9YAuVZeWx+ebUFRKj2HyqCW/rv4gaXcnX7KRZOZQS1AXjE8uhfnYXuP81aKnOP7F
uDmbreDGsZ3vYQ5lyz9odXhNUFx7K/DGHq5w6la36vXRJZ+PPq2kRZ9l9h91GDB2
bKaWVmaWl5LhllRA4Bd1Us+AlaQkP730PmuQO0Ke0mfqDiHGJEYwz4RAFRzuEnPC
TUIUlLtWWtS4uYMYP+4eq7lnN2LoO4gpol7j/kIDaIPdDwEyNOrlNZ2OK97uHgRC
hNAifGLjrAJ+Dz8VAIXR9cGm3FoKyICc25u137m0Ey9zHTzafmAAMFmWBL5dYw4m
/1SksfDL/H/sPZwXvtkY0HHeQSp22PuYhqqlP43NkjQG0dtbHe2E+UKQeEtgrqgy
Nn0HslBeD4bQwL+dD5DNGAF62mB6qY7IMRrqX8yGfAi6NIX8eNHZkEfD3rPSnFHD
OCCjdUcPbvEuo0D6o7TcFJBHkAD+14gQclb2lDiTPNzxnpDSVuIphmydyoiQfg/j
ESmQzkxEgkKU+n6JtN1qHDpyz+GqqkbpQiB/Qu5QOH4+SiMZ7WeJ5kyQb0FZ0ufX
+T9gk7Jf0wZeH2RWO/EMSgpRDjDWXSIC6MkVyKosSnQJ0ULnDdtpto8qWGJc5szs
k8OQxeX5xNlJIGkhdun5XKIzaI3fAW+n4ldG9ruIvP+dUSLmsBRFpYne7cxQ69Ih
3Ofnsqwm5t9J60QrGJEoUW5n01tgQGX/Q7IFvScnLtHjt2jDwWq0OPVrwz0om4IY
4sh4vVQ+ctwwZUVu9IXt+ZnUbsg2sbr+MH2v61/hBD8omVe8aiky8kHcjhF6zTDw
ZcqILT7+lGwVdLSmLqZ8dVvS3vVGIpIoZbpHabDrDjMhfrG02/qgG7++b0goOvhZ
4Gsqy6pp8KTOMuUYfOnAdgPvVdN0msnKch0PiC5L6XCnvE3Lwx0d9TQ4XkpRXVpc
4kwRkY29Iba1owoa2OoykM8FT6whcoPBgX0GvOq4lll/GLwMAMqOdxkPq86rZ9nV
bRyRCLbApT23EH8LSL2dzn+PpU9zgeGPq9npF05Al+3DXuCKEOt+EjPzLe6O6fGm
PopgfsKD92yj3SqPVANKnmgAgzUXyMMS97ErfZt4XLYn/HUM2ET/aam8zo3Axsi+
TxgZJm3fM0YTYk3PhVF1aINXTXTlLB/eJu/bMaIuU21221XNIOYlBDirlut0FKKT
ezll+La6eoT8do1OfXUXkCNv5bAvkYohRFAMY6kq0fzNwf24cPFgSGIQtiGQerTh
W3css5BuBywzWTvC6eBncYrEfQq3PH/yTlq5xc8FmHPa4/cj3xsSnzz4Jv9nP02G
EkZX5s9KSFKqumbkSYKILZOez2xaos/bhaJiJpih/mK+QVs2nbgOKgZ6duaswUol
Ibv5DsAxVG2BY1z0fzgU9ULxr4+LPfff3+Ot2Ul+4R/eli+r9czlfnEEGX2pTFUg
ntvI2OcG9UYAuUIr/zXXM6uLuHSNzbapoT8KCv2t9nob/1duX1BttCz94wpPdV0y
OST/D4Wrc54KPuKptIS54sZ632Cc8ncnLhWOSkfYrbeCrlGfGMqou5JxWqNbyZr/
1BtN+YEfZQ2WhJVwmkq3TsmPBNk/IlDXuEfw0ZCJ4nfsqu6PxHkRB9X9GY1S0uhF
pGf+MjLnIQhOLsBrMuE/OaMqU0LjsqpLkGLRM0x7dEP24CQFw2njmPZA1PqITPfh
ebS/SkD2ikZWUy8Ob6tp11Jv2XI58vFu5VJDRhX+EOgZzYxzda75/M0y5ZzJZD+S
axX8dJynaZSSN8FE9pRiGCk3bLCM3SMB/vJsvAbpzp25flXq7WOQLIzajJklXfMH
8Ub1FFrxr0iDfl6UhufV3ztTjuRxG8PMab2gfq2JdtstnNSr/lBQ/1krpKXs+UCG
hz7DDnioM5S0Xfm0r7C8E/lbJMR6ZU4eisPgoFXtWbHjLPA4r6XrMHXIuXiwmPaA
d2OMWnL5JFSYKC5KYm+HDKbLO283hjercdPiZ+dC5zyDx1+z7H28FbOztv+g+Qbd
8IpAdgeicr/TLBrX8360UM6AQ/D+RUJnr7DPYAop9JVRUeGBotEdF0o+bIGgXcgh
i75YkFSYlD4sRs2h8GpLdcbxrcbhdm4Td8Odg1r/yOm5Hy3utgQsfktYFVf5EYvp
F3tZbcPkiUGFaOqC6ssavlhXTLB2r15xKimyWg+bRIyJzE6PcNqLWpv4JapMahTD
zmTeSbWBndUly+xl3/yzM5NlyfFkUihkipR34zVHoIYr3ElexIyzijWsRX9Tlyb4
lsb46u+uVHPQ277M6HOutNmVMiqB+wGsNmcSNXEopOKAC8cLxwhQfscv9hHtdK/F
sOgoqPn8Kixpn+/OLhazJVYMSNVAVQIBwCt6xXZK0gR5wJAErmOSm3I21i3S8ykl
UIIiIYaWdt2GgOQ8v4OvizAIqFI1OgzJftBKyiPr30V/OD804i8chTE42Q6ASjSL
mnakj86SDj5BhHdtXGms4LB+7v9oAOMg1QfQbazfyVURS2MckEAnexSntKlhSI9t
CD06BgXS1BbPPOVmhBaEEZgYpWEdUwQNb5AaLBiSfLOQCLicRnTeJGdnYS8I9Sa1
V7sDX/qLXAs0wPzD7Qn73sprGBaShV9HxBIggvbEdjcLRodQN4VVb4KDE4NIuc13
8L38weuA73li4DQcFumI77jXW0xSjjQ9cBa3yPOJlL3IOE9qfVRBtRCfiAIaukzt
tLbB1rzgGjV/HcRLGBX2eLX4Gs7WVywtREIhRSjJMT/8cjY3n9j2yAlVxeYCxTDl
MMWPxr/du/xDQT1A+NZ5iLywsgGoFJup5W23TIlWy2ZQ+NXvrQafZtEbNA40wrY4
LpDRo8/bW0Vo5RDp3guMCbjWy3HgrwgdXxSbqYu9X1VzYQX62cNAbKjhVDUH1I22
q//LOtYkvZr+pZVA3F0tnDggROzeHfE5kY+H/cbyODUb/y/HjTqan9RzwRnwTS+q
K54kJwDPpoxBpVOswbyW2RSkTto9yeKiX+DSZAf1SVjI4osHQSMYCIKQAA/jUXXG
sHI+Cp/h9DZXBe+ghC2W+eOjjlP6SUhawSqdGdX5SjHCYx1eYOZStVR9+LrxpxmW
LsH82mh8ZtK4l65HnSBkqCMGwmwrvxWxKCiXcn4B14Aslz2Jku8eJIy4vn8an/8D
lkzgE52cz5wBWXg/ZzGleGebHdW2zmM+WE0FZSpt3jcmD8wMUSLQN31HfKbciAEs
9HNNbjWeVApeFfoBjnNqABc+29Wfnj+RD9sRyJyp4ZIzMxBUono1KNz35Zy+Qv5X
BqQ0oybKtQm0GHJTrgWoJezOWGP/TYVmYEPDgyNqhNJi6l7JBFUlk/Y8CLeegdze
6q3xGx+9XbVEMniaxVwu5X+4hSTthUeZZ/lzGDjpcLH2SFSaIBiBFpQ/3XD7fI7U
qeIlHrUdiPUC4lLGXV4evZaixpXfOPQSEO/rhR5sG+AKgBl2vJoCWwr0UZhpZiOT
mwkldfXCgUuc2QYZMceIwFQEGKjayFIwcT57k6lVFr9MVWNpQOlpT3P3+/iRq3PP
wpZt6ZPyGF2JRA6LnFjj4usGer/kPdfqmoe/67HcMRTP6zkvSE/0x2iq6PB4nv5i
YUweHB0AK0HccnqRBwfre67LgfYfPWVQcbUsuTVYsmSRLt7c0WDlSudugiOQnej4
9ACGsXjNrLaR62ionzFiloK6a7PwRYzqrIcJixoeG8OZkbU6X1eHkW+w9y29wAe3
YOWbXl54ooS6vJT12H70Mjhheega/PEnGGvqO/h9ggxOal2l1ws4sKW9IsKkyyF/
WVWHxSOait9AshfATbl1qS2jluXPjt6KLIKFZrnDRgQiEzhRmtvMsEHfCBhG6scM
FbVUTUJLw+fQbXcEwph7Jd3CnZU/1cikEIyAz0VKcH4dhBxFVaNoAp75VsBqJHMT
vaW569hlCFaMKSXXQ8nvSWEnyC/WMwS+yj6pNjH84hukQ6P29FocgzEFGBY/Xcj9
wJ2Dvqk9/hwAuwydyNFBYv2WaDobcfuWo/fL++R/WcQTFEQHKqWdqfA0YJnKF17k
Dr+VRmD97UtOAp9ZmoK1RBXAn6sSWyMBkRWOzFGKAHAWJgvIf9fMpMpFPJhD8HZ2
qW7xZbFlMT2qzaH89V8Jq3ROWlIWEQ+q2CefLxrLzN/6LT40dQNdtdyRrxVVAp3D
jhQsgIJznNB1NDwp+tzCUA8U/4e6dUXdaBHHbo8Tqqk48etUvRGSNQy/+rigL8T7
N5aZg0Kxjm0DEUhVDU7JYQ3ogUxn257wPn6PEHMZd0XVoLAlNvBihEdLg24GScou
NgZGsESsc+M/y6nMTrTNfBFEL/iqaO3l9aMcPmMVJjceGBCMllr8MSPXyYFohO7c
7ESAIzLIuJvKYAIuyu8P8tpNBRZ/5AlUl5vVmgH8+cxVecZMW0rv+RnPBmKw3sgh
qD2UJx/uw1LS7mWXIHvEmcYWraeTgwmAUDAMmvVK2WYUgwACmV3BRK/w3rSTC4bz
7gJnrfBAK1paVtXOFIFU9mhHCzXieEHYiHlC6t9S3tAqDSG79oETg6d94Mlg/+gu
JmcWVWzcIYkddeuyxS/8k+m5Vl0h9B0Guf9jJdemIxFrPN3O4QiDrvtd5M0sOjOL
jB1H3bNtvze1I9WNXNjmsvqRRl2F2brGewICfXUh08vkc6IccuJyEU9LfMRke9n4
+OzIGmmU8f/9g7LLTumtaiCEQzHDDeHTL5pf26Wl4MnxucBqo3lzw9MRj1jQpJI3
G68fANL/VOdpcTTgMJQkp7W2N+H72i2pz2Qlt421lOT7gb/+IYTeYYZiHj6U9usV
Fkoa3hdthuDLOd6dnWFFTJCutwzAdAnC+WqIp9cDwpQuzqoX8gYPqk5eFToHtUoT
4hYSjyQX2PsezSZWtb33rz++0UOL4hqKpLV/S4GpnH1g4wag3ZkdJ1UceZJ1DWTr
U9H6iC+QC+R5g1lFUuaAI4KSOlCL7IVpO7lq/YC7fBva0i/c0mlCCqmgjyzRRXjC
wtDIE8gtuJQtMHvqS0VQ32X5zD0jbWC/jD1GKEg7u2gUC/sHHVNYacbfChuIxscd
SQivA3bxCe8N5STQ8QCCp+d8EIcOx/U+QLXJ15BEkcVQhl6jYcV61YwAUps5DehB
ZsCBjpCXPCKRRzcIBgnyxUIRW5QuGk3wdhisF8T8FcxzWthRkNdQzkRW75KVzHs0
a9s8YaZQhe0v+2AaQLDYG/rTIt3Eksx+m3Pyetk807w3Ekk66KUhnz8Cnvo9Y+Ub
tkwBOtZyRkLwhCBeY/IopM1fkYMBFXVOd6KtOWtRQ2yuUELCzdwRoJAbgwcKyAr4
oOfPyGysJ3DjxPc4llfjK19/EkOs0WQjaymvOhWpZXEvxujjAR83Yq5yUtdpO8SD
aP7xhtgx3I1/nO3roZL/f+2F0DPFzSKUm4Pey4aa1FZY6Yx1qbjf+7zZxFoQQf9Z
4l9ej9Am6hPKyryXqxAUsisxlyOYiN/S+ZzGtjQ/EtI79EUTQ1T0lo/sVdIeecPm
ouhwR5Ve4iS53NHrP9mxtkHK5MzuIUTRzX4KYOVl/8+gG8u+t1x3Sl5xp8uOO0cq
alWQZOPiafiPDr5GSx8Nx2BfCDTJ29n6IbIOdwjUPOcJbcREtk+YfhmK0XInv1gP
BerOj6CV8PwS/eHoKOVNXfcRD0QXlN0k8As+57KQq4fBkmpnab0O+JYkHY99qaOa
Bj48Don4bIu+XWj2Upx58AvQ20ut+Ti9k/BqBQfO93Nu+MHWw5sa2Xg/gXT0Nb12
2zuimREUBAfT3RovT+U2ABbH3rbaJR7Bk3Sksq+3rVAN7Nefc3G2m/V8MxBuhiTh
cb7Ry0TV97o140lv381NhIuBsjkyA864bkHRkQOubzPdkvaNjGYrN9nUEyBpfzIO
Mjh93m2O8aRQ9Jd0dtP1kbbdPbM/lK9N44kMGnoJy+Bv2vOFDNwYXSbkpx6nXbDW
TZcQcuRsstMogzhoPB1+Rh8fPVDloURJ6X2nJcFqE6MU9oPtuptWwbZD7BJAd87F
2PN1tFh7yhuDLuV1u/Hdflf9Jukk0U9IXcsv14iPARQ35p9d76j1L+Q1P7+WzTN5
BDz/NqbvBduVdbblyXO9/79UT198Y95AlFlmF5jEbBZIZoCIpNEm4JN/o/UMHUA6
IHrNAItXXTIWUz4iKc5zchnEpahTfszcs7lu9jcJDxLVNCw4KcB7au9qk94l2Xv8
BZDJcLxUfuHpC+hkn+960fjB9RK2X9cYfOYguDwKrHE5Ak4zGMo6SfXoTZvmlrsC
HVE/+CTjUr3LXNNJv0qSLoxU6qpM9PHFUhYTs5wct40uGVkI5C1yyvS7e2M0AGFZ
t7T4KVzNhiUNzUqKIT9Ky+tdiJGgOvSauJEvIwiaxqt6z0uGfJxFYIAQoEUczzW4
biMSPjBTrJ63LVMFMvPAFt3BiN5T2Yerweub2iHqVf2R4MdhHVNIpMpTWjA4Cuj2
x4wVrC+T62KbSg3FCPttA1ubRlM38cQhnl+G2pUQRNwNUvKZdwvlYwnm+AdxqhuG
QrjQxEMopmPtTGoEVd523EyM6Rj3BhRPVNcQcIUN8eu3fWOpxqygntlA7wqY8poT
PkL37WA4z7qo/dXQTvvT/L3OfnpJQurwyelaOzdnxUXx5jzt1n10517uwdShgNil
v74sC5eJhBYuXlciuiOUQo9fiNX1peAke2CViMQ3693MPZAyKQlIZ8HemWtr3XoA
OtkwbbnZL5olt+2K9vQqnxCJsQnr8ASaH1utgTGV0NtY5+XKbC8rJ3hL2uBmLp87
wF6jQbWDiy0GpjonkuIQeeLlMM1eJisiJdvTXjnnFb7XlYrT9crRQbyguo2VOPSS
XhStQ9pObCpKyYYaSQFJN+RfJ4f6hFHbLTVHJdM2/FhNlavPZQBTwrVfpkviXz7J
3kGIdVzO1KiPENEfNWSGKfZjpAqPRJYdH3qZoB0GUcja90d5lIA/qwWbyUOgSWjI
TakPgN9Zg3LjwABUJ7RGfrTPc1hT5L1OKr3BiOliplxWlOfBAgxzJEryN5Y/nEWm
5+i9g9pZp/7jutGmZvY40oceLQ335scDlyaS60POZ57W4RnhJ6UDNy6BsVf6uMl4
ic7+mgTej8oTX+UbwoRiOIJFKTo/kj1YEpGJufH78DMLY9io/UXxCpH1JZRA3ZRL
VdbZUBTskSBGfdg1zMMunNS1p16zIjisI+gylA4XeK5eGJhSRAnjN308cLnAHNAI
Z+DjxJRu9aLYJP1c7VYzzx0GCodrYf4IP0Ze54zw+kFwG4bhmgj3MrINyAcFFs4Y
uN+b30YjfsPOeu38RuA2PbfCz939WhyYRJh+2tLM/9Fb/rUblnBPCzCfx2o7GBim
DGAEqjo0ibl/etg/REB+jHGD7C1hwQF5PeI3qxert7Sd20FEdrYql9TyPIh6bMVU
ALtPT1sW0gFyZAacAfbKHo9QNiT/WMmAiiKfTgSO1PfgHWOYVtVx2qWI2lMP7KUd
FJzIeyRGHzJRjtK/O8ckFGimdMVui65Spdns2Eq7GE+6aclu0LYfpy3BjXID3HmR
/4RFiRwhqUIFyKhxTN2p0qV9Ug7MnYJ2VpNoqEUbQpNjBkIatD2VbhzekJ38Ox4R
mV8yfF6vgubiizklGjvhwZWTkjR90weqx3UNieGonKNbenq876XwqS0S7qzcrCQH
iZ+0lkIdX1jmDM+EMwOzMCbuvKhmwDtHXufBHtWW6nb7AWNMO7cHEHhJj2ohkPlc
2azNpedQIPdO265s0PbIhRf+0dCwf779N+rbsTcp3JqdjaLoqgG6BwyCW4sXzxZ3
57voEia5MWEwQlu07ibmI5rumxwv/SEJhx8dhyJtnt9hxQcwrPOVBHxfOBK0Y94T
ExS+LHLBSUR+4H9kP9BQdxu9/s+4wa1GueP9lz38n4Ef+txsFZiOdW/+fzhSsj6n
iaXTpR7+By5xRtMhOLoZSrbi0R2T6XeEbz3L37uFSu/n+CWEm5vpdcd+XLFRzpuT
vF4PVsfp90Iz0NugIOkLqHSbq9Ecgv+u+miXXw1Y/U/0pfLa3wr2ZO/qOjLNrHgi
YEJeqIBWu7uk0JB3rf72ylSdQGpAwS9XSXNahdVLMWO8EoiQGVxLK5Gq7/AyZGi1
OzSXZ1qU9jzTpHOpW/zIJDWjnxXQuyrvchop7QXgxB83G/KPi1EcLuh5RJYhNdOs
+y/DOtpqo9nzo/eH43ISZ7tr6OBSMZ8lmacig9himLLKd7WAwCmZ1jDTP8r2uij7
VcPExSoHBcVpTMDv3sTo5ica4tODWYWvJUbSn3pKiJAnV8jzu7EMEigOB3MIjFKT
tTgwBIEyy4OlKv9i+bZo+8hfHEHFjtPmkEFQrpjylJugIZK5lDegPo7yR3VnDa7u
ueEsUjb78U7ws4vYoLRqO/vqsIBRth6+xRYEx2ulwCbzxEWqGqfrb6JV+Y6xg5xy
c4QFoRNCvl6oeTwRZ3fRB3UCeiCmVAAtp/55PfL/2Dn2Fs+uCklwRqwDDaWFpvdg
fCmpnOrtAjd/jDYAoU3F1endr5jlRAq+jr6yDy8YL5SNfSJFEAX/UPYNpcAVNq7T
q5RDDpaMiut/mQISs3E2w/xmZVdHPoVYOI1QN3gbN6740HJ0BcFI2756ZC0Rn9Ux
wLPuC1i6cmh6snPLYc0DqGr16fPxYoyL/co1CKFvoJ2vNXc/NgVflj0Lc7Ft35L8
B59pVtvM3tWM42wZg+mdGcYtUG4bV7Zx4FUyUI0sHT/wPHXZc7T5ktD7vCrsjGNP
hy0y22o2iGS10YQXoF6opLDkCZp0M3D4KCseu9QYhAKVgL9ScaY5OH2HgSpTbDxa
JpxGalicpaoIgGX2uAhQwjWjVuwtjpA+pT+GzwIcvbZybuvzsvBJkl3tiNulr7Kg
lPtErlSvkVz2W1obqkercFAxi1Cyq6UzdCc4YKR11nK+/VC0hvfnjfmQVD5K31M/
rlBAB5LMGtDvf8cLo92zEitj8tbBX9TNs//Z9GKRZPRDPOtNSWyLwGN9c30S1U4l
OFo02YO+ch+ld+T46/bqURkqC0lM5klfmsN0HfGBAFzp8VG7EHdAAEsD3eiE7/SU
6TXoQgJGfXrwLdGc855mo5phfjc6qYJSm3uv4aREkJuSIzJtoIAqz+CJmRpwSHz5
NmUd1uiuJKOz/SiMellBGRmeYIeQalRf1UldjWhFyHT3RNjMUDq4znxe5dkN1zWo
6rvA3lXXf7US6HwhGlndnJG2iAIL4ROJsadw0obilwiSUzZu6KE85w9EiuKdlshF
WQZoOIapw7bTih+MzBM2y7HpwXyC6SK8iU/15WU9g7TrkG2kLB1p5liVahjsSOfG
3zXD7qWSRWQXLgpZ4RC3cdew4b3XJ9K2yLAKH0z1czoVNb6QBGPuY8MLlaXsZ2MO
OqHwGQELW82j7NJW6b/S5yXuxlrC6TeBEM/anHGMPGeHn+nfymolbstzd3qr/sHM
d7HIZoaF45myJQZSNsrujfBWH6BKJCnkwzNkedbCnoO/9rbNbHEvEJqyOQ0ughJA
m5KCkVDDJhA7U+rb4KoA6LF/DEonxEswQ/3EkyS8Ovc6lvjNyK7qSmKQhV5mgEzE
vlqzZtTeeL35svOMCJGXmE5O3POHSrnxYDSoinigoEhaelti0LKOkSZhdhTIi7Cv
JFHe7VsU1OZxb+cLwOI2NZ6S35KZ4eKtnDQh10TkfBNwZI6jUv/0BKvUPMbh/5No
ySomTx1SJrUhFslKkr3QfVywW/pWs/dONYUDaIcfAtw5K5/TeCh8Y/QUhVkQOAzH
yeGf5NLQMhjoH9Y9w0tDqbNrs7fLJqfMxID3EvA1mkTpqSLaGsaHFD1td2G2U6sr
h86AyBrxJ7oAgJsX2wkRsfM12rrLWGqHekP6RcsxdDzU4BPPSlSPufNEi1zMtaV/
FvQUbKk2xP6lZpiRN6tUn00K+TN47dK0GcIvFMTc9vrFwbXVZ3Sb0Of1du2LR8RP
r4MyG6WPs1eSfrDhP04v8IsglEkr4lrR6c3WfHfYFK+rzURX5gCtGfeh63K9TWTm
kM/sAvHAu04VLsLpfx6x2SfPE3XMt7c+aUG5As5EICGvAc+UD6/w4l5/iiJVBTmW
aevTOMvktXOcI+VGmgLbJqAOcoMSgaC3PlPETZs1EmFaIK+4+7Yz8SU5dBp41KSw
Lm/QorQ7Z7aQAjr6qQOaX4BHdP+LlY+eXqjj0lTxtqoLsxJuwZKwTYxBuHk+edwO
QcRI+lYhlcYcwgYFYcN3Ep9pgmHT87hurJMFTANHleQoFCeU8+t5whADrnd6gykp
qfQgwyZMMoXIQuaxWgfT4iDz7VYwteLbdE12ajy8B0DkIG9bSjCq40Zuezd044wm
VA13jRjfTDavTTdNQXcDCP4Uchb2FtPXPjTu6iFx30Atbs3OREWh0SS5hlG8jmYy
/fSLMZzVa452bxqYtCjrNMzCIr8oV78rKa7GjpnxNEpMm+d6We48UKjUXNwNYQEj
/0jdxojX0VHygXTWARcxaz9xJ6k3oZAPQ1L2e3XZd24rCwHFb4cjXLdOki+fNXut
bVXGFAimt/sneaUyNPGSsee1XFEnr91q+iREh8HsaR64qdbS55u0tXx+jhbrV5bc
6u81i75CDYIdLZzAIgwRHQhlegCY05ATk1RWSS97PhieRRI5cmSq6ycKwtfo89Kq
PH4g1dbpWLDxmPZFMGNnxyH59aYC4AMjtJamuneVf/o1PB/AVuLOzUPUKJb4ukKy
PRt6Ptgp8kvDRjIA8Iry6TTG1ARp6n2WdzjXFbKhX9KGDUpusLsbmnChRqGOF0I8
go9DbTABFlBedZ00bUpD7ZV3LFAS67WwH3hudh8FoQ9+XBywlfLVu/gs5J3N2aFw
HGpECLxpLArhdfD6jHb51ZnuDubOO04xYa3wonFzx0o+E6nRixNlZvkeGcR3ojNb
6TuHI9yy0kS5ZBylgJG2T8RXNBoNTPjvv/V7kL7JN7+7Yp7xQfDoUZQeFn4ha6Zd
dDks13qAxTjqd1YYceD1VA9v3pZrmF1n2jlbz+Om/n2DwSCt/EEupps4ULeX7w5X
xyRvpa1pxg+bCWIg9jjUXW1AMvExjXkHEJhynBNjnpzdew9lmivG/1kn8d8bNaMW
vTXvF2qftJpF2DlVpKLWRPr5sG2hUT8IhVo71cWOuGAvAH+cQmQKIcCD9igN1r4G
/rQe9dWqZSr0hGx9nRRUt6rAdWy0IsGhz9nj1hNK9ZMxSa/sNDbez8VEQrVwaME9
z5jlhxaeyhRE1BfWmMgwVwNLqAsMrxZMEoAlnqDGPhvVQ3eXXXnvtBTVLb8mq+vU
Cx5iSk6zF9PxXm1RtGNHDpGh4TFnX2XhPP84bZUh2kYS36cJYRT3kX4fB0lfUho1
mwn0pp+dYJ+AzQ5dcKCPnFbAzH3IMv99eEuSk/U68OpNGUjBQWWHOs4/KkzrN9uq
UpQGwiv1+RBjVidBUWxVTmLkqHiPGBQL3NWNmJU1adTfggjtESqRMPga8QQabPVc
4CJzJx5iOhvl1/bNgcEHpfce4bO6p1PZw/Heae5QMrn2eDyP7iwV7P/LV3qn6JSg
ZUcyQpZd22BMoN+mhYXMC1PqenP1cv7iGVb23vYt2FMdXuWcAIr4HCOgpdsae5du
7qrmAgDGAPxp5Fwho3QHaGxiP/gWRb2+7wgxEkvzgoOrsM8xwEwsHE0T+3ikSYU8
rTh/V2f5x8WBJwSHINDB2oGEFrrSdWUXR83CjyM1zObKBxV1bGZ/UolTuFPlbQ/A
QLHyFQkVS1W2imZnz+vW4xGaeO+svpm1DzOlTdeNPJxBY/mVO4pSy0xssC5g3wkg
XwHpR260vXZPzL0qADfSFa3IWfo0WVucjXlAx1CIKwZFPb2HxJ7T6WUzsO3gixCo
/8SqALLB//hznv6v37Nu6B5Db7ZsNEvfBfzloqBBrT4phTzmD7pQlwfvd26pAUf9
UaZwum05pIdiyvsFZalnwrIyvRQYfaL2VxHsJZVmJ/jOgS1iKXpVrQmu15kgADYQ
MT2rF8SnUWRT0dcGRV3nmftJLXX9tyrAwXhMATAo6Fdo9OUOc3zKzcJF8y0qrIuG
d+DQvh7Jgz31lhS2/IF1ijhWXh6rgWjyP/5QsUChx4lC+2v+Cwny1066w1ZsX1Z2
fDYprhEEzlx7tnoTYG7jJtA87w+P6b74i54qsR6JvXx57uubOtrMpdASf0gu/IMC
gGuBI0wzzroE9WNa1d+l9nmDbAjdISsJ3PoQKs/tZPJ1cNfgMhqC9pnwzVrjGi6r
5FQzoYC6SPCIpbNeZSyxyR8gryDxv0FmSnXycMq5o44iSK2dfiA0A3Q15zkcfFmo
qwP9Tqy9frSwF2TWOOUOQzmvkzPt1DupzupyzPj4ZA1CQpfXIT5HMs/uL8H/Djs5
5LtCXYXSByk3COHf3AtMHtiZKBx5uKr67csihOeFYpF9IzGZ4PXJzR3fesE2X1BV
39P35+mIfxPEWlUFiFQyAnnqbeipviofyskNPR3/2E5Tym/l0x7aGML+oYAW/lEq
zUOG+s3a5FNtwPQEZQTQo8HNa86XBuxqPPgxgLINWTXrZCnEIa2uWiz01/gqnjrt
abblUc4kWftXaoQ1avCDLLIhNH03/gTJ8FSVWfAgw4eXmb6uzxvUDHR3zq+na4Aq
N9c7laghJ52FNWfpWdfIve9Uo7BAxJGcAk8kddZ0p8R/zpd3zgdyG7J9aFlb9w5S
VSs8Jfk427NEu2kz9GkYSuG2jQeKUCBeXVQ0PGblxRM0spBQw6flzJuLn/uzLJOt
lHuJR6x39P5O+ZmdxWbTbdKp3EFPsFJx7RjaJmGE8/dupdXilj2RnFWVLSpjwIIY
UlAneAIHYYzMyk4YynxIpJ4P5HNjasMcjnkLdg8st6k2jHVXvAbW1fh7d2SX3Cr5
tlBUpZRMUCBUVg//kgRKj+n171E9qj3KOchT2iTNhGZKIbr7Uk5Ps+bNOZbskijd
yGDKPmalxTGByj7XrrKoGfEaO3HybS29FbjrYNTQYvvLKyewbuCEmBVzqsxPxZ25
oODBKBTedjIn01NaGy6KmYdgqJq+3/y9yJF2VcjTwV/E8PsF810sUhpjj3HTUwqD
nSdWx0fNiMaRS68Tf1HQ7Ivbv236JbBxF2V/BrbTNevPZuVUe6Dd8Sa3r4k8GrJD
Q3ccRy9vI/gByHwVvgwaAJ1VBNnPua//+rMMekC7zh0+r4jH52/8h+raALxUk39D
jtYcTeeriakSZ7c/DyzyXUjVWcD3AqOaVmmdUIJL5g7CGdTIQFDAvRGobOgG4cqB
oddV5m8uob4wfGMqbkX1/Zd/2iN+U3OglcNNUWscTBIk/8CCw1XlhmaxBb4UeuAA
ljDGuhfhNDf+2i7ziHTICz0em7UMmw5ZQ4bJfyzRciBFsDdnxFdJgUIt3r4E0U3o
U+NmsIFVopaIwEl0RsuJN0xazyjAiWsNEM3XE1Vwqn1xKoI6nFrpwcElIQAA82RC
3S9eLnok1HkFrB2NpEkQaug2A1rM7397ymb+G2vy4lGZC8amY7LhTylujThqCGwe
Yd7etHrRLwu3pOKm8RRpBvVGIwryMIewm3rpQ3eVof3pDceBpwkenlYuagPRGlno
7psTWTA7cPgmf2/vsx1xYWtnacKyLQn2RefiJAc8ABCKwfddSZsQqqfeNlQDDHEu
+QlZeONAL5hlh5etfXLKpl/SE7EowhfNv3QeK1GPXYwjWqNprJWZpVqHd5vM9wDj
+TaxjSOUQ78AbVSiVjk2o29I4lyja8nSUnJ89MkiQlzmlTXVmLJ59COHHcQ6YqtR
5hwnWO+aG8QC80aK+0MpoinyKwiLROaEGkGNrv31dFXmHumBP9JHQxQjm8Aahaqr
mzT4jOjZsZFMdTnRCrYdFIAILewbuifW1PZiaCexryvL8ohQql3jwr01mBIeXPS2
u6pxBblfzhBkjAs5hO6h4iMm0J0uyb6cZydSVRC2u81upF5wMfsFmXANtnO8voQF
gH+fTnkkDtJFapFdP+mDZ/T0pvQ76byJjja1nDfx5pCCG4BeF8zIZapwZhesZ19L
VKUMEDm0IFAHXRNCWUt/riR+51UiIe5JIUCefaFja5HjpndanTQ8sXhF8NX3ZY4k
I+f4puUEIuyFfd/W67dn7Ediq5oc0tGbV7IX3ep6GMr36dFkJb5NtkoaVoUgB0Rz
RTBxDSO+aJVC58eU8jGrxzf+3YGmkhdu5Hl9X0qlShQB95pnBGrPXaeBZx353BPJ
jci9ejwlhGa8QiiD3Qu8EGmLGiOkjta7DDzQSrwh3613ZVNtNmHEeWqZlEFnlPx2
tR+96kIlel3Jehdx/IlMQcEzGn0xPTPM1uNwPPdOCV4MCWrXuGywkS1OGn+3Xm5X
nh1BSMLriX/ML7EtWOUSCWb48mVQ+3W7D5uXlHBrVUnNBaAM5WmXuHZMzWoOsfig
YN1Zq4imZH95sDvwHBxGV3gj2k+NG6kTxzUk+QNTCjXQ6lLKPouHr+z+dAI4QL+n
0x0TUWFTJ4ymybn4FIkl5IgixNcijA2anXnV8X9DzwUywHbmhKe7B2iK+1oyXN9o
Lq4TJHexGpD/rZ+ES6+7ej63ZjSwsvGEwIVhGBdQPxORuBoUZTDIZwsrSqrobVaI
rdo1IeHPnZKJ+kOI6tQcGfDlg5NbUQSlCu8YonqJHevh0lRaAjf+pym2QFStldnI
HmXl342m82lRzT0jRGtAsOWNldm2VIY5yLSqU/nYhCKpCMvSIHjk7uqNOl2zypO2
gC9SUY3JFfF3xsxzOFV8CODHVaOS3skI6KJf2NIobCkCyEQqx6zJx0DPLYojT4rG
CZXvLnJjWqo5luPNnQNguuMcM1COJFJmUV4ambDCuloJ87te2M80dZWTm/hrhScz
TDvlx9wuVSKFOaoqGAn0hJIBxuouO2Cb2y+ut4NOi8OLW42Oq3teCyP7rZ0X7ooo
mhGz1G9xluyPJgbWGFZefyR1G8oEhJRTQ//bfa34AcENKwZ2Y1CNlXkS0vGw5Ymp
sFblPN7diGbvl9ulccw6zJgfTxfs/ZIRhy2OwyIdnald/mCBXRvVCGZhJwFKxA+P
W/HARe/5zGKvw4O7KZK+naKJ0wvpJMSUrU+FsSe4JILBmplS5ww/zFSlra8MLf6T
yncG2esnr1IOq4vKY7JWw6Xu1HPI879D4+7H/6RmL9iNr34tHbC09yF66P3/btrF
hN89agxR2cXolzYcZqcN2z9q7+EY3BGRWFlGMTSJoP/rSYJ725mLEQYzCCDOUrbO
jwNofzkJaWwIF8D2it2LmuRL1GZCJpZr/suduhtNWRhtzdFrcpOPUR3uBxAFTXZ9
VajoV6KnH0LFjGo/XZK9XWnEB5LXJSFzti6qw34zPVyqa6uCyLJtwNLdTpeBmzxu
B+JwokF16Uns7K0cxbYts7fUFrdNk2BFsDTWi33yUATR4LkfrkKfFIR0JjudGTBc
OzfBKttEiOvlJyNCP5uHuIrY863qi/TZS9v186OlJDcHNrm+fNtW/vhZ05bT6XdX
z1PYBZaKNjgT9/tMq7ITY2OcfCAFBqUlx7IswFmKe8v37G73D8f2pEv1OAGjeLwb
3uYglj7yk/94ZLClgHDizfPiQIhUb6uZ+VyFaERSJKTJza7sJ6mt+h1XG3x4bSBF
J6Dwyv8fE9C02j6tUTJyx7ExuBsOnQjIldBrjm5t4Hiq/WLyhyLfRzcWrbemdSaW
zL1Aq3pV/N3vmImPWuJBV4Vwq4zxjJfggWkP8xE12t3Lyo7GJ9eb9O+4PqeqC0Ih
TgukRBOYGDE9Yp8PGffXK/TyzavKLXot87jEDh/Syfno3LgSAHPuJO0D8Wo+Dk2n
9nlSx1wrrIUhqYMG/FbdSbrW48tsImyGO7UDmrmUQ0I6sek7QElbZrXBLmrYX+Hp
V9yc9P2zWardF49S3ncm9yCexZ71+oRCGLzIkz7KDkK5RemE4aAwFR0DzePthTKa
52+NmAJHF+fKY2UW6gWVJ8fGJBrei3XPathqG0wrlyDBH6t5V5IsYFVpv8YhCRPE
Wr3ykwfgpt3q5U1ZM48y/uF0Hn7M23wm2Hvo1jDpw3IqnjIz29edx+U0b9yFOmaq
ee+vh23t21bpa/sBYr2pG8SwEIZNgBIROQSaC1BCAat/AKbcbKuItF+5LKTssvzq
J4ilhv62UCTN763GpcfpOesQOJOGZVtjTT0gO45s/DClaPehKkS7voRyn8miqBp4
pqmbMakFUSW7HFa8ABHFk/Si1tc7t9y2q9Kh5e41Tcf0N33ddJlC1gOHTju+hj4l
L/1nGuGjPU+QeUWU0BVQxCxnfUoGQ+1o+JjPMfhzw7bRug/4EuAqrMva0xnZtUHs
cmk3JpQQaSj+LcfhMaNGNpZcycBSO2b35SaumtmNlMohFQiDb4i9zhY0TS+V+e+u
RjYQDqUoTojq/wUlW/VwJC21HthDRJYCkGbxVqupxSlnhFX9vr00IxpdTsnnhjD/
y1doCLlS932F/3hRw7foKGfugrCOMdlm9tLMYLOiSDDzm8rFCH1k9/JUgHoLMW6z
jwwaoNtfNW6K2XqKVB0XtTbzt4QyAQFKwci0MOjAKs8P+Rkc2RJM5vuQ7D1jiFGI
otsp0kbpqOBry1J5I551nzBeLkVNsRz4meWxaYERfNkkFBfUECM6ZPle+smr0Cpt
8jqS11kNyVDoPbwd4hYjiUknZllH0L34xuJ1JeP4wL3SfAn32DCaa2CmXvLF9V8N
0V8hFX3DThzmY41tjhJi7A5BUsgW91Zc+hjBc9mrygUhQ4DiIYQxix6IKLtcMJrR
kbEyGKAvt7RYPrlkOl2EVwbGiHURTV4z1jX2gHOXqO0U48oCTQMrQvgvltyrpLnp
qP/dyySeo/JLF/783vrA2WNnSYBQQS63na5JOXITBLG6q0tZjxjU5PfNfRjq6oTt
Nn5cYzqPWKPHLaI+zozm3lLXWHkTBlZZcG+Nq7IdKCxVSW0x5PLlj+QpJZUcvJcb
4P6LLtHLqn5CKiIoFRfk056ci17KQL6hMT/lnneAXtQtA1U1MONBx5N461jBqvbF
wTXcXGtHgtWPL/4fCqvD32t8gFEFxoUd2lecATVE0dJLnB29LCLuc62IYrqGJQjH
uHefmjZgbPbECO1kTUM3osIKj2hMZ45Z7k6aqDtt/XDhe4yFmmXg5KgucdtP0dlr
qbYI8mqo3X37ShlNrhkpEma6e7OD/ZAmy7eHqwk2jfN7ylH5kI5lMkSbZnDjCeZB
fMuXe4m1LE/LJqCJR5ehZZFpSqpY2Iln9mwRiueyyi1Y3FFsi52LstB9YgJPZFTX
FRPlS4+OdUorDA9FbqMDdDsDTPdxTmu0ebc3JMd0gPbpQeEgREWhJ35GfnsSJ4gh
30GGh+hiEdsaZL9N/YWWdkeXHzKa1P95aSbc+OOYIrCo5rz+HUJhoGIjBZk7iAJM
yb5QRMIv4HJhQlIUMWz+loEIF7XeGi0vqpk+tkH+OFkiincr/xkSSfa7SLBW6Aqz
LlHNv8vkf56JC/U8zEnWHtrYogpXYbLpsyHMFB+tZ9u2qtmWEk84hRgNVAv8Uik9
t7jpSvewBrnGeAjl84qNR1NzIfNSjmM7fB+nYx2++5/V7NM6w5VyVRofOGFcpg63
YOqwyTdULh/wBykYDW0x8O/I5X5+oHvcfJahsI9kqmD2eP+qQv19W77VIp9YZ+Vu
232TRy0+thyCPI2rH1tznoKQOFl6oJwTMIl8EneHuKTJuryknyPH+Bykj5HIYH1a
gNggVZPRcqMt5KsHLeLGWlUWfMdG/SZoAp1iNitExRKt/RFRYxaWJWY3fldpQm1t
ZFvq4ZoD/4tpo/2i3k2nN6E09n2FP5RBk5n2ExN/EmjMuv8SxiKh5GDAtnROyGMY
noAYuhwyzLUpcRY8Zz8N39J50IuDPF0dkg7E9GKRytiC0uYMgp5RTtWV5+VkAGoi
p1vkWZPFkKKUo8ZAzTKZmeP9vL2kYWBCJtOuDaTvhYP8Z36q+Ty84df6OPt+B4PP
TejwKM2wjlMdjkdaxZ1Pot81mentrc2Dvr4AtmB+X2s3mTgtXgdzQZY7ZlP0xVxL
jDjVNCCFtxWm+986LtDftaIr66eH+d/lSmrHqCnpIsQqi7b6ys2eIG1/AGgQPDmB
pNAYjhiBkrlBJMvsLBgucQp75ZmjvIz27d8LTcQiq+QV5DvwxsPfHwiuTFyQGPCV
kiSKk+NxgGq7H9sOqKR9LYajFkUmurw9KQdeuWtaU2W4ozi3Ywc/uNIlekDOiRdT
op73BDl5vtbIDYE6Je4N3evXu4qY17RoLjR0JAdRS0osjYLByvy0MJSQYHxPVGPc
WUBhQ1+k/Qf35Whq/Z/wVIdHhWZdPBPv4htP7PomKqt5SzgNbVKld9v5U/xwg/mA
k9eBCMRLvDIik0X9Zpav7Qn7IXsL542NdTUnm8JGDb8VC7gWaRgBbp5T6MkXC1Cj
rXA8AhHNSHLTCj4LRGNBJa8Hrc9jiOVB2drlDHVrZlM+Gr5yUI3/QhAVBSGqojeR
8zy/5FwM0NZyS4GprOPyXIsPPrbez5V0Ut0L0ok9o92cWjbHgtRW9l6kZt1K31F9
CNLONoHlKu0wT5so7pKdupEpU8QYG2fKuauMX0BxTYOrcdl6KpOUZX+ZAKHRI1DO
Xvyp1sgJKXS/KgUipzLExGLWdA1dNlQN6g9F11F9PSUjGVeqJaD1CmtRJl5NxEux
KldOrRvTw0WAKgmDa1pnZJym9fZh9gfnvrIyn0z3J7IkeVbDfRJCTJqAUvEVYDOY
DvQwm7RA29QGdum4XTTwFn9tHL1kpzcAs5k1uBVh2mVta5JzMjD+didSMKg5U5dq
+lfqfExKF6EEoV0I5C8OIHd0qeH7clz3Ye4mIP7uG9tdXrb44VATHPua0bNjVhdn
IfZo+F/HH/LoeVUYCFX4/J8WYmXJYcGmsYXfGpmVpZ33nWXtusg+UgIkE7/BWwVd
IL8h1hzVEX48eEYZDvy3bYMe+nJNyaewjU2tqi/YE+ZDRQNYSbMJS6HzU+jYxarE
gUKuaxRpYmMTGDGz9iBZeucI2oxQmK58KQFGXZ2Hypklh/ekFIF+speaHJD/W4tH
5MpBeOJ94FIr14JhGIr4Ti79Mbqs0mSeNPmHGm8AUgG4sn8ZssQUkxWV7WKuwZkO
EniRZif38ve9tR3tjdO3Ux+QEjag+01iqih+li+WgbKDm9GTW97jCiUttglh3sak
wKyTUcKXMTKbfyvZun3f8QeYwm7dE6hwBMBcipUjjuHgGP8PmZYBu8wvRhoAnUqz
7u4DisD+7HHwx31qNR0oR85c+mgTGTuq6liM9rVmxTz1j4QutaaBmheO809vOJyO
RT86FNzPfPt9SYhmpF1MMN1tJY54skDyvmt0zqoTo4d4WKMvrrwkgCkbsC4qO2+3
IDvrp8HwrUqDPl9haPzCcL8kwnPIY/SBQN9Vd0A5aJVOoZ5yQnPwFsjCzNHGZ0kW
Zv85NjAuqO47mIY3MEW7XnNJf9wJjfVKVcV55+oYESUKJEyE4p87zJFJBaB7pu4o
8dvPmIb6IJLmig7CSLhVVFKikLVDxUWHsF7s1e9X3KZFAtHpTIpzqGluRVtQ6UUl
mqQMI08aKbtMHTo7jSSBt2KDK0d9xnGW72INwPQm1UaZCEhN4hgmIct1R54zi6Qt
J3so1k58XzUgpXoGnK1hLeoFsTOQPGyFEZdn8SZrtnzo4FTOKYUUfUwsXnK8BoMr
1KQk+34F6C3/m7QJmfUMXW5N0KU3rHcno+15gaKghpXJN09QEqCPxHKpICcb+2FK
xcoa53UgLVit3EQ1QBp40N9QPH2K151MQto/Voi7lDIWP5nfK74Ajx2uadTPlaEC
sNW3GCZ3tvKcIHG5MSulHrt9qEJ4wyCLGG7EQfREp9F72LV9anHiJDJ9HqG5zTrt
zSc+VLfkWOk0A6YbWVjjPIgPyDOBFBoVEC2oxb1B+GqzlflIOI36GCArh7N3EaZT
LjMN8a2QKqGemo+pOjNbWeMB2wpB5EgZ1zZevI2+qlalaN3WT1tqmUl83lvcfVUU
Cx4fcxiZsUc2X1vwCxbITcBR/Xuhy76k2nr76fH85NS8Cqm/JoN+tHnUPuFImrnU
hNysyzUoBlaomtK5L1Lm7ZyKZtcOUGdwRhxm3wHdfDvRz90qQDK7KehbF3PqkwdY
I88BycRiemkfVWG30Z9DtqwEwqkWMz5CnQ/ftk9Wli0ijiIHOvNSsWNguNzdziml
PO60rEW1XCEI2b/Zcr9SWCZKizxeZX5znnKJdw8Bp8sV6QDVAM1gIk+qHAwxEEVy
+KWucYU1Bf79Cz3RvcXoM/KZsVAINB4tgZteVdKRGGHmai2jiQpCKTdgoGaX7747
jMo7BsjSHFAv4SeoFBJSE54Fcay7A8JFBo1V1uTd3n4w/Lq9rWZxbVnrk5deyml5
ZZFLE/cYG2oExTpwxKrTwZ0BMAponUMhNmznYL/AO4fq1+Z/ysAkmBjsCch5t3Mr
2H4/o8e2zfJ7OGdBYgKE5q8oDimR46emSskFI6pmMFu4moDlr3zNpEg1mEjQ+L4b
zm61rn5RaMghNZGgMSOO+JSEtTf6v6ScKTcZ5o0i4tMnjfLRpXE6rmk+iWF/BEUT
YY8AVZSrMzPPXkKXEMdZmKjfirtpBxZnqmsKhxJsHhEWZBRR47f903Qy5DR1qG+r
IaIdE48a4CP/JIGWLobmv8SWab0Tqb+y4GXPNP/o3a6fEBw4ZkrCmFOvMDXwg/zp
3hK5Uplb2iLOxRWja7HYRhedrm56EAtayTE0v49XaJFP9S+55Ddi8EOBiY+Nvh2w
zk5gwThZqZRV8mvyutCGIhAxRWJoahgu0LJykNVPWKWbVV5DQfcEmFjydD5KzKtV
tqRqX7PaabyGYAOUVCTmNeWg1hulrOBAxObT7ImbuDzeKbjNyYU1WtYWZY64Uj2r
u4sb6AXXXU5lMmUc1q3o7yZy8GBXcK8O4HvpY1Pj8nIVI9J0b2OCvcnzyOSyWUSk
1vgDD3eGHPw5IsYo1kveapcZalzKLGLIA2V74fXx72KySbodqfnqpHCUlwQllPI2
uV/YZhBZXZx1ofs0CHonTYcgXtjnCeki+nh0DB8JZf+9FGBMv/9LplDYiX6OcgHF
77VAp3soN08Ic+6aw3iJlLU469biLKs0ZWjHaKC11eqILI6iUphjE4+drm2jH/ii
MtFlg4KxzKBmkuPUwybU7fk43fkFBFQihMTd16OUO4NWncSfbwxgmtfm7yi1ahhi
U14is2v9gD6U/yO5N25/srIgSxxPLLcfjoXwoiA6i1mmgN86GCzHv7EG5L969ED9
KYjL6YiqAutdnR0WCbaOBZvG3CrxzSBe99xLEAMVu/QHwO75NhMR6I63TCJ1OyEa
DhZj759nLt3+oEGN7PuTCbskn3uod7WFlfZXJGTx67J4kLUxkdYwZnD43Sohj3H1
nPFRren9LStBnw8B2MSgU28NLTpav1/ndnjhDyBBla00dXPVrHAxGFSjKxzL+KM7
YBkSqdM34VNVbdHKXwWY8h51tuloo58SKZUAOTs/SSNYm0Kk3CJ+FElwHHTmUz1J
yZHOtfAyRtpxPGnn5sAAhRYWHYsxUa4/Bw6hgGJg8awijSSaFgmRBqGhF1LqVW0J
4xUfHfSzXF2AOUFaLTXnIXEzYNgLqzGqahfpWfNHhQlqRpiDde3qQbYrI542dSXl
LMiBGWUwKzsKA4IYrnbsx10URRmJVo+xdzPwOoM+7kPlsRo+GBn3EY/4Z3fUwRb7
+WV631oLnH45u8mf2r33z0UMpe3jSLLl4p3h4vfCXbEnbyz08UxG9ekT3qWEPGIM
3EJlmncIylbqgaI1omN5Qdl8DUQOjedI1j8Hip5RjFdEIdkuXb1zKB1Vv2yjFWm+
EMm9OE+jRBNt4mNsSIaphJ51D1Oj4Jjgm62k+KLhWSzzbFUpyy2R8tYbAaLWylNb
go9kybHSbJgwJibV0/g/yNE5eaJyDxMG/KKd573ikDJ/r9s+kJwWts44L5hsaZIE
hFFapCsOs7Z2EKe0vLQlvU5bSvjLb579edEtw9QaNnDgjPRXTwfLsfU5lyDbfEgp
oLhP1mcJmFzjhpYzyBxDYdKaumNlSe+ucljHVXAWlQP/bXUwHXrYFcQ6PZFH0O/S
ndnmpkcguD95ArW/C1WG3GM0K3R1a5jPg+iTVzOqYUzgJZ1Rhkppv4EyrRuaw9+B
JvTcxl5Oht1zPAsW105QT5RplqzbsptcAj5fXp/qtT++kzlIweNOG1nR1LUxuRP8
Z7ueemOYMbD/DPBHtw2vxr0dJ7WoXWeBO1glno1LrGDe/HpmJjKCIQwLmORR/F44
35e/K7AwgltYRbY2C8R7WKalBUGLZ0fG0PdvrEc/jIhbNgL37ZHp6kG6sFBEyXs2
cMIwSeWTv2VDQ3JYpWDZKIUuxUri9W18o/b2oiwdl+aKO1tFJzXOdaH5AqRYPu3L
JK7qtGW7lfcgckFe0pLpMQRY1dTq/mljn6aoooboXqhMAn/QDAW4shZaIVN52kIw
3tge6eVtArNlWcs0fhJ6PYaFJ82Z2TSGOrNvgWVwWFqMewTZik+DrNIBHIuvkSHB
0vZffraX6omuu7XqKGeEn6e/yIzQ8nxJfC5dULhquTawWbfS5kY9vWHpFPl2r4o9
4ccwBfiU3bq4iAxoIDVeX3mymdIJZtW2J21bUAV2ml9YvyfCafW6194elFyFi9X5
fLAvg/7q8mA+gXq03rp8SABcLX6DDNw/bWh/q6mg22w+baEF+UxUxRqTV6Ce+T4h
ZX8VGMMPB0UKcPxaUqhfABSkPPLuricvhWA2IpFnGxevp8E6V+UhZuFeYnUOxBdD
VovLRdZLqYamL/wkVBuqGmcR5CqH2luMNNL4/aEPrNXPpLJ34Y+ESFcD8a6dVVla
i5VO5TshtWokgAMgm69mudIjC3mshNdZEO+/8UJCT4qLtRpeyuZf8MP2mWXE5+tu
tWrWuGjSCUr0QX4kBMJyuOEUpEaBUtVgrIkWkFnJSJ4dz2Z/2OmxjyAFGdfC6Lpy
kzzNl4+ybh24bzub+oHHPyCngkBgg2gCKf7vfbrRbv91fNozLpu514wjTslF4aZS
WbBliyZOqit8idrMBbrhe/X6YoeeNrZ1JScruQ7CyBSRJ4yi3ri7qmTzk4yVOJl8
40PnWlExN5SeGmngqbWPxwUOvizFKv8t+BwXMo/WzQD/sGk9b+bDRZEM+M8PwMW+
Dx4046HgVrLSGdv5uMGrmGvc4mfxnfl8hepw1gGtHYzcRfRsCNrEP2EjqsXr9GmZ
j1gkDduAFd3SnFx1SBIt+mryfMPuzeaK42jjTYuGUp96MlTRjy2zyjQlH2bzmTwv
1Md+CSXUuhduCxR2PGRVv3JlhwDuUq/tQZtL+gBs8II/bMkE3eHBzX8EJSZ2FpEf
0ZzQwX1mKg0gVp15sN2rYQKeOVVo8j4PnrtymKCnsgiSCI7WmGfO9Kq1rklztpeR
jUaSNnZGO5x0srwFfEu/7/Nope6tWVshgdZAW7B7n+uV/Mu2vIe6CRjO0o5B9cQD
GzoWKoIykYl9Ctf0jt2LBOr2EmPgpHwmLF8H3aefmlBsVxNkGXLscxBJo6DfRmRI
K4brplFq4+L4LX4yn5BIjpUzoAEevUeGw624z3hMAsc6TDOeFu2AUIeogZTcGBtK
LwqUye47Ugl9IHeKKw8D4rAdW3ymfO7V7pmZoWL/GtNMksyhuMEZPHkKJWWoV5N+
UrVxhHOitmxh8omyTU2Puroepl+aRV/J3kVpGD5QfEmAlRjEIaN3GHpqW2W1+VFw
i+UrF7cmm3n4KAJxyqx5wcfF4M3K72Bv+G3f8l93oH0PzQkNt3vaDJSmuTp7Dj2S
KdTAxQWUKmoaOVvNm0ip5Ep2RsdbBaWY0LoYyR0FCSkKoUDLXF3uWyHLPNeNmgH/
2JS2Mo1ckBMopF6aq/uMEh151406DIO64MXdQv81cFLZrjWDV8bhWaPFiEJ/M3+h
wI0tC3r9v+V+iKcwnKMpSn6jH2GUPEwR7jAtAk7MMYHcePEc+7dUVRILgiTxYZmW
jQ08Ta6fRSeA35AcxYCdSp/K63Jm5F3wyV05na72zbYs3nnzKgYwQ4LY9ZCwv/qi
TKR6EeExZpLD66WeQjExl9KttJXUFp+FEZo70p8ibNwyclx3yVgsqjkIVXlCVcW8
h3vfykIuO2Ota+IPgWwHozjeSsc10tsAnFrfrjgHHV6fakr5nb8LQUbOfO45f3lD
muDJNVFN3KW2/uVFoHWylUETeDqFWxAXVYIUHNvfkBXXezJUvSPg6ssljd1p8Iq7
FokAqgN8nJGyqd3k/bCT81P9Z2j3ev4dAPBnCqIN2N5gz1RLrUGgEK8RFvltO+3c
t908RDPkFo95B8b1uW3BfbfO4pVA1FqH3T6ct8Je/GnlFFp7WUA2d7vP81yjVBBB
/2JZLcS477rQ8xI7khcifHF3mP4unNp739nke0fPYCHfNH4PH0+zp/+J/JPZUi5T
xxtYpQuTlDljxJxR4c73b1RlzKDoCefxKM8WqVcqURSHuBEYruzMLayshc3AX5H+
1RYxecjNbfPVT5YXX7Zj72acmX/zuQGKaGj9WVXHJjbcKfJ/al3XGNO2LLzgJ0jO
1xNoBedVkL8RzzGyQaLxYvUvGSm9VxMi/Rd14PQb+6ONWr/H1nvZ8AbQaoRSlHFH
BHRLVL9rJ0rCWqUwfGMoUesfDCn8gIAtk1ASgPbjU0N4pSZmtdOmpaj0QdiEB6Qu
HwCLZZ2qTgT4H2i3ZKsQSkdqL/1eAbUq2pEULIi31qDN/cXo8Pejwr8SzaIS6LRT
7r9hmr/l9oUT8t9qBI+XHVkphHoMtMjOD2a3payghd0QJGPvLlzjByXu4TikwAhj
StWW9uZT4AOBj9RYRNxEFuyQIrqJRikels61Z8k5vMOZQak3wouH1u+DjRUPzSKI
r/saEBl6RQsA0BSvwPnL6eKfjx0ucHAzKFYcK3aHjFYDF/ZbifPeQOmjQ4dhfrJE
eG66sOJ3rDenZPAYMrh9lRna7xUW3wgqPf7IZ5jzO+mjzmIwyD9FfxA4KV05pM1T
n/r0nHw4SSU8Ld9Y/oxyWNAgtbOehT8lh7umvE3ghYYKc1QOcvb4856rUSIUgls7
1ZMLnWzRFbpPBQ1GvTp86EULvVbFX9M2Z4cmerB42O+EVAL0yg+qUhfMP5m/0Sl/
TI+p0mSJH/X5HHokyxW/vb9gZesJmgig/QTwxtHfCI99y4rxLfwpJbt0eYHtNVSR
B8mEnfrsL9aU/adV3gXzQq6pe0AeF6FiV4vq8EvPgBaWMnQJbExYfcPnFSMzV0cv
hn7tLyGVrfLmifGrfysSACDRwR/nhq9CGLbl/U5hnIqjfZfiyEORRYfCplzvizu5
QfRHFB38yZ955/dOrAiZiCxDLYzBfNim0TQ2SlWOlqI1QlC4xHCkjOjSxs1WagOz
avJgXkdxW4N6P/5qtRN9Koo6h56LKA7zd7UnpsBTr2HjXSs+rfLQX9W7Iopf7Cly
JSa1HTkG6UP9VISoTciIKukFrTEsTOS1n0MpHgHLC7XBgTkC175t5QYPlfMTAtN5
F5rqxi+vrDYPmaeR0BGP2F9YTarDUgVHV0c/mChUsLhIYNWkZ0rak56WbzHRICsF
rRjBQlSwHAk3/EPMO6/YoXVfcxYJUXzad9bYnAMzxsW4i2qXhbITEynKwWcamZJp
rISyxM7slXxvcK+cJ8n/wNUgD2ceLOKwEQbkHX+ZmFCAcVDFRfmhtRGspKxor7zZ
ANM/Wz9psz50EW1DddXczsnkB/SMjJr61MI0wnIDLIPKQGGfAOHWGpY3AVte6U6O
wzGDMDGBzUpoCXswVduDLegwtHqKtMOGbLhYZQy4vxhNAMd1Rsr9ZRAOPwzeSuQh
SOoCW7IzWcRZ2fT2ZaUUnI5/p0vtnowKERS16aTeTyVCK02VBjW3rhekgYpyruNu
ZD2lgDifSDTgceSBHxnk3GPPR7e5FATxy8XAK0dCSXZ098j3fR4IIps4OOjVnaXB
48TXb9hlM+YLmWp13xWwZB1gR8w+o5efNaJheky+F422LYzY3nkmmpglTpaaMRj3
bM3BRRstk8Tgn+06d+HUoIqY2yofDx/pf6z6NR7TuHa9eLnV/FUT4Hz+F1NkTEQt
7sT7OyEcmSqZmgGvhqtCk0TYCQdNRZJbQ6vaN9EGLHwUTeiMaE0wY94nbyfIGiqS
BBdd6WGezwLBlefTAoqtylK8GpM8Bc4m5d/kT15LjFLrmk17IfAItv19AFJZ1IYa
ncTB0it2ytqjjIl9t7mcZ3B+DPiXBQJItNNte1qeQhcZGAsNFgBtpdTXy34ghBr7
EhzGr05+7RE0/upblRCzX5jaG2/kRkSZ/JoM+sbmhctkKKxHCdgKdUHcui7e4tuj
vfpo2FAZyMTcH8YJsfYXoWafCHBqwSJNbhv3nYvMc8qwpA/nGtVETS7+g3ekA/WY
E3vPYvYt9D9ktr7d5Ft9ZC2p7hyk3Vp34bMwNKL+yLssZZzf4jEvuPmbABbrZWTY
CZBKCoY3oVU+sNL1NnrLbaKN+JEQq5xPhj3IP+TQNldSUAqpbIusCgkEtWrtQOQ4
uVFXPdpIYkHlKQhHB9wcsx36DpUJG7nVwTXVHbQWlCHcVNV0Ythhtykx7QsTF+6C
BD4qfFa+hxuPiAm++WVmvTQ1XKpWGVJBq6AaGRd1e/CLrHbaneHtI6LOXRoBdza8
hQqQYnGXzLM6SXYzt4Z0Hz9NhN1ye8v6open9yrDkQ+SxTmiSJrdbxEMrU9yLzKF
CgXO6i7stC7Yt+Onurnnif8mpGC8hZ5ntqc2SpWG9Vma1bMnV+2GOpuesS70+ee2
R3GXuT2E3A/BpWXAy5rSInDQ1qIcC4NvkVlP97EbPIfmmjtK8+Te7Ad442F3RqQJ
Zo/8HwSNLAwo1YjD3WsI5SNJlj48qOL6O9eK9DYHXk15+1Z7SbzuwpPI/wxHFAwm
ATgFeo9blzEZhPWsztCx/Cb44wmH9oURGdaKYQdf5Um2CS1E1nUGQM5hJUGhxqNM
1E69Of3vtLVDKmKKoRyFoMcbzxr7PIBGW0JepIu7d+y9MIEusVKnpapajiaGcSTv
U+mozFqNYj986P5tJUu4rus+97zEQKrIXY1ueYbz616HFdxRr0gPqaKt3nEjPPif
l00F1f5iVjNQujNjQcwQZavHWqBPjMrIh4UCF13TX8e4xKuuavgFczHZYbLpC3VH
qoeGW2+MUZcVLMv+9qTRBsD9gQjglWnB8Ypdc7aZRJb/wM8Ippr5V1ysi4zsacj6
8zqdG122XRe8dVEC4rt53RGx0YPnD1pyN1ZIh1obQvjvV6j+bhIEZWBMXxqb1iNy
y7sShiaDjAhRdwM2DrNzuTEUzUUaUXzLIAKPyyIUWox+xu9BurI8JGcePauAJqBn
JoV97YeP5fnjEyM4s0SRH3GUr/FP6Np2gHxdti08CanzKEEo9Rm67ssFaxLQKS83
x4gvjw2AEShF/YRHulCassTNDBc6zjbyxUixJX+q62P0lKq2XXsZI5ayuR0kdF3B
cutKWlLblCqEF/EBm53b9PGHx7dwT7mMIIhMFULD7sdx9XOBm1jwHsFT20Ya2klU
WR6D66mXedgcgnsQPsYQ0xeB/4PysYipBEc+ek6WO2f2jHFCD3KxmY95yzBvThEH
DUaEjRfhf8eREzP9g6gh77VL0NqGFOGUN1+jo0vFFwRc9Ujh27mRhjV4ImBAEkOm
9I26If9Vw+s7Jx3VULpHgNx0Fx+h7KGAKnNHdjQHBwnxcrgIksvokk9f/Mxav5Za
rMTfocQkb9EG4Zy9mYBXAaa/IjJvGrq1X2z3p4IxSKDQy3i46iECqtVDGZ57bCrK
JEchE1iqocUewb9g/gdN6+9Ld3tQ56UDGHtNqRxl6Ys79mWdnnxuxDgelg5qgCM0
xtWkiEq3pTfahsjHrhkPO0FveR9NvskHlj2cPQm+j/mmtfeVS+GOOx5XLyYluVYH
xbstAr8fonItvyAngf976/s84k+eeHXdkLP1V+TsnWjiDLPDjchs2GKeGEyDPNoo
KBiyPUWu1iPrA05gX4HA7oIDZWdDr49c9+Zak6vv4VkCIYdF9w7U2mO/g66K1vMv
JtGu+H0ZWFbJQrt24ak0FcL/aWYLSWfpWEmw/vz8ckCxEPc117zIKYMNTGA6Anyt
OOKkyfSl9RqCq4+IQYDuVkfudAnItYmvIBGkByCu1EDmnj1/bN6jKm6moXKOcYSL
4d2ZaHGaEcBMXHF3iroH8nvF3AtPLvM3tnspIYqwQAjNFweuGm8Mp/aBH7jz4YBi
aIUtBJhjtlqKLFaLKXzBpO7rv+pVuwejEWr5l5IG0gW6rG0vB4ImXhFjmGPaJ0BX
sN8tyPxH6Jz3L7qaesoUzWpqyFvHgIfUZ3LGs8eC3IC3KmqV8KwQJup8/2Ku3k65
BfShzZmdwu2+uJ1g4ffP3qboWf5kax49Grb2p0lM/4kjbcha356b2e4J93lmiO7h
n8ndZiI2rnu3dZqhsQD3hW9/C4mCYRl33FufsmKTuCZ5XgwGU4Rl9UD+Aw5lzml5
Xbb2Ts+d9YR/jfCJRqzFd9hJqSfPCl7PgdLjOZZQOC32d2vElOBkjTpqKPy9c4Nb
oU8zLFgFRt3k54fXetJ3Duwpn68cvAUyOrlmbkcECnS/BZGbCb3fXoW3aQuBxYjE
HOJcBKGVJymS2kVjRIX3p8Qm57Jja3XIC31SWDexWWBOXESyBilMTa7IpuWbTf4V
CyEJJmnxTp9fgJmJMFemhyvzkx6GJoWlKr0Z0YjZWC14f2PYYNcQEuSQCLPYYDAw
KlvTZTu8BQfKiMZquMwEW9NLzA/ztCiXZD7zo1c76EMXOilg3Tf7FZYGsXlyhiLD
dAA2Fau2Cis9lscy1WhHyanGIC36+erk5+DfuMsfg8XSw1pGrr8YHYPJiHve7cUX
d9k2D3lGU19JAPY3Xg0BR5PbzC91heZA25GIytPoRgppb8LGZRNodjYfgNhKwkYs
o3hJulAJRrEmFm1/k5yhyaFip+AaY4rS0e4kSkRNzs0Zt6cTEO03Tej7Lvi2NHDS
/2sLnV3ZAyyb8EWXBPd9n4cC8OSwb8yQepIjsfNOlRaJJuLhwXPPbMYWhcsBo0nQ
dJw1g/hZHA8qXPiGcQtlkJlX1ZUff4mKXMtODlt42QBm1xiGPBkh4Wmt6IeO4joW
60yFbX1xjNV5BqjFpLUuKquvyl/ITby46eM9VZ7CDuYwi/bR/nq5KsI2CLsuu0uL
tLXpcqmNamosI0c4FoJ7ImDTL59uEnMwkhIYBWYWP2USkBJ+PXmo4MWWylcIHpMN
q2ISuzdQ9H4ULFCRxX7qYEOf94S0b6pV12+VwOWGMoT3uuKJvj7ppaI4DkUSQqro
boKCNbR2hyIO1p2QNFSYh8O3L34AoFcM4cToI/YG0x+5Bv0lkuuweWopS+I54I5i
es7+L37bOvwZZhotbTuWCBWXi48GnIEgjXhL/9zqDhcodvWKyGYTuGRQ9Snh43Wy
a7jVXan2O8GKNb1feuw1HAGEnn31D+Wohrw/j1sOvAwLAh/3zuYgeAQ+3rzg/Hv1
WoU2WFbK268iOYJacGnrqlZlX4Ubhpc5cJ7T51PUsevKWFy0A8b1309NKLmbrpyh
Nu8rRzMviaWdeNAOs9TLLf0ptd2cb+43F3ZOJ45W1pFuR1e3hGlwtwD7PP8eWycI
tU8ReFoyWwfzTydoWkhs1Qde5VtXcsb15HOjqEaAue0Ee9DVR1WMEItzWQ+UNS85
7Z4/sImHJ8EB5ZkBbUktew/WhW6K8/u1GLDB38xkGD4dB2uWlRzuEfwGAd0j/tRj
xfii1UAzuKGufomR84DebUQpnfVv0EXEGSRyR3f8g3LDX2eFoVgScXXZwg/uAAkg
2o5lSfqsjzFI1GNUr+9i8YIg9SHCt9KNe6GOA2nwS9EjShFczpjWlZF1nwWt8uRW
gFaf2QUSWmhK2x5/UAMBmWZlxZl6/Rokhz78Ge445tF6d7/ZA/KrbhVAwqHJ4GT6
LrgfPu1EeiBcyelESLDU1IWFJSEtUOHTU/1jHKz2dqtBPFOBRBQE2PEwli6pStQT
G07nPVapuwp3EWWLKMAp3cLY1lIPelqxhmm8e3ItZWb18n+Ro/lc0GuFGIkFTJdo
aLQ3sRzbJmC2PCronclHjznqV5dwLE7C/TDyWtwXzclk1iMYPnfqqLj3iBsvgvkB
P6e0A9gqMvQBCX/xOrIfV8r5VmKgXlNfiNeSfjhOkMDCj39teqGmRwC7pLjDGMCU
ZFNdTsJzzQPb89Z8Y3bxYSX+SYKwtchxmq5WZ/G6EnMoJjxtb0tbNvaz0SBSIa68
8OGH24642U6RG40Z5OT+UZ69tTdYn82ZJhcRvYyEhj3j8FU3Y16jTDZWYrq6kEnR
cAbQLjKl6i2C8ImNAGrSh5hPAVUEZvryHXIMH46KN+qMdO+KqCzEFsLW+WXuHnhl
WQmmn8WAU4V1n5IhsmiSVrWmwtaNztZA6w936WseCpaZWwBe0AV6rRzAqZFsIq86
kKX/kD7+LGhmbDYPqw2UpoJTc6V+2M3YTJTSlQNMPGaI3ERiQku9QJIcI/aUXIPk
vke8UlsWyWp53gwxKIPX2fIMjMdMiL/3sfQJ1IgFyHJIIaB98Z8i3sE9wW5FmNWd
2oYOiUj0auTCyERO1VTct9N6Fd/4290h8co51qHrXp3v68pVfUaUag08moIxjRZB
D6m3HBApMGtw/brEhpH76v0rSRm7el/A8J72tAfcusgZ2mziLlJGqyGX/jc7Nmet
B55bGOOohMifdOewFgWhpIy62uc9dw8U2aXmTrzEZnDUSdUtTVgLe6IzH2693Ggt
2QtrSOujAhLG/kI4uTvayM3AEpynS5xRyTtaGUk4VrL5Wu5lDxVdeTjuvVVNZ2HD
o4n8WXEWn2XV6k2aiwLL4lxo64rlu+uSwPytKsEy5fqlXurb8mCJo5en5c4Xt7Av
orGbzsg42d0deAs0Dh4HAkIPOP4wOwRtoSH8LG24wpgv2iCSIgeMfgBetNO7HTPS
Ldgf0b2/mIthmLwQWvFk7iJo3yAq37NViuekLgovoMTLBuSgzfU+MmrpAxbRlbN5
XPdlCAj2P13Nb1beQRuW9NcxS/mqdGHdj+M06L5OWTVgAk9GUg0yLos4iQ4wUrC7
icMJSiwI2aqYKusJ5fQyUJWZR2P80yFjl4j0dQ9oxL3LYEDEDrpH/ZZn4fR6Vnwo
eQCu3FH2/AWLxY57eyd3JXglJm4ORudMYKmc3U5jCtGSpBSq7mbtiwqyk+wPpeEs
LaXC4RsFkWnrQTjk3BjRdhrvirFlvJuX2IB5R4nNnM874VV39pXXufKCvE3xAowE
hCOE73A/AJmquTHhPFppBl8sWIpthWX5NWNO+X8ZltASz+GZUGXfMp+xGz8atVS3
AUUWavMGOFChXGeMlyze/Dl7jfJRu14fybdfJFcnMTVN9iAmZTWcy6ZCiKLlpB+c
2gENpsf6tk7Iie4Ty941CU+b/hweJzijNLFpZyJ7mxKgVR6Ru06/37+7QXBqKOSq
7JeV+FfPJ1dCQExj6HlaCA0fBeYPDTAgg9xiq1aXWQdfMxaf9vyWrwVJ9UXKlJY2
HEacqyGbjomGRRsVISXSLBwXHtH9pS/6pf4acQWowfHDKEkWJGqFr6PAO6EDTEeH
hR5tiMDiJA4oPnRzN/waWYFkFXowsYwqDx9FbX7+7+4vsXMsaRQC/yhcbmAICz4I
A9XtRFGaMzSguZHFRfAHQdWOqXa4hs80p5cWuYZUOQXnWxrAYPGqGwv2uOhfUR0z
yvtbpYak7phZB5J/vonFU4/3+VExFygwj3QWAUjbRoSrrjZzox+Ch8IevSGqBFwV
wJyjSPhCaIqkIwmlE5cM1bmWCuYbMr6jbCz/udO67O5XZamAjoYmloXXnv7RJTRI
Uz5tAPw/24RQaqrwJmslfp6TwOuVGGlkn6XWzDGv12FJjAStnGHF3nRZdsLZwPcC
3WVH7W1sNnXLygw7IZ+WiwxzQRilijNAHHaWeudDppf6bD3hOvKiuTEFNWdcWWBL
E9zdiHD78B9cGaiCGCuJl7YfIjXtUc2y3W72nwLS+8uoLbqPOjVjpqL5dbJxm1d1
GIQJU/70VdcQl0ESGgk7G3h0K9K1jaK2mSLqw7hJXNmrV7/rpyjW2DIbnW+ZYS/G
4XdYKb3kCdIdAYdt6ZpFWqq6RcO8+u0hAkpYRKI9agfq5m6jWTaudu1cVKDmXQPl
fPhSMs8T8Y6NQZiVaeMIynDCZhDdvMQf7wfDQ5zr7LOmA4d4XaoUeUlLLlgxjbEm
EqR0f1icC7EEEwJVPvSiFAmko5LLjac6AsYmnfXc88pwJB8kp9zpqNpGeizLHSM9
xG0rJDCTmqrIjPerzcHmypDmk0p+6EzCyUnkfOdtzz5zIA8gOiuuQqg9xIcbpjX0
jni+Ik85zoC/ehr74eaBsBbOeEUuoMdmY23FyD6lzhunYZoqZ3lVrKF8kPqH2Z03
dcphK2wcop7U3MLQg4MUPbR/lrP69vjoZT+IpnZ3Mr8rw+y+4yz3JvVqWqqtILWV
2SOzjl7M4gmJejoTMWR8TTmKHCeiAKonQJULhhQNTSUxAKCvl14kPL5Y/b6yiHF+
GvoyWSbxquG3ITdTgf9o7ihlALgGQ9gtVTbmfryywEXxMlwQ/tKvccWijg2nEpat
EyRMc4XtWqiOQjhi0Y4IUniOBOIpY9ph/EratxxRXfzsQ+6Q7ySrqt9H69SZrDL8
LCsnaRMuzw4pQp4hGTHAsuQxqIVw3OflorccbEwgmeP6u/zPki3hF4f36efrKpa0
mxd5B5/Rr7xH+77BNcSVGVJdxgcbOTv10JqDdQNcjtnnlD3wmCq7GdxwK/x33MJm
EQVD1278HNQqh3B4LyctDOimgjYGnhuVg0Qcx51OfFlJ6QasPcdeWTE9Y273gf2E
aDJvKJVySMc5p0MfIN40hA5ut4wpc9J+P5x+CrPj1ChXmFcK8ouyU6rcXbKpikyk
eaw30NaPHPxRsMFowtUcReN5hPzJSAIi+ZezuqGO0GT4E1rXoWnsGJa/OCo9AGkI
IOwuDG9Lfy78/jYgTRrnRQ2xlxL3/boX8EHMWsQUz8QV+QG7ooIyWMqoVn8i2PRn
UVZ0vLTwOSFc46glG+e156UejG6m6tWNm0lPek7J3bP0WsmXukMoN7cYqJxiYEdE
mEP4m2w+Nt4g/oauwcq5L66pRhrwONVcha/DudSv881Web1qLbgA93yimxwdXaCh
b2J3m/9oMpszle/pNjAjQlJZ22pqVvT1GdsH4TpVPnO+gCva6dvl6tx/FX43DpGa
txsBNoGmjFNkHN3NcVKR+ZqZE5JUxLY4YbwvjUxhzdOI4gw8kOBZbsGPo8Dc0dBB
jLzlPrJF+ycthmWUrgruSZ0tcQEe7acXKCPkJf9IFiYfbJxh0abIWphmgSscKJJB
dFV+seUF0uyrCDxi2qmiJ853iWjxoGrdmYcU/KCRZaU38zImxI168K3giOnle38a
fFEg5VxpxLjrgiPdZ4MXwCwvaqrcMMaMTrUOgAXkQ1CTnK+8R66PvSkYo0tmDymk
Zw0K3L4Ll/waDzan+lU6plIha5Mef22hNB5HdvC5p1SVapp7EYoFfvzRqivrYt0Y
B6AXI1Y/qByzOxfYuKyfcVpue/t895t7RZrK6Jnurf+BqdTcSfCrr7Ubg57IoC8P
t9iqJWkzbh43A5gpVr45krmxkEAz/h9hsTFkbhQACimbw3sfau4lN1EuVMKzF04w
d5CfM1Rkx0tgJVg2M5nIilixdequPKQ/pjhr0ZCi/EjoTsIrb3+THGpXHHy0fN5T
RMBU5Bi9A1Va5MhSLlxevnAAyTgMNJ8MWiezRmu81OKEWNwIeuQOixSJKgbT2hkQ
w3I24YcIuAxJaUidSudSd1l/A/lc6kEXA+ntdfPLphCleHDvKUGZ8C43eRL5Q7z/
UMWXd9zPQMkBED46DvikiFeJabgx87XHD0LifGMh1Lfn0rREnjECKMcv9jhbQ6sm
jE9GP+6UgsKM91tfH3Nxa8ZA8nsufQrKIxOvgMO6Rpij/GpRubrYkxahAYmuimkk
pG+k0/3fpt7jBIAouKEHacjJ+B+z6gCa783WxC0nKXVZaCARQ4OisRNamDiOLcgA
z2n+vcgPqGEl4VTgFmDX8a9a1ua9iqOERm6oMLb7ss1yhX2J7cIK8nm5s9kfjyE9
AOEzHiYMjlPQ5/Zbi8U7HmwYTOhldUnayA2bHh1QRQ9VW32ZNtcuIQGfoXVlxGun
x9ntNQlevcnW+v5q51IKiXfbt4U0djZ6chk6oLNzNqw0uKeihFzDW2oFY671y46N
L0HZ432gezaI/P+Trm51nsF0k8BD+3MACnk/MDwh6IvpnxRGTEgs/AQ8YGgd2ZXR
lX7dB4z5LSPUTCFh2IYuoR3z7q5SqOvH1TKhSpMBKD+UhU5kT2mQXGcIjTd8dQ/D
nYAVJzuvlKmG6mU8HEsLFAjv9Ux954pVuT9lmybpWJ6Gn/WEVTrydlwcbhMugXEm
axDExBlCojWjlwwIKnXlSjdXPVZHnZOOdLk26ApEtIKc0EzIC2Yku3uFZbPua11g
5JPbP0OlzyGP+7hgIJ1dJVGmQT/jay2lBcRoFHwXPiBEHCRecc8mJE+g4Uivw7RV
PafWynZW5mI9mI9otJcTVne8uVQYPIX1Qna0oTTu4hBGCEbJIKuIWfSbNnYDb7EJ
4CNLjVN5iCAAkNdfbeJDIpQixgyqNpkBTkz+rYNypGpO48CzSw5VphKDrF1w1spx
UEbnhRLnyEhinN4OvUJWyJfrKNqbBiAZ6A1jCF60xYc1QETCityAP2Icql/uZz/R
KZRbHoiCQPI3ViOL0ilsxr6C05u94jX+flYORKB9JkUAaCKxLOs0hBrG2vdw6LP0
3VI/GItr8uk1vpAUqCW9sZZ6T2eG9e3XEhWUYLEAAlk/bPJR940BIfkdrbAfTNTM
TkmBQs44o+CA8mOC9B1eWWHcgCF9RJLdA6chZsAy28FBZkPoUf4GVBTrs/Gkk1Bx
lXF7q9GSnZDbqEuJ2CundewBXchwIU/PCV/dcEkJNOOCCM0xWrdL4POTuz40Ml4A
O7XgntJCyVUkQCAWgKF1KUVr9IDQigDropfCiIjeNRl4wEIuVlR6QepbfssDIjWC
vx4vWzY8xhS2i2D/zsKvBfTpihx0dQ8c5fWA+10Mg950+ExuhFhz3VEgCA2/5Awg
BqJ9NsaZjrV53NqtN4laCHlW18A1c+claEp4X3URvDCEnYtGSgOo8cDp0U05wQdM
djXzAaGRvFDmUtAoA/mvTqAHJ/uCQnx98VWwvxXkN/kxuUJ7r1XWydyVhaPWp8q+
IXM46wWjXyjipfnz2E6qpfWAh2PCtQRKJwgcPXqiZijGSy7lSGPenHWFJ86l62y2
rTIBRmo2ke6aKOb5v6LeLqmxAqcfgHUweWDB0gyV3NhHzscErbRg/Jv8fz2qFaaI
EyEw7LkyDzoojBveKrf4YutRgO/3Ekb48Dxv2TtJ0Qr4lgrvV7JZBbN8HeLlDpFc
JOLRWQ+7PjvR7HzJCA/Ts3Wj0b/igUnmEEb896po3mMxdzyA8eN+EG5MpZVg6VIB
wX8hJKMTQydsZ/p7Nyrz91ecL5TNSBTl4zNUrkepWdpJzU1C6HnoTFCgMzv5W+g5
FDvRVRhT7OFGBv33S4J9zTAElyXiTN+pZBqHOhh4PwL46cje+S0eWTejLxYvaVYT
lYRfX5K9x4FU2DEVRXY2DHI/LUASS4adUL5oG4nsGI8YD0o2AW7/pD2n1u7L8z4w
8dfejBhyZdoaOjqmYvmm2gRTK48n4zC4KzX2HxruScrRcmEeHu5tAOja6kBAei51
7AGavLiOGtXWE8xNUsQx/em8DxqFV9LjsBQyTrJGEZYs0J2uiJPj2uk7r9c3/jU0
EkByr659Onbfku+A7lP5D99XvCu9DJN3i6SzT5IHQbT2LllNnHjGuZtAOU4pvap6
tCicZSFTOMVwj274ydUo4Z4G0i5+ekaIj2/ioTmYqphmCrD1Pb/PqtnBh/DmhyT+
OBhuwwhCuBGB8XJGJDNV5CrwyVHJyaeq6RODPk4VnefzkTj7n2KPU1F5TG4uMh2G
QYu7y3P7uMFplrtZ+YqqB+yzbJihiJchbCd3sVwgRMOLYs2i0rrtmVVmqqvFgoMZ
LXCx9LgIa5mdkyCAQeLVDG2TLhAebpyvan9y4inaUzbfBLg0R4QYU2lmIIUYh4sd
Mjho4uc3br+Jp6TOhzkp+SUL8r0ooRQla1Js9B8VQsE+ACzdF/uaM1QU/jhcHhAm
e8N3A5g+vz2NeKI0CYvJIcmtmQ3MIlp1/tBTczbqPNWwsF9ipA/KObcWnwoQ6v7E
NG6ocYEgPxlrRYj1XC5a3LI2h4Qcg4RIU4JqpELT3EX3i8Qz7x9xFHphxBbPow7C
Wok9hFuh6f25u1miYnKtP/izETXfbK+Yy/4+2cAm28BUsIByiHMvzpk2pU8TeaZ+
+mTxPAq7jpkex4fhDArEVzm3B+rOPbvGFpuXqN31H9CugZjz7y2CoMO3UGcO9aXR
zaIXO3+XkRmKjqh6oYM7IsiiO2c9tfH5/4mArMDk8XJl0tkDOUBN5mactB0conjX
SghqKKCVJB5nDUvkoOYIMkJ5QySEzi+85T1mIh+MhhxcIYvMqatv6YjAIlBrpkxz
MAx1gQqcAr3iIjtCE3+ps89KwRGbhpema2H77u5uo/tnXhXTwRAPDy0t07mDuM1B
rX8SGmgcOm9MEckYrvsm916AuKvjGZF2czhi2+psUaV9/KvDvTsQ3s5iavROg77o
BiIdXe5JtCALYxTijlLSIg5KdOkuAJSD9RqkNIMJ1rMMYmGtesdssAFqCsnVp800
HcYgLyevH2hn0HuH+MPg47cBAsyZFeyPnzwjE4ayGAEMUhe8AJmLtesJN8gW7pT+
nxkGkfWpt4mVBjxdwO5jGtTr/ZHs0opGxj83icAbU29U3MS2a4OyltBsxAK2YqYj
cTyae8SFhAydxY9ALm85mHb4nturW5qxN1rFk/cGAp7NRTePSNsk8VPc3kU31cpC
iBH92y0iGxxNMC5ME5YgGJ3osGBWqYyHhkC35+iRWzbTlaeBzVCXNlFN3vDOaF2h
6++5Yf4xBsWT3USYiRXhs9AfQayxvg0P38ThWfjfbPUyqLLKhdxLsh3nn15tefg9
UKJkgMotdVBsdWb2Vzd+Ir5PSw7GFf9qabVj5QjE68AhCed91AoRehffmSSGIXyB
x8EMK4r/aHEbkwjVqvSIidTELvUKYwDsLeJvziuzl+fQQtEWRjHUzgsDg1oJACB8
4bGk723NR5ANYBdVBJ6o4um2THinVCLdit5IWIY/8Abq+pgJVgBf07GM+Srr8wAw
e/qbdYfwCSPShKHMTxrs3Oie8yolN64YVc/Do3sLZgOCcgfvU6smrUR0IyeWYWeC
/TsrhpXbxtk9njoM/6D8XHGmgaFOZeL7qDePjHgvxv+cJR5syR7bImrKTjukmwnA
UzxGZWUfyQXsLJaj/x+bvdpXJD9/z9Yn1B/69I+DV3+CHVQNj7MII7jeYG03bKfg
X7YAtt6g1bBhSsdBtYzNcf0vBS/4pSe6tjMmWpssFY0zCAzygSSS1qR2LyZ8bip7
NIBYT7mxGiKNbDf5DLT8fzOqf7/c+kBM5Vhhu9IBk60myjqqLtm1monNzNdXbI52
K9lhNR1lmhNDx3zoNrHCFMhAWIWXlazvvYRcZM00LVqdYOReaPtVdlBb0pwh2i9J
1KpHL85dciEs0fKkwAJ24hMgplZGjzrZP5T3IhLbSrhy4Nlw4guz7IR7by4WKMga
Xz1lD/LUeKew4u59x+0kCgAZn9oDlD5/V8McjnORV5d83NN8wFv3/MNs/fyWzN3A
sG3wk8Y6HKA3/5mIReWjRBkcLEsd3EccPkVgzZCGVNSBiRRe5RGDi/pl+aEDy1EU
DCANJ11NGaNv+Iu08Pi6ZjW2xVw2u9bE1keEqwSo8vJye51Ey2OiUVVqVUc355P7
0L2a2fQb2TDqr59LBA4ahai9mRELfvVhJ8eEftHchzYyvZZeB8ZtVy+YgMvqCCpd
GKVunVVsC+gk/YjkrJbukWWlshYqCrJ2VX0OhWMtm90ZJzJihVhQJ+HYiMHU/Xub
ploi6QKgT+gi1IgzloGp+s/6iczCt90JIIZDfKrBh7UrWt6o7ctoHMJb00PJpnuX
KgKoBst2WTxRNtgStbPcWPhRaBbB0RkoFMa7mqAe74+3nM2w7nqmHJ4EljD80RKJ
thOQa3/3WM7JMS3HN6nnCLSVZtvcIzkRu/bcVfrhA/TnrWvLOE4uivbYzsJ6lHGW
YmVVaN7MykRYlRN9TqqVI/EkSTe3KeK2RG3C6wmOpfpLUeYchRUL/+Zdm14OOJdB
X3OwgDDjYVECscbTFhL5W0w/p93q6EA7Qdg0kL1pkx5IiJDdNccpO5wl+LEDOC2G
1bb0ZNTLD0zODPEZfqwVPU3JlK+kxh81q1+p7ovUbYpoi2votlhkY0fv13d2XpEi
VWCTbmbpR5mtdZkisZB+1TFl+hezde5jv04rtcgHxzHacawFlX9zR/phM5uC3h5H
Qa3qg6F2zlzGeQvB1GOfgEBr7RBD48bGLrFJqkmAvz5y/S5y44uecxw79k27jWCS
873VFmeq/BjX8y758zvZyQ1JCPiNno8oPjFbeSLUOF5cPA6OBnBslIKPqxHVnh14
pbjci8QhgawDcpHoqbqAJrVp0xTH8uxmY2DbK92z7RIQz05XtfKJX7PeMxCwpMQy
JvRX/+kBQT2xrx1l6ueQjHJTp189gHUuZaEABbHDauIPfU8caIGAmOIJGco8KFec
1ct9vAlYT+jBRxDg6OEQCmoto+4mr0+O3dX/Q8/i8jaC8Zv1+EJ1d66MgpNzvGj+
rxqo/T/Dns2kL9gJP9vcxBCTkU5JwXwl7/3XnkGzXvNlLwQvc0Zofpz20Is5uiVc
rWekq1BEW++1xSe++feE5UDSCI/d9Au6t5p+6t/wciLakjKSR0oFTa0XWhymRKnh
lSBOdIph2VJINFpPxyhFKiwG+s09P1qpTbZRXUJ2kedIoA5sJ48Iho6tMWKwaDPq
8yDZotC+LDFaA3mdFRMHrIu9hp2ddwY/EP9BfDFQJlEf8G7S25EKeZlOBsuRIxEp
Tc8dMdulwk/H1s2HauPteaiQxiu6su1Ob2jdtw1v8mcyDdoA66rtjNqtmQpqHm9d
TNRccxb4KUqypk/p2SalGXKYGN+0j47jddReF8jbiQMXOMNgYNZvNn2K8cL0Mqdg
qedgM5zDQnhvkWo+g3q0w2XNmhC98JgRma5n/6DLkTSzLF9aExK5xfRSMgeob5zS
Un+NheJ7de9QzLPw5g358d+JZBm15LdVgSL2qLO5O8z9pkhYp/dFaYgEs10DWNLs
q95ujwntjRAlmQxYew/HHUpGeMvtKXc3j0ET6mVRvXZSPxzQSm68LFuNZ4zCf4Q1
orZ9SL1e6ZILiHT77d1neRaFNfCaDBKv7bYzhSKw0BDdYNEWN6HmDQPYmjST5hjq
RIMSVO8FGlnryZMSR65jTKymtFR7TkP4lX5rHsRhZnkPXky0UXqqHdRLd9OxwKu8
F9Fvx+2uP8lOBgZL/ztLzxhgfKtELxkUvcfjLGbsAV3rQWPTW0CwZKlv+dEO078Y
eH4H1aUdBh+yDRxXbNenZXm7SvRjmm3UUUkCq5wiXcnhohfNAH8uz3Snu+6vAkwb
G4RSf2S6Anzd6Di3ikH6m/krkF3JAslLsXI3GjKocL7m0SIwgBPlG6qFYU6P7YOs
M0mLqXrYbEpjk/Vl0pXdvmRPjwcH371d7ytvqA57cFViAmqr10DapbFXxcfHFa2E
+nlStGAHN6Qx7zFxmtlXhRASAoG9/MiVbgJwSYExtyb5VnUEnioJQGE0ZahCp7Mv
sa/FoT/M76ayLR+000mbYAaWbbeRP7cpVlBioNY+WhAja59AuqB+NvChemhiC4HH
stSZmI8FCLeq82hfNxYk/bhCUT8A4L1jZ+H6HqMV6DNyrWfYzm3w8Qj1pONFeQzx
xVY+em4o//RVWll8PXhSSP6rqwmHeN5QO/WJCgtfLhDgb6BewEjjyzvx7SqKFa3n
zCzb6JHbE2UAqUNNah6ZySaXcIjH1IqFrnR92kb7mIQE5/rKV5EjObRWK59tjMLh
wjxpl8Wlkq+Ob/VhEDk8BTtsCz1MyDmSpjt2fuPzASLStUe5PR8n0IL7sQPd6otC
QMsPGCCSUy4H7ZpX8hzz5i8/JsA0ZDNeQ3BtCAyZ2XSVd5mrh9ny0VnfpSk0Q2b8
j6lJ46cVJjqDs6BmNsNpnXnB85ybh+lmYGy+SuD0laqgy7a2E4wk8cUuVNXWVbhG
x1B7RWnAm9WPAyFUCDSrvoQ7fDTW0E+sogTnkMjXZOv6RAL2hY6t+kkyREY0Yrqf
cs3UINUrP9T/FrgM23vuzhCWifDg62XuGLs7/J1SeOgz5yPOqS7KoQyEYmVQERE8
YTgejrhu/XddDcozJvD/+FwqxDQGXS0l1C9bMS2oBpT377rtDmMsCQqG/fqadCXY
GXrTLNt1IiIjsD3YbIJp340hA989sul//UfdEggvKTKKoLygm1eT1fG8TMyyoRAT
x0FZvmeg9X+gxqU4hFLK9OLc0A/ltxBYwmJ4LE1/L7nz2NFvbkPulSRAiYnR0r89
uAjsJJHN0FzhXPC1O3S8kHiT4hEFNLOrSeRfbKaL5mn7Uh5p7PqtFm0/+2p79PVx
/lAogWeELh3v3w0TR6B40sgMekmOaef01cbY5J3y8HSHR8mZm4PRrl0IsIR2+wZD
Jjb3RYMfaLKEOaCjrk+T/lKqTE8l1JP/C8YOMrfaNnbfmkhUmGYMMuBPi0hlIAdg
e1BEzTJNdTFAR3Ib+ypJHfIMHRMI0qS8Y6wFH9BMU6i1Qivy8LPur+xsh38OSu01
WkMucAKMwA7IJfMUgqR4JIFB+0+G0yDse4q9YyiVAOk/FRcts9bUZ3eGjCUn6l/8
YsDmBUdla+Hus5Ld4ROLPs0jK7JhRkx+QOjKOXM+r4enlb0TJL40AmKPYx3ZhvbD
icceiz8Q4yveuEhkTIUgTy7y29Lkg5Cz+i9bvmYJCERo77DZ/OAk2EK98E2tTm9g
cKGYe1tOQav9OIoP0eDZ4LaOuNPn9vCDpUTBIA/xsp81jwSKvEE8hL3hicAF6+DY
lSyqjkKBnyRdF/UQ45CE2IYxQLiPlgdVqOLKFGN8siNZpAx3xelPLFStpttwyb75
j5i5hZUXmPYgZOgLnffNzHgZbzXWPAHyDdGK0VHtekZcfDVYWDBpJdkgSbEaNQbh
NpJv/LXF5vyUsrIQwNk+uDqYUElVUmFVBE6OILD6cd+gke6MpvOar/PZtskvxrql
ylZ5H5m7STNkjvf+DdMrCITl2W1+tWDuTKxPb08HeQKrRYjcpPL8h2azC9wEI5L7
8dMc4L1cnGnSU6LEVG3vwi4dM79ALsw8PRQzk7o7G/+LWnSu96XBOuIAvhrz9DuY
i0v7iPJZXS9SMsvtuN3NFnJCWChM8RG9eYo+mOxrWZjXI7ef+5XkIi7arCkntjbR
tXeQnTwYhtjuSY0AvFge29hCBhI696QOZtYeQjQpoBcScydXa0Ic8JJNofsEdcI6
bIafdwaGiPYMBeGVuuhvXB8WsnPoOZJkixJxLD/lZgrqiTR9bUA1jAQMdcOA7qug
V9poLbEmsQuJlY3gUeqh2XQPUBqgsZqPDMxek0iILqE2iUsDeOTq+SPiJF2m8ah0
57wcZ75h46uCvOJG6QYnklso6/rXJY8AdAjz4datWBtduFsg7BpjlwjjTa2xRm4k
1Zd+yn1cuBwMbdO7MxbrcsWS4knTWCjJVg6F9jPcDNtt/s3FlSVzBnLIU8xvYgL4
QbPawRECMe3cLGQ7JGRUB2PufP2f4/nVwEshdmgGzaRifT3youmiUq/PspZ7KX0L
Imqb62sHm+0Jz8gpla/Ovnzk6Q806BzeEGJYF66k8rZYLaXoI2lgYvxn84XyFS1W
uynq90+L2+h1vsDRdk83ZUJ8SDFJ7F0Vz6Z7XEZMaugS5LTNWgFaXZidRwEMvwUY
DXsVN834RFjNgQaHjiBYrX00Pksr8etZIDniAltQpPB/TTpveIPlwc26OhSL7X10
iboHFoJsxzQjhjnctbQD+Ajeubrj6MtNlBcRkspFg1HLQbbYGg3fgZLEtmVS4k7X
yDYxnDj3KmN3zKeSATiB1mrdTqsC1ws8qP4xfp0J9IO2+lxqicYlgVdNtPV4aA89
BGlkdZKBo4BRmq8eo3w3bOFRf7hmefxqZKEQ+9hG5HYY6D3S0aAS4OeYAX2GNaC8
q5ARPu/sMp6quoSQmnygKT//PAL226/LGNiEfD6HO9UpiYfDtteom8ajLsr1SLJc
9xgBLoE/NEUNpXifgOTCfWHiCiooqXwyJ9XRFaKpKXXyGbR5BhLz1+OjtEtjMnkt
byCKyTJ+xF24rgfczZA00G7pcR3F/O65ZlzLcxkIaWzrzi/HmRg0KdpXNnPHDcU9
+dxxCTQpN4Hm1mYssdW+9AQSUdtCwabUSNE+6CVsTj4gbcHsuTZgkc3QM3EYyZyv
ckux5U5L37iSs0EW6TNcm5YAm8V6uoitz7gbzKCw2AT5dVzabkK6PZm1cW9taLa8
4oX4Km4vhqJ45m3W2iw6EeozoG/E8DMLiW/uZuLd2sbLTjjhI+ONsAHuQpoRv2tx
1J+cQqFm+DVjKPDD7N33NuSVZFzKxm0oIv3czsDpo91SsqRggqAnTnQK5TuYWg+O
ROuQn9v9DtvWOYlXF4lPEGlkvTIkijL1HdpnmSgl1j6ydn0klg1WFi3X7tcAeNjr
noeviOcJzLvoQh02ZavlQx+i9/Yjv9H3QhtVHs1vUlz2DTV0o8ITXnhqmCKZFLqO
yiPraMMP7PFwiapAcdnhV/bkiAcvrnUdcejwwrx4ZG/jJigTumJuN3sueX0YHnA7
9vxAPM1alc3sSJJEEVV5er/+TCIfNptgdgIjvoIpNhryMtjCpaI57lCAShialclO
rRp9hxwKM4VUM1OJmuTqVh4dURqlUTjY1g+KIf7lKWhbWxJCP21/mCMwQ1JlpoqZ
x/WEYH+1f+hCNsWCulcj/GttyNKMJiUMwFdv2zBIUJM4vjtfT2fAGULf2L4oVxQP
q4SJ1qTN5RwHINUkrB6yAp38Epa2Nv/BzKraJ+3yhKUIeuSQ8QcUbNSd9fAdn36l
lisJBkoWy+k4hBNW61QjeaP6HU6EVr2Go7X3VL1+wmX9CgoaGQRRQ9p3T4x9r8RA
HbW6NveziTOOEMOwDGRv5bQe418+65QEm2pW0/pu3mfTbDiE7giX/uorV7W3PDlY
5/yuiMyQpQk8Jm4HOGS5EyOwCmaFTsCLS5+3IXUa18KzImXH1gqpBwoaqnh8m92U
e+yjEz9fIml4m6DpOgIjzeRvUP/34dMqOsAc0ZaOywUp+SyQzyXLWEn8gsGeJ5Lv
p9UTyZOpLhfyJtnwzkqcUnnsg4Dcftp+dAn3kDJ+9fBfZLrRDSeLpEYWbwwjNDLx
+w6Sm1GRzowiRYAOrzxfV8c4mOaVGO8I6ii18hZVR96/JsiqUMP7A61AnUH1cp9I
vTOFDwXraNXUlD/GiZ0GfziN4HX7Ucevgtp3kQkF7osY1Fkoos5J5wq4nKFOawcZ
RPnTH5jWsWFeAqnDrkr4xVOC21icZFfgPqq/oDDyZPp6qOIXNHl31c9mu3P1i85C
vrrFUTXY5Z4Je747/ze5PE4L3lKEjZnrNjyLzWaUihNKsu8nftQqoQI2kCHN9I+x
SRdp3tL6vslc82Q2LsRp1FXFnyfuTdor7Cz6K1r/SD4DY5wid5n7S3xM2EoC39gq
VQIwXP6s3arfA2KJwfXXinB1fb72vTYjzMt2WZ4vfpvTFXVdrHcnBbhjYEAddFG9
NPBFrVYfT/8EHnTPTE86mbEUnyb7/jovxhhoGePzZWuxD9Ly4v8B3VUpATAZHlE7
buYD92xZoeb2W9geA3zxNZPVuxNjxm5mDmh7UJRUWob4biApenxojKQZNjs2Ki+2
1q2lolZv/mBdqU1gF0pJ5hlIoy18jisC4atnnlyNmSJqe8NlbLY491nW3wYMmRUa
SYEBZchUg0Krf114MFoNR8S4DnIP13k+6S0x6BTDdSKTExwSfmQ19RnaTysrfNFz
46PeApdwSR5isYRwhA43CyExpXYX8xfKBzO6nB2OJrZ6fQJAPe0rrX8iy5vE+cGR
E3du8IZS8aZPGQyPUHecOFa8vy2NbDhaBONqaccFPNtlQUIAAg1JjyuQomdG8FNg
3CVUqufVpnXf8V1TPYLgb1Qf1rrq/5ZM/UPwDCR2gZVWJ3KEkM+eW7aq06dLdMFP
XI8f7/PA8pfUeeD00SR2YXUrNC9JaeTXJZdMh+yTQsJPO4WQ+aACtuLZcAJwBA8n
t1c0YmMYdVYVkOI00fLfZX7CyGRJvReDzYFG/I1q8MODuQHII3UtoyChl/nW8Cw4
1l4mLtpjDup/B474vZRNhbIn5Ytd7yx3g66kcYs37DX4JBPmI4FviDFaSfzwtdrY
vv9eZpFDB/QOvREl1wENmcon8xb1I1e4NPHkR9urp0QzyBmd9JaqZxuc5TvlhN7t
pCXJtL+E9VxcsUVenRGxzaI1b6ClLeLVjT5sNpn/1MjyMiHooW5koa/Lc4Kigotu
BC4uscKO8EqUgmNr9oMjht1onPtwIRvDZ2j78/Moht8Ag52yf5bkKiExok9Xs6VC
eZI6DXIEInWG0qj+FDZG5WuK9dw4I1NFLLLv7lhZ78CEnTKTvzbC1fLWE35Uw1fp
q+h5Kdn+WVC6UWo3YFcB4+IkhBtW5zblok0TzTu61Lt4Py0KD5U5OPxEB6CJS9gA
3CRZnPj+z/aPAh6DO4/Y9yryVx7Ths/lYa4MurKbLqPfaCeFdj9SMpvkrjT0zsbf
P6dTBtAtnBwTh/1T3SZp3b6BGQ7RlWitbA27Atb7rC4nAfdm8oabJRcm0E2By2ZB
JTl3fhwNIXieRbUc2L1tugcMEY00Vk90Ih3W1Sr+/fhBm9ETJS1bke9rhhatrFcx
Y6f/S8LmlFkisZdjazCCOqth9PuHlOIPVZKgCYZ0jDZgpI7qNCzRbyXpZb32GrAZ
Voqljh2r9ijVWTZde03WLmZfTsqT42VJeYnvZRmckktpkd4bPSEAsr/zV7R3ZFDh
3My86nKa1eICb2WI/ndkxGw3Pe6WmKdG1ofQWRRRbTJx95KuDZaWO7TqzawA3fjb
+VrrFJd4AZ0hBSqnoCflTuxqQD/8zH8mVn6qQVuT3+88w1eY7gixnvQ3mVMCFz+E
dkEQcqVEszuAOY5YSZjj64NV9mzI+GcvLAciMeS/fzPAB5qevc0l1g7tYLWL7mAe
UE89qHsQmZlMM1cLCQoqX406WeL18huA3W9aKit+Xsfn0Yboz0Su9179C6lkaDXE
IOHabt7J8/2Lug87onkl8m97fZr/Urx1yYIBcXYaFXsUiOhvGT+0q0ArFG95tT29
Ctbj/kzxT2lMDAHLI9Y+gh+ElINMOlS5XwINjKiXYTR3OUCVjRkY+parRgUf9CBK
7Zzj0ecCe/Fu4XF4/BJ9wtF1dtjP5p1J6Gbf7DmMZpz//qRl8w9A7drD4PM1AHC/
04JdjmLKaS5Q6OSj7irY5LWk5fkgvEExH8r9RskLueI9sxbGrIBZw0UI1ThpFhUR
IniPSDycUDZMmK8YljQ6m9nHMElRo3EKgk373K6qN6GkIetR4fU9mupJ7qnFTlge
HZAJFBorCpH9VLPg0SQckagddGDQzfbgDAJZ6EcvHwDGLoJ4WB2UcLDY1yapfGC3
vBNePaCPc7LStT7HF/KSJ838P7dn+Z4Y+f26Vcup2rSk/BfZPKWG85+SF9aUGBCm
B3OmBiYT6oZ3RhgxXQAKSD9LyQPibTJi0UK0c3gWrbzn+ZodeJkEDNWZ/9LugHU8
D8ZlZCdW6s2Lmm0pPZupHkElXmcYK4TBzF1y99wvHbVTq2a9963Q40LxuVJeIJMU
K6ypaFdsyWanXNZfmkpzxnLmIhCbSdUAdkS/0R7ym9TOXfPP78FxNE0T8NWjbxvh
DnzpgFTSFXZXPOMxNo1g5ufHB1jQCcmodKm8NgubaTknoVA1zNcC5FKfOPE1bHvE
4ottQUsjDQdXW+yuxdailyrW8/S2HHtUXUvOz49RflY7SC83TLlmPqIJ4oVNkgpr
qY7eq0KohqhVHV69zPkI1pRHoy6hzBdrj8jfgeHx8D/CtAYk4aelZ9WQ2Jkteesr
2Q8DUBBgbjmqmfe+jWc9cmjt639MeJGpoNoqbj7KlcG+m7lV66FkdJfWsyypZab8
PwCvCZzcjHgqMRG0kuqfRWIo4WHcRD9K/hu7ZkXl4qovm8K+7OSEAHXjo7vTmFNA
xRs3V8TjhB3eCQu/cd7/ZTleRlofRCpsO3mUSIV2WlQOCVlQsnU3D4o8jzW/zjoV
JK1kLoxh4DjeOS2WW1eSrKP5h0WBnIU1AwPFLAPte2PB3OenPUBhCJSjGuW2cjIe
0LQqQ/aG88E9lUX1dG+nvhBdvk69Zsj7HVi0ElzRkhSAafesvMrLQGGqmXmOm8wK
pMbVv27hMs2Dr+QpTHSFd8Ufo8UiMH7Kis/EWq30Nuw6Pq+h69WfIP6e+/FpV0Yw
p6ZYoIJkUu50xv2w0YWaNtzMiOurpujaAMZHOOCTVoCyh2zKSQ2T2YH57vLJ3Q0f
2SFKBj6u6aGF1pQnG1nYPcnAy+oIHUMw6tL9WSJugnGatkqvBMG/zeqBRPaVfZTQ
HLfFyTXHMSjfM2lJCPdLXL6pnY/dYXyHS1T2iRvh0HhvntmkPG5E9oJMQm80ZLgv
rNhGKAauWZHrhoNe50UCKe3hq+CtTxzOpLsQzH2i+BHwattgiBSkzrPnl3HB7coN
DaCZEKscEajF9MeoNTxGyStozAIUWiEMdYgzbXYKSl9/+lilcT/eEj42aJZk2zST
aI0HmsnhIeZnCi17cFMYOQ3eF+AUilnEjUfWSd/nYPYNGzqcl0rAmS4IXn/4kfWM
oDcpUV/0LO+HdhO2gf74WRTogqhspQNxuynPh88VLiOLFl0H30Ym6uPZ72UvBZTB
A72TFAXZH7nXgDYgPDstxmydwz6YySfjSifSVDjxnIAcK21nLxPtW+6Iv6TiHEpH
7ByNqzbdp3Y3p1FlE+d3RAGCsSDPbWLSxXjGshPd6L32KaA+zYzWpKf2O9G7hYYe
1RWK5qKD1WXZ+91oM/Y3DI2T/AOZJgDINIhcA6STDuaHsfHJjSQZ1/JnP2XGiw5K
lk0KhdVNb8gGr6my5p1YKIw1RyIAobpfj9JZrxUFKeqQ9R2i5CfCKPaqLZEL9prs
dUQ0kcIlc3mrD90LU0W8SHPPzniU5tN5w0OwoA+8w44cKDddrqSMiE/ZYwjdpzRK
VmSU2bK9VJ6l7CmqWoJZWg3IKcMyCAJXz5edw39gg7qh8t4Kfq3prnmk8DbYeJvh
1qZKK7DW+NTZuLTgo7R2q40TaX6yOzXji2b39kP715IEbhv8mLfFOpXNR8hQbVDF
A+BI02rn1Msum9MON9yrfQ/6pK8fWXnmWWMwNvMd4Ha3aOtULFDwsOxOu7IdRqP/
FM/2yiq6LwDFG71LrFK7nM8bWavk6S9JthJQNMtex+IXZtxyWcVSlT7ov6Yc8WeA
dMiUL3oqhpJ6O7ZwJ8FszLP8RU4ZtsbzheSxGe419Qxpe+6bezrCiY28cqFSbdtr
acPUFiExwvglepYoJ2w24SNewxThbVrY854tvx1A6x1eKikCiUtLAN82WErmn8CD
O3tSA2ZHmiUSYS7gg5VB7o2Wxw/wLo1Bq/F8Qm0XHKFIbPvoTGl7dOa4UAwYYlmT
AW24JHM+N0CUHFX7UvY/U7iI7Olys0TxfeqLcyZVi6K7SRJ2aOx7aVXOHXO04HtW
NntlK6tjYRH0lX6CojxKaNxJG/rtRkjdYsm0TML4LE/g/n8cK9nzgGy1XMq9EWcO
Gx5mx24vBwH2dFRAsBmF2nyL7NkF5nNBOw7q9cxUHHbwfrMavzos5C6YgZ0EwXco
FWSGdJ9i8koGjcs7+s0GinxP/uy4w/dQIJ9TIEgksJK6H4lCOhgjDRxlp0tC/3aP
J+SyklL2di0aSsb+1ouus8VP+vEdgZfIhsqWZVcuEmFqbK8LFrPHXoPSi1/kGh6L
y6DFyb/5fGB2NV4J2Z4sVIjtnqAoVnD10n5FyLIqO5GuqxTdQTEpHZTxC0TSNr3g
nlIOh6fa6LAbo6mcw+Zlk1nxRWuVX0Zat6HPCNu7GVrUFzn1syivZl2xTv/sYL3y
PC0wGLPd98VKalNr4VcJvLzhHHH0aOun3a59tvWLlHwt9Rl4+MzjiFUEMpigjffk
Nm2YSLLU+d0uhjGPWHUteC6tHRIxdT2aN+Jxq9+xm4KmRqP5CBOVRse2TAVOPJmd
ozW5tVsBO+KzB5spqPRXEtHzzN8HCv016DKmGZpeNtd8vaip43fLDZsH7AKQeKBR
04pYuVbcCeYkKr59C9zO3eFk+7wRwzxKUsYTRyJNCVuVZ/QLkTSoWYLVTJMi2iny
/dkN6C+cWcjIt66qlLO8+xybKtRGcSOvCyvOqoqZ4DNidv0Adwdbgs6jhxPmRx8w
KdZOfWBZqwmT4tr5spm4u0o6n9VJoKSTUbenDHPidBKP8S9HIRMc34dbJ+sXpuA6
WjwG7odjkK1wFRz/QyFQGyVtJCjOqdGy4F8DRJW6N8wrHDBZP/2E/pcTeSf0D2bO
tawRr3F58+nwMfyldYyAL6y1eQOkr/M2EKu82QO1Odtjw9Pb9vVUYZ9PBCAYDyhN
kdHe4J/69/VefN1bPiN2dWwCv+Ic6GCnFgwY+Au3bnGRnt7GNs3UkiRQDDvvH7NY
zHopu634x8i7DAPzsso9FeUiD36fRrZNGSXYzPQKtLb4fnrtbV4gMLkASYnE7DoS
YQPFdtcJW7LtZn86WdOmLz+G90zGKRSFv2h3860us5xu5kDimkKN/HT1W9Nz+2XM
gi5EG2UYa/CrEoEVBtVuTloZvc0VqD5VWNVYdNHVfHCLGNV6lOOh88SZQqRW5s6Z
YDW3DLYGZjqIXUvwJeBujJuDbCqVeg3vSo/hFYwY1We3M3TTn69LmJ1rx/wGaCoW
c5Cg0RPsQeBPn4Y4n9ooEsNsyPF0Zmap7Yea5TRLgPdyCR3gNzXCydQbzrVZtyzb
JCnD00jc5niZTconTCboZfLvaKigzurE/FKVzi6v8WhSpJqLPpgNeuTC7o2pNoez
/neVn+I5Wsjhoi98/fA9wRto2cNygDAvchEl1FJCTerriytMqbW3PML0NN4mcazd
gWQkZslyDVXKdAmk0KGcLcOv1WFqimjbJXpAX20H1lkzBJIDGzO7BHLa0A3LYQtx
7XY6dD/y5lU5pCEDCuKMSpEV7afqEM6PrzSkBCz/E76+3Dr/11RXbhxtZTJ5ZhRP
n8VathJ6MuhU0s69DF3aAGRIxMs9JS6VUxRpdm0pilkxkUfyb0Z+lHCg5KmTdPIl
msP9q2q1x1A6v0oKHjy3v0UTzvm5drsUwZgKMCVIuyql9l2N797iqeHwVMJRcva6
gOZL3KOsDHC5iP+WnpbaB1bjt+vYJ6VpDiJqpOo+LrFskDqknI5CadKyvl2f1kr3
9x4BnzNEpz124MZRsgU/IdVK3cbJ+lfHCMwKCGx4lJfzT1pBqbesd1BFnuplGyWE
AS/Y2YSNRiL6ft7Yjw1/WJ1g494SPsw2Ofm2aRJIEMg2a0+pNrMnOeZAJQcCHqY4
Wiz9/rgDcT6Jm1ITpA0JA6zQEhF9Z3glLahV+vvh7+6eMfa6g9GR6SM2YzaPddWq
HiP8Y8M4mTcwhPGmvXgn0alk/fH3szZ5/Qk08pqut4VPG2yeOIaAW8YUbZU/4dGR
fulT+Ghv8V7jCOecRWFj47wD4S+nfKwzNezeLoIvcXtwqe7QTXn3XRmMlB//RspA
VRWY001ViOn7zDrIEpFeUjGMrSxsdW45D9ZxF8tDKlNy6+v9ITfwzBU+5XWjhbMl
Ld5HtPNPphM1DRFWtr8X95Yo+MxEipfP3sRi2f3g/GxP4DisVvV+1Wa2gcnVc3Ov
J0O0fsla8GQsdM3ZXbHvseCbAmkAhsdXLz/z6b5+Luioi5uc+ExYwueuxGiB+VEO
hwoU2QiKZTs2eD3TF281MxfJzUCiIObf2MVXullWmpvq9NVELAzoWQyxqp3RqXv2
EVYMwrA5BDNJNLq+U+iAev2W8S6Tu592IIWuXvia6KfeqfMWKuaZDdknwyAYz5oF
q+0a0I9oHq+I6xfiy1Msb9DXXIUxQMcA7cWKL0016zFIY5FGC56JDCw+Z3i/mv5O
bCSdSHusojUosld7WFIVWiW2q26EdEyG72OhWCFRTORvaf1PQqIdYDr6nFlMRcd2
iRfOMfzKLwrW6xjkh26GKBRo77lqXybiAOVWXaf0tCFunyLHmG7rcTYH9wG6BnTf
i3nDl+YqAwmGHByaUan/0HboGz9Ed79bb1cHtU5NW+WW8rbaqn/aEb9IaRDr3YvC
xYUT2/AWqDtC5AtMnuQQYF3EaeNX0uHuT4TzcgDCmmKweQzCVfqcMAeDx37FIO2M
uA8uGdEQrbAr80J9E1XF0WsJWDZ9vEv7HsbfK6RUF/vwwdVk2MpoFiCIScioxgJT
kzjKrYDLWvfCSK8gomi2Tph85cjPZjA+qiswfBm11JpWjLZiPwiRhtsBLsk1d4Og
hkXMkKuClc6BVSG3k3DMQnFuMvqy5LDng7wpfgB2RQH+YfbPOvSplODTNBYWWAgE
5rxnDrTo6yNiCjTtLbqEq0UUcQAXLyqzsGHRqCwI6sf/73Adp8L984yiDCifiu5N
aRebdzz73mKhGNLQXNSI2ukyamREaLR+HIzHB7J18dj1/sUyNiNiKD1SQ95xyvhA
uJw1dJKqK3Uem8HBhyNsP5JYbvFcZpLFWPH52sTwmmDmKgBWSvaa/H5OaIGL20pC
Y4FuO9UFvXgNqOkPXsZT+FAXNEpWexu780+4v2KVkMfZYWQYVCw9O2PXzux7aqNj
YmbaQxh3n0pkCI5n5x5r9Hc2Ty38bjC6WN+9r9r5Ddeo0d/4Vl99DzX5MLxfR3P6
VaSf7or0kv95U9HqI4fZGuy/V9TQAjBfS8/J+Q0OI/yA83ZPyHYCQZ0clepT7nEU
nkBN6nbvPCgdL/qVUHx1QIj+9vWuPeWfBm9OENBRabdb32zr+fGTKEN/uOle/D9O
Hb0IRXax3ugxqIRv+OH4OVM/SMSe6jKp/LUxGoCahliGDivB2fqVkn9O9tgOwCeP
yV1iC8NkHtpqZCU15TKj/e0giOb5dX0ogsTay+vC70dBWf+NCnDiCySbuRk+l84T
8FG4OWdxe88tgNrlweLEubVgd5k5vImc+fDnAY6fc8kdOD242wvLjxFSaITtAge5
d2TS9PiZh1y0Zmy4UtyF53ncML/wKcL/X4SODHOUxLtLj5IVDoydnHEruvL9i+TP
jN206QjyRfbG1JYUJxtD+c7V4r1/zohHKeLZnHtCFE9tKjsCyDP6Wlh8MVYO8giX
F1IsNkuiSUTRqCHshh+83SBLnpGI4IqW+8f6Mld1r/l+4e1SMs3OTG4z6OBzRMgr
D5q9/DI7Dxz0ZtyVS6M6cAb8f32d0ua7DfseEQW+JfpA5ydkfV9BukUM/fEC/5q9
tq7UDuaruX9AVqBk+aRJGBwVe/RorXf67rZv7XMzClPj1XpT4z0am1tL4BY0Hg9P
tPjQPhkGEEXjMkcL/bDnofsbtO2UkmQJuj9542DLwa9RFYAv+KU0POSiwGhjJY5s
C15jKvM4NSW9tnevJoujv2eHyy4j/LCv0HUSZVg7eXtbLp8Twuptl9yNofZiKJT1
Jts2k1nwRSC5KqADcYJSVZwJCeogvsbZQFiJ39AfDSHKk+mPH/xv9oqe0Fiqga2c
xwGNJszFN1zXxw9lhj1sXkjaLVoJwON8TEquKHh9aRWgkEdVumlAVszPR4r0R5NC
VpBtvLR3+Ez9jstjB8JYoMKPO086RebJwp9Ji6K7xRZYRbtzw5IjjtJczh0oucq6
mMq+R5M1BCjH1sFFmNfCQMaxlGQ3vQ7qXzuN9sSiTzKQr//OIKZ3S3jhtnYYDrnW
bwDliPp+chayYcyiVMWd1WXItUYYiDebJWejt6EXO1okRPupDaRfe/HSON7jlH9w
bGWs+1QdJvR2eGqZxm9L+omYeoFknNrGz7X1q0ybhGkNJKX8Tp7w9vouyVPWcKoZ
wCXxOnDWB2+EjRlIcH4VxjrxWceqGlNZxM8XOKNiUanUNkZVBnjuL/MwGdIwkibd
otv5KVkeA+9GB+KhLUyCdA97O5Z290havnfjMi5OZO5tYJvoTlkd/MwdYBMzF7Gs
hgj7gCtSBYiq9uV2kfKipQWn1it93YjoRuBVMxCPy36mvOqaelBgJRrDzv6moXHc
4ggHjfkxFp1Y4JRuA/N+FPrOxHFakku0ylvT4ULMR6vs6iEI60C1RXe/Lowr7CzA
HUeWSySFl6TiGf+ebIpk1WVD0I2Ly7AcY5XZoXSJA+lhRatFs+znxHFRSVTgvihU
4ARJaq13B9IQGWl33x/aJY81fnuNWIwPbK462IDmHP6ZhbPDbWliFVe6NpYAXphi
NXMtRLeZ33N5h6y8gWCICy/+FQ8eC9QjjSyEAy+W2/edm/id5yob0WnTdNDf8+qd
fvckUL/a/0+1I9y16cRBSvy+bItTwIZlALxqTAFEC2MstGbSYP0+klFzxexVOUwy
jJOYbIi5+mnwm6iajBTstsIBIpFjxnVf+zaOfm5w4AhE3fqptr4jJ+aolNT/Ph+W
OXX6yByD8l5PJR38c7GNE4ZZFpdJztgE4HO8nDG1dJ0dfRShZ50gfMbgBU7wtDMJ
zShbPp7deSEwe4TcUryga1mhqnksatmxi6W6pY9ZmfG7tMsTrQsvRWYVFAI1+7ma
vyz19SnRsLBMfrb0ZEFa/RDdkdJPN5lfcdlc36AqJ9f9XpmS8z3Ndy3xV37zwcfL
wD0Oad7gzUEtFM+660g6/j6lTVGDIf806cKJ3FwgGoPb4ffa/n+3g3g8+qgYqn39
iCqi2NTGIIlrTEvlHJXuFc2GPq6EPYoCKLBRFqOvYprisD9Mdz/E679EEnYJ3Nbz
argV9IBWXDUkomTwsnH7GRhRxeRdJzHjVY7sVbTGyXE9x0j6lXW8tIz9nV8U6W8M
rFH8WssbJHONIyC29OEVDBMf4OGdRl3pvZb7c7RYkdoDfOqPf5tui4odGE8Xj3Iu
sofau9nZ9LJ6JnXzvo8D8P7fMW38cNeK4r1L4oN30l2ulAjxYfi2aib24iICnaIc
bMN/SvJ0m6PFmuNDZuNue3s2VJipRgnZfJw5thgc1rUy4gPpQ8TwiubLqSfuuo1O
63PJFvLEfewbCGAFkM1XcANjjWXXmELhDmQsxMeb3KYSA4GObz5W7BnRbMqCVLYl
N+OtUAm+2n/pxCYvOnZbJ1vpjg0pJfJhxpuoEWswXbHQIir1/1/rR/Uxd6kRrnQg
UW9VFUPqmH/p8j8HDuFl6kOn77xyvHgBdlvrTG/exFEJNOj0QI69HY2UuyU212W1
1DbzXjFcZYQ1PRTq2znIHwj+0Ho5aZ+8l/nNvnCTJpHoPUzqnTCeUyV3q2wG1rMD
ftevj7kjKf93vPpezz3s3BXgcqj5k0FWjmx5hr2J8fEAYWgWIpEW5r6rCDI1cDj2
eeCaoTQjKoPIlWqHJ5rDbkXScbDEq0x/jpPxiU8873qu8l4VkoBY/Ash+/X0J5yg
blpLEJuqfOsQoJW2xitxfMw72HVe2qhG3b7MDj8oxzSb8tUBcpSlt115jV+a4b4m
94RGOHxRvj7wvnNWdgOImaB6lca1d/oqvUayr8Oj3ij2Z/Aced+H3lLr7sJi93+C
mwWcftNFgiMsPD/7NGYvjNtS29Yhtmg8ON334VZWQyZU0J+0U84MkXv97Y8oNAmV
o0J3aisz0QRrPxwWI/lBC89YeG0qWVlnZhm9SN6QhfD9SUnwl7G8WuZC6gsoWdT2
uidOrbkTuU0meYHCVa+DASSTn6U2Mdhz7PV53gNXw6fKETIlAS5dYx/dNAllJBjq
0fezfurdW8pEakGnBnHIGcIlcGNMovIlbmmpyosZ9EZL2FzrrXemhEP0/ZwOxfqw
o1ElncO7U/T8Tdfh1xv+9mX603TCxwwnmoTb0M0dLwfIiDbpvstGSzIKquAXI91T
baU4j+Dx1e+REooofLcBLhi7CFrh1jpjS0UcW1YaWB9bBbxiBMfYvfAzGTfxoUI6
uYoJkjni6lspk6kM9Z3l2J9th/Hxk1rjsl441rc8xJBymwWy18UKCLPkgu5cU+Js
TvP4WctTzePdqL27V4UyXzsqttcQHgPcHbWZEfAV+11otdU32tGxD2lOeFGFnhkK
wZ2PgZnqBkCxH0nBm2V+izTSH7jq7VG4TTwSljZl9rcSRBn9gLal1d501puklYyo
Lyt4ilsnYaJOKF1TDrxxmOqwhwoi5Vfe40DZO5SgoPtKW3aeVx4E03+mo1JG+7fg
+U4AMr6n5yAiI9I3bBEpb2XjZ2arFeAAHTQZ5ikQmROJ5eoPAsFYxTkQ2o0ElKbc
uHTCU5ioU52jHxqU5UysmsMZeV/piB06PM/08PvSO3LKfS2U8KfKq2lU6BFfEk5c
cQYmtLwZ/MFnaUYeDz4v5cXFiYiYuKIbrZ09UKbFpIt4O4bXRb2KORurY4QxOx2e
7K3Jubml8ng0jT/MaUNu2Vei6E2sMLNeF/AFj85PMTduGfKRmUKg5AeYz9Itw93y
SfGeT8X+nJOcoBUb6jaGoV+wZcZQN4arVr0iGXfKMopKu7C8iNh4nfVH+jvfTrJ3
RyPaaX5F5TnCWVlBf4soKDjKzBudRFoCRt3v9wrLe9URqo/B89eLGB1DEnYAkNOB
cfWvs9oIuJCQXU1pdEL2jbF03Hb+S23SOhJnOixMjKL7nZFVGqrl0DknUJoKZjNO
cR9xwJsplnSF+jAfuLpKmZK5wuYnyR0bBeTEPuA9XlWXkJBjZinbJxPuMTXNtzrD
tdszXF2IxiRaT7t/qJv+1JOuhIxCg7ZzZ+LwONslsIFRsZ7fulmdZyAi2znAxY2U
yWMZbseXwOaf45FXOkQvwJXiZ6cqDAkhEHyfNx5gJFt+lhRUeamNk171XgisKW4Q
9gpM1lZtYJJQtJY52Tl1UHLdCHF2us0eIWHEZ066LwdvGvmQMkmCsroeqzJzqhYR
uD2g3TQ+NV43U3eUIM9aK+9JC4aVyIYvAZ3NBUVMW8FRE+Uojyz2mJwLNiTwPXge
heDNYdE28kcgUQYQzTOS1UbQ6qclWSRdpWr5BysZoKw2teXQyYzR/zEm96OQlklE
pwxe+D64lXeBDghXhi2yae2o0ETiiyZw3sotJ7FtOkbGBWMB3f3XijD4gTvZEqLX
xU3FRtxaxbDnLGVz0M5q8hZPtpJPxk9026AI+fCaENvhF2NwdTDUMb0IXas8MEae
gT1/4Qbum60pz25g9c1PO8A5imlsUEoJylJ7JD3T7ivQOUgnoH/ee/ZVXnkbBBwt
74J2UKKOsUQ6rm7IshLrdxmnw6VGgUsqJeD4GjoawERXZb1AZeuMyf9FEfdddJwH
aj8eLbQA7SGRuc3gsQQPB+coSYOyny3rSH6IkeH+xgmXEnlLP3dTJpCWSLJh0N1j
jlI9dFVWPVajbZJn1UVkV8W1xju5LO2nzkdOFSyUKB2tELSU+naCo+l6ZG9xP9oy
pxPMYqZuS/6xeGma47ynK4jznUtLvPAVZRN4tjSfcwr+1kMFQ7mBcAyqiUnv4dBV
ez95E1OrduvWjlXEV0BS6Mxy7EQ4fT37jlP01FxZ4gHUY81WQJzlssT/Jh7AOMn6
Z/l5wNM8S1FPb9X7u5NMJgbxepeZ2/I2OiebSuEoFDxhOzprdI/ZXTR47XvA/hKK
3PbllKEDvKiEg7HbE5hdnNrpn+3EHWoZzA/SB+k7kJ4ICtVoox1t5TdfyhTNRDsj
i4524btxlEJnAwt6r9Y8A7V0ueDht+jwrUy79DP8lhfe6xno3DdbcRm8d6xqNFpB
dF2SrVHbWhOAZK5jZsFhyNjXRy43wYlKGxg1xNfpvNrK7GkuNvuhouyJReyboXS2
eU4vJwFVQyU4k6h38wyjYJHl1+huXWOtvUDJ7KKfmoUm6UWkcCxQN263svp3JYxm
hPRTukSY/L3uo04u0+HDUn8bpy0FDcDosvwRvQa4w2qZGoHzW0be8oJSJbcHZZE5
KcEqrXY7MyButCwLM9QJFJklIAQvKSOqDHdXOxDKZjjglqmxzGdhUlwJF+2t7M5+
hrEM7Jtm4t4DTsJ5fp0nvqWKkroL90fU1UVLwJMvhx6KNKCZ5asF2H3+QrZg8JHr
GM6Ymvcib327xk/dws9UqP68a8h+fC7U3dIuRMyvxKI89hUZF2sz/2dEtnc2ozwz
qDHSh8LGUmCT55Tw81XIZgdy4zcGCcFhcQUpNy9GZ0CFPa5hZDinqvknACWqhcjU
jMv0nt8BV+153f41C4dLvefOmANdQZIUS/SHfikRAyN1A4PAdmgD3vlLQXu5RVtL
bbEx2clA1kCJsyAFOLeQSlmWuVQAfJQVSnyuvp/Iu+1YY8H+GmAVHa67oqpx2s2z
3kDJ0u+6BZSaoZ+tQLqTPk+zqb3h6G1rZwYxX+mZZF4Ph0Iq+7VFmSH8R8NynxdV
DsXtTuxse4v5K3wy/FQI88ts7wFcbjs8+VNHw291tIhiVlh75+A7xbubY9Z7dqgr
BjxQWjrCok8+HdmDTR+DKXl3RdYskialkuNOWkGI5Ze6piLc1njsiCoR1AOPwy88
bS0oeoCYtqeJa/+uNYourXhF3zpIfETl/5wgp02NDo69rchGatJxfXdW/SMmPAsy
cmai+ERFc4bY3SUd7JUUzzxa9O8gPGMuDMg0o9+FzygBpAyrWL7iXGyMpZWgf1K0
fYSll58qBOLi1yOtAPmE/yhIkqeI7NtKRzesjTVYQLrzTJJCU7+713QUqAxys8Ix
lEP0sZmY+OC3V/6jalb7XBf9eJ0FoRWjrajRI+WyVRlfPvyds3D3wCWUVNd9IIU9
V/MGWtf3iE4JF3w+Gcc110B7Jhn2KZz64H6x4VLaoss3mfCZ2qYuDwWx3JXoQNja
tuV3PgSLJKcHYReiQXhWEJZFq/k5au947Efia6+V16trXhtKhQpIWJCUjqBgY1cx
7uJeNWB7i6HRTCanlOci/j1KfN8oEAxOo/9FW/kLbaTuRvNU8aBcnfoalsKlbvVN
BsxmZKSLhsSogroEBxUIEECSfeUZolim68onceE8XuBkdKHeUJopLf9saLGQFeUz
Tlb7o9DkLYeY08BBYCSbedcPDLR9nxPGJYu3fdSBetLQSc3Q0Z9EQfYXmoOLhrmC
Lbu1JH0aIlLOHtpDvmlEB+D3esEpUffo0F9ra6f3vNi/sXRdW2gon0L34pRvIdWL
DVBjW1t1A6yaK2MnUbL2hd+RGiGKG2zSdgOt/qU+HaMk4nrsx4SRA/k4DMoqbPIU
190siWv/2B1ElWb4LHhvX2+MWhnteEWZ/bWTIo0MT0Ee74X9v474PczHVPRArvy1
HzRUaScZHGDVQkNsqJ+AtMLqb5jxOAijvbcgGJ5lXQjs/0yjDiVIBBfz7divS3hr
vSeyzcXyC47UakadEeDoxSHot5Vsd8IEFdylUfk+CZz7aMarJW3G0+Zh8lm0AFRm
jKyEiXZmtCKTS2/DF4+k86POIfS9hpAHUANcS/tfhYXnbepc0apwL6NUL9t3zpJG
YKnNL5vOJttWsJnCoPfdp+pW/bgVamE3k+Zjk9d/oKffpTrXvStWM0tcTwyb6CBW
89xE8FUvhJvxmMsTxdAvKzL7TA5usGPxKW6+LpTNrasepM/GvDMplTrMHeqnW+3u
7W2w5qbDBVg9TKDSjc/aWCu1/ZvAxzvQ93aMgHdtzv2movCWY4Ob1VrVreDfqBhc
xp2HLwgpOyAELUu8GaqopLEcHL+wSm7/K4PtuDBWnoDld6/BAGRgRlIsFNNHkC+J
WLbGLXnutrZisKwd8LFKiC9tSqT/knQLwy2M+jdxoIX7a8gjur7gfwia63SA/0RP
FfeVM4/va1csfqRtM18qTWRYtt6OtWEQsGXihHu7vSmkE4MbLFzg+RyLVkNYXDui
6ieb0Pl8/9/XENjMU12AS39Q6C7EEgIAK8NykLzyzCzI+kd6p4cMWM+34rS98fjX
am2JuoyPouOrcu+OXH9pqiLKhWkHrVXDjUbSUDiwQY5TsVGgvBSuT2dWEq3iNLZ1
Rznv3tFd4dhenF6+P98Jucwul2+x8ThLqMEPRAYWQcJD47DyUal7cjnOAX2UWD3h
BjBcg6VaGpXwC9K1+4xpMooGouisrQ0gggHYiFTGPc8lT/ESDh9lIE3EjPu5R8D9
6UoIY+/IlQ9Rsge0wg8QVua2gak5057Ak0iu+uY/370VbCpTqD2pF3hYpMBpzeDI
sQ+2Av3fjtRGpZUdA05GR4dyPRJdEvyawuX46XamxUBYnkMQUKDskybujS8/gN9u
IWeVCuHSc/KMg1o1JPWUEmwoUnsYlth6h77QSisPfQRMMltI08U+bLpNT2XMcnYR
0vksyj4kZyVKmv/660a+yJYRr52M5io+l9p9gj2VMxVCwCE7aZ09mDn8FoLm1yVL
BNF0H8lobFOEYxDwIeMItYnYTR+MY5hjlVHQeb+u1Mt8U3QJ0iXN5fIA3jcrflBe
pKhrqJ7sCrTvP4kKkvWgYExopAMiNO4VO2wNJafll9ZRStMXJ3Zs9LlbFPu9JS3q
TNBHhNGK1cY/RKMxMcPi+G1s+wGwTQxLSG9yjfD9c+bCZhnjMemecn5fBYlnTT4J
zOQSEbjGv7Sq4wdEUbv6DICcWpij8eFXVX01dT/qZ3VqFXvFj3EQ2AF3JWYXSxcG
ZH+ht28r8Ffyg2OA6hxzPulBFi2lIMzbyX/AOdL6xXydF6Mzv4xrfUWiHOOhJnbT
tApiCmspeA2hJnJWqp0Zlxd7/x3vydKQ+gA8O63WxDrbDrtQEIpCs8he2Qlc6xR0
3mPAOSGACLitvs+i4NxH6KozbPrF1COZ0dODYDqORZ2ooqgOCS+Wwv1yvTYy1t0v
maqyqt4qMnDAgSmRJJ+xcivxCwCPteZvwEfAdrEjO6YeHNtw9t1H8PLjoFax69b/
PMxGS6DOmwk65c0AiTjXRuSvqM63W+GCrd1DSMVCsvPrA15KhnlhAgVB5yRVy6Q1
oHe+KydV36uixYWwhbGx3GUIf+2/DVIfdOMNIGuUc921E0qwuXBP3asRsipsDbUv
vM6+bqsx6TddQI2+PhMvDARRrig3Vrnr85MVy95qdHncJ7S9d37O8+W/qeDjlmQ9
WrTkP/tUZA4Ivd3Bwmp5YRA+076CVnf1VzO5PUTFWYyjUGBfWAL2MrQ18STjMBlv
A+v59ClH/mf1nEY15hPv/7OUhO4ZGwyKfIopKepA2K1YKJrDP7KpTROqMZCmRKRi
YDsDj1Y/HaGThKhgxwscB2tWwfurC5C17ODl5O/PnqVI7mJJWE3jhwnxf6qKJrnW
15pHEB05X3AugU/EmBvQyvEw+lYJdht3Pzti03s0MDvbnrQ5T+gKcBxgz/tbgyYl
MhqooeoCIlfkWCAdKmN2RQ2XxhMGdFgp4f/y2OZUhjMUdBj2IW6eGVI3GAq82r1P
RqJ8nvGjZR2y+uEiXsCAzLKQ0YxKX5j+0x+3umearZPMiW34LTa1V48IZM7etsNK
rqH3Foo1HypHIik5yw3d7sbyFnkMkql8NLuKkrS1kfIT1rRBnxVq/IFHK/isk3kf
u1qZDexcwa3lN4ZtFJQJ3myeOckZoQWgHllyW8e1gQBoetxCvZfcYZeCjT8k+ihJ
9y9BqzOqnZNX6nSL2zxuo8pDxgXYGVNuMnwgDve/Nia2Sac5r6v6TclSFeP0Yzrk
+tgl1tCaGVQ/vN4Fos3vTjnozxwopj4DYviQgC1mubm/W7D0glnSqBCROQUJITjH
iMBaPIGD5QuTjQHZRrIyuGfiz6hWNpm2gpXZHjaP68uSghvqnK1ORuM34v3U+kxA
USwQ1sEOuM0/SQb/xsCqYjFLqyOLWQ15HhNXNIA9+b1g/MDVxj8VOOyazdmSZjlM
sbFb7LsUVwsBYWmK9v/Qg2JZHrfiXYZdF/m+I9RycWdPbTjggakmK86wQrhylk0Q
aTnfQvsWQps2lty1KEfeAhTo4vmu1j+zl85sicpoh6sFlXN31TMA49vrJaJcrhbS
jtX6Y2fhNHMDIBafgijJwRlint1dJY1e7vusCrCaocA2PZf1gqYC24XfOLWEbC2/
HGhCw4cjJLG4dVszIRzYA5jovkm8g8qtiB14Y8L+heTOv8oezNW4H+j5uBHzI9b1
AAQWCxljl/TlhaQMgvOVhu2/jKZkePSaVb1INQzENGVbCH/xX7kTSxU9a39Kd9Rz
qH0QbCKJ4ISFdqMvYbP62jPrKTr37F2ftOZg51+lZ1RoltO72mjYTotrrqadnXEF
Tk/HTAzcJii6CSeXvziipbGnBkKN/wWFGs3xE+K0ojt+qzjXaYDRQ0nks9zr/Byx
kFvJZJoL62yChIkcZ0dzVXZWwvFixFVDvx2+4wnIIXNcKFVZLvs+VYllEA3MNT/q
VydGXoUGI69ijqAtYdo2e15HRZDt0s2Cg435Y5VLvF4FqPXy9u5wEVXQ6rd5LHo0
2TLwyhVJ2fan0inWyRAh/P+V7UHfeqsjNPqvjh/MOUQKgj4f3lUhGnQ3itd7oBnx
VZADfL1zW1cHQg8RTM6NmvUx0Fpvq9ajTkmXKTu+sQTTN8L5W5fmgwtA0t2WcS30
Kpa+ljjL0tCyBgNGpA36SXTJubmNok5NEfI+7CHMudAQKSqxwMFZBkRRwp/wQC1K
AgBVC7hf0mwvf2DhBv/g7W8kBcC4g6C2rcr9he+LlvA7583RnW8cyAULQd5pzv49
stVDERXhpmeikmBpdu3z0YJsulxJH85M4qM2MGAK1RRxdJL9711/9YT/VJ9cY7Rq
OLmjxNl0LOoZ6545bAHG4p91TWPq8aUGzkGdiQv2BA5HBHFXvdpLRIJig3kU22zI
k0AzVXuQObKNF+pU10l/s5O7CUC9+vbjlYXJm1vMEKOd96gkw47WQNcT0MU85ASZ
XbwbHxT3vlj7R+KmE5k+Nr2kAEfslvwVrLyVWQpJxm7EQd+8G2lBq01yrzo6/CV6
gPnaaSnS+DbexHwqAn64elTYxRC99p3OcZjV58GR6RdW6vd9SJXnjoOvpuxHAnOF
qBAJEQm8bjXGMhKNoAVruE07LaDghP+jYTd9uu25t2HJLJfj7pZJzAXCSr1f3Eby
4bGKcxYha/s5ZE2Icyf4TyJNaQ6dSIdS7E2pHsnLNGXARC4pdh4qUugtcMEd5lCe
e9dGWYqAKbuuCItaIkWKTpnDHKqfaUxiqT208Wyb1po0FdBHHC7VBNpHysfayWGJ
Lx9jxBaoY50lwdf+CavttQQIHdLRSVD9E5DlohKEy1aupwrw3iMAc5DcKKkQyxho
MXq24080oLOB9zTo2YbaOCu0rJ3CuNIIln3Y26Ux1XzLLulmstmr/7dPkH9z9ABz
/CwaLNqgbme89c7PDnh/OBFm024EJCHtRmFrDA+cSuNTSGRtMhQPPoP+RLxcWJiX
fpmmi90TG4yLlshL2JofrQk4K1tADb5DnJnqXapV5ibZBGJ0DUfI65GiChExpZwM
egfrYk1o7LkNBNoBl0myQU97zBcel4aXE5IkM34+LMUVBkX90YAApgRm0wiZUJqK
N83APrfn7PI2wlULk1QCFTo0nQhIHwgTBbAVB9ifMEnOushsIrRYGrbG9l2425rJ
Gz7sEQpDyZTaNQPrayyCC1Yx640deBHeArpIoW9vytvYFA4aTYdyH3OWOlLD751d
rtU6Ybr7cHIHd+eBD4uFpB6Cd8UMH/Smar9JKFt0Jik3UN/zi6kVJE7nzK8pC00+
tn587l5Ei2ctDksYmUgL9yEz3R6RQRqrb71zHwFN6dOBcFoN09/CUJvoAn2dK9Q9
0d6/pdB/i8n2OTZ20dqyHmi0kehWG77VJapqq1bgkWPVlSfdAdXXbdXKp7SpAiZV
ZjR27ouP2fSZ6LbzDONVK/28gVI4VcNxZA8WA9xWze5noSAt+BYMO2o9munThdHU
PbwGRKfCnDdCCZP6YGZBZpJzc0gkmpS1ykt6JL6WNEmjuelTZblZpvEd2SMnXrin
m0bkTRP3+JFjwXyvHQM8WZuIdWgQU2GZnbuy7BxY3+MGwrUag9vUhMg1FB1tZ4ho
0dQLUqTmRxmHRiwjraScQvVwu5IkKNf1vhANYFvrT2jymtcFjPv3uCWPGsGsy1bC
XBf3YRfC/+NjpoqSoLGud+E9uSRGLnrNRWpbtWfkq5+tGeuZpn1O5Lq0TTNv7Azj
W7rczzQ6YeHk3JGvL9nVHl7LRMFHracZ4DeU9oubTZIm20NryhS+Nek/b/hhX+B7
np51fuLHVs3oF7nlq5aa2M1ZuHf6sK+5RJh7L4EyAUoeJpsomVNKj8vtb04xpgjw
uHNPTE0hLcOa0gFE51+mQ3YuGO48fYkGfTrNYrY71oynrLSWVeHm/pSSqkjJOj6x
+fb3nOVSJM+7q8vLsb2WWMuq1eNUYkVFEdUkVgCmi5u01LPLSHSV4POXsa5QFxtw
vMB5xglCQkJDCN9EiSVv4wy6EPPWITsslcMaGeOfCCLBfvOtKlnHjxj4ZC4csXVU
feQHgRUdFqf9QwrfPTLAOtDlhD76fRmf9S2A8iE7wiKbYNZAu5Epf2QQ9wSwy2KE
pU288fTyYebDj+RuLV5Qd4ZE+QCmAuNYtpAxqZsEfHfu1bGHqvq6RerCAhFDNgWT
GpNKWfQGNiSgoMtu/X55FLZYwXca+kzfjDoajpMUo81T/a8qxuT++j6uBMthTTzo
CNV8I24XECVPTqK2EgdZ8GBQXkhhTFcoyz/GzpiSz/+arNm0WUfexwkluLfdIb7H
x1klNwXcHgZ3/PTf4N/ddcis9zVj+pEmXHkIFf84uwRT+b8NX241FWY7u/5t5skq
Mgr0Tuw9hi9sv2D503yQ8hkr9zOzH1nycmGgYvr24H4NSBk7VSetadnNP7QPnUel
dD0x7+8SuCkvDt52DCxJtsJCSpDBfG/4Nxeg0zd/NLTXRbsSR4UT2M058N7BhQHC
u6FV+4U+V1Glyrs9/OI88ZlU/NkIv4+wqdo3TvmdDMt9RXiqZ3tNiWIXonkdtp7o
H3T/y7Q4iKgXK6Kvvu21tZIE6Qa1uFP2xW2pesBr1GcKIa3P9v4S7H6uO+nHtpBF
dbFhO1lKZD7tTtAS0JX1ojR6XP70B94tmrDta0Sh1sop+MGjOc0Vvp8UgbbmhMs7
z7TtRgJWQZqODKF38Vov5oVKB2OmCM0LdnwNrKqhu/9Th9vHuRfBQS0BeQpKgsqX
2Ylb+mSSt0+gOl2A/TEgi6pLQKGFz9CNf8wxBEDQeuBw5oIMQpjz9CfAkyXmOt1C
fcYxYcFvugQl2r4g4m+RL0vATnus08HvRzq0RcPc0sMatZBHd5y1QKmNopF+gyT3
zD/brEqmPFrOxh4VVJSrArYhPYXvK/14ST/hdeevdYKxKVPU9+P7WYpoApvP2Tw1
e9iOM7TXjP1Og/T9fyKTVlNOWbpTFL7dd+oiTkdHcwXWprbZNJcwUiZDdUBcR10O
3JOSqv5tPxO+2CeSp6lgpQg7FLgSicDAu4KSxWba8l0PAPusbr5B1JvVSfEx1yPb
8kM8BWM3yGGS4CAP8Y/30MlPdIw3xbEpuJ4bsfEUhhRLjpw5TfjyO/k2DoxcWgdT
hI7S9JpySCKQM2lJFEYWRv9wLkM1eSc/grKwQxqZpFaNMQjUwJG9Z8W/vog2w1VV
BSSkaTqR1P1fBMKkE0UDo8apbiAq0ndXrhZbFZBUkOEbi3AyY5JMgNN/nz7UWLGO
1dyAt7rUU3mpAcHLKuRmonyR4te44bYjSu8hAYx4ZbyQLg5A9CMsCZstwhi0rVwQ
fy4N/hs0kwZR3I0OllNlrIWYgg/VCBNsrPaopQd5kIxWf9eY0lKBz4SHotlDhfi6
QSlrSYn1Sxd7te+p4tqZ4CO0S3T9EAZm+cMqBU4/oRa1SPn0gU0PCYaCc/eBXMji
E56DqZQyOCwr8IAQKBKJP3Fz4IVb4B8ykiqOgitiw9NbCKiiapRQQZ8hMSUrQIbh
x8ze4qTxjCx1/7rsLE+/M71SQJvRUiMm46zuFTAdd8SFfSBzx4B3pkvdQiNfcGQZ
9s9Tfzty4+I0+V63uM05nufsWf+wGD/18vZ8FvNgybuHqtHFOTtG5/6cWcSp8XDn
VdnfgmI7Px7Z1b+D8v+eJt9oXsm16eTJN/Flzm27fiqUbROCfX+ctLlYPVBP0KFD
MGG9oGh8d9JBAHLgSfZxsvPO1NXiS43wcQEbxquE6pBQoUJwkM5UvDy9ZjGD4L4M
56Cm1y30+ubMaVuz/18IYNue4c0CaA9UuezAuCneJRayowqp4C8S9pDHKRY0ROFH
EpfXHwqzyF+LB+BQCvVWg9XsO5gDS78l6/ICKlUsSn3bQ9VZ47HO3J1ii42N5jwD
2Aw28zH3KPFEonJskWF4G7nETrm7x4QFzQrqy4voYHp+cwY2S1j4hfj3KPMLIEEC
KSlhDklpZbvL7saZgRklZmTNVQv2J/HMpNB+oYYMA2KvG9kAdI2rCzySIk+LgXHI
qDoqz8qd884U4TCOdU27PNdHVwaoMh2SjQqfs0f6Eba1qkmOub//cVYSpLlQJ7bN
u2+MLZ7UkL3IJv4zurOWPs6TZ4zdKVVO4YGt7xi5rnYTVEVHn/Ep2zRvo/r2U5rS
2MvRmOGJprBn0kHRylmdEJ2LEl5c5OY/Yb6eO5mgngpbzBCuJlBOPl+VyW6esSL1
ioxJxi/yumssbBxawL6Zrude0/VVGGXXy7YzbZ0XluSpdZ3hq9kcMIDqZ3Rdplmz
yNAHT9CvhSR5zMHlcBNRAWQRH1L46JzVg3cg0YP5dLkoRQaupB4+HIxN+58dbkWI
/HucPZpDBd6xhX2pVf7KYBGqwyYHCkCRCbsZo5mLI80t/xVxZ+8nWkc/WSNlZoq0
u1+y0TSkBDsgHSYRhg9N0YRKgheyFrAStSyAkrWAxPp6tZvKetJGmhnIfncsbVII
HkozahYT5/I4XGqGf1HIZDNsd7RxCuUZPg2WFHvy6HZdMeJm4kdO3ndG5s8MDLfp
Q4KVj0x8cwhyDPLsdnm55MmnxKLrzhAWF/0SloT4XUynOpBVGuzslbWF4SS3cX1b
1dhYAj4knLT1C1phlxZ9k8E3+rW0L5NANmEqHlLp4OX3W/gCKhgkANmcDyDPZZFj
vn1qJR+sX8gFAFnemlm645G53jtx3D0QYhAP2hwL1YGKhX/1cva3PCsvCUqIBiXj
/A80tB9tQJsBQ6Qej9x03S0jVQf2PED39YbNM68f7QPZfrBCaHoiBd4N+24aLKE9
p2M25bE83t0w8jhHYHzeGs7cbVWldJlY+/KBnO9qXsbZj+Gxh45btcMQIynWPEvF
jKtrS1yNq6lCR/uVxUNkAvZe9v0fX1+42KMVyLa+buWnPw3mT4vYzJxb9YNzhupJ
pLs0wyJtoAx764XVOxWQIEQogkysmDQcxGIHu16q/KWTNRq47kSGhykxNyvOwpjg
8c1eHGV/ab5L7pjE2MjCcq2j1FCES9nnCVgbZ2SaG6IwACM+OXBSPKnCEnANODgJ
S72JQh9kIREc56SlV/BDgNLVdtt9WwOp5x921eOWmoWAgBJg7BcDaQ96RRRorX8+
FaeU4qpsvzwAJT0RU/t/qqa4uFb9/3BfxwxQtGqjnfR7ElwIVzE0TWPl1+uwAnk8
VAYJuHIg2wufJX3pZp5FxH/W5nfDzGoZlfOxdHP/3nXM3xHmKkHHVpvVdyf9/4nP
NvyaEFDmNxoOCaiFFGsLjl44XanJmnxxV793iLwqTfXq3iVYpJXk9yA7Sx5FnrF6
r6/+B4FgD3UNlBLU6+JMUgb2/XV5k8m1eKavIcNpSyRBJCHRwAyPeRJrJXPaEb4i
JOcW3noXvT8B867z0bz990r6ZLPHTnirCg4bZK1/CpY1j0eFl/FMYw4yePq9607v
BPQkpMOIb7RV0INBqqJC9s8GueUAA2ZATop/HifISnWZaafiONlBsXGCJhL12dPW
eqIGc+QBVqOGOLF9+BJLZC+VCe8PtWmbjrGIVLEfAUr4lWe6QDijpmwHwPqbcbb4
t6Pa9VCKdNKGshqjzicTZGDU+bYVzzZ2+9RKpCUshlxc8JSVbmGeMPRs5DMP6up/
RxpxniHQj5aWcpPSH0n/uH76oLUS2uBc2mqr1hMTmEPwXvdHxWXLCibN5Bn9NNkf
ybldcYqHSWF3CidiTNW8unKo30ck/2Jv507djeYM4c1Ds5RLdiCxR5jNhz6Ji7ff
QiZhF34ARWvgga6zA7Yc7E/MhDFalY6ggnlgcR2wzm023xzlkhHas/TN2yIRIPr8
HCHilKB7dYwdSc2ea1qkAcnNKXbXh4eIBlp7HRdU1xATOBW1hg/Fny6rMBCt54v4
/KuO5qlL5NFAb1mWkHuPmeEhdO7KLYjXwSVPEYv8J7e9cQcacIZo6lCg0C/4j4RH
GUuUxgX+nIeuIDfT0QWll2YHHX7rtIX3vMQZioLfQAUjfhZDwsc9jfMpOe6Dxke3
Fl+dBdNDpfIgZFewbTeMGmiU1ralm0VDMMUebUy5iJojpxJY3/hyLuP0MLg1tgX2
j3fd1Fgx7PV5sTmRAsBnkNEXPV5jh/dAYGCCRc5nKsJzwFbRBIbf9qulbOKDzdqq
b/A+lmZhp62tsbF+cYKfZJOlAm8lLWY0CGSKwHYr8JJ4hq7gKLLroGDEqblSoBqE
2+fR0hhkpUuYWj1zZJX7j4tcAk5ceqfswpKwlCN3QfygqtmflkwElyraHD2tELPy
d3MrGXTpBKUlSaT5foGy3uHQCoLnrs6B07yqjOcHVKywrNu/SGo/YDcbpNPMVV7k
dKlZjL62Q6VkYa1k+XnK+fQbKqYHssxsJz7c7f/3K3vJedmETX80rpF9IVzA+OmO
hFXnP9jMTOvs3CuqClXJKZ5gw+0SZc+KhkfCf85UlNHxsZBKkMUtD9Jea4FgRcrg
/D/pb+pAuYWbo42EUMZ9nIZzq8g6jiF0BTFNUy6cB7JD5Tmupf61qyVgOoRRGlxO
s48JzUUGpAYXPQr8A8PsUDgqgbYko7G2ondDGhkvSdbRa91OKfbtlXpSNvjjRK2S
Y/DeRnFEcMFmwT+VnFWTDl5XD5dLJHJisbrLiFrJs/gYSGL7axo0DWx0OfiIry0v
QILSomKy0AV8qJBdGm2ntL0wThkyZRHbg0LJBsVPL1h+ejTXrL9GWEY733IJ5+fE
4yuvxEvU128l2CZKWHpLnRD0jSMqSeb+7DzSRhrwZJaPLI59c78CtxH/RXfnzXKR
vMGGNPj4tiqORXMBFYC91eBkvxB1JBlbpuKvE+40usqIthW+uW6arnbxfp39is4W
Rea8A4BFikvqvYMqmQ/C3vhJ2oAUuGMz/eVqM645ucOadG7HEhZzo60Zb54s177C
kAkLlpXw1DNG9KPSPBaoodfK3d6kfS+Z3s0ElzvIcrn/eLxAcEk93Y0uQPhXavg9
5/QwYimLmRZBvVkLH6PQPr8VS6BeADMHwTTcgifoBv9OwgQMaQk3giYC8bhrtdq7
whNPv8DE5Ni+atRl2i1ELOUMms847TJylg/Qb4cQkNGlItzF+IChbdW9H9hK+waa
24QmVIjsxShUr6g0G17m4S4ffCQXRgHLmQTmaN3g5Wt7y50QiO3jyL5SUlwFjiu+
KB5zJU1Uwy2/PS1uZT7I0ib4jm3B/IJr8IoSS+a/zR0wA6FjroAOrFqE/XE8pU/j
Ux/O92VBwfg00IOsFbQ6jGwhYd/8p5EDrzss/bP1PoVM/x1XyEu7ECD5TKf/A88i
6n5aU+qtdGNVehrK6j9iVdf/T4Db/+daUNtG4o2+YHJPPNORjv8GNbFOSkjb4taT
ggNqh1sX6atLeRat5uWwSp99bOQoYLGr+RLbVDvVKO4nxfuccwbmr8+HVfKmn/GI
dgFG5fS2Fn2O1C6/yJigOJKaZgz/kkuRcS6JSc16eYkotPECo9lPt3d5EG6c4z1Q
cNpRMSreYKe+XEOPQ+L5CMg0SI8uoRG9pWo9WKgQzigxfSxwc5sRW0AY58mNqmmS
L8Wixs3p1pexcZWg6UDo0T4nYYEM6+ivAs2weHAvKfApHdlgyjiBs+qyP9E15qWZ
0LpQCmDCShn9OT8/cTz4Zz3bIIVEXyNj4s/NSsEB5cgjRA3YHODl+ICMLPzuwsuK
p4gNetObzBOPJmRY1A7151JxM0//gswkh40uoGagrDuJp9UqsO0DUO3IHXOp1Ju5
tPxAfbJmzyKKTR7XW5gwm3R0UBkZzDc0Xi3NAAYvspnx2BiJM62ImaXCCXaxKMPw
ddlVMJhzxzHfQJp6zFwag7W8uxN+adWWI+2UhZhOQ4u94b/FXiJzdTtFx5F1ufFp
h4VDC0dZgVXRfxoR6oG3sqzca8ZK7uQIUDk8wAhiZnmAOW1tDKbt2rP9Cbkt9H3S
K5h0MioMDij8EUR2zseVVZ8jk/y45dkzJGdyHLoPz1s1H+jpull9E0O+W1gRrTQm
GZuewaQLljWb/dI6ZvI85kImZpXpoY1zuydyoFk46/nBwxuP8OW47OMLaoi0zsTN
qfyE0kPRzDMBFUsUxO7ms0DATfXik0ouHQbntjPoxSuJXS3YI+oWB9A/W/+Ka2Rt
gI9Y2KDxyLSAFumJcIlD1yR9DKCDAG8A5ey73OlqXsuMWGxmpX13G4RUxGay3NQD
Jt4vZvHAPk4L7wo7GTnKkS+fdWyO1lFBUwMnuq3D7oYEuct530DXAndpi65rd2kX
BZmmeXhey0LxJdaCqNVj4AHfSTiGQ6kkPnY6I84yyXhrmuK/gQZRqlwSXmM30h0o
bks4cU0dY6pxmzCGLgcvd3RO6LoePkD8Sflo3CeW8qjw1eGvYy/FYUh7bEtKfn5s
O0WJW/6ZrJQ9rj3/8XwKj8Byy/c2+ZWoRZNqYKOF3Sev9nCwPAae0RpTasfNTn9t
crT3ZrbCrwmSy8CwATyBw4z4MZqEc8xzoaKX3iQ6oGH6wC6ehKXW1/dRM3ug4d+e
ZiSsKUmE09OuZAAcV5SLFTJ9kA7FCbA95CnJtN0kjfZjj6qs/8Xj5Q1iyIZZqvyO
fwghdev2Sr0EjXTZjPFvE+va1ZDpn7pnFZ1oF385Rm4b9U+mHhw1b4ny/7UFCWHq
bR9P9KBNN67IO5KIDm/h3/YEMRykAADNYzb5v1LeUhvo2zcphgVpxIr1nIuIb6hf
MFON6px8czTFy04C0m+SFFMdkNwonxRKQhWn9yWpnzsPfcnKkvrRs8HFRW/m9MFb
21T8WOD5S3+2Ls3mMRnGyV1epXnAuDjjBAcdmj/RC38DADOJKV3NFOF7Z+wKp3lC
Ujq7jruD3kswWT0vwhgLrlwFVUzvcZiXM/S6zZ0JGaOJddY6rR9eVvPbyAaIDsPi
CKyZ5ksOU9zLT7FN67XLBe8zRMeiShQyZ8jXSRQoR505J/NSxgCouI5JqYDJp/3c
UuwiOqYK3QR885kdQaFVFXjhYlswI7+iSmZWDW0vpRlAhveLrckbFZiMI4Dj8uJd
edzfLIaIoMflnR0qaqMVec83+xcnWyC4vcm5zkbR63U/KbjFo/mu0yysKFrAnLbY
LuRUOOfspXus4bJnmxdMMbtCttUm8W5W4Ucuj7RRlzloOkMs6Km7Zj62HHiIRIKT
53QDgyZUoS5CdWw9Fbk8Ys4w8pT2MFa2d1/sFxh33EU/97gQmcA6q1301UVQbXQD
09ok2Ox+uu/2+VpXvsv4WvOCa4BVOwQx2jP3y4r9N72TNmdlX/Glo2MWGGxjFqQW
UkMTKhA0K1xAQ9nu3loIdAamI5tV5yJteVpPw1CEJDyOpr+lzkcbY4FUZZMSvUtj
/vnbw9sfxsMQD3P7z+KNXEbAQQ/SR34RVVeI5pxYVFs/Jqa/q8//gPgUgf1TiRUb
l2kWIlF8ZO5mQhoNiQpyQ7sMNjV5SAsZwgxbPhrzgOVvh2eVCqoIOJ4O3ArcsX2o
CED1ijU5XbZ9EjXO068m1Zaw7icAU2AYQtD1z4sm5QYoFWdctwUgKZY6qxqdHuih
lT1XxfIJQ489Z0lzyH/YHQvJ8unbyyCa/KwmxVyKUeGO6+HTNhvV11SntRxx7zAM
/fM4KHFqRHgoF5x+HJ2MED/zPX6fq30GXAjC9p+rUxStMCUD0KbWH0KRhCcRB1hA
PhoKpUzkzCbEs4yJK7sI6cop8abgwutyMNEfVuyqIF5coJp7C8EK+VmqDAwLmoI7
40ic+JbgSqvH53NvxqTJvMxlzM6OQ+2TrkUTfB/0EbO6mJH4giijIph1NtUTUQ3I
kk/GS5Y2LCrdNS2MahOjFvIlECnCJxRqfVVgWDbrz/wycvDjmAmb58LvFaac97ZP
fJntfOQmp7/Itn+aw4NeNpqLdyoNK+YzDaZxqFOTs67wzzqmv4N1r1hDbbMqxls2
zQkxd1u+q1fWP5FJgvnoDZv0PBU040P7w6eZaXMVP/XY8Fyskb8usmy8pnrUGgv/
8fSBxhbwfTV+GWrym/crTf3vB4bB0uYN3IleGDliz7oJjKwygW4sJ5Y+0hl+4apV
DJyDTJzMFVkbHFYUEiQM9osIZ3De63C4u0EotWMlsPj9XeEhNG9r3L2zrEkUYR6z
4yn1GnNE6m0coVHMNtyTSkKF6zuGN73QejnMC6TEeoXmnMd3ZDpfqFSL/BL6jCDu
n6qT4HMbCsYldy7J0mF9wc2Y9DItJyUgIlscwR5rr76KhM4RwzbZvJPxlWZXt/kM
ayqieHlJi78p0KHFQzApyWrcjwQ/US76STnWRa+WZFGOpDalPyulg5l7AdORziYp
8bfA4z5Xd8FgVpS3ha2hP3tBQUIN0jT3mNcvA6IOur/UEc32eZH7J4mgF5/uNv2P
6vfh7a9WQFPz7QYrwOPwD4P1eQM29ULqez+WY43GeejOhD/NMn+/BR8dTe6w/H3p
cOdv+zTRyMghS/R1kRpb8qaxfcQPM1COPm5fCkzw4GgXqJfuMkf16Aoq5OO0q0ua
Xyq5v8A+gDM3XqaFpCUOOpSLnrKMkmUKS13aRZ/LZfC/YVSAHrado8OT3V09oaD+
9CGl+8rFIe6S3+g64gyiALsWMuq660cNJQbgwJUoS3Hev4e07H5DKSsnj6YHgqCl
9/3G1U+mlxtu6NGUcYQzr3c5TLqXFmYma/jNRAx2XfdAx6iCalRPo43JOGfVhZD0
mHfZ7Ds65/Cq/8ir1sci7/jpFuAUah3/egImTERvJgTM5eeL0udHrLnDsqeS/WFh
yD5DeZLe0vgDfXRzITHhrCgwt6JlxgAEpzU29ZGW84fmWy7QKGWZ4kmU8WlKk8BX
kfzwMf0Xw5nlM+R3R1IPpWLlmqU8nzhCiFua8247j8ioHWYC0kOEEBOihMvq6drl
/nDqqoM0p002HEEiAQpnDLTfzvKPIsznbOV2B2xD4oegwtvTVLIdzSGs474IOBJs
oFdtYShrA6i1xla9DkTHoRKCm+jB/3zB41hbi0PE6nwHHlnR1u6SFkrsWrzeqwoJ
Am008w1RpDmjn6pMRaz5e/EGgomM5rDxLcb5jTKQaerEojNdmsI2NeZdCqJDxiHM
USTMEAZNd7YUXdqGG7zkJ4Q31RO1j2SP4xwQ7ZkeLK+yW0CpwMk9q+2y/GvPUdR9
flxsYfluLvesK3823/B053frr49FDpZvF5Q06sb/9YbJn1jM5Ji9XMDWCFeMb1OE
nR9NjEKZS5n0+qxlJeTNr+eYpd+qrzgH8DgI7cshWO6XVbTJEoyYF8oupyMZFB0A
JDRfqgLwqOukB/FP7o2G5oZHivoQqtSZkA5FiJYLhMQCnXSoMiTmcoPZBwTByxub
c7FXTJLyZ31lOO8sVtiQlsUNPl58kGQSNjE7QGjwQek/TgQrEM1Bc+EQOSl6cjcL
gfvVRFTpdq5koqVBs1LvDq6+8LpCglgj5UKkd3nROqWmrjnbAlNifSF7IFzVtAe3
8lCtYZ0Q4Ijza02mgtDsE6k8bcCxbpKPS0vj3trPNcS6bG0+GeIqDqnXVZbVO7iv
PRe4LsD8I8UjO4P3adnhKwJyM8c+XeJvtRqJA9h+avmre5FRAVugDA3cR1665LFX
eRD0pMyaaXoCeuu9BYzEj912ytKtOMYER7ipybN0nFR4478q2xXvZMPUolAT+YgC
tzUcpvav+vIVFv4CEduLc42dM9nwTWuIO7avFplQxxlz1Ji9o9N80GwzrM74/cbS
DxawfYKC+oB+HeJt2buMMfDfAe8hDJP2HYYKfdnBbPJTK/5w6V3toJz9u5/1hKf+
C7N942B8g9mc1vnNTKpgk2j4k2QMT5Y5TpeSkAf5Sbphz04x/FXS4L3d9oVSW9nV
8x1XozinvEEi5PfxQ2I1PfI6RvngGOa0V9HMSEol65iGwP9QV//q3y66WPNdTtOK
j8hN3nGLq0z+Hxye4CTThyOHB0JfgaAo+I1CIT8B34apkPa6gk/7CFIoCtsOau9x
BykuV4+GWRsh7HmGI0NlyODYJEP7Fn3dRjTjRYaS91D5dcYSIikDE8vTWR5OV3E7
gSWvTmAOBcZ3CRR1fWYfyNmTMEoMiVf4AGJTGbcePQyPbX6Wld/3MC60nriJPOs0
IxJELrVN5Sd+rXa+R4v2p2v6qiUpIuH5MRUXAXegop3HTUwaUGvndXQNLXu0D7oN
X/QfRT1/KJn/syxxsGkdRPVc3ykYkc39KG1WtZUX0UL9e6liKEqtPDERaZLO9qQl
Spuh1oOZ2HjufOMtlULrFyGFlZVb84p8nuhog9KDBJ3RmqxChtPFwqfCs1n+555I
Gtofriv4bq2xCiOSUGPRCm21ia/T5y/YoMKRSQ8F3nqNnGsW9nUxJNTwe//wVSXa
WeztaOLhoYsTpl/pT272JbLmVoHibMYWsQxVlnL+4M94rvmA6SiCxRCPuszPKWuo
Jfou3brP7XksGI/MP+RfRfBAZnHjdN1K5ulJpJOWkeMPWSs82y/PkoNCPBQMq941
vXT/mx0/ecKoajrqczFutaapi9fCsiDpiXCc+1FeEtdcR2hfHA+zILAXzovPEtZs
TIIuLA2J3bxeyzE7lPe+l2dNOMUbxca150pBsPFRIi9yQHfp4KrccJlVqAD/GAL4
bXFEHRvuLLm7ieV41T+YCe3LMryBmvfdZyjBQkATHVZmU2yWwgC2vkkgE4x9Ws0V
kUI8KjN9Ps7rUBBM4R0k26KOr+nv9J+DOdt3Sq2luPdwcsOicaYqORsltNT7/jAr
6u97nebkzVWYnXGDDvxeeg6nOwiziWcjclPX1u0IqiTXWU233wi3TlJHVO0io+7f
UOYTa3cYmi0y4s7fubHQyaWd/rZPklmRyYaXH55b0TEokMeHB+YO1s6rsM2STbdc
c8nQasykwHp9NIlyYSjwLZScAn4GJzbcyBUXpog/kGpyYNSWOdk1xfvtHhTez7hR
Xik0GfD4UZkTFYGeSHnV+0NluF3UNEZlx442ZYNv7Ci2/uhOZCFVNXfJIFKmPyGS
IaOTtPHLU5ZzCq2RPyd83WKfOcYEL0pFDkTrAGZ4usxH0VdDpIu6D9hX1U7cZ00F
kV8KMtugt0gipsdiOlz9+fIZfJfjw13OSaMP3tWUokgCeUpTIo1qWWhJ+mP4jPig
6WkUK8EdfhmcmdVpfPXr2k6l+WwEyOvTyMu5bUiLOv/1D+U/k0mLaWrywxNjFGtZ
0ajxIS51tChBP6/TV80jwuT4D8Hl9W96l83tRNjEg//N+s3oT9JNdzqx1755aac6
ZtVvIiu2pxNqT5qX+W8yGstVljaWWWerZiBonEXXFKEbUfb7zd4KrQkAqAQXJQrk
ZBniUcljjvi4JXrdRSEbHZBu4qcNT0fhfTAozs6i19qLlBx+tVaVU81Px+beKt9n
6QpRF9P1OQsZnW4OOScvMWHxTarTOqiApmS7LOE/BcvlcQWPSHIraKkdeIZIeQpK
fLxI30YpBF/Qigq3RcGieJYjPwWI0LEKQI2HGCqCbPXLTQhMI0sEeDhMq7feWyq/
8dPRIXvLSBIZCGYwu+obX8Q2qXCOspmBFyelIXSxoOV6eBOfY+3Qf6HEuUL5VNew
FOrmr71hCmb645z0Q/QQRWbJqaKKzBlCeMGGUcebV5nmQo+DodHDdE4GeJ57Am0f
QATcddhSx/vuKyvt0fOsjiqQfz7DdB7ma5UXURMnUu4BeiKmjXaZ0aebCpR1z5q2
a7hFMCRymQopeerHlgZ3z4FXrqCfDjyvF027ERNN2vAq8hKovEmvW4KH93M93NSv
ET6oWXlUrlqcNjEemUZLfvbntHLgTZAC071+bBvKuqgrrOp6cCJE4A0af06mYcH4
QQbEpIPtITHhpgpo0ctLIGEayUqXdwmyx5suGBPXA/2cX4bCYJf7NvLC1uiWAp8c
FZCTgU3qBmTee9hdYQ+p8Y70BzVz21pexvdpWdxfxq85XGatl14KAiZujQLlI1Ix
Q4uKr1F3a//eWrfNX2FMbEirjoJNohCRi1oP/U9Q+NTi4TUntOn2qAX5/B5A7OlT
tPY2LB0kUuS6GUEkNO3jlcVpt7unhD1iG/h8CdomzV7O+UNpgHFUl/C5wFlndrKE
YtT+KELhSzAUJU+5PMoOwldS5QiLkVSFbn6NyGoEmFMZzWep72bloROkiXRNRQjA
MmnPa7FqLEWXW6UeZ7uMSvDtQSRs/1woT22m6Mnl5738HE7+ffJlTFdbJpcdMsp+
2t6nePtMn8H6yDPPfJyxJA4ve7AiGE21MD1sLWTb9axzo0Bag/WNWn85zeLDlk+J
2RvZH9VcuVQHJ4UjiIUX74qpWWlbuTKvmGWBG/8R779m7TryU3LHmmtNjyxGCPXq
NEZTFrMxnShVBdFu8LBsBiHPoWi02i+FqRA5Co70U55O+5CXimcoAJfzg2j9x93M
7V5GutotTKw6IR7AoaaJIUpMsaclnoCNxZY3lkjLJ/r2hzGpJ1C8kjBNHjSHctZd
BXWnlNZhuU/AlTLyT217Hzw723gyOv8XZny/GOIJE1hoeaDiGr9c2dgX/LWWj2w1
CHiY5OWT0V6Fc3Jk6atKkxE3iDu+isoXMHQKVI7yCVogbJqqj52wiv+gX3eZermP
qiRMfYo1I8Ly/6ekTMYbECWaxAgqpnHicxb4+hU7vIzSEoqMBBJaOSIbYuuhnd2R
B6lrmGkiP7d5UZ70JRXKo2+prbPE3WanJHPHHS7PDcG0YkDrUSxrGsy7Qe89DsdX
HwEYYxbgUdNVKTwn4RJRE633ErFkJMEfyywCd9Torfzs1lHD1wvdFBsIpWo29ZSv
3gjw4g7mm56Eku+TZzjAepKnV7XxsCaM7eCEOSYoAejeuvtthiOvahuqqO2VWszY
KsHECox9japoeOsbSET0MHDIGpZYW7LXSUET4v9OZs0s7/FmHxMklmypjalj2jU7
W+R34pfQhh8y5fXBOTjGzZ/GnnG88p2kwvL/CGN6bo8eGVwWLbJhpsikxtlm8J7m
MTIMsj+9krj1vJZoVWrvDlzyH1pT7OVGArmGuZ0+AjenaJAw3vmOD9yP9nLKhmfR
fXCQP8RLsv2Dxf91XZl5wLDIcfqDJsAXmIgIF/wzI8RW3izuG//OlIhIm6kFQvMM
g2xX1esJZGYkyxukNHhtS5vNdbO270y4PhHGkbqoiICypD4xVkvPfOndWDSYDJkF
KVps4ftr/kBREcjk1oMlozeyOoKYpblIbmi1w+O1TZZUrzVohPCsYOph5eCD7zxi
npC/Jtm8K8n6gHuZPBInZKlXWlEtn5IXm/Oo3baBpjWLAjMo2V6h1urIwwKARdA9
3f9zx7HUaO+4Fh2shn/BbjvRb6oap1sDWz2JKCen+c7meYI07EK6LIUaSyxGTOG9
hAVLZ9M8yajW5N3l9FZ8D9NSjgHEThxIgot5nI/rNIG2A6fCclIENxOHTuQFFdUm
DrzpbcdFr+8lgGUtW/X91Cj8FlFGIbKvQxvdL3J97vRIMk7QpdzlcAjeBmdBXESH
7FaPWuXCYnRn3JGBDHYEkDqGYDSQHnW2Lx8SPOkL917sj2GiqLphFu3XZ0MSBdgF
QqZZLswfvfEbtyGRRaBRtYoKGM4JuofBfub/f7FHWHLsm7hyhqd6bG3Bh1dqPiEc
/6AijQUrjEF4N+vjXJLrQvI9PN1Vyw2d5lz012UXBJXOE04q/n44qLRU/wcjyq7m
CXF+Lz9d1cCCD3zdvk0cS1b/gPL/SORkXytRyzV1zXA0NaFBCzjjlqXHWFcZKm/1
1yuh0jM3pNGwBJueqL6HV+f7hDS007Is/vIpqoY2FpdNrqa4TB3wSDBTN5G9ks6Q
QKJdTsZmrvt3nFnNU2WaNQIm3nB+fTC57TKz2v/5b5G+gMPpcl31cEVcv37Wu2z0
uqBtROWLnbnztAA3+msDbW7ZU1nTy5f6YSBbjJd9bwicPizBl1R1c1CuBnWEVKzB
EkuCOenmRPRKPBOeONkX+8DH4kKw+TBW539mPI/HiAunFB/t5KSFErF/eU3hEuHL
+G9nMCiT782WrAaBlxAto3MQeizU3kLBLh8yy/BNYBjBVow0/RoWnFuWHyvEG+SG
OtM2NHdTdimAJyt9wjAkqEt0RKccGAo5w+YigGKCJeV73fWgThwl9oay0cud14yb
gZkBOFvN3/Wdk0+tVGIb+94pC8W7EWq0xhCqkEi5cHKkOGM6pmuaIEgk7NyDAwNr
/xvu7bSRV+30xeS2klDFZI5Hb/Rto8o8RiZJh2D0XbdVWaBFqpIh5ukVKV6QSY6R
yno9CXrvx/hHTl/iLWjY5oYoTg2aAdQpOO9zxvzQnx/YP1hHCTv1220tQtfIJjGU
+phvutNTe52bD9PVtTOpbue/i2QskwivQAwZhVnMVxPCyzKQj18Hhq/teq6R8Uca
A1pvSA+KTFyzYcdo+FQYBlYZmksN5W7AuSEuS3JaH/bFrbGIQbWoSwVDTiZNy9qO
cFPGAjR7/HhRV0btmcZFZB5VubOCV0YlrbPXPUBxNG30WnAnz58IusN5Ex5KGPnY
eUBc2nsf1cvF8/RJXBUO4GU0BXrGouB81hnCSTEMnImzpJU6nOXz7ifunIEbWTHF
d0K0cJZbLauQ9B4Bz5e3PCV+JngDeyt+ZunRlOvdIJuWzj1SaSUD7d/6n0AP88uj
7AsEZW7EpYNnqz5lW5PplrgPPUXsenCHBiIFGtjWVzyt+q8PZXbre6mzqmSIFXPX
npIsJY+fhNAJrx+PzzVA6utBkzIMa7cwocNcp1Fj79/gxejRkJ46CoUr8U1igwXQ
F2uU5fBaG6h9KwHJWltsy70gn+7tQ4u9kBtDQSkv/Anj+c737wRok1TJf6pp/BPc
ddSKMObkYc/O0SflFXWrU9tIoPAP5MyZRO2YLur2MPDalUlzQ/5AVV/Z9L0rgFug
DuadW2nER73PCnXrXNg1s6Z9WAjU+wJ0mfTjtkveVTwNX62eN1GeEsxnXeEY4bRZ
Zq4Bc+N/FDaPWsMOrbRvzmDguH07LdUtcO4eIqf8zNI0FlKJg269aSYlr6j32BoD
jxQVkjRKXqodylGCU9X1JIe+cVsgplLkgcP/O0Txjr+yFbIIY7H0F5Dyl57DtisV
Tl72uYW/wLo3luZRoFyiBdIJAa9dy9dixnaTphT+uFsN8yBgDrPH0iIatAWlWNPz
czIwuyAMT4ZyFnvEY/RAIu60f3VbvaseyUySUzXooD7cWQW5VBcaCeQ8FtPQVOBa
AeYDVhfNVigy/TSaaaY5z4yfxpXpBTs6KlR4LPbIYkcledduxOMrd8vUKbVKxGcw
KHHJJB7ZrWMFrcHjCbiGAMaBGV7iwdv2zK/MCaFr8N5w4bOmxf1r4+i0bKnvT4V3
1AdLCkfMTqSofhDOgHOK58b3pIQfmKKnClQPZWtErEO/9OKr6N55FOCVtzBKlJoy
8sa0SqRet22qfb4Xr+qTWufKb87ni+VA99RVAhMjE6kn2gqA2LgpS+6aZiaT2T0w
52mmi2KiLCVGw7X5lGcLY5WOEQm97Yj4ID4mcZbj4AaYQqTMItv4UXSkzW5AeWG1
wECv74Ig5TiSAmLddiQKrwnLfwxRvT2NbumcsTElTIXvz/efcV2hLsGUa1p7YtHC
azkS3tHjG/VzOFNe7jDf9f8aFdwI4LrYTXv/p7gMfPij6/18CySTkUjRog885eCO
tkfRDP93IrXm+qDy3O/Dmgw8ix0NNnbZLQQVRx4DSGG8YZ/vfkshiJMfbbY7G2Vy
BbjP45j5ioOPkaW0p4pasZ2376KdiqmQi4zdcNDB4/0xWaaoQRN64m/mfqQp1U7l
vU+Wi57JRyV3M3BekyGSEsdJggapvDaib53LG+6GgBOtXsw9edvijxmYeSP/gztT
FjRoMPX/V7WSrwTMVKbEan9hytj9U24RYjcZPFXzb1FfE3nipnXc374tZ7pbBhOG
hVAXvj0TP4EhbAkHPmmUib4XPU6DIbyhXkf1C18uOZI80JdUi+gpmDskFqlJWelC
oL9vUm0ZgCfqv8PbhW1ER2gwz61VHdX4Ydcpz8QmFC00MDln14hF2q+q84lJz6tN
4nw4vfsT+XEDqYgdquNpIC7pRCXto+4RXwldmCqevZ9Hi07iRhhGz1GKfKITm9aM
j5g7bWF8PPM/dMF75yO2lxnccLL8R0p78ez4NDYdR+8VDIOXfde256LXw5sHtAky
Qk9+a3hivUuowTElII9QJ1+XOn6EjAMo2EEQk8O6wYanEyoBsTQAfZ41jNix4XMQ
5Dc7ZMAb5FxNbzK3HSFP34J3p+0Kg42YeCDg7CK+oKSE/LecMxKKeFL2L9hKR7Vm
tBQc/YDyHjOUz9XC0r6rqhabSFRYPyQjyZGoJrKEW3cbNAEOFLDZypmvodGBJES+
xg1Fj+6S8aW4dznXj1e+H0ks6PL1JjLU/GosXNpTN3tv1AIOrpXHErrnt7JZsOPX
PDVNQJXnD35gwklD/wrWGMBLTRprMs+Nc5kcfnYyiU/LfzreYrMkoBKFOIl/JIUx
X6D5Ff6hBNY6G6uO85XXnyS0UrtoUzJYTt9GsDFbOMj1hhGuX6oduhdCrcAV4dOn
9QszWRX6hKVtKei7uaOL8MYJHy3kD9sezIbIw2Weeu3MB+aTgTGP2VA8K8Yz8lD/
XgIw+yZcrOQiBPyQCrZQ8s3W0L7uoSlsIqTG0vA4e49v43sWmFS5AGgxH6HZpEni
FJlOmsNfa5QdcwPRVfIm+n/Ppj2AjJ+9Gni9gGMWoC56DmKwwJY6/MXsGke3G2a6
t6Yu4QvZ7z8jNUnip6QC9lPJELZaDk5lM0ObxPpK/H0PBwqEJZSBs4BN8pEEfxBL
/EIqF6ACT9zgNmygY5rk+W8AY0Il4tzLFJrbKmS26zGl4BBA2bOsdBF0vXiFHAmm
tI6XcKiJftYUZXNVcjZZ31EYUsx4CqsIUGwUnGi+k3O4U2bdDnh3lNa6OnNMeRuW
EbSyN6r4A6KZNI2GwUhBkHblXQhvy74SEB19iP6Ns7R/0p0XbWkPR4tWBdZJijKR
0CXbOTin0iivOXBVZPlhzzhA5pIvkQaX8rGeNtUVzrJU2cH5gFhXFjcNPl7wSsr3
Vynxi9nL9kqODCELiRECzWbBVKjBNZmy2JG6t6NV44IP98WKf3Qq/Y1MkAIiF6lu
heCVv6xRbcFCCEEVnbBAoI7Otakn5TmHqQTjCaijzJdz1J+29stawGQQ/1rTKXIL
3lCk0UghySyeCGFla3yfgLmuPwWBoVe7K7CD9l6KKRwFvfSbg1VfQqyPVR0Nd1Wi
/uAFvUwGw8kp0lDkx08I09+IU30P2kzZPgLvlc3BJzY50kYY5yfPhIXOZFDmRkGp
rQfM2N6WpQ83+aiCEYAeDgZ8fae9M+4yuPs5qh8fVZxYQ6ssXb3etR9SfnJZFEpf
jlUcz8uz9jBeBeTb74FewpknjzN7mb4RsM2Uc6IqVC7nhq7HyrBlelIx7xCQ3i9G
hLyyeQQGZchyB27XbUZSXg2O3BbSUbtdjUaV54ZruHsCQRLfaH+bN4i408gGcw9B
SCxHHIxFapfTWko3EwK97bEto0gBnKAgbQPTZFSGKKhiJIWuoi8TpVot6F1UVXlr
+MEkaOMySFRxStz9CAjQ8zQy9lIkr2emDfkSShwCLQVSfsTDG5EAJChh+P78GkNd
cYjNwBF7gyLspbrvyC32xiXdlsdfXe3sz3yjBdcRGhSdMWoVhGXunv64bZOss06P
arbXXsSBHrSpnGox5zukx7Fet/BNt4uZRduXIpS2yeN7hyBQObE1vOnnkMpjApIM
P0y1NfPfSmR/KrgGpVjGHWFFp8bHeoFV30RWDS5CE9xCnbbKkjHjBMWCMbWqFiPa
TUutd91DzNlzrUsHOjyuOUUJwzhJwROJCRtIGGc6IDOg6tC6L4HmIXKCaMMxyCvH
b+eDmhNCnb4l9IcLHmb4mOVtTeCX9nFqadbY0KWUKBJ0k8cXMixBBJCJzu0eM58c
cLXSWSVO+oA8Guy9YDw+bXzcf0MwnYsM8CL5/KzJST/1FYH7MiH4jp/wwvL15CoP
0tRlD2tBNO5tFpmYX+iPL0v/CpBCcAFeKs3OYg2GQyiYuqhO+4+Wllm5ZvjM0EpR
Ek3uo2L64l6a+ably39gyKhIar1GI8G8njgm0iAEQLNrVSTnlH4Af9q0Jv9+k/s0
wxFibwWasxGwtE4QvPy9EG0HkeXoKKnDXRuO8hoVFTleEaeqifZFgFmSykA02F85
26vp5k9MhgVSlfsahU1+cbKMTvFceh1fxBtapDbDmlErNhya6ADhPDB1JO/lt2yB
SG0KJ8EauXuG7tesC2YO3p53kVvZ0RViwYurKFGPUjs3vFhYYChUCgthgaR7IAXY
z9R6k+DxpFCUVNtfwJdL1jeMjbta8jgrv+XDRYY/wTMfk0KaOZ1SByPXcjvo3PPY
4rLSnHG8FjzKI/FiPLfUlryRWBglLdgeRw6fidYgpj+/vIqyu8o8qqpS+oxtxQ2I
hvJ/1gMBm7RM4PObM6rQOzHX3ankP22XiiaHCJeiZbx/8humMiFIVsPEHwVXDdxe
IvEnWc/kfI+Z7TB9vy37+YquMv6fP6UqBYDkPr/y8xw+Z/00V5gNv6fV+9j+d8EO
u9NF4dmSAkynViEQQUu9TlxJ++m/fgUyxufOtRZ8p/bILsgDjFHTh1TaHbMeQCN1
jJoxjLAHtRsjB/tgkY5mwFRyq2P+7C8XuVlboEvLnTvQfWahsmmlBLEqcbcVImXJ
QpE0rpQ2NHFP4fiM510COn4gp5tTQ96zTqu30Ww+NEWvtEx4MiZFgbzdaWfJCH8Q
weJgsF6f+ijyNYipzXNUj+RwqOzXvpTlJE3bGVxGKM2gdE/veS0UwHSrbYatmnB4
qSxe+M2cPmGLuGRprE1foTG739na4MCZbpJgHroC3xj0c8SWSt/wSuRvolZhD0PZ
V8pytpsvWgogKV+dp3j6Mq2JB0HXX0BeEL/IajljHbnJuzGhOi6TlUp6P9ooH54I
wFAhOCgG1wQP+Qtg797BPHCT6rgb8oGGmH7gJG+nON5MJVUN4IxUFgTahH7jU+X2
zJhMT3BTiG+k3RgT8nv/PRkKgIFu5JuX9FgQDqRJm6FJJwRLXFgOtVmsoYgShj0y
u5NNA4A6JrPgnt4gwFVy+rSjzwQxc8dcAPnajiA+JEt3MwSqjJvMeXCk9mO+rqZ8
MD+gNgBDDP+fexjclOd0+oo9Pr34m99bw9lUhrPKsgAdD4yN/Qufw/9bygy3Xt+x
vUvKBYB5ECaEstFrQz/bE3w43g7fntG7P44NAf5o59uporjObqEeJSy3zW9vxopo
tMnrXVXDy4kSF/JiKHMZl/vEeWPVrFcLbnP0WaYYaCBE7aRSJc9bQ38Ndzya4Rjd
GH+fJOzAE0Ipm1WNED8Zi/+Sbs0CqARUuDR9mYkkI4coxsmUOoV52cTpzYX/lM2V
K0cOMItUUxyBbeZ8JIRZ1KkQ/gRo+V1tS1klEVBn/W/5B3xRFOZjRwoDZXcFWWbg
6n/3i0Wd1Pj5fAPpOfmm5czGBug+JJ/Qa4u6VTzG5YAh41pMyRrD0QY5w+5DGyb+
l07JaMwf1tjw3VwkYKech7VPEe3hAmHNv+9xT4j9/ltmV1EXO7ezL71ORti+TJjA
2pbSXlJRtWpeUdIh+LNLvjKqjiDXD5Il9Xa4nru70wxKoMcLIDY+eGDu4A17cPuL
8nx0nwLMupdAgMvZSGr74jYvBkeppQteajCLHxytqYu2Fl8G/D8O5i25poxClV5b
3W0hyYYx9rrVhTO30rUYdRWoBWVrPoEXqb4ikFvWBcLhOG6w88uHqOtIGDdQesUz
JBCIckQu+Noc44L8RFrgmU8NYTTFsN4jzTicLQbchgJHR6NtY8EcBRVh3UOrUAiT
A7h6tFSN7GqBzGQHLrItEWZCu4+KROTZntxH6BlA45YQVzi9h6vDDsYWkAuVNSWZ
z36wTCIqDTQrpgT1SI0rttSfoIOc1rdH/0VYW++fCqbmvg4TKcg8kYbNmOLx9WtI
zn5ts7gUP82ou547qgB0c+wwds5sWPhqJaN1yCwYWkvRobN1nnmtsLDAevzpZF2T
TKdr5m/TFQHyqri9BBmYGri6qCy9GN6g6/v4QQkZk6DcdQKktB1rbTweDRzt2G+c
+jx/BfImD845zBR5vzUxHtteHR8Oi5sxjdkYfXSBrMfxkpS4H7kucdF97tJvmEit
ikFOya8mDHuR7i+evJQG4xyEWFLm6WgfP3y8gw4/0Fsf/gquh+QcIkNlnGjBy+XJ
CdPRF3nUusXftJ+xN2vvHaMI7D8VWHCwusMg9XIb+xXGyw37SPb+FHHqjsGsLU2X
Y49VtpzW/syWq03GLmR3s+W7hg3i2MEJPOiR1BjGzXpQ9bt5dTr5bZK6lK5uN3Ll
8HpW4kA5dECDT1IVhNhj1ODmEYFf2iihDuxWYjK3Yuty405nitQGKAlPmZPiRbmM
fE4SFzf9zvQO+/8ZsUty/SqOAJWnJneE0RSqtixogCPP9xj1sm/vnLYcpVfgG5Z4
CgH0Qvxgpg2UwH+w6uHlgeFLIE7nWpiu23cMIBH7nj9AWxp65fdKZ+PHHXIv+swK
EipD7oMN6s45uvtSiVLbpssw7q7ajKGdnpcoCzadIYK7TN1PqJC3+PVFHqwssRVE
UPxgooCGr37sTDFwG+rhbV5hXxfFYkBNqxDzMjjf5k/gGgOfD65+kznnxQWRIQNq
SXqlplDAceoVpBicrA17/2ZIiY4gOGlIj2O+gFkhZXckMuLuNbTaC8YM6PHJeXJ6
YB/vXKGIdffQvbYWDVxEKjdVt3kBe8yxFjXt5q7Joloqgx63qzsaPXPQiLF6s9A5
dVglCH3MpQLL39X+UJPrRIfYCsrsqObJCxpXko3V6EpPkglQ8EegYCJAiGpYrFP9
LkNAQT5b48CQt/39lJRudB++IM+gCJR3QT1Ic0SeKQcWCR/3m/Q64TmXjDvTavcw
l6ZWuacjlqHgBcKoo21RgZvtW2DNG9PQJbLB1d7eVD1awFeQcKBjxLLMN3qFtxia
6PUzyCNFkjOXRlbXcBSoanTGMNsThLmpPLP9Bk4/q6jTjuCHOn4rvY6hi+Pdr9Fp
QRD1sqNVHErbFm5t/VVhqlxOWBeG/jhpEUnEBbPmQ5HTSCyIvIn0ycKyGZnD0JmB
/Zsjij7oPhCVDfivzpXCvnIinbb0/k/poMir4XOmuD1JLI/Hl/3e7AFxyI4ze/m/
ozfuhJZkLgFKur2psoeDuVobM3iXrNPCUm74tCjOr3SXz2IYpLHSxDBARcN7lVRY
L2M6PFeDxO+UR7nMLg7tZbePqHDFFO5aaOrcfMgDiWGDOD8Vsi5M7Vh0ysVwU626
H6KEJY5Izrkiplk+LtsOszCPPpplnXjN8dxqTfCOzrwT0ANQDAd3JYGztmqSZuNN
aaZJ8yejAvaGUvuelsxSRkCc5vrrfaMV+MBMHpr5Y8j9AG2IdPJH0iicyiPh6BVr
iaNYYc5jq3Ls9QY4OijPNJy70OrA1wwfG0CLGnuAXoLujSTMi3mnrJw6q28FkHjK
3X0tt3Z0Jo5I/kzq3tx5J+7BCU0J2Wuq29CvZJLMKb7el88JybgUCE5JVUx7lfBz
HSvZ+nKXgu6htVhWKdljJkcXYf9yMRex9pH1idl1v3WjW+At4kYfNO86SblA2L37
SQNzHD7vYZsQCCGBgxUT9u0hP808GaSzIGSqGw3116ZChowiWw5H0thTB/vcDCu8
GaTx0gse45v4srNmHhB44jwqrjQqXZmQ5S6CXuxlLqtoNdCK8whCdf5dwgCkPnVJ
JfnM4UZjS3xOwhxSzc/S5iLMij0xqh76wMjudQoGUp1IzDTdftMafd6WL5kZwDHF
go89yFHH/BGrIjGTcSF3S2qD7bu691TsAopBzMvYNudU5zpepqdGKT121zuTQAxV
EiHPzszVtgirgAEGFZBcDX+5iMSB6p3qTHZjraIKOK4kZX6du87Xr797xYYcAq8L
mO3IIyEb5HfR1VYddQlhZ7Z33sA4aJlPw1Xi+GqtxQJjccu3fKUaUYGJ59s6VAPq
9ZlRmK1BELAI2fDHQqe7hHBJS7RYBn9vYOP2f9N2Z4MNRTIyjQjQcLA6kPzQwcbs
LTIWzr5QlJmtaKzt6zJY5BIYg4PcffKeghHyJ20p3Q7LRYAWfgm6KuWTe4akegPB
wo7K3EFHVbtJfJCYQTWyDondk0iWlfKssdKqlbrOLeiHYB8/Zu3h4ky3vKjNZd8V
0Yd+Ph76cf2JU1qLutJzKIlYpcv9kGEe8Xdn4eU6VYGC9UWaK75hLoE6+jUZ7y47
sXinb5L6NBtvgwnyYSB+0BpGZEsSnpnOgZhNgmGdl0dselTPG7U4//iopBgyecaj
uwUI+QR89DM+Wsf3dV9vHUu5aYxjlfNDz2IsllfdcREEo4n0+boIBqR+9fg9wwWN
c6rpfjLPdXT1HF37hAZe+5mzsZUC9JLAgnCYBaaYSz9B692yAvm6FlgU6fwFxmXo
2/CA4Jb0/G6zXbrov2t6LfJlFCpUZmxQOnjT2t1pRfMilRNQJCme2WcIEeimUHiQ
qMD4ZnZZN+cdog4Nw7ACqALhsZH+2Oi+tC2isnid0FQeXWO0w5xT6iLUVFuU+5fQ
x1hiNUxRtq5+f/WJMCLzMNw4CRwDwQPDWEnC2N0YiSrTTfCzkscBCdPQpLflwbPL
PkP1K7wlRGLmmJNhngajqnuS/EGiwnaJthFQg/bY+20oFOrkElgKlm8laWxs2d4k
cd7wF4Rq+QIsf29lubZED5tMpLaGsA3vn/qt0HcwX2oaLFw5JM98dnetnXywjKrC
3S8sdQlqjV8vPDnItm6cTBTSMZ6rhkFqBgHvVrClyiQdrWSmQeE0PXhvyJOI1u3O
gb+co+4UKwulQhT1qlxt5J0WpSuCtpdAXy6i6dsBnrpF/6ivpblGDQdZjwONRJrH
DtrMFuGF8I6Gv37zkoeYhzN14Vhiu/l+qsAUfX0kK4WffiIY4NAIJIKGu2IB9BNn
m8fuz7s89vCjdgR/ybGq9SqwQiXDJwKgalUJ94YdCC9E3ymHXA+Semy1a9wTJTvW
wjBzQw1RPvKLEqS2+vlP73cTIUnsMq0CMoo3x8ARrnppoXJJKT/+YQKfAbYGuBDU
183A6e71/gcvR26j6EXiFZJ/EkpcDavL1aezzNZdukX17ovZTrCTnBg2CenfhHIA
kL8zmX2LfIP6AtV6lAxoo9PTdrwTDMDKeXKTE+2BGSS8WQsRgVs/6hE9qaBI714N
g3trLHeG4YohDdZmxSI/S7zlikxHbWVmIf0UPTtUNzKtcRk/y1UcQjEERxnEtv7f
Tl/y6EsYyf742FNMZcfMCcM7xslwc/j4qla4ce2pRYE9P5AOnP+BFDGFQy8C75Af
y3vew91LxZQe8uY+IQ68T2fTJ8lhinc2RYhIxLRs6eCgYGolS02oDcKJGdn4gUxm
AQ265hJY3wT+syUASojWdInAloIIim4UqhuQBvQwV3wPFUgKVpX3SYYV6nX3nD5a
GsJjRIUUic5S7C35luyGvIIIpLq6jCE/uiRWIINcLKgrly7rrbTJgh+tcgeE4e+j
XwaPYwUv//2S4wcEJ3EUd7IJb4XQSoiUavUG4OOD3qBhJWvRWkOJJccdxCeoQ7qd
4Kkc+zq1x2fG6MRSReAiqRMMNPF9uyyxIl2Z3G1zZEQnkWa6da43vk/jsZDdEXzd
lc25kiwCUgAa06AnblT4QP3gDLPmTloY77RejDvZ9LLNfVYMZwinNeX1xii1iJCi
A2C6z+KNBgZIGqVv3Ui8oCSVhd7YBmads0Yn6YZhDbhQ4mEGNQujZum3Jif62KJ0
0cdncVjRLEOmGAtwqFV5vEBgpVOwOc3rTXGaJfI4SOr4m2scd54vOBhpO3WlgrpO
I+BsA7HBo1Za4woc/e66AHmvl4rnfQQu/uJS+jxbra0h8KjzskAJudF0pfNiZpoc
V1F3rVTMBdbUq+qQy+xkWAjfK8Grwd+Va2BnQ8/drrF1NAPXRb90v7ShvoOsrcs+
izFIUXl1rRBRxwdCmE3QEZ7LQQtncDgZb0hoCc8ZFnNidkgm+4+4nO6H7cP5K5d6
CuANiw9oWbx9uaFkAkauu1Iq9onJk2cNk8aivm4JwEn7VX/y2jIiGN+XwiJ9uH4W
uGeZ0f4tzyuE+FZein2lSrLxl9tAr3FEmcZwCQV5SVcmMEEGY+NXrzKgCEDQV8EV
blm9tdgIBeW1kMpOBPWhxnz/JaqqX1LHrA+gDH/zAQ8FPgecV8iVtIt1OpjHV+IZ
nAIO7o1EHV6dnWk3utR1js3Z5DIQUIKH5yvNlKNMtKkX6R9dCDY39Kp7aMvJIcLK
tQM/jZoS46ALAUf/WA+9qSVLXwFtYk4U9C9epDcBahUz0ThBEI7yWe9fYGmhbj0T
sdkB7Ta/Ts9d3gHJviV+b3TcfSP8fNJGxU/xsQlND6ED23xNc0ztFEKE4yINSi03
z5Hm8seCs5SaISRckizsKEfbQn2Q+qRcF0W6Kc4sLB0qY7JFG9HmsBz4VCKobvF2
OcNohUH/arrJJUZ29C7lrPZDB897C+lam8b5f3FqN9WCa5w0Oc+X3JrOYKWtUk/b
GNKsomRVSb7vAjdyqXSAOdY5Nrqeh54qr3MmOQY0SVF9CO7enmmb2pmUz4ePSSR5
ZIeSoDfhWLr1iyW5TFjR20Lg1BBgdllE0E161FiqJ6Br9IsEoCiOnMu3zmPcftyD
EeC4Ihf0h6IsmfyCkPgzj6aksexNTYlTuc5czoANZ+HzglRwA7lsbhpegTSu+4Kj
rp1VutaXSPCW/yOqY8JVr7IP0xtyh0LV1sESDPvgLuw33H2D4IXs71OBK0LnbeyG
AV5myk/mpFq9XfBjSn96s54LZA58r4pWhtUiiD6E5OFabMbec0WGednz4zTpGHEZ
jf93N4/CsJ73l8LW69iw7pthAlpdomh7Jpryz8B0lWgIrB5T9SWxleR0vrgw5ON4
fsYWDNiR8x6ByxNGIVDp5V7zsi4D8H3UiIR2dQMuWe9rBp33UeJYFrEt1HLSoCEg
gaR8QsaYyztzlZ/J7K9hjfjmeRa+SE+Q6Uf6y6eiparbe4M/Jl/PnGhQXkIm6TPj
oJHeS+HQFRCK8H5SQti6YVGBG22W0WtPdYFteRO7HFQ2jzLLDQX5SN2w6AMYqJRg
OAMT1DcGZPO3v8r0X/cVzYFwZDUY9Kd0QNouWJFQda3E3gZfWway3xItixl9LT91
zN7ZnRj1DktVVAxjjiUNbeYkzLVmksBeXmQL7xnQ9k8ffndXf58d903fQNcTcjQP
pveMYSbV45tNZ4X0KSVFj8uSB9/p5cZM9dpYa6rNicP27j7ijMjrgbt+6iVqwA3o
X+FuDYrDbkiJtvF2y7SmDKeiwxTE2ptR10GHho53Ny7ab1m+6nsrq0aJhDAHOR9m
H5+VISzLhhZDBczrd4Z4QqiwAcoQv4dVk4kGqlPgO8Y7Fme7zix8qTDr2s7i8qJc
JnM2I58T5SqqfPeQPiqP2j422nGMs/WJgTBfSm7ASc1/1O4lpK/QP1w2JTvaCdwJ
QXFP42XoyvcxsHR2H84lPScJS/+WfidcPWwSkriS4iX4+aw3ioUwavnLTrk41y9Z
zi4O7vqdysJupIjQy0Q2R+dnOKIrnv+eGuIfbRyET5Oj2X+NXhNtPvgIPcuUZlZI
fuohb6o+8+hRi6fwYGJua7tZ0dU3xrsnBDYe+T+h0JKpz6vR6pYqBYuFNtAXdD36
5p6w98I6bzc3GhrqFRko86Pwr3evGETCnA44huWCW78CEUPanQ3TYxaKPTSfOEqZ
IQnNbI+hAJjSWasveGpNn9ktgksrG+MXaoq2qX0dmZr2KM2tK9ApqtvccBTj44/6
7cnYA5c07uhYXh7rwTfbCo8BGDU8u0nViXo1tYOqCy4eYLwbc6+pNW0fbL+rD7ns
uL+jYBWvXaL96i2kYQ0aItPpesEDfPu+pdQmkIMojwQA5X3SzEZTFjKsd9TJ/RfX
dBNDhp+psd7Xk5Pvxzzrz64AjSxfuliYN9ZakWdCHyVb4wr8YV26LSTNKCV0jqE4
aEAIE0Cl08JdhKf57YCDCWj8bWC9lf9hFBtF0auwSDurcd4OXB62nXeg7+04hkoP
0ySRCDpdwtHIEX1jahB190DTxgvDT2w2gDe6N2To0h5ogmmLZxNjo4CCMnq2xTFx
Bihd0A+SYfiPjYxCvKgf9bNiSu5DkTKYW2mMyk9V8xsz0TgLVf5y5H7cU4hMxqdB
T3ubiCoJvQiIVXHRNnWjY8V0Msn6nAAU4UPyp8vNch0oZsriVnmg3nHrI0DwCvKU
gCH8pHlOF5DmsjicGKhxkuVTpjYUJdeuUj21Fu2DYwVF2qcvYzM2L89yB4uqr10Y
EOikmxQFhkxfVE/RxV7aJgEga+uSbnol1p4Cu8E9zlaKMN4eKEZ/1/Q5O579SsW1
iSC/ZW/kCFp89nWUxsEAh1djG8TwT+wPqhyiyvtR3HaQ+IXeommlVvmahbV1OXy6
6JKk2UMy6LgiY02r+22+tVXYCoTKZZwp695X8IToe5yPCtN+BQoVG4CpNdafiC4R
THD3elM6utvXlwhZEQL+NQEQa6zNip4L2wBW7/ZqSCOpehnZviNOJ4ERdIcCHm3w
+El8DqC1jPMbJ7hlLUc2D8VAL+FKI0LFYwla5ZUjygV3QtZbxP1emi3zLlFtqeGe
jEMiv38p+0urXkTR0vI5qlY3tI7ZxRmg2SYNOjq/9f8M3g/HhvOzu9xegAOXF+UV
rc0O2b5OCNlf68Ns367xQA1mkojno7D1vpvFCUoemY2/ba3gwdba3u5wWT2N6gPI
pQcEPmAibx+I71C+LlbJvPtLf6ChrbnC5dalOu7fBJmYlwCbzGtWN6wninxjfUE9
NV2DbA8j3z+MLI5smfOk/EbiD/M5J3ZqjMCw6Akw+6jG6Gm56M9P4tq6Rpr5aO9h
ml5n8o1qWAZyiiGsd7HiERFvvn16OiYfI5gxhuLKrYidDmFike8HkrW1M8gbHvni
l09Jl+FOu/Xs2CF8tbebPC7O1J0SpjD1FePsO7NDOYuFmGE3HnERtMyQqJww5fa6
4PtsARXw4s4XnftJ861afeCb48A/hi/SmUM8mZEjRk8laD0b6hsI9/tYYQdAusjq
qmCvescvSl5/O5g4JYg/QXz6HQKY+3yqye0cYCYPPxW4G4SKkXhkkwRK86BJKJkO
CyAXgoGy6K2EFL9unCWBAIAlfWm8Eegsp42kj3cNgeyloCXhyDEtWsuJYSEV2n/8
hXW84PU5hhGBlWDPWFvJJXVi+lw7alDcKR+atimD0tcLY9ty8zmHVM6ySHrLLVGe
cr3AWlGn0mTuHazTKwl7AQUrEFCSitULq7+21ieUBWf2HLZcQJs4mnWDG3j5Atm+
8f+ZtEuV9caPNq5vhtEkLDzZ11SNU5oaRZqq4Og3HgPWdvowUD1vKNNafFv5RazM
DmDIboQU0bz74zX9mmvnzqPnk6SHSLfPp8Dq6pyDAl/UugtQy9qaRcUHkSvjxvrB
TpT65KKykTUjRtGyHwaEXJRcMrETKSPcJWbYAN9Ym7+RLU1v6viXKlrOYhBFvGIf
xPnk8HZ+IctZt7yWLkpQF4729R/Q+Tq64m2TP4nMpWz4cTOTkKAnxGe6NmLtSuPF
tZZ40lUbUx1c92taVNz6Tl3DXmh1I6Wjsd+Ttu49FXYlXtN13CZ5T7Tqhz5tKnTu
Cl6WHsQoRuiindUPNXOH1CC7KCXFFdZaCxRfku4voy5FVZc4qdH6owHEptsYJuMW
XVWs50P+QjFv2Bp8MlXoeoBs5MH1iT/gWR/2/CDxXBw3Y/XeYn/9+wbWeALdfAKc
kAKUxRGHzIJyX7qiwidyUH06wBzPdTdQjyKcp9HMK3IcHt2N/ST5tPYuACp+ca3f
eZ1bqPRhEYM1W8l4w2QFkAPjgNPEMNPUMpols2UN3KljKma4qo0EaEGl6fn2ZJte
PxKdFYgw27/9FEFLGv9qQMIgWGSGlyyPxeYxH1rKL6FATLmV3Lf7piSqSU/hDBp5
cZ0ZuMgUaP4n2pZcZykyKxsBQL4kDiSXq2hqJx7+z3QT1AlwL3I5V9hJDn22qamg
sc6YdmZlGLNY+1K69/oeRyFsXA2JA3jD0qiL1A1C6R6ZRXKppMF8kVq+SCeZtNNU
9MdMoPuhhXtxwFTq9oCj6osZ6UP2i7upbLH6KKc3p66ZjJNT9Ed29UqwC0wXguRe
52ylgJEd+bt31eL2p0cSpnmV/5aklrJv7GARlZ3mMlCV3zOIY9557BxKz1QmsW6u
0OjGkJqn5u8/6w0CDYzBkByJfoHQ5lSQ7TvWF2kubMlyWDVS074/FlEWFWBjLC1n
CLDavtjc/a16Fk23/qzCHyCUHkrc33b4MIKl3yqC6H5ugdz+YbzGENYmNbbQXAMF
6NSPeKNsFJ2BCxavXaI7NUIVNHYDyY/vdk10VLvUfSEddRI0eN0HdjCNh6u1nDAn
Y3B2Ky2RQB4nO/dAQVUgfljZdPTOaq7KpKAImKwy75T9wQwVy1+uP4jfnIBwawst
MocMIczIGa/ErJSIyiyJ3unhSzUsL9G9s8UzAxlAh+cHdlwTpvqGf5d1lj2Of6RQ
FhTgUJF4S7L5ifyBZ64r3DZfuHED1KH2eGTh/jGA2CTsYalfEMVZj72Q3VJIm5O2
t4yyqckEICKztLcyQGVv1Lx8/l3gnHuhma8fGRrGzou+kGnDG1+EXTQqEhdYl11H
A9BeF7ZwW5qQ/NNKcaI1BVJd8mncoOrAIv/XtvajiY3YjoiMJms38QqQdkF8SwJZ
uwZJqOJNTHvLMcic0+KwI/yq5Ei5aUOhANfv8BaqznIZM2G/Bo0Z1GbnMk0XReAg
99mE4KzBIDx5bZikyTja5wJkWQtXnLs+YjZYA99RdUvh29xIXQ57nKMfm52DfuDo
xpelVmgp5vOfZRAnmst/po4TUuzWqlIKYqdBWSb6ggRiWhpFy+1Qq3A9pkrleeci
aaNvP+X1Qy/Y3LdV5B8BMTZjhF9xcHSFah2hbnwWoZK3Sfz4taHOcaOzsqLXuaO2
ggklcz29RvHgT+QwN7d5PPqL92iN+iPvsigZ4ewLv0Ec2ZCICaWiNbRa4HaXNB4M
aeaWG2uTmC94GWrknxDCeYrWU7W8/y04zB7IITD48cLsX9mG94S1CujM4uLcZbNn
WyhfViAajGp+DPrhaALeWmJRLA/4rRt4UVkQ/wwa/DMuVvRdtP/nAzJZt0QI5C+M
aBJy0ae8Bv+jRhF13fD18E9HTmW5fktPJth45l2WmZQJonNvc9/5SQ8HtYpLMFl4
MSHVuAN24FHKIKyIydL40frvTxOATSg3gfrcLVOlARvjsxLlKrNlnjwMiaVFRm7M
LP21ZIEMcTrpco+RJxg9eMv05QyP1xLopxGhWVKe0YCY6QxrYt0BfecHI9OgWnU1
Clw+YEO0tdslcbYnhXHoz0pfOZFblZnQJQNWpAFXC8kLBx9yzXX/3xB1e8e/me3T
WIfvqtKb+YL0bqQHaicrK20e90s+ITJ8ajfT/O/V68TVC7oYUSI9v/oHtMJVWQQv
YXSAREUIQw0CryxZR31WHU4pFrJ64yCvgUapO6QdJdmG0bwOnsdyf+ir+2sdGzkD
j8//kD6hCH8R2k33yb6uP8DwKR1zGq2a0tZOYmDnDoLWGW6XxDtYCiK3jRyUF5EG
+Peu/oUpo10eyN5RhOiCLAGHhliqr22YRfLurM+3xjEqyKk7tq5abEHCrcUytSgk
UC7SHRvd9qf9EqJx3awQ65I7hGAnGG4OIkPmaJslisVmwYlLqvNIRy0NI9I4crl0
DtoqTMMZxVysHob5mPPDNaS63YAE2yXkp1A2JVO1EUXckciVWOQvZsje02IQwllQ
28oh+oczkVm90DQ80hV2Ttfwq3znzvaRSSuStock2KEf/+/Im8IVvM4OKhTWBxRn
m7CmbeeYy7dNC2Sz+Hjz9dk4UA2DFCZ3mPsloyvCn5JHXitYYuGWWY5Uvg1gTGnf
nNNRdudC+eBVJcJPvcfc5X90tcw6ODAAoPkMxhXWiaw3qK+ysv4r00MOScU7XC4o
TKwCC/93WCJtI18OROD4cfJewd7/2fkIOWrRh1HJpoda+vRoiPBeJ2z78qXHewtm
tcw7co9REuEc29CKV3vgGetVmmQROp2VWDRyLInKYF7yReE+BloCZ44hTlGblf3D
kqnR/Yt+Q2+a+4hHeYdabotrOGs8fExBvW81Qj132xPU+BVhbNy73OqiouOVE42/
D52kzG4fPSHqX8Nc/szYgUZCWo4/5tmD5q+RzQ/sQdMcwz+WybwP+dpjv/tgWhZl
gg99WEp0PALcEFRBUso7kqAqy9I6hA2/z5gWqRux8tVOOw+6f0lVM8qcyQvxNI0V
RDSFQC1T3nWdo2wEQ/vIvJRgSjtGUmJ/W0SRfraJ65Wsb9ZjAF7JAg+AMq6gzj4o
G8oxoo2Hyj9n+fN4HAI/Xu5FNqr+xACcjs7nTUF/a16zMefwguk1zcgS6mDnzXoi
RZBEhiEkfgiTSaTIU0Lx+wRuFd1Jvl33uysn+jR0i/BOmeb7mIfP27GIiY83VZ7k
yKAcsfZUsu4pvy6HyivXtjc83sCBHc7aPOGyskTXW+V6no7gwom/DBMFkhnDmE8I
OuwMueFUJqc7cJfroCD0OrQNc6Z8X9cBwjHDmI7W1HxU2bRD5GYyEo8ErWn1LHIi
WcnCtoE740//GyEjsxA8SC0Rt4sN1uFZrrPgrFlsV1yAOcQ4qksHO8JHa3KS31VY
fHR2UxqWnPMrOVPWztf1IOU3jI12HN667u1V+93jvBTUK1ZQEz9fQSrrC3ZH7RaK
vumdKjuhz/g26cCuTg3d5iHpPpNv+twy3iPrE49/A4LVGEZ8FFzfydw+E8YyjnWS
G7EvDrHKHudUvi8ctoeieRp00EMtCInPixr/2JFIdv85ntPCx2IFL+QLu3jGWPFb
z5PlE7yZ8YhkYq0oLyH+laGGCVDX0H0kD1IXEXUIx5uEfGOcSAar8yM2vU3E2vy3
hewn6RG+1XLWq8+iBMz6qQ+0/dZ3u9eSPGPcSZhoAp3+JxFhvLZVB2EX1YR6nx68
SwPhoJjl28hwYm32uYJT8EbCImYee0jpZTrpbq++ZE8GC4ilVBgokJbCLxYzFK9k
mEpcEUV9ceMzg9vgWzKrON997veIX5P8V49OwC64egtkB4fnOdy+WtQj2s8bSRzM
XskOIuYXWkP87O2kPk71J5gs3e+8iqOCPptMo5AQux7Av+2Nryx7gVs0cnk5EV+Y
EE403QNnmrKrCqqxlj92wTg1T5lD4VkMdXm9cWgYngg53c14iCdEwsf7SIsZni0h
NO8laP5Jc4ZULLz4OsC5SeSjVFPnlG8y7O89ltYVJEcMHkojxIepfoLRoEIOEG6y
9mL8+ONfFUBBUEfu/77VYIJedp9u9HxS59tzckhIoHdVFtatXKmyUmqy9lwgya+2
37R82Gr1s4X9jDk8ygbSZY8Lo4tOpdtvRM0456im6Z6SC94Sb6PYmLA983vmD1H0
sV+4cjPIwvc+XAs+HwPizGNOEwg+qEJIt43WLgqQKJf9vT7nhNq4Idp1gYK8c4nu
yTQOT0jTdOCANoa53dLR86Ws4Ewm8naiuYDrfsIE1ukrX6af16KUM25pGgBwNIUU
Ew02rJ5DM8uXx0HXNTqFz/6sWJ5UR/iyOMuJnxx7JoVKCzcZ0h3el0hsJIZbn9MG
l37uhxReCU/0/2hKWLY9yKj9wrwMzFQsO+ybd+WdStyKyaLivT0dc2dfBpS7lSnM
VR4b4K73u/S+NKj0fHWWLdCpPU3fXvvTHUqXf5Ot9KjQc+9coVrqzoDbAGcPWR5f
Vx9uF/NG9/78wWrTEIG/oDejvoualMwKutKvopVVUcsZNuvEXfmbhTrmtAaA5B3V
LDPTz+jz2Rxb2z5XpkNvRK1CqnT1Mf9SNEbnh48qRLcZ51UnYBzuqTXozTb90tNa
y0bcAPHbvDbFdg2uOLSf6fuFt0gDYAEtF+wXDTA8qANrKbVPASqqOmTeP8oQFrmz
5zGzREzBvvy5Z0ElAjmj1MOoTFB2v1kRyFwXkRjBjtS2QobW/1kojisl1tmfEbln
pQ7F9vWAKkQDUzbbS1GlAgCPh9OlkljZ7pVaTZDHNfYcMhER0yFPLdISl4R2FXGH
J6AV9m4gHCvSsdfsM1QobLL7+9/6dtsHU4QEOzcMIUWi1yBMUqT+t1pQsnbZf9iE
3cScsRA+lPwNf6Hmx/cH6aECB6y5YpsBnQFQtGjg2mFw2iOXOUvqF+3evUFIPmMd
e74EXz1+D8FpUgwE4uoKuxa4itoy4ECiD3emPJ/jTD4uG5dZmJXD4dlz5rBtjZK5
b9MyHKZc49BoywjXdKbvDT2IU+czGNqu3SGzDN80xT/4leMxUGHCtTU2s5X4CFeW
Zn/Qfg6u4/pF5B0hbG3khOMSrtnljnqkpWMYznZqJhbZqzBm68U0uq2dA3i0iCRD
VBnDqDmaKQdwAlJOYX1pOYBaujS1qzXUWXJABGjTYncoUX28tlodpaL7KAqaT9BY
G94DRNZFeGGaevYSyZPad+rGbZPdNzMgLJkcqKGzGSM2ZhSc1I6sdY1S2gh5YVN9
naBsOEfBUTq1i+f756YhcjdUbpwdbOJUTsrOciDuXjcY4EOaD1DuZCkxomedDolg
fd49icLfN/cE+SD821M/ZVK2DXdodkPQcKzFNeuQb6BghSheDIJ1uHj/+sWToGRk
HvuiRoVl7uP6wxE7JjkhKmIOpx5u2PyKB8aj4GC85i6qzyJkLQLfR3XMjzcBB4uN
bzQlxfy1ibxtoe4spq511B3NtEBa/tI7nkVYRRxHG6U6yQJ9P5+9UW5hj0Nr4cWi
w6YR0qkE8ltwYsuIqg2LVPGRtF0uQmIVR1xkyyhA4gRRBu3Pf8YfwZhLgqltlts6
im9n+jHQWh1It2Hn2SO9obrVgVqHCEtzoaeec5ahJYoM6nK2QN9AMg47Ec6v/ack
HyR+zau0UvszjVEehuZ2ga1mFbwOZiFOr2hzGvCbkp8qMC7XY5eRwnTRHD+WKs71
a7t4t3IMhgAkyxhUT5i1UnTgLnBMj3ywNviQVI+gQFfQ8IRlwB1QyagZ4b+I2J0T
3y7fIXQ64Suzs5FY04EjeFPhqI5RVQyHl/iT/fdEq5AezeQRh25r2x6nwVvwbsvD
oY24Ft8xgWu9Gkit6UrE3F0c0W6FIrECnDkru9B7/+fhUyUEt3t46N0gTn+MEY2u
4bVZ/ql+/di7glN62uhUZd+sx/r5zL3A9He2cu27BwzC0lVtfY7jvSYuQ3wq3u/x
lbrVheMLJxouEbIIaWXez/FU4nN1blmfqtXKS8fZJSDGQbmrsqZAPfS7JCbGOEWL
JgoF+4rVS0LvkSHJF7ELa8OuqhmtrYpKJcMtoAkPBtn+KILFLpoKsBrSOY/IoAO7
cQydhjvi3lQLeOMyWR2UPzBK9E/VQrIn1RClGp8Pu69VFoqGvH2bBKQYKVWRqG+P
MsLQ3nnT8RoUAZZTfrh7Hr7I6uS06W+rxT25Ljyu4GtMvQ+gsYgfJjA3d95d3ikF
dtbnACrdgasylvEt8rjFh/TWr/G+VG0ZODSdHHB3BzXSB7mQzLkvGJFGj0FEWLvD
qSfc5Wd6qQ2VySywKIs/DrJhp49m54cpVfh53ie7bvoG4LHxGuXgS+/iFYK4j/qX
eaOC07q+981l9GE9hHzA1vyqxeFpZVPybEmqkMZ5HWohdizGH2YToCwYY7ovm5/t
pc3oIpeWvBdmnf9H0TdlQdHdHLEh3QTKqmrDXKwtbJRE+U/7ICy6crVtvaA7UuYB
4B/lg+wTwxGTcXZG+JeI5pnP6QCqjMu+6YhGgYlEgXOGS6syihEs0NCoqjPplLPN
Rds9ixPwl7T4Af1FyN3guv6Aow23DyMGgGqdmkHLgCQW5XGtbkjeJ7Q/8fXX/cWt
ya5rWsStHb8ZyR2h+hqWznnSmBK6k1ZTruAolEsAEmBNKmnvlKmpwfiXeVpzMtlc
sRI29kNb3znSkx0rynHfuHeGhRWe3vGdb9zFtjwBooJvqZer6gZK/kVVCTfngI9R
yuGhHrm73nvgqZnvWJ/QV4SxyulT1AtiLd8DxWqtHn+0aWXh93O1WXnlRP9NCkkn
FeLeGrtXkBYPP8qsI61k19+cdZZSiQQEQqb9vLKRzkm2kYmC/o025cIByni6X7In
KF4Ace6Vwo7u9pduD1if0U4uLoulFl/9rd4tR80OJUtz6CJbEjrXU8eyNF76JtDj
dZAhsL/S7DY+9cvMjzQWwTgtHBpCqeACy4VfwRSih7FzJax28tEt1XDsN8gUOtdW
DdEWnXgCfzTpEVuapQRwk6usXsUhj6hBmR1ucrvmMvZclP4TjiSdaKF3AmdbM+f+
efp5vNWKebNlE+qIZ5uxY3DPxZbIK5rSSvF3556QDPt/EVgxkhuFhd9OaOT4+1da
gXPChFU3VAZv0HQBCz59BNyT+7wDYSRo2YmjARhwRifxJnpeD/7yOMl6qdhtv0Fl
sggene3FWxQIjH4Gd/keSbw0pCF+TZrjHUkd/5FYR9zm5nLxmhbT3+/1CTa4EtUy
CKLCkRECySJzMUaEWXqw+SxBg5OxAhoxpuZ4s+F1VWoeDtha/TvomJUw5Hix1/RT
0Quun8C3yWcGhA7QDW6xdJclOUX1/ZvfzoIRYDlXmdbNRy6pNauFT6NYGqzynZ62
iksHiV+9i/r2Ay1+oTvmZXsGpZn2rAvTxLujiUqDf7QYLqnYR59FzGr5U6yDoZya
drOL4ZZE/bTChiXUruKs+dqDWLZTj6ap/6GuaalulO9Cqj5Dx6rHD0/XGXnuyNb+
ZnmsSWC4nr7iyWuskMy3Qf0TAwb4Lgtgt0W8bOfaBeRUIYPTu/XVsrWbMb+DxhnS
ztg9qN2Cf5+z3uHzwh1zghHHoksm1LuACtCFJzKxonBZZ1GK30mwGk8FqvN9hX+y
mjOzrnqUPajH6jHpEnvlvJOQcIs1UdlpFE+qXD/6JmfJ+iAuxREtRkYAjUKt2pcZ
qVqbUn3yVltfnHP5y1wC0kXtg81qxp6tSWgLAMo1m6S8zDFIKgq2yPMpnl0G9M0p
Tsu3aq5PmQfZwxIoqxK/r41zPE6D3BHPCWvQ1LSPyqyUzZbqmSbqed9mYlMdRb00
EFAUgq5NLR74zJ00MlRi5rQ0U3QmS/g+a3+ar9Et0yMpedHhoXmbrURfF5T0MfLG
q0zP9Rzb8GZ0mOWyn+hgnYn4+ht7NfvKYLfUuCE3N11RAx7veHzvNa5eBRwEkb8w
MMwoCyy3cVVycEmibu+d4XvhCIrD+3ChKwzJCX+JMBNV9Xu7lV6stT7B34Wwf/cR
CXzomTQBpYBxcu1UtEGw8eA/A8VINU6O8nTurMof6Fn+1B7NTQbJmc/R3Z0wRlsk
05J8VdZyG8lj86VtKdP46Lfsuc42fUxCZ1kNJ+ukGjoVqtVqCpSKdUP2JXD8QFSQ
PtO7Hn/ig8bce7U0yaALVq0YgNGIBd5mDaei+DRpyZdpyT94HB1eEBw3ICsWck8X
V1c67uUTCWUBNCJf+dmEkUQRLyKqMv7uSQ2wIkUue1Tj2BLEhvk1w/cMAdixL8go
A6gl200fCekS1l3GzFklh1gKuF/caZ+p+AbOLN/XNxjJu8hErrkwIVVlgihpJpfK
cnTxozGZMadGUknjzltVtx+CAHqE3sVQyZieHTyTREbx9/4ODARYYmz0Ok13pr6+
UZBSnV0dTdhdR7/urC84eQh1PmwpO4WYbPJCOLx/+YprEUhD3zJ/2uvNaPQyGBRg
hxE87EWMwz2rdd5nsWWdZSCsGAJ7Uhb3SPwJNVel9LBh2ftFUqixtuMCdyJmazNK
zS3UACMjkJMi5Z0Nzrc6SMbGDcNhM4XHDkayBpxUfdW3+X5HhxBkcHeKOkSBrZM8
iEzq1avPsNRbSUZwtHC49xhpIOQ3JmilQDJx5mcySmrjtmmwMHCdW/FtRTqaj/fe
Pr9oG6h043qAblLSFE4PS3km/pvp2tmfE5ujopZDAfS4FhMhnxwoz+oa53X+SR3v
D/9Y+GR4PeUtbv4RjhIwetqJup0nlglxMCFFItbWCGZYbs5DwWYDZPgOxgs4PRH0
9esx4+5zdzyHIkcqCdv1TGjMNWC/R1+BKEU9VAP7gSEFIRJU7cYcno4ZjPQoC8sh
IPdANSe8kodX/b3qJKnb4bfPtRyhCPbMl+M71Qg1L7T4rMG1bFDs4gvnrHxpdZZI
YNuPI3TRU7rhB7bks+RVYAsmPFUUSkhd7mJq9TEhnMETS9NnhJLWE0FEIo+M4SCs
+5zBSdxVBtdteY6f6i1+/bqJddn4p5Uj3ULG6cBYlR2N42+h0wb9biH3YQ38xe/3
5cgixTmlUeCjUDUi8DX3QHdESx0GL+G4dDJgUxNtP01x4e7nFqIO3miIKdy15W+S
o7P1zSAQCSxTPSVtGW2cNW1SdZXCCr7ZilOxFB0W/FKfDm5f4r2BHmw5igltrA5Z
FHENF3UaJ5p2bmWrJEzPW0n78mURWjvdzh45sCRu9scvisIOWt9pwxBrtx301xjq
r1HTzzEW/qXfFU/+7/mA4CoxATq+DH4C1PXC7sQ3FWSW+QePGFq411eKDBGRHqhC
+6s07Mj+6ULHVwmM/j3sWvaUY3C/jj/CCQTHgCj/hykQag4jXIBdFH98RkiDcwlt
tP7/D3z/Dtkt7OsPYS/AK6l5Re0qBY4z7sbXdAdovNmRKpGTHFnnkXuEkKce+/DH
gOW2NWQvF2/+5Ved1IEAjHLzxE5tfxqUcZPt/FWkPLs8RraJuGOx1LIldvbRoz61
+ckUqlkMxMl7Y1APWCPgpjP25KxpNGluysXFN6LoPOUkawyQl63YqwxOqIhK3LsM
WDBgsQgCb3BRdW/+uwT1YS7bCIQ3Iw3S2B9KBI/XyRj1BcOaUsyL3iH7jEDs/UIT
Dat8KUb6bWpj5LWLwXDnnK4CDFypDbzBdWoChiUDtowU5y/svQ5l1Yp9mHaUJbQm
plxh3o0l1NGjqpYbk0AgPIL7lygEKqY5T3az4jajcENf6oDzpgHd+7Kcqc2aTSNK
IUElfCPoLoqXXRQjBLJ+YK+0amE0pwDY4MHVKMuwopcbkP6Vp9wdgHGtqBBZxQrq
CMj5xPy4Knnfpac9IeWS9r3TWzL4VDnF6G4SDNvqHGfHYR1PYrgsnT4wir7O0bPn
8EvzO4zbpzw+9oF0o+KKZzZfaK0HmFep/v30sDLjcZeL5KJ65Ro9w6eeqpMFDbcg
yVpHp/mPRzJQHq+PKNjdWAazAwNmVPVM2CTrkQdV/tVImRZz10LSMH6jwn+hosfL
mKJ8wvnaYaXhJTTa5XQIIzQItnQpX1v1v4OrIk7aC0FWpOnpJRjAc/ed23WTe1R/
rmvMcZnmkyLtUvemMS4xustr52S1k+nz+Buct9smuv6ysO7Gzf8iNovCHHCCbNeD
v8JHD7v3ljSfM0JtnQPbUpbzsxFCXAhWGmifTi6Fepb7JazgjDCUIqc455kE6HKg
5SmYSn8kx/k1tNMXr+OJ3bhzb6Qs1wMZj43rJTuPuFF+4hHeUfhR/WvO3kH8lyIs
/qb6k4STYFt3E1/q3n0/ijOujFPyuRflAwXsStM4Kj08Td9RA34EAvqwqaklxIhS
Yfj6KxGMeBvta4J+YLosPedtLtdJT8fMTYRhR9LSjl6y7HVF7iSs4l2jlEXh1NiE
nDc03OdGX1/VKsRkNGSyM7m+YgXe8xObbFctG3cPCivmVElUkncjT3N10RtVAC+f
jmPh5hUR5eHkxlrQiSR60zRNh/VupzMM20neCPVDXdifeSn4CgRVBUVGcSsdRNo+
bvFfSw94Sl3wVZVE3M8d6BwBI+El2aFdRCx9Yw62AdGkKvGqT8dsH8q1TtbqLYQk
FyTr4pA7muVB7MypAFusUmXS2IjPqrgjei5ej6ShtL+kCqMudy6DOUetEElA+qR/
TG2LoD2vnVD9HTfFAAZwHZrQ3e5ZvRu8gzBurQY2dvHD0Lbj3Ob3CGqYefhviP7b
014bfsOAmV7sWgKfNCWyjCTJRVo29avEl+BJKrTvQS4b92l1IPUlFyh8U6orTYon
mJ7PUrZhH8Y20dnhz8fuyIwKJLLgcS26PByyq3WRHgNC6++cyqdo6UpXRyzioX+W
xNP9AC2uoaD8HU0KNfr6FhNys8+z29/hvVnZUwps5K9OpfIpu+tMoGwr++1R3hl4
GHAfeW59GZHdYAyKyWW9gckvF+8qO3tz0QTwGVGm2xEB44bcFf7qN9siz4Jh7qoH
k+5/rCPae+Ti/HuqdOpy8KkzQcmht5LF+9d9KwymAwxapqI9mQO9alp2nNYtDxc8
MQ0aLJWNFA94skU1TgZ0CZCN08NvAxp4MMYFL3tmBfKVpMefzqKlxnmAYjAqd0OH
5THt6XdDOdCSMOrn7foYlbFskmK3A9bfDbKohdHKgELUgttAHmRkl9ic8DARUKuK
kFhqxkL1AeF643ay3puvg5MJefJjeQP6P4hrXtqgwzOV0+WEDmbHXhyTVXrMwXUp
VbCU+TeUZivt7fbzk9IrUmoNTmwPvJXw1t1SJpzR4sWCuX9G5SmZgsJOhtxxn3sa
AXUjF6rUmPHNhAXCgWxuV2QtfVbbeimM+b/uRuFJ46R05JOs9yiX654xLWcaq7fV
PRqWHLHqm9295mlB6NZPYEq+N9puXgDcBDxf9s4l+HZFrvnI/h0psr8aHxjqpb8X
4cMjjBN0TXG6ky7j9moLvywFLzLdo7mAcG0o97+sMWKk4MmRilxft56zkJefHgl9
b1MKjrszRlZ7/kM7sYGsIIT17dJAn+/+Lk8SFk/4gelvZ2PI1TGcbsrYIMf0mRAo
nUXW0W8RpxYZS+8kj9iUsAw+tP+PBKJgH5DRAiuWrdG58p9pzzsqpuKO4/mSncNZ
p2TjEn4R6DPa7yDUdyDJO6j374eO+av8SJu9hdcw/C4uEqo3u4IcYrE1DFjCwRD+
DV6ecJXhTDQT1lhFngKpBW4+HW7bbhOwRGZLG8rgMvrmt3nao/bPD+oOyCXYhXnK
IHkSUp80eHnMjHIDZnf/ygANHIdKyhYS3x5XwZrOAp2nQkVWantnZ9oGsfvvPC7O
2E0NPSIv3KuHaFN3yeydU/U6okBK/Wf64n4cHUfohW1DfoavtGvGK6gkORmVaZ4V
AM04liTTIpko1Ieegzm55o5xMzu+x8nNrS1fG3lXa7LJUGRsHWIar1FZ1B6lO9Io
iODTHkI9OwHE8moJ4OIlbhK87RPwe4ie1ifsKxWlRG79XBVnRdTSQ4F+NnAilgYF
/L0pQfe36CZeFPoyiXDrWOEJAl2S2oe2VO6IIsBwj6lE1/YU6ecGdQVEQaBxy0UH
W3MrjXrt4Lzy3jIZGyJ8T340M/uWnpCvqMRiPPsPV7u+PuDTWF1V3lu8RG+NRo1K
yCPp29/j+T7pcr6UcN9sQJsFZQw4HgwF00OIvhxUPGGbx5l9IeX0X5+CZo7Qob2V
BR5Hkwvp3hU4FMctDyGtK8OMYeh8Hl9s9JUJcWHHqRy8LYTBi4TaPUIL5KPExtw9
zn5pzCSev/ZlwcXYlqoRZw3jFjI4BPlxWGrsANhsABsS21j8PJoU5jWgdQ+ZguSQ
o9yvn1oinVYIMBxIL2WSNARC23cxzkEoXfgXjEveaChEN7+V+NvH2bqv1HKDfITS
bBBYn0oE3Ukd5AKAZWxxIREcLaf2+RFvkIAYJs+3WK/E0WH72qOZGqX2bqnZRPuO
AmyVhFxEBvmCWygm7Z4S7bblFMYEx37GZAatf8ZHur+hVd1LBlxdWf5NJfdkRSY7
ZWs6XiFVYhl9cErwN+3nhL6bVn6NWmHuzxlHWS3/lrBkLFBMdFh5FKGY86XGnqEi
W3YoyRWRYGHW37fvW8GSyoVLowntFnigkIwVMFBP7b8eMPJyQzqIMzcbAaAwPZ7d
R4gMRxx1+eK51e2bbHt4IgEmQcfS0Ez1nV9Nocnd0GqYyN6BbFRJ3h6njFyNWOwV
CqXCNB6ILk2XTai67i2ViNlUF9RCCX802YsbW53XuuCQyETUhqtDc9Wkx/xdm97Y
7ecE5lCG0hAJn01x26740zQ/sFz2Y1PQa2k8mMuqs6XRKL1IGPnoK/TKpRFHTFAP
m3qzBu8KwGECU0sRLSe6mixuw343VnsaZPMq7A3MuTbvuF5P3zN+MrftWtQkrLF5
TtP1j9PdAHKK/HaVT3AFPIlJms2Anl0L/bQAmL3bSEDAfk9IarruAqtB7q1myiOk
tAmj5XtZoTtkloMIv6bLffLU0Jkfm3H5IwbgMVzGU19/RFShykIMigNbk3y34Jie
fbIxDfWuTT5F/NYMtzy05xfG2z0TiWrF4Kt3o9W/KJR+Oq9maYZEkemCZhh2HfbY
OtSEEgxMNiJ72c3qvuAdimgWqygUhLwCzzaYamgK3Eg6SRFLdeNN1AZOo27MIW7+
oOE1m6ASXInwFTQuirHUP6MM8/Bd8djOcyX02x6w364f2tFmZOWxnFcaNTopmCdR
yGx0m4zmnM+qQ+wcTX2hLGcK0vZH4OIdZgNswOxHQqCIt5YPOri/3ROgbIk3DQF0
EQS5xDaMM2eQVrsei0WmaCYImPBZEokchmaEYFHMykDvGpAvg7azRe33Ntxkx2ym
/UWEN/A1+QPiYeC/JF2n05BYjX0X+qy/QWkp+jSn1R2bZDT7vAOVQu7qfCKgX16x
xIAzMmViqiZHjNCfbhrOGu2od0YFA78EYp35Hm4hphx5ofjx8noic3wJvNWFhjzF
pb/fxaS4P8XLlT5bTQv/Y0jvqhKxy/ruCstQ09tjS5ZRQfmih3WPYP24pdvscntB
C6ssY0BhbYTFFxWGVdEEO95jmX3NOmPrh1q4Lt0S13aLvkEA9nP/f/rOEKxrbSZ/
0RALSgjkOyG+OLg8r/nMajkSaNI7KgqToP+ayvlOeMm+KThNhHjivfLo5Yi2M7tq
ztkBehvBrCfz3zhmNKdhE95rVTIIF10Lb81TSMnVkhHumVnGGyhEABPmTVW0bTJI
NgJhnyiz8gZpdqa1SjT/7e7xyrUyQdbdfu4fjDTBGtkHowiroYG13be9pGu1PNCz
buaDw/MbM8b5Qs4IGmwUPrmzS4VyK/MUhs/KsH3iroiRILhwn+aMeHPnd8730jwz
2YIUK0rS/vUdW4fG/CAluw7tu/J27iQPiDZN5yiQxyc/p51dbxegMkZPCw2dnNHP
N+AQOA/ySap4KNdhIjKO8Yy8byW5PLfQ+s6nipegNODgJ+EDV7RgHuHUZxHrPxKc
OAajlsJDaNotzCmjCIL4mpgS80Lh97L0tld7TUfXgDUDkIPfBi/l0JskuYblRJf2
xrqzIoenQhfWhw2j/4PUdbTmes21dqTsdss3ABlo3VLPWgvkK8X4C0+me0rC3Ekh
BH/wMeowxuqCwTPWXc7ZDSnOLboV+hA0/IfMtDMeQT/XfF6fI/2BbrQ3jgRCBsno
zKoR2tr5DWMoGzYs342WqQ9oaFkh6GzdBEVRGy+iK8Y3H3gWiIu9ROeZ3tqoEgzr
n3KTdQTmaEFGJFQAdB86nMmoPp1VdtVMlm85lNl7mCLXF/GxUpQ9u2j2lhzBYg+3
GtuGrQuy+Fz1PWOmPRoIn7jKleJTZFMMgal2Dr43w1axXd2JayFi3O4OXUxfn5NU
SHJ9OAl8RFj2DmkhXPE6POLhb7qIjGZFb0QauRAaH7Yi1yu0k8FTV1JQmBtulp27
iqxy7AN52bAaHf0tkhxI9+3jscIb4kLFalDJScAqo6rMv0IttHy5Ljh1q+7LKDcN
+oCHzyrUKn7AYBGi1TNiP8IhjxgvBMZk2nmOptIqKrODWsRGKnDjWQRZgPwqwnuC
bkkXWr9ItPN6saPpaUeaK4bdgFP5TIAgm1i8mt5ZudPUdzoZhmJaurm4iYLx/wAl
lhnTAwrSVEBT6BI0sG70yT6o9nanh8RYUrKgP0YRzOP3ZxW/hCjOdxs/KKP86LAt
9EsdLIWm8MOPjhXAyjsPluqmeDHRvwXHvZvQwp2HLQpZ1gpPkNDolPogmqhoLNzk
nQXMsF57YWtMBPOC+VWWuanV5E9ZNVCJBvAXeA8Cm14Vpad8IuICE09zaf3vM+xS
0NMImVfYJALNuSooHqM6HEbuB/w0sozl4+cdPtAXkH+w1gePLo9GmwIAO4C/NJhw
ITWIbsoHysPgqj9Voj+KpvklXG2GxlRbpQ7VKXVgg2rcwKoSjGf1rsBKcTz9uhAG
061wvgNWYW/un+WtZy63NXuVN9CMS47cCWKaGrjTLqYaLzH/IQihuq65ch7+Y/Q5
JMcCQH4Mj15n6NBF4DHJCCCo9v3i8Rh599+i5OAYRDwDehc1+jdHJYJ19xzU7gNd
lQFMtkghXfINdR7pzxppf3K3IdXZEvM/d4tFJ4ffoiV3SKCsFgbQ8ZQRJuaMOvWv
o4URqLuxdyZ56w0g8/EAmwcr6Bjw0bs5sykqPutpU1gTHZKl3vcx7tt2emFDVNRq
WHjemgUlJV2QSMhxL60tv/nQ/wNK4U672eqm7+rYeijnBnLGD8r84iVEKt3htdtJ
q0+au1XSvgp4ebXB3DJlgwZ82DzcW+84/ySOiiaLmfu97wSND9MpJhdrR/YpTN5A
3NO2Zqmf9bXIbjsj8QfiG5kR/F3diijFs+zQRwhhdiFbiL0VwGrCyLl+NruqsRox
GgTn1RWigSbriLisXkQ7o81e4mQGtskJcJWIy+TFKSYxxpdFlQYL+c5iVkCNoDbQ
onMKdjwspG7Dr5iSl9HTWxjqOfZcJlyXHjyzhadGLJRLVy/SVjgOJWixhQK7Yc5q
JSU5ash4m3an5ynFYgmrQ6y7sxAGfhAXSi+s89Lam2l1OqD7x9Is/8KH9V5Yio3c
dbkt5I7jDvR2i2NCSiqB9mDpyB/nR3P9b1//3CkgZ8rZ9pZCTbJlaeeNaxAcOfDe
Oxsq5IPhqOro+dvmmJ+yJ1XkLbBHxNiQLRQWwTmVTyh2+yqCy4BGhkLKpCuOudYc
ctNb8eVxMxa3HTM6fdbnGgn5O1g1JUax9cC5mNIF2O9cCbAC3MOPJGS/u/VNmtoq
vJoFpNYHHBz/p9Z1rcEFFGe+03d1Dy7FVadeAh7XBb0rnddd1GfWAdI2YmONXEh8
dRO6Lg9cMKEVJ6Az1QOiuupxxmZW2z2WrI/IzeRwvDJm5lalFPw82NVpDzutoqSE
WnCssoRxvdviTOaOEcuURrpIsohOMBaLRLWqgi04xmHC5qzkBWfwDMu3SngZ5Xt1
3JsQHXG41qYNcqlyGhLBrEpngtDKJkvpV51rspD0o5Ct/WnpELP021NuAULL0ku8
krUfmF8zNkPgVTI44vSr3ZaUAF8AN2/vheeAPO/AZDuuXIM/YJ8+NkWBtWKFoSjs
HOG/5Uih0R3cQ/zqBLhCXKENR1jLnvC+isnv355yOFlfqfYFWz9LNr/RuAt6mOfd
gOpyloC8bx2qAICCnFw2QjN0zQVnP1u4gTZvr7HqCfXK7FxgR3RcwOgOIadf3Wey
lifnITwy/pS+IkvyXE2Tr3WRJQk2ewHbeTE9mGrpax7InvamK3vjwiSPcf/R2sDt
/sbmhBccOlS1+7Sg+0bOE0g7rBGBfQ17MBWDfFnh9BLoeUXIJV3Hz3c2MTWs6NoE
dOQD4L4g/ETjZ3NWs0MmCLX9wobrvv0p58Zv1mFbUcRBOTBMq8P2mudhdYVsREXC
qnWij+tSKJacPYDf7iuwlZ/IoUWraqPAxpsPLbXNfW70HVwKDmyA4xMoE1QdPsCe
dfMiOhg2dE5VywUlTaF5/YTuD/fELQcpFFm037NM+TH6luxN36ziIcstk10M1Z7U
k/4GKGrel2oyXGaCI+ctgOv3KPNj2CF2TSJKBAPM5M/GPyX+d+trswTdb7u2uChQ
gt7HHOJGUtUt5cbqUxtsfPk/Vb82GnIX7oe0WbliRrk6NTMx6VsPVpUKK0mOxH1K
CTPyqVGwmnmIBpT443gtLXYv161WqxoMJHvxv9iEbOgyLQpKOLkdHM0k9aZxiB9H
aTAvPYMno5tlP2syqD4VHwF5cTioZj5VuUdh4PZWsxOBbj9n7Y8lU5YW6Y5mq9C6
WYUjzB3+zcHpJojP2y6TlJI3AMMuljWhACEgm0aTDW61iLnQBoiS9HD7t+382+Gb
B/icKsE/mHUhBTbQe0mKZvntbGBlzRGx93AhHQ2tp1zAXIAP24oedjJcA6oyZqQB
PiGd3TMF+llb7ytjd7mr9crzN5Hhqq14opmrZiHzrDJClKDmt/o85+ewdeuPGUqc
K+tJpPfxZF2OVfEXdwLAXeA/CoZhxqq8q0+W3YdnBlFUZEe+s8RGKGo+4NXpXTk9
Aj6sjCD2y8PQvlGcpQxtUx1Dk050ubq04n6MqKkJUwtAV3h6PHI/eUyGkVdllYi+
0YqQ+SL4sMeqe/mJyJNq+p+Oy+gRTI/oJfxVBgb5PePzvBPU5iFQT5u8ZvCtYSK9
ecQ4RkjKT2VsvgG8BXZS4GP0H4B1MQuagmLQk7IlW0qzDmMX3XbJEEn3q/AlkmL1
VtfeB8hX2vPCyWMWf51WBiA+HHfGKYPp3chXuqB5cgWbV/DKD38BSuSjBt3yJvnQ
THdRP9nLnUGbOTpV48D+1aP9PtgfksN3xPXRGcAMBbCwgZlLiZfeBoIN5no4/Cnp
bObqLitvVj4PnNh5XP4pREmelYW556FC2btfD/POWCqnhwMnRf/yRP6+uruNSl3y
6FpZkpQ9cDA+cJK8Uzk0j3naETTZywesuBj2thrRGHQTeUMLXhAmQgs0Xi8xmOaA
4Pn37PhAe2d30lyNiByT2m2TvUcisWq/uro6V5WOE8yqWWU//jMb+7pT2gA0Qxza
iy7MlWmzS4tVeQHFZbIKyH0JyPn7QC2snac52Mi/HBkfP7js/ppuV0OwMcg26ZLl
0Gq+gBX6dP1Ow9efiBGgfuhS9tMGAFJlgmivviGGxneDkwmgtuKA6PH7uEV8Qw9n
G+rO4ZuMibQo00AFcDxRFHi9yTowGifXajIp//UPOW4daKRBG7oYo2N5/G9TURge
jcMOwAOEObMPiWRoeabCeE8dWn7roPv2/jAnh1VqBL6/yoaVopwP40MCwby0htCw
4Z+PWGJps/B0PJTDlNOLLC9xNuqhebmi8IaYZaouf8l+4yDQ+WCR/IgkppLy57we
2Jk5krGkgzWbxMcvDuRDepq9ul9JSMzkhpoxtIiTLKM7zuOwx3q37i9aUnaSq9xd
12injXt9WeUhNfuCO2nlEttO4aXy247QTtntLTlntiQ3qJBB/zTNwy1SSzUYJltu
PlBiVFJJpDkVDvT8ENxUwI2qjQf+7AFDDeGYOw1pJlHPbkDgPtpLv6mXJFcb9+ik
huF0ioy1hf7rXM+n8V56SIr1mDchh6AZm5XXQLKB6HSwoEk1LC7BwQaQRawnu4dF
Sl+Bi2RAlLSDxZNVaTRrLQJolH7B2bg0s+EDFCtlu4kjb+oHAYpYegKJay5DZ2gi
k8Y0dytPeh5//mM8scC5H7ffuQklCMG0pBv79AXHyt+XIr2RQy57NgKbPREUmkEw
t/cenLGkIOTdrSkDOWg0lJmJ4QL5x3+rez27FrWW4guvm8gQnppy11CxyxnlN+Jp
LYFujiwU5SAW4AeAAopluZb+FccXNiMffHVADLWJ0uSpbeKX4kxDXaxmIm6NAFRw
DH/h/12ugha7/U4pk8OAy1UHgYk4kUlqvbVeQv5LoAIIzpY/M8bgydmvWFLdShDn
tmUizNJMSLonoA0whrQzt2y3jeRJ3HUlvfct5S9EkU1Z1xg8v3HJbpI0I70GoMuY
43k5Cf6PFv0ze0m/SURdi0pld/JrtlHErtighU2ltGuz2yIiKl+Q8rep13YfgTh4
TXHX/m009RXRlhHHsiYewuR0+dgrYWuAFwAovkgGLV3NHBNoZLhDBF3uCocJchmy
8NI2SW4P/iAs6IWwjG1uz5obnpncILbPtBTsmtGMfJpAlq8M3wcHA7JrZod8NbzY
Ra85t6akOU5VypmLfeMuwVz4NktzaZtEeo+bY1G38Xqo/qNeTOfFAY/M/7hiqL+8
j/0pjHpD3R9RCvcPibIEGhv3EmO+V2/6LilZ4WfMufNIUn6ZPP+Qygo7t+uUm+LG
SIOunvp1ILS+5uqynEni2HkAG3UagupdQWB7azMv/adwLdo4gasyqqFf9oDJkqv7
msgmraMT3Pvnc4eQ7qgKNKkPJG5pSnVDwHuc5cDfTZJoMhnduzmTqP/1O4jHMLxI
EhfFzSiSO40IxDesLeAoXlO0/jwKyTG0jfH/S5v8SlHKNLaAsekjVOgfIrm/ZqVy
F3wuFIRIEKj/veHJaU1tsQl71pzxJHyf3+SIKJGey3uQsgGujHUG7tlRzHn2OJQ8
FgUcj5zj6Ri1eshNqd3oz0VMTSWnFeToJDRtE+myojBh1stvEbZgVKXbEPy0m19/
+1HnXwjEnWklEu2fCUaXARHjJJ5tl+RbD4kxh0BIXXBa+The7XR+OMEjLdWJzjeX
a4B9SNOdRG7rm/2t4lr0oWNewBHNQJdbTws1QewXFhsvHZwwXJuTuUFBvHYTgURx
btIHvz64ucSoaauN4ZijMpC/9cK7tEL2oFBtKxWd/xfKlYpaSQH9jVhtYnZcQsmS
Ryw5muQ2RR7uTv+F++PAQ5b66F5EV1N0waOYXjBnR/2bj9sVoyFwRTPuXAkDYprE
nUtm8mZF6KJ0tC3uRLK3RDNRrcvXUxNQzWiJiCMhe7bY4AJu9BHkJFNqqS7GVU4c
+tt+VEhmjSLvN8Fr1Zrfs7tYA7uMGeexBO9pgA1p8WnPGuh+ZDeaVIhyXUrC8W+1
/PkBlHdasUEPtFhNsjCTkziBeZG3bGNwL5ggMyF6DORW2UtchHbcKrr/EXT91MGq
Pvo4t0pCRui/UpREqp8ZZlFh3pJweBrKIRKeP5tHoMwbojGssbRTx3rK8T53Nv4z
NiK4bmkhE97N8onf4m10pTjhFK2k9xCGgJ7mN1BjLpaW2fwFsVx6YSEQeXqvjUtN
v0Ro5EB0CekryBgDjwTj6sKcjm++VWq9su37TJ2XcDfRjbwxDlrFSyDHUQ5OoTkX
a60zQ5CcWKXqiXAO3uhsZ5ZYSfSqQppXtMW54l5Old9n9oTfHKfrYD4E2dxR4eWj
vwMPbqCfEqVTanhq4nebdjm8EifqFsC/BlAPj/lwZ78+is44lS4X/0fekSLI6SrJ
hZ0VaaHiyN5zhczscMqHNjBVmpWz51ztmyQQr3ebkU2poTBvdzqMqlCqfWCSaRLB
IYtkMVV8Jf1b48NrupGgai0HJoQ6r8wXDzYBibF5QVcCvTL4wt3KdXpKUtW1uML9
bmgNEVmjbd0yuaVTM2RmxTLgBxTG25eUwYO3ZJZ0pHaB4LFTGqWXvuEdTp6R908F
UTWK80SzLMJvYLtRsY7AYkXBqyqOsu9gFA94EZiiI3gZqd7QGhr5uLVUgjXarhbf
5H9PZt2c+CVem4rlLqAp668trr3w0VPnrhS4RgyeTHyYYwVcGUgCPHIhQxx66H7n
bzMwSDOxpjF2CjC8ETVMTq3O8YoNSSatOE+WEjH+bpihUP7ARCv9JMy3Gq6owMKW
KqICBb1RaMELMIjVBGQsr26CkchBFKRQvbIrrVvykb26xr0Ik08NvSTIgti1iH2S
QvuYDQPZ3P7YuiNKhTw+T87K6UHNAEilEa+ujyJYjYVBzvjCcDQr72qNlKzdEbfE
lZmOB5c2pjZ98UVkDnI1hsrnb9WX6wJgrjiJWFVc5jSamWh95HKB8jUg7CAZYvgm
6kKFN1+7YfQQ6k0eu9oAG1PpZkp5xFYtW6pQ7jxN4T2BCzgOTkHqGd+3PfXFhT+x
erAF8f3y8oDCXgMuiNbMQjtEaD7ykwXiMbvPnUwScQQDw+dEwtAofJ/g3hWGM13k
Uy8B5tkz0WDG/wlaEMBSjBp3Qy2dWSSZBlezzmG5wgbNvX5BZ8DQ/1H3BIkZH+Ig
Lg1Nr0SJYWxGODu9QsiOcUmwobJHugIr9NCJjjFXMSKPoPXw6Qsc5vJxsLs4XbJF
FEuXFIrviTTvKXan9h4PW+XdtygjsoEHoaCNYReLJOfc8B/pOc4oPZ5Jm9akh3OT
taEB7DGpSK6eQeSv4ZffJolBjkwm7AJPvuJJBsW3/ZnlmiVNNfYzh7j5Ujma/9YL
wOfiL4bZcY5sH4MXUDNmIHqKgeHYlN8Yjo+g93anU5skfkhfhOMmZpEhQMnfg3fC
JAypwT26H8tTYOymMUJ0i8mNhsGvhkGRfH+ph4OF78h3kfCWQZf2R8zj6Lsecc0z
EXBBlN6VHr1Zl0Bnsn2ofGwtElt+SOuBR7gpIOlCNRwZ6q/3gmVMtXZwnvXAgAex
iunE/K+rBjfaeOZDAF38Va6Ul2I+9al7KbVzvS1GDmfFFkn/oF4DDlqXxmggbpy1
oucnB+yk/jFjSbKMxKU/fmVDKqT9yEIaQiXNw1hirBKrxVCY2ShQ0ZIRs+K7ewB2
bgWRQJKpBb0mswf7sW7Lj5eYRDamF++pJM2Bcx9zMbla5uD+LEy2Wq2oXn3KZynJ
YhABaKsxPBm0bQ/NbJUrajut4mvMMNw4Htiw0mbOSglPKHrR12hC1bAJoK1NCLTd
uFqht2Jx7IZxWI9ZBkzw1eEh3xSPJV7QG/+hcsN+KlH8dOfoAmGqan2OTQBIFoki
ypu8MmhNU+lwgu5gHnj2JdeMbIDm1XhH+1wjkQnysjdZxBdI1YqymDUkCFl1DdPW
an9eyAz37J6XzurAxn32QNAYUNJ4albh3QCKmLolwATncRZLZ+fZ/GhZI0JSNYRj
hD9kUE9ZyxsE25DtGypOS123FQjEhxYTLa6feENmer3XYD4zW007u+QG9ogtGPCG
bzTcBWD0eAxZv58K/sBJB2B8ULdQDqdq8TEtSs/fg1NNlxgEeRzhnv+cBiaybjQt
+659OuafqefX9smqKNHTygflqquyoUhCOxh7s1vdCgdR7gq7QUON6XUmxzP+vb+L
wrLM1YfF7vplpcEtjOSKuhsK9kq9CwHvafo06diGurwIpdgW+fzcA0Gdfd0AtfOJ
kruUbz8Am9oHTmpE6Zdpy5vWX3p84BxGXNOkr0v5v447wna8OI9DjT5f6lki4alv
w06YYTCjCK3/VqWN3RmsTz9bNsg8oZesKGx1uclQAxt5G+Xf/Kz19s22f4gTQlTD
25cv90PfG6kJ/gwVHQ7mN5CSC9wKA8WxGleLKw4ZqCOlYtrhdVuN8QUYkYss67AE
sbEcw83jZOsOW/0LmoKktwO748K8m5fofoTIskvbSqqKF1mVuhavktF7imnJKLlp
7K0kgClJG572pK90bfLJxl+8fTwnLdGTe2Fv5LP4X/ci6FacoM0g/Pi1qNNmdbYs
DuD0gKWYaicVDsPuF2DWnS3AXFuatHk4DfA7imOEylQkOgyrROYcbPCiwdNKbA9e
6bp65sWSurfbWtOaNLPT7QS9I9RAUAwiL4bsqoN8Oca/mmx74F22uK08cOHmDHIk
g7K8/xwpmKJQKv38hjVTLOQVgrGvLpfbYmn/F8DC6CEGdOWLH9dNd4Ol6e/lhurH
Jo5lgerooQyETDvQrF/IUfyZ8mrKEzqk36Tqf4ujm6ySusG/o+fIgwa/eIIBwcq0
qGr1O2ncceNlMMW/8Cg9zBtauORs+CufsnRw9d+koQ68GSM11pXVRHBFCxEbK6wk
JJhXOvLocvu2TEmT6ZQ6Mjpf///eMO5+aPt+J6jlPS0Od5Wsf8wxqkllV/Tw3yds
KGFCy36AwX2Ftr2LLAWP26Fba3Tfk6Ch0spVlFOpFbHE/ZB9nGkfrQA29oUIKx/q
37rwubq1ZwYGbsjCdoy/waIGNybh30tUJaj+0d92JW4suzQsoHJXz4SRJ47fu5HJ
xucgJu+dJnx8y9HI2mGmFOH6xX0Vi6MIx7aACaC3eJu7zhYK/I4UV0O8NtIOAlEo
fg+9bbIq2z13kBQEsVfbgK3Qfkmv8DZCJ/DK/0E6Iky7uZQLezSPEX1/yHrFYzyq
5GQu5POinghDYStZt2iLmuYTm0n3ZQXyQt/Igrdw0uwoUKDPudIa+ycLJ/8gCEM1
+IUc1CLPRtgb+gFt4VISrgnNOPN0Ds6b+hLjNUHbLVaUG3b/9i0zHRztMBARXrEJ
e0U1I4l0BMfnAWr1HwbFtZawkaMR/XL1n+3D9jWAJMJLN0bMR+aFAKjrKdQ5HbR5
FTX0jYHO1yYXTXj+iaEBx2SL2uUM2zJjuEIOH9vBMf6EeJmbYqjyje0nGq3M4tK5
42iInmUZjKf3P3jq90mlouHA8f+/u5FEubWa2zuwtKep5rgpfuEV2YVnQH3HZwOW
XVrq3fhvE/ajdCYEhjMcHlSVydYmpvNQ+NLNGmRe8O7gFoz1Fk2JcOKZ0S1DcZ+8
ur4+bhytRmBXN1FkYYjcb4EzoezR/ycuOnbP/yhuronPCcnpDR8brBX7SIcc34+/
ek8qoC9X/7GYo0NeqgAagtB99yQWZ4cSi2BlDs/gybmPFk1xD0o6wBary2sQs+pu
BybdsygEca/e3Ua92diNk3rx0ElfByjsrja7SYmmS21stgt972nfl1ZVgdizQiCj
yeJEbvybwnyt67qYg5oJ/jkwdj2XrzHyZYAry6kzQinmLiLWAw5dHiWekkxlxMjA
mw18GoWes+1X6MrZm+xCJSMoIu+LeXxHgSGapvriBOiGYfMno/fXLi4bsKESiuTE
2AlnQU6lAJUz2KhGroRGwRko1XD8rdkhX0r1BGYqB0ZQhx41f0cV6rHrh2YZk45K
Czae8jpPvJ0M09za4hzPbZ0sqY3tNinAKxtAMIVuGnjV8aoV7Id3khC84E4qOmns
wNI5SISPAxvVEhWNa5918eLaGxXvn7VES3n7KsoeMmgYmnARLR4O8l6qKMSbPFau
fGgiW6m0x3zkuvJj753DBKjrncC4qjqH+PTIlf9gYjM6IBpv0zpWucZFSWgs/YDZ
FU4fXZp2ykPlrO7nEEg+eXjmyKv6aBgAP0GhC9VIoveBVvUf+KiKqZ1OKuCGOiV/
KddB4eFlrQ6o0b2GJ3XRlwj9ImN+I7vSEbl13fh5cpe2ns7UEnfb88plawBz9QxR
blC3wq3EIj0jm6QAg8LqnPu3YHrgYl2spLZ4MaylUYtXb6V8eBkDDwmsi/+AB55P
/HLkg7Ikn3/yGYZC7ANUyoisyQ+IFkk6b/XRq39XbmP3khRwYJcpnTDVvdmw96Rz
PPrmHLLB4h6CrRlHvBoYcobJIq4cbg0RGXNhHM3VgHLQfljLiLMrvdFWK1LTyVGR
+c055dMYhMDOd7/Hed57MKqxeQ+K6LGM2UBWZm1mEnLrRoepL7TBQLHh6PDpmi1u
vbxAPinKotn8H8RGLw5Q+UPUHSH9Ga4QIxKPLH0EMSIwUTEKKNRhUAGRrJzrnZhy
ng/v/jpKKN8yRcubCBgKVHuE25hYnFyhE3ntuTTKBzx1+sjpTauaxS3HS/2M5zMv
bKvh91Gz4jM5hyLc1B6S35weEjSJS7hdi48w8qORRKHgsE4HgdYFe5t4O9a9FuHi
CstEU8kSQd8DtGFECHelokY8FmO/gDef4i48LBlQcL18169AubxQePUW+IiBBTYA
z0IPjCQX/KAa7Qhep/L+j7uxCcjkl0CLWImJuidax9IRPGYgyWHn2ay7WF0RZwHR
uwLErOYy9I3WuEMBDpZyC4ySBaDjvnkPeC2Hhp4hRjuDv9N7Wbx94DyLfbJiPFVZ
/OH/7mEncPWfvro8yOQPDg27FpQ90G4ZvJoebX33O8OmHd4qOWOEWRDbvANrLPKY
uiH1Fh3sgNe2sTP4Uv59BRoHjOEGwHOurNl5EridKeFPu042nzrAOe8Pi7PQkwU6
WAx50WJNgXSTbmCoVwoSLYpYcBYDEQ7wczrv8Yv9+B3ELlsOHeu4LUxGRSEJjBNA
q2aFTVsuIaZMEbE4VaD4sBV/sx/cC5dN9PgQhQP/QTfhBbk/3cWkSGwuPNsJ0C9/
bmKHuaMDNHYoZPdabz+MNEOELORXuHnXQPOvJ5fKzqxiAJiCL0fbOfGjfKPwVnpM
NIF22JE25SwC46USZEN0Q3eW0ywZyYPu0qA6mXpsbLRpCEHhLpbvHOT8c5j2TlT2
qWyd601edsPlWUd2uAbq84Gs3Sqfy1dotNhF0jz0lU3VzaMoMzq25meVfAhI3oFI
UvHv3JdIOS6KXARnRqXjaDhOCsXgB20XmWPfLjo+22CEobG9hSc2kFuv/IhR9Y5x
EFf+tWsmqwKXJBTQ0fMad2gcBvVvSCLFDplWCyIceRcVBbA7aMlg1nQrCDuAJTI3
EizQgwuHXKMd6j/s7RCGfUIiNzIq5vsDISHm6J4UTgCYzPl86QlKLubH/XXJxF6k
ByJ/I5YkrOkEKgszDfAlcwYwuXcTklfR++/SjD0gBE2XTACqrw9UPaWZU6akDX8e
GP136cQzUxUY84YN9gGXT/KwtaF4JBeyitppaAqW+lJgGTqiXIQhWJakFJJm5K6+
EyTzNeAbkJTahMFn0pAYpBN+k/mmRE+FYvLetk4GnSx6ESXPYIZ33us0PJqy71WU
k0FWNFTjoA1ioGZ22TqcUO5LxKFQ5EthheKMPDfRulx7fCGlwYoADH8mA/Kndtc/
tociovA/hBjEdNxKVLU/yLLr5dbizyte2bhIR8dHmzficjitHwBJpvMq0thjkAmc
1DqAZ1b2bE6kfGb0KD4qUTMwtTa57nW85nDAJmi7ILE7yu197MMLo5pCd8yVYmc/
yzOYomZuM6IVQ+fv9JpB2Wa9FMAnMPF5u3A3OT+71GGCzCu3m2PJW6DJpuvq18W8
rczGUyyC1/GAgHd9I4Jh8UZihX+ysB8W3U+IGHP5UnzQaW6WcZtFD5tPsyIycZRa
vMnji6W4UzCkVtgwPA/wdAAVAU1775Qgx5NZixB52cH2TSg6BhZaWOAhNtTcHR64
oQW7js/pwp2/LFkL3ZY1mIk/EAW0YJ2KFL2+WZlNcN5jx3WqYngWzzHxoSWuH9kr
beRbfzaXbZdew8DykHaDfm8uQDZ4CCnkJDndJKgcfotB3Km9AU3Jj+xipBgWioej
4ZpRIEzMEscx/0U/1SHTpBn5bpJ91U28lgxpU4Ls36YWgvczPmDcyaSvpdvVfEhr
6upunzz9iwMULAmuLeVnnNp1MwRxXNEJHcXxuAbQr/TYsb7RIOB0L5TiBcQGVTCF
CWtxD3Tnke7bN4ZkvshDZifQapbUjjA8Ikg4DsDmRbV3WIcM7pvj5OKfcc2P86gU
xsCYZokLtH1VHR/B9nJsL8kgE3xNxBQHqAgvZmqOLXUsYcSkoSbzDII2HYLC/YDG
47xIckTfjbNwIdNWmEwk6rIAQWT+1JP4vkM2VmjJxhHaDPPhZuGQpzF3MEHqi50n
hfVaFYDNr65zYej4nkyMXfbdCdkhIIo6riHposNF1c/h1rGKovOzc1y1KHz4eqca
O8nScUeu3b4n8vuv/oM6ZuCGe5KmTVFxRKQxQspc7i8VbUEMf3NIMFeA6dkKuyKz
LQkoKz8ueuT+mBfxthhtLzer3YYNCpeqKwD8Oga2G5aBzggsm9aoXfJQijXndokY
U90SuFcLpZ1l4CsqZwO6GPebf40Lzti/NpCKiZEowF/ob1R6Csk2lPvxfVxd/0Hf
A7PQy1ANCcspvt2OvO1n8X/Unrjpb+lIOqBqX+XqZjEU8OVmIegNDL3kYtn0F61F
tzdjjiAi7GXXKl9Jtm8SlNv+fvn8tivHS6sBmqSNUwxfr9cMtYi8ERGCrPre6Xfc
DftfqK4KNBsE2/cnn40H2JRWj+OBT+gs5jHWQkHGQOT6zBFtOMlDNzbKVCB1Q0le
A6rGI6ZUVQXZWlZJvxz0BY0+ARinH8hTx/UUWZLpaG4DXDsKEv/Bo2DmuSYLRUBt
owHy71YXC7xk0zgf+Xi3Ct+fuw6cOF9PvPWJ+t0xMhWxg9jirCY8cQgJd4dgsee3
XzQEkp64D0Ujzja33BZNGl8ljHIn0KIJS83fui0+TROI9yXyayQA20NTBK/xnvIM
Qja3B9lFtlkpqat4Lx79Efx0wg6aUtJ9U4uH5VBnDCuhphSrgZlAzQ13bJyaTaD2
uzGRhS1hR4w85GPjWIC/wEMAAsDohsr/WFOj28iLSqF0byYTTaA4JEgj0tOhzwLg
RURNeoYqi7yrkoQ247UbinazeUzCc2oUzpzh4oiKbztv/NXwoxxXrVlrdeCAOjRk
sCmarS9A+c5kMlq8jxX4ESFbADGRowRjOrVzbkTaLMJVnxs3eAzWSt7z/xPZPGtA
2k/cjopoPCvXxtBMzH7g5McgDH0sa18WoKUkoLNi++d2Hm4hSyFGrmyKkYQvMW0p
YVRkGuljL4XF09tZLkxOHCHA8F1EqKjChVVB3vPySyVZSkjjwu1pIXs2aEKbLlit
UgvIOup0pzXOVbvlCBueoMyTsFqTATp0jjjGI4OG2WaFkjqDcDytL2RatfYq3CoK
tzPTIkyN6PCeF3xuid/dHR+viFhpsKmJ5dily7e+puuCv2bL9xXHZyp+/OUjiuE6
36qS0rd0FPeJ8Z+RWx8w4YW1cVFitZxYEOm2IOyC1M2Zfl0nBJmI7yhfnO7TdK8V
7RIa22LuH6ZftJ0B0xLOuhba0tgMV/DyQ0Kmr+JOkMKD/qFU4gCatppBM7oTV01H
L/mqDaMISEQSJ8GtE4LCg2WahE+2yBvkAVk7S79i2sPIx3b2rCYN1uqCOJbiYlG5
Oi0bAwq8RkNJuEkLH0o+bQbTsqDk6QItBLp/n357JwXI17YYwmuQ5tQ5+owiM74J
bmoMOdNAWu/9uArbBKxemP7tKA+/aA+EgkohHk47qb6MV4QEcA+KULNJemix8mZ8
q0/OjDVz1H8iCfBgbggYotT2rg0lU/keXq4Sf3+Bb9BoqJv6UxQzyU5WEl09sm3e
kDRx/rljVlsbhYGQuMxQBsCL+DDlXuDq5AaW8P4I0ns5WvDxOHd4+Q3fWyx6dQ6r
yjlaike+ajjK9idSJAvVUo/EWbEiXUuv8HuUJYmJvLP6WIVSW8qhC25SxyVtxXlU
/9C/yGuuCE2spodhUGUoD6Kj/BwKG0dYbGQRDxEsXvc9dV3I7seicMZ1DSUhMcNR
jgRXc3rkOnjhpoxmWs1j0xyU9Z+l9p7qh372vJom5Zmz3J3DdXX1Azh0hNRUJnuQ
9kSaL7PemtGKC74DBds7Jr6IYmR4b0SKuZxkdqPcmQcVc/fvqrtxxeErEMpodupr
KuZ18O1JGA+4Lzh2NEqlkFnGeaEkrk9RTNK9xGhYLuH+l1H5Wvd07e6bBy+nmEGU
TlK3qC14m7ea2Myc5OURUBV+1kJBSwDFDnC+TatltoQm2EZJRFlD0m8uDCqfDRLe
ma48Mw+dkeMISR+DOPsbfrE07KEwE6208CvZ1IbsOhpnf6d9GZwMT7q2WY5RN852
i9I6DYTwURt67eH74LQA8fgbmVIPHwwEu/1Kl1EihJPIM4gTqj+sPXGS3whBYtAU
9A9snEKshXs0jRa068BLirktIHPCHgrDzxqm9z9I7wqK6OWjYJWDyyyNYZ97XBEY
gZu2D2J4rQDSmqQ5A2AhMEgY2KD8pD1Af3zLPCuSQko2wbnlfIssI/U/XHFMcipU
7HxMX6x+vxTgeQWptTLT9/oga2X1S85DcXejTX8pp81r3GWd9YbyPSto+08qzler
G+7L0vpbcil5ReDrvCR5y9/IjH6bsZxKQUhoH79jlVQ+L1lH7suP+zYOGeLGHdhl
pnR7znVf11VNBwcboQMJH/uMZ2/VZcO2k+4tFJmrG44p7Aj/7Opdc+qHOdpAgyfS
L/OeEmdQ+/fg/OVO/DgtpbAFrPNxxYIeussFqUNzFuv8RpB4kL+kTv3PITb/T1kl
8+SzAID9dscJAeAWE0BISQQcRI4+TyJsPrBNUNce7/AC2o30gVL5dpL4gihYACSN
zUakbZOEb72aIAAqNUtYm51s/ounbYX8LxnJwX4fvkfX6OsIt/SEIgogzvjsot4t
ri87+BZuMb8CL3+4A4GsLPnXdNDtuvC4ZzjRJ9Z56FQU0/p3Yk1UV9Tm9inh+Sw6
xHWf/UhVDKYgpGjf+g8YTpBUHirwaZs0wLrZ+G+0CsWi67YXHXSkCG4cJsIjnuNz
wO35MZE+cbbA2Xq7NeTncA1LeId/JhyOHeDbkY6bqThy0j2nfs15/Hm8a58rkpyP
DhNZ1Xa+fdcujkM7KVGAnlI6ETT2uG5xEq7KXfrAKkpiE/ME2qYylvVaTtkMVq/I
25nO7LnupZow8mS/TDLY2+k10pKP/vp0ZUOV2BCdVDpAH3fUnfQhq5d3OGYHvSk6
AjIhH/uZ9qpkaWz2C14eQK/vvndvQkBM6OaZuSc+H+5YX9uUMWkmOWqNlig05AjH
qmnwUTm9S+CjBU+pU7ICfe6div8y43Kau8x429hY5+PDJ0UOwsVIFsLZ/DXfeZxn
3u6v/OeK6O7E1gRKpA/8OfJN72dpStdzIIBoAAobQjtIcvfobKJPXNnfSnCobw2O
OT0JAufDyh42oyIgh7H6OH5yLxNcqqroi538K2OdePiBiDfkfXbEMBweFWx1aeYM
uFMEo5Q0wilQOVddjOGzemM6LL3hBFkBK0wyngbTt3w/qchc5iUNS3pR7UvWYXzJ
j68dg0ANNmMAUW7jF36qO0cvip9q/h/NsRrzXWJbOkmzf8OZ0HbtxpSdgLC1EOa+
THYDc09Rw59lFrHovbjkkOF9qP6KJpqwlWqdPMieoLF92YQ/n8HxEnalZIM4vOw4
zsx104pcs5MgxAyaWuq2tTyEH9je+TdPunNMiDzcCotPjWgptLmasiI7khXVn/GQ
E08tmf44Jph5t45eqAY6K2brcg093KUGHaZp6JVjVh73zloHFCirG9aTxx8oEGNs
CTOWIN4M3hWozIBsMxe2SBMWmxZEIprBIUIw3BzoyJROFopT0ljemWYCQqm9UOyd
xatMWffsg66fS3MU+fCTfxFOOU+Tku31KiSa6G1PEguZ93qVBGhC98sIG7Z9l299
qbt78L7eH5cNalicdLnSw9zI14MQbLrUULbb9oiyiDeSsRfP4dz55YqDgJ+EXWT4
v8kEgrnRJJkWPh8x242vZrRsJPLjB456AXzthLERR+8vH6WletxIeXI9KKH1pPTy
C9LWa7fd8AxqpFGVYCUWYaUhFG74NqJSC45XBs01HFvZwHxEr9j+DEXlnshIAU0Q
0F15UmFL3OBtj/DPpR8to5Nq7+JL499Fw7UN/Pnt7XrlPBqmhHT3CDSKX5k/dJ4q
YZ9ib+kRgLWXLVqRDGa2aCxm9rUocnpRhzyX7j/OvPjdYVokPoPNm1MvhiXVQJsP
ZuwP1RLsVU5JH1gKRb4E0Vc8VuzG5WMzj4BP36ECY9cAPiyiCFJwFWcDJ4IMuvJN
jOxGeH2KEsdKU/MfTuOUkBkLwbU9OA4jfd2dbAqa90KrsTutZn21Pirx9LRLp6/N
ZPwDLqHjGyO9ycaSBoPB/P6TwW/yUqWDbTq3q0GkDD9kxBydQxyxyA8rr1q1Sqwj
OKwuhpy2ATNl70S5Elt2woTzm/SjFTMAgkbq1GCLMaZD+qlFmo9d4MM5tUTV+KLx
0blhFulTx/wxbguJ9HJ3IJtMvAjJE4TXJOunniqlI9P0i27HJu5N8CREwJE8P9wL
X4m9DYbushkW75KHFb/u2LO5qIHOXoaJ1OG7INaasy21cSxVtOBw1Y+TI0zCwDHx
hezTovAbyfVdvbvyo49wlR3LC6RyBEDpRFWyVIC9TLM/siOQETIuge3Hk3UM0wPR
Ym8r0NBAkO+C/qkPpVuVqlvSVAqgXdjuP016rJKa5hnrIkYbgR39zsWvyg1mNT3b
RPazI9geQQ1qdT2p42o2aLSWkVuqJrpCnHBeVgsOY40JAxGxRhw4c0rA21Xvt6zo
d88US7gTMexxFQgFaG9lRfQtyI6FFFck1Zehj5PAXWmdIVfq/Y6/ebR+e6FSSF+W
S1XNoFjD/zsm2e6PqINPmR5HUS8HgWWK1S0kfHbsaFK526i/Foz+3IVYWpVb37CS
6TcqNMHHW3Ng/laNhooDZMffpWZa6auftYkFVNPkA7Jrdzppm9rU2JQzXXW59wa3
syOfiBNiyUT4rJUnHOKG0Kp1MNMgFZlK7LazsBww5i7SLagVL4kK5mK0lC7WlL2/
Bvea3MT91+Gk4eJRQfHjUYzACHX+yXGUZPyvmXJ6q0HUwpvrQRMseI/z5wam+hhg
lttVJyGD2Pxkx4CSlucmB+pdz/4YEzI4VyDJ5uw/XejLK+tVHD+OlH8Y1baoVQpi
ZDodUyaWbWPygvZ2mpa8H33s2g3OMbZ/po2odfX7aRP3cnkNF9jouXdNsJrNUdFg
rul4kUAXtXMOE4X5/psKSUkN3N1W1JUHpSx+dM7eIChIbHCqt4vHf4z3mP2yFHrt
9gYdvLek/+IBLoLQH18pxwNwhuQjiA8CNWQDtCpiGjtHvTmYdsMEwiPrwtMP6B5j
87DR0NjfX/yBcmsoZN9TDjelKoF+RoWmadk1Vu+T1+42uQz3nsz3NitQZGEhbDKn
rEfk6joGXG7E9Mw1WuSZSr5xa4lMq9+RUZyMUHdlDiaugOmatnc3EMUmG8j0Kuud
wcn/3QV63Jtng/uA5SdxAYG/aN8JcCg99bHzK/JTxV+6V8tGpkZnou5FAW288FVf
qD3IGxeCt8oBn3kNAbsVhpPAvJzyBOGUn26G4e5bXYEvMOfX0r+TUnl6jsGvj26f
ipuu1iAGQS3AeBfxbVjfK7cQ99WwUSOk3N0hyLzxbTdTXekhLjGazwFtvYsIw61B
jTAX22jLaq+eBF8Og5qEfTbGlpcGh7sVBbqVYp7fL+jgzpu3zumr2Y3v4eLdglpe
38PEPT4HhJjk06O4MopTw1Ol7n/vwhlc5FJzrXIdiUDvehSUVGCV9mIUswkYKbfH
utP5HBepoxgc6uPmtgqGpS0Pzu9iSbLsOBnE5wUW/c156tDm819vgGDQtPjXsnAR
8vdh495VdmDCWrWKYwb/BJ0PYS6iyLoLg07QszrkJQaqjwGt5XsaICjmSgEfbINk
W5qFXUCthrZuXT+144qJN30/97o6Ii9W8hvWkqytJ4SyLiKu4zAANboZENtgFXJY
ZtlLvNFdWHnmryGyNpce9zP8S9IQrbSlRLRI/YdWUo6BFXPORlaxLkYzVGn6/PiF
qHy0zvyFl29OtmXcwh7+0oYJQfe7cHWueMtxWBV+SWwgM/L40csJcCTFv3ozkVwI
AsslnrqcCvWPlexrtSmje7NGZrie1RbLwgNWpISG6quwSzVoly35bRNSb9TdhNO+
rAXdD7eLYQW+nG1c4HH9nQoCjDk/tSTRJQf0XkjBvKLZHHcOZ15wncV4VrULSGGP
CEX/TDAR9BPOjeSut2dJxpcZ46vy83tmuoU0pESinlB02D0zjqQoQZImCQiIXfB4
1irfC8WN90W+/gkvMd+22MfldDNpicaaLecAWKP3VQiluFBBB5OInTEd8GcpOEky
I9c9XlTVcQRpSAWeMgqm2SVp0+WnQ5DmoC85/wDB09c/zEn4MrgHiY3EGIBgxD89
CCTaczORLSKazSuRArDenPhDxO8etLIWbH6PvCHpEDdE38Ak541YZ7pqdF7MRe2t
wiLM2gZw1lDnAmOYfQdPofzxAkS2LBwLiqkSKAr57hX2+ONl3ihn5h1T9ILgN6rJ
kmu3DLFDq8tvBFKeOtzK0hgWvlCqCajCMahVAmdooY9uZcZbPc5Xc7LF9Q1UYs5W
n4aBbM2ND5Ju12MmSqZY+GH3g9vru5Lm6XvqepAq3uCsdNcEeoUnP3N4Yl1ZpvFm
c6TjouZh0Gj7b3qIpqqft4nOIwjZVvkIazuvEKkby5TQKYOiSfgmvF3lvoIVFMeb
TXjwYsgugvQZyM7JuIC3OS57moONHYI187ZSri/x7bDP/0ZYnSxBXAC6vciAWELX
0heToCY2UwAz/BdKuYn4bSoA/yYEAFeNcELm0CV5US9i9RZMTTf8eelRiVT16RoF
ZFJ1VptkV492EVY1Ot6mk/pPxnl5vGRESbH8LKimSl7VLiRzxq5pUl1d2BdLtfgq
QgTfQi/aZl6/n1ekYiEe4AlVNwj2OcFvq4QM9ooi58oOQuPKWS0yoLDbIyiLlOTF
jVNBnXNsZRQ+B/jFb5x/OVhhc5MUc/P0MmYNfqSNN9mrw15VDOqn+jdJSmvV+y/R
TLyw9csyAScIfSqeleXuNngyCtg2wvyuwOARBVoOJ8ps0JpXG8AniFUQn+ONgJ1h
dRynXiirwOr5kZYlO2QLj/3hZyTc4KT2nce3sKJkdyKnEX584Bh32tAjWL2Zddml
algtBbDMg+WYuD5HFcQEdpKDX/S3aCI5yVZsTJzKQWzmeqQm3/64gbCB88rgO+7Y
oQ8GG5wqW6L3i3KpYwnzX/IKz+FhpSJCCP5ksLs8jlwjAerZtmugDwvumR+pdi4m
K0VvR4VqaH4sA5akHx4ghPQAT0TEVbcfxQaJR6lKDyTCBwEylQ+p9KvAXFIpm2Pq
UGiHHteG+7QQp9qEdecyzUK1JyqTpXN9NrAipQRLDrrnU/FkLYuKmtRdJSZ+YIjh
cjELjDl7AUtL4u+kjZniHbwiqn0AcqUF1t15QX5cAhcsR5hlNwdYRdc3EiEoHdzT
z8thd2UhyenZ/xJolQ9VDco5rS15ORdB/ov4kw2LqBDfmYU+MZ+wwhM4tQH4GJqd
bhdZJjxFPRiLq8E3NeJ+bKUfrbxnzQZ8z/8VFJl+ZQL2FXk2RU/D/CJJ6iFei/hM
vQHucjfi6XUMSw0nGR0tIKs6e+ZYPxIsJASW7uo+Lb85L5TA/JZDztGzajCeUZ/l
kXXxIKM01VryifhwN9p6pBgApXulPLvojldogMhwWsevLFA4AacLj67dyS7eaTDs
OobdiCYrx85MbjsYuolzEB5MMArBKy1O3DI9Q3IavUk1Ctaua0Ql2PMT7xojD4wk
wCvG7H9OGC3hq+aPwp9XoD6cemLGZ/lzJmKZ37iz1XBnUSshAiwUaKCzO/UinSBv
y1NfmLfAOmdIvCJiY3O1GVDvvaaxsR5jpevM3+Ww9So14j0tFDAoz1ZToKKt6L6M
2wecEiU3GyzflqofCC8lcNs37DEf9AHrm+sMc7tCH8vpNdiJQ7cVV2paZRzYU3LL
ok4zvUaLONLikQ/8TPlsl8lAPRBIlVuuu1R5Rt50TKvOVr7/IN7nevyDIt2pVLAu
qSCm9LZPmC//cjAUdw8ZDW6A4rWfSQ7Tzaa0XXkqblX8mzWEMKGq/ZniSiYcVJI7
jjD6EZ5wO+GsGQIxbGLMNsXf1YZdiblLGaV0u9ccBuC4zmnFq0DrFxDMnC0TmA6B
jpL5ThX9iz8crUO4XTU0fNjMdNHP6onWakYe6r+otpKWydhDP+PvmDBqQVfzLV90
L2Ph2/KGWTiZPZuDc9uXykf5D6aCTXj7owT02euQATLLzfRECsE3tKoI1s0m3zlX
ryNin8NO7L+JCxBb9I14Cu+Ae7ibAXD2VUSqHAay3eA+qDiV62wlcoUuhWA2u8fa
Tj9ejIGURgxNZ7nwUrJsFU7uu/oO7belm92faAFFwqlWRrsQX7EBoNwiHnOEc0Kl
oRdR4PoGzdEwTuIAw6ttuiW2c4vXqCPjuXaOCsEjiZuxrxyf5Led4VlfuTGmcAXV
q0zMZcqdh5rfhyD+hAkCDjW9d6aQ4kXAaDllkVXkyJkhV9aaqbrrjvr4uQ71FLNb
2hPvBnQZrpnMI8WQNFe9gLo1KMzBkM/uv7jeRANMsNCiDWGNXGiqiIZPqpOU0EvF
qF5EqKcC3sBEgZTpZcXdyZAjE8NJrXpE8zG8eUK/J/PDyF62g3cmVh1JwK+dRQi4
KQ/J4adp/yKlSiKnHKiWPIKxCd9WTRNetv9vbnV0wJldwUiMlNgwJRMYuGPim9Br
J+MWM/0KNT3Sw6rVcaVgSjZyNjc9XgYHcYWrTYEQdamlGj5pMIe3H632WVlXiSM0
x9XHI40DdUVMD6U+bS64cU36QeawSqjRvdNUwUxydvoJWH1zajQ5tokLTcbHew5e
piWNz85XdsWdxFCq48aaMl26fCq/rjVXOTbCaD1F6H2dcvIDq0NxpvkKcZ3Zjv/D
C1lhCvlvGwJT8F4h2yg8QlkGRh542imTcuIicPJfQDdQeqs0jIeXmO064BDG0Vn0
owMVS594F4xCfjVroQoKgtkDzvTfRBcjTVpvhvBhZdiU28iNZd+Zs03B4kwPHbH6
UZLeHj2tFeVKb9jJpL2HXYP8uSvRNB5R6dPryvz6vUMwRYYZoX96zKwg2p1vzkso
tGpcYOEAUemXWYZCkZSDi7ZdsLxeB0r9o9jc+hwjs1nfKU4oaiYAU/hSqLURYLqm
34RGRDLVm70C5MJUzdTMNiqOf1IyTyBD5ectxLNuKbkD/s3o5Q76B4sJcq4HS50D
bQHDJ7Vw/qNDdtJ2ragNkYqeU3SFhl+7zB0O7CLEjyC5PkkKcXzNFGD3iiLMAqRD
2MSyTX8CTpQBFcg6/YE93CqAeQKmVP5UeDRBULeIZhJGXdM8dWRKqD2wgKk7JdbX
5BTzAkAje7DCK7ZhxNGQXThStIcJ8OWE0k0RZ3KsLJrC3u9GKlIZwivt1tvLDmJc
QrHfKef+EQVfXFpFtdDcXhFWNSqqYvAwCONMNu0sIEJ9xssSv2O1yBM5j1d1eEuq
g+K3CjBWdSSs1ndxenKZzgN10q3SoSN38JcBpPSAHb6RgEGIl3XNEO/b4D7OjnGJ
FqNUmNfQoAe9VPVM5ZxoZjhNsSq04vL3CQaRV5Ocrx6S93H41p2ZDQzqM9mytZSd
3neQHxGeTqOVDF7pdTxdeIfI/c03fen0cXiEQ7Ya5JBzkHNLElKlWI5NQ8G95FNA
1tKHyBRS8P0YY7W/4u3V3NkbgTF0Jw6j/nivReTbJBugf6vwYjsL+RDzQj6ymRWd
QVVwLJ6gzAd+UaYBwEAiUxLu4tuEyhqC00TgAY7wVC6G9n2CjvwWcAb5sU8MkV7A
mZ+q3Bco+6UdKWKCVtXlGc7n9VAIU2Xon87kRqD8UY485+tG/oez5no3xP4zfmBE
wv2SPr2V+JcitZaXi1C7RMbnt/QFNbm5pLQvRtWJkgzRPpzD2h9vgou+OB01QhKu
0b8YkFUrqCUQwO7omY2Ip4HBO1LrndjddUEcu5sbB9CnNGQMfGTSGdbpprbjAXVx
vUjO8AWOlWHtfTjaB3G1eqaRAHayiqKxbpgAnpLpLXSgkFzcqDiEb+8DWH9N6lJ4
LY7nQ5JgAFttswIhflEpF9zwtbOg/gFn/LBDv6ONK5y3WrA47kKRGQmYvTTsipyV
qguh0HG6fOvMA42bbycsX3QyynClFzaYTs6cT/nmmZk+M/gJDXnmnPLiB6jm9oUX
C8U5A6uHoHF4RtiBlt+Oc+2/eJq3MP5zbAZ5MQjju6lxr3TFDPQRZoJsXuqKAYJZ
jxwG7pd4neYWQjXVIcIvBWAiMLPsYXSDuBNTGTQgtIaxYuhnELIZg3OsAt9PAK5e
PDk86sJNOhcW/mGR0xRc7jNS3xQOzbBlbdE/LVM1QXfm54TqhuRqbjpCtJjdw36n
f+VyBxwqyo713Fgdtb1bocSxZnFKz5SkkETVtE7K+dEGz98RC0s3W0FsZHMONHRy
P5Uip8ZTS11/IB+tRdV7/bJDyoH66Ys2EhYvpU4XZD00WRK1RJpXEShpkVksAq/y
V7GJTSp5g29EUZbLs4rWRpkwhtyFKEH8ifuOm6eXfV7fchkTlHMf0r2zw/q2FlcN
QjZDX44DTwsvEFBaZd1lMUuVV4/hIVsxTIi8kRF1EduTc8E1UDJdMGrS+LUqO07V
Z5h7UjwI8Oed356NMaeLXsUngV9psoPi9oPMcVjHcc0qo02eua23dg73v+yg3lFK
IRu9yh4t/gkn66GqcdA+dCOYuToDJ+wRGKr9r/31BhC23T9iBvdgj6JK9Uzb0z1p
Z6zGOmMxsBK5YZn7Q6ncDUu0mIQOM4wrMx60+uWAM4wPAD4y7RhfFrEaisbhy5DC
ftIqVj7nk68ydRxRsl4fev1kzHaT0E0+a4ffv8mz7ccnfArwrrvYHeqdjUfyOfAR
rGkzzmCIpm2dsdJGBwI6RIj1KCrs0jxkXUoYiHtVbMLETaaJf1mp7p/4emSAc3jp
aMk8wRBkjn4fYccUvtvSvdU+jWtt0sNb8U9JAIDynOjMEH+Uv1UItwLXKvs4W2dc
XUo1DibrNNe21vHEY0qfLTniOoCHu5YuHzLsTS0PKRa1mbvdX3lFPEJEzyy6dFam
tGItwan7LKz0ufCUAM/GdcrHGBuXoYqkjpu3UwW7ubYq3pxvpnxUf5MEcddWU0M5
ChBYYY9C4dZE36pDuOD3EKtq3TM0OZJhucCUMIctKkY1QmukX0ziRpQKGyJJ+BqL
Gm3Y2OAMNzV5NwukaWiEKAtIgforBvRuicwNx8dfhPlpL10XVPUuQUKyRFoyF7Vz
SNfhU9SzJ22O9UC08JKh4NeZud85hueRpzkP4WHQ6ksfeNIlDY1gPiwhANzWBsmw
+PA8sfqK1bYJRft5sMk+MwOf0DdOG8yGlVqxW5MuGrNIRNUIyyuBiXevOadhgppE
cCWBh+bQxRWp18TZHsTuKeI5SmtcD2lLRA4AIhc86Oxx8P1X5pRDnfIEyqEJSgg1
qTo5L6g571CoSxxyE43aVj6J059fqtUCxwgc/8x2ew3IqgIBlTC3/zLvD4R3B0rU
7xcRM4Isv64l5Kb7Z9WrfqC52k7R7RoxPzUvZ6RWwIazHWsdlto4mukGbGZ3o5v4
cN6jUGESKwcSa88sL4rR0Pc4Ile8SZ+VFvdlB8r+IE8y6pOzQp7ihSe0frO6Nejv
MUVdaECWA0PcuUCIwtk6kgv0KpHWhQNl06DFV49r/ZdI3Z3hNsVH7i5GGFmYje7Z
wCnFMNb1bnhoAAtnwsJJyjv/zMHRKpytTt8TvalccprkOcBNrUCxE8+qI8C1aQwm
o1cjjLXLWI7e05Yu1bbdaIsKcXcA4op93lIfkiLIwi2Q+1mzznns+S0htLzz7WwP
VV4MmCDWOsfTiSSOKMxqaRSJlkhrSEDdQ0AOTaXre4YOdAvVw+b4H3rtNsesEPlZ
jWMr93VFCIWnRZaqhFQf8ScyTAVFoTLNlzT+1uty7T0YAJuzKD5RY5IUZCnwa4Kf
jNhyZkkRcquLjxdf+ZDt9dv00Zfy3Lg+yqzWv1zQ61HF468uSlzb/MoMZUdWbd4z
q93Z6zKmVekMb6KLmZ4y9m8g4/d4/QNQCT8a2Ze4uiKwJ/7OSPYUSniVcwDKZ/9v
nr/2a4XtYr6rtnvPhDHwmSAnhLhhRU1K3NG4ValPc/S4rbe3JyY79Az8zS/v1t0U
27D+xepHcZJ998lfJ7o60i2mV/lwoeEtrvXouESHTsDghyew8jjqM0P7en8YN4Om
m+FwhBBCjXbubn/hHICQ9LGdszEwLoMCiugw5Ol9phvFh/u2m6yh6CjKDN2fjMEF
5zTYf9966YvmQwUwtFWuSA6B225h1bYkl73uqlNPyDMWlZCbkWwxrL3yh+yl5yXw
VyE8gtHIuiwFIH9oNMX4Tu+KyV3WzQDdIi1i4PjAkn9i+QRYFGM+2WOrdJkrJxMZ
CO3w0NBhep4UrH5EYHYaPkkVQ82ifXRUc6HTi2QvrZB7vFS2324QZ/dbz7GTjq/n
7vHej5MzozqFS44yLTZY5Wrl3ilwEf3+apbt9SXFITVcSaq/emzXCBUUNpRpHji/
hAI1jXHMfCijGFWTLnIa1exm31E41RotxbdHloeSiXHWDtB/I3GPd04w92JIfhd6
cGDxVe3INLjqIGzNBo6wOWibkUJRxqs8CPK6KRv/f6gEL896eUuedfHC2W19QotA
sGK8FAf+SK3v6yETwtHYFyc98NOEEsRAwYMG2CVF6UGrRWabsJzoZwr8JKUJgE+A
AQ66MsDfuHJmQd0/kXIEjxvsBop1ZC7m21Kd8z6a/I3Y+E7tpSp89ZNZEdLS9Svn
RbWPjHPMkOFA4JZ2I7a731Kqsi+ye2O9PAOQ1AjIEVVFtZ6l82NUG6awjbPQgCxI
oQLwhHAILhP6PRoX2veoYL1qwbbNQdgfHEfHMzyvXQAdBl5ItBi2a39cxnYxRH1W
gUioYNN3iNFUGFL/whNBg3b/abUHfcDTx1G+Q9DMQ3ZxJT8P2CNQoHnFgVCHtTji
3TO59oWvIJqlPsDgMhzrdFmAue/gUyh6Jl6EX9lTd4uC2Sp2n3kWmvgfi1uYizvz
1e14KoLcLKypgg7RgGNYw07EeF28swO2MC3I0GqhTgefnqta/j9qDqACXqX1YTmS
7D3UfY0skSKDMXyRaJy7xU3AQ0c3+rIiztIrG9PiT1pq5674RuRG1PCxA3bI1OLC
E/gpbWi8qS+hwELidSFxpf69jUKwZlJBysAUsInv5rEyvfmwoQD8sfHKaZB+jHpo
mV2yj2ZURA9Sfy/XWYxboc1WiHkAoCZg2PZernyBCK+/gcmdWDgZHXRONXse65SM
E71ZKnpXkMo4A5+w5JHsPqD+GiQFCyfjc8q4Nw4VZ6zaijtgi6PpNytSN/gG4JYe
25hA+IHZIHJeVg1ltN/w0mTPObqtLe/THqZ1/p2K041yfQfRXq6+mozQwDU2dhkk
3c2oe7wz0Xm6WBULuOY4oKgA1kmKM5XEg5IMjWh2IOhylM1GjhzqiPUpjw7hcUa6
qRLzWrgkR28hnL+C78LM81YgTvrek+9v1wyfDsCtkSAZCVdd19khSTT+WMsdZW5S
VGe/yaBwidwyFfkqMn2sIyUCcK0m0g0ZEvvYXbldq3VHwxHIG6enHi4AxQQx4Ac/
iUMJLipNpPZKCoN8oeANxMFaXK8c3Wpo9Ey/8i0J2Z2kPd1c/r+jZ+UvzIA5OIvR
I88u9XS8ik1i0zPT5BtKoyYgNHP8J0E9u6T35ysnjW7X4D1w83HHdXq+4Xgj7hEQ
azRRUej9HsOMEc7a7A1MM5mGAfuyB3w0rIHwyHuwDA0FxN00NbiK+TVhVPwi6GPx
IiXugCL1Xl2ryV5mzmWifC0roYuleDaFgEk+LJ5wPp19dSbDTEgVsZSSBZI0q+br
Fcl7yz3hY9s7Tq0C3B42hNRGQHkTsJe2b8RNWXbioxHCu2lJoDR41To1xU53RiAe
IjljD7ZP37Dcs5aI3ZR8Pl8618UF2etWV3KDAwRmcYEa7MwesQ7uq0RJ4rrlzQT+
tJ+2Mv2hCOFvGZCDvcJludh3+4IcA4zEhNgEt24PoIXhFlykmFP0maZoe8A1J9xy
yDX96hhSA+fkzR5z3/VUmNcFsSfXVkqMmbeddS8QWsufwXFQGklG62p9WJJeIYQr
dVa8xWFgdy5OUNjBznNagTuLRvW04a1BA5hoc2WQnZO4FD/dblt5F2mfM+OYlO7l
wDL/uziJLkZXKLN8zi/YKUrkN/L3mAdm7C7jUPRYBuuK1oKBOjvUaBhjRc9Bb/W2
zqmkTeieWp6faCGcMdp3l3JGZtWSnp7ePZEraqytqeJF68ZVaOMG0Xplm0DLV7ZF
QBWp+khV65Q08ActzAM3Vn19kdSNT2XiUxarPAyu7+2PQbgizTWE3YHpnMopWWzd
z2I+4mEwMY8NSA35DyANISGY+T2el4YQx28Md9Ynxt4avJ2p4muWiz5fzfZb8EDL
h3ikq4ZWlM9u0Mjiw/PWRkDkfOJUrymhNisISq9eQOTWx2rFp2YQs8HZXBi+CrFv
aBy636teJkwHxMwGCaYrVgwuAl5YKCUPNyRZSUnjlUuwaljm+m8Urm71x5Vx6iIA
jaSGP9I4/3/iU4cTpssMsSRSmSUqDtvWg8k4sIFxCUTKmLM55KxsbQKVAMIQCBPa
xTo5Xq/quykOSi9LhP5JrLJ0f7HziskpdWJMDEZ5iq+R8KoflXf8cMK1bUvTsqQK
u1ax7itq6LstbtI3Z6tAvkL+WAEDQrcbKgVtznpZ/psh/R8N8Sg6NBYWny4SREdu
+Ns5DBnFhs/8DVG5sAhVr6fh2yxMKh1QPxfn9HB7srJg61vRK3zlh8UIcwRhFfI8
da+q1qvQ1h5w9dD2gRVjY6lZr2/A9btDi1ASHMtWO5/BQhUq93u2eA85OpvmYUvt
Fx/NTQGEvWWKl2rW2UbTau7fJFt6W9kTYE/mufLOmh4YQ19z1Dlh1LuWxP7lIKZd
jaGp7U7D2QAa3MtePPtTYH6ZCt8rib3j4/9HmjMhtfrxJtGltxgtokC/v94PszRi
ZGCs063kRbmMzT0uPZmbOYXP3dzE/kciHa7Kk5PG3ZlrUUUIt12mjsLqfxOrmWj1
uxHYgwk2vmktAONf7potIWac8CvmO1NY4BXE0eoSpAGE9iq0q6CoOJfUJqkRQXv2
y7/5W8yltQfNNq4Bl8mz3FYXHHaJS8G/NCMhd+GnYDEckocUtLZMF0dkfruaxxNi
IYKpoKkCxFqsboksz6Dq3YPg3h3Nf4wiDwH+vTvRn2SLhohHUPbpQt/gqiSeEwg+
VDiIfP8t52b6mpD/On9zIog/SN7MRAAyHDoE9SWyRoN1SbOGQ9Yrz1t33vIx0sku
1/isxHVzlpFNjU1PjvqXtnh11zb2SiOFdsnNnAmxUpF525k5EcZnWq7wX1F3z3Hb
u2ezwsLBE+0/vaKQbPiCfkCr1CHQA1kd+OCEPTcYblg7SWC1VFy42Nr8lY7Xp9Mu
oa6VwCpyG4/MV55kedETJyQcz3Y2+rsOAgefNaN8NFjoDCACIrSNawPfT+m/JUdQ
ErKUAXXbJWjQnML7AEDDksOiQsq61jPQ0p9x7xROANckBq8fyxqfCD4Fzawi5fez
jHB5E0FxnIXrjTfoqtuTUn/jrEJ/BuPJsUWmvidDEnhO8IjrLdTAO8oRPaDKt8Yj
Snyc/DMP4CWBb1OUzX4nO4bb7O5vUOH+hTMSNpeQfOaD0c4I+LDjhofnjFjCjaWv
6qGkd3WRVMvIRwbrE4CJxZtp4qb3ELO0n7gpEEj/d/eOazy9GieIuUSuMCkOcjDT
qrXJqxZWLDtwFyovtUC+OTj84K/7Lc/1bD4IGEOYGqo+E3kPJmQwdiaYPNVQcf04
Z6daEPDV8Fvw6N0Fmj6XAgx495ZF9VDXLhj3N1vCiCshTWhz2EqTCFlsk+6KyTLT
rfKuiaTK3NinZjiE60WtUmNOkegS78WkKOJeLS+pR24cWJGEHgsztYRWKc//bypG
5dHWh45EeTkG0P4AfhYbnJLGu9ktruwv5HACZ5q17d2Mc/avPhNPxhl0NTrhgIlp
MMM5kUAts1bnGQ3XhtKVJZtTmsw0CKHEb10z2QagQ0a9/+FLFUpH7vSm+YYrqwTM
zNt1jkX9dwGb4Z3x9Z7a169DY5cV7xaJGC0Mx9OU4TVvZ32/4jYg6Ib8OXjVmYpC
dhSf9ttbJS4K6GqeUGCX+CM6o1tQAbR3gKYjQPSzMxpSEYjsx8nEUd/9Tvmzy1n/
cC7gI2gF7hHOW/fzNfohaNZLksHczE59PZQZwStYaNoVgGSg860BBNxY4YHcSEFS
dTsse7xaLmQ9ZILU4X+DKycZt6eNbEVctQTCALZgWr517nVE8ZOXygISyftneIeE
98A7Cey0oo0+DqZQQXxdHh1jLlzlr3Dmehiw+AtJlZeCxYVR8fAmTyz3EefuCynp
F3rEtnLjF7ivWTgfTDJL+/tcRST9RD65nc5QIjTyVB/jeJ50UtQDfq0DgR6IQqdM
EeunY08r+G+a54tK07i42KxBt3B1ItUiuqPmipXhTlw7wp6WNx9rYcfVVWT0GeTJ
bPqM6D2SFpCAtDK1DpgpDzdMO27O2agS/qPMiAcGILjD5RK0Z10x04prBSsJsQ1E
xYZJMHiTIRhJ8Sfgl/4iMJ4PQknKvtSnOA1POA/0Noth9Tm4QsAUJu/QrWf+c/HU
xm4Mp3olSXgNvsjpQG3X+KZtJp/vCqiNEYU7dRudKFh0RoKfKG07K/HQzxQRZSNz
jSwXLlgSbcO6Q255gC2H5SccTeiJx1Hk9exktwJpQktHh4JZUvkWaSuDC0hEqtYH
Tu4dBNX7BEakENNLKv5NZXgyNpOppnlIgljk3s7yt6W4OvMOUVrR7s1NQGNQOnYZ
jon6y+BW92vP7TGHO/ECz3Hu9m9U5OQQgrO6xBPdTvTq0A+87l/050qwKV+8FOQK
b55gMYvF7yjJaoBXQK2cHC+UxnRTKocehQYL56LZ3iiQAJxJDp04bFu4gIp9vpFz
Kkzf5k7xJiKtR8XsbZMD1ksbcNSvJR0xVotbi87boPcGuB/nA7vyKjrzIawaYyBR
onZcJRFJ4RuhYLFeAg/lIBAphgqdNDyDIZOoBKlg6P+OOClu2645d+/SJleC1Cdx
LHH7zSAbGMMSRhHSNsTKzmiI8qVCcAVBCgFf6sy+2A2fxarB15Ix70j3VNVBFlBV
7ZtSUWtaq3Wuagd2KzKSN5GdUdGGp0DgBczxakzq/ffiTw1bQzBat9Q9LnzK/kSt
dOR2erwyF1PBSMm0E7ApHahtC1w4lqoGkPO7/ctF4UxoZJ2XgW9EA20aRjZYT8b2
d29hcSNP+4KEhzsrfq4Gd/pBob3b8iaotkn4uxt/6gL2+lZdz+sTr1xLy2MCOW3B
Y5jOA89mx3KP+/PbMYLfH9+0XJk88wJAJTe9qzqzI/Tx63fKdSFqHnbXalB47s4e
ZXME5AL8B5HRXhDOAsINm4Rxud4cULgjr334hByWKoEzBbymSX4qPImhkTXvOpEr
9J4B8+TnzqLaFALP3OxxHf6WpnKtmoHZyKGFmzZn6Z4vrojmy41y7gv/n5RlGFqc
2MF3WHpm/MO96lQMIgO+UtqOXdzqHawasNGZfhO+Co4hXKo8vWEnfr6AY6HwdlWL
osUlAnPgBE0FkDDksqAYfXIHPGtGSW2X+muDQOVRn+Q6yqZoBC+XkJrJqm3dZgl6
5CsJHdp7uYaheHcAjcRrn+pEVp749Y8ylxHE5rJgMQw6AahK+eZvYUZCc80lK9u5
GcI/kLy/WSaqgwWd/Uo0WpnZ+aDw+nES1lcR9rmz/7NPEzHu5ov1jOB4jOgGF/LA
JIZ2RCgfLPqmMy73/D5Kt3wJ7OkvbiSWOm1xxTvx1wWYo+qLtrqxYJbBtECg0uBM
imaK3n1fCpTdxpcK5+xCbBi7jwU14R9art+sizWAH/jKfeknk5647XGwKQ1aT/7q
vcKxx8/G0uKBna7w4trt70Phbw0EcbcGs2kNBWSaDUQPDWQfsRot0InG9nxjks1x
yXXuA0sYtqv3o4E0TlypyhJn0S2DSJ+G0LT6LYKI6YhQ00UVhedLT1nquZnnaniH
PwGjc9vvioXjxbESq4rs83YMbbeYfgMqVo9AZ8ohP6LioKJAtTE++LtxGKtkkmij
0Y7AJASJvUJ5lwqR/O4hfW7+5PqlhHHkBF3znYXP7T3ERAr7s4o9IEVW4PA/Dtev
dJCdOPQK4fxf3lEJgAfaxeNTo9bpilcikOPRmAXIWvXwfp/66QZkMnZ0TnmawRj9
lA3p+KMs0SXNs5/OAEbCjaUgBSwxCE6UastOhgHqaGLZ0rhdWg5mfsVFvkMWNBvk
WmYjkrmaowfNpH95wVzDuCxVjNP9BAq27H3LVFToWto4Tu9pDyYJPwN3/niS6oob
ivdARB/IF538D830LNtIu4cwSB1jJqyiXJTALx63o4zeb1GcA/RwfPZd6Z4zMbAk
5K6fhZBjdIiYQLi+qqqeJlKXo8nMYPFVbAnCzcFFWbUgSvNe+8FOkNRxe2uIx8ss
K5LQQSCsqNMC2LICSTjoXnSbtsDVW8eNoy/sBX+fEoHrPTsl9c1oBdqKGNcfa7h3
GGtir4+ORwc6lu4ZGjN7NcCdduyv6MGmgK5fzXEcuhJHhPg9h0VuCSQg1mNluxr3
r4WZoZvR21JCyqk6KBhPaYpzIXtgLI6fwLXaR65lJiMbEo0IydlnkOCy4+ZzjWKm
bXRz35gGU8Jc6N9s4qMdVl2t4u85PZzbKohzEREI4krid0GVbHKI4kqNKje13Qo9
DE6YJk6RwNkbze++l+254ZMfHI9gNKMoc3iuHunFW5UYZPTzAvVP9hDuO72PrRWZ
WB4RklCFdtdz7/5COe7bBel/NQR9CHyjRguI8iv8gGYj7A9MKIo3wzUzcpiC+8Bk
1zofduIdNDAfQ07+DJaW/lIP/L/nelM6Q97Y+OLt0x39Pba/77DSRBOrY8Hy3/gk
WZc2tQM7AQvl9xV3srkBC9nseME+hZKdAZK1QkXnV8/u1Ela2zYuz40MnduSxydm
/vgoqrVjOO765r/xVWxqAbZoKkaCYKyifsOyH5VfGWRVmpz35gyYDJ8ISZcBD/Ob
pm2Ay8qkPhZnAo4ddavifxTjhLT/JRyzzPQirwX8XQkqONDpeDwT8G/68dCIRI5v
Mrw4GDWkZEor4oYSWwoSoi3XryuByw5YOEUSwXCFSDeP7bBf+pTo2E4HKODAk2KD
GeSbRYYkzhTalawNhngok2J2PtyUOn4DKH6427ZWlLel7nPj/v8VppOEg2k8WJlc
RPVEFEn4cqP9GU1EUGQPP+QdTZpzzibTe4ckmOJPKntEyqr/eBrZ+VEZHmuRLyk4
coZ4bzLFpV85MjDqey4C9hmbCXSL6I9KeNLhbHW+JVsZjn8gyEY1+gMNSR6DxMUh
S6SeNO6H2gWyneVss0/lR0YL1VDnLzB1hME1vfhyYDBbu385QxckoAqmRcYU15vy
fqrh85EuAIC2fwVD3jS0Hr0I/6AcB+QmDRIdZpftReQ7bHc9aJVYCzJFeP7Nadxl
w8XFuGh4FRU7iUdj/vMq8/uu+aJWIJs4r1/ui+msxt/fnUtlP6lKhq3nhVKndeBY
MfiIX/0BwaY4PgHzgV9UlPhn3NoWK1tMaLZyJdaX2A3w43EXSBFqgp70SK3NfvCD
K4QDhzVkwSJ8XC1YL1nf+wi7JREx/8uBOZGaLzSK2TY7fKYNbGsXGMxRFENYIg5d
Gzk1V+wXzfhcP1hGJqa+GiLfcVojdaXBaiY/OidfAwgr8o+tbG0e9rLWvOMg4fqV
XaOzrlKGYXp5h0ZyrfxAo5lHahjV5CJSn810lB1SyUZSqFOLgnsqU/MZi3YllbRV
vm9I56mmkACsGu9UWVh3rlBOb+o7UeQWnrOVoe/VloK7tT/nPwGLBYIbwXy2Fl+8
b8vqxq3ZYZOHS5N3yaBmyENaHzkIDYg3URt+pBlaU1vzWA4I+D5vWDtgsGBIOjXC
aqEpMqAZrEO/JV4U+fi1JCb0ZjQswt3B4/NmowLkl1xMTK6yLTswFVAYhh/wFe9O
n4440oCXZJtAkjuwfvHM/Pq4VDL7UU9Cf6HUzQwZeHgJ96cTQVOWBcLkFKw2s+ja
oyxNMYH40iR0koedQzlssC7zpBTevnyDfo+H9VtJrIUN5v+aDGToDwTxO3uQbt7U
zkC1ZZunNcD5th47XjMgYI6VbNCo8f/4wURtaZod81m7OBgZ06bQ/OFVhqmW1CiZ
a5eUYErJ4veegRKJchcLENBLj+BhWrtE+KtfbGmugOAsukSAp4K9sbHdVFsGfkz4
P7JBkl/sv2E1Bn6AmSWys5/dflb12uA/9U6PTWpZ2k5EMmHTorPknEnB5xJx3Ro+
vbBiH3R6OrbYQ4FYwiIlGjje1J5gRkHF8YVH5xyH8Fxk076FHC+/+Fz1PJcodpjN
WaAubNawDXZB05nWJbNE9riAH6YVbGDaIlv2OSH6VkEcOcdqTiQpeHFD7QRRg4OB
9DXLiwLdzWG06XERNIbinCop4hE9Jn52uxN6atM0gU0o3h6IuvBS2lC5pgYo9gkA
FB7fbmulU4novtoeIEYUHA/Rvet+UB4XQ3andl6hXRTFvrRRYmSDKaPP9YyU2HAJ
FhI8fxincrI8/0Tnd0WoKtPkBo2ohdhmqqGOMkb+zChqsn5CrcjmTiAYKYEWwLuZ
VobIouRLlrqTV6xAC50bP1tcrWOt5DUOZcfvjzSN0rCxkJKQgr9PPMIZjCXUMD0o
B/V9X1QpvufUOoMQBBqFSog7mlX3VrQsbfr7JjgGKOCbbeUO8q2R2mQlN5cbgONP
gqOY2pybbsj112I4GVNb3Y6TRBfaeu8cTEMu+ZfsbR+dMy3mQp4aKZMokN/IOYIQ
GXaP4wPCBhWpFm5Y+1JNJ33dtKSYDteB8UdoD5tJAXERQGif9Fw1DWBkIDLuLwg3
e5wtIoNBEJKPyWoiO+chvGuEfXQqn+bobXoWc2p8+MmRXYM/t6f/O3zFM0aBTmGG
aKB8LZYkPWfC2CmZ5ILTmHA4KSHyWnvzaBfliLg2DyLL9SRDrkevAJ7E1v1T9VNA
JTSEE07lqVvAzyClrlkjJ4SoT8INxc4uOihM3GyA/VGvDZ+Ufstxbc38SdA7tMYG
3shhxptGlZkjFVaYAhIr2gfT69cDMUeUyqnhk9+BZhEgdTpAJhwni3BuKDlco6l6
ZOL2Kdh/drdtxuAReym52lrkvsx+NkAHQSTwYrI1c8lJhjXL9EtGe7JD+OjxWn0Z
TUQdQmHvmZowvCqh7jy6QQFja9aXLouQh8x17oXn77CdcAp2R19WHw09gpi97HaX
/WFGAL24TYw2HePy6Uq9zioFzAhido3ck+cLjdAGiSwIM6obM+yt4srcbs3hx1nQ
YbFkBYZB8T0mxdoUiCUR7m4BiVCNOfyYoTHjssVKNOgUeTCI29bq/CPUUBtkmft6
CaBFKTRvGlJ4e8UJ1Wi1l9dn6FJa7pqyOdhIGAA8csEu5e3+vYmyrLRCpDd0HHz3
BtB5ICKeI2dxkcVsFClSkSGQpIUL/qGBdhkggr3hU6uPIBnCPmp4//XtdWWKOADX
yTGU1oyvlncR4kdZzrNZgPgSWw9dp2N/gbJw/M1UQM9JoPGVigwAhEDTjx6D5EhG
6tV6b0pUvWBctrvddNo2uWm/kfawqsb+EnJDViyyCNqs0eVZ7OAj+T9KocxEYMqG
W4SdVFJ1Ief0SfYa115GFvWw5OnMeOTXX/dnrI8g7GWbMqTQZ9Cl8DCTcKnASNCi
ZSlvzw/uKGTpN94fyiX3uqQgrN1b3Cv+x+Yn9mmwxrPzH1udfhgjwV1a4pjc7ZRx
d40H7NmVmsyC/4kmianVL/m8sOvyxV/b5dosOmAbiyOravd9pUOpKJGwC152FZ/T
DRfoHKDE0GbF0Z6Kbj8avYCOwSlxw9qmGN3vqHxvZuST8wZtD4uSEOmbpFiwKue3
qQzTJ1BI0b8UMcrxi6fbp4HeMs0XUdWRc1EGraSP9kDHV3o46OzBcNjqUabFtUPd
TkrGLymrYR6mtJWlS+tfxf8WzB+2433jGUrIluN+qS64urMy+N5aSeld7gF0snTZ
+pSG75nka6Qru2FYSK6gFGTXfW++B66orAXWMdyjb13sMjzLhQZ0AZq0poCAltXn
HxmAoqK8i3mpCVTcGf1yIn0FyfwptlzpBmmBQh7PFxdrMchzseLmK5thAVAIthcw
PEShzJLvfBnkg2LNc8oB7yEB2yyf/NahL1vjAJpuxkF9xbBbLpJzTchmQESCWBjg
Gmex5e1tRMu0uRqW7Kgs8LsocHw3wuX22lReSR1WXxsXcIC7hth+ja5/Yqz5kwfC
9bxlOGVJeD6PgBg4leNLXtTUDCIv5EDNhPT9BDArB22OQGQgCkxAa9YrSyqzZLHV
CE4xYDFAf7wd1TGOZ3fG5k6KeHN/n7SeoivPOH0W0wfcb/TvVZNXXzHhSNSDmegf
57YLIZOAv2J7U+JNHE8JIHcM7KlYYcaw3Al33TK1El02jJi8jsW1OIksnsrx35nc
J3xjUl1z0qCn0rKVhs3l41Yjpn++N9xWYxKRl4fvw1BWgc0lJTsCQ27rcsGDKUF3
4cslGXs5Ola1wrpiOT8Sf7lLBDkpowWvrIhRyDDTu76kvvGphEQK2ijkg3aCVJ1F
oblHCGWibw6OTDMtta1PPIHdS9rjIvGXp5ahsl1E4cwDWbiT6u41W0iAj8ca8ZAb
MD2iHHTXajaUczglu8sM/fUvsbCu8ghMOw46zfZRO4BJHbAjjIE+HT4MWMg1waRl
uWXBTgCWgmYfebWBHlNcw1vmG3PC7+t3JWCIVEMhePVOjDoAO3FUDipVg6fmtRmK
5J4beP/zSTBxdorUXHoBPoL3BSuRj/xt4kgjGgroPNlb2dncH2N2OIZzVDmQNVCI
XIBEEepWegis/GaX0GMqVEDDlHLA9zyUyy9pfAzrx0sFS4ii/gt06WYkiX2+H47R
xCAwAa4XgPMwZp4Me+8QTILB5b5XDeXDm5y7P63o89aj/jBsNQZGgKYlQ/peS2H9
fgDj4CEII+HUc53MFY4SqEEIjSGjy4yc+ipns/5UAliy5NhSvwKKlBfyNotbwMCL
Yjvd7+lTP3/Ikt9s3eJC4Wk/Iy79qv0kLfFUF/hURVysUzgM3swxgCCaeNGVrHRG
KBCeJ4qI1SnmF3knSG5x6yLn9MimbdQKxOt1EamXQ7sNOtSRSqw5Fu/K4u7Cs6Kk
yhcm0ylupDsvyOxLY1KKhNRM7hDoKMEVgCE+mstmB1EuFgWHmoJJ/RxOOPttVzs5
GwOxhIU8QT51D7abcREN+DeK3oeeA6gii1bJizBGCxLtA1zU0e0ZT/bvsb/EeZ1J
npOpTAshgSlzxfXmLUz4aI0/+Q30ba4E+3+j1FVAJpvquOzEu7cEfVBNCFdvDnSN
ukA7OymY6IT6ZhVqI9eLZhTmORkALeYH47nW6QQVsDs8tCCtusRJZidLZ3gMJXOH
0aonZ1QLeWjzHMjZxpZsOELeNlSzPuB74bkHry8jhKPfm24cc+KjJhf79Txi20y1
JOnlsjSX3bUh8iyvmw5AoIjx/gCBHYvv1G7jXRr2F12KOMnMSda1XtmHSEKC6Ur4
MPmX6ZafM+zONYACY2Wq1x/cRYDbfl3LOn8IJePbIf25q84h9nzafmR/b4C3M/92
5FQVx6tKxY/y6g/jrg+9H0xn9BvEergikHqiNKKPxcVhGylhS2fOIMZtF8p9hHct
QeGmJtPRInGj6ccp5jNIRxBwjX1ts3TGQFmVUZbOORl9Jazv6JSiBOeBsFBXjtbx
SUxWynHuBcVC1Kz3wmIOWYvzxlsi40Z9oe/3FszMUH375ZDz006Y2XbOZGnYOeWv
9nKpSKpm0P5ocJUZrkObOGdWwgRh81k81ckkKtPcm8JaeEKxJlmc4O+l8gpLrFXs
rN38MfYQm7Oakk/fxtBlrVBp+ECcj+Vz8wCosnKRul+Q/d6m463633fhh3Y+ueDy
3YgcNyUi1SxJtF1yNczVJPzYOzlPW4xtm2T3MW8saJ22LvxCtS2Ksfb+nghPcfdO
vVnLItZhTXoubZqIE/uZiJFA9sOYYx9bNI1UXEEaCNqf0s1jFingLuGMLJW8e0+E
UfdIE3wP8vb5UrWa6OsFBBhxHOMLa9o+D5JUzdlXW1zsAf/iKYwy5eGWyycRKyPX
XF2oBfpbt359OkhNM1aixhkWxsn4k1IgOFzpF+pbBtEUZ6zbDILF1ImiQfRD0Eeq
oAZaAslInvkaq1WD6+D4s/Z5HKX8EAptU3tpv0a8bAPAJYNod4dSYVreusHocCYN
XeTYYYQHUMKqmlVYe6Vmou23kTLojJADCcVX/WBpKcoU0PzJieKDygONrgQ/y41w
wVtnJXAKSIWJKbYaRrjm66QD8NIavBJPAlXUVe/L/8afEB10M2zmwZ2qrAQ0xz9F
xN4aspfKOUW0EHdKCtTXIgmohI2kAhSgUgKRmXUSArCjReDhayAdgZAGARye3Mka
olqn32nM2G5nxv9CY2oJItd5sgIuNuU7ItYY/E6Aw40RcTph/CfDBZopLfncgbBQ
BBQWuvsMD1S8JkSoRPsC5mJg9zAFVrdQyKZ0YtP7gcIlMEClT2XVdLgGpFWtZF4J
MbcsGUAJUPd3/u5Do7GsCW39XMMbCzbpb2bnBYhXczpxEKP5RMeyGAAhHEo4QnVY
FJrFT/DUoqHvo4O2kdry8XAvzPJvgZo7/FamD42YnsmwZQQuGSLwqyAX92HNcyAT
bM2Lt36wD2b1A3W1GwHZcs45Jn93fECZkGZZbRTxMyqTYtAEb02Gc/BIj2Mcsq1x
jvaYNP368PuP6Orztd9nmBfYDgZS4/fVZKHYPNa/rCFvVoZ3bUpFM/sKa4B4/5ml
qQ8VID5VndRHIEQuL1J5Ia1EOUr/9sWaq0h9e+pWGFl8J7qEE1YLYY3BP8fqa47/
GBs1c+ehzqFT4nYbgo3CkesujFQDp7JInS8xskiRjXWDTAjJNSINkQwawPXpxZBr
2TqZOzaN2A9MglPlIvJZYqv5gUTiKTk1r+06LG1Rf36jE6qngJF0hyr6xZ2nb4ao
KTfafPOIdbKZrQ0izASyAIbQJl2Vh53cf6P9zGO/F6+wF4w3GQWwnKWCItbgCIsA
gIEuOPPQ6mXclqbXHwtd7CW0f5fXeIum6WUfs0aKdIpcXWCZ2oXYa1RGOUu0R6yY
LHHYXDq3OvBHxr7g48zjHAovNFTkPV9bBnVWwlzTv1LbecZj029UayktsytfW96h
aRMaGvmBJRWKzrhQVUFaO5wQEQkWomQ2+7ymfjL+MIwuwxSLPh3gkp5R6oFfq0AX
vUwSR1HQEREwb2+ZGvGuIjcNB9c1/3dHn4BKTnUvMHhNLcPLVAyzU/NgdNRzNor5
lnbZaCUSV33Av/0y/XMEtUru4i5lJlmeTBVpHSvTA0Pk3K5aH+rGkDCf69FJAq/L
EvaWdADnqyeLIJ/R4rQ3EQE8Wh6p0aiRSaOXlHQ7jDk6Ktk5vDc1Ki6mLaMSBz29
SzXmAdqeXPYMk+kVSM6hlZDLHTmd2Lh4g3u0sNwfW8P+v7CJCFVGmGlBpqQuHKs+
PxSuvbs1TckG8wkDInLWNubrpi5yOvUZxTRXxFn+1rc3LDJWcZ0XiwSG1TsB9HAv
Ja2Kih/NYY3Lhq3NLucPhaZC94c9M/lZRgrOKk8vJ/n4NlDDM75/QtbGxSAurZx5
GpblV3Qs7j7mD3jzNXph994tQSe5v5TJALt0xP0tQWB3UsLh5xiEYIaI6xJOzin5
N0OFq7RxuFiaWKwyy4ubA+/DxIBdUD8ZPL9b1WWNSxS8+awPfBgZ+o9W9XAqMG6d
MHhR2ADOIHieVE/Elf3RikzmqP8Ybyi1tLPZ4RcXAxSdw8AUxzGRMSqwj0+JczWl
7pH8UA1F2IlwvyLjc2ZdMpiq3vmHfE4kdkD2XEQfWClcIA1kUIwh+Pxk64ZQez2N
75puyyfHIKS4mt71vaX5wZIJ2pJYTaJ+q9R1BxwQEvHaZSy2JtcA2nOh17486NQK
6VzroCBG+NEsEx/dsLFdmbEoiCX6fpGtbAHs8y7nW/lO0v+vkJSYmTDAgwYELyuj
xPWa+A/1+BEuopA939rUOo+xmpskCW0radhGJbt7uTEKnnq4VGARcxi3XDboMXI3
phMFYTqle5roYwjqN+++7DdUI9FXyq8Zxx3zW51J0ExVshFuydDsJjjM7aToZKYT
1ACuNl4YrMuYO8DC+fOiAednd1aT2rFR0G7FdEq6bKFDbG/u/tkF1AM5UfahoPwW
DbxyAqb2oWjAbzqsZA3K09J3NzSJIs9S/32AOcOFWWoVihTXfgBtGRHF0h7eTBPg
H1HVP4FKTszMdBPDx7i/MR0UPQHv2MHB8c6LQX5l5nUgL6Af7GuhSiaKxRwBcRti
9saYglPSqaL1btRahAhBsc/MzKEtwpUtEs/TkGKxZhe/VbdnjCb7fPuZiV3nb7Xd
4YXIrphiQ2SAt/MKQ2nLT8eRPR/TdhW7xlOGruanmqUDDfQb88ElzGBx+est4xO6
AQ4Hf621Eb5REYJdMW0d4mN/kVI8ArP3gv8v05+IlvaEK6jmpwICxDV3IeE9bZtQ
yLDialxZAyQjooy4FVfFjrfs0Zx2bHcEn1a2esBNeGzih4xbOYdwUCiuboC6hX7K
SjG4xstutEKHwaa/Ovl5Rvnj/3YvCNK2k/tRkitw9AtvRV0KblSEIoBSYt3AIKZZ
menLjFw+s+IY8L95lDlaTg1MQC1TCxNF+0yUuAgfGed2e6OMMdFoexPvLjx+Gexb
nZ/sH5cwHD85R4JUL7uULrBMjmcHzlAp5yBQOBS/l62p2bG6LfWO/2YvXMd9Bb6F
/0aNW03xX5c0jw1ZVPV86PasqBICwnbDrE9jw3/XkCjowsK/XhI7PBgTCma/O4sv
dAJ7fJmPne7M1jpg9Qk2t0CJD4e6Jd+n5rROBXlcqhZ6Tkx3RloZqEtaffHCtvf0
v3j9kz9qFiBemAKAETf0DgSYUmGMuTw+yyAZQ9BR1zvGyac/YbX30E8b1eg2GPRW
OHvbu72LtrTC7SDi17P/Vai1/vV6t6vFX27MBNgBewuRXd8ZY22zSLAvJMx82iaz
bkTxXwrd4n67Oxttx+AmHIpb1g3IX5Ilyu9sAVzZ9L9jO8GTOdMxJhBkC4DDWDtY
RZNVCNmavtBREn305bHcyftAl8FBYh2uFMqI9tGnGmhcuZodzvNoaZMoGLAJJNSZ
SS1ecafHLv7QxoYyX3wKRKYDNE02OEaaZDYSEzPUvK9dxA5yZd3deicyescvyV9t
lGbyY54eFl1XuPxOrDMWblYUZOHh5rKR6FRQtW9YSjc8bP1SuQof/zIV2Z0nRTRX
V28F7O3kmP9qRJQR9aGhbfxcBbkIMA0woef6hgcSPHe9WNkaAPoVDa17WK2YDKDh
gP08lrJ6j8zRiN9/52ua8TyodEpHA2VyJ7oMXitN03CpNscVlfM0FAT0m3Yzous6
UJXjUaJKBsAt/VUzErFYc5Qrma85fc/PA/pthyZpvt9DvxDLmmDDELRC6S+7GbSD
o9atBf88T6rWsN189/c7wkN5Dg7EYQSnisT53pXc+Osm6R/PGryHjurpQjeHdwvc
iaH+Y2eeEDCgvPo0OlZzs6t8RnvkcXlOx20W/R0kA14wYavl9HhMt6T9qMrGlT/Z
HoXr6J94yITNb/+xCbNnuLXVC/MR9lAvQ22knoCqi4aGMT55BCsXHr9d/DhyhzJV
oFsGgr0u6Z1rnn4SrthdJ6K2gXRg5ZzYBryZZDwOeyJpjVvKCEdWzDp5IRJL/nRY
R4P5DhT2U2rxfVz2xsw8wcV3fx72ws2uIxiwAOZqxszEu2Y86d6iqtmHMKoH8fuB
DqAq2YkLE8RvwKBKCAA+XaTw9NwLLxH27aEQ3eH9VFCFe/pglv9HG7IMI0hjYart
2b3tBl5iT1FYbs80xLQdbTfrNOMoqKLGx48Mew8PCLiQJhGX1JtqtbUaQA+JMBEt
L2XU87PxIzpZjPnnw5R+b1QKRA1fY1OZvlF5MwIFCW+hX2qE6BZhkS/LnELwBaxG
eScDZqAsmFwGOTfwlEVh8kcQI/nXwcwYw8SnjCMF30Cj6o7xTd8aorgHCru7AX4I
REAewW2mkqop0kdjAVcfAkTlkIryjP8X31pgoNJzueFtVdRgyzd41ZKgF5JNl8Li
ueFoW8wsr3sGaRtcvOEMu6W2vhVXDDUY2D/SbP3UswTu7vsbuqOJRt26rIHUilp0
3kMBVn6TEfI1yQkW4bQ0hP4PfILBMiYfVU9ejzg/I0dos7fNFxa1whvXft19Au3m
GWmWpIsiuyh/Wf1vDxmCEnKWtUxZM2c4d5bzEuIjh2aYg4J/2tULkpuHC5mjFwPh
bf5v6aHs75H4I/nQMAH3w1cqvZ/o52yYvUxNsXPCF20iS7wc7sEBbZhtDKdr782G
QvAcZ4ERWVElBC+f0pkuVPyZFL5dAutYCuIGAwFhDPHSuZCWEgV8gemDBa9Q0Dh2
b25CCXLQTovCMWUxO+KZeJcb7jQbvPOFUU53hKseCzpSIkqxLxhFndIQHQ9dTSG0
nqhSmyxzxKvVFFJPaAI6zyaN6U0tMWptSNq6GUtyAiPI4YoI6evKbY+FesPW6vwh
v4TKzsHsBUARx2B/As39vva6NOyFCz9iF13q29u548YIBGHSiDPmqTkNK2c+zRzE
bhMfYwn3Dcj+oUSh8x9+E5Gd1fOIOJDkH0CLPOFqRLSCXYRk3uyqIBgpCWS/a1de
egnWw6TLa7aRZQyMJfUYC/aNyav16wrdeFAnG+lotv4rIt953qy4LXWDrOKsz0oh
qIXdtLuU+GyIIxIWNhoHKZkBgVaP7YpPnimSZ0+OukKfGUAyAe6M8R9lRWtKcBRp
rvaESoRBOuQ3kvWDjUZkt7IvN3kQIj7FT0Zn9yi2o/PV6tS2tGXf0+F/UCDDBldt
RHDMjT7ueVUTYNJq07DwaFURIzScNMijhPQi8SPmeJYrVr+BbsbS2kgpzDNyETss
/sNG/Ptee4n+f7G7VerYywEUEzBeivvdh+On3FiMMfn8HvwSpjYSxwwmjeAePisR
JnrRQ8LXWpy07osup00IGd4cO49rJbt9Pz53/SagkmL2UVc8WFqLl7YGe1pZQ3Qx
QzcWX9iE/dPIurGO4HF8hhgryNCr09MyTr+TpOXK9EBM6VhV/F4WGsG6OA/lc/P/
18UBy4IsVj4Hs20XUkm54zm/A16EPWpmKTQ56cieGJQ+zmERG1Mo6sQcoR44DEht
moCmIVKeDYlm2ck0BuBr8Y2os7SvO1Uc/KUDGpBrc4Hg8m0z1grlnRxk7by+gYpl
+HC2ac12C67NnCpoP/QFvgPobgVTuD4nv64vRUbK0uiToSx+27lHgurBKdnvd6yO
EOTENkyfdOVQ3TkgmVRhHLYp54gdnO4vF/JH6ddGH6KpBMoJ12IM17144NyqJ1tJ
HKWILe2e66M8PKccU7KAlz+PmWNRil5wKLuuoeV3gN8iVfx7BvYS5LRAbY61DXmk
Wk/s38bsEOkKPNzIHIdfEwJX5wQsPUKvBfuSfxxrZmRva1M2teO6Wie6XwnpDj9z
LVAuXPshTtRBhPI4uXkkv0sliNzygVxePQQVg95rMA5a2VJEYHI/X6/JLmR/j0m9
qorKvrk63hvAzvCzGA0/eS39WEhyJkRK8/1DdaGmKxLPGaXmHCTR24alhDTr8yyc
RM0Y5hspVfw8z417a/iduSXolNwhAYPgcazT2FDav/Md5fvImeyAuVrp76Inavz+
PMejwqxhZObVyZoAyuYhzqMhdiaL0dprvSW7mpepMMm1MNCmEEGNbSeayUPIJdop
6Xva7FNSVkZgQe38/Czo3PgMKXZaiKs3BYEtEBw0voXTey0ecWgyVXkYEQWWXjWQ
Dp/6zbHCOq0pgAr15Y5YBY692428ZqwxK09c6rpLLh6yO3/LPavYiNhjMFM6IE8C
aHGfRd52V1ifpJk4c/mz36+tXYohcpEH1qXJ2iEUofp6QDhMBMIc+U5MR3Yrfsop
poFiRqMETnPAaUiA0EX5JGoOmMtnZ3xlPECUhdM61yu7I0NqLQmv/fGGQT1CqsXG
nxo0k3gxKQVL+//hV4deDRlh7zYjt5IMfCCxMwUwFMMYoM0zvQ+CGrOWzC2CilIG
IWh7qJIzvdTROolqw2CFVS+xhrF3rFXP9Tl9+w/8i9v7zuwjmFhgRRxDRZB4Qomm
0pyWkz0vFuODXVREPNAxvArc2CGORt+7IxEpd0u9CCVcEi1N+lkv5tgW1HojWAYE
pwVHeF8ASE3bJu7fM+CLmuPNvq4zXL0gem35U6DX4/MfbU3X+JdNV00lDgTb0m/K
DhyZIFKAhin+nTnixIi4cqjg67jYsVW/kwGFlAZHct73rEX4oHwWxOSXM3eFBmQr
+o9dwuTUxhDF3ChAHLaPWxCZOVlvu+CIAUV2Bo2PT86rWjrG4t3ehpjByLKt+CzU
Af/G7TYO0sDQMXI/eOwLpsjQ1UK9l+heYVcT8jB8V+1oJLg6S17oNL7IkvPGLAjr
YTxvBO5ysUtIXpTBhnltztBWLc+hvAbrqzuEB9HJ/r6OwmaSfsr3IhjgmVPDZ8Wq
5IfFxLOIETT425VadbG+01l7gkWlRF8YPDwIjmKwNdZyDLf4JLZnBjwKQCGhJMn4
8QQIOzu11LwgqeJL6ebObUDA3dM+lDzZaeTzLdKpZ43syAEcmpK7dEGK2WilEsKr
lkq22XhfIzKklmSvnhuciiEhWBU+KrcPXKUEHxDXGW4R1o2nf605bJo1GyyBhWuX
18qryyyiYNxH8R200+QhN88GpR8gUdrn8nINTXJgMpwrbjJWXBDWP/qu28dpf8Qu
7qAlw1U1gpbXbkVLO/qSHTEipa8sK2Oz54XM91QkKgzqOdHXSr+pemR3tQ2I0FoQ
a7jBRjOZFJrBxgS0cLjrrs/RNZgdak0Gnl8wxKtNzjRIklCttfJDVKHby/vofJrw
p8n0QM1vBscwJGlslbpwjNnnrbS4kPN/bJOOKfeP6C9im6T55CRVfOj7BPo7PkqT
+clcIRKpdmAEJZtqrAQs08Z2J2FVpFeGBnfTK9MP/popkZ2M9nGOb2/DG9v6mmqK
JoXvVDs/+fW7HPEO4bP3oKTmpY3yAt05d8jTaXAlZPZUY3WLPU+7YvD6X7i+V6OP
ownR1GL01uDomH9V8gTIxAKcoNcY9E+MttuDfuiU3X+TVy22TBjOAbOs75VA1Va6
km639fgVtvbbO27sSIATL7iidH4wmijI/Y7T/hUcDul3lYwTqAohl3lSf44ICkhg
UQbbk09dt5uCrUhH0qJRvwTHSqJIccVRBDcq+giEUbI87KK0V2Qz6gsmo7wIyWNl
T1nl2LdPRHv7kG9cfbQoMAfHFRFQjvXxcRPYBEVu37B9X9kZ+6Ewudius/u02qGS
pf+KhWGMTFXtcAO6+uRLEySXxDPQ/h5K7tUEec08PCABm1gDYuZViaDlsOv7Rgfx
k+YtUSfOQTsqOaiP1S2PDG6HALRDDOA9+BakQC0nRMyHDWhwPz5G/Sdz2S4YNhvK
w+vKZHfU6HpfYnjmkJcZWr/sSaWtAaYlEr7DBMKxx9mKDqrbHC4hVaUkRNMNEJyo
3Zy2jFXBklO4myGaX3g9Yoxhz8dXyXdlAby2mNtc4muKxuB8uf9bvjEK/JDHtS3D
ZbEt6XtRtg1ynS7ChDCblrkuJXMKH44cfZD0PvUZkT1cobQfetpah9hl9kYkf141
x6guVAYzCmgFlye6DfRO/uVtxewlNwCN7PGaKE7n0C2WNwMU7t4v39wgl2M9+SFu
MmPGGFEb40UzfuZCy5FYgW4ouJXcQw4frGg6SKO8xTdKYjzFZbhwbqUAQ634/jO5
8MXpXWFFwNPSB7mNR2XyNCu+N1HdtVTZiQ/RYQmKnqhS/uNqMiF/KScMFpQ0/XKM
ZH/yB1nthofxTXcfoxd1scTMiXCSDld9kxTyIQXrzWoCd/zDHf5lRKA6YBdDzQkW
d1ywvzvJr27uxrA228PDlvoIk4wyfIw/XLQxxPKufRSU4ZBGl0pC2tLhqm2moZfj
2lfEm/OtQ9SaX2iiktZ+JRlNwphtKyQQAcspXIaZI4G+icfvcv3z2LoiFgfmobgz
t26t1PNlDJ6neEe/MnyndKPCSd71aPm1zPTqVFYuTRCFzwXotNkjLBMjgb89tSNY
ZIMOx+ynzuomBbxjEZY5HElWAz85ZPUOYXf1ydB6honZ4OBGqgQ3JZoAZqONao3/
wt/ReeRQRhjCvh0WxSuG2sPFPobfie55zXJzWW45wlo5DqQH9M/+ACuy0AEdolH3
yW1qqFayGUm++t4G4kKv1TjdYK6WgiZB5sDZ6u+RKdAGQjlf0vQX0RPRU12Hhfwe
SYzS4EnBWUjCtZkRzGvi6sEFIw1Qr6xEeGON+OAWkPGCfhta1wc93Da39/yYAXwH
ibPTm2Hdvt4PdV7x+oY5z7cJHQKZdT6jP9jzK2K4PEIm6Hg6peYT+yrTP0Eqd6bl
hQUwUCDrrDbBpYj9zrQi/g2pD3IEieXucHl68M6f9AjhVVFa5xBUNWDRe5siqX/r
VHFq/7bCC8NGv0s6d/5ue9yIBnNCNmXpQaiUddgI2wFlRjctph2ab/b2fWiL/YC/
W/D8WIV7UWRleLoMWMspgoT0811iB7IZBMNxJVNxcbTq2t9/nfBE7cWkdiD9L3pu
KFJh16djuS4qWHqnW98abR9TXPlHAL+OvNMnFGM2vLZOcgPop/0NcFhpqha2KUdF
7LC0soxtEeTUz5yTaw1K0znFxiZaSwZ0E9YUTDZydUV7ynHqhOHda1j4N/lLN+3N
VbGIF61dVvuIlsc0ZtljSQArf7JsblvnObNJSwaYN7R15IBKiU70fXrYkwjcu6/4
ZROfUExwMaA3exsXbSP+LXZfM1supphPyScHP34I1kfZX+JBKBLXcZF9Xd79gIkX
LFzxwaPFfNTXFrtK4wGHg9c6hHzX0akpgDpuheD+fCDvrNqJerNi7vtRD1pPxuZC
EL9IfXaciC4kS9kmCt7Dx/h2Mqs7zLKNktIJJlr9n0PcjTmyOlOkaLFYbywRfS4d
WxMvs74Wgc3KOdIG6ED1hD7/mRD+dGMTX2w20tY2cexKazuFQhaqaaGLkyv8tT4X
V61/TnAOP/+nSpRhSeEjd4Y5OzEftxgN3WUXXefVQyKz9wrr/5lClrOBJV+522HE
cM1/X3mfGnDTHaR28oC9+8tUNC0GVMOECeutBAYPMTjakPScY061tHYqTp4u2Nqp
FY9TwLxhWPStn4GUoeNyh7NkA/Oi8JkDkxiWG2/lNC3iBXX+Vy42gn/yE+BpH+56
W3Ll7AnoX9zBmqHy2ZKuS/VH46Zb7Mpq9V2407lYXVd57QZidvhhuH/XbnNNfjDs
0t2xB2f/lZdy1I/FS+WD3VjgFFW1y7NMm8ImWPWLO7dQ1NHDGn+3m+dBUKEjL3Qo
VNXply+2cGdRTjYI/T8kciwkVxUkRjGX1yUP8mrlIY4o46+nqPAKH3mxtGDQARy1
Fwbezr85lHT3/RwcQ3AhnVsieBpXIUEWjO66O2hkW+XxfzvOnztp0oXs1nts2EI7
KQUSFCVSzNDCuojkAHQFmld3sV3ux8VfKM3gDeu2ZqZbX9nhlPB0RuLGdDn2u9AV
09av0gM2XSa9nNcLHsLzezqawVBPVnhPQxHhav36OkIO+SF/P2Fxs+rQmdARvvZX
XFUAUmZe4fB1MRV0s0FgRfSLRbA3CuwTkUOnz2U3EbH5u9Hyvw2+cej+IgxChDul
Eltmi/JyZB77hI/MFDUkCrF4fwJZ3fNr0dJj7c0ywDGqRDCLd+dqovJcp/Zj9bpD
Bk02qsRiAG3fkzLHLnLoQAUS7NMYZIw2Pvkv2oB4TeqZJob2bCCl2n1OWHWi7dcu
C/TmD3I2DthwWDujxifTaj2Zfbu1AbiMVCPDRSLLhLpNCJF+AEc1hYQWO43Xh/c9
rbX5mWPrcMXI2UPy6PFX9Mm738bRZahRPxpkTuJtAicR0KiXoiN4wdfb4p255K0r
9TDvSKjr6F3n4ledaySRSULgaHKratYR0razHld3TXOHWSyLn04vSik0QtkCwsPO
2zssJoR9YxDivxoCqFJ2WMjE4+ZzQbmOyRBxXsEdYD0nPj6Fff96sw/2HZSURUw1
5uIRV2ovxpqOVGB1nOUS887dStaANBzwz8eNpA42XrsKvhx+fKVRddcwThv8STYg
gOCeS2lUinjb8NGdcQVFwg+BkiY7VDfsIYw/6wr2osQqaDUuRjuq+oxNiKh28yOb
rcpYvbWvjL7flN9CR8u+anG1a3bIB7PkcppKSoOM3BkdCaRJQcFJ2govX+Uyvbif
FMPHQD5PNGOkz6Ue//+pvVnvgd2yuX4QgnPx6KEJOy56gqjIiP+9IpXYnNhINF0h
5ghGBh2LaZHeweBl2nnbk9CCqitnwuVPBT54Ge8RE73mKJFvlK4dXV6RmyzsOBl7
Wu7aNsTTN1ERQD75nHxeVZqJHPYsN6H/orKCbo2iXyJRfQf2XhIp6zSEjszit2V7
txU0zqG2xRZgVwUWap9C1y7o6kNaepEhW9XOeUeYTsTzHP4zajcNVDVcZbUmcYJ3
baEBfNTYlpTa1KsxzFxp8JmK+LkinMFIy2IUmNh6lEa06DgwwgBfMzqRg/elwoxB
8PXjsXf/kn63t+RMNK0/lxAH0UWe0NBWT6ArUTJK1Rb33se6YAUa7DL4Vz96uUCP
htUJT+rVnfWAfJLqdgz1GG3YLdXa/jpjAilncXA3U2LyitCgjdsdLow1nKhPvfqy
vFgQVBS/rBSG7KbFehxn0yeqjJ5YoNT54jLqus2dBWBBvwtZVwuYM9mwofoXVyU0
6VBd+EpgX6x2eDJd371G1KtM79UFWc6kHs5XmweK8UVcZ5RPSNK973dbEDW5dbIc
CCWIr4GBeNJOYJm3h0u9dv9Vm13E9Kt1MwxMB9iEhbEFUbV9wu8+BReKZrfEDqCJ
Ar9Lya9BErCxxfQSB7WTuVN5lqNnuHXwAMWQXe0+rG2BC46ksxdYJ3OykgBCdD4F
GBO1drzQ0RrK5t/WNhAK/n6mmfTS6nIYGS4oCnwuwefPsk6qE1f6f4kdPA9cwScp
kYsTW9LEuAenJ0X741vER49bA37PLL2lkqFDwTFmRdu7JXfT3bLK2fU7Ff3WJdn/
LxxzYWY3HVzTYy+yDT0mC6cdpLltDy/qli3J0DjIaOQ0NU4H6hT63seiznWPVelR
+ffA8rwddFhLRWEiscVCvlEFOq8ym6KUT2HNPwTWVAIWuYUg5xZjGwmFH5WxxAty
or1Yz4xDI1RyMxLeNQ1dA6FzZtjGVxAeVRr6f8zVGflUJgt73IM3JEmXnR9e2/hC
wQtVqaXbY0VccP/lII2h6GYVdftTFTgfBoNJXZ88xNzcaRpq6Qy6xHe8vmeHdzff
FS4liRrSHCDZ0xu4dhsqCtJVEi09s1sK5fJQ9vSGlEp/jInKEsKWJCMtA5fzxnb9
K38+3j1tUY0PAxx1PjRIVXm71XdSE37Oj+A8MXxBoAw3vYQnNgLkRwxdF2ok2plO
ZJgytD2ZTThk/q50OGEMi6i105/APZg7sEVGY7Ru9Ph7X91rEeBb+LyG0gz2Dcrl
MvhVaPRIHL7qcQr6Fp2hbYD+5WN9n8rzMw1WZP92vD8aL73nguNQ0HdJDnLge7iU
kuIkKHGcNCXlqDCxXlC6IuUqjBayLxOD6oTlaKNk60eMKF7/z4KikRJ7elVeeexh
UZJutHMklxje9cyidRz4szpMFnZk2cTm0lFnFvQSygKXN63AMp8gW31F7ie9+gZ8
07JG7vS33lpo2YxIxdjK+SbnDLu81glgfTyCQu6Lkh13MxH2pKc/NcSEx9fKipfg
hmy2d8oEap4Bksf9F8T33JNer23lyuOs7M6TNGmbk6WFNF9xFS4EGxUCD+wrgyyh
IroEhMTSLBMNZN69dRT4sFX0gDeFu8ftc4eA5xMWUp3yNp4tMXGyW91aok62+dX6
oU51bnMLv5sF3HOLbmbnKEZvXxxVJZTKU9sq/GkPINEUc/gM6uPONFTV+IPz/Cmk
5uu3ND2Lhz+llES6lIEJyhSTsz4Gm46M8yiUMHKKdEOaeTjDM6kVeSbpBewjQLbZ
iYNNk6rzx6b0TZHSNEhQ5vPwyRdVRDDuBJ6R1QTwQMGGtTN58jiyNJFCf7FhDFq2
LD+MW5hlIS2IcQ9Rt/gJ19giGrQsgX1Oo0+0PEv2541umGo/ZdCPg14sAnBAc5Mt
3m4lXx6xkY17j0QepMFi9CxIiSgLHKpi9toW/WeIP5/zTYE1osRYKePzJIRk7Qxj
pHWnCayDY8eV2fMUh+wE/Lu00laNf71rE/5jHmFAHYTDgdHVxfb1tViviQp/Ec01
DRQsVHeC6SkA3tSYU2VMvExkZXpIbszW7+Ei83HEza/HZQJgD9UBt8uh0SwhyXTv
GRq8nT1Xl7PlzMLoGoX4ehZtWQHslIpnNrTtUQhkN2d2KlA3/yrQH45HgMTsDqRZ
pp5edq0aK8kP80PRqLpUuXmVSEkn5GZ7bKBXRc/r+G3vwp+4+meEEKjpXAhPVPv3
1jVE40xfyAKeKgk8CsqMt19iQ4D2a1LFjhWK56cx2A1Sdv/GumJ8N2knH1dP8PpV
KdbuTiRARkWXd/bx68fkjl7CqqyFez76AjFosprY6ZAf2m6kyHEQxpd+iXVvPLWZ
SkGl1jufSA0JD3sc8pvDCR4YtAtY6wJk6OzLzBQf521SB3HAKmRtQamqy4PGWCcf
zlo58j0o9VDXdxJzux9J/uqWoL57N4GoQQUQY1MjPzC9jWDsbcP4eKAy0UA49p1T
IX5hA97FoRke+xjpgvR2vEGrpSAYDnrtpWUFzSU/Nrd/qa9JRbORxlInwuroFIIj
xDKDlFT95k5TKzpiieUsLm0Dbwt2wamNqHv39TYdO7WTYNsmo05YZ/wK+JWfkCcD
Rbqb3aDL/GDxFtCmScukiMMdzEZBQeAKkOFL97jUqMYGq2DDPLa26crz0l5GJgtG
V9iIuQZ0X6YTh43W4GXzTItP3f9j2BjRZRMjTxn4qhJuBtvHvk3KYvfyvW0bSdCu
Kntmawam/8kZlIfL3EVFavy6OMdPCNXp+h2MumjjFVwvn3Mnca0NdKW+9cpHbtE4
qWgh/cIsz7qOlUsBxazqmA2hB8uwvQ8myEbXCFndWwIBJeaEYU4I8hbKNQuoowEc
b3+crBm9CLeeXsYEmgajvTpY49KHlDKLnCj8NbO05PD76T2KqbWu/3NOEG2MPKqm
i6pyKvRCAqI3+dlKsF4Jj7SntAg4LKVB8xsFQ00+riWgGHlI3JVskAsVI8akfyt/
ZxZhFVLxcdEJzmWEtFy4H0f1SwLUIg5siKu+VDVP/6mIHvMV/+03lli8+T56/CpO
3dZqmvMpNT2NVptA3ydlPLJ+4KtkYMIK9QfV/eXphrxGp38D/vFfvlWxGSF/e+x5
WEgcH/75EvIlDWbsBg/TBWkvlG2AWF0hIZvclijGx77ILYQfu6j12+hxoPj7sPoS
45xMt1IT70i8tbrwJiRCU8fjWL/GFA8QWAUyUAUE7o6hzM3yjnez0PaE0WkS+Vul
WWXqvwhXJlSrkKDZTZPwlwrZ4ayR2iacfgWkQ6wNV3YGnMDwL7//RxAtX5GGHQmt
4vqQuTQxusetl/gdRqafWZQ6dMWtqrkUoQP5ybvbsrT8okoY7sZp4Qbqv5Ms0/W0
udfI7zIlvMnZcAreKNaGycPYz3F8Ff1tTAoxBDJhSyIlkBT9Q+0HmmcPkXOzjZkl
13N9J5JUFFUsRMsg3xErmugvBF9PyWaANI9YAGoi360i3nPEBAz+FAa2vre50k4C
wNkJ9v9tzdTyQkmNF036heKdC/NyFkSQwJf95m33+yB9ePCKVC9QR9ofhsPd0Kyt
cCE8KZK5/BdM+eAzlLcWrbylYgVXVK1vmDJMdUN1k2DN5A9Fgdu1M68wfXOgkX8t
/H3O4p51oOdTbWYI2KWasunahLnSxNHBP7K+ScXO78a48m3Sycvu+D6r3VqMKebd
k90h3wmDsXRW4G+3/1JrKecitx4c5O0jcePA5+//Se3/sB1RVNvdC/tLDGsjDU8r
RnwtGFa7UUEsfFR907loGRy2nEEqACpdlE8ABJvfKHZyzZVLzm0K8Gve+qBkqvDX
MGnRaNqJ/nuaxcYjhaciCcxTCYFc+xMSHMVCUFkf26teVG6h2hhFruo+uw18fMzw
NgHN7JZlPQUGfUOJjTV6ZXoNvs81NOIH2gIz3sB3hoOwEWDf/RxlLktAgAeM0EX7
N7mOXHgyCT+jmuDei20Jo69vv0nx3Pu/blZl2jpJ55S4RfztsjfDCooL7mkXomqv
tmPaxFEys3+GL8eJeC1Ic2L9jLj/rQDK1fyS5adb1lRAZZ6AG5DyZyoNDP+HmlYv
MbOXkGAqnNutn8Jqe47KeyELHYkI/+6U0RlARqETkDyyblkANz51qZqMxN6cufnP
MH9ha2NuVlB/i5dTJ8FXgTtVmnVvAYBtTQ50xuEBcpuqOOy+2U/2UaN5hvZ3FEFx
dUG6XyKfyKtU0aButLRUlIr5M/SKdLQbT/lXSrShniOT4p+wrhhkmX0Au9b/foPS
krbO4xoFG5iHVG+M/EHMlmiaMjBcKjVriPNJfgXNHG1FCIg70PM0FqUUyTpS4pnn
FGDsF7G7J+mmBgvDeXVd0OjRGRePtBENeDAfxKUauAlfkFDedKnQCEksyAaw7xgO
p65NadGWd3Kx6NcdHs7wIhp7RnaUoz36ggeO3t4s/YvjjkgDmwPfGoYotTfeoPy5
QdfruNX1BXMQ0lqc0NwuZryg3Fck8zTfrsAniKqwmD8sLZLoc9YFuUL3YM6OWriD
bZ6byNC4u2hdw/W9P5iRWPVSeCQZbaE0SCqMzc18RW+VtEUBIX0oDQ+rjPbjvKQv
TMDBPhn2g4W9p9rUdiukXrQpbixy6AvLyv3ehaKyweQmVhhSK9uvBstFthskDjkh
UeuUNNacjLFfHyykKkZfczb4cNHsU9nRJlNmeHvTuZ1KVM0/3noP+F1+ZHIRqx1k
FH9P03DBnpWh+kS8QjQZaLukbpqam9p7K7rcwmmTz2lcgexJwSB89mkY010L+KbC
ocedRI4DMLQaFilbXtL+0zBKAFKgbqPV8/Zb4rRWPA14c8XppkdZqX5tIFNM8XKH
dRswdojl8JhVvcCqlBf9m2NZwaxqLmYsaLJIPnsB2lAygBM10X3j6+z/tda25C/P
MOB9fXbdXq6gf+aU7XnxiGoVTjTR901n9ag044AWk6eXKfn7YBtuum3b6oj7DCwb
gkqMwunD9EL42J1j+DAE+hXdjaIcRuM/CW8mpm2lheE13hv5rl6cALmLQ25FBWil
0qNetNM6G/w4MUURKtOVU9zEIlvYCUerV/kk99qkKwE9d3ghEg6jPobObdYwAW+b
q7KKAVAF0w9xwnxzr3caC6sjd4CKI1PO4DCWXh/xh+rxflSSibyuJz7BrFqbJxgU
iL2y3EL0oEdWk3USURbnBTU5fTwam6EAZdAP926QGwltPD6dwh7ow9AGQS25yrBV
2oGdfRTazUwmBZv6XsRlHKEqvqQTkpX1M60ow/SWuNPyzrPAidlNJ7poyxLVIpIb
bQd0ChhTXRqwqFTTaVX6nIIJ2mO/aZ3ZwkXo1vhULliMVCpuZaIBpP7YiAxHaGd8
kb83l4u53srY6dT08VjPZzMU/aXJksqIz1+X6KVrajYNskQonC+yyfFfdaYKnLw2
fChwhL/cbHIs8itPoX8iAnlqaLKwKnksbcIigPP79ejfyr3M6lG5Rq1tzQv9qYW6
Tv8Dtlj40zDdmWObBwPkxYvXx+WeivMuayjvacaYCZJ9iqz5c9GtD+dvtMjq6Fb3
bwARRPmviA4jLxeDXt73bSOlepy11gGFbc61PcMo/3XfSb1MtIIio3hgi2l0YjkW
WkVFn39LRieI411CmHOWW7XXtwpMv4ffeVQYy3iGChgbWIwCPKe5IVmZK2AuNt7C
E6zqgaGX3y8YNWoPTAYhg9XTk9ZOLB2gk9N8CkVNy6vkZW3c+0myMmjcvW2BRRNp
xTokqNLJyX4ZR63vAyH59DHtMmdC0B94C0FswDoUQNBi4aC3rhB1IVxk1q26ZK9H
wLSQ8UvbMbNPZSN1Qa2JO1PS7S+Uv6u+954BjYF5Ihc2yYjM8mFZs3npGyR9ofJG
WtwpwW9Y/I9Pzk5py0h49LV+Y3SgbzKyMR2oAtbccS4KNwJD7Gb2WNgVuv5ttaoY
HLrLqJMUK9pE+GaxkQvEmj9q4tHZ2+0QVzRS+eNnoVrHlgSgYWHvfSZV/KQIVt59
7tHnnLJPTeYsqpEyo71Lzt/xj7kVFmGOwjJxuCx3iQkfg444IQer56qc4gJGZUnj
ExRaUYsjIs4wJaZnmvnoAwwA/sSjZ+y86J8htQ4zKF4ZTALqaAm+Isjm4RLqRU9S
WS7ORd9SWbcC1PGn+vwZHpFdDtiyNpCnnPxLKFXxY7uhnGB7RcG0WclAYWGt90q+
SmQ5W4eTsXrw4gGhQlRo+5+12mI1DKADglpiSZSvIOlWMfX2SNJx/JAdgFbu8iYI
KZH+6EemzgtA5AbhaJ5shXl0BdrKhE5GMYk9LUls+HRb0l7JnPwLBRgI2TnZMVp3
rA8CUoR2AhoBGWac1hHNVpwVuGx1wyYXgVHWMOqKQ64ydKk0uT9tb7okRi0HxnDL
0H8MbTIXd4AsmOe0Cb89S8WidwvAYfqoDqnSYBCg3TgWywL4zjiWtWQgs5m5eBEt
kDNEAjWwQ8iqJoCa8wKnM9gsRruL/rkHLALxzI2fgzogiqRy2fxjDL35rmPthvcA
5ksIp2CJjDc1YF8RBQDVJcrE03KhsbO5LF0p4cd7gfU7bMUPJlqlJrIkEAdS3aHI
lWXXCHB5SueM2oiQSlLekgvYLIGnmBVsOrSz03JRXI0/9TKZcDCNDSr2cBkqIYue
9ALsBLTHy3SFWYldtTB+xWEqX+/PPYcyQ476moB8y857ZIiiuyLtjmL0QlqIBz/U
HRXDdbLW5PPJhCy8Djc5IQloYGpHIPDPHIgRH1r6R0x00YZayTdOHPZbWiufddGI
vw5asJiLaeJUh847djJ7X9SpxTfbuDQFG7v8VA+A3MW8JnH34/CIe/tc5sQKlAHC
cXEmDwAKXcrnRSW8lx4MLOLm9Vk//0hmx+bjhE/6H/C640T2l2I8JDcPCGuHmWnF
HTPLrA8UkvBkoIYoftQVoO3ZF1eM1Eunj71/ij0yz23cWeMybxe6h59sYMc7k9RT
GkhOymTVt7/mqItNwfmmg/mKveE2sP/1RwqoLh+QaHxPSDztGRuVQ21nDfUA1SEY
+gQ27wW9IZGOHG6qeR06tD3FFNRrY+0EvLC7pFdRLmieqKqT5hyAEblpEbQqjfst
CmE0kM8DGF/mws0yAxIE0afhdMI/hsxKDvyYD3VLJ16u0yAFnRN59NvPSoBtRDFj
TL1tBU1erm2MM5EE00Cct5io85b1N4P4CwtZVGJObeLGKbPmoh9A8RaIEdNEY/ij
x4BHKvNLfQj408NpWvRvHwp0DVeEsJYPbjx6CPo0IYirv6kjGDelm6OIOSXk/hRn
LT5xQBpnpK2ClfH68jtXttTYLNRSSorj/Zg/hDX4MYL6vfuC/cRCLMw33wZy5QmA
atxzvGE8PnklM9d3XHaV2R47Paj0dagSqqYRSaMN5W8RwNzZc9CR4WjfFfpnNOCk
kVCOXdzOqY6/GcvXaSNkKS72mhVK5ZdiEMgENjc9nJbi4tfR5MZ+j56AQ3Tb/AwO
IhgX9DwK5rR8SntkLhNgbwxLV3DQPgIoLRDqQuLwgSS8KmWYt9iWKVlnAI0OoLui
44VDxr19uC2FhcI0dd18cGMQxgg+YkG7lLXcsLa5Xv6sveNSkjOyg9rsXVsehgO+
k6VUJ2Shkxno4/vZ6qZSl7VRJcJDCsnE4davFOFzP/wVB+s9+pZ2vJeX9ZYo8kID
1CAGKoRdpy6rNpp+zIPmvhh1JTDH0mtnyPBE2PFAT2x38zD6hBv5JxVA4VIB2Qqj
kyBjpjA5h8d9NvmDXwNuFMqrUDy6eMGYA4RhJkFKXTVVTIkc+QD61dxFpry9q3Kf
sR0lK+Yz8byqSA6q5n+7DKXSmOHa0dxV9NMlajoe4hFCysaevTMMBb+guCOc5UkD
vGt6g0UnAXU7g8hwpjoK1dIAfCktYEMWTw1BcdoCvsoyHpaHkAlZcEkHcqB3Zxzp
O6tcBAAq7mHmEE1GOlHCB6+icQMzBLchSgNshU/QwgQiAWyoXRXJ5Z1bDIFudYUT
YGe4U1fsl0UOavNlFk3kjZhE2YdDPWbHbEVS700GGCzXXXZ6bjIWkOpvLKlK7Q+0
iyKi7rlY0Vs4s34RjepSReY1VyvXHU+Nl/6VRadkVMKhBkAIEj4Mc+ERzZDCL399
Bf5qKR8MWWE6lKJv9i+Hx3z/GCi48w4X0Zyc0fRFITze+Re8VC8Aw66PWiJGq0nx
ikrhOgpYgTKWQ2d4GIVtgwpIoK9YngXLcFPk+dMFe4raVeK8fogyZ9cnrd/CP62L
Hcr9ZFXVKUEi1gcRs9TU2Dek1/nef6tiB+XFteu6xvLN7pv5k+UwbunZKqRl6JmY
01v/R9KQ9FVmdDL+feKQPCRrjPXbap394m/1m3jH9T1eQ0D7rYoPmv65pBeg0Rp+
YcNF6P6oBoDnXaYSnF7Zq2NCyzgDhtDOjI+hj7iNBu7clruBtFj6CA6Xc1YB0DDf
mSpeVkGN+UwSzOQsoVLkdqsqJL4fzAfsW8W/u+WEqPhq25PJSuaD/eI5bmcmFFy6
IrWxswJbJE3JNcQmpJa2oKUTuUh8gSUNreAuJubRfcRl8xvb87xK2wQ9EoySMaBe
IVnIPDlLa69D7b3b4B8++OcvSKA90bMcw45eEY20rhb56kMekHwy+mWOCEYcrdA+
j1JsPTJsOBF3ARjnsXqWYKA6jYErfKt05+WuFFvWInUl5XTMWqMn/8jmbtifHWaF
BkSItK/gPZeLnIzbkOFkPu3ezn8cI52XzgkzPTUkuSQvEJ2Yt4Lj8VCoO2hM/486
6Vhr0GoXx7VP4SjbkZGF0qDLkapYeX06r0H7IFLDcsiEVHD6hZf21sapCavF+1b9
Zghk24dtWNMbGf96owqnLZROTrcTiMBN9xpjky6+VjzsP9PFKZyHwZkYuynf74/I
a7Fdft7snJleo3W6AhhvVbzFBGN24zb8Kk+YI5GK+o62sYlg+NvTgr60RrBQjscx
LCBDqZQ4LVTvkk224jAP26Jvk9e1fydoqfRp5+2aoWq5tG5q9TQtuThEAg183y+y
ajybPepoDZxGtrxsPK7OCrdVz4dzLavUHoGMDrK6Izuogrqi4IFiG9MRhP3fhl87
FgQUEhWcjqazEZN2ilWoMBEGj/UtHt6vM6v896zrOB8BcEynC7osbqN8sbbyJyEM
JdJHuA+N0ZIkOV0655SbOx7+Faia9bUTq1XgO95TlnX9yR+lL4/7X07ZP7kwd8dx
7mvgFkrg6GvjKP+e889WHB9ZtGKQVGMKmWx4AEJA8dgz2+rsQOFXEM35dE68o3vD
PEJlYTtD82jTEaibJ2xChQ9KZODD4Sfm6Yo4zfskA8tr7kZyK9vjIBuVkl8F6bj5
Ny7Q1KRFXkfkhae/S0nVjXHPTZ74rJ8hdit7DhHuXirjS7Ey2k6A8WeuegR3ef5o
qqBs+e5YxAt3wbLfTQS2zJdDqo0iDiCkTtnsbkE9FoOr4feSIVaOWwH13aa6dDlD
eKFxU+4Wm040aOfKF+w2BREHTpX0ql2Dr/5O4GxhLQVdG/wbIll9TyMmKU+erAbp
HBiOMlyKB4TEMcFcXriQjvBIqvAz9egSNJvP1jHA7qSqc/+m77B/8ewjG3oKUBQK
amKOtmzHl1Xs6luIa+qhfany3ZfnoDpfbHBNPBjSMhclQCF76IWmedEDwtGqb46H
w8cANREWG00gYGaT6HXp34dlQZIEsJdI7gUJzkVWb/HOfBs7J5hsKpwrKJZXNnfK
+QFqUd8nCgOcKAxnKxoKGAZoHuraYe+nYaLKmJkqoF2EvDzwa4NuzVWMg528f/HP
fZ7zE8rDkA2f4zpqMJT4+kaQurU+EEXBqcoPThmb2wx8aLPAG12tPQIXDAvltdFO
3SJmq7qIaF0eYHDzM8N5VZVOrhJ3EJwlEBW5ogAcplImZ43+kO2jjIkGzio3Xc2s
IDFIp5MMBOz5usoUzoClmZdKBmr+2fMZRdf2x4pQiJlWCNIB7jhgw5PkZhPntwiL
Iuw0Q1u+jf7dQC9nbFozUT84dG+WuO1tg/wbtdAEs8oUXnDNc6koxCfylHzhaXKN
Pzr13WLxDiNhBrfhzv3/Spn6AC6rN7C8de5wNB+UyAS+xWVvxX7F7DOg6GavUkyt
B3zdIpqM0rsaEtjOb52V1Q71P9VmYv1ykW6IFz7hCfrWwfeX7TZo1uOrWrL0wCEx
qtHuZPHWqH1Ad7FsD0c2D4H2Nnv7KvHKuzoQ1rP9bkj4Jl0vrGoENEVo1pmx5blA
jjFjkqkgQNljaouucn3cSprujCDsLc5EUbHXSVazHAyLqe0TCBkqfvS2DXQ4NZzu
Mont5DIvY1mT8he5cL5/QdC/kDuQprx9dRHSarCM5APFN4ESkzrm8IBSIq3lvXaN
o1qaKbdcySeBh3urUXxVSZHfB8ek42V7L2/apB22wqNi0BCt6k9Ri8/TzWUta4Qn
QgzxaHovCkwFuFw6JR58wLEulEp8QueA0h+AHOrwcSnNmBQTFAfXLUotDGxTHjGm
dGvbG3G58snn4WVVxTHbCxvdIOm5cjqfAJg8kK57vMn052EppfkKjdOtKXNnrWQO
z0vakSLtvGD15TpAJZwuvZSjefY+Bx0gtyeu4KzO6jp5C4mgquGtdiaIB1FHj5pm
ZNSwbICT9zlGNJqLxut7fJZ8D5tQP0nXdzS97+1ZasgUHutN2nARGYRGvx267EFd
iFP4CXPLjr3A4KYBttNMi1QlXU83jVzsdIjh6AFfZdU+j//qYvLWVZkK3NSub9JE
q/9PqKn5DUoWzXMtuOKv4hMLCL6JA8AjhGbEo2exiJfOavsFll5AcCxA6fNjr350
k/T9MeA6t6KgeyZrkP+cD3/EE4W2yQ1S6jD+CDPVCTLpNYrwnFpKTNW2QYG2wqXT
Gy0mAYXQiBBgYSaAqELPILceAQRGvsMMypk5DdM1fz7RAuzozSqs+wyiTVbQNPL1
UlZ7PC2u1RC0FmzNoY/Fk0f1Qi0GPn7bfwrO31yHUGhTPyeYGZ/dfpVcO3WsgrUQ
kZLnbnNZCE0ia73KS/jckM0zVg6PqV1rYJNwL5QaKXEKTqJ7S0vrcKkTdTrBoudy
B4qvTcZyCTC8DFvMtaVy8UwBR8gCqSkPCftW4Pavc/asTN8LxKdAFEk89SdKI/IG
JWpszGhg7ZYhM6aF8kxFTQUl8ms1HeCKRRJ7BoudiSfURJex5Pei79lOXfZ70vvz
XacxiVeGAeobHJv5M8L6fpGoXSLknQO1xxSTd6ktsBRmOOOqVXFRxOkEszWTw+Wd
YMDGJcQ4Zpkek4T9Hr48X93dFWPWgyVLLgHBnMJrzrsRUK23g0VywUr68JPmSPlT
6/i1EWoh4GzMoBb+I3Zan811jyOyvRstGPCEws9DpUEE5QZPQKxfuhjeEnVxNuWU
3bFTgRkP3qcn4gH4Irz6adu/5KhVGtow+CiYOoB0psxBvw99m2ecpEyP+Kdx3mYW
Rl9FqJta0Wp0IA8Ysl6wa//aOG192DfBtGauS8n7IOIyGxnqCXlWOgpAQLYJxz9r
ZQbW7z03DqeBvfMSdScO5W16f/qq4AXD8nKFkO6FjQd+ORStzZui3idoOnjnbINH
wr0dR9xQtD+HGI6s7ZKXqBFOSUe0xmlLgJEPhv8r6jZWE36C0FwNI2XxKr/yc4PP
HcVpQLbjwYbGf3BB/I4icXrujKOIXCIBWHOnFBbEoLgGgEbaAgY4Q8+nmoUcMnPw
kt+cZAZ2scx8waG29D7COv2ZjJfovGMNmneUWvA/Dd517oV7LeDudCBo5XCXg4WI
9XvgbEAhP2NZAcehdrA7oBYNomKgeO6QVE2BFq+xk+yNfxjJ3OSlUHHtAttP1QQH
Szl25pt8zWzARlFxk3puDhtvxQZ8hqR0F0RnPgZA4BR9OH+WsCV9XgUuY2Yc1SgJ
DyPwk/cAlkdSuvGmnFu5+DO2HdTL/cb8TQOVdenttCM2KeM7ARZVUvH2DbVQlZ34
PeR4lnCHL+kJ+1s6gu+/Mh4mxHC6gE69Kw6z22XamgHM/OE9tcMXXRd/scK8EwZJ
5svg5OfbXfPu/wtP73++di9lgpTC6i8UU4xa7qHxovSlNx93YvywUGAykaVQ0BiN
ucEH3v5ng+MyqEl+yCfbfag6Na0+WkvqB8EJgexqFzGvC3S4nakmrnXT+wXbGoRp
bHIV1zY18Y6PT7Nu1EIRaPSD77R/snP3JZgDeuY3Xtjd4M3jzro2I9mkH2DMBuyG
IS6Zo6AU1Y4fheKk1+zpQzJT+YPsf4QGYTb7j346zXilRNlosGkEHR5nTXIpwhQ/
rTF5G9K1j+FjLy5l3VFf1oQO27o9eadDcd5Cw5oNEQVKssL6ax+q/4P3cZiDsX6d
2J8XsyatZ+Bp4VUnjvD9iz1WHcnljfeBTZzQtJEMMFRjMR15+bB5UV+7AJzZI0f1
5ug16/j4KuKflrliY+IM7gm7QzLktf717uN7+SidrYJyX57KlujV9beq0R3e12oO
EIIfN8oEp561S9VorFVS0yOho+I1lu/+057A2h/pkjba3UVd/f97o4k2heDzFiVl
Wy/llZmNAoL/5jWVCTCTSrBL2wczux7fj0Fm/aDzeN8cg9lTw17EYzFyGZ5n5aRj
PHtMNeB0KquBKM2J/7gjWcSgRuB1YaCTe/Ked0ejCr6KZXO8OLxTMVhSU0UW47II
n4Brq/URMRtkNJ+366zr4TSfY+ILORfb4imUeWc+Hlxrik3+8kGd5pxixMqFXjF7
wBisqIqTWuA+aZheC0U6NzH81r2QxoS6xjOaWmWYqGm75Y6Om5Zq88jnvp3ox11z
AbZX319moku7k+lunpNlGLvLRfHyo70XH98X6MllQsg/60qmsxXZbgH3DFBCRtWY
3ioZ4Cvd3UTlG7/tlI5GzWSDsJhw5HWwt6VAEXgNnn+QPvEFy/rP8m/yNO/b5UJY
381+YoYZzI0UgN35yV/w/s2WTg1JFXyXz4kru+5qJxImjTlb1CLU/cO9VVi3ggXR
9Uayz/QqqLJ1hCZJVAYLV8iYBDUwJ1XiHcbAg2E9J+D3smgioLoUU9v/liwToa2g
R7BvxldcVx+aoikVxbbsBUyfg/N+7uALhzWF8p/6OlQFKsleCT11ELrw1An01xcv
2J0a88vOsTXqBnlTVy1GdfRbyKBQgIa+/WThsr1pqsh51RR1axyRH3RE7mUREg3v
oCYTn1fkat3VXYfL+KwSg7yqjgNkVxAOuKlv1Vjk6alHkIHtoXfaTSlb28HJMPeX
WYzPnb3tvD+iBec/53ninGkXBdXgE8MD0xZjMYSkPd0mMKvggiHYuwmSPtR+/ZLS
B5hzOwspOzb5Yw/7RUi4v0aF8i+jz3J1lZ/9NBUAaaqbxMh+IQjZ+aUuzgxVLxHR
Q/l5bU8fvogsvCSfNulk2xdKkn4i8mtAQGhAGtnl2Or+d5QS0oR5CzONwvP+we66
2pum9xijK0eeuWMClNaWwNS5ganI7+ZD1V0/qIMgQ8NkprQBHOFADQvDSMYW2Ko6
fKHtDYbi+xuODCmQgIX7x2J7Va8JKsjYXpaw8Iah6sgjoSQZ26yNnoRAmQhHj+3V
ydcQNmNuaIpVoQadNcoIamvGiIPPUsw359Dv0GO2IiNnT7AYQ1HkFflEdvSaMd/y
zOb5pL2kyzsrf8aXqHQhE01AEsdCTGF65Sj5dQMgxIFjD+4xEHu4nAd+X/CFKTgE
IbpBuWPsxGeALH7nO5xjAaheCe9P2RUAWLZBcgb1eHYuQBoCO4PNRgKyZUs8f8eQ
RqnugndMwhZiMIY8QKXysV3IIKgLfbeEQNRJmXqXTS2rAYbOwMj5meD+KzAdkOyi
a3HzuNntiA3LWLm9+MgUUsqSWwoBBpXJPJNryhFrhLQSlgz6d8Vti6FzM9p83eNd
F9eH+9q2ByadgglfrJpfVn/d2iMsMZr1iCPlH0/0YFDjvEc8Rje8OX5KuTB6otYT
UZxMAAYIuXIyITukuzBQx/KmENTd20NtOdY6RHHLkrQg91kcABdoMls+RIZVRh0j
oikhIi4hZYVSSFvG4iEvaRy6TQmD6TPLNit343UTyiCohJSdrafy8VkFV00Y70lY
ysyYMriIEiK+VOx7vtEXJeX5FbQAMKg9KTPdiQr86oQR1qy7CNZ1yNIko49cG3Ey
Gh7fm3j7cX0ATTBbjK8qsnnPDAgL6vdPjsg6s4HZOLFUEQKQM4IN7slcS+Q+VgPE
lo7whBQhsG9fP4/x+1ELWJ8393kNS15DelVwDCoPytGvEFjO7fko/l98eT7bWKA8
OFGKXYcXzqXr0Sxbm2JO7SZYyGNfiOk1v5Iil5hkAMsnN4eigMFbQd9lSfjuLyST
GBIE87iQKRxKhA6scRwiLNL08Yh5CaluIDCbfl2y7v/sOGu2BV7kD75WDpYV3FTB
xmnaz+8WfyotOAg79z+4kcK7VXwTaGvNV+af0NerSzmPsIoKG+acSX2K26xdxe3k
1KBOcJlpnOC0vZqE7+FPANzU3wmT0k+HMtY7bKBmrOCbX+8jAYK4BOLh4P+a5mh8
hTpBkzrg3fQmRuGi7+CkvEqTwvuEWw9B5ObGGFoVZavuPbI+7BVIYxm9bIkX3t1j
8Lmj+o2sSK59QCPLQyRk+/RBRc4VL6Q3WovkgaNloXg2RhLhi1X4DidsYhTjjhGe
ZtsbycmcbrAe1AmXUWWx6X9zsPA8mnvaIkyL7BEpSHaTSiTT8nchMc/BKpsE83yh
IzI4/XT6MjBdIxF2Fji5NMGdWA1xbWiTI6ZbO2XJejZ35goKUsTmXFpHiy0bjX59
i7vUnMYOmSxnjpvZ2bxIPSRqdRxGFxOUtM+BeezZAZuJO0zPp6CJY8F43GJ43/AV
vdCPueiu5ZkaxihMaN1HkBRUmso+zhtO5hT9rMTgitIMSyhvAwroslTz2bpEy18d
ykVLrsC62J0qmz1lmwU4J1s4sQNEQXqT1LIo+xj/VEjbbze8BQpvUzgBVY6fRS1c
2+hltjD43aOlEn6LTXNwSLNaWvRmcphZzpZbDQPtN0+kebPAEdOelf6FnRJ5byr/
3tCZB+2AZRuxg1iGabyRq+3YIVo780ggULoHt/SIAlwZrLtoyU0eWjrEI9JXQXtL
A271H6dxwpHAOjqtkq8nUEPwVbfO6JYvjgVEROP3qehWHnYWGrITDgZ/2LBs/3WP
QuTAO1pq9q7CnTH0Jj56qm1VxOA3RKh9mj1MbY6t8YYy0gdw4lz18bOS3LbDVs9A
SYs7xlh1/yRB61Mza3QozVWrvaO6iSi7VtAHYQhYBXso2zZ9M7jb6E0SoI3f2R+3
ag2OmiwqsZ8sP/UJ6v2jN1nB/fDubBsV4kCavYjNh6qbXqmdI0PZkibwi01oIkDZ
QOVcRMMouZWBvZGEnHH+g6+E1Hw1/37vP0Nc4W+XUn0L16G28Qohf/134/LbulHx
wh7q2yJmY5HH7dKswydATmM8wQcv/u2vSErO85O6GiUdZA5fiArau8Ok/QQeDsHQ
er7fhGv6v+zFRwI1IDaptFcGm2WcXFzkRuHe+Lm1m0TEDUV5GTOCE8UMEQ5PLl2G
Nw02OTijbFu/2yO1EB/e+gSknScwLLqsV9qK+X0kw2D8CWQgA5xziH2nIL5Vd4QK
5wr/OWxorQEIzCA35hWwcpUI2v0TlUM+CTk9n9igVlg7nY4vGwrbJpStw8tzBDNA
wMFajDnaL/v2YdYzEMQakBA82i+e1zZq/Di0Hg1e7RAef9QvC0v7Jj/N2gjV4Qlr
+reVf3WRbEa9KkeB1z3SRlBtPQV0UwcUORQ8lNga0ppIpE24FvnwXYdxu8uR5UhX
yNt6/I7BuZL05MAqpwM5G6b05pvMLXdUjXSHEz89XJg8FZfLLhQqweECex1XaJG3
R1NnKpPO0ljb0LP3bpoShQTSxt4wMdc5+4+vL2CR6Hs0WfJ1rutQ2YPIAv5tMD93
+e6XOfOqVzYZIaa9qZuGkp4a3HW12fZEpavgT/RnL1i1ZavkbbTn4bFJT6/xOpBy
Ftnh9QoHru5ug9vObLLTY2aN+o7ljU+eUUrET8wS5dYxA35DYvQ57fuIDOhAiZxc
yI1YJhPOc9nTGiT7HHezG5/R+rqHgdoNsHmby1ZxEYhTdE4Nlp1sTpBpKztIX+3B
JjJ3mFuM5+b4gW4QmD/10xEXgeW63k5d0GISB/vWR0rakufTcZTXQhxWdixW/leb
Rxih8xJ6+n0ZZwQhg4nVEJ+ds8t9yFuP48LpZTeo4QSG0Pq2zonqBg/nY/afL0g6
OSRBvlqDsoNfKJQJhzebD2Vc1iXGhJxsS/2Eb6TGMO9AljDHZJAVTgvy6Cxkpknw
nuTrng/ciu7VtVT+W5EDU7izK6v44a4D41YksyMu8l5gCnEwndOGmGVmamUWTAra
JfgGPtl+EfRSKl6qLw2ESNXHC7P7EwmPiFZDFFb4OGgl2OHbgDAh0i5TdDq7L516
7bX36uRC7FXRbyhaOyRwNJ6yXUyLYnXsoD3Ui8VcJIXt0YVfcXsz9TZ3M8AJdpMr
TcuCL05grv2tWo8HeXCAwteuAB7a2BdICr9/0YT8Fvj9/bbwZO6epomL2ku4HPR4
l4489HCcFgx2x+38NK9AXxS3biZygnUTfmRp4iGbuC/kqOvA02w6dI4K1ctwmce2
ibw5qU6CdL//4FV7JkLSaJrkuznCJCX3NPMj879/bUKrtjIRO8YbDarS1an+AezL
jxbIxwEeXGebeWARl6ND6vyJqrV/vWTdK2gm0YdByGUBolGYEklptSbJluxn8lR3
9dPLtjdL53XFJIeBNvW3W90MO/eQOsdAmggAfiQuBYRkxvDvxD78eWA4ZxS3sfSk
ne4mKlurNSAQUkTMB7vKv0rVjhunRQ4pmw9yL6f6Omdd28fjPzlsL/MM3pnq1A0I
c28TlhWPEQKXeZOj4TDQztXdTswOMevfXHGDO/TI1aWe0NPhZD0aNy/7jUJXo4OI
Jr2GjBikUwBj65zv65Swxrdgc8AVk7UrlE5v2jFysXzsnvbgpErRCoh8Hw4qErhZ
3S4RFNARdDyunE1QXdPE94e6iWa/lrJPDhtjBhyOH6it0SNQuJBQ7DOnWELkm1XB
c1TA/Z9V5om35T7HHDYee0IHdDZ5G/Sr6GUSVxzPFcm2WxM0BdGAg/8BXfb0MrcV
ypUyZ+j4Nb5jkyQqnBByFd9YaqGf32ouL6eCnCVcTNM4qOAYYoNhZlz1LnJlDTiZ
UJgxsVBK9eSLDzIewiGp+9qXVme/PRVGgB1qbfdosLufq81TVqmr+sgH1fuX+tlG
fXB5r8MIOjxNj5jFttCJlB39ht46W/Frv9dkg6gWogOOdqAthEVdN/R/wIfrWL8S
+3ejEsDj47G7JxNmTP1BcFD/5QGxaRSwiQe5qOhBi53tvXwI+/G1bLQG44bpuqNY
BuLXCnGa0hmYlYet1X9JeA7qLqbCmMV4ZOxS9q4oXAKIFNS4AnSTC+eMwKhF8/V9
k/6aaiJEI2mExrdHG/wew3Z8BARgwK7hqKfpcbR9n/BCPpP6lOqZxH7YYxTwChUj
z7gVVoyoUdEDMbXMXwCzBL9XxGdhxzV7eGQh7z62fPE9n31oeUGcyoUtQHA3VfYg
+a9fahcxytN+Uyih+XrdaekChUQvgwmQsDBhfi743iq8p2LozGYW+UOOcYN3nOYg
aw044vMqq+Uz2rikYacmT98wS9K3gnHFFW1pAU/pzSBNz/7lMa7nk0D5zq3AAFdx
uxu3qSxid+urMcgr/r++IDvwQd41V7UYZfNsSQRQb+1/0Z/WLbaRVuTJf+kYPppU
0VThaPgvoMtGXaT+GvxMCmAlZQ+gvxyUTFlGWZIImujefanrXcurPKaoKoTdzq7/
vIpDn9o0RTYMVMV/3ZpFfOC4CEIukFyajNdMGjAsbnY8K+PE5OCMSehjnO77ZUbg
SRH0glRvyTP/BAPG5fUJVQue9UuRCsrtPy2kU0m9twcJ04b8TbpwCzmIEkRWo1vX
uE0rM9hF6fyty2KCgW07g5CZ/9TN+w/wSmAHLoJ5u7ZzZLoEokuxp2xIAxdddCQJ
ytz4pi9fiP6/gnZenC1rsm7e18TvQAsv2iszkR1Tb2PXQUgJ/10BxB6cTsqSklZL
UZoM0pjdW/GeGgLBpjamUI1K/bJTAAsjK+ocHoycBfX13nvbpW+UTjSFr6L7/qtM
Vy2dFtEWCmdDnzwtScK8cCvWTrxpeSdIHtxF57+iUinZPbBung07IkQjGJywumoc
Es+HZjkP+1tlJ+Bt7eHx9s2Q+nKZOLhivTd/Lw+Gz/nFe+LIAloQNi7uE+uUB0L+
epAlObO/1HMFyTWWoy0R1NT2P/2iBWuOePMKBrOLNJ8LY6gTenDMka81+AOo67Xp
NVTF6/UN3XXakV6/ldWsnAYMBHXXyf8yRaIc4yrntHXSKgX/5QqfrNXvJ6O8yYZa
vLKjm1ALq0CnhMQ/+NVKbFAy02DXgYQJ43bCxwmnyglqGdvHcL9bzlN7ML6+vV0h
5Wn0khDX5fpWtLxZ94tHMxe18BIxlG9LpjPXda+PvRB7HPzc4MKCzyb1Qo8Gf7p7
4JYeVpeqbp0xCAQaa93Lw4+hwZoSn3m7xvgSMmzxq2wo545MbcaDrEQEL4OspFI8
sxsPBGMC0mCLiHp7SVVA0TT0Yq4B0T5NuyLeOOTr22OkbxxFRkiZ5Ov3LUjiMOY+
iYOxu0/LoCtvWdayhwzxW8gOV4gbsfkp4vtlCv+2MeuGRkQA6Mj/PoOLjLeM2CaQ
rVi3sVEEYtxKxwFECB6DNXtEsDux1E79AY+vTzMhdsUrQXJ5JRc7D7wo8/6yf0dV
ruZfCbnn+LziX4Hq+E3ZTv/p+oCbG47t1zWEs2AD49DOQBh+k4fXScsAWCeLjhWM
FeQP4w1gDGL3aGyYxipyP2VdwvIAinduoUjE9AJnB81gd7zInpsyhuzSWDLwp45O
IaqSZx1DI9D+ybqOb2UIvOr6/hWsLnYRhBEVUlB2+ykat7uZtzjaV8+OW0pCmuXc
fBv0J85ayh+TdGjJjBH5gpgcFpWDoLoMrPWCM3hplNFxSX9MAE7A+xRJk/0eTtVo
aL9cw0WTgCZMcOYALH9owXQVYYwAMo4Vyb/RoHlsboTzWwSd8xHdM5pAkXY/YLfD
OyJA7QDxMbT0qncWWBwl56NCDar0d28ONhwqiHrIY14iVa39TM1iEExyqYs4poKS
uEznC4RTW/HVciKTvH+vfx+3Tlw8J9+wACMIZymReW3doWX77mPLs6hgfB2uyKtr
3SmmiYhF6JibiNG5iZxjjaMraG0XkZvsTAuHyJrLsb9u6BKDiuBCo2Q4zRA6JOl+
Km9i/m0TA28+Pdr/bqiq6+EtlU9V0JD2iXApwy06/bsOhEf5IAiabSj6p+vofhR5
odJZ+PSoq+CECOUR36mq1ARhmS7FCe4SP4HjroNmsv+CuuA9AiDWHlCOToqKGsdh
WOlB7InRamgkLSzzTkSzSi83NsaAOzpFBhVCrRwoCdFswMO2Vqs3Gwg/v5GXS6Ro
s3vwE7c9iOgbx6pqjZwJp4qSTPCSh02DXl+BptMHFuId3UNds37DtqLR7RdVD64S
zECPUxIVEYVvg1L51QRrS4r3XhnC8SUDIWbBiq35orXB8178Tv6WRRPSutz1wC2y
COweH+vH9neAA7hICxgvy2RQ+0RTgPN7YaCznZwfp8zue4vKqzY1K7WvDwx3gLNk
jfHN+2/tFxsG+7241tP9st0fUg8g6zjG5WSEvyXmjPGGKdwUerV57c+OuojNWbfO
Tzlb21ps/xjPUyEWcpA5beHoWTT6qa7ubZdVHggk6REKxIq+vzRYXbMWXvf3mdgG
x6nvrjXNOaoqXZ0+ubr7xYBQaDGpND5rYWZoYncTxm+/54rQM9TqeGkAhmVcgdms
oovJkr4xLu4TQvyRJLjEESOdVqH0Bo2S15jsoMHoFnJSZmgYy3PWWCsffzk55JuW
LNeQAWT6O8e21ripRD7V+BH9r55vmjPtvXj/empB08x2V4J50U3qnazFFKdEEFa5
d9dGbwneEpoC/zTmx+y1+eBoKbOzeSQdpqOe/3A1CwseSAE9+fAlLkaCcDLAHHE0
pllUijjUUU02nl0njooIDywouNLc0tPINhH9P1cgUr5YaF2g9CSw204TaZT7I71e
LeqVXtraYYHzmV65xq81VZKMpEPNp7nNNr/3UP7ylM75CJ9AOiMMo9G26THA/Wfb
BnehKqJRMuTe89Xf4UNHjLF9rAs9vZgkDOhVlDVizacLbz0ahyjKhTw885YCsMZj
J2OLPJnjG/IwaPnErcV2KXkmOsHAdRoK3Y5sdtSAsFXbhEmupbkS9ssDbBHg9THU
h5/ioWzjQo0QV/O9rlsLz3ZyvOOHbtQRgGfDopZcOU0De3cpez09sOuDBaVxrR6a
rZYe1YEwdVDqDSVTL44YTF7ym6G3iqUCDZd0ko6eMFjHgYWle7L8/6AJkMiDuo7u
tqRTbrw7YUSy32H+mO2G1ff7XowqkqAgjqx4JdMtsYxRdNsNfrYy2+tJMp4jTpqH
dGmt8To5tP2JBf8N/Pfr9ImsBu0q1kRT5M+u4GJthoqTp7norfvvcsfs5xFsJla/
ba/t+57CLVarAqC11n+I9GMO6XVaLHDgAc9flUd1KdISl9DLWRIo0tQABGDRmf4y
XWvFNDhQipI6P/Mw98zyAp/InYz7IJeNtcJrtWRyrFBpcyO1JoefrNblvZJ3b1gC
GPNNnLhZ+FG5NnpQRxRWIyZDVs6PNxMAdKa8z0Fg8Bw1ocDF7Vj3Zq0Og8/7ryn+
a+Erv8ib5brMHJ06LHx1JN2rYovoJbRIbrp//I717g1n3n+PoMKKCwp5yMuxzWYx
1NgbVYXWtnUOoXyqbIjc/Io8YXcL35lOq7tnopKjLWMLIJlR29Ylr0CE/1XvcjY+
fJw1EU82aUxNDnHXExJN70z7/OpdbtaD0BNfTo2KoyICd5EU2t7Pn7W8Zuf+/e/Y
v1TidH0JvS1IggpBr4Mb+HibRAH5rW8twIewSrsrfYJB3HD4UMg1mua4+SjB+6ob
/lOHOxXJyta5c/1DWNQ4VZ19bOol1nDQHXiL+ul0OgT6V6cAg4/0YzoIR4Z0aB6p
SO9vbt6+78Kb/ITSPEZ7XPSuax57yvBf1SdwSNx6HmfnM996zq3PDc0RroExzLy6
TzxoOrUH4TP2opdfguRSYbRger30WZMaNzvRgIHpm7P329Jt0etDXME5HIvfl6Aq
RZmk/og0Onhs01N0Q1sfFqYdXpWo+qCA+L1WcQmQjvKA5gQw/3as2wJZqBWuogQE
IFpiOQQ6IGhHn7I7BXdxeuGnfhVWLdalD5+zX0cgdRweTBg8QDlsezjEcF/LBdPi
+/vwZszz5dyGvzGglWglK4WjQexnD1RHbNzB1WjIE9M70c65d7sA1qxH+KM+wqaF
qwmGJ22fzTsfDVrej1+D3iZE+cIxn4/8Nmhl3koqcHVIiTdnv7IDmm+zn/6gQ0vT
ryVbFJhHdthenPl5XdCPK3EpfbpMltZJS3VfOm0BdW+CqYC8TXEAoB+No3Eqlrz0
j9FvDoi93onAxXk3tkp2+JXSC/Es7rdNAWuzAeL5vTgrTBorLupLstbg0SZmniu8
4d3AgmWriD91BvwiMS0PKfEGBF18j8Kq7Nhm5ReyXUYwNzoPzWLyR0m1h1mFPr8M
BPDZRYzQel2EE4StRPJ1gfHxKwPhgGgrcpZEcekU+e6IXVdIR5vGAqCop55zMJaD
a41NtTcC8C9MFdZjEzdN/NWtxmKCpgEUsmA6zSCLlQcZ2zaLZ/Fho/8SL6qmSLRS
ZLGbn2+ua5AWjGx1xMPQT43uPhIz4/rVE6jMl0TbXqyiVmx9obm5zHp/BkmIuNz1
3V0Bj+/uWRUdzZnsQftWU9ixQmXjI4OFK6NaCpyWMC7dwWEx5qreUrG4/yzqNGXx
G5ZjM7r4uI0NsQUlYxVw8ZMAXzPRmXk5VWXTT+tGMFlybLGlpQEOrxZzWdWdPkBd
BBEdAFB0jc+0fTMzC1n66UuCxAx/ze1znxrZnp6ATI/g2vTD/uTTnOM8DCF0WBP7
uzuzN/5spAqH85vn5lgLFhLUEeXG2Ytp6uygqekgF/15x6sXFqfMr2xIqx4xMfy9
wCgEh8O9SIyNNmhLa2wJSyd0zMwh0evVwWk6uSU322RvQTfk7AnuY8SRCnu1jDBu
VImPUMSInXnFG0vxq8b9Izp/drRX8goTzC1jTAnBcJUQ0ezsX6mW8PZW+ydNK2ZC
Avh2XkyHCn4ZDsWhQ1VidFQ7NhFq6Lyj+EizpsksuvJpD0o76v+8RW7qxWfZDkfj
+AlPWQ+9PKnWsz/tJXJTG5rqsZN0q1PGBx6aHJXBb4Q4IVsKxlEPcoUutlPcixcL
iQKr/+vVt6gGiw70VmCI+BtFFboJZtTGBkzfVkyYtjU+UiPap2rKklybUtGrNcbG
Srne5vJjqFS7a97lYIqUsQVnUFQNFFRjVobWox8LvfYG0r/JPaPz0qDbhPCg8F98
0GOMpwP7OK/NvgSsqI8csCV+LaPh8AdwJLj0YLV9x+I0QJEKQoathrKX26GMevUb
LcZawqs4DfPxMTQ2h+CuLTH7Z6Pm9dEQn+IDTnTJKsodBMElU8CmooXxu6QPy2g8
vSNb8noLgoLGV0jPy2UTfcn80z9JcynZLlU8kCxXAWanOhP/WDqM/4sS+6ndRAUE
wgN5YgNkAPOr3HZa1jtYECCtyW7pRWh/aLM1E0W1c5decYY3PvEPFTAdf6pkOq5O
G0qE7YnaeAHd/0U48pg29eRBils3X84Lp3v1J5v+lzKZb6ivysxr/tpBENm/ohuv
7Ibrv0dc8RrOW2gKZhNOKOWl3kp+5jHe4aNBhJqUWWVYkRtAlBVP+yJ2D4Oadc5m
fyaAcmO7/xXjnjzVgM5X3lV+i9QcU86aqrC0FyIcyLIxD+t33b1EkjdUlMnVZ93q
Zem8QzKmLPxwpQL0Tc+QDLtuZOmwarAYNAWls7FEOPBxqtDMyb0HREgR781Gxx77
0oblFqodKo+3smPABqojugl8aVG9x4V/0e2Rd2E3Djpq9Jp6yune/zfGbrPV3Q1m
VUs+wtCs9ogcPMfOntdWV6H/60ahNH3XQKoM7CbTh49nI3Wr1WCCACv69+Ze9pZe
LO+r0ubqlSxyEJcpjYWoWeEgsH9ESDGmGam5BPlwM6wqce1SNpETukvs2f8eGaP6
DCwjuJD+vZxAMBlUQz9hA1gFbAZAZxGolH2cs7DXLJq3VXySRcEXjUU3Vk3iKTp8
HIFVaNkc5tVp52CstRBTKc3wQGOsW5aU3bEt3zQv+porI9sEulxh4hvuNQq0B6iB
poPv33ZteElm2OGuJK8i99Nkp/KwQQwcYIzQ7rJzQM24Rg/RLwtuVoWuVvs3WmjK
uR8hfos7vRruXgdWqaZxVBiIbUVcdjAth6zbTcBne30gnDjD70mC3skv11Eb88su
1Z7vEmhl7/GVoYgXnmeY+VpcDPTaZg1xl1BY7yOqc6S9pUeIq+oi3ZdgBgMmxmBC
TNsjxUQfXEbAGYDbDZP6CXryaMaU1TvjIECYZLSQNQNblJi9mrOpommX3h4xGu29
NkRq1wl0igBKZXI328LhT9JfuuNRVHYW86bYKu7QAsoiT2zszGXI3LVKU7taQZas
gVmFfmtPyS1gHnt0okE16bQVe0GFaWXxpp8PCbVR5C8cEj3lhSnpKiJzzRfGtj8n
c2Gxy75+JBWq1aa6hC8XQdeHRcyF83RoHoQdwbOUmvu35HnxquIU7JDTQj2HUeJg
sPba8Py2H57/mgV5mcXY/VD1UpD78QiAPrcZzgS0kaxvKqRixFqQuB61tsxvWMkm
QqoB9tSbWobSYZSDtyaAvYq8ybKz8JrdiM3WqTJjMfBmo+hDhpZCdrlR0GwIqU+x
TdXN0yUT7yvirAT02o0S9ADutm5Zbn2sGgg9evaUa1BFTFexvfVLDoIlV4v0Sm/w
5eRnrOTJfirwzhGrc/f6piFqzZso+2TLs2w3XhU1ssq4h4x6yM+UqUGSFvraC8JP
CePQqEn+x07g39D4zmYU/6UwGVQufIDFfRMUNk59FO3M7qjjf4v6fzWgpQ+BckNl
soGezRCT+dmtfsvIW5ERwJ4Qjc5/JAXzPLjjg6shpeTaTHlDZoUOIIz/4DWLvHRk
Ty8D4rpaJmsC84pzu1nBfz7q3bRR2lE9ucSTIKLBP3aEbH8Gnj4xo8HT5JfXdryA
WSFw1hTEV1kgqIAuG1JO4pbS49wx6dIhNxqKw3DwvMIjOxbO6Ff6JlJTjxStbMUd
uJOCcBX0wNGXogKjXEDJEa45/Jq5oZ1MABOK4UAJf8QOmi5nCxB7EZQaCb+d68mU
/Gwyn0KKz94i4kQWb+98aqYt8lMqHste5r1TxAuwldUMATkcl0MGhVj/x79F/80V
iW2/9Ksz9fyIUQGcQlSXiXUIU1OigH/U8SvfA2zfKKlykuf/mf5k0rSHuAbUnLvZ
clqIbRHqd2a4qKLo5lLU3E7nF9A2+vWRMC8QpHMKLhTP7lPHIGlj2f3E2sEUm8KD
zhhDdOEQnx0KveJtJy4FklWc/MwFTIttiBKHSdRnvVFmbJCtR0jhB2EyTMNsOP3y
Bo+MfxCQl3pugkcJlBKBOwzMLELPVDgTNZSFRMYt1w0NVX7RYWUaV346E46NiLdZ
Ne1FMhomEWpb6FUMuME8J6oXN+agwrCZJdryQrqaOfTEJluqsgpVTEzlKmOdyxWO
YQwG6YwdQmh25hPbnDa9jM940nN17RyG3ga4XGnObsHE6kCdFV8VXKc1oYglpJ0x
HLJJko2rIR+k1KKZmrN2pLyL3QrEIE5crPTJKzMd8UX5DAp7rGP3z7pQVZC/YbKW
t4AIS1GNdn2umGECEyjNF6u7dEPzO3KJxHkQQ28fKizMhitQf/ci3K/6kxm4ydEo
pb74YCI+hAJ510NkR3Q90UncSKk+cz8QzAP1oCQv/y3C3dr5mJ331CUNw1Bnf6IL
YtY8+BR73YUx+9CAkUpAjqZiLPa9CVtTRJZX6DLsiO9ApAsaRQ3e9InGMt69f+v1
nu+v4glTMD2Hn/NUtRC5arnF1nuiXgMqiQqaNjRBiHy1t7qI2HWKSmubTGIxhKgp
8+G4LUTX3NXa6urWvXLsAasGioB7JKVjSR0yAoVOZ9tQupujPOgwwAaCR1YZhkKe
teHcixDaz9TOpOrNnkVcGO03pmv4C1RjWR3+qQ2fp3wFxH6dXoed3v7l2bILjLJr
Tsdx97wZOElhtkhrKOJMr4iho9SyufeKaDqafwf4lkxUkMWEJ/il5WFrqrJUK6uu
NY68hbwDDgGki9wtMO54V7Xug8cICmI1dkktlDsvim+A/o0kDXf3zukuBxJ71aaU
tG1u/VpfEic8tTmeNWZY/cLXUkPnZZYHZmzS67k7ZiaAdCYyqAEldl2vGQ+ma5IZ
+TgTRFIxgQbLOEeQILvBBC7osOKU2wZDm551fTcudAc75OB6BvASSrpSfmmeGIjF
khIbK/PrC0znwhkhK1q+NgeMD56gcxfOs1FjK0dKkBkbE4aXRjwgUWOewZsIbK5g
uuhhQeunYbsgyZrZVVl8ajc8DuH+Fb/lPSioAGtTSM66G20dHHbVRy6oITX2ePLx
KkCojXbAjlNq2J4+/CmhKy06CMukI5wTbvSEjZuqakGAc/YS+61YpaDuse1QXn65
hXRFWBNKf7c5pVN+qDSDOp1vSN95vXb/o1SgvBIX1ARF6Wko1q4DyE1I2pvxD1Ck
UV0u9PFcwXtJxD80oT9JOVNuGSRtD1FQkig3qsq6rCtoMSOE0Is+GpNn83KpTo7y
s8ILrB9O4KFIe/WgdYkjUng3Okx8j7XYem3kBWPVNEIblxDqZEVSx1uybDChSOaF
8K6f+UlQGT1X3ofOf5DmEPlVmrcfcRzDxY88k47kxjmaVYffVYa4WV8zrq0ylY0l
IcYqyRICVXryosM0SqUmXDLZ1kfoPUDp4ItWz9yVb5jR05XFnO8nBeNI1OL2cWMS
yfxgBz2PXZzx0pqt1PmZyKvL6B6Q2olvKKFYqAhM6gy72FOBtHl1XLA3vBiMZfJ+
CCHrnGUksyLIDLz+NduvPB8m+RcuDXTk5botPD+kBjE78wvqmr8hntssdsh3sSoY
lCBtXnW14HiaK7malZnjwNb0Xl8vAPmPArHaCH3uVT7fnJ41XF7OFHSuLdrkawrg
CIM+IFxnkmYGWTTBsZrNs/Om/OnV7JkV6ZHi3+9raySvLV5tsw1ji8rUa4DYhsRF
kGr36XniWWi9TglanF+fn8VdguFOViqZXhsIGqyIhxCCLSQoXfRya7sVlLxjYqHy
1Xva0HYDB/b/uIRV1UKuG6WD6QbcflrljWdrvMLyfumzIfSdWNYAGxchDFZTinGH
FovZLsikopAbNbDb9CIvSv85AC/fzCyhoo9ESNrT3Wt9nVPtqBdDKD1R++dL1VwW
bBPpkgQI7spUOYuLf+C91EwcR0b62OOLbA9klxt8601mIMxIDbyaOVFZTUBoKjk9
MwbG8bDpo0XMBJiMhbkAe2i7IjiAYiGryX5hbhPtzLBk8lP1dFP5D0hZ7DEsyGFU
dj4GNyVIzG4A7fltEX0dg3NP2kXZMUMwAfGnNYcRJr75zet99BKkQkJXKowl0U2N
lmL5EgtU9p9jh047wt1gBy+ORI2KxOhdSIeKh4ePrNwOTa92fRJfVS7tHY5U80oW
W69Ow7bspOWEILlybbf5k2tOIXLXyFLyuYJrJPpxYFZWM1PIX1rpwYZPQtyJiw4u
vKlzzETDIBgcMCiHTc+6yPF0aAWsngI0xeziSfIAv1omoAWTOIGjX4LsUooHlMEl
aSwkANyedLRLPQQ1c7ApPZ0sNpRB0wl+H6Yzd6TSOhAISNrFfDeG8LSHnz+eAk15
4hwtM0L3LLb5RfgwFTufX8Fw66jNNCIW0wZAtm759SLAkV89AqfWwBN/5RV0SYv1
cY1YasKy3/KJEcF4ttNWzzXv0ZydUXcmkTLEz1SywxqN0LolfR7Pdl94O67Wt9dF
HdhvvdEYZVZVmFnezFIQuMInHtuPiqyvbA7N9CesMNlyvg7teZO0MXsHFPrsCBOy
2o0hmElB37WGqk7zP7vkw600qJ/y+hqVXiTDkbL6e+jqTnHXrbgvcg9HhXWHIuGg
y9ulEgtz3fmzVQigYsRBjbMceh1H8jIN7RADEAtzVgFhTMytkW+SxI80ilroH1wv
vgzjnoL2ga+Ug533ztO11Qoo4DGL0W1ettJqNYBpD+dloG0pDlB0aNqOixM4cbEQ
qOf46p7eYl0euTwCi50f0TGgjQXbD3z745XXkIio6nIi09ws1hj4SZE2Uvpcdi3B
5OpOmNIgVAc1HOAMMjalUwUuYu4n/KHSHx8VYd64qKJfXnU7JYlCeh+rfMffFs9z
2nbOQmCFuK8HMNbMLlBlUpEG1HoGyi+v+WHHDJQA2PFWU09psldef4LKyvRV+3iT
U5G3FUCAifDnoOLnFzVt2YhGSfyltivUxyHEYBs3sKhWoGbyDfRJS11S9envT690
BKGBkMARGeyk57WxfmgfSJxavMI/Tgf8fcQUxuYQfMImllmOSsEuLJSPZF9edLmQ
+2LuVuFLhjeiPoO/lNsi1Vb2zAL0adhbhvFtfUPqa4BPCFuSH9KS938yCbygw8DO
Cd2zjkEi+vqIUxFCJrTOJlWZMut6oT32CODJ3ico04Bnxm7zndrNH8CEAvwEMBH1
hONNxwsJk76GwG+w9Se3ocQFhhFlDyqHEIkY0bOYjavOKcacwOz4toae35bfk/P0
PC5M1BPG7vKqwLDOblbKC8HbP7yrx1ffdemeX9QXALlriIkie+romjmZJaleXI/c
UqxoztlwcRqoJ5L1SibbXlHN6FVWCeUg1Oi2+GhVq079yW3l06e+fP/EI82LjHtB
ZJ5Jp9mUFswYww+xPPMBWeL+6GPOUxxcCTH+KCyC2rWhlQFqbCK9jwBiy0+CkZ8K
GY+TzUrPXAzaBwjb4AX3bkLQKz1ehA+30ttfsM7Jr0QocMGSkvWKUZGvV92W+4vK
pl0SOUe9oHNy/78WuCJpjzn54vsfHK3BMEogLSnuxANVabtHpjaffNmq881qmy9H
H4361MoGUnvvj10Boe2lp+zwim42L0qSUfiycc8RVfXQqyoUYoH0xRperVcHoYtc
7gjStfCD3WFStfT9Ij/pBu3dtWocbK15ihQzzCXRMa3Q2xY8NV16PmroEDQnSJJ1
Nsb0LMHiV2gaA0qpxu/f/CBGZAjcZeCj1mf+t5SswDMIM7PSlAQaz4w33Iwqgm8k
Z0Er6NT/bXwaJ3SHSZmEFXXar4vw+FtJ1S+/wDzcEBHu3QbqVejkDvkDKFJICdmE
UQBaV2OKksgKMbx5Hi8IalTwQCcBLXpR9XMqx+I07vpqqyYbuILTcMMKw18Nrqse
sfEZLSqiJ6dKpraVaocWVmeLcsZ64bGOaNHkvhaHxMaeiNmVfMNF07nXPCOOp2go
mXOFzfGUJOLaFrgf2LwEfOM+/N4lkPG0RsGO0LAzHJP9CeX7Arm0rDdS/MZqyq+A
DQjksm98jr66HHr6YaJiTUnlI5Uw6DPUKkdbOYkKI488KPXL8soBJX77AOKZVCb6
qZsslZFMetkPTvR4ruhTH4rxXKG8TrScduz+HvRDWybBrf845cIgZ6Scf6aQAQEi
SE343POChHlXOtiD165ilvMJ3bAe5n2MylSgt1tAag0MyKNTr3pIySYRW/DADrkW
K/+izQvpIZPndQK6kZt6KGvypX6xjOQfnzqmFnqjFP/xvey08WOXo2O2Ma6FOPh0
zAVRD8Eo5/JzOJSepEbhWDKmSAJlIcFXdJ9DN1+8sNUzUsqD8AbIdz4bX8NpnXJS
fuQg5Cji+W85xqeT7e6EDzpRgsGUusQBMatrmsL9cWzTRuDOaf08HoLx0nbdnQwn
dO//DGlWcHJk74ST/PAEefWAWwtjyHR8xshcak9ejayr4NO/4cGbxa0cTlAd7YkZ
ay/KHLAeXpwjf7P4PiZmt+IUVKByQSCKM0XArqpWP0Dic/X7m5nKjCOfTX7LwSLF
w2C+1wFn54Cn9bT/d21Ey0SVGuHOVuwY93/uaFkS1Jxg2uB6GudTBF+QyPU5uE2j
ZA6cIZ8WhpC7Qlx7HuZ0X0ZRoSi4ZvEUfjS8SicBrTkV0KxOnqwiydsLJ8W8guju
wTjHjVkfbk9qVNunHwJ0PnxYN7ciAeHxTxOkGMsd4S3X91Ty/eSpfb00YNf4dbWu
P/usj+aPnAmZmw5phNeFaiArC8R0ImVyB8J2BwX9vsHrha44aYGavVjGofdrhn6V
x7sp5HmrkQk2Oa3/Jrol9Z3ufjwxv713vSI+mEEtjszG+FpouxikpihIb9KQg1M+
MfNQWC8YYrUvkOjEBTCMuzf3L1Y+BcbQuQ5uvM1y0md/hZg8rzmPwZMexI3+XW6w
S/nT/hap0jiPErXPfOXdCOcRvwpIWWvdELV5QClKgG1WKoKxyclKAD3Bst8vcgo7
ntkPCmrv2xhuEpL2t/0y37pUgCUf4Caf4xgn/ltTUpMm4QHeYwAT6lqk6KKCEzZF
JLcGAXjcWXFZ9bLymd5Upx6SProH2D2iW/qGriQpHxBAiZ+xwx3ncEk9mWPJWNNn
xLpNFa9TX+2BQZRbCa/XhRtzclbZhkB28KziGM6Tlpgs/FD6bNSPU0ahgHX8pvfI
LVtQRtbRRpS5sD1Xpu05TOVL1+C9Luwvp4FtN5sdGG7SSOEaAQH6jcecxNDt02oD
JSBVrbfLs5tXtc0inVDZbAn1VqqVWdhttoriuoMzy5720P9camhwJFzWmCKYgpcd
G0UVM97obthXgUGU9hm4Mex3gk2Sb2JCkTIier+nlOLXKm44ds3n9EXV4tDTvQtj
YN9NmhSfj5Wf3DqBuKdVSzxOiSZRvgbveTeGesqypIxI5eM2inDYbTPt2pyCUosa
0dq1lCgpo9xB3ony/JB+uUk5VUik/LH7AxFoqPvxlcM7qrwN+9BciIg5NFVegUnI
OapsMKQwZeO0K4sCAgqL3tCo75EiRO9DPhfAbjcty5tBAmDCsNgky0WzX1bvTVzy
DIsOeLolWjaNX/ScUpYlyjoHbcCTN8j8noIeeF/DAuqyfaukuMDlk9UlkYdwM6dv
7HhdvUGxDpXRJvijnxMer+bkBmhNYOdu7Cg0FZ9umU4jS7yGpHON74PlBjYT/m2L
sPglZlMlEQJnhj5PY7or4YwECo5wkpBLgfZvgCOeMZlNmWgp4Bvq53Bofhtzt/tb
FwnH/MfmEYV3O78XQtpyWXSfrFBawOHPgSD1OG6DnAs3mPX+oBjCl8XDIO1c+zrs
G9PJ+CBQFK+kTVpRJ2tkb/u+fwBm9BCRGMh49/lzxaVDavrMo7BARF9teTlTBK/k
M1cke5eW1iF/Dp8SEdIaBZjBHynYv43uoY4uoUWRWiAwtpILhALyFvpOFWKXEhKP
PLbqpH00jLUBRlQyLVkf7pnwB5JlDku34v3ybkljLzVmQQAeY5cIxUwnxgq0lcNY
Ack5KCIDBQ+JTqhieNbX6crewZ3060Bo243M0OZAP66HH5ZQ+QDwmGEo7rmpqyRq
PE2IIDekkkexIW7G3b4PxmF+FQCM7T1o8b8wpi6/QE+pSpdbQY0tDWqYeoyeJcwN
gafJAeSmnvIV5cjztLGxwFrqyWkmxn2YCFFhNKOKub8+/qkYKOEjqUoaysY6tLUs
mJzyY6EOy/AeojYrZZkxXMxP4690dl1aETC+0TbIbjoL2oiV7WM/SttsuMD8LJgt
ASi9AYvtj6Ex7sr9EX20r904F6RYieBS4TgZkz/kQAj23Z9H7CUIhWIbIwJKHh4K
qlQz/gDa6jLZbRDtl3g5OGpzbHrnRuREgya3R5c+GrLW3zE1ao5O8PGDlRRqTkpT
EG4GD+LkCOFs8itQYV+rmUM5FUbjnIk4kPV3SHHzevfUusNiB+Y49ZWsagwzvnhM
FKm5A+t8v1n4lDIkzllX6GBDWuuoY6m+UoXiYKHqyZSTHvR6meDO02cuF315tBaC
jzhwr2ib0ksMpiKeIyWJlGkPdQjoOH1lUDmWishBgwAvaIe7kfk6WunPZDKeBq/5
dZZVMYQtGGZd4HjD5R81wMqYNBX7HNLu1UV9myv6be7s5f+2XBPM7hxtkl/u6Lcb
I/jp/LC3JUBb1lEUvSigp9/DyFayFC88sOhRAa/wsaaEAR92D/EIBpys7KFfV8Th
nEzzt8jljR98Jbfe8kwNSrfmEW/eN42thkSyHSrpoWWSqT0YTZpykaJBT8Fw0LUH
4ZE+Y2lYtCKN4ua91Fj30v1KET6wIPSRoFt8sdxPoEsvOkYwF/J0gG4FHBREz6b/
RIJN/XXtYlp6R4OyAxvZ+yFQtezPvMAJOXLWcap8NcUGiDa187brod0D367qsM28
eO1axu1qdO8rDi6jVQRuUBdHD1gy9yr3wdgpV5a0mJaZhssS6K1HmUubR7Jf2+bT
Php1xFK6fDFU7nW5hkCKPhED9smh3wewXjbBlTaetl+t+BJb79PIYy+ssUaxqURi
KLJFGX5gmdPDIt5LD5rDou4b58g0REkodLZvkXAyPq4JrCQ4WGDQAXN9yi+VEc59
bB7TQKTW1C5x+A+AEKEV0Y5yFQ4+Cc7DapOrGAUTttvrOyg9DvPvDADq8vKqMa0V
R43oRc3cRlIFWchMm3pMlA4agY7OzMxf23ZdZozC+qapp0hS31JgUGxYNm/QwL9f
UPLizW3vUd/DGW68tszMgkTeT2GoH6By871CQNL4cewA/aZ/UGdQBua/R15lcCDx
ODLs3L9/+G2Q9qg1SX8nrpARjKeh7e6LT/CrDfstG4hlYDwME1rOnicv+X5Wmq88
ioH/t731360d4j5RXgE7uAXULaYQfIldtWBTpRJ/+FM0O+F6GXIECiSVUsoCXsu1
cXlAoq4xv8D0ewzfR60CaFrgCMzbtavn+EuhaZbXZZ7qV4k7ZxFuxUp6/KlkYxgP
ccG3HZ40IJlo8FHc7yaWjzopGSbqGx4a4V6GbC/DZAtg59M9Jp1EZqbhdbiz1Ma2
1+2eJJ1JnHbMc1bvb8zU6rrCVKCf8IvY401Oh4wbUN+bTH5IJy0nuXKV487UMoVl
tBf91mRdcdTER9OeyB4H0HmBuuIZP4DcwL4UY9CeEzqgSjD49dhSg1Wn3jz3Ucqg
lsVxAXamTAczhocXgquDURNwpoxC7eeEHtvlnlq3fuuN/YqEB4WyCyv+pW0MuMpk
c/KXEDkEpjvsuET23RAtBVsPMUFh/6ZZgQufcA7qCx75Ayxr0B4LqPNiBYH7TtJY
KwYoqFLGjtcgA2/ic7MK3PTqgtmrTTWiwZL6EjaNkhfLK5/BX7d5YXnnzv+MDxeJ
xkJrMmutMVllY1ai9yBOsSpE+lmqlFC/YcctBN8uH98yB4FD9sL4fftTF+75NwBW
j9kGlSaEk+PSP6COlh+ZS5TXtJ2YwmAuQmDGq5NDBhqA+JxVVhY5AU2cayyyoODa
S6aV1nLqHAZbuFxNO5racFLNeykhpC8+b0i/YfVhIsDuUdmSKEevTpjv91K3fGiR
dE46Cty5cdZndYXrxJZM8EILLzqAWOEL6VTPhlk8vOR4boAGsxvrv23hBYbN54yt
eEy7gjHgEHTfhAxUJU+U7u0ZSeX4umSQ6Q27CmQMG533bWDQBcgH7O6uBsONDqMO
8BWkswQ9NJdaChtjox9lkOGlxTM2Lg+VVcJDwG5aKUPMw5aT+iMD/uqFRjBmDJQY
AM9G6UqxQnctQCVZO58BPGDqoDQnBfeMTNbcpRuBYkyTHAysZORQGghoVeSeG6H4
8CKaFHjs0lMkFN6vWxgM82epXNRpcZAdr6NHh2YL/Y89/z8btBZT6+TIYanB/VU6
KxX328aZrDhiTk3M7HtETT35aJOyeJLzGA9f9+CLrP+RXlyq745sDuNmsSFaw5V+
PA9eBA/WaX5wYvDylHHORBxE7LeFeJR7CVFLrL44oiMN/SrPW7OclwF3zZyP+VhA
2yr/f68uLPIYQgPIgfK5J7YFyc2fRvCz0U3Bc6GwA/S/7DuuU9Qa5wR2FWOOjCXb
RA1ZOKRtCEWZr4MtPuylfR0MqFA1qChFhewyc0huR6P5SLMjfjNH9SwrYy0oiS7S
OXoXlj86+x2OK1TIjj/XcwpZ1BqGmWGNLrbRGXSYtBmRd02y+pHG5E/1ojhs9CSB
Me8AoADcPCXVN6l+c/+MNtI9K+gVlL94bkixZpt4jW1+VlylmlCGBAHh0J9XdkFp
Ld7hdw4l02ayjF9ANlZBEOGDV5hGy0NX8EiqLsKdKzGVPQXWjyukPEUp4Q6LnnUR
zp7DW9Zeim+4JpJYRR7NnB0FTz/GJnz1KJ6k+4V+oe3T/mK0Ig3Z8Ydm68vN1Qk7
ZIK/MSMvsNZu4dAHzEtMPf0nf10O/jMZh++vhftF7OUmoowCPslSYN+8BziysA3O
rAREcXaS64NoKOWZzqwBxmBpUfBEs/tH1GERsgH6I9ZmBdEdP1zo1f1/QO28NMj5
uu8E6NKHmcgSYNCZCSMe8j0GGkKhL6oENTto4j2q7C9Zw/0xoNrCaSUlIRUHItqH
IriUyYtTCh0+iR7terBamL4O26L2Cv4udBtw8uA7rP3UWlGJORSBVgPQAHwqMb7s
xVEwuMfZdK0EZKEYoa7uDfCmGbTOEi7rnxid5kTlg0np1OsiEGGnMpwF5Ml1s3BI
+h4cD+SzQ3P3o9tSfYI4sW8cePqJfolEYNzfqAeGbQgE6LkRidHVuPLq5Qnb4umM
/z7hD94nKyiimMlp/6msN/+BAvhWU9GNDxidBp/kNQNdNGMyiHbkB7FO/Fulr9YO
OcNoz6xHfiTO7jDpdLDYIPmY1Q7W/egenq9lQKRUDPvc5SeQ4XxFpMXls7/kKTR3
wfxWxsSi50UBWKeJmAVm3sO4eoNWjKeS22jcLmdEattJz3ub5ZPDO+u9Kp6QvhZX
ImbG1cdDJWaRXlRCQR1g6db0XKTXkN3q/DsDDtLOrHU4KabzgFiIIR+DPw/abbXb
9KytAIuTQH//XHt2eQWcGLa3g9zWnWemlXeMd2ZI5m3d1w6r28Ld0mcP/YzG6rKY
2Po7dBmqdY8PJl+tzw+GHJgso7eQFYoTw22c3h9VJN/Z+ekPA7w4zNXXcv1H2BeK
2o8pVINJHVT06jurbMnHC3o3VL16ZmneTh9vdHzSXEE28az4Hi1z9+LmDgAJyJKE
fOeh+bTuTUgfy9ULITH8ulC2dzRJydZcD1PmST3dsZgpw8I++9VnPOkeRm1tSGom
FVhSl9Zzyju7HHPPGGvwfhHOc4J71/hOFK7hFDBAeixwcwL+DsLzldNsnkbUIx00
0AHaWKb6+zixmfLORndqcou7paRKLcvF5/Iva0iLnH25TMa2e2XJfseUaSo1Dl5B
voQHxXJob49KK3Pyxg5vzJxw6XP3PJScu3Z2Ocf0G6rECCBUtBLA04Tn/riyT87T
G2UPHfvXIoB9PGtJuuO0pjYd6otKu1od/3zSMpYdSiPNA23UyjYIsvN8DMl++6m4
VpSh84RNCnaoxu6AtVmc9+Iw03CfQoS7bhGGY4WQP8Lsrkmp5SUO1rRw0+GukYG/
MKBkZN74ozT8rP0reCgWtJXfPFaas17rAXiMUXP1N+mupzM9H5fh4pPsVvHM9abT
bBDD4XhpxxhjTxlKuyKpfDuJaNIQcIwNKNAEz/xBhkxg11zzEub8hdLTIrS/CmKo
Rd0wSvxHX4a9nKvUNbFAJ00TV15E+s6M6008I4MrKeRk1pJc72kAksXtrwPxBxgy
EeqhyrtefNZSzQ/dRMYng8p4TbPMGh3aq/EjSIVCgpROVnVQA2NF1NXce/ppwBVc
qEW94fbyA4Tynsy1bCG1jbUVUq2aIzid7vEjUrwAOFG7Byc7Up+fjZROpSmfF9o6
5YAcLeyPpQa235HIR7ONVNTyjv4bIc6Kdov1KhzK/hkf5sIm+diygx5gZWlpTxuk
1E+tLUWyFtZemF6B3PVvOAh4+IFBb1IRDbFh01SuDIkRajDiynOlimidzWnMpmXt
NQ7d7zdhLZ8GUtesBkL7mR+Tru/B88jaRKziV5Rq++Y1+Hkk7o+4zuaU40G0dF9J
2yLxAM/QQ+32K5hgEj+9vDaSMzmBYgMPUelsywinw92HrgmEYqZ4N28yjhCAGcWI
PZn3ciie1pLbJbpEaYddBZSfoi9e8HG0sWSqKvp62NUIKQcd1I9fT0wMO7ZXCpDB
Tx4wIoe6Zv8SwlfhPFAYRt5YrHBh7mgAhsoHPAQnDFDd+ZA4PiZsSLyo9Mq3mqwq
8/atEpUMzaRhVIW50ajZbq0IgVpM3drzcjuMh8VdWI2gbe2dTc97a6PMm48CtNuJ
EhJvPG8alL/NjmZZDSjpWihKDQD9QqsGRiJdNtWkR0Li+qMqbljk4wqR4xG2H+ks
rBJ3EcD3PZNPWeodXW/uMpTYgecVTwpZ5vUuVAROwkW1cEnSz3w8T3RB4ULGVVMo
UEFZvqx06jkGjJI0o/wZdvn4kkyNael/YWU2abqaECelDEKBwb09VU4HHWUjlk1m
OCb9nwYQaGSBEvBzUfWPPgFccPgisZ0xpaMqt1Ypjn+VaB9Lqx8ZMSz2AZF0XtGH
I6NJqZfFxQ8MiuymzSmUrUFMJBzO3jbC7EB1RbYz8kZj//LSVfci5tet79a4rQco
+Cq4mLUCjAhQc9xKyWM6IqEYFTtQbP4VamBhDAcLbn0IyeBCcqlWDJHc6CBymRdH
GZ3NpmFKRjNELmj5tIbxpJUsYpeMzVNOCQYwIjLrP6ufh1ZKuNkcqHBAUkh3wsG8
YiuFs/GGvnM92OgdTmVNK/TqvleYtUbZkG4AKmhiabPdSFoa3nudaoX6zhk6XvH9
7hZPdAZqOMVARK7WEdD+qTMWq54+uH4IvWCyGtgV4GrrlN9K6I+W5qs9JeoaGp7p
Karz7RpypRNHZ1m7asYQ/JD25tfwThk+jN2al53MY169fAdjckRGwmtcV0L+r60h
jzjz7CyoOizBQDAFsxZAS6dvdGnuHT0C8ScaSepZvviJugqxHUgIQUu0qD4cw7fc
6aOpRfjdytpMxNqeXyeccH2ZppfUIIxUur4tcdfL8PZXXdfm6I+lahg+6BH3woH6
HUO+ZisO1+wh51k+o/Pyz0xnItFZl2hPZmvlrWkfuPuPcrfFyU7MofdNo9Y1G6zq
kEiKW28FxZpPRc4pbgIXJQzUX92XH7wRT+/Ra+Yqb36EgH8VZs2SM39yduvn9MQ1
A5CYKonrLUocmnqJQOMKX2u3QRZ9f5C5ren9d1X/nTepCfBnreLjfCY/3qu9hHRM
ycjEEaWxWb53DTXRIBoCrRzWlUNgRLFYtx5gC4bFT2atsFpW9KOYTBxHZ/aV7QmJ
I0skkbyA6aFDrV1N4NsJgth3BOt8IVsO2MqK4XD56iVLaPPAqDithdHTiaPUktx3
8ce9JfItsZW3wKqaMb7VwPNlqoGv0lu2+B6lP7ovQ5piAnqui+jiKj7h6wNgZHhf
8h6PTUJbOSv4GVwShkImIAkFJAb6s7Mmm0avDQnnvYEj/IK6Pxk5W4llj2eM9qPB
9FPvbrObvfdMbwXDk+gDrA9lad4xu4yCUZqciCNAFGpetqnrIr6lYW3D7mT3ApkH
pMIIOndnTWHmw0qT+6tyDqXTEHvG43SfF+yKEnSveKEwNaKJs8KP+D8omb0weqZ5
Z/FNO6DA648HVb9pyA/R6qZxLFDvOgEVj5t8R6AOAsTCfO+g+IAXl/ckBeBoaTgP
m+UqcoldPSSOGT51pFvIy53GzXXSeXpFJhldcAmGa+sgyE2uoryp49+HPRu9F7Qw
rxNT+KPh6naXpx1uMaSgVDuLYPt+WoQ8FAxTjhECFjzvEOGac/SwWthOf0JCb6Tm
cRDeLseudJKei8VIcIJDfHNCyFW0E1jExjzTY+G2+W0PiOYl2UcmDoB5QmTIlJ3A
E0SVSgMrBdZK/OQ/obmBEW23ay19bx6CIAod8tDsgTvl/ds2TrP8/f2FJpo1sbX5
96X8x8rhN5cQDe5yEgd+QUsMUfZBItywXn7lWVzrxsbrn+oFI01NhXH+z8YBmiN+
MlZLGzXbhsnQiqHRvOVKh7bjzpUDpOhqWKlWGIjtxeF66tWnf60An1W4LvYTlKru
abQCST91eMGKtCmzPnW3u/a2qp0Zt8hUz0cWCHCfmlme1u5VRxPwoifp94CyJ2cC
aDqI9QJxQm+kR0ibjfYs1ZVirISjy0vj7iLPgH+lm8lJacExfQFQ2ZG3IZfGLafD
NKnMysqHdgkRXaet811lF7nMt2HpEaoODJn1QajqTwJlpagBe/3bLvB+65nRv0qX
jwo2ojE8+7Ht+5QYkYHJjJ5cPpcuF0EE+XWh523L5QzJc+oaFSUHbhQuJVZC9hM7
iuR7yNFs6LEz+RoZvZcuZLqcevD/PbJVSex/zWUXf/V9zHxQkhtOAdD9HBQG/TKs
jQuSHTFmMq44sE2e3MUYNzeSrqnuuSxgDR13TUH78NFmGSPhjpu9WkISyJ2CgNP/
O1Bq6xiH44eygj5jkYLt9ORN+X3l7GBi1uFsShia1wLQKLyAulMdF75ZXyXSFgPT
9HgHCoJ+sWDw5i0TjFueJC7NzBsmmoQvzcojFtMm4xwCHuziV36G3MnLoWIXEp5a
cZNURl+1shfss2KIHuCrKZplu+tX+zk0nwzolSZahDb5ykjSXkKJGwAOBYafhSti
Jug3OmKn8osA9vJKVhC9YeSqgi9lNcOs9RlfD7dsjnUuKUpikXf+1z7D1CCxWgin
fCrlFjU4WIOFkKZU/t9FMEy/Eepn5MDvhgrAZyi+J03tjzBuhI7+02eHCMfDf1SF
2Ejc7yBk4/a3HHRaE7QhC4ANCH6UkVjJ8OYyr2Cp7/cF4YTVSbjF1Gv/Q8R1z7py
OEM0DqyeMXmXf+XJUiACNgsZHdLHx0CXcrG43O6t6SJ137tEJLlJiiMvXDePSaaU
HM1Vst9ekMUi3VhT2ZS9ZRkJVTgsUTMPTDuHar6iY/8FbGYddff+AdchdhLVS1J8
XjFgbd17JfDrUZ01MR8GyE+I8CuXUoEie92Q+sJsO/xf2HVt0uyj6ciCxLFqykUS
T/nnf0CWuRQjT99DJ6wCYivl0lM4PzlUyyFSw1dUCToeicZLi6+wAPROFShZYwfS
4vvc8xAJlXzJLWFRfrWcXCyt0HTi1DzS7tXm4gaX1ShjmagPtmEUSmHL4J7yaow7
LgtzG23i5H+0AUmSZMhVHu94r9+Yj1FknvDlaVVuFQv74606frSCzNrWfZYGTjKl
I5HiKoUO5NYExtmxtsUcqHH+sstQeYzCk7dhhcun/G58nPgeFoPnPpFJk73eZSrx
Ak7TQ5JkZTKTgPgl6yAqxDTKUUSR5zEY2H6a4ahjRMFVngKT0kCMoF13ixzf2m/a
mdKV3HgZ4vFMmAAmb+dC9EKqAfyVDZOtH+faJG5lH+AloYAp+mc0DxUaqlpzciyA
UPSoiVRV8sWqLnXYBoSTNH9RRKFrGd/HHHHu79cKT6WDxN63TztwYuyhWQZfWFTB
MhrOgjVs4Nm77L2z1WHZoUYgTGa3pj080SVB4WePEN0EvEufXN1eNOaE1LPhWab3
dQy6QdAGGrb/nnuxGAL5hIzTn3/q7s/6wyGURyJqPfLN1Tn8B/03kwab1hpiNMot
w+Ct/iAu8p67/upQVxMqMt6y420fNE1bbcXkNqWVGt3WDKmRvm9VCw9ILyzoCAUx
O4XluucSbS+OCnbya3dXE2I27Q5v9ic6gHhCAmEaI4x3VEYhGVUWv9ntUii6gmTo
4CL30/2JxKSmJ/wGGwAUmTCv5h2/Hn6KaRstYAcIuPRdsOPyDizAbDST3YZIkJhv
JmLH5HzvDHgO7icFy0BRFBed9KAp2eLthV0Gt/Zj8KoQjaoIfQQMLA9oabNr0YdN
5bPgZnpAXwYVGKkwJ9bhnVgLXmXCKCHZ+apmqGftd5kfUNvCGn0wYZguwwyhlWl8
Xi23BTFdWsFx6sv0KRIyw+ZMsIq/oMMNV1RjzDhZENA8T3AMVjh42fxjZ+s4W+TC
TQOznQrdyCLL4BXcP578Xsa/Lp1dcum2yJR0x9PnUu/1MbF8e1XEyz8H/XemAtrE
n0WjwiPsB6xv2cEtw2Adc8UwsZgpC2iAcEPDivcGI6AlVW1SudZmP4M1ROLte9yB
ylDG1oMiMdxAwBS78CVzD3Km14LG8AQ6FqFXbLGx6kTrmgV7rwF2ws0LOE93vazU
Zr8JBRLtndkOdwynYTVhOEjtVOBlN0x1bw1Hs3+28WlZ5CU5jTZXO2qBm4VDQKi/
r8GOeCiR4Cpdsx0vXDqf00NY8ieKJI7cs0Hr0DoNDHdMpnMLEOobISlwzZft8iGb
pjWiZU3y66pxtBpXAuunp8V5MTbs7Hyn2EJteJtCAeLtXlgk7zwl+kBfBgBNFCr4
83kFhGrJ12jIr34H+bcRQleHk9gfERpgrQGWWryGDDQ8ccEh9k8zXw/vlE+ZEwUR
N9qkoNeTHDYycXSs4ucpj8K9U0s5DqQoNHDaM3C7IDil4LdrGet73CdYB6ZFmQ3h
dAqc/PnC8Q6AzkkZNkhAh1vPvthm7w/re6xpd8NkFYY1rY5vuOQJ5LtKa/UwMLEP
8jd1AbWzGOLvpS/iQQs/UaXNRoTHVUpcqfYH4w0p019xEzfxZ5B0BZfjTncUAWHb
4Ztq4NVthPtYQK+B6YYeuhF6kvtY5WnHwOzEgoY3OJGO8EBxNp3ncZWIhnq8FQx0
oE/ntBYrsdQSH434/IqJWMnkbCBzLrSgEG41JzkktqItJ+U/z7HwWoS515hOScbK
CBAu9p1UD/G9wZr0ah3BGpaQq2a6Vp4dJHb0hpIBHef9id6pHHu2GnTfrdgSh/2f
bTehPhkMoYNVU8ym0LShUeCKsFhg3qElj5vgDqWXchEtzIGaC9tg2/HMRZkdF+U9
cE5JHNDJkvQl9CT1ABmhJb/gerPqIMc99Xj1sGQN5Izj1bWji87arhmuXzpgtHXF
z1gFt9PjZvmslWGzBbLLBHH/CTGXcrWYCdY2Bl8F78ViAdio2h19tZkUPFh8Om/7
wVBgqy3n5mrB8xiH8oTNLCCBnG+QrnF7hGQHOA+dUQOVmQKDSvHiNa2Ys2g3p4AD
iKYrvDdpggjE9VHB39YzpRtbIVtIPpfIcOZiLVpF6wYU4b2A/FnzXijYQXpLLMUf
0mDs9TaR/0G9VEZT87sUaRKpBRHzgdxrhEUW1vXvU1YL482IEx6LvWJywMXn6KmD
js5fEWXe7Jf0Z2NhExARiDlULm4MWSwrYn60BQi57/fuLvDtmBolQBIoSe00/BAH
Gzlgz2juqKMafLXinKbYtXd02nSTPv8fV2Rejw4e4yxcWoaOQBeDWTP3Z5IL8uzu
ajHMMnhBDjcAQAIhWd0O5Ty+n28SqZA9UY9cBg9EQ0F85ZurAKm7A7NgJBqyVil8
2ulRgQOxsq6O0N2D+BP9ThVwFN5vQctNVuK3fJ29Lg0Yww+pj2vQvqxd/uSNpXVe
PMwp/yS+Wc5K/Bf27kfKJHrDcfCR2Qf5X/MIacghYhvDJZLsYXKrhKhKJu1bvuQ6
SDlOLF4Prm9q5G2a1CFQxLmLtEc2LKpkGLiYjnj237QpzJeZKdiSFuwocv+eDG3e
zHLaANebzR6oOsYfI7V0mXwMC8Kv+3NxzQymM4JXH6670h00izndfEGXME7fXO4o
tT3XV+4R6DdCHg+AB3WQIQ+4XHIA/KK+PIqWwe3zQIifvA6ZZh5ebabmpcOKEP4c
BRLr8VwKiTskoYk/pIAEpET2WqVg9TlFyJMWwwzW+D4gsLDYzhiiL0FS6RQ5SzoB
ORvZslrMgtoalsNu9tQfWfFreIT6lLwfsPH1jtt8bdq8NRfj8xTBjDJFzOvl2lZq
Bd8FEpaEiQpmcDL9hFhvE6KDYdrCIlYSgNy52RifoI+1vVESrRPr7wqtkuyfNZ3a
LIBZTQ8ctjSQf4ZhmHQZPiMjmdNTVI0JMvqLrDGJVgy/aDur58d5S1VD4yEqcGKf
HEi3Z/UcRw8+c3P/1eicY/b7ebW86hVPt5htYoPbeu5bSZW2DZvrNDwMiPp5eQ21
dYnWNneuZq9bVETAsT3qJBVcCfH8HlbuuCU94fHtj29VJpmV8YAHAIfrwoV5P/sb
AYgbztxjgrBADmmDVaxhrstr4++BxGyRHVihersgjgXhAyC7gv3JibA5aHmIp1/9
FQBAwZSaMmAntE7Nb2panjz1WyCFmuHvAXicKJ3Qd6p6M9D2tXGngDxaV0YQ7GHb
FYl2bmvyr/VGaB50+ehDqYoZvqnVxIWZHaapgtJV4ZCg+hE7TutR7bElGljtyG31
+4DX0SKLmpN+5sxkE5ERN2wbukD0+U96CTqE/fGQgqUUvXFP5sdg5ljJ5bYtr0rQ
1/+3/9deb22Nqb2fpYni+m8emzz0P6JzE+rQqeW9v3vXHlB86gdG/U49kQhLU0ha
ycs4gnsLodbuQriKkZi3/9vLzUEzCkU4iGe4fqjR55B9I5HNlpTPZauRYDIrn4wh
2S2Wdq9MXGlAbwAfyrd9cM9CuWhSxvg17EO2HLm8DsqCSuDsF0sgRXFHufnbgdhj
1/lmNi5U9uzrTw+RrarJraNTb/zEAGOPld7clUEd0Icj6DL3Cvhot4SUlRhXEs8u
6ENCsIhbFqmXc/q1xMuyMmCI7Td/TIy+AXRdrahvmScR7w8sXGjhd/W6RX273IML
2iAsXTO32zCi4AchvH/XfIx25168xMwCjZahWwhkvzJfUShkwh5yLIN88+anjpOz
YUexBalrxm9Lopu/X3acKMngkpiBG+9MffLattYuf2mVx86onXoRh0Av9Lz+PzBc
YgRNaJYO2fDTNlHAzfrEGKMNSrfdcmczglFtUjL4/5T/QxRsblQekCEcaC4/BUFp
9PP28wK4yctJXwYIdCb3ELEmXfQP+PbwtBXDmjJg0y00pVSlUhb+SdQg7nilX2da
tdGkJqXdAimHWiV1Pl8UBRGqMXSoBAOUl9bByCcru69vLD9VvrQFDWwTYVnTcJfP
xCFMPAd8Qy1uoPb7U+TRbOouw5gRMOG+OPoMHAPyHdubsezilG1Xsuwp16Yf+hNo
Hifvv5Wm4g/e7KAetfX83t1ww2Le2KCV44diU0zSY7e0FxQLBcCUdtFwvd+va16l
MUoDewP9hkDHlzTzj8/JCXBAW1R9i27QpngL7ddN8pB5kQ3AIeyhvJ6pLjIPkZV5
xp4OUTbGASlmzx0ili9SZf0LdYvLFN/lOTj8CugrWItdAkVL+FMq/TMCxDw6m+m3
YXjPlaPu34TThI/b0/j5n+RAxzns/qDuDQGGkzxNfEbw1H9be/YFT/K8MRNitFfF
9Pfnt/L8LzWimr/paiu8RaUvMtFJjYfF3xmOJa3XJdtcDIrR/6Bi88+r9YJOWPe6
UThmiBlGFmybpnA/VVRcDNHXwhP2naEbaL8bsUQAlBUc8D95V4ehxI4XLea19aEj
jUgxHyIZhT+IRlJ5hWi7UPJFqAv+py3sw9y+4LlC95FqzypXx9nZsEi6tDptQcu5
C96P1wrwmnIy+9S24S59iX41NSz370HLaihkQUSgbWjOWhKxd6ldJOp0SXQmOXM7
T7y5oC0UQ2T+LZTr12ys5dlqjvh8UCObFHTztR6+TeBU2hOFG1+avBxFOsEUePKA
R/XNAlrGfa1ztkYi8d1hgpftk4Bpw43v4dVDn3lOTD6skNUuSCg5+COAnSXVj+Sr
sitmHy3IKj9bTkww8Lvh0HujNYAiihzkoaiPppbKmBFoUpuzNgBwLDlmLD8luci5
aqo0NDShTbN60VwWDVFEmkmav60EBvdJax6ejYjFKxNRqH23nr/6eRAZaWpYh+qB
Szd/OH1fK7iAVzA9IJ9k5etfJC0O0bTn54Ojwze1dpmlbtdnmZY0EYdNGkt/k+zV
tqP29Mnc9pjFIJN5MBkBwx32pXiK+uPPijtFhSOC8r38oExKmyH9Xh22/qw0GDOK
qFHj+b7GSItyoATiZLIbLG6mqFJRf2hqY2N0fTT/7SguhBtneP6MhBSYPq7SnINc
4MEN1I6yh6/Iv6IQAJbGO1eBzJEWdQC5V1Zv6gEEuOC8o43Yq+psGsEXPpNN0kxu
zc1Yj3z3nZ6kZ6Ir1DXG6inHWYqVdEh/9GfhSH2w4/hPDIs5+E8oq3C1260SVuVA
FOJWQJ3l6z5U5YS1zLI05J9oD/J+P6TznbbK/Jt6Bi9gOn1c+L/Fn3DywNXQ1Nwr
/7U/yvwK3YIG2nzpCRPn0jOxC/PPk8x2/Z73G1uD8bquC2SaHtyyIfT0RSUMEVug
daV3sofPBIqzxWgslBFGp+1zE90Zr62lznl9k0pGYN3BLjGdCNzmQApdkiHgJcSd
CFR0LD2+K8ku3H67x+FTEabtVIDmOjfQXXoow+Jf4Qampbs/jnylv0A4hoICFokN
BZ0UXASj1JaOhZwldoUqbfSaitX6saFAJdXVpjGD7i8k/Bw5F4Kq5ANcXzt/yh2F
yoqAJZTLX6dMp/CoUrYFShPGkyd+MMOYMGlpMoLSrqJzoSCduAz+z9e9hmCaBj4X
/44s2IF9LKwhtiFb4Mr+SORBXno7xBcyl8T0IHmEj00hnh/FUdwk60vh5N7hqXz6
MaRY3pMQjaAuzIf3LG8WkA7nt9NX8aRTaDOz7RrORX5VicUvjSQ8TLGxvzNlXAPZ
ta+IVl+wDuQ+x4S82vAzZZE3FR0X40JJHvdgUa5byXPWY/uTkrvBn/FDEtv4hYqG
3QjMDw/wETyUR+A5a8hAPHiJONt9BDYP0wloQh8bLACo42rVhIPCD79WHxIiXyKy
RrclJMjXTPQUugPVsTCTp0pfcWXJBJmNU0OGWE3brAb92ts7QMiP4C1CdQLkpoU/
hTW3mSYQ7PUEGWPb9nUDkzjHoysRQ72ug/o+WjAgFLvk81CJZkuzwW0FmxAt+nfa
GLfRPpx8n4eFDsFg0nTxxwlCXSdD0pG/9jYYSbORobIhwl/sBCz7jU7sTuObIjwo
Ttbjrrm/njHcLWokcEu2GwtOd5lO62EjRxEzyZ5r/WVCVOVeCFPam6bHIMN2XTiO
fNkm3z3W9S1jp1XhpbN3yklpx57yuj7c57PKUoJhcJH4QGjSkKLQ3QjMz7nfohbB
HznJzllchJV26vF5bmt4yBsNXt/GRxsytx/jXl7SYun8BLA3I8lP42oT3/udwRk7
nrpBcDaehhAAx1n9hBP+PNXzmAQwF+ZwbRuRRFl7/7M2R3dRPlp6mp9LLDJ9jKwx
4VGqF4MlFBuA4wQ+2zTOxEN/Wbbsu1lE0l88kSMLZ+xf9GlVKTu+v27A4OoSmc8c
Nc7r5wAgbQ82lA2BBMvZEcOpDzUqmMJWjjidoEWARjrsWMhngAKKaoLwLRmJ5Nmg
dfTd5lzVWMrdDi/aNvnRbtzamna29ZlNYCY4cH0R/jEUD2Ve0pWQtJdsOp4bXJvq
G4XILsNwCvqoF06Uz8gSSQNHRjIj/YJaYB8ZyiC8+rtK5aXG4twm3O40QzRLkJdY
fdqu1MXjLBoxXxSKqYHM9kWEk7eD2f31QigE1Wd/lJpk2WED85uR85B6KIFmbTqe
N2k6wmQ6mNkXh5G6IAnzOvQfWUiqtj7bViCfzHCUTrYIzgcqs8MprY+zAoZYV+Iu
VJKhAMWTnxGu3EHBo1YY3GNmvOBYHEnLxltC04KSve7YRw8GDYElE+AZM7trfbMz
s0HuQd9Hr6WgNVgtBb8wVg4pYSOkZMQn6yIghchvJanLd6NX/409ebufKuMPjtZo
TrmOiB3K3++u/6Mb5Fp7Pd2EJSwi/385AJK/S/dmuHfSja1EPCjDXK0GyiJFgCCf
chjf6V+BZLf0+Mky5OQ3kiB4B+UhP4AJPIMmjI6HGySIZIGme7gpGLvkQMTxbw2c
GtsxC8mKl/nQ7zS74ZgJr4UynCqaZIByzCY44Yj9FT6KOKFe7MTJAgGX0VaZk4uX
4cfTxu4FoNps+wHTZBZPBua9m03Onu4tfCiLC6Tl8XPUl52TAoicNrHJSuqfVLda
MEcCc/iAPyCcLmZwdQ1QxSpXTrkQTHooo2FO/HaiIPz7dKZk2f5uTAyaD7xpQD4h
T9GeOdXQYRVSi88Ewg4zvKF/WtPDJjLk6p47REHgB0opMW+1RQpvM0Z0Yrpi72IM
EVrBahrhD5WG+0MT9UdXz08BwXow7oHOzdjqyAjjAR6NLrS5Al8Pp9YpyG2tK+eX
c746vV5t3+6nYF0V2A2nnvDLdBwCq0dqbI8qNrXqL36VaioYwO4JWmPAKXPmpeVm
aD8KOeoRxvGfYvTfyK8r+F9kZPSrelbtZLq7bmESTZCL1GAkZ5GC8Ijls3+pJVYc
1i2I/LB0ufEsph4TYz0Wx+14VJ0AF9YnAxTFgkvCX+ILJMBdT2zUG75geFKFll4b
HRG2GVB76esmThcLPHP8zLNN9hJfKrHwG3d2iMF+B8eqS/qxCJcYCHUjes93I9bj
rxrAwCthcT42XBw/R7jsjhr7JnqTtI0QhNs6IeCmNDhTwVNlf0gbIr21Jdvn1GyC
RMUb0iXT99mRlc7qRIGXnyM68o8MRkV4v0d+FgRzq8I1AF0+MBzch2xKYOUDgCGw
Ym2qbEOR7IbDwkjrNT/xenoSA65IBo+wB4U1ZUiD3Lo9EEZ+nr7mfGLFvpe1JCYV
cgUoohhM2HopVdwrALoif6IjczdYCJbJ/BfNV1pkpDReVb2MFiibr/dPAtTIUjac
m9MkEp7bkigGU3VOz0cD5AdNzQ8nPaF/JNzlzZ2sqjdFAJMfPpfHoR3S7A8A4b++
uqJH9JqtTvmObw6gPgAoWTKIPogtOSNW+wKlqxLdLzdujVZ/3nWgTDX2Tvh6DIfQ
XVBtAw2vdYg0HMpx9G9HPUd/RXYy4HO/PVRaC7pcd6N3CrusV9HvKPHL1hKoWRlm
aSCGUATFNdaIlLSDmPUl9UGsDPAeMaJs5bkQ68FX+hQyxBi1y2IdbpJxit/qpQER
Xk+SJyGEPkp6K4wrBoihmywtXfKaLsfnabT66F4YTrf7QMxnIt3B4l9XSdpaTl9c
FA6g6tMK8O3fSuXNenTtVb6gDeNafxp+LCoa0mzySRpXAbrOBE642ZofcbHHXsvY
tCpsbwii3y3XXMO/INUt3wguH8Rw+bwZyShQr8AU6+KZSWQP4eGcU9l2zCVW5TQO
je8bRfHwa/6OcUGLN/F0vIL4db9fHGjecYVINBrFsp8HlZW79hy4roFYUic7E6Rl
9tPK5bEcA9536rCZUwjeIaleJSm9gRSwKzbN69GKLasDFQ32X+lZvXrMMQNZ4uVj
6/65Gtcx74MExFSiRYfRFsRRZLijqrNgaVrO1790QoAAYRve/U+YPcm1na4rpUIU
kPDtP5aAHYbjDXLphQpgn1SRIx60qeDPJLem3RuQocm9eL5uBKRvBerg0eKC7OCC
zbg7HWSidhtm3WAYm4OE2nYOJfviUd5OjCKWJqodUa7ygKmzbT/VyKvr0Jjc8a7T
85q23SIui/JguexABJbKkjZAp1ernUG4KZV8/mYAC/JDzXFVkNfdn/feW3rcpbw7
Z/x7uC1Ko7AFOw9jdYK5yU0V07+BB5k2Bas7MF3VmtHmd/FGn9vdLO4I7NnhCy9Q
mxldRNodizX+PCdz2qtuRlsSQJuLGwM4Br5GVYD3HG6A8VU18GftU2h+G/p2SeEl
YR8I8C53aTIdv3pv9M51g5mLu8GiLWkxPOqvoVW2sY6qHU+TLCDYWKHT9SPLv5IA
O8ZMiSQHiQnb8eBlUqRaFMAr/dnY465xqn+xoZqvRzXh4ExKDPmJtpDmmNwhkL/o
5hZP0b3fPgdD0Kv5mDbjZUp+GRE0sEiRjOd5NMLBTgKyWe+AP9ilc69D1EEfeuB3
2Qi9Db+u9JnCXQU2du4neWfUXdg7rdab0Svq5c2xZmFFne9kmxEzlkDpHkqqEumd
bMgHjP3b96AHvScy8oLvgmbFTLudVkZiLJINzt83nzm4gFJ6UryreY/5i5yNVjpq
uY4RlhckrOcJk+eAsCgvY1Y4Ue+Xu4eJqKSQWYvu1J1PWU83k0XBifQ923gOluLq
N17PZ0WIGAdBdJVAVSsm1MR1W1y2p0J0Ft0tnW0iJZd0ryY53wuHDXK9wt8dkxay
Q0UAo9pSd9l3GK5oEQa3r2l52yybRxyFYQOvUseHxq2SoS4aufMUCSEiLsCRkVNt
VZwhdgXZiXqAj2UjqaCjlquO4NTzkwz27g0/Mckww22rA7JPTdqPRLjWMBB2c7zH
/vg0JptLj6mCjA12fMBmJw374vejLnQ1idtqmXrdwswkdmL6fF7NG2Cy+Mr37czf
/wX4f+jbCHVAp/mPXZbGQhMBlDeiQ5QaASUmwyAMDl9Y+KHPSYZzYj8nWrVRyZg9
5k36j5a9mFKn9IMohgbP3J3VvOB1yK8Wu5LrFzJU9xL4chGPvmf6kJGlcdUOuvMk
okJJU+zRfQmEv9nj/YLA5bRtu5550txq2kbcxzaYHNYInrFa5KsOj8/keC9pHBJH
xgAU8/lCuZ6xkndNnBlEvqRyFZWgA5LSuh6cwt4TNbZTW/ASEEHkzk7pJtHHYxTL
5+O65vDi+2j5NKUuEuAIjctS4bAyq/kX0DOTLypJAwOpkRsWwG6Wnu6J4WahzMap
QHSH1T0icR0mT6kP8v/UvWivl5FHqjfllvPI5KrvE/B8SD0y77PIUqF5vuqIrGIx
NE8w8DAp9hcSxwDbzD66huJtgdt1yjmKap6HF5PcfLv1bLl/tV+jIgko/UZlJNGy
qZOFSn2cyGiRz7QUmQ7krlKN0gxnFLstKijPTwcWbcko09TG4BTVtlh6Mz0SMR11
I3LhfQUB91QLxhKmnaddu4BPYSag/n9JucCFt9DsXfcolSlCX3OydLMzmTddItva
NCFJY6VGAXetkWmFy/C9yn9ZNNmZob1NrW/bt88IvaO++SpA6nDu2zJCj76GNWaA
J9Rk0CDiXo5i2tiNWereHkFu6egZ95tH+eeFN+UbW793aJyEjrByZBYI2QgU7of4
foYSCHxgoteYWM4J1w5D2SQblVkR4LSm/rkDT8mxw9DsWnAW/QCSO4Z5Sq5J7j3r
H9K6A0lhlNkLvAeYLqgY0/tcXAkEMEr7q2kUNbiaqL5QLe2CiRPR9Qs5+z/f4BLk
vN2XrrQ/NmB8lApe7V9Iz2Qb6fhDdYjqVJh8r2O/J0hMV2w4mYhjuMfbtST9gmqL
YhSH+Q8Cuzzslwd0WRbGjy1ehKtiDSCKJZQSeRxbjYgRCRIUG8YqzDyevTaDRFPQ
SaZP4e3MPr0IcnX97PEyJ8xP8u4MYy4jDUg8IQER9dBSJkLmORSe82P/6+gPiAnM
a11rQqqgxfrY/PH18oFIcYMWyIFNU9MpbwYaFeMSWNAPVE1WcydvWDvQxvuOkjLS
3ehL41H/3gMexRHDheCmBHyeTWi3OCUpknOshwu2qeJovdv2uJPQ5ZmrUzA24aSe
DYbx9EX0yV51GZawIHST7Bkcxo1ZFgoUH8FKLYDmhFsx6JABKqlm+po0jjOjqzS6
UZNfnTeB1PUqmTYmCwl+z3zd0SVDuMWKEC2/zPek9Fg8gZGxPLsJqSNxQbS+t7HR
GRLYQkvowERqff6d35nFA6dQ1TnuU/Ovd+URE00BNvnn7wM6asSnwe8Bh0s7I0JC
vNuCtnIfr2bHJDO1nDCopmFAUgvWHVS0mbIUs+BnUzHxmCeLqu5tHy1PCN/36YDd
qv1DhN1p9oMIF8fXseq1j+XDPI6Wt0aGWvMNpjiAbsTYJexRGOj4SgPbCq57ARga
9afw9RV0wsliGL8eUPeYtBC25tkOKX5NOkHy6Ajh6mNq3wOGXQF1XblU49MpdonI
3rbbqj9QFEycZXu+3M87BQFKrDNeo51Oe8+BKt3NHzoUv3/Goo2YjLw/IHsBI2yc
XUhoBe3IT/pEUlsDb6b1a9HeRW8DmZa9ijyzJzZCnGWM+F+L9yVjAqKGdGK4Y0vk
FkNNwKIFW1NPwlDQcvhlUpgX7TP60hEZPUVRiOghD8h+/qqUPAVmWUCGAmqxzza0
Gs/GVBCa+Qdk/xgC/IoeTNGOWTTTmvdB3Dd93iWSKauFjDz6nEfj/EKF/G3egGfP
wLVezhdkVI4sFO2T+zfYer9Lq1kMyIaSUThTZqo7r7KpbBPrNJ0gH6bruBvrlIh0
X/i1IpNtDWhlgjYi3ohF3mIO9n/QmKU9k6S5t5pq2HNLNLVmQTpwuU00/ggvSRc2
tXxWgUaPOBewTTWjmT+tF3q0jKHXOb5nZeDLp3pUL+0SYM4OzmpDFOvSALkpgA0h
I0aJsNZuWm6Ye2E9ophi6hikmKtq579XIaPDSNKIaM0V3f9zpRr28wkXoM+hI8Xu
ugAmwnkc4er2mTi40C1+26Pt/ZKEioyRY68dcRukb17RTLWM9egFh3z+5BuWC2VS
mIj5bMA26vD46J2L6Gafq3PNReNPjSxbiYTnNNVnpwK16VAUqR9kYrJ/O0ky0iht
NUSXgsA3N+lMbhMko7/CFouM9UD5dmVBFRgFSqtNWK9MAvWABF3RRJ9aWsberoeY
N1ocS8KjUPbVhpNQlaWaIjXEiNnZQ1+7TgUxex/pKwTwfiZETEkIIkbM19LqgZFl
01x5fDdxiizVnntzvGgihS2aoFKP/nlTtt9h20kONFalUhY9vrLakN7Nr1zkaFO3
KzhaqhrthPlK8hXHSSTwxRJGHYpUzc4pMhhMgMaYE0w+FRJ3tUNMtWpScg6Mb1/2
qDd0xzReQ4sxxUrzIJwHYqK5XKuCnNitJM7i4i1Im/9x1GVakp75WfKWtpypf//Y
Hba7NBb1avhITIAdivgfaHm/awEapMnF89e88GqlCCXNbCyO6REQK6emY3sntefS
z/9QJw7LPnvsKlmZRMeVVYGZwpwqF56+4jm0WrV12StcFkmeqjIXVlCczre3geqQ
1sRU7/pJfIxHq/zEyc6yG4ivumIz8ftJdfazWHQtDa2Yl+TCZoMVzqMrqI6cgnjA
UBWkLb4sLuu3m8rJgPTpZqMNtDWGV0spTIMzcEoL8+lemIGEOQHT2hBPidtV+ZAG
Q0elhLA+3FIXqwsFRv4NBrnHWN8TsfsMVaDcyl2eaQz5+reoBOrUeNf2RBjjp/I7
nhmQRWs+b6Zg+VXjB5CKWj4zCEGzXHMmiqyzjXbj4wT5OTOayyuBmoz063zNsdos
xhg4G/O6oUJLchjtHm+n51ZCyeUPvsDDPwWYRtAna13t0XoJbVt5PLfm7RKGzoRI
7eHW2XXhkrussFqAXmjin6DerlW0XRuGejbnc8/SF5Lvqj03uJOsMcvSe5MHOaGu
7CLjLDaYsHSXDowUVGFMb2fXhsntM/0Vk75nAcl2LEQy5eBPpyew9N1gMVHPE/Li
SzJnKTzthQZJxbs6px8v1MYjYg9xrXQk882f/HnQosaVzjhtYFiwvBl/3N9fWZ60
nle+4MQXlGb4XfVt0vWYH4ABzYZFfPnCJlCRlt8aXZrr3O3b4fvyMgLZAhdtRdwF
xDMtlE9wQ+evrGqpStwejwvH6ItIpWyokzjqNGPdToWEOnGk6IaB3ts1Vl6YccpB
9pRNicogR9EX690z1aq5NqZIkWRs8mhIQEFxnVmvIFzbotUPo9LD5W9YwzNvSWAN
bBp92FiOQrymRGV9IlwU22XGVGXztfee6PHKFgcz1CJ+sYgJ3IV6EYhcTEAI449q
dQ5MA9Vkv/uuy/kp/GkVptmpgCPWUSMXHCRCf9KwXXPlSPR/f0c1MuOtDMDSg+/Y
nM/SqRkHq+WxJdeoInV6PeRIcuenaLfO3rqLhWZt5qkOYsWkUAFQdY/AA0pbxIK4
3HzEVguMlHrXpjxgGpr081SnXrV+7PmJpWOOw8ZxABrEvVLDEHmGmdygPa2V0+0h
NEUN/UUW5odjxHXXM5hWs5nB3oXlPnig1ECxhp+yTOTfOD5NgpbvQR6wIevmPKKT
oUXId34nNTguxL1nbBvb6kvoGkEs9MTjebTsA61M7s3VonExu/7M57eaYGCxjWlh
mNZW4dc1vmukRXYM4482PIdV+YCHCCOISOcHn8ogXEvu4Oh8QoyD1hsfDqtF42Sk
pfUQVPFfN2ITG31rIzGzQTyV0RQdb2SQgr7KyuYyh8fj8AurOYFvBQ7+MpDZAjPR
eK3VDDfj5x2Wh2PuRrVg4sLSTArktLn4UXQ4BtB4EQRHxxaidkTkGV7xp0MAfTay
pmfZBkUwwMG8HrdS/xDxvv7pTvRkL39USvEkK4rBkEAN7VyetMbaLhInynCWbl9m
IVWEEvQDGa4QTdYSa2UShpr2Qkgwrg59CHjQkud//ZLq6xrPeK8tiuYm7UP7KHkK
PjoP1yr3TXyQAtjiQCEYNU/OXfkahgDSlSNJUKPbDt/XWrN3FTdoD/Lrr44bU8Pj
H0bYRZ4v9hYwRq6AkK/pHgqBY+g1zk0EtWFdfN5Wr6QDxLem5O2TMJLye0muPcka
8bcl+3Y0udz1shYOF8OinoZ+SN61x8CU9stuZGfZbpZgeUkPog30mL9WQTCcK4to
geEVGOXGckeP6dwMtJ2fsx7Vds80mE4tjFv5fbD1MijP3pdhjrZgB4FAhnx86LX1
5NjntLf13v6P0taEysNwVcMUQCD4jUGo/cJcmEnx9M3UNWeuXUcGQYRwiF5Q/ewN
GY3qh2Hc/teeVXKxw8sXNrum1WJCZo3Po4rQ08E7NOtv1O9wEwwhY9KGv2ngcEH/
awtURAVRkENQT0xXPIDK47/Jc2+uGpAEU11118HzYRQZ1NDPjg7ZzNHxmaROOTM4
XTK4NUnveMKzWwPtRzpXacZRKJgCyw0BoLrqaROb+IyiUoy2Fq8SDMOVJMGmzO07
AueyeyRXNFr0eDkyJzKZPCsUaXbde4EYnXAe3i7zoywEIAscpjb4l/bR8dlz4NIz
eCQ0TOBZ97gCXo5Qv0kLwFn9waNMQXJnUil7rn6ZTi4pKtNEit1eWp7R9QsmojzR
CpkG3AaeKm8zBmlsnRov4W8AfjRz5/k4aQYwrBAxEsJxoVS0QXl9WNHs2UCI3xt0
CiiGx7XkegsaEOUkZ8Qrjg+NXd+T/f7iKZy5e2oDIPLe5hGCrgdpLigpjHjLV4fD
ShRasGo4KiTAeCiEK//KwbLb26dZjX9CM4E04TZyiyzOqkAzT862G0DFGDblDFQ9
CkarcECd7pJqd513tShe2PmiPbugaq2nUDpqCyyvcR8RCSXiZ+Qlw4sH+sFx4LdQ
jTeU4ErDMVQHmVUXWqRb+iq+SNu1jKbrdiZwk2udIWhYH3fIVWzkzBzn/LnHt82T
Bi3Q/1oXYAoZLlznMWYfXyU5UGxbntLS8r09owXt5EuybIMWCTUtV3WtldGxm9WG
+rW8R0Tdt5/QF6Y0d3J6r5efgXjP8VQoQBqvgWiZfRQOiKNW4NUsR1zHy3Wom0RJ
DfQ4Y/itNgicrdAAg5OFfE14oGgepZfWA3zZ4yQyeZ0yS481t3/o5EPXFIGwmUkd
CiBtEFTKbGF1SCSKVmcgGFe7jlw46ZErsGZKRas6yd6rxOVbF0WnoSFd5B3RAGwT
VLVI2nCuxJ5gYwblVLQr/5QGDKmZDKTMQSGDFpktarjXzfDy3EjWlLtclVYY7Rhm
2KwVXHjYAwtp5MVg53WuqLE/4SWt1LedoQN1YeZhYTbrPBIHl3BllooyPd2y3gOX
luvi50akULDeHw9i8Bu9JQs1avVTkbjzCe8tKCpUeX7WXg+N5Voy1zefCGCt2I+X
crcvMUDGfLFhTS67SYwNB7VzK/pkI+W0bF5PaFouGxM7soAqyDH2O5TxM+WvgaMp
PbUbglUko5sVjhYh7+KZVAnN6h2Zy8LfUv5c7PPWztgzahHRRGRjg0yvHlRN7wtt
/snD/S3Ymuz/ZSB/A+sGqWm8Hm5jXJSPlD1cZ+F3NnPhqkTzx/RvNgRQglHTR2zv
0A24KttB3TGv/gKWnddlK4BdVRQnGdhaE1UNNy2gCPIC+wDOXIm2ezbiHbrnBt5g
PLHwWV2ELO22DqFLtMTIXEYAnm6M3JGbu7jAw48ZNlglts6qhoH8nIt9y8OMPW+f
mDGH7Egr/EfXoLxqZ2mAC3w/ekl+a+C0s/E9FIsL6ekCRyjKtKCiN6gftTh7dYwL
Jm5xFwrm0wqBTeaqQHtEd33l7ZOrrDhFbkWPQjXBwgdNhFNotCUDJ+7EgpS9K5UW
EjaaBEE3lTpEmW7BVVR9WBcXtEYWmg7ef5fLPaV5s462mk4mkCYwGP366swhILne
2IFzJSBr3wSMMCdqUQye0jWZtgafg9oRzn8XkC8bsIxuCrkjYWnHo6Gnnt5pGn71
QHjm5czG7BgR3t4groqQjn0VknZhAYS65XDMndVIoaidqvAAGiYJbct1D1kucYps
It8LuYmP7YYefz6vOZsoOB9Pw3DMph38c1GTE+SCApmuy/aiMM5KOYQyYt8AZ/s/
Sl6e0caWl5U4yKdjG79lmNjcIAKZyvg4CIZCSkJ6CrKtTl6D1985y2854sBsQeEU
ZwLEolwr4BUPzRKzjytNcVl+7qdATFJ9fNAnO9eOO7a/frznGTE6iTi4Vn8xVtoq
iy+RBAQo6DAqDg0u4Z47nz+wz3LhmWpfOOKxNiPCjvP35cCjl/xCLqGBYXYMMIgB
qJqFG4WoekIJutTKXXYFRmRHVq0Fsv6cXpFAspgw41U2tSnqBMFdnWfrTbcku2JB
NXI8oMyiWvAYOdpNXQBhtZRuHhiTbo4BbgnpK9mIlRabGwF2huvBjc9w33h/GKvT
JTOFUwBw1fyEKnXAQzmdU1opg12rXwda6WMZvz+XSE+wwF7n/kuLFuD2cJMbfWhq
yIgJh7HUSvUz3qBfh096WD8npicvAAK35CxLwJPz+MU9FCLiQRtcTXSOjyBlEXGx
Y+jAgxGI58brJ62nQqXwhh/92Xp+fah07el9B06oo4dzKhfsthzkvV2oIc8WFYFU
0IoET0F8dlRydetUGNRDTx2KfeiJa305ra2Atk9jLEiSxX/aySicz4O2d0cqZ989
0Ju/CRoSU+fB22cxSxhqJ+LK1W68iv+k1P5pze8JPtvOJIciQVlim8Eys2Wq0clx
bVXYbPiLTlW6KIlgBWwN8/TrMZF7oLeH2usplgvvvUnzwX9CQRoBFQo4cHdq9r9X
zX4TJPGpQbBZUvV2i1ZLwuPEuZZJn6vzZSqq5EuZ3lUbDJUuWIS702GC9d26YkhR
4ZzbvSavc8D+kY2zp+roKcSRLu/rnVJgbo50fHxL/wX+ALqNoViiYaJ40ugh1s4k
kPEfd+t17MT8oTdAy7TqEDoZkREVXLrRcyczmdzeu4hEFEgowpbKOp3NbrwvXH+p
nDL4O6IyJCEGRf7dRN/HDCVQ0f2ccjewZ0vrQuZuE0KlTpMwtiIfVyfebwrsvQpB
vz9ac2cXhXiLrQ9NacA0P95fpHq+QhI+hKk/DivW1Q0FmnXNLikBEfWNQ6xnwhoM
OeonFGmnfbeFQsTCDrKSEj9q4PXqSLh3Vr6R7rrKOJ+ee32hgPwbn7DOXGTNq941
CuW+NI+QeslnSdCDCVMrZy8PvEgka2UGiBnza0JNh2yukxOGC+J71h8jabIrrMi5
doWk3unharw/3cpxox92FOX/BYQ/5+rLZyeVATl0pf358FoHw64822iIA3B5RU+V
ha5JRv/51MIQ/b3ueUSWaDE67hbl3O2O3PZ3nlL4DYPuP5wpuW7CnMWnghSGmNpR
++6gewN2mx0tErZet0RMbAp1FoxuP5DRi4lILGTNm5DrXuQsN93jIGlHPx1OKTQO
mfnZpQt5+Gn0eDBa3vykEhyYoYGinPCBFT3YRfAQCpfi4As0z50BrNfZEv+GW59U
aPhGRFD/QBPIdZ1zqWdJaiMdeTklX5AtOuRPzcBj22CCFdJW+aowYoLK4wfPoqw4
M1Xm9RWws/1ALkQZrL3ygDILwykrC32MaPeP4XPR4ydBKCQ7Z0+WUGerYR3x/YUI
Uvp7nCuDNLeJgsWIuJwqC2lOOkFh8Ubd8XwwdhWDZVaBo5FcBUVphpXFCsVGokvT
HPX6oiT3tzXb2VJMpuBVBPfHcDBXj9LsI9vC6IFaEE3XHyZaBg5dfKESwD0L8ytW
gsnwSQHW04XxvXDU4ZNT9MRcX61QfBLHIT3DyDB3IkX5xdiz8g2megXQwJf61Dzr
WPZsWyFXTMYYC2TYZnvscTYlMkNv4XOLy2LbYK2pUz09KT8KHsRyUQg0AsVhDcXg
j+GmJza5Ge7XyACJ82rTYe6tb9ipnILBMIKv41AO5vYbwZOFM4uIpniTviQGnfwn
N0ay8eNeDdklb10wlHTYdXynWHftX59by75nb/6qija0RTPlva0pgLIZeCIa+uX/
qWLw76JsqWiBrB8HVIp2dk4N8FOK9R3XBnWioeCPNjxnDtwxoIJDMCu7WFKzw/NF
viUXz28Hs1M3RLvHhX4ns/2tjbqdOEex4EgBTMRnH7jBhVfTzXSnxE8mVel1hMxV
MVpyX7YxBWDCJkuhYb2Sg77ReR4f8VGhscsdHAK21tjpODbYgcIZhX4eWvJ7Rmq5
c1HWfdVo7EkeeTUHRfm3HPyT0W8J10XhjRuXTeXZUcDWPvF3Xqp+iW1aJNhT8/Fm
JWk+5hDWNiQd7SRB4Stp1ssByjdcHAmMqipGO9PoZasOAZ82gwGEqJz6sluEEq/e
gy11Pbl1rm3oQyc14ZkHL1u/RLoWP2nqrGD79IKhAjh2sLYDoos+b1kDgrRSTXNQ
7zF6KPDOCsEoDhxCrV9yR2zaK1m4YhHvLtDqtNOY4+zTIgAMjox8MP0G3mV7NvpG
zEwRsychdTZ87SOKdiDCiyQG1sAS9lB/cz7K3lzP+hHrqlK34jlfORlTqjYcO0uq
nBPpPODwgfypRoyopel7WvhvouZXpnXSeWLTCmvjAlJiG12aqyzuFdXHdA6t+cmK
20BczCAw3UBOdYog6mvWw7pXP83eTFVVFiESaBa2hGbWg7ksecsONaV3wo7Uo7M+
S7DI31sD1iXU29+b6pNclZ19clgtqQsOfkaSCqBF99VByeGXyNLHEcIxAemA5nXe
hYqvJPqFUtW8SfSclG2voBdZjKSGudrx4VxVyC2OvzoWOC0ZCsolCpQYF0azWNqe
Ycu+BajpAdcx57gVUHcETyODoq5YxFAjxb5u23PmAn1QRpQW9lCphoZUGBl7cdws
VrJV4HBAnHCKvWZfQaCTIizV79jHpwFPO4gQzElaiDCtczlHR8BRLidcSOlYu3kU
+u7JsDRNwJiY9g24oTIhnEkCpHSCSnA8LgP+FLNjfPboyn9dFiFn++5dsqkAuW2k
d2GoTvqae51rEh4wkddrTa0AB4owyymi1Y3RORFS1jVNCRzR+6kAJCcJdOgbrVr7
AQ/8A2EvVC2vW6CG18twe+X3fyALz3nkfomnC6k7HBkdyRezn+3HOs+wFc9Nae24
22kxxaY0HD3mJP9P+9XYf1qqL5ioW1hJ3pKTYKKggU5ac/Gd4Pvj5VoMlJaYgOAN
HGxsoNPPFD1mJTNx4rZf99j9ZBvQIrWLdmJqSpSYkCVXrtuWCrMXJgBRfg2SW4yT
r4F02+18QSVQAV5148637y0eGoSvGgDfPbqR+L52F96ckaKaVqpOERqvwZ7cbalI
R2jwBDu9QDCjgsW6srSt/zvKLrCosLPuo3zfTjXvMXJyzA7dAX3E5t49at7BBAXd
P2feeFhdfl/s5AhMUqsolehNm9rLlaeM8Oinqpf3sAUadNn1XLZGFN+2k8oCPWIR
QwuAlF+lfvEeGBtkOP1513C3GCuomkql8n9d+6Iivw2ytHUw+6dF7nwefXJbm+Hd
zuXKncfh9+HNuWHmwZBPBOd6BOo9S7V3NMMQrwPLbp1vXcYnwV279moFsVDnNsDi
bMLjzP2mkhbyPPgakfEuwz2GHfzCzlAiMNYDd2REYc5BhGQWFKfArdikjMKG4ssk
b0qxUWwmNbJEEEQyFCUwc/+EWXAgl7X5BeLdbmAyYk8KMCiONLqCjzqGbacrYL8k
EoDHsrJ1ZQCRoIL2/FJZcGPGnZB9tfvZVnJav8IYPNjKtWcFKiiIJ8GlsoMuza2Q
Sz37h2CZLui27+r/W5Y7hw9pSaeWSYQIWXhoBhbyH4uEjK8BiPOQhoe5YweCHyQ7
kmHrZIS9B++b95eKmQlELGsXrAq/BnHAYucqE7kXKk3EzUCi52ka4n4LPoyrRdf8
mEcJkfLukqjvTeXGxyfr1r1TR8qiGaIcFlOrH/NvZHj4mdbiFPKRPUZivV6SY/XH
XgBOiPUDeYVgDmUs6FuXC+ym0YGDiWYdOP7RbFjlAykLF0YrcNZC1EimhiiCd/x/
2w8vAvvEOX8oj+vbP354kN0y+MtqNoxAR9gw14UP2T3auPzflnQhk3ZN5Zfv9eyh
qSTUiqbJpxkS+38bKyVmV0A2h3ZFfGiRkwtLju/mF2BgD6wH36lwd2zw2nac4zQV
zOONOUK6Yrsgv/4PBcTJzscueAtOtpfjeP+rj2EodfSWJCqtGYjpS5EZOCJOH1/S
3SJdRp/KjFRiJiaKyeVI0qIYuWQE0h2jm0OIG4zFR8Z34qdHHQF2vLsitQRUiw3k
1PA8y2rf8GQ0eIXrhW1HH2FuI6iqTT1tjfaaxCcHMX8cUaVfMnmea+PQLPfY3Ne2
J31HAb5cJaVXSkzJsZquJhUdiXEJX+/QYIq8cDlOGVB990cRlNUHSM+UtnX2rHyr
FdVuzTf1KmA/FwfDAlzSYVdaillsDeqQRhdJRCR9KpCviGX8HTZTkXYioCnjrrWA
4PVRWO4ru/3AENo4jS5qiC4DC+2FnrtfYwkhR6Byhll/1n2h+lF60VVBXuru23b1
a3WmkkDou6OhP+8J4MzxEDBU9juatTUtWtbOcdZNh+ohM33R3Wx1oWODJPwPJDCx
eSB8jvxjv1NSjaVaTXUfT4eMY8N0iqWPtuPLyi060InDSCsiXErjvGdr3gDhX5nJ
7nuskyWYPfDg0Hsm0xe/BzKX1DJrhDBoWtrTjAihN1xOpYTtsnCWze6d1LvpZtQO
8CMpvdYZ4zHIjoCe+KQ7+7MpHr8DTvk2hDTGAGbI4VNIsZTyEpwDSSWd4bKE2rm0
BqR69ep9zTr1P+LLx1tLuFxjCYdhHaUD0JYQgJzXp0hveYnnOiWYu9sW9JIwd3C3
/Wm9ZI5SASOfnAWNsmBxK2ASD82vULZN2zJKme71bYdnJm2DJhH1SQft4CXnCUkA
9vb/c4T37yZmT6To736n88is8wZ8V3AKsCKRqtGfyZO1qFs1Hk2DmSh9ZO659h65
YE3jAbbfUoexu7uxrcze/BAe5B5c+bhanAQYtbTYM+0pjZtbgPIoPoo+EZbz9Ppg
XHUuz4qsgcmaXFZWN5zStQKz7WvP2NmmuEmNtjYLI5zv9gyjSo1riO6Fjd8SXTWJ
kfX9fINxMqivfux1fYIs3VWqw48WcGfVZxF9FZfhq6GAD3WrJmfjDn1ZjrRlb7HG
LwGQNm5jTbe8O309ARbUMGg23jkazVnwC+ecKzVS2QkOYUDoHAvOrpMooWik6VN3
cuZIR8CaTMEmI4jBCxnWv9csIJuoCR3l5sPKOc/TiMln+YtZ4oenCzeD+ltqKdNJ
aGzOA2tEYM1IDdFnK0oIWTcvSD11IaWdF+QhNr8qfMD7UlPs+ProBMxLQIE110h9
crlcZPuOTJhMIyOE9vyLe0DFe5A65Uf4IQUfu62V9ITSI/7RPiPGwT24JD51hFBy
HQligkeT1rYz1QSB4ra2vh5ustgMcqKngFh5CbDTRo7877tg6xxlAANGRP8gPMhz
pRnBSMwpqy6UsdYkgTm8YxXLr7tj2ykwKFMLtPU0Hvi+AWsaBwyDQssNOiCaTA12
bxzqBGti5r1hZWyYD/Og4XFBsLl4+yXeHugYD7+uPQKSg/tDvdJeDohi7jjkXvCQ
8xrychRo5//YF+kIFGJLZqbPjsj9iyjABT8XieSwkj9K4vbc/hipHpgW7liz55uy
1gytM4Vq7g9Mb70EfjLD/jQrgm2SwDnGytRPzQygQtXNBMoDeX7z8xyLXl582xHp
5v9ZgxIsq9It7etfEa3m+9sld/vvml1vCtrcQ+RVvtU7A7xFEs9NlSKPnf3mtelR
CNIO4MOpeYF8wxmIez7UCmeXad6VqAkW//JF0CZzmeMFRocgMJDML8B4Gf6XQYDf
v8CtWQzY75x9AlbxHJWUmijcj588eMifwvOJpPiTSyZ4pXMFEIlLzCSY2vcX0geP
x3FaYZdKyvXI+O/Dr11UIWtiTQ8CS//60NO6f8HJdefLC8/Nzzr26DgbJCRJ2fsB
tLhSyE8I679PE1cij2OLVKVz7vZe0nrMzF9dh3+nCP4YPkAWkOcIdW+eooX0Tmap
hlyBMHnZyHn6TFWeI4UQE2I34/LoswSNrzmb+Gl3HrmZnE7fLeEGDZMQmJSIkySb
SQXr0JUcMXIAy3nOCThE8p6cWK6/BLl/D0XRWDDOyLlsWUKNHQmkNkBbh582IjFe
nQ7kG7/kqeGKVbI2SEbHD1h400PyQbkAYvy9sneBy95nhPYI+CPkpDCIU8a8BF5Y
/2iUEtBozkFUTZQVzDOHA3/UMmd5ZJyUt5GitWzOuY0pGbM9TGTTWGANuJuKDCNF
En9XL0A18oLY09TQJwR6p2Vhkrqn4Pa+IpAWdyFh0d1mHeiEAL+Nsi6X+c0F4dWC
TTKibtOfECfpLrX28Jzrvn94lzM6xwwIoaRppdfq8Jev4iqiIAFKtUOPj294pxr/
SJ+R7tqyYkeLqqRzGPb8TIlpKyzGRgYAUYTlfM/x0fi4OjjUKBKtP4+em64FnLCG
W1QD/wMlm8wTPx9M8/OcLQkV5BQR5wWpE/ITrhNoB2Nawd0SyyC3VoIZUGLPxsRP
OH0Rh1kvMcL+QSuf7ehgKDqJbQ+lLWsYpQBFtXAicP7ts3YR+0DykuXCR6Wb4JCN
CoXWt7JCLY3aVKnD9Pw66jaY3dLrnyNugt1H8MZlUkYoq+SHkXku0XW+xrDAQjCt
vunPhMmoXCL1qXmU47RLW0gb6Ozp+C4Ju4VvVq2X54w8OAdzRTfIp+fKU+tO2t//
n9jZoRN5ldDCu+fRhNZfBzP0JR15/zSTh3E7yWca6YOWxU/rj+oJAqzqZ0+8xq9D
EYH2paYuECklDpMg2ZJnc1qLSmAONGz2ghCKQivymyYh/sQcE3mSMrkIvXKa5ix5
1w4L5MlYJPYKjmsmuPV8ezWUkhpHSJaDGxov3cJESX8pIc/cJYrTKNC+d8fTa6ZV
kESp5yaaH2MD8It6/RHhyxVSAEiFzfX5yn1ukx2+F94vxflOIyr8F9KAJSUb8inr
1oBIsGCqm+Qba8d/9QkEGz/j1icRM+hoVjTJjHDnewYOA+pm5z5T0z6xCt8JuTgI
9dh9+BSmamsAN5RHMpnmn+43siSyfrgxiwItEaunA8HBr31FJE4tBz1X/9TVgPhu
J2vonuTuaM4vu1usTe4wntys6tC+hxBxxqOzK424lkR6lxHQnPKQI4XCWpI3CjCR
FxVG7sPphFVka7BI5/TQ0UtISjWpakKt6g1ZKJCc/w15lFsxybg+mbOcC9ZQAQcF
ceghXMlBAjdgcwzBsOK0k5s5nO1zZDhr61GRwYZ28trb2SJo9bh9wVDkpsykELgq
LKa1IJbUuGCTBeXhGqWUwsjL2lc6ZCdiFJyiRosGXAwAQSgCgIZkxQ1m5PIxLMcY
z6ZS08ooERQlbQ5RgZlCe8P+SLMkzyhG2zZJdNL5FH01CLZ86pUE+lYhFYncKa3U
EvPoYWlIQhXKeqc07xjYJECkRKQY7rMQ/YT3dQngnjeda2dbaSIwDtm0F0eo2hvW
MpyR9JOxkufLbEdxq9cB1wemq1rQTFD5PLIu/sHbWFFPYgPkIFw/TuUBnbA/Mwxk
PWN9pWSkTtZzq+/OY9XqWscLmqkdu9ipACpzTJxa+dg0OAx09llczhRq3W8Z7woX
V7kWUylwRDDIo2hYrFaQ4XhVDIlPzEhTkPUeV9sAdJiz7bsK03z6Ws0V+U7MEGeE
zjrH1LZSOoekuYAsmtagGfWdknhn0dYL2MUMvoisR8Kv1h4OGFVAQk3u6gCvJmiX
GQ0D/7T1bzytBqha0GutIwGCebuvC/5vOZZZxyY7RmrvBmkMX3i4MqnMHPcxV1jf
r2fttdMpY2Vl657Kim1GWOl5JMASASe6iq0V8wHOPr0gelsLE8L6J8fEEhUFDM6w
XgE+HYa+yYUX0c6jvkvooVJKTXQ7myrRX0wxsYJ0ZdSIQdWPXiH1WsiQhJKrk63X
qeNXqmdBwqlfAcA72zJ1uWQdam9frZYfof27RTTZl+2u8OcL3/kD6lWGWMvGuuyd
oF6oK4nAy7ITmLQl4Rc7v2jdBkLxKllwXtlHkQUo1Yng1uf77qFt4+1BQ3k6FSFf
aO7HyWbN7m2OAhpeY1IlT7gqX3wmrWKIEJG7FaoE95R3JfwJdVpews4Bba0uZG4d
x1jsAAYLRw/TmJcZdVFFBJq0afMr2aCwR8V2nYA1Ov6L+A703ldE4j9UA5yH5lVK
0iNEzX9vRMHr34+pid78V7xWlS8MbJ2fJOwpNhYC70KPhz4raQLwNYAh2/4kAfut
CrRcCJYUEclQk6orVwoq/01CNxIY94q2R2QERsrl4rGXXT970eag3WISIhjZg3wx
NfwqN4KZK4IbqQ/2FftNEO79PHh5AoauGTaN27t0nH/bAFwmwevcTpS+aX0zbt8+
ff8G0XlhLoX6r+wLiyjjUcS7SOZ4hh60dIqnhCn8mk7s7AQKqPaF9I3kspP8/Wnb
XCbCx1jWIlkgfcMa51XKXThKIWfAQxPs+/wzz5TwQ2gS7Z1lo2ySbD7AKXf9/WUv
NBpSCmOVzXWyTRbuA0cYIaL3/fO08fpeW0vP6GsWig/3MYytpIKUSdxOK6l+0lcG
4kX41MEOt9iohC5LHzuBc+0WDooj3F59DiXeaH4ODg4490wSiThgxADTjKAluBBS
OHO8/Wv+oGqzhGYCukqZKHh2SGekn74axPib0rOyD+lMP+eUg07H4C8MXa+/FTtg
TbggSjIq4EdczXlSNZ7WoHtVUu2RCNQpwPNZsvhhPBrOhxKcT5/JcN4q14O/hdZ1
JUPB3xneoMDZpPI/1E3u2OWwHXycKP1kfgrW43JVuG+Wg3Fl7lxv58pbdxJ8t9cT
giELf6jSGkfkdgz57n1Ejr6zK8UxoiBVJlffgGvRRhynYrGt8/HKBGUaHOvT9eGx
AI2lAP1pvLdWFDsmb8wRivcmqvVFcZ/G57Pr+Bp2hYxwBhCrW8asudDka8sKIXbd
yXhKgiseg1BxQbMxeL0LWuWszwBo6FkfPkojQqjVjeTvAaVJ/jx5ywE9CdEtVOho
NX9D92mj4V3dBZGmgqFVAvG9Yer6dRKb5k5sTNywscSAvCMc3Lv4Hbmpd7oNAlTK
CST5NyorE/4SkeVQupepcizuZx0VpXIRoSJF7RRHXbxQtw47TdpIETZbXBEMln+N
oIJgmOrgy/iMknFmypjj/PmGPoyeIHOprrg16NxT6hnQcb1Fa5ScFzKJD2DUveWi
3BKnTrNqmx7EJdKWn548IoDAfCeJvQRR9F31EmsF4x3S9AjA+BvI6Wc0DEgCW7Po
igADcn8f2+GLjFa5fWBGM3xGKOa10GXig7MLOx1hpvUwreu3lH9NWwKSfUT7A9Nf
48SWT3zdLqAMSuAJD4ocp9nKBlhzau+jsJIEIfRj4UugrNziZqS1nrPQofyi6u8q
U9/SL6UndRBHRm4os8G1Ru5TKVq8WsgyAbOIoGbBGnx+0/47cadplNhLFqmI7h0p
2HJBUpRMrdKft0nCADlREIpYVxmPdKUNCNUux7Gb8IffgC3aj36y7ffrKLBFwAT8
+pH9u+DjHBdFsU5CR2eOYsMmIdnJGt8wMQ1kpr326znMGQyXIH7L3HC3bj7u5cSp
1gTv9Dhp55zVavoTDnWdgrUfWyYtPCf0Xa1j0TI5QXT+Ne3e3cDYZA9AZ+pqjRcX
lVtn8y6qnqV2AWc+cfL9uJsdmeb771OScN8fBGfLX9aEWrmSqLd6JkxOIIvPitg4
JW7FbVQ/P5opHY2+YIHxwLzXWSIz2tS88Ex9wGRUME9i2ttIy5A0PDooa4RSjd5P
8cBVA6VT852gu2sRMvvEp45JXcNj2H+45Mb9xuLU3L7OhQR5uNIGS42+Yk6R9cfY
5N9O70kcbiiVaebIAd7BfO3GZ0RaWlZ1Aj9V820djmQc1TcikT4i83Hz5ZoFX903
aXYgXZHoClqrWJI5MGuim7oQzmFyfltNYDpQnvoZWQUoKirZVriJFBHmNT8EPCQ5
JqUSZ+eYs+szkGKfoY1boODTS3lyhsop5f/bPf1W/13+5PYzUx7dulnAGz7MxlAD
0HgwBRCRV1xVkiKwOn240vs20VuoREOIyEa+E65d3SMqMZxQKdj+I4WuOdCdBWV8
kq9tIqXXmXEWYkZpW3qYQwhcLld/dz1U/AqvAt5fRWij4GyBMHU+wJXRmAtO3YoA
DCwn8QaIDjLwdVsev8q2pANu+jbGlJuOnDbNKcXOad3FVpsB6mikFvDSofkXxHj+
M506OsOkrzyy/epFfwcz/SJCNN56yzWoWrmuRa90np6rJd9uPPvrHWkAFyr8p6Wq
tMgkszfakkqBKi+KwANg9bjqw2F6jJtMXLf6nsQvVGI1PPgpr22j5XYNd4i52G6m
k/Bb5rzgHn6z079ncJTQrbCOgtNfw3wZI3oQu3oWziZk5JPoYsxG/1pyx4pMSbMl
UtiTggtkVHefpiolxZvt/jQ4Z+eV5hsUmRCNoSxxxPJnWatuJ/aAJe9J1SQe6T9U
ynTerWUdlmhfng34MehENVUExk+Jo2p2E6sZZWpKgA/IYdxZjDKrKVu3P0KQhwcy
TdZd3eltXi0nPKy93/kDnKf/fxbz0jOIWwsJLGk0mA+/5LSwYW+Q+mt4G/xVicQI
MOOE6n7ue4WoxWiBdLxV4Chr9bS+freQtvBWOS8oSpuZ1WCr5CXwZJq6LyWwisv9
b864cyYwxWuaz8rjMhBux2iGrM6J7x0TEDHPmP/BvS1JW44+n6Z66T4ML8Yk9t3m
+2L0rTXyj7B9wSie284whAPYdNffTvTngLtSq5Qnq7DAQqcQnXMJojt604EV6EAb
PGjXbbXez3Tt0kkEJVyDukLct6hSc6H81MJDk9FJMNvRTItynEPKYR/aY2SZR6Qh
Cwu16cJqgRongaU4f+Nrv7hc43frmwiVWVy4mioUeDeHA5S3I6B9b6412qynUSL+
IS033bGe0ApBPatRDrhJYMJkjk4LH8hP4/gq6BFTmnLfurLOUnR84FHYn/dFyWVW
kNmHkIV1VCU9U7oiksQnrlatgOL76l+pdLnsgcLR3gRrFI9Rtqn23keZ48qpp2X2
Ms0cQ/ORoDzvISzof0u1ZdBJFIG+Mzr0TIO/Z6D2dH3HIvQUZ7fdq2m7Y1pXKCjC
ktsAqhZK5TZxBkLJVDmYSl1h/dA0d+4XCmqlQvAemciouPK5kY3uqkNdNF8QwXWw
gij9PgHT3wqvq75YbxLgdgfLUEkekTA0wC8177pPAKh39xWFpty1j9gFoxK6Ywaa
EabYgoMn4GIdJVT6ILo+SQtLmM7s48Zx3J1/RVmSHM0kY6m76lCcsv/CdWvnQAOz
C6fKv0sT+nmAVXfWWSQlIcII6+y2gOMzt2kLMSpj/UJntyZ5MD9xqX1zImPGG1y7
6UDbib1NcE+xlH9vvOg0bwn3nJYgPANqztng6t4VA1gxkt9hN3boZO0BPy9XodUb
EHpZ5hM73AxXDfe9g/KEfTcsZzHY6RbkMQ3RJjPJ6IzGs7z5rWpBXinH0afW1kpV
sJsiGnsbU74bSadVJVxY6l8if4CGD5rZC3UeWZYj2VUzk1eZkYroO2Ph1S81Qg4b
VOQCTJ6CvS/5p+eOwKR9J8KQar2cJwRaUFmlMciH5VvUHGD/gn7C5xpBrT5+JZQA
Wu8uyQthrpm4UsDfviJ6WWzUPxjVxxQKoA2vHKodorig6Ja+Jd6CnedcTqRSoOHT
fuYoHM7pBt5xcePcgaEY0qBsf1jrgASYe4UhFtrC4FiJgaV1+CivlY+MdcV8O996
+Xo9Vs74vKVcCKwm2aDy5ZloK2rpMXwiREdRftJrEnDZg5i9n7d/DWQ0qqpdg5oK
128pYa4OpqbtLKDmcq4bVvf9EaIm1E3wbnYkr+mn7Z2SPmwom9rtBMbpAyxi+0tK
OdJzXuy5OeX6R2FweLVpZmbMG6SCGVNsAXaugfQmOJBYJsyE+FPAUYt6Hdc5Ffyl
iXWXicxjywfOq151tK+UAWzrBfVoSbrOMgg3Jg/vky3jZptDmWjzRQht5TNFl52g
4U5pqR7yZvhc+MwQmDdokznadcY9NggnvSQtOFctSJqjkgG5FFO4eTnkqDAYIri5
h4Fk3g3USIVAFp87Vzbg1J3yL3hmIOJ/eJf0ZcJqD7SC89oUcPnaZassbvqBRhAW
oFSMBzmiiTyvOYbtpy5CnQPesv/TrUtSOkYcYkI1mdjoUp7ZMlFr6+nUvJ0f71us
VWk3uYL4chAtS62Yh+lmoghB9NAoAkDVcScad6+OnAz5vJ7EY6YA3JHNNnhCnR5A
qiK5C9C2gr2HYUgTFQfLkQLYck+s5rPOnBKqUYnEcLEm3Z4Y07SLUkbFfI+Kk39n
J31byCmqFBufZERVdxZYSBNv+U09Q0FH7cvgvlp6JgGWiyb8RVcxfz9CXHbtUBuw
M4/1gO3nfJoFhNLVN6jGa7FcPKkvpg6Vki81TGwDrV/64QATu+knrX/mFihKsp0Z
oBFtsAfofQPJ8hMYEEUi8xSxVGCLiZD9eUA3DmLsDVcaTJv3adFeIsGGmr/ka9bC
cCAUYerzCa5/5tL4yTa7HVbVNHEyP4b03rFCx19KXzN9z04qLRMgJCtrRwaE+SVH
iWpZgYNEqs2h7Wz2Bo7cMImopS+2EKkCgdtfhHJ6/YVS5/kVCuWg48X/q5v8WHPj
kVz8B2GvhWg5XCOGp1tm+TmbowdCDV409zF8uX/4b2nkIRM+yMSXY/v+34QT2Zus
90539X1rtN30z0iOzYbpi2epXOj9xOjWDuRxNIgcEfPF+hFy5XRnVPkSLYNUHydR
GIEZwBveSIiugxuGz7B9VjwkRYwcfdYtVICsvwi0XDvl9B6Lxi0d02hrS1JXBuIs
NRY2Rl9bfYSXSKwl2rGfaGxQu8AW9fEX9SJtdpch+3GlzsaO73T3PeTXRRaZwpYw
MKbv955PeOrWK5sPQ6HtKcgxrEPJPtPJmIsQBHNlvJj2b/9W3K/w6mmIAoqLBueS
yiM7QtKc20E8KmJ3+HwKd8fAM5GEROa8N+wV26U4ar6ZTMK4NfHKLgZsT6PBWCno
M72HnYMTwnm2vkvqu4SHNhojdW5LxPLoGZf5KWuPr4PzLn4D7g2zyfUrlc8Oj8EQ
xqDY4VBTL32eL1Cl5XrCx36kqw9mpow8WMw676jNvxRTxjYQr2yldYmUbnqRkMul
a8VvvGriHwH52ycO0GvaljmRcU0HCLFJPzeMzVRTC58/kuLSM6oatD9YpH4FdiCj
Q/GkJa2Z2J0fDAbsiQP9IXdcrmb2/IdbBxI4VAr2XDCnmSMMkDxgpz+pwcGNkP61
Qkyrd0WwXQPoXEsSsyxbD8vohHCr4kj2Xsvq9s3XgLASdZ2LFb/GkR393AG18JK8
9jCSjmllJWzY9HGF4BlWKd5AmZGI2+WalwRxpmRaVehLZy0mr0t9oTMvBn4aF3gt
E27EgSLh0vsR4jcznDrFdrQnm2isnpmvj7pfka0O6+aDiT6Cmmpw4UmYEmWE4JPq
tdDhP1Rt6nbTyVwKRn9HgJt3BKEuySUsfATiOjpGmdPBwNTb/UpKTNWBXP3uCJVk
95RwoKi0Zs2FQWoNCChkxSLfNPUuJ7QyvckO7/uNOKWF8hpQA8hZrHt+CmKxCkgC
qlI0uEHxguOmkz8v4LdT1QQUgVb1Gplt/tI6pt2hwqnnhllz4f25zKMqmcuDvPDL
iaTqZHUp6LyerMkOBgVeiRj5o7IOKona1PODV3h9dvlLkgffBhXEq5EJRlAwpeDX
B5NXN1Qz/vy+gsOkz9MykfrKHwxjQOy4DAVwNCLT9G86r4blLNsADZh4Y6FTlgUR
yyIKyWamWmM2SfXmJvE/351JQClz83aWiMN48ETAnzVJkBwuCG2E3Dr7HJJv+yHD
ZgToEDC4oNCBMGGm2T8fQVAxlnQzxIIcSqBlUCHW8DlNdhyU1RDHw7IMNHUbeG0h
FxhFf3xnSuy7vW3TZ3tVNXr3rPtJldQNR1WeJKr16AbhtRNS9nt7ZCKV9xtwdS/C
wCjPGHmjEQGZdb4pqIuiBl95yQvXmGuVs95/TPuB7HmFGLom6lOd9CGkPoCyFslT
gyvyktBpfwgJEVa0bbewJIyhCm8PpEvIKn233F+v6IAo2s5fDMDgxgqzG9I35glH
Oa/4jMyDX8FEzpKaJlZ2FwuwwxOK9bqSj5Xa7/IkP6rmv4+0LQEqFa0zYYm5azm8
V1c1PmOX6G43ovkesIIjMfmPuONEMB+IydZ7ABzPG8nZRANIdL7hq3KiihsXo/RP
VcycB8hLjzOJ+FoCIJn1wRE8F1WcFm+2ZjFva7KCwYRGIah3corjhvHxY27o5KAN
ddiYoFUmnmo/BUcFbcmwuC/4CZqbzF3nJLqQn7dumL4NobSaRQf4+PF0KTJGG1Ba
wnw6v+XBAVs2HYJRIMbTrPtC40azLmk2Iaey+b3YRlmJTNRqMNew0qYhRWQvPJYc
n3JbDyaQOnGB4VsItjFvsooUvarEjXQRQ0Pe59KttFZFt+/3rLyU8l24DseycvXA
lSwzGHnH+Xod82qTnNzh0oSpOBvxlR7wyxEoITQYKYQq1T0iwjKbTps4dw01MyvD
EUjJvLO7FayHJGGCLFww5HfAFKjhKo2JjaNBvvn46ocKPjm16AXxTK/GcS4LKDe2
pP31lQeGoV79Xn1+Z6dmomRjHVJ6GRlpCsHr3FeHBip6pn2L/Ce4XKRTQBMsnxNz
AOeK5ZfKoIEpJeigusYdRZ82JQCiOQtgpMOusZy9sgQ/oaQdW0xs9rF+t1S6PefX
uRozUew/qPISkrABimWQsN+ImS/USWEt3pxGShd5f79dfWTxlSUpQiwFovOHZuTW
vC2Q8My6glTEfoLZG8F2YDmgKC7sahCSexgz0r4DyJFqSG+fkzsytLxbd04b69Im
//s67uCEhXtzXu2DWLU7xAEqc8etiWCl2ZtEz+4vm/XIuhe6uejMGwO+3bpei55q
878HauamUTq3uVO3qiJbgAHeky1X1RXrn4FFJAA40D5hblGC9KmS/9iMNDx8hsl3
XKaZWwWHzXViukyoWE1u84zgaIggpqaTucr/lcLqaRTVJzU/Z9yhOnvDR7wdJrLG
OEJERGj4FvJh99opZY57Sgzk4R6QzQ+KgaXA+kJ4/d2WwQAB4siulZSJvyf8U3Cc
A+XJ3DMWR7cfqDjLPHEiX9iR8yLrKDsQsaw05UPW6upARvFhvuumhBV7zKI0sSUi
4XnCF5qtWdjhW4vXK/fX9Lsoncn/RLhJR7R9Y9vOTkKA4IrYS5lRN6iEobPJPQ4G
CUDnM446n1PyICsp4u7TVcLPUEqxAa0yT0xViirupboCGQO3gwO803rmABPJ03Nh
+cOQvls0/rppDuLxHYZPnpAhZBYzifhY8znQ01UO+UVKOlDiWqSArt8HtDMzvLUB
q7BXR1XrjcVdAHczG5WOnD2gnP2LTB0ctPVqJaiWkyevc0Dwmw2u9Wl6UMeExhhg
zc5tumUN5QxKcUwwdOaZwJB9UxJ8thP5chn8YgcOCNCYcgE+T4uo4qUaPujabZI5
PANEGKF5d1MZivFy88nHTztGl/JXVnYkEwBpzET/7RSu0IfEm6Jfevnb4gBFxHuE
ig4wIXpErId9OGCgvGg+RxjAm2NrQC7E71NsmmzZg2PBBxCYYkktsAufB2Akb9Ze
k+dQmtMi6vLJwKkQ+xAVWQzeGD5Yr/JmWUe4QgcAO7Xca7S/P7ZQLF/8BSiq3WC9
fWunzI8eaLm9K6CyZrbvblIJpkKhQNuZaBQPIJbWDWYSrssfb40EfiYPHl5bRi4q
T1uvH3vwqEUxjfCt9rZvBxDccqEOicwT8kAb9692/N88n4ral+IVYvZQy/ZIoNVv
cul6HmzrfOaxchUtEROFbyqV4B577Dcs6Y1uXrnyLCg/yqCskH2m+JptbqOx7wD+
QLzZgSN65X2sEBV2u80YXfWxNvVkpnmVuujsdVY3pvZxK6qluHxy2k2GDTQ5uQAb
WvCfokpisWNl2a4NsIsXz+6ET6zeXz3pMcxEBPM7NTf53RTlk80ySMNHTfsN/9nj
aJtqo+Qrdz1/718jt7hqyb6xTglwwK9RRXiA7ZLB7qs12mP19VdFBSBcnQGyJYw9
EC0FYlfEcOjUJE0bC2p2Tb42Gt1jlW0kMqKRXy5+gOeR7NuX1b0ExCGtkidd+n8Q
jw7joveEmYGdTh4buf/nP313kwll0XkHAhm1uZ7HCV5fzBeDUWSl+PPNuF/4bjh5
QdYjPf4Q3mT3d2z2yUHg/MqRGz1gn8bcktegeCU8OqQCJrAm2AqbxWQH068Gp6RR
a80CCKIMxYzpYgb0bLKOzXXAjiMYkvzv1TL+IXY2rzASos1uXS/WzAHtzb6E3hkI
t32BlrmL/LntBdP0YpPx56+qJPAUp05Wbias0sYRNTXrUbO87AdC0qTPOT6L6GjF
paBFFyqoplkHIAZtuwy6knoafw7sGxbUR1DalYBBz6UoDwOpDcDuGiZtiKI0IYW1
dISNgfTo1n2iE/ubimymKJCmaMsrdmgj3/1JCdVtgw4CZ9/TQB5z97WZSq8xWOLG
ZK4q3RLsPb+2ffaTClKSzTl1HAp/jN/plTkI/8HFSD2DRUaCmBGPxwNgWG/vbDIk
9hhUd4mCVGGh4ReFyNIh937q6vmxccu+nZcO6rvjYzuHA8KWlg2bpAFCWJ8UtULN
HFzAAz3VBVdmcDHtLuenoDb6u6p8C1kuOgEJthPIp5XRLdAyeMUmR7/V1c1BJmil
sBGOM1PCFOkWFyQv2hfKBM/PrBH5X8ikIBpHZtzYJBXWwYy+Fa5G/o4ajUZIy/1D
1Dqmzt8nvdBjR3brsgDgTYe8fd7l1vwblX4ESZQMmct+L2ryM1FpRfje63Pizh1i
x7XMKqO15cXRmtfZv56hVCV7NX8qYWypGe/ZQI+c5cuREw7d7wGAtMvxZnAAvBlr
95Cq9hgQvDcexqlQcEcFWTr+uUs3mGiZUW/+E8H/+dqveDytSxWesLwMm/hpAxq+
7q5C8SP0LUQRv9y8NI56Qvm0ZLN1NrhZWfszZvQyJWQ8B15UYAUfmA1O6+QoYGGy
AyWJdl6CkZdRXtLUdoGDeWjZSv/1fP02OrBfJSR3/EZVEbGZwlE1i55VwmQvmaRO
I3X0sidBzFEJAUkaraMozEJGOfUOKbXeet3SoYnuZtYfOdFN+geJ51jNFtEfcHcw
Ri7JiGhvsQeiGC/nwBYsEKGSBxlgz8wlVIimWXDTFPWs1lJyIg3rxpOyTkld9XPs
pjuybqToRroQj8W/FKOwIKkGgMiCKIg436CdJXDvWdDSuXb8JYZXB+sMrGZVL9U9
LUS3rQ8U7M2jcjqfmH7Kav9q1uaKJ98H/ojGqcTViOl+JfrdN397CR+K1ovhj6v+
06u5x62gotVJFW+z37BnV6FQgGP3MyacGEvSFniT1GdhgQnCdsmL3OO014KXcuyt
x7+owoJxBSWHSutkmPf3JrUn73OubW0dAdD0/aclzpvHWn6AHaUV6j/mE6lNLTe/
z7wgp9kgnDnX69O2PxKmCfFgoiuWdd+bDLnvcObQYDg2el6nCqvTolcjtKf6+lGC
z/RY7zNIoLnkMNN428jXc3HbZIOe+gwEUKyKG4ueKxPqFLN4xC6szsgbF82oWRJj
J3Qs+K/TqFLP8snEbIIf6XDfI3K4PI8RxXvGgxf65o8pCADRogVyRKDG+cjhuk0U
6p52jOWg0c5/6ugWjzzSyk7Ut3jTJvuHjNUBJLxe+ovsHNYHfzsVARgbkRKHzrm8
UjK4BsGbn7N+jH1+aQxpxTOvNcHUVkzzpikaStSGkfIDFkTAIB6M4mSDqJTPOtFm
xrozR3/9a00TbWUEfQfWdDZEcO88aeQ/n1nO/0DgjG8NFzKwXdDbJUZyRkp0vDhO
0E7Yey9AnvLiZnGZYpMfxBSp0z9a4Uf7gA15XvZTxTmeU5buoC6WXSgL2xafoiDp
k/FiaBHSnLmsmA+qKLupSLhHI5iofEIUGh8ITF7wcDANUdrBMBsgKxD2lbqxxw+K
hkm2lXdNjNLiDX+SwqpwxXDtknmpZxMHMaDZIH3vRz7RVo+7fmodVL1JpoFu7dLz
VsMDefuTlgSBjIcjVyOuUntpBxJIZwJpF3dGqlGwYUK+CYJ+LJnjxiAvSZ/ew0Oj
PbZl0kI4Wy+25HneCZ1CxdAVe17Ey5jjAS6X6GgzpqgCDK6R/G8wQs65JXRSYTKG
w3R10pT/HcpSF2DYoAkHhGasyHUnmB54na6GCGLTGLq+EabQRznGGO90mhuFWHyr
vyjj+UpWH2FupDwei+W2dX+fTRg6Ki1XVtMwQFbZrQVmMQAUNVmdx8XwgFj6mSRU
uPSdnAGW8K4f06zXfmEX11OmK0gG/1jg0Uz1GZpSB7OuF1JjneGhi5Y+qweQCg9r
ufr95RTUpOWSGBs3xd1l0kFsXSYSVE7lGOqOrWser6oBmC3F+fTgB4nVE3RRBY6A
5889gvI5oI1rfwwsvROgShyLuaGtoRuKj9soQfeAIXY/uD8cIj+7ebzLsmB4Lgxc
RRdaJtRhD7WH7eRA8SZjj789mX4pKyT8KFOZW+FmD+jnDCSZG+/kMhVAcL9z/oi8
DCMceEHuvgn2Xypy0N5TUqFo+l3akII9LTr0HByTXDIjdpD8T7UdRDWg+5Ib2ZjU
YLSTvts4xUrTbkaFRsJ931Ovzz5TqxqM2aUCDY4BQgw6KB/qpd+785iYIUrrNAxG
shl20vPsU2V/JtXtjtP8jzQE/6+LIWuJhYeuV2Rol/3ahOS64vda5668JYPl4qPX
OMdPrXzbHLDeNtj6jvTpP9rtydyDXle1wjtfjnlJzk0x7rDj9LSDWiHUwJ90IwYd
PHNiM0ha/eGYytZGmhPs6zGcRPZfaaGhZ/QSzKMd3zrDg7HBFPfkAGfNYPZWy4lt
x9vxodbWax02V0qIp+SxmdgtzyT6DvdD7fGU+QRNvyMJUpI5WrtsW18FbR6E1nky
lYv4iYIHNx+0I4DljxcUk++HVfSnQLQWxJ2RPlnDJ8+Ko9ATJ5a+5xx53qSLIjRG
g23kZ2BgIuxXL2Xk2L0VOF2KD+QZHg9iAJflup76PU78sQEjO3XpMuguRFhYW7wk
4K+sVgglLyL+zTwkoFtpM31aFwKTT5GPt9yUdF/7NjDlFkv9afu3yRS7uD/WMAUB
Q2sHxQlDIZsb60/8FB8mE/AjavkX0nTUE0Xj/ss7A2GIwSo1m1R7wzLcnJBLQ4ar
4oENUbNSap6JXPvVE3Zqlidmx4k2UH3Wd/pm07w7q/Bn/pzxxd6WJYAD/RKETSLY
UpSYn+rEJzIF3rHo49JFeIGMExSDMlzpa0luAo5FM0qSHyyLG9yQjDQaSzit/zpS
BrL/ZgYEPPFM+XLQ3QPrFz5BPXM5y8YhOZEQxd4upniglQ+57QMa95Ud0kq0QWhg
x2Y812UprjX+itSpVfezZhHU6ffTmEcmUVfM8AhVv6DqYnnXUjmQBkMUNQFy7ycP
XBqjksVrbuacyX0+/2IkRw4a2i1P7IU5geMq4h3bX2yXWJmtp11yCyxy2rGhXnWA
opK5SbmRMHgU/jyag7k+08OVpIfvIAXeXaxl0Zi56PBN0evWpYjq67M1vrmEhERb
+8pYjydySTEu4CAckLmCIgfT1GVhvr2BstU3N0Kh2VzThj7CjnTVpOzynHMNd9VG
5WRAC2mjYhmwT4KujdUrfiDvzS4njAE+Fre26qCLnSuwo0J7/n2EsTHEge6H74qt
+kBlsgbC0HyTB4/J3cU77ji4b7eVNDc44krOYk2mDBn1JUVnKr1IKUcbKqIUg8XE
1tqbqHT9R75+HCbiqe/evibKVixXYMfd/VrjFm3d3ZwNaEcY32Z2fllLo8r/XuPb
RA4VAoJB1Tcl7yCDXTUjYTB8XLXxS0GAoQ87flr7trqfhG/uJS3oXX1b+ZOlIrrt
Dt9u7mb0DCUcoCLFxJhUebVtnwa6UKyEXXk5ILcwZSBNNQwXovaCtg3TLk8yWnMD
JPpBsc8plAzxmWG2Ja+AjF9wBBK5V1SgqRs9xKyGo7ZurqPYwMkBzQTWtJ3l2ttb
Oc3UsX5HciCmEug9e9cuB5WK3YqfGAr3qT6A9Vt3hyjxvDP2ic0Qnec20tqX0aN8
46130jDQcc6BBAtrEti1ROz96uG8YfkQJBPYj9BMGh+tV1Jjh6Ak5nTG37d8I2SM
YW8nZDOpLSqMjISqOBuUpKMBf9mNfWtTQqd62hwnUnjVxhJdTJtDZoaE4HBdw4pa
5rDMV6859A0kS/vkUmhEyDtsrvnAkwrxoDfsiG0QryFkAdKD3L1kHMm3le2r/Qw0
8b1GDpkFpnb4bHhYurspAHpTbIL4JuydckM5lWD2jCN/kZukpb2t87T6oMIKqadg
KW7pRzm3Fzjsrfjnfu5WGv1o4/2OyL0OVr+7S/CzEY1aRLKVJWKlXX0hPiPsj69j
ZmrJ55Mh9qKCzIVKv3s+ZjoGyaKJcI22km48IKdxt57vKmULXFSnGyP7Rf5hRdh0
e1eNft2ufb+Fbo3lc7lp4gEIgk8+Ei2w9h0ZDr9/yuPj3YGWFI6mtW4KjBgJlIZc
FWCYQjlj4wr5eZ1MnYgd5tORag3omCxoOfIop44PURjzSXgyGlVAYzZMZ8tdNXlC
VgbMtA2IiQvEK3J5UQyz9USJHz0+0nBz95uO3079qTGr2+lZ5uR5dOjFjm+X4Hlm
y9zhR3C7mVNKMzOIVhXq1vyWPZWfVCTWeqgAKx6w/R2CxbQ6QcfZVOPOWP5mIci0
8/TSXD1EcCzgnEr2MotMHiZSGMAefvPb2noZep4kv5caPD7b7nkOsonaxSEl3Jb+
91XGdwfBpHKB8H2NsIBSloUrP5NmQdY8JSNxKrSB93S1p2K897m+6bGk/kEHx26y
aSD6JfgzJ/hT/lexOHgUwdaZIwvPZGU/g37L77XvE26qxTWcJHb9dKki3H1iGt1y
xcTG2IO5wHAdfigjrOtPCdGv9+UGKlDDE1yKvlyflEePL08tisDIdSdBjBSJMkUT
cjLnHtHLaAAyJWOgDkmEvBNj45yLHmEv+c5G5qfMyRI04Zc75On4xHPI6iWgtwBa
8Brl7sbgfrWR3aJzgS5RDS/SovPppR3fjOCiupP1/XRqbdai7zdkl03DXusTqFqN
4q2kLoLPVBR+pSb5mfBTj0T8gIspI+sNnRCAdOD45HS1aJHJFKUC8UsUiwL+Mzmu
4ZYY6CkPVLI19msc5ZISHygZXf9xPgPabKo35RBvzBmPiCpNsYav/47/YuYnckZQ
ow5hMGRNfDRcxXwTPoBMoYjVX0Gg9XMkzXMgmgL80X0wVror50UehuQgw4UAqXSC
mUoaFwwtnJA+DWvu3Vj0Sc5jgi7xG61Po1tLtsD+qQDYJJpvuIJvtm56xQvmWmb7
6o07TbAPD/3eH6vrT8vH56UtGGmzhbtf4Gs1l3gEdrEVyGrI05zCZG4EPD6wi7tc
t6kQZszt4SMy7Y7kKXK9EkJy1Znjo8zBAybymEiSSd2XLqdUUUS3ye4J/2VuYmz8
zXnLD7YFep7NAsm0uKzAwFArj9JH4jM4+7liZphIJPfsnU7WezGfyUFXeolHGPSh
vKVkjeKD9TZ4Kz7vkM8A9O7WRhGk0npFr+nEdoHQqLPfgvJgKZ65NbeZ52TEB3Yf
dBuCopzD0Carx8NFnqpxmXVm102UI6U9kSnNLLWjNNXsQOFDRpvprmIG6y7ZE5tt
9ITgz6LyX23HYgN4VCnYIvZUVukZY9eWYiVIMn+5LabgPvFyVLlQyC0Y6J9R6Ism
U/he4hmk7D6pqObGWZJmr2z+EYD/I5dytZXcLSsn73vrkhI+aN1ZIWJLym404v2y
KZ6Ba0Pz8PnBhd3ckN0bLHvwUl7wdopRUM1MPEYDshptY9blJyUyDsI3fPhOVDR1
Vd1vAutEpSCTucOAGNXldvwmZxSdgThWelnW6U5zsdWd9VTvIxh9KKo7gAKp4CXd
HbXjPeXQV+DP2/WgP8qRngBup7KwEhD0g0Vu/gv1meL5vn+EMw0RLWM8l2nkrFaJ
TOl+FR9gBxxc80raCU29cje3AgkaCQRlHHBQALbbCTNmjgXahFjQAqQ4CyVFNztp
TixfU48mXgd0a3jxeGbp1fd80cUADdjDlAmiaSbflA6Tf4kCWrlTdupXYtoUX+Lg
9NcXqMXCRziek4J8fdmxTbbkrnr0n4b78wUBqly+kI/D7eb1QJW5uAPstOGT/0CE
W5vkQJrWvamYzsbu93wk8KZmtnlYQ1DG55+49H8Ez3Qtpz76sie5y9mNFTuVg2xi
fE4zYrp6cSQyeXiolVQzEB/HJwZ9ogkdWBt/YkzBHjuiQy094ueO8C/uSMT/+lR9
c8gzWpikvGWlXNXh5tFj80iifCWmN9y1DIz5G0rjcWN63D2b84uyzwzcwS7W4KqH
wwwQje3I5Q2dWUfYnZWQxUjTWywOVCxrzHtBNvqEdeYj4vLBY795WESmTo9396Zk
1q/ON+MuAXGmYd7M2T6e+QPlJI1TtYdN/Etg/SgUQjwtGvtUqjpzeqKdzrTHF0Hr
+THC1xtPpSmle7UeB3xB6syzB6lNt5mitcci9hA2I741JjWyTc7FxdogjaaPeEoV
Ujt70ttNd266FQBEBWMQAoNhdNLLpH/YbY3XqJqL7OgRgWF4NZdPRmn7yPr1R1d6
qMLXpotqNnwQU+TSId19yQn8HgtJuNeKwFzQAbDyKAW5AphrjQjndyFfNwsTbSrY
97qO5lK1AV3hRWPyjWqwfG02T4PKOOzL5n+RpRdB+8ptZcThpacrwRKKZck1nrcP
XThWLIzbQD3AqqwGce36iHaQXwX9vI6FdX1TO3NkcxKb2YtYS5VbBe3NOkD9NHlg
yx50/OgiTgnPFNBSx+uihk6Vo7fwuCpVXruhX+9dNlWk01doMWI1M1usgD6bjpkA
2q0Bg3+YV5PanftcifF9wxKqLPr3XZHhzhAVguUNfDatYhNbTTi2/nIlcTicR7dz
SNNn40gIQkbn9fDnz8fMQAVZsKFbVlBWUgmJsVOFV2fIM2uMHVkDPB/VY7Jaz69x
yzmizkWINzOvaI2LIMqLyhiL5dsJxe4XdCG+dI6+d55uY6h++KvEzH580kgYF91y
Sj5fQdb+OpwsB0i632INRGnaBeuVZvA+rSmYzs5RLyPBnDU+qioSE8zkCgOWItsg
PT1A5I7rVI2Bs+HbtMASyv8T/MSn5bTa8WFJ4tkE+1mh0ZkN9zsiS+JZWR2Ue0g4
de6DUBHbfrCTo7kgytPG/a6zUsQDOabscu/QW1WGDvycVW2zYamwwr83DE456cjG
LpP3fY3MIOloE7wuWSiZL9b0wuxn30Dptx35ZsR2GS7n6q/bEmrddmiNJO5EZL1C
6HXKpjCmXnRo96zLfMzZJmypoYTAUVvhtROPlmq8Z8nsdGujDfrix9JscjaaPQaT
GLPD78UbfCABMbST8YDKpx5kxH12B4fWUKoGlQDAhS3FCeRJACzMCSsAV1jRuBxN
Gq5OM7TxyFb4TQoU2ivdcX2l/Exft7P5BFKZits0liLWEYKhG27UHX4Frvjy7olj
9ubLKXuyTaIjZZkLIWnhZXm5w/46lezym46dIYLxf5zb3rC8VluPqmTnD/tehP1f
HivTMknRenWWAF3Xhdy8buS4llrf9d+QmwjehO3ysbr+4aGJFVRDn6gP6zOXP1Qq
OMaP8SsxyYE94Je8ccU2chMmNwac3XYYM5ZPrOIrooCrSz9Zaq2JsdGKWqOFVOX+
NkAxymSqzpsz7zbGAcmfFfLjobDGzKZCB7ZvuA4zcU3DsqEVtAL1OH7A0YjRmqWI
kSYgmLKH3pbIM8p4lCbEXVXi9h5FID4RPnR3oSmZGBOYIvNMjLe+3ugUIGPoBL+G
E+6srcUPEjnWXgRi/Y9J4mmUvlM4CGQf1ylF8iSwTPSFSTykCWHkC0MDrRnKvPCe
XBlHJdvF4DU+ptk+rMdDxx0T4Y3qENw5y7/LN4vWN008iI6GBTJsUCYTnQVZsbCo
KDjNekfIu/pdhfxLx+oKUjL3FHCGOMlEjZUpYX7wNQUQ3HDytNnvSJjOIBYqg3LN
NdHk04WwIr6j04pyjROG5+c+JKlZ5bD9QkEgHl/CIx9nicJEteLEXGxYx2YnOvz2
d7HfECBLb34FuVfV1sWXGTr25363Es0S/dMKTiVzMnoRSMuk4gwlSXOwOqUxEu/T
KMpxTeWOipUrlHtEh69tbLyxKj0bMjoWlBhsdYa/rKrXEmaqHEoANP68J16YG+Sq
DNnUul+nxgNafp2YZLTtCJ03hWGZK3npG4ZWvoFe3imGI9ES2TXEUu2eNbAa1pID
zRk/VZpdOxELVQ+OtHqZZXe5WMpkTceV6a1J2sONmt7D20kKLco6VYYBFUXEyDNC
MxOyYwIBo3Il3E6T+iSZa5CFpto2YX7xHeDukJJMyTFqINys5yslwgrI2qfK9nAy
qNRkoYu2/2jaLZktu79CMic8x/fD4KpvyX/vX5zWPf296dNKzWMVPGc8wiTYkFYW
uqhQboiU95prxRd+0FB27k0bMvZiV2RNyZ+y69/Sfd1O8KUQyyB9YEAprRn2TdX3
gwplUFxbaLdc/wCAg/PbINGwn7syCzaUe7b3X6Ap7pzHxiYPuh8UljYJorvg3p75
PZw4aplxuWx0d0h0Z57BBcsP/aXEH9rj1DW8P6wfV0HDQt+7gPzKaPKNM57stlA/
BrjgVvAz0p76xduqLdjUyDY+AE5s8dff12/hSMfk+TkogDmGfPQqCQudUHDQ4FWf
sSzPtAFw9eAT3Hx1TPzv0LpsyvXjfH7xB7qUxFeDw53pWbZN5icIRF8xNAPmJeE5
fHsYsktFpgiJTAaE5OwO1tmPO9AdE/cqFhZaqBAlOg+7HT0hwvStVJpl6dnQAM7G
GLCbqcs6uRbglAP52q8xb29sqxQ2Sjyla5v25FO5M90jsDsH5Wbo3wBZ2MF8raKE
kgCPngMikEVX5S4u7UYvmxA+j2y9Mjse1SrY/An1GL+2bBSGCELofbl9FAAoR9DG
mw96/O9rOodVzd/Llr18Zo611E3NQFP56G7g2IfPKtkB3g1BcPgoAA+pODIHbeB6
aWWT7QK9llssKTJJPfYnGrzknTb840ZTH7c3YqtF1+KZsW87thZHab9hPphSRpke
Ff20WW4EyFQyZbRGXgMaSR5bhKCV9Y4LdfqN2r67pyaLk4816X0ULe8490bkm0FV
AVWyb4HQsfpGr2p2xz/uQR9GVDyhXK0coyZx84U5jt0gQUCRk0jyjH0kKpCkloZ+
3ML1Nzba2DQouyizGzeMsoFDIYke8vyh+lxAk8RQJSlib0KVE5/UVlP88jGeFIRV
YCoj8MYS/7L+D7gq+KTkqonusoLSRaerBRc6X2Ykz+xAoTJgkj0FIgPEFoFCz9WU
O2C30aSIOFYvLDJJsqulCGz/sWBM+TQ5+x+Q6/MEVQo1/2Ye+7kh7ouBKDzxOeqy
0AU5keM2olkOTuohJAk+rAQnW9vg4tlaFhSGL+9gtUVoR0AbxVE71FNeEjYx150t
Z+CFJVKJd2YH2JK8WRWJtFs6/m0dR+UqZsRYUjNrPZ7C1apNBxj4/S40dgHmDV0N
Ux9zVdxbSrzGAzHSJjGu7xkHNi9oDtpyim64YlBb5ldbnKar7Rf+vbxdHFtmP0Db
4Kqkx1t8wnSDYlNGQ5fHpRCeIJFomMEQJLhqF4e8ySe554R6ff4SGKFYmvmUcOqf
I7f8MfbIt4NB1VF4pWbHHYzE8FVHMjM+fiqlAKFa39DoItbG8NU8OeoeVLlarx+W
37LM1Owqske930nxQyEfLuvkXThPX8ksyvX+bqD54uyux7I6zkx6ghMjN0/EK13U
UQbXXurukQTbFBDNO5BtrKqZ63UETnflujMOSDek3xoiLHVXqH8sq/JkQpSct69o
R6baOYE1sOG4vwpmd4STntRty1HbLPTWgDev5/oD5IjEHBdMrP59tIj30/cLz1CP
JD0k11s58CCbVzhJ3JIL3yOB+wAENLXIOXQ10AjfEw2rMht/a4AtJiKei5ERmRqA
5xM1K35P56EuI1guwtdkJEmXSZCzmv+BTOUsDtBTS9eJlSJEcHlW7VmPuIq/uCNW
IYbPLCOSPs7T+FgxngOVJO662WuAR1Puxnp7PEkijUjPtQHvtTVPOmYHQEdAj8KJ
GTIEIHTqf2cJVLiJaIAK81ZTkG3apEIcbiWqZJU9GKgUEtlBBoLGIPzZPvqtH8Ww
tuoGt6IkZLvo6jVvBn+APkvefNusDloDFvMFY65dDhggWwuffG27fquNgvVGlCRp
vqsI9UApAIkW8GZWVEDs8zunnsxhgNf3CeAYjxFVWT4G1dBRDqP3UIGNeq2xjS29
oLlmR3gV59v5coRUtDhNg+JQKivS4RRXc0CGriwTseLbpfxlk3pqFj31xS+WwiYp
8fMp3m9yWJ2tNZe1+50ObG/Ied6DOautx4Z6+gAGrme6U7bwLau538jym7G4Q3dP
ruOOr3anpBaTdvBjDwhs9aoiqLmmmhUPVoQGGaUCE0EQwnqhjL+TboVtCniHwMWh
sYgVAnDI1DIUueqr75+yhLtFyLoF8dNyKjyEkmNotOPd1Fktn5JLPkxRfYYh2KHx
op4919RMnTusm7QubwBesKOpTa13jTgb9gFemUbrJEpPwVEshieWujqJDyfxz7qi
fwPAGWrLTicHntUS63sLScA9cKvxZ7ZsxC/csQH+NhynA7zaRq0ylCvW9lXHI+Q3
WzePV6woy/loU+CkmyMcqMbb5qkg9DHT1GiZdcUghVWs09rmiPU1qqQ1wUxnSgzq
KRULrYd6lkhd9QYrquWnsXdl5v9jqHAu+Q65kdPGFnS2n1OnwACWnrKl5Of+BScc
CGGM15vxY36TI0IjCI7BC7YFtW0byk0Bbn+k2t8QYHoeDthyU30CaqtNWU4PzoCH
8FzBxhHm4BphIk5NZKeE7DrnblZFgeyO1T+3Fo+wX5/JCQ82V0WbJxnCbmRJ5jOO
Rxde5Ep/IZV76NLE99K+V71iMrvnLHXb0PXbAdS6ZfXvQfJtPcHjvFU0qxiSusbP
2YJHW4nLfoNCSM2yCCxapjnlDrXmNJXu+94E0AY+0FahbOA5BmIDj5scE2aS5Ep9
PZ5iDNZ9QfH88ynvcW41Rc3Oe94iUoC4Qm45ZjXdw2yU+L3x5XG69LtHmdhnhKH7
djcvcxUceq2g3JU+EWePua9LkzERVnrOPcuVUYo2UdmrV1PP6JlK/PA0bJKpgtdy
l8Qq7BzmHJitgUhrOKMUcouGXBgfdI8Okv9oHJx6ef7uILLn0IL7KO+io6cNOQ7F
epEH9KsNt+o9sHcohgIbV7tv6hZMyjMAytdDWxMVSDj4MWHhKz8AAKpQ4lAptJth
q2bTxmEs2ysKoU1Ana0LGu0/IQNb7KUMtmVu2fvCni8JAV2DnNaxJTlvgiTRd+4C
O8QZN2otHHHFkcx4QSxgQ4NcBVjRlVaU3raS8845wP96AYTC2FqOlR7OaNYzwIRT
NAn9TpJkpeudGkYsDVVigx5XcTcwItW0MbA3L+dZlsJRcoIwFiAZQEpyCcN6G7Td
OHJXW4MYF/PesyXPlLvwn00BSVCyRbAhBKoKrtNXl3PCuI+25l1yFQgGAWIJTCTT
cY0l5rndVNGeNUVqfTvQkv5N7pCVsGAhEhFbGJhxhercsO3o0hPtoI6p9R5klzPA
tjbm0wEJoTWWMGERPjEK3o7gmQfmwQd16f86JHbZw89xzEDdMT0TKO7rwdQNzQZv
+g3nNZv2xAL+4KhnB98rkpJug5kDrpsSTNPDvjeOiICVrNVqFisFX1+uaa9gLvg4
cXXDiApJcxuHsDrM65PfyQKFRrkbGSqGdFDSOKTU232r+FTzyIYjHxkr6ONpdxt1
BypSECDrJLjqCFLCvtrkcGtnXNizaDkkOgayy1sCl+oQt4+VjE7ne5K6j+7F3UUt
iDoBwnTFvBEI5BEa5PZuygaD6L+zpI7vVGVY6ZA4e9zOMv+OvQ4ygbAflNDM+p/W
HIoqrzzIETgG3tlTyCxeJdrXAMuS+KUWEipG+sVy6T7Ow9Rt/1FigtY1HqgZZ64f
DS0Ht30e6CfKhVcZHmvSNJfp8N8S1J0Ov+UTdcjyaDqfISiAv5OJRsNver2FQKaz
n1dGu23S6UO1aQUJjMLf49luhdCM8DF8rAcuyLP8RxDKo1vKHebXgHhkAMti+K5n
wK3AhNor4NhO6B418rcen8ze5T3bEDb6U9TMXchxNy7/YMMwGLTT5I2LiRfB/L9z
tnhKKms9GOs4k1ifM0O4egHs+Tt9xNuUighu/0EcGzDzaVbb22+6K403qaiuE8/h
Cafgw4Ih5XMP7o+/Ocku54ljFEUqgi40q7Xy8qI5TY5Frwujkp5gyDTKWURNDqC6
yUd62uSg3tf0YiQpSYesDGv6IsWi7HqGjHiDLpGaIr9ZCJCdk6aAgdBWr5QSYhXl
vj8OKzTpmyH79jI750QSzMvHiHzy2dszL+mFV7h22F3dSmYdke3yWzNE5ywmVNfm
uYTX12kuYbSXuTfsk8LQvE6MLcmOn81y1s1ybBb0C5ujceaBMnvNuRPuwhhfbFuA
cJDRfOqWteaicgAYlICsbRlFob0WLlxaSoIdSF9Fgy09soF9bamdOXuj1SN0M7UI
IFGg1nWWTC4e2H3Ogs0O795TkzhyfFZU9JnbBUEKudun66QWlWvnCFzo7xqlB4s3
gy2FiSaVxPeDZXwlUP4CeDo3NQpb/ENSccmTAREakBaJK2hV2iHwsE6wtI0cUr13
hIpxlNySnguwxvF2a6CmKQVtlazojaGaCju6jtSpvUAj6/IRO0GFdqVEcQq+g5Wc
2xHgqY2R/K7OaNvJudTX/SreK2Nnb2Ir8tIzde2GjfNeJg6jKszfS/1EYn2DahFf
B4O9bWL/mxH+FGZIWiuL3dQ4Y9Lwmfnoyk3aIG/S0RDSsjdaVdxo95KXYp2WtZS8
/BAMYaPROSovzSdU+o2AwPNnDSyZgZQjR610AzL0ktALvuhPrXfw/Jto6CrKETfs
vIWEiYdtaLtcnRYd5eeJx6+lJxKNIwoZgBgFnfxM8Fd7Vp4Sy3cLd1Jl3OpfX7bF
+vMjf+ra8ITConeAKqygjN199l2gDzEYrZKqf4cAkju0siovImfQMEveZA8qx2W5
H7jOKT+K8f1IZ5NRN8HRo4PEhs7PWfI9MU4+blyurYsVh1t9eC5U1dybaUi4dspo
NY+XJy/T3Hd/0eofce1I2KKCdFveTTYHUWU8FyDBLKcXzLlHcGuCI/ox/PvHIRq0
9rhhEmRUUcqK5QC24TnTQFXvv+h7AzoNQOzsdlcGooSdrqUeSkEZ/IaNhbL2XfNM
9dmSqSwym/rOLMrrNv8AOapBkioCBL6Q7228kbXageNZFakxlOuxceGXOAV+oP5i
PtGB9iyHIRnIL0DkIPIy7KXbE4Dac+YH+7cpWNey8qCKm/mQAozFCYpDjbrcJsZw
h4jvAC+LEWR0whr4g1r680lfNBZj9GmCqnHDliqE6/Y6nJoB47AvAow/mNC4h4pd
awi3E/vrS1YQ2qLZGZ1HVPVGiibN3v6PjFNW+gXy2D4zOh6PshV9aEfr98BE5C5k
jGDE8WpXFJERXvaEjcBzApMTXw1MfecSnj7On04m5Om5pkr7CHRVml/frTypkdYG
2yefuhtpQc7QjUZVVgWkzrpEVBg4lhMQYd13Tw+EaoGZkQg1XxFIEgBYwIJimcs1
lVykupPIyYvAvj8183KlYjzmUwWGVg+blzMRzE3rA+eTwUOlweZBgu3rbql4QOnI
N1zg36SPPLtZBLDjjA1jYZ65p8ueGnA2bKEg9gXiLTtumOZ8ogkhfQMo+eLS7OHr
VqdJi3QXmH+Jgqg5vjWcrJGdZFxT6Vmy9LgutKJ18zazQtJ5ebfUEBYCDY8CyE8y
mPI72PmVSV1J5muGNguJQdy3MHNEGPGAI8m1z3lZTAmIST6wGJAQlPQI1jqZoXh0
q1jREX0E13Q0MoPxD+Hcv81AAjeN95vVamRSAz+gcq8vEie0T1Z7+1cZVLbvHfGO
REI/f44ImZF96ITBvJf9BPhGJiRwh+4RLkYErntBOzEHMwK6mNBqNZQflmG3t4Em
nB6+mNHRcM7RCc/5oJWk5QcbUsxwz9ruw1r8Q79MdiCmq0lOfBDA6Uwilb2N2oHw
fSnAHOU0FD9L64BuAUGwXirPmX67RE4MWr7tAS23XMiOxSgHTaf7lf5QZXbvOK0O
zd87TofCvLJRxvw391ZUnQA5/W+UqVxD0MMrdu9Vea52VSfZ1Rl6LlQdzUrMamLM
V21pusa45VZ0TAQK7eRAakTse8xb4TKlZQ92al68MUQi/iq0lTy2ZFizVoxyE6QS
cBNaUC6nKD4LiOsFIpEDIW1g3kbAjtIrluyb5Gz5L5CtujrSxlyFFhrDps1ZZ1MS
PB9NypL4UuzzHqVMFxgHRtKhRwoT1tNSKTovIN1Hm9sgAZfN3PfQ1hSEdWmsrwR+
PwVOTW9PjwRlzlE0/eHCIn6OLVir+YMAOhafAHLVfcjS4zWkXeuRFYKJin9RKeGk
m7tXD46bIRvAYDSYl9xRz5FeGPSTPsIow4SzrwFQDUOGuX1S4M5DEY0QbDfCaWqU
gnUB7GYpmNKI3N6Fs0QXsG5hLVsyPJh3UqHuoGnJVQB1cdfVXPFcYe2Z95PDpsgb
UUM6BOvQKFqfUgtZGMmYUEiPJByREgmwL2lgM2Kfyqf6CEoE3tVBZR7mm1KkCXVl
jL0vDHnzlzUQwT3n6xJXTdPg++EY81dUlDHQNFgztC0NzsJ0R/IVD/VraGxKxC7R
Fx9hiR4vZhFCqDlDIRNzWjMFIcwGVYqRU5pVDzerFPWHNPIjE0ISCflqVArOZzUQ
gWt8agQmB2F6tqiQaufeGFeXYpwGzLzF3LWMacQSbG2yw/yh1kD8yEAvsNYebzbD
Q4QVmm7gJIBTkWTcEUmLTzfs7OztcSshlYKSE4LxAriOB+vT4t06Mn21DNkJ49Bc
ebgW6RQwpKQhtciqUGSYjYVEVASd+U5ts2s1zdJb1mwwErEi7IdqB2WfhmTat3B5
ARdQTCTbn+8PrP4s1boCOIqCjFax053eBwaTb9SFikY/SXrqvQKhFeW6ADeZYiWt
PXjhURLBypPs1+B/eoZDF6+ZqDNCqXVxo5w1awjNY6lDNMKLSQRGX5flxGNPmCo2
dcS4IxoGrz1jYOstAsrRhy96z5grMiY2azpuyOZVqlIh/MIlXl4uIH8Mf+FMhkJC
JpR41vaO+2z1+JjPRFXYToZpwmcQmoTwxQlAVgKn+kWOS49bvhYjy64ldy7+Ha4L
U4v7URC7AGaWp2+nZSYsYMGPBYskAiuX8nmn9wwmSYohrK/Dh7kxKDh93HbJbsBP
yioM1aGIX1fuQ5KPEcynq53CgvEo5dDuAcEMk5uqgIZGx0Sen0PwK4bJbtVU3glB
bepNVHpyGNATyGL6rfI0f8bhvv8ZkrURAet7+c0eOFoBbLfj1KTOE++zKRXfSs88
BdBl/Z/8L9hicUkrHRAOkxOgIRvC4eT0O+J3ylu3edYnHjLZ5dAXx3nDne/+omzJ
sj5mtT6Z1Tsi+aQu3pJDhyJBoXZldw0ePgMr6uZKcTbOy8EWkUAgmDsm4NN8xvs5
KfHZ5tI1g2KpqnrmpCjzgXU0vEKRoTkgB/SIQtjj0jOI2fT7gofrNQgm0j0CTn2w
MVutVjzZanZUY5TE1IspiaLPEbsS5NBuhnIzniThE2qSTtCJ9Veybo/9yn7kUbCS
mZQwwsG+GtVbAbTO1P3ycVNBHF4kWN/M8r66bt1xYz16j8FtPk7cjrLpTafAXfIf
NUFmjLuCxFFfvHqs6XgRofXGk0mHjvTxPVvCvTtUMov2UxUCh28r3Sw5vePJjeBU
5ShWwy3B0XUimwZKc6vuX6qIK8vjBkf2eKC3sHS0rD2SvTeZCIWCUF0VfNKdceX3
38QC6FNehFOEx6n8EhRrIfEn152I+XxuLZ6k/teo1OFMVNgAJl01sdFCGkdteF/8
Uz/vIZsmGDH2GxzmgIoBdhCXSFma4VbtY1uqzp12WEpVdIb9EWB3foviRgZgabmu
OHCzyVQ1d1CM2Q7Bh6nUzl/7+aZKC+b3Vx+NzBSxj+X+Y0ZmNlj26LAWgA3y70Cz
SVs+Jc9dJm9BjfqT5/uBDmwG50fKZjWnz3HxMsk4XP33DD89WtNVGMCs4nFIr40s
XFje0zeWCfu0YZnQD0jdthJGg3Gzs7YAp2IblTgialXNg+qgKdilVlZQD189nUhF
u+4PKJh/Pm5VrVAuiZ200pEayhDAI0mX/PByMwhGzAwnNh5GRUk0nJfAeYkk1D5N
u7l7cYyR9rZEGpAJ0XIcM2BrfMGJMYTgR72rLhuS1S7I7nF2XHLmOQ5uPJoepJTc
A/S5s0ofLDe89V4iH8OYJoyoiCw966elRUGSt8sUDd8RNHqcg+OvEb17hiq3269h
20/4bSSIrwA9MLN45iV5iv/Y4+cfHFsKGSnGaf2nLHg4qsYJLrwOKasU3TG4ohZF
gqcvUSFyhGJOEtrJP4RUp0jUC7RpQgyPJOu0Q8ICI6aMLCIdttSwIyf6n1reb33i
WR1rtaILS61iaHQqMaONQt/S/3g28IEq3+RC1T0j9oxNV3QvH/Y4KDDruFg50iGf
EqsMo2Ipo0+SsK74p+4zS07x1uWDsLkLmv6ifxteCdwKGiivwtGQx7p4ist/zAwa
ekKiEW+Dpk1XYBHOh6JUf+JKx+jsiUjgVAFWKtSal66/MGgwv7sM4OzCfUiDeF17
jLWoYH2flNJCnX4RAiy9Wko7P1uZh7aqA5vh8TwebGlAiyK2H0nPA0qj9nM+r9S/
/d9SI2Tt7qrtA/xNitZSTT2l2SCGAMMH9bE2L09KSXcHZoL0N3qHgHilBLQxgrI8
gxaK+bQtEPons8N33hGO/sEV3m5KcviPvGztAPehfZt/PTBVTffNUPPp3sE8fQlS
d6//tkIxnCR/HdKJGsSuuKR0K8HDmZuMWyNg4QRFMxCcR4hVziHmjp/U6GRzxety
9GAc5hp377TE/vCug6W7hNDfUABc4p0RCRVXx/bP7ok6TaRMhQTWkNkLw0Xcb0Q9
jYg0rfc/GQI+hooJhYU4QuBBY5CIy00gfzm012AnZsORyYbgA56HB3+DV31LvIRI
hJo48wiS8b08JDNTps/Gq3jb/zGVHYOlJ5eHcbN6pDMo44szAdfE9oX5ck9Obk4a
VIIgHhvvDnnQA4OrSYC7Z+/51XV6X9BAXfmCsTa8yK5QJaPBKmBFhQlN+R1e7V8L
Dfrnt8Wu2E3j5B2q+tXHUBLomdr64PQFjjl6ZfGmwp9HvKmoJW+3EI8jPCK8vP7j
nDM6f52K5TpUiE4bClu53EgaSX3je4lT3mszwPlLH3SdRmU6Btujhea4K30GEU3F
GVVw/fGgkytxaPLGpuqAbYQanBID1za+8pA/OXDtDABKbIDgmIk74EcZZNwmGxuz
GRCfwqUMV3A/5QbERBtOr0tsH2WeK4qKvRlTLcuuA5UJGfpZ5DCbFwmGWfPnYpq4
BDOCCu5lTbi83mjpAjPubcruIBlzsdIhVnuojIO2kS6CwzVFVlsBNjP2uuPv4a0o
in8BHqgvFwct3qN8wrpP6RkBEzDpxVOGNBIDPx1WvuFZdtSzrpMmoikocKOwg3Da
iRGRrfMrW13fxaMDSA/G+KvLi/fzbYguxa/eRxGaILtAraVzISv5gxz6wa3jERXW
0plE7R5JrUQduY3UhKk/fZEBw5FsefgTyXONpANbTF2UYXMjulgwhUUsy/gTj6gj
XPVhzVz0WcXaM1kd96pJj1qRVLsFPDX1HEplBpoTr5LTh7calplW4KbTSbnIHGMJ
bzcmpFJJTitfLFWB0xsC+6iZ+/Qd366zpzDFlJGDTrN+lVANxjhyBOPw8ADuP/02
PDTjCQGJzPE07zKpp0bTeOh9HJt8wa/4fwDIVwmBYrhjHogNOU2KkiaQ3GY2v6kw
Pvw765GJvDAgobefIvGIuvjUDty7dM0uaxSWBBriiuBbcz+4gIt72G6pfPTsHLn6
N49HV/XLaIVvPK6NFJ1wM3s7J9Xncs8kwqsPUENiUT5sfJw7XwCg33wZVoLZPKiF
snM1xY6+eKkosaPFgjigKM3DuOUdTKpi145sbdfeBfAvygkKzZmqGFvZybqtnG/S
qAMiHsSjK96TR2leekzHj9+iCHVWxOqMjWNGE7pb5ZSWjfZstRrwMJ4hDb66b5tr
22Dfo6UmPUOZeKb99borZR48aZKqGD3QPupWwnBx/JtB2tpiYd+HdZxvUtS2Pdck
vk9bogKwaAf1SAUCb0rm7J3h72Nj2rHHe7Uzy170UVIXSo4ji+ym590GblziFomJ
UPcMCnwsE9e2mnJv+cUFEWZOoI3BW0+63Nqk5GpLpzRXJUEO7Odoei8oVfiFiSsV
MwNq+O8kzww2CTnU7pVKHu1lA3iV/CemeEm2MgIA6Roc1HuD2EQy8NRyPpjdGnPD
oKFguoE8nxc8c/FbJ5BLy27bxg+jsuoJl1+Bsq5GnuI+zaK2vNnh8V+v9/RaCF9c
yniK6cHyD1pk7d/oR8f1zaw75CfpdD1ZZH2HuGQXxLXBz3/TMkKsF8CUlKljzSN7
7Nw+dg3w5UV9jJB1bWK4l6PrMmyI7XoUFiP+QIzrqGiWhdPQYqMk3f6L03Sf0k0t
8RzCiHjn+MCijVyzhvz061V/GXxjq5d9ttON72Qy5vfSPmqNaTqdzgxVZkI0KOWY
/Ow0r0hL/6VQH6XeeRK6mg85wKYWOSHLXAu8WRqgSl48l9sJfg0pr64Dcyja1rgp
cSQ3b1x3Xkl4L9VaxKrnoTqynU3eTrsUJwjq8NDIkNiWrDngJ/VOzRlmimhxsJ9S
YaZ/RVB/yLd8PhUlbDAHQki/zsKnCouLDXv+3dXC9pMxrT8pPOxqPx0ViGi+VImG
qGGH7Du9GSPPSi5gelJEK8kNBfrQZwQQ9Bhwa5EdCB6AZ0zz3phncjGHrwdkCJtD
FZaOrTWEu8a0gLdkk5AI/o67gOG4sj/yNS555SB8PJS/tW0Uq/DGP6+DpLE78xuX
y2bqCACXbxBWARmmoAOTm/8FC/ex6jfkHD1eYoXTdhCsdDdQ3jXwBqc6+dS38UDI
Ffbvggb7zlbCQWLW5qqtKrw63SwXA9Cx6UTmHbwwg5ysxpVOx0UKbk25ej7eWHrk
3XjDcARK90fA4jf+DnatjFl63JumMW5PhfHvBHTBk3dWIVeO5toIZU9hmEpi9ujq
/s6/OU5P1n3eZ9cWp8iQGt8QH0xdGDgNQJfMDrSxwr+ASdpAiFzwRmKenkwKR9iY
y+5RhnyRCUOEt5bA+O1WY0zUEvVv43fHhmVhBmrZJ25+GA9CE4XlAJK1odOinF98
KLgcau5KErY2h2oxjVVh4RIcaO3rKglY4QmMXNJ95eH8GcMN17nyQG+iZhzid0pR
ISlsPKy0Rjz1J2mhCuw5C9emGUCifBz4fv/6ZzTua7gX6bkwxE279eABOyembqes
1LF0j/+y8ubPTHgKoc+49A1JK943PBNBvpjCUgLl50ooNhsvoZcQv89S49tpX0O4
b2YTxqz0EEMI92k+jg+LkR3gJYjpQj8bt65ILW6Kq/9DKexAXKNzdwyh1kwjJEos
loE41EdQd7qxrsbWw9S5+VH54k5XxEa7IsK7i0SVLHQ+tK4i9vBTL+w4pr3yXRTr
QKa4pOPMqSYr+2tuzcgoJRS8cF1U0uqCr6NjdSiC5sVUDJoeO9d4u7tNK6uTvT05
bv7CR7Ymc4JhK3EN3i89pToXpHkJWTGcABm49fb7KG/7VkLqoUL+vNJg0vwEyN1F
DPzxHB5jNnTv0kM4HU4fiern2HImJbuVJtMfx+52gLeI6GhSYbDJUOkaI1ut5HvX
S7Qtu53qEXBMEbhGRqnD2FGJm/FLHnp+VbRaATvIEgYg2igT3QWlfMpUyBp1ldRx
OZ9AEA/BhQO+/ZX8jK8B6W3s4i30o8Yj7hyc4rSV2CfZj8kQpfzl4bMWWjJg7CO4
544htTuiVVBH4erdagsXAkAKbaS6VVeQRbBec4jzbVy0a55prTUo9M7PjCcNtx40
FGA+/9DLOsvtgQuomcr/7TSNQaT47BI+r6iJdKspkMEwut6BwPwLunZaUgj6hXcc
A2aj3WUJTMLWiLeHlWeYEnasGsqk53Zki36cpgdKv8qWZ1pRkZ3fCieJEDp7vynU
moQu2DvUzjhQqEHFh3Bew/NleaRIfcboIQt1yNIbYjwSrybDRMf6X8f3f6ptbYFH
x5kdPWuqeUYR69RfMN1S/DX/66FlpjU5lmLENP2NXD2SZMsIcjuIwXbFzFpbp3zZ
Npm5mVnQvCW4rpYLbQAk4TXPs000iFO9FCE5kUNls4u0wD30l1RzP6Xm0QZHnyhG
YerUzSV1515TJXdW3Sm5g/WNX9MM55NbNkdR5mBi34NZCMBfizJR+htUcUpaQ7D9
TPaUItPNE8UTo3+nowlmn9gHlmFGUMm/2gn11mGGAaI9lTrlqQMmXcB3/E7wtLwJ
uTiEzPKAcLZyWRvVVJuoDHH4Bvxpyi0qrClPQ9y+QtTLiT7JZILfV5pTCCbZXvBs
pymiK0tkGWyy4mWVM4pEdmS7vLQikaPl2xIFyzLTqel7on9ltaQLsNnGyShR7t3D
1YfWqvtqGgh02/MzNTElOO1SG2WuWLJ7WZBXFnvcAXtlN9OpspbjUbL/6Czwb8Iv
tC8pYReQ+8OkRetO4QLGRi7+/wTw4AVd5kfyyR7+i4b9ACgV56uAqwjmX2pudlqe
/dTbaIXwj4ZlB8uGhVCGKLwca3IS1SXnxdn32VmKXqvcOnaCKUuqH4I2if0l9NKH
Xg3M76irQiVy5ubYAyKL0Y/+DkYeGmD58DUrf8UTgm5PZFFgHSgCQz9JNGOabTmF
yh5m6BaILgc/i5HjGrSGggS6g7YdOWuDKSeKzp6FLGIbOddbk63h6kCkOLmjRkCm
MsfBLkgL2L9QzuYYG/4UJpqNZ5bQLX/GEEfCLTOLoL6/Ef69XyRYurUuOfN6rMLK
rt7gdUAOyF4f5sdP4IxOyR4+vaZBpIu6/lwarWZdI/njjUwokFJAduLkXx/CPuis
1r8Ek8WOD04hp+Tr5fGSo4eEMJBStioP103cdt1cWk0LyuIawRqJ9vmp2ap2Hmak
O8Ge0kAIGJUi7MmIQhr+bc4h9uzaLZCt6BXUZRDNouEl7hFsjUTxAbcW6b/XEh0o
oMW9Z9PoXcudYcxMqUgw37EoThwCd6SPlLnWhRti0k/0pS+BJrfLovZrA8scnOPH
QVOxfVp1ZhNyx9NIdDjWqSMlSZfVXHozJSsCxd0dWlsS065zPsKULeGI4CO/io6t
cEcU4HmGzQ8fB2R0/r3p9XU2ptzhT0mQZgK53xLSxCde8R9zyCXK+IQIY3MugKzK
vtamz9upOcagqltFdqqpgP2Qk2Z+/iAm9TzQ5iWDva2mCaHy5WGgXMNJqDpqQzzG
YdN+Sj6kMaT3Q9XR3+vXLSc/zoFstcZd7OOrLsGy7S/ta4/JXE7jvHaPr+BS3BTD
u7F5Gmbw6ghaVBtejPOSsBNv/QHnjTV3//+m+Xymukc/cfbIuyqd7VIBdnodbfwO
NOdpejDeuvkb/va5sr/Rb9vfJeLpgbicUuAVNhRebHpmCZSWzsDAQE9E2L6LPZQU
zJsvsIHQXQuUE4yFBfiqT7FHBt4SAsqOIJqHDTrwxaRrxB4jiZMev8RVD9Vvjrbh
QjG4g63sESP6ogCucT7EOdtKW3+TCTx9wdniHSX2UPR4A2xnx64t0zg75JLpRChP
po0P1KyV9VC6H8SFwGTvKjnzhxncLpCIk1Vn3ECf50PEutyBv0VzL66z2/uk+vC2
uk6yTejihypFPB/ro1muGnRgKR2agfAP6fBiNkPlvTxsgwPdI1Y4pwipi+ScSR1x
Kj1aEjArxp72Q57zu3H5tRn1HfIIjKNWzc8HPocIzEKC36MyFIQ9TwCa4hTgzqqC
klq1ms1PyxvswD4ei+cbgJUVMDHRtOyd7JdJMEA78z614GWukiy+hr8B5IZ3E/rg
CS3lVrAWafW8tJt5oN6xIahfAib307jKGCwePOHW5F9MKrelwm8YaY4YCtjQddpz
QMUiJnAza2KIwXIC8sK12UQmLDFYqBwkWduMAE92KxPStcMGv5CvSWSg5kIixeWv
/mi4fhU7WTXEIaN7wO5s1gFqMeMF+V8f8n1rZFooO3aQ5h4P4OcI6p5VPr71k1QB
uh7VpBFD8FqsUDtu45fVxTfE7LsKtS9idq7U/ocSggZP7u7T8zLFWY7b430PEDHz
pTKV8zvYfL7qixIN6lbEhSyqp7A9IiPQvhJFt9t3FPrnuj1onK7K6URhWvjdvUIJ
hLzQUR8CK2upJdh3Opiej3nbPBGVZqh2fX9Kmp6dNFtyFYTMVYLXPY1lwC4bWtE/
649Nyvo0nWulxHWwx8iMu5KSOYrPv/9WYAjXvqxhDag+UMuMnQPmE8yM99r7qWZr
F5fHOnCDtIOkktsvrcIDVdQrz9xcdli2JZgp2Fz90XIRKXdCUaf2tOOeVLe8vF1o
WrOLrOcBPGNahk9+ghLvlREKCHnw2/biSq44/2D0E3RZzyl8eBkBw+G+r2wfI8Uk
/YVoEdR8aQxWyR7BJqcPLm0a6EirwppziMaDkaP4+4lV0Djk4KRs8pBZzXWemp7l
LREVXhzvXHOveAHxnPWPaIawIcpzsdFX7g+pQkK8PPX1vcpJOW874ukMmYkxSRDM
ICajYqpMd3JQ2gCoRtO/Jb0D4GPLmIMqot2r7b6Re7C1KBdJG+xlV5HeVdOta8Jt
nxYfUHRntLyVyCVzqteA3JJ54cXGw3I/1KGsRziK70H+H5Ye4jRcYawIYvt/6v1i
lUk9ovtDXeXT4zjW5u/VKab01gTXUnFvzNuDj5k2ZUq8dDAUjhhXuzegD/JgSm3/
lz422cZpbjUCd1WjoNbxieYMa91yr3W4B3YmbVrBfjstwgK+8Wu68rGEYVkT48b7
mYxzwcmjr91D6XB4Wcp28VRQI8+79/Yb5+yGK5MCZNNvx5/irdhmVjFJlwUjcfrW
MtBtTz0T8Fc2xg0onG4ERkD39m0WbMsMEa1zSBkeJbyzKTliZn6Bhda5n/nsbhuj
ioYa0Vl7W/bNL2rX4PrvKhROhBqMOZfifeQ0cgV83ArWjTHjpoTaPAb8yAVRDSUq
nS1CG8xqHWF1D1Nx8c+V8m6Ua3X411Id/0YWD2C37n7USGNqzwAi8HOQtcsve6hc
HqhP4YFLyeLH+gzNERDR5/OQRpCqjSgjo+TNWIvTZcefBi89F+09vpibcLUcPqVj
Cvqg4YYfpOTvxYMK9CQWJyyti5h3Uh1SEUHvr1kzDI5DeqMamP6Z/4ykZLwnAjJf
n+BjJiN59stf9XfT7uDcLMmu5ix60rMcqNXWxRHRM+bBW3yBrS3u7YQSIhmuJMgc
tZbA+fe0UE8PhNRKfWPi82eAyAKX4BpbvhqSX7dDdyYRSiyXZYCpVkN7g3EfNNF5
alcEWv4pQhdGI0cxvKOitbXpJwJYKgCW4U5X5uXILkVooPVta3+quV/5R64yXChs
VnsDQRU4T7xte9P1dc2BpXDniDQSwLDztPfjeI20qRrWDtDmjuOdV2zhYDDjAUWs
IfU2PjhyQ8SQ9GLlJITR68oSb+H3uQQuiXVrg5DV/g6P9i4WDra83wXenDHmXDmK
wF2/lXFgTH+0l92Fm2iRoFPK1STkG4Eqp3i1enzztnzRyO+PIogWI2S4H3ZWvOYX
pkCDojIER0A91SUli2hwfY9McxBrc6vYk3DELrpLLs/u8zNATsMfkLKCy789Z5CT
Dmkt+KLtkqj6qQl5ih88frMDxd6YbMCafuCV0eKWS7WH7QGmbaeiicvOvEEw9mqu
tJuAhy7FUzhcgZdpxao9E+DdFMJ0TvbmdxUloxmi5ytPRQ/d4KsphMT8S1rGBEg1
/qFfLPk1SnqoKdvM6qMRsQwr7sf5pxrWOYNawuKC1/+g54SnUvfC5tq2+1GTz6Li
VKvFpd0vnoIEDzp9IAGlLEjPqI6QQi0H5ePFBPO/sllnxRhJDUDuXc3rCmv1UIEw
u798UzNLVv1j8ZMfJJpzMufBfXnTzF9rQnkOvQZaC52H5KGwTQGEXGv5PpvWfYY8
sqDocASx4TydfeP5qNzS78Z525LEfvyizyIwxEQVx2qX5STSgLCYL7qQDw9VQr8l
MLy8ijG82dOIuURicaX/kfEK6c3NEw8Ajzf+VATj4L0g+Cbefp4saYEKy06L9j4r
LStGkS2FjcWRl54ly28AJ+//UgkaGS0+cc+Sby0hJRe/JEPBui2OZNeOO0ypkmbs
xKapAgxHESoSk91PeRvo5EgBwswg2+ITeL5SOP5Wsm/V5h/vz1ZMkzt6Lp6OhtXG
VjpVqnPWjd094NBryHJrDDv8vnlFo7StX0Bikj1ykAse9hldhfxuRtdkF2uds79Q
ZAl/Z+w8AyEhhMSgFFZUnuibk1anmjHpoSmMA2WXY/+X950dY26FG+/PJun4LcvV
AwguUWioTQUc4f6MjmOPkw6iuzYh+W/C9+BtEZZDnsO1anrTECPFqWMbkL9Ol9r+
vozgDJf06hDAJAkjPBqcAIyshrWB6tutIRl1DQTL/J9EJIoEr7eQQGvC2BQDi3v6
kCKqVclESOHrm/UUKgoVI0zyujlt92S8p/Ye4tL+vXcmz/rp6Q6IRr10pWbGUXcl
hdKUF0Rxsh+D21b2WrnA7NmdMoncx7NzmHfijHr08tU2ElejYiztyyQ5gCdM/C3z
LruZnDQaEYk+DZCH3ayykKaSfV5eMe62jTedaP0Q4XkuwQi2EKxFV9lBlhaP21ra
DjoT0CdnBSt4dhA4INnEGNGbxu5K7qrzv0w86zl7tQXEJ9ebM/KqsWk0gn67Hfy7
lSTu4AYKjl2T+nyohQlbYpnhMEobGLTTE2pSNLMQOSaELVotbn0DK+AFJ0HAdEBd
5ZU1EOyHF8gTK8fpntN66lJcSV7o1QSkhd9Bxktb3ZKOP6UcvnQwohzTTpqC1qDG
/plu0lAwLSVnedbfIvN76hDCIiOxep2AphVHA7Ln4bPvCsaoCFEseHpFYGDHiRjZ
zJ8G/b7/B9nrufbV77BlUDFdF0bfKqdVtbeIrK7KN/wgjJI43wSQkFsPHV4AaRdq
dVEoY8eLO2G6HZZ8/8nrnQyYY7emaHPNbOYMFeqYtjDPIyTwwApJct+J/fFDnvqe
pGoa6nd/vBYV1m3TlbaS/Hh5VUPeOhZYPy+KB1Z9E8jcFMv3xW4J9DwEtwF2o6Rl
W0KTWM3oWd6IBlqp29spDMK7U3zSLVmveOGSxmvYMcViBoqa5FR3qNAKowgoPvH8
bOvFkgAqV3izjs7A1dHW+YxqCi1uAYzNPI7XSo4ge3JJsLAD1K0qf890FFXVk+i9
yFCbH6nSgQR1jcq122XcCWvbsXASo8pZTi4jmVuhhvyeF6XrlYDN7FMiiuHqTZkj
y846VnDxWuWK4yoXVnD7vMFpYhX1eozlNM3H/J1e0RC8RbhhwwSk4000So385mMb
3GrEFR8q1zsBiXuuqrWlXHpeLio/RodlEsL2v6eqaASwWawzY9KzuTOD8q+J/n2e
kwrBojtWW66btTrDMDuYXj1If70bgUAh0m3mvfxsRxkKsqfut9YKHszszmGNN8c/
v7/46r8OSPawOLM5CLQhMFiEVF4qEH7uu87e1HQCvAR2WhqTqvNK8fgC9z99nRr8
b60JTz5rcndm8d+GKf0+hGNEfBoinCAMgVf3Z5iLaEN7DeDsMyXN2DQ/+nS52c3r
OzSC5ujTT8fiMp5Vw+2Czpkt4uvudpb+4v4hehmQ2pfgtkyUGhkAi67W4acjG3GW
9YqGu34Fe9OlM6bG1kVXG+9+PImSJV9ny9nJD66B2Fo89QEfzVBsj6MEjmSewvze
vNHvV5e303wB1ssABOJcK/SBCmDs0d2wySV+QR5TMowIMpiTThSCo7l0RFymQBok
hWFLYVh04thxZkyaKyVbWY6ny7Uy+4CmPfecz/ovhPnCF8gl7iSTeegL/229nKtM
Ngwtj3IJZ7dmS1zLaHHuXXnc8mimbSgnEMFksDzt/gCCMZ9LGrl1SFBxVkJ2+Iyt
qhKYpH6kaXqG9RUY8FRHDx/S7zMMLx2WBH2wIwEQxlvo9q+zctOzQ1aH4X/OQkm3
Myb+Lvou8LJhWuNnWtEV/nZPRuaJTEm/KKiK/H1GYymY5U+E8UtPlInti4cAY4Fj
NJgCNjkaCDgzvXab4UpNWlQZFBXCBig+qs0FIa1REAURxPuYVXtG8ISovntyOguS
kZOi3H/vpR6j6ZcYj1p2MaPgQ0kBgpF+vIS0S6xxY/dMCaCcGvxS6OJF2Wn1eZm6
c4dOJ7Zu+MHOJQL8H/UCyNCDwyy/fH2TSMjWuCpICsylasg0i0A6z5m1ng9B7cRU
VIuFVJIOpoQPgWeOfZ0RvZI68arJvpmVGlu7pPUz/krY/GzIOiI57T93dH+y22/u
s/EDuCTxbMp3T3Y3V7PplImb7KInIuhOXCctRaJtvdQjUqqMCP/864RBwRidmyxj
XLeZBhoKvNPJOg0p9ydp4F4+HwpTdfenNFcfeB1+OaOy4+ifI+T4DrBV4jU74po1
kUngcZGlSjES7lhJhYJXbyZk+Fof1pIAs81nKIq4PpwQfecVPXDYFNFVzGWlWlUi
JGfxxfb3SU0wFeGzYvtN7SJnZJLVhEQ0GZRiwgf8+ANZYjTJ9nUeu4objqoL04b1
zB3BOByz4Z6in5/XIRNmKQ09E3zL+JnKdYkZe/hMIc3UQSkErFumrq+zatuVZXB6
P6fzoASc788U71YlNsrm8uj/YNp9b9bta4d9YpfQSDSiwcHIsPfnIVy+ixAGPG4s
x8dYdoEVsj8Pm1JxCvtIhH1QhWcISF4/aYF93n7ed/kzTfj4ba2Ezmu85dNEfFrh
zGi5JvSu36hVB4vBaqRsNPUv0awfzxIsLYdfXezVPt0j4Wxqi7ySxl2Ae+yv/Cx/
KU6H+8XhhmbBOUVVnIG3hpF7lQHD8OFa4cZPhlOCoIA4fl9JJ56lyJMDKf9/hBXK
V6mdlx9q+PjKwP29SyXcVwiybrK4glMBA3wMrMi0ccIBNTsoSmXvyNiAtap4A0Fy
HbqG/FMukuecVsta8WjdbniYNDa7Om29uJG9YQ2ycHTTeXCVVD4pWenGiW+ZHjhd
26E8ifEeS//m/nPhUlIK3tIiUMt+cUNxnjjNbSqaojdrkXWqbaT26dpN2LYP9T9L
vMgKWpbMEHr0PnWyZntI6zPysN7SbSoUrAxDi4RewLw+uncdBBptmec77vxOtNZ2
02q4FHx0wktwB+ejP2e/6ZkJP3nsMSzlTdfKy0iHGe+FXicrliN4YG3dILezb2Qa
ba/73qnldNTrKlsTDchm4/IiBpyggIq86vxRZ7v2toY+EV70OqDBbTmFuIiMNFj4
EU6kdu16Jy/CvpzoTntLRGfeT8BK/M/egDkJC1XfMBYK0I3fE2gqdpmZLjIK7s+Z
aXlEEeOTqbGPLi0tsDdJvvwU22G02+PWFouERkemEgipVxtdUEzUcdUG1kPurhrs
5wd+YnBxIp/keTyPoJ9ih6MCgI/OI0MZqRyKZMX2QzYIf+Lcg7SbPtnC2GU7uKKR
KOzQ3TOc/VgMr7t9/naJu2R9FgLbztB6npgW1hv3UQCvCf5mbc6/h2uqFFZHK/e1
0XhzmamNEYaHvpQn5gyMO0X1XyAOJhFYkirFXZsfHXY3vwbzH+wVRYHULo6Crq7t
ODsg6F8VTp4N0zviPTGnRqyQxNINSIBUmHsCG6oxkX2InC+9KQeyfARtQObrJX1U
5Z5yMhwo20zKvI6GEaJgtMVuvPMzRV+bui10qM6qjlI0vQLpgdHhB4jPcmFBkdKR
0yRXAnvRzXbthfB4sj06F0VzcFTduPmJCDudP5VxDzkFrsDf+XiNFxfbT7tF23XH
OvBBBCKSOI++KZIN9wIE7Bbkwt5AVAPkgpLc3ci3fZsIm/k936AqdPPnco7tFr4B
EzTTCyRfwXRS/wLF2aukoJrdaumuS4iRXgnGNNYu57G2V8TlrI66YKTJsmCEeU74
2HM0z6KPQYvpoZ2bDLkLh6lhvpPiCwfps8n16UqMuvnlCrzhGDypCCHAjAaUpI7p
7cuoaJib2gI6jRzt4dKqxgjv3ulBN0tBlmK4/1hL2FbPTHvwkzihCz5Kp5/ZvTZj
Z+UMAtmRrR7Djv+S1HR83YVf+SMOcvdXwvoX+RCFCOdCzE+jkvil6FtqslsKEnU8
2gOqlJyd7WbRiXA/xV6Wf0QIJSrNn0/eflww+qFZZyESbQ5Gl0IC2FpJs0DyADl5
4plTVLSLaLaM9vb/feXzt67FxQJFRTIVbdyfHFINRxmjKxC2ohCODhTHyusRf9Qi
paQeNfubjZSrkc3qXpqx0RvVhAOomZNpFtq+uWeTWBGzoyDwWPeb3KULlRj1eN0X
kZ/DkPx42ctIXKlDNujvk7iXE4HUnUBTcGMLgdrzeAJHhRR9SAS6euuvRWuE9xvv
jFYTOFsOF7fvW8CFCVVNCCzDdkUWrbIYQljjsrcI1IBTZa6PwLg8kuhwmyhB04Zu
+r63nGhvSzwHLER3vBygatyBFuGDUz//8oCCoNS7Amacl/cbar+D15oEzewZKAky
VfCiRZcRV/pRfFmmqlSM3Wp8Mf9abvk1aojHO11DwYYuOWLybtklQkeDpbdgORN/
kBDuCoa/0AV575/xE/i8vmuT80d9bw7hG1XLIVrbih+bFzLMKZ9Ovqq2XJe1bkoP
BU6kcnBf/ad1N5tGp+1odmfGQoG/M1eaLZeylJUIQOE8ZG9mabhG45rkGhXHnTix
Iipx6oPvzDSdPDE5FDZCRyhhibjUXXHnM7uiPHqAxzJZfIDE8SWyYad084Hxr4M8
csVZYu2tTPWPh6znVQgzMx8yQZBzafZmh/iFvA2socoX0V45CHSuHKg31LwfRFXt
Xv4tA2t4EUiSamAbj+4x70l8Nv93YpENErjBqNOtxT9pjpx0b/8BOnJrPVXpGZJs
YLQ3yDrRTkmN4EuVOZgXNrBPhDeq3kcVZkTldhM/3gldY0QBDlPyQISEOM1zQlv4
0Ali5PjLN2NmnfMkCwWgqpGGzzf1EvMQ0F8+pXMsOtYZB/oJqVM8WtixXr7BrBkE
Ri9x1gmnzc6DdYv5Z3PC0lP4cHFuB6iTwQ+60DiNYn6t2xFY01wT2L6YW4Xewqe+
l3pFgfGESG/e1+wvS6lmDmjlb5Ma3tjnwdc8sy05MLj0lxb8VsumyhmH607MgkUp
ALgj6Wtf9vtam54ycpIbBFbUP3P9Ii9tXpppQTaGD+ozZb2ZW5p/kUMpYxe92TFK
I7rxuA/9b53W8JWbQoHq6kStAeup6TA1L7im4Cjd0HkKYjUZgv4/gB6Z8nLDNa9v
oo2DcW+giOZVAKOx74aFbSJC7Cc0IIA8TSvFVoVqpPH+h+HJtWdjUxcTrwMQkdan
PoXLSckN6KxueuGafJXACvQyazSW52Pq+YkNdYF3enTYUVcnrLCjOHl/a4V2fi2u
7uvdVSkUk3pw3bdKL1Mtk+i1yzbEovoc5ZYDRVy3iSfclkaSPqBKOxocOIU5HkzV
5TIwSjqFC8UpgistLpnlt6QUavBDwVwA0oNleXWvyRFvNobMLnLVHIvsilqDhwSX
SrEYm1D9U5g/NWjUnKjMvz/lWduCS0CDRAUMfxac4uvLyzwDhKavEpvXavJKCZFb
QMCpAsJR8HMXE4mNpcfFdOCwNT89H/RX8besVosC6XgpLL4VUtGdiZcVfQdRkQqo
Mn0mPDr4RSzy4lJSb0QVOqZc8RLl4DgqzE//j5YKV6QOpE/2tVuWOMgAqURSO2pk
SEsKkSiigdMrrv2evskwRnE+Y/aXxbfrRgWDjd2HXAtLAmrSVvUEO4cPTPKT5HeB
z89gJLSBsdvRCfGSzsjqelXlkgwwSozB7mXY9p2uRssxjFfnpVlDr9Lt8ZuGaKhr
x2crfI7FGRxgIc4quOjs96kMWEWz9AdGG9v6PiWxoJqkte861vFE1ADv9nMwiYq+
6cuWBRMk1c7LlbUxIKEe2j2CMjGSRyGCjdshobxTwo3fIIROWkhPPH1/3LqsiApp
v5vW27kfQveYdvmw3cTGla3vzuoePUTPabGJeY/hX3xYF3K+pQsjoaiAWBy40vDn
v7qAFRNi7z8CR0ZYPjc6+t+gA8/NT68LzXK3V9cN/JEmq40WEi2mDaZ0+edAcw4x
uFsLWibtXIm0/4L9PfMwxxYubC96WNCYYiS2DbxH8wrmgAOMdAD+guyP8g4siiWb
VyfEY7P5F5fkis4gCZu6AejpJ7UX17LMHejJvJrTURDDJF1ST9PE3iDqW0NQp9mZ
nvpd6uzY4kLRkxtQKQZgzZljOljI0wfer/fTJ6A0Gfxh460/rPQ6XANwkXIQzzBC
8pwyYFf0DWg71n6GguxomMDHfW+D84zUszFQsrjj3er7OrqAXFFYvrog6tEy6u78
dQEXERGMHqQltCKPLLH1DGroyqTiKABquQuICRYI1+oT3j+o3odKFF1/AaCcD6aD
lLym8sgD8HVVNmjNenRRM028J+padcHI1wLFLcngPs6wwY5hDB8PAw8SnAmB9U8w
lOU/d6MCcYBOWH1jDl59V/qs9/jvZHcxug2ZeBkgvrEx7x5lNEW1TX/UxrVlTrXT
ovRi1C5t7Mp5xRal2seX6Lw2o7DN1NM3Cdb2bJZsgaRGtqWG0Xnvb/CIPkOY18sK
1Sa/i289i+Z/789kp013qHanvLHE3rjwUo6xY7UjlSRkEQFlWWHrHiaBBD69dsOY
Ewt31rNSMTUQkMSmmbC3bwtCWOu1hY0BHWt9KSNmk4Pnjftdw738HMyMhPxhZnrX
6TXu5K+W9Y3jJZ8QzqfOECsJ9Z7gI4h+oOm0yb18s0ytQUo2DqWiYMybbIby06z4
+HkgzskmDK3NRm2qkS8j8Ya5fCmaXRN7bCbHVXS0oZk/5b4zh4fq7zlFpYqHS2oN
b2pbzKaSkQl4HIEPP41yN5DSKv5FBOpOUWoaeyP+0dAMYGlq60d1A9wXw0SE00yZ
CYuuSxhzwpWiUAxQS9T5a/hxgkJm98B1qz40AQbPiuvr7XU3tkRSbtEnpLoy36kj
IWqapZTQkb+VHGY9SEms+EiqnRSFXYudnXY8sLKJ46LppIC4u/A1jV5IC5NmEs/0
EVt2feX4Iocs0GjXXuFA8R/S3d6KxKkNCU+mKyo/bAeaLxVR4UaqonLtj9QivLqG
+Y0u8oVXsR5VYy+R/Pmwx7/12jBlqdyS2uZq6CnYooDw4icqFwo8ErvEM/OuOW4L
pDDgbajBx4ilj0qU/rUltD/+1HbNSlRUiMIGxwwr788YnYszn7a6dRukFDLtQb+O
odkI9AknQtGSfp0BGio3dSU6hlcFjP/i6GfrIGTYfglMxCGlMupToukAxVz3ZfPj
xEFDwK5pTZSuk+WI+yoKTpLhGvBoDHAiYyHTm0s3UmqwQRn54XjkHrJWppZwQNGu
MPN1dYhlOFYSo/gEjaB2LAi4RQPyzGQ2lAwA8FwilFJpVJTiZxY6RLwkHzjAzQ/Z
2YAqX0pg0lHCfb0+9y/xGwq9FBPfv0+6qiFUJ2sLNEUEGZW3dU+cHN1IYq6pgkZQ
LaYgFClPjW3E+PKnO6Vegs+S7jKf5PeYzKkp5OGRMSsorPLb30OL1otNCA3c45Eq
3iIiFw6yh4fib6EFZi5gBoygxC3MGe24MPJZQbnzZs4PVB1jaXlWoDH02nKWMHa9
1mfqs9iZS0DVGpGKhNdR7bt3BafsMnZ+aBt9/UiUnGZR5OAWPiMXGeBCBYuzfXCT
jcr5J1f0iJT53hOebBf7doat+8JBg+thgJf0eFmf9buE7CAS6Q24e0khMyuxAjhR
2SAHNaFYG1Z9fJAm2QDnlYziGTb+TZMYEoTeh5mLmRRzfXVUYJgv0ShldZAvyuPy
NwvFV060ECaHpmEb3B7gwI/uzKpOFbSDilFglhX/bhCxwtzhii2JaPAF5QwLureL
emugYNWB+AHb07OzbKZ8bsI+qieFZ9TfISs2zU6aW2FijAbquz1qGLr1rNvTM6ol
+6yODE81E39wcgBH+OOsyeBsDpRwrlKCzKOt6mUAsdCyCZEExh5azbiM0NcLRpms
juLAN62vIZdegtmpH45t67PpdOzXns4pvPPMdjqA3ewi1cAkZVDWDx36d9W+ZXWS
UQdVWh2yGCv1++trdGWTKTxMoWijPri8UU/PiZ/w7ZqzUGVyUe7PguZ2z+xhC6vS
BWKCCed3iFBjBU40WVnFe2oyZWvzDnyhYGQyjuY4n0FT6+hXWpqkJKxZBLVG2BCg
9dJtbjquLH7QmfTAoTWRry/x4X45F7IjGNyj4TilYDr4qZx+3+ouhhvIRF3C1n9I
BhQoa9uwFHCJn8MdVdObxpJlbRx6gIPKk7SS7qQpwRkj1SQ2VbuQdPgU4GXiuz8Z
QPkptz52kF7/DsJ5nn+nr4MJQdCOgu6ywTjcYCPdCRKceNjf+yZ4uJx6WFDRd1cJ
pLc6s5nOPgjK8+18d4TeEqYX8mMshvNy5IjY+f3i/pKm8tvln0N1fbMOYW+z5Kal
ahzL35C5YD4tqsUV1vwowrmh8FpiYF1cTK0WT3KO9zuzsZnOQOAtrXkUxzik0tyX
3iaIhjS4VVOjG+8orAJTNG8tXI4vCfoBUl/ucY78krP9DVtLZcJNko+k3SXx6+k1
iv3QIq8JRmgPDBXcVtHnAbS6C7hOv7F8T9SJ5Lf84Ne+3xf46xk9W5CCAj2aK0Kc
8i1dSmr9mQp1zHWnxhZfsWqKCuhNKJ+zFMNuh4bLH++2TuzwfttdL9w+uVp7ZX1k
Fw5oPZwG7YYUKMHQ2nurN/sqNZUFMVKN+20zWFoihJE0Obq0+qWrI4IWnZ8fbXQm
BtdnXTrYkx0IFy3c+OQOUBim+hGFvoRP0T+Xlf6EUzqGqgEjbFw7DKv0y1G+ffQo
Yt7AJlyJQQ0K4G5ifWxkYIC053HtQz3GDHL4Q7KBMKcYAtq2ygRazrBl9+41g5/c
dlGPUvQdj44U9wczScJ6bCZljhQ0Of+6TraTOgDeUg884Sjikw270HMWEHSqChlY
0lEsooR08nQ0uqhoQqz67xZMQGEA6E2PoQ8E8T0G/XP04enxeW3O8ei+qis+HhNp
MKkLxmhIWXu7f55BVEkXRMrPXgxRosFx8wPvfJKw+TOB4OKGl4kR6XaRGSKkXKS8
s9evYuFdpVYZaGYSyA5awn5XLEd4sdEqP2WGmYQDPoTHHJXY8Neygs0BtZoyjVLO
seeKKWm3AU0SyXCbFsqdB8g7sMkN/I3GDU/FdW5gHM4Isv+iGzaNp+huUbhORPEV
56tSZuIamlbtsUUKY2N32vPjGQOaJ5bxaXAyrr13o5YTjRV4xzq4/WxbQNiAD7Cs
V/zOIRWq7bQqlIEQ0XLbTizwt3uvW9/i1P7YWjQIzRyF28fCoh9i3RkDKqJzck3r
H+EEpurLzotl71Bn8W9sM4FbsVY5CJUc/Q8DDZ3VTXaUtvvdTscIVchc9wyGurlc
1JPSjY65DYuwjYb2CDTseYat+GxSlNtvebSw95ChGEwpcN1WM8qk0RSIwWABmOYA
NGjQxhS1hGwHKAU9yTBDP4jJ7977iIDYCrqR+5OayLDYu+doISR+4i1zU6gDxoFU
RR5R441tMf4/R9NsRfSrV0kzn/hSmZbTgLlyO2MsjtiH7mC0lyvkI9tOEJXGBCVi
G2VZq2EuVv1POAnQb7sKZ6O6GRgQ0Q3mHV+JPveOQgR+8eRe+I/zQikt5wWALbTP
9zgeJzjm+1gAsAfPhiPvlfqhP/h5t1uoa7XlzX8qtoxRBaQsIdf3x2PoYqnAtKSE
UG0InXxsamLXtOsEgN7kgC6UochQjW/0twP9Tq0e5Zji+CCWqAsR80ZkbROHnbc5
cwlk3y47ZIOga0DdP9BDel5wxzT673XDjzSV5fkKfS0FegyTCu0AV64nV0xwMK7a
/8FMeGyQOoV+TWQPTT+wZ+DvxIS+gFFexwbwt/dWcibcYPMnk68WIK/DTznbaXhN
n1ZBYOL1Vo2FGjOUJToIdyhBYEqFdQATEqG4rbsLMbaUUfzPTYlrkLoRFpgSXCgM
WMrrjN5U6da8DFa5znEgt0nPwP2W3PZuTXD6b+fI2XV+j1uUnwIJbK2ofsl12CDg
w0N2SqhOASnOrx+rmLKOmLv/oRHxhi+l38hG+kQdJbGQpMD0BrHSwj+3p5NE/zUV
xNxXGBUu3bRDG9nbO5DXRRWyAjBwl6IB2RoJqC8g43SGWYnBJcc3WkyXNUSkw0FH
5V/tOUCncQo6pi6JjfU0XW3Cl1ErK45tg6ySTUqmDUkidJD2gGO0WyQGyiGLOYcj
gpNEgWdCU8BKRyCxlotHTDGrXXCQ2f8o9drjUFQoCKRtOFSTj35ZjpEo+YwcE0yy
x5SK4vjdUdUmeKS0AVdAAMPFZgaqcZ4ZOhIoB642xbt3AUpfiTPsLNU5SOVTXb33
F2dKl36hnytn4v6jsTgQZO8ljycC62zDwcMPyCuuX8x+kccXqHBWynk6CU0FQ8W1
xch+CuOVXq7xXfqZwCvehvpgAOuXT4idy/qEst7WGxpXU1U/jGDjOUQWZQFUNuNC
VnbEdgJQM8tRHEhmCwhu/5Ril7dcwiICcP/kmCYgDHJbR48zPW1fv4noFfDbE0Vg
iwo3oNdqk93ma5WVy94e6NZcCIrpXEC1ICbaYAr6sZzMTPD2nMC3Cij4kCotiz3E
GCKhUxuVh/9qB/vawqk2Hrgf+QLgrh/zj3MHQNq/g3+4M6oPixflENvy85MEOe9j
VraKF85Vfoizo3fRKxVHo8CoIIyfOA2fPRRKtLS75X6zXi7HalPopQvhs2lnNGre
Cp1sps3vOkvAoyK1NfiiB2YeTiJt6yAf9cEmHP5AY6FOmpZuopflyvfeMbRLqj0z
Yb2oQA0vj2+UWswb9D9bNZPcBKqLOEQDM8nkfntikiCy0e0CWFLMepk2qYRbF0jE
E0eN8+8s9wF5FYS5n17l1bh3zvE6pU1FKp9nJgMLq2xuuQ9KcL/zV+ag/9y+Xend
/6K0BTSFraitavEtwPl4/1S2eW+mmK3yvKJ1I42HxLRtO4EHfZipc5kcLs7E69bz
SJTzI3FKwEDazO55wCJHC8SxPbxqBsIqVXdwQLykKrqk6lvU4Cjnt/mY5IC3Y3it
v9svAgBLXbkhJOF1IEQhWtqJZtl6UJnUEHUw3HL+9oURqqB6pc+cFVPrXwqozCNP
NjoK/i+hnMAGB8nJwr14nvC7m1WeDLB7klxG7lCrjBFrKA7TzRBjoO8rRFLNHG5W
QiQWwSk5pR90bcfKGKAHNMLSz/UIpQK4BFiXYDP/N1YqQphbmHwpmj2B5FNJxx7w
0wg6IdbV5PYnmOKeGJnoA23Wwk8INhM4XJqMfFwSwuJWjQze7I6Z26KiaATuOsgI
+JwjLMEPMmU+xkskgO+w/EhpTrrtb5Bgg/PYHwzVTPJr28HrcfPt7wB0XwvNs9jF
lQysJMOIYQ5RxJh5LH9dtAijXLalwka8R68yoaF2Smj1t5KhKVNw5I7LVsLh9SCD
puN7zjF+PtdwL/XNvKg3GqyE2P07f6GLLiky8ysTdkSsFjLPy1CX4gkf0oJ2TnZd
1gLCQx+HY0BDrOdRPQ4wsrDhcVmUvHimcQa0omWOxkjk4BmsvMcq8cCQpeA8zmRN
aaPbQcrZjhko3EDy3lzlt2pxSny4ImI0llv7E27VmbwRsqabb6RmIcPyT+BkwTwd
ifQK6Oxj8cQCwEPkdKSXSPiZIYbKxOTU+Lnh1vq/gp5JGruC7W6PI7yHVCrl8VYH
A414L0fPjXrpVKa7/vtE+jQvCOGC7hE9fd67TlkP4EREuVc78i44Kwg8f4xByJ5R
DWcT2YpL0Ad7cZ8yI0XjbIrLXYcmOpaIiZ11UJhJ3Tz+F5fSD2x8DKoIYg56SQyh
NMHTCJ1B/HKF2bJ4cXHpJ73tK7pYzcE5u2N7VT3NisZM4DgN4mcTduAOszvDuAR9
14ERwgIK1XTvJIizWgsTZ6GtU7Zy013t1Wp0Ndtn6ugBm/g3tHjocCA9k0dynzo+
d9zlWcGwXNK1W/Ag94y49kZ0Bd/H4wpUKPz7zn7xanMm8LnEnd4L5b3kpqNXkprA
Mrf6ZLByURYjw+ZXnC6ms/LSFyzKO0ywMbYIF1zbzaIn9ZJCBiQDU4esWQlUCqJ8
ybSbVOXCS2xdp24MJ1vSduH3jug8OxSoQjarehswpppZLtz3M0jjLX1cbf47Pl0e
aFf0YATnWgqfWT7xwa5XsAPLh7Scw1ltVlYDvA1xxLSZGr1riOG716a3rmy4plk0
qKvzUq9vCKtg0DQEs2kGLVXiXT/ta5EAoKjgkUZUbGpB4aQeQzcLGvVnvxDdr1Ph
Sj5J2eqPFQ0/3gE7x4KjwToK+niGGojBoqHYBrRMASiADtQAh5O/ueA8aIi2i5R2
MtY70ln1h7SPJbmI+OXLAOennfKsOin6AEVc0Slnvv4Mek8dkIdKuAqnXoSpd668
4yCYn+Aq5MtT77qls8sg74ALsFbabQj4P7YqnoQOOp8zLMQNxlj1gro49pVTUa/O
RolcyQ2yXJZfRpPuprlVr045fnb0Cg9nF+jQBJH5sM415RwR1Z0kv7uQoheBy0qE
0Bpx+0jbkMRcilY75yYO+AW8/kyValcxRHHdNhJ87Ppznxfcw64BfiFHdYluJS3W
MwgOPeBpnpGZpSFy/5qSIc4G7lOhQyvhDM9Q3n+3O6tUuBQ7r9F7/PfhSOr/+f8y
zOe70OZETEuRbcTexwoFVxXBonX72Q0NIuAWVjgAk17OukUx00ufwNSQGjo389Tl
uNyJ36pxYELw3JwXKbHGxbyxd6QFg10TQ43fORiQq7TOeaxxUvk3jcv2eU3dXjOk
rzlzlBftlMBiQWTQcawTXL5EHtmBDORwgbdEQe8pvamjnB3gaaV1jINP+KXJUAZz
O9FBykSBOAwm70/ElrBiOtLlplllbde98L5clkTqJ3j9nzTQbh5QHWQ7Wd56lqNr
i6rvEJQz7nQU7YPKp6EgzphgPth5L/yUS91jkLrGDFgYrDq1fVkHHZXqtPzwfniZ
OoDM75DeAnHhWZVxrGFhlZQUiN1oRmNEt0IC3+NDxyIHS6hAoo+NloZSpUSnpZiw
lnDxQvn0mn6kGhNz2yJIjR6s578cgUAc+nsQ9cgzAHJ3AJvLg9iQFGW4M2E3Q9JK
axwf1N0CHh90neRRBoqkzVOK3mKgZaNwsZhhnq2YgzdErNeT/o1lxEpcbVOKribK
otTS5DWa1J9pl/GGDUBGvTPdimgKqrq4ks3lMmrxJBbRbS4pdJ96AM6OSKkRk0zw
y/WVhCooHQiTNGTRvC+jy4sCELXTqlBkuiH3ZBeemMk/pFcwba1p/MljqimVfLu1
j31n7U+tephcUJlWUcpnTpEjUGF9atwQjLzvu3kYG4Lt7/0hBdLckX+X6U/hNG53
gR1AA4B1asX61Dbe3P+/mrY887OOE5h7HZVkoPtPlMWk5TLOohWlfapeLZ6z6Tzv
C6HAx5VwdG7eMbDwcuMPTJvUIoB75lLm7XELS899SI/0gANHLim4Ausm5r8CVsD3
x+0HrBa1avJJIlhhslyMmW2n5qUSznpw1yq+jcCaEg6U3byJL4FgAtGxNvWdCAF/
Bfv47ODIZMlbGyVsQtBNwIlHYFsscLYv+8X82MaeH79qQhVkxqojz7V4yE7JFrbN
QABLx/vAH3qXB8MLORB96S5kkXUlTL7tEpX9KKSrS0p3yQujpmYA5wGJHxjdNj0K
6FYzB0QYf3PY9UN1skg5qfoVoWpzcMLpPACC9XQH6f72lHeptGKp+j1Y/BOD74j4
sDRNgnzhGMO5YDJlcvB33P69BObUZHY3oCzc4JkA+PWdtlUu1U/yzu6ZJltY0yYv
hMljALIR/qbdp1EjlpdCEvfl/KwH/yailP3UGcNac2EZjnHRP3UhqzgEMGc4Qmij
TkT6FqY+m/ZuY9dfZ4DOtvxcyBw9R5TiLWhZUHEMYVHbok/T27WA8Jr6P7EQ8j3v
QXW86OtTsv21gVUcyvKZx7NsJM52lSitAryVrok9Ba2wbdBZZqoRWObN40vTWC7e
hAPRh0MH2Od66h0ol3D1TP0G48ip8hjYfsMl8QyeiE69+G8cw82b3+IoaDrpxCGX
J7/o093+qAhkCZgCk06h7Q2GNoshw90HKDVIwR4qbEBUXXlaKY8V2IN9Q/fDbflA
hSN9kifp6CPwKQv9ilRG6qa+psLXY7jGLYRmQONgcM+EVQcuMOeOoEuPCcc3nYyr
hUagc7QzL5kQX8nHwsLPnMr8/3/wNmdQC/GZnFfj65yA9RMf+ke7QfMKNXoAWAFN
KNSRQt2HuHK9+169gqRuUmNSR+rdQEpGBdKFm9rgIQpIvNlO6jyEUcRBQJNgZGE4
48UVMQdrCDhlE5iqk8DMaRentdtAoruOQvGpADnjQEQZpLQ2H7ExOiOYjYDQ0+bC
q/VZPycV1zuyr8emcOZ4XDiocxK4VPQU4X3zMsrmtPqdUWZfojtKv5IXFmcbkFig
D4o4hSv01MlphjjXwvLJyUvonetxt9a4oSuxQy2ku5Cw3xmn+JU4m8eLPUCCIdlk
K9hYnakageaq2AJQV8FrOOsFwNTl+6Tbz884KfvIX7jgLbava5NPYQj+C9r7JrVv
t3UZo2rUxAxEDJWFJcJr9V+3HBKqevFwlf0WlYcjfXQCGwwjyFSV6JsiERFIa8Qx
hLn+0M89gvQgFUDCmPEBsUYrjayFfswkEce0yUxZpTNJQCZRylURMIQadyHuBOv3
EfrXKtIACHvy9NPYApgtSv+LC7N00zKxNVzUFwfqNMtQGESBs+RzrSQI3Jf+jw7D
K+o7SYEvbXdymbag8YPBciCM9FQNf0filvXCtXXsOWcSfjBER04H/daDelRo4XPc
MD+rcZW9vFnoSlTQI4e8vnU+nqr4qPxJvJY1qt4CqXvNdc+uC8R48JmGLk7DiDAt
0IUZCLP11iIhLv/xpBZcofPZzTQ0AB2z5cI6eQD7b7sf0snBqMSQ5MdseClj91pP
iP01ru91hvJwKjlKZ+C+2/n68lJhP1y9/kitKtYaaCE5B6SD4gGyGCUULazfsdtk
J/33nBATt+I0rR7qANBp+p6fUZOWZdyItEKCJWp3rzI80kBBzVWSzbjhPhVBvkyd
XhGU9PGwf5Z3186uAjr/J/T1HV7mSgRTzqcuFX+X+SbBKW/b5eLm1PWeleq4IoZi
pxktW+MY/UxuIUVcagWNA6jNrjDkVMHGsXM+YvN1wSpljvIelsCkYh4b+BCAalTQ
0gVecjSsfwdS0h8u+kuugeglkIvIscRaA/yayyfsvjz9GOSd+x+dmpa/z+zuvQGm
LibB/uOpAweuOO5jiQ+iAgSBGDgJagZ2+WWIruO5TKSfu42TUJ/fPm2HKyFKlBTA
7/8JI6rEifJBtO5mG2wWra5h7ZsaEQk57193d7uB7XnLs8JsfAV3wLQHqAbJvAo5
XosEXcpLgEDyRxMoMyqv6HEWwW3re2yU1j2eucTyHWnzbPgrx52RMac7hls+W1eh
5Rmsy7YDgLxiaWCVzHu7s495Y6HPk8GGnm/EZkbR2Jo606FBrlbr36SJ3G8UZGZK
jbdVq0mP7rJD2YcLWlfOk4XoaSdVnV2YvdxnTYi2FwfZ/wGAm/7Zcp8JxriBDPVW
Z5vDPZ8ogWYTJm/ksDY5SuIbT4GBIpGowIyYZMJ2M8reRUfr10GwcYbJoz+7O+Sr
X3bkSayeLkI8OWHugTwBEMlUcq630y/r2hnqVksARtwRjBBNPj6s0lXxRFdRuDM8
oLeLLk6t3ZUZj/fWkdvFzoXXKLk37jgciCvAv/geD5yxFcVp8v3qNq7XBwB4WnS9
6nvabQsJP3slaHQdq4mvUkp1gKUUyinG8raO+9B8No/k5OziUK8aP+pkUVvml2tR
XQj3X96bz6LVMrkouzVGwlCtysSVRxIGhm4i4ekRiCEHG/mwofnWxR+fc6WXbETy
Im6VCUaM9EtTa28yget8ZW9iqjiMBMteiWSF5RyoOaGHrj9+F0KBcmGwgyMyAZxu
hJvu3/bkuTfRFJvLOd+DKmsLMcwQVvnw3wCipj3L5Y7fWWgp16aDKgXGp2BXEkdH
qloZcZuJOlvoX+EC4K5Ad1H7r2H+ZQGZ89H/iuc0CLlAnxjHiyFgoRNKwrKqcYo8
HbGgkp5z5UFSZIedayyW8f4Te44keiWncrxe0rKiU0jV4mA8U5m4/gRuOz/CNkSj
/FrVwVxwE3CY4emukhERgMiao4GMyCkKCIUe2EmgQDnQy39sjEXC4tfBZJO02/R4
3yNhF7WcDG7HlI+nW7k/XImHHmFIXNJEdbUOn4EijzsNe3IXSWDgQxfT/7FkfSsV
yyVYiLsIOltUWM6KqPtg4ou5FMlVtLgcD8erOqLvFj2L6812YXDlAba5L/wcHSaJ
4bkwpKlJbDdB5Kz4FFNn8Ov84mSgfFazy7yVrC/X60NdNbBGzYReV6XkU+4s2ndP
isvMhTkeZt1r8QAIwS7kV/gPwod0dvdSnkCXG0nScFAjsSflcVlerQU8EjfwsmfF
3/8S8bM5GBjrdS194aUrwZWQv+QyXvy8jzM3PfMGFPXudfg1KCKWRSZQbCbpXXd8
REvJBwjZkQCFV1y7ZGZH/YXgDn1LGrgEP332T2DZ10KSsr7JFN4sorU50zGowodo
8DlPLLRFlpV2BAlsoFgRjNZbt+62cUbqTZ9fUrtSkW3BNks1q48xDYs/Ix35B7Yg
5c5C3r/ObkRcXzsy4CWIlG1Zhey4nBJ+XpI31baMrhoPZVKLrLI4K0EbATaXSdzB
AbFvfdoo38u2os/u2AAKo2ayHDdl0CHeVxJtFCiBxxpu3wFBxhGNQgOxc/5yEKQT
sNE8lCMEABYFoDy1fxURbKzoOPVaD0LhQ6ND3DhJ74ZxJkweG8HMhqQ7g7sQOeEu
nXosk2eO6UtgfQamsW/LyA0T713KvK/+e72MzdPRZ1w96IzsfEq3HOHKMCzBwskh
qG4NuBAqSdr9MZPW0xfqB5ytmYGM/vyXIXgg50Cml9xwj1jbuJib0VY43GXGQzUe
G4Ps14gE8Kc6AuAXEz8m0QV9inL/UxOAoUbwIwfP03V43mcRK8sUcscUczzqrXy+
8JnifkfmL14SJVdB3sooubkamUBV9acn0SfYQbpAXn9uu4PpKLUcdOYSSADEZZfD
8EeZ5URREVyogeUU+5n+aCwFbl3i42yEZHum4DlpWpVDQDt6UHB+MkBgOMHvT0Tt
3/ZKz8+MnCQhm7cuXee1DiQgdxS6U8kpMiB70Vjef3NOrZaW7kqlMYefK2MAS23z
+9JCvo0Hdiu63wWP9O8er+X1xEFBjhgszjr0L8RxEX3c9VhBpNN3AdHu5FCz6N3n
ofFrpy8TH1pA9sZwOMrjfckAWO03XhT8efG42ipS84ykR1Io55XeyG4oC2eaiHfr
kTndG+OevKhHkqup3EdRy6VunC3R88xMca6A/QBz/ayd+vCv7IQYQtkMxMR7y12Z
p0J7RKvxo0H6ZwBCHdgXEBG1qSJSpIt5Ceuq7Z3Df8/bMXeGsNlDxYe/eMdLEkWF
MUvzTkCizsegJOOLP/TTQ2T+Dd8sNCYyKD8DO0nMljOEHHR5dBOkDJBuF1W6karK
0LqcNsWUx+Gm6NOkwYnWvjpEFUkfsbJZop3+SL7M9T3y84tUJTEl6uMEZ4gUy4L2
m6BYBuSwRUK3tgttFsYz6MgvxGbo/31N8AyzqQ6RAMxtHtovcTh5sS9jFhPWVhoZ
n5mTu/xhfug78nU87nG0fS5c2M8cYAttUNAyhiHtCChuxfGdovnkvlVFAI31N5iG
pjTzue1KVR8xSSr2QoyY3+g6iuStR92fzMCY20N0fBMXZapOXCgCJS6AtvAECWMc
slw7qsEqdr4orNGyj6UkPdWNajcjSRY3meb9FiObTLMEeZ2ibP8gbiq7gQrV+BSN
4Y3ROeTovWFem2J0b3D0mjZKzTNk8v9mvBaJOODS3WNQ2IReqVE7bdCEq3XiMCLZ
zYteLsqyo2BTKayKKwfGhd0iqH4kslV2NSvL7L2botHf1IwvA76C2SyVXePl0ufe
uFBj2sRUMkrpY5FPSBcrnSXG83gJlp5DIGyKfzyhJ2rWllvusl/3v3ujco+011xn
7SkiSbjSEo4iB7MroDc7miaZ6kw2PR30oGaNi+PNqPvZk77/R9WvtWLTi8VF2bPw
185dwVPdograjmUYQhmZSl7r0ej4HJpWufP+dlbzMGAHtBojU8hj1nWfSzW+ho60
8J+9rFrd1adv35LLiUjhZHCP8mT9B27ozz11mdiaiEIHEbXQKOThM6tE5YUfWtK3
nVGNZk3SmQ9xs5MFgPzsefU4MkTWk03O9hOLUsXF5yC38Sylc2iv7nF3yPjAPoGU
ZeF19GzlXj+UuTELDzgnStiTCmJ78vgOkOwmpSqQvS1vAPz3FnJjo0Bwn8sBEM9p
B/mggangTB5Cuyi05vCiBF+BDi2qeSRmnWZb9NahhV7rsBflUziImuq6NSnm5KvI
R48iyO0cSHM0AvvMjev0JW2egWOWU2Jm33Y5hg+s6fQvu7qzVwxGRqM23jqVTi+P
saC9uDk2lF2zT9vQGhQjmiEW+wMBw4kh2T9v7RLu3t2eMGDv21Dr5/OfQP4i9PMq
Yq/otPEWE6inBp+bY9RIXL+kBIxiNPbwYwS+WKhAAHpShqcE+dZoeFDKTFHfSwpA
lCWd43V2t1/QP4S13vTTqFcXRqd9I4yROsGND+bOFCuUpl7Eez0gxpUjwrOw40Lu
HqCHK9FayZAtqTVSCHw5D89k6ksdf6TZ/NmXgghcBQvoRuxshMocfKiBFCOOS69h
yOCvc+C07GctSfzBtMS/Oz61ILGwtgflk+q9dBJN3VlwFacCUitn/wHZsOQuKLmZ
qh0wI5+1tvB8rgG0gPx+eL6ZZax0Mf4isA4tYkxp+HckWYrGelfvCuO9sgm46oVR
OzQR5z+fX1s4hApR7k5lqIyFJY3Svmlbj+T3QWGalfEE/S6MXzHNDMYilQIZgdgH
AKgcJ/5hLee671H/C7XhSdmj1XqWWfr/HeCpZFpzvWEFrPXeJUFleHjVFVOw3dCF
m6AKTCloiNKPlm+Zjhj4oGP7O1qjc+okku45Oz2dmmKDcAiM1euopdNbEirhITyS
gAb3cHRHk6ENXpX36RG9xsTih17qTtyyhb/tDxu/SuJSPPYMl9GByxRTtH1FmO43
o9YG5ZwJT20EBUE/qwcPTWt8pl/0I48a4h01BRRPPyk2JXePNaJS36nLVQMxYP2s
p+nCRXqDYRtLS6Vp7PEw5STnZGBowv7RJPQqgW/ZVCZnvnYud5Pa48dgstTZVNiB
Ghqup8T7Pbw5bLanlacXDfBjIoGHSCNDdLcHbgMVMxHHigPQs7kT+j9c4QfzCkNJ
m2cMQbqPVZMX/plymOorKlewnFb2iWwLWcKtOn/CUiGwIYwbeTdlxgiNECKqzOIU
sZ/3QGg5o1faxv3sjPWpPM0PP6JyjeFJKKfEjITka0a5qlpdHQjbXP0VzaKDL6e6
M7XEQzG31IV4EeTfT1Vyoe6rb317tKcDWQXRSzmptlErvfFvj2TbK1dmsjsoi/i3
eP/rVT9+W7788sI0giUKqci5t6hH5ykO4QpDUz6otngF6FgA541huKuUGrGp/yd1
JQiCW1Jkw67TKrRhbMEzD5uYjNh7gtuwBbbeX8t1neN6oaleo/R38seY7n6KAxr/
6Kz/zPQPofKh/YaMSN2rf25Gyseh32HjvjeemG73q4oEwQhJ4Vedlqpz9q67bulf
bpW3w4ttH8ER4fKbOmWJJ9y211os9/+EfEp8NCBamV1jzXdSOsfTXz9hayd3QQ1r
br19puG1/olmHDNQwYfS8BR1q37u4NcPT9XYsfjmx84M8/nJK7jsocCjrbDpHLaV
LjZwYJLqckxPH/NRjgtenuLBU3ezHDU9Z5knkNP6P2Uy4BH/Dg7sWcXXECtPQGrE
vwRP+6yTJ0uM6tUD9Yy8ZnkLAeKZ1JMnTRIaJXwDHQz/0Dhp0kcxm54y73FLsPW0
PcKyg2kNpn8F4wgMDiTA/cmDwf1GL8qwAtkn/VKoPbLYuCnasNRbuzx7TufxPJMp
7PR+O8dE5xVn5tbOzexxYC8vJZISJlm0+t7tc82W0Ve9I1e0T32sT8g24Azqx5KK
XMMZQ1DYxrUdUnDEN1TLlY14eHii7H2v+dS9cbzsp5PQulf7838YJ2JZl8bDJSiO
C7VNNPx/ABalfmES8bV3vfVTLW7QvRh0lgX2VB4UE0kK8/EDGzziaUzB+WbJYmZ8
a87xhwRa+VvFDzN22bAoOEd70aPxFo2by+oEBlVhTOhYXqdmIUN90VlvO1M9ti1+
SdSQXByxVb6esX6F+Q/kOLe12Tn1BoJcP1Cg5yxyvtj/l0VZjfpAcOrPvw7lOVBn
iXfj66A85Vd+iNnAeldKdpYObfFWkRUI88NdS1RREmrRio8/JNFaMffEgQqki8yM
LMehIhDDoh9PVRPWcvEP3g1Ku2iHYquOcnIEJCvFPfoD6Y1as3FttqbvH1p3myv6
xz6G2DeNrP6nh2lxPLiwTRe/bjk4thG9EXwKJq1FjSEps+d3bDbtEHqUqITL6izy
2s7ZORH0oe3OArljCpdDwG2YjDsagKu+Ym2RWeBFprQQoNB8VvNB25JveFEGmSVp
kTvFjpgAWVKcMGMgab1GxPjifrVAt0sRWluwCLj434OtzSa7MCgNNeI1oBb1T4ur
cFxPoJb2DKF06icME/Ktco8U4GG6v25MvrZSxE5wDnItWLJDzRWUmAdlRh4Sw4oV
dCvajm+pTMjvG/RukN15GfVWmtjMQIAcbRAhusiqb8aKKmMrOG4RCBzhOY6bnGpZ
REG/AA3NoyXKFiJJoTwhs6jamwzYlTfNVcl18NVaZsJVGGq88yXjewj4r14mRUlz
IkTbzchyIA6qYA3yR3c0OZVqsLE1hkxDHLCrlLLZJihrvcnO3EaoW7ebqj/hKcL0
BVpxznwWmFZTC5kRBI7IPXBI+8Zt9xrcVPrA/r5DC4M2Ll1cggg49YPt1YEBMJVi
Snj1hIUGLXwr3dcftVJD68Di6ahMz95HM1lh3ajK3Tj2G1lJS6idcwoGHkHUrNfv
12xr0HboKte/ld2vEYN3VgVSQSUeawoeMdB8Nia4wwJrdcY3N6MHefUewSnqKJHA
YSvc8ys+gtjMplUTyuc3a96UkZJ/xY4wnyAEn7qesf1yZg1ORXHRAaDkiNVwcX2X
Ko51xsV75GVScZcv6glV2xTKnxRk8FNy5JnzNbFYuqUt23gzX7DnqMB+Xjaqk0bK
H7BebiEL0U7ipV1Ruby9AYJUUmEv4VIoxKcWB/vUsMrZAKJJLmY/Hcdh3caluWTN
jQ+bQbzc00Mvm4LGx+XS3PP+E/0YNb1l3xMUZcawZEpvBwo23ZQYeKHHHE4uzkIX
FD1hQm3ZxgKgwrLMCAQiqD6hb6UlioPSisTr6GUcXvT64z+VV/IpfTA+AAuCAsCA
pOvFIzABzq8Ww2dFr4Fq5zNCBsN1CAMYhlareMKXsKq0Boze5v3ypQBq+8DCIV63
8mx7OPAhvY/+lulITVU89lsaKP2BeZgMiTSJ3PolcAPQmVFB98qG3ZSoLT1KmOXE
QJgx0Q+Qsx0SYcMlPSdv4o2gYHZO4ATx3g6dZ2bw/pI6eIg6u5B9s8E7VrY/kl0C
hF0rNoP2EtvbqmnzluYUuOoN6+ylwfDz+Icf62IeK/23pZumbm00VKqqRh76saua
nJIgljhkNqWsrsjn6XshVuw8kaipYxgbgWSphzdms6/xfWNO3uT+nybfUhiWe3ai
jTDtIsqzhn9a1c9RyKpME73dlvZ1krxgu/R3eyrKOJXJRsU636ao8vnpz96FkAWr
WhIU9ZvkHLeo9ZwdQE0te1fhny3RGimGCxhVcJQLSv5+Le8/kHW2cXnpLQB1SNjt
31yXJUbJl1ggN0QvbU+Vxp1b47udpVeahFa8UZyRcCGSnm1F0ncNYWPVdObVufM3
+nyq6mSBH48FojXmGT9hpHCXRQn7Wvr7UKtz6hmu3QFdf2Bue/Ajgw+FD7Hp/vmZ
gbGLt+0lNK5YcuhmmvwKn0R2uMr163jlpNTJhc3k+Oq0L8qoUUN4r6xM/RRJdtKh
iZAL9+HMW2sdm6uCSxSEJ+9v+8FQXTYAFHgw+mX2OiJdx7wwXp09guHOHPwjlftJ
M6yvkjoyk1DNYrUJYUHxk1SdHP0Dlv8AjgCG/l0rPCaq1198IL0TmWK2TZQ66A/M
uTThyjnKykHQMOrJYNqU7kOJfgQqlUvSPmhnjjs5JnY+KfCAimwV8LPgcZqnR5Zk
ffkKZzOpK/BNshNLfV3RY7YCY/F3iqUAgf/PakUa+dJLARIO0y1ceIiGUDgi0eOD
lA9dLHROdcGpUzD3fFbnOX/bbgjUlhF29RvXJ1HoVN2ZC2MXQPbgN3pd3QvMjGm5
Nee7AX2l2UzVPCNnrexR02F4QnWsCY/Y2p3lAXHrX5idge/2yGISNpuP7GFXA4eW
qMLt1quA0XHUogx3DMMxiKhOgyvkJhIqeoKyVO0jKXTVuUhbe3Ffc/xiLVZotJ1i
ORLi3sjMJcnljviWQ3Pn5LT7pgohPXhhD1QFq9ZkwoOeD3Q6uOAtMGqbeW4yP5Ph
de06vkWxqjJXKwTPuN43dIfs049/cUPkKrhhZIi/nMb4yVDJKBtOO26Tg5uYcLvS
ukOVMHL9IH8uAxTf6y5on0zYuoImMUZ9UBLkEAJP/NoEFsZFrDiQbJVB3Lridcpo
j2jnjhghn3vQPHoP02TMPcIcHr+0YPZGpoUpIeAiTIdvDD6Uq/1jGzJuafXmWiUs
a5dGmNrDuUGtgVYdJbYmZtQqtqcK9w4zlacV66QtEbj4obuyXSpn+X4uM7w7h/7O
jQ8mV4D6I5NxVsWNrtZb8uqDQQZvBVSEvZJmFm84dkdfML4idIcqMA3wGgaftXo1
e96+5JRNUrwvQf5OQxqnFccfetEieA1vKk73LHpzGnOAGzRlCMZf3fiO8qQYM9r+
03XvA452T98zR56RdgQ/KdGVvU7vvBQPxbMwXDpCw1GcVP4MFI3/L78kEhqrwwNB
njwCbHNpYiVjyv2SE1JG/JhWY1f3aatp0daOlFpHPlm2NRmegYpQGwQsFzWTYkuq
+5rO5cwf7QxEZHWuqN9t2bcykf8iz91ooX+MCH6mm+Iv9WNivsfcjU9LcTb3rkmU
sw/vWepa4u5m8cGb4i6ltWc+2m+agC/udLafSH2FBxcJ8bYX02XREED5zuP8kPuR
wWwDDdaiZvTTNOSCh3HSP7pRQCkaf1kLgUwcCSr72f1RP1WdT4TRDEQ+WwoJI9mS
rmTsZqd+O5FP9CwI71FU2yUQGOTuEi6h9/14aECIPqRjKwmI3Qmx9wt3vdKRn1tp
lGSHlS8S3LNzCQviksu9vtT0xCqUmu0Ind6cJBtdCQ7gFA9Wb92fB32g3wP9CGLO
KLMPPAFFnM/p1ey3pJqyfBhlXWe5w/ADcIczjuDg5kQQdDnQVXVzMFxgIg/8maLH
lTPytFpx3r+vDjP0japfnEUSp6GQRiSG1ZVDrNtJIZYb6b60RMPLwERfUF68WHxm
GTrYsj/gnmNj8snvBRNdTcZdSLzD5qXx8zluD3zRDQcDI1Re2QOmOWD5pVkB7Rue
RAmqoaMG1PtgOaG4kvfbiSX9i+4Ohou3WQnCM+d8Yj64AWgUdCPQzxFhVQbkw8HQ
2+RW+XLzk6iZw3bhY7Bo5KAQjCGc6vZVktOnL2WrRGKvLCOIqTf2HrYs9Ok7AHau
QOJ6/0Xw/MZz4tE36qGOLJK+5PbfpghXtSgXkIoGfcrEy4mzsS2+9K882MfFJ5Gi
yM0MfPdwmODXiYT+7/vouZH6R3Z1mcbTzXPI1C0brw/ITCemTxRJQ1YY9mxFB4Us
gpVuNGDHsI2jOoHEQshT83sXeGQBi4N4tf4glDvqUOUxgSxo5y2bQ+YQQ661luAj
UMoNIFA11GYKea3ncAcpmLVo7raNFuUHmTgISiUhgYwiqukkVsEewbO3ZZD9/d9l
SvQwDzPBGoacxFw+bfy09/kdCZ4IijrkY9C1hBtUU6cDJhDClVfvx7H7/J6WF9eM
WTcp0PjLeNgYWBjdQ+nKMki5YMqbEFDUH86Z4rOcU664SyyaMlkq8KMZXvn9+KIC
/GOdjsiCApwl8+fgScqNfu0BL3QLcM/N2AEowfP5+OcMiEuHACyzKfXSVWInp6Wq
3qIDcliJ5VL2mus/iXk4S7YrCqBcjR+jO4f2i4SQhjQ1f+6G/v0PM3Mm55dXP6w4
Nq2UZ1BCUr3bTgR6ml6l5b6SEgCf+OGXJXgkHuvkZcCTAMAmuIQXBx94iak7hOmr
OGe1brS5ubr10lfwGDUPNbMqvvkDMJXjFnqvodF9XwvPoTV7F5nf9+SjXhROxy9s
eBDX6FXykgt34YtfrUHyLUBtQWxS8ZGzEiVteqTsnQ8arMSrpN9C2qsPU/p6v2y+
D/IChO6SkstWGgoLsZCNMMJN7MvbDMhuZ8uefBreoKD/Xayw5x908eKa8BTwdBcl
+kA/jofAF8EQ81KreRPv6yhWUmKncykiYjHuV2EvojAc+w7ZPjg+Ej1aFZTy/1Rp
QH7+hgaXFF+X1SJPcpxiyTpmSudBvLgrwPcQM3NcjrTYI7twZxl2WBNcauM+wNWV
EPPzn37RODjTrUlKa2gMevelWiLp0sSyjiSh733Ra+AoqUFRS6hfo8aB8do3J5iS
3V7j/1etV0UhduMKkAzjI1wW7HXwePe0+WXsent924tmArXhz9+iBFN1PXYh+oT5
C0fY7Ulg6QxrUtwLCBElNRPoau8eDI3DGjavr9rRFZ2/3xNznX7gy8FRsvPDruAX
UqR5qeI/FEisKl7TFQFRCnLuE0Rn0+DgoU1E3jF/8gIV73q5t0VotNi4+0rtKZRj
6OABaMKayKzKw7gCvWAxHu3+YJTFcrOooEoEdEhbql8fhUjPSeK9RVKlQ1/4Si15
CgFWmMDdf5WnvVzVNPWFzcrTB/oPX9x+H89oFjyc78RqMItoBmGLyiEPuWMCM8Jw
wa+XoL3Hd25QkNlYwuxVusjEy0D1aAUU4+/pdlQ7LQrukaO7j6/BFIY4YXdN9pnG
ZPXAfmSG2Q+nMz+X25d/iSRJJwizbJ+crjwz7RmZPe32yCOL07V2xxKiCcpX8jkh
9Np9BCaHzndlK7OEGhKHkHodTFMrgtu9Mrp4dNYZ7MmMHQQbjNmAs8kkC1LWLMTP
jQD+3hg8QMjSZzpgLyYzr1ECKR9Nx4su9z0XXwvmjVT8RsYn/NQg+cPrRkyOBV3+
Q2t2fWt4y1MT9Wx/NbrcoqNS4qpTgs1KkmwtTOQ27k/NFqvUe93mNZF5Sybsxdp/
D9TzhzXDYLF+tlVqvrM0etnbQZPlWcEQh+ZAkrSr3d20M/HyvDYnVUcG3y912eyK
4U+8lhLKF/QT5JusOuD3yQBPYBPAQKfHqKixiquBSUelKzvZjokPvqEVgG5cHN9T
QexujCwTjwhEFZljKWIw2hGhEcK5cVpgYa63ce7ouNciV/MPAxeiSbrH03XbJXMa
KcXIrMz2oLqN45VM3+hqRaLKsID+IvIMr5pNpJgJl0O2rjt/Z8lYQr3Hv3ixRVYp
Hx7AItQ5B5O86jwJcJXatcaEXHOpXY4R5QBjr7KORt2Q4BpJmC6c9FYywYMc1Fgj
dcauRT0F+tK89EHDGoQ7O5S5LqhJkAVCLYvyuaJAKE7LZ5/1q3KF6h6OozayZGEq
hq+MNq3+qr88U0MphMhQ4H2ueFfuCoDzYLWZxz3VIiDIMlEnaeg3fjhJhWMeT1ha
F2BP/N/iHvwZwtXJv/mmqutu4V3y2/fwxCiARw7bSwNYOJ+Ql2L6XMKbcsjpdUii
X9bpZjs2dV/jusJqpcm5QBuDbMXnLI+hXNY3QpeAwfVuJujNlRtrhljcq9gN3PZ6
ZldtPH1/Upz0H+chTMvUB/i51pft4i67OCV49+wzTZU068PKanR7dIvgjUsgCLy4
4SoQNavnm9vYXQliCZlzdkbc82a+wbaHV81g+xEairoV8uO0G/oZWcxpXvjImSM4
7Cw4oxjGl7tjGp33O+I8UCcj5thgLixxWLLHm2xZbfbnYUnlMREIKoInRmsyouWV
xGeS1XW67MZvP0m4xmVLHzk25/uD04tR1p7MY5jmQyYKuFaFbqzZL3z8qzppWvXk
fCzPcRIxjKPgL7tSmhGctPKnVUrg0w4JR1brcjQPQ/FS1RXVfh4ydqRNSrjSWKBL
vddS57uDgkYesEhVk7ntLelczkIfMkfDGM21GxKdv+2sT1QadE8ZsM3cEXvRKD6t
UidX8TzBOkj/WOyP+Bmc9qYEe6HtLIhzXToJrzNWt89qfWijVSjtBSLVvs4snfRk
IZpd3cHxr8pPlHnVW0TF5kn2f0Co3/c6PfFXpFsVWnuRkNhmS4MdkVGxyWHMVLow
9OT5cxZ91FTaATZrAYyKHD+d09gM9tTku/e9Q+j0MZDkGwCJyMluBCcwkT4NUxFt
MH6r/ydGpVYLwcsGjOT9r62jiERbLPn2knYlueW/aGG46ZIpy5oKztxE8vxqMYD6
81wgBefNkS3j3ddb86ratYids8o/5Dlang106HsPmplyCh7VvnnjVmiSoCcdqGZ5
H/7OxU+HCwpn1k6XdWQe/gvewDOC1jMY6EcYnnESTDtswuvOXz9uQhduv4ypBv08
UPK31IdBZiVYWnfQ9Nj3Lg1naLPqMR/W+WnPxPrrE5v4lwn2NW0J1h1WQsoHBcld
j89sPk1EdkwOtsTzpcS/Z7J9oFZJp9CtqbVteDlxplimZtuOFZy26Z4/ZSkRNq2a
1DYH5WRTc+U/AWe1868dhqLEa/ZNxChrw3Twij3V1EYg3pDhzbDjyuaXjYv0ra/I
AyN/6wuaCoiBjj3s4i8/dSf7GY6VfpmPhWEEYF6OWa22GoP5tSRWXcbDELzuV5yn
SqWuyp1WV7jRACH0oDK1hNo7gCEG07CUqHw0Xm4sJnP9hi9q5fadzBejw9aKKE03
Nf3kNBdaoqetMkixqohLBgiuypBi7z41JVFLBgcyUDomXgjv1ApiIds5+8Pm0sze
mz2ph71kGu9vyc3MfBJEIDKG4TArWNmNCSO9bEzlIXBlAxyscKqvnDGzuAnpgpIp
KSjkAuowikm9p94PADowYHKVpd8Kvu1Qke4wI/JSL/cm+Ykj29/sFWLwySQY94lX
QQWS4+2cU1st1zsLTgF/xOyDJ/f4ur10HKESsf8PtU8avlbpWSUS9agrNThqI6z9
CenTmuZW5Ql5F9MK/6cvfk0NqCcJusxS8V8oXqLDnWXdycLijeRWWFeNlrfED/92
S/bwceAtBpVDgYHKGnsxz0QDAShkI4jVptRoh7U4N/B+sAPQ0D7lUes7osLnorIh
1AoKiBhhq9IdNJZuvOWsZqOVQgmtUAG48U3EyfwHzC7Hj8xI8fC2HQNR/hknL1vU
ENBwPgrK+ksrwDHFcnhhdG9rl6dOJiIKDyVObE27d/tk7JzSZbecWf9jOX4bnFy7
GNO+QxFaic/qANaSOExhVkWAn/h5P+0mfmX78GBZRMf60o5vfOuFPBv3cqcYb8fU
DAkriKvs6crujUvChmlTeeFR/iYSt9lhK1GZ4bwqX212S+hMfMpjiNokz3hMhoaf
t9I8EWP6HCFDY+XSwBmks3Hh8g4GdnQ9FXIYTo1T0pyhgcZyzAT2o+HTy2UQvHcm
Z+7f0u/Br4wdMJNGe9CVzcvTAIOZXSC/DzsZ9TUdQSvpLDQTo9PniKHhbTSy2Sgr
1xyS5PoLw/yujVHhESCFVasQJ8Iz/SzWi8ixH+l2M39blCO1+p2I0mGZVNEBW6YS
8RRAWzOjWTKGHE7yIc3XkN48+Mzp6n4iCePUw4k3xBtnzcXxdHoRLMZnro4thnwh
MVGvQK2Hg7Jn9hkXSRceGMM9lCZnmeOV93x8lfLmq2S1s6t469fQiOyKE8oyR0HL
R4DPLdMqtyMmhdr08nBEDHEy+PFN0irkt+o9M13svhVBRY0BL7jdRjyCgdyu9hoB
pGVz5LWg5Gw7P8qilA4vUgmucuCSQyKIFH7DiGy77LaY/vxRlnZ6n0B+aKRzstVA
MXVsJN85eyX0ZC+KugoRw6u+zmg9atFCUFWC15hc9EOs/VJ7npnqp3nkkWYsTXDd
E7MpiPVjstD8wpcNYVrEuxNj4aMsPraLkVH1U7iMxvpSOTTzQMuoj65zueY2IVVE
1hzWs1uraCdmMQG51QVro2iEhzjOQQul0oLeRZKL5EtjdmQ4u58XGIv30trFP4hC
aZHy6+9CBUj32L9/fJ+YXs0EX8zc3UKdL0HsG08xm+PeesNnaziLU0dRc8L7NF2N
Ld3NjS8jKZp2k3+fgFaP8fxiro+iCa1G2de2pdiS7c872zDkutabTIQ+gXY4Gtmf
ZBClxzOxrarbo2Ra23fu3zHfQPszr4mm3zXkVLr19JTHM6A1PetOVXNlcsv/f3WM
/XFDngzICIR5ZdE5e19sAAZTp3CDA3aT17Q53MRj2woeD9kA3KfjapS3BO+XX3io
E4OWkNhcLhkiIDDhxoFfTcK2mCwc7XSyWgS9Ojt12D/ISjtyK2gcrWiUMKYEdfxf
WQwXvEwIf55mi6/AB2jJaBhTM3mjF0kGbSVCDxRSdj8nnbq5f3sfjkxceMKluAXh
upDR1+/4RaLYU919AnSbVzIS8mW5IMshrqPRrYhPYYTuO62w7mOgZFKjmmV12nEu
4oD/UGIbnxIBQh/5chXB7WypteYMvVfk1dBw2TwICnra1DyjX5swkWOvOhDcBFBn
8USuHeG28ZBuP8HvHWYLXR2AtHs19jGMxxd3/hbxpws/aOW2c0jl779Vha6ry1YW
CrCiuNSSqhC+Ii4O2oXOI60wnsFb2Qj9XB6mBqgPpIP3X2IOyFSZc2qcOpMy9eNd
xU4HeEwwbvq20hbrladbUOXpUpn+TkJJoduRQWlzGja6triC66QmMdvTgOJtudQ9
W/mJFPgDMQ8ixNBOhAdbs17PFI3MO0fjMcFl6uiTtkvDyJOEWRxGgjUNDMBzPxcw
ofo1PZicDdlBGredXBZNg61h9sq/agZFwLw9OmlFAAOJQFT+01ks9kX1uvmvopIp
nOxREF5/GwPQ6s5tNpIf7p844TLOb5NxZar85D2J9QA4aSy8TVylKkBGQiCT4hmi
WHHCuY1dXsEePcqUDiJX8MV7PJje6DufYcJYURSi1+kJtXjem3L8im5jnz3huUeP
T+TkWnDNmIBAive07GsBdLVIc+k5WoJ2/p084Kh0W6gtdZkzZ1S/c+PPwCKsHNQ7
Kl9lUkxWucr087tV9M5YzYwR5WRtoiiF64vnmeqMJtPDNDlGYs2lBekzA72iZq8z
ZY53mCtxSbEJCO0Et/NhK72MoRCo5pdxdU41W1VFYDKxRRnXCy7y6AVec/bc8T9U
OCv+UsDpYo+v6joHkn47EOw5Jzlltl5i6n49KzciNs5PS75tPT+zjfyQ8wx2ukqE
D2FtmlP9goVIzRvkHIu3J1af9uIFFV+BPqUNwz9YNT8aiukMzgtwjP2lKz3UfohI
NhyjSg3I7mJ0b6+kJaqq3baWUT2FMm7zF6XrCI45JzO8xQOryk6+GdQ7vhLBSitW
WDqLEJ/3dg6z+cz24HdNmWDFKzare0SLTaBmqMZf5vO80uzFnQ231VYrE316wzjV
jVDdlWRWP8blFy5+Ld2G/nj/URnnB1DSOCCGW8I6wlGKOzGA6YgEZ0MVaFUGcuzi
tyS0ZjbvBkZIAemYkKboGZhhMDC3FHyLiB8MckVGgEZMbxsUQtXzhRVyYNyVwGxc
zdYUeuhhhJj4zwvDxUmqUGFDH0W5D+TehmcBncZFAaXJaUNzKnU/NI/3knYcSc/o
exTXLyiaPJ62HopeDWC/Li+MGYQiE6J+whFCXNbO2UpvZNuahek2Qx0CEsc+ckuh
Ml8qr/hWasYe0M66W8YzzgR83lXwBhXxMCFnNaT/xfiPRiKPxNc7yyptM8VOPViB
9khf+EcAGaD6lJambOI359V7LWLSO730eHKkv/VZ+fTY7EOAAjspGIqIw6cnavMi
qOP6Y4mUQGy3Ytlo6H01mxRtoM3kLDAnUK75djIh2Y3JdysC5EHFlm2WPyoFoVOB
gju4BMVP5luvlZY5PZn1PhdO8+qlqQRRwNDNjnmHowKu2UU9v0fcHeb8cSQ02CAf
9F/gJVbBu2nk0kwf/CwH+53LVr4cyKZ9vHR2cTNAR99USpw+3kK7kuRV60BovT29
j9Los5LyqcpJ68t249RqPAsdj6a41mBWUaxojCZnNngjh96hHhQfgEk2/DcRDRcV
yl6EB6UftjppspxDK75WLX5uT4+ERvJVpYNuLdqH67mmiVxtFT5iGsvbSbVhljR8
usgwFIL+6VAj/U9hXYGQs1y9Kn3DzKaXVlwBtxJFUyUXqcTaGoVXPCRbySyc0Qa8
+gwVq1gVJJOhBIJLNGEyb2/LhNtIsodGbJ1k0PscEdbKAVla5lpiJeQJoP0yIUH0
8MiHbE11rjmrIbQTnahFn9zFelXCIbhLn44hMaGjn7obchG5uE4jGJqqYTS2H6G7
pKroulmxmQ1/3eHFfLPy+MI/1uYSCkpavO45ilmbQpeli849+dfC68B90L+HQZo2
T8h8Q56VQdrXzLBlgpjTZ00glavqAqJdiCplFpGhyEtZiSkAPek280CQQZy7sQBW
k7Q8amvXYKiWtzkEKKxQkpoBHc3KrAtY5iuRGLk7YCtY7Hf9jU68/mciKwftu2U/
k7WlHn4Sla0ftXk52FN0u5mxcwiipRxKReg7fSfTuJOdIYwW3FBDCPNARIpn5tHz
/CzWoz8RJ5v6PvYc8XOL8KvpQWUh3JP1uTV4jLRORcaEi2WOHEncqFjXAowrn5cO
gqWtIYk7qZ8qlqgXsd+LrYRe4SQdmILsnetyjtUfVQGhwu/VIeb1OQpPw2wswgN0
McEX5KHF04f1rNyVm3XbSz8jovkYibx2ssADFXL33W8iJ+1E19B7CyFVm/hxq0U8
qt+S8RKDRpXHUfwcgu1RVU2eMkAWOy8aJnabWZf/eNWgNF2TWlx0neT0I0FCleoI
NMUsm/X1UMi2G6KWARJtMiVI7aGjMp34KHOtiAf4rlha+OA6I5JZL7IImY9TLejI
NbI946aJc0GRhbYADYh5iCQo6OxweRvYwayi0WEvSzLn6qzkA6fCIIGqNyASMRHO
ZCCoqrOGF/NKOW3zgbZ5rXTRSGDlMH2BNTFdGs4jfdhYVvzUqXe9cumY7z+LJniX
2A2yN2OhipdB/dVApaTMdGRVVjog759efLL8y07sLL138r/2TWVHjmIWcbkYIztH
MkFAkyJTsggoDpoerHt/abPtXszAAkai9kfvFIYxKi5eODdM80f/ScDBaDxpNRgb
mBmIZJh6rBj+pvEEyK+UIwB1/k+vYJEy0GAQavUvKNh3WgCfY1X8wSGf02Gqr/IB
zvHWnh/xgXQxEC9rBj8hROvCyHkKc3Ebzjq7M6A0KI/TXeMfUcKYE1BZJjjnd9Y9
iFUNGaoT6IKVfAZuFq3x8Mpk+pXuYhdBEavThKnWmXxTr2OVorg3skzPY7jiWcqO
PIEyYiBHH9Zl3nT31s3YkwYPCGRGXMsD+dcV+T3wzBI7N/mAHRyY5pq2scNxXvsK
lnCmv/2nZgAdSC0hLJtCvVbdyrWqRDrXdu+dU9AKJxhchLEwM6yknzPDEMvhi4yc
tgFLwerrdWawj/3QHWG+ygU4VD/GrnWdo+g/UkopJpqAGK7MnB1my4ksXNE2ZsOH
llNnMHJIc+DH5MrFOZoqOpef4+c9dD7jX1M4PgSdVhKcXUl8+zjViNCisMdaBGcg
fxvU7F5i8q4fK6LQgrV+Wee2fBf251nkcUPWCiR/ujv2B37DG/s+ZbuSeoDAE21/
oYn3w3VvFJZsoAFWL9vTy9dZJkJe4L1nCVGXBC3ZdUKwUgrN7cmGejLerBwvUBj0
uaFDtCPCLR0/BgygQmKckSVEvTvQ+T0014M90EjBFOaR/OZV8DS2ms2N2HDfQCds
cIuNf694OXJlRnrUJ1RHV+i05pQvRUmSQvd2tzse4Dy/+tbIPBw6rhvK1jH+aEvy
S9Iz5GziZHWgyZ+sii6vd2q0H/k8oIyKroj0yhaAFUPu9W/wO54ORrsqVlDZ5qaw
kG88oKFcHrD+SCIkEGSMyA0h8rhxN78iFWGtktpgSuS9pfegN3nSGAeGdmV2yNR+
NiGMi++8VaSsk+j5AQ5eSGeKs6+iPy/7mdvtjw9ma80U7VGbiCG5bGd6Znwwrxfm
GSVeazx39vu/toSGYraZ/2DSHtvzOycGAPj5+SnztjKhKEAnp8AY+xaiZ/rKVjyp
7tjey5QMEAEdGsI4mYVNAHrMUfSvqhgVEnKcukBuB8G+zvl8xJxKJjUulUHB2D5j
BXwvglOPuVinqmT5H8DO++INOj1P7GGt3FcjYCtJwEAjE7w/dihZUOmlEjfPMwuX
Sby8VW3ZADe4UIdsfKb7/iyXz64B/a9QpflzgrY8h5enhOQhchaGrGuepI7oUjAj
18hyKrBTZNEF+04JTl7NrH0cCYopmGU2Z5fHfnZ74fNgKgaU2sn3FH4sW3pOwiCq
Bpj/n3VyX2YCYQm3bv2VxE3ml9GyJqWn1uPbrJQz7kBfD7eqTJNMacG9cAqwDzTJ
pHF6EQKV66kdvFBV2q6zCDz+A22cacPpBl4Lqp/tn7ZPtq61Jv0S+CLQXHLxKilZ
R07IbkOcJbA/CX6z/K35xGEcuS/OPJHX2OZxUbzwDs84MywZnWi0dCbUkVtFibAp
y7qfY/xeDbvnISvDJPUGn2RkcXjGcOYi+zm81Vd1Kirm4O5zjF4uQg0+E6JFijXm
xY6BgCdRAq1qubu7ZPVg3JpTQPq07gkvnUlIKJ9YqmNY6BcxZ0PQXtHcgxrQisg8
ZQJJd9cuZ0sGhnQWw8MgYXKDizu4V5ViPu3V/MaXA4WRniX4RvM4ZQ/bOx1I1bNj
AVbhhVSMZhaYDTK1nqVTIABXZ+zjOSuDZYjcHyX9v0F32ZHx412fLqV+NIc8Gwd0
jnF4mKLA4veyUkagEsljx0HyB08sDAgbdcqCdv3MgoyajbM4l2LWF5GRefudPkf3
wuOARamB5GPJKu5hfw7LOGp+yJdB4cfTs47/AANG2nE1GEPSbalTfTmgXlAQ8V6D
KDYBHd9qKxxl7P6WnkJZlzs0DL2Ko4fW6aTuEcKPwkjszJcVgaNK/koH+5O8v6cD
qMu6za5Y84JkP2oqmfI9lPVjYw4R1cvJ2v2BtJ/aHd2nuhWTTdz75QU178YJzPNH
ly8PYQviSfvA9uMyHXA6vqGk/r3FAoRU0zPHFxe+du+cJzDGiH8Uv/wDh61NwF7H
1tksXnT39/CxZljgwMLPh11O2U1RGgbzmoKZshBzi3Yn8Aa74c2HFHMLeSO0zz7w
KmtW0A983r7bv9T7ni8mwd/CT0y1NvxVOzleyRd4QNIF6OzOIdDUDdmmm5Vcbn/n
tfUvchRA+0cTDgiJQDZTsxeNP5zITAinXHdQ34mibQWfi69sBeHOl81W7mfYfIib
T6vdDZJDL9+noFsCGIGmPhQdL685O7kdepLYyiOgEs/dUqfwW4f5Y9R22+3kw6G3
sVCR6nZ5OD2j+v92Zujfd/CG5f8TbJlZy/q0X4XZ6Yg6TNgNvIM5Ai4B3L33rgcc
cKuK9gY56Z2QJJ9frmOiHy4QMWiWq+4OOU+fIifm9UriTFccrfAhvQPVzd5oSvxT
qca7+6fYyTwolH74cJ975WJQNKZiohp2dBYOWe5cZU8kH97BP1oq6do+prGlYlL6
gNstQBLUwaGVfTiTlaOvf+mhaNV4t3fMi38u+QIclV2ymvC1vCc97duAO0o9baxr
HXtaYRmbq1ctJQV5sz7xmEseyZfQ3F864QkLztFqwn73xI/kwhkMQYHPsPH+jhZN
RpX9IRqk+6VpqQqkPVn11AQE6so1R4Kz/5xiH59Df1F9AZNtTKM4BuB4eIFJYLvV
OVaLCSfG9xP2x6x4do50DKbZpVjO2U4wbvjKuHJCN6uD2vHX5SLow1rP89eK54jp
4JUWT/2JBSQqQKn0ZarWGqHOg8Xm6s3KrnPqFS0ybtpEOA8uvSHg4ekV5Nk30brC
6s+QRMCSWWH+4X862goNH6Omhc4j3AqA8Q6Ditvz1vjY408ywBDWCh2TghngXv40
oKxGpfQ19LmtbYEd7VDnc2R9e1NdK6OrsCHqFDOInFh1U+KAwsA+9GIE9vIpWxSG
ZkuqvxwEiKMU2QaLhn15ujx11GxvFVJAiHnLob3uBfjfEbotX4Lp1BmtxPU72fLh
/zAsoQ7RuBLFnfMIxjiUuFzE9kHkYDGFhlkSlc9aJ6jWxmJ566+lB/xvg+ifVrOA
otDpHUItReVQRtkcrL2u2uFzkXaJrCtCXdbBsQbLPuUdH+fTFUHpOgGlSKI+hxQG
zrK37pkuAXpkG/SIiSws7EQtdGxzDS4GjKYgo3Zq8msMWoutu86vVCj0njsjVs3M
dAsoiCMvvYjWXQHRkjDDlXeu/CBBMtlHkKWsEJHGM4Tg+zA4LPrploDa/+Fo5Vii
2g+hWlw2dkmganPD379dLORoJuK6Pr+cMQrWd8zDnqrCOKhFFxYh8tUi/tsHlnLK
n0bZ8zC384ymDrP3ueIdcAZvHfgdnV4u/y/JQeroUnL1F7jNk5dzYVxhy0v4tGGs
NSGm7tfoP6R6Kqum+F2JLw4rXPnoRpFhBTdLsnVljblpZvvhZpp7HLxuwRA8LsC/
R4qkT9ch5/VxDyoPlHMQDtA0IVJINdH/b4pM7PkHzXMBcP46zg38PtRip8LOP+H4
FRZm0Z5xlI7h6bPvPh63FmZfXV6P3ARW1ie1edBwUfn+9fGBJ4EOnK3iaHrk892L
bOShqGJPJFnE9TTcTm1/wJ9BYp8LEQSBse2Q8n4xokq4sBiNWKjelnFq6PBQkmCI
qSRO+RHj1THtZ6X7jW3jd7VALdJqna+ZAaQ6UgHnYJR/5OLoDynSGZBN/fH/akL3
dzdi0arEtc6E4QWXgaqHvBHUqQ8TuCeD4z1sftyRA0pgrKxCRO5PqFWVqYLr8JX+
CwBKI+F3ECb+/qkUS4xd5AKkdT124azAE4GHcM8b51Q8qBAujauZqqonQACScfvW
ozc8DkqL91x6ZyL9za6JXt7xh6osAZsrgDrHFQ3Vowfdt8uVa+VcdDg/4uNLmthk
eYPBjPYIEhsHjONCS/5C5AIRMxa0OkxgB2ANSp6wSFE/BgmRhPmmA2zt71v5VY6X
3e58whW10QEMl6Ezk5fkcp6sdGK58Sg+lbeFt9n7ME9V5HcbZnhEV0pvULS4lw4k
iRX+3Kjk9Q1wu3Uxb/1fRko1iJ2oDZ49kEjZw1kBJYJ+/ccScXiv7MEebKbjHP11
qPX88lIP07ToruAqCrQIrWmll9GYFHfsb8U+kTUELJFdEBkb6Ua8wVHgOwGvIirJ
mFE1SytIIahAIgW8dh5lnGZoUKyj1Nqo84m1CIagfBNRakMhl2orh7h/D+48d0FK
M/UDXrFrrZAFxggkxCVcrZ23S+raFuwTdWmugcCnoXHWtuGIX6eRCzKUEbEcYaQe
6mZk++3y+9xpkZpwfpQGRsQEc3ZPb1cilIdHfSy9QigyYOq5LQnqFI3gyMy1ZE87
b/sPlw34Q56PfsX77cYXYrPdA4z9E9MW/cWtZQd8nxDcin53XFDoiUntbek+TWew
TphktB1v8Oe9tyFLleJiLAa3Uu01y/4nKRahCM9T9RJdkePtdd3urvIG2zMVapjx
oy0zZpOVgIOxMt4yn1oiCkkzO1KL5PF6mHIhke8CV+fy+7I5l2+Na7eqG0Y4g1WJ
DyBy5KU34S/NkCFuh1kLqdSxtDg9lJD0J60ctAc/yS8uYKyoQooBpVzefdT6Aicu
bNkJO5rTwS1OCPJzorP2OjhJFupWmOzoTBzx5vtE94tHQ4DPLRGPdDB12DfCdL9U
a6L6DqkvZWDMMryy5uJOlh+5jDj3U20audYSpMiHC6hd/tOVS0tHmA27HtF68ZKW
MZ2PU/m1QEv4zDHiDFTtcn7UetX88bUG1sh5kLkyqPp4Rjv+3d1d4qRlD0RKpAj7
ZA33LKthRcJn4lEtL8pPF9sWH5zvfki8TmrvPCXSTJyo8vC0PXnVGcq1xCu7Ae9r
SnfRUkLdC0ryMmabIxAtrNrRpNInjfSNHukE02gjF3n/LKxbKx/4BlVpalTt+lYr
PVhqHvA3WM9nhhwWRCeJ/l13Bc4ylYB9K8m8KDK9ZFto8n/oRuEvV5L2wLYOYhYN
PnDQPGvD0fVrBoDtJvtZa4N9As283A9txsVEpHyqXgbi088QyhnEmnvJTztDKE4t
uQEllG9Rwkm2NEnDkNDv2EyQgC+WJWywpIc/MfixRYAZiC9rlwH9jPfuNc87e5Nh
yGNo1S4mlGi1zhn/ec+wv6CO0V7Sjrec2G8vKBVQNFkmzPsdet3Ch2w7zDCnYEPQ
mehzajj++eDbUS7KkxKJMIy748pMeWo3sz3r3Av1JWXrklI9O7pcX6Xm8qx5iX3v
kWgvFG3iOQ1q0TglMSugSRzsP7LNeMf2bCvp6IzKNGTT88JjgNM8Bd4t83rQNBLH
lEI/OHxngTjXc/AuztYv3SoMuesXg4rbzjQZYucNsyw3fTrsIZO5kI49WaVurgLF
7ZtcvABKDWSz6rM5+BGEz0vbI6XSD2GnkssaNZuIDDW5nvYK8AC3it9oBANleBZS
RxRl8jEfYpy6msm7cPqaaTMk/3VXwME6kV5HJYK9n6GlCOG44CfxJ96wyNB9DkgE
Kn0YwUQQtlgz5NStzxhwupqW4Xatgov9yZO1q0jL3nW6ZVBP9Svcx9iB7v5EfhyR
n0zO+b+WxIWNG4kEkWZFrBlgHg192PyFZQN1geEsEE8IbkhjCHuIHwxABQFTI9Gx
cqa4XjsWfacI85B+pEkcxSgEkW7/Aswgmr5bP1DiWwJqYEwnY6l8rfEGbTzoV+G6
nuSWGfRhvLckglIjOEKx7udBGUfRI/FXCz9eQyKdoLAxCaXq4HD3TJGyKRG0umYq
nJ9QHzmdJSCbUzcL+pxEByBSq2TZk7lw8H0+ZaS9JZ1Ry+BTOqiDqizIa+FreQu6
zoln/gg4nGZjMvPi1yW6FaQmAGLPwdo8E8DK662kEw35jsjv7/INbsss9x0nmiOM
l4NI0+hadOQ+ua9FlrNgphmZl1LzRVQNGN02B9OhkSH+GmJugRIlCkgIDFSq3VOc
pOX7DIvOo8pyHZ/su/RTJRcjadihTprOvYTDXr7I/q830V79YKpgWI85TLDi2szH
KIUx9L6mQv9axBRzHJ+iFAy8Gp6EJ2jkX28/QTLxbDx3CjOG9+48CHJ76Lf5o3dY
q4VD+rhi63PWa0w+khbAY/dzrHo/T8u0I09vx9XWrN5kNpOqbA4cu4kxbAFAVNQ8
dyld+ltIJFCnMK7RCKGbvtAuqaaSvAczzWbokimG+1JhTt29sI6r17foG2MJE+1/
Zkq23FHsJOQiOOl6mBbpRX2oejrX5vOCp/t7T+jQisKFuHBlJieoV2ZH3eKyBbzb
K54OsKK8PS7wocQh+4V3czmfyvMfNJ56JWNDtKzqjtLaGcclD4nFZdZ7nRy5ykyt
0Jh7paZwQCQe5cqUCnDWm6jTfhSVTSck6tR2qUGawGPXOvaPNZBomjh04r1SHHJ1
jzN/T5Prk4eegdI89KA0gwpCkMYmLgF/WMOdOFsNTU73HIVV7kG0AB59Aux84kzI
nXp61qB/Xk634fxTv8ucfWSpxM0o6x0WzgpH1+T03+UOB9b55bhWFCzR6UFeMFsM
pYyaIcZHuAOiRGEwybGMjt+Y91QwQh1d4J9EUdyu85XCbxkrAtAi3/ipwk7aZOr1
6lRI4ugSONKl4abc38RLHKFWvZ2ebdUuM2ZdFZG5NyRC3c4aZDgkjegI6jiAGV2c
BVXC8YsPwP+wMbSXYGaPcRcWbHpIbuC5b0dQVb/p5+B/8CmYTrdTmng+6YZpPARR
9EGvED9X9rQMPZug5VcAsNmVytG86DarHuoTFCpCZfPqE+qCKqmVlyGTEt2STFMh
Sx/Oh2m73jC9dTUPz2Kiv2lyoZvn+3tc7MKttNQVIMpGqsYyNxdLjJ5HEuODIw+3
oQGqMvmKzXbAYSFM8m6UEpmDbp0nHLxK33mGipuR3mQYSZAcwwpkQweRM45yPwjM
1GzEjXP9PpDUrtYxgKRv//F/fsfmF//hPMtq6slPfQcpSDYRAEorkYU0Y7BHPi25
0DBNe0piLD/Qg2O/ueeEEJ1pns7QJhcicObhLx9lG36oH7ZzQ4tF+W5QcXx/+/WN
o9z4ioIgInSkk4cE34u0/gQ3kWIIiGEwDadeYGZjavk3eCZX2MYsFr6HaR8Fo+28
ccAAJcUiJgFWE6fWtAijPoEEk5/VHf94eWIyLte7YD7lgTwVOcDrAgTK0PLir8c9
JE2d7NL4k2dZ3SpkUj06Y73YU42g7fbW/Lvt0rikkIPfI2g3LzBc5k/Ad5JRPoAQ
mFQFr8GcU1TbrPFRgYLfRBIPw0R/qXMC41ryjVsjtUrWpabJDs3P5MY7ba/VDrUe
DrMsA3DWG0kCBP8DRRoxW8y9DV+Jdo6kQjFkjaN8dWy1ChC3fEhBWsDackyJXXfI
DYOpw4vnU+wRzqM/82KB9XK/Fik63y9LY901lEfBbrgYPU7e71l+6dng3jNVI+RR
h5GJIHYYeMHPqOYqfuwk5pEwBrFDL6+SUifjBz0IfZOiZ6Qyry0J0Nf91izKVj1/
APsh6W2FPyqm0u8Ncfbp4Kn2De9lYR9cMLX/lRiTPhlw1KfEGWhGNk1ODOB+4twN
ijjZ+DpqdKdiI0yKVhhuwlAgZCybPZI93UvS5w8sLP5v/I8ciz6GLE1BGEE3lmCS
yIPWV9ywBiMzJSyCf04lVEkF+BPAlhcMJFzeGUDdEDi+xYaeJZTh3MFeFebTv4c0
8CVgN7qN7lUHz7IprEY4RgkgcMEx8B0oPFR4a8okgO2MOtnt9NT6KbJSeD6f83VC
l7ErYAws6Ri9CZla+WimrVatFEz6zrxOwKatoQsYZ9F6HEN+S5FfeOTEcmbd28Lg
FopRtrjWuEA88wlPqO2WP2/O4GKcOAS2xYedXKhiAcGshUi9ncBV4CXG27K3TxbN
vXmOG9yBQLvp14Ep9yFB3ddPpepguci4kXUQux67+8h8rl53ngKAe9tmhmNc/wTD
GeWSjsMnnC8p7hZPqMbtJpf4/TthUeu8qmTxao5XF6zOh2CqfADVRgMHpBwEuNit
1XGy+osAbvbo3WlvH3Db9hlu0JkuBCM/xPzV49IM10zF4g2v/+BazogKYtTExo0k
qM6Nt8tGqOGR+IlGIFG8RAng71Cnmh/7i44eg1a1bnpzQzHSR3ey6nhG1EZ6yY3h
R5b3n7wuS9FgoSaiPuqV5Jq5UcBzROWlE15FjYx8Yfkk48kb7solHAfLKrhnV6Pd
7f069rPjgkfNv640qv9HNIn60WonfUVGGmOuOKRx5AD6D5PXRDtzoPdnoOfHEJA+
IKU1DLrw7+8PqG9P6mtQVIuxK+IYv7zQJFZ5MwmaROqeHCL5SqgVW53vPfHEMiyD
iQB555r3EVXt5mz5wuKZ/DhSa3yBYv0u1S/BHTQi9Zb/nzz1oUXKkVRFXYVFTTJt
xXaiOmcilI2A1x//n4dMMXJSClKZ/s38UkZDRUP4cak82GWOLJfwDvPkxRMa++a4
NTaRmoJDSPO/U/YEMx60ZIZH/T4wu1LpXv1viykiF78f+hdS7DVczTVOeks6UVOB
5igg5fqfYpq6JIKp1yiMRxqNmgbTPO2HXiWTntchwAnL2WNiOwZLqzOK0Ja6U8Lh
PqkZrIgN/R37cwkG6VVAxqDH700xC+zHMkSOD0292+v5gmO57qEt0JnB2qCmQ0rj
PnHXfThkvCUoWKZZBoHfA1aZccc2s1YUu6njmk0xrYCnLxM50kj8qCM1JK37XhUu
PME58Hhr+kF3rDWiAl9wuvTn7ylpFQ+67zu+QzW8RJfyz2NAafFdiz5p5g3AEJeL
S1JqOvvALXX+370w3lwVnZU94adrvTpu2JFy1M08p2DeZuJxubOBbBqF2xICiYAa
2+ocvjJB3Fad/1FTutMQqr08eQJG9jrdPYyHu29CMhefSOCW95ik0Z7AQLVdbKA/
7jHMm5zC7wtYmzFl2fj90hmJYFBrbQuAJYD46Os5GRZzrCQdDBEEDPg7uni+x4Pb
aA/pvyo9Uo83GJ0NJsCsmCgE5J5RQKu7FB264OiKo9e2D3lLXckt9dLpQoru+F/o
gHoF5msCT08hkcWwZO3jm+fhdWTBoMr2h0HIAsjQ6T8CGg0MNSCr27jiCKKRWJqi
KSIG8HxZJ17u/5u0hycxhk5udgp1ke+WoaFZ5J25AMQ7o89O11kEaXEpTafS7LhP
wti0In7tmpGWJZY4L82gSZODPhCbZy8dxMdsvCqpw/WAsDa2R697v8U3uVBjSzlr
spdUS/Pvg8J4UWylG8CJa52YSZZ7w4d5RDxYw/rJFV5e0Z3xDFgo8HeEDg7rlDcs
JBJtMoImZZy00Mg6ir4HMmuWD551/GUcLwjzMagsuQXXZ4uWaqQZA9Y8umWb/G5j
J3coi7YNbMUg/Qu6kg+SFms/U3fpefj/0k6mydwpLvI+sLl6TPhPIF2kVZcR0CCT
pvPyDcxL+TQep05PCX4cx0NFKwED6GNHibOtjiaqZ9N/J2RPdN1dif4mIFH+PDTA
pEU9me7htySGzvrId2KRaUfi4xQpxdAUSe1zkXG3FjPUhwglDpSZboAhYGfsr5tv
ns58h2XWIDYFSyyjU+10DHj56K5H+BSVIkLC7aTrNWt0iPMEwoRB4Ps2N+G6zN/7
BWYrGoifAhdoEbiTyZEsJbz2IPplIjWhCBxGyghq+GYShwSyV0VMxLoY6fskU3rx
fgBZWg1KEWXX77+XhnglSMO/mtjKPw+ODcXTC9t5ye2Vsh+GPyKM1R9tmFWR+XYF
nHP0wz6C1ypxMuF3zt+rZnH/tJfv6KvEGnqR1HPIYgwJuY5vSXtevx5IhQwZCbd/
qgAato8y2WR5bYF3ieYZCPHve5SDu3PNDT5F5zVfeEvGkXfY7cu5Vibk+UjWP4Qf
sp++bfzRRSsWs6NQx2p7mqgkIItBexBkoiMCdy9iBCGgxdk8tHMDj1kyII7HlB0O
5RSl1geNCEYytic6Bbz3kAjgg2wIYDdX2ZDjOmaZ5vJ0r5vE+DX+KLsZlFph4rAb
kCoe269zmJossfwKNkKBxNnOpj+J6/VjPiZQ6ZW7GtxL5MO0WeuK0rQcC81cVWZ5
NV4U74Rd6FDxJsgWEBVYKp3w3XijkjKWkG8KDCz0igar5+Uo2lNKefPADXw8Jwqv
F9O9447ezqvRD/D9OTn/gTqaZEqvmRxUhsCq3AGAjLQSMQZewSEN9ivjYtPjh5Xu
k4wHbwXnWSChkXoDVuLJV8BjJ1fvOsyG6sn3AJnE7aNbLUVK5Vqgqy6PJX4nw+Rr
MfSdgMgJF0EB7QFFGFQ191/H0STVan88kNYUiG1dgPeQq7HT5/ta5fSfcu/Td1x5
7VfrmDorrHVC30oSb0k7zOa4af9slhKAS4OASfQtfBF2+iUoVEVG4RBKikOzyf6w
a7nuC2u5QvCUEDT9D0rhtSvNk8rHZ7v8RMaOJVSzUW8krL1e5vVenMPKagPAA2Rn
vP13XiJcBfshdVUCAZSlEJrWHnR7oKeN8FP8/dtdZvQ4J3zyIVqQILBo27VLQGV/
JBgOuSUADrEWn5rUshvtfy7qhJQIYEs4z9kckI0tloU6WKSy22+KLDZoRxByc9wm
vWksrp/n1DnPh4dgMg3XfORBxte7u7B5ZflIspRVEvnXfELdawHSQmgw3uv70aLm
b3VcRMRhbb957lzuAhSd3ixRly1ktEwt3IehljoJc55s9IGmhrzcrZXBCFqP5JnP
Yg75JddMMX+iD6HbplkkJUTgvSjK0LNw8VKdJpjC+Va6Ox35CwxJGfLLlo2cAGN2
gII4bJOCC1k7MjBrHEbdoSO2AE3gJtS9geqCZOTqNIspU5DOqqRQMpf+snTGZm7P
cGTQVTNtElR8iqUqqoxAz5GTKAngRRiOxQA/47dpO3LPiRvwuWzQuSIuIg40quPx
gbVJPnVMSyPZU/cwi+20QHTwg3dgMj1k+O/2ECqVP/mhipWwadKawv+RY/u6IJ84
C+WX29DkRE7gotabqFpX+Yj1m18+gQbsh7TdvZcG6jN3gsljY2E5w7Mi5FhKzUmY
jhWBJatp3+Zn0yXA6SgI/2vRwAalEwfxF2imZbPfdrg6J90gVgHVEFbVBF/9y/yG
kuNZm8YfIJnR957/NdN5NI3dDRM8ubP69EWAcSasb2Ctkk5OhgrihXqmAodiageo
xsN724Pziq3Js6TDBbdBqhf4sJvwEfNqt92kS1VEED6QeblnY/KOszCLxq9bj90a
+5ro1e13skyoNvLIsofbE22gS7pDT+jBDP+AV8bDEgMThQ/oSJlO5clTo7s4fQiJ
uHh70XExBLTtxtePOzQfPVIYirkzjf1e4OhGIK90Z87AACrp/5Og+QLsK8UhHDPZ
io7uIsY3x48ATIlWRziQlhppGX5QF/3mGFcCMLXJJXpavWc8alhR07Ruf3ExCnh7
/FvlLS1YgVscB8yHApLXvA8AcA8K/he6dIPP/G0BJHeNwZumd8VBLTUWXzMywz2t
4RgY/RY9ZXlrNBIgC1eGZaNAyZULnaCQQzvRFSRqaelWpwAjaSBKjFivzw5FJxQv
HVBcfzKiC2lpyZpRZm9UI8FwoeuMCkZ4MNHoUwEEt/NhfAlse36Wy0OI48HO5CRo
im7myjTHTQBVx2o7fArLV3/Mr3PrOBq+0iSe4yN3pTpR3730jmLTOKkH6bflRT4U
+FHU7mAMgbAVe/pPbyn43vJA6PkJ60b78Rxh/ws1S32cWra3920SWlK9C3MXAGVe
VZgAGyRaj+F0+YCT4jehj991cV2W7PI/8IfT5tTHd70yOO6PIyWIzsM5LFqKJg5T
WFpRVRXFCyY1yTFhTBue9mimAK/2hgORQ+hnABare2ctiRysDc593y3MHDvT+ojX
ri3Fmqb0mNzHgidQp3N0SnNJFVvopT+gMWPd8E+y5WwKCldIqk/wOiG0TM790omw
3oUAmKnEVyXKnb1IZizx44HvmTrrIeev2t1PJ1IQFf/EZxbSE9QMOKdhUL0qbLO7
zyyjFqzyV9yCcifwKEw+X+zXMirRKFhLRAqAp6h0OJqL+msyMpGDmvjha4DwHb/I
GnHGhzTx3pW2pkXapSr06DEI1K4FauKHTpRs/u9MHXl9BVDUgsaoMh1XrdUwV4Ut
kfCC/AD9dd/Flakwuz0OjgZ50aAgCVHut0vylYXq9NCnRP5VsSNAmcxNLdu4gPU9
SBjOfT/KSAFK6vPJvujewP0qvDdoQkXnlc+XILn62WCPLeONkbMrkUtIaspiQQ1Z
0LvE2Z9UfZgXItCTgpP0u+aAAf0ofb+TFnTwdxu9uLw7EOg6DUM60aeT9izhZmbM
7jahyloQBSn03mn5QBcNUQNgaWPUWKsyBAx0LVspVMeyvZY8xvCfUwt7g5UWChI0
VIIJmQyMwEI9sjE0mam3wcLVh0kKy61gOY+jaronjX1Wc609FTsUFekrj4kYtKCl
E9rIS7U0WhjpyLLJzlp1Z+BIENYERY2VdngJDDCewqLJ+CtZrYRT2Fy3RggHzOqt
0cGTza16lrHinTFYZ3dCc1r6eijClTOMvyZZDxb1q9kWZXopumBpMQp3X7xSlYi5
AV7ARnEdz1BE2ohkt6bHmoxCStu/BOsc973mRLHo8sTT+hFWy9yaJjXUwdoC9veR
y9lH4TxpZNsN14sWRmaLk3BqnltbyHFqiv5c49vVH6rIN9EtXSDdIIJS65LumuF2
1tZESHd4pr3nTuyMVU0w7UA3Ut7t30rVLXUkqwGsK2GQPp37zEl8I4Vv1g9sv5B+
fEs2hlvQtbyItjJNQUHzJ34iVFsDKzg6QiSw8H56BlQ68yHT7NbEfP2lct/HOnJw
whilQDBAlIuum/l7nO8yi9CHPICBaQ3OpHYkJzG2kVbGB3yWcwwkyOp9ygSOblFQ
HG5Owvlgfeeus4dOvkcZ+7964NWx+10pNHcyzKH33x3SsY5IHdw7O4qdwbR+/1cw
EilMPehxxAQ3vIdcFXfd+7El1EJZlugsLkJFE8QpLDGEEeyoGTncbm0mSiJU1KRv
GHR3dhIWBO/lymyF1WOvj4Z0e1aS4Zagp4Jqcd2SxWebkByeZ5EHK1k3vd+K8k7S
JY+2kWQZF101cHT5HnTImcPHoYMHzGsnwERg7kJifLT+x0OSAtOdMyXMsInL5LRH
qtRBJQslkcVDwQbo2G5UBm6lX19bhIYYdc//rhBoo/85vy3BrGy/t+MXYkItm1ho
rcZulRoi2W6KyDUkTe1vmEWUaBqxjFbrtELUpY+i1zCntJJbTgBR/LfICgmYw8Ws
XLTOKLV9BARpmA5SJQe6HmpI3Y786os4gObot58pGrOQiN2tMRLoBNK2eNWwaCsE
0BwzeQi7/RpFudGzH5lDKUvKRbv7voUHQi9W93bCP8Y2EtD73LSIul9h1zvLaTZm
cY5441v4hoJYuGOUBxr44mENwGdX7LKrelgNXZuycBGyeQ8AIkX5DB8sXhFQHDWx
oYO6kp3bnWlCuBq34ALUUgydbe36x1p5vTK30LTdMmdoSctKgwvwhf35LhszqRK+
0/7Tb1CLCZE2rpnaf6+H74rhUhB2wIhovcj40+u0wqRNTfS/f6QXzUdcSMhtqoxf
tPAyrAaoARUrkauODYumkJfspIh97RIdCqy1+aF5IyUDYuTJBq0L6fLQXby9NtmJ
rTNAR1u6kIkLeUVOaamWh4JpVrMx8KIPgZygSlf8U8QpIKnY9d97ZufWud/82cp9
i1irDydkl8w+OGCGa1pL40wxFJ3yHgXzy80W/77mrXRr44GRTtcLpD9NQgGaGmp7
1amY3FKMIsmTghd53A2WpLRpx5VtoHIJsBlBeodbhiTCwMvbEsyVBUKoca8N9cjL
rM+qWxXAFHD0O0fMYJ1cmHUeihcqyccylthkRyXy8+PPyg7mJnBkV6VObX5yXFem
F3lN+I3n57n7nNqYOaag7PZJImIiJ41SsfyTGC0Up5eV0ikMXFcj78yXYlauI0oM
yjgePkpux+3rqP8H8bN71kSej2MifgjXA1HOUKoCXGNnxkLUj1keCmAUj0vl2OC5
2swgGKN06uUB1FOmqgz8rvxpoS7nMgoVhLzu/KkBKO2wz7icMuGxdrg0Jf3OGQYZ
3clQ5I/6UgZ8NxjgJffzxyhI+UVIm6KBYx+ATkeUlAlZ1T+9cCRgKTUaxkvwNzyj
C+e6ypD22NFR2ghHr+nBj0hRzG4P36mPqjWQ/Ucina+Y2kC/vi3G1AgDOSnfblGu
JB2cmK9g9OovnskDfj0F0vwKfiu1fXvZEw3Q1SJ03abgecl15NQXoOdDp/XIw1HV
Urm7wom7RLh+rWvy23lARG0fVKouSOZZlnQjfyc+DyVrUFXhTGGjiRy5yvldrUwB
d4Kc6yz34WmIFsbmFakE8yce0L+Y8xSsfLzIHk+LdEGjZ3taIDYgchCOlJwuBDQZ
xenxSGgj6mKagdQzzUH0hAOMds9++j3wPphNhUtn2sDnG1kSsBf02WxwzEafg97B
YyOml4MPnyK++AxYksQW7dNUb0058OUsl7ZzIRxXCQubZ7ptshHbSDisEe7za6rH
tbf2WW16R7fgA8BUoCv/LqXEytPhSuYfsw3oEOu6cAf/h017BW9d7tsfMl1pDkbR
Wy36MOO6+SkGO9Ni+KyfqbcahdEtfHRWJFqhOAGvLgcXbqZhDnzTXXxOmNCv0SYS
SPObaoGJL5lNdYz0LKo4Ao4VSsfL9QTvYOAbPhLAndX61AryUUZq8kMb55bzucjk
GLWdxu9PSN84PgDGv3kxH6/KMiTWjWEGufW4BMPSlqoc1hwGvlVhGgs0sftArcLU
+u/xyCUHB0Nb7L/nt8wvf5RY05Ntcjw4Yi+XDB2l0Sz6zg0ff40wK2K/DZplYXTx
Zeerpxo3tzW8GB0P4LwfTEj3zel4/c8ru0xnqGxp3LIF6sxBgMmLrvskCg8be2Z+
IweaOmebc+IylAf3a5yMqxyLZMAEn8hpWNWH7LvRYK5oCETEHCVWo6ldX23XSWuX
NfEyjBDW3c7TVKmI5tzi8fc4y0z0UFG5ilMjHdtRAnhIDEkdrwBxyGuhOdOkH/d/
StAHZqPbSeHrPFiuZn1QHsCdHrMutvseofhY1j75XEc5fEptxw9ak27yPRcldnvz
dkZdJneKiZKh/RNBO9x/034VnJepF4LzX5HmlSZ/zCce2xh1YursFtL0AFJrNdEl
X2C4M53wJ0eIcABQKGKMYa/I1lTRLNH9O34VJkykg4KFSvvEfre8qgKzVUncuxRN
Ce/Tci5KHXKm7HewePWSX73tdJGMdrAwq+kMKrZC/9cTAUiUZvt5T3PD3yk6gbzA
Tgw+vAmgTbXomrV/IauvUwnLdWR5+KZQnblWjpemwh4j7gHgARFhlVdGWTwrm2IW
8zLtFJdMnMpZbF+8VlIiUvnjBRpuJRQgydPqaC86bkwZWcwt0NqsHMiJDJkZ7HL4
1KSL/O8dBjBWtON+93XxYR6JDUL9TMg+tNTVarVYv+WJfMqnSwrc+lL57G6DhLm6
+yIyLAlg+yHyK0TrCGO3cmkNm8TKRBAqI229AiWpCrlmD49b/zzlGQ1TwVLtOJiG
XTF2AhlqrbxDuni63YySUNxNNbWMnCH7egqtsYFoxlnWqU464vXSAeRPx/b+j9u5
iKoOfrN/4LDiVaKgjfOnKSCBTdWdDscNnt9bCz0Lu6tdx2nLZ+HNagVUZpYjcFqY
anSQ+95/z5RCWV/mTomJgxQrOImsqWXV6eBYQ3ufP7DWCuA1JYWu64mGdzxtcCL1
LQRc/CpiPZ9dxrg+O/rUpmh9/O2IuACg5RAGNUZMNc2tYtx1cbq3OXXG8wDS4vk9
NTfOINow5NKbNL5G58o+5itBAJyqYv2etV3JTWo+UspSrbQe3y19Yq7HzT/nIIzb
QWB3A/SLr+Zftr38nlbaEPrqUPvy3rgoDOHu539xkPyZ3MN/emgYKvdOzw9ccqWs
8du0qxoIkRSDVLZKS0ljcAB1H5toAzM8xbwb/JEzF43HIptRIRb2SYp2jjmYcYa8
bUHat+OQefqE63wnAh5h++4QUpBQoq+wSPQWIxwQIeHrOfNKlOIZ1NkYqF4H4fM8
SkjwLin2oARHZr2Cyz8FOgyrDmeOd6v4Z2eg7ZiA7ctR1J2Pp8Z0/M2WhqL3l+JW
GwU2wFIeqtQ6ZzpwFy6xVVAky5Enk9qnP8ret2XCieEConNp/UPyCac08rWFpp55
1LipMblR00FGtrqSsrhCZq4INbMNcfuHMpDI8jXs6URxML/eFtQ3r9xp/6DJrvft
hIIphUqzYlFhiIoA9cnBLhqPun+B6T8BnLkWDtA/oAL6B5n5mD9Exe66u+JLuEUv
m3JfcXIap1tRG9RINA5OGtJ+Me0EG6+vATdmyEynZNu8zSGIjbIPxDpP2wgEU7Pz
5N58kCHui+ShYoL2S3rPd2Fo6ogFDYOGXN+zl1Iudx8aiVGlhVQUANhaoZG9gmfy
oa/0kAVnA+SS8ipXN8iM8NLyIK3uubPjja9cqY9iy12FcMouPEEDnaKdNrNzHUmL
DoGJ5KTXRUO42KJtIRKfQn3qqXEGTvcTcJPIoABKzo6SMPKzT+iHV2r0OH2CQ2Z2
uNBFpx1etHnc4qeKSG3/HOE5EXiS2fAR1x7aDBUWpOwi5JvqKqyAQjBYcACjXPbV
JlQ+LhS7TsEUZCkiuMBJovxVvwWraTz97NND6gbY0b4vF7lbMc12Y3hQ8WA7F4Z8
THGxSFGCTwnBdCqyIZEYLPTg5c5AzbjG+0S0P+0SGAFuc8gLY5sNFI/UIr7fqfrH
32FGfVEHa4XpmKWAa682t6CLLVUOB7z2b0gPfGiqSv+CZoJFXPwndetnlxhUaYc9
6WyvWgKSy/tksv0N+uK7NnFbw1GH66ufSaSx75IYaS5oG3Hd3gBs5fqmHPUCO+Sw
vJZuncreGPidjN+uS8EPTKJTaf1iquizR5QCbtj1zUdd1O02pgy76TazUBsWkwTb
2Zg9FMBFb7aI3bxcy5iYPbHDBPGXPuL9gTSxJgITti24IQtnz82YhEzs9l6kF3KB
bA+iIWQAi5G/2uhcL47Epj1PUO4J0hVjlQ1ryHfZ9Sn362mNNXfh7rmFjZSxuM6U
Lt8AGYy8buRiYgt61LlLuiXpGxMJbQrDHp3tiJkYsOj5179VgMC9Ter/ZIRLqYrA
JmOJPbUgcVipKiFGwt2ellRB1pkpwsbifXCZ6JfyBg706zibVux+shZaYb2WTIUo
kCKa4WloTLB8PHB30aXaz+nWAy5xZtAM2kF7tiKy2f1p2kWGBKvgRAE6PKyteVu0
MYDrwRG1AiM8SeM8/6BEZsYrYptQ9wpHd1H+R9BxBVJNVBoR4xXbT0cbaCeWNay+
NqvAKZhIJHuovh/bL3vA7TxXhfAX1Haj2ELD0O93D/IyTWZ54i7pRwsJ2xbzKz6h
uyY3w0Vma7ynP9wvoXgmT4+b/QnmEmlsg9/DcQmhcP2KBf+J7Ne80m1sTX3oH+RR
TfAt58J+c+8PHXw2uMM/O2gbX1ChPDdAUbcSJP10yK8pjAInZat5rHDc/3kDTjWW
d2B7f8ZuWDGJto0UGvT8CVfwpN8ouSxaAliEwsDhTH3sFkOTsfJRSCK7Ejbt1vwW
5lfluQei5VF7nothlBkPtUiF4jd8ltPYnd+hPjmAcxAioIp22BhL7dFDbugSPsR7
sgAdXs8YLwUZU5/1FLS2e7z5aHMZ3CWpI4uPpRai2w0wR59TlQjv0SEqjqH/nw2O
JcWfD2Qsg5Ycah4c3Ex9PsLIDhg6jKU/sCOstxpfgWeqk4mczERQQAemF/gcakI0
Usarhd3gz2D+3SaEIHbMSja7gQ51u326EpQBWHpl1NXiGfG5YvLBlIGAX3Jc0ea6
pBgf59kPXH3XiWMRU70EKUhq5SkFyborduQkgE7xiSlAluqzZDMur6j3BfcqIyIb
5gA5OeCxDAqbKpS2q2Dp5EtsSsgqs+G324b2AxbsL71SrDA8vvPpHNn3vJMpSwoU
09PtBWU1um+I1kDYXx43U6QiJuTHYqjoVzmKaivQ5rcSYr5XRxPDxdgBNknHqtJb
mezpGjhyX0gwznzBsrxUWigcXaAialsdaO2wM6ZI+Y/U/b3llQxIpowSumVaxioK
2oEWuoQlOodmyA+UybdzX5mvYXCBXHzChZuHYYQRkutl1AiwcWJJk9v3ArGeOljF
EluVRN+bJDtMAM7MBwZCvaThwaSyFtkFAyU054yz6cAIQIQZ2ITCYiZ/iaiv+LwX
8JnoDMQbKUQz0AGpXYlmJa8bXS7g7o4ISZ19JEKzLlvpMDsR+Y8Oj4hXYknAnnK5
JanR69rn5LYQKpniX9wiwO7feoPwcbQgaOE1EPe3ypwDgF+peYTYrL8vjAaMFp5k
O88jb++GmKXGwlLi9w2ltDC7LW9V5paSiQJE711Kh3m6iq8JHVPK697DkKpmvh5m
TrexHJmIdwF7ifkyD4YB52w9oKcqfGnTvVa3tU315axHiULXSyTs0IdZXfFLXs1U
5/xNnnH/Sy5KZ7NZ7QKD0FhafS1lykRcWmEaUZy0BpAv4Ys9J0HV2PyPJB0QO8CT
58QUEnEZef9n7oORC9cl8+rE8S3dzYk3N00PjZzTrFGcqLLXhGX/KhEi3Gw1EqTO
ZH4OZF+SZkTr8Ek3/zK/Hqk5zPe5Y3QUc3FCCj/WuYgIBTgVscAWTzsFYP1UPFn+
PI8gwad9R/fdUKFlMIYuZHD/5lvkLmjA2kmlamifyVoSKAtqLQAbBC0HN9kCQ6Y4
QA8W0ShafF/4hiw1WeYuun4dTRIU0HuyxYwwF+51NYhXiHdoN5/8cQTXS4lurdwJ
hYnOBRyO9HPDKGzMahvTZteagLLozU9slyF3/ktWbhNtwMybCsa8o2MLFyjuESZ8
WuaeJQrX70qhMbyKFGed2uZToSzecnI8EAxkmhd/GtBGY1nNyLZWzG5GBOAxGqmL
lMm6RbaaYgjkh3kxh9Mr0SrO0LkKfZU2dWTsADoctAiKd1SUaU7cIGPaVHRBnqLu
6ErghLu1CxXSsZ/wo7LhMGr7DsQ+HT8/pUU/gkGO4pTuleJwxFoOWv9nVibBbhB0
kYP208F6eD7ehFosZA4+mtd+skwlEWilFjKK9xzvI5h9+ucG2k875lTU/gPCI++2
LhC/8oJvX+PpVLf/zvBXBj8Bf1Xyq1QaDOojs52RFg9D08/NMsmX8oK+Grzc0/hY
7d0oUy/F1x4pRu9n8AiWO2cCpFkkKcdJKd+88BA6FXDcesxh2d8yh52pw13/flx2
6YS7eC+wAos9a8hep3vhe285Ys70iilhyGYPVY1Iewds9pqVEPe6X0M4Uyhv+tCM
M3YdSIZRqDTO8DGbwgbaP3hL4Gmky4eeuRpujlBgyzTV/vJrHjG4eisYfgT4XsJj
RbZJocOD7jf9YCf2/Z+e1ccwmA7v/RgctdjrhgblPklLqGPct72SjMmdqQy5AHmq
In53UY+3oAbF1Oe1JS91X1tc3WrS6FLLJ3IkzW3+o6uopkpRXMkVL5qbP/mAVkrY
wKOVv1hJY7288+aFvh/E4VfIi/723QV694jer8r+5NYZc/DMMi8icLn9/hRhbnZu
IrZJ0CvojAzntyXxp7D0J9r3tkqODV/2cj45Le5dISMAxqLuFeBql79qLQ8nahcf
E1L468SOiJweV9wPt6U668PbspfOcgic4f7LI48UtoxV8K0owx5KZrh9NpMdCFBU
NV++r3Cr/v5uk6PhYnY5DzX9adDxjqrE6LB2tWn0MqSthuM3ZZJzeo4tQrGkreaW
iKzuUuTHkxALg+w6sSmawiAPOr6LPCZB9W/80vlLKqbpwM++HrynWSZFkyLIWnmq
1VWwqqtf7dafMGXSCqD1QayH2EJxEysHNNw72UOdGNAJwX6839hDHVwjE1//dW9A
FqgaYUrtEzb2whieoR7ozfXPFsm9MH2hM3uv2en1RnRdIuX6pzEYRu6VJrIMoDPZ
axkbCrJpr/BysQRF+HG4fuF6rUd8MtC6+dnOtFPjmEEdGUAsZP297JnlHq5KSbwP
Xs4mTCvZEJLWqioqDDstU/QL/rOW9WdJs6CzP4RslYLOf1MF2TNU5W9bLk4UZaDg
M3An2uc/5zWM3Jee92FjlFs+IRSMK5zmUrbuPUNiRL4YV8UniWe+WR9SwuSUgZKe
YOMkmWUumCe4bX1flNODXlVeY/iHnjsc5ypIzmCCsdF0Wias8qruR5TsKUeLMWgR
sFBsbR6AWySHpYMQV3WZfK2bwrkZ4da8BNeMYgGJhDS7VfVoYDYrt0NUvl5oEAC1
pnOTgxLGOS3FGRQiZZeMeVLNOrL8CvGOq9ByLtcNjFhr+btTQjXC61bsQjRsyunY
rwaErRhNdnjzKHsHVKi0GNkWGFNQofrTKFD8VzNj1bouPiTeotaXEBhksB/qbjCe
I1okezhhnfcut11EWmsVI2kXc/SrHN0MN2hhsfBEo3DBUcJeInjTZlDFDB7QHrTi
6XoUgDi/OoIjLNJNEhukFDiP3eCSAKBaZfwxz7KCYHI+OorcCRdI/WXkR9Lw8sqs
Nte87LEyaweYmeBbvsym9ou2hqjF75X2a3ot66bsPw+g2XzDplhlvTyl8kws/7mV
FoTDBcZvsvquV+XjtJadQSpnzzbAF9IH66HakKF5lbR9c1FjDX72IDdgK5Lo/tb1
vIWUDYOOwze3+5k6oWxRNUHKJecfyyk+JhClDjUGAKEwbiju8u+t5FM2zDW43ZBa
UAZGf5qZIRMcuLj07VQ7mINo5tO+Zt7w9zGWIaOBlaF8vgDh4omfSjj/p38v8voc
MS63U1twuX5PVA+GmTlX5rLDuLCaRqjOPt/fOGpHjI26/HmClXOP/xs6VtcshryR
etnvKRfdXvVBpDFffLlJEaUZi7bqWtN6DPGh5B0v6o6kN1fY2MjOdibq0xB4QKUd
3058YxUc6/L6tNYTlhhvGzKTC3X27t0AQN1aVs4Bu08KpTko9tvukpuxF5r1koMS
qtoQzhJ6lVX0TyGYkOi/YdVRD8sdFVLZQWCUXrUz/VibcXutGcONdK/GNQUTqU1N
xOsCbT8FUVFzifO7wWBDpvigMsPYzmIvMLB8o8PXy+Rrk7NRdCIDHOC1dWYlSzYC
x5HBQqS2s9o8wt1yK/MDYgz87UqhHNzuX3DiJhvrmCB1b1Zp5SLOXL3GFlp5PzKF
s1CkaUuPQobv0eEi/GwT8tizUPnXoe2O7b/Py63+ZGQ9akNX9QS+Dsed56QSgOYs
SLCHBGln1ibabkEGvUdNdy/fNK9uBGU6lv37/gL8oLr4ZNLUG8Rom7XW2pTXQwF5
DAQP+t6rJcmesm4rNJb32iP/ZECjErL5B8WxlHVP2BBm9rosKwgt6HA171p59lQW
aArGDcokjWcVswfph/L3LB9137XJICYLk9NmCjezB/Q8Pip6OuqgKHxk26q8gYBc
bg0xHsV1+Klta+Lp+yNdikM/b5CrMoRSSfEox5QgHu1iPilGXXgrt5cQj41xydVa
ei6YN8It4xdr2Bi8dHtnIM2H+byU3h0xcobJnQdzdSGRELlazaMxABV07QYbmcKf
1xwU7qLsOo7UD1pYmk0qIikWfNJvrrv4mOYxGHQ3yUGTY3Tw8KrC2XucD2AEWSq3
gsoM4TDzRPitjFNK6ehoc4mEuQ/gmA63RxzzP/IujltDCU1l8JrG6ZhUAKolYyz0
5ym6kPQVNC6qgOduBzh7AWpX1w8xYkSmnxca987a5wysLJyy7f0WLVFlKkSMg038
GZLw2SN4VbW9oi2Fr/3JX6hkbU0i2Mf8Fb76F3TQaPVrPcBT6qVx3z7wzuQP3vYM
2yV+lPTBiaQkXOHhTN4uihNGtrULef6HJwtYI1d4WZBie/Lk21x+tdnVeIayhTGX
xP564B+o5DYjksQTunFI5VcKq28E0lxaAe7FkJKB+CLVnSTSsVFurKmIma9rTqUm
jBSwVJcQCnMcp35aUQHUzHRYw9CWSdYtrH0hWmfSYApOrEZIsuWlVYDvYVqPMmLO
BS1U37DTSjmN3C0bnWaHCBFQU+ZIfgMXGp7P5Z1P+z/QXsa/SCT5LyBsUorpu5O+
unX/MsV9bp5ASPOm8EugHMapSsBXzVxTuetpNnUTwkStbT2IJRUIZeInqfcx8E0P
G+x/NGPtMiAXZn7+wJqSMTtpE279YLC5QPo6ijKXHFr8ngSpVlSLnF+ybny2Mb4M
kY1zP9lw09KU4JlmEmpKsdCIjS6iRgwgeF9bzBgSNLziVMmnLiRzy5SZDpYnddPd
/OTA6zgQwa3nK7YHKjDcv8S6PA8asvR/6YADoHNoiyijFzYfKlYQIQ8VxAjfER7n
BG28ftBmIbep0HUgDydDZ/0NdhmrB5+6nEzXfsc45Z6lCOXPXX22eXKjX7mZ3YO/
jgxzMjoRNdsycpSoUnMp1Pup9KPtFFyG0zol4aEpUlQvrneJH44IMuBXrpTV314I
j6aI4vd7+5CnjvnzSH+sY2WVE40+yyZ9dDDrsbXwPtZRKbrs3wgJY2MUW+UjAR1R
MmmB3DVCNS7bJHNo5bdPqn/XxieDYpSR/yRnLAYk5b86QtvDqYOipNgqg5gSNtn4
eB6WJIKlC9OdBwjMjW2NH+ooKdUVl3NHcYyrD1TGS0jD9hMuG9GURX94F6hfnPl+
ZR6qDPgS/0NYikcanpc+Qg6Z0NxsgATEMujq7yXJI9Uy7D69+mKxnQsD2YvX0RiC
blHZNBFy9wfNJhEzUGKK/X9LfVvnY/z1lC6h6H48ua1lNqvjeJA+f+r3nkDPJhT1
2MHAWUwPzeo+RwjacYW0gqFRJwkcoFQiUnnTRogNNGyqlhd1VjcvsJftp30BB8n3
rrIv4rMnhp66RvwS6k6t++rt7RTuwbF/rYz03C+/fdNh3/GknzkQTVpwUC4t5EyW
W+tPzlz8i7gIrIEyk7onHjzky4V4Mg60GSZseYFvZTnb1sa4uM1QOJX4u+I3+cA5
i6jha0zwcsQ8LschJ1cOL79p1B+CYRGNjPDhLixo8mlXDQ8ndXlzmp8idNKX1Lov
YC66c7y7I9KBBjO0z1PcSC105TmyEFkLEN1p4KtTgnc22P/Ycifc4d5jfpW6fyKI
A4mlAKMZk9V4+4AWqh2wv7zGIq68Dni82YlCAfbKgl/2GegGfl8DYICyB4oEaKRi
7WDKN4pPPbm/RmOFy6wbw+5kAbkIB2NSTuO/lD2eowfCWXMrEFcrbsbip4vYRXek
wNQdqtiLec21JoKx1AI6Eofm3DvmsQvYni2CZJSyXoFhAkcmW5M8I32PWEK2rpxY
BLrx7EzwZaAqZS3wJYRyrY7xjUQRwfnRtiqz2739Qy7tO8jVUgAbMFzHIzRo/+k1
+vArYbBwo6Mbn6gF1yQaGwvyOJJwic/c04cVx5ujFDl7b2ANmWJG3tUQDwYg72kX
/bliPxKFxzzhs4BlP4oSPfNsB+sTwyLFVNrLyFhnnGiw+fKTTVptEmZ7aCFJhvr3
osMfqyXNFG29msExbu+NpkKut5yr8UkZrDL5UZ1MqXiCp0RH5sgodFUAZzLwK5f1
iNgU7qRn03uxJ+nTA8Nu2UvjuySvqqkaHFErtYQ7GNjwOelrIWuzO6iORYpyCrku
nBSkcqgLxrDHWD5+DtgEGzIlXBAlyKqszxCwyoA/NOsb1Zl9gqMWn3/eH/9/LjHp
PuV7qeBBgtip2W9F6EfE+isWzMZiQq7REAEIvCZeV23jr3dhSa2IwXYigz5cW0Yc
04DECJePGvQAAqrObgy3Jc+tcfkSgEwZUsm061jQT97CM2NLkdkmmgVHKF3nNl6w
77w9srjiKd1dbbaoSN1uBCuWBTEKjHGcAreMPujunjLXipQrayPklosIJi3mr/mX
7Tcb+nskzsn3R/Ks4Wiio9xOjucWW6YltBhDXCgCMcP0FHV0kyfbZuo7bousgP64
zWrCcR/WOsluM0PrZnIRBwS94EfXRGYb95CwG/YUrhQeyjO6Dh64wkEdRqoJ2a7y
Rp3MCxLOo4dNOZqPHnaREjKkxo3okmVIYQ6owhg0yGcrPnFn+o5dYvumHGEKcWr1
EMQaL4AEORouQvEMgIdqslej6v+r9ZOmDLoZDCLHSFZ+KL77+JHOFYMK+cMK2bNM
2RX59+v/G+48UF/3Esplzrkkq/XvNuVxMIT7LOI8KTdkET6nbr3mWtlCFtPU+Tf9
/9Ai3fzgcdcLPQ53179sWvrbs1uvIyST5siTUBigHmFgCx3oT1J13WHLEkfi3jiM
++/RfS3Oi6sBSPr24O0HXHDEJbHq2DwoqkqWgWCJcOAmD1y+yBqFpGhuQQkxTY0O
EQMVv9/9g/rbZHhTPukdoeR0yDWCd+6nOrmuxm9hzdugz82ZsTWJYsR6jB42RfVH
NmUw60KS7ozytSru3X+uql9+cxVH5H9g+ROiVG1C+RNFXXeM5ZbypNNPF9mkf2L3
+q9PrNkisyBb53XgmhtGVAqHht+pf7+wFjsm2OGYJWVIt5LHHFWH3NuKVEWcMAGb
NbL5/WOceLHFLwT9lBGn14HZ/U3+ZPIZYJ7x3zU95uZm2rebHJSFb6K2zwMIRKtW
HkS3FWeCk8hjRcdFberxu4AnTps8x4YzYnbQ44qmLVAR4UwCzAR8QKrZzEpcP0kS
N70FKH6sRa8DW+zSWjDO+ffNqsEP0AGvXXlEhjLzMXUKwpM/yK+0Gwox1QGjNA/b
zqIrpbtSE4lHFJ/OI6hXZRvOUOCSWumRrZm/xqDwa7XZeBJZKFjLcU/DkklOGcOA
Yrdd5Ost7hvHmZyMILS3uTeUWKMkLmP3ZLSmBYMLYS5J5f6x/gQVCfCzhoRDP4xH
CodnvqZgA1CpyKYT58l70lesrhwJU3RRf4K6P8qhvLQIS2Tkh7QgoduT4YvwxQKG
aw0G+YGXXLUb0Hu4sjdoIOO+tTdSaxFLyHSEmnGv3e1ZEvYtqh/R+v6ZBCX8/fk3
XnAovSXJ+Bkz/zczSy7JOxVh+IXAZ5uTOJbDZWsuV4esJ0PCtc0wAsbPqd5xGFrP
CW23eI5kDGar3WgjPXaXj2ScAYyc2Lg4DNzCgwDjsnbC+nCfyCIGOC3aCZrAGWJv
5Vhq1nuVJNvtYHEOx0ReRAa8vFbe6kppApPdT6NGZ5INP7d2ad9k3lzAcoQgS2mJ
DmAEX8pcYWfSYUZMtc/TCs3EfS0udqrqs/H+DslFTNMkn1sKFxbk03LItjkmFUg9
lkUuCVsA43K37CHb9AUkDL+VWIpg2e4490hbsNgAk3yMR8XqHVCIGMz5KMx36xw2
4dvrsxjEKELYRvU+HcJI6mH7RTIidBWjnEVhxzQtdoJSEBjd8cdbDxiFoOFi0Uwo
+B75JYZOeidhbmMgMGIwvjpJk8rJwgtGQhVV0g0Z63v6ZerU5mLmB3tCt2QKI/JE
xomXaODiXd62rQ/U2AzYcCQm1zDOj/a1I/WrrZKB8LFKIBqSrpVhZZZ8+POU8oxE
JANqJ+DpTK1zwQtNtDTQbXtiFuPfMuzIiZdoaMoN1jlDclUxbYnFVSk6HiQlECyV
4F/jZVwNLyM8O2pncOmS79gV8e5NUMG3b4CYb9fRiXu4Z3gJH8bQhKPFrp8yUYVM
oAGUfRnxeeqDzQV5JrlWL+e9YY5Ank1qOzc3/oChuUMaZlS4uyk4AOLsn8mOI7mL
2L3M/rJedltA2o/eOIoO7zB9ZZ1qaRyaF98yxcEletx0M6iICz0KV0RXGbdLmeSW
Q+u4qZYaMmy9ZHpOoRvrSUCAIunGDE89n0MJdr2Q4sH+h4+M2e1j2mGCsDg7iqJR
eVXLhYfRSpay0ZeM1rSRUytaZXnPvGXFV0ebuCS/5LMB5yUK3sJRz/3IEMKZXLkb
ZxNpG/6RZXYreNNwef9EStqHJXBaN1n3KmBaScPU6QM8wf3eK2/swcKmqvvtVsTQ
qXXCEUs1KZ2JZahtRcAGSQigdWJr8LPV3KGLdwfm2tAtBpkTT9hSUg7H4Ls3j3VC
ioWCsIPTnNxaDGVYNb+g/eWfe+UYUdd48IJmCDzL2V6IUh2FMM9eTO3xkxsfRUYD
h9aP0CH9yaAzyMe1HRKEd0wls63We5ZdGIQ0jWLDJonngHkjqnPA0JY7EZQtZbXJ
YMixeaCQyBKm3xW0/ED8a/XMfVzwJ2hh0AuW9QGQ18UTsgt2V3MjUFwO1SCOUkPx
50jEddZPLPtf+OcUOCjy4gC6aC480KsOjDwTKdd0RRo9JWEKmljS1seO1B8i73S+
jGU7bnxhu1Vfm4TKkuFt3gHhhp17pQDSRAJ/y2H8njCf5vjSiG/jmrWG5ITCue9q
qrIWw7l5MQIV+dmN/l4olZVeFo39lw6c+R7/EQBq0OzfzQLFIlI9bYUUgRj+3zA5
00WSND4gWnJus0aMFiZYYgtr5MvTPaegY7tUB1eiFhX6MAaGzFkBdfZvp1iCAEOE
YZOQPxXvAssAHO+OePNidG9cbuksWvMvgbmAkxgF0vrWnT43vH5zl9fIcK5rdoyq
IAVROAPfxJvPLzhXP93VXLLXI+HqgQfYShYNbbV7U/4rPdJICo3w2Vp46iKG7cIE
dhqjtBzqvNBawsKYb3a4iQYPaFzzYraAMgoijpw2N8KUYWQrdGLjO3X9bjCqWS+k
X7c5l0zaDE6jbIH282BniwACoDEWOcSletgklDNSWDUBQxy15jYQLOAj1iPJMh1C
Y37BH3/32DOvBtO7k6fNg3EOw5EIy/W1wPH2t7J7zxVywwfyge223aG+Ng6az6nF
3IfThmRH44SEL/NeO7sytqSjzQH3KZQbg8jljBARZb3My7pc/VV0Wx9OFjsSt09J
ywEzi1yaPfA8KCE7eR6Ho02mkr3QuBKyUI/0SfqMb9GfnXtzwNJidkrYYNWzcqTb
DZp7g4FnDFCCyZsYk2pcFghh4Z9FR6affOCTP17lZRgJ4/F+Jf8ZygIQ5al7Uig4
VkBMsE2AzWD22sxqFiy3C1k3ApG7LII0o5wl+Sgl/nph1OQf+4ICL/eJK63txVek
DiOxeyPnMUUwPJhFLvSNxAWy1tF7Lddf0e19XM4K6JQrGLXRVGVF5M05UyKIKcoT
7OsBQVwc51Eh2sVuaHy0jy09hlVaUpBJNvwpoBo/OrXIOrO6CTuYuxUNR7iWC5BF
GzpXv6d1qMV6snl4ouJBrqqVh0pPmLWouFm1khjReuzG0ngBvVM2Tr9LgQe1tYaB
rrEY8MXzqDRJxJTRcKoZtkrz8qQihKstFo+lZac/OfEQqFPfUX5C/3tanmUP/F/5
VNjL3qZn1GyA/1EukJ/IUXPCoho4QIy8HBW/PuG6e0XrulmhOTZKJzlqhP/kpfbh
HKLe9KNtswTXXxqSEPcXpSCcaKvo5W0ex9fF5xpOg6uFZ6ADPnVnrrpczo8HWKBk
2NdBCO6VD7q9lzJWOoYTkswejDfeuzo9jscBkek1LcBLrTV8RD3AVY33DyzDTO1k
Nx5P2IZtCTZgKf5VdPY4Q0hVWK7/2qFmlV4m2lN4gICe1r6dU8IbVMbKiPGGY4Cv
/BPpQmEMEStbjmQ6PWY9lkaGg9g2A7SIq5yCc9m5HuvNDJ1WjfsJ5fFZjLnLOh6I
N3HKT37mbPiYAH5cKf/Kf8M/ixvNVoBW2QsFYZNDcwj/PdvIniLDYwsmTipPmSwf
ilwZoJBNgCoG3wh/BheFNLvSDQkX2pS2N4pfS7er46vQMfmPm6+C/tDGxj5MIPYH
awdmtBvDI0OcxbALxjFuhyifFOJXgW+cM3Q+YUVuaZTGgemLpPP/4YvJOe0bwNt1
TKPcaITr7w+pNAk3JAUbQiAUvPw8CSVTOhe91B8X3lQFzp/N5ZOYrwIUTFiZ+YWg
rDiPPqPSKO+Q9R4e9ddIQQoFYGB/LuJL6jdkEcG36VOuLDMy78zTx9/tV1orO4Jq
g9yJ0KvpO3eTWTHlxirWpGeC/9koXpJRSKMNCahu0cCQGKyqEbPxvIj3gKUOM/Sn
DFgpQqclOkLiVemXEzYaq+IAmhsMFauLFAd36u3mzIIhGxsT/4Bl8MyfTVLH2kqv
ziqDgBxT/0XsCLwGOpnRAYpJ+38w6QpabbgSq7W3XvqpSQKMQ48JiAZ/YLjxavDe
SxOLFFvR6bFUXGZWphWuZP/VVuQ9QZg60G3zsIoVP02yNRYsZii165W/PtdFRFPj
qop8NBiLHxEFX1jVvcX6vcRvmc1XrXGnchcHoxQ9rwexHDXpaF9biSMHFLhDTd5k
Znq+XQHwxG+i8kr7UgARw6YRqu0VUDPGQTyaOe/pvY6fLxAgKWSCsuXbqUCUg1IY
iN894a+hs2ch1i8LC855fed82LEzm6qx0/2OMjkQbMTitqqxSWo4+vToIvLISlV0
hutWvRmPB+eAodgEhbMZoBSqLUpW4CG4suRhZHdgd+ourFegUS2M7TaUOyLfq/ft
y16ZE7r+Wk+bWLymviIiK0DZSkpOl0tBqqxhQwZlIOkm5njPtXipGtEfYUIGgHMy
9cFrQIMoiKfpJBRBIdMmdXCyqbLMd6tnuB6Q1JMaYKXQjBb+SXy75p43bTFNYmnL
tvjnAgLlDNUdS6mFcgThNypYqc+UnK99tb8d2fW0pZd6FY2xskNDtTwDUSzGrvoS
0YWoK8W0pSOHQwLPoeJO7cHusrpFJSkNAVgiPj64uLyxkGqIfiw+osxBMZPIG9ri
d5qYP62KH5TP6SqsbS1IcZ3ugGn2qJVT3BTJXT6b3pWJBnDxd91NbdQZ5yNbdLH8
VHmrCHsjy6k+XyTQia8WNu2iSEO8bGiTe8Exm7mUjzghIQy6T0e5sXMI8dkjDavT
LQ1oiD/Rfb9fLHkywfWaq2i4KIn2MtCWy3ofgU76Ti4PD5Wf9XeXhtK8s/U49u/c
+UhjBlMvhtsSO/g+gyr1TxBfdL1FIVDfrn9LDqXSYiP2EYgmfElNH4S81z90C0R1
bqwvXXWw+alZjQHojIXs8AIL7Vk3qC0AGJrW1mKmitRyFql8iEg1RkpJxVmI9oCG
UiGzQw2em0+qAKA7+Db9nSP8sd6tqWJ3FwoKdEjo3NojyYhvcHBuLCU3nOeeEBvb
d//ardsh+6i1hmwrGfb6zESQWDXV42rw4XjpnXQZHQDJyf5wLvOk3HoNVTUJ+Sba
MvConLxRENndHo9pVufQVQOXUFlq88sOGOuZL3fEQeXUH4Q6VXSJt+Zws+A0B2F/
afHOHUprL3pLPZ4NzJbYNiT3t+aRGZ30lg3Tzh4P97NSNxHbSUmZLhuY1JvK05sj
fwJTeJ9GsozVdFp6AbdvzmbAJhc8n7B37ocuI6SR0NMV5/DwrpGwYjyQU0BP+Jlq
Uj3AZwC1MXLa3aCGYUWzofNCYM4xI9W8gxAVRcaSfxMEUJzHIJkOVALdF5cbSvMP
BjEfPmby0dVV+qzwBCVr7Go8u34vx6nMfBrU4P8vY92FJwKOTLZX3IFPft//G9SH
22pL04MUqAfIfhkZQ7f4EeYUmqUtsD7ckWkMV8paM4tR913t2fD2WafCdmMlFwim
5YqbVkWgaUrvjr15ibhPDOJjcXNCQ1jrUUz2WhWOtw1RAjMpaLte74wqIcODaMx6
Fm5hyZlDVpD3Eca4MmmsaYMOBivB9XvrJdo3tskD0i38FgJxuvpssJvI3+I1OgPQ
TdWsvLUK1HPDU2KariYifD8C0GlcaUZGaKUFugOB1nm/c8seA+H0MQongXhZ0CFs
vBgJq2kMNt2jP/yL7Khhvr4Duh4ap68tmKNGHnU3NfNhwhbKnt6/vYy8ZD4cxmY9
Aalk+9zGdD2UMi638mGlfdank90mUcfqQpbCKux/sz/UNkwxPRw26uDrpiyqsC1U
LmSMYkBnQlaG+hUw4q9e5MeKB5NolxGIai3QMYdmAD38u82dCfY+t2XzrxZd1M5C
Dz3WuGvC1hn1XxDuPoDhdX73CTzAUoKiSYh/C3xTnC4NVuw6QY0ZZHpNVD1nh4Wg
dGECddtfXDOwKq8nnGI6h1vR4euUh36BZC3hIo2wxEKh2PCmO2tjqC+pSbu68Xmn
BubkQD4oYo6fWVi0XVkETiEbI2AxneyaEjI/qaNLObd3AfoGPCcENB/QB0Xp6aB+
UfiDTo4kXPZpWOl8Jxu32NJcE6IJxutFBoq0V53M40XQaPWJr6u+CG5z76xJm6cY
7rCUqX5dE7TW89d+Qcyq8gFCcKK1UskCUwGVulL60np4vclOMrw3cU1xer4usD2O
2Ja5TUuRze/naB+psh0MsktEvH3rDr6q0iZx8SRlAYDbCd39lXcJFsVQ8C6z+Ike
HVkZvG6L74BOwOipn01+nB/2eLp6ccur4g3FtcMdCFPnxt0IgHWodrhzIgUXDMeb
FJvsGshQBvR4q435imOYJWuSUc78KLj8mZIPrTBucl7/vhihwxyGqdjm0rBpSYae
AbHS7V9A+sD1SnH4h7rgfXN4HxeQW7Gk4wrELGE4Rli0YDHUWoVUJMg0RlhtaS2B
/MySavbOsGCS8FfWUEx9OEwCbl5qXieBBpB7HYvONl6SyAnIu2QL2MLG6kAJL/n3
UjVKNyiF55439gecH0DaSYSI2DGHBa24WXXP6+/46hJV20Xw80louMUK0YMJuyiT
nAclGX7znrHkz1eJtIuz0jpbnt1ABvhfq4YElIA38hWW6FQ278q519akPemL5CAb
iG0Y7Z8OJ4iYuNSF9OrIg2REGjnhrwHPSeZNHuFK6BQX59g/O1ICkxcoLP1zHexa
6gjJ+NdQQdrW2n8spS43998bo7cG9mrRDxdi/7HCWA13VY4QAppUpjrRrBH8Q9KR
HXsVDKZWSWdYu1arhmWKXWXgsq/eGsPVcMSZ+2sU/Si7WPNf0hb6ddkJhe09ecg/
nMACo+xgBa0qSN90mYbm5FM+CsOy+ZPQ2ZM/1j2KzczzFlpRpjsDk7KTg3BqfxVu
LIccfDNf3IxxJSypc/chwW9JOGmMTVNYPpP/XhncNps/av2tZHFDS6cpf8Fbj1aL
ZVv4mwXYHl9/EIc6kLiPNkf4yEbA6r4dGEUAu+yzVF79lnC3KoC4HAQb53yAYjZG
AB5lN6CynUuUFkm1yZF6qFNdJXzWxT9VzY8cktt7ugsJBg4Mr86rveigbgt3HKz+
bxHevXh055V+g10p2wxkSZuTvznoZ9igSLknHJITb6QFFPB5IyBOVIP4RLLVEhqZ
Q2EKB3Y9JJnbCCqxPgOPoggP+NJ5XBAJdEon0rdF/8jufoz1d97nrw84Lb3PTter
JFLWBUzjcTL3QVCbUzlYU5CaA17SXH7KrA0oSwZv1ENYVmxVA1L8hoqZ6o9yOgCu
KRUVQnYuYr4fqGHlA9k9dlp77GzS5f5o/rw12x2NBRlTe2ddmfA0eundZoeq5D/U
Kg5BwpRBPHOroDND7T3bFqD4Y8JP6dZpDF7U6fxWz0ra1vgvMnDMZh4my2EcVx99
krGxwSHYrkbk0zLMu9ACtHAbqmTBVi9+j3S8RUcmXj9XThuIQ+0ujRJ/4tiM13Ky
9gcidKaEzT0vUrzP6XORPjb6Tu58PEaoo+g1RTWvfcm9FS5SvVtRsbBcTRMxid4w
RGkJyINJi5XshQKaQsw3nJepgIyTmpaabSXiFjTjqvaHqGDKjzn+qz10KWGRQDAm
irOrTMA2/8B/BmJPeuHq9kFANNsjwl+evrVhAvKCoAPFtFhpqSPXJMeLWc0VRVWU
2XgdlY6xgDFimAyumYo3ciAxtY6M8N941hdyrKI29heBCl3+QuvaGYVglATtnfii
ioKs4UGu7eW7hw0i/WXGLvxlgRGZTyjQoHiNtPFKLHVlnZWf1YGpLJBMali7Qszt
zoHCzWwpvjXYhWrfNUwiiee+lCmX0jGanBEylhX18p21w6R/f1dexkeAbY1GTwuu
JhWdei9xUfPShLIBaSQqoDgbwFqjnW8gzFJOn/YevURrH+Ju9Q8ZiTwouabMJyN2
Wk5XMzdGYlaR60fO1xoLkRFQ/rwwDjrTzj3AbZASvOZfb5LZhppVHKcpCI+vYY3t
56IGJtfRn+T6qQYUAH84BWmFUg48GfuczcYVPrttFmXXQhb1n1X1mRmtfgWciW/W
O554HFLT0kr//z3eYbXOwBAGjuKUdxdX6lSqO8yrHv57kO9pEYi926LJdlTCj+Cp
Dz/ZhwVWyJOXy24Zmm6lsbtIAvbxFnC16N91lp5dK6+3VOi4F7Sw3w2jQM+aMxDk
frFuebIIWeFb1J9XER8tqe8UKoIWyUR17DEAVG4kR9Ad47mdWGLho55zqI1Jz3j7
OlIsfkrJSExdkPvrafzn3TG9DDGbH48lzsFyySF2/wGD2RHzZWoZ/KVqmWzEP/xm
GqfQoF+FA2JEZgLMG4StJBR/FUZdeOeOimmeVuFSblyd5U9pqJeOR8shvbIFr8Hg
uASYi62FKbG+SbKdtIGa2Cbw9IKHpEOR/7izN0XOEfvRgVof1soeEx5+i9VBQI+8
b3vfKUo1+J6dsPnxsG4idsPeHo9wiwv7zcVUwFjBO/HG5K3jeW5zizQ7Ydz0c4an
bBVgWpUAwQH+0u0oGckOKLukXy/XEncgH2TXFcMp9BHge7Dzrm25uaJrAGunh8Cx
sJHB0ZiUPPtw+ZuNofys0gaD4iEPj6mT4nfolA1nK7wm2qc/PnPB/vGoqBKRaFlC
lHQhaPIgF1q8ObpHaqH4CtDfERKMi8f1PZ0CAKBNCPY/OsUddqK6q9AFxhXeswuP
OECpd7BOI1A96Cch3EyrexlZl6ru3v7cCtxVQBFGpaTjlOd7J9uP8XseLVJF0FYu
06dnvUr7bWEmaN1Gt2up/HqshsoB1j8hufyJ7hmxTBCkWoenQkIdHMlIi3pPCEU6
Ww6Kh9vkYlo4YwSLRiek3lwGScB3f0Gwk2D94hgd09Ibmz0bO6tZS3NvnYQzgW0P
+3mtHpDfvjK9xi2G04uht33is/0KpyEZGBrudtUX8iXCcbatUfA2f6tXIudu3U0h
vaEwbpI+EMGYzVQdz+nOHeZFY9wZsiz7AZKTmAjsFPJ+CM2Wng0kJMXZmdhtHvu1
Vq/tqrBTtQuRZIE1X2tJP+Uz1V3Qx64RexMV4U4mNDct+Y9gaZwPgGw9v8PE0m0j
l0KibQy4gUX65iuYkLHboUmYzg7IYDdWFITF5x5pUWlpALB6zOduT4xSGY3T6TJm
+QmrUauVoBE5OiG2h7LYkONxGtKIVfeYwTx/2boHkKS6ll4RI2tJAq85P+K1NOy5
83ZmmBH4NLEj4S6Z5sWkbHxUxTnkFiz3xC6nwOeQiE6TidI0ABjHSdOuGq+0UkEQ
k8RtW00jpO8DG3QbfX9nAWWD08LhMnD3xJIkZT5+NZ+xRxbxOTg783rn6LXa2wbZ
0MBTzffhmNjia5Ck/2QqoHkJFz2uJ6pDG7HuHp+n0zfeYTo2508357MtiHsOyjmc
JJVrAO/4/7c/UwRrTDhcB+KZ8BSFEWoRSELB1AS0Tbry4ly7q9lSq83GJEK3E44w
gfg9S8VEHaUfRFHTQkJp1iGaNf9wlHIKTiDTwIKWmJTzcs9ZPWKjQZZResgNGiek
2QNQMN0wzlIeJAdZrpFv612r/ZBDr7qDHrNlzbqF3JAOD801Z2d9DFeINqx+NpA/
GrhYZgfozmY2oIA+U6iYe5DBcmpAdilC1foPRezk/xT1L1fGN+DOERNJHpPMW3FZ
Y6ZNy7G/O7MYHiWxn139gMVN16fKyFqV4dTwggIqv1hL2fxptaBnIzWcdmzXQ1vY
muY7TKENCnOqoBN0AuJNW367AZwAqy0tl776zhr0sOW5swKGStFrPGdhAILBjGtn
IeLGEZ7gYAmIpwxDvEo6YscxkZmARDPBpyqPArj2G+r+A7hfjxGtIBswrWIa+i7l
imnSOlIZZX4pjvrnH3xC8wXBgObQS2XRnx7Lm/3H7vTmOvL8f11uvjJoqF4Omw6W
kztDOixFXhR4/ykxt+D9R3EVrwqsUaBMhkl4BHKT29AHrzdB4+M4XbXXdGv2eiYS
Unkau4fDjZBIj0YIg7fAsQ4OSwmT3+13u2NO3LhbT7Ed1Xy/5CCJ56sZNnRamooj
f7yGkBAY+r9bHOt6eApcwhHiiNEFS2lgkW1hPPK/gFOEtsHG1ZEk8p8TEmCjt7oW
Q56Fpd5caO48GC5Vht0ZKoa95JgZNpNfbLs0XL7L0TeI2uBFltkaCqmE8Xc+seig
zGsEwkKwgToHoNnptjojCocFtr7LF13bJQTk+ZfXufjfssipTNBmR62nYWORNq2b
M90TLLnS+NbNgawkBwH2K25UrJQd5N3CfYVha06tftescKkEg57mq+s/g/BtB8XM
ETBlO5hN/JR4k5lUexnziEOOiHtjTP/8ae2DL6Ikuv4RsYc0ze6dfIdkOgxoJoBz
+9308dOMwb2SmyAh6KKqFvAbp5sNWp5e57XUtKKPUPr7Mfgy9Q6F2k/hJIoxlDhP
zdJSSQsEKijhUSPWIIQpOVZf2DBzoqg9/fD+dP2gplFd56diSGk9wn9iaODO3nXo
w53byMTtmHO+bvtrkrcBZklEqitzwIPPtgHgqb1dOclONmM4Gt7MJDO2tK9VeOjO
9p+AJy7DE5a6OLLj/eYWwA9QYSX6zdUVAs4x7UEJe7ZeZQ+jl0qkpSeZTJX4Cnwb
Yew4KXJvClQTqNcr30ECuHMrJevqkavpQ/4hHBD4+t6HS8iw/SMRkn9q0K/HPe/8
y5HItIA0sqvdwXpQLxk6Mi0QC5dLikZTlclpD8ZSgo4EQuBBaKTsn9QvG3mqVIg9
b3rNyH/DIRTBC5ApYd+7qxfSPf1vHrqQM3BRxSW3QQTpnQJDfgIYa+kV44cV2V8V
pZ/+hhQCEi3TvqnX6fwReJJVohIqtWnzyW6L91kTd5SHubaO+zz4fk5Lx6V5ZVtT
3/zykP508onDZM8p6kH3bbVs4LuzmA+vbVS8r6Ll9QWmeuDHf6hCoDZ7FIuByWJF
BUeQIb2dMB3wN/V5Yasj4bbVTZKV6qs+jAvEtbEzzY+G/0gf1/BlphI/o92KqlIQ
AfH1s2zH8OzcpXj9HmsnfTKROWHeYJp283PZZ56snabl8w8qgBWUkKaUg7YhV6EO
AFSzFpLvvY95eBzv5k4nu6u2DNqincH5GkQ3zSmQzfoWxg1k6v/Md/eUSYTo9dwU
FpKD7Xx09FGifhHU5hZkQdpkhAaLLGu0GWpF70VfxPH0U8CpNaYsrvd5cVkc0ax6
3tD0CIM7d6wB1B5YXDY6F0+xk8cmiQQuYzlHoI5meqS+BeTp4Tp5KedtN5bf+cuX
LPEtaji8oPKo4ES19Nt9AG/tSLcWV2/N+Vht71bjQ2mnarQmu1Q2VeFVryFkncdK
qzDZfAzxzX9HGpBFP8avt3K3fvlahmb9GTfoJG4AURUwVjnzz7Zb91wVRvu8/bqE
LNAI2IDJP5uz7jbh8CVHMaFyp7v5+sFhfPbV/jXBx5mta2zG88T7l31CTqkC9/MZ
c4jbct0WFfu0zhUAxSqSiiGGce2I6S87fzRVp5tUQxg1mQPbP8ArlZ+cxGIoOOoK
CT2N3OFPMDLmcSN+O8S+ivXAiK9yTw8qm1hV1Bf+Ht+Z+PpI50Q41hddWBJ+kOoZ
I6TwpaSnFkYL86LQBZj6fR6hEUK5xikHXy5ccO/Dx906pARE8xxNK4rP/9hy3MCb
vAzcoQMtFOMviIgYDKWS51u7SkrSOxebU2V2+ppUwITblz/d4dh8ToOS5BBB8/kW
WpzCg02jnFCX92zgewZI0vTffR2qt5okXRIF9tW2x5a5v07vFpIO+PFACz4DRfUv
vuRzmVvedq9BUQWQdfkL36UTvLDYMVUezIqZ/G9vcJBLuuigj1WOlERrBxg+gNeB
LX0y3kfX1pJCn8wOhM6LT7h/SIlIPkOggyAV4MfyoMMnBEruoIo7so7d4r/NhoBQ
Uh88l/OhA6ORTAnkLp19tYPLH8Jd+EgD6QUrfVZkGwtB59saakRpG2giauk0/l7I
PzYRuvraykkQ4vyHx8yNlvw7TwWHZXNWd9TcR5C685aGDlkx3I+FTKAGrlTDJu9y
nOWJuIma8N1xD/Py05dKjrWcdu/KT1C05SmH1C8UKJ8rjA+66gbcZsb28FwOta/k
lGM0C4pU6AP55ppn0d6lelqEI4EaMFa3bFbh903mIw5IbzxB2RsKbtae5d3jo3M6
wTZilWTeuXEI/0zNMNY45aLZ3DRLff1aBWE8sB8yT3HQKXKsQy0TLPTITIdEiU/C
G78gFMQvZuKaEGqOtmNDIsC8wlzpJW0VyHKi4+wG2KfP+NrlmFOw8gLdY8BqGJLg
p7hmh6cMT00n8FWUC56h+KaVhktxhTuw+bWn2jicvJLWjsmNIyZfYWX8l4EV8BCH
o1bf/CYcRhpBWcA2tXXTrG6dnciK3lOA3P2KAdqTrZAqei++DHgoKkt7GDLcEaMP
YqFiloiR5GvdVRA2Lsa3GIzpsNi2rNBsqqoQFoy2ElLOlCB5vgqJXeXroDIFIGne
QmX0L/bcme7SYhLtKLDyWs61k7CqLtODoY1J8R6BviybiV/kzHUH3t5Khgo8xDQ8
Nxptq4EVqnwqx7mMXtZGXTrj8o8pbQ8ySO51a5SqYWgo7X2vCJqkAiiuXVzcGKqP
vPgSFphUSt/WsM4g/YogehsFrVCbSUwvGr1ov2oHHsNGhX/navwBiEAy4oF6Y5z7
FuhdR9iCusEgDGw7gh2S39QexLVQ1iSUYNoGzx91WLzGRUsIOYcOJv35qnhAAZpP
IFW+kJpe0hHk/5kmBdMgkhdyaWTX3FqObNQlxflWPrU8BKR0dUZe8bKnKHKQkVD3
Z3s/+OXhVVHFx9dorJvw6jmZrSqP1SmgPnEOclLbnya84Z8qZGiEmJevfVAwy2U4
T1g5biCHtSwhsaw1iYuTzTRi6W5SX9xIj59JicrPytHKq9Asu5WDapv7lxPGN2YB
dg3QSBC5otbtwz/48SFHYFM31WXCgaBlCghdPre1WQIoVWqC75WNHmlIZv+892Cm
JgawY0bNckT/U6dAcfhUsLP6dAUJjPjN0WyvufBoWM4y0W/9VTN+tptBSpiTdMFW
yul+u8do4JFmBKmjL0PANWuKIpCaI3MxnE5RuJrWo+ORgmRKs0u6/0sinsT+BhfY
0SB4WHX7PvWDDItNzKf4C6o6izqoTMkeJH86LU/Bu22AS6RNRIwnPyldj8EcuKM9
6US6TDucjaID6ESavpYaE3m2C57eyo/oU/oBH8b6EHgszFgY0sBTEwNbqND8Gz3R
GdbpylMEGCwcyrOuGu9vQC6E6vHZBqdD1BpW5v2P0KRUsTMpwdlkbWXFVxLlx1pJ
5Zqo9MKcUDGnrQRkvtao9T32C7VPVHZxOK95T0TbZNA/VfNvAntU/qkAJtEh79dW
lCMJGB+mLYxCMQWESGPvGp2Y5LmFFrai/dFXcuk9kzYj+5NkaGoOFZ0td4y6qpGi
gCIaPTd5rkCF2gwZYoHBPumkDs6ziS107Mmw8qeBXhCAPzH6yY8urextcVsHCLcF
DQ4X25p7y+dUe46d8NpiLff5LNTBJvYZlgrBGActz1avzWin2d6399MY8MXc1XAn
bdW3nUfGfvEaq6YWir1iM+vPTcyQzRxOiT8MY5iulkfmDYLWVMPlwRY0wRlELR32
m0dUCZRgu1muqjYGmEB59MAgsHVjNVfuB/R2DBQ/vkZ01JZYkROymQvkYHv8UL99
ifetiW9wIzExKmeHiPkIdeGAyrJuY3XaGXv/pz6vPNe2pdd3roayZ8HNj6nhFVsC
9uwuqIg1PhZGSMJ+sLc9VKY2NXl28PWO6wAsc8fmECWqnKhyE95RiRAUlMIAXlX9
GyvhtHc0UnJnvqPRPuB+FZbZ24Sh1FN/ynRcQxH4R/w2j942ef3jY8P4ueWW4K/B
3GyOH0tGoRQm96DCGrhcUFJ1XyO+qGczC62KPhsJDf/d4ghJ9Ga5XM5yja9QHo3D
DRW6yAhyHsoOEgj3sYaarLo7e7S3fm0EDrASbdl9NZHlCJRS3UQRvf/X6dAxtAPn
LrBb83CCOb7udIacoN3pmyUerazZHkaBZ2Ix8azmefJu74un/pZr9yDd6xQSkPnn
VhOgBoZM0vJAkn2kcWlBW81e3bAGZUwADu1ZsPM/NsiFCVoi5yOMNrvwTBdDyHQY
cPsp2DbBAh/9ZfrgyxW47/V7g6Tyyhuizp+xXiD/vpqBKXZ2VV7gkoPChgwsaHfk
aDV/9r7PHG27HfML3LYI666bPVlKX/2YO3Klclkj+IqSWu9878VBGisD9JB1IEVL
CWSUZUhRfiQuJFlH579Z+S+5tdsWL819r3FSe6m+XDYM1GESnLBjbDnxLWQyM+PE
Mqmt07MJ4FMGfmvQn6cHXLN7DVxGM5/qzoNhCL0uVfxee94v39XYbeHxYxpvR/AJ
B6jsrleAIuAXXRvpmm0Act5LEPr0pHy55R8Kke67KA/Is0swMpZ79x3ViOocyCSh
Cgp/PWaXFRN14NqyrC6AVo4/5SLUJI7qFJuat/tSSpL72JuLgYHC6O6dsce9d7yf
v9VGxokljuMo+04AAlnvxFTuW9yrUlMQ4MAl45EQfr+HT0w6k3uLRUPCJ0J7sFq9
EssdGqrikRyl+0sHcJfV02vxHP8qn+KLM8UmkqieLDn532fc+v6BgdmpXTFZfezo
6UUH6O6PddeD4wZxxdcU+nDS+thnbeYw1d6c6SPxKmT2OmPdHzHnShwRHREH5ga5
RkQTbuUqv+tWz+QpaP/ZmGvNqH9OcDMOm9Hup/XfWRKEIQ7wz2iKfYYUdWV97Ass
hsNpRSgJoWTMICddyNTNwZqJEZJurNUXWcBbZi/dI08HhMfLay9MuTbXy7eWZrx0
KCJz01jqDhUs/lk6A01NcrY3zcyD7LXt4K8XDkgMO9smt1XpXuXm0LksXQGYhmUQ
qFyQAd8y4VbKD/SyBFhU3hdeeJW1oS5APFxHacTMb7ImiyXJqziCz2CC2BtCCclC
CwF6UdlgCax/34YXgO+jdls0R/eoS4Fn/Arxc1PMcXyceQqvR3t82VN/APginuqA
Y0emh7Qeik6cvdkJDS0lkk67aFUpFCOYf9Xzvdyidw7G31FNQ+Pakx3q+xItBsLI
SjX6xsMNB/9uledWpozXHPs63O2dR397PXGuuiwEhh2jlZb9Y9k9pozgUpfxQvQs
w7oL1XJntrEGKosTUVtC5BL4i8pRsvldvaFjstOJdeKkt78JJrss/7faKrFiPrYr
Tpq6EAZM88lGkkY/GVwzMN+53Kt8Xk5ZiRuAnCh1Pzsg7+JeccPlztlNvxfx6mv8
adiCOcwrTpe0JNm2dT+EN84nm35nIZhU5MZpS8OFrhHGnY9Im7fI0935n8OJdk36
nY/reWLhVUO0vRqNp9ASGljsNPorfvGoqk+2TI9uCyqeuiYO/HWrQuj7cqRAFJBW
6TlcAbFFvyteaCvdYoE2Q/ohcyqvN8Wdsrfa96g5BRQJK0yzzJfnZufe2ssHtg94
S+rWbcXWGGkUPH/PrgEvLoYdwjUQAX70sUasLt4w+ZZDeKW+yAGKA+vfRytHR7Fa
uyu9+eENVTczqwagKIVoRi+EfdxNO0f2yckC5AiTWqRIMwbI1ht5JpYRw4IDkEg2
a/pOAEhZgPMQQxk5LtHzaKBAQyiW1ev5bziDaISNi+pRfWUQ0KzxDVYctHBx1HoB
lW+v7F+paCh/UrDLM+x8p8jg8Pdrm7jCDCCuA2XG2opM3IFhxZIqiOJ4zQwjnojv
vfU7DnCOnxgLV3WbZjK6AskCSdvT8KkNOGItFon17MDZQ7jBNoi9sWISDq7J9Lf6
wQrbMe9i8y7tZoor6vJ4WSn5so72yEULve3Ssr/Ifs59yN7al3PG2MYeIPzCu7SA
e3tjh6oWhMbb6KVcweRQmt+SD32l/9P9xNy8vPOUh84LuESBL4fQ1BFiwTYUlyd9
uI2V8QMMpwf1Qhebk00YG8hEpW2q0jBpoRsbQ/pFvN0BFt+DWQ/N6aEMal7wz4s4
/00Tqv9yBdU0cuQOnpZgF3xKrTKr0DbygLkMhlF5ui9UkOJSpzGu7lmmiTgppUp1
pR6xwpd2SkOu6TRQr5dJKqvarUE8s3PzO2JtwXAT3B4HwKRfrZy6b2f/19iac6qG
fIjYT/JXq5fAyZgleeuLy6X5v1FtRx7ms5UZpXpmLdcgSj6DyBAZdKblhUCP/P3q
AaliVsOloH7vvJGq730SdmhOK53jxpZGt1XrbG3PVEIRYPGlnDqUSZ//4SdGosH7
NGv/P5V0uc5uONFFkxkNYSx1/wWL3O1ENsezdEJDtVGjjNcrvlXKjb69bJ4hvHQq
v+sm6EWWpE8xv/ICdN3lDSr4o4gCI+NSNMxlYd1rx1zgDScg4iet3dBIlS05QSrn
Pp4tVcA5hx0cbDhR2bW28qob7ielPztNX5QSx3d1Ec4LhvPnHe2HukQWrKoUVCx5
ndyRAsZTae/DNNglXc8x6DJxa90qHAhoEQKpq8QgDbutW7GyYvsDVVkGzj1Tfcl3
5aLW2l5kryvSVSGduBddmudo7momKhRDBgG9jCFtLqlpGNow/qiLqAAOk3dcfd6F
OxkSG7zNkbyRRwD0xYvWUyU5E4QvB8XPo0S+BYLqQkCar9SiGmL25Z2k6dl65JJi
4zMYiN4qy7R+m8teMXc3vkXa/mhqorzcrD1imkVWesHXGWVerAH0CLvKVtSEjs0J
Ck5Dod+3lH80HQ492Qhsn+9d7arZClWUie5YIdHzPbwo8HpIg5XQYbzsozTnygxM
2g8YbS0noCu79p5yGkPUa+Wg9njdM1P8plhggvd9kFizRnGB3PKagy6lTLfSxqk7
cI/x2oJGdokBVsV4FKxA0ISwImbEW/rEvBjIA/0uhdxasMJgSev1NzDJMh3IKyEv
6MTelESCDKKiqxhlS0/aRorVC5RkFFiWKzrXuvH/2OCgK42i7V3lSVP9uu+8w5ua
wbLg9ibMV3egXURkFNznc7wAcNl9Vqg1vhwA8ynOPU4eCdWE+YE+2HT/JkVY8zAh
Dtyk5vJNDMu5TZIQ4sC2+z1NgVQ6p1+TLNWyzK4BxgPkQDp3hgzzZ64EM7Y5jz+k
ApyFK5Wu3JUKnd1nlWfeJoW14LanykXKakAaRB983IPlhRt40T4w9vzXJwTyOMNU
BdzLHRsk65IgNt9Yq7OhJDCVVYkLw3gDu1cajNJxIbjDEPbC/8IM8hfXxBFrHuQq
vZ4IDJwfNePDtgUAwVcaOIhxZJ/ZViapWKEJrJBq8kMAenj0iSh+ogxRMm0hnzFE
fZdczTgwWuJDRjiQKNAWTosH13I0TIaI5olCjFkjZ5ZWXv6pgsQDmAcF8ReHp8jq
kyoPbpYs2zn9yyntarn0oVp+Ye81jdga1MZHejz5PLC1rtvb270NDOj7CXNwvUFE
kGw3c/lMRODCw5JyjG1apRhsBmNhchT859HE+aqnb2Hji5qO1wYnrdcNnGs1J/su
OiTpx330Te0BYD92YN3Ee8upm9zFSaYddjUwNrbCW2LoyLkP8M3AQPpvPH9iGw5H
nprKS696TFM/sIcDvTEQuqQNX0i6n4NI2o7gJk996o8EEPoq1NW0CwWTsc/TBdGq
lsr7NVAPnWOsIAROpFTIeWJg9GkoQ0bZKoW2W6YzlwKLY7NNt1VogdDP6PnxHqux
rG2l8nuzquGHDFnnL89gJyZ3m095w4+3prby9O18IS4VpiIhrZE0ljK3BYqOp3m3
/cS3dRhnOCeqDMx/3rieYnmILXD0i8QiO5+HDsQ9tnIddgLmoKIm9OkxA9Glunl2
5obdpwFH6lcDxTUZDi1ulNGbIuXQqAvazT7Sc5Z/k+SEp8NHBnVmKYB/vsgdkhAT
+VfremLS+SYpfh/kUdGMnefx6OrxL6jzYZv5clKo1YgYzL3q9yJUzDrW02RvipDN
nwsjqqAPj6JzTiopw0ffxGZ8FQkGFPWkr/wARH1Cy93MqqKw2F8IdtoNocigIDoU
Jl4S8yn5/PRWyIYc6IASJ7TXg5Mg4GFSR2Mi1oDs1v7DmU0fCbnVjRY12KNOaLNg
sdYRiwH9DLcaRfwSq9D5U7qTM6unux8K6nIPbUdB0Nj0p28Lp1DBrzSSwBCHbwR+
eB04g8I7QxO7KAf17PNlIofYDoKgua9YvXqM5GPChH9fSfZfUKHIFAlAuCxUcgtj
5mmgK5dvAr7o3YnryiYHZOZtUoBG3hve+qxLLIaZDYQOpLvxxfLQy1/8W8T8o9/w
8jr6noYVO5U2CNi1oOlAGKM+gEpUpci8Wq28y+r3FfpUvrvwBtw2nsDfi1mKh8gH
+p+fh+bkibFSFxT3fJiC7Pa6EgVirc519tOwHfbmqwClqNo509plq7Z+eo0eANzY
zQN6dz7sWj4Vetb5T5URiLjbCgMCcEwWPiOaboNOgU2rWo4HZz/RCcP1/CLFh8et
zVeRG/A4l0AyeE3Ythq6nXjjaWh6N+WEWF8oxEg5+xV2+l2mQSCrWS7F6qI6ois0
8T6EHLgQX0W9FeCx0O/02Hn8j/wwBJv5VROh5PeEzHTyMO1+J9Pik1VHfWT/L5En
r6SqsFHyWIvO8Nx09T2nRa5sb3Zf5unra3HmoXBKneLkLk/qR/bUvkhPzSKwydQx
bcZTJKwliDzO/E3IzouHio8yC1qkvBGRh7neBdUiMi9tWN+0IYW453pvLJ/+UriD
fNEnG+HjJmoXnppDKLnaopec8421I4YxLf37QHkJVxGAs69lfU20w9WVCd0Bvi5t
5dy27AhVra27FJYL28bRSYQTegUcdIsEiujII/b5eZxwm4ffSh+wtwGF750AiXeE
VahsWKehl2D/9/TX5LWAwUblFFDLft+JI71n7Nilqmwn+gcRoHfnvSD71FCFpw2v
VLosqRBOGmJw8GVVRFbbz+xCV4SpvV3ARlYg4wmZwVqCGJHIolq7Uas9yostLPIo
2xIBrzSXy60cHS2hI9yYDPwdecAs03CHBA0fYhvSfETkYGSu7QW7o4zqp4pyhgxT
EDyvUSbb1eb2acPmVXijXlQoZc3GVsxD4tvcaB11bgZsEREdO2hbQhg5OA0HFVbD
LlcAbNTuZg8UzqQC7i7f3VwgexoLmWBZ94NkL3FguNtcz1WK6U5lbuj6ZHXeGe4h
Uv+oo30RsiAyw1m2/8BfxJMsbvSu6DwvlL7SVV0pRRHUavE595FetRGX5INJl/mF
GP02LaFgKCeAAM3BA2RTGmFeFXxwE3evV0cmnguZuQ2cukoSyQl0AkUoc4UWg+J2
7VqzaZkvK4Ox8FSKaRCimmqeIoZH7uFqA1s6nQRjJpkB1biSPVLC1mqUebMS00Od
ipWctOzskd+qNEkNtMf3q1Al+0+zZaErxciJaBiNp+V8XVz0+RgcYeLAj2F8Ck7n
s5Lq/O3xCupprjIig6Fqr83vIFfmrMWEunhJTTuXiZ6LWvM1xcvFefi1PuRrz1nW
0fAvI9tqyT37PCGD/xDRmOn8P0HWsxiKpT10gkB1aEAQvV4z9y+VFH1rMJoRIn2F
OSmP5NBuyOSqLIBjlxK2brNlzEz9h2RjfdgXuSmy693aKT1wVR02dQHDA/3KrA36
pwba+21mQ//OzQbY2CImAhTTgxmZ68ObPCw4gGVGwezJlFFV1BPWNMH9amtP8epC
Q607QtsbstoX3SqJxnjtsUZ/nNR0EYcGjEeohzer+qcsTu0QrRcXF6qrmETVmS26
7WvXbFoZCfCga59QkYvg8Lub5plnlrBp9vRJDj7aLCJ1tkAK4yQxovfv3mGzxPiM
jnWfLJOyCRDJtnmQjx/t4m+hYNkGg8mNC2j8SM2ezCXawaUN3jGR68YpH9e8YK4O
67wQoLg/KTFloO3DrJbQweGe7RMuB8VMlvOelHhw3t3k1h3dtzZDD28+SF0jP9Ys
kGBJr0IN8PHCU/FLXtHeLQe+7B1Rr7XbNEPVvhXlNWOxCVnncDRfb7HWT6rId9hi
JKJbCobtoB/IAhufoA2UXzjN0d2E126iQcfehBXLt0qw5+6NvLkC2vqOOn+1Rfi2
S/aSg9yWJ5VGyghm1mDyw/Ox1Q62yN++ilxQBnNJGcaEXXxT8JsvFtRwVnWRDoyB
vPdXBWajb3O/sIVKnqvleGujfzw2KOettMC+16DgD3UKULQBGkrCRqgsHBFR4YLK
bfH8Z9Xm7LCHuHkVLNegnE+gwUx7PQwWlXXwh83E8JmG5vw23ZKJIbuqBlgNq0Wn
7Co658RoaNIVzJjQ2lHTUsQIt/9E22QDLr+npj0NN7Yzw8ASnrFMr9urqW1pVXPk
BP7qRBYXqq61sTyn5cAfHQ0VcfphtLx6AwiPACnNbVNXyjpS8rjr7QoQ4X0SrbA1
rIYbpkMPMQgUtFQZX0cOr2E1RmAn+QbfmdNP2mMXinxoDu1XPZ8e1uaLmrQMJWtV
r/enXuazkUNuNHzUZ2FL3C3eFJs9muWvEv8PfuYXfj+a1Gy2xlXXRjIBMs681KeK
zL/jeKXMriu9KFb3ZnlYyvKBtBUgmLheUQG5+QfwFWS6UucJhBLRoY119gqvvO53
+1ZQqX+h4x/2dzeneOcwrQz2lM7/aLxLUk+NYum1JLatyNuI54Kc5JxZxNZoiWbb
tjlVks5Y8a/dFUVYvRxNy/TQhVS2uk8KLhFJplJ0E55dOlYSItlN6coNgpbEWm0x
xweQPlSOXTFV471HHD6M09UWF6QKnGBV2hRKn9Y9m2TZfcUFX3983Zb0hFyfWjNG
3zPI5TUKC4T77IqyI4a90W4YtYy+lvv6DWKEjWDXwCEcu9nKh8B/LiTlhW5/dT4w
CeOzeAQ0C0dkaKINmdmbGZEne+ityMU06f6ExgS5zrz2k/lnBvD0HEAflITJnNIU
4t7k7vKJvot3RyP4yV/oYSLyqHOZ2l1ECGJouFF14W24ddcIHnpSBSZMbBK4Auey
+NLH850m3wX0YZvn2o/M1wWbrhpNYIorRlf9f5pP9QdiXSLMYI7ZVgN2mxGUCmYW
AID9/aEs8aCXj7jhxjz6dy/jttAHbMznbQwTj8w7ayNFYkSoTLsATh86iK8BiL/o
7V4zysGroLSY3w9/Ei8ei7yXfo5vdqTkDhD9DwtXTkxOlIgXBm4SfOKJJ8SeX06E
OCwBas44ixkbvB0MoIpRAvFl2Jm09XM6hFjl26Ak6I/npy5G5hFU/4syFX1OkCx4
BF366AqK+TV8/vsSUXa8g4ZHsBeLe+FTYu9N6lIEjIdsGLDnbflOHsa6uKnRGRP6
lE4y+hybUxlNMasE0UQMwt/D0x2Kz57vrzt+QSb2iuLY3kiZgD1eFNi2se0CsIV/
OgaJCaUWmaEgtCj7XcWd2vhc2uNM5tLLor0o9nmYXF35V637g7Pzg9t2pG1cX2T2
qAD2A0u6+Ash/Hm4E0bITsjTnaNo3i9XolR90idmDGlCqbc/pOQCRPpBKd4OB700
M20wYrNd+GTqy3eDu3kFeDc8shRfETyu7/JhSDVjVUV1Ov4XLOCWv02OlNGezwaX
67hc3ePL/oYomtrQYs/CRZjJvcgaG/umhksPbvxsz0fOzPBlTvqOMQhAoK2EQM46
5/y6B1bcoAA3f/nnu7NnUWYKN3V7DZ1/rakU4TVVt9MVD7PigfnYD4Tg0joH/fPm
kX9DznrUpOTdlonXgrGdSxSujZzM+gpgKrZQko5LieausTAAf3y1F0f9swqZLpxJ
pgSeCSqplgkiPjeE2UUC2zb9EE/dvBgqja7xGV5aE4eRnzKvpEFGQqmqdL1jiM99
NyFhLm8Y9/VnjCXr/2wfsZzVJ/zhTnnrjs39gWbP0Y4rjvjPMYspLFTBTud6ipOp
xJ1RM6vmroNMJUjRVD9ljWIFftd7H8HQtF8Tgwc9blvYDAAXPjCrGWb52ylgpmWK
t1MwuVNYV4QB7VyI+9JSukubtByyX2HOT3bOn/K8P4sJk8j1+BFZjQeBpfUQFt3u
U+wdqGKTphYJSudvf9akBbPPFYiRfbfuW2Dn2UKqivVerQXX4xn868b15djC+AeV
KomB9BER40FKjkMiJqgI/Spc6crqqJ30KFqzkr8h6B0RUTKWlBpwbrtf9Vy+61gH
qXxeSMRQmIhGLDEy88hqfg+x6pZXWmjC+33LNVv7bfOzYzzXinW1nRSK5ib2RnFU
3Fnq3ZyNxiqmPg4HW+VSBZkLoRvexKWcm3J+0JBHEthdrXJtWMIhfSXpoapotNnT
XtdcMZuA7h5nqi/4QqCM4cu4eV+IoiAwRZ5F1IK238h5K/JKNaMLG5l157TNA6Ha
rmy0VRJCFqEgV6CD5c/2Md2c0WhYQsI9B+iLoyP/+aTbES9KlUcVbdQ6hi/+/OEQ
j4RAb3PEQcZUeuhUqQbYsKslEjnK3M9uKkiuTRS1Whlq8dJNhnkUeE4LiXAH6cc3
hKrwxIAYxkLKrKF/fhLcmfyX0HPQc3ihv0UyStFtjVkfuDCIhFWb98PK6j1OMNBX
ACSTT5rYmrQwJA8Q/SxjJA+tx5ReX5pnZeDRNxYKbpwWeYLYtDMTIBOB5z7mIC72
B8eioJYNI1WT6zSMsM3QnTaU7d9ezBJru+9lpZM2LFEfCjUEJyTFc5Z+APwUz+vl
h6qivnv+B3WEDhhQRut5Y/cAMWIzWvYawkxqHXkpGdZ8Qtit6+MoGDopUE4I5Xgi
Tdgv3r5QLvbTt2tvm4Emi+nWVsq8Gaw7DCCZd74/Jidmk3Dy7E5CKC6A3fQZ+ek3
QEuQdusdBA6bo9o81chfNyPeknJQhXJGQi7cqkDKw53wv6c1+bDymZ8AZ2EEdEAc
nV+rifV7WD2G0tgJc0FPMbcgAZUAQnTmeiBh9nDiMM9yRezkqZxWN1M34h54kzsY
UU/rw6XjdFhnzmE5cdWCfbcE9cQywBbv1WzExHuj2IVxBNJU6B2JSMXGXZaY8FQw
yCxE//R0CHGDTAt58/towYtHBATbQQKwYEZRnngKpm548ngOe4TWc8USG4i+IsjM
khhuaZmR0X0iFvkjl6uunem+T14RPVXIP7g6GAudVuE9l7v5zgX28rQcKrICHZcM
RQoSwTFHeHInDY6LOhoiCqQLH94ujln4PeQTcMJw1cL5v1gANRzekKQ8aers3YbL
+3aLDsVnCLNNPCiyGGlRHheLLuSiVc1lslHJefoBhyVhGGn0pv9zkFi/2mNSHYRX
7YyxFKNR41rFz0R6mlBMHZ9ZxasEPAGladN/mMqnaxuSgCCbgSo8X4VYWQfJYeq0
Rnl+dGzj+VhSyMCnGJEQ3CF2ArM2cpfsIMQf7bqkTf/PugQdJ9DwdA48G/Itzh2W
ekS3mVnRZv8PD3+oZnyoQLTylN7XHozFjUyzoST/FrAkVkjkwll37xmdaObatv7N
jwdoedriytFsNx5r1tEUXfc/fuYfiZhyaf2xHKTEXVUdonUu+tgBPxlA66DNoz3u
Fr5zxYsgqTuAAnm0AqUdRr134WtLXwZOKTJQ/G+R0PxsuWtqUDOjiDDmssg3Qrwp
CRE2buBg/e/oqWFN2CA+FMdeYsOtqzYOAPcpwGYd8/2MIXJ9gIPnzgbkdkTl5SaH
cQ1DXaoX4SrkgUR6VRcLCE/ixpUuHVeuLqr3IhLwIWQV9q1637ZhTwIgYPkT1aOs
OosfRmkMNDNhs9y2JR7VLi4Xfj9ggxl3fR2hj93uiBtTTCfvyIX2cM9+e0+a2GHz
P6PBK/CBgVvMDvB5ZA5tZUozBmDbeUcZ0TTpmJiJTv5MPP1mJ8LAEkPbHclkV1dY
88ymXgT2PwPYWstRY9HGJJCFzoxTGeIUcKCYxt5Iqp++V3GkVPyRvD6QAfwVoRIZ
eORIwI/d9M/TrD8KiDe5ioeLNwzFzAwaJNrVwP/cAjR56JdY5XmN7Gq8bLbmOVdH
gR0KJwbHY4SVGnT9uLey/ezwS6vyNMCA7RnmBuZ44XaLt2lTDMEoFCE51+GSGo7Q
vhks5lCE+KGokCThP0aOd7BZHE+GejZyQ66d2xDIFQxErgdhkIKjL7VPaHUgFJqy
XPCfA7HTEh8uEGFrhCCha7rS25s2btEq9T0ciJe2guRDg+rsW2eGABIYEU2BGAEO
qlcJlvPQsjJ+7Zx2zvKBaTuq+ibfgDA7hyrySU5xTl1m5yClrzhf79y9SgE6q80D
Nrjy1dHmYJaMvPyzHO7wy/8B6Q7b++ebKp17OrUxcXXz7JRQy3acoOKApprH0hQD
SAYE45VjyQbTCn8kt/JZSdK9n1a8/Ug6reGMQZuCscGH07SlCarhAmpYPk1C8nHB
F6o4/fBI+OksTejMnCm8I1T1Y2B+o1wRsLwwFdYs1c9s2gUNX/sKbSCdjuPVIzf9
3Ly71V+dGwHno/1tt8P5GNOjKQVEN14Jh597QmYGGfNDalGyqKtujABoLBUaj0EP
Z+F+Hnw9FTeDJ7tt7IuVpKSwv1m0BFkCTc3YZ7+jF068PhkD9MVvk1QoT8djs39Y
bJYGJZ0zpr/NNGok6YxshphCd0MlgBf8Wdwq8/9vBeWKmz6CKKi0lYHyZvbzVQM9
QBMe/emohZiPVxzwn/ZW7iOLgRL0WnmTCF2tlXHY4Ca8A+M3IWSpGWYHByteLo/a
sBjCKe6dK/TybRpXmJgP/gYT1kS0BP2YKm4UXxGyc3cedE7lJqzlKJ0iKApsQ3lD
5lnbCxlaCY1C4nxVTYpwMpN1sMLKwjlkSMiGyu0XY8N/l4oamILoRdRdezmzwhop
pyUJrHivpRkln28Ts1EyjKJb2TGxDcGAe4GVrt99NhKA8nXJOnRcm3xw59IS70vi
FWDNt65EghPl06YJZLXu2QPxqtHs2MNi2BMBZz+wPJarl7hJ1dudiRfiC5fxbUAb
lYgGbdqtxlF/+Lyyg2xyhqMbbe0mSSiJZrstZE8E+24tTGteEwFqpSGwG1hFmq8u
d6m3CQ7iljD44p1f3Fti0qRceWOUfRCN+cT8dHCOExmTWjjrTR1ww10WobHbDVta
0Eq2Yvs5+LnnUpJLQDmpIvVJvSR/y7R4sY7fRsunhPDMEOM2lqfIcfZyTlWMCwZz
pacVGPp4xqkPgPFFRFeSQufLCUIpLKeD0OZ+iPOVzyuo0uW20gzVo83wVKjlSzEV
+ywktImSQlGNlLM0eRcjVcwkHupLxWCSgdrVwVH4YRrHRS/ILNSnJ86npOVck96p
nWybKYYoIwIbjATu/x39kCVg8X2xTfws5kGsW1S1XvYtxU9v7knSDY9WfDd9/Oqh
zMtUlApqcI/fytHRYBVDXlBaTE0ecVi2IBUHPR+DRusS0f6cXYDjJpjayRAbVOC8
BZv52TLkY5t+zMBA/ARCFLMhba5DajJJpnjVPwItTkHWuMAW95iHf1ETE/nhAtN1
K2uDAun3l4wqezbNhDakHQuRzqFqykA/0xrvEncBpnsbtfnFRd2/OnnmIvTlDhEB
w5N7hmE8CPR3yPF8z9HbFP0wRz4VITjJtvQs6fNud0bpPOzjg2OYXu+JhSte5Y3+
MF7ZwptGEG9zM2y6IlPGjyA9xQR3EptjLf6160RDVY7b1GN0lAIm7k16MZu7gn6N
PUzhx14fl2teGIq//PYzQYkMEAMD9M1cAyeHVRPaTpf3xBBGAE66MQYGr/IyIx24
drbqKpBkucbZymWu0nuO+6RgcmV68FxjbVeisfG7G7mDSixYELBmX3Ot2kRvGCsp
U6/n78i5M9PVzid5OhdHOgjgHFpROBuCKqqFbhuP5P3ZUKKWjIn1hXbQjLv7HtAG
Rc0IYM4zc4KGlEF99Ia3AQrDAR2klL+8x5bdJHhMnWDhtlw15rG1y+ASfVGibLTO
4lKjwunmeHlDgvlUqiEiO14W7+vD6FNntNxmLL2BKKbjf1GKR6prazm5n5tOWkIW
CPszR9iq2cViaa36JVHm7Y95MMCnZpEtYDrGdW/MSuJcQfFn9nfk4FAa/VI6n8qP
V7Ya5LGs6x7sbsXpRJva+8w5Bp/HYnU0NosFeks0wZfKCREfEHQE4P/n/AR0tQYp
qVKRqMq8LoxaUw94xt/MtObSFE5SPaF9MJz2l99f+v3HjtKPHMAuAtlApZ//lc7J
Mfvaofk8sacv/VyM2PcfJ2gb/TZ680Ii5zjo4AuXX8ZDlEIXkaqFa2XgfpkJF2oN
ASmeTvqlBnmUJcgP66duRGODGX+uoqdx6MrEhNg78uANNDxDhE962hzljkDb5ars
VV5/O2EZvswtsymq7iKolNmUn5SksRwgcdRLU1ysf3M91oUXd93J3I74yi56Fc8F
bbC3Gtc2LhWs63T48+KS1Z1XtR0xmuimkLGtwZCvEsknOIr1DUU667T/ReGRYLVC
8is3mFlBhsvEXMI6n1Tr23zEE0ctFn9ujW2YDerRlIZhk1jelQNg5zQbYP8SXYe7
Qm3NEzdmtLDT4ODVgcmE0LSMLFNQbY1aLYaegzMMAyBGfeo6IjKXGNoIj5RuWUaq
su1VP7U8b4UV9k80NnV64VSR3ul9X10QpWUOw0Oro+V2Hk9CQehQ7ZUPT8FReqNV
H5CWciCtJZDAHjWdSeyPOxykPdRkonTZE46a0TsmiT62qBH8sCH3dG+xL7kGktmK
wlxtBcL8WG6mYKlKp/d6aH+xG/nIec4yjl/18KJAzVMiKH3Iwc6/ICBAjNqlLKol
7Vxe4zSMds66IyoeDqcin2yAjn3v7ec8vCKTIE2gfqrnMYc5jCpU5/YvtKQa9U++
Hwnf4a5vheGcEcaUD/vz/sfS4XQ08IY/de/3kjBfEbOlKtP1vKz5I4w3Xpy9Fm3v
7c75ZYo8h9H/37PHX+kblYNPAmC7h1ZdhlGFpGC+hcN+IG9Tj9tCDnwaszrQJe5L
W6nNMP78e80GODCYmUauLmtl6HzxszMZxssDwD0ZDeDCBkYGcHUlfszCQuJ/LIOq
dAaof64kcdzAquUoK346fELA9oA4eMKjnVugv6WxdGUfdfw0nNBO7CPO2tthqQV7
XwLGQQaNMjDEF3F6qup5Kb17fCCniM7E6zhk+ar0VhLlUmO/dBR6fHTNLKj0H/W5
5GgpXfcfzAfQy1Uu7/mKhUMz1MtzMs6QIlLItZ9kU2u+10b/DOWWoHOKXjTvJ9V9
ZZZKaGPAMsxC0UjS6/pFUt5rZiYPSN8fnuZEarQvOrnxZp3fLagxLvf0ayiBj0uO
yMiUdyJDSEbPrza9Vx/VoweFuZnsB9uVGdhxsxudaLHPxVLbFaz4W6xA9GS09jmn
pVjOveae5SM1NeEy9uzxIUU4UBqXc+B0OPAoFC9QKjFOpzT7qksbM6bFmBXOcIzk
bJ4neH6p+86UR/am0B8/0e8sTV80FeoH3OgWGVNn1mB3s7lxNiXdbzVQBVhp7ZjK
C/pSSHC5951NWY0yTbVL7BvCwUqPhtwzV7m2sZ1xuvELCY0kzwuRGy73kWFA0hm1
BAyOdrP4KZ4wQQbwuVuQW3I9zOIuabj3Pc8zcnog42jKs5fxNseAqj7Rez2xGckA
KSy41CalLjp+g3w9C2/NoG0VNrHvaGtDiqg7Z0IFgzeAnf7IoB50/2/MKjrY67iE
vYLAijIJHZAihwb6Ql8G0Res1LgGSQ14x5vPP1U8EDI/C+uh1MUOgTrCF9T1umo4
gJjSyjVVJ3AeQGZ0oi114+nOG9UKy/vILx1uY+ODj1PTCeZBPATTtjmRGvTBZ+D0
Pr0AImuy0dZiwTPGmwg4gpAEPgcC66FRrkUvh6zpA4sba7+AXQBgM5R3gGrpXfY9
WSX3m0rRGFpz4TyjhpQTGIz77a2NmutHfNfvoI79TIs/zDgaVw6B5bt2u/ZdGci8
o0OW4/ClBtDx45/bS8v8FU3bCu/QnmZAXB8i8yxv2MrKjZiYq3hgvBD9KIzXfLMe
BpgQ3dT53gPvGr8uPEBg4qN/REX1J+YnoYpuCyx3lXZtyqEk3UJMEVUFSkjH4pAS
TaEWh3j0IbSQOUxr+nCIZugJSUDy9WErhMmpGvE1vwUsFbdPRFsx/l5wxPTGjyfp
/1sp5tTydCgb3Z8U10GfUwDh4xhwqlSXVWaBmqm1mWlNkY0+am/UveH1bkbADtgT
THvjzPjWLTZDd9V2ctxQXrGNZApLuVd0GV3FlmU6Gz+fdn6Bw2/nQZn4s00jX/oy
E7vWhrr9d7C2y2hae3n9FVU7QMM/KPSJG3zFKCyzemo0fiqvmFLPetxC49pPRuH1
enp9Y5z3UZOQJlps/pph3QTaBzyl0p5udq3cMHVETgSqtSoM4USlNslCimeDRdnm
UVBFnJRqze8u2YtjWLkMCpIwY3NpEjTJplx+SXbmwJo84E9xz3wWeNrsZ51k9OI1
2cuZnCEmr3fuvipQyeoquP3IoSjiD1yi0c91WulucaKIiaYc6nh1YoStAPoY0DH4
+4vFgi4Uzt5yJAwjJesnml+QAyAwLN1dM6jlyoktr7KmtsfAphE6zIN4p1wG+toC
PvRiv5+mZ8IykTFeJONarMyb1mAqd3STolQr8E7acvX0He6gaeX9B5wbe9oQwuri
vsR9ezpyf456FQoxsof9BAhhr6MoITdXwGLxuIN/+1JEfwabMaWdvKIUx0Cw0n0D
k4AwHyHVZEMlfq/8j0mzV2Yt4PB6eL6lBmkBSCb3lzbI/O+8ltoyFH+6V8r0vDiI
Os8EK5fzIvxNhk0QWP1NphTQtWVpnNe1najNXiH4vL29nIpnqF4C6+Ndj41gACv8
wBDUCVPkQVQGXqAm9Qo9Zh0oB4wZqDx0PiEiymmzuSAk1cbo588lN7hQZWNINEZu
ortH+9cz9kXvoAFhgFvrkYi8umnDIJYy7APpLZj5rIF9ac2FWm1cSXSuQqzdvEfE
Cj+olqQPG1qS6jzSm2apG5ZbSIIvXa60DR+sHxYMS5b+nrbbZQw2quXn1iSCtwW3
q58Hd5gkeRA9Xe4Lye3rgJxTFD3MIIjAtjDCg8XLFp0MuqheFqRHI93+rcItPdHT
9Lnyv3jG7d1BYff+D85bDYjFjBXMyNzCDjZrnuGiw6NI+J44vKoMh+A7BHcczMKq
SZIeFF+JLvV9SSM9Hf1FVi9GKV2k9LPphCJG/L1BBFgOump6NxY6SIGLXZAVYEGx
0SdU0ypNoqlwbQLW0qDeY1lShVyJAAs9La7CSRjB3bs/HhYuMpHU2z6YYZdz9zc1
9GCvXK6J7s0b1SLjjhx6MF9rF9xkBY0ahGGnSE7uFWt28ScXuhyKYCrHWAs/2KBl
am5Msko+/3jLd/Ii/zT0p4LHZlhUUK2GkX08V8XblB6iccsp4ShNc5MH0CN4VCtv
NP1OxxGefMbJtEWWpdsmC/A1rTVvbyTKL8lqy5YDfCqtH3sCYL3d34JXdmRiBUXq
8I5bhoWDlBvU1eaYKakucD+DDCyEv/dzD8kl2OBpwMxddKH4UVDVFWGFa7k8gsWG
xxuokQscfDtbYcydddHboQAJxZErDkr/YaucwTDIIrbBK0Nj5dDWl/0CN+atR6Dg
BkH+ELoeRhMam3HLckGm0UuhuIckZdKJwAzJf0FPzEK9XmoorfF1lDI4ippME7mS
dmQXkBMoE3xEPUIwRyIXtqOnEhku3/Dh1Ljek7WgbdUEQsmlbz5UGvhdZRa4CW/P
AEKNEZ6IgWkCse+uSDga0pmzQpf+x1zAnnBozkEngajW6jHZscwlQiEIqO1pnF57
N+grXw54XaDTaSHse93fx0nOav5q6xyYKg0gfecm0VeVwB5RXJzO8jytxzO3TEyb
H2jsXv5+6Gw5oakLsNGMvTCYr+WcqVdG5fF0RJgZzzbBsfpKKh8/2FDOx2TH8JOP
zgD6sIHpnqeaRP8vrYCIPMM0ehgPHMaJxqQ1JF//xbNL1YeKVVjgudcGVSFUNBct
FKAEgR6SYcTvxy97Ob1vup9GxtaT7dhEP/F+m8lLc2b0RJGS7CKQDcjoN+xxYikW
OEKFMUR/74rrmp+tKg3zcDmS3en0mAepqclqwsSEeJARFaHSgoY8Ju2thJidqcIL
APqu3uoUy3oCB4Qq4gkV3t7OxMeFu5uu8OM3TtWKQv6Qpuvb9Yv/jI/PtthHppC0
f3DAi2F8wWEXYTFZGfqZjg2b7pKmk5+Yj+lkbttQ3ze5ZMOKGda0FsypnegEW4cg
6s1rS4paB/1tpVm6Zx0qkGRu7XHFSMmL4FPG3fk4QTiTCZG3XSVuVZKIBe5fVN73
Nv5yVMpW38tecihzj+HCwcU24xhuJYvGshmKPuC7VzM1XSb7+JyrTJ0qoRWE7VXA
YRjIZF5tf5fFLkMOZBaFXUlBbQJD8OzR6X3dqON0baYeUQgNT3xhjrbauWDT60i9
5WKbc3eYFQGuHF2/8QhOt+KjTK5GxlJIciOkcEbalG708Grf+fnk6yB4UJE1yfle
Jlhq1vE8KIfZq/EVA5GIiDReA6cN69owseLUGWJ6zJomKSzIQXoZ8GIwvffKfOyy
KY7uQBbPqIQUcMPkNddGwVJyhmeS/hdwI/MnGahsNLmz5c4cBWtN591fg2ZeelEG
ixTQ8qHb85/Kj68W/OV2yTOgBgBoeaFPCV99LHET4/Y4Hm/uGz+XpW/+Gu/gNq6Q
HegI6Z14mIRQDWN4mn+S0X1lpVWOEvgv6S1eztGm0mGcU/BuiaXAnAr1wqtHZoCm
ckLOe4c5q/sPoOm79vzNGTu92VbW0a1mlEHHpvtKmERn3Bh3XCXiqj1giX73MjNW
roATMFKFdktcZfILmn/uKSA1HLSG0Ep8ZKzShvAlVDD0cWMud3PTxeP/mWgB7mP3
fucblQaXaa9S2sucA84Jn8Oo4sg8gOKtykR/bWqyNHeFwX40/WPh5v5cDoGNn7uS
rKRr1RL62dJPVteTCnaMInhBd0LqdLGHXeYVrWwStIAIjpjnqhBVpwu8A1nipFln
/EKLq0IfeYalX503mGI+4WHIAKzFIEzFM5Rf7Bjozmd9jKk1EK9YGciEz91kkcXW
2/RGqiL8lAuhw7F2+y3olHRGtks4IXgyidUdXhw+87lMSeX7YGZ8sgsSqxvEJzX1
IVKiAnfHOJpFTTjFT7033nO3+Rp2wQm+FURPcd+8OxXsxFbAHUrMV5ls8xT4HrWW
lzfNIC6vOGBXp/4w5DAtwjEzGlOTOYCB1dm61tWlOuXv6y3lKc6QDmdugB5ZQImO
sPWvCzzyZSozAWytsGOkhMoz02Z21Olf9oyKcbX6imubKXNQVOzv3BhobUg36B6h
XDdqjFdaZ/zC4f7wmEK8xOfxOHr4tu/dQAN8LQzAOcSNLFyvJMzFHgN+i5ehvRFt
cv3jDsHC0SgTd6VLsX9qDFikITPYoZ95zFcD96d+IgzgQmTtmescdGM797Io6lUz
N2EmWHohqulrMNBHsOAzpqU2Nr/EEKzN5uaEzkt2oe4lFcu3kibj0ZgVJBYIwKuX
L6uieC2I0RtFDmhbY6kW4ilyIQmGXcNimA8nO19/2//aEBDGtg2z4h/yEK7buNIM
d+uHbL5Cjyd7Dq/7Vgh0hfX6UbUj5NKEnSczDET5IPArI/VqbLM5UThvR2cPu9DK
Lng2hEigbXsiUirXwLTmxIsgoBirUkNrhHbrVWuSswJuTMnByLofWojlo9D4EoJg
SX1k0YXQ7GhRdA9zFK9uyqnk8zcVe2nxKTpfxmrySqArKwFHPrJraeW5fT9X/Lkk
D0x5pVmdWAo9WUTnenqRL0okgJzAoXzEulp9b6lKMe5tOAFYYBBkur7ApGGE5cfj
+uI++ysFd40/7HslyHFDDIy0n/d4rk6wB+mTSv4tuEcNXicWGsfia6tW6wL8jROh
gZ8ziy+33RNmxNQiMBvwlqgnOvZQKwdhp2gVglJa8V3gyGChX+JR2ETnHkF6L+1X
IQcFIcdoWGPZzKr5tLYuYFsPb4e52Jj4WpDfxNPBTW4uBCG61wvpgDAknZ7hrHpE
J+DT7k8IFvfrgEF39GelUf4CrrMl80J8D294/nbaeDS7PLyrbKIoUiG95NZyxjfA
CwTJkYP0tkRB94bcCGXJiBXULheqQovCEs9DXw4Ak29AyA3nb8+WsgP+j6kZb9h9
HI1muW39ix6RHeVdzPKvm7ODo/Oi+w6orm4Dnpcn05mb1pQYKX+prJupLPT2UXD1
FV66QFsypESbLbW3poydGmNJxnkCZvWCOXa8+G11zzvz/4o1wkhZzANiU0y/sHtw
AUrm6UfSoAuHYyEeB5fqjGOMYSkG/YPhrDm+WjK+/pQ1OYqFtTuznCmYRWyWayBS
vAGCbOwawI9dR5AEoLvOAf7DOz0+pia3tj47TLYe7YkpPx86fDSsLhh+SZXFZw9Y
7NT/+tKY6imfvRB9kAcwImNFwkLckPS17WCBcKHPtkzfFGMNPVLku4AI9Q1JZ6pz
+uSm6izQd221o9x2zfEuUkbG8t3OrmHfmPgVjceK7/fiIAze1mBAWLhQGA99vrm0
whGYBDfTScNt2upMkagmFq+oPEhZjtYnHDwSFeUe0SL0UM1GpJV4RMa3dCuV06XN
6olyGU+eoA+Nh4xPn70+oL2esyUmXw3rogjBd3WUFEnRAmXggpheKsT8GxD6QCdp
teols+RlcP/ZkorDxjOnUCq66n2F7+rnlEyhYylKBsoIH3L7qMdieHQa/cJmF8Cm
YTG1lBjTntKl4EOisnJSCawErKa6Ts3fynoHWwyDyO7mbM7ner58Oh5IThQ9jzGI
d5JKMp0j3LcKolvEGFt6Oe5eQCQsIhJ0wy8Amw8uQmAkeg/RTZAOYyjCISY52Ofv
W2k9iNVoILE2DMeKWfgh9HNYTH54uD+98FANYBEGNe3K8TVfomVgOP08xf7JvToY
ijhgAcA4/dXCJELMoHx8lLsvHkIyX8n3sZzNQ7/2YQbJWL7moNMQ3xkIT7m45Ccn
XtIcR0BfZmJBnxEMI8G4CNkF8Fhw2pWyVNS0TzvNAEOZ0zPR/IorfHGy0HWG1BY1
GyIW9vJVq+WlidLDs8wXWk92YkawCR9lup99OpV4XrCBcYprtdYufcE9o7QvD30I
/+i++YmTp3QmmntOeuw793XPdO91c4pZkoxYArGLVtGkJSwI40wed1Me0bswe5Jv
SYfYM+YI5U4lK9QjF8OaqMQnq6Q9LxQaoMiuRs48jXdPZOEUS3/qYyuxCl1/KdxQ
2EZAC5qiKwtfJGiWvTpWVbgWdqaedf2xRShR23jdlZi/JJHP4Hy2dEGYGhLVFEf5
SgZJ7XigiSp/3mNiVeEx89JchKOObO5f+w9fmcGVwWCKgYerdAwe6hQfGg5UDL20
K5kKqJccwMrsEyFF2JihU1jZFVeRfnlOTAmn7ODgN/d+gfQkJ/pcyGmJNNAnesFc
HHx12IjQFnnY4hVDVfrceDnnJlbl/b+nSXNfNzS6WgsQ2gLygo4bUPtRuGwM7/Vo
l8OHysbd1g/4gMBS1SwROluxY9vbLhjTWiw9MZhtRQBiz6vyCvS6Y/YhQP3NZrsg
Bdzju3tlnH4C3dk0pBE6h3GDnWV3KN+4XCmhCm/jNzsy2s0Miia4aqCWtTaFkIP3
CAcWhcWYBiCJnQ2m68Oit4pheeCjoi30vWOZLpp76+cDUqcsPahpuV4rHbJImZ/a
hQvYGRaYd8jsLV9oRpjQpHuoPVT/zO63IA9mI0E3rGuLnpD7Jc86bDRbgFnNGTtE
EzzHBJFPljUn4Y1YVlWqotsuBT8IovzWAwEqqxsSy9C+nnogEVtSCGtwzQmcgcql
iHaw6plV0cnr2F3ZAONJDznCU0RgH7NVcmd9gkhdMxmDaytHMpENEfNm7Schv+fh
OSTFKRVI+OrJj6E/0GxbKp9DfOa8waLbxUMv6MiZqTedwD/OFd49GLh63b8kNLSM
VmBEQui0RcaCxLkMXs9i91/BYunNUefTB+Z8ruKdN1s+22e4v9HzLLK0BWSyXeer
COjwFZt37eGPPdicjP1VvQi04cIZWBOH66UW133JzJxN8TnhghVu49TaCfDEtJmQ
nd/9krSiMursIeMUWROAtbTfc03oFtL+Qr7HojDnZB2/HlCTqfJVON1uZhJLulzc
WAvpyU38Dfj/cxf8Yj4/kP7Gbtma/xOr6J0hMp3i60oBgrI8jlLS2SM9jUgFKj19
1/q26Wo4EC2pW4/nfKYEmdr6kVfcah2FvQfU19EY/XAEEXvtYGWRrfNgsjQ+Iv0w
kl2louDZNUgRLMByOfecWXY14EmmYkqkdVDUSWHZglmUuzqxSNYXkJXHKx042EER
kcRQKCaSfhbOHptAWQS/sVoAJtwTi+onOHlLYLcNv8Tk/WvI1W/hbKy9Me9fKU3h
lMGMf4tKXL0716Lj63w3+DWkgPksU+jI6R+R8ZAU4Nhyg355SyhOtbxQcu2bFoL7
9/L3ELma+8tr7i1c9/figK4CwC+zEThsbL9/OEFd0o/5+fJeGrZk3jHLhlOyr7Yw
U9aKTYX7ZRAdyUvxqgp+LfOqh0ZIb4BINT0FRcFmenWP/XKNDQo+gnDK3MKH1gqK
g03QIEvnfpyNjYsspZjzeGUzGH84QYCbwFqMlkfIv2/3kx8pFLTsNrFi8A010wlJ
M+yfB7srCDJ40uXV3YZZSGLNVx5zysT/3uErhwtpIQZCS1Uqbgx9UTyZju6GMRpg
Lqkw3gIGsegFxj56KFWHSP4zeyQVWofGpYyy3zNZG7+rn5HZ/4skOmzcq0NYUOdU
1ru5iozKwlqSG6hMANKA2chjzEENqLm4dtM15JER5XO63Iyw0F8X0tRQgnVdjY/I
6DgGuR2fAKz7uwAez4zBO2PuDj/3C75L7olMn2AXsKAifLOr/OmnQlcDQL9eufdS
q8kqQIDYBEs6fWwuVaLe4Gh7ImGCU0WjxhtEV/LlohbbXxMcFtKK3yi/4a356CVG
mhD9sAGApBjVjTzGAPfEDMSYoSB+lcbacEaBM+Y0X/YXttYXDiucYiqEa4Xr6Kzi
UWfEKlHDFHUCUWx/ai+14aZapnVrzc97sdPboT3ovBmhEQjo/ZtgTkXWB823SCqv
zczhFbngOJsJbvI1ImihEOXWK0J+xl9Dn6CqcipIhLjhg4LEZ6ZJSFiA0IrLfT79
yP6Epow1AtSosOWm6vmP12d8FXJZlp0/LeHJS8+kA/NUcExSrn20SnkrPeqce70N
+kfxYYrSA6Ox/XTEgCRwZqVo01ALqjsXSP/1Yw9BWo1DLBLgtTGs5+FxviRdq9/C
EEOtVTXMBYIQnHakwz22rcmABZ/3FUiK6iZjLvAt3x88zTluaGMb5G83FDHb6tDb
msuCYLoEZUZHy0I0k/7/OJD+XS3Mf33R+84EEeS7HcVvP/QKl+NTraMQAvcPKdSU
BhShBK6Ey5oD7eaAL/rtgOYSEMFkjyVxHL8VFFoPARIVhab4kZfbolR2BYwba/Xm
UuCixMor5jCarU0VXdC+oGwzZO6WuI2mWkM1ukeKkjgK7Br8Rrplpye0ubL3KMOq
VL+r+tyBVuFM9Bv86RMOQ7OPHXDeeSRB3EpEN6oIvlHtT3bQie5YEXwsrVdrx7PY
+StUqpAtIai70fHOOMd2A2MquDhTQHZrKwnwquODjpN6azch6UZ6FC1VRXh/MA55
57BoXU3rFt0EQvU+NHollK+MweiDrrBcmbMj+Ke9iUldnWoEWodUQFhl8M7xaZ6P
wwY6dTsCEO9x2UUJoK/V/enNlF1NivOimFmZYqbewiD0biTyiBA6hATTrU6pyMDt
+ByofdnDarYWFnulT63TjoBMX56CRxDkcCYo/f7r5ATgoxWmT84LjEV2RIOjTPVb
YJATj2gKA2G/yYOF/uqcYpWfocxJ2kxnyhQmj2X+aW2jYFMD7Cutn9RLPOuVJv99
f1roh/tFjYlg0IO1AIReZ3FI2X/PEE4NjflDTcK8a/tiunw+5GeqkrOd6qOj6Ynb
z1trLT6hF6Q1Em11jND7hyU5qfI/BRjHxe/RPz3RdFldeXRQGMA4tKS/vtGLQae7
WkkAcprgOcDB7XBmrXLwYHogddvbnUS2vjQbl3isp8lXpK9Gm8IcAxsNFfJUPIwT
MsNNR34mvHhj+eymrCPrEXxGAoSYSfwg//GUSCE95K8NCp0sEGJFvZwp/d7rC+TQ
3UPzXOU1PdbjOQBLPULoJSoRqWRnMxATO9D+NiVt36kgKkMsopkVRNSkNVoNTnCo
JtjJRPwWUS+Qgsx35jjOOzXnZdw7pSnCj3xl6sHL9wE3Oz4F0kxtremSgPzRtpOA
ltfpfGVZMGSM+Glwb1JPZP8PZlzHzaKHuvUDyJSqXCqRytdt0ic0NYW0hA4D3Nes
ndQ5epNmzQkeKqI8XuAggVadvJnIdG00jNZW16fGNtgyh44cfWroTgZaxTheb3OI
P5IfXSfPtp1WnqT6T015Y1Bpxrw/GpigbUT3ECIS+QMXhxasrH+6VhRtXhoRqjDZ
wxgZgEDVOVLecB4tEDyQ7bH8QnKRG+KAT+SMAxE1AGU2N6zbxG6W94Q2PIq5ptr/
Isp+1NqfSXnhxdm1VbBL+aOEew1VpEHveUIdNV3efTknXyUzRFscqWQeRJLZ8zl3
HISXtSLg+wM4O+6/3fES9HHSjZlthPQHx3Y2MZGzFdaYJLoHBMSLBIqHVzRHvFwd
r7wPDMK94rOQjmSi/wG7/afFetQvKeX/u+wUTuYg/9a2Wv4xmrAr1+9DMrSeYpVP
8hTXYkHCEH+i3XcDVqxxK6n3kbjGG/+UpBLvpNjTVAP85Bp6u5kZ7Rz/NxsaZiaQ
STtzfoZWN7RXO37PQ9z/dBOFkuRXs7sQ2cGpWzuwZfhHrOiO6t9DvF/8dILRxiJ1
fBUnun4aBdT64m4DtkktbrVW0GzIepwrAv01c+hzx1UzPSokWxQzkSFkN3X69b/R
uIJoN+Dj1ptNXUTHAYJGxAy2fhNWMesFqU0RkbEPbqGrKHke1LEItTXsuaIM46Fb
Aj0s8eeSAjTwh+1aSfv12oaQunfwqiQPLeUoZPmkJwQTZEnmPSFvEw3dsNjVnzqj
I7OsTzlHL5eEJK3PGg3Hd5UBYMMWlBR4Wqkn5rLXSkCpdQZsQWEKRXlmqGYxYJ74
7oSetbQxpodPA2Po5IB7Kfr1Hewu8d+aR8wgvJ8raFHIE6CMmOdFKIh/pGz1cYKf
dDICMxTUZBk4gNdCoxAesSBPOByvjoC61cfXuYA5uRFDx/yyvMHdUeNQpolf/eAF
UXxHlk7sKPfgScBKbelw8Hx/xiRppisMJv8RYks+i8t+p6QMjcxJKeuPF0I39AhK
f+7M2DERC5JIA033c3hGta1juu8K3X9uINul44V0RnAvkB3mfjsKd3v9H4md75oI
OLJI8jqKxsF28zINxI0TSQbYhdpQRKf2YSQuK+2aXzJO/7fjldr6mTRQUA8qOW6j
7yTVMpX0s3uneztnAW9dG4JxRy7aGgvQ16Gh7HZVaylfV8SVKJMMSEu0JF9CVWbx
a3eC1cT4A1RkWsrKK0r5vewLNpNBVTbej6311lAgpaHt9sUL1+9I/Jd+wgvQeHzZ
3TSkeQeJ9/VzXpzjH4XWaWvVVZdk/Zo8UELRAV2u0XEwA5xua1QAF89B8UVCXSQL
Xzwy+rami9HBXF1HqC4xRJ1TKCvaJW0J8s1PDBHrRh0JMztSiLvBZhdZ7vMHyJJf
tw5iiJ8D2dJo9dMbY7HcifXmLbvDH+67yy93nXOv2/EaJSmATTtp27UgC0mSiPUY
8akiLEf8+wyx9lM10JtuBHa5oa3ivr7EbHlGcc3qDk0VNBi5bJkxA4Oz+9rY2TyL
bPtId6cSu4DprS75Ihe+IkFvW9jg825NYfphpnrvdMlMYTGKH9dqd9gyQdLo3Z7a
14JVZ+rJMPD2sD07sxulpRQEgo9zXFqfOx65T5Nm1+ngXmrtLsEaNCz2YHzHCYAC
wJPeJYegjCiBPEV+hta4IqmXjYOZarjLj+QXR/L4Nqm5QCPA6UMOfBKVcB3q+ynm
AHDKIZVhfO57Vdd7e2zoTOFfFSLQC5MwLw+aNqwQM6MNnrb6NG40tGn02wFS3RpD
4xzDfF0qSFrBfNoIm+iN4gTv43hEh0MKJBSFBWNaX+tdThkTBskgAKTodNpZNo7Y
hZT/MiexFGYGC+4vBt99ZXJhIlVAmyG/XzpaNBW8QR9KYnEwNipMFzzrhXEo/nGj
0liCepKNA+/+gpfCOzXxwjuspOAvHnMlsl+AstCPFpgzFTpFe0DHCUuYJLrkwx2d
kyoe2/S286KJ2wXUCMIInN5oHkyzQZ+4pgvccEZzvOrZzanYkBYdZzSA9/xDjSRI
79TlRPsTrHUugz8GzmemRaFrQKTSP7JN9CHcwarr8eH47RvYSmMFNEYJftPJlFzY
xJftXh2BhLmd1+Yn0bNxMcnDk7tgYhW2zelfO7QzQpx21SxupRIR2wsCJvIJPQ44
Y0iO7dcZ1wz04vVY78IyR6JVnry4i7x1GnbCv4njp/TAFYhFOd8SY6DiE+mtUTDp
v2zT9shT2thirggDHxuqFJu/fjvj2mYdSqcq49cJJTXYgiT0tHx0HAG/7vkoXSpn
otBsQmaHHksDHuwldQED25d1d6pkdU70u6CiJy3D2O/534kijcnLI7BMQgGd2ALc
PTR6wlk1EoDag6+PZaVQGP32hurpnIKS4/S1Wusk5rOneb9syqI3jvMOpDKIw5mh
MT3LcwabAhacKZnPyeSXmIWf4c1teKs9X8R+CkH6N8+rmXMpfaQXEAl3ZZ1j4Swt
DWW+b6szMuRdBT1AyV1kzS63GQuYKAML+cukXV4Zoyosm/IdAz/aYxjN0236vyWw
6PZ1iZzLlvr2XNK/aVwuIYs1CjNhxyE9ha3j7PbgqWePXzmwQRv5lRJXCh++gtMb
a0r8eOKaw+DKO81VEDT1uKgmAhDA/tivJBmB5NC9QacN96uwCqT5tl/e02VPgtOd
iK2rAaFL3muvVOXym5qPvwrCh+6/bZpRgQqtQ5VcbWGlWn8DhLDVop8l4mSYmTW4
ETEpwWGBehUoQ5BZ16h+noGw6r2RgjXf1Yu9zqatCwkQ+p2Dm5WlMPCToMZC2r9V
H6Rg1mLHgpHb9YppkDosWgBr4yEru4Qm2I3A9TGtC3nfjoanSkewWy4/RZJLXhvq
xKUy8OlNoG/x7FRZFeT1OzYs+AFHnTMapaEfNz4Vd+xUhzSmEJxIRhkIgJ6IggcI
ntVu4fConVV2rcvan3YpwDAIM5o4ziIR0liBqnIDaNRz3FED7ooLpx026f1bNSC2
8lf0Sx7n7a39AYavzzBRkDgvohg9vhwGI1irIQFJe9m3GHbeqJpPEabMH5duAUqO
DG3NqFURm8KWEfJz0RbBJuLX0YPd/XL6QPoZGB7vHtV1gEOjQLxnuIpruBXu9SCt
HP3wCS8R5i5UaBT9zMh44FbdZd7hoMVoSFGC8Fcp0jWCE5KdNLs5DblBh2JO7FrT
Wpcve+XL6QRM2zKq+rPTe9jsK8nsWW/rKKO5vxuS9G5jpMlrVW/1yXYA4/zIt1cZ
bB+aWOLguxiRN8myPBzvhWlnapdGFp25gVro86nigBwdtqsM9j23zCT9jblw5gyM
7YKW5OKgB0eL9g6uPzbEt1y03pL1ouI/IfPS2Eh9lhvO3ZPJC+d0d7qDtXizwqJf
QegB8K8qQcqYId6TFPTt5Q5XdyuQUJwm6TLoIS7dr0qfisq86k/PEhJNKRJgOqk+
Ln5amQlSPCldlTInOby3VuarXGQrwamX2IFZMiq2upjiO50e+u+NwFa102WFfy0m
yEesy0Jv76/c02hwydpeC9aj0Y1JxINH6C6ZbD7VRU8SGL3jdalgcchbiC5Pbu0Z
qJMO9HkxVE9RYMA92wthrKRpUV2uTZOeYwqbsW/Lgx3UdFJxamICdlrrmxY6ewKy
rT4K5OP7sOo2GrRSlpcalqFYQxB8y1q9uW6WszfEpSmM6LxgzXBVCG3Mwx6GCRRt
mW0kflqzcvecXwujxJab+g419R3Ib5zcs2vwElfHO9BiCibQ0F6l88OBYfdHUdrj
ZXb5yZEsylNbou6c86fa8oE563siXtHOEu0+qHlTSUPgoYfsfwPq80Vab81he75g
Dst8NoQMWquzVOPN5PdBct/H3VUELtCkMPuM8wXjayh88gwbujfaqPso7FSkjLXx
WZGpPVZZgRow8S1VJMqbPh/lTH/Z+u9TyHGxOaArcAZ8fkWOfSldBkaID6RyNs9d
6Y6XRrtBrvh8pCTzqkiO5sqvDTenC38KIeLSuEZPG/kABI/1wHejyevar5b2uFP2
hxGjB3FDJZRjjf6G5Z6SdpK6wZa2J3LCBse7UdP+82LbNGkSdivoUmHZ4WovgcUw
/9IFfLPFB0JTlMWhMHSfugOBj6okpuI/gVukWQ/RWw+TGRNhk+GTDrZNfUxQOjKi
9T4wGkf5kgfTv4PdCxrdN9DAgCtdpPviJHeYUp4Z4tKozAVicnTJXOCh+Jj5fPO4
LVW9oB4kt2H1gx1q5dWZtAjXlHQfCfxY0Y8B79q7bM0zhf/cCpmGpKNuiXtA4nwM
zreHfnY/bNPy3c86ejaYRJNOi9Ts3+D2q7pQhxwa+wok4lA5BZgqricR1n2RHfc5
3w99mlmTwQ5SoL17c/jX4TCIOqhngSh0DvuMaMe0BvNkm4yF9dOt01nykBZKynsW
D/WPR9v94NKxbeKS/ZYGHYGsvbiR19dm+gPzr2bQduVqC02htt0a+ohygCIKjO4d
3HIMgHFyT1lNftnXU9ciQEO9mnmzIK1axQ5y4WQjYYMa7wYfIXedrcZT3jJXcxXB
SvnCChldbdB1kAnKLXll68DDTovetVKNTIHmCZjMAeAnJDeA0H0X+xGO+9HiPyLe
A3/7X2kuZYfx/8CeJhBinn678ELCyuZK/ONYjeZZvnkL5w4XlbG3wNdYwaC/++lu
Bkv1pOagaHoKP6dxuP6MdakVwDK0WZkn1HuTB8kn3Rt63tBzzDYp0S3W6MXHMGMH
UVgpkdXvzVD3BSAWi2j8282ZNBClFY4wTu8bEYRwuiKRSiXntDGa52H4t76CqEJx
m1KYx/MFtn895JboPT0xYfZ+xJ91MrOYS5zktGbhWuXJZBOc8kJaiZMLbRE5AZqU
K66TSdCEwOoA0iCjskuoHASx6c0Q8MHs/5cKmmIxSR/8Y+SlG1DkWx0qPgoKE+DN
Z+t6xMDdhj3c0LzHAg/BJ3aKoNSf+taWcjrolv2iVjg4+rhbgaU4mnaUi21fPJHK
Aykq7QG05MuUjPQPuel8C+sS+n7eL/afHGvIkzi/6Z5wuAGhi1HkhgpJXDDLOQCy
gGUGZHMJfPWYqnXujvsFgu0ATelPyq1NM31EKM84jMONBtRjzh0Kphr+HAg6hM8G
MRuQ+Z8WBt12yevRZq3YbgHnPASXgFyJpDRcnoAMtLdXDctwUCXWNEz6ks0/pTqg
MRJ/ForpR/n3CVU1fqUwqpSGYXIKUcu25qomsC45LpnBJxPBLosa5Rd1lcBMad0O
MdQoB5K0/EXYtaxcHjXoNcM5817Z+H26HmViRouU+ZqOc6A7I7Z3hELrN4Kwewq9
7HyWUEm6eTPLACRKWDeGh4YJmreMl9tUaaCDWAnShUM2bjb8w/YPX0t10+s3N/a+
4EwYae0ZB6yVrKlgiyGAmYULNPBhIHQe/mM1NY19fXvYoto0TeyopdfUnzcN/wha
TItuVkXwEr+LkhAGl5nGWzZf9h2qKkVMPLfjwWvE3zBSxp9WVDzY+BtSAlpdHVpn
9OAHqlYj01uwbPciejp3sbtNPxYrlqeBuqhjiv+4aNQ9Y2pUu+9o+C1OJhFBqP+c
jd13qhUsZi00g+Vweq1T3iW/OetDxEZxMnm5wAXzf26bHfz/ON8oXD8c1cfsatNJ
fdzafaGJYZOaoFVS9OuNGVtS9ALDjWcSwvMHJZ5r2SVfdeh0hgDyxe5JGV92Ylym
dd0nD+c6xibXfR/Es1PqkTMwr7/qs/SzI+trTW47xIey9TPWVt5rwANYzkUq5EQY
bVOnrRPcfq41RySECixWVK4LZaZfxC25z+Pqg2tq7eyeHobTI/32lfhoX0OW6vLi
wZkhzI1SYeF7RoMlhKuWfYMbkvFP7xioZovPnkWPYtEUEEmp8MMb1wjdqERrzO27
B6ZCIv/k+c4omzeerZ42GrkOvS3bbtadt9IRLcMGQDK3cwnskF9BaDnWGPQwnE8x
VXhbNC0ez4QrDOs/K797VjxGAMkKEDUwR0rBjMRn7JCl20SjirtPX9wnR+6FEgUl
yg9r5AzJiRjBjfWLRgY7qU6DpbXRY7G0N1A3Ob5nCY6SUvAeOUUDhj1Oq+86dNCw
H1ZfiAu+1zhQPQioOg/MmF3XPO5ldpsd+FWhC+G6s2gSuU0dm0IgbrqMUkG3la0P
QZppWM9PmQz3/dl/n0kZ4u4A+3N4s401jqsLlKab8chH4Gw+nzC9g4rWrEuY882G
MRKwr422uzK6eU4JRAZ2Z0ZL2NJ6o5zILPSgPVmDy78b/AIKs0fGZQmTPDz5xKjf
9iRc4Rvf2jNO/W3auonMouy56PrLWcUx3OheazVrRNOIXIOJXBtBH5h8jG1jqy2S
lIGZtVha8KeBg0lLrddA3ZfVwLRkLSYxJwg8v+UKLH4gRRsoMLwztCnw614swvTh
p7llxJnj//BAEdtGmI1ZnIqUjlH5+EH8G9x3brYlOif4eeirQIlVigWca4MJkH4w
BOxzyyxkwHlNEinWv5ZvrCubsbSBjnoHBVZmaxLvL7i2VLjZPnCJT9Jzx+1MX+oY
VAQ21CqPiyXAxA+TmDJ6ZMovrzoDyCAFCzZoKQdJwvHJI4uYZI3nkMTtddWGBT30
ktFwxrf/1P6/ntuWYVAZIh/r+VtveqmnjRO0ruv7jm92mN7YMVvvwEnu1J0SnDDs
duvmA847giKpeN+TIAHLVCG/w/JM90JcS7zQPJdaZLXSZvsLFwwVyKMZysUNZOq5
PpEmPcv3gjynz1JN4RywX9Q5Or4GtHZRYamICOIYc3MblsidwLZ+Y280HloZZUcP
yHtmmIij7cUj+tIoemNRfx6VXpGsG4BPdQhX8YSpOLLF47ZqNotVyKoJKk/maEUG
MAEewXWuVImqE9FtZeD4e6Hq6AzeXQYSSStLkButMiIeLqyt7V6xM8vDcEdYKatU
aC5XBmtyYJfaRWZYZgLi51M/ByxpU2w7bmXZV1Z3CxQqqDPubiBSIXuUp0Fq2QKO
KId59wGhwz06z3oMiAOmKks2WlwjAdvjdqHHtseukclPu1uBR11fYlzTBDDoHmTg
Y0dy1fc+6rPwb6C8E3xaThty074iLGApV0rZ31hL6MIsBQ6+jNpYex/g2O9VwoiV
jn6DaIjw7T6h/1kLqQvEhCo1QQMPrFfT+z8XcM0BTTIp0hcjoiXx+a0D6EGrFGKX
7BxOqoAtV5u7AItnxPrYkc10etD/T+j4+HDOCLUo1KZY2pDjTpGm0VHn4WW6GUDI
HLZTRAXXLJGrCYPntbwWDSHfKstPhVTPwUREnEHnQFvKbgrEcP00BcXLE2wZlFiN
Te1YaO9EgKL4EW7/3avo0E17hsp3gfniXikEOuCUwAhIl5uzDB5e9SLGAp4RuStL
JdAw2l9xXBS/8MfWzkHHUNihVPJPDDTcFh/EJxlo9hVBpVZ4eWZIdNMw2nuijB7g
0C82OmtPIaNuw9gN5+JOXw2COFw4+or/KSMHsekIle23NoXwQxyLuCR/ljEr9Zcx
8tLRLaNfRMviLDP8jOF5RubEIbNCI+IN+PWJalFNy+EBVWa/LxACjqRM4EGaV52i
8CWW79xr7h8dlhBp08F1Ni/kt+Y3sY1avO5MXTCuAZT2kqy+L3EOfOn/I8Sy1bM8
Z0y6yR6j6PgmycaJxq7w9w==
`protect END_PROTECTED
