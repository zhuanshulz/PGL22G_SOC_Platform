`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7NU3QynNKzXKXDEsA5lMvhpHBa/LZVbPA62yyxYPgwZE5bzBe63eQAIX1TSOnvD0
iwaMzGVr3QojcXR5SuM2bVXc72grai6lgbgvX7g7dGBaH1oW5mjhtlZAJ2fvd3HJ
QsqiWGiXX4erqgNKfm+XT7oUzCfyiVzKVLvB4p1+DDYdLzQwbcPbcSy4TjMjmaFW
cXi6L3wJsctesQzmwdLzRKzlutUSDFui/YvtJUvFhOioCFk++v1yKEXpvvD4bguW
X25r8bR/OQ99eODK4cYMnwLZwdKlxmWIXbIL6PVhhBp6m0VF+gYm8l2fZ6/70q9S
WRUkkmiAwMtc6+pNnr6lHi8foU5ikW+sa2qMs/01T65zQToj3+LKbqrsu+EopT2X
UGDtMHIE/DPwZnPSfWvSOgdSdEeBKWPCemhYaQrR222Gjk8n41MwkGdT/CakETLW
ZmK4uew8wV9w4LTXMzK/7WNqEHVCmg83n0vwUc56bxi6ncxw3fD95R8/91Mu5sKH
fe7ozBiC0VpaooryTohcRVv2q8mvj5FKlHZOcqh/UsWnF4IhxcLXSw0kfTqXfTv8
TW7IDUhGPmbez1VK9vjx5xp2g/3zm3491/4DxV0PAUHfuMtiBiQtDNCae2Dl7Tg0
n+SJaaVbvWYWraWqve66IqK4Lrum6tPLqJ0lILE6BN1QR184+m58KJoH8gjG3tms
vjLKyl0WI3/Pq+Rru786Z4EboNg9/cFWwCqIW8Y9kUjMBma+att/t2C42MWglR16
5uAzx98za6UgmvU//6hPplWDP+xQODbsvXZJqVNK0gXboT8FwgF1bnEf2jGBXpl5
EyAWC40mU1S7WfqdxyVdSIQjYRcXwW0NSDuqbT03m7i+nGvfb6E9EWHABnkK+M1z
+YCBInfqzPh7aPdsoN/h4aBA5IumcCb8ZonIky88PkuKeJc6xjSLKgpuIyjkzg5t
8TvSie2dnjLjRK4yTQD738bVBRj5FkZ1Wi/LA8Nf5nRNK3RTju/kpLKLu+NMwYk6
HG+hY8Sw8I5kWl6AYdSf0eUETr3KPTS7XGbpC+UBNlL6MUrFa3r73RWrHiHjVxkN
FYDlNWUqjKavTpys97gA+44QjJSrDYaUrRGS4CWRFMA87tivgMe6bm89pDYjr3Fe
7puxSVhdHaI39aGLghPYfSHYHCwrkf4U9XJlh0yJna+JBel07U7UowtYat+5km/F
2p1RDybAvkfc4/vWmD7NXuf4VwBRCa6Y0n52V8oEuS5ldfPwDeQr8jPwWuSM2xwM
2jwdc0X61sswWBjs/hiE1j7528p457bvDZNnK97dqrNeQ74cSQNmNz8CfLriDrll
caC/c2A2tBCF5bykQoemCEa7DmxN4r57MlWbrer6PTQpLhvZOBZus8d+BDFeiiw/
15CkS8njsgdEc7EyKY8MePh9Jzp7gZYhCdUMVyS9KaDGwuG/7N7gYtBQPSz0sOyW
1C7l0O3hxxXZpuroK4R+TR5m2C/jC42O1CZVcZoqgl7azFSQNlspljgSIA4X0e7W
qtUab6gTJYp+F7v3uPYP4wH2g9BpC2Iy258B6WYpUM65+zeT5ZT0cgHUiAGBZCN6
Wd9V4J+UMCu6kYWMMAI65y8+Qlyosu5Zti/1LVIKH85sSpiM0il82KGE6jLE4O8G
PQ4SAHY3v724zstqZ6z7FGiabOAynW/wvAX5B2bHZBRnGbds9/t5AvYtmAZjrUpY
s4ItPXe4tYDYlbHclVds5DgFvLS81/BJWy+WN04IUGUDL1Bl1L3cNZxOejXvOuB/
TlNeM5Engnt2DEz4FsVExCsYqw0pyetuSMtxkM7y8VYuepJe7AzZT60eL1AAH6H6
sagaEqlgpEVTgiZLNj1PGI3WPYvKmP1FBQv/LBJuNE5MQtP+mrEGe4jqpB0Xv4zK
3Jn1p9iBBlTeB/FzqJfOcNr0Co/JLXIcZGRmrDfpd1Lwo4Ffy31SLGMOz8CeBDif
3aG+iHgDC0SlcVtKamU3VYUTaChy4wqpI523CxqB3U8/38WR+oBM8Fhl3PG1tPkX
b1AaFlW9Dc1vRmQRXGXNyohHfMvowjsOE/zELKDHzGJ/zLhJ/A27AAN+Dkz1AQVa
ZXu/eORUhKbrbLQUEchop7cBx8rLXLnfwCMFGTZYEONY0ED2bCFjFFiPUzOzCMTV
kHQ6+oagrjTt8eaeI7PqvUXh1+ZFsLMAP/DfvN+Ei3lCyaiDSVXAPgFWqxT0tTW9
QVVox6gOIVAfbQ4hPZcKqyPUyuz5H3UUUweCFEnRhAz16FXMMQ6c13WS5LAdfBWm
e0z8qgPvDRn+3TKHaizEMe/XHAQkjxgmjSx8RpHXDW9iLmXQpU9d6Q9JdOWoNUxU
VEIrppxm78TIAeFBKQ6B32pEBfb+mCEa+YKsi/qvhPpS8pS2qVkish5ArtbwCj02
i1dvdzkyziUV8Hm4IloZ2Z+w4L1GTrcCFBMYXbbG4HZZpr8CWNTFpx6EfoNmBvcX
U3G+alvttrk9LQ8fYhqQv1PEN9nccVVYj9NmchZmrbg3RKwNTtyaKO35SYZhUmBI
J78An1ra9YHj8vbXBpB4IhhO1m1elNFqTWKuc8noPQGGrxWc61E0Xj7cKWTJMJDu
B2HOXWLLk+l56sw1TrmAS4rKsX8rSjPToVY/n7vMai1VQDmxrbRK4Q/WrILzEqr6
a/Yp+KdgNJ+aGTUrmWOjld6Oqdt0m+pouhR5J+nESgvBUaxEk9Rg9FjpnAorhNB5
u3fjcKWDZFqbw7h76X9Wq5NIsA2O3aaq7is81nN4otcXVvkebJiZg+YhLE0r64N1
u9r0aHPi/WgCeMpfmn3e9TGAWk/6yG5u7+ATLEX/Vyzz+FnfyWdwacBehZuBDS9M
lUkxHAcKoY0vBThpZTRgxjWJzkzSFA6tB+SVh0cXy4Dh1ham6JNis6DsEAcbMkeV
ppqnVvBPZvyBiJM76AgePtJWdY8Fk883SZU/gidxOO6h0siRdEkIzUzSAkhbbOvV
egRF3xr5PwLOR9f1fTGS5aaMKrwRsGREAPkEKDevBb2c6sXXxbnQb6461R+3Df0p
46mDxBNSiRkWAPa6RerxEgmMEi2x+1oRNNyOP+zf3PvtOopLcuKFYRhiKcyZ+++S
MU3/wguxIBaUagA9FJBWgnca332Uj9kMFWbTXIdO1jjeJ5PUkgLsrlGX+1akr2xl
7gENxgOUaHPK9ViTdiFgSZq6XcDu1XrH3263IBe12ZMczWaMRpK35DHHBoNf4Kkk
YrBZlCEOLnXa/C1i/ol/paErYehciG4kQXWZ/8MaW2DPCByc4WG9giA59oZ6ft0B
6KhsHN+unxZ9uW+hED2zSI4kweNs0YVTHkQGtmIKgjn7uktnA4GMLMOWxV7uE5wD
3+UHjwpcVrDwG/C+gkv6rLXUiBTX4TWrhBdF01ht5MMpqf2oylboPQdHZL2nsB0U
Zu6pj6zS0vYyUc2LDJbt4KbPJEPY/CfyZNI043tAvdV/ev752FolAajmRtDujiUo
1BBw4qbBbKwfvFfd0UcBlro48lhnkpTAoCx0ZrDL/INldt2MW2pBjd4+vAalM+us
6pBQnpZ06NX3ceEO/xpREHjyUBXaKqHlJQgo7/69JI7scjSx1vYWx4Y0M/PzUw3E
9vm22xNN5KXMRW4y1jj+GZR3eaPICRNTOiFM3YaYLKHZ49NY4J3PVA7wWExIH60T
5Qu2VfLpWARJC8aNjDyEeNJ525isGcxnK1L5d3YmW9k5/CB1voseEPqgLUhEb532
0VztlV7nKHWxcjnpugKLFNo0n9Z5KdJkmWafoHuHPtAbwLWkREYLnXSA2jbXMIe7
1UUEmjRhWi+WLrz50U1WN2KdR02d2yi1hAIENpsvyeBNmc4BEU221w7M5e6vcBJi
iMHwpWrhBZkRJ6W+fJtL4nQL0rr0CixDd7u1Q18GauKvBDLc7jFX9qHNz3egkGdP
EJi9zKmIioUw9nSYruFH+hOTpEbMzu+mx1uemyiNauDj2/bykIvCHuAtnNYi2iH8
PeVDCIeEHg3DAYfKEMZF6DaoIZ1rEbw3cUtWPxUlX5ydX2p2E/qcZSgHC2Q3jCRB
kfeVHCJ794BKIV2RbYTkejLhxWiR8FQ5J5+WMdBt1M44x0TKNXgdCYWFjR3Jscth
UQBNDTdgc1ebrFvG385QCC8RyBgG6aGW6ChB7oq03w72qtxFqlailxaVPfJ1uE/1
CwTEv2dnA5wTa7FvsIvCB6mh5LC4hneTPcKsd3g5xbwaUWjw0NSBsBZeMEJvfapZ
3siayy9AG0XHEC7dYYXWyTZPRt7Ar55hYNtnRclk7MIgJZk4p/cpnj1RqRk96LJu
qWDDHOBid1ceZ0uV5dNdHtSVLSo+rFAAhgrqFPUlh2jhgrUjSJ4A3G7LK2UvRKSu
iiFDa7qVtBQjK+dzNg9McX9nWi/8tMa7bsnSkWlr2LeyCWZ8jRtd37Ek2g/M8jIp
sJYbyedbKrVmIJiNb3kug+xxNpozjk4mSd0FyMNa7LuiTXq8kBWu6Fs8gQXmJQ67
T5U/YwDy8d7m30ipzV+i8qsvp5dzmTYx24s7CKoNPWmQbwQYlyj3fPRgvResZ8HL
OuM3pqk+jydqpUKRO6IM7Ly60GTgfkB9jrEB8D6x/RSItlHlkDeGsrSrC4EDvhTu
8KZgHzGhnZe5c0kputmtUZqYexxIVktHH8QLiV/p9tSG3bGwGwSPsXqsjSAhyRwN
+ki5yS/1rPtcbcQCcGJa08oEYyIm94K45teoMPFwWokcQJrhoq4qs2VogrvLN3Jy
DI2RjXZ6yCBrkOSDre4f6sE096BTuMeLN6v72VbtpEASbRxlZmmLWZWZqxS9ulr8
MGmeDdiu3vszsTGzZVA/QvVGvJ/0zLSyr1K+yaIjfRXUjZmKjxhr+dPll5B31QdE
ei6o35/Wj5I+RjcF9MgGr4nf5gFC4KucmqAtU5uvs1LuOrIujQEH7ny5DT9pl5p1
7wvtDtMmy60ZCWM4a+aCpKhaVDjGmmE8Viv0p39WrYTF2IlhqtA+0pAi/CnanJ/c
W04NvFGnY1N5zH/FvvnyDA+4/um+ueT27HQ0vXC0r1ZHfyl819uAkNlWMnYZlPqA
1znrGEeSYOBoX/Xa8lOxVnrutzI20YINQpCEacpKix9hH/U67/0MSsZUBia3T7fM
kUkNHxY3ydeWi8MDd7wW9btUFouCpqWWb3/GXsxJAQtRPY6bkClu7L3TVyPaqMy5
Il/Sd/CLdS1ccNS9QsSQsa96wD2fI76wNzP6OHZiYIKxlcxrodWI5h61wrNrThBM
n/Kew2O6suqXxlmAJ7dn16GTyR5H5LcD6ashKIU0hwvRZuJAFnXS2I7kS38is+oV
yU2Ef3Er7D+IOeB7ZsyCRH8LRYpPkoTPs9Fs4o0oUg981sWdLPYtaLguoZSwD+Xs
NB8rQE+qGjDfjXiMpcYMtn+BUByaU9xCqAEyB8PAiVqS7kXGQGFJk0VcRKH+tKXu
ItySAwkZuZb2RWjebX+9iCVhf7PZwNcqyCxsAVpfW3hQCQ9gOBhd6cv0iEtFlbCM
M9ne8STMHYw2gt9B5Gip2ioOJOrRaCP//NBw0Y2aiZ/Dgn688GiIfC2ZITlIdlxR
BIrLMB7oMH7vYb5xQmFbUaqIdC6sQq4FGjb1DCPQodHBY0doBqvh0v9DjasDj1/4
hFe7Swvcp5x2rUm9zrZvrHALDUAcSXEiERTBzI4ykoOR9k0I33/xj/n5o3CBKHkk
PBzObAvlsGKMd112lrMBjc2/t0YWEAA0wHKWz63d3EmU/4jhV8wm+RcvKu+wII6c
vzz2uDwLmnXcp3+5ERXEraIWUPWImACDOrF5p/B+UjDkj6bhSDqqnh9jjXkIa98e
3tChfcBtn8NgtUbZKR799Jefn29022YIwV5DPU2pxWhPqoW/cauI7jXNnIE2EQjS
4w0j47HO1tWBeuNSlTkG+umrS8510pJz4MTz0TdXdP1PaLqphCUlK+ZAxF4bwHvX
pT2+YpElxhH24ZPeqcpAiQD3bJ/SqgANqxMF9bXmk1vzpyAvmaBIPZ3VJh1RxgVp
M4n8Kv750Hk+g13FKG8Hx6Gx2tR/ksOcIC9u3C6GGJuhDuWIg2QdLQ80sH4UhMKk
jz75gO7ze3OV+7Kjg4gBh3TcwuA1l1NI3CxfFDZmsmTGJ+Op3Xd7aOGuR/QpA84F
ZRMexhU0OKiH6dHHtqgPOJQl92FQeTpI1n8gERFabQdJmVp5eVAHq/D1DLWQ0dsp
iW7zc8KIZ+W7ebiyJ0y70a7do8fk86M9zPC+q1zezWo2uns5fjW/WLld1wAEKeSq
ZdhVBvB/3H40PJ6IMGZhHRDBmIJtCUYRx0FY0ulQNe+JewVluoXmMyHMdrd8BN39
Kd7qTdiyCk3DTEuaoqzLx+ZBYsgZxjr6i/0ofjpSSObSqJNZ87bRFnXsFe1N8yX6
jAwf06g6x+0LxS17scINwz6tDpkF0DcTG4IVy8nkSFHluZoCxqXQhp6VPFaTuPOB
AUGBIUZtRfu8MPcQ75JyYOvisvXAzE08rW2AQEgFRC7EDJLx3wJLa4knN089TAFl
8+6hIRfHge3F8bw1Fpf6BqaMXL25dOxhePg6wDwn0go3dl/U3QHoWzYS83kG3W7o
uBFvgKlE8hjrj8BONAsBhqnMnvyiASmAvk2oefItAc7wc7xGtk2uPWKKpBWM41Kv
+6hEB4HdbUFSdpNNyq9lEdn/HOHY5+sIhGPfQ1MLdaXyGy6bOhZJjXJRtBj2W5MP
ubbbEc3iXd+heU1qcsNnirYrtgqoFe6gpBradtjK6NuASrqoSExpmqSsTwvv3brG
e+pNDJmcijh6xM/L8nTKfcNoaNaCj4T65wPOlimpTuZ6fkYA+jl8YzEs9KP+6Ptt
b1YXkWo11WjeLfbYH4iU5DyU4E58ERJqRKpwVYnhDS1VktDt+WuV9XgmJQGUDB5a
QfzkJSlXcmZuSzd4N/3yGXDribuSp0W5fy6i0TisfTVo5esdESmUt02x6RUbuIdV
slvvHAbUs3PmTrqvat+aeegoVWQgwUwbtuK2CSAhq2knVReIZgpPrWXxp/CXfuxB
qqVpKfGya7/OukQLuRcCK77wS8xOcvbXzJ31ZJb2dqo5WhajBlze7QvfFSpYxmka
gkRk9doqDTi1arOumgl64gFcvu56efPQjPLkjZ/KZRn7tzIWtpnlQ/r3aqOsR7h5
mNq/q3JpS/r8UjBWWVnzLpqFt8x7YpPhFMpHp09u6WfrjC7Sq2MrrFHIrNXI3hAH
OBfoc7Lc/DtVNYnx2KWntC2/esVw6EUe4nIZJUrC70SWYJMKV5mYbzLrNsOGgGyW
XRQQ4z4egqrUaGUgqbNUQCHJt7o/DYUvqRhpM595X4FNESdwDcKAt0K1T6vVlxFN
K4kmR00izmRsxR2IrFHhnz+efCvFumhGz++PR5KnZwEMXAxQ/GwkNPzc6MrWrGDg
5S38q0qlOOfG2Pi7Iid2NrxLlYL3N92UMy4WDJCCsKoZmMTLkcxuC1YYow/kFw6X
7mMx+/QE6cyW6sTvi/PmVa45z2w5bMHV8gbsqZsAMB/RgON8+mx0RVvtJtyBbTUD
b5Jkh/9/p6UPQJizqADruNm/uU/NLYp4LoNgK/pF9+qlCrU80/xV+9O6aFyujJF3
o0tnYACk1pSze/+FbOv48hIJiDM6Ddm0uQE9/5JsLF8zd69PllrCcY7zr3wdXwlD
ij1617jaMPhKa+y09qLPIGKHTSilDDprNC98HCfACj8jGoTrp38EwGWXFfZ8xque
+rExBLVW5+c2C3LKhxLUZV7rw6I5bcx6+5mtS6Y8MzvuZaXGL2ewsq4nJ1PiiMwv
t2VokJMCfiRi56LImjV4bj7d9sgJ6Q9C1K5pQqax7aWKRkvl8fwpucOnry5EefF6
sgS6aiDecA3JVwA0AmxCRDxNxBlyq9lDSZxRrINJ4j0hn4HtzSV7QMVgpDEggXUz
3P21LedJ7GA+4F7967QkoY9xPcFParD8fbEy54g1S1gVYDawe4h1IFdoEDldPLkc
50K1VRh0JX0zgHDyjVRb/0+VrEPs3LO5MLNBzbk3M/aU80i2FDfI+l2e14hlsVCi
K8kb3Y8e0MgrClcgAstk1HJCXNdeNQu9rjCs3XqHPYL87BrY+HpOWKlhKKUj/ulB
Ju5loFEFxV+zJ/ToC8b0hCdhneM9e5CqMnAArjLRnODHKy0M70kiUKKEcs56Qozp
fSGNkpFR0foOsawZ7fgNbr6RQBPfVoM7IGP3BpXF4/WFZLS4M/q4VcGQX1CHlaXP
wT6fy1F0curuUcLgURVuAkd9NEtXzlkIi4qm3FSZE8jDe7I0/hfflfI5ITVSJKrh
bgIhVs8W6ZMWoZ9amczi4DI1thX/Qb52/8QRJE2BipFmr1q35Ucx3/hUEQITTYl7
1MsWwLmHTM1eRATEOCUVCHEkMifY69BQPSZ0MW00zjkdQJZyTorV/4I57qrLPIIE
s6A6EeemZ54R/kTgaJwjoOQMW5OF++SlppAhvhP3HzjUlQ/f0JUEcSU1xYadPQi8
PJ+J9DZyEvvlLMXWlRVx5o0iJOs2ArWonAQCAQLUhWUR8NlR5uHFbM7dLGBxafxh
5wvnS8cZ6aAiX/zOrCdXHu4CXMHXGOZ1sIGg8U+Y2qTnZAzjzm497Q6/TskQk+OZ
vXPAdFOIHmDrSHSd6HoTCyl39k1AKFUg5JTKw97bR4yOwt6CTmV55uEyOFt4HFoi
KqnuvCvFJdPxN1oDvxVMxfd5LFXGIndkwiIlz0EtvfqskL7jEfSV8pkzadAlWwJm
XdAarrbZfQORxObznaa57sefJHr1b20iE+8s+BC9b1t2+9ZwigxO1ev9fz07Hwd1
8TUeILtC9txdl2hEPc76y6d27KiKHwysbKYUReCQOQ5Juo2uZXeSBzlFAr3sPKRr
Cmvfl6ulyVBIaSVgRTEGaqO9BMGs1i89077q3g11mUv3Z7rlFKJTETFllm8zJBil
V8G8ZE1FcvJumE3MPjfkfxM74bC38tMzCEUbB7sibmGDNql9TJrUMO3OR/JPHfb7
8hG8FcwYXPqXB95gty2j1A4rfzFvRTra7vWKynvO0t0BjgaTZ8U9Fkdl0WlrkH/j
75+6Je6F3H4eVT3fkS3xt3S2vXOur8Vf7tLW4K0d2YqE4jPgPQvSNVMCGFLSOXgG
MSAL9yzNxmauvtXwNvQwHcdTDFJNyTDeMtBHLTrFU+8mNXo/nBmfmX+/6PM7JNp0
UDnfUlFih6jPM6liBZVHHpjY6Nw5gsmAsA4mgGV4N5AsYtapzP7WkIXph7s3qS+h
NZWE5B3x1Lk7HmC9Ct5PNiN2oBhyxUz2pCRkzhPivtLgy7VGSICEwG4jNP0d084h
mYqUzEbiRVJsaxky45YuUQjUoHe/JVPhGtmgcae8I7k3x0LdRkGDuZll+UAvtz+9
FETSdxEuOzr+XoTIeLU9bNCe+NweB8EHz1riOMx31qdNkbDspvNMndyXhlhlQ7eL
NTDXstOWRC/PwnR8Arld8utqVkIEWnGWhA9Q4NWLJzcw8/jBp1hKvZwFs2ZIhNh7
AxDt5CrdadGtNCYzT2EFmjVIONOV6BDZILXloy4p/pEQCEXjbw2pk7GQAeEBImZv
P5H11IJDodUuEATkv2KX1bJL6B4OItyvAWZLl0sfouy2yYVJ66ovMV4jiyABTMUV
GXjZgalKQjvrrZ/oOSCYV/nSUumK0Y/muX1Xpajng4aRYSwuwmeqdfuugNcfXc70
bQ0T+59kDUK4YB+qqSUeHOVe6aHzni/B85X0IuItHeCFd2gYEXpTiSAP+0onytp8
Qjh3aZHqjMSUpVW85cFjSIuLbsaJKR6a5RUbi6R5N0EqBPa7HIyh373X8td1nHUg
xQvRfR0IH+JDs2Fk9g8l1XaBmag/AdUCmhSrn4lsvQnIh4WSWMk+FhyBhEIYNLg1
j+6rICxeoMDSBm3s3P8/MU+JwyW+JVxqKG+mKSGbvhHIccv/IkElgvY4gDVR9Ebr
ocoupTyXKqmFpMYhxs2RcmRQapvmZyi8zm33+BkFczAwZfxQ5Db1/OmjS6OTkeFl
GO8b+R0xpKb7T7Gws+q02oHlsBt4XXb/Lw1YTpnVPYrtvmJnT1a8KOaAxEtNeoUB
PdLz3CjV2iri1IINLxx78/Fmc22X6rx0YHEnrWK6yAFzOXejfmOM47FnuAouE0fU
3Yx9WCyZ7jA/jrww0YJwz90Zel4LhnvXpjOu9ZgdtJS1ckTCRvCwX5hWfvN0nE5Y
zYRZ/2T8A+N3YtgFU1KrkBOcRm4FCUJgSIFYIIFi4Z7US76b1oy7UFQ7aWcU5qvt
HjevZUiyMA7risp0XMih+dXZjx6zLsKaXwYb85f+u5bXMNL/fCLp42sKuGmrMAAU
P9Vqsq30I99p20uyPlHSNgFxzZ28ZOauNkUrvxXdUZWjp2FAelQ0B9MGyrvjEju1
o0T/EKv8snArWCD2qrT8WbYXuLz0+a4ztIS+sQ7Eoof0PGFGfZG6GrYbysO2L+1B
ACijkla0TPzKA4cHZXCzHoaxXm8qlxEROh3HZFEuM3NbdHAsMTCE52tuklfhqFZw
plpANXQD6Z29snApaJIsVlxUMV6wDqwpNpvgp6AQwbZiTK9C+b6QbBJeQPZBiTOy
7V1SIPixi3s2mcHIB0gp3Hv6QsZhqPeF5+1+yWW4d8/lcEk8LKAY2hCR/uuGhcbL
Twbr1tjlOfTt8XM/YxIPjHLbbYsf2cGiPJcZ+JEDYz9LCQBnqOWOoS6CBxK+lTIe
9k+nLT5Rc1VgO7JKscueYyBh/kit3QlMninsOBG3kCFHKuH6YJMwhemW8qX6aZUb
gAcPIK3tgB9elKHbeSFhb5EwnPsisOdlanfaeDKyfn9WBxCytXt020Rozb7HYiiU
hDcJvKyuIwLGhytr418uFpyEIfCWPjTJUyq5sBE4GpI5Glp1iHxus/qbl23RxQQz
Wz8f0bwyLHImRQUHzykJv+8SI3Hsi7BazWYHVnJc7v4KY4C8td6vVfp1ENH6wRAY
jDvKVkSUusKmi8jOOlA07nfflduRFLzNqKY3QYuaNA/wmF1WzjaQeVlkktv5G8yj
dfRTmn4P4cV1OEBNPPC3ThKGhOLQUE8DdpvH04g5JbWjlY7fVCTtK1VdEHvrz2CX
NiGKqoOjOQbqHv5erSjjhO218VfsYoKrAYMz8pPKaJIx2HqfAz6qCSAv3xQIsNZo
bDaSTxwckhQl6YbgpzeE8AtSonGyECt0MOq0THyOO5PI1bVC9urDbX15GlWKEqDo
ZVrfHrmSC+WR/NDmR1vPygh05h2Gfqv/MO7Ebk+MoUsNtkrej/Esr5xXBZO0+YjJ
/2aKje3ZYSulG/btNOnGNLcObEYnXzl47E2aNAmhA+9rAmJQ+hmlnzbi4eKICkBm
pN+KJ9+e/UPR8KRApFjBWUw1uGNN6di1Ia8g7AtOVanU27jZOADniYNN9X6ViKp0
m/CzSheKblyJXl2fLA7+yAzew0u/hlqK3g0bVwhd0OXAH2ipyxkopmQMDbvOIY5A
F/eIhIvywnrcbX2SgkvmsKQLV/wVtXKNtkjZEF+S2CGpO2RkJNpKL7H6k6eAH+hS
mkgPI3daHpVDnhUOiIGqt9EHwjkizgmCpIvmCJeHoe92z2zmVHjIRj8Kf1PNLHUH
k5Ot1x3gjv/jlqHGRi0y81EiAbPV3RoKV9PNYo0Hdk7if2NUVXduA9PI/md5KLas
HLRONbDp0HXCu9l7q9SXrZj+ZRBkg5tzQkyzin1pIK2SnsPyCFXzMA3bjNc+wBnO
iM2qS/+OmafVkaHOB/8pSWuHvd30v0BRu+vzSXX0en0cW2CqseifMMOXgpIG6Aky
f0J3m12Nfr73Gj7S23m+/B0LfTqFJzKO8gQaKO+A1XTuuyyTgcaYoNb1wmMAgk9V
wV3cyDUa5N/6CecLr/oQeMLKiNqA99yflHyW6yW3k7HpiKpvgKGczt7pEM4me1WJ
WzD1wXnx6hVNwCPPmAD/pUFHd3iBMWXkAfiJmn8PlsLQUnnn6JMtleNgOQ7xiS8p
g+hRY0JZieRsaYqPPWRTiE1fRGwbPCnjOSbeerosNRT4gc6CiR+mfF58bVVncJ8Y
X+Pj/gmKB9yorKeo5iVBYAvI/Ky1pTrXEOTNokNqGFpAbs+nCB1mpywB3RaWHrGY
kvMBPCC+YeVRr0OjU3UoHuxUOd5qnUfqmuSVXMMo5CFCmcZSUUa2/1cfUBEbssPm
saLpIQzAhRph4NT61chfZwYxXJzIOPl62JcZ6RH0t7PmzSiM0ybh1HRbWfuePQUN
IxnUln2T23grVI6/kp33w5zqhWQ8SgIWffELSvaXYlHrSbytXL3pfMykdtYMB3Nl
EuhB1Q1mh/wS3eC+iIx5BpC1YySBio54se3nogGtxK27VyWw5xPA1THG27YwJfBm
FKBJtZHIxnvB7cEduMAR2ebKhdndKSdhYRcA1wGTG76K6o55e8LRezReR+KJhZYh
Ur7YNr/6uagQYjDdYuCvpsh/t6BNeznnLDmNWJo2lkKQomCDa83m3CCZ8dLpdq4i
iMk72sEBTJTEsVQVds/SVMXgiUDr/V85dnUMtOrcxjsXI1subBByoYwybESUiy7D
PqbhkO7lPrB54hEcaUjd92+7WSE/uqdJmQCzu2YA6xRU3GLzZHwQnnB1p22XZqF1
kovAGuF1tkAWOELL8xS+qJGioGNnlCTwkd6BDcR/cFSbFUHVs92fcDmNT1QdPvFK
I29AtxX9P4QtzGU3vrePpOD047p1VZfOTAffzKSqHtK8l14+CztOybO6OFRmPSLx
JiUQKdkQH1PNXFtEgIJvv5h3HHybfLpDh42oHrDqpqxG38UaUPtrzMlf+r71/pta
tTAt9ZU9MQy4UxnDDNYDAup5C4Yl/SZ0WCH/DUQenPeg+LhyVQ+aeW/nKZKJH4c9
IJgzIsRhvAh8DxeHMwfKtshWdYRsoMDp/OBGem5Hl4+9bmuX34o+3AtC14wDv/tq
vcUoF5D3DjFIHXyyej4PuE/1VKYTX6wuFePdqqhNPEDxa36dx9pU2QLNa3aXi/aj
qJoCvAWe5pNHUVNk2e93rw/1u4Y8TPGnPoYvPeIPaBbm4XfWlCY6evsVUq/5L2gn
Aq7lHGPKM/TBTUUZH3/0SJRTlf/USt5jC6i4cnw9vJMDHQVUm8ZLhzPJeb0tzcqp
hsca1llbNVyPbAW3rW5YBm6RxkFvprYucX10MPxuEThTDBIIsWy0X493fHmTzQSv
N2svcfy4Jsbox4MoDiyyyf89cvP33fK66IKtPQVZ7yMzvpAkpplDzwnepFTkoAvs
PJRbRXPk2YkkV0UKJSKXwuxrHEz1I89mCXSyd3iBB4Vi9TLTVxn2JDj6d1d10EjW
EIryMu19yiOtDLku+O6DPbchkvnjpD9yTdGCX03YHyqxOpyLfvsjzDfpzESUcgYr
oBTTI2eP+tlSEgYZZijN22RF+3prxzBXeT2jztos2NxviV1wygvDOtc3u63C0HQK
vPv66q/+zIfvGLafRNgqXpkkqZ5+9VDL9mdqxWXEe31kjsSAu0eq3Rq9qLma4oIf
fOc8ETIdfamtGzcSv11Si9ZulHiTBmNwJjOOYce9/njObEcyH/FtchMHXsnQdh5J
oj3KAVeRQ0IJ5fEdGBO6MSeORggyLQSpOheu6NDIVvsEZ+z8Vi2tZ9Q0rQFaZoq1
ptjdcF4vhM7Rw3so7ehhXLFH8VIJSyPRdZoxFZqlVTfkPEn8plFY69UOLAkrjfZH
KfSSB6ASI7gPowNlon3DrJxSaBxv5QT0XyCIn0G2KPZR2oLHbK3+zIPXq+NviBtj
Ytuk+NosADItsR5MtG+wSSyen4ad7997Q3nbkSkJhXgsaWun81KGBOhzOQIMOZfs
JLGrOeBisbm4NEXwrk7t8vO9KNcOZCJRc6RT1vDUdwNlr/E3CfXtCcw6W3on0Nvk
DEeOO+OeaXeam1uem8gBGoiePBGWV4J8m9ttbpBMbfL2fLcPg7x8jhKOfASQWnX0
CFPBFCM5X1MzUIV+jmdbEQcvTUCYRGldqkfBCZev7hYxzMuWGWiS8wvQceUy26LG
sAla1CgZYhgmPEKYMhCjLfegkprG+co0+kMqs++2QJmpoVfNykazpGgwRj9catb5
P0v6xpjj8HXVC9PNl8I77zn1hwIjWd8qVkYj1U6itQmUoXzZp8WnWwUzd39/4mOp
v35KML+o8mWdtQrGRjnjaujjjRGkLnmX6DQfWZpIqgfBIcrMOR6IHhSNqDnJjqM5
OfsHrOx4fCJqz1k6SuWH+IveSANeUC2+DqLJH4YNaV2u0KlE49NH9Vopnp00APAX
Qk4cM0P26jOgbWvpA77QJBxCh04idMvNorVuCgKxYdNIHgemIn7bm7w/PVzLf3wb
AyZWnGyMi38mqdYQM4qXLSogj+QSLGttGz1Cy44JWW46drH0tQnBF5WChBo3aOoq
8h4qBB71qYAq+r3Ey8/TAkEX127ns+er9Mvtgrx6bfDNz7kd2h6/pex9d0GYTG7z
RXShY5x+lvR+anYuw1q8HYIKtIf+GtuG9QkzgEa7DDn67DsYFfO7l5mr5m70IVo/
n7i/QBA/PUVSFpq7y/WLwvX6/iBmHzrlZzXwR3zbLwKyu+liO0WSpuiX+9PL8+CH
G67gWV23ahfrnb0E2mIpimWyrAwYELJL1Z90kn5hiyTLoN/BnHID4WD+iKFAavcX
rKRVtCzFin5rISfiiuzA14lgrWEVVaM6uWj80kURlvgnGfTDcQvKC96lv1BZ8GK4
Lm5RPFwn1+G2v01+4u16wFh1dRABHV67uUjRc9AJVp/lURUNKDrGytBEr0xkZat0
s05eLgPgGt2rphqgKzgbAXRd+qRarfg4kY0kcT2r/fJjYuBnVO2HSCLmq9nbByc2
MaB9ec8M67PZ9RBmXoIidKAIN493hd//hMYH141JGmR4s6B7FAoLe/TaS1wPfo0z
9ZnWXTX/Y+5ZM5orjbC/atu8IxDEee95MZP3S+hjRBKWGHzhsVPfxjQ4aDH7NVpw
EZUoOvbWKdNivU1zwMZiO2dwEi5vTqS7bXl46Gnw3K6TpIa7fPM47egSnRiElA7+
m0skSM1KeZvgw0TqYJ1XSjEttPXHh8nEeVRg5oKBlpq3enOEkwYZcNH/iBg1FxSV
tk5tykNLGC+6Ss4nMvZ4TSxHeVDdUPP6Olu3Km7GBpiKuWC0glkWge2tKGP+9RaP
uqD8JFMvfWiHDqApk+AEU1AGLOhIWcScz6a/qO3myhbLqV4ddp0SbwAxSZ+OI79z
Ja+qEK5Vc23YuXhchqGAnmOlcz+5CkgRswKUz1qJ2dC71SPIIpbdF8BBk9fTI7qo
Lcge43bnENjSFR1U1QgGjS+PWjBLuNvKkLRF+mwzRRwud3qPELqGLJENRETHDJvC
MCk1xbIcj/Sve4eHcPhHhNuj5Z1Skn+Frtj/YHKZj59btdQ9RqhxdiYUKX8UWVKl
knZW5ux5TjoUUoWIS9UXjEpRVpVhSWiKtn9bVti8LPV+kj4fsj36ODnSHgawCVc3
pd80OBl9D+xAqcMf0gzq7BfaKuXoh79kmdss7ksVg89tWhjUUDNTL36vq5JbnwWY
W5oC1pvLu4FnRLxFGu+3eN+MEYGWyM3xAftpZL0VE3WDQZ8UoGUwehSFzWjMY5nO
aR+JWw2Fv/PMIhEAbVTREwD7p51G5HNMPydHiU4fqrqhffG/1idAebCMZbIRPUaO
Jj4wCQ7HeFykMi7276zDJ6KfMtnrJkHHB8nc4UmqmgoSMVttoTe+GwziLi8GkaRm
scQNLfGcjRnK8X5Bi4VppiZkvnGN1m0z9bRlQPqT0l3QCY9wCTbUhIRSt2a9IBRh
l73lfSUH0t9LfoeVEOjUYfVZDyYE23cPd1mvCkgrpC0zBhF+mqXiLNLoDwzSlq1U
q/syzjBUqPIZ39vRI9DA8JQ+KneEJqI+xP+ZpptFD6xa5HpmIo4f6vhhkCJZ+tPD
DqiFh+qzMQdEdsjts2StnUzvGnNQoTeE9Ol4oQmkqZCzV+mu6WOpHpMfLWyVoi2k
7ZOP+56Rf8R87BECv7rwmPikLwQnJSMojTBxhTWOAZYki51gRe64rMxRdH6pVR/I
80+b41788VS0mOSvDX3HdGit3I3XkmSh9s4ldsuP7rlLA4gTTWHshgfx7bD9vgdK
mu8xckTt8viXi7CdUlEwqbwRI3pp79/LIgvd7PRdiYcO+Hw+AjoWmlQjXv6TFCP8
6Z4K2hyCNC32ujAbVetoexV7CScCXlkXOLmBgk/eMQD7dn8056BP4Z1KKLAuYwtB
gBXbVm4IBNjss0L3ZoXfHybPCJh1s7ZPCEyzlCTR76SICBudkUEO9neu5xUZ+wCm
OSuAb0wQOA8EUPrJ6u3zCNfZnd1UgjSqgrs9V3xaR2h5gG78Iz+QalKOu9u2j4bv
rH2r9UYiAwSUxohOMeeYqo9Cl0ZTtqXimBMUGo4heaK7MewKDQnLy0wEUSTtL5KI
OBkT2+9aKnH/lSI056xmsrJpjlHbpDkLw54TqpHqua/bfnlGzKj2H9EsgYJnr/H8
FSfwGia1W6Jjize+oOqYBfh1TDuxJScwJzMDSJ964TIb7aEVF/7hyG07uAHlLCrp
j+z1YoOCJCgLFWngHdlY78eyo0n4ZlGCW4mixCHSf+cgWfsn/sLsGIIaMT5H8P6c
E2oXZZDT/fFObSwbDgx3MIle1DvU8tffinL0LRNKBt7o/0O4t33dJkwthRxZ7c88
xO+vbS97BBKBaG/ULAhZ43PpACnOFjehBQYHu5+8CvrkO410vinFzUxodyLF5Dph
IafB9eo7FIQqo59dOqnG+E4QAbdiXRTA86K8U8Z0Eu4CSubpd5uUNwx/eEnz6UyI
233H/3eCHN76JDCWC/EmWyu07iF4nck1cTjG+C5Qg5O0IaPOX8hnXBCwB7N1xAak
r1FAKf37xmWKtr5VzRg+O6UhmF6HQxEUFSNhb8O/Dt3DvkuT7+a83WlIQwafb30Z
Guv9hI54jUzWFfICsVK6cubbKYOQXgrxuw4u6fR1dfkrBa2T7nXV/NPNWoPVVLWf
qTr8JtVWlnb6DYU8GvgusC0KbVEy4U+Py1iy2EDxpwBXB1Mc/LrhRVLeDrrMOwGW
CDYOCR9giICiKXN3z+BYQbb+9GNULR6KcGoxqHO1tyXRFTp8Q6MYfGGtOglvKM3Y
znJ4ykqcw5vipEt5ozToRBgpap/NmA/kPkVF5AmyfQTYkK6G/ENru3ApbwILd/SH
uftTbu/GlQCDlfSWjT7Z/16JHnpkQOusvjPCFzNwoJESP3oeZF4skv1i2uY/QW+Y
w2CJRLISoYzKKd+TLu25m3YfNFjfsFBp+O8fL0b1ux/7JNQ4jpd5+Cds8T8oasvR
fWd8Bl1odIYl6byAQUKf1efsx4q/rwpw3eNdllYN1FeprDx4nLh0B3aIpgBukL7V
R3Z7AAn6ak29O4I21NHpBNcfu9DCv/beHuiTTwB5p92sgGWOlVKGwLV+GJs0GQH5
IirK+amDX4M0WOCT+ACXtCsXO1ovAfwdt7s25dxHee0t6Dr62ath2h3x+oyvdPND
3xHH1tuf6MLMCzWCZubh7APPBK5T3XTlpZrU/0mjVAwbRB+nXw2weNv2+FGApZEc
bhIxzj3UrBXf7ciF1SmZsHuhw49X1qSZ44icYmw4t2uQxkZUm3PbstE5F0YzfF0G
P9jbXFHPxb5NG2cs8KCioP9zz9JwAVZgbx5VW9aQX83JGU2olmdpmE0h71fLhVds
UlCIipeyPtUKiF2e/srPyazKXS5PdNLJa4uedWfpJMIpsZUgwXziSKEYvSyn5KGJ
m+zlfgyoUQVF/ZO661yk30hTi0cDAw1biBafB9OkoJJFL2qOTeH+j6isZsPvfx0X
iIz/jRAbn4w3UYjhhzAy4Jm6l4Zggckp+iwe56u6CfXlkB8svOaQkbr4BLIeZi/e
GxGy/NjzLSpHZNC56Azj2GHgHIi/YXqM6FkwUqurEy3pskRglR+/BhQUhop46rx1
lOrwtshMrFQhiAw02FIjKnKKXZy31UIeSGbGodUmip7DfSDfFQtAi9ceKlx9jyBF
EiH2IEXTBiM0KgrCJAL1vxUfW2VF8q3yumWx/Kv7IRd7XGpl5L4LqO6oSKnb68GY
PXn5BOczBzJeaaGDUo5eThaNw4nCdSOPaf2s72a3WZBImOUqBT8ZoPs3OqlymKTM
4jS52qoxo6yZ7ilqRDVunobGtZOv91PTu88zuhZdNKykNvyLJHHswEmcrRX4kuyU
Tn/V3oWrueQRraA6hOlfhtiqMctqFHllZF4XrXlCUt9HCI8mxYHEVQKIoyZd7w/3
sgBtFXfqbVfWvzizAtC+WuOrAs9RcB4hVkpHJyEQrJCv852uXZPZtZtv5E2MzSg/
6P2claiEnPMfsxNM2QQ3au3Ol3xKVlO4O05hx5xEhNIi8biz3sWF/Dhd9vmlt7ox
cs3Qu+VK0Vdl4mqNCapdOXRZwaqDW43/oQBX1OA0X9pWODKWIui8mSmKYmJcqfIy
O8r4EIUQiKzLLofj6DGMeCbfs3PwZKWRqwfj0vwKQsrxOFOLJVBZasmYF4DZyKMJ
S1P1cFBIHsYt9pLXIs1M6x2R/nyDRr7IuNIY3+gvUmE8Tyf7ncc1ZVr9JLQfjPOo
9Wto4fuSphCO+k7FyV/L7pXUYHFJ5Kgc2mvnldmpIcyTH2L406gfwPjoL84BgR82
BwYLvyjuG5eBVrW6q/a7LkjbA4N0raHTJ2FZQn0qxdTGVHyem6Jx4emYyVrFHUxQ
srUj1Xt83GXieliwGB5Z8HIpasP9CFo/mRZzorby76LPCwnXx5kU9KJ2a5z+6DqI
H1gn3G0xFQyTfvFZAIt298uK3UF/C9rSgfd7eE8XVaFMc9yNTd2iCLGKQ+BCWifD
7t6r3wH0AzES37jXSu+bgvfzwsUFKPdZ7iFw46iEN1bKJj1HrN7MNWHsHN4Bluc1
przpwyhiMUQw0VaYfebwdXo0fSezDS9MKLHYaPrXjbrL/kFp0yqDZopLIWGT+XYj
ccxJS+P8AzOVBAmeTfj1k7lPd9rlyjV67RrYg2wzCpjH7mcSE5MKBs/qgDOTnYCm
raaAnICwGkz1LqfFAzdT+0XQajJJhSLJDw8OG+fcfR/7stuzequt3zl0R5Mws/7Q
a/OHL9JfVRYcx9fne4wwBStxRN/xyHVbBz+k7cWluzDYlV2d828+XFJengR7nG0S
gSZcw11TuQDgnDsxQAN7Kn0sIwlt5mp3Kaxotd7wagu4P2L7dadkgzHGra4spg0k
vykhr7QDwcxgnlwYovcQMXIMAQ2/nDDOP9+F463thzqyonxnRvERDgkogZlEnwZl
q0kqDEJUjFe8IeKnrB5ENhozcRIiqWkKMg2V0LwKexqAqX/KdQslfdrVA5k6NAAb
NZQJf40ayL9LF3ouPI+wTTiA30vnE1SGXP0+Koj5+pKr1G+GDIdi+JsuIE5ouc9T
Gj4KlVHpxRrCblcA2Dq7rhJ32qkMeolV4jflumUE7m1YydWadyidQ1QblYgV9L8T
H35WYd3BwMWQi6mAQI92BDotQZDo5bC/Xn4PKJFygXrBHoWoDexweEo+6DNZhiac
bVpjN+4Xy0se7Yel6Osi6jYKo4TxCb7XB1myVfhOCN2MTvDxzOzmBl5lFWtHyH+B
Wuoy9U5Civ2RnDsQ8NY5qoqdvCL0DhyZ50LxHH6V+iQMl9MvdhLD7eIaQZI/ooeE
rH+eC+Uf953FSvqQmWpYr/LI+vNfLLxcLbvpsjNoIdzSO+uoAj1insmrss0/WBre
Jir7zP4VH5B1Sryo+ovxFoIpi3NU31YydOb0Zo0ylv6WGLZw1bqMTxPBfp4pB8DL
tHXZl7kx8UcYjOghL+wcG7YbqBZ/HLpkQGsfAANm4T+V6v4vQ4bhrNYGIchUU8+V
Dk9bC8CU4NW7sUU5LU4jPz/z9KZ4h2sEI9RxmjnoOJvYn8n8dxDbopuTO0tyCxNp
CanPYG7GIynSAmCLxhKIKC3Ml2xU4K8gcshMY+lGfSver9+P9Ui+9l1pRfeoJ4uU
YHTsACXPqAQvy/BEh369rXiGU+wchP7o160tmZTdj0yILxJ3Yj2iC/zN4NVt5wRe
o2NzvEtwI14wyfPQrTrn0L/ttYWdVhSqv41pgvhitXeARs1O4UmPoZ5l2LaVvN1Y
rCqdzqEKgBjo0YD5adcn/ExJDNm9fF01Y76Et0ueoHbR6gKx53gZCkDLR5FEfm8g
TVvwRDTyfk01P/PSdFs+r5cdRPniMDf40dpMmwMHAUUMwaN7Ck8Uz0NH+JO6SW9K
uLce5gxv1yjQFpxzuE/CpMzsN28cWRRMmp5BKxU8NVXuYZtWqci9zyjQ1PAwdtdx
kqUGQ/WrCV4EzpZ8aUtey7Wthl9n/boxoB+5MbDuF5P0c9QPoClhAoOLCYnJqsbo
Fjt6yUl82jeELhP/QqK3PvK7JHGHMeRpwZ0xzLKEkLZMaCKQJsClMFMcbUc3UYN5
572pJJJpNnVHey8QN9ENQ7Q4KFgQnLjBhvGT03aGr8aLmXFOXN+c+U9A2De6PsPa
6xjkRszdqBYGI0orZkeZOrKSfIy3fRTrArZCDCKsNpLetIGZpJSKTLl32CatyORb
sZL9S7J1gxcIJ9llf+EVMSd3Mb4P6I0tx+v4kU0KNHLQp7ppr8qmwhqcQg6sqP6Y
4GyCr/FNVizGzrF4i5rfeacm5tZbSi1A1a/1GBid/CyJUGQzf3OITJ7gAGDKHVGF
g1yGnkimAO0r0JI3ok4kLPUlNupiBjY4mOT1Rrc0cZtpwI0ddpRLQoBu6AXjGbTe
blNXFGuYkjVoSqSqjVhmG9ebZ5g3d6zVOZARfnPcRnjxvlVl3Ad/cKVkyRNw41Gz
6zyPSrMfjMrvhPlmfgemUjPgRejFNq8hddx5hJjIiCm7A+fesbybHrQ12QpM1c5P
3nG5E7RfrjgMIH4x4QJYoi4heZEPz6PJpX4P9KBTjIYL5LOVwLkJYVmozacZxzw0
W+8cYPge9PZuFuKilLpB20VMl9IUavooj4gHrFns4XuZ1Nhi7fAZil0miSURMXUQ
kPskmhSKzjFRDM7bor0cAOr5GkONQ76pAWPkkRo64J7qDH+Pah052Rwi4JeAbFY7
/7MXgnsgroUaE9S8tgknp/KDsYR3gQaV173ZBARMs82Ek8nHlzCinXhiM2dRuC3f
ZqmzZ30PSYW9LAqpbm+IScdHFHzr0SUPhJQF4HRQFLkF5olNSPXPHxbSby6I+6gy
ibJKO5Js7fWzHQ7WoBR4K0/bmWoQOXoxByd5bRqop1jQe0qWnUBzyyc2diQ44Vyn
DbFlmb24HXNhDWJyeJ0b70kv8SkKH3rRnCUzq7FA6BMsfp+K3D2kJXVVkzuyjZ3d
QWO/jh75CWHhObDzmZvU5j9ZnKdg4tDjh0f8NdLmtsMIIXVzIxmcZ7vN+MlNocyJ
oKj74npAodfdnyL1rgHfNlBm/MQUfVoz8Ht4vh6rZpYCfVcfCPsC5+Q7sKGTtreb
DQX12aUwkQjGCRqPx/o9foKR4YK+zhQYQW4Z/2/3li+PF1ldFBzMyRjJNnif3O5/
1siDi3axc2bjycY384SD4eVo3keuVeP7XyhBUq2VJfFz+B/UAruo1K1w1Jgw48aL
ngjRruZ4v9H5Atee4HC1UqyQqMJymwvWCHE6qXN2zz5OIEcZC5ETiL4htGZrKotw
qIOdx7lpkdiEqIiihE7aT0bwd5A7QIOpLSrfzvtkvo2+N7+dOLeAz/NA3Uqfxc9E
luSM357yzr24fPBslyUu4PvTh3p/ygRrTb8Y1vvyV6s0sFzZ/12TLQ0+oG+/qWLs
RpDF7hLoCE1aQnT5d4H8Cd92g2iYZVC3dyoKDZTo6+i+X7ehfLgB8frc+kJ05Ak/
dFpBNdXfrNelJ3goQLYOKxSiylaFNsz5xTszSoNIOKWaJ6ur+NHvM57vqDoWhk3J
/EmVme/9bvIHnupg6FCyb9dzRFH5zU+u9L9L7j96wJUhICvWlq3x2mEcNZgMcBlO
wdQsM9dPdVMBzDMyk6pghvdh1zY4mpFId0eTBHQUlqvSvTUof7il5FGTCZF9isSb
Z7sVFKt6LGdv/jhnBhrCNVX+6E6Q5ATaZ7PhP6BghNOatfCUb4L77xAPfewZ1r6a
WHHGTmzUZwwCi1wEX9PXVZI7DY/1qRPTteMfzcyctCbSynL/7JnAQR9oWsyL4+U5
B1o/f1lPNeAN/7516MfusiN/LCbi8KBj0i+rf2Imyx9AmNJZQioLMm7tjmMSuMWd
NVZ1hVKMt6pI8DQR9ATFWtCxoE7WDFIn2fPqxtbsaDPVgb8wFygvRxXhqwB63B4J
14wP/z+fSYFl1oqMVEDh/Dw8RHAsZ4wOm6FduNDmMNym4LMDtqF+BCcV2UhJrSrf
Top9NTl6CprnV+rpVSIm+4XbYBEjkb0N3fQZYwJKI9vAPS28siDdo+y9TZyP8Ic+
sFNtVcNFsalwRr9FnHlP2lFx22k8Ed/MSxQFP8icEdv8EXBSAUYFXB1455BcXjg4
jneMg1V2bDpJQtYytb2E9A5v2BradwYFEmaab8L6KVMK6DgghkicJL+bg2ETOfkN
ROmNOvtFCgeNud/6Nib0OGPcZfxRrycwCy92yJHizSSgt3AYFx8k5APdr+Y22RRk
c88yS9WnLruxoQKRmhWziP7ZmpkuvFMq4cmU21ehTVYOidfqMizFkun0oOnYOWF9
+kDJgilSmw4oS60UiYl+8hcbo3F1g5AI0Aaw+u9m16z6jLEPUkdKEuyjqeY5mOpg
UIxukFw27oKtOWA+0gk4V9Zp8pJ7qwpxkasQmmV1+uBcpo9d40JHgNXC+DhL9NlF
JC9g9N8MItGKbaKg599SV9F1g7ssB47U2BLsTzCKP0twmZvMT8m1f/ZAcJrWkcpD
Vb6vZNXg26OQoT+/3NkTKbOcRLVjzRbic5PhxQ+rDFeXdmcpfOy6mLmeG17NlvNd
S8yQvb1RpFpcKUq41zu367MyfXEyTD/sfPR8/DLcKC9CNYa47JddIOlvkus7Z3CD
4uQrQAmjAtfdyFbr7Nlcb/3r175AVpXO9q2nWgJb2McBQ1rqvFggRozzxBsMeMsp
UUdRye2LoKWGf2VRw3Zvjyxi5Tk+heZImGMGo/ZKBD+uk0D+HmKhZcRrqgiL5P55
LfGuGQmJlvdK9YgU46hQIZ1chi3KOZbpUqq5xlFloboX8FM7XyTsJRMdx0hk+3pD
4Sm12diTMp91krxRg45NYUf8rVJPMphNzVvW+YxUS1tylqKh0Yd1LoXL/bvS232G
2Dhu/RPpwt+h1Nwl5ulR+z2EcgkiA3PPU/xYNMc4NjkvPOROH43+8yMHwbsscn2G
9scAdvZs3rgAlHQYeiPn6cHm4caijbmBd3cJpO7/DC+ysoN6Jdj6NtZR0UKe0Hbu
+y2+5t8V0m5d0wvCbP4t5xNlSuNDl0qXFtka2+FLEtBy06yWTYjuMmFfwbFM4NGq
DrJpPL0C6pmlbHjizVdzVL3w8MDEYrMdfv873E0KVWRcczAeHuvyQp/39AL0RYtK
krI7AQkhSag4vIT9bof0pJoZ6qKq77erpjApKfch832rW9e4P3qlUUoDqdytcba+
Ko6EFIcRbgvBn7/Z/a891xHFnNC0m1nDvP/aToY0BU18pUQnjKeVL0lws4YOyxH5
Bi34mVNt6my1Y//009heof8cOsAX8eOZzT7V4SH6AB66OVlldChMRFvg6tnwPc1v
DehQi/Mg9H0xMSeBNCvsCVnhyAxaKQ5wuaxsKfdgjD0xY7+1QMHUT8ltIkkJ/79C
9XjQacHPsNQrENnR+wPz7ijD9K3o+dMmPKkNmN7hzhtGDEKEV28Qn3CkVt88Vb1R
iOYYaKISAolTAAHYR0iQ7hAhQz8yY36D3DBl7ukKqJ2nC5WUidItr5+m//jTrXdY
FlIh1ZYe3LzB2a7KhOk2Qrrer1/WmdzqVmcIcfraj6lB1XmkMyF2pxl7Xu1NmYo0
93ROR+75lb5PBd5If9UMjbKrvX3O0WqmvE/VIRuDiu8YHlDsavsBGjwOjq2r4LRg
hlSkRFwop85ehR468Fm3/+nNs750icBfaNeMvQwo31K8Jz9elSA6UFqHhIZPnJvG
bzJjDjRWcl46gdcn4egZwLNE2/NNLogYlkb5UTjuUrhHfSTkNnHkDYuFw5opKQlf
BY8/6Qmw54+AiwfBLL3ACP7G/VXnSexrjLx8k9LEgKHyrEdv2fu7yY0hb+EokqsG
SWbgfks3G92Iz9hbBl3lGAsfbubzDtAyNqKl1cVjZfdguXFACj+vAC69WYL1ssDz
cmR9AvlN44WuPE0QeZ4mBy64tOBjJCpw/Rr8bnUSkSPLfp7IXNPNhxKGIHIbhPua
tZQ5IqLzeRlF+k1IQ+iGLOlKuqBEUZFxQKGIDYqH747yeSytQQazGUcBuwd3ut5Q
cxKIbmZ6eIwN0uy2lpq+HqujW/2zjY0G7rjtNHxUwOsu6BS+ti+FDr+1wybaQta/
+33U9B7xh49coYjyIfqaJQV4PJW0cimNS3Fz5ruUQ8RFz6iB6cp91usv331gSgWy
jYYT3+ihRZxLJGS8jPtaD05IQGX7ElUuwO5PM5yWaH1i/2DdqfaA8oWvhZzHnYPL
HogcgOtuMIkX1ciFqbpcyyXCfPjGm+kKOi23w5x9EJN3HhYHTPRbnU9T+mwDoi/K
gJZ4KDSXzW7VO0G9j0gy+y1Q7Du4iUISS/uq9j3AU3ugaAvhh8ve17LfNZpHqWEJ
xBZ9GDPQwWKFmvdrXHF+f4sMr/93RvAWcO2rG+zwx/qmUJLyjIIUeXM5oT6jzVss
QHNDurivJk4sUtYJohJFi9YNTaM5PUEPuuCRe3r/PAySQAMdc181IqFkaDTEQlO6
W3RRUFMhj3g3b+REmEN7PLt9tYSzkLnlAbTFU5FAAEvIwqXMIlaM3q7SqYmPisQn
ewY1AVf+mklWxt2IS/wnY42aZkWzLoibezV5vaqIQxR78MBbH+WR9Kj2ubdzGQ/+
GX0XUeynsBh09VziH9SUDFkCtwq0+7IgXNUPkwxKru/N1MkGZeSPFbP0Z/JzbDkq
5ajXBP/T8WTVRy9oIUfToAgvhkNTh0Zfn6ba3Q0yJYWt+dJBAgYViboPKTr6U6+v
`protect END_PROTECTED
