`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nm1nzmQt//uEg5DkzqcflZQGS9tqJbSUeKbdKl4OADjjp7g+HvUthjbQ5V15MmX+
jUdrollCiN41BVYrcnmdr3g/jqqjw3T/3EMcYpE3pY2NYL0TstTZWTPGzUElOJO3
8sdXcnA/HMdwSWMPEEb4EiySQ8WZ4bkFvisawb7AFegHXx8Yg5fllS+sFOONw9sB
wZelg7DXpv6L3Hbq+dcMyUQKuUxCQt8XEFK/7lKvlBQ7j2rqY4xP2IrJug16VQ/5
SyAwPxKLrtuv2z1cVV95ouqwq/Bq/SyrJglueijmZBrQIZSVubBNHxYRveY4UdXd
eVriPGwyo+vEqjYRAKHj/8LZC13I3zOKe2/zycc0xd2Tt1V0W8wkchvtbgpoy2hn
2U8orBcpji5rY1VGsNTY/0iMGIdgxPlnjcPXHlNBsyLJT909wdiatZyiju6/lJIh
foJ7SsrM63B4lrQh8/oC72MWIqagrY969T+8X/kLhw4eZRDtO4uBnZV6oGjaJDIx
if4L3knbKejkpmrkX5gQZMDkP0+vYbxlBLjss+1rWOcfIPJ57DFBUKeWgZiroHa4
G6pS4G+uIZObF37eNEYaWG9ZBDipva1S5wnvRz1GaL1oYTlTkpgUrFonxvBaArw9
Dzl14ClnCExHNa7Ii5ADa6j6anQjRHNOrZroT+IWN7/XWk0+8oEBxP+V1duralKn
PJmHXs9oapfsQ9caPPK+p8XIFpAqsfZgbByvEaNoyrQeJJO+AYkhXlpp+WzARI2o
ES1rRAY8PHIPoYH1fh+EU6Niny8rzcslTme6It/NLhgTiNY5XG75hg+ugMkbYmUv
I3/019g2tfUd5Q+bHgnALFUoCbvP1pUo+V4HQ8YmeQdSoBXrYIzv/HW237iyUPtt
clhsvCxGH4Fo+jOPt4LX0v/uL0/+49QXqyLDf+VgtOO/P7C4iBznTSfI6vriekfq
lzWW6ED5tKvZ2u7D68SMzKGVmNS2nE9smsi8dfT9O55vwTykG1EELdAKCRqLHmoE
tSyqEhmxlP2IdCBbzELDb2F7Rn9DG2Ce/7yflPn282mvYvoKfNf6XxN0YAexV0L+
iLerPwx7r2vu2uJE9xOjZYTTGj6pZkSHLgaOni1UTGYWstSZwsNfnSD4eyMy6Jsk
C28Xo7FJ/vQ4mFvAZ0vAS3Eft1P4KrlxG0FfPklrrj4EtJ1u7eS8zJjfBsA4+Vux
19vAqgu3Fu5LWL0CDqVEWPn4wvCn49jUoDCVm3kabw3ENe7Sm02yv421T7JtQY5j
spf43QIHYBEBVgnJTohNxlCeUNWzy83WJffp1VQ3Yjg5ujesl/4IDbVbI+gOmrjK
8vI0k4kR/RakUIQOSrp/Ru4349YAVke6p+uz8QDMjHQzfvoqOBPi/dkFp7tZgJav
EafaCZlUq/PnWm2GU5wav4uw8rKTH9UJK+4jutMin6x5VopZ9sQP2UnewNQkMk+u
5JzzZBS5/iL/ui7jeBEDh+S0RyCDqBAjN9IfnvZftKTJNWLlvzfHM90vp62VOnpe
x2354ikS8sdtXPmTQzUKuxMON63WG3deN6h2v0ST3xtp5155JJE6bvsOdUwi3Mom
V6DFQwUlASmyVn7UdWNcFIeyjogeqv+BeBGgDoSbHgQwQlCWjK2TDlBp3665+r7U
9JGOjdBmd+uwkKClOdAih9JG8Aq90uVzWRYT1ZA+f9jugH1b3FCPuhroS5SqG8Gh
E68eAk7VFh3tyeI/mM1YjwDXPzb8/0y4aqsorQRB/SGG5T1HKav4oHIAOaJM3Ah+
mcc5lHGte+yDTXJwpo6K3o5FUxigZmX2vLcn4pEgQyqasIswMXvzOjdgcBlAe+Hm
RjVat1xSN3HFgR/5o7fBPlWzFBngYoysX6IOsiPIs6eqytX5aMd5xcW/lLXNu4xs
OaaomyTCcLdd/VOJIlFJru5pXb9omP7ijCSYHyFk5huSt44DGRJrlanDc9lzogTG
HshnSyjyBtwhX4+jYt8P4wd0fLyeiWVVPECBBT3tR/fsdcqeRqnxQHMtQRCUpYpK
wfnloMp+7p60ML3HW6pMp1+cJ3SBPW7k4b6AXwr3JZieQ7XQ/gdynrGWRy5VwDWw
`protect END_PROTECTED
