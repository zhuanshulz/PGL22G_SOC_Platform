`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t7kysVR9Om74dZW2Qtal7HoaAPfJ8wHV6BFYo0cNiUktxUvVFvdxqAWv2XJPXT/i
pMtolir1reRposPJiJvsmie4FlJV+nMvRIkJ8lWIrYP+okjk4jsSZH3HdRf95doT
bpZIcQx5SiMAYqHEhNPwkvhDzlvHQ/5dPrctVy6MYpe9PKC7Dg697W+NLWP+C8oj
TRs3iBaYZ7xvr9OZ9LCgOa6Xe176ykX0RVfKX6NWMl9Pkd6E6m6LGWfSgWk125Yi
p3JmTPt+TGHnmuS59cGZD5m96EqgGxV5SBDreMb4BXF0BEBiuXnhkdLP6wSnWFLZ
GgquIF4lagJYUq8sOXKaPJeedMvWWUiec6REvi6JgMkVoMg/WvCADLF6ehAUaSXC
pIu+5Fk6sJMi7SxPupJESZEl4W4jqNhovZ0g8ocPeY0IUUqE52u633ZOm8rgxeX7
/f3CBVKFAykLob7xWIZrCyPXqg+GEYdC8ZF7NLr2vik/7KaUYuiG4kxgBFD0coa3
gqMld5LlP6sgYuJkM6rkVwT67RJU5u4jeDgNVpMWuDi0H/z3g0TgT94hCG/KhT04
PCBihdw6VR0PGJTpsjTFSbZTFBzy1IhHZ9G4MhgqCBkGl4PghICEvFAPubfLV6RR
hEZdW464SE+rJCXAmAItOMXo4w+7Mcvc6tbGqMfAA0nhDf+K/s2VU6FAmgs9x9TM
vSW7SZauLfoQZFqosFfmR4vbLhU1ypjyIQatxO/4T+amaeU4Z1qEhdH9IpJSmIs8
ezfDffxnmS9FVWizDvTcUQK7WpUGG7KPbywQHHau6DF9zQCatll7DL8LDJoPd0R6
dpxdK5+nawpzxqkPNw6dnENI7oYjKBh8cV2NqbW0YTANa7S/Cew72BT8OCBk0/y5
/1fkBkHXg7qJ1SmlzTTK0Zg2n1SjNRJ2D29al0QF7vXQNk3TOy/UQq050IlGynmX
SHyjRvRoCWRYTjzIA8pfOy1vOYqHNEuXjBdeDC5L9p3a0/TKS0e/mNKbw05doJRO
L5Pj7TYydEOt9MtmBE+HzQVhtQsSEV9H0L4I8DwJAfk4OCsIMBEZDnGz8dvry5xs
q00hoUceylWM/8DPuQkDe6cjqFU1euRHRt3PfSZSKc0bEgeXM0x6iiu1ezKADMf2
zcMltNEVXTGzA9jfOgCvkCAeSCX4wW/nOK0zOZ93LAZanBfNV2phwC5n5z60+CIq
s0PPVpP+mT1MfxuZsCffLI4Ah/B3t/bcw2RyP+jZxW61zPrz/fYjhrAzMJ5wdSYM
wovc2Cu5YNUatmd4dqFhAG5KEj8Ad6JdjS08k78pNvphV092arBF8NXje/wkI1/z
2SkM1SU4nOQArtnB0eyAOg==
`protect END_PROTECTED
