`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y7952FNaHFQKvenvvXcBjC3QXLTlcHYlpO9fzjtctoXbPNLiol3BNjDkrIRR+341
T48jPUVT4IzfCGTPBNed1c2SveeJT0Mj/58b8rEYf3cqYY8Z4ZDy5xfMQshaNTYz
fegSDyX8oyhbWW8r/5uUlN6fQ8E+V+mI0cA0f1YXoEz77fppkgmwfVmBaNmW6NdJ
qKAi+WxyAN4uY+dLJEhc+mEIVCx0URJrpXz/nwFvYHzFMNesdxJecEtz9eLTsnHd
oKz0Ng1dh/sCx7qxVJVn/xWVEmj1zuO0hOgYyEzNRvjc0tvJuJxtNSWbhrA78b+W
xA/cMcDxe0iZW6+LczBTu2B+53+j84SiMFHry4gzs1MtsGSMZh2Qsc/1Ok+vEIrM
9O+c0V7h8Z7oVd0xFHmPsxs+5MeBTb7QLG9fsC4+GHntu1NFV+W/h7zSomdCBMXC
imvD6oaawdq0IqkLhOzT7FcF9VMLtUvkY08jsRzyB6D9g/sCw6MAbWZpiFCMi+cn
XRv4Zvs3n+y2UKKs19dGRoxOnIVWDfXxP453+EWsaiSoajwiA4ZcK8PS2CB6wemu
o8HpJZLSdKqHqRcqTenIZiD4abbqOlS+p48KksgbkMT63V9WxCWHsoxPDxhr+7EQ
FUK4eMC9pwh2B/PAqXkLRkLkL4zN9MvLB/kOeI1SM3D9QO4oa3ZDnL3058r/0FOe
XhwMXE/n2yUtd8eQ42A7+WHpTQIlN5oa3ESvBePBuTZfOyXRnnPXFDn4d3rFmAmn
67LntZDkny8FiMGOB6ITH4J8lRI94nCgPC9lBm7AJ51IguMbggDbs/O/5p7jepmy
MKN/JPuahGajRPwVssyYOcSjN6SJko8Pv+y+V5VyRMvFkTG9InDAB0eSVS2Gh6pp
cwEStMYu6cRqsFrNP9hGKZXKJAbJtQLPaTVDqfArjt14T7upmJLbf/exkr8y2zhm
3njpnpF7oBRgRfLh4owS3fUXzk9G/YdJqAAgu/xaQQYOobP34HGKV59Ed0OogqRi
WYI1ZXkE75yWFHnbyMQPxeQkHl55rseVOfxQjuNdp2lrCwnNZVeJR0HfHgEvCc8H
rN1ABym1M51eFT2OMxRakLv3bMgCVXPTT/HhwAaUyjCnzkn7MaDMCWpvb7SNIhj2
t2G+2acaBKEkKbo9D3Ex5OL0z2eJffKhdQJxqhWzUeJ+h4Rjex05p9SFJPU40W0n
T3MNxqdZ5CCeAz/nKSJsXM7wviDFti4upbGpakwifzenJO4L409V47WARaHelel0
8u8bZt0h+9j/txsJM1Cb3qUXzmRw8omx4Dt0LkPbiODSZXiHWSidzclunNpzDldH
`protect END_PROTECTED
