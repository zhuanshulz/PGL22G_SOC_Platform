`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zhd98g4KL2LssmJZrrPXJbIRjwHhA6myj5pqffaNzIzdCLIPnpumTjFMMjZ96RHp
qg9SKVKgMY+gg8lj6X4VOXuQasV7tfq6jVd10w7EaUJ7ATEps1XO4ksSZxgKMpOP
JhwGdz4wyqtfbtHsqtmIQp1rBmA3LVd18qqESZR398u1Id5PRFCJCdKutM+lsyQb
P1Du10PFIo0Fga9sUmBLapi57tvrwnmzbqK2yP9oCPkJXfEl/c0S5VrbkzFAUuoD
bta8HguI4c4vD591HXWwPhEPMctjVnQkSJMC7CqAAX7y5oHeCQXj5CYFXlyDgYPd
rhIHRolz8XcRimIxH71Sc2Lwdb3pOs1q1IgPsqPsUSQmyDzi+cCfFlr4dAlQXZT6
r+tPGfO2pD9RYMOYAYpMPlNzzPsFiE8kU3gkzhm5V1TL1zdAsw5nPpgo3wkgiNJb
eNHOSA2UaBxDcqkTC2tqCMvm5RzR5vfMwAwNETsaqcgrTBJI6vyZgM4PjtuJ2fyL
6km58FtsnzInIgcPz16H7O0ShgJc3UPo/RJEofuHQGgSNFIhuc/OYnWpaz4V/0V7
rlBj3HM/0VR80huMPG7t02OBDpacXlRUBqI6wMtE1gI7+IOVVtnsiEWnAvxtfazb
CpWokvgM7S1GwkADr2EH8g==
`protect END_PROTECTED
