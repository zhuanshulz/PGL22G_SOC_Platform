`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vbAHO66YRbbj2L8YJqvaxvlcw2DgOEh4c0pHnqBsRgNtCaHSyRo8vIXD36PdYSp5
zfw6oOQqKmqqZvM8Ok27yAa7F5JJhvN6/d5lr4VTo6ShpI/E+K1yZd3X6fg57PKG
T2rHShYFCas8tYN0VqJFFlPFiOlmkujJUoiLi2NAHGfDMsQMaYDn9sTR+ojNy8Uu
mPez0MvjjMd4HdN/NQUKgV5DXJ3XHNW03MLWN2QEopz2Y5OePUEnhSI1PNEemF+t
I/k8I1LyRlAvt+GtMsHRknpP1LSCARnPoN6Zzn16liOfcs/eby0k6F7vG9UTHNT+
K/dHZ0sGme3gL6qU2Ufjt6KKvhLp1HrrXLSM/wYztbI=
`protect END_PROTECTED
