`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wBGHKEeUnku7NTVeagpF1Kgd8W8IF1W4/FSomnBMWKYqS3eGfXgtmL93LFwZvdKD
UBueygJXQhLADIgrkRQGzVBQ+KfyQCkazXiW0dajshkb9ZQLo2vP5m8wp6CGyL9B
FYqHJEwn8YoDu/lqG21rHViR32P4y4T1cmV4EDmclbpICPKu5BbhWN8QGL5sfcoj
FTlZDYigIBe1WGg9GhhBMGg+eBHjPtocG9W8tqZ2/ZtyQZRfbZzTWgoFaEbS7pUj
arbBiiPeLqVtRQkqDcpLs6O8vFpWF1H6AmreZp8IDv+lDwpvA7X+wtYLujpQSLt6
l5ml1ZcAqt86bQbWxm7OjLvpLjUQ2VxHJ6oLT7wM99vapxDYn7uoc4kTjLnWV8YU
9FKjgKXiJUOm13NMhuGG0ObgLqHDBfaqBHrWwe9FGuK5V3tIGSTD8Em/EvnE6Roq
5S+Sr8WQxgN4suBe6vsu2K/Ij7sEm9O91yJ75l+Q2JAtC7IOpajzcsNA16zVQUpB
8z7yq1Nl7XuMoQD2GN/rUA1MeP5RtWT+sQyO4Q4m93o6hU34nQBin9y9WYDnK7tO
nEeNwjNwmbLWqfEHN3y+J8WqxQ/I/1Vrkh301p1wKEDp+TSWCsJOu9fCbv6VbF+P
/37N5/3seMtEi0KK4C/T8BXWKtfHDyYFW//rER/6Z2CIkl0a9eRxTPnCjlyYhbWA
kLdIVc7PhjpLwF2NkrOgedP4ssw2Z4web6GqWZMwfK0UW6xJMMrrUqRWgoTnrbBX
JaoE3AlHWyFtGuyqV/nXH28mzFDiTyE/OsvgljAn6c/O59/cSwyqDWVp9rSKGSMD
lWIy9KsHmmLeXUGHuD7tEnyvVJXWV6KnTSTyfvqsIYb0npVNSjh2Nc83N9O/ZCLE
LzGxt9QpBoksvjTn8KR4ymFRyIKKN0HPmjiNXmtA7I8Ak22vkJ9AVS4A7fpYfx/m
6dntqm2lnb3mGsiodQswMz9EnqZ6SsLfhGf4DIZkK+gtwVAkxTVNYDL5a8puXe3G
9Ou7yN4jTIITMNWx8ikFy1ULVX96iYl0IhFY8cFwmslL7bCoGwsP7SgXvjksh9C9
cok1D3lv4k6F4yY+2+wtkCPDk/7fPnQ4iVzMntBQ1MPJpu56cEa4NZCMlg4lKPHD
DkVoqZdNxbg3h8J0m7vnyMswPFeO5tFUvHdzkqZxPGMzlcmZEfFJWh/5dRGdFULd
g35CVqR++i0a5ekHcMLgnVwsagZn7vy5RVbDIxzn6ckpjv3uYg4aBpw9H6TWE4Xh
Zohb6fHMt3iJbNxkH3Q/0QWvDeBHr2f+zBf3mwyVNwHxQXMeetfjbAg2c6X6bC2l
7acpD6bs1IXsAGAuYsF1zFrzbhXO9FL5x1nFnM3bvCTS7GFW027zxKJBS9HZjN59
DYNnLS/HQb3L+TcYeu2QM0z0X20GF0ZgEq0Dzsck2aubuxrCsNnpYRaJIyTGXTkb
HXuE6Jaj3qZQZcdVech5YZwP9GxuY9Xe4hDLq2oDXhLvFAxzBuIdOKU0BVhm4+BS
bSIqqAf5NSHt3UFjbPkjEFrQC2DNN4shT5uo0CYhKrNY92X4Mg0NpPD/tVI2GVaG
VhDIvmMfSWXdjRgge5cvMPepvvIOgD1oIf92WVSPjnC+U0iCHQtkzgJ7WplHpdk/
TqzaTChxrCkFFCnWk2TyGLZZJ62PDlkm+igcSWJUVzbepPc1XZJuLu9yjUR09uwz
44rBw7yKK6KwEkVSgIUL0Yp/Ekhfy3SA3Jrd29E0vLbINsmWRW2fnAu4QQEkdONs
nnxKTDoSHBctk8Zae7OjqwHO/vkh+rL0SJ3KahdQoS6YUhw/XhGwbADcZ4KQR7Pe
vx6H2jnhxl3pOgRJUwR1wuBktNqawO59Z0Ul89gjgnsjz2zJx2riCMnIVfjUMKbq
JkxzVLN1hLbjXufM6NPd8v+F0ZcE1ys4yCtFevKmKtE=
`protect END_PROTECTED
