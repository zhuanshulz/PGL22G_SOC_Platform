`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NBdwePGmOMfAgNebzmurN7ngSeDC5VRxaX2Gdcuhw0VAWKdHvLO7D33LMSkGq0Pl
AoG5Hu93jQBC7Ygv+dbLxD+BTxps0YdxSfDCtFBtolHT/CgerP5QUAm44hdpL1Tx
QAEaRLsqXErCE99XKxwLK/BceRFK9l79BR/6quJbY4pow/Bbpo3LH5dynZ/hltA9
XaORUZam8zhhHtYJcTEAFJJoz9kWSfR0LDqLveos/Hjy9zjGpfQ334KbqgQufIl+
LkTQaekEORCt6VLsFxoRTOTBk6z8ymnoxky0rHdBe0bOmy4jegR4//pPqo9xmOXL
+4o7QciwUthXzLhyj/iB1hMfJYE3PzEaavW9hWMRcYTrf/W2svZI2yAA23LxQxpo
hB7kDX6BCKFwuAkv4mUDoYwKjWLBcykV+wUWFLIylfB8+LGymVmM1zoAqYPvsTnT
X9+nWSyWv0AtwMDr7D6vRWStHkEIftLI5dBDsBVwtXei9wRic8zaAKezpaIF1ojC
NawKJYMYfVm8wVAUS3IrSZagchcLBgoPaZTF4dJ/gtOyG3wh/hH72/tNokQlWM7K
fWlAfoj6im2sz/7cqDKUhxNlTSUnEqbh6WSI44/gwlfn/vq5U6tEkHk9L276T//y
bkHTujtJLYnp0Qed03YWI2ozEkB9OvZrBgA0urLcrYR967sQtd0ua6SwMQDDflfF
zDYUOfLVXUEmCdLrSLmz5P9CvVDyUEoKyzgYr9mN2luuVuqj4NbOs8CIUU1/AW4N
8nUSkH37lBxY/1Smqt6AvQT8PL/uQt63uoF1k1VhLtiL6Yqr7vJ1v/id6TaxzeFH
+sP5L2+zDVbavp8GrvahYrMgyb02iCh8sCCSs9Jx0/eCJyQYTbzigWjf5YzONKGc
KQxyj8q9yx1JZBUC5OyXzL0AGuOgRL1d0xLO5xHVV9QKvjaIh3h5xjj0nTXumJNv
EwcDU7dIv86veT4dgGuiV45GhxQOlvblqBVF1/ni7XPeWX6ZHPkJEmvRwr4Pc3T7
mMKy3F5LY778lPxR/PxpquCI04LxH/1uA21PjHwfQkVO+xDMvjqxhaf4Uwkqh0N7
BIUPW9MUq4ytSWYBBPFYyv7kaZLvAA8uYy8Xes7+hb6G0u3YrxD5SnsdiFKXFs/9
`protect END_PROTECTED
