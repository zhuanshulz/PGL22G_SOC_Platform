`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TN7bh8tdCDYv2irBxerzQ7TLL2NeW7wA3K4OuB1Axp77joonLbYlqIPsZYb/Rl/l
ERb5v5KuxmaiLa/Jh2DVZz3euI9i+Oso2EqQlbEeFTXDoUycIiev2hKXFH+jfU/C
47Dt8rl4YPltGTxFyWZIRIeK1JogHdkT5i1q1IiTkWBSX0uw1IQ4KtAY4eir9Agp
A72JM0BJBw74CTPn1jEy3F8uMkOMi7TgZdDSr++QA3R7No9+J4324fvHPU5OZ6rP
quatwlW9ak9VRRRBdk3rwCEG2OcoQCUqCFgf9/X45Tr8oPFcPoajzCuEunQn9ocd
VPw03f36VCEscu32sm2Hr2JyurbuAVTbhFm2hTVPExRYwO8M7ehldnyX5X6XTSMC
Lxl7WdIragQiWrcwNhUgckL0HGbbbKxn1/OdhJkefMw70eu+bK32Vc1tRUFQ2vTA
`protect END_PROTECTED
