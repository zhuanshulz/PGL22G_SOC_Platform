`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ojAzFYb0mZquwYnY8Mx94TRak+YMJ88gxxB2rX7mDRT/zvY9i60BmyTN6qg6lfUh
ExKVmWPW919eGKk+PolVvBvZ50ZdzrxPkWT18s5/WC1SplYlz8cPAGVgl0MbrXpD
ZzVcOw3E6BIgpuJdVSgNKp2vQdDdGq/J4whFOHyc+V2otLZgyovNlK2fF86fT6ho
wJZJgY1gzK6HyR63aRhuTEtSYQltmS66rtnuxxl/2mWDDYLSZpbEjqoPS68WH3RH
+Fa+c5091203nlX1/m8diZZJxrMd/J5GmY0Gwi4CZlF7gTviYqn9cY02KZvAYL9a
OJf5ylrHFysVLcro34WikveAKIKkqExxeg/VaFBAJijbnRK1MhWy5i2FBo42O2cu
`protect END_PROTECTED
