`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RvOKfTz9JgpI/3Quk1NZB5ttEMPd5GxeVHRwU0OZvjrPoGklOfiT/nXDrSeej8l1
0cT+Ez6MJX3RrwdBaG1nINlOwresWRmq2uHi5YyCLmtbLV3jgCkKzoLe4VgqRGog
NRYpBRv3+OHQ3OUYLGJ9LBzgyFiCpXTh2OjhekJ6tEKtPokbyLUSkg0iVgw2V6Y4
0BoJKiaWnpBkxw2yvTnrRL6XvjXFxzt8Ky9FGKeMYQ2/7p0GWUztWaSmbptSRhYG
X9BgNf+1Vm+dKMwn6LDBrAgvzwcOzvX7DhvVkhv+j6leu6zFeUYD/PxB+fb0dD9L
SkIR6ExK6r7EkpxA31tAJMG09rpTHEN5Fa0OAWAQ9XRDbPIK10r0LIx6GnCnkPOH
gIIEy7ZYHjR0JwLGaVDOVJ0GwnE7ZjlC4FtlZSyd4SIKcsgDmlpuDhkxzztxbLBK
1EALWDCf+hQ6IVqN8P2TLv3Wj7NRPWYoC3+0jAJAXxmqA9DO11aEKJn+nFw9RoQl
6tDSrxVixfYrdBqyMQ5kxt8vdyRVbP9RtWZLImN/r9H2KyvuRZUOeafZzb7+zIYA
ewVFWaSo/+K83TFrV8JfeN7KbiyrVj7LhcqQD271MTkCUSDybJhCHLEbj2cyJB88
rj009PwZwyF8nG6ryAbJsDr15p+zYIn9SuLMyL+KMtOy5e4DnAaWJdx3W2WpyT+W
QS6N2pP9tIe89MWWJv/SOLfEeyLOcprHNQQflI6unf6pZuIxuOfWooHamrFo5VqG
qJoXIet/F9MtcruNWcQ3+jjm4Uu3Oc0wbDMwwBPqB3lwnweRUzPbABK3uU/FfxFi
YkQQ3wvjkH5aU4KrCy0hT0h7y3qh0Opqu8nWlEvjtkDifyafNOuW3D08ADcSTh4O
vZLnNOSvuQkjOkbItpuIquxZUDV1jXVVS5Hi/70zIuzcpvp/41Or9nQcdVr1YNWl
BOyle5VVayoEsy+QcZAnMZfoPgWebJBxSjGbIjO9rKWo6xwo8ZDrv+RIZrZcThW5
aXheLa2d/T3S3qLb7Lwv+h7JobFokMqG10gL1TFjsZl3ZScsMTTN3EU/enduAvWE
knzs63wU/TzaSq8HS7NGzL0a5JRdMq8VFGQg9f7bahp2IFZrYVm6YVxg40U/FUmv
PfERfVP1UKlqCA/dorB9iFxAfl0yTab7X0UzM4AmCLBJY5v/mJJzzI1//HNJxlMt
jjSPiixm3MaFd+5gsPKKE7LmQRzZ+FnBVIqNEveGU25Dv/xH1jtIiCsAd8dfYCr/
mmLwE61CzPrQdypwl4rA/Y1VSfcBYwFrkSrFrxnhC6WJSMrXGg3NyVUT/UBspS5W
mXYYOa3i9Y/2Dkq7qafnIa4dwKECs8sNvpEuioQlg2nisl5U7sg3hihTn4c+Be7w
zZB59+lZReeBhTFOwYDVLMwHQ7LdvzHW1mIXS7/1ZwC0UOiR3r1gvaslmZqpdomj
/WkXvr+A9dMuQu9q2eQDD7Pg1cHJguM5siDIVFbZRUNX4LjxgPFjiGn8jkJNOk04
Zui1GcwWpi1O+V7sUebTBd5XaQmTmdVUR80kcflTgIq2fAv7aS2i8RBl8LQoZwbA
HtcM1vXGRUZlmF360IqriFg+CJYrRIs2r1Sn5N2rhdYdZKUnNZZjtGbq4r6wnPUi
x0+lRPbH8nmklpJCuUF9ZZzfZG7Ow5gWgykCqiENahagFhHTFuYJwXBB4u6yDrQz
JSaCNsmy3FPj6qEeOI/z44MdwzSIkYenBuRSLM+ONz9vf1QidE+OslTcYAeK1XyB
ldpCrZGQ0UAtOa5/un7Jms3VFh8fG/Qq2UrjWprIW4A3zVAawm+4lvif3K2BfyWm
6JTzGih4Zw0sn2IOaMs44R05k8P+cvYjQDz/XJ6nAdV+zLzYY09DSnrAkbvEQUnW
bojJkQ7aTNatsl+Yf6kUFyXutaqHSIG0bdMJ3cNNZ/d56DyggD18RTORmk+exZ6t
tmEQE79+nZ3iJDbeGThw3dMZopL9VNAmu9lJ35sE50baO1mIJRY20d6D/Qbpy9w+
u08/hiqSDbSgHcv/OB/3fqSz9uH3++T+E1E2nh0WZ1MTkwwo8bMu426vUnm6jEW3
3lajhJ98V1ZBID9CsWcy4HS6ZeXIhrLnom8QymCTI0bYEz/KP9gFft0YFV5xHL4l
G/TtkQfIqiUBDsr4SjIjNgFwiPJc7jxS2evDdZBrWLrRLvMBCYemzabD+mTEgYhM
O27l56D6Bpzd5uBFVNNy7YEQMrn/aSsrr+ZfYggoMGinyoC2DSFFx+OsczZp8SVV
dRwcHqfqC01U0pwk2QkbOn1n6iRQeBUd00vLbcOQAEGmaS90/doWM1lYxn0CMB8p
93uJ/B2pnSc5f/eaBg5Va64hv+xC4NpC8IGMwIB/Dwf3q3mnbvxwKn6RMduoQyh9
OhDG33Dj6XX9eR89AU6eAVDe1YCcgrtRsTkRbCdadaxU+cWkwsRWWKPAtEEXfjNW
H5Y8TEs0cEIH1GveZqyHl9nD2esAC909BhJ5X5sS+n1aC+VyVEI5L/os0VWxR95X
SO4Z9kpKAYoFpfhCj6d7GRXPhFzHkTFQoBLK07L/Fau/fmD0lpnUB+d7k6h+/5OW
tPxSfTHYGCZ8r/f5pP+zHHIVCCZ8FjAJBOjw4Herv6tpYQpgRE6mA72jo+WT5xYd
Z2aMndCon4HX+UAzJMH0tzA/1z6dyDLqRep3IduPuwCQBszN2MkS8/T9drh9PCyj
/mH7L4J4L13uwtS+llBBrI4ylJJcVNgkzulJKk+A0Du8ghHmwOnkeyvaU/9xE9BS
zr2E8UbEFeC6JbmRz9rif9/P7Cbpv+ehQ3MwfWPiX0YtNHsAlBxUqrlLID+H7i2r
JXk/0zIOEQ0Otw9j3eWRYxFeKA7quXxLRIzuUVh9x6XnSKt50XABmIVjJedzO+Wr
SL5Pk3TMKDinyUC9NNSdm6mXgoJSYjfP7JC3aE3kX0hL7pPY6yhBGCFsXor1LAmO
LyWHL5a0PxyiDupqpPzsWjcIQzDvnsa03upJBuQJhgsLqSrXLgM91xmjfkDVfcsC
zuRyDHnl+VrLc0DgwdfSTvaNXgDl+5uNW5Al1/qcncmOTJFQPE+vFUQ6G2TQWSKs
EKPW1fqeomQhckofhPcYt1lgJCqdq/risprlC9sroFzpaVgfvI62YLGW//S8XiZq
3WCsPz6fywelrRIZ9qsb6ArEc/CyOuuS1DKViarnUCsVcWERSQ9y0uKPAEEaqVAt
MfhgTp/fPDpD9n9kzzPR+MBaWFT3sUsgCZgcLS8gm96xRFGQdfRXG6BrlcZ9xbqf
2+zvLnk5MCaKcTjk8t/BF/21E9zgcsGtC/fBb4saHsr9B8mWVU3iUWISxtUzzena
sQU/3G6ZxRPIy0AMdLmLRqhQ9hB8/S0s0zU0M5M97W+0kcwL5DBA3afhnU0wHD+e
CNy6zwA9prlltzVHeHxVBWhG567YwJScRGRIXOok6z9KlSoDg2P9F/KByWIaOqJX
lcK1XsSauxaqpEddcQxdJirS2j3KNnChCR34+7VgL1sZd/YsDHyKegk85gMGIAgo
975FL7Vf4+4LjbszZ0vHBcE3qBQpreAOzDfXrIeNI3CyU/0J5I3JwWHgzRSctULR
ukXHUjX/iAbR1gra7rLB7JpNyqwFoZTn/seHY5Iypoq5eil+nHFholaYPbat2CBu
ET/YyKrND5TElRF26Lwc2XRCcndZAjYV3M3QIiMI8nH4olUnriKPgBsiZmWN5V/3
M2GKb/79oSpFO//7P7PiZcCJQofxyowrIztPr1PecZKlQFeAlmyZJ3K2o4d7zzYs
cDD+8OneL+ZHdfM+01QV6RUktuz+qVh2WZ0COljL79C7nDnEae5J7Ft7dg4xkCVl
J6O1W197iQrxQ8hlnWCcekkygmWeZcWpN2K76COmmPy0uPkRM5+OwoUHYjLViP+I
9993ZvwMPHhnL/iWRRpmsrN7RNmrCx1DDd+J3kHUqAF+NZ0XMgJRMJSVB2iD9HLB
9NYcX9K7Ny5siAUOe/REa9dCBR8FyUcfpNiZvrSaqxvEJgcRcI4NGcG+OT0534jd
OVjH9kH+WRgG5C6R89p/Pfgf+tnoPzKA1Jflr1rcgMLAsqlcUnzDEPtZgtkWgmHI
yQP63J7mWriewL2RDrIF1+R1GddhIOZvmGWwr47Clfb0tXUI29AQfAuwrx6sgMc6
1gEsSu0sOwen+VCJsbqpsgTZLg4boHFUB72qgAxqGXdispi5X9IMf40v0mMDlQLo
vnHB0ERYY9IvHABIi23pQFiEn1IGkygL+kAr28GOggjA/awzh9MWXfMoPs2UJbvG
IffrfFzv8ykfr2yMtKvSLEH8fu6PfJqa2NxdZZbHhu5YuqQDspcUIVuJjzZO1LBZ
johhuOZkWYU2rx4wdPi107GZOXq7cK9Aq22ekeOkHBxTp/0e89RnzyKaLopW0Y77
jEgMQzAKHF0vNEktiT9duVD6Q1W1DRWI+fZqbavnQOVFM3KaUt8K3cH8vJBK2Bqx
BsK9bt0Q4MNBCjFrlZxJ6oG8joGgjLnWiM/tOuLABLhQM01RQrVYnYtGGvOwlc/J
jZIVfAOoqTuF5V8wi8SORwGTciSHJJJ7OnNO19qW0ItbEQumJ+/g3z3ie+NazDTU
JyRRDJYF7sHw1adjR3GVMmr4I/0+6K3T3dEMxMj1yR4aoNBCMpLf6CCnJ9GZ7cJi
pFb1+YjxZY9zcqTjRKNT1Cheot/t6m227oKDW7U3lmi9CazKemUbrAH0pU2EHrns
ypMIvMIRs1/AS9eRJKJVme9W3CWqwFJP8m75Ksj96BgUYmom6DuXRDJny1iPnEqL
FO+pBsiAb/8yhgT5g8qgJX1V3AQwXdLePb8OTco2d7TsLqJ84X3zehkwH7biKZ0g
6TmVUM3HnVgw4RsF6GChlCcfPz3A6MXN1h7uSOh+LWl04wzUt5JTCEV4SapjvMpg
GNPMbhnPvw0M7Di1W42FhnROyMjdIV6k1w9GcKsQGR5VgsUClZ2rFZCcUy49Bfmc
oCl7Aj9W0JfRoSubbmHxFRtTTD05PrOoQfho0DSYnYo7SalnltiD+hVB8wZK6Ip7
D2VEaH66Kkx1ea2uL5bzjrc4JXvOWZFHeQs/x8mmksH5bOQSRR2K2Xl2aYccNjAL
xMXCzAQQzeU8WDD8dJtTQRQytIgKMQ7Y67+ooU+3g6lc7+9k8VuygXqrYOMhO/OC
2stmIOEpcPZ95kkO4qTfsuOLQ3dw750fuv4rH7A8jmcwQrqpTLxragXxHtdy5smZ
Pv8tCLv4LxwD1ej5cOfhAjtlgOxwFmHHpYIFwIxlmLKEhwQrZ47ElI4kCHfyhW8y
OMhF8zZmMah0FdNm5N4VAbBXN6juBPB25v/p8ZNTY+M3tC4p4C9WiMyb9uhRDFw0
zOqOJfdeKwN6MqsJZzZX9ImymeBftt/jzqvtayMsJFUGFWOh8bSycKH06I5yliyh
5mnJFH04bE/X50xOfV5pdrzRJ7mmQp1p/4cXB25CQEQv9axYw/If1iuD9sBqkxzz
yBxBu2tRozaRxYtZukwzVXlpQqSfbC6je/GjY1HFytZktehAVbFGWYWRx+a+atW6
ffwhergJdJJRWt1QwjovTko6PcbpesVbhLZv5zU1CG4dro6UJd0hGpq1e7sYbYPF
A9Qy7T6vuHBilN+Sjd03VtZznQl30nuH4qAw4NH8Ne1aD0O1HlifpG6PZc9uHa9Z
B7Dy/lWyqHLDt11rKJep60dva8qUAzmVgnbNCXRDFdLnExYkY2YQrIyxKosKPSg6
iP25DbTHdbcGSyTMhGI7QIDsmQ7sG7WBt6wCCvvf5zBcRHwJ2VkQTqbKIsNvB7ig
uuU94us1msl/fxMMPTj93dNM91lLNqhmNB+YU8RL3hIlRFwWgJvAjJU7/EUhom7U
1hIiUyq0mH5SSebLfRaDKgnXLgzO4wqxulULyqDQ2jC0C/Fjnk3cA/Fds7KCzQVw
bCVCE+Fwc2zEVPDwzLM4eVzHVUS2kWyfhp8hSocmQE2Yh99l9bDK0swkNAJPc55V
NwCmLnhorSVnEhj2IuqneypkgUmEW5oHs2D5fPiEWaaU20aTjlYbbnZSmUFjHi9H
NWrCtNkXrRTJ76eEFMKuU6saq9hdFasoE8XlqjtcZ/agkrgZppNLxAvnZ3XVLGvp
8enmM9H7wGeMjciaubDYnzI6aJTPDi7LSbM45Tk3m0Uk4OrfFqLaokU+yPVMFKte
46B3Gt0alVW4f36BLNA1rsl2EB5vMRE9PTd+B+ye20ADZVjNLA/scrXc8bYZToCQ
zcx8qo2xk5P4jOc+FRb1Xe5rrpntUwULION0Ge7D3oKsbrspPmErQBrtZN7xAj0+
VIkmuWRqm/1ayLBISIMkvEZPD4Zn0i6csAoeR5MffuRZrwS0H7CyrmY0jDWRyRw7
i/34TkjLF4UKPr3MLDjbZ12R3qAvqbIzT6Rkt1FolXfQMIhHRDjigl8BkDG5BUAP
DR6YEsQzqpcsmrx6d869u1jlNGKINlMAiCKREfmkUpshDK4GBCGwi+UNFUCmJ7qS
+aN29291hjb1h1NRyymbURqEnUHME0SJqRRI1Ez5MwP2cyK4x+P0GpIGjcaV2lHV
lpylO5A4cW9RwH2TxRxfc22ITU97JHCUPS0PJvUJJvP1PgLChyz/2Ct7XoAKcoN4
Err22dKZicZFf3oBQkmR8sXlAbinqCjHANoTN0rn3iFBwirHv+6BRdCjJ2OOaeBp
Q/MD4bA2pNH85X2+Zgb5GSe8MXQovLMAIubepOZMmQQKiqvExnecBJEomkJHSDkE
lQMxCdUmLV4FqCbmNlbVqZ7ujC20b/svYKGyujTcCOVdjMo2vTcW0AVB7BhuM1WE
el+zGhjEBShaVJFYU6TiavkTgvs6lfoWZfz+ArweN5Fx3sIWNgRcEYiZvHtr9a3l
YFP+KXvQFWug7mGOQjb5icP/vwDK9haru2JX46S7ixyJEsVbGImAVR+UutJDu/KO
cT/nOMk0dD+tD6Egktk91TOUIowvGjpsNSIWED0GMJE65no6vG3LVVfxghELmzfB
INggSuJS4f0Lhkw4XsQ0eE9/jx7fJBUiOcvB9MEgoU2a4dwdipcule0G8N6daDkL
Oa3hwT5HgDLF4mhCxRSFEt9hz+g8h0zbuQLjZWrncmh38mQub+p67LXbiCvihAZW
AqwL//ZAHPgSK81b/1cN+cvNz/RVxu0GtHiiwf0osOeMCYQd4qZXFH2k2s1Mvgla
Come1pBh8kTWHmuTaPaxNNus77aPFBe6E80gwPah9GYaJ2fO3OWddI00LBh8IwUd
GOlYXvouT/SdR9zpP0ei97Jv3iBXJFdvymyDMJVL5572ekIt0On0no1YmACfiK6q
KETu2Lw5quOv0ifgD2HsR9QnSWqXJ3qJ6el42Ey41EDU3YNwah/e/bIFpp+xpHrt
A6yBwUEumDVP/zpRReNVFef51pi6suDrGP3DzfqDbXJalQbCByRCsQ8MmVQQFCSf
vw0HxOvbVAXlx12jXxE8lq6CcegUCfjuj+3JGBMqmNJnpci2S+kqKH5ZEU+CNqcq
Wp4jRIr6DQuks9vKG1Crec/mtbT7gS3hF8VsNisirnIaWwbiARcP60Blk/0c579f
IrBivVLt9ZSXwGXDNWsfzQJixoppjgxyCCLMSFUbocsoWQ5zvCx6hnD8AnPcKKPw
2Oc2Nmrhv/PrtU+VkF4mX1YKPZeEUMOU3cQAq1HFa9urA8wq5RAGY2YonB5FVdeQ
Y3Bq0LnOPnTKeG8ijoBntlGDLu1qFXAWLS3SK8K3UffN+/c6lhAQk84no1yOmkms
SRELByn9y9/jgCP0GK9mZVfPw3Hsgc4WqbktOOkoU/F0yboYAFbEBjYwqnPpUGxg
R1ZrJEN1o1pAXX/6/DbOK4iTuGQnbsq8RyAKe57yjmZGg1jT9o1fHfPz0+Ebf4vw
bDqDKZzNdZRpyYQp/obkEBlwSq0A/J3ydR39xgvesyVxC35NzI8VQgqEFw0zKqUD
m5Vkom1Y8ramtfmwnF+Onc8GHpY/9ts+qCZ/v3Kcrk/djpEPSPhYrxZv29Qx3WPm
jnMGRQETD6UMge+PU/+Wfg/3E25VfZQ6mIMNhBbXI5ihw7cNPfwTxEuxt5B0AyF0
4n9fuPa+Zn0KHDahjk4NI3Fzjl2waSaXDu1ETCjqmS7bDMuIwCNw3yJPqNvo2jyB
0Agdu11kTd3RzbpNQ6tDqU5HTIhUNo0wpA03uGDMyOcLQj3b4wgwYMAUf63JFnnz
ITv5+hUBL2Xj15z08EMcOV68gfHZXY2J8+qGWIedJPzdMl/IYJIwzPdWH4rUBAl2
hzEdvgBWuiBH92eq2ZuPMmYRPYwiA18NsrOgmImKgPCMrSyWwMu9DkXJxa+QCpbf
s/kwvehiiSbEz4Cr5EnkmtFnkL0FOnc3rjbMXjDWsGlENKgjfjAZVWaFbpEChV3i
B8/CQL4IKpaIe2ZvVb2gV6H7uX28YSKlu2E5YcxLa6kBgUra+u0xr4tjtlzJ9Vyi
drfbq4nIxOIh2kW1PjZcs9KsicEPfU5Em5JWclAAIbhc2AI9pdS7lIaC1fL7cYm/
dMfslZt2M5hhM1o23zTl+wiwG/ovnSqNF5F0slFCV+Z5PtyPoK0ZApCmG/OBzDc5
gqqUvWJ1WXKSzVxa0YIPzarjXFwE1usD0eRlLk3iT+1I6zB34a/6/QTBBVkECbuQ
brym5CqsFlaaAIW3jnHfL68pE8YWhbTS8ubokX25goEwEriJtg2GG7SJ/uY3I5Bx
aLgNzHM5QlxnXghNxsaBNGCovklA8s6mysImcw/Jm8WlyA6WNQ+6eVHp5L3WhOj3
HY8j8LGh3kzyGvzc6/o6Lpep/hszImqTPWJPNZT7EyzE8yREGa5UlsB1EpSDWIgx
X7y9KCcmM/qjG6RaihBx+91p+39EAagjGTJuuYQEcHCxX/wzu6+xdCz6pdk2Hvie
wrLeEO8P540xPWsYoqBtnwLrWWK+uCG5Aw00JqLlbG7AVDq0Jy0HDQf1Fed8b9wd
7d2URqFSRDwJUEqG7AHhi/r6rnNq49ZQIcRUEwVv+PSJYIvZpCSj1gJIoBLC2pY1
k1V9cuu+dPAikIbZ38n/i4tglKrphF4RCREbTzg9n/vmlqSHGsgH0sll1nZcPGcv
eIzXeR+JWJJYqiKtV+uCWq4Le4g+fBCWiEsB+yVUThXCK3G6VrGV47Ryy8Yc56th
UKj4gmu8LG1JoJ9X8psDAfpPwM5N73gIcZ1K4Ai8tdB+mnE9G2bt4j5Ywmer9Vju
4umgBZzo0Dmyvze13Rz9JHCzEtN3NLMvidPy6w2hqwEqz2wlcVllB0Iwg57UDRcG
nYLIlsc+XmU4OnsK1HsAwQhr2NlY1U7R1AIpy7c4IYrADj4GKrkp/EBPYcP7fcen
zmsiXRtKShKdrENAYKpisx/KSd7MJm52r/bZCdrDHlNRrEX4RuqggnkBJi/jQPFS
Ukyfaje2j9ppTP5sr/nwX5LvjDFQsYpi9aNJWy899e8C4obTqI13cy+nS+1TmAtI
Jx2m+NbKozcA+YTzhNThx9PJXrFFEqCmqZW//BCmzJfEy0s1CFeWTwg2x/TuOyxl
iQy+5gxBthqR7BVmi4DpCqpF/DpTWozmSGus7yyLJ9ZBgRYdOxfOmD+p+nMSQw1s
EUUEJSK/VZlnosIgV8pUWYyVmUagkHDzqXsQbszZspDihYwUxI+FHyX0/2qk7Lup
NQujtq+TEqKTpxbAoRKa6QFFl5heZuaw2lQRC0dbRhFeEd/W1ydG7BYfhDGQN6Aq
O/ZTXOzRZrSmRHGPUDpkL7gOTeFg+D1vJ+TuAwGt1yveV83PS41kqyBkZwlhZ2EX
SWmpQRrhZSJoR/gG1oHHcIPKs5N3dA3YuNr5gNmzHXpGFepJUEojK0luXgy2sGxq
JX2WqytmZWvS6mrkvZa6ifYqTtgho9aw9hJ1DbcHtfqkpzb2barscZMrkzme172w
PRHVWr2UFFckS2KKdqRYqqH0UN7z1hG1aMo0eipbs00HJeMT3ROX0sHN0+PhfiUL
4yM0O69EpFKB2ebtEtEASi3eKLsHb/5E9hNPVkBImW0dJmmAU/osrSy2CibMaPNN
gyBWwJuJ/LMTY9CxMRJb1W9JUEX55h5TLKgpQ72tZPBMbD40MLggw4rlLxT259EO
x/W+6JDjI+kZ9DDAal71aiaTj/lrHWU6DWrmEyjOF9zS4HUhiwC8+fJusJx1FChI
jAwvDYidKXCDU0Q+EbArxJgnF2ySnQMe029E6tV/YljCnsNCcPWHsJ1hnk9wSzgp
UdR25c7OTg0DW8hdOUzbVOgOKlgK66lWvX4rLvC22R67m711/2BnavbkYJl7E37h
67nNRSlArEqJJWQSO39g2z8YPvzLZLvog2ZC5XJXfbhxC5Y5sw4AY2NZFIlz12SO
8170FVkXoRtBo75LAdgkn6w+92EGzvGMHu7J3RWvT34ZAcUekmBlckbiYqOGST18
bz0DjhxYqtT/SWOXxaoelXVKeiBJscKhfFhrDENXgqc2jN6awHHLNss/Cpd9aqpK
OAOGEqru8A9T6Vn7rz+Cf66pgHE1vDWqIrBbnojpaswcLpHPSp4XXPbOS/QIUGGf
FxMH5M5smFHtM4ZqBbW6A9M1E7F1AS1EBH5RlacjE27H6n0l6q5dkl3d0wKD58GT
D75/YS3efVvM/mXvkqy1ofuxlHAGg5hKZgcKudNWOm63j5hi5eKOdQooeIKSnLtO
7BWSS0YkSrvyVsNIAeAVwIa8csXujLgNt72jVlT+6OB6pwbC6L8AjhF32em7r2K6
8rb+eeuM1/3SK9ijZYJFGMLkj7Zbaj+/H2n09HPtHrQod/N2SamcoZRBNecsd+6p
yBEAgPkpoWf9eZBL4bTj5SCmp1wDCK6U9cci3a6TMuBv3jOLPwYwNf6xJjYw2Xx7
IEATBgzMOktnPi0oKkpeURpjzJ7JAe/ymptNzLaAkrOyAkshVsYouJF47etI2XnZ
IKGhMnCGC0e/1NudzNBK/AxVXMvPe/9YskITzvTx43vyKu4JZ+BeLLU3+uRB9Rk2
yw2vTYvZTmdbsfkMdTysadx3xIWnrklM2mfGHTEMAqbWRD++/yJ0uCAY1/0rRfZQ
zCe8ovhc4/bux5/0v+cqTm4AKFQ2n4CQ1dn1SOaTUjoIK8JIVsOv2OVcHGMsg1lx
W1+CmqOrj4JZqEn0Mf8Qy8g8kV32TGizEnn6RrH/CAXXBiqobUiTY+/uhWt2xvad
UGD5cgopwe1vDZ6YEvDBcZNNyhbVP2reTh2oOMQ35tEOr619UolUIcRNVjBkcUY7
6Rpx0vR5aNxsYSAgpSMiTkfA7ek1sRV7uDdKsDrRpJNsMOfFg0o3l+rIdGJeOW67
8X68AhKUj2SenDctwZ96ei56wQLgO0l4973IT2KoIv+6jzgZHoC8k5+0Xsz7u4NV
74YcCVpgwoivleBENenkfOYGzuf4SmkfyzdqxgZhz41T+1NUdYw17hMiVS6oUGLq
HIMnBFs9KsQyTBLUlh1InInIwTlukgrx1efE2xWPgufsggy5kkW+ghDXDGUfxB2p
4WU5EKhcYbM5OrL270dsmxXxp2aE9c6IBSa4/CFisDXlBtPw0e9MsykB2QXhQI4w
z/qRgOulDVeDnXxv6M3UEaHnOg12EqjKib1EHfYiyD0toZxlnETYYqKt+Lt7ir/u
7rnu2BUcqyBv2TJRvdlk9OF49uQrQ6cAj04PfJdRW1LpnoZzqXOMvY40Res1m+Ng
2REFyEFNUpOJYg/fvnjonniNJVZMCYG7wEj3tZDzZupAx3G1b/rP8thd7vVMI7Vv
eN86zVcEzveIPnqi/mSJpJaNK2r0Cj0iHPYDhhp6PR4UOaVsqpqygtil5b5/78CG
DvUb28FaE89iZ4QOkbktanaASoaPCKoQe/+Ga6brbyhcX64T+EjYFYF/uepxpJnT
EMr5o1bPysR8rkSIMAEDbvjfILr5DSqrwDIaSOZ5e2yq5bjN5r4wAZLgkyUi+rfH
2zdAgFqgj+EhzbYww8rJbaVTvqV8BiK6/kkRDGKH0lr4mcfCnXQgea2Nt4ttygt4
MlxxF4tsKqQRI2vLIkreHU8XCs23YA1U+KmLhwntCOxvJcdXt3JAbV319sndOjPl
vngaPni3MGXUfnUmBjtWjm1zumkbEwvO/eFBCix5Rdpy/k2dkcCdKL0iXmzWR++7
9w5HrGZgZzV3W8Twnem+h/TIpt6dDzAquXNh9XbsVn9BdPFGS8gao9IXj9JcONsV
T6kU3zhehuaZ38UmaUkwFQ==
`protect END_PROTECTED
