`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r0XwcUy73NlYHkAjGKeMqBXS7R/Z4+OZ08Qa7IUY2QGLvsUAMnSs2DTYXed2Ko8t
SZVnFk+q6EEplVaPh13vUe+yXD0vv62AreMpIkt85l6vq5W0HD7isqp60Ogvwbsv
v/fYKfMzxt3Gybz5oVULFFfk0dGL+ktphYtPwTmIo/6XL+nWZBUbSOyd2E1bnH0u
Q225wxHssxavSH9OuF5r8lEuV0dnX+ylaLwXBSM6dcB7K32/e6R9E+SnBtQi40hL
02axqt3zD08KR3dJOy9Dj8gi+bht13SCc2gTNx5eeaiq884zoCKWf8nZeN2chM9O
k7Cbuxv4DSTVbRHa5qUlecdjhJxQuFkUXGHoxMszfN+/220Qw5o78+deeKX2RYuv
E1l7uYnpmfBeH5P86o+y4JdC2GLkFHh0SUz3ODqAnNlkdQzagqSBj77cJeF713bt
oXaF2jOz/9aYTSBnkUmUEpfpTM0hYeWm2jFBTKs7uUSpf1rHzH/e/XFqOaiDCSSK
N/I5q9VxstqQ3PPjKMTdPw==
`protect END_PROTECTED
