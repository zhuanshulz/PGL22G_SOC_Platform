`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t7YCFOuRP/kVoJ0uuCUaXPdU0YmsvhrOAENEf1Lj24xjPcmxTVc1Cpg3F0Hk1JKA
dNn9+0yjc+ftEZUAsnEhTDBwU+hA/Drf+owaCrcFn6ttBbLNFr3nzRntXNplU5dX
sK6vZUNGULF6pSFrdtKH5/dheGI9GHMWPJokHwzv/7KIx7UeuudAn98+n9xeHZRL
Z+kh0wx1iCzb0jhFBDjT+OEUVcUVgqJS9T58bQzGZer0J0M/clh9NBCtRZXUhVgC
mtL4c7B5JhO77jhcxd0YZGNUIiCJat1Zye3IYBFdsmrwwxqOZM0IXD/BEF0jl+zh
pDVefxJlqGKfH3lkEiLjurr3oMr7n05OQQgkeLFE50Q=
`protect END_PROTECTED
