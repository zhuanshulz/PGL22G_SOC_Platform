`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vQLVU/uwRmh2v3tX5Gc6RrVN+WzlM+BtFn1wGCAzTHOELjZ2cuwTyUhSDoSgTTew
4I8Jx/QJBcTCpUxUo6mbFCfRHC5XX4qG8t1OTEeidvfIDbj0Xa6EIDwerGfgtx7O
1us9QeGZ/G7tU9UEGilPYkJX8x0BphIEgxCK4+127MfjamEVu/3ANuAQ8fCkGaek
SlTbO4i+nQbiIKLffjcxg86P5V4FkkZpasWMAZttXeP7RC3t3cCAfvvgEFjb0q7T
pR5OJohJyHv13tZp1QPreGbjCyoe7MKMPkMMSXkaAQQqMhPDvA50a8/fx+O9tkt8
VGLLKeohoadBYwMTgpF5ilrxiMFrDG2vObm1TkQ0Gp4dqqPCP4YNivcCUKTr/0kn
gVnAb7S8CpAVFI0DLayORnSmX2bmCahzPelCnJRe5nA+lCRXrU3R89eifiWopwTh
Hrint+JynZFSvyhU/QflSbTbtb3IxRCGAUrZFmm6eBfAbJV+fbI9ct4J+/2ry7bh
03wxGUlE/eU2XMlBS4Kz4vC/OXLIv8HSdlhrWv4dWDKQQly+egr/APExeUOfPCk8
f+A+Sj4rx4gH7tcoh5tSqDpqcCd3hZJuwFFpwZebGfeEbqfBwe/c9rbYz8ct3c/f
ijiGfe17dk48jknwC8M69BrGj+Ooi/37Jt+Dxdsx/q5URp8P1CJ3eiO3363z+WRR
PzHAK1LVZZTNP7qjUuLJX+P2nyHxq5HE05H0HNcrQyh1U/QXArJPjHb3nOzvPk+0
NcPSR/IJ/SLRMTLGQZfrZOezhe4k5Vj/WkxPIhna7pqNhOGrW6wixYJd3AKsfmXo
UkU0diOLylQolOfgqdqorndCHsqZ9+exehio9QiGzZgd6C4L2fPNMd0baoZILHHA
+Alnqq1Psz8Sb5qg7P4hQ6c/ROjfI7aLbvkpeZT5Pzs=
`protect END_PROTECTED
