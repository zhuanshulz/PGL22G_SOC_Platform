`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OjjE5MH9oLQvBhWdtK0ziQz9wlEXimJzuThQUZr/C9aQopiNt/+Eyf2aWwgH1aro
Ka8NA5JvHaegV/9/h3J1vlgkX/8Kk+LOLxPEPHKpJ0AfqHDID4fPV3E6X9fxUfaG
sCRfcATEiMcBv1o2zDVibORFbdVXHqU7AX0J606a1FqoUdh9WbuXjgsAzF+dZmhP
gzf6rhF9pjURnd0V+Hu1QY88c7rRujExCmntP4gbBwOumMpXm5GlQggaEyO7bsbl
ugwr4bHHAJJ/QZbzZ0cwESVtBaVyACAtvrw5A7WJRzXSFiHKni0NHEjsgjtmxKWd
hyEn/eIp/tyJ0/nqjboVNIZJJKWwTaLvC+1EdtjZpW4u++w1MYcINJybQp++bsoJ
izO1PxSefgOlhjXjvu2H2UFI4D5ocEpGa+3MznOhn4uhMjKwIwGN0MLr2EqEE8VG
8SDXtlLlzavXet9iei4K0vwVu0szWenG6jFB5uTTq/QjuaJmoDIKPeLNCMlB6T2H
`protect END_PROTECTED
