`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PnSWu4Hg4Li0CXe9RHzhv2LOKfsQ0TdZpBCQf6sDSY27nZ2H1v1SMfoZMbKRqEJ4
doFDJWFMCi7O3Y57EWzG1tHJWScLyzjgCyN/wS8e0W9PDRe8+A+43CGt3+uRcLEM
VijWWFVpklpnlImzPMWyn9F2HyMRwwuj5xl8/72vm+wzia0YpMOhmnUYwpo0oaEC
I6ey54EwEqSqsvwTHY7HcYGR9nAMimmlW9m/uaw62P03/40L2H7Kp6najTUw4syu
ozNVM07ZQDGpZnzzAxOyUw==
`protect END_PROTECTED
