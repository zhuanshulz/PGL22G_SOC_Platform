`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sCB8HRxI+wvP6MWvrQcuVAfPCGJdPNfjWV6ZYAMeMXD/U5FOx7ZCX3DyhA92YG65
Pu1LsMvsaukjAKwLF1zusjiQYWcKDxSGAzL4JB8FykMJ+HF3pMMoexzhPx+te25r
VUB5dcpc/axUrp+6sWsE6Fl0g59HalnFILU+0M26s/0FmgPKMCsX67W74kCyCm2l
PCbnaItJBL9xtHrg/TkLQmTW/mvJJY9qa3OiTxrnfb4d7GSegkeKHXhLHYLfC6ft
hxnXEX02JwP8aqdBeSYt1InyeZzysAJEJgVj0k1Ig3i2PvfGldAP9t5sV8QdATEH
6WuX28jHVyU+/OKByjkYkMImY9AmIdvp2Cq9lkpjgNd4MSVfOHIGc0ngRlCdM5N7
Ts0VDiesp0GbNBFg1kWJQamAC5fPYQv3FdoVGyAUfNi2koZlpMYUDXmrDx47kABn
OUraPSuZIPs0rf8ae1DTW5dMiNu3ml65WlrVpx2JL4FkU3NS3Fm6UtfODywG6quc
xqs1eR8TVEQVsMp9x7ZFQcTJodQhC9V4lE2NvbE8L56wi4eDLHHOxXmNrtlHtIY3
nNEWWCfOL8cY3Y0Wwfkp4JgNSfKXhyN/dDaL75qvbvLhYHBTuqdFftuZ7souAhsR
roi+9qzlfvzbE0TTpfxNp+A+VA27t1xWh7cqRpL6UeDDVnEzTvWeHBQKEFJ5kDMW
D6iuG35OHzDwT7S8xf1bXX1CaGpmNVqFx0ZqomCy/70lgMf+B8WPjjEFnUv2lLOT
W4in8KycbN6V0T6ETJ51qoxMtt9O3olRMphyXu8KSc4eLlQl2rgOnqUEpag9czfY
HQCpdRrl1dtYomVAmq5CL76+9X4h501H6/zf62Uu234wfC77SKmWTLGVPrO+gB0R
wUEVs/l0UAHJ2/kOA3OztPUJr6ViMFbMp5MWyiPK+ra1YsDX3MHEXiZGsoBSnHck
om83fYdyP8mJBz5wTGyBUJrUeXo1uB2ZbjZlMDnegPqk8AsyD6kV49hs4UcRnuFC
N4aOXNg05TWWX9WtsU6SD3ZKD6u7ST9yFsnafjOBHIj06j/yV2ANvnk49sCZnqr/
ciAo98q7bU7Xp6pP3byah3RT1S2Sl80xsUhcNeNW+CM2SiQa6fqNCZJ6vbeU/OwX
4WNQBA4O4WpluTXuC2J8+8plK6Vtf7SrwdlankSa4j6cHnInPJxHVVXVxkEv6YsS
cSyY5LlbTr9+63wTsjUmd87k3sJDHenGjlRRTxTbMJAcTohe1/CASgfjBtAJ56tj
UwR5L75qvrgJfjDOH6g9P9G00E4OWczh6NfIBzbKja6WH4OCgL+/ndT26KB7pOvG
LmpH0FSy8gQ8o65IoIqRvHshZFGmYGiYSqi7DYUoGDVSSowwWtS65aFj7GcSeWKF
yte05z7WNwcvDRCejmf7Z3/8HajZT5lEK/rhwRalTl95REhAjbYdwx4z4/8qeDuM
o5zBz8vuJDs88bSm/A2lxwohkOfBchwJzvm2EM6Jl8TyWOY4VzBf0onF2u5laPEm
3w3mVqr/kA2VCic678SyoekSZqKOMX2fA9nciP2y8TOOKcb8BJi4KTwyHIIt6aWg
W7fdMWokGP4fTW5mrLiI+zfml/XWb9Y0Li90f+NgKuhcKNTYIAQ6/NOjw3vH4WMr
4AdJ1J7Uw4YpZkDNi+GesHCSrD4Aj/B+QDPxhUni24RRBRrZ/SiiMaS9hjTNIzFF
Pd6qKKvsxpDNDlUQMUHIt/2FUrQKVUBvfgYQkBoNkoeMOdPm+RIgwwjRBg5SNDKQ
9yeCXpuy2k3nFwubmfibHxnTIEGjNwPeTjeeWA27r8H/GHpTnjlMGp97C1sYTkUa
lRN0JvM6jPWac7ZxY/bOn9SrNX/7J2nahqXM/06dKzR5aX+7YsS8quQyjeRfdlrg
5TvaUSSCMl33kqxxThjaCsY2YCHMi8F2VYWWxjePAdeuGpSrrRsssAaU5gBOg5DH
vji4j+F5fk3mRKzviXy8yE/m+eHpC+rY0VcrYFJBXiyPpBJ3QIBY0yA5tCJJB+/6
Uji4lt7xkfffNaDwEK+FMHQ9ei6b/82hPgrNDr6pEZWf1UUjTJ6OiDe0SOcQtzfb
svskFgwUFK6ei8KlS49sDrKFcSIhq+nWo1mtgwRMJx7fcOLUl4LSA+vrdyUD/Wn6
YuxQxProtGfjZ1C4GNT038wAhjPzWcI/t9A3LAKEDssHSm2kkngBPWcJEZv9jsHh
M0dfpgyLNdlGW8cwsBhd/+zqwdT+Ak3dkn+jctFhzM5+kldqncBXJZo/1f0dTLhd
ucn2g/IWlhiG+WzYkHEzX2J+TLV16wMyzhGwlemZH+wh4uShvGqsL/v0aghppJCu
Jf9HJys7aE7LXVKYycbKCWVTsomtDx8JJmtCLcHjmJIhfQXfyqLdxlVosR9fot/0
hf9wC4yRVU9OOezM++qTqc56OwjhCl1jwpzbPERtxl3crRaUycoffVOCInxuTxht
eH/t5oKfyo2Ve/67XderS4S9JpwycpsGyxHuxhCGw+hT5euPZ/vQ5igIQgXf7N4q
EsH74FYdCXIoqboujU/kdF2dOGurfTvIC5s2NUgQ6weLHWLJeFzk4TxRcbVeHKCm
CsLyf2lDzZfSuwdjjVnjtlFPTWDVeJMORVVk2AGhCD4sd+b069bM6OMgJQRXyPq3
KuyWYPSEB5BV0DQki3QDU3vTcbn9UDR4t/asiGXdz3i0y4oZV5+GgzMZEZ9whHW3
W6EYNTDtyYYRgp2PaqN9XJ1rSWu9zSKEFeQk0qPXL5o88XZ3/l4ABAlaMeVnBMPK
/oebTMGJEQ16IS449lmOHmjpr/6/S+XEIw7nJVaKDWTELwpPvn46TmoI1r1bceev
/ZxhhXtX3VeWXgRQ2nSoJgSsqE8qRJg6Qi4sj6ECh+MzMBYjWqNbe/BPAle4QhCS
KY1xMHpojeavGotDCGiZOos1r6ckTRt8siTMFx2l3GeFgzC0NP5sjMOp4nJ/yuKD
EqbW4W4S5NELQl4nYz/JhshIeP93ncoGq8o8Va6cRfAkFGIc1h/Lq9exI07amAuI
g3RRN/wArv08+Jq6J4P27ivAX5y46cOdoQEdyChQd9iRh9BK6XgGMllrWHziU38t
loY4qp5RF84jmiFRXGA4gsZvc9z9mkV3JZHRFu6leo9cMr9Be6t3Bmmo4dKWNoPl
4BYN5tS7zQJlPO7rQ+vSQp+O1AdrqjjsfXIxzRiGj/r7CV112LpHRnpgwGIM8s8K
+bWOq5f6L5fPd1+NdhrD6lfkh+rSL20kk6rQoCUTv7+qa/9V1W1/hj1l1doxzSVr
Z6bPTvYqcnX+73bAqoQAG3U0Alf7N3Yqj5mM6mptCnBVGYPnQmbpgalmZYiLkDXl
JOaK70LkxL6PK4rUXHVXL0PDzMFkScMLg5BbRZueDi8HWYGr9BRi1uE8/0WUD9Q1
pReu/8ZE7v71GZ1m08fujBsE0XgZy7nqSXES1ZtRZgVwP6d7r2yHjve6997hfS46
er5SWzcP1teDcYrPbzH17gWRprzvb8Fj/Fm8HhpJ/6MbjzkXtZgOzxR2d1WpllRk
lB9VZ0vSKeSEewQvaezRhAOGqTeFyheZ0N8k8rISyYh1Hg2G5XsZG4yHSz+ZzWmc
YAyFlMYA5SJKdqjw9JVF0mnu/rhB+X+9FjRWqvVlUY6qpL8nyhf3u5B88VyaQefI
4+NURWrWB4Mme0gWhLPe/w4Rcg4ukYSlGKL8d+25+69/ZtY3U0EFTBbWV8xk4EK8
y1RuLKVrHiBwcD5Ge/gE4b5Ld54t7k1NdWN2YbpFPNHvYoiXE0qCzr/Mtq8ZI0t8
fJLwmgh1m2LvBja6XWFQjNyh/9LI0+kGdg395u4JS+h1B/upqNHR7aI2w25rcwtz
gismFz3bxu4boHiIfOxJZ002ra2zcy3rqvT1rckWp4gVZouvBOU7Lq3ozpkQ/U7q
Hbe+Cz+3t+5kOcQn4rIL5IzfAdbM3fK1J7SuPuvH0gqQpT5FB8e3MWQEuh7iFm49
oSixYMD2f2ZAPH3rqkLQZmsA7qHhV+ZTffW3bh/8XMzWV3XaKArDKDlbKubv4vSV
l18YOsAEabmZahhKtzA62Xl34v+oPoxP5JkZObGNdI4r6/2ccyfODdd0pucbFsVD
2wHLkWqIN2ERVrVtIDx79S7OlP7zdfJ3JVMN8apOlX4r2ii9CmHscqgC6NuSg+2G
9/JV6sfFESarxb/pVtkFcyiZda4PF7OFUo9NnrhN+/mYjxEUJu98tJhsl8Zx2OYh
bUZTBbEbrz9Mz7PccsINptT279wVhoYO1Qx7XVi8+fy+s+75knogtcH0rHbgm8tG
TLfTJ8R4U1um0xVnI7NlG7s3aGvnsEdlkCoCuKuzi4piNdj/AHYpU4xGCC3ya3nb
xAXJasCgyYqmT87D1ZKS9+NaHxvpV6VEazl5QwYB08clsfvYJYX61LSIGwX4gmjz
IO+RxFp5TMzqepgLXesqoqDozzGuJk2ucZfjaUmmiwUiQEz0kNh91g0wJdiul5jk
N7lRAtGJTJDAHOMQO8sVgk0SV5FXb5BTxvG7B5n4+RzMaMJ5wk2iNIywYsRTkHXE
awuZqrsGlatmPy7h/35pqnGrx35Kx/kqtzZIc6oE6ogkP0binWhniJLzfl8DX+KJ
SXuMo95fdh7KUsI+/SUJkCx43z/2dO6oMzkjNTpB9Zcrb5os5eHd5RQgnJaPAaLB
kTJDT1YZ+Z3ccpr4l45dMqlvn16LXyExep0eoSejUX3UWAiMJgMhSFYo1epArFlC
OCoDrchgUUz1s97sEdOSjDnhWRUXudWsdn99T5xgoHzMo1nj/hqZFvUjCZvQtIG1
lfcB1pUMf6DYq9QAyuOHA9XdRAV0fGKAY93Lt771EHNaCuCgT0LrrcsWrDe76XYB
ouYjhaviLJQUnmNPNlW4spEK7PVH5w8V8fZ7jgBVFENHyl5cW747V3AXLo8tWUBh
TdEsKU8TRkozZumelO6R3euMpuFovMEWMMzYJphMGHPrVqN2u1ws0YIxQrUMud+A
cAV0eGMllkTmUm98qz7fMOO/Gj1Sj/qb1FSrSRgkNhZghAydUQnA/WHIxNC8oJVz
YCBnZhgtguQ+wwvtiP8mVEVDkNSGelm4/qqbCWZx0LbKfj3GLijEiQqY1GC2GIpf
JNlkaFE5ui1wanSUTb93VR9+YPQ8c2WVqs5dWH5zxjz55eu39w3YQwuv9D0jvlk2
DqS3+4Qgl2x9qcaVwPvB6QiFfvElgqwa6O4oeHMu2H8jy41r5afcJxTs3o5yi9DW
F/yvCIz4lxHVYzaBXwwB3417cMaVi406FZrBNztm27pN3bKcREMukA78DgyQ4yDA
Rs7cmP56S4MZf4dSmjVEqEOd3/xOuftMCGgBk8trqKMvjEHZJuXvWcXcf4+i7DcT
SQ6AEy6SuB+gnSBOLHngpk0oZ1Im+mVH/0NKfdf1rmxtfHwrkSbJThZv9XEa5fJh
6gs3o1ExkWe8uCxre1W1mRTkNkXFRV5U74whNSM20c5zNdBzJjQquPB2Eg5JyWUN
5CjvNGa1STIUWL/XsRiRZ57L822gYm6B5IhHEBK8Yp963aqrQN83FgDMH2U7iYQe
1N0QyOWPA8zIkzyRQL0szugBWAfRXLtGUxznVpsynyOzISYwq5mihftLZRJJJbLg
o+kk/cx9OjIhx1PrhcFHETebJ19VT5EgK9f0/+C6pmylDpsWi6Bbi1UVn27dtgFU
xUhzJkWzHLWqgnMSpzQ3d1+tvmBTZVTll2Yo6cZYDjQPe8S7itMQmAeGQa/998rS
stf20G90sGC7b+4A7CH0pf612IfTO+JUaz7ZUh2MwLNqu+EAFYpj7KbzPck0RQBw
Xe/R2/cjTOJblvNEdFQ+z/3ZW9yI5q3/7x5blC5XQeSnMNQjrfo5xF5zDBq1Svx9
dJAJ8Oj7WdcOyZaHmr7pdrwXUK1hQqzb4D1GKNzqI7mfzGCce5ArEMqDmUTFqnEV
FeHHZ47cT3tbtWKO1ToT+pEaVoQSOmxMb/YalZZumdMnvkxTnvp6p75qv4dXvsnd
A7//o/H1DYUu5aeYb8aeDKI8+zxKj2dN/6+IueKuT23gT9GGlIskb9bRc1G+hCX+
sf8rV7rWJSbKgV7RLK4T8Aq0RxTsGNkj8aNBy9sdXKwa240xpc9nBoVcfbdKms18
JKRVUZtMR1cG1LFnoyHg9yg9aHb8UxxPUOAMWhAAjRCKNpyHsL0wUASVLJtR60NB
TRiCk0oNR0XTP/ROQIsf7sQHbsqEv03Gb7MJ8aO95ebQfUW+WTpjxl3I9sMsyw6j
Bp1t22sPTWbTMYF0XcS3k4oV5GOtQ0xXrFj+JkaXXI5NHck9Q63JoGNd09p5M+fs
IZpTW60XYBstomd5QC/zAtPDfISOpwzDswFnYS0hFnX2YP0Bqkapl4YfWra52OZg
CgpVYVxbLXuSJrXBsa6d3iN4la0Xwgz+GEb/8QGdZqCdcqRHzRZUbexIae7sinwf
xyUVnT2XeZKWTRzFHz5bUGLPxToKwuVoFWtY+kQWClXWAiQbNDAZoSIs1C8N9fFG
2URXy796kTew+b52bclsP4EOSTdhF7iGMhaVAF6rdBy9qW7Fs54JdP1U7JvfzzVX
hTeHZyfVzAmHDlyYuRRrnoYLiMtbjpzIbQZqXA8d+ExI74XyzW8PcFU9ROkrQNCm
cWBGBiYrOH9nRnii9nfhlRXRP+O+OKd+5LqGYU35YcuzV/GEJwF8bror5hyGuxKw
/K8q/muxg/W3DBU5nsO2FIBtI/KZg2LTluuQpp5Mer+nxX4sb47uIgh8uM5DKbim
CSD+PSmev7TYLW4vP4Sb7dcYVhoi0OBSo1BN712PHSizGolMpwF2j/Uk1hdyNlY1
YpB9iDy8b3n7FqLSseo9HhXYOtVLOylchsQhA8JfgVqiEni7bQDdAHDhI+EudtDI
LtnKRCC6fHBHVAA9QaLvarf/I5yxCYydSIXhU5Kn9Hr3FO9vhGAFi7Sb1FsU8P1m
b7ZDt3bt1sUFV7G9dGLVTHRg09wf212dqhgNG2m/GYNqC/GLWyeLFG3HQLf/5Qw0
R9ppfTI2dSnTym5qjaUbdWO/FxBLaEEZh8nV66NElwGSehGTpDo/36herJ2KqB4s
1c35gGWGIW0T2dMIx9QVaNW6yHQbCkg7KcUHsfsFYpt5iuRrMdk8svABP1XUvstK
2sPvX9MtZ2mnx1bmz61MIBa17u16/1SEQo0Rqis0vQQ1FBeU/pzpLHvCvIm2pX4p
XtG+/3ku+4PCNgBYLIgdMkKv5/7evqiK8QlxY9J9QUVVzGk0b9SJhMW0Gk4PMk2N
TWExwXN3+lSoUuoythqgfE81V56/xmgzin0vZmgp5d6xTkoClRajkFgl69vSV2ai
tV476K6PjG1j+Ix+Six8hg00r/0dtB0dRVMd/H2PD8vEae/JPu2YX/C2v08AsoMB
Kt0eHRKf1jSaFWm5L5Sk8xddpR9PFNvJRInPf3zWvNcVeiip6f1IplL/iImG5Ro5
JOA+VNSov6GkGI6Nhz20JBOMrzXtVGOT0CyDvF0pUvp5LDukd6MasMow058zMTXo
NTr6Zw3z6x0/eYqpCobz2biCBZIpc4DV24KNJB4KHmvYsZ2tEqREVbcyfiFp9xS/
FtD5DVgoCDqPmlrSc3NqE/Xlpgl9ZOvjdVNCt4v3B89OgtyQ6hvyBzU7XZnBQ2fH
0CRlZPB3ih8ZHmfhduxNPXQwMevs8iw/vz9bl9eFeiCXfw0w/lEdAgHvF+Vbq2ig
h2fbjztyRqi/zWL6vzusyWJ3fN0paEDGhBikxVFrtHpr+2sYil6p5GFCjy6GZOpP
sO1UbzNKeC06KXZu/51LZ4/tB3brG/4/E9UBNAg1zc91HzHHZMCrwTSma+q2TMch
y2uOFum35F3xe0+1yl0Pkk3eVjHwmx7Uvtdo36/ugUpNmjdbkw8MutTkOMI0Hxhe
VuX8Uyee+UMSbaK1wnJMntbVQ5aXyGfFlNheEbIrZGGViR9X/yWmezCU7sw/8pCK
5IzTzlOMgGkkcdVOE3PeTVSC4J2P7QA2D4THbSst0Rn0UKJSH8Hkc08mytEvI38X
lj7mCIVfzVyD6TMP0puJgeZQvfCJ2c3vkPD36POHankNFmP8MTCpWJkJyTQtlku3
bgT1tBQs0zCf0T0zdaulV9jctAVzFmIfT6vKy/n2IcARl65pGaBYTqHPLmQ75zU3
XzZqH847dCnxAdmBiHGbgJujyWu3cDOuO78T8jiqO4I9xVlg96qcc9ZcxemLHhtg
4hJNVkDVYZO8Pe2cqo19ouW+9CNa5SnAvyYQKeo4WMQM6Bmj1DOXw+WXaWKjtd6y
rK6k+JJ0cL+STySbCiJRax30InrOsNbMHGN4CNX/LxyRu5bdua13iNtAoMjNa2mS
ZWPz6vsVSSd3XEDuDz1rAIX50x74HSYBT9HNvJqYza3uer2OlF3DDkzp2YsC5gG6
qvmQy67KuRAGYBPlDmvP5LikDiid/fU+6F7/x05IrjrURCRLW3AhkS9lfzqBjYJu
7llYTC+X8QCGofhFGo4VCPqDUuT2a5w2Yc3r4Hp9r+bWvr1NIR1Jf1jgjU9Lsp3S
5Lv2stoNN1YnqJB6hRll/orWNq0aSOB/TUgzdK1436jJ/6HKZcZdx7N1lQbpRjC2
wxtUNHGE0D3YAEgrIlB5CgaZvsYCBjPLSmWLm1cvafAy8w2MTUAv6UsHKAzbffnb
dPspMrLx2uKErZZlP3X7C0ALA2KObNEWP/yAsz0zFy9YlGCBD3kgqW6GFtIovT6P
q4NKOT2KmMOkw/8XvldEYrJ58o8xt23s/Sho9B7O180rf8Lc84Qp4+6g6j0GSeo3
pD5NbSAyJmhjiR2Fl5XHWr4wid3xONxBAuhDlSMyDNTR/0YwrSfsCpy3a2GHIW9b
m1uYxOGt5iA93DPuQ97Rbare5TkImcRZ2PCR1VfASVb5pINfk1ByqVqCFLJaw7Pk
rIzcQe2EtI0ecCX040WXkPvUCmg9uGyGaW1TV9sOW07ldGnvwx3mUhmCi5PkzXpB
bL+WHr6Bwc1PVfMTyQsF2Vf39fxi10stRuVhB4FeJl32KR4iSDqacsQFytn3LtpK
ukyG2jygeOrVtkUfUPbIRO04TXV7pJSqWpAu8OIaojxxWssOfnAS8/Ma7SRXflxe
m//HfHqUcJ8tMfR1rsF7h1K3EatgdoBwW/eXXOlJX1Az8WEQMyhR1w/kmPsLt89Y
v0qY7N0xfuH1+AN4SgCMi8FomNZCvk3b40yJ6ro0NWbnGQX4JzzhS7lvocqBgUHD
/S2+2QYZJJMaWekCNM9wHV0FFv8eeQg24rUQHeCA34bjIaFIkZYYpqqIQOqJe09Q
pMEtNE5gy3AkMb/SirxEQqul7kLnniNk/J44FkLrCi7/HYjhrLUZKYqCP8qsEHzk
IlFsjQoWHHnsASeEPgCpdt6vk8LQFBnCqKh30QDnyZBkSyDkE5zlbV7obVphptdc
QAvmiYI6g8klrDZ+g5JC1m+66ABCOLL5bC7KSM1/EE+EuTsszdFlJkWWRq7Aw0KQ
trHgtcEa+wxYx5Nu95L5pk23QlhnQ+zy3n1pco41VOCfmfvNoMWvmp/1OlIACLhy
HKEWVBET9fY93fOj5Z0+ZkHyJ9F7zjf5dhJ33bDECAbj/g2rRFAVnD71aica0Q1v
0lZOgDXXF5H89IwGn0LPAZdIZWn3WF8RlcX/eFfJltHi3BKQTp63gAO4euzIRchX
jAKoAZ7uNv5Z0jIRzdjrTIWKk2YCJDvZ/psjCS3z+jLD91CyipzGNNrBZTOV7Sdp
IIlEi1JLbiSELjOW50Z4340MriH5M13Ud5pT8/oTEIZynoSqPqtb2dVC5sR793U9
Nf5dE7WJd0pHmmUcpZY0suR/Ro/2dauohQR3FmtuucN+Ae31As+DQJUOs+MPRWSv
HYX7njnLH9qEda51QZuXxPLLx5kUXUBFMIgd3BkXZ3IHWypFO+dOdGndKUGlrkPX
ZBoVCGkARe4/a2XBzm+M1tA3UETNGJA2fC0cYhSI4ljr7l1p+tL1aKtur1aOqU7s
NeUI2tTTB+6FZm84Pg/UMG6fUr84SxDpwFFnDdQpnaO0VasXLj98BB3++lXllDwH
fQLBDqMgeCpD8RtZqCs/f5Haf1YkYdZBkAtmt7kyrLR6lohZpeQOfJo5M7DPl0Tu
sNFmuYFJQtJfLeK9J7Yr63NaaOQizy8Ov6lTAoMsp/OH2Pxu7+cmjhYZe7jC9bWS
c/oV3/vfA0aQmiTm2mPGbCUxZdoqRV6iB8pL0VT4T0j4Iz/99z1lQD/e5C50pISX
6YOWz6AqdRqCFmhp/sWT1fzsAIOpvWO4O48j966lyHN9JbXckn/K06uYUsBbVcaq
Xfvs7U2a36mWvaKCrlD1S1OQgg20Rf40n/EzqUKiYwuWyLlUClf4Nb/VpbmGN3WA
Zu/6up7S4TcTdoffI/za3qDYSQsDnJJtPqXy1/8UenzrJ1PbGjTeFINLMX0d8oaC
Esc6dCKh77tsfQM2nkMkk/lMwWOgqoThni7hDK+qezpQtbBO963sUz0W2cbCtIoG
hDG+2umwuzBpctLEoU3YLVqy00otIgk3GKeB/8GExzeEKMMgykkCUocxqeZpyfKR
r4kvKygdzZxw0DApp7FpCVUHtgyJzPEknt3QMazq+k9J71myCE0QhVi8FCosn+2i
g+hCdc9eUXwaTfyyvLAHYd7EaYpNelcjg8ONTEvTw28wvAEk9AlxUzi9cwpLpdBW
VLJDhbboqylOVeXefdRdmKOyBALCHEkL31ScJfODDfOr+mnpMyMZvi2zCiHN+UmQ
NLhoIS3SQ4xVOV05mrC+d7ydfkc+HGJLCk5Su/QowOAYqkDtfjolu4Sg/p4fInVP
h4e+upR3o+yDfoywtpML4a3Mp2A6xJpHNB0flFcWPdzJX/Q42tPH2TGbrycu2Qj5
v4L3e/zmyf0DCEypGt9IpOiRTLeDwzzO8nS7qjQFtVWhULpu/qoCzEOB7Wg20tm0
7dU5gDnUISx0LMc80Xf4cvF0+w0W9M9a53gtW8Mp0Ea6QtXqjA9VoxWuKg2MaUXa
myUzVw+6llxbTgnOAk5SmMqAnMUNPIInv9MSR7RGucPNN2yKqYL5TDSw4Z6jSMLB
lz5CsfRAf9eUXmfIHKnkA+WyjgC7d7nYyvvCrb/3lnseqFrpYQwt+KC6Id0Z0MKT
SszanBRyIuR9j3VVdFmWaCOh9NE51dBE20nlQf4Wcv4j5eCmzLLL6ozh8StauULS
OCITfhc4edCiFqhBfcEd3z9eLi4tWObCdJ7drxMG8RW+KPcks8R8exau+pwjXj1i
T2cI+42HnRjJ27v6zEtMpOtGkjIlZNGl+K433frhVaN4k+V4N/Mq6AE4uf39G4Z/
yliMoPCs24o5R5Iu99m+Y/3kODjamWfuz5xScUjENjXcFZOAAQWLsPoXeHgq6pXN
bTYswSNHzm5/2gdY/dLMcPP2F93sgCfR1/kja54T7ESqFoyoJ+nyfYwOEByMmwa0
iB6kpj5V5PBxvH5Hr1G9BdIftbx5wupFbsPDZ+lNNhvGYYPuk9j7Cz1prp61TBNG
W93seZt/PVZxqykmQrVgp7ul6tAo1LNQCaAJoDHL3ITdR8S8OtMk2bLV9zThWQBn
V2FDWluKVFmbKpt37XdF2ZB0y41LQZBYCozhBpcKZsGejQhmwpapTlYIcJDHUtn0
OQv3FRYlBOI6vZGZqI74CBVoDoGEIPx2Y0vaf0Gj/A6PweqqxxpmFbh2BRli/acP
K1yc9pnTD/qIvllh2pDhK2qGmuW5bGxSjZtYiKW5q+sxJjSexB8SB74jyI0OBw3c
a2SvF2412AdvdVBMi96hHUVKAzEvAcXbs630j0HsxtCkH00DMCP7hSw0F1p3FoNh
ezRF7OxwxDY9sJMmf9kkeioeI2oOUvmlFbHbIoctRoCHUndFj+0rgtidNgTGCvHW
V5JHsT/pS+wQqx/xTliPtY6uoYpOap7dSUJktw07yrfDQCVctoO+uRbxkYBm6Fl/
NMuBOIhFbHDwb7k/nx5D9G5xDCt1fVuduje8Q5hnVPiAF3HXErl4TEvQJZiiuFIg
gIcBWIYssrvLXrJApG5mXx6ik3Sz4+T79SuR6fqOWRPS0xVIIdqdKh032d16MBdd
eyRg/QmxPaErKs0J5jXs9WUTIDiUZfWJ49Rd072KqHT08cOVQ234tb/L9mqaqSjP
sCK3x/551GcRUz0F8kFysOU/651nK5Q1qplCKJTME0Ziirs/Z8oy/KuiLqui4b8L
o0bWVigEwQrb999s3f2jxlxBdUQyewWRs4l5fuFxN96M44xKV0XsENO4xzQ5ZXCF
Q8LF+Vll5VKXLkIUc5LpIGXIrjE7MxRzW0jHe1wJAu6Kf37CRBiHZNUv/Yemk+i/
BMnpp1l+OatRrUMrkQJ6Y5X+XG/i1U4TVuFlQPp73KufR25vr1FAwZYZpUEpQe8z
lBo/bicRYqGALSLR5y9VmFUZPrRl2agKc24DtwcQD9A5Dw+xCl5B3sS/AWKViPAV
T03rG4d1bN5d9wiWTaGphLePpqpGgtuhXZ8erteiS2sChFvB4ZRrvj9XiRF1ooA0
HykUmbwsJkGUGGrJceMLYcWR49i40MaNPGVI8eDlOpv03IATB19UU/80oTFktm4r
/CO+ueaFxsLN3Lv59xJDnsShDA4AdbccvgmUapswJRPolR+wPR9J7KKTD44xmxI2
oYDlwE4hbwZCzfx1Z6x6W4tl/Ht76jD1BgKFRoGKJo9CKZvF68yjVVFwPvJz+/av
ke55Jvi4ZLe+OsjGwqbOYbDjdp9Q4DwvQ1Z8qLMXsFogxbFsouFm2Ji1HatQLg/L
8N9yMCDD1u7y1DkcwWKqHEOu5EEihrJ3M/iOa60NiuS5Mofjk+QVLZD7Ed8+8i++
QjkufM/oNRGBya5fCsS8oi1cK1Cc41YuTAATueWkM/AxLytbxn0lK3oc1XENul77
Kd64EJ5v6gmJqI3E8HT5bkG5QtyVum0aNUtTE0wsGRqCd39Nh50AZDCZDSZgsGOX
ZsopuuSrh3OtTUYgfGTM4nnDmI1OXOQbp8B47L9ZgL7GA0bfzSMPjkonVZHzC4m7
Rbhm9JckL9d1wvlVJW+ieBGlsmXwgBDVbUCbg3M+NKMgHefYWCqJGRb5n1xDf/8K
/VyovRdKRDNH23sHo3TgwI8ain7l4ynx1NRhhVqqwEObakE57c2dluYvllEdHQMu
ZqjK0GxrJhn/uXnglmyvo121lIspP3Y2+6DNJ9rfA8MGH5rN6qzDrhM4I6Fk5iOS
Rj3OvkZLQUeCvqG1icLGZhA6mT33Zm/ZFpNBmhn0lYltN6RnzZNukQxRWBW4ovLl
ZSC18SEY7Gc4DXAsY9Ws0lJTKRuI9CAJ1iNbQ/FyMomHstiyWrT06GXWW4M7JSlz
aWrE/SgvJXsgmDuMtt8AxTaZvhWOnvMxqykTo57PPNncH4IA9cGd42dR+DO39ZDg
35QrzlkibGykhUkPGCF6bCQl+1Y65AxfodKs2xeGa21ThBBT2OS63NpDujLsw3p0
fELYNDykSaEjaT06a2PXBsVJyIWEgOzA3B88dUixz0VbHqYBt3dboctzHgwK+wHK
tloNy6vXaQii235f7+RXpeTQQg20pPotRkWrdk+5qekXIntCjMW2A9vsioloFLQC
9ZyrL6NiqyHGE6/KKyvRc4gu73mm1JHVZVJPjvAMIK9vPC1k5I1xZXNEjDyr75ef
3sae/kjO/EKIB9zugGyCwspsRucUznsKYqFpvjnKnXfHPhSs/ZloMB0oygiHJeA8
Imo8wng4i3dSxP0MbdykNoz+dGmOFY4VbpRe1HzfeYIEu7L6aE8GXZzNXFKZR5Js
2AVvJ5zxGdLkFL0wjxRr1SFDeoeJOljzWYME94welcoDatXWeeYpe/2FdkDqTyJ/
+iFLaltOgbIghGIorOr2bHLMMbChmWA+7uC1erJ3MhpIQLodNMwhKSV1qM3KagJj
fvB/Ae+pd9Qln60aW6UZ/++XvNNiXy3a3L7/gj9l32sjcuSx/NNI6N2q0zZEv0CN
LYBdElufAkkCyTpwj9QXDdgSe45zvAh4p2TO+9MCjVh56Et9iLy/5P20GNJ3D4S7
Nv6XwIuFPI9R83koa3rNG4WnRWggyX4XyjM1LTi5EX1yYbetgRf+wV7D8pm9XfRz
dFqom9X0uHb2IHapr01OAx45UL/pt6GjvT9TiVg7eHxUi92Vm5OwGr6iJbw0xX7z
N2wf4JrR7AIxlmJQIcnIX/hUorscw7KlaGjQHk6m0WQQ3TvqrN/IafdoS1pZI7TG
n9Gtp8D/5tRskA0XpgEmsPOHXO1M/YopBxnnmftIrE0LgQi5aiFe0zSKfns1QYtk
itvcJUf8nhksUzGqTAAP3XNUJV9DiHkdA8dGnu0HTASJCJd0714+8xw/u8xSpq9L
xZXP9L9oitfVlWNWfv++/uDsVzL+apxf5yc56ixq3/XAenhcZWdbS/68mJI6nZYP
uiHlel0T4K97V6S2LWfdISlaShqvNOzwy8OrEg9iTZQ16nBlXZiH72OzPEYi811X
AXsgWDnMaQLIXOevmyK+fucnRF6/GC2DOjfhfz5q/e28/QxE/uIrsz26JWPfr+8z
obCu1xiPBJlGbVbUNGwLbJ8Fzaqro4qrC9XYnyI21KhJTGmNH1YYJ9UxHQvZ/9A3
vYqqzcSQnEfZ/FZgX47hluKkar+4UJEo7fphwU+SLN7di1eh2y9lqhVxVmKsWEdw
1Mw4lxAxllxotFp0NgENLcLitXSoJLRVNZus5gIRM5IBYkp7RiEkE72+gJy0xhUz
0kK4GSk1S0rpRMxGqTOVIvWlToxSWwc5aHxVRuNYVU02KWHmCUWE9cUShf/PB0sZ
soRXFopnmWoVgqPIYG2Frs2mOXsfQMaUbZtxHnMmhUwt5Rqt5JPutud19uLEYVjJ
jCtEwEt/1RLJXVO+07gw0e8cRHBsDyjluNTOcXmgMrSUOSe+YLTd0nGI7wmeP2+F
4GjBfHagmJft+eOw9JxE+qRcqzVtglMOyxXxbBMMYFw/eqNn0AsOd6wf+szmSZu0
4+IbTBNaNAM6mdrRWS0PEcuNv921jtVqRsLOW0RqnWcxVGkCOucvKU9s5xzN5M1R
0EWSM4w6Um5d9W44f8BNlM6x6W/fU0p2f6ZOwn+tk95RXiBxAg54j/7jUgD4KLfp
5QIioiTRkJ1Q8AXJs9aIzKpguKbumCT3IdIGsZf4+qhzrpLBae9/Di7GNYaLm/dN
H1+wiP7RInWSuRNdZ1RKLQ6hk4dv+V5ocOy/Y036MP/EwO/PoTqr+v2RtoQCeXfM
bfP1yG2+WFeyMuotPxQV7VsVDb7HDdTPXAb9s2qJTsySTiIEnnUuyUZX/BNsbhom
Ims3O6fdoKEy4z+gp9HCvplW6ecojn05rDC4t4Yvy2UQwoKpI9RRqY/VCzf4CcRb
nwVjraJnSlbbImWYXisZrHE9+/6I+Vu85ypdNKhNQAi3ENWW/vM4nMdZBFTj1ZYk
jpGQkm397svX67o95Dh0zzhwjNZNal7SZgv8qu5XRXuo5oyc6YskCqQF1HvAyaR/
LNnXIpKdWorvrm+tj6QAFpGk/qrYls+m5KPxMkPoLRjjdoZbuS7BtZ+s3OQ2+sX0
+vtIZM+DGPAQMoR6T0GxgszDh+rROPmIlOeQ9FlGN4JZ664LW7Yki9EDoGPyVzB2
U0GTVk5l4jyr3lDDntyH/tyLj+Ypspmh7LzpLJaLnQWH9UrjyYYPSqO1yi4rtVsn
yzXMHStFWVD2mi9nDCfML0R/0UNEuT4UfrE6DgSeC/XN/aX/XvaMChM/JYqaXNhk
zm3uD0bpV6NRB9if9oJspjnX4/nW3OcZ6yfvQfK1J95j9iA9rQw24/+J7CuXzPu4
MBkzjBGzwP93IHWXaQghR82L9lrccbPJxLH0us5x31j3Qd8GygES7hMhTqEaPp2B
ScnBfJo81BCLdZ5PXsE9M8uJZdSXG++A8cDhmhCrw3gpUELeVl50CLh8ub4FBHkL
PIxPgbHDuus/7IxAyEE7O6grZdSfJmz/c1lWEb3WlWYzDuMjt3eg3ENg/bKi2+Ew
egve/ld3o+G0/nrwPgEw3nc4eeX/DT1hrjUId9G0OX5y4ChlcddfWNragdxWDrSP
ZuCTpb85GKQlmC/pkZivA20mwD+b/bNhS42idWKYVCuYq47Ds2JPq7wjyENDteoA
KACIZam6rvZdTXmIwu5l8KGy2ktMspneNqH/nDw8lyhLYnd/x/X+JMk+eqDRQ7AR
/O+EI5FzeFf2/sf7IiftVthbADH7tTZKf/sED2x8P/9i4jcfHP/ANn+y9oXqiTKb
4gVJU7cCo6aWKPHkUsQ9kJvRyW3Kp9olFr1Imq0yGT4d6V3OV3vdIDeQmHjnW5rB
sJTiOA668GWWHJAYo+2989pAwFVy6yIxzspyMdMWYIWE6dnZ0Zc+whhxcp+ucHML
CoZHyha80c4/svLJeazN+rbkCXD1HCJWLTcAUj84dW47Nn8EmB6QueT83bsSfUl+
+qyanbxx9/76STktJe8Txb5DgDRukO9xeFAmsi4az5Sz1h8cf2eWi+Ypsz7hXXu2
WBFA/0SUZvaG6A+xxSg3r6s4s4Yq5UtDQUMOxx20bs8wWsFm5f/LXircDQL1ghj5
12MyQ/BbHS+WcNk/phf5JePUW71C4fR6orz+rZ5WnIfkY7vAtvUa/I6WSDsIQKGT
6TnECozevO0Yh7PGj6AxAAsqw1sZIcQgx3CCGs6tAeeGUmF31DlcR3Ll7Yoa2RF7
CLZkWAOjxhH3Vhr6N8dvFyEpAFvSmOcHv+OcZIrbWqO3cH58soZlj1S8a2RDIN0N
O2G/lRpw6w+WF/QSmW53ADVM7r9ScgGfbGGBMvtzEJVZUN+i6WZkJIJZWa8XkdKY
zlbkOIiZR4H0BZZODrXNf/EpmXQGISI+hV4VwLfLix30cdPHgoH4sR0kCyDBmECo
6uwKj+mNg0F7GPrT9zQ3Pc9xePfDjFDCt7BWpvrsjlcdnWwbBdm3xZxNQTZNxk3T
y65/K013DMDeKekvJzWTmJeJ7I+vbG5gWj6oyniHNEQhh3Sn4osPD2/MCe+Nj4BS
kzMapai4v23oEVRCXwb+xGqrTftiulwTAPcN0Ki9y+aALUfRF2sAlLmdSL2Mym5n
JzHzuxMdOgisfxx6mbwCD2GR9h4vLY4TuWvkVwUWDvkO3z/nuZUAhUGMiOTa/PKW
yw7Fybw2xQB8hXWK5XbyNQ+q1+lzi0mKMv2SzWc8HfRW+fU1Diaj0ezOQVLcT7AM
2zo2HvlWI+qPZbhvTFOJxYkJA6vv3bkoZI3nHk25apvMBW/RuK6EmVv91Ln0sYrC
h3GwHJ5yNIL+GgAqhE0c9c0eEwVr2d17bvtTi2VjpkWXrm5XSrfdiuFUotwe4D4H
w5Ch42fWBnK43Qhxi3S+NIZ+my88/mnQdViwhpRKMDAZ0/src6+6EPA4lncOMcXY
KrnfFCi7hbEL1sssLTWuaEQf7RclGAVQjl5bFOjHCctPzknErN7A8uWVm9kw7bKR
0YYTq4xLaCQqPV5yStTkuIVaqeKQgSsiWyLflPcTwc+H69Qk+ISDcd+EZAKwTKpp
bkNHbVS4UvmJa6fBM72ECK3MtCxaChnfyChP8tuxiUoR1dftH9PDrTyunCD7dLoJ
DMgGkFu8dMBtdKQpNyLSt23nOUxbQPuuzFCKMw4uruI/mezsDAu+D/FF/+szJeqa
vnKTsVIzE59zahVRqd4nd0NfaS3WFsV4C/ufV2J/nZ97expbbX9kqWG0d8UbWvbj
KiauvNnXjpBqddoAmjCZNyNBhzHvtCXsb3+2PEkh31TpspL6fnYlv5KGvf9/SXla
ZHhMAZoa08DGz28UVwIs/DFRBoleD8krKxxMXo8WnjzU6IXic0gkGmU5Onx/8yKI
AAaTyiVulAnGFdt+MknbM79XjjqzJCLaECV5REy3btgUNblQpVkkRca658n9uLZT
j0Z46HkB+CtTPXCtgjE0KMGwJQom+tmFQ+9Qqr7pNniYqAdj/ZQyZ2tvsNOBkf+P
Op9C2p9Ai3dY1wHJq5IyF0T1Yxr3g+6GEF2B+6NBxOSfAQEdKcsBs9Fp+1SU6PZ1
N5u8Tcxrsxb+AZXnO2n6L/jSkYfU49BKk6ynROAtH+jB0oRzy5AyyJB0giNe+wnI
lkonbA5/Zss2na7LSX8SvISMZHcnB02QsMsqwxWhSvPaRzhgzwUD8137aW2c1IpD
Ho9RQ/b88mmCsYHhmo9B7cNOE0OPlID/Bmfp7H494xwSUtztMvSc3V7/WiwFMlVg
tzx6BY4NpNHiOT943qzRUxaaTz0cNLtqSJ7VYvxUsnd7k8rpWUXNuTjwscYc97X9
X+TBeubkiWw4bQ2nVYGFvAAjnBMJIVghIA/N6rhKfn+q7ajTT0TgvVi0VwhUOcO9
/5lQSUx/2bopRyrDFM8hMDM1Qf3xLPRofo70MACx9wmx5Aumf6YitBSOnZnX8wpk
KQXO3HV7JPQ96xs225WC21I6TTnTJ0MBIn7tqeLAyahUoKF4ZnHyWQwgIA0u+iNC
6hhj8hxMcIM30C4Aul639Me6B/+w6WaczXue8ONvMVZVZCtQy+gQ0AYR8SMciEMA
sCqm2Q4skFLziFZc/TLC0OWsN3bsMDsWeJVgyNeGXwLDqYctvAEAYfsYN2v86FY/
RhUIEHbGtDEAqNGf4RXZodm+Ph0wPwn6SRDrlisCsuooW2hmTeyehvHt8g2AhFaU
wyw9wr1lspIDDdL2sEvnIT4RXrYndttZ0+vWOwvFyuO+J/rOtgjFTVW1G91e3qNL
I14ooZBAfdsb7/xhPH1MHntuE+iF4oVGdVQ2qRaylSQfEw5Zdn00hs33ufFJ1N9/
LsalTZNI1/yQ8kHsQ7otO1iIGd8enVckWdb84I7hZapiIWSbvPE6rYqMlUrLiA31
i75PYjnjudKs9KSiz5TjdYZvutaXhrjbp9bSiDkfUbZkIoFUxaXth3YZ/u8rH9kG
SnVBSWQ3wlSIgDj12fbcU4n8l5Ibbmbt/075CrAT7DJ4HKxjUSmc2OUGoD0cPKu8
y6QL7rieU9whFEWHjpxsJUtNNDCK6cUtzozpBJRiP0uKT33FpX19LcXIF6hgo3rg
V+Au2QZljZ5lGj14f0UtEify5kveluKi32668uux1TpEmwaLl2VjgfYYg61kkIYf
yFxxA2dVspfkQsjRpxqK0pxEYKo76rtNpHKePyA+ZN1iQyPQArpOewAC7aJ0wfHt
NMxhiLSev8+V/jfEJeBQWaqBeoz37T9KVKXF6U2cN83SZA9nlVEGAHGEC/nh751n
iSoc8q+zsaj2Hv0xm/gsHnxcjGp0soqW0tYBRb4PA2LbuguEaC9e0tzrpkZuI4lY
F6rDyTQS4wppsJcfbLokSFIee1MB01srOU6Wl8lFkiAP7JisH9AYraeXKkBCosmy
kKSBj7R+tcWWLkYQtqrUw/bwfqoNa7LfHszcIbpKly9N9Yla8g88dfl8bgTqWjOH
GCOMGqfJUYePcK8NhYeLDfvVQqgHQy5pfntuDQ1R/0IOnh42gBJ6W1lOplAg6TOe
//Yfu57k0Wd1uf7kak5qjFajY/nXsko6oDUtQJL0NWF65MDgF17ik0HoOL24nYWz
Pr7bTV9AyT7ztWYiaHYfDtzv75KqV8v9+adJMdOykR94fXxxns/BTPVkHbE2sX1J
v5Dg10W7jMMBuZGtIl/piLH4KuZLuAl3zxZG54kOC0DT3RcI+0RWnYKKINkhnGRg
GQzVcXAneABNuwAWHZKmiNLojpuE8hYwNFAj3+mDPP/LOuDSqZGJFapYQqquP4c1
dbhetjBA3LAkuGt3EFjXQmXt99fegJE6uw3HtnJgbALvQFKPjAfz7SkJ33oYWO7S
mUJSxhKCaeyX0oCh2k/c6Ph6XFXaF/LEbvAL3x86VgleGUjy6HRd2+ffO7yess7w
H9r0xBkEJnn2IufqGBp1AhjL4qez04GopZv/pdL5MKPsYmbVA/xYuFVHiA4DJ8I/
cPSiHd/z3u2hNJKO7QU4yncY7/gZHpuGr7lifepxUl422/SQhPfYLbKWbP5C0tFm
b5cHAj3PrJ531KMNFUJkaI2ylrqBX+6R23xLy5qFWqQjWRMhlR64DomLEdfD61Jc
kV30qK3SEvCUTGUfyiW8k9FGWw36i8p5oBSNVTdKzh+PR4XbIYfyWEPVg2zwF3Aq
/3zdtZxgJu15SR7vNiW/ZoPko+P3QSoMcDkkmICd8uwSAxws89hMVpceYxY5rrUB
x5Lud4jWDtk0aOHfo/6zdeTfAZA7Ffd6AXsDnMLN3uEwKwru+vsc8reI4phmFWD8
tmOfkP70yIUBR0nN02ghjTeWqU/6c86h3M2FVBjn1AfTgzQXaUMTkw29fKkY13D+
bhcVIKmMROBUrcsI0CvRrpjQBcRjITMTQb44xBiYsehz6976ztNzIss6BMPQKy3r
d2dgu0JfDDtvila4X1jsfbImdIMzpTXxia/a68rABlCjW+773l+NsIVq6nAyMcPr
bJIumEgUg2684FhHU6VTSHGFanF2j+8AhN0FWWZghjt01+x/tqOKwVv3wORtfO4F
ZJnPTejSlngHyk5H+pHCsok+dqAwRW76KVd6ML0sP7SE7KqMUzGqLXcX17Hgse5Y
n9YsQSruWX3DVu9ZZKmallZoCpEJ1PYA72sbE1nrNOy4A0n7W5FlnDoLnBgT0fld
/rxhXnIuZ8kKimKGGlqK9PQQWfidWTGhI0yNoAnyFB8dSPQU/PSvFpHu6tjS1/TC
iFDEbtpV4xRNmNl3fa+5hIOGyer2iJ7+Pq/TVcBiZdqi7Q+ldJKOYY2CFw+u0XJG
6a6hS2hu+iyTOI/zyYH7LgAAyfgizDadjFyURkdsvbyBRnkv8xKozmBfEM4b6cOu
r50q2b7mmeSEpSQFw8wMxlFcHwWGZrFFAbmiD80DJp8eqJO2ThsXITnqiXwK2vLt
H7nL0JnKGS8IB8r5a1Xip963Anp1B63rPAj9468QsG0KOJDK94mO3Ow3L4GYsHBu
aA9y0+c9zAcBmePm9eaVXQ03CkhQ0Hq8ctuWUqvVCQl8X6fU9lsE85RUrd88a3ZP
p4cI1fShOGAD3geqBKsPdiRx/OsegjfXb+5iOr666Uzcz2r24MwkxkQZ4VdIyz3i
Y1LmWlXISZOyC+8EmCUhsn4CMDjQRzyXUctn4Y4eDRI6hKLbe4eTPxMrWwzppDVX
SQ4vArN49b6PnwPaCMzq6Z92RXkMGmiIkf8XIrE5D7AmjHP3ODTU8Pp2jiOyud7U
L1FZpM9TGBA6JscEENSYl6ZE9KSZiTKob2ty0qwTOP1v9/qfScDNdGRUzaaRdynh
xIL2972b0SAbpPtyUyjPUDuaIvLdogXnvKTou+R+d3hw7bugEfsGMoYhL4L+IJKj
OltzQ3MNoUKozhRS8Lp4iSB8ZFLxjjtbj2MbTMi89s71rTdiKn5k4QP8bzHZEKfs
AeHQcjWKkSdDGtfuUWtjWcL2hTF/KqE5vz25wHUXF/VauF1kx8ymw0lNVBYly+kj
7QdnZFmGTixPjxzl9A2jSb/v3Xz0Z4XKVWBFnTmKyRKbF++6h5BEFfZm9pHxp4pg
7SJ+a7cGN2Hgbt3DA7/TJnLTvhon0XdBkFAsEYqDsVarXCJLTYMzGsS3nLoQro+C
F5cObyAWNNCYlaocU5k1izsW/75plviOBfNw9QFN6yrMrbL68wvMYEd8NWtndM9c
HKdYzr5Yc7Qpt9kzzhp8u4Urpzj+RM0+i29uwUB8KsnOoRBPRUr2MtKcpT9mkYUh
9DBPu8NGVpq7ixheAlj9Z4Skr4YxS6s3/w9yQ+v8SPOiPzFjbLRTlI9OMgOPDHkU
cnQoAtoIF2iVeAUcOwtl7+Z6+A9G+PWsou+equikPuHbzJDAz2AZxvrT94yBYk4p
/WDde1TdeXLqgSax2wcmWEG9DfFzr3Ylzu+xsARn4bMu82owtnAJCaXKtTcbtn4D
okjiWfQ7IOkWhGgJsdtGaVT4KxU+wjTdyTjEwxnYyTF9M5Ab5Qg3EPYFuQ4twB7r
Id3nd4lrEWqh4beAa0Wj8BtXgRFPGKTMUxkzrz2BXzIWWjJCk8h8hMRg3smiwZL0
XGE1TLhwCn3zwjeDlVTdiJ1Q/CR+mf2564pmJFvz/9wPxxXh7yiSLRRc1FLVOh1K
xVd+RqieGriXy4NmGLZ3ubSoYAd1Vg8C92l6sWcP6cfIq7Vx668nQAS4sP4NXCQw
4bL2US4YAJSpsjwUmiB7jrGlbUypmX6n7z5t5qfSQ5ZalHgUCXghNj4L0u7D6UTX
A6419mmocdnrsvBGScs3qPzIdyMoN1Gy3vSFyJ3/9pBkyr0FYlBDl6mfYO1Xk15C
M+ltkmI6fPladR8RcB1pRhdD8/77qtY+MGQWsuj57W8D8aTqxDNByC8yO9nE2A9E
Y7ZUo1dKeVrZLmF6mJ4AaKaq+SsVLb0VCfgx7DMjyXWmZ14kJ+IB7R6qY3mbOVcS
gmYaKKjA1OHTi6s3BUoc/2F7F99yZAdAyFk9UxR0iR2nI9xi+/rHh8amSm9qxckJ
ctQL0yDzcOV6Gm19yqItpBqX3jBIMrOMBKNxVUVKdtScIxuMHzE5KPR7bXpH2Pi5
dgior9VuioJoM0cy6xa219kJ3vePy0QDiwTmn3Pv6GMjJFJtwatlGCJOEMYysgYu
F7LgbkfTSnzm5qsQUxqZDkAwgnoBOAy41XFfGdbXEyZhH2GCOKzR2SL28eQkgBVi
sQPJ9txE1vA/PK+qkBG7eTl7Q5VNBQH1z9fEblnER0yMpwqgzmaqajn2WpiMl/H1
P4k6uuNvLjZH1O6mVJOcxF/aOkyMuOrTJVk9nH4gNFgJhnGACvGJUDyueu7OZzXb
33w0lE4uho0Lh3sFaQZ3PTfH/7ZIQyW/E5tZbFKruWfHbwgHrqkj2BykfX5dhrMd
JUkgxFmkHPvnQLQJP8GRa4YmfX3MicwBli/MOXjtqYubBpALF6jaIISro1BY86Ic
0OkP0r6f0k7zPf7PobeAZ7xNgj4I2/Erk7IUskCQUpeux+dfHGTIJ6yN+8y2PtVl
ceWNKR1/imXrhvPcVXHJK6PsIlBcQk8XyLGtCQsdFt6ckta/2nGYLwsmbZY9vrtZ
ooGF0ixRcArzXW2VdtWc9ErcQrWaB3IQ242ouNaqSw000TtFfs22wN+i5En7xRmE
kjpDbbhBugqkhNMRiOPLmn/bcLGnENLLbXnmLgJgTfl0NnJVTDyIxo8wb59LgSO8
ZQ6Vqyu3T9R2LXo33j05lfxHKLyM2bOuUj64Pd0eXftxyfDPojL5/pTCMmSnvOPR
xklo3I2aU6LNGRSCI9u8dfS/wnoboGJNyQdq4egTb4nVob6th7BCZigyTGK28X7S
XDkRMmFUui2vdbhBRsHNzFBkyH7CRCz5Xjq0UWLTGAejCDJooO5D4N5UV3quwU7V
gSep7mfoTFodkRDsJlS5wfZP1JOj1G2cR3kcmfRpUFUIb3k5qYJgWgOLTpoNnLJP
w8NkTFgz9mlDbBXWZw1htamybU0LVM2WvoQrCu5b1XKuFbpB1T/zv2qzaHT4/3B3
vYGtsMcigByoRVYnqbH4G+hC3u/oa4vSi8fnRRG6bEqoxP/6xsTTVbp4Wi6zGFPj
Qat9LobOZp5JhJWprSOZr+R/Lunp8ZtTbm+UT+zfXO0W4RRbGmaZ3jSnTp/M8ljh
rFnMkv/XZ2b2/f69et4mR2RGeHJO1nY1IZJHjt7kyLmcx7CKSd4EXLy7l1LYgL2e
2yOhSwjp5l7k1/3HzWHfQvhO/gT6Jy7icOlpBfeI7t5vkdA9PwQtJgfEWOHDF48M
hUK5ALl7fa0KzvR+UuolJj0aSQCJhtJQFiSd3/gogani+gv87VsjZXglg5aDC2jb
CEDwP98eZTaUmuJ5alKB5ZO4MSMw97EV93/tqbVKXC5ZuInCYE2rbmqRywuNtl8s
TpnIPtOuJw3x7ngNSECkfIgQk/RProalit4nMYlAS1TQ58I2RdqOdmlMD+6wBJmW
cMoQeGw1uEpmXPhZ7ankO51xrKnYTdeosndpwLZ/9kV3ZTALapmg3E+LGeNWywNQ
7cGDbW14KEMaYQpQxVbOixL9L89rtWn+YOf7J+mddKv7nrG7pOgWqKjVlKuSfgoQ
hw5hjIQfDk0gzMjl1ZsfeetaPzhfKPA+2HyInkZWdeZHQIn716p5gF6eepRpIUlq
Suocz/hZ0L89ipScM2a1Swu7Zrnl9FKGdsf8m233pqCc7C0+OexhzW9DR0g/J4yC
5T5kPfsrM+CoZsxFqLulzACg3YeL2vtxLKGLy9c5xGB8Ew1AWFA8X996yeLA/Azx
mJlNacI7J9RUB26Z2zLG0/5cRs2JtHQUW0LKHMnH3EW7hlP4+UAdN2amUJIP/7NV
nKsyFDMqbCM6vcL4Bljp6wc6FXtMfLH/k+6korHRzH5zfWG2dgHHmnZl6XUjdFJF
57C6g05o63/1Tji+10zDTmILERmf2Ey4dfBlhJsHkVvL8k7KgBTKNjivPCukzwuZ
QDMvg0xEYqF+2XxlxExrjm0CLRb571p/NUPbEoT5izEhW0XLptijsqJ3ZR4moOB9
JhggNMkfVHwg5QB4AfQTihoOluX6+5GQ0XamYcnytm5Rd4gl7MDQHQKuPeMC8w0M
ZNb8P4w6EvPkrXXdFhsq6Pw6EG5LoyhgajV+qQ5xjYvkKjdFOCZ1ubLboylmiTqI
CC8FQpekq5elcF2xw3D/aSoJ0YFsBprcMdZF9J736/ILg9nbTVVII+MqpaztoHOl
UtTh6x3qqS0GcmfqeVT1VrrFmM77z3ThuVgt8SnjbQ14tIwr0R/tEajOAWF/1Xk4
QZS7/999Xz4nvtwEKkkJl8LP9+aGIP+CoE/ig0BzGnLwBcQCzqFosVPhFRtHzM74
EYSBqoBHvmjvR3P7BhyzlTvpJBzO5UQHO/TSMUiyyRObn/WZwcczK5RdQVZDLu/c
cmmqr2bXfXmcko+B/Wh+F6lUWsOXltOZZEC7KTStU56cTezvqBKqh0uIvNGbn3PU
rD2QfPJpIHpo9B5kicD+OjeyOSsVi/7CKeMTXBQz1/wSsoHvyOOx4PzUBVZpULBv
si7Re+D9kCQcl7pqDcW7K2obsW6lTe3UDKuOQZ4ziK4GmpyqP4GME0EuSvUzwChc
vfevIIAf+vwJEX+XutnqJDiFoVChJmE7CGGpF2EDafx4KLO89oE8Mo7iNVJKxGCf
AUpZUdiF394DWEs6c3s3pEWmc0liX/3E2jAvRNdyI4OIGeT/QpKpZhALI94AmcuB
4DmT2Id69pZAte0ObJMKInwmagzrflkxWjHRaswV5Z+YirG87huZZOrYqPpfikX1
NFpPYdlQBuSRja2km0qsXapgHN9UGgko29mzn6n3uJDufp/VykHwuS9mNoc+oE/I
VzbPczKawNd3ep033KO+FRiH3PJOAuNmxYqpX8urQMIu2P4SofAIp4R4aSH24Krx
+5BKW/sK+p8sMZdb+Z0AAAwwyb3SjEeZMjbO4Ur8ikPnDCk0oKBWvaBYtISZ+htH
f96gHp3WSmkFKsRXpDV0heuNEKWmg58WsIaWjF6LjrfMgHfntcPYFWhNkdzfZfm2
OOzQEGGcgnAJE/OTqQzAtfr8TL2lE9g8tNlCvCGH7zwTzRKXzWKX3iJWCEyw0ezg
t+lytgkx8Okkq52ucPiAhzhVXL7ZU6NAn0WY9EuIwri47VxVDJdKIy8TgWcJtLgi
iKhZ/2c8eOaoilEsYA4E3PqmbXz+TYZ/ldfqSy3Cd0/0uqGGcXy7sGgU75/n5JY6
xkULmAAn1typ8MdM5PNC4mnifiQWnv4yBkcfpbG9cYbe+1ASWoyyuX/wanAMe+kF
2htTG4+jvZanEQ/RTx6zYj2u+BawuB8KJM+ltmB74hPOuEHmCeKjDlICNRe04enD
2/UCr+VR5sPW4yV7jmurOkxYd4MRWqNsRZt28xu2ybCtYpXdFiNar4gFOhqEj1KE
SGmsbsWiD5Yw/tC+nzoX0VjxAw2m9lXGP+/2LyxW96Ukn6Yyp+GDN+Uhm1DTq2Bw
W2bVAnrA+W7E2y6s4Ptr8BAK4pKAZ02lguCtdJZ9yuVe/BRQgloZ96mkcQBCFkpU
x4XDnD7jxGw8xaIVlbvViWLpq377XqJ8QO8IuysstwZmQ+hqUnTmqMgHzxxpr2uK
/4DuYxxgiQyk/uLeE74r3DD0SsBxmg/3oMUaaCgZMG1f1mz8YAYh8p+BufbDnvUa
ZGWpFRU+HsNgpynrDUAGZU69zvh/qpmVA/FtF+dgM5ak3jSqC5b8AWRw4CJCqveo
F0zrbHbOBRZ4N+LlN6j0AJR1Jnx/SQ4PwcfZxVZ57Fsg4I/jkMTHQTDxvSI/NFFe
N6WmtjYoJYR5KuAALhVZMmZ28S/Udw5oAYELYGbWvC0yJH3inV53bVHPBJKPXyjP
gsY/S03TRU7g/JOJtXuOhZGjbfuzZKj5Ybx91KFTK/F/LST8rRJBO7e2+4w+8keW
ZyPtZ/xeUswvSSi4/WnetppmRLEoPFHUeMwkmN8GJSW9zkV6vVq53PzGBmv0Hu2f
P57xRUk9jEPxQTIL4uqn3n4okJT9rXsGO2OPLg1tLInyX6C/IvGjrdmuFekNb8aB
Gk0X4hSXA8psFr6L2LLVowNKlQ+6r+svRv6mS8DSIxvBQne5I+0mDlPMssbYCRUm
keZ4FdK3cIFfgxvRsGDCleHOYerE5O4n9YGo1Pkop6VzYwBIurZXAFyyryDKkfpR
irlHyDOZE5/MDCEl+0D9hd2SWvh7OJkLrEiIsKOyEHUcxy6D7qpBidJp+YbQcBrG
/I4uBge9tz6ripKiurWKTk0p/yhvR/ushytx69TQDgZr4jQtrYcGmQkNAEY8KQx6
qYBF2RAE5i8F8zTFrvd7RazHDVH765YHhFVBgSqpskegNqIbJmlGOHtwrNag3kIx
k4h+n8dtTBnwCn34KEG4gqyd6rQ3fcdocvHVZIBrYeMNrPyN4Db3syNmeslQ2Rnf
Qo9ULCKeMy1lkdY5AIctW1uw52Vbfz1HL6EThwkRW5vrnasvApsg2C4nOaUrgQZs
ZoRDC1SDqjBvxVM/ZFdVwSxKG8PFAY06PhmY625fUHrFZghSqxwPEzYN/4Xp5k7f
OZl2LbI7u+cf1hlqCExwkNx1vMXij7V8i7JXV1KNwHJ5psQwJUBbpyAeL+B5tVyt
pQjYSiJtUVg+dX8O47K0DUt9Q1EileymDw4Eoqeal50KYrIGfF/vh08PM19Dm235
chQ0aHCnyoUxYH8yGie+ahFGIZZ3en78fIXjmEAQYzy8ibG+0EyHLFub1XGDE9z+
70RgOcVmXvXKeWEP8ig27aOmG/Oeb00yIwWmowGwzR8d4MhkYsSRVug4XnxFqu7K
PYa8781atgQ+2ONTT+xWnzEHPjReXW49AkdN5/F8EkQp1nQuwDKfESUsOaZworbV
2dioEIpBVeD+l01ZvGEmBLEi1ssJvNEaxMG6fbX8Bj8RizE060CxHvb2fK20pZn2
boDhtN+xCjbh7WKNrl0zA3QS0ByPU7O1PtRPARmcogjAv7vTpM/w0nTEDHh5F4Qk
7bX8ZHLvTavCOyspYKjlux7H/UZcUHWU0CNArDRysSbXanp0Lmcv/RYV/FFl3zq4
YBo8Cur+8WsUcxqLJA6lsEobhjjBPij2+SFOho1wH0rnh1ZNiRyufn7pinrnGSxh
JWNeCKz5W5d3dSokK8Jon85yMr8ulSElbCBXzCSW/5WYbc83kKpZgcCjlxIUFO9c
nm+3pS+TjYy2aQhD40aysD5Faqad+UDXoFgW/KzBeI53LSJCqiRPcNRG5tsUwDON
7DTyqKCPExEwTO3+Vl37xHouQ5K1ymCQSydt8jheZ/lFlf0QcwWUgQnj94JmN9KJ
LRokJEjHUSTiLhLWBYcXJQefOMXxZHzjPtU12TK80ISV6pesjEJObO36IknmkvaM
EOvmGThY7WaIk/9n8TcHfJot5sEV637uZhPXgcHTdXoRehLsgYvegFPKgvXC2AfJ
dCYQHJMDntRBoi2wHL3DVzr9yzV4IDw4CvS8MOYSc8kj+myBMmqdWtrdZuFPW7Zb
nUUCcQU9wbSW+z1CJkzhVW7kioLu2xWWconTfBEhRd4hiVACQQ8FFL5U8NQ3CYJO
`protect END_PROTECTED
