`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TF4yUC1nXsBt1McV/w5jfc5CGPo+P+CM1ntgpLGqTQS/km2ZAYRde3RA4c/2/4LO
gt7iJee1+yPQhsnO7jvDMETOtJIojyS9tossPCzzHW8jv6gZp3SBxffh3PV1fht0
LRz3MR17P2mMz+t+aEK5UdW7brxxpWTIuc76KQ6zw1OQHG1cN4M+gTzWTG5+T6Eu
bTlPF9JyVe7BXLD2l7Kno/Qj6Ye0F/+37eIwTCnufpbtcmhQDiYoLXXz9avfW9T/
TdedQq3hYMmDJ62M1WMCY9nxxdQhdZzEQtWqDnk4TiwybcqQv2UiLWhGvrauZLH+
czOH3UnW13CKL3oCsSKkDVMymFIyw2jry3UObsvSXuN0aJZUcIrIu3dAZBusgqA9
m0A498EQQAfJlFhyYiRddjVIAqh8lob7v2rGcdo9Fkyxbc6REHaeN7ZSytxjumSS
yoDRhti6HHCaD+2ojJhli7yLOJuUt2T7RzieTAMIDi+INlhU81+2GM/U/BDzllSh
VK79xaOPQ67w0YMnHl0/wEJQczEQvyj/NssmRmzd51TPRJr+rmQ1uJUxIaWwh9Nb
hSlWUpr3MTa31GCHz1FBKvPjvZ7afpahrSn18VlmunWp9n1bVg80KhsK/U7p0jdd
YYXItADZVci2NNY+RV2jkA4EjeoFNFm1lqYeV6YO5vpIyKmr5NKRoM5ZYekW4Lga
ypoaAAnPryDuWFglvfQSLSAqYkjacKM+PJnJnIJwMW0GQbjZ/wv65X8g+5AQfOae
avmga2WtoHkq/Z/enJK5XCeh6kLcBO2/jA98vZm9/lwLTnFkK2cWoPj+WsF4IrvK
nJE3shFzz5yBrr4xOo15cL+qhe4i8jXQYfJi5zcO8UgIEqnI42Dbj4UJsaqMDhF6
CXF/Va8Khdm5uVWYqIDhNt1tzxE9tblut+RpjKBTJQAL6RFxclUj8qMU3gtG8C/+
n+5lJrEdOZqdpj1sxjj5P17JqZFjiLoORmOTqAQI4uUat2At1JgSCfPZTlQkyODH
mOieYOb9dJEpwfMyK8oHo4FeFi1ZAHji75dz9lOOWYIxw/6uAuV/2lC677MMLKqK
5mLksVvO40Wl2Jdu3x+Lpcod/8QNVG1OJSOKHoBujI42TvGF1HeI9i+FGLUZbElq
jkzZCHRtxL1xc1rnv3nJY5Zgz/5WqRJQwrJfGF6Ags3UHyMikEM8PHRmV30CGGAc
GD+44f/tOSTqrY8UFfFjX/UyDhbvYuoAdLGgSK32INRNslfNVPTn77RnwgpxnCyF
IpDylOP+7NEbcnOSRcLfzPgvu0Itz+N/6g/ujZKJ3Y9feJACoUB92/c9cnYKN3r0
p81pjn5tkjtUsHIVYoQsSMhcHHKGCBD+kQ36nv3dEhUNZjczMVPtt+/gFKROTZKR
e/2ZMM8l+H4L1oKLA7B/BsRuo6LQjhOOMnDVv6JRgW/JJUgOkAWmIYolEQZchQ9A
bWHdESl/n+XgqNp4BnhxZW/StNaBEA32OE2I9BqKlxtr1pzHXJMeUTsxHsTFqGFz
UOOuT+NGPNgLzOE55IxMR61IyaEikpHHlqMmDk6FJPuk+i5TyX0CVC/xgdQQcLmv
70aq4gte5Yb6RrC10UBhW3ypjVkhGeuYqi8P9hmqjVC3Qbrf5Bl/Z/IhmD3kKNgR
9UUtSW98QNmyoRonaEh0kvrBVeCRRhoBCrp7g3SH4HOalK8cNNpIVtoCYc1xhyJe
IaHTyb2XqKMJY4gEjCsdMp1+kOWY/9vJXO/O6x7oHghcM7bW1V2esNT1OgrbHb5H
CRyMUxdtLG/jMH5OEZ2QuB4eA6aWWNkn6m0EQ147vpX8qMzoBUn7ruNuNHDNWRHs
gQChokpbtje2uiVfUelJHfDcdLYHwkuBODnWrlZFMUo8dtp4sL8LKSbfti2BYq5k
bvcq/Rj81nKGJzXM+Za0wWrJrk4ZUueuR/9lAguAOwOLzDslqtvclCWx0tjMGvT6
oSmLuRmfZ6vZTwRrP8qndCCOzAcyf2OH7ZZ1ImRABfwTdN494pMwazpI7oOOHldG
XJZWsxk4OQriTRf8kktWjxUYIRISQ0+dj/IKtcX/QYoJNTjQ6P8lj26QO1rqzwio
4n6sJI84o3+jaHh4TdAKldw7WrdAblzaV48BPF4OTqgRtLXFZSxi5BRXMdtXIged
OkjOryhBVn6m5sEPkdMCJiffdn68JXiBPcps9/xlmvceEezW1VQ9VjGfxeGGdHyz
9lK/idd3lYyf1j+EOTe8bGRrrlURx+d2O6GoqtMn8Ct236ZY/e56VMykdikptdPU
jKmYZXh4E3OwHpFnRArfIDfMHrOaYfMCAGAU9DzBDEY3tWxdRpXH8UYNEEnzVZa0
nhynDhELO8YYdyIAQEFLgoja0t4A68KJmZyUPEa2JTc5TZUcMcG2RTcWtiLvvsUd
sCBVSdIgpUa4/TWMafgV5/U4mi6rTmXpZg0xC/rryK2BnLs5zGzG9NBhMRy0FXY7
C1+M21gxfce/dXTM1jwPzBiDcsdV+cXK+OUDsJ5w1XG0YGwqx4ew7DI6rjAsIS3c
7tD2NamK2ewQdHsRrw2zcQ3Kv7/j7Gc/ox9Qvvgsm4fNsIds6+RvEzZpNs1TEZU2
fJhgmTLiy1qMxRkrAjQIYBn14UxcWr6z+8nh2iQQ625+wb6xgnwuuuIp8AZFQ6CB
9LKY/rqlUr9QqJ3HyYOt1/dC1o0OkhGLKKPEXZxQMsY2aXIlmBN/bIArTDa/qZby
yH6E5s6iKdSlaIN0hA+/r3+ZTbkZw7Y/LCgeZF6jpfJG7CuWVhzDao5YK/lBpF1i
nmMG/JLBdcYFyG3BQSx37RVqjKU66iaWyrdT4Dv3ykUA8kh26ABfT7WraUEh6sd0
OmSIdL8p5cKQ8tUlTO6t2aexS5dXmct2vhwDD71rauVMTs13Op9EYllXyZ6banDr
W5Wq6gTF5/kMor9E480fRChZrzzFDfToSHFzQTWJO8oqnHsvlSKsT0ytREgkb9qT
ytK9QbCsAdU6lEfqj5gGQGeRDrbNNzcdmenRNf2h+YtBgW4SCeG6ZcHDQrTuMsvF
KmC2prw+ZaxTgZNzvG+dRI0in3xsTVzEFZS/GAJtuNPcnyMzP4/ZiEfJhaRi5YL5
VCpyX1FzkkQmCaxMznT55UJPupVLeWy+dE0fPESTs/9e7QPgTr98k7TVslrq+IAV
vAzBnheZFnTVhB8/OrPpzHkXfYAEIqYSusXTNcTWtTy9KKDdSmptIsV/rOstlCvy
wAswD1MPU0yhgRhiYmH3K6yIbUNzOss7+iYlchCnWzejz7/Zyk2fQcF+cczjxDH+
Fxvj3ckGbJsuMnrT24q+t/Bcwo360kcxLdo2C0Nua4kVizozKnIcwGdSj9wlKOkf
pwqV9v5aARFSoAIo+lLoJlshIjeVH6cLUsFUk0L/ab7QO+syCdpXsdZu8UAl5a7S
/UVTw1c99kIVqZkEe70vJ0AujlYaMaynJtKkNRp96r4tFi6uxjqxe0uXvXm5Quew
WeaZBxZwztC8PIVCADqI1e5RYkh22TR4/aGzNFwE68g1rHucYlOCgvlNp2+xkOuQ
/FfT/6AEJ2WGfMCs/wtPgaqaRcFBEr07PwzA87NjPlmt7vQ05tM8QC+HH4A4DG61
7cCBXEQQOqyGDrAHtUfwKLD8Perq0HeObPvAqKiSMIkv9veOh7FtuWoexYR39SY5
eRm/Ru7UfzVAOO0shks7e4mOesrm9PzHe2eNBESaeQddn3NvEZBgM4yZDaLUt1fL
XOdHzav7EEJw8jl/R7PWVSVhyU9HLhOgwjjqVbJJwoaLmi5bkJE9p7C3iipxKZeo
Q1IIJQ/q7/rlVquiEz15X/byefJHtDsQc9Thvt/7yvLF1gcdrSjakGDEl+2xttNh
9gHQKP9DEo65Oq3S/OWEaaAMCMXnDQ39HdEkIdZWLa0=
`protect END_PROTECTED
