`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tOuCtTezG0BQn3ef4rexdTnUZP5bkjG6PW3uTFrHAsjTjxPjsEtqURxfHWrQt5a5
tk019JpDCcbhNjsCE8MdN7S3Yz9dBnZzTBh/ig1ix9eHF3O8abA0QMRVLPW5sEhj
5NWTGcb8xNhoE7c2maFRAaUXNJdvbFrARwiSxWA+pucx64pMkubBJQoFc42chCHf
46fEQ6in8Ixw/NBxsT+PWcORn+0S+v9pxC7TLs6+E2i2YA/tRKe04869Zloqsak6
iByuF35N9yGpi52DWUJ9N8W6bTgjF8aR5e1a6f3KRZuZ/SZjtN1A32BqH7IdVCRi
oQ559kd4c4S9eyh1z+tP1xzlgTLKOgF5QMkZgtl4Lh8VJByyxVuJqGanhJRHxyF/
eSMkLb2sHFEOIF8HvbNT8mW2TfZqS4fp3cYgUieERqO7L9l1uFa5Ni+VVEEnXsGS
daFTedykNDHu9yr6Ssa0kA6km/RdiEW4MYk/Lxvb63VTg2+AC5VnB9v4CYoyU8fa
1fdAqivbH8CfRZPJrKeFuBrvowRhLoHfn11gMQNhq95zQwEs3n72NbMgCE02WFJj
g32nJ6HrRpW93JA/Kw5UQ0zHiDQsrtrE+RogWNFluf+2jPPHFuxh60yo+4YkUcLS
fK339hQiMiCVsbln+3dEuc2THcZXtuYM3gjIPueKxshGf1ILEufHrklcjz0UfNOI
CpZfgsBOpXoO5jPKMwy+2OVOcEShq/36TN3it6EuppoJrwQzQZ5BIwJXrbkJqKrl
xYqLOw4Fdp2zmshayVXlw7Pi/nrQv+45OTDD7Hlw9P4V6tKWlYdcnX2LVYCEhWEU
sjWa4j2ACDMiXzQQVh+tz+opv/2KXQSHglXk7YKDQ828zVXTwi0rjvUbYXrpYkrm
8PcoQFkBRgI5OsKKoqQZ93CG1dw2nK4331FtMTz1Qbdw590cwWZFGD90tK5YKaBr
9otO/pXAtCK4AgxnCnLVBOJjTaejYVX2WHLTr2KiXkM1YgR/iXJbbm5N0tVZsmrs
IeOOWK73DNXSCxThing9BIvU8k90XK/EiqdWFO3RMJ+ATDGg25lHtKxNPLd0ta1K
`protect END_PROTECTED
