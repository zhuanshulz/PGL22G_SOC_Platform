`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5zba+HlgejldH5VPq1FtFfQcd6N/l4UPOUgo26DjWl+EG7bZZ6Csx5MdGKVBlBkz
ouvf86NIVf5SqDp3XfhNJ81ZJcXsUMB2ZE3wFKBeVXZZ7Bd45Fc2ckS18GXpBQPM
DawdazkRucM91kr6aoJ6zqAXAJ41yZCin87oSjOw0Za9ZlHJ4RHOZt73NmiRgJie
JICEHhHxnL+A7omHX7ELsH6R71ZfhjkwQCkQ4CIueTkzw2MuNofpR/nJYIktbmhQ
lI59QK7O/S4Qap2OWt8ocITlMwImAN2zwJX5197E7UNWTCwZu0Sf8VZ6CJ9mxQV3
JxMQYCKCwIviRvbrRD414IRuQD4cPjMxJthg5sxiHX/zoA+YGehV2vhqyUight0+
xXU2xQhwKL4sB+3kPxCt4jzC+RdOPu8uv1dyNCGIMAKWKHKGO+blI4yQeuliMMap
x4gmjsAzVuuBHf8V5M18E1VzXWiiOcF4/GpThU8jE9LyPp23j8SVHaHmRmzDDp5k
LSi/tzI4FQmrU9Fr6FuANX+Ep9XSLBE99fOUQUgMT8Jxsf72rkfKxZTkAR5ddeIl
KWOJH9vN01VHR263qCXzAfI7GnYet4IU07mkpe71AyLNtTJWNn2ER56LT5t5U0Dv
UeuvS1l2shRtXQpc0fyWVc+oiwCYXcugCyde45LyBk3WSyhTGNAzvexbPx37OewA
9OjXiuBT+b/VrF9PVS2Es6mM7ESgPHt1lyj7uOCOoIlA++b9GnfNvH5dqjpaxYvH
veCq8peZsHkMqGuOvNMxmeP2pQQ1ti5sH3UhmLEnkJjeekVecl27NyFPU12vd5E9
YGSNoWpjsq4AP9MEj6V6x7r7qBLUWKP33WLj09TODlV2vsR3hrz4deMrbID64Lua
k+VZhcgBAm8Z2TYxb1B519qFQT7kHWpUPAiGLoJ+h1M1YSl+O0+6XtX/ahOuZJdu
pW6lJ02eBdoTzfEKsYcd86RlynGGS3VT/xQ3EYLCh7o0cv45oVU06wYHnjHc6swX
dtX2Bey6LWNfM/A4QUZdhrucnGq2xSzK8rchVVVIW3SISgmjmLx4oxq7FgmY6TUI
RVVRumEC10kUaKEH0dt7efkH8pLGPpXGaIiQaVz0IM5GSsXj8eCa10K+NFCDXk06
32p9qCDeQN91RM7APe6FqHkCg3pQITTFGyPWAKX4rzfU97DJFANYTBz+Ledc6t6q
sGTGc4TjhumwOkr0N3XPzuk7rxOMJVXlerAFTCFx+hBdLwCYUsCGEvUHmuj257Hn
xOq5b+bKngm8Q4Rl11j9GMwof7J9jiR9M8JncUUC0yFt/M2qdB1G6/t9LxDgZNPv
hcFc2zpi3hkxmcV7LzcKTfMHWDFCYhPkpSFN4ZHTbSvU1KeMDxulcKPYV1ffsCKO
AUw28g/5T5wqz6HAAFFFM0VUbmVh5GtvadLUDu8rDN4Hc/2njMkwMDbDUDq2laNX
FF0S+fTfRQCHmN54+0G6QSNBTs/164en9biVJxFmmNv0zygvpnJfUT3NnA+qAxGE
zX2MwsKsur3xMKurdVRPHBbU9n2YZ2Ni2Tleke3jRXgmvgRbnoO0XzOXDxVnq75s
+OXj3GOWbP/eu727M9wIQFOuj+mVRzOi06+7t9GbYaRX+jL8/MNp3htLZp44jRoa
Q43jsmFlSN6mLaA2O/fyPA==
`protect END_PROTECTED
