`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9dVp7dJ25YMKTayRsEop+mzqu8jCKZdrAqyrirkTeHjgzDkBo8O6zt2UFPs4rVf5
ioe4hoMNMMAvmE7OLhZka8P+ZyfNLyCwXAM3UhowrqKiAk+WLOM7KAVMr8Y8qZEn
6eU0D9ULlVCu6ghcC+I/35taX4mxFeDyPF2rlo1f0n1EBv5/zCVuJygvCR5HlZ4B
QONjiwYNd0Oi/AfPqmDY5JkJHR5cxlkgETLD/ZNx0Mkuew75hoN7P3+8Jdis2hql
FLR/5hTxWJ9Bp3Q0UAxzA2zzQpKqtPKUalWXfstph5Y9N+KrsRFM7MI67Qufsv68
bOT2EkRV3q7nlWS091eSEzXDvJVD+6pmPRZmuy4c1A8/bKqHjKl9m0P7SOhjRted
2zVBNSt1fxAg9pN6kVWGpX7AVy9zoPqkhdi/xgzSfrdkJ67uJsxXMgCepvjZF8rQ
vkKupwvGxtg08KyNlM6ya14HjmWiDHEdcQ44+dpKZpf/K8Celj5C31cDzKuqcfJf
3Fimoro3eLXLH6/l3NjUYRRBYaYWob0qo638EE7MrE2YkujzUpDhADMALl/Sdwbx
omYMOj9C3vN+EGd/w+kL0KD/0MCw5uyHog/ikHJE/8PEHDlyXb1yDXfKrUE8Noga
ATwLJJyocGvWZrYY6sL+a/2F2Wpdxy0EmzEbT46qmcnH/p2jWaeY/J8G27dseyge
F77ZpFoBaNblKtUQZPWnQimWxI5Pi//arzcd5ONoCDsPRtJ+T2kDOT0FX27dqnXd
9kwZaKkoOP4zHdlG5zXXg8ZkjUNpBsZju9i8EPbOBP6thkWzFDAC5IdShe4gB3+c
frQ0RLH/vqkewhGVLEhUj3K881q1nQTPd2h+/7bivO1OC4X6cYMhiqG5WKuhwYXC
799Tegap6/i2PtM/QhpDgY9Ts3kHpJ2mYYSzwhz2CvTIB/Wx0dyE0F176SqDWidE
djtCZxkPYvoV2KUdiSA+bczxhQe9L3gJ57s3R8RpLgCHNOQChb/Do7H5iW3JzoVJ
57tPCGguQJdOvudWadcWflRy1UkyHJB/G3wzjh+zBEEFSeWxwSgamSFQOLXbXQAA
s/YWcyy4EM4HwclJlxtXUbs6t9el7YnSa2Z72G0edpn0Sgh0vMRY4o7OqSXZeGvW
ZOP8UzoI6XS/E4rjmw/1PiuVxGGglvjlbJMAbbs48zzZCetWhogeZ42HmikdZFvF
O/eGKh6gTiZh3PcnamygiDkNBuKybmKwq8SzkUtDa1dnnoIe0Jm7LJKua65jXQ4D
np5wxFeY8ZzToRf8qKHJw7uHd7aPX4NlSSjoFImj6NmWarLTJdotB6/Tvprp//fz
1Nm1a71KbmYnXDVZSig7SAmiyChEZG4HHjqRnM91cVRXtjTAWxGt7PF9GoqwKpZO
/OASAUppdC3DDrr6S7IiDb7gv8YlCeHYhZHn+FBoZFnKcSCWmvsD4u8To7qiGDbE
gQd1yiUhW0oOzqLYCzGHqFZSsHDKB2ptg7zD77AToYhPWv6uR4/iRBVENoZSd+YX
/skJbiffV0idZWX6rcIJNsKPdI4Ggsn7/Lgzmh2/04sNWA33RyQyWgXQUPsD1Jk1
A8THt9xHw1S2G71vxBR1b5wFKUiYhqZeMlKp9H+KRMvpp3H9odbRl3jUZRe0yuZe
YGSf7dFeOhEunz/pSO/rCP9jKA2LJe6yipIicFi1d5O2mCM5Zr82w47MMKKFdacb
Rk7/lEz+2uYfKqbwqL+Fuz5o3f+iX1g84DOZoWOGLqIaBlFvZDiWEauFFGy9TWlM
EqOTkyJ1masouEj78vSR/3jm5wiPHEEOyh6dsN4Rm9mwRwZNMLoTAI3CGIKuOBEu
c2NDQDSL4ZayvFDKmUgSCxIQLjGy7LI5xXwwSF/YT6ynOnAHwexDjMMEjod9lESw
us08t3OkiarjEwi2OnRUJLnCYwno3t8bBiMDrXntcJlF0NRJj7GzKg5OatlOZ2OV
BzjCvdxb69DM1QQNkziuG10IGuZAyR/GdVE5W0Ge13Qc1yjIJAtBc2LKvyg5a7hs
bLwiH3+ZsyilBYG69vcmmyLPs3oaJVlREbpWipOiTqMLZSnFOpV6wmbNmoDQKJAt
m5q8QVkjGQfsWaX8zM8FH5aBysOrKBPaGu5VJ2IwCnTTqomYuH7IGivSGFTKdeWQ
j2Ik+RWSopL88uRxsYcCMRn1Wz2QobSYuC7tUAF+qs8AS4ZDOCwSFKQAooNB7m80
WyT8NlGLkvrR2gwTuFcsPvkdgHsH71KPS+qiFF7y+68MyY0ulat4FHOq2fMAf9ox
ho1p1+LPhFhDewGDgrh71KBKjuMVIQNDon2VrLNR3rf1xESiuMw3vJcL/fuGbEzb
d51yE58nc6kyYpvON2QXvQrJ6ewARpa/GSHV1jZfI5JHVeuXFToDbLPBw7LcupLd
RhxuLgEJvU2kCsVuglhArSnJO11axRKL0fuA7Ohy4z0dJEvd2hwygrPLBQI6T+sE
KtXvnprEjL06XLOamRcDAxd4rTUGQpEiGR76KiZ+KCSXuc1rZ49+zCmVn0b1K/TV
6LSSOFmqEhE0rjg+Fi78c2UHq37jOwLkWxpMFDKlvA622Kk6UICqukWZkmt7JyR3
Ci52NXLNGrlVASiVJp/cVBkqV4S0ho+hYjlajDTJa1hGi8Kjv9O/3BZ9PbC4l3dN
61ywB/iXqU6F0HwS7/wWaZ/YkLg+D1oCiG7VFHgaekdbpN1NF9PmbqSVBPsUiI/Z
Mk1nz8SAgXE7anO2ZPA+5D+8UotuCxjHutzTY0nitTF7BaQ74EySGw+fo0IXhJxr
uN0pL3/9wa1qjGSTjFV6Nlg2TJ8H4GUG2A3i9cfK2wTeHqxrlkMGr2PeDLXZ9J8V
hDInK0ZMXEvRvFX5Wx0cInusDck4VDMgRbGaRr/MoAZcqbL85NtTW0F5+L54718J
qX6hQya/i+NQg1oZV1M9Kr3NUUyHn+Wo4bw3hUWwpYjQWH2oA8ad6WcQlO0y9cll
+vdef7fOZTOlp9I9s+9iy77mXAl7w9xPZdL6KQ1zUNkRepNZ+PmdhtdfYQ16Tg13
EsqEkxSdyx6qogRNPnVsCq9mFpANan2okcLW5aGtptGj9rY0BD34KY1OtbGheb2N
tlXUjUrk8dPcG+7pKqqFhed1KxEg+KeKBtH4IuffXOPAhYA0KODuNv7Lbrz/M38D
dzsXrxaqA0D4yofAPUy18Jh2nPiHklIl2zKmjXCAyFyRfkObX4kblfiXqy9hnQ35
VuGNKMfEcc2BrR/gfp4gAtF6+z2VzVaFSgqlhS9bCYfAbWIe6gM5sBQj9z3Onmnl
agFByuDVqGEUDWjAatqJZ1BEHhQ96QWUxwacc19PSxsLixTjcy1D1q/NGWS5JpAM
tMcUFdv01M1K9bpX3CzClbbaJQifKhcHJd6O331x2R/7n4AdV1cxW6s7+5G3zAiJ
TezRXMNOwMbTmtWZUJv+R7KXHxgO0j0rNdb+zrb5cnHLzoqfK63LmmXdQ+Ft00lF
64gRvzXOru2EfsX2a77hCUUvGiXmL4JA8u1uaWE7qn+nMdjgvCZo0nC8d20ZPduU
eW/bB7NtJxIOxpTZGPUfO0qg0vs8VUFMA+yAbnuWhadXMpmzPusV1R3ejKNbeflc
D4LV1owmN9Mfi/NS5BDFS4jsZpD0jv+iN5o25jpD4V//A7hpIqh8jFNfecuVfczw
eFHMBB1Bg+qVrJaoWCICj8xfeP33JvbAZc6gbT+Dks7jhpPV0UKBJ+pnrU8SjsPM
eYhi8XPRkpQkn+J9B1VIy7c275218ptEqjjCjFhTfDA=
`protect END_PROTECTED
