`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XNhU7FmJemmErsJ3EY6vhRzYGcm5FF9aYaPXau5ftV6NtyJnorhq0iVte6F9Wzzr
O36jtvOXZa72qQtPW4YJTSdlwkJfGLIGZgzh8IFYpHLxm85D/Bg8jIKDMrm6l6gb
y7wwn0oZlArDhs2z7DHuf++dyc0FS281ScKNxtrlM6hDkklbavGQG8WW5ST2zMA8
i3dwCrkOq+dDtRD8mSyo7SIod7Hk+hmuEGh9HTCPMapmVZdShHcbJR+6PbW/p3jb
thvgSwkjQKjJ85VWQ1iun2WstJDNtuTDH8dC3ux27XwHcLAvNFUOS4x1Pij2DFbV
E8HWcX8/Susdzprs40opGFSK668kbccr1kown8OcpCA/KWsphGnIJBZHpKa47qW6
fOfuj92I/Cy8fnYVpY/har6m/pYu04xZ9sdP6KHFnjdbyiuBnthIJ6o1zw+t1rJP
P0YG8uCOmkz33CEXmI8EaaityV+4HiNS22/rTmhptCloYn0w1NWBDtyaHKeIhQBM
hLlMKznGoS9RGQDUwr7v7fjoC/bokf2NQ9avEhK758+Ehm1kAXPdaT1ED+dUMsYX
swvzmhEQ2MG9DWFLrbu/PaEmEloPhLq8VvSMyHAds+v4sMLCP2KWNxJCgnjfaOhN
J3KOmg3dPxzkYyRd0jMiBMJ4dCjUUDMa4ByKcWUjFMO86T6hv/+cDgWsstID1lvj
m21ho+b0I6EXOmfrIyTIkaK9JlZrA83mjgl9zHQ9WLetumptuTIevd9TUy0f4A8s
u7ymXDSl86AVrfl/zmz+4p/nQ+1vTvSWs9+YACxIyKPE5Nc1fBm0Dgu366EPrU1C
IRdGNv6rfXC6EZb3xvpSMgqZVRiYAF/OcaOt/vjrPxXqntqo23njrZ4McH2lhWsR
+lX23VQQ03UxPm08u3goJuwb2oFdL9qKvMsvbGADt6FsaQW/0VKwUQIb+pjiZh4q
MS5CbT4hF7I/+VzphysIcccuelToqb5ZtOFSxbTxTBOYvvbOkU8zNXIKTT6KS7p0
RfyX++lz4G6s1XsTjhxXd6qWSpvzqPv6oAdp8A/sY8N3AIutq5MUj3yg5e60XSh9
9V//hxa3+r/3IctiDIxjLKSmQe260oyfa+udmOLsdGy9BBmjXg4Gpd6OYRq0a4/7
kwR8m5ddKovZDSD4iGq47q/g+DGkqV42se4ENiycrTmiAqDd3GV9Q+5GPXhqKFxZ
7vJCr+orS6t/CqvAHW3lIXE+/qD783Rg/VngofS3bVZDV/1NYnEiL+i7OoinTkDw
+x+5L5m3kKFk7JIDhdb9GZoxqd95TQEHnNhAuBHmC5/gMkoPYgF5XFqx9PIa7hvD
uKvCxMv3qr1/xbVDHQLJGa4lLN1C3jw7HPjuRJJrRMSSWheQSsL1ao4ozM1WBpHd
WkEBibO43UOT/J8u3ODUeNH6jYSnyFrvjBorHORLGpuCSS10H1jt9MXgLv11Nl5k
Kcpd8CvYB2FPeMzhFZPvEv45mL+oFA/moc+37icBBLW/Cz9necJpLV7c7PN8Qery
nfM7vcVVQj7mSHMZWXkFFm72+ZcPIy5xs3CNWM5zUrazXm0bKXtjTLU/g7kQnoV1
n9mH1BgD8UsVlmhEEBzfE2JaQTnpDlC3ZU72Sgrvoc8RlBvI45ul2lEKX9BW+Nhl
/yP8ysXZbkVeFiO+bGgH1wOqchkLEk/XKuO2CSJAlYrRauPpd0IPLhzAvyF+bOW9
wVpHeYwqBBntv/P0c39MxXqlnKVG9J/xYFWKT+rYbGusMXN7GhXz+UMHB38L2aSJ
REw9UY0yEo0UYjpbFShSIoPMqazJXlCKAPG6QyRJa13ag5mOJCimUCQDwzxP+dRX
mdLlC/DVGWpe8if3F9EDDD1KMGhux9eMRCvG4I7BhYQE3y+kZSKJnvv9EJwdokBO
BtpmxlpnaD2SYZ8/rZgnUQllrwaF6T2NSsnUiCTAScDAbEN7OAIhUHckiFMvfBDx
zNEZcvotQqiSilA36fywCbYg779o4TOMY6l3KMO/k7JuHMJunaVpQRJsjxRMHQ5s
MOuWP/VxFeUmn0QPg2335J+/XgKuKHz8zYsPynQ5639vcwvQvIK688VH/U+JX5Cj
IuA4RUMljwv276qjdEzldwY2wrqzUwSfoG7hYMVPjmIe9JNSwJIXOyPBXN8usQbP
+kKjRz0McuX9UgtZHmX0KuIdJbFzCTLAn59+qOv9GFNtcJWyrKpONeknpszzFvDu
G8fFXmZO7FsCh8rFBCHU2oHAGf1oFjmFJS9DI38gPsJZ+wKvQsUoP4x0lrWZnxwc
RQgCjKFc1e5o12h29oPhfPSyffjd60GTGcrFmJnLlis4hY/BPDGwv/kW2EORmqsU
R2IihRVwVYgJhNuPhIKQio6ZvtDpFoPsokq9w6BXkndFZBoKYIh2sZGg0VEk4ZCW
rS/YGhFf7TGyCqLhVKsDFsbAHEw+tXAiVwU2RgIycq2YQBak/Z9rQrlW+npQWSQ9
or/HduRcsEfVQfxjjcOrmC3Ui9zwGm48Nkvj8HcTPSzD+L/QqJg61yc7tTUxBJ7h
LMPxXzAbLqQ4sUTsR1jGa50bEc29sAS09EaF4gFYuiakbwWaoDjZCc+60j3k/kpp
IQNGECCdxZAJRxJVZCJHOO7C2v7BSFOfBWXGIFH8W7PCZQJhBOirajukTl7AccnW
FkeyWwJCy1lvl7YGnJDOlz+zRQ7Oi2Lu6Bfyggr/LNA=
`protect END_PROTECTED
