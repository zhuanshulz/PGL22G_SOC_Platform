`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dqv69fLkYqXVWo5y0mgykE46N/lwIM3KsPLLr1xXhsu5Z1DuDRWer0NtuMHy+Fly
wYer9kOOvO9WO9KXQwLHSKchNpbWnUZ0wXC9UrJjbsOnos5ukA8rzSw3NQKofq1P
LL/Gz1TftwkwXVK8DiDGysqBQRXnGNwL5VPr0LV2apfYX58cKRem5neUDukgG5jl
aoxR0SV4fiwFYaod45AmrDhHLlY5wWe6F+fcR0YiKQQAZ+1NaWK36RYY8lUFCv8N
rTBfUhg75jiBXBOyI6FIfS7++bW47C/xMoILx5hhSgtVWSPgcei+2P67jM1GSAvw
hgmeJzkpCsqUH1+iPkye3RrmYAYKF+Lh8wf8IPYmECxFQJekd00FTXrdiTyjfJll
RjzHMIvv6f4hT5O347N8AJBXUP0cdPR9nVERqAJwVDduOAjDFp+TcV44EWTnOKnZ
hzen8g+trth1X/sm4naHgmQUYxr52gdz1jCgq8YYFJab5VJuF9lxA4kJTc34VOHM
s8VVCqU8hBHlXH1vOkk5LH1GQbqg+F2uT+pSYO1Xt2kVx5c+UiHOtmby/yYzkZdy
uF3Lfd2cDrQB4h9VM58dCeT4Mfif/Wimoiv0mw2FhC2cvd2Ax293Pt+OArtHaqxs
AmsDX/qknuIMA2Nx97ka3ZlwmFQPJJ2kWlLMd2fsxiPvO1f0eIwTgm3K//OmFpWN
SIBiWyyNxMhxLsBuRYcshGMUhWihXAjcj1UFb753raI4Ai5Qzpdnez/R5RjOZpTa
Wbghl50uNXixXsIMXledmvAf9SUPBrdwKuw5BM0LVkxEt3oi4RI4wfQlmyNYUk94
9hKXJ+e/peoawwxm4SP2R0rkAodmBMBUgSUI9TJ8ULrNGFV8VxrFgF6XcZOchwGQ
gTe1bBnRYhB/SCMFa3ioy1O0GRgpx5dsrHVmtsGU8Y549qGiQF9tvxMWTRd4JnB7
8cxCepgC8tKjSZ+ymbCpiCLRVOlseu7d0K68wETyWFo=
`protect END_PROTECTED
