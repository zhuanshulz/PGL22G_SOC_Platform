`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mCkHsR3FLvEEGCYoRS7Lj0vjX3W3V0z8SzjlaOzhp9KvqhawofiyLxCYsGDrH62Q
5P9K1vfAP/z/KCRaE/xOETOztNwpdWc3zmPRi/E49NLjxLTj4kGj6+uujZ0WEENW
zRogAFa/HAJc8US5GKpoCPmq0qJXu5YJbVWHxafU2Mwba0K8n4S64D0VNn/KuVoh
Epmf/hp1N8t3t29g6vK+Eh03d+H4WC9eW/0x2Kh50mQyF4pWPyM0sX0uTf+QpVPE
uhbvxCB56Irx42/JX2Jns+5U+4abcyIFV//New5OUtiApkntj50hOwXsZwr9iOmh
PZ8lxFpScWGj/+Q9dINX1PKugR9keC8snMTy8KMkpH/ZNEWrsSuHcv3rg1fDnm7x
DEg7Uw6oUzANa7i/TWnNK5u61g3ySFAeHI6VDenGtLCVqEZq3jZxNdvk0FpaWpww
d26Rj+ZpTNUsWMgUca2SMUafPLsRJyGFsvLxJm1Ifr6mjTIEO0zrRHAmxunkUFG/
/TKRe20IDr9Ium6dt2NmraDZPiNSY9wyRb9ayZPqYUO2hiB+lI+KfVUqcu59EhqB
hqnFX4H1Fq/IySUUV0hmCCzpOeX3jshJ0+/wkujcgMrjiOc8XJEVVjIRnueHLw/h
SuovQMtIdEAgpQ3KP2S053i36gc6JOu5lEOZsBrmbdfiZUUjRC7h3Fzcv9RzDIS0
1b12WLsy4stahR7Qx8x3ZeQBmgUEaSnQKvgsK0UG8gzxlrGPswFhP7ChWVYs2NJl
7f9o8V/erIVSbKrz66ReeY2d/7eUrOjEdElpWyzTxwPJlYNN7ed0Bz2aRec3gXaS
dSVDCv5ILkAhRUqb2yVEQDqP09tsYMI5iEikNYNM3bIG8zehjNKwvWmufIRpOFQC
aDRUwFaXnyxJIK7nw97rwlTGFwaiP68h3YKs4kUP40eW0JCbqgXX8OyUF9FwbsOu
dG1aIXkfTbwxONMYIr6uLetCvz8AZa+VtfsrZOyG2WqNj++dwPgcJXE6P7Aj3EFy
Cm5SiFwckqJTrprjKEbfb4L3wdKQTZODx5Wq0o/bDSiBwN7RzYqYAC+faZfwzbmk
pt3lnnzS/o0LDsFlpH8Q+SdGEWHDbnkOKR8oarRlo7ODc1HwsJ4GxsPeYOeJDDi3
VuCnNvRkB4IK3n1c4RtM4NY0jsKt0NPtuoBTwvo9UY09zkTqyHs9rJ9qHfxOHSfn
gNRfB6NypR6n9e7wkIqkj24uezOz21Z/yd48iSCIyP53ls8ujceKmPrxy4QByHqo
1w8ZeqQHJ2CvgRWYoMTrBqZi7wQjAa5RbEa/mNP2jQaZhDoFlIj0NpmVsQznuNsz
L7k050ZMCU7PYUvzd9Xs0wCU+wk08sDwGjW8CEwBP3kLqXiSMI++PaKnzHGeCwsj
XOw3RdiKfRKV4dktpk3Z+9fpq5Zeok5CrdwmYWf4HgA0LP0fAB4+EA74MTU987ek
g2XrJzT0CZCPIPffxweSWTJfsWbNH1XKbc8w1mp49QF5U0Lx1jpgGudHPBkCLLHK
d0U4H7eIiO3zHxerE7rA0IEGRGCpSakBA65yOf+GztNkub1sJZLvjo4RQ5MVSJN1
mk3boAst6rnfoa/P/KHzqC1PSSdV8EhkR9SaWxglFyuUeO0rrtF0Btf7RY4A4e+5
2LBmPfV38Dp7ik0MThYxVgzjEzoEEa3oKc83kCIs5HYfIs71cQpWxJTqHag7aG1r
PGZ9aLI4vtSAfIbVrzfk+3lKcjybrttvUwlx9Ymv9ZKAPI7l/0bWWQkBiguanux6
qGMo3KV4Svqokqdhj4ZWB6PVS86gNJejC1BoUnGML4x6CNQS2Qe8wOsr6PUhC/iE
itK+aHrIIj6gLB3RWjsHWdI1RmwevSxvt/bSySVO+v1zozbohXJc/IewjJhN7doc
ZuDXORYnlUV5GWHZIcAB8Tagp8PB6Q8zELF5QOwjotrMvT3084TS7Yzzn69CChA/
EI5xMRN4MG31fT10z3MCkTlqD/B+oR1cAqSTHjOonaeHy7tNaBAmIz/cBPgykQLx
uYf0UZuxDBpCisyRNmEuEKwAA9dJG7dQOmzW9TxtvmMwaUmZK7yTYMMl1EDnZrSQ
oDXnkSQSxJ72XLJnPM7Ro4sC64hT9zl8yFDnOaYWRrg1l3Wvex7c8UmIoTK3+RTh
mS069jUrhRRcT7+86hTQg0Dim+2qlTu/9Pczv+ss6cM25a+vAPZ4TnIDKRQdF9wu
6lbeqQuiIPjGjL5Cy+lmew==
`protect END_PROTECTED
