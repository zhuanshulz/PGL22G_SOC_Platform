`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0fJfpYT/+EKeTcuV/2vyAHRKtXvEdO2xEmlcNdRnJjRd7ZABj6nIzUbSGDg3pmgk
0C4QfNu+ztAbac/HgUgprkV/yoAlveX5lz5QDzuzzcnLbHP559Z8X98edOoMBsFx
tMASQqomYDbIs61BzkggjmaVm9w9knEB5fZwhsuKJvfBxZswRqxRjf5Ghv0i/WeH
Ho4wJWA9r/X31JxhrXRENIpqWTQTJEFc5Sw9uKDGz71KDRHiYAaQQFMheA582HTQ
TklhuWgWFEBlH9+admZC3YADTDZ8PCYMfh+O9JK2gV2CB1FZL+aqSYavD4JFelKN
KQTp/hTYUzkGCURrkrCeloUjjYMM9NS7w7qrRlIwcrkT8/RuMKSg4t6FWmSjmnOo
XmkWPJWyeuHgYgSmOOAK/l3qvzlsY++wDQezdI/ijYevu0Y+4t7EMMT0HOg94rud
PypKAd9zKlmj0SK9YEldB+VErs/eA3jfrGWoh9V+icWGpwf0Npwqu/32WB52dG37
CTTcPrP5WZEAhfygYiyQGKUTC4J9FewDN3zdGIjts1dIRWYicmm9Mq+c3H8B/G50
haylKv2cMQciQwXR5sGxX9VwLNJUzKzoM2GTYdMi6bE=
`protect END_PROTECTED
