`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SsU8zRBGdY81th0I4nXS9pwRczJochITiPVDp5MBNE32dccIPgPiAOyONJ1JU7hu
p6XFrMPpQSRKtkBGlCGdvAzkpvgAZl6m8dsYl7rZqFEUCYr3WQca8snCmFAIzS3g
p22zAqVehFU7ris8sG2FNMhxMUM0sR4+vWfrl/0y51+VEhWgsm5164FGtJiwSQC+
V+LLmPdD/qmgqu53ycS4nRexUkJLClX52+sSwsZEVFQQor+nuXWLbKQvV5R1yape
uYxAbdJBoUf1/UzwUAPPEmQQ18ZitdLauLkCQblCSGI/HJ2nvkphKZ3P6LBAxTar
UVEL6AkH7Bcr7xEPOriWwhNZcfGTiR1qCpmiazG/8x++9JEYg1YcRkmNCFzTemWI
53nTb1uYEf7DfY8yJBgYl4hwjI4VVTtQWsiMlPgxQYAD9yTW9m+X/Z49wG+EtJ1S
ptMyT/ydq7HfvfZn+zDrpnNohy1uEYilNtf/k67fgPhhxIu9xEHxqyHisDA54wgm
BY1LiLNMNiy4vVDdEJC1ptnWr6OEeaTG/h2MDRWkd6KnDbnmVZ2v2s8i5tN96W2J
P9tsCzHSuNueCy7szCC4YhcycJsnhEig63MyZd4jr4ifO7/ka20n1XNYZNuNHlWP
1M1oB2VgKlM6HeHMFnt3ZSeeRwoFe0vQ1zP/T5IaCdGQ9c2a0C+PptwwTY21ix8J
`protect END_PROTECTED
