`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UgrOSD453xv+zWIfa8NYUJyCWaDMYK0PsvV+x+4N5mf16t5WPXLMa18TffSj2oeV
XB+L6WdD68/5O8UM9mgj6dbwa0LKE11XBAAPtXNrhqjZ49Jl1/I/rATLVCW9di5g
h8DBdTtEHIbCbkYWgsAMteTH9wLdILUE2UE7hioaidL5hpIgr9FuqD2bB1oqhiMa
OHUVMHt6puGh/nwXX1jRrLcx3etamTNzCQewbwEZDXHtezIFt19yBIDIiAr9lfbP
sZyrBtfNt0yXPz0l8eiRDB6wbo9xRR62D+XrcCAlCRTDNqyOgOwLuVObuuzvgicT
KsCrkJDc4M/pdQ/AOKESkKN1ZzBb/plphZEeWWhgd12dVmZuXQzWJUCkNH+Fwv/p
mNLbMz/yO/dy6RO+Gf6Yw+cVYzCKekk7F+iBJCuOKVg67pR5lYp/VZ9ctsCp4GGV
CWiO8kA0cuUsAMyTKH6jLRsAX6n3AnfNtrC2jUSEFG2A7d1vvVoXRpvWdl3VwPCD
5zOAWxALHqOzOodqDVVW9AmQ6YjXWuROlKjtxQeN2nqg6C6km0w+1MZrttlaf3+r
SNeW5nxzkAOoH6qM2tx/5gqgqtD6JzvcxfP0BEBIfgMVk3Y6oGjazZUZPZt0lQQz
NULBt+ZL2vRskxfXEVV18u96+ez99EuBEmAD6XXxVZRLXh4TjHIkbYv6v+q+LimB
qtWIw35jlJN57l7h5zOPBD4kPvIJ56DUSF2fPdT+WG+zCbh2nVBETddYvHuasnUL
o4rXfasHudGCM37GOXtggRB+QE0Z11TPQbmk4aoCagNiRpnvjspgW3J8/DVgxukt
2+dnl9nltIZ31CiqFNrVX+KWOWD+tbhKPT6sR9jFhLD8Pa33NbSvKZU7IhghVUkf
zzm8zQz1KBTnx+GnyC7FZP52oPbNOT76OTJzf9dwKiyjl6ObsUrIbIM9dw948ag5
pLWf2DpqQDgnbnHgQ/DSn+e054m1uXACnx64/QV9OlQm7qzuDIHNSyYVZ9I7Q/9h
pNXp0MOg3Rp0SrvieRdOVGgoGzxFiy2+HbuHyPgk+WNyaOfC94SfbIoq6LxisfJc
vAf1qnlbHxtWBb4AzvjDQS1943r61pVcRTLgDipEMDSjD/fh66vOY9K1zA9G3QxY
09Yf0Wap18NSyJCUz3kbb2Bu7HkoMoYRKAVaKJ33n0ITUBkQzmbFlPWM7PpbUaJf
4AktM8DnvKvoOznR3rh3fna06uTKnJlL6chk8FyB9DscKna1dFLU4kZsZuvStulO
jL/+3OnZc0vBzFPugaySrEqwNdy7LgU5DV0nN/F8FaOATgX1i1dUWyOzI3nu3grW
l3sCuFxjlsiVz/KTd/OtOR3lY7jiPeB7/W7wbIDtxyDKRJQKkAuYYaoKXf18/BvA
oEgzZespHgrmb6pqSIyJnALm3euc2g3jMqRtu493onIRsXPCwTwqyY/EUYdFVnf8
FceKzH6GtEsW4XKdgNj7jlXirYXkmwl2H3x17Cum8tdTK76RiRcap3+fUb2bPl6S
I0VDce32w/PddLQRfY1x20B9RfJfVHuYT8yJoMob69MoXLVAzWakOJRvZ5bNE04J
/VeW+0+ZH411QK1GN0GZb9z1b+FgrDHVse0zVhTX4+aTp5dByOFPjWWZwXtlywfK
eGzs5L6VWyfYH8DTpE1KKRe457xSV7euBuLfhYUHATLgm38nCdZYLd2iAhNnVVaQ
rZus+C2ONQB4fx24cQ/Z07wOujRf79ja1v90dMU7OGdNAyL89q/iBe/WHdmjut4d
Ud6nIm/IZUsTG3Aw+vYuU63UEbpfzO52qUIpw0wf2hKntQUQMQ1DIPrKg5BneuOa
1Z2YjuTuGp7I7lL7WMYJstjgOIwvnn/bszD+mnUkfXIj+2fljIhbU4xTQ/MCPqBR
tJEdoM9xF+xm3ZVNPhM7Tn8Z1xLq0nJHbsfcbSIuaLMbz1FTIvMAFEiYMl2+W6fZ
th+obQ+X6Wn/s7KZ9aRLJsWNXkr4Q3THWpK1rHRTi1szoKCX/T7PzJD8yrj51Xyb
fkjMVAj00qzM2+17aZZh4BKlhw6ZDX4g/oWd0hHmwyVjT2V+aRrH22+FRIW+Tuv2
Qct4kMT+m41Lel2tMVvgM3vSL0x/UVsdlWjAW9T10PVZlx035qa4IV+rsnq9fqT/
wOJ9nINTl4r0RwbgVVtDNpJsY7J3Sg2qs6kRzY+jWXz7ubwiE3gTeMfTHp7Wm9y0
sxbt8+26krlLwbQ/9Ot/1vECcAJr3EwYt62BOT7Gu5ADG/4FJ5cDZ72s8STIRt3/
UcB34Lo49nLsTM+g1gs81VeKV0tzZr4yJddwSj5z41rFGyJc/2lYpRRxOvgi17VR
TV7Mh72jLsqBRa1yxkngxr9296hRdg9UiDzJmHNZ9b3FYaspFXO7fYycEGorxmBd
XdyIU3pcb3VPTIlr3X8FS2TwpE/1YwAMZDNDEFQRHXuydwIl6pSLRwhCAF/JmcQ3
Jm4awdc9jRgynloInSJeTn4Ul1ophxgfRkfck6UULLM/UeQIHD2eATnLmmdg4IDb
vYSSvYTZH2SU7xRkXVX7gdfFRFf8cl/f848K9K2M20w5+CB1EM0nGqkMz3W+ubWi
IXYEJlz6vocvpR8ENg/XeLlbZVt5pBVmJx6ck7pzRXlnzgnUHwm8IXVc/lEA2c1+
6sdOROzKRM/g6aEiJ79g3Uy80uadbtmTTjytGWe0YMmygpSU7JPaySVN/d/N/Yl4
qLyGrUW5/Gdz6Nwrdv/Yv5p2esOyYMC8Ty0SHu+9nkDJ2s913aa0D2zInCcgfK9G
NPdtPQLQevLn7UDWI234wXVKAOWltebzmfQy86T9YP0JoI6wNz/ERFW6VsjoJawo
5u+m02luRvtTpVnLiXU2H8JIIi5Q87vLQ1PfesRAeJ1Pq60OU23muOkB/tOh+vXs
uif2p3O/MkWiGVaVaZvv7V4ibDELiLFb4ScLFHc/Q3wSHw8sFiLBFGJe+eJDcYgu
+Dh0gzM8H7/j+m5R+3XyRZhYBKZXlgq4PRIjCJgakr4cz7ZGweHfdyAibFakV7aH
2qIBjxL/wtK7nwpyWnOkGXy3o5DXHTgQJljm+NSxwtusa8OD+NTJbooNgUhvXZJP
xFNNy6t4veJJJWFOzXc7TWemQ/T2+kFJc3U0aXrubNb9xV6vRFgI0YoQxNAfi/5J
7WUHbGQvPN64Pts7YRuGMzwhiOZVYVp40ZjwIhUBTmub7RZcxZKlVOPGVb4nO9fd
bXg4N8BlxAbyg3KDBWnLtPwJqGjwXCLh477JDiuSrpcM/DeYvXdXLw3uyGIbxnJp
TwMqrR5RX0x6/lzJJhReBQTQfZzf1VFJFqns3q7TWuu0/jy73wBYB8G0LVYBvCVz
65EDtRK/0Z+YzaGG69lxVuhk3y+PJRA3FQjUwF3alvIgAnFdxl4wwxesi6CRByPX
+/ytNwLCcu5B5vwp3G9rnaLm4nJX2FvvZSpx95kB/D8s3DoJFXPvwUcy/dSUBOwm
gyaS7znDWimomoXv4Edtu+5yBWUITSSf7B4nSp6OR4OUtG/Q843jCqiOyN42ctX/
hBUnNu12iyFuTeisCiCOEyumWW2FN+BylBD/o3Q0sjAJDm94hPD5hGTD7bk9fC0Q
c5mrQmvYHsywC9I8VkVoqdP32x3lLV1PFqKdAWsZuxQwh2Ne4qA5gDDw1gxg5fsT
/9nnGoHSt0v/hKXhRv00XL5Z78ocFcSv80RkvgWfuTCpDqj6JMhltuphmj8yIvWh
Owt60F6VPoyCdWWBNNfG7cRhoJ9E8knThwF/bbMQctLlAUUscHFo8KJveOt7F4ym
V7iPGzLThli9K+PyAvBbLBAT+KKbmc9oaX23qzYoa6l08pph5DDEXAMlTlPDu85A
`protect END_PROTECTED
