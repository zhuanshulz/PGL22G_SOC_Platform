`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CaLY37GKBx+75E15yuZESTAKGrfkEMgNSVEOMqPfRuxxAAhBmQXR1IkJ/Wb/VJG+
qu2mt2R0qsdYrQAA62MJI5ROGMvfJfukMLCdkMJVuA6ZxrhMCo0buTDFguBqzGEk
rA4F8mi2dhT6W7RaISubzJTIpWJgEBKz6LUkW6xMZenH7J/f4NsbMGbq6N/kvGo7
UGrXkTSuLfR5XTOkkYpfQAfcJC3HB0uQkzuRHTrUDxo0gZ9BG+cF6+3gmV92wyzb
wc+VNif4rAiPf28R/rzwm5lGPV9P8UWlMOO5qLNSG7BKyvmnO+peFrn0U82hUjqT
33C6hs1kEIUEqYVWmG4rnkDXOLpkIrbYFuvhD6086/D4BN/4hUzM9Nvm1rXg3dg1
yv+N0TZjz239lNCaVHeVPXDTs9NUHp/NXqTP9RyVANz2V1YZHot/JzCmhAzDKJPR
rHmfxn/P1x2OMhiFYK9HwaEjina/N6MUGGjFKCQ9FYgFEPBMWqTlyfQFmxiy0qDJ
hJaZJeWED1i4vKGWU8NW7kAAiFIViwZgl+BCfAgnxGWXOvbKBVcHk0empPm+K7Zc
PuUwlAWc+RzhWBx9cRZpTNoih/q9lIpFT22oOCD2+bSeukwKLU3bx+1WLr/CShFX
prdY8c8y/3XGBzSmqCn/xM5GBK+WyR6NaMV4V1WXMiUvBC/eToTZpaGU9+qwrh9p
1WPyaV9ogOehoEScq/HJv1YI5yjQ+V8piDqQWZuTV39aIjFs6eadPz287gIJ0xPi
MwmCqPanwUqD60NcXpb1aw==
`protect END_PROTECTED
