`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qR5vxBpX4Q88VPU+KW4VRnxB4kofyYqAqh5K/WiPIoS19IUPsRB3eQCICjL0n2+b
jB85xIedk7wCM3uzxEJrvXrX81xL5/PMfbw1Esr0gTJzGgx8u3zA0se+0kAjzNhe
2bZmAymZzWvjv+uMdA8q1VE3rWiXe4/psUe0LuhzBG9ZjGGwtmXOS+nTVJqOAsLm
BMwna5angtz2yZ8iTQJdMgHaMLHvCGz6T/dVg3jTzOmQ6nAsRRe09Q7e5oTJ7lfW
364dFIMaVTJLqTGAuK39Lg==
`protect END_PROTECTED
