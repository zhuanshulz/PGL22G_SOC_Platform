`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
boX1A83uwPWfrFrWC0QfosCMVz5UZxgv0GHcbzw4oshA/v8wcZqs1tGN+gTfmQL/
HHP1skf0SXIRTD9Y/FolElvn3TAREfWB+Bx2vD/No4jKye0N5gq5LmSowsGk07Hs
evhAD0YjTAr58w0YRIHiaT6VIWdZ5ixgBSXV0HGC+Q0w2mZ/vP74/THwd5jCtGH2
kopDPVaR2nEvBsJeSUgh2PVhwASSaqxGQ+soudfs00Fc1EJ8ZlOPsqZutOtrdNMy
CiwMWwSyPokFKZ7bSw/GjPDh/gM7d1DFRRIwAF/fm00IR330z2abT0wkc2dko0X8
kvfFM0BtGqooWiBqaIZwiSJhVL59PNQEiJXBdWeLOzKGT4huH1OXUtaMlrgf7BA1
THlCT0Vk59O7ITOq2RDRSo14TywqF4yaA3qZMHXrWBmolVqGoLA5cKjphsMgMoJL
tb84byfUQ2r6RoOKNwIXB3AZ8xFkchxjiCILkmwdqp5Se/WvoSBpv4vQP8yTGTOn
yhKXTZ8dPD8Ivq069N3o4q8YiT8l7/1K/eE7F45cTtx5YIu7ucMS1lq688v8TTIT
8hYes4oC8ncI28anFxjNnskYDnUVSrpmqUMOEWD0z0qE1FoRsnGdCphBgnIRmjdg
RJArQ69z6df93ZBcQO70yPJhevQNx9ZV3JdY2B0X76XLnhCwuyd7qYjCk7C1O84w
u7yIjLT5P5VeTKhJTZEUINLk353bQWB0OgDs0ofo8GohX64//oeakjWpZbGMkF66
K1oNdLg45gu69WCmRIOKi5zq05EODGrogXwFaO5HimxRxcTof4ygQQmrQQySezIv
BAjf6OhMpP/0s7huVLcVS1JbcoHC+jrU5BmAGm+jJFRMy0DmpU2wtnCeatLXX4jp
+4Ic1KM43LqDo8D58hB+q7PlkfHbPFU9DV/8juUoh4NcsdDZp//euNsqQ+I6TcYF
uwq5BG62EyOhQqD7Wq82uAePYQaisrf6s854aqs6+XmFC7iM8ncAKsIXTwYO7251
kRIosal4pA5XXk9Hn5MWWZB98nMH6h9/Gd0QiDWzOzK0wSeVe0QZcWYmtBfWcYoZ
d9y3BTh1LbMTFKjsjQ1nFmD621KfzUNyLFQCCm2/We92MoJdIdVai39iPo5If0BG
txGinJ+5WmrO2BSimK/5bRtu4OxDrbAE0n/feybB2OEu+IcBdL6NRlu3G4eMcjKe
4+siuWXQDSkGjMR7+lHY5BWbKstq50HHMj6mMLE+M7RLu7umhB/7PHqTmyOFY1H2
OkH8AEJa7DRiDhY2Q6IkDvpOqzFeg11G97jgDzrssUvhIQMak63vZjNEUXG7O0AO
EYhPu5JTL7OHN3Bu2ViY6dZOjnIWxOO55jUr74ZE4mZsB5q5w06s+l5Pdg1VKcMa
/M7JbuLAcwoLxD1TQa/AbkCW5cgECI8sTS/vbX5hIIAYwpzM/eDm0wI1+45kC/cr
/0dg3HNV4hUWG+uvGQjFPS2kHpoR9CFzEDA6OuxI0cyC2R1P0WkspGFvkLxOczj0
ZS4LyUQ5ZQ1JGGcvYOIR4i25JOWFjVLj5J4/faK/s6dgpCcAoo65bVvCwRGo+YV9
+36yGmdahDX9RTeo+Xl5ga+PkUC9FJya+5BYviN/nVY/mAEzKSTAFvhmoYmVLBdL
vGHw4tkPRWnSHxZ+lZRJOXNuX4lNW47apT3loQBwNtk=
`protect END_PROTECTED
