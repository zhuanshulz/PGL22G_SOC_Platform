`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ShibPRaMeRHZB/Kp3ZgKnmZbidQdRMUH4cQQuHTpc40w/xO5s0ig2rU5z9Ym0pKp
3FawPuZ2uI80ecCAoP+Vv4pSKydmBFRPltD0RMYSpLIYEpRDlNif8yMSMHbdcDxZ
cP88B6TODQCzHNB0zv/ZPnPT4/Drp0MCabpENEJo/K0bBQSHCjqmm54bbDqFjV/e
Hp2lMKStmxqEpMSpab6Sqt0EaXNAhE8pVznNAtd+eqA3zqAKAleg9dhmHa6uv2yJ
m09Sc+b92Kvw933ZdpBa2xjXYgieB1T4bKFf221QpMKA/lppgIlsFwzSxYeTsNgO
3tA8SR8XW/hKoQGUqGVHMzWWvamacMecRlY+VUvixIIfAE3CIrM8fyZylhhYO13C
Ks/46JW1XK3OpXCYug/41knJk8GttzmhnGeuQNSTaWnKawB9SI1JEYGkcLdV1f6s
oZ+m7qouVFMAKRlgXVpRPpRyIYkS2VnYT5oo35Yiio2TQluSxCsajxeQ3IJjS4V1
sARfvj0AdJ9efwG1UfXWEL6UaJnh3QQ6uJ33DqFvt4BCm7HVH+zMAE2XQP4HohIr
L9sMvzHtPebDgHB1InSmU3SYGpcjhmvKhZdCpaRnrMiG7SO9j2TWHfhf6t/gcYE8
WgdzbL9fke+BdKei8eocO6DQlZiMEPx77vkZnYCJc1fxzw934UL/FkrMRtslub1O
7FknUU3Ck185qdySX6VZdQbMoXNJNNIKTfJJ0sx4JXMc7NNSi+UXUslW1/RaA0+V
gbSbd1WIlAyUmGhOFuB2A7epXGNZGvJ6mEUE8DNM39qk69AenX7TPwztEB4h5Aqg
h4OC42/AYRWibNeIT9ipTjZCaOkkBNdEXaSH1npGl2uuhUMr1qLE9SdSg749Qtzb
Te+wOHqoxeYIVbXzPKapa2AuGFWc+tC1y0q+1o7S9XRQhFl6xJqPdNzk0Znng4Bm
zGaJWvNghT3G4XkZhWiU1qm43cYvKbkXtzEvVtJ3E2JghpGcdUH8INevf97GNdu7
kGFGWJSVGWng+GDLp9Wc3sPiaCaVSkjAEKXQuRHFsVe4T5hjSLI2dvujMFLWlNg8
R0pvvqd9Kx4CbMZ6N5OgfUCXpXIX7mGmuNqyyE/ycHAFt2P/EWIHDUfgJL0pQxtQ
xLmxl71OnTgKkz0PIM89YMWcNVJustqodCSzFoOu6amM1xXLP1ko1CSdeMdwOe/N
K1M/45N+RnjNl71Mc43fcy7uLe4cjXz5TgG8qWMKgG6tQGD9OcpAW77GClVAc/lA
6n3hFldzZINH4fYQwKTThswEVAOa3ZuGrLlLmGHCHK9RMLI/3Xa2trNgFesoXkfZ
ENxPewfk5jRBP6RKp+zKD9HoGqPndn2vVbxo4FyjJwUSD7Xrtjw42JHLE+PiRxop
fO8YOAhNpBwH7XrIkZWGPSt8GXtB8S0kxTdivc46k3pHbTQdl1EdAv6nKMFZGpVm
9tnqDEP6Q0V7iDZp973FbDvQmytjldn5NPFXYNTQ6sFvO8/Jd2xN2buf1KSMKr++
1GiR6aywvSvGFVr0cpJ2jQO5aT/iLsDHYWrkWp0X9uCXtaNcDbwAp8aRO8dOZ9Hz
vl7gA6IU9syidSk95xJSlkSI+N54T2Eaq1sFhYW+bUxqnnwt6zydz2HHbQqkGgwO
CUuJiJ9zR0cL5mc/6W4PTggx1nPhRApTCORfam0Qt7CzQTDtd3+FjKsNnOPlqHPT
t+YHs/5J556e1G9Rziuo6w9U40PGDSGQuiHz3VSHiihLvPHAjnV6mPnKdV8VQB+C
ro4gP6nXu4kJrzuYO2bJY5LzlNNKLR0mh/vFoZgMtUUXsQomRw66sepmeBNJnBO6
+hDZeHOfXXReP9sD2IhlYv4rU6VM2CN5MkRdmYURLIIv1WMPegM2z/mscrPtkz+B
NCPdAUtegGU4yY/e7r5tfDRGIjbENtPrbNesv/dDrowh0PDLqLFEwCLHaDLqq25M
2HsTrfs39GG+FXQs5xd0AEYiyHmWP3r9syGl3lQn3cZkFQbbrBBdwM93KhMXdH/H
h0LzBg+Mv3dAS8kdVa2Q95YRya++Lax6uLH5kLGnhqWMZUkvwEYX4t7hUu5YQfby
oay4IMlhMmsUiPNkxWgPrNwcrYsitDSy9NnQGGZWxI69Vdf5YOoSWoba1sDmoACd
vsAexD0u47j3vzyUfEpdIRQNQiJZ9u+2rXTGm5lSgW6uUy8RDDlU0mnWwZ6MQASj
LaY0ERRMIZ7Qzqphgo97MYycm5S0d8v26LqVd2ZWRD0Kfiio8g55TxJIq/t3kZPz
EerBvjnDKIU/N94xTv8uPsT57BlMwVf/r8Clf32+gS6AuZTqPhd2E6Q6bu9/2zKz
xryaIZqa59zSVLOzJkSWtEflIioF1VFJm52ngMChy0D+vLZoKXIC4JIqoiCsJ5Br
vMXGTQirj6czoC6lzdQwt9Q2Z9bnbBtRJK5XLwRSxtPnlrHNCrIFAbppucW5Kqwe
KQB4Z4YuLWknZwYiQmkf5HcKXu7UiFy7LCJcObadgiPOoUwWVX3GtrnuGLyjIAR4
kByfkTBVqAe9yO7hABl2USyLzCTgin6DwB+Wlg26id7ZXYOW2FbIdDaV+olcto5q
yzhO98EmK0pKd603UIW7+W1e6KWp00+di+lNBCaea4t2QS0ofTmXUWMTJiMqrd8W
NSMBXMVwy8SQ10ztoe30jDPl15RVe9T31gDjrnmRr/5vwG6a2MS7NSB+XL4OAvtR
tWD8JlgjVPn8PCC1pNouz7dErIN2SKOK5ViUXb2i17AnYhOjRz3VCB+NWuCPh0im
nHV1imY8TziynEwmp26vGg8w++CvXu6vjKvE2XISZhVEtbvj+RFbi9SKXEqA33hS
U37TdAAosZPP/2x5oUt9p3ZXVjM0FkweEMJfOubXL/Sqqm0Gi+4Tfpra8Jz9IgSq
rR4xPKCIheO1sxhWWtr4rv6a9ZxiFA7dwwrmuwIhb6f6zJ/lhEkPpPqpfecCpMhf
a27yhRsRYaSl+fHnR98kvspBWYsfQiaWeoS6EyD66uUz9H33rxTTa/vx35IDCcFn
fj6hpE1alPvlwHpbfRXn5w==
`protect END_PROTECTED
