`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YsZfepMZu73YCeSBMd1e5nGdEYIsLuZiF4gWInXqttJUX53FHnQKKH4U5TJAfmjo
ZqVMZ2Y+5qRar5U4xDs+L+4VjezEg1/C5nKfrvX6BepFjNmBeWGYEvTMOo9ag06/
cXN9smAgTVcxCf1cqJmVmFuWbFYEohGCPwG6dn4MRPvCtu83XqZ07gf4dPyP4anv
sPoJNA55D8w7bAtpDFhMvnGDeJ/dAyETgFaAZcvRYIUepViyiZdyV3ulGjgH/w2c
rTTNaR9idQCn4UJtCwK0Ti5icXAnNh54TAR4UiV0R5Q8i3uny80ZkKZaglGGHI9U
te7psdwojAoC/cXdEalMtGBrCPY0bTkbs4PRk8pnabFB4vX/drgST1rslmnXbANj
mW+pGJWG7YKHptiAni+ecmHVcDpHnQCCWYEfJ1sduEw7xRw62MWnLPWtxxffwuES
Cx8XXNCBeDp20Ycs2T14taj5VWTRYDm+ips9iwi8i5Bwr+CyHWmze3+vmjJrTRom
Trb5azcwRTB7abhp1QFdGl/os2oiDxhixlKGniaQU6u40WhhMTYlVFnB+ia5rREL
DtdjSP8uQyQ5OXYCFIPO3/zKLOShXsc+BCo3qDgl/tkX0kp9aOy8/m3TALok7JPz
FThkwJm+nGYeKzIGIfZ7ZF0sXh130iB+ZMBVWUVVt1UUA+5JbvFtd/oUed4zBcaE
nqY9wpjE7ur33NB50H0L1nIop28YwYRmEfrOUcyJ0NONpHHB7nkL8/dEGOwhFBRE
EkxytigTHgiCN1yc05bRqS2tgG7SPzbyqfgaHzdcVXkwkobjjF8azDv2M70DlJj5
53h1Ismsl5H3h4INO9H3YryOLycHbNq1YNDOUEWVeU/gD6ED7wSgJ1B0v/6sOmfI
8MSYh+pxir4Fwre+fKi8DP2o5upZBqlt+qN2/60qZPSNXX1knvMBLZ6KybYVTJNU
iQgBAshgxAIlKO3+a7l7gkoZQUC+tyrQ1N5XDrHmri1NXdWRHljteWQdEJXAmh3a
Yh7qbXtggOccc/BR86PlIof8hOW8q2pkjKGkMIdmn2asIfX8K6FIKeN8MZO0P+nm
Sly03YRK0ZG6fu0caheeU+qRyzZPzkPaNd/NEYvmoNXK7uzvBSE4zpciWtUndOkN
S9bCLSFJfyOuyKnEf+aUcnBDA9pU1KOJ4UQBaChodbtI4jms50/RXa70UcOnYvM6
bUKcxY5RHYz5mHs7triQVh499psfMhfdFfzU/kj9ExUdF1rpbjLjg/Ix6aVWYyEl
qWSXDOnLahwR8z8ITL21mG4RGMRg44L9khsrLPqSDq9wa0xr3iF1r89Q4m5XBfw9
UuXSEUx+JfPBWlR9FG0H/OWfavSVl5krzwrPPai9MqaA+CYVJcc18NUBfRwqdy2P
t0h2wxvzQAf9JBwyPjypzsACyWOQnBb8igpAPKDUnnxSCSo1v/bi6ayIn9hEqxOL
ZqkTbwyWu7Pgt4felZm0EnyTFZok+ViOaWVhZ17MlDGVPgMmtTZUsIIm2eUdGz2z
t0t4Mxu7kV2cQAnnwqaqC9078NQ6j7exHoftoUDmCDTiuefkKdgzqG13CakGKoAx
jDpetkiNXt2LHWpDdCIvTJfVbu1e1UmmoY/90h5wiAMMsxVlB8nWjy0Xo51dRBh0
gX3+l9sW5P13fLDxBYryMo2oMuwuLZqYbuhY+psT4ri/GDc238jgaGqeMxETNcF0
x2kVjg9jsafsUZCW5du2j+/uq2g/TnCdqL+LlnXBeEdU8/Ziqzy7a4qYils3uvaY
OK1kzXS/oPOfgKcZ4rXsvtaRD1DCSXhN9Y38fD7UI7yLU6dXicM0Uckh8HUXsoNX
ummbYGJ8gKrgSwB7THziNZtztAoIUGQapILo7u1au4gkRjmVZmyi3deeA2NDPtBk
UbcyU2u/gHwg/+gUfsR/gxrO2bqbXyAUeRlix7fE04lW+HTrBg8h43NO48X7/xAz
+VLomocvgDZBZ9Cg8ageOOMsAGOmg9rmUxSNQTRmYt+jQlsSKGI9QmmlBZOJNIyq
25XCLfIyClu/alI4YTyYYLGmStnuUMC58Uz22s8+96QC8CaVIM7WZ3mlVfzbtSDn
iflwgkVURXbQ1An+ldBMZ/Hmm98qTHgiW2NbDT4KIt4hW6XzStwTzbQ0b4vEkLQw
/GZUkCl4RzeJN/RfX0m0tEUMcWOTJ5H8NgnbK9EBzQ3tz7Rkzu4TXPfvtNx5/UhE
78B2PiPTBPeH+q+f97sJkJKpsJZ5D65l2sMeVn7wbgHwEa4YsuJwGxNhZvuG1f9W
p5mI6g31MrHRwUCAl4kQOlj4XlzS9XWvU+/1/4a9EWdXurVbbiuKgKutSGY/nBkh
9aefAHIt9xq1saX2jwf7KwLwQtT74VXYior1lt8HTP5dl0P/vdV+UmLlrbb/0Uh1
zJv0KPacVpUFPI9aDA60o8pTdqas0SoE4d/ZUo71onFk7+WXq0xome4mxd4qnbG1
IVBnqIr+cG+/nhedzO22xGQYG4O4SoEjEefOBGy38UzwtUdZS1kUJ+tVrpK0ZWxi
KGD+UouqaEevI0k/icgwq+pLFrEdvPQjT3YcyqntJiJgmX78tprur+2a4tQ5bKLk
HqhxuJBKPZ1IU3tfm2w6+E963t7xv1zQlyZTZfJ8C9w4lhpw1SNryXRdxTx4S1Ci
xNORlsE4w5QKfD/bYt1T72A7qDe2bERW8V/OH0pWIPq7JR2eWQlTUV4ugfOCMBJ5
JljThs4lyMoM5bOIbSYV2vF15uxje8rK5iv6NgTJf7fidBoTF34I6gd8jJiwz4j5
kduTDjzzmQjVCeR30u15yPy6L/JND9Cs/gmSoPjAlOsPGkAKBzRI0+wWvDtCF9tf
bu0jaPYiWqNXAglGJvTW0wlm3YqO854VTeRqLxWi+VaOo+DY0vHjhkxo0F/83xBc
hJIgitiDA9Kx+hGcPTGtFR2FCDhnQ9T5D1CnnebiBQ6+rCzQVeJck/RH/eGtHA5v
0oAqRuOpPs+MQ7SeFptx4njgGF4OrCTt1ueEaY+87DLuSUAKNXnFzj18lp0uS4DM
tvgiB3C6q3zNf00f5vST89vBNUuXjjhbvCyM63NgRgrCLyWRX4ZjUPyJoFNLbaJc
azX1JuU1ip5f8wSwOkn4Pobj0h8d4MlVPUxNydFI8KyWz9qECYTQknqu1E4p1swa
fadlkqC2g8YisJ3pUfzLi2fXlehPz9ynjIFJDWNbWWMa/HWRO++sduIIi1sXJpzh
sh4qdKp0BFEXGrHMn8qJJYukO9ROsJbBRVu764BBm4qFfdsnVl3pXDN7z1SbCkDq
NV00hl4z8eswxsqTNySCjZH5IR0LheLKUnlSRd1tnYIgweRaDBdhtHaTO0PKTzK2
6lgpMa6gRSLH2iwFHMm9Vw042gH5mfbILEliwtKMCjJFeGweUO+tX+8cAml5MLIg
+w1F+H7ohchrBCM8e+cETK9+4r14+fPgU/qpmtEIu+oyFApDLHdffZUy3a7i2kJ/
5bUqH/RZLNk+DW4peoow4aRoqGD12iBuheyHiOCiS3NNTmr6YcrlGj6a8kwOrN/H
46UqIAbZ0rwTGZMXHHlhmOtOYloF6OV/ZiMal21OIWDiPa6uD4sR87736diRBUWp
I5VMLU7S/2J/tXtX88B76Hnb0N3AvVS0sVvJKIae59PU9TVp3BVcPoJgg5LRkoG8
D1pnOZQi6AgSUsX4zdfG6nflO5GLgpiZqiT12ywBio/x1cjl8N2Ubqc7fInSDS9W
Xu3jswncM66imEYyC+SpEHX/ZKVY7CzLp/FTP+MQIBmx7MwPCKx2iE9zm18fwYlV
LghIe0QW7ZDf5Me91Fh1vuhZ5kDDKDJs8rA68cDQtdWE+JPLCMvWoy6IynQyjvsb
FigUDSWJlpG2DRCUq/K+jpuCOeoUgviHph8jiszmh1Zi6WmwaxpWoIraO67OHwIe
UJnChaXhJ0hJQfiKO3sohlNxBWFMtfr9qCM1dRyQoEjBPzp1mHXsAIpKazHS9akE
XZINt2zxMGwpkdJrGTQuwCyIGcfUfeFOsHMb5JAzcmcxqScsZsitgybjTUJdMVvW
VaxD3q7tPdJqREDKzhyep/6KsySJdtQp+HB2EFRZqVrlpwrhtnuRyO0nz4JwdljB
XK1wE4AIvagvN9btaKDvZU57dqgA0EhDV8d0/nI2j6OenICcsZMtNCkal5oAruTF
ulyIYQO6l1coJet6Xg5QyGwndCCRVQCEXSE8FNj7gMVp01b2rV4x34HNXSBDOvYZ
k5yk64jJKxxVa459Uh+lz128+T3X+dJvPlv57mEeUE+MjftCM2b63cINfIMaiNYG
gdRsPoytcmjpr7eyUs5XNJS6Umnq4vgVmtQQUIxD0AHT68Q24EFECj8dmas6GnyH
LOmmeTN3Kbf1Wg99Wt4cx325xQCHEq6dyxziXZcnoSFTncaJOVHsNYDSBjJYgE+K
xG+Got2JELusscSVmC/Qs/Wv4KKhwK16j3qPYCyYNix8LI+EbzHYfeogwYkgFmNZ
zDag3XLz3ctuEIOYyDlgL7KTPKlAji7lLfKeMWMJniP9LkV+JeA3Ma+MHf/d9GJr
z+fL22HV3VIf/eBkF3o/n2d27ZnmCPMemriJ6YVW/MP4FChnf8t+me087X6yz6lk
0IDnnoRlCQQ13pKhHU+sLMcxaZpt3S3bw/IN2j+Nzz6TY3N6gf8gRxfN58+qkh4/
Mb3uHE7X9WgNiBWCINNng3RW8/QU/TCMuGJ6rAv36to=
`protect END_PROTECTED
