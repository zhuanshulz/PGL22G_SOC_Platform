`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sUSl/zl+ECXNBCzXpbOJ0jiz8l53EJrKGyqNSAbv8sTp+zm+2EQ1vKxvTcsAPseQ
FmP6y08t6rlu66epMMOJdkE5wVqmDQ/q2bqbymMPgx7x3FevdvAEQI6RbsLWWTVY
cFT9jvS4b4q6GWDfWB+P2KJMvAU3l6rzV8d11CWchguMA4Eqsyky+1UtAJdYVOGe
Cx/rXwYXySddAmkqYPusLZSPWDpFqDeAu4+0we9v8B5fqhCtUq+dm3X/b2HjT0h0
m7rXwtLzwd3b/oySviml2vkmaqHc05feM+8eYA1DhnOnJqQaDx6Ho2iqzjuV0zhA
BvOuO/Sq4eY8kJ2gMO4JWrAv0leVMMmc8/KWLrVpMkXX7MgApqd0Rp4nlS+giiLM
Mz3cBjspa6G1OMiQJyTH5A==
`protect END_PROTECTED
