`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QCzWYUxfuENfInZcRkDevAdHszYjezKdy7G6fSocwPJzQXk0fJvTOZmAeCA3w4o7
v5qyOA2ZMLr9Hegvz9hJScXhsUPb/xXj++NL2znLcf0d73KeaFGlfi8Ual3W7S6y
1PE7cea6d1bQK2HQ2eqDUEfbN6c5HjGedpxqVldZQCISotFy8zU1nczcC94qCpai
gnkufmwRPDHh3onjyD+eOBEPepy5LIWiJjOqXKZp9giC+CmuO2+p0NFMB3wNSF4t
b0C25UfXUq13DP6yqo1PFd09Vmi0IohLVxsLihkoGuVHNdQJ+CQwSplrJqko/nzK
pxoDNXSPOSAl3mwi/AiYIL8rGvKgfuyDEy67i3ftzOp4/xlHzVyg97LpcJ+u09uh
jk/ekjWUjaj0PDxRd5iri/30E2S3bMW7uzoEcaRn0KV0bU3vBi9XnpUJeWsq5xKn
l/jnn3Ny85zmAKtatHEr96fSKvHqLNmbp77TU3VQiNgjXDn6sap/PIHYXhlQWbvF
yTJYd3QfNxnPAOEMW3JCzV4XbM6KByawWlr+xEMkXJuHPKSW1+V/LG1uxMRpt24H
q3Nfl8TTDhlG2pDPWgT55FW32VHgCBOOpMLN5xfaiARCFluKaHEOiU62IyA+x5PU
Qh24PGfGuJVfCN0I1/pIISwG5jLg2q79HKEsu25Xae4aek+fyALSbnJvx+y+Ei+R
0pxQlZPk1rBO1Igls4v8JSafZ3fXuNdqebYD7Vv3g6gAlB2uWKIvAImhfUxymPdy
s9BJvqj+JLdq3G8tAbbCOnj30ICxDvPJ5hZ3u5x8rnKCDTzUXl15vCOlfYf5Wfnq
S1ccZnntTA9ufU4YgjsphHaa1rJ6GK+gTGQwvYJtgClGhjzZahncprTB8mkdg8CM
f1BZD5LQt3iE7dm+Wx64qS0KSmijPHjQx1LvNt7WT9WXtySOJ8pXNuc5dRhrs7DZ
oTPyFyY2dtturMClNBtsA5SYzEOU6+o9nfov5yESxNLSpwr4VFkAOoIyRkqLa95G
jv7TTmRD5OTV2OsLADWdJY5h6biuL6llAyLZsbqQhjXzLiVDeF31vg394z0zAJDG
m1+FvNfMjAlN9ZISjzDq7McJ9aSfPcuF8wnbvIB3wwABobKFm/DFgHczv4YiZVlP
hDsUUjoSVZnQ69QO03qJBjXioOWJzMNIoYzmauYKury3/Cd4X+IxIHvsM1JSDoHz
JfP/RV1m9spS1cKFMxOiDmqGh32WWBcih2cCJlk9t2d2+09g0MQDOiyuFN1WGulK
5FkmusrnWBRr4qi66qbtmZD1yuKG8X3qEg8HoHNWLJ2rl9SBMY5V+6SeNODVXC+e
eLiVBmVBWxHfmYmy+Hv04C7EoFtWfzmjgWXhQLXPxj2UoVYERsEvzSbs270fZkbM
DAEUeZ7E6cNe06ADlbGOt3ilNXd0WrT3ER4S/NEvxueGV2DCLwjEfUMAdcTbisH8
bYB/gWtG0MsOrZrBNbChXN68ELl0xBnQLq95MA8+SRWgSai1NzvJ/KDigw/7BIog
0M5QpqAmQS5d92nn+rspnppUqZHJpwMb2i6yi7cX4Zankx4Qbs+wGll7TRcx5ZJk
sTqlO4VhtL/UivPePn+E3U7PzdgUAPEfcKM5COL1zMhWJSThe2D/CmzN0sisHRDA
LWsrYXsjV7G7lE2Iq54nYcog4P51pc6/zFJXXACCcubDOxTei9lQA3tWCFThvYwH
yyw5lozsaICG/A4pfYknWvq3wV9UEm68is/zYaRcgWCt1sB/PpuSmK5cihv0Fxtd
Jb7bzHglqD7v9jJuhD5PUkhRn+qw8cxYy8VtnAQeR0apbr74WvD05KAFcEYaPlXB
wR8UnzeeA2316WPFPx9TOpFHJE0kFax8KwMP+Foc8NhxJaXH9wbVbkB7yvhC0Q+i
e4J5kMGpjQbT12NkPVgGV0G3JztAkCJQOVBtJRmm0RkHM+mjYqas58Zrs/r/ZT1C
GP/DegiMhoMm/NrhpV0Lj7x99RQqGQIHEav1DgWR7a4t6CFSQ9seSWajKC6Sd2E4
qC1YrhxCM/R4/TSBie6HNK96KsKYIfAOJtDFGU2VdL/gNc9acsUJVPRSq96oNkaB
3DAEGkcQtl6H/fms2NgRU7rXWqyaXbzDAdHJssoP2C2bNBHc4ukK9EbzoUYf95SN
sju0vzeH9O2LAdFKOKLggP75Fs1MH06HsuH+NkI3rMhVqITTGgsCcljn8Tn8D5N7
YYEe7c+Dh+XSqpwg6ooYr6MpoZL3W/aCIiTkipNzJZzf7GAtNjOI2WADMNueRsst
4uDSclGrKB2t4u3lpKZokLJIKteULS5qfO7SHaGiZr8tDtSkw54eLaM7u5rCv4uv
ywS28SkXd+erDXRRQT/n1wIPQQmAyF7RvcWzm1AExmMm65yiO1FqiUnX2GKehy/9
YVMYSx9CdHQJswcz9tbwE+rMIKTuT4FSN/bNy5cYEKYT71L2lvCqsLHEr1z0tX3o
zik/o/yc88krlqLh3wmn3lRR7WdqeYBcqDDLLhXYvX3IewMwTSEG0TUXVQ/ccf0V
oZCOZdtL7nssBgWSjwEe/6fUdJU5kMtef5atgcTgrNKWFpgxWrK+8YPjxb82z1OY
ivEg3hYfh7HUpbbuFHPlwEEwXqWFF7MRuhzXLwNDvWnbQaomQ4khThYN2yiYGBMl
PJHlDm9hZzhabJtsURA0PIAcx69cmTfaZL+XJrPruQa2OQ4E8As0ZGKA/im6fVEc
7Y6pPhThWViixge3cp+T/6Jb1cHparlWFhCXsgV8OCT5VVrBPdE7xn7VFztkMC75
2qn6M6qaY1SayoymsXYiSDyWspWJHgG/0inDuOaiMYb8Fd0MBI20Ylo7p61CK65x
QCrgt+RBLq2dRpj3zqLfd1jU3lZTBPcSJPRWGoGqvm8IRt6TuIzKEaChLgaAMEIf
y9ouj1STr18x1mGXw+LNNW43k41OTprFAd3Fn6vfCbQCw5fJdxzZiOv7bqEyqwUc
jBJoVMpA6/lOf9ZqSAEHnkR6NvSyNrbsw1yiEfL2+CNNODi/j0nnjs3B9/3OQeyE
O6Vp+eFIXFOgRYhyKZmymO+d96ISmBIDe3EkMYrsIk0=
`protect END_PROTECTED
