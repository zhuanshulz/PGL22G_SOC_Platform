`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ztbd0REiTVeEzT0GqO92UPr3inEkpJLl0EEjdyBwK6ggiBJ37xPcVyofP9bZKlLI
W3TDrkMeZIc5Dc/vIzMpDEeAuAbQnVbiwugHYs3IqAtzSUWRgZ02MpSCFmPWXxmY
vLXN1PDFsR9T2XyAofC7ymtBaZD7w5KGmouHXhwh8sMpQVAqa4flSMee8KkmILSs
2bNhChZc3tb9daNx1v840XeAsFrNwj34vwHICfAMNJeIUMcrh5BJkPwD6J63c7PZ
ahDH6JHWlC82d+5YLixWWBu/Fw/bl08HfjG5XTRzzIiT9OR8+VWt9SbQzC5MHTLL
jhhY5iZlEyKkfOPEMQUE05qnulHpnJ/msQIU9C1Rk63S6zBqF+TxfMg4FAikcNF8
KkubgJLePFsTqHJTkAyNjIJpqITQLhQ3rghmnp3bo2kqdPT++2UXzXAvT+XO/WOu
B5JqUJlVxMCo9KO92bTVx8xAi5nBD25ViJ+bjfCjnNf/gIJKG6FUy+Jhp1W07sVS
IB87M3wdhF/UATrKJkd0Lu405VJgdPYs8sXmFPhB64aEHOTwik3yfZ0xxHkxFQff
ks+GD++V+Qlo5uq+W3x3vRICl3AgqLy7Qm3NB49m46SeeDgg917ySyF6OaezWdlv
5PMw8JIvB0m0+FyZfYW6ZnGuMJ5tIl8Tt8WJbIfTNF+cpafDMXZaI5aEsTgI86C+
8q+JSRdbg++Lwp+v4EXkBSe9rP5MF+y7gL4rdfRWExfjQw8Y20p41QUNA8sltVr+
yaYWxNuAeF92G38rJnv3CxSBfprCoku80oAdlvP1ttE76RewH0d2bIJcd/gK3/tM
v0rEe2P2q+YHm/bmndVhIyy6vPh8XvpMpEbP8nA+m7wWJAQ09JkRoOyH4CUkHy3I
Q+KZ4Q3G/UuNiDHQbH0mGYYL1W7YHIatdvjOqSwOS5LHFbaZQLqVPOs4ChAeoUDP
+HDY/LY8Y1OtNCfPRecBWD20mLfOrFT6Gyd8BlJ3W3vZF0h38V4Y4hzftnRj6Dee
IR8LCZxvd82nULCSxETIWleVk1mdwj6bIX9Eyj4080p9QeRNsX5N8EvAsOGZrsrM
hF5LT4Q8fjndED83Yt6p0npe3PZIwcL57gvrXwl4yEieUy5x/G3QKxyMVW/6lcqf
Z+sC4uAvEYVGe6ljyZYh8fTna/Hg6qeIN5x+5w6t6dFSjaVJM7fcH6v5CndW8xJi
xRZ9nBH3XFeuqs+CsyKxQy/3a0LlGXG9+NU180wSJw64xbfZioBlDK2i0KSNIABd
TGcJiNAF3xtI1amgwnN3j7HRPNN0kRjjMXMzTUnaI0baqpwXuIh4uWU9y5wQb1gL
J0IDj/Y9BBpCwg+zbau3vlvmWms7FeGebYw15+XUM1IsrWjOva2FmDTLUrAfSwH1
C8uoS/I9ta8n1osQUkuGS3+/OQVfULEcKVpHm3v0VVRvHRmN4WFH3JKH6oY/rIgX
M+HxBt20mwefoxGLTJTPli1TXEvidrRYxxAN3HiJfItRv0eKQbITKxMxeOm1RrV0
mjBdLcDu2Fr7Od9R076yrG66+tGyymArMYI0nRp1KRjq9EIudiqeEDMqL5fCGNnn
MbuGzB32bF9GeTZbeMSIjuOsUjplbldAfWeINdrhmbZtfRnFkCWxLHupYqPHnTz4
94vKfixylHc9b/92Ft87mfVoKU6IJ5P88ZvRKLamiBh6aNbsguIypWbPDP8pxmiY
VPWPBS+p4fxZIC9cFx8vz5hCXalLr+mFoKV4zI2QMHC2LCGUW48AK/ofD25gIJc7
ImubbEVH19hhrwkMGDoETS8ZZkmyXEKVF0pV8T5zTPD0IlBtmsDHcaYD0Q4xilfb
ZztwvOmm5v2s0QUTSdnX+qft603ajGaAF9SVYGksewACvHkhso2tBkW+EaiDNoDN
EMlE+LUrLb2rSIcGdodTB/K4no7Swj3XcM7AbWk575O+QAGhRNnkBSmyQYmJSBFr
59Rfi50sAfjiSSABy7LyelSwqvdUh0M7U5WqogLAFL7O8Sqv/JADiq2SyD81kKkY
ferccKXsDrVlVD//6OMn7wCvmHlVqJlaOTq4cX5nWor2k+jzmoP41PBFHJQ3UxVW
mwY57exfPFyndTS3QCgxEuRAfmrauBVzkanc9vej8bByMv56Leyzjs3Qa5Odr8+a
ICJBbGw/flxmpdtMZWxhBPB2/hVWYiN1hesSWfJx1kKgwRZmXQFWDwO9/tABrMnE
bRRyX54H4/MkVQcV09gYn5twOcxHtS7WPX30cJYS+ckxwXsLY3MVL7MaNp/igvdu
sRvTyo5QAPwL6bmO0U7SxysZn9ulSFsa5K2IkVGL6/3eReJ/dEo6GZASrxwDNWkM
ha/f73eF+2GXZ5mfQ462dDL8wwHwZaCL0IKRHM0UFdG2K/x9/FRUAACiOzdrj5pQ
etX/6LIVP3wYvuUTecOi+ue2DnZN4HffJfEp2SBMt8NoouXBdv+9w0HtQbhalqXj
W9aI0Bf9UYfgGmvV1lBhlqHoyxKJ40FhOGZqJA8R7Q8oBLFZ1ue4dzQ9d79WsbFe
1J2F+CxRiUC82TPRXn3jlDJStf6K2FnPV7oXUz/j2NzaPKEHO8YxIeWV8dP36vsV
jHbo5KLNCX4qRJXsKvTAIMlh29xjajBxXIbvlIdmlow8lJtL77WjJvhOW/75q7m+
RICD2jpsGRaMLQoJqTIJ+gQWsO73lUNNHlNcS7/6Vqe/V3ONhBR/lJB5teJl312t
EPCNZKsmSMUVHBLk+nYiGwhEOfclKdUPLB/6Ke2X6Y3QcsdJGKdD7xPfutVHHYoe
wEyBs38/3gsA/D8thy8/jfY2CsI8EACQ+FNQGZ7yUpm46mB7lpyAI99C5scdX5Tq
dzUsCBB2J19ZtBxuoy9u0kfLIKsfOoMWKQNVuEhrOa+wUNDTNKqaVtbR43EpoDfs
7sOg7mXhVsc+We59LesxGEBRpPnlUhB9Snwl6I98TTIBujOvnYKSYxUbvxC8w9xH
paUpSA9rQTXQ+QNzKPb3w7DxebRBFZS3IXtEWDWbSB0foI8tAro0UkVecVagu8nG
HI1cWGQ+4Ab+c8ETFYmXBW8fvqS34On/D0edxSGi8T+RY9ZgY+hjy2k4CJNGQRKS
s6etAbhcTp5AGoh5hd82pyt3muHnzJYTLh7vKw8IO6WCs8wW7N2qOXCJa9aolCOn
`protect END_PROTECTED
