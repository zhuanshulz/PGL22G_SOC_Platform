`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NQ34uKrHKG4+TC+5LcDwOKY1dtxhFZKozNFOHIAO2ZgGeq8LGJvVBVZUORl0McNV
v/Qasr6xijG9Aezm8qroEaziEkoQV5rxIP76ytbjlT9FujoAejkDsvZn+ZWJMFIK
T1w/tXZfAGFziYyJS2ABT+/UZnI4/F/Mv0BssdPje0jOys4cWzBjtp4YwTOKXTsW
qlk5AczrwTqVSYkE0nZgjYR5BUhBYzrA8Gjy3Ac8FrGcgkdBIOztnMFISo/3ZVVd
A0FAR8bI0M4t3BKCKbkb64NM2JurxHFKbUNSUMpa4V0gRJROf4EJN/Bzc/aVdUpZ
RYQ2YLAVxVguHHdh8We8olFFYU1z2/PCNcQmQ0o+XjcNMuwzcM6jvyz0VYT55m41
V3YVNYgsfG2v46YlfSLROK1HuSRZtjf1qZJp7XKXrFwYuhpeD1ccooaRPyGetmsp
tzg2A2weQ9KM9Liv8tkY7yRmv5U5gFYLGbTBQF5BILubeQTpp0mbiL0EjJrH2WI3
ZQQ8DMI23UEGtvdN3wrS0tuMnB1tm+4ZBMtcd4J0zyY=
`protect END_PROTECTED
