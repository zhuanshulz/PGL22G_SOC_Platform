`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UcKEu9GjXxW6nQvAjaUcgfulujFGjorGXWFq/twzvWzMZabF2rYYicvKhQv0YaZQ
jh5WM9gKILApP88fsfLtDRJ4a+fJSHxsJ1PHRUtGfyTWLk99YHwpExpSvF/cW7F+
VMnhrqMqN/T7tKcmwj/n0MP3D1D2XwG5Kb57+Hp60BEtYu2w5qWsumLDnSGlxMoo
Dz1wCPGBbrw5CShXNuY70BteTT8wIOOaBpcvWJivcLeZITl3COTK/hcO+Yzp81Sq
zK+J/XD6U0ngovpmCTX6+pvCkO8j3n3y0/4o5E2L0UBlKgo60RFt0nDKfiMVkunz
ZPgymL11+xa8aTnFMRvSr46lp1YMMVfM5HHzgLhnAtRyyTQaQyxQ/DQeIpHULIbZ
x6I6BT7iWT9bBidaTHNkNPxKtg5D3xkeLBMdI28NI8MCGG+qHDUmdt9DDI1KmEy2
4G54Pu189iVxBs4WzUuFgX+fwKamam3+CertvjDLyW9xzyVqIwjABA2W8dnJ4k9r
WFIN7IU20FWHQLNZ0F41MnUG5yfaPgcHszZAv37EEOuG5XhFMhleqzkyYTl2gnkM
3tX9pUxsRRSE5Zigq4nUZA==
`protect END_PROTECTED
