`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+alvb4SnDuFBcFamn0NQJDDV00D9q105MOZjleIY/rCOnQR7C4c90s7XVPEIl+QR
JqxkQ3Q8JeRzBwXh9Wz5W5H39IK88CQxDFlWGurOHivGTgNVQwdV9WyHRPH1eMJ0
6//J57uCVOIoB7xBAMfdRwXKRp0/uUQMzrMmbMbxdBq8Q0sh1wFItZYDq0bUfPtL
OJ99h4BhGCol/vopmjyTb1QSwGqfyQrF/oNVl5VhR0DPC2vZSjbwy7Emzg1TbYq+
0LOHi3XGhowDAK5ktZ0Zl0M/QHisfOmEulukjPWzvdVvDeGrETxY77/r6C58rw3K
7Pwf8YfJshx/6r3dzMbsv4Ics9WWdUmkaAhoBvQFpw5Ihrk6uuNFriCfgVa4i/uX
zWOsYSya9X9sc9Pu6/4hE8p/Fnqz9BxXRkdilWr1qB1OKQFs+Fw0Ja3mtOzjtHyK
QIC/KjUq1r0d6PEafaa9Xy2nYatcPk8hzyvLRF6rQu8myFFDy8gW56ZfHB8dE6gi
SJL6C5zEoQwOM9TFUc2iamyzEZbLTyHoVterVeKtzEpf6gC/+RHLIvd/WFxL3ibG
P3Fq7Z8o+BNRIQiPbFaGpxZZ3CoRV0Y1CyBGFk//c5omOmtJ1mFPqdccZkkX8Tac
`protect END_PROTECTED
