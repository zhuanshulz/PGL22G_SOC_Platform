`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tHmSvmqsRtnGmQcq63vmf27YTmog058bIqMkk8jz+V4k7UtkF1pbWDGYGedtK52U
QzlECKxqKDpvN/8yrAvU+UW9bzSFsHgNO/PuotWyCtdohAKu5CqqmWa+tMtaVdcq
cJbwEB63ouFoblHgGWCqqUI5f7RkcnTXTfLaxWAytX8PbFJ2TZxNCx7jAG5jCv2b
UHn9JkMLa/1tF3SaT+OuefDKcC3F2me/GRP30ewL5S4OJgUb5DvIn6N8cifIrMaM
ySKiADzMMI0NtLJJqIDGugDkNvEkFbJxdzTIhjCYXqrSoSGKl3z+oOrRo70jki7T
ROipwrsQboQy01HKMUkBzCV0Mavz9eTgJZnKptnHV6Xb1cMsjRWIW+4sXfYM0L5G
WzqZoi5PgF+Clh/bhd9Ds9GF15HlolbcCwr3vo+xFvXf6Hw6KeJKaQEkbJudvDpE
75qN3ksbXMjRAmrLTRQlLQiWsozNq8jjNPebSmiC69nEVIqiJQW1Zil+ixPywQMe
J3aa2hToX4JYFq6nq7WKbH8meMbJRoHB/bmv7BzLpc4EfZGN0S70Ss/tRRFv+45H
oVAUDco5dKof6sIihUqFlYTJujDihizGzspvZhIaHjg2RwOG2K7PyIZoeqGoHSr+
aKVOAsgTFFVIcpU9wAMfuHkBJL7VL7lKVw7Ud9YWL14jjmdY0bQc3mQ1PA2BQXQX
wQT2TUqYtKpKMeIqx+2S4oLRUM7bKi1bFTO8BI05Otn6LXJ6A7iys7kJDldGnsqu
EJIajzi7PECJ3LhvoAoUvXTumoXmjLNv8rU2mxg5JrUDRqcIqhBe847aUBQ+NSDn
UQv5XK4SUrVZsfN0lfAw5yCiwnbSS4aAvsfB+BThtpJELSv68mR3DuIRE9gLueng
`protect END_PROTECTED
