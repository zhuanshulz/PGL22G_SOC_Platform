`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
50zYJjJMq46oGwAHa2cGZKCfZooSQ1U5or5kxHt8dXb3wP+vEgVF/jE0M4vjy1Xm
H3wc8KhtgHQo4oQhjSY+UrQqeN704VfgFL0XRizChZVxtnHoKWEY84bBjwUMkJIt
JNF4DPZCXu31PbrjukgCbY0wWrfDlZ7rAwnLS1hhRWuqmtIApRwWQcpnhGwGLgV7
eaYW2pa41BTAC7J0P31SBy1BGK3yf1Hs0BDOTwDHve9BVfUFOaGPPYFSEdm+Fcb0
fugDGkGGUY4pdWTRNQOm4gldRoUTfG5UWMx90DZg2nHND4wdr1l2GAMGyndaCmUL
2jeV1Vr9X/kQIoj4oOCx79LUdWQ7ULvG0WOirOxon1Mkqn6CDalMUFREGwT7FCaN
58VS2mFxVy0XdbBr3eTBHTmZOdyWgLHuWvoJC2E+zOaMHlxtJlIM63niBgKhix64
ZRpluf4gONl3zJaCzkMTtG2VBwi2yDNQCzs7YhSx4NFiLkLgq+EW5OJujZ4nwLwe
Zee4LuM0WbP+ryGpX1oPPhMtu2+WLReYwP9lQ9+dqKvSP7v+hpUvFM9/5VToq45e
yk8Jq0AMdtQ7O5NO2wYUzXdkEKEc9RhHuWbb7k8f+Y4AzaVw0/eIM2kmy/L8/JOx
uV0UEyqa8AKNSkSULY4GfDEfTYaacaZDomTvh+aP+GfhlT+O1QgkGCnQtN/6ywgh
eBRY56mIxiPXochpOqU9J+2dxhiQf0FcyYSgCB5tX/dFUGOsDPCBJ4pYaAXGNl+O
J/Y0Qaw3aSEum4cD+f/oluLNdWXyYvTctWkJAaHeVqUE15a+IEpjk/FezK5cdsJ2
mU7qJSYUQPpqH2IkLn7mXW++aYyJI4CQom4aMZDQChnJQbuwhwTgYlycVPqJ8XIe
XQiHdoxnGQNhi1htEGD/OPwq/eK84wEbYjwmsSUDudreXGR6XQl7SmO4+nVk1vg/
Bct96sVdewdsBKtlNxdfdedsKQhgvNyVinJYkWGTSyqzPBofSxFxralEnZk14qZp
bXjR/LmXlYEH58SS9+3VXXz4RcZZZoO/tUVyafp9NU73dc8EEwsXDURH5bBqyZ/j
SDgcScnC5xH83QUDBf/3DJH1OyPV9p/DzvMufh0Jjs9yvgVcGHZf/ffGrHfmpyDA
fCs6rqO+XRCetmOChA3iGUJa/CP9+5jnww2Atpgw4V7GNOufzzr8bf/L5fGDuO15
Se5/Ev1lu6lKtB01rPfTHxG5a53iyxz3fhTPegQJO/HEOMI1GyaLD8UNYZIs0R/Y
G5ljx0fpoDtE53HqaUD3qvSnTQEBrmaMBA2H0sP2e5qz2jHRz9THB7nVddKFWvpH
KY00ypt/ufpMu/Aae1vRpiSIgCOiNj9k8uGs8zZQegi6NRfX3yJcJaQxjsa3N9o4
LnEASvvEKvhyNjBsEC/9qLm+03jRygmXJWMUTMsTtz1YHv1bMXEglGCgehCtkDNM
fBr+T3VLfwIdp3etbw2n3jV6Axu0BG6TcBZz794ez+Cm1x59xpC3CQs78FlTQn8f
KXAZLRD08y6P3rd/RObFNvgyaiMkrrixfVs+GADiQlTz8De55/n169A8Q3dto7jW
+E6CIgw4Bw2dR9JzDSC32MrgipPk/nh73Z8v7IIV9gU6jPp8Ql8C07zpkyVTmrEU
QBgTKpV9gpbya1NqVY2SBbjRTGM+4utsYQ6kvdikFu7JEsR4WtegV2rlFhvDRcJ+
7nDIJ4Mt9tqJLxcmPjCQ7msllFNULlW2Iu+b8skGlHdttpQChk7F4C3VCx0sVi0U
wIKVIX6bc3JrIGNhUIrDY4dHhtN007uAkhM+FnZcks6EB9fvpAci2syqzyeNXyPa
BIXAldebtTSAR+k/1CaQpCtWPs3Po6+nftQP09Ni7YNj3nCzoOc0rsM5drqwGPgY
df2VvIc7Y0bfO05Juc1J6ER0nFKKrVhcueyr8gJpwgRujY3nhD0dnbyzuhPi4sIb
ukjs8rN3CC1iQwYExtu0reze/y+Jg4AuWN/QWEA/iRrv1sdbuvhGt1vkxb5+wWNO
vGLjmTAspCD8O3NHSkiORx9t88azVwdn4nfBAXIQiFfTrwoFYkxtsmHOo26JOf6W
HECoXVSY91B9A6FvMdNw4blfIYvauzeJ4X/rtDPc+5zvNAS7NqY3rnq1g7ZGq1LI
MgbCbhtn1k3vTtQCXPsDRwALd1qnmzl4b/eeHpqv7ChV0bS5cAcqH/HQSe/smonW
KCbw6F/WRY+RIZBJ8WLI+LktcB9nn4c06qnZBkq9okWQ5rmSnW/LLtnkAhNrUEO/
bUsvTq56qTJ1aOpGOjwRU0h1649+dX0fNfOXAU4SlmN8ayYdk0GGiZ4jujKxCM5N
cD19YVzF/TdJ3kmz4IVdZByE7njJBMlzpUfDM3jvnkpxRyQrZ1PGwZOzMkYYwH3G
k/U4866QDamOsRiKH7F2/1NYCb6jdLckcpK1zVr5rTfLkH5OUb6gjM8X6ljaxp9M
LwCmlBZ7yfXMC2egyZQzgs23e9ahmukjGAi7PowNjxcZdiQpYk7LGMo183l5RrH1
A9+RgJ0qTLLMPdZ1XkNkOftOW5/QX6914Wm3CcG3Mm0GUiwKKu92ZflPpecj0IUL
hXIIyqERR0JbGwpzNcwyZSktSRbwh4dh9NOYUuJ2YLuDG1yb5ssEbMP1Khve0ypX
N8FxkwKT3zemMlbagg7uoUb3Uca/Qw5xN98isj8P/DoYnZCAW0GzjlVtxX86knar
9SsyWu86LEY8BZDsImKjBH6r9SW7bRFNBSlBxBMaGkYsvEhvrs7EqylzMABu7umw
OulX6ObWQdCu0nGimGurebCXA8HCWmshpdfPCO8tUuQCfBRyGQZnnhE+pxa/B//s
Dqw5ukFubJpZgLrEbGtSKlp0hJPcQJz8BNlYZYWsUMIslBeelOiVR8TPJFzFRO/H
x2hdtazGn21+3v8EPcMSlSkRZlMSFKrMBL6YBIwKYH3cTOmBmMtLCXuqG1XWFTIP
obLY8yMxCjkD5UBYfFGIv5u1K5rfVhBmUpe/vr06mzO8wB8acu5Tzr1hPJJMMPL0
ttXjpBjfeK6wTW/arAdEAKYrQZNPg3Ft1D+Cakw+kekCPEeGNetCBBcWwUqoDNx1
Rar8tmsHFl1vPHdnzib3mcHWR8RAALxF/nae91t6AueROQhIK34tINb7y8xmH9sR
6zrqeY6/01MsxsxJQejP5unTuXv4XiY74RWaH0HcPsg3pvMFmxtvkyy09Dt2qVoB
ngV98ChJzZdywpt72wxgrAE/upqu4qD4Qao/e689DvJ/CtgrrPld34SKBBwHx27n
yVI3KRA8BCEwxbmY9b4Zk7IwqRG2Wmf61KlnZzs+WZ35st3+48V45tdu4Usqo4lr
AkG2ErylnTsuGfkavPjbFYPLODdeP40sVVrBzCvovqTc8CE1vvKc4+U0PEC3GSS3
zf3jw1LNHqr6rLAykL2/+2lyXYOEJ1Q79+2d0G/ouQdTYVRsrIwrfS72HGr5ugV8
NS89hQfg2aLpzBUpC2zzBEVng26VqFw5jt9K+5LoLncKFPyjdZ+JJ51LYmdfzkaZ
1kQqnJJe4pqv+bmYlmGALlQsQ+EVgJF88y3TE2FT9mHjt8SbQHCbyDJsXEQi3Rbh
y703YAwmvkEreE0yDdP2StxDDJ+f6TxjYJqtMAm/+G7BIftHWk/Qwk6ZDhvO5IIB
GWJhPgvn0m2950mHjtjjF5XjQh1KDigUmPJ8uz5DcROMvRSWlqpax3ouMHETXPH6
yetqIBH1vzk0gfVzdr9EBY0/nrFcaRIrTZOZ98dLUkbAv5Uz5UtSHu8Dd9Jkujyt
EoXviUZ6C869XeHX3BtnfwZfQTtLYJCGfyY+9Rofafw9b8NIHMK8+4NMm62MiPX6
ct+cQXD4jCeroeYLQSamF53xnU6G3yMC7ynu1Z4sK6E=
`protect END_PROTECTED
