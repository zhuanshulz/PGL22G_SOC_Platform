`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iaIoJvdWouyzmUAyt3TuNZ3IAvd0xacV07q+4yutC8X/wEWdDB8lGYQhoV/ZHJOb
mg/PWw+jjdMqrtevBU7K1p8ZB1+x16bzLrpQR+186kamSxuCojCVnrnzTSC4fY99
3BSuOp37gAMSy0aU0jh3R7hRCM/be2/EJ50I2GVFwMQtDSXrikffmyRTAwnm0dE4
9SfR8lgMz1JbZFb9cLAlg0H9kMswT7UoDBT7zqDAcriygxVCVqvNuWeEDznwin40
xg47Fg7gcMGUr3Z4kogqU6wFziB/x3LHYemHrFbMFymuy/8lX2EDNHdRMByiB8vc
kdjg8KHH+B8CZqOJqB6va0yQC5M83YE8hjOcJD3ThDWpHMmoCsRhzEX/98jHhWIk
5bUjO9YXHyPNGVbySM35R7QBe3GmbS1vHHC7+94nb7CcDP+U7z6HjGRxMFXDQOnL
XtwIGG1+xdbKdzvIlUhbKJrYRGyoG/AEWDS2jPvzTKU8KYwZ9AgmFoKV6UWd8nlY
ELDs80mf4ekDlUr6/w0WRZrXw9yAIVGHK7c4sryE68njhZ3TfymiKyrFRPO6hN9B
6LEyDKqs3xyZzmyPvnaWVkOnPiEHqhRyI8Vb6A1Xr7ue8JxHwdtG8CUE2Y2ew7WC
IB+kN2QfIjnIwrLTsuDUHNCPYC4hyOYr+/KFd/XB9H1SqrkZPBm2wqcjc7bj3IEE
lovDcIUOXOvBT3VZoNuhg+qBl6CP3jFnKKc2maGQ+juKiVR+WyrZBWdCbEJk9o+F
ReCqDZ2+U5Bf+0A5Vz82H/SYRLaG3U2RadNCfTFy24iAdFzwqN6nJKgrSx03c3Vw
83o56+072jYztZYh/t3sxjuOuLenGtvsnUZHNV66cfvQrzMFKktsQq9/D6O7WDq9
aN24FcE8Cny0HkNCudU7peBRTkxfNMLECUcmCYiANwSxxRH3I+XIEAzXr58jYzQQ
QVEyxzmHHD1K002t0TwFdIUt0JCaUAzozzmQKwxhqaPylcXQ2f6HJ0qs4V0yj5Fy
nW+1lHQVioWy1tSMLYtHZy9WIzXo1QOnNwWckGYaDl4sNfdaExC0Qmg+4u18JkqW
Z+2G7xfGgfaOGVxdD3joAcBeR0tPq4kCV71oPV/HAbpP+uoFrk1+Jh/0T3vYBTHe
Zl26a8+4yEULeYlPKoCvhmhc9j0L+2/FDST+SxjgSFOHjCH6z+Opxyx+0llxk+Na
tkfI3mGB8vOXpUzdukHuPhrun8nc6H8cntGObcWrb9YjtAekQJMERe83oFGXHhBc
cmyXOEdzobvYuDCZZtECgY5t0aXBl1e6IpoD3uP+zREqdLA8EAztn0+Gi6It0RCZ
IitBjnxZlssyNf9OTr/dA5coSDiqJR/Lem+p/VxhdBe8pi+9NrOlrpqAhgBGT3Qp
v8M5HOyDmjnmjZMTFzgCwDgmcn+UaQTCYLqagPWk3IJOqUuCNen9Kk22YIcf0nb9
lZdLF6+jTEygaDh2eosVBXBN0pyzZTpRYfI6jfB9IyIJKcUmz1EfnznxJBkhf/by
/OEPGNehdqF20GTjgcMCxFYOpyFD9CWSIZfKf7jRRyLIzNnllJYFXUtpfTlnrBYS
AWOdlD/qVJFFb8PYGbleI77ZGlnC3xDcJqACiVU4YMLhRkcga1p61wX5D+iTBtWq
9lcRzjhb1HYyWXm4y2dY5HsUo0GbvUm34sSwLWmmhCQz6DZQjai66V0zdeMemMW3
u4bQHykXyUI1cyr/1TvCLiWTt9WgRU1gKTdVM2EjOtkKaN/2YOts2wFyPEG1/9MK
Alqj2NO5eAauhnUAbz7EXFPlhVTknt/oLn/GYqSD0vc=
`protect END_PROTECTED
