`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5bCFQQJlqhTM0jgFyTn0R9jKzW0ruNW2ypms1nHQ2pWE41KlwOPKTPdHToyYmWui
fGefdGchWei5RS6r3Hj1Ub7j6BImgFIXEnOKJbuhmcHJA0pVk03ms2fx14zwa09C
d0Y1nfwlqxLuXVckdqVNMwGgJGyknuvb0A/hw4lK368FobWDOez4FOljCnFl2xmk
3ssbPR/I0Guh3j978C1bT+LLImtytygGNUE12/+/0aGSiVzqRiQ/L65t/xlH01Py
LTqZIeMKrdbECNKUgMkew2fP1dh3OkEElBJoDFJR95ZRLRglII70tCJBpYlv2uI5
70mIatnrNmV2CdCBresAwPMml5JfZmkeFxGBenHN0IseEOrAADvKSD+vBEg9hkSc
4mXI+7d8tT6mKPwbFMxFRteBmz1r5/ptwfzbdXEielXVFY1cPfhpqklPpUD/+j+T
slDz4TY0LQmcb+r52QxmC5MWW7GKEeJ5XWDf86ZKVMKRrQYJKvbLwDl/hGUSfkjF
z3H9k+yR2lYcANwJu0u3R9lTMZfgAOOc/ifhsmQOUx65neAEmaFwoUyroDdHMI+x
axn1GPXJJbWWkirNomdqOJ8jSdkM2PGs3AK/6klONX1+mQDV30/F3drGu34n/L7H
JVDoJDGWxspKU9+M86wNc6AhusshFW1evvTWNtYgKG1l+MmkhHIGNF17vCUdarKQ
xs+81BhlmtBzBDIPgjCcHPnePm/XyHH0znGTyu+obKZIJPdrZf9j4OYZF01Ml/Dg
H6I8P2zPv3zO9OYDfelefJ8jW06wPUONXWSPH2wHWenEbKRSp2OA1yepHpx5rzeL
V/7P28l9wjbMMFI862JZRVx8UoAVotuZStNhRcGh9R8nyiRXIQHdFNmFgU27hcrA
dyvlsrk0xDNI8oRVx26kONUrmgHZhRTzAYFvMN3+30dz8LeXIirm7yRxNHUAtlhr
Ll2NFTD4cIDFpM+z1qdP3N1m7LTIxXC1Oc+aE/xLxRo=
`protect END_PROTECTED
