`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jY8S6uJmnWuaWwKtAtrQ2x/f23yHN3nhRq3boFXznuopK/kwH9hawkd2OxGExt6q
nX0fXNsZUCR31RfrcjKYrRPv7jGcCsNlAIVff14V9WT9zG97B4gJmbznt0vvpRHy
lmR03ekoOigxajALwQOuHh4t/x0TvTb4OLv6Aq7w+RHMFx90jeQffIJ4bBO+JCOs
1fT/fhbQQVRe8ECWTYVch1OhUPVlg7V2TaIK6VZaPFNlVdDHIfJA4vohuwsO3jSS
mmxzttmZnp9g7BwpG2RbUcaHFkwtFqVchqGUwDxRT/CX6iQ+7yorgpGfEUlx9VCW
/5uB4eIJBhbniOJ0i9/pkkpxVYREuwR6pRsxBY4+Qk2Pqrhx3Gf8UMBBUv5vozP2
4GtPBfMgp5vLJXTQtFxYF5lbwL70otY7zJMPu3AJNvGys/Iyrywik/TEjGbndVhE
gTBVM5zXXJsFVd7dt6TFIy7c7syx8ViQPZWr6nIn5tSlD9tG6TjGUFUThbwYzjAk
gXeYeq/DfxN2TEPhEm0obp/5+nl08KSqp9ZAV9fCoEKmoPBoUH7yGGpg6lVcAsru
CYO6UNHUALckXk5/lZfNrDJrTmJMtoOQ9Tz+0dK6cU1XgQZtqXuB8bd7+kTPZuHH
`protect END_PROTECTED
