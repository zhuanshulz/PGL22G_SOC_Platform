`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Fp+vaRgFw3+lFIoETosBg6AWMs6qrPa9HzvXT6cQ9m0wLuCmugxdHgeP4mrZvZHY
FNi/1IgV96fr1HcauMWUcP7JxwPR7dAxkUFGfbYV8A9iV54LxiouKy8RydpmEISJ
9f0FGKRvB4C9noIvEZdFbVY3AOxeZ53g2gQMOY6A/Lg7Fok70mOUJwSFt7+FAZJq
ifSykWdtY8LYwTnkaJNAsL4ZqH9SnAHVpHhiL2wt1GotVQMIPXStzYh/JFGIIYSX
osW3GbBBlp7UcXM8UzXkyqre9OwweVj0FwSZ4vVOQd6qYZtHwyleBAubODoy6kk0
zlYVMVcOgZvc/2iRXpBIUA6+RcqpEE4tN1C32qutebmN8kbhb+QAxm68CQH+qb26
qOGCgBAJGPDoS1SaQHNai246rmtVit/yWORyeQpCvsk=
`protect END_PROTECTED
