`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mn0Fa6RERed8KFZM5T3t5duRwjUWl4f3I27vAj1L3go/Ya37EVkAbHESC1cIrima
5drK/EZWMMnCLdFJ11QPGZhGjTbzH2uWVyCPK7ecCdN0zXYDoFH6wRfd+oIRvcfP
OCf2M/+rLrqMamSqdQtW5U/QK9Q7hoNcMzK8Nfc7nx3W8iKR/fvjhBt0zac6cyuN
TJ0l0pDDdir2HBwwb3Uw9K4wBJtHjLhnDjRthTa1w021T3LhyG++46jWAn0a2+LF
cmgo+pIHDB/hBdZDEnmuvw==
`protect END_PROTECTED
