`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qhTZdK7y/KAQ05n6dYmcIiT1UCvahToGkAEpi24XABnFTtCp4P+b8Wsq+AH2Wwbh
+6vE2Y/X3CA82Lwnc4PhiPgeyLPEtGgrpjiiR0pgKJOmVXSP20JaFqvz9OCFrcbe
h2YlihcQqCQAS+BlStOI1nMFmV8gxksfOBEIXo9H9SopoXdVlpEoB9SZ+i1yIRGk
yVJZudjX/hnq6kUpq+ecTID1Lwm6lP89jEVwrjVPSjEzGmEGXO51j2IV6Tk1MHRV
6KqOwWfapHwjZG7ym0c77OFuOzpzMOt31lC0/MKur7wLsRKzDtiOGkudOC0dVREm
TdayPwxBjRhrjRomv31eAsQw3vWhZXiuKfNTSF4GnrAJlJ2xB38pjJqBnjupIxVw
vO1mN8fP7CDnAVMocCtbHh6wLflRcd86oUj1e4KsTZAckfjkQ1o1FEYtRrhswYE7
tNR6Bb2ITcyvZDYY0U90uj14gH73stA0jc6iKtwVk3dzOkS350XAIpw1sKWM4kCP
5IZVhEUaytoYq8lSAvTpcKCVXLgt9BdYNQMRydreKvA=
`protect END_PROTECTED
