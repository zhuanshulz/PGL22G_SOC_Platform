`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fiVwtX/onN3JAsUDOCr7LBp8u5+YVEIkHCF2yp0P9dnkgG7ZNFdFdGdwfvXFco2U
rPzK1NbBE4gaoUMiPQvq/bKY/Y7YEs2MUX+akFE8jlETqXZxbSHRlFxlg8II3L8c
YBPr7gzATA0oemqP/sHVTp4DTJszCWgq9Wb6HM3wlMnM8JuMbbaO9t2cujchK16L
dTXA9qE91jUrAuRDUAVsmabFm9A8ghV/d1U9WpWdYCdW1IXXE/bXVuuMVU+TblH5
mHZtSuJlGo3Yoh11B3Y32fz1frZP1vKJz8ZgI7JTpm2clqxk1MsdzsNxwJluYqQ7
gDBVL3TkLoLmkOSSBN7tN0tA5PkbK48HDHD50UZnzK1dFg3/uM6oApvJXoPKzhRB
7dD4GTFWk9tNEKMYW1hhTVjUD4HveVNRWrkEBtIxYRba+K+JOyhqxYfpZtz3ooH/
8gu7XFUHsVMIknI/YJ3dOaPetufE91e+HHHxMmS+6Xys97AtNxTABm4rveiYQg9L
CzWEA0f+aI+BRSJzzc+7qSCXLSKtjMcMYV+ecN1TdrA+6k/OguZKZXl7ZI8Mk2wR
7kDXtEDoM3Z9N8HZFAVkOA==
`protect END_PROTECTED
