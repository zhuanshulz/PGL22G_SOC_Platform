`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C4gyT7HU4UyNhuKFz24sofNk1rr8VH3k9Hwg0mRJxXDf+yN3qytT1H2DsUqY4nCH
fpa+qPcDL67db7yKX1Rv0WzyqOPMA1uJR9oC7kRGXbedKUFYJ/IpYMM4IVUp7jir
aCL9JDzPkAYcmW41cuO7WLdjDBkNZAKys8g4fGlUX76EX9SG05Ldm0YaXDmFH/UQ
pHD7Jp08MZXrIH1NZ8YZs9Qd8zRBnDhMTGWGW/ru9G3fJmyGn3C97RTFJ8XqeK5X
w/XkO/7VvtFya4jJeBZpEC6xIKrqRTgibaVz/jSw+aj7YhBePlj7MLsJpmQ+7zSM
er47iIE/ljViyz1ryVGx23MYeygF5RIuEnHZ4Iu7mpiri5XoIVe7MHNVod4oS693
iE2TOmSo7xPg9Aq85HC5KXON2Ksb1wUzUfnZmTAQVsEzmpILUS1ta4xJP7iYp/wp
IqBX+yLQSZkEWzcKxkbIBREKpMtqIuTvEt7ok4qhx46ZH1eqkTli05x89tFr1CG6
3h86rK+hft9+fzv/u/OtWQdWO1vim9IvqOvnrC5EwmZep+qFzsDXPeiuO6asqnmY
eGDy0QodnNPdYSNkR1exl110ueYG/2xOYDPOeLbL4cPlkpvIONcHEDvGQnSmhdOH
vgtfMYx5xkokyYnSZnt7q1QXQEoIFARGSkZgzv3QvXLPPSatbXFAAggiSi2/EgY7
TAp6VVkBbeb9K2/u4tXB5XnVTWHZM4AjhlcJam6YDpyPL0L00mxYDi2LOE7vAh8i
VeI/rUK2iaTB/CU5IswaPhad1LbRls5DvKnK/f/09UF1VKiXuNH9ERFCeHM83E0K
N3bdtwGsxC29QLEa5Vx3G6zGDrB1CR0TSK4vOpvnat7zmmCHYom1xL68l8ng0kIX
yLhLERR9+KyaEbMlbIRO4l20o/fQlbkttzBlAyilzayYu9vv3acVXWMwIodFiBdH
tqP2TTgm8f4sxP8hMkPo8kSQTBo4EVnaweWKVj8u1RgoZ99TUZqC6UG6DV+MlHKN
oDexSE6pyGhnFLgoby2rwMJ8UfFKbihnsXzDWniFwEkDN47LphPqtk+6E00h9YHr
utxxqOavQD5Tq2qB4AtocZfoPsYu/xwpl6REE/WeevQg7arOHpFErMZ9WpPyv7r4
VhRVLHcXWsrZClPsQPTI9rHbwxdFsWblFXlccWu2yTeOvblLBmYG/R2ldfrDVrGd
4rYaHdQW91ALkO9mdTNKi/mscqQ6rrRtRSlFkgaGZ5WALVgAxq9ibOcpqNhPhILS
6wMDjbsE5yJPM3UXR7RduUZXOY7G1MRbv70mEn/TszDQL8GiGZZ9sFbabjKiLpdi
Hv/feuLgsydq04H2vt4TGHuDrESYwhMisLy1mnU7ydHdJ074PujnFvKbAQcwT1lb
02imJh8QHuWraF7ZdL5MKVqHCH6JvkI6ouVhmsQX+cQACphfMnz/bNVSB5/KIa71
nKk/cs1qdkut5SC1m2ZSrdu3rZetv2F61cv6J5P+gfY2IAGSpMNIxt/XerfOG6j1
rDm3Ir+qALh5uwWPE5M7iwwFBOrQnOGGjnKlF7tRIlVlTl9BNVOuhXTXPSX70PZw
4Z3hrHrDS9jfo1WOlwlsXGVPwdjSBFj4enp/Q0p2ihFbrbX8xpNx78edTNUFUzWH
GF31AuDleMep9tXURs1lk3zLTerDIuEk47TAs317A0FXngZTssbMe3dVSBvRT4DE
1MZq8ChiB8uCoE8qWN/bEBhXkVCiddkvcEeffEhd46xKSNfdapJwgh7guY1N/CAH
570ab0no1L9Hfy0S58INiXBb+sGYckipRHvlwvUEdD5Tb+KNd7tfFCWOQ6c/8OxM
xPOs5oPDs276NVdSycVLVw7iQp0oRR71t//ioxgKvUrErTIFzJL8FZymf9jtgOh4
UsxS7bSQlZuzdvB+G9tf3AtWvEQWyQcNs1piFWaTGZpUpEpcf2aNjTfZvWOu1qw+
Er7scTiIqRKot8KghHB7nOVCAjvXegADXQ+zGiyLV3hvgtqzU5yJUMOfawOu4EUP
GE8bZxH8HCY9QuwWJZdCmJTGA4viBM8+O8JhjjeAMx+41cPgzcZbqdr2XU2Y+x/k
8Wtd3Z2bGJfLh2cQj4nvh9uknkM/P39iORHyrqEc57wc6Goby4EcDNtRS0kfzzfD
rlshIki9NT5r7v8+yC/gFoWcQKzAPs9tBn3PFD2D75ljDNZBmsQ6r3I6m1l1CdyJ
uYbo3sVvCLdxpMm/RkbDVbdjigp0dxM3bvDyAnFA2clS1mWZOMYq1u0vfTz26mwT
MxgQAmbVciHJ12MuNs1Ly126YmSHWHswmKZk2q8NtVvaUVA1N4keWRkPv9yjVbeC
QzMBfvvV0eNFueNlddJSfwFX9gQvpkEWbWLm10N6yzcHjsESRrM1zkWA90BKw8Jy
fDnGoHml1sxeYnJsZ3iyp7ceZuKeaFv6PafvK+YfhafScXFKDM3YmtPmpr8FQ9Z7
HnOTah+Vf1YHPn0r8MCtMlGq4LWxiFf/TdY/WQ7e4ev7ataMUxRgXJHbs/VFxnsF
BjzZt7vxr30yxJvFcFfinNuCl57Z0dz4PjNIsfn3J7xhT7wEbOpyZO0VhuaG4rc8
wIvM3CJECgy3igr3CvfoPUXzHxjb3jNgCyzJKO1zAPQt/VVlVB54AydXECTTtfSU
dKSCO+8KyE+6+gLP+uM3KL0U2VDtktSaD1S1cBmESZ8gqMKKB+Y0jOPOvbuJY7UY
G0qDNUO00nwMeCFPVApmFmhs/+5LFB+HLNimPEat1d8nSeutmY8F7fbJFv+7QyR1
ZOleiBsrPWn/V3ukLoMblX6J1HHxbmtSa8BhPaE/gXL4i6TW163R7eXjOlDZvOGG
VNotqTly4cvn4aH3OGsRhtQhystoPndwVmfbeF3e1pnnIrlIjLJDXaIADXrG4oz4
TubQeDg147d0ren71ILVJRxr4dMyKUHnKH597PhnJIKVCybghfFyKp25meuxc+t6
2XLUDctCEAHGaSDhFolrETnmV9kPXYY43kVM4LW/CNinnfwAHketvG0mFOqJpAWI
t6OduqTZoiAHyDUw9jd4gLBTdxrOujuJwm9/24qqmBuYuRKRNvNvGMjjYYVZPwQ5
yJ7rWeBY6aXPPlwwTVWCwLaKp0B+fgL12t/W9iIHy05HAdwM02zTHBF7bnGfzWIr
ez5+e/vJlI8VqKPQqLC5rFuewjjumTiymlJQmLKMmOlbMJNeH2RENTOzh4otk/+H
/wOD+OXN5zpgYI9Srdbx9CrEx9o4Wdgxwm1TCxFltqRpRRcSvYSqPKeFn3sJswxq
zQKpH9uXl86osu5/PCPgnXofFOfYuX7BbfGGsTlcRnLICK4ReC2ok0i3X3b5gEo1
s8zou1Rn2K19+M7Q74H9XU7QYjVk1uqEXqfMEXlENvp8ZhHuXW2Df3xIKXVKau+Z
yrHNnkJxW5rUkrPd7C8EBJiP8v8mcn1wuShno83GjEUY6mfBM0sSOxfLCMKaUtja
2+dEQyIS/KCTadmBXUHr1HaZJr+5hdn8/4mpXD1xCbmesk8BOYeS4M6VXPflzK/V
c9P7e9MJixgCZOEn/1myNwD6IIWsWPeWDJPnfkZhpos4YHAXMHfkygLl0JNmP1Kl
GErWwH5lK9E5LTAkBmqrLRmk0xpkM/586yhuRCe5ZUJs4SyBDGmmM4nt8FVR2GJo
yuTMt+O9aq+XkYPG7BOFaP0DdMEp0zsj1upCuUpSoITcis2Op1y5CBh2Gv4d+1cI
OcWiAC9nATKrYDqWvBZghHgAz7xeNNCwC+HOueLzdzKavs3LulBK9Ymr654WLEZw
J5F0Wix+xc4PnEkIU3kAFQfqQpOAFlEz74CjWio4OIeb5RkNI+1ijtB8td6Av4O3
8TcIrkeHb2GDyytHShE1C/UNnbWHACkWj0/ABPdHOchbGjpecA5TIEnvNHhi72Q4
OcnjN1L0/FCAfgZJOfEDqaQn+DH7vJgIxZMJe/IkNc+QSh4VA20qI8KtYdcKJ0vd
lCbSYxBOoyCu8lmFUI20koCsoXxC5lAopfjlTPrGPpQF0Gxeot0ZP8TbL9pbGFI3
K+TuPOstzoBLcIg8v/+cFCON3J++8VCLxhIM/bxzEDFcCCPVxvIuRuIi4K0DQWpG
luC9MiYe5fvdonIwqTp9QGjRRWmp44ar34JfZkX4bL26eaW0kTKaBAt6OmOSuzyC
`protect END_PROTECTED
