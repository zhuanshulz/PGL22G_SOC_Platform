`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q97OV4XcYO5mmxLSnzGvKbVpSzsD4lDvSL3/mXPR9HXSC5ow2+fsvRs2eDqYyKcy
9etMFsqUE2suCymdEmLaJ4X16NqOOVgXHdoaEFxtXW/F53Jjfz82AJQSN2sa190+
Lw0U+7YUh99YHJacE1r6ZgdkAvGQ5RDj51pOmApp8yOQ1nwiVtgi4uZQ8XYedES9
S3WQfMGCy25b1ibRKPwwm5M+Ug1cdm+XVyAnXYQosFPqfSiBXILVP8ebXNlQmCAl
e4LH/kyz1+MdjIjVt6BiUm5E9SmEuMfp90FUNCaNLC518uORJ9pzGo/0RjH12Er8
ZLjjxKapsB3xADSNO62P89F3Xs75uk+ljrGJDAMFyzo7DNzHn/9pMCFFWhw/G9Ke
EQCGvcYYBK2RwkKvxKdgKBivomUW0MNCiANDdrHBF9WgZ15bQNMsFRffI8Vt48oC
jFTpleNUiKS/Lnnjt6Og7eXe0Y95MyByFbhvk4d/B15bv2QnjCVWSc4l1oc0oFL9
7jJHJUW/QMz5iJA+nRf9T3R8mXQAvMleS6c8xb0i1MqVriF9xZttDtTKBnIvykTv
sYTU3nIgEHOlcZNdFj2ut8L9aEb31qhFq2rO5pR0Nu64yC2Ks1N6j57o6zCty4F+
EFrbNTIKnrqHgMVdDrx3LkAlbTseaC22s1eutBzm++gXayouqqP49Rk4vuCkZBXx
xe8yKgvuDDz4t13hyQs9j5j2lpBaz4plY5bw0YGUTzAsAPOQWax92udCjOfX7kMG
WKS3DkIL/seDCoMsUiFvuXsNwqKz6VxHDWwuAuvvFjUYaZep5NqG/NcddFhI1LAP
HlbWLk7zvsIkU8LW08NiWo+M9RCFvhkrMSRBoO2agrqNYe/Y1XsCOi6Y8xKhPU1V
dLgPwQgfvWlov6ut58xY7+qQ2bwGPi9f9FeE5d7boTmsOq476/WhxtEYhO2PUepg
DdpsJsyoDBTFhhJALN8bqs5Cap6eb6mNr6JjdGxR5P6NXfEcpzaYIDllLGK87M7Z
eYgNbY2YwsIR9/YHS6qn71M7emO8FNKD1HGLpaZ+F+qGScY+NacC68z9pUVeI4S9
`protect END_PROTECTED
