`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0bfv3OYbYiCd/m+Pk0t+zTFv/RcN/R4Mi8ucOEeI4g9lPjoG7ein5mAOCjoWYODN
rkxD0LG9x+cLfOl5PZtQ6BiF3Uyd8ezLQR7JtInwddlQtaM/3unQcateZen0+BeZ
Ya/+6tWSXhsN5vRu5SnYnBNMRXCmk2T5E1RoUzJ5o75P2np15yPmbGdIGRFzBOad
11pWR/WsJSgwKUO0D9IAW7yRAJbkM9HwS756JgR1wxnqccxhtqui83/PVTFKYz1A
clod6G2RQIFo/wIFBbNjpgNZWWWXgkR9MU06mKXrnpZ/7B5VPXbXhzwHjDOGiPB7
kvduf8RyLGp20RKh83rmTlzLuAeBloDA9RPpAcfaDgmkU0eatKwSLoy3xN0SzZlb
RN1zPIGDIjwbwW3Z6KoyG0aXFepQ/srDgJXMwuXa5iJIx+IZ2ZLkexyobMCbaScx
CheC6Zhd+8bS0FRjKJe7QmuiyRXYD9dOFdnhqpM8/BVj94lCLwMKw9j0NRxgDn5H
rspB3fMg/iIQJUgPrd9p57FHOmjzPuQn8iLjzqhQWDubH1N/xYD+3oCN5ivT4nJi
jG4Woy7j2DJWVgbttyqRvfcKmGzpq05KHytHrVDAQXcToGF3T172kljtbfAs3L3d
KnEMLf461zBmtPnPfW+WZ5ji0YwSVTj/iTCNtbx9QunqyegWqY+oIAX9ALnuw3zs
G30fZ99NbAWDVPKMTg2Hn2WuTMyCkPPYQiluH1KOplGXrnP8MdhMZ135mf/KZ6L0
eJPymj/In1We1gT2x+ewWKNL14IzfQTWEihBF5X1OrH5qJ/KcJFEW9Px/FgGZF9u
mHT+em0Z/sAnlY2aKCQ4y+p5BWdfuT/0g5V5Z+Xf5eyS5Fnc8Dq2/9c78Lg5mE7f
kPNjez/KipBAhW9j8Wc6moan8jCknUcyuVlqb2PMgrbL6LiDCvslzqGM3R3YGetq
JhqnUIITq5TcrvI6yIYQyJy4MIKdCciA+Y5qxuAmqXaavMEXkJj60176pYTG87Oi
NJgidhi8rlvsDGUC+OqtTGs87e+D/FLbVrIw0gpIfUKIYdK1qtjz67GGdWzHpK5M
DOHG3tJYyaEpbnPSRdjA9/U2P2F3B3r23+r1T9Sf71Zp5L9dLFJT9Ns8auA7U2yK
QrCsgFE/tbhtmQzRvr9piucOmRlOp0fHPqnK3Kc04CZj+Eq89h+u5Iv1MV3x9dLZ
HEDcjwjr9lXl15aQVwpnhnPT1dJUyh1i+6FRWUu+VSgABTJrAw6KwLej1fo/zJo2
mMFUuA9VbyyFAx+Jh60rtP3AuaKpcqc/+vs7duP3vCFqszcGLdV9iGiEBQLicp4P
ygkn9q3RupfFsY6/TGBAKkY1WTg1TgPeC9NWjumauF0ITvhKwPyxU+n8Z+1pVtXu
kzCljMkcRBTskDg9TiH7vWRSQbvB3IxSOc9ZIYcIPuBL+dzWIxgFemzyoPYBbFcL
0JCM0Bvgx9NzZ8B9Kt4kfs2ZvGmebh9JXHc1xfZe3pVj8/zwhrJakvGh0LBgWr5U
BDQa/zVarHYKwXO4Gs/d7yH5S3t8LdPqtCME5QXlKQNGi6+ZUIpW91gx39vrjJN3
hHYuFUanehJcZiXK3PjZpmMtRtq53BPH9Gk4Ss8cbbx/e1UiJ1ouqQJdnTwempTi
TTH7S+e1a59VZRyE7N5o9d3oGBh9Po/0F04a0LHk2fu/2rSZYJyIFMFvw6Pvm+8M
YoqpaJ4iT6iM1v4Mvir6kqHDtEjiI495TKFMdgJQnsETlu9y369oLY/2irYPJK4N
3UFWSDM+Jd08DjUXfhDBulIYVTlC5CYAg0z2C93jvU9zg1GQJj7zVwgHfXwkAwWv
IqSLJwoAE8pr7c1gp8keOu3OI2BqP7KjJcvmytl4dthCa+85HFZQoXKwpp4TSZc2
8ahiBrDwl4jxogN2iUR+98GU9BXJaPPmbTDmFVnfdgDat8RoHZY9HtSQbrnvQTiH
7/m4NR6v3QjNoUSj6ishcWmEjtiJkdbAWFZWDsX2wcsqt/q5+VXytvhghaGjWR/a
BhHELqv0zrbZIK3OTtoboeiJYrHdeAk3Kqb98N/Ov81doN2LzyxiRQSZPM9QR+/K
ZDj8nAWspY4Yi0NGP8ZXahDnvzXtzJ5e5Uo5pf7r7E5uwCeYqKEXGCcyMPIYacaU
6adfCM021aZ4aDoX5K5OeDsnh5HxAS3bksbW88lscsjVy2qs51ZiUVkrVh5v+1De
kMwQbyV6s5Q/MosVwAH8puowZBWyBQDBcCc2vFWcvvXxvB1sm1a3JQZNrL5pT+tf
e/gHsy0J8LGar1Rw2BvFqduoWtkzXs+ZApRhHjltMB6uRydnC4sSM6KRV0hZyo9F
sMWoMb9PwzfRqJnRfFsrYqH8SaZxGU6WYqJclVQQUxz6eA/DiSWqjl51jjPK0CLj
dD4420BJn+z21cANbhTxcp0A4ewIyybGZJQqM8jmnPnxGtO8rCJ/gVpBuj/BM1BG
XTzql2onE9yL5/Q0QtyYUCx0XIyinYfeBRignoL8IP9k5a64U6qprjWI3a74PQID
btKBPRXdXb47L+9jcWhtD4GrIcH4oQJ4mHm7gJIb4xys7oJxvHvD8gYzPmtNKvE+
+z0WYvV6ToklDfOZyR7GPpj4vDIJWZyEnPpcLmpcYq8O6zNIl1pDd+NbmOUjVNmP
K/ACheELWHd2NfeEkcN6DHYGv8AbaPwlVESuucPU24zUnfvXQ+c5awq/V/iXCvIi
H4oUq2Qe2CSBmpTlDQWSrM2iLJ8g4Zctie7bPPNIKataf32AZDlreiS97BQzAIyM
3JTrCvi50/tyeJ1uUtOuodE1jp1FBZNTNKKGhdwoaXqTA/zJ1/54LYHWrEPwpqbz
mixQSdlf3MY1N1szA0g3dtN0VqaNxwUN+81VSPvn7OKrC8tHNnheLGp7fuIxu2A4
5iQ/A10Cx/WW7pFO1ctOmOfOZoFL8TvkH1A9bLBEO5XfbmA1CRwIrz4s1JG3BmuH
nCLRfyzFBWdYiYuLk9tD3LxoEzJ0+usM2o/VpQQ5pC8tOm9jA99qR0WyEvaIzUc5
W+fLblQGiOrRMtqFCyw4NI7eEm3fLTrqUh+FtvdMc2scE/LV/TrbmSKidDkyzmP8
DJV6Mj/DTv+wvW3B7AA5U+HuIuQgvqpuOL8toJin+lM366qKV7XqetmEpv7UtBY1
g2WLF3LjF128bwttWqdcIaQj/uIJQ7c+660l0DwfkxiVtq5E/rQf326bOoRWObz4
5MHprrmeB5aIwKkvastF2+S5sGauaWbTtMSCNjG8okSClPzkbX2HlKKYtoyJYFE2
MWFWHL9DEmmsQRG/MwyPHgtlrsEOn83AibG+6guq1t6KeJjgvDP9muyatJb3toCs
zLmeVkCV3N75oWkIWx9GYuO95Y9dKcww1BXOGW7xBZVqab++YWZLMipAZpSr6flz
IjDBGQ7KO4oIerZeh6LdrYYRVtnxFWrJi2f8zC8uJAc=
`protect END_PROTECTED
