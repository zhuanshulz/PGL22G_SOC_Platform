`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Pw39BS82qTReExdws7xEeYyTbLj/MkBNSoH6hZ0FydFPR9SksXiShl4AHeWeNrVO
ISEHYVgZhCa4UsqpBcc3xVWcflw+xh7AsMb1XfGFGIRWcfzg42/qtcqXI2XL7pHB
OcPefLt3dTPmxiCQBdcfxN38Hyw45iTFfgipK8voEC6lQwa5dJzN/oNJIJBE/r3v
EzwaybfGs50Jl3Nc5ZYTpKFHepL3a9hvnJaXSHcZHN59rxjCuS4swvNa5DFzCt4b
O4IppqM06V39/sVzKA8QJBXG7lC41v6aJq/Ou5CdyXtX+QYuDg8ovmIKDLhNZOu0
aISl9di1cnbH8LXBl/gNMQ1WSZ50hj8zkQqIaVVfFqCBb68JBuCAxPlVOBLi06Uf
wJSyj7acLg751TK3TM6u2SYpjbDZksNK3hXKpTg+s0ykZWHfnoo6gSxo3p40Qzun
pTJp8kYpnC89uhJH0Xdi71Hu1AMHi54tHkxyEHb9/ONEKJkHWAlzMd4u+CqRkGMD
2xSZrgyXscgV4sZ6tFhLhch/okBnkoeXENfPJSxVkvqnOeQnswFjdzXhQhQLRec/
oPSxNwvuLms/AGR+4SSecJcOwk5ChKk2IPtx/EnGwDtBGTvrrfaN473ydHMFPYsL
ZOKycfFfbWEVfNdFPv/g03v48ob3y7Ff0aX76vvaIrXGhfkB5K6YjpLH5M5SFFyu
7kRMethrnfhDsRHoIcLdxEiWCQsToqZZZTDFYRZe7cYn+mr6Hj+ei0F4/ZURUoV5
Qwh5Oo38ILJXeb+ORnZdNLp4MSl3N/S9JLH+9+HNMeWGESG4HtB5KKfBsyf3SJOx
yHnGPJ9Z9cPUQvEuFgdD57Se5ZGJQLWmNEspY9DReyxA07ysyxiCYEaFshI9y4pI
LjXFLCyAwOb+vSoRGAXhqcMFmE5nU4PHNJiqBiB0JXnM6j3z/84RH6AKAloHSE/P
142ZZ8YcWkiIYqZOHNOlyVizZYEqa+s9KTv3Rw8pXxvxDNDnEkV+injDlswts7j0
8BiIjYkifxjScaYtNSmilslAF1pUFRl5MOw/39dy2uwJgWOuT3D5Evei4fAXRrTB
1/YqJhfa6W9G2f1Bvc8jpSLYM+SjtoCuJ6kcBnDdbERTlS/RycaUW5Ol/zOQPV8Z
qJv0KJ7RtwNj2CbyvhPzQzE+UhsG/Hk817SSoIwF/Sczm1eAYaGe6RAhrGEO7xVJ
WxaauK46tqEZy/H//nNP/KcXquP0bll0sTJHaEMbFwJkzLmR0+K6KSjaKo7wlIIM
+PyA3z6nOCOXFYvjyAu4H5Xa3dZjM3VGC9XGOfyARNRgPAtPW1r9G/nxbTzsrTvT
QAfJe0j7uHdKg1Uw5Q8+8eszuEn0QISm0SNx0Y8+WQFbcz4I5L2AkQqmaJneWQ1a
5Y/mLBYjxwPe/45NAMjSbX9x8NvIZvfwqlWnS+2+0O0/ZYPKAM76tauZhvTpwunU
783yinLrDBf3qshNvrpQCrX61QFhj/mpow1KGiVg+CaB7O7MJvbjQzzFohyJ4Fan
ga588rL6/U8yAzNytTcw8z+/iwLlrT4SuRomtvwTSVE9tOeGMi/4f5Fie2JIZqce
ohiQWNZrvy7LGhLKwW8MDTbglE7weTl0oVlE3avHqhJ2X4KrzqpP57NCGytoZmdF
dUoQJdp504CRwFkt8S4JHXr1HkA2bfzVRK5VBAg9PtrQ5X7FVHMrSpX6VOD9XhFA
xHVmYH0mmubVjTlNfYdLLR5ghzpIEAP2xiEz0xwWLA89TDnS9Wpgm632DWHRETtz
ZZW8x7mER5LGWREGyt2xgmEmfOidumdM5oCijLOqJgY7xuWfWOnGUUUiwGNyG0qx
okKo4D9pxT4fUVREofbvnK9SRYIWDT5gqXponVcVXbEBRt2k211oYR7a/Ube5FnM
/K5Djm9NC7hU8xpLCZuOQe2CY/Jlg4IoH3wR6r3vm2w99uqjDhaS+0cBltftK/yN
5qQ8voknqGIZiP60ryRdFKhd2qwf2oL9e3hpLgyFm8p38k+hc7g2YWadG00O1X/e
3xQ5AcKf66Adtg2LaV366qgpy6uw/sC1aq0NBC5ANbFV/TNFVQ3mR2U0Kff5dUie
RcbFQ5n2ZlgDtfE3F3o9A6OqwEEXI7jt9fUfpOzD02ifEKRZLwb9Q2v4uDzLrCY4
lkDE+eSfYnXnh6E3pAEOw+a8EKMkc2C9xhD5LVsVMM3sdAb8V9KGWWfFxmK2i8yp
DeK+OArqzrjUGcSHDD6VLY1PrjSfjPyRuiSXO+SKJiJdp55MEwnbA0PHim0ZPoBP
4KLKrHDj7gyjifhIFkNEmdSisDDJ1wD57BCn1DcWWhVNIA37pPe7CcjWb7uVTsbw
UqlBBL3xclJOJjsL1867KcHgbiWcVfg4It6WMFiVim9y+v8CIZuxqMA5SbHj7JaW
lACuQJfHttSYiCmJ8qr8S310DDp+UX8EerdthLH13WaYRPEYeYaFrCdogIJIgo+e
OFUupYb/UPo/sK2HTPofh+b1aPpYezFG6Y6b0N9R1evyYm90BDXyso5CZ9lTSgMu
NtKc3HhD7o4A9zj7gcvBlb3ikCPTLdu4/+02Pc86yY8N9OKCk0ryaPQ9nmZv0OoJ
DPbD1LV0dY3otXNQwKIBLfVNX3YIKsN/FzmOGm3pRwBSyulaszw45RHzVgZ/otUl
709Adlqg9Xilfx5cLAbiMQ49Qbaam0HhYpDqq2XOFO0vrVL/Cv9PC3Wxee4d99+i
e07cfpN7U+QidulXbxwufVgzIzMeWYQZBJGuHl0DjVCgPzsmhD8rmzk5zFQLJKxE
RO94zfV0LqKMot1UebZQZwSR9rESXYsiLUYGZmlo5CdjlVp8ycMaKW3K74oOnpau
RyUmXVTwS/G8r3X77Wisd9HpGA8D2RVKQE+F3L1g8Q/fqZLqWHhfDrSmg5d2V6+K
FcIKHmjpcgKswb5tz/3cGN4Fz87dc6JuVuXKPv5Dd5LZ/JeA3vsK7GYrhDKUTar4
mhFIf6F6YF9HN9HtmSqz4I6RYwHZb0ulxHbQAHeRJKebKB6FlkYJhoc8Eq1rGn/H
pSiWO9K1vo9V9eRuXBfb5u2t/gUiRJObSd31qlxwYCW52RQVubk+hNlJqwEiWwjh
MorOyRT9d4SJipElwzZJu/bi6b9krQNzntqjaX8zwso1LCbC7I9S1Ja4kEj1K1uX
3443hFf7019LBe3fIdNcVgSPFDOa1+m46Kpds71MwiUjME7RzCvZBgSksQzEluoV
Mv34o+Qmn8db8OYY03OaupqT29EKAboeNaf1lYotx891sJ4SHo6wJGSktJTTaX6q
m1TtJ0EiKLwy7KY0YrhQMLbbleNF7PXeaoH9W9O9ofznS3B7XuI61KgFd0bdWm7C
yS9V7dxKMYZ37dIKVLrXrNfRqTbzUnaNK9G1gdAoUC/UjM/OsT/l3fC1AlccHcI+
x1+tM5AYT+JDdexZGL31F22Y3Ylwy+QAbWGu/Izu9kgv08SKjSWZ3QAVyDoHNMuY
lhfJLKzToLgYHSN8hO/lntDB3mbrDXm0lscBdDA1sqFlqZDM6wZuZ/mZkb41Wm3Q
292IWI22gqILPh9+yI9BgV6brjzewwzZ4pXbhF2up0icVA1IG3JJ3L7pGA9pcou1
IU+hsm+fdvWwoJMu1Xk3K0bxV6AXVAd+WAIyh2EGthwMrG7ZS+2ChmudIgGY6gZx
xTndYQbcDK8693WW6LH47RsMF43i23zr1dEej8RoxkTk+0qnA7PdccaQPXXJUrHR
Pegzlmo7sLCVZF4NnnQ+Rn+kxceMWnr2SAwO0d/uNKDFmdLMz0ieS0rnqAyXvj8M
YIYvuiBW4fSC7+8AH6EsI+B9l0bfZztzQ5VNRh2oDC5wIqZpav6PeBh1KlV1FRbY
nGQ3Scw7Up6ulSkYrMcLSOSQb2QsapHChS4xcb8/Qk1Ubm5NXhiE9ypWLF+ctQF/
rANP9OBzofd4pmKiCYcWTApY6OCYW8ehvbrMW5bVh6xgMuHgtqKCx7RrUktwwHEt
wT5sGo8GrRssBzbb6mXnVGJ1LBQwQ01I5kYuXIUAfepvDJZYrR/QhuOqUtUGD3vU
bpPXrKON0OyYrpqqUIyllq9MyyDrcd5PvvsUmCflSUynOpJZx+W9N4yoe11OqOzy
gjfFs2b39IJ/n+XRX15N4OFYFAG+LXVyX5EdyF7FGiUUtiJyQXGYVkTRg932ogpm
gxGRYpDnrtA3LUpxcD8qCJAsK69ouhw608Y+ziCvlkUGuMaOxbJ56jr8pH0nKOmu
4Ge5/PF8LFVCROOpyvGLk4lTAtSd6AgRXAckXTS8kfjQOBMcKmLmuMpgDhHHduJI
m8ZqMSbB/JQcUUXamdB3C/19f8aK696OVePZ5bm47z5VS0VYN+O4G73wWBPouGjQ
UhQyie60DWEgBKFsAMN6z455x7Seh+CeFQbhl+1lNCFZzTs5vmNnPvvbBVShqYkf
lSLqU6U0Ef4AdON98ETX8N6e71C8bdcnyBmhZJny/kUbzxhZCqpi3QiaDDIq8hf7
RN4oULoMuSgScEb5ZpbVj8pAhgSWUAitfUT9WLuJZ2BurPUuM7IbbKJLx0CZNojo
T5LYWPnX3/1HViQfW+cBjlDn8Rjra5jdzAM5F5UfHkIN3CPbX0l9e7c+1FcomO9K
eoU8gmCsnaGBLnSWc6ieejLbY6loCcnTZBCnukyxTFZJp9HXBbZn8waItP0G3Hdt
adEDIhYA3ShnxLiMqOdEGZaL2iOBcNZvdXu80MoGjf4/Kx4KRX5iZCaYgJL1qq7/
5ONQVlWhN8h0cg1QFD3lCLr1DDOspIMGg4hn35HWgZdqGAWCwp/5rDBD2L/cs1nq
MN6c5b0T5uFGW0asEcr2jFyKB7zJL50K6m/sWV7UEb+R9WwMdftGzfR2vfUk4IJM
HmcGdqxyr5eBZIrpaDD1If+crEIrxLkJpIHm2AczlkPDvIOMbxQ1o7uLUtuU/qFG
iVxQlH2SWX8a41XThgl3VtSHHfl5X/uV8MMIH2bJ27WdKWbZ7+7Eswh6+b74zIb7
P5pdiKlTGNlnbHY2bfyVEEOraJ2qv1JEvPaixRIMMdsUON9l4e9HAhsxk9uw8ngg
BiYgnDhhVzRl9zS+GTWq47sarXxEaFfloVhVVQm2XWX+cN7ssDfpQveX2ENmfaDm
F2CknMEi/6ABIJWkvqkW2/2600iuMdxjDWcYZOg7p37tLFS7NMouC8bkAvcXboTK
Y/hquuzgeVktVMGd0oToaEQhCkevKbFpdNQMi9X7KnjFg0qsXhjzS9d0TFnvNn5m
MFFdyrUxbet5SkCL5zIM77s7pNEO+McUT89H787ktdskGSuj11BeffvGbQ+KETcB
PsZvBUUfH1XEtDbBhIgoPtKJ4nIIdeaool2Vyq2i8XbDipugUzwDC1V2zCkk/I2A
MNjQh6yxzH374AeNZl1U8u6ov4RpZ6iMYcFRqFFsMRSLoqyLvrFi1Fexk25cIARZ
il96/BkubzUuhqQO8u5ePhZY6NU9bqWEFeLxsVN+GuXPUVc6b9WMIKEAz1ulQDL+
6V/L+xRTI9VDnqFON0gH7qcpqjz8FreKd92J0U7sJOlbeeuGPg0f0Qd95O/yYd/1
6Wf+7WAd7ZbM9c8plFvn2vL/ijYqdQ0rSvBCRVekFtprvz0vqeJWSyhtSsEJQP2z
WI/fXKtZ/fm9FEGSKMlYbHJBSuMxcDH+hpcR77JL3Y8RyELYcx9IHyKIgaqwTEns
EpD2au6eLQrUWDATS+PdDU0INPYXOTkcAa+Sc2BmjCSc4zl22vzvGh0Je6bE+03I
lAiYWfFDHS8AoAT1/Bc/GNCCmnqjDAkl9/qyENJZ7tJSggLvAwe4HuKVCO3BxhcH
6rrlZU6ggTh8OrG9qL8j0VdW+DEc/hDFrD82uAi499I=
`protect END_PROTECTED
