`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TTed7DbvMNGRgSHKmQg76AfPpAvHy5rwNgWG2AxwwYF7+byduQWD8LJOpZl9vwHs
wF4GTTDFOjGAg417rfssfveFoimH8u1ZKpRifG4un/slvuXKugPp2SuSXqy+xtgG
DWPWvh46zgvYsZm7J9b4x5hHx94wxXDCfieL53Ku5Oia7H+HMLoVqmsPJYgphVpb
RjtjTvMo8n2WI9Wvb/7ElRrYcwyfOcICjlC78FFfmydpR6UhizQh+VvaChc6vYyi
CTKl8Y6+aiTQCURR684fCt4lQdaNtqq4A+/z+NZOlz8rzPxbZxAYcl9lrSCII5KT
eM5gIK+3OBbh8aWocGDL+p7WnI8vntRJR0vaBYCq/Nif1rz6gG4QlSZCuv/JLj9a
mD6SQqBZTIuS2rIi41kBCJlfB4i+GZpR2vSCQQ6v5WXnsAWIS6xzaXsQ5DpUR9Q+
FMX6x8QwC+hHKC9z3kRg7EVi8uW86V7zmHDoTJUw6wzR+mjEGoisoIKtS7a/S5Bv
cZ3Uzr90kn87LHCCWvs107+0MeWNM2T1H5ZV0Y+K+vn7g8mtPcZN3lTq47jU4dOT
R5S8zt7XB74rriViAGHgWc3YKgzYINP3Z/WVBj0VGizrEyPEGDKnvAacCkIigyQT
0r5la250ACRtewqmNEMzocesS33Wurhd8pZDA+6btc13fUbdsk8DdBuzPx5lfvIr
z9ux+L6j3ZI1j+gaeDGfMhyCtg5nAg8HWR9K63I+PGnjZkXTNQ8VAEie8vwUmMTi
G/L+oj1ptjz888gZAYuGZzwM+ztALU49SVFIQxqaVmDO++SJ3send4WH31S+lBX5
ymef+rtx1smRb/fjZRe5zQ==
`protect END_PROTECTED
