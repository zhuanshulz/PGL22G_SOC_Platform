`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zXf9CM6lPQ4JtAv1VoWNudikx553g5OQWk4KZaO7XdXniEsbOHJBjmBE3S/ioCxr
tJPgnPTBlUUAPZR6SRCOX9hcgG87TJhCa2/pfSvue4+YgW54sF34XntBigjCxvKg
CESmfikRGxo1ZpnNyALRbeKTkbYgVI0gHDlH5RfEr2ntJHwZYTH3M+aONJMH56P+
/pSrFCUhIwIqBD7usk68wRRc8yyvRyVEnt+aWsNutsr8zxgfBSeP9x5TyzcdXfkS
budXTawB+MQE4uR9KfK4ZvHqX3HUWSIDAfLMJG81hEAVjL35kvGNSF38X0xB/pkZ
5qeCH5uUi+CzjiSp+pXtejKzicrPoHUWq8PhNsD8qaeEGYr4zAjO4t6a0cSSOXkB
tLdS6WgMc83BANUCGU97CQ==
`protect END_PROTECTED
