`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jLbS90WSvJBpvr1R9KpaEjUcxY66fcPDi/WOfP8MuuxWzW5aGIsJkBweg/3X6tM4
pFQpKerAW5FOWtQhYhG9CIik1IAkGHeVHFaqPEKWjAB0IjUdOVFTtLC3TScWPKjt
7AOwTllZmQWm2dhG11tb79dj/8Rgf34EoVlFJ5dmkcJIl5x+habKl7hetN6p/x8z
NdhpoCB1RY/tShY7ZAJfsmWCqyawoYaUqqEBy+8FnXEApb67d2BRAqQY6CIffqHr
le3cy2VovKEz4HjnSh4MsdorUkGRjynnVD0xzivGIJvtj5gimN4qeHcN7vemHTqa
SGWqeQzvbzx54yanGaHcwPVgwPWs2NJvHMAGPl1+MZSJNw/+kug7W1WEd8Gw3F57
8Yrjxo8wT4jBQpw6YdZ7FLHFwZ72hkjD7U1gaOwsscBGC8X57UIKFR7PJGI6sU3q
TP/Pvk3yF7/5HVvK2bEsq+dR4fg2l3ApAK6whT6oF7YKnFv/euTgilsRLv6xrxAJ
aE7w1US5EzWk/ctzvA7S+mLW415C6mTYtWeu0QAkZ1s=
`protect END_PROTECTED
