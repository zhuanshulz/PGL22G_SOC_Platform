`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1LC0PY8lK1pgDSWCQA2wG0BihMrhhY+vGfFSwgE6/fE5ADVP0BmdSlKQRJkmVnD9
z9X42/RpsecXsu4VZBE4tE2Oo0024Y/EC5JjecpF/vSFTWEx+bLj7vcGp3tP600r
hY6W6buXR6rw+aqzogsZGaOu/gy0j3VKiNUPebhvAqcMsnT1yPv02vHjEx/ul1AJ
M5sUzqaxGpDr5wH30JB8whqQXicYMVTjHK5zYT7/uWHsr5e3dUBXI5FxlZhvlySp
yJRsOWx616s+e0QQfnd7nhmIkVROJyATx/SBo/BvjN4xxylUe/lAwjO9MO9aawNA
fQRZXsTncjKEYYGUBjCB2xsXaK7D0koGY6ZvMFUi8Qy5BOQsdrol6+hw18/hyTUg
ZxX9a1lgVKtcSNvMZwG9+VBAdpi2j61lfD/DxLWB+XJidxRgltzXFgeiJappR8NB
QyZsyqa1vD4EWIFnBPgPfhoHCXo8dbdzAzs2k5Kyznd9T8g1F9b+g1CgTDGRIISu
kZy3su6FTaTivdnXMruznl18UAUe093BqQeoynuVQ6PcClP3AMYr9Jmcni/1xi5G
3pIp/0LkkLdbkAP3iyIsoQh8WTKcugUiyNZxFrRiBII=
`protect END_PROTECTED
