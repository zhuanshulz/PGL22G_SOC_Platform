`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/2UmuGkblqQZrzpLTbBI35I2TxPijDJ4oWm4WLJUyn7qyd92mEGSBZmWY/Ez7IXw
R/qkU5iZOBfvvApHEifdRcpgJp2hljW03yOflDgFqIEJpbhj1gFGD27eW1buhTZ4
iHulAosfAQ8voM1hm3FlrzMGTrygSoxfMdkQO2x0dA3n2cAOHLLsWh753ePKnCGs
XRoCy5pHx25ugJwysl7KqUSi2TuLgzbJALsheov+Evk2wyfvtMJXD+xlIc58Ciit
9l92elw5idSgYcfhmV7rwOkcDQN72Emwekrdf8wsTOad2aGCbs4d8JSwjj0Drl3q
JLAxy+4puyiL78ah/Mindcrucq+cY4RaXOtFFao6V/8mzC2isqDqEY6wS7lu97Kk
eIvgTzP1VtFDtT+fqUAPlA==
`protect END_PROTECTED
