`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tkW4AeEwL3wMtwm7wIwtwkyY+CNsCocdPVLX6ycbqybwTKei4aZUUbOTm3zpjoHr
rAp2miM8u054FHXxA6Uej7rxq7Hnvo8deBgAK408CrxCbC79FAYp2bjC+N7Y2Y+Z
dNEdw23WOh8gvwpwzHWOxj2Dlz6bVX2oSltBM6SWBBKpISZvBcCpecHqU60XRwon
zS56HzA5CliaGhyzFvj18No7ae1yG9GU+Ou5rTp8XQlFdbuhqYTqhAW2zQjikQ61
CYavMM6Y9Iwunl7E5XNdP9tE2N2ZxfFLWrtEpFZDnURW/evIAK+Fu4RPAit2EfbO
PMQfS+jwC6UsBX5ju4/8AJzQtb1Jx/+kZx+9nUIrpqCWKxkO4ityLRAUrCU1tNOy
jeIYnvZ58gQUyY5Z0GD9TCrRwxIBgwkLgHX7PUFaB41TQyi+DgwvLTgJ847RQVpC
zJNauhBX9fZKByV3259QxWlv2uPQeyqxcn2+gWSOuQw3IgI6/IvRvpzajjHNwit7
zFHxPGQk4ITRwxZZWDVpsGKopoQ1Dtn82mwHWbZE0e/vWW0ctSOM4qQd7o9HDMmr
vQkZZzcDTnc404/OS2jPLmowpOJeYu9AOklhEtpDv7gccihNmoDvqvPkjugY/zxa
ZrcECXIGiWF5RpnudimGlaEH+gh6nz1tXWWVO2XR90L2KPIPXlkjJJmIVY/+qLe5
dWZDD6Tu6EguH7elrQKK8bEpO1BSN51KUdjQnhhbHbIPFAiybf2ee8nio/KUfuj5
PlkF+BTCawsl2ZXMG2/9jg3CEnMg+onCKVsn4riGlNFipTX/2N9mwlJC4j5n/d+r
`protect END_PROTECTED
