`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3T1ul9cJWdLTZYiIDGqS/KhPIgdBT3IHi3t7d5H7pzF1QuG+tICIT6muOmcNcmon
BUSxvDA4t4gJSjjnM3otiI759tKgzmC+ypsJFngRu+Ob56978QIk45o2368o21uv
h+DnsK+35NaQ8Lxu2jYWKldMjCrRoYQqlr1zIFDVYAWuwFRqKXZzFE4wjKCXGPhF
UD22nAvDypl/M4aQV/DRuQomtyzY0+1FTF/i9+ig3JSgUSM22w4v6F7viuoo5hm7
oBWfmyBhwLZMiKnzRsBoDFSsutDq7fPlD6DfQquwp0i9Olkwd6GejQ5NRoeqn1jb
OXhfz0iNofgdzluRVOacDwNUoeuuKvL5FGOPTnJudtS5asfAovM9Kxwdo1hmyKo4
wEt5X/ceAmvmGcN7HcrOwuRPWlIoQeuOI7hGkxF57CwpWdrYVqP/mcd2be+SycvC
ORf8uFIhXSz0GFU3wh97E2HMsJ5tUOBnfOnBMlbmOjmd0AQw9o9Zr3VmE9bbPt6H
Wc4BMLo8GHkv3oz3g6t3PdmQvlTNHzIiz6ZnwerMxAsMo7qxYfjHLtoHV21dO20/
gmGx66Ana2x0aAR413wRXfeGDpl52AVRQg2k+Jy+f7WA1SONZV1YCsTh42O3cesp
RwvZUkW/H4ZPCnEZvZq7GcNwrDLx82H+53N4TFfvVpeYfZs4e9D+FTZKhQQ2CRMP
sal1YPbpjdtab6drasdTddIkmlO7EwVpYkHOnizo0Sdi6Its04Du5P4n+VBCrwNP
m84BepOBa/BlpF2AA+XVBpdwJ9YbJAmR32u4ULAqSH3ZL3zQppDD4luVRjdsaZU2
IvVdSzEML54onyHX2u+Ia2HIEF462HKcCNXoTZPQLdCJvLJ7b8HnfCg/cu/88vQc
FmfUTPxGf0+O0XoYwDIGb9HrO7UYOs7QXhR4JViVp0+1+f9nHLVLZKsT8L5m3hEb
NljsTGsKB4nTqh38m9QDeh9kw8ux8OLZhihu+vcAStPJSQWXBKL6t1kjWeEWaFHx
s5TJJOaDdl+YQl0eTwoIT0tgK5bxUcofTcybQ1G/WAL48C1noftJ8q0q2c514+Vh
BR+eqJz56U1B+fDyycjMdZ1LEewTshDif28ssTNCIGevbfg8WY34ln3UX7Mkl1iB
sqMm+lCZx0lNQiFUSTPw3wKWKnensQEOAyohNtP22uqNrKkfm64OW+HJbIM/fHLo
csgB9Bp8t6tF4U8YBHJPrrgAhlGr0uTIXnGFkFXwWxzTonleP8/uoP8mMfeoS/XJ
d1qBGLNg6u8s8iOuSQTavzfIvx+p27ItXSGSyXmX3BgDV/cTodqKz3Vcg9qKjZ/m
1oiAZyNWjJKqTAtTt+AfuN8A/iRyxCdLRNjEVRtYqw/RlOliHWTsQcrsiAcISZyC
ymkdsA17jsiHW/BLQCIpP/iKjmRwBZW2WXFNMydgtpcWu7owwfdX3dyF1vdrDL1B
/UQXCdIEflUtIF+gwzJlwxECyZEYGF02MwuvpTZ/20Tns9sWNvyRzUVE6OiUTsDF
DQhF5BqTrLaIbLproaX+3mh6nCaFTBClQoqOAJXeFmFMQt11YeC6/W/AS0oyEfbS
eYPhIpmIWhRyVd/5Qdvfa9jiZLihJzuz9l8P0nZ5ISNqipI5JDRSU5ROVqDlnh4n
o63NvvuM1pMwsidsJb5nsB+RQotVLCHfBv1Ob9PF4bBEIJ6510diIPa5GGFVpmfM
6c8cvEdZzFSj+NW0PyiAABkzd6kr4ImYFmWKM+dgh5mX7ta9PQL6X8JuRVd/InFz
ynATMLOoLY0U19XbvDpVHxLnK7JPn8OiIO9qrfPbd8j2cO3uoVv/eLz/48hjsjKH
GWVMH6VWIwb0qD3K3Un4EDyximSXHsCjRuf8ni9ajyj4luO0EwSUAxPRbBb29vaT
OwOGxsI9RuBm3DKXemVnAHBt3O+UuiR9jmHLsH42w7taJMmgMt8bzeG8EX/uHPha
HTq85atffJ5oqWXgCGU1z/ZTPlAFBQVgg5uykbxjOPOqyhMOZdiP06Z5U7vK2BBj
EbdPN72YPrCHdIN4oWW9Jtej7DiiHj4N5qXRU1Yl2HChkyimwz4fJlpp3rO7pNxl
pU0ANoHfdWW4glA7dYXpSbbI3acXB9yzJLp4/jZPXRKP0ly3q72MUVMYM5JXzzA+
VocuH0mattggeQ80S6Sc4TGJLdMhesFYJEG4sp7qkq/Y+UvjyjXlpZhuBCs0akCM
MpLaBzHsKKcmqrbwryXmGD3OUPZzS8RLWXnRGG569kwMontHzheNDg7ZWbJn4tQo
UpR/sRi3k/M3OEX812Fq5I1mwiDKyDCeHoRA8DkVIGSI9AX2qF+NbYrqv5SYBZGu
A7mjLgAM/pAEvW4vjMP9MrEqq1XxbsiNDN6lHRm0qdXrJ4KlbbuwjNnDQs+v90c1
tMXYT3fZiOURhTWg7+8C1BQxgByiyIVWSXEoKg/lVjOcAOPBLYjvujQkjW3hCK5h
yN0izUoP02SqRanLBvDszkUBq16X7/f4lpvU16TnD8VOvtlq3nC+cMjdt6u+7KsA
sLpkkDRHeRvSPKMRPZIdl/qYflApmZPGRodJmMiheGCrwZq5HRKNa7V2Wx0Fx/NZ
+5gqM6iQw36jVpj+ZQHAdOHDe7zasUkwAXd5RVkg+j40Dr0UvT5B/twoqGnAq1Rw
1Vun0JO02QyWnLD3+YNw3/WTcmd+Z3/DQ7J65KHOaSPhuagFnUyCKh+0QR1p81UJ
GhgI6ooiNAP/8eZyNCHU+hCH6w/9sPCOe+OvOj0yaFeIU8F5oGzEc4iQkrn5xM+D
3KmzTx4zaA90gRZfbWcUOicMcF0ZMbPudZuQZlCmoN5vs+fHG0gImQKUmQqXdGCA
E0+YuImSuOSW4nKY2FBu6TZIDsBeWGKLaKKkO+ThLtiycjY6O2VYSu21txPHP9RR
8Vm7a4IVVfAf+s6yLd5qNkTyp2WKwnkM6zcqenFyzaBYmLQjZUrYtcDKlTVnapuK
2GYdwaH9d59E4034gJpk2nnYQ+pVNpxbipdQcuMdIBy8+fL93a2JQ+xB8t5EVgbl
DuA304c5uAly6V2r4HrTTVICl0yzcJ53oJmBFmopS6av+uDnWc5ve4AJk5gtCtI7
/GoeLGercLWLeG24brtmkKQdKZ5OipP5IsRebBv3J3K2Y0j+LPCpwAKdg52BxVWR
nINGKDM/9V3VDBmSO4MsEdoK7sDTjYtOkO09eS1pihj4v/9TFPuZERKv1WGwxuLI
udRvOPg6folMtMCkfTxmdj3NrjY+vS0I+BJmpoKB/F7cbalvFcJDYRRJ08VUOobg
G7oyEOT0/sgqpzrjNszoXej8yUO6uGjZqFlZgPP9XfV31hK76SJHxaLun8nZBmtx
WmxH4eyMfcBIlAMe/d0Yg2Kg0/719gG4mE8e+JlSEYzEYjRqp/DnxGMu/qdIULy5
1EdVnazrn9b29j1qESl/Lm4gARcdkOIsSTylcSYPWXSKOPEuoyKWNPse0eaGUKs/
3p80CTMlbxxNi1gN5pPNA27nuWOgDSAuV4wobsAljz59NlcSCMUB09ZeQt2IhWit
0Rzvi67sbxW5SPiEg1hY3/sz1V/nVEIvFSaImljDDGsMJmExjJDO6bT0WWhxhk9z
gK4BEdPgXD0YMwpSX9jMOL0eLsLi0NVjzq43rG1gJosT33Ul7Rw/cO1hc20YEijy
oWHUtKBM7r0psv03/BlAinD2Jo20In6kJf+7iS6kQe1ySVVBjeY/e8UVj0Et633R
Qq4ntQkbHNqd77dZwKutyL/hIftM5O3RIXYW4Lei09BYUz9x9EsGqzbyRkUC3hmW
irBYE8y9yRjVxoW/HLN0/p+xz6Cp1j5nNfjJgjv8/SyTTCf3LbwhWA0hrbu0RxB5
rZLHd+962kn1hp/WvcgFeFWc+YMRD4JZLgvzlLJRhn9l4mVrSZXDmgxtNDZzPoKY
H5YnQjpDXXzMZEqSdk5VmLrq9KPjZhPNG3x/eMStlSZK+RlFuGJ/GnxOV6nNwIUH
H698yzSruBHHHfKTkLTgncFaySFf+wugzOaU/oUxptBZzDO55rqbzjBnRRkc01xP
PbMPMJmks2flDiKTGSE9wyciZEs8Sn3FBjybn2ksTJ+6T8T5On4Z/RAUaI36o0jk
PmQsCjQhs+3t3W92Op5Fw751j4ItDX/U6pMIR10sBsFz40s9VUBn6viIOMKvIPao
lroW0xQfc4AjS3gcPtG/oo8fQ2GNCZcMPFo9E3N9E/vDIjmkET2zhw5NDJ74MOny
q2NrA62kuXiW2xgQN4aCe3zroM0JqX7i1/YnupSYydBIyK/f+2Y3kwIymTWtVuI8
g1hnjmfAq56lciObkduT3WbHeTMcZNmpYWUH+Ei+u0lLUECWglIrod+7iwYS6pfj
72YY8xFfPyxc9mY+Y48MKSUnXCiT9wJk15aprtkV0Qww0AoYMoi9/RjZvJzLOgv/
M4kP09CUKzbLosXjXsdzmhV2swkgNSM42EFQIuZnhx2ECs54Lz6A+dNShxJnjWlH
19EjFrC/VHgXUPtyiWluL4gg24NSNfdfl9B82c/aw2fQ6OOwtK34FRxkU22uVqRx
t7L9z891CpbzSzhkQ5w47qvV/BEUwuyekcf+EX4v4adjPKp5dX9lAT+8n54KHcii
7A2YGJBE0faGQD+5mGoXQvatkKU5kBPP2ucDhSsBgBemiKh4sRlMH+0fYQGQw5Zp
msRJ1A0L1OSYkoVlxKKTFYUklBYcwR5gN46xNvgWIgWEoaa1cG1SWjrs6xFNNDC9
5ITuVzfVmn614A2qsVXpvCGlS2tVh/m5HgWAeVlsENw6cuyeIEyauQIsmXHZPjQp
Fm/pC9dtCt1PcVqOjcZfg2Y9FR8zpSbfHYeRgM3VyqugvjZp5Jcb/otgebxH/k+A
ejfvHVvwyf8zboiwKnEGLgA+bvopR6PHg+JFeEe/CRiOR74Qdjf4NZY8kp7oOrm9
pECeB7HN+/paK21zLH72e+tn1mJ8lFAkjn0o3v5F3gDHLqmMiZty+ruWxBKkZOYG
ehPapOT1f2GscdITDFZdUVp6wgO+y5tG8j9ooZbn1Rjm5NCtykQRj8tJWhKyhysl
kSNBkir2cqveAD0tn/YI/T3Ep9InMJY4le7ogLJLwOEsNcUbyAlNwxz3PTyfvBWG
HiKNZUAEY1P0gIMvXBa3j6FEqmNaDIsaQNOIZfYrOvGG2Tmyv7vIkLKP6qJg9CGj
TxwgzY2Bde/yWayDyhqfz7+FG98ntqpjBE4Gjv/H8IovGcvAYLyP6pUO7DNg7ZBz
2JB+x9+DQGLhFgSlPKaXuWIHIGu+26mGNZ7NGgypBpJjJqq83zHZ+4SX0jJtgafp
N4c44R2BM/9/9lkBtZGopORSB9yRkn7S8ixOMIy2g/EP4J/KmWSOa7uFdCKOSuBU
nm8zU1gTcTmn+lJdv4MBm6eQXro4PGw/Dot2QHPm40dvvXB3JMgIh2EjBv8UKgBG
cVy9i9xsafGezA6Z4LqumTW5+7OtbNMPpYyVRcUc2KawFteOdprWyb7NHkLXp4ZG
ODsP8SVnxSY4WC90oRQFhLBEEUiRaeLt2XfWr17gEA7VbxM/KqZHfStMfXNeJ6WV
d6Bea5cwhHvJ6QiMSMkeOGyQJnlsitFTLh7AqdD0srHpApfst/cxAlI/cPk58h7V
iJAd0hoS1anaEKeU8CM357nUDJ5/fIwzxb52AUBKdHIjzw44SkaiOVMmMTWrDcJX
vGOwhIzcDeMkJss776H3+Bc/nCuFah/x7jJNH7S/VpdsnnMguWObocKULo07BYIQ
2cfWZtteq3CtauN8DH//EQv9oX+qbwtI3U4bJyxXrFrt3++ZAuYPHjjJO6rdh94S
HT+i+cJmK2IHtm43Yax+Awt94c4Ho/gSu55EYR9Hs/2BlCVfht9OssrJwmZFDBzS
VXn9nZ9/l/4KyNdxd1RaEofhmwkODo/gl4L/rmr4c2+H++MHdFYsryyeibxiL8oy
6CjlVY4vMVkCXgDCmQ/WLd6QrpezrVhwBKVBtZgCxAd/3QbokQ9Jkfkbe3yj7HoQ
P6CH2EmEhr2NrUUt7khfkNhIJXGqjFq1A6fOOoTZuTAhBi7h8iR/JvCR6MUDjpQB
87n+IGxpdghgcfg+9lTBYQ2eTQg3/C0RDdyCd2WszFJSA+yEg9xtwx/Tfdtcvczq
5ox0gEryQppZ3qVSP5+hCwBwiPQH/bkrcCBZEPN0n2OQRmW9Winm21tQ5Gn2Heax
HCjQfu12Lbqb/zg+pOLtwIBx6oi1sHb2DOWeM9avHUkg6N5ptx+IZKh86zuOkGS4
oyj+PkmZUwz7Af4q+5gcQ9MQ/lyqPW9nDwDvffQm/v2Hf6dFqtZy1Rb8FVL0YjYx
gZF8pXOuX07JsBB4NLNEShHhUJK9VuIltIc1PNQfuTAFB65VUTuz4/fexdAEf5Dy
koyYfvmEWtZfSdLkda//F7vQlgsXHG6IqLlFszUPrt8POjwER200TfvjNpChbj6F
cqimwiHFqBYuJne5rv1YCIJjdnXX4ufht2xz6emd095T4cgV4ETeKA7ihOCQUUVa
iLepSqwgdUL2P4vxy/zHDeVM61IEVhxWoLzoi1NlgqgLwGeel67Mro/KFXNfU9Sw
p4cEHwVMeBR/ovmf53o93wGCm2ofM2Dbf0L3sVLQd8V7Z4AUv3yPmmBsREUUFRpU
tI4lBf+2WJGPZtc0nOgGgrNs6ovT9PKvG7FSNkWUX5IsPsT6tfgrqmjAB8hI70F6
JbW8InBKdTMtqZAoPzSvy5De5V0XWUNTNYzA878zEXIJkJuI9CzEPjmjlSoJv2f7
WWCUVHflnJkj3LkAYpsCYcfBEL15GkiTohZMk9SNoVY1IwEEGMGkxhuFv/CYdK/+
yYnBQ+hjFvbnlM+KkKuVvrXsB+lWhT2DItz4WUYeN+aTFJ0Wj0gvlJvvjvw62T5f
LOTTfChNuLARqaF7pCmNksJQ9LTcGul2iPFcDTipZZ3PDaOw1OleP3k4xT2A1Fhy
rAbqKaZFWE7gi3s397YmLPKvx2JGuCsctUYy5KjHRm7AurVSgSqM+yRHuOzJnQDK
kITPWg03c1B8kjVa9ZWP/8hCjBMY2E4gAtCOF6iJzMqiFFwAyPJBhtwrxXPOW5JU
BsgnxFgdhJxTW9h21OKOLuFq8OQfJVeZ+muLswNbm4buL5EFx4dpa7kle2WkxzrH
UjKWTHCWwnPFM7vjr17bCfeMOpuWZqfbcasgJOX6fw3uJo/tpKGgHhVy4Lk2Nxw0
lbh21xr9a9+TqsIYdVeAjMhZPVh2aYSmlqFEPfrPbgYOFqrfAMJwR/7W9oKEPb2k
6UY6MQWFY1G+UXMzphmFZ+oA+tXxL03j3nWiT9ZaBkFQvbPgeq4ow8y+V0Vi0erM
ipNBv1YAA8AbGOUoLQhSn+j8vmTArzqfWBJwIuPOhkqrjElqcF8oynzbmWa6W+7y
rEsNiYAs00Jac+Jg7nLHi+o/+nqwcrAdNXBbxp6DNz99P+g6gpCzk2Y2+HBNMBWy
u9OUedACx1DZBJRgM9lF6doHPU5p9IUDCgyIef9DzDZlbhdafya5PPVIcp41OrhP
Iz3Pd35REI7Va8W9tjkEJBCWP3zydEcFyk7k7g1ESJpCktu2/Vr3K96+nq6uQF86
ib3P/pkqGlDTkRtg+HIgXE3d0EM9x0lKc0Yz4ZjzrhRDQcuY5REOV4J1AZlgKUaT
D8tsKyhHmFcHR2ffQ6xOc4Xrfn6G0gC0jYFIPTrv41P3nKnsb+ehH5Zrx0OgHZNd
vfmlo1/A3xgKbPt468fv4ONVdXBG8HtcVEvlqhf2ADcRJncEJsmW7AVYvZvkt4em
SGl2DlJc8f2orQsCql2oKp783J8LcbrQ5zKJs2Ys6CRzJ6rJWcIf2lPK8Dhcq3xB
X9LfSjEDleMi41faZ1jsFH2preRGWoHzhquyhTthQTFGQiHAgTY9utsxvXaMF3O2
O4GOK6n0e6LjiUyTSB790MtoGNYxf5q6HLQKfHHgl/0TAJUrh1QLs+TpJMpKM8WM
wVet89v2CtfPwkSYIYBbt0t3z3jA/Wts3ueLaEtenj2lAlxDVCYWDmAzHp+3kiI3
J9bRI0GVEqsnLcAUj7PtC2H/7wL49bzXQ2E3Eo+e5mrj+pHh5fvNOjwBv9eCm/X/
Qg0mocsbti7oSUYNRCMebd9PN7QZZu7QohWegYUib2ZJHG8//fCxjawMGEOkiTeE
Pim1EhhTYblAMaJ8w2Q7SYBcW9S2Mj9DywCOEtUzbylXuKRYnu+yTs1nyd80i8qb
wr4r9lXF/MxoqGML9ih8gMoqHtFKAsC6Xo1aYcPLfR0QC5T1815Zs7lC4ae3xHdX
Iy0OsCABkvN6yV0iLnH2eEV0gPpQP7by196V1UBE8RqJ4XfXAY928LSqjsI9F9GM
z9CuGF6CSyzI4TKujIlJE8kZzgCbZQooAOqOpcqAvabQlq58V8n3OWkXLZiiiPrt
4ADWnqeGmYWfR+BNQKqi9NkF6PIM+oofmz0Gr2GzL7rcTCLXgRi8VWh5QDmPrrfj
E/kqX4lZJOIisdg7vzcsVV1mOa1A1zYwbCyzSLh7sBOgBzEhaoFu6iJonHGdRvqJ
KgkQ9mhI+jiLZY4MlyHsVw10TCkUqH+PzHE/76r+68Nxt4/Q9bZExL2JQR60HyxA
LGDn6lvnMVzZD5HKya7dy+tqAYhXNQDJ8D8flOlF54rZl8EKfhIq4aP2bSOB1NRg
UGpOJDyzs21ISMCMHyRRlOchgntAr7/c90s3CxObfbHcyz0IeTAmzgne958ddNhR
3QIg5UN/5fEyf7ss1DPP+eaH7TPITwAOtPkddlmD1cNudoXAtNs2+QhNMez6GJmA
uoiXsABySHN/nw9B5L5uOI0fYPeCrOqMnnXPE+2ll+q3F2L/pc1OvOPSuEPxU1aC
1YmvY81GC12XYVTSAl638PrwHUF/m/0kRRHq3MGdh6gX1+VSbnfAI9T29cqjoUcs
FtPmT3/ARGpXUwHYIkBZqJOmpkCndQWAzndDV1AEHS1jVd/hcGfoRzK24jWaw2TR
X3dHcv0GW/b+hRfsPDpJkXv7ReCuwEAVkEj06xJOwOQZMr6uZjxzLs0l7Q0YjY43
hrk4cO6JCD6affKg4N63IjrQurL6n2XzMuIqylb46K0QAGXZDcPhm3rS6t1r9g/X
xme/gy0B6WU2Xrb4FQ+56w0kjQ6qysFyE/gJjznIGB3XgM2iXDmL9mU9/VDKanlO
40mHkXDQnwV6Ca3y5Clq/AVVfmEoTwpeaP7fv3X9BRQueyMg3VU/iI+nrGcOSg9v
GgWv3N70zEc0xBwgJE21PGiGDhZpsLlscn+ki3qx4v9Qyo7jagDcceCU/ZB1xtd5
TVw1io6NIbfXSYxNjpdOqht7bddAe20jknnGh2uQ99hrOAKPy2IgINYMnQs22OIt
oOiZCg/YVg4UlKcE2jccTFsNIKZpU7paDo1frusTFiZETtIU9NDYChBabkkVVi7n
ObKpF+N/8kkR7qNqTKsJoIgbDxj8k+EIUIexCx0oTNLTc5wrK7N8Bz6kLiGE6G2h
1+3+I0elHoU/66dblodNaZJHKDvZJjhsG+G6G7N+xfjj7c+4C6IdGCFb6SdGxXpA
uOXJXq73sWTUge/lcnVuAViu3uf17CpR/EPQQTYZXFDK2giHIDgOLQhUbgHF5hBo
hWA/RQYSo65VhmEA9CiTyC2/GEMLy6VpvzUqHm3ikpDB7AvGX64AGA+JecUN1Nl7
0aJj18PloMT7HczyttW72Tvow5fYWaiflCFJk37RaXB4MNLEw6su+HL5wQo4nrUW
ylm/ESoEVLvZOyqiF4OjYL1RnMWup4PfOpiuXu4ZsmxQa+/lYOrB/smtOVabKHZA
TZlKOMuuWHYLkNUfUsjrnwABrlYUvwotqPbtoOXt7QTxyoiYyYuN+AWPSRXNIlIo
jVzx3p+jsNKvWSXirgD+CDXajDmmiE7Uhg6ZHIu6kUvgsUZC8DrWtgpUB/1sK4JA
H5dy9ceKTN0BaYrBoZA587hZR7O80Qj6hQO/MWnc+4o4Pi+a6V8DIl8DI/0ljUbS
9Ia/H5MFMXe8z/54Bj3OStwlQzpRrYI1cHU6V8xUAssGXsCGwUggUWmqwJsMRjVM
7ddRj6ZPRDkD/Koqa7HSjQ==
`protect END_PROTECTED
