`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
83FwrFRr9c8hN3jfbDABL9JO6zTEzkIlWlkMYCk+5eOZV4G18ubc5pquNPQiaALR
I7XXUJRRRDXv1KjEK66PcExXxGQauWYR6+IQPE8X/wVv37F1c8cKfcTz3ctq5UG3
dwOWuI6dQSocsrns6bQN7jIgK/IzXOoepj2y/HRew8F4yKotHcYZxuxj1w0EvodN
3S8BUJEJ2Fmbz+WL9IKW/kSIctcA2jb+dzYRpqN3JNx3JIcAXXb6I2pBkF6vl/z8
IOECXot3aULMx7l8pZd8VZ9Fx9ff7heTkROhn3aNIUw/K7D/n1dAUvoDaIsWc4mo
CLaJiV8R/NzZ0pouAIWZ5dfX8zQ5o55kpSrUBhf4JxEt2KHcaanNAR+Ov2CBHMQX
jJ/f7bePro+GNYStrsGLdCAjMbjH5zjKWRwTEYcOUtwX7VGljuf1Kyf5IXeQIxmY
PynWwkQqZdO0S5WFMLc1eWA4QyV6ryp0SAblaGp1s4hEVgIrYpkAbhrrb1kVBB3E
M5BJ1Fl0cHaHU2rcV+k5tF0yYBxoc1fR0KEm5mNObHX3VjiUidTaW5LpSG5WhUOe
6iMN1WFZwHmZXg2KMF/JU6FT24xTyYqIRqdpU8O0cSt4O1zBI9L7BvPSbAcjL0dv
lAWEdSh+ucoI51kqNjDZ/33/NeOeTh2eJcHNcyyyVvRgXQltP1MzfBP3YaZxOgFy
KgUVzRldL+Ec/EMweojNqO8payHSGCpVTOQYxFaPU5eZ6wJhHKyMEbAOS0Katpl3
J5rfQ6nbaVY3i++iOPQZIu8NMvar1nSdg8onuQaIuS4FcZR3HrXMR7Ask+kJKMxi
HOHVmbTchY9jNb/FL3te/1auR14ecRRbgG7uuuGFwvB+EWsVXi+DCO127gDaAi8U
z8fvjBxQMCh+csdXZwnCLVh6etk9pMVu6SZrTL7JQeDIW8QJjAyTQCOHqtOU+pLK
7AIO1He0wrBnu3nRrWa1PVzbvBzv8myB41O5kYCwhBsAgSFgB5t9ifQzw8ukfIPp
CpexGhBJOZxJ+T98cQy4/SMxe+5sZxet2ZTZiGERHkEP3a6lpYPzjH4Aahg+re1N
c9zq7PNgCj2EkSrwMccqVC+luS3nvjN9VDmaveCeofYN2e5VT0SRHIJBSNleJI1Z
jUNEleXihDKKFkbmY4bdbM+1joQC4aShgqoUKrcPoaA1h13+dEILiwFz+PZid0P0
nPFucrc80NviP1mdkYPtIU8962wrouc52LkYqfySxbBvcG3dEjPp3N7DzITeqQ3I
ZlbiG8SbvtMXsYmFe2Ieaefwo6DvVTf+VEfSh3t/CJ1u5rZhWLDSSAwksYyGvrGO
GF/IDktvI/8Qr4mjnytk4GanHHNU9P6NZkPwx+JOZc83rxCgJg8TtrkxujJbN2xK
UQSxn0eEa99Cr8zuheO9tkj28Qn/q2uilsBrYfKkI0bntYOZJhi6n//KxVAMq+tQ
Lzmh/AL6q1D8j7r9JqRRGgnSWGL/LCSnXGHPmTwEZ4YphVb94/cIhqeJX45qBBUi
s+qfJpIJLoGkTLr3puESrc2u8FnOCTuLa6sPFE5cjpeXEFy2e9M2OVdbao6/Movp
WH2FR/rmqcvpzBWOpwOW3rnM8Ih96l2v4dhu0I4HBDutEySegif91EZpCOIr4q94
gcmAxiFAFO7sOfjBakge2GrSbvH4fsmQhc/hh2E7vP1e9lVOZ0kphC+YvVgTeb3d
AFIPXhj1QbPqa5F5X4zBYGaWabl9PmLYokx4WU9cr2AO70pkiwcnyXPWRzDv+Z+s
tR9crXCzvbLX8vYJro3F8qLKy9CekuYJETP01KPwLhcnr9CSlV29f4KIsSgj/dPb
GSbxlFLDG4b7y+lIloAuDgon8BW3bnM5YoRVB/hx9BVcKXULpVNQmXrgbLRVZz5P
Jfywn4a368AalL5DZNL0vMUrhbhhAr95kJhPYCPbUiBX2KZUHWKN2j10QURUU8fe
pWRdwmLHofS+edcSVJcSd3WdNE5iIKvktWIp9tIDI+SRVSzisB1RcgEsUN6OFV/f
QSLmQOPyRPRBgwMX9yFxmCbDyryongzixjb4bJ0zz4unfMoeyw3/oeHGaVSMZv+U
x+41VmTRJWiESs3HDQwwco7H5AxMKnuDKsaWCkZ36NDMUBKeP8ufyRfO0fodhiy/
nRXfDg7ZZp2drTJpNrh60Y4xiZjDT8IcvRYaXvibH1UugMwACg98lPNTM/1VIslo
L44SebUZnLBXYzPZdGIC5LAnDYB/m/OQps1sNavVqMKIl4XjWhqmuhIqvrikqq8H
oyPJhRgfpO15kmS8lR2kQK7NQPPfzn6L4yqcMwM2g8gps7h81XAQoQbcTKav/tTL
OL/fRXqUvdQYwg1ereupBF4ywzlNVD1FzM+m2msHwMyOxFsIhJWPaoGyBSdxEj15
3qMpuHBvUi7iJWb4DfT1Z8gcx09yDwWHJISUqCny3dZI7tHuT1mpaK0lH+7S2T8d
d78DWQWinLQK+4zZ5Os2tsS9U+CBB+IsipsoNKKOmT0cCV1P4PEKU7U88FOnYlzZ
BGT/bPdRgDGXrl5bcJUwbpnGAQslpgAZhZjCVySFKw/ygVCKvErECmKriZl0qBla
cFRWqwoUG0J1ze4LEIl508Nf7ASzkv6XMoxAxMwp8oM1LsBe3v4CRaCclAfbR6ya
2cMyrnTax5VeraJgRyboHXXrnEvs+hz85EaaPH42bQsuafS8M7tVU64+/KvlKs1P
ogOElhEZOLK5qM250ijFIfh4at0jkTDwKSTmAEY1QM2sj3MsHl/2UzoLm2SH/gUs
DGiZlmETqHn4zaKQKMsac1UpZGQpywuqTDdMAhQJJumop4MdCsgHB0Ow9RPQh6T3
av+jW4+l17Kcwdj6EiykUxrVTSfAndT2DBxiL2Dfi9XWDPO91n0uLiYPP7q3GWUe
5KSnaPuUCzVqDXEm/dmWl8kYlo0o5p0OEnjDIGV6HMq6sNCQ96VzMG4Rzzx7hVRG
ovYs78uDU5zBuPlFHmtxsquSwV20cbDDbsv1WzZ+BoHzVzcKZfqVZYBBqSkQ3PMM
CMhnKlCTymd++LLh7hcrYn7F2qAFHxsSkM/yosq94+qlqkYlj61dcIu5Cv/GHNkC
QjIwQF334J92spwAs7r2p58dXh4xkn/NS3IqIzGaotx94ZDGiYjHZY4XD0kAWQ6d
MSHMT6O8UUgzXs8gmsF4h94H8l6p8Ps7MoBh2xOyC80Os01aoKdVv+RdIkmacXY9
ViEvgUapV28L+SPZmuhTK4p49a/1HO04i9ncP0hCZZUI71hpMzqTG+QwA7SXClDx
fQjN61nT6+jUNV7NLJjNeJvt8uVWTOKHXPq/tUMzzDBCbvyBN8SdtABuu0CY3acx
/WKjy1lMfnDqG2O/avWMvm5Td/8Q3CHXWexdTeVtBOZkG/7qSYg98ORtD+twy9f4
2qgmTdHu1yFcDOVkRGwHBEH9dCooYncXR59ZDACQyWhkuvd6KJWKQNBC2U8em7ru
m05YVQ7V8FyKQafI+49CnCDDRt6LDgXmz7QfLTqnTXDAme6h9NzRhCQUG9jTWCpl
bqVX2fYG9Use4GMZ8E0jcdgUcW6XTNH9juMwDFHiqKPwoxdE/7/p41oS4b1Alyum
tqizx5z4LOf80xP7icdx63ILWyUeikMgr24U5PEX30bse0nX3YIclPZwdSBOwgs1
1/Qt1QGa9s8Qv1L4SpoxrxtLJ9t9dzk38xBmRtutAXEuWVadOFIHCTXmneY8emLb
8SdC3qwniJT9JB3ekEIXFScUOPvi+zaCx78Dgw0xR+jknz1c+VKsAxFBGqvur0Vl
0mR8INcJmnB7SkTHZRpGjwKaJfRx4neRNEwEhOT/xMnF0R/a0NISUQKPIKxdDUW0
swdplzfqfBhrPAdSXsgmtchxWgDxZq808yGu+yV94QpTHRaWlQyLxJDqqrbEMTRd
E3JahaLAlCjt2aK9VosIe5dv2p2cQqkH/MD2+kn3kt3tyhaFeht5IAlFiuqsixbn
5rqp0zhMEQeqBceq1LwbvKhzXGX32q/DdaG4wE7RWk0ji/Yml+yXb+BqBWPB8Bxl
xReF4whYRBtwc1PsTFBArFaaogtRdWQ0UUnzKUOrPV/9JI6DNiJzUh13FIjQZ6GY
g9RE59PPqZmIbiid5PwI3ayUxEHBcPOZC4P/EBZBTlHQ8vc2arukIYOi8xIaWyP4
/jJM+KFVO/L7p5JI3hz2zXnVOjT3L6uaYnOD0yx8Z5dQMMaACZ8JgsAb5TUtq7KS
h7n41d9xoyd51WCvruPz5xT4YH11oblkjUujDg7yx6FOEeX6Uotuab2bFNG6R3wc
+G9nLHKsKyqy3MIx0jx580U5yvowS38x6EQ93hvLJAb7U06Q9oGNr+Ev618rp3Xe
+Yv9aWD7MJqaoXrFfBDefhS1kvLsh1M6aV+og6cq2FzOB7ET+9ZwOaFOZadwkKfe
VPEYSqkbU4eKBRAO3lDK6PbXO0VWNAr0XD/M3lqk4SVgICIwAZHZiKEjF9Ns5Mzp
uCMxtn/Ecyt+6MlEz9WNf1PSyaybbr7KzAagNLnUOyTNKAEWpcZWbNVYobs26vbU
RtiLRFNtQgTKZXE73Gw2VofMvqziOS4pRKLN6DSIhUhHT9m0HE6vjv+kR0v0XmDz
tsR+Ue4Rkw1d06do2mPyH+c4NRD8S2M+oZs8U5L40KyAp666TULTl7v0oAdxzf+1
sSx2qAPGsSwQy5IBF7TFXCDtqd9G1A7LCV8kzxkPCnrYiJxG6U/yisQNmYG55JnB
hlZffo7cW3DVUKl3i3f2/RLYAJFX5/tU6mOIH8hExKRmMfQJxqVfEZTCNulacMoM
zv37eLSObi3nPx/jMDFWp1Cy0UuscWYZhIGz3g6J8c8zd3Xto4WB3i8M3tV9Iwbk
Bow/EK/3UB13Upig9+Q2EfyQMfqdpjXSkz2Mf9n9f0vC2o1T9UGqg05gYzbhLzZr
pK3Q475Kg46xDgWew+qOPhDnpid/advgqGdEJamUi77bQt2785oHGSxZo+OwcX8g
+uqxHRdQ4CrFGoqDGsdzKhDmc8FpqPs5zwHB2I8KggPqzI6smeIFqq0dzRW41Btr
ftbzCYUKMz6RbcCl7OkG9lFsAPmITgSrevR50UdiqgrS0rOR2TPkZqr0JV+MNEf8
SCuV/PRSzMzLMCouu7JeJhi1qFMjtm8IDCmJsbWe04LD9iqWyJCeFzgx+zUMuihq
wZ5HzY9sd6KN7X0DtVHR/qsQ6oo7OyUknzd4AkSe7maLTr3N0IZiaHOHYsRL3aAh
wHloHYIs8rNvjcJ75ailuiI9uxNZ+cHXEv4DTG/kiIk1QsX1iIdQ+3T9vswCYEY5
SAjGxHMRmAMR9cDqQ1RZN7OqsFGySWuCup6cX1f3n9NAz/V6Qj/eIvci9pNP7MY/
t5ym7TkksNCH2Z27c84m0OpFqwrIEV1v+p2L2fhTOoflFivx8RqHK/oOIRhibqy5
xTmYZzU4PPCSk4tFTW/kIbJ36HFMcrfwRSUclxZreWqOII/MtzTxaxPjCufdC6aC
CxeZE6DUEeZ8xJ2NYMEA4j1MnswmvdT+czda9a9fwP/naQBvKkP6o9QDlLVM4jK3
EzBbkO+4LIgHX1nK3oqIFfmwChOLvkIblb7J+FHmXJWitMO3snnTTEDZxvqtyB4b
yBZIfXD5m1qPFUpGyWQsmrqSVBTokiivOtO4tka83tsAg+cYtOh++p9A0kkbFIky
DGN5ZByoGm8OUX/VrDOxa4QuVtIVasUfReOOFwuOZWBhaLDtx03iwBZERIqw/wYJ
7eYXIffSl3FUwIXxHUepUfzhhZc7pPmkjLVnvlv8xVjRiCReKnXZiCHoVNtXni7w
hSNQuzHhURlLvZlWHe7ARGnJqSgeXBgKSsQgZKJ6s9zFZIftAKgfCU+F3Bo6OHgk
NSWQxsqOMLYbKpcZUMGEIjJVbN+ZttbcFOXddit63s9mSW72zY150of8JAUQo1P7
7IGUpf0DRSVTEgjdFSs6/qe0YecWqANadKhxXbl5YEI4VX4jwcotuspn7CO2R+iU
VP6SHJOTVb8A67ULWf2ikTQEb6qEfXCjKapkZAnj6tgmr9yRnurzlgkV20LL/LbA
kWc55TMtltfmj1s/9G6c/kg/HfGwrNdEu95bdC1gu4Qbz26ZiXzAWBedQQFr3Fw7
b9luRViFa7BlOh8iBw6INknkaJzbUt6S9DI9RivHs46nSDaiBdhmf+gZ2hP6275Z
qWs3IK23j65gOA1Y5YsioRL6rvN68Lkceb9MWrX2hVzyj5SxY4O7x+HCjQabB34k
zV7yNQJ+kpaihWpG8TFvvCFf+ccdoCizcAKedyq6df4BXIJO+ax2TVQyUZ7Hd55w
VqNXyq45GuLQG2aJ/pD6c0gxZeeVu3sQAyXGnDW369PwqLTz5M0YrM7UzO+E0HWC
ApMDaAiFXpr/3BK5SZQsewA94LPjK6aoE6P9BRu77Efy9BcGDAq5b1LU7oeDHzq2
7eOGAjYY6iWdkRJtza8eG7Hx8N1dtWov07SIblKGaFRcQS82frzqnaPuX46llOB2
hDKtb35QcMRKZ6yR837BkdcNzaDSCyp51fSmmqW2UcxGCZSM+nIBYxS2bAr2TtR4
46+y+dR2fgSaLweWqYd3gZuHvOFt1uSU8/wQ+4IVQv94twlIAsy8IgPHHDsVWbgz
S73E/SAklulUBq5M+WC9u1ElmT7zLHxgzjG6Hjcdaw0cT0wgxWp88Xv4CP3yzHHi
AiBu2Q8rQcTOUSC9Cdrxg5v4iST6q9HxQW/gTGCamCBSn3SuMqkWQnwBv1cLCROK
LxvN+gAFNBXuVPNSRaWG0zGUzYuMsxZufabu2mdPhxZD0FT1BEEAL2nBuzSxTfZS
6Ogei8TChMUwbeHK5eCQwC7K1AbOgewsWrE9Nc3t213JKJPhK8JXXxioEMludVGl
0jFrKN5ySa7kEdgTeGPaH3WyX0EpzH9DBCQ/6CRZ/tKMfgCKHUpwJAUXoN3fRNHj
EMEDP7+Q1wcQIvABB6G6F4z0Q7Xfkr3rIHayPvNleSVgL5X8rir39IPsvJvieSPZ
S7LdxRuilTlVHK4l/DpyWN1dUUMrb9m0o4Emityc+peo/FYtGOshulqTS8y3Zzms
7WPy07BwKEFiMmsGX4SHvXhj4FrTmSxcNcY6bSOS5NSvO45sKKHaN5M3C/5NyZPU
oIvL3E1sMn/ZDWYYoESWdPtrFMA9XgILoxSSb/sCb+XGbJFlZRzXr1Ijrsup3jC6
G8wOMEgW0Wve2FE6zvK9N3+S5lQuf9Jmjq3ylm6KLpTW5AkVgO9cM7XDcaN0TTwb
NxjApO/H8N+WWk3vNSZwrvYnv3BT071f94hKOtIA8w5TGX1yqzUYNQaQFHzVwE2e
kumKnGDxY0t4aD3C92hR5aoe/oU8hyj3rLd2D1hutNf/E7RADsDnGKSZper7yr9i
d4cI3oH42O7lsWEy34NO8omsuQ7oFGGG19bZP/qKFUFo4ZNVucekuB4m2TehsGFC
zPnw5x5zkDVptgni6PegYGudJVRUfmqXR/TRujvlMmBEGsMxFUxvcOqke7vq64Tl
F7QNxY7cWHVkFDK+cBeT9rqSho0ibixb4wSVVMQGwvv56gi99WB4jSjjn1siuiVZ
dyXQrBcPCcF6wCnYrCwBnS2zvOiReMrnZpA3T1Na/Jt/PDvCWJcr6zpl9HQSc8Zs
bi+PckkotPEMZNT1/cX1fa/TUWOKBIItWz6UZVta/5Y4XC+xQB8gqLjq5qT0zsmr
uPFu4d4lPcg6doon9XIS5Ngd+npRY0+5wZy4bFjZRi+tiIifaTIGW2dGi3nQI8tm
uwPNGhdB1oq5w3KURDWJgva2IkBWRXvzfaMNCQBWLK/IIq25Xf6PCNNQeBw3Nof0
A1cathmJSVokYAY3gwZTRQASMqjQqOIDQBiUwgx5XB9IuNPf1OG7ZemQMCm7XN9N
1UA4SBUI4Yw09+Oe2+B5uNmwy1fUR4AN5OTHhKd15x6pleZAcLZhtlKjHTHuUip0
sY4UtzX62iI4g20zD4ZebiA8tf3tQOIZjT8VMyF/4V3ul+Dw9EcJ85jG+Ep1FJ2j
H/XfBH0BtfYfBGQbuj2mEohvAUfB4I0wMEUufzh53xcPcE7BL/Wppp3kKXVn/nq1
P3rwlSo8qQqKxLQXkFZQeNXrH3Uu4fUDYKKrnNi64+B2W+OUCUxe0/sbG3KxMfz7
Vzf1LGQq31+WVYhgjKEfeGmM9FTvouWwl4QfJ5kvTOVg/HLUZL8h6ZEAMJd/03EC
1lXCfBaOTFGozwN6sVcw7JWlTOSF1tXw94xukdn5DhPghZXHujgLnJ68D3Bmy4PW
1fs+Blst1czElKUgwCrZVr187F4Og+GcG0gBoq7ee/ZyC8/Mkr/2BeAR3xwi0oTx
khPWcF2Xc7dKz6rv7l+sKG7xn5HVfNhiOVz5zeaeFSZggrnsyAylMJBvL+qgxptH
k1q2GhnbgSfIi5K2Gf5/MOVcVbxSU/pl8dUAqkTV5F174EjHgOLKETaGiKh7Ea2W
xmmsc/wdNYgvyUnbMuvvJMKywyYj0x5t7DR9Kvxk8AWn4xW5qyo8l0dtbA4zgLaa
ThmOkqFqGugoSYJ6aYzrKna8OAE3iaMA5Vz7kWfq4YzRpmuD1wqBqRzJuwftG6f5
zSJG4GnW1pkQVAK04oez7zGMy2N2XHWKfctHbRIaqFfMPV4mGgW9jbvoTE3f74NB
h6bdUhns/trAXOds7UHTH4DqMML6HUAM5Sr639mpH13LvsbA+4t2s/DWzuQBgxmr
zNdVt6CqozxPMJwilfiCAiwHMbdKhO9i2MaczmaBVqeqBlz6BYEc6I4r/yyMNtEg
7PvJmYGN0fHEohvbzYEKws6Ae692zSXhU4KTWz8jpa/UHqmAANA4XiBT1fcAt7D7
B1zg1XcbA4e0stFbyh2hugGelyWUeXiC63QzcfMWdaazHunBQVFpPNiWf4vDiUTi
43MjHnADDfnkVtFjxwwP9MQ2rb0+KoKukzfqvV5FN1YzqAHYCfvG8dKzClW7HksT
dcXg9m8UhpEzXut4ktpP3zFm9KBPRde7kAyy/c6HGHJX/fl2BiFnDgDYt1Xe0raP
xGietQyag72cK+MKRKCiHrUrmMuExFxDAC8hMj407MnHxPPTB/hKCyel3C9pepUn
/sarlfyyPguqLSylh2ubth1dvVbBpnGDG24OhtzR7OvEqNAHH5m2d5DnI4foAL79
9PFcGEvuxX+IhhSaqknDiQJbO5Jz3/PMhHWlynEbvOQkfhGFGQTQxjJCgr3jxe8c
td6ykpEIG4PNe93kTkyfFn7ZTtjA6H4MWi8XejmXCKRr9uJGE1rI5n6tiAH54GU3
NC3/WdHdCEnqupZrIPyeWUo5UoG48Xo+GFHp6ciZ2gFHlWJMNsRXiRsza0J6aHJE
ip2Q4ZDvRUgF0FC2mpjcO6nzZO9KsET4j2tzYSaEOzYCkWK1LLCUccYkLA46W8RY
yYG361X9ck/dQKTMNMbXj+TBS3fvjJFtkdlBKTmYOElMBw6LfGMAMkYqWnwyx11H
p4ClV9qOXRhq/mW5AXA9ZyytDSdkWRMtbK09/Uc+IItkt3T2geGA2nI80osh83mo
dsanFxhxIan1wCA0Bf8qoWY3Ie40GvVrDTVJqykX265LA75U8Dfy1OZ1/sU3eowF
Ddgxcm0NEhoDNuC/Tc0XEsMxaPYfZtoHQUylPeQDMSRAlkGPzDDMkySu4cdC25h3
COb7lOZRvUhTuYqWSwK7DsJMioqwW955FwFRhIOgNaPedr3EgwuudVYiJwlI4r3q
e4ZKWiCMnadLeAeR9vdqzWw3Ox445sRy25XqJtd0U0smngwKVoE8o4lqr081HrO6
Ce/a2YIF6GrTU3VeE64KaAVPNRB/FjaCbCpJzI3xhSiGS+oZf4W24oLgpwQhzI8g
XTivEC+CQw2TuC0XZ4RPVAqSAhSzdvSzn7k7LInESchPmxWYieqdqL+stUg4OjB1
sn+hDeKwra9n1MuWW3nhl5osew/QlxaYxi2LePZpcquPc0fFReW7gzWvOHmgv2+G
uXN3pv9USGTXLPgq0CSIRVhMzLHqjnltTQ2XcteATiPV9JnXD3harupYKTSKPAqb
AEUa/0uTMUxOV2GCqoiMCE/+SjjnFZg0C8q5sewT6IVHJscq718RW+oDWx68rqgf
Byvda/wD5IWz/9qY3cPDXx0OinrK3R/hC6oI0TK/pFatBhIV+dsx3VYU03CnVqCQ
NJXkS/WkpchKWlV3Hz9qACUKWLAG+OatycBH/2wNg1snwSl+6+5uY+Qpn3S8Gvhx
2hfPpJb99skCgneq/UBXV1BOGrGgotDP+KmVqSXpJVsjbS1ZZtqCFfgDLR30Ms1k
gVZnmzagtipeiFkW1Q3T7/fkyDdpMmIzPOPdxSGWA9bAGphEfmeoRz4sPsqbi8Hw
yRxY6E4ZrE1IPfrsbutFxb1qMkEGjifC1h3+WQxmiC4SK0gjYa+sKogD3km+XTrW
pb/mF3120Oks+LWqaoLWHgW0DdAJguSU077RhYAXyF6JtQ6JjJTR/vivNNtVWnZt
DqhM6kiAi1k2Jae60sx+Rvgi50PDvH80PwY4WVY4IxRBcb7Y1SaE8FQ1R4+ru8Rt
eI2yBQUMGMYWgAvjYT9dUOWSkpqUiIK2r76pGIMhj5w+Uh/uDyCCjk1rPxttjW8l
pFPMldfmPuyJot5p9vchtNw25LKbf1zZSLMVi7xxZWKMiu7pwPMBNcG/ulSp1aCQ
ijZ5FwFkY/9BiymmnjF+O6pjuVcN876VCtXLRm0h1S8lMiLg58gqv1x9wrJcDy4R
Pk6Ty/qQt/oPLYdIT2oDimSmRJ1AKurS86H9oZQFquV+8tLFipnMUFAasAkCMtA5
X5i4yv87HhsQ/8sceCkdw21Lv8Dl87PUxsZY/XdQbQtRPaW92hTbX4kZTa4WwDxR
2cYQ5UNbC9lqoqXepVjAKH2s3HZhZmP9zJ11BPdExBwxRtzjPUkhTMBoZNmnNYui
3q9TfUhDk/w9ALxwnh2FSGQ8I/2+ZhqcAxy84EiWvaOAcIEWe+JE/SiiPWqHFWaO
fhHXInMQookhfAtvIcEX/nSY8y7+ogH2mV+PNCqPx/RUSyPhxd3Vk8kmyJ7gdJCT
92l80O4mUD5R7T3ztyaimf5eMxyVaMA5DhR/Ije3I+8WnG9xeKQUfmgiM02f+V5t
yxH+x6iZBCRwUPWHYDPZs6krcSzErk2zWgVdlLEo8PhTtHowMZ5nQb2ADtqlyExX
r6CWu/uDQJhd90NYXOMRbLpOLktmKE6eEflQ3TMQDcUX3tNbQOQxymrRGfBP5eCA
Ofd4czu1RovkaReKAGnbl5f7kJhza6HA+sgnsUjJzkQbyhB0/poMdz1yx5AnzVGN
RjvkXmI0hUtGDddBnckn5yAlkqCyrWLa+Q+mobjRLkinbCgPdEN0P2fgQ7KCevP+
ZLFYFHobJS3JRSui91DL8DZCcufrvpNfgy9mkXXHk1/Y9lQ9pFTYV60fvsqYEFlI
i/gxYapl2MYlz1JbxCL+Hovm8g7XKZ7b8+avL00/66gTU9hvdx/ZVqpKLvGJVIsU
7QDr/wgwdHPwAnqLUGgQPxXMvBGBRp5JPl3Ykfzfd6o2VjN+Avj0GaYtwUkUz8T2
ohJgnS4TxW51GL55O4izI1rujYlerfZ3pAl2pRIJ7FWA0xwla3HoALXG8OF61eF6
g9eRHpaeQIXo0RyMBnzLkwt2BjBUexB6DufNDbe6qwgpLZDbJATopgjN0nqxkv0C
9+oAuZKJfJnd1L++qOdbRxVXIu+4UfnEWzopPT49tRYIyMgXnjfreVCwJyKtr5ac
d5Ddj50c0ckpIxthOxktzXlBUU00V9pEprj95BhfWw5z98GSH+w2AD72Agdk/2XG
4kphFSYzAS2fANcZZmzpbA==
`protect END_PROTECTED
