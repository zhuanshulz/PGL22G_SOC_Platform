`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DBPfMeUCm/JB0Nr+sFi80sWOeAlve1z6IirF7vYxXOWpvL47cZ7tfKYOB8XL7fCQ
eG5//ig+k1QtyTAcXeNORpgxvguI5oY/gvB0FB5Sqftka0Ov/t8kO+sNkU/jfa/G
4mr0yXlSMmDGpqXfLw2i1a/dbRG7SjE4En/7Ye42q+DRQymle6zBz45KwYH5YscG
kkOObur2voycyF6V/bpUJR6z4nLd1MWjqGWemvNAiV35yqJ2wMwk0/DCQiwwADyl
bjFZDgI+KLSWDhwxsO0KOGJWRKGOCB9OAprEv2QrnXPteQYCYeqNz39XFP+fd/hI
I/O2jZRctWOevhYw5/Fpcq8xAbMtoZerg5Of6xYwkjTTBhCHQt6QCmsNFvFUIiX7
0kBLxWTSOPHomT0CISEnqH/EdkByS/ZZIQGaambD+j2qcDgDGXJb6IGBjrNn6KLK
SjGCyh8WdMTRoXBUAhZgjH3Hvv9OvAVbWoI+22JEOiyOOLsh0T9vet26BsgDRZAG
nrtj3CUuLLyUGV5OLt3+lIS4pkhMDlz7QdhZzutfRwbnB/uSwg2LsRP523TW6Evk
z9P7NfLsjk8HsXONQT61VbSIkFSkgGe3b1C3IKztsa0bfpE2m5YAl0sor4B9tIx6
LuRLkG3RJK1vVNwhHXodp0Z5WiGB+Yz2qZ2DXgaCVERa6vfef95K+kyaK7Mc60fV
oEvlXdgM5wJlBna3Ce8ZjHqVsanxTw1bv3OtsO0TkPjtuqJFJ7Bebp7GFdOa6LKy
3nLQIpqZYO8fn4MjxQAKoqo/zGqK/Wfdlp9BZaP/c/xJqWDz83NmFOsgWk8urJT4
D3scW2a/+DEf38tIyX9xT/v3OZY36BlU4UvgkrzNkDDjq3/T3x+KKh3uM0PxGiOh
TXebfg2qM+XwEmbQ2D3loLA40PBkCfbPyrm3ODuFg7dm8COeyndxJeYJ5j7OnJas
gMdoZvBeWvMHW4gcxWQjqUhGFRsaWLeYPVUadq/xc3WdbRmFmz3+L+HJh+WwfFR0
jbwLQfcTRTA3LyYMOtFQnoLmGGdJHRispZ7CqzJsTmCayf92QVgpqo0YQjxmH0Ty
IsHo/O95klYAVE4PYpWaMmlse21xibXuSu/dleuIkTxYVp2t9DHjoSrPVTxIiGLc
OHZI09wNH4LweS1Mgn4xLgNw8BFmgKLEJAavFkrY4Lll8Dqn1mDLEtn9pyqISRYp
TASm05v4Eu4FuSCrwki1fHUh5vANpJzf1R9ENimjxOin5Y+CH7vPqokdYmrcSyUs
j8ibPhMyQkIQEAGMvWS6BWJSr09afc/y4oveHxh7ODV3Gsc0A879gvAhzWdqoZOh
pGzBPbP+1KUZOZUwXUMub3p17wCoYeOthZnZeB4rj/3Qj80UixxqPWazA6Q4k7Sj
z8Pgzqw6zvEs0TeUx7w+1effhDhLpQt8fwCkH7F6Ov7aQoD2Vbc4S8JBDKL5bF1e
ZqrO3yXmH8p32HNIDo6a+D/V8PJ50D3rNq5czoSXoj1F4twI5fpwjJyFM9YWFO8S
sS6DOfxYFFe3XcU1WXdyp43isdFJNm4IWvhSR9A4miXUdOzTVBljBngnkppMsT24
D1wGo5BjQDOXomqHilEG/ECl/dZJryPj6KR93qDykfAH2gMfc+tvE2x78UrWr+ly
bTnFPbRUXeTFpaLnScKOve3PigFdDOGga4+2fEdLPfqwVoAKgNIG87voH3ZrSL7Q
gWOl0MHSSiogvH/d7bH7k2UNLhuF9Dk0cmauM2RiZmmFLQn0kyPvSMMzzacFOhfd
B+QM5ShTtQ2gYzSbadtnfiPuZLcISgukHebYK7MKowHFpYzXfVaJcEoQA0LQLreb
yFhseg2XeHyZPIaxGSKwAmZTFvheqHd08ke+FPqNb7Fxd52Mn8Hs2MWA5FV93vC6
okkHIctjpFLTZFtyquaqaHfCZsIMkT3J3HgNMSQ0gWDXqY++3227TWYizE4qABFJ
dtUKJOJeIOf6iHXpB8UYjoh1Y/cOQYsfqxyX1sBTPn1MjcEP28dLHMEyYU8E9Yl1
cUyhSszfikqGuYM8zd8Am7DMOX166sSFdnl8uiUMWbiDBGcyh72V7ez+zriV98SW
/E6/S8tKMcJ2iPVZm13jk3R99yGpQYlMQKiuNZpEaI+/XY3e2VNgsvKrEsQ4cgnp
c6zHXKu/GgfdaZwwOhh7NJxCe8gwZUK66KYQVOExExQVEGBrJb3W0L7J4UQ8k1fH
scY0/c41UpLw4TXUJZ2u1BZkTRdlvnVB/STtp/OvrHZYiWUCBuG58Eupk6q32U9z
52jnkkwcuSBG+Nyk8INOQklVptkCoW4RwX5uLfpW3/FBumrEK4/NzQL64Pp6zZjl
psxPDSi0NLBlCaPljFpWK2xxy7BnT2G4cW7IkkQCP1H0IAWA9VPjCUY8IuRnqixA
S1B+39WjWQzp2n8OyQiPs8POET2ApZ6cz1dHWcVlHXXUoCXza2UdEspbeh/Hemff
ucwYi7HSYSX3QGAKdU+9QL/u2+bWLNZ4SqPe33hQBhAOaSIhlhhVXNQ212EmpLB6
Vo3xo9UKM6lStSBlBmwMfqZROqIt35WQKAFwEIZuZ3hUIgj+jgsyRIpzclYfZStz
yGE98c117JQs52kB2m2mG5MboZd+W4fN8OthsP7/Vh+sadb4Gk2LpOx12O+naAYq
HRbrn4usZE8rH1Os7/5DRaKYRDH2jTR83lvi75yrFVJjwW8nEQ1HnmpUVrKm11qA
BjXRiPzMrwZxoX2N/vSdAwrMDIy2/2WcvrPgA9azNMs/AqmS+Dyu3vW4Gc510bBM
Y7SGlmjnmY/lT9w2J/W+Lt10YE5E6a1aDxgWHiwUnr7u7lejmyHWuylLGj1dOgvy
BONd+Y99kFR9I2/ZYim2VazAH/vEUjqeluniarltFbnVS6TyPAluzRnEjTGze49s
j2RgvqN1umFIN943UJKsm9kO+Oml8CnnMil2SLzRblOoz2TTpONfPUTEgwh10rkt
BCFesiIcwtoD9htzcBWCIAEl3yC34GTVhtLNYv9KRHuxEOv9OFso8l2FDB/ileKD
Hw7ht9/T54TULCV6AZphdhaqPKKZP6kT6Ilg2ApdW8KOzBaXFiK00Oc9XZyt5orF
nIqzNSvlJlUyfkRCKdleKPhywMtmuKiOzRiTBgsrzRjqRI1Ie+8i0gIEfd5mqPn5
mmPHQVwh6eVaIJbodEKIFPvVP+bDH281/RsrT4rj/5BQGyPlmZCdOjYpjELH3Gw8
FBNQoVGhbIkNS+FDTJ8pUqPe7qQIgBGD1TaYPxvtbVS+2Ad6cOGC7JgArDkoHFpw
qSOH1bnYCpHGuhsgwnkfNqN+mSA0JKtIAg4CKW8rWy3mG3rqxMd+f/gZ7XZF631W
xEwZ3ixAXETg7JjSO7eOCE42LwSPcrHppZhzHTkBgzC7l7hNx+UkKWgrWglrElNR
Ep6mRZ1RMn4ydK4MqMYrjpYnDZAs/8MrDVb7b0Y31r/2QWK77VahDd7A7AgHjM5x
lRNimtyNaymxdoXJQCYIJbTxcvF4UlEQjs+x8H9fFwI8awCMFaXqDdBGce3+v0sb
`protect END_PROTECTED
