`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mDkMvxB3S6OnWI0EwnLUjrWMEsx042iLB+4Kx6iL/cvvx/l0K03GbUkVdA/ENwqN
WhKX+oPk52gb8X+8lbJITKaJaAS+QWMHwtWb6OLP/WVKHQ4fxphtv2a5GD/iDznE
FSyMRtcXIhVXUZ1PptWl8MEtqYYs3tcYyQnZiFRkrSuCfkkBOISSNIdDOSgOnQTW
saz1VFRqwv1RH/kb51jvYP+AoAjdjPx/dIuBHJU207+qPC6pPn8QlD/AEtujHdql
glPVA87/s9hD5VOz64ciUBUFjsHNIokuimFlKfUGgR0fmm9ehbn21IHlC1r2l8bs
LWmHA3KN+jKTv8w2sF7RWvI96x/stPcZ00b9NqH4FnDIRpKK76NT7iJlnJH7TI8d
wqOJT7HcN+Ymk0Sg/Xt01qGa62i0Q5QOLDmvjxxUg1jgC7vGqLyYtYPose0gNbgx
urbaMbtpYRXmLV3Vpq7DO0B1sgfq55xQ3JDz/DFCuFBssoW6IVMtedWyaFtaQgIi
utdN/YX8fSrQRlWFQVfctwtFwbnBBO2JWYTsOdJe75UWSg3ObXKfaV75+P/Uwtbd
Z/e2BIaprSqwLTS+ErCOEgs+eAfmLEU8FuzVwt8KAz1jviVuCX8NkFMcuG6oOPNh
rhomWxO3AXVgP+66cfySF8v3qe3R1NFlj8oMIVs8GnsuhlQutnuP5cYXWPmn+D3z
mii9WUgWhw7y9z75OmJ6CN+ahPJpy54Fz3v5UkXHWb2I+1h74VHWtn/qU8LDg5dS
mEsOqZ8Yu5dYVHmwPl7ttCxtavrtxw3LHnyqlniBW3CEq13H5k2cBGGgEJPYeYgF
Cy/JbWEQ3Ga1nNwwEIxFT37wIT3Jr74PpIGUffaebn/HSf+NTgzyv1oPsaQhwVS0
7E3NLw6MTVqjAhqaIDSPyduvRMz907IIawn3vTmCUBCYV9uE2kRakBSU+PM7cq9Q
ZUBfc3l2LzFWYir7vHHI0U4sbnOqa6mJWu6ipP3rC3E0X5mj9LQiCed+JoLvhcfs
Xu1B4IhC1S8ZkWFbPu5xodVNP2giSxUNoUXZjsczU5BVtcZoNfKJafb5v4ctjLuF
46XmEh4cW1Nj4b2NEq2RHUDCxPbm4PwSvoIE2Bicbtk9m5NTDQspmTwBclmoLbIV
dXK7Q18CgyrjnnS9uWtkQlXI7IG8BylFgnAN8ueVueWwLWzlkKww4iSdkbqTknrL
kMoM6QKcrbhdvUEnSOJnoGjetPspDcZbedwfXMKfM/0+CrfPVAd4dsN4KFyO0CSG
kMW3OpHrayV1hA5knylUqwAZoCShhQ2ELfZ5hCJuPygOp6ElwEYX8UdO+UEaq4Oe
32CSA+o9HiVNytMwY045Rz/PCxA0VhbEy2pfnmblgaRPus3s/CLnPZqPGqSG9iPE
xiEyTZc6jgApYbLGIabxtGEgqk8Ph1Q3BGcpYcsZqug6/Tg7JAKcZgRQgjgGExjs
9SH+j1yiVmaBEocm4p8qRkoc1x4B2uXV3QnX/S3TT3P8dqzspQRC+U+5NI1BxHM3
`protect END_PROTECTED
