`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cFXMui+7/rVwk5c/URilC6uIPeWo7TGPMjE9SPujk63V5uFrJWIJPVW2IdqDyDFu
haRZtshlUmp+5urwF8qZZkcZw1dcHcyMA1l5weh8DTdsi+T4kXZcARRC74AWnzk6
IJXc8R4JiIDscIZ+csy7NxX9Ry6LtoIevUc9p5rCCcTmUGplIH9Y4tbu0y5F/bKE
Ev33lCxLRK1wOP06fppr4moECDmYCL6Rbp0hLtWzoPvbdrmq+M5aROVOuNf2zaJF
aoWUnpCZ21HcupSzTzEU8x8Zmj+PYv04ErtWK1nhieN8HBaelMldobodQK+20fDv
fC4ItEYavbJB73dcyQAfnOWGb6dd/yLbaN8RHWArMEjEqRNBkTLGgI6cXDugcP1q
8BwA01sD+ehFGEH7YYGH+Q2KQiqgrlkoBrOn/Z+AYpfLXNBVM+Sh5Uf9h5nTxXLC
LKYtKw63SemQwhaTypUaXrFTIH09hf1m+yKueeVGCsymF2X6rRfKT5dIcVjGpXVO
19au91DFwB8eufyr+TKPEMpr5vMuSHF4Xa1PMQDB34sFVdNZizAQejVcHDdhNJzv
jKfamHcMTRJA2QF0kSGNxrRYyuGglJU6XPx7/PQvEZycnn3Mf3JGl/p7HGgp5OWn
CN9Ds/WT52QE86yYdNHJ7R661v3CymbHlrBComfS6B5u7oLQhC8KdLp3J4q4uSt+
BDuW9Ot1Yz4SyZosMPeFSO6Nmque1s2c35WX2Yb5+L28xwuVLwndFprIe9bO0kQf
CQ9VTqm4S7isHfFwP1y71aHyRpGi7wlNK+YEVwquTFPTPFeVVbKy1qx4axILCo9e
FthhX0cs/7pax/DiBJTzVzzK4RPDkrXlulW1DqnQbQoLrDGSj41ZYeVMm9IETaZL
rNDHbJ7XFqahuLgeidVjluOnXGiSmDQTVWMD81AaJZdtEVPAMQ4tQIP44oh9M1Jg
Mcdn693Znm3Dl0khOE0mdr3D28jLRdWu83K0jPFDg7eFnc0D3Lqmn9L0H1VDcbmx
VOs2LkAJ1z5iM2oXY8q5MxqWFDTDA/zpc/gGSK8sYFRw5cUw7H0iL/Rw6II2WTy6
M+kjT6zLqpvh4x7djN3jCs8LaS1evGI3zXIx7LiB+QOAqWJ8yW1Ozgw8mYs9IVKH
GmvJrJaAykCXj4vkhemQgJ5jtXXd3p0BbC15vzNZiRo2W5PTT5kXbzGtwkD8y2HM
nYNrCZB+L0leCzjYNq5EZHM5oVttV/wGhVle2HSRU432BlJ4EsfYzlGM+yCEISSk
UYqfloKsn6XSwYbQfSRphB9ghUjhCHQANA2+Z9dnaPDTBwV3vUdnMSHOVP//Y6EX
p0z0jXCmdAz3qk15D1sOhLT+9flPVcOyd5563j8jQ4dnMOMc7IPVU9XsGWV7Ubki
Ipd+V+TS+Dq1ag+QmVKgVj9hxqPvxB1uweS12dwZe08Vvks22TWI1m9zP1yIl18y
EdsEoeteoI3T+UUbXcL9DTmlJEKlPhHSRmnBDcSFV5iAJngqIu+KLal4gvfD4IBe
21cCZw+H9qYQmFhsLnI2qCBLdWZBcsSlTUBQxt0x31pVNB+2Jjr/WfOh3DdEgsmx
FjOceU6FyLIipbHctd72jmCCwnLfRCt3/JLC2zevoAyMFcGCY1wg9P1JhDzCt7fz
sjSVdJ3hgqnAyQS4qRImGTXFNrNKfvgkcb8ONY3CDE27ufaUjQ7quUYOwZv7wzGH
BrgTCdFjuj0y8TWZ4ReTxN9pSZltExGx0Lttm2PZB3IV8IdxJwjJbmqxetwkuH4p
W61ID+2jTaAlRgSvaOjc5u4whJ+CyTt8qHPNQ7B3SZgJBjj5wAO9m2jzchb3PMPz
WdaiYbSD9ZMk82vahc24tQXrFH68Y8t7pydvArHiCunAsZp20IafNocp3sk7B8N0
IhVPP67MzhboFt8R40NmK9ntLn1GxJax2bHgRJ7/KSU3qaUkXmYofGNyfdxr5z1O
LIdj/BQrYf0yB9kFYx+SLYApcRYjd3m08SNcFA8/Y3ObeqxmVYnr+FXkQ0Whmf5o
ixmgogxiB+syYApAbPL17B+rFr6zlXK0p4UQA9X7z+FAhD39K3HB8VUjTTXqWWsn
eLS6TIQ8GUFOPnQ5vu1aMjKux8uIDM+sXnZRQbENAjCsMicHMwn6y8NnBPIDIkx8
EPRoLnYwLdHeM7cDCtcW9iMEPDSfCluQEsevGsPM23JYkPcJN29HhDDNozrY8bcF
IsxDZ3h69c9NC0wKohEg8hLHP5dE7qh3IaCwKwV2gPy6639KGZwiKxUvkWIS+DB/
LyS0zA7n05/EiiF0hZLHYrcGpd+zoIdq4qe6ChEWiMuUp8K7HLcuVhkLf00JgnzL
OeAe36o3gQklm4yebfDeslCJNd8dSoRuTxf2iYpNJyzlMtGo2nxTWypaZjohSBuj
eQsoscYU4gAw070qjC0Clii2cPy8+FDI3VgEWdtH7ZrhbaMfdxlnpbkFM4dy4oYp
tLwieyw5WO2vkfi7YrvS8A==
`protect END_PROTECTED
