`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zCZXiKTsQnjciBEhHkxxMPyVYwtpGzXEHHepbmeuyE8WgvEzRRd+Z++fZYo/gFRl
iTDKzdHZ7urRyI1N1ooJxSv2cm/MHH2CTYNNBksNPsNIrobvk/MUU8fKx5jCh+pT
c0eFzH0VwebmHWLykAi4qVXBAclt2su3kEWArkKwqyLkXBC3sbQofjbtoqvpxUfy
Wrr9GiPfLH15FY//svYCGKSsv5zLzpBgAETDaU/i8UY+rvs1RRU61esln69Wv52V
QHEOh45vTEUAA7e+dTxdZw==
`protect END_PROTECTED
