`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lEzWO90dbs8Q2gONNculsHj5eZ1p9XqiVm8OduYClaPvz1BguvC0JxW2aKNegX0x
+IM+nM3vQ3xOVI1t+MsVOpuBGB4ldu6vnywlST6ilXnZ6+aPxiRdduzmnSkbpZcb
inSTwDho8uiolspeNuvKLgv89ogwgx4i+rVPV5mCfnsSGTnZ4EjW6LcUmahov3j0
1FyQO7+ro2SJpesO+ppYXdNC1jkIJ4x7p+wSbII3Uu5/E2yRlavcLNog8uTcxty7
GXbIFiJ1zNMknNtN/eLcgFNGWzMl7aX2NoRPD5LTxVzm357qSO/zt2rKaR1z4d4P
8EAn6rB5AnB3ydBkiyZ5tZ8Xo4Rxq/xB4d7b8t91Hlp7Q/9bvBzidyCB/Dt3T6EL
QpE9DvzINvY8x0S7rvs4SE0NdAwo5lsz0adMbDwds3X9fAfhaoS4glzWh6qwVhQZ
lSTelUBwXVzb4yMpP2l0RKl0xFHkWeM7OEdEdqBkjF2CQNcYvbqVDOqjxMaW4PVQ
8tge8kTh4rFgBBaN/1mfm8jac3ueo9vjpv0HFbhu5dw=
`protect END_PROTECTED
