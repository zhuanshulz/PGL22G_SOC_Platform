`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j2pYE8JN0mVVKcRPJZi79uIXBS6F31NzxOqWVWF2OeiPHxCEKSWbr4b/KEQ/IS7P
nJcEhNvHJd5vpT97lkqp3/U3x4ruetbMj+RMiVptfRfaalB4NbsLST9luixIUPrD
xMZEtV888CHC7WV/VOLU1xaQamNSAgQgFaZhbsLpTM8H7i06v0VhJx44wfA/dU5P
y3ftB4mU8HB7PUgvTOOZHAJNKqwp0ztg8efQA9PNvwJZELtRgC8y6SiUN6etefAC
jBCP8YVoClH+MqTItLDqExlYrmP7PDYLCUcjuCDugn/whgW4YQ9onCU6+7NRU8/l
u4KyiM/352NrmnTSwQnIME180X+DPaA+PO7CsDrbO8ngAB+A6EvLHf87UhToRqRv
eV0CnqN462hW0tL0oh31AOaY/jDFCu+kGua0tCMDJdLGMkxt3gWAFwrUMIwkZDU/
6KQD1eE5oyucRyssfbpf0om6rc4GX/W2cQu4Fj0z0kbgZ/E+TSwNIB/HAw45dFyr
gzC5aRDjUefuUb7whRQyJw==
`protect END_PROTECTED
