`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
19R1yPeStJpjr4n6PPq03t+T16ilvk7IMYsKWhwM+/NXZ36NZ3XsyjkpbShywpTk
KBuW+0llUzJ5xcvS8IteSO2vfDT/izCxtvwaxxBjsZLOzyMYGzNmEZQd38FgQHZf
GtqKsRi938Rj49BIFJimSAPBSblmYJdY1v9aK5ol6osLXtiY5fw22M74ijIfsnwd
W6kH9nvXRrl3ou+1eyOUnOItHj1WDxUFYe+CKJuPbxUZtwteHX1A8Ntk8iZblNDJ
+Vdsx18Rxafs2guKy4LB2PiQQkVAKurlpJzHKtPVsMp3iIGP+Tmd9t5xmO//527g
XPRsb8w4s/51i7/lulidzkudF76KpDKFYOZ2//aK21jliEB2XudB9xwNRDQAHqRE
HVsb3lVkjoimKBV7iZIrOorRu7/XIt8Kt3Xz3U/e5TlG/VR5VVAy0seyDRDGiL1i
Z8/Y33aMzHLBZ2+izktejAkAYjyTo+I5HRYfnofDlHQJT9urKcFt7XI1CiGOYI8B
JwJ576FWTEpN0a56s0Vy+47+xG8vyxZ14HfAgUbeJncSBEOYCA8Fn5wOfbjqhVIS
ImUa5jpMqOpvE0JiRFxkj8m6+XgCELxXT1cPq0q29kB066XF+hr7/+MgvM+ZM8hD
PPUKBKhqIpRA3l0I7Li75L3WYtFzpY8sTiXXUrwK84te2sAiHSLhnni/4+S2kT6C
daoFO6IYOAHozjo6khf/RVuDZM5H/97nNnhZVoICC8hKfK79naKHaiXy+/tCmUFS
q+I9i/uFZDTA1vE1p/7KGU03fjv/dfPsHX5n/EbpqCC2DgCkXsY89R73atNam8/n
i2nK7O6Sav974f5SiClzcyAli95Alnak3SH+6QO/eQefnT9ypErKK9s0xvH30Zro
o8JMDpCzGXpmzSYslsPeKHYTFemRn4MsXTln5L4K7JunoPv+1NIoPJv6pb36BbC9
vbrKgwzsmavzqXtZ0idZRg==
`protect END_PROTECTED
