`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RbWy3UKlalXOP4+Wi6KHljz7PyEcSMzhGd/4hNjMpiEB0jdOyI7XSYF8D331AV02
C3yL6Jm/IuhBkkluPgO8cggYYhrJBwnNHzpvJxA3Rio+9dF1hyEz5r5kEP8qRV6C
pQ9y7hg1W4tlgb/JLdtlw2ramBneiRC+9gY8NmJSMklQPbhFoJNBB8niogn6iih9
QcivmCcHlYsh04PtR3uLuktT/IRHy/LQditSXhXqDtmMIZMhpyerWWiSeitEioOM
8rEM8s90c2tebj69aJNHDquwiU7SuFgebRtpxkS+m0w+RZLehiNa2bCeh5/Jw44e
rvQmFdIpeBnuqevw6fk4isK78aZHMj6rEv+tors8nDIFDpcAxbOQTOd1cioswC6Q
Hqhl70MCCp0OSkv8dmA5YZysNW/Nxgs6fplw2rmRbbGSiJAzmnijqS0hTSaUIBsc
OiyHYk67YpO/c2zTdR+ai932KbwzF/8k6DRAH8Hbo71805dzG8MwMkAQgT9OKNNz
SLMtdxjWfjJNJUhEvYac57kcNfexY9VH90rroWOcCmMb8buatDFkaDUaZHD5EsT6
p9dtEuaJ7I5zDyelsOA7f6DGxO4jPdQxlhoU0OUunG1Snz4nKBwpVqUvo4THtPRt
KTwYP4UldOUZg1yuXXzyhEcCaWzzZXxCrEtCDim+GM3/Jm5PBT0Mno5FUdmPh93Z
MJZWi2/HwJ9PAp6W8xlvHAcUKcsYFkhYDuVYmciXCevymf4bxpR9D2CZ4rOnUJkf
9Nj/nS/d65eENrPo5tqEGjrQ95rwHx03ri6LLZajDHkfKQ5rTl4fVFImt2dsx4AE
EhO9GoVALrf7t7T/fApHDljHzKg2++8XjQxHy+t+5Rn+e/RDf7izdeLmCM8s9uO2
FW8oSMAZTRgIKs20vEQJq4pRazJh+RFiRh0Z450p6n0=
`protect END_PROTECTED
