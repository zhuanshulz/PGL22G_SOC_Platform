`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XJX95JKwdbL/GBVKOvkEK2gX8Gw1LtnDGgzWFlqVOW4spt9+iKao3qgCQCn95DXw
dl1nIYXmsI8HC4JFwvlnPk6urnb9yGzj6VEreXHeFT06WCio/RQmGE0C/YX2A3K3
0dGK5ZpyKT1BO45RAtBAttPj1L/IkS4TuQfLPKsZ5sLc0KxxDQulJ7OuA89JNkMs
7/bF8wAPQwrGs1NkXkejNRBdCAsLqaA9QpmnGjRDh7GKpAouj1tDh2/fvH2ROIEq
KPxMGjgvovZNBgdjkTLFG3MmZqVa9xxOUxEK09ba6w0oUlHFrxerKrxR08BYJLmV
DZ9IKdzCgKJV5YpfuN/RJEG0pLHywbvab1JqSWBFJX2vmYfE0NBxlxnnnsbdFXo1
a7V1dzkPw6YXH8XLKXdcFPcT/mjiajItnatg6JcPdyxeDJfbXxB8YFsFNYYWScYM
i0zDgy8QrxEluJpXGFjz+PIVmiWMeqMpA2ncKZCki+aqrzNfALHzH2ZrYjBeC10i
f45CLC7zZlP0guKuLbTb83q7m56b++rsXl/XqF+YaHkPNUEHUI7DxlRjzFYCq2JZ
ibl74XVFCV6rau10f4utvO4axVhGGDAOQpjS3WUe07EzxmHiwLH3+OtFSQ9WuIMJ
plWZe9VwUB5Bd4KfksAEPug2cgxn1eRf8II5wFZQV7Uc66y9UzoptIvJYqhp06Ee
RkI7kjVX1eKvm4Wx13hmZiyaUATdID0YeLAWH3oVY3a1pHuLt8k3PxQ6xzzgEvGe
Oe9aoIb5uq54cJJiqYGmReShvC1F59Z41egfwPAwrFJ8wzkELa7tECeb5EDkQ6c1
8tAHXn58C7RbpkV+sAt2d0ijK0GJCn1nvETpO+4FtMJaXolFKr0fkat771QAwlmZ
oi/gXt4jgWyLzJ8o5hAdl/Por2o/q5xcvBxBNZ0T5Ul7e3xVifeSSIv5mX4XsveU
Zk2ytRH/8lQ9H44ir9P3F1wCVSP6zCrwOuo7LEcXLTuFZjyhx1DqASh4UaFTKhuU
+bfxHY2d9hucsuwdyzpD9bFeZVJ1I8CE5eNd+AqhRYIHQntEgSsZEbq0MAnRGQVQ
n1ucYGw7sQ0Eb/LJ/yP4ewChKavFBMoahNBm68rEbryXB2CnT+4B4FC5pXpheGTh
Q/kdCVhyKKc7fiG+du8hyOvyEyjjpchW2A5ZmjcZ9ek4Xq8ayuF6592S1oSutEJt
duMwuiMaNKBCb7mfFRdXnmeH9753T2Xz0If7J1dSvjeF36loujH2FZ+fEoeHE7kW
MMjqnst9YH8RClcR1XIEbyIPIT/9drHVQ0iHwIOTPyW8sKy6G7BBtIw7Aux4ZTxk
gkuneEkozb8Oa2gcDMki3EefSpUfXD+d5qwJ9fS+pCZvUyyR/JMvzmYDjdx4g2I5
IX+U0MoLTj2JNxgzhqWYTnQrhAde6qvmNIldJ+iJqUNWxXhivxcnT/FaIpMFREGQ
jCTmSOLZUnccQKi+ctKt6/jhgrU/gv+g/SDJ8HNWWTULg7F8KD5KRheGmv4KXDjB
YnIB2X9mXdvDjCC8u2ytOriIZm6eWi5RDeFLjJk6mcXTZLExkLtCKNrV5z1CLcNz
T5vqcFyKF5SCvU5GbgqpUFDqIRHXzV+qcXgqzfEdoi8wArGDRAniuRKbPE+Z7SWI
+ajBvRDGmbeAd0nJPHWPZ2WF50X6IQ/5Qb81R44NKdEQqiWkEnstvC/u9l6HWWSo
OUq91AafLi5ajAsKujcXcEX3N64t4U1yFQ3DVl3aXc9sKIT+RvpQsh4lHSCyu+R7
I53f86ggcniIayPePoUkZGVD0ZOIFYfebZaC7jVkoIomF91gGRdIRgebs7ZWT/ND
b6a5F/CLyIZvNoERSkPMOWT3ts7IgNnZvNEzfY+m1+KzMM4HBnPvBItnVGsx1dmv
INQFau1H0OOmM232rGkEFwiu6tDgXy5arT1+lI7oA85mxgVX5z/L2oP9E2SvZrmW
flQfEMkj93fu38uSXYp/gb0BpMvcqU2lM+Lft30yNnOXGkJHk/H4hY5mw9se0dUZ
FBgeuN0OFg0BYiqck8+5bcpUVEi3zwPa3br7JjtO5JanktIqcIM7Qw8xFUIYKioG
HKn9L1b9tPhzfF8tF3z8Dsx0FsGHKM+mDFwFgMFo524M1mcTwSyM1SbA2bNdmTU+
`protect END_PROTECTED
