`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hfJgFAtiJpxA3604gKOB/+cXc1RtnHQrWUHHhOl0S1PR8d5Dz9nFx3SyAMNIuJPa
GqeO7b7iA3C2KAjP2Yc+FjIbSIDCEgEWdbsLktTXZcGczH16drNki3R0EUm6EO8n
nabQ6lXM3EiEbBLFCmuzT51dnjinxZyRt0ojhALW2XEItCOoHS3WZ4nWmlATIzZ8
LqtQJAlolcMwkSpxH/8VWZd6I+E6OZZkDtuNROLqSQnA5C8w3V8Pk68oZPn+bGr1
6KyB6UxynjPZkT7LQ5X263lduxDw0XkrKT0VeN2mBQZRDWrFmbpE2v/VWNiNXun/
XFr0i2PICoyYtFQfeaOUFLPqkiLIipG2pMV3Hl/o9eN1ax37k49kz58AnIexFkz+
MlRxtZ+qOKolOYuSwuQTyE4w+y4hboEVi2poHPRsNwQYSbrVrd0mBaKjbAvDitTT
tdCslUoMsdneNV0E4Elq4KzST/cg4feOWSoyWZwArG7U2Htl8MHp4QluAhSEQgCM
QcOF8lEvfIEm32YzpoLitQpNXYVDyXU45HqMkBNk1MPSKLne8bVicSGRRPgSZ3+B
eQXgqfUIbUIhby/EEi3BnBFI8RU51fLNvO+9wCm4sdEMIDMLzck9+KqWAUR2LWig
2hqgQUn+g2rnwgNWzunyDxyQa6S9RWvAGqUcJeZxrwQLml1y2e6l4+ZdEXxYn1Gi
/CJmc2m89ZbQEVhKOZXMlEVuJPlKcP2Aq9ANIuFkNiAZqTJ6c1h300XSQf73+zch
Sf4IybAreTonsT5VcWtou5dL2WSKYMzaGNlz/oCgYt5W9bU0KDOokf303KJW27L0
thYaYTNruv0aMrx8hpPz+X1ACC9DnT8MHhh/Pu1BF+zo65i7KXQNEbltcEMZCq5Y
U5gb15qRceCG8xWdVoZr19ekvxPtCvd1pbQQobqdToFnnCTkMO4TZWE8tW+PZGPv
6o4xekxya4ixTo0/kSXfm3XGWoFfBKy9lyWQthQGh+7nTfR6jccc8dPFk0FaRGGZ
hBgweXJEOJ0Y7/+JpjzksytNXl2pB/glrVB1eJVDAQfxI83SbANQWYidkF9Pf59M
hYI71EdwbLvloFp6dVI3+dLseUPht3pBcRedvXqPndxIvFpQUbYDXgLPMgL9I5Lv
gBxQCnuJGAEh520VuPc02aztopgT9FTS5JAnCJcIVs0qt0qbqVTj6ov6ciyFDuz4
MuFZVdcJmTXGURJvIO0tn1bJ6ioAhOrOi5NNInjTrAmCXO183I9zjJbimum7WgVL
zbQjV5Qt1UckgCeZxQEJoWiv4tz6O9Av9k3+uo8d7PPFM4Q5aNtCIYujlxS+mBmw
smauY7BgSLRDF+ZNTQfxjJ4W6FaW/3WurOLI9JQcWZtYgP75nBpqcYPT9ISjA8Jx
kdO22U2nBoF7aGFHrD8yr1CfbGhAV74mBeWDzChuf7jC52aZhZPJDnmTLosxY/42
spUCXDfbElnLu0uh+1dJIBhq8NeYMjPpCBinui6jekQ9+dfplePObiTySVJH+2tH
en+1GqxEp8lJx+Jpl5EFjCVcv2Dzzt/gploiy9AjMxzzzOEsTNKakjKdCK3z+psw
bc9J7Idy6uwXcadqNg6SzhP6pGMu/G5HkQBnC9WIi77JPTIRuMRwg/uWypTQv2q/
jSr3dWFoY0QmV2gOkUHeNcdrDdLWLzRXRSdKICC+DgbN9CUPYwsuemIQdcmFd3/K
gftBl2Wvi5dgqO9B6Iohx2lPsdDBBlcG45zc/hsCXtRv7S3lWhuuwVmkSKjv3kIl
z8rX2Cdi06XWZCdahqisPTjBVSd0Dvhd8XlRqANZxFtziASJrgKiUz7ilKya6qQ/
B9SH40t3OsolYMHNxKXt08peYHkyGsip3YRnaG1z2jhG/93BIR/DC4+zzRdu5qai
7l6poKWa7DEad6244G+nealGUINArhQbi8MOm5VtPyGidfaPn2LfrTR01o8bxWT8
om4mD1e99kqBNmnaQhzb+cULBtKfdfMxcXv1P5pzjzNnOMDZopyC8ugYR/hjQBSV
NmCMlQGWZngTjz+F1TWZ1dCATn10xQB1gQtZ0hVmhumMzdGvvn8NE4S5zb58EN8w
u+gPISUdQ+Y9lQP3jvG2e4iLBo8FZZeRYUMOCN5Wa+uk0lZbh6ahN/IiV/zs1tTV
lzUt3qoOGFAvZqcvVXg3MgrDrW9fNJOWbXkovih1Q/CdqxJTmCLsE57mS9RArb3I
3BdPFxDIqK1dcLHlwXBxM3KAA5dl8fwW7YFi2eQNAgFkyQaRKsW640TOKRLxgdI7
CHxMxJbckzriw6tEAR4XtQhHzWHzpzw3LTAob+Y9o0TfRsbzXttC/xefnBZB5J7v
`protect END_PROTECTED
