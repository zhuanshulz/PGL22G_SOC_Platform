`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OKQPte8zX/L2J7IJWLXwxj5VZGoDxRolrywgs8cT9W28ukiDtoXwqq7Ha6QBgqJa
YiUR6c3uQRSJ/VcmRYIk3JH+3kQc1LcyEgKlu9LKkGDrtmFvfdcd80uMkhAeRm+O
74gS7XZhm3n3nClW9DXjFcI6KERAWpbTLiWMVWmtZ8UgVKVw7esr3rfOv4PcMjDr
JPSLQIVsI+eVx11iSImWZ2wrhtBLweI25A/5z4TL6D0qnoXRk9PvGZV2seL6/xF4
IPg/a/uWIjZnn2lPwP6oiMGVu0h8zWT6QlBTSnWyewlX2oMwclHkH7m69AdNZxT9
DMJ0+CO7tj+u/gxm+l5/SPnlziMvmoOBaMVMDGnqvRU6N0KbmEzrQ9eV0iqvk6qy
+8VYhR/y7NUj1fz9dLTbc3VuWJE885t7TS0Mb6hb47PDpoiKwL/oUODyYDxM98iK
`protect END_PROTECTED
