`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0C4ME7oCk7Hl4Isl92EYUYRS5BY+SLbx9qEdEopC2Z10782ksJE18iVKULRbGuY5
ob3GavKrg83bLRu7WTLBwg7LsODSzuwWM0x5SSdIeZ7gc4rIAesE87JD7PmiZLj3
+/gW0La4bAGt5B1AoasVKSdFe5iqU8wWgVkCu3NAe5BuQK7HiDjZzsYFiFHvEvgj
BTOeVcV7limjYJZQmM+o1emwm7WwfXVZqvtqboJ7gzmhyYCqZUGkOwgpbEJ0HG4t
4wQfTd5z2ORtwrMjwdRrK5LomA1GxP4t07EE6gQiq+NjHM436svYWaJI4xwSEdA9
sygpKLq2a0gkRziDEMlqage7v2EPWxxwwRXJd9bficD7fNsMLTksGNd/sqUb+ueb
5GlsPHrzcImceNy2tkDnMtj9DdQxuPYhdHvFhZbkHA19ka59CbNBc6Xywcx7Ln3v
hOMwib4fEn9zEkEnASSkQg+1iF3u4VDeBfWlNqC2wcXRa69uVB2lB1d+odKK7KiK
hHYeKFZxYYfYC9HgnyQCQ4vRvcu6SZm/3h3E30uXYdp5Ss7XQWQwcg3GoIpqxCjt
1xjyK887bgyQwh3LJsVN93PjAWh3VPDjeIGrP3xtWF1X8mkp/Xc5mIz7yVBbhAFM
N5zAk9uBv+ZQn7Tq46sP0FI01LeQPgKx+7icMAywNIW9rHw5QrRaKA3gBbhnX0Pc
E0hfusYQUFuBLGh0DrWGk0Dlhs+mDgtFb8NXRdYP/SYqV6zv6XuShOG3JifYoTS7
1loG7rDZnJhCEGuD3FKzUryJTxRabp3Iq9/7VL2zkboOdf4XVd2UeFmCW3R539xK
9C5vjr9W4ebrSG0UsZGivJ9BHlACoZM2yRDJq0mHfvfSH61aJtO2AeisHg5tJ+MW
1zosyODkskBnK4BMJArdFjavbXJTaNNG3PG30s/MksbEzOWRh4FvjeZjIHmVPhum
k9UWyWnj3x4JAR+DTOJSIlkCNmrE+uWDhITNA/yc7/0pIy0duwan24gNfMTW6tf1
2ihB/hvwBNMIDPBfJsrKiUYA/+aWMQw814a0ECCKG1b+vQkyqw2fy9DCIZZn3hd2
I8TsujpZgl11+dm4iEGibfpY7QuSTIBhgGZ4pzg4OWpqL37QmjVYpLMuZziuq2l/
cvxQgNlbywZ0K7LpLRVHmm4Vtyfoc94EYE9QZy8hVMbLK/frgyvm/u33/FtWC0pn
6oiZzgDtxvRhxE5oREVoMbkabi9srJRXfFqASbzpOb2iyry7f61Pmri5B2/Sh6MZ
rFxRGz5vFL5nnMLVXDo0MjmxYtiGL2cPvIHz1R8RHX4=
`protect END_PROTECTED
