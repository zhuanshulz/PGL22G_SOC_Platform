`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8GufW5dhz175uNhNoQRZqeLgZi6U2F/3wxb83fCQ2TV0g55x3/7nHInblDN2ajjD
mzs5j/vhDRZlTYegi9HSSgaD4n7AbB4ZXpFB3Ye00YtmQPKR0lgiLXo2237+zEDH
02SVRRAts8TqOj9C2d3g7EfIqY+DTFp0NWo9lVgfKYJMhhMcy8D2oKEiwV7nu1t+
u6fi7lga44QC1saEWDYyVS8KAVbapFH6IuFGugJwj4z2D40t6dT2xt/U5WIJdzam
MOQwqKOygrr/gFSlVp6JVmCDmA3P3+Yq5LaMdEyKxR2bmMUa3zxCobgPe9UKKQGA
cKFu9tL/cgJe5JgwL21BowXyCJ1AmDaSXcrvR3o090ay2XtHVsAafw2ovYPtqooE
Cnlazry9wTZI+EkajCWwpGddlnuS5vnz7Jf6+lG9HJIxLzOhOzo1EgT9C5saBLqE
L6U4l0IlIzZwZpdWlmhqtcJqTM9/MFuYwHSqthzsiX+05qVzklgOVOejUXgYFc0i
x6mbJL44rijjYQx0DUhdZsGoGTvMjg1ZYtSev9YLmsMvvEJGWCsYrwadOIbOj3VY
tFeGY4UUd1x9avyh6/5msh7F+usBOckcDniL/IxY6b44NeOsGHUl2ry6ZrlWRv+i
uzjuxom9R82fR8WqlpwIOkm4M69HvNvaKwTFRM7V10SA6zEGatN9JKbMZzszaRzx
3SYkM6TjnSwv5xn1kUXQCOWNe1xbYf5hqY1IfZhk26c=
`protect END_PROTECTED
