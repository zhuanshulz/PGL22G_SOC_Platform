`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E8QmoRkYXA5hOoDd34H3J2B5NhjwtopEHr4gdl6TelZp0msUv05W3ekuqkC/qY8t
YhhlWLVvtdJmY/D87Jj2zBKvqzyj7eUCU1y85ChEHTjKbPDIN0JUp0/TO0HAc/Dj
LLVoBTZVmi6Fp0DHtmkCJG+KLE9GZPrPqWi+oXndfYUKfxgtvCVTtkBFzub8NJ6P
xPH7MUlHjyTi7WaqQt8XJ/x4o5GfCl9uKytZcUntXQ9/vR8bg1JFQn736OVukeg1
nvivAr0dl3rCCPlUzhvrqNIF/QjfzjWg7lEEZSlkV21f3VVkzN3orblXys2tM4gc
ACDxL4xaiY0jymFShF/zZU7Q9PQ+LMWEx2whIu8QmDEjOWYA9ugSJsG5b47smUPm
5EBP0z/+cjK+Z4Qe5kn/pSfUQ0N3RsLLQNpzBGz9cmttmlEFAIi863SbWkCLW1FI
wTkdYd89SAfVWLPF6s38Qg==
`protect END_PROTECTED
