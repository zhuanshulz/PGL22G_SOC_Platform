`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KV2j8U0Gvy+TsFlOJ038Qi6+pSGFyuH4lhuGvG+APW+pNUyQjDSU19xR+w/qoaHS
uubMKG0CvyQ3hf/kH1TTkWvak4F6k2ofivusEQzyUvcJPhfG/a5/MHVDlqfpxlaV
ddd53qyKbL5evazqsn/UKxaMDU9ItaId7Ys8Gb5/IHtgzf5KOZBIv1axjtk9o8Wt
znr8MkuagOtYRBJ1W2KDUD5dHFeu6OU5ZrZ4dKKksyunkJ+X8M5I1lhL7xmZWOPW
Fi6RX4+e1ho+OFq3cJGXiJCU9BudQpHSvYkNaqoDEk2j7zRMoXNPHpyL9MUFPH8f
tuh5ZHQcMEaSvshEg2KjcJYDZcgu9hIyr+JVwWcNU6ogvBwqZ6UNsfwkG4V68StM
wCmB71nlI0PLJAMdVytF6A+A6quo7dIGmGf/Sc/5un3jk2JV5mYE/WUlodahmLMr
b2s/K/GsStI6DaEIAZGKRS3WTHCl8tLvR3KLM7T13AZ5Svf5GuCDfsAWNA/92VUE
ttSKqzqXOgti2D471fXLhZymSX3k86rXV2LW/jUtVlfZJzVWpTBPnvfXNzo0Uw7M
dpSXIMJmtozj+RtCuMujWnvyaIE0Lgf+3jgKeCPPsRk6Lu3d+TCeEE2yi8b6DPAX
mA3ioR4MmK3jncDY5a+x697/gU+dgL0iTK3b6jCJu9NEQQhabXgIdhngsi1PPH+W
r/LWvLYbZ8+o39awfgdobWWAycf/KtY0mkmRv81jhOLkUnjgWcXorzpMH4k5q5HN
83ZYd6BtZKAsgW79xLExrA==
`protect END_PROTECTED
