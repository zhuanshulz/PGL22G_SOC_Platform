`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LB56K0ENi220HxHj74iicVV1r8Gs3yVVmaJzMTNl2nFizppyONWfojp9F5K5f/W9
tSSpIWNhOTTJmQkm6zLXd5LnG0xN7ObYSvnMhzxR2hXt3nbne4oyPkpPnzsXfFim
vjbxUmHzT3X2Wx9Ed/P5+dCxedowzptcgv20n+2a+rqh+1Hb2EZ3gNbmZmfNjLL8
0IQ3JBw0EtDmgyM7HalvHO9RMnpuZoOB8NFUygy0UTOnIQxbxNS3Y/bdgHfLcIM9
824dagy56qZuna+E/RDFaSE0WVeEPSNt7DktJKwvCUDXdwa8agamwfLzHgZWovUd
0nA4vyiaqjfDGrRyiW27475ZvcnFhFpOiqItmRdS1JslOj4B5K9AC/oR12CfDt2J
w/ASeFy/uE/kc29iAAQ9FHk2rSD3ObJpIbuX1hLRA9lT56LdnNXFFnJO004ORmIF
tbX5SKczm47cK9X0V8qsJOd//+WadD5jYB+bnJVHW4aNpllSu8fq5qVb+e9s4tTT
EqPWXA1uGgDGy63xJKnmc7eT0ENFHlTNOJ1sUgVaIzm5LoDtanFXg+HSb6zXqztn
Xdp2Few0JCN5G/SE9j5wIVlVoyHIrDhXnMSvCaa1GHw=
`protect END_PROTECTED
