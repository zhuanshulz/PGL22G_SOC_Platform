`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MzXRec9tCZA23crf6RrGCzYnDAO/fMNNBevrcBnCw0wH8NUOMzmRa9GS+0dfYN2x
y1KZgNQLru7u16xwdd7aVcAbOjH5KiST+JZ5fQbV7UYu1x8iZdq3IGeUDYziDIFD
4z8smHyUzIIYnlga2XgVUQ6YGYIFy6jpgQ2QO5z0pLMJjrZRAw6Jy0RtMwum4q49
J1mrz8vm8KHkTBh1WbHERzAVc5cq81dK0uuxz1qUTdqxqYkL9wCQDBwxzDRUOg89
xcHo9LAKzlf9hZm3iR2xNdI8Cyja1S2O7VCJD9Vm/9Lb4gn7SEcCvNhZvRBuzgVi
ek9xFrKUdZG83YVQpKXd0X9FtT/6JKuEBd+mKdROY+hxIR6+kH0/QvrjRaGHhneu
UExFTJupd35nvEwbeqXcAnDeX8zAdY6KTl11vlcJnyM8i0c4agL8T2PcEVJRwNOI
J/BLpGZpbbZg3ZrFmNFfSHve4fMicNKoWjK0qAQHDm/xrNXFD0nXAzrBSw4W8ul9
nW68R3sv9P41uLDD6Zxx6AtIDDlM+FXiwIjYvdSQ/aTQJmRCINrf6qfpTRzPDg4s
LTQ0/B4jvS9JdtPITTcEZtEVdbnuUZrgkBt7nnmQkixjmF5rOYAiZvoCjerCxMZi
4QbqnPva5ocJMP7LkzDA5r1L5c/rYeK4+2kQHccHWPKP4QmbCxy14zMSrfiqs80S
pjt3/SNU4Fz6vWwOPcs9Z7FrSAjc0gr9m8k/K9qyld6rJ7BexActfPO9L50uYg5L
TAlJTAktJwhlXNzpPETyLGz4kL62V3e804Gp9Wqf7q71oG/9dVGJYzrdtT30jhtJ
FNRkhUNfhyAQ+QgmXlKKK4H8N7FGq5QmDXXJfoQxdNTEA0S/uIoZo0whTG3rZNL4
CxTJ8VDMTrZirH/5zJcc5coZBDUCStH/9mNiHMwXgFKb0203Zcew+pscCFkqB/8Y
eqtVn9/QBseTXTvQoMsI0WL5WOnTm8/Pt+qrPFsKlZa+trEZgFWHVMHlcX2wQh0w
3xY1kbUYCGCKguSMTBYQNpPnE+tK3uNfw4pU/7Rj5mmstpKl9sB9ESfzHuwKEz2j
z7kgGM4kQNn4gCQ0xHRo1ojQn+h6PPdq5EKHp/3y4GX7xHi2dygUuOHOBXsISkU6
Lx5NRyiCrtVGHw16zsTYf/6wW6QfbCG0GVIxKownTCf2WZ37xckfSKaY6QD1ix1O
K/HjTYu3imMflzVCfQ2jTSy+Die/DesYCqeG+r8QT7xXiPB5j0RLSIqmaxfuHG3k
uczDRb+Q+O2pxqXAONyUA+bZvW5irzP0vnS3PD1B6nUEBOBKei4ZZhRmlQ+k0F1Z
iZzriwAQVPzAnYqUiwrdd92ff2LT29awjKGYbsZGYVMsU3B0C2V8NcyrF2O17Sh2
xdEqrkvVUjqmbVQJPxHZaSlD56enGJ3GDXUfneb0gKCaUyvI1gyAg+rbu5GFZ7jo
jx3NMsykxga2IkM4a5Ipe16QEN884BHiK1/4PpZ2Adh3R+qEItO8S42LSjSCF96N
n0Lffs0h2FpGqetDOq1KOqSCLgfvYCsm6iMA8zAlOzy1IkiCbF8l3V+WrH4J0bAf
tvIMNc0alvoq6xhEi6dKT79jx5hn0LI4Entw1yZxFUGryDKpiqgGyaBVbjGXOx7s
XSD/3EPo/fQcqxT2R1PYrGX9GRmla9UcFgjX5iDgwuE/0pJxYBiEU9Sd4AlU+Wgo
vhAOvzCcOb3LQyYHSulrDPDyRauT0c7YoaNcZAlGFBMqpdM+eVxnNKPrOjZSB8rf
tZCkFXM7e/Ds4jpPNoWF46Qq8SjPVnRsbHcZcX6ltmle3tQuVugPLhiQZYlZurk8
WnSdQ0EAydchYYbmM4InMdB+0XN2ltCJUU+mlG1YakxmFr0Fz+df7XxO3CltyGdQ
IJbgPypZlOEBrCCdp83/zZXQk94b9WLE452sWt/xw8ygV2YfIsW9h7Jh5/LBHfmP
x1pULz3rgZPZ5+YxQHpAMcnGZcFEo4gSfe7/3Z4HGrGCbHnKfgJtaO7mbHoYjGWx
wEwK87FceEcn+F7RVdunAK2yn9msa5ZyGPwcqmFX9Cb77wt+9P2adB6ueuZswBtF
K9BFFdz9umiBk0CZPPxePlQaMC24P9X3unLxSF0Vw67LCVSQKZK9gXtSB6c6UOZG
hl93s8YfW1H0ZxcUQ5QumQC9+imSwdaLRsvNn8RmPU04eQDXBBLbPGf5FjfCWNzV
H97ioTH07SBmq4yIWVu+Rx9wUm0mjCrHeFFTDR/lqmZvfxFVTcawfYWMzxwfgmOs
BdP7WyfTNwphDtmnwxrPSuL59wVPhJpKhVnEXntsQUKnbOfbmtBxEcjNfzG6/+q1
qmYjfazyiK3Vzk9Pf/8P8sidJdrEnXqYtfLzmmPnMJUEW9Lo7TdUAUREijDJDOpG
1ASmfpWASzU9ib093JHeH+8qcZTHlBsCFn/8TZazfuxgKM9Uh+Qwy9sVPxcmQIuT
fkYBVZJlbYT96ISzwWed8r/CidAvuyUvVqv/QYVuWXeUfvAA+DAQv78DG+dU+zdr
X0jDeMLDEoA5pVX1PDYwntaHv9xJMMoD8tnzDnYPTZBRpZALLa5wxrXIiNehVAYH
aE/vh/KbsHmRyyksUOXdNUB3j4iZ57IkWl9hFTTGqXWPHgu1DBWfP9C+qaX1wb3a
R0dj9wWgWh8rI24bUbGprGyGoj1l7lBmDp4nWaQFeMSl72J9dEGex2dz89I8TkKB
XgHhqYdoWmf93bz0sjf27fsNR3pEWNBdtwmL9RQLNw4v87rfem2ErAAxL46C4SQP
SIrLMslSrFDYz4TBwL7CxRmqKQLWbYdjaV7AHSW3fjQ9yTW2MRHNF7bBuFCgJygl
PAjeECAtOor/yAPdBWicTODdLe7Lsx0hh6P4o1K6vE+NPn1Ya6+IQuSc/VzBYqwm
Tom1AEeDhORsZw36Vi99y5dyYrcmuwJhMn9BQc3XRnIFUymoZp6RT/+VK3k1vRzU
KvKBoypa7qxkKZFR1OYE4ZgDrPJqBi1IS88m7pxCn9Pt3/RslWjFLeqe9drjUuot
IMm835hAfonPYrYBYTOkexpbqwQrTm8OgEw3Y8MD4G/RJ1C1VzOkj5sDJ3Fn5dhG
kyx8tsJFeAgoZqoI3xUNhljORnEJ6CAA6llRmWwd2tofk+kxDWB4zQpM9t4rIWLp
dvesJiHf2fOHqFRxTGnt8uRiqLDuUFr0hfU6Y6HStpAOyPoo4lCwE4yZYjcRpTXB
A6XGL1TeL9N56Hle+E/fvbaA/0zfMKDlgAJ2C2/MyUxtQuSffkqRbvHK2EexgxJ+
Ku1j7dIrbhTme5+EK+74j4RccodFu8XS5LkXqwx58wSFCdrsO3d5FwnYRemgP/A7
tkfs3/wLY2lmOg5X1NxbJkn+wteWSb08YsUzwrOIMCAvl9xdEyvsVSFYYvmbt1Jh
yMKNJZ/EsCeEBoQGgllOBBgajws+P+ZZiJUhfW6AThU=
`protect END_PROTECTED
