`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pxUhhA9jIrR7oEaIORgACJRLSUs+HvPXMKKB1KLaFECFmx1/PtA+VfwB34JBZ0un
L1oxty+KkYFuzQy2jPZJJN35fBEioLEEJdXuzxGQUVfHdV/3T4KFnM0W8jPB01Pw
7Mbxhn5Fs0lzr7jGR36ED2aqmh5FE0uTl5PBINwN1sAOA4WyF/nyV29C4ce9SJ2k
k508T5C3RZ7aBqDBUOkvHpgSYRjf0ONXTMrvqMlUyrRdqLph6/GURih6oeZkIQSf
NcvSAhU36QrpzQvSIFgqWOrnIeYPGTfTGHI/tNnGxG8NLqQisr/BiFvFiOuj9S30
AriQ54I2qVnt6nzZGelUow==
`protect END_PROTECTED
