`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
68aDIE/35/pC/aJBnNF3aOKHM/izKqgCxi94u2VEWzH+qdYA6tYv4nubvEBNehil
qxZDZexl889rfdQ6XsrduzWnd037TWVe9mEWJCEgyFj6qOaXGKupbRsYc00XwZ7z
Xj+LnvDOPvJGeKzcgMB7WIslReGA+n08+OVt3Ikh2HyZ6OxtCs48xZD4HaSSyRit
v/r5uC5E9zYXBiFCzOs1ptnMaOsqlbPRacBP1qVxJvc0ssz9t5WyVg2FvfU7mZl7
zYQS6j2/RpqiiPi7jNGaWfMIw7mqCcOg8tOdZjgw88gDNvntDl5ZZPBGvGsn5ELF
yakBmWZbVNjQW2m4N67B95eiGA3ItQZiS+4uUfNC0n3SECeYbwwEIFAL0vU5b6PI
y5odIXtnRVNcbIWm10m4CxKfwDVRzcGB0bbQodddQgga29rFPdiq2YfAKXJNohoJ
mZZOD0eqhqO00KsOnLfa++b2vKbGFTfU1LATiLnbvMjIMmLr6FkVSwR306XjaDMH
VVN1WopZw8NM+VQF95YjRQ==
`protect END_PROTECTED
