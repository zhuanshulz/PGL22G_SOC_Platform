`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t/t/1o3Lnjpc5E6lpWCicSzehHBRQJSjcGtMwl5Lwl1NEppe4BEcDRYp93W2tRwW
mZs2EgVXE98aHv5Mz+dmI+7xdwTbhOuc44ycc0CUzk1/9ryt0ncEZppDD9nWGMJf
4/f08CoC0FfAb25WPbdUyfO95SyBMcLxq0zhl0u1wdSSuHJ4wZl2tsTfJEwDgV4v
UHCNCqNAN8I88XrTM4POWHCKaZr/+6uzDe2Jb7mHk5m//kRf1+MTa1aY4fpIl2cO
nziP05uI/QRInaUgHjq0PWv9PBri2XtexNKu5YYV9IKY1ZJFjdr1RhnjqE9Q1DDU
2PDv1Ev4IY9wSFuVaKWPo6BxA2ugNrJRcS15nI2Gc/RpG20BXOk4JMwUwbYd8hzx
lFd4gQg8yZO+dilRSHAmFLjoisdqcS0Xu12cVNWnhndV8hE/knxQPAz3P2DGkKlO
82aYzlfKlFHJiNC204e1HW3vG+VRCcAq2biEDtXjPRmFqGDFW4W+6/a4W+k7BAzf
1rNgSiQcLi8hzDlztHgCjWwJFABiNA3IQMCT1PEvVe1RM50w2rf55xz2zRKhHrx4
HKX5OXfSDps8pyjnRZI7hv7HordDUkYK85p4Y/a+f2Z0GPvdBKza1dWjogy+vLlL
U51rqEsvZJiKw13wOtLkzZP9AY73v8TLuTWqXzqqdGfofYH1rjcjhL483MMsET4Z
jHCecVqhvaSgSt+0mj/K2yf8ltNXvcHmcTdPZbpfLILPKS2DWG4jA44xdbqx7O84
fsL3MnfvF5SvAtrIcEEoUiD0Q6hrY1ABDWFkbLcJl0dgFvWTrFHsC73P+OCGVBGW
PAUGSHjBrCi9bOgUciPYIHZx8niK4Bs2T+dn9CNL2+gK61GrepmxndyOJCPj916L
+tZQLEjKZo6Rw9Lghv1CXsDAgxsTfh0cV9WF/BHfsVKTIFsO54vP6GVVqDpEz7cg
DM39fyW4dyoFmvSkbvmhQ90Wc/66UkmbkXnq9x2JkX8nri3hh0qo1a6F/D+IsSKC
Iyf+QvRnaya3hW3vJ6zFcGi7Q4itWYa9mhnZxt3Zr1KUosOzQ9XyyvGpUyo1bZ11
88k2Xc5S+VUVn5R5fQSXNjohvqcJE7sYfWgQ2PCM+BkQvx2wfqQZQnUTvbnpzRef
iqJoZ8fdbip9zSbA/uTySnpH0S3oE8lCv1zM0J6mku9KV3xtVXpApWAcgl58wWPD
oaGSFrPHu93EbjecP8IY4WirwVhYAyhRgnIPYEEgVZA1ptsRfeFDMcUJtRMPIOUV
TsJsrJEMpyDzPBt6QZp1GALMZk5wh4FHNprRXwi4QJPJnoDjjPLC+zkFZyyuwvvV
pxQ5GIlyux/UT/+nzVBOCTgCZ0CsbBsTgDO60cQaLRxUZ5p095pm5gUXPOVnm8zW
MHHUp/FUaKf7XDhw2qE2lzn4S2XWzHmYtDDDOM/yqC/slOgwb6ZfMh89QgtJ+J1H
6aCHlRoGvJ44RVPSbZdkaKRaaL0A8rnCEsslXLksveGOajABphuHATbAY5Baiiug
lyH8uIAz+VnQX9EfnViLm8ZyAMvvzxOZ+d8zNR4I8gj85r0DeZ+3RpGAUHnO91ym
OsprjYeoGGAiwiM8o2rYjHXacCBkX9ghVls+uavLkvCikjvN/9KRksb2IpZVXNYZ
tKGembeTs59TPOZ//QOOnm7OHivCDh0Ea/dDZjmQB24WMTC1zY1zjNsMz8ipuaqy
7uun9/OxYkuBcQqyQFcOb3Uhy3NF4ahW1uKonrcksBKMrmhZW5hl7Nm077Bmriuv
0y1dt05aglxDqZNYS+ytrdfv1z2DQ4oCS4dGn485/whEtA+8poK+1wb6lalq9Tq2
G6QUKKgz0AH9qZ6TArFwoWEs1FrDWyOP+JyAtAiwrobAfvsQqZgIerFNQ8ujoiL0
zc2JF8Q+32A8ls2OcecmWGYtiPHDEWH/bsB5NghN+ZC63MYNJRyJob+qhRmnoMCk
PoenBA+smC3vOmESFES3Ccc7sXSH4393AtBBJjZ9+VqNh6CuSFYk+pVeljdTko1s
NrkJkzLU1LPXtV8WuJTBXaXNdUun/wy7wH5YXeeoTuSXSlwMPPy1SbsW22s99Z8c
mB5PEctvkRrt53DvKebICYaVB1hM5396v4LLASdOIlRd5fYA6Hsqv9zRp/bj5o7s
hJoRZ9wjXfZ4qYosspRAmdEiPNgmnidixeoJj7iZU9RGNbMRIWHlArgRACD2WFkr
cWBPbvSYrrS+/CxtgFojUzc89rFi+Bllm97K9PnZAnzjCOyxwFqiUJx5uwe8RjsG
ZeXWvw8U+5lXFApLHf/vP5u2M7d1cFQUt6Bq6Gr3D8OBGlqxRZY0dXsYi0dw6vPX
QkadbbX7upuSZ/uPwmD1LhCcFl4bft52aP2uc80UbXJf7bJIKi1UrH/IMBhG1lwO
RhbCzX+mWp8OmlTt02QvkQUjC4wk6TbUR08Unep1o6ftPojriLZrgW2s/N4P6Stn
ldFF1oXrVFokYUMEz2BAWJoQX32mLwVmK7HuElrfnghcGh5RA+P/gc8QyTUt8Ep9
SZsISgs90Nq2uHcxIa5mQmOdNfSfMFpEEyVkzE41cjIenmnfNdtiubpZwcvEGaw8
D5hd4dLPABvYRjmaZAX05A4KA+yx3zOIhXbvfg/0MoErphCpgkrcMK8yv1RCA7ES
fzAEdA2mwhlFhY4ZTbDRCX0UkWD50Wk3iZ31TMYh2r7AK4uF1tvgStPlkZRaWmZE
uVSxwZwvGqW4Nq0Uw0fr+UXmbBgwFUSysc9S7dhP/snOdd2jdgpbHQxPzEhKn280
ebi6i01CmeXxVW/W51TlF+x5NK4M2ZlZ4FldPVXFtKIVuwrVeR1kXugmTXioBtgw
yjcKtUc6aM7m4gEubD+qdyMKKaWgo/FU7rluVfAAg4NYOuvHB63NVKezN/MZrnsx
t3R87dSwQD+YxjvdNwOua4SLqrraQeZchaqqd04oqTtYw8am+UcDk8M3t6BgdZx7
dj3kYOSBEimJBiaujbuc3RpFpn1+KvaXjpYJZhFdIWTnwZkYQawXCd+8lipgkSh8
RqWMk5yb3e5m/I61MQg3NeNZw93rrhICFkk+tVbVV12Xp5fWEtKsL1Tcx0wMGTTu
UKyj/jLU1DfSISQ4bRewGYDVHzlyuVgInaN8HrrptJ5iOT9/P5DF9XlJyrrxoP6j
4Y60RCW3jjA3hDMbc1jhEwQtQhBnjqBaLxn6/9EwdlrDadYjcVmZcLWCwqT6vH4k
/l1MENfDFvDbJeTe49kFCPLJZQKgbIUh2n2eZ9UTE2/Bna6T+OM+HyMN5jWv1u/W
L8aq8JjrzUo2x1zLEooTN20X0NBFBKvMth1nbvyjXPWng8x8X/YsLo4qPnWibqxN
9s5nlomNi0fmkWi4JrdvJJjUBWZngOTUlJfnyHdImuIPdEmuiE0nxbLMrxOsEmfS
aESfqvDSqYYFE+pPLKu7ZP1yEPIRCGw0YoHrbdJsHlRJqrafa0ioO+XoGfxc80kx
XNizFOLPhDn4KmELx6Qoc9WhVe6DUKeq4YyxOkc1OSDbpf95Dg0CNdPXQCqC+oN/
0W0AEyUuPCXBGaz1QcKSq+nhJ6hZbntuZDClrkCf9ZFQZP4xc54LeNiXFtWTGbpt
dFj1zI3ZE5Z+RHuUNh/GJZ1EnOP8ER2pYWBnJlrYe11NAxuNZSXk9TX7q8cB/9zn
pvH7mgUQ5ZovVJ6thm+WCmn1zuI8X4WDLs8m1JQ5aoaX6QCfRgxQP7OMxUz7KejD
TClYQc9nu7vhanA4nTK+jlWxfwSUMvyzPSvoAInoXdNk/jR7dbIYC0gSOrePrgz2
o/k0qEhweOPCQOsRO9vPXZ+8SdtN1KgKFp+MTGdy2JspQLH1ccEseybZAeKKG4eT
oPhIX7OcF28QyaVItYjKhm1YPsA0+EANI3QrtU4SfOPUkA0UaGj4i2tAV3WTuTda
sImTOQgkk9zFVrrUzw6kabP0zMLK8T5xVaTLCHmVCHtwg3aBQ7Hm42RFLRCtq0MW
toJSUwoFpmihWGuCnxxd8Xguq52kxC2INX6WydDex5EMVoczoHKVMesHjA11OGO6
KLTV/Dc7zylUwiPbZUnDKEqm4ZyP7VBWgStbdE3YgD4MaG5jADqqc+7CdQVREM/w
UTLzAUSNmdbOn2UTxG2AT5PuOeX5/OfIm3yK3NptasuQjJoyPwt5qntsO9WAuQCG
Ml+QacEVEoyYe1sOn2tQHrGqJ/KX9nXzUREjmDA7hgMjtNfDB7F9WHixtPhZP77I
fbSc31IiM92vmvOykqrcQRJFCHdYzPVYO2MFvFWDjU4IvBLI/btaE/+DEg7PkQbJ
+j6KnZFJXH9gLq9pJo0m5wirkPKxHxVOVhsyjwe9oUnZwhiZtU6IMLVUbocTPRmJ
s6zBM9m2mScQ+hgH1OyU+cYBLtNUio+sTcEisczjoLsnq717ZwyzNnS13zRyFs3N
7aF4YY6vcEl1k9LVKdU5HouowyHL3tT3aNdi1fXaWOiPPkJPU3WvnVy3LkHZXmJO
gbLstbFlJJukqDT40F2pyUTghZz8R5ypFeHLHK1sJJhmzfM0LRmz5H0HD2/1blwo
t4FiDMTXvMrmdQhIDeA4Cj42VKeJ7D5rID5I9C+15PcmhtFKkmgR/dwdaV/xQlEh
jmnxfB4H4mEFAEopGJ61Z/3F4bYOpd6NSxyoT9SAiMkxrV7i+dPWS+GW7TcpOPK1
bTpRK2QLpFkryBnL1scnZjAC7ui7yK6EALbbuPpS/kao9uoEHkGBZk0TCBjuIFeq
z3wmUKEI76hnwgA6512U8LtGEwOdihKf3O7KEKwM/PKJY9x8DtR3CFDs5i7OMf+S
2jawZJyOncQmO3ekKLuDixFkOpnMb5JI1TOKnParXKgWoOuRwLRCnMXiqE5OWhLh
FGbanaR+2EO2MS/vZbMMeZAwnF1gt92swmg37F3HZM2kXFs5F6hPHhNrMQWOzawz
Cupu7tnn8+gjgPgT7sUHF7f06gepTQ5RNbh3WSjDAWXlrTMiq3Wf3znr0BqBRZ6c
e5UrM5uIJnZhPHL6oQ6QmI2KA/e965wQxfGTYzD0srT2LVaJTCT9ntmup7X++YS/
+LxbJjyaHoi9heLLIN8C9EWaQstUlABpJtdf4a1g9rjlNpWZdZGJ88WIlklkhIgT
1RmE79JV1h6tdo+WAlbBO2VaB7H368Woa0MtC+TR7Dg33mQzFF7+D32GHsjb/5hs
vgvEtZ4v8Lf6bsyRq/RuNaPdPBJLLr9dQ6PHw6i8J18Z9ED5ADfbKZ+7s5dF1c+y
T5SQg77Pm6rJyfG4+92FDIA+VTUDfskWEvTC8IpC9YbT66V0O8VANcwKtqNTmtFt
uahRxtYr3amJn0qqPuaWQaab+M4oEE2t7SI7uO6ItIgIqyZ3x+I3cleuRPMd4Dum
kPwly9JJnvJBUpUipHk0mOYi6tZQVIuhvnoLwNIU50Ff54N9IriPmIoe3ZVPS8Kc
k6v3zMdgg3g92/EG4wJHO7vAqfFnAMe195pPRGXJ7QGN7MEUCYyylrmjO3rUuuhf
KFkXS0fmwuYEUWsYnoGDnhvRbPpIZ0/+bxx0+aAlu0KRq2wwyO7BemR/9tcKQDKc
vEoF88bpPf3DW5pFaUvtkmOAdhO+ckW24ToV9Xu9LcwbcqM4HprC4CKnIXj1vbha
RnNztGajkMsI1C6JYz5HXbSrrJy8HpO+YT6brKlTbcVTpPu+jM2WiGRa4oJ7LbFd
zVrxvFa+ttJehlU6/oDW55Jzozd+JZNGCrX4KDwGrLUjWl23Du1t+6CynSaOJVEq
1ZMXjUAMkYJBy/5+PHuYlWLSM+O94aMnCpjGuzCRKtoGrlEdz7xSVI1GMPtT/YPb
`protect END_PROTECTED
