`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1mv8ZZ3aGazwzi0iAte8uy+R1h/cDZZd+oln1F4y6fQDCsSCENam4TtAv94h/64k
jObSV4o4YA+qYCdl+7BABJpvmZ6x11DdSRerSJiB01eGktqhcbjfYaR712CliIJs
ixQ631IDYKPDY/sQosq0wvsGG5FqsWD7gsDrgrJCaOEqim2bZRhs7sWVHoRHrNNv
sgpLP28zY5aG8tEHqC91Hw0b07ob7J8ep3q1hAR6Wpc1lKYGQmHHyeITOkNjInR+
QmYuS0jrF0ZJ2st9zzzc48fsZce/SAdyaGH9e6JToEJsQ8TyMNknbZJIjRVdROcu
D/s4e556fb0c1gLXBL526Gg8ijTYioC9yqAQIAMkWs/G8a49Z85u+/+B/xjF7Y3i
xwAUeLZXrZ6+91Y0nymdjKM0zoS60UbaShKfh7C9mk3QKat+UN8cyKEmPZvZJpO/
GrXq43DJnOYBGn7ALpq16IRysUg58n/5/pUR+bBYtMHwLvnW3dH8783LiyET0tH2
v3iuvBOtBW6Ez/XRf0yZw4KX27skLrbi5V46v+Pn2XtVm6plUPnnqwY/RGx0Log0
`protect END_PROTECTED
