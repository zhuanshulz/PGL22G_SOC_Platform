`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zitvZ0D2YSj35Vb5SVPdbCm03sGFHuTyVb5iNRVpEM6DOHKMrgQiqEtCjOpTADCh
3MricGzCyu8ajCUyEyB6wIRckuWHXMaYmx+j4yrFxu8EaEUZ0T2bdlfDRRlxS8YO
4ZpXV5yZP1u/eK5C6B+t9dTqHBh/1x58hAcTOLQFOmNfOM0LNkQp+a798FClI6MH
CJh9PYn2cT3SM87eTQPBKLvjnGn5flPfvVUDqeYfQGLK19CUmsBvsfq8G2hWEEjm
6XAAQHmedeI8c80ESamZ7Gcy45OV5D3ijxwe7CnqLjlVxFWlRttwdBnidmH/77i1
lHgF2iW44i+umBtcSpqjBPDN+LljidOTIJ4KbNnwbXpgMiwcCfhlzpVlhLJ47XO6
QoLosagQrr8SZtoOzQdFmXFMF1TTxSYpKK578HCztvjCBdvpgj11sku59+RMejkM
HgctT/98FRrV2ssZgZIm0/jxnfHQFVTNjuRGKYUKoBurmmwDuCjmR8vpT6Ewe3+h
4viLDXrwc97E5qb4ZiDOaULtDBjU+JPDX4HV990c/6dneci4rJxdRsyMj1L0Ur3r
EcGbx2KVW0EkWRI2Q1zqpGos1j7zw2R2aUv6tNeh3y4A6eXO/oCWQ53pF7oNwvD0
yNvTZ0fQwyQ0V/b+W3WHNuWLKuoazyqJdy6igwCAA1BQ1GH3J6EPsLmBVRSETeBJ
f1PlGXdulK36aA4ir6uGOhmYO3I5Ze1pXs9IUtq/L1x8wqOss5CCGbxYHrRNrzNJ
ctpxm0elNXjDXe19ATIPuRyPowias49VZvci6qN0+kYDI/hAtDu64LUiHdnBU5vg
T8eJm1DBfgVhlqSGs7OIvN6EBtpVyx6M+iNqEav1agHl3EkwIZUlbOND8cw2AgWu
W04AXIy6d/1PHt2Up2j0wEIsokHUlaCydTRTlpjvlY++uJxkdOGUmaQ4qh3qCT14
3RooOsPr6Jw3Ob6j43p7+c17Cut5QqIxSpZeBW+dbvOh5lMKl/mn7XhQLmLQe8sM
tiFniaOR+NGivV+aL73tnMd9X9uxm271nXNfdB/EPW5TWGXNvU1A+rG8grzqXl7W
xssUgNDmt+rzLkKV923vl2R+OzaPmB8z2ggosIQpuU2jPeiPwX7LoLeGogEcBsIc
SObdzTGyLz+ULCFDud6zZTFpCg6lUBMZvMAyOfx8JjA3LA2L7JSWALAOlK06TAjO
l5Tz177XdNYx7jVYO4yidDRuBKsPdwt7Jumh58Qa/dBCdZVDa6aLz9BTyds7Iu3r
00ICZiaZDt4x77g0SqazAP894jdEUoCaxuDkaSzDK+HLh4SoHnJp8SQgTDT6LLFW
E7M4bMInuTXUDtAQuX9GJffWhZkAGM7Oyq2WLFoR0VWoDt/t6veSEbS15oyQrLNy
hVYl9asVvuGmDLA27BMyL5qf0fvfrDZldsGFTToSHiYgK5POMHbqh4S2iNG0h0MC
Ca3JKJf9LrAPB2R3qAdbuFAVTUKDz/WrjKDyym+VeL/BKVsNQxPnuyKG3Om9Sa6K
EwgiKKtJedA+Oaqw0xCa2Zcg7qW00OH3vbSwShpgcLhRayKOYehuXbaD2ms4AgGS
ovMxsHfXWmsJH/0qM4Tsuing23g26j4B+I+16/k/jUeetNXKYs2ZKwM06c3QlEib
FSZ5iagy4bU2uCFWMwsT3DXV9xNRk+e+IscGdIRI1I58lJYM+RA0yLrRvtMRNJy+
JhXwYTvFXOzhtbF3YUO5LU911G2uKtbPXyeKsc8gmsExzELdi+Kdwv2dvoSBF7QK
qUzBd57NcRKXGtkuS+xZQXlJVPx+mID4VB855GAAKNVAPmMd2pTyuHJhuiD3cDrw
q5c7u60fg7PCkdr9NmQnCWFBeVyAo/W5Tt/2Vx+mJZe6q12eGlX7YHLWbQRVarzU
7VHzd8AkZh5dWCPD21p2I/MYTxr/Y3QnADJd4VfErO7Q6ZmCKHzalV5ACUX3ZUpf
DLC9Gnfgzb2jzq4gbf1jBwpNt/QU0sZi1gOISR9oH5IJp/6HukFCb/XCi6fZ0jiI
MtZCRhhGWQyK5o73vXUdLEDOTJwS587h90aVJtpvcWyKofugPyjigRO4YvivFzuj
xlg8mEOxJD3n4XuT6cI87NTxMj0giUHsYlt5hQuRGPv4EnZZCntYkCbO742eNPnA
aLxTskP6hMl/MZ5v6rZH0XkLDm7qIKVt9R8C9yURc8YhCHz8hrlh7TvzHn5o29Ic
+qMmu1ieT90e7WN8tUl+QEV1I7oVA/fvlOGxp9uvieI6+1Nv81BLGX5LddgR4MME
N9QZk396oJXuyZRKyNqNr6AiCsecQgOOWSNX8sZwLv1HnrIw1nHIOZzBbOW+UwVx
X64FRJDw/SEWKr9/tH2FeTeuby6rcIqIOi3MJScGD15VVWVNLQ0/xvhw2WJehhJ/
FgEgMNRcsD0OS1f9Oq8kXPRW775PFGsRqYjfjuOTsrCgPEEu8M5ziJ3tB8jgLJAO
MTwILpVB1eTwbpaY16fyqg/YVe2dI9IAw2wsKkNRguqd099myIGdcdTArY6Qz0LI
iPG1AdPmIEAY6E4Kuo7TkfaGxQPzG3kF7PWFCVqAXsQZJ/5LXlnkKC1tO33ps3zU
S2Jhb5p5d8zxyfHEUvQxIwnOkngiZMpUvYvaDyCywS/X0pUWUD9DpFxe2OlfFYM5
Dk3vRbjyI/JMRApPHLEigd0hLYgAf+SkXw3X5Uhg8e8xcsgYFLX9cAGrKjwKUSXv
Xs1LtuCXn+7bRfLz1qJO5AHqSBQ2oZJSPmo17BcVrHyQXg/4S2U8EJd+kt0jMsIM
8wK54Gh3IEXwfkwSTwhTIpW9XvMDQSn6Qz6AbVoMl5RODkshwKlUWQKRC++0kL1v
wSaXpHlVeWK0htD14+1Ou5vtOrD45B6nofdzLFU/G906NJB8zJ7jaY5PVuzeksZX
bxZjqTWnwrTuYKqJChvP0XW3kRNXb7pgNH3x2mr8D3PbF1ZVpDB9z1CwXTtUjBE3
oGwT9Z+3pbOJpfYtMJI181q8u2nfBzRV+bwRK+OTFxsL+ewqI5P5Rjkkvo2q475o
SvLRb4YobGVD4PgkJvLsnp5WdQ8plgH1d77czXMRd/nbDlW6hAOEuTpUoDQBhcAF
PS//h9/hRXht8Jv8wFO2N76tXbS8V5dax290M+jdgq8b+LpbNLqbgmnA6hwmQ2VB
OSUCsBz9+8YPdrVRsp1juzVd7lYxnHkFqWCQK7oQnfEge5m+cIAv2DjlpV/rMDV5
coc3xtkTGmF6z63hdCHrQ5Inhuc8U1knA5WrtP/IRSR6BLrNebe8ZH+n6ghf8Eh1
1mAZYoMJ5OT4J1YdhpYDdw==
`protect END_PROTECTED
