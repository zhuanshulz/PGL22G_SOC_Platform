`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lURZaD0yfXLjx5rJLYcAe5H23IwnV4EFVd1DZfKTCCEmytnD5YUMe5dyKpBRA3A9
f53ZtZSoiXmVa+70c8T/Bb18F4ay+pqxhKHOg6u50AK53X9+x570BZIrkIK/8XEx
b18pL4CB+KEX2dUzjJUmaFISywZozkXHc47Gxj25VK1kodqkY3qT/N96HswoP7/m
0jzrqJlB5xmvcpYNI5LGOOu/StdYu5SC/Q9ZizTboNCDeaSko0mpxkJAw2W1ddnO
1Ci0BiHhEJILv8tZ4nR5Xn0Ff8DfaX5ID/wp1d7FFLTA9dY3r/bulaxdRC0EsnTw
NFs4ZgkawN5YXWD6ktzECuddi4K7g8paa58XG9nvmSF4vvlJcDW+S2E6EdsK0rfB
abQpO6rPVbxouYbY1nP2kfKzhrQK72YpNeu2jQZTueNIhbgejVI86S0+mmZlo6Dg
N29BTPjsudPxO+sOjzNrGPo0iylwuL8bfLrf2ddP8lE3HctsUzhi5KI3+W0uEiRr
0eT7mx/l8zMYrlWkiTBwgegLvL2lVnIEh50JvyyWkgo4kaQwbVcQcJOd7E0EgQiq
raYSAsWypcqUuBY62+eWdIECpNRRr00JP8nEF95n7zs6O/rmDZEZ7eJ6EwkVNTAJ
38B15p2BM8neXkm/xZN/OOuYNSQBwjCT+V47VFJkYt7x7s07G9+wt8EXDe6dkQDT
nVORR/+Uv08zZ3dKx9u5UerenlA1ktLIOd+uF6EuwkvcuB6djc0fvR2g8j2v8PkK
3wPsTTKZezo7RdSh718sTpNY6Fcj8iMrhbhOPk1yNeEpe8yYnAY7uEEMUWUfJkaU
VL/0zbrGMU6ldeSEUiJ/aE9brf0CyHaGUnqIFMIJIZQDVrLQFBhTYM5Bh/Mdv0tR
BHLwHadwRB4fPpQP/oqNHnjJsODFJoZ9a3iNjwRHPyOR5DaGNPcHb1rMxFhgUF76
JN8HSGJsgDK7bGbv5Taht17q9fD6ambi7jVjafMzmpu70oZkz9uqg7pGyyCiGDTX
G1ZeztoCHJSkmAW+3othRDZPzTU3HfhR5fH+ESqDLiWwTzgwL2hIwK1ln7KzSA66
7nGmVMoJPUXDomk8gb/zjY2AVOEHnzCAJ98d8lz6SGF4d/Af9BgBnnRMEUQfsFcx
rZMyURVunSrS1YK7lJAb14m8UsD6QsNQ6M24JytjDWQHpOFmHfm8+iyI+FfqxiqG
sKfDcxNlDNRETIics5MnKkwkEkdUMSYfLB2zeS8fV+LmQSQy/3EivDBZYv5CT7OX
TJalTu4DihDAM7StSC5JD3q1I9ZHAVPHzMMfJrS39kiAwDXsK1qAgQcGyDYv0aMe
7DsyYahKZ6Pblj/YobNh8UWsBC4+aKEH6wMl+9hpTaGb3P0CMfXI+v2uY1Oynb3M
`protect END_PROTECTED
