`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7mRHVYUXapaS5iDNiq2rjbINUbdjH6LJ8ySluxg6cetuYcxSyyKH5YKW9koFQVl+
w8YJcHYAN/xatG1BJY+H1uiDEc5vDlDXkZ8l1nGRcOY/R0xA2DSMr9kN+7JKxz+W
tfLdrcRDqBeT4mwLzdTYmHe41GmJQMZeYelyPgnpJYiyuqapE/+iMviHv1Hpyf+1
PJbLfSrDXNkYaBz6LTQVzWF/KDoP18Db2YTI4CzfI6mgMI58oKGUq8+nx1GN/d/u
uOjD/PgSlSGII5xWOeUxmx1Wt1FRMyntcHeJ4lm62az9Fhy//lRoVGRzt9kEhGw+
ASr/kly6NMZLPIWEYQCLIVgQTEo43h3RXIjkBEAuMJBQD1P5lcrtliGYhAMjrHQf
ISgp6n0iJm2Dc9k9J/++OUlPlKMMmN6SsZiqZtFe9XGelLFs61/MemYl20FIwdnv
Rb8Mkl1BNlmbMD7djmOK1PObpzADPaJFEL5OFKcuHgqv84i+bVACVIE09dsST+I+
DFdIfu3O4zIHDlkim1WL5n5XbYa83WMMJmExI0z4Txi1gS6aUDcucMLUfd8umjxa
z1v8v6ZiDFsT9O0Wa6QX44cDLRfBzL5OmOhvNw4r3Abo3i/pwp2gzMqtvYHP+b+5
duu6CcGViVBQKQMwYFGz+NCNZIjYfYYDfFazsRpHcANgn77QGnuUXMdtYE/fMLm6
ni1a0Ps/YrSmvvDYvrLju3JSUXwe1A088Bu6O2aPLZ0YhSdli0im2PIKgr2T4EO5
XmnOceKYkIa+P51t8KJP8Zi6B6GyDhV/BvJb9KyAuamevMsakgUSKPMo1fnETvCT
x0jMdBtp+UirKY0vJdV9q1CEDVNVoQUd+d5QDSg6mk8kyEhQhWEykU9Hyc4LJ0v5
eQIYl1RuANHZz9MWRuVLuz9XbOMSg7rB4W5rVUQUoZK2HSgbeGqnzOtIVJlfjB/y
Yx+IUH2r6ZUK3dLXxP1P8tNodo+Uadkj5rTqx0dDH7S6WHfsQZCVccIuFBLHKyi8
ha1Gdd1i8NbeDFBjeSmynah7JaAY0Khd82SSdNC+jfuUr63IPL+EChvn72TJcCGW
whBbmJmKhFOq4good1xPtacawjpMA1ODYRmJ6iHLAh9pF1L54c/OR/1D2e+DEr9i
s53fwf6R2W2ZInB8C02MZVFIl4x7nZPAiB6WYlHJMk0LH/IJAmeW7HQe741YO1mG
foRsPzE3b/BohbzJ8L2y8p24pU0WBapfYSL4YA/D8MVLqhjiGPZ6A+mlnxLTHic3
0jHwRhZB1S+HTPtFEp4E9x8+3+CSiDQRIUl+jaYX+8W1QvMMxjNHIIElMeTKUDwY
q3Z8bpi51BTipuHHXR3FvINmyPu4oL2ARiN4rojpUX6UAeWIaMqyDXgYGD5yhD8o
bfCroF9DYYD6bxkItFZGrfDMzp31xfHJswoRJue8FNLOzLlOQ8D2bEfEIThDm+sa
hdDjoWHAaoukGQHQd1aAyF3xIAPsalhV5tx5P8bQVRsX0QNFuEN5Q8W4sH2dpEGn
iDmtL96Rr7w9SheNS+jXI2rydBXl2X5+JT+7IzYwPQNX6SR8MFIzfSiD0NaBc/pR
7TJzUPkiSFiqS8W8oll+yJ4A9XM9sq7Qy2mvrcflv2vAg1lAsYcfeEAD0monrmUB
JqTjLREsRT54Bd6QgmQSGIkNgttyn2WlZVCJVPqJ9eE+ftcNH0IRAoKYArdVbJ04
0o5JhIZlssGIyWxo7+zbbHP0IkeBmyIdY1BLD8WOIFcliYiPPBwUUVOKnkJJ0avK
6T/7qJ+N246XxV7IFLbkCWQ9U9p+jqghCY+1NL1dTxHN5P0JU+a6xF+Dwdm2kTFq
bNn8K4dqoFNpBG8Q5aMIqBNamio2sATQGdFLGJ8T8FynnekyqiqXGmLojI2BE76E
7f17cyMs1j5DygELsq7vINi1+4MGfJDrItvfwkmDM4n0yZFWyN7TNOGR5tdgmKui
7cTPFntFAtCU2y6eNsgXXZHZBFcfIFAwmcPpBu7pjl12/4gMlV9vOvGB+DM9xnx3
z8jLwy+jVdB/G6IHFGYldToF6+zmUXa+5pzNuTftlOR04X7uANY1uLiKcNSVpDpb
csiu5nizrg9nH3ka3scraQTQOOfIC74CG4i0hXweZTA3OEMU58zxgAQIxAArG+eq
YPDkAT1pBNutNjJMIpYU80Hy0GZ4vi3KwBdya4ssdBhoIu5qvXy7Ka127XC57xQr
sqeeT6MJHdjxuudmURc6qwFxj2mloJJkgQGYXcXY517wvlF2a/Wb6W78ZbUyZepv
++QiVd6uTR0m+iSPLQWJiZsWpBhaEV1QADeeYVpdnos7oJyuGLraui6YA/+twhOg
ocswRxC7UVt4HEYIvgXJqw2mXj5jUGdXdvSkm5+opWVxYCGk7fuqZkGO8hos06ZM
QZmw5d+nHHQRe9FNusN9yjyv1OKIa+6ACQhK8tIOF2gIhI1RJ0YlAiD4L9joHqwW
ErEXYUae7rvUNXNnB9YSY8T3gos/j811eUSs/gNjahuknDooGO5LmAmFoGLfn6F9
pvyBv4WViy7x0yQsUbPFC1KdRyM/NIs0BF2Nv8UTvguFDk/gOmcJwsq0VEiNHVNa
fyexkYccZwEIhZ8yd3weA4xqSwZjcceFqkk5HsCDESukBijLA0X2Q1ANjfI3Bw3v
noN2Qj2mQRh9x2PHoDeWgwiNMLSu3+/MkV8Mau2rFAm4M5f0zGWdPLf1wopPqFNO
XRNIL9IHvcaDuWhUcbmoKYmyNDinYAqK8wngUSBj6d8K0sHqG+3wWNf8+4mo8XBb
KpR898v4QDnny0wKij+dwZI2QcI+GyoWNe3GbwZWzvFHAyRzq33DBFLHud9BcFxD
Ijq4oR+8V+X3cmYbIh6oLpII1Z7MGgP0iaHYTZc+7mnVXnIONr80xqnJ5gGigjW/
XQrIIPxp6Keh4xuNn2OplVH3fzPFJiPB+XQIJlAlR5Akdff+gtCPDH0vycsFysWQ
QEUQZdT0IIzuM3o4TqVVHJeiWi5d4A7D+TbB5ChUNPIlb7ZBZZyx7vtxkqfqtJ4n
1llicOxab7ceXw4HV7M/HQfgd3Tv89NkYj+yE+stZpXDe9fSEbEI/FAaHmqcUTWV
cKpOLf5jLWKjzj7gdlE5tSpvqoci8U2GviWWl3xhgRrB8Xm8Hs86u0KCC9YTyE9C
wvWo1Z9ZAnAzgwmSBcK/6GzP0vSpHCjcbBPDl+IcKoI9G8OuzgzgiBhSR+t30cMK
cQuv4g5lL2EZ9YAVXJ57pbYGfMSpW6g2DmZln6cbMCC9ZZtQRMTReh6BggsSdgLz
e4XQfJGFCJJZMaQ1ObE0PGLypj84BuSlP4HKT3Jbpgzid027LPPBjnPGSkEltFQt
W9VjrojzmZ/Ro3LPjr55AIF7dnZGeGkVjQlyhbNispz5vfgaXpe8010XP4QlLheP
L7xb6v1S/F5QMB8Gb4b37rKE4iwhxd1ymGdP6PRXz+PNIymtp/abRJYnEZZmBix5
kLFA06aPrrGBYdsNogAijtfs6hc/45z4REC8YRJJBISrEanOrNcjhHfZovD3TIc8
q34rw4Cr0VkvqKNlzVWZlqBcD9+eDqfcQmCoNug0uF5N7QHWd3inRWNZivi6eBI5
e/GfaJbqoD1shvSEFJPBeXM2nYnF1WYh9lCpye/s5mGm64rva7GJMSojezkO6vd0
OZZEpQSh3bBNqePb47nCzFZi4Y357MrKZPg9HEMJ8I9mJR7t/A2vgWFzgDUSJFEx
kuWF20Vr/dM8ePpiXOy8aiP1/jCW15/Ndk6AdtmXj9MMpqwghgjXS5MfuIlK8KxP
+T2Ek5TzD9ehua4vdoj6j61eEb69/jqdpBL0usk13+5TyGJ12UqoRmxHk75UG5FF
ZpOO6uEINDGZCzi+85CL52XpWTYHI8FnWQfx0mrSSNAcejV8ugkGNNxBrYW/YQx3
oZRyNS/mAwV8E8jSY8YPyCuq9JbtwqwONIut8mlNMxkhVqtcEpaLHkRNfPfsC9/c
CX5wkAnbSGuWPMva6NoOr8XpBpn80M4tmLzWtL50WrF/rPPEyE0dbq6DP8rMiiQs
TA3/kBKB5gjv/LEWXmW6XjPE+cCYymuWfz0ijg2S6iLlQhApsNTyWeFywaMsZCIa
zbvzGYAJ7dNPr78/GQ59NRQRJlh8PD/OMlWbFWKw5puEg01KmBhyzru8wgLytTwY
JAVZb3ZJMPZOspa4g53uc33Yd2tV2Q9jO9xIc+otrqOegX1aWuXd6/eAQlT9rNht
94Yte+C0d4rBzlInGdKxi7CZrvjtlC5dY44tIDaiDDoTPYBAXK/c7viujkd8JF+b
fY4JaYivWgx0hJkCHiOSHBErsVX2AGNYplVguxce1VLgOrfuoyasmzQX7anFnZMI
KDwRio1MxUcx/kgQqrq+4EpnBM5NUC+jIDHQLyJOCeVEz9GCOqctgBz4dzdHafjJ
RC2Iz1CJuWO/42LEIgq3BFrm2k3gk0iDVvzNKar455UusiIQj4GwAN+hie38vjTK
NdJcbyDWYwK2sTMP0sSNU7uBu6gyTYsQeFj8H4Xi5HlXaKACzPCLzLqUGnHJSXXL
BTUOZ5BNgatdauByyi14EJsqIh460AYXKGVflVjYEAGz6u9uVIJb/ZPndSvz2gPv
ugCLDrRYWGFdo5LiNrd8XwVt9FsVkPpFXuDb9aU2foMHafCQTn5pMdts9pgtp1/D
cQzc2iJnrcOUQQkhNexAG1FB0ISF2GIbLVcLSRGEFK23MnDDDvD5SPxwB/RbJdZX
onZG5qqmeEunfi6woVSnMlHBKfj0kW+IuqSvwi+xXd9by7iUWC04ua8e+HcO7eq6
HvNpKE3d0YwuKrw7mqjh4unesNOuqaclE1V2/XRO+IW8MBn6LOM5VM+m0Cv9lZ2D
T0yN+qCigUVvdJKovyyxlH31g0tAZZfKl4EcTRnJXJkkbip4nn5Z4JnzFZu692cP
fhl4QZ7XQfl5f7s+4Y3a1bgK7+s/cgYOj35eKmV4LeqvqkNwgHY3RrVz2T8IA8Ze
VoqiuMNCZGzXngEt5zgtPRL4LVxXzp4Qs1uDUQ2vJW56JkddbZnHVIoJKUjCDJhI
4+aGbrOoZIiMVVX3KmjHfrBqadlUH99kkc3Fv5Hq9zOBKW0BfTS2R1W6eOxRQ6rh
Ksvhq/c+6VFQSO5vs84beiySSb4grhdzHwMIjiDwAevsDV9wy358jhTPI8oAAZAo
uFmnbU0qOmBtHq8ia6mfWztommnXqKOhpGBdaOJIgNEg+7TgLfbM1MbWHnOKP5KK
rxMUy6YdFmfjSPo/VI/aFueAtW+Si8gbx+X9Blv+pKaSx+f6IlYyAUFbX+1hxsDX
BGCLH5g8oCHTZv0dQBZjdaTCre0Gqc4YeZIzwrAkys0jv5nwMjLGrnCneVtPsYUy
S946ev0wdWzyQrnU0gTv7Nd5tVhO/0ZE0HHHVT3ob36tFpYEfDPx1R9CqpoZi5sb
85gbtetTnFk+apxVmHMFp8rGznCRIJQiQpv0fAebll4gIzYARLGeDfiwL25SMHSB
vODVMd5k5Yi1DM2B0PJgN457j+DHYT3ILprAglplnNWUZINRYJm1xKlQ52H3cElG
vYbRPf/ruing0Dyi/HU0i9/74wbK4/RG6jNUdyQD4NGicprNsLp3BgGIuRyhfNFr
mW4vZkvHyMgOpe4l/bl6vlAJZ+U9J2wlNA/zBaQ75ZS1NeVlWgb6jinSqlRJpUwF
yoJopoFWlXL6osg1qvdHUiF1yR6jmIEy8zQwhsmOaLSvGcd5CoZ+lJbMJzZKxZvN
G1IjEz32Cf+8rD+xNUKHHMK5ESYttJknYylVLFJiE4A0c1FkGM2Agzxgg+tZJRgj
n5ArPpYNsT72ygtzduuCUE5U4fEKto7ay7h17sSDcdPJEuqPSPYQrbo1gcoaobvi
Wp92B2Gomy91TrZfa52mTnjtcb5VdscZJ3LbPvTFcq5N2FmEcNBT/t+/zfW+nftA
Z8lVjN9ND8pX7Rc2Kao58B/rNwSOh4ijNpd+kpDWZtnPWz/McnRK7vazNZAzhMVX
HQAup4WNf77IlQl75d3do41Ci62LQaWtDP0ORewSUJOoOORPNjpzkT9dWxPKuCrU
zH5Aje1Bq4NNupYK5g63iH27f27UMYQ752hoqHBkjXPD+0xJTKC5nO8k/iM3RvBe
cGYtdUOhIlNxBo08U7tlc418wQTOB2/9mCTld3JxWHCR/4J7CTtAcALTVKY3xB1s
iV/HNldt5XrUXO6TEpt5p3ubas4PfY+LjIQoix8jpeSs7I3wECtwDB9y229zI7+O
oT+z8iuSCuHUerBpdtaL5bE4Bu6dRXqmpoDNfPz1xzNDc5bOfibAHrzLr3MqYSog
dYQPS6a08vjSdmbaE/DC096wYAq4Y69NhrpJNPJwdPxKH8m9CGh1cCU6Oh8GbLkD
BPaQ5MiGjHMozxhxVqyMxliC4G/H3xQ4XaRhKABykbJicv67UY4EgGO/KjV2ZbNo
hbszRBcRvjiMTPyCGUN9dRy9tV6r8aBNRhG6zl2HPA4G4lyIliDvRZhANWHfJDQH
o4a2JDW1faj3Chs1w0VxRrlK207UdSM4hZ0PWG1a8WQ+8fAjIXxLX+oLqwmHNfhu
stQTBoDxnK8NvhOK2HPT3R+7wu5+PRc2Dun/vDyU2uKhPziEeS4o+yxdPXgDe8Yt
iyculthyPTwlPCoLhpCuKgBJtjJvR2b1XYc3zU5L2SHSzTYRe1q9y6YZr+av3hv7
UnMsfnr28BaWU232Ovhsqwr6zlhmrVPHPm2Doj2lmGu8FlbQTmWa9XcaMo0bDjNr
xyMqliu1cqBaYxzdTbY0bh4aw0Tgn7B3FiylKI9dIUfPwr6iammMDY7sLmmQak+P
fvQ+z1wwcua+iN9UqCWr2T6bguU2pvdNZ+Qq1vnkU+T5+UiU5A+bGw/vQ0sfpLSm
oJ/uAw3kPPy1+epEKx5ssZPKHxtj44RBqGJHhPsORyCczM2IE/3toapt8Nm1Fwrm
tlObiHre9PUa4pSJ4j6HmX0iGheq6oEgTd64gQKatwvCGHjwz8Qa5VP27VVuKDTZ
j/LhHL3qFpBbZ9j8ivNjt3fVe2z+qafZ0Pvkx1a5UqPMsicXBK72Xq3GKGcGlIXx
p+aamwh1dW8fGOrnPf35aNjOSsCfTa6lQt2Cntlh5ODe9bZxcirQaKddkXwWCIFZ
bDEYSLvD4C1Cfxoiq9KCFni1Ns7BpVgoZHnieFdLADG0iKL7q1FF2+MmRr7XPlNe
qAsDKpLX2TX/bm99i+TAAvrx4WTzpo2A1IW547L4pCb2yhFvKV6boWyJ/ndeueMt
SiTJlpBYYdx005LTOevnC6XCGwrO2ngQsSkFxoo5krlS+Rmk9q6A3utC/h51yrOJ
1STkK1o33XqvCseKCTVdx65AM1PDs+eArAtt3NfT4wLFgcd8M530796HYXJdLW0g
LXdzOz8acm9zGJjxB4BPr01SRWajHugojxZL8vdvsJXWAdsmC/Yq4ugVlw11Rp5t
hnOfUr6lPTNgNf9FxUj6MNKsPgbmyt8Yyl8tF9khT7V2dr3joNv4VqkYPJCMP68S
RpZHLQNjHYvwCQrELjfVtC21zUfEeh+D8tfnzjv5DkGMeYqnym7sDJQShzYj+N64
aLwwAxTH2fbih1ECLkny/vkdo+ueox4zPvL+YyNQLjD50h6nKyqI4dwRvDTSDgZN
RZFlFWHxT9prYLuj9MmIYTOr8hvQ7ryRAkITWglJgmt7rvjkR/PbcsisEOthqZib
TFH4SkNU87PLX5J6rmwBtkYFXDVg1r6gSqK9KNaQ/nUyIiH9q9GErasJp2BnKEGT
nTQPsmKwKrMhqhDZFKs234j2BUqgG5UpBQBYH23B9bT+6Je85UHibDUqsncjyuTH
Iilac8WfqjA3F6XmGXQzURpjAfxdCIgMxYF93xRzY7fGTXVgPGK5CVYdYP5HyDiW
JQeipTYUuqBeLVuToV8RI7C23LD8+S5FaZxFZGDjdYuqQ1aCpYLAQu3bPDT+OqjD
xX+fOnEPQoaWt9m5xRqW0Skv0DBeOyDC5q+wvZPQ4fnmGCqZjOS769RohIopX0vV
BXs+p02b+/VbU9VXrLCFYsgRg+Zgsz4mwv0Z1iiAqGQctwFgipUEunV0OxV00vOc
udO21qn7OSStneQlCFJWbu70B+gK6fS8+6o/GrDFEPyTLz7ngTEiic7gWq/YSrSX
6EQgzO8w3IUN4J3HDH6TcxgJrDHf9/W5N6F+yqZchiT0TyTlxqY0KLkscEZY+3TX
cl4tkPuqgJzQmG3itsdsgiXPj/p/eA2vUjWBU9f01X/JsVkAPhCtDk7KBo1BD2/k
G1X0vwaBDA7O/ubspVdaYFMICJXS98JsCjG6aeqymsRvuKcvXU0xeST7+Kl6xlZr
zycnGquwSHlY3QRcxkSrVMIbT/qzz2RmPUDvgdpefTu4TdC2PTRtM1Jm/9/AIthX
ajs8Ex6aEe1Zs7NjZyo/8MlOwO/GovonqEy4J8vhATC7zs5/0eoQ449FjT9EYAMk
otPTGU4AavSkWWb4Hei5y4H9k5LtBZz8fTdLluY8BCVbHH/qyRD4puuZUxjsAEAd
jnmMgvLk2wnQrol5yl01fA+EQ7kf9cEJ/UKx5sosRCfvNQig0risRSaLYBic1yq0
qH96B/2AKuf+UQGumY5P6/vYzthTnFF3hcZ5gBkPBxphbMe6s89AviNaUyYtlsL9
/3m+fyKPsEvlLuf5DMuIOlRjPHA2LMcbrThIRJS2yEGl4q1z2LzVSsjhXr8mVsAJ
fpnoS4PIUDAGWVuB0hM3o20togQsc9WnziqjqfnrWEy+bFpY5HrZ6PJHVVJPG50Y
lmCWXp0kghI+dR4WgK1K62S093DeY+6RFKcs0kPCoDhc/FsYjA3DAPG3IC5prMt9
dXRng6Yjo6rxSw+pmiL2/5JrcolzuiYFp6GNyyYxbYj2w0JqTo0pcZVsum01vi0c
k+bC6djxU1SQiv6mclBmhb/BqnAW9MH/yimkRiQvoa//m5QejLPMUgotdPDHcGg+
bqRr38i89xMRpAdJxkzk5K/Ze7dQ8H7aiainpXUam/PZ2sd2d4HX+gM31tS7SKTv
M/aWHLeYSsI/fR6ydgEhJbqwvo513ZVIuN6XOz4xiGhdhQSzLbTNFibkfhZqtM0f
2mNQ/Rd12of+ff0YBY/+ElveGyFSS6mIhXXjG3LlU9g89yIr9ksHE5OSEihN1LEB
5c13DEnfSeaAVlDKtdm/2KiXrU76jugR/g+r46SfCPHaFNH7lF+ax8dLlAyESkeW
oHQ+UIkYZYZF/shyLGhFUuGCwu6WH3P6+4Sr12Az87Mso4pvk3ilCLIEDuvJ5O8A
K5DMaMVqtyYtXoznRARWT66ZfzITB6WZMkb/AFB5a4s9h7OC8305uFhh1Fk7C1Je
KZS9o0xK+0XV5uwp9BpE26xl5cGl8DFc4lVz7k+kyDurYRs5sEpWmAIoRS7XTmm8
eTWmAB6if69TbJ0IoULETgvhkXuHQFL7uF5ZQt50L5Z8euhdpUMdRqc+NDGMdbRr
k2UDi9MSDx+Mr95LuvYmanEgdS6v4WdU2J2MdvhNMrDEF1/1gAvwT6yQZrMI++03
2Xv+Hx7NGGZudTXyvhC7tULb9HQQ7bkvyIVfmMIkLu5JiQ0E8LHTKWXnlGistNSp
sNSWt23Q48fDfLO5YIQSwA3D4HJU+shqUxr3bb3FZYq1sXLFBJdGw1y5mWfeJ5Ld
EJjh0IN5f7qqPMrq9Rm3YV2weFc27INaNkcd3d/CZIgp97metau9MrN+a9pd/yyP
iN9VgYECwt7z/NW+DQ2e8PgnCD1eHuq5yWzFmM2fbntA5Ge4crhb/vyITW2+4Jz8
QBkS2gs3Pz5+nuQ8ZDAgxmZ/EpXc4eFs7UUTy8oBDjZxZH2Y/bQmAyvk8rK3GSw0
3zF/3+UST/3hxRBhm8EtO0KpjZxR39yZAqWp+EJ7g4Cym+oUYxLlnWo986z9DC0A
H2z8mEKWgnAIV8r+02RZRGea+DPD4cQi2RudcKVKUfQPnOVTFunE2BWLKFUyLdoS
XVssxjbmeH+0pgAX5BbkGDKksdWyYrNlm53mf0eev6iTIxiPpSrEl1drIivA7QhQ
FWbZfV9lrIRVYds6pw5WjQaWuzqFjPTzpFdOEfuyZnEGJIYy80B+ESGkr1iDVM1o
MCisXM85+1fXo63AwdyUvKLYQUpc8VCAIzVDnxrnYoMCjL4N0oNmjTK2xhK9Z80T
Y4j4IofnG97ouTdzWHn0gNG0zz83IPNnirCBC0KFUAD31oh52LOt5fMpSZ42nxr0
dxA6UJ5HQIXzhsfQ13GT8RaqxYdndLv3qxur9Q3VMSUBUD2Ug7HvgUGKjmWVC1hC
ii3Kat8JJGn4H6ycI6I3/e1RaVtWBav4VEdvnqrNszqWppGL1VlZUljnlTa+GhDd
Ccz/QRiCDim2724+avM+W135Z3gUbTRpieMnGw+pE6OwoHeJqt0cZS8fZkkg1hwp
XAlBJ9PcuHdqcQ+/Qh10Ro7VcJcZsKMEpZRuFeDRojXzxmcff2uL33djpmkMwVHL
0HQW/wUh1HQMDyJDttLOxVNIRM4UOiCg7TZYJXDvXLlFh8cAKcxC8DMvqp/ZCGlV
MnVqcBb0HEd2UE6CNYm4G4xraXmDAjfY+KqYmM14zh0yt4FDf8ciJCXfzGmFIvAW
jXa+bq7fXDQms+w0izeNR1w0lABzEWp/AiXh0quWo5Jz4WDhH40/PyK0+gX0Ckmo
sgBPvd6T2SYX3EsQwJPeHMabBxtXEnb9wl2OCXQgwjoElEonrdMrV9OE0n9AyhVI
3E7QUdInDX9Z1Fp1zvRVR4ECrBKmt2uvO1I+mPhg5JVkYwl00VyDk1F7fQloaB4e
zsaJ4H1uJuXk6G37qsSOzIaFeAqKw+H4TM+AG18dB/g0FPKfgqkTSyLmi570Gc8E
TlhM8S7TKoMSiacZ6vW9OQLVrm6+ueEs/Yun3p6750In5r2EXWbeLHrMFLkyDg0c
21V5U6nFch+OeiVKgEdCdZWiID5RlMNRjhhezclWuLZnRPmMciAHqMCc5ivrlsYX
jUX/FIQU/jFMFIwiorIqunPHgAOIvF3s8qNrKq4zVomTucHNRsIVuWWnN9V4pTHs
sumtajQ9qsOiGx5EZW2ohNJXCDe8ogXx8IQsvddbOQ3U+x6+55SESEXzKD4G7uMl
m1/29q9j4YReFo14plWAWKMXOU6+DN+6zPrb+l4M1Sq/gJLr5PKf8XJ8rFw5ukML
7sUWbF5gliO7wlkXYzcmlGdvWYParhlDQwdlh1KJ9mA49dUMx5gNzgtl+hOOAoTo
MJeFuXKBXw9WLbXQG89Hv4D0UUdweeoZeNybcBpk02hXG+EOXdbCaJJNKcqMpk/V
zKldxJHu4AR3f5QnFo59lFIm/gir0UHWoy6YMeY7UgOoJM+Xv1m7DLzAw0altyJR
iIGqw+EG7UNCGuZ++lyoPwQjG/wULi8Q8wFJKEGPszGTctI0822RUNe2p/A1GZfe
rMPMFuZHRYN1tLjJ4CkLTHuEG/4/QpzOG8HS5lUbS4G0n8Zdd04WAUtMPINfIfdw
fcaYHADLSBgoAQN2o0tdUZePr2xXKqNdOqBS3eZ+1j2LB5+hrgwYGgh/sbAJOnn9
zeJfdV23jSMrKUQ6uT7F3u7BEs7+MrZ/MSudKlDkV3Q0IMFuM8tNoMBuj4Z7Oxya
Ar5xofPQxMVj4TKTq52VqQfQkJbLbaCaSOj18lPRBmna1w5kkrmiRdzenBujxCJe
1Lj62P2DjcTEf+YWa5W01TFLEYqqUAeezYcNGRwVdHnhA6aCBH8wxfDdgdVwd6OR
p7i+4+8WEVI5SNi1yaN00BZmX72mka0/l7cgMlSquxgcXIRzHx1ll1bbyvZWALiQ
wgYpjEaZNbZUboeYvIKRgscC0+EdfUXSiyFk5b0spAXyyWKgavB/xaRnOOrbqruF
bg2qq0bMx42JTmrd/nH0Fh71GietWjXqppjyQxn3n2KbEd8ntcvIvYemADnOgzKG
gIYcC5Khpm+XU2V0wiiS08Yxvr99zgln49KrLzUd2VddIi4aZNHh9dWY2xw0UABr
Jopxta22rfbBWKKPdy79We9pvYo+Z58Y2pYiyTJTRvPsl5dUjU3MQqsMK8FG+F7O
nCmxiFmYQRDvVsEtz0BHk2v5Y9JG0Ba7yFG2LAST6g8YDQvPXhocp2giNcNbJgfc
3yPgeprEmms7clF/4o+cHzFrNXkvFpdNE7T8X+wljW2zbsqyo7gJ12Z3DZxm1ep3
sWHaAg+sv8/h3XeceA+JRtmo8AAwgQff/K2l660f5KxUm9IOb/9ikDVHzlSy7hhr
TfIh//mU4y2FjMo00pMuFdjDOm9X9UkfBiqE60lYMqnj2pVQK5M4x8BroJWA/x4i
a3zokWeOeSX5ZUQMI99wtYRqK1ft++edgfBqRQSKW1if6shHgFTI6IEz9+jJYwcW
IozDhfWQ+TzyrD+5eWzduxJLeBBZzrNvp4P5vOQyYPtc73h+zAxZo5ps58W7IFWm
nirrR+rABeFEHVVoofc4vqUOSRCQQjHAr2lZqDvEw4PTl3YIhUf7FM0BMwAitf33
gEqJS6egX+Bit4VeXsxXTcYDyfaKdANQ67xEuWBLtMJ69uy8+mQIAOsTImncuuQv
32Ixw3Q8phkYC7IDMouKDLEYhInMxPAJDkVyHRcedMxz6mgk7X9hZpQJFbOLsYid
rl91X1PNqqBCodgxOZ7vu+3KZwejzQsw+iMgtPTiHZhVqEC+TJSxr4JDhHz4F3+g
sWRZYfIcbfWNG5+6gACwRyVIXop7hfx1AOYTIrFhx70b6GXhF5aQWfc35AUZCOYo
8loOzsEXMz4k+CjaBtxoD17WwdDP2FCGNJifbRLQthG5zo565/kYE+vkXVHdYqUZ
xpSjRDg8eL28cIndk+uNdCm9tatFELRCIs6xeNJSzuY/Z6BHabmEMD5c4nRqlSKM
4NfGp3APg/k4TNs1XT76aALg2r9xZNW/oS483jr8ohe/zAjUvJqsnH4+WVz5FiJo
CVEGwrO4roFmvkZ+hGvRHmi0VK+r+cZr52Re7N46AzLY7zG7fxLicb6YqdE15J1x
gPH/QMzOTKHByNT2kUk1Ot4bXjhKZf5jkTzMKdsg/emubGCdgw0hzdtff8vQjn0E
s4RFdmjuw4z+nTS0E1xVU/qhrFKvtHs7bR4/Pl+esy2RAZRlVI0cd6IiT+CYBVVZ
gGpQRbBgZDmyHJvyne9WVpIeKVYP2P3CmXV9RGJwaVOaN7YjrjDLYX2nAQs22GKI
9ITL9Z7SUHtL+w7VxhlyVSkYB19Cug3oNnnW2/deSbNKUroHGQwOb59DpgC+VHlR
qo1nVBq1ZTmUz0uBeI83NZvGPFlbT8kuNQ+3VPm51u5Tb2/sO50sDnUDKLSv6lDk
rGyHen0zUFXS8lHTQCNnHgLhDIbS6aTeAxNlhTxto90SiCOsRTxxFinpDua3dqbL
SoQrNNcJi5kYKuepb9Iv3/4JABI5g+hBZtcFhm4q2+wMnfPnGSrbYoWEYlYsnl3y
Lxypw4tZltrJrl+ZW75/s7nAcM+Atm5bUFrWhhDXoFC3lglTe6IPBRrGf4GfbkWF
kwx7r4uGoSOByEMBcR+UGRfp4ch11hZ2QA+7YgrXbDC+riZWjD3NFD1DZTP2FGix
T/IUs1Y3S2nA3FUhFteWs1QkQqN+5SeY25Cg96krV3YYNZV9DLo4O7cZTeLw/fjU
i88WOEMQgJnQi2h/l1V8x1Y5snbsddNle0/0wPpNx7byFF0YHc6GerpsV7cTQ6IR
DllX6BnDiSJalK6TtKT0l/Zg9HDdtXwaoWZSUJ0i2lEw0VSG5iuD2SbVVFK8Hkg+
3kV7Uc+KfvZzempJsthyVkeo31o6jrCVGMJMNxKKdMqBy57+PsibBVMAmomQN+Tt
ZPVGVUhwsP+KwGy2LMT661qzmx2VYWUeVSvIA+ZJoWwqb1vV9RiS0bkYkNJKHdIo
/CR0e88YELnKGGVN0CYdMZ9sCHoa1b7G7T175OO3uWdo6D630Uonj5oTxOOpMN/a
uX5qolg65okqWzxqDNOGFK7gqW8z694LwXOcB2n8LWClMh3XiLXhiqQBQC57iMyJ
+H9UiLOKHhYVsuIIiqK9M0gKHSGKB8hTNwSOVnSH+cNbvNEo/L+lMl+H6PzwxY/6
b729kViGTV0WuD++SPJ46ISpfaP0uZSojFfEsGA9Ro3a0CM9PpfykoXGG1PclVq1
A8S6pbu47FV5w20ZbRiYN90qjQXwPnkX967QxCygqeMZMJ13BdyzfLsMwUMKsA1H
7DtvTmwtbKzu3qHbDYZ8nxw2M3P9kLJj03hjfIDa/MHZDtDby930q6lhLyHGrfZZ
0fuwpuzjI3ZqImm+2etKEzewCFY1AEMvoBlzxhfvNyzs2LcTD8e7GQl+7jLRET78
qJzp03VEk5Wenc93xYpzwWZ1y4IHPWE95MItTqVEZ8jkdPuu+ZlQ1Q9bNxXPo2TK
SpAeX9bA6pXErqxpu3fQuShWPIEhD/VsfKGzC8+gQvJU+bGzT3MDacocm8exXClm
7+012TvPTTVQw40a8crashYR9qoFMjlZHU1CmbCGsUahjnoGkb5/Pai2155u0crZ
R+kbTfiOOZPQNYpgR4JLmyZv0ZiL1svZqM0c+BqlmjTVwskwAHEUqzNmlG/Z5X2i
TOC7ePgvxoOBFT1Cvc+nVnxWzZTsfqbZ4ouROLquV+94bQk3ELIDd+8k8QpYFKf1
REjopPdh8h3+PSW8lDXFka6l7uacROrx9LhuCQTrwIzhVnJv4Q3vg6NI0JYh2/tS
gT7wblqLJO2Hd9fhahcmrjZF1vCQyjP+D/GED+M7getWx6KDbxcjFSWovmCxfIe+
uyiBz/OXfH0GzssN0URsAfX+GVJdusxtCtD6h8TELipWt0HM1j9hXupeOr94aOW1
1p9NIEuQqMAhw075HaLH2xYjspTbwg58xRG/SPh6NA84tAjHk7g8b1m+upFt1MRy
HAfVTCckCA+xT3b93B3zfJ9JCsRka4TT+GC1XqMEkDW/zY1XMcp3oAi4dkNIAsLe
2BzhZjh0y40nDp6siUoB5kwHtwRBmMeTf/np6i39gpmOPKmnAIA//JdPPmxnC1jX
ZBnK/5XikFFly877qkGTLISphlfo6HeC+WCT6WOQeQ3wgOa9Mui/PVoPCpn1/VTJ
Cz0Sw5NSPEnRzFM43W4qbbYrwi7yHn2O5odCycT05prcpOC+n4KU7pi3GXdTofoS
cN10HfGVgID6lWpABBIlITdFlVQ4EIlDn+H0MYfK/JcrDDuipEjMvdQBI3Z4dof6
6taYivhvzwzuYRhfHhmsIFVVc5JbIcH/OxR+0vl8fUY9RAcVPAO8GyLAxerl+8fC
SxwwWq3QBf1jBOjzz61tkdEl1yWO1tbsXVxSLY9Ux3Ri9nUG+vdqnoGjGMFrY2O2
83/5zTXTKoF8a/0M80OgvpBXJkxXTIBZaDc6q0M/JHCPTEvnxCP/Zr5xzmjOIcPM
ewqN4tS8W+qp4Z1sGfp0RSyiPj8fwMG4+Grz9Ss7nZS3ntASGnAYJX3eD7qDwtG7
+9Ns04p6fpHXW1tAs3LwYJJhN4HeNdAyRNdt/g0QZQxrZsgcsqHoK14YM7QiCKDy
iUn2kuP5rTPimZSmKdpt0ivXj05owkmUg49U23q5n5BG6HM67l8KRFIpnj2Nyjtr
szWPUYW+Y+ViG8xP53r/QMQdikm674WKfkoczb5g8z+JZOJmQejsQqisIrPGKxji
IefVYHrp3QfSUV1RAIrWIeYdpMB21DvFZjkYHSh48VwogeyV0pkmm5P3DwfpjLBC
d2fP4S7GNVekdCKOs6hufeyq5sPPmSJfRJ1OBJNi5SobxNmb7dC+G89Odjcs0kTf
ELewE529yMXXLOetak2MsN6Tzfdcc84W3d5V8gE0hvowUeFRKu4PAiVNR8gwAILO
QGBziWXHYqgOFGX6cPKFBVAC5DO2mg/xdEnlYyXC3X9LkGkqHAdLvrbRCcCt/8bv
v0A+ZEGI/cIgoINGmbtLDjVvGWJkBLbCQeFVNmpuKX/a5bo+CKqIpRpMog4M4X8X
aGWFgyKzcO5m0yVF8MeZfH2tLVTSp3MJ31xUk0XKkuC/6mypQ2dHVnNizHQbI1SB
YGDZcPHss5gYuaoDwBn6jF2CxCEgvf7i15mrlnh37j2YBvhjPJoPJYa5Mv7Qxaj2
KOoAhNptan3atfkIzekI3jiX01FKov1id3W/iM38a7CGgoaGxJrS0h5hHoHcVkUV
hcFXInoZunR5QIuVUVRRky6Fq4/6mzMAB24YGMfwVQJJX1mJVrYi6G6W/VJjRA8u
viGv3yt1EeYPg6ajTZLwB0vCMJo+euNkoE4t44TlZHY6aN9IZD6Q55PqQm9x+eRB
fERoN7P29ZBBkBznpHyTn3CbRKhLVA8TsbRsczmPcNjJ9H5WM9VxdIFwwr1kNi3e
MOnoV4Ay6BUQZgyE5ctdPeOlYrNmjNOS4VbToUHzKiRduIzKAAKnZsnch+rcHjDZ
1Osaf5p8T9doSnodThNCDgwb75niea0aUhqN+rWl3hy5E3duaKRcae7dg+GZn9rX
fSdikVOliXFerVRJMKu35a7M1ct86Xo51J0ZQpSbAIJWMIVIqiX/RKMU26R5DX0I
fj0cVUvKgOSG2XFaX3zUi5okxyu5XcT1Rg66EcmqJauuRvekxIjeySbgBZdNsYmo
LhngWVxVcYB/1nOb3U2DNtQqEGz/pLPiOOcva1+QyYV51jQDSAn5oRMJ4J5NlxNO
LQfW8boJLhp/Hza6Ry7yN6P6VAfd9C49AGoQiAz3ftbqkW6koEh92TkQcXhjHWY5
355hJfiyKGMTyFDv2FTfvlpYCGnATObYvaimDNKkvEChDXT02wBX1koafFHTkKmZ
YX4mxlEtcBGh51cGKTK6jSq3eYTYncWeGtX0HKqi3hWdU5s1jrHoxbJ8OTd85wPu
8H08NewxZdiEOgxNnET7YbkFRGLebC+yeu4A1QpyEnYpulnsOoCtGVB0EBy+G89M
pCjS5KgvgVKGi60eJvYIhVfSNPfriMcQtJLoqp3EtyjQBP+q77/1iLz0cUSvcYir
QF8BJ7PommfP0AV58j7IhZzG28HRHR+5bwGHCo1DSWydfV0C62lwK5dLFCSJbs0p
PURjK28Lyuh8ck2Z1kty/Mk4bTwPJC4TU45EWGS+b47ACeaG68sK+8+KqzQ1Ff8s
PDKxd1NNH9YDdHA+5hKRo+FmY9OCKjM8/6B4nXHDTXTg5qBWhYXbT9igdMn0iNW7
Aaj4N6EJLfDOc29XpDCqQ4XeA6oBfStgos7MebFosne67jDV6So2ltWlnYkgBrId
0N15H+WCvJFd5je2ec+2NRPGb9h+9ulOoXcIYtV9YasrVcAy1Xk4FQ2IBjB7EUmx
yG5DeK+6QTaijSBuLC2/3sW+PGm5fmsDNYT3IMPbT/YNLyaWbcbJZyzb/6Z6Gv3G
vEkaeRlntAZ/f7wMuQf4sus+cfyIIqeV0hK5lw+3tfjB6RaVBm3jF/jrulb8xhwl
c7MjvoeQx1Ak+Ipl9+OOT89Roz8J+pbxQl1HYfIqoQEMidsPzZ0n/0J5sGxEHJ01
rm5ektT6f6PqASun+mMRethG7ACudPozFSqci7Q6/Z+oVFtVCASieXNXw8mFlC7C
t8blmxGe1EGODWTrBPIFznJRs5PaxvhQmDEH4lO54copRSX3CvNJtRgG4U3lZACn
t97GQEIyvLJ6DE85qAZjjTs2o4UtqIT7dgRMWOOguv0=
`protect END_PROTECTED
