`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bs68QYTZ1pECUcTSxkblwt7XbjX+In5gmO9UOsH17qEV7L8p9taOBvDK/dyYd+tU
u17oHZVGRnXml93jCo6uTEr8BUl3hD3Ef/F4v7XLWle7o8YFvmHwFFnOYXjatYLc
8VoWwqfCVBLJhC2zVW7g7Mj5eD5uSeW777dQvN+kEIJvBia09aOjTV74tGLAnNcI
vHU6H5mRmGALlNtrxcFQxjqE64c9IquvDIwIjh8JoOa/3AnexNW/IBnG3BHX++2J
uHx3Mg/M2lEGlPEjJLzGv7UMwuwfFMQQOx8hF+rSD6CMFAW8FKQBUjxGN6RC2YH0
VH6DleFyfTiIgqIr+GR5VTPoF/WplfXv4zyNHNJ/CAsipbqqi23+XcyYg0T2ByAa
/AKgj0ts+/neCk1vjAD85AgisNs9D03mfSDsh4xpPIJlSeQ6PeVgOrgLL3HG+T6Y
hrswnOHeA5B4Hy2dlYE2Wj04gbqpkoV2zrZieviOFbmRBWvAkafgtJi1Riw3sDUM
WXaWhy/V9/yu/YgSWc8/Ynt0t0gwrDxCWjKOsRLsju5Gf9ovor9SSt4lw0MurrI+
5cgNC2Eq65bDTCt4nD4iQsE9rhewatpM0j74z6wYbY/SGYBhzaywQu6zyWAgyI2L
nZd7xfEun+Tle8tyrY6V1DL08CF1ROQVfm7MEfVT6W9yle6I/JRqiU6UCj5rzRkZ
Knsn7+4y6vWSXiLoU8i/OJKH5Wc+tOqbkOHE3j1Z/EGcdpQD2HpmWzShE3cRoO0j
YID54A8f5QrhKS59xOhAYOla0Gy6AspG+Yg/Y9cpLkHTVpKxO30LFr+b11dpfApX
SyOCTdHtaUj8ewnPjtdgPgRRBtfWfsLbVVQNgSllm07/bTmv2BDAk/HudcHhqJ0u
1NHGoDF4NEk0Xcs/sNAWdiL04QFOg7iWrr29moXbkuYM92Ocnj4LLMW/8rkTyQPq
8RzNb9dj9Nfm/Tqxeq+pTehCL15624qGwm3Z94O6Y2L/snOTuG9KdXXzdP6NW62o
oz0oIAlI0VijPTb/I3HRIzYwwoBlocwpt7fBvK67FVJGNCMkWHOaKvBSx08XvzuM
8qHMvlbYmxdAS2zTuv+LH8Y1pL66Z8XLfewrUJexSE3fakuxIRr+mSS9RFTgHaJf
xCtMpkjeV7VIhnUMQP9uvyp/nmKFve8AuzJq659KFBhdCJyc7Qn+1LJXPt/Vv10U
fgn9EDze2h3z/KRP2VHVUeaaADyvoSvkyBowJ2SaPfuXWdyk3I1uFYUYuQEwmAd5
yzN9mq2k5XU+mr4qEspEK3JhBqzKvHGzbB7RTGba1LGxGO59iwQAgFyTgEHW/u2Z
hUoZELYx6kMHv2c9VlCEazt9W5KPFBjt7zhZ9jnn0k1AQ/ag9yl0mgjYNnQBiyNW
LXseHPzZRSDxG/efXG42cQ4hkZ4GHmSZRLUC1YZmgCLXoLIRBuQtgCgBZrZdSgDQ
ovRByDM6sx7a8Z+bcXCKULZhpMZAK+/fLxOWpT8oYyuhK3JTFblu4M4GRIrTkgxm
nBq26n8IwnoffycuWFt2F19PYY4XteMARSWrIb4JO0hQvuHgbVlZPW1oNXiJNs4j
G+R8QOa/SiDItvxk0R2nYv9j9egk3R3inducDh+GXmTxNnIIEj/9zHS0Kp/GmXeo
okvHxdo3uakw+7h2By4ZBOJVzWyi649WazoLsypPd4MDkMV/9SrLy4i7F1ksF/+F
ovlRTro5jfQ50Du0sotZmQdrmIucGp1gXPZSY0ZDipC6XbKcowRStFX+XTRAn4Dm
ysmGb7eY3CusZYSSjK5HgEwnNDvweisYuPwiJQpfNXZsbYRD226L8Bty9r/52VO/
PlGYa+APwg5qsn/Q4xSedCW65cbosIv1/fbbOXlvc82ELMz3DKqwoZEMLUTS0rms
U8E5Lj/oJymn6lRAMnnvlTDpjf7kKsW7W8Fih2aECcZse2CXjDduf+mByGSFA2LB
78uUdBzUy/JSiAuHzqfY5dwc1NSRMZ06NoIxsNAmxjR3pY4MWYC1xE+r1qQFmStA
JjfMPfvAkmkupfQbkYvZD3BHgp6n/PTxNFaOw36ZhbN/L4wbH/6wh/fHYQlReI6b
az9kxFkX/9Ybx0fYWCU6r2mrwzx8rmBMBrivGYOFbmPNB78dZjDpbm/83UBFO80o
guA9PyCoTSL7p0QIvySnMbTAhzJMvueZ8iKupj+ja27tfooUZ7869LGXqX1xpbIG
CmGprBu1z3HGdg2xQhGnTIvxjtohZu1uUlhyssIPeKveLFJHxTJAFdSxv6GuZfBQ
eXftGcpgxjriR1Tjwf/eAUyVUzCMkKOebNHUvpdr8j8KUl6auRyDfdG31q8scSQZ
Md9rJ/dor/mBI49n7GVuyRaopYHjQfepu2RMcLgXOP7ReQEncyKKevwOS9xfzyDZ
66WZLf9G4QwX44+HAEIPpi9SmltlDWymG5x660eWGVPXOGexn6TZvpkfbjwrhcNa
Nl+luJfq4MwhcF6YFwJPNfto/1g1W/1E/uaqtn/S7fi7VNQyAwUu7VrFyMQ40KH4
VDWLF4+/nr/D6qwaJ7nfbdM8wr8qOJEDGUdAyycknWyhFvFSrnblLIHOSQA1xA9P
K4TZNjg/eyf33cTNh5UfCDiVGTkYC+RluLSDp8H9mjCo4lcOk1v8x807YPftI/eT
Ujv2y/fvkr8dSdKBKRdcQfo46pFnGj1Pt7y8UB9cJho0z2AJTWhHYEEBG04Pcs8V
QDtNV9LrcwDiJH62niTW5BNFUTNxYvZXQ7SRDZ/4obJPLSrFPTHye2mqohs1HJrx
Xm1VSjyF8pa55U+3eaxQTKVms6UVr/hbOou5I5hCrwov/376Ix2tJ2geUrfVDXJm
ox6f6rYqt6sq3D52pVfRe3aG+MHdcs4SlooFDGfZl+F8XUgL8WYE4MtnANTTp6Yx
f3bYCjQL7vh+Yk9V2GrtVDDREB2FkyH0zrJ65lxw8HuewSpz1ef66mEozpC0hy0c
6873ONqfKFRRHV8Tu0F3hRakpiWYJ/gAIyZS7gDvQAMRj4K7T1+v6fUHXJDnLrkj
wIgdMXQi7XW4XWT9KXz02ADqZOwk2nU7OlDYPPU/VWz7hgGOR9lA/sWhhAZixC+a
MXP9OpKfZEAr6IWQ/4qB49KOp4lWtVwtZaJ9ZhjYny4GOxb1Cjcu0KnEoOFIigYs
7etufqvgEphX2stlkMROl5k4yQvB/a8juq2OwJk2zUL3x4szUdUwLMspBdxmH7MB
FL87jGFbxDG2BwNrsusdaQKDaXYQg0GklgOH8Bwe+LYsYej204Y1QssDFeGW44U0
GDiiYKYnbLJzpDTwPhaRZY+E+8fUFZQRDxRn610BFWrZxQRsxXA9XhATJdH6DoC3
aNYyOQczpoWMPg9VANAw0IFft4RqJlPLQceAm/fVuuXfdkbuCFgrNG4Rcjy/pPA+
aTX5pprOyOeuYYBE1KuTX+ALiotkJA94ccuJxRRXikbcW0cA7TDO91S6iy8YvKuN
CM7hNwLmA2xWuK/jl/khJB5al9dhCp4IkkDn3w8RW8yxY2F4r6Fm8HFSyWk2T5Tl
Zz43EZnTbLadzIXGAtpk0Q2y/JGItkFQCan2Ui4W0uRGBLoxiOc2graA8WyAbIPf
6nvRgxSgtY/2hI9EDolsmgsbSwpO1mH/8Ox/tksmG6nJUV9z8r7eXdLBg2ZSfSTQ
tGZOuyyDyqogq1rSqD3lKksLbX4AyaAx2KVg3hupyejTFXgK4cnmx6Ij0NPxY6TF
0fqbQD7bPoWHDsnKOqTebvDXtrG05v6mbVJsbmmzIb9Bt+QZBQPWf+6NEGDNv7NW
OxYeraTB0wbOjF0j8dVT8W9HDTBlzl6H+jKzjrDi9q0qbOGEBmw/HMVlsJdZpsF1
g7Uq7X1pMl++oN+QBojl+fAaFfiJhrPPezvjxUsHc05J7ZcSZ8lXKot6BN2ys7TB
x0ZCZ7cEyRcz6JWKA6fkI3l344/cQiKqmPW+w2hMz67yEds8Me/XFrbRtgD7hDnL
QJZ6Iav5NcMGqHhEdwMj/TcED/cHpjxEdccdPHE0laNdWtgNs245TXI9eMVxKkhU
lUB1RVK6KC4lII3q5u8DCUdPpdtZJGCrzlsoipospKuOQtRfK2YWpnb32c5DwqdD
63xYKWn6HplEbYj823z1kFgdB0zjDhGAj44/7iDYyWKEHbmvX4YulS3pgEHuSHAJ
luziKzBSOYlw7zzHpRneR44gKkoNU8apgAhxAcOuqztnYLCaP5FMPCKGWQxwKlw+
ZTYa7rKqBo5qMK885jp9d5IXIKqrPd6iD7VNu13k860nAYrsjV1w04iX93G7pUqu
T5QSVKI3SEr7FY48oqBet/5icnRH3Ki4hUMpURcfjIyWMPejZ/x0eGpfy7ztJlsN
D1FyUWLJLQYnq4Ra4ZVXsC/M13xafj5gqbiLPOfXHzp8Y1U0Ihnb2LkfgDkkKxu9
yWsvQFIgUpETmYkpqHi8jXXNNZQgXfE9FYHnucyEtc4ROS4SHav+QxEsTISCLetm
Jo5r/4HlqVBZrZz2BF07rbSonJrcRpQRrrSL06PbTeD+kkhz+dIZBndjUDqpQDvy
P2ezxKbThhW5U33mGMBhPqbIdILhk2ZY3wbAEkxWnduhIIn4s+3U5ZxOCFJ0eMIj
tW7Tj5FboVYLPu3q8mPNOSIH3w/KMEEgqM4a12hZ0oS0NO7z8YkVdG1IpnMHsHfZ
oixX9C9QDwE1t6QgIWo0xpUPX7d0d5MseTkRoK1WsOPTPT5zKbgTUFBuxsTRE5+y
iGk1LWeFQJPBhpYS6y3ZAOi0zmg9fSPXM6thgc3O8wUWlHgE3cChFXPRwFBGXvUh
ajtTjl4d1DXngZ0RCZCDaFcVyHetryYU92rplJgVTqjjXIdhjT+nC6pFZqnAEMMw
YnpjsMxc+HNnb3RH1vgurvAwxhh5lF1lBmoy6d9v5rkLyvxxhU+yZBw9Z6iu1BAH
wAOM3wkoTFdjKPy+4H/Wsn8tkcb0Ip1pPnBzdz62pABkrHXhC4xzeFq6JOKDFWfY
YrTmCuxDYbJc7tQMiTud3nFx7D7gZG+BxAzHQkTNEG23Leqimbm5nctULJShIqu6
JK6LEoOsZiJGqjQT7yC42+6NzIrfsxcvT4poW8VjXl57NjEh8z7BH8p0pCy8rQOf
KKeCbv735YFPWo7zii6nd6pWRzCFbCgjpaWQzg7OyvxnTTzqyITt4/TnZt6RFKpn
zpQ341gPVowK7MaRb0CFw2odBGArQMvXcpWPKMmJtb3rFPkG5TxKLtGxBNvKTGKV
8W0vhBTCqzNbjPwvV/S/CEmZ/VHaCK7ZS1Vo2Xj2QCZsaqPG73AdamMvzk8f/dpc
/HrjfohlvT9+yTxu+ZkJcn5ozUlBt+xJfTxuUxy9IvGXzcwQCVJOxie4hn4IJLu+
qY9T+tiHQzvvh9XOSaO3RFob5ZLO6LNU0VjeIqlqqMXxxG43pFyaAVmdHW3pbIOG
rQ/bwIDuQCMNAL0r7uxIs4lWhc8luOgi+ftsicXKXt9l5vKAkmsi8x4DOlPKQTxY
AI0EwtPFttxV5uTRqDIjk5+LqdHzHMw2duO89U4T5xvckj8r0eysXAtp7VGF7Ecz
k+jSKYr18AIpAhefKWMnK3PZ4kQULIpIBxvUghVoA4gmtWH9qYYlZu0nHHeAFfcW
RDeaEpoKZ1wsqC9aWgV6GfA9kO0y+TKMgIkdpMMRLhdty+HEWVAsoFTUvNFNrPwO
LYoY4A0AQQQHD9jmOYwRoEO+5yAhPUt3GEA4O5r50FGq2o3OuGnR/IzTS7VHIO1a
z8NQomMpXH0Y2B5V81T9BWMQQjB7wPxufIrFZUWnH7WIABYTYgW9bsuxbsjt8hWV
Dr4kX/FwRO9WHMdZOhG+Wze9uBbOhrC5g4ZQicCOJWM58ECF5D7DgB46MEJ6BLov
9KEGE2zRQUHifiu9iN3Kn9XAcJqjCPJlroqcqjR6G+aTyMk4/TFjeDcNTCWwacBe
rL+a6ndAvq9n3GD/eAo/BpkCDbkBfbax6FBe0gWDRYw0vdFLpCJ9DIx3HKb0ij3u
V2TyffNpjZnjUl9P65uFqJ1YIYiOP6fyZuPmH+BytqjDgL0bHfpQR6LtZMH8j5ww
yeDgd0AdNkz6RfP4kvE37PJEKlS6SqcXOlwkSKL89yTi3Ip5UEAiSroFRArU7Hc8
u2BAQl2LJF0MuzAjdatTIW/2Z5JituEhrJQXcFhIvAUwVQWEYAPYLC+MbA0T2Bxs
B/2rWZ96dFoGSkJppSwcnd9H1I0ji9RB2D/b8H2ItGmwbcQ7IXkFY3FF6/F3hzYd
9UbtdRQmuvUy9oeMvE0J4KNJ8aP0VRF9SVcIEiXgBko3TfrP8re4HEYbYwHXTddr
XnpszY2k/Tuhs7Z0SO4GYFVxqD+dbk0uguad6uNX5DTjO/5pVuwcj5JnVy3jJTLn
UDq2K4U46R5pjPCVsplmXlrpXXEZugWxgqt5UACV+y9Z59Jq0pDbZiVdoN7/Iq4/
J7eR9SkVoOO8j3aTc97pRoVKD31t7412ivtoBHcmLWpJ1pLkXhIR8YcMssKHHWOX
iVrEnSKpx/jTlyfRW2BaefO9DgAQ3rFmNr9eP6srzSx7hRIm0rxEgHW+JrO8wRZC
FqFCyALfJqw5fDhgDM9tyNbLvIZVNOnlGFhxJEWErXjVVJLtkMdQos+rtvUsyrbi
vHel2SReMyz35U8oQFdr5ZFQ221ybGw2A0J5NZ0mM+MU5VqFCuiGGgLNqyk18J0u
of6ntZc60CqJqKeqm23JCY5w17E+3eRYOr1k2G+L0AOdPfzYpcy9DyaDhpdJ3Bo4
ai9SpHPcuGxmCueon+DkdXtGNn44+sPMbEEM2i1rBQVrsCRsUIJ3AdFsAfDC1pwx
yEhSoUkb2Pv+HtbTlxkMh1R7SdjJ19QwkqAj20pueYJSGyrKMfPxAyxughemoamM
0QqSE0qZ/Jw2T4Me+ntCY1K00imv53tPi2LLu0VL6Tq1q2o8/QS9dYlSp6yeF0AE
awziOzkt+p9JaDysAfopkevhrh6e9sjFmqq8n4QORmCARl85tzr/l7sqXlrQpxIg
jcDf005NN6NvoegfBX21CJfLlm/YGLrd1yvQ/XWAjz0cZP8ocr1w5HcaQcBmRj31
hckLhsKwsDhD/W87KdoySRsFWMGg5Gqqr2+5QgCD9qUYzVEE/cUHLF04FswBxW1e
/n+3i/OhHan5Dc+/Vs9dyN/ynx1v2SCE4Eqfg0P9ICqzQjN9I56F+vqvGLCEgAoT
mea6uI5CKzSgQc7LijOaaAIfpPJI2ZDXjSY8fiUtEVf685hjljoARBHcZXnc+jXN
YsEZr3uhUwWQBgl0ftcQAMgfBJ2oftAtAFXp/LcLTspCCeYD6rmgLjlstnUpWcZc
GqyH+pRHk9ZLLq8j9aZvLOUJgy4VR304k7JZf/11sqivmJQrgtC9yjGseVjwJenj
/YuksHz1Ek0Jpp00YcLVVD2G0Ecb8Pmi0t3axCXeukEZy/tbS6yQCTlrvkAYDL1N
koz/y+rrtyCf5OAzxF0h3OJK9IZAFz5CqVaRkpLlyTMJiTadQ088P9MPpo2Ln9KP
TMOhb0I9y1t/E6Ij8bGwVZhM9L8QfptX2T4yR/jn9RW1Q7tt7V5+6p6508NQ3otv
SkJEtQ7AFzf4xwrxC4RM4PXN/OieZobYcNi07bSFrNT7qu5i9bmnJFGKCHm7joFD
nN4DA+SGcQL6uOphqxj/IN5fGz++YXdS2oYHh8jcfQMweqIUmjHHbX5hc9GNVd5+
+BilmmrgKWiigYPgAl7TBy+3ivNXSSzIzqhqXxaWaqO8NW2wLNZckbt8B8lrw5ON
UncL9WOpn9xsm0qHTPA63tBWapvWTbQFcgiEaaqxbOIUJSDzpRTqFn+AqKYmXPZD
NzoaVO6ToomZlXEGvtY1f/z/iYRniXhBiaXG/mm8HooZ+V12vjuayyfrSTP+lfKu
or6e0A+J/yG7Elmz9CUnZquCsNJl+My3SApXo/GihHGcZV2LzUVJYv0hqbDOeZF6
JxCxKR7cGty7qQ3pNkyeaqJroiq1eTVAYD9/0UOTTpn3fy5LKRrZfgcgL+AXU7mL
xFni1lrL8/MqzBv+tF/fYfAnRnk/GVrdnV2CwOXNvh0EaPOK+p+MQqH17bpe3SeC
u4qRpU33flPZ6ywuKvXsA5Y7G3+Ri4S/n4Y41cM7k9jzq+4M5dEvvzPPC50bUqvT
ug1tH5i3JpRiEgX6rxUbBhBUwkS6k/W5mEytPbY9okMt3k3Skl/qIPL1gMGvrz/5
GwwbsFCcXvTl6HZK2Vhtwkce9awzV0amxfmI8MzC2PhmqTTP2gLN87kIwLgeFkzi
ZUfG85zAtRl8aKvW1afMxXUINuYj/PD16sOsYRgxsEW5IdFb+F3MJWf9pZt1/0YA
IhBeb0NZO6fRbQcuaekvqZi7y9RZJQ0zIjGcN3/7+5mxOcULiuq/Yj7jHVNxL26y
0sWjTR+Scd2FMfTmiO4dpCA2qVtbpCnt5mNUn/cGl4Ivb3X1VVERx2xcg/j31QL8
6rVM4tN+nvwbNZk6vVwouPFXFw3/TWfdbC2JmUowbdv9pnAS7pp9r1IlB9NhFJji
RGIhaHQG1LX/LGmxg76JzH7WmCdLCdOlJS4JwiV0l5yakDKv7uN/ESJUmMQ9zaLL
Ji3tof81QaGpvQJMsC7Nc/gMtr6vAhNY/QhUSf6DKKiuJrPG8koGklfHDiejzMqr
PSbQXhdlLEMyyh/miuZQnqA2sKcIk4+QxhFjkESZRkXqw56SC1/s1N4aTTKhGqg8
AYCZtShAAPFHYFnWA8fYoeKRes51+B8El1EQI/hJvPiWb+T0Uguil+C0CBIDcr49
eFc3TufcmOqfczt8eWhO3+uTRNipUk5PFhidcDei5fCQJ/D1n18bY02YyZzrzN89
p+a7U4PT650mOMsdeE4rxFF5Q7rvYMXpMizkK+cDv461h9R7WHEYfubpb5iHyaTL
wRu+XvaIoiIDb3aMcwgkODr8zg5OzkzMYQXzmb22szkeSdQBUC6dnd/v9YWXDEk0
4N8IeBlaNshpocIz++jXIUfKtVAQQQyWJC+9yIB+IIl+n7FyqGqkC+i4tziTh7BU
TYaLRtsCbr0VB3f2s0iFXQKDgBRms/O5SFkov4QTD3t8+01oDG6Gsr9aIHnO+1T/
4K4eXVjrqmOyZzPZuTYrNS/Vixl4d0JH4+XYfUq4xDfNkrUcA7rgO8RtBnV0yE+9
58PVT2DiLJjsgsN3csK/Y3VuqsmLbVt3BO0f97y4L9ZvXxtCNASHQnAdn/dOzSTL
AYPUSLTbHDowjDqWkpP2pBkpMBMLgLyCmDt+P6EmBCY1zwfMEvZxvjsbSnI1ApJY
RXnJyuNZ9US89kgZZon02+IZHk1m6xVVz3egs3+D6fQDBSlihL4RJZAMkcbAiIuR
i9xTbhPaTnS/q/hqupzVpwdhI1/9LiBmgdV6UQPm1fV5QRNOGlV+p0NJU0DI67jA
FcI1g7DqUPI5SRpN1oj9nO5RirJ/G2mIiZ8wKNLlMzmSUU031I/Q3nR7aDPp09SP
dZCMs92ye1onv106lGRqlCDO9BSluML3n+m88f666/N9MA8hYkCdrItia5AVNOAZ
o33yHR4BJg4mktdfDN2rtIkOcnBoUcGasP5doswotxJCedtpKbZm7qjF1nJKlcCG
+l94lUgUiHure/vp2Zf39luicpPXYTfdCXkr5eKOzNLF06TZFP673BgUwM1M2574
WRgcPxwUO4b95/+76YapYuRglD3HRjYXIPdmal9WKNTb7qWFLODCPvt3Zpby5spt
IwJNEX16fSc6hF8iPnM4845uteJz4kUykkGqcXwl9NNjRxRzFxGPt0yVYvEFeaO0
V3iweMz43Wr06u8V0N0D+wRU7DcsL66yfTJLDZY2f0ugQwxqC7xJFNndr/2SbHRa
Hpqjwcs5vk2GhZx8gcqZBaTye7nh0yh+oo/3dyMHark+61P0fxGA4tNTmMTp5Q+m
h6gLHaMmVtRprztTGkpvzxnuTgPrUCaVv36frl2uJVSp9uZcWM0jjCAKnFK8aZjX
+s1bdGgTezuz59sMQCNsY0K6kd0fKeAm6CxpKRrejWC5XJ9B6bH8wrL4WC+UnNoI
0zWURle7jWamgZeFfZ5KmL/XhAom6/oiGCDJyQ4lDylVOd5Zuwe6bSroy3R1f81E
z2p8fLgcGEHvKSg2bTDbe+QoyYd2DGakwzznfl4ijekuMb9gpv4KLl414sAeGnpK
OoP2gquULLWbHX6Rwdsp/coBPeHJo3OFtDUbUv8YcllVKl6rnD5xP0fGAwZJB4Ip
pNgCLRiSB6ZX4h1QvyvSrSvQlRv1rdcIVe3SnawxsiFFNgFUn/LWmFgi2E36lv8H
bw/vUeuuw/0xNpcPSZjrM8CQll9ug9032Ost/6IqNENLcXiKTdfevUxirQSZF+zw
43MNsN0kfifp7nua2oHg4bozDBVdDrdg7yU83bB1hTDmigW7lWStS1xtT39spxv6
6UArukLwFcrhlCiX8+rELDwHkmwchH+Tc6E4wXVfM2dH/kSdFBDCPklj5oMkyJ4w
ySVGVe1rdjApnDhG7kQCidiQJCe1I0S5zTVcUHOLrHPQcu+SJKtwVPjP3+X6KjXI
grnAZubKlggpLItioimoKTa9xSWq+aO+QcQn4iMk5XSrN7MqDYF2zW7eu6JvcAJl
CjWCqlxrnRhpScBSnPppyBUFII2msLcy0f73o+HZEXOREgvSZjWLYbhdAOXDHvVq
I6NQ7Kl7N8oOgr79SD4GkdPDZJpAthAFJYxKMTA/dbyJjQqz5byryG3Q20PvaQcK
uDYpKBy+bRSiykhIX5TQFlka5g2iiyqHl8YmHd//E581zvwCnJaGqntwzIVzJy92
HLwPmkVJK66XH8y0shsmCvJhPbllNDmbYjJxcWWH2gyKsEmpgTlvtx6W70tJjkC7
8yltjFGXVpjI7jOWRRZemorkjT3KBVFzNg0gg3s3Sv3slR/X9TYfZ41X6f/pIO2B
LGo/n1sE1efTleNI7dv9hfhU+hgYVjRAHGq86153RjFqYC+Ta/W3SIY+Cl8TjdSl
9gAInc1Rktas8A6C/IVgyFKhWNSiZrmOuCIRDqZVC5O2nSzHAyc4jNid/kMFMUd8
Ldv2CZ2R2Rbh/3d8l1hjWHY2xWAR+oyDWRok+G97WPBMLQCNGaB5eK3W7W5dE+3+
Js1dGoPXlc5XiJTyqwn6PEH8cSTf6lMp7BX6PfvS4Z66JIBFKvRHeLh6nICrWQqc
9MXlGRAh4nrqq9tYckTpPuIDFSVIaMhV3IWqUnNpzg3nIQNIwGDdfccoX8pBuNQb
aAbLkFXG0CRB8bg1+a1jKlGQR0WYwSJRKupwasawBnc/UxhMbk0Hd5yYoktbZXYf
6rpc8nQ4QMlTWeTdvkgofY1hp++LfKzIRD/gxgPudxl8NwAIkmWw0+NLC1JzCdft
EeiJe92PpyzdItytii8BsGGBgY4qkdt/pKJ9XAd2wFRqjaT6WDQ5ch+cTbLD//+s
UvCgbqyOWolPoj+TBVYIRGN7cdcnoFrPOkohCZYeMuHAKVdK9Jt+21/dWV1K1056
7PDJ4cargCLrcoIkqqrhbDPOmcYeMTQWtUa24olCAQVfIwsh/VWSwWBxIn1DtaZt
2KWY8G+D2wxOHSitSigrRjR19y4WpILmGBLNS+2+zkrUfv/2uat+RLTgzzWMSBrW
JaleDGOBTVUThVYV3A2fOMg08GHqGjQcCJ8e7beFhTEUuCBIzVffYBeEQcyXnbhy
FKyncKQa3Vo48FqCNvHRKurGwDMn3Y2aj5P7iu46i80cW/Za9CmoUprmpEoOfaUf
KSY2Kc5hhO4OnQcJocdtAHQC0ftrXtwfHYrcw5Yq27zUACoMNKBOZ7aElNAxA6rH
hkAXB1jqKVq/i2YHFktKLSeZCDsJjCxz7rDQ9FsH6NT4GDAAdXjHVLb19YT6kATB
rL4Y0RZKv4E3xO7pS6Bi5kNZd+xOfSC4QIqauUYl5t0FIrGbO2lZODaFKa06rez1
1dCLHaBJFFDm/b2bXqLYxpEBoe8HkQTbwPfNbH0dNqzQtVFctowhLtb8cEchMfzQ
Mb5f32FHSy+wbeEykPC2YFYz6oMgTIRoR2NUEpnGNRd4pvEwbyIMqOUC0V6ef381
WsIejwDEoSykJsazsMp51W33tKtIep4L7YptZE2dZMLLm6aOaV2NgKoGwGfqIO61
Cz9PDrGb1GEtEDBNCrVBVOJwMiM6QmGoPpjlUpzsPhAkck2J6Z1bnoKdu2Kp/hB1
Q1edQv//qEeICweJqKsCHLde6XId9R1q2XsGyO11TxhR0EybV7w+pjDSjuVbalqt
7dZYJC3Lz+Dt2+W/LLH9BsKKu5XYGUhEIdTsBVs1cAKhOrSdHI4L/TX0q9lbEx5y
fH7VMb2EYSbEHuLfTQxv3F7rcfqy72SOYE2J4a7Q7J4AfufyVhtkUjw4rpVqpC5d
hzQgaWAunOYiKwk4M9H8WlsER5rhYkzppRE1Ix64GO3KcL9owl2vSaVuefJG0WEr
XkK9a+OYTub5Bz8S4JbLHFiDJV87W9VORewDG8AnVR2UMnU+0Dasw6hHRHpclfzt
3gSh6T0HRKR9D7vQOW1tQBdDA5yfJo76UY/yJcDFatyVzPB0/z7Kqmt+PB5YhFPe
DVgCg/38N3j/UOTJ1Qw43MrRqiBsr57DOvVFqEfillvOymqHIhc/fOVk0BJbOmCb
V5nM2yJDzjpMxllkEfkN+5Vkut368wGzG9vLhaVt15ZGQALpAFkd8UVqaYX6LeuY
qg3+FhteJBcoANS+NyiiA0701m9RuWnI+aAAU5vYWji1PtNO53gkg924imGTPMWK
2VhCmziVouI0epTgq3OjUCYsRfRlSRwELotmqcaVWiOmzfjR875mqzZ+/6yxGlZ4
LRhSjjLcEQInQBgml7pjMjbAjGqd6iYGWU6qCcuBg69ETsZFApyCsPBlApbvT9/O
LvoGEBTzi9/pk9QB0i2kf6YX6MBhwDExdZTPzgKv4zAlJRZp4bUg2NUnecdM/u2u
cvTEO+srhUjkwRXQKUfR3dugY1S9P7RV5mc8lMd8BFZA7uLxu3lmsDIW6YurbtQX
CQ9J5ldmdiIYjhdOKKnN+R2PwMR2TMQAIR4qX6p27iyc5Ayeg5WLxEC8sNHn1g0R
NauzhAziSM27/ucuYwu5pnZujtpvMbDZszj70xsHswKfZv6PALbfjUpPOVH8IDSO
1m1NePCvVgNETZQbI3sEzIF3NGj+r6JNieWRMa7KdDPHLNZrga7kLh8Y+MDYPtUM
xSctbhBfJcdFCkkccoLQE6IL6nbQhd9w5THmsTLztaeG8sU+N522NzyzVDVMyiBo
Ex4P2m+5LhsK5ZZpxHBM0B6mYy8glJEJiO5OF9xrsvKJjEM+7OXbnZBeAcbJuJFd
l66gGgnkiOgbEg916LbAeMoPiihY8P8ss1s2vKqNAr9+8I8lfV71ITe1lldYkJDz
KbnWViFRjPtX3be9pex/vrFG/4x7+rl0hSEUKmGh9veh47jsfVzdJSu//A9TuSg/
PxbjtcRtOEAxO61QEdXx3noV8n6mMvdFb/JKsqz9m46GE5mGaLw91MVLmmq8/h8u
d1QUoB7wPDKxonugR5tg8J7s2mHwpUwGKuAQXi/9Qk0e1JMRhjoIEMO5hvQhh5kF
Z3/2NU9Axj5W2fDcM1pWdnXTrom9ef9Nq7f+vq7SwHYp/865SGUbikmJ80UYZRXT
ZYxGC1UCAx2QJ9Sz0UZCvCo9N1dEj3Oc2ygRBH8RpXenprlIOLwOVCLC8QTSLQXk
FwbEWW75f8L88N+GXH9Au94ScnEqFpV9JmMI/ylCDW0bXBZ5YgfqUGzm63YJzMAV
CX4SGFmdAr3bsF7wSjklQ2BRvQTVL5N8n1+GZUl78vxPBZNIqopW9GWO3pOoimnI
oedhTnR65VwrsNMi9F3gafmjF1L5ByQZjosAacN4Li3fMycGO4MG5x98rFNX1sop
RpCoOsDDDIsNALmp2OFhbJ4xNjHY9/MNmjjPzEn19rCwncItV+jKbfkSrbGKV6gB
Gu2vOzpRbPQB2RlX0cRMgXj2DE+XpEhANYHQBNURwiW01oz94XVLs+1GnnPbQvo8
CNAKCQEccAsLh6FzM4uGcbCuBJY6UBIv6cutIgSAJ3i4fn3Sr5xzt7uRuPAtMQUO
K+7eH4Mznk5/szgRTegxucYic4gnx8IqzNgtz8eSxAHV/LEBAbzWi4iKu8COUhX8
pl3O40BQbet9A8N6+KMSD03+l+s200OhGMW5NQYWPxZmLyGZmIv5/WXYlLL7Kj8b
JHqmhTkHDqfkMisSsbQrTw6CAWFcxpBXI9JXPHJRaoGwOENTrT566GkYi/3HZ/yL
C1hbcqYs1pGLXcKyF59/+h57Lfsx4MygTFJt39Txj+OpvH4QDq+tGav9uupJAdgl
2qSQ9GOhOqbkFIyoTa6Xu7hsmcIpsH1SUIfTCdJEz+R/P6F9zYw56+ju5bRQsiVy
/tMHm1TLq7TERCpUA2ci4mxD9hZNEo3KxvR/99QtORSWXQAaxQjfOzV/niWGp0CQ
zi7axjwCPo1N5lMYS3NTRIuTIPQHi/OsBd+4ZbJybRAZ9fgJcr7ZAG9L1JjUbwx2
gwhWvgVgWzNWflsr/7XgICsFSSmo85tbqqshf7JSS9swZLeNlTIU8UArdGCk40ny
Y9WMU0NdYHkuvBq/NqqvIjGB96WTuic13Rb4z8ADOpuX9wmqdBSi/0WVFTtlbwDo
GJurfSKn35HdEN8fbXg82VqOPgi2VIGNLRoDTU+ASxGWvmnimoTQCes3zeJjT9fy
OfZyV+WQEhhsyTgPVy5ixQgpQQDxkVrQt2TnC1MkB05utc9ia/rJNNiVmggPhrQ7
p68/M6ahnLKRr/8kEN15OmpeVThvaMwjPTSjxxjxDJmHvVO2QqRSCv/DCc9ZjUxg
xcOviFFbcPBgIkarTYxqFy1GEbJpfOYHgsRC/4/e+aspNDDRwT9RPw7ig9NBcyEN
/kN+nfRKzDyi7tllCaiPmTjEVRgnQ3pshz/lHwEjxb27KZQsTNqu6Aadmkv1MppZ
xywJxaKdQUaFVxjW6dsTJD2IvUvSawV5aE1c1kyce/W+O/A2bf5Y/Tsco+7uleIb
bWcCfaQ89KO2kz/fHQzwqQtd+cFx8GTXOTdWfSknNf5IjkUZaWtGvziq6hySDUa3
hhU62HEBz6Sb5kbskhN3Jj1FbAYnmfn7vObE2NYdEjEgyc8/ewa2Vo1HCJpZrwYp
YmVxWCq9z4PAR74Jy37xWzll6yK4k3ObcbF5Od3sBGUmKBKS35LgukD0BqOPrRZp
b6LYrHL0QYDOpk97Y9cecK8LlfL5hRMcIijBTQz83YPY5juyW1H90JP8OWdh6N0O
GZLNn2hKjKTl2MJ5TtXgUIOwO0Xk2zsGhLwilqZHITRYgFjgFW8zo5OgTEfXSLs9
dy3aZHVzYZuLY/lxoZkW/u7qBLTNTu+3U33mSVsnffk+6iKGdMctHpdVommpBrYf
v3yBZqIjiTuY612lgfrjaBNl0f7FoV4BVQMEkTaDlnxjR5QkLMNqHX3hNzAXn9Ji
zRRrPhENYIe2+EUgj3XjwWmEigf081IEjdGFQHL9NadQUwOnc7lIiFUYakY60Yc1
MK5mjNfJNeF/VhaIcPBLcgBU8t9qWhWx+KI2YHJdatReHbs4a3u/6lr1uk11oaFh
psJwOqluZJXY1bQg+pqvrDz/EfS2gBeN5mLFDxOgCWzgl4PSn71MqYKdAGD0ZGQU
+GGRKWx/7F4VRxXcCcwazFAxMcNBEkg/1tJzQNazMJ1FoR2J8ofphRfYIbnSCEb4
jM3/wNLKnHQa6i4epPz3lsquc8kOz8dG5oXRT/e9qUV5dPIiEEvznhWFV270iWBW
+kHgG6Yd8zGcYfQqBiLyj8BdG3vBAvr2ra5b8CJIdKyMVFBuFZW0M4/eblD2VYnC
tsLqckchjalVTeA7v9o0KAH8H8zpNcndu7o3u5I9Q9410y5+G8N+iUamhU9Wq2FD
jbTe7eTOAzlXeRTVu+Clflh2vuJRXkVKXjl8jbYLyszilxo9zPUzqadEyeWdAQ6n
SvllNjh+Ng1ETClwCNlZW68bFOUcZsVd/EZo3BczLm+vTZdKohJCpNSjKhpYN/k3
SuyqDJOlqQOxX0zMs0OVv3RGNSZtwGjQP7md6tbFfJUmwv4H8rP8NujH2+jmuqP1
sUHF1FAInmvqSyin+clU/8OBgLgK3jp5hdT8IgsAY/65Q9iL6dQrcw/ddn+CBh30
B3yHcQzZiGOVe6EVKesdI1pPKUHknPmZuw7egNQ2vLxorzrttZSgtheX58uF7esv
cnjwbuyVHjGEixBn/RkBy1UXyf4WoVM2TNTje/C5uPy3qos2cleBwPO9mslV3kp3
aGgQRyap8RT7oGt8Sa4O9GeCNTyZhDdN82BWVE3U4mwygc275/B1jJp2CJwhDB02
k808N5qvXR5rhi/jj2cSca1A0M2GXrIY57AJvsrHvIqU2IbAHoDw2lyYPa0Txsbn
nenCM4FaFUtdzEd7MteiLeH3LcjCAuJAZk6Iu3lOOvDau/3ooqq0K8vlSmmtyoc6
dANNm3F8kBsudMcWbcLFwr/kusnwo7OWIPILY5aAe1UcbVijym8R9IZjpJa7XHo1
fw5XriNfFZOvUQU2WnmVjlauY/2fTQFMgsRUxf/0MZI4HwOAyJSxsTAs64DxIcNf
X3j3RMWFIgTMVQwfNsN7Hfpw261J6nSN/NDdDwTzDMaKezkxyGyPRZ0Pa0DlgvSE
odcPzrLINOaecVy1s4zADGexi+pwfqZ7HCsJTGcALU0T8PaDv0xGAOhRRhxzyUln
AcAHBIywn9vlv9j/e7EGpDjtlaCJebc0QtOklnuOByOL5yPhmNTw+P9f8mCWYQek
kIjnQehJXOfD+36//FG3voaCa9+R+f3qK6dVf3P46OVm62PKo7UmSm9H3juM0YyV
61qy0zhdcH8wQdhfoO+MtNXceKe/QGWidNKEWxdfxgKz6njfKckiF5Yphfo/zj2L
MpeXHlYSnrBSEFCcs1ke8LMZ8SZF98uCdFC4ZX1Gejoz+DMEypZwacd0em/UN1eR
VD1erPDIMSVE9R9kyH+rdwiP1MPQkvmxumzN43/g859bFS5dBwbZh0q2ng+U7XKQ
OvmeA+gV2V1po/o+fvQ7/lVF5An/DWRtenmiYJUC/pmsX2lJ+/qf9GIpr0mna3W7
5TdtfUfaxOIHnY6FuekGfvwcZR6vIvKwu1lUdKPm7MIkZdo5vVCjciVu1THdABkf
dc66svM28d7XG7yTxKPXPiDquqWIRt8z3bmD0r6N6LxvOz4wXbY0LR9ouLGl2Yzo
MUTs74V9tZmRQUoDmAcDM3bvUCpwo8xjxlR2IJUTdW93mQj4Jl69KZbKhAbfYSWJ
IduKLqNw/8qT+8ZnL/62DtTPjlddntGsAJvlNZShU3Zh7qAqYRSqzKA7K+XvN0gv
v3S/iVrEeVunzLyT3tWjcKKSy7TNoKTZftAlpf4OXL4wGsYhHEWPlWSyt9mvrpLJ
KCwB90Z2Axd2k0/2QQFI5qYhwIuC+IJxfj23jkADQJce51ZqpgsFProrx+xY9G9X
AAlKHKHVKoiXbZUURCBvfW9Exy+tUgATW3k7LAvb+bgMRSserd1Mt1z7zruLF9Dt
wYFypNhx8z78otD3n+rD7kTfyGnnG2do26NI35uUh8dC+DAVkn7jGW9mdpr6+1fe
/wQGaNzp7NBPqr3J8OAk9nV4jvKUkZmoSw3uINYUoMk=
`protect END_PROTECTED
