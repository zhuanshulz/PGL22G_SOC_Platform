`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0kWVG9jkWbKgBWl6zOjnUSsZJNJTyRgGC+EwUWxKQhmU+bcOc4Bmpdl/wUX5olHd
ChuB6fw1A+qWTWFWoUcDswjeOQgb7n5P2PSu0mLqPZ9JM+yRVQMhGjN5uZ6Afd60
3Y842U1Tm3Ujvd1rJ/o0XpA09PGjmZ6w2xwT0NUzYLRXUu4v8LYn0/foxW82pEDT
BSCdAOPxJ+gGdXtecybuC/CdOBy+mY7IY7tPK1F1p2anUbdFir2z3Dq2KuFDvucO
0aOgTmOHRRKzG/Ht7NDbHRLke8sBOaVjNI2p6RNY7dL6ws3CumKu4Nq6fXlz+TR3
jjATW7zmCFGaSZjtyje/XD230G6+2vE/6qDW3xH3sTuKBYc+2Chq5zHK01SxvlR2
72cVMq890l4yo8E1rTBbX9T9ZE5rZphoMOfzO9+6GbUWVvUzlnL2fJQ+PMGmmYV7
S37MFxrM9xd590yorH7JWohC+Dzt7RDkM09cFwOAtAOSMfGZrda0WmFZW1v6am/W
SZoUOjWq4jdr999AHCzLHFIbr9hT6qFP8sfOfwlkDo6gdvyPJDP9ujouYjvBolPh
0OfxfgNRX/nqDJGxbuB/dNOpbd2CM9I4Nkrm3zJE/nL4NS2Sa5IPn9bnwqNMC43f
78mJx0uvhk+0ANAfxF4KxLxcKY0+g+Ks6RSn69Hz/E0cReSw/H/s6y7gjC4W+X4u
E4xI6iVm+IsooTtKlXUUQ6D6kBV2z6X0kelylsRAbWwMdeqxQkHA5jTSe2kuaMot
SPTRA3WeHc8W6HmE93lyQl6C+SeF4k70KIDGGozUCgDmaYR8+yxSPs8KVLyZzWaC
9ee7cRWJ5LBH2LfeB3vep6OAIXrzA2eQseEOVc0QhuwPftZWUJZ75cYKkPNom7A6
s7Xx88WSmkaKoqeSV42Y/1kcLXRpsek0E/IWKy055pd/jWj2a7/kXKwoCUpgFkni
FwfgpUaESD5YINsYjeeWtquCtKU7Zh10YHdIPoNukJ/fs2bsRUR7u8lFspCErzu5
RFFd0FpM8u2M8D6BxXG4cTFr/GAnoZt3sP708TxydQMg8Oa1NNPrC4ZeZd1Ur6Wa
d8ZuJHOtQFaRaLeSJaFIvkqTEiSNjhajAAY1up/VaM8ynECQ7WQh/XsDM/Vz22Cs
XcQIt3JWCSjS7ePTpwiqABz0Vsql9ZxsJ413ue936i3hnUvcKHSAjtRseoGUaQgS
sD+RnL9jk5eSq8hxOHilMtqz+mLSeUeuzYCkGTEvTgQ39wYYDPAK5aB/Ua4zU8DS
jXHvQjXqhcCYmEsPvPuNhJF0w5sPgPlKhldqyorkR0hsKSFV5L+AY7zlHzJXshLz
UNvIM5PZcQqQwfhUdYQEPJfcYr3d69bVMBTE9gwgf4wtYWPm24eaGiCEA8YffwYa
FTH+VxVkdxvsfqh7k5vIhuOFbJQY7xjx3Jpdsoc9bVVRZ3xstrBX2MTqZ4Y5O+pK
oANKxhTWEO/B3dk+LMCwYHUFB1/BiL/kgjI8jMs2B1prt4QSYhlQHthvR3P++uXo
To1f1FkvUjS3FVmWRzcntD+awHrCfYIxjsnczW9fTDpCo2GGE73dIhxwQOWMPVId
/ZPhWxhC0aeQ106H66MuFHtQyncoMq8DZYdfzZuszlvWRWDm7XCZKQEdi2+2Hi7j
VKlO1DqXWtXAK92Ly7uiQH7qjN+X/JOQMQAkasKNDe178EXGE4M252/gd8NYiVjz
uyisGSiJ5IaDooH8HM5HvehYvzwjU86F6sJn/5VasXv1oW4um2VPDK04ON47s7Fq
z8LuXjXSDrKt2GpCgbxQGbT3qghzUaGdICABH3e/QbOwTBfMwvWiKD3oUxEw7eJv
8BwBhbX//0kFDBcYuPjG16oZ1ENe5bsnxCq6vzauOWaefc08IgLTylZ2y9tLQmkD
YshSEGCqvNbN29eAvm0nEtEwZ1lE+D16JL0RyjkxdnHWyJXqCM6D57qG1btibVy2
UQBG6JYhstr/H/fqWHgBE2Ro0cex67o6hKwVNUNrgqDpbv6fZzKhuajHjoCM1CxU
6z53wufqsDE4sKRlTI33alyWbnkQTH40V9hN46XRwYMyUtYNDBpkaOmJp4WzuJKd
mLB45oXFsCxv0Bh+qOvfzF8Q5YCQ+aILdBNbNPkm4oz06FaG7Rw9ABEfY+pjssUp
hS12GlDPR2qUlO6G+6N14j/85GPp0MZfr7nb0H1J9WeYwtr8v15p+HYeHHPr4zGk
DO1ZbTd7g7yvoQqm5WC7VyhOfZ3GuscyTVHSwqCigd0iIvWfn8HO0XTO7T5sAJ4E
XkqiA5JxIpuJzyo83wOWlXyM+rwpcDJhXGLqvA+d2JTNJ12LvzRozugNgAbW1d+H
mHYf9NS89rShBp/LYBZgQTAf7Nx0QQGK3simYvPSu2Ss8t/zFC04UCg3ZAV7bMjl
/XC7rwgQ11KwTdymCD7K2XmjJloJZj6CECrlnqvzZI0gCoMg/+c5bz41c/PimeOx
EXmNSSWDULjRHJBCoDFGQz7NypbyE/CEH0pBZlya90Cv0Xgqu+XN5VVoUiED3NBi
DpFOtaOcg4Bev365AkdpB9JavWDCTynd/lCMJFXAnvh//r1Pt5V730FCNzEHyN9s
Nj30BBbIy9cZ79OnaqDoKQQ5HVmmgQMCYPtaW+IqLbOwi7hhcuq8PKj3b424J6pe
1Nozj0o8mnYm9IIGiUccjIkfBs7CwkXonFTEc1dBeMW9iYeX9F1Q7MMuZFixux7I
j+pTE/DGMZkUKhYQyEYryl+8neaTs1Y30/4nA5+VDJP8+Q6ofgxBvsdlPZPLDQuf
m4YFYj92cD5yPYXM8Vw0hBzSj9uuoNqPzIizWRo6yMHeK0Pj58+w1SqUmADWSife
22yVFOtMel1txmotKNtNczTKLyA3gGy4uf4E9aIu3D3B6xTKxYDu9hcbGschtPqc
ua415Yop2ox2y1GFscdEaH61JIOQmcFl+3TNmomqgtCduqCKALCS3JueYDSkGDfT
dhrQI0nSSBLFX+q/JMr4iH++hkiZBGupYs6oAAcZmzuKN5QWOc2YXe/VTrgvglT0
W3jR2vbu0R8u/g8/u5r8jbwhf79cNFF75FBnbJSpr3vg4yEZsMU8ywekx5gFmiEB
c1eTnPHUnIznLiGhiFXnCKod856j/ftZaHqoccZKF3clC8lRBr4UNB2oBBPQ5Ck5
R8bgELqG7PSOg5Id9uNKNrn/K5S34E+JbDcrLnd6+9jIzSOcnJThfqN0V69M/EaP
Gt//C+s3kJPY2e+ptHWVVZLdYIawLD1TNZaZ/vJUOhrNDqrP17NBgk8JDld2/5ev
BJ89qwKencZ2757lrnWq1xVKjpY2xY8cqHkuhJh1ZwolmxyyL+KaRq5pr1AiS6tJ
w+VpVd6vuQ/ECMfwk6xJ8bvBqp+ct7/SBee8zWYmQzYoMg+oHBkJcNz7czGKwnRJ
WZ6GHFWDfjVe/cLLggPra8SWlcw2HXiCmpYXflPnLpt5oLLKEbTg27UZ7CQzJGQb
hZHYiXiF89Zy//m9IGEwjBaWdXGOhridbhD4Lr1Ev6scqKDg5VhNVrwz6AkGIuJ5
hvEjZEFf1NEMTBQtLKVtbkHVSRVQukHJe6H4YRILM4YLWlgs9Eoxp565si7K1q24
hxDtyt5XJV4inbZw6qmHou3qNORVXH+dx/WQMGjObZE0ZxQhohU/gqBDmlzdH/Lq
Zj5UOa2qjulEkJE1nkOvZUOtS2fcMNVTbo5VFEBDiU9OK8lQSRPo6fueHS8W7OZo
Jst1Ele9IYnhpJQKtkxxroZr0xoA9cpKy68MO9qbTQdJwUaPAmtl3asNKHCfX9D3
Q80ei2jgUZkLI6qLCAWLy17PTS7cX1LOY+x2ELoo8ByDGCIgSHQNXjTGpfd8EVSg
uoDWWfnrxvbouIzXU0585yS0Sib9mK/ZCIwZlRlIZ9HlcEx5qzyKayl9M2qw5/2W
WlW/F3DPNKBtawNzMbsnTh0dCyaCJuJJHOLLyAk61WYfCNHbESSPTtGgjS/FNIm4
/xFNR0IyMu21s/f47FD2EnU27cLc7yomfivrkc/HTIEWvktm0mr3rpjNDwPQCbYG
7RmacwJdGBMqdVs9NSi0gKFuh2VabDxjgLlEAsh4qBe+TCFCCpbeAHF9e7decDjK
7I/pJUVXONs8oOfQMhdI2vQRnlpyigfsloPW+9G4xob+3Zs8gW0iJjwKDuzXXm2O
+IVwaQ3YC8NPComz57cD9R1+7X7gRSJbA5J5fAXbLnmdk6wKALOFSr8CN7W+nwZN
Pmale5VhJWd1QD4tRilxZLYrzSMVTDs7XhYFz3Y7ov1XnBdX/sr3djnVFawXGY01
8QXX7l6l7+GoT6/gUJA+jS0MiVNqLKeLRPUDn8Uyq0N9RgoYei/hngV/Rzu23/Bv
77QpsE+RmuDaFArcP3sQsFeVZrz8CIZI/yxfXgOFwXciQxviIBTuZIBuGPfGTMSq
VM1Cwp5XHvoNWgqwwWQKVQvkEMUOamHmofduKS3Ctg+rbgLrN7ZjmH+uz8PX8DqF
MgT1ugxX5a0vuKc33Nk9XBEwDVXdZDo4gOw/umhpGFTrM5fUBzZVv2DnJz3IW9w2
T/Zdbt51j1IO3AArF59+YwRq3E4qyV8W6eeZRVHpdaQEbdafkIa/QWfaOPNuhaAx
SOQPomMgqK/LUSYZeWDy/ZYSlEcZjbMrD+HeR5WhKOuS+GBMyxqBRX6Mh1j9k6LL
p93WjEH8eS0Nk+w3FcuvnAVHOfxkE9acyp3zf3MxIlzkw9X0s18Emo5jVOX4rmAn
nnI9o7rjyEk0mCvZLjnAK2qSw8CTOCJjp339cb1x4lWEUQxOeCDX9J6N6k7iE7yu
6oWbrFj2NtnsxnhBoRDmVBqWRO+VgOMMWG+pL3iwW6yS5wqih+W5xTU126pLu9jq
dRQxDwrHsmQ7hS/+eV1u/v6SO0qxelRPReR1nyBM5tb1cQElpcQNTGMQxUvkTGmt
SXzacjZH9e07hn3oNPMwXBbePsHtkD83jquyT/f6S/+zhBeMJcQ6tEWRF20WYQHm
5PqOCI0zIBYwbu9QXA62mKWQztPFRrL03ug27TN9TpPYVqgWcCeqLFrBH8UEbJP1
hGltQDssP22Z1GJbDxkCptwnZ3f+NToZqSHlQWnp/y3UCPXffI4cqp2DGt3boL6U
8NzvghexkFFU9vEJXTJjCFZryj2PzZV1ALyxA6Uiyg8LtGc/q3HPm6kQELEhebsX
UA4sAFr43V5j0F+59T3YFjpeIvL8oeJJBGOkzNCoXInDiII3LQtyz+QmQ3kST88u
KXPTSwgpHDWEDZ9PEDQ5q1/NSMmDnZWvNOE9l2dgFQUsOKMYD6VAPIEnTEMHZL9H
8y2/m7zfXxUPSLh0PgWhsmReADxGD3MctKAn3WqzhMv5tsAIVonxu195Q9KcJLZh
HnjyXpKXi3UFoovWxzWaGma/wuoGvJuMN7zRON2VDFTTFgmRRwHSqu9WjlikCFOj
Smz7fM+cUPnvRo3cafK9KtLn7dB+9IRdmb5VPoYf/gLhlz/mIkYpoi7HRX+MA/Ty
7pNywuPc2rf+YDlN/iHNrS7On9tJUS0m3b6e+qgBeG3w2JT4pLXZeypkVN+xxI3b
GbKv838uk+G9FXRJwT8kuG+SMUuTXYM+rZ4MSGpfG/HpLtdCkYZnII2Nhxl/Cy1m
DztMXZafIyeyaY9/rD9Wr0SamFea7bw6sYRFJ1t2heuQMcOk0beS0id9UGKElIZj
ES/OMK4Qyx+ix7QhONaI1JDuCrbVWfi5B4r3l8fRcxo5az84aG7lS0dEm94uU7Jd
ACngcrr4dwFZViR1DiINnuHSH+CIx/im4AHgEjtxTCS7YFAPuESgR/VGxqn1v8V6
PeH8J1ThZU5pYB9PYOQs0lQLWSfn07YkruVHhp8Qk2lfgJOGSV+ZUlj7/SdWTyQC
llfOnnaW1jakctRak20lkGQ1QLRJQ7xCvYw15qt5gYGvYEXrEy+w+6RjAL0S5/sM
YclrRL1miNQ0N8+KrmBL2iyvNRQnOHRDfs06WHnOV1pqVjlIxjxeNVj27SjcjJrO
2rfffoIaJ8gdp1cuxjo2pni52a75mbb6o9Ouoqlg65T6PzawmO2NIWFyiDvk0BI7
q8OaFjgX0LNNdKzUlXdRhSfAuCbJQ5QSmPARarZpFGNTLOqrBM4NkNp8Ffg1EO6C
k/6we+XaKN8Z05S0J8BDvjhUXZef5UaollhXjxnSCICQIqHLCJVbA0vvHZBUU6B3
1mLZUWORhoFzeQR3vPnT8Li6EiZzBwtNMhaQbRTwryTbHx6BykWWtQfqP9IQIjgG
UjzARtx5HqIgAQbfQgtUirkVQkKgZDsf7vbqNVo1wNPuwX8htXgJpZMeaYL2A2+Y
MWuS2Slz+jH4HzlQRrzs0Rihs6AXsOkxFDZ/+NEWp9feRfsx5UOQXdGE6mxpCl5N
k6RjzAQYDw9quQAlvMWjnFw1CYEkCMy3c9kNBtywSDh5jtZ6Yux6tc5eAyEOeXyU
aR8XYiiQdoiAZbCUeyjiNVXPVkarNwSEAr2Syxm25F6BUqw9xNRTJbvyTYf26DSD
E5AkOdwZxzA5qqupXNmqvGuItQD0MpT9Or93GrQFIDDbkjZLQBc5iJ+hSZMUmRoF
7I5B7KaVv9iF1dlcNeAuiCNWROoWEFE0GU+AsRrDuLmRmuFGVMAYX9Hy6nBy5XQq
rgPog30sJWa8/dSY7U5aWg22qB7t7vcr75n6+ZvMxDClVdydzYfevdKnLQqobxY6
VEEx1jsKmqxyfbvA1QT7VW/LO+SFD0p6VxhRqGC1IvkWQRtKK8Ibs6V7X37Dions
hNMHtYpUWytLK++0pQcYN/TI0Kpi5YFHkzRZDM2osMm/1G88ActLoiTkdEhoqbyi
rWBb/Bid4dIUJK0P2ilJicY95u4i37zqQBEp9rk7xibmiX+SE5W6m6lwkFCcJpTW
AiUNdS9ug6yUxkIxLwV+hWNXEzhbdD9FkIUJDcgp0CZwRO9Swyt+XuyP3/LzAx1L
S69mQlK37T2aDVKIQAipwfeNyfLxJyMdEbEGEImXzz1KkEU/koWVj87P3/VzyNEy
NLjkigOwBFqyfXCB4HiXp1ou8CTXlWXiubSk81PmmCIuMH06OMF5QaU22tUbUlP1
GYZI8MOaHOwjNQImbyNuZl92W6c23pqDLIjjSCSsX+/V4kc3wyBeFmn5h8xIB4+c
5Yv0L1UwZEeGxOOWFaqvXYb1kcVCf/AKXUP4Je5ayDjjtdbxerOLseebMkHP4xT2
IcR1CBAXkYN1hViQQExE9yo8V/5tvIHWkB0t5KjLeQsREH7ONkbgCpFVyadML9HY
KHF30qKe4um8WLNIg4UhHdfVH074KgGS06SBwMmCIgHO0Her8RW3mtDLOOSLkTY5
3RzYpKDyYCDFIJShv/aj5Ccz0oNVvMYnGRo9TbfJDpG74ajRAoaSNrmtBkprwl4D
1H60/UuWStzbpwLaoSUs06Gp6/kWNibSQz2KbRKcI9HN6+Ot+x12Nvm+OVJuwoEA
MC0fuWvpXz6yuIPn9krkP7gE2hal/vmxn8vDyJugsNy0rHJQaUxTFD6JmyJCPYOP
hO2uKQNUrw40Q21Bs8NxEaoMTRg8S9Q/UfI6BIEp+Tar+N5qro/3yElCCRd4PS+M
EVdStzDhQpSSB2GLO7BYMeiA4ERStzv3QU47/uV/fF9WMZi0Emqd+6yu2ML4A8tD
CEV6Cw/TcGX2bBO38NiCVA1lxFgD8MPVxCScpf0TiNAmMWQPoAobLEBIeyp2yeV+
gzwW36Q8jjEeeNus0TKYxom0qaRsUxIHuGamrA5XN3ezGENT6nCf/WOT/9tP769f
Gq/ugPBgNZMgpNUgnx9/G4Dx9N3Lz3zNAYmLOicZKK/hc3jBQtHGhjmlAgGUbI4A
InpsNI0OmGfFZrY5YH5GcWZioP/kdbNk05esgMsFojw+jJLLihcUXgnDWN6Jtzyq
3Kx6BIZaV3V9jVowPk9Ew8zQfR+g1WTQ5P8UKjxuPrxtdbVpwzogpRa6oAu+dsAi
vczR3aOcxgQHxGwyk/dYZtun5MX7Q0+qhz5lnoRW+5HPkR8GG1DCTkESg6DC3Kq8
io5vl5w2Hbh5X9YjmW8rq2/VbO39TRsIAd5bnjXahOiqd5AAWVMZUWokfeSa2Tf7
RoLwJQN0YLblahdFcbur/ZMtmfHdjttr9FI8Ncxmy+y3W6xe+A6/borLQO6hli7+
0we8BYJKBXv3vz2LVYzb6i5cLAG9Nf7rkDSaBtaVP1IjM4CvDP2AmQVjhqK31ctS
jLshUT6gNxVWPUz3LiRkn+Dz83gPoB4JYWB2cW8sAi/FPG3Ckr05kWksQhD/0oak
gi90j2ws9/LIqZ4LQq7EADBeiAbU0afyCX2XCv/bSUi2inI67qKOr4k5Hgs+n/kW
oWKGG8L2H3NWxLkw5PUA0vqFR91f2B5YrS/Fl63NbClQSyVYJXo8XAAE4PBpSBxz
Sv91SzJPOSFAjZgK2lNbCTkz+yKxAFK287lyMDqWOqo4jqyNMjU+rFd7ILWQOD5I
5f4tvDfn44fjTguvvdCnDPpI1DKRYQTPjfKXITvYMmbCrL5iL64cHc0xBeLQazPz
b8nNziKMPtswR6r14KTs82zSSWw2tnPaWU+WHyV/NByQTjqfANjoY8LqLjAJJRAB
0s28dkwlbsdllu3waO7WC4PZxkIDZWJMqnJUx46oEEMpi10m3MdHvRYbD1pbbh7F
hP8ffHp8rJnxLmKFMg5MT56jVYOK8V+jPX12MXzdtsnBuY/xVX3AVx5hOvXgqBB5
hfslB/o7VfohtQMLqQU4ss52+FTuawem3r9gB04qpsNG+0zZCUhU8midNMZY1tiH
Nnnp+4bZc6a+9Tm+ZuAhT0s1Ph+gTaUfGuRjZe2o/jE8upgQkJfqYwqSb1EFsPwD
cYC8Df4aqA96bKuaDvrQyK5iR9ded8L7esEMTJkpEOe2qAmDre5hewP0nH3FoJuO
prvB+ffJLnuydQZ9UOJEvCWxCzAqZ2akZ+oKxnu/oZ5s+MKBP0n5K3vREMRshqDm
o8aF7Rj0F6OUhnaT6yiJJUFut5XVxLj1PJ+7omqUgOUIuD7V8qPiCH9u6r9yRWzt
Kv9L2s1Y/0t9JAwgxD5xZ5VDbMBKKdtkShEYmK/ytgjbwb2ZASvf0sm7fC4kLdDy
mKvorlsBAobtiq4ovEyrN7xF4e13oObpg8rbAczSQjhbqNLwuPr31wO8Ry05Hado
C1gyB4UQdjeLyKvsUjDkO1g5BcfAu31cnfIvOjq000tTJpgEsfZSix/06UxHfqCs
ptRS+m1eQclcUX/CkNNdMLjJ3kQ56k6qdDOcDHqvscCWqNwWr3TQJijpE46CXvCQ
F6Nu/yl/n54foxq6I057kbk4Oph5LpKIBfybk/8aprwq4kUmtVIhS0R3qQOQNGqa
5mL2a8WszRVEJiIYhIFhzA7peGNQM40/BU3CxJMSrks3ZeAXfuUIrv1olqz6+mrN
Wax9Rkw0KGsg4jCPsH6AWA2gD7TYmN3jYuQxHSgmGxA8+SAmLI6B+Zhoey3RmOQ9
EZK71PivAAEKEpTwSmaIhBMcs6M0cdWT5HBNJpA8b/+rHNr/Tn/6cYL0J8/9m8uK
8xgr3+9x6kbV/pbeZGg1dyjd8Bbo39tFGRsrp2mXCFURSFemBu/T8GypQjICPg9b
cnKxyqQblsDY4fRrqPvxPougKVQlpnWdxNMfL9758MPhV7E/kc2Z5t13s+kRw2XL
iT4aXsJNVbX1i/u7883D7W4IWz6H4nTrnzoTIafJmRb+jNf9EM8rzZhYU0BWH81T
Bf5rLSS/upzfW0/j+XUJTVfvIIyZo2IQaXvQT74/5tQ7PqavSs7aYJ2KiVni4qFP
SeuDjblzTGdE/PEcxPQcf/OVYzof0h0K+auvAoU/TSbWMUlk4blEhQZB2xWYKjUa
mEfk+sc5p7XG0B34/wYq5QjyQzYNj0d4bTrJ/bhJ9G1SxXDj1mO4ZUJYJ8Apk607
nIbzDjWdV8j/QneB65uUhaECwkEgky+M8H6zlnZjUyOcurv+5Uxu/4Uu2kWOt8Kk
i17MPjFePeoAh1AYoB2qqURDJgma+Yh1fw5+lclxCv1menpT+jQazUkfKDuYWCrR
KcfMWACvXvi0zshITry+PbCp69Oy/mAeW9El4hLLiK6RsgmHCo0u3WvBsNEjMKm3
NMrozQGYbh3Twq1MFJfqb0jX1wpbwps2vG0VzGkCI86AgqzVBaWRPtP59OcZpv4C
VapM4oi+9rsV2t4xVLvQHYe/vSQ9Kz6zXvkLfVGo64vyC8xvcKMF1/y7brj12o9w
XsVDFtUxuVR3dc+IddaCB+3tjehMyGWpacwWXDw6FeqJZF/vaDcA8lVfODBaAcHh
ytFOy30bKh2WGPnFfO/nUD7OunDy9VJkh3hgqGZm9XV8E+9JkL2ryraLXvJ52oRP
rpv7NQW7Ok/3Oxv9hQTr3tP+BNAOcDZ2NDzohAr3uVwjrxJlfKFm4jQssQ1YV9Mx
/zXj+Gb4gdecRYuSZ2iJn6hFyPueK2QG5NgPv65IHwRjfzaIP9L1E4BGlIthXmjS
pF+Q/IATbfkzv+PpwmN6o7IZ/5dI2jICJB31JhN1U0QUJHaSBij6E2B0wppktoXE
wDET14JfbIkH7XQvgMe9vLe569bALhq+jXYfQ/ewGhgJ3gRFD1832BmDXa/lKMrg
v1q4gLrU4JOzrlj8woP+S7K0hUrMQEJIJmrgSN/kBRQYn60QAEVtI5TORxjF/ZOn
7/ZXjaNde6Suu5WofNZfR8u5byeBgGJFm08ybLZklci7sUMDPe+TrtuqHsm8ldTg
hk51MqT7bpM977wGvY/7PRHcBsAnRwDA/z/0YQo0Hl+kUxV16Xj2IHb7LgJPnGqF
OS+cFYqjsBl/FV1lDTaLm2pOFYFVDsUZ2YSBGvZvuqxXPWhhd9dkrdl+cHYTvEWd
ikqG79RNs01YksqbI7g0DqMn2vmI0m632Q0rAUZ9EgZKCjBYwkp4Pkh31LyDsn9i
taIs8/DNI8130NbTyYOR6oJSBZcLjzdk3hO83zA8VmsPeLDjjax7JcRMXnl2fJH0
Gy8aU7LxZz4i9uqab+3AEWnD74g9td7YZsEbdFeH3n/WXmOVj8SxbyJ89Z8haA/W
7EM16dos566aDIPmzLfBZAxdi8dGDWanctgxN7beBzo+JDRrMazTgzC8pSCAir4e
TGCDXi7K5smhICB24YlmkS8//eAAoJBQ/wMswO0MmXzp2TG7PCwncnQPqjLwowFm
rs8rpRAc0DYYEPnec8RsjKVbxh0kGYFn+nfYFfZ0sQvjeOzLjHThjHK95/xUbglO
IGlySLs3Ym4fL8ztee58vQLo0ELrC3kmiIqtP4f2sZM9umOM2vCgnA0HmXt9I5fB
0igtEl6ElZRRQgjOppictGHwJ6Kk5mpkzYHzEKOSgx8dOOaL36P5LC7Pj6Vr4m8v
FeAZ/HwhOUr3GgpLQI11ThGFG3v0ZqI6S8SpPRMBWUEjKxiX9c2VNHF9MC5Qd9HA
5GgpeGMZoK9Vv8uY4yBfWDQB/oSIn4a8u0HUnQo0bgSMrgDqH7YsO/OQVNP8uC5h
ZfLe3n4yyat2iba47IiGIFblxLBwyWVPj6QGC7fq2Lo13EuLprmM3Bry2j7Hb6hT
Uj41WwYmgqv3I6MJQS1ba6eEaBA4U8pBhqFuZIrhfL8MMfiJgwgMylbtt5nYho+G
ynUpbwbWO4rg0bBcGZeHQnBBNJeMjGyg935Jz/vqq2/DXcEfBPASs7Uz2UAnDwq2
6ToarP7TLwZhOibEd4j/kSfx8eofO6ubiPaHyIa/mSh7Ek8NErteWj/vmT4vl+i3
BRu7inVyUOkc+JtGUk50S39F8ZXZPYmVcU8+DOC+riPy8iE+c3v4eSvzqrFsupgy
RCUQNuZHPI15zqJMVa5gWNrfDcYf9rAULMWq/uVXn4BXQXkhsgJCD5pwOev0HBlg
2OXtPY66JgsJ5drpcb+vlUv2aFFz0RSRNSPegU2koeuEUw1yLP179zUoUnbMmp2k
JrtWbk/XDqxr+n0dUQm9nvH55DdtvWASdBgvZPXgdknaYIyo4V07zQj/ZBn1V3eQ
aLf/UGi6H7xkgB5lKOtOqJSjQSsS5ADx8pm38zzZ0zJwt7qqwX4OsGXTCCGoMJ7o
vCpCjS66uYZGu6U9uOvGSmNE3VtlS8JrZ0H9MvDe2emm/lt8hdZoDT1FPOmGH4qd
9nreJWXhvu+131+VD285x1eXCA3rlrBztlW41JI6/eypQaczYITChlzZihhxxcYH
/TPjruaT2eAmESe+L6683yznegUfRAM233xhqHve7gCkq2lFOtKRz+t4Du27ZmZ6
i/5CbXdOdcv73ImLUfqSc9KPCQF+LP5+gJMIDUTkWM/eyRe1Xz4X5jDkF21oo4l/
C3Q/IavoST5jlyVWBIFIiemF+loog2oC3ACpELcxorxCn0xI8p/0vacBLylP1bEW
gW9SHUlhQxpbr9fydJLs1FLtBlrLQ2h+QrewVeD2XvzWOlXU8l6o8HmhCTSJhHzN
DadHqqdH5mShMRec2XmBNmavt/CqfucKPwqPlVTJzRrcG5Hd0k+QCEFkCoKzpKG1
JUS1wOL+cZYpChsX5L7x3xNpuqZ3X8wBnUCTb9bb5ZYalFepje/WZkkJ4F03mNyh
TykHwPSeKtpDSs39Afy7LdYMRIBC5Ubs+VHAhdk2806a7Z47ntgvSrlTe4mT86Rl
Tmkb+VYHAHLt+GutnTJYNAINRViiGCsSJumxCNSPCeTSe4KyO6C9r8huVJAyG730
0nHn/aDz/IcsLoNf/X56ymexCYLNCc7Aw34RzWrukD7K09SNndGf0KrRpZ3MiA+v
iNNteFwDm4CkqgxcdF1nf3I6PfeRp7jhHsubr3kLsbG11wcWgDto8rSFt0ncxobv
eRuISF0SSJ4hGRRxmGmgsUg3mUsoMq0fqPwD+vhshCm87IoJcjAlB8OSSFiEqPMC
Um97N9p4tJWkkRBDUQFeleAl9BlaXV+XPzh7QJko4DtAahcFgdFs8Dy8Z97vaq1x
dWbDPq0Ld6gBlrjrPXUbXq4cfggskx+qjIZw8DhaHrkYrOTZ9EBbpP4/eqGGJkW+
ixnAX9eQHYKwJcUwTkGuNuR/51fwOvU8tde327Isi8P+rkGQcfV02kdHYQdAKSnJ
UaW8V1vi52ah7S06RO8f2vdeIP27kOcM59+NCJlWKaa6TfHzD+6LExUNoOqfwyMA
BxwdJYhwe2iDhKyOR/ylFLaLvws0p657dLCr5vNZmmWQMy5qrMWi7bG3Astkyb4p
d0m3Sbtnoh8jBC9GEbcp+kRK3kC+LMf1iUc+9JXxC0hYPbE/bd5CRaqaoEflQaRQ
VOu7c3Ura+sBFLzbrm6x7vLeLqW5Bn6LUt+UHYTOCdZNGbCUIoZQrON/0TzEoWVy
tb3yHy96tEQ8NTxUjeP5p0cP7glH1W353JHbVT0eufafo7o6pRBrXUFnNhJgHCqa
iK6YCduMxMSm8QnJ34NP2Jv1GTZCs7eJYHcb/iIjAMQkvMKZ+lUaRBsSumv23q86
3dMAJWxh4kDat9lNaPOJgewj3Hc6WHQXTtKQA+eVqKYXRYfcK0Jdf47eHrL6uHs1
zMXYE3cxb1Mi4/+LukZdEWev8DLGJxiX2owikx8XQ7nZJs9xg2xhGfXFrHOVPYJV
HoakcIgd+A4m3+FjEe/1P+Q6D5wuQlwM+CoyzBi/q+pMMuPbFDZxWgPpEogOGluR
4gWpb30WreP5XsTmxTgwtUCxbXAhO7SUEcFh8eM6YftQwMf2lVl/N5wUy/MZejpU
yapfkOYYUY0fV2nYFtDfCoo3o4Y1hGhc6xPoZH/zsDAnOr/RQOy9BJ1huL5e+Kad
5x7sKmFOJYqWGRXFuR5F6My+atnvVFo8AXKxHeMYaaRQvJdaKgzalN+W02oqWp1i
qYk4ZwoQzSUSo5UBqNsPulwWG0hy+T1yPWfUhgaL23gQK9msSuSU4hugsPi+5pWg
tEU0pfI3XY/0LmVrpQYjC0AVLEk2swDrZ4F4HHcVSfhnFxKzoR1kFt9TmD8QseCP
kiAGPo+iT7SW+OTOkBGmFglyY5AFGybnEk+B43buxkRasjGjXAx3G+rkrLWjcUrT
jyDUAlQSA9H2eLmrr0hHKAEWW5pquP/AcmMnsw22vNlI3IqJvIhfheBJQM/+vTm2
lfTcI8D9ngQmbiy+F/kKi8vh7WNysAob/5+vjhVGnCI6o99sbPQFxFx5ksq3sUIb
LUhO49/Ocp9w2aAgUxJELjgjawZCWQFclxXDmotVm7fi547lrq4cw0XO/a8rhJfy
eCHb5o1TwkyeLQQy3AUNpryGWO5XXX9C6+iyrNBTink215kx/IjJ9AJQeZCRRmfq
Jz1cpSL9ixcsuRthUkIky1cswz/uuQdFtDQxCXv/9zQnvdFqz9AWNl76dZ/Ni04h
EyagsScs3wTklnG9D0WggestJhQJLJId2xPVwFGyut7E44zyYrCA2T6Kbluj1Bx3
EppW8u7mTroZopaCb17dRPCk/kpeQVQ6kaaYROHSQWyTk9+T1ttF9b8a4cYrivsl
YoqgMtuHjXvnOfHP4PAp4VmOKAgHGnvxFYIqCSVieClAOU/FhtmUJzaAx4hnK1Wu
cdDt1HFEavg5Kj/Ge6P8EeU3fJWlcD2B2GGRIGev+uorJrDjzFdVS2sQQGJWcO6r
zYvqr4or42EOwbHNqnECcz69/DNRy+/5xd0sxD6EZBF7sBZJKJ75LfZs/x1xogCG
L2czOsfFzQdbnEMug9Li9V30dpsF6WYsPYdqUVoX4wCUN3gxOEfLiDU9qws4c+ND
i4OHIbDUuOCtu1nsFhUqkoRhZ8xkIqmaDpj0LhiKPp+E/KrZqoK80rQu+npadI7W
tf9FzcAkKY8FROGjFIerHVc2wdGdy9VyDQ6djyqnOl6ihYyyRXEM+9BKmgrhxQqn
AEbnpSsY+2M/ZaAQMtTy+vOCXpDgs7RIgSPVucqq29xc01BJ+/bKdUUqjt6xhN9g
29zGJrAsKUNpYuv7m5nQt6FkMPG/loEWJ8yYquhP1PpelgPCtbWgN5ZnFFuPOeY/
sV1lXZjvVmTB92c/kEggGtFP2v6z5delb+oVAuxytUSV0MqreigQ9t0FvKo3MY4G
q/Q+Qw33O4dpGev9adedcyHKVg46zi1UMei5uhPdBp/C4d0VR8JJA+Ngfpe3f1iX
Iee3t0QYxyYXhsjCInsLqU8LH0dV8KOXcHTa6iGsZ1J5n7CzZyMAif2QoQhdtB1s
Cha6twbCKTSNr4wn03tEDmCn9M+C0muUd6FNWy0+MB5wSS4LytrsFKyR+A++k2tA
6Nvj7x12Uie2P9E9qH83XO8qasUKm3yP/HlvFa+0XqYyVRgZodLKROSuRJvgioKu
zhhe0DbRA02o0CaweVg+3vDaZ+x86Cwqg0T8dmUNN+ALoOJ8pS0TB3F1pz+vrlPj
DqjdyCyG34h07saeJfz9wnFCece1K7ksmbl8P2dxnx5YRycYIzOBRuUNGjQblW3n
HZK+lHBADxXuYx7luwllanleCmCzCMbaxAaXZ8Gx3vdnG+zhhEZkSE6SlxuYjEXA
iQ1ulOEQzmij2SDTIDpPmO/KBFL9ke082f2j/C/htq5kF5EplH++pyRPtk0qDiOv
fWmOCFS453nOGUzsSe4wfVigWtXdWvRsOwJzELMYD3PtSd/vBpSjtO6V+uxde/by
ghE28GInKAHoJdp7/SUblPVy628ToMk40JbAiwYg/8dFadF3DDeIf9QKXvKnB/PU
MgrM3w/0017eDO6Td9QzgJg8FILqgaKBS3ZUmiPvDszwTyvHm1VRzpefnucnB6L8
aeChBmJltw/ueBrmCt+/QNh8/aW2SXbCT2fqiSZ3jY5zVp1mV7YkmoaUWHrljAK2
uEWzrj49gSTyUCnwdVty527dtdi9VZKIh41QSwCekw5Z7FB3OHhV77eEGaNR0EgR
72bdES9oDhM/jkZ1/iCE3RAxmTu1ihL6rnASYQJi+i/2uRR/XuI1xxB2fYDftjUN
e93yrRtMe8jryZ5PYjwIUNJsOLVo7Bmio8CKMcEIrgCHAKdq327X9hEdEY6fI8S3
ukGIxFQBY6RLQueTCQylBAmsTxRj9jZ3oCwYyzhjNaSwzzrULMZNBxwiZa6HkFbD
YH4E9jpexSZc2jvFKFw3DwUa39A6DizCrhuWwKX+N+OrtfJOLT/reWlUsGDTgDsH
0ylkZtFIWj0AIoFEL7bYe/MYhMuyT2yQmP4t7szdO1A6CVtD60IFNnHox286MilD
IIF/05oFW8TSR8fpvmS0QrDtoIn0xEL4mlpt3ypc4ZEsPYHRYaNJ3UfX0m96bySc
ew7v1D6d2hrCqVu7T++n4sxoDVlgKEj/4aDU1p4eOSmQEN/jqbOMXpg21NNtTdYi
`protect END_PROTECTED
