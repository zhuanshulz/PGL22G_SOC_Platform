`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oyyNuXlvExOJ4vF4LPI9R7ZWbDpypC3pFUDoAN4kNIkwfQCRUJ0tYZEpgiOXXGOJ
5EhgdM8xE95Enj95HuLNTEQ8EdIjinx6AuIpXTLsvL7T6AHmMLaHBcKu87Dbvtuz
Px+VOC9ChhJ15U38ECotYy++GBJtZeUaSzQj3EFGNU2WpphZFIzPm0QKCxk7MOPA
3Rzr6gQrIhawdJK3r8KtZVYQ/ryCdz+389jxPsnOfvIif+5Va7ES1e4UKWEPlNg6
JrTRCjx17VzYmI8pjj7stkFkgVDJoZtrukse6aE37DAh33MkQm4mQucyJVWBSSE4
mXpSe+sS2S82q3H0vJor3dVURGBrzPKt5zk4d83xbACQtULI1S5AedWMQo6JDEan
mnfPzSRSdh/uh4+I+UKte48BxnjlWrRh059bPHALqMmoGsc1HwUJt8c1BwoEPGAh
2yZ2CdiVwLcGUcxeCTagFfT/8UFUpOvnLLBZKMIJOM97OxunPTEKQa8kEaERJcC/
Ln/t2PEIQxVPe/gJFzpekzVJptF512KInMrFG50oqRLk2LPqxCslLSCn9hFAAaJF
OiIzbS7FV0DSvIF1k3dkL5bRoX9n6c3+0pfwIM5g55Vrz88HmKaKUra76j3bSt7C
qDy1FxqFCQzoc3epR8i+U+ECtNN4V0u6+vIZ7sXUiUlpEVvPpKEVzTLRBlIOwNTw
XFMZZIGCU15V/1ZL/uvL9eEUt2EIh3pBsfpLJy/jV1LciTCK98MlwJJEp9NdZOO/
OGXp/820T5Jb6GIov6FJuz95gDgSCnrvy8LYkHFHklaqjebF1sCDdfwHjpRmTo1q
YASSw7qyKm/xcYbSk/1lQzSbyGKe1ah3AoMZXkfSPF9E2HJa51xE3V/wJs9hkF2n
D2fv/JnPkPESaQigwH7foprjyt7+QqcZjBemcH/kJf97vyrP9RvT5tFiUT/ErEaH
qcBBUWn/R+sjFABMwE9u3op/5I/mnPH8q1DFPMAjevXn2ICP6W0XYC0Or7UQrxVn
6pbTDGkb5lwJ+5g7zBkBwMrUrMPHRRGL7n8dsP4iZZ1wyyZEB1cdFsCf635Q8x87
3wfHW6evhEDeiTk36sD6YaF0AFXz31HjVugOFLHJxohACkwyGx3M3ZpDp5YtT962
1VSbJPtkUoreKy3WibA3zh6X+TywFYWXsQU/dFnQoitSrh4UCbENFfdJOV4FUCYb
3672fTCYaUGxpqmdovp3KsaNUO4DZ+Ggb4/Llyk1JAI7UyFGv64vG/n/xMw7ds9n
gEBs5JWFwd/o6KVbFX0ntIlN+p6JhzIg6/vAFZHIvflai9zWdLvnS02P17J7nYsH
cmMo0whrqLVnMzuB3fI2AIjFyG6DjxdlphMWGJN28jDvnsqOsi5p+1CKCld7KNeU
luduxRXI79k4k5Mbr856YGMtxxlq/mNEVN9UiHCMju2XOyZrm6qCNaD4SzuA4Ai6
mDEsMnDMHLDyZzSJbGvh1dh40kmELqfKF0HWcTW3ZRIgRthkulbWfRZHdmT70abV
DuACgq5ZMHU1ybRK6NNPt1/VGccmGVIAtNiWQS5nLl7EGrKg8KP0bNr2lA+49uYy
HxDGWYKE6MRvAx6xUW2xTgakClGnSy3hvTMjZbiIttsEirc4GJPNK/X/8tpmVM8v
1CH4forreHdzzv0USjRb/lqiUjJ2Eq8tDLkNDms8Zzk/tYsItzrWt55PrIrs2u4x
8fQeHe4fd8TxQZatmKSFfYmru8Ep/j0rAdg11Qp67KvD7pM8SouzyW6taTROompo
psErE3/trV6jUbiO66AXdOMH6D2L3iVMeAadPJUCs7fo97Z1fAo1GAfykoJA5QnR
mAp4NaKV1aAO5pTuFkt86isTFHwZQlRp2oHW2Hh/3Bi3yJJTeFfe/Tmglqq+3yIn
Fic9ZhPTqjaHYmMDi81HX4qRdFoybxT4DTEy17iYkI00kEZ8u0C4OJ+QZEKUmu3h
XK4YKlyjg85KKDYQTUHA+w+mzbjlgCMaaMQt6IKqJ435m6LMVh+/qE6xbEIqukTA
bqa/IIlJhLGSj0qifH0P3ISsXX9NXgRR96iavDfGWPgJTKJHQcJeAdjFeGS9iIYR
CEI7PBqHsLpjfO312tXEf4YCttVM5MLg9IvtG6UdO7KNq7fjWG/yg/j9Zrp2DSHm
Irzq1vMUQnt5roiYFhrWpXVn7EpRiCg0k25JTV142qfrbJVtQKCUvaY3P3TUBnfw
43BbYChJdBu6kYiCpXk90yHtDV4tLcXSQThms/grbXx+y2CaXe/a8ICuQVaLUWYY
jN+cQLH74zzgvCzCvTn8lMzmCvIGEaaSLxT4e9B89PBmk3Lnu0OCcNDVaax2unFg
QRynQ2lGQ9fjgFQboAk0TzMnd63vz5/GJl/y3FrG7Kyghq4nDoVr8q5C6IALfSjP
Ulz+R1tEEoIK9Mqgp14DZ48wcQ34btNCkmyce/ewg5X17LhlCRUXv72BhsI0b8n2
jK/iBxfk/wj7DD+RM/AFmjfCV7Qtk/JBYpT9B3cAHcWOB+5i1XAZnQxigdLrpe2S
4vpDJD0K8yakIumvlJq/HDJoh1cgictH3bHwtkdULUqGTUeMUTIDd12uLCfBjkbf
u3M7rxYI6eeuoKjk1NQ56RtQenFjPxROn4OgSdtHEwpab63zfJmrob0uv/eWfwzQ
aGQ3aoiEyP4JIzo0r0d5hKpG2fIX/Pt9xJbaW0iuFe0L7Cv/myJ6IWZmZDD5NCJu
0TRffYA6uVNG9xfAOXqI2QgCrzgNksV6GgHeAczJT70178LqXXseaEClPm22NMnQ
Zpv2SmL/TOoA/9Wk/y85kPNimbrJv+ZjD4BIiyPm87CHcHcwlrlkK92WNdD46FdH
/PD8qUUdHug1IeDyzt6mZnE54FLDImi5NM/trPu0YFGF027aq9Qxm3lBnq6Rf+bH
Q97EJ8AGl4bgucDKfCG4hYS3NeiX6EyrM76T8NDCr5aDFV0o8SCMRZAyowXCp7bw
OAkFq1oINMETc6i+Eox8ehYFXS91aArsoL/BIPvyomJWUh7lmxCxEjDRpkzugneK
pp6y2+RPzUJCXVXUIEl506Wvwa+RAv0Dc4r/HIMWM7qfCShNDjVO7LuSN07gpsyO
dQfxtnDmz4uJh6Qw9Ddk29U9LlWH7mE5W0M4g6lLekLH+GhPBmefZF+qwsC879ym
hFRsu3kcT8T7IM6cACv2mA4MmhuHjS1SgHydq+KOCKKzm2xUwSDZZc5X1nsz/HUF
MddzVMXF2Y6mwQ/plJj7CBoLW1iWrag5v586L0W9K0FCBTjmXNd5f3Q0QGeoYv0/
0jTI9o7x1wrUPxPYOy5zCn6rfDUt4dsRokkg1JNlVBA787chQPpdpnThVzEXJLYF
/65flvNtLuVoBnwV4KLB8rC2ZI06hNl9Rg632vdYf9LqBSgyz3EiAvAGiKIm8ZsC
T2WNHhzqHdf1HW4jyPVG7NF9kXVO3t+UYKCwKZu4o6SYGwnqemiBOKh36lOGCtzE
pbfNRHQezBKCdw5I2tmc47Qg+0WYuIcTrfLqE494VoBcjLfoHXaxhg9JVZmaIUJA
AFkPPRwjOHCVyk0t8NqWW0ZtGnpeclwsRplOZhS+otE8Vq6pjRlRUtC90XS/bymB
Nm8WpjzNJY3PF6UQ1wu7xm7UVHf0DNHFdNURih/jQBRFpu0oBiC/vn5nIkVyraqg
+SW/mPF8rTEsfmwjkQVzY+hDC/OzJvLGACD4A0D0E1oGRdt3e21ZXi3SRz4SRFuG
EM6LV/Qe8yCk3NyW4dJOlevLV3mrma6R7Tr6DIz0kyr41slTIZqNbvUO+t5mgVeY
IH85+Xm5ZYmYX0PqZz1RXjGeV4KUlZVYkMvqa4fskBdmfFs+we/uJFLa6Uqa2Ut6
OqjLnApHh79ODwcK5qnE2N2LHozDUnapMzP1ujhwdSjRPU4s+VKYov4CdQzYE+AT
vEIuOWR/faC1VjJ2WjBCdXICRPW+MuD6hzcpXOp5xnMNBldShfderBsNF4ua2nuM
BUgdQU4yB3+duFroi3SQWRjNCJFKBvf47Mc5YMxITQLRYZtz8Yzsgbd03J05UcqC
OR9IR0ynv85SsrSn/ELVpuU16DVqCGO+R2QaA3vLFy/4Xk2iqts4dKyNJOefGoDJ
/iN3uwzDLSPqvq6J9CibOLf8uy2HvEYwEzIEfxPf7vJOGQRIYLRU36PDhPuJsnpo
pBfGn2Ch0VWee+Qdlh67XKfslAwIzUEt2wWUbhsxdlXC/vqjRNkb4UHGpBsSrmiK
VgGPhosdV8TsRrQCHaTj6IRbEE3DVKfdwxFQ861hI7wTw+lhWE3mYBUkPzueSLpe
a79l4kubijNVGpdlc9yguWL87Nn8Twki2UDP+vt8OEplnUqM+KaYi5gVtLl9cXkQ
diaw4K3zNRtOhGWL556BrzT9Gv9/rVfbtFu4y+wH8F8j76uhLpHkEnJffOjJGRC+
yYF4GdDMJYD59uh5XfEgv3sU2BnRZm2WGxeD2yJeBb3Ebfr1sPeqiMofxotATsdA
613Nd+4K9CVg8uC7nTBjJQkAd9pyXESJieXzopWoaijQYAuP4HvzzOEDoacyfI2l
kFmyK+us1Ex4F3ZsVkxvDpL1rrmQ5kfFzRJa0QJmLivg61qA+DMvkBo+V51WxVA/
14RA9XrTmgSXlmvfYgDBr9XU/56aN6mRHexltTTb6mh+9pydD4xFM6fAILnwPdnR
tUMmTzzotUBE53H8GyVaHBzDbLJ106AdO5j8ZkYI78/KeVZpzno2Uxmy942IB2ZG
ZhoK2TVFDFhehP4/CeStx5X0SsByiRB7WTOy9AOEESfpslOq7kHj8e7oEM/7N8gc
JL/yzPQvzvPAp+R+hKqPpLD753G5wxw6ENmyoJyOJWEdvCqQPTwCv3HIvf2LAMGX
+4p6jHn9xWl6dQMne5Kg1A==
`protect END_PROTECTED
