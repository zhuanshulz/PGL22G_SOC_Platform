`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VyogRrUjvhVyZqQWaYWUGnJwqK44SvaN9khMaQwxfQH0UcHcU+dYfjzQk6V6mNrs
teKrQQgSb5gPHxz+4C7Q3GXktrRZZji9YU0W6QqJEhRO2JZFu4XefGlJ/ryr8Pfs
or1GK9aWY8g3huFmJ4vNgGxYNE9wizu4BW5iHSTOMVD0UGpVzCWVSrEfIoIzyL6C
rBc3ZxiqGzVVsWO1IUym8SkwvSZMILec/MCvUXZ4VqUiNfLoLJ/GTcAqd49jh36n
CQY09416sW5kuByAxnVnYzEcs2dBcEMS9mG6cqkOH43wu+DrCvExzr3AV19sy4ZV
UPtELQx1HsEaCpE0+5TwJHLBYddhvQoW7bSQVwB2nEvdZfwars43G8eVDxFL5nL9
JwvfKJuQRKvDySk0LwPzw9P0hGzTdtIbMg9oiaO3Wk/2p4oFlUn6EZaKFUdzt78w
+XYTrG+4j6K9VNpZp0N4UnkXmhWR40Akke4jmYs2JDoz+vlROZ5EbTuQ3p8aiHIZ
EiTI7iOcFdc1u+rHSEi8qxZRz4gaWtmDcZ7dGABwvHbJjJNy6zV4mwnJDKuaQBaY
FH/NWBK918KCLF3OoViV6GOXed5l1f9rNbwpakDXspGvRA0+MHNdWRO6v4LWFyVs
e+giflB+/6HmcG1l6cPabm/z9J5/TUSsVWDPuFkbGkKkHDRaS1M0RFfO3/uicGZP
M6uun5cFeTFFNyTENOw3sUQfJ7GhFkELY7axKB0rAxykBP0p/5MDVLZnPKPCajCS
o7Rad6pFaXst79WcMdv0pE060JUXF3tpjhO57FtxmNeU6B2OaQh3TUAGsP3xFi8X
bPxLncb/08xXJJZBoueh590FkPhNEydfhAwWtXULc2u6zdr1f7A8pnLcLIVxD5rD
3qxa9xWoIm8iTtXCaax3q4bY2Qf2/EYIsnutFO2CUm2nJdtZlk5BRWHHc85ORrCE
Aukd8q5HioP1BOjSIBA5reUhB/awa4/m5gLdHmaOuIZPspiQsJK44sWkDMD9/xmg
QLcs6GgB4SMTxSXZ9LxNgefalQpgf4PLeaTiYhQ6JYWJvNCekEZamEtkW41H0YRw
jUu0cOT2O4YLfY0m8nSoVqrm++o/TJWelLpfaW1DCRZHzFmkJO0Ju1lBntwG0Vz8
6PodJIvSjG++5EAdDEYIe28xh3gT0IqE+zki0QmLKYpYcRY6RPHAkkXlthVooIrF
asu7HjWr4QVFdt9i3McOI0G1ih+ZJNskHyQf5NAilsz7em5cL6b08q6hlwFL7aW0
vqh7O8/neHboNvLFlVZ1WVlLBvyb+BTobSN4XltIJt4A+9EQrgxemdTmdqWQPed5
coBEhfMdu7YVp9Tqlu/jEXVyNvsCDMuZjKsdX2dY0T8kVpPmocSvt0cQB6L3OF3y
8rWIrPCTSgjnDe4mw2EAaLsVXAVdSArfp+ZRbOCckwN5gNSBV6BU0Q43BAcKaX/A
DpC6nQxFYHMsLUvdOPHqSEJfPWoUcQgiIwy9vP8myLm+M99IB688pfmXze+KqWHm
HueV2A9/c4lp1y1Az9gZBAvekY29WzQwbvHu1Ptn1J1CRZeQv8FMdp6tJTOsqPM3
xay0h6YWlNyFsoCtrgVeaq6pg4VZB8ROO4RyMR8F1fG7UdQt6MizipMOlc8ple18
QYxnMrW0q2MBHMmpGm0mTpxP1b8H47ieQGXqRF0DPifDH4+6WQs0+rBeeRkrrlwx
uC/+4kmrJm9CiL41mFox69yjWdIHFm9g2+9xhNPn2Rhoogw+iQmAzIL3mIWIlnTK
E9ZjJiApRoSwyt4/NCPZxJd4Y2Kfz7Yh1X8Kz6Mst2lcaQjo6nCsz7TAHophNP83
aP58EOww4GF/mQtJxzZJR8UisrU+kB1JhWrB5QunXcefkHJJIBHEnmqV3PD6IMf6
cIkhGP7Am29HMDlLNJWGbImgCidHWZbbUoZD6z0eBQgtGCk8D8MVlGy+q7WsftPQ
fapR5XnZU8ZZRebuydv1dRN9Bf2SObljYb65bEl++u40aMRvH1a2+XJ06ueTH/3F
WSZCgdifgLiSfq1T1gNOD7Q0Uuw9fggCIkU1BbPeeASCiBwZklnpJjIfPBfyPGGW
v9fZhfz9mQV0Ce2gU9rOvnVmkJ+3O2x7OeKgIdkCzTMf5nz8yX5e32ej4Y9E9aNr
YuJL8OjBlzMDRVAb1UdDgs1MAOGx/IpTKSGVrRju1Pb53UCjpN+0c8z2ysZPUV4k
DAAadprQXNZAfp2UgoS5EMQ4Fvv8vi45OS5LO22aYJ1Ml/dDkoAKVMyVgPIkBXNg
kVauG7gEZMHIFlFvGvOoDjQhl8m7qTNHoo+rFhNWWYZidhIhU7n6M4FK+vANt1pD
YCeLzYd5mq7Sb0Ii/XJYCTQVmmTmdd1ztnmhube3a1htyklDbZK7EBGlKKl6yJnV
4Oi3nv0DLTxnyI5gkZ24dAM7arN6fHALPmhPYeHPlT+EdbxOa/3QvUC/fD0inWWX
vsRWUnTdI/tP8E5zA+1haigmNbQS+//Ml2KFBQd4tlQ=
`protect END_PROTECTED
