`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7bZss+V9TyfYsKMCQRlIOLwvMuZtRYRNn8dZZLki/9dhNPXMmpKtAWlwW87x1fdP
xYLX5KMmO4EiEw2cF6hJKze4LB/XLBW+6Soxcd7pEyxoQq/uyi17CD3KzVAtIGNh
ltcjwa7uw8fKjlKizQBjXgpqLDe7IZKUhlqbK7d7aubFg5Xha5tKuOG4sd+Mb66D
VlrXaK1gBIv4CLnlF5KWMsK0Hi1EapD3k0JstgIIp9lw8O8JFpleFZAB6MYOeZVM
uL9NwkxPeErDqs87NBWke7Z3hq1YHMX171ZS8qL+ELDcbAD11CxJLisQlmS1bcYl
UXRYwBkOHPZrgr67pFeyGodc5OBZZ1eDKrky7d5IoLBDCdNW+QsXnjYBbKqz/XP/
FhqrlG4MFV4ql4GV/4LgrBb4V093LqKZR6h027cdDQafDwNiXVfb/xHLz1478LDi
cmN63hPTg8Oht9y6zGcMvxIosWrU/gIMaITHUhibroOB5TncOXUqslU+DVYFl2H/
aw2+BUNC6Ou4wgJkvsfSWoGLALVXWdZbnaGpZWmW5IRjHdv8lXdL8drcyhUT/qaZ
IlqLIpwtGJntbpxaqVaXReWXx6tEgoJ6VopZ0lfencNdjx2iL+ShkBXYCuyEtQDP
yXLfuux15bAsbWstT3BhelTAYw/ggiFEI/ubwdDMe5pQKFjpnTUOk6PMBRKIWoEi
EK8TnLQVF8h/tIxE6C/D3sXCYhANu7M8LuixOvM7og+nNer/xTIu2etrw26hu8KW
qzIoXxS/wTTZIjmVz/COAOcY/Om8I1TSfl2acAPjCxC//7bizvUIwnmzqkwOgzZ3
cTmrYlPPA3LZl4QmCepRBEXlDAwIqyfY09WR4aT/ZH8jIPw88nLZppYqiHlOqTiy
ZXvQsBb6sLVcw8orADk3xDJsCH/JMdlZ6LO37Mj6iWIVjLzSrGUqXl+Fv/DfwNPg
NFtWlK8mOwIqrXT5IQLIpUxM2rqxN19y7Ydtqe40jAdf/dM4MAHLDHQFVasJmKxF
tnzW219hRJWwnmPaZ/CiUy3i0bsihFjdZ5R7Bvczk0Hj7XBumTDhjaY9N6WaPiEe
i3x3yHRZu+eth2zokYa0GWSQW5J22h6T0Z779KsfAHHIJ+BqxYdGwcyQGhmdLt+y
rPeJBqLc7ogXxcaqxiKl2t/pdBJqPcX1+ClUDAguMao7J3txr+mvqCHUwL2bVrIB
PvCZXi+wMj0sntYp3fXJSAWYa4+8MWr4s43Cc3peo/2BAEtJ2lLKCHz482prhqdR
tCje3ajaoUCv+yLDf+mmajfxySJpfz8YE7NTUp0MIRFh5ti+Bh5bxF7luqkhAyd3
N+uEHjamci7s3/6llmhTxwtUc3ceKKWZ4BsenBwxA7ie0itzpyiskkbdKoF4YgKM
sYtqD8jMBT1TBB+u4sL3xFy6pdedtE3691cH3huTPIWZXTXqxoFuh7QGcbp9Annf
PF9x61UY7ZG7+4yxNgmyEInKpbP4z2mQs6YhFB4V9cM6/bhp9iHsjBp+vrj2E2Xo
Cx5Bf6ceRlR6leI8/tPS+f2PMr8tGC/0VC037AlfLWrkjlXyPXCMoIXWchuckD4A
LiJ3JhvfNXU830kOJd54d7uVsZCzNJy7fEUOf4aDhHQxableXtzPfkXFL/RRclsg
EJBytbBs/cQZ98SMhkyok7j17Y7/b/HcUZBYbj2cd9vyrxvZzsyrqGs2i0Kw7CkZ
dZsafNeQyGdFspUq/celK1N9XuxFYByBqgoZOrXVKdL3MhAkZSvMiGEUetLSdnzC
QGsFDPEfirzv8YwGLy7hIfiip2gsIOyjuRyJ2mxKUipAuu8U/gm9ByAnjcrTtyHu
NCUsMHgSlv6XFlr+iZCWYb7+Yu2zdLt4R72Tr5GiuYkIESxaDNE6f5dUns07gUQi
bCFB+WbG+a24p9JtSu6DKlvsbF9CXZM8VLCjGdLDe/z+J7e2QXNIqQbynULTOcf+
AeANP/j+HSvPNjPdjgRj720QfcklJiR8tjkeAcGQMdQZdWE5W7Tiv9j7/kKuj/0O
SzMCpX1qxophdEWPQhrT0PJvyiZ8ka1F25fecgV+2sQCC32SZ8UC1yaKSHg5zsdP
if50g63rGzavGPNdSzss3O8fcKHza4fvzpj4dVOjwVjK+iIpLyda8e/agRMXIbF8
nXcQH9oB2BK/MCtW7I9i8xGN8KVop0reJoNLHpev0vGJeQKrbyHi0inc5z/y/tqo
a27m2+H5J1WwiesB0CE94d2/IaDosujIjm7OCazl8ZqBvh58GR45VO8sUgcRC3Xk
zc5qb58sZuqQK91WYj/Dnlozn/7qpNKRiFSItwSAfVxw+dlMgSkwjnskjymMj2se
zjUMTmv4Us3W3u7Zf7JEbnD+V7kqJsc8H6mei47sUy9siKHkLLzs4+ju3wPLJYkQ
zVcLpZ1cPubiWpAJgz+L3kpgKRR+z9I3GkjW4jKaFPy/hXJ4f1t72GM4Nb4NWdYY
0zXvtPQ/FmuXfjAT4vpHF+LdtoroW3dWl5jsxHnf2ya/C3zAPsReh7/DKZBF03ge
`protect END_PROTECTED
