`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zdYzdwEdNL+F3DVMT12i4thAG2jAJLo4zflKNvlLqJ9VHNyu8kkdm8jLtd9nRG6+
hxcWIQggtIKHBb3XyYylnVObwd7idEq9B8mISh8nD4uzR4GL0Cu1nCOKn9VKrbFX
Iwb0wkBGVU0T0zONc41U1crlHQLQY+3XwjT8tbs2TqVDl3IWM3B1VCPqA/+fLICc
UFeE7TYuTi8UxIAsLFsGKxlkuQ2C55alcUbfKgGYF0T0F14BP/UXIG2doHuDFKXM
vRxkOTjixzp59PozVzrAd2SW9Y1+e8vf1X4rSfE/l+Jb4LK+Awyt5Vb43d57ZBgQ
wiZ2G4r9E4t7s+BUInvX9AGLcHhMKKfRX2uIbUzjHNUmGyu9umG2HfDjAfhmuQZo
IcmpA/1pMWVUPuN4bs+/UrkBUaz1L5tDRRjPsTmACtbzJScXB97XaflYUesz1ZtH
MlL9mV4FkIV2jGKT5YIPjtrZ1DEHcPcJbj9rLwIhEo/z3/vRiaJ2I8619PJ/h24E
alMi5kQs38x6wqH0IpRtNXVI+ZQcWI2YXGzRu1uN4SUqg5bvg8jGJ8AIYZh06mQN
+i8BcW/S+fvFVJlAGbZb8/8QKZFPBBUjMFx9xvbfRc70vq1YE6CcluuSDzqaCRNP
4ETuxLw4+Hgz+AznoyI3su7a9rnYwd84ylkUYjSz5mVEq0rgVj8I4WYfN1WtAD8M
M2k4yDM+PnT9UsWkFCvPbvHnKgp+94kwnPAv5FhI0CQYpn7Y+x1B4sHdSAJPE7xM
5fgYS0VYbecVM0EVn165YEsDMB7BpqlVFpStMVAlS9k77Rx9PaTauv09PlOz9oJU
JNm7LDyLLvsa+ZgSQggRWI+6BGNR5b4653b98ALdLGQ6WhkYFzOQuiBl+lJowAq7
1VgcfIlFgwhGWY7CeBVKomdUDIkduIZYwCbtvhunluMQd4S4iPPJ5tS1v2ERjMJX
od/ze3aMwjMja5hmv56JzUMzlsHLiXDpVtmKMiREiaoX2cV9+/ben241+fTSKVgB
zyJ2h92t5XuQd1CTDLTyeRbuXTKHlXGn42gM8kRp4mX07hXQFUjARsNM2KBesxLi
CMm1X5L6AzWg4gbQ4AwSP0LjI62C8ahZSYOdquUgB+FM/cFdEjCHW7pg/5DkiBtA
ipSw+iMYno6xMHTNeNEhzwFQhYHUstYPjaIJryPnBHidPVdaphEAW1HYa6XLpccq
3pKq1oGFh2nK9HQ5p7rGLbWsIsxslaeRw9yGNfPqybTYgUPvdTU3HYamj7rk+xma
nRbnlPk1WdqhMY2pRS7Jfy/iFnlKYk4cS4S8PKVkht2Gpt6NYOlhQyWuSw4dFhvy
BV6Tt37rmfHu4QJIYpposgWU8v0uPYwj3SgwGmlLrVl+5wGFocZ4IwIvZpJm/LI1
nZIi83s61g3PG9fW/o/23yW8zaKIXI58Y3Dcn8KLsPT6DV9nCY5Bg5jm02plvBCA
ub8W7e+/EzvLl9RWXTJGPoUXMiV40jgHStCio8jVdW3VhjlEGdeJIZDdYmAi1KX9
3NbUw8yrtlAmWV6yWUQzbuJdKQJEP16qJIWwIUvclpCnteBMzyHdj8l+5okMCgYX
KYJ5xh4h4owBcS4hLBo+CAHMq+2K+iNqiHDEtTasxjqAcXFAz+W8TUE+8lBYo+JT
g930ppRJ/OYOawG8E6YXEqAKRAGGIipaEZ+FPUavhvmZw5wRgRGv/roC6DbEK/ZE
6PyVnyXuD4mWY8iiYCjokeQZOq2q+gtMxVvG32mNOzmufBCQb5pEdOfDo9XUvq3c
rk7rF9HKX2kmpYbxqwqPszG/OYHtn2/IGpmkINYX/jcQ+Wc/0f+gnu6gj0Rk3VN2
VKddjdk+uDffaG570C8USoiU+JGUczZfm2IgsWa/cY+uUscL5tz4qJhnrLtNsQnm
OV4EV/22d8KVunX3EdfnVRvfEkCfR0zER4eXm9vicZ4=
`protect END_PROTECTED
