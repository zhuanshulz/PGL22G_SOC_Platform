`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mo0YWiS+PjHbp1K9Z4YVxSZvXgWC2PylHI+4X30A4+/X9/2aiHIVBBIY0vdC1g6Q
tSpYKTuBScA5ZlX/qPu4Hy6i+xCnZzq1P81r/kYUqcvMLSVV8yBhQpHY+vyntu0/
n2rJECg8lXptDBAiEIk0PZZ8vUGmVQXkbQChzHLU1f0hw9ZnjRR62BhHS4O2+Viu
QGNXs4F3bZGta2Zlk8jtEYzQdOjuvCzMOdVnijV4KfYqN10Slm/3N9NtMSQxO5ug
MdAA3yQZGnBLOrC6QqUCZ+zy1S+IIM9ZJ16ToW+MNCWUamX28W/ojfLJQKbzt9Up
N1qF+29vmfB9W9vkonV0jyNpTSOI9+MrPknJBqKwzXkoGWM0+ySBvqVjohp0Ks0Z
gqPiGRYmDZeAYH4WCohQnYAee1Dt5NR0f+UnLmPD8uMSlDOwOGmkjjzAYO2slSz4
C3nisUUH03Fg1tVPxwBpMZwWVz0doygscDi39bEjFUha0otwLniZwwys+ujycQ0I
WMYCzC3LpSVyFxhOAwpuNms0T7sAcYgfpGY/1ZHR5Q0lvvnKuv84Pj52rAwPyRuG
LLk4T/Yx8o7YoxGH46XyXWqCKKYHKGewcFVhSzA8L1TOroAekWVDY7okNoB2EXDb
Mq2IGJWj2YgleW+iTk4/aBRhnK3RFdtU6yPR1tXL2hsf8keXmzaHSswN+iHJn9Up
fSdNe4iP3CVw3aNos0I0XeSnb/Xww57Q9M2Vm1eUPUQmXuNr3xQrVxo5wYNO4tuI
iN7N0bzcdlvb6eBQA2TbTBsdPzHZU0IdcP9Xrd+qYCcpIGgXvW8cZsx+LxaHRcQk
82RqUiMKxG9CWzUm56FMX8NY2FJWRnB6VGX/GV8aiqHS1tVYlonVKyIq1D2hsc7w
hYVgoGfAcoaZfeU4izuYmW3eLr9IIR15512JWebEQCALiDy2cDe1LDcTX82w6ANh
YM1xQTryv2s03EdH+hsiwlLOvIi4lM5Fnq7VokC99SjUrSC6c7HToTz8advQrcFZ
67ZVcdYZwgdCP+OqQwlIAhqKuIaR8Z6DTCdSjMZQ1Ywz5KS033DlXE233puYptaS
fAYbZMrO7GE/cFd2twEdC7tlQn4pPneN7Egm0MrooFURu8eIkc8nVpPEi3+3hv84
KmP+30EC46t7KsDGyEoFyZU2lKwZxy5j1pqeBowpTnKhgl5Fc8zJBZYp2V22FpvL
/ML7E85KQBBQhCCBJfI8C3zZjp7XIqYBudbWd3dFLi7jd2Z+YjvnQH7ZJ1MHM9KP
uzU0oKsiBJzVrrzpdaydEVR2GKKu8PUvjnTCPrxYF0jKkit4wVMJU/8PPLhqRW15
9Q+bPf6TAZSgN75/nFm5usa0+ndS7iRJH6/5rSmxOkA=
`protect END_PROTECTED
