`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cp3flw6asOqDgvc+LPMyiUpRvi05NlO2wm7rZDrF8enlTLupd8l1/9f6WyRyy8/y
kXbAs6eoF21qKfI9U39xmM+cQN/98IXt3dqVf4fEFJvFJpG8ZMbdvYz3vJj5lFld
LFmZXW4zH26pTzSrc6uANgrba32btTRIirksiUUs3ENGVUSyqcCM1pR4bdYsGN0w
+xgauQFy9tE5xk/xPzxoKAqReufWIGWbMmHYE3AYIVtjR2KXPawimP7M6xRLuEze
KOa4heFKjoYWSoNux3sPtyJwSk61Hzg4wPbyzTETSYiQFzjy5LWTezmq9U8Mplhq
VggssIXU0gvFzmBAlH/OVi4dDxbD9umjVYe/fHDoepw+nb4f/bxlJjy8kkkMEP+p
VG9d8uKadSDEFfQRt8X4MqpHYfCh/xKNqaJisIWrK4gE2xrz4pqVhhjlF7iDG067
hTDo6IKBxQcIUID8WZmyEdFwxrKXUMAlO3vBNJyrQ5lTNvT0RlVZxQA9VNsf/7mJ
8n0jjHnIuu6aapYVKY57/AihuXGZeec6AQiPjFBrVYEZQOTPOr3NmULHbQ0INkVO
5nmJa2dmnQuGK0cZomh7ElE+cD4mogrZiQR+JReX4DNdya9EhFpPojYWp8or5Lmh
o9i5/k47OBMhkN3yeLMlT95IIBsYZaO1CoyvFxHB6ZbLRZn0BFcMVZGF/7EUbm/Z
TbbTBJFwp0BcbhWnQsOVBGbWZaQuDjHWnFO7iNGBjs+Sr85N9+y0JjpcqTBPIvjj
Zee94Ke9Fbb+b7R2TelYLEus4aYQERqdOhi2ssFv7GrenGwiFVz0AkIUZNyf3j/4
b90xXMPVygPFLh6f9Z4oj12QefymiU9r9tqUGGPwZafOO8Gp60j3iYQOSmTZN+ET
5qsXj/MxXl5QCFxg14to1aZLEtnBfMT8CkGi+G4J26qrqg1lQ9NIIR+bALfy2bh5
0ss3CEtvPKqDEOldSx1SQZmuUKiqtnK4mlWfEnsdXZs3JIqgwwR2MO/CYXoyuO7y
gPJemmd6rxxIdxM7mO8dvgUoMhYEUaKAkDYwwH2MFiPJWB5fn4TbESlCmzk6WbkZ
s0khH6/M4UubQTGbm0LUx13DmuH+USn6qOcSdPdUxB6WthIED3+TegCiKqnnUdw0
LSYvzEawKTN7UqwtdMcXQm6Sw6GsY2HZxyLKzNENBwCany5ehZo+p7Dqbpt3HJRX
YV52jfPTnlzrnRzH/fopyVr+eJ3P2zXiGotX6x55xFJk2eAOU2HPsUvwh83dicgx
ErQboglLBNNV6qS/37BPGj+L8kZ289f3nvTURg5apjie89mXLp15ZB8xwxOlbGlc
1lJa9r5WrVNCY3DFWJTaw7x8Awla2tq1B6+kGpT/sBYnrwvTvuTtvwa1pH6CLTPm
IyzfT7sZVLogWaEKCHC3hs0uRNKIhLClP5qRnrF63U3kviY0UywuKm7kywlXGPK1
MhEUeDqwwMeQUnE5jDjzTJumILuGJSG59vZdx4bPKzPkjErKTSqkYuEuGYnj0dMr
H+83ZRxOaA4QtmszQElD9YOVJBWHTi21TXAL6RuHs1AUPKwgxCdvZCTBm0U/PHE1
xR9fRFVEkokyQjKO1U2HJ56+2pwymPwEDlWrO+ZtsSu4RmRuq+Bs7tQewCv1LoY4
s/1bdm8lwp8Zk1fGS88w81wNOR9tF7sTn/SeuMLQYhQXyifzeWYNVIA8+aoN1Oq1
3bhh0vsx4VwHoB79cjR57czR3ZFux49TWkzmRCAppWny4G7/dD4GUNXITHCUYkxi
vJZbY4NU/2KvVIPEc7IlYkjYZaqVEpMBTPUKFOpcK/uVxSo97SU89j+VuyHHb9OB
FTNH//+y8DEWcljE5SPvZB0c7IMU6FeFkzQHSyptVXzeQkC+Px4ZD8KsApTPr32V
sXqXI1sFPgeE2+/aCFyQ1EJ2c34cMvNM6NzEs2z43HsuEtimszetVpTe4TMNBmja
4P2A+OCr+00O7I7wOwOdtJvZM1RbK7IpPj7fZCGxT1EgnCU8RrCIEL/OkLuKpozm
Y+DhkDctO/3iCTwMQTTv+SzJw0PKRi5u78Q3DbesaDLOfXQChkIErtxqaXrkQzUj
TNXTWDpUQ4LlMn7i9yClmZ0JSHl6+/HeSRTN/fiR2u1pZIveIeiL+EAqpZtmD5NU
oh9sv7Ffzil6lK9xUCYagZMrNQgiwbkcNgwp1wLe2kDLA/g2/xYVoqVf5jsuZFc6
rvpydqdnt4IRCfG98zLzSeVGsaLiKO56UHu5RPNJePQOfVGigZYkanRtsrDAKaa/
REaa903wikRnF9JmLsMgV7BpTxRnteUSGX6rT+NR6disIHQp6uxDYqlIPKGwN1zH
3wZLmyMkIAMtqsDwpsHzdW1UstiTgKRrQlZak15OfvDvcy9bOEIpUL+oTeDWQodI
4B0Vc6gcy8EnTeg19djoLnj4SvDaRLgsaNhwPYyzEZ0ASjwH4k++meejlHCLTdO+
0MXWHwF0a4UqQraLNdT6Y9WWaRKqf22jvbaQ7IGIEilcEjtRN1nD+86PhNPV88jS
/RR9KNnVGiEALihsCTWtvGQiQVl1u9b+n/dbI/3phIenjVUq/nr0C3ZyJIqoMCNv
mOcd06zxTBX8RA9yM6INv0jhghsahBQtAbcRz8UVnCgDtIC+irMai8H6v2ozC1NX
gPKdnrPZ8TZwfq50LRPb0xJBOXwCnQqamEQ6vsuRUe3F+2AWW5E7WawCY8NdPJ4J
XjPuI9pipwbUoQUze6yM/qpl4gyembESvjHC6zNse3PGWzmj/6NkKyovxaM0rNnp
MvTaTxaxKecZUOw0lNieK+xb+lzkvpXZEBzjrLvgXiYTt5TMGeYR+QPBHcFRCsKm
4zp4t2PLfNbQnfuYQTMxbESJuYqVkuzkLAcn0NokrXKzNkJJzCHc9Kp2tEjINe8M
10w1hRqg9CGQE+0e6bgNU/1wZuTWbz7ONFF3sMAg54nGhiU2s1XShkThTUFBwFgX
8YBHFB/nEp/miBoBxabl3cvHWb8oouFdWEoOULEyMsyPjZGU6E+kGm0LD+OXrNR/
VIt31hpfEjuzWKFSxizxIYfN7lhDFAXWdh/08N+2R+JqrVyIY8qh2TBhGbeVnMdY
ot+xH5jUqrf3ycT99iAsKXdQ9IcO4YCu0507rnTzvywUDxp4pGiPhjYwsN3yrvxJ
p5I9mY9HjClXLEisvPA9gl74HS2v/b7cuHjMYvBmkGyZnr1B48NTZBeQb3UyRKY1
IOCOFMTFLFR3mTCx8ehkgS5aNA3txKgnKs3ml8cSlyzzWNIqjGbyFK5d9n4nUf3O
m3XRTr+JQir4UEiz8R/aKHVFcSib//LOBo+CoZ6giBkntgEwh4HtLvcJkBFXIgRk
29rZDxYN4SLiBIaf0GjtrY9O46f/9kit6g/asujEoqVAD38BjdnwIZK7Mo39G3c8
Q+SugB71fkZiIZMzfyTHkFWWidpqKHNXW2o4GbfwLmUDUobRS4vwYl5+Fr7KcpXu
yd7StgAYag4ZiOOy8mJl0mCxYaVglfRHMY58/r6N2fTk2zNZPLZT0yL82By3bWdG
jo+c0M5xM6QEwQ5DwFQUVoUf+D7X+gw8N1DNu6HYowmTbJAYa1khsgynRvZ6dVb8
LEqCO1W3M6lchi4vT0Zau56wEVJC25zebAeRqoIK4WRv6cfWFIChzEV3jVyIuN0J
EWwWvOSkTFf+WzXpUA8R/ae4ekdovpqTCLi1BuB1DMB6AnB2jypCn/I+5GHMA5Bb
FmA0ayIbCm1Y1Tlk07Zwd8O1A0G6qXJtLT4/gmB78z+NqCoRPtfpophV1AFqdq9K
AImVgR6zur+1oqks7i+PXUAjzjwmaa2WTOomtSwmEIX6aardIYQCb6LO82cf4fNk
zJqQK6nLt/NyE2pelnqMuFiHGf9M6iQyQI9T4nUY1sOiTvwOzpVfn+B2T4i5EWAk
MAFLA+dqGTBXtq0LPz5/czA9ukCEhEc0ROPU/s4x5JHsOzPEV6KnAjbImKqYpv/a
Omjjpmm5pMu1adYCD+jmdtK/sozjIn0fovbWd6wtYVrMOykSZ3tVqp73kHzSk6+9
IB9c9O9L36UGxQOkS6MzrfdbYYEjmhv2tgURnSVpksmRsSFR8EJKXdum8zD6OgsE
7YBJyfXhFWnjzlAwD9qewpmZ6rP29Pdk7PVtR9DBuDbF8HfZqt39aPtKxIN7DDrs
WDRMxti2VO/BHgQ2fC2BAgZX/CoUCEs6k+9koU/GZeV6hdSt4BJ0hsY96DGOQQRT
zFEojl/BFDfsKKibzaarrvYVK/hQT7uMTkuJ0zaS+FTCtNokfiw+9EFe3JLbZ5BD
M5axB8xEeTioP8H4IYD+qs+pnnaQNLN2xi39EM52shJP2V1lYOx5XWGGs/Sbij7j
yLafRlOwaMYpeHkGWL+eO6MY30qvsFbb4WnaEIAcQtHemXgYZ5WuAyGmOZq8XYgN
xx8BuYPqj+EO/dXDg8ELBZP0O7O0TDx9GQ6e8hka0q7W2RofnaLfjgMz+KM31Q8g
UP2XTSEIM1fYDCddV94qlq8tRCYXRH40CM5rcZ19SM1P9g720gUFnXrpxSlTdfjG
mzu4IiY56kLXCkl/p5qSQacVXOrceKCPsUByyObRo/wd/b9KgGeEQG6wWkb6TtwQ
lLEEGVf6bqk7dXvvvo/ptIC8nUEqvW/iumtp9gnlUG/fhsbYaquplFP6PeWnsGfG
ZAI4uHjtxCXktOYaLWh/MOvZjbVXPmqg09uD7oa5VXya14T8gwJCUjS14PKV6lW1
V7/RpTdt9l7uyiPyars5cUwIqB6h62jvXdTMUR5xwDKArQW/L+1Tq32D3TAMcHsW
bxXS9Kw5ziM6dSRPlgOReASnIe17B3FTYqO7m7m1oG5RO/SCLs8mrmjm1uea6BnX
1D+VnjlXH/qopsyAGIdAACD35UoMP33G2yRZA5mKGmb3BhVl/spzAeLV/8FgisJY
yzOZt7U//mCmAUMVH5mSQnGi2oI7COPuOuTYkEYn1Zjgj+YAd4Nd37iOMzXWmWk+
2G8QzYcI9QhZj/XeNL4UFg3t4eMuwYQfywBWgC/7dncYoCblcAHJ7kg75yXER+Rq
LM1JUXCPVGfUjIhkbc48hGNGV5a/aE0OYzawPmRPv3YHlIC+1a2WEAaC9PZA3smp
C7b2XK4VteWQ8WNGLkF5ntyk3aOFh2ZgURCic7joCKvHrDSJ1gkv08vx3EyeOXtw
tCNgFtg7hvgBBu+X19cQl0c0rXXCxBdpB9/0j5zNMOYcIEDfziB+zO7txThP+/D5
yW0MLHQ2WKJs7smEFsHxyu85t3rFmXasuDwxFH4gctWRbKxanlI+wU53Md4pDsP/
Y/BfC3+fiht761IGPG2mBj2CuQlT1RkjdapAgb2z+2khxtKsApp4PmKfdDmRuyVM
ldLmzH41ScJmgTTQ5idqLoM0IL+TLyJncZqk8mIqG6CnjTjnCKgtZKArzAfQaS3F
0dWf8MgtMaevVffYJa3HEz8qvWtOxSP0rfz6+FLUow1YH0Pi28Cp+uI8Vb5uXj38
XVVnKpyC2bCxigvZ1iFBXEQKJYb1/4BI7a6yqtTyDtHt3KYvpswR+NmGukocnm2U
z16rZPzTGcSaiLAe91VB4BDEvbhRnxXcHH81021oCyQfuvTwNu7YToSkuu7zU11H
hHCZ9Hzt0zIc3s9faUX5vv5NcZZNhAi64dpPp7LWRR2ZgzYFOyqEq91yRhMojIA5
zw8YMv4lO020wk1dJse3JmwD2VeokzcihgfLLUpitSiO+4kkFc8PtPpSW2zmFZBH
MHEzI6awBQ9aBq9bCqHCiH+dVSpbSKiXPjdLq6tXvbHWVFVGd2Rgks24Z+1ymtsy
m7UnWsnqJQ3bMN+VzmouTNOHCZCrX98/cAa4NmR71v5C83AAO0jIUjZLw6NoHLDI
dI2dLXB4qijT9d0j4NJRcNDg3xdeZhbV8JuNjjeD8KKIWqugzHxHQCRkBUfbuwz/
k2LMWwUU/UkSiRt1hEQGb6BfCpna6CyETThyLOgIP6b43sy0yGoWYlZFyhnBEOUX
MF2mpfx5s7GfYZ2kMQueLVpD+Qv7WigWrEXJgTGScbqyGiDqHAkW1kmC0riZUhMo
CuD200doKiP6xAIhcn27WB6q0hQyZf78W91CjJMo1nxb6513j6jOCsmhrtarDMcy
D4VtttZtzNYdbXdzEXrr1Nqn6CF921mXPuV86FxuWdzSbN1vFtcONOy9+YbHpgRw
DFF8lbm5/4mgYURgsr0Pw0lNJGVbm3BjCNJj4poOMJ8zidAKjmLu9gQT8Fae6N3a
zaBgT6EQ7CE985K1l/lz9+wN7Q+txScr8k4+6DFaS5C9jksgvHOUJti37iBQX1Mt
BD9wtmeu2rmsPEZ/jwBLKSGYOTvDHcfLAZxMSfZb/F7epFIxpq14sVOGu07VotPf
ckpoeWrjzi1F7t0GTcQrjEXyBB0SCg7d3me88PJ9OZx6TQgw7arL2x7ZJHdje8np
IyLjLn/bYvnbnYXNfTB8gxAYFJmMWHa0pL/DgaP778okocIRx8UhUBEIhbWnzf4E
DZR9gURICSGogM/BPlp61sBRlOluTH645TotEotQwp+CqL4MXfLibIbzS+bk6ANu
MWn8tJ+9dMbIADHEJSr+7oPEF+fkT8pA+NIJilx3QfII9zrT4k9bVsT1dPKLgudi
FoxPhpck64YJD+T5ThWyz/u58D8R133XUZWendBFN2M9NNaDQ8SwsEowj5H+EO0Q
e9jilfWbmghrkR2MYGn5GQ/t6JFRWk2YLgvlpHhnk7IJs8XYuTtwNgenJ+//qx23
0YSjrqczGR9FMUXT0oTOqRwaLjRmkYua0srF5IQUkIPyNemsU3Dv56xRSEu9LGvL
5dq53LstaUxGIbga0bxMq7O3o8fMemo2/xonAwJVDl86rg3rpDNxHLqd2eJdbsZG
pTZN4GGbby1oXbfzb2JxnJ3Yu6u24ByaCjbsUKcjK3PVXng3+wrva9FJ06bYx2ke
V/32ww1Hx8NW/V6dbZJxHkUi+awsGj4+dMmRHfGtdIvY3KZb+5aojDfjqHq/NhRJ
ozqJuYc6r7xEUmJR1NlN0PHNx1OLvGlnFQggXOuu27J3gTgs1Viq4erA6Q4xbqTl
5cW8EZ6Eq6a43watMOmNpcgK3XOKV5V4FiZPsozF4rNse9f9otID1X/qeCdsn1YQ
BDxQqt3/HPoHbo5tuVklnkzkE6ZW3SE2gJmFywUlzF0RPTkW3icLCNRuEVVxS20r
yeQRzZ1u1t3LYw5eqjWyuFnIVVlI4r1Dnu5sv8i28DIbCelDQW+kk1o1TqC9X9gq
YcEzUCCJBmqXnOPQgg7TZDpPxcLPSXjfn/Qu4MoCgz40p+uHY8yEvYZ+DtBUqjSi
qdTPxEH1s6enqsiwC7JYpcr63M7zSRoMXtJw5I+avkqZj/MTj594ronQGen+4mRu
N+U6TsVmM2zKQM7hj9KK9fPVN9oJ+6OjQgh7/xGC7v4WzhrN4jpY69IIg5+eZ+N9
PjJW+YzL8ZJ2bAzaH4p2KsPxySxYsMa/ZnQYQbiUKdcGMmZrE9DG1cFsdMXtEmy2
5Zqgk9IHMSSfEaTvZ/rrVdYD/fp8L07EYHZLytzIcSNKeTBGUa9pK8PkcltVG6rW
Tciv6gMeLpoRK/K69KbSzJvcRcoTXhhGSHFJYtpADPOU5NIzNlBHs8BoarBk51eh
vtePKbKWOSc8GEm7z9P+BGn3x2qy1egJD4xC0pDQcUzow7w0xs1bwds+o15CLes1
OR6jw7si4VIUgGXlKwmH+ftFcFdtIp/nQ+Ma8Ih9oGYjxSxPWAAAFIXs10NxOFAF
dl6lghjKsUKzk7z/rnBd9fU5ZlsA1jNDImDCkP7oV8SEBmz6yRbwC2tXjc1wjxW/
hjcHnJVg9jbJif0g1Y11jSf+GFv32DJUuvwPKUV2DnN9CwlOH28VOmbZXKl/bFKg
/bRZrZUF0VHLvoyDJhOjtOq1Nd28WoCeqhkIK+h5BF7oI4gC8gC2cFOKpTYG31tz
S/Xu9dsOzSodr1y8r7jVIB7MNCq3G8TBjhfjXIwhjcRPmyyl8593sFPlMOVaMfZd
rdftFcgIFz1kq0ukwkna3UAkIWpBXNsE8AkKoDk24D1LIf9nreS6Le5maQBO2nXI
Y1rlmBbaFFMDr8BqQpbm/LET1XWeZa1Zfpo7sEdNXkI=
`protect END_PROTECTED
