`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/Cv9rUYTDPvURpYG8Cv8CNkudly07MctvhhJwQufY26kt9HrloXzrCJxPH4xxoS5
aa1bMkEDfUrzSWDjSj0hfGFBod6DAVqCAHEOGG76rW42Y68UEU7MQFkWKXEIXB9M
xYkOmOhsqW9Bs/DlR1fbQE0mrC650NpCCacMOEDFoHh9N70MpVMeb9rsdQl8LCII
97XjYyRw/SeFlJhxUWvUB5N/VqsT8k5j6dCc0NqY4a9yVYS2ekf0a22/euE6yyGV
EBG0XRxl4moM86VnGB/4xwpjguDuUACXiYtqd3vB7sjNoBpZiO9x1AjkYs+YF+x6
EHsPmCdvoS+4mIj9hQuD7GaJrOcQXiE/4oZA+ZQK3+lC5M3EjuryBUQ2Ya+TFZ5F
aTS78jU/dfEqw2tBgKGCww==
`protect END_PROTECTED
