`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1tGoFsq7Hq+kHLSOJCgekpols4V3TpVzT1HNkpiqrSHBhNT/rcmCoISjSro2pbEG
GcmYDWpaVx4P0O8p8rIiqTflL+QNMnOqshTLSskXJPrRYjhX9YSXO/CzYISHcF3Q
gYXLWGZehXgIG/Exu3nbfhkCyISOzizC2asA4bZXEu2d/gWHli2rRLkcnAQh4dl8
/tI3Pt230dp47cTCOLz/AqtLsyRGTOIczZmqu1ggHWafTkVnjvU57Ae3cY4D03nk
yk8D3EaeRIYvJwWexyo0t+f+wAw0rsBOjU1zKurQ/z8oDWLv2oWW5tnpLf4W9brp
iNsBZt+GBqjTqxkG71UGPgHp93Z6QUMSNjXbu/0cl4sSl73+vJlQG87eC0Nh/RZN
RS5IDBjHctfWvGk1rg8uFAQBy5jAMyB3VMkJghYzTO64xLD0xjhgN+TXWugeiwsX
TEaYQf8sMQSlfQY6ZaiwimLUVsT1H5gkjp5fsiqzV1YCYRJATII/b97eqWbitMlv
DmjnVDeYvasWx2tJKm2iR1W7fhVUVkUMuWh9g7Q3bxAp+Az/4Ch/YCbhZOqlLtoI
pcXxnjy0HWEIy8heHm3Ir71PGwVq1naryMPwv8GnCNQB5MEjXuxNDKSPofDWdjjO
rTXwFtMTU12LQy7mMgOB+z0+FNS7UY093FrVUg/lzL/n341OZcApEPBJ0DCmGS33
py7Ns5bBs+aLOcYO1MrJ8mpCANLfyfkaENz+cYVkI4xNkqLeWUaPnKVqGUrPqfI3
TQfb+qgTUPVOlVJCcuniZw==
`protect END_PROTECTED
