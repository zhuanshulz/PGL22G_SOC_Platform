`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PjdW1XZ/O2Ibq08TzaEb/biMM9mM7S1mnSfgIqgm9vvL/yUjwzbHRfY62Rv/cnRU
h4Iro/suAwkEmyEkD/woVbVDz62XzKE+hCT5oVmC3uf9w72ArPWc7QzjlLqremGE
A6F0/jHfrYhZ9VvmqkF/3DciXKR7QMZnobv4NgIJRqPrJYbe6WCg3htpp3xGUVZC
3X+OuUcDxII4BKNqvYlUy6hn7pbGnODkpd8bPCaoEtCJ/wqoUU8i+D22jHmiZ89X
diiSZ9WKAIQWC67Qodn/44kqugsh/1tcDgNr8oSrw5DxLHslgji/kcKIRSK/f/iD
qmmE/VpS41RpwQHfCon+fSdxXYd+Q6aqa4GrNz31dLqUzQtxJ1blS7hQgyUjfPvr
fMIhy9PiQ8NsWz2O3O9l+VmbyFqkY85sQDT384gyfJCATvkcFoDoY3uIAIs1sSqV
pUmhQ4gHELC/u1EUND/u2dhfLsAD+g7nhFXZAD2Wmci02osjbA+pT/yj4ctnqRzV
AuhTqNCBr6PM5a1AzDE4olaIhAoZCc16rW3+4LCMM0OzuF7LhpQ4iM9vpRe70LYw
RBg8WwqP8fLavt741++P8DSoevCmmBQh/sddkECGlzNFQtXpajQjqvGD1HMRVDyl
xACBr6Mid7iC4B/e7ssyBbcXLTAxQnF7x8+eev1qnwZhoKA5+/XOgJLF91tO0+fz
KRxYqQpTPEDbKkKFguuld7QHrsliHtXophv/QQcxeEs/5b521TjWh2dt0RP0Ihdq
7eyhFMzVokd+xyaOe3I1+IWt+ZGOGLCXlCd6NuB4SKqDBR1sygsy9fgz2UQZuPVZ
Q8WzFy/E1hrTb/EZGL8dxswednS17XlZTsU6TPly+5R1jbzVaghQ/vBswQjn11sA
OMM4ELG0dcoMLqj+T8NVTDVrX02Aks7yll1pqjGYfEzUSz5HOlSF7woIbMMe2H90
uDlp/sFBKKLWNTOwtFjK3INnioU0cRe6lYqx8G3b4Z1t++NMk1ioO0lbl7/P26dJ
A+E4cR2N7pGuj0RXZlApe2VI/pj1Fd2wS1g3ugOkDXg8egEtwxTO50JK22ao2ojs
CLNvQlLwDZ19FgAUgTFhg/sWx2+IJZW4YbM3/ZHRTERNAR5cXqqv89TYgUIu2F7l
g3OsRnWSy+Uvkkzh8C17LEzu/bqT7rF0/gABPxJiQX58lo5+n2myOH3DmtjUykHk
lzccYLB3xfc8oAxzFaPHYu9rWFc0HF9h+ZIXNTBaebbL+/gEs1xi1QEDC9RFc5BJ
dwNLkBxcuLNcU+uF6NOjajJZWg+dgOabJIo+xZmccwR37rETL7RqMzsH+/2oC28j
cRkQnbterA6Ibi3rZ7rTfI4qAUZdMiINzDRns/HvPKL/aDju+S1qpXPHuJdUp+TI
hS5XmokqBGIu+xvLvIa5m4Ggs2oOWjofbTnwTnJt3PLh/T6tpwCtvCY5Z7WpV7Kq
MQPMwIM4OmIqTJWLXpa6HYejEuZbYm4EE9gvvVQVEOue14HbwnYTbFfDz7CG8YaU
0Lh01Aq/23RHSk57NS7RmrdbE4+XFGgqF5AoMVlueOJUmvtLEyJRQyEm3XcoEUDW
gX32pmF0MHtYYhtja4k1BpFdtNn1OpbPTK/wigoupkC6EMnds9XkkmqzPXmUZZLx
P4/l+u/EYAWisXk3V4MpmK+vvNnvSsKlFua0XtG7h6S3aPsQpBtF+NSEVBZFF055
HDFKJN+M5oMWHCPoZwipdLHTc6S7uHYe7PEhOw/3q3cYliQFVb/9lMnLfrnN8d3a
m5qJlSPY6HL7EOP+V+3KZtEgrIUJ+85LA5JpjeQEuJ2UgsTtYQt6pIPa0KLZw93q
Xtrhx7OzSDLzwK3oNhnr0ueyKfr0xny8jDzMjba+dcj2sBRSHrMqv16dvI7hCMGD
ghZ8chr7n2bG07J9gYEnxaKg3OyJOORLgl/XUN9Z5VjsUr0Kc1JdZbtGs0inM6w8
d0Nk8FXq6nkkUYq4B14hariqLaT+cLD61/fpySDwehryd+ADniQ0WPvrdMSQEfhi
fNh7UJLN8TPXgpFNbk0nWeyfh7qHYv+rHclywxHyhD3pv73+M/t/eFPWoCKIFIiW
OQiXdIV4Npg9P5fqv+kp9yY0gMw0UZvOLn6lTbX/27TiVPQ0CBBEVRCYqmO+G3a6
yleOaZew5kZlHvL/qrjrUlaCJiIEUJYllIopRZV7+5MCs6Z30CeQAlhaID1pKc9E
cyzBoYdNgUdC5wEaeep7mM1eUnoEdbpfsMVRscrmXtmuvJks7GR1LxrDLYSraGPX
lmSJt3q0mfM/vma0MeI0Q5gwAcVVPfxMKvUDWGRvYyWTf9eYiCs8ECS6cfjAHFzu
xt75iBoJkYjqj347zzNLHYBEok3dyG477sKLgpjv1ReBC3lj3DmA/3P2RmPEvxfO
xb3iNfB1M0jy+YOgmWnMgD6Ter345ZR/+sHOhWMGXKwSSL/8e2bGaTS10Sp4H5qX
8LOijDUe9MS4dhfdYaeLbByfXKcanon+fMf1x6V304K+BxA1eKAgPYrE15jFtxX2
S6haQiYNGQvm4iwxWfAIEqS6jLP/S7fVf45YM4IJVvjppu+DkjQYCTbyqw8/j1je
/nUzarcN7ltt2pHhAGigQhJbT7d2yrTn8pFwBkicGh/bqWz/0ryvP20Jyze/p8jF
UEpqmjTiYSHY2KLN+kVrhBPSfGhXgvm+qUVYyHVyb90BUBt26UEIPGMRI8QSpfmQ
xLQVuMEEO6JUzkNAGTDaWJjYLLI7HUWHklMVraNjm9sts8S79Zz6gm04xlRLcYph
dmTJuycgx91GQGnzWjfcOhQaYw+Gq+Q3ojMHTdLS8WtR8cHKELviNAaQSmDQ77Kv
+NSzUuwTfjKnEE5M7cOQ2gymlVZVlDe1JdtA5/vQhdmlZK/1wW3x3tJ+8yhd2jbx
xESxriT4RJi0ujRvItd5UUEcCABkVhiURFWARFqe1dXT4NpKqBu3z+7kR6XV4DzT
m0lHA5RF0FENNLkEFU3y9bwkjyUhKbBPSpn2dzdo2kpvDxvbLBw/7zBV6TQpUh4J
R4fofLi2TNjiTPckcFHQPamRSCW5R+1W6T7xjKz31/z/+jKAdViJ3eVE7BrvJgsb
vfySQxSIxN4rGh2hAaeQIt6LnlT/ELD7sasbuMhQnDq6KbP3RrDNw0J3j0TOgpRl
9dKNlnJg/j1GZRnXMuuAbH5sVql1PMcZKP5KtXbAS6Rn+nUrAUDq+EPIYsH+iYGG
TGWixl0KAYwaKUx9unlfhjiUz7LefSaU9Rf8dtl8EkJ0qtM+F7VdtFgWOusfZ0fY
CcA9cFwItLdqX6JaRbgmNW5sFVA8XqFPOL/yiHK30a1BpocOeGjvj/09VQOCrfzu
cjazFJBL1KmCiUSjHzo/1zUiOjyCDfOhQKZV49fr2MwiAOQhHh7LnKaJBDYOChij
PnuCd5PJxE4jzxNjvsJSXEsNu1Qul1J2qVq2uj+xau3CEWsY8uUgu8SzaRojVD1y
9JzpohW04z/eyFVs+7vrAtzUb5Vwyg931DRXCOkJaLGXQbdMrBl974H/AuX0nehi
20KEoobUFEobdte9jEbNRRmQ9AfKod2mZTlJnpFNRCp68TpUfbUIK92v8vIc9J+t
Wz1uC1HiHSB341TMWhxGUwkTlPNjcv/NCMlEVPKYle0ZmQiYuAUbHBfzPEQUvqNr
ueGUPeCeeJxQwcF2zJRcLK10xBnCp2q8zooA5xOpB2haRt5TIAOkw/iVRZGS/isk
grI7cj+WUP7s45G93I5hWGKOglzN/WRLSRk2z8ZlwL3WK0UfwnEOt/+rEaggIPCk
0A74HghWjdTWCsbJKgNA7Pyu42BI6zLZtubx6CFUg3gu0SBhIPmqocKXANRv5nki
oDH6Wt9KEntfCwevNrmn9l2Ycrg/RGh0abOIVZ5ZuS4q+h1TakmftlI4zZL6k4Eu
eu6t9P7urbI9vRrREhcE1oTA2sI3b+QWJqMDAhBS40rsX6bfT046DvVjJuF14cXw
U8yJljUr9JfBP+BI40kVzs7nsJGun9XObLd6p/qE6zQzzIc7oSNp3tLOI9Z9TvvS
0W5AK0JHu/qFap0o892vY4PEf3gNGpH24MXUMnd1oos9cmUwPGHRJLxFTe7V2R07
5XLIIyF9wWdgPFAP05JaU2VCR0E6B/nrYnWOdJlmcdjLXzNNNcvODOiPomJlJCCt
tcW+sAfNH6CAZdy8/gPskAuVMK9uRvxA3TTlYE3/CjDP36Ohappp9TJtm+1nFL67
lbGyaC7QoXRYerZPYfDf/FieviuYxLlEpBCjHy/a2BdXevOrSLffjiyNWN+OJn6x
JXMdUvhELjiq4iZXqWDu7KTgY3Jn3k2iADU7n73WY2OoldnJrCKRRGJYAen/zvTq
OlcTmMu+2zJUQxQvkfwZxdfTRIxmrgGZSFiZEMr9AA6U/O8ypL3nFpZw2/7PAmfs
FqmJg+Y+NnUIPYfOridDPMS8klSmYIFWknB8glz+wW8i6O6i5g3bcRIOFasJ6RZ2
i6ihPTgQBA7gcHtpTEPARC/fYPSJWQfHBtxhzUXYgI034wPvf4yIln7rWvm0ts5y
n/lBFT2WYtY6GRN963b5ZLlgNbPE65NyqtSMKQHJgasCsP5Ew35N79YAjyW9ruTr
MFccIZUhOWYiSn0R56W4VkmTTTwL8T5nSt6ZPXKluajicQ+x1dIx3SJTRjc8wvkt
nCjTDWW42xjulmB6osZa96dlPmqU9JXz/8juyCmXpuBxjZ23lSdY/MH3JAilGP48
Tuf9XNc/p4izf9ya2+9pf0B4GLgyjb0FcKy+ebSJ9gBFR7epgJASXpNBMJ/qQNWf
VNto0Cr5elsu8+/6SRrPVURqufWOprSfPFxbGHEHqFZHaVwWwGovV+tfYEIoJQO4
ndiXoi2u8kPtJWh9M3TlnOJvIZ+fxGpPeWaQ/o9momOPj3JOu5zp4rPRXuFv35I3
ZxqEruJONYFAa5H/eOilpCZDVagGTlHclY5i8m9hHp0qhQeRrpN3bzQKe1DYB6J9
mS3zTtAg/noAHMlTNYSxJa2pn5uSYUYxxrGyFDlPwwA8KYMxnFiPSNnYaGiTti6d
3mutVvDkMXspBNpCZ05i/AdCPsbw39J+2JwaX46f1Eom+f/nzbeKo2LDei93cGOE
yncRkfSVmV/PGIsuEAG+H5lnZUWMsQreDuEKd6XNz+5DcEH7Ks1GvpTiUdKG/OWC
cgqfNAug4md5eTPDVbBvn9Q00XMpAe3lMxRQoiQTbFullyCkwbYaHctt5rqHQyzg
xjcTvCMJWGqGi+EGgNuMyL/wnoNz5WKmuZ7SWc9SbuybxtwBV5T8ZDneYDgdZgnO
LOYWu80P/6CYu5GGIc0w0n1a2z/h22KyIjU6SEXR+EG6IOo0ZcU9KxOWO9EGkBDc
59UGSMQlrJ0Ipkvi4Gsca2uIgsrWWE7F0ll/NhaXYgYAqziOZqD5KDUd8W0XLqEe
r92FLGjpyQsuDgh1cIYhkgoc0aHAF0yVOkaOSCGBPxIrnfNcheWi+Ygmxv1B0+bD
Uooz8K7M7AAbuWzHd5bkHs+Ut/o9lVmoFBQ0vIZf6PjgDvO5ex3OoxlcQ96W9cT+
Hx2laqblm4uz9Hv6Aa4HwAJUF/yjzygzP4Yp19e50EcA1XAx/jrQ37VqVHqUbkp+
GjFqLee8E2pX0YQT1H7JQUdqVDsQznJQTGswj/qCHGsxcxPpAX+ZVQE5KKzMxU03
T6vDiN7BT90W7t92KDCWEIAskZyZTLqQH1+S783e3sZ4qXqF0fUAhe7QxDnpeFYo
94DhSAZHQMLcEDbGjZ1tUx9KsXXkarrRXkt7oJgSXoIMfNxjENp9R8tm8HDbIsjO
kalqXcDHT/rV2Li+NFTuQ90hDfudTT2vLOS0GVYXYBdRl8iOgrVDTD4Jf/5aL6+W
aUvGErPciGtCQkljd7ao9xvc6aIz039RdcEds7RLXny0hPRCck9KpEwJ9prCgFS6
5sHLhgcYqr1WC2UQGaFraKVj6vQcanssBLb7xfaQcwT24ehUs93axm87f5IHlEwZ
tmXLxcN7zXwN4z3PmYFW5p/3RbTfeKcoSA+V8StOi3qXyPihS2L09NTEUMh82OIB
ZKfVpH5igU6ji10u+kIuboEMeii2Eear648rD7aTzuSGL7vY1SG/QH+jCrTktKlA
QNRgcB3dCqAhUdWwsNzpuN3YpuVYBuOXtTAcJ9z1Hq5e8vX+IXqNxOkh+aXy1qvt
Qyqy+mWvgNPpWinGW0C4wsZ6r3B8moTosIowpJYms1MTmO99bZVwZMN2cpaBDjoR
pbumOhbumCJzHJv1a+yYOPGJFnLsxB1vt3HcgJzj+d4/PEwpKucLwwmbgZpLVITG
Z6PK7BptvP+c/dmR3tsDGTLtRvbd4rQYUPvqpjX8BP/R0XhAP3BJU2k734IjAj5t
qPBpk2AKVutn1Rk4qNfe+JXZLKfJC0wlZmdtnwgiixsLKB3UJ/B4ECUHdeXPlPrh
KrND76ZYDvA+ZEEdTGNZJiE5+xla4GZgejbU7UyNujUPMnLHZi70qj4xVW0+cK+C
7jvhrfB4KmMP21+LnNR+UYdZJH9HqX3wEyScPyZnVkY4NmYqqvKoljKvIKpKrehk
vIqpBs7kVJbQQn1afbiLwbz7KBBH8eZsV3Rg27sr2xQ2/WTFTVkJs4HJ5mF1UZ3n
jl5sDEmDViM2CTBaBlpzzNDK4L1/eCp42j94t3+vq1LepswnOYnSpwPC8Cy+eIjQ
ySAsmsWEyMjh+KLbGINJlAzEGXMPSx4rg2ngZPmQGgqNvUeZGMglFS1Clhaaqv16
BeiIIqE+8EeYxeRJAEML0CKZQpw21c5+VKaT27YYxgm8Le4HlBCIapLcZBHORsbr
bpgdkx+yGrho/OA0SQgHXygHN3XLE/AxDVUX1QrGRHgvipCvUq+ZmHeZenG+furJ
inqkaY20LyJHvORc2hCfITydmXJv5dmXszXw4KnvcfD2Oc0v1kmhl6rcw64IENx4
JZ5onZjrMUxrICD9ZUO+gRABP4www3XGD83QvNhsvikahLb/a/NIHBdHpxarQp1P
R4seB5Dikmv+Q38I6Er0qUn7TtG1yRZxl0kshdfbTpMTyPQUQZJSmstVtdKzJiUc
tk50ZHpyD3HV/6m50pOc6xcRlkVJhL8MEjCg7m1vtykijG01jU1oCdTx21YMuqGt
JkJoblKnG5YmnqafuNh7OPFToPMy+GdYl8xKIY+Le8M9PNyjylHe6OfSj1I44MQk
8nmqRSglrD74pGY1zd8zdqrX63m8Go+By4frmyYIjNPY89IYOoLvz0owN3yS+Leq
woAAqukodcaWR1+t+vESwuMhJGhifxLYa9mkDc0DgOmPEFuwTdLktCk9UAyBBXnd
t8aXkaSiTc99FKuZ7XOoE+j2mpppQxNwvD6xI9uAq+myWaHzlWERp21lRxQ9u6ls
R3wY/k4AUDDvB//HyltdZJw77BWHhfU7CPQGKXaAc9hQCsrUOfhMK/SWsYLgTQua
CXyJo1FDUMrjaeNsMmGuPkOPwA5i5a+Y0Dy+BJsIBWImtSq+RvcV7+DPJmxyGjkc
MlT4NUxHzMhUPjMcFYS++1KwMdBVvM0AGyVlGb4NtGVOZOzhR1vLxt1eEIhdqhiP
hopanz6Sa+gc4HrwCdt3orpSi6P1T5D9GpU0gLMeaQohAoghkjoj+BEQqNqPUFfr
y0r+ZtDInyHZcouCJCb44H0iqG3R4j3Ait/Au1apsPZlF7rwQBQlTt/3g/OHuy11
1s1OGNVB+Pp/KsL0gSVH2RmQ7WYuZHJU2bVNSGCDdfmyWKdeK6vCTxhwKXx/R8ft
/4xhLRY+unQsu5c4xhvBa/7HqRjybKn9tgYR+nEaHoEDhxNghXpVAxIK61SMr9LI
hpndFDrnHeFAb7puEjGTKClEvLqhKZCpWXJ2NA2bgB2jgnHdkpfZMudHpN3KhSKN
3T4pkeHKjASUlPT9ixpRGOfJ0DgJc71bemmGAzuVFBMjEXm9lIAX/oXLmM7Z8b+q
hUo6oCsYfrj1mAo/kiFxJGdWlM6OJAwKwpiuiDEpuTfAOlt5fcufgzNbaCI7Sm5y
WVQFDsPRbYLT1Z5sP3YWOOAn5LWZHNR9FU7XJoHIExDuYOAiDBASvvZagLl3T4Jy
vdbJGQaFLt8AUb0zoVliIk2KXthAWRAsuTLm3ZJ8phWXVUNBRwHsSdaUSywKwxo1
SBa3C8ieOXDnG/Eg9RyugLypfjwpFxN1NW5Lxxw5sSv9OZLhK9c6QLczV3jVhxhn
jvMoIaneFzOA/Ga+6MqpB01PtYfvDEtA61e1tGFdQ1u8mh4au1OsjVtJ8/ATfCxA
+8LsNH3/2QRiMmXnglmMjPj3Eh4zec6vWzSc0eL2b9WaapFEOy0ZQ3SuOkqG6Y9A
GW0PGZSgCxQ+/q39PXL4fFrkz/il6aRwN1YiavLyLmctM9RgJuNS0Dygtg+DgKag
/9F1F/BBIOBIk+yB8Pt9XFKrUolhkMX4z6E2SkoV+i03suutO9j6psdJpSuOZJMb
OFlO/N1Gg8TgDd+7e1HMaM2mhgCT/wVf1UkxCWfWtjdJo+A3PI0A3Tl3MruMJeZC
/rTa9NxCuMfEqGuwyQ1gxaBmk/vzJ+bQQlQp0cXVQMbhW8XLItrWzc71vA/yxZpP
hP6pd5ilM0IFyt1KLrAq+OWF/+vkeL13wBHTSyKxiMgnvzD+xG8j15uGPKMv3O75
ioWwMp5eWlGPnI9sdGVO53ASDgdDKJsBGRS7dRrqqpau39SR5+23udiYqhT982uC
Y74YdhLWqbi8n2QFqLt2OB4C24YblWwslBi4MYeqHBXIEzRwirNZ6MEqYCcTsU3Q
YwkZo8Yz6co48WwyCrauHZl6bSuIlEfNvBNX/wGfqIXEL6eMzlaaYKk83MUTZwfn
OTIhxtrIYTX2jfZHx8ZeQJC3QpUwTEU9U/ci0Gz9kDaYsNBmbqtx04Yx1XzvPino
tKKYAdvoRj1GwA01ZC/iHEI7cxMAkmKWWOw9A2IExIZBEB0x+O2b69qsL6NNpjqX
KffdimHk92AZX2PfjSgNivPWjDgfTkakhFR3mimmcQ594WOHiBGvvmvhv+S7y7W5
YGbAmOlVv6J31uJrcf7i5xA8N7DIn9GyR/oO6bOAFxRIKZf0HDODl9hpzPdVlwdS
C8ARsxDr/z9Ba6T9CJ9kDe9XJdNwCZ4ZVmfn0R4zeSDwN7ch2GZMOcRVkKEpZe19
nIAvncIzlV3spG9PKozXzoAbuTVOLBcJ2pvHCcpN3X0t6bMHk4QJjFah3/ubgjUL
tVjULwbzjMThjqYOArJ4pwug/pECyZ5T6MAFB9SkwwDfVFCS8coQa+FLfRmrxjgN
jYxFvM4QUF/CVUD883GyXjymYuvmRwZ1fIpxi8EjkCXDS+yqmqhVUXmMyNFKFCCN
V+Kke+dM+WcuPEcvhfCh9zMPcnzPO9p0uR+N1FgSMcW9gS48sS/kLv0vzF7ADaGT
+Q9Y5Vy1kFt6Ry/BeYkqxcWKLCHXTz6yVoY+Wzmavs9neDubsUCZOPUAUTLho0Ai
LLqlteNisK51r6kvjD6Jj7OeG0dUnPLmgWoioxwUlaSlkdhCB4dP/F2EBoWOSXyA
J4ZwKXVM6uE9LvVGqW57Xt4shAOf2jCMh/xIl3tvjkTu1yjwsr/MnbUnt+fg3hjz
a0SaX1+VXKKx2PeRyunhodjOlq/Z42kVG0dNFaBpQ0pMBdjTUIThKjjKzHaMwNIF
onhGmvYx6EEeiYb5os/3rdXdIfDFPYdmr5KjhK2gakGubAWVPrwoqtbaKMgtc6m3
iVhtlDGNHVWWR5ELxg0+ydcecm0QZ7OhYz1GNoPcl98fjU9OgGQ+/j1wrM8cX/TD
xpBDFUMT6eoOaOp+qQOIKozaYgzBUb0HHAglU6g4BlT7EInwZ8hSZpV80p/oHPPx
nkHRW1pmaNC6FLsHRXPoNdbuI6RUwNZVSXSKt9+A3wrecBpv55EKNBlpIMje2g4/
vUDy/+YU8f5jzRttDKZwN/kfJ/Sktqk1MKmWcY7wNEG1GFkFJbJQBaUVDIjRmnKE
OVLBXDHtpYBzrSVZq0oxF0l4QNWeLftacAn14P3dJ6PhCXdy8F0PaGcLWg0vSW6B
682FRGvPSiGdlFt3DGYn/VlaB0xJtthKyhpfxmuvZnyi8FmYRh1c9jJ6JtJRuVRT
YnN4mJ93pDEu/Sf/CTDr40hJdEpQEK1SlcuBgDFUTik6a8g08Qqa+hU4LASMmR1r
BW3tiDn0DxFUAr85Vs7yigjTJHE5Hzx4UIMvPOVePIJqHA4/qyRKipskmOkOZ+Qz
71+bpWU4ymTOKgrcWc/Xx1MImvucxK5sPkKLkVlVkM4Rp7BnsQx2DEzVEsfh5WPg
JgvvvGu6M4LzHQit6lxdWyhZVbhcCgDM1cZuFzNJE0gHFaptDdwKDZ0E8UH24DN2
QXQrTqKkSACbdN6WK7ghe7Z2KSY0J40rHMRk5o/IwhSLmewPjOrgPxL69OUQwnSM
U6k0VgXIdmtVgyjO4ufYOtewOYAEuIP5kVD2eXrinx+H4uUYEpBZI1HCSAtE7PNd
kRH5hjoiOCMO/3SBBSUcJF5u/mxpv2eyUjXrZOLhwc23FNXkRY2ejGUA5N7rWUwj
dfUoDBG6OFR94mlJCCYRiJBUtp7yla0/YseHMe5370ZVhcRxwUag5zNoq3HQeWF1
XHT/oFjw3K+X+eTaab67uiTR7JCxljL2C42CbDw9plWI7ZCG7Kov1WhsF1A7Ul59
+aJNXWzqs9u2Ur+Ev0dW37OvuFUUyBYFKYj7hXkq2j99O/9AHcagifPc2kTD5iaI
qK24hQ/cTPTAXgdS0kbkizq067pCIhti3zYCjhgKyTUf6MWwVLs1eH03NG0iRQgu
6D9Lc4wFBplgOrMTeRquIWR2rkTf7N4AsUkD7fTABdZmbYy0X31SWtyGILImVBrD
+tZLw2uyWGnU8R+W4LOmEXux/j9I7d2yZUvwD7qbVLICi65CUeCw+c6la8Ym68i3
OEgPJq17rjECyx1pFT/Hy0lOHgAUErFuEuiUyYCmX2gK516EDmi8Ohn7vKgYjVbl
qCpDZaVHHPQe7626BlLI8w==
`protect END_PROTECTED
