`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HRZTbGC8RIPIR9dI1MdmBdJRyupMaxMwl/4T0y4RYpqMl2RcEcgmNjD2Lvw348yj
H1ZJ7Ga/lPkBHL1ZqLryKQWMDAdApl17Jd5TfqP8yJT2j0YxwwRChDD0OJ4697Ig
MfdWO0QNMevWHuLreCOe4c7Mv5uTxLj1oIpDgtqTOOpWsLCPpngqcvQvmbc+evfj
p+5ccrVxUJLcYxM98a7IFHGlT9nMZNH9hsS0TV6GVxLCrwaZRyWnQF8kLk834JvZ
j266B0s2ddDTpQxKonyFHO9E/OL/kNiyQHgmU9i9AeQRA9GYS4+MJVHv5JYcl17u
27PI4czYTpVcFPArH3G55kVV4iUaVQOoGBUKOej30Bpo1XHl8rYmuY1oUk4BNMgB
J9pV6xFikW/wAk57xg6jWL9IIBreTqVgY13o0IowgeN7iGlMQPAzhmlqCjxJ3x5A
o+F3eth4UCTRgLeJEey8LvMGtTVUblina5hCZRyd9pAEiAZ7KMtycFckg6zZFv6U
h4xtlRtgBXU19jBtf1MvrM9Fm3Jb3Xwvt7yifQ9htxo=
`protect END_PROTECTED
