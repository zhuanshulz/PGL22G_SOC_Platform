`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O+4bq27xhxViLCDDtRN4chn5+jG91pftUut1FTQFbsVMO6RTeFEbyAfhrHsMJVwB
hiYOffPqYDw4AAF7AZtaMMYvKC01mjlIl/7G8lH163Grl/HgPiiaSS/o6cXJUNq8
hu5x4djD2MJhcwpaEkiACxBN7++GkmFjzKkVvLCTNBA1aBoeXelTduxBF1x96GIm
YaeHiaUrDT579ecyAbddXcJiVMPUptKE5rO2ICnBgy3B1VjeaAlpYH3Vb3q1/TVB
JNiYxvqHP8MgCgofY1VkaG2irMAAHOTNRceR7hnVcamklkqBcByvGXHJRbQbUzK7
15zes4QS7WjkyUin1p3qbE8+PSTYNnciWXZaEZlnoPp99e89TvkgEqz79eSYpDuA
ABe0WyJFprJtJcjHyPCBZnK8CCu2Z30+BH82JGRfgGqGtsia+fsOhN82DbT5q/i+
Ab1IvVQ3Y1ITGja9n1YjD8/H4dZ9Ly6cyIqdzxNyqilTO6UhJCstbkTV77VXG9lM
ofhGJEKulpouN9Wcr9f2fQOGUR83kI+n+vVtmPc49F1n5Q1eapw3A7EEBJBw5cmd
KJOCWwHGTLs3t6iVOkmGUCIyFxvL2FtdonguO0Ef0ijm8f+uyI/hGSlTMRe4lzPv
BmltyqMlGLxBXJpE7a5jyQYbYPaV8zk6QZArwFT63swveGExsjJj2vFTB934MSst
Jhgz8tIZsNkWPp1yYHiJTI8oYRqV8QmSFuHVnUEPj9BDqY7IzZmJLrea4lTgi/PO
UpGyLV/yrHnp/ZS72gAWGTzxQN361+HJgOIil64weBIy28UT3K8tPoU9SWn6EzQe
62NdXirGC0ucL2/59Z0fx6devBi39eRHd/QCjiVgsgHaefXIak8dmyPDnZbyP4Lt
e/3TcHECs5hmv6xGh1KBdRM+CZG2Bb1eaWIDGZVfWomldnvz+w7D7NvUP7M0Scw9
6yvrFozB10tCPTX+k17sZwffWdTalZX0fsaTUvkX9MqmdgWZAPBF9kl5XIaXdZH7
wvjc6f00kUxzT5C32la/3bj+nWlIvtRwuUMpnj7hXA2CmpJ1xqBFR0rTYvbLSHKl
hiqXSX59PPA/xzS04VuU4ATKmChKv8lkMrbZCrOAveQ5N0UYwVpQvT/rBXi7+RYh
Z8eeV7qRjbzISLNWp9JpcSR1nX18PayiU90SFNzaYRq1/YIw3R5MJu+v0G90FGEx
muuULaWeOQ/u/laVK4EcM9UcTAjJZ+7rg5ZAbH9taiSOaXrG5AhfBvfTLfAlRVxY
`protect END_PROTECTED
