`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tLYrmlYMMNCwyNkI2CtmuLZ3e9shSSnlZ9YqaLj1Y0sZ2pquC7m7zRusD3QR0d+R
cAlMB6d6JUBWz77tdLM50BQX8/ZeZ9GeSy5jKx7dZHZ5bk2yuRa9G1VRflHRhs71
6EE4gECVaZQFaxdcCgSi1KFmuI/ZnnLZOeK2tTPzfZ9X01aI8rMztBK1cOfUeK6K
R6OrtKJ4X0xcRIcaeElfUjZfNmByLwcR0HhcZbIprQZJd15eIErSAsevvjcYjgOn
e/OIS/Rlt3doT0LXtE/nBqhccIKUb9PHgvzxfZkZG9+rm2Dc6mqQDh3zSlhhCJNG
PzWT+0/IPvyVkqWj+dJS23F2RqiGUM6xAoczVjltZb5riH9b4x7VugcSNNSkPGsM
8THaaRFAV7/v8BBkC4KjrkYOm5Q0uaqIZxlrZvGZQX0hpTlM+F4zwZwwFCVJ7tYu
bTUW3S3o9QzUX3jiBJExKYXsj6Q/KjR3V73x7rNGGuMLbQ5DLAjK4zHiZRTg5gOa
d6K8uz4+j4OqTAGl1v6Odm/L46XdTW+FibVfTjIFjuNUzuja6/MLOIKBOOftrSxn
YZckivNbrD7T4hJdv2uibO7/q3mLK+J8ZJpvx589ZgMAFCRLwLPD28RBoCJcAzkn
SGQvR+b5St6E/RMgWaskTTQ/zUgHCSemzZvIs69VK2/tffFgQyDQig5DY4lF7VhZ
KfmI2WNVgIb3q2QqFFPObcyS9dWCz2L2N6tvQ5PdMpCrDHReyRN6tn6RcBLY8tlm
t2y/q8lYEW7Z892BPKIBtk6cNA2zY5aXq2s7/0EDStjNbLdoFfZ3X9fJNVKw8Eu5
N1nu9HKiTi20VxD0VjXUrrlABag90w6xdvW6S09cBGYFb9tZmCG53pe6IhKZruEh
feXMVnnHrofI5MvEBc/yfjBtB+l9PAfGrE/OWrJUX4HABrHNfEeO9hyU4W5+EIlU
/VUr7z7CFnDLs7zWgST6Q8LNG1STaktWHrXMH09Bho8zfIr7HUr6BVfd3NEG0Z6+
bRqmeTY7nllJktiN4lOwHYqlN1jwhq3jnY8b9B9EB+pAulf+yIJqGg/W5DT7WiXZ
L8ZmHYHJZCNwt7yVdFhoFpo2KWfmM3E74pmsuG1ZrIaFEVVqYh6OM9dJXp6fySct
+rgVB6c32D4mqmJ8BPY4fRg1ODEK8BjYTYL+iDWymHfv3iw/OzwVU11xw0V9tiMJ
nwUC00epc95OpvxR/fKzZViyOaH6Cg9H/4gmVZOPoM6WJsG4H6ZPjcoTxPTDWlqd
FmC8dp7bOLBS7OXYw+EPQ8NxsgcUH8gTi0NxCYaZW5C7bDTb3tdDMdWwB3BJRHJb
FlirqawdsSvyi0BWLdsYtC1TYXOSiKRDSEgRSBT/6+ly9S1E3AV12h1ieF1c0zD3
ZuUdTqCBUmHYapCncNPKttSRiKY4n1x7MpE2GIAG9AXebsyTVr4xW996IJM+xTpL
gWI493XT8BhkyTQJO0XVmZAB85AE0MeswSM9d25fDFaFn0205dG1EEUZgYmpb1u7
blvOBCIH6LSwKWWI939USwISPOKbBsfPET/sbMj5FAGeCTa7jwTmKoe4FgnHtSOe
Oc+9FbWHcEkGWUMzhffqPsdqbaOreTaLrpqQblFj1TBoWEE84KrnmzFBudMFqMOs
ClRXApZOI2cyZjpKrhdyFxzuiQpPFGVgjzvhQTFSQJ5NxMgRT3tqmQW518fkiFra
VO9TgszQdL3/gR+d2slKRTlMfZDDgooOeutLi653yWIH+3U+Es4TkzjzzsFthkYL
IqG9mwF2ITblAWNZ82P9EE0UiQNuG0WrcYkJGZeWkbb9f//qF96CDOPH+CnSnt0P
l96La/IMyVC4cznCd2dSieciBje8LMw8DWzRJXeeMoW7XyaJfcqgp6CY7CwjNCg4
oNZ86k+E9tEggxRWWvyK5DMC57kOsZLndRqoJxEFlMdqwqQ3lMVpbJxELv18io07
jN2dTMvRukbW+AXzmMEDtSkKloS2TUp7kWYV+1RtJRoAxPAaS2zjb2Gf5Cd3P5sZ
nVVclJd0MmKfwMMxaQtqBjcx5SQ5DAMst2ngOsL1/Ok=
`protect END_PROTECTED
