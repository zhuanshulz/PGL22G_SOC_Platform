`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nrtxMbx32saaHvY1Iod/66DuERmltdHIEPdFkKbtzM1A0FwNhFVEFnsjzRWdmKEr
ok7wS4VkvW322Jp4S36IrJf2ZoxeYDjIcAgSrSneru4tdKdRgogCZShbic/LRg1y
4OLMQ3gt3mrbmWhrbMVrJRNwUgD/SYknDCvXKcNj7SdL+Wokw9TsSlJ2Ly5jg4Pp
a+1goNnHqdXhDDdOPZb+7lXZDP3hFeGTb1Q6ssyCkPukS6iQzsaA6jVTHsx3EYno
iHuK/MEpgcOXjDnTZOE+Vld3bnshpPjZxy8sCY1QEK0oBz7KBg/qFb63MkhQMp8R
LsuLHvrxoTMvDzvXyKrAKTayLE05qoFN7CtOuXipbbEVrWjRIuGctv4cZIUWVQPJ
w76Ysz/fh8+yI2H6LWW7fFt5CSuFh53PbgjawtvcwfqEJRRSJuLPouL8AGYLG54G
PqK2itRZ4/uVdXKdACSOq+b8BKF8eVo3d2/9ZeGHVqw149JYTmdX38QmPOEm12hM
0TqQXepXFRZtVxulbyN96KE76k0etu04BUrH+gdCc0M1+sLlQNEFo5ZghX47ZSAb
JFHKIIRyoyWtpn6wHtFJzP2a9hdo3yhw8Whw4HqVMbL71EKDNSbpLGJXjMivP+9X
Ui8Gl/SPM6bsNW8hGIyLf3k4xuYeFzoC1+5xFJ5ZKMqxV7KWSwfYxfUOPC+ZrvUe
bCh+TeTEpWmdUco49G7GyIqdXyMhp9/VJFsgS0pni2OylCbd3mu5PdpNjkTnblr4
leJWffEd36gyfutO3bgFEW5qRg/YKSdggBC2C4EE6Rv7zdBToWNQRYt301lr4XCM
`protect END_PROTECTED
