`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eBkHkVgOog+ek5EWstE8Wt1mPQMbp5+n/OJ1FCrBMbOrLGqSkLRIYqXykFS+Ld1h
P/TqEDBAHRMD69lCVJssYGfvOrClXAo4uKZ7kcqdqersh2uMKIpHh20asMxu/whX
oBO+i/w74R6muE7ZyVvBNueQOzRUjh4Hnv5pyr/HMMqvEBMe1isFXvLnbq1Otw+L
0EOIZgSYw2Z6iivsfSUoqgXu6XsCK4doqMrWr6q08jLs7OVfIJrcWrW1JZBaKwa0
TktI27Agi1gRu/OkitrUyBUE92cI5Q+75Ffg3hExg1DO7ZmpkiKh5/Jo4y+XyVbk
0oteT+SjBLO0wi7KUXXrBq51tWNfUHfjqCHrjuU72N4Nq1LiD2+Y6SF6mF0hXmxf
q/ikvAXASS0FdimMW6F1cGqHHfb0jzfYW8vDWIn9d5gysbRrOzgpqicBqgSK/Rik
5xIWKW9GeabzBt2YnDWyTPq+vJJ9Mpwir5oN7hM74F/CO+5MDdoovUDOJR30jz/W
eHlAtQ/5jLSalB9o9INIXQZ1vs9ZQQQJ0Yxo+3tM4MGnabBZ+dzscm9bKnm/+Wh0
8S+u9lqQaBr3s/oMNK7Ql0FlDzMJD5+wy57IAwPg4/lkDGcY6kd1WoxFJhcBiJuQ
wBin68QlM/7tseyzmYR1fwyk64Ao/R/fmzhVFjXNvQeSBic/t8yLHOd/PX3L2fjW
VqBVQnDdlry5XdAHesDcKI25wRCFrefeBnZ5qcXkFsFQBJQF2KE2vPITOA8aHQUT
PIqrxX1FIUEn6WpIjU3aOeNHR1VJE2n4/iSuCYS3oCsLurom8krWTXICAA9lJGEi
`protect END_PROTECTED
