`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m0O3vVswV4OfGEwl38jAfDHQOFdUJ4dkCpO1Wvo/if1knZ/yDMIXayHXCGiarQ7G
zTSYVCNN+Xmo3abBLTU1v6KKSaIqaqDGyXce9SW4dpsq4W+SOhCFveO4bkL090F1
omoWhczKHJDJqN0+cjeSU0uuiFauRD9Em7gI63CWZlfa2ovRB8p93akdon6rA7bJ
MQdQRzCSRu+RV6lfquec5npOEdq2bGdVxjiA6G5ZfhWatMD6u6/WnoD5yOz/aB+Q
ZqdQ4fJkHGS9HF/YdkMCBtNWQrw3RrqAMZe4/zB0/+fQkKDdPbC60aYjkwXdSYoz
Nw3N4l/qH8u2WUm6SyV9DAx05uBU6SnCjMB928slC7h5NxGbzcQXauz3jG3sxlzn
dhHw+bwMizk9eEHBmf3XVKKFCv65r+CboZN3Ioj5Orjz0lu0JsjYyNidDgb4SMsf
wPl23z15ruKY/aykUu+CEq10w/MGv7YIYUtNqr9SXvZGP19DMtJxu+94ezSMGO67
JKpXMFKy6AQUUTL5vdltRA==
`protect END_PROTECTED
