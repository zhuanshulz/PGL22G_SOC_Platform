`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TuE7uZvsmR//3NOMwWeCwoZj3jRAGSE6057D7F1acO8HkF3QdTGeiZ94R36QV9kT
FjGB/L5/bpwMH+H9amUeIsxQPJPrHSPcWaT699rLcrbnRw+4BFSmuC7XX1O3rVzk
AJTWMAnKQ3MbILbuQDyWICY2QBiuO2L/i+AHzFinMSbbaG5wb3LTCePkj8y67l/V
SdNssxkNAkIAyFE0PYIJSOsDryVtK4W2phbC40A9fmm5gvIj2ffgKcC1Iyok1zCh
RVVloJe50CoMqbMj53Dux2YudTiQaHVIL/ujq1WSwOJUyuVBjRm8xoTDzbdIebhr
8mH6bvLYZrk54t+YezF9oyKOPpSmEnu8IjBV6zCHJTMoaHOSTjFBUdZDli+jWQNv
JUDaUO+YmzreJ5ChYAfl0iJqJCdCZ9X4/yZnotgVNFTKMEb7GDgaAuE7pjWgFqZ2
giqFCuMkEyTvh2Sso2nTiqBrfV54gbISDx80tIp6XhS5K5Cqnz5Q8X1RgeB8WWCZ
jzx/r0pOlz2tqKDaPMo4l7cwO4BTWA1N4mrR6BhtmZHDERSKDJZwpZuE+e7d57x3
pC+RB78z+Zx06KdElLKT29FmXTh9Aur8ovPgT+4fxv8NRRg6+93rn1HadL6ryFWY
+6oSYuQQNNW9v7E6EHI7t8JGgyG/c9NS1wxZeZJZfPAF0v/b09QrS11t9HfNw2u3
byGD12AmhRp766vycKRuke3FmCPgNNH4CN5vBjyMi/xiYMaRq8c00aTRshZ1iqM2
DJegxUZfyO7YsB1NJPW+PA==
`protect END_PROTECTED
