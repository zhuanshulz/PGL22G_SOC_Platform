`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hXMA2ZqhZxfXZJLAAiHh4KtnbiCr4fKV9UgnxazLoq1SUrXTgyMrfwmSvfuoyxOU
P4s/EY/KgXvFmtqPbqRdmjSgHc+PYkaFlsvPsm5OAQte4vRQHiSbi2W2LJfyFcM7
6gt1LDUy4P/Hf310ZMb3m4bE4qgxTIQNYTh3O9Xig1NIZum1NFWTAgGJop9iPDfw
aGqJFw9Wq9rnyVcmYhN9SYQlezinZ8cSRZs9spFdlNTXr0Mx9sWRN4Q151bx75bM
C4uEB8qGTYLRqgn9Zb2fyJN9XDIVjEDFby09V+UcR5KQL/iwZ4Vu87Kt4cJ2Kwm7
fB1KLUbVJbKNNHmMYi1pd/EPAGlinE26W4NB2nwvF8WmQQGecTxibQcforbwBoih
dQKQtfUV/5XDsYa16NO9as2g7iqr5Uo6drPaqi5Kt+RQfNdEzNznMMQF8VM0VAkc
dsTXAJfMoNbk2Atcq/xYqQD9KvnbekfP7AY6dtutg8UPMbvCd9YRxGCe1Iip1NmW
5X4yiOmxlACGD60MlHPI7uTi0Rfnk/3pQMb2JSK81DedP3uPzxll6dA6G7eAX1NQ
UgBZxzs2YbExnqqOoApNDDfD/r0jW+Vx2O+VUq73oVLKtHFGkLIeYVN94SpDbJK5
RtAKu0QvTkIYzHObv95djdRfoVqr8rH5s4JMw6cUmUQW3wd01FuoIT5NU4TozVMH
gzffWTVvqPIMZDkbx1lp+bCE7ZMFwiaG6hyh5ImGa0fUELOGi/bbkDjzcnzn3kRG
7cPD55oIWPQFV9OoDr4mhrp8mPCd2b3hkjw1KSb9qy3ITUdGTU5rsSij7SuXgN85
gr2SGsTZ3V/xVBk5RwR4J0oAf8byOh+zEGiQAOS5l6tufk4PkCWFLD3ipkhMp4Zm
DMGtLw297FrHNTeirv1gTaTApjgSaHmI0SaQT1Pl3zEFfib797aa2NR275mzChdv
6WbVvRbVgNtD3N4sHG536ufTg6wY+fXByFFsTtAydzDmsWu5mTwJKxvXzncIJaYC
vsNwAHtZoGmwSMFg0ftOwXIicrqeai4GVLXAu9pUEvGGWVqyZmq8urHmkuypy6rd
YST9OQu4UmUCI2HEXumiOjBOhi/JPi9M6ww9m0YdkkllSvxYIwdwrFeanQ+0p8jP
UwJb5/RMuxlEreCrGZDQ048Ompr33wsuS6DzbkrcaTyGIZEAnqImnt76CZEmE6ou
yIpg548tkIOr0q3X+A4FKpf1VbL+7so6Yu5cwvQcUy6I877gDl1HBylvb4Geco2o
xGcJ0zhahmgkb4inSJes+3Xd5ESJ74uLINM0pAEK9EX/LbHeFWa2dlupvdl03bIV
XUbl5h2uFEWoXxxt7enhoUjf/Y+KUoNzeLFumECsAmn1rigXY0aBZOWM5kJ+atA9
CYABnQFTUz9JnJL6MqN2xILt4AZzuepkp5CjeQ8pgcOLF94Io6BPDUQ3En0iB0bL
L8zGjZcagtgd5u8GXcxuIJvtGjz2NwLraILdM/10xJFigmsZ4aWB7teOUE3yriOy
23w/prBxDxfnc+U6zCfQHtTYwaQx2meBYBAg37+lFXCqGby6qmLtauTwuTohMzm/
BQBe002gPRZYzADayVsDFqyuHerOPcbAtpS8uhGulRo3kLiVm2syU/53o53UxsH0
2YAt5zUReUNRDYIZvOnlCm9oCKTCaRAI0JcHm8sU+c+/ZsgFzG88198PsnLZz7he
Y7u+2bygMnRs8QZkZs/4xhyqbbv2PQT+9IYZlbFBzs0=
`protect END_PROTECTED
