library verilog;
use verilog.vl_types.all;
entity V_HSSTHP_HPLL is
    generic(
        PMA_REG_REFCLK0_FAB: string  := "REFCLK0";
        PMA_REG_REFCLK1_FAB: string  := "REFCLK1";
        PMA_REG_HSST_LAST_REFCLK0_SEL: integer := 0;
        PMA_REG_HSST_NEXT_REFCLK0_SEL: integer := 0;
        PMA_REG_HSST_LAST_REFCLK1_SEL: integer := 0;
        PMA_REG_HSST_NEXT_REFCLK1_SEL: integer := 0;
        PMA_REG_LANE0_PLL_REFCLK_SEL: string  := "REFERENCE_CLOCK_0";
        PMA_REG_LANE1_PLL_REFCLK_SEL: string  := "REFERENCE_CLOCK_0";
        PMA_REG_LANE2_PLL_REFCLK_SEL: string  := "REFERENCE_CLOCK_0";
        PMA_REG_LANE3_PLL_REFCLK_SEL: string  := "REFERENCE_CLOCK_0";
        PMA_REG_HPLL_REFCLK_SEL: string  := "REFERENCE_CLOCK_0";
        PMA_REG_REFCLK0_IMPEDANCE_SEL: string  := "100_OHM";
        PMA_REG_REFCLK1_IMPEDANCE_SEL: string  := "100_OHM";
        PMA_REG_PLL_JTAG0_VTH_SEL: string  := "60MV";
        PMA_REG_PLL_JTAG0_LPF_RSEL: string  := "20K";
        PMA_REG_PLL_JTAG1_VTH_SEL: string  := "60MV";
        PMA_REG_PLL_JTAG1_LPF_RSEL: string  := "20K";
        PMA_REG_IBIAS_DYNAMIC_PD_7_0: integer := 255;
        PMA_REG_IBIAS_DYNAMIC_PD_15_8: integer := 159;
        PMA_REG_IBIAS_DYNAMIC_PD_18_16: integer := 7;
        PMA_REG_IBIAS_STA_CUR_PD_2_0: integer := 0;
        PMA_REG_IBIAS_STA_CUR_PD_8_3: integer := 0;
        PMA_REG_BANDGAP_VOL_SEL: string  := "BANDGAP";
        PMA_REG_BANDGAP_TEST: integer := 0;
        PMA_REG_CALIB_CLKDIV_RATION: string  := "DIV1";
        PMA_REG_HPLL_REFCLK0_PD: string  := "ON";
        PMA_REG_HPLL_REFCLK1_PD: string  := "ON";
        PMA_REG_TX_RATE_CHANGE_SEL0: string  := "CLK_FROM_HPLL";
        PMA_REG_TX_RATE_CHANGE_SEL1: string  := "SEL_SYNC_RATE_CHANGE";
        PMA_REG_TLING_IMPEDANCE_CTRL: string  := "125OHM";
        PMA_ANA_COM_REG_142: integer := 0;
        PMA_ANA_COM_REG_143: integer := 0;
        PMA_ANA_COM_REG_145_144: integer := 1;
        PMA_ANA_COM_REG_146: integer := 0;
        PMA_ANA_COM_REG_147: integer := 0;
        PMA_ANA_COM_REG_148: integer := 0;
        PMA_ANA_COM_REG_149: integer := 0;
        PMA_ANA_COM_REG_151_150: integer := 1;
        PMA_ANA_COM_REG_152: integer := 0;
        PMA_ANA_COM_REG_153: integer := 0;
        PMA_ANA_COM_REG_154: integer := 0;
        PMA_ANA_COM_REG_155: integer := 0;
        PMA_ANA_COM_REG_157_156: integer := 1;
        PMA_ANA_COM_REG_158: integer := 0;
        PMA_ANA_COM_REG_159: integer := 0;
        PMA_REG_COM_PD  : string  := "FALSE";
        PMA_REG_COM_PD_OW: string  := "FALSE";
        PMA_REG_HPLL_DIV_CHANGE_3_0: integer := 0;
        PMA_REG_HPLL_DIV_CHANGE_11_4: integer := 0;
        PMA_REG_HPLL_DIV_CHANGE_15_12: integer := 0;
        PMA_REG_HPLL_VCOLDO_EN: string  := "TRUE";
        PMA_REG_HPLL_REFCLK_DIV: integer := 1;
        PMA_REG_HPLL_CHARGE_PUMP_PD: string  := "WORK";
        PMA_REG_HPLL_CHARGE_PUMP_CTRL: integer := 7;
        PMA_REG_HPLL_LPF_RES_SEL: string  := "5K";
        PMA_REG_HPLL_VCO_EN: integer := 1;
        PMA_REG_HPLL_PCURRENT_SEL1: integer := 0;
        PMA_REG_NFC_STIC_DIS_N: integer := 0;
        PMA_REG_HPLL_FBDIV0: integer := 10;
        PMA_REG_HPLL_FBDIV1: integer := 10;
        PMA_REG_HPLL_PHASE_SEL: string  := "DIV2";
        PMA_REG_HPLL_CFG_7_0: integer := 3;
        PMA_REG_HPLL_CFG_15_8: integer := 0;
        PMA_REG_PLL_LOCKDET_RESET_N: string  := "FALSE";
        PMA_REG_PLL_LOCKDET_RESET_N_OW: string  := "FALSE";
        PMA_REG_READY_OR_LOCK: string  := "FALSE";
        PMA_REG_PLL_READY: string  := "FALSE";
        PMA_REG_PLL_READY_OW: string  := "FALSE";
        PMA_REG_PLL_LOCKDET_REFCT_0: string  := "TRUE";
        PMA_REG_PLL_LOCKDET_REFCT_2_1: integer := 3;
        PMA_REG_PLL_LOCKDET_FBCT: integer := 7;
        PMA_REG_PLL_LOCKDET_LOCKCT: integer := 4;
        PMA_REG_PLL_LOCKDET_ITER: integer := 3;
        PMA_REG_PLL_UNLOCKDET_ITER: integer := 2;
        PMA_REG_PLL_LOCKDET_EN_OW: string  := "FALSE";
        PMA_REG_PLL_LOCKDET_EN: string  := "FALSE";
        PMA_REG_PLL_LOCKDET_MODE: string  := "FALSE";
        PMA_REG_PLL_LOCKED_OW: string  := "FALSE";
        PMA_REG_PLL_LOCKED: string  := "FALSE";
        PMA_REG_PLL_UNLOCKED_OW: string  := "FALSE";
        PMA_REG_PLL_UNLOCKED: string  := "FALSE";
        PMA_REG_PLL_LOCKED_STICKY_CLEAR: string  := "FALSE";
        PMA_REG_PLL_UNLOCKED_STICKY_CLEAR: string  := "FALSE";
        PMA_REG_LOCKDET_REPEAT: string  := "FALSE";
        PMA_REG_NOFBCLK_STICKY_CLEAR: string  := "FALSE";
        PMA_REG_NOREFCLK_STICKY_CLEAR: string  := "FALSE";
        PMA_REG_RESCAL_EN: string  := "FALSE";
        PMA_REG_RESCAL_RST_N_OW: string  := "FALSE";
        PMA_REG_RESCAL_RST_N_VAL: string  := "FALSE";
        PMA_REG_RESCAL_DONE_VAL: string  := "FALSE";
        PMA_REG_RESCAL_DONE_OW: string  := "FALSE";
        PMA_REG_RESCAL_I_CODE_VAL_1_0: integer := 0;
        PMA_REG_RESCAL_I_CODE_VAL_5_2: integer := 0;
        PMA_REG_RESCAL_I_CODE_OW: string  := "FALSE";
        PMA_REG_RESCAL_ITER_VALID_SEL: integer := 0;
        PMA_REG_RESCAL_WAIT_SEL: string  := "FALSE";
        PMA_REG_I_CTRL_MAX: integer := 45;
        PMA_REG_I_CTRL_MIN_1_0: integer := 3;
        PMA_REG_I_CTRL_MIN_5_2: integer := 4;
        PMA_REG_RESCAL_I_CODE_3_0: integer := 0;
        PMA_REG_RESCAL_I_CODE_5_4: integer := 2;
        PMA_REG_RESCAL_INT_R_SMALL_VAL: string  := "FALSE";
        PMA_REG_RESCAL_INT_R_SMALL_OW: string  := "FALSE";
        PMA_REG_RESCAL_I_CODE_PMA: string  := "FALSE";
        PMA_REG_REFCLK0_JTAG_OE: string  := "FALSE";
        PMA_REG_REFCLK1_JTAG_OE: string  := "FALSE";
        PMA_REG_RES_CAL_EN: string  := "FALSE";
        PMA_REG_HPLL_RSTN: string  := "FALSE";
        PMA_REG_HPLL_RSTN_OW: string  := "FALSE";
        PMA_REG_HPLL_PD : string  := "FALSE";
        PMA_REG_HPLL_PD_OW: string  := "FALSE";
        PMA_REG_LC_VCO_CAL_EN: string  := "FALSE";
        PMA_REG_DIV_CALI_BYPASS: string  := "TRUE";
        PMA_REG_CALIB_WAIT: integer := 3;
        PMA_REG_CALIB_TIMER: integer := 0;
        PMA_REG_BAND_LB : integer := 0;
        PMA_REG_BAND_HB_0: string  := "TRUE";
        PMA_REG_BAND_HB_4_1: integer := 15;
        PMA_CFG_HSST_RSTN: string  := "FALSE";
        PMA_CFG_COMMPOWERUP: string  := "OFF";
        PMA_CFG_PLLPOWERUP: string  := "OFF";
        PMA_PLL_RSTN    : string  := "FALSE"
    );
    port(
        P_CFG_RST_HPLL  : in     vl_logic;
        P_CFG_CLK_HPLL  : in     vl_logic;
        P_CFG_PSEL_HPLL : in     vl_logic;
        P_CFG_ENABLE_HPLL: in     vl_logic;
        P_CFG_WRITE_HPLL: in     vl_logic;
        P_CFG_ADDR_HPLL : in     vl_logic_vector(11 downto 0);
        P_CFG_WDATA_HPLL: in     vl_logic_vector(7 downto 0);
        P_CFG_READY_HPLL: out    vl_logic;
        P_CFG_RDATA_HPLL: out    vl_logic_vector(7 downto 0);
        P_CFG_INT_HPLL  : out    vl_logic;
        P_COM_POWERDOWN : in     vl_logic;
        P_HPLL_POWERDOWN: in     vl_logic;
        P_HPLL_RST      : in     vl_logic;
        P_HPLL_LOCKDET_RST: in     vl_logic;
        P_RES_CAL_RST   : in     vl_logic;
        P_TX_SYNC       : in     vl_logic;
        P_TX_RATE_CHANGE_ON_0: in     vl_logic;
        P_TX_RATE_CHANGE_ON_1: in     vl_logic;
        P_HPLL_DIV_SYNC : in     vl_logic;
        P_REFCLK_DIV_SYNC: in     vl_logic;
        P_HPLL_VCO_CALIB_EN: in     vl_logic;
        P_RESCAL_I_CODE_I: in     vl_logic_vector(5 downto 0);
        P_RES_CAL_CODE_FABRIC: out    vl_logic_vector(5 downto 0);
        P_REFCK2CORE_0  : out    vl_logic;
        P_REFCK2CORE_1  : out    vl_logic;
        P_HPLL_READY    : out    vl_logic;
        P_HPLL_REF_CLK  : in     vl_logic;
        P_HPLL_DIV_CHANGE: in     vl_logic;
        P_TEST_SE_N     : in     vl_logic;
        P_TEST_MODE_N   : in     vl_logic;
        P_TEST_RSTN     : in     vl_logic;
        P_TEST_SI0      : in     vl_logic;
        P_TEST_SI1      : in     vl_logic;
        P_TEST_SO0      : out    vl_logic;
        P_TEST_SO1      : out    vl_logic;
        P_FOR_PMA_TEST_MODE_N: in     vl_logic;
        P_FOR_PMA_TEST_SE_N: in     vl_logic;
        P_FOR_PMA_TEST_CLK: in     vl_logic;
        P_FOR_PMA_TEST_RSTN: in     vl_logic;
        P_FOR_PMA_TEST_SI: in     vl_logic;
        P_FOR_PMA_TEST_SO: out    vl_logic;
        PMA_HPLL_READY_LEFT: out    vl_logic;
        PMA_HPLL_READY_RIGHT: out    vl_logic;
        PMA_HPLL_REFCLK_LEFT: out    vl_logic;
        PMA_HPLL_REFCLK_RIGHT: out    vl_logic;
        PMA_LPLL_REFCKOUT_CH0: out    vl_logic;
        PMA_LPLL_REFCKOUT_CH1: out    vl_logic;
        PMA_LPLL_REFCKOUT_CH2: out    vl_logic;
        PMA_LPLL_REFCKOUT_CH3: out    vl_logic;
        PMA_RES_CAL_LEFT: out    vl_logic_vector(5 downto 0);
        PMA_RES_CAL_RIGHT: out    vl_logic_vector(5 downto 0);
        PMA_TX_RATE_CHANGE_ON0_LEFT: out    vl_logic;
        PMA_TX_RATE_CHANGE_ON0_RIGHT: out    vl_logic;
        PMA_TX_RATE_CHANGE_ON1_LEFT: out    vl_logic;
        PMA_TX_RATE_CHANGE_ON1_RIGHT: out    vl_logic;
        PMA_TX_SYNC_HPLL_LEFT: out    vl_logic;
        PMA_TX_SYNC_HPLL_RIGHT: out    vl_logic;
        PMA_TX_SYNC_LEFT: out    vl_logic;
        PMA_TX_SYNC_RIGHT: out    vl_logic;
        PMA_HPLL_CK0_CH0: out    vl_logic;
        PMA_HPLL_CK0_CH1: out    vl_logic;
        PMA_HPLL_CK0_CH2: out    vl_logic;
        PMA_HPLL_CK0_CH3: out    vl_logic;
        PMA_HPLL_CK90_CH0: out    vl_logic;
        PMA_HPLL_CK90_CH1: out    vl_logic;
        PMA_HPLL_CK90_CH2: out    vl_logic;
        PMA_HPLL_CK90_CH3: out    vl_logic;
        PMA_HPLL_CK180_CH0: out    vl_logic;
        PMA_HPLL_CK180_CH1: out    vl_logic;
        PMA_HPLL_CK180_CH2: out    vl_logic;
        PMA_HPLL_CK180_CH3: out    vl_logic;
        PMA_HPLL_CK270_CH0: out    vl_logic;
        PMA_HPLL_CK270_CH1: out    vl_logic;
        PMA_HPLL_CK270_CH2: out    vl_logic;
        PMA_HPLL_CK270_CH3: out    vl_logic;
        PMA_IPN50U_IN   : inout  vl_logic_vector(7 downto 0);
        PAD_REFCLKN_0   : in     vl_logic;
        PAD_REFCLKP_0   : in     vl_logic;
        PAD_REFCLKN_1   : in     vl_logic;
        PAD_REFCLKP_1   : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of PMA_REG_REFCLK0_FAB : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_REFCLK1_FAB : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_HSST_LAST_REFCLK0_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_HSST_NEXT_REFCLK0_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_HSST_LAST_REFCLK1_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_HSST_NEXT_REFCLK1_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_LANE0_PLL_REFCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_LANE1_PLL_REFCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_LANE2_PLL_REFCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_LANE3_PLL_REFCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_HPLL_REFCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_REFCLK0_IMPEDANCE_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_REFCLK1_IMPEDANCE_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_PLL_JTAG0_VTH_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_PLL_JTAG0_LPF_RSEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_PLL_JTAG1_VTH_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_PLL_JTAG1_LPF_RSEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_IBIAS_DYNAMIC_PD_7_0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_IBIAS_DYNAMIC_PD_15_8 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_IBIAS_DYNAMIC_PD_18_16 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_IBIAS_STA_CUR_PD_2_0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_IBIAS_STA_CUR_PD_8_3 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_BANDGAP_VOL_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_BANDGAP_TEST : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_CALIB_CLKDIV_RATION : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_HPLL_REFCLK0_PD : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_HPLL_REFCLK1_PD : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_RATE_CHANGE_SEL0 : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_RATE_CHANGE_SEL1 : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TLING_IMPEDANCE_CTRL : constant is 1;
    attribute mti_svvh_generic_type of PMA_ANA_COM_REG_142 : constant is 2;
    attribute mti_svvh_generic_type of PMA_ANA_COM_REG_143 : constant is 2;
    attribute mti_svvh_generic_type of PMA_ANA_COM_REG_145_144 : constant is 2;
    attribute mti_svvh_generic_type of PMA_ANA_COM_REG_146 : constant is 2;
    attribute mti_svvh_generic_type of PMA_ANA_COM_REG_147 : constant is 2;
    attribute mti_svvh_generic_type of PMA_ANA_COM_REG_148 : constant is 2;
    attribute mti_svvh_generic_type of PMA_ANA_COM_REG_149 : constant is 2;
    attribute mti_svvh_generic_type of PMA_ANA_COM_REG_151_150 : constant is 2;
    attribute mti_svvh_generic_type of PMA_ANA_COM_REG_152 : constant is 2;
    attribute mti_svvh_generic_type of PMA_ANA_COM_REG_153 : constant is 2;
    attribute mti_svvh_generic_type of PMA_ANA_COM_REG_154 : constant is 2;
    attribute mti_svvh_generic_type of PMA_ANA_COM_REG_155 : constant is 2;
    attribute mti_svvh_generic_type of PMA_ANA_COM_REG_157_156 : constant is 2;
    attribute mti_svvh_generic_type of PMA_ANA_COM_REG_158 : constant is 2;
    attribute mti_svvh_generic_type of PMA_ANA_COM_REG_159 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_COM_PD : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_COM_PD_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_HPLL_DIV_CHANGE_3_0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_HPLL_DIV_CHANGE_11_4 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_HPLL_DIV_CHANGE_15_12 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_HPLL_VCOLDO_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_HPLL_REFCLK_DIV : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_HPLL_CHARGE_PUMP_PD : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_HPLL_CHARGE_PUMP_CTRL : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_HPLL_LPF_RES_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_HPLL_VCO_EN : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_HPLL_PCURRENT_SEL1 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_NFC_STIC_DIS_N : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_HPLL_FBDIV0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_HPLL_FBDIV1 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_HPLL_PHASE_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_HPLL_CFG_7_0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_HPLL_CFG_15_8 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_PLL_LOCKDET_RESET_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_PLL_LOCKDET_RESET_N_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_READY_OR_LOCK : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_PLL_READY : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_PLL_READY_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_PLL_LOCKDET_REFCT_0 : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_PLL_LOCKDET_REFCT_2_1 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_PLL_LOCKDET_FBCT : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_PLL_LOCKDET_LOCKCT : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_PLL_LOCKDET_ITER : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_PLL_UNLOCKDET_ITER : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_PLL_LOCKDET_EN_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_PLL_LOCKDET_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_PLL_LOCKDET_MODE : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_PLL_LOCKED_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_PLL_LOCKED : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_PLL_UNLOCKED_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_PLL_UNLOCKED : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_PLL_LOCKED_STICKY_CLEAR : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_PLL_UNLOCKED_STICKY_CLEAR : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_LOCKDET_REPEAT : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_NOFBCLK_STICKY_CLEAR : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_NOREFCLK_STICKY_CLEAR : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RESCAL_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RESCAL_RST_N_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RESCAL_RST_N_VAL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RESCAL_DONE_VAL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RESCAL_DONE_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RESCAL_I_CODE_VAL_1_0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RESCAL_I_CODE_VAL_5_2 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RESCAL_I_CODE_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RESCAL_ITER_VALID_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RESCAL_WAIT_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_I_CTRL_MAX : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_I_CTRL_MIN_1_0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_I_CTRL_MIN_5_2 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RESCAL_I_CODE_3_0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RESCAL_I_CODE_5_4 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RESCAL_INT_R_SMALL_VAL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RESCAL_INT_R_SMALL_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RESCAL_I_CODE_PMA : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_REFCLK0_JTAG_OE : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_REFCLK1_JTAG_OE : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RES_CAL_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_HPLL_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_HPLL_RSTN_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_HPLL_PD : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_HPLL_PD_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_LC_VCO_CAL_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_DIV_CALI_BYPASS : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_CALIB_WAIT : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_CALIB_TIMER : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_BAND_LB : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_BAND_HB_0 : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_BAND_HB_4_1 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CFG_HSST_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CFG_COMMPOWERUP : constant is 1;
    attribute mti_svvh_generic_type of PMA_CFG_PLLPOWERUP : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL_RSTN : constant is 1;
end V_HSSTHP_HPLL;
