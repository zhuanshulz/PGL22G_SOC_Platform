`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M+xPP6IpmgOaEb/nlee/oLpk/EcxWJpVZ6HMXGuhtFL4Vk982oyQPqrI1pzxtBTQ
WVEoPgY1M5k5rNyVNqx00wLMq2ugW2rt15gklz07GLYjakfRb/nEh3/zM0196NOq
X5phAovFewZ0keNt4YSZJ8wpEz14OcDB9QFHiPbJbcCS0w9MfL4Dve9TYSuNtZFx
nodHV+WSRhxXS1wAJfFcoNMXnODTpMMiBkUu/5K1dU+VpB/XcVo+uHwj9aZePcau
jVbbGRhdiwcb1J+JWl3c1EKtZPeG9OljiTqvrsHmU/WsODWRoDeYFCbRCFJljRU5
kMUUYppW3CHn1u2obBgYBw==
`protect END_PROTECTED
