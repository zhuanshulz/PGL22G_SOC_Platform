`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eFRIy+z9VAeLYgPJBbTY+MsIGbVSIO/XMbQwuXK5RTNsso2WVjroh/NdpSy92KiV
zOPz97Z39cnwtSC0vTiWHNEEybiAtL9D9LaAXO/kK7UXI+cN1fJfR7/3F7lXVaKe
n6OgJDFSRmhviIbeTKO3Ovy10Y5a+84e2WloQBscrvnLBHTZp459Z7iNGrehicPh
t2feAe4Y6TluCGKF8KBzAzS5OjqJwdzaEsrf5PCg97HaOCsL6uDA1uLB8K6KxqNG
Jv0GverT4Yxltk/kZK/Vty0tRWVEKX8S8BLmA8qW62oOED8XVEItRJnfHBsSJQW+
Ub9rNbkoC+pl1sEnvHVwgb70gm84DpWHCB0YGgaesfYnFtl+HEBUn/b2GEQ+SBMr
XZhrEITwbEPotm63oosYRAbc2e2GkE0hDSye+47mBufBt4sBV3UXsSeqn4fZYw52
3HRuj6T86ru3vmwrFHrp3pjUr2XroB0gYy31uZncseL4dRJmv8Ca0sxZSwtOa197
qjXlC9XJ+mmTvdikIxeMXbQfasg7Seqq7R24+8elDkeczCBVtHkDUX9d801DM2Zh
+8WAnLy1bG00Bl3OudJjznkXsSwLuNO67fZkx2+fnLMDyq2PNhXD+oVgNpB/24R6
H7js6Lzt9d1fsbdThmTcHUWgab83G4Jgp5YcGWI5imfqljB0QWD8fzzfYhMUMYfR
XhgqTeOu1MIt1fYyWscwUTx8hhqWC/wsm7hc1k4Yh+lHL8tXKDmHv53bLZEw+mJA
gcVoB0/ZnNF3fcuuTvdgS+HnaQSTWkUhzSuyXGxvtFfihKBWTrcrtUBtx8y929CH
IZk4wDmdOXfZftymeLX8UaHFU5sx8bMBJVXYrmXMaajjBtX27xjVu++OFv1czB12
lUHz1XED0Mqtam/BW1iUTblBu3xMDbSFkdjGfEqfAGTW7bwzYF+Mxkm6M57yBUck
MokN8VubnARCzVZfQgNqwON/tRWxDsGBddlTEyrLk5vE2StILCeEbOxHM6s70bHx
wenizZI0A2AP5pRkkSTEiY1a4RwUTKk8Nu2BY+zg7xpeDjcpm0tRklwUcLzHTESC
0mDvyvyuHOW0aelSay1mQkTOgXHM+hgoF2XjuMVno7Rmc1GUF7HrKe61dOlKhEpT
DeKuCcxTziaS7fzbPIT1EFncNb18R6Qhw1gQh5KQDe1EB+yBhkaCfdxYVoDtySyl
klk2MZOT9v4UL1MNmV2YwQFzPhhnAq2LaUwMrddgObZNuumG/zwXTUMKLnXQRN/b
hxIBf1e+LaJjpYOR916l52WBEElnXyFi9woT73ycjA5F9U4uzHDAz/nPCVKY+IIX
DCNSCQiwRpZiXT3SvOdFuv2e2hp40LB1tTJhJd/Epiw7K/o3ETf8sa/M9LUGaUdZ
PV7A3hxDWbe/yDg8OTRJBHmll0FJ46BmWTQ+LHdEN8T2TnCTezbKCgjsnp+H2ZcD
tMa1OwSdpBeONidLf2zAPHbIDIYnBiB45etC+42l1bbxPe3vMXEGY55rCfVpKaZK
X/QtOhuwxiBrhF5G0NDZqr5pRwnc9pnfX50LW+/MawNMIEGW99VFfcXJSZsDXDT5
n48pAnV1TD7QXCRYW6vTT+ySnSs0dVpFxyJ5Sd3rXqdXdEq71GQiU65wWlVzY6b/
RC09oDFylBdz0GmdqU91cT8xxAE2RlkQ91oI2tJYbs4rYJGfzlYKlae6V0SENGNi
BDvOX6rSgKu8LIdFdXw/0ROxK5hq/NZTkBjSoSl8RrvTNU6QJJPkHkgpywQQdfn6
BPoy1fZPQFfA5Lp7bNpP/5Sqmi7bfXhJZbbG9eodvHqDqLtNo5sYK5TBw0ZEvhpX
mwr/cn8fhGmt42abcctAmCMVs0os7w2b7p6e+i1NUVvZl/PkipvgZ6EE5pRMmkCx
q9fj/CPmUUryAYgRMaBJHLPaEWRheiLH4VFqIfdMSBdWzwQHMg9nG8GebbmfB/mS
7q6bfBIoSY78Oeo6SUlJXoE8jY3rQDrd5Lh+4bx1HAxb0F2fGXJyg/bvPoceP3CK
`protect END_PROTECTED
