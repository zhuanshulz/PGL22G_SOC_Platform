`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lOvZbWK7QdAzCytMFsFZR/itUbs1WAPWxMNKoEwZuw0Qv1RBwNZ20CfB0dtJ/95g
8u7BqN7ZvKsWoPdp//fGDuBa+0cre7ZT2kPu/NY0PIKFm5ftr4NUg2RuqszFOCoD
VMR5YbyzyNHvwRPXoGSjqQhp1bL+6L1B/iiNl68GoLW8OLKLi1VJuiwyszGazGN8
cxQzevmnrLt6m73wlpTu42mvX5DWV+O0jaXB4E6UgyYRSFmWxTWETt2N7vp+GChS
WRIzY7LgViNpmD0CbK4yrBdwCu4QPPhvV7aiFCAWbkLwx4ORg4juJwbFOI3qDu5n
bfW5V2KNOLmMFm5AKRtc7pVvJlppnN1CEkDMVwsI4BKIFHx2eBlvl+NKK1SKMnmd
a92JDGpVeUsbsk+gbnpe0h20jBgv3xacy7HZOoR+7pYRcvJAJlSdOJ5ZYRnaxHZS
oIJbXAjI1Vor2/p7DEj/VO+3CU5C3un8QzEKxSIGWcx1eI3X/uNQymqrkN2NxvdV
LjiEz3t0dqfqzJmFzFLi6+Ik9i163adRyNcCygOnghnqKDcE0E8Xa8XXl2AHx2V2
x3AC39V+06NeZNZ2ZbsyW9t1+XMr1b1bVn/npolSgEcRMG2nbQ9ai1Ij6r47AhNM
nyHXfqeo+qTEbK6tuAKAhl1EEOzkXTSKIHtMUyo9tos=
`protect END_PROTECTED
