`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s26GZ5HqXBR9V10jY5HgptcDuGFaFdvo3YpiBLczjcjl43ZK870KszRBoNqYb1gf
DxrQ8JF4eHGm0ZPjydFI9nNCPAP36sknHKgZG0J8eksCHdpveWmTf1dkcQIskgCL
q2KnDYJVpF0F9SM7Vf+evgAzLBy4stfWSlb+QLU/N0ufuP5lD/at97Hrk2gS8SPw
7WyHgJkznDPs5nLBgQxUwVpvx44nYTQY7/nFqa1zUf5HLGl9vCdeOLvPB6ykuQMA
NMRdiisTSRddYOx7JS5gIw==
`protect END_PROTECTED
