`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7FO9axif3kPQo8Dq2PtmzQzFDW0zqfa3BPFyF26GbuuRm7EOoY9A1l9Ey0qIbZXf
KBCtWr6OL/6WXdmAc0w8Z5jeJnTL+rxTKybLXXWhPqJuT1IbOGwxqhZhAt8VFUj6
bsasOIjoNee0S73uMl1b7CgLSIV8muzG+IWfJVyz9SZQE8Y8i2YUtlvyU+CuqRRi
ijrF507MqPsXRDxtRYsEuGcT/51zC1Y22CBpSqhrYJh6kngO4v4H5y04n1jos7lJ
XLWjEqZGxtH6L3RbWwGMsie/8kLDiOpyOe48nKLHaON4hfoGwTmlA/QvCQjCTeBE
ScwuJjeFH/GHFjkx8MixiFaDLQnRgPz3A+kzgUUjPsVLBv/rd1JeMqf9WFiAO2jM
jpwf9KUA2v1SvS8TX+RZ1LuYNtNSeyFTmCgvBur4sVvKGasu6vDu1274oVxTDsoF
hPnHrAvyUDOcxUl+hGs50DzBQgOTlcuNFs94SK8EAoCoHzg82r7FQvFEp9GdtSfd
WAHqGXBJ7tQOGdGR56PkFYym7iazd8dKVOAaDndHobjdLmFtOWYQX/w7HEqvjrKG
lZP60kp/dPhadkv89UK2viu5QBprOM91gEigmZnf67+n+ZhS5U2ZmoAEnaTVMkVo
8kt9E/wzNycY36i74jYrt3tfQ/zlo9HKIRzZxytcOSoSEPgS3aLZ6BXovKM/DRTA
CY6Ngu/OnFHKxCPUSEvUgqNBJf3oMMXb2bAPI/b5wOTkAXmalmxsz41gVBqSg/Ix
U8CYiFjho6rln+HXGgVEG0XuhSul6ftsm3NLeK4wNKrShoJtlIoZWFlRfaqa6ruT
5v73vekfCh+lno79His0F9cW5QSSSxfgxwzqdHeWm+rVICFukqb7mjmuUdEfekh6
piD3IdLGdfdRq3bnvh/FYD33PL2JuVyzgLQGeAe/WTYxLwuw0FEJGNfgkAoFRoYG
/5K6c5h6izVm1JrPzBnmdRkKcpKek5Yjkv8+r++6oor8wziRKqg3kJYxCRWaSi0n
FSjKQfNCAP95dPvvJsKz/6nzZariD7PSV5ZAcNK6u1kzMNWVSIotT0CX2GGGMk5O
NqlYAPzMI2OZYxsYMYlbjQ+U/6aL+E33Hd+kimMrl3sVhY5B7DSTObMWwN17MdNo
ntR+mwtPB+ksxQLJ0OhI839s+j5dyNZYo1mPwgFjNxuOd4m/MWv5tbHz7PZVatpZ
lkPAJkUge19jZacivjRJ/BaGYqWd3T6MFeG9I18WbGtHl6xNPwh/eQ1gVdiNsVGE
DbBrRMH3lOX2LBl/k7hpEAb8e13zlXAwKXkBm1bmL8C42wmoOhuEfzC34tUiY38K
glyXGsLrgmwbfIL61ecsI9CtgmAOMq0CxrbaW3QMC+kakg1dfIXuMvM2XykVmvbf
eHN6ckUyfkCDiO1YiVUEhtyc8JYX7dJz3+QrivF6gX0fysb1xxul4FyAXAovqjlJ
6qeF6xOD7u2IsE8aXDDV/JG6xsQam+paSSW2VuN5WkA6VTOsUz1BQy8Ecdw3hMAZ
TulO6FoJ6gfSqMaiYTKuV5keXTT7NaNMdXcKiFMtP0gtcLjVJSxIuxIDYywk+fs7
tJfOjS9akDbetFHu/ar86pjH2du8PBsfRrrSnnIolYQN3l9YLdcUjROKl5AejkMC
X2aL2eYlzmL4fSUxYJVqbKoY4ovhe5f3wCAX3sAmdWtSezQgCOYLSx354bz4Pr31
8c9HXTZrneay1bPQ5FrZJToZWBb0JTDMy4Ef8yEIMWiXAeLiTnqsZqlgj3Kjjj4q
kbXezn8G3NosG3vCmy60hSibbFtMOfuXq5ZcMEvitIgzX53dXXpWOyUmFQBpAEbe
QLwZkyalwZyFY8lxhUHtQNog02BWHv9tOGRk1F+hdgjXXbL2sH0nlKKgNL/pe9qR
024SHiUtXY8Bf6NW48P0JX4vCZo+Z0KZLbCd1A0tHPUROu6iqJ3hB1sL0Sld7l/A
0jyhUKdRZLkYS+AYdY2+EyVetLfVHQYyUOr2UzwnXn1Y3D2Zc1upvCQgIY9Skz6y
NnFCTMj9bcOhVq6UCnLJMgtYMhTPPEV+a3uytOSsMYL7nNe/QPfKJU0TvZy/Tq2Y
wZLwS1I7Q1bf52GnuRjU2jVU/Y4kXmmk1qmnkkH+BLofbjhFXo2TxXG76Cdp8Zuv
HU7ctZtEMTqzzJy3S6k/gqwJICwpzhBYyecd0Zpp1jMdgWUtYjd2CQ/OTHFEJa1j
j9NbNeHhdeFEOqmRJDw8646OxCXaB9IJxoZ5AB1B4f34rzTVE/CcyU7FZs29BaDz
Let/cjNV4kp+XAUouA3b1v0w/kdoOJrkJdNDsIIURCr1RIHwBKv7C+5zvQdrspne
`protect END_PROTECTED
