`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zUzHH4Owei1eY+/kFWHXOK/cueGmD7pGNjT1j7eTH/Z4GkxIUnd70+D/1sh1v/5v
+5nrwmV/nCkJ9eezKCXLVawmn5T/Rxp+8ZhjbW8ikfi8jQ21VzqKwioYqotA6OoZ
m13t4Bw4cZZAFcpJFp7mu4gHx28sE3KFboQLdKHeg0PgO8X7pIqGNlo8uMGqav6g
lsVuBhr//b1y6EfxD2MUEikPFAyprxiG0a6jczbojWUfWZacTGdCzR7nZLe8Ozgc
9e8K8rcwFLNxk6jC2/xBLnCc7TAdp0Eo5q11J8Lub38o95ajRc4djR0Itu/pbpiI
rzaicq2fFHC8LRBFYliqDCcmZ3GYdcMHaV2+Anef25TBfuNf3iKb/3IaIA9TrgW2
yuLlbn7tUBU5Aj9lkIk9KR5ENG8ypxy0h59vQtXiIlH39ZxW+hxgx+FQVcJESiIJ
`protect END_PROTECTED
