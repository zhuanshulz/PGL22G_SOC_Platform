`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YCztfYigABy3pNtCXHm0zgldCaFY4YxHVqkenaw+HK96LuTVb8T2IowqYajdxUZQ
qL+ru9IDVbvwlYQVjSb2jzPaMzY/9tzIZl2tPBZ1YT5PvMeWWDxgvpK4smlwLjBg
+ivFE6x00+Vg0bZG00pFlz0VoLbwzdhx1uSA1WKdaD2oboaqEGu9HaWBUrOCzV7v
UXC7wSH9qKBQCVim1HYqVp9BQOFm9NC3CdqmAOeWbaaTMZiFAscc2348ohFDJqAV
Fgzw4T4kK2qZlmtkgWB9+5QIu9raEbfU+Ghyz5hjd60BKLgzgjL1KVLhRaTlFZ5l
NfVjLDb1blHbJP08lelT3slqlwoQCjV1MT5khZqE2rSFqquOmBDZ4Cfd2fmGv8bt
GSR03z/SNFi8l9Q9tamwPPeC8i6KOTWO09MM2iI3vs4O2GyOVwC/HJ2zxxLQceRM
fL7Y05lFNE/hxMxVWmXo/DBopea7p7a15zhK3pJyyxL/CE/t68d1TgULcH2jZr0z
aZTMC9MeV87PyY0E4LPAnBVRjxOZzdzvAm2WJVD+jI0x+xq6zUNk5AYevxJhWw3M
VOS5n5uL6wuyU0ScEYZ6v3LgxuXJUhmYa32guFM5tXY7W3Q4eXlxSsNoWiQun5yK
yB5MzY0LbKD8gTgDwc0Glox75uzP+5cK8vDN1HZdtU/r9RnD/iWrwZKKaFOmZU02
qokDn4cM7M5rcEA77AcYdv33UOAb3MTIIMJFwFy0Se6PKy/Wj5QyuwNQigPx2eLh
TBBT6eiC1GBvUARkM8k65jvQuyE9h6TC2MtNcagtKv/oXdzxe9ZotlPzxwtxi7WF
xizy6+LcbELJWBPamu0Lsw==
`protect END_PROTECTED
