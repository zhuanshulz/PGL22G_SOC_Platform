`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
28+4P+HaRQLYX650AKY73POm3PwcXcreNK2VfsZex54tqvezS0XZ2brLBq63m74b
wZw/gIuS520P5GhgN+wOiFOdKGVWO19+6GS/t+8pK+wvhAdstHgHB+brlRtL0IFR
ZU/jUG07HBn3fnyWGegY3w4dI4zwPLXrrjtqu5fvFmQl/NkITmlv1PcMf6/GQEZt
5+6pwA+uVYLymBPjbJguwwaRpEKFpxoTC3R5a9J4jaWUojk1u38wsH7fPIG8Wp2A
z3U8DoI6l8ZvGd+zE9nnIGCVWHgMqx/lGWvxFK7+YkP1JuI1DcIJTDyGubXwboyk
R+f73YQvtNi+BmU71dNYn1TCSZGGw89wlDSHHiUtg6bfJhBxIRzv11HS2Ntq8HlM
l/Re1Hlb9Vs+KOb9EpN6/VKw46a4fInUtf7FT7YN5mlMmxdfzvh2/8sMmpMSss+f
CETgCuR3kf1VSe2NXJ6pGH2WPC95o1Qq+nyvzS1JogdfIxI0LGhNTQ+nC4lZXetp
RXoussdMDWEWuPjr0m2cQZEMM0SyxXoO9SpuvEg//waXPCP1EBn0w9SeRRDkfshK
sLU7iXGIkwCnO/pFjEM8hYFmESSMpEQi6CpLMpBuLOu2qCphXqWrQdqVkbBFo3zg
q5GuWjZwudb5Z01I106pR7ePgZAUlg75jtKzNuQUd+wLq69WbVyBV6tZRHnyoFW3
7AUv1MN7mrhw5kEqmGmsmqMaC3gX3clCEi0qUo+IBgytdMLNZ9ElUG1jYy34/zHH
UBi2JKlYqf32SPcaE5T2/zYjoctTZ6XFRb19FjujbxeXhHLJpkB0eBgDlCp+4H34
gJwx6KLTxg0zfZN7zPkvHtD/gza5IUUSDsZPOb58sHhq59dlFvYpkB/NdPkgYLWn
dz7R0Nvu7pm4MmOjOW3FoCx5OEUmjftNI+/1SIkvlFLrBsDju2mUFkjuyV0iZXdh
n/wtBGyJwhw/1TWbXtIqVobrtaBvCOtRhqyRMqBP81NilS3vc5dp9Jq/KSeyKwKZ
myXCUxioEt5FUjK+tgXin3fGZcOvDApjMaZTSzNh6cjtIPgLTa2KERZDOPgvQr15
CmLxeA3G+EAVHHugQ6CSbymcK8xS1KIdg9KuAmYXcLawsGzckta8E9mk2TP+t2nE
pLnvC1MvjjVxO4WFMBbmpec0yMomD8GfUCOz7aqDMDzsrj4WNy2wHXfLp+mAWok2
QBhtIot7q7rha2C163cXIrWDMisNU48hxohie1YKzv8iAQXDWWlywXhvX7AzrTm/
v6YHyh+z5u3ZPeVNKmzDwqvpzcAhyS7/HnsRhsA350hJTOWm5QgxFJht6NAC85JT
Zyb8JveN1tHbHGspVmmWJdI8IdGCesnJM14PRRYDAe5ibrcGutFt21DygalhEnXu
65Du1+nZiZ1ueamwapbeZbpFKdhc4G/0+7ysIANLIZwqd5eD790lP3W0OcJHEf81
Frq7RoTPWS378zLH3BCms3tGanQ+aBKD4Vgle9O5OIRS8Q1qjXPv3NBk7M3FLgUH
4GFuI8/yudbWghakQkO1aPjiNqzJoR8R3fQdXghRzZTzKpkuq6q9BPP64jvtjYxN
24ZcMiFB78KWzFUZGzaIywV27ivigviucBRFd1rqFGOmu1kkNnIkjJK22ISkawPK
Ewpm+ZzFngHxevSqQH1B5zrTyY2nZfm0MHx8anNcXmjnHSD14Ffa3Vorp7zPfHuA
+gNMKsvqgkEk+8W5Ogkz+N+ywgQwlp3gmX7LqqBEQkkjpUWT+7OvLip7CASVZuIH
DzLeD2jnT2ixGa/gVzrF0EOOJ2iWQzgwTrvz0lfHw9ohBzPXWdh8ZQy8F3PcsBww
h9ElI2eaFw0vSZv1kAYb4y7eJFd+AA8Sth8I8g9cox7O/Q6cvQ8Ho90gTxGI8JQ1
L6m8Z16W2Mt6K73o2bKnPrNW6w3JUsdbB40VshmUMQK3zJpo5/iagTkPDJcZQfAb
FRDxPUzv3qZPlTp41BCc7fuEnE4StOB/3GU2ptfTtaSVQD/CnpOdftPxVYH8e2uL
V94I6KXNz8RCB0BbZPy+DLR/70DZ4Qtq0AZs02a8nPIaarrhD4LxLTYxXe+Mn0ws
t/2PahEXt7lt7ixKT70sqNDnIIehVhxCINST4ax24bXOdBTlYLNtMnGYsAQFIlcF
I8Q+5SqiL9Gbj4oNLyxgw43SNCGi/znhZJ8Mn/D2tdQ1A2niIxCg+T3GfCLIibCw
/sBcfoyZPsssCh++5EjMdvaI3f16FsDiP93rz42XxlbRtXKDHIGsfF/LxLUTTwN0
byPk41bJ3E8Cr2PExzqSF84yUg2rkuHkcsVzxBz1yxDOyJVpF1EORdjBr95yPaYg
7+BzpHV2ZzLnknhv2wnnl2d3+G4NvQM5G5sKfy1+dcb8ymrV8f8CPPr8+F6QjuPd
8yc/VpfumKHfmPrjznDcKMlgHWpyl3B/znx1Oa3pVPN+nhG/n+MjWLzYfpsQSe8G
UKIQ71/9Ilaf46kdahaHbG5BmajnQXCbow+jp40BcxsTFIOg8NEF3vehS1mr6jvo
XQU1DhutJbhqZDGK0XooLXE8cWcPzq9y+8H4hfpHLw2ZlZNhlRl1Jb8Z7uQwfK76
G3fwafA2npse5jRpcgQJx03kz0M/P+jbaTP1A5zVBPQ3a+toq598LdMvDy+sXLIx
naEATTdxh7Y0D+9zcsR8k4pFIH6IvXykg7UanJfDS+r5LDwJoTaafNsYpqqIgvu0
vrW9c+J7AP21Zf6Za2FyYSBK38PKWv3cK6WhWilTjEEF08MXAtCvtIYWiy8BTYSd
H4lwbuE9XyUjzjmKWmjhtv9kkWhCfUSEMSdYXXTe45yTYcD/tYgnYqRH2jPPd/1l
RrAwxdBEaktlIrplwtVSi9MKDBykjCt+p45s09XO7emDPifzEqr7QA7rAD4YwvRn
dWLlG4D/oAhme3+4+HAPiJat6kkx93bA9zv7Rtupp/HE4sTC9eGMDq+QE7uAEw+f
r1RjI8LPsPR0R9sBq7aCRFAT8QsIVwmptbRok2tiXJmHNAqFE9qENpO76I8+Kvz6
RaGMurOh14R7c1tlE0VtSC0+UXs3IOY+Z1eVCN82i6YyO8mkCtdyWJUtc6OJVGmT
4x9KJ6JJ0jtE37PRjFGq4zoOzAldPmglMVTWA0GUdNbC/lvWiHh9aKAowWzg+7A/
/GvA2ogSKydohaeo5drzPZ/W4qI69K+2f8bfRdW88uWpfYR7Eu0gvWsxRf9BwkpY
MYK/iP5hwrOuTIQW3qxOcMpQG3xFOtm/NN8BRHXGFeCFwRUBGmk0hZQV8Hi0l1vU
KS7n74rFPscIv538FpVRiz/RCGQdGHg3Ub9M2liEg+ilJ3S9ECx3Mc+h8Qn0v4Pe
VZvI+e+bwvRwA3a8+cWSRiOXHrTmyBdIwQp9fHTtXM2j1RBGvN6Gu1u9/zK4yGLU
DYRbt+L03OPNgZ1g+dehKBxQT+DagF8X2cJ6ig67SSr4el8zrawsy2dkFW5MFLKE
Mk4PjYgHKGQ7n9o81JRmTJeh6Zh5Zw5FkjM6mlHMHayNTMc9sebM8QkerQC6TunI
tpmSNbsgYmZq2EGK0qd0SKBvx+Cos1hbN2AMlIK4NcmM0RtNPmgjx3/ZyKb5z+05
lEe9ezRcR2TbHu+PQ41R2ejp6ClsABpCwLVQskm0ZfqUFBFhzgtAEEZMMoHmeeqH
FrDXq30lYJygF67FlikonFb+wQaLhu5F01JPVaUkGgLsRz5a4Jm/M0SKVshHefF2
oPaVyrM1ujtFp2YNNoo/E5IHnerIjsIA2IkxGqqLX4tL1uF5bFoDXaXxod75fjuH
A1nEZX2j5jLYYjedyV9Vp0v7Tt1W/Ex6/fbUOXzOUV47UM7YSbgGJlqbQdjnPUf9
WdbPPspY4PfQAboP2FPYfSK7yu9267Ymk0EJXNBPB4ftFfO/1Qd/V/dHAFhn4OJN
3xRktjDIj316kd0UM58ocQslA140y9izsP2d077QBa2ukmidek9JTGUHa3xR83xs
4O8cYIqyANHS2BGcwwITFHMthfsCWDzffmWIHHPlrTBRoU/RxGw403wboQcU9T58
xjuJ+rW2QO7V1gU3DNmWNdgEgzH6d6Wcwvv1n2zFEDPanNF6ZI3VSGt/OrP74Kfr
FMM7y5x4u4zwbkLrumsQ0JaP36lO+bNnDa/tHoiiro3mkQCDOWBWozr4FFc/N5do
8VqshmpV4NhzLJXtR1bq2MfhvGldveZsPvlyHYuaFbi9NBmERfqmoBLYRARwlAU7
9xzJEhN47Cpp6oTw2tGy+MxrP9VZoDxAdKmrD57KUb46La7x9+JyZ11dTShzA1xI
dG0Oizvzp7B0Dm76qao4ma28ynYUWZpp/6y3Re94z079GW3rFU5M3Uv3RPogz1T8
CPnBTPs5U8N3udd11F9Ukz6KM+2dP1MpvKWqrGMbH3zsbCvlMtrtrNrerP7r0KMy
3u0fVsx6ezmwx3M5WJ52EYQHnt/Ul9e+PO3xyWkRuHVSU/2eHyx8qjZUztaiciFS
4Porm8X64qkao0vSAHkqf3ZHQWEkmtsilJ0Oh5jVQoFOtdcnyd80NnoF21LO2i0u
00YS5iIM70e1muTEvS+ZtmUCDvAx3boiwXCvu+VBls+2ZngsIuxHepxG0t2ykBWh
K+bZAnIYtQvBfDeb9nqoGM6gbi8GZuowc65VkUvZ0pebpuU+0WwtViWYRDZKzGA2
gVToThDjiOKOQMMASxq5RmLzQvVbjshyx9BRJBGMEZwT4jd0wKvMAqQJau1jQhIN
t9PhUO0HqMDXnCyevrWjhF+pp5bklzASn7TNeXlWzomcxTuR3KAsTnwV4S4MvWrm
LlnMKnpu1X1fKGPy6V1OjoszhGJ0/hv+XLjbSck5IGyQnR/DuRII+rd3aVXlMZ66
DXIbYjtiuzLKqBgTaIp2gt8/CyXuDBFRmwugboFakeFOpaIWN3SCIN4+wHw7xRhD
Zm5wz1qGNNjBUrsomy4ktS22Bmimf5mPmeVsU3W3Awm6fiz3UpxOHSMv07DcmMu1
/MOL3zw89A6crlLgcZ0o+tuQgOCJJrJmEtLbENXk5gkQVhklWJlc2KmXkX3k3gUO
yeMlXJWQ4nCupxK2W17QmgusX+2G+Yj2zDb/Y7dOL8WiCbSsXBXcKLMLYMuCzgQl
0RhYbvpt8xM/JVGElMYLRLz+lcUeaun4/+Te53EgTZC/wFQSYSjLB56DAqHrmru1
uSnM1BJ4zs19txPymhUkdVIzIOvCu+p+QP9UMhFDMosOzjFINXDSZUXltTYn1nNo
RmcP+pU+ZitM/YkwhXMzuhg6wSTX3F386TGnFQFeZWLS4O8ZnKdI3u/ut1jQLBdd
a/Y2Glj0raWRqOFFkMbct7WF9Jf0JCXyTXSfIq42iqRBUZrVosV062nxNKcLEKTV
JYPHOC/RSwcFX3LhQxAkykhhxMMsn+o8WYUTLr4gzXvlQiEoMVc0+wFI69KoXjx3
WgI8/wLHR4LoUPS8oOITaCXLV1XbS1smVl32NhzeZSXkq8VnBLAcyLiIHZijoLRH
0TzrpDLa0rwL3/oOaQTL0la9BPQPAbH/VFHfg9n+KmYpN9gyl9YkURdrJDu9ArXB
LYs3RyNsCp/lXfXQRB6u0/LL4aJ5n4YxIyDJheoODWuKl8doC6MyYe62O7AaxkQl
YBRBceftWdSlaXCGwQgzG9HlmM7NEqdLfhZHO6OK6n0mkkA70fdEr/keaKdyuhlF
GKOZHRtgfOV/wdc/+TuRtDKpP4kxGSenqxADEGqjHqzKybdr+J8/dMuRSIxHpOZq
5xvYDmbHiWWVMXz966Tt1osr8CA8YCWh3wD1NZAq2UjJjozh143ucm9v6HLKaqD5
OKMN7IFjxbAqlf++JPjg5GituTxX3my6DnvyOlv8M/Kgb9kEr3B+ohpKxCPpt15H
+/fvaoXtHYj+TRYkzHIrLonvLS9c7ZNXYuVmD0ZhJe6xUQ9V/sdeFIoVxdlCuqYX
af0xvI0+yw7Vklzu6mfhvoFLDfTuSYSi24QU+gODaDQB7dDTdN+EZ/PWPTOGdOQY
XLHtpNmXq2pN5s1/bipo0yBI4aDvPUJl7NdsUyMsojg969cv606qkyvdCwH+blNi
ZjVUSv6zDdBeWvzBGMhA1nNKe8dDGMfScbn+JP3cNwcmlAMr2oWtfoC5kMb+B0gH
xsF5jEQMUs9UR8DymSsj1m3vEhuNTgko53gqpfNmbhNTG5Pt5u2mFc6tz3sx/JGP
FtdmNtRQYUP1J0PEWdtUfvy07qKj5qMwQb/pYuQHhx2ByKF1pJmbzSUUOvHYtg6j
j55drjJfn9bjQY2yncF2lvszauu2z238c+SUvdxDuUumLHTwyG3wNpxkz4XB/mQB
qLw4OhAsXPA4Hm4y7y0LSNqqFwbsQVP6aZJAkI6jQ2nG7Zwu7AzjmHL+EIQ9lfQ9
1unhAejsu5JbX3PVMjJJpITSxaePJl8bQ30w/4sAv3rFPDIVt+jEPzHOTY6tv0Vt
UIWpg3vgRZFykFwBKM5Of9KdZ6gFELody67uAgzf4U1wz2qUf+8keiv8OajwF9iI
ni2J8YEOtuAqKmXNOIdz+q0hZptGJtPIx114Zuu1a/rcpPFbLJ0Sgd2KqDQKk/UF
LTqwKl0ANyZwH7UoVHijMH53HO8GQ06EKzuDPIRVlcgHSSzQYLkrI3ubZdxwNq9u
v9dNvSLQlNxnZpIsI5ZWJqQ2qihkKpGQGqWcyisJt2E5pE84EysP8ME30aVUwOTa
B8RP/e6rKk9ilpuw0/WKuWltuGTmIQ+37UTGC7edCDZmHK7HXdI0Oogh+irlZ0IC
E1GXtPIst6ChzFJAoPMpLWNGAGseY7TeZoEdHyTp7+M2qa4JQZxvoLwLc1PD0GPg
Funo7d5HygpM5gY33MmslUZfoTZYUhTV/J6CoD8EJe81wPmzX4CNzbWI43U7BnRl
O3YGz7D/TVeip9ECHseUelvgmzcziHBUYDNcV8SN1MFLItwi6cSrNBH57sVSMXuL
cD01O3r1JqLCe2Fxdw6TmtrVJccvocGi5jI23Ge0DaW/OaHxspU4Hgbo5D6YMY4S
jBHRDfKpawsuBjJJNax24ZGQjxBW+CceKlZob9RWaQ1560vUPotePu0UeWcqAU0Q
nUf+RuNqOQGgxXzKiu6GVDR1XkARzkoT9k/CBLfpBtMP/xZs+NYUq0leEc79f6hq
EEiovJuLlHE4jtdALx0iyUm70emWCaSxarGWYTAwEDlD3/oV7Jwbml5RBJQzLjQH
klHxUBAHGoIOQ7JKKCIR93Jt9pPLwu41KD13dfDmzya5NRI9HwYSPalYFUfYQNeg
cKdAnPrDFkHjCjkAgcGxnmslwHyqCIVV92NbTa7uSDavf10ff7I3gw6bBd9ut9zw
AwO3EwZBbHn7sBovCC+iV2lPisHDUa1VLiEQ0CI9prJGnFI1XGtzuJ1+FRHUzr1l
qb9OnA7f5Y2ZAWT9bnZR/Gc1ceWRL+fW06Ka6tJt2ryJiGsaBvnk/3S34cydqVDC
WxmG/2dzsMQsibLo/+rXfjhf8iGuF32oGsujhWNOzKMgexyGd2NGk4wLZQvNy28P
xbJ6NUYwqsu7QjHXaXtQGHMVmMMcc1kD+1kFjSC3jxUwdHYQC5bif9cn99qWWIEP
N/8GdrCLcQTjYBt07LeLHlXkrya280qzHn6bRVBggFdhe/0MSWZQRv/tp+LOUm/7
3w8umRW4hEljT68bVN5mTbx41I7ndAGPT/YDDJSm+WXaOYg2R8zBzu6Y59ykqPcq
QseofgoKUWHcpZxAvmY1xjn+weYB42CuaMAXUDkzPFcOYyof9gz3OLNkijExBSIy
NFCK7DKUm/iYU1FaP2+0DF4hyfpluw6Okam3kDi5reaYnRg2n19/kWugzn+ju/o9
qL9cubRXPZLA2BRXLtH3osmgMFukUsgtCEvkZH3PUyIEcyVgbN+8inTksmRfUAfo
d1rdhYsPCa78j+cc7zVqXCDF7wLBzSIwqDQLMnAAmO74SbywZmEwkrcmZzYPQVYt
u0f8zP6HprH/H9hzpmxQVNkjgF/QKcx/nJu8+XqlhB+PlBaG0oeBxXorj6A6YHlU
kE3f2Dc4/75KTt70WH2gs/KRTpuWERAwPBZKTcME1GDBBoEBQk84rL/XVyHVK8Jb
s2jJHEvrSfnJvaXu/exHYORyaMEFhClGV/UA3gJIz8Ek4AK+MmFsTe0mUP/OKmgx
is7cPk3gZC5x0AuecQySuTifiiUgiD4YEmLilVdA2NV9RZMYgAvIzyHDTWQpjdzc
FLAl45mPcipgKgo9R/GT09Ewks4LOMJbxH06E9AvTsnw8/2SxLObei+NeXP5Y+cW
AkpGp61qmwMw90mm6iCidKAZP0KoUazM8vOPws45yyB3czoNWSZzvM1mZ9crh9nZ
2iHVNbiMLBfG8ih9FX0d2kq1CPyim8N8FQCVuxreZbp9Y7BYyzvh2tvRAS/sAvr+
AG2OAdvWQKrDDsg+lRf8Td9aW9m24vh856ofPrGR7r3LaIklAiigN+ddQT1we9jk
CD8ZIJSIt/yEqQUfg23AJFUyDvghRkm6rR8WEwmOWq0j1wE2khlJxPMlQWMV4Rla
XsgpEQqpdVe1a6tXTrb5VonfMF6lWmG6bf5e6SIO43WgWKD2L717Iv+XTNlGxSIp
gzXFdb5Dwgtu9jWhHIM1/lltU0m8cB8RFW+W4VzHCfpyfxFm2jEkav3aCZauZMD/
T80z/K57eymbcWEdFlJomxFB/UACHME0yBkLNWkqqpy4m47xXlSzMbOhhV3YC360
fVQgswpRht5Dvwis9bStXxpmQDiYCJusAqLkZUTu7UPlYSHO8ZheiDXcSsRnWhPB
3bj8vqvqc3zmzhyDs1H6YfX+LkrRVMN7rgoPhC3LtDbKF9nOFwV5p3rAgHoCwK+l
VjKDfCmjyPuy3V+ZcbT10EKXW4CseKTAigorBDp8MdLy2LDUud5i77S6Y9QCP1pL
oNmy0dFh1dRVL0hbrSV8mAouWDTD2PsntSDWuv//ZMHfierMBZw/7s3x9e3euzq2
8OU9+Hx0DFGVTZ0VEF+Pbvc0tEXpquqYVo/5rXzjC3GAiYPsuKJ8oCga6dfd838G
f1LWJss63KoqMnKDUU4KoX2S+tMAMT0OTyRDJyAcU0KWtQyholVoTht/QYwI9wuw
topmNxhcUfn6ROJ+9GFe+mVxzXPQ6VYZf/iXJomeDuhVYF0ZKJWCohJf27CG/A0M
wAoSTAtBfyKxrNLk3CdpUaYHTAJkaC5SwjcHxSLdVpxc0W0z4jCIuPvlA22L1wGA
gks7FNsGjGuySL2FmW/3L1yjdS0HG/NttsgXE11GCNQvMXCq+934F6jLj9oxzE0G
XOHhZdsmtz4kQMUG/BLEVuq5GealI+4JZB7oOZZzpNlxL6oNlok/sbMs3/M46KqZ
fKUhq8QE2tUn0L2tX7/kIKmWwU/vGItjQ0/4bsU8/Sw+q9bmWugv0EWxmnBDyCdY
C0cgV9yU8TFKNmtUwDesl+7HzKkjNZ+KBvleRHxgYasW0a0nWwZS2Y7PLftZJjX5
GGLHwmdSE/xodnDidIxdo8ujRt+R1XuRu9DJ33hbFvtedQcrUf4mbY7RpgHScQaO
NTUciq7bripKqeQyeWoiPttTJo/CeR36TbZy85scieZeYduIG0shO8YhIudlsiYH
fZSFTXnMbAfvDMa7/A1ZSW4MR1nVn43UgTapdA2DeEoVet0JuMJjajSq3vhfqn37
yVEC55mqowHaMg4AuUY8tNbh0WVqXORkJA+NhzlH9S7qfbtq9gnRiMmxtOmdBFZq
FRRheIWVbplJjddq2Rfphk8EZXqJuEbjNU/Q3E4wHKxxHvnk53SgXA6tFQK/oQxf
LrZq27XjMU4bXCCbjzgjLhXXX9JSi6Bo1nA5ueopN1AisgaUjqBYA+oeGbUVXtGr
bGN11CWPzPksuZFaUlVP8f0kbHhGIulMLQU+CCbaut1ShBtQBj1QkD+1XhYASshg
zb9bDKRiOwZ2l0qrw3/36stB2+Lob0ktq2wrQLrZu0eC99JtcIcnfjjh1yYHQs2z
Vzp08WEBotfIVZ9eb4bQYY1Gp6imX3O7/BznX3SuK/HXG5LTc4tYjYof86Lh9j1x
rCpWd8Ei7nk4qCByhE1Jqa2JmwEXuBq9qHLQmYh1kcIGmo6ZjC5HddkWi/k7xvSc
Xb1KM/NrAbvwFLrAWq7rYcqMhzr9jtJcjS6oBfTaAcF1ijQ4o2NjDZwtD0jw1XSr
ZEBl8K/PiOPKRJkBqUSQcRoKikeVQJ/NOPZ48R22Euk+56ng0B1B6Zat6sQOMAA4
HjhYkjJqWx/tz+VHKtE/3U6w69iFkwLJMqSezWllzAdcsIh2PASl6kh0EL75sSjT
5AJI/2LZV27mWDBPsN7m4DcXrhD7g7JPat7p4YkCe4PWhIZYX5oQpq+EZI90kBJb
0fPKKtbMqiqCqdAX4NPvzhTuULp+YwE699QBfNfAJxTQIfP2wI0h5evSvXb+ratw
cssvkge3wrBhqGSw3nHRSdyWK6pTVmgYGmxSS2tBkcQCNITwoMwvkTmBMhnb+kbM
EI2bheG06vYBj4KrtEnqTmLf73tw46bWx5ONCTy3dQYnxOBW7qfACuvs2xUNQXvu
uri0j2MZt49/VTCGMXMnYUt8c+Q6Hwih42TOQ67rIZd83ESOom3e710X1ZhJB1sP
z1tn5Ke/ijK/G7oRBkCjtcitbMpwSiuyhUmCar1exzOgvTtQr2IZ6NHj+3bkxKy0
Wzo2LlAolDx+n/Q3M5kPKH1FGcaZvvMtJBLX2bxVUhKaf0ekk8OWOkSG4Yg23mNE
sQHTxdmkFQo90lYRwSWss92B5WQ0naur5uoYtE9h/arx2VNC9XfTIazlFAvWgXwh
4aSEdPS4969LG2SkWcByxxwR4tUDy27qGIHXu2hbaWtANdNMGjCDME84jSoeoOie
xE+T0qrGo9mFtCxsVEYLeurkUe8znVuH6bVqExGU6BhhnbGZubgGpSedIZs7vnaF
dN3eW/TTnlyHvtP0rGuBO8rFY6hRbXmTvFGPFBxy3LLuwNxrhdBMEz6azrcM3KCM
PpJIg3yF2Gi2vx+EIJfU60NKkVXccGTqRv5zO5/vRzgAOrwBvaATH5JkURwPwY07
0LWfMPKRGENvgQzU2OZHybeRrbUq7+ZXAbEAVKrfSEITFV8YYdRF7Y4Iuz6Uz0ho
2W+4BMk9m7zUXnz2mp4qDgx2KP04lBywbhXf2CD9WIOzby8JtgNjHG7t0e/rBbHd
S0yY9FjKwfbrb2chOTmLJQWThX1eCUGZr6gGA4Mg8zlsuuGiYgbfHEpuYK13ZAUV
1rlA/8Grls6IPF9TZqWUcRUvc3ymffPfudP8RmSRUynK5fzX6aSi+f4eTV9ab5iB
tDYmfkyr1qhOdVX97Pe173sCVrSaSMmumScVppXSZBzZ/IBn4LsPcS6gTequgLN4
Upeor6OqUgfwfuS7zAAAPKkBpCqX5gSR3e4XuO3AuXzwKRktUwxUMjquAPHjMJ+Z
FHs0lWxE6BeS++REoL2M5ekPc90kibJll1nJkCuz7icw9aGoCOgJ7puYXkneEgcG
TMDM7ZIssjrReXhMbT+V1m99k29KeU6E9NIURmMcRYL9kNZ9vBUOrWwmgMb2QwOY
Dh+BcmocL0AjUl9Al0aYDo95KcBbbo1JbG0VBjbSJJuFfQ9OvtEayk2X23aRyyRm
SfWQi0UrV0Q2jwxI45utR/WduwQQjHZgzdb0h0HT3SWGOWXzrzCJOdr1+lMfujq5
vRlwNDxdg5HbivQdos2W3V6H4R/q/RY8/WcHks3If0FaOqBoSkN60kGMnRYhB+Gr
/uzU6gN2f+K5M3i05ieV3dpL1+vlvn0Cqf5s7tVav+BOQ5jecYRXRz/eIB5vrHe2
DX6ROkaPEPnWRREIKurskK17jgTmSP6vl15Tl83BLoU6TOZmB2SPEP7bRiV0h8aH
0qqrx32ne4h3Bj9wUa6Ch87C1W70RkkLeqXEbUyORcbEVo3aokEbWjYjWLnX761O
X+OA+xc72e4bpgfeMan78ktekhnVOOurAYzakYRF6dU02eXoAQktUsUZFyl5kvnM
T8K2RThlhwhDGOVc1zBd3sh2a1OXN/PQbxtMhBieouE+2uUPx7r/b6QOsEf/9hiZ
CqBk98ZpgCJiswFBqcIJ+pBdDFSYgNTR6q0XVL8YPQeQWSFmyeGBOSerdK8bz10r
0nX5c+FHwh2cBO2wfd/Q75o+yM9Hw3k2UScxTXnGUe154ne95CwddTLEG4+ds3GS
/a6zZH8VtC1lzV+avgVaovJ06WoONkjGTRCh1KI/uYLglR14kVdgCEk7MPx8rTox
WMdhbqcqLvQ8vBh8JXkCrBqK1SY4VDJGFekG6vdGKEnoL1yyAi91MfEBcB94Ozet
K7/6/wSVs5UXBBsolLxB0MiIJsWifv/F6nt3IIt31U3oAXEq0HRTWO7g+yVn8Qt4
R2aXY6MnyHipoCw46JtTjqK0AzB7Ers5HcWmM+/TfblnGrx6wY7YlffvjDhOHpk+
p08A9S1OstGBuTtO7kKdNhQRTeFaarRllKm4SoLyIOx5FMEmf+i4fPZVLfy3wTcl
Y8gmS2IFRPZb+yHiaaBxNJHr3Po+xcsVpxhWMQyCSrLKdQEE4sc3XLoTILs2fbkK
zpOK1Doq1PeTeTOmu5JI5Npl6gXMI8UeAmCfrX7ZkYENkAT68rd54inVpVJqPfQM
X9ihvgfpEG1hjyxEtAq3ss8dR84iGuH2RWIB4lT7uI5ndZ91/i2gFHYg4FdoGSn8
4OJmnaEyu2cpajX6JUv3IWCJpZt7Qqnlh4ZTztRRMVWPwR2/5BtjqKvH/a11Z5zO
pVR4vEqaqVUCCpaGbcyyaCsI1TzYzHPsohNjTGlOUKWaPJPxKw5m1BgqausRZQWD
obriKKM8PxMN76j6pKYB+GctifJGO5emCPfvcy80SX2C+TCFiQc6ZsXF2ShwcCh+
CfbynQJwibG7LHIi9Q/g8NCCipN2mOhTg7nwmX/WadAsrzUQEcHBAzNpLeN0Y91T
U/1LL2Y53oJK3+ICJ3NyHV57oFV8PsxItZuZE7iXNncotx6VckCTxzRIvStuO33J
5riq7BYMNEV9usAs+EwFPmuH9kW1PVfJiAj5jCWhPVMaFazrYiNTqrlAkgcfKoYC
+J+s8k1zVl5c0c3r642F0+im6MCPYmPRHxpt2tVHRk7kADVHmrHZ18gZVyf5h+aB
tvOGUHoUW07Bl9fl1mu7is1OzYeJUx0VW+LQqheEDbRp6DHszK+DKEDMeCDecGPT
yNPXVDquNX7r+pZvfhA3XvOVghsq8zXDjgZnZNjNuqmVnRe2914LjvL47tvoIUvn
C0HY3RmSE90dP3nqoriPUipDAQCRAbdAAnvSa7TfmeoPg35dM8rNXbBZD92xUYel
K+6abq36Z5m27XETuC/lueOldq3ucYsD2PVXGdo66Q5bbwbUEcHmEEFIhJ+mi8wA
oU/AVKs1H6O5KIhMTSx+fDk5/jNNoaYYGor+e0/bUgHSWBMgzlQ3shoHaX3tL3Vk
IShPhhr3Pxcx9JXv4idtiYqUXL+ya3SYvGPcDn5CMHrgeMRPIwfIcaj4zWJC6jlD
Xguldnh/Pr9f1Eqt5OS+sKfHwl5kAjKFe3kNJ1l/Ccfod0HGma2xwgkZXYaxspZx
rYqCX9TXT8h1lhPOqNnCoTIgEkPch0nbDZqZN48wXQIMbTozqfZ8nVeGMMKZIVP9
o1dPe1UQBs8udhGrJUq+GAGSVpoDAprDCeRqen7b6dBAUosnhLmxPA9Il7LDDerk
meFaRb82kdSyjPlBQVpgpUOplS6Ox3MlJhiU+l2D0B66qgC8VBVeMHLryUerlA1S
ZjWjS3Usgx0NCdBlntw9mlE2gkmZOSfDxxbaWLebef7m/q6uhHRArkU+OAGq05A8
zZQXrSSezymxAFzCo+KLXxpUeLh6k3GohGu+FRWA851t3r+qzetc47M/jYkwWJOP
i/l5NQIcbzfTjLxrRJ+7JhBEOiM470ynnP+IBCZwNKyYptZbOjNOKfy+TKfOCwuL
XFqY/G2hHKR8oEipTEX5U5ywjOZqRrNAfSNyrFN8S11gdUdVIa66LGYu1w2aZp0Y
ufJ/DtBiNdHLNoFLowcwswobpBVYrVvoznbgF+YRfTOIl8t3SjkiPSEStmhN92Si
BRNOcX3VzBWfQLDgjFdKrmhlJZcClE/VzEvfb+LksfSpnfbB+pMBaz2Vvi0LoxDh
Rc0ml122JRb2dX3WFt9Q27y4on5hXB9kBZ24TX4xON+QqbvoGyWV+jKOB/ScrZm+
V1rRFJ3UNKZ2FhcJLb+yvQd3c6Q0CxATFf0DMdzlwL3HQ6vxTtrh9QqvkvytrBVG
lZvZRIG9xUobpGgvkqfwdhRXSsZO1KUhQoyEvD41LsR/Zf6aioBROAbcnysjQrxc
7VWvPEPKjISj1UEtucF3fuVHpGpWM7c27Q8T/JOK6OpguPkFc6IsbZHnF/JhzQo0
GYKcktM8VyrqD5AibQWt1YLJ8arVQdlwWQUefKD7pv9gGWQmB+HHb9xi2wr4elo2
QaFC+mBteLEZxrT21euJVnVNpuZbrhdOHYNB4wdjB6l08zy1fnqCFwAwu6Djgnlc
qGjvq/qsH4i+qLsGGkArYPJ03i2sR4ApVy7sjFzgVK93mL18BUPKAeyHiGjtItCI
/5BSypHgNOnLx2xmO+UmTkPf+FmjErDuWk4FYjVp8fKXMjrLoHC+h4xDX0qlN5HP
MAaVNRuDTbDcDapxf0hm0z65gKe+cpriuDrzZ2D7K1w5mqMN9qphOaTN4haGxfYa
olOpElPlEXWUZPo0VXEC3P8aHV8a3Rt9T0anWT6xjR6EyDrzaUUEjLSpLzwCpM6X
hcsx8FUyoeQb+xrgElCi6NLN9ElHKv+eOCf+jPTqjmTUUO7BOzPwMMFEIbxxFuf7
gNyzsBZR/9vtT8PKdLUS2BfDcb7s99ewWI1U+EzFdFw5pLOrpSchSmNcFQUXcmIc
97XUIXv8vByIm1RVLNnd4M1lg2GBvt1z7xiLYf1gSZiabNt5lnYGwXSSjvPWUKIN
Z50iGOYDtSDqyHWyMgMDDh5WUSQlTgV8dHShp0o460/AuVLExrLK/aDdmEjlwbIc
7swNBDYOV2dvYfhdi4TdMFKqVPP3B/fbPZKLRpPhsi6lwo9YCrxPMIr5cj304wOF
+d9wpVmMh7Jj06c8x8CAjzHzxsBGmWkoqWT2PiSAbj510lpwbP+Ip05C/v8nv9Wi
On1HJVGJnyW5mFaP6sAKNMq5Har8gpDhcBh64eaYaGdYsDpXhXKZlXmzQG7ltTS5
QWhate1lhB8Wch6pK1DsvMuKj81vyl0V++vjYUVpmWK15vlFXryjAXkZdACaCq+2
RydgpEJ1QhD9SxMw6lbGQrCqw/g8egV6y0Hn8/ZQFNetuTU+qzAEk3J1cRcP3YAU
6hOCsQUmoZusQvZyUjao2RTLPRu5iOVpkS1nwKNeWASZTqZDHqDVX0yR578Sh64C
gvUvIRxrFUt05JWmrX7iJIEgoupdZrqsTxyNAvKB23iQsDYIyQYVi51PBYTsQH3X
C371NeYWakBScw2uO7K1a3gs9p1/7g4zejbeX58RtJLkhjyRAXmtKDROLnmm5WKb
y72lB8/UX60XH/sPgJYQR/mVvPeaxOq78+/VXny0pOVgRCp8De8tv0xqwxBE5pHY
M8zlng/xT9IuRliS24glkCI2O4h1hJfZcLuattuwu9lKU7BpCXdiOco8HB2jGz8t
J7MXe42esrU1pHwA7Tjx8pfkiMCuGOY92P3PUZ26k9bkkOHK8aDnlPPDwzkRtucr
Hrgvvd8X5Ubfzs0LjAtJKaEiLYsor3FBjbEKrmdLLoDuEULoJEADavwleZgzpwqO
6X2gdPLaSfrlFugBL5vcP2T4Gr0ajCrjZMkWX1GvCUkPF5u6jF5xK84lGfiV3khS
5aJYJvmJTkSLoD8PDDTv6vc9CJ8SSU7MkCAmh4uhRa5/IQ+iaGuVt1o7E1XQq/YH
zbfYcdlC03VlzF+BcnqOBWXOYehQU1dRk/ypUV5yx3flQNgcPRoXNH40XNPnCPR5
eEMETi0vKVdMENWsj/Jv+vUV73Lt7ovxsh5586IgyfqgBWEhUS1F/JTvQtF9R6/v
xDry9zOIgvDzKZ1mbhPZEIg/Cd4LGLXa9PKOqFd6VaaPS9umAxgm6WR6YTz+g47R
ICZ2XpzCYFYqvXxowI0w6d5AWwl5Zx/YSXn2ESzoC9UAIpey2T+RJxKCF68iPtOG
nnyWyn+XRzZK0UqDRxbl3Mt4JAUh2tJ+DD5liHuYsV65Evg5DCN65bYw9hwlWUjB
enKZsb/ZTndtS2QhYxJvHwfmadRKnOT9aznCnebj0ssxZH9D/JsTDuOr2CbtMv7C
WWZTM2c2F6NJ1B4rho3VSYvItOBopu+lcHTKlL32Rz8M6/3Mswspjo+uYjSCPeAJ
uzE4AUqpnXHnOwNZCKgqks83UBOTzOvnipiodQM1VRO81Lx0GwwxQwBtJ+cdEdXU
1ex+Oh9I47kVl6YqABM5bb9YS9SjpPdiC/k90vss3OsIWlEDy3Hq7WKPhVmCuB3Z
19AWyKKmCseqNIvbWuJqo0eLBdtV6dih/k4fayN1hzhfdCQ5Y53cem2U23tjG2fc
ltCeoYuprt8hW9V+SACcOyRSee3J0mtNtlrq/mhFbBBlQmQG2YyMt0cC0qkJoelo
RTbfaiAIlNLgjBMRE3MwECqDwNmP9stWuVeC7CH+SkdGEEU8//82JGHmr7U8OmYk
CMFb5EaosoFt2bq7AE4dxvrd9A4LwQBK4cJ+YQjxWrMqRzJfUGtwnVVs2tg/drNm
YeoWe5PQbO3k5wPWHky2F8rp/G4ZLmqEKdsiljBoyGRmuKZxW2eWg6PBQJgL4XrG
mMZipwRS5hkfWHGcl+8/R36izbl1/RQyY5gklPB+EkObpEYq+hgI9OpvJuaJ3YdF
JkQUh9cXRyNwbm7YWE6t8Feqwd50vxOsBwvxulblCXIQ9faI9pZkS4AwQGaYTGwv
OkMKSvUJLgVH7N4yUXbZEQQVrFCJO0vv8BjJ5m1NJOfSx7KCqwuG1FZb/OWAG7q4
FN4hQDNqGR52uozDB1NibBAyTpm3RZttVfpiE25VEMx17mrcGncTebu4TP15A9fO
RO1uZ8frW4YlOlIZGFEa/eq2eCO9mxmoMWUfcRDU+6r/DfHgtXZnHUFp4D7GpKdC
DMgxiZdEs9A4N7xkV1lDMkGYbIebRvu2KPF7lvyTYYLHIu7ana2OOSQHU+fK10Hz
JuhnJHBv4dIO5ivd+uYWwuv9M2Szf3CaG2QiUXNUeu/ujOLsZn8D9O2ecoHAzERc
ZsRFRMEenZuP6VdkOgHdWPfQusterob/X+43RfDUZ9Zguw7KiVTF6tsTX1nI+XFg
xj0MQwsx0xWYGosEZfHjROAccyhRbq8Fnjg8PpvUyM8u+v4JZwijAtHBM9JKuwrc
fymNKRoDJakMLtCaAjB6yjCihC9GoZ6qpiPHUEoCjwmMl4uSBQh+3Tl029M9r5W+
iHo4Fxbwxw5aoaXzPdo6xn1SVPhyJ4IfFaHGX4xKqhmkyDm1Ie2b5t0sA3P5pT5k
cEvhDC4Tt09MUh/NCBMHJZ+y9pXgmGyXnoXRlyoyyOLA32OxTWy4kqA7ZMevnBvo
OmZmdiiBuePX6si/7Ak0zZ/EqtE9XStmqJlx7bWGhc6wcNqi9SiZEQWFHr8dWJf5
EsOOenCPl5A/5P2YFFPW/bACr3J2jjWPFsx0CiCFD6YSY/R+ewtk1gryWYG28EYd
XEFRSB8BKTD2n/ov266h1QODYkZQVi5Nv46eVUpgG+WzoTeIbyrRnRUP4I09u9lX
jET+ilZ4e8BWONJsrj911w1rlhhwl2f39ohbPYxzniTTjyx3lh2vsTxbGSgRzdvO
2H18QFCa6Xwzl94ZLKDnETxYl2F/l9uXOprAKjTwaGSc8Kceb25hiCIyWKMTCMY9
DoKbjxiZvV9Yyj5b/2M2mcAfI8Gd52TP++fugz8mJ9h3JML1ncinX0FzsK1THE0p
Iusv2ITxqMI4yeYQ9JzVa/SmmRU96Ah+7GYWCjxPCRtPTERPde/WtoZYHEb6ctPD
fi/xlPkoGB+5p5eGELlyc4Es4p8eR+RbUuVBOQn6TP3od6/f4d4lrcYQEXtxEFJZ
sEML3dSrEsj4e+CsOfg8vrL4wRgSWY/NP/JeL5fBMtaIgC34VQE5atnRWLLW0xS/
wtzncyEDt+KCZzu/5Qh1CCibRLrfjtpRrql3fJ+5UA7t1cvAkkSFOOPTjVXQwlR3
shNZFpKuh8RzfXpHBuMGEzerMfJRqV2i41f2dSjpXDd4T6yXv0UTpwP7PGXZiM2G
Ab7G6fQUW8GU0zimPrUp7miB2LZTvxSyoWZO6pUuzgIsvGkmoALUUL8U7vCwQw02
UJ608cgE/Or1vigsM3rSM232I8nfqCBjraNyUkCxpjsVm+IOu8zNbwuucp+TCUS9
EJoLpXBh7hkgD2PF+Ot+OabAASzit+miss1B2dW9cfjgTuvN41x4nZCdAdJKJxHL
1tsm8SVM+cI3kjy6T2H0/Ug/Ri/1aiAp1Z1YqMkJ8WSBXUjtf3UBwIiaCo81eosF
jIEFpoGbCxoBTCdplRUTdKJZuzCrafgYuRyLUyCKF51n4OudvQUDHNXZOmLrNZ3p
hyW2de78aS2zbNWV+mH7u2k+CpUMXzNwx6rYF2j4p/Fkexu+KXybNd0XFyiN2m47
T+VPvQ5Y6uXkIs1W5M6YXYASj6AZvidOhPps3cfOQnEM6u7hzSH6iFItAbxxOktf
LBbPXAoU71f91Au5sw/g34YsY78Cn7CYP6Kt6ie9fHt7id1iB4Qx0EuamJhGV8Q1
Jy3GXa+KqQiaRyw7s5yq3tmlqhgXV7C/O5KSsE229ikILkkW+epb61/Z5x5CtRZ8
6ZuBRXVMF79ah4kvwsqQU8EjyDU4lafl1/ReJqmaFNbQzjvwaNf128Yy0XIQqm/h
iNVDyW63jf5HMB12CaiuczTgcRN79xKcDOcAmhfa3RUB6ZKNF6lFo+wtCpzMIDsi
N5fhXdQvvR+DNVWDIHWnKnrr22Tupne6B7rrhXiFx50c6gQn9rD3zCKVbCeUH55H
joJeqkWKYInfxxc3KopeBDnKVt2cu9m6s5nJKSV4YKalOsPXO6Fv1bJaGFvLNbOX
x/r4zjrl2xILmP5MM4seesSwxjDWSIuCc2IPPO3I/lnYvJR1BlFQ0/rnDaPpyZ4w
61Hgbt048TMVAIWB+19cgF8WO+mxOSggdmOg5y8sCbQf3HEhKGVsfaqZnwMebqwF
GgKOCMwLMPAtduBizup6byJefJmWq+fbAmvzu2PiUPKsKxs8FhzpqZZC1inCNHNc
mZJ4ODyCBhkOAtV+hzvttztmVjhMmFHcaiE/mHgLHUiGkNFC01bmdOjXbWWm8ZS4
ZmKeGMVFrVHLjZ3S4DgSJndSampP0YijrAUEr43mowkjUdi5zyl40GMR6PrtmSBl
JGNXMB8WoVdGff5dIbGUJMq8hf4OWAsZEn+P9b6P0vE2f82cK4aXKOydCZpdvzg4
apBr6hhvOBKEWMxop8wj1yvHP7C2cdiRy3HwYiQqwjPhUQv41FX2CeW8ijHZpGDb
6DfKMvxLXnvi+JyyzLfYcurao5MjNNyKqv1zkZoqdjBJopjBO0pniN6elFQZS4tP
2erjfCvGryY4Tj39z3fEMgu3T7ElcDB3PJ1ZZfr9HQQ4TBaPXwYit/q8D/o/6KoG
NVa5O/TQtLAefD/FizbkoQ==
`protect END_PROTECTED
