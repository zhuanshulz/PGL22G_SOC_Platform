`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iCNF300XhxdY/Ak4p6QGLtoU67MYPKiuMGTR3z+k/96/6Jk0I/3TdQ9ppHMHWomp
ZEY4Ljya0VsiS93/HAT+QGMoTqshbtKwhQek8lI1L+drx4JGqYBtqgg3u4/ryPLk
tOHm4GWIKPVjCmo9VbbbYWrlvmb2ykNDNURIBryxPMbyxYHn5pvar3pMNzOHuIuA
+9xbIzR+wd40VhGPVMFFt2NYyitjEcRAWe889spjrZYsnM78EI1D3lkricBQhBT8
ERBVeQayAF9cJpeQXIUJbA==
`protect END_PROTECTED
