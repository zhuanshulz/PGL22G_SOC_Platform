`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F/eSJo9iBSDi0D6bxGYgUCukPyfA6TkyrsM6peA3AMUSQRnlDBZbjHoYHHHRjbFZ
mU1+RDwIezTbsqgfbJGThefNSWj+4a6OVI/mlSt5GbEzrlBSdd5PySQUixVICaFa
qDvuqvj9pDKhY7rd5L+6JpeWOG8YW6+DBA5XkgcFViDEk2CHkPnfxp6JmRmaJYf/
Xq+WU7CzSuyKY84aHaj5Ra37wtyAZ35Kh0MIZFq6D+SWXYlAZRQF5nPDyG7TFZXL
ysiW+UNpu8MH21uMoxxNVoY1xdF999mJilmpiDIP6aFwAz0a2+pulpEcLAjbgy1f
2MW6K9r5+x5BA1i5IGoy4+E9RSBT4fPvZIA43kw13PExu2vi642cv45qix2xSx6Q
QsYUUn43tdpgZcySz6t8f7dfBo0WDKgagQMJK4HuIB7h0agMgNub8+yKxXz/rjDM
omt8mzlmJ9+Y5ZbLZYJmRvhgGWPrf6Mrt9OzHv9tu6aBMwNhetfa36v7aCFhLPy4
L9Ady3OCxhk0tDt1Jg44TWx7REiIpVbpwqX00D48mcSo2W9AdCCY6fmjxpOLYJG4
z6GkLxz2ZbYbZhVBsMoyx+cFn1C0QA7PAn+94J8OJ9Qo3oXsW7D34xpfA2euIifm
tPTB5X4MOPBW+ID2Q4Z2N1tmdSbukZGFgbfCALBb8wSJubz1RqHuqN2z9ykSJjaL
QUhS6HOSYAL66LQzl5D7hIdRX7TrXkYCQU5qzoy7bb9OEnVFyCVZUF/MqoJYqUvK
LHT2oAFuVy+W4G4qoIyOjI1OxgV273h2qpTmnp3Kj8cby2CM+EcXQf/42hua4TDO
1OkenypzP/8HjoVC3oDeGfYuZzvY8fuzE24/EDm9N+lAmnuO14ELWOA7zAyQ9zlc
StOvtzNO2dJr6Iy1Wk0gWGaFRaqcHtajJ1fwFrxVBYUHg6yQtQSnn1UYJpMtP2g0
rhDrQ5dw7Sh5mXvdDh25AezMjIihkFPLfK7GUl++Hprwxx4zGdLr3HksxNkwstel
Fn44O6JDztYTy6tW+XkKRK9xbzYAeJ0VUV1oKfSzU9Mis+D2W2tcvp/tQLUeOap+
k5h5rdJ/XnV3LfsJ/p0UfRaA4c/lJtySSCrIZOXokmKiRuG4js8ayKkrBDYqtKPi
3/VkNBAQMUQBr0KFtBLqYNmeiVAWasVjr2j7l2Ij2RteC9BKU2xW4AC12dLCIX1l
4+W6Uwi00im461rBFOC0vYkaK8l/dVE/1TErPyorYzytdBwQYIkQc6buzR3SmeGr
v7hQpfgHinldTYbeq6Zzf86GWm18LQoPcYPrBs0M3rtyg7Pgytx1o92biQFgl+EF
Lfb/cuBKivFPQRgLYvWxgO+7JuuQLkx7TjAMXyBauG4Nm89pLxXO+j5DWwe/Lr71
dS02yLUjW97nfSGl1nCkZFEolXe7qfeEMCbEPhw8vetlItULuacurx80x+KoYz6y
0l6aACN8VKvokGQDkHBWOolNkyFCbu+3WLw3eOoWx10PDbBTAZKvEMUobpAtaXeZ
zRk3zG58nHOaZtNYJ/3JmKBpmMdOT1RiXCvN7dTpRvzfm42XMyG1IYLkHXT2/et/
Q3/8ye+VfkZwrg8TVoeWKgnTT4bdW74K3e0V+rXGl0/TPqQokyFI/M/lXlTNfsKT
S8Ei6zAtBKk0WC3dZNAY4X+ZpdB0LPtbijOxKmn2QGI31uQuOu79KRvduHrJ22+a
RiLwHWZ+rZ8OB5sktEXhP5Isqpe3yUoe5aveV+BhsQ7NO2ZOgdrgj3JHZF2R8kMt
NLkz7iERnk2BR8HPWkDL6h6zaWhYsxtotUMvvLugqcWAJGA0dgdGUjkbKuUkhFZ9
Agqf8gNoRcYKer4BKUqNRl+LpCI830Vheon4TdbHG8PO/BmSXkoIQz5FFEO4Iyif
ztYC6eqE16+QNyvAiDHikMYiQ2Fqnq5kH4nXL9WyP5a8alOPU/g37wUkTBDURWJm
GLhEelWi0TTfUdCiwvaLiobJIuqFXkTfg1l7nrBw1Nml2KQ5yYb7hQeLs6C3K7Jy
TH7x+IoIfsnjl5cVVkFwAeURn/+X1GG+VLbQNQE013rZja+fOdUgZ000yeaoebep
NUuhX2KxfU3JiN9PguMoj5rh51IQwe7ObbfhPHZN3xq4ahL7p06DyNfIV9w3y63N
oUOySWS8L1PsaSq+17GdCLsRrsXASinehzLgyEmwUifwj6UXWKTFwzef8LmWOC1y
mxd3nR3LVFmBRC01W1jBWGW68FlOgcowAexd8YajOF30Bp2wmj6w+xGpQ/QvvZLp
pyxq1Id+zWcJPoC1xv5Kb6bG2qJx2kd2KN3V+KY5ZWukeSaRcnqBL4cJJoOCW/tl
M8aplZRK4U4E3Cmk7GJr4nLwykcO39+y9blTa4GU9BcR5OkzNLFJLwd/hsp1hM8b
spa2PA9doz9NNP4DzSIkc7/HzBI5aarnAHlvSKtAvkr4FdABbZCaSbcRJRK6AUH/
OqFMEH6sksez94f6J2Z0sgoX9qb2KdI50OE2aQx9dHbWkmsizXetmlFDl3ZMxlJw
6Au7pR4NWyUH5m6UtFiUxnEGuDOCt6oxOZJYXllslw5ZcD0gOoHcqdxx5aofgUl+
FhXE8ZRaN+QAIXIbuBXa2ET3c2bCNOrIzqKbpsLRsMiTp1gviE6leFRE/xKLTdnM
/4Yke7wfZalXMaiq7p4uxf73XKCY289mUjsQREz3KT3+sjc0UlZ8E2uCpSa76pez
nNOBZGyDraX4/gl+4+6a4qloykpAdbEE9ay/e0ySFOlsAnXAjfysKFOYkt3VK+6Y
ZskaQZ6OmjwlN1hQ3fNnijw7MgCLQdVtisAUxVUWHCRDNV/NvO/5nB82F1U5Qf60
dq+OySpIF+CMOAg+ws6gAPKPHAzgkuXmlnLqTbS0bn2y5xFtrPOcJbicAaNZWG7s
8KKz3wTVeO7AxRfwZLrsSrEKEo7AduSWulMcEBGjw3Y4OH5bfeAKfer/v6DSNyMt
VNk0oeaZFGLcoU1xWec3uIWF2R5/YUkRiI9g1Ej0tV0waSBqbBRTtrtA9VJSOyIo
YSFkyODjCvmKGonryYFzoUmLHnsAcLJbKAVyKQO5JMZjoYF0T2NxTmOw1duVmhK/
paxF8j47pjgvbFv23pOzGYvjSzNY18lu+TCWeKJtnnWiS8VfEe2rGA3C1/z6foUM
TjRYigYYenM97mvsE8Yt1CNOD2AHeJRvR9dqjP/vw3azLguBKtN7uEb2McG0HXM9
2GvL6kiN6+CqEyblBMZadLieeOwnMbdxMC6k4QCnPmUeS+EY1GL+QVE1P1BlkUic
U36+h7hL2AnmZA8SjTortpQGhLohjl9nuyauilOLH6CSe8hCfHS1w73MhYa4yhsU
JzKYMz/LHs0SHDi2NKvATuFkUIn+jBRA59B9tW/tabP80Nza5yGLxW1ElruAb2BH
7mPZ3zDhj0ycFsVVd6ej9f5iRJeh1e6FyxmfKRs9/bCccrlzWL8wgbbJMOAPrVHE
zatibR7HdtnZBJJGigGXqCGYsx8XSXt19rI/FTrpsrJSJV1L9gxcSshMqmgPYzPk
Slfkrjz+7xd72Ejtr4BC2P2MtJdXrCq6qkXkub8QfKBkFUwzAtex6k1poZw3dtGT
29NG+XBlJDEKSB4LggjjEdoAzLHP47nW4Ix2Zgf7Y2u4mRGtLk5+6LJm/DmFt7z2
4VSHnAvpEBZxJVDOtqMB5RDPEakGRYto6Dxk6s/5jDxNP50MWf/pEIVhIZ8FhGHb
qKlzeMQOUzHb+d1ae60tK/L0Z6kN/BEVKKTt4fEeryzw3RBUNfjrgtZyD4jOpCyP
o1PrHpuQrTPtW7x9fACFpTW8pMpbWdi5Fn9wFxQaizf3QbrQEizXLZh9l8Ck1+Th
fa6Lp5HklfyIOdHMgtslbdcnWso5DIZvfFLTG77ROLK38/aJLjH95PcPrTw8n2sH
Ku6ItZ+T8BP6JxV+vN5ifKXVTMxUusNDb6FQj5rKvc1ZMt1XiIm9I1Vp6ze0c7bc
lA+DNDWa4UNJj+O2TR9SQAtflfuS//9T1xPxN7knxDzqkFT3uMi1jpyVMRohTBLm
TQ0sdnErjNbX3Y1A8oub/PC2w2tQiBi/02jaYCUTvqxGgrm27EutIr31Hpn6qKI0
8epj5XUmhfSTjxS6SrOQBYIVd6aiMiOsxqm7G/IXVgPfsykdgVe+zboGWkkbR/A/
wDwYo3Bh3ezSPmT785Pa9oliyz51vaEG47TB+GK06DBQyG3+ANZWsRXzJSJEYjPx
/w4QmmOGvTmX31Kmg161Pq5Fi+9YGDSDfD5N2mcczIqhNAYxveNmaB5AB6Z8Q4nf
59JYYsGRBzAvkJi4XLVKDQCQl5wdEg6bVA3nA+P4cLpgzpAGPWcNAIh0eAjRV/u9
ZrdKDe8sAOin5fAw/3zo5aOnxV9TROc5i2X0sdlNHkWPsBvaVbJoVsTM5/HwpXyC
iWsQ7aMcm/Y/sEpJe3TysBgOwZicVdvw6nExr8AcOlmBa25jp2zXBK9fZlOaFNNO
dASW4N2d55VoRKyPGhKNeuiVZlfii9Tdxm4XL5xFywUDrRwMb/GJd3AYxd9hf9i0
11+NrDDMd8bvIDcwtz4E2Bcaa2vrTjZqjQgxmyRuraQCOfD6+JKfNRsN42RWHi/u
Ivan+DC7L5Bo4Imc5OHnOiZ5iNL8oUTmJD+6smnuIl6RJab/dzeGntCLBA9/XppD
x9SFbNZegW0MvEyehonuQGRMddDzmOVF72Rmm8fTctCZsD+WDfeSyWoXhXzxGhDo
diX6oPQX5ZHiQ4mrCh08Nn50RCzuT4zkoRovS6Yn0NeLGHHakgdDjG//AuQTs4M4
iqoIzmW8mMHkblwwlRdyAhb9QYhAWQv5d1F3S9SZJrMGgcYG/lVbtUScOUYHdRv+
2dFH0rcNP4YG5j6ONxBnLM01YoWNVZ1hnKaAG+AzjYSznKIrotD11sZcv10SYM3G
KP8YZ9Eu9jUe3kVLauHQEVQZUcvlMU3BcISH03S2CMaJZpIE3jRJLCxlHDaozKpE
l9IYFkvNzYXighx4nLrRCS1KDyh4IEmVEykxW5ZW7wJE2mYjgkyZtbd7vGX9XL7m
LwZEjd75T32wgLgMcKJpp5JOVqCUs730UqLvBwxVTet0/dpw48R5T7mdxGP27l2d
TyXOOFUdOlB1z7dT3QcM0nLoBY4RTuDgsjeK4M3k18F6OOeCrmKMyO3txjeHWdy1
qWY4KFPoioovsrcOTO0N+hZCfU3d2JBPZpfTdEg6tJqDDX7j0WlSVW9OfuVu6ZJv
zzHPA0ajdSo1c1mZcgFBzJutKPcIV3ivQaTwQVn7gI9g0gD1oczd5rSy7qtCkXMY
S8Ju0KwzlZbaxamej/2mMnXZshBfIAJ/T99ZfGuF86lzyPvOXndvr+Xehyq0bQUb
8hNGTK1maqqFDRJpCznpqhj+ugwuG8WMbofbq+eZS444ZSvXg4NaXzoBuKsZbsho
ZkdU/8M3cJwJWkYB+iyJNNn/RgVVCuuz6fNQ6Jmkk+F1GbXqoLycgsyzO4y+AAOT
eACmTkK0NcyCXI9mTlxnkJcoiJnc7YVdEnsc3ysToa7tXwehKhp68kgVsw7eSTkC
vc1ES3GPBOcqsLWpfRSY9YO7SkGclL9Kpce8763WYxtCPHmCUhBnD73d1MBulGm4
WC6HPOVBmXeXYkyp7CQTnHSTVESARA+w+5YblIw0O3TElfsPvlXxyMGkj55ylSeB
k4juXZrJNAGMx4jRs3Cs/8GCMAr4s6gKpH9VAXGkyr/+sfaL0gej8RiQZT0ePwOg
oz0rTaQm4fZV9h1d9mnXaQ22YAoSEhu/kyGsi4kWbJJKpFEXHGcRheaGxpcXwiMQ
CTOhuBu1qoJYBuG1XnIalJ0bzcQBWA/EQOJo/6Mn/kqQFIp1u3W6l6EQGp0ANNdg
g8dUC9IRHvEp/do4bWSp/73QSBbbil6mV0w51E5ml7IIXBjkCrSdiGh2d7i5WZqf
stMGwIOgyeg0sVWt7l5XDj6CSK2GCJ8KM28TUiyU6zWKnJU36WaxME945tBCP0aP
42v2s/Hta6yA1NilNPOCKAfYp5ye+WWjVPaSkGf59rYPxplU01+vgwzs7Ne7vwys
v3WA4w1Q27CIa7ObwI1GmiJYdZif4BNOLeg80G2moKZ0Xbz4iE4dzwApZofdZzKX
GmIgDE0hTWUBrsL9vBLZseJoLjO5IWP/EUvmbZBYhZs77gG+sb37ehGzlX4yLcoZ
7ypUSousA5mWcptYPCO5QniLM9SugCYHOkdfTR1t5Ncn+coNbSvOGF7t84KO4AGa
TYXpjEY0oLyFUZ6HkzhXSWzdGzk6njFlM7Rl1PAYGGVitJNf1pYE3qZVUrPytbjJ
V0lVkxNx1LIaAcyppuCAW3AX4ogSz2o5EmNr3ROCdMh+VCn3573GYqLV4Kgcsl4k
bUxXzujH63IGvAkd8loLPUbOGsGHyo8Bmwhl4U5gu5DZ9QHEMcboKm5BgvLnaK7P
0+x5i73IlcMDDGy9vtdwZlU0Cx0JU9nQf2rhVV+It2jAQX+yviM4S754JEGg46xv
MhA6lAsXSaNPhoWC3RTQ9QfH+ElRhzIKJ1FWefKnJxarJ9ylIYrc3VmTKaEYnrsk
sUiMg7DC4vuA0fYAUP/vfA/gohcMOOfJw78kQD01uEv7Hs3Ogo7CX8Ojfl5PQNEs
wdPNE0IGnFtNAKv+AHOD8FW65u5PWKxXS/meNS9j2CrfZfGp+crVA4O6bEQBT/fn
jGUyK+uHLjKHyk15B7i9Hfuo1zuTLt9/VzffFZwL++Y=
`protect END_PROTECTED
