`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S4JYu7cTa0bZ05QD/ws4uR5UJPWzyFgPuTObOyg3eF3ZskJ69HpOmyetUBPB16Fx
Zj1Udvyg933yxWn5Us1im920bRsjlaQU5F2xfRfht6ozYC6zaEK50ewECA5j2swL
Smo8Zcx6ZyFoZcXdxrrB7mQ2uWtc4t/s8ypSoHjO5ThyMKL/h4NrKCfd7ydnq2fW
Mjwn+S8n/4Wy/Sou0rCx1grto+ew5pflhfU86VOEyhn8BU1a9XQsOkaFG/EwCRDz
B+9zuyL2f/lD1z9NLGuxtWHFiKxmvl/XrwrfgtZ6AdFzt+eI2OCiCYWuoAz2ZzFN
Nicf+8QRfOFjvFdzykqGw4u4EOOEgpO6YAK47u4FMFjmaLmwnoEXPGoTYwmbjYa8
9c4a2MiEypv4u7KoO97lMs/k0dJ7wTg6I5r7MNIMCu/G+UOmT4dVY3/lsJ2LCAny
peeUkz3ceO0gOoKkGra5B+sZP06v8jyMtq+/RiMoDkfQALXkWP7Fn7mb6mXxc7DH
v0/Ad/TIXvEBmg8xW0I7kjTmkWGlZ9oyQNPRq625h8XRC3unfDd0Wo6jtVHreMBq
25VL1KJtnyokYoIqiLFHeX9njjICTriBMi1LtMQbC2kdqY6BDatCNVl1BkQVVwd1
PseQg+8B4SpBvjs5j7ZExR4D9H05yO42iUMjm9h/BSzgPwMsZOyZnNlbW1afU7m0
+htvl3I7ObZ8Xzauds5wDp2zjcVMkamIp4fuqltXl43dqIUwR8AEHqS2osdNWQhm
0kRLoUo8kk4LwT0JMdZ+TkV71ScyCuxk1kY6lFwbElSdkcrznydEYzBf0tXsIJY0
dKEFQFJKQ6SGztG9g0alhX+io/Qxwx469a7t1R2c5+8iNuagN8RfUdT9zO3GIqXX
bap9NSZpkVECGvXSL3cpV3uNctepGyj79EjdbS5OWbo7J6maIbS4gdk7fZg2JX4s
DmBM1IxUfpqtKvRhcs07VbIFFUK1vG12a6nSWC2EBAIJY3B/pyrgqetFKOoDBQTw
IBZ/2BZrVNm6uTDA89GSii1+ueMgLcZBouSzeHrvXVYp90FywviQ3SEVyznEmtBi
a2jCdQ6RakYGa/+UPIl1SNYD7vdWG3u0zwNBH0h0odPMHCNsbS/zUwKeGB/dC4zK
Zhu9zoLY54QH+w4wfdvGv+cyj9DMw1H95aV2NLhXz4up+86L2Wj4GNvXGyxRVR7c
twtmOCvnQk4kumfs2I3eRK/y7uqJaY01c17/ewurVdc=
`protect END_PROTECTED
