`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aTgUY7E+KFtmz53XP0uTVGoq9K5cf/Y+rDg4Hv/tAmi+42lcJqpq4cWl3kARJy4R
8inAnCF7DOPv4b+fcpw3vCCLmR+gHoNRQQ92GyRtTxgG4rhn9now0xUQXmTGMTJv
boUYGrbonec2RouGQou/VLIbfkFcs6sECAuBEc3t3uWw+N0G7xbiwmkAqRBaHtUk
9V01w4ttXqlJrJLgosqevW2vTZNfe9U4/BbQ913jwS4haXSVgjhEDZZUvwHUv7jT
xDDfEPGLnWSjqGU1/B1bUYyIjmjTvHCfC50pCOGoHbhQbxu+DEJ3xp7JT9NrZlOl
HoEPRfnh2pJXoyUbKKJG0lZ3HUfubRplxBGhCNgcIA/NqSYbjmpeIBfXD/paIxl8
Whtq0cefTUX3N4bjF4xddJVestD2kBDoinAP5Lwvq22Fe7wIaQb7rFLyD5TYjevF
DX71jwxoRsUgIyswVXgj9ezZFK/rcWFfq0knY8npQuaGMnRjV911S40Gjw3nrH/O
B6eokrN5NCtatOZR3NTv7HgZTMIwJI+qWgI6CbJwJjap65/3B7Sg6eAo/d4Rvl1N
pSRC5YlkiTuH9EbfMocnBUqxrbC2tN6h7OsAWMqLbYd1iNcMKkuNXIgmvGJjLQF6
OHtkbOtWjOxDCJAa7JvlFyJ/Ob8lQfFGGCHhI4Z0aYA=
`protect END_PROTECTED
