`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kubebmqMhfLBEh1BhcGpFlKh7y/kO0WMunVdnrpnrotrcC94GE5aZ79p7YY6N41y
QGhBR3yqKPymiKbcSPt8GR58UNm+HKcmp4ApBA3lvRP/XCePsmTAsJskhTmCDLXp
jRCvhM8qTbdKZ1VZpSO5kE8l7pUuUo61Xf/iE19zEhTwozr1xCkPKMyo65UTWtFX
H8g9nEOP/s3RZ60rG10r8D7xqcgLeyvaVm/QJg5IDeWhfSIdmc5bhyAimoL3ZJE6
uYRF+1NhzKP4X3HyxOCGjAEApfnQ1n5nNxitU3IWEU+jvsuhhF6Heo3F2h0qCkdx
LeWUo0/VCKwfsoiTJrXJ/+9ZZJ4cWPRicBNFvnfcvg/hA1XoxxKdCwir1FJ5fMwy
/44KxenNxD6pTmdI8RFPBs5c4abaMp8gd8b4eKxM2ybztOPbqL1HKAwgKBMZp3tl
cleO58fL4QGlLm3vMyII+iBNVayHOgzNrV1naAW/bmZafxpEC+qeWjcxEmB5xrq7
DTdwn6UvsykRz2fclaac++OHIVnPkwlemazrVjJXJQ48T0m7DOrynSNGIYWUE8wI
ffmhxrQXbAfeBj/F42sqOKDq3cbzK5H8rsFLwM7ReI3lZrLfDtdD2IWKVgXSioXV
5Gxhn/tOspWCzABVx6og7dVvn2SrwPd5s015RROPpxmjoDzlCyiVhQX6pI5Wh8n3
HwxFJ5HiRApPDbjlI3FEy5iaOjSoS74YDmW8ID8MLA8ulFzZ3qBTYuc/TNDfNzqP
`protect END_PROTECTED
