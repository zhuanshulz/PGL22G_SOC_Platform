`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OrREdqSe9ff6ZTGoVCm2Pf519+0M+GvlhO3sDRCSXo2+ZvB3ZcP+6KSdFJBi2AU5
p+g78GNkYtkitwszMp03gQO726b8zssQg9PGE6VAc2/RI0w3TNsB98OLgPWJhRD1
WH/PXkKwCBCMFSXdNIx7LArI2xQFqSsURx9a3P1O/GNOSlKDBTCuj+18IDL3ta4v
czZ174oWqTQf5bg3rzNoJiU4ndVmIIUDSCzOBOpABXsGdiqa59vEN58/GXhRvAUt
TSEaKWNyF1YnkDsMX5mqvSY3aVSW5KI+YIaYYy1+js5cxpBJzmOjwdmYeXFvWXuV
EFDBuhQVeRLWbt14KqMAcrXDxnQ4cZojZwnefAZIHdYeApuYxx/Wuq5c+Alu34vC
AweUIc8PE40IBqQqmyboQA==
`protect END_PROTECTED
