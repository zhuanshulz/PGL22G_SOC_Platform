`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yEo4nUi5uDhyedHdFsEqrMuK0/mtHxlNT+VZVtvQKnY7VuUPtroLWEQjY0cowRQh
mU6RFW6sYddU4lK4RkoA5V5fCzfRfq8jM6yrxoGaGigXqTTDpiRbTmEXgfGgyu5R
rxiyArfa+nAS79KsopFea7TvuRbnEYvrnGy/Zh7pUUorcEBMw+WhTTJidJqhaBkv
hLqEAVEBHdfDQl5B/+NSp6l2+A1NKW0j2rpwB+Xo2YNv2nqwF04CbiDIepgcA4b8
qmP4LarevZi7i6nfFCJp8EQkqLkU4CuCE5cLekGI46aQBRTldNFuOy16bGwCEuCb
YeOfBRyMhb+DM5GC/M0CbZEquwjaIZgmSfwM9PSj9h5SgJqBYvCKjoVYqWsHRhgg
QWE61nMz/PRM9s8iZms+elDvz07QHs1UgrzfnkDIv91CgzE1Pi7ddpmkOhpQKUEa
WXxjsz0lwETcD5aZ+H3x15f6o5eLr9GOXHUhaQHIVPdACT9tj1h5ttGSN23u7niv
DxWP76SvkMZsgInU/YjAjXJ587GMv9ZL5KFiVj3siQdkfVV1mx9rNi3HnRrqUYOD
XNn3Sid/dZnnzL1cz2VLjX/iHe1GRFxzPxwFZjLoAc27WCZi+ArdpdBcA0f2AxOH
/LmQ+a/aSM1JXwza2cQkuqMRzE5ug0jmOR0h0v5WIAjq/HySh3r1wGldByMON3IN
dHpiPE7+y9/2S0uwqrhkOw/Hbb05P6r8pUtyVqYq1lvyC3Gg1ICF1RMCS+1YVMvs
I6CTMz2oAWPld5srUmOqossb4iu6c+nB/2xUYI89W+douTTsPdwcfVQQYnvgLejO
bGcZndPELwz54GMq7dlP0E8/E28OnrOOwKd8JFzDj5OQl54EguvjI+x3atu6R63T
e9mzKkw+Kszx5ylyDjX8wEGdAXMOqbJxPbNuP/q7B7juEB5yfNSteVwD5O9UJyOc
s4Yam/ZuldR7HLf5fuHUXJPqyHNIWPYB/WtweWI7wy94iyPxCcf9Va6YDvqxwVeB
CbIUd9sH1Eip6oZSo3k+96CE4Oo2RhhzwQK6PUfd9Rzi/RrdFucgtmtx2yfg7RV0
B/bIMPU7X+7UIsnXj4l0sk1rUBaraS1kdpzbUNdhJ98rY1jGcYydHu2yCqf8bLAo
o8RLx9P7nVVjoUjSQse/5mU3Xcmf8M57YiehgaC+x7ekUQI3HLUJX4nJBWTGJrfe
h+ms3oXgZvEN+xapzqzqodZaSuftItrTERxYienP+MEBoWzIuwiY1DNZ6Wj8Rg0t
APGvPU6qJDWNSMkOq6WPmhvv4bZTp/R+gOF21+4gjIVEOBVUYXj/3PiPA66CU0mK
G51HegvYXzAwxWk0CeOXZqrpxRAtsU9fmfC+eUnTRuFrKo/C5GO+5HIZNmJozADV
YJWkyvikXJV02D1OE7b400xOIqv63mqN+C7D+wgRsQttuFWFyPenjMV+jWtAxZoo
Jm7YYOndhbH7wsfF9wcvyW2pOT5lHU2idHXN+aqiEd53llo1cszT66ZF1WsNzu+r
CC6mAqVjbodu1lnrlTrbuV4wE2VK31zKaTVZHfk7Qll/5gF7UJQMlKcZW6PBRy1w
8bECHmiITmVs3tJCElaD3w01TB66ree7MycUKaFSt3U/neEWW7IkyrfuiTKjWzPP
dgOh+NfObyYN6g+62xVPRgWjK1XF/QwNhHVTtCFvwltKApyJJYZ9kss/d0fcX1f+
XL8di/nsAVMbGyeeDTEHOhFbMKlEu4f56JAsIXB19XkPiROKfVXqWNlkF/mbC4kt
AqXnHxbQSzNsSjFqsc6D6A6qxPuqiBc/vBZ2PiGfHnz9RTrS94OrvZqBm5ebOxSz
kcOHyv12ruMQKcVi95auTqDa2vpj7DGarZiYmPxZ70HxRnBWhDNGaqP1176W2gOm
MYs2i01ZRJi2doRfUL73mmpGy1YNzdrF7WTc1S7JqDrUw0TvHXBjiqSl0/kL76wF
G+7XvcUF+SH3dpUrLsPiSEcA7iXDEmDLHtYiQnsrZNy4va7YUQa3XXq9DT9bWpX8
+MKkXpgfdlgymIwHx91tR+kFZ7HIUPc19UM3aboYSnOBHBRNmT65fZXD8gC0ib11
8mb9fEBTbMH4N4ys5lZDtZPDeY836Oyt2Sj+5fC3333VvScFGktnq65PYFkTIX1O
aWkEnxQshTfqbbLgaOlRyuFkBl473Qpn8LW+I2l6KP959JjM9f5ZmWfQ3u++iouF
4FmTGFvaFBg+qlLTSwWXt/AXX4VGdZGf0b6/UoeXURJ7XTuB5LmgfWi8raD+mzgi
awT0na0iuGKm3RlLXl/2bPu+oyX7PexQiRdvmgZJOFcT+ydkL17KLkR38wbcRNTI
WdbyjfkrVym1c2tmzxVmKYFkiAtO70IA9frn6BdRfPkFnkkhssmbo2qaNTT8ufmV
17oGynyvvicjlVgaYaxe2OIleZUTjFVJVMSgCcJiFpduS6lwuViyqYjVe6lpSrmJ
ELCvp1XaDXXGt8eQS2adP8+JHpolhH2gDKidEjV00RiN6Hfg1vfXyBxyWLQlVubj
naNRGgxwCv1TMC3D2iD07ywlJ/ooQf/YlXm6fhJsBso6nqXxPBcAikdqz4exuK8o
V/qtiJAV2ZM6MPCVepO4XBC20CPspnDi7pB0+JPkuEtc7d6DcMJMMoSHCdehg4up
kV493IZuETiEkSZXwEuCf65B8Az+XA65ScQE0JjIBZMv4wi6Agevtsf3o6YZ2Ump
EFxd9gUy/4kou0GF5k/gru9KaDCwcRrDHpvkC+FJXXjCIOqHJBR0mntjDsV1aCxD
VnIulfZpSJk4lJauxREyJF67NH9lRjIWETULGkcl5MPvNaHm190aTypoAX/eNFIv
d7OHHT9hOVWIfhLaeYudPPIutBAxNM1/frow+wkDG9j+fwtOGeHqIv/ndGt/CbaI
C/gApRFGkc0rgZ0Tdkme0Uuv+dGVxPTWlUi1mz+aQqDBaC1w7flAWydndBRSJYAa
meuCKIP7WAY56Fd4Yshn8DvnKobafjJWMjKU6fDKxopEVhsvE6bDSWb/FT//oSLI
uBbBaL1ZS0l4P7Og1e4c8g+fXgswtgliFJE2igNZt3WyuYK2wlORBoRN1qo6av+B
uKeC6AQFHi1Pm5xy7BWGLiXxQDLgXRcEeNSdS+ooWTWxCxkL9utQHNIOKxWT0VuG
goQmd/SJW4LpDOStA/QJF6KYCVo07ugSkRqAciEwxt6FvImkIZoFoox6W2LMdDY+
zQjVRhigQ5r+mEHrm7Td8AfZfTeAmOM7mWI31H89Krl098VpedrqoNLXgHudfLp9
YQCjrrbFsBPoQhBLyGmd4ezWwp1lEGrr9c/S1/qlrPLiDVN0A9aai60C3xCI6H8c
UIt6l0nUcquUhLQjdPz96gk4WkrHsJSPYCIMxf1FPEgpmfNNouWa7h1/JBOg7Ka8
6i/u7HRw05SRomOfhgXNAvgE9iJwlQHzkwevu4hn0gHyao3rxSwd/Otk0FckPrhy
XkL2K0rUaV6hdjb3bewE/155jDeeGzWmgnM+DGA+GLsMMj4siIeS4BOkl0uRdC+M
1cUzGwKnsjWJhSkFNpRdb7V8FjHGww9eLChYeTwyxWM5LZLmQnrOGNxYlp3z6+Jq
pMg7n2k/MeehGexYbGjgWRYlyu8ppTfmwBEtdZMNd1GA/zZMwmquIdaY6XBcpsX9
FIrwicw4KYIn+drGTB0KIrr6ujxdlH50KkMTr/35FZkPs+9Rx3XN9wKydIlBzozi
S2hzExctIoHD+r746KhF+8LQ0L6wsABPO1MSiI+q38ofj8xkLZ72T+ttQs9jmnjk
rA2Jb57MXCyl1AAMsagTmMbfquiiEjBWDjKWGV/PgEmpNC5c7LW1AxZjFPGcbJT5
yRA9bIDCZNUnM80Qw7mi7fYDUon+ipqcy9e7TEeWxtgOt5NiyoOLOzQ0cvGvoKpv
a9HKZBmGuJ0+N8iWvynW2SAVYKVMX4vvVWDrWfY7tSt0c1Bf8+tmtUF9hFMhwVoQ
ISsq/uawea4T/H8pohi89lYw5sfoOveF7sOQ5fMBg+xyNtxg9ak81k5NCNNQ5Woe
BoIvyUeTJ1JYoC7K855J2kyVjdqgWk+6C0ypo9gTNJI1TevpiumocOWEplh0uWzy
EXEA3oGJb2yl1k28o0uY8VSAmNNmnhbth2r3SoaWnshiRk4OTC6vlWGTKX8PMeZm
UNT0Ci8OHm93SyeX33ii4ez1HGGkO+fn6asJ+zzkbGKoYUduAVOc8TA7nh1kY5An
dnr7mHBPSwpOOLrSQ4rKm+RcCu1zxKKQOl3b5ZPUmcA6Sro11ypFHukM5tPEXz8m
qYnhv2UQLimnf4lrK+49wh/oTnDP2S1Vskie/tzI7QQcdzKLY/8naaf4QZmS8EAQ
34BTPGflx26jWbjhNudYPiU59XxUoYPYlnuw8hSnRnRIBVTlxHYftcu3oXSQP8jr
0xCjVDXEsT7XahQsRydbeXDKBdpv2yVuOkljtaXtgMr/toT7r8XQp58uanXIrPjU
QBOI1OeQlSXaqKQVPFGw8gjToEKtnSoTMfT5hH0TBRQaBbvTSf2Ch7INsmGNAKGF
lv5a90C9gVRA10Vbv1sCSacR6+twT4PPICa//mlgf969WWn4qEZ6R6vqJmWqGtVy
M0LzRjShp1Sl44L1EzS8IJf9//jvCJvNe8dT/aj6lH++bKJKL/HubzY4Hh6slv//
Jg9C0yRMkpTipS7yeGPxXoJsjL263oieRW7bQSNXThDaNGEbS89sHONkHqCkjQhR
SKXFEQyDD5gywfYBCxQ3yOd21c6rKND549O66kM48py5FGd4uQSvYuOh4VMBW2p3
6x165pgzyZBpX+tNGxYNGDWhkmBrygVPO8D9t37Fsn7+3TqP4esEPuYPU/snCxRO
Z/30HRFFNKiCiYxvEY8U5J4mdjOXDCMHCxIOaHlZ/xXbOvGOb85BTXDW9WP5OPdo
CILrjPw7M7uAc+KpznNeKtuXfKThimqCWIxL8BCpY9WAKUKUtQGUFi3OYTsvClCL
c06s/7eeZRx1jqZr1Xx5fO1cjKyoNbuWJmB55GW2BEgU413ASeUtB6tnwxcjSM+V
36RYTdLVu9Ek5TPgJ0eAobkm7AhdMqd+Xz52ZyiWXmHICn58jC8vlFCMfR634DiN
ASWOi+1yKKstT3mIXxOT2gG0iqqzo190hnCuD+DC7ERZrVZdnL9ReE1ymHKzZjXG
oolZH8WBSj/Mgml/9+eJc2ggc4AX3pcIqlzdHjyEWVZcgXM2O3dreCUuib5kvN9T
rVQZUYHUwsTzNGBlZfb1/HWju0LSJ0IUJv778ah4G16L1/bfVll1W4UsnD8asrY6
FTmEaxOdvzrahlIBboIwVBzeAkH+Det0EXS97EGIv/04MxGjkksjHOys+Y0t2uaQ
H5b6kO7HatSjzpr2wc6YAeXAJFntk1tQ87B+WgC8nnZRsUlcSuBu0LzMhdS6QQKX
OoIAerS7zHOlCqD84amQcRivsjH8m+JICOoVYQoXedFDaiyu1QFLZ8H2Drxcn9yJ
MgMg/NcULup7lfFnb0F4aQQYnIaNTPpx0PnFyoPq7Hvgw3FGsuUpBiP4SgSVq0qg
t/ApE4cl7BzYydbFM/2GTWp0x+I1IUp8m+kZGrdEJvKvJ73k1KLaBTUshsgt+1Ps
4MNJWwfj8+dmULB0/CsTn5SZqXh8fd/FZeFqSojsMP8qVVFJBDqyBGmg/0I2FHFl
xETQGcjYeHbh6NhyFuro3l55uZWvQRxZ3TdZ0G/c7oR0nA8JNyGR9DqVOfCGiIFD
ZShYW71UAKu2H9XGZqE8p85WfyakNZzIg0CH+K9U8XNS4XeB5oz/uAJAEAcXe/PQ
waKgfzK4dRv7XUYFpPL/bTJtwzdmByczsW7+EHpfr2ZOTlKDOLMfwad72oeBwBp7
SGjiJcWVBLd1luka0tH/Q2AwwJdUW/HfdBJ5lZCXc6lWXcqW4vNvAGNAk9q0+Zqs
PrgDh22kgL/mnILEfEqA1qH3qUVk74W0de7zOEZSEWC6SJOQ8/zDyM4EyCPc1POm
76B3srwSC/5UQ9WRHm0ibeqhkCfP/WLTfhLlui0dAUyzLcXF8n6DpcXVLhGdXzsv
d+C0fgDh6WDjIoZeDdhinxHHC+0YgbGjs9tTosEYc/WQUZbrVZRZKYWRcpRp5FoO
ave/NJ89GB/lZLoGYpa6JiYSmiVdHfDYffTQGeq+TV4eawVWw5LQzQeOL9I9yhn6
oMtwFulG+K+DrN/ltRJgUJUIAm5QLX0dY5BLw6pPLmUlI0SV1LzpIrEw3V+VwT7f
B30AHVUySYVn5YHMjG3jPbzaoRFxYeBO4JdSCN+j5f7V6MPg/8x/WpKMgfWQwBbu
aD1FbWWjin9TrWpY1nHf7YfrwJZGahvbL2dR/ClUF2Jsg3WL5LmCzQcbfY4uS6EL
yTcoHL4Yd7l8nps2n9yT4nBQy2sZBYE5ErMsGoxi6fw5lZEkltU1NEi8ztfWI1mG
hEowePCajdQfCpAW/DISqrlZ5XMLdGMCNN6wukeSowaQQRii/qtuopfbSesdqzRv
fqUfVpbXa4FNyE9tgzhp6rUWSaJIaIiY18Ws9CbiTKhKZbGxusB3V9tJPd79HiFU
jCdHOL71TFzwL+CnLOSXFU3WYUGKGAkYjYo9xjONDHGOYx4tmJDvLYixzcf21pJx
f1XyBnFlfVMRX0jHq97EpSkAChjMo1euFKMWaqm7iL0fb1FTqWOJU7NpWVCa1sZZ
OdAB5U2E8o5XrSJhQ6Ixfs9lcNVpjCsSpJBZjX1PLNTtKDkrwDKMK5mO8SxRyeqC
GvkBaQ1Qyi06bkNbisa7dcXlzNas5KzVPaGoWhuuXwi3ARmP0M+W6CPpUHms3EWm
6+EVqL8j+LNKcEOw6AJC8UDbNAOICV7+Li/E9CYqh2whD+u+puvgNB0BNGkH5gKQ
e14xQT/I8SAqoQm1AM2LzdqG2B+QBzl0DQ5rOfnCBDYZagUin9MroKbvsNB5uehu
/DE+CxdRf3KytgcV8LB0vI6oF4h00h4U2/ua36RDk0TW0ol7U64GJIZQoGAHpN5j
KxEsvfHFKM5ob4LUsvPcqFZMvjcJjzHHMJebtXPhyHgnyap4pRRWBsoyDOFaudPC
K7w/ezH3JhSCOCwDHX+DfDfmGALN2uaIlAT8q4J0O6+/5lPYDVpQXzalR2VUnk3H
pdDEv6ivyFRXgWhpx6IpLDnImtrWkxUy1Dcy273ZsWFGn7bjgj7+HmBI6DyHZpxe
P9ps6AjDG/nVmlHAmUHodVcS+iJLSF+XuNOAnOX+kL7e55jZOe+GFybJK1Kra7ss
vR/lAZUvaJBjdgugXXirZ0C6ezEMIR9vAkdIAccrOvWAZwrIj44EmNsX0X8sj8wT
TiLUZ0T+q4UFRRymuocTmjmjjf17NdcVxFN/uIVAUdBioqdHgwwYHnwhuZaKREsC
hwIl2Xxu/7dgBLwzja5e+KZXHscZza2gkcK67PsDWzcmETBFiJHccVlIFRrG7OqA
HKV0ZGt/oaxdqUJ/cqLCoUS5TEiyR2ByuZ82YbdUguf3qjP8OqCy9OS9De6LakYU
9MEo/6n0k3tdde5flUc8zs/dcm04dT/QKg5E7mknpQvqzQ/UYZ00ly0EPjOg+7Ty
5HXpNtt0F/hNvajXMHE5iI6mgQ508yPx16ARH+s0Sb19rQk2IYxIzHzwZ8Dmarae
pAscLfKhdyqlCytQQxg5V/wgPWz3dno9Teh8mqLTh9FtSOhowL4oTzI7eNAPFYJ5
ghL1Joaktkbt8A9mGvSDluc15N4MctDtMFh5UH1AyuAl8m+0ofVlgkLzepyBfPHk
zbceFyqw3kMNSZpKLx6ZmpFUkSoEqL2uS1zQ1TExPIKUBRPy6JT2UvFi+650XYRK
KJNS+5CMMEeHgTk+8hGudf/QeQrkrIG3A0XsCv66VacBDvkCBWwcylhcIbi2EV7e
7rby4EF+EQVVtmUp8OIA+MF6tGWjQlQrwWt4KPwovSS+sK6Hb3uzcWT/cvnkg98D
+m4chBGvXhURcD/TYFpZ24c8YgxUSglyTXke5WxkytikkVrfXsGECaX8r1JIdbM7
eDE64vF2mab4Btr17GsBix0t3It3pLsMbi8DDuyntHOcwEJTcD1zpRav2/VRKt+E
EV85H1JUfmCBsoX+y+nAQd4IQGqX//Vg3b/pFvA4rfda4x9v5XJC2SkUztSag/w3
+3rMKr3yyrYWOcM8X7n1SzzI/p4MmangF6ESFHICFZIBmBWiXjCU6rFqXk5ChGvu
XhdiOTwJHPTpfpX5TPu8Sn9tEpKLPScoTWjOV4FFM/iic7KRkyJnIyhJz6OSfk0F
rDxMI/ZCkIha9IBI0y2uf7gKdytP6d16XWpFrEkXhl45oT1zMk8fK+eL0W41kHIM
R+hui0DdWNIakuRefxJECdg9agDFMdFGipXoSXUAWpN3UW0AXuzMkNkxRb2Q/qFk
xIe/G/OfXgO1DPV4LY/d6gckVQA68mw0OzyzGQxicIzqsgc/pBiyHwel1oTBCMiO
jy5KWMXsSWaH0Yli0knKhCnM0gubTo9g3wnXQl/abTLfJpc5DKa3+MHkLHwm309a
9+Rg01C8mCBj/yEeK45UCyaY47sbJC8wredvTaj4gwiOGPxz75Rmqvgv8drKhuOM
zVd21bLDctTGNJi6Y7FSxhPiKNQuuJno/N6zxSbuACwP/WX4No9Vb/440Qfw6Rm7
310JLekPZ4OZbuELq6VI3KNHX1AAElNnsBjSxhRocZE2WjUlTK5nTMWO3aag+syw
+xJ2xULB5k/zC+qeZQ2lumcIIudYZbEo81Q0ro/JUyyl6ZwD4WGqFTud5Otd5Irs
eS70oOBoC3wng0K8Dm+5PR4+HG4vmZd0Fn5o/EdjAwSb6a7FjOnHhivwNwfNzpi1
VzHwFCAdehqI+HdH4ZMn0piI4Cde2y+iD+MRbsYiZAOyQslz4cUdmBQCyxdKzRSN
nFFoeVtGnTPIGzVo5qVGlUWEQlVskzUlh4sLK9HPoIxkWKHPuB7XcxRwFlMwfHh4
z9bT9Qf0O5AqIaaFouf/w8jD11lRqkPsvGxY9OptKChkFe338od5EiwzBd/BD0sE
+jRMexSNFgs0jU/uzZeaJv5PfycP8P4/HgwA5H/nfoeP4eGocUrSaaGDd3LcuyFW
3u0Ri8z8QuG22UhM4NfcrU507xDQqko4ESCxMWkWA9a0dkbXu9vHRhdcLLqWztfd
4VDkb+v44eCMpCZHJsMd3PPfo228HsUP8TufpOZN//5AyA5/fsBbya7DogSu9hAT
1JttV1sIXfZNjfXWs/MITkecHX//PbQe9oYHu8w/3O8cD0lDBO9AHgkckASJw5Po
5BqhK5B7AgRK+A5kkdr14uT8bv0ZEK66XWfYgOzmcxDNwKdYKjB+6Otd+mKk1E3v
lbDNT8ZPvZMIwZCdrYHbnhfHKvshF9RlgMWEC7ZJnSkDHs/xL2pwqzf8BkHZdR77
Ri3uueVJVDVljdUzzzlM/7lSRQkmVSBbrxORkL7bClHSpp92C0rpbLIHBtszMp69
4GbSZSbi/yQ7Yr6quGlZNXE0QGHFc07zzDt5qYcr7hPtTzvVl2VTizgcBTvVrZo0
INlM5zHm67RuyUBMkxzV5xHjyX6WmdGHzhTMHlyZwHMz+4jcdSbHQ2IseOKuoor0
jFFlBMMIkyo7ACQANFod0Ed0RSRNc3gKTCN99vxvjtXMxoCSxPFJt0/+9pV4lXM6
9a/8bX3LS2nKlsZiLVRqCGifPIF/syY3t+67vNRPOLxyqfYI4M/SFLL0q90EJnyc
jdXJciW0PClhNweJNn/W65W25wIYa+uHvuZ/QbEfPl5uQwfVJSgGmkVR07D24FmP
2RXa5n+p23Sz9SpNh2wYH6NrW2CduoNKL1Ns7UtMVgHF7I+Lv02f9zKRaUnIpEaE
YxpQ9zwKHf9VVA0fBfrVsdX3pqS3rvtYC7hBucb5xgao95rS4u2uJwk1MRl59FWd
o6ZYT++MPx/1D+8egvdT7wDyXL39Zo/I5hXwyODkv8GGE6rIczVoh9u1lnnWXGqe
AdvkU2Ne8x4QUoB2y/1O1F9Iqba+DU9KQRkND50dq3piV7jMcegn8Tj7gH0EU3yL
K4gKoC2mis1UyCMUdxkzvacAkunLMhr2xZordHqfalwbMG1uLj0sr9grhji92utR
JB0O3UlR+kWxhoKIOFtP2TNSo6c+SVewFyTRqrmA+hvedS6NLRlMo/9U6/g8D2zc
dEGD3kU1CdKpAysnrhTFM5HYo3hoRZM6FAH+pQJ5ZdriISvvGfX+gWYvzdckLcpg
47aBgpODn8v9OUHexGUOhOYFOScrd03wbFm3dAxGjZP/hOEyY5qdvpUd3l5qmxgz
Znp6JDRoiYSp+Sw21SeNjSpTvnS5g6our1gnjH6AX0RAQkmfhVPNyHzvRYBNocBa
1hAxzTJrLzaRnwWQ+1kyXRNgPie53DgFPOemZ/vqtbKWbcJMdHP4gEmYjOLZ+haI
XmsSM0EjRcAEt+9YaJqKgwisyVHh3In1Bxk1DxdwF4d+QCyQac+9V8pr2YKjLQsM
kNBNyvDeC8TmogAEolfvtpWpHEGAAENy1o9np/PdQH4eV6/IHVTbdTuPmPS34fGG
avyeZjdS9lIySMR/9fvHgwt7tBf+yqhaXYOhfnM++at4XN1CrgBfL4DCbOdkKPZZ
oslFnR3EOA8ong8fFgag2iImxL103DI7ZSPGT3Bx3VREoUgzYEhwvVHa+xe3qfQa
CLsfAH/LtybplkmePNSqliew5M8VcXW/nTLFsLrFvdssZLmzRp4HJR4S+orrtvxr
15SaQmqpJz1+sfu1V1+XJCozx/rQm2JXI8dS0z6CY2PhLnTMIfpCVsLn6o1jMwAw
62/AiRl8xzGBs3cvFPuzlUEM9eEYIvzMQ6KJYm1QmCXVZr5JL18+t12BYeb4T2VQ
z7jHbQBZjriYzpko7nGNzwXJuQ7/5oU7KYCWrce3qFmrOTy6g2PdKUyR557ZD2xS
E7fnAkDJnlBlCpvypEKeqZsQEbcbmZLMdhzEuTP4eKYMzT2DlVCeiwGOlRpGHpDz
z19tsff7bM9gZEK0AknrlQTOJO/JbFNv2qkDPfVCgDCResEFi+LfsdQfE2qoDkCR
3PDnYNAO/6l9xUn8OCFXWJMUrVcegkBYqe0j+/8eWfsFXoWDpyKJcSjPFTI0BOAS
sImbD6quYW0UAHUwHsmntWbkbkNJLqJecqZvO/lzx2ZrgrF+dxhkAR/Ik3LKHBTc
IPjaxG8RBSgZ84HGcTKziD6L9ksOyAYshR6NbpVB7jgGzOLTjNFiFBRzW9Vjt81N
NeKwio9oikdrLAyZwhaRkx0FSZ9NLDvyeIhOwIfRKEQ9bC3WhoxXM21EeI01E36v
DKc4Fl8pi6E+Vpc24EU9ARBl0wZhGOD1cVTK5MnTqHm3szwIuLvtS/rIpL4A7LC3
8imaase9KXE4IKgVtTFpkZBiWKV1u/PihUgBlY7eoAYjBIxQNzcCd07f27JEetN1
xi7NvWa0TGwJiOibm2BKe8yASY6ueU5xn9fyuk121lQkxbaFBSRbDg7gWV39r3o7
fwoj8Kr0BESmwZXLsRo8X7ZUCzsKEDvHqIVe+H7tlC6nnBwNwjLdpURen5gQuOsd
fUUvKGxwV8LU5q8OqO3SsXSVhPGP3+BUdzzDhbi/Hxa0mx/We15l74Jt4irzvQjB
e00avdVp8Sadzd509t30Sd4XeWXEvnkLFTbEUeHJQIuZrVJRMuUhjFjEvpUshp7h
E+T+a5hXvNkfulMUXanuiyajUYMWqJeszbwxiZI+jwOc8RRExdZaz+otKgCWr0Z9
jmeLJKgBHo+chEh+23ixu+KF8NuJX2QWI3n/2caJoox4ZxfzttBxzv0AuHI/CZf1
Is8CdL5qPkIgXOzESQiKLYn2D5R2kLLoxk10/1cu5d8/4Lgdpqc8VL+haGSvtsPO
0JpZOLV8ym5Z0GbiV7RLxVgip+tisaYCbV8PskjL1Yu1sVibtf1E9CvC0xLyXEET
5u3QRod2Qg6T+7NxUKjCnqONw3lGdJZzUSPOxqTmLVPKlzVlcJIkxrKZ7KEH8K5V
vCx5SMeYoxCAGqgxXARv0JsbUPgE7EUDDMvn9g9ABXn1SAskDnT3Xmwh2v3F0+P0
+ZkJ51BP9d1PKaa0aSOC+57aBB/ibOQKw6GzYzTo+mr3iQoCic1zqKcZy956kz+4
s3lDyeu4Qmb7JrnFNzOCAd+DF60kmFX2cB97LDHMLCDw5dkmnrAvm7Ypokz/WT7M
dHASb6h2NB+3ELiVa35IyB55TVIbwOrvLpA7/fu+7nddDgfa3GOipK6Bzn0IoJjW
nUZ27YjMW9fKCc8J2Nrk/AYmouPkidW3hORG9mFJkSA4cKRK8hbGO8nGi0vnR/DP
GCqI3zRq5QdTTgUIKYidV1VmkV4DcuaPT0adOsmrHpxvLELL9HEhj91SMhDBcAxy
3XULvbHoI3H2dqiksyNZbB+zJzQPts4KbkHPT5U6jSYwmR2E5IQ7dV6ZueLF9Idg
095Bvo8dPtpnjv+F9QUwTYWG8Cm/iksbC2MGOWonDoc3fxCzAG63o708wKreIu9+
iNXe38PYs4iWbm0SVWFmI1Lm7f6NlY5lWmoD1jNG8IAW4R3O+loWHgJykRMBIM92
ZMovg5kTF53JypPj/qnaxfgRPgCWcXWcYF+G86oTIkBZSn1V9dsSbiTNvSGwg5DH
Z+PVm8TmS2Rdy/N4/Y1Y/ZGPiQLBhgtkjgs3nwZOgeuVBwT45EpuGfMbZHNEkGXO
OIZTtu7mlWR27pLVpFGfGVwECV5spvVOr0EKPiO6xGANCfz1fFg7WkGhKjL/lgig
3djA7IdFP7K38rtBhltDoK7R/sVc/nQrKDryda09YWFJGb0jT4TXQoXNlbFDhJCM
1bg2O/U4ufY+PcldDIOGItL5GQBex7ZQ4Zl5u9SymBu3Li3yt8hnMTavNmK9XIez
7Uc++0nI7QAaFR/FK3DY7ab6fITrvVF2nwc15vQVaTtxHNx/A9JBJ56U4swBpVgd
xyAyx1JKHDV9j9LH8xmvWW5kjNjBTe0DuhSMS/ElOb1211JpKiL8QdqOtrHdRYln
zsh3Z7TdIbl/wV+t9yczMYIpdfkdZjefKmXn+bjrViyXMW9hw6DVjUQlw2ZI0mGj
4s13HF+JtptY1RgPyqqqVXR9JMvfB2yIF2KkE5D9Fb9EX/y7zF3uONK0g3BGcZ67
YfsA0pM9zDH13DZXFFEUoEVOvV5ptPn3I4MrWSFRqanlD7EUekmgSG2Y0dqgzzJ8
zuvoA5/ZcivFR9dB7H1dB+DK1Vo1AboeeA2mUnVRtydlROUHire2Q6ZuTv37AqAB
oytaMCBcTOvEeMHG1ZgY2tgihjlx4KXmEAJ0dkGuRxWqfAy29kOqB71wtVv1p22h
wyh+wX1vlVXk3rlYKfyblIm529z7excGlXAIIO83YKLmQ64sskdLq5cioOUJORUH
R7xhx8ZreYYxfeZna2FCkuQIBNOpBjjd6mlNsoc4G1Rs3D0wRGP195K2Lz/6fycO
aIMlK9j8zjYxGVhGGg5aM4a1YePgcX84LD3PZQMFbUo1mw8iYlm9PYdb2gvrw6QT
CnJ2l6ocwy0/9E8xnl38Yoxb0LKOdKA6akAvG8Lo+hkauPb+AhmBoz3f5TMANaMk
Wkl86f3jY3GYJQ6OLGIggKqtqHpa8UYnqP0NbwQLtKzqAq9fvJDd6hGVZ/0aYj2p
77vwT5gFuz55aGNXelfwnIrY8FYDM0qYZvb+ShyGU9VZRRL7Zzny+SIvF32yVa2N
AevbdBYFFAbkkQtkyieRqy/DnBSpiqIh8nCLF1sseTIGVO2EFqflpkbF61wUNGHu
938TxMlnYnhmJzzt0l16gWmeIB/TEqHC4+JbpG91LCQxBNINWD+OeIP13wuxWi9H
zG4UKGa+dysyPEpW/aLQsSSDb+VUL4Zf5NhHb8w4H1k=
`protect END_PROTECTED
