`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aFDUFRGj3RMMBC1VJlgDyO5hGyzyClP9XOhuTF0czJOFGNb+rBbVALR9ic5msaZ8
TdUdjlavLTfFlSl59EBJXVhcyasEErxpiX8ZsJoamxa3FYUiaTu4+rXPS9VUNFAt
l9/S266M8DWOgqjYjFv/v4VAuC2ad+RDGYGwwdn7/L2wjtzC35J9uO0myxfhiaSJ
lHtI2+ffB/PD2Y29WCJy7bcZ1nJR0hK79/me1b5ZUZvKt4kaB1s7XPm6BialSzay
uU+JIBfqKo3Ytnzq8SAHl2gfPTqFqq/IYbecpHbgW6jZ5VKsp7XzLelEPsCb9S0C
S65F0bu1ZIXsB/+OARShUrKxf8ov+nKjfdYrYG17RtgHCuCGb+d71yKwuKvCBAnt
mlCX/4ekeIZSPCUYJ9EIu6iZSMX5VhXsJbdw4GANTbI0/jSDmTTBf73IKZ0Gfop9
3bsOaHjjwmdDdOV5Xhjg6miI4ofPpLFIzZn7MsW7mIPa0rwia8Ten7TiucOAGFto
4JCg2XyprNrSRncu8fAwGk3IiHLKisL5sjaeIVQdftTm+k91jThyGUv8s0y43D9V
BbdmHOlMT4Rf01tWXp6D+ZterHlEuGXglHDlAI+FW7YdGFtftXb8d2QEO4MK9WQX
ImgF29PruuWif8/SF6wLpQoUGEBkBU3Pl5ckxx/BxARgv1nfRviKVgaxDcKxm1a1
JyULUrdhwScDmoBeKb7+qUuC5sxHYbP4sQT7oQTmOUZ3+dU22+VH165iGgbWw1gi
4vQfww7O3dhniSvi0fxacseHIr7D9XrhdTy4Q3Vry+5FZr++WrTqzADh4cKO+71Q
Fh2t49AwNczCN40Fbhtnx8z5PmxLInu2vjbUI4J8mIaejkgmPF0tIAsn+SjRx1uN
aATpNJThfn7LNvUfMoBVjDnKyJylUN29fHkwSVATT0qW4RD17wwYS/h5UZY80ZJj
EP9mGH6qT8lgkNaOPEsU1UhhyImR1IzjVS69BjRkTracZSDtc6IQprNqSmmEd4Sc
K4wtCJuFXFi2SsNjpPBmGBeqTXM/4pQsLvVtjm4pdWmGdxS4WY6hARPr5OR7PYJx
TkIZMHhHAJQYYUqm3eE81a4uQaNptZUBYOaXy7qyp3o9rIvukVv9XVhCP9q4j8HF
Q+k+49gcU22eF/1OrIQ9PaJSNqZIzo+OGgDiK8EoN4vA+zdwBFsJgu+GNA8yH0XY
hHssAMeydd035fW/DozioEZFhtWGXP2AVk0BdThwy7KlVKlNLOhm8d/EDob1bbTo
aDkGYcTmuqN4BfhQ5EiH0noHF1EQ9w+lTnsvWS0j59NZHh5E7nszW8T9h5KXmyTS
J+0MmMQJ16ePBjol7kVQRBuxm8N8r7BFSdsFvDFgyjP1AMp3iok7Ls785wrsjzYC
IxH/Pz+YAoGbi4318naUMR7DITw29phfJv6RLLjHMNAbbkrKPtXrD4kzVSAoU/BI
8oUGLEd0L22MGq8l3Ie5GqkKD2nKOQZseka4X3seFzDTTTHhcihLvPxnjun6EAlq
2kzVv8fylc+NEJHHuFMES2Z75EQkyFvAirxGnfR2yhXMI4o6ixr3yHN9gBsTqG1L
ygX7ZkViVhdwTqB5+z+QdBMaT4KyIX170icNuB2eYeQglaBN5k7uwM0t8wkg9gg5
/7MvTrs72TIf38ZFmTke0bmSFUPnpcByQ9Belfj/CQsOzHIKXE/Op8x+GHtEUjIU
0/NHi+dysAR9Q7rF9my2rgilJ22jLJm3LCNb3GwvP+wxrTDiEMEK7/IUzTpTDkGv
SM0naspTfPQQg2GAYT+WO/VR/ShUZtqDgL0LZO3ws0fy3AjRT0kmrxFENyt9iEVF
HVG/MPQjTbLwXoish2ZKn75+cfBg1IB23Bj/S6s1ykVU5fWhe4gS4+pNcVSNYoUs
vTJ8sgACJr5kPzYtHzJ4XqUKqY4/kIm804yLq1zsL4lPqRAgQ/VICcgNj/Mn2MvZ
qs3UfXxpWPXx618/HdVi/Mm52VK6kFIV7oNw2sWGdB9YlG++irGzzRIU8GOo3GeL
lx8y6ltk5G7ZlGV9aIdtlIXXfA2ok6jhv/cjLZ4JaZgVdVyf1ObjWJGIGyncul9O
9+APEdhnjcIa6FCmfRLc5SfWDBQJqkXp0fqZxHz1j8N8IWjadTTQA8WR7bhv0KT8
LF++cgth1LI9z/+qQH7YEyMEFdi9DFQzna7NDuS02307ESK3e6zvGvoF/x2piDJi
kY0rotrsZePqdEIy2JrOwUNGlFpgeCYmHLBLUAaXwcjhb+PeT4+zByTH6ClG0kBZ
rwEcFg+tQbYhoFw96Ez8ZAY6UdWr874DBrDgbwBxsE6yE0hXxyEpsbN2G5u++r+F
ZWZSuF2KHAd9ewAvm5SMKBGPHF/OB4gUxZCHZk3f4xuz8hwcdljBNZ7LnPWSNvUz
I6KfFZz+wVwS3VWC1UZ23pNa5Ft8R5fnzO8Dk0zPK1R55pfKy3+lrYB/4lVYTiJw
+WUA275vtNUbcy/TeBi4I6njV07pYkHDDVI9hXztBDRP+rX1rkTrxKNeHrIUGICm
t28AZ7hJWY7xO4UwM8HSXeB1RHtUS440Z4BXyQWGNEYfAE3i8qU/Z2+ul33lGAoJ
dxzDBv9nwtycZEvpsruCcXssJcJb94f22IWGcKeJqhaxgsAOpUB3cxr1/VuZ6XwU
DNqyn9R79Yu0syB6hZofxWGlnRik+ltJxm6SLCegwhm8thuA1aArE1Zvl83B4M3M
q+c6rfx5RMcNXvU5AI/OE7gt4tTwmVUhhNYNljlUsXkke0L+9xyeHwpppYQMK6ob
aazPCzlPEhRY+gooD5DHUJdazBAnQ1lrWKn0Rb1iR30eicXBgDHTYLywU3916DxJ
MZ7TqOYtnkfUrxU4M7lWgKneewYNJdAlFnzOW6XnWies5ISE9UaeFPb86eI6++Ub
RFyqb1/Nnv/FvS2EJpbIXJaoeaF9MZLPol8m0PMM0Vfm0mScqjoBlSHhHxTukIB0
9pEx9THj7H0VfZPm0E7Doh1tPsaU9xf0TdIqZ7+2Zyhgg4T2e1jiRKKkvAFAfKbS
na/qTltAZsYwgMEaJMFh0WOpOI+pAFvvS/OUtP/PoeGSdAFaelL67ceGxZSOzq02
zqaDAZRD5wXvIqEiMoftAv+064Yx7bSyvE8Y97/5SwdCScIKrw/MgEyHAmQIFJ5h
EArXLKPUEezwRjuJCt+HbnBG6xobR7QdkkjdOGsJ7NaLksr2qx/6Lv7hf7P0+nGJ
hggv6kozuB9IXAaN/IQOCeNfpHA3KXPeeTv0GOK/WquyATXlKNLJ6Ue4lbsYmSAc
0IPmw/qGmV5/F5TWQ9tUvsf8nG7A/yBevjkm/3HR1h5AvySjKUVYRyQxwOxUiOnj
/lcxegiyr8hfnz6NxJ+yBZRJQyfdgWkaL+EgJaXg8x4/atJ39nld7XhJVtVRR87t
MtDalq3jURapZUIFK8AVMeMFn7+mWflJjgUHbW5Ag8OkOiEYWhKR94xh7yzNwCIc
nK8trDn2EBMzao26MpvDMyZPWLKvmu9UI9Ac9tX4X5WMkvV06u0kLwIX9y782aFN
tVexZR4LBCAymS1e6Z6eLhd4+vznZkAee8iLqQB99uG73NDGG3aWkSa+XooXrI1Q
SWTExRrtpcKcl2T4Bz045oi4RnbylJxLiYNw5o62YmD1dZ5l0domXoX22Ost4r7D
+Kyu2mVK75nLINpR3AnsjWXuEIroPdmdCuSsOJDIRqC4F+JqOo0GfrjDD1JW3lDw
0FAMk6XxZgjQR7br9um7QWycbojDvspzrYIbABVzLfu3t82Abu442lgXiaINFFwa
pMndbXIZHyo372pBLAP3lmb432aLk1uxOqNxUu8WZeGV9Lr3TzXWEe4wfrpCNgX7
StmrZWbZ9cPWF+lofBqIUv9HEykIX2MV1s7dvXLyXAKwsrSkRcnihTBywt+uXSwG
OJHUyyNWmVkwUQVyScTt9FWb7N+RsebCnT4uYvtDjDfZ+qbLU5EQeBOxuqIMixR0
CXMoaMCVyKhSSYy+0c8M+VzeavQ/kpJgB6jAZ8FolHinJPoGhzJDaW2mipFrEUzx
Hc3V2bbWLny2vfo8NilklJdKnE6vf5/fKGu5Z5UvRW01xp4aUyWV+Me/T1oSHDRv
3eUz2ZM9aL4oSG7ehC4JF+LQDFQK05FthgdjdvH2mrkbbJqOSXFW/c0zc2znPQ7L
SxXQ5YRtCtd6cWmNeBD6FsQS85FbboBkqXTJpcicNOeBCbo4Kenwwgoi4XN5Jk/0
gzdCmuA/TqHqmOdujO5033HDM8/p1Z7q3SR8aH+E0BnUkd7IVlRI4hxLtPVhkuz4
3RTRX/TPIy6DdymWzZpmdpuVIMWH00NRTaiecrJRW3AAKesB/He7oKmU3vCkW3Vy
NTKV0qTHsBB5LybTAQUjIu+ZyoPxgNWIENlVPqW9N4a0N+05u5KfqKD53JPvwElH
492g/Mx9iDmknfhVLmX7lA+AUAMSaYkUkcBnGQrBccsIfxiSuN91KG+UTbOt2KtN
724/4KWAqRMUbstz47KroQRqprtO+H4sXojNmUVKIkytvnCjo9O/ugsy7GK4OSUE
UuEJHDcqGDp7kvkJp17DKImNjrbuPhgCD8KcGzEr4cTCPxhIehIxaogUX17FWChc
/Wa3338wqpVlplW8jWB8SLupBG1M2SlZSlCxk41Dy1hBiD96yDlhCN6CTf9b+3Zt
SPJnlEe4mV4MwyySAG3z3Wp/350enil8ih0+rdsmvZH4P/andDKRbg1fKhnDwY8J
ZkCq9lxPEhWBCNEcQ9ALpVgF54s9Gv8krbvNnBLXqAUi8meYuLWfKrhbUbcg/pKG
87ITMhfr2fPygxFC9t2ESdiDo074HCQMcTlOKEv3UzFbrBnulZYgmmGbVf9uwabs
f8QXo4wSHglqKp+187ryH6Vrt2ayKu9dhE+Xau/ICJcwafFFWjrOZDx4t2B7uLZ0
siWo5diMwNicnyP3TV9kz68Pp7Av1ua/NwH71ga0rktuITbJjXoEQmpbjLW9TLDt
O9vLEf0cLikCKlAke0NCYXH86uLJOGhWlyszQlWp6M5WW7yZBORjKckzrIQ6Tlai
9d2GZB2Rz9G9ROu4NpDZ3GM+lny/pnh/oT7zHI6t2tojhOyINBfK2DQoSdxvwKpH
5EeXoVvZDUyKuxqUfPbR5CRSwdGXU4huQSsuOcNtsakMHbo5tTTL7kCxAOwlGdYv
NzOmk4VcqpcKpX32NiCp73vOWyKTbUUR7pq93k8olMLp0u9SqhHX1Lze4rRaJliq
ESpRY7MtqAgEjGKMFZU9PpBwebz+yCfWdc+llR58NBKl8l4vD9PM/w/wtIVhOP1c
IWuTs4kOy6SQJgVi/06LlIiFi4n15lJTkhuq7YuPOnqJo1ItRLEZ9/ISMPljIYz3
eh43y4ZHEFrVvy+ewpAVsb+Uiny1a93kKvsZ7aOmlvpJpxwm+MTzgoPcvV8bxe2B
Af3WXKEjsUcEUaL8jBLI6K2ysEMFALwPGhd2XCOsfdoxjqhGpGjZLZ72TieFAted
iXX5r4fWV4vHBYVpybQgVIkzDYBUT4+/dcI/jforHH6dnydhWCi7+E0pzaSXxO6M
vrUo3TQw1cG6w120zE7Upq3YITDVjumO8pvMSN3rYIoJrmEudBXH/569xQm+RzAv
ArJADWhOW3LDLvWdNbpUfgjKcZMpzmk5fk0SPQRC5fj6FDmfotQgYOpSUZoeIQK/
KEFAmPOZUEOu/3pnzbm5c9YRq9brCXgwt5Wavg8yvjJQISoRxibpuY760DfbQTIg
Ex3Sq4bEqKFHOJSPGlu9Ugs0HAgM9Kez/4W23KiIi90JoGcYVPhjFFAmIiKBpog2
OGAu3cEVGnhLrEEdK2x/GVfjISpKcM5e+iIiPDa920FX/BN6SpWXfHGKLJ09AM+b
R0okvcbCDkVx+2DzQwPzGbpvrgyw8gfbojEaUeXRpUGGxkDFz8mASUaA8gODPQ9x
IaNPJIlNaxij5nhP/1P62l9d/eX6YwmqhfDYp7YpD2tAP3iQvKjTj5KVrry27Irp
S0z+oSTq0H1BTYWweu8BNgXkMIDlsO9uQYa62Pv+yLxi57ghkTb+lcMKs4H1fEmw
Z+1Gkg82LlFeox7/OP03AtgkIdfPneVKbncfxH6wb/2Gr6iQDzpszQTKrxKZYKoP
Y3IOvP+1vqa+8mB2VlMiz3BiQVoWs9w9vMQlM8yJmzdMTl7EdCRBRVnXfI7BQgBo
JUwZQkxlJAq8sAj5/A4pozZ0C42ocrohI3KjqhpAoQVREFJuvcViA1nBsgGLLk50
CnwYdsHM2NhGjWdA5sHhvesvsZtNFkP44rPs4pahMqzKEvv9SLr0h1VuVQQ0fw9Z
PlpBqibrW4Gtfqox84tZmyQa82zMa+gXJidwaa/POU5LRBecA7FUZyyzjJgYC8az
krVj8aodrYv+oaBa9P7peP5Ahg8LN9P+7qn592cq1zY2rQ1Tpby1HFu3MIycfOkd
82QHZx0i0D4X7qiJoZ8TldbtnslMH+GB4h45lEWU5xwahMPmJDpt4HZje18ChP6p
0YEnbWF/e/F4mn/JchBjqnY0suEQcddMwISkySxc3sgPTUK3A7vAEw2PDdWNRGLv
YOnTVofJQpw0ctOVkeWxEMpiG5/dQVaP97T9BkfcJiAimHY9/4RFo/6Mta7TNBqR
ibrpR6FBdAgxCjwND/CoHSQxYhVFdRCj+iYeJUUTqDEMQGlBKdRdmNBNcjcysDSG
9nQX7Ez1SLWUSAe7hHUyQZVhQbrziZPbLdyeKlPKkKCtdh4QTCKK4KgTQ/ws7GiF
q2lnY4+/QkJ9a+iOfTVxb00zyRvVsbCw8H+xomVxdQ9RV6Rn9+spp3joxm2ZKqiS
ps8mkNSZvD/GHYSqs0hC1ZbLO+W+FdBF23RDd4674jietf9uAebAP/bXSPP+wj9b
AHuXDQ40yBKwbhm4yW79cJBij11mmSGvS6Ev2s0OLp6EGFaxbGZo2SXhYEugMe/b
aL3gNmbs9HlJlyztsmCElToSS1ffAk7xwbTIeN09ZURf3aVeW8/R1wUlBcpmHw/l
tMO+0KNM9g/FnrsCMWhPSkHynCowxSiaIOxrUFfui5XNZ+xrbYbLCn890h3HEAKP
67C2SOS/dOHxPW1qhbi74/e2Ip6n1BYvJqdLnjirj4nHdiRsmhrQswN8G6BOTeMk
7Nor8a7CET4XGANBU4o/Hv99Gej704deqwuPUP48QMBI9seli+JAV0rmaNk5DZK1
+IXgDVJMmqQCAPb4ApI5qn81Zj1o3MuRx5Z0LJWtZLJeMWaqxmfp1OY3IvQuEU5z
TfOSTvmGnQ/3OHw035CXPy2P+nSdpni+CW/O5+JBjkctnc4sauE56jcl6FDOctEe
Qs+GCSR84UDQPbjXjcmt1sYvhVvbkdAeekQCBwinM5HrPt7cMiB9xmATSyFvsCUh
IBaS0qZbWchnwmI8wWumN17Zf4MPWhDkrW8e2cZ4TBM5KAxkt4PRfnhUH8gu74Sm
AXXET4xUpZ+rhwzekqVo+8iKi7vuL09wbI9Q5XJId2PFvywSVBtdXegegGs2kM6D
QJDTI99qYLhAIjtDQODPAu0Ni0l1A1qTQo2IeXz4psbp17oklZcZkBwXOGpCPXpk
44fyt+sL+2f7khEHjxxmXrsVRA5u7INL/Yh87P9yd1fYXDEuUX10LlB3iwpo+4IA
miC00//4BA7yDgOj5ohUG6BCvk/9/4Szunif+ZHFj/wV9s1b64gMpA8HLMiHb3GA
MgL0HOHPX26VEfoDTZklnvwogj4/THcWq7mB8IPm0+dqh/IvP9/xbPTVtzSSR24g
GZZTjBDNtgAuHAVkeKNEt5+0aivdZnbDo5FHn9tcUuM71Qktcm0Ss7ludj8fgp4c
ZhnWRrO/l+4hJhmclNVj1emy579aS+qi1hS5synzI3CyiTgUXrjyB4f9LpQu7W9O
Nz6jkitjK+dsdYUIrkz/ag6QJg6FMqlnnOazTW+JCkfGWnGci1y71cKnlDFldNJ+
HQ+W8pIHoT9gyEgMQ9+pSixs0prt6u5zd7parc2pDJ2IneAvODM4BWlG19IK4qmF
QXgITiJ5xEe+3aLoiDxTY+ATJkHNx0mQwg9ixeImdPxeiA2oj3+7iEGJw4HKJqgr
rtsvpwEsWGd45mNkF/84b/4d3V4zBpQ1UooGE8RTlX9xaDg/CTGIKWN6M94BDdQR
2lB8ZhYq+h84OglRfQnsdBb1+rULy/Bu2iAuquC/9AVgGD4VL/CBMz/SomkrhA8e
RAR0ML+yXZ0K1s8WJHNx3fB0Pr1gzlNN/hTWNBR+kg53B1HRFqjbmdLG1FF3jx3v
9S1DgrkY2jD6brMNRzKzqU3l5m2e70XznnaWfSglx7WfUMr9GU19k/dxnMyS9mWU
JyGal6Y7+wMvXQZcWZbDRkV1zRcmD5ET/YNH4KHfG4ZHbLqMbzInaQ69JVEMWVWd
CNUA1B/sDXoyvULby1vGXVhd0ua6GGH2ayrSqxv8FoiAWwfPqtH5OxcNM7odK9ZX
9P7qsNgO+MuqYU/Y+Pg4Jf2Q/lL3XwhXymMYC4VDgyvY0dx1oXFLXWnQ2QAS/Yh1
KN0Fjsj9FZ9quHsFb4VLr8qKjTGAIfiyyq7L8vww/NltMEzEJer2YqoVAznVxf4l
2IoHMlc2bAmnyy/XoBwxoBJoT3A4XsHJGgG5j7dZ2XzkB5xFieYSFx7yBR9DKDyg
yIfku9RhMm2TgbEeLpOIeeohb40fJpCiV8xTrZBlpiUhe7SOjxDAyekzxxoBkRst
xVMSLBvoHxGzIzh8MllLsm3mDVubOAZacD10GIVdq9C0AF4KdSR6TyE+FZnuOJPG
HZnXJcgsSid2tdIuMt1AR1O4XXRoL9Rik8YpOQPLBDkQZMygMSDwNzohxU/ZRZDq
NXworokevnhWebUXlxHUqa/47+zhC5Q1e5iP2+immLzAs/rVgAR2eY2MW5EhqUlG
YLs7tYQwDC9DjeQLcAkeOQrx26dcp2HE8Jmx+tPje3KwwlKleYdbnYaTFkLltc0V
p397MI99XNPSqeTUsDvVzAuLaIDckpI+tGioxnvhv3utPRCSkyhaSs0+Gd/trD36
EabKJ4Df375TOw9Cy7QWgRRve0K56rF3lkZ0kBw3r1dWR1PcGJexQ5Vu3AbcEUFr
7CepNI4VkuCKgFmPS1QIS7BB1bqH3lyKpXUt71y/tk3HNgmSq2xgcmv15P0tRW75
sB96IhhYkSCb4p7OTUGEo4F3P0+Km6ZrQgTxnbX/0Ywo2LIaySh8DE4yvr/ItYAW
rsXZ+o/E+Hk+Kw5RIvWUlD1jnN1fY/CpwQsaNJuU+XkkhHQmSHKHAO4vPyx3XEwt
zzTiMtMFSw9tAFd1rWtCxZeYut+Ow9/m1Xw9E9l342sm6KCDhEHeSKQgzjnz4HEO
QoS3buFll3OZAx8h38vxMiA9qKtmvhH0nho6A0n0Dl/40qv8fXusX6txeOpUtItQ
Av8uATtJWDE7LeLO1eGuvyaYA2CXJzNVDi5kx+LkeoPR+MEl4Zcko1sESxk8vKNG
3QdwwqYKG03R/Wu2uI2KvHCELs62lQpqdalSKGnUWC99lX714ENAfROoYJ+axpky
/Di+kipvV3+KPzr+ptQWsIv+U3RuQY/Ltb1zyDz6MxEXw8YVRQ3OjZsREXTNi2wh
cbB7H0Oyyr6vKLGZUfNAXbcjHUbc+mbGwrR0RtXBiS02gEYE3Fd9y2B5D472KCYI
0BGV5ahSrTfULilgc+hcE0rGVM9DcagY07zA0DQygFYW8hV0LsjC4e6CdG9UxWuB
2GZIN+Zq6Kfu2DgnIybeOZU8cFhHBNm1iRGirHrdk7IdkUqvZKhvI2DEqpzrloCK
8dwncSJRPP69V2E199UHaabz/UXZr0wAA2ic/txIcTcUNsDdBn5Gj4xADKWfIZ4k
w8//hofmmsY8ltoIDXDlkTJ+ZjHe5gTHEdmSj8JibteBFv8lj0Sg9WOqCNJEXmPx
xLAPsadjplclOCklGZ0AvlER5PDi3sTyoTiAKRKEjR8S/nuEKSM1hR2+zkmcPCmu
Ch0q4eeE2BijPgroRTK1iIOH3p0ejQI092qCoGuBz891Eudt39a/8z5DpDtU7S2o
/S2BlI+tW/XRRINeoIoE8GyaUUvZdyRQ2oHxysb/ZT05G6benBah+Gj5VzLkHTTs
W9eL1gnMlVDVrxKfPTq8kLZ5i9W3I6X/iKt0ilFLzXZy3HOAQX9HoyPjJoglTcw+
mHjFs7WB5K8c2LnwpuAEs2yQPYaIh72c2+iwwFNxQRc++coEF8PE0t3bPc0l2Q+W
xcaIA52DvggG7ga9B9ThoXxQrERG4FGF9jvklrYfOvX2+/Zk3Fr4HrF9XPrHBJGZ
9s6vzv2mgrBCCjAyCPRMSudhhtyVzymTWkVi/NND0qiRKoxJycsaJ2JRW5fQnaxv
EIeWV/2IVB4XkARgSKgKiEQOuCSELA6EKrWWhK2d6zBfj/3s3K2LZCgGacH0jZMC
rv/f+zjS1/y+6x/RtEJqSE0h03JS/IUuLmwELiCx1nXaAxUa5nDk7HfYtOxEPxo2
yGVbRrUk9goYdRUOJuOH2lQad7uhQnTVWDJvwkL7ug2WH6ygrpUPYZTWlPQmwleh
KiIPWeiuMnJhOvGeST9PfPeMAZ+09uyFKv3KPRVaOdTF3pMSShTUlLPIsCJMOeg0
tj8MjXpf0maaAolKjlGZ1I4bLjSrqI7i7H+/VCrJvVBWaheIfdc4TaXqxUgmgRNl
28g2Eex44VBRaF9/mgybhAJBjhQU6fJ9FrH6eVljrc/P4cekFMHMBpznsvHRCzdd
ph3m1TYj9AYFrvPPaWW/eNtYZ0P6F3JeYg5HJlaYwCjQkpQx6hJ0f3L7t3tFEXd3
3w2gAQ4w3RGUqykOt35JLPQz5HPr220CHWd5YlKhmJjCuMNjvjX/W4DJdBLS3VtV
x3YP3Z7OK3YVohqlws78HqPUPAvxPgRE3Co/A3c/MXxFKqoPPUvQJd48rzW/kBdN
TQMI8NmIbzXsVp0CT1uY9Pl94DsigjAS9HjJiS9H+XCEVpu3FqcQchgVP4Y2KNM7
LPgJTMxCfpVEWHBUtnK9naw1eUKBa+R5DFP7/iXbklxTgEHdB4FPNk8PNk5KLSaS
gikL9uyaJA5Pb0aeDM2KuQPjPYdyeiA8qpw5FpMNA6wCpG0vghtY5U7/I3MCCRwg
9kP7KFawGtm547xzn13UduZQmb6S1vLthQXZbbgxlRJAgEqzcrmUpPqGOQ946TSK
9CUESV3EKSLu+iXGUPq2VoeOmK4I/wD4oMwkPC18teKYgBWApCAK1tJBgl7UsN7T
iZUaYRUCprHir7NUPgMRu8A5lvbDIM4jmcPhxMzWaWTkIMTXDX6REIq3TPtJ4euj
0jXDEkHo7W1I3E9B4iALTZ+Twdt/FFyeC/Y3JHWldeleBbp493MFmIPHXf0CutFC
URGy5LVIJAW5+tpoI8k9sDCGdIjsVmtqqcsLNCbhl4GG8JlsrWrILjAf/iO4sfnk
JQBRwgwMOrNy/NmdCO/1Srx70OmFXrVc9eatVIfp2eouXeYcHTeK4MqAonOsoZY4
sxU4wRMMvpTBPbnzKYEJm7qetWBHXX/dY0cmRtgUYHMmXKozJ2al8dYSuA1gt4yM
cqktkfp4qfKqxCisLMNRXcxeT/G6nCcXUK5F89AhYPHtCNnzwK3Fp0OtXEIpSlMr
YTMia4AssnOEMofVUTIOruFnd3cXXJtpG+S/TOBFPCNKAEvhgYj+xqMTbR3BlY/M
wjqb7oJoMxP8SBF7Fxrq09ljQgDo4rDdQGIna+w19xnkJC05YvmnPKYTmqptcZkb
d18v1afB8qJ7lIYt5j8ku5ctkc2odMqBEoGCWtlT48mXoRvnDnopoSZFs/goJ1U+
RrxFYXDR5mM8l+2Eb/1YS6ACZQ3WBu3j1ByufuruIJmCiOeQh1WT5AU4yeVlzDAp
AJ+PwScGwpbSE+UHvZRuFrF9bv0bE5knKnDxetKhEOVaYxqUmOPXo51LqVDJwlqJ
cbVEhJSI0DXGqbcovOkRaakhpeVaYukvIFOhqgsfek1rypV79S0Eujbr9pnL/1IO
t6U45lAEFMJcsundnYXb229pmFhUKAgjhbAqocf8v9wU924XvntArEvxtX+Mg/2H
DxqlAVumknTBqRiJ0qusW7m6YgW+NsolHxsyl3S/YHPtfo15gop0dH+oZqs6xIhy
K4z42pdLaNAb0C8RLyGNHWmBGDfe/TvEnDhEC+SAAwthJ8lRQb4eXgdhM4EPsqVK
Nwiobh9atQ0bJNMTjm4OXwXO2HGRIdLKI1yQqDtedLHJCSUKh3sfEaFUdO17lLgE
Tv8KVPDsGrJHvS5fMCoz3zBZ1r4+9Imjeyiyb3l1FBkj2ID9dlihMI/xqjqRqpAH
34QZoQmcqZ7ag6ExrXox4hCxQNa5G5c5d9XOp4NpFWr5PIJveVoMRUTX+ukvd0qO
bfEF6K6e8G7KJDtzvtPySLEQ4yQ1O0v04Fp1C03GTCElEFFBExMIUMTMr3olSXmz
2QrH/Q4/58mhlk0T/uucA0WhC3iTfUoGYG0rVWgYA+VSlJBClc6Wp87imlFAyTKP
pBso/9wXKq10lrt7sXcL7lyVzYcxWs1myDSeFyKSzWMBoVwFoR23guNu+PPusI7d
LvEh52xK/llPiyR0DOav2VsKtWX0Fw2X1vteEZkroDBOeqoIWnp+szzq+gdBx+xu
FeJl28XcAYy8uXm1zAtTERZHmpgV8+MPvoehTLQBN7LFlmrTy3kNO2HxWi0GZjh5
pR8dhckHYBUa6oXnlsUeAUlnCNtlQqySVrIK7nPvhZA6Qjty7FErUFxwk+48cNLY
ytkS1S3J+hcIai9jl8vhSphQldGyx6mcMev1u5qoynuwOIEQjNpNjmIAbjjKyz3n
kLa+D/6+F3foJ55cP5DYtRUyptj9GpZ5fkEOPQ4ZA70enfKfoKALrDWkUdXDmKUe
sOEbSsaPNNp8m1D/ooyxIfi5eedfaZO/kZzph8FhLGndZ6h5Ow4J8SuSmnpd7sJX
oVnOxkSyhphtgH9pjYi7IUe1sExKz9kL6UFCgBrP6WTrgu5OQVmNeJ2OIcHruj7u
e+OF6198MzRbMudadLnY4OFWj1tKYqGpfdSPybPgTjJ//Lc2ytm0xSEOmWiTlrgi
jBmsP9PYLdHmZnGNR5fni+nvAy316Yj7SjjQuYppRp71EsrPp1TGDj6wm7ps6ibI
mziuMzCglDxrj/dKarDx7mUkHWAX52EzsIJwOCnu5QKAv3xXGb0d/Ic4wfbJC9zn
4orte5lHcZpXtVBUT383L6TKiIavwwX1Y6ZGlHZHOg8R/vxNBCw9XReAkMZZTx5g
XS4Kz+VSA8t7jqB9VAUB2kUq5+j+rVclYIsOaV9d9u4+2jSpgEFCWgdUMnGoWI9W
GLrVBXktduqBFpJ9EApfhR3s4SLRRq1sETJW1iqoHOez/EjKBybEVvU4hHOVIdyi
HFyjs5qTbs5XdBszihDEewRrSFlT26Fd1x3BqVYPw+3+cQ14QwqSSq6nbszQNKZQ
OfQ3EE7MilGgoI6DMQmEoOL9hiYMn2eLZlvvuc676GY9jTURYbgQO1pAp6qZNFCX
92STZJTvhYNjeLwETwxjUTmXBhsHk39r2vc7rQEW+fNLoNYJN4vvtW5s3ws1V+bo
KrTK/zVKhrKy2vXIuHT0Uok3c3mijQceLKna4HgGgqLmabtbYuNhMAniFWHLCteA
ta/1rnN5gX5RuRrcvKScaoZQBQreZGMu07ZD/sfwteVhC6PiLx8ZXSi8XrHjrm6c
7F+8BclSyjjup7Jajylq75UKwZe6soWk7STu57+V11s/iBmnZKsUSijF6qzuCry4
c7QqWtt5uREQsNvkonrqomt6GTh1IlWIzWaodtRsxgLm5dv/kej6oQ7z7DKRzGsi
xjkYWxYykF0/SPj9O2sVW+/BpUo0yoBhrAa3ZN9pQyYNUdSOU2pNo6/XDfCYzzyt
9fvB1ygH7ewvVfuHCv3+5LhFtrmmMX/RGQajUfWfmKQWD2fNI4MEwV9dP4IomFK9
8gt0OyxiK7GwPhVOTlmgYlrlUWAMAGu6+SB31ldC88AntUFEBzqi0ovn0WQwSeEC
9HSO2raC8NKqxWhbwcx3WQnZF8fqTwUA3MqMleSar7NwQ78jITpRMSqXOGaKrKaU
ErQojILInYDfOoRMIDNpA82TW5G0sLwbvggNKoB2Ku5fAmjGZqMk/Mml4ExwEIuu
WnNrrAsWrtz12lbwUNZ0UbVosvckngUluJjscnQDsq/SIxeijVFF6dfwOF0wN7yg
WlTwI3n0Oj/tNle974EBfP0ajGsGxMz0Qw6Qr6yj/Ev4F+2Hs+aYH3OlRMO+wbct
QofSw1P7q4ohZNJBM/oZc8UOlYQAVDBEc3Q4ny65nR/YZ/9jQxis0Es7mAgQgUTR
vg1hzJxF1T0gD7zvv4tYlEXBLlbtUmLXPwG/bsGA9eyMBwpVoYI1HhvAw54VnbTm
NBFdWkQbCmMYQPFIh5LB1iPmt7s94sKEjrWb6QkyGPLJe0ceOEqravNQ9GaD/fbk
Wrh17OzwyJ6t8il0ttaF4cpV63MgD4Fvsk0c8hn7xq9MhQilsY+LHl3as5a8EXUk
bzS+1vM9lrc96XXlj8LgHzNHe7le5s5NyqXk2m8l0UCxj/ziTprpZuSuOzxdHc7U
YyKRlTg/UGViTWzUn/PqACsOi9XfazVyRv51mrrhJPZe7cT7DbPvOOGOtf+ffXXZ
qi9nq2LaTd2MkuszPGhh022Y3s72tj2MYleXd3lA7uDoulAAJrdwhw7PKaAtLenL
PMjHzL2xPZ4F87YA7c/b+XHuqfTVaW7btc6Fna2eWnEcIAvv3zc4UizJrJiyQZ/D
dOW/TIHYR/ZvyTgXn9xEB0lHnF/iqI0obPkiC42IJYXacw3CERTA3ZeE0tgThhzJ
2rD8+OttNRGcyhg8n2rssKQPiSy9uqT/5nFOgY8C58vUPRTLwl+SH+JTGKooCQsx
TYPnTLDR5+q7cQlUeLflsSE2jqSVThPpwTCJNApSDQiBD9GWNj974AaZ9pj+dw+S
PNUSwIggLGbrPgvrUEK+S0tIMrjp/kAxB7Wlpc7VCvJmnk0QIAng1uROglBHpYsx
1IaJMbGuledJOqT9u+Dvaz4og5gz2dK3GPwmYtyVGkzcndPSN7S4ZctFat7N/5gC
ALqv0yKc7NhXsEN8tq6IS06C+ievHqKTx77AyTq7871nRxyJFdRs+W622zte9whr
wCzNa3wmFiz+Mwnc+qF3FkPENfeYjkY4RmMlsd5AjPfhOurkR/xAR+kdu4YJL0ma
XR3ME7AMoOslQb9frnG9LWp+fbcRUz2sIqMz3Oes/xjzPhaZx0Xyf1E+rDPsJw2/
AaJiGQPsRaHcQGeGKQ+JGXf11Z3kYE7bJXZbYp1uisOOe3KBd6u42MetV6GTItxP
ZCGEYLPkku4sJ0pduLY78fM00jsmYZasRhyTFgALFGjl+yeVc5lagaCqx/hLCFtS
QREt6ZCqSbPNjT24c/z78E10KdlVtKX6r4y1qKHHPeY+xCF3Z8ltnsx2peFh3eS6
AmtesbjfCaJjEx895jeTZjVBFRdkQqAIu/fWS7yQFwFrm472FAxu7FO5faVUta7f
d5pqTxHajlB/LvZ/JWhTam8uTESq6szPT3i6pOCR5tEmYH5z6w+1dLWOpNHNlDJl
d78u2f8c5VX9i7Sm6K18GF+cleaWUKYK5YK6FLXcHCH3Zimw63dbzcU20aVOg1vF
r4nU6cyCtGypDc+Q0mb6aRnDIruQn5GgPCxei09lVICvVhlVFgSnh/6NAP9gUhrL
+FUTQigBM8Od+p3w/tSCwPfMLhW0nj7mpzYI3r2IQM8Al5kk9KV4Y7jsT71ZVM3+
IfoII1mN3/r6ZweluELxuPBo43DrUM8M+VmtMylN6W0VaXw8XdGHF2YiaejfP7z0
cUteQLa+NyBDZennrnNf19WqHs4l6LiyyD43baQYSkAcfsh1vEojp0VcOLc5cMfa
of1+A3GiGGuQ1ZNLJbo+an/IaneYRUSmWw8gSPVi5HkHFlh0hZbXpWsE1aIauz01
fk1c/0s5ku8Lj6c7QWDn0Vay1uW9R/u664LAzwSnpzy32TPedMdauh1561rPuTQl
2kJuLFcVmJ0K5ayW3Rg5YXLpMj3ZiKp+4WkVmFL7xXZWm9X1hI3iP2cIXgb2vu3x
/0LchwNPsPyXI41JmbNZ/uj4ixySMwPiDcdwQy9b0SxJR1hL7g/6h6Qjc+5orDxV
pSMnE3aJNp5AQ1uyPjfO7PdgiTYT1Gq5UNhEtJcSa+awv1A2CThMG2CEGx8WIAdc
MOnGQNYZUmMu1+ZwXlVfi9VcJl2g0Q29xN7QrpHwAUxrvgyczXtrHzGmQIE7K1tL
N+4zHQpgj1+QYK7EzoaSuRu5cFlPGWMPlH9gv4ZYmfANG8Yh00M/Wz4lNPE3fadA
2yyK+FtHs/wmvNlepkRsVcS2PLd5p8PlT9lP2Zmdoo8N83PcQunyLpgaabHFOmxm
KUuTHTEkP6vYEUuMCWIlOYgtpgaTQRkM4ZsNIl5X4thxTwZF0amxjtbMyoE27CrB
knTXFyqqxUnGttOuGErRGBdzVIRtFm7xZkJyxiaqrQ2rhufGRV+Pokx4P5izwwBk
K0f7xnoZOLWSM1FwJy61NLrKWXY8vyqKggASSn6PJ0/rTLF/NfS/W2Q6VD1/heAm
t7fRJ/2yy7WtQHtodYUY+3saM4E21J/OPqmeSm+GYAjNBVT6UPZN6XA5Z+2jvPjN
5FOhpRTUXCVx/M55yUdZa89JDo9bZTZrKIdTtpgl1n6Rl47dfQVHido1GSj2QX7Y
S8Tpftk3hW4sLjjPvE27GvbMJWDJRz/CgHLJgnl51cRMJkmne5XUNRYOj0+jE64N
1OS/wTw06MOTHHBGtNm0sAHRfivGxGM6MTLymcmYzRD/mRJ0580dkyoA0DmkLW3w
QHFJdEO7pyciCCRI47OBy4SX3oglMMDYmw/vIw7B+LCdYYt9BtAADIN2P9btos3v
33jSKFt7qXW9fisA6CUXSAfrUhHaEPeoRhIH5ui/FGMdLA9wuPlNiE9RGZfcutrf
wCVYGTNqwqVd0kljuuBOjGNA2dlDxZeyKBNF89nPOIlZrgPWmA3IX9NSVnEHIU1x
dJ/JhSf45pZYVn7ZFfRqEfxqQMQvPdKVHxe4SbDRMwAgAz3YSGuZgZw73e3NoFaC
0PBMw3mVKKevi1JuYE8ZfbLWeOVsnzsRv1mlheu0dUqwuuYC7NVB1emL1uAXNXJ0
IAPvRv0cF4lVtkt2fjy330u6jToGaD2eKbFyRqssOY9aGXk6WFtQHsASwvLjJtxX
0a1XgeYi8dPSCihTc4YpW1e8XanJ6r6+qD+2BCW5fBXv/INjEn4bBgx60BakHpti
GqP4eWTELs1HWFkMT8owOdgTRnPkRgN7hP5nVaYjcT3W5S0BXHiaZa8BdL2JpChv
B3GrRD/vRK8i0MiinTAu7SvYuW8e2iW16JRMuiDCOEIaJVkepRZdA+JnFSTecVfo
KVuazJ7XZEOjMfgZh94Kv8J0eOe52TrGBzJ/yfRibBoxefh4UoulQLPDHwgL4buU
/EEYX8TDLBEWV2mVToe+9RJmTWqz5TF3RPFPQd7Zkw1Y9BOslY2u04q+rFaQi/yH
iDoBmUEr36L2toHbS4dRKwW3+TegrtFjPjT/LTOSvTDRYXkvn4oVGWdYUJFKNlth
tdhIr8i2Clviqtq3O4FZRfNCq2yGukRoNLKe6lHdBY36anf/z1BldWYH77NFRUPI
oGB9Pfwgso4ruP187xrq0zqQN/hMxyDHj4d4FFDlnd9bcDc5vmO+O5Oa0S1ACqEj
3vLRZ3oMa23w3bqiGLSWDvcM9TJDsOMo+lXkP7kD2ZHZzkzpgHo4iJ56L2kPEPsj
zCntlAjOoB+ywVcRNszIs9fQfnBy6BYbUnfo4M7yZiodJcx1nhcMXcnjb0Ls0leD
/9HQqTkTM4sm2rfX/QnCRTStlcsAkNVrHytQiPUbSjzY2TJFVFjoYbU58hXTcecW
i7JRDgzROFQ6v2N45pnaaUF6eziaXuvlnc3WiI8sqVSIPHauMtHxH842niB6b3WN
9rUpcUZzIsrb9njyCwb5N/dhOQwbGMpkA9mvt8CrAWCv4HOyYLOVcVJYP885PzGn
tAtP5SSjGFBBVmrfe1twP0dTOsaOE2OmMWpS6JV4fyGRIgpTwzRwGEXjkhGZH6MZ
NY56Dus/1ln7WGFTHE2j0SQ4lzuK1ZuW1Sx2t26waMr0Bj3gqe5ztWcTP4NiHT4p
5lU/I0h4FDo8NOuENB2yJOPTTdjTMbZtRr+leB7Hs2S+xAX7Jkm/1F7HBcoBz2eT
xAC2UCDlhMdD793LtMh0avrlwNsZiixdcwURqpq6+yhpKAv009PyQKR5k4Bj+ynn
ef7PvCPnBSQZvqxZCHNsltDAWSVfgw27nvkhOcURz0MYsazcvalPN/N/eRwK0Ald
NidumnCltl2tU6YRuWj5UVLi9oOvWz4a6d2IxjRGNCrqKWkQspHYT8TQo+DfZYzW
68QwjhsFFdgKsxPucXPwSD2Sk9KSw+neIIacCwItzPXHlHsAFlLlxQd1032sZ6eZ
lIgDKNCahwsx/1ELDEqsfTh1DPJsAlFeWUhitCkYhpz6TFrnM3Y3OmhF6kd18ALA
O2IzXAleb0TLuWprXMp05fmlET5K9PbU/rgkInah94trBWhSPZqLe/Isgy5hpyRf
M/PmPy/D+fSsORSWdKToT1Eu72tM8ZP+Nu+8vFCGI94kS7c60i0HIGhnaAVE0cLA
+F2IoiiX6LLxvOG/Xd6LxUaQ7l+y4Jy4Ucb/gbsF144gH82d3TarQOxOeH5vn15z
YYqn+aLv0qcG9vmmzL7xDFVIzWLaaYQ8f9VP55WSMG38+qrPMgLNbkV6BmmQdGN/
0WFZBreaAf/M+WKMvQ7FFpJhQCG2BLMPkVXV5dn1/ynyEZo+t6NNLFOPoNvnhEK4
309IyFuC+EcBEen2NUHNNDQHopVRS2Lirf+D0Kcl/kvQvDuXX0FlIXtn3c2Vgtkt
hml9gb+/6pkeCO4ieu6Vp8CbehV/SlcTiwSoAzOBSzFOtt9fuPRI+IGp3U9A6swJ
/df02r6zRHz3rYKH9PnFGKWmMO892zKagPnjZYPioMVIMwj84oALS5W74auIKa+W
ZHynqi0Hz3cKCXc8yd6xIbQEi86V+WcV8hHZjxEl3lALfJ7++0SeKs+ycFbQIo5s
I/rANoa+jeQWjypQHfLt7YfzHZTuhr3DeB0r5hXkHJy6hhOiTYDF49C0eBHeu0Af
L3aO3JYSv6QQISLW2RBEbyjGcUdyhaYU+ZAIcnL0pNbErDImy8NeICtcZFZEKxgX
LwXylRFNaWt3waDcyFgO8ozfgteXMriRlV+IZSe53cABAPz1xZC3h2quF0OMa4o8
C41dSV7DJzc+dgvz+mY/wSKSSIzKXk4OHhFa6527h0MZElX5JU/TvnqUKuJhfLm4
igwig5ktKwERMdkPEPNl2T70LTU5D/Ul3Hm38459IJH9xRR8MbcV7HW2hLhR5F1G
U3pIIjbB2w8D+Ke0b+4zkBTaWGqXE0UgP2N9CkBaXO2TMbYHAuJxVgsLzRoVuZS9
jRbqPpaIvZNL/PCF47PYukh522uph0XzLpy0FxPVEBaPmTm/af1kUHIs45J53xlE
lZX+FFHN2nMwcIlzMEmUvIdr6xdDT+eu+nNzhm7/5EtOxq64enKYEK+NxSsoagKM
BnHniZEMJAraWThwY8B3hGdNi/r5zaNLYfoAUTRevJ/HN9jWlub5nVUCMCSXl58N
HAvcDdvhXugs5M62wmAbcbShQEpWfjKn9jm5XszzlwFgI/GQPN2h3pOwmVvrJT1e
PjwXVCpLOXGNUPain9E5lpNecbsfXaTu6a9h7M0SVKHAAOSz+xmJQSXWcnF5/6hS
NTXodGmVD1BwPDV6xkx1QOOBOaPjPRnln3W1VrpTNzmgLYz1bU+gey+tJz2n1jhS
toIR9YVCDJOb8Pay7QvFuGfW8hTwurXyJ91m1faPz+UI8xtpMPDsDo7tYA1n4ebQ
kDXWIGwK1MHE9635fnz+94IpA5RWEQjVVEUsMB9N8d4p6+IDGWi6Kpie19aUS/46
9HWTmVWcEHbhBLNzMDwWwOrwySRs8B54nWhehAclZtmKdspeR8+m5X8KQkMcFv6q
gsesFKOdjeZhJFqGR/wLh2M5Ux47i/d81P4S5YImxNiPIzFBKEuKyXU3DRj6E0mr
CaEjj6fDWVA+JTifsEbOr5aK7MIcnZy9Ca/MhXJ1ZI4KOVBDsRnCBe5J/+nPWnVj
rTqIIwjmyJ8O6/hRdvZ7Di/KajZN/pFUnfEyTd4/OhQ36mgNBGlN7YS/Oc7pDMau
ObH/XG158CHSoRpo2SSzBGJdFqAYPJSFOUHFCN/XjUrfWvhrHDj/OnMFGHSNBIHt
L/vC4uWN3QojPlMxLFJuI0TDyd32Ej35A5+13F3M+k1wI4QHO+JJdeqVLIgr0VsF
qiskRJqovOWIdyUF1NM/o+2bWahSe5jf8XAIt/A2rvfw0W/qKyjQAH6Ixgo8DMXs
mmtsYtIcA9sj312o6yeeh8ZeuO5pU+msgvZnrvOXqr1LVa1yzQzaLYMGtVwkZSOI
uPlbyd/N5oL01s3G+BZjl3GpOuELtlz8cJsnWdOKhKsLMeVBqu6quj2C7QRVXVos
0hGJazl63ujkaJLbmM8xiPn1jUDcjOwosNNqtwR0fbt6cyVQ4Kf84KdC9OI2foY2
tqWx7vGiVn0ZJo9h7K0n+GHvf5ifOSzAcxI8v/O8/0tZL5v5YWGcFSp5jTZph3p+
/y+P2TRW5zmX0F6yBdDK7PRcBWm7HvF3S+qmf/OEYnFVvG13Q2ticZ75cs5JGECn
S24JLV5RcNXBpAdlw57cU2Zm/eGvHdiFDvjgInjUqWI99IwUTwVBsnjrUKSiUH+j
uSU1ZpPF2nfaP3ZUShIga+pznCAXdFzjbn9ERK5eVvU4c/7dxgVSCOGejQUFF63t
oZ8dH58erm9rQ6E7/yTKM5VjSFNHV3ikU2CVCC4by9HzMf6nxa5+cUKf2TQZmnlB
hQ3Ia8pE1BkMFRMa0oCoG3j/A61MNhZ4FT3iu3A4LnLxPzJlomtBhaAcI2QKyKR+
Cz1Ex1hfJsv2kQ9hMF0N7RyLmL7kB0RESqJKh9YxhuQD7iqr93nTCqiVUmnG5WE6
Su6/Mk/8LNY9gPDPIM6anqF2WODzHx42ZmYHotLt6GugHRImHu2LCzz1glEWAYUf
o3lrL+8dyUUIt0tRViX1nm+t6ZntTZxWuBiE/PNkdyUCkEUO5V2rLnfAgQuCF+HH
i7rQusJgsMvR0MNI1scuXwg4ItOLcSdcZ+wYwtH+/gd4imKLh00bvx+Jmzfw6tXx
8HYrlCoBL6LLcw1Knvz4+VmP/K6E8H6sZwAxX6C+SAg/C99TPi0hNaQmdB2s3lYM
5KQ2cuoWi1QtwLYW8xwHdLvV7wawbpTgemUaIv6PbQ0CkSOWdkkvBMBQELgXWNG7
2IDRZyXDJN9/pKGAlbUOo0Q7fYfq3cp4vV4oRBPlgKkMIW/yKfbQySzIg/umGgV6
LnvC4YPjR3M4WZyO1PUwPmtMKEjKsv0vP9kcQtVRhgqrhej8oqbAINtOOkhLM9Hp
tSM4gW4e/NZZ2PgyIiayHOUfaJd7BfyO3PqbgBNVSSvf/sqGRfA0Y7goVSokR83b
wvH4nqJRVAqayqaxX6D5ePJSZe7QTfeFAQL5b6hKgClsLoR/fVhk7d6WdXAk7j+p
hBo6AWK5R3iOCfKym4R9Xek9KVWeNHBAHrkqb4J4DMFeespLm51TCrKcqWQgwCaN
K1fYpCP9KKuLbO2W5HPNzyTL6gVl/tPDjsP5zjg66FYyeUExV+uFFEo7zWu5gkGk
HE6erwm9EpvC0+6bLl7tuNz32lfOPRKNzg998x6sgMNsRTwgXeqeanSuxAwdXCBV
1cmXtAI7ykVX3haH05KLRD0xtMBR8uq8jSQniWLEu2oIDWMbGgJXlXidh2TTVL9P
p5wGrNKGF3szeNOHThLrF//yleYN+mS689HK7bYI8++ghL89g0djfvhLVpeTWR5M
Tfj2mBBIIeQv1Xs5gKXNTdsKvZacyrH0/C6CdCbmWZ7x9UoE05yoN7qEjUVuvtqB
382TV0h9/htb5wkt9cl0fvqLxV22PjDSfBUONJuRnSEayeZEju6qACDHijL/dNsv
8GJMoqVTgDH8Rmeg+aBXAw7DGqiS+g1o031DgSkqO9B0DAA+ZDfGRr0bNJFWhBA7
lKyzQIHoeuEPHySrFLq5D1A1gjBAxWiEPnH9JoPOrzKdL78jX9r8YMK8XgfJ5XG2
2IGEK961AiicUj5SZdfn/9uTNfSZkn1mOBEBBYaDDCVa73GCgkE+bho7fS++jZve
rmpGkegeYVgiFV5eTu1vESoas7fErRcAjB10H135LIjLWFvzlSPLxTL3/jaMQzER
llKF+Hng0wFxDTm8JevDCLVGAlNv8FxUPjsxumxlTLlspvQJzYstk09lwJZ0c2Zu
mbDhimt1oLE50eTX+uTp3X3vigEtLEO+NTUTHVPeISMtZ2cD2oOkmT9Jx/XSChug
8OCGNEglpa78zbvs57rOeKG6s3sPsqibMDqm+SZIjTqQyxZrazxYuNEJvoErjVVg
FoizgFTohHsnYXgjWRvMYwRfFjCdS9wf3/U7HlYK9yijSZzDCq/KPpbZqAxpkRAB
NV273EAvlqGpTK7gIqtOygEjayBKIv/iJ1tmKkFOgF8SFN4/18N7Jc00JhltvIh/
PgXFC4E64Konbbnl1qAO80KLg0LllISJDjYae/AJQOYTsvWZjFkP2+ysBYH+AjqK
e32wOszlDyAxrHq26etIU46J6YVPGu/nqanQYnpwJx32IRb5z/QVVjKVDdrKxlri
OqBVZQs5g40iubjOvVELR+6v+BSqQ3YGQ6ntJh+K7Hs2KXu/6ArxybYKgu7fnNPB
nQaGGX+lkAlCC4c0OvUhaLrAVNX72/4OWFmiYM/ANK7K/XilSZb088NHyGuNbSu/
qm+QAOa1TBOWcM/VI1gVy573XtuRU2IxSEpgKcAD0eW74kaEggq2wqrjt0CJD+1L
bI60sjsknAuyK3jmU2W5m7fO1Z2TbBG7dIH6uhSNL5Hz/8+uX5HBkLlFbWQ5vbrG
Rj8yU5Aps2IdR2uXoAcsPFJdcxmiQSLqfBWcXjtz7IOfwxTX+9EqqTHTGDNpBP/M
RlJSTAUrxsr4aGImomgqDox8MEEQXXfwjHBcH3amxxyHeulcPtsx3H2XEnJoxd8g
p1HkdbzUBtsC0F4Ga9nB8iuaaH1LT7WbGuImKDJ/RlhXT7xB+Z5bdswlJCzH+ySi
+sVsC2owEkA8Bs8Zqctv5shWycvVxjh49PFBmVIdbKEjft/bjjtXPzKXKhQLhucN
ggwv79T+b7HB+kQvnoinVINJ7ghw1VVPDtu6Wldv8vOCtOGYQDtXi4SYm+hz4Ln3
3qHm4g5nfV7Q5prKIIG6M+B50kIMbT9P0I7vkvx1gzpToncJK+nXH1eGn1xSSJ20
kDfPzWhvKKSc4ZQ6TE4q3NHp6/C+OVxs62TUgda87vY+XmgfpD++fPGUs3fuUY5B
38q3wF5rnL159q0deBmBeCrEZrtxTWGEu9FUb1hBn96LapznT8+Mu7lB7G2l2ZH2
w3PMygViL7c7ovFVYTst+lTXwcgNLugOHplMP24br6BVS/s4Hy2VraszInGMxdJj
rtNqiWJ4SeSWjsVQ2ySXcXJQIMjGMrR0YxJYaSHbe5z5ScMVSA9V9ieFgbGn/79q
02B/hTcdbiwlxhBu5hykYjrilxBwVSydDVXDF7F65j6rOofymJvO34/QsecxXIWj
bDAxW/ltqdgPFuPSUI9J6WzKL3dSyRPwV71Rfx+kB3634NWAE2pFAQQ2WWMEM9qC
paV/Gq/1BAged9TpPmM1cmqUlqwA4UNnN6HamPe+K8/UxMQi5K8W0H7yg1tUK/7t
CgKuOysvmZwmaMf625s64v3VXzp3sb86H8LSMHZMKw7Ni0TfLk4zDjPKigNByd7I
TmXDT5VPNqCUug6YXCu0KrPP96XfsJ4hKMzgFeLiBemFijumslKOqgd7tUZTN5jj
Je9oeDKTtfxlKKMKWIKFc3P4xBsscdE9/dWLgB03LhmrahG3F6ACZeHoNhHwOGun
C1dYOTzIT6k//tzhaYAemP3WtN5r55yNDyaJvFqVs5ASRiCiVfLgXezHFX+rfZ6n
WVwwQYuvkK/4aUKTiVxIsBzTxCClYlkh3vIf0QTnJUXHie11zKmFraBWvD9Ky9KX
drOEeHj5VP2OzQObI2y9iOpaM3lWko6U4wYw6BSZHb6D3E2c8eYJBmwljVxMk4j9
fUJi2cQGCtZompJX0moU2+LLnuwd/ZmCxaD62jOOlHl6agVcmtO24cTPlEZw3MBa
npxbBDWWWhMQuBbHyBTclJWrHdVmZxkZ/5bp7KBeFt+szUexhrjDPA/4vjDMXyUh
Y7xhC4hte2L7BgJfeKRkWvoSWByMopLFppbCSAQJDR6Pd9k/j7/03kRj2h/E1h5/
JeOExbvDJ1HmQQq9pdS5w0qOJcggveol5B3f866kfRcstTm0VjR2nfg7J8QqJK1i
Y3gzDvwcCHtwvObwXnDOhpspGdqXGizeOUL7scYTiHxTWJcukhQLjGIO/7oYcTGa
h0qn8fZ1LZH3kQoY+ThZVJ930+8RzyWA+ywu7ARDNSiZiniQyLlfzcfLGyHRb6Sh
3RQq7OVsfKjYVbId4wsEOBmeN7OKK3u6YixGCmDi+CDMb8mRopMnB2MkbVWlgGYK
fFYrODXMafLLbuqwta9BopqZ2TaBFS84DgY1Pup+SgjxOQVLdoj0RbRW/0TEvB9h
dDeISgkamTx+sYwP2HT6Z5AJUg8gx+QTfWTG17gePSPkxzER+ScI68WX8e7UHKTJ
YT7FteQN8OgUhftnMvhBPwvfvtOEGdQ2t0VwZHupDTbQ/AErFuKCXYKtq3ey67Ez
SmSCQox101jGXxGHp1kmNHl33qLTmfI+4UqhBvnEsvyUVmu15FCyc26GuUe2mmPf
zOIxfLlUzk0edVHuWabw/lnP5zYeJ99REsrK5b36nzxoO+H5/sZql7j1l1HYxXNn
MB1Oed2sowWtAvUvXiDQJUeVXxXgPe9moXiicC3mWBgVLv7UeoCpvTMYQDSxkCYf
rOk3+RO/lwLTnadn7oSnAg3+WrueKjmOFqV4x+xiy7OIYCKk80FeT7ij0eoGAJ4A
pVeB/BHXm+91t80P1UavcZJr/Xpx5TFLWkKmxbZJrUWfyXa2CRNxerYd6Yz6wLNZ
zY+6f6CUwzwtNQJb+XgiR4x1tEN0NZl/HrHuY8ZyI1/w1I3RD6hCHC9JiyJW61r1
YSvfkcAdIDg/+Zqld8kofQJ6dgCjD7noNPMSU8ch5jKQw0nYwz2U/w/n5RrGnji3
oGVFge/G3Vm4donmF6QpwwywbPyXhy97jpnvWpLcvIICisttaTz30n3dMbe3/0cg
uXZNcBm4cvYilKmktOCMDGBqvFL2mrXic5LcgSckKpuGv/YHA9YaP3ccNvh4vwwp
oqi0coMDnq+FowsMRwNTD8CBr1papjyW0I687zXkMAQfh2gWF2RJHfdNXpFc5kJk
gSf1Qc4xa2zrxC61C7729vx77E3sEj+PqmUQH4ah13/1trr5KeVuuX055SObpSDl
ll9SD5i+oUq2iZW6jRst80KKNOZ33j2h/CcNV2BkxnI=
`protect END_PROTECTED
