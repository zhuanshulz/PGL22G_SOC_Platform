`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FeHwlmE23MN182tYVpHuUbnTdu4xA+3xN0yGnjd9esPWoH8c/uwEzW9WTcJChM6p
l9oxEkmd1S85xhDb9pIRHNQLEMbgQHugj1I0jfAYhaannSvdPVyqX6iFILPFScvp
gyBsAIBBKrkXUp8ASFpB25aWQB9BqHxSFwxFPmF570sYB86GdtQN8jhR2wyOEUIx
LTwWxjNrmEfdXXo5SKbpXYtgcim8otvWpHoo5h8fnuTS2lLawTFaLET3bX35kqJY
3/efpr+bvp9WFleZaxOeAYe4bO4P4qAp8OOyZJg6zyvWX7MVW7cQ8grKsjem7I8j
cZ0ZvJZ4LLtxcHDW3ksZNAgNNrMaYx+/fWCcPyOvVH7kg5hf1d2wOQYyCXu8/xSB
Lp+WyhWOPTXp0JdATQiOacJ0ELAUaCL2qaEgYaIi98R1PBuYOXzGHa/ZFeW0xhje
5Dg9wzlfDXNJagEN5nQtYc8IN/HpzP0QOVqAIk7HTvGD86EFe1drlBfsDyYWdfMw
198YXMvz6gvk72r0eUROfwkyxUGAb7n5VlRBKVSi7DI434AfgTd2alxUaS42KY7c
RreHiQzJRMLhdaOP1tSEuoE1HuADqtnE4RNIe97TPtdyerHHwmYjDIJQDpRL2oIS
MpINvIq3tgLD82D2E6vrW2XekfpNdcqDnEw0q20rEU4GJ2rsw4DggMdzbHz1Y2jn
eNVonZLWgggtWrAql43vFcfPHGvFrV2LdEFY28nKwOXOy5erd6kJM7OCN7MQT9DV
Yk7n0CHzJr6EzsO5qBWVp++K/jb18dyIl5FwPRcjX29KXbDzm9gyFAP5Vl8srrfJ
A8QkcOi48wPVV9i+1GWPg/RZ1tT/mRu+0D6DdaYttEJa3eEDgGggtKy3gSQNPkhs
5X3UA0jdr20nsnUmnOtL5BJYB3D5P64c6RdeBaTgDHWnEveFNIbUszYUzu56eevV
kO+BWr4gmXeKoHAvfMu0HhBEp6PeZwtWEXXxr8uG/2tiP379ag5p0dq5R5ZRNwjd
04DrQRb8SZ6c28NA1Mg32RloQyPWqVJ9orDZIsMDZtlyLjTi6W6PIC7YROONquCr
4+3o+mfSxda8fo3PW6WVR8vvfGgaLtNvmaL4i7S9triAcLgsEcUrQh3T5D7TQS3M
IusPfRDqeJ2EwV9CxerB2+jVDyTXQRFCqvThxfB79qctj0VRue7srlXYkiZhRdbl
j2Fl0YIrBxBtlrwDA5VNSZR8DEYjHAnypmxKrkdsCGlZQUJEMNz0CVmaqkvl9t7R
T+ZzOLavhuZiuFf7J9Idnia30n8maafOaeDmarrev0M=
`protect END_PROTECTED
