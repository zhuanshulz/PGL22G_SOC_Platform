`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lAznKSUJFBfVJhFJ5XJ0Pk0BW7BFlk8vEyMBHxgaBHXgLz8OX/r6eVCm9a6ZAudN
K3+WTQ0qpbaYUFOqA8bufafASZJWd4aBSWCYaJTjBbqNf8jAzcipnWuPudl2CRQy
36Wn5a6bIuxgHWMM25e9XMpCItlT2eKVgwATy64+4TBhCfEKpCLN6/jmIcAacdIt
lIQVTIcQgHMkrYueCOochF5yyK6fXxbFLecxNwSeuVyryF4zzyQfzm3ewMIRl9Re
wT0ZG8Rvl7yMdkgQHgwQROY3FuPyEEK93K8+J3V9Cj/qiwZRHzi/fdC/WPY58dQs
oQTwx8LG6B9lG60IQthUPKKtdgGS5of9PBeCzwc08R6uic7ZUybbY8PYDI2FAZNb
Z1lmX4E8SPx0FszcwASs3PCgCTkezFL/azw5d7vytJ5a9DptNyps1lOkdtQBjl6x
Z7qGXkBmYZiLbyIJaIohsRmkhnUEZrzt9YOd5JMrbvIg5DAT9qhaiUQ9aVEigMHU
WSnypqoPZhNYzYw6nYCS7V9ASyz2LGNhn3ZpCt0qmIUpUf5pmocScVmEYwTse5iS
b21AvDGffKsy3XsXu0pHxbcO9lNPBZi++BsQSKEes555H9UqINiq4TtMQhjJ4N/B
CqTG2oOj7J6ESRkOcpZ5tULnj5lJ3gv0n7tcLeQashv64cwKLuUowmLs1MR4dJyt
03i7uXycclTHxp64j0RkOYyQg7Z8BRphA1XEN9Eu6a4MA7MwQ7lm9V5caiITxy/2
YrZRckOfifNVwGQ2iHLjUwPAap4p16VxMMCt3iAunF+TgideEb2IUyIeYwjZJsBF
YjxTVwloxvv+Mw2tWON2i1OunUjaEitO5D665ZGICr7DVQOEpYvfiW0Ad9lKHLFH
A8glFzU/ZbQgmbonrPU3zzLeqdKtnSr4DZD+28CGl8S59neRgowF3jgvV/VPPRq3
PWbqqnoFr44XJL9DNlp0kcLkib9e2MPj/vUohpcSkUs5TW6Uu3ezJH6glyuRYDdY
ZPlVEHSNcEfJ9szdRBgl31j8WQ8p0K0AqeWw9tsh7JMDbfqWbRcBXLhuZTZ0Mhft
Htkw9XeqvO8Znpb3+E1b6gm43x8VkhhzB1a43BrJELw=
`protect END_PROTECTED
