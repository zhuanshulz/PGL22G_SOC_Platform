`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vaPPtjnSTViWxeskMM9s6ZSibtabVH6Gt+B1raHcVKWEuC3mEZ5pSkGywIL9vx3R
MgsUXLfmlx0l2IeFCrL94HQSP6mTIRDXYxxz9HzCOHuhh9a8igQ/v7GGtF53lLUL
399VpP82rfTx7Vb+0j5uDuEH4kMx81lllOMKVqOyBe4EdrW5iF1dfI6jMwKikk6b
D3CoenOQ8q3B+wOKWVljxLtIBySOadGrbTIiX3mc4f1VBINGBQrdMTf7FCB5JQ9b
/s+utCRvkMBAcbWNEYiRuEQiyQhTk6Ec85sRd4oXf6Hp/QhB5iGrQep5+9NopQDp
AyprG26mHO8rq0M+PNwE/hpW6AhhhVEtIW3G+mrpek70+5n0xYBXM0fc7EIqKFvM
7sQVAIDmJhRJS5wV6KPpktXKa62b503kUMBp8A8Wse2t7VQIrFeKwnf8uA5nD6eQ
2VnAUx7nzR0jvE3tBvoV7+je1TduoMiZ470pwH0BQ2m/IGKdaSZRcwbSgGkyOqK3
fJstKhrsiKZFLun6cW7f4fBGp6V49Mkt7m7DvFyHbMl9gU7QmghIBVwo/P/JMJTr
vns5gOF9aXedx0iG5jIRkPudMY7ZWvY3Pb0RbgHEZduOlLTGwTPdKmvxX7GtnB/I
EPBgzheC5ckqm0EIxKUHFI7GslXDY+ykgv7NyyYZmxvhjQHSJraRstQKCoLonpmg
srnY9+ysSLH3lu1wNHR1eGsCIbxp+fE8KqKqb6Ye9xaar/vIH9Rv0t4qwrntENrT
5KKwdOrmj5fuZejcYp2HgLYUsYdELmUxFO+MQyd8La7ogYeNkqrFayXar2M92pPd
g9ceMfirNAbx5ocfxrebX/yL2hYFWp0duebMqWwzV3eC0hb9o3Se1DEmS7bigAw7
TYc0YenOJJ2bBLqLyboi2FBdmECM4YfqSvfAxWbiolKhTTe22BcRqlKFtD14z0pM
5RQL0cz8nnwcCXZvNxg+0x31Mr0UJHoVI0cMn2dsZKtka5I9hBHozMz/tsO6qRsO
YJ3nzHsVaqUW78XKmfXSkg==
`protect END_PROTECTED
