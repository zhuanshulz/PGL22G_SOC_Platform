`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RW1HhuK8+nwGawRk+ST/eP29547Odd5cao2/aOVylZH1Xgl3FcXR9KZ1rZwG2VTu
EfaEsWu0bYUSh+rrMyNtYov1EaamNc2XVJ8imGeosNXmk3JEGJluSo+eCJSXBrza
TdtG8ymd0eVaILwikI1q3yBBTOrDWfueEyKWldHLg+z3yHwJGRXF4knC8yLN0rSO
rAQpB7cPfY8vZb3X7gyfPIMWnq3vVcaqIIm40RTrH6NTBGu2NFF6L9BQfzprR2Dr
b4RryCMratZr7YzU+FApUJUACLmWsVSag77SHhEcBlT/OzaTYdKKjJCqfV3g3fJD
nR9D1gERtF4VWE1fWFLesb0XyzlJba31ldFkbFG+26cL0IU6nOiDmfdiPAJeSy4J
3s1YZuEpLf5O/beHAUPlsGW6TpPnGkgPEzKb4PHAd0QDDnfc58j2PQRt9sK7Yu2U
FvNWTwHvRDVns4kzCzH6gFpl8H6L2lUGg+hzfovrmQtEqEslyt466NekdVxVkFqb
qMVK2U47K2eJ2njE5KMx0TXzFwLIbywQ3bEIn0Pn98YAhpXGg6l04eol5dIchsff
xq7gcYSMbWtNxU/wx/hffeQuoAaxEQhbkAdTdrAzptYRfrNLO3s7mvhGieGdYA3U
`protect END_PROTECTED
