`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dOl+yCtE41V4Ky1XkuVFuLGtifXkR0mav2ULZjhNvSv40qugCREd4y+5/J1I8d+R
Fon01JmJl8l+25AMAS12OTsGZTw4xStjkaqxcaYMB8qb5x7etBcS72EZ7nUS3Fa1
/LfQss0DeryNejwhqvIWMavHNHdtfoYWxyb7mqeQkFNbneKRSitbKzWEsejMs4Gi
FrnSf9M8np/VEXl9/WGR60O87N4ZZAXgIEyHboyBtgwvZLtP+bsjDm17KsOpKTmC
pqo3iDMTDLiUqwqW7P/BXvcZbk2KPeii3RfwP/TaPTHGuW+AJYV8OJfFROJ9Ijbp
kv1YY45zmaQs1IGl52Du8CvidBjcJxAx0w6huUb28O05EkfFzXDkCA8BSi/gTJAy
j+C9NZiCH5Kh2aA0qLu2mZRVs823yDyWSiAwrekc5mfCyDhypCTf+KsHUQp66V9x
o9z1qwfreiV8T7rU3MYlsOWLYClbrBKGxvgyJONOz380+RQcyKDGLuF1wO6n1lq3
/ls3bstC2YpsYyb2N6g2RaAGJ7dk7ySpuNTYOEEdlkGQBMgKkPmD2rvWMVMrWiio
GwqhC1fdg+qU2mcJXJ+6oibFshbnUfUmhd38xso10JICE3tlJpasZsGxmZHCNBz2
MWyFgz2hBC8TUNLvwfjH6rUr/wpKWV53qjar73gdXP2EYeTSMwdkhs1a91IwIcvt
SmPXQElTGgF8sofkr6Pz2XWvKCfBXA5GsaX2yGDPWxJq0IqgHgh8ul+p/52S5Vu3
0pfE2EOGCb9nmybbUUdP5MuFWSeCE6F9B8x4vstotM4mHgMliR9PHZs5kOvQbCYE
3OygvTUnR0rCa7kcW8YlukzuBaGjLlb/jivtP1H5cHpxCdaX+Q8TKbggm3VxBqqD
6sTq/F1TAXSHkqeqSfz5sCdAQKduvlJnq9wur25POkk25aMdr50SZzu6SEBgys/G
7Q41W5p0rSn9ZEnNGWo3fT6mrCTxWeziC8l3sIAIYRz//cE352+0mv2rlgG1zIzU
5L7Em5ixdDlqrYxqDa4tXjygOuTWOFDW61u3U/GN8pvllt0ULhlyFPv9lzxL/4e2
32Wfq665hmiNgEVaE4Rvogo611CZuV/4wAtoXFpe+VhdtFA6gLZzF91KCQRYbCSM
Qiik2cOaNmzM+bTdcbNO4CTptFOWpjoyQn9FybrsKzuQ3+a5ng5TFlHdQXxELId7
iZRL0e64UqiOOUGswagj0omsXn2CdsNhX8qp4F5jnZXIjjWRdWBJfZKQ+0FMA1pt
JmS4Ff/1cYfC3XQgdz44uQK2EeYnIsFkhEfM5DtprsDPa4ag6dG2qxt8rFhnP8Ao
SCR9/hL2DfIfRLpCZ4jG5s6dsfoYW+5tuXPp/4i+ASWX/7YRx2hSI22pM8Y+25QF
/Vx4eO+aiKGLBPFXLHWi1jwQoNHECy41zWTlm1mE5OUDTVQ/3Xm/Xx4awz+mpMyg
tPy3iwAha2gPbLqTMkc70RfWVIBmMxoF50Xv15PPATKosQlLHRNozsSwq+TYn1A9
CDgrzah+gM8/thEEnZsyeC4nhtM8oG4KXmTiEHFKqd7y2HpziNXMo9KMsECsxGgn
T59TtR7I4lYzpv+zIVy3QPekDiiybDJ9axWEvwTorHeBcf+4frb/yc5qpYClrxW8
2KhHF39/vgRQ8VY8gm+e9RR4tRJrnhG7/rsq/0tuuP/bvkCqnB1QvvE2oLLGUBgQ
KGUycEYo67JWVmcfjpuXIyYHETy+egkqK12IRS49jkp092yvrjsW+ZOZjgZnOCO1
Gd2uAgnmHZ6ymaWnNvsHewcsCt3aECDGTR4yFv7UJCXas0ZwRKj5pdEIhoAYzD4q
3O3zAU0PRAjpSTtUeCx8GnNr4TCttwCut2ir5Stl88iV8Jg0ykjXx7IvXp8JFCUm
3AwLL87YtNHeYNZd9QqykljWryuvc6yPzUzZvYrzNnU5wN0dfTW/MTzXZPJlAYXG
acl8T656ICZpBeUJf67XfUgORAVp2Vm/yVT4SsxB41z0kTiw4n7llkOTuLkz5vvT
/OMSWmFBlM+9g5RV0xthNbiXMlDVr88pRVPR7hZU497XXTSzluXYDH7C4tF9H44j
UvUL+9m+0DRthUjBnhRR3/I+l4QIuB92ROJ1AVIYt/Z/+9AMvNaBtn9QkhNh4JOd
49MGZMq1nnv3k9tHvdiPuVQ1CllTIDVzBfDLTrfbmOy47YFvQlusYa+ce84fmD+3
M5QB36PzLd3nbMurcBI8bvkqVAxV3IZlj8O0YqSJe5lJVvghppCwm0029e25SXt9
VOcs1esXHiQGTkaeVgJVI80OqFNXVeN4JJITKGnFGBdoSfVgYxFwdG5c3G39zpu0
aWzUvJ++eTY5oveXFqPe84xqOkt1zhM4xxW0SgJqspoyz8AaAElx4+nEr40wevgg
S36/XZYENCOuSda1VhEb54RioZpcQ2q+vGKT1LfhNjC6/5JmjkhfguHRYQe1OM6c
Kk65cHOkN5RmPJ+pusUBIMqE/QxjgwoIVlqRPdDytcr1UC5z8sFdeaczYzw+LrBQ
yC680T3RtPQE6j6w9LyLmz02OMhHzNBibvD6MF+BMozK7/obQY7x0LGF6nupANL2
98nPPjITrzfi71/H0qn92EZ7ip9tJB2svHQEJrLA6NLFKH2HlM+k0qYkbKPvwLT8
k1WFt2GJVcxr6gKi/Ar+dL7nlBSrOON4G8zeBoGks8v5hqioIuWqjmM/RZZUR+59
2frSQXd1v8y4yKjRCIlVRUhNj07VflMVTjyOwQ9GlyO+i42HJ4cy3tG09b5TDNvx
pxYwSMlmPIOxybnbezbmuhjMYwgOQXSEFQHgpSRHnDKGhp5hDB4ovxYNcSELYb6l
upySKMphcIYCHELpe/QR3Skiq3TjewzeR6cAS8GzCv9s+Ks809MZZdnRmkN20dF9
Zx8ZwIDPFAQZ9s23G8k+LxsHR/vaFWTlIT/Jb+Nzus96vbZgUpzlko77zIu8l1HX
C6hTa2CaaVhboVl3i/wx9wEt3eUc0eYEQpUiz4vXWz9MpFvQOhL/J1FpIMW2zTnQ
I56o43O9EvwxfdYgNA9COdNRGahUe99Jb9JLG840yJUgZAW5L1uwKnsDMWDbSpbJ
fo89iGA0IQ9pUa6WW3KNyfp3tns1t1AkS/BtwYz6DA2YdscQpcGohJ466uEaE1nF
vDHzCO6r/1/7vm9sTOCz32brcv0N45gyDM457J1+HNJUjef5p6Te1H4LFdRXiJRJ
TuVdGlL1hTQE5UVbT0HZ3AWAEhZFy8/GTCVd2wzaoRqg8N7iCd/LaAPMOUmyooPe
396tYvlKvzS3IN2CBqHemWMVcwcDuGfsee5sICtHgGfELtjpVqNV7Rct0qQK2sx2
O5Cll7PTW4PD0yd3s8jlYL7TDlrF4ILU7ha+lYoqKaGq5UW0GK5OaOy5A2v3mrNr
E3hqy+/QF6AUJZijlgGvUd73u33iIA1nW1j8VAhjtGklHQekYgS9kJtbwje2LQPE
W6l3oTklV0d/jWIWXrwl4nJWkDTWhxS/dnv8TbLS/1XulW4vnrJflpcy2dOWVWdz
2m1KkEeQK0AZ90UjHSgPyplO6vZxVrbRZamYAxIJNnFa3d8NvTQuoNbYBKWHINH3
gaCisfg6S/s6LqI/wNcfwdiYPjnrRgII4q4QxMYyYgwd7xPcyn+fraUE4dSWGBNx
h9hbdB3nZKqhiXOZ3S430EfIqtqoXM43c5PCTs8q8UjVKZ0HPFQO1p3BqEtFQa/k
6fZ1OI4RV6HuSQ6i0UvwVrNMpBTOS1NMlY8krB3KKkOhAHsgl/auuElmGwCZvQhX
HvwpvdkILA1X+CLFKapxHPpE2UbEu6qI7SJuvvLiwBvpPNuR5MLU1YlTUglxHfHk
v3Xo7K8gblNxbRJs9OjvwlRcTC82IdBqLJzZeMuy4kHnOMS7dhxvf5+Rpf3hfuRx
6wVct+4al19fKuzWgKtUO42TnP84hp1w5xDW1qSkLZD1s0vqoaJYmPdJ6yMUNtai
wedqaSUZ1SQ9FFQuQ26dR/0TQEcThXpjrgn1urvMfAlWGfhY6ZDXeDPOVQrdP8oy
xjk/1SGNwI9WA2ia8F4EImoSHvabjHewrJHsbKOL0b7/aW6yeqbowu0l5GkxnaAT
4JoxaCltBsB3u4obtBsFln20wQb/APAG3RXSMdSABjIBDqvteIWTF3JN8yUKT3Q+
YeIFWayZj943M8BfQXASrZAuM6baJkUZkSfWkMlxPMKMlLQCsiplwQCk+o4MMSsL
a9QGnym6E1vJasDDPvUiMEFSQaIKaFrIDapotgcg4+E5hnATcNeOH6RhlyxogyJy
Af/lrBg/7/Tl2SUGJ2lEjNvmSsXneoA+ANWZ5P/odOaPlVbJCL0+tfcHI36OSKwy
6IYXasndlvbFfytJuAjfhfkyTJF4Tg/CDcZYHPDdj/egyZ80whChuIhPq/SMVe1u
q7BiA0I7vqRnD+mi8LIQj264PJ70N/5/Y6S6vLFLlrRtY8ODNlJxTNILfZ3iHK5T
AQu3ScOKfuUUyQ3sJ/tMDQ==
`protect END_PROTECTED
