`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xtomc65PGTKvy6MRcX21aBLDxmYW1YmhowLrGokyqihFAhyk2HGpydPxOe9TrYHz
flto7B304jV51rmoidewsFXlEDxUskUbSQlK7lzYm3zOG8frc2g5C9xxt5meh/6P
ai39Z2a7g1mc+hGFzVSwhmSRbzqcolMM41Z3o7vo56BqPsQp32bfG7hjBU2ITXsY
aDyK6UHZyeuOgpK1p9+PvKL+/aaW/D622MoaBb6drqjhyeD+If+jDoe5N8tDRzQE
nQxEY4Lygm2VQaM+YG7kg72/m+X+sQfeIuojF+nwlw8WRkwTLLTGuSyWDf67oxJ7
SBeF+i/OnZA30AH6gLEklGCOjyvEj2dUzQRpu4ddC8uw/alM9FSK5pt9cgDNI4zJ
nocpjdyUy/WKZlv+3TTrHuKyyRvCEkAZ4SSrmpGzFsKIPE+CRt9uPo005PP6gRC3
YSB0VdmU5fkkxK39SKJ9xo+/uU8f1KYp44qNDVM9Tmkwvp0JGxT3Ae1+HQWMWmdr
eLFqE9YzMhnqQk7CkWqetQm1oAHO395KI7GRbU/UYwRURytFcws+cq8RKJViuDta
y0W8lkNi7ph2GlfcfkpEn6kFiHbIB7oow4iuuW5DppiZiVawsEYuKdIo/9d0T8ma
CcanmRZKS1gUhOIVVNNcvlYs85IZy3iNh7nLFJo3c/vWFECrx9EX8n1P9FwkkcCZ
XJp2WKo3fI4ii/z9J0K1G0n7pEhWjr8PKQZ3FGSaNmxjhuK4BRM5xsdrqbfPLcaG
OUVX4GurAOe+5gxeDbMKfzzW9gHQW3yrqCrjmD90ivYplDHI49pRnceCh1TP/GQD
7bqdbKqKQ3P5xPaHcUOdFEnOh+1Z104pschqRL5ZS+h555HyMbhe2qeAaSRG03+b
`protect END_PROTECTED
