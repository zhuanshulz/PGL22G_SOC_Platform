`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kheljQ/pX0SQh26BVxSpRliBGqgsET7H4+2c3KhSO5d9qjjfa4DooXLBUEqodoXQ
cq/HBwL6bV9tqzAOeTv4vyydR98gTIMMeGRtCeID5tITa9pxTJD4nRZmcFvdDAKm
BtqSuAlPr1+2MFD7WsFF5ypo3ggIagdDOt1SOwT7o76slUljvGvDn7hotN8ZbSy8
yBSqbTrnywjOt9brC3KBJA4VM6cdCsdPvnR9lTD58Q+y9ooscqjEty2D78n67W1Y
7J/C0NaoTbKsjycso3GUsL+L8un3UW5TELF7O8i48pE7+xY6h+nMYWsmNxZiewB5
7kr83AlUsmoUK2Fh2fDMbe6UcgaedjrpaftbAY8Z9jqGUGaTuIHLiVcNI7FK8aC/
n5ZkRkCWnK6437xIOmxpIPQ9pbk9gSxFKpLvoJFDULzKWojnAUgWI1qvN/QMDkx8
C2ry8lARPvSFcbohj68Jj4xxhHYxljtHjX/ozxenEYYpDYTBjOzL/oQzfvdffazk
5BiNsweetHBfmI3fpsyqvA==
`protect END_PROTECTED
