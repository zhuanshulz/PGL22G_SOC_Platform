`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3iIr30WUrXaUXU3ImNyez7PJdjCHQAy+i6Vff0UufIz09rhe6+9CX7f90ABcEguU
zMVW9pL5SP0lPkc/ITmO+7GpPSCwAdQ1ODgYMZrnYUc7SIzcVV3yLUcfGyBKyX8J
QjBWEjFqMZ3KUI/CLnRAg9MTnkBg3XaN6KpiMbGAbafHncqiJ/lKGa5RaZpW/x3Z
g3uD7IUBKrrEKLWxjLicmYxNRnq2SW1U9ZvxWc1BYQo1/VrvZ2MCLQl7zS3mFx10
SGrtoHYbiqPXDaHwsfbD9fLVWylYWlMsgVxfd0XW8tvnZ8sMrbNk7w2gkDEJGLws
EFAbPJ7Zq9fD34ngNPD1Myco8gAZceA7yqX+uQ+VAutCvksHvtjxew9xwA41qGvJ
Y0JVGg9MucXkSXLjsrMHvzLDBt1naVQxtF2EWqptyoxNY6nHiVZX7eezM4QQRG4F
POLfFYnSp3V0ta/pJGp9JmYrXgv73MtwTYRDBCw76r8ViHBSLzYomARVWRLUZ+mn
nmz40KES6xk1kZfY6GyYJPMhqGzcyYGXKH6Z8/QdImY++WjWu/qicBdoqtu28KDU
vvgc7pbMDbIRcK7lUyQ1N9VKtmFpM+YOat3yVe9M8YtE9QSyOpwe2L1YpKw2TFcF
sOxcxOl6yTrUVKxoQyHoFSwR/ikrb3SWSR5w1qSwxE0qHFhdkqLyQ9BOqJVQ4hKn
bT8eC500w8rqd2agS86aB5rbpMk1B9rP5Zyx4vLuKLmmy2e4bvBA6ZRHC7c7towr
BXEb+6GTMCxOgKhzdr9tBY2AMwBWaAXl2fy0cPV+fSLtxnEvJdMwuWTtvg57aSk7
gT88Cqei8PZK3MAmTiLfW+SFB2KvdUQjdvcTzwt7+fDrmORJ0GsZl/YWcOE7IIeg
YFCgrIx2LKeUvDuoRnwkXrhFiyinK70oVFEZHh76fKprkIZuQy+bFIBt1Jo9PPT4
KnEs2ilrVp5kAGzoDOtOuT+984bDXmyr1zhaA587HKkRT7E4FF4kV9qPkjgNinSZ
Kg+AGsM6bmhTbbby7RWWOqBXNeQBoOiG1zJ/wV/ILFTnszc3e6mGZPhI7qDxnpru
9Dmv+35MPLeddfR/DbGsgZMEv6O4Jyi84koJ12BiLBq/5xjV7JAxPirRpkIL1SLv
QkdQmoqV/Ewm+HIr42Y7QLtUklWswdq4l0vOX/cj0uS8yd5DrMoanO4bZZ2FCfmb
iFH4MPrR1BQUA/6ujx8KLFRQsXWiizp3HDpBLxv1eSLgJtYZq1cCjB24RA8zlqdB
H19Ugy/xmOawG6yUlfGw+Kg4xZb/9zv79VmOOC9ltlrgI6SBzyF/7JcEWztHR7EX
sgv7eNJis6lmJbkaw7kfpZuHDpa0+R1Lal8StSJdD9FZRbmCGT3WBDSWTG32/sO+
ZajXRXw1hwgceXS72HTClwJeYVYTEEQ3+ScXYTihUNZ43WJQew+i5t76Vgx3EZaM
byJT4c3y8782KGrgjTQICYgSLtRHlrW1lm7B9MnOQg1p7Ev74Mw5JJnAbLJw+xTn
p5jTq63nsp9Khdl/8nj8ik8o3uAJed6lKA74jPQyh2CDa8/xcWRKDt8pv9ArhBMa
PfyEfiLRaXPuvIdG+ixn4UuZEPv/A2szuV6TFI0yA9WG+SCN7EY6OqKWBIQVkqwG
fxASHXPj1qeSsI1klTBkWe10Jso09NLNb3fIuvsaOOKMSrfOBJSjjqanA4rdluS8
iHCLp4XYsBxO4U042HW8LxOMEY/T11Bu5rNcsK1DdCQTAzHytlWJ323rBilyrBWL
7LU50TkZXEXXrUMUHiykELhSknS6TwvKz/pzvimr3zgdXqaingmj4hy+Gin6EVFG
gmSopiAAuijfabtGykQZ67SXRqPpNQxwT0/ylw6pMhHBvCVTx7FsrjQKchWV+TWd
NQp6xXzcjCuTRUKgLAU102Xc0yzJDIlLgP7bHYh2WT17K8PFG4IvxKdZadJPgCKD
I3Xy4mwutiexc9zj1lNYPVrUEWiSq4MxBlgRyk6dKJILesnnfy1X5g8WkSOEmNzH
p3743smo3S46oY+vxXDCFwKfGvLXno3hH7h0EEt2OBgkpPcCiC8UoA6G8rWXbHcA
WoYWdbbvJk8pZAleeZ8qD1G+cMa+Jg8dRHu1knejaDCtms401bXX7PyjT23+x4zF
VJVzT8nKgQ8eVirViIx2usteWvSZB3qoUBT7aD13TCYm4wkK6AW9Udd/WyxE4CTV
jvAcCfu+eHj0WU9bOamLHzJOdJWA2b5kP6eHD+tTLHoYl1pxMIU0bA7dG8F4RGXm
Aae6doIUOZ3/Cf2I0iQTEDdFMs9B/ec6FRFaNQj141aVWz35QFzKJC/Cu1cd3e9i
VJ0RfIz1eBLBo5Au7MgNpA2kf7WRDMHm5Y9NSPZ//M5sz8NoxuyNIMtG9yZD9dLD
jOpuOW9hfpW0B4RyjULFB8KK5Fm6k/V9EyMBNpAuEseHlcKIC8wdjbzjjWD+E0c/
Jo1+yQjZRY2lBNz+DEgklVHRPNnrCXqfT+mH/ZRG0SVigcdZU0ArPUNps0MpugEg
/NcXLbvef4vKYyZGsR4qocvXF+dy6behvDW2tevTze7pHWwBwZxD1xsJnHUq1y5p
lrH1dvyy8JCO8ubZhqvmjlSEZjXT7JLAHDX/UiVnU/fZBOxW6FcdbsPQvDLjdLR0
V8eH58q/2Bwj7FJl9q0ndc+asf+0SIs2W4P7et9CGYaTbDHzzvKbBgSpQZ/EsmZ+
gJnl/+SyxvHQEXNRbuuFaYhdS2JHAC9xvqctydZeMIgnRQ4AMrmAJMSeSBdXkcoU
nOY1gwspYVHfO3axACu6dZK3zQUyIlrqc1Rnl5dIiDliMO6Wav/TLQdySd98TY1d
XToaYJzYCl2FPsTgUpbijpgODXkF9L2QBtvi7BgIDHUvSHL2jkoQqg6SVXvKd4s4
xSB5HK3g+EXwWdJsWfOH70O2eL/yx7viBsdBl0lNDaT+suYevywkpwGH64iyFBm+
vXJ9Iiy5+nC42pKbiWtk/WqYUboyD24KShiJ1GvRAQH7K49rAX0HprTJR1ExmbBP
0dURAmRMSNKsqIvBDRwPkIsS5ZpVPH3X28ScSu4sQ52Hg28E1nuKfS8fUfntRDN8
gzf33b2Y6z5GAJr1eNXoTVhF4EZiDqrFA/yluYGBMEqxRIvz2W7W7u9p37Rz/RUL
0fbfsaQNSpOKdqhoFZV/rH0xPy9S3xgYTF+/NlaACIM6xIqmSPbUuVhmI+6ZddDo
Khz5JyB4mQBFY12tCE6EaahrLec9mWHxBhKyKDU4Wyqn7oKQXzg2pQqAXNPv0BRK
yF11QLmnFBrOFqNPt7EF3V2hrS+yxtf5HdeNKPg+nW81HHAl18vJPkXD29aEtcof
57S77W7j7VsDgzH3c9niLczQYiIobbMIVwUag0rOWDF2czvZ4bdsMOY2hgyeqf5k
EwqZCUukFFotWyl01++pOL/Syy0WJtWsYrcbLNKkDTjOP/N1vKTe0Ll4weWOLKZE
E0EwiXn+tTbBHm+Hqr/urVaqI+CJ9hvZHjvQZNFK3Ivi5mwS+UGa9mot/el5G9sE
0HtO485YACAxWx+hfg3DMMM+iuQ4aN9Q7lf5o8i9oo//bZKPH1t7cEA3n+iaESRe
sKyxRknSrySUOL6ZalqJDcERelvH19ioOTLaUjuGBTlA4GmvDaJTwhC+KfeqHnBy
Kr2Rc3+Od4/rPoU9AxlYpFEYNWerF3LvOIUFHuG9vq/sX6mqpBAOoNByPGc0gEEp
vMuCqIgtBcU3hebywqlORIVVN+qQULL/1CtO1+neMNu9pvd/oVw0yR+daih7vhHp
omQxQiFw2mHlemJX32vv5M8RnkdbqEIryhLOMJUDgDfd0njt52MfoLin1RACfP7q
QDg5QRjtM0yM/VbQU/LR0hlD/eznFNwTmA7XO7Ce/ANpiEwjP0H4pLlB9rHBeG/t
AmW5uyDrVymFA564gAPL4rLdPI2hd1kj04H/qFUOLDdRb7MfFz7jMTQEN39AVuZz
Ywaf0VJ23a52m9A13JMKLAIvxCVvFsywqqesbgUnJQpiQtY6r2ji8n9SysaweIP+
v0L+rFzOYHWlzaepC/IyBT8yRJElDxsX5jYrSvyR1xZeFtlD0qy9TwHou6GPCMWK
hT6o98NHFj/ZpVqEwIWfTXMV8JxQZ+fTB9k/gacaoMQnhBe/yTdkImjtpva5M1q6
kKpj4IdOrnt8x/8/qAZvulbk6wUwXvDPkGM7evjW3v6wh7+i/uvE/mtaYEsUoSLu
tI9GCwmPa3JgSbaPIzLdAWhy+7f0C6BtfE1UXN6cDySz6cxjJpMUbDc577w4Poiu
hHWNF8I4bkZH5BrENIOCt4/uKf500CTX+zMHmlRUSxDk5kzLFfiBzW/ije3odTo5
TvMZXxVYSORJSfAAlUMqwihYsjGap41InYzYuaVjyb4rU/SyDCnsu9r/oryZW8pJ
JhiZJnJPcOFN8ONZ+5kPdue0In3cLlyP0SDsrwQuyMccnpvcma6dXFoaVQxidqsT
ptvvo+DNMJt4gFqdhJCUqFwPb6EZU58Wq3qsdfpCkisdRu5s9xktFEg70c379VCa
wpTM06cRlJfNp3qRBFW6bhwLvIDbffYQEXgo6X3xBGOl0eAVhVdi8SjRS21eMH7g
/nPYx9NiVphGZwQyLcJZGD9Qsd60+rdhlwnuv+hldUoQDOnZjlvGToyUU6pwdAsF
PdJud2ZDAEwPZfX/xFIPqbrtEDwplk9LfArSdvmAwmNBohU042I1aIS3MGSjhOPv
iaMXW1F6FRk7Q8v53Hm8DH5hjuFyDXFhUiZ1A+RpCelulaMEiBvoW1b3gkTa3n3G
gvOmFMzE3RLXsas6L1XmpaPcT/9MEasA+MDQWyJ+8K3SV6K3R5RMu0rBkfcn7Vc5
Kh8uq2s6BwEL6yYZr+cQBXrbzvny2qKSud1hi9292IS8zSFZ6vS6NtjUGAHz7rvB
0tG52dMR/cIoqmlQeeNyAIQ4Q/Ybzs7zC84YkS6CUzUBzGsH8jeunKkoAvG6IFdh
dWYj9ir0s5H7SKmf0dMbUVD52WzdwDa60O5a92BqxhqitNf6ioJPmzkLi8WMRE22
lzzVR6qgsWYp+jLKhAW4cbDnsXlXIPEhq27rzXjICCZ/j/MHg8qu0peTTEx27ytw
N18bDa0vbSpfH9xU+BdwPxVJqvmLtPUZAFDUgN8IUYa6nN89fxViFRX6kdSQGHoG
k0JOl24XRgxm9VhCIy3dtTdh5qxMchVIBS0yZDIJYTRFKHWy9d1xIRSYimJRY1Z9
zyyir9tFyIWswuf0C0HUXsl4YMldXe6BugVmGJ/2QkaSJt1NYAM36QJ/9XfrHJno
O/fefktp+/kYi9ACsCWZ2BDYziqaPpmvwYCWgcxbT8R2X7FcCWPLA5qwqRqx9K13
HAfOBbHDWFGcwa/moVYXKYWRaSFn9qkhCEgHS1xLpC3y8/x8j5uLYm3mr/PwenCt
oLRywKFSpCUbC/4Op7rjX9Lmggleh/Ejo0HVR0qQwiX9yR+jQVyTJbdUV+dMpbVB
hDY39tpIooJkhjGsDZ8MR0COkH+9OyeyJ5GZz6p7zP3B82VAhvspSAgSXwf5rKA8
sHPrRFL5spOwkoHEu9ya4cNhOPHgMM1x0wa8v5afuRONAL+e3MTrEkQiXC/FU5Kg
rAz7/h4cOSinW9ONdkyKmqw/aim1JBqq3avmQXeSCYw755uFEJ+FnNIgf6wx7hds
3F8fb0HabMKVgk8noI4KwbpYEThJHL3VMLyeIAqwG+XJ/GoC4mhnpj+i6sr6lyEh
BXakwJfeEIaF8QEixyVXpUiNMEPTScXQy1P443/QXhkFh4MymRVaG7d5Jk0E5qTu
bEjizaiAL8Y4NS2MkGTe/WdD0S6cTCTYgWctaunZ018jk2SvN99AyIUctbk3byxW
Y+Jl4oF9R05pT2/0C4n3KkfemqKqajeANlTcH2nyUUx8sJeejS6xbRpdavPMnJpb
HvQL0E5WI6AEjVSPD2UFwyZkBD/2l461NgKCjaIQOvJIrHNqinyiGghDkVslQfT4
ZsWONJPkw0EvITn6Agf/B+AGfwvbZPcVfibJ0TyyqXpjBbdn5zyWQnvwShZsCqri
flewnZ5fF7uHbldnLLO8ZrX4SGa3eJLMBYYVcUsgNw9d33ZohkqJfDrnXqpY/Dz+
BPK4yzhOUWAHOgv6CfJxezKe2x9eA3/mR/F/gxRFmRIqsc37tVAkT52n35518KiY
uL4/YbZwVkoGEIavRUE0KK70o8wRZoYVAUH08Gp3rv2URSHyEo/V9uoFBb4rtNe8
i/h377U7nbr4FdqRSx2uC/s96mwDdLyLTaNn0TqbwjsRjK+9Ft66OBi+m3q9KiP7
KLBndH72uPqYUJx6vgN85bM7F8zxrOsGz350s7LghTyU8F4B+iqlD4RrSA2yl+sN
UU3+O63GjKZbdGeMhvlhNcN0Ph0tR1LWIAxBbBC1KY9XOa/VITI7EXec8p1Yrn7w
Qp75frSTkiLXtunfsgqpaWLKyZmO2HbkgQFv27QAFpTVKBzPt1zf3Q+YBS1PWIqo
bSAbOjJkEPyy/hdRW2/7c9/KpMqtLmDUnQETwkGanYJ8Tkdd/uZahoqBpstoptk9
zEIDijchzuM4WJB3j1IygNN9fhYG2ytpVM/vgi3lPIPHL3s9QJZA5jlz/EeFMBok
MNOyAAxgRhJFMOCM+haH8heQG/obYXeU6m6BEEuOeQ9zbUJrl1oo1KlqOLgioYqg
bau62gLYVcxJ+zwOpzCeyB4+/PdDK7QPdtsWZ/29EbepwdV5P4ENyKf/vV/3NWWA
TXuzEt+V+HJgJunVlXnU3VCnm6yqIGmivdRVKwYRFsG9w0F2VlsTIca/V+9bfBIi
rsTCNzj78Y223PPYLhrv0xbGqQ9BEqVeUk+UleeLiXa/mxngtuGPrMY5pmHrASr1
Yp/stZ19f1lMnNsM0OJGi2oIeN06J24TAq/PkdWgYrZV1/gmJMvSBRZoUdEGsR4z
bb9V/e7TYXOB07JF22ff9PEo9SigzUuWkqrBG7fxBKE232F9QuQDY3Fh1jRGbSLe
sB2Kx365GPBbPv7iQ4KJPlIgAfL+tRoJ9hCC08ank7JlTF3ZX1Y5gZ3kmqQGVcGs
ledH5POdwnSI7ZTEXe59FtL8mPYGweBN6s4BMVWi9AGPhmxhIi46fIWDpgCQbRt6
pVixCElBKAlPW6xlB+tojp0JqNXHMt/re5YE9JJVHfnmaXufsXE8z+dXh8mqo9wv
Z1OeQiQ7Yb9916xlAIkCD8fN8azw7la0MJTs1o2Cu/1QPXskO0fLXhz4mbbgNWLD
ZpkBjAeK6FevJhLTc+E3eYdUgd1jUVN5b2HS504fWSgKDkZQPi4iCtJ0171chWTY
PZo/uup1TYXdEKFwPAWppnIXsfzXLZnIWrq2jh9mJZqoF2wNx49Fev6s5oekR/h3
NLLxHjDHQLbQ96IMdysdvPyr7U1u6ZAaPJ5aldXVy4nVG6kTMZOsNQ9nIytSvLlI
7y/VPF1r2KfdQi5Kw2jO0lBH206BhBZf4+9UbTLnBDq0lKHpvZua1/czoRKGmqZ6
Dz55RFMlwjcWYheYO6Q78M0S/HFQgavV5UwHkKViWs4=
`protect END_PROTECTED
