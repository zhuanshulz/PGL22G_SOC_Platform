`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FuXmSTW6WUaLrp87sX9Eu5FFf2oSYJrFOWb4iqCln3TQRXKF5Ul2Yk6dOn1XLH0W
yvsiwBTXLkninRE4iOgmn5FPfFN5HrXtAgs215MtS9qm38D/qGqtg9wGYDvgbd6w
xUa95q+810Ppxv78xlCixMtfZQCYtWcN1+Njqkobc48LGj1MHFTmTbOUjTfbXZfg
StIUeadw+AzemufTkGGxGHOvget3PBHU+1ekrqkxGWUTpO8135FDalyx4xwQTF9L
8eR2Eld1XxWUyeAeERjPv34kuePGCi5Q4+5BUZMuuhI1S12MYDA1nzmDnJV4m9kZ
lfApCbWo/Eb8yMi/DyPKoBqSVk5YMVOGEGBDH8wPk5uncNPWpEgIUxfOQyUCYzVM
5FDqkXmtJf8vMQlVWbV/tiXx51j9vtOBRSfYneAYgc4W0FCroLdUEeg5TwEo6hMw
QF3oheDdNhqrCgwtPAd23qt5DB5QGL18pPAd71ohdDFjiCjdVYfzrUJklWehydAB
v0dTJiGzGXTz6S25iMzvY9jsJ0cEfXyeGRckNhT1xhLks3Z7mYLDY7SSZFUGRqD1
XWsY7ok3Dzpl5LH34WwUtukO3lYpDIgTLD0xole6sXSZ0ogcjAoiLwO4ntnjp+pO
C2dOL2nlb44agKNcdDrOiqVGWTsDBtgBP0NgsAExKgQsJ9LU/GEXuF3NNIadrdIw
MVG0hCoTAa7NBOQYCtgRC3KgAk4dcK5PEgzHS/UDCzqIs3saRaWaDtfzs2YGHlaZ
P9my/AwhXrEVEsEG5048vMaPfuxTI0+rq/ZolnWTaqk563/FILqTlPqgZeRDz8vr
HzGlcXviwWU1Ai78QjbGEDPh0hVIPBBqUVshYkWBUSUXRtsurOn3BuS7UX6UPKV+
TqWkFgQo1muNEVMvNhkxiut+OxMVbVu1OolazACE9pvZ0yaRa6pUeoTCHgODSO3h
sfZoY2Q1GjOJ1iTQwZ7i1iu2Co+MzrDNTrL3DrqXU884q9nGPD7gDA7bcXZHj7TQ
2TRdxJXsor04Jd9IpwJruR7NZa3KiPsa/Ab3aCGYZc5itQQieHkQ0gUC3zFcjrrO
7za7IHZSFzP7JUwp++bsOHE2lAiLtQpcOmQ5MBcm5sy7qfbyVra4np2GQ8nL+rIs
kq+r+e8L8RnLTzRmApVlYVrY+NmYlQFvwPif6co/9JCniLKgEQKURfdGHkTFIy7r
hxsHW1osTSLC6PuBIrSgCeC9VP46ncZuIQxz+JRIOogVvI/7ZrzacT09x/TZUKZA
/9bxqNBx3WZQMnjFOqdxrkbQMS62EAe72Y9WBN21QfrD/M34pNaJGgrDanfauiSO
hVhwtCi64KZhM8EkxEGgajHxOvNTshwv+03EZAH7Ix1eW9oodMFH9jRA8H+8X3BM
J4bynY+Vs+l5pcOVW4FdIN33lek9h0ZSKaiW4Vyjvfp00srEOpstYVJfMpgEDECT
Lb+5658oOHxoSZA63K4Yiv2RKlOHuB3ZyC6IZtJKi+1Q12c1iTwC85DkRX38efVP
FHEtRO0m7RoVUfv+diJNU9p+ftt7STWgh6eYFh5hXUwDIw69oPcc5CfkJ7uHiy4H
YHtOiBWubb8rq/UQvtIoa5Uh9S4BWXiz/DgCuvATOifIJJl9116z+iA3qA0yEmMd
Z4k84mIS6JncFIiv+WkapbsohdKUMhG/KmO/5XTlo+0BOUtWHlEf20iMo2LTkwgG
7kzhW/bRuzVJPobpVfNH0MuebgV0SU5FXSjff8E/7j1Jv1W/nbZd2YpB6Fdng16p
Ywg5KX2eWLMM6OPO4giwUsWbmtj+BndNM8gINasXAwkIUZOuadoL5xfAEhpRdOuL
vgEUykqxFXSF/3oVmtrdKdDqkZIm1CcohsxwsHY+My+HCHOMFE3w8yUboTQCQbKs
EMEeSqHaX+ZpVQfJ2TTUDzurzn5S2WTNZ3Y1TPo6BcyJcnnKvrFM3J86NX9Vklt3
LkVWyruKzPNSfgOo+mBgbHTYyenqQDEgk3k/KIRyu/pyOSr7VvQVCqCPqCzD4nXG
/n0IftHykdyd70iMqvQis+5QIoViaPJKz85iN594GoNsmV1YPRKtF5uitV1OzvXp
Hgca7ajoJj6eIlFxblynODoSx7kXzz3g4GZ10Fgv9tiwSBWvgv6itH13qTbD6GV6
hmlFCHnyAxCpQlJdyhHF2Cc3m/W3nbAl3+o3DJ5dLUkRjHXk+K4jJib57hwDngKR
AweMJQCS1ULbl29sdzLBjYo8f6q3/EtDUfRGKV7iGfedlHbpdTaLkxqmt9pHf1Vq
M9UNgffGGphZkJ/wP2V1rGeCMob1630iyANFPoGZwbH7+FWTKC2lWVY6c9TqnvBo
sO8ME5AGoxLeFuUvAkKnf+c4QZb79evboNl1Rzaup+jotFwDRtgiAVOJGowzwNQC
Ag5UYzTgyFqxT8dS7nTq5DuN1AvlMXFf9/ek0aeQQXSfq2oteZcbIW3i2sSsM8Cb
E+9LIl5nPHB03gq9HKj28KBn58q1+Pi3+0ihBLUgFVUyF3JyOjGGTNXEBi/FmS9M
bROu6EVcZx1CKkSCwUuXbZd/xtkrHISBZUzJdicOKj0Z05yTyT6C8v4+21i34GBL
c+dMla6r4OjM6NUw/ahtgLMqBLB/aKyThyBWlYH9O7kROSKlzdP/Ivjwg3OEe/sD
O5KdXt17f7li6ncBvqHxCCr5CrGPyigoFzzo4uEyoTDiqmUH+fJSZUQBVf7WCJG0
d6pjNoUHu0V2Dm8yibso+A2LDEpRFdDCkvmlfq3V+zFrEUZuGyhuUU3X3gO0GLLh
new6ACFnyyyH6A3SC8SyOASqWtN4PjzNXlfqgdOO6eu/2kea+SPx0+UHSvh77Ejy
ePxowkFccv6GmSU+37JOKSfWKizrRBAWHDCeV/x1GLfySak/8AtNjK//AC+y4Ufm
VZZ/YDz1bCUL/ba+EYJUV8y6hwQeNT2cCiU4p09gWrwZi6qMl9mhlPLRpZpvGy6n
nDSAcyjQrucAI0iTU/E0okbbgJAnei2GaLtmfgDe7HL0kMTGGnViDq9RyoY0QrSi
+B+vNDjxWFP6iTwXTI7XMA80x6Cy4vP19SkShp0jvJHBGl4O01DKtOzfxso4A6De
jiFzdIbUdwjL+vq6KgqZZFMNZRjnXPHtGrY/bU3En/4zuVZRQd6Eop/6euWJ3+ZH
HIrNELlmZ7xXAYUGFN22Il4avuiY2n0NCEK+ygYLMSkF6MI9w9dyRQPHnXMI2YBb
DW11SYrXXFyfGjj5/h+U1pTWAhRYbG3XQYB2/zpLsm2UEij7L0+DRGNEd7qILPNq
H57joNdHYPYS8mHA7ezPwoTtRIrruOCIEhbXcW9hbPnNM6+eqRox1HZ+uW0uVWF2
dNSsztX6OxSQv8Q/K0Q7S+J8Qvl0mTcLsmE81aeqZ5YIy4v+Pkumqj32vAvNa0Lp
JM+LWNudEIjgmYzbflsRymx1amfXSjvPNBbWs6p0EGBmVysgeFpuErqlSMPKVR9f
2uMYR/5jAYz3ECUAchkhYW/SU/6eyg8t3IiPbD9YVowYg+upcrAGZJiVLSU+FufD
znnwuS0/UnPEykWwTlLm4T6mTvi0Eht4MYUw3BxxxX42WqnVpd6OfsoMbge1UL+r
dzsMFuV6Umm98e+9ZmBFGk86a4TMsQgPZ5B8gMq42/x5sUKtTSbAHtirq6j6vnzx
XddCZqrgEyBURePyHLUrdFk34XOVLWbx5ImYQze9gMiYRdgfFxH8DvPsujnfy+Zs
nyaYqwctVBNo+j0UMpW3S3vwkUF8jrwYTHnzeWqQuusYtPR/TUp/yEIuoHxFpwi6
rxxMDD5qQGCi49VjQW0q4zxM3/kdJStr4J/yO57IgIoBq94NYR33OQCnG6BScCpx
BtL6pF4lU++svl97lshBciN+8fT8mU/SfNfNrTwAVnq9LtKGm6wH54EBMsROSdQH
6SP+ue9+mAzOA9OQWovkAwKqiz1WRpIQNkBpAeKCIRdNVz8sK8HYa9M+qGv3HKDo
dzk64hTKRUfpUC2MzRsIHPdt/zOXoGAxJIXiE326rfuKDqZ+Bt+F9/uNekteCq2v
G/fNnf+9mC7mgiZyEZcSl4gMO9bUKXS8R/ShaXs4cwBXHVV8seagPHD1eqDgoTCg
4KqrqTIOWO6vygihl++BqW35cWy8yg4V0PbZ+JOTzu7WpdNkiAKX22JbSr+V7BYy
P/xLx0sfaVDuWrbdq9CbUXbb59Y+LNt4baxsfc90slbiKu5ST9DA1yQ2tky821yC
KXqQXK6tWEYnIJPyNZ3cYnioHHysaTwx4QyL8Uk1PM5P7Ue8JKWQ9AjLslGxPEjY
msVc3E1BX0ncSRcdOx1lcpwmBhKVObic6j+JR3ikBvTvDaQ2/6jIEvzG1sx2Ml+i
W271zjxye0+MG00aa8VZ6sGs2DSLAmZiQC9D2dIj9pzK3TTxA+il9nFgkYKUnaga
9wcgU8NacTjEL7oUeBZXvUtVo6pLCY5CuWEqyBALhoWElVFCVF/gEXWMSr452ueZ
/MJ/zAAjFnJduyCoQka+S8pGPvmSpd3raTO7aRCmtoPO1Ao8JeetoQtGhzbEM82T
SSujpvPrxe9HrTQvh5OlTxTi/HcmB/8l/nKgQHk8UGBu/SLeN9uqpRTEL0rZTHFU
Yjy6wNOyCfBQ3d9DJ6yrz1oRbUoOCH5tO8UJwVpIjo9p7r/C6fQb5ItKnOtDuoC1
yWOdmNTiUW8rrbDlrEwvMcEv33nzV8nHZstuEpPujIRQFwlLDfs4QLef3sWrFPbl
IVayIFeG6qw3l5Mgz3ljTqPTqhy5ZBLHPhJ6r9ZIBQ2qsz9zQQe/mFpbsTp82wdE
hMiYdw6YCabEqe1vaMdAGc+zAJKwW4MwD5YrPdE/zDtLVk5Dg4Q2o4p4rXdryV9d
pLACv4hy4jH5WqYyff9DXKxJlIL3SVt4a2wG3aPu0ylWt55dANV7m2oU0iUOGs9L
u82qenHskVWByYLBARcH3s93q3CYqpYW9jQpNSVevVWkBLAHGsuhzsiTThvvLZia
+LaUNiTf5dlJir34Ar9p4eeg04DqJ5Ue5qgKA4A6uqz5RnOFjX4U0V0ozmTuTQ5x
S+IzlCEdv8yjr9K+43Vc9s0qm7vySeTlOCFwQEIJ+Q6nihjJpfD3DX2oS3HTPF5f
3eyhExOrM3HxmBXu35yyVHj5bEzJGbcpu2q3dHa/QmLd0Mq5wVRarD3Ah11XDsOt
HrRC/Y55zGZ/r43JE9cppMSUYUsjVhH+s14Nc/zYYjc5Me4D2zhivyGqpr8AYjcD
SJpfEFT+oZBBqHzhCxUDLA4B+5fvnpaMKdYkf8pKycDRNY/WdZdMsb3F37BforGF
kqdKGbFejkrfrX1qE4y7gx3+9YZCaPfrmm4czsq6XJ0ylbNjJwrE7tnO+77I3oot
SGDcwwGIzxyzsVErwNyyKGcVfKlSRe5nmFmrm3xUxk1HfmHsumVO8TEeBRwEYhK7
DCR06PoeV9j+SzHTCkXga5gRrl7uZuEJ6K0sVcUeMjYvc7vwqPTIDl14JXPvLmuo
78BMDlejJEQJHYFLzDHaHA==
`protect END_PROTECTED
