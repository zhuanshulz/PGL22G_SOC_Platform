`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Cg10bBTpOb5IKQMFv16KpwUsIOmMbu8V3iua2tm92JjXRj6HQftbCxFk9TigbX09
EVrrD/pcQRpefDnErUlgGfXZyyfTYVbJLgtNsbZvtNoByy3TUBhyMFbPCjobomE7
wc3tGO3mXuVWzyW0yH4E8g/JGLI1S+1W2nvKzVUg8Zx7kZU0x//CwlkBFSOHzqH4
Y9nFKohATqNCbQLCkz944v1TI8+6hxFzYbTzwZ6cghGrlSSuanvF/jmn0TF+yg/J
YQPpb/Hum5f1k8YLIMlucJCcZsC8+1okssztQ/+YBCE7cajl+aNQzpLMPhEe1eLH
o3eRZgpNsLRgidVy3iFWgAwZR0Xp8gzA/0GWy1OTk/gJXBINOy5aSJoY7mfBjXAQ
dCqIRUy3UAZnKl33meWtZEON5xUrtUNu1GfRxByk0Jfk62tdct/osf8uKnDuYeUj
N1VTwYEa7dfqqXzNvHTyFc/6fCDRT+IegWOejvf1OXgziZBkaYR+6pMaW+TepACr
Gomi2vx91kF0Lwf7zFckj0U7Mf8C9w45ltTH/TSYfPDy1AARsj6rgyaVWpoZwgUA
`protect END_PROTECTED
