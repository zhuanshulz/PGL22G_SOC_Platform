`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a0Mw950tKr/e579k7sFFzsm/pzv5PPauIlTvxtHKpoZHSMZ0OUqUR4XfJV/5aMjE
vdaw2hGXqGGTnSCHr67EMdJD0pZn+t5zBcW/h2fpGCURWlR82Hk5T9fHzptXGlDp
WVeA8Ojnh4+/4oALgpCOfksnpvILlSxKnovCAw0tP+9nTfffwRrFjY9KIJg1fMcw
O629mwgauJVcKZW5yJReAkliO3fPQdYdwbyi1cSgiqPsMVVkuA3mX3VSVd3OtI9c
5C6xtsDR8LMBI98WFJPBCj2zEPYqfI5B1nSNzYBNTPcseE/idHH+VZJOR/tn82zQ
f1Nw3IkCeXJnZM07q/lVnmop81i8FxqslDo49ZDY4xC+lLdsOtu3n9uZehZlD+RH
0QfhG3TyUL4lDTwbJvgiHYsADllrHCawVnmriL6zwvRsP8vlOvD3z6wSHKkUwYNw
7zFNjkaEobSezv6Q+5cJFgkGrA9PeoXiImOtmwOX1izBOYlwWPsE2d5atGPEB/BI
xEpAG78sqWvehayuzoJgbyMrb8ex1OEmGkbECvixP62eolfbCEjPdYhwLoXg70lG
+jXWDKxxwNWFnjb1J34hPnTnfVd+RsVg63vkjePpHiso237uxYQX7PYzEl7zpp/8
ueRVPqCK5HVfluGorop3zUUUmHiYXD6loyYlIgt05J/UGHqchLzAwSpS6AgWy7CX
McUa5kYOXekrh9dEbjqzA0XjdPFa7YeEJ3S/FRnTkqxxz+dYEjwrJ5FuI3oOaMVx
2sTkIvgMAD0p9OeLtJTZpKCbZ/g0+ZARdejrUvd/nhKIrK0iLjVQPUZNa5fRBCCR
sy5070fq5T+zRR000Sl+ufYo/ef6eWyHmatRFd0eKEbNEjIHGKZiVOm71l94I0HO
p/HSIWxMgQxkaBXD7J+9B5rIdkhbRya+BaN5UA2X8vzvswNjl0bTqhnD1L5p5c8h
zhlzziKrLKE/Vierz9uy8we3R9sJeCS1NVYJ2HLKYyNmHCcTMEoC9G1sGd8CdjcA
Q72aRBghUgpBezFoQgFr8GFLvAb8DlDz5yxsHhP0jVL1hk8T4Y8m2DY2oPyWcvYG
avc48xSH+P3F5GzZfBYjEgJk4H1YYZ8JMg9MOcyw4qxUfzqkrunZY1/Tc/MhwZVk
+vKQmZhQHLX5+6sstAUFwZwQc4bpd2qcUm9PT9JDRrU6IxkztCRmdugOkIIjmRQX
`protect END_PROTECTED
