`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2pfPqXmYNnLNuuvC4YnLd1ZTN4+Mey39dA5kGFbwMNTncuM+hyT8Ix0SjZtf0hGv
ZwsPp6wDDGZOllF8zqiZhjTh6st5SsJUOo0b3P/r9Ej0GDJMRJmpWuHTW0fFnJP2
XCYNeC92w7X5APtqicbqPx+e0LptL9OsJjlYqV1iD1+W2CvonMNsz/O2fpI4Mvdr
DxcU4tlrPXaPQ+l5jjPnoeuNTUO/nGxa68etAYqhaTlbwSQAw1rgjKUZJEn8rClL
M3gRXHxvPnV0GP5CoV1eSCjIXZqypFk1GR/S623Ao3iaBpnd5IS+SZ525oUBJ9Pr
z8SmwKhE12qmf0FjVOCnw9kUjDs/Qp+oL0hz0NcLMqrrOCBhl1FiXl5ARZ6QFEIZ
UgMoDoNTjk9x2UAtrjzsRI9fIpYL+S7EmpitdvPxgYUM/6QUB9j8pf4e5Gxokuqg
OPm4GXDYOhuMN5W81GjAjSa+G6h8dRaHdrNW9DNaawHmm7vT/kAjbLcpxyQjm/bL
QqXdeoDNbGXSzFqUccWYog7FPTxq40CspWBkdsl16RxQcHZwT1vmfwMX6HCnge4z
Tx2q+RpDg5KpDuSo2VlF1miNYkrlU7/Q/IKrbpBe9B0q8/ZV9tfYXfr7iHl20ENw
NN5fTGJG9VEWsX27u/zzLkRmWHsetDT0xUsnN5ziUw/nCR8KKZd/gGzCn3KE0D9g
mA2t2faMyK6pw80Loh0xqXm57+nzm228xD3If9Qlgk6oXbn7dZ0c7yrOS8AORyIC
X96qWvx2ZIgFB+weFCnDfTIGoIXVFiEwcomNi8U2ntQqlkTc2PNDlyugHeLYkGCy
X3Vr1360ppjTTAG7Oe3HgYNGVcSHEy/CEaeurD342Z33gyVfUcCY4TJE+TW6buMn
uruDW5IDMpYOsLyDZYAPfvjN2Uw4yO//n4KnkzI5g4/NVDHOgaUaTMzEAZunuiGQ
k2DY5JAI+1Q8nNRGoKW2EPYgEdmmB1xwVf7ByIR4h1o=
`protect END_PROTECTED
