`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/C6UMrvbt/PFXHw+1+CcOAY52jhlamiZQNTaUOjeR7Rpp5WXJzJuMspLrzcPr6KD
9P+X2y/pZnrcLr1LiAvr3oArXg92QEpNKE/WqGTu7OpIghhM65ir29eCYigUx/q3
YrHfHbEXSMEFrT3EOaKWQhgoEYThAIyQYVZfNKToUeuXqlibVZ/yppW3YDiUYWSR
wPaeucIcl3npIFpRlql2umechMnQ0Cq+L94vuVXbbMeUIqEjWVQ29R6no5+rrKse
w6WULgMvPnaFsrR7zuYUdCDAfjYUKHv4DVwTUHTCSplyVdSDtgRKl2FV83HPWtVp
4k7Lxn/z4i5ZbVoJms6br7TZ+LXDTKsvP4j2CzekdOKTJ3wWpZqOL6krF6AUf3SN
DU45epY2bFu4kmrtisLmw5Qm5msliwS3j3SlvBn+BF9a7c3dQV/RaUPXuc0ve3lA
kQ2DRdRtFOrELM33JMxkc14Yl+D5jtiCru1JtQbUctZEDT3bnQuJhjEaOJfnTF/O
crlxdaDH6cm8WQKnFwiZ+mcPF1HwGWsRrnN6mAgWGwMeRVB55NM4+Ldr6/qQOquU
Ekhhildi25MhISVh3wQBc3gOb5ohwtfvpMLENwOQ74x/eBuYrALRhBOK7HYbstFG
vioGxIW79Qxj1qW5M7ZXPi3r/wQMEMf87Vj1EqagZjpdlip3qOzPtc2AeHrj8V8G
OYB4wtGFDLUHPjQXvMETnc1j+kZD6ux3bXUWyQdORLuLU96mhLsshs0/2JpbIqiL
ekPHt/P6lHT89B4pP0kEtCdtnTbL+Gi22jbdkDaLzdvfIIY9eIJLPu8jcSnF2YB0
dFx6stpm1kQwEoGdaHoF++mBby8U1euC/FzUTAkX+uYcj2cogGqjxcgSwDRzSAz/
d+g9J012SwHSak4ZrAh3BxwPRqXCGCn3ERf+zenGHy2ReuSa1tdmj+A/zx4Y9gnX
lXkAiXjCD5dbnun9UBsKFKM9cqO7sSFf5r/i0QUurnuXHvzkZgvRPQI3qBXNymnZ
pTV6skXJO9prPZgMpYXJKnC0qPOGDbrTqDxwPOY8HoIeSceJGbV4ykEMbjqZPYDj
KbvYQKlQpj8o+QJMLVc5odw1t69LINxb+r37SBGu8/MjBsPMm3vEDQiUY1r6uYeP
yjDCXLa+GYpRZN2LXU+xEw7syzDoREU1NzTdW2VfTc+IEFHhOF0/XAOeuPAwDd+Y
av6cTT4UwP1Nb8WNf8kFOzgp4of+X13svteBbNFa2bF0PNK8UxUPL8AIBY1v+V4w
+xvo2dleNtJ0IS+NffjfhBW9heDZ/OIkPXBXE6Cr6SaYIK0qjuRFW+omN/uVzaeh
oupm4AvYhOqIuwPRXIYcc5AAnbSa4cQCay/GHmrQk8N2nK24fVxXH2TLX2wmGUAi
SQvEPzYTAjJzhM5wzZ1Tgm6hqcnqzP6egBV8YZzI8AtDRWYOxQXM34ia6+EODGOK
Ybo8pRsMva6Ij6+nTiBemsMnbbyzr8EwyxfVPoV734G5dZG1QMI3KVJyaU44kWn8
m/0LqbiqPuWIfiuqw3gYpax9m6k1hMltnqZibo5w6Gj+c/W7ccSSNj0Ej8jUbaug
lcf5lvazZKe5kvwSvyvWAVdbmoStkW9z+BBs2SAterCQKJbWRJtHbA9LBgUu26IB
YMq0/NI1kvhrLy4F7Dns4Hz8euWC/+nvbl+ZB0VUDE939vsBAsaHEu/1dfMySvIU
/PFvquOQmFOK4bFjZ44QNjweKo5yWRN3rMt3tj+34Q2GE3KycG3/9zcA3u4mpZGn
UZua/fJxDTL3mlDzb/jHq9rZqFIn7kcWbLOuEYikvgvCT6b3goVHHrGZeUnOxmBa
7gjIRdHdd9Ois/7QMXJ/I4MuZ+ZeC/mUpcAx1s6fBHnlSbpgEYTd+lVwfwTybkAG
cFvzOmM+D/82UJHtoTJHv9S46OB3eQmEYPiL5FwZAlrs+aryhsh1PJjNjjZ/qrC3
N0bGlFDI3Usu36vt7pn3QkrkOq1bV8KXdlDLo2RG46yj6tcXMsgxNrVuI06BNHgw
J8dKWTgV/ZYrxd8FSBFCuENWRUY0JQJA7hJc57+qSm8hoEOX6xVTC2UBRCMl8Y0c
1TH/rVPrkOLwTN64sDlELbZqjPT4q86wgDo9yGxPDzwraPnqr1ApzJj/YSz9OvrN
6IyJM2syjkWTA8LcWW2S9P5gqcSGFzEb10MifLaWOaCXxXKjzhRyyqJX9w0WCFdm
T7V/oyUxDfB7TYUH8WTi+U7NH+w3T3dCZA79YhUNr+2tfoL76GVLxBDJLcI9FbLi
t1E9n1rscTqlC0qg0JahA86GMb73IQnr/w0HXbfUHcpYeqhgzHnewgRh1B8OjckT
HAcemfCoNZZPru6lifQPac9THjH6djR5I/QmPzgtMt/TQJPsqG9uvHmckIbJ03cg
rnIgox7cBO1r6xdCkVvFRO1s+h0JXAIOfEVP9X2SbrQc8YPEM6is2xvrOQTndRb6
qK3nuTT/DHBWaaRZI01V45AZSv/R6frfqXsFTvYdX69IzwuI/vLjmICJtPsIZV/g
ZLbfzD00kOSVjQ4EK3R7EsOI9eqBTj3cLsU5GVSAMLBTMWu/549KVwcdvwSQhObl
+yGPOcDhkr6STvQYR32lNDGnPcjzWb1WUeqlLVolcqfF1NBSDb/nZquEFHaBKAEJ
NJ+tGDYaFJf79/+QmTARft2/cvMpi8uQMqspr46ODf8CcT2IqDmu6hZMf+1jymbD
jD/Swejo4BurRt0c90z/gXNPhj3ilqoamSXtFVbO/Bu7YtpFY0j4H0u7dYGScWYE
9SaWexDVssOxwYoQLp2NHpCXqRkBdQ4y7ClgbACAgE2cf46HexNLncFrNCoQr3h8
RTlR0LyVIe0Z2g82ibX3IMxlgJ/goxVZ7On/n4KLExHYFmRQxWhCE8yHgkqAzgiv
IZXBjDRqPHFZNvR4JhVNKrjpNNoJO1BJNXsxvh6gMcPsM2RI+yPNMN7La92GfZSg
9W+3fpyLeJhx37/BHR6Uae2KheY/6AYB+AWOPISe3PkqMLBsVxJBfh2x+S2O1Jv6
p+XZHa3zKuH7kYKDzP4An93W2gux9tQzOcgzLPK+59NbkBo0nL1dt9taXgFNdOEl
gyAWVfDTnLEOP1Q4dsLg/tDATgJDgPKrHOCZiCtmCN4P3Q9zl3QKtcDuDDaNo6fr
eoiqigOX5K4zM7I9/EeO+ZuK8DwEsdHBWGeCvY2uE3ddpjSHVKz6hbAtcd3znzxq
QIBYadc1Jx9qUKxzmaey90k0GQ46OXIIySW4g112ys6ZkG32vRCtyxpRL7O+YaPn
U5aYa8LE/4cX2BtEbotk1NAb9U43qVKy+54pwMNJAiSqpJqjgOqoAomlAaq/l+iX
9EbnyoHFfSxZXNtOv70o+JIPIoZ1pyQh9JmI3rEbbnNhf4I+HG4nzKwi+UO2tGNv
CvYAhjuNqkzUYauXamLU6eWjRw7trjg6D4FQVZwVVCXNYEhkDvPA0qq9Vu/nndK6
4s3kIZ4KVTkdxLpu0p56aa4BDSnh8g0NfrKZzj25Aphq2mYce+0NJ0404WhEkqZ+
FWS/hCFV11CNkXXExJxkHCryFfyrQzDGnC2vzKUwJ6Pmq6BsOxMaV9d9JCh0sGYS
YJep7spcFxR8FQ7jpzjsv/0T/bDKkbbTrLIJHFu7cRJbAwYI0kgs+j1LCjSvIqER
U33ofJ555Pb8t5oXgCyrzZO/WUDNOIUEJom6XPTIARiJFHKI4kvh3xjQdInP+P5M
BXKl+Y7UkmNop0Ea3OsvmDZ6QZ51clIZEbiea7Bi3qQrw/74aJwfMGdGKpMsagmG
+1u5WxG/nS+oWg7F3XtBM/6OVN6+hXbP6ftMvQNQhaXxRvk8Aij0euHs82zzaofT
suxcvXnE/Xjf4XoXRQSxDTES6FF8rj8irJfpk0xzwWiE1iGRVP0fwipUO401cJVa
vRzi+2sLM4QcqG8ZNoZ1g10WoEilDrQIVwEz2O5mduxu3T00GJnx2rqX+Prd55Qh
OAngx69Nyj/mEjVvr9Afl+zU8yFpJ6QdotTvDjdzV5YCpItOqtO8nEVZmKgUDwrU
C4ILjSjEnYLNUQF7CQ7miwjhPB2IZbLZ2GyAsvxAKPgFPfPWPcz6AKcFubJPt/7S
z4sSno0c1+qHSNTxW5/dVDDnBst/xUWqWeSLizJDYvxc5uFrErOKkMbUyLjbNfCm
8/fFUrB0DxAWcKWwqBfWQTb4DvraFWjdebqrx1tFBauCtoHU7KG6XLRKUCkVmBNk
iwBt0Z5En8brAwKsfkA3/IsXgOaIIWFP0/YrwO51m0jZI2pmAnxxHKSUsEWs+21L
ypXDM6R6ur4D28tZ3QtzEZgwBxNbYjTey5YJFNV4ctPi72r08Z4RejYx2U83Jc/r
CiiSblpIfKiEHX/owBwbgsQdp2U06hxbR31MsEkxxRttgC6sEtjjHOVS9JTvqG3I
Lz2BEqfF1IkuZrgokVIP9D+6YXrqr/tMBvsN1dIIje9GW/Fmm8P7eSGV5O82EHMH
5I49CVrbrMuGUem+np0dwqFGdZQHd8+UpC+JTPwRyAu6zksD7ONICDxUED3z0YZO
6cULFbkETcoxlokCu6XhPvnknibNY3GaiC51CGhvfd9IjFKbpshcUP2ic4ZngG01
q72plwaB2+pt9p5ATXwYJ1nvDu1lP20OlJma3Bjr3rQuytZmAsQJ44K8RvWqvYzM
MfE5u3WVZFoOwXl7FC9Xpo4bWNI+fz0sAMy0CiwES0R4PH0+yPAALWVE8kxKrgxi
D+vouwykc7HeJZXcofKesCxrOygoIt0cwEvZMMfJeATsdciNmg+poQy2I7HtLT79
tVz2F6AWWoEqdypVA70NklwsFzrjoXMeeYbG8Sht1DEsP+LjPtASJ25+01c7ne6C
RGP8dlcn95URfy3pkjYcMkXtBfj75/51b77LKov+9xmxqe79HA2a6P9d97bF3GGA
L0u7qCrEMF1tGSEqs+cF+1I2fcXzHhHexQTJnx1xsbukIHuvQ7+VK16+Ol5etryj
EVtdHuBok2IiVmVAQcRQYgxWEQtDNirXNPdOLfDNB18wzIxhYN/1A+wFQ9qpGeI8
riHrgCjHjC9T7z5LBaE4lUJ/7gOdHr5pWO2+MVgnBWozk2x9vXk/JjHsQRFdjlFf
6Q7kT++szo03hrfQDrcF4V1rMLOzBdLcLQP283GBrHDzhmwCdxQUZgKJSl1rkZ88
aB8DEi/iXJyy+nNFJpPNSKWjdxh4Z+wB5/pip6JtWTI1c2IWaXu+1h5DwzMB8C6k
hmnZf91Qj8OzmQYJi5w00KjRRqXy6tFCBuZQ1eJSyujy7zq899KTS0Caazu/rVDb
qKkIpE9Tl0h0+1X4fFDLBg4jJ4V1Zc+KpwV+Tu8bwyVlFkswYOx0RWrDYkuYjSUy
NEVyg+Y+0gE065ZhDX97qfHQKk3cPEcgzSTD+36bcsKCRkH3K5zcqQ64dw0ywk66
4LHt1JBTjnas+vi00FyuORqzJp4j56gwj8laVTRlqi+bb9SCMtfbYCDnIASHWTyA
YfBK3BcXEhrgbqzZUvxPI8qbUv+Y2D069ShyVS/OBWkFuN/sZWxNYS48rXBUHPSt
85oW1SKDaQ9pSiw9h+B7uTUCKdcs0l08NRS/T50miYOsPLbYJXbiEh13/rrIBiOk
d+Z1Emi8Bpp+JLHSrp7bfB47HFrWCjlJ4SdtMBnQhHXabSXK/RfTWuXCssa+0/uw
/4+CqBSf7eJL+VFp/PiynrsVWXSqp5sJjXC5l+odqYN/Kk7PYmhN9MPj8YsvFJvL
7SgINezq1uw+cUEihbrTeXbkzSe2Yy0KgIe0iQqC/75gIT0sDFuKPYow1fpQECJX
dXApE4kFsJUongqv2P+Tfcg0ALOs2EYfdsUvjOQeWEWGWDjx1g3lzlNmn/0AHCw2
SlhBowlYBxY3uMBiLOCyf+8yrwT7m3zZe4a/DT9TMR0pZXsPkrz+s8Kf72GdI5qo
NRgZuLtaGx4KpLMqX783E0RrTERC/GdwkKWaDWpAJKzQoQCP30LfyyuRqn4YmLCO
uTqEEGAOcoYcDB0u28WvuU9Dv4n80NkicqVIIvxWAoriKpOJ7GU43RardD9d7u4S
l456FFdV9pcrvLSdec+32rV9EhHqAX7FYSxiqJkU9Jxx+v/KAJMJSshGBpHsbIIG
8ideB7elaWsAztfoXH77eo9pDxzupPo7DHrNYQLFazDcF7UKoKPLzda5lPW+k8bN
W15m9dDnfQRAq9cFxVHWmfoMR1vsRQsceI/XnLczzFGM+GCNXzxQGn832lHnVRiN
0Eb5hxRXf587ru+0MDnRf+Ggk2lGFRJ+PxAso4YS6dkB8eidRjKMkaC5jFg39+Ay
NK7NjBGJCiLlFI5XqRBoEN2rTU3EQbq2FaC0iM7etneMsAezqMil+vDT4J9FVLOO
mxUevcEf94PotrPMLg8APZPXt2e6qFtUiyurkPnsS4zb81KxnmHSkqcf/gDW6Fn+
rprlvrK43VlfTPXmX61PVdKuVGtQG9Cs8H84DpRzgxbV7GALI4rbn35LwYv7B3nH
5bwIm5ja66HWVXyFQn8+NpazJtGpfKczF9pR3DEpcQ8yHyfebhpYMOnJa3ta2Y60
w8+SuIRpnCaEx1NwhfY+15MhMsO5wBxIQfTX+xc8/Es5BcZGT9s6tKQOkZS2SzZy
mYibJZzsIg3CQYIcP6wMwxp4pIPJeIcsXrq5fw2LIBhkNiFQ58qLENrxZNhy/WeL
hJ0RLHVCU0KAXNY1TfsvaxO/K+t0U/7G6BvdL3eprdKJVd3B4ScEIaPoMVRc+eIe
djp4WlXPqRzag+mG57taR90co3pMoJj9TJTAGFZOEa8SQiHqwnabcXHXLWlDq4Tk
vTgkuZgPJcK7V/aznBVmgQ2uenu+qky7W4bckoN116jrInCuPl+Lo/dWQybklN6d
/Uy1+xTR+MwBGhTWJiP2W8kkAbtmrpPgYSWsaowD8zYGARVMPxVQPkwEYIYfVTJt
9qWz/1bFNUtQJJX6YBDjKqDSA4bWlZwwCNDpotjFfGC4mZCsMxG7PCwtlJQXaaJx
9C1wR54k+oI3cWrfT0s8kP9f8VafPJah5MdXYbFKdQ6H7hJ3b0Xo0XbzBjP0WTVH
ZvlVkN0UoCYz97JN3rHv7QFZuE1P/yL0gEPECmoZJNRFe0Yb3PjymZMrap0HlHxA
+vKzgrdEk6cpiN7GuRU4v/s6zQCRkUsSxSNeg58XHCbYeC+ETnlRNroxdbImyApr
siVd1C4VHqKq9pO+kLoSobZIHqUFG79rEnGLHGSYxxwPfZJOxCESrBNIkkpaivBH
B/pErC7QU9jluZgSPykXusm8elpmjo3UjZh+LLNhJrwRY8N1lwkoR/wCwTAfPl76
xcbQEn6EIQ3UJv7AFcH8cSLLt86apNZQI/dJ5isU4OHHezwCaosJzt2gzihymL/c
lcJ07sjmCWwb26W48p6OPcKqraroxQrsOca081ClabNDwE0RASnDuq1u3SB5hnd9
kdFn3XfxqNsmWVX+JnNZzeCo7XVzR9okOGJ12vppEeXGbiivG5MwZsfiUFAZbuKA
VuWnoeqqLYj8IoMANYfmDQlUsEWw1K3mWXDMAzb6vsJ+52C66EUU/Wyfkr9FWEgy
EQuu7GBN6+vfLnqnueyjXs9r9e9acdyFEb2oIHG7Uja4Q+Mwk84E+WocmZEAGpOm
KFaGZAxc9OZ669Yn7ro84h5V+SIy6nLrwrIfvEAeycckynQX4XuVX1EX1cbPTHkF
1MVkoUS3Lp6rGcUfHSx44MOTkFiKFlaASMWDkhaDPyL8B14BiqqDrIJTCZJNFInr
g2wnkBTiFde/D28tlCDOkIrVqBEfsUcNiOKM6yiXm+yfcrGxYHUI1pDY9BGf7T35
7gnIX0hmhlcd0RvkGiot02h6qs0UONKjr7eTG3MeJht3xy/iI15d3uqgkA0X5YmU
rO5g0LL1UFjBm1u5mN0maRU8A39OL0C6zt5TGPj0NukWupo8L3H5v11pyTo6X03I
BFSrk66D3HRXzWM2ATXQGNBABer25pGvTEYcijgW7ME24mAVbopic9EGtiRR74Cc
pwFzypeB4YVt7JvnvG6gmRCCXKJby3rqnH4ueKdNTHB3nq3UQGjkq9886ejCmF7G
f2LfEMHhDKIHto5fvg8NSktmjC1Ta9JfNuK7gjjRBYT0lfvxZyZ7kPSiN5khIGKf
nSGNh3/jYY4OtVYYXHU2u+4yUBrIOU5FgNpJ3/SaCskC3hVhgs+/xw+6V0pqa3gA
V1ReMDg+tyex/HvDBevnAmrPOv9Z7Y3bj6FE+klAjEGBJghYfnxsho1h8vZzAJkx
i2pv0HuJp1e2JIZV6DZFQLIIBceM6PV31aGTjhYfipuXSRCIOjFUq3Zb2bOxhSp2
cFez0mJGsKetn2cOOwWRoU1xGf1ZVHnA5jRzddT4YWwn2JSw8uukS0fEfCd/Hnx+
oRMtIi382eVQQkg/ZgnNqmOzCeqpuxntsHIoge5SEwZwN1Nhu+vvvrFCCzGNiI1e
AI7uxpey6iRiqDP5Bm3DPEaMe95ogSM1HQCxR5alzJMQPrqYlc3hBBT/6dyYTO/3
medhMmXmSvhGemThper0+t1WVKvkPPtEPQDUG9Utuy+YABjbJiOzB/+fd7h3wJ/E
uYfv4LrBVHAn++d9xCvnzQnYE5Y0jFuQg2RcGlofaCu4v/G28BerTYGMgR2M2N3Y
jHIqYe3jIx7mOSzlh4VCsEGKFS6NL7yGCmNlXGmok0d0XMSpj9Ffl5DPqbfXIjoz
dQPcAN2T7uLSxs5suZGfstzSdRVkAGnJBPqK3Dys+vjH9RRZmUxrRp9BzWN/y6va
8p3ugv5tDcUHsxqfPbhpSeY2kOOJJ4z6N3JEJhnQ6nXf2J5DojalMGyeBH95yXNu
s1BNTYmH3rpClF+XqVks0P1w4Xeprgyc46tbWXRlE0Cw60j03yCgwf/vMnh7apGD
MW8ZLmUHvMOu3zZkNTispr3PL+IIJ6LDXyCeA5lGk6651/LW2+sxXLPUlsps4XiF
VAEc5boPHIs/33gNJ8Oz9lDOO1AgA34m4xy7CRkb+9fS98h5XvZcqxCYjqty1F7S
9A+VgF+CzQBhhpkZY56NSRJquaRTf0NKnzc7FAed3ENRss26PgT1Cr3AIG3XEu5M
D88toui3rmIy6q1Ew5PgxcHkGgZA+iR2c4/98KtmVQ9Z/9hwZxqNfI58Mp895d+Q
mxqSl8k2gDrPHKD3/zR2DtrllXMwf32BPntWr7fKJ9lk3lXsyKDvLc8LlmH7OgAk
n6DIPOZW2APPx+55dYWwkys3LAL0oBHPLL25umH438ueGae6emXU4RBuoTiw+/SC
l6+PXYVzMC1Bp/gcDkc7eVgASrEMHlcHGgFj/XtrvAGCeWmkS72GfmKOgjZvcxNl
XM6cXB0ziFGGisv3GWkNNhNLdrcREVHMtCLvwBdnFIMD7OLZEhD2mx36yf4JCUtJ
sdscMpB1d9+Oo9ZwJx01Hl2b0/EPDlkEuospdp4wWT0BMvLzua8WxzSWZwtv1ZVU
AKiUwF847Xs5yWttP18jWULCJUg+cnDvwVbJjTzPNtVOt62ct2yTZjHBVCOytgXU
1PdERh2io6be/z3Z3rpX2Wy6R2Br4fKV60EXl9DmVouqv24o0w1ac2sjA9rR0iTJ
9EQEbHj0yArBmY71tKsizmumH0IbOIkAWe3KqIx/DqY/6bLZ4GiPkBrAKjGpFAVj
ck9+1z+lYy9otCHYuibLATTQsGITMhrlt/grLY83gvaRX+ENDS1E+qtcI4ycWw5H
Iu1qFN+zZGA9tJdBG3wyzmw+gCIo364wME74M/+IXFk1un08FE77k6v+75lxda6b
2nWA/ZvMrcPHSDBWPi+9xl6sGnqlrQ6FS+bqDcD4cdVPrs1GHJ6qLGyAZ0lLsGfS
u0LYIsIqE1LAPQnYEWQOgw==
`protect END_PROTECTED
