`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GNYOnLSOKZ9TU9BZLp+bgxJq/X5kVOyimRyhX4db3qG/Fag39Zl78FTaSt5Go0cf
ZiSJ7UYwH5AXNrBH5mZkQEZBM4sGl487QRAK2QTVGWdyJS0FackxgL0/a3YxIpVr
mtoyAP+ANT/aIKZ6Eec8sryaxWuiZZkc1QsU83g02UoZ1ECAMPfMnsmfN3b0h42u
ZPkRCIuwmBgraYEMtSu6OUQLUZ+DtoiD/feDfVNDGbB8YW7JXDAYBvkzEn4w8+2d
kZSobnlDO7cO/pWMLIFkgS2NQps73A+L+2oDMs8xrAUTXBkp6QU7XuCd9uHZsFoI
WQTiunSutWacTRCiAX5YDbL746qTHS9Ta+avdMjTzpwu0bl8W5hN1rhZCe/nzk5f
KyWwbbvBwP6wJKyxcyvJ+XPzmu4G23t2Qjv1qWsEupVskYi3DrmDhAkEY+zL8MwQ
MO9qaLoDIB4ToNvAZv/3zECglZ0H8uYy+9CUUuPvbZg2BuAbyE5xEOI3uUiCIxVo
OP4rzB7GLgshHhubsCKlZWF3H4lKJLPZFxMzLofvHdzY66Nevk3vmdVQjdjRZJLe
TRLbXb1jAGf3UhL+3Vh3JmDPcmUqXjXof9oDysGV8bf3QNBJcOEbKQOvNEx388cU
WS0vbPTmkjLuEsI8E8HNz7K0t8+l37HzwBb2nA/8cOgWUYzj+DQ04y12EAfpE9wk
4GbxR/mrM/BgjcTaWNKOlajwHPeElyz3j2pRt9tT0alD0HJeHZCT5C9QW9A3n/EQ
ICmURMtBCZfjZb2+Q8vTjFs9awfb6Fi6Z7LWGkViZvjFntqcn5R24fwoKqBthmG5
kMkihFJosIHYBW5nXiOX8Zp7c+TD4ffm+F5qIT8lEbIvydeRlEJswYojj4YcPGEV
WK47Al25dHnNJJ/uOMwTyiTe4k57T6CbSvOVRGqRY67lC30P2DlVumx6E58Is/ND
Vg60ZhWz4vE+HCSvkrZAKMK/MwZkEO1EO+wwAplucaOOjta7zWwBMns8ABtyFHoW
w416VUbhJVeVGbgjJb7Uu9EkyQsxQvGkzvjYoBcbZOzDhM7oHLyvcGghBCZdyP/M
s/T9z86SKFj9ZHCFSoD3+XKJ1ULFujZxW5IxUvhL0mvomAn5BZ6SXnEPh7BJDQ58
lYaq6lbWfcXbKWWwVQPwscP/PSmozv78c1lkPCoXVO/i4jjrXjPNrnQ3b6i+Yldl
ONLp6T3XH7d6vxc9ptYofzXN6eRut66p+6vtqDKb5KYy9cVDTVyMPa5YR1ogfuYt
rMsDoMfJm/cDY6OQ84IT9TOWjAa/1I3WvhT0OV7VUiDEjjSpkrhLLcPt588ZAciJ
EHcHwHJ73ojrK6nJLDJjxuK3bOyUYBrUb/vs620fGlOnCvKTFBVBjmCcrzhHBfLv
4N5rrXhFmmywa7Smp5GSmLrsGNoovjp3FjXtDDlNRKlzy+tptuzN8SeAeNYPIaVN
ku50doVlEJu9ZE7qc5RoHu0Inm6M2nnieed6AT4NXJerRbBNjEEjL3RHE72h8Zw9
KBAkuNWp4dmWZY41JTrXrYxpSgitK0oIOlW2nYlJZOfbP3mTQKQNaSxffHzh6Xfn
kmVAlbMpJDANHDxUpU+njNN6xGNKiS6eKdDSOnNkl4Pv42PhTdFmRDugoS3XTQ6T
EtPQ0SFUQVR6l+YUH7XgEcsUqLLNDEGQVWyHkK+BMhMmKpMUzuAA6OxpyrLSJJkX
VW1eCH+jO2e8zybMChlNmxBtvvpUDe4Noj2wvWmmaMkh0nCUsIi9yQNqa+iTgQQu
f657f1NEGkysk4DHikDROC2IGKDwWwqrZI2JZS3ukLmby4gfh0ZOHZ8tkqnPoctc
EsXk3qJ5iXNZqZ+OJan7NeMDFXhVdB3Ir6E0dfm/VADW/VPji5d6v0eDnakU5vdK
ufjLi3w5MFFYZMj+KR+SlUWB6/Bwhv0wZ9KIwRqGf405WsBKz7fVpnM/HWsD5cR5
wRQd1+ClnxZ95zk8FL9DwChzE+UWAgjci5UvEyuBShsnbhhYXRfoWYyy+KVWrkr/
9tge3k5W9zbjA/fkZRiSOrQpD51GBfwd9HxDVwZ3AGoaFmN8IEQlPk0p+/tmH0G7
cVJbuejiUqbocQK1YdQlfw90iGnOp/ID2C5UyiuPPMleJRPSPSb36E1fXUwahTCy
dZvMyW0zAFjVI13FNNKQe3NYh3SnV9AuEweDGj9iPv/ETrLns2l4QS3QLj9wF6wK
fvcxiIKnsQQvEsfL3SzxkU8bPHqUuC7FUWmmPcN5Kkw+6QP5dQM+t/PSnGUci9ZV
jH6T0TP26tDt69SWU9+rOu6dGI/NzU+fYNLd0vRiGhfCVUUxNuVPEZKecK8/9O6/
1DxsNJEqtC2b6K1dtveeUDggil1tkKBCLw3EVYbU5MOS7vy8d0c0ql81HALOlrRE
2yZbpWsBaBpPRctHHy4ZsGeq/5bLT3Utv+4ViFzwRgt/t/ZBUcqNy5zk8y0FnKib
kb9H5GqRYNKGDOKy3ZOb8b9U/HLk9XLZ84BxJx2k05CnsIASzgbZQBu3jlEoNYq7
ay+SGTqAPZ/4JK1oF7aROL9iPkUPMcG5Ms4fo/HLp8IRdPy6AgwYmQfwoHPr+jqh
z6V1cFvfYn3OC77crTNMh5sDaB4T+GnDa1i41AqGi8MHNQZ38CzQrAl5hVBva5MK
WwwS8ZkS+N1rsjDiPB+7oBZwj32fn6k1at4ySR14Q6n32rPdaFnI6hLCERyspmAh
IcYD6zewr9YEVgrSLqQNgL4AQh9BNPvXcN1WjTjB1wDs2iM018dlYeFWccAoglC/
3jY2R0G7Sc4ySK8c/ByNUQyqigqu4dgE7ZAb08yNw3kmSQOnXp8ff4FoVIyGoWoK
HUb5D+7sSj8pYWjw95cUoH9jLSaaiWr9sgXjznPA5BwZuq3YQxLKb4aFvhHMjI2b
g2eetXtlQR9s97leoDAnajitLN3DMHVCHU4BuP4QCdYVjrfiYTaeKd1DOYbhyHiT
/gEzfGQQVQ30f9ra6PIOzA0mxFpnve+14Zwn1m6++Hie7PPYElKOVI2Ax59x4Gf+
ZLmjKQBCKVeCoZot1nXhhiPr34kl+s6Jmka8+ilNTg+Dr7bPRvOyrUeTN7DFJPjO
wjggFKEz9b9fMR5p/LyK7PDoQ6NKcwkZ98GXk4HBADmXTp2xCV573mwKKvzNJxUl
T4a5OgdoN8TLGCiY4TBasBdp7jjcXzeh/F7Y96x7QVRsm5qBjFoCRVkW9wk6qYVk
1tolVjxi2WX6bTlLofRKBmZ4Y3Ui0obWAJaTvv5VQMx++C+zetOlGloC57c39KJ4
1nQcBNE39xZhYtj6jaGafBLhUMY138l5szFisIOKEh8FuVcuRL/Z2SF/INXg1Cx0
tz+gQApOb49f0I331RLe88ZKkU0Pk9E7xeHYzW6Ni4g0IU8JcmG/emb0sWmWPa47
RCIByn6dfiFvKGhTLqB4X4dcZwlF9zIrkK5f9gjk4nkdcDHYq6zk13IcJkPy30Yi
/YfRdQH/UySOgAoQxRej5vmN9RmEib+pGT7bwqIc6vkYaOko1xIWqSR9E2eLXshl
OiGFe/7KshI0ZwrL1YqctANn+Kf3DuH89iIp1l82dv0cOSWE5tx1paF8ou8XGv9o
oh5pM2ZH66EGyUNcXTl49R2Uv+RQfvm+Bknozu3Fc8B+nEk3oGZQlPTcpxJM3P97
4Zgl/KNQesT4xSmUjAITdstm/pMYtR4U03fb1IdiOIkt5S26LOEKJdX9+wHO931v
UYPF4wQAPZzmrsPUilm8hDnjx61QMWU5IxBcN993wE4oY8g76afDYFH6ACqU4Yxk
zH1McCxH/HM+CMEmzLNfrDcqE2LppzCDKeedhmGFHnvtliwrtqtjkh055j6F8pMZ
05HVNUAnA//2fhNiYWcsQm8Ma8fS9v2I2kPwZ66eNHE6OhrlsJhqkrOKjYatWXH8
wgHKyFF3DFMYwQO4Z3mHo+Ahxwopx4S5GnzgY46i2mr3I2v7KqEQ7j8IK1RcHtmA
SGQfSRni07KvXbmf6iDxWr/83qrxPW7A/NSF2V6Mq6KBawbJlHM1rGnMkFgQLAWa
OHcZqvhpSPnDa7852+W3nXEV92P7vVXXwuJXMQgJtheJYQvqu1W/TAlVMeUmdGCS
sef2LRmJ2OuksbOrnEjHTvU65+2y9yDxxQtLksoj7G1MlxCe4Nv6r2KVTAMtdKi8
8o+t0EmhItVe9QvWEDk1ZW1wdexNpgXKWqLLa6oZ5BkuSlQNEN7eEHeeXdV/rsSI
fPDG+9uJN0k7bt3oIPrq1DcY/xzfC1Jul1tvSqFcXXaQuhDTqG9CWYt0o5BGqB/x
6EsfHzh9DijME/5iLiUT9WRPrbA9mV15Xqn0HKwRBYGlz9g1ECLbsux5RMuYEH8e
GgD2wfUlI39gB+GDTIGxl896GUuNqGGzhxnyjbGc5QarHTTy8qvLO2cK8kEcVXSX
Pwrwkx1lZAPVcQPOaOrFWBrrlYzikT7OJBrI1V/Q4GpXboliRau2PlbFAYaXBtZG
j1Fjy9aj18oGaVtHOujqhCmR6wv2Vcy/Z/qY9QHmYrZaenFitPYAAifqDKR4NCR1
aVa0SbB3DAZKkOC2IYKGNW+BNpWkN7pocy0v1LenBJGl2euDrGxzbDqH/1dRj8Sb
w/cRnkilk85wN+aFSGqBipq6wv3SDplD3CgBEDhBoStowZaMNNDT2PnuL2QTN8t5
nOWisArgL9cU3ZHehIGpkSjF6PySQdgMwswEci40S0majRgD2H56TXDwT4FfB5rs
RXO6OcZ7uuwJY9RENoxBGAp3pMi1T3DN/kHIt8rfZlmBH/sitK+R15D5xHSepghY
lMY/Q+Mlxqkn+8CYh/t9dkzCM0fJKvnqIBa1cIs6bjh3hSr40VTl3cOncKg6lAjX
MdhB1AvcizvCO+7RFoSqdQaolRGcEZ7wYgnLVsIWEN1brP57eFuwqKB79bgn8H3U
rWj2OeT5DYRXMWX/9moySN2F9y/ERyFWXXgThyWoR9Iq5lckIoR7LuYJvo2z0q68
DbzuMPHXl3Zb7TIQpy8BDAyGSOWyOGcA+HwEAAl9tPLkCJc8+zNM0O14DIuK4uwz
Ln3urFXoGQNrJfnC8FlLd+UQeeFKeTOwfKdj9z1cEaj0XJULEX2RK1ElBTtvLaC5
ZJYIEjmknb9ZazM3DQ5/Il8VM08wFlQLmfQRDPFXuOo8lm8RLvRgja4fsRRAhMUy
DkiA7lWhPCT+7mAGGbPUT/2Llyc8p0eJ5YGy8qVGUFK8tK6NVWlmgQ+sk4tIWZPQ
xmHzRT/WYEyHibkv8daDL3u5E5XeWDcabXtofHQ23pFoLZ7NQo9mUvhbs7wokGiJ
X7FnB2aYRhXAJFgBA+b9O1Bjys+PUtzQRZdzH3RJY9oVaocYhm5JEahj7iMPgsYM
43XYNLM2jQ26CqFmUS7wMdQSiiPe/5iC1emqAP3P0r2TRftIg8BURdhGUYQn1kO/
OLU68WuhrqQLM5acQzSuwi1SrcUyGCDvhizcgg1O6447DH7IA6QtJu7RV4X8VLcn
67IAFgVoclDv4Bxg8OXfd1lZuhyXqgbVWUmlxxBZuh+MFHyJBFJsiO/J1leiOoWV
Y1aXTrD7424HupqynYFosgxrnD4y8VrQi07Uh6+a9luYInww8IqDcZ1Up6ADWKE0
7YOXHq+uxa3j3V0hJ+/k3dSNoJzIG1p8jGfRl6X8LBg=
`protect END_PROTECTED
