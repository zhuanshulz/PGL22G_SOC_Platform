`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Psc+pmVJ13ry5LXONGPw5BTkvqVUzcZ58J2P76Mrhh13S71hD14uzj6H4ALAJhKO
CqPYDIsc/dOny0J6EYmM9us0ceUkN6uYXVj1muD4s5HYZKR21qZxlxCfVUUOsP0F
DX7j3e6ZmY7fCmAOdNAwsNEXJxXexRAB9TZv1M0uITDdGxk20ix2ePFjTf/uNWBF
ysFsCaUjGaN3cVSGcTmSYvqUqUX/bgbkIJVEcjlLpaWFFatgzvUa4sKUvdysBlnx
9EILlpg7zu5uNEyKuSs0wpIzU0RXDSlk5ZpstB3Zw4WQEhpH4oVj+3ylKOiWPTBn
GMPIijWLRoQl4Nchlfeg6U/eTUyrvte8QdcfpmOI4gvG1NhM7eLnqHB/R0ZMIl4S
z/F4ifABbUvnuYRTbZ5K2iTjC6bdVWySDxaO2IC3QVXO8jFILZvFu463WoN3BgJ4
M5HUPNR1WVk3Jf9HTTtaPCQB5b1/iRbWVtraFNvzwMJVRwW3q+7PPhTy4CNiN9Ld
AwRVsSE4zEiZofPB1Rm2d8AiJodHkC/pxt1HyI/UiSBMvHt4BINyzf3GSsfZViWv
LBXOCXhTzkjMaks1iVgwAt/GSWHk/nHcX7ZDhPiiBQeScpRJFfrKKJI9fhVxjqEi
4j410Ujttszxn12t4SBCxZy8Q4Y88FgrV7OP52dJjJdEAsbrYbC7J7wiRqiKSnTx
C4DTHpjKUJhYqFmACy7nn6OAUpxMdztBhOu+KEKW1QGc7c1V/zo/aKy3rpt08fuU
OnUeKIT1XnXEvuCs2/GwKovRkhnaH0JHMRkEirdEFKnatx5bX9YtgFUZR97pOyvR
mU6QLwIhPM3lA/XLG8I78Cl2D9EZNMOCdw3US3bCM5nsr99e8WBSM5k+uazGYnx/
xRbCTZnN/cNiln00Bui22reePSFcoFc9SSBBibNuySaeN7CZw9VJgElE1TYlpoGk
uGgyEv0JwaNo1o2LDpgLaeUuCWOM06NCbyC1Mib9mCGXxD87FCgoUPZ3ql5PwLYF
Gi0EvyMfH/Pj+UvJ1SDbU05SUyf1C7GXltngAorKRsmGUXIHgEJw99/DpONh4qPC
TTo8mJT/8miP14QOmz7OTuGvFNHAN2pZFOFjhsPSfyF2AdSR/yyNSNbgxS5SBWjG
BzGZpcIE1nMjrquVPEBb0FlGW07MKy63C6IGor4oc5hkbLzTHdBRbeFZ62wdx0/k
DuBXrXlDfu5ZRZI2VgOF8iAV2r0TrnjwhfLpj9QKnTO809jBAADNvjSGRcNlIrD5
eqx6gk5xJ/f4d1ZrpLbHbXEQuPRjyNMzLEOFcVKL2VYvB3bLpZDNVXl99Vwpna4m
hMqhEQfDK/8Lo2H8L8bitktu/qmZ+YEWJL0OK8IA/pIN0QiK6sXDzurVx/SH1/Hb
Dj0XlYSodA969P3RnQe4GylrE2xbER2RPPF9NTcMG4xpSZFCFjen5Ee2rSZiRTBJ
S+Fc05rQb7yym8HWJ99bc/GnRV6CtiW7FN/7UXj81zo3ISspvUOIeDDKl5iYNPpl
86538Chxy7k818dx8aeYgdDLr81I05eSShoa5idIh2dqHkIBQQTpvAZbujtHWLTn
1e4IL2qtOZdYya+Y/AhLq36GPm3+2IotGo/hCTA1VOpInfKJQXR/q4VsTyqW/2NT
RE7M4Pvl8jecMakNvQSAj95WWD0kSr4CfTu6kXF7NOwXGqSMx1NvKns+KfI7Rbx8
1kAFCZ4TxSPaHdbrA4Uod/uzGz/2aayt+HYchFsinWKRf1U3ueNZjptx8+m58OyL
RIpY/QpRxbAEiyuih+Dnum70atap+9pBB5mCwagm5mzEKwG8thehAGr5YiQxSc48
MkkFGQw9irefu1XHLDu6ot/AnmFnGY5CCta9azDxXX/0LS/d+k3FDcz2SU3YMenn
ozlJiIYm7tE6gPcSm9Lodjn9ni+Vws6BPO1b6+uBESX3gZQYWlMIRtiuOzE+X9Ce
Gdz6SxsQMs4PQZmmJyJsx+tgHYBexE17rbsXq1uf24iq/uE84R9rRo1xlJ1adU1e
b6UAmBqIGzKhbDCpp64GqtRNJ/IJZNShsiZUsyVwxZZECmLYYlHldOH8ttA615z+
sraFEmwm2AvBbdKOTQwYOzwNeYFbHCa2MFAPljRzFTe8Vs3w6/gOtv43tz0K1jyH
cU5QxNK2DA7bpVfcl8uS7b/gaiOhCB8haymdddGZbo/tYU5U+WoB6GhaXAs9CL2n
y6012iHjqYmaOEZ+2p8LapyCr+e3F3zSYmvW0LtBnv5IhXvOwaYiz/8uGCaUyepY
VNTBwetUKekNQEZ6IwTMa5zB4Y+lttjZ2CmNSNJnOzOJCIlihaIo4gCD2mP86V4h
RbFZvoUwpnAVQJqQrD7AsjN18im3qX2QdsaTfGwR5lJBsE/rn2As6wRPInJIRtsl
tDugTRRzR+qIPsiCrO0CjPc58X7BC3R9ZXZmaCF+8j3shm/upG/wl0rgUKy/ZUwy
BYRRUs0MjOQYvnRTccmEGZc7FWHLfXjZ4TEbgU8lscfsnpNKg+y6pNtrMoD+1UVP
RS5z9DabuOtYP8L1F8kW79PlhjCvULh944JZb8q27F+2TwKbc36EkTYpdSBiayfr
L3orTgqpZ2tiSTRARo03jXHA7C69wTGjussoWR2jz9amhzmt8dso88CecF2qCwtD
OZ1ke9DjFJtALZmEetuZfwHeLt3xsaZGtWBOh5x05qNtP5WhXa4E3UnH4xeAAe0e
AZbbJ3bTRN59mAJvaTsaUTATnml+ZVxf1i0f/0JEAXcn9lTS90l40lCNpboyCfpA
agKOw7Hs0xh59BeMewlQST9Pptr9J5a3Cma6mkPTU3297Rx5Anp/1F4GhYWxG8BA
uzVDAUfIC+/esKa+Bq66Ca1Y4wH1KRcBDQUaAIyu8Y5BkOtVOKmSVO6eBVk2tJee
62re40D8MuRQL5OCyzu6qVs3HPd/DEL7YAoYFRT7WCwgbTLdMy9ezjx4Fgxbdwzx
drkwSFg55lCt9yANjPmcY0XR+SmOpuSAYGJEZG/n5sfLOu7+YjgPnjt63UJnYF8e
6kUyiPBOlSYT9OBIjtvysFNnQdkCJZ623/wZ4UsVpvvdRwd3oW+B70NkhUc/GVMq
SOCcfsLyaL/QYduIHKzLLzQl2qxiQ7fHdPrjBtGcmak8QkvSC75g1/t/6O3pd84e
4DbVFv/MrBWN12qhLPTdaActrpXCqI+sSEanvIlqUvmLcRxlbp3ZxSxY60H4SsrE
ML5S6PZ7KxrQhdnMu0g9U1IVyemxFH4B1QpwqnGzrsd7+R9A/TjQJUM4c0sSuTZW
5BPQtnflQvlSzw8ULacRVoKu5XDb30vQHR5w+3FnSJ5KJLSa2g+Nmmty3y5i08JN
DXPn4yb3D9JCEECxQuR8WTdKdtxtHKJpfHpV+YlCZ0xMmv/FSP3Ykl2pRc0T42FA
/S5kCrGdXIXbQnik9YEtr7OHkHsHSf8w5bNsvqUkXsW3wlFEfHZTnb0le2328yXi
QoGYFC0evlnlgj/yR4wy2KU1zNIfVfFnchiyPhgEhpy8QA5WI25xXHiHU+ycbuAO
3ExleGf0eEJzq3epJmvi2SwJxCwdEOW3VN+dpnsYjeKMlQ8Keznt6dH/W8Bj78cg
Gun6WJu0PVsnKRznCIddAx87/VJuNxIX1+NZ8nwvPbyOok1learMpz5dhotdBHKP
VzqacoMMFSwTK/14LGW6Rm/ad5TSiX5l4Gylhm7yi9cznqm6IGCcCzud0z1QSX1I
7kgdRxSW6rMuuPuqJS9fMg+7LnDjnUtlx9iYH8uZRahf4+stUZp5n7dngc2CKW0H
cYOf3lIJpAD+t+3C6Iz46RNxqY30UE1C08dIkblPiGePJqmxZkoEc/ce+XAZs+IR
TnkqOwldEyIHGgvySSpzeFRkXIjjzpEh+unJbGEO4thfgd6RA17ZwkJG8wbpWBXt
T6PUxvgxSiY6FM7hHvyJBrJgqZ+TUYWZs7vyNLV5dOcgwCCm25NcgF5jDz8gJx8G
iBlneufqSkHQG1JvpN62PagTn2EQ0+LlaZjW14tWrCxBUclTFoWoT11wfGLY89No
EumpBJiNrRb9f8uTAHCJWeh57x9usjFfseIa41TlkkUgoJ4u3XE1HnaHZ2HA6PR7
iq4/nJlC9nd/UZvJt30WkYaTkLXMOFTqPHUQDA4b0/f686WijVpj7Dl0eNHHRweo
1LY4e16Fb0gOADVvLIOze8ILMvX4oky8dhMNXxDzQTPxDYGmUj9d4Ecg1g5utWwl
HeGwj/FjilxM5ArypW2E2x65hoT5hXYisTutCQdtkt8S06qwHKikuhe7QsuXsELs
qLBkOseiYjzsBQevX9HQ6h6jLZOa+tBz++PWuO8KWiXyKzDSgPcEuRYWLq05w4uT
lLvhyQiKNVf5mhGSn45umgkn+eHBdtxLhEIY4nRUVT0CcXS/6PmQaU23vA/qf1zl
HLvBtkEL+3lhKxq0eSSHw5kgg4cBZgUPHRKH3e8nYsD4XHua1OK2oHZlpX+oC7QS
3E5l+jdyQ9fKEutFgPNk/cSwuoKAY6NnVPI9QJZSw7cm8oOsBA4/e/wiD/rAyUe4
CemzOeuE7CgKRWT/4uVuIdItov8KaGEmydvEPzWhahXXc9t3r4o5KrYbBpGrepu3
0J5iTZx1I430vKsCjRZWIcRqnGpWCrBE1m5TZX8vlkQQqMEtw+sPwbXmSwbNDPvB
DrjkFpRZoHKeaAsHMIfUkBAHh+jKbSKMkHN7VMJe2AIaN/4u5sg5V4cpioHsDSLC
MNBdoCg0J9H7Q4bJHkR8pInmwomppFL+qGXhH8CSBYM165prndr+RDmvJ56Gcbob
heiBWgC3E2PkLoPrvMvWvVbCD62bmWnULkXva3zsXGk4pQC+Ar1itLWEm8LXM11b
+Kpkvd4odw1WEJ2f4O34/TWlu3S2Ot3OzDA08kvTEpwXhwl9ncF5AQaXYBG6lp3s
lIWnR5Da2GoD3Plc/wDWcwPVruXB90bSE0oZSZl8ugn538jvokuLSEqdX1rM816M
kW1nYLfsf6vBqeLMdaLEcy4oV2viqT2sqnJg6WHXfI2zDLinPte7ftGIbaa0virD
WI6A4NGyuUOwTiehOlqsVeiLESWVI1LLfleuH9qN9RRMXm6Op4YCT9V5vmUtMhrL
cxPHJFpr7N8xMxYW2pE4B4WYHLmhGXms6hRR4vZfXbBE/i8wOsul3ZZqmZN/AhnJ
Gmai5KfKIZ4W7RXrzWan7Q==
`protect END_PROTECTED
