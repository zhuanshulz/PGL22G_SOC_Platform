`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zj2bgbIlhIYpp61YZuXXFv82TISCCCPWgYkEEUHXaLMp3GkJ9hpl/+jYvFVrh8H9
LGzKkEq3R3h235ICiS25ZLO8Q+IIZwCdJOq3g2cQVVS+RwDauy+Q3li7vyXAJIUU
GEC77WQYJmxN2tyidbJcJT6MWOR5eqLKmQPBP3W9z2vuVTPNcppm2eV2nn1e+rFH
QQRgb7XxhgtyJ6cryl2OFz1vy690oiNzQrMMPBSarwz2p12J/2bdygO2muZL8Jm/
0SqOHeQhiDlWk59ghyPRuPX+kvouxumkt+sFWzrqEl0iStp9tf+mdy9pVW5nqOBO
jkMT25x4GO2RrbvzLHUpcw1wZkFr5ncoz4uavmcOL+vBxjkMoMqX9rDHK94xvJSr
Gpg/QgjFKQvISVlx9dnYpTnvg8JsvObQ2TO1+7+inTugdXQcCfyzdFpBxOasna74
owa73f0SG/nOfgwtQVWyIEk+mc6vEvRIstuUFzNqnQ+S2ZWmQynhBNmbNd8nWS1c
UH0sk9AevmN0NuxRxMrPYopx/M0FRkelHTNFZwfkfKRzw9FMFdvdprziZo+bOXsd
`protect END_PROTECTED
