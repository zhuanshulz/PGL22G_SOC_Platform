`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OKSx+1DIKJsxWGEsVuSCAEZSlc+JoLH06w0COHY3hWLAl2ZnPH8CxhE5EYI4Bkcs
iNBfF+omOciTZBEutlbDRMk9kjF/6P6WTSHOwr+Vbs/nHEVASfUOEqdyz+Ig/rx3
kO0fGABeMd3+z4vxzcdI9LOrTs8G2wj038gkWDvV5tKjzHXipB9Vnj5XC7//VbKW
/3e3tL3fiz31chXGH+uFEaLgJKn9ExIV3Vt/yHX6eAsaH2rZMwuSe32BM3CH9brG
qFsKHX1vys6RoP+mWX5haBJrZm1ug8oX0T7e9yN1kqT92063NKpKKgzLK+p/iCdl
MyEcqvvQLDqf0eVTgMzhar2o0EpG7lWkpYH0ashMcn80drfJrJkXfFvkLQqN2rC/
I7TZVGZWMCGhniE+PyIHjAGG6UXSjCT04fnoReKiTIBUUFtIL9JtVa36sbt4t2j7
4VJwQexvadVT2T9QIEzt0arv8CXb1WJmltsHda2o6axLwFU5QcawEEddRYWbcker
5Eh7943zjS4Jt8AFgIsFTKA77DJuTYgAwdQomFOn4uhT6W8f1bG6SqyC7Fj42bn7
QOYed10ivafJTY/pVNHVsQ==
`protect END_PROTECTED
