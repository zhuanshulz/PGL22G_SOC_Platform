`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PpqVn2Px39ZVZ4/1wlS8Cn2MvMhckiVGp3azsSUmrViItwMRau1HvHopTJrAmMRZ
/3UunC84NzZk6U9+aubpJbFU77RmeAFJ+BHJUuGy52BXTWZ/qJDb+lr/5v+BnaAa
K4nARVvPnKEUFDX9cnH3IZBLyB6LpTFQhlEg3U450e16nZNH7mhaxWX9L6DgR/GO
0gvl/K2At/tb0Me6dtTxyirUjaTyC4P8pus2LRPef9c0Kvgrqn/uoBI3aehk8myj
LQzt1sFjaHU0XZDxUiTel03P3yPcWdmo1ItGu1AVexCeO0yx9Rf3Y5SswCUqZU2u
ejdRPGwSqI1YNK5m/JosH3L5QKuVQjCuhMa/9a7aP8tSXVbddrwr4IqSvnMhzS4F
LV6by3J/ImKawp39fq82rThV6avYPuQVDpuyvDWRDPF+f0BQmkHqyCTr87ENj0Za
94nHXA0i8YGEkYkla7LhdPJmXbwKplgDWdre7O7NR8jE0VPKtMHgR/2Ubjh4h7+o
XqJUDdzDcn9QQAf9cmmQUnuou/l5pkuQUzT1L7bkxMQ4TawyTrnbeXRtz1y8bD2z
LQlvO7GOoRfgsU/OX5XU2sl3RzAVFKo3Xc5jsrOiVKCTmGWoF6RO8wjvxM1a43KS
mP4u9Oerx03Jx+SWpVyHTd2tC5mnL0tyJGtiPkikolI57fXpvzyxDZvaltDmxjHw
53CbZG2n4ZQqPU/e/S8za/6Hu03CRBZq56WmCOYJ+D6RTKdZDn3Z8BADLR4OPYhQ
8JQ+mkyh0o0faXl6BLhHTZMis6vjxSjQRm19IOEu7YmaW/d/63oPHH5VL8e9Jkoi
IrFLv3GLRuZr7zk5dzbCCRq1Xqfy99ouO3EoxOT3l38LeRTnOSeM8w125atnWJAT
q5o0rLQHTdFzH/EX/0I+eo6+Yt2uFFLijZ4EXGo74yFyPMjXZQnUzLQmaXolfvcE
nKH7rTvC5kAVcVe9n4COfsIcaT30G/JFG39uBfS7GbWZmtpQtSm9gBu9d35OWJFS
mltue/V7E09oAbfThOsxB2r9fqciOpA9H/CFqdlku5RKsOX+k80F5KKC4xSpu7kt
VLLfiVdQuBIgLgYtjJWUpSA8c2NdPZYbHXYIO+eOukQMw9HH4m4yyWPbhj3cIEiF
Q2rAalWx633IzdvYb8HDKOFg2/gmXpgw8yDAvWRUKNnYRY7pVjB9wBVGK//RDR++
3olA6fWqUskQLo7vbAVQnOxuEHC5tR8DlJB5LKgJEtOQm4pHuPl5HdA8+ca8/5WD
Xjrl4ke7fRBpiDXpvkRq1tJmqFlzbg9xFEaP2PbbBi3MM+KL9KWnx3uUt6e5w1Mh
Sx9S6CzlQuDNV8E4cEfbzKvDbCfQtr8etr1/CFTzG++2y2qecdLR5QyszjV2+mD5
WYiP7AgCGWBAhYkftsOqV63cY0ybY61N4THBHnuDyneSs9+7HF34ja4yISX6pF4X
on7dBO6WZy6qv7DfdvAfAtmwYAT9vKOXX9/oKMGVy8Mm63iO42aUQbXgjZdrETnf
NIrnwwM/8V2DJyDQ6xDEtBl1Y3mSqSrup3a6tAw1U1OYMrPO4opP7+mJt9FsS0cs
oTNFvQbnKsbjrUBUn3/UkEoNT4m0jvvs6isFySczL24M/gc9cByrzoF3KaXgcuLb
m9N7UwgT3b6WVANTYT5pOR/qO8qE0KUQQoXgiAkbOPhCnrZhsmLpXkbk0WjGjkk+
fKD34cMylg+k4s/zMM/CJXocRVenQwtZWj7Hl5do0Od6cIQ4byM9LRuxiJoihtb/
uiilpUYXWzIxP6XZI5n6gGiPMfFEwWzLinADVLGo2jkroodHR7GEhsnXsXzBPvdq
j5OnI3tQ2C02iGEGKG/3D3gJBKOqM41Reg4sXoYvFsiVthSfeF1tS3bps8z3k7RI
RK2Dg9j8X5aMH8U37rVH9sgVCBV7c4O5q7qhGzM9SIBk72SfKx9xnBrfMxDaDqAn
xepIDYKk9Je50J7zSSsjfw==
`protect END_PROTECTED
