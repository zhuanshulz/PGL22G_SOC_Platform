`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hDCIWDrNuAoF/j42jUJiOEoiczPiQA7w8/xR/smDL7zHNn6rqCxZB2yLyXZO3r7W
fL5xoxE5I1or1AZ3YQ58TRA4KZNihK+2mn1Jc/dRRJCSlxaYMXCdQWQnI6Z6aPKj
fDqgBerJ6EIl0OivECcJgle1PZgEpzQnHuhvu1pUhBfObbtp9nvcqgA2zbMsqrJx
WjIOZ7i3UImpy/rfStihMgrHYaecjg0Jof8I+7hwW3ALGQV2ZyrlxPFSjsX48yeD
uFm8hrdhzqfF6vg5oQu4e2tOtaW4VekO3h+q9/5mAc/4VPHqgI9YjJBuQUo65KME
DRPWhiL9AjAyozLWNBBP05fGp/stbMHnbVeqg+Dg+tfhUYtn1mxUqa157pDNwc9u
P1qnJqZHsnzsErvBOkyw7PEBm6ML5KaybjfLFDTL28wnSJDud7YpZVz1Q3ohkS4w
hcXZOHYMjPO5py9ajw+7hupl3rifOteYh92IVlPMBETq/0zC55SzdEe7KTiJyk5S
`protect END_PROTECTED
