`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WbnAFL4f6iZAunZQssLP6P+EE2J+1h1XyXFViIO/9gBKIWHTnuW33aF8Np0ptG8+
/3Qflxa0hBw1AUVF9EJOEDEQzQz9o0ZTYbkMrEq/jigODh8P+itA3h/WTL3ljqw2
19q7T/JXw33rGyZpoMFFvfR6McJmFW+JCuqIi+nX+a15yZIW4c0VSXrLREqgNcTM
Bvj0T9qTjRkw+7VNfzm28YqR4xPZ2DNX1+5z5CQXr+WWv3ZPhbAD1Bjs3DFqghPe
A5XkyjMyWfMXBlIYixQ35eMcn2dVLhYoqZOEBGvPjvVliiX5O55bas8a+46bO4qa
qtzpxV1On4J7cTlGkaykvf8X19Q/nGq5IMsXOB4TXVWfrG2nNHw7PSVDOhSBI/Tc
J1drKnJBnbq4uZgXa8qEJpe8Ge1rii4KlYWnD9exBtgGfMsh6d9uspZg5XlSEOsV
wdJ2xuhDvct/Lh+KNF9U6bk3x1dWNz/xzQFnUMN13S2bSkCrqgh0oFgF97fe/jRW
etERybv42dTctGhxQiR95eIZTfDU0PZ8wPilXDKqnCshAEvJZlG25iv6Lvusmjsh
pu0kn1yV+D1tOAwib895zFWW5GpiG+oVaEa9o6plOx3OqN01uduIz20+JOzLj7E7
kMwJz+/+A+P5NkgpVZijRMqahBtBR2VjFfTViSQvEipuJ0WRGucBrjeViSev7t83
5Ef2bS570ROF1IJ23rJVgOK8MZ+TOOOZkmIzdYfiUyF41P2zg/Cp4QjBjI43ftRt
XTpOS7dGh/sjyjGZ1F7KZ1ZJR6cEc/IRUIBswiR/X00dCBhkcyW7QLHu8JfRlfRJ
Bl/avEBSK7/zgT6AWdCqHQH+Pf8wRtq7WT3Dfajt0k4CUOJK6MpKjkAFF1fC0jnO
Z/7ABera569L81Hzh1rmqi+xozzfT70yIm9OC9v3dCLpoCRax1LyahYVJNEh9NmW
+0ycp1o1AL+pCDQIXK7bTc9izfwieAqfDuC9BB72WWvibf2stMbGG4hvFk0X6a+l
WVLHLoU6dri4eZQ/f+AOXeOoEbAPSPeFcxd69jtT3Eny/RyI//o94w9PwOAOkWJJ
DvuGB+P+ujZjfGGJD3vlPISh1TqD0wTH1F2ZgGcKP1qIVL+uuaaBK7hZIktlxz26
cZeHn8uYbw+Z5c90UBNae40Zzv79Nx9awPLsRGZqwspnO/m5UBy/7eusgchCDA8c
xl8SgcTVTtD4KowcXw++kZjHEZYF6Ze2pyil6HhhAlCVnJwbKR9hg4EydQdOdWaI
PZ622AgcgAR0JzMDOm2heJRWGvTjKzoDj75Suc8AXbfD2mVX0AvS4T3mfqJJvCWA
MTGJP3AXyt+a2i92XDCB99tqwHwrJbjqei5ye3+DaXlbPCGeXnAeqrYraSgJpDB6
pulnfXjhotJqmu5EMLVmwr44MRxoKTBWJWXFv2Sl/KAbgGXBhzLnpBQq6TdLnI9H
SNs/a19mwqi5TQNydEh30MUTLX3f0od1V1f95PoaQCIEOII/PaAWdpxw1glku9XS
yEP1fDU3q2e6Rzzb5ssz5abFOvi8x0Nvr9awI0RJxbfPWCBTrPZ+xWVvQAAQkLeL
rWL6h/BdBJeHHmyBygAcYizrKN/41IeEbE/6rr+6o4suOjoORVzWXZgzNo17Z4iv
hccz1mqCPcJJlClvIB87GSTxCjyokFmdI9Toi6c0PkMK+2pWdt/3+36+qMi6G+Ne
HK9xC44IYq9CMwOSk3+kodcAcuaOphry3nx56vzSGOXAiP7/Yu9LE7su0dWIJjKu
VOSk1UJ+iw7g8Hq9j36vBH7frM5MXhchKd3y+jYBFw9xNUHqFcARL6F+Vg2iIrCR
kZNNFRcCJ5xNkxFHyfOYqmZg89toyklac4d21GXBcFHo+64ctizLMzyj3NcqqYmb
RK7Od0vnPZGngyXxlo9qAAMMwb14uDWu0UD9yEQ2R4rO7Q+dpuow8ezrF9FqLzm3
1zAYezgvjvSarqodzwCm93H9Io3KeKlIZUNdmniDinUo6mjhhVn/yboenIZb86RF
7QAXPe+MSEDTav5TyW+EARS/RPJI1gn35rveCgGipziHqNFYB31b+41myQMlsk30
cWzYYcxinAAYcr5ngXEivYQfHabTVt9aJBOHkT2UbHRD7OHMxyIAgM9KFWc2NwWM
Jb0GjEhX3RTqI1mYw6AUJB25y9LmYUlaCtHv7ec+sfUB9gIOXgfIxkFdXTN+qHp9
iQUGhVu2wtu8WDgQ6yp0p+AS0o3Y9+lIkGd1Msa/1AeicyUZVg9ev5ciwYBASHqu
+f2zLoTo34r0RuMhY7PzogSzjOsBvYTGwRpPZORVVhEsa7nCueIZ68LB9siP8FE1
qjuamS4GmkKsZWgQ9HtfEvZVqpHyUcSS2N1xriApnmufxgLLyE3qJokOatX2MZ/f
NrMYnhsTFlyE0yZ7SmDFKgoG6K+/nQmO++N0PwhRD+7fb9XyfU9qw2hlaaVdQRC2
d0pNot++zWM3jYhDhKlhaVHRYf2VWtxy97HbHcEgGuaXiBcDmhcWa2GQSe/lsOv0
5rIJqqf7K68tlKNCdNCCjxHin1yxESeYRZ0/6LBFzStJlB+LugGMdGMVkRXodlAt
jAGU6hnDowd9K8eg6VyCJl3yBbFBGFFm7W4gA9RxJdybtSg5f8VmBrGOPZHnOGru
IwwQLpOFl8vlI2o+NPpIKVJeMP/HzUrcM54hURY1CViszAR5qIaA5R6U2aDAqRdJ
Keh5Buip9EWnkM8W8DnOJcXlWaU2+Z+NOUhBaOS+2M+Xk1LHN65T2hpux20R7KSb
NTuhEFe6MylJj5K2WjeJegWyhrqEJKCM4/V/dcT9Z8REpmPvHxhO1Z2c1hvPPYX1
RGrtnTyUhKNMHAueGHqhdz7WupF8r0Zbe8F4NKHficKx2OOp0N/gtQOl2hagio6S
CPwNOg4vWCSoVuBrNzmnw+24pFs2PdGXu4mCZ93taPsJthNo3656Dk1gGhCIK3EK
zTtDx2tmFJynx+QM8JgMMV1yKnS1Gkz0sWxMF5gz/jTinLH5CXz621GfRVyN98rG
igzkmiOH+pnjram2KLp0IjglJWrAuBBi5eHv58o8Rxkmmuv1bPkKnYfxN2h8dF/P
vLz7sdb/4FJNLEJ4ZdNJJSuSPgHjpQtkGxYYvHjirYzl/vQkjlcQY7ESIRvlZ+dS
8M/5tq/TRNYSmaEjkmdLnjv8L0zxqiE9k5/ytccvUU5aZ/ecWafy6KTkRrt3Xxby
pXgjbVzt62LwY/R5CNVnIysDfok/bRb9skLCYp+Pg008ttXhfBvr8ChpMYbfDfbi
ToUPtGJG1RDUcC7SB4CGZiWmmyDWJ73b9mePQVbupbqorkvIbm7b0vDi4HgxSmCh
ovo9vlBovHaxWJjO0q5aRZOo7UUrqy27uJ4E2WcvegC13s3ogOQhyDiiHcjoXSUr
E3+wAxkeli6rePnYechJBW2LmVQfkJtfrWFP6z4e0aMW6R/WX69p4rU6IdPGZZBH
UBKYunHUyAG493FNlUx6DTggzfuA5QDHYOXBMIMzvPJEu6bIYfw5yXDq2kf6sFvn
IbB0wt0TCEPhIXL54UyHoQl7827PBQbZy9i7dbFA+qNc/00MULq/6aaqB/ii7ah+
W585biJAKTjiOl78FfwHie0aNeuRqc68yhfbi4+uZ5b/LER/66lINkoCAB+9XVhH
MVgxg/6vVk5Q0ipMFRtBJ+4PA6v3tL6zSnKjJ89qQTF3Hk+U1J16mQyffAe/YJ56
WOGXJQhgzUBInkGrLmBWcK7Samltt7l4ZQp4DN51WhtsIbnVx+LsO3d5RWvaUHsg
q1LCq3JIIIBQ/2e4hIk3JGhl7QQDBOFKt4D8wmlhXp4UoMwVVJTzEsxroARvx86f
F2zTZ6uSAwQbn2Tz1Fq/pBBqTmgm/yebojq4+hv+rz0r5IgJqWyWaNhoBG5GmImT
yTa0HGDnzpzJQPWA62zoJ9hlU4x8tHvLOFMRVqsjlcjYPqQsuluTU8+HltYu3KOh
GOqPS8HfDydI61QSaYb9ryIQbDXS8sYN+lkhYLpR9oynATDpagcqq3xFWyxOrPPa
pVH8rzCW0R/j8yyPuXo7rW4SzeJjv+1tP7+palFQy/7cGmSHS1ii+2G+6uyLG44i
ut0+G5+zBXDJ+4l2Zjnv9NdpjOhDAIXOuPNNOKiwDU/kbh9WVVUpGRx6vorbsSzW
L/7A3JVPkvZvWfo68VxteQDm3ZReItBjG1q/2tfGU/xl812cxNnNAuL2Z14Z/8KV
oFIFHSKCSeSvuRPteO6oe3vgR8NLJSOE5enCwT7OXQGDUy4tYSbF2TeqOpt9T3Ck
C84F2yYU6X3m3d8JBSxNZKXQ3+2USCCD4Ug15sgKKtgAmPGkakDHhXpoXQRvklLy
9xFPGzNuBo5XkEG54droS9RCKF6r2T4K0f8Ac9yICjIYDdvEVSrCtalV6llQm/El
eLb7Kl6+xzxBhiI0TvAmurDRT8IN3XZrmPigXEGtAn2GdOm9uIRrvdbVi+1MxNzT
ZXnU3ShHwSQPPEHjeclryk0uiGF8fWf2c4r3CyW0fObnIDdMzVk5SwY6qzdtNNiw
jsoCUZtFa05M1Ugr9sYBsdpi1SsEE8SIzoy5cxVciciK9Vcb4pbsKEhQ+hkVA0Yy
kJDaewrcAk4Hxr+XP7NMe3mPn+FAcSKk43FwXQaGK8CjBvicEnDJZ/fr3eMyQXMF
fI2DHbXGgGFZpv5FgkprYJ9e13+DxSk0LY9J0YJuMhb7yRrF6ut38bsuTe7mft+q
zw5g0bA7v3NIj4AcpQOzI4sLpuVsRMaglQu8zR4wAplG8+P194e/g/DqrHhsuiVS
o1P6gxFsW0dOsck/1cnr0oMpaqIsduQZmWhKuOD79WLgydUCN6/mhCurvK7NAPS+
J5mYzBBWOYGy5B4uA0DefzggrC9AK5NN5uanOQAGDNshOjAyf2Z23ZgyX3SieYa0
MQem3AKL2dl3JOcls6Kp3iA/4rE32ezRtkYas/NtcyCuxgpw0MLUEXbhODExKgrO
UVOe0khcRSwKeLR+cjd0EM4gpwtsWcgHV1XmPm3J9gAdoilnmhuWyrmfVJoT6lsD
BcF2sWBfIPCeLGHmtO7GFLfQGjiPBnALDRY9Arx+MI8c8vKXjW7dYn0NDkdIlnnl
whS9+jZTxn0PMnIsErev86Z02873Tr17Q0QQDj/VZn84QBbIPql/QxzDsnYexw2v
XcL9JFYK8HOQpLxoJ9dFfTwJyq4in3huYHYhwuGgSR5sailXiShizUXR0GLBBLOq
VCJ+cSq4+RRFx637Z4me9gYrSabxVhQY9QK0WIsEUddUoejgMJQMdAWMJJ0joEUz
z+pkukhsu7yxDtb0gA27Xs5UpFhMbUPeAkOA63Jn1lGJosJgSnaNIMfJS2NGYjkb
7gjXMQ34AgagrFfWvP+2pvkN48DFrTpXU8ydaS873zlavbia2AU4OGNYITyE6+NZ
qPVaeEC3hp9QhBZL9jQyjAODmEGUaailv6GBTsKS41ZwirdEvimdb2BrS5vPhEzQ
/d435Hz0b+N5koGSTiWEUKjiQlZKJc3aX/7AHyPEbyreOQ8xwSPPBBJ+se7ID1HL
xS/VRB8jyPgxgZQ7mOrf5PR1V/eZtBAVhdB/oA1uz/HDK2EVEF40ixdyiwqC0EiD
ZxRNlzdJ3iL6Jdn01vmmhI32EzjwB8HTDH1IQ6FQGCGbtfwF9VHw+8xmlkVMQu1G
AQmRlXz4k8KcABLGcvNEqh7Uznrg4EFb1I4l17AZHixbPSwycFKXmGqCaQHJxAB9
qIRowDIM6QvZqoJRPhiFM+eE0G2mpkuExKx/T3ikq1cl8TkRoXPwKM+joJVRL4oI
581G6NK0O3ZPrTVVQb1trmg1s1w/9kVm5uLMtV+qMfA=
`protect END_PROTECTED
