`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bNjXepF4+v6r+K3jgsK6yJaiXiKfZGgm1MBz2Z65bgDeRcAvmzy82HaG+An0Tt4L
j2Mk05zRkdqycmWRX8KTSvuoEuyw8rIVmG1tuoVVuQIUfY+lBoPlI6R60ESOKyvb
mrrSqo+MSObZqczbUEl4wczu8s7hgKgyJWdKlqCMKNGYT9iSM2ykgXbdXk1LIb9O
KtOY4+vDjcDRTS4bY16MFSZM8QlYZzix7uPCpwFgJsUFKClkXnfwnBqDFVjHN7uA
MxqRXy0ulE4R3u12y8bi1zOfHExx2GFDAXObBHJTOEpkcOpE2RuY+dr0nR/l5AWm
hnsXCg9UGkpYSK6lDXWjYPYPDWIpJ+/DrxNTa9t53nIkyRyXqLyVKJ7Xf1Xrl+7Z
FZOeqFcGdy5D51qSiuF+UFWwUX0NFX9+iJtPKWBaX5Z1sJ/cgDy7qUac3ZNmeJhW
phqWczIqiXRt9QlCAxKupDyrKSgHNk+bmYkqNGVQwFYFxVA2XzIcdf4KPjRd7PMy
2rmhmMT5fyLy5SXCPNhogufJRUutpgiMRMFZFq4zF8u2kbhX/wT8tnTbTLDaKzQ2
NCdkWE3s7ACL8k+z6hTeE6YwWB4qTWUMvOdXoEO2/nDBBIrwbqc16/+676dAT39P
SLH2AmoEFTK0veiWkHjY8WYGm9ymoZgrI26Ba0l2Jry/1DobVAQMc/f/X/sA+dY0
ne4GNgwMPdwUqfBMUszwhJ6rpWFNFCns/NaUtCsnBYvO9TdorvK15TlVDSDHGggX
mV8XUdKkuaO6aJh3S9fnEPb70oqsn4bLbDy60NFAYSznGdavHb6Mhr5NwBFY3cU8
3JEZjopaXQ+3gjwEKZ7ZYUF3JJaMmwfAC/pqFKt4yC56edZirxJRs26BJ3ItDEbT
ZdAbc0AAv07R/DSD/bgEu8IlM14NRew33odh9RzrzjAQ+eVgMjM18dDpSEKSRM1C
+xR03zKt3wawFK3p2T9CLSSfpHcvZQeeq3SPMU3AQMlpIjYMa1AvXuea9poPACaN
Sg0joAxdclgrKGocM9Ry19jdacREwAWFw4s+n9kFfUsqRLPgT3jUBKSKLSo3KEoK
8I4mbcbrhS/nSQOpgA8isbI57DNyorPv6+2A9AdMX9H9/xoiRYu0YnxnnY5LEKRy
txQucRSK40xtMczGn/ZHSlaP+InOpWlPQVQdr7CcBHVLmN6m2qGHhzoxF5LrM4ZJ
pJDauMexxnBJcA7o0gmrdZUWCh2aLN2Wz1uNaYdZMTeszxg9YSaGM0btvpqs1u81
8Skcm8nqCHsCRH2cz/4zgR/kXq3Lf1xCCp0xVifFcO4AaeuoTcMSs82K/NSFZ91k
EhCFxMYVELV2wS0zs8BqEZUH9PD2nQCboT0i7kYbn3DRUDhv7vN515Imi8gsrr3f
VHfSMnS7Zig79qH+63dcIPFONdl6dnndhQK8AxOer+vJ1JvtEU5DcmY0WBYAgTjZ
//LTpjpsux0ddmLy8oupkqCevPcLARhoeJxUlZqW77wLOLZlUqMGDicGpkt5Cmfc
C7m+OilbVfiA9OMVFPMESfchF78fFpedECdYauop9VQ2weJCgsvFJUiegNPzYHCH
h/IZXKOYLI7PT8+k82xZbYEWjJADR+x8jXDy2J95neAQDNu1K87r90vE/I8uOaba
1lx51pRpMVuecchLGRHNmiEhMpv58Lk2R3TQreOW/rSJDTLrouFcKBkY3HIFbWSe
Z3WGHFigMoDxynhBtEz6YDrGerXyQHJJawSLcg/sMrKyiuci2DVpiL/WYMlwV9R6
DBbWSswxJf5k54TW4q52svHoBvHDw7e3GjnFFTXI3m6X+vxqdXOltnHSEV5e7x+n
kgHi9OyG6vECPdLcbiTPD6j5eLkBejH50+XmBTM+tCPUj97JYoSxbWGisYFP0QM0
Ini8ESfnep09IlO0SIs9F4/+RhadX7Ngr7cE7TjKG+8uwqi5HXIUVQJdaJ8fUwO9
jcFdzhgzCCv2kbg17DZR8Ini9560KTfMAy6rQFb+lOFbQrDlvAhu29pLeczzEyP+
ce59Ru+87TMP97O1IBi4ozHbm138RZkLKzEc37TFICn/8SdElLfFM/4Gg118YMVm
iQ9wqRinS7fxuWozuEH3QtsS9ptkjdENFEUQMReRnS5a/yJ4AlIfe8qbk+Xmjh1b
2UTE2LzHpPyrJY7K9432GPlI64c4BfUs2z+FH1TxebL87C3y+6I8MhgnlOWVWTRt
L/Z3luim7B9XiLNT3Oel6m6IOUtGtFp40zJckXuiV0uTvTGcCPPgoC/+IMRK8+Zq
bVLAdv1i81tGrYBRr/ZSys9GABzox6qNRh8ccl0eJfAuNdq5ggFeMzXmvrV5hcFo
ysF83P2tDB4PsV2JFAVrtnvuR8PP6n6pwx0TC2k2ML1xFziIg2iEORFeA7+d1chY
FRMM3BKmTwlGD2xfrSqlgLUtyl//ZlzkV8hJPlZ2iSL8J0ZyL8IvHRjf7W9UDA5x
V2Q4gakaMNs4CSYk2L2zcRmdrP/1ftOKSFx0Hb6AKak1Yh5HR1WrAiQFjdKCBWkE
n6OrEzZmwzpN/kNAHWlR/E0eJAqGk2sOtwNS3PFVaV9zXsZy9n3KB0hMney64siO
ophE46ftPewlfGhxx7xYhmCAQl4XbdtJDUzA0AVNC4K3i27zaktOKQkW2vmjKtro
1Sx4TxiAuKH81xe6NMOyD2bKvI4NZXfXJFdRMlE/fzlnmsPW1FHTg+IYjELjS97Z
Hl+uqSXeKA2postnN4lE+a+O+T7o35l9odYrHZ4NEFeJOaSluMmhaksuSp4A8UwK
W3AndTAqQ81nusn0k3l8Z59pwRoRltuL3hLFPX48XKau89jP3y4rLhLLZjTiPdOy
A8mfYdVhpD+dfd/PiIXeSTGTxlI9rsyQUsOsAIyeXeMpfxj3nDXbgDc7xcqnHrjY
B7oZBwMALvO7S4elpz26zC62JJtSxPlmyWoJIyVxY5o5v0OeeMxrNrANBSjTUR4o
QJxlc34v7NRWjeYsSQntzzY4wLi+E9UAxqr9Qj+kV6aUViNPqfGTjesrbgNTKPSM
G4UHBbL/XQoEQOTHMb7zkN4O52KQuSdBNzFtSmMMn9IHtwBVQFUaXrBx/Xv5i8oT
Gqy9JPqILQjaIMopF6LoBU/XLN48gFEf965uPNyyzgGj1E2IwStUF1n7v5SfDKdS
PpvbxY0ECcJl8GLcUFjaAfzvYeJgEg32QS8DzJKXxgjRhwPjXwvNA6uV4+uNZW0l
eJWCzXwck2nFeqL9UblLjmLWgcI9EFN9nWNJPX5xR8M49WC4wnke3HQSqOeVDwwG
U/O9uTp4SQ+HUcAoieebEVobwYWYOUVuvLEQv6Zp9gZITHoca6Q905KF5m2N9KSk
hbm7MZxbBpoqKP5mzKaur24mbEgmwjFAeo909TB2rh2nVeQ2OB+TtHz3ztJ3JMHC
rn8mC0dmlk9UReXJ0KgSitC2Q1iCLiaJpFU8S4aVtkvcg9pjbXT+jCvICIWcNm91
FrcEv+4IDKAT0Wx8o1zIaKjE2oZ2gLHWYY0naM6QyrdupUMbOtIAB3Feo/2xBl5v
aIvhN3ui6ugvdggfqop1veegluNKYe0FliJt4CSisRYc0quUAhgH/kzhb4AzDZKt
xPwm4hFo8Tw71rWVx7vFabWAclPl6sHBchhWRXpuUQauG+I273rpS/kmu8dRrg2n
z4GsHr66FMORW3XNCawXBm69gmkU7q2hvOIVd5yWhCfwvnPFNFr+IMsdjbhk+t1L
TCrvTKsb6wXVFjslvPCfHw0uC4crXJpiyRHFiiLbFi4I/Imlyhsb8MekIENeRoKJ
WhDuM+srka/TQOz+N38mhhDdvxlT3sYBwW2bdS2+XdFLrKv/x4mmMPjT5vZVs31g
G2qVO+vYnaj75UqG3/QgCV257cd3SoIo1k3Qc/DVC3ebRF647g65HQ0ZJIH0eZr+
aJuePW4BhtfC72wPnaD6s7ohCaXtSHVhy7d57Rf8YHHJw6iNjOXJ4y3T09oMwTdP
nhYqs4z3H7kNnywzjsib28mlf0dZSrkQfK7hv+qNL3ICID45xFOMCzHqADNzS+Ps
OdJEz1do7FMG7icVqOuRxLPS3JS2cYIHEhcQjJkDkQgMzaL1MyljHjxhQKku0tlT
SSud3wZHdFu/u9ro+xEuZ6Egnz5YDvad1mlo15mD5KAfmFRvObbmPIVuDPBzeZrw
uwllK0H3SssH9wkjh/fan7GRNok3ZAABGfAgyO8NnZrclNvc7GFzSeYUoNvNaXe3
7witl+6VEBJDHoUxomqd0onrGEUfVcscX/rx31ci0wXnJI8Fdg8SpljWUZgVF64B
HcEpTwQ5XUCl09mcxgrIz5ze+j132miHX/guh5vspZmIYdsPzdFldKX42dCxQ6nY
`protect END_PROTECTED
