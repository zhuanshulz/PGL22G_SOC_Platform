`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
URDsZHH4zZGrQ0VK3Bgd73o390w7Hs0pOmSK4XENF0A5G3YwsqKuFYBHQnBQvDuL
RXuXCrcdhPxD5jlDyoTi+aCtL7aLh/MrQfyMgzcu8nelEBIx02QBPTPWGTdqSc9t
smSKkNyWeeuzMdPWHOuQfDvMmsihFeW9dY/s2rMlQjN6itC3x0dBvEWQbBK6os1Y
EWST0GRglXlVb1shLb8K2tQe7eF/JTJgKNrABE0rq/hyctl0lpDCZbIoB7ob0f4q
KNPsPrN+qwbSnCJ4+NLF1qBrg6C4pz6mOptNItc6docsRjm9zSVxbWeaXPW4ZhC4
cOvGr+NK3vWQlhJztYIW4KQj5k2KfBrCe2fqVn6GUy1/zRbezyjDyzaeITP4Bmk7
dzEOQFwRJ9lcMg9N7lVXE2LaN/dzB1jFU7Q6c1QrCUFSNG7y7oXwCiuOl8Kc6KXc
RlaKtPJ1bCXn6sL0Yi+YkqKor+iwlUKqL/A+VH5fNAjHVl0pypibSOIMgTK0Lrqp
zdpKPi92aIt6ulMrFHJnHrJgiRrMo6GDmoww6GvlMSP6fgdh/ugiyH1GvzxxYHD4
gPoTlBxTSG+vREzwTS00ui8+XEmk/X/wA2sACaLir7HFtbLHzHNq3+QMld4K8zMZ
iiseeoFnPJ8DDv1zX8Ox6Krods1xmOYEOVG0pPkn01zxi8x7pHvtE6CA2KrYEdpn
Ls6KiwnsRWBFLe32dtsNWUuoUxs/FQb+H0QX+SUBYv/U+6W88ruYhv5sClTvFFcX
/Ad3ZlUGp4EvKaly0LHb8Za7pAhcJKPEOHmAGRfxtNX9A11YTVnXB8I4jooR6yUa
`protect END_PROTECTED
