`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8qMpGALWRnuMxqW/Av4UFRkZ3o9MVPlHKCWCiapuYGHbPlNJH211tzTciGWMkBMZ
6yz2cv8JPRByjDST4yKB2O0Ts3ts+PJZ1a+hoXSa7jIgnkECVRTfL7Zgp26m8oAP
Phubn5nfA3iYF7fwVfXb7Bl8WzRxiCaddIupdMlDicpZe/Xa5KeTtZTPF0NJaOh9
zDANMQUwZTCuZ2SFqCHICwda7tlKkx7F8Uos46DTi6Dz6NyXc4P2uQiT9nu7A3k0
L0ajDA+vBvENctxjntLrYI+0T5Mx0lTUeGbn5j3Zyj+zKXtu6XL2AMevN8lU9cJh
2euhARzyYyO4Q2YJtD8FFNyhjlfC4alDYz9aGKLWFiy8pjj9XSUo7C7zDEwC7Vrb
Wn6U+PZyPMKWIn24olFyEczHD1RtrYj/2tbAbbgqWsTGPDoS3yFQKw4tU5dtLlFt
DiLEltXABPLsuX+CaJhK9g==
`protect END_PROTECTED
