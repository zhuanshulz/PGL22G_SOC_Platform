`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l5CtG7SnL8Ed821bVGekIbciG44naEKMKRlnkcPquRPwm2zTztbF82bIhK6NLXrZ
AS8FbdYAANkxjqoNERB3VjtFS3T6cL1SEcbcY3hswc8zPUPUlplA5ALe8rsZ8WII
iQChbw0uenBTJ7coCY/zsLUAyUAgF+GmD6FKt6pDWdpyyfwEU1T6GUQx79O2lbej
AxUz79OpfZX4uS9sATGYLxlg68ASM4MnCOCnniRSRGUHhv069MRn5P3e0+i/mCC/
wgkjJ3Hp2rPnc/ZRDCbLviYnlateVIlrizXLWI49x5PoaBnO1+Tm63tCngiOYqqs
X2xrAnsbFkmPNhnO3o41hH176p/rhrbJUpHVSiDttA3NDDB/c0YtLLLfmwo/7vrQ
yRmHRe/XoyA0FGGQ5PdGVeUsdJj/zUruNNiDtiDL9aRq62rqzHHMa+7DGmewU87m
q8OyDviJW4Dr4RSAdOvPX4EPCFRrfoO2UHiMXIvseqli8vYgLj6I5FAVr5eoIca6
o8Z+KFwpWZYHhBGBTcLXHaqFegHL/9jNfWyQLsXblCGLpe7rgExsdGojNFvBCt4m
pY8HA7TOaICeeExXEO+CPRHzvG79SeLZEB4K1ADktEWwSzTXEYFZ0+eHiJ1HiN8z
yYOJkyntFW/PJ63KKH4RMS8eena19yzi4Gx1mRhsVjZt04Oot0MMuSad2Sv2yM/Q
P151p561lLSQiIGQHVGLwbossQMKXflUCiM/hFb0gKzvaJ0bnskYhkX7EGG9aXTh
Zi5MLmeOqQe4z/D+ZqADwzXopf6hPcOc0nqqwclVc3QTFUWQapRE7KGYm7mKn5QW
ysn9ddoOF9+a0WYHCITapJCDK8hh+aFn8CRLtzGc/oAk/Lh+v4iJbF6RbPORbCDP
rq3Bkq+eMBNsMGxveLe3h2okaf1a8tcBAcjvRkkUAj6jn1p20wT7I8fo4OckeZ5W
7QY23VCb3RNWg2qWIVZeQBbHoEQ9X7lHEEAHW8rIIR9sZRydpiFF0m9fMfGJkGEo
2HHUsGOhOIolLERlyWWwh70KnF/YIqKokFh3cuh8KCr2wrn40L5KExq8trWDYUJu
FXleLdS+G5D5U1OXqu+RYa0cf15DQn0Lt57wd7yr8f1WX8WGjAWKPsA3gvtZYiVM
JjHl6Nuy6Ea7KsTdkVP9ll7YEbK2VIpw4VrQxexIMmGUdTfJsHWhttMixi0rWDjg
lwMvvPK3CLwblkVIynMe0HYAE+KkkmiJOmydGupTQf44K6QhEwbG9q0zHKvvkwtE
/u4A1QuPr/jYvz0ohJuwW2Bnb29fPLm4yd2oXFcaC+dCBfyHFe85G/mLa1MawDqu
cQmhZa3FsH2Ll8Ti9cFTVrG/2nKCxVBG44iXju3nix9j1UqB50MLv3gVf2HXigbq
7CCB3FsqgG/igxDuz7JowD5vrx4PrtsDNwpRdsqUXGh2OCVwfmidlsf2FkxYdeGs
BxAREgN4O0u4WCrtBSGPoOsWvl7E7A7djuQmKUu7pPRZ81E+GjR1eKDemC5w1piL
kNU+zcY4e19NphezmWVlHFb88CYsi3ihPS6QXqlrGZBHyQHzdEL9qdBtj543xqLc
F3bkTGMf2Q0UByTJ3segVyQ8tRqYTGwBD3eSRle2LwarbY1VcRbLGK0mzZOn1+HF
ztPW6c2rDJG21UTqtPildnZcGh7mQPaMVr7fWiLCisnNEdJ38+pfhQSH++z3STbb
N+LXnIH9zr+ih5FK7Lsy9HxLw5ZCuyF+FWi9NbVkBUtFcmowZopPmdJPGY44vZi6
74PdXulNXNqE6LHaThBLgmZjLmoq1XlxvGpGCX4EO7r6bV1Bjf5Ra0MpNxXMODzS
aM+Vk+0i6icykazGTluBpiEr/oVmD41PATxZO/nxmiBWc1TLUC4OQQZ8GDYJ+Uxm
D6eU8livWKKDK2W5RGFuFonctVm+G+vk2Cv02dVACjkBBVc9U29QflY/PgMHyZAT
aFEaUclCGY/FKD50sRt8dn2yR34WYSE5uV/GOPvLZF+vFC8BQLTxq++Z6aQrpgcw
hzNlpmM6YYZFKOd2nGbDJjkKCJPgyaYFZ/Dyt9K4PpQIBZnHkO8tQ6QBUilP5PE+
kRg/LvOd8Rkzka/jDah4ooXV/rHY2URLzfcAayzFP0v33uus44tvxXniY5PhVaef
L4C8lrXfGhKLwyyTz7fMZgJ3VF1cUhyXh3QX0tncrpX3bUKvuEUvF0x8TLfpMkpl
sPp708aeCIeuI/lnGweBAOz4rN4tPyt+wp4aN355ythWSrL3s/I3YB/RMQh2fPmK
d4RyiJR5Y5JVloaaOmuxbOLYJSiD3hsli/YRUNTLyqk9z5Zk/SW0SF3V8QvdhJm1
zKNYEBgOHi20y7UKUP6AwthKZks5U8b3L6l+5CQImXK46tpAv9acu7H+e2tXSBkU
OTVjNL3jw6KkSwC8befTRilfcvQtnz0Qxg1t/KpQyVH7pkXeymKgCBUzVQ+5y6qK
VpCVZgQIHuJTIpmYZjbSjw==
`protect END_PROTECTED
