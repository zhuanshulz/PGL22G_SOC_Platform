`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0phL+ii+MDqPIES6MlJhO6hu0Hpn2RngBza9Ae63UIKS5u1YlLpLvFsMqwf+3swG
BN7gPwAH6oECiKYJAe7o2wl35uSbYy5lKDHnkIEqzxtFWH/OaWB3eTUSxb+GQdw2
/xe0MputAB38NQg2OB/47HGHm1lEgfsysFXI/ORM3XFOP+f3kSbS1qgs+sFH9v4s
5mhcG+M8eBqo4ncXjaxsXld6uGxzvRArbOmSYLYUBzD9HbuxoD/PiLmQbWChSzvE
eDEMTN9dboBFTidOnQ7nuaXTpD/jwYJzZfxfl7wtR+EGO1lBlwP2/pAkwXyqI6In
RdTbUZ1GBDcsX9jYcEjztg8c76MSjGsq92tzC8I4Hn5cuncej2edweaK8hY6IDFG
SF+pZDF8oGVXYF9Olp97ps4Xqp9VeRaQJYI4Q69OQy8gpI6urw0bjnwQm7mr4qmU
ODS51mMjx54s5MehF5qPswE5/cjgTfMBK3ABuEtaJkyz/ldUXZFiNdoYKBpdSuFX
j/8My5b1VS1SM/tnFf0aHifgOXAk0i6tL+av3BcDQoG9llO+GFhdajL34vL2F0sO
lCjO4pJPlRcDZX/wS6KmycyXlaQvhLbOpUNjWW68ZFi/8vEksBgtKBumgFA0uZZ2
KRrNrL+pbGSbbMa8ciUCCWvu1KiohlYB0OYDp3TssgrxiQ2YuFPDIXyzfDmzkMzy
4+stH2TciiLrBs1KAnf3Y1awDeudXsLUwhi3Q7qft6y+xTh/HGu+9toIcl1v0tUq
rDYJBx2t6FqN9dThcCQq5xpvEX9j4aG+qLAx06RQeWnXfJ1p5+1Dk40Y0HPwt1p1
tNKmd4a4hXoQJlrKK3N/cAEpE0Z9tzl01KcpLVAZS36Ej4Q8/8dU1Kw9OMivpffa
TeA0w52tIUieON7yiErO9d9NH82d9vafBvzq+iy1GtEoOXrTS0EJJWea8zCNRjxt
jk/NvkfxzIfzOWOOFgCbhwQXz95QsaEdD6gy5dMHIezwrIyM9h8tbeJIaU+HWACT
TXm1BNZMEJN2Xsf0yGGt+TVVKXIfykHE6XzP4vNXKDOsm4DDFkBu6CgtKdx7pdHR
yjtx39pS3veucTgad+Yj+b1jEuRWsV5vmGFu1epevoAeaMvvEW72Ujrq86NAWlJL
JSGkFb4pRLK5IIVQ+oWHvTbDrragygk4k+ifF791ONFppTgDQOSu53+dAnEOH3I3
N1+fvFpRcokHP1N4/XLs2lOmmErRPYZ2tV9mJydRG7KGnhZR4CgxOAQWLBw9/e5k
GZpref7K7BMYPoq4quBsfLOcldS4qSq9S/phEc3wCPiJ31GCfiFL0tvz4F4yPkNC
V9l3/7BkWgIFqOex1dY6GqdpXt2huWTdfq8m0yFcZlccpseTQcTG1/PxF8ByJuLn
UbGg1f/qllzz8o+rYQNIXE5peXssVt5ZYIe3WK1R/6gocDW8EHvbjbAjluFdwcfd
Dp8A9YfkngItAqLbWpOHCxDGBGq5XduE+aZBoKJMrSeNJ6TKabJ8udW6ma+5kCcd
i2VX7UsPphXbuhCn7JJ2Y76BhY8ns/OelS/mLaBTeETTKAWywB2Blhlf8Md/Qh1R
jQ99KtIBek9FmtrydnLQ5pb3cOFbuWgtwgTuGXCowFAkWBfgP1/EznpFqS3Pcl6b
G8pu0b0Zm7++hlLYs65trz+wA0WK2IxPn8zmOOFJ23SJR/Jg0KsrGE09n03DgiE3
hxHzuK5MoG1FLOlf5vPFeacae0JAHOgmdr7X/PhXVyI6+Ms9ufLvov09size1yNx
HBto05YsfvEUpMkZFw71vK6Ee5u4cvzklrN7URUlLhR88+L29MT3tKT1xHxJGGpy
S9xYq4GJo2uIdeZ9l6ZkjSugWsPFolAIrZcHFIdauLFkZXdz59PnItrmj404ctGs
ixQdY13vmR1imF3oToiMhNPG7zB94EsLISc4Z6SvKG3ygl/9iMLtNV9UKcSp3MJL
2HasNGl33F6SHIzTPn57MC1MV4MwUeyBH5YnkN0GUq5WzAXijQ5bTaAvyzimCAqj
ZZZpSiPh0IHlgQwwFNpiRG1qPoLnEXOKSz60Zp4I70G97pQQezvq+IO2jEmi747H
bhsfM2FnCqDbcnHCoGD6NNyevNSXxncj40NnhW8N9jPSv2Q6mvZkr/+sSeKR8P2g
ABRfJeCoo+O+T+HZYHHRHIc2EdXJbTcr4yLsXe25tGpGjh1Di3h/YrZJlXEZ7eni
btMoeHmjuCOwmsCqa0PruFLrLXSmcCPi2yMUlhvnsvVE22bChXk6tmSm9/xPJwXg
1gY5aYpKkpg9nUmpC6Or4GK0g7kBgrw/hX298+uhmSCReQ9w2C/NINY7W8oujdln
Veakl8XAa4/2ZOBF5fyqoK89dQlZhXrFlht2U38INUbC583sdaMYV9c2IcLm+R5L
PZxjXqERO051HBzEBCj9F880pKi1ypry7Iy6h8Al7VJiIdbZAoN9LqMlgyB4SR7y
IqNbyMgsoTVHcUEYoWwt9a8x03HZFKPP3WHNjxNpvcwmk2UwWX3E5WKUcE4XFyRO
TXDy5gVFof5KLrNT0PGNTbS3TYESy8hJg5gMr2DuyeFFJZfHeFkZRdmcpriMryxD
dgQ8/K6xSyzz2kLnNdY/j8eYSN4/izV8zUWBCn4vS10P81mzzavjeNXyNzV8fYL/
Sj+Aa4WIfqUA2B8PQEYb0KK5MF6xZOjtkkcv7/iWYJJ152VESFpiA8HiNhiV2pQW
OGsibmVMTeQRmwCuwaDNPvIVnEOxd8RBMLAASCyoOP3qRJYnvHaXWIM2l8KAGyMB
6AAgO4eycBVeEzbuTPjWG9EEoGp4zMKH5wD0TznMYXPBbDix/0Cgk3gMbuPNgyKk
wabnEvgONO9182ssaS8ARiOJ9legwAileZyF6z02j3ovbGNy1BvtdD1opPD4RWmr
QKGOQdBAmaz9t2uFwtSCuHxMIgr44JLe3Ncl+iEx2QiQxEhEbDdjOG7JKHMhfBTD
1dJDs8KZFdR0bvMLhcupWh7/4lkioMT4arbLQw6srFJb3psM9+KYR5ma4gcJ929v
haYCtKJP0qyXfbX3fVwael5aqcWPSHWCG0RGDtcEFxAjc/97d34qBs00T7Haoxyd
4cI+BwfHuysrvW+a53/AbNTWFDy3dg1tw9Yy3WFTNYY8Xu+4NKGurPDs2UBT3/j2
emea4tNqMujxFfyz0O3+F2LG+x66TZdkvflG6d2CJHnCZtWedDq150VUEIut/PP5
rlsmYtmw4FBOP1/aqF74fevpnRDjcQMcJWAOJLIjQAVzpKEieWPxsM7qdnXPpvr0
xIye+jvlBprEcbCk21BKuc9g9zZbBwuAUk0ZXLscCgQr3KpwUGTfoGddxKFF2M8R
WwVBcc915IVcamYYmuKzO/3pIRipYfd7OHrY8uNX0HdhVN4hQdgfsi/sNGs8J5vy
uCc6kJ7dtuXd/evF8AhWqhW3/pfWjw98SXvNj4nRh51r+/+5tlxivrTb1NG8WWj7
Yj7pPpxrsdc7CDFjcZ5t7DkeJaVARjAXChJ06qXy4oCtpDYSdfmm1B7+kvVK0wyv
mcQk8loF05cJXGXkswvA98314NGIWZ5N99bwprzKRrZ1hnpCUNSJlPBurDAS0tDQ
c9DfJ3Hmdrymh2cvXfFR7d/uay15dS6KtKfyosP1Ce3xsx6mT2jcLMXdzMZnjsnb
VrQmU1D8WZDfTawRCNhoaplLmk58Nd0+WZVwPu0iLD5EaogxpWwHfT7bUlj3asYJ
6lGov04eESh6U394NvQzw7nCh5Sbv4R+ochodTgqfagttJS+AdvXhz4JsZstQV0S
ljrsBCi1VZPemkvmdQMxLJbvBiRkzYs3BK5p8Wi4TRwm2wlslRD7rKxovf2jbdms
N2Gkl0w5KsQ0Y3nUebQylVDAbGMYMfyoXmljoAb2uAIawTTU+QRXytF3anz1Ch5b
SSAj2R4ed46POzsRHjfh4xuiqxApXOXbcm0cefW/sOpMYg85gxEMkKcOO9UiOwlY
AfiwAHeKMT94US5TDLdtAN9oytyYovLUvi4ZFrXkLokhzKy9Qq79DRh3gT4g5XqW
sXvfvhssVvhssceezdShPDRv/YPFn+cx1QyfTfqjk728kEWuYqQBfb3qm1ePXLli
Evs/KvvjiQJmnSHnsGc66Hj7OyR7wA5HAHQVCh4hPsGx918C1BqHMBaTuDUuL6ec
ohABVEztGxO0IqAr6dHhHy7oCCPe1SW/jMeuG3konEtnuASxEpIG7g4tSSZD6Ll0
B/SPFnfLT9b5lpm6fx86sFgvMaWyq478uKrsO7D7rSWQglX0dWOHPBJKvQKv2bPr
fX3+DPiQ4Fbep9txcTjCeDwqwAEuymKpqlTwognc36a4DL/kkIUHVHLtC6VaIU/c
k9vrFeOQak3EMTvbmxvwVdx4WbfAz0NVUfza/D5XMp+ZzHmZoKaiKLMxgTGjT2ek
hquUXupCPYxZft/fEzbh28UN0XL06o4Bdf6TmGMCcQQnueLDuK8iIkLxlIfUVEpj
PAQN3xHXX8La99jzMQDOGYitsPzZtKS0hZO8+aTcJ6M9NoSnf7HjwjTmsxwa31ER
sLQW6Loze4LYMPKubJmJwRO1WrDxxn9G54141gIW/A5F7Wh5QvDQXR5fBRy0Wc+V
5hiiysbH6Qfvz+dIPji5/+isLRgyuz0BvhNHrYsNXJ/TnVHGwh79jFsQYCWOd2dm
JgBb/QwBMEgjuKBqe5gnBTipyqZGboEsfo5+M2EIcHpxtngIvgbKN39rl8lJtqwr
sNVLPUbPEMQ3eU/k99ysAe4l3h9GNud0RUutLrVqy7xTCPWXkJ6zT1wUM29/lcmW
HEup1s3KGFO/tJlxTchGcU+f7dH80VIZz+5cSbemSgaCDSI5jHKbbfim9n/xpn9m
mfosdjUKRtGKXtGKkVRfwjuPV3IGxQArh2uLRbmbaV11EXKc966i3EJn0v2DfoCt
wYTP42WlvKhxx+rGPRIppg2VWdyPKE4AvqYbxpNh2hwrW4TmqBQw7GqCmeeXHpS6
RXQiyKZfRDHYdIsz5BMiSo/f7bGENvJa1bdku4Z7aaGdxwRwMcrVJgY21WfKeAh5
SRuaFfM1NXiO2hNL2K3T+pZZLhN2zlvdzQaqIkFbxbWlpVRQm6wynd8tRxiDUI+j
nBVn11z8uCsIu0zq/27AYXWLBR1dJ4tD9iaCPPacl8KYXnqOe2qcipt2hr4lJRDy
tNsK1oiQOf6jwI68/xlQO889fyEhDTcQIjyzEsfiPCYdmzcCY5HFs2x/SR4G0fNR
ti/hj0jNex18JonvsaWi2bi775qIl68xH47uQVb3EiGHesY1ClUlmiEhmYiT1G6o
JHHVrglPMGzAW6lWVFBfFWaADhi/8/qNwUFM51IdLRpwQb9ghzGYKIGOdvGnHxvG
VbvFvn7dA/nl/RpDkHa7u8Om8LxBiJTPVhwEIhLjSKfJa1BWR3eddTxbpfKP2cud
pLnW+8o3rntvn0OvxKypqjhIfvE5ywOouwCjf3Zl/Uijj6+kCMEIjUoL6P0geGcI
fU+N9kCCk8GSQiHw/kzGpsN9ApCfu2HaJAh+wl7ctYyEqKRrZqkuJm6NcYk4WTsS
FoFL63jFcgXFDyp7M0jTtCdtlKUsWIL7RzHjhCnc1hTAZTkI1MjQRrLDE+imuCaV
R4n3vD8d0tkwW3Wp8dSEC052IQ8OSVixs+/014ejFOzsUNnL3m9gad3cqt6cU7yj
uznimAn++iCNrET1INVunXiDsLOQ5KPROMWe2Xxfy7mTH/mwXWqTmuRyhbbwjQbN
bp6+ZFHmYZbJBnPWMNx8ArDu+CKmC/SAaewLxKASG1kM1aQkqghUC4p4USiAj316
JZiAfWIShX2EW0kyI8tGs1nwjvNJ/rdTwKAG7aQF07Cti+x8IDdrW81HRGmxh7zz
mvs+69z12d6JLqA5DiDa8m9/le1ZMOBTdvuHqXchD6otf+y2G0xrMixjL5KhZZRi
u7Uq3B6Xe3EIA2cbLPmntx8InvSdEx0oUD7pSdC6CeEBWRm797mk5VbFG7LTXf3r
63kDBMKCPcJqsIOSCdH8aNhvyp7CEONy8JFB9e/FWQbqWegEmg2V44arQTjiZT/C
GlWVQoLDkAeQ6ox8w9UyaCNWwnMiGoBK16hYkIHMVtDb2MRdI/acIVJA41IL1Hve
hEUQwQclAXUHa9gk8WNt2C9WAsxjEEwo2Auxmtf5Maroak7TCY+Oj42RKcl22wQo
JvSezuNjN1MLapGIfRS7KeF+I1Ph46eESPeJW/eIjF9SgMjK/IFm/tm11Xfq+z/d
2VJuIqfqucwQiY1vozaVgs3Cmgims0r+oxSzTgMbRBYwbkWZyH1VrEJcddlQdMBb
Ke7T7/C9A855uctO0shC+iT14LwIQWOXaYAvndlL05rhIo6Lm6atn2kwD6twK6P3
JTqg+K1m/ljNYoj9Td9Ox/O6MGS399z0Xg0gxnFpWG4iN3DbahMtPRqTdz0ToHTf
y1dDtyuvVRVx+7J3zLyvG6f1WutwDIZr+47SibXEdtc/6Xc+TogshZ8ax6d/Jv7e
g38P61gWXPjGcWqC0FhY65i0F9mpVofoBy9PkVQXUq3kGdULMLD4pCWxUgt4KNlm
HoRiqH/2U4haGdED+gU4pPDO+FjvPer1T4xW9QOE8P5f7N2gutIDAl9UfTo+qqy+
wcaJBrTXqCMLXhzF19XEqhQQ8+uYJNwp3f/fCzzdgY4sso9ET+y4DIKT7Zh4Vaca
ia9HJ808JK7rDVxw/3i92l2MkgYZjkWmkOrMg01vWN81FlXUq0JMo+xA2zpgrntd
8KYYJd+P1eCfh4b0tCWhQgHDJINfG2T9WRwzhAEcuhNjzW1E4KZnXggrQRrUHsnW
Cx/XqBHt0lmq8I0dPO4W/daFNDyJ4jwfpNOWT4ZV1VCVUAKpMcIDm4CzCKMN70L8
w9WNY94tgfz2dQ7sFCsipUh4jsbJft85M3THdPLv8nNiTparCWhY1ZUPOnPpf3NU
DLNI/I4/ax8EL5uE3mcCvRvTGnRNxVUrIfg3CeU8ElcsYDNLPGG0BMIAG7PsFMww
oM5IGKkkjtGxISfaJLvUzOXJkeHcqT/L3OozdbxnkTxI+vBV3yvjai3LB1KH40zc
4L4hMmKYfLw8SDuQFED6EjpQNuT3b08x4AtMwPZvpykmpzDb09HKKHZ+igCjodi4
BI5x0onlCqXczJtG34MTZZ0l7yD9URLE7EKDu9/8Pg+WCRGvy7v/v3ubl9KxDaMi
HyVPuF5t7xPab5rJSO7Xwg==
`protect END_PROTECTED
