`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+mSlCv6NNx5YR5QhimpATixnbXv0Cc1RIEr+c5Bpr8WwolUKyjXWWcEgTfmijGDO
b8/hF0eLq3KsVbY3J6RwZBC9dUsCoyVwPgOh2t+LkTYjXo4IQQ2lDfyerbm4ZYmX
h+gDXq8tJn0I/GQQ7+gkc63n8vU9uuwx33FbCYUawDnnOcW5Nl5E7TfRAk0dA6bS
tAJw3hoKpAIA64GzVum4Im1M2PHz1EqEx6AevvY+XZy+Gg6oxulEPfH01KHIpNnQ
QfEVRZ20zml+/5iHevV6zdBmxaAKALF35DZpACgI5c/2cAf8lMIM7kL2Dgmqte9f
1P4lx71j2g2uTYXtD5/7Zp6i0MFeF3C8ud6x9ouOsmH51xzOYoFUyNlRqiMZvHWV
tBWc2QxgiYNm79fvP+RuFsAK6aHZy2E8qAyReomDqYiPOLfxVbAKkiZQwFNsg99W
wUSqHUpzObvBXhYnZ+P61zW7i9ABHBLfK2foco9PrdrdCa5bKfbGKoWg6YzosRGi
Daf+LrAz97teC7NPYwEoUeuIAwEmP7fmpH4DhJMn8BzAKFoXjILMgqq0dswsS8mU
O/QZlNbukoH4eXGpAqTf0kHddyBG9+fPgwzi2dq6euoHHvppzs9MUYHBOl3tIIHK
ui+jFCbY5tc0tY55Z/251XDQeBFVanLEZrCRYw078ejkObR9HUC6InGiLTcl+j5Z
QOxysEbqfDhiOmK1jWdgokbRaGXKiZ4Kj1rCGtl4LJaPtJTPipgjpDdb4VB3H+9r
o4f6R+sbaV030qHGGWI/hqSIXvfaSf88TJAqbXHoYg1ihfvx9fNcLGiyeQb3CNHl
aPAMVauK9XMD4TQjd+sUjtvoqKmABHPMgORRA+ez4+PQ5tOsXIVitl9Vi4JvtSjX
+rk6nCvXLMxW7C/r4mD0wDHMszaMuEnjqRu7Er3lgWWxgMOqnoUobqGL53hh+/+6
gDxbHKhnLEbxmlaYk8quVlU2mP4NRAk2PEDDSX8SLcJMb5SHRm5YKqF5Y8CbkFGW
aJABK5OlKddbTqDA2oBVjULsc+TR9KRztlktkgtGkdGABC92QZ8AAtPuBP62TaDS
qJamudDoBqL3BqB4yFHXLxOk90wr7IYLAbknlfOKvbAoC6KBjKtcuXQJ7/mgWYjR
0xRcYAQvfzl8x0T/MFjhpPhnio3PzdhpIDPlyXsoezuNRdBot2ad1nwRlpEWQ3Cm
v04vnyXwh9Q3CoVbq3GKVaQCSjuSt/kd0SU3XrTvVl1MkYNeM94pXX87Trmz+jZg
ZxeUe3LXwZxl0DBouDEzGndY/Sg5yaV4XB+s0b6/6DFRUJV5ocGOsnzRsPzpu7N0
j1MA0ZGDmcx/oMbHYY9CX9Po9gTNWGwelgzflDSKofrNUQ4Eik28iL2hQsXlRSne
gqf3yUI6fXns+qgJv9+SqLPP4bP3LMmFBMLsVEZFiSnHeRGuf0aYG7auYQQE3a61
rEbOr1z2tWk3zfm9+KImnLHwdunDy5NQ/uYiQ/rq4WvJ/AX/VA0GzSBWWk/dIqck
L27yyRwlyHeLZN6uOmyzMde97v7z40SBF0gw+7fFCdX3C+Kn1bqu3fR8TDUnUA1/
kXasjxUTx6sq7i0jPfopjYhVcFr4cWInvaWwcoKlkLww1bG9MBSd8/1X8YvNrU0B
neW9zy0dQwL/Klna5M37igZCnk3YhRN6ExNs1OABKuYOg1O1eB0sDxDUNMSZmR5Q
cvayRPtV0cXg30Rf/kolB9kAXX69zu8dIgxwPQNLozH6CaencA+rqNY60Ov9y+uD
KoNsIAqsyyyL47Jcna9EtQ1da02/+IlkSPfgm3NNkPN0BJTnOa7+ee1ZMJTIwqke
Hu0Syc/ynU5XyPH+j3dqP6X1CZ6XQY03Y7/lwCdS42L45yjeEqbr7zQ99Cn1YeNL
ToymsFtXr2AoXyAzGUn2LXC0g52dUKdCwDKg+8w1qfnVigagttLs9BrJ+rXRcWx8
QWNXAH75TejmWbAhzVFEYMB+lZsbLRN2Ed+mwuy9IDVEcEgkuTrCrlQcJH4RRm87
Shon8gjzr6EE2Q4LilKsdlyKPHNaXpT2YbweMt+G1oiMNCCHP3XTnOY4Y1jsFq+U
y070AY/oPe2dUBISMaS061T8sVb1PvlV7kMny4oHsr3NS9xzRlOMXvE5C+it7B6h
srZLPED4Zw3z5/eg/9zGGzZbbFueMRcYojknt0GDJZfDpSes/hUL6PwalV1qRZ7q
O11v5eZWpAm+MJToPtBFMLYe3mZrYaKWYGmhP+f3d/dOcLRrR4cvgfYk1fwtzn8X
lCb8+KlnTTSoQNTUnArzTb4WxphxvuED5rf2FUGN+8Sgo94UlhmLf4GFk0FzoliQ
jvBo593FAM6HM8TEaEPCYpBXoC7ZLpJMCPcNGeAEJ+JH9lctYVUPeASmybD3UojA
B0kFsyw2FB3LTUrkh/Cqq0e3XfubStb8H4boCJ/Xwo81gU0KB76aOmENWhAnuif5
lT4ZoBnzepiPEqrovU0WO8IeDz6DD90ZBv/LBbLSn0KhQ2heMOUrhiOZtm7aSuvu
aEyW+fGRM2Z9ByC+GYWG6Lc6TwC3lqaQvo2JOKC+Ng+r9pzh2mH3lzGTX/7ctAQS
/I04Iox+j1HUcxw/beo3sm8eb9ut3s1AaTPs5xT8a0sjAOwcnoyY3k9wu4kIRz0z
TYOzu23qCxLUWhPPGOzW/p95TJyGlkLxlG3BnVG2cV+FyzxyX7wPeFf9DoacuNM6
B6ziN1UGcE7Pt0rbV0O7K5WGVjDBfWs/wnFQ8WR5H2OJfrn7Hr/qXe/02tNmbJVE
oT2WiOXjNBdP7qP/dLLp/lNvYpe13eE9Eo/vmWFME+fZ/zwz86UU7lPy0pVz/+wd
dlCO8x6lAPvwJEClcD1bL7anV5sXh2rk16GfCtI6XtSaB/zvOahrcMxDHNe8JXE2
wJ95+9z1GMipNRXiH5pHo/RYlgPVdvzmaNXb1XT+VqmWOKJ8ZhcU8Hd5aX0Y0yC1
PBmc0F11GGr+c6Cuzn42iS4TN05fq4iKzbrmdOOwBzAyYtUa6DJ4d5s7L+vNSUHI
IarUpncULPIh0E1qoKAVkKa/EFITzcqIZhPnvCE1s8Nnqc/8qRxEm8VglHula6A6
KJU+y8vTqWeH86jjVT4bNHRkc0B+3gbOSSKTFr46SjuE/eAHpkJ9Lfv1XzeQc3N3
fpmTxLiUQqVfmLtwXA1lw+DjUP7IREwnqUXwQkmOCC6gJE38NKdTgruD6FH1VdCo
0NXX4Hj0yO8iTBo2txzJEEbSBEYzWstp5QEfyRSaQK8oIc8u3jI4YS4lUdi7coy+
wLDfYh6W0uz0A9OL22znFMd+iGdIqwoipn53QJ/QDLksdmU7SGQym8A2eE2svBSb
BOVm6vnKfnpgiqZr7fhr9W1B56ZFQvHgndETMQpdzopfImUyNk+ZQkHQz7d6ROmd
cbrss7lroq1J0ET0iHe6XzmPYhGMI93J3Rjpflb4sw9NkPbwKXIsnb3jUM0lR7l6
d6vz3oyJw+AYTq5Z/hHl6MwlZwKVJJYjfQVHlqGUpWk/+HSSyaiZKWel2GZP+PPU
dWqrNaXjDQtBBdwJOee/J8Sp4YkpbftA9ZVxId9kR5A6VfQOyJYhvrOEfX3x/rMN
vw6IaBzUS5AYkXF+VXl6wLx8edtVAZLov7mcO9IpJ0tOGwyLZ6QbBnpKviH8wKLn
mfTnsB7nCC9ic4dOf/vJJV3F4gFCGIfXltZrv9bTnF1L0u4n3VnjkDBenP5eYGOW
gBlhL37pRN39kSpfQkuiVAM5de4hfqWJnsjOVOInRhA0WTyW5iVL7eq9vZ3de1ii
3ICzSWGLU8fal6qweaMW1QZejpTYCx1ze4FmlAf0pVpzKEWuOFWivuXXzwXAXjAp
8kwfRbTHPS0Vta0Zd52JiL4YuwjnKYhwkm+7mbYjWLOxgSalTyPUSpXjYdC2v1P6
8q1v9+G/P0epK01T22T/tRwIuFO2Cn7/YQZDZopaaYkrczT9lbjThceLbiU2EVXz
jgd0jT9+atBIN9p8bgKF+48zsbuYEkbmNWO9gJR4p/yi1O+o7oAEwTi5SGcz3p5t
Q2VWeJY4ejzPO1BGLj3w8JP1sHjJPMewxKIGHmMlHD1ZgBHSO1ulQr+2wNcFnn8Z
WFDu+JlfcM5SN10FCVOon4jqIMUDerTKuSVAmnKSX2z2ogYcNSRfIB7OWZet8amh
zru7QVhcaEJrIR5v4hmx5w+njR/j+hwTlnwYV25wtoEkJOpAQEAbek+O2tnVTkSS
7JC0i6Sekn2NzPq1zYtUUAoZh2i6Byb5XgpzFoQpXVqUaLJha39Z+W+DsQXB6zTX
/oTWjN7t+Mib4mutBJC9NrTYn352k7Jyv6UQo/ZY29D0up3Zoq+RSWGJy8xb1U0G
Y3Hd8/4pGAMx+oOQ7Y3wQejaMP7JCV52Z6yT+NtU8Euq9nUX34fP4stBb5p00N6w
UzY98CgCSiM/uqILFadIuTGcHhgQOd0l1jwSpJIhWVuH3z/1+nAJdIJQnWL9JQtX
A39AOwmb9kPKz3KU0V5zBYi+WxzMej0WNEUi1opPMtXkQri3zX74P51/q+9FjZNQ
Nu1MOFFjc9XkEWMfBfLM/YUSS634atmnmHveXamrmeYIgl4RJlEi+CD7a/Jeh9Yv
Suj6EfOiQeMUhF1Dav/eTKI5ZFD8yaYnCtWQLmUA0Zwp+KXits4Rnktj/skLEFDu
fOdYZFxdNmXV7kR6ncel+xM5yJP5ePK7jjc5MBw2AozVl2HVL+t/z01h5hc0X9X2
CtjkbX8bn6YVSy6pqf/LZ+LH550Fa1SekGsVuVOlqzaEEoghmpaegrdCLk0E4v4z
WnWSD66KYytDzL9TtrUznT6eNf1cgJsLOvT9rhIVJqwVprEcoc3CF1bQ4lgV8ruu
BS2JR0PXBAVnC09+MznVLl8IwPYdP1NeR0Zwyd+FEHKU+CKpS9ByvynKCLPDlStL
pb5f7E6m0QqgPQ/+IZQAzOwALKzCSQlrvGfMbD6pXIG9lySZIRPFh/4hQ3/0foS/
/M6oe+l9BHgRKAsHdO5aStVf6MGlmgh6E/paomaSuhQeMGXR0+GJX71pEWZZzoGz
IKiZB/uEemU9dmtFSpTnfssha+X7Z8dh7cBSsVPTV37MxG1SrGueJYPBqcS1G1/W
P424+ctVfSnZ2/Y65y/swL2fL1uhStky/eqnUDMHP0eSEUtPuLuN2ScFNfF6AuFW
9SF8ouIGCAuh2/OReogLaUyKkn4G1f2Xzd8x9bccpqxotBK48V4i0GasGXw1XvRM
dj7Gs9ft68y2RpKwvmBHXJta0pPobfs9cWgHiXetDeu8Xym2gIiGfVxAnBolmRx3
R47237yBlK9Nk55YTtIPN7pnmAMDHOIychQ5PwX+iNDEPYhNVfOh1YzStOicDLsc
YxRVgamM0PTkXUcnfwMyYhUyCxoyqwuYCn4Az74p9/d/8OpyYb/CLwwaA3Bgjp50
lGta4C/m3fyvYccwvO2bDyb2lUB8/wJjnPzhwjD/dAjK8aTWHFTQC0/jAgb7h1lE
4IQQY2eN3P520zw2Dxs8cFVkBMGxAoSW6IJaJhT681toSh5gCCJIsy5gQswb0YT6
yvf5+wyL3DYKm/jvMSbhkiqI7Vs1qFLH7BZBO0DjJ6beMO/IExzXgn9la1svMNI8
5xqj0HN/JwfZnqXeGVlR+c/PbFtrcifZzx12Nhta+9UlTSZkLuOKeKvpzzqL7FXL
Q0a7VoJ3gavF/MWY3n543bLQhqhjbq4X0PET33Yu/mvSsJVWl2EOLe+kEwVSoD+U
7C6HdWOpzE/4+518JgMg92IB7eSdVN+nzgCJw50gcJIh8own5rqe9pR0yX9wOghq
DUQqfDC1VwEpgjBW7nxPDDmO141pk2vxkJof9GZMvhYI8FVE32luACM8xekxochf
H2bdhHtUbwqTn3aUxsJk5YciaOlzExTdotQDbv1e5dexOYzTJ5ZrH6EWvfoObX8C
aq7thH+EG4ca/W6khyswv4mw3oBuPyPXmYKAdKIcFU0ZAE0oFAeVHYALKJY9Y+1Y
X/FT8pH1lpV3YaA5RE2UvR9SSECIDj+LVYmwcmxpVjwQvfZrvQvAdTNZzTk1jT5t
60VagsHC0+CL6+8BpIRMhx8W35Pqxf8LJ9QKR9OGAmtXlGy6Ezl1yiq6RBcelDIp
UEMnUP+Ehd707QhcHgBFtD6QUh429FAmCVUlzvIBaWqG/zIAhaF4iXa4Hnq8Jb5m
7xGYw5NwNSOqSKAOoC360v/OqYM3KZG0KL7fMEKob2tMQvqh+95Ru39kWxCNiRsb
vr6RT65MA9M8c8RI+vR2yBpSUHS7OyTYdLXG/iJNc1VL4BIqS03fpg4AQE6l8Z++
f2jthNAOqfyuWQDCHBKKz8IzXvfGK5SPe7BVJrvheAMFR08hNoBgADKJaEJVT0D+
Xq1y6Qmce+7HH6ECPrDgU/MdsXjBmY131dAErxuAOhDaA5lTM97Ot5HfnPuCUUfB
FaKRQOmE/kmkYDfVtlOdILcF9R7fJCQmhGP2BNAttz+2p+TzoUirbpSTUwPU+SAU
t7nET8lNVuLqSV4TYRGtw+sgZbwwfmRfoyYnLkycDm1rc0ZY8RFlBgULZ81HR8wE
LLlgRXprarP2sjbBE9UqoF9wED4oSx6iI9DmRKxxoM+HX5JXow1O7dxEPz13x4dI
lOb8K4T/pLuOrJdncZHUaDsTfj9AfBv96gZFEq+TuZbryRYN68dRyADFt5Jkryiy
Aj5f/kQjCFSRNoFs+UJ/ZfsJoCyjWkGdHOWhOAeS2EHOehN3kZCQEx5pIdTwJX9H
empN443Pb8BwkntMJ8GU2g8WWhoC9mMoBfPciVMKfcZFFNs9uHR1qO+qOvsC7+Nk
rM7E8esJJ3znJpYyPEi+5SGGBiHzTcam5Pvs7THN1UAPixRgQw1COQL9cgaHXP/e
WtDZuhmG9N2qfJVLFPV8ehJCkpmjVQZmBNFBXrYzsvkC1HckCih2vbN4NmJ4T0Lc
63RNh8IMOuaGgepqKeyzY/18JnPATE7LWDKvcxlXwNpb7aCZh5ghU/pqUXVVuknT
5dmqo5Vgk3iyIHRDryGmHG95FzoC+r6ZlHqSX20tL+cMIF6e/rr83UN9XgiJ8Hox
7t8tiKtGWZQBWlv53tN9RQsTeWvlx/r+xoX8N4LHL+s6VSkrPPygiZuzkk/CWHog
XKSHbITR0o8YAUitvueB0QeowLcsKLE0EtSiBwa4hkmdc8hWvn4HtP9B1/ayka44
xic1cAylsbAhGD7oFD8Vh4CfAiX09sQ+MaRbIZz/4KfNIUpqP3LCkPbeuqTz4Iff
oSLZBdvBAWaxIwiCZceu1yeOHULexpW6lVsEvIygmMJeo44chbhUT/BJY9knhlml
3DeA/MHZ8U2ydMJieGnrgsa9rZCbiic520ue2yj6kKtM93qUEe6OZX2MQE5Pdyfv
IQ/HwgU0UfG84EkPdP4DyfUEO7jnzQdQYnmMt766zAi3B593dz5eRY4POuRptitN
3+qmkfQAL3paLc8R4qGIi3mEOG6rVBswgs7frV1iNfCdxBBN+8punJqpYdYsS9Eh
5vtBTN/mOyrk/av77PtsUer9uXWW8RKXhdPQ2L4Adqiv+Ahf4evsZk1KRl64zC4k
PbIU3c84500B2vBOBzErlOoQZgG/C/nk2hcJaA125M+1fam+MeUv8hYXmF4MXNBH
sype85mqrpM4RUmz4MCgQc3R8avIckGFdpZBBp2nCoZlseuIOXGan2rPf3jsWP9b
+UQIAG0nuRWxFj7+5saBxTCDZr8O4Bw/j4IFBFc6ieCfgBODblGnblFYkR+L32LC
OgregkxbbYwe1bJKa671wWVyF5G1ZOr++rDk54F1/cOKzUAt/YpeHXGI4UtR8jss
Un5WnI9uM8UHi41xNYYOU5bRp3Tz59JeeoELC2Ct+JsPrth0skl94RDFQLGvTbkK
7Im7OCH+C6DziOoZnmW6/lOaXzBPard876k3WkS2giLpeqEHmsaxWGedjVOv4csj
Wx8HcTnlAOwgJlV3OEYOgUjiJAAC+QovMxoeHjbvOFHwqGnTrxg86lkSBc9wzlaI
kfK7oRXrpa98i/WzajSGLExcafPZ72wIwxJhLXvTbIFL39E3+QUm2rFkI2X4GaYq
Ho4tGJfPObMIqNiGM+csD1FNxDa3ya3/YzOjzmuz9HZjLt6ZpjaqIcODELwWW+D6
i9Bnw8JldZ5I+CNP4IS7OcWeanOWVum24RJQaHZRg4Izfjg5XVj6Hm+0H/+h3cXA
t9LqtigDzGlleA0it6IEsCTFozQD7fiSLXFGtfApARzK3hAXl4oxWVvGWTHBdx18
PMEEmycEPzFo4+/8iGL2CumO0ZKCnhgyYwHU3iNzEIkUqcgeXj3QXQGNSx/uoD1C
79BjH+3F3vbg+TP5SIzLp+i6wIBsc5NCRxNgmur/9vKnjTRW6wDMJg6+9tlMgmN7
Y12Y45sBIxOf9DPsEX6Fke76uJstqvAEJ9G8BmLzHyQ+jcZaZaJg2KOlsymwo3AF
pnXPQvou5ams8RuJcM0vrKttRglzZWVcWzFO6GnRvnvwzGNpXQhg3l37KxbS2iU4
LmWXonw+9N1JqzlIArQjaBekdgxtOTTJ9sGAMUySQEfSrho4hDfS5hkq+PPJN9ar
8d8Do1hQr+/iv1tAXy1DQFSbWDhw8KHCmBhL+JkYEreuN6s3aSLgLCMEVvUFMptX
/1UHeBs+4cG9EoGMG9mHCc04gaWVq1z/aa5WeWirnnYC0wf/N4ZycvFF3WClrDLl
Xx5ABzgzOnwxqMob3W1LVJ2Hw38U9RIOLt58xjHVb0QK7f4MrOiyFbhPajof0N+a
849D8iHbVxf83ujfr06DrkrAyOycCBF8/06J7mqDTZDx6YjcKlr0VmXxL2GEL2b3
ZI49r0yWt6Q3VMZhWhEuoLpJrJUOui/OoG3sTITklYt1D1fP9bkZF/6x6eaMFnrD
KV3fKT8dlUiLZOT/qjZtjVfLTOZTHECM4RdRQG0WF13PkQWGL/lcy7+/lnk4RA6a
5f5grCxMSo8/fqkYYiKxSWr7NrtTJB8n16Ca4ego4b3SdjW49uY48qQYRQk9zUq6
E6adb9bsLStgttSgSc/UU841PerkLNCkK8trAT8f11VBZQJqOY1I8zEyC9mmF2HT
URuFGLW9vBIi01Ty150XLZrTTbYhhcC4nz0HR9HQCCckJVm4sgqRQkrUSvH2kboX
BUMskJ04/i6G/3gQeU6F/RL1fH2vCS9IHyrd6GHVCMCdnE9g7FH/mekZVCN+8qI3
fYG2GnNjTVRViO+ArjZClqDHUU2NmGuc//yR0Hc57nhH4PW1XpWJG5FVGb8KtgdN
Wz/zGWUet5+tdG1p/r2V40CBxSuRaMMDqkm1wqUqRJUDm3077BB2kB62ZtBMd0Ii
K3RGXG/NPI9DPcxZ4gcx2x8PNuk6PdD3sqNhwpmxetm/dE5BaLtDwrbZAhFPcNKU
Bc5IXpJDgHYj6B8wLhssRpJiBI/pPAcZDvWr58zyFDpixBMqRMQxnAOKabtwnV1+
/U9Hsv2kAK/SC4p1em+zhF+RRHt7gEJ5poEr9r4bS9j+Y64ifD+uzJwznfbrnngz
VVH84hQ6DfSt7hFMqmh98jmUqNj1wGzDFUQKmiTSniPyh97gefxIoZiaI/Qw9KZ1
0byj/GE3TDBLbAydw6Gj0lQskpp0ZMUh5ekbRbIn7iNttaUbWg3XUNdpRCFvxo4a
FhDD0GNGy0dR1tUq+R8gIuelnfagF09BUXSwfSF5C0C/nBll2kipuerYRIrQ4770
TA5D5FkP9GhWFagcM83UEAk6bAQnpgUulUHkhNzelr2irjBaAG4DmEY9uA05uCHP
gqpUpmuwGTinWo8hztDY8PegvV4Fr8RORDbdg0IXgBp0W73xdy0g3sWi9ZXbu++H
LenPiFnNM7wHytUD2XshLl+fSlXd6nEvG/r479/NtOK8gdApafGTz5JhZwU+6Dya
yMrrh1qw7bbTdgYMfqpatlkeEu+XCmxsmth+QPvGTwdq7IjAVO9qoly9g8LUXuUA
ir9MXoksA3Ke2pMsEsQ0N8d7sir2xb9cWvYz3QNrhnX5o7+gX3Cvdz2edJwYywou
U6yt3a3uJ46Y6NWZ1kwtkAlY81AiH7IGnCpiAAc2ZTomCfwu+gDbmUVPkGJT629i
OmTThMURh5IE+iKUm60kxHEkSkB008USRZKAKm/mOaOQiQjuOdsffso9KywSJ0Hn
MdCg3h5yfyYab6VzeFpcf9BUjne+9vzgp92zftpKQcI4bI/kQoHKxjbku7r1C2PD
JlJDgqFiorc8jKu7R+GVgn3M5y906XYobMfRtoeiqgpDnPILV6pPGkZSP+hRIUr0
aAPbHnKQecKs7qQrHB2M3CHT4/FWumxA7jACuFQv4yyWO9XdYFLJdHazexTLanRV
rSBHZIplGQEZnG6wlecLVDKQQOJcPooB3OLaKTcQXFxw/0y0CfRejM8BR2CGWsng
W2X062JNwJ5dqurkfSlq6itpulUN+Z0/QIg02G7a92R+hoohb7yHOfpwLA7UuY8o
NlW8IINFQ0q7IfrhLIgUnO3StDzUyRj9t+UQFrZTGEgQRs88rDzbUucvpcYTTaoy
GbRbJKbNUVmcGsigkQp2gyWwYaMkOL4BxoBfCWTH8ogLw/KfzBpZA3lsFGIu7cEv
TuPbeTpuQFmSbVtS3hikXr1rW5F9HJc7y1dVcmox8MAottzPylcw5XNoozoJiXUL
hjjk3dUCNdkRVTidQSjhnuxb6ZlDnxNFlqrjTkfojQ5QWnRJoWREuaaHxw4DZkbM
iaY+hdhh4DMO0m9z/MISIb9M7VZqSaL08iUYEKT9vjkwPMvXaSe6I9udazU1Qs5h
0ivQhbOaNJ4dF0BqidkcdONqvZTS32NsRb5jTgDo+HmgwB82ZKYplQRWTPL+L0ku
g3R4oIv2L3vZkqmhHjVzezinzGtzAQApBMBdIL70Rdf9GyNWQwO+njNXivVuY7xz
MccnHqjeobJip6eYWA+pC3YOHnsm5IIFwI//eusp1hq2IUiMYoHy+Y6sgvW0xjzL
lPFHDEEgws4eeQQZjq5rktiwpchHRWPsYdhvZXoICnb1q2vXGe3G+fIvEe8qHr4/
Ioh1RlWcha6EFH0+JrYHHymap9A3wldac4MvFoNqb36fS6BsVLj+MGSRSRQHKB8h
IlUBdWY6P2z5L2cMG6SFRCDSYGWAuCbuRQ0+dpijEXsV/5ODqOIQY8ZyxbWsAJQf
0/wd8qFl3WFGlZHl1qY2BDsK/Jb+EfBP3pj4EbrDi3X+3Cznbo4TzwA0X19Ngml1
7Akj9ycWQmKuJl7DwL3/v6gztL0DbFWSOeuzV53FPuYE2kxMuMxMTS4f3crX6UOM
0TSA8yX8IA7bsgDlJnJe+YztKFHyjNNRyj9jmagFvVVh6KxM7wa7NQYZpn5TvkSf
nSjB14TFmZrQcawONK9y4OMCrb+7X3JAnji1XKgBTJyt262zhlKXV5wL0GjIXue0
C0HyWh+p465ysIcK+x5bAfyvtrfTWKwO5BhDeCn6r1e3IMfv4HdWC5cLy8AtLkWP
7sjXR1q1j0vxuDLNrAIPlNv5/8evfISEJRYj4k9akqfKm2za9/3Qf+Oj98mKFOlM
G6WQMXZkAamv1QGpKxo9N82XITIL6wbVWrIcnx+66k8Smz4NF13/UuxykuNM3QDh
ll4H2ls9csm4H+4UvtAA8tzOgMjjoOJEw0k2rY3/srzIWOjXMgJgFx1sInPdIc62
/HJqUHIyBzOox2XyPs02xY7DBFRaeG1l1u4wlpaPAooYQRUC9B3V7Jg5kYt6/ahE
A/la0GbhMmRDMw1vEdHOEiaIcb8FppTMGXA3mvB5ONiETqBOHwe+lL5U7jkduwKb
+YcDEqPHUgbTaSUGzKhCPH1tiNL/FtlwoSwl1BautRRXYn9M6eLtjtoQVdD6z1ed
V52cn+h1yisdy1HfRjfb7kqTBm4N9bZMpih0zNy+3IZmAVZbAHxPCVdzMc7EY+v3
9q9qA39hNzryLmwsjdEOrSBrYb3GAZFGf+Jp6y+HFEkJIwpt/F1U5T9P1hZBaMI7
pYhAbscb4RSVD42mWYkJcBNK2njl/zDxTYtdBJh+i2UBOH8nsovwGkIdZcQ02omM
CWrlugr5a8G/A8C+l23G91dCCo52LFR3pmMd96kUJ2gQlYA9jHekJOIsfXiFpCIE
6DPBAbnK5bvaxBkfxukuzEdUv4PcK1b+Z+2dHRaFkGz7jlNwTCv/S7tpy2iTiM+2
BcD6Gy5bcBbQRMhQyjUKpdRYOJw70yDHzicrp8ZcZ2QpjqQZohqASZXOXL5fLhbq
NE3/p1rSHD57Fu1VTnDA3cLv020yUcq+kkg4cHuhbmUiYyQsZWpUK2KSUKJmAcf5
z80723ACC4EOvG1lawzMmbyBktuNbvFwOo32ViHF/5WZ61uu/dgYNlTP0Au8h+NO
9HRxaWPERdX75+QNHz/eb6xFN2s/1w9+kZP0hi1yG2LlfFmAMhc/203E32pJnCsK
YLvq8o94LRVJrGIwM0tp/m0Ti6N34n3mM8AOkw9FDnODE4HQoBiZQweRW8SeDwtL
EwEjJn2loSSYei6GLiFkdmcTJ1SWf+c+zOSLnwkBE+xEZSrCQVn2JECyC0RDcn74
KHmAVAkVA6Kr40HI4ZILCXpFOsnaaHVMwoV+K4gUZ1DTJU9sjk2OHk5M0nwAMh+Z
KGezFezWPTZQP0ginT7+hhC9Ylw6JBFSz+YfHdJQ5I61nLYJEnvx7E8nhcugZAih
sWEHZx7m3kcUucowH65bFUTwZIB6zkawkr7b1lJju7YyUJrzeMI6iVKGaOgpMAkM
6iNhig//4tz83RGnlSU0unyuLm3WzDXq4Lu+KKO7NzMLCyQ90NF4q+Zpm5K19t28
lSZD4P4V0jDWbL1c6IrrdcqxDgm9rcqpVHxeLeNCufl2NesNHlBOhdpq0gfhNinC
1QXtTNgi5KKJW+5EMKbuW7PutjzbaOLoM0kUw3KxeNx71bq93FTDOi0qwVLlnsYq
Qk6ip+d+CfKvE1plVa1QtrX7Zn8eyj00sC33QG/5J2k4TnttddX7R91n6oQPN3hp
TVCghJ16GwX43z1/jt/HdsFlqEne9sWJ9S6IO8FvvCYsrkJQAKbbEcRNoHgZi0cA
PExWFoYM+GH7mjOq1SeP53igqB8ZMdUkZrw61gdanS2ZEhE/uy6S/WRU/D3mpukE
JIeuNw4s2e49GxmtS+iQLsn0rgL8F2rYsFOp+NweNmi6/2IA+1TbeFjY8RBvZyAR
3YOWXqsfgD+XRas1HoqKUzysW/fs0zoTcsoXHqlCZiE228p4aYda4Knmhql81fB1
NLGkfAjbvruXn6tj+hfiShnqkqxeV9lpQMGnMmtk5NfH//ph+GOSZz09XGWLNW0e
JPHr2w0057s7DEDRK6AMy1jYZ9YGcja2eIaxVFvSufwgPBusWEfGOtc55O0bYB9U
1ng5zZcZByu17m4k2P9fgn6JnAhCl6mZg3wZpgl3Hj+b63naq80jynEJkm3s0XFD
T8m7z+JgMmLlb2eBJIIf1z6vamAY1uJmu4cL9BFEVccURWP7d4CC4aLA2n/Q9MSY
ucocDGvsuqqmswwK8pykZpAaSSNJMKen+Q00t3cIPb7HgqPdDSnDpJMNXCSSvoFo
ayfDLdD+lrbvWFAPnqeRbPzu2dBDq2XN58bBTZ/QRXJtfgoFMv6gND62uwH9s3fc
0AxxzS/EwBWIOABWKd+/wt15hZ81+OizD8DrdbwCc7Mhsm1+TY9ifW7DlcOgJTxw
/zZjFnIaYt8qvfTUQpjyTJwoTgRbAOgxEbvn15tUQPAmanK/o6nt072ATUsRHG4+
NGB61BnQCisteMmAxOHn8oRjYiXWjnn660C1GfRpnpHMGyGemm++o/OGfxCPiVm0
Ov0FwcNFHfgtDKmGTOFuxhUTWpv5i4yqLiDhfwhJq9RTKKfLkolq/vvZjfIhCCtY
9oUOl+lvf7XRZwZwcGfg6YhSWh/UxHngX5YZ2Z3ZbTzVgSEm/W0qpamyWEzX0mTS
pSCYHXwe9hJrVNc6/wF6jfeAlLXpTsnK/KnawEs1J2aFUHlg8Q/37MA9bjiXmSXc
2bj6LlM7MCQK/3W9ytnrkP+ZpdZwbECY263oPlzMPxPgAU3I5xrZY6/TjCJuM2WO
K76O/ugr7QeSDZZf9BprvbCSG7UVgDLONqmGJ+PbGc5FVpcWvTnVUd5jL0OeJx7n
mr3mziShDVhoLwjIDOAehWvRv2S3FGWG2Bbi2r/k9ikcGyA+OpVVDrjHzXbycBwh
DlDWwQLnMpS5Ntqd9hCieRsN/O6OhLy42i36+K0qQFOWkSZ8e7cV+1/sd5c2dLfZ
aCJWpgIqe7mOsTKLySdYNGTP1MJMtu801B76CzJQZZsyHqTUp8orSWACwx7C/DLi
QtOAXi6TC5CpJqYiu7Egwzdkh0KSZa3U70j3maJ9h+TmQnxWWd9+EJHklLMh6U6b
iHIKZz3FrSOlF5sCJP56Vm8onYqeDayi9QA2pdDQnrUP3cCAnCALrJeCQHKCUk/R
htIV4jioPsjk/7WgmLNX7l3gSSJXrZn1qMqsew+Xr/7Gp9c4TbtmcyBNTF9s7PBr
GaW5hMjez4FB3kezHku3s8wWqBl9YCGkHzLmSxg97hGiPd8YWkUI6r4uNFnBpUTs
7EX5ro9wF3/XeUMHxtXQdn1ssf8mC4LdrWvTRxEdiPFTuA6ClU/IzB0ObFvTWCfC
7SRWszFAis0023wv/NVqqOhi+I99gurgdE3f1PlALTAWqbNphoC6S6oOyGI2Rkt9
AS/e830rqPOTqA3xkBVRKRHsOUt2tdKXIxmMnceOnbjuiKyswW2w2mAA3rMP39Gl
mXVP/S9WCS22rEjlJ6qZ9l4BgQLjgJaGIZihm/GpMr86E9Q49DOZA25Ipdip05hw
heYk3pzt40/blSTeyS8fwliZmQPqHxbTGhuTfRRgCl83+I6TSzpr2lP6c5Y5YaFB
GLczBDYkgMnGNDS//T9b2K+gBv4eg4CQ2AMjuSpLC3HeUXqgc0l7FNEStiVu9nOe
KXMVO7BCvXCKzCz2KGurNOlKioEUiIwlMlaGsWtMKVkjXbs/hgY1NVkSF5jHWrE6
a6/Y39yPh9HtTndY0dpo7km4UHC969UvFtqNdzRCyyUTObdHilk/zEEZOZhOUFUP
jrjKO4N+nXyhDdHvPVAhhRH9OTa5IDBWUOTFvf6MEI5ekaagoqmC4Dz21n7Flq0x
C7/b0AXWF3gK8jJW5ezpqg/VSKA77TO9RERe3XLV+ply4pHG1LBpeIXuyo9sGck+
8Cv4nMkR4zkveoypWT/bb+mSMjXar0Ot4ykxSWmdkmN/5gKnubLAvY7g/3CB1YyW
1BBjFWGNXSvidc+0gsYr+KMevfAnXLu2mtY3KGTwIOk5lnxGgGYqZRBRdkA3BJPN
/3ZgQ64OYZVEdwN2fxa+M4xPJFQGI/sxf3R4xkkw3bwpIqEWO5Lh4FTVXUVucudv
XiOCyQIxPwViUxNpfGTsY1Ptmr3pGPPX33wvbuma4WMpN9RkJpL2zjxc8CCiDqT6
wOyVA96T7lN1u20liji2xpqMRQLzQ0UWcq4mAixEGolbceLQDtREqGLcz1dN1YEK
gdMpfyXpGRoDsLPd51ODeiPvjEA1MGEWJ7uUdehu2LUrJGkLqNrfZ+ZTWAj03PyC
9ehWHGr6GDF5/kspk5VYTmSou3f7R/zuh4cGPHkLdctb05ZUWzUDt3KJHf0ws6gt
YubJmMbN+iSETdIbpPg0ZI1ErHKdJU4GJxuZLUDmvTzTvQoVfNIAfOVzCIXUMA8W
PGvsyWyLCSEYGVphJGmHwbMJECCJf5MWRvXdgCyFp0FnkXJH6IT0mUlzeiOUwYJ5
744rlsPoAzhHse4/VCLB1Vi6SOtVcFQ609hpy222vJbQZ0zkcPpE0uJYJg87YzYZ
+MJDghrGij9OZxVgIv1Lgr9kBSBZrduWD95BRwtxa8rDgDonb0f4g+ZIdW5+foG3
YUXfucsP4Xv3tBQRMtzv8Zdsuz/tIfr7zxoCZ/Vddrq4hm6oljymXnGTvOGR204Q
TbmRyVQc5Hcx5CIOx9XKuPEBL4lhaSwgnCrcNsKfD6fcM1L/zc/GYslk5grPuJ4S
PkZPzxszNjXiy7HJcd3mhFkLm/eIWtjBw+HgaWmlE4QuErHNIDHFbeYthG6qxp0v
Ow1mr0cYUZ7/u0RG5gZiXvU9wLenyc7oeV/HMwGYCYDZqTfhjMS63ZdG3pq/yHQ4
dqAck1S+sePyXCEIK4UeXdlKd+0RJO0ObSxbwtq9nENZyUgIo1g+TnYMFsuZ90iA
9vGBEzeSrlckYb17TOWUuI23pd5EhxPdGXnUKfwGN7FlH/+tJuA0K+zGefJFD9hm
PMp5i24K9w1oOnuRtLALMs6Xsru+bp2UbTt4rU8WhAWXga+O7HJRC8u4XNJVW4ZQ
5x1A9Nl9BDje1SfSbhY4OknOJpT51E4ySGZa3xS7pkVc+C64+lCcSCGBhUaeTrtq
1toB0I87SkEkpVr96GcLbya0c2sTFMgg3SbHMmu9ejRzaNe1I3VdHpEJkxjDzOCI
UkhS2xbGqvjpJWCk2uNDplEcT/kZEQnkkJdc3C4iTPG689XA2PW2ATTy6ylKzhBL
gd3K9NUCTjiG7WF+YUpNSAs4aNB7mAyMTtEftpOAopJdv/DTqp6B84Cqou/X7poo
aC1xonZGptsvL27hDYF/JJLVR2i5coJJf0KYczxmnpbfXf+pDvhwRRliFfJNXqXV
X9GwEkDH92abQDDnRTZ04unhCz8Ulh6C82mENMcYZqCwmD8nthY/WT/jFxwtaDc9
mrWGMG6xFU6gqmd2V1RAhCa2dbWfyrZWCD88C+llfID/tnlFdWCgH0kBwDfPBe1c
i8TgAVbN5bBLVJPIyGVvwLLSpVsNEpWU3wHUiNq+DWjN7WYq6T8Pb0jxKg69HBzk
aXCAwoKwtnjj6lGVqR+QFdvezJbBjQixtTNYeG+S0AgLnF0ZTVslPUm8J9h4GYGf
4QHeKnRUzqCAWx48pypL9asPJNrrBB8lDEUqTeX6YlE5IDONtYrhwEbTJS0R0x80
um/yytfofWGq/FNYc0tOVr5PqL9ytQMq4FqtDZc9ZbFgWY/ImwGgGLf1pV2AsPCA
NePpQ2F7tBeLkUCb8Hn5OdIexS5AgiqRsnFfBexVHN0xRdhlHyprZy5pAth03v8w
yjD4cDJKGPeYcJA0xulpAsgKrVXWsqoqWg3QLyPEFXwf1GIUuiwuT7rdQZzN9l3D
1y5BL2VizbtAWIcdNtFahd0Fs2h0E7P1lr0lQ5NxzJ2nA6sAQ90z103krRqlBsoN
HB2+VI4wj6m/mr8rwVqUFK2nxSQEaWM/lkQBosCK6vFxyG9Rg+OA5ZcZ/Xd53vZr
Vc1hQdwviCNx5BpdfBQI3Qz3ySn3a3NsW0+YUIjeusHmlUQjj5iinlbeovFo4WNA
8EgyTM524xf3gwFI4mbu4xLigN17G4h9dHG026qPvxBtSajYUbFDf5V9UtItjRnw
lLKz0BwYeG0IFeWe07H9TNSP70SMdJ0IwXQkn58RFPscUplPn9E8eDa3MPiZLFwv
oE+OKWE9ypV+utsg888xQ9vDuIVWkzrN6u9Up5hRIzW/Ew1uLlJLgAaMR0QIXr9a
rF0uLYiY7PWjWf3gKMbNmOrUVndhfhb2JjELJ1L2oWNdLPJx9kBGFFCr+FqaowZT
wLaOs7FyxsOg+nkcVsjRHHfV0OlmoF8jkAkvh7UrFCXlperrg8mLArFO4cM6Fd5P
zi7LZ9DPrup/MetfaE8J9QlTKdLjONsvYonR5MNaMe4gaFbhlluaS2B73THb82Gw
1fbypfo+jT+4Xukf+T0NaZqARovlpkoYK6UsjyeS+svG8WXDqaIw5X8H6VhcA3lI
AOSXugpho1vohWKZE5cox4SlddPMB5DrtUmSwadlzu7Fv/3xVdZ9Xr0wgG7DQuy+
jOIVvoK4ceaDjazxlViOo96c1TA1kXMGm1W2nV1MWlB30qa/7GAvbmPO94sQqqLK
1qnRNkEdnOgctehB5lI4VCtDoKQD6Sjf2uL7ViIq1fmdxonxsbxVrCCNdZ18mwsA
dIxvAQNy+SGZwoQh6puipPnwU7zzMazfZsbJrEAujZb9CgYnGyGzZukfUwEcETvd
Wfs7jsYsKXdyJfO8qaszK9/foloZN2jqmFqR+ykNg/BG+BJiLaQXiRBBXUov++o1
81nY2d4pbUGhEN+XDf3zek8S6TGMmOyBGSpkFKKC6i7M0MB9GOv2myPdYMZdgJFN
h7rm7N/AZdvnn180Np2xXaOh7q5/BPgRyx6KQJGeL58JtY3EHtGhrs7ZivHLD8pi
5opaku6UrUrjSnYaPMSaSrRZYK1y18WKr3+g/XufnDd0uLJ0BYtNSjpCjrVoAadH
88eb2RM0xjIsDzfMy+VVaF2UUvfJUViW39RuK2E9jaZE+czXV/dtmMq1tLMwIsK4
+5rr9MClpgkdP/3Xj+sgEF8rnUm6/sCmp4LJp/JyhvBHmm7PCcd7pl49Zdyk2Ieq
QWoF4fmvTHANlYHitymdHG+RphgDaNPf3q+a7zrQhJNmi4SySHf8uN5DHOqgD+VH
p0BSZdho87bfWykT9sSLbDqqK4CfdsjWDRMv4YOS8EkzrG+EAwk/g+C+kn0K218x
HBc92IjHQ7X0iKnjlMftnme7otmwNLjXCOffiCiClyqrptN4c9JBbCQgA0GqJrnl
68GPwUCjKxol22L02ahiNJmHfJ38ycnRgoxGTCmzmOUzrHlOdj/DeMbs/YVR6pd6
5XF4us+23Q2bidoGr8a3tWFK1tIinnEa99wJRORJZeCgG5PqTzT8+IFcWvmZaaZR
9YBu+b8kKjI9gGgVL9zMF9U6dpFsDWzTdz1YdPCK7vx1+pUZ2nO/ABQuf5lIH5iv
T3anAPk6LSGySwWNSa4/giLkAGpntg1p+WmuBpOmTRtCKcjhMpyRruWomZK92chc
/PX4HnPf7HgHiAOn0gsc1I0UlSl/TGB2b+/oJmaOCs+GP+eLsY3mQ1pgutYZHnBv
KLOHO8xcrkNuhBJeAImKJCPKzOWuiPZLK1kl//UAFgPdjTIk5IkNgVz+ZFwOI0er
hIcoz3LbEOB585YlCaRsYlOFgzI+hLKgnNTqVhu1Hce5il+cIsgCmf7hd31gNtU9
I0pDrh13r1fSZEZUgMr4KlXpSeJJS1nO7UzDutGo+KrGWUQjBM0/TE5HtBvkWVrV
ePWpOlZ4QNBfIJA0T56aQrF4mElz03h5W6vwFwteahyB6NOdnkhL8MmLohCpBWph
lJxvNl4jjZo0aBKS/8yZHpJL9pZXg6jk8PiNYzyI8j7bowCPnBtUURgdRo5hlcXl
jot3OcABDt6sepT2yrIK6296EoT3oFGKM0uP00bNrJI49DINeYtFcRxUJG9QFvMn
7B64cu/FyaBEwv5vlx8f1ZQeywqeiITPbwNF72MOEzKgbJ+6wGlt3ebfhcxwRTCL
r7eOZSws7KLF3ps5zeFIK5tPWcIrcjqTgSjZ9xZdvZujVNwKVJhbyIt9jKYT7x/m
5Jvzb6AgEchA07gpbR+2sQvxX35kPwTShEX0YbItsosZ9xzEY/hZTdf3EtjQ9Y6K
izJbi0HlOv1QaurSY8nXZ+sE454SwssFP/aj7RYAsLfE1aHHbmnr2+9lco3ewfil
vCZxMYUh3SsMtbmRi8bkWJiqXeK9jkmvsD5MnBodtUckcNz00lssVHtLWMPZzwoc
Iei/06Arnn3TD+kcf3i1huLrDOwVkJpE308JOfLldiGUgZcFFJckg4CmeDUHcwya
atku5cOVavz+p6dd+FrTjVVy3n0JqYhUsiQo1cxsQrWLWg1H9oiJRHfKbp2bRicd
a/jN3aCXn8aZJWaM+JkIPNv/tFrzk1E7uVgwrBsvpsBg7z5fMEHq++NUReDOUgAh
14ee68rLVwCjOlq2w2fXRm3YnWnnCCVRpaQUHuaJITvVlEfZjV4oCoBSfgTdkR+q
NWzpIPLIOlvlmQIdcg6Z0tY5f2FgSGN+ecuLWQLr7KaIZzdmuwvWgIrHUZ/YAQeF
eKtO9yxlZvvhkjSL8LBkEr9CKQh4kjyN4byCe8zT19EdBjDFFJxHSfBPlC8lBqdP
Klki+eCxhTnmbvqnsFNQVoYEBS9leY2xk46M2c2DIZp/otpSyKFPgZ7iQCvlqreX
lFLXDs0LcxIssSh/2okfrlkWK2lnTs8U0ymVq0nztkx+9Qs++pwuik2dxN1DbSX9
MCWiJ5r+ZiTKNdS9wb1/fgi4um5dmt4huD/35RvB8s4vqtDf3juUrVUjGyaF1/sL
I5Renn4K/HvbFAGGgogX9eh8pgNZhbArFThsdyd94/G/aTwQoVxZ53SEA1BANiuZ
2z9pUBhtD55g7zt77q7fcpwqRWvMXSzgS3sAmdF1BW2Ix8UI6v7LDx50ojnpplLn
Yosd1nEjmpWf8ZfAdHrwN2EMOMPR9RaaHXQ2jBEgC+QOpUOXZSMdGymGABJxf08o
jFdAvjGtYtfUB19NDpa/Imf5+yp4QEYmOxR+vWUu+o96MOqOfzUIdgd9roO84ZFc
7YHqvRzHdp7rzJSrTVfrm5JiAmJaBUXB8krJseNnDFZpO50TcBtovNL7i1wcpvjz
otbCPbNcifIShZm9jlOnNB9aqaHzxIq/wJRIAl7mG9J2feTM3yENhj+7jA4Y8NrX
T/S9Mth3wabZ00RbHgUNcVYMR9GTkUQV3O3iaxgmq8kvoka3CGj50jOzfn6wgZVo
RSCJbu2BPVcY3JqeqN/Rs9ZwXsCwjA2s2y+nrxOC2CgN+q9IVnB7tZjGT2FQGcoe
Sb6wDSMbSym1Q1j08h90S/xEXKfYvhwheJAUr1m0eVuX+2anVvxS0eMpjoFK5nbv
xEK/wDw457/phLK+oct5MBRXdAMmXn1oPWlzXeGrx3VJk4WQiLP2aTG6XvYQmfVk
F73itWkOYbqqnyxfqzmn6w7cg6wuq+fLoiFMGut9VeWPDy9Gn8MtCuWp2JB/Qjqa
I9It+GHvfnmeouh+6K4D7AKyttsHz21ycGrvuWgFubnYuAk3AnumW0G8AqzATTqg
Io5hzM7gfiviMOD42Gxs0athXO9c7BfKMhGb0hR0OtvyXSFg2vkiw7Ni/+1zolly
Mzroa1WnAaUFZbwyMVdO+r3mxxvrw5/52Av7TqL0cx7yQlWqS6HfOH40WrVaYOMm
EF5U6+81sBwlM17I6ih4KtJpFlJNwBZlGiRw5WzGMmX4Uh5qw+jJvJc2c7aekeeP
P2RPPzxJ7QfnBX3LkW7DmC0xWvLpzgDxY30e2BsnWpXvLNAJBagMaL5UfZgmb5so
SojHGiAs8nnIYszQRrLNauVxKphaK4dSj41oQyIlpP7N462h7K7iVxx94I1/MuWH
0MxT0hTar1yKHmLmPd1A+FvMXDwza8NJJHmhvji3+Layue7a+0GBdtp039p59cdn
CGt9L/KFOCeFx/WFLUpe2I9VEBz9Rshn6nxTi3GrmA2sVzgPa4J617uT1AOzu7ri
lvHPZO0TSeF3x+B+Pf8cZCjnRl/ebojMSB2kh3Wce1efnvitJGr9fOC2f+i6+r8U
fImmp8YfR+3wffvBn/XDA4pzUXMNeDINdloPvkfnZNc2FHdlB9J9nsgt0llzGGeF
PFgf1uBymFcy4X6JnFjjuB8sgw4YGFrGxsy5Gv8WzsZpI6WcskunLc8HFrte3nM1
T02tcruUtZ9v0uNpXPbz3pp5gxWcmGrtFfsFwqmcNb9aazfvwVGveNhWaAeOHXNh
qEf5G9toUm5aEjD6IaGKhiDXE9gdaF/jGz9XVepJi/1whT8cU5jjA4ps4yc9tGvC
2FLnBFzFnwxBuEJZ8mu5qEn55V4WgWFqFZsoxmffhiqywBQb1Oqtcicm21cD7G4I
PdcjFx5F2n+Vos7kSLHlFWnlqhqaIrZ062eQK6Oj7WEfiCZDyYzqKp5d+XYzt+fF
TdIdb6wXNgRVbrkV7H/rWy5swvQgghHCzQcrBlicddDedeFuB5Hheby5fHfD3TJX
RwPaVOFCIg66tuFSE7p96cXZQflQxIgx4J1rMXO8+WV69FXQUqan8zkZ9sQ+cd4+
1tbOjUC8SzoMy4qbGxwkRcSkSy3aDvuLPrKSUyl3eCP/eNoq26cJY4spZ3GdmfxX
Bh3HPHUVqqAHq6rIk961SfJ8p+e9gLA8tsxAdb53D9xtsL3TYXcYNAyyLqbFUVXw
WGB9u68ZauBlmsAXeE+ElumivbZ4NnLpSrTS1I8wqxgzAWn2YZhwdbd1bKfWIaKl
1HyvVa/kc6XpKA/EnWk5gF2vEI2Jwqf4LIcaDeY98QZYIR1KRqnw1zlM3CEL83Tp
q/a+JV4x0402u5xNdP+iaL7Hppp/IUef5CUjVbrN7GP8iXZCSCzYUaH8gzy/Dy35
ZDNOAFDwwnHl1AHnokwrwA8MVr/PDPqJ7DJoDg/mZulIBzKWPrPQz56AHEbatVYl
n9hwJYnB2dkUi0ORocmNfCnqWukkVzZd4AVa9jAIwQHf7i2WLsJDaR3IwTsUx2i0
pe5Ea0eWKFtU/FiYfha189GUfUm8PwFPGxXLpTLXGMfO2nprtadWmd1us5jUTjYQ
ShsMNlH7Hk9aXPUoOO6QAYZbH36YM1s591R7D+5VWJAq+YqxwPU8DDbdRbT4Y9fL
Oqe4RnKKFPJeVveLjvF5ErVPDphZuAdmsYEBiivvTzXxSBsrQdlp59jlVXhd2SQK
9DEmvNFJdIPYOxPA6CYu5htCi+fs0kFvyk0YxUcllf4GFRptR2bAoDphBy9Y8WDj
x9y0OQ1voBCyXFl3hNqmNfPqXVTupbc7cb1P05Ypki0EAG0vvpDyVdc6tVqH0Pnp
hWwo6xSmjzyj4Mse4/HdDvb9Eka+bEm8q3jV4cdlehvb9HFzNG+h+TtAATN1c88R
4hmkWLva+bBHeOM5sytLrLlV5YApmbYH96N2CZHxcXI9etunOCc7hEmuZjOU8XLu
EkegHpFM4Iz7Vkg0sGFHPi5jAnLmhy9esAezeY7RBUabQ2sFDw8Cr7TL22CbZDBn
XV4jPSGVSGJBuG/YfE00oi+UfQJLESm7GaNAZS+gNVSmwxa2Uz+dtP7IwFGTB2tq
DYfvjn0TDe8EkAbDGYiQ/aYX2ooqHeHUpnPLpkKKwmTBTZca3A2jB6poKX6XUN1Q
8tepyLW2MzDEv8DGdB2yeSotny7tdUdstn4LXEGcMJavz8bZSxzMWmhHYWaKLxBP
SHpG62t1KfADsPGOPT/d+nX5YzIUjUmxyYU8jPeWYWG6pM4Sr5eLPoFKzk8RxBVw
mR1eUeND2jX3E7lTrzQo28aWgFDdJmPArO7jCnicp6WXWLvMONKdu/wG88rWmIPH
dUZ2ySxZ9hCeZFgh+QCStnXDhbvuNf2xWJwAOLwq+K8OyFxu7EXP1rHcmpnr9B8b
0/ekdPgPHkyE8hf80PCBadi4RYLx4B5ZBE2FvJ+nudXsiVqO0p9cYXasJA5PVhhj
nbtI+YZTirVW5u5QSg6VYI7uK8ofNu8mcILwC4XQfGNrB2D2976bjWXEplUadq6L
7AzyDdPqFPCjpHJkDfBI+L3BeA0rOdvOqwi2nTYBz6HGzEt+Nlmd1FD4P2XPeO7A
Vt2qoXuv0y/jhXzFMalGxnOhoxKpPvGcfrBSc9oL1qYZaXfTfXswfJ64dES2wIUt
J3pFz4FTZIRyw1JbCZOo+Ky9lJo6BSwUatjE2kagYmkjCEPwPYSQ/jlnqLLsxqBI
d63OVLbp4adlthPw/3ukoaHaY4YIOUZcXho3wq0LyqsovQZJN/Z5J7lWKdLMjWXl
wwirMn5pqmjRzNqix026fo6STIdQHMbPLFrg7i2U43r/J0E2PjiEdRu4zqEha4uC
VCW72tBkqnhl9uK2RupSInAr5vhQ0axmvPXbPOp0ubZW1XiJCBf292pFoaOfbzzP
IY+SxWjN2d95dpMDOg0EnwVq1/W6oL9XnZATlm7xA2G/vS0uq3/Ro1JhXf87c2S6
0xExZ4OAaXZC0v9YCAF1zWl6nccivmLBhITef+76Be/rIqWNhJsAchfRFIvU3Pf/
+OBj6VmCIR41+3lVHF3igy0LgrMQ1H0KPaj1MsWJJEr0DUFV1Iol0rA2VgfLjLIc
68ZcRR0zW4RYzfehV0naRpa0pM+34uTKOLn/qpNsFRSSWbakUHrwGi3gnr51aBw5
qQJHcSEph83mtdiZfTpjCx+dwE2sb9GoS682FOfWk2nTFimhcWFINyhPYSiyR5vn
p+CN6A78YMoiWBq7J6U+brnKlz1/fAeeajK+kmog6Qv0DP0S7L//2Gbf44U4wooZ
BVxA8JUWwC2NyL1qFZiM3am2zA/XH29s9guPwoCgh2zY7yZXYvMV5tRTdAEe/5Mi
YHh1C/vAB06fFlHeqc+vq++g6CXzvkkGekuw8N2sRb9ourQ9768rddLAkDvG+mUz
U5pJlOJK3V4gAsJY3jgE9z66AbpFh8xLHqJUMjbc2hfPsFBZrm2z3HxHdq+JEPF1
UO9IGyCQflI1gunDOT7LyfCl3kVhQCETmdMJDkRQeUXK3IZBIHN+2ecfo4cxy9Vj
QZ76jMzrDVfTtJEbAqVwK5cgjihWJDPhfgG8isvmGF4DtHXtxQtMF+dmH41E0Xo2
MKCM4d2qvyOWdiFHxDy0jFkbCPutjDhpLBQQwc694UD5ZPULBwXbg2hl8eZ/zh7q
ZjVX2I20m3H83SrDMSt94cXbO1FGYbjBkvcPrOm8kEdj4fO5/ZEbentmh3E/cT7a
F/OhlOrGl6UJJ2cW0hi48rJ+QmEXE+hTjEOpnX7mJ9lEqvOlz6mSy7NkPfBEzddh
4713qHa3PgCgnjphUe8WMqIP/rc3N5oItHqapb9Fk/lxx+ra2RjrSTZQym2kYvMI
ScLMYWS7INh9HAyKLzmXGIARwIeYlN3yjFPfDgrF6QjsEAhJ6x25B0qRmrdYe1o+
8ehmlt+CUn9hfRcYcgfk1RktB0okP7AcAJn+ZXe8t/VzNmE+49PRTQz2sVk826pG
jA/29BSVI1n8t7egojYGfDAw3hWExEJ/lcpgqUV6fx49ukddbRUnR9qgY+bXCBx2
G2BaDHn3m/2goDFExUd5CarnjH609ADwx3RPQ26aV623OBMeC/rvlTVMkxZReQIm
lMtNxgE2XbkyV7skhJcOdDWBInGi09uXyhFuXAupaC2UI4eORGkK8Qz/9RLEYhVA
P7O0b1FGk6PqoCucHBaJ2N+C0RvVACnFoH27a0qRjrgo2ofy34qvXNVAvXEyOTt2
eTELan3pfyaJXpYUqsbh+1m+PK1Eyo0pBnVtwlm+sY5zF6V8s9thO/pALD6OQwrK
thoss0TqE7t74UKWRsr8iv2gLrtI4eypt4zTTuX8cwSYD0yp8ye0YxaSQWcTvJ0u
0j4sGF5IDc0SFdBXiKTEV6gCwI5V8OLnL4UwJXLCbsnfgpOvM/eJtEYwtnRlLgS6
g7mSIfCOBMNNBsISEvNjsNcvGp/3DGwbzIButnlOceSJdTE5LUKKdJ0gh+pA+Pos
ODgmbknBBQAPqHjTFv1gsQ0jwY20OvrvI24lHr2RiEQ77tVVw0c6vgU98cGAhgC0
rNuHRZQRZwge2zrPYQBgKLngcVTzHlqOmEZdUqNB713Nv0t0eWQiKrTqfakCMyNK
beneBiu3lAi1veyYUIIWzWgVebAGylz2ff99RB9+eK2z+twIKiOjYc+w/VFxNg/y
ff1hkZrm8SxriaEdvYdJEMm2SpHdyhpehvy/paCNPCsjF/R0Bu8PczeZ+Bhm93sP
ZL50nYI5tTVyE/ztzt4972dpiscvUx8bpknyDapBFnwGUrlGyX3zq0m/dE3HoBeJ
u0bMzFoDOlUOiM1JHhFv+oXqlQNJNAYxZG1vq3AMauWEkcmQ+0GiFcri2hrFFmM/
jAccIIJMnopyDGtD2KKKoN6p0P1LrS5MaNeMoNi+aw0kUU2966mXGbFvUeqnjiBv
C+aMjcNmzRQwBvLAxGW9V28JWluOSqNlXB/uZSlfk++i22QDjhGqMPJhjw2DRdPg
qRtEefHtJeYihXZ2C89/RhhQ8Pn1JufdsXIczMZjjvC66pwI70rFqPL4hmo93yne
9FmgigpuJkMA0dszVxh/rLIfYtaImWu1j8iQ3DHxcX+PjeZ5PI4Lsp5w9EtGMtxI
h98HfWjlQEwv1Ihte3sRuZl746KqREFQR4jfDmmJcWpIC4EPG2Ckcadht+L5/sst
PQFTCKtlNADQZvpn246VJdRfgeR6Aub2UdUedUtnBCdzmjkvjOqDzOPyRxCbsTn8
+sOAthwC3sOBHgBSFeJHK7qebMn01Fc7VfnLCVX1NQBgWz/cyHZb3tfp9+5uNJGO
W6/ML/ALLBAhEu9b0ZHcpsBzxJ7xY00SCwtWC2u6TXST3hNZeUNMPpV+yo5MuSvc
cjsNRH3YEd/0ok/5/yx3kxSOCAEtj4y22vgzs+zZIZWepr2qLcIYQVsWxkTLB28y
XVI0Xi2/kr2mfWVZPZ5fu3vrS37KSrik0LzzT56rWUItoTJHRshmRErhl5vZ63iS
3meH3o9G/jTKq39HxEgtx7qGn5X0yjU6lD4h6csTwDD+C05gGuDDtAEwdBvlVC8+
zymyZtshGRsDjR/SREm1zfZdoxoSI/KdzotlPpaiFpuEdVlF+kQFHCxeJK5y7zX3
OQXmSqaBotxzs1wylyFL/qOM58QoG1xOBzou/draW37zf/Dqjl5w2eZX6FYPS0m2
A5Ca5HInN+O/vbt3HNUEJOpsSRb3DV4YsLjyTPADRQji1Q2Dog6mgOyglawTPvnM
AGsTsAonjddin2KCpQMrU7QfxemjLUyqvbx8HCxUNRZSDLbxfGot4SucEFZHZo5b
Bek+m5Om8INMrbCsuOZv6mtZ9gpEoR6vLgUJt08lz8EgoRJTcaxXBfBAO6K6QlT+
ecbifXuUESlcVWNzSFI1Y7epn1W4a6NOAKPkP+jno4msgwWSrm+2kDNyaEezUaPK
odw3Rc/GYZcUfO+RiJa6M1RJfTfazlUYPzFFrie0iTM1RyKlaTChaGdGFSKiyJ9t
fAdbpVXA7OguuHyQJtQJaVDOvSPgREmgAZZwHIIouUvDyIwJ27daOfgaiQogQIUO
SB2G72pEsYN/Mrvl2caxbd/gjUEuNGzA+eCBFyDGJkmjlgxeX+JAgqEoozH5S2qF
GsmAgx4HMFKuaqeuMlBaAkBr7E7+ZhbCJRSY/ZmPQOVIH7VAh9VBZW2CC16EG+qm
xgmmpfLvDq08Ws74jm1wE+AiO+N1SYXIj6Jhc92VEDspRYt0IsTG+eEtU59uVf5w
aMHxQ/jRhff+V4DeeYHxAurKRCON5G6mBuRcakbx+igJoCBCyUXaIncJsg0Fq1Ru
2wwT5EcvNfngVlpxy24kBdcQSZ3Z6ta1EVwj/yAhAI2Fbb4KqLyaO/ST4F/nJ892
bVXjRUCyjbrUMbJ0QzPWZRWxrolH4Ic76md5ZVF6tmap7Pdn8H8Fk+c7+RoysHHO
m69AGLON/sdF3DDoUQaY76U0kUM2GIxNiDsJgGiLAFfwmRw8SQBiRNNqoRG0+IwI
L2nEcIO201vnvF0N5tQiOc9nB+lbhKI4UIwqgeCJLJQaCP5VsVY1p0AVfnSkV85s
fnPcMo2Ym/gsNYHasXlroKy9fL/qkRY0ZefE0R5hQ315eJ16tIQgJm6SAijCroP4
MF7oClbJv35/fdwc5pOzXCAW8o1NSkiTONQL5tvu82GWRAK+DshdkcWu6KiLc8J4
DOragL9eTRQG4KCJKI5732DEp760X0ALuvxGmYhFqJ/lDrxZO3bYMxGym0MuZ9Zn
dUwxFVQ2+OUVsakWp+oUgdjfOfhyxcjB5Un7cDL9zktoIQTb63B8msF5tr7AeqJS
8Reqp0JkrIlJjdiW3PA7mVstMryqiNGn3eT6+hFv759qrI4wJuEmezC29YZpm4Uc
4WPf5eP/1hQ2NzCoipZHVh6thTG41tIudRjMgABEi9fyAqXJxUGKDOMR+NE6DUs5
ddlsW9F6Mt0Tjp6qiwfaiIw4dZmz25uQzo14yLk3APVHcNmXCOh1lKEtJKT8H+JN
xZxSaSvKJmqD45TbRkFgSQNnJmjFfDi5eoVaXyWVghg12kUhIsAZuUEOHk+xupnp
03HNTGVrAqy5n4uF/Alm90eWFNU0Ch9xypKRiOerdFEgkZ3W2JNUfA2sCLOaSQS5
0Bm+d9ePa8iNJmazuM7rd+P8eIhSLL8uJXg9HAD4zzIumcxmdOod7n4JprcMB0R7
huAHs81S4TQM5Cs2y1JW2kBHohXfh4LAWwgM8JOgGPLlx7wzY9y9NfK4BlLqmigF
jiCULNaO5H108u7x7d/CSBafCwqOYgbENTywhsGobHkj/QNGbOFNY3u9FRcjMzeC
qJHigLmdaKvBVATGAFniR2wRthFkNAI5t/neTNEuJ2xRMk1HHunBO5xKqVC3Sh7Y
WjDHGYDKK7WcDEKI8a/GQwbEE60zrwGBhIzwVd0yy1aHzgK3Ip54uEUP1aCBfexV
His+RE54vWhDKqARr3dRsVQXvWJAcqYk+e/cSpjvi7ptCGoXARckd2xAx2iddQkh
IcYUc3G8G3Jr2zowq5Hf/wGiBQxnOFssYNPYp9dTF6fBxGxpDhGlU2Mc957UkcXY
S3Pw+4V/R4+vHd1Ak7i3kDELl/kWPTRcF/CO+34A9OA5fPjHc9JTr3yaR210F8G0
0VZnb+T+Us66gSLG67fMADC6DYAnnwPjEEVgw7f6vUr7CLzTD1Prdn2iWuYUgEWV
xhdhZjkh9D3Kj1b+ECL5bz9uX5t9+deZMH39XNU3pZ9yaA73Db/9cl3fIk3YaQ8S
eTCwswNzkpcS04Ldz7DSfMIq9uqHHscyk1lggcht8H3qyrH4PHVM/BYU3KbRo+A3
1hnbadkyz9e+A0EJLGzwqNF2PjmKPBtYpMLTFXXb7srRx3mlsTCED2Y9LBex+z9q
YMkNXYM8GqwaH3ZyNcKgrD+1b9YEFPha7X9BR/wKh1/WDE9rtghWmzhLmRRghEs4
lzdF2CFwdTN1CRBfzdMWrzbE0bxzKqZaQQjNm/7n/ZwB/KEm3yWvMPOVc26mLb2S
fid14SSofqS+xvDYmsA9h3+LoGSowfzrACDaYWx5fcbEk31B05TJF+ViOm5LrovX
oF63CgyU4Agke4PiobeVeglpxhFcp9YwLPFsxGO/N7mlnyrwXQvmADGEDj8Mg4Hj
n8HwkI5YRKFN3xZleJrI6LFXDbT7+b+j3i/703PH5xdyniRxhgvmgyIodt+kkMhy
fwjfS3cuPHtdsw3W6n5MrrT+giQvvQmN0Pqzcz5fbuve0Ckle4jBluzuXUHMpI9i
UzrWP2KzXe2FecXIl6BjNvunlQpJNEJMPezJUigl3HFK5zREJUeOxVH7xN9YtWBe
uYqxyw/dLmfCDgTGX9xY6juj4Xv5dsVpEwfroTYp/D01eBpmVy21JOihduOAoVbM
xYb71iNp+n+JDGAM1nQ6EjOZMSBgoHKEDRJ2oFHxJUNMrdGnGD+lY9Wy8hYX269e
qmWxG5b0Qmm84E4KyP24rAaiN/WlAtI1xbCnJbADxfC7HGCl2UWJilEvoVsS6u3o
hRTGwFXNkVW71qDX8jBfA4hSkHBdl3ZiWA3iTnjHNpsYpzdqD3HAzWGSG2eDDWq1
NQJ8nljWtfxXOYQYNpKhPKVKjrmIdrNi43V5p9SZHpihgXfyhAueK/DRBKNQIoBk
5RbcQn3Xv93dpWJypvHqpYN77A9GC4GRlk6m4fyQfEyIfpffl+FLewb6Yqr1SdV8
HSaxDR6UaUUN4dfVECuu8Q0h2WAfG/N4OvSzrAdYilCR3wbWrK1h8MEBrbLq4cGc
+/9cO6JZNBJV8+YflO467b25ChQjoHa6NVIVTpeF6TaJDQpROxR75t3lSrwKyh1/
aYVO49eN0ZLGeQo04P0ft1axVl9Xz9KX1hq7zBzZxE2vtLEd/YHR422sGntnKA1j
bZ80KK4XAoUERvpKy6DuHdcYgfeh9TgzuusBlMiQpgaLAM0BW6Lio7J/rZB5bnuX
Yf2mQnDSP92k66aZD/1Phf2R28mvfP6ZwAqdwwRJU+JLeuFMhGd62Wvl5eXq+9Ud
f6g7/iZ5z2Q6EUzxXTvinKt5BqOwRDM/hKrfBtJz0KyvudXer5PovYlt1Z4KBFrV
+Fp2le3bzIBEm+/2leVhu0prR7SRzm9UBPPoGY/SDpJzzEfghehd6QpHK3ovInqf
ivzlIpemtoFI6oRHsabn8SSTqbIR/QSAa8qwqfnDpHv2jtR+KYBpt9HxGMyYZZe9
KRuqJvZ787NbNPYZgKO0oMI8j55A7+WFCCgApX9XPk21V1dJUZDzrHWjBOlmMLLb
Inj3QK5HG9f16d9pfntwMv1YJlTEVkV/gyCqKosqfDL+ioGqTETXy8aYc8AVpaYr
nQ1jKJ+O9+/pwWNtD9pG/R8ezIL20eWcLtQ2V6r/2Lp4gdyp3n2RvZcq7uhXxQn4
CzkHBVa631b9XTPMhkENtMSm02GwzIxowTZ9ZjqUuY5nY2J/edain/CFBYjiy99q
Sm7WMPJe81KMuQcIQxxJGzKk2vurCnMzxHfdvavrHTOx6jmzqvwcWfHE68TPqMvb
acS3X2gs6tKqnZFdszyID06Kuo773QBcb7nqCUVylML+oV0Bz4zJw/bAHLowlFfr
e/Rz24PT+4f9QcB3EJiTshX4e+tlpsREiXwTg7W2A05sbr/8lM3jLxCqhetTJGEE
cIzNXN3Th2ilwQBHrBRHAe1KkeB944+30zV3mk3be4nmdy8+jXJ5j63d2bRA6Jif
cVqt5g/LI6jQSyj4eoE73XMb3SbH34LukKPyC4D256StfONvNyTsAGRxgWTfLxxk
lJG3T1oFYN6sYNp2W96ZR1Bn1O48dQUp4noqhpMlP4gRDDxn0E5a1OTz5vS+eXn6
M/9xbFbk9TcXsbObOFCtMZBGQberVvhXfusv3t1GZPHHx1eWinoZHVTfPvzWjkD1
Q/lETV4mXJoIwl7zkEHdLmgR3JKyM6mejQF2QJbj35VL+Ma0KkoIQX/812lW2Bfh
/W6myv5AA8WpcmxNX/C8CIri0kkqaQIJwjkTjz8tcDfnMRGgMSFX8ptQaIOwC+7C
GeN4ic+3doXBaqoV2pF/so6g1s9FmgtT/wkGh1XK2DPjIhDYb6/5FLuLb2IlMvSx
fE1lG95a5dAJoyZIa1e916x/n6DgXrF+dSnedB67bIdWpBiGRKSyUX7GIJPSMnqo
MLckv/aUhLLeKUBDTMr2TF9KiofxgZI2Yzg2pFrsQJmxCgFSkGz3oTrzU8tG0nCL
J+96wQy1ihFGbwS+5Aw3nrh6PJGHOeLzN/T78HeY1rdIrnmFqJbb6VPag1LLquLH
geu1pEMu8xcOQaNOvIh/Wne8m2XI8+LH68PP8VJ5cB/KUod+Iqat44F3fuZkwsbq
S+JQeODemA1ttx9FtSiRS2kYMwYPZlF8qRrLbKI37wXFU/8Wai01Ek5oMb7lsH8z
8ehzYqCV+qDGgKg/wEBt1vADJMhP2u/M+Za+WqmtpSp2g57Re+zpurfoOHW0KJcu
sd+3nm+q4Tj3/KRoxPMWH96Qh792WwrZ9121gSsxfmrm0FVsw/Da0b1SVRMjIKdx
8ARhFTPMrJ/v54SAZQTCdCevHBOdUE48DfZmKpvy29fmXy8tFd6ACq+ep9xqcn4/
RMsYlevZIYmKfJ8Us/RiqLdZQ83O05EnpYCDk0LtAZwIrT6nvjiO4nt2dfLY1IiV
TnqnL8yPbt8xsIl0jut7lzHQL8lGzOay09kZkUui63AdmExAu0lhG/nZyY+w1KaT
ipoc1pdTKvU2AOTduxHW/IO/KKY9pnWQ7Y1m8c3wM6So+jcHO7ZtcDzs9PYc1+MY
YgFglcwMnxwucXzFHaZ5wXG4LVi9M9Qo5U93GniO+TDjOvjkkCluXjENSnPnHpUK
9UkvBGEYYJpuhQp6XVjoYTPqjsmW/s4UE1T/wXIYUsvdQ+UZRYegC2IDZY+gX4Wi
PSy5Ps/M5UAcSgFfNoiaWMwJjsJltKbTsesUA+4Yq7iu4rcnFPtQ1PqBS3Oq+EFb
YExas8t7absuSN1nfLdkI9ifg22ZbkjTPpYUiZQg59KV2IOqG/ntM3E+wtddCpUP
BnpkQ3YeuVobbqbDDB3lECxcxtNBnEHRGsbKoWTIZ2BAC4tXAJ2Wfa7nm24UcuL1
XPNqunkhgpAIJtWxsj6t6nf/pGb7LzP/1SQg7R/iLE6eUhJYYi5tiJGcVcPySPZd
puoSfeowmuh3Qw3sxEmXShbe7BtGLVHZZoAYQspaHnkf3pppJZoajLU0PYfzie0X
Ca0wuemCW1zZ1NBeIsYJAv0U5JirFroG5dYH48KTaBHTPCRoN3XuuEqjFg3YRdN1
93mkMZDwkhZs5K8ASZwU24c6IaU3sVrsCAyiUJH7mVcPvncMWr+8VJOTVbJP7Wjm
5pdAL1UdA23oa+PqJq6xnM/QsJq5WARt2g7IvDzQUJtqFhi4cN5xotDLBZQ1AjZ6
c2bTe3orCE3FLHQspicb+PRrN1WH/nFdyWyzHj+lCWT52cRzUXEj66cmdZBdsdIY
3xf2u+Yp5tFRhzZFhl5Za8rZhPF4X/Ig7pVFkYvCIL+SSlhH8nrff0BsRFtZdDEq
dRbXlkpG6gD7XZCv748qWSniid6F30Baqj4d2zWugU1qDSfdfc+DTADoYeJfglft
ZDs54m48XhNVze3XgXEJ2b24Xq/f10tO42UIkLejL9Xz3lJQY/eyrHWa0gGtjNci
KCGXs0WYbXvdwkhe/LpCV/mDB6P3MkwrkoAPZZ0hVY2N4iJLpdsZA8VWEy0pckH0
BJf9DZnjllUSjsOoHWqAFoBTngW+7+QbllsccdKj91/NlHCuzyHNrPiuAGXg/tY3
5Bhffn2qzptofmMdqiBeLwPwObgFVi6U7XF93sOhV9DpeDjy/Xkzcmt1RLEBXG+I
citSlG4FVgzN4IlJ4Rc1liTAzsqMQYwTi/tOh2ibwPeTgJu2j/PJxTToxsZhIbZm
xJFSs+2bczXKKCtdYNs6LPf0t9BBIMxajAszz21oghnWR3201u4b/sXooUEpefQu
QhJbHjLjEzEpoKy2HEqxIEG02RZ0t6+rtIBl/go9pkzNFbMNdOPHvZLlFYJMiMg0
a8cJxGrj+BNW0duYFp/yKSCcWa71RgDQd9aBQV1egjN3wwt5o0LW53PQbRo/f3oa
d/HNAwwjzSYrkyG1T/+xGTUA21YG177555POJl1uJxBjGM+1O+dKR+S+awYzgr9I
+PibgUvnd3Bzbv8qdvym5zcqWIdsg9QoTvyCKg5nZlgFofApaRAXJqtpPC0V0FNf
LojEU56j1oI5z2d2uqEVEpoYXDjfx63OnqWKnppFNnpr21otQ0g0eu51HD3x6KoT
XhmcVi8ejLaEMT8I38YRTIrzh74vFKEH+TYe/KmYPdm7hPueoxUWG1eijhkA0RoZ
D7vQVyyO5Lexlg5erRZUqcRVes6UrhpJ1vccycyhfORmRBGsCffwiVMToGpJHbkP
7B/I1/IhdPsTdEHLNxxH1sZSS6MSGl9BizRzBfLOIV3gztmab0EIJg+mMLoRgVST
QxiXw8RsozvJKhSN7/2A6iI8jGkyX4W2tLYWPkncHWSuVVsuMJpLx+HIkUVicbB4
Ga1l8axH98YjR6QAPHdcpcOcyTCXaL1JLxNmgheqCRuasfY8CAxQveiPHx1vwtKn
Z/n7L0cXyOYd6iEvHQPKADOo/KxNtz9aciwBcleDBjWN2sg85885V9YzOF78cCs9
k0kBl4FfNK8Z4tTB9vw2dnQ70kFXzNgo8Xf+pL8yTpk+ffH4LT5wU91Wm8vL1mU8
qcAhLmJfXEk8udU6gXeQQDAUBXkgTON7vyBMpJyZz+YvoXrwpGh2NY0+4fCigE47
Nh1MbpChLfHefXje7tfmfL/wzzcw9sfB++umAPkO2Ql2Opt96ZhUxUO3q/rfoOeo
RPtWda0Le2JOmWkdWSNY6IIteWPuWKJdtG/reinrOef1l6dcRKYC1idYq8jsOzy9
5xAGXruuilnlVZUSnwonvSqoa1HkkTjA4R+kzLJ7vcsNWG0YaMg5yWbaJRNuu1R+
Iq2TGFmChV3baqCXzsbbCw8o/kj+3kq4j190ecqlq8U5f6rBMmj+VuOr4KOCC/eT
IW4B58qd0eirsga+OKxkUXtGjRy3t6T58N3EfzwZsWXSVDD8KXqSb8HnAO024vJk
c3ZZj84alaGLdo6CAjqzUPS4Px24ps6qL0PAIs7KmKolJICwJXemARZ7J+uKSquK
UOEklmLksouz1nHQCF7Q9HH885GgmnwqxQUDG4Rpn8wD8JBoJGI1t2PciLID/NnK
cXhNoyymzBshZzACapgHCCeOuUNm+fe5RRyOSwLIxY5cJITp0ZY071l8Aed6/+kO
Pf/jGfp/Do3LFU116Gs5gsvY+cRjh6EKEzY9fGP1kl5jIeiQfNcK4lJWtC4xiu2Q
969qHk6vUTCjDIn91/nAgO3a9GkBUZLGFfQCd7jAqzHrVnB/v0fn0T4NnVG+A8YV
aUq9Nx0oSQDneYk7CeQy6sULkC3/JqvrqdSamwX5Olfuk72+0M0XpX9qOCYk8n2e
AUQWv8PzSc9A8HJ/NvbVBhDpyW1HZKzeV15xN0Q5qQGuuG6mTYf+gnRMtZ0uX5rR
Xv1ATSQBkKsYOM0X/bjCI+tGGKTreXi2WoiluiZhMenJ893S6PpgSdzTp0EJQOv2
m1f55ImbU332Oj5xDCOICYcczeqPcJMFc/c7kzRRxja/MqZge0zjfrFaOFf31+BC
WnNbHpkkwdm4i20vmXFIU8VyvmrGhYywXV6++734pe3xtNgOC4WAh8+Nuxrr6Jpp
2tuD1tLpIj8wouLjPklJwD7/ltquuzf1Klfz+nH79IVI9MfThU/noKcbfk/VLZW7
X/tu9IR5cxzYHAtpexV/PHxmg8dCk+zRALFxjF2/ZxTZysbnfsiJ6x5hKkbKPsEP
j0ymEM1BXPPJvMLMHEs6ch9Yi69ou4dNT5VWPliZEYoxle8QHsEEK+Mgx4KDwqyf
6n7vadiyHb0vpEEGqob0A1Xp5r/vVUGzg2Rz7SsEBcEgT59VkQcWj9gRJhMLyrqg
b1YqGIxQ/01iINyXph2GFsIjny8V/bsrHlT0nd3kjXxc+YOdxbbqh7cmGl5kQiB0
aj2DY/gOO/OE1rXA6TdT2jMlbvNS5ELaDZv/KqVwUXNm3hUM/YdPHMssIKeGEJNR
WEU1X28vL0BzbpRF4PO4TdcGiKFYUrwJ6Y2KT+NhB0NUXD2BDjYdv88p234yYXUQ
k2OafPB99+88SZ+I9jUSnOLT8qTnNhbkHevbXjZzR3cBkTGw1WfzZknnASqafmkL
49Yg0EvmAFo2PjdP/le2lBXtkhJgiUo3Cv/HE8wzSgM8CpF0JekZJcpOokGkjr6+
HucZDc0Cvab1coadeemwMLFPzeianTL0voY2vHOBOzV/sjQYJNihlMgxWr1mn4Oo
VgRTj3L2FeX6M+1kPVx9hZVi/XcVKHq0amNgKt8Hv895P459AuTYkniEVgZNTnPK
29Gb6p3OJFHi9tph3sNLZY+44OsOWMmXs7IwBgRMKLmv6U9t4CpO3w/RAUvq3lhu
M/mrt/2IHs0B1TWakuGsIkjnQWFkg334o52q6u0RIiMeXKgFajCOcU9cHrYQiT6q
A9z2yY6uOGFQR9vmNZDPTqpI82Ur3chIl/gldWA0OczdIr7A4I53GMSWMwoSIlXV
WAj/BsSoIn0zPA6zpyYUkdXtahOusjY3pb0WvwltrAhyVrQbOJYtZWIXJv2dQdaj
d2xQRsG/oLB/VlljDSTTxtp1a4PJKuP1J5ZTI94oymnVfu6hZ2J8jd0+Sft4Mxrz
lUOBPke2nVIrcSzsIRKIlCiaM6P/JvquF4HbcjGS+1gz0sO5/5tYVi1pPKunGhMI
IJpU/kD3PJMZTyGMy8lydnCsOLTIPfzcmYqo4JuVpjo4bWmfhMkgrcsAhybt3OgP
HA882QgqJHCkv7uBr/Qps7pkZHoDuGZog+QpKjQHomwNXgimlx1jIkzidO58gR35
VkRwZQ7CjY6/Ti/74fgG8aLh+tNeDE8g/3A0WxfDfReYxV33kRsX9UO2/gzVmTVm
fEvLMUEg57kKsmXA+qXyMSmiIyzzxZZF4/9TDfs1UqnuakORmpW8LDpIBXPzP89f
R+aMpd3FlWLHefg7sq9zsFYys02psO2OPhMw/OUiINBAV8QcUPjac2W9fhKMMiMW
HfZwWjjbNJRVQi1jdrogOzS+4VFHo9iJBF7eTwqfVlaLhQ02jBGZ3ZKqVH1sJlkc
UMbNDnGvMThhlFmzPanFQh99p9df1Wc9Bk45Xd/WOd2YKx136F21cpSrCSCv243Y
aAhpODbbnU9i+AImM+ll2pk91K8qEoPqIVGOczshwal7qhfsEBYGw5QUv19TeuGZ
rmRQbipGwqbxZnvDvLIDJtKPuuQYy3bFM/n7MagHhbQFJjoqxRIAEce65Q4UmrwM
JC30pFMWN2k33Iyy7qvZNg6MKTo3R669aULUqBcJRQ8SwPnOjR2AzRif7dMjHqgd
h91NDGulmfwMTh1feEwWwFkO2qwxCkfZJqgqB8OXsBPzbLNZA9nS4NCD5NkokFND
44WsE/mJLYNB0F5XHbAlQEBUaZAuyI8kS79kU3bf15zHE/DVaLDz7XMLYh0LFJVc
zKcjD4CsFNNhm983qy1p+tO/LcKdqEn8Up7dvV0sJlNFXOpZleuN8+2klczoPgcp
LGmzVflB5jPkx2tpKEkM5vrN1z7Rgeq7K5xEvMz7fGdJgSfMYYavSCXipZZ9bVZJ
MJyMcoWdm4Sq8ln8QFf9J968IGbZtAlWTju/Vc/gRl70NhR4iYzGtc8/23rZ3/v/
gHmZ2BtTeXR3+CGUTtm2BA7JIaQCFOVJzGsSpTOL9B3DKaiEeO8MkBZkMFhA/c4/
Hho6QahBp/oEuJKq9j7V2xmf675Lz5OGujOu5r1LXoNvJwHLVZKWErCgmSYI5Fv+
WXAO7bIyuzlAlHCQmvZ4n7Qx+45gncCNkDuVol6xmwiscEpvK6vFvnxAxiuxXE6S
/U3wMoMyKbx8eZ4V6c+mTjM3IFekKBjPSeCQCpYlUqdTvUDGFQ4lLuJ1wEkqxZjK
RC55E73BDQXl+icLIv6DOW+rOCfq7PTDwy65tiwt9ikxENvQlKHGZt/zRTSQHLi2
TIIwnvvzPrcpPVVZAggX8drMphauQ5lTk3V3ZOXjBGIYVwy1DsAEtQ9sjD85XbHi
XEJKN/x70voTGy05cs5kzKigVEkewSbCTYSVMbpOhYU4Ccw+WN5YxVzRaicYbzQo
ioy7q1CtnkcX1mggAXI5AxwaKzczw0vGHSOADdUu97RUFZpGOe01UuUgJwr+BSio
TEGAYY3QX25361n6c6Wx/xT7aCu6uxqg6qsXDciwFEpUkaQnonQXOVnvN4bJJi+b
DzNY6MrY35GbR1sa/UkHma75myuRt9Om2Gfxw0ZLwFkoddAVUCkSLMzjnIRkzdHz
KLZMIbXlF7L2Yos2HKviDX7NrDhVMCS+jG/hSEyiRKbcyjyEEVRj+btExpe/RdBj
O62SzD5VJHEciY7iGQXRLo8JIerB4VcetzkZmiUs74lPQotb6UDWfS6AFH2n18Si
VpyebOdabHxI75CSv9zBl/FZgYUKleP5q1fFjNvXgfPO0/nB6k3b/ENL9PMKz9g+
YOb87Ezy4fAKFbN4V17CIsDTXhXe4i7t3VEJJGy5Fe1WodUqEUPe3lf4+/HrO5xO
1upgliCquM9EUmgduPh89hfos1k7DiCVUx0udBookXRi2XtbHZv/ogTnhEPXzLiu
bzSWj3lWcoMMIAUPcZhtEheZtAu6yvNosyWJM0lQGDN9jWeIokXmNzSBZllx7L2t
r7yv7YFvK4cLOPaCUnsQbvvsO0FA0ieQBvsADECG1WpGO/Z8NlYM/RuyZzBPfqBR
hlTzFE0kyjeWjpI5OsjraRuJoPo1h5/I2mcnZps7zzFAo3dgLYIqlfTinDa5StzS
9cxLiPN29EvWVBNrAy4E4zx+u3NaETj0uBbU+Cx6RfaLsZYZtY3N4hhdndkRPGA6
ODVCngQZETk2PmjMjvuqG9QU0pNvYhfur1WXmB14ieMfkIssMXJnSawP7RCMCygy
m8o89n/nJtvKmHnFr5x4THX57VWQai+A9PYbRUJpYEew1wx168OjDluFMb0aDMdw
CzR7AvR3P6EOvESccxuoQQGvbpC62lB+UN6gbxSU5MrkzWF+YXxGlFyJ7z9TD83p
IR1l2i3p+3Ygrp/Mta5pojilAVFAK1JpYrctfW8kqStyji0dwAyZLffZtXhKJC9L
kEWaoNMdq9y1QcLTgZZlO7U7ATJltiyyJ35dyHQN+ZDS4+cvr6k6k2BuAkfTL1jM
DVWKYp7i53ywvG741ohXQ22HaiQAaqeTDM+GJHTV1Oaz1hUUq8v9rZSM35nWxB9s
O0kNoZ5pk9ARhvdnldLKG0JMRTv+EaENlvdzo4b09uHSs7pUe+Mj7AEdk7/Lk7ZH
F/He6rW8K3qwzEjdZOw4QlPQKI7fmFUrOgWdIik+k7LFVuugFjqIkn6Cp7tm4Nmu
0Vk7GqW0G6voJhbALs5iWMlnwBFhXkPtOucHhPp5lhGzPQZ0G8uvLqlA2W3avw2m
w3rU0QSEu26gcxborwTikJm6Y5KMdtnN54hhE2I1lmWWTpc/3VZ/EyhYcLjrn43E
7BqQRcJ71hdoJ98TFF4SQ7A7XKbBKkx9M40Zh3ouNsGN88DiMxS6jxlTFPa0vIaZ
ASO7eTIWJ/kVn96B3XAMZgGTRLu4jvueift/JVCESryJJYvuVjJYyQKPcu8dvPdb
gEFkpIAwa1ejqtGOAKy0HSghGxPxqJLBDYXyRzOqcdCum1ZmnBYH9o+FX30hQpM5
lqJLDDn4g5qy8TQMWOd1Pw8rAajlHPlIX0LlSlPghDZeey1A1KuwBmZefAmcGtqb
KLr/5XyHTsQBU3EWyvEUGqjmmWOOdswl14LsOevIvwNimjdGtDGuS2wfd1+CROnb
ene6PqYGgPRsRnxHj/aIz2YgA37yl/tR6KOo7hMTCDy0dd3CU9q4h2Qa8LXhVqWd
S1CcVX8vpTdPzO2PN1rT5IbxRRHRTS00iT+l3QJUWWLnYcgrw9ds/zF0rBp/L1j7
4Pg4ISquvi3wUqQzwunPsf8F9mdwSPjnqFwoAjKcq7KghPdhr+qj4gqIVKdH0IGh
tO+meWr8QNNxTNEADHayC5NJo9ecgLrHZjlpHWlogUmuqz3DMpw2GjJZXsOwCyfx
2zehbp2xxNUbrShZ2cWf/T0M30lQEnv1cUfZtFREK7gvxkKM6IUiHz6ya6fouw/k
77gCQKbT5HELyxjBGj0UBmRGKLPXx3MQzvkxKFz5a+Up3vEWCnahg1izIYthmSEi
n9M12Jjjrq0sW+VXx3FxhP4yVA2HwwRy/OeQHk2gaIlGv2sfIXO3WfepuoYQtrnv
bfrWb173no+RiPbD8okiP0+zX7sRQVI0eaNlDIyoGW4agyTiBVqyaRL/qiyKO5cO
awWs1CIYWMwykJVikAbqkzRZNmnKeCgqQwsbMd92Bb+XtT26kCelmng9BrgS5vBK
pPW9EOcIgZ65EtO7mXXq63ykulVnhVIuEWBtcYfXZExXYVehB/8rSkZSkuyp6FoP
EDKJdwfVsXO5TTP6mExUaPhj2vks/+C7i6vXWZL8votp8sJZR9js00MzBT9UEFpx
HJiAaOlBdklRsCbvvX9EAo5Lc4/iJoXRbCmCOJudDW7GGDEsPs1lnDMBFlTe+Kx2
whcxZQFfP4/LK8cEQco7i6x4NDIadg2nBfiW3f4LgMBKPnRDVd3LdD1rge5W999I
NDkIlNWCigLkJp54g6qtJC91zRhkCtKeM4wv/3HJW9d5n97wV7I07qPekIk0I/FJ
IBV/7m572aDXBC74UDQpVTrHOHJbDzY5OuYhDcDHrxe+x7hDcNEIqea/R07HMn5u
5VyuG1e4UoAsd2Kxzj+QPVsa+jIRC1tw62PFvgg1PuBjB2oaxkBz46SLk4ReMXdi
4zqW9g2w99DSy10FmLtQJbVhDU/gQbeBtx2a1xkF0ZA4d7cGMzw3m0Vs2ucvJ4SM
IyCjxGwaam51MDwxEMY6kj64GwvHnOyHddRhcqT3vtLV+ahrlum9TAexPAlLQNz6
Dcb1OFOnL7RYPJ4AKFj5cubk0g/QUDy0hRkwF4i8zegHQ7ItEWVJ79JekxjtQnRE
Hfty9e1t7cjbzKtbv5dR/ElmqPF6IEchfTC2ru68SYDpYo3Tf0gec7pVB+U1js55
sBihFF7YegR6eS83sqmt19Z1SO/do5J893XA1AP7nlN3u36Ca8FvyCU32Ggn5TBD
EsfJiz1vdgKP9MtL9epXadXlpvKpLLqVGoY1k+SMfjifHfcx9g4XpfXkN5ieVRhZ
QqkeqbdFf5Ibl/DQgwYcDqe1auKhrAfTXuabGOXDd/1XbvlRDcb0ZihMQxV/BAMf
ucWvLpegqqSchG4kyZdDzpFNCcqw2tTmFjthBcGwUo/M8cB5SW5ulDQtPnxf6qbE
OHc5hreJdpQ356igq/yhCLJFUgs0SsKMA0CetgMkoQgXMsb88DhRduXS5quKTJg8
PuTB1bHKscZ5Y4/71895pEoj26Hp7b5Zim/qG+3/yduaGyJVqoFajMryAoRNACUu
8uTL3nxbxVxu3+yUSxO457U9LJ/hyTa8BSFVXT1FvXWBpHyHkk5ZeYRSZlPHsMQj
wYgIDdWy9YudGMInJiCRMv8vEF0i+IzHB5894RUi4jUjvbBLxR+ECDOEpe3oH8N5
wKLVy2upcRTyhKGfN09ZzBP6rqE8WhC/Kb5XCnfRUk8u2tP/7MFvquMFe6mIYeeN
35qQAUVr0J+i8X2i3lIPEjQsKnuaC6dJqGTWdse5+6fP4hmpWKZ7GvgpBV/1hL4c
35kgK+/FeXcMBrTx6hCF6yyBjDewFPsl0+0MAjnx9+33NHQDB3yp129J6NqTF/Su
4OLRma59Zw8cTwt65/vXXP7mQOe9rsejJunI2ebC31L7jdd3GPpA1qN2y124HL16
lgOaUg5JEKHIk8e7gjmgiY2DvxVHW45obGL02jTlm3u7SNNSKW7MPyn/t0H0GWM8
g9aUchjst4B4t6J5e9Y67kTEBqX95i9OUD/FTzg8J3tILJx64eNjHocjGulgLlsM
7ou72ZHfyiH3zYxCLInRlLHYJigXQ2puC5unN+/Djml/nDADagCwOeIEZZ0ikkXa
mX5QEr+4lfdJehqQN6r4Hk3ExwONyTtMyCYyNsNFuN68ThdrfrRvKsbwT9BtBrgy
Dg47x7RbzMxnmlH6f7QqiRlSr5ctPqiIrHxKa37Y5KQMDHiy3QdYc9ywjMuCUXjR
hmqGG/OmCk7UgSKCDCzRZvuI6KFZZ1gZF4/XyWQVk7kCuy1eTJcONiXzWg/5xpsP
GJdeFU3T/n/dotih/AQAnUDf7D86RMOVhQ4Cp+9ZKt77Zia5qS+XFSPEMjzdbLLM
QCUYta6IqeNnhNLEdCIayrhQzNgTURyAj51+k7M9wW0+57c6ZWSVV+xe//AV13I2
1cDk88tJyupFbJbBrRJO06Ns2lvBnZE1D8H8l444uvjAIEGOasxBq8p4NkVMOe88
qjO1KXhAdZ3btUYaMnEcEl1lcx4jTwdeFAzT/kltFpAc9qo52ZRvLg1vQnVPk7ff
oh2X1j5UdhHe2g4+75optYXaMdJzDHeQCt5LhOpyvHqyC+cTiXoYU4Ls7iLg+rXC
+fToiV+oLzd0TTMl5FRSnL62Z6LyASkr+FbBsmixyMg7+Y5ORuCUfdUo4XyOImxV
yPpv6w6Gus22BMkXS4EBT6OJgV794XRquhA8hTdl5XtGrQGSz+JdBDa+gGKhX7R7
x6nHPSZW+ybbeKKbZe+2kmq9cH3yM2BG9lkeqbAxJuEGc33KJm4WPTshDPUUmS0u
B1hqXzzYOHb2VhCvCVvkxVqNMmw9vXR0LEDY7PYzt4jgFJHi7SYSLBUUXUySN9mB
arFq5vPwNjJEb55Juu8IewYJakPGbD5HsnzHjGMmWTuA0Dw17PcZUIirCjzx7mDw
94E+bxGlU4mu3wP0ypcxvhFLVKcHZU5pljOImBM+fdm6j+4v6LEt22RCaY1Z01XQ
JuI5qGkGo+ck+dpkpDjXdtSYy5ADFyrgGN/eszc/60X2J3bVqrEvPcJS50vwXwMN
JM2io7XNWhidhZwf0YdBA2qjWXJ8V0Ixfo7wQ9adNYqK+shQxpb+Zv46X4N5n0bL
IqyWSOPpjUtJi2SDS2xLEcLsmflDorK+UEx7yunMl4lsMD56K9VupCwqtT2J4G/M
FQz751W1uoU/iNk3SoDHCHhi7VwPwXt+//yTPnlnxMeoGm+GCRuBt6xXy6nLawRI
gcevN0YDk9zbgVq/zCQPq62NCtMWB5M7q8lKYlSCBgF8U7YSqssU0fI43yyoPCmJ
X4TWKBUGjR9gE7V44hVT8prXBIFWYc28jQGxen+aoudtycUl2GgqXXv2/1jrw4Bg
ikSLPeCkHNbKXytU9hdGeCObEJ04qR2nYhKz9TXgLQgKAFVtepJC8w6DGjmZTx2A
YYs2fD4KFoqoUBtgy11HZSkgseU/q+GZAQ7F6cDBNZjD+/hIn+JZvKQRthwR7Tcd
POVES4pAkADFMCHY58MLgTSDrTluIdhYJSi7mWKP8gwa39cGIi4uGYIe46O8Lsz6
goBDN/dSaWMoCYh8zag6AyDBciKcW5oGjwcSELQBnBaGT2wYUjIGoxRwlYFlecXQ
O+ZLSM0SLu3bzloJ8kNysf0M9qvOo5I4N7fMFER6bn4heBwLUoNdvNPHjVieRnWl
QEAoPW0rhLENLhSLEO5lbOYtKrCIMcDeNQAE6u3JQyB+O5aML9vtVoA/UcHYt1eL
w/f7lU9G3xNqIzNiORaESvg8fpgAw2SmyjNFQv52hSwIYTx4sGCx7ZUTMZok6+Ph
r36ycH/+A7Q5ezjHFJ4u5b+e6ky7gbR7zVh3CRN4Wic2dGrcl+ILgPqCLoUIJEE2
mdoRWjGHLoOy93vgh3xhH6sFDJaqvel0UeQXyZnXfbqHsz+nau2TD0NeyObUF4wF
Hf9dzGll55LnQQ0Ye2xhnaAkWs2i7Qzg+3WYTI5ZJdZdgDD+D+5NxA5f+H3IdumB
523TYR3HnqnjBzzY+Wt8/qykn4AgIGraIZRarxAWbeNSZnq2JjV/ssr9qZ3CeBj5
zYpsYZKN4U9GdYOrl25AitR6GGfKVYktYUf1gEARzbQ8tfJKsHDH2NcLN+mez/I+
oUhhP1++xXViPsVoXdeSn4jTPt4ArWrPGN1VCrigmN8L31td5O5nBpam5VUPCVFT
3f8ru6DAZy4WcD0gj0qy/BBCBqBhjg5DZtUj6PVxVz2NLAWpMTMW0xX9QFx2SpoJ
zqWdwu8NQFTjb3hp5hEnGEh45lyrDm8BgUrUfWgiJCGgsAQtAol2VxNdI9Xwt1AV
UWgaaN78vFF14daGlcUIgqyj36l4RhXVnBMdlK5wfEG5gXLbYAkAXrv5ICN18axI
06au4P77Bj7WprI+7va61k5pm7ycBPcPS+7Kiwynr8fQtyakqfzyqBsT9/U/eSms
pK4+IYjvW4RoPR/dS938670wk8winuy4LUZY6TZxVO0Zyrgx0FJznW0NSVXkdU6r
lvoPqVWpaKgEsf1hoC4r8LeZXpU4iXGSzTBSlI9OrmuPzGUnMv1q54z+TNS4yM5L
4lVStEZc3K+vN3qYmbIXjiMGlVtryBV9vWetQ5PLqphgV0tChaQEayNKGWXJuMqa
HAfcRHaNp/4MEZR7f364/QqNNB66auJ1qMy+WZhVsTGE+RfL21M1FF4I9UvZwXW1
S+SA45zumUugLthp6c3TQ1BEboQ4B+xfzDOsr7AMC/xn7qyMEbb8G1jsviO72ZIw
U6xXzDC8h3U0rQ748/D5uUTVmQF393JJq0SoRqgjYzoeyoEiMh0R7MD+peLRNcoG
mO0I2fbimp8EdaJrwvvnnRi5Xb9R/b6pV94Z6vsmzdq696A+p4sCtffY0/f71Q1l
Tx5iyHOkskMd7eA2h2PbnruQZ7h8/7T+Ui3x/c1l8MUN3+kDj5dWqLcQlpImdY8y
uqLWvZtPvabBUSd0BOOQytdOmqciymKkkalkXrSJBR5LsiLQmpJ4mlneWDqo3XeU
dI/jj1q1V/Jc+vai+vnXmhMl2GU4fz5quriwTTJbE3DpnQXhXHhDhIitP6EtrXux
mS/CUR0VKpBWWvEG0/5FpyLdClXuI8Ydoy9PDLKf0SkQoYKyLNWbIDjEUY2+ZgYb
LjiuC4dMrJXkumhpGoKbSWnsPEiW6T5UrAI7bPTna82vb3/ip7OVvaLv/qDtHNGd
5PYCr3XLGbCBrBFJuQQIwcQGF8whchtFCJovZ28I8/gb92mDJLJfM3xGU25vStYg
tcC2m4WRTP2ftS0mAAaTUEAS0/A+eKnc2PHcW2Ugrw6hMVB7uGmnfjqz4sX6ei/p
iYx/ajUptKl+TuEMuNTPQchGpKu0F2MwYxbsoGrOFOdf5odB7WEisWJU3f8/xU71
Esu8O3kPIt/DiRzv78V/8F6dsZBE0Lm/H7izydauOvxxHyZpE/o2rTKG4y/FKfSW
KsX4p41jMvlUqPLCXcXCc5vvckBfObnZKGAYWhphF55Hq/4faczX8i5uDSl1XLJn
tLz/8O/y8qke/tlIIXCSrpOAPBYsGpSfZ/Gxl2TOuRh2+oJS46SrBuQDhzX4PqP9
eBin4kKcllTsYw0mqe7UH2WHovYAfSaaLwAIDeqjVCLmDFKYUoptTEgU/HU5OzxV
wSseYIcsUal2wv8H9s4uiH+QDGqSaE6NNU+CCKMZE9t7jL1K2xWbHLdWhslzTQuL
Gqa9/2XPYRyWtfsRQpHIoMOCwIDTbYqHDwROpNzWuHnPoj6tqjJk/D3iwpA95cvW
J3/C6hZPl2RgxMCqPwaHFPryslq+9GdKsN6kzcrsfjNOEMDWerJIrOK2GNvP5K4e
z05WzyUSW+AQhzidSoEpBKa0GaJ3rScmzcs8EoZZNxH/6zuFd9MLDfpxUndyFY66
/vfrSXSoTuuJfW+gq0YgQ9m8fMiXtrhxbL+/zDvwK9fGk08V3r/FKp9j7MRXBFji
DunzAz4E9KvFCrApOWQKPCdCkn45meAeWb9dGM7tgI9IXo/iNDwy1pvodxt77wqU
O1vyd1omUu/XjwZEY1kyUXNgn3FCVRNXK1IeJ96wGR7TcNlo83k7ACEVGgDgwUVA
BSmJE2UkktbzJ8cGNLnAs5kWUBVzCn5JQN+eFlZee1P+5O+Q4inpiBUD+sD1fsHw
ycvXNWQU4AeG9pBssrJTGpZGvhDQ1z65ayd7YAgH3FzTsraE7wM4Ip0jtDfT979+
WXDFR5ttRvcwnGvNiDBRU3Hr+VSUrd7hPgCzY2PR/Cn0StEP/hoJdFznYDl2JHuI
sCa0WjqWa3D62ZMHSHvM/gB/5zZqwM2a6UbTt7wKUtZgjunv2TZDPkznZXddykfx
jqIdKXiuCj0MmdmJapC39mRFJBMJtNfvDxMWejGvodEOqH/3HU+zf9j7H33LIGir
oBe+2ZmVEm/89JfsjzSs4qgsbd0ddvQw6x8+nX+IqepDEw1s7Vd8RrpoUsbcuKuF
zlc6skpR7kNdcmB3cCLsLEzgY/uDchGhHjXfvblIdieKRlT8TuEUXNpuVUA5V5gp
QnfLiVaApKTDsbcPRwLdtRS8sBedcaAjgAAju2IzKt0Tuk9pvOW77oi+u53gLIoZ
LsrppKpT2cbxlL6LenXroK1Gg4reH9BCv4hkg2WdhpM+yE8rFM74lT4yHTsEAscx
nIWRZtR2VzMEvMXm+R2ultbe1MHY/Rs1hsrB8rrhx3zzKpnDnHzjXuLMSK6QkwBf
fZ8LoP4eGzgyi0n7n0zPZBPVI5AaZNKN31cTV7JYji3I3wsR4Ak09JxlEMbZChOL
CGhE78iwvoRkHWg5DbG9WdHXxgEhfm06lughQ562HnAhx8BQp2a9cYZ0j0nmEigK
Rku/n97+D08RV42iLC/wI5WHw499lhZZBx0MWTXSwoZvhOx3qfKepJWTYjLR7Bmd
jM9j/TgsF3JdOAlrxMyjsBZAMOA8Lqt9ZCOd8+4XXYI41jC2WR7WOp1D0pa7fVku
xmZf1y9PLJvM0jWRLpYFOdNqEdbnD3gUf5j5R8KQDVn+cEQ27jxMXbf2mdR93+jW
2/63JD3dXsQZ057ATHpXRaHNMvP6mUgvr8bSPlBzKAlA8PyUWQHxtv1t9l8VdW0J
wmR+wmL1xBSp3tCDFbRg94pN209f/CmzBQ3+lsLrBnXqJh33ph7t4OTWMwzmPPyn
XgtxjDnjqWZgg+y2V4B3Sxsa9aOzwkd0t8Wm6nrMLxaX2bcj+8kIAUZ+y0tno9bM
V+SU9ai8j6VP5xc6ywTOCHqYOzd4pynQzZWba5E97+2guQ0ZRMErLsrDZeY9GR44
IzvSS2VdpYl3I9mPapj0ZJCtQkVo8rnxVPpAx2epYEkLxZs5ietCCYT1EEf/BSaI
ZN2HCg0VumI2aZoe54sP5udhwVQhC8R3cIUTXjW2wr1ALfN3uxS5DPqHqbEGUwb+
VLS29PBfh00tlUEARNhsxpjRLiAoNY0SBgFGdZ6Xc+aRdP8GBZiyfCakQ8D8WuO+
UoEuLOBm8afG3IU3VV1l8CSwMt7TrpRmo51Qx+NGyH8WmVNHwulsP5fThqq7pjRs
qk+1z4ND1C0IsxpQZ0VSobJTbwKTb+76+kM9qXZ6cmH4hvQUszHi6QUflfHsuouj
re8Vb/6RlyySEF3Ksf7DpLSBCt68I02Dp5CbDV3C6bXPo/uWU/GWmtcbDzTY0lP7
HzzvWbEUsW6qmXu7sJ9V3EWkhBoBgMiyFk98FRWWekf9bOsFxHJQXAgk1GbMdVro
/v7kKvkOpzPhOVCx6tJHu79UJOg6MRwQIeXtlWrXxTNRvoGLvwTxXgYnQWBrUWMf
NyMDDBjJjbuveygXjI8esdRuHB4DyzZyqA0YEGUhL7FWwcIfh2m8xixWVwLG4XpY
aLWZX+xD8b6M7a1Z4T/dv6ZCTt/ths/mo8VgLoIX/Jnr4P9LNMESc/hD/WQVPkoN
8ez2zGsxn/CP1RV2uaX4/b4Zq/H8rXHNheDIr2OOYVw0/pNoNit7d2So4LD1K0mE
U9zxLnV3GlJUiBkCaIdyzamHZeMpTFTPSU2gMrUeJNOx4424+NMpGRvzW6MtjcbV
QO7nhdC+/r588ZgcadUwRy45NHGZb9Uskiu9nwQFS9Q9KlaZmaI3gmI0P+jkAmM4
+QYFoO6vGRDQv4bXziJK5sY7j3vQqZqmMJHRZJW8vhEw68Kyta5h3lj6t7jtdlKG
Y4whOAo0tnSXaiYk8u/waGkgOF/u/hoA3Hb9U8xM65kCGNEWTSSzplfSk28QnzdM
2YLr7EGt9KBp7mzHan2ikPpy1LyZMgyL/WT2FXHvfb3Ku2qrK4YtGnx5QRDY214y
qBjlzRDizU+jj47617Iqj8KBsFayAOe3wvYOpHckURLi6NdRLSoFAgjn4X0KABBA
4TYkql4tNqQ35eoVXIoHM19hNxIZb+m6D3tSFFHdEUb2o3fd+yPoSvmWhR/14BS3
e/Y+Xyg+d/8c3DM/QuO9vidoVG9CvUVuL93buoRL18B58xkBQYRxPFNA8xdWGduH
b/8BIIEGMBt0GzsEAET7/BnvWYVYBPK52aQnKc7g8frhEtcDWLNvkJ+Rj0W7Yo5K
sl1MizAquxwdDq0Q8NGDLHADbXVMw0XmlsKgV1JTtPidDVyJYw0tCVTPJ82i2em+
DrPyfm8dxw0qwX2knenfhogEMgv5Zyb7bQaC9NzArmpsZc5RU0sZrBlGJbliEihe
Bb3P3ItnJuAfXLQCDyGLGkLiKOrpbqL3kqLvlHrvFf7muVr/d7dFJH3Rzyl67aGy
y394YkWiEgZapOmIZh85B2V96/YWHEotc0trDfWr+KhRo8GTkgFUwzpLm7PB5kG7
sObX275xxVCR8A0xmy0HG1+dFNUUrX/24NDuxEIs3Ly5oybk2r0m/VnkcjtmfhGK
CiFplfJ4SvMFjlx7nZ+QVX3yDQFr4akM+YEuD+Tnefyj2RuPNdWBrOWz7euWCjsm
cZRyxSxJMJ4lRFTpvkS50zgOlvPsWSdsd8izTG4e7dcbgpSCiKzAiF23AHEFAOg5
08j1tvtijWLjeqcM0AaAM76Vd4Mh3TSGoUKTH923lPqun+yCw/jeZ9hSxq+FmiB1
+/MV51fTqw9xTeLB5WHb357gOuxUDzywbQn8uKWw2UkbwWknIldFAqjLra6eeAWK
bvcPP50FjkfQg+YH8BTgaQms1jK7nEXKCJG6UN/6X5n3zNgVZN9cYD7gpaqbs+kx
7t3ovQq5K+Nmg4XHDe1DlYPWDu4GNTd+X5pULy59mnUnkIpJITGkh3OfuOsFe5AX
8x5FdYBUMNjDUktPLDzfudTxcxL+iDjSLwOrZjqXb6cQTDaQkP8C0NtGE1C2rvsy
IIF4Sb444dJlNzc1jYSM4ocxsoh0LgKjFyUg/k3ieLohFlUlG9FRTJItTnhOP10y
HM5M0fnkR64FW5wPVq5O0BhWYDB8av4OXVNW6CEVY+WDnA1bDwJhY1+DAKn1IODT
G3Ku3j09i5Of76DQ0eyCoa4tz0Cl1vpR3f+3/xtdVaHMv0qVaGeaOEc7xFJpTlS7
L8DfiB4Fn7UdQQwXAptMKDhW/USr+O9a2vlNGCM99NwRvTpnoN5nNTQ/4wm1VOGd
rMVbywGBYMVMys87i7vBTI2ifW48Ff0lO6SVtgrVVAGmIP064Kmg76/keUOoj/f0
En3blSZ7hoUhIB0ckjBytmHhEJeuKUiClSHs32m+E1cCAAqJkm/fkCCkBQ38IQq7
svlkVzxUnV/4eYw7psC64kTiBu9eVUdsjukKiImLEvL3WEuAIiG6UA0ERSoL+59O
G+uizDdLHYgqk0QmGfzpgxra5icZobicrQnrzX0D8STyqY9JYOtVRhL3piwCZIA2
1KTYEXO+T68/eV+uKnSVKQQzg2LHkf/omxwywSB+h75U0KmOwVN7uL/w9a0UVdlJ
EN1dzS0Ijbpw/ZUMCliMxD35r7kMk42wQV9vKYmWMsIKd80K6z0RWYcJYsM3BSqn
8NcqsbeCni6YInkFdKxhlx3EietBuDQziR9pySCl2ky1/5IYsZOALhQ0x7VDkw1N
csT3aOQ4VktDnQLx2kr7waqMAUzNHxjRYWd81Fj4Xtuhu/c5F9+ZnVgUVZEgq7Vh
O12ssRkrSZAppNarunroE0w7yPPrFH4RgMTFbywGKQeVu1PX6vfTluS7pNWgaD1w
rYHrLi77TC3zQUO0uU/D7frQN1YcK4COr4awNlnaUDs9K2lpDuMago8GpwpZlVTx
FMR7M/tTf5nJJec+JScgRBhgRBhI2z4kAFY286rokxJSmtabhEMbxgBfjG/nX6j9
/sXeVYWBnGFPQoqRROrn4940QUm23UX9QTUBp2ASWD/1GajbvvqGgY0mW4rJzIKj
XojgUmZ0ZJ64xUfrxbgdiY5B3mo/aZzGkFjIXiSQ5sMhg0KMbgWWgU6XlYy84Obz
I2wP6JYEyZNeS6pCqJbspNAC7Y/8KNaS8DvYTvJ0JqVyUXKZbXCKFAG4QSSKUvPQ
cYbu2CA1Mxw+oaAclURPDJ0uRTRSQ1nhS+kdfLeeluvGv6h1G5o0p+8r2Lo1Sq2u
Z2rIW3Y94K0kC15cvHGy0qKsQ0a8laCU0l+8B0o1Wuwkw/MFKUN3vFvRWVSXphs/
lHpHvyFeUPXzJrQOauNDIkyTUZpCwjUPqU6TQRzu8r0HuHyZvyqzGTxIDHXs3RE5
IcLvBYX/8hP3oYeEoqPGoUhwGefWN6B6TX3jh5a4rNoXMX0Eoo5gnMehxFYjlXhw
W4rmsVAPoyB/IpbDKnRyI6PgLXVURsmJ5Xu18NFJLdRSGkNZ16ZlqhnwWN0EnM6A
6kBr0A+XBvk0bhuz5NJUAgjelfzfwAU2mgwd2K9AsB1UFS8/7YJBQMEi08JX8Eue
8BhOLWyHcpcDyJeBA79W7q7Grr98+P1793u7cR7ifz9cBhb5DgK4idKgnOQug315
/zQSptkVyr0ZLXMCxl/mH9MLaMHhbaEj9JjL7ieCNKYyr2FOoxTnfdSwMVVklo4C
3x1MQjySfsUCQs4gwFto02juZFvfCbQyJr2zYUx+vWGy5UPCQM+rWUJBJ9nzunHl
1VMBuoE5aOWnzRs6ls3XDxzWslHxBcrWNUWgmzv+FSSSjNIer+5yODCENGQlnlK7
pKHcpDB4q39EoQNMAjD9Iuf0n49grpFQh8JQHCzkOfsdHJPc5dpZrZmeBAhEBpSc
s0aw0G4RpjurNO7P5ot+fATuTM+AC6kjUEHPa2XiYi94sWAePG9sI9SkQnxjXKeo
3XMZBVBQXCV2n/6BKLeKQpGd4d9CG5euyYoU69WYc+LaTmp5bLugVsNViNWbBklx
bAA5eJq6j2viqKqLuihFTI+dtS6BScVnFOgR0En4RUe48sbnDgtYHWLn50mt53t9
oNNsvt4usJwM+WnWiFfAfUDkcRWvxM0Dspfn2eGstYgrk/4AeDUHMLr+wzHIko/k
LSrv58HqGTfLgCWZ/FeWfZ0SkDGQKrQ6/gCgi8ZxUX6BSCSmZbRRIelXIzC+9DLv
ka8YzOuMbMDf+xF8hB4Ri7zGKhoUmdA+XQ/eumxO5KfM+kB74Zt4uc1baTE1/Q5C
BE12eT0GK63TcOyu0Z7NSWZbkDhx59bdtRutNPkOJmfit6V7UxSZLrCxneEuYx3+
cLHJ3+DhsEjPpZRzbMRpog2GIoxTf1Wfow6F0KZsNbo06Wpaz7aVygIEi8f090wx
Ti5ZWkQA2rODz4r6mRh1ZO2TuOsYShJCZtVOfVLA7Dx/+R3swGr13LeBAqj83nK4
amDwj3VUsnvkhFUr2aDO9PmCsldWncSDIPpCCrYr8da+/yy0ErRgWGteUFePE64P
H6VrC1dDe9TCw20UpkHGK2tpHV1zsJ66ovEGIYzrYGI6hfLRh0kTJwvXGINo3dTn
8GXTti06Qnf4StxwXiF3piPtpOwkHaiaeLt60Fk1MocJjbkMvYRlCRohZZGx892j
NKfLWAyihMSSYDrU8sSzC0NPhvKVJWyyXtPmreNWlyGiuMHvs3il5B/rfIZ9DMjI
wALxRjK7ZpwrRPEJZuAUGhWDb2/PD3m+b8HpnYsY3pOR0LF60O7sMYk+mKbLZt1O
TSsfm5PDZBRvkBhB+GYTcyRxSSKsNN+fsVmD5YtJskqfPJ9ZMLwh81Iirm1+amim
/rSGfh5YLh7nVx7F/mo+uV7mNyq17m3RqLJDtwDpfR3+yv6wCedqGrEhE3/A2J29
Qw9qtpOztZP6qSF/tdlpfuwmDACZ1Y5Z/6hxXpdnsU+sq8+HvsoGpzmzxZaDlDhj
BJ0IF3ELA/Iy/IK1bL4a8QwQDEabzNM9FuW7T/impV2VNxQiMj43I33yQSWAe7Cv
fYI3JwL/ZASndXlap2z2X2DFV7vlDlja543CdxP1ndA4BzCfrQ4+VGWJIpVsQg32
24Rgga6obUkSGhV6hMntuft4oRFfT+klyb5s0PXw8nQckEhhGpdMr3y1djXUgkcJ
lc4ox6vxDYNAUSaArUtYv2zEJLNj92qnLomRp4+rVg3vz/u1AKQvdVwQBn5ihb6r
nF5xdSO6LNEc+884NyOnPnxGXYHJjB41FcC8PCStabE9V1Ss2X/Si13xAqTndGJu
ZVzqEq8u2ajMV5+jx/6v+Defy3Xeym5bN5OUiRZHiKzvPjDb+/WHymJZMP46bKIi
PEezK3eR1NSjyB+BZwRr7Cx5isr7eLNdesy7ISNiD6Lzc201vz7S72fgrxwFvg1y
5EIY6fnrQjRsNbmadsh7WlG4q/X1PukL2K3J/I6AhvDkHzw+BgRiCsrfTp+3XHl5
icmA/2LjF0qdtUeG46Vu+bR4M40+bcp8ZgyJMGEfQiotNuW5usnJveoFKpu/4s00
1Yxq/jlO3Kw/9SVhs0qSwLdKL6pz7WktYBtnYmIXKMkgDa44TCC6ZRHJqRbvZrxS
hBKgAmIaBrrvjxLduFILVVI25GlnT6UYrJ3BkryhtoU92f6Aye5k06q0n7zT9H2j
KuPuBy0xZ4gZZ5G/rdQIRvFZ+PJ3/F5RhKA/Z5dRXHZo548HApa/zRavzHAsvYuU
v1U8oME5UwSbXi+73D3P9/XPjlbayn1oqjV7Ex1pvrlQ017MA78/rPS9918sd5vG
9p4QqL1MgSd090O+njdnY8wFDal9h2oafKT2djAFig0cESpmrY9OuLFw89MoWlpE
8kHObKJjjXxDif4cKW3NDpQQrA9gHdrKmJYBjEr8N2JLCAEN+Y8BRhor4XcMBbsu
lQDE1YEzFv4nPbfireCf/PYTmcR1qCoVCK/qYFgSe5v91zNPne6cq2gVTVqHZUN5
a3ONLNIUD7xsf0iryLuK6czs+kBS7qrZLrUJ7Fz9XTPC47AYtKSGsyTZMnC4VoH5
fitRw5bM4fZWQwQFuH8jYNL7RwUJwpDVuq/6MXSuO2Xf6xVR8795PJQcIDxCkIj5
QjFidxwOW8QALIxa9QYR0TqXNkE+0LDHwmlScIrH6f96jXkwndghu4eHmMsBPp3K
2735PtNOgdjAOn4KRreKhekJMY0lt3togS0cBR7oq1ACFs0CWDTkzI/24Teq1eUl
h2y9QKWp+XV1CpcTRO3bn985ZUoQuuny5+bO20HIJrB18NuDWIpUM894FM9D9anZ
2qfvaXP6mNeF1tmt/ABsdnF3KBAIxh4bKKYDWWmoBvhsd2Gj+c+mC0/GRN/zjhzd
S9Jy8uRNjo3K7Y0IfvFvQ45tRfT+IY5FXhRFLYMaLn+Bq7d2sPp6xv1klXTK21vP
wdzO2VO8YgjEyf9Bes0z0VeRFbKZFrbeMMMbsLEuTjUvtr0b8X8ZTA1IOA8x0gMi
uwrCQ+2GiF3esOGxv7gRyIOCo/9rkXTlh37o0KZCzgdt4WCWvzTm26ng16D8AOm4
HgCzfXh9P+1w7XszrnFiRS5+fkLCG7/945PGzBpNOPowi+QNZj32nEXFm6oueU7d
ylLj4ikLX9wNC+OdwKrbb1LvfD2aIIxW6jwD0LogOWZhYseMFAOS4jNXFSBKab7r
zkBb9haGArm0IHF8UJB186CAHESICh/AK4YEYWDTEvfDmkNrkMdmXR4UQ1SHU2Q3
H4yC16VOEXJKzEikjTX3EtgwbpK+SlUMEDsu1NLudidWOP042ApoP+BeXu6YR1nu
5C7HDTJ5BZfVTbcAkA8wwgZD2rxE7+a13eCYwg6Ht4PCUzayZwveTG+kDBRm8Q0/
0/NkPOWuAabfKMKPp6MqAnY1JiSjFI5+UhSJu1Urn007/wgJSRQQfAuPHDrHLbSL
35HDB2wAybytS5QnI7TrPv5wcf4QMBrZ6f0RgemO48Qj3eGE84rgwwg2ke7h1zfw
DBhS8iuCSNg69x5KOUtaAw+ICbdRmkww1Gw6CoLdbyyhe93J9KQm5cDLhzfWHysT
R5XnGB4j3H6TVRXmhgpjejExOHrzLnl5ksG6vtB6v1OP+KOlUyIdf1jkA/rOttxP
95URe57yG3CdvMD0CVqMPagQXqeHGePJAVtyoqPxp0sJ4Qoh52aZIZbosUUNc2R8
nxZFDmJgHhlFSwlLBqzQ6sVQZFUazYrm7oDvLN2GWuwmmQ4y6c7dexmQUt01GpBA
+ZlEHGfh4cT1rf41yxkCOy6bwKP+0oRTChENz+jdAbabBKsBkrX9IhL1X0H5Z/t5
1GZORczcdiRWw7Q4h52kzthp+k9GoIs1eCnJS5ak9TqMOFZaMsKjmZNKIXxR+aDu
RYcyd0+oFzLKce7OGf8V+f3lEwAkGYwMgVvZusVBVGMjB1Cd0wJF9pfX4arFXwRF
kvDh0+C498LUpvM9uED83KtB/OfSoGJd9ApRDeTc+PQ/9IikuarNX/tddqAWJdOY
gXbZEWKhgAwmK9I51Eu5c/AoYq519yAKan2v4a+MItJPAR1lhj6vlTb3pj8rAQF0
Hb5iVX2W9QBPAq8q7RSLQw1NiA/VvEGhZTXMY3unSpEsj+XuAxEgLqwZkzm3pHm4
N0mGFIidTLaFuNPop+tBHX9P3Lw/6SahYvaJ5Obu2LD3P+zkALvw2RA5cEBQSa4l
YYWAbCknOPn1Qw6FS09wqIjYBUFi7Yj7q643zUmOXA/m9KdC/ea0hT2ICcWBiKAp
CzqoJhReUneZYW0rVIEyGcqoClYMz4GeblcTvckZvjlN1fxIdFBbYgBPzRac+oUW
ixXvizrQvFMHzWxthV/AQVsccmx3g4LbH8SXQ0vsu/A3/4vCGSsr0Vds8mo0Wdo0
Dpg9cYkn0p1/Xxfkt9c9MN2sGna/KnzTKQ5orwXV4lykOUpC+DE9N2vbdhbIvpfL
LaT84p+J6IhsYMpAX0XvFyLOOTZYXIvCXDOxWgP97CMiQ5lDoLZEJ88Dk6ukagM7
QdxsC85CTfOcrWMGz/42Ob/eHMDPVEAT3w4oeXOmYJpE1rYNR07AaxzNW+ZM/53I
YORJk+7/WaNj2fiPR/LHhOEHIy2tVbf4qJ53y+NWICqgwqH+koBl4xtXBsa6VyKp
nJM03muXwsfi+KDtwl3FZMJAXzuDSUVBiX9qtIJ10WY1vxN9w1FjkmwrIhsYPJY3
QcCLkXpfBffufNfEJacre3pGDFmq86ZPSVouRFcXDRhviUM8p6EnzkT3VcnMd8ao
csw2p1cUAIA3o+yyARP0CXsnCzABWp/PqBrX4UVAQf5kGp34PXz7EimIQt5NxO9S
AOo8X63dAc5u+TuiqhYeRkxvhHX+dP2keO1Sa9+0SpjnWahDBqmtqh32w6BskjFH
1Q+9r36utpBi6jZf1ChNMOpWbk3W2pbe3WzVwi9ttF6C7GFYci42HDlbmtxFM70Z
N/UXlrW+8elQXUqMlcaVIV8cuIkAjCh5dFr8PLVWrlBbxI/JZi0Ofj5FlmqG1TkP
g+edQc6r+FZF9vmPqedhKgqSTuM+dDucMLzQ+r1pTgwNWGD7u+fzI6Rjd3jhIzeW
dqv7lBjInsMk3LPuLoBSQ+WSdyKPkd7Nso3GtA55Qlo/5p/BbLN/72PvNsCuNKFA
ETZlM745IKWjw4gCyJWgAzayGLyoW2t/fJuUrPZ0dGXmvr2fz1uvaA4MrpNZle+/
AsDyAZY6FdKpq+ffFP0FpChIHPmPvMgvcnaCw85cRqLZKdMahe3hd7kRCHySQSRB
fFJZ2XY8RXSSFyhvmXDBBocqR/9jUvZ2kcJzJM+tE2sOW3284B7kHROQA7TKiZrt
7hRvoGivRRwabCvPcd1XlwxzryPOHo4YD2+ysDWyMt1HiJ3e09S7MHYiNzyZ+N0w
O9876pmyKqspbpoOj8dlp4Ts+ED1mIzuFcFH67dgAS0QQSuoEaysst/QosAZrvjQ
ZlIlz/ruQwX23571qJP8fRGitGesqpxlAYBO8jzf72WEsp25l8rQQwb3eo+gTtKu
9+YRhC62HiuIvaYAz+W58olFq3vGguoVprPpMD9CdT3kGH7PM/bOBEVFURuaMNUF
mObQe0x6TiW2ggksf6PqLEosMf4uppLIQimClM1Bm0E9x6IT6LWWZqpomx9UAYGP
eABrWAmD6i8tZfil1xnGk8Av3Yc64Y0X7JV8ry26qU8YFhj4WJ+wWsGohJUfZYm8
9Tsd67isBzPUb6NK59fic1FA2I70K4TIDUpd6fvoDZqbJq1to1jwS8OBgYZ/vnxY
b2FhDxZ0xfzfswSgXloLITkS9UhcVn/p8YbuBGyV8zbuZcUCyilk6h2bSSr54lNW
VigIW35J6w7TkLL50oV6G1HpCnGcwhqvvn3J5onPkHqko9WW9GS8+Frwj0AedcVz
XZdSjn6/cqInVS7klpQHlKHKq1CeXodUUyPNcZYQgdUZJfekgp2zgWHayDxDdQmw
6+RsqAmv2AdgdEuSjIXdq8j5Yu9p6dIUQvxpeimv8W3T3Q0ZBxpd+w7a6YvaBt2T
qSgTrxlyb2W9GdN1/0mj8iKpQUYxz8fmkGJkB7KMQPpHsYpRrxpwuWGSjUTsm2qx
HfOA53sZHj2oWCGgZbBHlmu40zWN86TtCh+puqE8di5oX2X3JpzsxzGJ+CGgn8l3
/u2OnGFEkyP9qUgT0fpyQ7jc6sQGbGZP40/rWDHB08soS1zfLXmkSg7PLyFVPjzU
qU9Hxsl+SKn+mZLpMyPR5qD34Wwnkw42Vb4aOHe0bF78CrqZPelSxck2Kizrl1sS
3lOzREeofB5I+eEBJYsz+ucuRFmvCfjKIdGumOEwjKDPn2getS7MUlZTShpWo8QV
dNhkL76bxjSpI5vro8oD14j7qSGBosyyvtuvRa+wZxol4As1C39Rtbye5Ane3a9G
puKzEM6tcn4jBD9I8fZRACbwzi6QFOR/2BU/5InVR1IwznVmYkPx2Ys+FPiCLKbD
xmiMI3iqpExa0ir67elNNy7grkB64dmwrg8MKvWcKoznet9HU+TqUm9mdECuNL4K
25GNiers6vwVkexl3Hj5hgEAZFDO9Ut86kElfVGogh/zsZszU79lXIl1/TakDJNw
qYA9AogirvP3H7FxDurnvheeD+NsVYfm+m4L+m+Egx1sxYEyMPHG/zR/MRrMEPG/
CK2SI9ExOUpU4tLlF1hC5K3D+KzM2i4XZ4b6I+H7T1nn/Pukk/2Z0FLm4Otw1ZGF
JStwte7L1dNIhil+8ta82IkliaqDIcxipidUYyTtV9FqEGqT5xNKg+j/wkU3aNz0
IKls8HFglPXe2wO8E5b/y9E0yLq/fnZufB/p18tAR7C+5Ooo/9gPlbYn9PToWeJD
OVZlFna2w7aC+dQzfEr6wOKheGu6kKMu0zWgBzCYCqxF4cx3IqG+SJkNGelLNFQB
QV31cDhn8Jws8aqfkVn9l9ABWk/FvwVHNSRbD0MFzWJjddwLJy7AWh/mVL1d3aI/
Y06w5T5uyFt3Ki88uZNBWldMjgZ4LmZtX4VM3lVcXSxzFSTYNeMxDoaqzkfVP4ic
Hhe/ekbxai5aDfh6CUUhdHQ+DRRSqnAaUX9YbqWvBEQwIG9LmK6Mug/VU/fI99Kp
zNNumoOMPSso7IqY+UmM0LwOpA9iROZYsBbT7+FYI/dBH5vn+t9tzOnBY2+amBcP
pqEEEJuF2cu8n0e/QrUl63eJFPhXfZa+Rl5vBVEsL4p1jn027aKfvoiyvtZkJ/7s
nAdSam/emwMXpUQGqZQlkUiBaB2L7JbhLxlaBEobqsxG3zNp0084x178sgSzE4vE
ztzwWbDF7q61n8zIc3iFhFQ0NJSPQSiYc94esiY/vqAZhj3Q9YAlo8vUgWSmenly
7sfYUMfDkJCM9MGA9mZpVldTbUtY/Vg/2DsF+EXkB7Q0RRA10IfKp8zyIn8NFWfS
BMlspr6EMf1ba3RO2oiF9WtDKVXLHGrr6Ufcvta96bqbjitjkqYmG4Qk0ENIBKXx
heFE3O8KGl5BwAjsJXPGY0kqti6QG1qSujBQ0RaBJehbQ2HEgK/HvQZG3LOYpKTh
ZekdSkNk+6CLJKdDzm6vKvzt7D9Lz/8QyCnke/3hPo1uwJ3cDAbIy3eUhkdE3qQb
U4Ou9iG0el0i3SZe8JqUODtl4PCNFs6UU3rm8IVGa21bUTEM2V3UvgD7RUXrRgb8
4419DP86GqsM84UeX1g+qsrwfKeOfIG8MN+cFdWDNzsOOvIUzwkN5F7SaUBxI9Di
e2m98T6Om7fHbu4am2MBtQOVRTFLFw6xUEaxWD3McFmafK/zHAU6obVQ7d8omH4Z
Yvo1489KQUm15XhD0yLoW8GJXPRl9ROKCL2NMameix0BAgOz845fdybXV2+ts/bH
p70NFj0WWhDHqDOkcnRtMIJCa7GzuPQOmbtyKsL4N1bPyCQm0/KdY96Jeqem0qcS
AicL/KOjFeb8rjSnPZhbll4c+B/Haw+5/MTvxiO3vo4RYpNUkq243XY2+f1nfhik
DG/fXvd8wBdAiKPkhQxKEVfHCsZsLF8g+d+slKw5PZQrimusM/ZZN/YN9ghW6THG
470Nz3JrZpKgPiHevlrA0PyQtp6hmlTn/om+TNJ+Y3PhXsn5r6spr6td6Qeh7tDR
0yMquCnPvJFXRWmfofOCaYd+//nf/32FNlvIeYTby0EhHzbDblQ5Sek5NWjm+ttU
Kuf6I+9hiGSZfwqWWh7f6oEhyFoYQxYeG+Km08AGvYHJ3nh9xwNkqDqj/blNbrER
3I9Qhn2u7INv/7EGSDX+RyQrAtYrEFTKAM0zcZjCk0k/I9ziLD4U501EsUKXrIs0
J1LvzCeSgiL8idie8YdqkP01pI/zPgbAYiQZif8o07W5nHRXaBRnpUQ4u6XvQEVP
ZyoKktt6RsA0xhd8Vj7zbtpotWgGXZh/NehC9bw/ZYI44JCj+GfDUz9N8+BWrU2n
n/t73/NLBZe9HCJEkZkyWWYcK/SPPXHgxtHONRNyhnESL/aIJRWMZapHVUin6pJb
RaBMOI87cSJoA2uxhEYhhFrRqZIwsDngvF878+zhzavl7b4p/D57vnpjDUeR1K64
wUMUfNBSWCAHaxlKcxh/ApLsKx1pnPMwhfT7r0IySg0S5hQ0soer7S4PYFVdrA9j
c5+xd3Iq651/Jud/diL1IAJnXWa3pX+FrbT3wLPYJG7Lm5CmPngLVMGQKa/XqPOd
8SNI1Vkn++cNTMo7wIVcK4ozqibwqgiV3TdPLshEiCJ8sM9jI1qUieR+Xm5hlTri
d++kiyksbisuobIKOkuIeSjyo24i2v7Vvy9bqf5U8JOlmKGWYtgI0FMOF7iv1QQ5
bAO4vhZl6g1Y6op8SpogU/6M1jvRHxhKcsUmqSxifnWJWEkZTPuWmW5IRpOwJzEh
oGoK6OaYELZwqYVDaLosnsb6enq+JFENAO75ilMflMDPhU9Pzof7AnO6E5OxJysM
JG4C0l4zzkqDtHUjaPksy78p8ZQM0nJUt1Nchs2W3cBUw4tOMMNRuIcGd8vqhHBn
Sl7Mj2XkMgQcavMbJaSiNXw4uuFWY59FnhDmdz73bpoNrpXjKsIstuXnyD25Sa7V
mabjyZhlqK9pfyT3o9/wSAw5bxAs4u/B9Uqbq6XSCHHqVxnIqe3CWDaRzMBUg5Tv
3rpvnk4Kj0z/qGGCJ26zM9QEIU19Uu8ghRwe0huUG8n/byyWY+oz44RqfhIFuoyJ
UGAS3kk/1+Jk08QcS5QM3rpaFCo95mdflLxtgzpoZ8P8EifmW2AhWSo2aVdpV2Ih
YyFVDIJQek59HeEWAj/hLuckxdvWefMSxxAoS4H0ELidiYhd4gLP5FlI8C7jhrEK
Q6SE7xDeq95plysQvYPQnGkW8+/wwDDshqyW8Wj5LyNLIlZ/RYp+NCzkTzL3hAQu
N+l4q2/ZcOT86XlKtS1W0Rwzun3R2d612z80X6nBWGszQJ3MoKRSWXBTBaV3lJf5
vE+J1386XJw4uHjF0OAyTUsVUzK/Wj0UB5JvdnPhsAUnm/wm2ISD1pUwx2YvaeC2
7e6fu2DMvnCKR1Pb7bABbiCRkIIHcpHDL0cd/f7U2XfhEaWyC4G5mmyk0fGPy+1H
83RcIEbw+80eWwdeT8AGT1/3y8k5iYOnbk5YeT/J5cnpKtRkII1wwe0LUWIBuijX
f6h78lute//bF1ZnBTq80f9iwVqN8VK4JUpQZWzWFIUVtshS22dtVpwCRrlH7YJ0
HGajVgesRp3jzCIwSxld9CPoTc6wRnzmdxERCJhTf0ILxqWqpFopDM7ZDABPTHAU
nCoqNIV3hIO4filyACZm6RwMnb2D1sIzaLXtOMgSsSpNmAw9prM1ijB/dfxSl0ka
LMbd+Sn8CjD2ZflOgqU6L1Ve4kGtNgIfNEF8Cpgmr3YNJzmFi5/VnrFwm0Phy1FV
d5YS/cwlB2EUSWnElB2B+TrL8f6TPPWWbTGd1vDkHN9Iw40bWwVgVpJnVhRLOxJ2
FyVzrs/8rdm/l4MeOuF/umdb2s+9sASX5VW8P3n/d1BTHrJ+QNP4aLVOtp1NwU0q
FiBl+jcx+tmeiKYPCQA7wCDa0fJZrm0RV4Vq8gXXnjefJMFg2gWxpOOW4Kofu1yj
iU2JnuyLyy23dKi087X3kJd6AKpDSF9JsmEzUNf+gK3J+kOaHtQ51tXVSXv9xlgz
hzSbwL/5goA364r5wTkak78HKeYooxgf0+AUcqaJw24yltGa3+QzOMgmxVowW/Mr
qHEeVi0STt1pL9GOXQtk60Ib+hGdSkPdizBmpC7U6B+QPfomR/I78ihOZxErd+Iv
H4oasZ8zl4Jm1BEcuPpnDr380dtPS9h14Lk26LBVOL1O7ZIgZ0Rj7JoGM6QMc4xk
+6RtFV0CExpRms1WlwmDO0+u8WmUU4HmvoGes6+zx4PZ2yfQ6trlDTjnKUCv1qI/
+waqmuvHpeVEPHfysM4XaGOYCwnaG8OuTfdUO/2TEfIERtNln/tNDPguu7HYDgA7
9tr4kWbaXjARREMZ9dUf9BwUDZC7g9trD9AfEXv+K63WqUk/ApJfpnU75f/IGbKK
wfXaW8F2kYByKD9SyjlVUfvVETXX/qW95NJBwZdsRDFJFfK2K25f6JSvqSiIo2cg
z2f+4s1J3bfdxUhGd6qxUTaMDFn9e4LKSgtzafNmAqAd/dyKYxeoJ2zC//JCTAeW
6VaIs4Kt7qSczjSx1/SsE2UlYMvQ3g18foIuYS73lTNU8EAusvSJSxGKMw0Br1HX
O6C9IFXKlv8T/TL/hLXOjGxRpvOxA4xJeDvx7wXH5RV6STLJAlhNTeCwkrgHLiIB
QqU8tXQ/+gvzQI2R6fOTBnviwDWifzhnhyvdTl5ZW+ii2hyi50hWA1iglRGckko4
AuEVrd0hcm3zZSJlOVFtFOD5s6jEh3wI7oTb4p9H+ZQNGzlSmEhuS1GSN3m5rk2y
6atABRKzUC1QHirqqyGdcMarh5M1MueJluLSb3M61M0iQ51VtO3IZkv/l2qOitcs
Fvq7cj+hrQ508wTCi18T8P6ypQJVgN1f+4goMBJ2PzFFWyqD5vz5qM583iDKtvEM
23iRKihCLAmtccZMi2mAxkKmUXZSUox10SoRNNegncCu6XFOGCja4J4YMr2BPxNt
9FYuzyNyAS7PV2ya6POuS+8XxUa5HEat4Q0u9SyEdBMEvbTGYtmNEivI96G0VGHx
0q2B1Ilc7JRRuclbig/XSwDBSEJ5Yw63hCwxnPwrdiyF21kld540Fux8MlChlVCR
A4AMACExZcwKJrsNrhcnEK31WER4PGKKnzMK+KZSQU9Bnv5GjTiScdlXfVWb9kyq
v2zDNc3m49Ge2W68+LIJvCWu7+hJEO5MWaTclwpzHwpb3oJ1JBFkngpSVq+LkO8o
v+8zWTnFd8TBxxsZ6MoBSj73+PwOuFgsm2ELXPZk4qALUQk1cbXpmUJHAyw/JVXm
NbRXGHKQ76whjRc3LAyTn2aJgPEOWq7rZvw/5ltR0swWUGmD5y1ggVPdBpl5083Y
QrVSU1hrRXXDfgAztnAPd8485RUxvqExrtIJQE6+Bc8TxOJCAYy1up3LYzNVIdeh
C25orqOqYjNP9wc7SI+QtFjq8TxQ53NtnMUpkH9q6V8qAijF1zyT7CoQx2KbKwzR
ftriGfFyWygoRPOFBKAFm8SrP3yTRRf8WMfRrLy4I0IKrjRPcM0QA+sOpV4Fq7K/
VUo+uR2x9/pW3G8Jb21wKIBnhrd1OTkQBdrDtdaQuV7JYnwSHnmwgYlTFtR08Qpu
EQiCZ3+G7YVkPulEaa+BLrHqRp+5tZaXs7sRmpWXeOSKcyixy4xmGRhl9Qh5zHLv
GrZ1oFY8PXGGtS2ON9L00oN41NVfrJmqyShg0DcLjPyD5mboGMvfnkfxzQwTTHb1
ZRf5PfuppM1dRwc5SL7Y2fusHbCYWuzS6HwYFN1mDWN5RQtNmLS6vIptxglEtVXs
rjoq8SvQ6+51BTg6tpFntOR6iB5+rtbULvS/L0W//GduzrelSMCSx7uR+G19Lnwe
tRfKW0YrITYoUnzr/auprAxj9kDC4RSzEEBX4qHe6Q0Rvhds3NF0fdk1HZwMAM2x
Nit/blvb2avX8VYmILOkC+VXA05hoUixh2LErC6DnBLFgCokAOdvsfd3hDjYdGhV
qXkqOqjnDOFn0SFN4JsdG4Lsm6CCi8Jthl5wucb8jFEtNRirQa74EjJEpmaE75q6
jpnNwqWsuBeJbIEusT0ivcg3rFjMnd2HanACWYWJy6tq3lSD8j1gLfh/buWqa1wX
sS9+mZ8P3msUU/hALcdSMQ3+k5FHjqx4NgSp6ioXYmNkf3WNklEA7qr9l7P1Qo84
H/ULTieadZrueh8Q3AOWJoHpeJJjBygvUorJQkrjo/WvKyvpo6t4mtV812y7elH6
Mfjmiu5dDAysYBgwYE4HN+0jb535qYB+v97mZCwQ1gVO9jM/CQm/sRAlD5Z0DztN
VzVbIKeZQxw4R6GKPg1YznNl2ZV3JnDQyEl1KUx50uHxD0POTOB+mTy3a190O2Ph
DPeQdPnnyvcFfskEuH96071UieUBHQ9OEpNKKhSNEZq9chHjPG6cd7ZLJdw0/2zO
BZ0ecfD1RYa8WnzUt/jV7jqSf70TqbtpGcsPeCtLrjeN9zyt1PnE+8nYIO0HPoGm
dkK7LfJH1h2JYTr3vHtINke/dWQeQVvNgz4geV1gXvsGxXS1cOUTpfvO430eXj43
VpKiivd3bfg3VA9KltDama2tgZP+dwkKMbzFx98ADDEU3PQGIMNEjrcl9D4KeHYM
Rm9GmmcHtBZM8nm61UZ+xTfKsOvBNzL1Rm1Yk5WVt78j/mP9v97HB1MlM0S6pSwS
0V2brKrYNRbOAKaOHA/f92/L49E8b6kpM0p+uw/LaX8P6DpbB55VuUSyXPWZY/YE
1txlplBjfJtw6XSbvzFOq8t1z9MpHKUCG6aryavmVHIDagS9OMiq6JWRrbyxT3LD
KxJnzlG4XxpmhdrQqQkyRGSWg2CoKeC30vLiwbBHGRqWcWzqn/xxa+9vTH+7lqQF
+J51e4J294LIb6qBvggD9K6lGZqhskq4THcRGHjlwLtPVuBuXEz7phdyFO+XYxkF
c2HOpSdSSXxTWTCIYgGvCi6Pw03i+r+Rr/AtM3EenDx3TJ82gx+a3wWw4dgPA9El
rNleXb/SrEFYiTjXDXSbD/rwdSspWPG6HbxGXrW12noypNWICbN7t7MYAWrsJmBZ
g5Cw+2zDEjzdMyKrrbV5kJJi2mUVREwJYxxwB5cJtfzyY4ZiTBZCoGUkxBxTSc+v
p0NY2CSrNcWN65JlpD3i8kYTlruTq3hC3TLa8JjCQmux7OAUKWsjBe5xcLVFYBYA
T9CRE61II8u/2fghpB5R+McizvvFtziT6zzBSkz1Szmv+dqOYrSUEgfhbEeoPwdj
UR1QdgJ5Nvuk9zA8OjSj2l1xFdKFIxyB/QM5rsY2WBBWsrB7MALVCiXJHWnv4427
6JpiZFxLQ+K/WBg2kwgtLEYRBmVO8wxs6F17gWDW/Y5EQqsGgJFvJCrrtuaEqas7
oxZ84WSZKc51CwbSor/mTABhLrURXZ8MnmbdRVhNtLV5Q2QGAq6+bMXi79XkhBsD
v/+kxfS7sUA8PA9PE1uaHRH9Jy4Mjw3qtSwZtqjdD8RJl/NY8mYM+UicU9MZBaiF
paJGmAiR2LdgwkCojwmDhaoeKq2IJDiGEnrmJMYLcWl0SnuUlBdXcYp7tTj42+9p
6iIZY1m+8XqnXRx3UpyahWSSV7MywgERUSqaVhMo27B+F7RCi2KMFw2MZYhK+6t/
gZC+SZeK9STy4Dj/L/yBltUgfRM0eseZLmElqGwmu0nmAyvyg1SoWqMEy72eyASi
mpseFefTOWFFybVUR/ssg+L+zrKw3BgkuUVbgKRa+Hxjm8WyXJaUeRd52RGWR2j+
X5BTJJFwMNhbrDsq6fdWFdESzbEqPfR2Wi0sqTFujdom8w6MxjTv7+9md2N63+xW
/k/YxBG9FpvPmSaPtE62NV7+3vfvOuYr1Wqs4Ahr2VV9QqEXb8VAEsBGH+vyI8Cu
w5ngYBINbzjk5lt9DHIG3iY8wIBGnanWjDy8XedekcEdWD/4fjc+tuF0IwSypK0k
gnfqo/u/5ErK+ds4RRIQ5Xqtfyxsjvf/aKPh2HmqKRyuCVk0ATDX1I0UDkLCNnIr
WY3jQae1mfEfK7VYgvLBIX0S+VcI6Spy0E/PTHugfmcvzcxFTsSaO7i9XCupkGV5
0xk3DgYOWfJNzakP4AX8CcqSX02lTh8KeyuBf0npds9Y6li8U9Vm5G6Ez6EP+1IR
wmHmvoFVuKw0iSldtomC4KAE/Wj99gqoXHkfmlWyvOyk2OUjzgljvYagDqNsjuhE
1fLcIjmdncZimAjzNxOq+XjTlmLE45rRFmToYldtR/MJU0SaNrciblEug3pEdnzG
RB91qlBYCzW2HJ+oIy6SGE2s/bXA9W++Z/o1x6PwuURtTXQtTXZGLzPe+qNfxSgw
TgFXjcorgKIrm8lIr7KlnJ7egQVeOkOaLO9e/XQfCfQ3zHaqn9BDx3iK30zU3xpu
hs4Z+afYaBX3bDHhhzUTOBTKEEwuOm44xkP9d8NWOPfWeSCziXcpZuoZPViaqVsq
8oC/QKp/Otlq9u18Q79VgdRTv2lcSAgk+bnZfiuXa6xsoabC44Z/9AvvUvg3vBjO
dfIubGLjkoU424oC0VsqrI/3jOCs515FR7CHr7hzPYDmVDcalKVBpfbqqTdtXpKM
GIQiHVb9dW7Ebmm6NcmpBVkE5oI+Af7elG1WlvyCjjnD27MZAKMGmItPgelyOi8T
cgU5aaKV+Deo6hsVvblpZoEeHqU4M/g8TXTixANNQnmtP0xHcF29NiKVsCgx4X6+
S9hJhuGQVStmm8SQT+piRFabBMTHAHro+cwFmX1wkWtyiF/C3f5T2f+f8CgZp429
sQsFZJXjDizGTYp/LPPbSSwDz00RdZNEmrq7VmDykz0U9wB/jCWXa3ZUoaN9XSsY
J/524lEU3pBJ6ik4BZvQ+2S1C3RSEmnFHamtJ3rs7GjcNm/ZJFtLgZ/9mB7iQOKA
WqbDsXWzeaF7HyV9yzG6V9V87zRE5hJ9LXqriD6ha9FaeL8wc6J14xL0Z3Y5O8Zm
2qEtbCW/O1NoOkyTEzNaDkPht73zlkFaHEaLfxTinBoH7I6JTkzZnMsW8PDK9g64
8GImKmR/hJLNNS6KaagBjGHSiJLAdQ5cwk8z9AVYqXlC5XYhwkh1adMhhFyR9EhX
Iebc164Qa3KIpXgQ7Tz9PE+GImKF5LtSWFq4awRuBS0+bwE7ynd4GogixNMS2dC8
uVgpPC8+nVtIBwEcys+ZS1N9iDlaqm9WLjscWAIRqS9ZkRcCdbKgiefmFbdVNnDY
Bh2vg58vRUshG1dH0A6LSioN99r99Ad/nbQuEHs5sNS1uyiOrYvkZgOC6Z5mSqo1
xNqwmkQIthWQu5wtn8fMYL1UhuM4whooW10wFXe9d+RrGSYOfJuJVtSvliVj5hsX
Cdd54lDlNeRghLa+AYgorcU27IqmelC5oKAtYnL0g1Uvn2/I1sChXuEtXoTsssVq
UZp3JyjP734/LP9ijevlv20r8B7nZxVwUK/wVAW7SfuP2zxOgSgjtp+o7sO/9DNk
2IfHoykpd/QdVhAoWzkAaIje/h7l4wV+LPKlcLAuyuSPZlLBrJ3ZfZosXXmDlK25
eUnC7TYlwl7yJ/2p0IgKjbdKyYdCa5KCdaBd6HkNFqWnw92jaCIdP9sNImlEAxTu
rZ7BbI7Q7MJ6plBYpYEbAGH4WIHymehZ8EmP+W6avEF8yo8dVVmL6X0Gvled1d0g
rEGWDI+gPXUQlPX9DMSNuPipTKArbQrIOrSAD3gh1Owo3/SEQGKRbY0onvbGlarQ
cmlHc1tXwaFzgGaR66ejuA1jKPdkvFsCWD8OcU+SEdF4dUVlkm8mo4bGzXw4at0Q
M5Ix89+fR0TQ6fJwTidlUBDCmRqxXOV0JpoUlC+r/1lADxCvvDdAJ4zZMvKeUcZa
uG1yjdU8SQs9ssPXV/zxmV6kmnFGoUraQUG5+rIk0RGSXJAzVCtmZzWvo06zzSfW
UtK717ywTLk7Bi1y/amhX7tr7X1M1IOgbU0lIwawhHZ5af8RQmdOKZ18tut90oWl
TggfegNwEk0xbWDX0b48MiobBOxxrpf58Y6mI+VoqM3OqKaOoyftZINrEm0q66wy
oNNaOsojagmcJEr+mzUQccOQrf2ik1aOmmDH+vJMZGO6FPMa7+m0QuhIi4hvcHHI
LvNFFZVWFzrvoSUnyr3DuRATmv933TgZg4R5hfYrotM3UvVVrDWHLZHgm/tAay8X
FEn8AGn7liAQNtmCi0DIBKhXV0EYXoHmAUmubC03C8bpXGtky+9gee/dY9C3YBqC
bcTJDxkd0ye1doc7bT+X/S1R1ZDWq9ZlqSEdgyEAwi4872WQfCJUM0bnT0wmMlZg
pUdQxvhlmQT7GSq2Eerj7SUch++vhZC/GN+VAPZftcJzb+xQ7jGky1V2rS9SAVgm
umFRcx09SplJ6nVhurvYazXQPcAAPXpxfwNtD9aTQxyYMTd82HlUhUK/+7ySPFGG
LOlGjAeNpzfEkLQHC6a7Xj7bu9sbfJqywnaDXIpjJvFfyiYTsuSQXii8TFyNLKo0
CUNbHien2ZeIhN6hbsYmmZ/XBjm/HGgcDxtaSFI5WbELbnjyR75PNI7tyPrBBsTi
QNbVuyP5k5JowbgsFiWV4TnQ7kIA0wc/DpslfMxbJw2HaFrshvx2V5YaqkTq+xja
6BGkfHmQaHp5RS4GZVAxL5MjS1tNqTXPKohlCsNz6MwUj/qJUXbTKXSOERuZyiBT
HAn+CLYz6POJsx2KKgtZzMn8tf9wL413+F53iemiyoQf6I89GNdnD08aiA6EABxc
UlysE+h4QO4fmDwMhOOJ3VHPTArK6NtvR6OxFhOeDA4Jogak5wuzd+At2Z+KF5WF
9aD8rjYC03Exk8QIXoe6SupLtRsf9Exw67p2vdH43eTbOwlVjqnOcdOQfVeSNDg5
SbGVs4hMADZwWCGoT4RPdc0BI1J+zUGqXyrbgbzJK2gY7E/ggtF6ufWJB+ZNvdAq
6B4bQE4JsTijj0YNCRe1tgw/7ixORqClIUWpZVLuvF1/4hqvm0CeIZCxkW/5EH0N
NTVQ4hVYfBqFgdckDd4g7fFSdQklZhO9v3qfV3BoWnW1l2EXehwCAkS17LXxSusT
TFRtfJS1iPbM6GdR+IB8QptFIW66Ud/3yAtcMopCirqS8dy4FazAwL0FU7W4wx+2
nrSGPenwhQtK78ibCvcnXgenkS1noZcYi0Tl3bl3BCcapohJXqGS+24vxjjYprKd
ByIFjsZTJpZL8CSraPEUVpWydy2eyp6TX6T9nQKA2T0jYGKxWenkqoGQEIcZHwR3
DkrmvMQLKRNtjG0XOtbM8xPhQaura0keUQ8PoXszC0u+xdsty/o3PLMBds49tX/R
kWyDMxRGB89quQoRNreuwqe5ZWZocnhMtVy+qVaHzHbOyGmrbR3A8QrJczYH6bb1
fn1KT6DjH+b74n5EAP1URSvGAcvTQkJT9hhp4Zb5U9IdkwhOQfdEWSxayhjpgbr7
/B9bDRooVJi8jEtagSMQNmHuv36etJfwEImgz6OC24lgneU7WzBlnb91cEKoEVtI
QfZpaw/E2tGV1Vh7eeb3fu/UVran2w3wNVZ0r7n/31ii57tKOuO1TWUEnNfxAD0F
awpjx7JrBfAf5G4l5JqIeQopvscdu6xg0UMMMiv8PNlC0JqT5+X054AMq7w+JhMz
7CJjxyTH2OxT1d86fGqoie+Xs8A30HogwQ9oqyhUhN6LBWe420HN5Wv2C48ASwCR
TZpHa45f0zaJJFfTo6nswWmRVZKYdgqCeriEEjosE8zB6uA29iJ1+H7YoOYrlXZh
vSHfIM45SGbLUj60zI15IyAaceaei4eyLpFK1jpqDNhlhtZo7byuRXTcPtmeENIR
LTtYHsZrxBIit0l24+pbtu6kinLbui+PSeO9sdPKsBz5G7yxo1XRkTGBrxDQjeoP
8ZLCleKEo7UNDREttWSkKvc1yAzYO8Avs+gkSz6dU57YyVlZBxJAtHTpF5sLW7Xw
XFxLRK3/DaZ6hmqcCyjSHU+vKnI3grBaLh1jkvJrsUlTV6gBshQuixYTKaB3NvoU
Xh0+dIc4Du5E4Cr70YXINmnJwXta2aMGg3CBRSMKu+d3iPQRYyDjyGaS3ZMj9eVI
tqI5TcHq1ifIn/qVWQm8heKIrLjXe35vkefbdPKswMtxhGJsN+8Naahpr9qfW40y
cVscNFsO/50RZISv53ALYCTaaNkAjj/nm0W73sSt8Czn56Rzwy2g1nuzVwnTRWap
RlTqqz6RbSbD0CfJUYRxPj07oST0I6XHOyN7s/3tJHi4LzCnVRN1M+1NJqc7YJVd
ufBaAAX7UZGTP/286c3yI15gtB/HyXU5mJBZ91OlZWfZ1an+NhlJk4S82zAEu58E
RkQNPxCvlt9cCExahJFPay1bwyAXP6zEWTvPUh7x0/8aEtCPGmRSDtsDHMSQYYC0
t3J12INhGAO/SkJRF90jNrBg77Oec1N4fMfGOA2YSOxoTFgqtXWAv+dbqasE6J5J
cxwSrfzijHbrPdpsLc9wppxzWlt8nfi2oJsh5SYSSHqCowLC3nA9S/vKy1giPrkO
grjxYIE4GM6QRR9Hz1pOU6/fFoZkd64puMOf/MjZdWwwHFJiFI1Q5WYyw7UKK8Jl
4Ml55oScA9cSsIeoPrJdKUtRkguvSf69kFlvzszz0M9jwdiMjBs68gzVETN4Hoe0
nIYW3tzgAEThVzU763sK4vSNdmj2Hii1dRHQgLM6zLatwAwWONCP2zQXRzXKuDGx
3xNF5usyro1zDTk1kYFLI/NADDYpNf+63UnuLvn6RLG5eZvrlo06RszXto31oFgT
B9UBaTZypUJnbRkRHuz8vODSUg8/qtJv8Egh6XnAceabypzJ8UpHjNhYTXVMu51N
00U2OIwkv2unetibPxDKs4ahSUAJTm2okwMxZ0XMbi15G/FiTjZ0Oy6yrfEbFD0J
n3yUv8DgxBUvPZI9+TmDmVr2RxX54iuluOA+bUeIkUYCx9SiEOKDz78ozUzyk453
smHpBVKmdMBB/1LVgmx1hFXBS7fUcqh6R31YOtRiosGlVg9havbJ0N/3bPQG1PIK
mRBODubSzyn3KqR9XZoQFzolE4IvD9w+8a5E29jvl/4rwUrGhvEpprHI684t8ZPR
ePIAY1CVBSPTKJOVlhMNXqbnmzkRX2RR1zjgw6RUKcHoM9vg0AL1Pl0PP/S1LvPE
2MmbUwG116offM2R/Vqtgwlf9/Jr3AhnjEoDXwiwWnCte9tSoc3zgG7P9n5eC/v1
h0u5rxrEbv7wPS6N/HUr/lJf1n1HPb6Ti9BZcsiYTpB1qU/9Qd3CnVy6PRrKI/yz
9eIFgLqJoDm11dktAFD+9XfxqCZhMec40PeUKdrD1yeOtEX6I7Dsi/PgJ0eUYqF6
5cNZn1Ahgs7ZJJjeDtV4Ihkf6WCm7hDfaxqQCb15p0S8zd+mtrjQXBcj13oemLBu
B7FmLsZAcKmVGJUacKkqagIcZ5S7m7fSjyqzmzLiNljK97O9+kTeWDh+SmDvo5bk
lT6pAO61+TDJZJQ0gmdOUgaA9nZf5x+LYsMAq9LH7YTld93d2hXG5jdtdfxRc/5b
TepOVWPV1y+0haZDiDtJWJatRJGtlerMSEH8xi5/0JvMqGyH/gGYnNRyBxAkH/4C
p/TCFqA35SlXJeU43NUZ7G/jhCesWofXVh7CNgxvN4j0TQbi2/hh1GV/mOIEZb2C
8l6p6EVxZ/vZlrfqOKNIMV0tZEqOEHt115V+qr0wWiotEECcs+UwnSu8mS9JKO72
l+pUwuRSlc4Sumv8BV7FiTTI2pUrj1BnIrKMmo9TlW56u40srZU5tnO5gjGrCuy9
7RY4zhFafKhaJlE9Ip/leCkGdOimwa5x+StRJ0CVWSyO8MpK3Qvg1/YBAWjLZVBd
jlIov6h4g2VD3VevqFpjhRIEXni7aP0n9LUyOW1EQ8ZoBQ7iR+iXolpQtHDhLqqm
ioSqxGySoCPzZ8wGYODaRvpETLaQhCF36l0zJf37YWDK7NMPjNuX38+KjEDQNMnH
3Ov/0OitydqCdBlqcrD288xBbvUQOOy/QfBHGUoXAz9wY9vnzP+P8n26CYeAohmS
zlPh+jDpmjLzompw5qnI2QGxfitjgOimY1gTWXbrNhYNfScQ5yxzt0y3Xc4rc1aV
09zIHKK2RtTxubqG1istHiONN/kM0ozP8wjj8Uh4zOjvo6vFh+tQOc3uxesk5I/b
6Mf/HSI3XDowkJwE8Pn2OXuNHz4RLIscNTDe4F7LfzLbntQWmSrzeSmr6I7I9mx/
WdxQPAuaho3Axf+SFpk8JEWUqeqeiTkZ1iVs5ojAZD7D0WxLMbVkrwi/4RH0UuN6
t44c5SuWQUKMYU4F3AA/ce301uIzA6kZirLSgJWtG1ULI88e/G6OfG/dzOxrdmX+
F3VPyc4lfqPa24xjCs4Zrd+vye7Zx4+Gu/UiCCYdX8cbo/3wOgOqFndbWhbWxY0t
fh9kTz766lbeUSuJ6GPKPs7LZNwGgJsJMmtgCQZuhb31vbRtaD1obJaJdAMqy2nE
NFf4cd1JtmQSC1Jb0h9S3294DPnApgdhQo+W/cBHSbEvsxVtyE/aDKk0ET82fccm
rUv77z6M+NmNc+v5IjqKEqIH5Sal1Z2Gq0nwTOoUiLlnN/lk3inR8rDUqq7nbrHe
6zlc424gpgIXCJMFWQRwpSS8Gnnu4NAfRsXhXcbicisVJDZXtXGiut52KK1eU6v0
M4tJhcKJVGuklTRjtpVwL/uaDaBDpGZVci/uVV1+vYnNBXhDSJ/vWVIvNzzIcoiA
UTVgOBu4csMQn94xwPcvwyvkvPp9JUbPHykRqw6blVqjKVYD/ORgyJ06xLbqf1qi
6RSQ1q7nDudGajAdk+F3vN6XmKM6NUccsrlc/njJkDCnCFDeVUilLz/SbriZytez
dqDcAgWgjSM9TEn5kzePSj6Oa+PG//djVZ9+x4/mgrzV539Evl5NzI+zdGhTdXxq
+h1mN2WSqSrs/hSnG23fPuFePCq9UBWWUKqipqV4VgWmhE+nL2V++XHOM/eZ7tE0
DUXtpkmOhO8LGCHeOkClpGAaQ9HMDmmbxBnfQA/5njMeDfkE6b3nv6Wkqa9c3rie
85cgCHYa55KnMmlJeBiJaBv/eCZqG4BhyTA5/wZeo/wCgWHZBT4xaf02NoEY8l9b
kvRwpBd8DCWCv0eiHcG7WPQy33znHseBo9UZge3P2K/LmbFuVW5opBMo7PmhzPQJ
gUeNKr8GcUOIUMxVLqjM3JJaAZCnhW0X4pa6B4XMXTQ/UEFGY60pdyqSb2Vk/mea
b4JktcwwecRiiC1dXOOI3199oOqOvD2/rQDUKCGKWfOEUaCotdyNdiIUSyR6vQi7
NjSwj6dmwpAE38IGWUfOO6/ngvIwNnVpAi52RaDSdBIKAetrXak6gXhz0kPEIp41
krJD0fhsEE50I+bZ14C2xsugUWN/01ASOdWNwPHkVa27BHfpO5jGfUVp8at34hse
xb/i/gkn/1o256vt++ySDTOKFMXErismZSebOXUc6bjDFadgY/jqrGMiWUMI1WYL
v3yxoev7r8jxMK7mGQ3R+wxS44zvwRTJIF4vfGJ+T+y46llStpKJ0xCeSZV0NhAY
/1MeoBqXoMgw3PzxIp5PIz89/MgTIHeIkSXEz9rMJnqbucrgv8HDWEQwhYOvaaA+
wU/UEyD32AsaiUcPkkou7mCMK2i+iiozGrxHHBst9F4LvYzncmCmPd3WWMPoUNos
s53KQoTAw7yFPrm84SLhriGWase6IHugoAI47crIyFuWYhhsWzAqQ57JJ5ccLpvN
IS+E44J+wWWbNvKX9jOnzrk2m6aRcG7ONm49zoo4lN6WqJa5odIi33PtjkPrE8dU
hzWplaCdANHYFutFLvWtxhgxGMUhXsurCMmseC8jE0e5g7Co41GDoWlCXphz8dQk
QEojg8Rl4TQho/ghf0EuRFzac8/0mPbrsXXX6tnr6PNhRVNK697w1xzy55+K6uAt
Vaa/ymy7pf4cjMXUOO9rrWHl9CDTIMvoBnEjepmXXNRQImpj3jyyZJkZSWc/dKW3
15QkKEaVUTxLYV2NwwTEuiLNqb4PskDsTZJDM28hYmrspzrfql0+rODfTLgKtXGG
WuCXNF7OE3IrbZg9pZrqeD+T5wR8h1qpu5LZb1qsqibwcrgqyusxAUAI9kfN3+pq
k/4xjH3meE9ccnz/XGECK1l5JG6tw1g6k1aRbymEoJKB152p9X6eXOtjmzTrJz56
l7ENjFEAzI23AFaA6k2KYCR/ge5F9FaiJYTbtoFvmTqwff6ewfy7Cbuu0vkL7mOd
OxhL090OliPTcLnNsI34Go3sIv3MisLn6KFzNyVcO6R0pUtgb+2MA/H1kUPH6MT3
v+lfraxrAfRVm/nv5mMA7UOCFFt5qmiONVz0jXHj+q8FLzBITepAjVC/b3QCbXgF
wAqEBrU56MSl+vFE+Zn6EaslLs36D7SOj2VintDobRU+DKCUx5mvNtDKQ5YYnr5R
AY6TFrH8nCJRg7NrTnkASaQBxNXKuU2EAvShVbLcPKR6rqhiftAj3hDG//m1KvhE
Y6ITbpFoqom5PRITqw2TFjIwLy37Uttsin/yVXEXnbzvuxCBlhcFppNQgU+drJwy
NeZGfwvG5DN5gBtDA3ozQanOAmKUoxNi27+RLZd9IB06e8QGNUKpCtR47ihaP0FL
8eh2XYflp0UJZEJ89fCFauHctXDfe7oUfKfkZ3KMHuyHanMcAsbZK/7NWvWIXAkF
i4Rs5c7gDhAYIgV+xEM3m8ybDsiRXNJyF1MHRdjVWfYVO54Nu3iaodiHjWPTvrTB
fR2OMDPNuvSlke8fPhv/NSkoq/C+6EJQiDhPQK0InOytMZ5EL4fxriNNojVFCs1f
BcxYIHgYCM2Gr8lesyQg2xMoYfapkKSXU4FzN3JbGigjvyO8Mubgt/0jtKTekguu
gYvVOie1+mx9L7EElJAFwgiJ8Z0Iz6C6Z2s3BnsPtQDRx+96qikgJVSB24pH/OSx
V8Yke6W/wGwINp+am6Ticp8HqMvgi2pkayi2jJoEIM8COMVsRDdsDZRJsGJ6emOK
bCv8oVxXdtXUeVBVA7ZHxbuXOy76dUcldACH2SzdV0xQjBzr35ivm33KZNDPErtC
zQuAFnERTlBNdQRjgd1Q1nJuFe/CjSbId/hHyt0qJfHf+9sX28w1amTwqYeF7a1K
l6V5sPuJ2GHMwrhhei2XICVgFYMggvS3lZ2B7Cmd7uw/2iMKx9cu0mzEQMDsLXiy
8S78s4zgp6JGqFzPdLTE4ErU3RIX+6iMirchuumFsvKbRxSA4eYMH+rxDmOkHwbA
jwkYg6f2ey2GxAMXcEgMAD6VIWKFYZC7PEYGjVV8nsdktpzozBW3vjq5WJAAJaST
2h7Jxc7zJeLVrysdewPZzX2FGobwLVc/SuWbH9TZX9td5oFSMTmKIwr5tQ787Jm6
eScWNAH8M3diFWbJrhQRtExEGZ92au7I1Qh9CfG+7UeJLkhCv6buiAIPvTH0VCQ/
NPZmFLS2t8HiPfl403kGGTPC51iRj3s7YUtv5zyzUoiKO7K3TXFoc3LKsowO5AMQ
IAJi8pzkhYLzbeasK2QBWVNyFrCFTkboGDxMfEcrGaRdKdeeVdHQRNL8p/WUPUlw
T5+yTMrj6rz1OnUUDc5+G5espq/vJGTM+Qi9LP3vHqskcNOHt/pVhe2x9oSOQE/p
8gJxUUkBeIr8dZRf4KcpLf2HLWfOrb85tanQU5p/2qBzXCIHUBd5/o6XFvhvKhXE
PFlskjME8TB16ZJWadE0SoFjF64MMQrmcuwNefIWePzgb1Vrls4xwJl6U4q8o0Qx
0Rnaa7vo4s80QVnQzBkxEuJZ4mDHGtRK9s753jhAKvnuBXyD0JV0HhB1X7KcZfOB
/rq9aZD8nYSB0LUfOkp6e3YKe+udpFmQ9VhXCouT+60a8JjfaLcqjz4AU89Qe2j0
zA1o8x8dyG+JijAmfESnd3oZhxCT8451IW+/n+uKw8W10ezi6eXb+ELjfL/3HTaV
YxEgkUU2zGlYoiOX919Q/vGHfIU0HMix3jJDwYfOkajjG+TMHh7q2Zp5+zVoees8
aBrXg+nhawUBUIJ2QaNptRvVofmjCMQ21WHwjqt9BTMNL6jwwOKMGztHvXtByGHM
7piromQI+wixCWmplWj0ON/fiKCqG+GCq7dH0zSZpnUhepx6WC6LbDylCycR9pYI
02o4m39nqxa+bl0mjrJ0yWAFYqelpfye563nB9xg1nIjuFk4KOSCQrCX9azJWzOA
/nF8oG0IMOYGu7a2tOwGghUAeAl8ziScjdprIisas6+WqAS5306gT/0QwHFpmnN2
0yLJMp6tVbPEdFal9yY07zjPgpC+s+AXlUHVcDdkfCKoUScjPLX4q0aSImDU4AsC
gyZZ0WZGYEP8QnuuC7U5PWDPQIQz/HeRNi6pVK46H8EfCHgsNF+r1KXd1X0RzdHF
OgjoebkWnFSv+cDu7YRSopCLsaz6XIMTUDlcfFrXCLm79fmA15uxgCPxGSX9MoLk
kigmDR2Br0q+yHyu2oOatAM3vKRveOzVs0QLcoA9Ew4t+n6J/czmIkamlCYOe/m+
jlKDAJwp6RVwux8tQ/jG1u2SWxn34IiE7sXzYrRgr+xvm/0j+JM34dELXr7ywWKe
Ak0Zvo8HAzl26bFJXgmxRVqoiL1g/HZGd5qgd46f2yRWrxuxXb8pI3u+K3p/IyiR
zruhAE+Crm1ABlM36cUO3IkiJgMURfwqXVIkv2soGR+30ZVpv/KheqnGSFb1rUdE
8+Qx0ZyO6xO3xDnwq9fVijb5lWktCV2CLpMb5Gpvdtfwe9BeapYoUyd1EK5Kh7t1
RnD8xGefHiIgKtMgOG+pkF0OIYZAw5eJbURiv+M7sy2pvAozW1AYjF9B25/ExjBW
OvgrJH201qKFHtyPhK9NSMzQeuZaqxo2LJJS5hslbUpV7qA+UmDnEhn8Qr+VXou3
4vGr2NRDauSdVNpv06INzzDa+Zl6wpBENbEDS9nly1aexaMxkg02EGnwXyRtNVDs
7x1TdFz8bEu4ih9vHesSf/wSM3xM6c1+7uLR0XUtrzZdT4ob86HojWTxyPRLNg8B
EIQm7DTduPx/FUBA3xVkXmqua4sTJc8bExjfeORcOIiBd5MnAz7wO/hBS3eIcqoG
HHZrPMADQiwxZ2Eb1aiD+DSvlrOeMWkQ4Rs9+zH1GJnwP+DI8mvY3pnWU2E7oTGT
ATV/ThFd4QI5+Xk2Noiq056NSCPFcifLkJG7j886lh+A3Yj8G1bxUrEd9KsO9IV0
4JwKSbbLncQl2GSBqHtT2//kdBNqWVEO7xW15QvrM/SZHEQzP7qEZdY5/9ROY67q
HpRMS9oUTS0hnqb94TuE3PPAKTsb79r3Gy5o+UChpZMKFIH+UX8w7jFVcaOtxt4P
8HIdhPsdQNKq0cuwMG4RezaUGnI0Q6NPNtcl8R9Wm3WAgOsmVb1F+7BFrpyuOLad
/autWIoNzVRWalbOGwY8zq4WjMGmYynTrbRxruH7aAK+V6uSDW0naETqAEm95WWg
O6BnZyZh3Xbv4j6q0wez/AY0TfdIgk5k0HihFbOQxEOafx8dkf8LMgb7OPf9FJCa
ZmGQcwrCzoJJlwjKOPkdHPGp6ym/iKefHRg3PliSlN8RagLe45hQUD0I+2SUDSah
ERR5OinoPLXaf8KhATP8IqsRqMuJR07WLlyxxGx5yAvXXgl9a+oFRUII6JaJ0zvG
lVHXqbSkyblMhl+xhz46vdB5u1qxgPNeP5KB0SePndFeO07WCmpT8j7lJHON/Q6w
OrUF3bGff6EudOM0siJFbcQYDWEUxrBVvieUtgep7C2DR6/QdhsHOWjw9Iyqowqp
kWuqPhMpBo51VAey8cJ1uioyiBkLkiPHTL/f3GVKRxjo0j7tOie5t5oYgksryXlz
kngIucZpJoe9Sli6TjSwZLUNSMIut4e75Lp731LmXLc0OAZHxUsiHkMaI5XjkmBV
Twckidzusxd9J/Fk9wkhlVC7pjv+TyaMg8rkYGiVFu/YLiwn/VU56PYtCJ0e1OC6
CmN/1TeavMRH//hJxTjTyVXT/hWtetZr60MOSIs4PN1r02xO0XmzANChA8vlukVE
cEzH19YzYNetOBvy1K26cIrgijDKDVKKvNlzIg1XzUmktnYrOXuXbnzAeUTgu90n
QgS2YbkK17x6oR9ypACK1T9L6pneoalqON/3+gtED9Xqf+TyVBKVqArWq62469eP
rL4z5nJcQBhjgaj1WhMbBGIcq8vpqEQhrcLL19coPPQuQeMszLjQpqChG4GZPN0A
irI5+bIhIBZjLuVEk3dbxaI/ULRHdMUHtsWBsamUKKeGKyOwzwHr4+V5AUha8Qru
24EqnGneUL6A6c4Jhsj0pMtkspVoPTdg+Na82bBrHhdSytwggAnsSrvP4kZ2dVF2
66OPqcQn5ljiX63W3211gFiOEK2gBck1dPfHgxpdKGkV6ubHT0TfAFy2egRwt5A1
30dmMR/GkW+tpQrVIfX1gmLGnIf4JZagxP+zCY9pAOezH5QIsjhGtPv2po+OUhUn
CUVuKE+fpPv4F81hEywCbfGI34pWNmz3v9DqkzppUIJz/ozpPpXF4tv2YM+OFOSM
bTz/std2m51wdMXjgduCreY3W3iuLMV6Y16NuB055s61dwnnlsPsf0urmjTbsOcG
kacQO0DyQ6qeXKxMnQBzKcquiZKRqrF+/olKcO0M254bF4tzmhqUgJeGT9+ozyGU
EEXpp/PuRWEILMciVhr/L82O64Rc9N/b8pvpSnAl/JCn2fOC2KKzEbIl7cb0ft/q
OgOFkZaWmQZLqk0RXVVmnowCpwb8rU4xtgCv8C04e/hcsvYC6CPA220j3zBq7l1W
/JdguoIqQImrYcm1o5F5hoYl6GZ/SwZYZiRYjymcNMPW+7t3aix51EGZx898yMGa
awGwT7CWCkR5Lck8wGH5Lwtj484rWOgcIv9zSp3BEAu5eglDh1+QqVtNckTJpnlh
xyiQY/c2QoZJlluEr/atgFk+rIta/Xtm2ACPlXhNDS2kP71ozVfzkiRVlO9ZSFkT
y6uTCIRkpWlY9SVNMFX6bmNYY9AbBIDMF9HTVH6aFliod2p8dc+3Z0QErh6sqZ32
kpOJr3eB8gWLUF4AdE+6NL7B/5gS+fhI594d0RPP/XyqbeXPYhV7UnX3n4hw9DMK
SOUh6iejUonz9EA3H+mxsQ/WNMqlbFlFfle238cxaENlTyxXU0d05bgAmTftw4B/
JaZp3oIw3HokJEjjqnrJXh1cbcOgyh1vWORMD5IIxCEuy2ePyJVBf45ZSl3bBM43
y7j8zQTdvprlTHmviSc1AsH2NDPj3qWTPLYk/qJE2HtUtr+lsNSEC8ribZPgc8it
rSknX+CcbvgF/n86gysIxvqRVcxBdQeOmgO6n1sWLEQgv7eaXubpLB1bHWmLjWng
LpeCtnZ2q6IEBZZnWpfVaKrE/U+43Lkvd259Ph2OxweJ6RsT+TBIwGy+paJANKsd
gkA5AcYaiKvXTJlbBkvQQannflz0YfiWZWY0FfhoEz4paD42ihVCfLn0EFO+HMrg
frXDsyCS8PC+2BhXgIwJFmiBCMDKohb8gLCoueBQXmRND6cPlvz5+hb3n8LL8eHx
qXYSEEJ3rcLmHCLPENoRyqzEO0YdtfvjKaD8dqTqWYNAXTgfEcQQ5GIcAEMCTSqw
iSrw+LRACPxEF2Tn1iodOazoCg4dEeWNlryfbiX2uxUbHFLqL22wjkL1ZE+MpXAh
6GH6g3s1pNEA5ndoapAcZYsyi5F4tAo7s31TkHUi8ZP7FyOkxMxE5XVfBmK/dJh8
y6nmyZEY26h26+XtHxQYSWRIGg5e4ZxdttsVKI7NW11shbmjoLDIHCb9hVFUoXew
kB1Cq0VTn7knoMkln/8KR8ghTgx63jntnlMwVTHO1+xLk70CCQMiqliUNmdnZxpY
/WCV4wFrpoMjxoLK4S9l0dXSzH6MiQubkzMBWKs3V6sZoQzuF5QCSDYp+jPoJ49E
Fcj9Eq48nMA+c1Lf1KhPv0gmQ/bkxXRL1h3o4Eg4laDSw4wAhg/O3XlI0WtWkRa8
SNGb3zpXhJCqd764bnikuZh5ssdjAb4SWgyXufqIkDWMFKlTdM/QJdS7CSSTbC5m
j7JcS9vOMjtFWekPo+s4Tox9umCc02gzNGuXYIY9TRfPmTKKyWmD3yGy6xs0TqAt
D0APOrUB8a35+ZpSSXLs8q/PqkETvDymIE6wWOXFi0gklIxc1HJKBwwDSWeM62BH
f1XMFD3B1G8qXNddljnvW4koMOR8Ahj3UcsWlJovMo5p1sMZVLJWuLx9yNbRI+6M
JQGsgYx1EdlWDrU1MMFUV2rakVY6AgSg5fgpKO0iCmAGp/SHZueHfVddwL2VwNoi
Udbr1ENgMX6CsRVfdtaUXHmNm6wTew3M28YoKe16w1qGo3UpbpeYirJYJUJXUVgL
k3HfBXN5krWb35x+ILrhaZsQVvXMwYiNBYl2c++E+xmwvfA37Sjd9bUzeUyljnf0
h+ZhTIdANHE67uuDfCXxv9yS9YyzkirL/KxjShokegBDd1o0F8LFd8ToHt0q7KA8
Dc8eFveCszpKehk4Z+XfQhu8en8ud8AcZODcDg+wiSjDRtlb5+9fdfkze1f8CfKB
RjS0w7HBwKmaePXvvdfCaCP587HMiSYYLZdp4S3a1U0kRI3JLNbSctqoxuMBUpn0
YtM9Cwd+TOv2BXtkG5wkZeot/2t0MowO9e01mPUoiQ2pDuTmCVh6BZIs2k/Zt2KE
mQznOnLQUW4Pbs7JoIhiKTWu2BW8PMWHNt//IW1lyGbLjIes3mYpg1x5OJ5YwPWx
wZd/iWCW9JN1KBNN9u5lyqjDKHHiqZv/yg3IwS7xTa0tbeW66odZrECVaHKKLAgK
5E55kkINt9Fn1FZP0XiwsAwQu9L5QyXJaB3TRI96Y/qh6u2Zrftl0dBXju4b1odn
1B0WM5IM977lMJxH0QKixHQkxcIVCvlSY/9xmNjuuD81TXsG5oZ1tRXWyrZHVJbf
iLn2+l0ez/txfrfjSHMB64TMdcatUgwFzg7b1Icy6ZDWKAbchi7lEl1BqJcK3ilp
vZT4xQOF1hXkpQyRilmtIHBZWY121sK1RZJ056grUqjWq/356+jhchRJqO61gQ1a
koMKa6okClO+ryszAZ7FBBUMbkK6AtyJK0jj2ykh3n356K8D6y0odsm+j6dTB8S8
xHQjUZ3FsI2t4tbk3ldEJP+Q5MkyVZUJIyRABSCjPl4Tom1dCTW8FK2DP6Lf3OLR
YY6jgIhcAnDFoHe8Svz2zbXmAM3dD2qxfULTqStVdoyUfSx4t5sK6z5pjn6bSyfK
j9TA23F9rEbhoQ/THmslygthZZh0mFU8gnUzfKne19Bro+YZWbKhx5x2bdeLNs9Q
//kWkw7Xx6ejj9cOCwMT0S2qxQbGmi7pUY7qGtAMixhbBSXcTW3R1FgVIu293HeH
beVbPu2zqrYXl7Igk01vtHHllosClMhSPUYlzim+690LUJA5ucLno9nZ/d97IEv3
1Nv5/p17RlqtJfjjOqen3ux6vIv4yWkqX6fQN2dQf59GPT7S8RaypLzSfl/AuINV
zN6Dc/EEYVGDJJRod6lwmHC032rg+fcLc0cIlbqD5DKAlEAvnLm4hfqvL+gwRxTw
/jYQA9zVKSa8T8oOIXcpWna+xGmQr9MxHHKnS6qA0v7aEwma27ih9wVmuOxAu45O
+35K8jjk3OrNcIQAuxkWTgyGuYYhqfr2ctsiOYyf1vxvey7HCI3Z5vQu+MEk1+5s
rMUqvD6INwcO7M15AmNbCbugZ7igRiGV1o5dtPrTNFn5SYUXcf0A2qgJZ9J0tE8F
rUiPSBJygOPLaTARctKMM2p97rsQvaSRSDtovj47tRmuXETEoATORQIUReykuTAK
0M56ce8/RJ01erAJQEdIRIywWQVc+Ue0GEhVhaGcZY8zaMlXHbgDQCAhh69LnBzk
TNJzAwExu8RGNR9EEAIR7OaqlHweKdnJ+gZXhEmpO4w1xbzEWijdPLHezVjv3vG+
tBbtEOUt/ps7F5WR8lTVGrws5CZ2tCyZiyECcuq28YNn6LssLNPaqjsmgBhEdsCS
iWPLAR49Q+QTUvlfozKXHi460OjUiRDK2+AwFzDZM7gaWAHdwICXTa+rZ9wPTIYt
oqngitFdHJPJICZ89DdOn03k3d5FyyBQeOmEGG8ma7Izbubw3p0fdXfWEJz4CXpJ
AAwCH+3KhzJiZs5a4BmizYRXg6/vZxQQWhGCFSHGQA9VV0ytne3sKNnYMQopKGPf
n/QDXwBKEpNVd7Hp3+wuoT3LsYjyIAedNgxsw6MC3vc2aO+kit3vhfSa6a442xdB
ISVcithS3bU4c6K75itRfEqSOvtvLPpzUs63ozqVj1W3NIG0aABTn3Qb5KxoIY7y
95/IyfggRCGVpQX3vhT88qnRlFHTM5+IkgICYyIiTU3/mQAgaDlX4BIShdLhNSk0
gVckc5eZJmkFOzpIFZ4l0tRhZyYUH3IpOdhoEMk7fsc+XDUGVLg+vy682sh7qgZJ
NB6o4Wlmu++EjqzPgfKqIJxJGALVJqcClhJBGMa5DN5EmK5Mwo/dFcW+BS9Vaxy7
LEGONhsA/rXfhw2krLmch97r3kYSRuQUTb7365y9siAC6zm+3sS4YOn1V3kEprur
tIxWD3HjlWfVQBTW1cu4e62FYxSlUJEtMuI6eHd/Gp+1/yTcBFruSLzx5THCIthF
BcwudK5ectOA06isckUnM1/MMq4AcXuZia+wr7UAQbCLWHmjQatQ0lMW8VhTHDxX
oeF8OGTE4/Rt1iCw0VYCtHVdMw/7NfCur7BsfJJlIXES4vsMdT6o8usek5yvfHHm
mxunTa1xd7WpAU46eXEJbG8lKG0HvyBBQa3hvNO7wDTfFWyVzdo4eIZtBK/NHfE7
AN8jOfmjVnafVfznAOQH9fzXGhH+b6wtoGcE82SIgarewW0vyyLzTK4Yj7vJEkqH
/hyf0pUjZkE+lsgyW1UKelXHheDqvEwpIO9kx5Fp+JpBeYP1bBCIBwQE4Xhl+HAk
86uxkkBqRgMt9FQi56vqZQFz+y+1KnqHZfq07ycYwBa6EtmJcw4Ayg1btDg/s9/w
+jiFJ+a+CF1c8KxFywLjQIfuRVb1phANyjcjM0zx1XtyEpzPy9BLtkkyAaG1CfE0
cLFHXxN45lVF18JiGRzmUxTSNLBHrkhioHsgMS8NUErbPTC9mD/3D5QxDUqZSr/b
rCqEWJNdarw5+uCfldFDWJibi0nQx7N20SBrcy14Xs8JMweT7HpdnyXZ4Z5+WH8G
c8CWpdtCYKBQHz13aIOrAtF4l5AaCWLllkAF8DP649TBKMSjFlhiaNL80LligR+1
sJb+NxashuRf2v4RYVYpGtwa4pqdAj5m8Pn/xOTHDNP/41vTsMHzH6z3dGbVsDjG
LVOUiHHYdCagoBiZ2ax+W3FyIAmetdCWrYAd49UeXV6gnN094efJgELRLObBe5Ai
wxNNmVdtvLio3VPWJ09fzGW3nwgAJQLjNgftnHW0DcKxeXjT4Wb+/7CuEm3TFriH
JQLfWitzwL5UmfoYt9jzgxi8YruprM8pEM1hNyD52CEW7r7Vr8I01h0Li7SA4Y2C
p8bzkM/dX+wXqTH+hphTpwi2k0PTAAhKKvdviMlF02al+aBl73PhinzwCEiZsU4Y
zN/2f4VL9W20W17drZhz+JHdlQmw/ME12h4C9s/Kmcv57VNYJsIDoIO0Eo5epC7j
+y2W+mm5wB6/TB4x9Dsm54EyT8GIkpZDp8KoP0YOkSyUbaMSbBZxDsdC/si3Ow61
j6TBbXcirdX9WmJWyypE9qzsQoy3BWouu1k20B/A/MUf/DE1+mM6flW7qk1CV2hc
PcUtBiws43Mdwu7Qd94cTMOceNWv3gMvkJ2fmTp8dqHg4Xj1CgFdnfqUy7D0IsYF
w24XYnmr0Ffd6zDupJX1aPMvYdVT8vpVEg36mIYcfuBf9PjvcS277WXouxZo4aMW
ccXZeTwMPoJjURpvIpP0SfMBM+oJLllmRlX/9Wo06NVYtz9U1Y1y8mtJ0y+BHdzs
q2Tt50VjQ9QWDhE7T1HT9GVMWiQhc+X3lJmK7Twtc0X8o6ERyk0V4Mo1z9b9C5bf
xUkW9ZRThsbMkaNEgDBG1BG2XORDzlsj2TxP6Z6P01yO5jYbII8ux4hbbNtsU3iv
PgoOXofZFMgvNffo/JZaxII+JIyHUoTa/tjM/DhjkfX2JGyY1QZGZFSWL5ukpWmH
qQXyf1QZICf5tIkv/pI1tdrsRWnau6cp5QO4QxRfjnW5mD7w70zs2wawv4x3NiFd
22x+mjHbWd6m5NgpkBs91N7hXvmWWzj+2QO+D+j1W+1cSVyuzpy7yGCBhucVbFep
TzLLmFgUOW1wZBtu072NUrZhnjxsaIiu6B/wjUPTdmD0Oml3Z7LqvkVE4WDRcc0W
6Rjxy6hesBtfoYMJaf4XZIW1U8otgYb4xIrR78VAKm8ZAzjKlJQJGyXUflUPgV43
sTq8HK0F9la7Z2SPZNxodqJVEwBwhupepKSc4JUJJ5ue9I/iLMMnJLIjsNQQpNeJ
eoJJWy6m7iRwVDDNwZOdlEbuBqEhG3Mm/d78URG84zCKOCB369kQUItNTa68OnRY
IqN4aiTHMOlaVP4NLN75SAZb3eEelY5We0m1v99w0q821ezCuMD1bs16zrUf7yNy
RVb4yvBARIL78YXxfW71JCivt606AZ6Tr+vA+fMb11NCEg0ZnkcvdRFGLX0M4t7e
LWhIcl8n2Vjhoz362lHpkgWXvp2iIDdfBCAc05O4Aa+jCoz250ys88vmhrvk8Jv/
B0GE95UpgQruPrusgNkiur+Gm0ZMEJSyeOic0JSh7UIAvL5G8vCZuKSDU3al1Gqe
GbhStLbtt4tDp4w9slLeqg1i08voNx1V590WRcEP7C3pa0e1YeHQjgMnJLtz26XC
R8DEkYWMqWESx5k0z4zYpBfH11lZyCV1YcxEiprS4nO5G3N+P7CDTJOvY9tREP7+
RblImU/lB8dHh5FfdpZlSZfZ0fLnZobSHJ+8j+3XfEy+/CWQS9+eOYU5C9fK1f79
H/BPZmXuxIENBoUTJyM7G+ntZ70Fm5iSph6BGsJfk6vxtvT8fni/LqJaEo//vXeU
HzeaZLb3Pg2LfQ7Khj2m62fRGLLwinp22bGFzptF+iVCv3iGjMQAa3GzYwM76zXV
XlbqtdJ6E0yHumhM+boLsw3pUEQfst9XdQxewnERobCqN1I3iM2u5LZ2u58e+y0n
DZuV1yxd1OyiUAFRKwtsDZrmGjfZGnieBXN79zyl8tzQXK8eoc/tGBtlrIHDl7JM
DXDXy/6ffKykVvhxWhexI3tGF83NTEeLFHBlyptHF+Cb/52K6BUQWVn14RSiXps5
DW4sz/dUOtc+C73wh8wprHEahLCBfONy2IL6zx+3MmSCg9LPt0lgvOdqa2eShRL4
fH9lzJAYrg0l9YZQJc/Byz/X7EarMtEHaE38qygpQS5mCv3ux3b0fToo1AuuPZXs
SByknaJ7KpUuKNlPzi8K0dypNSRKCN1xEHUOGff0PhiSCAlQcOUOzdL4z88PjHrh
tJeJfzatwudhvp22mEJo7ArHnfFfcS/T3zO1MUFz+S8FOvtpnvKkxsPSOWyqZ8vw
cP1XND3orqH5zumL2kdUGFE+iPUytYuI6wLlYw2WudiCKUzYdRSDVfbbQbdVXIzB
z9akRdcl9SPxAMSp3qgUcm+WFuZf4sCLfW5lEBFkALHQoYx08q42ORoOfFcagCDH
pALjuAZtrO5ql8zaYWezfKt//fRI8QcgADU7Xd7j80jinDoFdcZS5h9/D4CrJvlk
PM8fjy69cvKgxGDBc9J7H14OjR8AKuLr2VusE+yAc+DqdsyRsnLDLJz4/CxhUpui
Wk8AEMdgvUog5RDFt7WqnC53iNp7Q8LFWEvi6U0UgO04vOcIUSbWqSDYh3wVBo/w
aHOmcLgMi7lpJ5EzffpJe2Aa4B4E+mzWhJf2J/KBnFSpEdhkiz5cg5PxMw4xO1uz
akXBUvwoRRro6qroxNLwfVGSCtHh8mnWlbqRSy7JaDiWPn7hI5fFqL0+4nAaco9g
S8+PcHSJchpZUzJdLLnlcvji4j3VKYNNe06Mzz0bEyMrd5Q6CXVGLk+eE3YXGdQI
0DwUBE1Bi4XHWplZTZdlzuANFDssef5UUd0imfzTOUvUAn+ZIDKrS19Hzskpn5nZ
9C3r9Dv3S/FAEiqmUyFM0Y0vEPwgOrSpWoxjKZ2ODuKeYPr5GDK3TCDEanK0T5kY
/aDa4FQ0RAF8WIqAzNWI4U72LypzeNjKg7Vjuwh6Ip4T6AVSOkbG6x4QfgaFrec4
d6w3ukyuaVZecKmnBaaVQTUg5SDP715JL0b2IXSsxufqlebslGAyQ/qo0vSV7DUo
9tvDrlJM8gj7TyCORc0bdSkmU/IZ84Z+P2piVWFFejv3o955O8SXeNeGuZ3HLqg5
3Ga2i+s1zCZGheFMWU2Fk5hc/8idusoPX4kG8Yu6HicRf67/Q8TSEvPrnajJwDX6
alX2G41fT+R08rvlQ6q1f7XE8hgrVqeXMUg/Sih35XbyQVoLJHySd8FVUdLrNyV0
PosmqDXmOo4v4hfmg/pW8AR0iPBRUOm7BqntP11PwyVQTYnCRJ7J3huIovHZp/bf
22fT2m8aoOhY1+PI8+aRSPIJRkEQQ7KMR9FehzBWu7m9SUIoxKXUrU0h2xveC0XZ
sSvGJT85UrDy4St6bZFnxmLLwlsecI9v4QHwmvf1I3aXtZzQXPKtO+grdZ1Fjgz7
Ty89wFWS3Jic2AjIrPs/43xKou2Q4vUqjD9BmTGTn0tqDpprCqY5gflusBCbwGrn
56ZvAiOYqhJJLNLtfKLNFfYQ41X1F0DR7WB6FHppnroYp7jwkZ9EWyEetrToykq8
ixK+mL4E18pf0Kxg64aCaEMMUCePVnpMu7HKFK6gctm5NIZmc3qln+jEjGqrBRuv
G7AxldSZ5yREbjd9sg0kym4ue1oQLyDZwIFEfbqhpq9D5U9/+ZJvugD7lR65pSaE
w/yxFqZwBiVJ+WYObOXEy6Xcw/+VTWUH2wvVFpq3n+Yqnajcnd78/+xgYoyeJoN2
ANFoyDaCs9jyx81Mnd2DUFnfeUuH8TasEgE2+p4yJjdNyfP3W2EzziGAv2iXWcTK
tzRpvWXO69Hr3AER32gacxErUANPhprsJ/ISYEgrLUS2JzTPVD7PVUodsYkXsBHq
OdFVtd0RhjMXbY50ymdSGWuAwJQLmloflNnMm7SXq8LKgmQQqc0lnRvN2cOq+GrI
hsg3YSpmc5tGV3uvlSTjWSOTTfrNInfW/grFM5J6v5I0HRvoIcjgRhJ5sc9+KqiA
mrGaED2GDsmeBZGRulI7r5B0bcwjCgCGYJUeDQNIIHFxsqGXUK+NhoAq/RMVIQsB
d0h8JOgKGMb/8rEe/79rnZAcuNchHF2ZEEPskOGPXUu2Gt83JkxkYDwyQvsQ0YKC
VWeS5/2CfB9Ss4BN0PngYFsRpHpBvwMojnz5OSgofWHfnCrQLFgYfV8I7wZYtX9i
wkVuXGJH6rpkPXqf75y5kIk8tvPIgntiI6LfR1yLXUZE031BxQVxpQE44aZ7x/49
8GVmLl7LfWV8xoqfLSPVxE20ydSWribiPWPw2MKm6ID7KnwRGxuWAnVjMnUUyrsP
gNThnDBoF5I2IQT0geK9Ep2dmnhmNWKHtq7WiUL+7cmqXMUxwaY72IWgw0QpkHgA
8jQ5AUfB6j8v1Sf0ik/dJmrPPrZpEvTrBlh0t1LtWutivxbRgUZCOh8vJHR7bYXW
dN0DDVRkbvi7c5z+X1GNqsHuI2SJ1z0ml7ZCiRF8ati27y+YWkFAYumgl1eZRkkO
J3k984engBv3uPZyNfVwNtAaKroQWeERBfgsPNTDJNwqIFQOXbDujdkSCBIw+Cbm
/1zNiAFEVBlXDH8UnzOv5TLroTgwooVV3XVmdORDuBCQk7JqTFV8ZrF65R+MoXaK
k4AGMVGWRwC7pp6Vp4z/xQRQ6HXkwCWbdgr4Z9Ja+NJ91NNAr9YRAsFEb272yNg5
/ZlmNIDN60/G1vwFrE632YK0B4MKpUScvoGA6GVDjQeQOayFCYbK9Po98EoNtw03
oTdbfdZONBOFlNVgehz1her0JgQnKYyYxfSUP5WmM4G1BlYju23i3PZGku6lpDO5
YjzpB0f5OibaybTbaF3qMh4TOmQ/pEnOGZWenPO5xNHYSbgCEIMcSEpvQPdA/s0L
RnpIvZ2NSTHD7tSTIc+dhrnRjBl5A5xNABagmYIjUi2a/I10SN5Yth5DM6j/moJs
1nXXLt5XeHn/IqCOnC+ffkfwVHEyggUOIFpErQjpR/DojtnDwgWoWnW9tt1gkJap
I/Gp87c7O5VE+FiuGDW8/NaUDeXFNo8/clIkhtIZSPHP5yUDkZaCMx20EVqZgdh9
9r3jif6PAK86dbe9S3b4NX8E/78ml+Qnrin+Qo2GLk9ZfProXXILiQ3TlCYavUYh
vljC2YHz6QL8gBAHt03fOdIvxSSp8HBsCWeLlV6dj3TfSAEiGf9vfD7UeocPwI7r
uCiG04QVdMqDolTA+UaCwGFs5nOT54scx9+f09lLhk+Moa4Xt2n+c/d+FZkc/b2G
WIgzkTPPVEveMdCdp6oB+Yn8bwHMNymNnolvzTnO7yCcWYKMiL+jaA9kZ688eQT1
K4V0xCyIdiTl6L1FImDbL/0znOfX8D+0m5RZXiAZYHzvbgc/O9HVxYOYjhwFDgEX
0dNBE3pTvGpFrNnvVZ0BidznyN856ahByTD2S0hTh4M7v2Vy5j+8cj8XYprLwaMP
p3WF/WLofDgXVfS3r2Rbjj8EyDqY9662E7oIJQ6sGW5FAxUDcjYzA4d7rEba82rk
+jmLmGnogCiDLz/GFeT0rvW9hVy4kJ8ZUvJ9F0KQk5q0RotCrcos54Yyid0zw8js
xf9nSOgmJBjXaww1Uz4MCfSckNK/FeWJQcFKjSkRfj0y0663jK049Vu66L9nyoPB
hSlQphsZTlTyWa4n04k586/uwyHP6hvSN3qozLi8hoGnAxjE9j+GPNmKF5TDw+4w
/Z+nh/ZLNxc99Sw56p9kCCsmvoWHCHN/9WA7h+CdNINVUvuKdpEnlTPWuqUI3Q8J
F17XMIBmeZxjxd/WyAoWpHu4vUAJXmcF1Z5paOQJptZDk3TDe9CqZR+4THD9wCNO
cdy+mbwQNayrs7dJhLuAB2HMcRRcoEu2iDYee+y7UIn2MZ0P3G1yjk/+btfrw7KS
XKkcdl3exCvpBjqkzHMQVrsz8YsE0bKzuE0Gtjr3dGUWF40se+uTJ7uhgcP2o+Bc
9X1di4AXonNsgTCdZZIkEMR8cPnoHDTLkm3zYMxAxijognS9PZgaAmR3k2QL4Pnj
7s6l5ku/ZPOisPXMaE3t0AfZDePgKGoDtgkfFlDFA9KwU6PREzTMxf5ZeyeWjfdB
tHl7iBsXiOAp1eMiJ7zwcUDM1FuIUGdzqDtbjtcGScFcTmT7RRg1WjPPgPDoUOvO
Jv2/XwNuVI1NB8qI1Q08SgF3Gn2PMv+/NbHeJeLl8VqVPUP0U0RtrXiCtJ43JTtv
RJbewAnFyRK1Qrzj+iGnrxcy7NC/o1aVcwGdHIyEcuRtyRbuSrOZCXTgk1OLwbC9
QACDmbRJxcfQ+dDKA14jrRfZwIPEd34SgT0l4YeDqPwOtTukGBSCz1S4Vhge2xZn
u6pnNP5xPaTPGIdaws39eIPfQbc6QQzShfqo5LrOA8bVR1KnxRjY/QIe3nru3ODp
rchCuXocCdgqOplrBPPf27RNrs4WVN2rlWvtYRtWuG4W8ZI++wE1L7cn36cqmCjR
C64KNbp3xYjPCoYmFuD7c05UNC4eVa8zhNDp6KglLQRjwMpWhZ/L5DEqq8HNQool
i//fsqI62gISH6z2PKCz/BlvtFE+6SrG1tKitlFZeDa0zbFheKv6kB1aB/FfAnOU
9F86HTTtSKDhyfDlicfVYJj5IVR+V+s/HQebkJ7XxrkmKe9KrKowOfmV/lA93ycv
VTr0WuGA+8d3efCM3U/E/M2kkeRg5u37UeOYWRKV4WO9UisJf4XqW4y7vDm7jhZv
GfTFBR/BvCnBqvqrdLnuCLm+BstItWRf7g5k5Y8hZ72ywnKxKcmqkjqUk81XvEdo
7jbiJXVaytGtlXySxB6MR0+D+haKTF7ZkKMhKb8zSmbSOXaq8xJBHUOaJ6omcYJD
768N7NIx4O4eYitxCuc3e8x50nPlztu40PKk6KLBz5A05ElGz9w+D8PFxio4/pqz
N+MNjCDoU1z5Oo9Nf4aj3Zq+stulKtjAxDReauOa+VNGG5KqijIVlFiEXlhIKgQE
PS3Aj9ONhkFZGinbiylUzZ6kPs4kNatA47pdovvTLlJewYLSx8fxEy+A2Tk3Z80d
6zEvSO5EL0SSxBPLe4PUbd7SST2BTeMu4uz+4IM5zFlkS2PGXlAKvOv/de883A5S
s/GB235BGwSYNQRLZ1cKM+QdBSIOIJT6rXBQ/CgSP3KVKPo5mtOx3KdfP+ifdGgR
mdDRUhlSfbyIt1SwiTpPumMgmNaPtjF/DRMPshzz7Eoe4NeR0IJoE0lNoEqAbx7f
G5ebLI/WKqi6y5TEefDY67bCIU0FCLL7rj5Z5FJVl+RBoVmyRXAKmdgvKsdGYJk5
eqJ/+fA6XHlAURtHKW1/oNZnL8R4lPNxPk/xZ387ERKvNB6eA/jawv+xyElYIBRe
G8rMBH1An2vHUK9Cy1pMsnaAFuDk4o2zUga6JYkUPh2E2cYhmSy3xcXRd9RGwnar
8HoxUVsoTvEPq4OJBMMQwXYPbHCQHVJTLKLErhiaru/9CfluZiNCcfhC+NGfv91Q
yB1CcdYyBxa7meQlL6YBsyidgaR+YLKfrg16ZemwRhCcr54F0Huo9SCm/0Vq5DoK
B2la6E7sYZzVK9DqDcw5Ej9P+ZvN5kD57/dF60Hp+jZ6ASxKilHtJI63Jvex0u09
lolwnch0nBQIawsZzH5rylyx/7IdBc9qmvAmcjJ/RWiulofRhgvhiXzrM+ryc+y7
TYURlg/hrsyrI3UWPcDQOHZaPHb/7064azAYRPnTbhH95MJAxpadESIApvICdQq5
vx6JZMWJPOFdEA+qKGVEocS74U/qj/mKpWuwoOrPA4psmoB2sMo6l/lQC5leFXIV
5vr5bgrQCK2csl0dzh1K21yfoR6r9jlK70oPh4Qw92S+mYDb3bhx3rjfgGxhQVoL
3M88NJEX1VTmgP40tW478KPgTvvm8zn/JMfXY2BmjnBN64n0XTHA++YLi8nXNhvj
cDFX74xN1t2Hl2AsmATa7WSLemESc0spAmede7DYbVLPWmpcF2/khUKL8N5TvRvq
YSOgp+Unn3fKVzNRSP2z2F9Kg06Ag5KZngJksUcm/fvUtZucZMdtpaYdu0NGO9D8
AsQ7iyt8SsRfi8auARE4FoCwh5S0FYGWAeCZxn2NlM5/OyvJ50T26RjwDO9eiiq9
9kohsjqZuK2yKj3lby+Ljq364sVWMRv/pTB8nhlL7a/pnweChJROgViz9gtmBRtW
CaN9AxxM+8STsUuKcSAJ/ZQbuYyl72TKia+rnENWWXIDCwPTzwNfL9zxN6FUu6wE
hiA9MiWIhyP6o7otg9f1llcyLLo9Ky3v5xVmqAjyn20QL6M9dmQNe2iIvW2G8gfW
NpBK03PmJdvxozDQf7eews4192fy3L4VNabl6cqj7lod0HXYYjFTbFZtDH+c1Ak1
1PhN7cDHOfit9lRKm9wjwTkoLZlj++36ZhXrk4sgacqe5AshBZAIcLdUzQQfHdgU
Rd29jnADf60iiUU3fuuwyrxpmu/Uw//jhlzJUWRZsboNwvC4EWo8Vexw7wz/Wlt9
uWEmcyIfMg7bXKEJ/qvbzvrN7Guya50iXXDFB30thMADlFYi7pxVyISdrrdbEKvi
PRF+PtxxQmQdu0mj7KPGPy2+xnq8qhMa1on5x3zTN0RyvoHeWUzy3/da293ZMW7n
IzjdimVlwVszNtQtM9Tj/WStSCE/41+MsIHnEuqFOf9RVjdiDCVi4YCavXCVC6JT
+CnocabsPMyGc5jpkwn66Ouaf441l0JfghBGCRHbk8Fz0dB7oqHNTwReY660UAON
g7P17AsDfZyEkwRriFjn8GLFZ6wp/NpZ6d+zRrh+OeUo/9MOARgB0obBdqlzcrqu
UuqF9NxyLjwCFT1Q0bD7KfJxLGxZZCycVC7EEW1bgXHOY/g7l7OkaRB1aDwISmb9
8Y1AZx9tx2P7UGQROam/9jIxuCJxMvF2Urz1kY375CXjR+R+5D2CRKLS0ul6bSK3
Vh0/+lEKyoIraG13uPlDECrwgJO9Wkp0QMjUljnJbPYYmOq5IK0pkQjvikJFNcAC
YflZ/lqobmQlwuRZp6iKdxexGs02O8tEANvxDwx5pGpsCX3guhALhYmseAhqxN4x
VuzaDZnwiayFqzo4yaevOkQeYO3abjw05RokYWtoK+x6yBZ9OihT92VmLZ4MbmqA
ur3HS8kPwGek5sZsiLtisZpgr6/Od2SbMfogTlIqMNQT2T1MyxMpyS1cvpT9hSuz
Mn1Ih6MN4GJJ/XZ4uwVGw8rsIqHrZujZ+0kHIu7g9Co3Wb3fWR/XGgSzi6SfKS/D
f98QB1JdZHVqEcOIIB0rQaTtF6nUTvcw41FZHkMMDv+nafO/ug4pDGtmeSUtCL2a
FKp7XfYD7ht+Umr5DU3jtlqKLd6ycz9CwIwy83izhX1pqMxwW15G6uR6pe9xdr6p
3murtANLmbMBEBc/4Wjj7ID4b34cPRURTsv9L/NB3zas7xgBM3cgymEdAtbURnll
AqFoJfpMd4WbTT8I4ogGZHzXRmahkmBwmgBBS6P5rz+2efX/+Ogdpsj1ZSTibo7f
cLEmgR402EdCsaQlpu8Aint6j01YIR/LO2Sg/FmDtCRYdX+s06gRVRjU9LG1gE/x
joYDhcUuaBAqcmUkndBN+zfekBWtp4gxgx3aZM/fCBwZYUUMDHGLaLVUjb9k0oeX
gj4QkOIGYkQUh8I2J8iGdjulLGYXcED1pviN1USRfIt0cZz2kUs+pkApOXIt2fan
ID63zeOLJ4dz0MXvPXsFFljrQQyTVTWperVxPHp3PXidgMosaBPyaGInfsyFKyvX
GiK392MxFDs8xBxe5bDf2IA+t3zQZ2VZiBCdj5cfY4y5qz0OLS98St1rs/ewauKb
kZtytrM55YH9sF5rmLJbgElXSaZFkax+lo67YfpXoVhskxcdo6I7HKoXsK3D6Oan
RS1x9vzbiM6ENSBQTf0h6kwaxce6az/HXuPobSEd2VRBjBEWSwdVE+a8ozSgDA9a
Lyr9SgmaOvGZPz3mGtHNGpjUIxHzE5kdW7G+SyBRj5vFAiMbrQb8R/+w6hMhPIL9
4wwaRRm2S8ixCmN07VT1Ea217kZ+oD2y/nBZhggLbwAopEoMYLOU8rzaR1FGOoyi
C/yPL3TPCbow3TuoRyMuGoaUkR4E4O955UK2HIDZMpy03m6mIgRrbRu6fE04V7O9
Ic3QROAV71WHvSGcOkLMOTT5IkOKtWiM56EqsJdNgJYtujxMKJpLU14c3pRuKS04
XqEf8iX81O6jceSF8mv8gCaShGiZifAx9pGaMhHu7ukO09sjmsYucL51IvUozXwY
mCBgXgrZfwa0Y6FJ4JSUYwwosasjGAQtL9yc6x3HqIQ4La8pZsmGXm55PkgcciCl
gTP8KX1QewDJ4ut8PM4CLY+4mGxAWo6xq0Za33MfKSQ7kbKbay6KDNg3G34p6zRg
5NbbTMLJdNEL3wqNVngKcmqx/+ppc2zjCZGeH1UUf6bdDXckf66Pu01wNvbY9zw4
tHHzKQ43V9sxSWxTYZG2QNPVjXOdLBEfa+ozVzaY/Fzzjs6GUdW+R4ZibuzxGEwT
NZXmNYgKUj6Hh33cJzEGUoSkVIV7b3zU280C5QWY4O8q5JU9htrSWkTOUOMXzJ2q
aU3eMCViWE47CapOOTALawULN+Mip9/zzoHn2U0BlAh03I3r9pAHouCEIoQMBNFU
wLtatBK6VuvYu0k/icgwjVXt+tmP8tzm/03P++RoCFTPTBJwCSP6Q7ngDMvHcD1N
2DYBFeHk+qISXxJAKnCHOVWgVm8eIgvkXT3mmfzLZ+aOhsLzla4O5CATy4sOwYDY
XkH4Pb2WoehzryadMe23/nW4duQc/46vu6puxfJS6dTvyKMCVP5FEX50PmmL2Y3w
lKxOpuMc8JoNi6v5/rWlomOaxmkvFqlZPHZVc+RPJEZxetuXA6KrEOt2Zjskdi0Z
fYdbvj9yXdu03r8+ydL0/RwM/ox/NxTXMuZkF3CD/Cn1zA8q57WIuPeXsFvatrll
qj189oS9oS75iI/FzTmK1WeozFHcK3srGwtriize+dOMEu79zMYwZg+qbWZQF+IP
whk8FmtZYp1xC6Or/3sh5Dpe+zyizdWF3ZYMOj7tY9vqL2ZHVO7FIaRcXKX5oLvN
dQDDU/+tKyTHSXLeFKUFnZKkhBVg4hIvi0T8nRlmoFMwE9n6Csuc17CFhp0Q2S+5
ucHxxA9W0QgeKLM7CvyKkpU3Yoqx0HMrwtIG8XqF7B94bUtAl5xlnR4Xx0Pe4NI6
Kfqo5UfRJ2ZjMOf3qTGVOxF7HfgEx5wUcqKyGZrw4aZ3qw0VYwDgbjkcgrjMPdRP
7+88zFLM7Ba26ChVzXxWFFadzAJbHoRsRWv+snS//Jb8iC26prUnCor/CgxEqL+X
+fpvhIFDohfVZFVwN4rklkiElIGoD/+1c0UtE4gazkeYnmLnIoHFlfkZzW7IqgAJ
vb7x53lqrE2JwjnUMBj3fmMi4YCZbrqLXovoWhsVnGEmv+UO0TPzYMLl+KGp8bAQ
+QyZNZLPOeVy84Czgeq7lyRF96YXX5E8wr5cy/Xeqjhb+kFTeLm2feEGo/HB2xhr
hEhrcPnw3kay1/WN9WT/j+Rd5Qzt3q+E25twjzsC7JSdt3bWj9Z6LJh7z+2XGTu/
hg4nhdG/Zw4At+KOW6jpm6ZZSosF0GRj1U/qPIeGc03uC8saCz/6/vFVD6C9tSqi
BGMKhUf5VKfYd3DSPI8VAhNT/xbV4nnw305iHHRnqq84oBV96UNBpBCiO0LSOuch
s03YlP5uCjURfx6XkX2xPY/Llfi8G28wjrJdsV9+5VNOEEqNii+wLCb3rS5HWRR7
8hLhe6SPCttWbWjcdu9OT9oHL5hkjhFqpStk8XPTI6JaaSPa3axlPc3l6d9g0P85
CW6Wz2hdbNkTvCh8Jg6a7/BTsxQt2d0SBRtXNYz9dbN62DKxcioxLHw3PDmD+N6W
HBZvSpDWUuWPhZnIdaQkP1VdJ/d0vw6PmXIeUK9cxXSgclUTB5SCTNA6Vqj53gvR
njgYEa6pnH9+D3MQlya04A5Fq7LGf/n7WaDMshkQHbyzVzBPjpOwFLK/TrZFsVLZ
VgTG7kimbH1IpEjwlludlYC2GP1R8sPgs25QqqUYuZcC6jvFaqBM4wntVIM7FCPK
S0fb6qDkN9yGrGz42LT+ujwI7q5BxdxeonipdiIxqUqZYeImHtxPZMda2RCZ7mdc
jeDVi2AQNkLQnsoxZGN10AwoVa2Bc5Y1ya+D2zSHMxBbatN0xJWVlQyX8SeyPwx3
37IKCrCPS20bDFjPTMEhTbysfYhRjVwM7DwTUF0I8xwrQzPZVcKM9ui5DQmDX/l3
Rrv1NA1cH50sBDpy0aOiuEyfkCSIbe+AO7KnKxAa6sJ0CwCO0sy372zdgusfXU5p
xKdxAlnqnSEbmwm+/jtBza0dI4Oyw/z5I8lRivG7nn9VUIha4XY2clv0/aFQ9SRz
iAZdtZ5nTze6YDgZmcUWEBqRk/g1vT6E7VRb+B3LOVSfEWE2WcdwiOPN85NVSq5i
32Xyvo56IgUuusTUZ/szcOFnPa6BuRDsqULj+Gv4HW6RZhvZYDf/48NvYk1jfy6d
dMIuIAI+DCmEiMMLtzK4luXxtx6XM9A5yAtsWdr4vIDtAPBx08MupN/Jftx/XikT
u+0eXmpZA6nzhcUDdLRgFvS5VWXF7N2z48qvdmoeuMnLFEtNg/1iK6SKZpLqO431
erCb/1Sil+59TXgTR6h+PA5wwYrTVL7Azw72VWb6reSndt64bTmARnSLspzGIVjp
4raDJ0hOGZziblN44Dg/8FxCHgyMuwsWgYJ662AK5wLlUxRrzIbvEgopIAczVkat
13RcMSr0B0T7oUFq31B3HP5pOTVdwl9lT3n01PvXI5FFwwKod/8xLE3/u9v6X/cJ
A0kXLH5scRYUsTT5kjEJWI58W9zFMGj31c1EnA9Y4TtUtcVNnrgwHr9iwxGmrozK
6snXzykANyZNpWsZUM+vJRpP22p97ONnNX3tQLLEcH7kIbsCKU5xdVGqN8LwdBf1
se0c3t0M4yv+37cE4DvTUCLAyk4vlmu86mB5CrsBQjrX2+YgOWjSpAiEvbP08Wrj
kW1/n2CqVWyDcWl6xSxQ9mMv6V2nzKsa1O7N+8/ukLIQ/iGemNcZVPjdw6tNKTW+
yQGao6FKVUTBf8DwuWZZf9czC+zuoUdPXxif0UwbxUtR/bmcUD6Uev9E7nfAYHz+
cmO6Tw1ObXQPysR17Qedb51W74ZYLWUupB3PglpDFFZRhSQiJ0gbI/q6MY44mmWV
49jod5ntw4Txvsrt66Fb8JTG7uF+IUPxkNQ+NS8WshVUcvORdN81ZuEOklDAYdCi
YM0y0LpM6G193WWKJE4eDOYCkFwXIIKiHzBOWKnONBaB7lY4ZLiir3EdY05IBI7R
vgTXwEBY0OdztjuQ6ZQb9CsyhaN87OT9N0i1NoKIT0Js+Dd1lwTSAwE/LhBfuPap
njLk5v6TyxqTp0+aBe0+Kb1LTFBSgnFyUXnpGtJXi2dRi7CeQs2jeO/wh4jyiuoZ
TrTf6HEgTy0Vj7ur04FDfA/7CCLD0zHOVabEyLrJC5XazvKSUsE9gEDYtJsqeZFy
AflbrnsX2hbiEeyVQjYol6GzOzrjFMTbp/tYYgQ4l68MYtknilIpcttzlXhRTeUu
b9Z8cJ9NVae1WnRNwRRviVz+3k1lU8d69s2r2NMOaC05VtNaYgnq617TSPIJZ3Ju
ugEjOGVLt/XvVp5H1NhFRgtZBAmlW79sO0TcfK4+Nwlka4k0Gj0/DNjUOXdtLXWd
sBM/C1x/5DIKqd1f+1o3yLtpVFqQAxbUDkyhGT5SjZNSb/KrbJ3rA36GsLrslm06
EJwB/A7PIe1Ij0J+xuopzG7jZqf5Lae9dARpjNOGNxMyvH4hmRbSSrA5bOcBRt0n
cVzG8WuFQVH0vvSoPCA6ngRSqIzbW6iF54O3bp8UGhiWKU9yVrC9wIKpmts8nMtg
AL4L+4Yq8O/1EtSsrGvLi1F78EnbBEmyPPMwQTH5J6fkAdUS5kg07LEbRha82r3f
1nvl0xRYOT4SyTD7uecsH+Xra8XwulzyPgCvwGOeCWmBeMGAiOwo/Ebi24Iz1rYI
AYW3WLASKLMFnJtNtmZgU9YhdO6XLYLrLYZ219Z5Og8uD8LQ6yUepd+VsF8voLgA
4SW2hb7PHU6btkL3nlau865V78IF0eG5wwXS9WLKDls4RhNvXE4ydh2o5T2zVagL
EGv5sr5qbydDT7owej9BV38EfGehLFT0i/IRyY1JkO9yA3gzCcKPqRofzZipWTGt
eSqogjTU6dIj33dnmoOTs+dFn4k5He2U7BVhiOOxUl7aakHoOhJKWqnn6ZS625R6
HJcfM621bLEsThCbiVWeXVpmrowEbr/g1NW6KVSbi4RuTMjwbl1VxZj7EmKbxX0v
+lj0qRttcSAs82jk4VLkGmJnPPeGNQAFTG4OenEEEpS//IYj0z42ga3ezsdoh8gB
oOS0+Hlb/6CrxzuK299GMZ6pA49EjDqOtfq24ZHk56rUbVEun9V50rIecNvUESRw
ZOyudgAyN/NaQkAptPb2pBddVhrS7F9QcaP1E7z+1q3ZnTEaqPPex5vFdzly3ldT
5e/Vu6oL1GaCjhbdSqjA/9a7ypr7MDaxXsyy4A5dN/lQl5bK872L+gcO6U340Sdf
XEb34EXrPpjvnJDXVjMSyO6IMz+pOSTChxLJp7uT/jXzI/I0g1ACrxBCVwgp9rBQ
lIxRTntsJ98S50ULAP8mm5Qep4598iuB1cNphAnPkIzSbjNR3oQpgAAqeGYcOC34
Oy+Ud+kqcCKMxDdHeU+39Iei1JjevCtWGNDCOazAclFAJfqtRIt0LpV0rJYMQUij
DogF9poZan2N7kINAquCQ8H/CAZBVpZfFunBFUAvN4vbcIlV2XkrfKWpn0QpS2QG
Xv4P5m1JUScX3NEVsdMRyhKNPTICe2gnpYxCXzIwV7fWGrCLbOe4CriTKMQ1VdVp
BK9p9ZDCIFvLuFhuIq6QMr2s1bq8rwAQsXSxHol2d+lkm6qFgGAwT8DxPoVe1b1V
mTqYlPurL1xK6x3Ew17g9En93GYj/J0WdNDz1the/lsXy3O2W7ESvTAmgj+LFeMn
lBcoj+I3z40jawZibbsAQ4z24GU0/0Uv/9YlfmIKEpLqr9Ri77mI3kUhZwgHnbGN
+n3L+E4oUzmTDFrpdtmiRq/ZAhnwEHCEQHeyT/aSxnoxUcsoCmkoaYlJJjWVu6je
WwTzslgXvFA0WHiOE14zqi25tYpTp/AkVvD9S9sYyYFHy1K2gX/zxgnS0CBZnyGT
4vvA6fB2/4P8r92bpS1TP8L6dPxPejmCGNtQwBZtvpP8MLPltc5P4nm7AzcYbB5i
6wWMcxiQojvaeQXpDNWSLiqCJaYNBh9opsQ18Bawnr57pT7+pLuwtMoMHDL2GnZe
76z3snJD6zwlribjF7LVNxEOMVjoT52R01iGtJ++4bID7NMXPRqo7S4EsYh1lM0o
aRxWcFOQpIiWXFLhgLX61M3rEoWVj2MFfGX7Z5DF1GXboJ1HaD5pX5Us9fIJMOzu
Pm4g14Uq3QiyE6BQyqFssluLlSVPSGImQe1553X8+guqKgjRHm8nrmvHDCgNZAcM
kYp9yi0+T+j5XRjZcQpR3CkCqtbOKOIuXsQ0qmrdZZh1bnv62WvPgwrynNmJ8yc2
usnMhcis26bLb87fkw/wDnM/6i9HhvtmgVYdK+VXgvHazFiBuZcFsGhId0BzjRPV
xLs9IOCJtay7xQjBe9yUrDP7T+WSvCDCkjBptkQNxUpC3++swGWoPmG3xkHT4pOX
BkfqE0PHwJhaJ4jLNDy+4W2Id64n6mzTrZ6HRsNnehAUEFLbQZ+ASqu7QcYJ/mPp
4FNPiL1A+IueJE2k4jNn99sUuwpOv70VHdTSsJzxo0dQwWOY/VDqSaiN6eKJfcf7
+YbEc6xoTMgbynMEL60DTFGtIOUF6JrEYQIisAGTazOiyOpTFw5CgMV3oIfDjgH6
1qP1AvPOxaZrW4ICoynCKK4rpzDTRsR8TrIUyrjEN8FrnDp67J4AyPpLWWWWqZj/
xBXFVEFlFesXepQWBW7IU1gRT+Wu63F3lj9xt1Rb5gmFtqztOUyiwscH/bv72ZSq
Mrrbngv1tSthgamU4l2ieyzldjkxQApHy13Zcetun6d2Zp+JP6XB0MUX3+osoo2z
W8qnJr4TsUqukj7e0/OeLDSXcOmipj5KorKsy+f4lxRGpimfCuSjODKr/DfmS3RG
Dv6I7IGFjEYuu1l5TCr+CwiDpMblHSSKOxAMDUlBx/F8jVAgMgF671HEQ8B18c9B
332hepqo4TuyYNLCAuRFgS6Y8J3Xa4N3nq8LW5LTM7uu/H/HZhoSqTxp67QH3uZK
CElm8iY1F7vXsXDG2vv6rAYg49xVyxiDySNCp+IHYldryKBDy6BdxqHhpAn/Dj1+
+ImkapiBYdB7l/VFCotsEk8o/3kuYQnrn1lrEtJ5yeeJGj8R6JVG3TVMW+Op1Gvk
mQf34OMq1vQ104RGX20qtgQjuT3C7fdOLxocS4+bYP+zY/L88FQ3taaB+pPoD+hb
YtUy2RBH+7Y+DIBEY9uR6pyyQOHE9VX5ksV6muxbe8XflJ5aVwInFjDJdZdG4Kg4
a3Wab6pSeNnas/zOtAi6BD8gbwQEMIzPzsEgBe2brqn3psqF449KSm3AS275dB/a
69E1OEOZGpesfhP8Qc+R7nHDUe8/AoE//yePnZtKsX/mgruzWu61G6VMn4j6bH4B
TkmiaAUWDGpokclNpmC6NYJtT88TfocNJV1tkqbP+/NGWVnrWSpI9HIDB9oh4Dsl
fhIoVBdIgxbEFFZyY0USHwogpdeNUlAyQLmIg6nm9otEa3yBLjMvc5Njv7Iy3XLm
noAIJlyg3D5mys4GqH/33g1xpk12IODLxfR9NoxR547OqYiu8EmndujzSqV58Jo7
eJ7kDZFLI55brqZTYNUArWaRraKjmXRjJDdfKiu/ONeDjxqvpffdG35L28tEnwoQ
YtRCA/R9rsRYBzOQWeiRVG2nSUQevc2jcpx6PaEeY7y/xNAYMR21kSiUOao0W7x4
npwTc2UNgoAlXDRtYlTYYs7QDBiMfkLXlfyHisRwGzqxgTHhg/dfv7uRsCn5wuqs
nEr4hO+HQs0sAzuiZLqPv22SmwRFrS1iQ0vV7OZlb48Vt+aNV50Dursa9xc3Zs1p
3NKZtEPWOYu/ILYF1N73825u/nfiaP1cE+zIdpHBYDAdA18HPgHq2nk5d4UQ48Sq
+sNcDkjJ0T55ZN4XYPispe9k/zS7D+2GEtjR+BK5QkTcBAkTtd2AkwabgPBgxBXd
0WSuajH1u+/Y2ZRqBY6dHSOAXlTArUHpa0F+Z2uTg4S6n6ZSSu/8vPAN0rdHGrYw
64qqDCEMIOBtXKinrbmzq80uM5y534Qn5lO4SmN4W3AKICE82vrNRnuRsNZMbxpk
RZAsuSX6QATBiQCgG4m62B+jq/FJU6xjhcAiOseDT9GpM+2M77UaGc1/5UzCvW4C
WDWDGJBY76WBbBKe6AQBK6wWW17P2AyTC3Mhcgr1kpU2YppiZk9KAnvFlyh0PsRE
zIWkoAaAKtMApwAvdef/9Ku0iOCa5XsHSQdLP0uVVoyoJDNTg0LJYQvWPS8bvUI3
YaBsppymFNtCw0tL1l9ySPwzEjNcxVEVD6ecNMg0M9oC2HcySdfln1uF+57G7vPd
Bbujl+vaavog8IManLit4K1ghi7VqxLGszv0r2RzuFsI2EZ5vT1r3wHaWLZ3saqE
BZzQvTh+L99FXwzXK9jsrWEPliS4uFVjU9KbY3BysEHjECl9fJMhYrAnYPo2gELF
3Deey9tb5En1/MH4I4rn0a4PDUvJDbYR/CzK41c2QTklPb+bVMBRXyK/+SxJNkSN
IXB3z4z8NQpRgnvdYCAziPCyGWTS8UzCF908RjomwyLvsLeqqZJOk6qlwYNIbGss
orfZb9p8aQ1zZe1LzRfTyoPqa9Ki+SNvLSdfZIJqb9aBH0WMzWrerUT890WTI1v9
0vSHWO/zpM/Mt1/YL6gQBhu6swvCh9W1Wx43IiiT60nJFRZQy0SwZUdpzxJTFtAw
OOSTH/TapLss9cxF0Q+Icqxj4hPmHRrUzAxkR+zvMqvX+RCQtAk8HnbnSEhSy5Fv
q4qVBnpVBnUQMg1coea8G90+zfgcDXPZgQ5zEJ1gnw0HNJ0ecQtT2VMWrEMDfci4
32kYF8DrZpVZWwGDArdJE0TQLTOVlscVykCVj5OSdG8i+rFK1yiJH7mako2RtPi6
jBgJkBryxGzZqpGF+BnbEGQC/Yjf0zySkDf98tCBPF3FKX/lqpFJxmPPrp9TeTkT
WO6qvOaF8b9X2h8ct0ifObmwPgjQe98FtifA1FjB+HmEobUsVktf43WEqNG8Irhr
J7LTlzCX7UdQTT6txAY3UvN2h5ChyvSfLGZmX4hIMhVECs25fHzWzsjJkVz/cvCQ
wWcyGfBYEpk56qSNnXgjEs163/5ETy8vZ+a7pqOOXHROrHma//64wYQzAqYzG/Gg
mw/O4kQF5h6g0DwTri8RnXlFcGe613fyaVRjigR0rjNqvps8H8QDOSud1OPDmiS+
X1rb6foOD/Gw9pyLXdl7Uf4+fa/Uh6C8ILIa26pMh0ggF0WPtwXznVC0dVMyEN4i
fqiLB5CBJx+Y8rCTRwzIutbGtldRYz/zVi7ODoizhQCBJ+zBXgdCPqYaQ5ssxVR3
fIWr5P380sE3rU1wq/e5YJ32b7AWL7tOzNSOwuSg4OgXP5ohKu3JqaUabt+OXJkx
+ojf5jQ7D77JAM8xzwLriRdjqAnu2KIzQ/oWvqh8d50ouBml1t2WZtRhxpwfx3xC
IhPkFIZvrdzThz97n9B9PYVstCG/CaGLMfdj/741+kF2pj1AMl83UktYV9wySKay
GmNdAvrH7rm35usda81ehtT7Mu67WshTaIRUOw1LtgV/31i4RwZJU99OlzUBEzam
2InGxYHrPNJ1CfNheBJKAqdjRfntCdIHQ8fs0a+UVEY7TDlZ4JFnc38cNUcUD0FK
Ngb+3et4jbf7RYCbchBjfY5GATt1mDyK8sruiQ7A6gkiSIIgSVb3kwRf9WV9N/u3
JLMD/AQfYYfhX74FNboJdieR/iDobmQ15qwArJi+lEEnM5NxeFxJlfrsm+MkYLHu
rAnn0FXtA76I5uVgdjya12NSEq064Qs15tJxNdKzx4GzkX888M33v0kk0WY3AyPT
/bFrN2LacGitIvDEmVlOShRu7N0GfQmqeHvTkCV2fxK2m9SGNF4VJdqrsNu1IsDR
r7g9TT4yclHu8WM0QVOVVjRpfg33gpblmdRL9xjhuJnLfDysuYt7+NskBT/ZtWkr
Ccd2lIAhoHTRFvsRUMxgdUzFfOAULhJTpZqzBwnCXgbAGOuGsrLB0UlC2Blep0fw
SWWrKV7h+IjyfuH8NSmOVQq9t+cHgF8AZPay8V6D+lKY0omXaXW6cY9ttSSnD4Kc
lVjUIp9VO6J0+z2+7ZKle7lU3iuhAkMQBWMS5yHBjoN+CldcCLbmWlhykDFKYvGa
FahhYxIsDa6X1ICBI8UlmOPFr/UYcILNbj2gKYLqWPF5RpDId8uqVb8MVQ8O4cbj
mkjL46pMVJpMUdQ4liqHgS0GCid1oWbY4Rw/YOHbHm4wkTWzeKNXRtq4kX/Q/Vhp
hN/otRL06b9FJbOIcQpitmuXm4jVr/175OUHB2lIQnUuoPLkU1QT2a/YfiM3+vH/
ytZ+exsyG/JfEwIKv3n9j4jLZPFY9f5FfNEoL0rAavAY2adVtdvgMv/Y+0EKrudL
RN5Jt9nz0+F8fdchg+dG4RSC4KSyjD7kIMQH/QVz9OSjkn08UoMn0jFr8htkNE4S
kWDfwlFduPQCMuT7wxL4cCvhJF/kJnadg+TFWZuNke2EuqgxGWUsqCO42ob6DJsY
8Mod4B8BGjg76HaCmTBDaSCFsXNF7Tu8azjMG6SrmPZ4FcwUC6tijkPTWyu/VLxC
fOJ64CrpC2sfDTOEyxHbJiJVANDGyVoy1Hoe7rTn9tUJEOir3bD4dbDC5BwqD+iw
xUwmw3X/wSrzTmniArKG3/bScpRvMVfxjZUkJuMrpZP33eloCKx3/Jxe0vCAmlhh
NZW7UI9m8GiFMjWEARrTgSPeppYcOW0wkS9ShwEvMrhRzb+SFsNqzlXpWSkg6ZiT
vPSwd7oOlGxtuxxUOrQ/U5pc0Q31/IvcwyO7kA9bTiXxU3+XcDDmC0sX1te48DI4
4MjjwkrZSCLonISBnyV4sAXb/gOaihkNRDGGlm3pKgPliq9XMnkHcOPID5I7HNKh
xzsFLu31h3fphJBmbNX71LeQyGFhv/RyeLy12EREGkdIGnXzrQljAIgUAHi1dGDL
Ly0P5rXybpf3fFlc9lfRSe2npit/KKwJQwZ5/RJVzt2wZ3jNBxj79F8yr/6Padz9
Jr1mVynqnui+JiJzI6uanXEm74Ge8N8Kzez9NA/aN2Q3tPHNX/SAS/UNXOUfXsTN
iF7qRBSMQXWyJqqRxWGq6I2g9STTTLMeus+jJKXEOgvN8P3r4t867aZFlX44JZep
aHJXR/Q/xoJ+ZPDEiTHUpS866/I2HTfdyLJoXiq5vz47FFpdC2zV3GdHi3cKbS3h
u+ABVLwKldvZS2dCXHo3gaTYatnViQX55lf8JyWyyQW3p/oIgFHsrEAJiWm/q8KN
ACeqbIICtUnPPGhvj739u8xAOLQ/dP+vKQKmWoeZWLBGhJGIssXlF+sVzMvDFdDP
RIQn42cIysfHM1d6T5i+phhr8mRYQnEnCo5B19L/KuA1aU0oApZsMYAxGmkTfx5r
7JgNYFtOYWnXE2+S28RR7FIRiYvY2jD1UdbsNi8eDM3IuDE2ZkuxtfPQM0cE8tEh
06JFqfgmcWPPL1aYEvUq70rW4xZRYqAN2d1Ssj7hhdzVftW/q8xIy67HB9YhLmu3
HztK/xDWmoznzBo5YC1LPZbUwx5pUI1zyTEnIrTnPxXM7y/IOkuWiz2smfcjHp/S
O/vSLwPhOD33YUE/LntSCz9KW4N5AsMGGVQUMy/bfrWwnENyJRuLYw3xBHKjGY5C
Cjq6JmKpElRbEnWz5SsUkYrElngXDxGlcx9QjffwrOO/A9u03AGKlqIEAX3CgLeP
NqkPX9gln+2jVQTL9LdSqERnlpM64qJQA8nMb/v4FsOQ/OWwb1oVvqt2jG5bie1P
E7/jW2hkB+qZL8NmT0QFjzigQaYzBbfQuanFTeKaStBwsfdAIbKyA8pBYKfL0eES
9Thm5vbuvZC08nbtClv2BoK8dEJQf9Fq/WOY9aJBEKt9GjlhLUwJcx9D/YeLjz0T
yuDbyZG6saolT7CeZS/rxEtq/OmT/F0XghtTCjZvxhhnFmum43hD7sxmZfHOrQ5l
vDFSUqkq5Box8xI3P7/3QTDZgDznpOBgnmCZDXWBsKoIw2nx0Q8zReBGIIHOlbpP
mPCnl/p2KM9R7IJZ/HGK0CvNTR+KPkyN1UfNyoRGYShMPLFAyiwX1Vz6juxt+l2d
64Z851vVbKs3/HMl3M+WQDQZacZgdtSePloi0suPCB7JgTdjabvL9JKkIXrzLOvH
XGchFBpHFmbi6aKPAWgP19xVCWot9va8t8/BjtCJ+Zo1qa8Fvmr8teAqEKnQYfyd
5yFqMfHuoa02gW8OOlqM1mg0mxDImniMry8ORYcV51YgP5NUSNTVCUnOncvJtVX5
peqSgyI7p+hurFGAlWhDTH6VVXgftIa9owbXQp1qp0TAcglgi1WQhBNONHkcvRl2
NhMmPFGPPa2FJ4w2PamVL3O/lEiqJ5rHxNWtXS2iBH3EbNFLPRgVzWedQrAOwQbQ
e3BfTlvMv84demX1iSt7tBBx0wcNbfvHWtdUm9Tik8pAAnCg+hwIO3e0g1AE7P6+
wpf9+UiezVi0KtOrvY0G2r/3R4xGQaCLTWrjt4cM+mO+gvFsPZwOMC/HXrgr+sG6
wiPTpYr9yYEcfgEq2L4leQ89Z46EgJvrsX5jJB3kcVPhQZXUwZ7tdfaVFHO9w8DQ
yyf7G1qDFh0bMVPxARzhClKHS7HuFNfsGS6Y3awUzQvUdIS9eAGGXZSYMVK9aZ28
SwtW7x3bgo0IqiU/g1qT3bgo2n7Ch6Jae5iCBVyyNNMyh0MW2ClrGZp+AT7lrG1X
PO12aaHhZJ1Aqvbg8lST3BdJk22b+zv2pApZq0yYQXAEe58swaAzxeO1m17WCSIy
VxpicPxdnPtt83YoRHs/bkFfK7gokFUZXHizTfpqFH7odUS9QNVLaKTQ2OWZ+ukW
f7IAzeCmArpbTFzdaSp0c5aXbCStGwP6dJevEg3bdgPLt/qjXdhJes2zEU7R2fz5
wkLFCR/BMmlzQ2mk4nJm/LnF+vjg4B4Gb8Ci8KVveIHrTqis1UhACbRmC5u5QFcz
hkERW2288x5DcytXwHZe/VsjLCERC/RD9yc2XJiBw/yjlhHcF9nra3kSXgmPI0J6
EMH7pH4rNwm/fIp7702Ymi/3Yw9UK1m/N23AqM+pKNTR6rPNSNFXQyxWF6xqaGFJ
HstPaFOWV0N1J2rxX1cXEBJlJeBbW5jNc6WduWDFXYTIUetad3qL3q4eTqgKYhr0
Y3hUAZpEe8yFkjB6hqxAkZ+p+2w25z/f5U6PlvTn2DpeJO3cJ7EAakkv4pL/g04N
Fb4RwIotpKsdDD4JXBciGBQ0k9FyZab8TJAWraqMyOByN0hLWI78n6BZmoxBkvO4
MQLSvJ/V0OHPjtLGJ6LIiSt6MmxEba9/FnS++8WtBMVsmMuorIoCGdNYoN4j/5EI
cUVIoe/c0QkcVKrxs1wbTEsGSscZ/5lIJM8GZlLWW0LSRdQrSLyqmTP/eefZTzl1
WbPewNcdH/BkLmEktm5MJZhXdfx8EAAk806F2gs5kUk1zwN8Hgz+9iVSwmb+6yRN
KcwJihagZp8TBt0hdvZGJnEiMQzVrM+kZFZ3vmCMn93O/Krm+E/ZoL/vUw4w1uAb
8nOIP2edWgnGKxIaQJ541WwOawKtvW4DzxJcA7YE1oCXpFFATRt83bBU5I3EZ2Jo
IrTCuiL00Wkfk6PolMuo3EGLme00CiExCqi1Xds361JKCtimSr+jEo8zFKPYutJY
jFpgwdgnc6cKJUrYp7BFjuWCUCfvDPjpchXmoV8M+OIDztnYSE+z3UQbxfFrjZS8
tM4I3751ev2g9n+L9h4wKlnfYWTgKdOSJ2DUJSJum++KGZDj9Cvuy6We1t1UMlW2
jq3PW6Uuqk8BQheJhOd+grEQNTx76X/HNC02av0+fsxFU/0BQIneJIkQWZC+rBgh
8eq6dYeh4Uiyt5bxGFP646WpfZXuvIhOLTj7p9a4Bxes6bX40MW0uPwwDQ0kOf/O
qsbg825sxg8/edX93V6SbsU15/8xRr7UzkmiE4uIp9MtxU2JbugI6itb0+02GlWq
wYFyEfGm/jY9kyoQkERSBmo66IKlCQtUBEfWK+njs+RxNJQ62uJnm5Y8KKfKymW9
CnGbaHCO/Iq/LxiCg4AXmKm4Me8GVs56nXm/+wRUTfC7m6Q4QQN49xs9u+za3brW
O//yRuRhyBhJI2JQKqU4eTI2e31DZOX4nd0I+pMPKPannI8dnnfmh1okYeaSd7Ue
t0x+UzwPbUtsGuwtSacgFmtj/2GAzdwFD+J56pvluNA4L7Mr779MTjPx6a7Grtz6
2JOmgAtiXOIGjp7yFTeLX/k5Vgi84b88A4z7Kpl0q5DhPg6YdFg3IuXRIGU44XJ+
hzPHpKKbRa7Tmg/iIZmP9UOuFQUxOQcG6cQDawf3XQ64DPgc7q/KuiIAA+q7aiHD
DqJ/Ms+T/B2RePeXsWC4Zf9hPLwzcyyLDQWTQHcUfFhl/qUWslQUCdA3C0Cwoa26
9+RFCvnsoQVxPn31FS1roINExciP4KF/uyaKlGl+x60MmWDtkb7raWkLp8nUGJwV
YnQzQDuozNCyxSDaMP/qagpD4x2pCOryR8UGC3EzMwQxbiXKaIr1txcK1I5NinUf
NGUhq+6arwPmv3PVJhbbBkZq0PCDNhnahS+S8dfMdmpee7yG6n9l+WRewcozHXy6
HQS1v65HzSXO4+1aSGRR3fO7ZV/7XNAYdyVbqenqN/FUxszPhoF03ZcMBNCgl4LN
/j2dHOasdRmy64vSdxZ6CE6fWra953R+l91PLgIkvTyVStUKtr6Op9Gterq/A/Lp
hxTw0GQb8NIEkNxnWv52Zme9eWhT8PbJrjv+J+UKh0B5Th7WGYAdJwSCKDnaOV1d
S7ducOaa9aJ4ZHAPH1AQpv3Zj46wrWsfI0eUTZVlspkQXzQWg3+RAbbQ/ElJ2WRm
VtjSi2UmTr8qPgS07R+m2+8HS1XmjZZ21l0pUjjHcwPjHB7dsrSlL3feBekweLvA
8aUybITN563YxDRXfIWNCsaXrQgbi60eJN7FRRKMz9KnBHznRKROytTp9HY4zoCp
arYE04x9Eql5+gxAB2vXEUYWBJjKrVT8Kz0P0NtGl8rKCh2tFHyQJpSvsXnwHFW9
9zUQFZSOpbOS0DiQRRy0WYbld8iiUz/4+dRgwshA75K241nEZ6LiqU3WjdGa051y
NAYS0t7B91Jevc89Pzq+R2RyPhw0jjC+vAAPsflw0UdQ8yR9HiDUWGWY4+t7jGPJ
Iw9DpQTviFLaUr5TcFZteK3fomPzCbTS5m9BEqOP9Vavn1qmAYTPZRvhBIt+6FqX
lwL0DTsBs31rtYdwjSwbTQhxXqHjEYmduu6y+4FRHv4s9xxm2BUzf2eUIaC91OXi
BQifwiXytHizibr8ymnL/87sELc+giOgiTb+U7tgjfrZwlN13v0oGdXfi0Bu+90h
8irH4UvIqh9qHbJwwr0jix90F5wD7KVuKdtEAIAv/gcSW42Hg3T+VpgS7wjbs4PJ
3ALPZWD13y4xjqeE2rOUKqnY/yBYnLFLFvS5iXORdOfdC9kuN0TjCLRFVTuCz5oE
O2CV+Rhz77vFoKNx7uagOHQge56bIr2IxfbeunF1nC4ewul3sSoVit5utYc7Xfht
vJs05bZ881QUIz/PBS3EYxgydELP6s/LfRhdaGwbBu0sXQgo1bV+c8UhkeEcxhAB
81GwEdnnH9sr+VT7jtpvs9Xw9MdilFpRl2QTGPJvFj1MQjDl2hDUU7AZxVkRABlu
IoglA+csTysxiqb+9G5cR/beGO8FmUMmK6NRE60k6nqFdxMyOYinljzZk32a+cBG
c7333osJcYxeOFEuoIp+lFCics1O3MnELtnYKg3/5t90Vm4lb88FWhKY7J9r7SlA
MDP/4qBPhPY1JdLljcvyVzaTxmxbge2M4BRyzIDbwJ54L2rT5qmc4HBUM6AzsL8h
8Y6X4ShIcC9CdWYokAIOnBpR9up20dtg/6YV73pIoGqMU1lejde61oN0ZZR2z/CJ
KzR5N+JEkm6zNN8RIdYY7MEUCz5b5oTP9uMzYapqS4jx5mEKmcKfgQJ1fgnuy3hH
BZxWr8GEg07vOB7tWcPK9F3VWNK4+RSLcKm4xQvBXr3jaxqNOV99eCM3f84wI9TQ
pcvMbbcx0iUhpmVdHcT5PlywTccj3ox3O8Ju+zOUaXywdmd1HP2alZ3iq5LgcDda
RFaQ08+dkJcU2HqmHNln0nkUziqrH5GM9souNmTMBk34GP9kCdHBJaL3H+ree5Sw
rKki5oD8p8qNTeWMDWM1DvAh9dp5ndEa3oiaJZOxHXdSsyJ00K3Tz4RKqFEsHI/d
4o59+okLvBVH0FKZNvJNi2DW1ZEPqYRPm8D/2OfvYmvZJszvnxI06S68haGpiJHo
F0UBHPzTkCBM6MWYtth7ex9eCijJK8rtuJtSoHJX/FUmjagPiguUwnAyMIu6Wydh
4upZSv0kOAioUEnPAtkJVfzJyaqwH6TD0ncM1SZtrh51bE4GnlrvRhNfZjjHsPZQ
xbeMdha8Z5ljA5AIZTmXPVvpvl/wAjhJLs+rmuCtVPfQdDr0+UX3dI6bOdtWt73C
39dZAuopJhaUndjTtb9wj1IdAWVH3o4ZICEfzceYxcmUtXgzJS5Llh3LfAYGrJAB
WvSuK7VjrauyRd/ByQ4hp8vx0Chu6QNCePKPwSKUFDfzR1rQFFL06X/SeQ8Jv4pQ
7UjAuCpeHC5TXS7/1uCWAjwAtugGhnAy92dEl/Jb5SCrzxPgDsqMrmuYKl+oBrNq
Ep6CBSJe84QsOHZJ0WBGZcUXe/7MVOuesmQFfY/snjDcZ4hLpF3/Ia6XX/diQTkZ
Z7hs7z9h9nRLVjxUaiEIXIrqgrwPLSM2APofekD+lg02n93XxLeyn6JatmM1rPeX
qWCHBbU7OQLqv+QQmj63IS6T12GJAe0P9COhtbAdRsLipTzFdSkBZ/75zK1u9pAr
rZQLxSLO9Nm18My9hKqM2AK++7wBURqqK6kPxkL5zB3FcrmL+x3BkL/RVa7/Niof
myBcE4c21gGcXO6xjjqY9PeTO/put96EkFUSV7W0sCHPq3XL6Yqw247pDS2RsJTt
wP1B0sxdXucrf6z3Peuc/fnNs7P3dMmHX57SZfj+xLQdpQICsczg6y01HkKaMoue
cF36d5o+qFsgnvjPAavjbV4MiQnW1AFvOrLfUdu8pLChv9zyAPWUdPbZsTbddsZc
otvYbKyRBs10MCHyAWPb8I6FBUAgHgW39PetuN0MaV1n0t6D63QPDXT+C5GoiGJ+
ObJB0HdtCORJ4NHJKnpHWhB785UC0AVJXi4cxSm4whnIAyBWhPIvadt5ssAPkbUU
gga93+PIw2HfNnBkaBRzno+gJQbks2Ipa4GQ3Nd+y/R4Yr3R2WGS5GmyLYLGeEmJ
oK7U+ebLWSJxhmH1/+3PBzcmNOwaNtWkn37l11EgarK82WHFvcCDM3VWIQoarMX3
WUM9fPOpsli0VpKATqT1CTIqEy6hi+m7TbDO5at6LUVar8fhRkieJPiem9bHCvPv
UvXhUpNNQtMNdwkzDvw8qxSxd2y70A6Q01CRbJhyTFYKRu4ferYrqakBjBw2PER7
4fxATUs/EaSokBHKbv0yjv71YvwpTDcHL2v3K3ZWWzcT/Zuhv6ZT2yFr26kq6m42
FIo5WNoMX371hX/m1q6Zg4kbARxR0TA82UkSG5gfLFl5wJn6AwPSGsFp1WJagr69
iT7DtRsFNCp7YZEAVLdSLOtQwQ5zcBQ7Wa6rDk13pjfusTMXh9IhIesnBcUeLKfn
rVrdO+IdUTH4qI+sc6tSO+LgCgB+fuAHi8UCnLtHRH26yasSNIF48IZbdVpfx9GV
vqoAqVYwr9/8bwc6BD4eqPxqawtrpp61FQXpJiTCe0KBoGLr06PIpVZBHHLMrLgp
WynNggCSm3QlL5FURmeViHT6qHnE4cKNsFVU3W4HcBXowg3MVFjDbNoiEVVzM7ed
ZaH/g++RF+FG9am6tWLYAu88WtFJ0LrdGsEZv5Dj16mgHqgmQSRh49lVH71+toXz
XYCr0z9bf3v82QaBJmBXADb7o/9GYYrt42JcDq/7K9MsvPU4s8dtx6xn+VSI03iD
+Rk55l1jldKBHVaV+45crkWFruKW/Q/O17mU6JTQh+fEOIQpbHsEKjYQiO+1Yyb+
0jNur/7PRrQCtP8ten94qmSU1TcxobROUoW1XLYkFMtTmf5pdI0fXD0G5slt+8x2
ey4n252XVTS3v2FOq7H24SxaXhAPVKeH/jHUzFmIctZAJcAk9MLvZnwJmbhBGmsb
NJ5jr8NofslBJoA3kl4ozRH04jVMP437KiQ0mk/EhuLf0z9vyMFGWueDTJbzAomG
iP+u1MY2+ZU07Gaimth/bWNJhXab1XsvHynIMz+xhqyMggKa07xTUg46n7IpRh+V
QmPhS9feIBgFYdRdNE+P/x+5rpXHvnEnQKd8ih370ON4g1Rr/Z8pkE52Jwn9ZcnC
fTpDzKnCIwgUGAjiPblIa+k1yOZkXoh8fWsPOMpQA53cA67FJR+ucb0Lw3wUZpXG
gdKtmkeNYyM3tOZoZPFTpnb2uT5/wUAqC+m8fWyA/TA8jrynfmtTVOAz+ffGB1Ha
Q302rkJpsRqEch+KHZWNXV0Fazkvco/8xUOc8nZP3akSzJ06hJjURuKyKhi83EAd
VGp5wEexm+L0vo9ksbA9GlrDk+avPCvGgS8YU6cQLex/3kIozd9pYCicuWM4PS64
4ceM5674aLqBZngV77hx6tZ1MZiz3JHHOq+6hp0YV4bLkTObVKIvhwxiKpNr4W5C
DBwCdKAlK0vtx+O0Ib2c6SRjt2omsBome0mjbDmVhMcPekgyBuk3BcJ6deWAVHaP
6wtpmov1grL4vRGDZP4EWd8c4F5jviEch1jA7IMDuX2+QSZHQ9jV71GRdPR+NPiB
MduRzxnvOubPlfvuiJ1etHA2s4ZG9wZJOhnQ6dtiEGUai2nsbxW42zwpkeCLIBUR
y4PC7Dat676Urh6RpbUdiNxTZXNintoHan/LPovo2ucUoHVP96Nf4LEtcskmFNsb
mxvWqtawrLkKyOVLmZRo43xf67hD4h7tkjmq9g8l5raVFxa/cSdl+TqXpoQ6e7n+
VrYxsLvy56jdBB+7XGFLpflKnxBuTUY18Y3HpFza5FG9+zEhudNhpesz7q1BUAuY
W5Xi0WDkIHcgrzJ5ZJvDH9Ch35pZ6e5QnKEIvD5BEGCKwS11m038Jah+nuesA7ge
6LmjfiG5O19VHWKhwPwCllJz3ue9v4G2I+RqUJWXrrreJSaEjRH8ckDUtH/pvtIA
zy6bzf52Wya8DTpXEJU8kP8/E+cPMAWYyXEzuq2cnZmfNXpXSoY6vu5JWKL+mzD+
jERbazxWNL9W7eO2ksqnk1DPaZ9QKWGo7QjCuAidaOq0j+K4uZEIrAD4/R/yBBjm
Z6VPbo3KfCEcjkLyUTEY2WyBuNBJZ13xLC3k9rPOxR8TglInBj0KbniBzHPuRFZr
Hncs3Djmqey8SesV9SjCI7PhwuQTHbgfSJ6nBlmLRa03xhlCVz+NffUxisSobgCp
frX2NLczSKlGPXRrQZwq3T5S4tY+PFWbOWAkwFtApJKAq3/0swN1oJfK4VoVOuqr
GI9dseUdcRgZqjzOCuwaEu2pbSyc5T9sXbOQWp3r6SpYocBVGdHu3+mE4QYkF6R2
qezhKMg2J9dJM5Yev5JxtbEILCR7mCepDGt/NpIJ75X1WeYWdaThHMpawZnQYNKK
9Wxt+coOOz1TfXIh7IsczqAK5tBEZCk8ReEm9gMEFdNGdHgp/JiNiX9BHcor20CE
sJE7V2U5CeK8qZ9oqjBrw65DtVs26/qo+ZOIqPtKlJV1ohijSHlrpaMeuKrb0f/q
MbC81Wdjs9GWOxpz5qtLdcfSsO/FJoc+opoJoiO9Wp50zowprONf7CSEOR6Wm50q
wO7bPmOIyJ6fNiTwcrnpABnlV7yITeKNlRPokHUPzmxDUxenBYH02fjK6V/mQ3C4
oAEYNgym6ZayDl/b8ANMLUVpkDj5DCXuDAuWuD7D+0ur0qWoKNm/8aE38jsUJmUX
tObsgkp8fB5aJ+J+Pqp59RbPg1xyG7q1krSaxntYVhA0nXYqoHN1+rhBZkRqvCQN
+DXAHAJz6MCbmXAj1pxO/EzaxpLe1OE5AqLiEl0TXQz2HNR6UbYjlmUB+7aoecHy
8QH7Bv3Z376YN/R335FQg2Uyt/QrncVZwfGlnXrlypgUFO1DoYncfuPNOlL/Ci0v
hrY4SoM4YoATo1JjWOGiJ4RMjIBn5ctRqskcC53nR0bUZhPxC3Ny16utmrs7kSHG
bY52vZyoP0VPYWbC9OHt0Tbl45DmuD/MyrL39YpukLDn59MFGWZeA/3KllzdaZtF
iRIoyCOknRSY4CBlQiMuGm+gU2oWB9VRxTbgJ2DGQfJOJacEzV6Fjerlr1/0l6+v
CgqC60tnxvI9qQ3Zt0NHoD+yVnX/g+9nuor41lO8gzoWytBIKcBve+kCpI1P3cuJ
1ZzmkDrpAGHmBEFVX1RdVvm33QS96thMb3dTlNmHf6bY4GhopXxPKouENWy9g0Kq
AZv/yEx1cSICDdU9qY4+EcVfmQ89Fr0NXQJ5b5VFusterAkR1hDNVBQ3Wgt9DonB
BfOfOYo8BqVNMhQkwEQhCNr9U59CiAK0MfrHpPjWyvSbYF2w0v8OFaBwr1LzHbla
zXcdtoq+1Btd2J+UrbIFs3Zbn/EIkVnsjrWQ4rQR5hMQdY9Jf7qGWSkpDut/+V0T
6OuexMmH1lNpEsW24KVrdb2iduv+QT7PuymUbnc20vjATT8kZYyEUFyG2ETkKtsg
tb1RT5odfPKvoOw6qv/R/piyJLfag5eNzar9mjJzZdxhuaTDWVzAYgjzj/j8mhpk
E2FOHN+Sp2/qjXAEGtnfSSIBQlxoszbjbVFDhn5olj+jsX7fG1zixtYylilQnEQl
/pySmY1d3GLE4t7PBKNWCarmg5H+I0J6GkFsF0/IwjibDvDI8tiuncVz9a5B37ic
3oujHUXZ/9YJPmCCa7ZK7ZbL0TzmU0DXCylJSG37J7DokK/tf8IfdvOINeUlsAL9
Ewo1cHvTIzwDM9PiezKSCI5tz2Qf/IcNRF7/8yLn0nQl2WmrySIuH1dlnZVojrnJ
v0h86KKof7bs/mW5eyE2bfq7zYFekg6E6dqZgltDYOU5S7xCbCw1zfa1k3/BW308
ecQx8KvqNiBPwvOftltjbO0aAv8yTO8uE4Jqd0mERkTI7x0IvYCEmlAeSQroLOgu
zQpdSWtPpEVGmdtuNvTfSMMFpWeMEGHQW/SSU1Q4Tewsk91/4B2rdq3GCCyL6945
ZgeIlVIKAMzRypBQl7RdWBJg2gQboawoAoPcjK2nlxC7isVzh6xbNk1IGVHKikWF
V0btOx0QiEf5WZEx1RfH72dppOgbniDUPqDSNyZafk96lkxtGSeyUQzZh5kiJ2wR
6Y9PNIFMFzP/TAD9YsG79AdA0r8jZqMEBzJixX6YurIyYRSIE/36nkLLZ3DOu0ii
LyIvE3HmRrS3Y1YMx8Xjp5z6EQsGtPAHnpU7ivu2+47m3//TvYf/LJoEZlo1Q/ul
pEvv0TycO8Kch6R+h+8fYjKX7zVXnhieS+QPyUgVvfM8UsAyxzqR2cWhBcStsYVA
pIim3AWXD37aT4YdUg2PJeDfR7dHRDYngSCkJAjlWbhc+mvSQwWaXOFY5EFw7KDC
B7k2kcxmJCleRIa5kUqIJff3SvPPkpmkmDbjPtrfiBIQqyle9q5TV/44VQYbVu74
g3zW6MtxhLbLU7ioDF2MZHyRx6N+gXVG0SxhLNXxcEmAenORv87vOmYRxiY5NBAd
lXeSCWcTNYUHr15bhBvnqk17PcY/H1DrjxjN22T10NSHcHhey3ddEGqGNT1bJ3Bw
rF5/Rdk+GWTiHoWNYC5z008V+Wfj6O9nZ/g4PQdDxCi596P4WtHX3T/kSD3zLjwB
qzdoJHa2IgUOVcWlblTZWtQK8pGyas93/pkFgv8CTy6NhPksP+Sw93yp72oyn+G1
21T7EjzlJJ4MohF8SAGQZlLHBbrxmBwtzA7hbgUr5lSuv9RF37h/CQ0Ds57mv6dC
z4pl/5AHvsprAG62JBj+K5Fim4hECEszFUJJDVQUfpFxLEsTQXRn4LQEqyTN/M+I
laQ3mDSz82iTyEueZeKlbkz2Mqj8erWHZDGt+0fZ9txLh4Bbac4QUQLhju/0xHuI
TWhh4e7fIwUGm9sf+ZgBpRir7mmkWAaWEGkmyeByJOe5Ad8lMcKFrG5kgqsJ04tk
HPMSdQ9F6TqK5KqdZRcdV5T5KuiwP4AEcJhzMJ95Yd19OTTcv1/Ak8y182wqkNpZ
giyRM84a7eWZy8nFNF2MKOCGFxlhfRHPcNsbygoQbMPAD7eFU2wuB6u5MtBChz9E
GhWXZquKVHnh3GltvzfSRrSKMll+6xjgDgoahgiJhd1AFzpQATVJHmWPlEjwbXpK
LpzGh2ht0gWtmJETFSdl7u8zDM4HtwW6S2J/H+dvi+UqEvSrHuyTPTHC38NPxfLZ
tJdUA04/w/RCatZKZtxHJ19RYph+6zRjjuVuUcV69s9ZKZ1TWBZBjMr35KAkgIaJ
WqDmc47Ut3FZ7RuNaIOI0nwYe2H5zNG1hXVgx+xBiY/T9DNvU9/EFIG/dRLKn8HF
HIdPK39eQNM3c3tkx/p5y6dgs6wH+7vXc/rmkxPmMmdYBGOqnCpThA4MsE/Xer8i
opnvuZ41DygB0lgzhE08QtTZohfEXN393Nlccu2591HD6jxqVx2PYVUs+LE5fDH1
CJkrx0wh5sBSPwzNE0hqPsBoD8oKZE8usJ8JzpFYelM6SpUvNNFrqhzvu3irAxQE
wOvrIq1pcgDIWY4salIuF5/QpsOMmU9yA60VPYMr5nGKPZy9RDRiOCBQZ5a5U+s6
RapLfydVYIIBCdSiddqC1NEEJOK9fkdTfMV0SKXpgHCON92WGxcJOjveO/k2acMN
1hHwQx7a8vlODr7qbXhhai60IhKnMDmXYvaa/zbAwY1yss1jgwB0f3jKoPBh+qZ7
3S8RH/3v3h8Ak0bdeYiCIGlEjntG6NWRVdQ+lqDQAKrY1fy1OYuDHfn63zLegLyK
BasBIhP0JhF9gBj8jqi3ch+Dog182tRQiP+VAnvYxfFmpmo92mvupOYSSI1ae84F
oY4V/8NN7yBrSIq608gbEMmvO3VSDPwq0l0taiQO9xP2NsJ3wdHOrC73o8+hNiWh
ma49WCLdlGAVPDJf38F2bP9wBuuuXxRhsNyku9dAoNCsG7CG4DHf+DKaCM122rNL
CrInZttLiHi8dAuM4za/qoz6i6tuOazdASi2CMDnnt3cYgKToZB9FPksEB5deXvs
6pK0znkLwPyeX5hAixd3t6eMwM7n+a6LmZh62yHS2I9M/dXwlg4ZbVZNt/kSvMU8
+onkSgGS0UgwcIOwZxTdZUKsU6vnIWe/9GYXRCDlzhsicfJ4ox9LcJhjVErWF16F
vUFWp6uS9HCg/NTJQitcKtL0gqA/RVeu4gHagcC1hMuazPjNM+gr9ylO4BxvWa8C
l46lRDI2KrZWXiM1VVUsoYVmG0MXblEtKW2KPKzaDZ5mQAQc1NvE3quTDjYHksXf
RmR4h9GqPJMT5f00avzVZrAYLMFoK7lNxc3UUsWRg3eQdb28UXt6SYcztZnWTuJE
irTBuvRe74/TEJQbL+tShelLa5ysUD4WhxA7bAu1jM0NfLzI0wWltYfAi3rxlGjh
dL+MwgzsBJzFzw88uu3CLaObildvsosgOp7AsH9BEanQj7wdPaPlsnnfwZIo138w
CM4yQt62UC+U8YEdmrT+HcWInGaxcmZeMp9XenaFe7CjeF7gZqFzWetquNNVS2Xx
leRHhKB3HDEoDBLUZcu+KttGWf/fPx5iD/kT7L3YLwZQPmYhY+Pbcd3rWulTYIMx
YdIY8C5/kOe+VpL2X9UXfmd53o/iq0d2GR3H3tzHu2whT4yH//HYbctv0Vr71Itu
OuJWheRicPSaR60SzzC8Hxejfi2M9izH+OX7bxJJJazOeKn3rHqDueaf3e/z4LX5
YlB1/v3GtYZ/LhKBi/i0WbmKuEO0jtePPSrEZLH3QmcibatP/M5l61y9EWjA7NqH
xynC+WJDKu0etO25MIZZJYZqSZ9aWF3WXOMfr1cR5ph8He4y/IygFWWiAzOnUD8a
Cx4A9L8ZNYSR/+2kq7hAHYkfql3N+35ammjwHf6gbeWGE5V9x2LiWdD1tSZZq/Qn
pOJNerHy9t2x9r1lgVQ5RIX3hlh1iQTSZqV4waaYIeuuHO3Gp5KpDMhdk+hnuvuh
6J+XxQcozVotXE+2AiQUrV8ku5HE11KqgJXg9+2W2e2YN3iOIhJF4a4fYYvXqTvi
kU1G4DYDiDBoFrKQq7aKQDXaBO4pXHR1cHJPuZhDev4Zxs8xaNrZvXyrwLz8xOWj
+u2la41m9LO0YCj7wOGVF/cRZNyUbWklQUIZXpVxQWBj83cUoA5WokMG60OQf7DH
BRHcUhfEhqjUNkS6QNPudfebFOvrdB9/tvKt9YQ/GCZX2Cu4Jsn7X80cJDU4LtaB
BMT9ZHwceLu4umSDHQosM/bmc8Iw+/ysX7Rl4IJLYVhURATpA98NExdvPrLWKGfE
PTaZfRsMkknrzc0+4p4gAiEWulT3WDMe/JhZbfTYgN2R76EFNfyVRwkbmi1zdYYr
Yvcb1a/6fS0qH5XIHhNU5ZCKkKY0ErqIFIEzDA/mYJNoLQLTbsm1kotfJ0CtoRzT
6FXZR1UWt0kg1weBcMqRIlhmQcMKDHxZkClApvihmtL4eJOCdlY/qD7S1myifg26
zgXrzfsZSlTzGjoE799FzHzcGvusLJOztEgAdTgulQir1U5hhBpHZfKgBrQy6/th
ca+ziSTBEs0MrJYj67H/hL4eX6cqkoFvJIb8rOcG48HNPeSrrvMPaDAHJcAQbC8x
lLAXQTlX72THW7KaV6x1ZZ9AAfS5HYMHjxIQINxO79R+8SiBnS2sM+YAQKvUt1Yp
hlslq9mSH5j5BhrDEdsT/Dub9pYl9+yZZli0goLaLNSYw0kPONhya2sZyDr7e5gT
2v2+kWz5S8Cd5SWJ3fD3b9uAkDQDvrcK8rw0RmlLDyGllyq9iQPyhBhZ7lCXq11t
EkzMZ08mkXsfqSN4nYoJ3CZEZq6aW/iogaEn1hGvIbP6bxDQP5j67/sREJ+Uj/vH
xW0jdL6fxKEKrpVCiNVmHw/hyLWy0Bz1BVxl6WyKNW1UKo7raACbjGeK4xpU1ECh
tkSwQ519LJv2cIohvR1qbG4mJu1iSDkSzrbJwBKGrWo+tsx4UKX/nJIpHJidqzru
Hj+1VHmJ1AQ+/BBMDQ+6A6JyjUWNH8yByZ9zw/WyHt4p0gvf4dgiBv+GglHHY4WN
W4FLsCXpl+SpbpxOgEn54BRqPmWfN1NpU+9XLieU7cxZQrZWWHv+qvsg/wWp2YHi
sVs9Skf3/uTTuhvuGntN5FOPG+dN+uuZsq9mC+TicLx44O+XOekgmQwTpWGjBViG
9+nbT77EdMZIkS3qD/OwVfkhTXUapy7YaLELAExKIbRESyu2FNqsx941TCRun1F1
Cqee2zMm4jOaCqBSdZU4YTSZjQbej1vxl6WhFPzQ/GzMZ+J8YN1bNzgoSt0oDZFf
O7FdJ0B8aEiputivRuLUeQ43/81YNbGW+DK/wpLJm5M8I9jkKAF58qtWQgSLxuaj
rKKfHkBbawPR2NOKklVCM8TgNPeIoa93gaGmheY5wIu4u4if/IUCyKPc9nqVyJsR
aMl3KBZk0lA1natZWeNKgOjeQ9yOJED3hx9yj3iXvFJIiMqz67ypwvfrp6E2Si+t
FHgouowm0LgWyjO9OiAAnndtKzABeDp1jPnUbknYuwqMY5S1M7GiuzkGxyvxG5dm
Q3umnMEQKxZkTk7hxdwYFykNb67NxO3g313t9dWZVGO1xFLIdXjW9Nc1rFQZ0MHk
mroFPi7R8PkncCXXHHgWOywzWQe2H2kUIxFXH8UGFn+vjZVshlCuYT7pHmI3VuO6
OEirNAlZyEtbxwID2hGtV+XazokrHV/gTQsgdMygVJNnAPpJY4hIbUtpNHFR71w2
T89xUNxuklC7uA2XoVV4WHjdE/3mUJLvg+vDVhxBqgDVDHk6Jc0bX3l1MLIVaupX
JLYgUljJoNIdOEcvU4zf0+3Os0EFpzhiN7Mhcsky3M3FXKcKvFSXr76Gp4bRRRoh
/kXKOu7x/AndBwtO/qoj3eZxEa+G+REpSUP99yMKz5jNouPe6iDhn7sirZ6/SHpK
ICibIXUtkI1rL04oWeNxe8EJNphUgHGyjM/wGYE9xkZLBtix5JiZdXwA4ueFVqwS
93QGLsq+WdDtxrbzajoX7TdGyXcp4Rr7E/gyEE1yd2/6S4NlDdMzaYBfYVZVP1lU
9l1ze/8aoDVJi1wr+GJSsPMabgR4aVAg/kig3fHhpliFMh5zi74bqz8FxKJO/Lmy
4Evn0BDmOmhOp23mAr8Q9l4+07K5ci6Qdmdmj+0IU+mUvqwvD84xuLp/IndNx+f5
/pKUBV+x4gTj1QwCufkARa0zhw64o48QzuKQUQYLFItFkAGmgYohYg2Rl9l23Bcm
8vEdSJ4iah2MuJ3f3LaOUMAw1B4Y43IPlDBGjnqYW07fTRNIt5XJxj5T5nJE5pV4
ElVdii4rEHCaAuS5ptH1mcRzCBv+PcMAmqqIvPRH9A8/afVNpg5OUjtukD14/eNX
K30widfliN6qsnbefHw7zUCbDFlZUFtHA1AfYFyIQJCEKXWNrEmjdnCmuccLEYvo
WptYJ5+/DD9PKZF5rSvmUdKKfrI5N4/HRiZJgqhXBLpHYon4nbwnvmS2nxSdEkbS
2miZ6+73+OjH34MpbArTTQweXHBWYtIOTCrEieipjpBjUw+IoqUwwB5iEzwkZ0v8
O2U4eHgpBq4TEW56UV3D71Qqef5w+hrEhaoSLmfoSISSSBuKpalGnak3pJcUmShZ
tYjv0shGNJJFKCgqYnK05Z6R93fEWySv86Y6FRCNx626PCNiF4Zr/lPPEo70jANn
NvAkzUlMTWZhSDTBMJHOgZG1HOxHJLXc3WXyleZd+zjKRYBG1T8Q7OJZzUDg1dXE
JqW6tmdQGrVAxp24fWOkcjFKuDquO6h5eYWGVznfpMNVdD+XPYijMwL1LxdxMW9E
l8i6PtO5/KCBkoEXRRw4ENkcMpHSrecMkYL2ofWKtn0QiyEHiJ138BsEo3+3btxW
H6Yv3iwxjF3W5unuCBJyOYUfHql2i7ammm2Zc64nK4YSnR8gqOfRPiJzlAZdHCli
mfEM25SliPyDvwmtw/eShmL/V2gWJHfU1fGDNjIqk5Hd9MbURL327uVpBtl0BZo8
Oyl1RvGlzJhLexkVe24QsSLOG5swd3Sjsgjwzk1CIAOba52lXnhGM/meIggrsJIp
mL7yETetFJL0Wk/5N+TA5g007UxzwpkU6zafeNQpUqiJEqjPbXP/TtbFETpPlouQ
NpusozBCdIRr7Nx+Oig3+StmE1da7gcAo/96RmT60vQH3rtiqDKzWBJp0ILMlEcY
gzvT9MHv6aNInS5rgt6+Xs9fUGxMSAhV5PSzTGsAwbGi+UHjAb6DOrl6GoDkf/Yf
AH02JL60EaAfVDipvrVKIDW5qyY+UwJ3I22bGuJdW3i5iZ0Q1m+OS6uBozO6D63p
OuEDk/m3nXyHOkTQojuT1mjFn2yQlf4AP3E9/s0kT9SVpHSpMD12KVWKTio0s5Es
RUtmlOVcwqICoTMUEL2BbIFoONC9/W13y54+93caeQZ5sa89mA3g9zujnOr9OW6N
p8FayisUm+qO5rQN5Nizfn0HLd8PmmKdJQb5XXSHii0p/whWjVOi+r+ubYlu+akJ
Z07+Vxf4WXFUM5A+GBoPTN+Qz4Nupag9TGGoGQlVbTf8En5SjC6E3NYEwBB/76Ul
dD21MI9dZKqBVo05b2B8Y5pBPU9wBNvumiLh8Vc61N3YVHilw8Iai7E637+0CA4Z
u0pcwZvruoXlm9B6TUmyQHIJGp47knEpN9sOCCNgB/7wovSjPNdJ8MCQRZL3u4z6
Adi+naKlxTl93jjTFVeS9A6Lr3Ap/0XS7To3BxhTQxoq3sLbdDxfeWGOv2eG7Ksc
mes82vGCx3eXv+4Jd5WX+nA6j8+BknFwB3++gMj4LGmRjv/D76arBTWQnGkUWAfl
Uoo5BwjgVeCI/dLGn1ikWcYVECMI6aJOmV0Hu7SjYHyMFJUPMmxrRzvNcJmwljT5
3tuPdE0Dc4s3zYCg2/ou9iE8HxF8QwZRAwhgL7zRevgoT4rdSIpH0Ias5JMUDFrA
cYiLRJHiE53Kta2oaRZqvDx4dbAYWUhSjEYPQMAVhbslht2sRsTMAYKidTa2yYUy
aGQgtGBNh7sSn+csY1H+PbZaVYvwBVZxwGfnn2Nox8GBlD+Qe+xykdyB+TPvh9kl
tcnRBXfGYiyq31RVdf13LvGmPWD6jWdJV6A2Q2cbpG4oq9RneKUxq88vJhL5XGvM
bjMR36zOam+EfM9uVqdaGLEyQCwAJ9bftbTf6uI3SL95K7opC0Xnc+zAWSB5mvsa
fUwplmsC2NrjLpyB/oWTX1j3FdgUA/wlOWeHB+k0sbiKDNVTDjY+UA5nbgh0pNsv
/B4grwQCFkIUWd2S6PECk2tGkOpHcrE7O1dvSHQvPZimJDJCcqKwBjlulrgor/vZ
mF9EnGs4bBAHAJaCuOffjuCOAxVZ3d1+k2BZlQF2MMBttWSIufA9wj6FAs3Fwauo
yHSj9+F/mGuaZhjPzsWyBXHgfRxgZRsKGy869SzA4b0BsjCIAgD+BCV4Vl9s91zh
r/EMmeINXRyZFdeSaogmk9lUxaJhBjTeCHUDS5AswM6tvNWFuZ0F3+hnZzCj/3wh
kQWsywCH7ioQrXcW0uJ+DJmJmfr8XSX7BF/EWWxPfyMfuxSUFsRaydsHkmPHSmnY
x1FOC9LiQnB4G5RjvHEdW10cJhkQbBTl9ZqzKe+Q0eHTUmCZ4xvjP3R/XHLFwQFw
VtI5m0CB1d+8o0T6dxyHc06JTLT4gYGjg0dGTWjGZvG7wAt7zh7aaI+h6LEAWFek
KcSVWuioNjMhQ4g5deXwPXkwgsyLZ0800Jqw/mDkkJvBUhSHpflMXGsd5JqQVKrc
0t92Le2HlDQXlr/wi+vZeVsYkZd83S87Fv8zNp85OsnPM3BEOpi+n8osSPiVsM23
hW/0ovlHfL70+D/K4+ppH4GabWGy6WtWiZErJiv+ELSz98X2yIO9iQ6mGzvEs3cY
J1uerbdSqJJSLEtbNvY9pzIOH/Buwx+VWqFvKa0e/0R8NGU7bZ7e8vYdfeqfdMFr
6xnC+SZF7Ih6qGmX0YNQz2ChGLbjgeJ2BtNuV1m9lno/moxPklqTFjE7LPM+iVNw
jom8bT3ycYIM8wwI/51KHn6v45C1O3zKpJBLpTM63VNQXeFvZ/sdOn31UW9AXosq
fa62vQQ/1+Ma8hS5NntYKyBL3kL5aPJT6yMkM4A9ha1M38mE0/20ZjB+0q1dVTpR
AbJ/OQdOXQGupoAqUicWvwe1y/pTw44irDmhX/78Cqi8PwLdMm7eV76avEy4htAq
Kq20HnnDCj4jrkHcYmc920AOuXasbF9xqErqTHikj5nvSVxMCGHdNuzH+YbkHp8M
lunF9GkpUEUzrFmUV+FujLtlBpOsn2l+iO97ZiiMgzAtlEo4HbsPcMGsTveF6XI1
VRJgoUKkLsijPmNiF0lknPVUazBtWqdvK1t3NHFYz14ZvtxDzqSnvBlGhnEX+7/x
U3qZkRPSq0B10wCFHS3XOIsOvI3eA6Dn0S8/JSl4qfeHibObExtFvGunYg2jphUd
Dq054kna05uuEkq3EnIxGXtvc4mi4wHjD+MsKO49kkeGhxi/pBoyQaAde36dX566
gAbw9eHmjFE7ltFMT8cjP3Ca3Cj1baHeAfAwA73GaQ/JR/eNRo8xVk7as2IljAQ7
7pWG/8ySdTIUno1MMB2PXaKKczZ5kDGExr7zCFwWkjLvsTv0g9CvW0db39S4g/wT
fl4fiyd2c/vhaPdpP2TMX83n2siPi3OddATDuZ0LxlrSN55eMP+zR38HS3CGf6/O
dYaNcW7YtLxsEQ6GeDcsyNpthH9MRnGIB9VAqZNWCWBgomn3btRs/aw9d2xdqBnX
DJS09C0DkoSoUyegYIJl7GmdRQ9gJl19b+at66qPHY6UxmXRMvSBOnKOketfBH5s
obKruPmNi73VG5O0zfxv4b6Jfs0PVy+OvKL9VlMVys52Q3A31ERSEEyLGA7VQFcr
XYFhw1WcZuN39nt+/2fGD9SaZv7rK8ix6bZ6NGVSoYEGJdo6hAq8aVyfm1Hc9DRM
vDzG70TxaSbhEmLp1Rys+mDV1XFFTTSw+PPmtAuDPUCdk1EtQye0zMfsZmCEYK16
DhBo0dI1rxzQNo+ib0oguH5wT+bwLDkt0GgrO5u4ID/d/Gcr04QwpOdN5wXEIUvY
ihgMXn+Ta1cuBn+98to03MouFHaPV8+T9lScaaNe9/Y2omJ+0OmSGRcIi3+hyglc
UDCWqOU+slvQWH2cpPnCG5qLXcxkEaIdun7qAMaRBP0qb+ytUBiS5MgmOuGVDm5L
tN953inX44Ot/e/7MmXGrQx5Y6g3orf/e9Rnm7T1Xga9jeXuw4mim4S5ktcBbh/u
2nuFEERxCZUNRA7hZlSfEFPqQQpgdSiW/8NZDe1/DN6XWAl69lBJ6ngTTRASltSg
BBEZweNilnI4JTEzVhW8XIdHWR5Kp/WblYRrmj/HCCXM9uMoNzZBugQPX9Tb2jOq
Ug8nywzlUkJZTIup4LRl0ZFk1VdG3csnwwYzx4GCzKLokywK69giqNT2IJ4QLEjj
8PBXmNReRToBEvR8IGhglk9A0Iw6w56KZM3sL3hmwuBv8C9KWP8j0Sf3zymt6d5b
SBwiFCtoNOOFpYYSCn+4PsQsIcR5XOAlilFDPF9akpXjtL8FJvuM5QYHrQo/F9NN
hsw00GbYoIGGP5QEcIvHHWNz81N2fIgAVtFQJDLN2J2dMP3SUmKdtZTL2dN3tOOb
z3VzuOfNPUCKGMH3R3L2BeF8dO0B1GzRcOl79zgRkeOzF6Y3MhS8GvY7wuxzUAe9
+mGAFC+easHDEvmhQLRnKKQzt+1gjcDFjOhj3dv/VrjlmKuenIOlQKTUAz+peoh4
C/sFWGHbw88r9DvNjGwzTRmL7bAnX1ACiDyFwRfiHMG9HXKVSEUddFtSDFAaKikU
vXoE20WfbcoXaG/+SeKWoiW6dQPRz+jG35I3gHSf4kUJLKxYoO/w9Cng6pGxBhv+
tPGn5fsmF3Mn+Ld6vQI4g8GLig6qjUI2Z78ejnjqDIiySEkkDu+k0pCXZ2JhY/mu
SR94AAh9y79FtU6lGwIlcF+0oNXkGOeoWND4eSaHqypMihwLHOXrgBXwkocWjs7T
/mpKHjtWX4GM9l6SMB+ZDsY/HSsPXJD1AAP3P/fdat3ZSlCiAs6VeEBSRhO79T7s
Tg1sEyu4TPtkmaglEdqZ5RKMzitgCYZ0pyo7PbQSfbqd/+cTf5fPsgBuktbNNOxQ
EeCzwCs1Ebjn020/DhxmJozP+aeu2FR0bXY1rsIGe3h/v4YNJJBPrvmAvp/Cubox
9fwuCEK76aaG5MuOoNe9RWpLWwotbMZZNfbiAK9WCyLgz8H9LK2uA0VMZ0prnR7/
MoaJrTMVUeZ5vRXR/8u26zW/jtpT5ATdAIAgXgMH3JbFzYSvob02vMRbyC9+uXOb
a1OP2kHPcVqg3H689uPccWZtwQehX1csv1Udx0LAdGefoEt1jDd5yjBCCV3HHzsO
ET/hwRdv/Lrnmgr1A2KNZEqpDy7WYYRykaph41zQZ1wFeOHQpx5ixpPLLpxKvzbp
Y6WfsybnbOe/L2uB3moxxnOZk4juUpGK1dtTqLDg9OkXXT2XgA54/xwOw4m3F+Cj
mRhh+sLbVqkmg+xiulK7gZxuREQoMmIEQFgfzouqiA/+mJGA/9b96nesi43yD6Oe
MOLduLZQp24OMWYdA5u9Usn012rsO3uWNkLyBkvd/3b9aa+56WbfcrRrNnTDG2ts
RBut0OR+QVs65VIPFM7ST6lqh9hYls538wCwioa3tdKIe8q1NTRK7+cNQsueUmis
wn6eh3M74xdwE+7rlpKFRFVvdmdwSB6zbwLCWGCyldCOX4ujau9fo+Ua63ihrv7k
+uEQihU2XUELSaV1H+anXmJeuOmuOX1z5WpzXtXW41ABdz/BwTzdoMSNhs6eDuhf
suh5Zo4CdgSf6zHtyMHGrbDQH0XCcfq7c3tGwo68blCZvvkf7dTjfVLIVkIakVLL
x0yLFDqIboAOc7Nl8i+QRl26kLHd80RSx1zFgZiK/q5Xq5lEOXb3bTha8fYYznk/
Zgi97A+wq+RyxlA3h77y5KqaAW4t0DmI7TKONYr076b3kVFYwGd394j7Uv4AAaql
uz7+LQfv2zb6gsHhQyBWQL2JL1oyQe396T0Z/Ay8m1Kq8vzeZ+kvMJaKX+PfzE7d
af8dzVSg1i2+uJrZneBlP1RhMwcwTCxnMlQdgz/dPVAlSWV6fL0wrA3+KIX/OreH
1joM7L2a7MDapvm8x73qq0K+u3kKP3DvnQEvsQhedktBFuOFUB6CosNqcdeUvrBy
lwXYgir7Be3LgRplqdH8SM7elgQi+0Ism4NuMlm1t4nwOOyir7q/SwQ8DfY0dJED
ojmnbUYEAUcOpzFBwnNE0LXS96wP8zQUo7aTZdl6TdxFX7ywXseeHWqXjkfjB5aF
qWIMA89XwpJfWQfIqAiMaGVscOV4jxd5lKUgJZBcA0mmfUGQGKR3T8y2uH4LyBKr
GShh6nABQxBpRWfA9JzmEdFqKngQspiIDJM++tQveL8Agm/bUN5n+WizJgCuoK7J
FQSO/kDCJW5KM6qs499IEoxGn46D7fcz7mqUidxiz2yLYaID0KvSdcvNoJPZJrvn
lWoF5ZlDqVoSy3IhpENcPKS/N5QQvoUYR/K4Igs7MKwNqILrYoSnY8Q6MjD9bms3
sOswRbhjYDqtUlZb7sXkOXUz125u27+blxzofYpW2GSoiuYPsCoLLd56RR7mcork
pblrUzmC6bHZofTjDhhCviL2JdQzHMAoP6jqIj26rCGPQ1hB1x32AhJFwKHxtLod
XP9jr90MT3034N5jsAmLVShXehvhARibMxOU/R84DehupmLYSDSCIIJ3N+zIEjPB
PpTxIK/0LkiwWZifzBCOC7MsOmzXhOQA50nQwaNQzl+FDw1kdWlTIvNTFXh6MlDW
7rd+7hPw3mIbPcuAFqrWI7wuqPYQVcrhuPuKp7ZCTP5lmPc40PN88wKHvp0T114n
/FkkXP5dFJLb81exbCGljy44CDosv2bB+CayZo3SKmPDIuKFFBzPRHea0V7SMDzq
v8uKhFH5Rrk4gb+/hVAszwAUjkcTOpjYxgwonqYPF94By/UoQH7VjACCE6u2QtHS
lE2ydLjIjEGfTsiaH4YT83eEfNcwbaHp5qbJP95RNt7JDUjrh1KuKmGDpbQPyjiY
BPGQoZbp2R26nU+OMKoFuENOMyJQOV5YZGATzkpwm8NpRkMV89SPqFtCyda4S+77
RjSVpjpJLLvxStFRCHvCtw63zK4bbUqIEVhcB9ofJnXSc/98n2h/SNSsZh0Fn5ts
US33zvB1miX8niYPvO1CufE6w23jC2yC76f6s7/6EdrsdakCZxb4x4qb6yhE5Mbq
rDbOVw06CGXmg3L5LFyfWjme3vFXiFM1y1Q7ZeL0MFEKEFhfudrh7Q6j0K+PX1LS
+WZbIwlJ9PXsowphDR0lDzv13+hK8Tj3CJVBtb4wWUFcdcYfLEKIKFuA0ulPzHBQ
iqs6QIZJoO15+U3abBb1YTwd4038V6KE/3OcbOTVwGOKmfmWWLWQiGhFNumgLNsA
Rk7GzpLvz5l5Tw6aLzFPBCA0xRovwVcE2kaxXduCLxuSIOqf5b6GJUWHURGiMVpd
3St3qcXJ6Rqv5uInOnp5qmLbyrwyWPtrpU/iSscXh23v85umL0UvEk/2pYiDW8s5
USMexN+7vgrkXF2rUT9XnK2u6nDH8eEBBFomdZ/uzcIQspNiHW0yeALZ9yuulTZa
/3D9nfFvcknpZ0ZbmceOkf0matN7Qb1BAJn4CaMtFGaBsn9dp/npvfj2cv3eap/i
LUZVlDMV3IeJJ9nKxkDuRKjrpO2m62IyyILWqNan2zIKL/VvKIme2KOJiNemGhND
F/+V9eGmCPX64QypEyQRFG7Hcy7iAU2LmqigC4YV/ObjSW7viig75H5J+ENBd213
oelDr0cVeCPsTiSi5me+0t/eK6NnF172QhLFoZr7EJHuOb9jCIIujmLvbb4Fbx3D
vj/vkrcC+RiDwT0YgFB+3kArlpZQ3UeBhlxTwDg7+PAr73ompe3wqtJugzSaWARV
Site8wCzGhRChxMXfYrYNHk/eB/Q3UUeIpuV+tWX1Dq+9KP+NDYnlvlK6S+R2Fl9
1TqRiLLtOXrFzdDDFTY0CWKwBVt0RhGqQJmk5lz16vQ0u3fZImnN4s9EW9fum7FK
lN/T2CS0YM0SFH90B+YYw0U4VWzdvPL/z6OGiMSulDPS3j7NzF/gz/rAj1H8uSXI
qf6mlGknlLIF7tuoKxUfPKTHQPzHAsugrc6aw9xWpJZ5dQNtBngNZxADJnT+0OoC
VhfG+ATx5J9KXk3r6ix2v/0hoWo9ifmnTmf2QvtnVW3gy8OyelmwoJ8lJchMUWSD
ifuJIkmqKNRwO1p6SW9BjfqOoDzD+iN24ID0JmMeg/ZRfNQcjsBhoEs9ONm40/z6
jYIHYhLONRcGCP6PLa7RU+UHDlZkVY577zxfgq36nfFWpuGjt3TBJWniqMH1Red/
cBa3joP9HMTLg8wQwyLJ18nxceYvJBj43t+jQwiB3vS79Tt00RcS0QaH6d7mMmP2
qrtdX+AcujZq65rFlSakS2/YrRzsvX/VdpClc81wF0ncN5iK7f5Ulx8WZcqZANnk
S446oDFMdnjaEwEyDEHKjYDW0ixLznpluCiRoFGPlN0F43UoyP2beuzHb8fWxYvl
7WoUoAuykqFyQhUG/Z7UvrMj8CI55varxbLvgOCueHKiKgd/75YFGLVVgtJHMv6I
HQKter4R0ADcuAWHP85JX9B93P9vOtiMHhs3ayH1zyS4Ahy39VYhEgkDB2Mvblla
EcZZsYfa75zIW9HRS183ILHmyasS1aLRYWnHd2yw5NVVK9oshBQ4hR59xHZKj+bk
B2U/EJnE2isjVcwMnyIYFJclwGTC09WER59S/fi+wIiqXUQmdJns7H2DJZaBfakW
fQCb4WXH8rzRr3GdQGJlobMSmtig1WJDo9ff3ht8Aw+6xyoVc6VR7RgVwklbB/e4
lCljUD39stnlacU/T7L1gZ1HY8kMIUZ0Fy0AmdmDEhvhpKFZ060o3H1wHVrazOUL
VPvpdKApLGgGW23uceRwEjcsEduFuDlkd7y5FV/2BDFl8JeGeRSU9ur+3sQpi4RM
HlqSdh2Ag5fHpsMtkgYIbjaoG8ZzLaLieVGWnvLfiyeupWkCVut0Hg4cc5xHJ6si
bhfoNrHoykU4wH5fuom7mlPbu5pOjzwzZYOVPstSBjry6P4ftXG8p6GCJRRznBY8
bBuXECClbwtPjR2sOJ0XYlScHZp8gGOKfUv3ktsNIr86UVNWuVIXhuGDQzCez+47
zbtJfGExL1Sv6FnB81Q++ax6p7CIXeUOLw+jBbYezYrOEsF3R6ArEtzJ23exmi48
IMUd00Td4aZzUkk9T3kqDxIjUVohovPDk8hy7HDCpI8gNCvoBaJcjPSa6J07rJ9B
U/C0RNIE+GyT8TtfO5xTLYqptN5SCYlun0oggSYwP33cTh2Fa22VLO1BzsZXcwFy
09fd5zCoesnEjVnU+c63heKIgSGScwF55KjQFXg3gqlw0Xn1ykEs/NwJty/jHCiM
ugO8k6qp6Rxf40+k4o9gef43SLm0k2vF+7Hpp+lmQOV5MzRvYEILPE7Sbfwme9Zl
TQOSb0uvpRUCq6+2KYDni37zS9DvhdWIdFuEmhxeZD5B3OmfCgFRgTroOXRZ9lOu
EJlLn1Qz080gNd6UbrC9dzS/zmr9iJ67LSCIfRVNFSlvnOVRty+wbEIEgV4U80SO
pQ8PI3bjZdQ9u4okeFHAPDJB1CasfDWS+ek4BmhsOybx+qHcxJhHsy20c4wib7H0
2P2+t9Xbr9uSA8nQIf+Xx+EXXhDP2aZ6Kln2xcffZpLUuXh7aByN2joG3h4htRqW
mhMEo3jImDHAjaFgNgAFZUpxzEMGziN4hKf3lzbCy7yn1vDOz1kb9niukdnYLLbI
FtI7CdSi0gKdRnfSK6EvVLUOaweXGD6gYRtVom/GK0Wq8plr4GSvAIyMqmNYbrq1
UnFa4j3X1cmIAFSJ1tcG0I2yjT9lWxmbzQKoZiqkpTAqyTNFQXstc+qXPyUwypRi
v+EXymxcWEUPk7y7i0vn27s9jGTMaRjwIWjvNr0NRHSS/CA79a7ot2wSbinQra4L
/OE5CZBMF7PSOvzR/LoQLhWMjamrkcCbW/+OBn6DBkRI5a0aafqi1+LHXQDsSmPx
Dwjkkgq0HUH7hQkv59lQPbY+naeEgux3X0RM1o0aqJdSWXwSgAyWHSZFYVL6kJNb
YdL8i6DQbKVtIytKzM/IV6pkwV29LOOrvwGVupHpHu737qj5d+LZrmLsrH1rIOPT
X+HnGE7jPrXRWcpPLYy6PWG8zNplBBfnxhpUIFcs+8rwvksVrKH5zQl4NuuQr9Wp
hdRU4lzxGGVhJAfVZBHftJ6aNdswlyqsOxpy+DMNzodgOnctpHBxh0ZzXSELaD0H
phBUk0mXx3iVXB7DQeQQMcmn3CvJ4ja7Rju0ol3bQMjW5DAnwEdZH2duS7Zkm4Wj
YlGRubfK1xaZZ0JREdMz6KGNrNE0sb//X1S91ym3Ox56uvEK/U9Ljfncg3stmxmy
995rp3jnBnQkGUtc7HuYnh2qV7XLcn13RBDLf/D3W9YXd9A5ELyyZxIGmkLpcbAj
/bzRRAkxgMtVQptQy1qfEs6985lhbcupsZqk7L00BNiJC+/ZLe6b+bj0iH71utHc
s95Y9kEILvf5UqqtGISUK7wWlgucXw8xutePVC48qC+BdQhMsi3lUKrTyGKD/S8A
m1nKc4Od5j3IFyUMhcPsQsYrnZB8FEDKdN8SRdZsH3tB8l4jHpP3HIAUbHkX/3V9
CvaT/Od6C4PV39+W0qFYkHkHMrJUjtioDY5WVeOyHsPL9qS9G4lApn58YVYEc8iC
wzNKbTmNzfb+c2dLshNhGmD4ej2GtS6JDhi8lUsgSW/fhnf0zmG9XyWmfbH+H53N
2DlxpbyyzjU7omWSa/xZlKZLkbFE5PGB7r4j8s07jkGRKZr5xFy8sajvwyki7uSf
irzNxUBl+hvnS6zxrvolGJmymbUBtD2kiucW4/O7Clq5GsL3S8DrCSCfE5z6Aodm
IYU6WMGPFU/P+m0hNz/7QY3iPtq9LI0kUxoPgctf+4mUovqZGJYyZQcCLw6IbvEb
vCp6xyJh9BTSqwwGbiOz0UQsEGAtz0bbnuhy1l9qLnLSBUVAOtCDxa9YTwCw2FCh
3Hp9dFvFOeTESayoYW7sMKiVkdHdWIszaelBilUBUQYuiJREdGts8+oiecR0ftR5
pbgDKjuO2w6Eu4cGkCyLADyeR5qrMT60XXYZhifbntK5P2qDyGaJvxOSJ+Op8V9U
YQbnP/JUMzIeWFxXUzDgZliEu8vKsfmXucXT5J0zatUBDxLzOqDLQyr9ZOQi85Lm
GiWFmR3sK50zw/pSE7y5ehjb+L7subX7TMDjSz1h4g2Sn2x57P8zl20JLLdGfRLF
g4OMulO+CMpgTQI6Zi/e3qdv5XT7GBIieWVwkAiylTjB9jnsvPtRA9b/65EXea7R
xxMyvr59E63v7b0RoZrWakmy9rn2GMgJdH975Q1FAeAHgctv580ya6WBdtKSrzQQ
Nkti/jTXdDEPamUeAjWRTuQqqwAtTN0IL12Q0groZIVmLvMcV43IDqp5sDK/a5cR
mk+x0pcg6mMCtJgqEjKbB4sweG1BKXvPIjf6ktnqjbXfnv8hurnPKhUS2c7SZlG+
49KuBC78ok4865hiDLwt9OeQ8lG5C39OEVLTxtuyZxhQXJvwpr019uMS3qA+Hj0s
xzkhajSTNK6KsH1Ao/+bnHVfAU0t6p14foqrdClurW5272du7h5DQV8JwIJgNs7/
UXnDb4SV6PcvGM2us5PLl3Vt9xy0l3xSoZ66qPamxtrcyqbUARUUeHD3yms9g8Ae
4enBD+X2NejnFCTdttiSe6Iy8GislUGIbpxEKJkjv6Ee6wMV7zkY5zzvuylAPjvw
cokfXPeSv8BzeUPm5lg4z/68hjyuLYx6K5vHvuRSDbwXvszZuCK4ZkfpE12jd0s+
a/Ua46F0hXxTFkNua2xHapkz23p8xcPPUIKHb5MAnDNtrmC+rkxX7Io6KZWTO0/0
sDW+yAVbSJcpTycV1TFAsJFklB8AcnlpbBh9LvABU9CKdEVryan59ugvMRrf6cKD
MzdoywFkyawCg2OsKNA7nsoTywpym26ZIhsBSP1B2OhXo17E5GPBpQuX4+i7nTG8
soGP2VUN1PRo/sbIU4xi1hz8276F2IRSa/DhvFiiQwj509NEkLv7NUlLWrtbzmcq
EzlVDDhW3NOaujTozFn+WLO47jVdAkdIRQ0YmSqSRflErTodbtZFCisGcUylSQnx
Jv5revCThhR6xGratU4Qrp0CZS2nq8pdRrmfwC3pFTeSTys4/ceKFJlqM4OxX9Fy
BI1hG1CII0u0qgdsVFdmRwu/Kdd21fu+Lh79MrBHkYlwRSbNltnUW2EcvBQxxAp7
Ey3uiKQXhTrkiRfVMLM+d4HUyd9tA2HzWH8mkInEUr0EFgsQCNVD0rnsyOiQFguC
6ce0+mvHrI3cY7zovq3zHZuPXN/AQEOgJZ7mDGAnwkvB5Tyi2t0yjuJwdzj20N3J
li2IrlW2hd8l83e6RISGFD1d1DiOrvTmpEen5BN5TP7ZdX2x/RrKAioGribOsUr5
9jq7yKb48DtqmWM1lSi1TfaU7bQhGPWOs4n1uZb/ixtSMX2Cvmp+dCYgIMRjUoql
PqxTdRQFiFhNKQW1NJFEGsKTH+verj9SV7YhDb4qtYo/pzwkTcbhcyGzzP/68nLc
QzK5Bkk5qMnZEY5YcHsockn9fQBVFELjSe67N1m0wDpJkAwY5hTC4ZH+/TSWKioF
tAd4MoRdVt4tiSe845LnM1rUQgE54v8Z5SyzR7YkX9QyMRN0E9/bTLe7Lb/aJTCb
cHuJRmjNqDCuS3CDdk3vh5d/2q9mlso8mH81rV69Ox3xlOrLzMMuPpFQ4n8WFBfp
+T43fn+fpH4PfheEGbrgrNVQv65UVRU6u16/ULLeIRmT2pI1k+FB5JEgi/rkizXp
6qWIYQYyTaUkwC3Bhttd9hHcpKNi/28ZbK6sh9f/czeyxLK+Y5rqDpT3sDLkqlUx
GLmmCK5DbP5ip7Wgz8iaU7kAtahZW9XgvUi+N+vDuFSrH15uUljyje8hA1/U53xN
HiRBu+PVU41oQhcH4C18uilRJQr0MT0WEiLXSZtDqQAzgM+RZUWQGz56d8doIGcl
1ZZuHdY+/5w79tVWjo2/iQG2IeSJuXFEenuhTlmnGZyJTnh0nda7QHasFZFOuTNx
cPglVpooaeqebKQTsQANmhDnnuaggVGxuoxaWJM6s3qvBB8UyOg0pODtCiHpRKNK
0Xcq6NZiVGMD/dQme8wgPVkC/jeQJJn/eE81cpdbY4Zr3GZn9w38FAHnMmy5Xe2G
e4hRsAODMVRxXNGawI+eGrPE/fGTLxdounYCxs2H4ZNMOp1/YRg3gqeRA4c4fASL
htEqzY+B88R4MLrieI1UUVE+UGTDwBaX9y6DgGLEpumLYi46sriVFwr+5VjphVBO
d9aMrP+tgAXuh4EcqonSDprLYKBeuNUASJyKuYQrt72FVZvj7ugq4WW5OutyMgw4
rH/XzRrY36dIzl/ult110LSLmQpgRkI2lYVF5357r2SOewgb1XgaYjL3PVtx3Mkh
K0uyLPLS9EE871bfO3UEyaxnUDReWj7KFc7cNvjwK6kg2gm8nvcRo88r2tfjh2qS
A/XqjGfCWAq0RTv/hiOL5yAIu/QRcbNr9Rcbd0gCu5KY2wYUYrT0Dv472S4fzzqc
MoOSCs7mmPS0AA7zA09oZi7LJT6wKTX9xSw+u05Ysgh3Gtkcw4qxkDdcXEN/EDQa
ZgSmXNoRH/jeTndeH8ZdTgBaH25mPTj9l7/5RkodzcBYGmwJG9+9l+nEcuNo/VHz
wFUVSdNZyJWwIOfrN9i2vh1bYo9kGZprKVx19EDl9Z4FGTBnU0SyIZA0jkVG/w8X
JcuRmXLoqYgJJrtyo40m/vd4bXd/WeMkSCZUCV+zOlzS9vNEuRvjjFRZMArpuzlO
SI/i/TQ7Ttu7sRb/uEVEpUPU+KFoPE3Kk8tNA25z2JrDoqTEVTqHxNrDkrsVqbVA
Qj9tJvtrJKhKHEThZQJ+m397jAUuW6tE8eUTgUc3Lrqvh5A9cSgEZ1L0vGlvS5Ws
cFSMP4ovwDVRURRnTJn3SSd3MDVrnlLS/RlIuDg6KHqZLMexm3dASY0pMgR5iFr2
gETxEn1diEcKruAG2+OwgbGp/qkx2RxRZLQgwn/Y9+Sj8997EES0f13MCJe0C0zj
FqCiEXTbcVBxaVFnOosqg1JicQCg+eKctBz4S9b50lxQK45W5uwCGhkh/g3Brvbd
XsEEYK9hfeRjbNbLcZRUumuKAnxBIS+BhavgxQQg162NrnttIYNoI7PW7u/hMfJt
XshH9El1l763w2bYzvUsv5pG4ae99v4IzbXZhkpyBSwCol/tqzuFbhqta4u+ofIy
pGJnACn/MV65FJdES98s4wCoxr6QAwa5d2JEA7u1qjLCVzvoMKrEYhQ31MFDm6WO
/s3wkGl558dKSP4avJH623Sx2XAt9qUk/FEJjInfxSdguHvGAkromj6lptXM+nn+
LEKpwx8lTql4VlaXUL7LSbHmF8Jueidm7usEBpMKDykrFqJFhm1U3zz6Ecrh2Bj5
fI9/OhGjrp9nB1C45Jo5Ra5TE+QESG7u0VveqJMFSki/atINSNSSDq5XU2H0YTS8
DPEEILcE0OYVmuXD5ufNRxa/1EFvfy+HrpClfJyJDihc3W95a/QVWJNj8yhfTHwO
qWov4albVOEyybfgZOmoRnRxBvdqr74pUCX+JUvZPBZvdGxNE5CrRH+9TT8JftvH
cTp1UaWxCzXoK/ZwBeXUD5KyHbA8PuTqPYgUTqNFI9W9wzHL3oM6T+FXfJVzc2Pe
xyqyloQACCUPiXOYY8RNiW3uZFaXmdd8Dd9W9Xt4lYbgeFygOim/ORK5l5nW87YW
6kryhDif7mG6uqoAxgjF8YylUrp8DK2TIm2Lf1ZjZNfkJFxIhHFrpPA0g0IJM7DV
wv8R600FbxijUVreyz0Z709bTrVDRN0PETccgPZ3ZgrRdnorrMtPwnTUHT1o0atw
PDg2HIIHxEdruGgKucPS0fYw+8CH3WjzgxEXlU0HYNwrnQxFO7JRD+gtkdD15QZ8
/7938qbyXmTb90IqI95Y//bCCRgljfNhpySav0kO44ZO1rPQVkuqrfRmUschLmhk
XvVXEkdUKvBX5DOLap4qDYIwHafzOf3XQfvw6d0g9KoObkx3qJPgezoaNiEV/0bI
he+IF34lhr3DmWJmsDA4tiovfpeGw17U5PrHavlHiYjZtSqDKUeTQ+cM35MKlj5S
OHsauoULj0Gghk4c1HI79cr/9OpYthjhcNahrCbO2Opsja71Q/dBvZ0BUEqTRNnd
lfT/1O5/vvDe49h2IVMgSyCdYXmbToes65wXazKv82QfaNr0BSOcVL/RSvYVNUiN
qlx6dgn6Oi6eScvPeg1At05Z7HvhKIhjjWSVyHnm6lk1OXMuN3c+fr5mKpmbbNb7
0ZCrdDj98zMEwpcdN2we60t2GvywJK6+QlmStJN2xoqDiHOZ+weRfACPhR/+QeKD
NUx6AOQK3MSjU1Ph6svq+fZNaV1X2jpZ1KEs91t1x+qgaNOwUdMFjZoa/622xL9U
MSc3/Gg0s6ERKZH42iK/x9TGC/ZpvQAYbENe+ihuJJ0mIB6V47cigkkPuwzqwGNI
rEeaEW9z9Yq8+WjqHicIt1CB3T0oSJGpzkk67q1wbSesgeAOyezayeWJoUck/12H
SDIcDJvV0ha+YaUW53JoSJ8qwuL2FTwJC+y3gx9VDeeXQ3i0xJ17mgMHtlzFNUaV
8VO4iZhaEjUoB6R9jmGdpLWOcRNI7Qdt6jc+ObSQnrF6gbLcsUtrJhm2YBmshWL3
mJkYMJrFyQDI2PiN9s8q3Ad4BXPFEE24Z4pwzQi3W9NFtG77ihlc2JW5eWHCitOg
mHi0zuB0VqwNHbFPYNepAuCtjHYMesgSH47NVpsNOqC4ehCVh9bzxOYBbgOVpnr3
43MsRIRO3OdIariuhjrTsmoCUgcZuPbzsauHp1io3uBLCmc15QkUcbZXdqS0DCqB
QUiy77OVlTifXGP27c9+GDDZZUYl3N92ncmLImlljxHfequWwFIngrtjAdpIVPaY
MdkY7FGQ4NHifRGLdE2LuTci3YlFplt6IHhY88w3soxsCzjKGLAu1OYJntsK2fsj
v8Ri/p37q4oA/J79L18X4GmV3BHTeqKnf+HZqTDytbWmEUcAi1iF60qeERmJxBdC
VGGcEaNnbNCxY7oIHALRsnLsEHA6qis1TbsSFNHnhCGiQuEPmeUtwt6Xvo1iM9on
MZBphBRLOiUnjtf+SkeBoPcedsdqaY8iM4t/bnqmKGT6kWnJNryR8ZBjv4+2HupW
nS0+MwlhSw5lkjRbX7uT5/LlLp4nrclJYJE38dq5D+Wzbao0+IIUHPRXGqaA5r2v
V6bIPFBTlxEKg3jbR7WSVbpe7UfAGo1pAHkrjTArDG88reblhzh+D6F5IZNMQ4Nt
DNM+JR4D5rCBW+4XyI87AXGHLXJEvfwqkw1/WFs9T0eGL3WuJ7B/ULtdhHe4o2f9
bouGVIIC1agTxOs3MzwRESa5x9Ro4UxSmXBebe4vVGtCeLFZKOHrF1VgE+4aL87E
CUBrySEbV9Mv9wtYCu1SMRCZMXqP4OKtLdhVfvx9ySckFcqnYzkyWmSUa5DBd3Rf
/FMtWgsZy+ma1bEyod7QDPR+5JlYBPXKO7tMn3wNFh+oQZFDMgFBbllK8ZdeI3Td
7fS+eeOSKdYs2MA6EMgI72qFl8QrtKhAtmA8wJ5orEgQMG/SQdN3SeajYbrS/CYm
mfGkJgwkTnNt3bSXbVkU136XC41SRmDjT+Gu/uTBA6VAEP/qBavTAq6KhduY3/S2
VXLeo27+Mg5VENTWuseTUNQp0ljzDa/yrAEiVVOifRYiQd1LDs84tlHroKoIRyeL
AStb6z5dyDho/rtSi7KQHH8SJwKDKjESgr6hDOjT2o26xwArRuRxYTFlKdz2gtd6
VjPfz1A6SlqPknirmv/3BWnox66SPj3WMpYwLX5x+RFWAsGp9dPa0FXa9rxnAcXz
eBpFoDjQ4Bqg9NaAFzjS6zD/R86ENy3FQ/rgFDF1filZ5GgxgAZlLf1aaxfi3O7u
02lhJ7ZkgAP3CHDMr6YgUVxObHunLcauyubgbgCpwkuopJ/NX1+yC2XCcVy7wW11
nx4RfIGczk0glVm8gFvwYsWizu0Ga10dwKtt/hb6Hxj2zmoUXHPHbl3bJfQA1Awe
hih5vQpTdZ4d+UJNTu3t8GiltfrAYLzqz9+jl/mmwuc+CtEnlOcFzzjzEy0Bay3a
1L+E/aKd3e7sQpJlaM5LmZvftQIDF+mFegQVw7LEda5Hp/aomPJCVP9EqbFAMxgo
JpUuD6D6JtEFMcamGmtZHRfthGqarimIpfwI0PHnDRvFyReCqu9X3OgRtldM4DGx
3oR9bMF89zw11klxBgIpiWggpdtDkvwMGay5P4KS6mXd99H2HxbOCod0uCxZtypf
HDz1vdGV9XSwWmsKIIuYrH3ZIFihlp9pRfMEivpWOqkjDmSe+NANjRkn5YRsiXEE
I27sZei4Ti88UFuNWmY15j4kVl923mltqao5BcggwNRJgt/KMVmSdkP/hR4xnLcG
4B66ToTf8Gh+mQ6t0wMzioE3mwo4SiCjhJL/V6QtLhZLP/a8VBVgxmhE/Y+v2aqt
bTRcR/Cj6UNeB8A3/iSIdcalG+YL8g3x/y/EvveC9q4eKZoHbiBuqkBTSvidbbl9
R0spKESUB2iH4zOc83BsXAOhmc1LhQDuMl6YuPwbWA3+jwvrwW/ZG0VcMU9UjwJV
2S456c9sRjGRuLmx9GysWiH1kRupITacRkw3qQplwT7NqLiMFL/OUbNOWI/tiEGZ
k/JkYpkp81T5jGNBdFw5t692L7+Xalpk8Sm23Yyxx01zcNtObY1XQC08AHKDUnss
OJ84yCWDfbAlRF5TAswCzBf4x7zc+Ko0zofvQQW37Um8019DQ2dz21jBL0BPsx/2
it3eVsaBzIJ3aa6l/ZFuTwna/rsc7Zjyv6dxeVTHhLQw5uaULQB+WWG0IjMVE1j+
r2+ykn8jc3ire+uqNaerPDwPxya8HH1zoyqyeD77g/sxEf8GhkQ8TPmHF70xiFDE
EjwWpXGslEnerya9OmpQEUgSXJWTB59voQxCKxWK6YWHPSVmMjTcbTSBkBIUMwoD
wucqRcc/Ej0lwqz1i/ZTAFMAYNQ+kOcl8eN8+RMPTgp0kQQnFXZoBBpApDpgPysk
q2IjI84Mi0Jdt6+JvwvpsS6DnmilaPzAObV1CLFUiYeTrWUBqI1wDaTKRiIXG9yQ
ZbCIqCVFXYG4iazntU+88tqyEfaTtwqbccmibqIY0/hVgQvIker/I/JH7MfvNpZu
ZOHEtYo4OX8FHufSvVtJMEQWpWXUxoo2C3JuKYPRXY1SEGSOFvnDj2LOFX1mBQft
hUpwPD9r6Q8A1qbNR87tu1Un78yNfchFaytQj5TStXS1O0470ELe4vkjDXLlstxm
hIr1RS7ExbjdqxXk7QPIsbC+07z+X5q1iba0kuWcN8LweAul6Wbv5Oj4URfRGk7E
Ekz4vTz474SYMoyHSclDP/YJFCBuKNcHwrvxSrKc9B6MusQwnNQYDSkzXdpEfS80
5xy481oCXKxemPbAHXCF951pDJBipbgapuXat0HTPCAxDBTCt/I2p4xI7zG2r8Nw
B3bQeJwfGb8eE21iatXk9Sgtt2XybqogzNyGGHB3JWkShT8SYvTSthOu5qjVZsOK
DO5JXXvG2+8yWqdMDQkJV443HShSRTfuSjUT9pRvgxMPWW2wooPl6u6betJ4J60n
5qiBMTy4O4PDxFMch1sCuulbw3dBHMdYIrMQH7d32Z1sfwZ5HfmawPwK0UTpSr6s
nvsQZJI3a8lK/hroY9lwZkKT1etLLmdGO+2ewFhCCzjUoAK+9kUCQiMGYm2YONdw
ygVVgu0FiZm4o7I77TwNqT5uwnwenneee3MnrP+N1dM/UFBgi8nEz79W0vzixIPs
KXbh3huXbCc7JbbCWfaAlL1dN1D200j+aPUBtQ3IqDU9thdrzJ2QjJ88IhgrmC2J
sP+oMB7H7DqKMOUXy45XNJFFb5iVh2WPRQXPRj5DGVdL1UVDhvwpNBgzB2FtK7Jz
mFeGYgPq0VQhLdM5r9/oGhxckiiLdD8LBVyLtyHoUrDioXDBHhhSJagudnQ6JuWP
iX7gbHrETlYmCct9QiXgWuihMH042NwYHFRPCv2vMrlXPO2A+sYvshFMAC4InGbC
BXRPABzEf9imoxeHyictxiqFKBh4xXq4KmDoSukvnZZoubeiHUWA5X98l4bhyFT6
oVsfWaDoTszX1DrwoDOmXKTbvwh8Mo0XBgRxNYqKlu62UxM2P90j8hyR+h4HfItE
BQgQgnCLsa9iOKkxjUhYb8WZ2XRqjTOtKgmrAiuesutGWOGRdFuxGVIXEbOBiYZ6
Y2wzSg7F69iTJDQRccMdcOq0VQpZXg13jXx4p1vj0E8gMXQVvOHBKANVuS6frC01
abkP8pKzbwX+XhGQEJtAqH44n5x4beTPUxxuJIehf7V7ZkPuVYd6iOPws63TKaGV
vhRNwI84l1JggeM7EKuokfEdgeuF6PAEHLQWo9tqT+noM8dd74qssE0kYfOn91bR
BnxD53/9aCSqNtMaur5Dns5WWiQT6hf3OVPQMjJn1eYwc2eLrwiyDdb/Y0qhYH7s
QWCftVay89OekrxGT+fO3uszh3U+IZuUCZ1VxcuMoRPyhgYxoPwcA9ANXTvZ01ns
2zufi0WKxvicdljSrPmWQXEE9qYR1j3kuOVjl/021I9Ht997YcfIN+ssUhWKYka8
UbLt4ngxAaQ1G8Oriy45I5If78fZG1tGB6XbBU7PUNG2lTZSpijYupINmgJ7EFDJ
TYkAgP8JymKuLy+GibtVyhpp7WxTXHgPKze3mplUvFaNcHkBL9fvI2JgO07qKAJ2
CKJKSUrSFqimddUh2lFh37MJsOXr+wJXqIWQFKf+g69Vc2TC1ajxI17mfxMRfUOz
lF4PLaGhdelGw6PlaZ6U4m3C6qtap2cOQAnAcFXtbx44ULXlrZOoQQDLYo8qnC8H
iqLdTK9ZFoI4dWGxRHyiU6uIbYHc0kuSjLOgwE/CayqDNNuWTl6vqe7wgDj7wWW5
dDWm4a9tl+dvXSXbi475eMfEWdGzLUPJ3kevuW4sz0QHBbbmsDYyyCfzBPBDAR7I
jAXA7fsJW3Pvv9e9+fTbjG3siGaVeGW9/KMciQOM2J7tqoxvwEhusjttXzWOhnGC
fYnRCvV8xk79AIxVBuyfqZQhBJtkl4L/PNrIjqtBaVqVfnVdofLZ3OZmI7VrEgxp
YsYZNXOWRcfOV6hpXEQ5UCiMVCMOCbEEH7FcUERdIh4+ekBysd10OeMa+LIPWPEI
cYNzMcyMzZ0F4M6uaKul6NaoswyQL2ZKyT0GdO9RGVx0PWUSe5rcuyIyEaNu9s/k
s0FnH0cfmpSJaz38eqHIooRZEnpXj3UjtiLlH8jLgE62gbdJkufV17UHumZjSOTs
LrHuE0S64rsHUzU/xv+oZspoLhv7rdJXBGSUKG6K8G5UqvHjIzYZ3WmaiPd5TIzO
ab7hmdOiBghkt9GqpzQUMJFLYYhIEeEidRr+8eAfefSgRcVrAOF7EeWBqmidxmLq
5+nXrsLliXbanhR8rEo5cbFjWWvXkGnFyf7k5IdSHI1AKTTr7ww1QEwqLZpcpkOG
UapDI57CVuGZx2gPHOWRD1RpeD4h6rLztv4FkhkDWbCk4pca6Itf/KYFNanse/cW
DEecrzklFFjISbbdOEPqGK5plroIKqcFrAicATUKe9RhzBYY4Al8xbl8QjBsyJta
EUiX04BsfjkPbS3BbTdpiShKKWtMhQcPO2vC/k6Bfqx7CYdfgFw6ItWh4qF1POPN
ye5hPAgxYlgQAOvewRKiXYraWIm2fh/qMVLOYgHtiXGjdaBDQcqP4xOw0aEKVV12
r4FBHdw5/qiI8jX8SGYnNHg/QoYhC+rqfUC3KWmrDgnAptIG6wXuauJEQrW8Ce6Q
ABJPazAwBe5VW5Vw/j5UsuVuvH4BZyo4b21r8P1foVXj2kFhZM5bibAHrZFxbRaS
ro85kPQj6FRqLUYFMaU9+YG5MNLZQETR+zf94ch4fvjWyAfLsC81w0CImf30IjKF
CyjGIAUNYdIOysU0p8+FmVTWOP90ONgiFL/CVG8W6BY9ZTs8U5CdlYjUEziLqJ7p
NMTpez5kzUo/pak3xE1YgQcd88YJ5PNeTWJhDqyN74wck/20pRBcqirBMrlWXZ8y
Fd8OtrQo+3D6hrHFO/5qpp+U244zhuPGrrURH+xPOE7jHGgq0vcptqvDaCaLPvMD
l3RIWd8AS6CL9xDs2GU5KU4oSOkOZ0ohc4pHRcBp/yb9xZm8D/fGdlubGRh97UUH
mhOnAGKJG6BCJIsmjaqGagGa1SJP7o8lz8VtsJ4gRwJWplr497AKJN8wax/n+VJ4
KgGHqMpIqQssGcQbQCmVnoq1iBTWAjYknHvvTt+nl88KN2mrYDV5cJFS/Kevw/o5
voLYpVmoXQJJoRfw2MNevERU1VjL1eL/ikkjn0iRP306wuHxjwkZ36DQSMGKmGof
Xi704oEBk93Sv9hK4yrJRw7SNoCcnsmZt7lEIzg6RjLcH7VlvJYlAuX0SNMHqoN4
wUXo2UtItZ4FCUJnE2liLGZ6oC5DmqxhT0cUWH1+yWhIEHP7tukG4tgfjr9jMNl4
9fMmpwCctFjq+DsRPj+oYozLUvVReDhTY9Cy67d9BSpJJRZowhZrFgrfXBuY0E7C
4iXAKnws9vfbkYT7B0G0ilSW2H9RSdZgFyxwV4oCmfFgVJWY2VxeEn7wde6Im6kb
1NcoEEdB0R8B4zsYcqrQHpBKrwGsP0pXEkvKlYPS/a3ICKGk/G23rqvRsLJbP/zU
Wf1yQ7PcjC1CUNqLWaiWt5xvcC+hb60hMUCg4whi9Ga+P4yOQ+/LL/qCCOe4jDau
GOZ8BIQWIs4a+Cb3MqtzTRunWcto0+JuONduGfsz5V6j3lwBmwkrIDBHFe68uxR3
EVv2Dzsn1/31EWFkbqM7JCnjG1+giCaomLl+SP2xbAK0NeYz5xYSNRwTwaEDxgk/
BiAHS24oZ9yQQp1K2R+UPbcVpJxNCVWdeoQ+aAROLQdMlJVEnpRstR2c7rMETNUU
mTYCCwIopBf3eobz/4P/cOHhIoropi4kuMLFH7Gc5LcL1mkB3ZEVTO4KrcUBgA3Z
xr6QxXBTm8cGa53LEpVRMyjJTU0l0PsiriXSEg0Lt2SiPIjLkh9aTiKKRNJMWMw4
DJ+Jw5VF9GEm0EM/KTDaJgd9WPnbi7jsGbZcuI0qC5bQ7FiAxec24/R6wsQJzPKa
enLGefH5iBXGarLXhmitSfJseF0pqPYnTO5QkRYk7RRNV1PlKyek1NciuHipuZwI
6w9FqUQ1XksW9/VB/Y1MFqqFO0TUBoNYOFgS7PgjgG278j59cCYE5PkoG6pdSI1q
dnW2IeWg8ipKKSjvh/gE8Q5UI0iCMvhTgs5HXeQACHBHeBMK+v4ow0iIADEix05S
IF/3yZMy/Bm9iJN9Mpb7ksNuA+W0WUuLib1ZK/NrDDezrqJTWjKHLDUOC+Rbumkg
BqcWU12eHzbBRHoDVABHPpGXvAKrnJrLDdshUafCHLNadhIu2azeGvu+MY4pWBTZ
rl5keDb5AQJ3wUrFtaoLZyMe7zsPOaIBSv2A34Y+dI67O+sR4dDwf+xLSzRNwwCN
I1F2sD48STQmgcv9TKhU01c8XooGRXgS1HE17t7mOmmXDMn6F2ynKNZ2wB7C0N8Q
NXi0BNxjqdc8VZ1cXow8lM1d7mvCcK35fFX8Vtdhtl/E3tgDhzdpigqtbF+HERHA
FVFyYJW7l8Nl9Nw2j8a6Ube8xhj0yLlxco0K1T18wjrWKIW+aKlwGI6h6Atuz8yj
gv9qu1tf1vQCsIEB2yY6fTwCPCaMA/VjIcvriD85Bi8MJE7eRALe15U2ZVGRRawy
IZxgFh/OlhnKuH/YrywqXrZ1ZJEvh9zIroaAMPHMNwjl2xeOu8J39+itd8a6w2i7
lz3bqC5sVqGNVR7Kdo5QF2NbY39ee38KMTr0+hQkeblXi0he0xfkayOC8BTy0QhZ
Sw7V7cFmZhOG0kkFktJWh02vkhSg5NC1ZDKHub3WGJ5zbepAGbAo6YjMKEbf1k4c
2fdarXNaR6Lm41KCiJmYXFt3R2YFSMszc+aBs/1VbWqIjKiFRg+uMXCV4C3r1MFw
CNy1QZkVrFDwUg20lPPpLrLEIR4MaVarrXL/ZM5Q+b00N75OyDM6g9rKFymf3Mwt
DFhRNpX7hyNTgwMLMHel68MuG8NJU2Ly9qYIoj96+y1ytym7T+VErUy+4XInOfWC
vUERIMkfu1N+Lf/d8vNMSMk7u6bIPcHNUzW0L+BqplQxGQGnfME8lCQzbS3ERPWb
+a0Br9OW6zJ0BL+64xdDcxzQ4c79yg/GFlZwP5GXBxTCsP6IgsQTaceg4hQgJ0Ff
SbnOiavo8LXF1KRYSg0EWuaM0X4VOOlu6tRjB8i133kQUz9NgEkkSQE8/4h1MyTw
7XukpElF17bUGcSrbckBV8DQsqu6LFoTvAUif1DPo+KQNqBEbaP/CUlxAOuEjz9M
G+F1Ep+FMtv8Hy60aLTGTGJS42fkl+gQSJRIo/uYZQCkkg6f8XF/6MieMcvXeuac
cYag1FT2Dvyvjz8vmVUAz6odET1wsEo+6NTeVWHvMB2CpOIR979yHPc2jZPhB7N0
j7dnAlVKSUIsmimXUFj8gCddO2m/vH7/+Hc2NPBNMLpHywA2m5a4dSMtostucWju
538cvK+ZdQ1nvEmt0HAuLmOO2UdlK0izEPK6CIDjRgLY9YAZSI7wWy0eJM/fxPp8
jxbgc5eToJZbuS6alvsru4bajVKeYYNQ5TNeoxQ8zECuUEVvJOp1kN2lOkLuh7Gc
zBVCy2i4Tx0AT0XSNtVpB+zC/OemfeueQ35nPPnTmfFLcSX8FO6k/rb2rKVjW/zo
S5AVebyCBTNejvLEdDJxLkkJ0OKdRh0ABvWDV0ELJZT6Dxv+yaD5YyFDL8J5l9RU
mgNF/JVorlapCvQ6iwiZ/baaGeErZTKfch06+gZv8FmWHrVIipCTdr2LzZKgymiT
zx94cPlUEpBktUu3SmATJH6916kAGptw7YPekYwMSRGjixFbUMhTlbZibGMKwsdc
ORlNp0xMHA2UNNjjFVwahqeMjBk478sGSCCPNTR93DIR+uCl6a5mRRGj4sDRaUDT
yu2ZMoAd+NrdVjNKuLEbOdsOY9cosGwg6Qp6hGKyY77GVj9TuGBWx3vQcNaitVAe
Aw+eiePDwp5CdG6OriOOWwyzR1av+w3Vu7cZ9me6adu+OIZMks7gu2R6u0nc5A0S
CxA9JyeIKU5Wh1kDvhqvwDmvMNrQsosmOeXBQfML5skhieF9CU3prS5ruvHD/yYx
4JBqIl9byEJK/aPUzYNcsHnZV2DdgiEE6wa0HH7mCUEQLlagZKH72SzhreIT+KcL
CO1iyFOFOqqLoMX5ABVQLN3qfMf5lldYiP3KWXfWAutlNip1nq/bhIRLffVZyYlO
U9roXZsbGuHsjVKlcAQsMr6K5UfS6cxvUh8qcushL/HIEyK4gahEDSqMkTDkr+Nb
9pwML8R70X/qf89viDwRXOv1MWMi8zYHrJs8EUaVPBFgXWdsCynP4ZibV9ZZo5Tu
W14D2Z+0RpJdOjKTUcMWcrdTR1dQaxJUbNk/g8+UKGdBxVqCAO+riMXxGpBR2K+m
mQGGJRd2Diz2oinqYf+Q6JWfqDLgxNBMiL+Iw3AysPfMkx6uweQCym1P/nwaXUO7
KYcmzp7JToSTmzX58/KnFLWaQ+YgWBFU58RhMcWdzGca1oxdF7dzusuyNyNa34NM
ytN105sfX2UojnzJ3K1vAxJrRfhPoEJ2jhh8YMfL8Gib9YB4HnkdDFP5yYiV0Dcl
NwEs6JiKxpAUGdH+oppqQlsMsGFeK0AVE52gKJzujv41wJLf2nb6X1VqoJYtRqq0
4SarKjAoPy8k6EL0LH3ku4jAMsEOeX1XnJest5RYgC3e1kXk2ThCE7wQRWNyLEGU
x7qgvDE0j08wR1O/bZ00+2tdAkjW6sPXieDKYGflR/0dXvDzBn8UThdUUiWj14oU
Gr42dEuaxbL/18dx6sLLmqATejYf0pxDOSL0OiSZVeL5/dbQ2WERJ6m7X0CnXKuQ
K5a40pnmO707pOkCBD21KD1/M+SQJI5V18X7TL6WRSkX+rsb2ZSxHXcfofzOmHqf
/DVcj3E/2u7lSUF5f3B/Wdx4Tac1k89rqCOE5d3klpCNlZF9ymseHcL5+F+uamlP
6mFbdxkZDd+PfpmYOt5yDThBxGa6rjuEx42q0kn0hEh7Aw0N4gxEbjz/qNZONnbI
gkhk2fWDzqtNnnYNM2o1Mh9ykDIpw5jmR5R5e8NutsQN4OJi5bPP1GmMLPu0QMbH
fP3TopNwt7RECN7H/Oy95e7iPH2ZUYpNvV5ayoQtkFDjPnKahJA/7U53TgndxMMc
MgSIaJGiaG4xoCGF9WdWk4aIdrnuy3HY8Uln4+MgEuE19GvpKm9QoxVdkG2bf+jG
6MPu0FWH4IkEGcLzewSScxKI+W0x0n22/9rFDDCp2Dc7NMzL4aKr8vnqjIBCf2Nl
kD2rADc3DEBd9zERYTpDTMXRzC4PuYuEXCydQFZ7zkQBOXfPpRQO7KOAhX38fh9V
/9Fpgj7XjKLULJsNrgRY3MHjcLlkncwS2SyRBUGsL262+mRleESpI1EoLsPTK3qO
Dx/tt8v5jeKSRkiXOb/wgbbm6B9WltCWsWpgYrX8YoG9/5zAbZZ8tBoCBW0Tchb9
Wg6/b4qPeChYClxqQ9iqIG7kpJtEcpVZ76Pk0Yatkb+5hHC317V7R8KY4idyY4ZC
OzHyjcc+ljCapSCpl3DoGdIoMXgJ1C8ak8YmhdoWJdvL4HSGm3/AYtCiLFC56KMG
1jj5BpCpBCC+pBaTv3PcqXpk2J+DN8VaCQPTfYcMBqHVIfSJPNfe9U3n5hbLeGhc
SwEQuIrmztUX34J/YW9Arj0OF61RIng5PdhJKPjJ2ZTuyCpuFzF21eB/ts7H4yed
duuTd9vQc5aAB8E2TOKhspdVVAgYPRMT/QJXa2+v5Ercj4YPGOvbKF7CVcmQJ4vI
YJyGJqCvTstpIsC6GmGes1CaKxX9Thp5+1/Mr/W6t09sfZOAOucEygb4/FlnNk95
llkAJblMxBqF6DRdw36T02bP9YNCwMfpY+VnhnEQGLzSPLNQiRUljhW0GbhJcJPu
fNl/usgfLp8cbE29prkal26g2VEqbjbUPLkCiweBw6v2FD+Olrix2AfSd76rXaT+
/Lrfc/gsxDPRoFJHcEsh94lIhudrqWEI0g4mouLq01eRU7IMA8QfOvSGH8hufMrm
PlN62h7h2SXG05gg9BR0RC+w8mKw7ToPpknSYBKz+qh3xO/Q2OlU9BaXH2tBiyFC
SN/FapW73HELw0xFmMU8D6IkTRj2PLYBdQhLftZ3LSUBGwbaAB+dq8qO2z57oSAz
ujx3/AHLj5V002iiRm6nV64O7deuHE0tiRhUM0T90UhEqqnh0lK7JNhxqxGnveXF
9OrIRrFRrBXdhYxrin0VuNft3wT6wt4kk3BDds5Vlrzrs/9ffR+EQZIW9wXNypm4
tvmTNUEytKHHWozsaYTtd+HuVnKzKMR1wPFZ8CfDCJ5dOUQPKjSDqfIahQGNwCL/
1vrFpeWv/FE+VDX4vMh8o8qAjlDlUIsBnVrNswVdvre8qfC0PEOupffpplUPIhzQ
NQnDGAff9C0M1b4UXH7x8SDghfV8WyOqM1GJby9sXpcUzDpVWTbAUdWVTNlLKGbK
stJuBiHXfP7c6l9/pjOL8ChO4c8RZqUZD/06Myr6/bCDpxI9Z5JPdjvat+trPzgV
q5wJP6a3E7U3savj6lbDi1ZFNJ3DSFXip9zE5FP6hXbTuMSyojO3xN1LJWHIFRGr
aocGIEXIHlQzLe1bTbMejMGdq4n1d0uJxxVYBlTWnv3QJDqfI9WdxZYodd1EjShz
Em29KKias2xWK+tBzNXLIYe6VEox/SSBs5XByIMcBlHP1jFLflseDHGhhDouKM7L
qxSGK/s0dawfeyhwujQVu8/9SdONL8++4MxZ/6pxZuiUCaNUbW72Hjza4m27qdOc
Lv5EYoBVCU0nlqjm6gqYtpz16dPb4jzAV6tambIT0B5eQ52UhK+fX+yYVMSdi3m5
GCHzJeOmRkuAgPVC70cCdIZx+YS826P0gz3ZYOreAR9OBhgfi0akbnVLIvhBNnK+
9z04Zg4Xt7w5yuSWFzt9I6nBQl3kQw81sVKKfRBsb5f9QNragiLMDeeQ+RcBmO0B
TcyAEvDDwqhMUFzuGXnZebuI3s20GQWQakUstLwIHgpOhYDGc26CZ4HE4ul9Kiie
d/FyYNSAW9bHExaqswC6gAEfetemcoMydU5x1k2WCImrttWf6k/Dj99tD3pJh5Nn
XUAuZ/mHZIWAbhkMULCM7DHzB1d3M9z2zzau21n4FyOS6JHJQw68rESdr2PWkhVE
7B+na9U73Qy/sGxsIbQjcu4/57b7OKhrC3/BhkDwDf3fOWoJH8rdYbU+43ixg30J
swCCW0I/r2ft0yNatpG0czM8xHxxJiogqOUoG03IT4KLjU8hG70PWq5j7BuAOQTi
nXQXOqdZalkPvebrmhnAI0INVo1uUnj0MMJ8ZbqLS3Cbk00IIYta5mdaWryyZPHO
46SsTu43Z10xfEF1kr1ei1Tixj+saTqg9u6go+aK2a0LgAY7S6BBfrJhM0FyAxz8
4uAzwUee5M7Nk5YjhU8Sqw4RCc2Q2Qg0ad43LMpnCc+Dlag5yxbgtWY0V5YnIvB5
3wcx/YDDd0OtCCnQpQdODk8mcvWSTHDF3Y8vr9KATfhVLoJyTpUARPFCi7+AeApn
HnZGRfxiysjTMdcwZLUc3LcKPHK2u8RhxrSS0IxU9DTsTFl0rEzSdro7oSzBjgyC
jHXpO1zsthZZRXcT0jVnhm1Arkky7q3jY6ll/+ldT5bRncV5xuYv6jhSiYeqg0Jn
RTdV5SrouaSJNLY1hydNFKGu8kAeiaS3pMY0t1hA+ix+Qbbnyc0dR4QfdhNpjG78
7ah3KWIsKZ/XM3mQsQ+J8WFEsqSPIUedX5bF0o4F/S2c5TrUqXFgcXqYMV4x8Cc8
JaaQJkPXWig4ucSU2KGfl4aGjwKWdPl21h+iuq+ZEA92YRyDqwTeSC218Hr1VhuM
CZzDgDHa+965NFH9G6PopDjlsqNik6zToTZt+C0qXEkVlsSN2h4F4TcRxbNMk9Nl
2ANXrRuayytK8hUFAtIqndODGKtfXEyiQZmtakwKcYtqgpczo9ZKUou0KNv1orGk
jitZWatjbAUePpl0a8GNm+dV5U69knbPvCX8yRZ+OM4uF/Z8+KnnlTW6ViLYrhzC
vLXIlpR2HGLUilyJIXX6QSik0Ff1AmHu43oaPhsBfdRF7w+Dk6jvohWJ9LrvvXUL
nrOdDGKX3szPJBBO1AZV+08eGbvBuqxsyQtzWUN8owhBX/85euGC+yhYjw7+xnxe
wNK9c/cMNb1/ZhQN8MnuVCNiBESkWod2gAo0HHnwXLj8mRDV3hRU74T9pIWv1L5B
Ejc4jzBl64zi+H01/u5rHHH/Xeb9dSfLWiWRvi3JxMa4rKRdvIZaeIKaAcbnVWXv
jpXUi2H3JspnxgOdtiTB9hicXUug3xrcuiyVbdLK8OQsh2gZ97EpUfkFzkmIzcL9
5NHKdkqyhryrUB6Qx9Vn+REutrtayRGLBB0soO0EbugTT0ocOP84YkUkZcC05/pz
RHaK5CX3IPJqV4Svb983AaYRqEYXgNFaqrU3SZQSiiPQ0ZkduUdl713kohmMAENw
hSUDn512QdtQlNupmYQ2rguHvmDhps1aPHSB+A2kqQHUbFoExpx/k2wsvdeVij6A
SLP3S4FjXrJmONlSe50d0jCYfYk03ML5+4d6botmr2rmVKmIweFaVpSjtQ1tL8ue
hV2qJeT653hJ85z7MAUHHdxlaLhVuKjaDrc6zyRSoMp/IRtxtsLsNcoSWsVWhhce
QkGgFv3Zg/ljoOmBO+K9BR95AELdymECJCmjmYVyMO3smlsE1V7X4tAH9OeW3ySP
SXm63zu1ifzEDuEfr5tv9s5j+bMvWlMNqVTv+awL8Kc7eELLfmaKadLI/ujmCxGb
hZRujVRUiXyv9XnYEFa12MYYYDsqKqLSNuM5ezp6GV2XaLIaP8DZBC+3T0veKBTl
efnX3M2X9gvgWDOobNCCxXOY0cWZwHsfTVR+5o/MZmxItKph8rScR9EEmi8iSmpk
6GwkNKCNMV0v8ICr9GTCRA7lhMsNL0gMZ2OEXKWk8C8mQetDxeNVshWnv4GtxdKV
QL3cHsho8uthTf5d+cesPjA4dFRJA+H2B6UVGjR/zhPQiJtBaiyebyjL01AZB8Q8
RjolP6ZAmY6AGADnw6AWHJQGN0we8HBFTNZdrmZFts/Y2KpW7fv34qIf+g0/nEsD
gESn6YfP1CuW0dMCsPxANBdaA9IoLJ7edl9g/7xJp0ifbrTujTEk4UFW8yS9zenu
MATaKgCevdjwyP2YEjd9BZsGwY+WfnL8S54eeicOxsmxrYqinvZKT9ox9i8JOL7o
oAvHLN4/2ynvnZa/ECnwoRhwWSGdCrEHb+Oji/npuVAhCET3g/cKv/Eak4PxNx+/
0koe4zYqABIHjuF2Nv6/q4grz/sqiPayN2BQDq362LPWnpeVJxnS1kytPe9vlzda
3nHI9jMYufyvwewXXGaTw080I9S/QCgDRtlNMfpB8melhYnV4VnWk6PpCILK6dzt
yKlUgOdeDeEVflSNeay/JbBT2LbUf7JnmG1451HQvlaYxeU6rp4BT+cNEd2avCwS
ptRi6gB6FDLQJWaW0C8FzOVgvICxCIbq4pZCAmpaTez0q3Z606oUwxea697BHxkc
HhKwFsQEVKu85b7u/xhXWIsXYr60dUKYZ6jFohIhrCuFqMrd+OceU3yTMR0cDgYn
yHfayIyIPkAj4k1AralWZraIXLkLqe51K0/KPNi2RRYsNGUhaJGM/2B/4cE8oA+n
XsXZisqwEBQmHBFxAOP5/IxElSBZg/OJON24JgbLEH7APCowN2whZeDZRbg0LeLe
ydfqAF8VRxW24jM/vfPfLkbcZRO78UCDyMlWct26zeE7c0j69RowtHyHgzKlhwRe
NZIKIu2stadJzIgVYghzC5sO+qoZpgDH2jeeHX1tjOxFDIMfGNxulmB5Air7gr8v
WUrepkTaFfXSJdB4Abwd4E/SLnHr+Uo/YiNe1vduzayjh/He/LfAiAeqT1BRnoK+
p0q0iUQRCk8rNgMEMiRuyTqwIsRXDwe1mZgxgcurZdI90ps3uuHhuocUOhDpJySt
u+3PHNjgns82Oo4zSmNGtctum1yBppziQwXkaMpuLYTlR7OFuZWNc2RT1D/nK6fK
AONpzwoSOklgBA6Ux0M+nXShem2WQNUjzYcAYyMrRt+mw23zG51qXe6stmGqYMTN
9QMsKTCNx90mv20xvSpib0+UtBtPVPeH7aGCtj4QW6OJDrcrvbXghBMe+AuAM3vL
5u6MlDDEEsW/M7nGV7dNtbiK17cWuocjMbm9dO3N3Ovxd5jzqhq2v1RYljH4rtiI
KbVlBGkB0CbJT7dIX+9nx0S2ftXDaSUpzAy3A70+nm68vd9EKGurj5lfZm1Ptez6
ikJ03C+gWriwGwZOxy5wngw8eFC0CQWU0dLseUI7PM1/LP6MMGX/ybgxhlOkkOzZ
vm/I73oq3p/uwmKLcIbAdlZm82VJ6j+m8XDXW1hvak6jo4fgwlzCyqYwriSW21+u
5OdhDGiLDUQkZthrf6e0nx2RofLipj/8AWin6eC+GYScTiyLtCU0JIq12S8H3nsq
dehTHu9bsv/HW2WwyhnePzZUlAMrldP971xuiokizOXUcX7DUceOOrAWqfFX+EdT
T9uqesfq0PziJVUYe41izEzGVJuBtCsFLlZaBOnrXYIDu9yBS91Nd2kBGyTZFyXa
K9tUggYedyfCjNQkCA2R1taz237bdzGmmI0R6EXCIYBKkUh7oqk3dSxBJh++FSXf
WwnxAdKThh8BSkeJimp+lRxc3hxW4s/rUotL4lDqrZy/JLFCrj3ML0uAEhu+5Hew
lcfF9ceI/h847pRgxg3g5HpNINsjEIdMtZyFsdvqqK8NKS1kCjZAovFIkyD1GXDn
61dhjH/HdmHdVOhXoNI8x/ccS2bNyrMY5AsJseAhdKC3uvsPicP6+OOjEt5Vlm0A
OQZl5WxfzX/1+RsDNg1ZSrYKEGQK9Ox+AocgM3CAH44HT/EhUDO/9wxJPVv+aYLk
SdkntrgPA6jYh6zLIo0o44QZ8Y2dBN0c/iIZmqnX1aO9Lut6/jm2UyVQ9hM/spHt
c1ZURUwXMvFzwTI1kjamh97qNQp7ZnNjpAJolbozsACX6y7gRVBf0fIA/6sDJ6+5
/NAOtjrGfLj2UICTW+8V1tuVNT486wgsX2K7CjyckGJTr9uU2hGhqp0R6BMapEhV
yoS6QBqOFBa6BCkE2lFSp6jW9Nz4OKavMhf/S5hgmW8k/QoqDRe19YigNyh8Yeg9
1VbBshYgmefr1xLGEw0EsoXRx9zvcPJjoeqUzrpm1CPdprtj5YLsK0WES/+iNzUJ
9gR8zRndJRkA5fELAIC6J2wGU+K8MEpTPF15n3XJ/VDNs05Z4QBaDIeXZPsnOhIY
XRaL5k9nW1D2H3oqnzUi1fCMhmKvhxs5VjuaukpU2+gJ9+6syQnmPumG0FZBx+LE
bkdpM9/GS3G+dAsdr8kLbaB0IZz2tTQBN37hoI2MsS7LaMfozTRl1Y7f7GT4DJo4
zHRvztdger/mtgZCqnB6SDYz1LM/LRj2ALERA8oYMzyL5ATt6Jt3dH7Pr0N/2pCa
Tfqiv/wSpRcMrL+l94382yqbjcnxIEC/egVt7Q8ds+426VlFSOrhHz2+j8OOA/5P
8/aadKowSQYmGgSzyq77pDha0ilADSI+HaDMDf7YVLUVnHQmGFrWlKlMdyhR6u+P
P/RXr6a3yGS8ElQq/ju2eHlO3JjTtUgwb+cvUPPgLT+c3jeMPDXX8P5RQeCA3hP9
GGUKCJF/yjbYPQfIggjVIkt0BZNftYTRmLvODex/7a0/Z/xbUlT0jWTy1GLJK1Kg
QXwkRSsoTeO8d0Qpq/B7cIEqT0VLinxJ3USFzFQpv5Ge0TLzRwl8jG+j4rIYDrYB
C7e9CJn117FbmJ2qwZOREc5DdP20OT0iJSyhKWDbT7/DhFNC/NeVDnZENZfgFfsK
yNRSVisLnUdjWPzvcqKG2+0wTu79FI6gdfYBZDhDShsECMrsaw1o2pOafTIo6g4z
xXdUENUs6139V5KHLWc1j6Cb/YF3frta8kMsm4SXBdkQn9PJTCK65+e3lLlR47rJ
YwkxQR/gLQaPqK5Tiz5mAAjh4bZHglBr4RdvDPkxqGzsghY8fy21XMrBCti2tb0o
wAo0xQ94BBmBj+ISzKBaS+7mfJ00OyouJgfxQLUAdGTJh/UdmLpBXqzizt/6hlHr
gY+T5khRySSzTmbDJutivbARN219YhA466f90ToPOpbU/m8fItUKnUCazpVL1Tok
hdPbpsNGKXz/N4uWLXp8A5FEzswwqtLi54EUCz7clTggdkM/wtf0ScAXvu4slJhP
Dcvzw9Cd1NoUsD92TewjDxr8VPP6VWw/bszQCNS0gI46vGeiZHtV1WOWlWoTqaqS
CMepEQmQ5ocdT9gtCTobV3tquVdZs1M6QDzxMPNAeST6yKS37E+LIfiMMoQWmU30
JoJH1gLLcCMyZUzWmIzI0dgFqG9uzqHNac7F+45TXO85H6M8GYOgEXlKOuAHpmkE
wI2Co1y4gxlzLyHNDLjyA3GGxWOmFwSwAui0D7XsoLJMYHnf8QYPhFwCiOq8NkP6
N0iX7yraGfqm9TSlgL0UsoWCxCzYyOo66RrXzv+Sgq4gvclhxX/fyQaREy259F5Q
HPcNFcg44Sx67CJllINnSjKjBo7qzBvm4YPQEMZ3cYWFHgFL0/fFj4eLrPlhoC13
k8jn++SmC4tq7eCwMTVDbqyjHIIgEQQae9y+YBc9gqv59gBAY07x58AjJspY6/T+
iWSW80YfPkjLYwOElz46nxAXEhJT494tZdFdjVRHS3lyI5pr3BiSLKlCKvc2jvEr
MwuVgn643WUix4jl80Rb2e9v8+agrdqYT1NTdHZ5YP98DcL+2Zd7eVGVkT2hd/Hf
cDJgZgQa6/eBwmV0poD3tkuO4JIEVstdgO/vf3K6YTqVRdEkXXLRR87o+fpVPW/1
Oy05+ruiXGlFtDMN4oGk1jIakeWn46Vm5g3cRE7Nwa1jsE2q7cUQfB1H/Dx7z0hn
iYMFbfGj9NLL+yTV1f1FouAUQiy+o6KCYq3rYuEgRB9Bq0+Qh7aC5W0uqwN4NBww
bmfsYY80G1x5CGSLWuqCPRcUnl7KsWVAaPUNK6AveKobRjbiPgyOeg30spT66Fkm
eOqvA5xC3FNxo4Yok5wn5at5RXJkY/tpzkDGwUi3pvOHcV/A/Q1kl1rfyttv5KDE
cCybiefV38BDr1Zr0qFJG6YosqujHawW1Xq1Tk9ShGHK6/ihW5ZEMfel6IMOnG3e
crp8U2017CHwBbRuMjulzRpfBu9pKFlPtsVHoYrOnDwLAcirpg5frlE2WEI6Sml0
KhudtNSErn5WGorSYu/cGPgj7hdN0kg0HJb1IO8z3DATSjW2RUitUwlEZkJ/gqJ0
AunQ25cakk0d0NSVVbvFkQKQC8vDgBtHpudogbaFS39Cn50FMXjh07meJplMO8Tc
Mm47XnoO+4cLbgRDnmacWwwolEp+HrU6iX6DNjzLM7zv5cJkkCuItRQyI0HndtHd
/JiG/k6baUZReS7L9/ug0XLFaEXkOkRu6ffg2AgGgwCBVRAVSXmyFi8oqmAaX7z8
E/rnJgSIVXiUjdnhJNDZKZcU8qOqR3bDaEnHOwpSxKkhbF2UyiLnPkdrakfXR/Z+
zfMvlKqvJCzuxnHDCTf4r/u2ZJdULE77tANDnxYKl1QR28svsdjJsVmH7HXEwLtp
7omcxTFvM2DskQzM8vgCA0ihdmxOm4wpJuve2Ou4X655bwhyuZPls6y4jIgGHOkk
fZ88guQP1tR/0MdQPEpwIs2wknAffceMqcpd0dhD16XSVZnw0pGhaYyFAVKRVmx3
hpsUoHB4KmYAvhB0wubZso6QHbhCxZyvE4H21GzFVPdzhUirBKZaakXg5/UNpTER
5freaz2E0ZS+18yRbjyws9veYQHmgEnqAQzDmAMX7QnRry6FBR7RqdA2p+3TGxEA
BVXcUH43/3TiwNzxDcQfEjjRcQnqTzf/F7fDtM0xxcHHxZFjg9KxukhHgS4i6BJM
IUFvYmSNmPXrSgIvzK6B6UTvULpLe3SibLyAZcHu7IybJZ6BAzFwYOSzD4fMcrnU
V3wF1AhMYKrdmhRIHLYKZ0pYZOMy3mYTswSuUjogLu3pqfqsm+9vkOkZvhKHQpku
+vGs3glgksIymg6Gqari2GJ/gHn+bu7P45DcUIPvPPDKdhu6y1PoAaoBEoDvvDOm
gW649rMblNcQoln2A6NjzpFRiE9ul3HVmJ1g2D8paECuHO5KDqz2wccTHj7g0wLN
zJp+Ow9wnJt6Hs7VEFNy3Xwk0gE3pH135+Ql6Bn+C3eZEThX3S6ptvSlQpz+ofgu
iyS865yGLyqIb1ew1xPJvjbernlBBJjrStMdOaiKkCbCH8LeoovBVLFm8m3cCBmz
N5+Q1geig/ERO83IeU0jLX/avNhLgaClGF1WUcWr9+VZdJX7Xrrd1TvOce/MZ9iZ
a7geAp5E7MnOO+DgaqDO1Ay84q5AzuwJw9E6MtSgckGcb/bu3Ddq8VJmQGIO1Zsp
GvhVgpXJjhSq08d4GBQK5Jx2+aIzX0lSkf0ly27Z+N55mv8ZJFkwrMromcAiwH7P
ZDHqdHsiUVj3tMcB0lR77/x1Ybj7S1qRtY9mZNflqOS+kJNi8ODMxsWJK3pjzbMw
gkRrD8iUr1/oV5gRqgC9Vuo4baMekaVobhmOQVS1Ghquvd1QflsTal/E3owNxOW/
dHZNpAxiE3eZlT01l6QuZxouxkzPiDQsmf3wPmZQzevITf3zVec7+2SqeXl1HCFT
BlSIzRNKX8LoXP9A5c7gNk7mBYGFOT6liG+3dXox6u1KoB03Tf6oUt7prrlOUJee
KG9Z7eLgbGFByLvZqeUgttTrT7WFs3t4MIiAwAjy7LwxRa7v4cZUxfGBybFKqizn
IWVpxDqxVo3Golr5yCxTeNKmKcSpZ98/H9RUZSa1HerYuRCxVa4Wg6KZ5iHr64rM
IrEE+TL3NqmuCbI6Ank08bPniGf7woRHdecVrd28F7ck6qRU43APnSpyAAzrb4X6
nVd7GvPFaQ4DVQK5MtDR5L1mch2j5yM1DSIPfJ01huM2tKc1VRawNbQXVbS8AVh5
cBhqNGH437VZkF1mVh1ssBEYMmynDU5WR6F0M7iHE2Ha3zBvNMY6kyUiFzMwOgcZ
SqfWzST8O9Gbwwt2x7uxJRKRkMPX065ecKszi5lynblp5RpbqoTx2g96Hs7ONfUB
jzTbbZjRBZ7GrQLPKkHW5ei+Ih5WC7hbML4LI10rZLInx6BZzD96v/EA2k5llX7Y
9Lugwa74yfqv3crsRYXQsV2mindSJ462zAE99BuCV/yaldvU2oAyrhLKfBWwWCx5
0MI7juFybm/bziPA2VvstqQdnWHtdl57KcyR3e9LJC4j/jAXaucU336W9qXv4Xa/
KHf8qRuCBzjpP0ki/rbCIIVUUb72KsrCyVk3e5k5lZizzcsl0rZoyRuP86tuJeXJ
Iza2gSWwj9I/ZrVGydjpIWrmM21HwtePaS9iggxA5XmOGyfRMVlwxuaTjiZ/j0oI
+x4CvO4sKDKyyKCSSathu4vovbJdUX3WWvZ402DNowjyOQnfBbbJUtHfjfq1cl9o
zGdPjxfKwxL0tf8PCwNjK8rMOH5AtwcwKdZsZLmqpb7sAeEOT/R7Jufae+zeq1j5
y2daCiJDG7DJKsXfDya2ajto5lQbG/WueDGA2iHVMoUnjzVDujOzsBvYXulo6+s5
kxh0G1x1zcmET3kc15ZUoL9BZKGoShiwdHNhO0QW/HE2MsErV1AzgU6GrVcYwBcG
+DbCayKrnJFS34qZhbF+4g246BaJ6fFzqp/Gz44ZjBToiyxvPhi9i3F6hMEjYSEV
hZ0wFVR8lT4jttnyA6LGvzvDGj07DiGNOuQs00CDWGP5mH2ZKQ+cNDWLCYnCd2RF
BOnPwl2Y/xaj8zj6YlAFrHsp0EGDOZC0eRDd13s9LX37W8+2ktTCPThO76Ewtm6M
7/IuQL6bL5uvk9C0ccXBaRLRoeusrv4N2zoPUND0RBELO8whdk64KqImyscEJlOW
BQUrH4y6qb3oJ253zfvwYky/3VWeBAFneQd52V0EMzhlDX8zhUzHsbALt+/X9vLG
s8XWIqgRaGXK6T5dToNj+hjYN59koLR56DA50kJIn3u9UVlfDnjYWYBOlLPSNVTN
8jhR426VDEN7UKNeLGRbIvx+GmdVDbMxPxaq6HaqvGLorT0k/NFJUTZxNCGNy3jQ
/XCT3JKRyE1hYYlA74nf9zaik6W6DV/9c5AoFTGL27w4iglinApicpntDaMEiNA9
6xQdUi4M0DCNf4LRNfeR0u26Gs+ydL/rfV6R/dq5tgpcOib9ksq9pN19UD7Mk85Y
gYM/T69h/qHHw1w1oRZM7dw7Z1SumQ/zZiZhgxlw7E7Y6mb9MT9H8yXcmq9EVgNG
ZY/615JV2YkzwRhF73yA5QKOCWTldioyJIxLBAXRgrxkgZbQdX57ox+ZOaUMHONS
42sp83/sVUuVVCglJIm41kDn6xKMUKXl21qKx19Rpnh5mghGB9q6VfksDEiTDn7+
cH34zdKZIDai21FHf7wClYfFpO5OyFG5Vaa/QZYZ3vgLwrJhcf4v0Us0ohN30OK7
J8cLzdDcV5s/rGtjxVeIYbGYpfUA9Ig7dXjqUwu+N1jjxkTdRT1OZ4duRc802FvT
MENxToDHWj7dLmGzLTer0CNVpcd3MfkAGrRyzIc3VgQsb+LdizzLi0ZZT7WjmF86
weaS1iAVJEf5NznxtjLflpQgm778ZkAViOXQJlBRki+QGPGjsZysbYhfD9pZgL0l
++2iJPWuon32wyA/5aaQfq5GIY4y4zPGdcgXwP55YY3NUoNf0nlS8qBX/11SOrFD
TKPhvAL4WbMpxu/l9PgxNy0TcDs5eBrTJ4pxTZg1Fya56MZKwjUmUrJ+hJkQA7vQ
M8+Jata36CaO+v14mnJDE3J0X7LA2W4UUUViHKtDjbbRo9pM2A5YRyHuWqpqDumw
I6bzYosamhZIhC+MZWuPbOziB9RMestMB6Mbm7DDSyuo2JJQ48ruLvw72xWA3trd
O7btpdrlWqYoWqKfL48eFXTHwMbxZTaSUlMOxf3pJBPCaN04Re+l1VvVp6iwywYI
6lSoEt9JW5ZR3w7SRF/WQbp2wnuVEv0J9A0UoJUGZR2gJVYlXm3guBD9qQ+n2uaX
TD3ZKylIovZ6pnVJ7Mp4GWMM7qU33grM1oHLycBjs4xzgnd/Ag8dUB9HDvHP/f1j
+FEiswAL13Uegwt0kaN3uOXZmk44pmUNRw7vL952yRLaiix5RL2NpEHm3Gml3+Gi
vkM07pXQs1zD/w/SsD/0SdzxMH4W4zHi0vFjdGm8J0IzrUXjJ17S+s41R90tWRfh
EsuSjS4LLFl1MYu+8EvVIJ6KN8hwxIW+nqWvJzOs7hkjmcLjI5VJboI3bmAsp/ND
H/LUebIW0Nl7OGlZlViuofQGje75yojPqxrJ68iSDY0oFk7jVBS72X1j19dxLBEf
w0jmueeN2zrlbCeKrKtLQZ8ZDVA+XD9gBzEKg9SJ5ebeXJGcuuezNZLWuWUmOKYK
Od/lg0MnkOVuPTx82RTnVUJS9S/em5KtnxQhALBxCZWDyTCPNeJaPQAmfbda3LMZ
QpAWA4HKOiFIyRudH5xbGJTcvShaFu/eSX0Q1mKrvl0beQJCOnN+9aNorij7z69G
0zYA3ljy8R4OYRMSPb+XR5Xtc2CaeF07+ezfa5xzqeka65tWDI95PqGRYCIwaZxk
pTTTwkRjAdVLLDBZ2OyhM7nwzaMyNVm3J8pSbgQS7w/1znZq3JAOO5NtZqV0f0W5
Z9iy8YU3nVwnOROQT85omSjvc3hIQZHucgjyeTvAMm0zha7wi7aqJ9C1TwnubPb+
RruCpBgWwwUIaAWPFvXNiQ4ayh+4a3a3vQ9U2Xom+kU/qOhpBy2hYE3AFnl8ob70
DgSnL4dAKz1nxuTEzlklcOFNxCSCdVPURnQAq6e3CQ8uG/lzWNQFEFHlxToIwYnn
f58/ND22zdGp3lsSjzazYq6ByVCnZU8XBHFoxW2ipLVQUR5r7pz5Sd3+CVWKD/mp
kje5EO43oduiIxxtO6+/L/7KRMq8DQW/CL0ZOHi0VYRqy765uiPyxvo43QU2vaTu
eSe9g7hhMSF2ehzO7IG6XDmsZmX1HQNrkFuZa+P6iwAfxRgZwa8oofXNlSbtB/7S
eWXzL1dBHqRolVV9udpNubk+sHso4ybHsnqfHu2y2wIURsl7R9ISULxAqWe/DjIq
N9cfrHY8aHjenIJnVFTJrZB3v3180pprGyvVhkf6za70DWIfhbeQsLDLmhihisaD
S8GE9z/d7URfJI0U1TYf7vtlVOk3+gASsR9wcjXTyuMSKZVbB7Tq0nZ0/PEwL36Q
eNBUeama//cwRftkNpasckguY8ikZdC+7IbXWWUP06/ZQHhEkDUGvBcCHbprpgMX
ykPh6aQYCSwFv3h0vL+xp212xc98P2yAZkv2w12cRtD1Fqt1S4zaMwfxT0CJXSpl
p5hD/4LpJthYSLUbcyXilfqC6QKWvnBLCga03KHk3sxKs5opudHzVBGlLGqEdp5O
7CmQuq1QPHv0lGMU592wNTtY06C+5McsGwDD+fOYFFgITgNgJCVgMeeJSU9YdPbZ
XemsD79pBHpxk0yZmRKVEr391jZKUfDlxIZhjqgOIHp7hmkSgiJioXvPX8zJ64lh
gKfWbdXW2R8lQz5QT8y1jGcy3HQAVXS4GgPSAo3d/QT7iWRxGQBhh8ibmcYUJNMi
2wxm60KoVPkKcaMFwczOl0dWgtT5/BbciGQaLQuAPypCjFo+8PVctPr2qZIy1w8Q
2upY3oN01qHjnbuak76KdVBy6YKvoo4/4BK80CX/WUKoWPvWe0mhunhGO1MKRBhH
BZ+YjHg4inbch/65i1bBvCC639RnXP9BOi9AYiNSjgippS3BmbVqTT/0FZkADu5J
T6JE/vl2QGcjkOxC+WccYWw6BPhJx+Sw9VMwKLMqgU3ZFA1XQgzaNYrv76UQo9yC
KzCLwg+XAVpw+t815yFm8a/FdESSTl94ohti/OlOFh7DatBZRu7nKglkwFhm7EBn
GiwrlF5XOy2QJFATpBpu5fV5aipeQORbaS2lKkke3A3M0FAD8ry/AgTT8oetFiBm
RCcWxZHi1ivC15B1nLcaHVDHykvQ7mKNziS2Miv7n+rFOY2hrGkWXX+D6ZMWWI8p
8HW5aWXqTCkZZhrIjhWiXgMcOxChNdnlPRtpixq3Qz98W98Hh7N6GWPqmN3YZBp7
AzDYf2LfLBYDTpJf4Uh3/kNu2SJ9nF0nbN1ndEuXMEs/9Pl5yi1uarS+Q73zuKH9
rb9AHxhY0/NyCRLActIZun1yLWLP1v3VLO0yENhBOTDt1VlSHT2qgT8vrUX5bbup
Ata+CnckoJODJtyJqktaRkZxK6aWpYVOKRwV6vp9B+dNzzf0OCZ+Nx49H6uw6vYk
blqg/PmCJbsvnnkFRQ6kWbr7cmkXIhs8hwYDt0NJWdIFuQQ/MfKXfOu5MAWpJaZT
Bwuc59JlstjBqM1PIp6ivy/S1sQnRSFJ5T8RiBbfo6dLyqsj3pY8/ujdmPXYreVk
vNHEcXYS89TsQ+df8Gb+LNOD7r4QC2NOyfXt8fxyHVjCb1y0hWt11KFF89v19Plr
FsBEKcefgtho2xsGpiScQ7rOswRJT66FyBIKcbkJzusRkh/mrmazlduc5NXPyZo3
PBUHG0/UpHpK7fFyZt4WxbWydWPdzNqxEIrnsBeKfch0NukFuLuwEzk/y4C+LqWL
fXsp9MiRb5lPoiGAnHtkE170aG9PqQ0Hj1m3BfZZwMGTTsWktNVUcCUckGy02LiN
Ez+QcDuySjWATrfr9gVmWF4zK2zRi73v6bCs3wSZglIUDArql1NUE05+NdNWMD2o
6KPuRGOwq9AfY8Yz1742XHSsUgSa1BQ3kInVQh364D8XEslfmZMN8J+qEyVstX/j
7yRmhNJ13IZFUqcH1nhznaH2b07I13hocrQlH4/7hagTbvMd+iihIQCW6IfVsT56
W4TZA4KhWheb1OKAvo5Q1NHn9y89Sb8684qh+1Qk1y+3ykE16EeGjyBV86nw8cku
UA7W0tnkwNUPlSQQ17ffrkUrGDPn9K4qHs6nxxc+YnAz748Z4IP2lTU16IUO/ZJC
o3ryzed8unVtGeebBuU59LRt/MXZR1UIvfanamGWxb+r5NKZyTyjjCy89IptRcfe
pFPzAOK/S68TT4OO01dSZPficcz3Zr9fs6fMGWOtGQuj5MO8k5dsmIqGUWzpcRrg
gXD6Y2lN/cFYtE6/eD/kzz9vwl8voxnqJRyZtsTh8/57z/PXpXxvm+7nMfV7igLb
44afzONwanIWt39T2Oj+vn1QKLalq6LuvWZJaJHLAtExP2ANMRxnIwVrrN4QReJI
miFmWKg0z7fzpLVJmjl2zX8NM1YwLxKRYrkTSi+L9NLWYxsIeLh/xzcTtSGC6YN1
UGqEjMlZEjSKz0AQmkJdBAqVVVJC/zTCT3nfpqW85bWbvxN0LakduTSZp1vM+4El
8kCxJiPm36TnLWtfoDE3iBOw/R2qAMRpJ735IpXwSA9ZuV4JwXrgb8Q543irISVy
b1tqPDxXiTqT/WfLjtgtblfD6HffLpJeR+uT6jptnvpWx8oWGddFYORCfiw/oXSB
c7Oqd4BU4NltvqBCv5c3dqoFvw5UiSg/N0H4UUaUDgbMB1SyjefwDuapZNCXKgb3
EIRirr4Sj3qhTOu0gJ1kA2L4Ej3UcTJurrIIp4aqKS/MdB1CXZcqBMOcnZzfyAU8
7VGIO8U/6lLZW5iJb3G4oOCMRCWYR9jT0OC8kqyPyeG6nU+0odH6SaNJ9204vKAg
2bxUUmXE2wc3+Y7+4NDt2wd0tQJVBVPKbW1GmWWrvzQXq0l5Q/2vJz4Q/YGc3+nc
rL8huV1Z8/9nv1qB/iGR9SsEPDoaRSqoHGEjYhNT9yS8EomhSa1Ac1ZZ9NjfTA1q
kCeAWwWCyAVcGPnFNsND7tKwRWAfZs0If7ZtJQfSdN4AV14mM2lfh5cBvyp5IhVG
aEg5njvAmfFWrr9+fceZiv02Rmb/MPE/UOYMBFV8taL8ViTJ5F4mbvY5SesaJPx7
H7SiikhDMi2TCsefxpmisC1QhkfMECdsgv0a69A6E9TxFoFcDCzy/OxR9lkSJvlx
5G+MKi1QCrT7jzuSDcfBVUTXAYJHyNfi84Pbdy0aqb8UwUmLMJgtLIGmb3R2gONk
fM/iljql1zXO3DOJzDYpsgmBt8ErKJEE72QV7p4/Pk7GySpp0xpJ66XHu9zgy/9G
eR/eL9shaplYmthhD6jRS1kw/YOaVv/xk3gynCf9T+CiAr1Xj4xmBGLvMQRCsnd8
kFbPSIl77hXe4Ny6uEug07+C3Z3zofH9FpBzw5iS4iyc0b2+QoLWfRbUtPPHAkwT
YzYLpKHUC9yGY4rJvmFI6XhCEc9lTLOEgjw5AJAdLM/Jf6Zd4rAniYGhEdjFYjgU
Fw81OdNMemlVU7tcuvdAPSVxheEkwYLAMQlXcSArmCoByqLTgKQEiQcsjm2xybw+
K3efpcTJ1uOoSmEyCq15/fYJQmjCYKWsB33BWXNQIuKbLtnS/e3+nFjq7Ljs9buN
uGb7Tw6q3aGWLqy2pllao1umLVu6/UDKyZaF2cCKsESy1NHhihyDdQKwWjcEN6VE
rSFDC9q9aArI0CIwm7akQEFje+qGd8zUlVSm8Ufq5ADBo7XDaGA1JMFOcJbLXWFi
LJCfNY6IERrvMzyZohrWGt8k/pfu6OS1FeKxjF0hwIKHOPar5vyBekWdDq+7PwfY
w1oejFgy3ZaHgzMYnZMn+QpCyzpidpxor8obS7HiNzYxKMjnN+mKsA5LWABUayOC
D1mbagxIcWTxIissq/3ygcOiW+OjYfpPH4pk1yPqc6jWoZJuXTixxwrl/Baue1GP
eFrySNtvSrlyJUNFbcdEkUtFTUSO5WD+hxbi6lo+vNJotB8wKIC4x6iWQd764lx6
RNd3gBaesUBUsBLWUEg7j4hGz5y7Cy8qcehqH4fjb340w5rpRK29wSErB367utsy
agxNVHPHTKmGZgiMiIZDZhCDuupuo+WZualt0o2p+OUVbarJjDABhAyJ0smpdAF7
5EyhM3D7EDqNEh+kZVHh7EJr3eEQNGovPNAYfI0+a74AAF8pFe7gE5p3QBf0yHAf
G9HeNmb70wgUQXIGsRa5TY8Ik51wAOox/JGBjloCIJc1jjUQihEY8EnFygueJuOC
frkwbC2r1DvD96aOFNlOFV/Y3DApyIFIrOvpjMQO/NLYs4igceRHFTo8AVZ6AkvI
sGfXB5CMtVxsX6JjumH8sVJMtphMin8Pq9c22qpiYu6zgrpok0diIyDvyT5MimVZ
T5Pd1kdf4j3yG3U+DEv/JLcZJrmWXGYIhV4doW6Ra3oqxnazBCs46MtbaLwD3jKw
aWfLThbOPVMerYnkasc6UvAePGG48j2QgcZyrO+YXAu9rqh1mgeSl8A2oYBzkA7P
fQIfYVRNz9mVkhGLur7aNG7jKvZks7WLuwR2cahuKdN+lmcb3B9Ygx82QO1h+Fh2
m+eRuVqWlVeRG8nJUeKu4yAZFoZui6PiY1lfWNIJ8d+ogUZjZ1U12EiQRDvL/fW3
m3gQQUgDpynV2lrAqcrQHuclVMVsfnw2Nb9QyqEjdCGpNcZQsrTjw1k1f/6gYyuw
n+iBzmrHeKbYncFPAggWqe4NgO5wtM/NrACuzfrQUNqr5tubIb+rRuspXCyOCwsM
wlsvY1fi9cS/UwSazm76m4s5qX/YU5TArkI2uXDQyfaB5kD+AEaw9Xs03gDmX97k
Y/X0umCYERaPGkb+J28wWcIhY5XZRd17eKlABDAWF0TSKlRbLCwIw1W9tcDWWrWV
10Gp+NgH+bWrjxKenYCRX2OEHYC4WjdOMEnrbkElWVgPfII86S8m7HtTXMqLSDVV
lcjzZghO/qPLUBHA4RAQSk+dd84srk5mp0lV3siGC1t0kbh/r4hsZHrZBv791ZF5
iwo/TGbamAs7pac3ZlFWspd+vvFrlBMSo/2hf/79RraIMERQBYqEnBgiMeRZMjxt
flLELR3wbGrmaFUxVYhLh8uH+HPH+Fb8P5f5PKYL/Xana4BVrtZa1FyVytkvTH4X
AghcpKl40A/Ot+XCYIrjYQnCUqpUjehtsebK45fHfDy3x9SjPyxnagt7u68dKcNQ
22mxUKJQZ+hL5rf8QHwhfIA+dsCqlqZSKkcn/e7MRO3zJtfhMswaSk73+VgysG4r
JzthlZs86tzOZRSxHwFIdKFAjHBMx6RK/cfISMW4NJIwTksR6qLKsAT8d8vIearS
tXzyNaCwS0QWfLyb738g7EDGJbXKZ3fcRElTFit9h9/i8ak/XU2mKzEvcsf8K0XY
UtJxn4c7sgDx6U01NzI+2Z7DCOrWpo1xnOM60RXnYZ7Lbcl6CD+2eFmupDOxKA+0
PGwm7bjO+GHDyT8wJqQ0iIt7/vtl7zsSG6iOAOm3oHNszhCWYrKEyYv2qDlMYd40
bq8svvu5aqJGzdfr7A3nV1Jg6vFUF2o8zRqZXe5FtjTLWeFNjiVLRlsVcppzvntj
EzJ/HS2BAPfdzKyKF8BtUsri/t/1JMkqpaIcywBdS4zLlatj6JviAMcgi8Z5+X09
Uh7qLMcwcsaaGAb6ZIL+c+A1QX+EhJUcFT/BysSu2O99CnEru4tsl01B2FIHjGTx
jxrCsxy37UMUkNrrlGTJHBnvRKQUeQsuaGI1B+oisxP8XthP4jRV+J/WufyRKcs+
v3cxtTqFDjYo10mQK5v6C1+6VjqFpHykvRKX41W2xdXj6bdnQB/FtObhv65ruWoD
7e+ggbtFIqsgCSCsgatey7TJaLmD5LSiSsz6qxoGGBD/Yim4XWBqZrru6xv79I+Q
POfpzHVl2q5GkMpIFZoyzxQ/kcPINR2BFlhUXbg31oCb6MqKbWni8RpBn1W/0ms1
cjd10YPX+KPL6nhSnWJJRkwBkfWWFfTgaLJ2hedWunjbGJVlozIwd2n8thu8I8ck
JtyX+oRYBT09CknLJXUWB8xW8koajWeJq9CTGqE00Vq3Ha/Bwn3gzCALYupMY0bP
OpkjCZpzPLFR/MGXBD3mU+CMjAqJi9wqHNHSNTEhH9Tf81dHkU61n+aPMhWTK+h0
1frt6/Yx2rwLr0grs/icbXxuN4b84L/9zsRJ1Arvy6mYXKgDwhAlu8glmm3EDPkY
rDYI4iBgEhTldvz3ORfjmJShgooy3X8sZY4zBubl3nv4t+/ZZ3GAdAiYn82kzdNX
4jmI1wNK2nzWMQTG0UDMoULd6UBUoM73elLepsliXYQx/7BbyeBXJhWrJz8GT3dE
omLzFQYd1DBwfFxgNQ9vza3/Rfuqgsu/k/cfn8T0CJpcy7hm5Vw73Awt6v9hGLV9
3Hp0bI8Wf+TRoTE3Q0fsMu81PtAJGnINsiRKnti4XIL3XyQBIoHY4szVGILcVggb
N7IaUjWXajD0socNxLAiYntb0SaETuoE2PhwZuGB3CCqTfFW/9mDbUvdUNahFZ4C
ZKm3xhW14vsAD/bkVm88pll/LpG/KksXwLwY6vwo6QkkFjpFVf0UWd1qf23AoA9s
vErIOHMAL/mLv+HS+19SaV9VcPCOPAPVlKt7YER4r/e+nlU1bWHxE5Oq03RZyHLI
vDjrRPYfRiH6XRBHVtrovu6p11wXIKum31mr8MUWr4TdKPBXUkJEFE9KKRJJqgAf
N1Da5ccQQKD4+NPrkH1BE7fYE4upvwR7UwbtdZtRSm3vq/Od9/vdLf8C2WmZIGdS
612E9BSpSEaHZfuW8cZ7FvsmDrAx+cTcOtCAsUxr/OqfOhlrb2AMxEfPFHgP8zK+
WLZw1vnKa2pBp/OhuAiqZFiYxBafhsOpGpAfqyb/jl19PnyiGK0tD+KaAZF3C7p5
3CoPO+tS88NQobjpBrEYr1huMWK2e40zqokG6NU93p/1yudMatr4DVm0a/raMNSM
p/7FpVXa4hxAkL2JJFSusfBn9HVDdT/5CuOUx/DoHFPeudDrkAC5IhKhtbOLqZUg
7llieGUjgqn56jLwcyEz2t6rguPfUpaBgEx9F1y6uCkPp8gr5BfTUfTjFjrfbf1G
8qzEQOUK7wFhW62uF+pZZj/j+gyuCu0yw0wJrobK/r/wwUtxOruOu1Hws0E3G2gz
ziRZi0NNVfeSFD7mModHfFr9Nelrl9N1TcBz20HGE8kb1SIs1Gh0CGe2mA8+N6Gy
VKC29t+I9/X0tzNSctA5yNJUFH3lef/4LWKDTCCktIyrStmGgoRp2bRXMXgytVq+
qyZuwggmm/AVyC5XV09Knn4J4pifZ/bMt1ntN9SWD2TM+Dd+EtEQew9fYCBqWRvM
b5kjhuZrdAZtG0jBfhCdFyeSlyzpn/pL4HeJNfLgWvlxf/ApO8YZgaFVypUJuag3
oD7Exxusn/COi1boVu9Djgn/VTXJi8ck6N6uJDJfARdHFrDNv1kUFpOqMholTo1j
hgV+atRF3vJOVCBfB/hOpiq8AfnU8OgbGwubUyQR97YyHJ1LiYArjAv6dsnohKqp
H1lGKyG+8TIwVtMbjn7Z4D2Z4lIM6MMDkUvXxx6hUIdJUoYVLaCC9GSkX+uXqCkF
CVZZTY36FUfz3wMe+A7FZn9kJoZ1A6bzSWx+1TfIfGcyuLpqvnGSfj5DC/xc3IDf
RMQ36iTB1GjiwrGZ4DkogXLkMucSw4aDgWTTTT1Xfy7KEnESIddpPyB0kDNTqQ5/
YMea5EvqbCTKxeZEW/q0HFnKgu9VMn2BQbWVcI/gJn4OLvcCK649/HUkp3hzTgDp
6eNPqzFvk9+P79/Of6Wad91CEX7FsVS5ASgNQi3339YoqhO3/Kak5zuSM97BLLcE
Cf1tdxmuu1HLm6OFD7S5J47RwWr2oLaRKPyYlkmsEvp2fJx2qF8ZyaIbn8JZJwC6
DtLH2Lv376bwaj5sd3vYdhZi/OUXx3QeDToggZZhvI5Ji2HS0jQ/CCzcyqcfABY6
PWXbxV0TFBXjM7ru9HoCNJdaFwWdDipZlQ5+M/Q/4Y1exkJLbiKB1elLtd79ZIZM
Wy0rzJz6130FyTDBREHqNPaHhzU7bmoLAstbTUbBhRQTbuSSgrlmHarnUg4pMKG1
gIdfQjd3Nh+VoF9GlzAYPl7t4uuKKTz/yV1uQ5z4NXzG9lMIJx1fQS0TqDMhnWSY
1K7EgE3bAXaQG14aECP12J1u0z0tuDUBlTZs+z2c0Q1Q/3uho7dWk5P6ossoYWbv
Jw63HInTYD5uh+8hCBxhWCNsaGwVpUGnPC/PnBRDyA3XkXD21miv5KV1DHG3wOCM
JIgXoTuI32YRDgixHYlhszN78Goa3GjGRaKtZSnuDTVqBZoFungx2VoVdVJh1ikw
DpGbk1/DrQzSTEBZHIJVdmeZzZbMC14v+6xxxUEl0JT/U9g72dykMRqEdSDINKol
8y2OUPR4gugLFWVvyyNIK5UTK3zduYr5n6aceXuZreb7yCkx8VSVJ06kaAcAnCSe
qo40n1yY7jEuTuV5NH9xJOP+kjTM8J6VEX+ynwNJ/4nPeDfv1oHeFRgmHRpUPtl8
rUmm/voTc2nXkWlkjmp8t6AAxuslT7jXlz30rN6c9e6/cDZDhrdLMnFrEABCC9OD
+Sk2x1N863rlxQWZcdBz/hVesQNoi3kQpXm7dnrxS+fogDKaJa4MUuxe/EPDx6Bw
g90cMTDw9LbzKb7xtzKRz6EW0i+ngaaD7EO6QOUVO5JtPbj1D1ROkODMGVJ7Ph9j
Srgobppaz0JTuzWH/wnUGstz+i1w5p9aESsd1Ny/aMT27mBEv+i4HoHbJzI2I2U3
CTdFPTKbRs+4ZF6nb8wjhL7c2QUJ2CRSYvw0yj9sqGW2OxtuX9VdDxIx58it8pF3
VHLkXFGO2rCQbCkM9EbFVkxpgjC/2S6GBlhT4NsOYNilme5J0oz2bwzMb9W4kD2Z
fQ3xYfqOHwIy2Vqh7Yg2Xf5OrWvNpoxAg6xLzkocsbfxARlub8J4Lg6W1jJ6JexX
097VOLBmuUnGr1dwAES6m4dTVUghlwCN+OqvDkd8XN/pa7FhTWC1j9vDtMfHKvTk
JGmJbuHo9tNxb2Mqxx5Mxp8kSIHGuNdYXcasM5Vc2EQ99TcZBPSTKyJnKvoll4Tj
j+BcaZI6V8hOxWs1i44U0dywQueZg4wEGx8IKKvcq55c8OhPo0jFPGGcWjYb3XrG
utU6nvKR1yWmLMV+jyvXj+9C8xF/laQkekXmpSYmkA2eDa3+xVNNE5KaW5rg8Gia
5Cm5ikyitMErzqQi99HQN1Zn1SnkE60XDTXjdDfeD3AMZIhhwijwuXBIiRerv5WS
8rgWYa38N+4aS68sY82i+7powfe2U5SO/hIAhTZegrwBf+V0SFlK8mZxX1S0v6+g
fQd0dvBmkWrY39LfNMULhJua0V97zULjH065n/cnrnhbBnfqBGYM/3SjxKWv0uM2
nbqaDUG0Rgugr6zQqzXgaF9IPPYfwBCFaxKuHEj7MHJw4aIQ2JbZU+zoj+fqgqYn
/+YlAsgY40e6tdLzj/Hh+zTU22d91d3Y+Yml7t6fxMG+Xf82IpZDVa/r1G8/sied
dIOWNID2WtPMsfscQEB7cyUzPqM8kzHZq/TzlnIg6eiUy4PxAVm+BT6yjmwa8NYy
zayUS/34BJN2BxFzAk3iDnfmhDW/t08f8tfJcSaFEQpkgMd6Otf0Rzx7zyxJzjaw
ewJpkpWUIiAOQRDUAGCniImECUY9ieFYE/niT0RYgjLiKYaP2eGYSpcLZttVWP2+
Ak9fLFdjh+gMaZ4pFex8tUiikRrf8O1s4Mm7eoQlRpghG5tl0jxLrAOM4UJhRJZn
fk+BCRkZjxJNa4yJdmVzdeNNB322/lW72SDqBJUwQhEi+moJaAw1c3sfygtsDH7k
oyxQt50DLph3oep9fpv4qZe1GvmZjXlBP3xue3NC5whhLlcmpw7rp6J/3sLJwqbE
4855VL26sVy2AvD8GpNf9S7FeCWY+a5gvvYwmAumh7nQPwfWokwvcwMtQYTK4qOP
9Q70XNlO/ym9LmePxuUVzknYLR9xg9vdTlEWj/b1umWN+tARDmw+0VJpfXpZQlU4
fDN3COK7ePXu2maduCaz18nG7/H8pREorrAejWOJP2OLWWzi0GoARuoLbHAoCYZl
I0SYCNRcakpNc49FtzLrxD3zL3wN3t018qabIcR/ZCfC7cJDUgy1YawHfFu6fgLi
Tp2hAoyPyZuunWCgRCbdhuaqqrR4AaHx8OCwbwmNvDNGYMCh07sksxioDj0QOS+j
y1nbs0hL0T0/D8X1dsbGo6k5aAMLu/qbAl9C+4K410f+iSzr+ypK0uEVZL1eAsQ9
DMJ46qp8quI7TqLGKtn2D1YL66UMxUq7I+SVHwrVbw/0GJp81o3hbDm5WQlsuwYr
LW/tBH3aDqtAJKJaisvN+jycOz1iMFHB8yGrfVax0TJZ0arYaq33g3rV77NHhEUr
TrwR0SoT7ZE80i+7AFNhaedS/wHbaPx+9uR28Z4k08u+yMc4ODgfNF9yypGaFeJL
nAZ0QCPueuALtjvkZWr7Nf1Ch7RPp8z+AuAkfO5HJ2AcZQZDnR03gooGnUkJgD+i
ExbqVhVonKriquxV+amkjvI9ErVmRAXruyMbyoeHfCfsttMmitMLrvV+TIIPISVh
31QSoZ1DnsCfo7QA53aKun9G4YGNhDwlCrmFjTXLLigvazGDfQPY2202Bt29mmda
B+WOzbvJt7zZ4qscsJTOioKrlsnL76HkHfvJFiq3s1E03tJVpkAmOCHw/1zmM9Jy
WfstmQC0MNaLn6RG/UhRLr5nSPeDhNA2mqvN5It6rXMDqnrL2UwHP+m68evovBEg
+aztaGYzirWPzuYoL47elQnWBLkeUxI27MSZwLcgO2y9bumAaa8oOubxQuiaa7mf
M6Kra+jXbjJEmTxMD7wSH867qCRKh10omYIhHlWS+oqdqrjkafeKr7sDPTzV1Bli
Kq9BPgjLUWLNeK0kbACwVlHK5bPm9bgPUhS36pUQhoBrTp4IiU9ymbDMOgHuqSu7
DHGGzJVC8PRWxQNISF8KBYENhEPuJbJUhM4gicIny2Ifx7JRT7sZI+CLXsgTfPwC
CFAMpwmCHSUHVQyAgCxJDGYYPfzoxson52awyss3FDsBe2Os0qM8Df3GbaTw8Gay
ceIhNkBqlr2/fuQWC8B3ZNhC99S7xUpJMA4Ea28DuXLDEf9sppbYgYBJTqoqbyjC
Q/JE0vE2sQHgHtNhNVbKx0SKhfDfkQOvBcPFUBmAP+jsLnd36X42FSFbuqdiNzqj
JnymNVb3V3hpdpCNHoxNCdGA9/dk1DeOONrlJXmcA2eddAPh37gxwgiFT/bqk6pp
LHDLCjA3IGLZCL8TtZkwmkxT5iU3YuCBTYD8OVb6lp9nB9pNzvEVw6DVkcJBNATG
HPW/MZaB7BNkT+uyzlPFjMsPkDdp0idSkVQmLYa9s9Vtt4Uu1kkGHGSHnzhD8EqY
WsqOVHB8gOQsi1nEmmEf726Us9ChVeYHUphicgdt0/8GUssPXuHp8wxvNOFkryzi
E/RAXdSKuds2x/62Ig/qEPvCZEJdcRIytSt2m6n5fdQKi3O7PBKf3LN/dQkzQksR
UEp/r64/pmpOhDg9yCOETlPkxpeSWDuSq0GcIAHBkWngIL4Sb18XwieQDxVVzKgW
FXim9L+jGhQKHqZUGuWRsUjrTf88EJiQkZn5vhKLOqtIDFJfCrfudzyUG4X7OUin
bpNURpmRU5rGKorRCKIlhiJ9fDruOruGuv14I25xgJBkH3/Lk6d8rFwOq4ZAjslt
f3227y0YBPlLq+Kra8jaVweDUkvP9IAK5NoL59NQvOiHa1Mud4OQBBYzFOZjDWgV
tyjoZp1CYLZeq51HV/ruYw7i3RxJI+YTn6e4ZU7GoZVqxdKDp5bGyL1kuBzUpkOd
C6PDETxMAVRVP0X6fSq2beW0c51JfvS2+B8644kcyKEC9eMG0VG9P5G55ujb2Y9C
rmZcRr8hd20F+djtNmyeHjai9+zaYymjC9Y4mvD+A6GMGKxIjDMokhMMocCnJkrl
MOelCd2G++jLOUEh/BjvzHoxUyOcPFsTLeeXPc4/65y20P9M1wiuc3bUfR+m1LZt
YJsuuUQT6nqb8SXQONtMZthx9bN2X+5E0wy9azVgn4rmkenCUh97ZlmG8iKf3okl
0MwqQMD6Kv8SgfN/jMWRu6F/zldh+6TZN8aYdTiA4eYGlWSsydEYJvK6sbfjz7eh
Ir5/N9Agikz+ao6nw9ASIVZBwvT3eh440+VvMMV5bj03JQvHPWCAwFHd/fZpQ7/+
L3Y/6UC6Gk+rsrGXmL0uHmy0TVXpC7CpShz8dH4aZDz3T23pLqFKow3EsvE1kxVM
pyKuFbVnAKAQXdikNFaA9hbnWdGN3082zSVEohTBVvkZxiRNoZEaNQBzDdDwpNmE
UuTDwuQ18wxF2QVVtkMGCwS/4MhHNBytA3xrnC3XQ4uk2hKSK71Sf3qbCbAJPKP5
r3P96K16y8xaJ8JcRsCodonGHUvN6/EQLCig4uroW/V18Y5LWNehuQPdRfcOHE43
E7xJqwW1UOs2TgOYceQeYII9dqMacZ9hutgPYpQQSnw1Bz1jaYB/gF4agNFZIhzB
Nx/e/JOL3VCCqXmKV988bfZnIfxTadsjfkNh5Qw5SgHf+PjnWuk5ebDVYa7SQxp9
jdcHbkCDI0F99Pk/UGHEJNYxPZkJMy+gHs0DmFSbWnEBIY21BpJv/Du9tVkfzcfs
kaKITvHdYi1NZHVmaLwXoBboHeo/tqZcbZFuvrruhUBwy6A9csFMVGm6mG9k4COJ
OWC/2xCFvbbvDXHAmz27HZ4WULEQL4Im74v4XFQIRXUg2LBWxRCRoVP+tnWIkB4C
MeqX4hp5jHOs5UDpslpCMFDfGpmjM/crgQD6QcQWyHr1u1kQEqlSRJNaBdzlibR4
5zjAQEiOMGzE/Sj3VQlzrQ3mPhLjEMCiB+t1sC7DfIh3mFIjyHNNaTH0CW+envOt
oLkyS+Q8hruE4jiQZVGC0gRUN/Du5Oj82lfi51Kc9jin7NdUAi9+b27sPWxj6FRc
QmulceGJ1pweeJD+eDH+1IZ4gtdhc4CvhwbYbL1CIua8V5J2IxIZmSjhQ00XEthn
lgjndB7tkx95HJMd+4LugquJzbgWQ60ysGQ0m42Vcp3QwqgaHeCqjWY4uOs24Ihh
itXigfiuW5/teH+3S7372wG3bWl9BwYk+U0Cfkv2HcjR76+nTV6DLquqdHTOxINb
n4HFqSPnRFHoHt/+YXTHVLJq5AF+eLGrIw3fEdnRr5NUEovUs2N/+kFU/bMQw3FE
8kDhassUc+RvPghonreKjFY5nRkr3K8jMlJ0dVU6fn3WD7Q73yvyJ9IOAJ5MHLf/
7X3ujor1+fiGYveJXQExLIs0XPDzxQeOnS3f1skR6s2td0O2/G0pp8m3ho9s4QFs
NlnOWfAE2C7g3sgUeUV71rC8sU32aAk05EEgcqX8p7AWqn7R0lne9eaGw31o8GNW
xuk4bK3/ZDWhFlAd3vBLvqnsa/iqaEkZoiO7vm6bM+svIqM6Dc0i3uell++2ZIGc
RViGf6188Msg7pKvlDrfv0RfyL0WVDU2EBqmuHiMn69gaPPtUzft8eCF5p5accBI
Oh9UCrkW7qA6CUJyvCCWTrFVxUOdmZ2s1dkkJmQc7f+iX3Dwzh/e8uNMwrAiz47w
6iicHDxTaOvitsbb1uuYtad3pVEUsRYO8g+56jJSfl/hRWa+/ZGdcKqJPWeJswCG
EHf1yDwhVu6tHc/ulh1HeA8sH7Vv6wIp1LH8Zt5pOcBnma0MBb+kiimLeKK8ZRFE
kEGDPdP480Yif2FSCsoD6LUJ/gTNTzF7WX0e0F1LlcEkWVm9A2Zs3vWXwQrbhJdu
MNOvXeFg4pFOz30CaOL1/wIsKFJNkJ0wHz+zN2DGh51bKdxh2wy9tHtuTN681l19
4LPvGYQKSWXYDRNFHC929ceAhBeY7KxyvQ02d0kd3Auk9kqg6kPEwEETeL8Gg30y
1inz2xFwMFDs0SPZy9u+T7t3z+bbBQC753sIkkC3BJS+tUT/A02Dhom+/QL0B4gH
bDFxrHsNVQUZ8ZaSOmT3Z+j0ew+pJ7RmgzU5HpHsd0IsbXoQOZRRq5sUpFsQXYQF
vHXrW49cS63qccNTzTPT3PVZTtLYd3Jhg1BNC7dle/+2+6226VOHPL5di37Cc2UA
xz2qTy+AmzbFf7BrNPfWwdXjUaMvL0A/r69db1YUVCggdx8r/Be+G/02Y9hALz1p
soY15iEdrItaSsOxbkV6tAXBd0QVAJocN2ejekFrDQ/oadbaiHXqTxAo8TXupFry
KzS03FwmeWxuR4cG7SkwmuUCDEKHN1Nnx/NUuhOaD95toPpjPpg19LeT/jTkwvn2
JnNvchyhV/TOou350HhWOzF8oLI08t3iBaSTjd3L5wuoPzBEMArSSTybHX6AftYO
iHmYPiD5BoEw5+1Rw10x1TDo4K6UZVtVFuFeLBwZbk+y38z/z5qzK6R4muVGQpuN
hpLVyLfaLIotU6F82cBDYEDCMou/MYXueNIGyLMC6EjtsWDTORJbrM1JZwEjxewN
x/tYVeOquYOvsWTY2LMSRL81z5PJKlAU/rgeLqtQKkTEKcATXq6ykW9fBeoRPhNs
Qqo1wq6X+BKlewiNtI58EinedCps8OVtOszZ7+viBkhnJrMMNycPufVsIiDFO8a1
ysHk8uAG4LWObbk866i6fPQRdZOzn0DFt2GabcJpJI2dTaxB1kLGCbqryrNGmLmx
0z3vO+wMssQCubxTaAT7VwTv0rliOphHdiQWAnMc0tkyrDuEO3NRHFZBoHbHKHsB
E1m8QQ1ECNSfkbSF7Y55KKfqnldgmwp4EQywQT5OLZnyLILNUfDifiydTp3Gy+/J
BTSRVir9HXiVng3TcObER018kuhysfOTIyW7EX9WYzy0PmMHhkqFn5NSCAb7djgG
BY0k5EshKFEFMM5iGMm4xLqTb+EBoitPzwRKK5qoDFn26TnT3mnGw+ujzyzyUptb
+1RVFvoVsklXWaqATpjMB+DbqI1DZ40VLExuvNKgBDK7biadiULXaL8qPR2g+BF7
fCKekCV4LstSDQTZkkFToR7rqQNEogXKJHpdt6KgQZM+8aHerUA4KURnC0UsFKdo
j+NyW32x/2ttaczPTqKFpjj4/yz2V91CoSjFAnH2xjvEm8R/WJ4A6DYUhrIj1wLW
AKCelvK950+LIh2iI+AVeW+yj0t2A3YdPKeTwhId2W1wVV1+8spHi3gMlMSSNWZ9
d2BbJ1OOdTnDwGIs9CtrnS4YTcErR5Li4xf9BCR4JZ8JnkVbpCJu6jSgImLvq0TD
/vK+MiL1+NSLXAmIxZKvXnoE7chxC4r5cZvLCKESiDtoZvpO9idMHaSUbMBRFdlz
t0Ha2pXeZOsD9BO+DotaxCZ7ifAGOz8QBPiVVhL9KLDf5wU9/t11cGDjHENAElhY
zGXU96a1kbYsD1VziOxqMtK+oSZucwwErSBkxb4IF05p7/WV9AkMyK9osWbnMrMc
Yl0VB+JksP2LYmQB4YsR9xVgnWbDysUglG/saPicgDC5OqafKu9oJQtz2g7Oo0lE
M8K7aX9mGaMiMgAOGUL9wkwM09/IFinwuBxP8/VUjeOrUotP/2AIMOdvLhQ0ev22
w2jc8eaOAVksyP4TL/O3RsArmOIOEPwM5EQheNMHMySQFN33si42JesjPkkFe4MT
+VOO234V4vPC5NAYpjcG8pacK6OMuaetQGPuONr6RKGYC9dMnLaIicrCJi1AKZzY
PtlQ5kajLpleLc2vRh/kvyUqa01fBQsP+J7WoydWwSWXRLt5r3OEeAQYcdwzaR8T
6oxi25WPMFZ6d6wUSQ3DaicSRjgaLzJndZ821SzG6/kzH9Apt4CnAbbnqpqSf0y2
xAS4pR0r2ud6v3gkikDVHQId1weIOvG9PF1OPYONnk7kcKX6DtkCuhSqlNIWECuK
ooQWZ8boYKIpqvgp0gNDxCRHYrHOpxjcLhIavILZO72igjHxWqeYE8VxK9buSKIY
T4jUVwhuXU+Em3MFIJjfAMT1shtVLZiZnMTJ+qHaYYFQlD3y0ozIU+hcnRbpyRIo
Fhn7z1z4JxqcpQgI+A8bNahfqSof7CH1NRSaZLSCNpI9c1FxMoACyi9xKKb9VLHV
xc0Hpn0VKBQpIrjhP+XXoZ6BfIYBaMp9eq89H3LbDG8yDxGuU1eTfJRhutaTVFEZ
T665ikSXPrY396yYE7+yMEvrTN0Zw6Nslu7CYyTt8pU5HsIkgZx8vHF0QZob3cIZ
3piKhk36vT/UJKarQauQ6KUc5gwou7tKA42Mocf8XzL9Yj8RF/X6GS7wPk5b50p5
1tPD2Ne/6M/YAKZwt4RYP0cTu5HS5be3VQY9Qzbc+WWlcw3pi850sWxAlZqPqoFL
gqBbvV6o3Sd+QdhyTSxlCIHeOfF+exKFK2zFmBIbDpyg41ABpuRqnTrNR8hyxhUU
j9u51NfRHHtIxCtN8xqXB6yPoe78GpwSaZXw6il8TdqY62H7VSSZLpo0a0WHMgzD
d30/yAWKGwmzXeN58gXdfbLfuglzTyJX54TZrSqVcXhsRpKfbcmvpysCJncxpQ5e
HcAEy/bNtQ/lrH6/eZYroCOXz5MJQAM53RwMNncBzTTPos2/ujFUQzWluzLs+kJ9
x6C2BtlY7YHejbch/YDqk6Gi3dycpdblm+U7bH+FwBLy2TNB/3h971CrKCHbPgNb
wiWQXfYifWe7jxYI93WtU58vIpF4LMX0B6fh6P5PQ70VOmAsfEgKcUGAnF+s5+Vz
gcMU9OmjQrmAGDzou4gpy6rFyDGRnczhz9ozoqPkOLuWhv8U1mBvBnw01B/mwOUD
oUE6AWx2MgHPuI0QfpIhyoIzqIPLIWJCi7nbtkmdftlsL+Vp2J/xMKSQ3OjJQcW+
FVTWaR/+ZJYuS3N98zpUMCWqw0Mu2TQA9To+9t1L1FmVIGpZdc/avWaU7NYCxSXQ
i9HA3jNaNLU/iusC3Ti9mk+wzN+AeyJTHVoywnofAYOOd34ppksRa7jA5sB0lr/o
f8NQCsWa6FWsQRur5ElLPXvtydIK/5qlCxAp/SnmLRvcjtgpEXa5RyJceV4vmKFh
fGt/LXDGyjaVszn0sKaomiXFG1CHJXW9EzaP98md42g84PLGo1GdchwAXoNGuLtO
pIFvZr2MFs/mJUbrhxJakpfWbnwDkC+V1zDfEFHTFr44U/J9TQywIDWtX0k/iJlN
bw5cBumBuQWZYxR8+qw6DlVq9dHFEhDa9XArEIDIS9BsrrTyG5BJRICOfv6C9h08
Jzv/jpPpSdXvhl0QjHFO0PtrnM3rXKlPSozeEUhlDNafFggyhc4vjz6dqL5Gy+3U
Lln3LrHnkFfxjHrn1M4T/2FEgc21fIDkWjye2W1elat5uxhmw8hRBRszMmfuEweY
jmJmFq2exoSqYDJ2SJJiy2MAbSWYYdPS5cnLalZPjxYoQLvV3OAx6wpDznoCssOu
lBjEDD/I89yLVE+RJJ5wgV8PPMDcYDGCSqNgiHSRZ1VruRjU6649tH0bKUUyRF8k
o8eEhEExorxQPgSMq2jv7WSbt6PE0cS0f6XouEV19wybQRUqb8ls2hwknyekn3Yv
NkMhZuL4mBQSN9jO1R9GmxkB8k8wZ90ZF30DiSQUlbNqLr2ChSmwACUCNsq/m04G
4DPpnfLlLRX6+LwvZhhnuCQUZ5T5PML0aUis1U+10J79X/t6dayjOxobvpElPvnV
lanuTPUwyJsjF82L3V+1913oH8ZGhxqnXN28PaV6Q4wedd0CuE+udRi4dSNiyxwh
pFdObKX0Mw8i8VmVAtH5fV6TQLZ+18bfIx+FPR7SOkDmX30HtChOZdj3TlBEP1XG
Z6VcplIFLbDc7bWGIMIhEFt4u7rHcTVBEyo1808pwT4RyVI1LeirkAzGontvXpqA
hAnf6wRjnThfT9UUO9oJr+VKDNDZ3UzLE7eUSOTK20g98sSacSknCFo8BmLuBH/P
tDrHms8wyu8hNSLnpxEFVptuvFlI5dOJOG+WQcJHdaCjgkgPPTRROV+MS0MdNDHy
SV+3UZ6MV2iyfTB8AjIK0cb/pGKlz3UvK8XM7mFpggU4ML5OIxAiALWg/5IGcAgR
L+MIlfaWQ4iCEbvJCZy7cN6rrzMkGmvpPy2S8qUR7bcHYpL4vLvOnNP8I2YbCDAU
7K5pUxgJBluWyMC92WIj4QXKMTMo1CvUlIPG8jkxcu6Fnf5unyEjKTl1F/he1cBD
FbqeOajIY2VG2IH8qPEVSTEl4uwMBp4rsizffWKKXueWyJEJpSoh7dLHAJ8sAPvK
YBMWtsI+8EbNSOF+KVysPj2SS1Mc+ValYN4mWZX/FhU88gSMM7hPVt9nD7R8VbDg
EPWFleGSpNLcVAvqvwTYbH1og4mrILUy7J4+z5EJIxOrkxAYRbXBeRYU/mhaT58Q
Qz830cE84i486Anz0b2C3pkKeMwjQA1lGnFiyE1kl22jH2z52pFe8sqY49PtkJh+
E05yGp4q/PejkW3a+UBPlDfhLWpGHScJ2MhtDGhAGgt2cyh0/9AqcH290POdeQ5D
ecilJed/lhLwM8r9u3PkT6oyeZFBRPA392edgrEhneJUo0Z76SlibSL2mBhdLeBP
ZWAcfcfDWpn5Wuu7gSYDybRpLfyrK7stdCZp0Tu1LP1UwROvcgLdaElimAV0jqcL
JW0oDYf7QNT5oEB/7OuwGt39SOAtOVOZNIOMCyPKIOHqwzNOxZeiHes+Fm4jeHA9
nmfv1E+AkyoWyGJnOXEn+e5l+WK/xMLsAKzAEQM/bU06YXe8vlj6lh0vm4H9Xmg1
coD0z5QMTzK2N2Eox0mTPdf+9kcL3FejQA8qt0LjCW4L23DYZe9PCaq197MrOg4X
evJ4IVKW5tCd/pq57swqA6+cS8tYlro5DY5j0JZHCU+YJAY0tdVCku/GwjODwaWm
oe2P+AJ+1x/RnLzjDCiVBbwgcegAdlmAZMfJgyvVrG6bjaTP19qw5NnWFCPIy3C7
K32yIqqwZ0+MOWW1NbVrVaFXlmvWhHL61RKC++7XiKIgvTgwIatlyNn7Co6mKth6
2qC0tFN0pxfvCaiySC0U2x8US8UJPKo5158bER7hrqtuUEq433ifnow6Ut9/Mtzf
fbyL7xRdhaP30aUc20vOS9K7JZYzralPBmSgSijO6wxypThj/LlE/MZZi+2qIu3/
DRXdCU6P1lB08S45aWA8c1P1ZtwO+fIlH/uwPSW62KZAXhbkn0ub8W17+guCS5WE
4AEI9sSomdpzjroO9D6YcsvIJrzkV4TYOYxvdnBqpROx9Ymp18OfvQtgbC2SwEq2
NGGzqB7hSUQSehZvM1s87sDcKPkE8tRGQfJaCEntjDu+q8JXSiC9uJltYIeT4hlu
yAEv2IlruEcCvIAjZ1ICoTrZgBJAR57aYqcR6Vu8NMDkd4YLC/5I9YFQoEkyd+KN
OUyzv6SGTBAU+9zAsEisrR04YHnHHNyFvzMJzCUajo9FAQwzJ6VjmV+dqeR4hZrt
QyonYECxQ7RU0p/92uB4semfVT+6t195bYsYkTpxwU4aGeJRd0RUpcZ/gCdKJWia
4l18D2fTFVjlOpcDCLy9skbp0V+4MBOgkimRZ4EVY+hhMzj1Tv/wmkamQDKPYyGx
inPWuWPT2mmjwuP8HQvmz3xyM6S35vgYBKlvppRei33b2p54OHA+weiHzFwEW55h
1yQD8S+/xSQbuzRk3zhZh8a+hnTs3CZFbA8E3V395jw3cdLQy1SeI0BkmwAngwYu
SQG1uNhZflNMu3DuwzAPKDdanZ7wUlYizrkZqo04wbeBHg95aX1LjxuurM4NV0Hd
mcAw1bjUaiIjR9fZ07mwS8T31hPPMaapGMM01AJNsY5aoNJ1708tGmE6v/eyWWmy
oCeTZaTUGpG598dyBsit85QVesBIe+Tcq+TvLDBzTSRIqeT0BX/fVVxFbUOZ6pLn
SCAEhN6DgO6nD/Yc9WzESOV1xB8Cc3PFdNK2QRHdBdcnHLRYJ+3DhWxNX6fEZJzE
rO+ucBzULM5NdJ0wUsbkroAib4odzI7b3TN+qkMufKh3R6qCm3lGEjxSU0RpjkMZ
L4oG0hpvPYnmrtUkh8sWm6048DNZAMHFzmJmj3eX39wTcH53spmklIm1LaWXIujP
UUoLaeG15WGirlYWeeai4CFhCRWT0/nJXgGHAGRlyDmcoaFKCnuDSApg2Lxej0p9
F9jUhpMTYo/8a62RBydB1QG+z4dzZ+OgW864UEtC09Z8BBLeLpc3ZH9/G2maBdmT
/tU9Zs3CYitFqeXAtRwAbzEbAfDHJgzOd7emDLe9IGAIizEDZEjWe0Ob3JXN3sLO
1GTqZ7idT/5TlT9J2+sXf0R0nhAEoYbg8B8/gK187/OncmlMaW8EV70WiLjzp92b
M2h8Wk6SKjsfJBbQh09TWwXTz+GWObnXoJeda6nwiOQmBFYPQvgBh65Hixig/WBc
Cyi4VLSLg3WWK4NZrgokGjtBLwkoF7YiE0TypXtwW2HtWZg1ugNLRQgDHn5F24uC
Zj4hNQaZmM1BhoDjyFmRhVdipVvH2cFX4Rn7NRoh9xPCQ/10i6e8UZPFXAgCvypv
1sCobm/AvCoHjKi7x2HQzy7zgVsIeMhDkIk0DCcIr72+6VFje/aiChK1e5/NWvCR
r/yTfOAMVeCdaHqiziON3pl/Y5jfXr16b+qaVbrAgcEI+ENH/EKqXEXzpNWNmKh2
e5fliB6R80UOtFXdQrKuxJv0XK6Y3wJ0QPe3Hrywo6ZjpX77BBq9yW/0JA0juoB7
YYNfQKsvrmRJ8TdlJ/XP3JaALP9e+H6m7Lhv3xpmvYo0qTa2RRgoOdPavr+Wms+/
U7EhV6VJKhEmv2cQAj/Q2eqjW9vPRLj2A8BerYGnVpSqsM53NmaVB9mgUGWhXmi8
+sUyS6Rj60eeypC6PFZQMCwnA8nk5rxDJnH6gIqyDQ7TqCtM6DyXzj8tmY28J01N
k1wUkC02llP1emZ5GRQE41H/iocaTM5wMMNcMzyW5gUsU68CtQYC+Fiq/YIavqc+
jZvRPmgoVLwxObmyD7iRUrpBRS71a7VFvl6aGMT2W9oOuhlHwA3qtGLhHZwc8YuQ
pmdVWKEw/KtZQ3RauncdyIawEI1JLxAVctkJ3V8+OMxVKmmnwchfpFFk2G+umst+
bJhQwgvYkYbW7sBYoD+uZ2A8rDj5D8HC32EkaXO9srzEll9Ujdb5BxYTkMyrX+0L
NRHP9sffg6z4eNQLxBtyNEd0uS9HUgstNXtsPiFl62oB1V2pNpNhtX6qj8tyWpkK
htK5DrIagw2JADbBRjMgJXvPMQ+4y+Yy+7KBv4iggGNL/x5bUWJFRhCCnjXvZ+WX
p8yjwzjctPD2a5huH/lYydTghmH/Bwa8aMxQx+60NpYHhYAl0ZH6NF8cgL2GTJXe
gL5AJqlNniT2ugEMkLne9iBrb/FJIXEa2TbIpJ4brJ74CE1S2rV/4LoafJXynU5w
PcLIFs5mGa6beHSaVbosR8ugw4cPndLR7YFOi8xE0O2uOEaAEEon8dGtO9KXVe76
fFmHHikda3APh/HCuxAmJZBR7oBWykam3BZyviniesx6aKvSB86OtTJHdtnRuMLo
vbj7Bbcic3nztYWdig6p6cmmxrSEkXaA4LEcEq2S1rfpxhZLA3DJfMsbJWxnIGOb
oHlCVpJWByrjDqGk5n4nRAyuQl40qzfPws6vbsozuQEv7GUI7+zKPwIwlM2h2R+e
VbfKqb6OeayhzydFl0ZcjqvxMzS46FroETGnxrbGk8YneWPK7XggW9V/T0TvRgRm
juDk0EghVAELED/jphSo9lEAB+v7y6R2Ktnf4ksoNUuLUZw+b9ih5ylAGiUncNWD
iqH7Q+ch8JphZg5dj0tgQVJx4tefP0XBzIu+ycUw9+2HOH/hNC91n/Hmb8QFavuO
l4F4LIVBxZGvTlpSGZQOkSELrEK9YbgZ8G15r5atrPAr62s2zwDcXUk+9PxYm0dg
NWhQ20VS7BnR6lzJe+c3foBx/Yc0P9OwQ5utXH2gS0n6f8TNuDUikhPAd+DrfJXY
OugPxuHxIw0SXtZojpxLM0pQjTVkmw74z0fJlQPptfzY7kGeU30psqkVo/XBTEAQ
PN7+q0QRL/5AMxHTGQBf/YdaGql5+Weh2FuVCOhdX4ty9DcbbcpitFVHOEwtKTz9
TVelJ+nQEMRUeE26rBbqcsbg+NxJoWu/7dHXzWk2sTjt9BeqFFH+UMhi6l+k4Cbm
P5S4MdlOcwjYCITYSO1P/tm6Npugx0coQm3JRGlKpAXNPAcM1veDrsLN9uSpY9SD
+FWh9R/WCPhV8AeMy42eDtUkAU0V3qKCnWr3mjJiWkwMykr0PNT5rc4ff8LykWVa
5oU2Pv62TlXTfuXS5q433c16d6I0uNUtM1/39iEWHi9dAQ67NHTyzv+g8xFxC2e8
ePKsU52K4JmfVatrApMUYbawaRMDfx8t2E+YGEeY2/OtlDNzbwWXfV6hwuHKYg29
0epgQ2fCN5jddyVX9Jd6X4QC2IQka88kieClKZci4wnlqJfSLA3FVS+szIKeCOZf
38QliuMtEDuYc2KcBfouTEd/h7HOGurb/Jedu0o/fkOvEzhpDGwp8prPjFzvi1R3
majiMqwHDHSOaJOx479RGMhJxh4cTUK9gqvdmXBfY/KbDpHRyDxKVSeHb/HhKcZH
5ISkGrsM3OpgwrE0O5wVDrE3qI+JVtU1CuP2AUDPohgkOnjslILp7PG/5jG0qDyl
UQoVJos4G0DlkW+3ugNryOeoFdVQ8q2IOBGWWhQ3jNUVUL6Y89IDjyk8/9hTSwbH
vt9LRt56Jay1fQ26s3DDHEmClhYd/sPEcCRF9mJiMlM9vG6GaCEKeCgFylZgnfEt
m72UtkUGcH2MRUQto/p3iIpV6R+3D2FyVTqTYGGYJDtdzyFTmh9Su1r67uiDEkWE
7RArzvyPF2GckBBalhnoGKYpnvzovgQXVRr7WBO3MllK01VZcKkmdD18ARygT9p3
gsgdhrafy3iLbMYfb8weQf+Kz4WDL2ETW+2cJGSjFkAg3Hsb0djk1f5uDg09mvtS
vtewJydrrMhdDH6YmfGMfpdXuOQnGbLwJOp0fkNPWf7janY6IQqvhYC1mOO2O5hX
Y+bgV1xN6FMqCv8xMwnJxuA9207DAhTxgyalCaxpS09S7ks1TLoOWg8Ste0NNkAj
vODYIYJRCPTS3k5uoejnUmQSlQsA6/W6a2/AeKmzKL8WFZz0cWx2sBebxSqMhraA
ztPQkfGhnvv971nfCiIzR5fgW/nlkv1lp6o1blBPiDAOKSmC9m+w7/8zHDgdqFvb
fN3tPzKn6SzARSt3b+Gbihn8FxA8HE78MvheVmx/bPIM925414m3svPgD7G0rMVv
fBZkt3R1d7sQ6BiYj65MUiKyLE3X1rJaLsM01YDhr/7ondSbr7kbqChlW0xLEWs/
vnxG3YiEB+3frcDtgUxF2Z4fdaudp1PZ+bW3R2/wO7HjBmCN5HZaDm0tHaimU/Fw
zbYRoowxb/tnP0mOhaeGH5BqfPpoeS6rxJ5Oj3g4QAdICIY0lVDMW04UVFiJohnq
zj3WGWIM3bnaWGZcYCgqshDqqKtXy6y12rXSYYQm5uODlV5G3Q0NdMErL/oxXnAV
TPZrbgH7zygefQC9/KlwWJqyz7un/CfEjjXmZv4aFe7iZCJHw9dIwO+rNVdXxoNS
SE4XQ8SDP6FPsvuDyXeJTCjOxpfoDh/H6oWjmFjuaQW9/unQCSMwu1RYEdYmrS1R
5+6QI2IBTawQuxuH3tAhdwuHn8Ti1s/IKEddmoEg8xmtmbtTUjLoeoFikmAZnkL1
uHj65TW7hS8e0LkL+NxvxA9Xv6Q+uWGRX/Hy0poSFzqh6kg2q0f50ZvsqXxBKeVp
0iDIVKtkccxS4eYVukZcNvDFSdc3x3U5jJh56N1ZCrPGlkmspF+qkBqVdpcKlUfz
wyXWkx9TcLDxWDB6P9e0ScKE3gQlEZhSzRhnKix0+QYNfqkFeogtU6FEEdJrltgr
WBscrIq6v5HrwIIvz5MFFWzH4YBJ99fUwtELKvShHFW1FK3AoIl/kjE6Is++xjQQ
KsvM0UZZZT0sMbOMnelx2GORjBybK1KVax+v54lJADk2ACXse5DL3odC+TtWBIxF
/m2qXfum/bznTcCxJrJSq5Zu3Ra1zcpLRsHy9A8DaujboD4v5Iv3h2yY4LddQg7A
vf4qg6HCXZJLXUqM/qkhIObB6weNkfhEJsZV2eh9fG6QfJMZo0rKL/OtOdWZ4huT
MzLGuurLp1kku1P1Ni0WdjXu3JZOPwEqJ1yhMN/jbhU7LpVY7INfIif13HJQ+0Tb
zJvrH9m0zqwqQ5CHFsLJg35qvKjOxf9wAiIKQIqVBWAZ95yQvu3KU5KlMExegmPo
+96TVJnxWoZoWBokrMYguc9erAFuzWpy/f14aydeqqis74D22iLe773jTxyUmnGM
d02t5IHeFcGHK6ng03OzFRmSPOgv+g5on8V7B9mkLbcUqEi0ZP6/u1ecTYTv+xQj
6QormwmMQH1LrQpKSa+kROWdBjLDJF45VQ/9AF9MNCUgpGyJEtcbJog8sjnUAAkv
EULqkI1ypKnPdZU7+BLcOHqOr05rJiO50XbvIuIdZoklip7RIJEi+8rjO964ncuG
A/REmbTTlEkskB/TKu6p9YEg5Aa8zOE5g2dZxxc1qM1PeqR//A4L3vGgmZx+Z9nD
kEfy+xsX2jB2WVZ7fX44zTvSuqQAlzlZmWoaZBz2Og+qtcJLtU3ZlRELFg93VUsZ
PDJvr4+5hrUf/PqCSEUwu0h5Ic9RpipImEjQZqvrn+Vm+dYKKQzHFlqNRFi+DuUW
vA6uBAGc97yR+gW01L4csaaFu6AlHHjZGjqfzu1RWJXru7TAfN0IGyJg/ja7Pu2E
rO/vhWtc0xqEVzSWZDBO/ztMkGGTSs3mkCFBt1LEims3nFQbDnUOtEuXIziaSqq6
mRTUYa2KdjwF959SGCYjH5ApNb1mcNanKU5suOBFpgZFdTBUH1+1w4+163M6VjoI
f43G1VZjGPkQ7Q5PPMQur7BRIEFQoq6gNhWez3m3Io0Y9R0lFXPsLghHmd9+KYf/
D2Lz05R5PtMivA/hzo+oEHUQJkuO86rsYC2g9cGa/sHU/R6wG5qK67Gf2bKwMgx7
LOq6qFADxIjJCEbtCYU7fzuXmQdx9oFHY37VuKMhbDBcdpb7grT6QcS1Yw+pgtSx
MHi/4GgRyvHvQ6GPIEVw1bTXmk7Boy/vOVQp8Gx7WSBP0smKsnb1plAkGvKO8bkm
2dJ85fwfALnqg4OYV3nQmcur18Z6MvZNyiSKY4Wy/n84a0TMF9Y4eD6U0an7RJ/V
5mFKmfH3ropKGexmit8Puk9suWJEwtSKgjNRgUYlmhbTe5BQ7FzKkLXFt3/7XDCx
3RIpvpXYc9ETX0P9ON8GFcrvz6YlGx6uhvyKdTxbhIk3++M4AxavOwNhWNtHts2+
ni3PsKISxTUbk3KJnUMPWfjZKkR7+3OxRu4bWuNrsZtYxRUd6wnV23sUlrjow3Xb
Ejr+FYwn9QhDBrP3/Dzez/35Ql8wi8qCnsRGeZTENEyxGZezB+bTFJsymgXHG5QV
JFC/bhsK2U9L6NE7XJi7K9KLiuMfl2i5WQy5Qx6B2gyDkUuOCLeaUiEkx/dihxYR
E3ot4UTqFdsLJ8pPSjXcIeMnX6RYvbMUZ9zQ0l1CVhRg4UtsZi5deaSiD/30DdWZ
lHG18Xkoj6+lw487AXfCjwQXkh9G+TneNlR6JKIGPpSVwcd59JaVMFMEbknCu99E
1sgVItAP23+SW4JoTNAArEmhZXuVgOqlAhNlFoPlLMGA/1jJG/Pmsav9ILyjzKOU
g5KtFsRC1ie1ZwgP6OUdElGDVuyc6cW8B9A1DYtWVyzloe8zlsLlJMdPUWmFqegP
palYnNU6fHELAMmCgT4P63JyPDboV/QmJC0otA0Yd2P/YRNwoQZ3K/9a9u8/wwlu
ghKJcXlOEIEWht6ipUWGA+0KLQe3JUiGjL1zbkLAp0Lazq5WvgvBFxgRu2+kUNIC
Sc6rEiMg4ZjpfCLdMTyTL4A/ZzlCZt3cIqbw851oEZVyZyZFa3RJ346LHJ+UycNN
4mV8knlSF68rsyXkp0aPsYpRVgNfI5ks53DMktB5u72F65mqv9EwoXoGH9rznWxG
ss+grX5FSCnFu73bhBIW2muGKflezC+SLGVY41A7SCCtDeKzblJ6U+i0n6nAamdJ
1d3q06GkaqMk/7qIYI9Dw3Kk6voIwYoYjl1iJ1yF9NFxYWMWwPNIisJvP1yODEHB
TuDLpM3rerUbb00CLXKN90SIeRkK64B1X7D35bQxFEv7PO6U1V1+yH0eY3DXSktK
SKw42Ttj4y3dyjhjHC/kLn6U9NMZQu9CGyMZtYR0i2DSl75KezhXXUcwhJK72P7S
uTU2aQ3zMyQxYIX3zRzETtWCVpvLzgkkXs40+d34IPHmyHd4+KY8YjJF0mPxC77m
f8Vrk7l7m7nTxxFJ1Ur+Od6kozrDY9avqPvjNmaxX2+cGFBqqus/sW07YeDDaWVk
TeJGEVIAlkDGmtNPK3oWXuQjZwQz+qpz8fc4eNktbJvD97tjRsazEEYUHSyBAZwG
QupCDowc5JsLjl5tW3pVutDRchWTJBR7MMvbcH+ppR8tooNyqOD+scRo1A3eXjBX
CxoIaDXSEt/lP5LUfyzprs4294MKls+Yo3W7q/yEhMHxg0sP4Uz/ChOiCizdbUlU
R+uvW/kVJI9GlNzjKLz29FAAP1V7jtNKVRJcybeo3NOYKfBPpovYBKOXUCANGNe/
KEXwzjnxnHELhfQE6uEyTbdI4gCir4tuN9e3JOFLUmYRnHV9qgAGQ09AL95OkvVk
oW9aSsbmfwBHIz0rfHD2quTZAIL3S3/1rsRKMvGLjOlf5ANGvqS5wEB87bwU+Hg9
d3m5RmL6MxKr20lqwf4w7hK9YRB+GDliXWWfQ0zmR/72UtVCAicqWsA82o+MvPtT
zi2LArYk8MfyceEtepyfzqmNsQpCeWkWbVzM5i8fjLy8lr4MGxIsFbE18hGExLBg
FCF/bejK0JN406zTs90rvsUPc3j/uF0IvGzgknc/JeRtbCB4PbP8mEi3xmvokMz+
usGsY25kahizyigmE5rdR8d3VUopfDmFSOlvs3Lbfu7xJAc3GW2FKL3YRVw5F7tk
GjqxDeQuo7av3L+Tt/0zj0GbqVbmUm7oOSsfKcxcdYwNhbiFxuRcKitg6wV+2R7E
Dxq07wjpleDLca52SdzVb9fTO/Bgt2HOebQa/eYPwLineqyOtA7FubZQaKRM60aS
Z6tTNSXzNfwe0ZrWydGTH+gzgrKdz5RHXwpjdSEFBSgmagE2xjlqKbE27YUlqiix
/xdBbEItK/wRa1Sn/gGZvst9o3tSbBaz0vZhUZkkKvhAHW6upFLhW/FGRkAvjyCv
zzxrV0Dfl643aD30LKqB6v298k5w5cMtfp0xMtz3r0B8kZD8FBcEfU6DTFZ5MQlv
hUu3qSAbLp364NHOlLFxsDd/H95lFrKTBfb/zznnpSyVAHXrpm+v9abUDSehzaVr
EXtrFB6Ok/7g/pqQBaU1LZYMVmZe/s4naU456Gx2A0qPAPX4FY6LEB+sYn02ZI6/
BP1Ms0hD9VKe+xzD2ICbwpB5VIGVkfxjJ4h83JP3rMHWtfhR1jBpKKYxLwiv+IqE
TFM+R4ebr79/1bAau4kG66kGJX4jXB5dtlMA5913HY8RK6kvYji0p8V9DeszPmDQ
D4H56OvrFhtauxSmhiL36+6FVNk/fzhrRsV6fZyFF/6tYp79DS0a6R/QleEhmfZx
9XcIlaMisoxrsP3Kkdjmgmeb5ePrt31La95gBQ0k3J7FpL0fhBHRQ6q1GmdXcPzz
gPSEKkr4vjYQoNbiB+7iDvqFNHSuczhgEYE/qD6SUmyTq6YLCwMQw2nOP3QDAKXP
5ADsljFD+C6rlLXTmV20hOkF9nQKDlcxxZnZb+xEpucU6KN9wze6CnzBeLIwVFQo
NUKgthb+INDbexTVAVLhWlDNe7x1N9YgajcJf6gfDI+4Lac7hR5upsWTBsvMyNYT
YUon146suLuBc9Dru3dhXCUQyPLkVahGX8ypHEeDbOYDIbb1so9nggyCAj9uFlcc
4+aUWUOjI5tpFP41ynX7YnjCttyNNG68Nu+hy6mRhZzr2QlTLmgB/iKhhh5vo1f9
smtsHMxN9RLxnmra5g/A37oDqcrWy//OtT6VhD8X67vrVBK8mHl+szfbp7gmo5Xg
8cHTd/p5R+YLyrU9Wk7LJ0BFMLqVgO75MEglBOJjGYMd7x1p7OEdpBtn54/i9bzo
tMRr1LtOnSHvPZYZFKWF2MJhmgTZP4ZnHiFRWgwZKSV3EvohUdqs63vEBt4IT+Zx
ePgJ+dlawLrss8EV3N3rmuF/bV3/AdcRF7Bbaa08g//AyUTDBFeYzLqw80UsQSKT
dv8DmpIgAg3RJhwEjnHhkqYEhssbId8nxTpG7pVE352hIzGlnLJTfggCGqKQUmlk
FlWMb2nSyrDQLVg3G/8T23O0vFBEsFht/t4Ufn2sdlffZWg4AOVRN6X+RJkj+dbj
MHBMWmWEpBLPw/mN5Ep8IIQ6IsSzSK6A6ALt2GbGWVm061NiFdBRt+UJ4Z48n2SS
wZrQ7KA5oMHDuVxl2pl3h+sQyknH1HGYxRZ57NdUq8iIgWDnSIIC6H/Tr86s4gg9
RuCr1z998DarJnRzwoX2b+Y5Uf0YKE0PR1lyzLgDCHkPtmFkK0i5RiUrLgIbaCKf
UOIv2oxlS4u1c8kQYmVwObTJ2GLr+wopEO7bWq7SuUk+Alp6h/VGvZbPEp+VXK3/
yDGKEYA0c8rjgp9mr4r/RiWPsn340gDySf9avV1SwA08wUFO3nlFmhlYhgm+fYuE
lEUNvmq7b1cbYhLTN2Re0D/xmVReqULmvwV7tFhb6tJiUBZOPyq3QVOzyRVXmcT6
1kAtYhQDTx04o/c4oRgZZ2GAaQB2mj/2qmk82cNT2tnxolj3/iaiPKqTB2kuKdzM
CeticTIz7UBtrFLcMH6rTtAmRwfxP/WJVSVc5QxOWrCUreHwy6BGKeoupXgFOTeV
uRDoXkdOgSppw1OMyCWNqOoGQ0t1BZCDfoKltbqS55mot38f5qMvzLsS2NHuSEQM
gg4YMaJwEu3novbjT1VMlnvCOByJHygxF1Kcpuylfa03pPnoAZFoecOVcWukuWRf
gFSB4thEj6hDTiCZ879V9odNie7QL+BGSt9L9hUJVzeUgbFO9pwnFJuu1uNcxlvf
vmo9kAPH6p0kqDOwV6w4HW41tZ5hrN9CLk/PXdXb4o1WAirg4fifVp0bNp3j+oi4
H/YtL5mPTmfKSBxlOGqgBTCGGXsyNPiRP+TQNEL2Z8mji2N/qvspkx1G//9Rx7Kk
jcStypjumsjp9f/bIqLxLzcEvS9T+kb2Ug2c7D+YT5EE/92UBABQNO1KmpVGfeWw
NrWmOeAlIFEKyC1dtd7+crRj8lYsFhJPQBgYiNE2G8KKm6d0BHGBPwEBDoCMoV1T
x9Cg1SyIDCySGWWh1/6FHVHapeHqpfTIyqkfzOXCkviGu+rrNB3612waHd1YglwH
OJVV9igLotnP3Xm5itWtMnzzlp/n9MJfDxDd6REkZU6+ZfwYbSRE/7ChSuAXhFQJ
Oqa+Z/lwzMMuSbx001ZL0qYUO5oF1Z5wsLZxGhxVpPhDC9Eq+/DIw3FJgWiIlgqq
t7N5OjqEL7/pOYKFXjAgrzsMIgkYwfDYytWpMHxnLIMAC3LFzmxElYlEn4Q34IIO
iHv4serEVlBIgnEGNg1+nhY/JU4+Y2vsPt85yU9CkKtao9mWgydVtmny1dfgd1se
H2feNO/NKt48sO8D0kWEQAa7czqnT+oXC0Rbg5aVH/dsYGsTiLUDSaX2tWHfM5vl
tGvtygp3vesfg9UvPfiYACEfzW7cai9yEvEzasK7LMQ31YSLSn7w3uROvMtnlFga
ij6PlDu8r2bWNQRnGpfQbu9ij3dWKFq8JpAROu+mPE+EBh26znLOw1UssVMmtnyy
xqVw/+bYWb9fi9dEYD8Fly/MEjI4i4MYI/JjKJBE2sBgeP1jjUVRFxBZ/88v/M72
a7zqR8jEV1lhgLOctP3s7kt5jV5+kodkt0ewcDOr6rCCor9GcWGqAZU9jSrIku2S
klfmIgufsK0UR/DB89F1ieWlcwuQf/QgZMZEHDFtL5ph6blllMfbPdx6QOV5yUuw
gLPr5NpUK9a8QjjlCq35eMj0wDzNL9RJFu0IzSLJ81JHU3haZdKxmvExEaVZJBxd
8JM1349nlIbfREVzGsYRnw4UlYcdArCXjGZ63ZuBCeCPeHZuOihlh0xcTYxWeOgQ
uQ5WlHHGISQKKeKC0JSX+ch6Z4xMZrAfhXbKruaLDIlTh/DfRtKJD0oNF4zqgrWG
gNY9rhLlkejxDBtEPydt8USdq/bURXdQY+Yjq35L9zszpKgM+N50aoeQhRqbSefy
urw1qVQH9ua424qdbekxZ8n49Fhcfd5h/p5RE/hzB6d/xGvTkDNZB+Qp2ZwBtIjO
PcYeqLC7dXbIPVY2zi1EfZ5v2dA5fhNExsHI09wQbNhUaNRymHH3iw3jGatsCnAR
hXc7xTNBdygVrLcfCBFigAIBjyUa+kWmoX1lzItiOK9j30N/5p/t12AxV7KgZ1BW
kx6+oB9HXwu24epGiN1Mwf+Uw0KYxRb1dOGTNhnI6iub9gpZYkBKlroLGM2FEuKV
nwNNB1Tu8yCvRwKoBQ+Gz6Dj8/UDQEB+GfZ3/nIn/OuTvN72cy4y8Ce50M5Pnu+v
2jHofhGn+gAZBPRc0uK/5mYCJnOIJTCMjFTHW1j3KIUy2v2pf8CfheBsN1QQgmDh
RcJkj4dX/en8RjYT1f4uuVTRUi0Zt5qIMZN6oSem+6vi21AzW1Onmrdq+zOJSkYO
9en0FXRPifuy2Q6HFzp/KJZWT28MN9ofKh7RIuDDjnXBMPUoPQgLsnwc1OMdq7DV
lB/ox/aRPhlO3vjW7XiUxlVu3l6jc6fbHIYhj6SIRyK9kb2QKpRw0IFH1nqXZtKB
xqW3iLq6b4Hy1ZtShDW5qPEArmUNqXySNYJ0/AoaOyeT+YZkNNxyAwF9JmSVlE3V
6e000P/VfLQ4O4skAXbWHkHOZVEhmo0Q7CUWWbAc2kY2LVOKh4MrJiQNxD/fOL1d
VGgrNeTOlBhw3yn6dd5IF78aHRm1CMBf2m0blzMEU31CqCLWYKnM73JZDR+/vz4p
9yG+Oc5iXNjB1dYpqrsBbkJvl+6IS9i61VWNhttgqdoWJ7wJCc0X5KKVclswjhku
Zx/6g7mUoQQ+nohMuAn6u78XCZExpUYETU6miaMbHw//GmmqoyAOV4afmiJksxJm
4pY7NU0Uaiun3H1c2dA/8dmv6RwXnOShgUp6oHIUAM+XcSOwTFF/IO6YV8PvltWt
DxOKAFQVDtvlksgKMC2fCongnN/z6vJy9p0xuO9DXL4s4vQtOdCv7Xj3jRTwx8V9
Tib6EMtfXfAEbDC811aFIwwXbtj4fSka+3VP7HT2SurU72B2HwiAZgn9f/d7SIg/
j3Req7afchOuG3Lfr8CDia6/MuVIOjssG53qmHr6ovqDkpQrUpRzo897g5xpU8Db
zQ4/UC7CoDt6CxqNrai5FXVlfc7ythFoLwYNG77akxK9pDJ8TS/r4HMmkXo/T2+d
zj/vWXtaevKcYB97iJedPy9SZW8RSjANUBaRgMxG74N29KYkWFZfVv/JYcDJaNph
WuHYfmsNkmyQ3LKpqew9X4TXFKuD5RXX2ar4av5xGk9QiQ9b3UJGVjKEbM03yLvX
KD6EFOFyzQjoJ5WpFKaZYNSirL8Xs7Rqx8MWWtFjWs5jkfSIz6B6ea2b+/3T8uNC
lLoqo507wWf+wKoq5f/0u5sRLHpxk3VV1wkwSE98ouETbBCQNqBgcywzXTW3/GyG
oRmUeZA8Xpj/BbqxlW8vrSxkRS6LCN2qggrnAsKJVBhKJOTPtnAgnevY4fdDojgU
ygoAC6qFM3bICNzfIw13P93mNxGsVv0FvqeSk/bFErgSH+YtQL8Vqos2ml7A6YkE
SkT1X3ThzA9acqoF8f+t3U6YDsUi8GMHZsGcj6FdbEL5W5muRFiFfvllJAOhrmQb
30D1ouM8Egvce4hUgD148LGQ7umvgu1ziS6nyK6u7wtQ8VNmNbjm0Kkq2J6EIlAz
1ACq8BCXL0GCgS6erJ6qPWJ69dlFxZA/HN8IV302OAEFMOA9Uf6bRtureg14lZe9
pq/n7qdPfNdSIVI8LAKDN6L7xnKSLBjGUmk+0G5HnQAY5ELWoVWtrSb8ZK53pCGn
rIvyWLr7olzY/aSurRlWjBWTLeBDKXpyPiw/SeiqAKnWh5wl9zI+UIrqvji8BRdv
fYUAR4YP5KbXXPrmUMBx3pf61Wu6/pXYZXoeyz2U+aFiOC86/6gssVyU51LmwYLU
44PxwjFzRSKpmkrY8cswAmlci50itXmAe/5ol8Qw6fqqCHhJUe77o1McPxAz7/fb
l93YB293n+MuEGa+y4QU1cXpzd9j7btFql6pbAuPvoJ6uXBBBevHFPCPxTB8uMLW
NCZvHdwclVRhscBMTlfpjx0nDdPAEs+l6rp8A/zVqIp/LDhhpC4chtFFrdT7C/tb
GAXv9p24DnnQHdELsThdY+GgoWL0OCdTo30JyoAyDy3WJ3CHMDuqJT3gEqkb0JW2
N/1lrFRcZoAST5q+hulGNHu4kwQ2F8yTJT/jphMQC/t0Y3Y2EkVfEYtNJLIprqiw
2PcMGf5jq3jqjehrOzhHrscyHiZi8I5HCckruPsPvgN3yCwPsGoLYYhiCz/hdHL2
yeROhddiaBffXkb7+ggrdvMwR7Sh5x1O2Isn2ZiIki8sSjzJ8BUBqRJtBSrU9Y23
Q0BvHi3SvBgPVz0xXdqGJzKJd7VUnbOV6Vlebus6jzjChAyZ3+sh4H4z4fRIfurK
3UbBYOJOfLqsx8AYqUi4mWpfKG949v6z2Bv+g0M48CLZwwGXrBiHEkjhLJX10Ikn
uGan/csxshxEDgiElFZ7+BsQkIqhxJUHAxYmVp6ZBb4L4MzjFDJmxEaR9X8saOpA
olt6Ffo1+OcKVbDzYFeSFKtA4kBUpoWOTLaCfBV5YUqiwu68wYvqleGP7sUOdaqt
egMca5q9lxwdReE9uj/qw832YSx7Bwvw17VZ85Nx3S85S562PBbpZ/zsHx2q5Jcp
bY+WbkoQdY5RLOnvhUCfrf4dwxEFNb/DExl+XFjlLqszf5Wee/cE6FSdiQp9nl7O
DYfsPw1OzF/JwuyP+LOsbrSV2BPyKLMitY0jdC27Tt9j37kzDr9hZ5k4UTOjGZAy
FhAgVx19hgT6PPpqLba6O/guYqzwous+kCwey+XCEtQe66+iiUC5s7sO3eqbQv8m
YCeqOmxE+EzlUq0e0+tigJdk3nP99zUcL2sG8Z0cxy6/rExtB/WKXRQraCc01OtM
bYlJh4MMl3eunBaaukhwAmV/Wgz6xxLV4jk//MhElqjIboP5BvrtM78z89XPAvJS
g1WhWzqcVcBMGkeLkNfkzJ/0+8S8zxpTudEP6+51reaOEfxm8lF71XPIkGT/WAZB
kcaf7LE6W/nGbGAQQXWd9+M5jeIJjvSzBsydLhEhtzHvmMg+vVfD0ANI/PwEXIhy
SWdJV3weQA4FcyGVE/6qV1VT9aBd5cqFX3Wyjw/YMOPpnmYIR1U4O7sKp7qFokeS
CBQ+GfzM02JRmO4e8mYdR/bEZwbeVsGWr76Jm7+yWGH+yrGjZ/yeoaUbjpL1OD1+
rr8ALL0S7u3IMc86s//95jgeoQQ7xQoBXnaWK7KZhNM4V3sRF58hAvoOpJDKHYY5
OqM8Iyg/dQT0kXOKtLEpimce3opbewydwINSk/1ijmdCWQzrb6RHog4xq0GAT46f
ljUzKHefPRdhpYph0UkLbi+Kvx1lpHJWzKIFqlCYyyHb95d96VEKcSaZqPWhbZFW
EYKEZAUGsqKJ/tcUtxT0MDMRtTlUHZFWHbi6KYCd6SWGZlx6lfcWR1aKRr81fQ/Y
GxPTsRNejSzxiYsohbGU4IJjgl9O4qACrY1s9egIfiPAMubZLF0W3wPJcT8QRrxy
lUD4Zar61aFkgNmg2HO6VvoO9qzPrNkBwZAQG5IegW7vSWo2xgD3k8ucuE0IQob/
8rRI7n5Aus1WxgEljRJI3vgOB7EAz9x+Gp33nnX5qcSfbk2mSNa1KQRrRn86a3Uz
C2/PvCiKbSLblVDXQVFL5m2aPkNIp+k7vLF5nAvYkhPlpuHe8FwC7PUZOrrNje7g
pVcmCk5Irz/K4eE3dySXSi6g7miDF9bDt65e8ZSvUR0qVQuEM32B54BxZqsc/BfA
VByx703qUlVFGGN8PQQ5gdoH7G9fVauKCVZ0njVV5ZFQ9XmO2sF1dbRPsErt3szq
Cl6V84INqYv/CXm/41tbH732K5o18NTRCRmexxUpQDywjTKFgLCN5m3zi1Nt7lHb
zoAUrxAUcRsRlMAbzokbTbc8M95Qt3CnttotHh6MREari98WBaYgXDHGfF3pcHHt
nhvLg8JItXi7TYIPPo2vwGn6RXnPJMpH85xe1G9Ywei0plAQ2+FhQlC7v57un/3M
qwTW/WiyhvaYPMdSBVrgTFizRNZ7e/eR/FuFYA4Of4+EoZk6+8a6p6VUK21yfgKU
GeHIhNJDjqwJgQzfg60kGDZhFlWCqImQzXOcJvkloInzESaDUH4BefsGdsOU/73w
a1GccUfzgsrs2Ln5R2o1A82C45cFvZMJ+Vd8Gk65BQu3xcoRo1dt3KKz/MJZ+yDu
sWxRhoqVGgSh2rXzmSMJpR5+u8YnM2AFSKe1O40F5FxMxsg1S82r9eGYujCL0LyV
ckjMlxN+UQsASt4rfovWPAhg+6KWLfIpaXmuwcCRjrhRqz2Gjkrwmi3z0hiIfnJw
ETrjJNuHzZQ+4lnUJtGPWZvvoGJiaWpT8ZXQtNUDKThpdjbV9CZboft7s2ARN6xs
fC9txLFPHpn3xX9efKRBUBdxbi2SZcykh20XZzycvo3GuCau7RiV2n5uPtf0+Exo
CbsgTtfUX3+hx6OfCBp+7x2AOEVlC3G0/vVplhcty7b3GIduMDVhSGb0pNwdTkyU
zwLtgob32566OxrUSh3AuMJs4rUqMT647KV/tdcLNjiymhJBevj5HCtRQRC+dIPF
oqQS3tyEaLcNMaMpgsyXaXTDhvo+M/UfQN56W2q7jwFX7TfVcqlEHvKqtQDuqdMD
k9jaChtSs9w2+or7Ih9cWxGFSkSksLGR1GwOMTEuxzkKzMH22TyDvh0ge8+MLiF+
AjiHja0+uBS2nwAWWgv2j+uZ37u5DsyRle9Lpp//VjlTN0YbZ0lzBQhDpc+/JbP0
x02dgnHX6S2V9tjHHjY75iApcwky3WV4LBknDEEXUPDUiaK+yRcNZDkJMbfDAkF6
gVDiTXZd8iNO8xW3/+PgvSf1EF/pqqW6ujXuxk8FmTsERVq4e+kELlvMb2nTHhv1
kUYyV6mIj9jqm42dNMCR2r/mxTX9UpRQBEMGTywVXpy+qv6OF7Ewp4lvvEKB19Ew
kwbHBBpH+hsNiaEa/J5dEA61M9oCh39FIHWj6AFtVO8eNO7MbMqak7dXMS4J/ajU
nYOKeOk8uEHdIW+VmtmmDpTRmvjRI+U2XwuDH2gRh6+DWHJL117gQY1l3uiCC6pJ
djPSiASSypikgjUkp1kbu/Meg0h+fU24zsta8gYMUwZxkGUEomlJLUmg7U7QF6+D
J1YiyKmDETczwM+DNvMBEqkYhtKEvzc4iruF9dZO53QYUbwLKnbZPSWxhZvszVbu
zHq+B09arlatK//lHTZwyfMqgydRDoOKxWNa08ShTnoBdv5ZqPu0EHvB0GBkfGqI
2yH86bk0vyK3a1fXFfZH7fcvtD8E31kuZ062R/wlBjyUGoMTVBhsL+f/4FtqXGq7
jGVQ6B96CXhUfN/DcEm3I/J6dVErHrlr5fYUQI+B3PEWjZFGk8tG1mL6eSVlZ3yG
b3Cw5jtUR+We1rnRbCBpq7eN6FT8aub9NJYEjlEGuKP5SEVA0wlHUL5W2lXwM92l
+D1kiH/8Bcw13fvA1QZVigIvqqbY7pGB1agi+sIRowkzsOLDpCxdZDrfDVRx45YB
1ppshrNQNsRTFdvFOtN4Z6oWmfh+RI08ThFfg34BI+X9Lq+r9xY8mjQRp5uGVgaY
T9IXbMppe1heBHnGfDYidUdN/O8d5ngBGhCkA7jdhA/FZ2QzNCI2JqjGpJCIngdU
AjbncHNvMCoFxOBkgDpbsHWIpt1rBG1unK77ZKuPSOZJnJO4u320gCV7q1lgsqml
Tcd0qQAxVslRFT4W8BGqOdg60tpn1elUrQAZtSTq39Rm3n42JVDU1FSggOG/HxoB
Txy7kcxVzoIrVRKkl0FI2mGcLH3q2ulAuECyIYWD8YiWeypu43yPA0hjzdb+Cem5
E3tEtoFocfhXY0uT0ME8KH33PenxU635qgemSDrVg/WibdbjmMxw2dG0wJ07smdW
OqdtmZd5LzLCq4fRTTcRpAxjNpB4Th+iavdAijJYKAmngVzhRWyfzWX/8K+zdoNs
ZvTZo/YrFtpOJQ+OgUEGHHa18s4l4Y7emUto2HC+rYMgCKNLyOo/IzA8EkAuRV2k
JkFW/akDl39A5jSXZ9QbavTQn1dvOOBHus6Go0nYegveSXnauwbilAsdwmf4qSTt
xfVAQ5Vpv8trQ1wL2VLSe3nXHNkiOIV63Go4GDgo+rVodpBuKy4minfpOlyKowUj
BK8INN4vI33nsQb6d3xebMe9rh3h6QN5rnwB4tah5bhI3ICuh5ypaZrwUAD81Xtz
KwOQN98F0vxdN2uWUE9hAeaCzS+2f2sOJFaZ9kNSPGLuN/BsuOLNcoOZxaw7p3A/
me+Hf2fv/35EHux9qDck5mb2dEkUj28jpdFZ+vyPxliDmWni49AZ2ZBTX/DHxpKj
YErm3MeABtMGnDdXwpSRgUwjS4Y1nKAc/xmVrxJrBr0+Wh10OQ61yuVCDAvdaimm
AZF2Uim9gnfxUS2aQZt14D4FV3KcWVkcPx/QkA/4ddDfCRaXFr/FYDh35iOeKwTn
A+9tcYFL3vP+wJxG4SDHeNLsEND7BYO2vwBw9wC2NF0ejfbt/G1SDKkVyLI1Sfd/
BXpVzpAvpi8x9Zd2XWpSfOnBZ/LGZEqe29w3XZjF8ZmYzhn6BRQKVClifOJXS0OD
vr8QWU3S3oIEMIlfYKsQeFcj4Sak1Kb8P0QS24ywFEyCLhd/OCb+cq0mVGYuDFJV
iMp3W9tCCm3jqZzX+eiQeHnn0mx8Fpzj2fvv8fHtf5shnt7LdQ+QrGNJ+FTWhRS1
TWLwU+iZAJYH2Eo8lYMb4y+CnejJMKJb37wICKCSAIhHPvRfbryzWKHS/K+6gYA2
vecxzFiL9ZNURcAnZ+XtDEkgcDnXkvSJQ4mmtCz5QB1n8dMBjvjokFyL2y9wcISR
lbnYO8pqqpKCyEC+u1PJG27S/MV7VZ62BhxboOfiUatl6RjT6V0bvUmDFRpXyg3+
1JmGf7nzdUUJHtQYG7hGc7Q8K2eePBC3dEIX6ahysCZ6DByEaqUCClZp8g9mixax
Y35SPD1EGa3yTtZKhg6V9yn1pw8tj4AS8UyFtq/0XfiTdQiox/g0znvwjYmSdOrs
80HJCkXzA2RoNWIH5PhOyDsHvNaJZRW9Y69Fm9ABmzu66NXBc1AGRdMlOPi7NGrf
DrljjT7ZeCrodaxCgFr++r3bb13SXfjlocmoXJRLkkiKgkWcdsUtNBGjqg4RjMpY
uDUPqiV6bjMGjjPNs44KvaY+omyp3mkN6eRIAJwy9qXp1EkiIh5btGBeqpBFXlxV
zeWuRzBc1G3ko3JUZMxiTVahXbcRzfbl+wFAq0wwSu1UYlnQ1EF0FoYr75Ema7b4
tVKJEK1RLFRrK75VwiYJAWZIQyg+6Umdj+i8S7hKvAyb136jQN/Q4vZWL9Bk9RB8
0oWhBE5GUtxm8EI+xKG4/L7vp8lSkNCYweQs+0ytLziirP+MKliMlOBQYS26j/d4
/ChYdPyZKe3uahpaMCi0FW3V6GdZAqqgzVlC5r3qYa3IUAo6C6kJlNBg/2r0+sOx
bu3tclUu/aXYf3i0gaWEipJnlS5tgrfUFrzx1eoSfVILVZwQWdsZzBTssBmrD0XA
Bvq8nvnKEdUiuCg5Yu+ewP66yCGPzDAKusZrN1Iqlfhbz/W1lfMbwu4qqFF7oIa4
8SJbQsAAralzdHng5XfnU3o2/s2z2py2e6J3qRd/ljNFHUF5mljFHxsxddwNfqj2
BS60AVRs1S57e/CFAFkykxPH8jsIQjL0Z3ozAelQuaPaL8e9vOCRfnB40uo4vp9e
nhG0jn4NQdLWemqCOE/XZaBhRSrOPYUpHFSL+iv1iVZWuyWiDCAZklis0hBgWIwC
Mx0fHDisGz+Xf20LkggDMjJY8UPEhV/4lMuhcJ6RvDwJOYoS05izmoFijekN7zV+
8DfsqT++GL4qaMWdZTxh6I3YCa0U1jdzdzE7vECmLFJ/0TlI5RuKC7qkPkwyPlEP
qAUyJ8S3U0KOF2iWD39PMg27uvHiXd/EFXLrJ2q9vwfeR2n+aomGjuo4RX1h4Nt1
JSG+jGB6YYq26BzIVn0cPYxpXydMgU/qxR4geJFh3FEcDRgqZ2FZZtXGgXlymSP7
Nf689NYGsh1OagrAq/RjY1ehndgFX9NnUhjZrzZy3ctbSyewuv/78nuNYiJZaBKj
XGayMcGWAk5TtM0LGxLfVKaHgphqUqRsCegHuRvsFhcFYuGPyYFs0S8ZcRm3vW+J
3pW5tfaXpUm7IchP2nT3olyeULBPc622ZGgNnHbt4Je40OBqarHl7NI0fDxBk/P1
nwaL1SLPddGpDylIKv+A+/88q0bKT2onYaKcPtEB079zEaCn6Jx+cqAJ1vqyEy+q
J4jpvwgRoUfJ/DDSFuWlURWfuL05+gHkWxst2DsXPHU55V4FYjB9Perkd94LQLwZ
SJIt5K8B7ZyG7TVAWE5I7PiZmq1FN0ZJBKechQ+gMR4E5dq8FLvflyyfeGWVPJcp
cgJJ6MV12+zuduxl7KgwHysO4Vv1gPCh1DMS5qI33X1hWXqjNTLUYiV9Lr17UgR2
3dQPPwVR+Ps1uVauYVY9OjYXpMcqVZjm6yHVOtf+a/1DymWVbWuSbNxwIcJ22XnJ
bOzSa7PY8N2Zx1uJLvBeRvyQhnf+ZVCNwqmEFlCn+CHyc/Kubwp8xNMeYqY/iVEa
qZXlgpbcHKmxGUostTm/qI9WrhioaOrwaBmLkNwqmMTJfbZHHWegrGZvq9kUoQs9
H5bLsELvln+oFdGKCsINtll6Op9qiVFg22mZcgM7FeYGj7jY9/7QlAnpSLMbIr2G
aMSkBTdc7pFWX4vtLOV9Ts+sr/n9kUfpMnyQADrm3hyI0285lPAwUGdpa13RPG6d
89KvPKBd8GPjAhSKxGLcawd/LzrPiPd8/AX6G38tBNOI5zaER2sngGxBxuPipqAY
oRpupkM+PUjk7B7ybc0ELYptrxYpRpsQKhveSI6Y3kR0NJtW2OLLnQhP/Bfv+GG0
5EU5FMYCCpSp8uh94+9cYylJ+aEtVfAb8vuBZZWTgylkv0rw+iDdEL69RPuAAl4o
hBMhajqEkt2AbssI5XosMuOQzM6RNG3jq/nll5pnnU38QPwOSI3WMi4zwrKeCEyY
U6QLZCV+inuYAZ0jaaYCcCcgYqN8pOmwXv60NGfmaVnjtYEg9XHr1M1sSogBypkx
z3zArlOzST4N46dUEDeoCQFV0XBGI+O8X4J9cY7TSx+nZ4PQW778W9vzPnJs3tUr
+E62DINbNvJnY9yRKcqXSZTKsuOZpbJQV7c99CyMvCb61oEvXE05vr/j+OgzbCCK
+RbwhMYfKPWLKe0e5pQ+skxH85FtWlegtMxdoQdGXVXBFzxbeifPXKwOHFu00hcs
EgH1TQBcKeNndhjDeXyTYIDTG/QsNdQVQcrdVKAGIB38K8pZuimr1UgPbcI+FHZb
KBZccIoHCGKp5ZuIy52KzlKwizZgzu23+HhUuHtLV7+h3lshV9CmC27UHEJyqKcT
fXfTuog5RShhC835Mb9Ab3JeVBlb32H6o0m93nSJTp5IItDFjwpLEByC5T0BDql0
A7i5uOeKfe8oA1Gi/nKmOezauK+O3AHMaLDgScQ89PrujUzDLbT0msGYFXvGEFkf
NB3wZwlQxY8pEZOchnZ4n/MBlwHHtvmzOApWIaPyaUkx81nPnX3k63P2RhZSh5vG
U9OsYqzyVZYiG0kLSSQeTQclVBaIAGMBufdEZTT6qPUzva79EaoTNp5vNZqDblSW
7k9BsNV9WMw3L7VVPljyex5Nd7CEvYz3uVDH7Q8znCswcI40YwVFa8psRzlG/Cc7
khGCcy3j4nV7CnvhsZyBO819FC3P5R1KEhM5gHl2TZW8DL4ff+OG/1A/01Sugv1x
WmHHAbLFe6/yKis9d0f/oiaAHy310e5ZlClZ4jcjpRkpM2v7wmqmO+mZWpiNOYJD
E+/dvH1HdldQxHLPutmV2EpphrbJ1gT3iyEKpRIR+DcBxAIX7f2uIg9TURfyV/+x
VyZ39UQj+SFKBpsINeG5SbpE4r9XA80ehMGgxkeGOcFl0mwafiDrKX2sfYNFApu4
6oz6bCHp44ZGcDpDp2c9grxFjzE5sGd620cjn4UiQojEn7Q+3eaDBRC9d0uZY/2M
scFCXiMOa0EYv2cUWciSv+U1mDdkwF6azprX+ZYjJWnpmiRh6gYJM9fiA//b7+Ck
5a0M3PSUDFoafqbaWlXjfH7IrPr2R+RYGzMTW7ufv3V/Umwy2atpXePZ5B/vtxLY
GzV6sY7u20ZxAHZmcPP5fd80UFCuUCPdaRNtlyBb1dg2vV8Bg21GeryAaGkUi/LX
TTuRLYJ2nLPa6LhIW86ObQf79mySIZ8Bqub5d9fMFgu4BQXeB1Niu5GV9rbWVgYp
Jqon0JMbXr1Tx3TqKX7GtKTh384HM8Lp7jvIyTobFm6OKe2j2Z0SNGt1/tp1H81j
JAHb5drTYy5xq/LL53r645hkUHMz5iAaIReHos0MgRondSfNov0ojAPMjVyymmWA
i+whIcHTmcGfNEhwJ7SkkkiytNT04NEddpidsE6yG/gUHAjMHU5+QxwfGh5S1r84
TBG4zwk7o4haoRqL6ze6rDs5cmGdYA9xMDq9EeoDhfs/OTu81paCC57yzNK3NrfO
tIJ8Pj2DL+b1KHFPD6msoFs6aTRA3JLeUa1ZAqgt2HZ2bHtbIAEDgiqjxBCM+2Wy
C7ayd6AFmonmWE7avsr/3dgEfTb85CElrSDhGcHC9Om7BnCxRL16jOfvpttxWbzw
jANrMKydj3zQ/JgIVinCSpKYZxvoh9fUMv7q4oniRTVlqvXgNfdmhtJYjN1ngVAr
snHUtbz2+Fl0xfhv+Fv6cog927/KbY9ueh2Pybv4/+IpgS+DdWmafKcxaMIKemfI
dTkRI2J+IMWc3CKEuw3SuG0rzJgIUCbOXqQhjFl65UQgjOVd1wjb7FidN+24qTVr
M7Wg0LETxC8hV3ldG+cpAEwJte244+nNjt1RRkUOpeTtBJuiZ9EpIFaGq+vW/As3
ehMH9BNOu3YwddR2Ogp4NmpW4g7Js5NOk+RTZX49tG2iM7+CwD4OEwgl8qGVupLY
0qvPCklhOpjwNmfaqt8sjtMhkTCww5fENdXHROfdj/dsXAcW+XRpTDbtgNh4r4cI
QziOOHlZZw4nbrNCA5XVHyie4yaqBXyiEyyhZHnrZbLc7MducV0aD/Tm7UC7rwK6
u30DyAWJTH8xHp1lWBuDmhX3Ix3eyhw8cc9K6CjIGmXhKiVh8z2W5LhNDSs1ELVx
AOvVZvxlWfrtSGe4fKrET2dkuxh5JzG5+iK3vLBSqgQ556lHVFHX7Bu6II3S1bFV
tfN4HLan2X65u1TcpSe7qFsBnmpFr5K1hAIz0al2irgwdFcNv5becxWb7YxuLT/j
dsZFq/Y7jYoKj+Dxv85m+qjJugGOeIAhpyHrHUTRicmR8arEgaVVS0xngDXdW4ka
bLt9+Q4wKqLRhPBWfvc9kg2dl1mWVTs37069KRu+haS7c0nsGonoTLAPE1XN4C4Z
UnxIODQFozEGvuZ/zv3gqpCJDX3ilB9lG/qsUtJV3rdOxxqEcJuCy++rpVuqFecf
uqT2+acCOxOWL6nnRzCt4K05Z2Ek8PIIBWwd9ldlxOgan2/RrbUUGiPR6iiZUh+S
+D+aa6ketfAH3RpANJJH8ZMGK8wH/8ST9fxrlcdyA9K8hT2jQUqMy4TPrdC6VHYN
Oo56Tn/jLPQMQn5gvohVlXBp0BPJUeHybHyk0B0AdDOT7UvBFWj/YvOfxkNuYhzs
A3xLKcrumggMsHc+lzcyG9hW1yGoVgE+P5gjhqFihjasqOqzmqeieYn/hK0kLYEB
R0S2Mv9y6E53IavT8BJB9OEF8mbE0RrbzSF38zrL8Hrxghgl+9a2AqRVYtVZyb+j
DzlVPi3AtLIr1v4ntgILyYWK/0ZQNvwsI6odAa+QC5eu14Bx8hlB6B7mSylqL3ei
il1a8q1S9QC18OuUJBHdxsuGZTYdRHVXEZSGVr5iEoSd18MfDxeNKhSfb8JLlsBO
58MWnVnUuz0wLgGZ9E7vfpl+QJ4XFJ8zs8IQ8d7nGn6e0hoQ7PLTGLdM5NWrujiu
gtSg/OgGLm1JqifNvX5sOHaqk2KiHwohks/tdyp30veih1pzENdI0M2PjFElwkJi
bE6Jar0uSN9+2DAvbjQ9aHV1YuGA38SXV1cXYCMz3eNyldGkGrCv2SF2vYeHngWw
JAT2NZA6LXsUNMRgAM2PCHTAQLrywx8xsPXTKN8110HSkmz/jXwwH5MjVqBIHSEx
2yFKbMevYX5DrBIutIYJpYzYG824juPlPHLS+sskC2/byoCmoq7kyN+LQa24q3B4
j5dfuxmaiydGyn/brF24kAtRB9pKbcXMrvKkwZEx0EEyOlHE01eLqiQ7oVmrfEhu
61z8qkd3k/4c0xdsIs5B0/GwK0C5nyD5u1xkhrmSQI+DWRi7eFok1MJJGVeGE0jP
zXk47SJo0SWvfxuNEb7rXObKesmi37jAXLyQD12iwwG2+2lxsYLIpJDNldw6j4sy
94SkCj8zlv3s11gL2hArUTjwscMjwcIkvA5fAvWA3WQYEFTkMpZu4NUxN0iSwYHT
8TDgXt8BsR5ShnGe9rG9ZpYIWDwOdOzcq1Q96WnhctJ6U427uyR2gbU0N/dxDY56
Ua8CaMVqvRbtQi6cxUIaspVqa1tAhqwzJo5NsuRw5rRCcOMriG71IBSv18Qqx+0I
da3Fgth1gBHwKLOfuYnqnFbSuDDIa7Pb8E43FLnpRsv3BlvLRYao6BGhG+Fotfe8
2Kh1vPEeJjm0pO4/XjD4kOd0Hs+TwgYmugBtjvXRkqIDrn731x0iqw1/obgRaP0L
OJsrKlPtgMCRD1NcXhPpT4uanehYpfTM0hD2tSzxZBiLl9/71NZ9oH5rgAzcovjm
/W9F1qzokQt3GfmfV0okJJQBIZPVvchq+annLycw6y0gdjzRPHHhVfNQp+iCcexu
9PLVo74s2bvZDOa41Gd1Ud2eT18aDj0iQzOaoWoUFMw4Y+9AXW4rcs6Nr3pE6t8f
mLHgBzQ1+THLCUpbvtq7F4eKKryWAovcNROJuWypxrAuJjNfqdrBI3Q2glcxkFmj
3whOwW0v1J0hKCQM9r5Gr9IrdoF5apQHBERSahTZB8mmSS1I7C7P98+DCp/dVh+C
5RFTYUj326PabRVATFCnWIaRr48Dosp10mDa3tkS7kef5zjt+YOXTf3LJ3UDjTdw
Wdc8y9Es3paq78FnSCwSc+8G9KZeQYJKx6zQqpWfEpxK+O1ds+5aO69zzbTANvVX
aPmKdTK/z6U+LE7nCjPXZ8GtfLpaaFTaWUu/kj2ZmmhlOtLrY18oqndhztYlgGi8
fiZxIXNPNJ1WtDSujhDqJrKhZMIUtefjwMGr9BfZ/54nAylQmlb6hLhpFfbQPvxD
E+AFKlkJt+0RiKIJkmCvJekCll8G8ZupxGborg9HtSixVoUCARgCI+0baLgi9E6H
JWXHyqDmxpvH0Yv5/40bGhSHCjnY8CSrI2d2mB4DLQ/54sxzCe4x62jo/Bl2f1K8
yRRaS9mYfACIUUiyXsSFoqlxa/6Bz8t8eI6aj0td2vyIip+z1jKNvJjN31LvVuzj
8ccQVKc6bEDdJ1i5FJ6LuJFroMKlkxniKxmX5yIMt1cbzbUvL2rsgqoyeqDLfSyB
/eCrgzfSoeVjVaaIj5whzZvsGvWY6PK6P6pQEZ9yt9pNJ49911h3lpPy66qgD+No
5m4MGhiL9kU7MfB32UfXnCfmD1rzda27ZFk6zn6FHdjQ8xbCwNhfFPHDQOBepY02
G6yFyIP8p9+Eg8jz9bnnZSttMAuDm1PpIUM4+/SNko/yahBj8YpJf2OW6lNXCHZX
clR1CkkyF7yawzLLn8ZEedQt4CYCjPo87+w0U9liLtxP5TgyRtr58YaTVTx+Z7On
RTm5uCjSvU3lTHCx5YHZTo1hHO1pjaEr+hvHwjv4+fI+xJ5fk34m+BaGLozY24nY
jebA83JmYxiCN9s0o/RMAJti0+sx8GOzknLflbknq9pVplNpHUgOoNdaXGkB17XR
mnQCxbOCXIcJjsa+jS1sfmlXmqFa0mldULjaZnABQHDef3DQSHRMPW4WQDhZDFwY
nrJy567/YJ8EZWD0fX71/f2Ewvs3DjqKUurlNA/p/XpbNrfoshX7lZXzgUyfm2Ai
jscBFZaRAAA3xqAt7I9Peuvhc3/vbO0wSdrmLnI8sfA/OrHTGya/Ab9x4TXCR7Mu
hTeRfeLCoBDK81WbMLPhJeigYqk7PUnsZzSMv9zif9IERydgBWE/ifFd6+kUH2PI
VdpCwWJvhQ2gZjTb/MwpGkhN4MfWComOIxUF4YJd5Wd1JprNF/VIa1h/stx8zPoI
633giCC6f/UgiiocVlbDhfOrEBuxPGBdubxPQ7SRSjLl05u3kouLLiILJt8E1wmQ
qKWo204/sl6rLXbDLTArEqkh3hFNZ0AQeta2xboYDkfSs1IW4e6w+lc88NJzYg7e
Rl//rvgZ2xUIWgvvVbI2a9RWnRzFjk4sZzpzJgVCEqxxSzCTGHNKUEMrSbjE2+bh
Oaim84Codl4ZR1/VcBweEI0NKIkFlhSrqLBfXSQGq1BpBl5ufDmWAuZZIENnrmuP
W5pheBZfnKmaY699HSeiy0R87ea9DrtwdCrOxbaZo012MIE1BEANp/eBZU2E4N2h
ev6RX/UTe3Q0NgvWgzROt84AVR15sWK/HTTopHxTWX8F9eU17sTNz7PXQJ6PFhWt
SP8Md2ySSKzMnkYBb++KeIgtBnuXS1TpOmuMI0LCruc2LeXtAj0ae8TBeZ9xZO/f
NgWYy6aAgdmH3WbexwqHEfYW15z3wZ+98bF1Qv7aJuw9Yz98+4/oFKkbJb0EY7FN
fMnfMLaaIzNK60rxatrqskyR9uqNGn3PDOjY1bDFLEtbBLzFNSf0S5pZvGEekTFB
WNK0G/GMkkUrDcIsboYq1jIj8rQcVh74imytQcokYbJd7bV3rDP2DuhUjjP5V09M
+MHWWDh+lvKXcFpsp1j+QLbRZzC17KNh9jaGxT18hUo+0z5nY2aq44u9nP0pj0Pp
YtsQVOPnKhO9EjC2IXmGMTnp11ztaUM12IWq6NHNY56kj0pcfLiUH/gIxGnUhJFa
kPOhSvoGagqcLOycG1dDDOlTSXCW1rg0Knov1CSWmG2abDFpWQCEG576KoJeuYFv
jeKJJLY1YNscsRQX5HR0RVFrMV/uh6b5Z+h5PcV1xeYcAeCyZVG+nI4QfvVUSTic
iBF8dEhk/31rWjL6yvmIKCowcABgKNJd+e/wO3Pp9ANgtmJjfE/Cb/kH0YMFSqer
kex9A4IVhBkDSfrhFy58cWaehlATY6lR1T0ZAhe+UFD2zaCjY+GwoBMXG3jYngEL
Try54AifjwyHUCBDTh/llr3liujSec3rbS1v3AoDeiEetKRdt119TLx3r0yTg+CV
0wUom4JXuRdkXcz6ortOmZz1r1idTjwmI/Mjyo9sXPY7ndpiWTfMK6Qu87Fep6T+
gFL7Wi05owToiolew/PnoKnaduce4HoiNisKEpMw5LSmTeAYDLerlpzbusDILBko
ZHR909swab8fMe5G3OZh12+i8ttyqrzzm+igWyZ3gInU/c176+KdkmG3Zv69o0Oq
xKtv6VYWfq+M0Gq0exqJqnBdGKcjlPLzIOkwHagLWdd6Y02C1ewlry+NdCnCnWip
eoPAAYb+oi84B1PLRdYorJqkigu7X1p/9Ymbx5mSX4GfnWf17BgNeMXQiXP1vpe0
44SjwTl88bcJpmxRV5G/rmhCkgUmi/rIfF7DnqY/+FDSLUJovBk0CRshpJz0b2tR
8JXFlL35A+uhNsEyxURsPhGcwRoAveoPH0ykDv5yMhgbzDp+HiW7qrflVlJ5qMXx
4SWkQOQ0jePED6j5Rk35ID2GMaf+NWMND0/F4Li9MqX/nWxElpJVPJI+RG+ZLolD
K7fY/3RwqsXKOmzJxOCD2vSy2md+yiDTVZ0ZvP7vZC2Druh4h2PuyyRYixrs8xT5
Qgga3Mv+rVUIeokexz/l2QC0aC3QGitEb6nkKoKNPwLrtfbOD+ScH3VI5APpi+2h
FQtKc2cglARPRiS5iWz/PHsx1zaYGCsZ4CJg+XrvvUSjhSClhAKz2pX+wTRKxX+G
plYZZxeAkm9B37xjNBxiNVDMcKZ9vhq58I7opPR8q0TLxbTHgxRsvBChXHBWkNNQ
fJCf8SCUTXVgTizKMIj38WCG6AmXoEYRzpq+6g160R/QTmg+1EDO8xh3bjTiwH+W
Ws6i+9O/f2ymLnMnBahNgBZtXYPF/l2CMD7coAy+ZtjmTTtrFhfJaNlUOqJVDHmh
t6za5OTqyWmtkEe0eTilSq9zkSqy8vhXJYTf+ySj5gix/zP/2Qimh5I2NZ9aVNy6
t400T3T0UFTmA4KN4AcuKyIl8J2A/UfUzHAwJV0WN2LGFRzokYsGX59nwt47ZVFC
U0Smps9nliTd6FJz72ydt+uVzRYB8l5ImFgEHmy5JIQNCbbm3ChhUE5JHEtOzxx5
oxreCBB9msnO/68t3Y3CYAsZSPeT58dvra6JcsTgxu5nRB5P8dM19wXxZK1kA06s
luiLugqpS01iAmkJt/Yuv98hc4ZznGW7zNrbyk4Ha6sMGfxTLdALMKu5Y1O7In9J
JJrPOuFbp65h3AIyttzIbdtwz/AlktW9FiYCx8uE6TNVtAbf+xg/ISxXtyJ0upal
8jfc6IhRqEehJBku11ImBHpr5pe01c9c4Tf764lWus++HFa7Weci+6fH2/v8kXWW
0JkL0yigBUKxAGVtLcAZB/9WrJu1/SUVPoW7BYcqheo397wIZsX+HHgNs6tZF5wF
0Qd6xH6ibrtJeDUlBJrnP+08BSqF8HQlEusZxTofsmOcYpkj48W0iXuHZzdmn/f+
lJNlshMGx50mIbZ14LUjsSV41NNF/l3RbqI++oQr4avwJi6m0WNxrcy+k7SIsIg2
ayDz+3LPLO6aGii5YG96dQJfN8eXIF5V0cDDPvXMlShbTH+HVyED8zuHx359albw
4hZoQcsCgZfkn6KLlP0aXskzQy8YIE9YU2/rd8gh4N6A47CsTYf/k7zBqH+UAIBC
XYXQq8Xmv3WYE6Bc8ITFWwQh06mL1XufgIDmXVumjXek7QK0PDx48dH3gcL5z+E1
yuT75pEpzG/I2k54nxBOY7J0vHHGlLFkqaAwxDw2NK2ZmV+dCuLqVx0Hc/T8YQEk
GAwZ57UJV9baQakJKtaZ2pGtB4rniboISbiMhqwm7YYdnWnYiwiqHsByg7ZWBBFn
62ZjlllBIxqwqCidEV8C2Db3E4+OLszOx9RTkXHY01E+SqO5LS0reKUui5a6kRAu
UykYb4YwqYtwkwDdfRUiiVafh30Bq3SaY7tJOeV5GZ7d61YU/eEByH7Xtmn3cNNL
y27+CV3Oq92EJgzh9KQKdYRfFB60xMg7NQDyGd17YsUUJPTAy8nBbHX08hqg0KuD
5uaTzAoKpK09N6QVknzzXg9GegJ5VwYudSMshR9+zCHBWWBqU6FKd6uaaDLPRWUa
1ZXzHKiSrnkwUYEZpZ2nJmKvumSOOpxPoom1cRqSWbwJas0MK9BAm3X4K8xnORi9
UNe63o/ZjlLyfAncVDiaibX1H6tJB7WO97J8MtI++f8hDlML4FgzEWifnuf25FEb
WJrqW/7AqvwFPOysvRBMR3juQ4QWgQ4idPDQR2xGzeo1nW4q3C5PUrInYeyAlqPX
1VLg3acTWmQtx78AQ59ATxyJrmX9SYe44K3f2FYK5VKpbb0VcBsdZGjnrnjKSuTn
wX26g0UO7yNL1nHoleNagjrXibyS4OX7RGSzgbhOcgM9MPJiuYU3UZzfX8d6tqfS
vZIkPxn5VyDgmkO5LgO5jiWriywV1B5qWuE44v/dt3jS7CKKnlBzH7YaS1Nex7Nk
XKPTuwa8//wVCvJMVSVOuk68fCjGDEyg5oumxQmbuMdx6XgJuj88RgATXFX8KPN7
nX3/y6O2CHX1Oi5hUQbvBvp48C08fLwg1Njh3yHEN3dstlxg1y2cK65M0fIX2GS2
D0MCC6vDLpgNXTZO+cNN0nBdGLuxO2HOeKfLry2C+ISRH4jXZaXjz03RKTNf4dyH
Xv2LGDPLl6jOASeNhS7q4o5eihZaPEgRZ3PvCd3teUHFwIfQXtCD3s5Dh41tpyjB
IlDEfGrzQyhmUKv9Vpr6BP+2tJrPDEWfdUL6TFFqeHnMZlVvPK2AuKjeZwmJZFjb
+3xR77IR0hzsge73+xx+PSaAF3Wf0r71lkSzEANhsmAetEUhOywDVotYjMyJYWpM
5mTP8jghByKDqRpTxprzJM3R107npCbPRl8iNE6FdA53aL5E+7eT95pJRveMNuFF
Lu9uwfXC+AaiErJ3drUDntPRBSpHQ7tLEoQyNq1aVCkQF6DJ14GjJXKefGUP65Qo
fbBPZX5NugtWfafdqnmmJ5KXLByLEcSeCHnvdtc2m51k18poOxISvo/fP5tOeitf
LqbMkzpTGeBV4YCIQHZVxGGwXRJ0sDl0pHSRQaI+VYkEO1oHMpEuE5kbgPAkEOuh
3L1eoVerkKlUV5FU9FRMHf9NedtS0fzREqAYZSoZoyh5CXtF1Wf7/JXK0M97pmNl
wR9n2uSn4uAjOoCjVSCTpnRXaK3thaAn1/mcfNXgUiQHZj0AVSMlGUW1DObUAh45
fSu7rIQtOu5dsz/nyYt5LzY9mx+8opyrUelx/QOjA7x1PvZFR4I2d1hW4bTa3Mw/
RJhHrp/fblrokHzI6uSNSHUtzXK/ZkeeNvEkPtiDhQxtWv+RCrM0QdwC6uxNb2YN
KtPYiEncwxLxwMV2arJPNXHsLrwe0rOMSL0XrAYMjF02i7MAJvDzHVChItArSR4Q
vO9CaY8mifb0pWPzZ1JYdxAqQ3kyVtOeb7j0MZQA1EUk8U3I1EE9prclC0VfdlEz
xbIdxf5dPzmarPbjVjeea+CSr1aBchs5hyBWOQYPDX2rAhQ3AWWn7GQW5we/Ylcd
6DuVzPfAEf3MiCdbhGSEBdVHgbxnWVw8pFDJjixm6p/2KqcuB8U/scBpDLSXwnt5
gD+5oHGcGSfX118+orYj0SRLdcvEDXNEK4407oM6cke1F2iWga6MZQLN5Yx7ij/o
jNSEIlKYPESRl/zp30s09UPPqhpALUi1Ci5k95Tpchs2wLYHNoNYoxan6RCbyjfP
jIjoigDnRm5ayb38XZjWf0XGj9BimMHbb5zgZbbflgNUPWAw2hTfnbWlc6wTYVTZ
jPcG9c4CWuGZBjwci1ntwgBt+tVuWdlgRsPazT2zBaI339PuyOPO00HVc/rcQGNq
sWrpHLC7I/D/If1QIp3YwtdXik4S+z/cldYrx8h901Gj2x3bNc7WJin2KJQmIlAt
J6OC5JWUPZXwuA75ES1z3DRXI6S2hGHL9iKgMH/aWE4lI2CMC03Ck20pPfNm+Hf1
WPJyex8+VPFMEjsUb7J92JolKRColnyMEEt5TM4ZFLQTbtPiP1ZvnhVzE4EJG9+q
y3XMHVojiK1Jcg2wag+nu3VU0pIMKiQe3qvzUv/t4bbsKye++rx04OXB80UIFF+/
s/F678QH/vmznhU6e7QLNV7CAQbvkMQ44MW7JwQ0P+dkMGdSb4nROxm6Ad2Iqpea
s90rbdrhSAIted23hAx6J/ZjsQfHYb3TXFu8oLF6KSPjB+jO6BHV47Dokuv+rb1e
eQwyPkqd/a/b+w9BtHmb8PmrqXlft91yXdm/ZaPdO3+YloS1bZMEnr702UPE0QM2
rbntGp616Tgy6LHq8xoqwX7kj0PGLd9SNe8Y4VyCD9vvmRWS/+AXgbqCRhZT+2ym
LR0c44E1oDMVjUqhgivjmUzH3OjJFqJ6YlQJeDLp5GtdIO3Xe2upmTOjOsvyvunf
FNu3sWQ+Le5AGGF2ugfuLrMaqNhoh8redM+dgjA9V1DHi22OxCcrRA0jwa6t1NiK
xMve6uDuoaGTcs7Xqb9SM6Itzdjt6/nGncFEsi4Y1yOGT5YKEmMuCAeXyeNE1xGy
HeNqevl1pZzeagPa4yisL69+aL6Nt3Qwg0QAU1fkTZdrkkY1ceiFQc6PXvhVWxxd
9og7Ixw2RnP/9w9M411ZjqdrB2kfcdJTO3Bd90+ZdVCPgywoNJjHzHXHzhLgtxZZ
VPNdCwW8OC43QcAOhwk9BCvIWvj2+kgnJIvIg8o6Q8VKwKZ2uqFWuyE14VbLRNuv
acps5HUAHMPExcHTHgGeG+NdarVaFZxXcZzOjYWNLCZasgoA2paN4JWqxQniZu2p
KJvMKgc7JvmcpqhDAJu4OeKuA3/1Pd3qHbL4X5cbm1wzhk5Lx1UrHhHR1joSRVBv
kM57dLDIq1yVgPtTxIeBxEhgo19hpT/HQv+AgfLS8M2QxBa/KNbMwRQpsUG/V4gT
6QWvYO9IH6Vlih2AYwoDQI63KLxWssO0LnpqoEKywUvsRuahpB9T/d4xorLBTqmY
lH3Lfv3d9qrdMZOYntVV7RkrrcAdb4R+lsbW2kfcl+JUnzGNYyWOZiPnKEXbDcEc
lxBA8zEBNsHmk3VzBQhjTdcPnt5NGLGoCbp2SVyIWMM91IcHlHfJYFxFlC7qnc9x
3gveOh8ZBdZGl0lw/FawFPad05mtJ5MLIW+iswqmxd+qEf155s9rC/O1b+OhRoEt
j7UHmas9YgIBzjE60I+479rYtR1Siatu4EZi7ySVphYQQt6pao52r0drnhhHB0zw
vQFHuWBLL5qp+gWGvlyDwJMuaJcehnaA6PZYTfwT2g1pPaaayBjrgsKjL4w3xsHo
rvz6o3QwVth/iOBgy28Fnl7hhX5kkrYFFW29hR2rPFTtbq/swwhHoUumSXyrkj0q
wEH5BHBs6T12K6l9NeZfD1qN1uFZ/mL83vqAv5mVkjrbsHQcholhOp2j10/ct+mb
+vVjpAl90kgzphi2yPJxtrzbD79PeZjngtjTUIsPFL4Y48ISEJgQYZ5e9srKribj
rKFUEaxiMVDGcwvbNTAmacADuNMvYFBuZ6xyL95H7TSXTrpwvltAZuXafmCB+GRT
bZ1CmlSuygsuRVd8UYHvZeUhokA6HTWu8K6gLoZaUCEfgfZYvUAB0uoomC5Lz3xO
JKi4R7JchB6imSypqLIdfHPa0L6vlbA6HD/2vQ9mUdgdajLDRTGEbyP2lqVXzY5D
OA2aCosteaCdn9zBTxfQxPG8yBig3zWeX92jy0xkm8EvLfpifg7wguyXbJQAJtdX
wtxThXOicOCdgu1UH/tG0pnDBHoemboHJVTWH101b2NB5gIldWNsZlnROgzmGOJx
PT/Ga4yW3Y8S7bzjpquDpOzmrRkyCTWeEjW0TTrifotVvzH3T1Vd9IMT0WM4fv1t
PFSNM4d2SZZef4Fz+zT92+waHZ7JgEFAjHuHsr8snS72qElKEvdnTzX0ZFU1BX0P
PTzR+RALSCvj7VZwqQ4WNKGPXvBdi8BmTuDD6M26LbG8W/rq9jth31AZvnf7mJ5a
h6ZU8GuSZWdL1KEzeZodDoZ4JMbnzm5LrKb7qELvT6HGVhjMDV0+JeZex7zIUOUZ
SD/tRjdTfkGXEmIQDejlLJbg+ptXzWF+uZWhrZkC9v1Dt0PrGNAXPxR+nfivjDFl
L4BinbCbWBJHG6w4iyIZzKNo2chviR/KRgM6Nn7OrHK1J8yY4ZNFEWQhW6jPEk4R
qZQ06CWFzn9YXKtYA34XrE2kuCsP8jpWOy02Iqcjn8TL+8XMTjcjaWEYqiM/3GcY
S2Iio7GgSPRMqP+Iene3Z4qCJWiBn08oOGNLdzTLcUGqD59sQEc44Vx07aTQttLL
l8v4az0v1K3jLyH7qb1rLl0E4cwM8ZZjh3okfo/iOlUI81ijSS+zXhOOPItwPhVU
i6fAIJQ+hMx3cZDo4KVfVtLnx4bkpMNg89cVj89H+/4BhQs1QS4xEoyjy07t/d1z
0AAb2BPSx6kuDCx8jJk1glI02qIM5d9OnH4Z9WZ9JKFN0LioyLTzWNL6gx67vbtB
vor/nBmr6zXUKGBB9Z8aAQkWvaDbs6niFqdAbCPltneLEQXeXLHaxrB3TjcknZGE
vWHdEQWc8eUBn535Iat8hfG+UC0geTuKo0NY+00e/GqBmsxPWf+WyqtjNzX7Ot0C
6WMbel7XjGglotcWcAcTMz5IdlU64mVU8jChCuuBQCi0eBydwXjqU9O1JFxMEyb/
Y6UnBjyaiZBtUi9VfatcvgOJrUCXWwzNRp7z/Q2oMHxxJXCbCzXs+m6C/XzVue/k
z/o1F14s2S2RdBJiJzXVxr1YW6qB8HpTdxyekdNzAEyzuS86bj5OXd96nVUZh7R0
xiCUG2c4wTRhKlhtVZqA/MsHedTm8kswi7JTa/b2Sm8pOzviXHHL7lrWgj7rZB9Y
mGgIgBLgZlU/aRcq2AAeH35DUfKhrwI1r1Wl3rAYzd5XZmg/6FL3vZDmWCUhHsYx
UQps4ODHOTVjs8FvcTAYLzg/NgIt8PCuliA1hq+hzscnBoOvBTO6Hb4gpi5FcroW
5+1/NKqOK0M4ywCgSfD+C4wJR3Zb75DMvQ2lY1gfakFKeVZbc0xzW1E7SDLrBNio
7ab6m52L0+bOimk+xYhF0w+V90FxtNBegJw3Pwg0BvjrcQ8mWxe/B4z5vcVcYS9n
VEJoRrKjB7dgIZKbjRO/hAUjQG6okiFC77lqCneBDjWk104j9a/lZTKzV8cNjviG
C/t65UAh6LGUATGQDREYdVv/DUJrFBARWjxJbrF9D6wxB8B+tY9b4IXGVHUtfUgC
xd/ljfdGUikLUODtsc6tTA0KhjXf4siFqZ4SDUbRUrGq1gNJqKfG/a0W1jvpIBvs
bIvWVsBTfAmwd0ORHMCckb+mzFRLTIbWyAcX8iBlc4w2150hy6ssBi2m5Y+7aN5d
vinexsdVYDItcIa8iz/EtkPvAF+ZV6NMeKGIzFguWzItqf9JqJsScYdn9L2OB0IS
+SHPbB8cOyfSxwlRTirpXnvC6Zu/Dm4GFsIYnsUAP45nNMaevqcZQsanT6jmEW/V
TOAmWKPRgFXr6CrzpFVAA6E3E0br5ywg9oM9yXzYH0q3v0tf7RHW/oO7QDIusGn1
n2caQQbe/ZqBu+fgKFIsJ+g5Tv2rYSpPFEuzOOsn0LmMF+CIRj9V3IkdS8xZBE9E
KPDU3uvtGujLoLZQxz3EKSBy9PmAeMbawTeIz+KXNYtJpjw06NOO5ky+r0dEW3P9
CfUjbY0ID89c1OZiBN0PtVyATuPl+MfJEzjExTJPr6uBQ5xqgLNqLjusQWKOVvNy
OZoNyit+qpdCdsRYhIQ6NfSS075uhkiqjXQzbuASGM/6NnMDPRwoF634ESe86YDR
kHzoELCjwZp7da5LB3i3vn/qE5mobN6FQtCspPIuNGOjvp5Nix3AyAAa4bi9089m
0jzVqtHCEvywaDbU+hOu17M1v7svf5OAvajga5N9ov1pjG4RmuTkir3IrjIcPrwN
GXYqtTrIQfjvfRqSmYOuXPflsUEx9q5AvOqQlxAR1udMhfUAcA/5rsiXEvvwrSMI
GLmIqAnw0diNtN5t9rFSPoJSL49E9B7xlrwZ+0713A+Ft0t+mCVPvXyRZcxPm8MT
qTJgakyqpU0XKT1ofHJrwXaWyvAuVhwFP00i5//uHOkabqrDjbMmyOi/NkVMLGmN
LdTWU0p3YtVOCvMLsew7yGIYeY141l6OwiwOlehw6ogOSIECpUgo2YnydRltPJPq
bYQbW2Hz3KzkDo/CXsUnd/wx87MiaaCmkUGThbXA95Dg8ENFDFH6VaE9Y/nQufkb
QFJV2DSeeA01V05lFEXkVep7G/ix7RgqFeslsVzIlj+8AxQBX8PopiXzyjsfkcXi
1zxtqw3hPF+iuodS7CpS+KWEuntKlLydAy5pqYu1OAXZz6JRStn+M3qxfFqXCkP+
F4m4YOE1mOOSkhUZAo3sW6JaoibTvKMjP8OcVQeaSZupdyIttTijivd/H9sKCQm5
IR1YcMKn5bIyAD8kNRThDRbLe1jbQzT26tcpXk9CfASQAfm0/MuQasJviaeN4aNi
hazIUNX7ItvXVDOggrQMiQkJNI5S7US0MUUeSEDudcTUhLTRz10QoCX67NQLf/fK
81uFcPZABhTR7BmquLB9DW+HW2guFf+tM251eTA0RGdnmTm5gTDF5MxAtThg73qi
O7I5HcQEvhMVSRR1hY9Xzdn0J+kTMohGY+wqNXAgV6jDErJ5QKHTBxk8QFzTB2ZV
mxNb782tO6C0HnruqEy7q4t/rhtkVZJuDVYefZ/6mSIMvIh0tsKhiWVtIVH7B/T7
DukNOi+ydw+7dRj199m/rIQBfg8QwUVH9NAuW1kkJ1mQkCgg+ZkvP3049OPTC0lS
cb4kgzS8MO6AzRPRdgohohQ90Zc4v9T7gJiNMHIm7ocrJXsJd2+MZ5UoqrnLJEA7
1k3EmsRwvFy2JYMenn2i6Hi1x/OWbEzvuaxSygygYHH4lJK9buCLPaMu+MHiR9Oa
as25cZXG7l/O+jCXGnrJGtQpJifjC51jnqpi33fpIIoLByIIPEEW8qBvT1QjLCka
ag+OzrJG6mGSwTuxtIn4CD0IONz6d2+jOPoEd0u5Og+Akzb1DvVmf98CTGwAHsIb
h2AkVHqbXHkP+dNSp+QgUEba4FPOsjR89KSBu1ur+LrPqi11nIhlwHHFt4EzHZX0
pUvD4zr4AqpYBZahyJLefO6d1By8YJW9T5XWLpJXd776xeG1c7FhbQC7O2+MAIyD
9L1AOorJRyyTcByi/bN4Jmin35E0iu6ZQJh8TC+HgDMjlO+tU6SJtep8MpV31VmG
SSjEwjEFcFL8Kc2PZ26dXV+ON/+Yb3Uc69u4s/sgL7LRYWGNBFiDCe/oIYhBvttb
/mKRBtQfjH1nPru0zRdcqN6+EYEWpa6ONu5gIsULgBVaFXThqk+g5IhDq8EjoWNM
X5WEBL/5Sxg8jDh6U1n8lXygtrzJMSqkd2U2hYraPukCN5F052Qv4Tp7F3ZYBOVz
HrlRBrAS9sO5b1ghKRkwL2Zy6K1PodxkUQ4olpUHbE6u5czh/DL1RC3UA8z22wex
D9svFqT+Ayfg6d06rixXhd3T6C/DFEoe9cOfs7OWzroko63dSd7CPMjFjft6R12c
A4ZyMmdcImV0OKj7LzpNXG8Y8qti62YECvz3u/un+giBrAd9ctNM/3EBOnjiKuyB
Qee+ayzIyEyiYv7jHKB9kEBreBnlmnclNJycSON4dy23IZbDpyWocYIzX8AHR5Uk
791BvXMg39GsFqYOmLtPZLT4ADxdZLQujq0OZaBoTIuGeBD9j8DoBQShnBN4tedF
UWiv83rqAWCvcnSVW7a7eeyLvI6bLfiVrx8Ed7jt47XSeXfM+r672NhX8w31Vv2h
esJDw5eBymMuf9VBXVVfA0hzOYvwvPhTqmHGt6CGl4aQWaVtzPi97twbyenYTgiR
ZJncfhFUm5cugETXdd8YfSrMRLJYLs3HK/efwAeSyuUIr4qOf6amWGDZHCySUGoM
JU6VVhFzets0QR+iZtVKnL2C84SSEBjmJhnXOYdLiaW66lvJH5XSOl4vnrBni5nB
ouXX2cwIaguZu4J3GEZINc1HAr5wRhgzn6pHgWxpjgRpR/PIJ0b3qKQ6yJgaSGgN
zhQCH8S8FR0HM+V/hrW4Me5iEd6ajrhQ3YFiFlLqEJNUqwiXrNQzpvo0hNky20/K
YzEC8X7QLBhEh20+jzZ628x8nS3BTxGzb8rvhnIisvKlXWwzs1Z08n3ooPPxhzj9
YBND8zhfTTVFHz/w3I4fFbvhHqP00OFCndAF7hVMY7h1e4yhsr1Pbokp+vBk7HFZ
tyA6TiJASuCwpk16UTP39DdBe72KmhN83wRVNV3DB8lemC1S9z1spqXEFv51CotL
hXulIIRbT04MDP+vc5XGs4vjEmIJAzkC7qsFbcrbKVEiWvAzE5+DkcI9NCXGR4lr
ji1Daf0f+pbZ0r1MBrjZ/64FojlyHNxp/xUZMUJcDwhFEgntGqWy2bdIS+On2bJG
8q/5U3fYVD3Ar40th7G4kaPtqsSTDK24YC/cMsdb1E+WOg9FIVM3ZTs0d1WDTmTC
otoB+IWgZljKeekPO8DXgqF3EBIt60S2LMpMjZPUHI7CXrbLqtkdBs4vLDYpuQTj
GMhqvN53KClexHnZs/7iBoId/DdOTDS/jm6H95Fxn5surJohfGIWTvotZcBa2D6r
vptE9PrXfd2SUuZCzD3luRzjm02CJs+VC26mJCo05Xi1sixdbAcMNDimPveTKGC1
yufXVOjSxQQOkdGeolaOmG45JcZIIXTJGrUfEK8NY7J073GgqaE5+IwV2G28rvjf
MtUBtm/QMl7k/OpUcUeE9/Mzgki24eLdDZsJo/f8jG13YK6MijTeb7QGLggkZ9hv
M+fMa56fHfve3MyJSLqFXcSz273S7FJ30wsycxZ4UC29Q0TdclXwhtuMaiSyGkTz
W5kMQfp99Pvj3V4Dsdsr38pTEZqw6LG76dbsRyNKMeH8uOo7gYt5vMITtpjSxOd1
hWx07kSRUFH9A/FsvFSp6U1VNrrGq/Npkhw3e3JOv7XYRxtJhYVEXaSeCtIKriw5
VBcmC4clN+8unUYaNVqgP3DWxa0Md5V1gmqdR9XFIgRYHSHqOYYbPaw4BSPSH89G
rmLhixyFjvR1TXLkAs6mSqvEI6O2s2paH2dAWjAOpi2GZVc6MLBLYudFW2jnUHd1
VrB0x/OfAPlHIU/l4rO94UqoWrnXceIqUevrFF7ukFFws+GxTD+02+tghh6ywsym
I/QSRv/NkL+deASk18+6AUJfKoH+aRCO/pMDVnqUSK2tWfes9EiSMsVDC851bbg2
fsPiXgThBdqi0sJnK41izh+EL6YuSW1srKbKBn3v6aLuCAifeWgA6LiF1q3J5k0K
Mi1DCq3tdrPcK5cHfBs+iwK4aQiuOIE/BUwXrUBz54KLo78sEDdnkwhV1BLbe8VO
Me6TP2saRiYuvj44gDUTtjPUI/zUwLRQV4Cj+KaOy8Ga/pEFqGYLLQ6mFUkLQkEt
oSe3FBHHxQXLEcis01j0RJONjQmY67zm/OFykGUgOXn/HNPlEYz/S3wE4kTXKVZN
n6YqcAvUQ/X+Cj6HHXGiBGi/z8N4WJ8JzlD5l2hLSCE6vVy88SGdtalnIxaBqkuN
rfbBNmWY69UAeH2nbk878dpTkRkf8ylXG58bPsS4b31ZFUOsPUaCycJkZdeE47Ay
ETLTD++HYnP0WkiDk+6/EEnVljaL4MOhj6Fy2eoTYotk22++RW9H70dklHK1KWEw
VNqKcUZ4cdgbw9ggLA6HirQYQ787+CcKqZIk9Bb97QOAZk+8kjeiqEcHeQ42cpne
Dkq9qdw4tamWxvHLv48NpW7bSJku5DATsEqqdd1hs8vwjvIRcSNJ3h7iioRjGmBp
Qi7AKz4S6paxAlUPYt1MXclODuUvjJvLLatQURXZyLQk19aIrZEl/i8E0bXVTYEX
at1t60CmWXY2NUUdGd1aBwfRil0OxmESyP7cwZyES14i53yyX48Hayo7nQWO+vI/
d8YumvZ3KyWRZ6QjUMttFRvCmZ7CpOXMj/+ppUn/QKgTHw1lOE76+D4F7ea2XneX
Oq1oJkWbFeFDK7E5nslUrEqQUHixHTaLH63BBrivC9HaqmyVzeaDI55+J574ukp+
XDK6zl0Fqfjs6eXGiRCfhoB0AsIvdhnlZ6T8hhe5TXW7Lv4gT4x4x0sLDIHiTLjw
iiduu7Lss8XkQPFjo2a5I2xIe6gN2trHPTe8avgk6Ac2RmrZLebWxn/Ob6xr8nGF
POIxbovSRslyU5Pc4QVMwCW2XHeqzKJycLoBwaQh4eF55lp8y7rbUSiU0zfmh60S
kw8uL1S6WBN5xAD0gQnBFLlI4cWMCV2AVSs5++GqQU3Ok8hMk9iXxBAY4TNZNj7P
ICcHLvHy0r6FWdYkYYdRn9JT2ZXkHsRujV7bJAnX7VtMRHLNQki7/HiesVO0IGdm
Nfy2D3amE4/56n6cpm5cssCcVpcN0j5hqjcf39JpYqxLyslBh7zuN9NhKMasTojr
+xTRRnC+3P42MmxqNSUrVkFMtELH8MT+a1ZH64MArrZjTSNib6q+MLTDVIKvecJz
YyOf/KJub2CMQC3fqEiSJ/XgPdkj+iwudgLHYEf10BkW5tZ8Pw8Dht0STi8waTD+
94urOC92VozJe0FAf4O/cyh72nC3d0SHLLReHh2HHlNjAUgCwCPFExU5AWTGpV4A
H+E2QxvyDl8O5zbGPeE1IZfyJmt1bThCOPi6XZuepG3FDPEukOwH6vbdJWAR5X2O
UHvmM4cipIMRXJAv3p5lwQdINcmrnt+AIlqljsvcMMMy9a6RhhZ/39MMBnEnbHVG
PDXrGQgcNBhqmcQ3/583xw0tU0Z0V1hfcX2HzyrV41xNRe/X0gvVjJX7QXO3onhI
4M9FEjMMRwMrvNuP9jcjSLasvcyBgR/+wkONNI8k9uPkoUnOwotiaXSAXS8GG/UZ
tOdRs5gBVLAPu0RM2Ehjc9MH5T5RJLJlJt//iSCbEFkxjJwcpZX3mZKyUr/d2o9v
pLFOI2opiW0+phOr3TR5PGskSJY8OHEuBmIMhc53MseuSzYmqFf4nGbe4G9993kI
Ug1DOCYRhE3ZVLOsjX+OzJxel3bZruOVF8uEiMRWYDSDdKFC1XqQ/Txox85bnxno
xnOu38el6+39GoWgUQRUz33ZmyuwoQUvshFQIklSIAiYTcqbKYYHh9GzkHKWCvp7
QfeKKpNqBnyZrzkZo8dAS0BQT4seNVVvzrG3Ngienj5BCzcvtiPnPFnd4qrDI/v8
s36RGj6QaNYQNfLUK0eduyZ1QBnK2F1oGSpk8WmZ2872fu/31MDoODP85rIrd8K1
EHz9+fUkmEkd+CtJCWomEUcPnvObxMTpYy9RzQRsi9yXsKIyW8IpITglYKOfQDGP
6X0fU9TJXFVe5Ljy1Mzlduj3L2uyhKxN4cI9cs+y+QHL/Qfq68BcoYXojumfpX33
vUitwCkq82ANIiIKZ4xrnrWmew9U7Lyw65TGGSRJgZdjTtNudqSiMBnG3io+pwjj
CnCAwpGscfca7D3uElHSPDaVkHJjUH6CTGMAt4swaa8ttfckG0L2oDgLJRwpdukO
HDMkqZJKo26Kn4N001EU6b26/gILHG475BetoSsyWROaR/AAa+Fcnn35DI6ql04K
N+hr1DJOB8pr4v7hEe598b36uCXyiIRa+iuYZqvstzSlF/DzaJePh0C6MDRRgAFS
7fGuBzzSFFUadaiMbQYpasWuOFGRwlDihuiO8tETO4trFIY+ZFAUZdftadeD1aeu
JgN2rtJ1wgLOYTiiQxrx5Xc1m0aA0ik+DpUhSS9PCr3ix+hTtxYjiLqpjr6gHqAb
uPuYIq6lNyYxDVMi0wN6RpPeRvuhc2WHByNgrf1sJe+JoK7KhjA8AyVoepVzWBim
KlkRtc64wed0saHiYe57kod6cRQUUrJfK9gsA8B8SMRN6YRtLFNI3dMbRvCQrSS0
IJ2KGPbJNaYyyIuIr3y70clK4kvml6mFqqduEKiqNR7niKS7ib++ejcqrMEamLln
RtIo/56tFUjsOp/FaDttHgpRhG2WQgJIoBbY3ULtB6Ve7puCkLqqJCAbaxwlv+Ej
AXiokq0aq5UuRgQdY/GcOkNeqIo5eHctnLEuKLt+0AB+1O5J+L1a51zuaNYv9Gdq
vCQX6rubfK4g2PTQphP6qes3cuhblsoHtimhbrQETDRW9sQPH2JFBngK1TkAaHl1
ibO9jGDFhh/5DOvsllgUE2UU4LpuTqm74tyuhLrW8ZR1ABOkyhsVjN2RuDOebSz4
YwQ4zQ+zOr9YTb1BwXY5WPAJgiRPbqsZicbEqp1rS03rXs4lzA+ViCHwo094syLp
gnOQz11acLhJvqqmuBbz111xMp5ACrS1o0iqTR7tkvsuUEDnjwREISphIneUWKc3
V9mSjQL+VtQzEvHXZoa71IYwYx2Jr325jQG4atwAwbxe2jUrnRayvZ9rXa9bbyG7
/nqWZ0oHHCd2KM73OqaCysE0kp3y+n8jsDnZKH5pEo9q3zHDp6qs/dzmW2MpZ+gw
q/j9QyKkEWuN0koibJg+uySl8q54dBrzvU6vqm0VstASRoDSYqtRWF+zhXFUbNSM
7AxQZgh6GE/UqvAn1X5K+hNZmSS6NW3xEZh5KvTpB2wz287/mos8eB2am8YwVdQ2
EwlSDhjJRvyrJiKCtY9j0WtPduxrJi4VZy2xzVlXiGU2+gVeUOiEIWgA9jUYOwM9
SJwyV306Jg4+h4f4xWUB2zxRbqEH3F9RTBKZcev3Tz1FkiYldIZltC82J1ecBfhU
02LJHLXlINicOb94+34u8ohWEYPo/EcQgROOJleLyy8aiCmORT70tfoiEtRXsj83
l7W/dK5yTD3Ob3G/VJwwOAiho/bNmRJBps8GuYrSeywesOTLMDnCEDQSuxCaB+UZ
6gB0LB5m8e1j0x+O0wXWk/1PlrfjhDuXURksxirV0CmgrIYha/PIU56sA9cdcWNw
aGmSnDy3lnvL2rX54qYEtqF+T7+hI/KOnrZQhiHuRb+6alSDMqD3UAqeuwpvyvnG
ujw0Amp19X2dx6+LexOkpnPAQPFBpl08toliBOdGh6rALSwjofrh08kUCA2VXIgG
cai+kdADklZcEHMPo5BgmaR8DbE8Lh39mopWnrzbIMV51O0AQzzdvNtMMNcXSi+n
26f0ZPoXBtTFL4eY31e/+6zks5ioil97Jkx+V243RyL7fwM1UYFiJF0nZlLfrkGv
JLh94BiKX5m7lJTEpXdufhaL4gvLN25ZU0TauqBDkUJ58or9xNqGbygXwuo2vBA/
R6rf+DXbofL5guy3VZtutBHyyL9TvwhLontjQIP/y+jMLBpt93IX9Bw/zOYKqLZN
ln7GJFvBwX8UQCnhg6B5fM1igJXg+KwwqhaUXQAXOmU4mk7TFZqRgZUCGcSEsgKI
OPCRvcMkcXk6viOwMwk4OP+kPWNqWf2xbPSCADZnVq4qlanQ5Y9j6MbQQFsjYCBs
XtUqJzD6ZYAgA9maOvYRa0acETR2cRKW7rbkjqW+7KNNMgBdGOHkyRA/vlRsxIF/
T9aEb1XXikjkNnqRFtSeEgJ3fTOTaE+24q9fMa9Ud6pnGkmGfR2bJSQx0hrUGB1o
QI4dhPb+MOUZ3XG3sWbG4/254iv7P7yFcwm5J3Z5v+LtqWrinGmMo1KvsHgrZ+XJ
T2Zr64+1w4sY+yQASlRp1/MvWzQSNe0zJGJdS5Poi4kSIUwMC6NExOnSFecrgXOG
sqqfPgygglsPhqHsrkFJYj5LS8tdHhi+TBK1bKRRM0FpHVKSwOz1j+L7uecqK/CB
uhtjRg3/WjZNsA+tmUcpf8p8/ZF5wy9YTWMf6upUZFkHiOkaB0ukVKZeQc9WKfag
VXlBpMNKSiRi/biX+2KC3CayZQwh6pEQr4eWHmGvT8b53lFRQI30YU9VaNpTbOxA
x8DQObYD6+zsq/F+pC3q0usESSaFuQGL8hlB0tKy5xdTn50+BIQeh279LnDl6DCM
+TuveiSP+f0Kuem5BtpOJMJZ9NGvUa/zzKM4f10KbePWv5VTiAUOrngiGUbHLIuA
zlJ14N7SAJK7woNH2u4lcvAndj82RSYxQU4RG6OoMM5S4dk4hhgTZsbeTtChSxxe
mWJlcUgD0jSPlk3/ZgtOxTGbUzocSr8ljwOr4wFr1Dgmp22/8mAmev5csK2kcjaW
rZmgzmQSXi0fAm0rSfWzxBs0bCJHLc08BhRa9CLFE0zSByytOIsJGf+ekZutU7u9
gHdRFciYHT2lr/rwXXuG8bPzyzj/zpIzeWEv602I6wsds3C2vDZVXk7t3NRU3VhO
Dj/WkUojFs3byLRsG+OeeswwILGEGmcmwy1Sy4Aj9fW8VMZgWC4sLWKX/ie/vqvg
3vUwkOQQBc3kLa7UZ4mWyQxmBqHiIt1eePxNbC20w/EqTQsH836VNPNTJoPMh7lK
4tzbAmlU7sHyT9lDMROfrv0JBLCym2vWLfvDz34yO9COu0l3Vp80yCgwqTjqQi3v
lO83sLjEevWZ197NoIXNS97ePP8K+3Q05ocZGd12So6U5LAIpU0HD8kgeZwCz1Sh
x9xzuuA5hL+Ya7OLRXUqU5ZGeS4eC3KbqNGfIVIfXkeeqJYSs31/eghPZIaQIEF/
qOzQCHyE0m/5r/oe6CYmo8/pdUP+QoEaV1/zsz4JUfrZ6OU6K9RUx1BpNjeYKZqR
B/Rc7Me3zP6xxvtU9Eby1p/cGEU1t7mmGS3qDKgxa5xTNrY3B1v6/7qKxPLuczfK
Ys08BrK3vf+6uYyfiAh9sKMmPANPPpGa1XnVpvnxIfYqav842zmWH29jSUn55Ilg
mqLTa+QtHBdQ0x36jtaLBj3cAiVDeElGipr862KiQjKYlBMDoZtBxQfkzTl4CjdW
exENTFXq18laA3uu2Sfu9NRPNDBUdHebtaE48bzaP+wP5xMHQp1Fn1T56Vfrdkh2
E5DgP2M121BB377iJzGknl2Hr16azxwwGfSKmKABa1cnSvchEwv7Ee7FACRih55r
g3KwLLHd5Q1c7Ivn6s5A9NeA7hYd4FmQG1R7h6kcczId4UUwgzP/F1hOzGLvt+u8
WWCSxrV0TvNGtKqMDo9iK1G5S0UEKn0UmKEL892+/Y8nAk9x6fAUmjxWkpPAE6YF
i/Ebc5xbk7SLR7ad7BI2PRjENK+xvOIM/AT92pkNWH5SRFml/Ood3X5hsb1uIRcj
L7Uthd2yGVxkkJmBasc3THRmBWa0xh6q5Tii9K3jt+s5H00qMFCOpFZdcxc34bdo
26deUZdds3drkAL20HMKR2VG7V2quSLqn2AggaGkraZ20OJEXPQHBXXiENX32f/D
ckkstRhdYMfCdt0Rf0P2wiE8ANUsqxmCEln1NC7wyq2DjHW1iBSEKkkEttY87uRN
JxaqAED/6exVbFyGt0si6jnhDrc1CsFOwGj2dXgY4RfZvJCntzKEFfUo1Kx/9bHE
P3QPsQFJdFGUhwH3a5FA6Xp+OzkEydya2lWW/0gpE9nYank+S9SV1tqSs60BeGTJ
zxX/B6YZv0/a4PeU0tRoA9O+FZM9jgy7U7EK+N/uVDmxKa+tESppWgDcnRn1OpST
RTcK8S2JQa0QlD/HxYRt44pVmpT4cEVyiu22KcusevxTWcERJKKXtvFPg1wqvRVH
8eiXvasefOyCjtEDM908g+mMT5TYHrFJTxLI5TOwnE1XvfX+qBoOPZNaPXZl44va
qcWgP39rNubEaUFayAKET8Acbh/FwanyHJWYR5a3Tk+5mLiDriI36b7bozBUX2jI
hkrSBm3cX68b4sS64IV22y5PfPT56QJWSjD91mk7gV2SQnh+5c9RkrFocWllZCI5
dR7RUYOYkKaSufVrAeXd2wK+Qb2B7H3Txy63bRCxlE/jaRSWiOD0VkspdGBkwvNT
bPdcVWQ88Q7ja9LIDqu7LpVo3W99gITzUtE9ken0ed5h/h45ezwcZiOr4D3+8PNY
BpnCEkWj7F2nuFQXZ+rWiA2IAaaC17cLjEdsfwyvqzhn+gsBluvk7Ftq/2zFMMJz
DYOEcEuPHq50RSuSIJLYwluzEhzJZrs8Yl9uGLMiHq49Uh/3tDVPqODnwzrvSAt+
WCuasxgXHjs/jRawEr7GIdSOIWQaz0IGX2jTZEXnqM5nXCqUngYCPQu9/2rz7+E+
M9SbYA6VdbtFpqrUaMWJtPaubAZB/LNFkwaQZzFA0O8ypBCjew4qCfqQO3HWIcjQ
rMg/vk4iXxAg8XRInxCtUO4E+BzspigDFfNKbsvWxF013eKBZN6UA6HaBIMwH1rs
LNiHjIxShaYBT3Eahmylb/uAvauSHrmL+c5S/ZYnncAiqkb5ElFZg7OLB5Vrwuis
ZVuxO4Rodwr4Ba//ZprCJSYmidvIo27Wcn1c7A3no+dinA27I8GOr0rAvuikbcZh
JaujL77kLzpPuIPe+Eo5eqCGUXgG2gYyvv7lLh6et+xYDpmEFOss0pAfu4/YOx+W
k0a7jkgfqALelHlEiLNu0owVJHKRB1LZ8Of7RfHhcrJQSN6e6yZJZOjRPxuKKreu
lOdqmCozLRbISbecs4JjQV+bFdH5qCYWOHAACVCkyZlXkR4oMofLwcZqUCAE175b
OaE9viGv8rM6h/wRd5vB77bql24gr9gU27x9QVBehd2xL5tsi3g84PGtq+s6jzy2
+JIHCDEEX0TPzv7MSD+zEdfF8dUUtX4LUeBOMGUvh4XKT+WsnDBe/YZNZiOsdjd2
lpFMfHHkS/FNqw7dAWFod5mfzm+Uv7k4yCJqdPeQSa7wlyOM2otRYqvMrFj8UJDe
crxgvOYOXOw0LAtagwviQp5OdcodfS5EW9JgH75ka7Fa3Ca7LlJxeTtIGfyb80No
/dXtfMLYottwMxXk7iKVKrisu+FIN6FS+MA7L9P0/NYn4sJoDMeabWRWrLCACm19
YLrccT9prq2LKxyBpWUmZsAGaPwtlQTIFHTroqkZpPWcYMSmpSDT6miavYydMzOJ
PYkhW4ZzR0fTm3llauD7Hdxif40VAC7CqchlG6eEJK/YMT0mmuhgp5yDsIze6x/G
/PfyGOZ1Arlx9uxOAJgih5HKaGJQbJ/R1QrI4URyxijVIGuJ3zujotGPQgjG28Vk
gL7kUbl7mPW5gc8Xqj8Zciux909Io4+PU1baDVgTjLYtbEb03PiVHmloDmxcXUf5
rnlGxvnD8FNQzgToiNFw/QERN1JDBixc9LBrqim1ChLtIzL30osLaQ4Op96jcHt3
3oUQlXV+zufc5oPd/NyQ4ksnpmhCRaarnT7HilWrfmbWPM/sIKWbJSe6A9EkE3kO
GdaeZeYo+MNvuRb5+WBfAoKUvO94iudJhhmD7gUSmvcPIYqhLmnbXlzCp4trGIKj
6r+cr15kXUe5PP+vw8eWrL9HWs1QU91GvMEmhjG/sZafqTvg6v+gI3Dvr40D583r
BZMgsDNs5lEirowH0T64IfdYAUlvhE/TgyGAPhXWdrcp7WVtxfX+z8NmaiEKS94M
VzB+ZB3nC5Xhm5qD5WMC+fps79tdl8Vwnn5vVFbVwTJsTJfK6Sskkw1uBRLeUPUX
TsAnIGgSse/VleU6PXfykig6rE9sFSa+/BYwRzhTqMTu1bVD2EgraFVdT5JnhfXX
CfeMYgsmchMuw7s8N3yZqGZ1hyP9py/R1o4jzmT8sjCDrZ7INGIILIB/Dkcd/56f
m0nBcujCZaRn56IzDmeMdyKXGasRyFtjYXuPnPf1odwYX7U8TbRsBrVuBQEFKSwh
6JTzy4foG1WRkDkWd23hssJWybLttwN6lWg4wmYWhl6S7F4GLvtnAz5KFk5RmFal
qHId4A86K2feobe3BrCyML/IcaCWgyb3SSJtL1LRsATQQP+bqfl3dQXa+gVKqRWb
eFrRlVdMcDXTolPNWHYlHbsJrWEqonYbRZ2Xzyc8kRp7MqMZY4jdj92uFC5kfqDv
9yMsJgJHeE7+BP/kJ5CgI4PqSHowjj9UrsCaWjVXbolGuwMx8hxFCExfS2q0/DMK
J+P6H2vWP4P3KlpiKf1FraqeNBvXz3LuYqKBpQqI2q4yjLD53ch7LBup0LphjONl
6Eu80nz/X3/Mn/bcL41R9FBhMVwNv6aj2M1th5aaZTev/nrZX4EJCO8lPGY6nV03
/Q0kpeFfpAQSCLBPcDi7sPMB7j2Tqad5hHMIRREzUisQs2fJiiY6uJ8h/PLSDf1a
JcqBLuR+MFQo2uYDZm9ksAmsXzs0Mb8bPAgkSjpJ588D4o8lDFew6unUDsXXsJku
7NKnglWBk2W0q7ypDlTUt7XTAkdpvIYsUBMooipC/LSwR/UkZoFYGiRLvjTRA85j
3/56D+Ykvk2neI024UeM6/Mr/Ck/QR5xHG3i8spIZvoFYnATix23vKc6Ksdi5WCM
OfJ8nmcRL35vaBfj8Qg+LSd5rFiF20aMRvsBes6TZK+dTwC2mDn3IYxxPkpXL3so
Ny2EWOtMoOQ6qeKI5z823zNQenzEHXK4TQOsNrcj3HeknncBBYHFO8gsP0SmTSEV
hSGUFmHb/snhN4vJeHOhtSDH/qpNXGe0DNDgfAFKNusjgrRkQqMkf9zRaZZrav20
rkTMC4Jrll/cbzrvgDw1oLvneG1TEl3oER6qv9+jd+8M01KX1N8JOoqoMC0vdHkV
bCDRt+5mJ8S4iIJAEBXjGN+Btels08GCZ9mNrrqEShY2C2Xt+T7jnRMtUiAl1Ghp
SlIncg8EjkvnFedaKrAGK6MyN2G76l/4YvikRTTmH07zzkrOt35l6La7OD5pGGiC
XT4xSjgykRnr9cJy/L1k42qh3OBw5f0bZocoTwOP2lc2B0ANloztTIZB2AV6VpbI
thJDQHxKx4IZNQzq2flvHtjzW02i5BM4woUrcNk8KmY3pyJSEl0aU35DzquywKA4
CWPp/iXAC4bO1cPKUaYmcOak6czi+zezVBHg0XyywAUYiC6PXyO55uouNrRE3NB1
axgrsQexDhfQpzhi4ykEy6xUXMNlP3vmI4RiHBEYaFP8FKwl1zqCME/gs82wwZ/g
C/5VvktVPWUSxZp/w6q7jSWArgqZmhrd2sKEY5Yh6GHCz5R1SwAnxclnlpikEnw2
LC2+m1tIVeL6hCbgRcTCKk1qwT5F48PuHraQhBUyCEywx+LjPBDtB2/boWxnhi7Q
Sw+TcshzBxrwpyrdWQzUSBxUun5Rpc0VKFng+BQu5rVIEw8ibscR6ihpEHFAowF6
0i9LMHEw/LUqfT10r2r2i4HBfBGuP7BYaRknS9KaLPRhlZ6xH918b4XqDMC+mIRh
qv/56E9m19Fd91j6EEAusflueoPO4IT1vYTBO99csofMrbAIKqE2TOFIvcPGu5eu
/WmwiUyk+pc9VESS0QqbTbPNqWgO5LwVJU2LZrH9niws/vHgJQKh4YKpT59DIvv3
ON8PD3pHkcXZtu0yDY2XHnlYWjSGcQSTCD230luJfUl+unIwE8BOmYRgpfUPPC+A
yPEV7KW4kDpi4X8nnKKR30Zn8q75mejPXYalt8EgRPhuEmDLiysuNKF6p539/251
/pNam3ImicZbTxK3JClJ+yWXI6bugmuK7YMWEhb64HNee5gTWji/lInkN0AhwJkW
BtfrDFbYfXdONiVJRZ0Q8zlP2Q61nkEq9/qhKy84E24EX3sGyE/F7ZzuqXECEydi
7zncI6iB/J3B8lcyg3T+zFO//XulBUx+kfjd7DpVuqQKu2FtwqWRbOqp/KEXo0Mx
nIypcriFzQCY8jYbPc9XMGYHqktXkGv3dlhI8CHTG1oig0zEpcCKe3lkaYXuvANE
xfIEuoj21dZVYQDZau9zJtjjufb9SYWxM5lLSYAU0cvLUR74MJbqyeYLJQjWAxwJ
3EsdXy2zlUvFzCfGV5wKZ4y0EXoORGlw1SgGM0A+rBKyAPg8h6AU+oU375ZfoHCq
9GI4zz2ZqedVcgDBTkM9N7CL2AzIR6uW+8o8vEk7M1XvJocs6PdzSifyQlEOKD6a
2yAcgaatgB9BLiEWB6M3rg8QE2QJFtCoRfv6XfDopyKx8oC3P+CrXFoO88cMYeCJ
7fPYc1VRqnQw1Qj997c+2u9EfkZhLsUxSQ5Q0li8otbdNNQasUE3JHAOZ3JMY73a
MVrlzyYkZnXIv43zjTotQWPLMYLdlKrKFJG0Kf/OguL/eaSSl+Yx/50REKi473sK
CYwKNCZ90mssH+DxITqqji8ISBCratCLqe47BPK4/kAsE+YzSHejfeF4ZjMAWtd/
svhB9sOJw07bs2R/iKLUTWEcZKqjgaLdr2jHcKhyrUCZGaJ9FV87I0OIvHhQ183i
0fS8mYHsHA71QBYSdN0s/iayyrGUYpO+C5w4akEJtiBZBom5kTC8gPc1Apq/cgtg
aOnb8QyqNxe5iSerFVSZlfNKkN2naxzvt24m8ZGIwCnQ0E/T7U0CpJrLIarZ9Se9
2qTnenw/mA4gUOQIgbW/koknU6tyo46hzKH0pB69Bqfqw0C8LW3jUif8TeGTYzlc
euZjsArEwKpFxBV+/Ka3rdYGtiPpYWONNsKk91Ybh84CM0xyqCd6I1tQfL5N/7Ez
hxnwWaP+q9uP91e/K9ld6rjM17FJTLX7513C0QqZz/OE3CwtT+igNrqh1yEwbOVG
BtrKDkbJgaoJskvmjTjYl/kGak5RWgvc5EBpbsNDKYTq1gVMxg48Oq8wYr0WmWQq
Byg98H5y6nc9odWTToVE9dq3o+q19/tUwaxyYjQp/xFte8cQ7x6neaSQu9qa2ly8
N8GG3ln6DAVPRJz/0nWhWt1SGOuwASyJxeozsGJw9mHpsG1VSFLNRVrKsuCzT22w
+m3NaCvwH3rDI/0ZjWXBffvyG5IgLOiUxWrzG6CKMb+wq6A2KWbGjmHDO+3FjyAs
M2Jhn9UYRvB+N54CfzT+ySl1jONziVoTlXxfptlO0eUlDpW/vuhuY+AKhNutVpHF
8+NKgZ+/fEdYpUz8vvsRMu6SPm8GT67o6FQ+WZJcVZfoxQCY8sivIzTtsLHcoFEG
xVQuINt9dU3D4dj7pRdAzgHNuOFOsRKp3B4OI7WMwiK7WatJWfLoAi5q3E1FrJCK
d+u8zyO948kSYDRQ8VOfTZsjlBkaeg2OyzV8J/jYw1Q2ftQAnwnDRxScJq/8ws31
/GwtqwpP+/AFzV8KGistcAxdNuFve84if8aNDETSqvKy5MYDyITWWIVedzE05UsF
hu9Ya3M59jsq5bGOJB+SOS3fFMoKzfLeROaPj/9rVO2LvO4ZBtTJvuThf4YZs7bT
tTYwxDxHjMIjzRNMyP2QxWccr+kvzPJ6mn2OBxA4V10kT9vxQJ2q/yo+Th/VUxO1
qTdAZur4kRin1Dfah7C+7ZIHN8ZGV6quDZcGbIjHDGctUh9vedZl5z7j6XOl/BL4
oRHiKNTyG9PrzcgELnbW8vxTGjc6YCWflw0HSLCX4/1mvTsyChxcdoj4cQ1i6FdV
k4e+hDFRxCjt4UwOsXJCDC1zKadL9oG3oXudv1nI9hbaXHGm1hYuSQaxOIrv/n75
RFIz90v9uVGIrR3lF34ZqHG6tFMaPsQO7WuprYV7EYqSj0wn3Kx63RIFcjWB7/nW
T9k5NHHRDhqVvKWfq/0xeXBUOOls1w99kMUGTN6EiHvm934EQTzmR21V4OToNa/y
w764WnaKvBnanRSDMRG6fK6fmQUhte6dO+sVGkmKcvk0Oy7VxztEWNahVCQ8jPxC
G7vFXPa0eN3SIxRmzjrgX14Efmh71XQMsqHPwyD9zxLL6jpLwYR5PZAeZ06HgtWK
LJx6fGnRfA12Zu0XIsTnpcjPT0TFIG7OInagUt90YyYFmg12xmejdfjs8j9pftTd
pMeNwH8HRZ1IlsANkrjwiTqBbNAb5aE7AU1yWWpJcyU3girvSaRgRsv5gKlrvPB2
S5RRiGeD96tRY16HWvvGM6R+RqErOvLE0m97XFBv43At07JUrsNqSPXSLo9Anb3h
EtBLCbe57174ERjKjkPsHkxYhmBKlCIZPIM79nwGgBezdkZCo0mp2wfETigSNI/C
O/Tv0+7T1IEB3T808U2Nk6087PGK/SHoDCBYxPx05ODpFDckN6gGye3792VWtX6c
j8MAxjz0CKOLsosVFe/+ae+3gq79GrEka23bo0dqmbHPXx7d8/6H5SN2HeOswhaH
89x+aphv284YEb8uljoBzAgK/rv6Buu+8cwdFwmIphMsOr6VS70uj+s3aCNThfSY
DSwvKm2P+fwEgWOHTWA5CarG+fL28HkflmoLFpzIrmFc+hARm+vKXhSysi3wt+BT
QylW2Bo4jr1KaGgsxSytDeCyqK1xwrUiHTlVECi+FnxpCocHnW5XCgHd3Mg+RmQX
2Zs67mD+/qGLyN4LFvVznuposajbjB75CC4Jat8KCoCRMsugQUxWZy4yzhaZG6X9
FinILoc7zahq+/fYxKlyws9WNqX+r29PubpkWqh5R1Fp9+2KISy8DOTybX7BcAq8
kOmLkBKU72esPpAU8CLmY8ho12xSiz0fd8v8oYG7HNgtCKcT0mkxAnTPWv/mxuF1
lyoVgwHl2SkxssYV0mK7mcee40aXKn4mjNOMSUCMxHZwSExTIxWe+BONQlCTdt85
wECr2yJDjdpSGwcIUmI0iZZxWFgPJZXtWbuyWu3JfMjdIuvHhvKZrinQZ4atlvuk
hd8/2hy4BIJhMTQfFTDp8bYeBlX7+5b9T+3WnJ0Zy7uFxbOmoub3E7oSi4XbrTjP
299Ag8N4WT4JvB+tjfobkn9cMFrEqQlp0usmn0VjZJRQE73Bw5pMXjKoY8HqF524
Ck/uXI0U8owR1WTWnEaE3ZB3nmDJbeFirZznjbHODT2GZWHLlbflPpygtYw4NGos
xYNOGT2Wq3lSQiEEREFE/L3z7VrCpXLS6pU46XRjXjgL54uoYm8RcmziP1lDFVfH
9E2KG/dcdeZD7VTQD8jmbS7+de8LiSIYIdckuQVvPDBxFMwgUZJMMj/Y7icUxcUB
Q0tJKHHB+W3jk5iq3D1IGZXDPSoy8v28xyW9JdUNcsvzqGlLR9epqfkAjndSkz0C
yO0DRYAy/WOyY82elEwBvU8wu8/d85H0Ede1jVOD0ZgVAi91AzpGMFJsyoZWrbCW
y8a0Wcllq8XejuumKvFKK7uPadesL1+ZnJHGhRfK9I4wOW8qDYQPThETsc7AFOsL
VFODJ//PmGLAU2u2ofndppPxPmch/XEup+yuwqATs9s6qJj/T9zjlSL9G23oY+o3
L2k5JHGYgi0PSbNwJBL9391h8J0ylc/GSd5IGdIjHyHlQ1U9JM7sOKxvoiX4/u3P
7wcYsvNEWakh+4LTU8xO37RKW5ysqFSESJgPHG6NvuF4/L2uGnru0wT8mBal5Lkl
IQAr9rzi3ux5SP1QK/tmogQ1TaZn9reUV+xHndNLqH371wWt9TV62N8p9jjriBeH
SceFpmWvcI6BqeFI4eZ2T9MZMjD9LRvFiVkpXPNTIi0wt6nXyEnAoCRNVoDxFiAP
A64yh4LvbFzz/bc4IqhvYJSNF5ZPmFVszSWKD4WtU2J+2Msso3kUuHDchdfF6/RL
NZNoJNQcQSKZCk7oH2rdrRPL2rsotnTKBwsX2xmpPs9J+kkmaDXywCCxf6h+wErA
WOEyUjO6IR4prJwD6NxPMjd3xA2n6eAcovoVIWTbZJeCJSk2wu+pHDR4cL/gXNI9
JJ+kENy1VzE5M+/7EqPoeDIdfDV1w6LlV/9hk+6CC0fA9PsUKnvIVdnmYaV7jZdN
ZA5jeLbDW2Xo6aGS+IplpDYP35Zo4s5N2O5dNRG0FGSwPoh4K5U9Mve8KbjjCkUK
wSlxb75uX5qq5sWZ7gXRMT90QIaP6BNCrZUkOdGGqQN5DtR9UEXOZ0RYFSLzNzy0
g4QeVdAsMrTnQ1I4jWkDUB3qlwP9sIiwn0XsKVXlziWp8oTW6maYUo4lne4UOVmf
hMTyWquO5/4kzGZaNrCxduJNzDsmqb9/gSL5GRIQZthTwFhiDM34X1vGt5M39nom
XvaI4O4j3LF1r0gVTugDKxCbQ+A/WsPfBYV21x5F4otbZcnyQq8hFoonilwxiw8g
MZAaK3YrRXjuCn3azxH16sHqyXDbi0AlESZeX3FL7DhyuKqYo4mspfoHlVIQUFGS
hCCFyTx2x7HRZaDW09vNAVdI+PkfROX8BWfaH4gxWVfSaQ2mOwMASmvTJn/1S74a
Q+R6v5mYugiUv7MitjXaqaH0cvy84+31g/AW6Nqq4S4lh/xOAGgn5d166arEj1ey
ANJPOvNd7N2Pha3/P7qebV9Ps506xxwgh1qoCB/QyAf/Fla0/cUggOJHSsV8V/bA
VoeA5WMGxm1ztx+IxXhjTFS+nSRB2s+7eylhD63oysni9YwfCh5iaPtEQJLFgUz8
6UPmvSbSB0O2vpcY5Gj5hx6cImTw87u4ifeWSAimF5FiS36TnJRLuv0zAtc78nGq
NYXBwKPFNGPhInMES6FVY4NqM8+8RWsgFI9GOSaqTgetpx60DOA0MWWITKbfV+ir
CxVoIIlf8SY9P1xRyudGbmqml4s9zYxqVnJmudyC5ZrZdCwVbIiHCjeK3TdaqdeJ
n7wY96M1AYsofz2z9SUvlNhprVsuHLHHWLrTWlmwBAwWey69TyS2OYV0m0533xQW
/6A061mCW2DYXhEt7Rrhyz3ke0/J/xHfm/dWGD4etbmw7j50ThsgxF++IuEhOTOT
Bfl8YWsAVhEz0ePP5ykxTLBCkS+5Rb+5+VuWVjpaSCB3vTF1QIGxGGLD4YXH4gl/
fYu0QOZ0rgik98PTFjeHq6zx4WeJjfMgx77kJvvIC/HYFOl2zi5F0gpwY6d+jPrm
9zl4wN3QiHb9iB9kItGgniIr/ntmMl/wkyMjheXJPKs4UXsdt4fix9c/0MteZxrT
In0STe5whHthKJiM+VsVTFvNJOuJMhUme373ztZuoD8AqvpT2R4bdO8D9nWBmJ04
3AfGF//EM82Vx9z50yeRgDqrv523nyRLO/0k6og732lIpP0A8jkPKxSHFQSKrSV2
8YLfgSCpLn3UqCOK/2aGbd0x/V2DgR/+K3/l4OHYSRL1QDpqVoB7cQ/51imSMqyq
6mHc6L59hUVvJgORF7ybdWkaKJXgPbLY2g9d+vm33aOOb18Kv0YdXB/ZMDCmYvqP
zP8PMz4GMHuSloajdgUmiJ5NEt5TfXEQTFP3fj5Sh9x7PAyz/P+XPk2se0QAlru0
zxPTMoWHX66Uf5COP5r+OPHM+xC3+U0z+gZ7301BvKH+oHeAW4o64IbH855xTmwX
0n+w+3htqJAocsXb+n6acrv27VdkSfEoQxlVOzT6DvAxwJl73uNblf52V6noqSsw
+E7BSJrVAy3bXVwUt7IZkVJx/UD7T831Figtl35XUWMOIasVD+VRmujdlJsHNqAF
J18chhLDOA+X0uN+239AbGJqqAj2TaTXK4+FRR3Uus6ppR3rxxU6FfLJimLczPFT
R3CApqWh+/oJ47lbRVytkEId0cPn/XNLP800GwJRZyTKqv5X9AQQlT2JdLuOPZtl
IgOE+1am4WFvASg+OhHF1x84hna0xVo/v0u51Crno8d4s7Q39MK7AGcK7rJw8NSc
On7VnnJ8WpFQiH/RdT6WCknZ1yGWdgng9hXU7KsrFDpAG7MvASLf6H/OEegPOKnm
eH8SA3zhwYNQe/nUGd8tjhC/gkGsWIk5dboGDqe+C3ptbMm7Z70AXGCbJoiHC8YZ
Ubi+2QEQ5lZT8hOo04hCQR0MbEQHAYkN4pI//q2lqWq423GPhrK70GWOcW8pfMc3
C9OptuWv1dOQPYKHkMPr7WLsU/nyGQ8/f0uFsGFM1Xh8lBAdKuPbOIanbuC8228p
FvhZC/+Gb5B//8bZDhafriwa180kxgMNA40nJH7NuARNJgjLzJEpr0TVTml0hGxt
XxF+8MdtRert+AK1u+P7VIfWYELFhNvn1LSiOvRUfhcb598rL2Ch/c7oPTMVi67N
SM8y4dUK0MsZbyqhgPmvRksqpi8LfMnnnWjz1lSACarzZNrHaQjU1RJdN2HfmF8j
4EGTWnhe6mvJmfhI85DBQnfjFeKelzuX8STmInPKeW3P3zwlBvF34SheEc/aveW9
h5P+r23Xa47Ycxvq1uM5RWnuGtDomgNJjxgOLIisyG8aC1+cToWmStrN0jxLu2kx
2G5Ojj/v8j42JxAbXZ704OvVXSeBYYWt190mqxuSJhXpIUB/uoi/Ne3MwV63yR85
JFk4JZaK0XziP3jVrNE1gbL2/J5H9iT0a5NLCbMBBQB8INgnpKwXBk5p4BLCe7en
QWQseBwXB5eM0pYMdax50FKtCKxmor9agnIN4DTVA5pEfwZXNDMI4f4w3+751iXT
rslK7xmXt75V2jughGYkvDo8ogwfzEZiYrKnMtE1RekWdi27+t5Xud65R9FnT02A
JP+JH7Py1gwzIp2Mx9ahPaikwJWAMqe9kO6shzHT44i9D6AIcBEXD/5ec0p7kGV5
17TCfTA8K9Zk6T6wxVHt35j3in8WUatPx1kzo+4bc3t3mxpllsikPBkF7YzyxJ8J
2ppsn1ZPoUxsQXV9DKycRsE2HuM/fEkKz25yildYEyo+UgSui5LnFzxxgn04yhJX
i0pv735bNEa1Jtc7raka16YwhpvKX3i2jjA1blHtRR55217FHSqj/DAqVC1zvZvW
Dmtn+TpgH+MQGv03lA6GdtueF/aQoQUZdLv17rYj4Xh/BYEfBZn3Wf4fy4aM4Ggr
qSeM7iAkXwqBowzKFCwlbv/xb1UHTqVRZHu4MurdER7TyhKJ+bC4rLze8sHk/woQ
4bYbmcDLsiJDz3kf6ArGWYqDYeN+Y5PgiSDkvdYXVSaJT1nZFJ5whYvQxjuqi8qO
rlpG3YaPZ5RRh5kQxMd/r1FFlR22g26iSroZGU40lyzrxLI3jZL9r6/AGraPf9LJ
TEPBnx1r/YOh0crv7KbC+VQLZuhz1t2/ixM7uJljo+Fngq17XVgxtnEHDFUtmKb/
zsZiSO4BeEA+xrV7PP9sgtVUWY1e5w+sCUauXi2RaIIlQC116gXt1q9TYMHp9VBb
0LmoVYfbph2EPoXZOsWsE44MrSWHUnYYWrPwVsIt8OUGZNrlyJmIjX72HEEcfbgV
P7KPsW7DZUW0Wh1qBoUUsJfi6NujTbBDcWJbNKwp7dFebCR9v5uJs3HsysGtM2Hp
cr6d1bdpZQnW8pPZCrSujSXm78IbLRCUMsC4qNoUUXqsVxgKnOcclHP8ek6EgbV+
TACJSA3CJX4eGASD1TPzGLEo04YY+RhY3cE80PRb/ARw0ypm+kSc78O8hDl5PFyA
xeSqKORvFejml13U2VPKpJbHtGwDSHgwSdlQRL1VcZKxnl+IBy0jhlNxz6ZTOlTI
SDFd0YtDJuvIgIbvKLlt9vo+IGNoCdf8fGDbW1RoDPgMHpGh4l8nIEN1mgNb9wi8
8+OBb1gPkYNjOEg5sc+CPGZMR4+1gJM9C8t1YLDAJFW6qeCEMJeJ1d2DicTb9sUo
vPLbPd1ts/c8v5qU+tOXEBUL9LiWW4NrtZy6zTYocMgp5EU6exjl0PE0Z0yuiMxc
YF+T84EWQodCBFgKJM80/eW2fmyQOYYShhUDv5LqoF6Zkufmz5NJvHFKP9qaoNvW
vnNh+myAicFIFKsJtsiWNAbDUt8OTMJR+d1PXKygRacXANz2KV1+wOqGvRJyizEy
PNty0DkG5ziyFMP7sMR4SOBoPu+DSB6iWHkjLdrvb3wh5wCMMMfIoABlcavgZgS4
yzBY1GJ5R1SISGLUsAh3DSTeI9VY84qit7/k7REKILaRYkv9lyLFljhycXr+YupA
nPGhCQC1nc9fyzHT7JhFQ8SCeSNE45lMHNtAPtJxOMvNX9ag+0Dulx27cRa40Q62
+Jwrht79VBShXt7o6jfL5WOJDJbFO7lnmjw7I0fVkxEH4EC3neHXGmYHJLToqEy2
h95y+kFSVB5bNp3zW1/78vCU3raJ46i53APCa6yZZjAlavVcTSp59K3OVJmHSYHi
cdBl0RewyrrY13DcuMtk6bDpfaJgwzd5114BI1Q1xfo1efEsQ94QuGwu2XdZB3lA
BtmguLS/AH9yhCJLTsqhr127zeaceTpXggMVeuRolbP/F1+Ben88e5k9Ihq6dHKY
s1A51oV5H/8Rrqj/9CCoyK0Is2ZnTUW8LcNatz+l/asaCy1RrfIZ/5/FaFj48Or4
TWguv8kytXyLXKgtsM3N5HL5y6uePkUgRKOmO44VNINlmAnNGwcNqGzclb6bCwIA
DCwB38RhDuSvtfA6GdSlvHPdu+7XadyxQZtNEfUlZXvf+idM6yIfCLSjeAE4iFeb
ajGosc4qqYaF52ARrATctqhgef+sj5tl87B+CEwFotwSPcsyf32Bp1WdjQE5iyPy
+kcbuiNuqnZtIf049xl0knjYkrvz2Q2eW6ttcp/wVN0v0QJOwQdr/3t5xCbAj9CX
2p50xU0DxhNLaSTszq7NmM64aHpJh2anNC724K/QfrXzfLIHsONWpPrqpcPeNl02
R4pJYsMU0S4w43lRjyY7RSCO5jC8AklcGiHHeds8OgNVKGPH82yFcR3sicwuNQzH
lcMpgt/xHhuQKC1Y+iHGcE03zXuDgVxt5R8xRsxD5cZmRmmVrjuZz4b2R9d50x7+
Zud2W21dAz2OC7c5ejeUj2i/KAzKHldamalEK8onz2LLUZnqOA9Ajq5Iewyo+RqW
jENULAYCNMTIp7sq8epDfg1tVlaSwdPmLfaEIQ4Wcf5BihAHniBO0IsoMgq5GgXW
cEIqn3qn5g8r1wOSg34u0gl34v9QZJnD9RXXA65ijNF2VuRphOq8P8mVTmrgW7jX
mCK7xnDqEextUdDcHIi1lyQ3Z7FXONlKSyVN+ykRXMQ+XkTn56igJkwF32PNKIAh
uxIESJ+ijclcCUnSiwBDmXz+w9UzJy4VZjJrBOIFnh3B3gu1jm99yhXNnu49812i
+3yjjMQ7svdNXtBvQ4uWUNfsjnWTe/oj8kRgJhj3PE3HZLXh+3yVyTn1plnW3R5U
e8hCKagPCEoBlRnnmrkOJHjZlzcAtmLC2QV96kBVZukTWtolYLLK1604KTfGGSkq
1ZiXEqSOCgi2Z4euyKMYF2WMf0vhziJBrSD2DdWI7UAF1yFYJjM+7YAjAftyTJRQ
Me20ZEcVZ13viHbmKsk+SUr4NVuD8W9Riw7UNDpgMPTPFP30amEFPmUvFtKZDbP5
Gl0Ldj6DnPi/KpyzavtDcU/s9EfaKPjgfmJDcKU0l60lIFiv558DJk77r1xEHY4Y
Ai8FWyWXE+4k8TiW4K2qL+y6wwrazGTq5idKZTpFughN4iUOZ98PmfFUs0cCk7uO
l5NujUlJ1Fd+KJykxNrybNHkIey7bwv7Fqs/NsTA8lqj/SEBzYvDHYO+UE+TQBtG
QhDuoaftpzDLQwiytAiqymvvHcTWwD+qfJh1rLuwCpWnoleiDxvGBs9MtzwMiz+X
6k6t5ykMDmTFc/Zzc6kg4Rb7G/aa9jvj2xfYxElH7OtDOTkGDc4jZmBocRzZtI8/
hSav6btvzv0VVhB9yColOv/C1BLlc7waAbhaq5FlV5MYHrFULGw1Rx3YF1coTaN5
0uec9Pv8NBgcDzjXNyRDEfHU5mpZ919wEjgv4ACQrAHW2nucKU3ywNNm8JOjwaqf
gGCu75frf8ZPH3UfNkrSmGg0YbPYpFEpvwzCiElpSLBmt+k8bdBQXd0AC2qA9+9M
O6YYRx5RCAcwoYVxkTnhLTmZ40GbqtmA55WWK2O4is2n60Kjg1PGWzAFTgqCcN1B
snADR+6BDlgaHHkUI0XWqA8UuE6w7EwgxwY8dvd1xCsNVRprUjH7MxWcgr3S4BLv
+alBLeMTItUdqxR4CmFLwtCSI4BFud9GITEDMIH2kv93I96BRSN+pOA07f1W8VxW
/vsDN2moNU/hsqVE6+laHEU/6wR4qpd5KiKTqhxdCu2BPBzCSTdB0YTfr3/zjUue
P46+aPwh9wBR2UrJehgLlOkresOJpfaMoMU4p5sgguYjOMaSNzsdpBPoVxJkKkMT
GJuhTB1beran2Zmb2+G/nwswiYk8NESnQf3ORvdVRtA+aaadptSkLmRO6wahJz2A
CbkPruZhPelNFY5cd5oHcMVXhQMnp/FP7Ys3/GYfVUh/VDKSNl4XLrsJpXridVPR
xM4L0eio1x1CQkYsjpoefJzZzHchCnXpk2sV4p1nL4SlYFtiubIS5O4KcJQX/fMm
Cvw2oykx3aSuZ3Vas4UM+8yKgepaNLGVbbQ8kOTTmQ12upj/5gUO0DTxXDQ61Gti
VfUiG1iwdZGbhIojzI+13Xv7/mReb+cVZ6yq8SrWGy0xehmaNKRcGxuLdXpigYBN
UcGOyd2ZHcDgmLgSbFnz+mrNJG3lAbT7f1k8KsCVr5ghK5TjtUe3f817a+Mf5wxX
TvwcEtjd5fTItcxf3SkVNgm2uS2lCgGdbgi30XklN3Whbkh/9qEv9t/aWrjWpdEI
Cqn1QbTh5EMlxS4dVA1GTpL7nqcq2noEOV4RpNJw+ajn9V8+Z1jt1C/P+44QmfMG
TyYNaIgvGpePwOlGCrI/AwBnT990jgEG1a2YYfIhcWQg1i0xawCZI1/JxFmWCQpx
u5znBCCtiIon+CJRW7Jj+tuqC7bJnYXTzf2W64cPio8aO+3nKXmL40AodlOXeurm
0UUPrF4hehNMMfpYEIwZZ6GB+79rUZsQrWnNnSa0aP4L4+D0WEgec2TRF9GsNVsM
8Nb/VH8dRHdgWMu361pzBwto3BCypAJ75uCmG9Tmiap2lhp/ZurRaA0XFaBjoH15
uGVT7eQ9cH/wc4kP8hTXt6ZM/wVetIWKFE01S0xItoia3N8WDo+zB5lNkmRS1Nl2
chTBsPvwCecBXRjia2scauFuLfunsUD8wjJjnf8GPrMihto0H/6JcFVHeeSvMH8Q
rCk0zvfF4vtIjqcLMEe7SxpD8/DDGKu3ZbuOFDbnc8G7ufSkaEgzFMvdaEkOm1T1
w7w2I1xHccqrKhAe4WWBBs0DsFE3sybTpV+vAkynujolYzF4ketNixG0pj8gHs/p
6CyL86JzbznZhVEWqaTbYUKzamBfSyaiARCQ3uO3DmgstURnXXK4SpXEXySDlpBT
qVzjDoL5GxX2CRLMvHHAbMVqnPQN7gWYrmDSzYr5l7ED7etNogc8CZeJzPeSltKQ
JDQQzJYPWeWVreZCGeOU2xulM2DrOXF8gfkzVR7Bpm9b3pnnv5Qxtuk6TIeY0CsG
xVjMLxM3qYZgN0dA/3tCgIZTFsxA0LMVjPauEN1pgoWZL50EGTOGs32tseQlzNyY
EvL7cBrl5ng6gFcTu1bz3bckbC7DYPnWkhxSs8y7MH05tiF0tUoxyNHkELku1fbR
MtMJtT8fljhx1FKfHdWm3mKOBR1FUKfjO8pyL1LCV8+ii23kOrQ3mK6gGTQzNuT2
7rmxEM2i2CJujOwQ16NzxoAUL6QBFVUVkuWtD53mBUKNAoqQ4aGXa/cP76wrmX1I
SS22Y/zdv3OXk8lGw4hERdq6G3HrcWVUBWAxf2kyJoqwWIIp4u3dSmxgavns//Sm
/VQzr0mAUO4e5qwp5tOtxylPVE55zGPPoUL9Zm6rXIFNFKmfCKRP0nyZlvmlWeBv
83hjTMVN44tseMbDASfaHpZTQbsv3UOaZcdK/xROaL2zxfIV4ExHoMgKbf3fWahC
aYdSoZCynaRqHc/1OyfmhEhF1UKCbtkO8bxFl0KDjrInONDMTUVnHHF+w0i62+j4
SbSFTlZpE63V/kgQyMqxbzg9oyqmk3m/CkE96T49NkrIwR5jbBu6nJVbOw00xgma
H1Ozcz3by5qmVVljofbo/mCj6EHHS2MSBIzolbDY4PM1cln14b6Cs5XvRFAz24mH
sxIXwd5E+e2d9ACgMz3yuSRsdpTf0Lwx0h3znprr8TXW+sEmALp+cNDOQWUHVQU2
bKf+uR1W1rkdI1SqymmnJsHkoPac15x88+HaUqXnCKgYb3iBvX9dn3zRdfPIx6up
uzE9hiX4o61XJD85rKs1Qe1QqAl4CtXUAHQQ25uQMA98yNYktaJBkVNXTKTKKYQ+
a2oYr13HJOZLWUS7N/rUX3xoUFSen8M08SG44VMj2P4N8moW7Ckjiv02FSBo9Lyz
yEBqJ1pLWCwR0hkJV9aVy8JXEddum5WEdDwhKc/W6vPHQj2nzQex22Z85bHKbi33
ch5ZcqGh6jwBWm1IGbWneLtJzuaY6vn7l47u/o6zhECPuX1KQkAgyBlP9Dgqmhaj
bCmStlC7Ff+zsuVVU+p4OIecWcEQts1EwhjdTSZ73SjXWwoF3rj2lJl/qUPcePvk
Th6bZBA8c4u6RQzj3MN2B3tKV6viKdPj+4PLANKqhJMyeZR2y+Nqvt1XpJD6Px4O
kr6RBtzEJFY4gx2S+bdqJMn5zKq2Xvsoj+RyDT7RyE/3KluvyEl8fSaJF994ogcp
Gd/t0UndyqZaW07tH2psvpzpcR66dRjtCeU6rrpKVAjw5Q0vETjo+hkNTuA/Gg9D
s/e4xWVpJHXrffH/GTgSSXYMyBdHcwGw3zIF6jzv6NHhNQx33QW0L7hHnhEmvdyg
XJhcxGjoN9dmSbiGeSXsC3YLOFMP+KjjiSEjFQeIOcEf7uUFkC/6ExYuo/0Bbg0k
dfrc5z7NzhQMB0gKnjVhL3oH5aynxstrqPlEP2yJpclvoi6g5aup+FJIjW31P4rl
gSQMLBie+LZQwMZHL5MngbdaaU2AEFBRCY7GcZK5JWPIYKhcyruV8MX2QLPHkxLs
KFf+cF8M0MmTeDQUEbCHKprt1OzgFVVjMqs0tLPDqSan96y+SzVpLrfogIU+/o9n
cwW4XXGrsoRlxIzwcBq5wN4YxUwILcp//uCX+3LooggV9ZRVjIrZ1qW7bgtqneOf
DUnAaTJnez0nDLk6edMpmtBopthoS37ZIama0UAh9wZmw1+u5k0389IdAJYUMHmH
YWJZ+EICR7AzFoC1uwQWjmXcr/kbDDKo1M1fbKVs/X8tLgbF5TxN0ybJIcaQRNPC
vBj5i9S1TRhnWwzIlLpgyl0Xdqz7hwzkgvo7XZnVzlmKystdxUwl1ghF5Ihuyn9F
5pL4aQy3XnwYt8BnMWTYso16ZkvIjkCNWVFA2sRs4G2aSagbj+P2VX+QmWSkb8fE
JiG6SybhcTsSgRscTeFtspY6gknLTuBaQoBA3H1Iwq+NQ7l8N7V646xC40OKF/OO
kETNqv7RiE/DvMBI1G2zZAtDGNqDO1QHS4p6x7lfd9/wSpl0WEU2ygm6ANXTOg2Y
RRwgrIcTEt6/67Hq0J7Y3txO0PPNeUmdDpXMVor/0ymP9UzXxhDs2h4q+pdSOm2s
XqNc0i4IiJqT/gh7gfmrJLgp9AjtHOEAQpoRHgWgqHxUP8A8lrGWJTjOvpJPJHw4
1/xJtj0QAGdXfuFViuzKI4aM0V2BD1mlq0fsS0xiSV6c92a9Jefd/XUTMw//V/Rd
o3upQcuJo5q/d2nbTeezamsxIX8vFWOe6f6fZ2dGD3NfZAqtbIyrZrf9m3yUINqo
ruX7ONGh1INLLM0mQGJT3hryq+dXoolNeBpT5ZeEHL3AIG5dfAK53cYhaEUDCu2j
wtKLOGjNhCdhUM9Lx+RgVtcA6yCTpS6xHVX13srCdoBriLQlmkLVErOXInPzUl4u
nO2apqYsBD8LJJ4d2KZy8cJIaDXwPSjInF4nLSihqndMt9qKo+rM6QVmhGdUFEMs
6LNXCi3pnViaRFhHXrfM31CuHHTK6aZ94zSs0dShctCZEMDzRzyhzJMnUCYEYOM1
ywvNit7ialJUaQM+N2CG1V0a1h16kL7m+kE3h71F4125wbIPTrqi1jRMzuHDHVYm
vzn6ukLUB3sNvleCer3SIrs4Q5LpP8SB7johY9llI75SBmZe9+xDggrWoXIGb6ts
n9suOzZsofYlQTgrcQyASXxQrBFiCJefMDqNGvfaBeS802h/FLSI/Sb/NjaK5eAb
UCjMqqgKbKiPETw+COdF5twwKrAc/jLHiHdKfpLzSMWhsg7zF1kWsSEVkDrQdyJb
HsYrqVguB2hRo6RM1mGeTLwEKWC6kYDWc+AgIz8Li3mQhkuj4sHhly8ojFc4i9KU
8EntSfCtICb8y7mkMONysuCkrKfvRyWxd1cdBFJb92IWjI2RPoPfX2YG7vkMu+LL
dO5rVq8Y2CmLdepfGuhBUmI0g/KFBZd1rZSsCWV8iYBlsZoTATXOmzcBmtKmqgIc
VqbIUc4EJyJ+XFIFkp8SvPmNM0miz82xDwS/MWKKEQ7gd32ldXrsbm46WKKHSnnC
gIhbURyXDwNkwyARLXhAepARzPAyT855UOq6UluykvtvyTmQHPVfbtUH+useCyHw
AP8qck+p52DSiKVmIoDDuGB8LNgt1VFd7S6+2yi63ulQ6hzNG4DEXeOi56TMubnJ
zc4h7PUxiF3MMmU7zaQIuOmp8K4LJ1M+dIQhl9SH1TwztyG5Qy4zVxyuX4Arke7w
K3/A2lF3m4C2OG1/Ohl1raj9DGa9sunpHvVGeV8DhpfK2jZiC1QVsalK8DJc57EL
aoxYRjm5Fbfo3wzV7VLHEeVgaPAE2SRlsuKXNZ8AWTdvpR1AYNV1D1FE1yKHAiGo
cnerN6RDQlYx0ZTBS1vSkdOcRo+pbCwkenDd1AVGBsZCXb1worcnRyIo40KckA9O
kF+Yzg2CkawppQ40DxUSjqh47T4+vE6WZ+JFO/LViyEd70sWhl/e4W8E08n6xP6m
MEz6MidCwnCgClRqC6m7wGbYelpr20v0zQFX9pwdwNw0SQU2oOFKyfNbFDk0uwaO
qDyhGfK9cXqecjygQ35is7WgKRvJGBaK39xuJT0nGdvX5b4RCLcWyLPi5aQBFfnp
iuukRxGLXmeGfvU0Lv+wZaVo4tnd6lDn8w269UK24ATjc3mkdsSAgSi91PANEOXR
jo2X2uLHrIjlWCu/sWyUfa/pIuIf9PE/0b7227azEBLwZzTbi1eqFIAm3iJJIORV
0fdLlE+FRvWnPW00rZmS+wvb+Ho58RouyCIkfkwaNhMfZdQzLdt6XHZqaLqyz3GB
Kdlhh4cP+vRi5Etfb08r5AHsDu4NVNvvbjf8plX65gFIq2A5hW573+f20+wLmCEK
miMGNt/4t6Cxag81pjXVT3hbCMRQU65HiMU8Wc4QjoaNl3T75Yje0babo0qiZl02
XK/5z0PX377K621knKyvMvPh57ayGRQH5HrlO3niBzb9La7mO6gzPmVPrrZWWY5g
ArTJM8dhhSbLsnmEUVPw52eQSnTiGjCNiok4kIDV/Yz7JsfNW+BzP/WA6fEPT3Q0
jSyyMtRcBHdjbDanm6OAMZ+nVD05GaOTJS2tINU/1BOuWAO5rXk6jzrm2b/L+pWn
LP1RFDB4Ao00J+mA6jyfFKVzqBgbDTyWJBHRGhlnZ4Jeee7DnkUacl9YAU3xnIwf
OvQR704lMMva1cCfQv/dzF/g+/Zg5GYIBpMPWQkhxiwttt1ijZI4HXfWaTNfyVxQ
L4kWNqgYVky+DrK0zwaBmucAdJJC+M+wmx+do1ptJAd21GYdsUBlfihHQzg3W1jg
jUcy0EmkhCTI+a7ThH56q+0g2ykdv5VYUPIiukGh1y1ZMzGp8tw4ks33fCD+u1Cg
r9cCrLNO40KT3+2ArF26CNsSu+kJpqn0uNC+TRyi/8x1kuXRjnHrdpray++HOOR3
nl7y4YcUXyRfh7Cvc1niaA3tc+I/GGvaVaPy2wgobKryX35nbcWqoaBww3mb2Jxk
G54wP2G9tzFCjW3krJVA7TvhTl61+ExMh5SQD6prF/G7Htuvd/ZW3sgk+Drb5GDP
STk30ylbuaTIJMgBIjXw3rUmGhH86No4geXMra2IwNh6z8/csfxTyRv2qJBoP9qJ
1l4Sw0MgYWkwZ/5A9tYr/s3k3cvY8qAGD7R5lyFNPG8xjxim3yR9ljs9yQxZaWC/
OzyXjakk3HMxPh/9dF90YxjWP1JVMBhtnLFQFBGSOhGhn9fiJhQwWtMUkz8CJ4Db
jM2OplWqeQgfd3X4CGQB5kxcokYHbE3Pbp038ZcFS1jfFVJpmfNN1qceZGg8tYYu
4U25MPNWdA8ZciYUhZQ3FowBSzedJunEplrn7R5QNvwGf71j4nZ77g165G4Ipum/
eT/Tc5UgGhuiOvG9pkP32jA+F6OYfcurxQ7puV1gWM6SLCM4hzpFGOdU79EuCugg
2iIDlgb+kdmZoKQZA4ybvllJWbonjdtSeBL3nYvR7Lzz4vd5nO7dVfK+ZNpEzqg/
HzfvowWPUahZBF3Ecl3hyvjLlyvXS4MIH+QMYcqNNngkNHOkbk123qGNvJjq0AxO
kDB1nUxp3Y6W29WHRENnvzHkNjbi8ler3zRXTouSXO+vvQ8XAbjHK+vi04TDAruW
QODivDS7BTU9mkgpPUdylo2YHjCis7qhyLOd2JgIVNZsDSFpm8zgAcYJpLLpc9Xr
GWzixvrXddS9JqKbbL/GsGmG3U6nOT9PYT7T8yDQwCp8YxsI6aOEUNDK7NFtRtrg
eb+Rw8G2Ivc6l3VDYssUo3oC2VMv7YxamMqutVMa7AlczOpIJ7rWklV1ieucLGbs
LYsWNK2QbtDQQrKCrB/Ea9CGtd8FmqfASEMglrPRpMzFqx8pRU2FUuRVpHctCFZJ
1dAQcYvu/MgI77Ta6H0Pg/4S+dHj0H4qTdsc0cxhQ7+q4F8uJdr2NZSp4GasV4zo
uvyRZvwCfFsdHSSM03o4jrizorxiqV2R/I1HZH9g07FN661M+1p1vHEimCSKziiT
T7UNbud4eXTzITCNfoyaGvXBDfHR8NhHEkVrDTKd4sD8vKIIA1MSZhBitI1IL4fT
jdcNIJqQd6WRcYdd5upOH6YxdVAsteqeOIslnS0KWQj7Sj+JSc1X7scPI7NjhEDk
2BUcNOFggdXMGQ9UG+Lw5Zt9PDsGwn/ol9w/R2pK4utqofRGJNYSeWtPILdpSG2x
YUMYRUUl7mleS3+fgMQhzLLzewy2vhSQlsqqem0OyycD196GUzMLYferN7oAH25V
soGrfaM7WuvkyH35dn7BOOYa5eylSAapzXyeIz4URMOAYsB7ErIWdPi0vbLgaENk
OAVaOGQccbLfbz5p3I4o+NU/mJXWGcm87hWOa7o1yFyuAspX38WibBYv9AHgxG03
14srNIhcmncuFydC128Uw23bg7itG19tRDvibG1PCGfGMkFPKuWWpaGOaYIcQYdO
3tvBPTjOe27qAikF6DoLluDIh7G0GqGmSn10vnW0DULudOaedBumHaBAnMpro+D/
qArOi9Wf3/YOk9Z51fSKTrLvYMSRVsAuTOqb+6xinXuh63IWxYToWu8NLPtBjn8T
Hq8JfGqwComyXVoCej3+oYeIX0/DcdLgmD6BvLQsyEVxSb/oQbm7Qt20sZk2gqY4
JIWAgvkF4IGHrS5HMy5yXwYnYWLvCiTJvxS2HxfYAsCppzk74yYB3akvdegbBflj
GcfxZhhCWvBocE3PzwOqPs5jM40LHkautfQy1Q26LzETeyHayxnbfj1fgYz4m38S
NklNAFtX+IibtKrdmqfcLftBEn39DyTqDlIYAonQcJDKf0naGmIDdkfVvlGrQKZ7
fpakHdYLeWPe8SgmA4Do8dU+ZAW0zRrfqchvlkPyAQyzEktcwM3CARgo3fVbs6VA
cEBwufF4xe8RfS/366xUXlJTkr7ssV/AuAlqanaWkmM3i4tcYTlEIHnVi6Et+r+l
Tx9BHSXNUXzTF8WMIGcSxRl4YWNG67CIZBQwHW2cjc7pJhyP8u2Xqq4t3e94WmMI
us88A30encG7b1UOXxvKVP5PLT6nBUlMeAZh7nARl5v/SG12Zkt1AxqOXl2tChto
lAa0sLf7OkKseav+Q+vSzo1bXw5ZXpI/pZ7W+JYFsyFr5aGo5Z6diS4jMmuCqyLq
6STmdy15rXTYxKFUM6nb2BP+2pjcBQZqFhwN3lSZTxwYSt42F/1sBqda8k6qfXLo
e/gxtFwPx5X/9/FC3G0xhyvSqx2NlzCGGAAmFrm6LoKh3ycjaFjivjbSfPNe8iJB
15UZScI25bT2pH+MOMMR+SjU603ZxIPQ700ZVtZgMiwiaNjBJ/DZlEBHkLxAvIQe
ydXBJq6cQecOiJnkWErlALVd07Q0srHM2EMuFCVpTJrs7MAdgfj+UQPYdvFKwDCR
qpPjrUH5LLcySosdLCCWYB1YNUfdJ9FZthxtDDKDvHQpUrxhbIKVY+iZxk3oHQEu
BquzC/rh9MHkFt6xoBxrp+K6FHKx+25S1TJZfPPITPiuijg5EZvu5K8bDWhCtmi1
2F0uflEyQPgjPwhTKuGiP0nOpt6rcE/5Mk6Hb0ZEDF6ic1EsWgc92i9s9GQpt9rb
nk5XqlyAYLY56j/OYD2ABv+A51OT0l+6k4rQ/jPALfGe9k52RUvf6SZQ+Oklxv4C
4iVNfZr1Q9rkU2psKTCdPtZri6KdeL9/vXQA/ERHAr9zi2JYIzvTwMO8rvbaHizo
irFstDSsTSOg7ph4sXR9wszmmr1esCZAL6UPk8zqjxbYqAKS3ErDFEypPOkl6iGe
jGfyYpwpXe7v/U3KizaSeuYirovkFpIIY4zhpY6AlBbY4AIg2n6FQN1oz94+cVKM
3kGRDNj2OXSJBokZWEOw/OGracBMAPZesfm6jjOTUjiHlQTdq5jhHyy2XjLhFWME
sKMc42ecdJXqj2MIEh3LvsO8HZQqFST+j/fJwNAT+eWXOL2JbSZPu6ofQGZFzfcT
8lqC1E/+6mu3HvFzlS9nt+ZU+JqXJOXqORov1Zzwd+pebUCztFnIIUojNNS7apC1
UmxKtVTemJPgaa5zzM4YctA5wWlwO7afIDb/99hHJET2Ap04JGLrV+F+chiTXVQX
jARxrUd+Z+sb5/iEhsuKj6m8QDWsnaRxVJBoLGDt9n6tDxbHNgm7YXEMnOXVVoS9
wcZAqjjmvXL/ttGGvzIOx34yEKwh4rAv/55mvXE1GuaeIik7ztYhZmbOdVdFCgxt
yd8q0G0cx2tK+sLngTXIiSVC+hbFRMgD4/n78PF/CyciZxNIxQ0sGeOUY0TxiGUT
prlD8E5woqNW4lMIMh8FnKgan8KIo3SJOBZVqxfXmGhq/UDLhCDMef5nmz+WOOtz
dVQLe0iPHkURNzyU4gIYrZer6f16ADNBWrjE8Mtywl6exRGiPt3R7VmTwAILLUh4
j/vZeHis9q2p/XDbDHyoaU7OJ5vA5DxvSQWEVVD+JW0ddQVfnSwXL2Fskc6iv0Dm
k3+CjmG03MgxDx+oEcYRKCoBAZf+6NTss9dExT7qyryMiJPQCJDUTLLrgBb1UoL1
GDN8A6UyPRNqa0juyXPLi7HzG/r15Bs5IE5rUAwHEff7KP5dGPs2LSSYwwMPA/vE
Z44egp7J9QaiB8BtWaOmQ145Ljjiv+CYnezCaoXWMaxNGQedhWr1ZK2A9rYVgfF2
gjJTKMpH0mlSTOrspGPyPXubgN9oDlp9k5zSI6apWP4/JdSCBFJnkxDqhX6wuk2Z
QLc6njHv3dzZ/+e8vGpYQTLXUVwjhlZu09xmdI5ZSkSGcu4htP5LAPEXurxMMjiY
2/U3e0iS2xhw6vdzVpTY3zhtXmPeTpt9yZi1u86jhdIZ1CpMq2RnlZXSdV2R63sM
jPbF9MzqKxS9M7x+HbbumKtO1gDK40eX9sP0Mfk8IvxpXUmNSU2YPMbT3pSlyCWQ
ZpaBdIy6RprdM68xWzBlGcdPNy2g5gWHiSzxFWQRwomv3rwcCotgVNHyEaGTyDMG
ikv9P126dD7mlPDHEiefc8sm8BWV32bhdONO9CVr+3nzzX7Kh23YXRXQuKYjrSaR
+fj9l4BvZonsFtiOy+POUodCZId/0ML8p1FmndmLC8Xmm2cuijKSzC+fTaE6Zi+C
hlVsv/myKfiAs1LHqsEc7Twp8i5XqQTiOhbAT1Xnv7lbUi1rMBl0I/sZgPHRD39w
io0GMYQQgVtagdbqPO0nU/ZYgCY5xGtGPbrLYtuEQRBO2SN0wmv+XcCIv1WY4Ex3
V0zFlh30AwiD40GKnH2LWZ0ZRjDogHn0a4OjXG5J2ICc1VUo+TUqxaHfrK7KiAmp
ngksujg393OO8omSDPRMyTf38hKPvy1F00tX8kk/uRtGvR3KQr3rSVlzNupqzqqa
c0/4OcurM7aLEaOz6Ddyv0PYHkoHQ3sHF8TFqJGygg3ggB1n7DQ0PqV1jgRISX4E
Cndeo5LD2z3mO2+8KuPjmNvQp2peNK1Gj4uDPhBX80Mj94AV5qIwSJ4fZToaUdKI
1Av9cu+UU8b+8hA45/rtCSm1F8WlUR4R9CAVH9s0U8D+BPWipqQLsZ3nTN23Gmvu
mRVjWYopsDeatkul0mUTRds1EPHZx5/ErvyddaFxuXEl8YJbpkTFQ95l13Vv/RA3
IMDkR8eK3BlVn7O1weiToQY4XftUeHOgx5z18vlxSge+VEQB48ZsgG/8dLCbZJ/X
WvNpqgv0kyREMS7tjw7Y1cKGwqneosFYp+VYPfd34Ymp+gkPHMCiTEGS0YwOltqz
jnlqqdITVop+3HNjPhyDnxC51sN7VwL1s97sVeyMawxsJTKzgc+ziwCE+uwo4mB3
PM/7zL7eUxueMkgZM2PJptsHj6DuxEJGqRDNFHhOCQgBxmm6NiuzzThgZGSFz9xe
XEfy2oIT57dqOIFRIunH/oEYsyoAZ+CLj472YWAJNPeRXNxY2EMj/9BvmIatfbuY
it943jYLce7LT65Ty9ND3MOaPV1f5PFYvfIFKxOxPndRiqGSKndPn2o66oTaFjAn
87cXrQ4Yw+CUp6cw1i3Xs6kVdBjpGA3dN0tTjXSaJURhJfcauufHNxOgP66K2QjX
Y3v3SRv2TsMjVDmmi+OTUrBRalP9aSKq9N/shbfojC6WhVCdcNyczCafs4U76rNV
hNN4pRbe+KxcwLTSSwVhPH5A5O+We4ujYe+qs8Vrjr0D+ILNtzM2wMy3IGqVLnsl
h/EAaqy5sgtumcZp9TXNNefuaKbnuqN1zXz/XcmeXy3t6G6gSklFrk3TNVIoFghr
NKVRao32xYihb4gsTrZtGn5mAGZbj6toRzDpTCyxv2Xz8H7FpRKunr412/5/Mt3V
dyPmTtYcAgRtPfN7VU0WlEXx4Tqf37yNxb+oo+7zO9LoNX9Y3mA0skyQ/NIYF7fm
LgZrth+dprlvW2yAlFYieJvtwsmpvih+/+aUWeTgRtLUwj4FPKYe2mUHyhzOlAdY
g4KiYYHlCXWo0Tqts4IOvL9gHbOb8xWEYxbvnIK+xlduY4H/+rb1LapsoJ052OK/
BYvm3S8YOR0Xef1saG36HXytv50G47rSgQLazf5HYvFtMZEE2XNZdhu0eQJMZJXp
b3yhZ2PRw0uan3ZfA4bYWSEPDBXLTTqb08px4rV5iT/Ojlq+ShvLBxqrhhvWL/ZZ
8U1bk7morrnFhHsOOD5N2nf9HmD8pHes0rqPcHbNZBoyM1KBvBoxyqp/pNEc8fj7
JBfh6vz8yhGOjHez9T4wi7o1Tw7dbnTyZnghU8ZyqDeDA8jVHUYpAdm7aptlyw6T
eI6g5kAg04FMcaJvgNk/031PW/zS+yTXZwablp+bfzQppnfAC9GzeMLbpi/rUH4N
8o0aNUZpua1INOsy3rmEUplxBp+gHjRWmXlrvunhzfu2SLZqNSZgryrhx+X0aqoH
BOnK/rkBq5BR6Yd2RKkONM9wn9CUHSvbvywsswvUvCh0RMCYJYso1U9idYuJA7ob
DcMppzNDLp0Tl89yUe4c8jdLpBM9YPLaMwB/a5cabLXHRp1fPx8R9uHp/wEXruFw
PQ2uy1wLlnnwFFhrG2z+3P7QUNtUYWKKBMSiNCg8WNBXqpNz6UWPxKGbKPhSchRt
E8WXwGyCxfOicdbMVzMY6Bus2VkADt7ZB1KF1kD8oZSGlUgzw+lOCph1YJMMU/Eh
dR2gGetTyb2cx/Wi2mRmjFN4oPBUndGxIuGa22Y/Na37FEudBCxrOn+T3enqGI/H
15T25JKbmK+eanj6xTEtiUBd/3TlZTeJkcvL9tsl0cxNGiJMcPtG9iMTe/GkQN6o
DkMvj6Rsb1MmIkQuL6wOOsPYQtw5F6ekQ/3WxzrwHr04RQYhmAxs0HJQpMhaNX36
85xk2+66nGODVPC53EArmfiInYdhfEMeFbbR98qW7e7B9QBNagiUgw4HI2BEksxg
bSK8z8bl/kAl0AlTWTH8gf99EVR6Xj/SAVGYoVqfqR+xq6pUzqeyMfHQuPE2SSHJ
dxD8Z/U5jvcs1/7zTgvm11tQFUaTcp/hHvKdQabf67SpPEhpgcsi6KB6g7wR+7c+
4Oi+HMZNi58TkxLM7nYTgO3jHhGmu5+4/xwn7PEiqFRy/nsj2RwBfwTtzq2/KiNq
B4Yfd/pykHSdlNDzWwvpD7OWEGVandsZvYuQUvTUS2+cOJsTomaY25zaTE/qKhHJ
Prom83iMrN/WgRxdM2uFStfG/K2pBI1pjC0EHF7SIJTa5RJa9GR2El4BBBOTWfQM
InOQUCXmgEfstHs+49JJbxB6xUYGEOSQ77x4gyxvc8ld7muGNIFUX4sgxRg+W0Mw
qHVLbaK5jd50sdWjVU1WiKb357CayiYLpZLrDfwPCrdTDZcHGLj//oh/r/mBU6wM
vZPhhxiAWRfsnfoMnBqrpzN1IpidcFrwIneOooi3P/K67jHKNzMfCniGU5ExGLsH
q6H/2ThoB13cR0rzaf93q1EuG2kIuZJRAjfnH//u4cnfjXQ2QKcxWm96vtQAGr8X
EvTUTMd6rLfDb9nOlMoZe5ENzyj2DOzezj0VZwcWAjRaYmyxunS6LoPB9fStTA2Q
DvUTphpvuo9RqvS68xVIVjK200iF5PqVA7KmuTs8c66X/Il9kWMqXz4m1hGt9X+Z
d6XX5/yQi07akiW+z25UcyfKRuswrndJr3AdPVFvcGRRYRNzWWJ76O3Q+5PH5Llf
H+H5z43HJmLID1Q+k9lzySqJ7xkMkPXfZsuXZgG6YjzTYvm+YAn+i5DWgFbSt1hR
d26LLbJ2LPbnvJecja4rWPOumytE2g8FiaKIFx/jOi/7/70bLZxGUmDGDKL7Q9uG
/tIM81OjUBEiyfsocrxUjG34nuGmCTQHMMRzcu4XeokKx8g2POV7Qudj3C2YW0QZ
7kGve0PCZrpx06QEOlNaOP7E1U8smdhXlRklv0q+pXehP3jY90mnR8t6AlUYDGde
p9Pdii4n4698A+AsslkPupr1rarW9rjVJhoekF4U6j6hG03SqjeWJpRoGw9tq/z0
bxXmd+Z7S289wfcyzTF/TKjyPm72DEKP74qVif5SowpOXKcGhiPKbeGiQ4ftwBOU
MxQnxDRmYVp46dShOVtILiwh2C0EkdkoaoRvwImbvksTimkeuTuiNW+Nw0XM1uAI
3Xb4lbknQOvzgiIET2tGsw9yuzvzTvVORy12l9cBVV0pmLZjr+KGUrT5Oi/ihSIF
uu4FoAzGoEP2V2wMwC4NisGCTe5yOPITVuds10XebB/5tpr6CH3+6dhFkmQyQsv9
iHpVhVnESieXGmgBLO4Ac+J4xUOUXP4hbT0CbhxQpkdJTT17tqZSfoThWIvdJLPm
7nxwHQn2UL7OgjKh4IqzROpzNQNte0Aqn0TpY7I7Y8DQqvDP8wCBAN4hbQISMna5
LacDNk/1H2e7Ee8OeCbcVrEbQqwS0b5ehgwToteFjASq0V6hGMEYrFM8EuEHszd7
YB+HW3s2WtasJ5z7ahHfGAehv/M0cCdCywhLNbctMetR2vVC+r/K+OREEsQYQ857
3k8c2OSSd7ukFF8V6kwbi7JqLII/ByZ0Nw7o3FtCGdddgow8oCo5LytJ/p6LNJpf
dnC4BJnnBc3wjhw9UGPJtoxcRM6PWIFCfYZ+x60V9p86MaFhf5Ke9rdI6tdmWl7r
BZQ/U8/D12bYQM8wU7l78ag3SKRyA7wIYkhOla9P2vevtESDlcaQiGHL0mMZFrnh
ty8ktjE8PScwetP7+J55mK1lsmCB01eAWn2BPyd9671u62C1IQR6KDj6z7Mro7S+
aCa1GYO+4qcNNrEbvyqCfDMIM2lJquxz47EG+o3SlS6b+RdOJnZ2cOgKjVF2YeLB
lxhXgIh5YipGYLE76rR8iQ8QrhJOy3KfZ+j0N0vv/2JDBKxLliX2SAtVyCThZ08s
MLTdftmnn0WqdnfdfBnRL0DEU7sfUK3YLkMqIP0lRKvTji8OnEW3eRRnnVBkVl5d
QZ8pWIQTq3dB+1tLAq/872AOVqMtz4ZSWTsWU4BJkERYi8+QzvHItfUilwYZMbiY
/yGN1P01oHfZwvBsdZpHixRJnHlCRZwPOmBzm98epGgx9fWun6ssll5T+7mgyzE6
vj7tZRULMTuqCMIUi3TZwDpPLRW2KW/+bftZXluiJ9TygwI4IAPUfNQnteYbHRpk
jJBfgaoOMPt98JvGqBpncPWrwRw7forlQLpQoTHSDMYcoGCS9/r0LOI25TyF4tpz
IELB6oIiWRpkbLNU97+CUYuHYYpFDNkowx3hIqljPEHlWGwOaALF8jqWKISGoQj4
59GR7qBDFP0SYpiXLagA8SDr83YIMQuO8ScG646KdUZK0fjGpuiVdiNePfye9Rnt
Pwx5a48iOTKpV7wLOPjvwKH4903SrjW27JQEy0/IU60Xi2afbsQDzMNXj18NYL+E
yvwIQ+xZWQ+Jg7OYMgLL7TdIazCGoxUAH3lGKejQRiUL0jdiXclEvMdteMkL+xox
bdPydsmzNmTXDo2cCM4D+MRyt+pTR8brtmlcXUiDbicfAOa5Frcnn+dICLyAYFNp
0kO21UuWvYCwFMiqX/d7NH3ua12NIMvCJksAPWO3ev++ndWwBB/4FDsKugsKzoo9
q2r+OHURMq2Xr7o7GDV1yTIR1PAQlPiHJNVVqvaUYJs+ZZwB96EgpVj3V3iBQk42
gAlymAMX/yRUNCE9ERSMedTQNk+dSWfLWRWr5Fub/uOtuK9dM0KH8SUna/6Zr6Cc
+GnRQ7w9GRz2Yf6vJMf6LCQLNA7i7stglOqVcJakVZm5/T63DxtQzhZqvzV6miha
yIN/1utAvvFxtwEob9CzEOvgO9Nwzv3S6NuzeI3/yILP3Jwm4Dj9C6qrpTpWv/+Y
XN0U9vExBdshUeFvF8AShtC1YLftzx2pA7TLtsiVmnryLCaAX6wRl3imXjYA/FoC
gIAOIPrPtN/hlwqiMsUq15OTArCZL2zA/61/4lL2FdN3gNiiqzTmajgPBALI7VNt
oL/v52EUV3RcqJVav9mY2yMPeg4P1TnDKU6TDFthOxzJ9qrzFh+TcPzxrUBJDP9h
HU3ztdPN/0L2O1aGfavn3Zb2/RGZ+IOOQVrB1rsgPLmkA9H27YgH5i1rzwTZBqW2
aTUyiTioYDwADgxc+bThgWGVz6Ch/9H94ie5PwKOKNXTiK/ac+GmNVFpEsNqThzP
o4C2quxi7/kXRz9sur8sG0/wVTY6y+c7VMJhtjp0QgV2iRwv90mAimfmGr47Jwbq
NDd/zBzInXNfXJQSMNnC/mEwSgOP1Z2FEco5yAsIL8rDKLOa2pWQiKgOSd/o2nWY
EU3sudHDgT+vXiYZ+KaG/Jdz+e9IHbWfSkw6PDfvKJFuzUKrYKUkPz5lFdTZjkxG
G1l87LWk3Bu6L2fxKWkxk93wFFNlynwnUecYrZOR1tJnke7XOrlQQyfsDdtDEz85
8gDgdWL9pUeBeYOJ53TcdKmatJ41hXhVQkAu1EYhS3hMbd1jt6XTgno6x0aLF45Z
31Am5UvCQZksGqke2G6uwv3C5rY7yr05HtUEp7Fzilpkv35+8UCOKqDlZm2b9ghk
FVUOyn/EgV84vxcDuykrIIu0NO7lpfCfLiJIaMe6DzgGlWL2SOYo0rTSb0hNGiB9
5GkxrXSvvJeULSXT3KVhionA+FKHYDgUwEWT7FycRYcm4wkqEfg6rEY57+wew/qs
RMb1bQYQU0akshCPKWUFx0DR+P7Y0wl65W/yulLm0oRZaOdxZq6cjr0KogCCPGNm
N7LRMWd/I+pgmlxxY2nn+vOBiXd55efJALQ/H/tuAckkQWTQbeVaaPRc38X9+YT8
V1dEtETi75tXbpFXSM62rJFHqDEjegkJ60/ew/jlgJuBRZUOnh6R0B+xV4osBw88
x3Yu4GPJQ4TW936PrcbqnoXmPGLeP3NM3KYTjh/6to22o7P2FMuUsFlexsZtiYn7
MvHlQPd2iaAuMSBLs8kAfMMqgeqMME8W+fj8kIGiWoLG7Md/IYaLgDAqas201Ula
mZP64MG8ZKzyM/fFvUUts63Uo+hDOtkCxPBGsAwH6XJS0lVQooWifOYUkRb/QfYU
qIRxV3pwegfgm5B/8bKB175R/bmyGX9zdoHj8aVt2k5NP+UFT/jaerNoWGfDXy6m
s+YSinAqP6+84OK9+xr+UNA1nsplqLZu6uPvTPGJNGhKFtAU5u3JYrBgPtMyjmTM
4TbbufLCF02YCEsrCmp+1c/RvhKYw6N0YI7Ab7tzSWjLYWwEfjGlY218eV2VwIlp
4JoJa7soWtBRwLCLJkS/CMUFmJtYP3xI/C3JQMeXfooWg8L2tb6eh+XSJse5pYeh
DIm69nEG4rUNZcVPWtTFAXXZFYgW7m0EIMl2oz0JSO0EQV0lisSkZUEqvcv9aISH
1CzYhnkA4ypNau3Q8N30OIgQxWEGBza8LSZ12+jEGDhKPP9amYmLJO4GEn2SU0fn
bBD1s6V7zZNgja7wnD55PZZC+gh6TlV7tSRl0VoeOOcHz8UC9qwOYtwenNifuEk5
ctJFalPpFisMx3crfQ1wJKBziElN94jc31dCxDKYYSD5RR9r+NpfohdGSknwpWfB
+CIOddbd/CyvDuhK51JGxgsYWnHF7C/1NvSW9QVXUwqDpQSoUtwyHRhufn33xJV8
QRelV5sGsJD6CDU7T5zCDGpwlwwdhmpgBuET7HP+D1n4kaxQ7Go58SLQi5OJOqp1
jXV1UQrk53bzzemyKB7EqH1kBE62Nq8oB5PfUIF3qADENfiVH+9GXxGw7Gmj5SMI
pGBvB1lE5t+hg2JtMdT8i/VRfcPuH8OfJNtx2sfXuzMMVedJEDt6kIZUCP1kxUnh
JYoT+HgH3oQiwdpZQbcjk+LNX3MFxaB/aj8mhBmX0e05d9I4yjljZZiZ+5t4l3fR
cDgBBzfcqQsEbhxYpMQKTHKkMKFb0u64G25LqEGDY2NDWgnMV+GCHTheRFN6/EG1
R5zfKwetjQotJjDOESrt12CrnuOVezwKZROLbMYgSarjMe52wWzXV6fDCLSOLLf1
YaGJtSAlrvPLKF3BQ4iqMeogyVG25iPnDz+Yxa9ciHiHpudZ4e5cHrxO/4OEZVjR
D17Y24InMdgQRZXRNgXEkoi7WdvhhLDv97izTvoXHgjsSmiPmla5B3Gt4CBiHglc
CIoMXwin0rzVoVUrpCcX4irJoYu46asT9aUsnBIrhTm9mkxP3PJSvM4xvjvvMwUc
MkIDZjIeJsYWhRtjWuw2evHvZvv8lez/v95R2tBGEMA76HVXCfz6t97qx4kmlBCo
h8S3Q+6bS5c+Xs17ZP2M1cuUZ7n1wAVRzI02LyDZggjMJ8ViSXGBM15tSrubIY9n
XFr+W/bTiDJNQ6mKXTbutIK7ZqW74mocnvbskfc54qwNRsC3vOKg1l34iS5hXtaf
+JZooVjQz2poIKKjtDkBO5eEYeAzNo60wIMq/2MqOGyonagHU99uT4t4YZF/v3q1
FVy8izUJY4kADmZ4ZUsJbOs08ApVux/5Axlwb+eoE+WIz4XIDvua5ORtuiZchrcX
mWgLJxVTgtugHuaXujPHG/q4T5chJC1hozQAzWj3KmLIdpRFsW/2sRA41VB4AWqd
crYK+YsB77wRcmN+YP52aHoZdfqSALM38kA/+/T9C06FEWp30wJMDmJHuIISc4Dc
hdk9QSbEj/mWBJk4f7AFyN9+WDbJtSM+M+XFG5Wu33EpllK72pVYUut2B1/2xhjp
FpTJilKtPV+hyVUiSHjpDlrF1jiXWezHctDRMVx6Ao+SX4QNJQY1Uq5L06L6fS8B
m+hB9Yp1H/iohK+w11xuv0Afr2ECcnRckn9xmseqoHOQllQz5emtjgueQ8d0b183
R0NGP+t+XSIjPXIMOpfEmElStH59hwS+Yg8/3IXu4QpxftDfb3NqlTu1iHben68O
AQ5kcELbyQwVrznpekdES7gBE1pH59qW9LB6JXsadb06IIuYhmFqc/sI4SpZEzmN
QLyEMCNZm52M9VEUiRuK6trSZbeXmM0+O6IAwlNXbOLc40EnUFT0w6HTD+0wsBnu
HlXq84Csv+Cc44BprIdPWNn+S1+452ln4MJCyoSzvLFDpoquXaVgJnU/iEKjMeMw
YF51DYGL6V0bH2DsKkQkFejhtQn5jw+RjYvgGLnzvKgCBALQWX3wKtyDZ16bGJcZ
e7cMcho7kQWl9NoU8+oWocXEBR3wt5RU26smj/hAXZu69FVNK+24vgSE3ctO5qPA
LurK3hgHY8QzVF1NrJqJE/KLdGgbRt4EzXbU97DVG0Sr5OrNlLj4wKXzdoUeP8HV
XM9FoAjA387T7pncm1SoQ2q9EyEwOF1C3lEkPbdEsJUjXdmyvIxZcgRhuONRbodd
puB81kah77/M2Co04Dx1ps0msACAYbY/9z3+Iiz9N/iYFyBSQOK+aVGn2FS8JVWI
TWc7kVLnWX6Sn2EOl4tP7vO78nkE13ZKgsNBeurfV5s/vQxD0noOwiBLqqropvar
M6WjeeTWCply6cjNkqwuwrWcXEixS64In44EJtwu0v4frjerMa9yJRaCwS0mNAI1
D8QxS7EFyGgQ7VfQ0Ai965x+KNv5Dl21fRsmvDJQW+/M/ooX8uiSu9Foer97ai5n
uMGRZKEU+LUhkqWzpL43wemUxWCdzG4SvGf7QcvMaGefVBu/7J/rNExIaGUk+n2W
bFV+didsku5xjGGOKH3hsx7oIMt3f4xBKiL/wAynhEDyMNW253x83txSsgZ5Qjsv
uZrtxPunoh4VXmmYtq5IG16L5lqar7onthG/R/kBE51GLV6XdUaAZDFDmmlujoJK
C8H2fGIIJ9vR7DUnGDek/uH3uw3Vi7B2BjLl+MCSY8ic1VJWAwN1p7uqLvHtkEM+
mH67Bmzqvvq55T2uEtGqoQDZB0Hm7MjgXomf1OAedz70mowOPUlKhYDBKiYzj7og
OEQ+t33PcvKn2JmWAF+X4Kwxm9DDBW/UO5t/bVr2HZMxUZfzHK8zmdH97rBJNsNE
J+9Ba5aZ4vxnDiVD20/3Z7FnVd4HgPSx23OSSdCv+G+WLgc58+9zmLbJaDY2RJZF
ARc3IBkgCU8dTA5/pW1I02dTVCn8fKdi5iQNRLpn7wgKaOyuuSCV/IJ6GCiivUMx
Pq6T4608Za0z7tH/9rK1tGUNAob3zb6xf4uK8VRHqOG6owyFUwo5rNyjO0O7E6P4
Gys/06EtMIB9655eLmOhNuIsln3nmybOhW6O+1cYsIdJHjNpZ927mPRNqki9PxjN
Y4ZunKUmYYYYqE5WjADMcqt98xn3zBhARHa1OIcEsJJT0jKwpywXHwm80hpbM3+V
zLc2Wfp2gLL2cgPoWOtdPSq4y2YgNMXqd4ivPObB8yUJpxg5YSKXYbt0Hb6FC5jA
a/SHdIJDEdCg+oZvDc3L844xRc8unPTI4NfQUKh3OSRVm70poMCvIJne9HkQEVer
Q6KpFBKy9DFT9PVd9MyMlo+Z+lsQ51luOK1ktLC5ZXidANp6IemwIURjchHvETYj
UickpTiKQYkvO7J88YCHo0GRZvRcYlKtG8k4sXpxXb4aLWW9CvRg78vpm94rNHM1
6nlCrHdcr3rOlA0pqMgpmZ55ib/ioNZGCRd3qrDGEm5iz1IQBhlqdeE4NOOHo095
MDyLmzJzX+G/L0vNxeiXIv5zOtElnNnSBurkZJjt7V3AuNcwgMrosaF8I+IjqPS2
yyVxRhD8rS029qtoZegUP7FFAJpzEdBVB9NNsZVWBV2XDE5URrZXCUTLetvPQT61
8nccFnRrEKaunN67OHVcwDaAKt53oF5ZivkrqxbnRroUTZy/r/PsNK4ntEqJiq/P
jFq0dCSc0dhRQ096ErJAau7837e26q327Ffa8SfC9cV374BW4MAUNhMz4h0/3O//
KSvI53YcDRyCCJFmxmEDeskBc8ptqwHXMbwmOSb1TkpFBwDmYE8dsQU9vvQM6fn1
ePjzmHoTd3EQZyDy+7J8+bbtCeYMb9tMr6zybJasWozawW9Xd/yMX+j7TiYDRLvB
HKA0cSTikoEJdPhTneHFs9o5y1iBWMx0BfFMLIXNODb15gZtoASmC/GXPer3JOoB
XbsbHbEGLGnzQOQmob6VykArTTFCuwgpha4HImrIFRDIeH7qx2Tq6rnLX4zTHCaP
GpWF69FszbMdnPKlM0SMnnDkgsPK2NsWQUnRgfUcrbukCsGjY7AHmOYZfqGBLEQI
zqDDFXiz41xd47yW7g5bYuVqCBFZ8lgC6SRvsgJGproWEUVjRvZMEcU5RzKMD74/
F9BwU1UkofkV5UascN7/oS6OB1QHl+TX1CpD0A7C/kN6mWFnqarIBoVTE8xHOJcz
KZwTkQR/xniaj9xNCQULxkhSJNnBkTW5/5dJbjEpeZ6I3KhIKxGdgd844rP/TDo/
Yvu3oiyKxU2MObubcWQHgq4dbBKIRb2Nb/CxaNMHzhnotlJ5Zj9tpCbZtQ/mBH9k
gAsvcF3DjGxwDRt9zWif4qGll8TO4YI1yhuzJy5AgIiqL2Z5ItvIXlEIeN01uN/8
5T6he59XuLbBIjAH2EhvBEFhwEL0Kd8EKxBapaciKQUGgWRorLGSthBrg6oDzmc1
Nft1jQxDECgj5gN3e0aK2F5wUJw9mq0YdecPthsDHBC40fLt2JFejQspF3Ymw26O
mUUBVrRRLQA0rjaECRrWwAqk6Ugxu06Z4JtCa9IP0SyHZaoa8kEA54qAP7RMCITe
2uqtn6UnuRBLhbR1Cr6XpEhVk5FIfyJ2eRBMldbbbcfvGQqyZwQxs4SLRuBNYcTx
bASIaoy+fs2641aEtkZVLJKZlDU+R0OEMl79JLniH7+bGugjM7PD/4NjoiuDkI65
2Vux6izBoWIxAyUv6UtXtCELd/fovV+CDfx59h3K7d7pqCc43CoOZab5hzpMYwhG
Vyak5lXd/GS2Spjhfb6IvHM5JwxqdWoWjez0KhmGVjYJRV5IQxNhXMTVh740f3ta
Ngz8XwZxwShJ4FvIaP9C1J/8lfAWiab+MiIUZ4/AX9FFLJkMeDKr6hIvEa9xcj6n
TTRaXNsg7R3GvKJPm1uM5/+M1a9WZq36LmBjae1/vvxCQciHbL6jirgp8XpusrDX
Y4S8Vd7CLfJ1jHryel3RfN+7wZYzUUvasNjWGTZEt4gsZ3Ic2ASk6Tsl8C68TtK1
CULrhieFc8/iOze2qwl2/FcVzKRPzgYim9hXGZ13q5HF2NKri8sD4x/ZAfA8puSR
eGumw9YmKuObzp+PFtyFrwV5/Dx5O9qovLiM3uYbAbMk7YgPOtPTvyVKM5BTnTUf
M1aedoHnbKqhWF+dpDlTAr2vFBuC+Pe3RVVxEURqJD8tMEObMPxs5hVKux1bT+Rj
zKcuKqhkaMI4wJwJ+ME4AM7jN4SX5TFvcaCIigBMPby9m39cHXJUtoSCI9VeGG7u
Oxctffq/XsvlCKvZvgIUxh+p2OgWqQqkLv6wki83s58KAdtTuu2CbIYMLRuHqPJd
yJRaU+6UxbeIOEa2WuFfJzzdyn9Q4OvIkxiC3MpTW4JOcC4jzi7v8uQ6snwr3Ahh
CEkQGWJmcitvD/H410vtzOzaL0phcD3T8fF4z+v1Uwhlz3tuTdo898PGxts+fn9b
6MP1NWknGwuTQrNvSTG8MabF7SyLdSZG9TrHEON+fe/hviXeMBUlCqgJ8wbV6lHP
WAqs6m6oFXwqBXXNFWUNYskHjqFT8Ky8rZWlLC1VKukw311nC9EX0P9uKL5WExBO
tUz/Etf2cn5S28vcbA2fWDFnLpq3ZflReK1IAgdzcYXab+ZrwL7kb+tRzkL65zse
ueGYWWKb2jU3X/xJEfZj1chyz7hQwhe9cxDO6zgPMMmv9+W5zPuNVPMe9rpo7zKH
oLFxT12ZeX0Y1gp1dDxpXuE4y4JmW9TSzyHfzAT0I44b+UE8AnMLwe7zy4wZLsYT
jJ5Mqn15D+Njehc3jHfSmprQ+bFYM89o+RLA+26ovEeNN58Ex4PJK6qSIGt52srd
IA26VTVx/l5vqKUAbZzg4J3vDKncXHvZzWeyRgyWkp+1zekmFO80gxRtz1CoF5tU
jfIZ/XcjsL3M2TTvRlj2Arh14fJ6qA4ChG5SxIWxppU6zxY93y5pJ7RMI5ip/3f6
xfGva+QPwCJJhVJWyOIAqFgJoV5bTu1WH6FFPD44xHdefX+Si9Crzg5AN0ud19mk
0aE1Q79bFdGcI6aU+oReL/Fq7Ya8KHq7WmIR0YPD9GeHkMUHf9oAIpmR7mhrwla+
qMMJ7N/aTCQOUJn1ljKciAQ/zmErxC+JV4igWazCsbG1EcKviZG7M+lF7v7aZtYn
X6jNSvRTjvoaxNyAB0Zsu6AkZzhoLV55FZC3wjiIaTlACWba3eYa/dIFeJGGI1NN
VqRJKpXcwWkLESVLMNwe1kxGUa2NIEkmT8HqdAYGLw7y73PRrV+uAJSXFkEQpeQg
OBpRCFGq7/yJwdtRlH5dELXtbKwx5mFc4wC97WPWpsgTYXvQ4Pb0pVlKoTPJyXRn
O7SeGRxDd/vPMlYk6YlXGDH1GhcZ5VLBRDf+7kVnKfS2TgUiAnbu5sr63JjzMKJG
sigpVdUH9uOOe6F30JNsNBS73JKI7OZRz94Kk5P+94Wqt3g2jK7WcGjaek4KyN5p
7IRjcWjbMKfSyqOCdiHOKg8A01SS0sbCSN+7QDDqAuWzp18W+PRSLSfILV8d5mdV
ncpTO7H/xDgJZeFd4E7FcguQN387218wJA8hxL0zwZmwOazB8ya9UUYQ2sNgW6I4
ArjtuOOr3Jfp/lApTMUWmno8PGAERrCNvF3o/Dj6v0ePSARpenf69GPKtMHa3Wjt
d7lvSwo+b6HNtPpGEw0DYMNFyObGpGq45GZazoh18ClJpIQ7I7aj3E5cB4iVhTpq
EbvRLtkLdoNma9f5UfIUsoiyiHza95dxlYftAqn6OVLh6Bh2OyiQT78vj3CMng7G
x7T1DZ/9xFQXTqaXryLkr96S1RcH7Vkw1mEtyIqnTT8T3E4DadeqfkOyujsXj7b5
Jw8++9re9tlgEzSGYmRg5t5B2gRZ3ZTSfOL1QtEJsFoWvyNV6SgImwdwN7l5l3Pm
gSNPKGEb+r+xlqF1UPi9uyF94C1M2kCzFap2h4F74fUy5vhNKUzycTQgw3LkpNwI
+hNTHIFGkvEFAcs4Hc3Ivw+LKUZFH5aelYOYulq7jt/S61rXAQV5cAdB4Um06MG8
FgMcUiwCuxCRzwOFrhFG0foe1cXKwcYzNUoV2vwzeiz5RuhWOVRzqohO8VN/ObSN
E5nKN0LHW8RDjyih75dnQwfR/yy9Uf0Hn6rMI9NLszYydEP0IZyjUHfn4iovNg9X
79zG8ByYoij9cGLZhz8Gc+SHcJUJRwoez0bWUU4BorG+0duDC4bbRjqLSgfNnXBj
5aub6daPxXboGxyw5Q5lWJ9S40TE5PjaJCEhHiKt9mWK7rJ8GDTC5eaYlMEXJkHM
Vgyne2sbTplYLS/7614pQPNO53Lw82IF5wXOPl/guLTRgsiLH/gtJi4JuWIfR56S
5Lh6Iv64KgQs24W7Wzs55lUbQHZb1yqIneg+VCppKtVAAVlSMptTuJk4zWRyUP+Z
kfpR3rhSJXCL4/G/GPIfyYhWDB+fP6FPGBzq1pAcTXoXQet7okDtj6k3msYzG5Lb
LZVz1z80h+gi9VjqTQ1sv6HP+zZIUAfbds5aEJNxasBgs/uTDIod8BGNVwq8My8N
xX7n8W6c6TsZS9Rz/TQjH4PPXDcNSVtkb6jb/K+aW2ges62HqR91EipEbtUAFvE7
pc20P3fu3bvbUQ6whCWRZKj9SaP3csqHbWdolzXo37CijpC9LKD/jHtTpDYc3r6U
29rvRyPO67Cf6gCK/BFcjJB1gbulKTPFT00+Vbl3Trp+ukEMrh4Y4w92zU94jQDY
8uACzN+9EOAc2KRjv5u+u2HKBLPIYB0emh96l4+HUSQa1HI9YL6ovBlbdWtcPo7h
hRayYcMJyUJxUrj8c45/FtCM6hteZY6sHHAn0AALSnJvxdUdgzK+sh4vLKxn6iOh
n7PGRydYqHQa3z1RT8JwOTCU3nWgpTqSUN1+5UlWJOT1xirDDrvNLil+KGp5HVcm
RM8s5QrpiXuaE721n4U5lrueE85iS09ZEKOUF8G/UPuQcAemBLOsBnxH3JZ4bHtc
FTFRWJBrdfk6e55aFtWAQTi/5LolSvxcIcLElvI9VGH0Psmh7SRURh+nYUr87cYj
pnoKu3bAp8049p4sfIrfwYo+Q6agDbs6P7KQOfzvYUsc1jybSBLkHJJM2knqk8TV
+U3kGnpItSDdDvORtZ99VL2mre9H6MATF77tlOWBtI4E7qXPVf2rOnvIu1ET6q6d
MdaBmieEuaNKC4M8q+X6Wgo77AT+5ccxxKcWA3RcPxfH4/wKWxXZMKx7LS6xHoOK
oCqkMIsFEAvEwS96Ak9krpZiu3fBI3piDMbMfcaretp1XPM3kUWxe5bPdPChd9+H
wP58sPineSVo+iMhUFAL+embW1talKtz18WgrZBj5cqXaypRECRRxGYfcd9lq7O8
sQTijkOsOPw03StU1oUiygahZT852qXT0a6FNWXiIrFA3fV6bCD8sMofew3AJn2E
gM65kuZnvDSrKjZVwA6OAGorWT76c635iE5v8YXUQwfaFra8lT8IeDHUqOp8y8lM
i1mGwkDnr4ilG2RwShOhqVNgf7gmNKRa9ec6s8P3NsnlIIl3VPDhQgWhr+J6x1oa
uF/lL7sGY+fbwx6iLDCATSaeJ3yFAPK9bOC7/iEM2Dn1Ai56VmI0oHBWw1nP97SU
TPc9ztjIkHUNRksANLVlL645IKJqb2+l6xhfk+Ed5M6JDpMY194VbhO9Iaj1tUjl
osSQT3Yn2nngJNnY+QF3pWtslNk0ftfz9nvlFLJAPWMNZxeb5UvLvVDWcihPuSMw
k1JWSfuviiYD3C39YnzOZLdd1OzKvtqwSVnYOqP9FF+n7w93XKEx4TrcOYLc8/Mp
ItDaGDurnrOcQiWT/IxuNLrhHcMVBcnXjy31uiqgAzuZLxRbuWJVGwiaQIJd+47e
j795OxzlZOJ8KHTKJ400i+nMpfYhhz2jBn2aMRxGSg1hlamACKMi/dPMyZYaYlmG
eardW6t6BOTGwUZQi8Tz03VMnAgiaWfmFVJLVz0PIFODYQ9v5+sOUOraRunvwLW8
/j9MujP2Sfyh0MRf3b9ZFmRFOaFI095BGhq11U1a78ZiO+HKYn2hRMJXoFeux7tg
enD8Lw0UhUkwfqVVP8fQHquk9bppkJ5QTAoaWf1JryqLZyURJMel4U71CE4sF1f4
wjV26xPQCxZBsgf+C99Mcav4fAGJLRkY24i78/4t7qDqxCvE0xMPf0kcZsJ78CFQ
aB3Nxb5PkWzTNUm0d7ieV3QqCrU91Z6jTYNdl6oNUxxFxIvPDyhigXsGQ6v2gKSG
Qhdv35ULDA4XhavSmZ/r9t8ryUOauHR5Gnopftj2Aa8uU3100VoWrd8it7MeL1v5
IQuI4cdpkk9dwMS7LY7yVeg/XIZ5mt0QKH2cncZ+kIBFTpmhzUEDJL+/nCtH2NTK
h1M3lY87N8BB/eVs308J1GgJcGR2VINdldZKJT5Zx3D7cYMusc71jq6CkzTNNYwm
yowrNp0dbv+x8aS9NnUVI2SS85O0o0I8suPJqtJh6OfYMphdyN5huT55cGt56ZDn
auOSL8xGZY1WmGurtzqUMeAEXuAb2EAulyEiyhze+IUywQ+hfnw7wQRvPaPsxXxQ
gJt4P57+AZeYKxycKLd3ynZLmLzOe5GH4i5vsLgeRFYculXd+jgFHuCVywU8R0mf
WE2lIPrb4KA5pjloZVtb8Oy77PTGV/Suo4MRPcB2w7wh9r+6XnQLzM1jhDRbttbd
bDpcoGlCvNNRSgOV2FpiVmF4A2BeDSTqmAiYtnl1otsB1CDZD29umL+O0MgRmQx7
9vF6B+TjJpnmk++/CCvlFulzQ489VohD/ZXEEhjwQMyTkfgvBIZRRPzbMxBLHnOB
ZSsGJiAkpnEo+otYiR7NzJBQwKHbbBLcvQpDRyLx1+9CLIxE1RWfJwFEjg9Bb74u
R/uvDb3qNQcbOKMHtYDMRKLquDqsof618xe3K2JZsUxcm+b04mFmA6z7BcxM+JXq
asDF/jVVcgjzsRoFldnsHSsb+squ9Du+qpkbH+wyfzKOb1Qz4/x4C9xPQHvH8oj4
SPlpL1R82ZTD1D9HUN+FGz5XHoZS8Sf5KBjuy46nM72Q4xqNpkaFUsdvICPoblaR
9eSMZhdkZBkVoecIeMbWT4KlerhtYVjKJDrzyxvjECm822QHIM84NMd1nf4+vS7d
I80veJD84OXG3QqgOXXl4rEkafHjFZXReeFERIQuekjbcWu0q92CeQokoVXx/EXz
/ZbwmaSgXMeEDo4F0bPxKlE3AROC2Z3h+Xv4tCSaNvcOsAgX1/ZKJzaBjS9vo/jH
P9mxVpEpeSksOMIEJPaZAvqBR07auP5FMdrtLPeX48bdoYLm+X0MM1hJedpYdl3/
2HvHcghjWXO3jdjU854P41ibPmsABEEPgfuvgwDwcxHXE9DZZMyMIL370WN5F7sf
ve99bzw4cgh1+vzxGc1LczD024x272JVziXjq1NFKfD2/O17+rQeP4O1zsAuCQuk
197CEGAP72BNq2QGCe8NgBtkQlSswzWXfJoECYZ8Y0JBmdIxD1A5PcrgINyBNYDV
c6ifrcTS04xxBYw5Kc+HktpfgRLnL/uX5qvg2fOO+1Vd0EZcbSyGyft2GxHCBQo2
uwKPB9teUvuqUtAvtpAtozuvvdqX0rFiR3r8IZ46y6N+GhWg0Geql4Sqohph5ALT
EiYkb4tMgFQNW3NnqBoijarqWPCmSxpGqc04hkqOlkMIQwB5OECOHulGa0sliYGr
ioBjqjrR06P0KIzC3lRyW/l4p0FofFnCj80uLG30qwq8tEJqtNWIT2108S2B8TsR
7+VtPsaSZR17G55eUidzfm1JMF+kFldXlxiEAu4WdSrovQBuvrSJcTcuQ/TMJ2Ke
sZty9EJexVfMXSuWuKjEq5x7Y+HmlWnDHo9Dp0BZ0wb1Y7FzdFgwZKTRXKOymZW5
ZxeM26wCQtNwbPkupKWzJiLuZOTjpqv7hICObM10I8PdWX1jJgryWbl7RGmJw4ji
+aYOSI/c5Rf82X+N9J8gX7nc1pRuILNr9n0iNPykUNGag0A5fHCqI6+FrReUpFtK
OCDh+rm9ZFAFNLdNOnXBp+qVZGbx7z0/XcUmrlVTDtb0QWToMK/T8qJc7173oXrE
tuYxpwp1Iv8KJH8Z/zNdKuGNaxPFV+gau1icX2iQE0rVgct0SjKhJ8d51oI1uh7T
bhnp6KzNDmboijk+iIoNAixilfFhG+8ANeUTLHX3uYt8p1CqAMgf6hHdwb9zCkiK
IOQAoQOcFpJSpKBhrjegsqQBLAvkggJEsBbLiTX1acXWDLXHm73tTDeUXrXp5C6c
pRNngaCxmGFZN4Y4pGOsP3ouPkTjbMD1F/IZN7GnoUerhAGQCK65h8awn3RVjDO3
m2mlFgBBIVNwiAGbNnqNSrI3bHOXqGsJa6RpmYrZaPPJcWsd+VUVGN0X4O8IC7Nv
WtBqYpz4H0BhBOQMvtX6OQ0YVUN10j3dE3H5sv6kkYMaiW/YDrJ+8TdjLuVGcOGs
+sKMHdRhhluxborwsR3NYwFHjvMEhfknkE8V4AhHtvjoTf+W/Tv/oPpSudXbV9ET
BLjrypQclUYYh5c1YcqF3MeUbKdg4cQYnFGgAnSRm4zGa2nnl0k693ZL8tDuFyfq
9O5Rvt5F4PxU69uZpZ3+5761uwD7fkIKua1C2xHu6UENcRWyvCcIjwlehaF1JMRZ
1U+cxqr/Q874uUlH5f32GXr6VnYAuPLBCXYmIRs0KMeVVo5E+/ZxQETMLJD82dDe
+HIwRcOu5lgcMwvaOSPA8voDXTPYv8NwJRKx1sfZU5rVK864Z9RuZmRUVD2OMp5m
hihDpmymiPuTOTDls3ar49GOW76jCtMxZn0GtBTKwDVsvuoGiBbdDk4+WBjVTiaQ
q3d81nvPhHx+M/c9HeiJ+SlQYh6b73SAQYUG4UiY+BEkQr5ePbRkkZA36JHGil3Y
OBmll0xmB/4jAlBw1lsbAddIYReRUoOhxtUNms59/0AklULOAjc+tFWPPTrZOOPm
wx+7O2qG5uWv0ilaNgMdZbKbZv1J1zW6Z43TBJSpS9JsNRfpIK1SCBBOa3Lx3XZG
tdRkrLHrVT7pj5NTXpbasqmI2LkF4VtUR5Hm6dDPvWvhdVA8Umy0+z926ML547Un
tJIS0UShePbkHkSwOLZ2n6VoGqxD0IY8+UHPyS6Vn81wtT67l+mzZEC3KdwWMKox
2sK8RSREkEPDboLm2c1T6rCSWUPQwAn81P4A8GnhRzSpuHTvziaCn8GtkyQ16ZgR
Ni8QQLqSVRAPc1kBaMoSpe5jEiFla1sosP+Gn5qebCGn5+BvVX/IDhGRK3lSJ/sz
MgwO4teK59YYNiqxKhldHrGr7zas4QpjuNo4ckTntr6NuW2e273rDcj5fzkY0t/1
GGzanGJDInPXJgsduk1yw6tvXkRScUhEDm007dElbmt41OOawQO2zKMQ/86inACU
KLq9dijZhXrS8084DMJTSTnZd6FAmsAxqRp49g6Fn0A35PaT79U49/cr5lVI399A
Um7p2YI1Jd5vuhWSJoD2TfSRe3JaHt/V6QUlO2dKqbt9TKWl+kHqYaFNFYgJdobK
N0bXkrJCxVHexhXpmsQH2zPWXVRmYayV+mJK5Ez3+WBg/KVPtENhpjwrzubyRqQ5
oAs4sDyGz4OP83Ud/Dc9vYjxZlYM11ec1+nApW/CSHzrEJ90xbTbIomN3yQ4fQEI
8GAoAoOloFwb6y9mQYBu2xXfY/a3gh4YCbYJm7E2YHcrges5RJvr5ehTqDEEgIZd
rCamfuJYBTZnRk46ytthDZ9103xdYqQ+turkapC1XntXL3hiV8JiiR3TEfCu5+44
PLzm9lDkJXgwmgWy+EobJnJRJFmuFoiJ4SLYAi1pX+eFvvzfKuxuQNSD980do7kR
d0MIU/Ehrho1bAg6Th1seVNyn/TLv3eJeDpzqLqtNPPbNm+T2D1pWYE4LUItPGVn
phszSZ8iC82GA/odPZ56j+VO77o7R7PR7oxsfKPVV9QTiGQe9M6vMTS421ctht0+
cMT6MaML7FM5jyh3hlDN7h1nOZtqPKV6R38rEXBxefCdel1JBigcExxSVgUZsQ51
OFokB1CQVXaZ0uyOxXQhLMaKwG+nRrgyo7KIIffYrQqEuYk9bGSjINW2zPGoYlf0
doYRdcxqwNSTLcVyZPFEaQInVNOkQD4lZNjCnXy211YeVEAt/0eGK2xNWivm+Tqz
30a34rL+opmHBo1XlFMae3Q/JnDY7jJNC+cWXYa98q3BpUiJZwsyqJW8GEre/3k1
6qnqmmJUSR7BegEu4Fblp/5bJWPypTmUy1yLNYq6oqZ6muC4zR4QWQSH9DkYU4Jl
UlEijLLgQPzTnGZbzrxjDiOyGouA7aLPOr41PT6cac55LoX3GjRINmwKm61prgrs
IECoIaghNu23GCn/ECaZ4RSDFla9pGzEMsLbRza9WGjAltOcehYL98QA5JjGGiTs
eZ5yY9muXLGNgNIShpywHWgkRSy6k+qctpy63j6+oZApOmM69cdsAaXDL+7/qpoI
qdppQ+rkpOTXT7yRT4eyQluMo5MRVnxA6oUulwUAO/ZcK3+yNGa4ptlQPElb+w55
TlvSiOMsSxtUfBWCxQK+NK8VnqqhKepqFhBQROeuEwq3dHiiFB76PUwdCTBWnZPW
g0G1lKljE+0Q2QcQdjIeT9m8Md6VsjrZr4p+WQc+B74gmtpvzFx16ZxCT3Y8K5Ru
VcZaiR+wAWmrZ3p3l/i2M6fWEwy2NuRXpoPhSH/8AQxWvvu4njKURsjbEhZXxYP2
piTAg80W6LBlDOAk0i1Ie5RgHIBsK1uanRLB7/+E4aB1qd7T2BoFSdqYXcuAoGHE
D56vDeFBg3XqDOLv4e8V9gVBCTgs2B592zIBFgA6/zZrmEKF2tn9xxcBIHyNDqhx
gI3syAhLNSyEsWPWa62b3DGxrESyyeTS3WyAgL1OVpWsCSSC5PpLBInWrj3PNsfg
72BkjuzPAEia9TXMIlPvN0o3oXyimf1isUw3iCRCP3S2r1hKkG17JnMZOlncmk7q
6RGfpF35ZUkU3lJ1KHx+zjygPnTMDIcge2TYGWFjdqlMhYMWKM1p8lWdcVdjbQmU
bKC3540BmuX7mN81lf7ncXOlDcDwWYRqR9Fa27dvXthwfvV3JrFvx697T8YCFuOM
y2rwTwAChIcDPwkA2P4M7uN2tNWoPhqe+JFsoC1//rBNevGejxKQQA/BcD3ByL9/
bY7yiY1xnIDCjU3AhAuNB1+X+DSyMeFamX+jLL/mm81VA5dCaZoW7ck+jyVPzGBB
yIolbdh0t3yFwZaZBIDtT7ugriPIQOvVkgD1Funws2Axec2zoXAJZs17tR7Ovm5w
vSjNqrb+jJKO3Wuwah2OcuNcR5YOWS1Ce30G6cjlDW14TVn3N4PIA9divj22sRq/
HTEmlQXJ2j8ggLHiW58fwXqjihIISUPM+MAJxC5Ushzp1F515+iNOkmW+jyoEeRV
M8T0AAFyUIBr5aKw0wwdzGoYrvTyPPcCEqIRikQB7gvS1dDwtxCT96Bhkrmhgrz1
uHL8ycREgh11D6T37iSZN6UlFLHUJDYBx5M1vTYF0Q6tLW8GL+t1Yk3E2s9WVebZ
cQCh/qdgrzTQvnCSiokWnwk5ItToI3hsvz26kM9e1RKpoKfwTDcXtBSKM7pCZIrT
zl3eu3NeHLh0FMdhckO3ecEILmDC/LXNnJSOJdUE4vsSUShp3OHxeNe0ls54RyZ6
3j3v0j9M3GZsaRzgDcSU9Q9ZjfygG6SF1bG8IJQVYrPpdDmETuNR5FUkVkTWTNDN
x0PInE1LqFqf2Mx8MRfMDkwgLsR9LNT+ySzineiRkIw+TeyQgZ3Ad7ewRAxVFi0b
En+0tYnIDpuarKPaNVSgfLC2imdBajHVEf9UGqvoFV0VOok5Mk/KjwxLzvpLK/S/
ylaohBkBr81+PDMY88SIzYIiv6orN7t2Vd81VFlbqDUf8pk7C7riFeF3noIJISlY
oDcvz7hPTpkTYV1N5EV8+uN2Vgv/jFbo1yS5djtTnv0A4fCUUm7PdkTTdwHWg3E3
yZsCpDVTwYqYaj5oeztA3KYKroAIf2SqhhSs+/vTj1Jmz6Pu5vqdr2562kpi8Fuz
mQHSYdp1uE3oRplTOyXTAcai5x9TirrTr652GNhJFreck4cPIaGAyJDmJ3EyNnG+
7/XdhpaZIPyv0Jgnn4pUJS5gAg5WKTKEw9LC8G7BULfQ5yv1E9j/kzaWPBi84BK1
9iI7/7R4uLND0dG78EIYDSdapu2mh5Qj+UhBiPxdfpKBr5UNXsQUXr8hszpX+W6y
29XDnkt7wkTp815V9tHShaAUOVmc2i8uFFJLhOS8qvXaNFcS7mCy6549NAxV/9QR
43Asm3AzkH1kPuKw+imAzVdGjBcqhMgVeUm5lkOPE+JnGmteiu8CSF3y1v/78U7V
HMcgk3aCazfOkVP1nKO1YAesTl5jxxekGBjHVql3K/y1GYTWnCOvHI9urhvH4wKK
YyqMOpkE6r6QHmVuxl9+Xcyahv2ZAyh4N6bYgzW9cFdi5jqSaqZKmWUxHRMvTFqp
ykNai11HNQtTxEre8StZ7ZGb3gn8qnfxtCKfdm3GDzDp+V4Rwf67W/NGKeqkCaAj
yALnlaP87wYH6lYwVDSeJHivpvN0AKUD+15dESACT7a05PTkfViW2W9UiLyX9JPU
Uw0Faf4F1MGpTRtdtDiH5OVU90Ca5xxf+Ha7EaaJK4UpfY2UlFIUGeZqUjDUpsFc
LQ4QR/CxB8/5tQHCdLWtOD8swpI3REQ+4ZUjmsnu8ke24LUfVfE5kCXrl2wNP69Q
jRx7xjubMeuT+v5W+GVSJv/jTaTJKgxZBBANASZHu2TEzrVjO2HEjrHYKgZYRgE0
tgWgHIuJKlecI17iPsNR+joWW92LtzLvUmJ50mhbt5kG/riAtfB5uYUF7LusyrB4
dJq5zYuiqKLY8Gh1TSeD7E2efcBqSdKdeyafs8wgkZDLdpwHQwAO1XE7duf+ovPZ
yZXqbuKGfhAm0WENj1awv5rgbrpFVHKQBhXSdxEu/vtdfDG6BE5yXkyMtTf0c8Jx
IPmBNiwF9qn90WbUS7EL96NeZ8/S/72J4HhWJjgOqsYSelTRmj74p3RH13pPzLhR
ApkU7O5+Gr8wTChtuGCRqkF0H0gQdUzjvQ5AV3VygpHuYlVDXHVKOvQixuuuU8V3
D3Q51FXquQhsAhtiAIV52Hdm/KZ9cGlqrF8cOJ5h6nT/mLc2Dpbece52EIwr5/KQ
jjXyVNCt4L3TAnRM4Jb+0kFrFjTWgKxI4/cqgo3Q3f3PlbKAlrPUJpbSXNgFli0X
DIIWr3dmNw9jekPlFuRsCh3Ytj7nry3eClyUDGOjWEG0ppcep8MdJRz9dUGykT8v
F0SWT8eczaubF+12Q8PvgIZh9+VjSeajN5RlUc+O6LkYrz4Yx5n8cmoLTCih3llx
D9eXku9Onha1hCHrLOQqCW80KLNFDoxwXu3I7zr2T4xSWKd83+Wy11pMeC5eY/NY
uDvqyqD4jy3En/BwUmCvxssp0CYwpl/ClTfdsBwZKsRMdCT6chg1GHnsEc1nH2WU
5KTvrdmpNJ5+l5qwiyipkgYHFaKgfANb0beHRW54BIZRr913iA1c2a89FvSGolkq
IpQhFI6WBf42RcvkR38gHdHSdaU9aNnCZlvjjAe9HQsNJbbRoMXyUvSIns5Z5Toc
vV4bKa7RPK5QNM/VW8lPHAxaIcUtTTwP1cWveEF7AqAi4CvsY+qdSJpiHHfuPsIa
q7TyI9oK6VYw1kKmUgZUp9xxA+uGbatOLe+i1XE9q2OVlPFRPYJ55J6gXEcT85y6
AmnlMc1CpdvORraGZfXWA0xTV7oZxZYtrIPGlAvBjoNO/oBo7TxKds/m2GPe9P5/
a1E/KWpYxgka0xn1bJvb3pJqAFX2RqK5VA0FA+FdvCoPrQwPOLbmFWbJrsQpxskx
HFeHCVahCmbELiawxzh7EREetHdm8Ks2TKRSZLfN1k/HUmdVPqIilh8B+Zkf+ksx
39cDdSJYYk5Ay55OtY0ee6ezqFEKddEYJgALHPzt7xbAfJ/hBAbhNoajJKgMBVh2
BiXifybxOu5npWKK4l0bwY0he1Zab7tsUD3wdIy6HaHyrwEUixl7EAZ8qvRC9CWD
uOuZAammwqHhX1ZnShEEsG7u3H+P1zommQgOK/hnKQQUz5WH2zZynO7ENwBTGOgg
OOoXLKtcxcV9Y6WtBDAh746MX3f5gz3Ho5PqZWgFg3SWvIGkXgtnhM6s49dbEZir
i8LupTysczscqVGwy7WigxDFmR5d0DTf4TmdgkTV7OftBWho7payzwseXxiExd1u
DMtLBBgfyQhghW9rm+AUOApXtxKEullV4c3V3zGNMpHx0cHho7zxP1tmMtVngDTy
BnC/wV03qsjPiEPFark3VXUwi9EWTHnQ/UtTIwujrEduy4EQwMcH1bEX9gOfcDhY
uL9IeHh6vhxv9kWNOjGS/GQWkBjXtqoWtQpc/6wUJTwAqGw/JpXYG+obxmxLHWhl
5kUN/ZR9k1H4jxt6MTAC/xJKi89h1rfg3zHN6vrWv5+MwKW/G79ra/CftYtbBnSF
6xpKrbYG79KjG9/teEnm2kV0pizOM+NmRlx+z89RYXiWJbsgWnNJzXbOevc7k6Hg
UuRNPXXUfdzIKX2GJk2BbpemCVyOt6xXHXhjkojocUWycj3rNAJFmstbU1LRg1fJ
J8BNejzr3H09MknG8RHoRq06vgIX6Hh2NJchfaIwGu6NvMkfra1oqN8l0lB4UlLw
Jo6Nv3CoUN4jfjVG6yRcGjbg1cqN/snkPr9G0ezVjTG87CPIvXZOwhVnc3ipG5zp
guKu70F17XowKdMLh3bBR81/BFMC6RBFly56y2fexFnE/RiEIcbBdPXSkkiGP07B
AhlEB7Lg1mFW75BR1tgUMxyI+dlvc8GlqGdX/WJ8F/6buhkycUhD0VgJ6E6kmnah
3g+N7cXcfkfLeutZg4xicR3n37wkukTAJykMSLZfE1b0O5PRt4VwSGiUONpHH28E
qu9cA1y8FL+09jzMp0HQXEAjQc3XuYuAe7wR+I7J8hsMg6ApgzHQcE4h0+LqfkoY
pezGIN0Tm/V/7MDvDkFrrQ/wjId1LcXhQdCqp+SjXSDNesx+0t1vLGrgC4T7s/9l
tmkU7VT76RMactG6P8GF0CP6T6/L1TCutApQL9Vwc2U/DyC6D7iY2qpRFoKdv7Ol
RV9oP5TdyXB5+VyLsHCcTUypd07l050U8ghK7hg7Ltp7cXpO2g3hVchoHzQ2PV/5
ushlg9hJwvz6pFe3PCCKQ+1Yc2HhiVA5lSuc+GC+0uwkUtmhiidTIFVv8nH/pbfy
GpZbuSAVKiyjhzNk6CUaHkESIDeWQXny8xFl8uuP9r9Swq5fdk99s8KPoa3Z5oyl
Uvi4mwkwrDtY4VfPrzoDfq+QSu21tgGv3djwFeSGfj58/2LihnuN9IXJbo6118zq
BGifSx/VF17ve1IguugB6yUUJXB5STy1e10y47WjNjU0zdCg4e3Q2HCmwwPDxIwi
iCcXl/g+jSpC5ezqq3SAXI6JTzXNE000x5KWaDHHhkZL5f+kMcoGmJABhteg4h07
yFQZmKY5DkqmbBZv+IDljb5ksL8uLgOq1hmjCUBM9fwEUsjvNYLUpOsW29sCaMrU
sgYjsszVuLKu+/HYUAdF4d8mEgocfa0GgHLwamvFs0a5ey9FCmb/HxUaZ1uHM22d
J+sE3bHv68U5TN4zom1S7jK8JtzTTWnM2nUh0kWxGUq5I6LPiiMFL5yeWE/j/94I
RhHyaad9VmpjF+asRY+mLw9fqM5Dr1HtvqP313hZf7Agc+g8G90bXJHki0qQpOrm
XY9V4/AJ469yIIoCfhewLe3HLa/gOe6Q97NOBu91RlY+xtjNjfKmqIEgi55VyBQk
F6e1LtWWikfw0GFkNoTu3iwhzu2bBp6tfYRJ9er82oWrVaQJwdtCVfVSlmMzuxA/
ReqxzA5U3rBN41DJsZsMj4cHQsPhXHg6/su0wV4kP0WatNOYWX4eWAn1UQMPPTA7
NisQ8/0LOvMV7Aaaw7gObe4sJaFm9dZ4xRPfjXT3woIrrVxgsmXaZrNwrO5Q5qRH
4T4FTMeQxqSXWLNlftRI6ZS0C66zu1iRSFvlSGv/ppSCUlmyw8hxGoyV7UkVrw2o
5h3YGRSv0Zdq9hKQFDfyqIypraN2EX4cxhTOHQYloAwCi+65Yy44yxU84qUt5VIr
e5fX50B9ad4zcAfN9Zz7oS5m9Z0+NN7cOklVnGLIgHOCnDvCqlus8yvtEZemkDNU
PfEj6IMa2CT2pt754sFVAU5WWLJI50ymaIEPVgA2pxWSj6xqkl6HQq5VanDGic2A
FwZQqXibnbYB7XLr4f67qtUEU/yAmo3SEWCseAyQt7qJhW0q1ZYy48lUZy5I4qkL
1uBU4yUBpym0IR9qTRVyD/+gHtOmFzEi0FTfbIO2yu1tG0GKhHCUvWNrfkTvIUh/
+8isO+m/wF7qKEveGMe9cfGVVXtlSgPmg4xVa9PhOZFkBgL/uiGCia33LGq3Jt7L
K8RCFDp6dj7I6Bb2xGkMiX2eJbonBZ2yYJYjDvlaTsFgQPk2PSFqUwnCYK6XRxlU
XRXsUvM4LYq8C2lCvaQ9wMHPeXVTg1Y6befCEtc9jVKdQtjL+T3RHHrNOCINJuYN
Mx5zUI3S39qyOoIuSkDkiE/lbZp5wUh1pkwFEdEaV5wFMXb9RsoLW7mhAXEKHyA+
EFH7GofVXUQ1KonBmQvAU9I78aMuZWFro07kW0qE3kJkJ/R0pz1pcsI45D04Tloo
FAug99hpGeM4UTaYfBlXjJr2JbQWrs8jLfUgAmhYhZLtlsWiovsFB43RugZx7+4t
9clWGakSMQahwSpQ6amdOhrcHujPY8NGWMDsJdO5TJuqD4jloMKE+Cvo5UgRJdrg
0uJijO4HAN2A/NWbyiIi0DZrmHm6pW15pKZuVqJxEMuMC/H89ry3qyD0n8qWBP0w
+81MC2YP0+1fmPxLRTsczXqFZJMgUE99wo/5f8bkbfzIZ+1mgbIo7AqjKUBNXGvk
EYLmmdCVHV/WY66D2nT1D8yWH7H+lZ6jgf4zZh0hAIZRmdHXtyGY5hE6mreMf4i/
H5asHMbcw0Fg2JP/3r0TUuOxYrNG/cPBT83U4+wAjmt8UPjh3EfARCDqhGBr8/Iq
DqIM7VDGGNBxgPRqZ4WfFuE44SgP6c/AfO1fXJZsLFqr+2ZuWC4E6A+azcJd76xs
MeXm6Ytnp+9MSYwoHeAUE42FfaonFplAJBwGy6pPgBNpUjJ53w1oX829qJOg3OGB
+4ZvE/l5lEDmDMmanCSt/oVCKZZ4CBWbvA/5vtaXxMUhRgF6zi/euZadpn6iB2P1
262u4ic05vONmqK8JsWsw9ufDkgWAVP8SP6MekvdU0HbalJ3a0HqVENkpvTxZ9wp
2yFwrqTHI1ilP3CRzE6eVh8ptAFktf9/fuMJ3ncXe6oRadBTKMey2pbNbns9BJR+
h0ufLmqaVy01zVz5oWyzIWVtAITRxvUFHEzFwMIkX8HrmjT5Wd3hg5M4xTsB+YZ0
EvPGBrncgcDPFoxmdyDSrlGAS4sjAlvEuELRXOZ4ow2lvCey/gsS1i7PpV2q/gQf
JRFmf3L1nC/H25DqKUXy906D9kFB7KauBdLMp7PDaa3kuC+W/HAAQYiG/wL08NGL
xqWyUgyUYx/lSDsrQ/kkcHC6e29XNStLCCyxON+/fJ3kFf16s8ylBd01dSySluHP
4R+m19wOCnDlBIqt/DePP1YqZVNBYQ7LfoIRTodUXZ3d4Rpj7i5x5iV898eGqE1U
MAQKBoRirHnRnlnijFiPIuPWnnMqEX2HqnFGEDNgRzwVCZn3d2NsMjdfnTEbmDjY
jG6793pk2gPpArsnkOTe19tG9k0G8Lt6YI1zznBiZPgs+jeTt82qE8V6u9P11o2U
EQC8n02nPhMlpveIPCF2Nxmmo4ZTmmxbqpduIZ++vna6uVOdPNsVWXT4FpIiYR2K
6zd/ArsFvI05QCdEL3DmRtpENnh5YLoYE3BoRBGXpHtKI+n5OJVcfgsBOTWsMfob
b8AA5kwqnbTra6YTlV0yZhwCbLnI9NDOrdW8OGYWz5Ojd6pC32RxbIoyLsjr2HvU
Qxs+72QaiMT8ZoA9REia/rolE6CCnNpfcHByj7gDWf2rQ/LGZ6p8WKwcZgU+eilG
dlL/+IEJyxyjZpWbG2eJXJ1ZlZT6b2hzIXT45VzRn1xo6OX3tH7+GdeJktXqHG/i
bFJ7NQ4qe9P6DjpOiHbM1c0cHP80p2v9OruqQaLvucxCEyjvnG/pINGd/IRhD7fI
E0FXnwa9wamw9sV/Vs3Wr09agPnbsLiWFshLjT0Z+lgM5COT7suBh8tJgwTzsb8P
pZPcZ3uOWvaLA37MaPM7qX17MHY0WRsDMXjmWfMfj1gcg/g4rMVg8u5xsd0GJG7k
C7Bmd/aYr/AKUhjK6BGftTphzF9jMuWHRAV6QI8MEKlwDDyjPlXkgAzI05ZXQBCE
+C5DMfszzsrpmUBA/RcP47pdF836qZdhOuPn6MVjb1vMzeBIYyNyCEAaFumzmZC/
4s5JR5QJYTkAjcOM6t6IpLSs2/OImUjbZKfOFv+ISFsPpWqBUERuHjZCAAhRGloo
GeFoV04G5996vzjg511CZ7qfqXJm6OLzXOfRsdjfRPcVRRwsioLl7b7CVJ3cqlzo
4r6avZWZfZpqLTT0olw3uNFK+37cD6NtEiD8ev0yKMmwUz4jvRiz80irjOEU+apu
14xEySpLStLwy1nRSePOr665AQmovNh3E1vVlry3pdoG6lKl8+GGzuf63q3kX1kR
jYXdjMpAsWMBtMrEBNVhZ5RNfurw/xgBDsH+O9OOerRkLoNfRf5qf9C2pknN5C96
K5K8dCy8ltPD5Nn+TjVYxOz51BmNw2Bc1gdnv/kk1JwGqyraEjBY+RwuAW/QXiR2
siG6fVxxmhLPeDvhum9+lu82qzTiWYRh7olGvlboCQP7iElc8+yKKtXNlSb95syt
co4eKwWvLK/79Q/tJXENNIbrL67vY0fXpdobbsN3Z2EysbQBK/DwxyizWy1c7IUG
u3j3k8QyWuNGKy7CDarQhgrn/spH+MaaS5UTbQ7JOkqM4WNsFAtIUWuff2nYGqAQ
1RUa9xVLs11Vcp4dvjV7dINtpinyEXWO7Wdb7LWDgBnQVNQ1ezq8wecOvo18/Zah
AUVZKzbDVq5WBNFpJosctWo20gQcf8gFTJ+DUpdRoP4gLKU7CQw8SpWIyAc9bDM1
jUVr3mlMqZAPlvqZNgM2mLQzIPdwfOous+fkNLVZljdGMtxpqPhKZ8QDdFd1jqr1
31PGW0h+izB+JZ7fwQMucJon7WCXqE7ItsQcJtGgftnWS8SeRMqaosH1DHmTbNrq
BgXKnH1VQP3+xIOXKVkzdXyYKweVptAWPPjv5izjX8z9iSovVW8W3UuP3+Ceu5hS
QQfqBCf1qNxj3F9dmp9GVEO9BvM23iE66PGHT9l6FPrWnrsfUHVMVw4y/YPYW9Wb
XNTAd3KFw6VuGLoWdhnfTaHB6HRZ86HxbudIk/3peyJ5JZMnFQrjUJhcYsl3W7GC
8FIJZdTOQJujILcHxXItbIPxNqCEJtlw6WxKglMPYkMZWqgO5fxh+aXB125QuvO1
LiVkiI6BnmfO6barD3Oth4a8L13vxJM8/s8lIszbB2vjbCg1hbFvd8oOeP32OzhF
KHsq1RGCv8CNLGNgmH52vLfU99SjiBSEFfoqV6FU46inmlSJHrNkJLKBGfdprTrS
2jspPwhSzkf4uzy+tORAaQYIfcAO0469lcoKUxkC9l2Rf7ADWSEoReWaSoWnwqxb
AdVSNb5JJiDSGWfjObH5iNT6TpPivh+Euhacx9Bs/Gx1kTLtYA7c9wkIjkBMZDVL
xD+aRZoX+v0ZL3RNlBd+0MQ5fJRs5Wxq6EUeXdiA9/Xp7fAGWkxRoGiMU/83+4YF
KQrh1XVRw9JnjGGengNxpzX690vKZRSzB0BQfI3iAN/sSBwpLkh1bjJv+QYY1kTd
UqFcEVPlFEa5VXMUE+7zv8cP/N0OHMh/mbRFR0qtOMr5Rm9v3ixgm1IDesLT/r8O
AMer0g776inYTxZ+w+jwXnwLxnlUcprpyaBDONBjeRE1n3xylnQY9rqlLYkuJhIX
/1FDDZz5e16j+533zjQtlAAGLJcobYDxWY8rm7tAKJNRy27wpObIhdTPCMHIIIBe
cAYuM9Py8OxeD/aYkO7FeLLzkS0SJv1/3pu2/Xh1GXvKCbA5x9Q+FVFn/db5sZeL
JChXnl+I1CLGznuc3zBd9NkCsLHsC/vy1whFWsVDWaCs0jXZZDdZKxPcKAzo4mpE
8C1+2nF8qx1/8PnP1alkt66bp/bunfWmX27bFC52pJzx1vqjLysEK/Kkm0fgGbfm
9PcnOKYuKwixIWdcTmcrLx5kpZBY1CZjd9YyHHd0PMgrfUQjzmm7WrpBwiIfu5ci
dVB7aZlUDJQD/lDwY0AE1ph65cjw5ZCKDNdPkc7iuj+vuSINTGFgqqp5w2JLkA8j
EY1E9vzMT5HTQQHeBBq49xJgIj6p16DAUQnSRRL0abBQrN8R8l+ZROx0y6BSYIWG
Gbll7N4pgr0zzwOMZxLkcdJwjbhwycaCcGl1qHN+aK+52/nrEM/fXa+HsmIIBIp/
6iTDeG4qb/Z4O+FRDz2BJrY88vP8zP1KAuMi0rhPLDhDK93HtyLYXRyU6OnKUos0
vq4F6ZHkR28KOjS7WeAlC9iVj1RJ5myWeEL541+OatuW68HKYR4LhJ/dLn2B2v/E
0tSXa5pPsyOUJzpRpiBnbu2ZvGNj6/9exnlvZswacxmaVkSXSeg0ka9SSh50o9fQ
Z74KNbQ8/K37YXQNNGXoCPmW6V5LXBAA7njjwOmspdyDfR1SosKwrheksBFMu1D6
wzyVv5nysm+XHLaEeeLPIV2q6o/dGrerK0W7htUeRR9fD+Ah62GO8q2bl8ahHgUm
2LNOGPHOuc4sVTLzVK3l5I6X94joBr5nCXQDKZ0jj+4HOsOEBWLoG95vrzyfghnn
YiZPjAtqDAfyVift/XOFyb3YCJP2SxkMQoCiz3Xw9JZoNAJMWwRzF0MCZxYD/1tC
fIMcKJFGlqwF9glHhoXp/MFMVCFBmu8WMe0kAehdEzUVOg+C5JlPXYXIOmKy0ssH
ypycV+NYURO/MeRFumMZyG/+eo5B5qqfH0KKqsHz7tDanhN8oVSIDfe0S2WB1D6r
imB+cNv500ew+0TClz9d97OAM8qMPe/gICF/gZ1c1ecAOYVBX25PaUtiiADmNl4m
tYjEs6eTgZNOOzU3ahIuo6sQa7WKOvhxjAPgeJiwyNL0KSxxWR1Ne3O80eoCqkht
kuxjlU2R7WZQyGY1+VZFYmoSwJSlYQ9R/70jqpvAq3pAl0dqrsIlXGH38Ic2iRxs
K+EQzWOs3hsEJAHijDgfoc9DjQgRIaAYb0tTkSHfThrw+TTGvdB6qcOpTvyQh9VC
TlH1Blr6wlaoUg4ZI8nqlYlSEA9evTn0Rwi8mKxQiDpV/GBeue1xu++19XupblO0
RDsscvXmfJlAYulnTB9KLrph/qhztB4M+jbHaCMIVDW1t1LQwwqm9H2PTyaEoblE
u3yC3iN1Woh9DtY+Sdlrxhy3xcr1RDobBMHfbmSSYF++QZ23G8q5VNyZO0bKQYvF
YlaoE2oHCpMpufOluvu0slDCuytH2w562e6pLGjJy1qp5/A/eSVlXRsI6bSYrPWp
dLm41Erg9OrCRiMMjVY7ByOaUmxlc0gq7GLhVYs0nhCEeFKHd1fBOwL9rfE96/Qc
tr1hfWjiuCyioVdR+zU1//WOeZQ3IEgdRjDlr7F9398OWyuxXe5A8vzvAJxN7btY
R4A4JqT24S8C18LxP+TbKmFNIio9MJwgZWegBsqN/KKF5aRHbCwi9XWlAVUuEz7o
XstiW/iny9U0km4B9uHbgVUTtMLxJdwVtPf6cuIWKSyQWwtE0jV17h8hiSYrECZw
gbTQv0wJHnqBzMIpotytWt47dntw6daT7u3qDRZfOsDzq7O0Jo303wzqIu7pOWAA
V0DgCj7x+Qqkubmqvj+3MSLykZNfrbQQCSl+HlHZMakLn6FPKhDGhG9QQ2Hdx4O7
5xIgvSjwh+3tjdaz6uYs0PXL1CM2dKy9laS+X5nddVSzTKK0s/SCYsQzvRiMau+N
/I1IaVnl8UBctz5z7iho5T+IOTZngNkUXwZt7VU8wYNvOSV/3YD93WWqZoVQ09oH
Cl2saRRBQYwfo41NzZA3wr+0NUPX4uFtSE6SDIeOEH3t81mTRqBFftvwxThHAOGb
h9kvGek+ITo9evMYMhymP1UmQbo6LQrYk+GyBcR1QhDLibBiNi+CSeFA7F2A2O8g
9fLA9V5pTaJLvzCpTurp6V8MLoKiLCNUhGz11h2tirLzO34+hZUZhwAyghA3TIil
8KF8/R1E3HOh0+h+3TPd8haQSkzgSeWIek5mxa2RWW1C/5/7r2ID0BkuIjTfTCoE
RAuymT/UVAkSjsTden+uqUaMzCPJaIrHB2Nz15QZ+TuBV8oE2khc9Y3aQVUEY9pj
aJryXvUizGjxJPEwUb988rnMePV581bMsT6XpePyZbHTfguxYgooSa6tQwDYtPAe
H7C247A3GfL4n9tVG7LHSmUeMKdn3jYZgyu3HMaQpU20s62bljoxwtHwCkPyeKQS
24uuEP2GrCe8ttJKjj/g2P9xMrEeI4X0Cod2TLNIf63r1CrMfP3HywsD1WZO8GjA
EBZ7ne+iglODENDSY8uCvkrodPb9Fxta5GaJc34UnR6mnf7rJhdgJLVV6SGsEjdd
Mf/XYHWQo+IPo4l7eDPNeSfOfg8S/wJSIIWpejEUac+OzWlKcIJF9VwcKzizsHUs
BtVjVpGuvYaZttDQvs5BiBJH8Cq68ngOFISAeuE3O3VFhBppEdlqMOFvdXDBIS+M
cDnDhWC7JUs0jgvVD+7bG6jsFop+z0asioM3uY9vYtxN/ShOwkXlFQltLHU4V8wB
teT5079tyq2eAaKLY2E4hWOGNXBecM5jSSZTO+cu94x1W2hfvOZTkSTawwvbBDfg
bwsjgAF8srhkY7eO8OdKXzqTnV6mUCkAiql6SwQ35AsXNc+430h5veUXkhTvpc8r
HjBvQl/ZcClHYUTwx+3z/C4NSi+aIHeYeVNjfoZiN8C2z851b4S3Dkrkfh52nMAl
CHZJGJ5wXaYnjC+LrRAk5LlAQKG/jDVVXkb+WEvmoQMWKPd6rSqF8UHRr4wIm+SH
M0Kakb3el2oPcEdvYYrezSa3zEpsJxtPs7SRiJMHIMZhgV1Mb3gzJSnNW6+eZNLV
Gid5Io2g+NpwS1ctVnfM/h2JxKK1OvnFVcX7QrC2BSWdfhKT+/7eujFJFn5CT/pp
vo3L81z3pWe8i+954kLPDaQ0Imdo0IsENF51Z4km9fV7FNLFyMt0AFiouZKC1vi1
S2aVqDLTy381eGYlGN0USVv5mvD1AGEyGSFVJdHfXS2eCFEDOAIQiYBn25wKs1tl
W1ALV09KeCKF2Ba5KQaHfHMuWoRjDkz7efIzqRuidJZjIy9s+MHFIcfz2K8Jx+v5
IYqdXkIheHCD3wWFSOcbbu+7KSnaHJghMlhbTM53Yp4a1SB0Z8UCAeZys0vWlPY5
YpyCVN6IV+KT3URiJZGdh5Kd0Y/12vlujg43OdZAu9ZOkhwnUqQnZR9cnqlC/R4k
VGiIpkMhfLco1SK7bj12owhzXnv2n4TlEsQEmsDP6zLWCmXh2O+lUwb4lIZZPzBL
0EpdW/q0ZBmnhqYgxNMhtwjJE6+u7u/jnsEowsAJb3uLfFbVq+iBpCnWUsWF72II
qZCN14T9RJDCBZq5fPYqrJcdhyaIOvaFSl2Ob4yO1EJsx06amm4LEi41WE6/aB6+
HPEER7p3oAfBJe26BPA/Y3b2JGrQtX9KI7YfRoX/GRG5KmxZpZTf6FLfuw/qvj2i
0CKAFAF4BvNnVqzKciNf6MVGv9flhHql6kqWsG1kg5137KdciChk+B8Li7l8z6ik
MbIuvHv+o9NZUuA+IKN2NAIJTKgYlU8iCBjHQ2NS/WJgqIeLsqIxfnjdOZYeP+9p
YXbxLFhx6TBtYB0Kg3WShISn1S9pO2NbTnhYVm4O3Xq9xwty8EYauW+1S5JxOxas
nWskMMJwR5PC3qj2iPSFH94bV3NNN80o84ZjVa/ESceK6IOZN8dw1+Xh1FeH3BBO
pLMr8SCO7n6QYB7DXcthvVG0m7THCV1t3D/tQHy+Y9E0CD+M0BxcdcFgi1jq6TL0
X71wvp6ufRopyz32F/vuMPHnu/7n9HXsgaJnKhyiiamZfE1mvzf4onJOgGcUdcQM
5/oCvwXuauKJRjuVlZ4d+99CXCSjveMAFrXnELKdP8rjL2o3jC+tlWJNz9TsarE6
btfw68yVVA1JtDJkJu4VMn3e9iCQ2/6GqFykD0YGtXgwmlyx282vz3ILUVNFdNqk
M+ZZqsmv9mHbbDuQrQuFqtKYr472h/XQ8vHWYzp7ogvH8LDSCmRDSHQUF840+pme
NQmjuZr5nwRMnU9LUE5eVckJilHaQxZi/cbVLUbGW+e6DAJ4M1HbKUoLyl0Z4czS
l65ggjzem+eZd7VpeYohtPkTYk1RlxIBzIrvsR0iCeWt1zZkJDZf+XfbSg4+hmJ7
JpPbyNKwE7MsgGk3LsUIQiZNxJrHk3nsrmq6p0WNfxgW1YegHKp4uIdjUDXtq2nk
u6N0WMZoCE2oXHJgHrDJb+83v7yTvRIHmI23NQSjMKt7tAU1mc8HaNekAxa9ChV1
AirboiuGE8VYiHzkw5LBJqgNZaqslDZK/G3UUJ8KPBZnGuUL4XBTQhaSNdc2cPJ2
MM9zKCg4bQTaGIRU4BMSWYmipGIJDDf7pXZ4L7o2k31gJI825WYL6DraRA5hacLT
9DPSJWgEKsUNly/B1fBfPC9JQT2WIfjz5qPPuqmFPVElluzSbZItM4f9BUkvPvKK
Fu1xHuYkzaERfZu8BHTV7KUWUN9BU0gAVUdhPTKci3XNzXQhX1Q0AjR3IRyV+ZNZ
EixHFwMTQDuVSIb461K4E1G3wPKXKlHuK7cg0zEvxNPPwV2U2NTHkC8L/YKewDnu
In1Q982LqqPxXicw+9E5dNHoo/BiHimMDyEqq0Uh0hT5GOGf5u7uiE2hSdn/zRc7
LtoUAgXFMOpd8dGYo4yCwISxHrxSwp1t5mmdzbKDnsjYWR6AND+exGZ/zbsOqSrH
yDkNZQpyEokvtg8pHbuxztIRAfs/pirE2ROBlHioF2KIDcwRxKO1SCc1kNlyCymv
+FV3m6V0FxwCHhrMd4K8m7e7iVtD6GL43lrBGYcaZEzTJk9CjKfkcfzj9jA2U9ej
XWYSUX7MavgSUuQFeWdqvxWwmQFDcbj0PUWjaxii3zKLF6/VeB33iZLm8sk80zI4
yThSRlp2qWfWOzVo5OzNr4uXJ14DXP7+s8V/rku+uPz+sTXyDf482io25OXQx0us
TJyWspfXWtr/HuSZZ7ZJPRo1I+Dwj8L7JODmufhIE+R4JP6jVNno9eGvyZORT3j1
73Pt12b/+vo1TcZVan9gbHulo2L1s/Yq8BPPN4iTcHxxO647aKDywCrIEtpwUGZJ
FznQqeo5uEBrAkSsc+KYdLE8RE3dB+eyP9K24aEPuN/1ougYQ/MBF3YM7SFQY3ED
EZ/lD0PErn6Tv0sxXrRYE9cBd63zXwM8aKxJpUji2mbV7S9TY3g8Fo+6M2T+UO41
ECjueGt4EdHd/HhYRZYIkjdGe5EPjiGFmGooAqDK95HeGBaURnSfrBiOHevLKfGl
qHMmF/Il8nNad809BlTy5hGjM+vzv5QsWzGyo8/FW7/NlZmaunrvMaMtBtlgot52
26QxRo9nECPgxD0FldNHrgX9L5se+mFp8EYYdALGBCV88UDhRLGF6soCiDNdt4Et
KDVxnhSjyw6fIskYwDvEIwJY61MxJmfcIsSRdIOkIuLXdTrF5dHamzcUsTatBe4m
dfbMDDTJVIRlKV0ttSJAyyNTQsKKAiPkJMWVwMaU47ZlN2ek5hk8O36Gdf/Lca2k
7B2uu1RCBSemvYRntJ24On2t8G7C9/NJYD6rpIosOyke9zw57nJLXbt7JeSfcPGE
RirBq15VullMUK/R8ogH+brpb+G4aGRxLvaICbFAACdgPNgQHQ9jKeDcklPVrYz8
XYY+kjvkvxZfPnL3Qd6DkJRuaxSztJNKQdUjcfNXqjxHqqnDazaTiSe96ZmOsYkg
EDCIqX5JE8Lfac2nB8qf52QfGzusRf+z/KypVda4nak94BYCyK1f8x50WOHI09Mk
LuAx2bUKyELYZ3t36SxcM7eP34Rgnapkz2uAro8UQfoZE4SGdupRcba9+N199JAT
DF2V8tbfdb3wQmC4i4WOQP/q+6FtBTtq60lAb8u5u7FukXLuaelKARJHD4p/UgFq
caIqECtFukMgZufN+kQfvPqvhJrQQBQplNHweoKRYb1cdjINefJUH3Pg+IgTGLef
6kHOMjkwsUZzcArcRgwWsvF8tu7fFuenJTNZnq4ED3EsEiwrQIxT8sWwJPI2HIyn
TaGd/xTTiEsWEwcTn0/R9srPkNSIZd3qL9CrmknGWUFDu5GKqHpd06etPKU2MH3G
R+l9abM7BItL/VYRsEGGW1KfHD83uDTKaUT45ybhDmWq9/cwgSTrgkp0zQCvoZV/
CA5bP8RFlxcCa8C5e12vnzGj11oFrKjbXqqQAtjidhV0pEZMBdRm6D/yde4Dob61
BYK5uQ4k1m7lLsFP99px+Ya6tsayAOPptCt3u72mIFkOrfjIo7HXyAcdc0SFWQ7S
qNblYcDA1IQ0JNxDfO1YZHDmxh+5WR+HUL+jo/OSGNjwmFm58S5vqcJYc0HoWVpH
DxnB5aIdSYhVlfOMNFoFdRXwDl+jnqX8HRypqJ0Y2NjSN3dktSq3w5idp2K6ahWn
+yilHaFupbMgR1sm5HlkDoRlBV8mZuIqVsd8s9fzMGpNuNWFNvuiu4a8VPG6RQvY
U6ja9GOVTvYOxI1B/TIKRkvStPxPA5RMe1dr79xlDOQlkHfdtVphv3FECFIfToVF
qIYuP7uTFTLAPvPQjKbzA9XyYHFmr4GwEmP9eZTHpcWlCkmvmwVOI2OT3BTTY4zk
9KtlSTy1VJHRTv9448vqZIYcShrpLowg4nzlAkFOGXqLRrg6ZaFW6ziuX+YIduDq
uOVpuNntsKa04K2VAy0nNh1mdEV640PLCZspFJOu+FSLQmcexNibB1d+FmlbJWuD
r8U7+fqt70cgCdPMl197moKhaQxvMplUE66Mc6uXu1XCfdEQYH62rSRV7bXBTB6s
O2GvGJkQNvOlYkw9gvwxsjTiOdT82dp0kBxD2KfvAiNrg2DyHYDa3gtW5yew9qe9
t063TccIZhwu7M0LvWvNbb+eqvqUiZiUXkG7wdVFyCsWSpBRud/DDPenouD9RERN
U2FUoBTclARQUSjBl8vxs68XJSg72xnEilbVqa8CRZnPEe/piyCdp6ekOEF8XNYH
KZgC/ixetA5W4ARzV0uoA3wCdT8AIc+/ad0LVSg9gW6OjSZHwNOgdAF3wXE+yBAh
eRkU/XLINiyCSE/uYSXaVjm5YqN11C7Z9Baw6pnwBHuA4RuQGD3ZDgxf4QyUzcCt
U2/xr+VhnMvF4FGLLojMYQITSJfcOBRuGAzJJ6xyEr5ZzCYt70R5U+6poFa8ZXtq
l2gXmIfZhO1Qb9ytAnowcYqCfYlWpFGt7qru06HgbZAJck8qRQ+F4ek0XE4ukl2A
gq3Vz3V396TSl3pl1Vf/LbDQSbVQMuqmZmclOlD/1lB/jUBPF1QiXqcoq9yj7YZD
jqV2YA9os9mRc5I7VsQFA+P5R0AzzAi/arXC+kDqQtAS78Gzlm8ZAd2rwd7lJdI4
ZFIrsMeo8h+isJ4e7OxWG11F6Nop0OC+3f8iCDSwFiE8nZwAkTOpP8O2FoD8IRaF
yIU/OtQTvGvyznfFn3hzfr8wiLmghbahgGXmX1p3P3kNHjG0jPlgoRAwqJkjM2JN
mJu5XHts/omKmuf06xUpL3tnC6+VQjp0H0JzZmlg0IRBaBuYxaQfVK+4Qvh1X2Bh
DiHgiS4ZutQH9HRSTSrUQCUbix7OomyBVt1H6UMn8AzjuWPnIplOFnNn/FFF1Caf
778rmhfbZ2NL/Bf2JWPu8uWqM5oFbAO0v1m+HTk0Y5M8yrRpfIJXiiFNteWxMvUQ
Z2GqiMy3bpZ1vJjqPgRzMriO8TOtJGdCBmhEpNaryMehDK764a678A+3QP1F9AZv
e2U9OK4I4l+qyhSFp8MNf2PNElByMI9raX7Xuf9hDujFESKeKVxk6vfr85Gu+6ZR
hef/eNCiW3xXIad4EqUwwlFuvrS51jnfo3TfQnkuyX+0UFt1S8pV+ljOUqJLl5T4
Xr0Uzg9M2VIMO6h0XUTtPph0hVEAV36oMj8uWVAh7X/WWeQHjmPcJQ929kEuO3Yv
oq1cYdInNK2j7MUiIJV6DfxOpPyqT7VsZr1AB1xthswAws7yMbmF/v7FdEaxT9ml
cAHTnPu6RT8/vwcBUTPMmC1FcZ+6gA3JuaOXHOnyMI7V4sDZx7np5BgWiczSSwgD
oVf+f4OMtINoyHZ2YluYjlPaSu9qozKQW6rgXYVUgunmykdTaFrEiYJ7LHnKdcQR
fHzWGqog4EwyT4cZsPEOd0Rk3cJBjmSEqM5Os/L8leLHIo8JrqO1Q5JOMFguD2mz
7TgYoXOaXjLXD/aizuoocKPwteiF/oEoyYsVFnPyiNkxc4cYh0E49BXKA8GiEX8c
g3d0ZN+2gYks9syqe2IVxDSmDllBBpukNcRUyaMM366QufM1JUqobtxG6NVxYi7c
hiSRpJGuk+xCbCRyrqoSQ8ynbk8QRDXX92Up7dDguqpZWod23jqRrOUr0NsX3XfM
ZPFi1GBs8KVXY+h1tOAOyy0UJJwmjifPA9BB168Pjqa7c6OdP/F6+W4dB3njTL8O
PdOW1RHqaI1Bb8gbDHOxPIwvpzIWM8e1r0XqWRs8kxbzig7oirHbxQj4FldyIGRt
73Lgukyn3FJb50NbqmZ/ATy7fLXiX9wwl9iGlVlvqPvbUeJQbcI4QireQbtdCePM
/W4qDug5CrVWvLLFhldtxHzvhCGFDdt/B45p23DD166/0IggKZeuGvUhEK6JSQwQ
WwqQKBkTRZCADyoZfNh3bdacHrhsS4pwYdlkMwuX4dlTqVjqRJOOE1Ftx9OpaqrA
NMwZipifmfJewkvp983mU4envYwPfu5kkPIaP7BxITMIt7/Lds8n/JGkZDk5abRR
zosM7D1m9ZItMF6ywFp4YT2U4UrshkvaO9UJrLDxJ8I1WRJsCwObi8HPNXPAqBTj
YDy3rKXUWwDVh4pKRwdVDl9vTquxMkcg7gUVts+MAAoDgNGKCKypysh8KE+bWchw
IcVo9SQ/6WJDaYjrIGVTMrDb+JPDGUtxeE9tIU6q0bO3ZgMkTG4wEuh4KUn2bggd
7Wd9tRcqnY8rt9UPlPSXvDN5lSIupFxeLlVQJEpa5ueFuZAJPEl1OReBdmFs1c/r
Fn90PZKYv3ZecHaSfdKffz97VuvcWgbNKy5xjE1b9oGUGkcHLb53qDR8dz+cmR4g
xNn1lAjynMnK1molQI5uDx2ZjBzCym+wnEUtDWXykXCaurgVhV9WMM4Svmej3TE5
afoqDvc8oioY14VSALsGIhaPvrp/C7MyNvzS15QRGnLGrLtpyJDJ4OjzQesIg7jz
W5b0heNmvV49UKPXXdrzwWYoKsZoa5UyupxIWdihJxACnJwMHV9xxKvi1qzo9GQF
MdUqRMvl91qfQDEUutfhAe2SJQPgr2lIiep/Qvtr9Yg2MZLCXyF/RtjAB64T1oqc
jrQA3oN6AX9TMKL38u+SSit32nGH0pCl4QRJcZEiZvAhue6O/xCisHhe2Tuy6Vfl
5lnfsOCisYfKxMjVI/0Ir6Qpv1f85KB6Aii3a3zdOZCfrLCliQm5xkIsztrhxSwk
eXEbpJ60BN1MX/+XijwTjBfYOIvQK52r+1cUWZR4l7+W1UW7+xqWWOW3wuZ/EVB+
dxMX422j5GNt9hrQmyIqv0l9KweBRx8sKas2etKBwNTeLYqucHibnRexeGgRvDgS
+o5qPz0KiGYddVDzjE+E+EDojgnsklWm3rCefTOQvZLCTSOO0KmBf7MyrF3DrFp3
t4EZHKOofkx10bU6yjgTipzhkuk1cEYzoPf/ougxYbge2cAehg+LoQpN/usAQMKe
h3p23mJAaQDyvMadWJmvtNiiw9M0tDMMwMAWVdRXNBmI4STf6Tn0xi/Kr4fZ+RUc
k6yqBpaNPKqH1wgg2ZVZNeMbHFrvvFA4dTfloxn2XiNPOWXqKzSI56/LExVdsDrV
zK0+ollUT7UULJ+2F9n5CCoX5XX1D6Nhupi8JMsQj5wK3VTJn/aR/T4hO7qg9iul
y31mWPXLXGIBOc4CitK/l+ulH9O798z+zZAB/c2PTqShMbqzohObfKXodYh/R8pw
TJ2vty5qIWI2MEJESpmnebv8SWTsrTkIu4MOOqA/O8dguuAmQ9j/Wmk9rqED7JM7
haS7aGvFnHbHo8ktxR6O8FaAssofQL47Nv5vCd0MnQtoyeEgRXll8JXpm5rQNlGE
NMG/gqXUWzZxBpRi8b/dPEfh/+RHhNv8ixsmPqAwpjLP7Dsdg37h+nN0nZZMrtvK
RCmzGogiaORFYIqjcamD1ICb3B9FOpiYG/1oNG/nEb0dn1jJ5I7NnHXKZZzP1SpD
85csM1njnENp3uv4jwo425wwIXE/MWTweFGURnVbQe2i095lDsfv1n2YkMOzXYvs
8gNVj6Us7vS0T8DfZuYjVZQ+TyXp7MAyWJ9NTLOqXk7seDCVVeYpC1b3RLYUFW/2
6afgnWGk00Nxd/nAluJP2wEa4S8liDeW1KwGiXmds0O7P/oOAR1VB0easjV7aLDo
OprjNPC056EwkFmK6F8CRcsF+WEFrGQbk3+FOrB3htWPAkNxeTPYM6TabI3DMnFw
rp6i/6y8makyUnEtEDXMm4PSgiVV4xrzJCIc9Hi5lhbFkdUeeGMAoFlbICLzc96h
/m0mhNFLajC9Ppt9iytEP2bnFl1HEeOUhb3ZKrxB2XDkkfZ+lZn+0g3VnPNmV6sq
LNhPYgUlz51pONSRXHaiuN/lbvLsstvQm6FFBZwVHo9KTvWRtDj5xxuat4uIyvKo
11nSOsg7Z7Pg420RQZ+4Byeu6Teq2sgHaFG490QzhN4OgTp2T2Xw8YUud01PhgRK
914ui8p0eR+Ef5dAPVBtGLP9l1EsAY+GdnUbvIvYLeojZJZKJt4R692QgFnQRG55
/hHWQ93LfBK0K+9j6KsfhiatTuOzPxolbzVGGYZDbgUm5rza9bNMzvIftMvMfCGA
4hNyo/kerAhZlmAG2L49O5f8R7zit/GiY/mQjsDo+7mu5ow9aIKA+BXKt0o/JIVF
54163KzqPxFRmEgi7xAn5zKAZf04Q4hNHASgYuTnuhHNxpMQcQ6jd4D1qB7/bUUE
epNGnMwMAI6yjEp64364CBEtE+i7g/grsjwk+0ikl+LyaHDeaEsI25hvRIPLEXq3
kWL6BCJw7YgXTrp83jdiaDGrflDbG/Qy6TRJjoei9GeQnP/1M1M9ctamDLF5Nelu
lXeky62SpLsFt2OoUeSgMB7uxq7cNuwzhMf9OdYQEvBYVpuu1U9ywKynjd6heF1h
cCYZJdi1VtLZxM4sBLhcJOK2VQk4JrfbPMwaCsNXfYixTJo8wfsokv41f0eHndfv
vGKWUHx7eWyq9kCB9SNtwOc/IhjFCTnTWa+Nky0RQ8grROe5paWJxwCD6kbMw9pO
pt2KsEU05yNDfbXblveVmvEoOt2kAet7LW9q9NKy492TkPz7ugMrl4KfnYHi80fP
JnKSI6BbhRokjHsJyp95kTO3YRKLBlrzNSCV+sFeZzugWf85kXvzX6dh4phYPvDe
4Tfn2kZnXrIeNHiJENXaOF9FZXENzfthFWLwjwLfwKgWbz9Kx1zL1bErkLYGhVcL
5dHv9vA1pi0xo8Kk1wY6GRdctp0203lwcaHJYLhKadgdVBIfAGCAS4DWMNaB4Kiq
1bXH0pU2AR/srZ8ty4CsLsI+uqnGZgubxipuo/HdsOkLMjm39BitTuG+q/VyL1+w
6dSt/XBNL9RujeyCs+SomxMxIap2y8HiQrhWcUC16WpDLmiLpPLdAHG8mkH1A28J
TJELzg7+YtCwUqBW0qafGx3F4bjvx9sCPsLB8hbE5W8QG4OgV0opEfyiRhOU3kcZ
CPpjq+h2XZjbfLFf9Q/BSqQx/dfecbID+WvhTCBMXEj5s2NkKq4mMAKekgym+tdA
xT9VzMCh3nSswfPvxChHAMk5VJ1QBLffPYP0YTntFipiNGlQ4XXTe+LD1lpU6FXH
kq/sVjeJWYpIRJV9dvdYQ4y7E+hVcHiJw3HchUi6xmk8cRCoT1Ddi+qzuUYWaeT2
oXtD0yYAWJVqha9m+63KkA9DFREJAzNCrKjOh7lCGhONHD5dhzztsNWUlBrOYEvA
y15tWH1tXCiU/SX+ILFRBbJjKgWf9nzlMMKPPASuZAVyNfKGuiBXuorp2P+3OIf1
H09WyPxXgUzh+bLR+e6jaKtnSECNiNZ1xC6Jl4FB2/Kfi2PkwA3r/DMB30B7xH+9
Ke1rmbsEYX57rIeODzEyNq3LrtYwBNLEk0S7eYD1n7/pA8z893Gpn880EHKUjmoS
jl4PxJB0NPPSto1/Bt+sm3wnOh27qXhV3QjirqKlRq7vJsUNfFidbRCc7cDiFaGm
c0deSa3NWavtLTWC49WAZh+51VynMUNkl1PfnwVKL8cM1CBCKrMs6n38eUBghYhm
rf5hmP09Ygi0eqbaR/Dqgx5Mi6/WIDAfcCfEwA0lSNiOfEYK4ox/G9HQwct7WuF7
uyKw7vHSKmMjvgPfNRlieDaO46wAJi5uzp8FuchMIHjo5JvFc/Isj5iVDPc5agdA
s8deEVzJXAgbyRaclD0iZi2uzwS+adhUjqO/luW2PC7HJDdD+d3hzDKksJowyQSJ
X8cDxNI5unj97eUhL6xb+lyYc1J1ORMHUr6ODVFA705VY/1dgHNMBeonfO2kDmUQ
3qZsfbjkb1SZZDbfACZZWeCzlTuJ/KYCjJUGQSj0+7oytWcZfh+oWJ8V3114ZpgO
CqtI6xe3lS0/zq2/sQ0NyUyTSX+B9ZA/e5EN9+l9GKGevpyT4dnVIgNL2crhN5jD
em08MK0oGrLjkRP94y3XY1Ee4fa49R5a810xwWOqgBoz6Se37aQw2KxGL4/4iId3
+MWXBgQuOaha6lZ8LFQPiP/gFFZ6j9+JpYqT4RRJ5+LnJxOqeeuj5Js3x4t4f6ES
w/fM3yFTW3IbBlTVs8Ib7Cj6Wg5xB5hH6yD2ULKuz9z5T1otSdxjz0ad/GQKaNeW
Jn+pc4rmN6cbdjqvvR4AtUAzyQ2/KLfxrbbarg84wyup6jcysdkbWDwwnFez+Di6
4WPdB4f1qiQpCkrbw/Xo7H/TcpE2LHldfEt/ueROaowbxeopNDAyitGutgkDsfYN
47zEBB2kbo4UxP5K4NLjwNAHqCH5QZ9CD8+TrUu7li4/+g8k1I04euMjrR7mgfMW
EsGcK3x9cCvsH1CGFpargCQxuxpG2/XANdtdaoqm0fIhIxqbHUnVdMVbdstyE0/l
/aehsl66iIUq3WUjBvZ5HnGpQgSQdzTgVHz5rniZOdIOd5Wkl+vubpvZ/8w48XI2
naRCHHL1GjM69bFA0zN7IlOSCDN6EslWhoRHyzzlT6VNkN+qvEktKN7Or/ypfau4
F9tv4TDFgdc9XXloUqiQW9/oHss+EKMQ1a8E7NfNNQqagMqqbUFb1w4Yzl498HQN
FQ+Ar1xhJDxS2DNaE31moSWZoFurBAJOkTzySpcwku2/CW/qwEq+lQdL3hSXaGIz
4u6N82C/L0O980frBv1g3xXc/bssH2C4Ot+3GiRrCE4FeIzeCdqhSQizaSUS884+
T9bR6rwsoqjw/yjJkHIMBt2wXs5EyVNFEAX+xPXXQK8p/4juTW265DNLXF4GysCJ
t0wK8dFX/Z3xgocEdw1nXFt5gYmWBDbX4jWV6BEQa9dqVcBpvJhYUUuXHIkR6ydQ
4t+Jtf/BynnacFnSZcDTrKDACye8IFzZdNDy3hIzgEV+WUc8XJs8ru9CQaulekMz
kEv0zC9Cy5pFzkc81Grl3WVuxaRqEKO8xv4BNOV0KzERGFTlTLuA6bF2vyzeppJr
lt8oHZxrs210hfGhyknhMxXgsF9vAazeJrjGVxYCxWjP7vTE3ZxbEeLqqHSyyW3h
HZDhpdCeFzEZQWzprCDWoYn1WkWA0nneNAXfmN+1Iw96I3DLAqPExAf99QbCIuAm
p5h//bG+4rP4WtCfy8tP8opM7FkGwtmO2AXJpbW0RDlItKNvsyj/GZ2YmZOaIaZ2
aAZbkddpYVDijmpJVsolzEWzSa76XkjjvhD+WSFxF24BnRnEtBvnD3d7noonYTnp
ZXFne+o4dD6A2yMcXBpfYZ3rwwP3Ye4F1TnzK0nK14+tnVqvc6dHuD0E+xaRC5Jg
FZEeQc68Lj218w8fFPZF7HfDkeha+eyrhWCbStvWyJBLaQnfqWuJU0i8XUPye8Kp
sGBwwToAsrcV44nyK04gg74KVj2UBT+Qsaspl9hAX7y1yyzbiYuDjUHFpvYpn02J
ZfzVea+nXK5iLe59dwhNL39WvHG1B7/OV8YI4nPtYXWOKFtW55+bSP4U/+LyBDkh
ZDRbRck81qWSyMlGcDa4QvWi7D7Q5wgtYpjptd0a26nU9aLbZcQsF4TGP1XEcpZ8
9leLoglVn3h1xx6/5WVAdCs/4dunelRFOzgxX9QDaF8bjFZgQgkd0F9v0Bl9W/Yc
OULRqVpe4KRFKgt+09qj7cy1AxVt4F4qbqAoc8nWbA2vgN8QfiWsUTK0rKmRrpdy
nzjR1svOc2iMnv65AgEBr1TkYicN1bCTp0yyP7V4oHV8OF9VyCbfwWzBoIHHc0Nq
EneogaE7AYRi5pVCIEkb74t8VrlXnAMpE5NaiFLzjbAVngEo8a8TYQfmE4Or2dP8
xR/Gr163aHT/BRm65DnRPFcVwty/TsgJEYACFkF78d3Yk9EzzfCRvH2RXl4Vvy81
4DU9P1aXXKcLODFzV3V/lrpC1HgscLoI35yqlaIkSNFbtJE7oF43s8fCeSgJBqVg
UmycG6DJOCuXVqQFkEv8H56K8bniebj3yzBzueVJcFTkrK+8Yic2V+mLUOfEVjki
7xWbSQyeMq3vqOHXcCcmFi+n9OgdQ4kC/M0h9F+VB3OpkoU4WUbUu2zCfXyvGzOG
THCoTmIPJGuHLWQs2h4s5Klwu8OGtpZ7Zter5qb2g2Cc6hAgFQkNE8qEOrswe8iF
6YG3bzwoekE5dqnThlDNFFb70oL2Jrb6isc31dAPEib4pGVbBzZB5hN0LmcAAv36
tjTEbKrEpIBWcZ6eEaNqL3gPG0umnN7YVJgCRu5FUlyWicbObH28UOa4kyXwJP7c
6PeEpAqYZxG+5Qyi8iIufr4TWAjk1mA+JbAXbsyVTH8yiISKwucLKQjJL6jBPiaz
8EQqgqHNaZQFxzdW+gWpRNcucB+Ug0IPxkxeBz9yk19AaToVkswnGdr+Wz/qyJVH
AF/t4J1Qk0RsBtOZMjPBBwVVpCq4hqrWQx/Pgc66/wkUW9+tPZ+CYHXPOugRgNeT
ZOQjokgZHSncd+ioqrCiW4sXnz8SzHO8rNlT/Sih5RYVYyPig8jU97lripfQRvzr
wuPC5YYelmc1JqhC6siUIndVHuycW1N/cbAC2CbQURDnCrdoHIIoOpGDa0uwc8AR
yxgHbftJKGXzD6+xLX47xh6gGeQFr7n6HWNVyenqV92Wpz7lKnPM22NGp/3lMP2h
IkiZx2RrJT8pjncsepzL+ncL0Vxum1vGmYKIDP3tc4q27H8o43erIA1JOc0OxLA0
rCdLudIkwMVVWgZpdqFvuKvtbQL1PSG6uoTl6K8r/Wft9XTD/b8/jYNCwIJV/ZG+
vsyHvznJy8Z6yZ/UfJ6XvNoc17aGu38Pz7AeT/zpDtc5LbCeY2vuKHmmgiBjraj9
H2pMIcwsTCWWE5MpWpJ1MXhB/6bp8bxqg6CpJcywvXj56sRJ4MFhVkRQ6RwmkNYY
FZAXihn40GNNgr5+yVtFJVxR9EH9PCKoP1leJBSRLkaAwBX1koNKX2/4qIuc4CoH
EQogcVYDCC4krx1u33QlwvL3T/GI50gnuuMhp27EZQysHQAi2NF6OqNftGfxG4O5
oEStTj7fN67dLKQ01d/ooHmDBLnFAcL1ZUzmyxDhqHuMk2Rqu28zDUcKhyOdAf1v
bv2nXJtA/cmBiuirLM5ePrFxxtn6+eHgACArQPDVzIAFt7s/et1o4JMWhScoSuUz
F1Oup2ZHXHSvEKy2Rt07od/43oGAZZMZTBeGzglQJRHZT6MNTStWa8ypMnY6GDNC
o+odDJgnpBJnPIylyhTBwdexW6fHu12RMTiBYEDcgT51K5idnAjhhk1gjf7KFQ8S
AkwsbiB3dobuWaslY6vvP6FTz1X0yrD8w9n5mvtgl6B4av+nQzAbO4fCr4PXU5bC
YIzpIjnxkdEegDDPietDFM+D4b5w5qkpDaiJtEGosBjPJugYQ0V58LgjYGeLil7Q
LfZSH5CYY9pqaBQWZnzu2folIZn3eHJYtMdqjJIDCEmJiDwqjXq4d0HiU9eUp36b
LSsvZG5H2euZC//b6XFLZYa3NUcMhC3C7fOQTOYGWvIkIuS/h6IQvVc4eC4esUDj
Gq7WZ6d5znkoWHnKr5MGRZMBaqxyCZcGRIeq6Dm3GlEIoNxt0vOk/iz3l4TVsqhb
aQUEeG2ZhXiM4P5faP5ISRGniCBEVNVq44eG7lC2PILI2knw49D3fumAItseEstq
oNBJnn9BkdHPCW8Mcvvwtq+p9UBectGLuOoM2WCnGwl8LZ4KRo/nNcsQ9LWMRGwf
VH3fGDf5b49/S3heoj/b8N+y9gJ8c0LYrdBnffbjX5aIAsJAU6SJ75AhhwjOCcq3
BNA0dwwQHbHsvV5aC57AcEccrw4SlHUeFrf4Ha5tGhWZg4xMoRGomXJ+exKigFvR
wIwj3Pjlfm4QwN5zZlRKAP5T/NS7C79rGBzPqDXkHU5sLP2vxIVHpIuWfzy0P7Ln
EDcIMO6eJKY2uUBzW6GGasr6QVMKV3BdqY6WetCGXGwI31o9XWUO7plJUtYPrN6y
piDbumpINbfiaNzrxBAQCzumKG8jBt/lKc4OkoQI2oNoPunpDff/2hMs7ghiCopM
7GsgDQ6MeavZkQCnEj/m7VqnOfwstGsYxrfOCs2HIxhifr8MvTeAkyBioV3j1AKr
daZgioQ/7z4QPKpwePAxFF84DCvBz9H8eBTDnrilJ3kqeCMePVtgVTFGohNj8X6C
HjLvQoa5YEQerbBh/uFiQ0I4U/1U4pMdr/5OKienlq3FGOXJp4O0LamEgOu27J1T
LB5G2rgP9FdQzIZPnV58VF7qklNsCQodXpC/WP0cNQ6RV1JzvzRUG9BOG8ePse10
m6VmiSfMeGTCBqeljzyCSDZbqswm+9bDK/qWP1slRC9nwaduCfh//dZvbK30/WOw
7q8AQe5T5bjP8EIQPVkUUDSnqsDN4ToEeJnN0+iYLaEfiHVwrservOLBEd62TVlL
BM2Ov55dAgtrxq0wtNrQUXQPLOgyBnLvN/OTJgWPMhUTePMGtVOkYTBFGCSnvCK0
nTUeffz4fO2032PweIiEXJtbyvHNiG6vIztBo+WFWncxa4tmGvWvbAKlzdSOSKXI
pIh20X/e0enMwUEY3bMFQzUv0IzQcYjkgA2MHcCKJsr/bGcvgFgxHpI4OHlJbTGW
Yo3xJaqldGWbjubt2BC306MDLAHBpG0qkQy41Vnq1yRjecDL9UJqBkbZu7FlkoxL
LpftPlrKwlEZezamqEd1lzkgB/Nod7Ob1z4g3roeHHLu1wnYgn2QNjuSkqBkjvOJ
3dnNeMLPElCx+r9fWRKUYs6gqkHU09xFpCwAjlGH6+90WggCSknn5Im5mxkx6dv5
X3lRZ62OKzz1m8FrXVYFY3XXjgdpNiWbR9mO3bBOoHKFtHA1xxqn/vrsuG1oyGew
h/HPKc9EGQZCpzUr4TnbCaRttZ4VZPWNXf+qfIdSv2EdNot03kv4kqdtMdLwjY5V
BXeJ0Wp/NM76jpYB24LaU+IvBN0rxzk1BKxl0Xui0+wBs6eBGm7wrTq4QTsutXYv
7D345tyrdKQr9OWJED9WQOB0jDqHSvDKj/n3jFNy4dRq+u1GpxRdh5WTD5pid4bl
B66lvJbFCmw09PytpBQgkXa7tAWUk4B+sRvyiV3Av8mg80/KE6FWQJeQ1Fsn64n2
tvJBTPCFfeVQSEJyrYlq9cbvhuTy/lYA45qQTGnI6vCvD5/ob0bkrl7HXeeKW0A8
xqFAUfSJ/IJu+qV73lOeX0Y8ftfcBSsj51NArQBJrExW5lyWItWdo0vHC+I1eTA9
zhkgb4PV25A0DYvi1JNCyrZGlV5jykNqPFgM+RH/cXHmiMeoE2vmDOsgFrLHghq7
XSxK3jl94E3xTFjUDF+IAJOz734tUxJo4Oy69O9bgfyQf53K5VcfBo010gJyNJGM
oQIX0qt+yFSUfTCftF1t2vglQz7DI6+fYWXeliu9PEMqPEL+XpUuz4IdZqtlIprA
Yzt8AxxNf81VjO/DFZdN+r51H8zZxZ0x03xmyfkPdXkfNcfEVRD6C4HJSR6UTAsT
Xp9K021czEuBvIsJ5zCuJewFbx90Lh6CPKgfSzsPl0+rlEdMQtUr9EMR8BqHaANl
AETBd458fdT0fJRYrGcFdFyAbdlkkIFLzxVMV0Sqg27RNBmdyJf9ba33Fs7aCUHD
jYiw6BsB27Qh8upfw+6oiN/VodiilGVUhHjbIjOlGbxBTwap2RTMydF/wk7nDQ9p
OJWZqZFFNGD9PLKVLiMJ3VP8cCzY3JqxEfplnsh/90IVFmcnWMaO8dkocc/51UP+
sG8tT1iO1YbSiJQKcy2k4Glm7pVkcyWAD1K1hFRGFD33SV2OD3VlAw2mjyBezk8F
JdfoSxe5rmUJBRP3goB/9O6ra4qhKku/MkQfqtDrk9EITGZBf15T9DxYT6th0ZyO
QnrU/JXl46h5ZZQ5iicCH0VA5ee6NiVpL/NJAC430KYLzxcvGOc3iy5Ps1+r3M+W
68UUtXgP8j96Ga2brO2EnORuRo6Av4wqYsG22q+1rqJMoodoMXWXvl4c02EjpWYO
0VArCflXP+Ukz5x1/wnuSh5AQNFlrrNBSV2YosDkkG5TRVW2+7G16uYGI7L7rCoJ
ARabkIAbmpiXQYXuUdI8vI4cG9ZlJiG2I4xxXz7V+vo2ULRFf8r9pqC2ccDeA7Hl
ztoRAwONy/IPpe+Q3PDAKnrw73YFlcJW0FNmunIMHL18/25rFv5azRpnJSsYxSbW
wJXbJH+Qf6KtZJdhnSIugUj/L2EY0uNhoos+gkMruEC0FRkNeS0UcjYpC+1hC9/S
pDvItBAz6sVddI/lsbS//RZu0u2A+vg3zLp1c8lOJN2RzxoHIsgj8pUOL+8tUG98
e8o1W3W+eEaVEjNAJArJM5QSbU9O5ru487BtEA3BQGxtI5a1gULmjjpDL5OTezzc
9k6xzHZRNa5JtfUEyfZzr4LxXh//4Bf9pv87imnkc8wzbBw+uzz2DTaH/f6z65df
ocjeYGXoZfO3X1JwOUYF/roXj2i6sb4YzvuSsPHA9UFRNM1qGs+ydsOjEnqnXP+O
lYwOREW2RlAy5ktJiXeW8p09JTsqTwTkkeJ3Hv3yf/5LLHNTb7A4J1+Dsj/Om3y8
/eWrR1929HWavJbnNQ7t+1RP6DenA12nyqp4vDBHDVCISp3ebicQ2ey78BXCzZNP
Id9hHjP6IiOw7vBYZNKBacScy/GshlUiOgSEKljZXEZfJFgVfpCIM668Rkbglc+m
hHr5Hv/7fAYAXyJyXWnCCr8Qeo7DL3nGe949K2mOGI/jgZdqFisqaFJ2l7nWT07d
4zc5ISAfHd+25ylPmSpwpUgzn72Nxv75N7pWt6bczCwHZ9dFYyWfDrb1Ix4pLLao
yQ1HTQUMQhKmEpSWYbK+FImVu1keLRwfffmZpicu95tSE0kshh6FwRPK1ClWxUT+
buhhASgDlUNH9OeSmDrXXypy644Zrg6+HnmrjybSfFMTII902rXCRXJToSiGF/Ng
eh+vQoDdMffBLqJCoRWBFklDhcO293jwRYJMom4d5MnLXDHVAeRKs0b4H7EwGc/i
VdYQi+BCpFUium3F7F6JIVkztcgweDnAIvSo3ViOAvHG55FQjqkFTnKgc3nl+kw6
gHHQUsnMkYqn/DtNWw440VXUEz6EyvJK1HW9IVBagfXE7whWDqcytRzUX4Lq5bH6
XpXi5ft6hKa22jnp/CzeHEBfSXx0kvdukNgb891AgiE4VqRVGK2mAB79zyvi/dmF
jDK2p9BSC0eVN8+pp0nKwWiMyhXVpxgv06tEZ3UPDbKwyugJ4euitYd+T9MhgCkx
liHnQt+XRBMQbr5oPzru3QHccCLvGatPRTKtvbp6Vr6YOZtqd0bpmV1ybWUjOcQF
qDL55kdPTSz+VD3q5C0aUNmh8GY2dFOPZs2xOwpuREw9g7vqKercZ17cmZnW3RiR
yqifAA5jeWcFOJCCU4tr1n66p/RZfhoPYkKe74CqPOgcZsjCOYZa1p8dahfw6sXY
ht3M78Kq/HaW27I26/SEiyZLI1AzZYkgzuo18LQHtdxBl/EWBFOEVylXM+eDhTCD
l2+5IDf+w1/KVbfAFfuhpbA3O2hSRZAf+kI9XkW9OuBVVDBDN/4KTgRUuKNR/PVC
3AGrkRqeXCgfEs37r+rJIUdO/I4vjMGsVUmMpoKlucFB8xLfOPhMOhJeJUW+lhSG
bByiDTisQdWkzLUPosN7VdjpVTR9pVOjsJfIIRWNuxR3dwmrq8MeZv5hZd8+N0AD
pC6jL14o5nz6Mrcwg68XBWhXLcz72+BKIWiEPfOZfnSkPARGZKDYtxGkrh8EaiPn
YWd8td0d+Goc1zxosm51B5b+zjJPXBlS6kwj9tWhnRliQOgcq2tGoADzVT2BTxY0
m5GmrQSp7Iz+Ia28zHws/bT5VPq/JGOoZb+wZUnHLS0ZW/Kx6m22jva1seS/yS6S
07LKtrUifJ7wEEoPM46C9qATkNzFUADtKqrIe6yHNR8XW+E2NlfiSx6QGRIb0AQJ
8jjto9xOoL8DeGMrR+IDy5Be5IH2xjPlYRK9ekxtpWwUJ0jnEA56X4dU/eBPl4xJ
06llFARuPBpdL9uP5ey1uwpbX0S2/ONur4IbIhf4WGIQSh/nym4zsmkZJAVk1ma4
jgHltxPaPdSzS9D4hskYULF9WL9XAriI2K5cXXcGpbMReZBYDbllwRCmjyAJx9T8
h2NWebWq3kgpS8ctW+jMYODH0XBxO4SObBI2RwKlNy7aMOLwrRjiLPiCUKBVPVGI
j9sF8o13IY33bAhYjVpO4ACq7hrptkocyx+o4WtvkqSc9GjbgWHg7rggQSaqSSC1
o1Se9SVfPzH2D/NEzpDY2BZzBv7dJ7BElUx2fKQiVt0XREOY1dm2phJuScvm7qTD
wv6G/mu25w2Lb4e9X9HP/T9AEfyXw9V72YJUF9oOVOOTgLAA2aQLok0xwmbwwmef
ZlyK7N37z07tGVnMU75WyjmVxQFCwXUk0qHnDpMI/FHENu3gtVKrDHNKI8dk9ChL
hKKM9a4eanlb7YCGG/LHoc3x9/L4u0uBuk5xgYj65McTAgnugJs+uJ1p3ZPpaaRU
DcxYIVXIDWmZP71GazbLN5ezD/OnxA1hOeXxpP/ECHLVXKi7JJEipEkT27heV5Ab
0Co0eJ0gVKIdADbyC8T/fruA4HSSuJPLcQ0egUvXhOq0h9hyBVSIT4l3cycSebkn
jvwB0GApat06dsrYzftpgXI79aFuDHUig/gsmzopZD/hqYO8Bh7kvynbutC5aSBd
N8/9SJygEcOdkw9ZfyaMgj1tDoWenHhFNYLjNLKpfzNuEyvDt247KnrN5xSk4NhQ
UPN5tOHcnllNPdIWG4wcJOzoBE+EdMgEbFCNNkjsNnVONB61mBJQuXW+Y0I8LrU/
6fWuclN5riL4McNwCtN/wFMz4PURIBJszg1TvmlvLlJ0p6ZJdKDfcAsCmBNqbsvc
I3hydjuQCqUNRx4yhAH/mayiIjlUIknGi/w60AQHF7MSSn4LscBykGUkIOH3Te8l
OYbTDV3kGDotoCrjGWKP+Fga2i+9EQaYcFxhldwEBQtoW9dj5N5O3ts2vKyhI/95
uTwtdhAU4HjSdXxd+VxVEAKtUTRf5SI2EKrkI75KEM2Hv3Itvv0G607cz5QJTEtF
IbdEn40gahHI6+Lh1+wS7xQRzGVnLm+3LYbrn7zb5D/M23kmt4kA2Z44/7qluDhi
/Zu2ys5WEXJ1R+yCAhEqP5vMYyzgJ9PSkm/kQ7f8nJi1HBi8Eiz2pFsPqVIym1wU
Ua7UlFRle+bJCDBvQ04XhcScfM6B6+aDOnMgyANAROzFl6fIQqVRlTl/1DNmoG4r
35kXmHymWeSdmsrBBdRotGZLXehAOv9/MmvoFiu9asPA/pK7QuJw1lwmh+dE5vNp
UP0Piuulj2qc6dzeCinTwxkMsdmAxivXaWI6Cq0UJuJ0wWZWAsJfseZfX83t9D6o
nCXad7wGRgb8O5Kz44KpWdtY7IWCHzMlvHYWR+lZSiLf8NNUA1lFaWwS3n6rr7PO
J2jgvCrKpehN4bWK2Kh+jaH98nh/QO1XnJkCEscWqlXIk24CF/NgdXT49hZBnqTH
06HO0R+iO9puH8xGRQ68DV0fKzNWkzoD85UHZJFKmSagrt2OZSUUSxkyp1WPQd2z
AyKZ0kmzg9aJbaUu1KU8/pPlzEYXfhCqUfBGdrTKuFcfmRTBxliYjmHIRdUd64mB
9oddRrCYJvAZ3gSKKfP2o9yWsjF/ZyStBqHX4s9sqY7WEVTfpPcl+GzQxR0Pot1Y
jgN9AwmQFKsdLW1zCxhobtqTt3sqbBg2chrTZ/9L4KQP39Xu6Ny/30z95stEPsZx
rddWapXieXf+a6yZIOMIXvDaM+qr1itrkW+z9ddVHewa467mJNFyvthxDIQoCgDQ
YU375Tq2LGpFRGi6rd73gR1Hu0LYsyvS0lQIXWBHvboSKzm1itjtCoKCdOwb1PdP
YOqWuQHfocDx1cqUU85SsmhnjeIlBc9pKIZhpcGCw09IzPe+sUCw0rvNcPGpj9LG
93FsTiX3X0hHZtvQTJ8rNAO1XLusgcDZy/AFFOr96GZs1Uv5bJPmRb95j9ODfm9E
k96/rAi+9Z/dh/UiksF1SSN3eLQGEQBfDt9lSLSFYK9EnqZMuwrxCTu0p6M45D2Y
Se4JLM48S8B7WWi9xMdoIxL5oa2oPLrUuYNQXez19nup1/+n4cp5DAdWwY8dnJjp
CeKFG+A6CEHeDa8zhLI5noD3cIjmy+O6Ef0zLmilFGfv7pX17pVyK6H1XF2UrnKo
i5APC9/xlF7DjOzzEjj/0uMHpqm+ixo9Tzhp7Fe5xE39F7Qk6GHPLyU4NeMpmBE+
QPcYC6CXyqQdYYWOzoelhLTCKkGZtieX/fxZcBeyfQ5x2907JYmF/b42UaZeT8up
LM4F3eQUPRdDCr1jn0CW5TQKNK/60vvkPmKJrG443PeFQjyGCNgpJ+HCezyPHkgg
F60WeePLhJF03FzpZ5cZvIAFnsUWg452Ki8XXAQu7nCvEpH6qjVLd6vEzp+LObdl
dHajCMSEVT+8sSjz2r6Tlw0Zhk2/jUR205lQPFUdSihr/ApwMcYtcxfbSyqK9thR
YNLuXiPP6KsDzUXIY84o4ruaQ758y1AmtbvPoTfmNHh35Z3hEMaoHnYvQEdVqpDA
1iZboUl3vWcIz6YTJG8Rdp0HaaNu47AUua8HGX0p9GXM8GW6XX/jFCwNdvsJxfkH
NpRLLc5zr+8xJ5cEyThz2B4GsEfvm19YQd8vUSa6QDOYbZ9EtdAK5sEMjpxdWj5z
s/+TndderUfwUPyafcIchL5MhMv4oFdiy27c4JrysqMSu9D7VW0vG6w0KJpilXut
oYi8z4k+CEWW3XojTJpQua7uayyESO0jwz0cBxoHa7FvZReTkEujcLJePzG6B/BS
+dW4NC8ild/wOZ+y4b25beEqlNobRHm7GJaDJIJxMVwd4MVaI5ctnA+auiJ5MD1Z
9sKP0aO8mKDYyO/BSHp7LbL4CfVI3w8qx3A6EtdwjaFilIQFe37WDI4sfaFSDV2i
jdLV6PQYq4EKAZ8iq+H5mWgrQY59ill1dyDarHnJH+C/kXTfXq4f4oVfIvPUsU1/
yltt2DVPLgOYqAYwVERyX4amAc+QShJXcRrt5cbyCala4og2zzeaHiUSL4BC6PEd
XWMC8c9sUscemiD7/0rNt9+maJONdbNC1Zz7NgpXHEPlvKNzNw9gjy4GDrE8XOz6
fI7NraYppKj7Rbz7tjgEekMgfCxItgJ8aAveG6OQ95PwU2isAARmssIg+MP+7aRC
YcmXVGhYj6i7cw0Hani20W8682kNyMZHZ0GhomCwEfsC8R8qP+ThBaxuFuIlH0Yj
9KA6lvUE8Oit+QpJnyjIElv0lY3hwDrlzK1a8nsFfRGxjLphf5ILir+Rf7db+H8h
rQR61UqYHJK3z2QXnls+aSyQBxHBm5qfvb4RiBfe3XSv0Hl7wdtzLEAjlL94aoT1
A820pj98Dcm0RmbB1MnLlsIeFi2jFA+P2bfOvEegP0AYftuIIxZmTmpRR066ppFa
j9ygdoLlyU/LEN7YsMlLNSpdDQ5i4r0SimZmLKWPP/5FJh0Dq7NNiisUk/NE6HbX
82kk2OzBYdr0PMGEpFgtVwDOlFDXyzD57UhqW6SvF5fOz9ofvlikIwMa1MCydiB5
prE42d4F0kZpbpJecmEEqBZggv2k6tMIGfK8YZTl2A/wEwQwAQH3piMYRlBQqVPQ
kIuzGVYR9b+mRoTL/Gspuan9bV3HsihTtDOTBc3Te46SllwSaZYxPKM8r+wFN2Dy
YgLagXhMtdfZjbUw4gvx1cBjTsdHtZBQwlYvATc0A4NasS46qgtrm4eSdyWGj1CO
nHRqxsQJ2gUGZygVriolu1HXtsINUPFgNVdFwcn6l1ai7uXODlTbj0R1ZrzGoVZb
h8jLCXWm45GNGANJ0MSeXZyKOCA2/bEg8Gnw3MDpUtd1BbfdPApunGnDeGmVlaae
VQbe4Trtph4uJHw+kKzLYtR/EOC/R/p0T5JCKJwQyEZRUwYG4gCoajpGx34rWOHH
Y8ZbhS+Of8hc3LKk/ATR7uKBMJP9YHNyraI9/mj8mZ2hPGjKXqG4m9BjvA841Gi/
5gwVVh09WKrA0iiZWrGMQATYntdiT9BgOxRvkGN7fSUv+C/cpvGFVCRuAii+i4rs
FqllnJEMVhKRwUkskKqKWFAk/Ws28JHMLqr/KOqW2aklI42Qcy8Za9MRo6zQCbsy
WfRjTJTfW0qdlM0hNGBQm8QtY18ejfiEaBLdr8Srkb2YOL1x8b5hcMryRN68Wt3d
8IwlG6MbXRi8HGfOxQaVs85LI/ckOA2dAUKRv6EeUDwZxHjKSo/8KiiT3C/zwoOn
uvLfKmSBTU7Vd88kbPnVlmVNgnAFZdUH/LlKGKQUmdLXuAox6Hemz5ctV4xG8Q3w
Twh3agVFjUhVWbJnP8FG2MF4GqAPxgu0cBKJUUYP97Yxa02ZUHYQn73hxXn9wuLZ
5TYsy+l2QFQuZ2JqcFlsp+o7E+aPKuZyU1zQSm1cRBl1BahD7qbakcMvEhop5Psp
B/aaUd0pDyVTWYVg/D+0QguTQgVr14LdhSza076HL/Y7a4gBvQbS0cXjqtINswLE
RD5oBnDV1XohyUUYyHqGna8kQjb21c8fPzRcPvfHg+FO2Y/vKPXlZH/DeDDjSTCw
hFEN8y1Nf8W7S+VnsLNsM0oE6PDoclVG53/yZAE7Yxo8ppQ6RqI2DkZ6Howzo8A9
B5ry/kmxhdinwo7Ph5/IR8tw/Xh8zq453JOf3slY6UvsJGioHOGdgY31cCqo3Zw2
kZbscBjlogrLBv/UHODh4/JWGWvFu9UkP3idtdr4czid6KQNeP5EDmKgBDOrj2WE
JW/1F6yt9QlDrAiUYprVq+BQlFdFpN6I7h8vu9Ejx1DQ8a2m6C5hhaUYBXuKZ300
+WBZ8aNJ0Ge7zEppjKkEAGLRpZIriamdBBxO5SP6KLlbxP6FtomiZInRI7RwegyL
JvONSXsZyJXWgXJ2iKO1Y6+Uy9iXnIwlAnHuMQaoIeK2UW1p+HMkKMnID9nri/iP
zEDBE4G7PsBB5sgWR875Oaw1YL+rrqP37S7F2w+IDbpccfictSaoOkZMt1B8f8u9
oGoe3qfgWEm35nP6bKlOgceLKuhxr9pQeHxAFb97GRhAny3XfDEvoiytBAEax3db
twYqsCcCl4NxiwWJ0B1J0b/5SxPmgagCsqftE97CJQv6qBCm1TrIis0W3UGV8rDf
yKjxBhVwtPEej/8kTUSWba3N3LSL7Un/Tv+bQBXyhx0WYnnEPhNGGGsVfUkpOvF/
0mdJtMNiRG99Sch+GYQdBnpebbxaFnsVzEeBS0c6KvA4JvUFGH9yMErPp0CcR2p9
XMOwMu8F8JyZJSmEKHherjewJQk4gpkK/q4TEI2HSxWwH48UXw6BqSQs0EycSpK5
T2LxW2F97UnW7qlQB8g+dXx12jlROdgWi4tXU6PcSzNd71JvZA0pTGHrkAVVjmWK
1NiqIuNe/57NytIHfS8EeUGnj2s0A+gUHN8EdGqjF88ADF34Wj9++np7hugVVjCt
NBFZ6LhINO63fGA85DC0U8YH+E4Cy2uliP3B0te2F9bIbEjHOh7Ww4D+J545sD/s
xGzc607WjVqsTZvl560Z0mU14UHlspz+T9BahGRU23q7MiHP/eBxf0NmKKqBauM6
cEAtfegKwE8m95AqFtlh91y3+LxQvg65fV868S6Zlf3g1xDGIjq1wpyv0hx9CfUM
UbQTv2jmU330i7pwwnLmm3xyK1D3uJRCJjy3Ob76bUJntapyYl4ncsq+LpnaJfku
RpdkR4AItydTzvC2/vh+AzrbEVhUMs38O67PwcG2EvadUxR0vAFdzIwXeuXTS5OZ
luGT2jpgxmq1BBChPnepRV7HvTAA9JSMDWSFiL/Ah7ZIdHU7FGSQpVjEd7tz7mpv
2OCkVs/tRWCvNp7whCBjx1zghhkgNMbpJoSsIJER2qNXxUteQ7O3pXr5JBMtMf1b
YsYK7YMBxIeJh7ecTw14tKR2zGWrcGv/x33p5FDGaDxo2vsXT5Q5956Ycury5igU
WY9U7xvfgCSeAQ+zc/gk2Se5yz7EgwHY3ir2JO0f6RxToowU7T9ZMReDWfBlZrM6
0H4nwHtlYgxElZAibHsgvNzFlE5kjnz8uR4LylCLvmxSZ6P5596ZwhOPCnRXKRqW
T+zB6wBtfAMUKZ4Dkub5CGb3VrUpu+WIQK7dIBCcLMWaBK3402bxP5l6othZyW/u
QDc+46wFAaVnfzYdlfrjgpnwLKeAk1SX/7sC0JxqvyDPfWPdSVOnnL2S1WDMikCX
D4lu+fhBvlhraLCYDrYOfyfUz8/jK+LubYwYfqEjTK/h5ltYXsZcHEw+xDD4U2uj
9Z4dOhobM2Y/vqlFyxdgmNUCHS6Qp125g/HFqBHI+pBx3RlZBxH/w7ZjW6Sxjo7B
WdHXvKylU7Y6eSq0hmj6Ibv74DWqY3o9rBV9/58lvebxUnQwgW54Nl5Ehnsumyvz
1+RzlTzgPhvllFzgjZShbUqjYk6tcOFmobSuNlVXpk+Tm8lylvz4eMXS7QhGvrhJ
YU3Kd0uht2qxjiDissNQ8DYnKKjA9r7luVcw8UY5j07LptP8IRVZ0tqS6j1nsT5E
jelyPh8UOst/l+iyNMGRQLPSWhNbdRFhgbmgaOm1+qrZIsWjN+0TOX9XsYQq/+JD
VE+GzZozCK9aZgyAbYB8dDejjGgQbwNHtmwJYPHoEXt5enKxMghMguleLw9gKoxD
sM7sA0q2unxCDXTreK5PVm6Yhp0qBKZi6yWOCDX8+i/3NfXD8jMfZv+nDVbiRQ14
EsmmH3zOxSpL9ks0tdMCTqW8PIZtokLQCXrPO7zWGRVimfITyNAGdscIYw0/Cvmf
eiL42JXXYtX1QnlIkZJyowufQTqP6IOqWp0DeouqPZeLjUbr3U2/XBr6GFDoXT4z
LMlOTMrME8JqSBHLMWT+NrGAZuLzACYCJt5fJTYfgLwkL90LA5+MLcPkEC5ZkXaj
bBkHJ6Lw48U8MuBfqq9FyFZSVmApqrEkNU/4brYSyiWZMpzypSI4BudZa61HT3vA
ssgg3cSwDRqdlEJEVE2IBRifLQmVs5H52G0flH8hKpV9xt9cBEO1g7Skk4Z3BpXg
86JMjDVt5vQ4XmmQvVmCa1Sg2QloH+Ze5vV5fZpQ479I1yZR3GkKtFXrDtzjlYCz
oy0k5q4EYtOcZV2odM4EkOD5qHN7phID4/drUPGzI23/xHEQLbtNh9pK6KFNTHfk
YYn8dW4NeATUEPy2NX2JzNE3+bLPE5VUlWVvQCD77E3hQ3ZGiz+vh9boLSG+wBx6
lBr4+uMTfs2C1U0em3Hoq/wtshIZPGKgH1cdUqKT2TriOLeuUWmuRTQMhhZ1MjDo
atB0mlvarehwGhVv+2CogrXRXygw/ijc8C5ZBOalVFTFPosf0NvOxYDmAttmaXTK
By4kcta6d7VzckrHUuaj7pUHbXmZVEt2LkhAjwsfH42J/t16Me4A46KCo0iw5UUS
k8P2cIoLN9hovslGOMxOd2Qoq6nmEBV9hnpa110QXkAGQS660BhT6I7lqSyfqWVg
u5W/mQzXosFo8qbEPdGiEy67ukQgHq3aZ1h/1MQAqAWvlqw+IqyRBA9VjXedZBUK
YlbVrSGdbxzR+VXVMPR0PjCyptA9kc0GPTRXi2RTkqHJ5Y2P/nQltjhkQEkfq8lm
Lq0WBL8ztXTpZCUuhLqp20/5rK63iosTvxKHjgxbswTdVDRaPgyC7eztjIZ9MoZH
vZzEFO/g/msxRox3M0Dd7hv+ll2c6mYWjiM+cRWhWXD/UKilNpkX4cSrRE64dGGb
D5yZb0Cfl+au1WsjEAbN50bB2kYNJm7qA1euO9+b4QaWPWVjUprhFIVn+MokH0Ey
22+gJHy2Oyd1k8jZmi2iW+yj/T8RBaIQbY63NKUZyJe/W4RyEfCf7COjgVrliMNY
EjpfQR6oSJb95HqxwsaGLcQ817txYxIvBbjmnQ5YnF/0nmfnMiAQPj91LGmNooHo
pFXg+AgdSP/qr3PlcaL0ansydtkXr+HMOAs/b7BykzpYICqADOKhOr46/LQXUC71
p3O6+FVMmU9W0YD4cABprMLnsZq6SucxNZnzDZbTw/Le0CgajiPp+wRZlcz/QomU
bIwKXiFvx3aGpBF035yALGCVAsneuCPKxpqm0/xpjUR/7ysBKYd2vG3dFci+zISZ
G0RTgY4U5y+0cKsvTsUPqZ4TRzpCgglQMamtaRAZWeR9Qb15eq0YG6L4Nh7SJgS+
o0L9DXoMBpR1Jxkl4twNOSdQQITNdAKjMzos1fSYw5zJgUti++MTpRKbdMTgb/pB
peswr4+0zuNI3mxsHqLpn8440ctSjFCNZxA4Ol/e9sNQkVagoXfTQth83F9OCsOg
bEFnWjUG6JxSXC51DAbZhaZ8CLy25A3MIfeI/mqPVILqzRvwt7lMTqNd7kNQ4JqP
GuNvLSEWFEQQi1P7r0tOjR/NDzyYV6vvJSF+U7OL/eylIbd7AmFFOfyuj+8hOfFQ
ePAefrSYLqZ8mTl5P7jdhLlqaAwhyQTGQEtAV81cN5QcOeXoYeQF6FlFClWws5Jb
SXTyLN2/DWcry0c+imtBnDMeDspPEmQRiAMilQ7F1V0fzsn9vWNmCKYLhNnVD2sy
tNiJee8vI3a5DlECeKZwFIZYSmb2df75lBNR97ZCi3UbXLPCTIdvyCzK4FC/ZFWQ
iiS0kYHllH/FIjPCjrcEsecGEHeYUa0ghFijtRNDs7X8M6O0OXfXMNLVTMOPyeFu
wd6K4Fvysl6TkmdxVU2/00ZqOGztBIod3rjbb7v4INo80yvUrQW/h94AtanMWY/l
9KQmL52dcI49hv3MS0Q7iRxc4DywY3VJLVJrSDe3cpz0yo8Cf3fGSvljsgOVmOv9
YZopP6MzmPE9cK1HKjKBc+3hFsYhBn4jXbHI1Phx4goqA8cnf1qwNN3I+EpXTXMr
iRwUfTZWSb/NUdSCDXLpZz1NiIMdkw0hgWoIAjP2+bWqcargKh/6Odc7WVWIttnc
ZEEr0FYq70VpzsoTDIdPg4eNKzgZ563ATQDjq1SioES6vRGkYlvtZw69fmsFouzs
AYRTfPfTrwFj2BHoDEEnacIJyjalIHJnRRqPiFfqYDkNjmHHLJc30qDbN2D6azxx
69SIOkHqfwV2o/yO27aD1saQuXtwoAwQCYFBzwcIMNnPikNAn+NbAycEjqM3xZr7
6GeKHmXhfzZYD+COAp/GFXKo/06KEbSD7VghC4BIBxphUJYtYdaCugUZ7SwRboo8
PIZIdOuMjGST2KLCiwr1NZEMQ+Qa+BwFvGGak8MYxY5MVIRpRFVpSyltMY8cpRB7
sb0z6BszD/XxnTvmJT+lxUqKlhtL/PE5l5smRU27cjGuA7EmWnlTt6E8/bQXhYci
AgH76hO2M0bzHMUXMplNylUjJG0Xd9/5orbgWBkgzaSiOxcSThouCF/q9vekNPLg
`protect END_PROTECTED
