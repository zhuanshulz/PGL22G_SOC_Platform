`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pl+hBs0NMLWG2agXiS8AlTQbQhwEQgyOWjao5U/hOuxfEhcGuN30VnhJFV6ujROJ
/bwRezgOflL3n5ICT91IsboUPc7hDHso0fEV58ksoV02c7Ry/4CHAkbnNlVjTLOR
TdHITwQQd3G4HcpXS3aPadg5tQ39iTL8fkRQAmtVxda5UJGRVEhHBgLNoNdFjhVK
2tkX/2ddlqHddnIg7S+5BRURf7WYYPOvfCo9kkM1y6K6qexujtDURReVYfJ8Io/M
X3+sCK3uYrph2VSKbEEE5P+uP90u3ug+DGnTu4nBEIJY/sXeekIm4aA+1ksVwuee
i4XDxbmFOkxYvdpxum30+dYFHLHgpsLrtNcEhhiU/VZ+dJBAkvUmhWGPLAX6zYNL
et84ra5VgneC0rM3Prx9dAbFZyOwJB143M0z2jo4dZbfnkGogTSk91QSyA6lSbUC
GfaiFc2wC0lJoTB9DsJpvhZJ/WRbNLqj5Hscm7OaW1W7AIUnVSBGUILcx6JOiWfq
brxRE8RGmwLrjG9as/g+FWu5yjZRbzc5LeeU3AYY0l3U2aW0vkwrTfbiPqmxrc5S
0b3LKUMVOhrFOWG1OYgiNVySqwy2z0LvhnhGddLxysWy5bPzRkik/0StWXcAgn3U
xmrvIC8IU1nUzpYjORd91OF00nmZZ5AvC5RduKZfjWSslAdIWQtKQC8MDjYpIU7S
Q4zYvdwDJ6D8eB59PZegTFpZSfEs8+BWhdOroDsFYEkB442f6dNz47qJpuVxBd7W
UxDoAkiDY4Si/YFgfaZPycGWAS16c31oQbpt9fiH7PbzF3CJUjn+AoBAWFwiCx+h
YCxp19daAoci5VvL9qikLH0YWo1vKTsDWu9pFbDwQRKSvcmOfxRPttY4sTQcz6WP
agZrldDfJNzXXo9o7CD+LWAd/FnvIFaPNcE3xaF6b9F8SVhH1oaV1SQutbbyl/50
+N8HtD773Fz4AgNotyikigoyejErK7pzMJMAA9H+F/K7M0N75AxKduVtPV901/SA
jRad5dunBuLevLW8RAypfkfxr4KDKN2S2YMwEkJMvULkunRnOKQH1bomxAcLuKtm
gGg/z6TnrWCIMzgXAnQttdotQm9vmBrCtI/eAEB/gsIq5mDf3O+x5ayV6ebU20ls
JcGfW2/LMJ3gDasJc+bksWKI60qF0Zrze5qCp0/z76yhZXqqwrDLyvwmpm4MVsEy
swCSLlgSP5vpQO7UwCWQVpeZ7uoImozVQp6gxG2vbMc8sk49MFyVDUkOEUQu9HRJ
mtrFqXbXNOo1rafzjZQDWijtjh5J3oVKyAx9iiKgvPQYezHEqQ993AR1hgIqFyTE
uibtjbzFdi+xpd0KGdACgnrG48SQukMB5MhHwQBrlrO1d297/pEbDIvn7BC4xPvc
FnyjqInRfftbBYho0SXvsiFityVrfxnXTbfzPD1RSVM6miJ1xFg6yJvezqAPRMz7
jxKRBG67aBlPsg1S7nznaXNFdJpHa+Qs3XsMaJKPY5LBMk1B/JmQhL2oUppmp3HI
aIwVf6evawCAJnuA7djjBdhTtNdEgn+nJ0sFfkQZnFLxdWKh10iodKfqYxcdodMt
8kOn7pbnjNg1Ze2IFrhumnkbfEYJLL/Eo48fVI4GmQKQSFszzTrOt+Wh64JMkNkr
B054puT/CJel6UxeiURLXhWqaCpRUoZlw45YqAiYAYjOU7UeJJWOpdUI7F1y42M2
56z67Nh8wFlvwIBpN/5iwxl4od832Wcxzj6FCZt+ZRj9jEgLAuKAHOTq/JdJjelD
LgtnN2C79GylUZw7ab63cE8YuZ4ma/RoZAa2NVTHlNve22TGPrBrbyN+smNIm0vb
3ggvK3W4n55VyF2L8Hx4pgBecXGOeNTEHuXbFFKNQMqADovlgj+icLDRqsxc3fIA
xOCkE0Zwz2RdzPec5mBN+5thUOAJowZlaLe3zRdQXmYDox8LmwRYj+trpgeyvkJ7
hsb2yYHMXBXJ+WVwU1WvbQ3ibSmOCv7c6z4DIPQMsz6rkD9qXqoTmEfAUaohLETV
OuFowQxtC1EaKvsgC08CGJjTWm5ZLq5FdretIBbScL69VF1ixidlkzrTkj8TTpus
V7SkOX8cJYyC2A5bnJt9FKPKh/BxnfEzhiriRn7ebjWUhaCsD3KJayS2slk+aB77
FdVSVpsMAIkZWekcm4AtVSlaJ2uiwvGBB3xfS6Gw1jTLAIe+Nkbek07ZvJ99v3wH
VPYgGE9o0LpKhruDNLgZrNdwTLe2H1OGfsE0me/Wm3vAzlVD2kQHvx620O4sW0LX
6344VoTWfERP6kaJXTKbtKMKK69/twF57IMXdk9spHKEx8orgSzlQosAcK352shR
KqLvq0IxwzPilKpBcCCXBA2l4S1A2jWg3bMJiKhxTDzSuGqppey2q22PGlMddK1p
EieDq9PKA0PGc8jbfTwwSi5xQ54TmC5x6X3RHQ47xYdU5PeWgqThQ8Fo9gBFT3qy
1Ivja8E/H5V3km11weVu/Yspmm5qnyjpHQTqdxOX7dVA6neWqx2Qvb2GuYJUK5JW
CbkRkmIqHgX7TsCoeHV2UxERPSir9wrlouLowlPakNgcqJBEUVaws6f6YyzCjiay
6iTaWD84hSGH7t792Spw9wF3LoNjCKEAIvwx73BFojKbqyRmYuINm/Sns5XVbmhh
V6j8J6wq7bb2uQ9arOOEniFuAXubNK96q77SJb1rNjU0xFlLbDaWtzWgjf2UHYUF
6lK+RmKRdYZT5brMlrqP90+1Fc8jsEISbtJgXQO3tb+xwh8sj0JFWr2Y5YUIHaMU
aZnuPJA6nxY7oxkpN4dRcV/FUYf5nS8QdJVHXpqE58EsBe6n8Kc8xAjbXA5FO+NR
SgR/nEOmAKD2nIV407pJkQeEXp4PWOgHdXH9croDAGHLSLkaCs6FX2IY8uR6ZwVa
pRabr8Q9+qnBsbbdiCi/icnNtOuetWIcFfY0sKuqXGk4QbaUsdeSjkHqHPOLg2Xc
CnRLlyqDk6Sq3LpgPSrJVH5rOwfUAznUW6Js4+mFZE3Ucavxa8WN5qkdp/+FAO6w
t6/JB8U7RPI79LCecuBcquUuJtlhedxrSlTj+fci05AV2p068IbBMjv1gFQIInrx
UBkw+T/RSevxbFpAeU2Llrqxtu1RVea+Jjf37VubbbtSWPVUTgKmRIfhApsrOsG0
`protect END_PROTECTED
