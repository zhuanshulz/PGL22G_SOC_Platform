`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6rPffVTzRMPXOIGehQLrmrCZzRm1kAEKeYYahVkbCLt4FDbNb/aPlHUngoSdJ73Z
HCpqzdHujyJm4It8IKUsL8KqpTar6o6T9B334viBNYCUX9Pv4dwgKOQ/z3DcRUOm
2/+icu00BMID2SpZ5x3bwCq2gz/Cx/BH/bKf90oEM6GLBXVr41d20E9i1PWEqymc
mWF6cjn/TnxHbHPmurYYMuvq0I+1GRyKV+PcDS+kQzGaqDNxfDmXO2pM6qsHtYX2
BxUr2pd6xJOGxqPTFQCZ4QY0/a8iSPjvxLCvYNn9aShGBKgeOqzjlPpferJ4rpIR
XGR16zyn4b1FZEPTDfkJyi2BTXwEOx3g2BALJUVHNTLBZJrienq/HuRXyCQoVqbD
+C3AnUk3DOmfraytnNGQN4W/Evhg5d7HBdIb3UHIh3zpecq+iN57Sl25nXWpq3nb
xwOfamUBalIBCm1chv7+8X64C/zgy83DCtt3xQ6RrTN1wDXYmlCd2SgzLU9EenOa
EfsrZuFlHR61lf0uElOPIfMHYi/E9eKYI8ZR79E/nDNcx/B1aWuiGynypovO3WkT
FQ7vCpzZH9caItwN7KtW9Sq299mlWk0wFy/3nr5GkBOn16ncKxxbjfvoxX2O1z8T
QeikoyloxLVmkkIlUiy0KACG554cJDd7pRxRzqGnjcyWn4fsniSxa2t8WgGLSPtt
Ts8TffqfRbI5bMLSIPsJTIbb40UCwH6C61FVqeiyu+yL4ve7Fg/08nR/59cN0Ejw
4e/Rsx1dIIDT8piy/5WsRpFXLBl0Skq1HCNLLL2JGJLnhPcHNRlhmnR2uoAmPmb6
iyd7LWAZ2OPPspfm9qDEpFRIyzpe+2/3Nie+y4bxF197Hx2N5rZ1EN0gs/H63YBs
wYxAeJeP5h4IXFAs8lnPELEjooxUY6MSNnMdfr+fCEWPD8apEO7aMVg5NWpcW04y
cnOKrSYXCOjnYY2XvW/OVLgBtxFkEzJn/aR4Gncy/9kRd25AtuluTypRJ5BiuNxR
c37q8wO9e7+XRgJZStYMczcvvbv0eRwRi+vmcR54bFl2j44ksH+td+MqtDcVOzQP
dNM3LMbG+jfZO4qgp8KZHRqyCUbvo1v6kttPTwnEdJeYMXJZM+7A7mGC61i3nwHa
yR/3MSEyyKe8Ks5CoEjtK9fZxCuNLkzkYfNgZo3Jw4N7Rx0nN1uDwL/fDxGF0z8z
cFKxJJu54cVeJLoGyogP3WlByFlQuJFHDNggPqyuzWOYEwAvM2oV67J/QpeT6Xt1
K7I5ocI9ecWzn1xPcmkMNth6kbMaBNNgcOXCCT70d40KSilQOC5WxGaU1UluYWjK
zNrVyxkbSCIAi26oo9c2ykQGnuWFKkSjyOeP9fQBietrzv4IkRavbfvM7M7ND6Iq
PAfpCYZuba/arfW0DTm+1jT8yVuk5u48dwYohHThPdxM6Ywqnx5tdtxaV0qr+lch
InhfvOs5dIBuKJnHgX890WQwOwxldKb+2FNTWF/vToIgxLfe/yvsJ4CLeW12jhlo
KQq1n0cW39CAOsSFcSkcHgKr0udgrV5p0ri008JZ+xISCZQMxqQOXFhw9Y3V+zRc
YyPvFp0OleK/3ZUn1CjwtZZRszdAOGXXDMSvPnMgjTzYfpTpxqugQle5CmM2V/5R
vmxM4uap9WkIvJ42+2Nw/Q==
`protect END_PROTECTED
