`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rlz80M+O657kWTqU7o4Dqp8QD4zaCFDVR3rpsznZ4yQlczh3nhrgPUQwPDgyrAti
s1zUzrHIxmA1iJfUWzHrk1y362QHCBnHj+ixcnEH9iNiXOfFpWDT7Vq2XtLAsxTf
kvx9oWqm6qSPCjhAJDP7Mnr5pvSD9pD6LpkIu8zHJ9ASrYvns7TM1YVG0WxMktAD
RZxkzncdJiYxZPTc6YsoYIb79L6CKik57WFH74VkS4NeXp4p0YkEQ85UEo+RBWcF
QYbq4sTFVnYPRk+br/INH6ddbrnYYo9CpVLwcmvdCVUlPY01tIpEMC0oOjgc2V6e
UP952jAgQXWNUFu3rZIUOb9z6UuRxUlPWyyaAtKmXFjMY2mDfulu/JJOT8J2QCYJ
g+Tkwp6AB69/ssQrMAbqfs0HRh/m4aBSVAuhZymlqSGDvM13DuwcHPBi+x0RT6Uc
IBpFxXrIPRYQ8kUQ24fTVPqRVbk9cwpNregAhfsDVABF3tlUA38yDsF9lgwPdh03
OzT1U4cNlAxcRkkRa1l9e3nZoxLW+wnGV8R0wF8FayRsmBRabwDmiqIkKHR5QpRB
OnmeoHTt7+L+VB2tJ4b2seZweAzenBT4gJ44QrfgyBw6fOkZQjBIorKB61XFmzi2
4VZMI/yCL0SMET/9YHZEiCurgDUgIIRo900hiY0Fpq0Ayq+zgtIPtpWwrr6vLKgP
I+JNb0wJlLxK/Yr+dkyEjwwQ6Rw2RjDrnrvQYsrG0Hr16tsqC68ylBdeRxRHgjQ7
nr+tmGkjSrnff7PzVskqsbFqbfVUTzdMSbiQVnSOuADF+rbvRLj6aKgxUqIkJkOE
yKhEnB/NLJaRXj3M2p+ZA+8ukXWcu45MtSsU2mZNiSWeTE6/ZExQzzQX20EkFdHz
2j5dNFSTxVW49M28ixT3yPXGeYeAnvSvQethaJ9n5ajEs67cKKx90DQoPzvhBUwL
yKrkANe3f6TwHkj4qZdomG93Ys1qvStqbHr8BzNCKOo5lfelQ/Ete1P5Wu6yoFbl
nPY479dZgvdytXfs7f09Ym7Dx//CBuLF87e47yGB2s4vO6IZQxFo5YBPLPRuL0wo
ha8OH3PB736rcrB7cdoahc71/Qoq7Kl8agsp4MPApBLgtDuo0u1ON/uuRojsRZps
q7yq4QEexYjtBfT4GXf7ikU3QewA52Z5Y8mUO6AWE+bjcD0WAnD+spz8B/DThMUr
nQk0yiWxNWg20yNGNgUpx/kl78F4X8Gsq3c0jS13+t86p04Xw81LLdpYeiwB1ZjA
jsBaNmhvCFiVAA721Bg9XqCPf3RWdhvHLNg6uAgadlrZxJP7z15FuzT3rSTZa/in
YfgNyOVjlg/1tZfm6w/58dhosNqSd4yPI8nKbr7nsfa8HW1j8Pc/UERTX6RhisI3
tk0Grn3ovkSXV26J50UqprKW3Mc7dO0NZEx6hu4dTRzRufIm5ZclRmkVq33nxWHT
ID1wu04J3p0Nx3Wv9y+0mHI7+8v95eZ9iF72BSNRozPejyfmWzWJd9PZQv0sO57g
QNcqR5Icnw8zSQLW67yI0ip3IniSAJ9X8rs7xRIiJmrQIhDcYvEiYKZrAyZwhcUq
2FH3getP1XICA6hoi4ke2/0BA/QpSFk1f2eO0fih0VIWQn0Fc52yGD9C0XL5hXk/
vGV2Chy2F7oo89vRKwEuYnCQRafnjnZjAHY8G6uHb9u8Wla0zLx+QHCg/gbVbNhS
oI0LJBfCE8JDty7rByIhbxynU4qDIR/YQ9PgwbTTWdfQD08VkGSNJog264x80oU5
3gQhV/fFSx9VHb82ii9Mvi53/0+Aw1BpnNRR+8w5kXH61HslD4Emso0mXXUdyn8P
+8DD1Skz+yQq5b1jLm4O65ZVAXS78zTEWAClIE9Qto7mOzPJFqcaQ1VLAWOUS+z7
tLupaKpezXI6G2pdN53vB11P3n+KEMdtyG0yPAXbzfeMrnfaohw4KRRrDK2GhlZ7
AKb5QIk6MEJ6VxcpFA56CtCrFnqy67BkMBywuaKl7ATIF9TfEGDBgG0A6sUP3jOo
RAFV7y4bSZdfnh5rBkzCXJSxK1g8RByD2m7GpVAdBuU2oMm/snSZqXkbGxHHJS2A
OYFCNnhPIEQ52oT2n5Z59hGey3BkTj36e4TkpqsptPrKL70nIS+ghBQjb2rUjaey
syqJ1yOdN0TJn7imOckzLorQB5Rbr0QR/+s1M9l/QzWbttlTZ4wzXOFq5N4Kiomo
rZZtp+NwcpturKmI4zuXVp2pp8LDGaasWY/Y3Ohr2QpykrcJqV/J6DIupJfLYJ59
EBAoXim7qX+g/+RhZZRt4pN0m70HsjWBOebBhlLLXsq1wuxfXt7dKJWkzgF4G1+c
3gMlgpYBHPkYV2vTzlA6MG84NvquMHfzfOvR6Dunm4VVUORL5cB51f1rjHddfNup
za47gqIDL7Fbfug05knrSEWic3t9/rXw9BCoiVrZ06Y+Zyo9Z7p+AXzpFthAO5mP
L0wMh056xQ9UmuTRuJcqpO1IWcHb0qD+sYcq9oBXTPqprEdBblUFyTV97AnUHBBp
Oxy9p6Bb3pbgU5w++yNaAPijxL6eEJD2tIA3ffDDKXYKuI34gueGjxR8RQa/k/gQ
5cHIho8ndtWyQj6L0XeK8LIz68/wBsNjOWj/SCljqJM18SoPCZp8Z05hC616F7Ps
a9givWwWRKkPsdw4K6LyC1EyoGQmALG8r5WbL5jD7l4csHBnQCYn3Fcy7Q2Sa0Ph
/26duPt1u6qTxA5UK3K/3upjl9aBIn2tldkOcc877CiP0ezDplyjXw1jnOm8VVEG
YuPA05DW3+qKKXrVNyJ/rQ1QE9iNES+Y/eo1N9ZuZBh4L/l2vHBJj5QEf2Pxr01N
ChDnvTRRiRhrSSPzLT0lGh0dA//MfikVaXEArbtf7tleNmSWHVxgt9n6TegXrVJc
eRA+GkYZDC5P05ys2iXjBAjH3yNamcbpMqVj9MYBRr19C+R1B5J9jWm3B+woDU3E
Y9bUGac6zhlha5QjJTLWSctDRvaZt8mnYimGM+wLRmqIusgK4lfbz3AmjM3Kzd5B
8gxfGKdENRgculo6PT2PQCbikahkIGpbL9IMn/mIUD1CPr/cmiHvXSo23SUcccmW
d0p9YKyztRA2JmRYvpsYnTzd8XInS2Lt/AoW9T/02I21V+SaFZdKS5TzuhuyeKpD
yNxq32mWbtI9hA92YbVyzgsoZ8EUczy9C/dRsfBHSmpVVvtm03s54zqF+gr22J4f
GkPLweiEGoJKybSR8z9jp5QePNlBMKXdwIewAegmkBJFi0zciEwhm5zGEf8TXrBD
PGPdLva5sjs3Rlh4SNQJMmtNKJehpMQgkBUQfcRwgZDX13bPZXDnJitNOcaZcox+
nqOzbAoRqQZoX3YYwGaoX2s7/5D+Fiy8jv9Kd8LVKKKvj2i2bBE7mhugvMS2EEpE
V93Zoy5+eN2IbV8n9Yn284uyp+wyHVA8Oaum9F65k0QN0qO2rQQ3sP6YHBsC4u+p
0jh+0P7QwZ/q9hQgSvyBYPuIy+wsv+7qk/zlcL2G4XlFHo4vndgkvK+JjhscwoDU
xuJOMLOxZd8XSCdrMWoxPzfzZfxk13wTGI9WCsTNd+Z8DTYGpRk4EBOr4un23W5K
yHSTT+Hv+SxkhvSK89WiM9Y6yNOleaph6J2u0Qnj6gSu7zXLNarbG3zdqrIAohof
GykT+61FegkdrQazFf7ee+oQcunzBPoDqatGgxN30QIxT83PSz9huY/Tj8N43AJ+
`protect END_PROTECTED
