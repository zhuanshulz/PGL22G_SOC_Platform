`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gqvs6QRCc0TMmuFhCrfa0tQKNxc6qyiVvMUIveD/UmswgmJHeAROhj5baFNPXKze
HoFVaZLZSfrJrIdI/DSC53Uvu7fYtEnpwaNZ/OX9ngBBW5hXd/ZtyIU89oaWP9h0
4rUC4DfbEhPSXP2d8YeDgApfyaBlK+lkDhwA+zwqKr/Scm3UAa/B7aU2vZfYSI18
bArAGrA7Vbv9bBne6Q5Iv6Z6KQzkcjmDVE5ITxkKGJQrPaqQhwtkE9LUYVtaT5Dc
bUzD7RZpvP7AHnhS9kr1mG5n4+sleOGNEUAh0xQHwyW3kB6nm/BD63vZoR0TDzDr
R+ftxydRs9wgmFk4N/G1ztcAEJJLYcMyWBb4g7uJEkMKs7t1FNM4w1RkvocuEYhc
0sQiPxHlOSWtghWLHPx5iwxXe3yusHiSbjTrG7gUiJzxGhjoAQMB2TUKLbgGyBOx
udkS8BF1jRm8lzQvi83IPtRSDeLusi6jtKgf62JiyNoyKBAfWFZDNBkHubGTFNyS
MqdGWx3M+EsNqPwhkpKBqYP6mRHkM0n2ccrSDgBA5/OSpwI/Uvzk58m0ZH3w2Gt/
+zn7T8EyCIyQ5fXDZd0gC8RPoA5cVAuvBUaVU2BvzInKW5wMxf/Z3GGCIHt8skWD
3WOL+obY0YseGtRg1UXooJLJG+OlImJT0huXty3mDhZKVXKmNkGbazMcIEouyK6R
PdMLNnuDb0bkHI3Q3Ln6+wIpt0DHoKZ4uJl4d2SyfHSVBU/NYQqN4SLRL2EJ2Gal
Fsmuel08DYoGdowaRlsnwB7d9DonaSi/e8u8zPrtSOyMT+LLD6wp7Nsaz1Fo34hZ
k8EUINCD+cq5AQa/7mspgt0BRT2vL0juVlcCHP5YftknQnXPFEVzCoNW3mBgyh/f
w47E2vEbTs9uXCAa5Suf3SC/30XExyA0RGuWCMH2nP2tpC1yx+bxA4NC42H1ISV0
mLQ15r7LenCiPMe1rQ9pufhUl/Fk0mqluqgT5pWRvH1yGXjg/B8Dx2k86yBnVfiD
tiXr6T/CADZZCgnOiQgMZxX+hO6pOQ0L4OO1ufApnDfPk9ljzKyATIXErZW0X0mi
QRbuS46I64xXs97FQmIn3w1T8rSeOdSetUj3fA6FS9k+GTvlbRH3wzCxnlA2P30u
e9Abl+RGWIY33k3f+WjgYeLBjMRJS1QHq7qNbpqUl5qAE0B157JW89mRIVKh8ztu
CJvOXxhCPxsJH5drpJP6y2Tm5jx1HsSmUcnfYyrBdeQHrhTQmCBEYbj2U9rzl3a3
CZQWImWOS/OIgkO7ttgBpOH78xlxEqsAq41adEnQGXeSb5n+UgLVEHgUuwgvikcD
vqsm1Vvse64V8DAVuuCx6oswzb7MIvam0ERLXHUOTd6zcEQpXVUCiRKhgHGlRkzm
B6yz/FDdhnQTN3mFFMxQzeEw0pOAbfTs2bcXcMZsZoIDr1meGgTo0ntRyb1nYfkW
UFn2ZJ8Wn3HzBkdm2IhndtlyttCsHdjFswbKk5RtHhhYzqcKjFoo7dbQceDQUn6+
EgAQb8mmSAHA1+ODzKW85t4vuDvA1snWRj+nVazjQWB1AhyOtD2NXe5/SEoOFFnh
uSHaYdlDT6FVR0OHpa3gCh2ZoGf8IfbcFP7ZLDg/Aac0IlihTUVy6tQ1tiQceYGf
PIxhgYXVoqNRXq37N+nQD/VUJdTk2VDtIrtXSclWfuuwAJ/iafkMkgyYnXgmgWDh
K+bsL5RorHzG2MLTuXpD+cR4nNPeWPvf7l6aXMwr6rp6JK5HYWjVZlFrWxyZib4v
W08ZTFyiCol0c/vsFodxzsTnPL4pTqCPhKHrVjEPxXU5PomkwSesxKHMfcU4vmVS
js1mITvS6M1jED24eCNBatT9ZwjPu2F7MzGXRlTCsZdfnJKznUBkolemEGUJCSLS
dUuNLonjF/TtYnPRIQQK9A4gYUg6kor+2MVYo9VcxwYgaxAQpUgpgfScc8D0aAWx
LmihYiGGS0N9fKflMW0Of/JU6ldC63jpC+IRVZhU908y0XgUEvyvKckHG93DTiHQ
NAizZKinX17+hO+n9HDl9ipR+exUvKc7AbK5sgio4CVkj0dKUQ5LniP3oGiZG/pq
z+IzZJNMmHVFUCJs/9aS1NWLu0U4dVWhfmzjsKUNtVMk19yewVSJMgzHCeYzuIm0
sVuMZykC/Twn/PyGlCfbYOzSu9GBawujZQDgtMZLOUCseal3tEsV/gMuyVxBEkzB
wbuiOmTt7U6DH1fGZ7N/pTuV+jp6WQU416bnRhMirSIlARVik9Vx/LhE2kLQzgTr
uzJ00bLJkPIVDYzXrsk3GHfpeq+IRqRRQh+Q96gJGKZ/FLN9dzJzaZrIj++iQxqm
rQ8zmPqQLzg2Sfcp1OChuM3S/KJgTiT1Zg75lIksHhzNsW6kextqL41n/ETcdqwW
vmYQLQ3zcx1+oeMwQN269zgfAOwV66a41O0V2ETseeUO6lCz43cxpnOfJ/xNA9Pp
q3rSWL+pyAzbjP0GIYjjES0XY+9w102EynYdMbgFBzqdR8NwCTHWK2+h/0Tn4I6F
nZdAZs/W1RxYLiw8Ux4PGPCSPoRIgFtliydEo5y6XZ2/oEBdB/u5uyPlIx2Eh+ra
ieITOuPmcdNc230kk2D55JXkxNQJtrdzVd5xFuIog8SY2Mud/V9YDlNB/RTD/lbp
PwkPXO4Ipjf5pJrvQibn2yZgy+rvDdNQCXFWJ+SBej6HBPZHuafM4VjeWkYmhJNy
CXx4XSaYWT04dOl06J55JdchSI13hVnA2C34SiObedJMDRvcqpjYuSj1ZbYDudC+
2DLxr5ygx7Hy+UY7YBpWaTmoZVdYMRA9TAHrD/L5q373tVQTJy1+Il7TFPbXh4wz
LB5WCtKKOlLfdBPEiGknA5reea+KOxRSNf7fMhdt+LEoobqlRUya/+x7W5aPe0eB
PrMB+I/2Fv5SdhzJUexB80EdroyfRglj2ySJPHwTxd2j6WrZX4DxAtbTR9J+iiVD
ubiBc/uUsmu+7CB+K//x3VK+zar37uJh6xRpGVX+6mWmI3z/mZDSu9VWvcLqXeHT
X9ZsCLdpAgfln98JBw4couONzNfsTwgCFAXpZ++Y00z7g8HTbezxgjcwO/8Ei5uk
u/xxdcNOazIBZEiAIazz/HlTKxHnAKTis3CmTrf962sm7jGXNxOQBdkfHqjsVxAj
g2bt7m2r/C7ni3a4T0M5CPeveE6l43zrFDRdEimgpp3SwrDmy+sThbFHF+CmzrxV
1kKkSmvqIsDtzRP2QW/VxsSqvZdqp1cton8xVpk+NkxGZ/Dik3hIDmMYamzgYD2S
f5weevjLdcQXsLb3syF4iucfdXFcsHVxKKcVs2bT6Z3rTq86vw6vF50bzPcHFe/N
oZP7ujvoTxFCo9bt63sQLae+102xiRL6tjzBN+Vi3ZyEtNqAUueGHveHKoJaS8Lb
j2jP3c9KyvTJrG+dKK2iqpOOIYIV7W/HqEYlPxAHI4rv3fJIV6slS8t/UkwDRDeU
9+zN/cIpD8CPUU/ZtuDyZ1BsWhm6zc98pbqL+HmyNQPu32b/0oQ4LT6BmGVgSHHG
C7YXFIGPW7OONLCSst+MDf7BnBGACKTJFTqCf8923A4g6dvKY8CL3rUW/8XLCQ4n
fcyGA/DglXVeLd/5XP7AnIo/vDJSA2l1ORD9Z20GCM+mQV4MRI4MmoVFbhWzEApw
eVO8Mp8JEIRVTrBg5JeeA4zelCTnt6TNRXio+HAEJxwIWjBhuWTgj6SlSaXvID9J
JTZJLnPOm0+uBLWxkj3gQISagVySb/dMjAssAsU1/GG8Ea2/1qPf1/mgmLBppMz6
NDIY2pBQql3ZIdK68MWhpMPbRN0QXNKcuTZNLgXDjFnbXLCDrsUlT/1c7F/Qvi67
5LJrVgPgQlZmugzdph3sY5kOF4NIQyGQlXXspQ0/7+Q9RCkkpD1ZxPKIU5PEftVg
sL04XSy2X0BzgXb2AApS5raF/8vDDpPbksZZY8MEa13o39F3odFH+i2BVBVOLerP
QQH6xjlQNpETKbqqOSzqSO6VZ43wlOnSPec7DDm+RZgBrX3087m4uS1HZhIr4tez
Zf4+xEYHcZ16yqsK58+tqFjVaQ759Ch3BfsdG63ju1n/AZ2N5llg819wEOVX0LXq
6ZvWZqfzM8+ml/M7pVZ9P4sghTv2AaGRME2BVBzEFJkbbotGoB5qNrZ0G5YmctX1
hhww5r+z7KgOuJAJdaIBuNtU8y7W5cf88vO7R3qcHAAge6WA72UVUUQtyfrp5Qqn
CCsubUz+uuaI6OHC+vx/XuFjMPh1JiTXVzhu5dxzWl6QlnIZMQdaleTQuQldCpbv
rkKgcSV8WJadzuDmfKL13d17nWYuXIDgtbGgulbbUOSpqExAZO04fIgGHE/BtKVJ
3urlKr/AFmF+7M3BiTtM0FJrYjcLgo9bdaCu7vN4zT+BECzCUDYmSpWY+AwqH2Ul
5V19Q5rx/e/1E6DVu3KlmEnIl/mkXV8csV2RoQ8FynH9RnPgwfckOchuXgDBfQDc
JoBd3THUax1eswOFWyiB1p3tFgl29vkzNE4JqgvD3Kr5TEztT4bCuAYswASn/MNl
A39jsrHQxhvM1F1NKTZoUplNq3ArRQoLUpgFBgQIa6IKxidw9xcSf1gf+AR44ngx
miw/VftCtMfoJ73+3pu6BwzMI4Ls6VRe+WVdvE4/gKIQc51s3REwTyGy7wbWNv5S
X+OG6uq5x/dLH8ic7JCcAwwbf/1X6FTnQ6GrAKWHhQeqAQFfHu5zF0b2+CTa8w2D
PwZSOAvEVNlJUZPC97AcIbPRfP3PQm/W/nqp94+lo8rJ1vLfBT0dEamWy+JWExPr
CGjaXgRA/KbEDQdMLiybubGY962GKPoS1R8JgeMF7QpNAj1ztOuiQx4n72PijsEt
eXDRyAQwuX16ipIVsoKnkVMffHR0IsPraZkz0baZN9h2BYVgVEiEtGFPVpRxEm+D
JmVm1buurK3bsh2Q8JOIuQ9h7DzffTWgsmTKMQ/ZO15vy6y8vmaW/2l+lIndHtOB
PI+PiEsbhS354spug7LludG2UtEvB+l95CCEN8NIOOCSVkQ4TCLWiPOuvRx/R4v0
gTHpAXh2tp/Mk1QZt7as0MIiwnhqf9dPE+8KNp3jn4tboV4HR88DAZCy1EL6VyUO
LmjNqVxzY9xQ2ne2WacLZFaXI+D85OXyIBLU0SHffumMN72C23T4BOad9UzRS/E0
zVX7y1HWCXK00WTFiHHr86OH9O32BbZmRQD+U9B87k3NNzv3NZ/cm2GO0cqhgSOY
KhVsnIV4hOBcOt1+FVtxbf5prU9S38nmtRYpEBsemhOk3npxUwdU32AdhCRH4jtf
B4TCea+TenyKICSyuN87KuJ8G0+4ciIrdgYPanA3Ye94LRgr2mvtHegw/29FJa+n
r1bTaw8MjDezwEhnxf6bSiJUAeCfRtQfWD/fymNRWu61Nsrvibbr9EBW1OSQ9mPd
fzxER9Pp5sPOnRcuY3VTCA==
`protect END_PROTECTED
