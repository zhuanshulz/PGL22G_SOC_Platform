`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ejuRkNiWoa4hyPuMBzRXciQF4Fo1Xjv1hxahCQ3njDRnzDriqYdlukGzmfY9YZ11
kDlJiwM5xQN80SFSDl3fjTa6UPGfphPIsDQkbd+7ZWM5/Vb4fWt/FP/eaCKsIyII
qzZW/GH4yl4lWTwud6jlHs0ql5+7zAkG50mjA4cVZxoW45f5coVtUfEs+Um7kAqu
H6Y1rsDDutiJcFGJjg45ZeuG92aQW6Mpv7/eYlAHasNJGm7bkN49JTJ7QqkjC+oX
YE/F5yfnKvAYwg7Y+U1A7/i5hGEgwC7nk3ieQFrbvhDvwIIV0OsWD/5XrwW128qi
gx20rZ/h0aqxT8KwNjkzcdSug8R8FXM6ERoSmQnytFyxrK9MVAiuVlESEgJiPHrj
SGSPGDcocU/d/kFpWX1nCjNSUBNQB9HJ+82oDsFDa97/acCnLnkSGOxlrqTBLfC9
T+GEY1Ey4AV9mgV9lDohwzTtVe1vHakA16RzA7ihneq7AES58C1FASRukt0Tlps3
kBbA6bG/itdSd10HQned01ZS6jmk1W8l/pV8NsN1c0z2y97h1UjvbPgcVebnw7Of
FSj6HvSDUZrFVwVYnQ6QOMaCWHLBbe/Am56n5CcYXHs=
`protect END_PROTECTED
