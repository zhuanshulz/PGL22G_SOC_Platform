`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kmweCMZTVA0xGuT4KHu9zCuWhVyxzqBWWPKq2aO+uOlrbz4S8R5BwyXgomCIdlzj
BKgaRqZuoFpA5sQuFBh1ouWZcDlyM7K80lB98/UXEZS6zWcfUG9kKtTNqdHZZ6ip
DIAYPS6pntNQL22SQCI+04VE7EgZ7jEGRcdvDjCAOkDGXO7KDMl8DPYesPcET660
uJN8Mpd7qNtIXst3fDy4BlCXjQT3oy90IPYhussfG83l27D9vWwxHTYefhWWK0Ar
DFr04fGQU9WNr/IsIt7K2GaoWGC8O4SnBYXOMs3escZ0MyrzX1jf28yUekDXUIYS
8SI/BB6aHx+9H5okPsP09ybfnWypTa8QyGErTHq8CxftUHgc5KyQYVYPqW6wHBKp
nw+a0E3AyAjTPyPeuMRKsAdw7gY8ScTFl/5BUsRYXatogZAEr95g93vEuGEgGObv
4QZ2AefbUjPXbVhS6fDZ+ohgQC4T7iu/wp6wS1RUt/hNxD/oX+3d9jl0nBVsHMoP
uZd7IjM3fRcdtyNVa80uzE1NFCb2SQEBD89YUexOxe//WKc/JJa6LZDMWT/Ik/ao
VB6s7Ocz20h9pwdn/LGRegyGNbk2QwRQBH2CAiiR9PY8EUsXFpqekRMwD/yOxh0O
Vd2s9sUt0SgvrO9Mnws5HT3ZUxqlCQo2BVFz4qE/0D4=
`protect END_PROTECTED
