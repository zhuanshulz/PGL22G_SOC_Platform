`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HFC8OY2sybVOGfR7UMI4a/pt9aPU/oGSSiS14uBBaz6gMi41os+iOi2/enAgmjuK
x9brvqLyQtA8imqcPjHuyBz5eDDBCXcCXEPfEBd06oDkI+0uew4+bP5hUXisYs4G
+jgeftvLPiWlIDL3TMnpvHbsEKuXVWE1HgEdiAnAcUrST9y2n30uSPLVFNjIfOEL
w/bzFwxRF2uxqUI8ufnqR5Eot2H2A3obw6xUrgNuoAECVscXJUEjdegwu//jxbf3
pZOe/OHtm3osWY0WLXJ9dFBBmBzxghIARztD3DX0tZ+FH18v6DFWZswbaQFfij0u
wh7tMWrqKLmkzUK0v09t3KtLwfBx9NptKGg8+OAID6MsJtmCnaGzDDtKogqeWqa6
kmtDA624Mc1D4e5TnaATGAz4tsux7wQHyjlvvHzMwkc=
`protect END_PROTECTED
