`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3pPF49I1tCthtibNL6ZfvYek7JsY88PrGaZneAFEkl4KqJla2p0lwufPBZjwCAG7
9zCJF/y/HuvBAEh0q50xHhp9VCKq4VXbXeHwDLjreAkOE0Gtt21V1sXAmm74+17a
RLhtU3R0161I0Mq2L7VIVNzaP49PcbD2Lw9OW5bLMgqUvBJMpcq38YaNmcwDM/8J
fSxTgn0z9MoipY0XOxU63M6A6/w2NY58SHVkOEdE90tw9cEWEoF+vB+QAiGzo68c
DUvWwiccMJqbNrjJ4Zut69eMMGhzlGA/8cSWVZjbPsJm+8bBDLwRdDrB9vWgdW57
C5GldRemPtwNFH+V9TcUaufqX4quxWpB4w+16g62npMov7CcIIpFLcEtFjgLxvsq
DQbVKmBqleoCI7SKYv6CEQNqKnyFxMIU3dSf11S6WIauIE25UhFcZabNsEvh3ebw
11jdoRm93erv2gjt43vu0jows8SHTg49OrNDtdqMP8ZDhtIn97zonrGLc3Ad4Z8f
PODU+303nO426Pq+aELSsVgTty783uCal+YqHyvC16vMWe+zLFVF3uIhlIj12j1S
`protect END_PROTECTED
