`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LPHVF4cF6TR2ELxnPh41I0hmlycgc/Yeht7YgvkJ+FeG25czkC4Y1yYGD4XryXg7
dIbocth3LRjMz843+ZpPRrVv0Msk0sVY0q+whM9jE3aURrDYpS68PKZOZtvpOwhO
975W7cfJvDZFcqlKQi/BORYzVBxB14N8SqcySuvpzBKVuu57NCa404n2C+WfUCi2
cZqYXOOHCWzNVa9Fyk+NvKVs6sVcV9s4+p1KyIhEG6VNoxgDJa6iwUsDGIfmqzSO
NnLB5wjqyU7Z/vvBxdQV+rWt0MP1DMkBp6/1VwHf/vRSZC/hKZk9EQzjfeIBNeQ3
yx0Vze3L6q2WEA8xZK556NHromX/3wUKxyVosplbPBKD3QxU4DYAmfSw8VYP6qLD
IOaUekq6DI11MERY2DdY1iDgSowGdSbCOou09+yBvRxLgQaddGe2ZrkkCqHESR7q
gOoBI0zqeqOWGdD6bvGtjpk9mVjK4ooeoUh9JuPdoxWUid1dOudejvz3gJSliKyU
orH9TZg/v5Mwx0CRiZ+eOJIHav/zyKki1qrJKjDtmrEL2m7/ZxKyLbB0WZMESsES
gip2hNrrI92cypx20+6kpGKUudbUtgTM3uO7qPxjUwUWTDCuYSaRd6goIdtuA6Dk
oSOIKr5vRXnMBUCo8VXW4ZAF4FLD9zXdFkV9H5qNAeW2i0+m7NQXG6EJD160um/b
/dI1FpmNWDA18FjhabGjx5SerB6wfxbZTgdronkp+zXUmkrdLBkiZ5EqkT2iJuYw
JqlXX4RfZYDLKH7WyiQATR9JsdLi5kjFa9IUBAkKT1S+XbxQ/nnj3tWmFjuioWqk
dETzkk4RRv9j75rQVewb4Ty5f7zjjm1EL0V2k6tfnunVUwwFNsXzfV62rOMEh40U
OT6E3XMzqpQLw1AYVDO5M3pjkgdwKS0bDv+qar12rnvhcF+ODXKBi8idrWHOw7O7
MjPrv9LOUv74Wbld1vPUbZrxXTlgQG4HJ6/HRKmVikaNQ6O0PToJfx7EZLnnCCLv
K4P/rG/AgT4InJo12ybcnWGcJHLTm+E+4ZU7Aco+5woSz/YWKEm9PzzyOfAmICt/
AyEi3F/mt+3/8BQXK05vUEiDo1hJqlClc4UwU3dfNpX+mF5xAJeEsRa5RqglRAyV
W4OGSxrgOkJXdFCWI1uGnKlS8xmx8ze1m18WVPQu8Y7DlxloNOi01sSdgrYaM9fa
sg3TgCv0142mY9AY8iqQYQ==
`protect END_PROTECTED
