`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0U2M7QCZm8AIQ5kYff025R4TRvP+qLQNHq0ReKOiBLNs0fdU9+vvQiiRxbIiACmA
7ILm6khgSuCkmpk+2KWFvdxIgcLiQycOHvCHGgv6Y2qyUkCgD91WK8YFEuSZGCyN
61hZCg6LBUvSLjElQYlFwPVCcnVMReGoZfvleLAd/1Q8jb9yKB6AZFXs+Bs1K3A6
T01N5QYIHyUr/qfd2HSHnfV5aZjIn/j8I/zxJs5H1b0Mx8Z7dzQXgHygSIHQCrsx
33IWz97bDNNVmpn9LdBVk0L0xLgXjbaOKqZTbIrIb1gatNssa36FY4AA8Fepynab
9QfLu4LBM9hHid6dSJaut89zF3p+AOoupVwrCjL+/9JkpbxzXBLWjh/ujXJlQJeh
kfXyy67YGDHhjR4mNLy0o45ZGlzM6moIw78nIXudr/g=
`protect END_PROTECTED
