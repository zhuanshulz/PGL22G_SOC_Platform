`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d/GzfRLdUhq53DL9PZTmw9Hpr4kp5SjaMDvMG02F/z5Z0s5ZKISSaUBJW2fQ1tOi
3+zjphQHYUiHhhhCs5LjkaowhRnj0TY+0dLuWofkxg07y2SD00lWS1zAHe21Lrw0
Svy0mAItdMAmzSyGLegq1o4DuCIJ9FE0IEVrvutzBqaxB/jRe56q+6rWRpO2V+Wm
dohBgltlkF1X/IHfhADY3UA3bdm7vMISh9tBjAnCf4gNfjrMTjQf6KfFKr2AmQod
cvXyVgMw8CH02/expHFylJQflZ+8kO6IUdTXxL5SaH2Yb0Rk88sCtjamUY0X6dKw
TpypfK7vgysyUf23wY9qbCFVQ6ft8PV9wrGlgezJQs3StiQyvdzM3XCqd9EC2X8x
qU6j4RrETyh5MRbBmpzt5y9DVr2v5HApjcgjR7qLW1flkDqX5tDr2H4tAreIaBBn
sl/WmfczFaVL1v4SWSLcQfXK2zYqQ8uOr0anJGAQJjCRORtyg55VRayzQZ7pKw7m
n1stni58kA29xSeH4WPYrn6+WffMUU84Ab702jMoK6BWEIQfoA2jzGJp2N+NaQwQ
pPeJnwlzMlCQFQcUi9NlaAqDGCKM9dxR1Q6jqChTVX4QLFBSpF69cs9cjzHJwgLx
pdrTucVkHJqhJ6EQbkaGwvOg8s1q2hwau2asOxpUGMN+DjKsRnwBheU0fG+gvvCc
dKxaEa3dXTXWI7hlM8Rh85Ls5keB/eVzMjA3Oi5yPT7m2P3PxrVH9dc2HHWIhi3a
gPk70TkT2MB9lOl1SdHzvadj9fYy+P0jigWiFfUKWW7dtISQYE9T4hKh1D+1RmV2
8ahowOMCME/2cd7JJ7wKzNZAYeSSQigXIdEO99hE05Yx89P3NRbMsOAYJgDcToLq
Qu0TFXUYC/6xTkAzf73nd3j5Y414OOF8Uq0ZSL2ZLiR05ZSvDFes7sSIwMeo1vLX
6per2Zy0XQ6AY95d/k5TMahy0b27HMHCOh9ITeBRkxI1E9EbzEqb+jdEc9s6f7lg
XHbY3Z1soXWUujm1pn0a/CakZ1LrUPM5dFwiCtorYaEpKwONEkXT3ifsQa7lQriV
zNF74SwEwUwuDAvu5QqBIy0XoCdILZOY60z9Zir62mftr4SBejr4UkAtcl1tI2Sq
6auKSvpmztxdLCo6ekMFii9kDi3AHCZChHY03gNKvc88WOSh41ODU93M6jrWsyMo
j3ugUfZAVkswAks0abchJyFluKEV7iGdLazswfo7nvbZg+cCa30UgN46z948oraA
0EOOdAIbqzz/oxr6h0E+r/gu/wjfnDLqA8wn6ndZhtu+tdh9hl8BIQa1Scxz7Cdg
vfcwIeVGup8glcBfhx9b4C7xBfxpp2yqRqCwZNqFt6I30GCjKYpky71MpxQgyge+
g0+PBnoe/RtxpAvSrsNjeZHXNu8yGpFrYR//v5DTG6+UjDIqbNbMx+o3sVGO70lA
Vd6SigcCuJHf88mpQuBRTV+5tkNP1ue7AGIfGrVritjJKkseaXN3nkm2tiQlzmAZ
LErtaKsZBZ5goqWEeUpBwiLtmRWjQTnQBsdtPQu76iD8elHSAiwZiTNdC5M03Rn1
WvfhlOwtzPg8sfJeRuoaO2Wz+OZW2oFKnw6X0f7tyCJpB3+AVbx+cnNl0n4QRzX/
uOkGSnyBzQp/GASPZslUUgeJOczxDQ9R7bo4JtX2aEGFuG+JXO6g58bBTo1jeKp5
1qK6EzcFqeXGDemz96UYMTK6Bs5CT1mqbiT8uB/G+e+KyrDxUMGYpjg2x0jdN0wx
yupDe9X0lv1QF7BKcPR+BKKuZhJ4YeYiImg1adaIfgl2l/Ka63omg4q/0+aBM6Ln
Ho7gBJDaH/3t5bHVDIKCgXXGaJChVHSG0271e8KYRzfFjG4za/xDZOse4febN3oQ
RQ1L2KQ7UhJbdOshuV6UWtopp40mb4rM6Y/RbUE1kNfEUIuqIXx1SH0EuvTVhe+M
yna6GKosU/yf++oId3gTxQcDhypbELkcR9uLfgiTMvP5sa/PHau/HFtsZwNJY6+m
2PJtHQ/xxpjxz1ZSCEW7LAG26ZXzlnss3r1dxVhHTeyWAEIsjEVHsWDHW8FnJ4QU
i/ijpn8/+t9I6I1W7WEuTyuyyXIhNd0dWU6Iaju0FQodgc3CtXEcnIJDS1CUAKdi
+Q2BysqPsfQiOx43fiRBg2gC3JlVX9xdW77PQyZhoJoIF2F7VCJmEqVk0ClMP1G0
1SAbPLUOin6JOBFhQ2mdbM9mQ65JlKLAY42Plo9rRt/0P2tdDKmr7NHsthpKLNZa
h/n3pjrvM4p2+g7Nd65OzeoMQYQwSVtrDqpkwXdOdvPI8/h6v58bC0PcI0xPUCYp
POgEWBHFIhGSKbPpoRT4P4RJ7WdJ4X/kvV/TmGlmjowqiM4vaGp4hLbY2ab7YDJV
fscCpk4d9hhl8/aNP2cgkKAZUvf2ynjuX8JyzsKNsFRr6wvMpdScmoA7SZGyi/W/
OqgTmX7+T7rDcGXxmk/GS23BCzyNg/I9yF+2Op1ilQhFj8jtdkzGplF0SaxzIi1O
ZClfzqkv73EQSFsePe6Ll6lJ5a9AH76/MZtwlrJ9phC8EtqVjwJI2c/Br59zKU0g
WsDfH5tQnNnYfJSnh7w8L5fiarhiBVVLQSSzSgicNq5pEMBjzks6ExQVpCQMeAl5
t/l9pOde97sJIwhJmDKUOmPRdTo4Hkqm3OcR9bVPpQVgaD9jPjThJt3VG3D2HhQk
2oF7buSQ3bQ3+kLz8wrY70WJwCwXOjbc+4e1XQH5d6pJeK0wJ+L3HAlF5MotO1zR
m33nUgsWCw+gICU9+N5H21qvlGLANIy+ESP8AcTVIIV1zgNNiVKB3lm0Ep/jIxl7
Nf5TK6XAxjD0FG3peS+amameCVg/wcIj7QJMVuv7jLBX1IccKYFGhksYsbPiZ/dt
Q8UFy+lGTpBBn7Q4pKDTKlisyz+yrASHqt9yFk9H1i8WR+bGZgLOTRV+f8IccOLU
nqqU/XkXlsR7CyZUdTF9Trck/YG68GCkzcl7NSXxHMS3RCr8hB16BXVClgEcwIFM
rM6KizGA4xjIKuxs0m/kQsVuYt/IMHw/yaM4sCYIASBWTVzHX1keRTitOfOKEQ6H
aG1EFfdlm/hBupuOlDN6+1t0KYvofakUFG71hYNNGEGdjlvzfOYQaZB4bOnOKXQr
XY5LfPcsgItipfVWW7mu5B8zHn7r6VWZVDk3rbzUpRHN7KdnKObsN4yx/OMx/2BC
kUzhrSQIHGNMMRB5Xpbj3ZEpcgiUAKAVTanqbVw7Djyyn7nsuwpCoDMeuRoomT5B
YGJy0uedzw4vgGCtevEwnxMUhfx5EHXcBJenAhEvyhDwcS2gWi5xqLlNtZjOJoRP
XpiULuNV48m6YYpDK4LPmGr8ODnqJXie/XQoLUvUVDx62PbWUPavEbfOgvAFMM5Z
AXjNDpfxMx6i/jWPYNTCdbuA71IC4SK5OJXzekI6lhXvX+L8MdNu4o5KXrf0k+tc
Npq1wlk1pqXKlSZ66vsi7QVEKk2cxnsdKHysyRi/SdKKxQzCk3GUORdQAGjRJs9O
gt5Cd19TxjaDEYdIxGVbcQrY0N4AGtF0SthBYLtBJbWtxCyZ9x4ZDasLpdNUtEyS
42XKdB66wm6exs3zkfReCRoQsHbV22/UjQmjDs7ylTHSwKCGv3IaVn+02GrtOsiu
OPB+Qt0j0f7+/CkKziD/kRXDWjlmDNvpMbmv7ocT8Kias1NUydvSjQ+uE3BCrM/K
9fN0Exgk9P+c+gxIxlKUbINMc0rbmxfLdK17MQKWCu57JCStmVSbGtKBy0p3ztdy
7BU0q96iN81JkSa/eGKNZIUnng8bPlsmyUOmOitbMebssuwMZiDjWa9oYnlbBKdL
Tbz9xxL7877y6KxDUtoL1iRCADX7STyk8OhLE+ECy4qJAmX4wJn0wrlceS3AqfDk
uWUjjcCijXcTh6GleBmqFmwTJEvm1N6J5wpb6wGXgUrnG6AXUhZT6eIDu3wRxGcF
E5nh7ss/vMgpB5fSI4D1ImmgkhfqqMZtvjWWv/3R8HkadTO68wcza0d8MxKL+h2H
5ya7pJXh2FYDxb6oQNZ0bHx2wi2MhbGkfLvSzqvhURBuHntqGSopMNId0uKWoH6M
2XstR1x4Qhrh6ytgk1gq3FUMH71Y3HHxizZQih6xJeFNBlGG+06rxfMGatmCwd5U
02cKak5n9S8uEgYjh9JFq82Dpl8eqBBDO/Nf4brG3c4cqvYMdP3N3iLK6BZ6Z8UV
Va13U1bquvuAM5kw8BiDNF8ggZK+y3xqW2VLpddEBxEtcx9J0C9I0hitjePMnxxr
I0e3gC84nKxDPVNsAh5Fkku8HhxQnHze9vGUWnNssch/0ggSkuZ4oldTnV8dpTDj
jHr/UhdMMNqXgydCVfjeWwnBR01z+VOTt3KajE3YJ9Pv6Y9zuyPV5bOJW/Tgd1LA
dNr0GXdKOybaYgsux2VHocPEfloSza2JmLLwFK6iprl5fWxVuhMuFJWXu2ryWqy7
cGMSIM5qDKyEAM8lskVnuBGfxBdbGmo6lumy4WY+2/KlTST02oWGTAqi2QNBcJwP
Cy9fgytugNbHHqsBwHxB0mXYPw5jPB6aWX+1nMzm5w233iuskxVWP4Vn0w12xk2s
UBt4TiEJdjAPCg9W03+ytV5KYA8a7wedWKxbrfmtF2y7w+L0pyOndObnK/lNbNk/
YdYd5AIPBfvldrUMZP1TR0WPuR87GLAVi2PIRpVo59kMMm8rCEBEzfhMkVSx2k/f
Koz0xsBJJklhPkSUxjcuXHaXVq/HyMNIaYRnRS2ZSmYu0wn0Jly/R/663HnGz+vB
/qDgCmfXNd9BnIEACzjAajNfU5/sgnZRvrAckkgTeP7Mr0NIfyJjkszCw4FJSolQ
FrPIS1bK/mGSoOYekAKWtosI9flnsapZEM0Wph6WCNdO9VmFENVoJ6Ay/mJ8eak+
XFHYc/D5l1uTMtHXn2NBw28NZL6FGOTdQMbdSKeVynwBbQ+VCzLuuTbVxTKHv9Lf
gtp6YD1PBmkB2yxxngOaZ4zauk/a6CSutYq/UWBE7ACx/O7GqOudoy6OOK4FIxKF
TcqhTjZNgsKRNMUATlR02mPrd6F9rn0JUYA72OMhNHt/TO/+uXuQ3xsLTbIERW+W
GTVMzWpN4SxJwAUpY5AyL8WlH5I9fMo6KfwhIB3I/6AHNXxlk10LjT5coX1RDxE2
CdB9a+DT/00DSMbdjKBp+6HgSxBN7yQxvdhoik+ZMNR1VCgosCp0tfLnI7QAndAZ
luRX+l4TPLmiOCKZ4IJpDUegMhGHhSihUvjKAOxa/azVkWKky8HMhI16Aik68v45
5QhKUFJ6wi676RJtgfiLVM99lDVUzxhO6nWv4OKiF5UqbKXs5/VP8ZuQVYNk+N28
uLDiVNYsAmXcMXrNAhD81Vcz/OsZh3XyCIZeYjETYvuSZzqlI4RPt2zNVUcO6+1x
UmMbK+5f5e+7l6Ao13vUhI5g/ahhWUYIsdxmc5xHofzany/mYuXO5rLGK7M1ZI4G
xu/KRd0WHfePUjToEYS7cejwsm5r1gKHlsPMTQ14ODQUI0PKxya1dojgwfeqEzD5
D9+TQ9Cab9bvSR7jbwxUwOzUSswEwl5jNhQbspJuMWkMuLjdMzCU4jkNL1cWkYns
9bZnt+fzWAMgYGJyFxbkUV3vknGRGfU8nDw7j5IgUI5zOCJ5VZdzx9mSqsBQ+T48
9SeOutrsO3H5pdDl5XT0/zT/Vk145WNIKyE9BJPJHvBXoPFDnCXAVr/XMOSXYVge
qYTWXAMs6fIMzlPBOB+MiR3AUOwZ0Wt+uuH9goId8k2IhhUIEpLSUQfiXEPXbHxy
qp5kRoAidBD3dzzu2O0Ivp38fmuuVTgPzBoxr/daLsZdAd4fGczu2m+h8zoE4a+z
KsZ0+TFLkcx1E5rKtSh/4y6KdC/d09RnCz+gl0DZKBVcQOWuJlFlCbrfBUw3mFMW
gZVAg2qsISEnkCxmUryuAfjDxx2NtBfHH2EOlk4Wvtdjuw7J1Wl9PfKH4z7yuw5z
40aUUU3BV3LUI83RVEk6N+x3C7cxIBaguk+NW30GwMnSTr6dwEEf104iO18L8gwV
xjLnaRu1OnrudaFM4A3zmLi8/BpFk1VFPaaTD3UnR6ue/aC8ULr7fgsr6k6T2Svs
0g8cT4XB8AL1tMDL8f60roMqPxTKUGFvK8wRFRqsyJXRz/5mrLPFzy6xyXte7BJY
5lgDSLLWtGPjn+/kWTPF4OdCADot/0q8069xrggMSvKaWhKzNgcemc191OJddKGX
Pan0iAQhI1ycACrgs+e8riN2G23plG0DUOtrLqS6h6W7keWROeMQ4Wz9RmEtukRX
0kuEjq3QCmGjePJ2EAbNltN86J8LYQ/Wsls/+lmNz+nDtbogFB4C/nso8uo6bDgY
WS/vkuo8bdHx9GXqkeElS2GnMl06pttFwuzRjYLfoMwzoKiS3zuYmlvj4YQmgfh5
zeRZephNRicDy4ibgdqE6wwUaiG6f5/+641U+Y0Xs4slBDgKmUs6Mc80SNmgnYW+
91llAzvgCdSPZbPz6LWFJcghNiN4BezyIM1iqvndmCl7wbSPLpcXQoluzb/ZTrSH
DRIaBoRzYqrNPJ7AUpAEnSOGBh1sXuGFOwq2urxjWXGyI5tQpUsvvaiAT40L4/3M
gnovXimTuJnMPk+APDUTYjxBWToEFlWAo5wpF12KZJ/4Lu1b/YEzEqQOArLhdOjL
uZXKzlcpI+XSzpHsGMs0ejRLHUvAuXicjIarD8zJbEW5u95h8ThGCQLrBjA5WP2B
SjHnoxyxvMkkxOrR7pRTz05E9QthlNcNPpjoPCki/W0A6h0vf0UOYW1X+kEkMS7r
vH0bqR23Iv8R3bJn/ptW1z8GrB5JFjntYiHGy2AV80p8M0Drwv02OBw8o6orSuv8
+bbbdkVavkBrU/mEGf0NzH6HSlPlWWU83+fVxA8a9Oim7BxPL+5IMHYx1gaRD6tk
NQRDO2s1Fw1W+lpE/9cZyNwjEWXMqdFSKrdr73CvKA5GlrM5RlEdIk9HDcT/16BL
6iFiAGgnObhGvl5Ssy052nAqGyWWrSCaBAS+gcD1nR6Vl3A1IUSYMdGed1HFli6j
ok1UJYy6PsTGIt9KdfNRw4WuS8aF+Gmm7VsUV0fp6IDuw2bKDhKSPqNiz2upt7IW
ArWlueseaXZvPPnmI7MFZ6sa/umVnr/xXaqa4qmpeZ4OMsuVrOuf956QuOQez41l
Fs3CpI2mtIcmuBkOFVmiYLfhEVImPLbxudszsydnaZQQQ32Wyxx16LAxLeSZPy+p
GtJ11N7KITuC6EvuOxFIffnukBu90zGKvGRvzYwY/0VChca7GU1vlsxubMX5/8qN
VYYJZummxyJQi3R505/EVkJL8074PqrSHVviPrQddh9jAdbSy97AOlxo7zg/THlr
2Ll0EH8gzs4z/PJDIk3zlJh/IVaYjdjTg+uhbWkBDAvahHgOBlBBWtF8AUi6S46e
0KyupDNaA+IE97uFTkNa2V0bvE4hTta9vE6CUzNg/p8CEAd4Y2qL73dkPGKM7DDQ
POz49ctrC+OfNLnvM0B9qj6+7H9WqeWOUla+RJcNuRW1TTYwVOkoKCq5Oae2bTpk
Q60R7Xvc0/0rdN+Lz4JqGPcnfWxlFd7WUP6EpiZsOEWOWyuwRvsaHIoNGQCwkYTm
jOMRmRmksRNHmgMdAZMXJd5qdqhcunggy/N01K71LVUQF2ira1QygACBIpYBDlQ2
ufEicDDaeSA5A4VhAupNGgtbHvV6KfyEcxgSSnkGT1errNoQO5XtyQaH5Y7ypiyI
VHbwgG9KyhwsdFPNKfpF/x8cnM3NFjnXoX6aaf5oWWsUBRf4XSkjZRNOVx86LYyZ
4oJegMxYemopy8lSDz46x78oRnOkh/IRG3jJWO6mRIJ4731ypyRBGMwhXb0ggEpK
Vs4HVXg/fG9cmh18mLgJiOcQ/AiPUvBFBZZCgzJrFuv5xnRUxM9/gqM+LX7nglhE
F0o7v3VntWRV3rBN9qVRxqGd9WHY8bWpdWHbJGXQaigtdyvS9JOcInUx10sOYqgc
2FCzOvcBXc3jQSDqnlDnRQh0OwE13xuetRoMqUzFhTc2+2DQGTIiTwhd5EOu1nON
jdm+k81A2u2I6saHC0oj9pjGnKRid1p7Kc+EAh3jbAd3X7n7b2rrCBR8prVnV1ky
k0z+LkccfBNPtxm3e5RXnMJ3dRD4Dieaxu7IVRTTITOgdmmmmba5YgXOEO5I408E
g8dVBKV6GV47L3rTfa+cW2x6Lh3Wsc0j4jpv3TUQbmlUukOFGyl5dfDzicgJeNi3
7JZJiHe2CCn0Vgy1eOB9+bOjfAUor4thT5w82MwEWU0IgD6RXQgMpoLWlHcJ+Tn+
eL7e9kJ3ePFiArWTfzsVJ7H4umDmjVoVg5QqJS1MCqcyqYU5OfapKJZWfzDZEemN
UTvvCx1Zc8ySplBkjteAfhkb4rowVDdHkRPKkfn0azRb6EZ2dF1Jqp1YiMGvDaQz
LZzXlYg5A/+zNCkRj2jZ1GNlDzIBLQW2alJTllt77lC6iXTbiXrK0gkTVT/+SjGp
DdVp7KTJc6gIe+r2BPODygpeGQhx9YnSw08UH2VEKUhDSmwBX40m1CY98qWNn6bE
ecsYmvqqD8vY7iNKV6RwRlcy00/SjnPW2Lrqoy0VvxkpWFBrSWhYftlPeZbriU9B
N+606Nncf7YPdC776Ci6iRHdq6u9iXk6d8dHGdpm51QXPWfyLv0fIpsdNAJD/5l1
yVsdjMGqWdCYeCY8OB42NXa9kLZ1HgJlD2o8wuAxcf/HzK67qXhgYiXHj9XZLl8x
jgZQB+0aXaO2Ekg1SZhNfUOSm+3gI5oJv/YemY2JXDEbeozjaOlWF7rEcqSr1rq3
KdeYdFsUoP4kNQ0IuIZV9odTGqhkfi1J15GE+4s67T6g+eWbptjGAoHJnf4wb37W
mnITL81QN/dHpPYQL0n97VUjAZsVfHDWpHtOcSx3hywS4Mzoa/1lPDNjcyTkU+DZ
HgQtGr93I14L9cFBRvDBXR+6QSMkMv9oH7XERDqVHI8eap0iKnyTYuVz7zqvlBx2
cEc6FLjJEKipKi6EsnEVNrcpmv93n693fbj9wHe8FwelT7laUxZxNFLiU9AWbSYU
mp2wGOl9bGpiCAaKGHbJcWbDWECZIcLLbZHiQZ5HC30r5o9pIZH0OtsjNuMuGkuD
MFg4MnMR26e/tNqXC0FXfjmjnLd5/Y1nU/oeTzbxNEQ6pOiyD6c7Eq1IKAexmp21
T+hLAh413dVT1RkxokwvdB04UN11USzmmOqCG2pPBQQQP9PJ1umErMfzkaGY5FhK
EhzRb0ZVaK8Xv+vYbSkkHllGVqCfOZS4mE6QqQ0tdWJ5PRQinKZxN3qXLN/PFB9c
XkuiM0SW1bnpBoUA2MAUwBrt7EJYqgjVAd5Jojq5+/+xUncldVO+P0kqKeRpYlBi
dXRb5TglYdkqghmATmb9oiGYmPwThxUsCA4CtzVBO58AGtUP0sDrnltDqAMTmukR
5Poxh/QL4+FF1lVTDbarvZlILECWwsqNqRegA1pvfGMbNwy/9T8YDCRCQx5Cq6VQ
xNnCJTpTVIzRVYfK4JHU8gg5cCgU00pPpikkzRZsOtPuzXzqWD6xgZgESOPlmV9J
gIRtF57Vwch5I+lhZnxRGqLFiqSI0/ZFN9KFQfUlNpRWzOoLy5TfzCqJUxRGEz2N
AAMa872TkZgj4UwHAtuvvPRLFrV/jLDbIz6eGPyxiC0CDC+BR4XDcqxJ3RzpdeuD
Y7vtIf/KVd/m2mn+Ry3jamlbVMq4qyeLshzn5KUNLj/7Uhc05WkQGtTWEDncrJIO
ldVSC1nqLBVw1L/VSJWBE3kqc3vwfQAv9qFws3PXzf6di5ajNXvBEOhozxK5QHKC
wImqGGEuEXDhF2rTVHgI51PcIIlOobNzLHfgoBxkBF9iog9d/4SW7tfwD0bRsCLd
Ao2D8QZHJYMICYUJnzAh/YpriLDlOt1VzN5Zf5XQtQS3YVZ0leg5IbsHh+kF+Vt0
pS+RqdJyyQB3EbIvYels34hta22sqKBl3monaerZZTud+rgcqo8NtHG+qOllwSDT
HOSbCiNgrfc41g1l40pm/4k6eaP8v39/7UNVpDttSRFmrVqiIMHfGCybqgOk936W
dpVjNzBPoKJus4vnb+vukXnBxO9aNcnqGn9EhyLuPBlT3RhMcXyYkYoKfRao1SQx
+ro/Z/Pyrzp08H9otWL0f8MLy+MrHXooxW9FIzYKs9bCbAIwHKtosR7PstWr7lMY
ZwTkxbVFygsik7pc0zRKUo+F1fYE6l2ffaxtqxB/ZYdXGaMxaUQtbY9FI8/dB2N5
57DJ5Hm6SO9UFCT5OSt6TiTelimBFmKsRuhnJScN+CwlJGiAAn0wOGSUz40BLreS
8TMFb6oOPop8OZEsB7NUXCVAn8B6l43b9A5aybu+mEbYZdyBrfl8ipTdoub7Zp4u
UQ2UODETVRmfFo2Avo0BDljKGArBlZ3QXpxg91eHq47lRJDazyTmooHLMNenvpLn
i1MXrn0IUD+Xih8bBQJ3IPa0Kw25N3QWAO8gEsCRyWBYXZ/+6MS8A5SD8V9yQQ+8
oSTljqehC11YUHeiRynYTeJmYYzwloBHMVwuRHRGnNdXDs05GipbT3rbg1HrgSC5
8BjmvPiFkMid/ghXXayOKG/rm4aS4yRMpVp09osHI4DvOZ+bcnJVRyLJMiLPpP01
sWBKCFxaniCx1SayH9nPYE+Bxgb+/HUBmrmbhBVl1eLhXqsoPy9vtWGG6yniQHKZ
Zq5e7kvfG9a3qYZefR+ZyNTEX0sQMc/3MEoM0/TRH2GUuq5FWhsIZvaA8CBqWtHz
5V4hUz1J2iBGCtXDpsEm3Jetc179xZJ5nDuExzvwSyVRPhnjTuqwT41TAjcco0/M
DE1yKMnug3M4q0IR13oSOhimwxy01MRHSzIFF4TMBjXrLSX7dA0duS9CChVMC8x6
6ZzW9SWQOMxWd1uQz1MnICCProD5xRVmSRVi2F48qk0DvT0lYjcpenSB/xyPvfdR
2PkGOjr2XYHpgGQRg8J3+ilgD1IcDtElHceIC9z/XFQPdlUbArFdcQWs8gpU09e3
l+A6ztp3QTJTXRfwE8Qgy5ydY8j+elxLTNWPgNLvbNLXZwlqU5S8cNu4wl+QKGTa
kmke5APUTmldLWJVyH0E/a/0pVJHMoQmmSnMbHrL9mRAnE/WlanbdHNc23GTjg0U
aodLI5xWAWlmWmCZNXFOERoXq++dBiqd8vcjnST8qxj26K3JD362UZ9PMk1U8g3B
OPfv8USYSyRCHdDOY2UmhGHpLr9p/2geUjc7IFI5iklIOMImDX4YiUImTVuBxKDL
XThVXpLEn7v9eWMhAAnqUugZK250Z6swrKXE418MODpZDohrEruNKVqzlxcipZCg
G/tW5uZu4H6PLR3WkAdUY/ottvvAZJagCWVmZioVQPe7m9xBLLYXD+slMRad4slo
HUS1Xlu1ym4VB8KHAooa0pSWUOrjlzxw2YDBxTYkJ+SS59Lkscrxq+tbiKEwe1B5
C1IziHZlXdKcH2s59/90/Lct/y9r8dZwvYclEfssJMXR0UsnPi3au7s5Cj6edQ4Q
wFk88fUGRGmFLKOGSGTtzCNA2GVh/uUtRu3fw1VdVHAvkO3Q66LXYOrzvJcn/6ex
paikVmNqtnSBnRqxCbNO+9bNPO/7mKAabyy5xiBYd2Rp4XtjlxQc/PKndBpl4OiB
zf+mpF/iC/oTGH3k3LvoUdz3n0NX9HQ3diJsy14o497rf0X3EqYXaUNpdFqcnqZY
o6iyWcIPAwPjzICWBEzyiCMF/eSNAPDaC9PSMJLXdgFbhUVxa1UEPcYbAnsewNWP
BR6O+KVhLoPUvz5+a2b3whL9JRJ5ILZsE1ZUufV2GugwXrDFmajYH8/Sci5I/ndF
i3iU4A4/U44bsvGVgIwqdfEPHfGlEJUlThsp3H2HqBD2xGwl7G4zCvkQM1irNaVQ
wt3vtk3J/OSC8T41E9ST9VqDArMFNk4mC0wXNrsRU7gsijIHz87K2oiX9GbIIdqo
wMC9S3emQld3nEdsLbZtlPjgVnm3bZzdcZAq6ozHmLxfMLmZm/XBsTvCXDm6+AEe
Iu4niG5w5uBy3BK5PZsFqFMKg2vmoQrIx6838HBsL/gMoz04RDUbSVY8p9G6VXQK
JXRjEow+j0YOHYTPnGDzqw2waAbuK13+evgf14VRZ7TFNuZ0rXJPepFIX6e+bkus
EaH/2e94OO10ILPpKLXsGTrOI1rHKNh+KzNb+INmL9RA0+0KbTOBxmLgnu2XYkuR
7e/RBbAooBDBCCuZS4hEm/6jPM4uQt/EDKt7/K8Msvoan+UKxZS2e9R1vQPyDqkf
Uo/MjQ4AAMLbFj08f36Ca88Skt/DdbUdpkSFAXKBOZcuAh4/19NoROfyqsQnlGuk
suANJDvWXaFNKXdS2Hh85RxOxkdhCweq6uC+60Ce6Cc9qvAvOEAlSNNS21y1xVN5
5TL8nIydcBNG/7noAQogCrNoLqc8RhAtreGI96mvVkWV9LzoAGcMJdxyoFdHDqdt
gu0TchXVz+htJ2QkXuwliZMvsqn8txvsKsI2W5bhaj1nHp+D6NOT3Rv7xJQvyOGp
uLCE6rjMiidJ7E+7iESm/JHAujO3VX1c0tJBKDGSA/5XjjMBPLPpWjUfow9kPrpq
fv1X8XMVEi2i+wvfM8WUfEv9nMSlrWpxTrzYrCWUf/yO2QNLiX2W8fL7QgvEV18W
0fqJE0FiwXB5hBbDdgJCZuxcvCX5VEQIG0/FAsreVnljBhEvtRRPJ+Q+tl4nrbyS
6Ct2rLLYpMgeibkX1aUdSPlWpYpUdC/EQfuosaRPic98Vim9dTW/oZsQORznb2SG
RNx2y36MeG2lrhvvnzvPCCW01Qw5WAEuJf+dcqWHTWL3hEdFCdqoZ/x6PjF5Wmwn
IsgHvK1x/NTFAi2ynT9ph8M86ycuKKpS7hmmjxchLRNOO5DeO+m6TbnfD/irjLT7
nCSRyOBbqMSeacg52LtfPgt1T0by+AlPMrAj4H1mVTvxrRYjLKck/pgmNDIlZEVD
uBMaSL2eKkqzTZHhCHb8cm+9RnsxW8Xtd7oMgfm5YRY9BGKVNODXrr7ahKJ7ZP54
EwqBHPdINVlpnSl/taq6r//8Qre3cE2nYGCSqdEIkqRcauD0eQKV8G2NNBEDdfze
sotJpTOZKNoU5N+Ce4CzkWHrp4im5xv4fhgRfRVjr58foMCnH/BOLkhh7sQRQsO2
dAxoICzQSw8fhdox4mxsbRWEkvKfxJTv8VOtNZoYj7c44x0/70lSayEt8A81vxcB
qNTIJOP2ivgXIxUJFhZye+Wezlssi6V922OIGqcXoLyW/ig+F8AY0edCsEjkbEHl
ioyGXMXku7RAdGeKx+Pv0yCumNfZ29YZENuID2KwqI3HLXGsThB9/Pq2atU2jdpg
4IbkamDwWEFX7Ire2PGrCfbLP6i9l+6rBlXgG4znhRflE6pFS/x3+Y4YYBeGPkEC
YBn35QaBv+6mzcL2eAdhJVJ5X3tnktKQ5Zx9OCCYo8ZOsMYIXGYg7LYNZivfTrtC
P0W356egrHWgHgUT8Syx7V81aTFFDVbL8BdoCOXrXpyEyWch1u4UHQV4L+3/ur4x
+RGev0B8isfpA+5m9/SkIoV6lsoYZDnjMS6npJY6VyEZmqfDMovM+2skkibWGof9
FXHCB2QeW93nKTRehzY1TGpkc75lCOyVEd1VNqR9BFZnoPWFK32kpJVH0cuxdkiR
rW58Looj0FOhMif0Pm4AxSSe884Ytf3eKcfPQkgzXzXkk19c1QiOk3i4kirV8XB0
jus+pUJQLkxYf7G/jnVQ/VQuoITZaKues+MAGhOHeDSq/rAFsmJiKKjqDdbQLuvx
ODxlNEGmSJs0BiOas3LU5IWA354D88dN2QKW2oT0ZnlSciHMgQvD7TVhaj+otdVl
cUF28NY5ksjtHX2HcXHu/MVJICPZ3cQN3K6xoKyVIYFbciuEvSFvmuERNAtN2JVU
fRDVu0TWs+jds7dHYMOIGdNWbMfDytj5+XMNQGb7/OkpPnZIWLZ0xmMQOa/58Nzo
vmVE6z3p2MS2+U0/9VxqjirUs0eGpcVBNg5ZNmb0ROa9lbiyMQbajwRlwNWLfn0F
uL7apQJX8X/fcr7hQezr5Fn5ZLTfcNAXPMCHvEItQHsEJSqzzTZ6P3iJ6sibgl1c
yt1QuSfPIUAi8B0Zi4lnVjKr9pKrLbI81k23WyqG+s7gCoEkXL2653F2J9apg2GK
Fmz55TWezsbHAaFv80+yzkxZ0rK1AuWHGsEp7Y8ZUKmvCtoIHFTGPLeP4SmlIWBD
zpnCXcDsCGTIZOCV1umcmd2mvUJagmFNtBKL/Sa//uRKNLNDVedp991KBwi9BDxU
4f4wwGIp6wZS/SvG3I/G2eOd3DEzTN3TQwgLcf/W90fjc6j6oBVe5xiV2dC843Ro
OlETyW+uG0ZnOWuh6SdFPqJgVx/3ZFS2NdbU/yoikj0eOAKQiO1QpNqVe/Ji2aaU
VvlWby3nwPG1/8FDqjfV+qUzqakcqp8BwoY/v4lC7NRGC0GoNjaQsBF8byvVk4N8
GHROqeEr4yP1z4etS8SRB4V7OsOzX2SxtiZg4f+fq5sArqZgfUSsHoLqXOhXb9B2
7ie5sQVuyK7shd28K1nEG25pWf2yLHdhNqCtv/FMClvKWvUmmcQSpAJVgv3hokbc
M1MQkwqlMeUBRcXy66ay0HO3Yrj4f9C8Z0PxLdY/Rga0lZsOab6S9UPDxCJ6upi2
IW8jIbDw4E9guFo+cZtpKL6IiA0eauo6hV0d5SB8eKowotXVope/n9xrWNaK89iR
YkM9z400zFkzFFTvnjyAOLzGYij3pQs7pjak7MnAtrB1vs6g0qPh8FTxQUq5/Xza
SGq/eLn47HqQUgB1rULZA7MdIQkmRecHfpwmNJLFQ6U4lyQ9FmKQCYeTi+lfg8EE
kt0Ti5uEKYfeLATRynrsIrpb/17oWC2h2/fOQsSQfVtyHvixqE1LSbfgCdl0KZmZ
VxHQK/G9ljXqWCTH5XXnRIxS6Z7xJH0OR4VUiHQp20W7guneHmtoNiE3hWctb65w
WAD1LqdTxtsczT5LW4SPR4wN9Q+9uKWQF+Mg/KbCCXzSYiZLd/6WpJmzZO7ZkwGL
Bes7aJk6AiH653SlICogdzLNDViSSaaJttDDYKFqxl0VLAgD96L8QjOPxPm3ik2D
7T0XNT85Wqkg98Pm3MNHJ9BLselBXmWiUy+icjx0rMBvQ/GAC3VVFSN9QOzYAMsG
MlA4CB6gze9Wo5RvWFqm+fBsyQdlbbW0XAJ09419zka2/+AD7ItmkoggzaUplaux
rDmY70VrXq0k9i1EuKBob9RCUHE2e/gQ08891hWA0KS7r3AyhmaoAmNCq3jVIJEb
gK0SbqL7Hen+u1Xs+ALi73xzDsA38kzSD4LrCpfQrubpwqbcnG382ETN7GRdSqZx
M85q9xRd5SvSbTaFrqId8Z3JtBbyym5MEIMRuxelwTGUiEw07eIDoI56spc6BBkL
8HHZfg5OpWQUnmEgGr/k4DdIwt9qYMe0jlFCaTgJOvrk2WjEW8P+KKrVtca77nno
xE/tC/5vQE7VuEht+vCwlGrxdgb5ox+QPF6yk25ussq+j1bBdCdb/lMHP14MvjJx
tn20bAStVqrhCVGmXaEiUJjlxtizXqhNXHD7yEo42rxYgKf6H+EwnMAHdjjWdxy2
UkzcBtIX63h8/dpaxF/30xwDiwlo9kz8cNb069qgkT7GXfO4JzycEPHVAoOH1c8X
R1KjZ+rgWkicS5dMJvQpfyuphY5qyD2MK/vgKKzcFtu2eOGoBUUIVEkJbvRLahbj
zXYJoyMVQtOPro3mOqcHmEqVxo4EOTinEj6fp4TsnozV1IiDVAbZxqvdXL4NNaXL
i4UYk3I8YQFr7a4VNiHKb3vc4FiDGSdgNm8wx7HA44j+FQfElyt0J1Z5e8yGrI2v
SWOz54BPXIGJKkZE8m6vYu8s6QY7u/Vd1RFaIThfDsDN0TEOKxqmgA36AojyWar2
/rSR5WhB6tc4JVda5wp0dBsfNM+uBsAJ6m8PFZbV6Cd5CDS0Ln8tbwe0POibT8UJ
eBF/9BxzXoDPpal2miQLbgps5EcHmhmNktIhWCYA5B/cYo4thl/puUPryhD/iqdP
oZs2z8vJBSY4I4aWGelN8YuKeXYIXiqjj5PWKawflmzvmeSteeKhDheyuIgeubSk
Rnabe2BD7tfVOctmEigXjznqxS3aFqQwKtaBqhgEO2a+HWQxzi/1+lgFpJNHTfAy
d/5nks7IEyZ3jJQlzwdJNqdstSeC+zrp2hc8hVDWE0z+ygu0v8+/OtOM9Zs8VOxI
nW4MuthilxctTbMGod6+X1AdDQ/MaEDMlKEfJ9qwObxDO4WIIQ9NWpt+yHBxYeSx
YJbrve6m/rMVFhXEsF5y4o8VgoZVvtflfKkQ2PSr0JsCwgUoY6uH7NO/PM3blhWI
WcFsNzFxD2cxPwBR2C7AtsFo8t4yE91s8275K1s3P4pQyFJGvtPfkXt7UY62GbjM
ZhXWz9gvKn5XZTz+8xFFyus7h1a9IEbQUEO5aoCpDQNneD8eKFKMDUxJOMJn2PAQ
pwfsMVM/3Qoge+s38qrEINdLkb6pAQFZLgFFKYPuRWhNnQpfGVorfQqrmz8IObbz
Pdyg9yILCWTHv8Y6N7W6rWNtHdRE3oqKgE3C2j+GpCbYbf3JiViaf1samLeNKiTR
HgZKb2N3MZuES5knQahXUT+hgowVLc5botj9cvZuuDCT9RzynIKDfWf7TxGdjFZP
XPPtwnYs91wos1Am0eB5xKmGAKWZ53Lb3AD1wBe5TNrlM29Tw1RyrpF5h1y/qJ01
x4BKN++AVnJ1ejhOgtyHtpAo1KA1I/Zkdl1ahCAcSRKZUCP0kLyGjifwzgva8xdC
/OqXXetVhroYx07HzbzAMR17s4EMktVCBPQUsnkO6RyYkWwND2c8QtwutV2LUER+
kN79dv7XpUYUud7GJ2f2xwvzP9d/QgsB4HJUZYu3laolm+7j5x8MkoUlh+US1YOR
fvC9ztwqV8xtKEmRPJlforhur88LGWG7L/xPZqWxzeX2MMfDjNhhnK7veiAq99Fh
UoCsgZK+evpM4jKggXQ3xu1AYd5u/DXyjkbnStKRo5ILnNIRaKCANvXma6O9PJQb
0ygykl/km/1ib1wOQJUK3AaT/sYTHqgzl3K/nnhRI0FQcM/oapBP8XDEus7ay4q6
rnrX+tK/Igb7hLw+e020FFRNt1pDLfAmNpt/NPU2Ia0BVgXzme8hHSgE/mdQd0Ku
9ibSR0mnyyg/pWCbw7DQqhiJg7b1Ks8/eODd5qR+D44zOcM6cmI81xA4KTl/6J3I
1pkxEkPyLJeMKUhdxYn+iaDpZt5/W/6Lhf5TApeaDaArl5BRND1Lz7TbHFvA6u77
73zBGW0LUtJ5q4c3eLlHgxtvPFfhJKuUibm86QP60Eu+Q4n+IH6dsq0KVX4jEHr7
hdmWwcLYfxqf8NTCg/KRD6yALKkxAXkon4SgZsDj9JDaW1n9kom+IGtiBD7QIXSI
uqgLHpRohme/JQnbl614K+1dAi1yCt+0kzFw54eZDtR1F33U+hj8IxIuaTbH0Ur1
ATXCbW3elgf6KFIDg9i88QILL9+0JTqSjt0j13A08U4oxVB2CjTTdn2ttwUKoMkA
dT7M/3McjTBoxU1T5ROBO565/D/ljcF+NNQAPaEzq8dlFWVXb9S2Q8fYpvuqpuQw
wyQT1zMkGzeOu7pbSTl+lE2o4CO0k+NcOIkjTQ1tkMvSkG3qwOL2zIlZ0tcG0E95
p9fPNPUZaV2g2cU7mo/7XZPVUmnpyYpLCQj0dZ8LrWcFEmYJMRn1DYeeXpHcAKLB
gx3ICSxx5gBpk/YkmeHbDkqFr68CVRKzoHc+M9cPYYkDvChC5sACSB7O/5bKUgkc
c6rSb3YnQp/KArRuIj0sWM1WRECBgp37fk7IB3nP82B5NB4CnBLa6nmKNxdTndeH
XP4Y/fhTnUOQg6RsnumaZHTEJ7+3EPrhNoX/Upq2vncamMAiDzYS/3Q5BjOsnvSH
zwBJgkkOGTbVBzn2r4g9+VIYJCOuygF1OSNprzV/ZraE9wPYiGnP7whwyO5yAq5g
x4cTXNysj/ft4cQyEL2B+SU/nPRL21j9/TQ6XPPmWNHge72z5/jihx7mFcZo3Ux+
pf0vigulCHgpt3qCGBtL4SMGJIGHnrivsX0Qj8J05qdymATzX/vKaqh+8A6I4sDu
uUSV9Ucj8zYdPjd108EVM0oKcNFUOaz+d/UGIE5KjuazZ+8zSIM8rPZThCTexBNl
QoikfsgAmMYFDJ6HGFy2mK7u3o0krUoBKHO/YyRRLlW6piUJnrzp3pWs3XWCDs59
P46k2juPWgy088gt5eKNsHNaRnrOdyH6+EF3iQAdiHa22Cw4IVK1JqOgg8RYlimd
sQ5aBs+KjAYWKTRbL9MaO2y13otCf5/XjjJD4No23zbH5r7EeHeZKPZC71sYfYpX
0Yk/Kb8N8xdRRf4ZLr3d/OcU4z/oKOLvl8//Slg9aKVy/M0zzqV+8wELpP5y7O/r
ppgPvYAD2rHKo7pRMLTdtEtF90I3UUkQy387/0wD7J47dyPvTeRKG9wLiMjOV2qB
wd/mwq07VbJbtZUoJKfGo8Psuk81DE/4tDt85Zle29SPKBBYyDXCuR8A/R1MNBHY
BweTaFtRIYnzU1hUWZz1k7whoqLDryDMe9ct6I/uvjHJ8xT50ffFM/e18KDQn3bd
4Met4qlHZ7vGvGCHCqbWVB6EWj7+2WJu9eiCyhajrycNgnfZm4rgZKwoMecmDjiE
3/Idg070bkPLsNKUJiwpzCfbWizKOAJrNc3O9lk9v9GBMZGQMLZdPUyXoiOLoFk0
eacwnJqkj1Vfo3UWXmXIu4tfJaFGSPF/bRInQoiwrE3i3wGg39OGwwv+j/tNfxxj
Kr0bUs6qSsbgbXj5izx/1htBWcZ4d2aQx1p15BU3vB91tmMOc2c96ypFVvP04SIA
t+KA50cFCYnOXTQZd0TfomTWmQafCXAz7rfNPpe5uxaHtZXPw5JTEjNR+cqQkfcM
tNHMWOe0faeusP/8ppMPuYzfHl/EGSznR+mQZ8SOzzW5v3BCSAkW+jqdGGucZuts
HgTNzEFNCFHwH0TiuU1RINdoyvlY/CVn+sGSZmFX2BT/JeKOkwVo+fjkyu1UhVs/
fMuPmQuCxHCWiSB4cG+gE3b0dwksW+h8X4cioGsHgaPpWvZz08qtbeDnEaKX1A5T
qhHkxERQa9FK5n12KkiKrzrcL1BlJw3VhWPSyRVN1u7NGsO/AW4m9tew7F4OBEdX
3g+2JzPq3x/SWpX/rtMyBeyDi1kN5V2NBHqT8p+tLormE7gy/MGMqvJbJ55av9YZ
nMzGeb66aFDwk8M6pAv38m0ElY/SLrafGnwcn9RWLbmIL5pjhsLaj++A2CZVj1jc
KAdfyrEz9MnNQqoeSPSOgi1gqGsDobompW6lZZnqUxFdjvDfcV+8I+74byA7rydp
f9Jws8xhWZ0KyfO6P0+cdG4l1IrP0j5gTsU2faK0KLpV+h4CnCc67Vpu6D+rNzmE
jf+bbD8AOZBUehAZLDdDBqzuqux2D31BfXoZX1HmGoPZkgUoX3icK6wh8syHy4or
dAEYIFxv3Lt6jbuwAoYG2VzQZbRpVwgu/q4HkH0XI4KPjyZj6UKX4ZISyX7ruXqe
ZMdJkZNsBK+/gUYcsm3TozgwBkPXdVWA4GgZXvFQOYgOsj03OfZ28jkcAcVl2gP9
8rwn2p4TghI8XCWIcg61iEQ4aknapdob3Uke8ml20lHkQNh6gZi/hF2UygPsE+JO
GDUTXpuaytTP7vde7bScsL9HiV36DXmTBVEmZD6B+hMZoRDpQEH2f5kACs0X5vWv
izt4SCLhXji+QxmxfRhfrdmrL6AB88XG4V58TingLnNIOOhg05us8DGaJbLbIVvW
v1qqqNjY8vc3+lkguBgOQMBn7ehKSdTqcVDGwPLCDzpAH06MQGd9pizlAI2zVq7X
xSUNL160uEPCpDlroOSWWw7xr3KSKeF0XbI0Xafj3ua3tvjhuPShT3OoDTQ3prTz
mmepOyKzswjS6sPfrTcH09WCR0+AS4l2bd42HYJ2JMENjozPytUczzzv/t414a5F
9QASPYo4lDuora9F4ZWVvv/9d31jScYiVxf9m2kLPIYjKWD86wLJFg+aZqM6bsfj
uAv1ujQx0bn+GsAjeFeMh4Xn07DOoWVT39WiGRgC8Haz42dSUi+OigYbNnweZfrL
owcPyvrWw6X8U1D4fHvji/jkcfv/BYRWmMCvFg6b0OSHrc9uUmZxQHNi/2ohIQ+W
cZYn8lo7yV/B0oo+3QzpIe1eoIV7oeixvO2uYaCBkL6jByYrlaOn1/zhhewsxkjo
vSIamyKN6B2SZmUkDIpGD9cKGH6y4gW2cPPlhXUviJ8oPcBtyIj99TgmVoSmlWuO
O0HGBiyq33Rkrbelp7KJPRwyMAKwyBK6hUVoH0NVFceFSFpA6cOvUAMHf+Kjj05r
hi1vt9azWDbR+mtpKbJ7YSdpqKgWTgfAKmCdee+ahTzYJzgz/PY+x+0A1ekDh037
23No94tkGhOQmbFuf3adxocnDAAaYNdSupmmEbM/ymTMBpvDt6S65VJcrgj0sy/8
3mr2kGIls6U7fWx6BPpDHizFk6S/MBUA2Gf/JW1wE8hiq9Ntu9Jqs8HANM/EgDr8
bk7rvqFYixxkOqgyY+cdFaYfEkPd/ZloHzpWuA1oK5OkU7xfT7RMSYhHU1iulrU6
Na5I0TBHCWqPPEHY9uB0PWtB2P7TQzQiNdkO0iGpg971mXjmwYVpoxD67Qsc0Ec6
PKNWmuE2nCbqFzEOaUpnWndaSberkQ71eYSUPiKHlFMWN79cXcNPpxcMsd7h9Sg5
Nzbvsb434Jzz1wrfcU0bMfCxofl03sk2YXgMZxPitGAHelZ/M+j9uE/c54aEeGCu
n/QXutbKs9hD6MmEmil4uO3cwzBEVunEw4++mMGo/QFvdODUVnO2Dl7EQehxF8gG
gXBIsH9rYLWhhexfOPDblzes4212/yRHupNvvgQTT9bKJdD71xq6ss7Bd6RHWOYj
7LZ6LQcGPuFhJ82kpF4ag8BvRE1rLvmeScPqEb91OmQjmR9T7tMVJ1HVWb+Xpba1
+fSJBmesehrG1lHmStgxl+CKZTVO5XRLCbha5Spff6p6rhr9z4ooaJ8zmSu3luso
XfaT9HYLkKisVr2qPNyvBjqDRshTPCXVzD/1Kx3pAwVT4mc2APevazpihYgT23VJ
2QQrnzswOkFeSLgoTSgWolCNyTo8Iz2aAJmZsB2HMS7uYxjnRy08VM/WtdjIaUAn
XUtZcpdkicyl0AKuR36SwS5bw5qR/hEFuQdixT0reTLA9cMgmnEdilRFKBvzSy/E
rAf8SjTgJEDYbhS/rwRcC3ppdK14izTWbFcFOZp2m8HoBFmQTSb+pclz/qcBwNn0
`protect END_PROTECTED
