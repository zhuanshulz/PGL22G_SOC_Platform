`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tbgzvecafgEJ+MC/ZWcnNRI8hganico9y3E43cdubJqnIQ4nk5KUKWURaXCOSwei
a0qyYns1DL3sn/G1mjvZy1WNCcUMZRqmqecdVePpSiN2zm+u+jnYJQ3lcZ9KIi+6
zK3sn4LBjZWhdH0cWdfJTWDmeM7zGnAmYc/DPXHyJQpcRjQNxlJklwS+zFE3bK5N
G3uVdUVI19S0EOsYcxfTPNyZxFdRjgbi8R8fGNYbvNFIziL49BMPLF2pRUqHSWeH
KOsluiMJSlAYbDkP6OBO2TgwY0tKmI3/q2Cwd6gWM5e2bm4j213y7T5B2o1Pk7qf
TTFSBYUISoRKP64u4BvyJ27Aggl35rPpJ3oFnqRXGlmY3E0zlDGcXV/OOPXekPsz
P1+EXZEw+V9YNfEwJ5KEp1SFZdw6gaOEXNIGHdjqT24+0fMTjc+uszwSiNGybOq3
M6zm6iqnVpKofo4/rzwIMuE0SHaOk7ZPV4quUly81pJEusHQcOsDFam2IjVJhk2t
TTB3tUTpSBRsbnwqibOZ0FapHwFUsRW35aWnwmP4zt2OFpyZwM14hZ3dho47KNMt
GnxUtBt62Y02OrFb1ewRrLwOdd//GVAqOf4EaFh6zh5xLHYGE9mNanKXZ3zBq+H5
hJIR9qmASu0AJHmBm33FgTu2Euu+opukukv8W1QNE14Vk+7Wg5sEW/W+ds96r+fO
MAoqZHI33jIJ1ShBaroKkVw91MDckvqW1ugy/3rgIW6d/7RKyzDkGq8zkb4Q483o
wAleDMWJeWwSurLstg6IRVzcy0nuqno+tf9SkwKAUhivYupW3vf4Pd3h4+H5Dt9H
`protect END_PROTECTED
