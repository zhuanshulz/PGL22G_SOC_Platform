`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WcZbZw8GxigNCxhWd0x4Za8TAnwQKEUwa0/NkeUSHc6TIv2QlvjH301cYfJjnK0z
kg3j7jmTEoHkpm1bXkI/R1ml70kzx79goOahHounuJTljSu/AHX3oW5eqB33Gqie
tjvVjiGT3sJzZsmPqkEiC9127TwsH+BMU81TByP2IF7UOqtg+kbX45sG4EoJhXKW
h/J9m+AczG16t45ZKgwL5czHHCDuds7l/ab+vXFCb8oLag3hWhhEHfz8XZVNzECC
z7VvRfmjuvEDwgXKP031727DN5bC3KtzXJcmtbRoXRYj1koukLBlWmKewG+E9e1d
O5U3NG8WtDJt2uEASBYncrMko8jl4cxW5FRoq8EGHSWVgVubOXqqqVF19vJ1DxIZ
JEl0mUK3UljEbes3Rrwa7w0W8RnCBiwXTvw6TVmlb7kBg6Kg0hVYCrQXE46esOsJ
g2bQ9SGNhem84zmdQdJhkr5b8GvzEIvj035sgWAn4JuKRquL/dJcoLO+cQq5Bcjh
EenEcIV7evZUY7AzuOdsPFq+Pg0oL9YAwHDCJslbwhAQo+njpiQthSt5yFT4xYMK
4dxkEyzQe31ePvtqOZkXvLqugkAQZrNEz5RYlK7pM/dUU/ysC0qQjN0+5q52/rKZ
s0h6D5v3UPVbTB7GjOAqMmIFXcHn9YWeXCwW0kDKFDc7BjAUSUNv4ldoDxwOWHkv
gBStkhAtcEr3cKSMq220h24TEw9COuYmMazLGjd2LZyiJVjR0nAxx6JquYNoxA6t
96KRvaNC9j+/bgoA0xrmOIMd59pniLeWN5q7Uzzb5pVXeBwjQ0uR7ge1uCqlpyZ1
lljQ/H358x6Rjo2mwYpAg48dCVrHPH3S5/Hu1A1IIGiLh9uBgDaZgw/etc3lgnxt
YxAK5mBJdRrk5vehk9py+UHbJqSdeDV2FHCtQD4RHwXogXgHGUlndA5c8HUvLMTV
zE6xjlHui6Pyy8lA0q/5b2OYv1fXFtokkyD0aLaprRp0BiPfGTvA39uYAm7FNBxn
dzhSlJXb4ZbmIWvwzvkZ9CfGxGvQnZ86pQ8g19f2cNzyn9RjVCJcqUDdQcWHX1+6
RxGgan8akx119k2IkbxtSM7NqYrVk6l8E+Ltj0HVojXP7eAs/izvNgI4FY8mfI8h
OslzCjHDLhJhhbv78SWAET6XAq0gYxjnJs/ZEKQGCaOvcE/GqgurnHkSnLETDK2l
6WMa3ElZdnQIFjIZ2kw5TwFTdbzpKmMe5uMfCfAZuvRespYvtf1zHU94nzoCEDM0
jeH5JbxE5e+8dxRMCt3EjMqRsjSYPdwMq6zWCKdGfktT1fswyQgKw5G9Pihw6k5c
vnNITYj1Gfd0kB0MAIuJHJaWtPxlap+ltffJPbQLeo+L2M0CEJRmYASJkZNrbHTz
h59HLUusfqRJlmgHK2MKuSh+ihKmD/IfpMa5TaZge0SRMfpRprKjS92teHm7jlti
hLx4iVNxdEt+Ksp8SnMNBhXL3GD6sW53kLoCC9g7dxjMIcTL+nbk8KMQQuSPtBrE
u3y37teIhvRO8UNnmKhp9WA/eJvWL94PQWOTbkIJ7maw3j8jBElFz9y0AHzAeJyP
jNU7a5bbAHDcr2CY5nZwsWSC7RfdSdMpoZJJ9mH8qiDsQRK7qivOaXeFT0kOnI4n
jrfgP0acOEKdyRbtGk9Hbc0ymw/Ys7M1dCkfbMAURELbixyoNk/xePAYd1Ky6WZ7
OkY/ICSXBXXrYhu4BT8igTbcCPf9AaCjBqb9y9zOjikCny0faCzQb+YLfQo9MN3q
XQrJuqbyaRqm+BgPhDJY7eOVGZ0XzmNbMGbaRnbdYvc6/WrFCdvj7q/bZcEGWbmz
pknVdE8osKFHTqaUztx48S5O64oFBkg3KOxq6E14aO6NOBRK87S5Wpx+Vr9wiN4d
wUY3k7xRqzmr1fF4dYL9OLfO7lw8iMhYXvV3RI3seUFsQmlsSitTw13lbX3DXpGY
RJ+5VFtEf+NQE6c8+f8JIVPU+4t5KUz6Rrhe6CW61ofkKNInwTTR4oJzP5ivr5Ks
uB987PhwA/O933mMS7t/di4Z/TIu6LRyHDGg5I7vsG2twQVQCAWJ3b9krk3gPQb2
YbquGXXI6yKPB63bG9vdHB2BzOXn0UufusYQdpHx2fSU9ZU3DrhBF19yIYQxYlzx
6V+WFVgyaE/rVYKtTNsXzgGzybhp8+pi/6g+3czRxvmMwX/xFevR4VlDrszSP/hQ
caASuI4L1/zm/lL3LMsmjfz3qGkkGDQbCs+XHG1RLmOOJfLrD8Nx59OI4p/xLFnm
tbGxq78XEIOIsq+bvoCIbiIBDYEsUHQ3rQ1oIjBRFIZ6D9oLsio/vYpMHUyGtJFb
/GVYgZL26ufGXStKI2yfdqbhAlCUDJiVGHlLPyu+Jmv2TGmf+0/nxa9UHZOqFziG
EhWD3yzo2B+uRNuRDXLd0LNTTEZJA6/OS14hIy7wC+0T3uD82rqw95Z5o4lsMYBo
QSZf+wGWljLL6LAUu4oIcG+P3kBBjxuHBKfO8XFQLJIo+qoM7R15avHtZhZ0/7rZ
jN4m4K7aGLbJkpGWfIAulP9Nhxe5K4tozxm3B897Fb/PlrWjobjYBZ8rYVwx2AgT
a6setxr3zGTdGcfVuBZ5ziBIe3M73qKXR5eohS/H7Cs4Tef33T87pHj5CFOmknWw
BPIcESOcvcLs7ekM1oX64Yjtv3NpMmpdgzfgXKnsULCSsH24+8O3UDOYRSok4FkY
yZyAR4noC8uJGtTwB4TKEzavlLYPb8D2ADKmw9msitqXXYv9Gm+WEgFdFTP69LUF
yhbgijltr7IjRYHy9JTWXxjH/slptExnNpOFmaOjsnLbsW69E3TGMA+JBV0lyw6u
rABtyEOGnV8NfQ7febNwshG571ztaury67XLsjd4d8ff1VmJ7JtrBT+11/24xJxd
QhpJXQvhF+oH5oQfsZUCubYfHBIwaX7w7cTYkjJc6BdPseE47L75AucZjpSggCY4
zk8JzvN7oHilKS1PrvCAHIZXFCretY4wdPQe3MOUEMx4dK1hdk/7uRmrKr9siu9l
uxUzRG5D7w8WksSU36ZyxhHwXKb2v/NGp7xjjiLeNE90dgnDsIkx61rekttittHi
mJiAKPtvb3Uv2Gm40DUkLrsXyF0O+lFXeEw3rv35m5/KFUkwCFPfb4Mi2c2A3teg
XqW8DWbW0VqvpbeOaQMrzImY8oX2lESumMm9t2idKWTxx2rGWPh7dxevzmO1ra7C
aEtgTr8Q60Uivm8mMWujYb49iuxnK97aXJZ75XElgd5vtCvfXLKKF7aB0GlNzIqo
egMlRlV4+e+qHSgKTVzUwSNmO6rq0qcGVk8c++NkkzLKLiGevLOftYE6/V8mfbVZ
CdPKY7w6kGWBuvGuuwhFKXUq/BTpeutwMhqWlF+qol4bZBuAxTy9MagKao2LiPSQ
YxbgoT6c5RYnSijNfoabAcP6ubGhe0mlsAUlqPNQKBj+Vh0lpElwla4M70PJDir8
ZVOgu5VFu/w2xvIVkK7GczzVvIp6pUZxsP/wLWoSCtYrzDARe9sBY7Rrt1FI9F9k
1YeCaK7vFBRQThrHqrT0y6kZsiuGIuROX265SpUfNxdNcBaTLH3ZwFK5FEjcE5Wc
keDJR6uwVstqz8X476h4en7TFwFp5hF+VpdUuVlVB26SEupL9uGiiL31KJkxp0LR
RCTBSrrK1R38kZX2ShzVXLKx9LILHfxAyYLzyoBXySFYDbKx9PnbM69bW6j/FQ7b
pLnzyB5ZbOjyTEPtcr/UNO5uEp1UP7CjtH1XZ2pybY0jGGCdBfV05HPwKdZ31pgo
ROMWJo4pPV/HHEiaC72dE+ujhiwz2vQ6fRLoZZMk6KPp01AjlDGckmnuDViRaixn
gBBaWvKM+TS0hFZLsHW0JBliXRY4DtwqLtpFXN0ifZ36qDVVh3Sed16gHKy4s4HT
5+i0aCxjrXk7YMrdnnyvHBUMfxhGN60a+ofV77LoVagQMcWRnwx1Y38tmBHeDrAY
h4GDHxoK/gyDdlkiOlLwgSGJkauItixKuT733z90N6I0suvGICWe4AzXlIJWgXsp
beUfqYkJnXiTCIksxtaDspzd2Rfz5mArizvQl+Wu1UCgVdlmBwV849lmHoX+40ia
ntOwwE1OLu9pYj+IvpjGD949EyTapJAghzuNhMNN5vXhX2f2txSXyQ4bR1eXS6VY
eg55BvuWiCDMzfa1yf39jWV/5HxANQprBzZm7xKgZMYPvTTIX+Y0xakcBjUC57Et
Sv1saiz9oMnp9b7jAKeG5A9D2EFR5f/Pi28MSbytF9GfTSpHRxZ8uVNBaxev7Q2E
Tv8LRGlElkAvDtskOl4bvVZP1Pmt6jyjuS45nccBJcTxwB9aq3YmstP1AGUccsph
n1bWw0EvtB7aXh2asI5Oktm2Rf3rhbjTpTBsqHfIB+X5F99LEEPet7IZCAyg522u
ehzQdBNxsnJ0O8weXS5hrvxxfJub60VCmS+kYO9JJ/BYZOyHHkalAydamiS76qoY
H0UviO9JAsfu3TYWadsVHMTKuwxD2tVHn+DywtnZKMgzMqV2qMMpc/xuW2+s208V
TOMmEUDJU8Zp3JaQ3/2E0EnN4KwwYLMVyiU9YWM/QqdVRZ61JRHYUhpOGm6m/ugq
+o3QjHEi5Pz0n31hWFXwm28dZVK+BVp9p2AST3TQrTLNIp5C7ZvXM6ff+XF6AYTI
Tr0hw9PtnG1CVhvlS3hVJUUCq/OXghzz+dUB8jIu+i3cxzQ+gBLhezVAWT6I8kQ6
vZMtJ4AwYs4bUgGklpdJ4SzV4jue7W7ThI+d8Y9VFJGg8f44YOEszNmWbFTJDWsr
PC0CPZ49qI7CdcCnlORGqS0fwqoqtfrrPyZJ2ydCzO7IzgZFjmlm9ub7MqKX/J9r
/M1Sno+1VpDvViKCajOC9PmP/HsT+GjtJ6w7wDIOpd1iHqQTFR4wqToQMjoKZs7P
ByQ78KbL2j2bufoXBaKCkpSTc+jMcI8/WVoSKAhrFLBYIcFXYUQJyA7v5ZZ2Lq2X
ATN1JTUjsBC4bjoii0GbJDhewnFLdcjSDrMLEJSpbR+RkNQABXaJmGqtKF35Q/He
vQ1wGLOvAl1kTYZLsKBbP0y9Hrrn9ncCI4YZZwK74F6GtN5/JIAitTfoT8334NE6
mnJIkSmrqZHCD2HIdBwPrQF1q6HAs1X1WEu3HXUObl1p+Y2P1A94Nn7tOI3cU/Ou
C0g1mH0yDQS2PZ8N8wgRp3Jl7REx1NPAGq9ZGv6gMl8C1sT1TgOwPE0IidREkuM7
9wrx6LvHiG6nMNfS5Wa3LMaq6rbDJfvB8guMH8RvV/ZQ1E2YkD0ItUyvHjFibkQh
xTURXhYFznDjZGOyNNYL9gLnlsCLEcYRAmgBCRfIHwpntpOGorV8y/jLFhXQEIcA
lDk0+W3oMqv0EnePUybKopCgb5ALl7+VhHY5ppKB75Lw8FCt4YDOHfxurGnUHf8j
5ZdK0Z5Ns6/Shficzmm1bVA/DPLU2TWKo27Qe2y+Rf7T3EMBggSm06Bu4DBtS6pO
l2u2RwbcKZFrKUymC55fAWuJUGoupmrkHm3kFBlzLuWgsi52/bDf5n6LiuNFj9Nv
4GAa4ozgh1BPfQdpJjWoVUSJ/TnLdQ8Wp9hzGgtvyM8TMrn25HdXcch9yTu3N++l
GW67lO6Nb5R90WiWHpNS2UpxzZU8jSkgVvXw3Xey8VFNnD9tQUvR/1OY/GxiVpWC
2s400Jv9iLw62rWDzQF8sw==
`protect END_PROTECTED
