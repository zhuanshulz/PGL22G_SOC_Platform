`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HLMurSweDE3z1q2C/r/NiwfklArO6DWzxS4VTm8J44eXTKnXIO7tkqKWXNhBEnCS
JFur+jE4NfD/SnwuYlEHKAaILsGcOa4ksymve9oktTO6ce34OtO8kFRM0Ld3Ickh
4V4rARYCcM4fKMKL1q4MUTBtIfHeIojM6yraYx3H8lcRlsXfAvg0CPBHwlyyY70h
OqXx1y8doLdmlgBhbRaIHEr4kGzFRzyG1ujGkmiBZCOWJ1/e3g22DeqAQEIguI63
B7B3t5r9r+XZV7Y8x508ngkBFMvH3lxuBb2FpFv9GJWQRAIyyAxJ3uwNV/J/TB75
PGm4ZzbmRXnSieB2+b52zcIwQkxKOjC5JP6u/ncQChpuoisYtAwuRYNbMYHtTINB
FeXJAndxThDZmHl3MiSR8qo7w8MaF3EzsSoI2XgbtuommVK4Dc+HmX0i45sbx3sf
KX0SYpJVOAvRNiHAW74K3JD98ULxCzdhGOcJPeRSQSHBRAqV3zDuV6ou1Nibbe80
a+GUiU4YF2sYAJrJCbbXzuT506sqeQcw170p0ZHcPVaa886CTFnBo4J59IxY2rE3
4AUAVooHPEDtWnAwNw4IRQRfLh+lUQ948QMvuO/AHYV1XyRqlMw0VmV0wb0fmwdK
DskDXxyI9Yd4ASWJcakcFUtmhSuhGEZFWzVqzkdjKMdIsGHCn8yiOAGT91innRKd
GMcnPneRC100cxvTdI3IfkYoh+SIJFhGbq3z0vb/bRUaw/y8+DF4HO4V2XPl995s
2Vy/ssrgyl/cjuchxsxQYkim+y1NwLFEKei/degWhVMMWt/hWARR19W/CwnoOcqI
`protect END_PROTECTED
