`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jK/2ZeGqhr5wR+Z/15G5fUFslh10Rot50IA7/vk43B++fa/drgX/H862VcwiNw3C
wME8hbX5Wr15R91dj5gVO+tCtsDbquksiY/LZfy1ISp/l7SIRFSJVNSjG1LT8QE2
Ldn5fEtB9t6kT8hnhwIgQAHmwdIRWoAMAnQyLxHIAStnxeYEckpui+Px/6cMUgOQ
8a6Zk8xBxLl8hTSUS9kLt5/Koq7uOdv0sB0OZtWbbk5F4ewSwCDpv+HIJZSDGJiC
M93TrgdaZ67Btf9Qccng2o/moHgVOvsCEfVRNaHIrqlHdTlxCt5mBS076lUpfS1/
opF7LSMtzp6+/ZAYnTlDvXqr6UewYOgq3p+UsGmJMfkdfRV+HY6SCuAAXfe7GubT
LVNwluIBS3RXpLHm2GVi3/ppTkj/AGyjvYlpgCR/oMAApc45/oI2G6zb4mW5ZLAy
eYBObMk/W37pI2HbzGeh+x2fzrOZatqznVwrAMzPxr7u7ipA6juazOe/ujq5ev0N
CMlnWf3j3DPNLILinU0JxQUO7phC1Jb7Eqx1GfSsbXbS0GtlItZ5kKkVJr5pPJAt
jnevtLmNUDuHRC7FU0iCExaSn2fof+SsIpCDOjpfwhsAqebqWsp03L2yq/0BSKrz
cFZf2GzyGqujzZy4wfvtnJJtyPNV1O6jZOI9S7YTBtJZemZs1jkAV9ExCJXA0l6R
ExQe9lf994AHLxEf34GM8c+j5IMhnJyJNdC1JN+DETph2vQlkVFVoTacBrm5Fz62
VEuXmWh65WqpnhttKwLIbYY1QOQ9EzLHEDMhAA4y1YaM8McW3c34QNPsYhBZFBK4
AZDMduTTEtUqRdvAYKeuEw8HdMqKYpKO6iD5u7FhdfHHt+cryFm6UBAUjSrGzV4y
O/sntAjl3XhmkhUQtfwsVe8+LMNFvI2fX2OoV1FWXXe6S1bEGeeMHX17Vh2UHh6+
Bif8kurhvuoE7w84w+X8yVYq8dQckOoE8QAoqLGwIvJetzgDRooyfr7vI8JqLqFp
2yzJnmHJSGOic8pL+1kknXjJtElM95KNnZg4qMdy3er1bmfKgeZ1O+B+3+lG23OA
Tpe2z5ZPl9W9Q49/1QSEHFOho0uOUCTtHUY7b59aKE5KhZHi2lIZ5awGp3v+94sC
uTRJNsXyMUdydwa+di4sHCfabBBiCjehD+X0pyXcIw5inZcUBR9wSW1V7aVtAf6q
T3HwwHsWUIlxswKKHpnyP4cTUfLlF7j7uYOA38rPD5HWJozwfgwzgnR+mDU0YbuZ
8RMRe9YNTgUyonJCUtZa04T2+QA9OfCA32u9IsPjwu2LW5YOh0XOr6DPs3ZlMkow
rbfgWOhEtxBSolyne74xeGbZjEg2eUDHHP7S5IvC3c3fEvfOgnUVUf7aC5vxOer1
DfZahoztKpsME4tHCIiibOyQ1fJwrHxaksY58XbPs7Jr97LeLKufJhj7DAE2sNQM
yAZkmI/E1ILxcSYpIgiS/M05UyJon0deRl/0toejl5As3OTqxr1tV4lJ/ZUxZwAG
TIL2AnlpREaBH6mWNmFppCrlhU0wknGJJhCV6tVOnHdJqj8zh/hamVcjUBuyeGyx
h7HMySUI7kj+UDkPdEkS5UeJr5KnE1XLTJ3EmRpqCAQaT+wi3qJzUC6OMFnlSmj/
kb/QlRswBMmiWyTQe9RE63Zr5KExHnOk9LASQfj26+SxArMF73ZxYnWCelKT1m2/
ESnUpnCTByzBrfs50XEzEkEsVVu/l5Fkjw0jVmy1D24OIohSlnwXfh0siRhl0Tkd
JfIRke3JMb7KLOuRtMWZwQ5iRKSs2GWd+dctrVXxTReB6aumVEh92wiRdiMf81AP
+CaaQbKn/a85w/nAXpCl36mHUUvH0aAhmuVYRQ5VYO/UUhK73QvbXsvmhgVa1GEK
hMv15wdeahNJpEzkr0OY4DZAmHOkxZ4UbZ9RCZGZuxc7KzTXipW7MV6Oj3rYOe/d
HV0ERVuUe52KKxalUz/BWxbfOF/ooRUlNTWifRbcR3/bUHfMfHND1k9NhUIMhGFA
hcBTY4JpctsuBH9armfF4phtFx28TGxImoQvl5J/HtMgCH8e5rEzCmwu8nQGtyay
kBLfj2anGRndXm5QuTuKaii40bsOTq1/6rbqmtoZQHqPlFfTuiIF/W2zRypwliT0
qyarRNB2b2vFCEIzvQ/D4UGfrXAJSjI44txGrffJGi+Gl3VmJv/EjcePRujsw+5b
fpTRHpYYRgktkaiqHAFUq9Hz6kp2m4m0h7t5kXLt7q4tXiVS8vrb6HhI3BSaJsDI
ejIeu9Deam6G00GK5BS7VPmkO1QdZ+NZLM6BkOZZ59svJdgM4lgLdljYCZodC3Ag
I6sJHfbkizv0fCXMRzo/5Chj5lnneK6+kQ59aWvA9HA=
`protect END_PROTECTED
