`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xByb8/6bfakzlMb4lJFXIcp60BDkzwlGDoZsrQwos0nKovIo52uH2/pnesyLLoL4
0kdhka2Z8GMy2eOb5YohWdDGvMPIIPkbMzk/7/+ZRDBHyHhTkNeIEYk2K2iG6vMR
CuONazFtVgPBnLtUzTnTbN3JoV06M6iRFt1aF4w2KCb/qSBOZp6pourZlzDjAc49
SpwvS9d7XkLYrX5MeewH8poslVVFmqsP8AbZCJyBVqARhFVbDpfkFDzO7CQBoXiU
5PHgnmGXskovULyVuS1ci6jQqBpeg8D03whUdK7JuqAj7gsVwKy1gC1fcBKkLtAt
TYz4yEuM9WwRIwDnSXpU+ORzRQMa0VihR3srJtfuTLr6nbK2XKMneg6qGIbgumgh
DlF2TkFtBFHuRNQtjnBSbaTma8pULAfWyKGFDRuZBbD4k8NRXz3i5AsqgoKBwsW0
rUaCNBHDPT1/FE+nwrWC3puzBTJ/3T96X65dy20BO0pEwyhQgdGKOafRBPG4SQsk
0slKgQF2pYkCkWZhbhjJUXvj7NcIFsskGXNNVEp+qevqgV1cLmCxhOwCRlgYRwJf
xHRWHaH3qNljc/brrsF52IvSBeB0Oc6W5d3d6UeueCQsdGuol5+9I8p8SasU2L60
IC7NCktgJE5aJECWDUTN2Sf8b4b9Rgr6YX8iPRmN9kdZpXgza2LuEkfF2XdMex0A
4FsHamTwVxGD0eOz0cXPip5NUP1jn5xJ5yTPVWfCiudLXQOOrtTAmC0374iIpcnp
0Otde9x+YWJMjosS0n8669pGkTPO2GeL34FnvPtelkPrjQc34Ro9MFnyLcukXqww
Wp00M/u+Uq31IMvzfPL/ukl/bDmbKWRtrW793wyaUln3rCv9V7uB+g1hAg+R+QBv
iSx7uWGs+HR8X6IBJWGuYnTq1t80Qz5kKGQB2K0u2SUmDAaZMhDidy38ddqGh8ZO
wwJe9gdoEdiNhuZhkZW0Q0sESnOrT0OXaAHanTGsuZ8Yi+3TkgI/8NUYUgFKkRBG
lTGBnU/fMRdC95EnpbvxLLaPWgYKRNrTiQIkD7lo0CLYOM+ANZ2NbhPWwjeN+2v9
7ILzltBqyOYgO2aI4z1Gh3vNdDvK4egE9VWmAnp02iPwYl8OlIWb774F/11J0cSX
jNl8DHQLd29Z39OHSUDuZpfgRwu3yWY0uMYjkK5GiT6FfyMar2ZIlXsiM8eKJTpt
DKNf2NLKGlGr3BwDY2MJjeIeYQIMjNYMFgwH47vqOdRnztOUDSBJek/kvLVHGRxt
qGCTU44klAvTcEJEqRTFpJQi6LKldt7bXaUVH/v4MF4=
`protect END_PROTECTED
