`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U83feVWj285kZGWNdg7Pn9jnAvlF0GkrepINk1Nen/rGdb7F3br89dNtvazPNK0W
1p0/yyOM2tqXwmBvNnN0JPnAfaqsOsujARDe1av+nGkFEXmQK+hw1khm6c/V3+Ap
e1ajvd1Gg+j7PFSzn6ADcPybLuGQfdPdWfHtY14eVLZl04cH0yTUeAPHfPA0rb//
qAI3d/PalTqjtetG/hpX01d6mIZmTf9FSHz16hBq17Dbb2cG4yid2Ycoo9WWmjsU
9jM/vhUWLzHVzOx5a1UcwOcpcxL8eow1QpNWGvi52c3z8gEtfZ2iAMeyLnXYqJBq
fLLndr+IzHijZXp0rITyfIN5RjGO5CM2lVtZwPSCnqqjPmGIw+EkKEaUWizXzkVf
C3ByW0/2y3mnE80eqwMXe562tLE9PWJIv1zy3YiNRFqQohCdvyo1nxtyfLS6dkWh
UPB5cQKmBKeysmBeprArxR42AMy3O3aX5Go9yvQKCym37pF5RRpJzF534oymdS4N
fDmnhZg7LRGkULdso4wfS1QofMgYqCwZ0g6d85luLtueDKLWkp1lF/vFSph1JHu1
mHf+y+gpmTDzYhQZcA53F6z+hj1Li9u4bJ4oYDCveuZCLBLtFbshIj5g/TgaHZGV
H+WRgfEHGSbWi06TDuYUQgcxKEzAUv/JaIWqZ461VKtht0Nfdtm2BcYwuBK4Oo43
+/zz1CTpoEX9BMG82oj2fMY/dMiX5Vx0Hf+zCyDV3gKJa8XOBsa3KTR8DlvNf/qS
r/2gZ7w9Sikj5z0AJDNTNipuuTxuRY9Y2f804iMLDfuUcR79Lz1fX3TY3RiwmW8N
p6C4j2PwqpN0tHHc3pzQgep7ws51EqlwDapj+d5bLnUHFntwE2W0uG/7uw9aL35U
Y6SSENo9Gb6gYUiLKASdr+f3+BVjqjdS4nX4if1XL1BBn+eRRQNNw9SynB9Jlds/
vLly0uZf1VaLYGyWO0fZ6uK1PS9Eqt6Z1MKwW40dDsswmol7QjRyRyXJdImElRRb
XkFHpi071D3pMkzmgihJ5qFJp+I9NcBheeP198IwMD0V4DDlcBxxTrPwjJY8PR4+
jRYKuOAvmXGuRcRS1j9JPTolgSMts9U99b2Nf3WZzkafBGVvQpDh0XcFCKLZmGw0
wiPVZFrEHq1CjhorrQaldf9j+i1jAbCcEt99f+40IoFBw2m6lFD201BrYRDcFy3w
7Ks2Y5vGYq+dm02HEQVTyuD0VCg//N7fgQE271tAfMmrSO+AayJGoFOn86cM6XM1
rhNF9gdY7udSLUSQEbUjBGQzSTOqrzkt3khIjpXZuOBaJ/BFv6ZQKzHTttcjJA6T
xzUCgfLeFbx2QccCaC23ljtAWZgeadcNnnRfVo7gs4apYA9AeQBch934V4J+QEOf
6THfJ0AFneVBG5luSlYbUXMUgQcCu9oe4CQZno2EZHLTOhbn0wGYXlHwQiMx/ioa
NhhVGLXd+Q/LmV7G6Xqj9YoY8gNcFaNHxmw48udmlCjJODJbZyygCrAAJPg7oiwM
weO6ElRd9sT8ZcMcR6RZDaFi9VSlNotmtj0zKtC7P4qxIY9jt+QbIujuhqr3z0re
UMWx/QnKcJF32ZW34M9ZUqQcOwKP+o4QxPcuDfMEaMRfXXU2rIQuBepjvEvwQf8B
PWOVLeUYWuIP6cmy8gpSFWIK6q9wc/QivwrM31i+5NFRwSbVpiz0sXFwFnzON+W2
N0ElsX4DB0JPknuULdAFUXElc8aCIGIRjN5F0lpC42FJkwSwIiZnb7iL82vEb3Ju
dfTxKuLirXSExAnPypGI3D60H16sneyzafA6st6rkjPCVNdsdabw7/ngAtiLfMTE
hJHVY6p1Yv9kr1UFojre0sq9PwIBPFGkniVy9rnQcBMFNrZ7f7nn39ZoOZnAvEEO
wdR99vElHbmuW9TP9+h12UPmKPerSJnU91gMQbVh4TCmGRBFE0NIGoU/PoEBncGf
ux4mpZl54+aWvGAfaUayBPl0VMyilJI9lDlWXq/DdiA9ibCM+cvdOHjjngmKDl6s
RTFYnIqy8zdSv3zwa2jCvnf6KmUIBvxS1KLH55e5sjjF8q8J55iN5pE/0pw8s4O+
JXTu1qQhKzbu+0gOKDW0wrB5lqK0VbElJ4UErr75WyKIb3ACsVehQI03UYxcioXB
uVdBXBf2Zt0dibUqaWSulLE0QU1eFDJs+NnTTX6owbUqUzXtFKnIEoU9mp8LmSuy
rusYrxBtzjYbZ3UkZF4BNARYgyxOJNYuwbebmAm+nbRcjsvvoL9n0CcqV0C0+SSb
SgfzG26ZZo2csLudjqVJjgA3vNHnfsPiaBLeKxbVqURgUpegLsFQhOsZGp+Hw/Ra
tQV40LolG85VVwC7wHgQQJlgOmy5H/d9IZBqFbYnzQmDswBR4s38+5B6a2R5wDut
39LDSmduWIQQ8/204Wr+/52W8wuQLxeUdbWOH67V2D2Ut3xThd+TJ3QG8BWCVnJz
L3oyRDy9MNZuOKG7DD89I2XbmIDNdvxfzB5WJFsidEoF3Fe1zOmAnIMT+XwlAFsv
ZnxoEhBlGuR0bh9mTKr/Utj6VK/OHy0MTu5l6rhPKFYiIowMWI72y+zyntx5rCk2
qYTj3WNPiLBn7nWMHBLxVZBxduAC3qM3UvxieGZ0ABMnNf1XWFS1hmnzU2PMudH4
gIHcDTeur3whMNgBoE3sAcL6QkRilIBbngbRkmIbRStnjs5LN3CaHBYgURrv/mDV
WqBkw38S7Ryf2C1JrH+AHY48b6USdM0ST02ozWYhybDLVhB9Y6g0rm39cfXnWhes
8E32lD7624m22Cn3AfAFejVSjC2gpuRARbssnk1f+mrTCFqOO7HDicysWAZ/DGd9
hv36FMDHlPqCUWnMkbPQla2i0bJ42cQVMIiPHruV2EN61eo8ZRIxHSzLBSa4hNbd
hvR9tJpl0gbdtqWcUTxjM6Ck9Oj2PRi7GbmjJ7rP6ElGz3vi7sJNvh72enGKlap0
Kd2ERyt+ghOnYWkWKQZhumSGuA73DNvIQ35G8MAcFSFC0FCO1oxtpT8Kh4wu/SNu
cgJWzIjnGq6ySL7YI5+zhvO8RlGRsu6ciA90rY+s05XQs+RnZbIaUO/O1EN7XjJu
3z+92cclfTOxzryihI+Prxr53CZ+7Ql+Tlo6LsDC5qZQHiVIpZ79nz3sHdOSNLEg
Q3Hv1rOOhOwK5wlaqy0al/QyJIKcmflNuDNyBCbqieZU5X5zFuBKO9MOVLXGiGK8
OkMVA6yM/mFspN6uqgWA3WHegPI81JOzgdtwYgxIORx5v6G1jvKAssfNiHom+ELJ
DACd7HUm2aGMIHihW9MkyZuEfpqYmBZfNufXT4dZHHuz/OgniNesMGM82ORpIqty
qzhLoB2pIFLx9TIeUGnVSbIGAtglJFwugXKp2NdkG/fby8m6gJ6FTLsuYyBxRvo7
Htw5FNfHe6jUBK2ye9GTYZCzf1GWVUH1V1/PyxV8w8BikgtYa3DW4hLkgUphHC2Y
+x5hEudKN0mnUaVzp4KY6z72bwR5g38k2mZfM+M+2jVTM72Y+pZDg2i7hxCoVvnH
4CivtkyhDktVlg3zUQx3+K74zWrJJGVpLtngmpltJ3I6oGTu9uTCQ8cdaWmNLm8R
Zc3Xnx6bBZ2/+voPSJ21x5++dvx+oQJqBucXc5SViGOORMO3i1IB/uojpINlgq2R
L2w0tTXVNSjV0Jp7h1Cuj3xnn/s2YAU02a/VwVvcN+N2R8hFUtQAJWr8zP1uz786
Fa2sc6VwM7NKkthGeTCMJzYMiHDLYRZbizNtRxOc0HzccK1HT6sU8iKWwAAwZ6zZ
UHnM7jvoqWgnzfXOxNMAPq0MJ9irGp62nDz2Ixr5nKpbtZ0ka8jozO6/ZS3WWr5g
PGokTyC+1oFobb0tRRscSF+gokx5brE+OC/bRBd54G4=
`protect END_PROTECTED
