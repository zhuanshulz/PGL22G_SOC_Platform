`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8sMhKwFs32s8SRI3UYA4FvXXtFObU6YtqG6hZg901zzs+CQKupfX2DXI+fG3FtAF
QE9PTf/2GfDjwXAoNPnN3NBRq1ZAAAIoMn4SIgcYn932o7ndZGRjzhPoTK5Udyi1
dCDkSJvEt4MdcV5YEbEdGBvjuZbkjpx84xvF11lOCA3VdNqcOHiX2bvShKXkN0Gg
KHAK6I4lNM/7czQb/TYUC39rClaEUKGSIfmE0zjm5G4QRfsDc8nstXrVFVG6Jpiu
vh6H3/6iYCYhWX8SzPS7BHBmIk+/wsS/7Fv7stuDeOwc/X+xjfsifXJN8rzeZW9X
WcBNg1fre90JLOypjFCPv7QLoO6Qz0azd7O+SUx1DVCKwh0t75feZkh7Jc+skbPz
MlJs+iDVQYo4gvU6pjqT/gpD5eubgB2tVirdatwGZdRtG8/DqkOgFSH9agd4+lOu
8nOGzpfuw3scS/E+uBE2E6dU/PBqqM9Jvg4eWcBQfUS5fEIJm0Xhzhh9vBCvi6aZ
MjnArjA0vJwwXR9xB6Z/ocFWlaEQzjqVc0H528jiQgD2p416dTU6vrhjoDUGX3rk
HYkA6kw/SDzOyu13eG2VkFCBXl9zoVBl9F2YSwWY5Ek=
`protect END_PROTECTED
