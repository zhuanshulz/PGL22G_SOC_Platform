`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5Ej1kAyN/AU67GGQaqL8D2WUajCL/CUEFi57ppw42Txn5ou7BPSylfZb1igRfb3V
656muHYaBOuKOCt5BZ0lz5WBpqzDJ0a0VZLeD/PF7GG/TamPslO0ye8UjzHPUUxR
P8oAMO5dTc/oX7tFzMtRBjSGmh0RTPVBaAoIPDBhj/mEnZptFecgKj19PNrP7uMs
JbCULO/HydiU97swkkC1ivNXH16wZP/wY8hsmiJNuDwOjI76bgfv/fbNg7lUdGMK
pxERJR1XkUVWOBAT4EX+PQdWs5Rb6Ip5yHkptjLy3iz9GJAWQbyxfWbELAvb2j2b
MBBskhkFD5TpheibFszW4cWbF220ga6KFNijeQ3FhMOeBW1X7O30O8uadaEm5nfD
+N7cSH+LvhUDeJVSQzoZIWKz0zjEiHKh453m+GsqoO0zEg8Imrgj/eyJUt3N0k1m
zY3/YguD262Ku5QTCY0+GqxNSEBcIUKUSejId0I2MPxPmoNGWN6/Y+rnp8soZZeV
FcbOkEF/IamRgITtboR4s2TceC55PpmwtHs8UadFNVxDgh+CCu45Dm2AqOPgY3QB
w1BoXgRP2v4PiSlDTX4LENPtrPY973RP4xe+YBIycZ/83j6vY13VGevUOkOPwEWI
+FMXue30/IdBZ05JbTgfkEz5zWYNMjdQHt/vI2IwmHheaJKBAx6DCdTS37z+Wd/O
BKGQ6ogw9sGpWAWkSl/RcxbRn0YHCCLWXYU4kp5o7H7RUm8O/5+rCVvQrVKRp34/
L4tmhGr6UmoY7gOY7lML31JoZQz8+t7cjet9Uqkscpyww8fP9Dc9uM4WyvHMnPIz
MmRt6ZZdO6esW36w6bW2E3hd74dtSaLQkzST1OM9zF66dm6m69kEN8dlGonn3uVo
/jPU/aUby+Pt/SM4hrl3wNm5G9wgcUptPv33G/XAga3vUGG6dq4yLqUllaTJxhxU
JnNOvIXFcW9OgGe85u5CbT2I2xd1uqeaNcdIgI03Owt32MEpZ5TXKH6c/+vOORf2
sy7NqiWywIgK4aO9uvcIHOeu2bC65OKbUPcC1PxFvh/f5F6VB/0E2M7kcTbK65I4
NpO/sE6moH3AWEhLHz825ZlEkuGTESky0QRuRknUlHF0JZgNGq58citVR92VUbEh
VJ18R+5GiU4XMefAntJK428weFuKrtWpPioUM+Yd59MZi9IYIbAJ7UxwmPIR6tYH
X1UP0EGcQyl6UnRXVV6n2EFRAm21v8pu4MK3gxk130/hY5UCvmATPJV5OAK0p4pz
NNQYk9OboEudQeSP6vdyaXIQXUG6klmVpVoKnC9XVjvXZ+NcMacFBDzjOvLUDBvA
wGK945+spnxu7X9WGkeTMAP3fBasbP9FBaOHm6/Gg7iUXNW7J2UnQJ580bRlh7QB
Vov5ev/L6n2ONxhbqcJ7+Wt5dELRVOShT924SkghicBNaxeMKvt9I1F/t0ivFfrw
qs9FVHMGH+xWfVK5j+YexzdLNDLVhWFnSptdP3Jhm+d4jQSK+kxd+swaGYkoYgzp
HRLrhMhdjQD1dFcLWqcOj2fVh7ZfKI8XUTJ6mfjQmcLzmwz3wfok8qTuYPtTWUjf
DoSWvddws5tb/QIgk1KVuRRXYLhRW5leJoP8yHPuVi2Gdn/WEJuWuizkPxMk6sv8
3xKK7I0p+j2uUOpjJkhkWT+kkxKkoPfhRUePP2Ia+cjaK1bQTh9Tbfm4+B9y+FGo
hELDaOYEQ7yvNgwjOTrcca/9tXbjwaS2FW5c087RIvInMs5ntRWQK6z+ERFP0g1/
AZZiCQARJHcpt6gfpiFLVUF/zJt6PWtBUI98wbEVqfleptugXShnCIz1o5GhstR/
UoTlwJ6wzgQs284hrGEF96MXsnAJ8H+wg+GupZtk6OqppJsig7dEwHzy+Eh6nHBz
AIzPLbrp6aidcWxSYcuDmf9dnlDEc2T904RCVGY3UjrGrGXCifHlxQhbafm8H9l9
x5TIxCPQVFKmKAwkG6plMYeDU7TTiDn7HMpkOBbLkTYyX8FaxFD6gDhzB2+fI+wC
zses+tPOhdARZEn3ADpxI1qD7S3CGjaE5DkD0emyLZeSZJdOxW8/LZYcgmK+T2ES
uVJTKrNp0cW3hWk/N3vleZDKkd5rwquzWRHfKdcz0gFGXoByIsssSFyEyFZl6jK9
y7HPm5W3JCbNzLha/7zapS8y4iDcpc5TJZaQK3HLxq7siJOKDPSd1mBaZoVXmA7g
G+EHhKzCKnBh06Q20LpPE0tH2FjeT34X/wQvHL9L7awsXsQecLXEuOxJXhAJ9QPJ
oV0+8KxArqETkAnC3l2fdm7ENCllTh6qakfZOlLxAVgUl9hIvikencRZePwJytNj
x0D+Z6rBv0SwePFSpeaAEGNq9aSiD3+Xaw2jEV089xIxb/UcnyiNvvmIutW/tdw7
jmymxNoscxIP293PSJc2M4Pg6PKAO001fXt6FtIH4pezEMZFJC++RkVC+1eXz9pw
CJauviSHlyOWwoZewVCn8oaM34bGCuUS+aSaQY4h2eGRgBurO4APveBe2/25OrAC
DyGibGQ2RHVZ7F1jU4b2aVxikkV2kCzOTgq434eeWfDqgZF2lPkDqihh3Yh1dU05
7t01Gf1JHLBhocjYKesZO3TrPcANOErV6PGus73vuliKi3ZnKFczA104xdjZdJWj
P3LETK7s7wioA9y2olpYu6ZDkkPcjn4LcjaCT8Fp6X3Vhj9bMdWnzGajdEH/2tfC
bMN6rMDBuHauOofIOzH7FFjbREtViA+bkZg6/97RSgzvnpMBZ1sSPg2msn4ESofC
QdsLmPGvSxP2DcpzEGMv+pUp7458jKHK90n4ikjq8NFt3fiiNRoy9j6bE8E1EC0V
kzVx1zeNDaNVZax4023h18NfpCXsJI1Y8iYnrFksLPnx0Hoolj4VJGxiyNJ6w5Z8
Wyr+YQjb1w7XL3yBuCJiT5DY5BuM4n72JR8qcKr+BMFUrz8taUmPiv1l2hikLt+s
Uc3AI+LzJ7grLHhavqkvPh8D85wxcwVXFFnNg+cB42eWU8cbXBKkNupW5LZt9fNr
14hlfAfEFJKbgQ8O+7jYMk+Y9p7bShZ2qxDfHKxynDZgKVH5qMHcK2N62ZOsgWL1
abEnWCSC+4+b1W8kxalsQTh0Obn7Yel1p27BwK0m63n+i2H9HR6dS1Dj4q4R99ih
RXf/bQJkyM6wehKDV4yZcsVVCN7VtTuH7NoOrpGtM1I1LNtbYmHOOJXIgavtwGLv
Vm2PjCeSpzkh7QyEuR/gFPmmFscjT/QBCiqXK7tpd+EXKYU86g5xP9JPYvqHyVmW
4wwjTWSdc9qD6J1SetnCyQqtGBcV0SZt6IahY40oXXe72VaAbC4lloxulFXR85dg
TxYqq5flQV36/j0ncFcOo6GWgDimYzLc8Qwv6MBGXIL4HEsO74zoBL+TjP4D+k+F
YPkMunAa/0Ff2MTuzzHPAXtseBdOuE8KAK1rkI1R/B+RSqNSilEGaMa0H7CQ0Opt
UjeDuOAT4+afy/KUnYYyKYIzh1tl8uFxNB6RtGERmudDy+yiXZu+hKWcIu9bViJP
X5GrZFvKJK66WoLX3KKR5hmCfAqzKaw/jgOtk9rdpl1V243gfk6GZFoZLV0lYfMZ
KYQ1LqoxIZ0frGbLnpHMB6NLVkldIbv9hY0GK/h35OUXsEWbS97nN+osoV+2HwYo
JOX6aAJ2ct/PfBrr8PhjKAn0C0+mMYk//syleW5mxtKbYqoBvxhJb/L99IcGDo5B
EQn2Gycn+Ry6B2R7I5umR2fGxAwPfnjT3Qo4ojBqW6ZwOZXdDm4P8cK0qO/4Gc5g
TxyZg8RlHdqcQx2XaTaSS2jKDNcYu1Ins7QCf0NpmPPUG5hWI/7rLof7qPhOuGuQ
7VqGwoujSxRSJAfvNgvALm5cCmmprxkU/ZaF5h5HPgUrVHOAmlfxlspY2DtiMRQJ
aHns3UEBThNGEnVVTv6XP5QctTBR4AraN4GllEy5jbe0XRSfgLbiXh5WTI5KMTMx
3lzblzvR/Tvnft0dNgixu+EZaKXrp/cQTWgJTWFqSdPxC+QAQGuI/rh1sYtxXACg
eNOpKyNzNJxhgMfwvsK6pVjJfKyw0bS7zGH2/vIWk4TxIkj59okh//3joKS1pMcX
J9EQgJI4InFxZgOiPSq+naMXS84S7aM81BpcTaADzmTpPKyKghNGYAvukTq91bLg
zg06wvQIrTLoAoP/ky2IddZRB9visRzeQI8Pdq6HtWftRfCsvUv0L0mqentOeT3K
20Hoer9Tvj7hnWroSyUQdPwZwLBo4kHJi8Cv9DY024ANREF6/cbIHz6CZrDIvm1c
zUdodtFuZHtQSZ3NI6gwlFNLs1pHx+8EwM/iHCOjPT5UPq3AFK/NR4tXLtI71c09
i/2o4jZnh8tAFolswLUKW7keoIwAgn46hWkExh5hNaIFWmbqZiNXwlnX73TrQgui
eiR9n6rY5VF+o4X0/H5WyKveftB+V7g1NV9AkAmffJXGfrQqdlFkMtK5Idd4Vdr/
PyZswncgc2K1OXoDWj44h9EO1vb4z/yoKoleavKeFzigZ3OSyAXkgIjLMvaGTYsO
rb4nCtTIksbq+AjnZBjQsDejUCvzrKlcWh69SSihm0U4j62bSwLB7tTyVRBGV89v
BiCUrAaXMNCg1Lg3AP4Tl0cbwj5M2+OGQcDgbiVcIPq0wuxZ/tel3skrOsUcxBDe
KzlC7k3hapL1tYXYU6aYZG4QilW4IBoF3wOY0aQUwmmn+vNj05c31W02rnYpi58x
HwwODh5/K4wIza9+fqW+qqdmZqdXOxdyB+k6ZfQD0l7cuKuyru/Q573gvciJZONO
Loraq7rJ4lIEEYGZDiyi/oA/KXC85/PyKUrThJXTgRtP3MtLhaenKbBSAcAwxlsg
hBL4Uayy30Ru9cqOLEIgb7zlYazUJPZNPbl7wv/7RhSn+sNC5jxBt3OEvlkuuRvW
DqvvOww9DtnZZmIWC+LpLNaFzld3RRo0puO6Czx1jwuXoKQvHhQuZ/Z6uJ74NBWH
OMQ8sTrcclhg3C5VIJ5ZQ0jFUa0keg0EWZHL80idystqtPMveUtw4UkRFN3/mZyZ
R40nE93lf0KN2ZDehpEgmW7YvN5JwddGEq4Ox6S2XJ6qkaMg1IyYSpmOPm9MhSXS
3iXsK/synqDMmWlqDvetIpF+hqmuTSXlggvJ1pqJNBw+/DSMgz8OiUPketxUgsUQ
+UDTKm8OWcfoQEtNWrAEOHcVCI2TEHotkeSS5AYEEAL+nOq2a6CvVP96852klEnR
ZRTDEEDhFm9LJw3MG0wQSsogOLtXFjvOUp4/V1nQVV5e4KxQoCL/84j2+qogTYHZ
3DwIi2bghZIa90O68O7Dz6cMwErv1nehfdKxOGIZ3JDxXQaCG6DpM6eSXH7ItNFk
K4fLsyqYT9cheEf1IOHh7Li3zFv8l6oprjngGbhPhm2aiScYBUshxsMM3jFQd+SN
6Xyc49RbNmb3Zxis9sGiXMaOu3cDe+LBHKI1sjPu1bKd/8onxtgHl/JQC+NkOvIH
lNz89ppXc+5rLykBz4o0YKHLVitOTOKGEjKrvXfaoC/5whAilLcsQJ4yAIcc8w/m
1CxzBN5VSptphMLdCX+FaPLSdREaTg7q1HfSw6hbTtKB6MjQbUgbEcIPjoPkcW9W
XirDQ6LXrasfXaT8nK0cc8AU/KLFkHH+7kw2h0m9/Y8LBCN0rb43lqLZyiEFTyHM
m9M3OfIb9N6wMv7cu3W1Ia4m0xFXafkJTXQwLd1LOQ3NUuMd+vAHmd2OVfpmvwCs
mOHXLR4AV6Itc4zlpOpFKp2udHu4Ka61WekjfaCnHVJS0CIaFRUyqAEB7BoLNZPm
m0un3zxzWNif9IdMoI70QkfnMrFnAFznY2PQK8VmKMSKYf1zV+UzTipqjUdfIHxk
kOEglksacLudr6+HcMOs43CI+MnRZDDMBp/jc5vhL9JsjojkCc2PPV7/DwGNFezE
tlpZwjJt60lxWXutsL4BrgeclWoVbB7Dm54RgGdbtwmcwbq3TvkUk/1c8STtkR11
CqrGcrgG4wyy2p3p6MA4M+dAOtFwYh2/dCNyMZpBGujptuO7uz1ZtSlY5LGldCax
REzpP49TUvh+FxR+o15ddT7To5sCz2saZI128Vp2keUGkkE0sfc9awWAk+uAFWIj
JmUSGbrz/Vj9WTfRhU5AZjqtkAv1S86G+gWIrSQ/AtIquuQe3++K8YF/wLu3wzr+
iOjzBSQDTCIb3YEAoXz86CUPUhQ6mXW+jw9eUElXNVOKcdWZGaKFh6QWJNJaAgYo
yWzqaJbJt3/0CF8wwvTdMGmpy15TZOX78fPkzAMpfpxrQKif1nrYY8jfT+WuE9sZ
Hecrvoava17LsnkWXAlW/7eyuv9BcYshz8JDLKCMwpLI1QFzKyUR9PUlBL+Z0SaC
aUugP3fJqGUgmdlYQthL0vhPi42MpDi75Zp4cKW3vCLQdzhwZY6lpZ655XXw9gy0
h0+1pMhCZMPdDc/x0SnnO7xBHA16JouTLEBkkxqvHNiL721iZ5y3oPky7Zk9FrVi
a4lSoRJS3ovX7HDQ6uUGKMrwf2tOz2fhoBgVLYGpHcple5YJTKNoRi+J0vqgjw3l
WMqqrW2oF/imHQ7cKrwH2aRggIhutV85o15lGqDdwTI+zSDtlB8oei2PZuBVn9We
i0PyHnYVZByZMeK2FuxMJUg39jwCoWnRui6qvynzfbF2KF6em5742JZ2RODwyxLb
RbwKV/GoiZF41VlAyK87tHN0Ilbr2g+EtPeRbqbeqp5I1hEawlAemgfZXNM67fBV
qfrdz17NWzLgvk8Zl7Zn2Hm5wmKg8jTd3KrZVDe/c26n8Ibmlq8P8AJL9Y40mO9F
AdlmbmmJAPIibKPA1aGHoTUpc9CkahxW5GyUUY+VczSTeyDJre7Sgb/qiG1e7wfb
I/2mx+7/dPEhqDVTQyNeYQz07/7ab89guzhYJSZ2XitYNX1xccLvKxo2Mcox4n8v
Od4nXTb2EE243+ShClLWyk2qf+uOGXmqrcuklADhgXKBxcpyMnR6JSt+i8PENCU9
23wciKgN7uZLDdEM3slggmCsao4sTt/dOf9Nin3EI+YLU6Wu/tdgANSA1T609/Ti
Dgu0f+BeS15wfo05J3KbpmR7zm3SFaA/q07DAwVkbzT99Yty5VwjSxDfF2yvSC9R
rmZLc2N0+CBizwVz06luSO9+RebAmEUVMHvAR82Ks6tLrgf5YRGi/HEfkgD/2mkJ
h039VjtbgYMegthL3kANTtuEPxFkT2YviH+vrQeiW5HBOZokVWEKvFbePC4pjJjj
dsmNcDo0KgGtO6KTXxkL4o77RTKwjdg9t9APYNc3S0Bul9Kmg3OZrnVXfJdbPW/y
ES/COJ8DJt3OA8ShLPoIB1A4mGzGOKArWTHjRBXQEhXIikUloQDtHA4My4+k3pfR
H/Tla4iZaAIReCffz325iy25Et686ncZl45igcb9EAESkJhlqdxxV8btXcShWlcZ
UIVMvWdPZgeEMrwumNumoAXq3JO8GdA/oN/64om7LOGCI4/epXrvZyFMgdWzQfMR
5cnayRLl3hthM6EXhnu2aw==
`protect END_PROTECTED
