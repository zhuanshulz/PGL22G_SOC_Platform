`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u2Ljgf/+UxBra0qwmEg2/4JYATcPtVaYC4DfIhk34N1d7rshbegcYr90+YywljS4
2RJmnAzmMaEZIjDHxIi3cympNa5mHny8uIcsPGs3xsE5uDYW/gPRGmLgYCcfdlD/
+cDjSdE4B9FzyItLOsybD6keiAEI7W0nQEFMM09/5R5PgonLA3e9hirkv2FMiHhT
KPNNdp6APmr/M4qrpmGxaoilr1uVDbGUE8PnFv/4sPUFswqvjNxti9yQWoQcweU2
6dANtZpSE8kHw4DZHGzJCkQMq4h7mf1aSK1AbS0HBZGhkI5wUZi91pIrXG8jLFsv
MusgCKlgnkucIBWCNb7ecftjrLGNq9i30E3yPPmdVgbTTPhFUqCFM2RRGNREH6f/
IDbSnPeWDYC2f0LqMHEG+1A3Q2Ssg1fjNSveFgz5jR4o1iKJqzN+Ke0xaQrtpSXS
rfQzvPwuiBuwsVfGjjHEQXaMPS1zw9VCn4VNGFkWCjr3mnqO9OU2f6hkPSgZ4wUy
FPfQyF2bTCovLm9ZWQYbfJFKwGJA1moV830Jc50+5KgcxuyItZXHmvnD5J6r6FEk
zW+v0H5hrFjpoOaM7fCn1Fy5NFCNtVXekIkya2I7NIlK28riMd9v/rJF4taoBLQy
+w9QKJKY5qmr9KJFI4BRuNWGRETvp64ppgVNy+Lb3nnolFBqRdkO9M5f8rkj4Yyb
ovzWHtYps0E3O2r0O1T5VhC1U4/brHt4/ERHVhN+U7yj82Mv2sAk3MJg6nUW5ucs
qPlGUxEVg07w2PMnLQDmfaLWuwvqBcy0vmNdvr91+z1FScYDp2DPsYpYfSU8GgL0
GpdE/OUANiFJ6M6RaB/aYTr1NPKVbMSIPaghpK2DffgYhM+qg2BNxlJmai8zwfE8
xemyHNEbU3X3VKIpe/q7xKeGNo9QKXVWJIKm3xb//NIpn4P+2j/WnvBv5empIwqu
svgGQuk7dPACwuIHD1JPTCU1IvK+af0AZ/Gn67hUb4NcTaU5C+7D47tIbgGIST59
uiNq/r0S+bzUYmemaf/0pEmKykx445WI6dEQxDznsiVKRsizSAKiRkkoyPqBAjfz
fEH7sWShqBYKJM66DyrxNx30cefGHHfHvTpKd0uAy6FrngCaf9WXil9u0ms3+mOx
bvsLM2hv+U7QkxQ/ImxsTtgN5MsSTg4Hbm+0K6Wk5xQp0SuDpwtjTP52kHs4mxNx
xSndd+vNMc20U+Z1b8COH1yV6ZJtt8ZpVH398p97K6zVGF3rm/JO/NGrSRMBo6m8
ytmpb3r3CEyTvGZbpRx3LKQU9vNfypGGaHHo8+ZWfbXLEbFZowQ4awDElY1f7uu+
ndMtSQefzbMTUtTwg7JoKxd+jZ4n5Zfw1uiaEXGdrUHyr0c/EoG8ltyY7cKDkeki
ZoTZd+ZnC+LjQnRyI19Ds8hix+DglszXhR3moTJaZcniAxEHzPQEEFH9AcLnLMbG
84TQvgyvNU5DujC0stOFrbKL0DkzsNGejM/WGFE6+JEhyrP1+eQyCQ14yRwUTZKt
UJYBbiC3/2Io8Djnykv5/oDww0UdQdwaeeh/0lD0zFyWrFztV07cHdB6bEF5qmhl
cAeGusJXgky+1xYk9nuPS+lgD6lywVWGISTt8V6ZF6q/Vuujxiiwun3E1SkjLjT8
+cWaE+l0UsAtElvlPfo8d/erSKv6f01JLT1aSxByi646Q3ry8QoU3RumxDbCEnUh
aE3q29oYdVcRztOa1jRW6cF54CultveH8LtwosuNWweI2QIDQA3vmMUQltwJWOl4
eMO0adWWHEKDtlg5F1M9Gn+vPbTjsgvjvZTLc5XXcAombE0iGTFSnKHDEShEgG66
nXAQpjJrzLte+k0etVfreBVi1o7EvchbTVMiEs33KDGYw6VtQr7IzPMXymNovDs8
W07BqD0XTRjLC3cQJVChN0RoHkBXPZoWvaWjfZYJ+7hkiHN3DKf030XtFMwbIRG7
dwhF01Hb1S5CLIfYBQsyC6XrEjms/8VYw1tcv5iHflXw0MnFjlFlPixgilUlpiYn
`protect END_PROTECTED
