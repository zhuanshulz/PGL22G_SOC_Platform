`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gxsP3tDdhzH+hlHCGmarsCvzpyWJF4r1juDInKnRtS7N+yv1lsBZVNVoqWBtS1sS
Xt0v6Bmq3zFC32+2jKU+77C2mc0FbAWfi5N2KR7TffVyVl/oWOWpDAvy3GB9qN/P
hJmE0cfbclCgCmrYse2XSXtfEGS2vamN30bc+J+VRbGOkhBfOxRlhMdbEVFxfBUD
OycAnW/TTDkqCpu17U7Qa5Nk74exxlyrZBbVlTWUrq25PYgkEunUb0dQQFiwwBvl
hK/mngqVty1kS84LtusuVknk6QoTJpizWTQoB9CJZXAKLEwdjgSjptCS6sehuara
MUib90/CK6InxispG6HmGBgekyjSIJiV7lZYBY8k3hDfhJMF/ze8U/dZN869Ru+S
YydchTFGT7DkP/y1Oet6CkaXDqqvfNgRHPcfvcQGXzjExGmV92F+R7gUUDiGkl4v
FRQ+nD35/5CfN0W6EtVEQhi+s/+zm5i53sPm2hximDBJMyBqnnuBPOfOqAxN5qmh
mQJxUqrq13g/W/LKeGde224fPtaxvU62yUIGi+BXNGwouRXAy/UF2cXABhND6wcP
oGzihRtxXWWuPh9kjYldTcMcevO8/L6vb8B7x+j8ONbbbDELUM/KhM+ntc6D6zfK
qf3FvIrNpk0m5K7C5rYYK4qzKvxPCk8GzMyDFspQlkzNfQhs31DM0IGLPHyUkbQo
EFXe1/iUEC88isAb+2C8SFMUkGLY6I2x2iPdITyzjr8PsT1Upmsq8DVtwOUSRR8h
UErL8mfuwOQ17dzAHzdyLMa07j9NpWQ6orDptUFcwsA50YoMmQyED0qG+ac8TJFn
75trpZoU3OjfaK0MLhhBijQxS1vABcYfXbY6hZ8XKaYANE8pRJffuKaQq4pN09jy
ggnf3P1nRt3kLFf8wTV0id8USU97YLBMG3oD6aeSRO03OTYStZKleHcdeumqPao2
HkTru+xxTg9h/91XcDHwbplb+o5aIiblgZbWo3JRztMODlrwbOdb1ugyMrTMFZDg
zxOOb10QuAU1ZBdADVrqE2m4Fp4QuBji2ex6eLPHiz8yFajuwmx8x4AN+1lXLG52
1S0AX7ctZIxcmv43fqsl1hfJUrF70TqKXpeTIxfcmDC8UdRIBn0g8CgC/FKW3zfj
yKT9OmaQBKEZWX48YNnEI0rvaHLO30XEoLJauvE7+ltA18+j9Zt5yg/LtAxWldA1
3797o80JV5Tbr07H7Fu3it0wa9oJJYoOFz8NcshAtcabyQ56YGoRK1auc0eK67ge
m7aY3L4IOQkrSC2hX709MSdDIS195VG1gxOxtUJtIH0b42bnLU4p6TsDoGWNg9zD
sb0Wg2T8v1JwuxJfYTCaHMlsvidpEZdCMQIX6XBCiG9HfF5cAjK0yCnRW3jyo1wo
WA2h2cFjen6HtyF+OGft6v1C3KH9hdHDqN5h3J4buSEwNuLZypUu351Yjci7asMu
U56qD/uFzXb7LTdPs3dPt3E9ON3v/P3Qm6anbewqhe1TKscbnYmXVFWc6/bpXTKB
MnRXWmGF3TX5qcuS1CD1NoxRAuk1HL8wGzGamKDdLHmKJS21W+y+IE7R24Y75udX
YuQqBw8m4A/6Y7RwiUt4AuhOOzitswkBUDB4AV0XbwXU0H8tDeArgbXDNu23V+Yw
mbbxVfP7KSiQj6QWqvbGUo4cAX70h5iJGbz6XOzyfg8ZLu+9HFHZ0tVxMgwkb9S/
ye8O7WysB5DVBStK0MdkhlMnUYPEl9kPKfg2SkIU/H8gUBjE86EIMU8Mfq6OdPy6
aHnw6pQy+3bA9090DxUYahzk1qH+75RlASQxPpH3oMzF6WPacn4lWa5/PQZdIipU
Z3fTtzP39LQpSJbGJUefRV1oo5msVnSYGdE/v6ygWDLHLJ2aFdRcQfUEZdTEFblX
8jvg0qGqtB5JQyR1Ri8Ciu7XC0PLazHQkqqdFMrNrOlehIvSxeoks8LJxwNuNSmO
sRxY+/LIddO+YdD/kgYIKiBuYDOQc6bbqmQm3CrO4+QYgVlSjPPSozTIno+sEGX0
Pz719tWfXpsEra/+tJ8loYbUnQqOrN9Ogi2VdOZgKANcGGvV/28g3y2YcMWCM/PR
qGRM8w7OwAOm4xbFnXC+Spsbg2W+YPgDCnjuWnz1cy70jSdHWJUaonL3/8stOzXO
BNdUnaDKqLJoVz0EE6+nr5BRVGMyih6HMZHh/axedY626matUaXLPHCLocQz6TJL
78fNFOVpyus56yj+SvKQ9IVwhc76ZISIjwaK6FCx+fnr09jmgqHdeBdgI9wSr2WD
kDz2yctjPIvqLXt/tJ7ZCTHeSPxBQ6ZH8qKTmNO0W3pR8eNmsI3ef5pMdcKTUcCb
NdNkXxjKvH7+aTLuTx6u0I46bgmeMXEqhluNddhDl2dEvFA1L98DAPTeTJilWRpu
x69sIFGKTWUyG7dz31Zxwhq1aH5jQ1+kTSPPErgsvWNokQviAEQjs4W5v5ngVscx
/bc7ps4l1hrLjWq+CoAaiDXBVfDFPj/ueEiOKxwsVSLr/OUkjCpTjP3PPgx7UNIf
QrkTBdTsLa5frDvIszcUEpugPJFIavU39mdyJp16WWm/OY60HOdTFcSEHctOl/i9
mE7LejU4y3V/dVCYAuVvP12WkpYNe28W9JMj9SJaqi0p4bL4J7hR+RsslwGgD/6v
xJrBPXbc4Bzo8UMsVNfNF4cB520WViPbXSKXGFN0RP0QVCJCLxFu0B0N91TYWMh9
03hDFqoz/44xHRokCzeHUP8PNx9AGNQKN3I27a8m6LVlRpPdAiW3X2Mfb2as1MkO
5RU8v+Emal/DD7ISUee/bQlHbtXkDOL2ZUHTgYmzMvX7wYixl4s35DAZcUc2b3PP
JU4Xo2AJiK4PhJ2KzQGKCMB70LsPmTzQgmyY0aRNOj+1LbtokWx3x7BhR8kTfLWT
j1q59udgmuCDs7TKiD77C/yY7vjEK1KD/dd8vsACSHzORrHJGCUYsKVkibypBPYm
tncK9Axsmo/3o7lx17uo3o2zpyTQ4prnmjVRyl/4jZzFfzq+s3PI+yq2JVtvvAgp
cCZzuYnAkoMIu/o9mta9p+PtWyZFCHWI7ww2xzib/Xwz38R2IHmGdlSTOITFV7lD
nH8bPina6EjCZ35rK1KuRs3tfZQN0wZd9QASMbroR1PzTDUD08Rg6YMQGeRAcZ1F
2bw7ADXXAqM0xHH2wNLlMjVLr+tjToKol62E6JwRAki8khZKDLpekQtj4sekgztS
6t2EXlkORfRmif0F5U+cINk0Y0GQZIeOBlvbS3reHmoo/YxR4629OLJ7L9P/ObzQ
B3Cn6LtoRvmAzrhswPP1TGOVaeT4wzNeMZParPqMxVLEgI/yVc7C3RRz50QF3BEt
Bm/a5bVhlOFEDKokq9YdfSmsQrqXJuEnhmfjTaNehMqiJ42hicmPIcaMbwIrby30
wNfVB9mMh7hZ/mwDu4j/+Jz1AaFmpMSlv2qOnAMarOeLnkQcKtn1K7KUAEmeeekK
luz9o5X2UFAquWJYoQzFAeVRqq7+PSETNpFfnhP48F0LyPLpaobbCIzxX7i2GEef
`protect END_PROTECTED
