`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HX22V+Ad1EJ4snpl0UGVWyl17LFobrHo6dAQwAntcAKjDpWbKtdMv3DyueLlBsVr
5g661/dI1J8PEyVHhpnNHlWjnu5W4daiwQ30i4OkKfu1/SpuzxWiCuZ2+A7qHHxa
gFLWWTp+EUGJ9rR15gcVy8xvNFh8Den7haXM7xlWCpP9S7P3WNIfuX1Yhg4oPj7N
GLTdqNH7Vdu30BMQE3A4QeQ+4sGzQRd0j/O80nSIyGGpOm8BOZAMLX4RWw/YTMhd
EpY8T30js/1PQsCb4P3abarCFaDBV0EAFfQ9GU5QFyjB0lbeNhV5N1VjzFEEEyGA
XhnOtNA9+XEmOelHL9+TU+zOELZbIVlWgOGlJnV9Ph9ffBSSaoeETw6BL9A7o1Ov
o7AT6hnYu/udZmOvHAtUCV4oOLwj75mRYxUDoA11gDvfREsciBTW9Te7AcUIPhoZ
JwyGmw9Yl6wKJHh+t4rlWYZyojKTHQYVjGU+y/O0liJiwGs2ToXLhL1fCiYAlrU/
IK6cRf3G41uBNYOiyLfgkkIgGurrErXC+AJd7r89IjSL9or5XbyPmHHLlH3wbDZp
I3kPfu0U/Yzh4oFJ6dEnS8vsTFN5rShZsav20WxYt+3OKWNVpaYNMUbSVMju+URq
YsOw+Vw4Wj8NhMSwv25w4cuKVccP0QLbOohlMYwuVW6EVt3mH0uDSlaL/78kSWdn
zpJ5WwD53R3TpdYYJmhiYgZta3n+Kys1GIvD0V8vcp6xeg+MEx/Q0Kv/QMgXtt7K
3qSsWNdG5WnOBdDhTQ3zpv/XUYo+ovXn9OdD0YvRy7zc+nHrZeXYJmNBLtHygoYp
bXSGo4qICXVhv3jpwW+nXt6tC9nCozhomFty5XSfUlsceJ2mqCuC9xFxb6dKL2MR
bC8uzh3m7TK7fDKiq/SlKsnUsnYqKqzgWCqy8EzxhkxsKs1eLv9OrACrGxjvR5RF
4rCl8ucTLmBT2xwD5itxmrM7/HC5L9Xd01KqRlmjOti1NNd9gKppscqobBD1umKE
xsBtKkrYjgV9ZAZpJWcQltLpCsi5dmtfRjk0Tn94bXrwjK8C1L/bLI8uvjXAlqI5
7X81zTC17dZx336E6UB5paQcBZguJD89NmEt3oO9gRbbojqUdjVn7c5X26Z5C8Cx
XHzPp1GiVGOSYDCR9RHBEAYPD/8BTyVKp1zWE6OSRj1S7k3YbpLYbf2QmQEvAkua
ZD+rMlzgGS4Lk31VUijuglCDv1hLVicPGrPbsppn0kTS70C5LikhO6UmCmP0uLqQ
+6s3p7GRIo5tkGe25C3zMBh3Vrqz5myJaDD+JoVBJmBp5BGASshbOgYjScCGbiDk
EYB7X0OR3n5ED4y2uiVq+/3Lz3HPlwlGl3EAmt8e6bihMyUbWlQjYujivubG51Be
HQIx5Ia6Y9AnOm5w8+GoPLtGOUkv8C7W1rYOax3L+NJRRBin9ipF1V0SNd5Nggu9
ufonaTi7MhnSOHmAlyqjjjPO+CULpZpF4cwmS5BgnkfsYxuLt97m18vNpnhQHgZ+
eVElmckAvEpqgsEz2d+wiRLaboBlfLcz7r8VvALSDymCMGxDn4UcUhk1joOc6IH/
pXDBly5h0G2kOZCrCPbnGPnL1FBP5LtWPAJdoDpyzjVH1tdVHBGev4nMdfC+l8ax
Ml48pT9ZahhKYpbZHyVfI7bdK37cNLfWGzzSoeBf8NtHyejfT2TE6WL/A0jcvhFh
dfrvFoAiE09kFWq2q6rYJ88/JT4YiNNpX1y3i1JBG1wTyggkqNF2mihfNTjigrRQ
V60tVjrAhXMqEYumbM7EOtnsh7Ut1UvU01P1XFXRIOi42vubrVERliZo18oLYRHM
X4KeRLMg+BrmfqFP22nnF8/fQOhTK7fxUJMcE5K+UEPKBjOVh7KDoktw4qDcRMNy
v1FwI8NYJ/DhEEhgc4umyR+d0NxXoduJK1jNs+K23igkjFdKZ/ajxE8y+mz3oOh/
6a5f0fxbBVtKmzCQgA7AXmN2A4aQjTlJVe3uSCiglvImx8FUdHqZjkCSNy6yYoaL
ZWkqAv+84cFA0ZwSwp7/aqDGdLH0q9o/A0LduZtV5FG0EXiEGdFOOE6rpXoIRZcn
381XCH5PPOkjUgu8pJ4J/cXi/5eK/qUzoj/0fZeefN6CZ/7+TAhMAuqSOkVtzptl
`protect END_PROTECTED
