`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cv3fVU3FBWpSu9pk4+wIn7fLGnfnTqiSsz4DRy/Roe5m6Dp5v/Oue3UhmAKuym3b
DKC3SdlM6Cp4gWrfzPgYxBn06bHQtRytDk0fk7zFljUZYFSJL5DmfiOsh+ZmplLz
XQOVSgQPxL+H2BPAzZBAJfcOEYwaL4o9k63w+id7dqBBtTcpkGvrs/mtL9L5ClGf
Iap6j7r05h2mVPp1OxJNozrepwFbTFQgAX2w4f1YZM1RXR9dyKWji94xTmOXg9/r
h+uVLakD0Fp24Z1NXPQtvseP8F8bp8zAvrTWz71rj0VNJhZ9fQaqyhV0eK4+OwLm
2IaP0yxx4ujWU2txyLjCs4nMar4Rmq6NHs3VPAzmcPtHyXbw5geW1B4QkB4ssqIu
VPpnc+zkyu67sHrHIivvc5KhpYk1kXT1ekAqhWqz4m/+Fq5eWruTwe5yRv0cEMiq
yYDT05OZD2r+Xsmzyv+4ehoQ9zG/2rx1sBKitTQZmveL7tLpBbfk8ywuO7klERFw
nwBX4Z8Ss/nszQLPP7U+6S+vpWgPblZhun86p86p6/1m9tbSVMxQkMPqf65TeHjx
RrCLCVymFTYIHtkBHX/pT2AQVpSXrDILq+Un8Sx/AxubnXHudYThqZ3zvroP9GjB
xEyVOq1fSiUuqEAfHUvU1KcIck+LNJtSXqRTDpJKN1iyUXhmlV29GEoVfsTPfXwj
KM+pxjCAdIP3SI5skCtJ6RRPohJPPxBKxvcNU+24bEdmEweJi/g5aKi/tYia6CLO
gbpLQMfznEfyjid5tDhp2nQjvsbvLuRSSloXUgCYAiTSYiQOapQG0761/ar1+eim
lg+Ifo4PRz6hKF0i7kTJqKkaqJkZjRdTTZ74pUFLEA4XbZXOjQ22Fvt2/1v0FlD8
5gvu7/hY6ll7nG66EDItovkLdYhQZNxlPUkDd2T2nnGDAwNry/rj8iN5KyimoVmh
qNSFmV1DiqgRdRCpnMuNJrTFnr/hNukz9NgkFpZkSk5wbS7MNM/XS2PBunBVdMvX
gKdppu6eeDWOP4mTG+BsBbF3UVwSv8nB2mm83LebRGjfHYA3vhCugmJSYd/43HVZ
rGmjHJMRfZuuGdMHeZ8/oKlGB0EthLhWWXFMGnNgt5Qsm99VgcRjLN0Gz74KeGof
idD7Xr2344rNZO3PPYh/2BhQR53mkhiXT0F1SoPVvULFkKHP3qTay6OQEDgjAmnF
Ef4g9Zi7lDWKw3Xa0qgx1AOCBPQnw+0znvNyud2e38esXxLeO2z7zSEcpPGDshTp
0kEPDOoifBoIt1w+Hx6keZRlTe74OtBxsEEWrmQ7iIJ7+MsgLMxYn4kRCQHeRiRW
o/kUvZV4HTx382bx3xDP0cIZQKP7I97VzWzZd05ev0L71r4cI3IffwhxEHR4P51p
G2SuVuaOnrMznkVTb178zxwLWL4uRW0b8o3F5mdEYueBKVFMr71IkEBsVw/AG9I0
3Kbn4Q834ar8VRdMXUN1bCa6aEgixsdwST1dNoDCgUvJUx/FrxX20LGixD3kaVBQ
XxAwLWT5rFB3ds/gHRH3jK6TJ9UpE/sjxEsbcf5KAnFKs4leG+/PeTFNfpziGLW6
bPteQ+a9JH6pkh8J+uXfF7bICU0F8Tg6mrWxrlihAxGK1+nzWSlebWG9eBnBrI/q
bXW8fsKXQuu/VqtNX7VmW34M/mE4DCu7rMTb5Zhl4USRNiMnsZ8ivClkBzFmWOqg
d2Bw0RT/n3ccCvwr7JdwgkSv0KgqdAQKJZlLMbaP85F/k8xljKTVVOO/zYc94wuu
JKWF8oBAUaI/lJ0vug7RxJ0YNLZmPUYlqGcLO+jLR9gCMOgwwIrVtTG8GRl0+CRf
9JmEc4PLFUtF6HC62BkXZM+5W9rP2/e9y0dyi113Q2B7MD2f59++F9bk7qQPegUg
TrwPJrFDvZwIO60+1LGZvXfXc60ZjMjdUMP8bY5DdFoUL1eqBw5jQGnGaDvpmsck
q6IYuQLzvHS+g1558gGI2ObAYzK/EUTYL1AohMtzUFu9HzUN+txqlYaqwAtIA1Fl
g6Ax59jA6ZzRau8uS0nJOXUzWqUCDbCclBeT6qPHGm20FJEdoooysI2Tt8diYtqb
LmaGnVN6lCTW2P4vphA+YUmuMDT2/NSVObaCFh4ZytcLw41UalrshK2ZFl4VT9PT
HiM//PF81VlWRdkTt3LbVw==
`protect END_PROTECTED
