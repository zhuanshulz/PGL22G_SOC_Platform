`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A5Cv+lfCT4E+7/7fmPfgXiSqXQf7QqZ+5vxOx1vX+wFK3J6xZUyiLw/iGdO2viJn
glc86wZjalx6LTbWYbMDmfS13Nuc+bX1Ek+WW3xK5PyH9WVDILfFOZvHndo1v5sq
IhRopU5s8hH4AqWTYXSmBjRmCz9M/8BXp3fuW8jh/2bN57o1/b4gWLbCAmQG3El0
1p/kR9Y4eV91pszmYBV+Drc4D4n3bnaX2p/W3nyd1mk/SCnJCi+4HQ8oG0pS5HQe
C5sDyb7qTzCDYhKH2jg9tIT2Z5jOkHELJCSZhaDCmOgZlgpp0e4uZYHEe8oOBF57
qWjK4+5gAhS9pODhmCITm5Xgyj/vn76F7DyEUIY1prjxGYXqiTNbxVlLjItYDZ+t
HwY8d0c9ovKtEfSK6VKA6G8pFI9/2ntWSAdgEZ4aKxSfbW2jA21kUS9xZow6nje/
ROO23LDS+M1T0DoHTxvmTfVdAfXTzm4fAJfDmd44vO/Po8UBqx+BylPvBVde8tZ/
mYwYM684NJsOuM9TQi68q6DEVz5D7EIH+UJKCzMp1cLIQEwUsSaeI7Wo3rt23ZyZ
CAAIsbU72NahRH3bsHI19It5r5YGeri0WPrcQzG/WgbGn6U1BYJsrRR+HsVGXGFq
AgBeWfUoTd9XjPGW7MqS65jND8/Y4qVV/ipAP2t22gFd4ikS+GkeV6FRtnuN5jYB
Sg5G05sXmojGo/oClRK+Jw0+mAD9Ph4ljeo6ft1P7tquNXHU8k2emGjZp7OMkwFp
mJxPmV9vgGcIhAIsCHU3SeonUqfSv1HuoSaKnwP/j7K+p+PWJbdEGf5hYl5gd4AJ
iIV7pu5QEJMfefHIEmZE92W3tNHdM1DSuezuOVjGuSesbtWQOj9F4+dFXvyMQZ6f
KRrxsGqN1/u99qt+E5Nm4arqHk/inp1ioZwMVQFNOWzjoJ/ZpplMc3ZFHN3KAJhp
v8tQeUCUDY7AdC4XN+qjKMNDBsFBkBQN4VAcyjH8XIiGomORO4f7j0aLeJv2KRnA
EYb4bd7+BXaq/REXnLCE3cNpySpm8LSOS0HXcFGkmZGRG2x4q/wNv0eIBGSbpn3s
DpDVS+LGpH6Cd0cy5FK0tsbMTVMCo4uwI9WpHpmd88IfYKGI560EvtqudYQABJ8c
N414JPGh+HlkCWVL1Ud98mFRvKcqpEQtqelgGbIFGiNPfjzorH3XKT7oEUZP2QuZ
UBR4OkWPItJBJpQKIPLrUNwVzBYsbTo/nJzP+ONEbdmmpyW8Y8/lBPkN9IpRvn5R
Fw/nGfe/cjN21ZLPdFbMd8Y331xurdePrjeGWx7sKw/j/A06hO/XOFufA82/GEkQ
VO3GXWnoWET70WWvembrV2W3JgiFk3hJsE5wLwwjGVK34NIG+EL6kBGidMiqDpSG
QnV0ex+LAVq/BrYX8D1F3rukZFFcubn6UU4lsccp391taXvy8DTfjJEH0Z+dnBvD
fFn/VyYyZwi/Mh5/2XcVo3X4WkqpyD5aReUiMeBcenPLEBa2q6f9MOVdTXmZW0OR
YrdPLjiik8Mpw/q94ePXE+SwXi20qIbz3WjLn0MEwao95lfbbp3oP0itT82nIUTD
xdG3QvXKjbzWmzfcWSiOAWR7sAH3FcXFLqR1fA29BH7uY/v37GDLNVPYSl2pDRSo
LvB0oEhSCaIcw/UynCWc/cJmfszTLrUaqtqiKpLX0cfGnhlfi0/msWzVP6xcOA8y
ofY465s4GsT07vg52f/xflnxrWNvNw9cQRH4GShLfo7T4lhjb0B5lQvndxenm23a
lJZViA+siSfbuv/WJ0ld5PIrcBBtidRrWaNemg+76nPOt2yu72gKu3DsrMVrQxMl
MGQQXaacmTRpyNbFmI36Lf83+SqXkZTV56BQr3LxhJ1MEggtbZQD4B0dcHfc92Lr
oExGr6QwUKt3NB+P5Le1FFyQ/oseLWbPyfUW/sW2D2zX92f/g77jthODO2QGZyWY
U83DV4vRczW0rRbxZyrPXHjhN09hYCVYfE47FLbwvsrode76y8YntRJBfwhCFrbe
DFBBhxf5aespHklQJT4U47xT/CYV77g7JQPY67yVLU2b40LDHCUOerfen2LsWzoV
XMwk7AFybeLUtC4W4PnJKgk7ZZ+a9YVXxSDrlZWhOX5im2cwY19khj77s+yK8PDS
vzQwwIZwwwwNm5i7jObYh3bswE8ut/wdKmkJRCs5SB4x7fPZF4a3sw+xfkD81pJX
+lOE10bpdSFuAB0F99RDgQ/fEipojXUeh3yVMYxXOMmuK2Ie4zbxVameC3R4+iTz
av0J5wrm+qKcUIovhj7qUvJrkpwoiYa4gDjVDYEfxBp0pvtA0rCN5cPeoxETANWS
qrxAoLm898Z12oMGYQplUnaPNRiiksyfv0J6iR94mK9lJzG7mD4aiol7Y8xxE8rN
t39nV/CgqDlwx8f7Hozom+zdjOdsEVKdypknC6fIB3lLR7yc6u4ukPknIzHHrfCP
Lqj8so1Y8XI9Z6jN/JHrWZyYsPUfIsXakHlBgw5E0XgrK35hMpXI3g0pEsNHTE7N
pYfXLL1X/vahtnBE0CabtR5x5Klc39XZE10e930YCtJYKyAQqKXasAqjw4NbiOLS
grj4+et5bPJQdzgBrVbG/zP6x+xgSqBM1Iph2ut0fHUMY+S44mN32TepsX358IiC
k1+fJYTwIqk/czRMCPZL+Bqk/L9wvDQIW2G15oHcpbozje8shcnIqo4OmixwVUfX
noOwwRSH7nerSaAHJjppjzmnzEUymKaupvufaRYhzeADbXNzsICFCJ2kuoUutHrj
FkNUoY1l2T1xkq1J5es1W71J4AnhQYoaKmbyO7/KhjO/tdwzbjr8VQVbeQ+6NL9g
NW/uULT8CiH/dKLmvymtQQOv/ARJ86CV7CgPfaBeuWJ9oej6XYf6MJZljGI+GYUx
Cm7Km0wTfLDlTrMf96JC8w==
`protect END_PROTECTED
