`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
INyOURLIaoks3CmUvKvqSyDdxNwZ/hKegyPH8USRm60USacNJqzXUH0yoGOgIbh5
uvuSjeAKJZfkbT20g4SQocXYNqEEDCxzBzTNqqMo1QC0XHGPWMf4WBm/bQSZaavZ
p9wj7OKNuEU4vD3M6Cj9yhDD2PZ9I44FovjL5hWNVi8CuEA9F4+7zK55G9k42Tqk
wNgc2p+2AFMEH/Vzy9FYkDdqrD4kV2yTJ3SQoLUVnyn6ylXBlGedjxxZuLBjzZce
B5B78/Et27+EWWJUsFoAd4VKe6jHHeUbC7uygj224fh2i2h9G2TCXliosUvTbcrm
LPS8E8UwQUd25n55deikWxCCJztycnWuHs8QwFRahJn4i3o+8cIwN2Ra+ibS7PUM
jc70TLuMHCEIOGOyMGy94SD1GmyP5B4UgA6mbDmkqETnnlJwMA1PfWjb0+PEs8n6
7WJnJRy4XEenm0iR8I2E8/uqqel6TSNSdf+PFyTkiLmilTGoBClHRKyZzZvLXomP
3pcBDXndTNkV2OgxF/28GsyR4KEA/+FtRXH49WD+Ox9eS2zD70zGjyikYiFcYSje
XtIFEPgznyb7TghB8mfey64LiXS3LT61t/thlkEsKbWthZR3gtb33Xd2wEz4rs0c
L/FCFmeFNqpu7K8L/ll1Zl8jS2TzZ0ZCBnj+2uCkxv2FcF9xFCNGFUPGSn7F5K/L
GclqbgNHeO9AAuxbvAX7bDJRIJitsopsM7Je/2rDHUWo0R/Ff7wA+XVHpNsmJB4d
WsVaboT1DMNJAGTNq1cbUVYNxQlADHScg58rpsMj0T1ZN2rD1NZ2dcFd/9pmL63H
abgNLxOxOqTxZLAhWgAHS/qaiHVKgvlWJgLytND4DC/3TPpGC2178J8bn2ZtI6bh
wJVSs80sGYyr3toE5qI+P3zSLEcsZKmIrY8nUAcu/hLupnjc393P2pNE6LwlbPEp
vtKwoJhG69ppWpqBBjVMeH4XtgMCPNVr7k54p3r35DjyfQsC5sVmP9FpV7w3CFBJ
NuovSXIlXl0T1683qHbiocqKShXefcbj/s7m6LJffhPfshwEIpp7mErHFIVlRfk5
Q+vqAQXqi2SSF+fYQ+24rZmWz3Rs0qwp9zRrsk6ncG/QtW5gldFgd2MRtjejzthD
YkfcmQ3hDIKgXS1TNr60HMvBPxUml3mBB7FIkXPLWNFexM6JtV0axJdy82qJtmfM
NDtFlh+WPXwHZdC5XrKV2laTKbLsIsPQ3NVL5nuoBqMcG00D6Ta4BDHjFJ3Un/s3
`protect END_PROTECTED
