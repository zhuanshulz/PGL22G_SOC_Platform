`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G788ZIx05YLm1D0CQsDL4wbhzMHjw1GjFTVoaAW85XOQSyTdOb0zEdUCdpBE9FhY
WrqSwOOOkLeP4nXvqqr4FbCoNmMPNYwS0GRY1oQdY734Bc6gr9yD6FvCmD+uAxrW
Txw8eVs2+VpO1k/nKMBM+pqC3AOpvQbpCTSwbqZZA9MFi1ritaEzvErkAYWe2tol
9omckznyozpfAxZks+SVRJhqSMRTW0AMmR1djN6VF7TcD4WoTn2GPbtIzeKdxFyL
tTYoqTe9zjjiHdmgvQ8mwPSyJNjfyoI0qtnwqZ32Yh0hnD4Y2V1Ly2rps+TKoCjL
9z0+G3YTjpAz0Mbs3y1mBlc7s/L5cX9U0Laxv6zsXHISjxZdUnyAgeAERYQA5Ike
6ZmuimQPO3gShfHjT5gcCsqcZsP6+2B2v4fjtFcw4I/G2gKsGlf6+wqrB6kWxwvR
aovD2GaCoNtPQCTQy/YUw+loW+VNArYUukW+q1AEaUXsAdHUeu5LLkZsqmFvslxD
fURuF6gVh511kKKnGpuC3RiYlWaUXiLsprLwfAKCSgRoQlMJCYjBewSW39NP9Dsk
FKrmqFsMJ37AngRMBXLeI2++5wDwfZeOGMSlNci0avQgjJgF+6uqln1xsjqckszi
e2l5lcAaTXNSkHiANOzRMaoZWhvGWTJa3p6iC27k22Z6xoCBDn7e3quVkIKv8eGf
3JtDA32/GPa9iRB5pytMUTP7GKYwkFQl8ygeDkVBS3nwrzlrzIhA1/UDZ0TN4oie
DeRy+4GM2f9K4Ry6x6g0R/XoOahWirW2WPQXXvHGOe5HtrCVBFIVri6MShYmHMB4
54Xff2YC/XrTvBjw3T0VOX3ptpaUOxlU1gqlkGpbnokR7EsHJHjfkkwF6c1yZyGR
wzMV7TJw2PysM4V5FcHwiMtHxUiMmraY8Us6lrXDdUelTqvRVc4dNJHbBASIaeoT
WD0BpbHhIKbidMTA9pHu2UNOARlKSob1sc5q7VDQek59/QPUFuVBC5pdkmV9b53U
BRoQjXkU68pCbGl2snjdSgWXeSG/5kEU1A994r/jJKDw6mVTfySLoaQa6UinCwBr
JK9ntvbYzcFMND3x36blJao+ZRbSVMc9060TlVvIiJeziZojImww8XJLl2sJoPnU
ye/f11ifEoar6BJOeU90YVAwbTCD7LfFqVywoZIyv4+uENxiD9RIECPkOkms6/Iu
SWx7wGGJQ450qmhip7+ymyN5Pa5QzCfDug4Gy936QvZYCU3KOKWvP62y6zzRT2oj
rY6rKTtHvh0gVWGlhbldZRRzrPBHbffwexDuBhhY0xZsy2GWXlI89eW7XXjncSMR
RrQxjnlAeP1NV0fmC3OkJl5K0RInz1LsHMM1nlVKIwr3ol8VtfmbFf5FLhs2lC4c
9vZ3hx3k+5tDR7PxcFfybubeyIM2OTZmxLPnsrdGZtko62hQR4IxC1m8zOcD1oRU
R1y/4L6MiktT6TyjOKa6DiovHnufpiwSjwM+Hqj8SqcwImdJBJgP4ms96X+z4UNe
sG2PYOCSbXmgpYyikkuruCz/kg+dSmjiFdbGqLhgXQuC5yivRvARmnOKGS/VUXAJ
uLwd6CyMEjMRkVKX5gp+7bmv3hpx+0esEQXhRn4vlGv7RLS4IhvcWXYsGEpz1YX4
9a+V7ukmv52XG39Aw2hQU2ZAvJb381u4xNod8E4O1h8rlohWC7QbsvHYwa9rpZaB
Ds2wnbzrJLItQJa30pCQtD+VSCDAMGlxdL1Z/I/X5hGGpOqgU9/4Fw+ikuVNiY6i
nR1kfFiTv7lwg4ko25MH7YPxxzOXKBKNcMfgd31/g6/6LlhplQXs3qad6BriBXVq
XuXdV6oKRWuL9kEo7eqXLmJyqPPf39KwtY/l6cdi02OHu+RWXtJ9FDf2HN24qW69
dSUh2BDOi5VY//vATBcynoQ0aPQydsXS/o80u+NVnYvnS/h0TPjQm1oKd/DLiyY+
3Xf2jVDXlbw/sLhNZOhjCP+clqQvQvreiKXDk/gVnGJnTafeniWFzKaYRu3UrB5+
fKzIWebfkqoXNjexkPbkYdsYEZnoeH06b7tFijW6io6DAXRuNZn8EFps2SvEE3ou
gpD7lZx8nBC7T5FRobOF3JYiuNhTX0LObiWUEWiNdas12i0byHD5qhZJG3za2mCX
RuRadsq0EU4pYmL6pvXRoizdvOzctZhtHGX/BwHMQWdZ4VM0hIiXQYqGiXODQV9g
GguxdCqfLh0hoCGF1RaNWMFdDAR3KKSWIzSqllFRFLggNbGPoTEiy2UYRlJa7IGv
ZqElvWrbTEWXv0t68sfC2/xgQor2lNTefxxYSPMo+rZ4CqNUsh9Kbyf5cB24CeEu
UTNp27Aj1/fPBtOiTv4Gq62rTZ1eCtE4oA7h45ZRfQ6hMADz4+NmNt9w6MxBAFjn
Kz0KkfnN/ZEYsH8f+GxhpOxdrINunptGS1BqqAlieNjE0MR9uAd4QNpJUWNYITJX
9aoj89NLDNdRsNa7P0YEcXher91N01lTyw60NAFniOvABRqMig1sdABA25zOb8SO
1FZ5z6tVT05HuqIMU7USCAGmVv4TssK1vPbscTPEQHpoX7P4G6yZMtTUy1Y0GC2c
oEpRSkU3AAWzSNTtPyFFm579p8JyblgeFLtbcxnPyPGuMFNAiEizaN0JbWeVz24N
jDWhrTrvwihZwBQ4bVFdaIQ8wVGmaB615ssgdPPoicXU+kmLrTnawlyZvT+CBFIt
fQy6vwS/aGhNqpSBYL/wpFFw+5icT56IrLYY8uX+f5J0+agxuTUJEGWTDaoJ6pof
3Xdo3nPU+3FEnC3SRMsEddW64oZiYsdJcxLxCF3iKwejYDXYWdvwEyIWVKVe3fd8
i3nqNVPqfRNQatRp8NqqVoLPk1xxUYTH6xS1L+TgKQeYnCWUf2nO/SmMphY2cWij
ye3++uwrAQ5sZYDRhekzxcRB7f0y48WqxwVlzHKpstn4ewllzPJU+RWQCbMfq8OQ
i/MMqZ6P7pHNg8mDO2X0n4MBak8BBdNuniCo5g50m5PJrF7fM0NGqaSo3/rxAX2y
LyMfbaLjnCazAwRq1aOxB/LKZuoqI7+353w9KHBSXwC27hOVShCLgHPic+/5VBV8
EHUFxEhCoxKwH007N5S8Bm0rFczbyZKCB1t7xBpPXzxDFFBwzbCYhbufumnz9XDv
nh888IVTUXqQaiquE5/gML9oJy73nM8mc5bWK2CNkjeV60P5O2NqFWidHK07hkt6
xSu+ydHqX0FFyFp1x2IzHZzGl1GC/Ok2nq/oPZqvmwgwS5NXmC/ccVI7lJ10SMas
KjzRKGlm7mTdiD2M12NTfFSCchsFxyqSuQ9FzyiLPJHiOgP6gJXeDmqoCoOdL4Lm
YigRl3cBX7RgoOsfiPG0d/zM0WzLwLq6jbHM37x6TOxYW5EvLQ+jCC+ZtlB5Ky6a
fVp4K9t9lJNL0nH1Yg01B+0liik5zCGJFYXn766dTZ9rUkiWX0V7lbPuqAHOZoV/
`protect END_PROTECTED
