`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lOpZPzxIqU14lhsZpUW1roH7WWT3FZQ2/LfWwLZ9G9g+SO99vQO4bfgH9Tok64pI
mOklIy1iZ5Gd84wNemgOwbKBmqSS7qfa/qO5YAXEDZDcu8RcamoMhugsZ5fjpPTD
28qOqnu1zEUVwb3I9f0jCdzdZMGirIbbU7LOKMpMuIBdlcryPCsbCzu5S0KxloZl
PT+zY6BS+04XxW/oQ0fZmzRJKOYCWUQlTG6YwrkIxMBDlDWxrW6YvBOZcEWNhB5T
o1hGl6K2rSR+Qt5jQbAlJKlPec7Kk/SNYDi9C7lk9PykT/4j8Shh48x4s3GKs6vK
2RTznJuoRlU70gffB09p55MJPaoGqouicIUHuy/NGs270bpmdYUph8cuuNK0Xey5
fEpgHGVa1JubBfNyA8fBxkIcgl0fHKSMTYlgAUWB5bnezGFLU8PmhO+5/M7NBM7g
dZxYzWKdjb4lZoY0BGHYB1K6yWGlbLnruH+as4mQCekv8uLh71KmeukzP/htJhuz
+TxJ3wvr6P0eUqx6+nDS5bfchLywRbPzlmLzQK1CBjDjsoR9k2Fs8IohLUVf1FoF
aiQ8arlxLUh8q0TVPvXa/fVkBRSooAedG0z1wiFWYoMjaWCkg015jy3LSqr5IeGn
JsYaqxlA4ZfVGDKZBmBJGHbf1oUe3/SRusJYqE/2M6tID1MSQtunDeb6oUTH88Vy
UYWzPohA86QxqJgo6gt+x2wiDcumgVeAUewurVXrcSGEZAAWH1Y25dqSd+mh5mMN
qXkq4ySAJDlQDQfasFFrKd5uMXu/F606expkqOgq125XQPqLmeQUY6V/kR2h2dse
oKcYCoercRLw1sqhqpM5wxMDah1B+5F/ksGWcAXCYtQC1p/Cw3pJ7l8VjVXslsND
I3s7mv9X4C+ZtQ4OQhF0GXOQ2j9btgHDp2ezF9oOyKXzJ/abvnK1YRP6n/EukAA9
ziqkv7ullOZx8j+/yGHTJz3hVrbLDwb39WiFtwwd0bIb2F+b0XLVWPxY9YWSDRZI
1OibjBRrDSdDdqfeso80VEuLkRx8Agn+YsO+t4bnzZu5QIXiYNv5QgC02wH15JFe
jfTaLvozc7cJCxeWLx+h5ukk+op7aHqjrHyMxNb3OU7REnRipK906+QRhcouhTmF
ccVt6Lt7VQFwj5fGc8VbcS9rCetsTDuMBX4E3OBabtu4iukvvMnmtQaVgYnXsyHe
vXtl+/NLdIHFLcFyi2MdmTJ3p60c5Is4++cTLBfuXiNmgk2U5q2C0srBVWAFDyme
VK8+QmsoNtqZ4s2ZF21U+cxY6Dc1e9TH6vQwRfwSxgkD0JhdWi8BN9xiOLz1HcoQ
EUo66o3hhRtPEvQYRAZKd5afwiaxPY44ZcS2R+SRY6R/tvYGioxCiCmRU/BaLLyp
rVx4Pz6njNrdzyn4dPlYIg==
`protect END_PROTECTED
