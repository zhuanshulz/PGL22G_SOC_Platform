`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nTgj/gZr+6B14JSURaKA/J5wAoJWON5IuLQHA6WTMVLeJvLE8ZFolVFfx6LcSlpu
GJoSNJW0GuSLAWi0I+cDiT2Es1jWDn7uPOd/wH7VPl3KBjkKoad1YFeRuEDWHoRG
our+0uz1jCC250AoQibFZl/m0l429lRfQi8x07ZnoIOjDuG3WrFWVKS4aZvW5D1d
uMrrcwtZUY74NrRDkJBvkV9kzUuj88Ushf82zUlUetrZGJIaokDxS84bQFrT1hLJ
vkQGkvEeJBzD5A3ghB5F88dAShA1DZmPW1YRCq+3qLxhNajLlLKcITctL6R2OMy1
/eH6x4qIjweCP9E8DTRFmM8Vh7p9F7pirA2d84BJ/T8ydw17dfitEe+r+MzjZeAi
Ll0YulOQwaikcMSLSQLoZUskDQil6n1GdpQfwW02uza9ELp7tWlTT4oRIc9yCa+l
lHrcM6hTvXrjs/ivylCWewnSTOwEi/xmxXY9K1VHQ0YWxwcaBue4ZTXFbjq3Gnk6
0cSmO9m4VKKnjByCiMRXifOHBPPxK/D7G9HNlVmb26c9FGpD+lKi+I0cSZUY4Bkj
OnRi5AnAEfCyt1gww9pAWjs7g8B+klhZFLvC1zlNqkktDrflBes73Ibp3ufDf24B
icP6N0m7w1dzMXT9AW+0ovIamZXl/MI9S0VmLJkcKyFMdFxGcaP/69Bhl+ax9QHd
GnBmPazW7WWbyw5qSVsInZM34CWlr+o2buC3MRfQUHl/S2RgxFfIUSOliPTiIrR+
TCXr8qRkgJKN2RMP66nzdQQPADCL1PmGNZSNKV21vNQ1DkfDWSYhHdOG5Io6pzfC
9T5VB2uqMknZDrkhSjDyHklQAkJ3Jru5vHqUm1yUyziPTtePv2tu6TC2rW7Qe6GJ
bODnyPwihlUdPJSIiYiPMKH14UA0PXqYA4QpDh8/xXD+1BzBJG3Pbkti50FULPrz
phKIL/7H9PrrqAVaN44BTF2bjP4PUXPDvHxK7bzGWjzZjt7BCAPkrIQHyKsixWHZ
2sHkGfv5usAbhG3++RZ2H622qyNHxulUGyLL8Rzvif4FtaHZ5UJaRBYpM5yLxYVu
S0dQ9O37LLchEfGW4DhIrzCPXQqqZZ80cESmqX6InZit/Cx4VqHoy8b/rnWXqWYy
vqW6iKVdd74aqQaIqqGz5rUvzKsYWoDwHCmL+HcpCEonYhqZwokSRSGq/LJdR3VE
NcLzXKGd//IcyBDeDsuIPaavLrII7r7j4wb+sJylEJ61XEaMQdrlb/SfW2JdH/eX
x0Qt7u2NwblwBeLY1OyZjkqteqiD/4JrjkUFk1bEn+VYihwpUqfOm33AKeXpLDIj
gb7LPe5pKILd4igXTVVUnG6I+EznJ/W4OStjyr6T15CCn6EPpmyuAwsRmMqpfdHc
8U6a9VoIpaUG3X3CyRzUYAmTOc1bIc4YyHIwV7S6R/1lsQr+ch6jZE1XBVB2S80B
gaQmb+7hKfSePDtTEqL43bEasFwFw0DQyMnP4F2vL1MC24JHOtShumvB1DQsaL3t
Hy/1aM6rgAdsDdHPkMtICAJr5DdAjSqwUcloDLOAnpTHe77XqTDoPWLL1I8ORYLc
WYVPqSN0g8e/s95+HCwhDQpYlD9g8a7mQbbXRGorPj9pUBq1CqVNa73CvRJrOUvz
FkZtJ5SzRQCqq/fdljzFgY+KMWXlQxav/09qVXGgeI9OTroDvdhKDCqoCVnw0vO+
DPNWa+OuvGicxIHw447Ll0b0cymXyBzCKu5S74bkkbNHHIuD5K4jBT+/p9yFn9XD
z+BMtnY+mnBFjtfgxg2R+3RwK5I4bH5GgqVIFTAPyV9OgoNYmRUD5WxtpgROoFSg
IgTpdFWUe60mu9BAgsFT4Lbuyk6t2Yx1I3bXJhpXaKEdmoqCiMcCDGK4CE5pGpMi
/4m7xfoZBEOlnmR1HnqtXNbPCEeBIhwaUkpAZDeBiW8GZoiD7L2zOZAiwXilaD6w
VmXrGILVD9qqcMgkXe/9vY3SwfgURIJ8pqeAeYLUoTgEzbNHwLEUG929V779K4f1
SuthfMN25PtYvvNbymNC0ia8JmV/YnKIiz32FzsADb06on88qzc7Pol8YqTvXAgC
iS87Sem785OcpBPFRCGtu8T3R51NLE4S3bKX/X5l9wuj3SVFXyxhiekw1XNP+ifH
erj6tfxY7hb/QdXrsefoQ9CCigOHa5EZDybO9wbFWicIdviIJCgvwoPHGDrgzg6T
WBou/PU8OLyoKnoKHNS16g6rPzVPxHo/BlQsGXKDU6AsVF53m9+VWocnqQ4/KqLv
JTFDyTKKhgxAVPtHOeVk/VHS3QbgsDxuk/o5GfkReSFGEAwSboD0wXE4EUYcUF3v
SXaKxYr0LjYLiyg3AEmY04Mws23vdHd9nyqV0xzBd4qRakNW22RA5IrzuPZn+H/F
L2Ay7P0CqGBU0iqtB7sgJFjdGyRy96u9wZgOq+JQDvR6s0Sl9I1hy3WeGccQ/zbe
gV1bj0Ob3aFN6a6nYEVOmDkTyV3E3h9QgGBfwggR8VNacgxHUe8LLazbUvODRe0j
G9gVhzafZ6eXMIE9bPOIvVexzDwWfV/u14TtQtJlJnmqQZSADhjCbr+m6ZaN6xt/
whVjriUnYzzPYljPbqq+3LnHzdhpR3+nVzi3Kn2V06IrdmUcIDEmq9kEMkUq+uVS
OiapIWObw9BHTf1Uwt3loBtE+3H7XUTweS6ensvFHzTpT/jlMzNu6S217B/XthbI
nhIonfDujndHq9AHdl0mBiyotzk+1aNuOpkaqSPXhwaMs1WhKjYNLvPIZn2YtQHY
XxR1HkmQ5npPp5zaN2ig0RD47TwexytY+xAuOdQ+hGCxan/1ryOuKqVu/mj/tcKq
U+45xvPgDMc09bhs5PT9HRQt9WnhWyBXnO9a7BsjaD9Gd3vd0L1NbKlVjsZOGA3Y
dEJike/+KtRE8qAfD08U5KyEQoWAIeEYooH+1xPLXR2tYPlUfSd2I4S5YcRkicdz
ouBYrQkA1LHI5msTl/Y3WzIjJSncAM38xOuXXtXEPsIKzLyLY2zX2xu6GIviDVbh
EfDjkYLrUNHYUWwcYGmDa6pir+uxKdrGmMf7mmC/pRZxYp8cCezmwe+/KP0R6vdr
LBtm0Vgtifx4lW0TuYsLyToCe8ZcuXfCaKPZfACGrseaDWW0Bwk89sF4Aa7zN/PA
erDpMDw3v2PHKh9sGiDQL1k6rDCC9rvkfL8fXYDmU5DjbMu62f7X+MgJvlkSzHJT
vBnhGb8TQtPl9/zW96raBKf5tOJSrR7fxu65JCqrEptj8fDFwmrli6LQp2U4k2D8
W2ty7JCIZwBFSg3NMzjSe94dmLqtYcv5OXcTBTZdCDEL/ZHwXh7ZbQODH1M0P+G9
9BT9ymem6HT4vNW9JEwpdFhzkyKyH2209gz2r6JGPRkx4Gf1WWrarmHS5Llb/rd7
YgMO9nEpYxNaoqfYnp7JhJMI7N5VH1mO+Dst+AR4FldYZpUcVE407nQX1W/FIIUe
zNJ3ongHY99Y1SvI24vYFk572YcVQKE9x1KIGPf3Ah2qUMRhfAAfHZnMfoYYkSV0
XAG3NAadWHrsXRpaqFuKzkPqj6s1Sm+K98D77gvFyAeu3X2NYncchysg1Fg7ADjg
Dm3nkk9VqiB6IPPDHpcVxU/caaWrWWhPMZnmqVEF5FaR6EBAECFoeoC7CncNAKQd
S2JHFZI8iYh58W0eIb3gzZ+WetJ4lrBJcAFk4CrK2tRmscqxKwe7vZG0cHH5v24K
+Sc2eqOk75pt/9PNseNMd7RhbGUr4isc6jP9LOGnx5vfIp7eZ91HUtsIT+369dGO
gUe+U5LwJgmxKI7sfK1vB3nD6yjbXEr5B89FOool3rE55WZ+AD1wlpGXioFuMc9K
W4WT3ogHLBbJ0gQ0I5VBpqen9OEtgQazjFUJU3LrYQAbURAdUAj2uKRek2KKrGOk
Wa+zz/L0NSaRWMGTp+k+PZOZJOdjw49dIBCWppmqCxhVX45kSrG1GzIhJ+nsdMVt
vSw+U/87ShZ9nqX1+IC0GuQtn/5e3TtcNYlSWIKbnm0FwbpYbT/2N4T0/IJ2zBSU
4Vqe/eWhIM8Ged8AEDAQBS13EW9LseRKJMWluoo1Ayq/yc/6C/UoLP4N2CKz81KI
XvU3TETQRqbewYqUC0UIYQ6YeP7ISq0nmECJ60XurhibXJhgOIWIYW/IiP7//v2E
roBkEmz7B0he6BbkvnsruZcgMTb8/Kv+ELDJ+414cpSjw4Ipp6vvKJsnTAokF6E5
4Nut61Kj5NHHkB48pLSn//1fenNkGTWV4HmslO6Xv9rxOdvi/V6SRNaa/yIFgGxe
ir/0A7B9OKytEdYSCy/BllT3r41Rzu1Jmuk15sOhK7U5AEj94r5BnYLvTKABRgfq
Aa38rNcIdynkln5HSPCyk4K5hNmOeKakQa0Ld3iukTrOM1kRuGbOt5HDIcsDIcvj
ZatftFue3iITlok/ihnkum49a64kuoPUXzzthk/EE7+7pee7E1x6Hc9oCyrsF2jT
7fwEu63LqyNm55/7KnfMxggit+jSA7Rz76FHXb8AIn3xNPV2swtlU4JvOm6Q5KP5
xEj6RSgKjm7Jp4YupH5iGEoRM4SmpM9wo+xTSUwKlMyTYiom0vAkyER3fCCC4JFM
Jl7FQ4iEAyG5IyN7t1bQXVko7tlbpB8ly1mbKJfttt4LurOQEVJ5uli75qeaCa3E
WAIazLBn8OAeBYaskuOFRwc6ZysnA1l6lhf+MGKwz63sdUB39i712Nfn4UzFl91d
FhB5MB0tP+JqBDxp/cHWnUh6sQEQx4q+lfDpFc2cxxe/WAuWgClGpUYom1cc5uj/
STY+27Ss5X+De4+rJlVCYLPGH61SSPXwxJAbrwMgjOg1Jd2b1OFCkGWJHyK4V+ZP
G9ML8YOPw5+XQhW4cWTmEBw/fQ1mL4TI4/9cmnI5rMRAAozlEq4OuPtFyfkUL7ld
UrKZrsQUuSOi8J0EePgZ2Ua+n5ms01sXjgxvdAr4pbU/xcB02hU/TrsAPrEAJZ01
U5/sr08/uXz6T3WzSZz0v8lvdsD0LqzF3fA49K73UUlJMlhgrecN2DRASBAvDGLy
sOHj/4DcP1gXz+XCEMKS/jFoFfoamezx9AA/IZIE4fSfWegsk7PTaB+4BKyenMGS
NZEZRKsYpazC8ZhrclZx0uGolA8c4j9ZS1TRaL/DVwQFNAgBL2r/m/kXdTDu/qN2
ikj6xibtpiFkuzmTluKC7W5GXp7pJV1VODKtvYIwNNcNBeLVzFtWbuqKLQl+6HOh
QyNh30nk2R+A+xYdJcfgxbhkY+WiUpCFApCeP5V20JbDgSBfqmNKXt8B2bwInrUd
RFTd/+KZheFImFRVLs8aM6SE9zfn0NNT3/YydnTZJvBgb2sHWJ8vwI9S/0RquM4j
t0YoSX/J0x+zIDZtbrdPKxGeI0KMqAJEk9D4fIHNY6pgw7PHyviygzE+WvRM2j85
M7k4Y4KoK0XpWheTNyNOaJWltYUP+ofMppZy7VcykIuY94CYFu374RTnjUfixaFX
cH3ttWd8NVt1cX0ZYntq/Zvc2Lx9hLtV1nzBBSHzvjdArp7LNIhyg55NS1VPZe4L
KTG2PheQGrTwbBqFkEXCzW3inRCEBjmCNB2Criip4MukdhvrlhKkqIiMknDk5cbW
nmVIG8blspwgrDZZKa1nbmN/3M+MGf4Ji0RvOKfDmBTT8peb6kuQj0341sEMXbhu
2hVM3iHPPjTIlC/LoQ86YeqkH69YghJiYM3PmqbjaxFlaGdIDZWjBfUuCTCmGFfU
V4NPO1yQSSqhxMcADld0RXp3v+vETUYgl4c3jLH1v4p0g4m07Z5C4pKbBxDK+xay
IKRQzwa/KiSIlYXzq6PiTZfkzBAeEOBpju21JX0cd8rqHdoyWDY0Hc5VgBwskY4t
6u9O9IdCbKFv1XTgEcNoW9MbgFmyr4RlTPBv8XKe709/93ocm0HGWxSn4QQGUzf2
4746Yt1BbZWhV5tPDdnskHhoghEFy/8rCSVaR8ZLMyaPsFVn9tghJo2ceCTe9vDG
yIXP19aAN3aOzmNy9xuUB1wWOFlpVpOPUQ+JbjNahz+Qm5c8YlzR0G5D8xN4duGM
ydR12NwMXj2E50rW4pKcHnY/231ouVJ5jlS/tB+8gupZlruOdZpDgFQdyRKBqu98
BruS6DN9hg9Lw7AiOsRFKeWwJWGPjtBubG30IsQW9CzK2GbkXDCHmHuffkQsVrsH
NC9DWkoR8JKcqMwd7rYpF0IsWRH9+435lfiXq0z1DW3wuPib499LJMpcqM6O3kdL
cEfwpBqVuyke+Ut1W8UKEWbZC+I+x3wYXAOo52zPb7X5VDmtF57YfxXh898m13Tv
nab0ir7AlzIrtFI9sc3A7An1FSSLkHGYk/1TLY1tXx/XhzdEXkg2Zs6mHn04OVm/
wlQmQ58iHWQUaLWHyM1onibI9j9uu/UUvkT7KFQzP9Dhg97vMr0+lVWmnOk4dTRl
dh0OaBs+WK4ELk1+kYbm0VIkjz46fgggKc2kmk6i58NE0vU/FHiHmEpcCMiOYuya
ubNF43Mx06q/umLvAv7IhQjTB9DpLi9WF2uVc60sYXGxGT/ITQFu8pNRNRwK0Iiw
yIHRBwV2uWCXosFICZJPHOTotHS4FVWVnsKfVjZwOsfTS5kfWVBWxgoJHquvnvJw
u9OZvH7d/eYBNRGz9lMoic6FqY/LjRP1+ao7LOFoWOS4iCVPyNhWftiQGAnlUte/
NL+iuN1OAb0npqC0UVGWa0sAdColSqvBPDNbV4DBMXAy7BbdwNGj9ZUqt2d7RrTg
rP/a50rSe8l3yfEwIRNdCa46J8qnGuDjsYknc/Vbcx09K1oY6fK9el2FP0Z1BPFL
qe4eQh+aQCT8MKGS629kW2j0+FfO55x+gzHWMZ9ejWSq55Qygv/HLMCjsckQucq0
1jdwWa1ZAiBIxd7hO4ceGdniAs8tQttbwaqhNO5CX7UmHqvAKo/NBXiWX7g6vo3j
m0yjN2pUcFRqg+RUtCoGDcM4VYBSopGuGZPxmCNZqVjeq9XijhGXFvsP/SjXOa2n
EfjMtK8gmN4H0BN4H5OazMJ472mHqZ5nLxw0Mfz350tf92jRvGHF+mJAcGPabie4
9zozw+ooJVxc+Dec1cmD5RUGZt8aD06Us4gu8tRP8dpJy+9vNFXlIbtw/+AY8eq2
Qmfi8rgoWTEa7UtboWoXk/I/xlaTMUcK1VFFGZ5GaueeTgVwj8LVZAFgeUqflj6X
l1UlSaHkDTJiRx5JB/Jk/fj/p79oyNrYql0WPC+elgHr2ME/wQEJy3dQImFmegIF
llKR8yuJiZPuh9xPyO5fI5waAywI2VzEi+1psyF1O4HjKQS3FsqCmeubOWKDKJgM
/BYWlpoXRJnVnjF+3meK9Hy0g/eM2o0f2/6DxFv6RDFU65okE/QsrkEorMh+tqKH
fQ1NIRVSWW59mLMvsdq6IvAW4MkDhiUNAqXDhnEH/fYY4X163H0LMFggKCWsEyLA
DOA49YtVH5ts5yI60VGPYlEY8xx4x2m3zxYpq29H5grLYI+GGup/aYHQezzJ0JPi
Y4qsCbJAt2mhuxBAqwW0Pz5O8Heck64DZZbdu1KidfSE4ebZ3ZxHYYr3lkfKWrh0
GoBLGOtxWQFz59Dv4V8bvPdauuOygjVnYRBjCjD/gHet6cBlTry0Pvi3zVlnahZm
Bu2bZ+PPufsP3qQ3KiOEiXYgiepTkx5DSuNn/ChqOmuQ2g0XDCeZ0i7CK6ex625m
l0LizlEQ3Xs33++Y6WIVh1fgbvAB2VLiSFLcXlHrqFeIhHBf2K0q9FWRp/nAqkpM
RiaG7qmIMUYu01b6nwUqj3RBMBwRdH662TfL986zMEpInneqj2mvb0Te6LLJ9nIV
OGZJBl6oc7LURd/DX0Qb08WJA4tYnwvrapqXh7GItC6NrBdl/ZEA44qpVVQd/Hvt
9f002TwXxT5ETeipBmbrcCArgVto+WTucn7v3LesHvWli0Vq/GwTzPcXz/QHhghZ
BDnbSWbloTIev7+YGs0q0HVqJcwbPCvcyRX/PihIhF5DWs4az0ys0d3Xjfq5rPG1
VGJYW29gpbZMSysl7STIFCy398ZMlu4yMVnrzy+A73yrSu00Xo5lHvexTraXhkZo
0MiWS8/paCstFnnDsZswkW45p+AzsdzikcZr3jlspThu53aQm/fqjYBlo5paJOUR
6wZWpIFIx2QC62Wt5RVSZkkNP1K5WXDfxAltxYDjINXAgBPLQm/dnMmkWV2mAVki
ShaFIC8kDI00mfBTKdM8BbeY5IlKP3YWXi/F12m+zfx9RhhwC/eGvOE83w5TwfHY
gMHtOW+qysEkyN63TX202G/5XjPJYxybZVMkpXbjeKeFsweg6dR8mb8Mtr5mCjrN
/ze85ZE6dEXbVqrLPIt47p9FvPQDfAtZWsTJJXxPNonGm/gPxPKET09KU/AaQtlx
dSS5EnNBlT7wDXKLdmWvbjyFhUn7q3ubbKiJodganj27EnFpIwYftIw7BVfaaYNT
w25hHSG8A3C90zFd6CMwt34CU3Glo8RvLJJBCBwj1E7f5t6yskNE+5POU3eBrrkS
ayLyV/vZRMRDcQj+MwDK8oO3+IYA9AzCUwp3QTzddlGvXKdkdVlJ0TDqdxEbSZDU
AosXgfjfTQuRXJxmBjk7sY6C4eIEXSDGsT7C0RQ1f08xID4ydhE7FNk+R3+foQgF
he0Oo/uFX2az5C1OzBA4T1RQxQZ+DE9NBaryjx5PiEDz4mPYRNM6IISlKjYtZmBp
nvSPlqemfK0NbgbZgyBtOIa5iTmk/JdLwKgBOoUQZdA98AtwIacXClA8WSRzaJzE
jEB2oNn3YOXSuDRkVryvUs6PWnGrCyhIuAYaFC0C5TrOIBjQR+1lWihQF5qjGUX6
AWxO/vjMUE3wjGWhdAYtPE+nfi+mGRhJi+UhnKw2l0T7k1gA3qQhaaI5MA3hkV5V
2M1o69dARzbjYUTc9woYLIxtiQOz3/0SuRw1m24+jVrA5n7zKFbtIxGkw1HiBxc/
dEMTGDkXPx2M9M/u6RaNIOrIdPusov5rhVk6ypPpAHZQMOgmGmdwm3SflaFVR4iy
NmY0jeah6EG+SKH5pJMtXP2LD8ku1g3nfqlCV8Q2SeEpYnhOMSlMgW4QI5DLxAkj
vSvYO40N2F5+yaPUJlpO7E4ZyTsoKwVHDQ4Mpv4OPwHLyvaOrIPHrs5yEaWKBZZ5
Ge/kdtDw3QeQs7Ybv+xLqN/5ZaJ9dIoi72GuEjD0coK2SkEOjsdALtnVdxThlIvL
yY9rVT/ocvIry6z9uljpNg2SWwK994EECGzPFKkisnCiVFrWcnIhoWXD6lEBViPA
w/3T6iXTwv4l8C0q5sXCa7TJeDlkPH3uHr52DcPLP76wdnWsJQChmY5gzbspXPmu
EmSuRQGlHVb+P8FrGEBrVSiSOQ4qnSIMM+UrtBd/R75692j39yAPg0Nxfrgp1S8Y
mjSmts02JHvDiNWp6Q+yApYoV+xIfk26gD29rsNF4B75pXbSVlIRb2pzF5RBpCNF
6q7AssBB7cSf4hIcscothYRA0k/l1MCB28fDFmRfkXmLPYCo1nQ5jLk0v0b/Dm0j
cOwlLXL96LAMJ5u/7sdIXDcZ6eMA7dHuGrSgo3uZxmzBiydKs/unKmN7YLKiT3KK
/71E7NNHZM0ZuSOnztE34moKSzbDQ8x/dfl6E55K3MgXD/xP/3OsfYXn/sdQWU5t
caZPHMI3DFzIgO2ftKJ95P0EWxsxg0RxFa5216xZrXN/bPKAxoGz4TBcUsPoHs+s
rns+hyBSk9RK91Ta88odSFQNMD4HPjvkdm3vWiMhRfxcGvXAG36edHeE4KKKkJ3r
APCDcaAtza4PIKanqbOciGh2R1Mx1FoxlzOxjZ8J0b6PvF5bLv580rvicJXl4tsH
wkPZvvYR97OunSFZfXLR2uO9WORtiNX8GC+AUC+WdDRFPFJnMBUZkMOGaKPPYGR2
5yXw2oOICftOLgf0yssflzNy6u3mnbqzEJEIlsTXOpaIRZ783IbIiCSOd32zoPWA
TzOus6QqvlqZM6ZpcYvnEwO17CR1Q7KERwNgodbADdmKZNbXz0gzj+Ls1XrK5hEy
3HkryhVVKHNn5L7Rv35nSTawjk08KloI+nEjS071mqP3XLAV/JJWMZzjshn3R5pt
c3r2fzobzMuCmIOqZOh+BVpuz8ulHjQ+KGDaRPfWoj6myq8bd/lCpGe5x2d/kXyp
`protect END_PROTECTED
