`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CoxOH72J36L+vwsBou25QKKRw6DlMDxugkeGXeobSpG1vHbk0HGhC86ghNLaEl+v
bXUqHNwICgsaBDvq/QVCwkQeLwAYXkoH5uRiTBopETx8CzRKkNkB3lzS74VlMQ/u
teGdw2BFwczRZaX40EDsURUT7Ei7gtslJaYyAW49jprq1UeByb2RF+x8r7fzrN+S
JTYBRRvW/iU2WqKFvsotPsr7ED8S663H1JroNYT5Y3SXc4HiDUpdRSqCG2XoLeLW
XlT0c22P8lNjiA8grIwX1xXAYGnnrfkFS0UT9ztTdI+f2VyUs2qF8YszCOQUbZNn
XGNcH59Tdtp7QMehIF5QflEJCDX3TIpO/8aTMDdcJB5KvSZ7/urAAsM7UKQzhhiF
+sB0U4obmRZcYFgVbhvowYqqh0vcP29bYshb/99zyvRmYGvWmRJ5/aBNtaMqHLOM
gLSBD6ExJn3gfyIapcwp76Lg5swPX3l4RTGizZl0sn6H7ptKyQ+xYmDHS8seoV5u
eYnNmND23SJPEArgHDb+JhRhd9oAooj5xDxvXRJ0GiZFqlFOCJsfeve1durlveT5
0DAstjLy7g++KIOWzexdVQ05Ojb2aQ0CRU+S7dO/+4RfYe4tjOT0PP3IYygio4dP
uczCE+hEt3g8zOQ433/7sw==
`protect END_PROTECTED
