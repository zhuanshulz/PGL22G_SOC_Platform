`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iK5u87mP+3uBxdfqPyoO6DZEaPvou70ynWz5ky1b/kzcnmAbyFDLuKpu7q8W7igM
9Jn1dhlL08JQEsWtSADaMJPDZkhKmUZUt5XTgDi5SSvU8S75s7t1ljG60MBrwFJA
5leY9R/2hNB0x+EIHtExq5nYd//zVcBEMmN/2/6zfmxAGyOxvbHNbTNPvWMqCfnf
ULzG2NzYR3rEmAws4MoZFuM381xy1seFrk0U8zC2L942pXyMPdC0aH/hixbwGIWR
m6/8bZw4+DjhOoOrUE0Zx+ta7SBYu27EsUsxmbbFqU9m6GnxLC5cMw/LUXaUuvUq
t+jWJ7EKQ+jCwLn63Pd5lUfhic3Ji0XVSe6aZpVGqFbo+VVyMvzDUSB5t8R46kk7
gx0QtfP+2hpk4n90LQ4KKPpO/05ioIRmrJwmJpBLlLOT8dikZz0/TOGawDhGTsvx
XAoSYTOjN2lx5+Sy3jcrFRwaVlj0tFvGsT6e4hngBFaz9RkdEd+q7GSGo1s2xfEM
ZQzcE/Y4uSobVRQyHLV3Ge7o4QL1mII8tC74Q0b4iijMeXzKtsTjhiFhTdEY57uB
kBG1+LKA3EyQRdmxCZChOLwT+KiB16KVks+9vOpGow8BQhzZtmEpaYS4PwZkOYgA
eLerVB9aACHxpnWW2EMDBqeLZ3gtd8u4rrWC4NTv8tYk1NwW4TxFJ6rd8ByXO4xb
Z0RSFpWUMdlOnXAFgmDTb8Tklra499qyGZ4xBrWsls/BNnBCRg/dM1R40L6REfR/
RIgKsdwaXzBguAySTJlrirE6ujm3P+wlQcTwagvbzIK0NSeg6xEc4t7Ym4Nci+p2
8MTKKfI/sj5FPnP2IUMvuk1hjzQ+Hn/Pf3s0OyvfcJHGm9P9OYxwu4MSHHbnmRG9
I0joySxuCYcDTdUdzoQDTJo4mqxS+IUGMLTWsmzFfT8uXKNGI0dPCevB/PPka8+S
6sjNhJsB5l8+EJObA8d7GPA3vlpzCqRXm09IIqiwdREcW8heCnt/ZgI+06qyf+ma
nZEkY+NXS8rvSeZEiHP50XBltvL0SQWmkk4/fISoZTI+NHFIKDLa5wT0edq93kXx
SbVHnuUwbUz+cdhNejDowN0zhhD2rQj8+RVte5cfrT7KONe2MGcq2CItalqZkngv
j5Qy9oDCvvzEYHgFbjl6PG07nbtByjRhPnWysAvP5Ii7fkto/Qh+eE33AdHYlFxe
19zffVLfMxgfZpVlNhav3+Ut8NdKX2X3/7nOm0TPR0EW9MmLI8KT2SKMjEFaki9W
RBXsMeLyBC7NlXn+VBFFjMXUfMxlQyns3cgdeXx0PQ1u7P6qBAtVsqa+bprX/VbL
Y8rbgCttWvWA9ZH2mfDmd2EIEPjpxtoCHx5U9nREXP7pmQDC/DTRjamBILd6Kae9
ZP/N4j6TJKRyapvHNvrxUTqX6a+JYDQFCeVvv4MclcFZ+m13md5nVe8WPfF578Nj
YaPjvyP5gV6YWpoCHoppEsi+FyJuzX6dsCJ0iTMpIYCbEPKpt8DFPz1ipaMPTJIg
OFeaRvDanHGsAAqbAnwakgDuqQey66yPoi1isMzroRH2VARHVPb45b+nFQiEaGrg
QpYTf78S8y9Ob5yPCwnehgQWCTqU9/CU0/d7LacSxUgV2fFR7w2X7naUX2jAFMgR
TjGfSYQFNG1kO9yqmOWffmFryzqENodVMuZxvDLTiw0CMpAal0oOy5+UIQUQ/zRc
hYwGsNe9bB44vF9+sri1c85ljt7SWzGlmZ974WmZ7jsW09GHO9MWBVXlZE8Nr/6C
`protect END_PROTECTED
