`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NnTEwV63D2mPlH5cuUv1TRc06YFk/GeeP8oQWs5VLSXPpeB+kapwsOJ9xkr+bSwg
zFde2OywiflOTeyriwhbziFcK3i6KAUzQJ6HFPcaHMHiuU5F2QP0TmSJMYmPnU7C
ukFGkL9gOhL44WdKuHrlrmi0jLPO79g9b0pk7Kr7ZUr6JZtaip6lb2qEWOgNTO48
EEEQeJcsx43u6awi8BqF4WHrl9sDgeG9CB0SE4q6oR6PzGvrRzkY/INAIqC3B8Vv
vPcSwfwg9bBUjVilx88yxwoOmLYZhc2aLmgxAqWIDgtJGgmghS+2mzcLDtJ89uP0
7XiHt370JSM3hO1wiDy6HRk/ClYlURcyMyROJMNW3uon/tk0Kcut4/ZbaMDXaWSO
lCn8CtwUv9yRmjA/ylfi3YNmp3kIERgOoAzUz3kSFip4TWkw9KXbtUdYVzKgFcCL
zs7ch2x9FcaEscbDtOOLr3RgEIBQBFbDMcs9IstoyhNMkH8E5H2t8gfMrLR8Ew/w
VX+vbensGMtaVJtDtUQ5mP7YzCyI5GbgM1BTYHpd41agz/IxLCBbzvBrc4aLBgz1
LCz1rDhUxin0krrmwZhzTQwBph+Id4uUC52gCozMmectDE3Qly+AG8GyIsK7Vitn
K0WN4otvguo5B0wGgqe86NwIkLWnQnzKs27h6FFIl14=
`protect END_PROTECTED
