`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TbD4d5ffZRPiDsestnKTq73Q/bCWAwNoEFspG4d9HZkiEmWLLZI5XmeXrQvx1u2z
OKXvxKUTS8Xxz6NHr+STdoJdjn/cZPs64snW7VlNfiCoENzyj2faoVndNDqVLiqt
Ythtd9yq1XPcGcEFgwVivppYFXWoozCIM2LYarhVoPOQA8uZ449hyghJTwW4qEjK
pIkABvqQKDZQGbRf4EYcZpXBIX6Uuf8goRUwIBCXmoCImHZ+B8yQrTpnWGrvGYAt
HWMpQuPu2+89STCfNkTCawHmZ8WCOg7CS8MvuEPnNjqt8r7CRLMl7IbnvTJzqj6h
UHUCF8Cmb/gaItlNIGq4zweW8ptS7osSLKPwySwtfpDpdTZgzho/3XvO2gZDe0IP
8p91BwCc8EYY/xv2OAr6VZuxsseGK9g6HHlvC/q4KL3MI6EozBjGB2HIQlrzgTWB
ZQtsUgF4HLz+vOdGdDSiGP5IMrdUTc1bGEHXFClxJQ8K8o1+LeVMuNjxZkZVvj0k
ZgjAW54NHZ5NaTNg2JNMIygKR7n2jm864yca55N9mQBJDtsG3n3s+N1njOVc5aM9
LSMFaEW1HIaBUj2qaxmIRlbZU4c1j9qb+t9vFAEri3vXgC/ElV9Sd5t6apvP+Cir
vRhblvVoPfJSSj8vpf0dSsPAxErmZTXGJFZNBfgYffPWteYWCbwrMPNVhDY99nrH
wYijI5XeceHN9mGluL05QkoXoM9YbOK0ExcBIert/eOALdXEZnr8mwC/nPCYDhr0
+DNfaobS1Tu37+/vo7+dOOwHL4jPP+ZvbGYmFrjb4dmn+Y9fw5Sn1ibzm/Q4mOFd
4QwBueTI9TFqc/W3ZxTD5Mem7ojQS9o9Kj9VVlbplXtmVnMBWupdOKA3e79oH+Ij
`protect END_PROTECTED
