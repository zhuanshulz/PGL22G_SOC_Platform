`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U72i9aexYWoT+dWipB5VupSEAe3hWrCndtM4brs1/5gceK5ZyL4logWm19J4d/7k
MfhflZ1d1Wms8KmtaFAuwq8UKGn/qqdbwwtWY38cKHC77rxQO9aoJGc6a/+wdDt3
TePhAxYWXM5bnX/VAIRYoWJHtqd2pdQCD8S5733hb6dLFXmVdK3cUhCAiiloykWX
Wpo3IlGQklBbVjhtxrkc9oidQ8RqLfKkcn1j0guO70hgwctVMaMvahvvUzsCf79T
SfXUoigvxvev8g+G+3yFq0nx4/0yi2d+an1Pp3OY1J5OjtwXJGGKnjzLi+DlDdhG
HSYio34okPva6Hrzbc3VrW4zN0oz5KXYvfzegF9lcGc7VO9DicjM1YLwI6uz+qcx
VytwZRKx2RPffKVd+iWpvGAohU90S38mOuvjFzgq2KX5eVZPySLvAdKqf7w9+2Bk
XijbPaO0LyKw8Pf5h/1SRiSiFdWkrl5VtcXeW5wP3VNXNA8hO7tlIG/Wzt9+3cD+
T3rfX/5HhakCW4C+46sNFvDEIL8CAyVFxlxB45i7NUaVV73h/1pHyeMuRMiasF7E
5jJva6HLm0BjcVsWdjROboFd0VT7YEnxAAir7ZJGNQcwme9qb8uYT8o7XtCp/5cN
tbUN+Lc+PIR5XFlo2aX7r+tKdZhDZ2+/CHKj3+62ghG9DB5JaAheNt0s7WUdTmcs
P7kTbLa+8ryRn6MqfV41dbacs8WNNjVQY+WO+gjfWN1HrSZgddTzKrYaksLSBTF4
ydJtnXh3fLODOSMcF51zi0/CSfTfrEFRcLkEUEx8ND+r3hEaJ+Etn33SwHDFrwqn
6iNvgxjIL7ZBsBzkS2Y1mCrNgDq5RyCfYSZlGvbsDbLzj1ZUs5cHkTgYxyzq3pSM
EkrBwrxuu/T9tHrGq0wmdLFJv9SrGDK2ys+y3YO8hRhYOVFETxcOq+H3COpqOA5U
mWn94TxKJ2oefkAwp8mv8idFTVipJi1O0c2SaBgLK9EVRaCeJuosPucLdShJs+yF
QU5aC9pjPdHWhB/z53fcwplbctPgVwNPWdV0bsb4FmbLlmZR6Ti/kbCSQduO9hEn
bqbeD6GC5U2eyRgiWDFX+a7T7YRtrCvNmcmaS50MbrL2ijM94MyP3XTz45QNCnY2
oJovyCM4wikX7EcJwitrcG+wTvxKlC+qcCYeX0hvJAN9WZM8Pz5g13L/0BtaxfpU
ausTM+Y1D/g+CrPpt7CflLSiNNqqVqyYREWfPphAWSJjWABvChgWxBV29GnvvLy1
Os7yXxbnDfMDORePfMHm7hjlBY+Et2m5IUmUi/Ky2yPlUmsAZotiXwhntQPrFGFQ
OwPPSuIzxfElD8BKZH5MqEgVvvMkdOP9OcaW5BxSI8gLYIn/MTbQhw/aUiCIOsUn
`protect END_PROTECTED
