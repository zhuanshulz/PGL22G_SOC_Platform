`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Sk6WthkhzwpEQ/4GE4YEWcPm3vfBKhpI8aoFjT0i3hkalYDFE9b51v3ztxpO/sTM
2LNqrYhX3VafLtHsNA2alPKo+IfV93UlJKjOcK0qYKESBtdSNnFp8xPowcJL9vaC
C7W0xWcWOZGMZplVC3b6Pi7JjTouoAIae7VsLgE/UAoE1BaWe55tb/oDHV0rKIKI
+7E54UGdWiIS/9AHVgJo5iGhzslGXHpXIfXGUqMS8+9qYgM2kpPMIM7x184PDgxv
eCe0qyxSx96xMcvwGRVvML93hkMpkjNCade4wc5AyALC2yK2D7TveYMXGJs3aEvV
PdorTX4OwUeUmeQQ1AcQsEgv35prqZh/iGx8F4Qz/cQ5xR2Y/ftWvse5O+e5KGy6
rSmz0W4dxIKiMg281zazERPH3DNBDoCRYpDFXerCuxw=
`protect END_PROTECTED
