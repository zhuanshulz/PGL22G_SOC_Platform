`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5b3yhQu+tmHdLbiirAQ2wyDLHK5+CcGrmNR2CW/eAzIjog7FUtC60Bac9l6julxS
3bKAeV51lejjBQ7uWxP5+2ETbwMDjOtqqGKUnaRM618RODdj9gSWwj6q4X/hBdMJ
ztE2ZfYyX7hSVI6eP8Q42j7h6IaIpk95h2m+eNqgeFjo42hmYuyRoBsARIER8tvD
9ss4wUCIkv6RMsPA6HYOMEIM5RJ47emgykH9tEd2dmnLw0ymU/W+IaHhEPPh6AYJ
7dkJpPnB4n0QN9gT+lIP0jzcLKxPiRICy0s8Pz/Uc9hesecswaKFOaitr3L+fEkJ
QaEafohbypo446YqyWpJiLKvLRBhGCsxWRI+jXJP1cqMBRFUm8qC3r4rSYw5KVYK
3ira6VOWQEFuZcFi+TyGCkB+/m6wp2bcMNdtRnsdag1bKTO1jQ1o1ge8aq4dDkz0
nSvscIPoo1Vb/gZS9Hew3+P9msTaEd5MGFUMmQYlywtopQuc+zKoQSWy/eHOltGG
LAArHDIN6LaaeQyzEczEoVpg9AsPQYqrTcAiMvfxZQpse0BsXECZWzsKen22/UeS
9x7ZLARQiZkexelCT4c3PyUzAhHSEbMPlTWSXIUjzEZo00UqF7dSWgNJjB4+vE4J
22uPXT5kLsKxVRx4BT+2sRYE0tSzVAdn8j+jyLx94bwrAACpSgdIQluFtkaFmzCQ
J3tEFvXRcq39/PsmsVK66HkAXCwNI9k9vG2qzFNf21DsvE2Pz+83UcZh6qTESDrC
01KMQmuQTQpM2IbkrPuenpGAHtoCQfVMLhTjwv5TvGHjsbXoWHk/7LAVREwa7OSM
fe6c/iZRGZWrYr0FvMqubi4siKEvmU66M9zcuJnXsk3YzO6/oWBCRano8RvoggK7
Vmn2QBomU6Hd1evHybmVKHqX5xy4N/wM/lg/b6iWrZY9u82OB2nCOqb+Os8RBKB9
iMM9X/ZQFL8e7TyuFnV4CoOcaS+p3ryOJcVWNDvvFln5SNs5zMrAIqhf+MHgj16B
wRqKcWV0TB/6MV9bH/QkRufS7TOB80dDamTYhV75kzKBYeyx92vDvR//kstDm9ha
HdYI8MuRl14ql1C8MTblp0kcvyoxqdeQ4/FbvEkRdMH7bXH6zu4vgRiVxFD4SwpK
JfSa3WQTsDnxl8IU11BZchHfC4AN2sK9Q5NYCDKzrltik0/NCLHaHHjigy/dYCxX
S/WqEpYR7180rYQTA6dvM5G7CiMi6aTc85LQLaGkN0ukktZ7TZu+9c4QMAaZoxlR
lR2U3pUPvsCrpiSx9q51Mp0cyWutchmZO3FVK82FoZXpK31x7oOE76VdlSs/LYpy
f++h/A/RxKNY1pG0h8kCYyynHz2cjqvEZ0WygowTjIBuI/9TQPw7+D+y9N0HCGeW
mzgHeCKMaOIFdOQOVgAjs6Hj+LyYQdHM1uiDF8PEevuxWD9gsqtPD1sNDYamAHSd
AMuwBh7i3PioS06rw6dlsoYkJKjYFSKz3N3hpC7aTKvBFPxULorfStUm2EpZlGVn
MHRiPAGlm5AsBp+q7F/EZI/zB0bL6kFldhRSl/Sb4FH9OUl8f3Nk0bedVZPHfkRp
vixQ7zcUNwHsBUeUrJ4ojb//opfdZFaK2EG+KTI5oga4mwU7U36A3X+o9vgimSFg
11JEtrBygBau9GzvKDGaH/aeNkKURcnaQNKa7KnNAmk+PcamH8ir/KRDnXnVGsIl
lRxnPL7Njlfajhr6u9EXXlkvwp3JpM5EXEqk8NpvQePPlNJXWSVBvDD4ryrwxPrz
4GN3hU4BnP1dkCoGm80AY3ms1jSz0LEXcj3qlmDGdg/JjrTYHtm7wEggp9InyXut
CaOqUgdl9JuNvk5gPoWBw8lqsIqBGapPsoBQ2PYmNFcodZuMuHGMS0Iryh2aVlLe
xXNj3/ECaTkvwgVrJe91peLXDqnQl6t3aEvLYZMtU7gx/sXpAu3cjlFhXcUplaKf
bAv/IQOiMmc2maWic0U/5/KaQg0jFsX7Iekym1qGjS0eU8c5+bNYeak9cuxRe6n/
gHOUTDROe6T7d+dq05grvcjGPcTgGej5k692Zv/SQdDrDch5k+H2+rXYAhvwnMvL
NjOZesAUHPzAeOA/epj0IrwQbSJjl33RCmiTE0iW6GMDi0jzXsL4kgxtnekSkYdt
r2LNUZP5uQJqROK3o7rVXiHCPhVnUMR3e+Z9odoaHfssxEvdlxIi/yVs2f43o9w2
98wOiQyG2QcA3ERStZUNZ6hPtb2TE4lODVS3H4uNisvS21nEneycWHF4C/2S1cxt
zCNmC/AVvatYVOQifHnhnJYN9BenDmC2qZExJRfR9XhH6QtpAcaO29JjstfOcCVE
LhccIggpheHLyGhfrxzwtjsaT3jIZIrPvImVDX4p8s0wet8RwGEjM75z8tqECFAP
6QSOByvz2vu42YAzS4Nm1UKwUCpfPz4+JbUsBfl3o9emb/ZwJ1Z5jYrr92UJOVEe
e9Ydy8dtjcOPGIPZdQEQRg/skOadU0bg0LVD6VNEaiVgh3K8JyZ8qcfCDdmdCiLY
WUj29DML0n4H8fRgG0XZbyhaxQb002TcTB9yDbL7eaWT9uMNBOqrv7NQ/Wcmbe34
0IIFwjEdNZLX9s6MTPOX3JmOe4iaw293vevYXAV08+mOsFkR7PCXvaZCKws5TXIf
rfwe3EqtigyoIz+/GUiLLvohe/HOvikeqw9C37NlXdAJnssEVy2v0nsJBRAYmYfV
YWOEzWW6XB6w3I50JdbcpLKI9QgSQnX50ll14UFpFGSsmZH1J9HH6312E603o0wD
XSK0z6NzEQoJKbd3YtdyvUN+c7H+2SogszprqXWK/0u3qco3fopTqnJ6mXnM+CnM
Wa/QeCQjfeAsvIl/BVhBM29DVSgz3rsBvnfvk5T6OiYaNtgVdYwHHdUkJoi30UPx
NVFGGLuox9RSd4SaxWzPDMtsITP8TslmuLn9bM0Eud049xb8KM7H+SkRhL5GkZz7
swgsCvRCguivFii3QxC8uWdVDl0Azh3SokP5bzMcRJs+OoNNkP3S3EIi2eeUpmwI
e11xR3O9sLI3aeEMcQPd8KDvXao2DX+7JiVHNFhRriVfhKWrc7q6PWcEXNh+n67F
lPGfYakXbKfDz05vwexhSk2mb+JaOw6oIsxXsHnLMGlrAMWYnUOE7jTn8gsn88Ny
ePjIylozGtVfqUIsHUljOofU8+o5F9HjMzEbYpDg9rCQVICV5AfxzdwVIUhsaWec
epiEnQdWUxEjicsSIk4Kak0/iOroWhU7bCd2SEIbLoyjBAECUE//gt8aEkAs2kJn
Mh6//NJRJ1jx4qlVBMzhyKu8hp9PGCcoygEUa2TEjZEHWK8geUwe+Gl0RCA7M6jx
CbkHQYJQ0OKGP7NpfJVDxQe9uF9ZXf/QDnN05ifeVw9iy7bbMaQMkICQVQUejPj3
UkWv1VMwYoaDW1dtQ35Lt1PhxZ6HuNR8I1XeM3xs8/9cHTdsjxIKxJdfdvhfNsx/
eJhcZNVXr1TZOMZUKO5ktfSgncbwls4ZBZgcXORm0SLUEL71oHH1ZvH0xe8pIwe4
xWyTZMfUOf7Za0orykcLiJyVDhu6YncpP4oAJeClOfGy9c9ea7SpYtEM9LYC7vgE
+wrKIOLp+CuGxSpoqOrweseZxDu7PJkTh3nFNb8pe+1cMG5NEi5XTDCvuMQlO2gJ
56HknAe3oBXAvmp6iqkW/A6LAx8FHOFQPypNrJbMpUsqaw7S09XgU+N/rWUEiE3Q
wUGAXPBdjBWuSsSCqmJpmwdLBrfY657UWkUfXgZ8SEM7Sh5v8rFYATFEkN05UjiP
Vjj5JqKF4oVv/9RQefWCMFIl698sLe8xHPz08g43nENZ5Y5wcZlcQsMzUfyIPxlg
4N4YRBv4IdEpn/DfTAoDukdpAdOn62A45VEwJOUUwW8KrWSc32RO7s9sHEe2bbwV
0/Caozx1dTlaWUIqvbycAv1awT8e7G2jbDJZ1hUgLh6izT/RWN7F2w4Uqwzacfew
XuzoGbIGVIw+kodRH+W/9x9x2cIuwZRL0U8PyGLwHV3fgxgMnIFmdpiyArbc5D6C
jjyL0aeZQtXilDTMGZCpeR6oyVJn6zbxBHbXqOZIs2+HS37gAYasFGp+jvAtbxMA
45CBAA3twkfQKmmNypCtm08YdNlPQ/L4SmAtc7VCdJ975siieBgwot0vB1HyBtrQ
hLngue6vC7UeGliI+hIYX8mCVIWIMRYgam2PtcM9SEHx7jTLwevfYlujCNAx9Lgw
4kBDRJng7ehiA8jjrg7uJp9IVj9vHnli73N1ltvor1FRsx5SIR13Y/+XjBaWm3sZ
P2p2ylR5qM705mqwjlMfYGhJcl8XhlauiOQ7ribm9WSz80lYIQt2kcDvxw4Vm89l
4NQEJIrHwlRL+eMeecmASuimcttvjB9VoUDw1PQ92B7xPoJXtJkTsbUWp0G3IVor
6/QhUXbZtqfgWwwY4R2ncJOhQtoh0zfONBP6wLmLi/gr+LBUB3noMc+w7MQJV0f3
`protect END_PROTECTED
