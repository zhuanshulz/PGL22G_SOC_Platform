`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
twhXCYmoqIbjdSx6jKIipFrHNjmgjU7KaqFlkC3LW40HV2KzrYMNzKxSZGaiLsPk
FRexCrWVgiI1BT2c8qK25pYa2CRH1uF8zQfCwG4SCcPDNzxiatWVZnIBzagBzp8U
KrjLCSZYf41LhZCqjtcCHm8tzKDHQck4zip9c1pv3dTIo2mZ6svSgRfRjyr2hyfx
a1+agoQy92wF/Pb8aynVAbK0ePoKnMzBuNoI2aScMzEqVEAg6kvkn9mrx9FWv1Lw
4+uwBJDQo735sUQoqYWklUU2fHGwXmpqxiLFiV6rFBqQ2cjqYAd6we4CGQlUioz8
/2ioPQiQzN2S/7zHGpNy3F0A85u2gicv03MA0Dc/YCLeJOCo5FCq0hpH2B5T82Ks
OQsFozPOrdaCC5oIRZ5X0GalTruKgnIMUeN1FI6q2J2eYurfwE8D99j7xHkaMB9i
oPWvSt0WiogeMTzMTzgKUaIsFKrpnarVWbDC5rReCaYvbSUB/VBwdYZpdo7+rm65
vvyFNC5pklV7Tms9KNovMCcu+0aUvH6FDhFGFEgdu+YcHiXMom4UU5OExSVe8tOV
h354+xgFrAvwNNldTI9G+6V+TnBn1kifSkt6vnAASGOlRqhvjsCbS2lp9DJ8M2Fh
tSY88ji+r2+va8HlMBtGjaXpTi1hFJGiSuz2yZBmX3O8M+ux76lHGHtgY9D9rBMD
YfewkqY70dGfeKnmSijGry+q7OJrHJvP8oonEHU75UunaN4Okg6JMk4IqWC2HV/P
TepDrqZ+Uq8Fz9gz4rffdY7ZPOdYDUvTKvAVBg3wMQ7JLlYamHLIVrb+zS9fOhfy
8NECj01rKxTUu6vOqH8ho/L3HHixQgcW0eZJktDdPO0JDNf+J2qz/EFExSUM+XFK
38CWzK0LysmJxi1x+0opRS89m+xTZijCcl0E7rVQyOg8qqxc50EoDg8bpSY+I2Zl
eL6u8iDZ3T+djhtvN3lxL/nMM/Bi59VhLYNghMquang1/5sQKkW2m2tIWHrm6KQ7
4RHXuMOgdtmIdc4ThNdef3eEdmIuxs/fpQSlKjHTjXFXjrAmgqw2GjdeYNBB+BRV
xmiQRCc11r3zSN0A+gfTvL9KMsVasRzvE8oOeBlSWj1om0CBgmupjHgpGgs0vQCn
3bvvh/v90J0kFY5aLNrE08rq9zsF6qIeK0nVzSV+Gg3lodi4bMkJQMKrrlbnlF+3
Kctm9tJHw33JU46JrXPcCf8m2OO9BkfUaOoPeZJ0hUGBlLgdBouAzh+msZGElCig
nk09ACrPnzZi4gXiKaZe5yVjJoWG5GTXUsidqpyH1GCIRty/BmILXqjzgpRjwiHa
nC+QUH7pp+L2EaheqA021bbK9LFnQ87rnwkfrJ0wIvsX2U/qS25bbqE/R1hFTEHE
dPMYFUlTCL3jOTvP+n+isQvhLrgJ85ul+/i69kmmQ2TdWlJnXBBl2xHFBjNOZ4vP
Zxolttjp6WNf5H7OFkPZmmzh3uWL1+GjlBdoOaP+CRLt1Wdjrcn9kIby95IXArAp
5EbmuRkTh3nWxsuh3r1Aaya8KSKxV/z2OSN9zNidfK069l4c+CO/NuVgeLF3AswR
R/yWNNShuIWd3TH/YWj2Phhye9URiyTyScIwF+2GZHSh8KBXLk1bOL1AofjMkyRz
SxjravT8GcocB70ZZBKn/ZKUEWpB/BczY05NOa7Tks7FnBon8e/OQpdb68wSIpiH
38WvdCmTJTGtjeaCgTitPGNSAh0YAWLbE0PJUKxEdEHObhlX/F2uF5d+h9rF4PMl
v5US6+kCHGYRcZ+iE1G+ANIkZmbH7MKkzJVD4XoLG6Q+bFR4ut+T5TD1RS4daLlF
WzlUcdmLzPUia7PdIlad1/XdLzdaSMkdVsMuLJtxkz/kQm/PzZuflSYY9jFzBL97
`protect END_PROTECTED
