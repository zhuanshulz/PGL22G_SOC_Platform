`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
odGyw3g3iLPoQjCLLFHeipFg1f2HQxoiFztkqqVxfxm+xUTv8CgOA5UfVwLgxmQC
x0vUfykesBWT1T8arjKdvPdt5e/ZtfFYOiBNLDe5LqgX5JOeTTMgj7OHQL/jctMN
4nN2e4zxyEQ7B1bIYoQoFm49uqrIHwLtEciZNoK/DdGNKxCBB+Lqqms/CdoMMMSj
IPz1QU/aL6LCgDo2MLz25cCNPBrUcTEWYvZgzwDsmCTTiE5jGcedp7nyzGgAg+1A
tkVzwXiL3R77iizYqtJH5ERupPeLOIDuMoNWJAjt1jeGQ01MTbrZn+RKvrs7A3qX
w6aitKh1if8G2Leo+MMNcuYxCuk4CnnSNzPJJryljy8w2jz+jJh1lm/ylaSfeFAB
+pQvekE3x4Xffu8ID2GSzcmZDPPuszTk9VttLT5PymPTdzeGDE0C/aloy5DpHwHW
qLFLvqDKVa0lgcQRzCalyr4Ipuz4ULqzPYMlMmFQCi6vRui3hGLw8KJsXxv1xWgF
4bJY7xhZismVyCJbrpeUCjsLXPOOVqIu67+tuCZ+mMdG6C1naMdZCng1nHI/nw50
1TCfrHZpEojXyf3hvqjMau/OBCJurOHDTBny2QyVzcJN+30QA274FoeIJL3hgSg4
nmHbCxRRKJew4o8KQI6inJCXa4gMjs1DOw7F1LgeyXJHAticE1LVzZAuoCLJU5as
KqzJ10eEiz1vGAsr2ixT75k05fExOrOKWaSSisKB2kdOaELuWDMVmb+vqt9t61+c
R02F/hN3AxH8gZbSgdjXJLqAAuWlcNEZjikvR564U4w=
`protect END_PROTECTED
