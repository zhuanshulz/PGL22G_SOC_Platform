`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UuUIm4GL0c5OvcP6nKJVqlC/zoD21lhOcJJrQOkOyAV3QB7Xch7EPMtzIa+gJ74m
P+NL16NZZdM8J4rSUoOI1H5si92zF8oZEk7GnYA6jC0STn+oNsrGakJkW8kMc0sn
fs6x5GaAYBXUm/tVZxlnDo+46Kn5WVSw/tetDehDA7GcTUaeH0yLnsw58n5sHyW1
/S29hn0qK2twPZDqxW0YwrHqVr35llGCypgLKUnh5QM0Wc7L8XTHQDLWQGcRnOnM
2YI66ZwkCS8BL/lV1rNaIy55NJzOaiJ+qG7eTfm3ZV6v6rA68LbKWb5RYPVVv16l
EBFUuN9eWtuH3jRbF9GnG+8931XRATXUBTiR/bcScSEtOjslyyWr0MYBGtEJ6kid
OGeBrm1sEvVOkBWW96WcCVzfzq9mXxbP3yUAT6fwhC5QJaElIUayltH7iLZ+Mvvy
cPjOml9zGEKEkLE9XZj0Fm9x8Syma9FQO7nbru7JXnG/JwmNN3Ms+GezMH5KIQgn
B4Vy02stJZ6rwteqBTUU7FOPqFhib/o7ZtEt0ZB4yyoiFW8ytilK/iErFUUQk4eC
r6Ni6fqm9S/zWMuCgVGZumL1WzGLeaO5PKCaK8zFjIFZbOUhR+kKJe5SFZc/SeXv
JFkBN0LMNu+TyaI4fXBvrc4ih7Wiox8jt4EFwT6+kUi09pi4wzGT1TEBS7PB4itH
Mbtguy+s3wkY36lvLgrsvyg1TdIO9rpkzeuSo5eg8ps9UsK9fl+tDFKmkZ6WGAKc
JJYjlWoXMHcxfUrI+yB0bX1WHCOPU/KPcafy34yMNG81NgtVjFklmZvm2LUYbs7S
`protect END_PROTECTED
