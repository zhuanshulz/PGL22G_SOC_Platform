`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tSW+54PJxrtCejOkcz8192IZOp6kDCxXIyE8xEpNejyIbCEn7Xx+gXP3wvqDl0SJ
7GmeBwcJughkXZdkqlNmXOpTuH5+uCF8lj1e9NClANLIg5LfkLR7FFedneZXJM+2
qCzFY41jYBOJ5BzIY7Guf3Q8uwgcz7x7lFNngWaPHgfnyq5Y9AFYEH+FCk82E3l2
h7pfG+HMlaLe77cSyKRx8hPlf1yYSOpCj9L/4Dw2F0nFwLX59/HqGhRrV92QKUKu
az3cOUVl65wPT9Gzg13d6OLLeOGSbUnnGNtKyuvf5cqABljp+mWgCVxolPD6ClWN
8/2kg6mHf7DS22Xiyx4i/ZqhPxq31E4MagOJEDtZ9M7PtJFPTfNY3C8x27J1j+lL
XPXS/YUAzHTwMAm7d4raB7PW6LWvB4ZBePnwJQubnplZXV/2GSnfv1tPBOAyNrnq
aNL7N/AbphDBKSCIzJE/ZxSe9C9YxxK/morrh+l64aZueMuDguZftBZtVIUM/NEd
EZ5oX89w2TMag6Yo7Vax4HHXuNv5vEGFSCWGA8TO6o+YV+RXoZG0SQdnko0zqVv1
Rab3h3zbomyN0IGiyJy5IPhT6dr+pyUG9wOhUzIdxppMEZkutIPtiwB6x0cWdEr3
QBC1qsDixsPP07apeGT+Tumlv0973CS4rAPVcX5Y40ateljWoCd2bh6xhAof/rGm
tO7zEx9UjhT1fkq2qPurKU4/ydcLYS10cWGGo1sxAD2ils4vuPfR5Lr9H7bW9Hum
4AzUBF38hJwWM+jo96m9RAaM9HApI//H9B5WZo2Z7eDuew2AeWEWoXXn2v8VhkJG
kxgijc7U0Q1+uAWNu5TCrrldPWC+xUG5rkhHcl9bcTeUYB/yVYU2zMcDhACH82+C
OQ/orxH/H3d7S0Lurbe0U2EfWNHpvbfFbRvNJkSJFOmwLTB8J5hhnXppAAEu1TOM
/LTGdspu6TRjKxBfu/p0yonsy03EAxFunARRmyvdxyFFAVB5NuBPkUarGa+VzhWD
1YiaS4KTlHrZ12viY21xTspgykwRtWH5wL+oGC4HndUJXUFvwEM/eVrWOm+cehc7
VJgMIg1202YdqR9joqv1ijjMXpNUMxh931lzxTr6jgD+hK81CjTEq+ORUpVEveFA
zFhU6A/x9LFA6NPZ0A1tGKrKmh8pk3TxqLtm/AsehuvjuR1HwLvjfE3pF3mQMWS+
S1b3ktPA+kbj2TgWDNGuUKWgce4VTIe8yO+jhfAFmPdlo4VveNvqcuEjgTi+GLlN
02BnJZePbgR7vBbAy27D2FHJvTMuIVAn/7UT0Xa5ES69gjMWUc8XM1QkfXcOEctf
1WGQaamYdXs4kf1TvNuDHvNkUQK5TCwuRLsIu/crdrZnDjRZ4xqUjvYP+TxfHjir
nK6rDhgWURJ7MltqTXZBxJJA7aBl0Z4A+Im434MKAgejTry1aBuxZ2wqH7aWoLRs
EokY+JSXj8cOUw0nNgc3sTCt+8AtZe9YiUpOy6vZZFOu7KcJufv5mReZb8DWy2wO
tw5LtgjEWyLPG8SNMPnQGDzbDAB6JLKEzopLzVTuOEPU+HQ166d4iqnN/bhgBqHO
cAYNhHRSCqZiO4oNGVayzx49Qa1ChdcjflzBcVIgjS1aLPlLufuABnuorX90ggcY
aTGhyNt/na+551LDKoHlnjCebTUIMX/kdAf/pegE8X6OcTXN2rl+uDIqkbJL+rRo
qNi4d2c9ebUHxpF03Okuag==
`protect END_PROTECTED
