`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VWiySxGnHr2mRrpRlxoA48vS5vWlNsERr/h/W/uyN66VNvSBsjOrOwLbdJpXgIpl
osNjz8lCE+8gEzqlMlTJbOe5V101Yk70QGZjS+da7N5naGf26gCDcKWkFwEjGAoV
EyM+zb/nVOxcRxHpO7hx42hff2s4ahm5OeUHrqrr4goej/hOBAI1a73cdksnzTms
uENLBlrf+ewMc6B4GWpSywKh58rHj/ntZpbJz5XkjBUQAx3UrC0SoVyFy4rLRJ7X
jKalfwBcc0GH6qgq0KRdPatr804dhEL+fH3uB8aMU9XHyRMTVKSAuB72b7Ih3jXj
erJCpAvk+UNldgd1cYup5+TOTu6Jsxum2j6qPkHL8ThZgJNiwyO+2mJxQc5ecZaQ
3sB9vzSPUBHuPOFPl3b7U3qJP5Sge1Zg+Zg8b8s16RfwH2NsVCc/Z3wtvBomI6AP
sHJGw84/Iy5BmRlTBdin1CgsHlb5eFgLs8iZuFsamMIfsZgPyGXeD7Uj24rQij8j
Oi6HZLMSxRMsgC91EOhnZw==
`protect END_PROTECTED
