`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zUAhoREpi8ZqC0lm6udvm4ahQDaVvObGGeor9JGe8G+MDkaJ505+99fxnbnu+Ulc
wF/mQ27TSC7mcDFhF+LmGgUM+YdAbnMntIA01ObRtFDw/7I97PVRh+XGnHDJ2eVo
UjRuZskZ7SQo1kwkBKpEVihXzUxali6ocI1609+seLiajLlsLreh/mfmnuqajjqe
EhlB7SBSFkS1funHBSLlVZJCNxyAeHJQBdVfI9K9HqosCElt3wDjp8bli9W7ty8c
dyPHX6wKO2ZIFvSH3WV+ACJybFiR+uwbfaVMcEKT/gLFlSyX3dLT3Rai6END+INR
Pj/yAbzCWtGA14Uko+3NecymElgvDPcohcblhH08wRw/lPaJoFoVC2rETyca8Yia
c1E8ALaBcilkLTq4gGteoqaatKYuuS650hJEkCc6/Am8I6AtTTgCd6q4/C0x8d9B
SNQWURik9MbY0WW2yPg9v8eY9j2Ml9KQ7u8d/qfzyHVCihfI7eanXgUnIocq6hVb
wuJWerJ1Dl/n44zuVTaer1Uo3Grw7f4YxQEIs3DiD6CKnphgFTcHeuIFL55cRJnR
fwJIokN/U6zp/WJ0tqQ1DyAO1L5yc6OTRsIHHFMJr4Mul62HDN7G6THRVjbTfSlo
UKVUgspTZ10xBdWVKXPDdtcsMnNDln5NMs0QVh72Z5lA0cSDp5tSVtVfD+7sUbXC
LStVxth1JF/AnsijwhKfx6DRUG9pnjnc7GUQ/4hH38Cj+7vmkyRA3tyIrd+WugDU
JOTvW4sapUBt+33H395qpWBFOFN4ns10ZD/qDG078ukhz/zxq6d6gG94MB4LnlbY
i9qNiLS6Y5PeM4RBEUK++yVICSvhkRnzGv03vR1+6JCtbW2daBwLjtteYczJzq0r
YYidFB2gBQdsLV3uldTy57SmyU8TyhpevEvMcflZd+YUVWIHfO23EyxZTdNTod3x
7Bkia/On6I/C0BUU+xAWvZFqHbDBpHR3CNb0i/+A3YmuZXUILytEPK3CpxS7eSt+
vfTjl1HiVRYxK/RK7HUA8oskLb+GhBEORBEOwHuVVSz79EGAVP7pi52Tm1zDRgF1
BRtRGK8D5X5ap5iHp1BV7XeS+QybWqDFSDag4qNeyRLkXiXeHLt/RUBAlXeSQLGG
WPf2UZfMdiXE3MiQE8SOkixSgHPAer6kQ66z+MH3ua74dmsxSaTlh/oy8HEKktHz
CA+c2rRcG7Ly9m+4A2+9nKMG6UssHWEzDxXflErc12RDaBQY41sE0m+jo0G4u1z+
wOuOJeTD/4IAXnQ+GSFOfjz7dTpt23PLin30KDR3/G0ZxL95xqRA7tQE9Y1ZHiwN
CepAkHr8NkZnteWVMGDoKU1vh8cV2+WyM5HM8brKdzurA4dWwJAbivNugcyueA2m
55tSl+gQwEqAhKjlqAfOAXBvOnw3rHNknHM6fmpiDydkmyJw+crl5kJNXmMou9Il
RA83odL2wOumGGcd7z//JpzlPr/aDcEB61v4ANDilnb7eIb/t2XYnptw/bY/BQPD
hWQ76X1wJmAMVCEtyGNpddO2oir/Yrin8GwcRO/443TOC9Lp7j999lC7Q+2te3Qo
qqsG5x0HMojtZFoK3NZ0Ip9DnTfnmARIrpJdydA+eDJDpYgn40YE5byoq8c4xPrG
`protect END_PROTECTED
