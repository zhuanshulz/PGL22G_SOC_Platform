`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z99XUh/PaqAU8Six70A5sTyWWSWZ5rNQuSXmmPr1Zoh08NEl1y7dTtcWlXA1LU1S
4fDa0pDjH5pXiAk2+VSlQ21Av0jUD0TW2dBu+CWYZ9+4MI4j6yMxAMY6J9Ks+0eO
IX0Epu3lHtOUPNDPL9VNuEh/JiSKrx0oIlee7P2r44sN/wsiXZOvR8pvc5zfuDU9
3zUYt6Flhx9dAKxOO4z4PCkqr0khRZJZ0NESnDMd0iWJQIIHlyoNMw0WgeKaoMTy
BIUalPuKoPb8WjSlhbZv6enCYRRxdGYToyfgtKik68p/gbg9kCrWsHZO+3QeqBWO
vgv7hwWYnVSznNLwfUVGLl5A81pSLtIw9t2sqWl/qfVQR7SysyXu23kge+IdiPYk
RoipjXnCbgdIZKGy7FfmREEcbhovDizpAg4yrV/L/q8a5L+P+DkebyhWgIZTmWgX
XqfiYLXzKgMXShVkLVSh+X+EIAtxXevfE5JDzpGM4rwj6jLlJgQpAV+kD6UO48Zu
revcvA8Gc0Vir05cGXNIpsqgaaGFzTmP4Z/wJGSpGHUyCkJHFV6lkeFmU1Xf2YPm
h/I/ShSlBiZONzHudcZNIg==
`protect END_PROTECTED
