`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nv17UKeBKNCje7JurU/PRbisJQVF+4gI4olmkZZ0VnZY0DdZUTVxpp2cJA99kPhI
y84aZ9mxRr+oD4jto8HJlFhRUfG3Ffh8ZXJa+kN5Wn3BmH6p3hFEdmS32dRg/N7x
h+IwzSFSIgoqkhc6bN5Kl9uD9oNDkKyJophlplNL5ks1N4+KUp99I/M5XltxWSjX
0hwAsIN29tV0CCGgGwwxmBxrr5owRiRLRl+DC/8WOxg+WEn6ggxVWvyI+hrlRTPe
qwSaFcX3PMi3JVcWJi4LFuzBSSc9LmjdMsMLDFJd4FmEOIdil4ArhizctugIOrW4
kCgIahLXH/OdMkT7Y8OLzR8cV/nW85SaYgNF50CvvyoYGR9eV7GawFYDF9rLYikC
nyP8e/zzQkLuulkzJzFs3tz4vIaQAtQpeYFbWFjyIP0pdYv+9OdEAxSyqz5b3EIx
OkLTmOb+aUKRgyoNirogpFYhu7AgrJ1bmmnQ2HJHxku9K9whfWMVFeDtEGtxwcaF
p68rTMwycJSCBrPeET3aqPcHOO3IR/tLIMaqSAG9XGhbZht5ZOEOHxoXALUcfFl0
QRgpCuddJdrlmIuwe/JabsqjSZ4kmDA0SOS08Hhly2sn2U1jCyH8CjAZvVKvtje8
SWyFOzu+cS579U2UESDADe8LfP93cg2DMJPU5UZlRMZJtyYlY39t+wYOUdM3KydF
lci/zy0ixheRxkQvNwVbXfNAT0IC/2og4PYK+XiBGsawerpxCF9h33PD3U6FbFV1
3goSZkDoVG2I+vA+hqy2/AKRyPJ80IOcdsFM2v/kAgU553h2X9iz9PbE9z2vaMpz
STddAOWp/pFM01zpHdD/FoXFtCj0lRJXsY8WvLt8CgGJ8ZdEoiC1+Xfdrjf3IRfU
b6e8oJ4bCnfX5r2yoUqUKt0sNV2MWZsqTuJ5t15njtgeyIR/zK5Jw9RtmktcGZSX
k3oPm8Ugok8+TjSOy8Zh+YbXYwFi2swhu4wdkiMfr86FyZ4nmWPYxnMtdSIecz5p
r3IBc7D4AWAGIRYqXV5zewjG7LXr4TrPR/rf4pOUApEZQQZiI2QTmQFl2/fY6gPZ
Qpj43hZkSEnwv4LIOFQwSqxXaBoqItfRbLIqZtXxuBMdeMnJjfIJs7A4xP1MKRKk
wfSi6r9PZpSu9XO86vcPZ97L/x9rgHegbiTk1LnPaNbwE24JVFDt7IOyXTvDE4lV
zpXOqJ2KvZKqTggsFfcgVxMZ4AF+gPFA0sH88TGDGkEx6hEqZ4e0yObjPXXE5F8m
yJ4T+3YAvMhxaADfsbH8jK4bQd5aRgHJUPtWlm7HEkhQS+e/tigyRffd/gXjnQSn
agRkvJtZSYgXV7IQKNaCyRIbqbOGWK5ScB1BEClBzB6GjuRX3yi5AR+xWhOfDqVF
SDF+nOGHxfL9oabzJus0Quxa1sPG65vsg9ATFHHwpvnqYAGEBFU2ZJwa31mwkLHu
3EaL9KpnvwedBYGaeC6NVA==
`protect END_PROTECTED
