`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JWv8vmRtmM4IpHuzgFU9tc7YZ4HtOGy5oSxpl2SqYVS/QLjsWFbxaWbrRVmQlJME
wpQyG/7uGGFjyisFUWDKazvY3DdquY4Jr5wZUCeVNFi6sJoptHqp/E/p8EpiHgPl
AyFtUBAH0qSfXVnDNQmWi61jQlouN8spExBk/j8rci/kQFIng73gB9oaINVSqrqA
gdKNQzqWjJ17+SzW9EYk2G4unuZfyx+/bZ2m8ugnoK7VONP/Mfv7CrAgR2z3w2VU
nclNV8CJLisVuJ0UYKZ1QHAw/wC4BNgDHSz61ZbDFSZixqfMKEMSz810SiHhlPZz
rnIgMgBSWYzhwjB3p7sMtkl62eIz6Bezb9pbBZX7AFpkuTpVb8h58EF6Uu8TJ+0h
/sKMGRw3TPi7JZSaROFDq+G+cX7B//zbcv6/ib6GI2cyKAo/+HLVPngHour4a6sM
ty2ltj/7vIfK1UPONEsGimSYxIjeIIAnOxFv700TzngEOjGTp5wAVNiOApw3jpu/
5vmpAybaCvwmx/CO9il9wTb5+PovmJmbWJQ+PSlvHpvxuin/jgNLlEYD9GIShn6B
Z6rQqID+UtALn4q5orYlUml3C/mKC6KMmJZYm6b6X9XKmlft7tOu3P0yZu72Iuxj
qR/9P6B6tvDkB+pz95WmjFTXqTyI4Fxyl15HWYlyQZXqBK0Wov3IpT08kS69EPVO
K16tvdWt862t97Nk9VUqIDX33jCfoXe5ebB2RnsF5Xg7eNHtirgsq9xSGH3CT316
vxVtNrFzdXL7i4w+SbxckLOvkd8n4rVsST8jYtcBYEBFiEBf7Sc2/4wSk/CRbLxr
2ylWnSKKyY3UC/nUg2gYZFAO5Ab7FC8MOfTD9I3pbQeMcSPoN7zVfdfBTEYrs0us
IARDn829/Qysg1iPNag9x15baI/lisdgRlofY345ImpnS9Ex31OqXPQbGR/Mdn4T
q+g70oUzzpRq9qqlw0kkUpj0iIT3R7ylAAyxvuaHqCJDVyr00CPweH5sM8sNgSrg
TnGOsRCBw6XFwrArzOkRJlHFSvjnIwVIzreuukWNAol6iJpJBt5MVu1WM31Y4vSP
ntJqbcuTt1jdKV1ZotoFYiRGYIcKxPVj0YACPP1VoEbkqUp7v2HLS9Zjy8aP3uox
N9D7C7guV6X9svkdeVeTQOApnbkH5RkOaJOK2Ds82IxZ5uvfgiUcIoM1xykzqZJf
9eBHqzsAQ6r/xMs89lHNsM5h7qpgbaoWsjFRCMcd0aAIplazvjZZhLtacwZBEYLN
o0WcxczQ8hC/rGQHa8kVALvXcGh/SwBvhKeQ5PQGHPgqioDhpl1UMr95LiYp0+ph
RIsQYxE8CVGUeDmScF/jmb+TH0CLUQmXLDiWjQdl/4mVDLaXhwXfr+/AUzxohm3D
IFW6iYokt/JCRsrwdKnlymL+O4zSpzJTewKDuVBubRVmgZNqcyjbITVeiNGMSBfP
TH1K0ZDu/t0cTTaO5uOuD7DLCqoPNVW8YcqOfsI+X6VHwcbdBH22KweXMNyl1H1N
CkmLvToU8ZarjsgDIkfSCrDXTpHTAQ7l0kXw/gNPO45rad6Z/sSZ11IAKW75KdkQ
wU8fA1aWlSHwu6kZNSv/iXa5tLs0PKw1o82o43eQ9RxM+qg6mPveoCc1myCiZs0g
+P+NGUcGvohN7QuYMsy8si9wCliDFWT9DFf6E1UrGlo7m0/Q4vUepakvUZ7RP/60
gjKB1kMROSineVDOoHO08KxR5mWaf/pp58a0Pd3t5h7P+GGezmoYogzKvYWM0D04
Amt8mPJy7KjrfFhGS1sxZSyY2Qn8WKC/7nLWecTRbaYw3oSCUTr7j8M1fF5cjBht
JdRmGB7WQx0UmgVit5syI/bVpaZFT8GELyG/ayZn778qyd+bvRPZXsk3yUjiaDs+
G2R48KXl90M+WepwplHDhg22Ea/IsbQC9ximKhe077H8F9ypSO1PdgKAARbJKPsd
DkRTRGfzKRyMIlLQnzx/m4+SXYiuRM1WPlI8ZWeTJGxqQ2ZtZ43U0EX27F/hpIGp
fgRNo3kSNwIB13AnjpBVNgO6YLnUo4UF9nufg/iTARq+nxyaHN/xezNskC9u+h7O
jtHDT8iGowfEC3iS95e1YH/eTWw2TxdsH4G15i479gb2JUkMcsDpjLmqxhgHJd8/
+nFY9mnrU25stiYXBs6DB6on0pjv8a/SzWsWyDHgFATO6SIw8wv5EFTND9kJ8FaH
Ej2TP+R7eu8rExAji04WpaX9k/U3UKohdyWTUN0ugnxUq8oCZb/czWoBXOPk47cz
X7VJcoHCJMka73c9KzWcC9HBA1Rs3/aO287vWa3hK49MaaIdBxpTmrUxUmCaYDdD
qz8bCDXvvw7e7DCaYui3Y278HoAS6TtOoRj//Mj5a71l12/Pr3XCPaHP6WoFi7bS
8v4oRXHBCQ2+Aibcoh9JPxZYZrnRjVocGc2xtSkJadMY4lM8oIUlKD6KqYRUuSbn
EP/HDz/BP2uRjeN2+18pDA48eDgF5Opa4BQxjIDPmFZMY/hs34+hIgzpaL2tB2tu
gVH9ots5kxRGqH8mkBdS+gA49BbJ/OSVSxzeKy2I238Y9fquzGIyz1qWv0+ZQCcj
TFJs/t4AdLnSJsVfEbwnhLYXVHFfi2c/wauGKI9d06/zgN7axv6fj8p1Wcu19T+r
b+QHRZXdCSC6GbXfJB7BXFR+P0FDgFlwbW0V6TMBCLL3Ou6wh6FvNDLoXi4xUf5D
vvz0om0G15G4mDN9LpyIFTJdeFs1IbPn6e95NFfTGPYoGGfHKhpfeW+NVjf+hC81
wxrwYgb3FwBCEK4hdzZNioIKQQuntzIAToMo6ADa/6SKGBeUURzKrI2mbKLc2a/B
m8c0gbvVn1PCKfp+oaJjQnH5TGY7cJfg8g4wDn6In2jmGYlsXYq7IMw6GgRUlY8Y
aE8kR3GUcB0a7PcdINQkRsYHsPmRkMMQM7g9PPyEpQtFZlIZyVQnymhuuafb2YgM
R8X1e4Tjuih8Ey211q17ZuPxk/WEIxD1nveq69w2CCNBCne7/LrM6xKMQ3LyO29g
jSy/YFHGaOeMLuH3fXDoOBbSB6wteHeE5MtOLr++OHXHwvlY3ZcGIZ1P2I6xEdSH
LU4TBCR9pW+kLblF/R+M2auJ/GUrimMlo2gzBGzJxz6tNJ4tgY3Poc6XGOzryrT7
L+YyVupicSbY/RKnDe21xX7JYEeGPSelkoCKl55/b7QbJuYtf77AtLmaanAnUEeG
eTuEDJXRVBb/4sT20sJQyXrYOv4/VuQvTi5fEJwTlCd0EN2U6/sOCVayu+RzVGcL
o5SHJbUaAG/FVf2bTW4T0utvRY1PwE4rVTYkue1rvEKToGo9yB1aXAoJIr9zl9qM
vjTeH4sLEIao+8az9Hec1aUpcvNgrn1ycY0uR5Ld724pqtQnHFyKOhlICKighNX4
5qJjanR86I1Q+tXtAOCPysLI1tGMerUJ0HNk8BzKoNa5mOx0qp0mQGa8h/mH7Q24
jX830DT8ye8rxmD5+f6fzwf2myH8ro6nulL4mZ6UnDNGu6Vg7qmI0mxTanjy9W4f
4fjnGz2ysG9oyPRgp43zsJa0DAqTboG7J0nPbXPUp05d5B8CLEzqWhwwOpRR/8Nb
L0AYGX+ZAvWFIHpHcw0NBgZmMWx0sPXJZfEXVq4xnnRmGVrhfvryy5V2mk8adTZW
wAy2l66YbmBvWhEtmM38KqnjGHDJOq9DqB7pFWM4AxiakQM0OoQDgmYBKgwLTele
MLiNaS9PYCqXf9/NmVAgtmvSzMHA59Phmu6Yjd7ua/r7aVW/BCtvqFK2sdvSB3Va
qIiPA7s3N5Og+vN9K3Jj608zbmj8Taw33UaDC3Xq+0vyylVNtuxQscDxXt2azYld
7yvbW5aaIXPBWJ0jECZXwutHucwh9wims7V+Ne+BTTOc7PAG6EO46Ci7MvM6z44C
FKz8bbK/dClFOQTPoZ5MSu4mksnYEJZ9ACOjnevnBDA=
`protect END_PROTECTED
