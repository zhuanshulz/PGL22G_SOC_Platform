`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gokqWtOnKBUIcwpkyta/DOsY8zh+hbLz3Ih8Nc0rmqC3/6I080eBOYwP72bYaOjK
1EVuYzwBcZsMjq7RoSW5v14dqDdeNVDU0276Z9l+tAdwwL+C3PBdnTnRxE1tx30x
tM8LQ/UdD19ffTIzWDOhZhpD+UR/DU+znXGLFylls4FLYS3f2IIYi6041XleXaGQ
2gZ54z2GuQ473sqorqdKEJFvWuc5LsRgUMxoLfEb4lZ+ZhwwPQRx2vyuvPP0Y52P
tSchvAGXWP8QgKy7eY6uNf0+FffxvhonFmUGlATs3AhPmv6XcngEDnL5RmtQYboC
8XdzTOKmd/qqNNfF3/Ki2Bt37roWJn7ftC/dJbrkJF1T4L6RPXPtAJd7Ng3MRlqI
+WbTiTlG+teFWErFalG1B/CVJE/6oFQGRwyzGn7mXy7O1/bSF2qy5bKY3cAyghbe
hjc4UBUyTlctvqTkL4aIGQt4wCARovnJGXKP+9CqOTJaOd/hSs2ZNLEZS/cAdfwt
VIn38MMpIjRSEaWAfsewfa0vsvFn2DEUwfw/o7uX9+VMXEfc45SrEN0Vo4vyTPbS
xm89Y43pOQz2m3raVvI2dTurSUlmg11lLkhipod+TSwSjZk6NZ9uHW5+4Vpvimdw
2JH5G4Hs8DwRB5cwZziza57ZLPY07yNnquQn1QgnNG51Eel1cLbMnoXV+6FiHMI1
WoTKyiZ7U5TshXMf2gbI/l/vdgWH9hBXYnvrR1DeOVuTItniHq2vn50O37t9c1Eg
/2izZe8p8stQlLUhKLtGb5aHyfkCuamF9fCi/uLUI6Zr7S0GLtvtgZyK5/5l/VzH
9YJaUtwib/aDwChbLKiW1xiE6HUMASCtxf7nPd6GY1ioTXVT8OkyZ9xfBo0D8ZLQ
imN4PUz465t9buF1w4OqGLCpojksjDLl7IqTOP9+OOOdWvebLExhvnSDQBwgS7JK
dXBIKLRCj930CyfIEKxN/5Jbj1JV2l8JUTiC9ubohsvQxja6hmFeNdR2K8kVgHLU
iieTYgFD6il7hrenoMLD1OZ1VYabi7dnYinJWokkp6MvVBuIYtRDyrwxDFgpnlll
Q4DI8wbpjUE/as8PkueH08uTrkXOQQpyvABLAAwwINSeAd4wQWOiZJhQ2c1imYSy
jl3aN3cWGBkH3PaUnlIVEyHX5dm4oD///vB1oDSocbnWDjFYWFZnLglzaUvUxA0/
3utA/zqVTovD50lLeyGaQaKisat56K7EBRh3zvdK1IspJGd0Mt3rX52mw9jP8yxm
S/qnQ6x43JW6Oil+9mIGoNCqkl/lAP3FcKev27bMJhvTs+Cw+7q33s39vs8FSWq9
YHH1hEswqX25NUEs6dOKq1SpohtdrfVYWz51cmdIOojtiNlHxAtnXm78yA1mGbw9
BtUgZZTdEo12m1tjOJV9AZ3thcF+FJofaAL+wTMB/n2wftuattIgQhmziRrC2fIF
7wj+CYLRrLlC96RiyqM30sCpHqgSox6751bVrfoggV0rA1tqDhtuidJ8mEklPV1d
vpx4hsheEJReuuJdencOw+jcyqxMCxLeR+RUs98dulCQyaEJETbLTtgpV+VoPzi3
bbJMN0bT3iX0+WrXdhFMRf5BSUXuxN2EhYu9c1cFwyRuAXHdFIV85Q+dyRQb08ZH
BUQWuHzLwzXZM3qbmekDdFAmUGdUJccaqFNdyjP1mv5v+BP08Q8Tr/ub8xxzcTcn
7uKRyMxbI1pEm75kyXJBuIptNrPoyhwcfLryPEtLmrLlSpMPQQGFR+0YBdPFmtbe
6bzbi0tI7+mCcYtU3Nm4A7UXUzn3G059o7E8iqsAdawGT36C2eo3mL+b6Y/JZ2Bg
zIGqhzSFvURR3PDc3KSe51EdcKEXTDlefqYr/L8NdCOUm60pVQRet20UFj+0GKKA
2I1Y9Bj3jfkJcV4tqjUhxZQa0c2OU5Z6NXfx6DiSIyF034OLuwcWMtSwkQ64n+MS
4aBZWwFAfg0a40IDJiKCVGkQpulBxaEbbvKVK9bGgM+bjK5IYIMB5u+kfaxf5YPh
eVfAEhgCTJKoF8hC4N57KdNxjQri6afvpog3cPQd2lO8H/qRVz4abrI08ezz/Ik4
dCSdFfwB6X28Sz1GMoS1ehO5Ma1p3Mpung3Rzch0/Tiw77xxfJMVTauelAIZwqTb
H6jeSv3WLTB5AhI/BFO3XJcVcFgBfjHj7v75YjbaETPZxM+3JQZW65OjAk/MfTLC
HYEDRZVS/O6CVFksjWGtFfpP7QJOZUKjz90BSLZwQHFuFMacrUDv6cume58GnCIx
ItPFrfGCn8Z9XvdZN35LKUmPUJ65uY+EfAmZbySL2+j84UHYh7esvZe3fK54LTjJ
z+OT5RTMjEDlOkXrbGDkTL4UztghSgVjsGqe4yEyf9PcHkF4z3ICwj1Wf0P3y/O7
vrHKbiozFifvyjPB/C4nl0jJfAgqZcvA3k1bg/ODIRLiHt/6HanmMp+mUuW36pWg
AE8dvfF8pTCVfULoWuceMTNP+4CWQJbPpdmJ0tDWkBLfLKSnx61FA1UOnunZUylz
8FX2KjS6WcjlqwuNoYRWn1oHbD6XMcookhrvOtpkIU/4ajmZkO2XhDPPlMkti8Ck
GXdmNty6JSdtI95eDnrWzn0M6MLqrwRPGQ/hKxe3M3C+QGiKReX4vCiodG30LOkw
HwJiHEcglWhREc8uiZX4m2+x4S4fNZoTU1K55KJqwWI+FM+suXjwVE4STrlD0z/O
Fvi1NnA8TpK9b0F+8U9ymwoxCddy3W85mDUzfy7JsBSz27Z7dGCjdQE5LCXXu3Gc
Jov8mnNDwI6E2l97Kd8C7bTPuF1a4QdVkOBu5PZYANyHhuCX7JOfzqD2+U1FhiQx
Bp0F3Pmonidl/oT5eOhcsMZqSRrbTyFTsFjv7AjuuO+wr9JUwDU7bGZ5OHn4dyXq
791/SzinI0aL3W2V0doU+DJUAgU1z89abL6GP2zFhMCx37t/u25JSZxctPdu3g7d
vWC6tAbe6T6ffE+zYjiet3d8b94PzOvXvWRKU6zVXTHm7QN3BggN1m42NUM5hdKX
wj5nBGUp55a0qmyfhtVXmB9rgHmAgkCHNJby+E4+P2Sv88xPQvXv8qBcYc9Ium7D
6kl36uzzS1aMo5Zu8Vdr4w98eKuHD7lB1HJiF/LCRbazR6E+SfHMA6R20NK/MX5m
92oDrIMqJLy5h7OjO4P47AYeB5cdu4aI9uCY7Pzbj6Ig7skPS2trEgyDz+dFpcZV
pHjEdkG5oT2OC5q3OxAJg8/x8sMbxglwNKkfbL01bdOgUfmMw9Y0yjHY5AOHdfmm
ZUk8azV4I4OM5/xY3XFaue7F+TiG7+OZkEidtql35HDLFh6iXlwVrp3ykCnNrQF7
G85lNQGG8CLxgga3php2jS3RmWSMR4FDqSYEODZkfYOrf3h6RDjw/u3Nb5yA8ubA
MZXrjp82dFqGf4WcA4j8stCeDtuheMMNJeY4o/bycc8u2LuS51xuIWg+gy1hAw9Y
cdwKRAVpxeKfPj9TyA1r9fX6O7CD9xHzpJGDYtPb/sPySYmwpSEQmS2Fq1OS7cZx
ENmo2//AggBXgVwCtrRx/H+/kfSbI0zxQdr7XopDo4iTCi+9tE8x+UhsSchwO2eT
U+gZJ8yUf0MFQa2uJ/sk3nBbET1zQAXQs6vXScxFkIFsEhvev88UNJLVhOMMqyvJ
3Hvu8mCuGUOLMOEe1RRzs/w3/ij8wW7xN6uzS5kEioLoC3tMOT0LPWuVZ9PWcbL/
WxLrcvgyyCqHQCO8LU9rvWVwh8hehttdrT8F46eqZ9qT7RvlWLT5oOU2MibeObqK
4OQII7YLRwW7NUqaRQb7V0Z7W1G3IHVnOWISzogtJ4Kx3SUo0HTcAnxQsFNFs4jq
H2eMaUp2DEYXFQr4sRtEPXfr5dj6pym8eRKbJySbWgaFzx40Cg0ngA2DIRC5GbmZ
AAvAzympORoL+aQwekcjMaz+hgx7bzHMKFkIrWMNyCtN7LruDX2hgtvvZf0AxrX7
9w0MKs5NTsde+B5LsORWh65VyJBYBbKJ1IphvFYkZFNp42ybXV1/GplkgI/PjR1Y
uMLa/jt6IDqzfq3rBIO6hnZwUnyZz5pEcPAfIQaP1yFjRwZTyNF21oqrd6lJkejv
MZgcG91lKPnSbEfOURSBC+SKG6tLA7rVl4A5ZNhyIxybKzzxaHZdBLQDSW8u7M/O
n2GoYsBRAVidxJ26Gx+FBFU4ZuoHsIctG4PBmiJnhfaMQ8Kp2awe9RbFhbS7LMHk
OSvR1moqq9PKj5YXcXEbnMHsU0iIhMVolciNthlvRnTXHW7TLQylpSCa4HMCfxrL
TibrTNNJCyK3L9zTF2nQKPPutrnX5vou1Gm20XOceVKa9l+2EC9doLcD+hHTN1LB
cGEs4BIJV4/y421Wzkzse/ZoUQDJt3bYjuScJr3ygdqEBw5Fht0LMO0v4TbZrhMt
F/CWUn3vshm+WjwJfErxOq741jiKZ/ycGZASby+i51I=
`protect END_PROTECTED
