`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WRlGJ4KZLwb9LCRCFARs2qpswHLhfYM3vBTZxzWDUh0XTppYUvnWssGhf3yVcJ6R
4BlkpAasGiZzlAHJO+/KIWvpfXElAUUA2QKeNFQ8lx/gF3H/ttNM3pJwBJOC8AU7
Z+2UyUQadRjJAMXFgMVEtLgcOYfvazHrbEHiP8gWnyL/LwWCQfReA5nyqTK5e67u
OhXN6acEzWVoDIGA+Qj1vUhpG6EGY4VLLNEzbJ9M7g9v+IbiLejFLCp4HtOJV50p
akC83LvtcWeOjcVhAVzjP+efAOCwQ/Ke21UldvCCbOhmtcqIj2OEsIGIPmg7gJ++
FAdATnndexrGLQgYV0lLEhyQBxt3WjchiDziJ4huryI7RIkr9KP/UHGpc56DSwvL
13sLEH9RTfSFnwWjz/KNwn7yEPaQPo6ODMDv9lYq3C8XsP1KnudBWl0jDdvr+Zfv
VhUn6nNrLPeQU92+ZWhqtnNfklDt2kgTsKidQ16vYtjIR9ztrczZiQp8LR5HMmQu
ljmzvQFU5+d+Nn9jpZlm9lN1Qq7rlEs2QUu+1CYSy4D6/t7Jk5YMyj5vS5Jty1xO
alUj4koI7hhez1k1CHLlx0z6mYD2RNE92j5ZAB6QcJm1kN55KQXOvP0V/uAgNAJB
4aFXt5na8Ypa3kepa5I85rflLjSqqnnMV+bSJwmxc5oVKMpH34JaLf4efQSn4NvF
XASpq6MZEX06MH6rsU2aMNwL4tGo56L+VjBOVVaqAr4KXCppWuMz6GZSV8qK3oI1
pCupv5JDPRNiMU9UtT4tSgbyS76m4RbDIni3+I+2a3dPamza1boue9i5qp1grAoc
ceAwXCRs84pDJseXUitMr9fEY3TkrjQAzHcBpXnMvVs1ZfhSoRHWUlTsPg0jGnwv
Q+WO0NTSIHAdo4XTtXYnFDKRNP6p73KzAKaa/nSBqzALuM3UyzrroajPuUKkEXWy
`protect END_PROTECTED
