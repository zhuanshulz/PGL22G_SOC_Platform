`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e+GY7GBzjHIHKNOX+3ne/2ePYYysqQyY1xX8JygPMTYr2rqGd1mMZmGLkjp6/j2O
7p0+/6Q1Pu71JPQ+jbuPqGJ5lk4Qlwp2eai6YGk/UBV4bEvGrQLVvbjkFZgw8Jt6
4Dcff7kWXg4T8BS4z32isoQVvLCK6y05ubbHVY9NuLlP4jZsQsitt+rpZv4X/HYE
8yoF+wYUYyXcu43VR67i0FOr2Wa1zLhb4p0P72ksSt3R8NMYt1IiLWK8xkmeTqTj
8Ao9nYQau38uU0PpioXk5tyZEpLrcCkEyN0nB1THSOy3t60NoYPcOM1Aiwzoc0AW
JU5X6E/53ME16VuDjb5hrkXLy170mAAREaSclqqAJIlzk9nfQGbcwX1pQ8aqo+ow
w4fZkxBuiSetRZsQt28NgWmL2TZXzP9NMzmFrXmw76zCJEf8NnQ8qkS+2KE6n02D
eCRfHHg7+qtqg+gYmhYRIXdTd4yHdQgvySxSkzRL/8iTqlw72yDmVoedrDl5xeEH
NtD3R4YVjdxoOcswfv2q/aord+ZneFwJejOzB3uvWCBsBh7bC7PhQnXWTJno3kd9
d5wBymiuIxb/BxyS2y/ehctpOPKEbjn1RKJdDu5/xncgruzqYHhyxMGltmxr0YNz
8NsPm9+rdPLPdY0okdCqqrBiFlHEiGZasSthivAJ5MiRhEKObw47fFUAuFOqhZpO
WCGxgDfRMCjuB39mV/xuvgbbsAHNWqfEkHLPf4k+uc1iabM6q6dCt/YNqOpvkwT2
U0EvNQJuJWvryhHD6HhNDsynDSOXHZXZ7pEuceXz6oocK4TnG+0pmmgAzNx3Lc1Y
firXrjHszN1b5q3CxZ16XfDO7+NhLnv98abNztrQ+a4=
`protect END_PROTECTED
