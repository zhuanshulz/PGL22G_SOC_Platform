`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7nNkTyRpQ9R5UmrcAxkOrO36z/tD1UWoOAOf80NB8CdWG4v9GO4AqkV2vRItkcwV
kcPNy1cUKjzYLudcv7ar5X4Cbyxz4GI0G9nV4xldqHRmZbAcraMw9NIQx8mcxtZB
LKznu7QrR6WPpjrIpv/yp3oRLYz6aRDUz0mmXKvA6iH6Ds8S+GeGnlIrmQsgKvQC
VtiiEboCGr1/K2ScOy9kQM/SUL/kln/3ggjds57/sYF0LG36zO4fTYOH1/h5SGEM
uaMwH94ITzCxhRKl7ki1wnPCq8hXs3QeEPnFa3YQm4YvMOrNhMNezg64nwUMqvJF
yqbWaC8faKSNfi8QDDfmxcem8V1nXl5hYko3fSlusjD5DNRQhOYDd1dmOxur/d92
tgdr4cJ1UGvVnxn0q3ESuk1lpRpsjwa1vD7lHhn3EtdOi2yWNeXtQXzqXQmsGA3F
1O4tKrIO+GP+VoQJELHMoQfqAPyW924XOJF8Ju05Ya/HiEPdBHc0NBrygYYl7sqB
pX1ETmhofhIAc46ZRT15XkQc2X3VBHLvaWCFYFC2yfdPzS5Rd0d+Z1dbnuy2i8ds
xkMObvKevT98IRMFQ3WBBnSGxSvjWGVpt1i2p6wkdaU=
`protect END_PROTECTED
