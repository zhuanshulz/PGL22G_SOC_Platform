`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GHKDu4UR+xateopqwl8eSOw1zWuDFOSorwt4lZTnIpoArSMFbF3pLY9mmpaXP/uA
sUrw4XytF4C0u6r6oXLASEBAARzLbFZTrNMvQl3DO5y/Ppuosw4qQ/RV6rR5r/Fm
NWLA3XjTOyz94bN1KNEyhleVkLpg2Q8G50AA3pdJjIg4khYf1SFBfyIdMeEvEQCU
Cb2QfdTVViVvja0SJ4D2D6T5flt+05ETsvLgBkDG7atdGj1afxBsSnFxfdeLLFMK
788Ek2WFydKrzopBKdaZLLmtWXkfMElXxNYk2pA4dJONjlpU7jWzkXQx9/2ObC1s
dB0k3/CEALyL8wiLS8RUnko3KKf9FbZRQTLe8ONJU5/lSxZLzS7wPK1GEC39GFO4
0beLCqmonAkj28VgTpAfn/B8rTbcm1cBoDAb4EJSVYNWhU68Uz0NHBnL9rb7jvro
hfimPPyJBPAZWRcaLw3IWhqxSdD9mBmRxrB2QrVwd8ps20dNI7qy+zbB869QXoNG
2sl6ffqj5BCySxoeYbnyLuju3KKOQ2hbHa2ctQZ7UOuERqW6HcM4Z7VSdswbVvd/
zxf20iWvnS+KCPjRGfRL8KxkZEH5XchdBWp/tb+GNK6JDQBY0juNKM6gsUAXMJdK
qUYqOLCIg/ymbPdEIjx+HdLy0LIM/kxhAnXvhgX98+hGoCkzt1MEAo1zUoT4boya
/Ots3zK+F52KC2HkF5fKN52ORlZzOEXXI2xd8IePtVpD90qnwOHAKl3rlmyjb9pz
cMZ0xro253EdN9hibTdgR+nul8cICXkSS2zNXYJev2h+sx2LBpQfMal66Ih4o+VS
/vz1MpqWHOPhMc3wVP6JkLV9dfsIr4YfNL+gfT1cCUGzd3/CqJCP99Jd+hN9HiEv
+xNwpWohvmfbw/qk4yXE6hr0AGx7vdjhIrovlEONWKGxmUo0PGgWkW0+f4FvqKAI
yQMwISN8rUkEFGh2MsPKj+fyj1IMa8IyEQFCP97NfpJJxKPCdyD4OzC/nVzyB3sC
e5Ll0LTiQHuJFsAj+NEvSSeX5bxaMzc9owHP7642a78lx15njd5yxGILQmHUpN/h
jwY40fN1imb0Bq9f5VWfd1hwyax5iJmNIXp24+1BhM/maC8kv6X4Ny94PnJgJ8P1
fk74m2nWgFAT5R5+ZofI/iqu8R5bqh5dQWl77lEeEgdTQSvLNNa6DFlPcDDNQrqz
ucFlQTeiZ2syG8nF6sRcKqE6On1CDnJfI157McEvf2XmyB6VEhGu9COwYPa3NeEX
wF0FfwSKCxLQt6MkJJ1PSY8+ILR+JhIAm8eVUYZ4x5CA0CL+4HtV4bbN7eSNjBra
4QS/ANyD1Ujp6lFFtxhLKaLJ4oH+XnNDYJVLjVYKaZrlPU9bdbLboxpQZWPbB9n4
rx7MSXWRDJ5Q7Ob0jFufOUGubILMc4ZbN4CTm0UKDFM98Z6SEtQRGu95sHWGbH4j
hMz3AyaScv5acOmj2Y9z9I5cHVlq0KzW40BtekzUPWchHRxMJm9/zmCp/+Poi6up
ayFv92CzYJSw/8IhCahLUJjKswoIhN0daWeR963hZai7rsSCWKa7F16drV0WPQvs
BueGxMQAuN06p4Qtpl31SPdCawLkQgDLNKqCzw0frX4Zmo2bU2qmsyEhgOYrONRm
Qky6X0ptvuq7iA3B3w/f5/R8krN8du1WNs6m1f1QlnEpefqOu5YVd5GVy2oVkhh6
fmUpFTmlydOxZGszqyR9H/X6QTH2qLF4dH+IDkkniiZXB3DbdMdeKwDWu2dZrk+s
E5+efi16np266nXHwbJ/Ug/wkkrGi4fZB/RBvL2pvvENofPhSv8YW2ICykqb296l
Ia7W2Bct+n+t4a2UFBmXIMGnq+5+duX1zLqYb4JRXTM0Erjb8KCZ7U09wVQHPqg8
shCZha/OGh0EsGqiKp99t5BSfK92cUfwNKmftYLP4VwDCzea2mpMGDore9xI+ErR
zFxVq0XYsie8oom/Uq3WH8t142CEjjTml2AB3qbbyJ0ABqS5lM9djaFpibgdkacA
AAjMsSBnS5yYGkueeQ3bf1WKQex+XXPCFc3nvnMVxZur0OKLjAi4dEbCgkddzX2E
iRF+7ORIH4KQUfyLDHGIqiHa5DOpKI6wLspjbbA1j5R3GLhJu1/1Xz3VFY9vVQDd
J+fMzZX1TgJNvPFjkNfszCRuiBbWLa6v7XHkfh7c0uY5h+VwDTDkaf9PPxG89dXr
JZXqIIlpAMu2sU1lDQLSNRJWDCUAcpa+Mfx2XJYklJ2mm5MBevq03ScL/p5jiOpD
4Fsf6R1VuIVJ79iyF/225XmrclyRY3gYlhfaL7ZGiDEMxAVh/mKZGvngNAiDBWRn
LZ2UAn8ajrPXxNJ7blETdUZAYtcLbyxK7UfcxOfcQvbvDlFU7Lrz2yB6ilDSalFy
YaBuYywekQGKORT8lMF737dZ5nrzUv5zorrEi/U0RtncjUr5hrawWWJHGlLf9BDH
x+SMS2VdcXDRFJJCop9WibutRc44YKXkpwp9hKEW4B5JW27UELiluGXYIjsGeUL1
uo3sSczF5ZKsi3htmo1q2J8gYJqDRnO3uEytJok6zumQitsokv/YnfvMpNd+YlEA
MybIYJ3G8odaYHD9nuSHiRYN/Se3xw6XFaWMZC8eY46L4e3by3exz+wk96Yi8Lym
Vm9Ui+3yu4XfkOUCs1At4EntA7wy1sVY7zRkXhFgSREpRVhWBbsHzU9go31iblW/
082EUvkK5PIdSeXp38e+NRiH142csPmDvzs0lFhuBBQS/SKicvPCbIQOTdAiNXzQ
1XFkfBnEh99AZF6SGuO2cZimI2l0s0ocpkTMtK1yTwbg9I1/HyYeByygH0PMHJ8C
s3o/lLTnpuprIw0pfms5AsfrcjLaZWC1b+wi/Tg+G9Ck0u64cvtx/635azexdlg9
aR0GJ083/VkGtSm9397BQf0VG+3v2oTE2vvlm6zp7+PMN2TXBzDaQA0G4wM13agB
0bRPObW9fixXT48TaDsmumsLvgHGhvauiLpxT2JoXy/SeI6piALpxkFOEmkODMNg
HvJop54VYzRI3YvuUaIy8HRUvVNVtVBX6+tKM13375ga0avneyweVPx+oiCIomhU
8aUX6QgxvwaeUQ0HwZuYWjYVSHBZ7jz0IEfb7PS5lRoRzMo2WtAYLIXehpypKJH0
b4fvDsRFdATDV/uxb52IzcDyuwnzMX9mlZqCGFX0UiCZ3c0nbkYFfL+rlHQq9Okq
662GmZFs3Kqu0UM0eyuLv+T/y022JFn5sDFgD+TVJp3vmEqsNIR6P7SIUkxbPnQN
BVRHqCMxs5xCnRY++DbQFofu3NOJtsgqSw+2Fd3fVOhaf+tIOSaT8KJTFvuqJoBV
AxMkeVM2BhqBl5rHNP01Tnsd3WTfaMp1WvuYZOzpZhDjBdLjFjzuw9+7vZy/j0UY
WpZl1T0xpg3xRnj+/GiDduw71/2N/N+rmgmq+scDPwHyMsIp79ZR6spSEBEGhwc6
xjfUJsWQD363kIvM98bcdFHuBafF7I02xG4A0fWYQv1AkFgYZb+hP9m7cpPZPZuh
xX+KnVaG67CrGjHI82T9qGr359B/W7c7RCk0iOw7Jcrmq5XqFKWwoXJPeveoY4E/
0Qrr/I0ZTM9clMle4FwimB9jvVsjq+phUC+NYKLgLvcvTXhang2gL+rZElMg+w/a
PRt07OrsREsYiJ9Oq3FX5YgF/6DCnhwStdh3ygRDRlxU7sYS8a4dBI/bHfeabtaE
XrQZ9y4EPn7domYTmWOMD2+N/tnyNtB4/ta8QTl7WYcXZN9A/zVt2HZz/9EvUM7e
SiiTxlrSmwxmS91j8pEw7RtPLxZhRPud38pQjBEi3TdoobiTtbjFqAuqRWn6Pd2l
/r62i7EmabdFC7ihR83hnxTxQJ5hv04X7r62kAwx0axJQsyZK1cbik++zi3+ELrR
WDsI7q0pZjMl3Om4Cc/euDcKR5RXJOK9sp/iH4inZzoKPdSCqonBBfYloiE2hrki
aPi5ckPWWmSWyBxQOlHAwOP9BTrsyO75cC84Xqt+FxfKNVIZZ9QGnwON4j+HwBQ4
GTiprxoM0yyViVo9f7HfJvlPcfaBkXzB2Hqq8xnhv/NUqkgaI08Ehu4ZzpSSu4/z
lS4t58kvV2JSZ80w05aEhvfCzuD+L+lpaHNQZohucMOCwMSqTnuJ4wYIPxMNG2Dn
rY5YI4S6OtUiZRFHdbm4Vs9elhb6rANQ6Ah+jo3GZayi9wyA90WWGdXjL41kTC9P
LurorpGPKWlzcGmYyI9l4gkqOG7j+06+ec8fkbGxXTUKKHtjfL3Fb/98u7HfSYXs
LlMljrWP9YFOrgZ+2PbwWZhAcmW3C5UqTLY0QtvhUCZYfPSoBTDCW92RqfeFZz3I
w7X01MmbSY44Jt+hXVIUTjgVGdpTFAkY+PbLAR5+6J5TQppnqpI9ETloS1NOpHNZ
Z6R6FR29Va1hYMl9sAqmeZRyeiEMoM1b/EgSQzwp/yLvB2cwwaUpGuDpXzQ1Xwu+
oTfPGAjmYu/07cjyIYIzmpkPeKLzQj/SjNGVYz9Xcxll0+0e19Xk0zQLYI17aWUi
H1YQFuCPi3S4jN2nqkGuM8UEunrECTAzR22Ygxvtrrms9PR6EbXolnijqSXBAKBF
GlP8VxIYg1cpztxtluFkBVB5YhWPnqPbQsn4vA2+nE+Ud8ZKPFonuPyqGCfD+oi9
83CapNXREjdzj+eGFgEzIZJPcFWdTtpdMSLztm1BRA9q51sorX9jMwxctAnMrYin
2fnTo8F4LgV90cO4qBky3Zy9jPvk4NJrNMlAxtCAfsXLKFw4+8uPXgFE5674vyZJ
b5z6045rGV7AQz3usCqCnD+R14EasTNsFLK3v/RiSRiQI0ne01GPP+F/DD49C8RA
JMOLTYNkA4ITTj19YoAoM2nfi3NLVcOlxQmlqCLFM1b5e7C86LwcGT5uJQr8KtC7
VdhKK3g27T2YERq8cDuKka8iPNkAbfC5+YzBz5SnxBRP3SbX8BV1kHJqdYXDQ9rE
hBfBNvA8ybnTbPV3kqQ94/w5J46a8LgxWyw6AmWXihmGAHEnsqoSJYxGEg8K+P5b
GlRIIvAC3nwXv0+afCYNDgSXlekUY4033PQA15gaj98L9wPaQRExi8RC84v191SK
vNXN29vE2xd6azNkl5otMwqCWJLlhTPHRN/s7JEBIRXLxh5jqtnlZ6sdSCVHyMYI
JAakieTo2+nrT4ybRwmt3p0sbk9DT3z/NDxGf+AjL/lN0zJBpUHsRM0HKi79Cxfb
5/hjGqh6PXjNvW32zjpgyXd+AQAvpVL2LykM3ihF+83+0u8iJcD3iq66ijNhD/u1
808/vcOnpsSd+GvHoAtc6t3rGttI7NT6DmtIGpPh8/bdfT9dvC84GYTTquMnnlPM
jxJ31EdCxlv6Bd0T98TunaDUfRNdK5IKow1fBJwLHWwhGP/ksey3JKZxwCwv/wjU
RWutxz7IISC1bDakZtRNXrfLP+ypGgTYnZzq8BcyATin/tHHFgX745WjhzXVH/Jf
PrT2e1PGur0zgz4BvGZWFokTFOZ1NU3uchJfKKLgAZXqQCnqE3csp1OpPaOkblyI
SMkh7MDJG9kNvOWBGMH5VWqdIvIZUS8UktHziHPwINT/TxYvl1w53mhVzDgbYTCH
7UCZ/qbkjqTJydYg8hm1aLdwb0ot1P8ut2ReyBGfeQs/DKtve/8fMKwl9zpPKDiq
5uZAob/C64J8wLw5w8QrppGIszVsJGe3Kicv53NlDldVXA6SgarxV/V/eAC3ql8f
yptPLxESy8KvOyZbpjURl6wOw4Maje9FFTdj7L1NvVCAuH9v32A5P2zR0B2GVEuO
2mtiCz3bcInWub0tKE/4mb/+Jdi1XKOQW865pUygDVYZV0eJNxHhiwKLh4QmoFAT
csid2vr73pcB5AC++OyNUKEu/BKQT+mG0k/09kOcVrZn1sv3veAAyXOFKJEfl2Ck
Sgu/H48xqHY/ukp1FCjwYhoAKvewLBsvJwVnYJ2O30zczyvzTZx5OonleMX0reuu
4CbnpjCFdz0qLWeNWHL68vtnIGr2m2ZtzXAQ/wJlTQonKuKOnDg1OXw8+cSVqXY7
`protect END_PROTECTED
