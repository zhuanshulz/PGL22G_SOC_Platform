`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jltBvpACzroCZ2/da7Q+J6nVP7SnHU1djD7zZhFF5Tj6+1AU73v3Xn09ovwmSLIz
omFm2Rjkz8gmLcJZSupupDms/wWQM9/746cSU4KRLQEmxXKRPQzrohaGhvGuTVUz
qPknzNtqrzB9X3l+/lLz6Jtc0YVh9jVneHPA7DYdjc/Pd6Byyl+tUu+l+3Dci9aA
PGBxw71Rwy96wuKtvQtVrRgOXkKDyXNSWrQzJDMw7dNq5gv3DzRITAKoun7Zx2mg
IUTM+v2v5RfVxO8fzHz2ddadLSG9SfIwvbZ4JkGggNL4NBAu/YSxn74L4oUQFbD5
AhWHSPYspqIsDX2Wpgnfkq+Vt4miSLRZ1Dbmqto2u/fnIzX7iY9+Eo/z8zz3GhaA
OMBvKhtfZuHbfrP1wRNfi8vpUBsn9MQg7R8dU3dIqCU=
`protect END_PROTECTED
