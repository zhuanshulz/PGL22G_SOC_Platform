`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D7NgPcQs1JyaCGbcH8o+i7UANsQCaHK+RgG0xn+IFLxhTZyAqwGJJD80fHeqRd6R
XeX7qHZUd6x0StrV14Szf5L2A/Hqtrz8HlousQxNioHJBV/fj5iPW5Gvy6Cpuocq
Si4cp4RHXhj81Y01/kgcQEOEVlzHsYJUBkVDyD6/FrSTwtMMbaPc9mmuAD12zLxS
b1wVNcOTRHegbDRcrHGjcoOEcJQ9BBKQlSwcslncL6I5sCavF8k8eOKcglJql1gB
2LmwBn+yodNFerIZtIja0DNEbfGDPtJZqYcmIG8dxam37/K/z8czFt/0A/sYb9fn
VtxqzQjSJqmfcjPrI6c7pcR2ncgLxDXW9Trl3YTnjZi69n3EElmKNc7BxaxZGq8M
IS+NcEgMma42IFIbo8hIFM3l9Lqcxf/vzv9HqLiky+hsSC4aVWLdqFDT9DChmT2O
425hsfbmNts2GiyjjjwKKVvPLlWRzu7aN89n5mKqaL7BCwSo8LCZfftXGlkEoRqt
3igtu23Xa1dQoJwjrOLl5FZRivK1JC35NOSkHV++h+tl8azG7oahLgrVHTIA7zLE
Aka2f5wQRVTXS0BQzluHxzZBq6wupyQsfokcbvR+6spiAt4XkeslQ8sysLcom1Uj
F2GOZoEEyU0TIz6+D3AXnJ0nLjsb38Rbm8NhJumE8PJkgxOJ/BT4CJAwhx47Yzq9
ITQ/DKo/d4eyP6+fOJ8+Ha/XEL4DQvYPf/YXMdtQZPOxIhlvcmsTn5E6wMu0FQhS
sqc1e+a8belknOmZ7cOIJKJSbAgeohulAJdI2Qbx7KuyXUvJn77VRokGOF4lZi34
Qxrh/V9hNVuLkAph0llsvsypCGaaxnkGKGKB1FJH1SQ6N6AlepJwnAkbQQBaq6XK
rjWufR4cxt0UTrAsxoF6bT+6ZpSC94ja6/qazQNwdJ/ewR3ORqaQOHtIudQS2yvl
UzVfMylQLRJw6lqidVRzQN/xI/Mb5dHsJf70uSQm048+tjzASwehitZGZIJuhg33
jp0Gh+bqPyQwbiooM0wA062JThd4k+dU91I80DfN7P7r5zFeQGBlsp8vnpmR1RPq
qlNlT+s6GKMZFa85gFZDWTto65jM8Da55QmymesMydMBzsZ7B8akrbXdMmIuwxvx
5VryUJ+AkqAghl1OJsDnqBUvimPCwTWiDD08LvZxiJftO5NADlxr8lEyN+v1Paxh
OALbagHiNHw5pWRxeJ1fzGeeQyiNZqthYUILtSD5fmc20CFmdsHcdw3tUurc7F1N
qi4rtmbbPUi89CPMzz5Ao88uA/KlyahG6/C3o//MrjfoqhAoXFkBJrARQzzcK2Ob
kk22B2s9UtbBANPM8xGlj0EEofzAy98dSCDB9w3MxujModTN05QvPPVph/zpyTl9
ab5+ny+8WQ8C/9YaE7eyU5rppcbMQ6Ta3ICJ342NL8+H0DwPgFMVaVqWb82YjPOV
m7lkVO1faKR9NWNuhIdBjgugsLtRBmf+nwfFcKLZME7NM6feNmL7WxzyLelpYsiB
Tmeu1fEJ1payHVBaDbxqbVP65rb2Wfu5quTqsBf5jaD5D0AKxgpOwyiMbzi4x8lC
KAl20RDrAPes+ptt+uw2hthLRwDGmDlBGk0AmHX7xpyH1bduoPDv/7c+TAB/0HYN
gGKDKk21eZGH851tzz7g0ztqmAhLSjHFOilcu+/irV5EU6X64FHwqspPJJpA0CxT
Z0mO22ZMrpZG15oBLXQsHzw8TVC58AztqKFgVhWYAziA/IUp0CVqAZxT1Tyll9CD
abjFn+lq0cJxZkG1y3gBDeAbNperc1XvTy5K2wg10wl+RPKAYiJS+XQUIh/ap9TS
3K8clRNFQ0OQmNJFhB+itpdzZjKcpkeZ7Xi5cqzoYAoYypONgJGvVa8UjzN+t5Ec
8z8cYkIriXdOmFPpJ3LPZAnsO6BwGD0R0bsrYGf1nik7M7uRUu5Fs+/jY43KLHVK
KvhEV+CP7KFnrPvdiKEtkKv7iK9awqt9ZWic+4jHwPGZM3vf+QJK2DwNz56hvRqL
9g/VAjgESYYjZplGGTD//KYdX3UnaDANR17A7MTkzMGb8ROkxdHNG7JbRhuALFzy
vucAD8UmME3NuWE9orNzLl6KxEBWre22nWbbaYEaiZJUxOJEwJDB2hHdDIYdBCrY
gGUAWiL6XhLEGnv5/hKV21hm7zJdNb01tloqt1wtKuztxVlnJHAZwD87gJJpDMXV
1pwDvvPouQ5sATnGM7fmrC/kc1Niu6hys4Ckl2j7dsMXahymjhlab6dV1oxk95ud
qtoq2f44mycmLy80eRqF8pBprjaCq6FgOUIIgWT0hAuBF1sdswVO/XvZXrAAELb6
OSAfsPpR4PaW5nd/hkSuvCfoUrM/uu+G/qbavDETOLIs/yboAyiX6t7i/nA6RrSR
VsQ98IutL9tu2JsjGFrvxpGci7LVZXhb4x+OLozsFGWGPBqxtgDVDwsqV2vadQBc
76qEpwdM1rrRjvbU5wpTdmkBOs3oVhSvmBJTHAsS6zJb4KW2NigSV+X5cE9jvK2e
9yVIou3PhuJBVXXZcb9tM8x4WkXA2RDeQdtAK6BPHBHrsagCrQnJQcc8sHtrSCWw
Y8c9gVC3cfa7YucZ2iESUCWpGFLB82Yx+SS/MtdGNs4gb5sCyHbowLhapftQeRXz
xQ6mdVtGfzoXvD3273xZMnu0oOrrmBWbAL8pQWjAN25zi0hieI9Z5jdZeMAXKSug
0SMAkSq4nN1sQZTxGYs/Fa4vX/xP6Ny/vyt/DB0Oxn4lzINeI7ob05Es9YyLW3Jo
EdXJ5cvBLFwgmylJYS22QV186V+lRGehu62F/p6Yd56xttMNdS7gQyq41wyrAfcK
mZZZV1LXqryg9QQOOxTzrV5vhzo16fMMiV47zgmpOX7svbCeiuWu0Hx0V/GpumUV
3RIvYRVYPYC0FT7q1mlP6bI7BHVPDGaAFF80zB2n7r8zZTZh27oZBPgFvfFvkO0o
T9b4VuKVPB9soGCZBtIm0BCZFx1szttEIG8hQkuByn2/qu3WW5Q0BCoJcf07Kwhb
HpHWccQkepsLmiDdIjps7N3vgQdz7kHukU/9QO1Pg/6XZrcX+wTnFLBdpabHrLAI
9GdLz8skVsFQ2hxQQmC5p2RDOY1I3CAOheu3iIO+gLXJtFBhrtEkKgwOYK540Ome
VxiHIFu9EFlyBfcK1MWnaaqkSzdAZ2SC032dx2MCzpKegISshBIRauGuNdqNzQXm
dMM4cOnhZelbdUF/0H1Z2De3ZmKr3GbDZ+Fl6cNOWBoY5IMoPfEWtk3iJfc71+BV
Dfj5HvoNFBXpQ03UqC0xhrK4N9sP/SHojip7REqamWElePC0BQQEt0DUa+hzs8N0
gilzp5kIuxNYBQD6F/PBBh1+MHy+hBwp6pp7eK0C4Os03uxA9dPMTr4dlNy0PkJ/
xofA8eykQnBS5OFwU4/XlyHua9GbjJ96siidl5RHQRsh+IdI37QyyjY5ULo31rTg
TJqgmJIpQ53rm7PQgptHiCDcx7MJ9pdyhAF+IpVHPhhJqdpAlgayB3afRDdP9nDx
JjelghAjZuq4qsq0hQef6UldFjpz32WC3a3/on+bJVMZuZrqZViBFS+Dy88m3cWi
MGzP21IC6vhBFi2YzrNrPQCkiwaKBw4PHOsa3PWay9M8R8pV5E55tqGXh6u1fzxe
vVeuJLo/bd8QzDQHijJ4TqGprPl0hCtNaT/js0uVSpcSdkI16HqJj3Ndzw0EfLVe
wS2gT8Bipx5dOXpr5dufFEjLQKyrm8QuRUmw0atSclk3oAFSUQssodUax/WAQio2
i096opwdIz6dZn/gobaLUA==
`protect END_PROTECTED
