`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AFdUu8r889/Lufu0NkFGeMkhTSTxxX6JI4u9VCPS+p1nF7+hMr0MF24HIQyRtrce
vehcuHdaybohXnjG7cxoTVT99i+QfmzzDb0a2FFgZsEa8vKPipNBWvfbxCgEiPrR
4X6S9JJV4vbNxOwPhjxfAwmPygxVMrq6F39fam6lxrISuQS/6jX1jeL/yjjIP8Xl
uku20H8nOCBqsPT6d9zuZqrj/aWLv2BhsOQwaQ9Gxoe58RCxHOmc7cu2sGvcv2hA
YJk7PFKnxdwZoFTm67Icy1hiutlsihNKiE6xSNLJln7tl0fNGD/AzruCzdn8rnVs
UXR9LBBtdGdAdEvDVI+CGp6wXahumTJElnlj6kxQ8X3CAsjNCzC0vWchp1s0Yko5
kXK8tjinDImwN0PMNVIEmVBkV5H8eLnHBFzHLMv9nm9I5vxABKtDEOW2Tz1jBePC
TczyX7D5lcjvjKHQwXeYMiIPX16/jdC0TIwzhuNkLNkc5eIHWFGPpV+ld2k3/LT/
uplM4pib6yboNnlI8dDkm3lbKOKdtIDXwMc1MpSeTVrvQGIwclGQ2ru77h0u2AxA
kki84ZvdMhFujlS+ZvWms0IzB2zOr0oNBLjbNje2bR9GsWjVOcAAsjA7L0z0uu2h
ERNcoub94HAvQ5lbUo6J2aNvaFweYiSCblYcSuFxUoc9JA21fmFY9shBKYzIl4gL
4qVZ1B1ktGsWCuThAuR9LQiVburJGTNTZ9SM56q5W1g1a5ijOuv1tA26KjMr2gcp
GXAn7V746BcL75sHMVLOTij5DfPLU6LSwg89w5SOk/5pUizL4Woq+L3vwYT33ubp
b1Q5CphY7Oo9LgzWXbqcY7uv4QSnTLcoPhE4ZlDhwjucR+S5ne5+Ng95+TofuDTL
LbNxHRPwckDfZUXiIkeWGVVO3DSomMj622boxcUI9fuRwc8UNH0YFjb8zCXM6K45
jWJyCig2EF2GLJzKeMolfdmQpqVUCuwYsCmD8Eo+U7ErZTeowlPZxzd+cVKuHwXJ
D7Lc+Max3uupa4pafTMUZhOmssJWpE2eVAzkXMu7DjroWZLUQKZvQziW2TQnTTmp
5oCgpGpzUq1wFCJBjjbB3goULFHiJ4pgabXQjWo5kcM45+e1JAD6MuV3ZCUNzA0n
qGUdS8gGLGVHuNOTXZhhrNbALFPpvcZUh1kRbe+U23l9qu71Xnj+ne3zLLwdsxlR
FS2/+LIuosObBBNQNROz/nrRK5ELRSTItHJtIYsbrAPCjuNBwwqwO7iXi9QUCR9V
4qasCpapn1djj8zHUmJqwW5pEynJYnBPNYcXiSmvWcj77q+ojjp6AFx+FhaomL/G
WTCMO7qey2oO50NBJ+zbrYN3X8pcY7mauWym5McZVHk5aIjilDnEpx51V34z8TsU
8CVia01BQsBoSSnuiH+9y0x/YPDhFuma5BjeaUTvRTosW354CQ7XAHRvjdqYLfeq
zEzaioIoCWDwB9Cc5/QXjsZccLqLen56ec1miwDdh18710CC3M1AlIQ3vIK4CQyq
UK+t8BBqX48gCUyIZ+EPa7uw8jrvTsmYpTMhAWPBRzcXoUeWxI28WdHRJtjeqoYX
y20ASKaXFbMQCDfbPrPKerAcKGoXTuSpi8QOhq4tbvjPcTVCsbgAhQ07ujnuC9BU
ha2YOIZFOXb44f7FUAPdb5Z3UKdc6BrUAtQxX2yirPqv2KAP+r4/DjZHnHsnIVKb
obrIlnSOfuo0XZSY/zdXSdRIMpvSsUlx2mmEygcBa4ClaXhjfGfSKhm2pzXKv6hi
nrBtGR5gq6RjGDxlZQXzwOyNe0+Js5TUbkksIn1IwYnXwcHPPA5nt8NQQOVoFsEU
JCeXc4CJfPwb2VMg9Y0k8wR5zQHYueGXqHhiENh+4hTXLgk00w6O2UwFA6EdddqU
T/JsK7F9YjJ+cq/aGxdjI3KzjDih3IVU7l7nVQ43gi6mOD3v1wiP3GiGuvDr6K19
MNh5Id3X8UykXFyvYlxx106i7iPkpqepPgn4c4s2LPso3DRqG1SgngulghrNHjAM
NmZ7Y4+WEzuZD/2VH91HgrIuXcQkZNxpYhJ/fWevkqV0+RF966CY6apR/5K3pygE
DpqW7ADlJ2OybiR+goLVJZVwiWsbnzCsn7IfMox+NAjP7XO1tM95vMLC48o3OSpn
kGgqanW2K35emJyy1r5NPLRHAjcqgyD3cWoYMOFSMfOuox7uS/MoyPEO6xQ+mVrx
jiIJzaH4MYjWZP1DbyaXb9XUfQvSowdTuIlTbe1/wa0hWa/EM9pkDVUqIF5sirw1
i5GBVQmhphkQiiorVU6ETP9RRjZeNuJTAkUbnPhXghbrtvgGvnLkxOCQBaRXDEfe
yAmnUM25Rv3IsCUqpbcvo3oW535mQobpsLi4jzfGhQ78c19q5JrFD+ueXn8R6VNi
O429qWcjrjWHSuW6rk9xbCh+a3wM0flQSlbOruoft4yPJgT9VIn+dD16Du3AyGVO
SHFxEyBpbL2s8J8p0/MsaVDuIRu/Gn4214Wv8TOgzxcn9XdWwo+MAKiZADgDsa7P
uJaRdy9DpN3OMEzxMu6b46AGZaRn+HFmCmWc9K75Pspuv9dbXmPxPpFJakL2FNF5
vvECmNBnHqcrSJdbqXQbS+0EBd16o3Qn+yJ/XKuONWmBFfTa17mi6UeWgMpoADMe
eTxb1Qb9YwwbivCMXhpj1M6/f4cYOKdTAafzmlHHxNt6z4fRwjktG1UEhRp0tYSj
/2RdUaPp0a6VHPVMimKB8vRxDH12LqqTyjFYNNjO5GNne0BkEtzjjHCgYG+ZJboY
UjoIMU0XdjihhlCPeuA93LbytPOI9W9BkhuXN4DLSH9jCYaNDheki5vKjDePHGfx
GkXuZtQRDTIT7FxBVGqVmvokVDXFjqc8ug52wftiFKHVHTAZQioFQDz2+wfnoqmU
V9735Eg9zMKmPylG1Pa+DiJuwEuZ8iWL2CpMimHqjTQ+FCBfkS6pNQxFNK3W9YXY
InFC3f+8QZR2GYWFdvuGy7XZuR9I13xuj2gtAG47mGGE9Yx0wZ+5yTmt2sK6tyv2
NMbkaLKySt0vWx5sS5C4Qev1BHiad6d73SseraahI8U3eGymzLBc/sGNykid5qUg
yg6uFV1WoSx0IHSInMmNqH0ksqfDebI3eXftZPZwhh9M7EB5DHRJ6eLHFYQjgDnX
LPNdG55/ajP1Ixm1elbxfsIN8ozdarm9qpmyz5Fov+9s5/5oIwVDNpHFKBnuenSt
CfHYbOAnGENzpBgW6+Nw/qVxSYnPnfVI8go1yHLTwvLcuFhmCjT1ryqv9NmQelqn
1d4LWZO0VEbxqkjSivh0Uz9tvOv9B4og3dEraR8m7m8ra2epdBnUXVu2LmtQ33+J
aRDVADfyQtNcaxJ3zu5Ib/QImajBdccroy0E32fHAlG1pD+kwmjeUUAwpILS7kdX
G9wh9T/Y3qUH2EQCfm+f/aNZ8r7Oqy2OGAaMg+X4h0INJO+sVXXJAcmdfbXppngM
zT0Yi7lM598ADTvvShiPOY+tQ0A5Rq3samduYJkcxxOp23sj9h8Yd+IZ9/DOZAH8
5Xu5frWm1RKtG88V5XolQtEE2+E9RT0HtZWhV1ODil2AzCeatJTHr0m6YoeS5djd
KHuvAQLwgSC8CtFnj7C4IFpo1ZuyPRz+wnGTMAs5lFdxEdDDIgNQ6g9Z2Z0bVoaW
18sWowdwXrNrTIVOKPVJS9aPqXBvSF8idagWwcUJjBA18+LHAKnRnq2kNpowdUy4
kLRGuwno404oOQxs2Bug4lj+wDvRPdfqKV8xtKgoEZ1RvcSD+1n4KTUCxv5zJY3O
64wPnFWsy25nPOPoms3Wl8hNyvbUK/DWb6czjFGrdYxJbKu+bLV56fm2oiuODuGe
Mtb+7w9PbDv030GLwXxS/yVeo02IXAPwWBDrGAT8S7Qt/c+1dvDRjxNpBy4U475f
YTZiBg39QUsFB5Fo7TsJHEwCxHQUrNqPMnQFl7mevQRj4Fuj9qW+zQrZadk3WjIP
9Ma/Kp2gU+EfBKdkG3NsreO3FksEfNNTiiH1R/y3qKSuV5vx15uuE3FQ5++QjuPI
5r3esTkB52NWJ4RbWCn1ClTYxVJyxKRpH+TtLrKXjcAEKnyPeM7iapQ24jIgcHoV
fdzA3a/DeATmzBOkoKBFaXzs3PXuVWks6tPYKt37EWNRh/vEQGTk/AcoVCJ//4/A
Kpx0lv7SkjjFCPegLLLC5ROSffcw4pvgO1W+gl/9qoN2tFbGaFAxUYFuV+JE2CyK
FojDQb9OHaHTluPedeN3Yf7+ecn3QA0cgMf5bnkDlfWOso/KJeZNplH81ZLOH2Pl
amkFYWuS/+NECdcEL1u4YXKtDG8WJ3AJPhSc19ujlZczNfIeZ2YPpxdt+Qo9fqwi
CQar/MemNhmRusxPN7n0ejfZ1YOURnKrDoWC6qqk5Ppdn+mR3JUkCb3uWaIFB59Z
2VsmlxjRr/rqTW5PKCwehVTUpD/EDh/4KoZOgTrrGLi+ugilFLaUGdKtU4w350b7
3pXY1xyK+TBqo4yLrpfr1LHXmmV2cGH7XlqaQSX308K3tOpq7XIscHXMblMpRM4C
M+Cx+SMreCLhj/76NDx78DyMawp5DZuQhqcnscdEWx2VluRQcs9pILY8NCrM3Mft
DSTs7QbzGCaP1uYlB22eABcQytqq0P2vGjrhgNJOLPYZfkuqlyRqlGiBTeC5aVBl
u4HCW24lj70T4u7tbvMiCZiUeSIHaWehypkahzj7C/sI/RXc1E3g/3Uk77pulhFu
IyvZFON3RMbPBtW9whPkjNaI9zNosWqH9monjBSALwOCPVqdlGfJcTuLCGbjyWkc
6L0h0m/BZJORlBSGkVm0oxBen0o55v+Kluw9PHrD1tO0Jru+wBF4Go/sn4SYPaWV
tbTpfftk1nk9J7XOMZHsqxIn4QX/hRu1zi6UlZK4fkm3CGhT3e3bz9/un1+dIMd1
3GpEtRCn3yQ1ZYIHuy/p4XntyQJNZ+e7o1gjJKKSyqEls1pNFkboKOqESHsBf+hC
P66C+vXv9hav9JhB/pRUwcmkUYabWztwWhgevdTCKnetGH1ZuZ/eIySufSh8KeBt
M3Xeju7jvnD/dBoPISqIGQaO0pY30MKE/7LSQRl7gABFDicb1uv8OUxmmaKQ8N0e
sCk2iOGi5VxOpRtgf3zqFjb04iRJHehL+7BXzPvMCQ7GuMR2dv8B761LU9V+ysKV
jRufH4VSP4u7WjC+XemHcBEHfQxvTmGKr2n8Q/SKqeDdRha0czNNOptHBmvYOhCM
0Kui/19srOt3mvJ1hOhi6Yk3g0QfyqZk3/f+VPlCqv6WfjlpKdUIxIjlAprSxY/j
wdwO/9afCkP09Lf6Pb7rDxB2Fkv6RZkePvOq9i7rAp2Mz+BaDXMrJauVK/EcT0cM
usCJV3BHxEOFIV8blJGuAcCo3B+pM0cd/U/B1ejWHm40ViGaDQPSjaYHW4ZQZFet
rmEJ9aK5Expq4l2lZ8jzw/TKWXEAsWqA29mVwJHDBk83u4WULG7q9tPkoRKUdNLe
XU0+VbPe29P1ClEGNJ9YA3j4pFjEvDdNP3wUR0dSw0o0kQHT1PJlnCes3HLKFE/j
GNBYqzK2+f4rwKyjRnOoU6Tl2HAlfvSURvjESaimiIEWF1dkpV6lwsvgrVCIT/r+
0V+GB13YeGMdkS28+vS+2YvUFzQFSVZzn380N3iUI16R3tPtL+ULTqgMDJKkCS5n
f3VzLBDbAUQE+HkEjQcfYIA+uQ2hynCJJbKiX5gMzi/9LVfl6LbLRglo7gw6ajn+
8RnGIY7/jts48v5giteom5htpP316p6kYxU39EtgXebJcfUZIk1nqs9vOMiDmtjJ
nfUTjVOt2cGVokWwcucw5BTkRUzHsyG5Sz91ZWDjr7Dehu1IUhLwzU/HoGb0V7LC
BkYiSA89D4Y5U2j6uXZcTqVvuZz3eAAfjgqBr9oxpwWtuHsLKb8l5dbr2BSrT8ah
GhiK/4akUyWT+c0Plvh+F6TQiOyfeYk4PQxSJaptwwQdjGmZ4p5QFjwRuCrxO7il
uOl3kHC6XR26HifpoQe9/kYh8vKxDY9YoBKkxV2ib5LmneuSUyPTV/EDtBig18uU
6expgwRUUDDZcgMmcku2zKIISTi71JKUJfSYULFA3CdDSegcaMTo/GPqDT45vL1f
Hn2q7KL2xGbFBX3OBEt5c2CG3OYknxOOOX8ccUWzgIgK+3Z+2RfL8UpoYpOx7evK
GEoxF9CRl8JLc397dgH5Tl/tnIe8Ji7huUhmk9FQoztGpMksbRpOZg7nUFYH7/ox
uAQeRohQp2U0yeek0nWp7zactysn9yp7kndN5QlgNmXP+TFRyljJ2T3fDvfwvIk3
PS0f6xvmxqne7mXiQRu65meK2Tue6BLHm9QtO18bWnpu4659Vy3ZSAZl8QGfce8t
rdkFMlheiqVijQfb6thD0pfAC47NElG2iq7W8tNHjYqCc8dWQP+IVOU0H6kemXL+
BhvzcDc1Mdh7UbD4Lx0IJrJZpLCnVvMCwUGm1svxzLzOyc+3HOkOD/QjZ4d5sPT9
Nv+AfF2Lwz9sSWX5g3fFUzyh1mJveSC/WTQC8rw93mubpb13g/h4OmBAg+iSTHY3
e2WxRElUSbojzxcrwDk08Vs7695QXZ943wgJ7tRK54nTes9o2hVup2E3on3lxe9R
bVA1f97uGFEJHokn98SdaxEDHoR2KQ8DbaQHjuW533wE6RlllwBxRVgHFJI10+9x
UZ+7o8mWqNv/zxMcOO30jGq54LVZmzTMA7BnTBO4JcMa1jIdJ10AqukSNE26HYNU
mJMjfr9z7vXS+QpUbRnIUpm1cfaoWbdNZphYFcnhF+y+lYPOjB4Bujs/0leRjUPj
j9SsCF7xrgtbEO4H7C6VdwKAcDrhbcU2v6cXyDR9NNeooBiJFg7y/ulTmqbNoZRD
LdcPxdAEwfPROyGHBohOETfSrKqQ9mUJMKvusyYGbRMOWWbsEShEmjZ/2QA1PDqa
ih9LUoifA8o1wdisaopmm++Yr/gS7mbCjCd3eyhDpmzyjP9OeL1V7Kb1qWeVgQ5c
Wx2YkeIl0u4kn8q/f9VMLCLhmSIew/pHH5OzRYzzjh2c7ju90vUQ3+rB8dcoqyc9
0de6JK+oi31Wld9bUmVSWXpfdK4U3h5pdMhRDoyC4rRklipHeZvuNxuWRTyCET9N
AC2KclGSm3YX7tNDcGHHUwSryuFMfybQhJS3Ch/Hon2vtN74tRtcziezl9FtObpM
LyWwut7VQr/nuOpDkGetNjTFgG3fHVGrMPEz1OqvB29prvyUQDt4gVhx+4HLIgrw
SpTQZH1QLgbIM1RkJfOqyNg6jbs+NoUZu5JJ/rK50H0tmLMU3jUqvuAXiTUonLeW
ZU9GC7yVtMUvkdTSU2gcd6TTtM5W63zryLBKslcdRhTlMSAh/Ohg4wb82Eg9NzPo
1WfIhjJYzsDAhUtSnA7t6ASVA9RGR9SlagblQMpCfNZtD1jzHUJxcz+ykDEUAFA/
rdCfvGrML90oGK/5L+rUDHBtPnHrkleqRRZCqzHW4GHgBzNimVHK0cKai3qe0DXs
Kk8Ar2AsXQkiDwUdTRht4gPPklf3As2IIGb2SMfA5ySXFv6xeCtH+sPHOnr5Btg5
gcCnuAiCRxb++YhONpIT6dVat++Zs/0QsaI1SeTmZ0+ftmmV2ES+8WkAU9XsL4OH
qbIeAwgpRQqX5ZUvwDs9UdJHuuecMOK3m4E19ZliN4EXkaN78PjPMY3QcB5CJZkE
4TcORC0pMzlV7Aj8vXW8tZOhtlMkaKlcK0P+kS1uOw04vFlgtcChrpXF2zxo3wxZ
crIj0srn5Xp+NbfeNOI5aCd5vKZ7aT/y5s18GETnj5iHyr2YlJkP1g2SI+guQCVM
u0gIhJdJfuwxAMEoVfNamKyfH4UsHnwM7AHvkcN4OTHsqsR805sM0BVoRTpWGFGZ
X39YSRDZoQGjLTLDxE1ZZcc3I7Pp7DymmriQ5NFw5UvwMOYgudXK6VXj2iX03Myp
q6NZvXgbPJvD/ogubreWssigmEMfvKtSV8nz2lLWOuot1eD8pnYCHnMei5TUwvsk
NTZMjuKdeM271yjA2OgZduL85m7dZDuuSQsN8Teo/KSPMhDM+PYToRrFB9VNEESN
joaqvyn9Q7Kr2+LXokr9DNo0JNpdZEoSBN0ddOSrI4yVt9sDRPjfZywf/mHHpj1d
6CamzsZidCUdGzoFlWdC16CCeKEvzC3ayuA6xizNMc75P9iRnNSzIGbdkQUYmVG3
pSBpE9MaSt78aPXpW59JfV8+L5JC1cREHAYm+IfRz7LEwYfdtcjlyuAauuHZ6Zgn
Kmb2jbUcs6e5AFeEoTDQVzoWNhoUYqiUjn+6hkwaVaQKzXMbwEGiplqdNO+rOAoZ
IiIeUdIAevpDLg95Pooe1vqhODNRjpezwJKI4d04+SuSOtqhb/mFJUo/DO24yt4k
n6TZNlkmuhSW6ShFttsfeWduwb1H2OEJYjy7B2WxQ1Cp6cPg0KkDYAHXD7lxXqSw
mlooRpXt+IMKLEvSegs0chem1swSnLgkSBh85b7HLA/aCXdjObNAIYxi86xPcHiW
0Xba3I+OE3gJTCdDQYtmQe9jqBbIe4rgiLq3gAzAjmO1DJFh3bQ94gfcal8/RKgO
WKoSAvkjWl204jlyRQWZit4pgiK7lSMzQazcxbrUfE71hwY+uZKvgzXXlFJKo7+d
Br/0EKrrwixLxJ9CkejSbjOmi+gztenmlLWX+MN7TymKg1lonv9cHIGleWdahTuM
+Gl/vzB8k7GLY4+oOnrmohwbMYbRT4bv4tpR8nVxwXqYzNHDg+Adqu18DADH2NlG
QV40aj8VxolG8Ys44UtJJqsqaFJTimMFyptG283m/+Atu+6C/tgdxuHgVjlWdDhJ
g8TXdfOJ2hXtePBc7iThSKjMLGuTQ0N7w5TdL7H86E+cj75ZfKbv8GC4pe0/p0iN
8WJCVfvCZWrK1cmeoZkSaatmvSO4IJiiUWXdjzc8h/UnLgyJmeB80B9rqMAKqFZN
oNx3tdunAKrCCf4uTTTSBeGTFF83/fFnHC2kw205FuTjkAnaZBcvR6Mdh7tNR5xt
OtGetHZJlyyVEIzF5Jk2GyHmcRx8VlAo5jImPFDoBZrLVq0KifIXHkBs0XnLVcan
LmvQDtT600JCQAKfxq5R4rXmBwineMfV7JFGOagqJQcX2Ez8PNEBz4aDhPZeuSdv
`protect END_PROTECTED
