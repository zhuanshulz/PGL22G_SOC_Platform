`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TA08xx8nnfBlX+lBVtQko5FbB3vSjWAQKwh0sQA/HNQ4hqPhdAj2nXuX2VNHjYox
jvONlSmWhXu+ELW4YfmrnrVD0n5nZTwc7jrfx2fXrYEqx4MYuMKMLJquHFWTBf0s
sJsYLsDfcBPxrYjb2qhRH5lcGJJOAOOg3zyAI2HWs+x2VDAtpgHRZyxHFcJmKt6E
jlsEptEAW8DbIImJFUNqBbCjnn7ocKpJuJHrFOoiMzluzCgDcMfBHriLNE1bGp9E
7igJcJ3307agKtZFz5P/zQ==
`protect END_PROTECTED
