`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PN3IRzGQGTgqeVV3z899vVBLVYi7alAPr6gXOBnit5jrzBQr3TRtfh6gc8o6gKt5
WpthdaR5v9DI0vet/KELg3Vdi2R1ZnrZSvMmhpVSERyuqbhyPaWFXGPJEp8njMFf
Z2XKwLVm5A7JiOcxztJrk5Pe/q9vCNlkQlvDp2SjUIjvDO+LHaOLKmXYeiFBbZdt
kJjSpx4bKHR0r5xqy80uPDhe5IwqmjVVeyoaFLpchpgON18gbHb2d/fxl9ZjVALx
2nAPxX3Xlr53zOrjCHTY5mjI+WNjJ+9sBnB2rBmqoXkdcmWJpO/olJZiyB9Yehbz
zUD6d5STfYNN7x8gEx6JXlaytGBHCvfEsvgPT+7d1Hsxrm1KyZLC4f8FXGbWrEQG
H5+YUVnD1To33ak6QV1ImKxEqBytxKB105B1NKtZTYUF43TTujcWUKntwtcyggrT
AvM5b8IfXizZiI9+WshLFYNMbfYJ+1kV9CsQLXE+ll4kuF2R6qoV209FERMlWC7p
z9iTqAs1H63/l/chae96GfLJPzDq7aYbIJm0QzelT0OrYR9CsZAKTGzIwesFRYFa
PXc4pUNgh2j6RoPHubnW6w==
`protect END_PROTECTED
