`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t4SyK+7BRh73XrOjvb+3leFgLq75/T8L3NUvoygrI3ztfTJ2qZxWUzJk3h+FhHIB
KbQBHs1AswT/0FWQjz9BfWDE02lcpFxc6J/rv5auPGL4Z5HSHY5XTpnQZVlfr3hQ
nOVcF9ogpTwWP2dYVbPnxY1ZLzKl8sIuTqt89A5/HsYPputXwLzbdpJE1LVD/3/B
XpAVzMLFrTJqq651O8J4MTxd0Gfh7DYlP++HdxfSm8yfX2zhMMXPtYM/1TYFs3CE
2CDsQP8n1aXVE9RKtKLI3RmUIAH7pXxpSDPg3oAiU1SF5cN7IpYg/hPKHD5UYILD
eDzpKKs94z2KSoAtxcT9cufNnaGvPqZSbVWWZoD95eR6xSH38CUmcssyWm4NJ6/H
en4KDi+9YKlE/lxlqw5c9PYgz+g0DD10gRhk8is2GtxK5A1o1GQN8Upf3iE0Ed2U
yD7i2Jhes906rcAjFxc9LrFeapnMG6YgfC8LGpP7pBQFw8FlZ6QFksYVZPKrmLKX
tcASLsdfEQ5QDH8VoGD2Kw==
`protect END_PROTECTED
