`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tTWwA0KbwGTaiurILgne/HKPgJzNXfJZuUPSTaOmce1J6ESgRFDWtov588riLFbs
ySvoKxonzOD/LO097asC0LFR8ZJEDoCxKlbFLReWlw2htFcP/CTZpFgPSS6v4ZXu
6FktO2gBbDo1bc+RtDD/i3IKUUuj5uGb/Ut+6KfV4Sqt/BpiGDeCYIWlINaEZZbf
emPdgdifEoKK523gN6wvWa9lbrpWPifN7LaBATZpJe06etSg5lofJFrvhoKOKcol
rZew3sMbiuKf3z2zOli40+AcMjY2CQ72l2Kvlu+h7MRlw1KMzNBrIXjEFNLRz1d+
Ed24yDN5Tn3yMNI9CvX4ZMbLFsrM3OBgU9qcEZ6W9V/HYR3h3ai7msuNYxoPGwuo
HOCXHvKzGM865jQO1JUPKA==
`protect END_PROTECTED
