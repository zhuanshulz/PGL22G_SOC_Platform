`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rleawmJsCzMw1zIqZYvUs0OH7iL+/ZIsX/N67tZ8QdVOTmP9my4bboS74s1G4+iP
T8FDJDIeMGhxHUa8osnyS7OgjITjcuKpk7P2ygVxBof5xalJ2CNRJTmQHKi5LQyB
EUr42NvyQq3BCDjdMEJTvmCma/JGbiPjOfWv1gE4CUd8yJc33O6B9p2kPpT3ZdGL
99YeOhoVxqF+sYXzwMXDH4oVe/H55/nzrjcVe9fK+eoMRdOhtQYJjGVgtRb1z24w
E850I2v6Nhd/tJIWs5Vwco/E2uTNjmWzLLaUtQDl7srsprIP75JzpB6O2qw1E1sp
wHvF+l+kz7NgFxvwI8RgQ523NFW3T0+2Y/gv9ethx1qZlRDRTAgwHVLsDIqjsBn5
hY6jvVa0rPXhp4gsJPERNbRP0L+FdLn91mJ3qxfjbMIjpilM389EsChxmsUs62L5
CQ9StSEvUW/wHMqZBTvUhKay4da3rh5Wu8gcbf82/5awcOb4PbQkX3MBYYJVWdOG
doliFyMBgSSBDRXm/5RFwh04JaK+K8g1Xv7qihbyqP2tDO9NyFFiApCOF5wwWGQ6
5C9cVYRJSXj5IOO1HS2+SQJcdeMg4ScAPFZdKAYpQMmapglFB57JvdKQP+76XYRw
G60uPxRmbvdQbTCn8ibHqTSwtNEl9g8vkN0BYzdOMp2oql1Sj/htX5cZfhTIwSEh
osLq7lTzoGvOkFBZNlFYuc84uhXyPgugMG4QQxHyPgFfqQ9xLVwSSfVRudd0Sfbd
YZBAoJKNGcGDDvTVGM7oi9hY9TVtNVLUmG07bE4vkXR1XkNW+K/gC6YCzNfRIr6b
xhfSScorz/bdJuksQNfg9d8lGLowNKYmvxVZfme5KDejojDIn/JwoBYcMhRQqK0J
nr1DIqpkT1HUuG80nw/kgKL7GQX4QPUiCSjzjai9OjUBM73cTUgqi6SjJGOHmimD
Yt/P/ekYrFmab1tPC+5c4omxu0tlh25zef314NRJ6ISF4E8fgKQRRB08DoSUK+sS
bSNOjftnZ/8HwLP90pdjxA+Xs31zbhImm7TtyJFgPDLfaBegwZ9C1EiHEqxQPFtk
pRSBg99k9WL2qUcuN15ckIy9UTERiMygVUaAbe3ByHCsLSBg6s5/jjuBzpL2BFLo
1HVi2me+yOVVytwcNv5gHSp8ETm9L8nozWKVYmbgg7/+NFdb9M26vGiQznweWeBz
mOqDl8nCKWh2OQSlnZDUkNka3OmEQYa/mdJbLQIsN6QsVqcQEyvOndKDgv/OswrG
eiX7baOHBQkGXchWM4TMtTjX/5Fj75UUCYvRqubQa9UZGDfTsh7ljcyL2b7I6V7p
HNY2Ep3vZSs90oILV4c1P/xYHx8j7/V6viq4TVk0V+B5AMGTaSwlHsjIObyvr/C8
FihghcJA0v/6jYj2053ZzsXcheol1jnVpp3vY0oV8GP5UkasQn7KL07OXFpIJ8G2
`protect END_PROTECTED
