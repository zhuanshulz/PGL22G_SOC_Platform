`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sq2e1ri44X6hB2/2SuWQsBBGG2hCCxFkZz1SyLj/XjlZfTGDeEmNkNe2arIg3nyA
1MxGs3esLwS2shQHt8aLL5LDfp+aTQekKGuK1xwsloiht2sPX1L5elHSzogp1y+x
bfhmIxzArwxAGna62On+T9+BDvRcsSlVVSb+LWa8wZa4FBbfnB0osK/+oCBLIeMN
TfoaFdI8xswJlTPsCi6nqq8OTkqfTrTp0zho9/ONc/cdj5vakulrbdcx58lizTn6
oUj8OFJs/+LveMYUFr+Fwpg/zVn0m/l0uQL0PYLn+HXTSxqh77hmTokH3iOsOjRw
B7NqrJI6MKly1xupQVN+MaIGOQc8KYQhdIBffVV94FRsCwYb6Xiyd1BsvMlhdRVl
UqulVrj8FOf83Skn9q9/gBssZYVjgj2vuL9K48V13Y3PUozkMSiTSMl30IvPOQmj
1arpiilNNAnriEcGrz78yzQ4TcPdYlOdzQm2YPCgm8mrG3jt1JLIU7MhsbrMBtrm
yJFFtXWv/v2s4tjAbWuPFOHLKd1HBceySLzUFlXKx7+utaUpL6u1Eb1m4EyTz78F
uFhhYI7d9uipqORPf6DbqcqG+iEYe5gxEvzytkpI6oB64JTmngKz7wWFHcCcz0EH
2AcedOG6WsBZDUoNyJ6A0s4ihzLicD79PDCE9IgRpYfKajvZi1cbJq0ecl8JLUQM
ybYTDv6+lQQLmQQNDIAJeY6/Ss4a12slE4dna29UU3AEW5SOTOA9nc6+lacY/W6Y
L6kbCib4rvsakvWGL13a+vLhyWOQdUJjadrpwOTZh7Ewe0pxZzaawy5sMel2r44y
jBG9u5SCDzmXfKTls9ZhILMq26G12otNnNcMIE4jPeFi39wHB/whslKNYYb0355g
vqT2pmGbCLNqtqx5S6fnWrPhpo2wutRHr3tf1ch9Cj0iVnXlkQOjhIeEeFp4BxoP
OmzlMwO5mpxZWpZSDUM1sw==
`protect END_PROTECTED
