`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8Sx8w8vjVRDmZj/1uM4E3gXmj+/uVoIZcqYC/1Dcrkab/MM+2WIKaRuppC+0VqfP
QbPOa3ACn1cK/XmskomeBQMTWMVVyHkkaFXMR2TfqWzkiiuN0WZ3PhR/8YHD8G+K
XPxGsZSoWuyVyEhFX4y/0E0dAhqtmUpJ1f0D8DFbPkDlxFVgCHV4RldbPFfMKEXX
b3MLleQobrgDcr0NWl3bZ0UEwFUcWyDlMJYR+KWExYBqVStnKiBV2VslHoM/UEh3
PJIGq4MPr6t6NCKlOShcUORnlVTbmkamyZ5qTpvjsAbqL1pd8jQVGGskfWsP6J0N
kCSvEkgQLqYwq01KK+ZIJZrljsprRPgPINRhPhSThraOiEX+Z0ZpbbZHgvKDKJOo
Rc5SLtlGjGAYlvQ+9i8/vHsJ770EsbLhII5C5GE598RodWCJ5eNljXgtbTgPSLrR
us2XUFB+4yiRML9jvdpyfEfiJwHykU+LmQNZ7QmVwTvYPmsoHmtPrx1YBomyazZO
z7zVdy3JAbHv8YKPy9V4iAxdwdYsgDpG7nTvB2t/9cicNRT7p8L3zrzfKvqnWlrS
nRb0W8FmnZMuAw9SwxRMKptAHZlGxAzyCRGjMiaOvr26st4JBrYPxh8I4x5T6JfA
rdyB+BjKOxju2IiD6vrMqRuPij1/TXm/hkc9ibzEu7kYOSvqylP1VAL0cAbFmEnS
GwI3vsFMPE5GcETNWeD7lm96njo33aL4HIY3KVFEkQIXRQ90m9+C9CHdwIPyJ+i2
v7VCFWCvzXZZ6+4Zx1PZapQnPsTIBSZF6B5oSbNtoTaAa7gGGLYPWsH4oAJ/9Frj
B6pEsNk3XxriDPg/y2cFiA==
`protect END_PROTECTED
