`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F4ejS2OaEMYA2GL7a/39aKHNIGqgfJaZESkfDj8XxrWnnNu39Yeo7oALSdxmaHKI
ZlxwoJTDA/T6u1m2jwChUKIB8G+StXGlB1HgYFhZ1RI8ocoedLoyZKBEskFV7T8p
KNOcvJL+IPwMDKDqFyb61ZZECNlnzwXvvbc1mpF2d6MjgfmOS0ebc4u6IcHzZub5
xykMj+kzRBL+hSAxo2JP5SaAtN4EEYrY28lklw4iCwq8yF8/caB/aBpHD/nBIKc3
QoI5h6VoGLyirc9xLTuXwTSzkkINZ1Ojx7AIo1aN6jpjwOGDT2m7YqQIw53CeOFD
eAlHRYvnq3xPYeOy/jBbY4I0IlcLk4TyAtk9w4JkDNez7Hpn8R3OhLCFzotQzFEc
H9msnSokBDi4iboMMhWAIY8VkvFgITUW+oqmMKiUloYFrHoo+WGi4faRU7gZaDPr
sB4r2HzlhIPzX2cPoGn3/99ZtRaN2UwK9Y4ZmN8zs6XcJlWgDrqwscbsxcZSlzra
Jkzx4wW0gvk7UCMw7AEnrLtHieie/K5/LGD/m4ImHZWd7JPkfqiSOq6GL3pd6eW+
Ji9vyWy+Z/8LG3enNRiAiedrEQ1NWHCmqtJHvp4qRxNHoZTPGsiBJ+j4mJ2h/d5J
DHqUwlVlk4yuygjpaVpPorAE5F0dd7TUys51d/XqL+ALxOCTvjmjenyhhh2kdIEN
/SHHtdnRHrxhqllGy9b7fPCs58LMOdhjIP8uKwlJOIZbu00DJXYGEt/JSZHoDuX1
1YvD976kJgFK1SlJnCNEbbL9Ap+xJAgbv/K16Nv0SvG6n5FZ5q99uDJtW64FqWzy
R3TQxw/Nn9PRGVMVZn61JhEYfGM0LTyh3VWP+82G6Qn93g0fqbxeQ6nIM1L3TQ1d
lysduSVSilopjj3QpMJojOgiTbx0CjfTRg1i0CqTyPWDSBNzgKmbqOya/rIzgfft
pi5YSn+F8g8ICc4NzlX2eAKRAzYKwW6Zv3GvqrviYhmOw5sWaqIQ3ZO+DNRdQlIN
xyfBq+etznYyDsdQgZ/g3chNGstVx8uKJBlRV/mzfj0XC9eZ6FnTRJA44Gn8qeW3
8gIX11Bvos7PobLX1cWIZmIVgSph650eUAwHm9axrao=
`protect END_PROTECTED
