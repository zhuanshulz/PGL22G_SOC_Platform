`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/hG7aYdjJ1e9kKrAyKhpjIBoQGWyk36qqOFXOCLI+UfzYfx0n+mXuVKYo92Fm8vl
z3LOVbDDaKUGBNtnj3xLu4gVzM/BBlTbbl3eZ/qyh6FstQbz8D0wgB/w4+IeQ7bZ
7b8rs0B320LxGue8I2CivjrFk/G2u2SdN5Mg0NesWKRvoPLAG8zLsEJqEcxaCzmH
6/mL2WGGErh6zathojbAoOW708n14u9tr/XTtTVF8hAiisx/1UAdDtWq8hTPbEPb
YX6BRWGFNpp8UXTUttO5YlGOtlfVcvoEXoaG1zeSJxT1L2Y3E3UNCApxdnrXC6X2
xV60EbzPvH9dbG2UGxrER8H2VTDbOnks/xhwXIkF3fPgyznfU1kTPYKOkfoitOhx
OUBG0gc4fJYHp5ltp/3FrSjmke1rLFL9WqWKxFZvBtmIYXREsbY1nBZdvraU/OJt
tA2m58iW4nIZ23JZ6zcpmBsC26TGLHD8cZ7YrHRYnXbDLj+7hn4HM8mvmHlPYsVm
I7SkcBzdsH7MAlr8ARlAW0e4Np/wZlXFpl2X8EE2NS3by6F+v0nLNdW3ej6iLYOP
hl1mTBDGu/R6sStBu+p310lw8jKjOj4FYcrMkONFa40Ed9DiewQMAZwtrBjHLUXa
ysAHuHLAtOJFxd5bkOsatXa52Jh35xCBGFR2OmP4tyPd9+Eupna4NFMhLSqVjt93
OuWdzTeO1POO2cAubE9NtHJXseWxh4gyCXz3Mnc/7uYDb60U1SWSHhuZ6Ra2ZG5V
Pl4MBtI4k125tJUfRX5KkGERWolUJhilEo9lewPB+ScY/nMY95vexFTfGCmvp8vT
Is6TUN5bj1aMQ0AlPeEm+IHvkZVmDaZUAhuGnepKY0miA4YSJqVIwK9uhlOEDXe6
y9hJkQtGrXE74xDOCYr4dQs/0sJ49Az2Rbw2+Am9Pc7A5HBXEZF4lRZlpFD9Vsus
Job4kvVrtqwXXC8/Wrg6LNm6QDca15ha8BlABSD7JTUQVNW3UFq3b3qx8ysqfHnW
VPrNXJMi/RtoXg5/oYtEBE46FSvSzwVnF48DkebkEOr+k821BpsX5AonvIvMa+ZX
829i1WAaqsa1GLCoQ2c+wDCL3rk3FHviLKiH3MJ5mlbXCG/vfcYx7hZna2LRdwBf
39M0ULviHGrBNorVErgk0N3tgunn/fRhRQAkkd/SvGwTUZ+YO4t7kAK4L4DQBTgw
Y3iELH7RfWyTB3jgGfaxA6s223mQGCkA43K6p+B31rm9wMua1kquR20nDhs07W4B
Cq4nfTyLLo9T24UYlrYMBvJxG0wnuUu011IrVifsktjnggw87jnDU9zncfPMJER/
/TN4LuB1OqDv9dFfwkee4m4vO4LPnvHt4QKXdgy81/pWxwnYGXITwmxkg8S7Ukyb
ww/Nq1oc+hz0/M+AkM4/CDT2aTiAEwUuoU07cvNCIBJXeJy+nnGkSY9vKIDUH+2t
K4WRV44CsirCzbQ/hlKAZhwbe2lIl5cK9rpEo62kmMon8o3OerTutpbW5mEN+sVw
d8O4b2aLiC1Gv8zcyxm7zbTpHiOU5gpysMSIam/9kY9FZ9VuoeZeHlNvdVEjMcSg
IGRMeEeaAsMe+s9QQxgmP0gyU71OKJf1Iy9mokgYsyof37VzAAeWznXjeLXBo/0E
bO1HtGcFpz680x2b1JjZm9jI2l+1v547kN+hwR/wU9L4osYgRDXXfxlKKc9cMnFJ
cVsi28/YpVYv9VXE6HQ/1V8UTo14vWOMsTlQhPlOG/MzjsqX5blAw79frQ4lh+3B
HjSA7fyCZRkVtiLf0HIs85FCU4+UoJoGH9v6dYpXa6wwXZDC+H6JUKIv10mrQ8WU
pzI9erIf6jaa1TGrl5Ls2w3BX2CbsA3TuXgQioC25GiyORxi+K+/6fpPrC5kcQnd
cqC4qZHcFnk6ztC9iD1RmnGf1OVIoqUjWc4jJRJ4JT5+1IkKNitsnr6Zwpb8U5ha
w7CbmBhLf+kdSSJ0eUYWWjMgSdWeCrXdHysh3I2QVLjDSRyLBLAb5FvFf1ZnHs2+
q4H1ScTZG4qqr55yneqsDyNzlPHruI+zbRbe9dhsiGiCKddcR5RAYhHgBj8M8H8I
2xRVWFKunSrPfsc8mE1JXJXldKPHLdB+OCZEyHY5+I31VpdLljys6/edrcu+V8yz
RIdad7rWfzb6Jm9Rq/kE8e0KgIDa+fEZKO1/hYAnOWirzwIjQNRTGLaNzZo79Z8M
RJVwg0A5nP6Cbj/pHd5cR4XZ7MIpBdJfx7sPabBSbyLgrL9v2vDC9VjZ6JAO190T
lnqNToBzEDS2Hp4R0Vx+hEZmslhiIsVf6C8etO1KjLkwbJdgUi2rrPHYKJIJJdzs
atqT8NaeCLFtMmE5NlxS5Abn46SkW9l/bQfJopctXCZfvvY55xhqx23aZgVYh1oN
NV8UOGXaD71+WEHktENI2bh+4tlAhk+H5W7pDs4+QtYc9kXTe4fBaKe/ZkStYzWZ
Ibzu7jOS3buqq8Qo4XppqqVlp7C4tKwCGJ088VDipeV56zmnQhTpdA4gLa0HEAXr
W0PxmuSiHZuehQBFNLBeHvaZIZMMTpiPhugzyzZShROkm6DVnCaQ6p02QgoqDWUM
JV1Xr4zwnSHugPwpQbdv7g==
`protect END_PROTECTED
