`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+s6nMK6vCQasqjc1bZ6jBc3TyF04rRPfHX8/l5IWhcfGicMU+JL8AQo/OVbduzOf
sBlb9uLr4NpZ32h4WmZTGs/Fx/jusrKFqikzsNTYridLJLjFGP0iUrYEebFaCIiF
5LGMLyk0uKzyoN86+XhA48e6KeTXsQAIKtlchMQEaD4sW6SGCrL7v4WsLTy9wCuw
WxBaeo7TMsY74Y9pjWfDXu2DjGfjRKGnLBgY3wCuYmcubffu89qhJ9smFGWExha3
g9sIIkmZS2Z6WZfNwUKgUvoOOlNXzUfpL8xrTC/d+iuWEjA78IM7yQVCHVlrF+5G
8dai4O9+KIAirYYTsvBxJCcNGHgPNAdK9DFNiUhaxQWSeU5Do83mS6/cDxxOpNLD
CrWvLNHL9FXeb/jHApcplkfdn4jnCCnp2brfyYAKyQNtJ/JQaPJJukEYAC+Cj6cG
PeK+CbUNsxvaorf01qEQ8xufGkX9a3uOtPp5BVgBf6G9aUmC+XYeJHe//bvq7XmK
J56NFdNCVmSyYYBco7pzbbv0tQGoFSv/+f/nQLQ08Nn67xXHxl2BJ7wjiJzn0neO
rzdKNHIuU2bpiy+EH9Yiwq23rWGXk7KV6cvGpb58Wc6WFG0ZsocIGvAydSWih+/7
VG86If2xuonJmVxlNZ/h4Q9UAfQUSd9U5KBTdd9bHXdSR6J9TKxnTuT2wsmbTG4c
O9FwEHym0UAkVZnt9A7TKBVjxD5OwS4XIjWE3nYxWZ7kAgGX0qSkbYK8ALUXgxWt
TJ3CjMHYyftv5nKt114qLOPYAE/smeNLBO554pYWTWyO/aaKt9OSu2UT85djcQ06
`protect END_PROTECTED
