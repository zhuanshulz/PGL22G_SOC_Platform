`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aMI8/V9Bd+teRAxoyz26PPhc7I9cn75aLKXuFE7ONEefNx+oVt8YDCfnwTYpLlOX
CWWu03YTDLZdRVmdKyCvfII6AtggdTaJJfjOjaiHxnUX80dwJU4DgtQKOjj54hY4
xNrAW4jRT8UmI25Xc5YeIJRIvoNRYO6UfMB3MX20XpcLLxZ5kcQQg9+gXm4SvbL0
M2SrXBrCdh0yuu253RcxDnJiXH+ei8noAPneOCY8kRM6u6vWNlN2ReFuW1ShWhQx
FI9o7p8uMfJop3MwTgirAxFD+pKiY/FtZNSt2NxO/1OQ3FyjhWMLwzGAYS4WDxbR
9Js5Nd1LqYrhdMpMtmFNBnCS31/7l1UrI/QSR1p+bru2jUUNGjb/Sieh1wG9DG/i
58xr0CQVpNMuAVMxUTTEbNJe31bcm8yzoZ0n78msy1cUm34EacbzmO2yRlUNCGig
DWdszEUi+n+M621JwfcqfKzx3QGMg/ggD+E3NPbMrfaeZ6dj23ADUGCI/nKxHRGJ
sO59xe1txcNU1VK/1sSGLUIOKTWkeOJTUkZfXElncwKjpmZCrxZfu0poWBAGfFHe
sHAQV1fZYFX3fxBQm92CKCqEKYI1AUkfZVrvlUoJdE3ILOKHgEXk2eYq/opRfC/c
FAF9hEcemx/DjQ2EwrGbOjqhl56yhEzVouspDRce97pa0D/UkbzDSKpuk9e/Pzgz
xPsUiNvTxwzusmzCXnEW9tE7Th3dysjesLgkuRWEbnYsxVzJybeJYsmC3bmQEyJ5
dohBZRORfwAAfTEELCNCVCModsmh+G6nV+YpvNue6nnCQQ/OCk72G1RRHVQ7q7HX
VKsgxx+jzoyL9I0+dTGsMeEtlC118BrWzjwyr4bfuuVks9TGzMuZXe1VuoPTqqoG
d6SDS2ot8OIeN9mAKCYrLFHqEYCY35hgTApji4njSH6K78sheLm4DFZGAguOugxI
Jxw0gYlfcUiPD2gT3q5nM3XFScmB9FpeVFNFmkgPoywH2rOtPpk3OTIOCC60K7bw
yBxBAEcrjzolLrT6c+QIajr0y2+2+M5BFMjqq052Gw8waJwI86J28LCvJI7VkNaj
GHyTh11VkrkS3WM2oERqPHov9EIf0qFWQy/4tNSFw+ZlIAwoXdoH4idtLFN4+wwt
bL90u/WUQ2cKHCgxbVL1gR2ZXMamWywIHyFrUgjlup8VmLC/M2da+v4b3PWp5ZXc
AFADXeLAjNyXhKV/5ceMx5dXjVq1WVc8eM35au5wTmsiFBGGgYzPVALXd3JO9f3x
rbI1P7FQ89SHhoIH2x7irj/p2pyqPX+tujIAw16QErtJh+TtC0ygxQH481mysXko
ophIL9S30fZsuMk2//Xd6AVByAEMrxAQ1T4SJtdyg6yR46+PUp+uXJuZqNcd6CBm
w9pzDpC81sRumkw8MC4wChbl+2L+3oiSbvxJ6VFxkIAnXm1oADSGY0M++xyKbwxN
4ktp16E9Ex6zbF+ZVsFRZES1KptrU8Dab5MY6qJ4otGAcRKgsRUobtg13hVuR6/u
RZATqDbHRyRhzlnph5U1o2T2ZkMImOYgWN9TszUHxXbORlEYvVOPUKEEaBoDWwkf
gq2f1yZ9Zgk//OuEL3oisR9wbX8CVwbW3dCu4AEywHUowBTjkUOJIcdHwVXAvSsv
YOteW2zNTg/6I0wBLl8htDgVg2OsMCVzncO04lVDtUE2H57yD9XXc91f1qWle5mb
Vs7o07E69dpuIE141FGovWvBvpVBS7PWtsKxggzkhbXjjt9K1+AOrQTNi8Rx94Im
sOcCK4AfFLQS16vzThsO+UUXX1mDSrkJcf21aeRA+ZYlWu0fJRgx/1cG9N5j3Ypv
dE1w1pyXO6hZ7t73QrRWXkZ9uRrkJri5rB2aDxQlqTDq5o9j9e3GLfo2TvIkODSa
zM8gxzD9oRSllg+pHMsrajw+LVXfaezGzcmqyKpAZygFEPeolKpLQBDP+Ov9N5SI
3gCwwSCVnUwATMV0LDBfMWeCjgNeynN4PEAPLE9nXzTD1A6UgbN0VwmXeHP9fJ6G
w0K8i3Dvn7P9Mrz634Nl1lR6aHBtP6c+WJII0U3Jql09SvxI/3f6WZ9+6B76/USR
iVaIvwwxKFEgso91kbIsgfsC5DYYHMUX4ut6ah7gRklC0yUzes89S+06LXMH3xLy
U/6b/ezGKpGmQdxL90f5+p0Er9SFJI24YFBj5KAphByfnbahB/TTATY4kitduU/z
rXCwwUbplIZShhoXStraO6lqDZsPjRo+Nr9gNQGIJAGzoyUoZ8Xk87vYQ5eEaYVP
11abn8MqIcv2zyXp67vXRFxD7B90JA57IgMJBOV1cnJeq4GvVAPCVz7M1eWbHXxi
U+Sdw8XAMCqHA73P9V6oP8S4pPg7eX7qWM9AX7huvo996ZkVxIwVpTWi3fnLqqVf
AZFnjd0fJ4HppP/b55Bguud7HIeXH349kT1uaYeq67IjILdHdrPcoqR/BhruFa/7
3PevGnrFx1FNvtNh0NQKxbmFTMLL8y0pw+E1EMKYmHovGdqYytD5pal1EkxOuQfX
zGO8hbM+pD5NFPXXXLRDSw+gp9L9PoPKFzikl7vIR8XXlAfUSM4utaQEsOErtfz/
K/JkEJwxyAuHd8oA+BXcrD8m2qnZcvfAfex+KKq0BK/uk2tqLVKris813rTkJ/rN
WRdA5+HNEkmBr7BVf5+DtD22nhaw9rXpWpYKUlEhGIbJdzvFRrwuFm4x0iSyzcN8
iZpmlhcmQiwzxeXMrxv4eiXdKugmGblGydjOAJ0hzpSoBor6IjU+NYSwnSSB8FkR
MvriQKlNL1394ux7EZ9ndh+WQcGkQHZ5yObama/P8eh1NRNwiR2V1TD/B5g2gRNV
mklC7heJZ168jf3GG/0eevvQxxid19ZC3vA/zCvcVTKVGXthvS2zBflJmrFSwgfG
kpqUxBOvjANX2qr0E2g+cAoOzDKS2zu4oBzWqdBhsdIJd3TLEWBCv1J4iL1rqKTJ
bCeWhfbqF2zJkK374aRpbAWT/f+BmOlTam5BE5Y97BzlnBRim+MgTJjmrM4urpA4
SmGjtnc1+vxjC6+/iwpGTV3JoIZulwGIx0+o/NfsHdTuOBb/yDoCKmshOVt+4tTl
Vv9TYvXlrxgtwbWZ889R6OKxwtVZMHCNcEkjN5rLvegCJKIWqwGxLFQscIz3Fd9W
DVxACtVpfrvE3hrh4MMNP5ZXbM0udqLGhAUVD3iVTS1ex8rMHmAE7cE23lvT1bAt
PCqccfTQX8tpu6iFb5unLuWplptovHbZuJQsooVEkLkWge6/JpUlcB9XQMXKMsMg
2dOJ0UyNN9LYEG9L/a3aF8TUNRmAwYt9VDHC13+5hJL+8gpbR4NVaZEoZOWEWH0r
WiU2WwLS61qBgp+tflUtC2wYOwu2nfH8j/y+PXy5TOrrjiIB/JmJqARJvxILRgxg
RFuqsezVzCEzI7068/y2Ema3CQeAplzzXCtCZcN6Urjx/V3sDUqYKALK7RJOWmPB
GMMsQ85bl7pTk/mXiN2og+tApLcey9JSD4piEu6ahZ/bSZ1zT8TZW8o0qzBIGzuw
eqWzN6BdVSLWS/8uLdoa8EWqmgOktTgsnpcicVMQlQi9aihYt2aVDHTyJXJcKe+m
15mAO9r6vI+Mx20Z/muCY8V3aALgmqKZB8NxBKq8zKdRdOZwn7s70ud9jENxbbUn
isrDIbacCXhyHcmkJe2fgPveBdDsp2lYK2YQ1yxDofsjeh7lPYarNDefzuzZHZ86
za4rxLT3cAf2z/lBW2K0xlYfr2ihV5pLML9Cv6x/bd3Hc7OBMnfsVp/GV8EYu+Zg
5neWg36kMqnnqiMiSkq7LqjLsoqj0cdb7HAEosGpW6XXHbl7K0vmYz9DZ4onNqvf
/HlEp8iWhiZK0Lyc+BABS8frXn0vDfwVfNxD7lnfvEqOr/zy2Pyx6l/Pqkg0SFxR
oKc20rH19dy8ml39lnaxQVx0UW8X/LA3jxr/dfvDx8zAQLEjrEfOJa7XmiOx5rV5
1xM5m3onb2fy0Qt40XugMxzSTV3lyrQX5FXmLMi2pNztZ/ISU50A8j8kebUCDYBA
tU2li5szBcX7s0rx+V0B85UwuRJkN2DBnTCLes6m4rVZZpHEpfyy/8GUXaeG/+r3
2uHfVf6HFDItnFWyFDDYXEseIhaNXv2XEmdiREJLDRqo170t5BwSdgIhBesEns+R
eXm3rozbxNdAl4PfofbIRkPwkjvQ+zXPmb6Gz2Fr8XPIzHY3G57YTO6SkHeX7Qjo
OSguEQVLxFfffaGEAyZGf29HbhAO6n1LRoxPQ5Y0uHlagkIjmBqtTUzP2NZ2zFuX
JCBJHX4/GZt7tWUUm0VVfvDOjAdlAS/T+QR90FvKJ0tfklnwWiHHNV2TTIwL+r5k
+YT/cnhjIxfLQG6tJUHPx771oKvX2F+4UNFyTPiMsmgrr12sDUVC1rrMUmtgFqMM
CND/AN4qfNEHoBcsBSc5WABBQAGCelmZ6yJ7DlCweSaNPqaZxqF1xgd6AB5BYSA+
8z2lyieq7f5JLTZDQEwLniZFuKEYA7tsPlbINK5S61ULM4JPejeVG5IkGJQ5RX6G
3mQvAfi+/79aGzm0+ERffw==
`protect END_PROTECTED
