`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cvfOOs9RT4mHgqbKHIJjawHBlTlnJu8AmTlfPxZQ8A3GuImA3s3R0Wwbr4TN9nEX
jBtDKZ0WxN9B/N1C7PE9tUJvj/zlfdD3GZyp7BOcGrO+SSuA5yozRmYhBhwMJLKW
jK5akXZUtlIjjBT47PcEogEHW/EQ0P8tAo4jVVCovWHWMJPn10DQssxvWgG8RlOj
5EpNJ98uP9kExd4yLBn8m6WyKBw6mxO6myGxR6IYq/u9vaZee86EtQz4BrnCBNmk
Z1THf2hsuTMAwr7yUPAJsyc+TC68HOH7oeSAdyUBbgG/H/bHDDi/6PxFSWjv+AZo
JNu5NkMRSIxkLOB9VWEo4eUDZOSA3HaQJSM8fCnR4gDzATHuOc+s3sLwLcXTnR3u
b+WtQshDLA56B8010u/P1WT8QowCFhC+fUXpgvUlRTZYdZHLtW0NoiNJw1OTy/hN
TdY8z27lQJfw0NFZWXJL78v1/HSbMRZGBxrTUsqkhh9S9xEhrLWDPxL22P7pk0gE
lHSXl3qVOK/ZybNDomR++aC36eRXSQ9pGO7Tpcc34A73J3DXB7S9h/r984Z2xZl5
hjfHjfIcVUdqsmWGi7batchviF3+Sl1jCc3VUYmdfyfYBu20X1w/oHoyQ19EkVFP
B+vPRZ9UJRDfy41dOzmoP0w8UoMWI7t85fGvEhUPmYsCxcb/xGdlJenpIyvrm4+P
E+58+6pogqAIjhPVjaRMkB6ROLBNesBZCshyMevlOLkCCNcdNoRNr90ECj6H9iGJ
kCVug6G/Zu8ZPwwuf5Ct8Q==
`protect END_PROTECTED
