`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rVv+gjPcwM7ZRz0kNjN4XK8ii1mrdpRtzfg62zXsgcNxvXq470zeB8XYK62TPR/w
uhqRsg4f4D3p3iQh2Zo/kYFMsBo7PwUcsZhh7Jffwi2T0BYUNuRJ4tAlBUxSbIay
nw3QVwGr3dbYIp5dsyjCDF2/bhDQLIPXz50YezshTQuB2JGNLyyoiLTJU4fOX8jj
/ZFmktmJBFtsyQ0+C3YZHmWgEUBwCYS7/6MHd7W+SFRciRoad87Y1/yW8KzBw0wc
dVsHh1Vs/kW+YPxAtWr1zX2T3LyrzWQ2Sb7ayPGZgCe0raMbF11ttb2XzQQjRCXV
v4XzPQTLccD4StFbeQBgwwBRLe/vYE/xzJTgShNOWR5euumkIVx9gJirAfCDTrTE
5VW1DjSNjpGA6fS9BrG/DgJ5j3vSqaFJtOr335uGf5M9mm69oU+IhaXeMSJLqeNY
FqxiFmmfJ3J2n/fjcTdwLWSl7zsGV1uIQvtKeK1WWDNlooUpXNPnWDD5sjQG23TT
asf7J/aipAazjltw0m6ttjA3yxvkWmYh6HKIvsisv7E=
`protect END_PROTECTED
