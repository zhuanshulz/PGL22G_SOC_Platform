`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BjaJHCRr7/ZX9YchXB3Q8sPxm52+EqoJiH0q0xT3BDHRAzwkI1ec1pD3higLmL1n
rW3nWBRa0WXLBjcaaoXwbFoLaX9VeG2Dhca9KihxMtg/OTXM+3dAVYHOVf92hL7j
bzdBzda5+qxAw/3KVpJjUY8xffb+ETpHCjkFNzKBh2RFDrYkEyRp9Jq3rG0k2zOB
0ObAJlgrajg2sAh8+yA3Nzszf/k7IZxlmi9swhM1Aw8HL860PZzCKHALXl3N1uVO
2u/eCYUs2J4OGSa5rqEqSPdDwqsXSXHSiWj4e/74ro1S3i76/UXJPryqOVrI+rkJ
S1iiDN/3upsGz5PrOtSTmsdQy/OQH02GVkOgXlLmhhYNIKLz/IiH/uQYuhEUw1WX
`protect END_PROTECTED
