`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vGvfhJdNb+e1ZLkDji086S1Cks1QfRqrXPvo9QI8IwTNBb5CHZPzh0ZgwSXDBc5G
qNzDwh/H26vPcR39wxvPzJ7cyGtJmzrphAio1bkA029fNw3H1KzpXX5eOFeyRZmI
ff1496Tgexvk7/S2JUdNIV5eKNE3c6iYgSMwBy7IhtOo3BgmHAsroQYC/LE3O2Cs
qKmHnQh7LLxE8P/N0ZT7iCW2HCBme/ndFGhfQKvUhKTHv3hI4zwfztRJBskIRRl1
91f/0F7PeRZhk2NvJp+XS6iCqI4n7JAcOL+2YJkN3JzREEi8JCv8FWgUZT+08RZn
W3qzDlsniOm19p2rHOvoyplfvP34jJvHhFieX0XLqIRE1yR1mg4lB2bAqpzpExiA
m/zliA/jaHd5Y2ePMnUKS/my6F21+40doMKvkTf6nPGXBlB13s0LdKLIIklTxXh4
q2x8l4g7M1FGGsyAWNKhp6hHOTN7O4qn7mGH9WkWSn3DTbLR69msihFqPVZiOF1h
L1U9MLDY4PpNRci9/7aDZ4GmbrioIlQhdHyHRq8RYKTF97nVYPjFEcOVj/YxqWhN
nO5z6/h6DQMHb0fbLtw0z0JWVxBw8a6NowP+Fu8U1TMy6VoF0ghCH5CqScMjwotz
OuNEZNocT+bCdAfpm8+i2PPrswQFIH8Ez76lFMo+QNaT4vcYNexEjoMqY4YWsNZa
OzZTOWk2UyyQEp53XEiCzEwmMVdBVc7EgkPgVFdq4wBGro+328BBK4J01vYq0q1O
YSaCsWyn3hQ+y8/pFTc14g==
`protect END_PROTECTED
