`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GH0MUOM35fozuyZehtOgF0ejYU9eZJ6YjwTGZWA0CHQ4bL6iEWeLfWThg941OIUh
a+bw9IrNa5ry0hpu1tNXJRLiD2oaIAYSMHZWCPdxix2eQFhINrEvuXlDjYhlsslX
MGZgmzlRe3/Mx34afKBhCuWaq1S3/yVliNEWnsynzoM2mGGby9vu7OVM5u6jKG8J
PlPyUTc2ufi7gZpRbJk0BDAgaFf+gxHW+nF2rMnhP0jfDCWZMu6r0/+gZybks/rb
+bYoSyA/ZZIrIhV2JGMrOqU62AOwI2pmpGHFufDWDyc=
`protect END_PROTECTED
