`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+32MTywm7Mg+tj5zxHWlmMrfH88bbw8OGCyzXbST4bCrx3rq25mVUeF8FmD2r9j5
hbnRFMoxR910tB8sqTuITI04jeITo2fXqoEiQmCYX/YIg6jz+fqJIS5G8sqpFN+/
WZSuF5Kip7Tw0h5jyuZjvEPdG9wO+U3ZSJBB0J6mepiR8WV7wBV82NltbMyDsSU2
nP0sonWqZkwZmpk4TtG1pUPtakXQ/Dx3rNHNEeVc7Egm+dvHDsi8vEbe17ioELWf
SNJhyZsqcebjIZcy8NJEFUY2oqAFBwaT7xrtuMgsNbQM/ow5YORqpI+Pdntdb44o
gomLd8nQkSy7JfeuHvnKbi1kIpV//dZ6oG3fmWg0i2BcMlIgcOP9Y+P9BZYs7i/x
e87B0gxJlUC92k+m1cHsoKY7gotU6oA+g8QGuHobTE3TEeXrohdaTaODjzhPkW/H
RdNrn8/Sq3MzbyBOyTgyGIsBHfFPP9j1xiOQ5Co9kIN+stqIGshI3EBYAR1r1laJ
k/MRY1iCVoUebxKvWPMiPcD0xE0gm1vG1JkbKnL27qz1013wZY71qp4a7aJJTq/v
uF4F5ud9Lj/AAq8x/fDK+JmlEdCx5yqa4AX3a/N6uMUAE5qPKtHXf5nRIJZ4c+Tx
XilAHTonau2jVB7VhEEI/YIUy9bgXr+cwEw7w2w6Y87G1gIv6tCLrtYMHq434GVj
zfdGi0XRuUJvtIyz+YN3NGeDiOH4/e7Pz6FFAibnZJiSQKSMiyuA4Fpxtc5ewNnv
SkHme6lKJMWrCPihno60tIwxBKQbKAXLTSKa6Ws0D+x6uhtLmjHr0bICbAX0a+12
A2Nq8QwziY4ifKE2LiecjWK2ahjQmIYsISqS5m8NjKsEPC/eE/CKptGc+B77eU8w
xD4vzkvk2HhRbC+iD1+RVG91IbWn5aDxaolhx+HNNWxNeU+nEa1dUMB5LVE1aJRx
z20BGhwuyyO41FPyX7lJMY5isHZeUwpJ4+778mP8e0MZuNWkubKU8NnmzEj7jTQJ
xjcZZJKo9MwyTfa4lpFtdJVayomOxx/Yo8/s6i/cKUi5L92xcDNFHS19hvZQE/g9
j3d0h1gRuGgmnXdfuyNmCanwSzHXgm5p9/CBYMeeXhLBRDDKQM65MjHsqidN9L0Q
SZDkXLAWe1q68i37vM6ChjeHCp0VytX7/uxxWXYGp3JNuHbJi/eKFcUuU9SlxCuQ
l99UoWelVn2Izj9aMuddViHDFHkp5RsTVYdGDJGutfNktQH+icH1y01EBC/UK7UR
RUgpIVekg/lHXwJBD9Hwqh7BXf7OQ+rKnt6zRT8oRd/Vmg6Mz2F/kgXPToq1Vcs3
xhMhSPXbwDEmrtq6Aw/nMEGUvJoL551PkwVdd/2HgfYoJ+Tts3vEtMaHh8Y+lvkB
r6wEEc1no4oXRhwFyFl7XcsPf7ORd6/McLgx/aEESFvtWsHwFXZsD7SS8eqjQY8H
pyr0+4eNQ7bHnElD28BkN0cza+PkbeTnq/dmfOf1wUMl7jAy5BGUGsC2bGShYQKO
zP3riNzmLUp2uFJqWBcVKDuUQ8krUCx76vHjfapIKHv4Y5UzDXgZszm0f6uZguqY
iBG5bpfhznLAAnGKbfLrv65ay8RDyauun6s9EiwLXz6pKqTzJdL7NRDNUS5s++RC
V+P0TgSZuUK3aaCJFuJm/3QKeVJBxK7HK3t9txYdUOnX2S59NNQXsT6TkJdxQp4W
Y488zfQqRXGej0jkdZhZY/Fq0r7HQXCNWxMs1WOYnhA7Lou2K3ieiowJHbVAZO0/
Ybbx6uMMSrS6zH9JTnoX1LGUuD3rmBcrwjZM4xJHZ66xn/nueaVkOFF4Ut4HPq4M
W44EXT2uJyNTccPwO96RMB4e0sGAF7+TIHtrfhClAHXs02RbFaiETJNlHV0r51aM
zrqSZ9Gp/ZW6H9b7fZI5Fg==
`protect END_PROTECTED
