`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2CYjNWdEWTWGPpILPFVjZsQQiKtbxPfQtxB6sbYfa60RaWxL7ou0crVZeLg3xtGe
vlBoEotjOvXUXs35eZGzX9gGJEhroOzj2bdveM/OlTId8j5in2m8zCmWpOn4ho9n
cyWh8xxp2GjAtfTSKv1H4lOCWjoGjG9d9g0OGd67d2UnyfTYIC9NhVf7wWrtFYH3
DFES8tQW7PA7O/g3h+YX2cxbav/Bp66mXBoaTFzG7eqWHeeE0Hyt9yB0+XD/CPWB
0k6uyvSmQnkn7DyE/exAmczxMqkPbCXqZeSIYpZXwPTinOn2LQRpWP3nWR6OA88n
EeZTPOnaLPlpShAsvL0Tpr8jFcv1YC74FkPObVrmmx3arHv7UyIHQvAugshuVdlQ
7LkJxqHiB2jyreOKkRoaqFmfL6c1fgne2KcRJS7HqPjlZxbMuUMzLHbrAnwLq8ml
7QyWkqAJhGziDqN1/8KbNG+hm0YgVux4F+e2DCMH8HQ13lRcD3KP/tOMePvv68Uu
HV8yNTJEXBpgdabr35tSHSDXZPiI1Zhn1NXANc+lfnHT/vPNwa+2Ssn1I4PgbG8m
GFZayKOaK12I5If2Ni6XuuB8jQiycPCbpJa2xmBPxYdFW/FrRJigV3telKY3Neok
43o6kBy/USflIa9IcaYog5VWQ6cOV5TCvrjlnpPyEksDtdlxtkqUVjdWRnmznTOq
ctvUDDF/pFz/SDDeF2mpop2sVZHwk8gFN6xiL5zyzOz+MVqA2Ft7XP2s17KA/n8s
9dgRg9IN1WO6jjcw69k0UbnVBiH8rjnjJx0J0aiDUiCj6zyfRnRLTJFQee+2gAII
5EhUei4OeLjBPgIUg01X9F8hUPpiw7EImoHB2eE1rTUqGu1ZzNEt5nIN/x7IwgK5
tVQlch7ieaJ6A/ZP7eqMApK7nWJKTTHxJMNx5RY0CLwTr6iKllRCdgGhVX0uYxKY
CogJ3/8PX+hcSIzUZukqomMwymbA3NNJrgSU81JmkSdWfVV56sBAqxBtX+DlcmSH
BDMd4TpOn/hk12WzFCUulDtpGwtLOt/0rvc/cjtKKf1YFRMxc3mJy05CsvtH7tBW
kcHzizkrXkkQwoomBv3GdURkEQrbVsXZZfBwEdmtbmrb7YFiTF0NOPjBYwN5qHMc
Toq476ZHN3Sxfxb3jSa8akhjrzA/TSgfv3DJOBGrNdiViq1Uyr4BtH+t6tOw7DJo
mmULyHLSHghAKnbjTE67tzGtH0Oi3z2LPgM9T3NBEeaooOw4J2AF44k4CMaExYq1
RyIIQcsEohK9kRMXirHaP8x8mV4bn5Wgb9ByguyNwm2NpX8NaeMwf0vuUd47C6Xd
A3nLZiOJUkeBJSZu32MSV//FUSLfm9VtXko8aDCL0FTqh7S6qz8BUY7eu4p2+mtg
Ho55mR1FARLlJxZZ5ulRZa917xv4XyUBIR72Kb1LD93wnnL3rzyIzsEvH8RzgKVA
PZLYNyYhKgTTXrZmX8PP08KwfTGoWXq9mWDFilH+zzWDDsHyouOF8IiN73j9iwhm
QyQd5qEalBDa7DbtSUP1EiXeK9ZVPJhyzzw6iJpi4czPGjeeO2ESbBXpApYcpGK2
aPdpBnfZMYZLfSnNqjm4SdgjzwCbpbkBMFR+WDEiupOCaP4p4IYgnvlFKDzczgfz
LJplkI5sCFGmUTQWi2iO7k5Wkel+HuKiyceYEwzVVBMggMzXmZMons+p4eAoWN14
CTjD3mNpNbWZg8jj8vNS866ydLFK3tqd/PspNN2mZsRrimY9LJqzuhFWV8K3mfmu
LOgfMK5r4BLINrR6qVQVIq3KNYAWnvz9/BdL71ET3uqm9NURcrgl9/lpix+/8XIw
EvT4XIQjTBAO1bsO7ycHKU0wGHg1B6aGrOdW1b7Q9sULgFr1iSOHSGh0c6skKuUs
XU9xcYPsQb0C3FcKryEtyV4y4+5O9HNztGqlZt2J0NpQONtXwkBUGo4h9AYClWwj
4Ci3bgb9t4sa8wfSPnpINLAryimyyY2A2NiZ5/sP7Laj4P1IYKO+om9URZhffbjO
u0ynneJHq9vFkvN0ZWrxtQ+vB7CDh4Uokvn3uxBz9Hkwi5EPsz53x1zWm7cJYVXt
zp8RAJxx/wpeiyjGPPX8ySsBMwX7caywEWvyVZvPQWWx0Y/A5MrszVMgIvEZV8bt
7fwidCHJzGqZ79eQVG2RxkvtLqRqVO31lDucbh+b0Hqd6SbgoBZlJbeF/aO6jVd3
GtGz9H4CLYtbJv1dyVDWo0C1+Dj7gu+uLEyEAy63yvKoFCrJh6SZvx0tbeibYvFd
YhtjwDTdNXYdMCAGkavbC5Jm4ipAeaxCScVGzHTLQuo0qzD/ysD5sW0rV74OlAhw
HQ0M7ImCzfxpLSRFOpmmfdOKHGMaY5ja4ZSIq2CqT3FREwRN5IHx3Q5IFOZs689U
uRH6dQEiuuQkPOQnsXiZdIt00DoriDF4gxrCQ6TAvyJLGnUUBO2NMBa3gJvQPeV+
ncc5mCXUfpMASqcicaVelItXO79d2btzQkEiVjI2gyaEftX7LXJWbdxkC/s+lmaC
jvFBCVzCdQTXxfM/3qCQ4MnmxhEIojzBmgC+IT5JqBx3dpQid0cs0u4wGzR4A4iF
Z4mMHjdQUEXC14D5C4fav0mGOToP/sx2UH7zP8uQScVKDCWGWAcieXCrpon7w3Ax
PVun+ayUHJcHpW6hNY96t7dbKfmUfqvNbNEYglJdSMrsPacqTOoTlfNqRopv29Jp
FGf3DzAuwu42XZ1sfV5meWplBeEIRbQKcpcF2jsttd6ikFeMTH69Y/51kRxhsZRg
Fncat0Y0eiuRqZ5ocd+IFRdVufj6OjLMmq/FX3xsSSGoWRkWq4KGXPFZLJLicC4q
p9KkJPo3EoM8/UBLorWR0y5wR1cxFwd990KSiwLUWh3J+BR/cEsJgeHBXCrMJeBs
g0TEjO8VO4cwIKeTqbdOvWPehBW163xSAYhSjPR8gq1pakC4oRW71gsK3v+uMAy4
3E8IBNo+FNLx47HFiZSoHfpSnAK5/YruhuRN2LM9YeFifFZHM6A61viFEYTswVHS
EanEwv2Z4N+YT7UEOO3CqBjaq0E/Y7/1SXC8eFobj/NUU9el+fTUmWPbcf9vcDMG
Vblf5hB3U5pHxEIbCMqgb8SznLJ16QabsseBETNZhE4VEUBMc6n2AWkwqJE2schj
lt+a4V1UFG/HahWB5e1v9bYDICe8JkL2HlSP8p/HCU0XUex/b5vEpFqkVdd0/lsG
7Gd1+ZB/Dgj+LejVjggINeFqcUb+iXaJz/lFmR/b0J4Uf4/f2nTgP/8/kA3mJwTA
qdnQmmp1rWflnShUiBxB2ykU67TT5MSrb1APSHCa1eg/ls2jEfyE/DIhH9B0Q6f/
WeuRfbPrKU7D9G41hYV1m4b3ObomfVl2GguJl0eeeDzkijLnRVpVlWXsDFMEeftI
jVMJ4/yAAWG14NHndIlAO+VFVh1DHsHZOIZY2m9mr/7ZJg4MM5b3HjrsASKvD+oZ
9IVjptr2ma+cVYZZ+kw9ss26ifffDTZDpU+cxVDbV/1PAAupir4WgTVZw4zaGFXA
x3tUhXb5hBjN8IYEwS9ra2RCadI2j80jKG/oAldMr1mw3BzuKYzfdWupubS8cDaZ
jQyuiWtNFXW9ULpRzR+mVTIfWRi5UykgYRM5oh1Zx1PJGLmkfMrtpwTq9mgzTtZr
4GuKXUNH5dJZKTnUWF2Y7ggGjVPlVqL7E39znlXjlstAarKsj4wNb3JHTtZ6hwPK
dXJAqFeMQHMHu+4b39im3VFQBC7oxAlw2wDpIlx1ZCtOREveSwsIHHtwGWZTd5oy
wkNSj9BojtDZmlqgoXLo4ncEgFG8W5zbqIzEPoON0kycnm4rPP0oNIEhIvscH6ZP
TYf/yOmNFHMjKnSRSaZozjC0uWERy+qRUuu3fNYXA4YnklBXn+0ABeXjLFmnMzgK
IeJQX2TnlYmhmH9uCsgRKxYCecbsEj2fWH0AcIKOzXDlTJ4YPtIs1lKrqufDzIcE
lRNCRo8AlGdmeyqWlYDg1OaYfx97jg8d97Cq93KdpTbj8zCqQqiRwUVT+SQMZdp6
W3hNkMgX+8Js7HbT3W3OsvEOlNkjTQ41paJNNBRyAiSi63rdMfAGrk8UZ6i/jOUM
HYvvvZqFRikpZ35L6rTAl8T/EUfK4rUoJ6nSpTrOgK/dOi/XyFoCVcOEzY6CNFYp
nZBxHHBqzRMVDpCGP7Pj8KH+pTKIoIMmG8qJ3SMOUFALXwd6PzKFe6q4DIyR29V+
VU4ljUvxM1tapbjhgFVjgHarOO3a7EAOQpVVZAEktMOPBz3hLxzuwoNVc4np/RJQ
SLhFFhDt2pqBY7N2z/cHDmPmXab8xmBrUB/ihPaTL77N6jYhZtoeo7rIp+38wMUe
ciNAZZg01kSMsNgoaGYJ4yN9x48PS+lxM0zj+I/+hiEzSF4cTw5Jatl9XhmMcbbc
Grb/2faaUHhYAim4+LkXpAimIia8rcuNDO07BSge69G8Z/d1PXCSIvHYjEP4VhPB
RfExFQbQsJCdX5IxZpMJ2/c8GjAoNscn4tlcKNBl4GQ5HLzNNH6o3eMb5V9xz1px
dPG3iPjbrkmVX3iB/QjrZBZGLGrw7DmF5CH7vWmSkvZ7l5EZ2pnTX7NnWhtz3noF
QMTowBu5O8pksDBxbPHAuRd4r1pMiAfAXsICResTZgIabUiiKy8FSCJEQVzaKIn3
p0M1MJQOd7VD3Ce/0tmRVZc/if36KRo3CIv9tfCE9rZlLhR7FYHwdHU10GSOUohA
lNHpo4CG6HunA6C7sof+mjM1EsUrdvIX1P2sxbDRMP8KK6KccBQU5hLjCWOxPMwT
IYnR5VGTZ+Nl6xtKLPlWjmz6A1zy5o02l+65vuAaKdrN0zaBVOTGxaLeCd/XvT6S
lnZD0ZqraAiePeJYKZW5wbfO2mdvwCfvNB9tgAynbuxa/UK5eAyAsiUoDEpUj8/E
FRl+Up9E9v2IG5S/cJZA7fHJePOOhh2PubqzKnH1hWhQAasA0+n3G0PNcfhI0uNx
RrziASSZcMiI6/EipFshi7bSHQen7/fUC3t7ydWmj6EX6VNNj6KD0tEEkPIg/Nrl
JNaSNcydzK37dF1rIDBM87+QW/fejTh9jf8qd3KvECkD55ThfdrORYd5fY5DRP1P
Ola4qndkb30e6piO8pT19UzQECy7PQZzOxnC9y8VPUw3G87BrhmCEi4o1Hv1mRqu
5+iHYIkHIAAy7Xn3D8O05Sn0ahM+Di23g/O0BuNAano9AQ3RfNvb/2EysP7Lbku8
/wpAw+QhyuVGUQfjN0NyEL7FdQ2dcBrrYpUqFk8jRLdiH+Zs4mqj64XaA3gwKiYg
vIUribOm/TaXNy7nOIMYDIamm+5AfbfZkAGoRMw/3opIquWCitGw7+F5gyklN4Y8
ajvj+BoU/2wbSHSO4MaVv+1CR7HGcNINzKO2ZGKqXijCsbolHunz40ZGn2Dlu7Qw
AN+Xk28riOOMtBGajnCjQ8Q4zLSxsb20d+DNP8cf67EXZjOmGV3nMlWdVpkW3Fzs
N4Kj3Qz4luMiDf/WOYhi5IOwE41/C4ajZy2y/IAYSo4jcDGKZaYoKequl1cyP9um
zgTBLwKPf7cVoO7tiB6ZkjzTQz9hK+/7c7Gspre2REGjWEHabDMuvp2jECZFjFfC
JftTR0KL1ijdzDCSfFskpHgqpDEQtUuGZFFGGl5rEMNkFKmm0dEDQXH0nyS+VTpk
Q5+Vs8TvV6vNAeME/KTXwYl1poyPVN8baLEdRKrWfU5ies05VI2QxLPgPYSvO9tC
vgOJ93sQw/b07bbiLzeIOruQe8+WA3POTjy9ZnQNTDRV/acxGSa1+e6YOPrQ1HCU
SMjK1nnNXemDA+jjKSS2pDbuASa70soIbtGk2IrXhK1I6qujhKthLLm+BCKOunE4
pdKqAlIXOSgNZ3FgYa7bm6qIgMOuNCa/fvnM9FOb+fty0sxODIEvZQm7RzV8o0Zx
+KZobVZv8yS5/Ty4ffB9fBN8VoTnGI/7mIPJRSxn/A7asj+jJQoNCkcYDIli8p8l
wPyjMfpdt4t8/vws34UuVvBEYBuDO/Nt/TNFLzVa8i5IFEhMGuR0Q756Cycr5u1l
2I2R4uJ31fE08aIwiCbKT+rJAOY65wtacRrSqU7TgN8FWIVcSIh7ghSCm1AVzEr2
/ohnA7wzO3RcF3T5tycmlS56j7S0YLDrPAeCP9mjB7jcpwOo+8XhnogdlIVl87pQ
RBr8aNxqYYtKKeb08T2L+yTBRVfAXZ9zGdjLHPiR+19kWk8izOUEa+TAguHHfWws
aa5zAxDagVanjiaio3ixVl2rks2D8hWUKPPhyMD8eYEc6KITQ0rtTanafJtaNygR
pu4qbcEaD/unxuPKZsJ22SRGpReIWfV4exUYrWDeGdWSescVp6zjrZBmyd0oG1F0
cRE9g0/3nQCADk5BigYw0w8V95o7EouMEw3Al48HQ4OQngD6xLB4RMQik28wyUiE
6kh9pyfGbM8khpnKQ4FYLCCKv4TzE2uwWoEJaFeUzDcKbQ1nUMbeQNlLffNtd1P0
e5X7bW3UwHsJJB0xlcf8sEWzxHz2YANWzsQHOBnwxiQmduqEREQiFVZt+U/NbO+n
aWYoNvNQcSiPd0hXYIE9vvhm+Yanq9eBxeFWa/to3YBql6VeMTkZDkZHIGPk5FO7
4oheRRoKI45av4YRVhXSm1LbmOYWCI0rSNV7QuDFGO9zpJgtJ/5og6iYo9IGm6OA
veO/xwd9A1GOlOpot+VlvWROW15echr9sP+gwNIYLF2bixDpxiaY1ZH7Zq0fzXVo
ZNnwQZqsrl5Y4B1w23S0nw08Jbb/tmbDcuUBE6It/cE/CPxguG1MCcHP71eGDEdw
KDgJZrrlaD/0wxhn3BhNzwz2nKGkgsA6Ay0J4F9nypdAix/b4Da1/8qtrkERGHpl
VYIiEApkLDYeLZGXuDtCTHvQGYCe5gB6SvyF1fhP/F1P8ObJON0cE0ton1gbxejo
byIi1+QBBWBmxEKpClxdji6XqwUMHkNbkhXT2GXhVEgIBCuY9mWz3HA3RST2GeI3
1sZ/2b7zw459BR+hQx9d0GkV3c8ojSex1+sSZOFZsqe7wvI516zq/JXSuFVeGull
IQllos3++55vHN4QzdligFivSjWmItpA4pxFCtNej0rThC1lAoz1cBoiRzg9VNmk
YnOD1TZ1VkQMh4KiTFZNgEoNniywPkPRDMVe1OM/A2Zv1sosGipfzXUdfz80+1Jf
ZPQkVbIMP/DOfL2H/q2/O171P3JWmzaTalMWW1EsVu+PqbmPrlgA5rXN9kRNiqEx
vpxiQIEzX2yW83HtKzD7s4E0yZFgAAaMGnmXSmVdmZ9pMRC8Neb+AQjTV6k3zVp6
E8PNMwT9XRwnoqjLnYLrCD5HL1hSvdekDRLBcjueEz6ZHfU/jQwJvUvorv7KVor3
HYkWUjZVwZObvYzSG7mzDjRByzS3jUYNJGPCziUiF2QGHK6IYVfrsEgG9fopwqgw
3gdDWr45jT13gDWpTQbF6UopbyalKWkwzT8NTpQ0l6ZZq344rY1n6uMUJtgHKqMv
MK+qsL9TO7kcQipjWME0Aj2JKQhe88nuAUilx//fccd9roN0YDXBvqBI6I+tJTRQ
+iNW6o1rC2RCJKGBvcWma3vE69Wesv/u06kU4cAVpc4tpqHs0bymkM+W9QlF9+Vq
iGPCWV5c5I1COJE6nuXemiXCLWtl7RiNmGT7m7SHpvoT1LS3k34vzGBorlELKk30
Zaps2jEVWsxgK+a66mloDT6dJlsO2Y8ywXiFcAuaEz3Lnlde4sevT0cDggWjyVSn
qm1ENjqVKX6U8ul0A/F9yKXVhpruux9uoVbij4PcbXOxQMZp8/vdql/tcMLsaYVI
D0C4kT1N+lfH0mBaVLsYqSgVPK3PbBB2eC8nDk9DHt7IFj7QstjL52vxZqOTx+pz
/gGIj0TkBd/pMIqedT5+S+20sI1+XnQToHtavVn4SuDo14lDOc8Od4TkxNNft2Sx
mUSMWMeQeKoIJCt8k4VmB5v1br09HYFUu62laXmtbhmnoRg+TnyB58MQpE8mA4Jx
D5X6S8eAzPXtSO7GvtmehcUe3FfxafppfKjrjWnMd1tGtqLgZI9Ldg/FbEJijVFC
JNsdImdmBIeRFlNPbJSKbNPFrODbhciaVyATOAOHxv9sECCrGpwyEJJJcYHNcpM9
VvsYW9OgH5yfdBmlgzvcPLk1WmcJhobRFmdb1Z10uwL4BbOnZCS1QgNwrAVE9KGF
LQsBJ0LusUiFYGYHUrtp+QA4RN2kt9z7hKhG0atA/gsYrHzLWa2+/aLZ67PqnbOZ
/lIrEhUbyLBK8dM6KivC7rGic6X1iPPigfIooU00sGUBppEDjOLuT6zdjZHfYJB8
FklBHPuC14mJZTaTxS3vBJb/FvhwG2WqsuQdbl+ARm5IbPD++BgHAlPYw9LvAsMl
hMxwR4Ah/U//5FHJNjetSHUCin52PPRGeRuhCdeVinrKgqznlT1dT89MaAHrZhW3
cWtiLIR2WcRNTVVcOZ5EiDr97LREmp6tPE7n2bTKUXmf2O874XppBkgctPYtbY/e
XXfs8slXfi0bSrGqYGJop/lmCykiOEQ0L/IZqvnC58i93PMz+XGQW0hJMIfQ8pUL
wZcJheF7cBNkIBkQoZnjZLKSD6vG8vfC2muiMQBfNk3o0EkqnEP9fbQz3zvzfAU8
EhOeZeDUuPk9Qq1tj2yD4x7/pffLHSY5OoslmezWeNrG9IURKFtilfxbaRbqJvfn
jQM3GIccENVNXFSnxPtUUqcGJZ7tFRR8qwhiskJnzAppssOcQvPU5OAMqDy5d2E8
hW7JcA9eBIhm0iCEADoDVj72QsAl3eN+AOIncM1AXqM8CIjo2jgxSRm6Z18OaIzv
yt8RglB/S+3w6iFFHWciDH6iJ9ns2sevukUYkiFSd2iK1214KK6xUeQRjWNGfoLQ
OrNIebzMUIv31eTqRlLzY8y0x4QbxVePfSb3ykJ7lzKwZ/yLoaqGXx+bQNTBNbLv
Vbl6gQ6bNJh+O/k6BWHPcjMCmCE0XJXPkjTdU43rzV6qIYownvOzAmxjUnbqq/Tv
+BqG7F+EzM1JlhEV/aBcpnv175MXBmvsgGlb76CytjanSxfj0Scjp4/OWHXFHZfd
DYlsP7brzxAipFBEHotHeJfz6m+Al7HVcUVIAM2lQkBUmY3yNo77ZQg4xJU2UCWv
KqTJpv47M0efqWjjwG3WIAbW6EaAjRS5LIhwGOowWZVpwnQwctIR+3Laje/df+z/
/oqHYDtuSoIF9MHsuppGINEk0wC9An5K8tO93nRLRVFWyM+EOm8nlcXyU6ZC5mV/
j63wxTNK2thX94SNQK69WFSjC9MuGzWeH9nEYyq/dnpZdhRuq8WfuXsR1XC0FtU6
4pC7Yjuo8ZsI4UQ5VF93C9K9JCAaw2sz8PGWrqGzdnJBYg6WU0mC0oU/UYugYg4S
B8ESQVCyWLQJR9ZJaOXG4dBv8hhd2i7wFivfKfY7aGhmd9ptjYQeDuz1oAhbS+9h
kjmllrQ7/ZeNuA5ac5jXauJ0SQ+KJFdLKVpeO+uUhq6D6oiIqysZCs7+D+CMqupM
Y6J1vJEt/Bcj/YrAa+vmTPSdz6pq9eqleS8YyBgREO/9wArtDghTejI0WXyIyIBr
DfhBu/9y+zrxj7fgyTSNGoxKFD+/ccVIy7uqxIvWew1S7hvAV66l10ObyHJMCRUX
v6i7fFj9l3oy+lx0tGOj8GeaWqLlkUz2/t26r2qs3vUBBoTBNvDFEkCK/XF6QNso
G69OPaCj9XBqiRqyU0l3xfo8N995YRzqp7PXM4QdyciVpvXIOFWXJPFt1sZ9bimz
zAEbVdWsA57jIxRbmkrKxthG3UWuhAk6TjiI4Z6/0t+64YEWNv+Rhh450U2HG6Pk
CjdUpdL0JtVu52mi+DjI8rHElTvbRGNPHK+aw7rwTBv/8dbrkreyNwsD/b6W1Bc6
6iwVkiOk7V/8CN+Pm0LLTlf7Jx3S/px6wXtIDwt9rxc96WwFLaxve0Tth0W1KTpt
O5c3gaHIvzoF5Ww5V+lt9CfXENuaRg81/oOe3VBqLyRTBhjWB3KO35vETXKdHMGQ
Cjwcl52mLSkrXRlwmpeSNXvSruGfY4rRNgezf4LPvsvfdKGBOW3Uburdy6cnEHU7
XzcZ7OunoK2M8BpJgEg9VDC+wg1kknp/xamZzMehhA9pj5+f6372oC5L7o8aj8hJ
vzL0hFh2hyO/WQx3qtu+xGjNWHkQIBy5BIKaXfdYuTjyfy5wv/qTu1tVqUmQKbd5
sYr7sKL79DOn0UugvUpggnngUCzc4oQk7YVSxIxWvRH77rcQKDSiaoq4nqObPX7w
RJEg5dvIzq2RuDeQIREfRAX0UBxlyW/o35YnyqybdvC/4VT8wKhNfCzYiBRie4EV
MgPitKEVKd4B+wPcyT7RBaiRWzD7s3Q8FFqB4a/uK+DeLBrpf4ehQ1yYATPnpSD4
BuwPJkR6ERjQOXE6mvHjmsnAvsHhWxnrx9896omH6bzO6hcT78pUffgOpclubGl1
r0dhJewViZLqg23WS2U7U8djXmLmKp3NNfn8SYrfrPvGipihu36beyAoTRSFzmLr
+jgziJLvxsLN1bSXHLWlFaMstFj8NzOms0d4/i1Su2xkroIIyKXOhfTQ7QGeQGbI
Ynek6HI0W0JSYQly2xm1Rc78QNxlyOmIqJw4kmNPvknGx33z7JFyU97CpPRyUI6n
vw84avxoqkniv2A/1zT05oPYK4ZJE08UI2f1xgu7TTi2r14gffnGX0lAF4W8FZds
aXjGeTLeZiCZp9pHC1KPKj2D1GO+EZoL+NPrdDDsA1nekt/5JxfyYnHzdI9J9Rr7
OEYT/NbeuSQESb46/dTcd5RZEKuSxukGYWqYQwiIF4OkkIef4cak95V0tcCLq5uo
2DP3JMf7dBM6Wf8UXt7J7W23aW7WIOfg3MrkNvjJKpU27n10ZVvzFRuPs+d1ZTaP
GDmYHJ5e8p5xVuVbrHccMmMGyyOLCkgB2ikz4xzo/0IQgn5c0zh0n4YMWhF32ij2
q/SHWcvnDVkKL6K50+jfFqIBV4B7ojmf30kTzCwMw281tf4FEh3GNXrFUPppLl8u
kMRCWfiiiaHkJ9LkKXG2gdy7qvJUgB/WTsHJYoQuglO37cubzRklvZuhfddTRHHI
uc1SqevU3vm+6ZKkZuhD3H0nPy2WyNI/7LyUK+OtN5DPurAY+StMX2xhrg2o6O4F
dqcP4y3+9mfUQwTVRHXZS8rAh1hOR8iubCDuhIHL+au/JM+qlw93ymKRL9Q/BGoa
NHkVY6rtQnO59HnK6lIpa6rek8oQrruj9pAG1iIdLMMF88u7y6jmwAESESmZVHQK
37cxojUUwC4bKda0QrtWmJC0iP892iu7p1NOg/Jig8P/Y3mz6TwuuBdH+RMaIE8q
JFUJhGYTr4KNb+9qJuej5fwZryVh0/rb1/xMCzw+IJZ4sV+4jKUR2bU3Gvg+Eahu
fQ8GCWTtXtRjzYl1ZmU11MPuFa7pyUpSOx2NNLC+291IexZ2HuDVunzG9XOtQvKt
ZeZ0k2E2dmvp1qBaJgoK+CJ/d5gQoEn630MQ+M4lDxxckTrw1GAv9FqRp+U5wpoZ
NgPct40WPsQ5u3mHOGBzZcifz+QMYkTetuhMxJontdF687lvzbk+OQ3PnsBD9P4e
9grpCQAGJr1z/0e/ul56yWlZDV2HBcXDSGdXp52poOXWpzgMIDkdSBfAqWqxyk+0
SmuLwXmIF53IaFNQ0osHCiShU2/69JsK+J5FMw0JEEL0/Ma2ijbVyZbquqbOkGwC
S0gU/mn3iBWJNiinb5sn1YzanDavE4WlnpgS/2gLpqw6w1CcjalWshgCjlCLKnj9
OlsihhMGR5H84YJNYWGqTSh9j6/Da5/KOMHcq4TcbChA/ongdKrrfHP7AuONQOWi
WvTYcK4mTPbgcgHAcGWLiPqXmxuyDMVdcb8cbvc8G5k1MVKIHSAbM9TceSKC9Ju8
ZNZZU3nE6oGfGTkBKLhrUL2/1aX3nvj94y0xGwGEyIjPoR1NZ1899ObUGB7A5Itu
VeJDxy1iPBy7Ql5U+Xft9IsbzyiPlrDWiEyGxVAAZq967VoN9KWczhZwE+K6Kbx8
d6kEOpVTkuRn+x5O6kt9BcBst1SswEjz4WX9H91Ohige6GgVX5fW/4SfxJAy5eaj
mqh4RVOKvC0DGt7FaKelCdwZdmYEyO3dQkIzE4yQkKyQvSCoXn0I2TwzdghNyPju
5nrrSG/xeIJlZoheH7cHtCDc7WVhiJJhjZSozb+/SbSPbs2OvlsWB4WXEVKEWPhw
7sUmpFW5I2quo7FvQDiUIsr3KvXS3lmE7LDfZ0hEymjlJN6ItWdmBql7PbD8Sg5o
AnVvPLFMOPwvqIXtHAJZU4tCyQlI56KQ6/FpJZZz4PMg5DLP4rQkoqZ/qZPMGLyA
LoNFRGptNEzUQ6Fvup4/74u+msuHnyVKxk/8x4iITnijBb8MVk2b267ldE9l4Ln6
f7M0t53wpRn4uV1SPY1wdA6htp0H2mHWz3mnDtAYHCRvt/iq3LPQRhlIWgJpwOF4
mDg5K0Moz0v5XmakK62oqVZ37Ml/vHn/k1z+SRsgUcNSAj6J9F/d3ezPQCm4PFm/
n1RCMHMXQ8r0+Y5yp+E3xtsSJLO5SfzBQWhHMB+t4tVbPjx/uPcx+rB1PmA1lCS6
+R06qEIpU2+4O4Sz2OoXRmOgechDHgYat9nVPbma1KYgoBtpxuwCTd4T/QQXxc2v
9IACnX/7giSr1Hpve9cmRXf7oQTpMaKKd7XT2Sd7dUZQ+M3F/1KhVIwplOPLcC6U
DD93GOtzke0+qp4/vRsRC7eaAfsYDw2Agml1+T8wuGgjWMWW2e8FRcsCiEX+SKBT
a0Xo5iIXc3xefg165nsQDinfxK86f/veSwEE0oTjYAFJSl34C6WENGWL9IqPmB9T
1pP45FlyxT0e4KUldLaUTzE3yg4xhURUqNxSLMvsBpQgW9/boGvNB2/FN4D5c07K
6pCHNEYaJvHtHo4i/yyljI+J0Jyq9iJm+SS5eEczxDigvtgvck2X9OiSlX59EEF1
TcphRxpdDRDHBKGH2BcTtUXQx+ZRWDB+rziNSUoPIUBQYObHQ8FJyZEjFXhqEUOg
FK44EALARjQClDQbhb61IuIULdxeyKz+P7hfkOc6PMVJ7aEYw4fX9uY8D+lYmQC7
rqIRZwsv5ZkGqApe9+eJjIRMrMkXU/PLN5YbcV29+frkTnPKJxbS/vwgbxqcytMb
dDaIqhRVX24LoTa93Tb39Pc/yYhCf7xq6Kpy0u1t4VmukbxQo3IkwH+gjoFZZ4Sx
0WRGVW9kr2fwDuQkCbwjN5XIq+792QaST6sJhQut/EDdeksxj/jZyGZAW/THjFZQ
1PlAv+PWt1tNDYjrT0SXyA74yHRf4yIRG7ESMy9ZUsjuUUbxQLyLsFEAFoa51bkh
1hrIuX8ZQu+fSZyOJiRHC+cSBAubCaRMl5pFiMgnZr0Fl6QK3r9bQ40ZEbRDfgQI
OBvhgUzb+GIyplrX4VSpxn1V90X/ECjPv5DnSp+WEuQOCy4pVjAiCiXKCwvraebP
rrqaVmFWmsAGF8KXeEq39577bqnFwT+Q+dA+XolaSi2Gp5363wHW4LlO15U3om62
Y/ictSFYHAWNHeBAHJbGt6ifKCZKtgbgbcFHJHhsj7NWRBUZ6kJpk6CrQVzysiUl
QKgd0f4+OKevzPyjeLldvGG/Kb5xWI+MOuyMyX1gq5gW/d4WQ6g7n35aGSqBbiub
7FpwLCL0mP4XEGSp44Dgp1rlGilOVXHF2bChly9v+wpvNWDY+ZKPxsbkPle/MTCa
/o6oskkgmUcjmR2YzetrUCIGXUOBo3t3kyb4cOxYwd7GEx8Qp7P7VVre0R9k2vLn
j14P89lhnY3/KQlzkgq4VtKvxCjL55IraNeVUDsatWNmlqmIsXIZsN6MLiI3wl4G
gsnXkWLaW0ZGn7hFOtk0PEW3wgyR1xfumJsPkXauIbVCeH0WBYQ+B3V6eD0M5p+u
nwp91iHDjOTZ+LlVa1fm0kUc1jdAf59B0TSuqESDXxwy/f6r8+mV1/BfmPQNKlcV
TWDRhfmDGvRngJ7m2onkazPmmCbFDGJ17x4HrJp3jprp+jb4yX0Fz3pWabXvHHls
thguiEnYHHW/dF0FI9FveIFd1DHp2hOC9sHjA6wXg9EpY4xH8+zvyOPb8jfvM9PT
bo+kd30Er3u9Zh0LBmGdB+So7TXob6of9vZzdZeJzE7LzwKQ08YVR1vnbUzgvDHN
wUdsqMXHP9claFdzhJpD8vp76lloZNVMj1TY4gjWBu7oZyZcAkmxUGuZYbp0UufE
u00NwlnqLAE+Sehfp6SSrjKMAr1TxDxRwLyQUfV/4vojtQXxb8y1/kAWc64fBRdB
CRUexEiQj9wdFYFRI6hFBY9wXGec3Mn2gFmH41F48DCIaY2H5C05TKIHPmO+WAeZ
+eH1JQQvPJAo5XZMXYYAlYJvgi5i9U3JPX6ZtoHNnCmflPzHOBij+I+8jeAw6QyZ
fNi0bPytNaFlhYvtwtLDQ3NhuFkiLNPj2Ukz/mhdArz+ysrzZlXP+BEB+tQriPxK
Fhrc+rVsqtTAt/WAxSsKJkwC2+Tb2k5MN38kPBKmHbAH4eTRUtPL2oifcDuraRmo
KvpCwFP8Fga5zH2QMuSemQYo8nKNQqbDOicxhoFG1SO1e0rO7w0VgO0OC1scgk/a
dtX0u3pLN49U9rvvxGrpjeqUJ1+8/TusbFgpJjC6bn/3itvLYSzpPl5hzjdkSfoe
4NKm5qCslOImPJzOoa+kUqHjMY2O6J4kt8FsvIDanl8lQwp9/TigHO0s5RotXcSt
q5xXlCUzAMq8fVbxc+TyLBbvjwNgaKbVAjv5ICPZbNW6w1My/p6CNPXQWqZnP0CN
Gr1iXAoFEYQ80XgPMtpxAav+Zr51iq836iBU2BKWkBz6Fadr3Ax9E9qWcQruTfIN
dZ4QUl2WHExJVC3r0GdMAddDjsN/2C+I9KpmzsZqVGAZOCUVeC0dM0H/KpzgxzFr
7CezjfdKTARtDubGbAtnR1wjYvIBh3vUlbS/QIjLQMSsuUyjFgR6Mh0TaE1PJvq/
/+EuJMi+6qaUvJtsyYjeX5x4jZsU44DTXYIs42WcS/MJcLLiZmzu4Y1YyjZRvTi+
hCJnbgCagxm7Pkn8eendeBAHl+GeNF96HV68X2562G1kDXCUDex7An1eLaybHkDO
ugiI5G106EXrwqV6B6AQpwJUaHPnvFO3jQQ5dGjWddpPMCRzs6fqXNba8c5rZ2T2
prqCtVE+7kpskPdhWXtAyyAZcR3lXs8jO25V60KoCXtWG2SeRjYTjrn0a5ch4Mi4
cyMAqaizAYdPU/+cqngLxAGLR1pv7jjZOmVMYpbzD8XeBQrSLXx4WYQMeHVCSwnA
0IzffiD0S6uYAJoSbdIadMOxxqYGI/D/SYa/W5NEXv5psRa28quP6RN/pnR/yZLd
/oRMHqf1Mqmeio5tx8+f4dylTWpsW/+11PtAP2yf1OvZQ2vabrVXFXrvXbMk1mzc
2oHHqA5FUEkGXNDACWlVorPldqQb+NZoYzeCLyN/qke7zdyOJlXmTVFyidFyJrfL
K7+wvDyAv336NuUn+4ehuKfrZUDySRQ2vk/bmXSyUj6YNNRb7ZHLviomDt56vmzn
yfZNybeW9s98BGrIyQ/T9W57UZMYs/A4Qt0UUUwHIhzX1KzFykbS8ZmgNsLvbeFq
O4Ioud5TcarD2bHZ48uXKyuicGNS3JiAdwFc1qEZdgzQJtBcX8FsIo6Ur9T1vvwc
P6lpAWnYnaVpnhCK3wocpDIB3A2vrOQZZdYTZdguAVu5zjvn9W/N9bS/Ii011UCM
AKvPRGPU7JHzVJ+Bj7DT0bBmWK03Rp4UPxzMR8P8FwJTGYJe3uIiFzEtMwBEiNAE
w+KcKt77IgkjwPogFkyr8US4aAIwCi8hn37B8qpncqK/uQyNuJIj6G7QZyMU8KdB
ljekNuJT+jJWr1UhNl1CkkRaT8QlDGQVedIY5VYJPRhlCzHqWxNXz67DXt0o6iqM
SdpjMCZfRs0W7/9frvDmeODndUPIBuxPoD5qbfJZCG4PYU667FnFge5BGF9WijDL
BjycSy82/pq86t2oWrORNg0iu9kbs1i4cNVunZuDEs/1ayLZ5Gj5cHBNpmhLaA10
jc+WO4RHbdp1HYh1+C+bPRHofUZ92W5QAC+7xyONPrMCrtxLrc+fbdQ+v8o/tWST
qqAMbxPvodUunRr2J38+fBZk9eoxD88W8APNZgBxBALcLDr80VSJ3stjuOAI/CSo
9Opn3UU+bYLssILS/KGBIAqAPahN+Y226vHXsP3tamfC3W2xNIxiVtGo6N/2oPaU
QLsylH9X/T85n/PZHziXa5rRwCy/h+XL8c6EwILsgLUOlluYCE3aUdTuOhDhuF4v
5tb520vNfXX4HzEIgBdrlnA4tplohaRvQxxILhTuiYJxNrkVdD+451fGlJHidjgT
VKKN4Q2Uj1+jIk19tFKrX3r2uBg6PYYIyZp+EehtKyMo2wC5o6Rm9XaFSN/5w60R
fIr1VPLI4x1+L3bnSlzhKSFGW0dj7xgg8tt78G/Sb+l1ZTQNT0Yo8QANHKIqrxfo
vpqyuBwsyvbx/kzr3d1DtSk63psMEHQJeV2BIW7Qx3olv+k/A3f1Ty1BckgX+IJm
Wg8IY1mmHcgYPy7bJ4KzMvdHFFKP9MBr0Xn33/sozkIbL1iojYicr+/z0j9/HgPz
B6nZzx4tXnQLeaJyn2y1A8W+ffg75yXonl1hXbF59Icyp/DeF0MU71D3VFe/kk9p
sqci88h0YFjPxLmDgoJXy/LKRzMgl0YsJcD6nAbS6Mii6OngoLg8RS9bKwTLQJU3
e9EQfHCCm4AnG1cBh6ZrQGMn3p/zJKRiBmNLtPyQUe73uc6HD4KZdJF32js2bEHu
GiwblecRY0xkrIeGudXbZop0xYgvLmi7pCiGM28SoTA2sVmQQCWoMrXqkD96zVck
1prm5FE+fJs0TlFVQcqfLB79VKX3iNszBx286KsaqEKAxGJDU8P41M3jcVAKjALD
7MsGIPPTQQ/3m1BjGV7+w3KhFjufDCCzhoYwZT5UXSDKXF6QXGVxSYbcN3g+QHvt
5LPJwftvHGydrqpQn34Zj13/sHlmywTxSIOP4KXBhusWZwhAzvDlggHXRSnZWNIw
gjwSna5bLrWl3AwM+dpQmEECIR3BrpHox1V0acF5FdkkvFP5Bt9+z0s4T8eP7gX7
b9WxkXKGFyOiNwoEjm4jB6hmo9tfwhYvrJ9F43+ja99Hxkc+frler6+wHuQyxTvH
hGvRDO1Q1aQlCQxcK6hcV3Due9xpYaRuTMn0FbKUZ4HTE+1flF24wHFfp5g05P5F
LeJpRGgIzbx+9P03JKC9Bq7ZNOWpqM/ZSnudILnBLjIl4c9629ykLqlHF48ULBea
OMIs00r5lXCh0/HEoXxZufRCzJYbh8WDVucuaR6NSqAKP4jS/E2lsGU38BmUIf8F
thOB1t7LUPVUelf4s2tTSPH9AuPv5ATvwAZp33JBRAiXH+WwDpNIl/cK3QBsiavh
9lW0y9j5ux1mXgwLFH2ZGcpkGdv3DA7dMXHyAlK2GI+3BT99uwcLD1eNAjRy8AiT
iKKfqwzlY2ETy3ohLCM1NVl7ImdDJ7I8aWSlpoRQquTpyEv0O0aKYRuiNP3iMAnQ
NFMkXSdl94Lr+jjR2KWir08oXqEAQyI/T+uS6zdQDf2JE7KWql3pEIJQ/kX4F+s5
BepJdU4A7wR1PbCE0lUVJ0d0F6iHUeeVJIy6HrtfaiYnGUugM0R5IKKA3ZXPF9PJ
qb2V6fUXzHKoUrHJ05uhLY38QM+NlmdIB+O5SvBBKXfBOgtxKls0xa2nTLbs7eQl
sTBLSwd+mibGDv44lGiy52+QZdz7Cj0iwzDQ2bMv66sGK25/TtSV/RgbQ96wZW1z
OVC0b8HuOZQGuNERx98y6Tl8fylOsdfJ768lce4NQVgUlhTr9UOARaLxPMLtmlZQ
C2WtG2A5wqXWqrjLNKRbLue1ZUtJbRPnlyIRHZByL5TwQffljZEU2JFUCCVNahHs
x+rUJ0nOc4A31lzRtaMVJ1COEawavsbLUEcZFsovIY+CeYiCPKCYn/mHwJPaXxA/
UOKutYPvbxyxZOTCD9UM0h8iDJx1g8HPtiLFQzLzQFv1ZbGo1ltWqM8/KN10Z7L6
QyFv/FssaCuynQWCjOiCqqZ3MNjkNe/AYOxWd9U97eBydoN1lHLl8hnIKieTKuEn
+/hlvsCAB1/mUZQxuH56tbMdsNY2vd1M+UyDfiCmgmh5fERHob03qxLrgQHG7TbE
oziyT8U25vfDgq/8XlGfd9eONKxC+vPzYPjWZ8uewQ6DWgOtQBke/ysplUL+rWIu
sgdexH5cfzCd9wxYevr/OguTxQXo+sqoHyyE/UXRDUak+GqjZkoCyk8PeUgJKDBY
SdKxh06eSPaH2hec0KBYN0IiKKI6ZsKoZoVDl1OtS9cXvfScd9cHrNr1aI414En+
AenQdxPo0wt2gB2MBM8bvLo4EU2R7DE+OAg3HhA/YL0y6IPGNJDACsNxYwAZAfWm
1vI58+O3SQINDnjG6vbU9RQnlTz+UoX1QKS/tN3mTIf+y5BE42E78avrjUIUxgHh
nE+uggxUAALaCzsQd2RymTeR0Y/RG/eCCLRRm2DvvG7o3JEk6yPJZoUh/r2zhtgv
okruXPxZGN+oMI/esFWeIrC4cx+tX8jCB6aDESPNTQOXzgUEs4vnIU6WdVcMOWen
DKVCpTPPh43jqS+WYA90N6Smfk2LTNCbl9rsrTfwjdgNiX4WzCy9t4oFBSxgavK6
1LfdfpBVfPxCnxnO90eDAOqTbyN+ve7GFJuw/j/XW8FIE77cnKc2IpOOXNmCXecQ
0EsxnQ9xZm/wuqj3XDivXT5EwZb5s0Fie5xd/v1Zl6c+3KxbyIyzIH/j+Gid6Nz0
bq5ilZlqs5YwJKhsLFsZWeT47pRvKmTG+aWtoM7QwOg41URSDILOv0+y4BBk1yNg
/ZLedk+fLiyO3xlyxLG2nFWrYeoG/WIQKreI8tmzy5TculQeoIDQmJlklBLuTudR
LBnetlOzkzsQH9R2ir5mIvs0xVZ/1D6CFwdDDrQycNJpLT+mLBrD7wB6yPi0Q+1n
6P3SPIp9mTZGWYg2x/8Z3rMd+W71kfdRy3tsReswJ3x41TSD6S5qT8jU/Cai/HNt
UPobeHIYK0pmJwZeWovpUxXH8Ctt4RrDmib3GriqiMXPMI/OaWBzybqoB+nnM9Mz
uybP6lplRI2Aq8QjCzc2fRqMK/3qa+LrJuvNkLIC2y66XOPfodf/wNlHfAlzsH6r
dGjw+Cow2rNH913+Fmifid6isE0PhR1NL2s6TKjI00zcRfKdTdez0gTKD06lVlkS
Jjuioi7vepGoON2hbQPQm+Qf6PUJIRHotqclL74zt8C6HETrgEHGMjGXk0xo3J4P
kQEaPmXCgkwC7WPLPTVqFivbpTelYRRvG/Zpw5ET9P0prpNR2RbxgkMLBgqZ9Tb7
ATpNtWn8XvuyRFCUky2J8A4R0V6QR0hhZKQ8sES9MuyeRtZHQZTpTtKNwtR9F1aJ
VoXqr3TGIB6NWyc9dlqpfW4s4OzNFBFcRgBksU7Y7oBygO7Hu0brgD68gDbBRUK+
cAtuxADJ8vkUvGGHe/B/oUAc0QyhuWr4Sh7O2AvD+mh8fYkjTU/f28PiPYilPO5U
J/NMKOUPnMs5qBot9fVAszi3oIqYshVuAy4Zw23oebuzHrK9X+G/lGEp259s7AST
e10gJjNvqaFmyFGw2/VMEy8GhN81CjRoCWXH/WEou5HFpzmC/mdn/LtOsdg++IuZ
Oh/goB9U63vhYlqJ84bILjEl1AUp+Zq5bY5H5SD6+LrBmOWvPMO0pctQnnfPokGW
5Rkj0FJcO+EkPmUfl6OQ2bRu8z1/0gLpsmwSDf1Mzsdvi2j7w0fle7CBHWVJ2nPU
6dpwOL29jxo5y6UsyYvk7hrYQTeSiICZEXFhnG/IX0UwpO3bLasXJGRJR4v7rQx8
XqLSgcMsKu26AZzaCiDL/dY81naM4BTjp2LN/mckNJSsY0ekO0sWpQDRaiPGy1yt
q/XhRbo8B3IIJ+9Vsovsy62LWbpB2Yp3QWUTv+vrW9dHjDPt6fc4fQltdjyUkDk4
wuANvLGJUjcl41qXReKu8nDsjn/xVJfi5K5Ncs2GC6BaFuTBWyOMr6OmmYhV4ciW
qc1W8sCLE15nr8WAd0WWcXfAorcV53emaxSYZHivk8gTVX71LAdjfYGj4+U7ub8r
Gt2RhciPFT3J/4qnw6UGfpPGSP0l2mVwDWeZqImB6ZacT989srzH8cVO83b3jMNT
oVd1yESvJmmi82dC7wZK4YkvRwRp9nJEPz3Pjy06f/D++ywcTveE/3QaBvqErIvJ
c9ygR4nMMRcatNx0tqjJCoo16FwTsn5w3EtB1QVHlB9MTc9kMvNwMvEHdfbbLheW
w8C6dlv9SD/AmOtd7+Tmu05+RSp1wUKaNyIKzWNAK3VZwS+I4fN+k2yt+EdTo8pu
5rkJq8OFW1rjSEBifmeq0aqC0vH6x3732/l1naXI3TkHIWZb/dDl/7dkRKEeHptX
vThtujmsGFHZ93bYww1h9sps/LXMhpAOpqsagZnah0ZwyLdw3mjKq9vocF9QTodl
oHYvBQA0SvvvBrD/g2uLn/v188NP23ZDdStjPnf1D1dHCaVBaAWq17mdH9aVRZ8i
9mMzpDpvWbOGt8weAMsXy49i6/vc21sp5r18SAssDs2jTQRdr8wAeq12ZwdqGKp8
hfBtN/9yMjVkm7gIXEO2w/VIecon6gPM1WHHnaPhRaNL9TXqLNFgRBLmxBUwV9py
rESct4uh17abflAITFWTW+EJrtO7Ujv+sxCshxhlZaE4tQJNcIQdiXra0n5y1J/h
ezWixmjBveim8bs/VsZehLSkShLpWOXpKDRVL/Vyz8Hf9eAPiOJW4YyPY95I1Oa/
gXKPxsd+E2hxXeTQkn4PBaW+cDQlPAyVBQoc7oTTxoBcwZpQ/JMxVC2LaUmY5yAl
89dpGZobVXQHmZvmEZ7BPuRHiR6NI7oKw58uGqQF3nJvN7gSG7XR+4yC8EH3hs6m
pThWRywPW+ZNQ8xpUgLXQE1b7G9sSUXm7J9FeuIQ+diINkPzZ5mINORvZvYGtzto
mbdfA6zB/n0WGqGP1OfcwKNwgZbqGvTRt3z+HaIiuA1Di4BvsCuUtsyQgztP+syQ
d0s52dl9nXqlq5XDrhOxIT8c6tZ5gHwHD1qm4eB6ek3hxG5aevzxv1a7gtCSqWz9
N59s0k2uyLRq+5AQcb4KZstAAeG4YL9z/uMPKZ/q4G/5bHhf6om/yfB3cIwJAFsH
Lw5T27J/sv2c5E2ms4BK+pgDDRXq1rUdvgpLoYOaDQqbbjtstRWLPQndfLLp8vlH
1qYNH1S34nhqR93mrSQToGCNnzSi7IL/kqBupRBQXc2aDT+qc5juJAzzCU4RH79a
lPkWDg/e4STqiIewCZyXuf+ie0nhoComrsEtNkCiAwb3HqeTMT9dgGm7b671INdy
pS+MVH3dLYA+p4fSEQ1tfT8BwJyOS5592frmKdORd2bnRpP3MFHHcbiZln2EA8oO
fMSXyALziOzEpkDu/96vMdMKl6d4ewrywmpYEHglwXIO5yxRRJvqYqgjoGdWiIUa
1YVng9A+rk1WS2Gk2KzPN6wc7ZeaNH7VEtYDI1tvNyIsX6rO43CKkBH3raJ+qr1U
U7T+GTFFwLbZrpbcMiryLQCgbM0nukgM3R0WSj8uTXaVCj8e55o/0T2Q/ugHZKN0
gWqdXh+Z1QDirFKJ5SPHvJQ6YoFZ4lCg/C+hrUZcgH2uRgKaQViJyOpVgMn8DZuW
Yh43+fui0WTGCnMxC1mA0RzPvqWlvGCWtXswIczVR4w7slol7iDbhzFOU7hg6gTo
xxLe9FnroTxZ9c6PQIKvu0tiS1Hd3SnDSNLb1u8epZUFozVe7BQaGaq52OfKCk32
Pq6ABd9//aGIuj3I89dFn4cCsMVUJ9iapXdb9aAo0D6bHiPL9yYQLifYNvjm5Fv1
mXkdwTkuz3ww0ZiYPMTkXGnFvB52lS+bnCabcGPG8i4JkmV3QRH4dJzJxpwFwuQh
5wk8RYtbWYcYeP4yUlm/pZTGeEwHg/I4GUpTd2RTRQ5CfwPnfMtGoqVHSe3A2GH4
hdXmk3API4LFBYnRP0h1R1naSzY756GGjNa9bGCqZlhU3D/NjSIdqDC01wKjcSlF
tR+TU2AplY0HRcLABKq6M8IXBaZBnZ33+E5bkaH/T3iNCBbzG33rMRxfcr6PvCCm
mQpIDRkyJNgJbJhKsG377t4HJ89ZrqoY8TuBR8LLsVbX7sdad2HAzxoUjEauxBVZ
3o2zVULPKgv9UsDsGFKZX4QE7sWCW/qLrT/tjaBZGdF8PDTahaq9OgkAtDfH/w0N
seGW2KZgeNcUIHOJI7BAcBtqhAYFzfajlD3CCI+CDEv/bQWKYzqzLASGpudOGto5
wZbjqYuaNwIlGsy+6YFmHme1iZ/YuT0Fh5wKDBloRSIIdcCUGcW5gmtmZV7kbh1x
jC0vuxkTXgu7dsTitkXZD6RkcJkZevosflXwLg9ctCR9ivwdbo74hWyoy8q4YHyh
QF+oOFI2/BMiHTsliJM7c+KefB3k2HnOdPQEudB8jKK9O0rajiPobffATsual20Y
ivu/SK7jqq2SmqOKzeVk61uPvTdAJm2ngedCEYhUnTloQzWfjVWsAyKzotRvSCSX
fX+Jlk9iArYRiA8MwDjDml25xBsg+G+d34vG9GcQh7w72ZKebzpTR69ah053BHAM
L/9gau4EKkSfJuhCR0MV5x2yf+Xw25CrHjH3ABfqxlW3KaTu8DOcW0/F437zz8hg
cZ5XOXlMWu2ykU0QZafseF5uhsq67VZjbShMuwR8nYEwBEcPCztW9kpFHFhzy3nL
B0/nWSuPTg4LZTrfPDRXQ6rfiiq81YCJfhYKMJbFuVOx0JDhxDs/c2vpwcx+3/IS
PfnTTo0WFpVsqiBATKRSYKB7/LLQqSF567iXyWbkAkGzGu8fQwMeko1UcxDSXio7
UfPy48vrjCbLiFdjwqGLwaaNjeOUhEnYjvXC9q0mvfmFy94L9qZMJ8CCEjEecw+m
LMEFSPk0PI3mGG6NvNjARI2YIjrFzCPVBVsfyBhchEkBdon1lXwJpT0TGkEPZCjM
kULz+LXsxisriDAZ5yUttgBjU3cP6aCmIgqnZJDN7kkcP0SEQ1py+vX8Biix1mNS
8HO6KOoNmCeK7o8m3dC3QzGcWmu1OzfNDIY/pwiGPLQVkfcOrtXHZ1IZlSeqfK8x
DK8k7lZBBbA8IlQuKe7BiUpIBb7jdxUWbFIR6uGV/qoTGn0a+XaEpJmwLxXfnwKj
cK7wa4gkaAO9r9igZHWF25rZMaskRYqOlb6oC5PIUVp478URFlkQNPR9p63O649T
QhCvGFyfhCkigncSsc22fGvLhp+AoNB3O8a3blQ6Lj8sfjrwl7kZvRTk0aB3jRTA
utlVT4L/SsaqcsK8w4MofCdGQPbcWo9lD2GvCy2Y/zY7pWYaZUxPfAN2VS35I01y
V/9FjIb44JeW7J/EOC5StVbv/EyIkFOcqBcwTTM9OhyXHNwdgw6QhESC8pPiF3Yx
F64YDfUdAdjkULDtT3TLZJrpY78y3aSo0TkUqz4tIcFOOYrLI9AF3VyjjEdP8KvM
FqsKGadhAKuYZvmGHgQQi2BZU8sypGv18N2t/QY7dg2shV15gpMueo9NrOImHsiJ
eMYrc/fX3IFdZuII9SS/OCZGoRmcbfVQfsECx8fSQEtjWrWH2QhUDUVxcVvDx5cf
E/yySGoVb8W1r/w0rAbsRraKGqTJn8DGZLz5Hv7TYhJG5WVTmIm8K1hWpnER0Na3
IrvXapTE+WCNVIYI820bc7pVSQ9u7PX2yVzv8Lqn1cDKkLP78J4+emjDfuVwRj5h
Kz3HZjtk7WRSh5mrBi7PE6VGLgPc/nG7thn7rr3RScTXUHcFxHIcmhQxxe3BXbCG
utCmpE54fFEAM9lgiubbXFsy8Fx8WntfzhIZytjxlnjZklodli5Vz8I0P07FybZ7
FsJtIUIQk2+exlSPNihNaB7vlFmFg6nns1vYsjLmcsJAcJc4lsdrtbFGTU7tYNK7
kpe4dJuxQvgnpXbh3hF7B9e5TpyCsk0f2P+uSwKvie213Yg50Hs6HJtu8GdzFlMA
iGCJT+oqcPkDWjII7OPuEwF8IwibKqRlEbDpw+AgvmWbSK9xtEWwjOwCwGNm2Btl
Qv9S9fIpz+FqjQSnXL2C2XCyVDhkDzexX63QAReScu2sedhQmlrR5rRp+XQ8qGEY
nx8WXYqSikoxXZ9Ds0CxO6A3wGz7wLGWfI0Bdr/SSn8m7jobesGMoSBbYb+RD/Zw
pN23mBEUtVHBlWb/b/F8S4ZGKUF/HZFH7NcyGTfF9pFWswdlFvaTJTF5e9q+jXNZ
oHBbhsls6oQ3lVYuNtrZ7mf7Xh/i65PIEzFOij/Bx316eDciq7v94GyGzlUnfziJ
NAot+ZDzmbwZ4p4a8X3Rqhp7DBgG1GNnoRhwe2RS+Wi2dM3fKUsa87t+NK9Phl92
ym3MJXoHzBoaWhZyKOwA977KvVwzSI5dS7Ma5GPfp6r08QsNPW7qjsCB+WTKFwq9
Db0S1Si+YGc6s50PK8mDgHQDxqZYLWI2cp1lc+Df+2T1TG9suLuefVc0me8gqN5M
h6uWVZcNkc7ncPRbSklZrgDn1gvNcLkLR3I4CFTv15Y8VH+Mcp+06NHHRmOSSrqK
MfIRY/HRSVCq8o24p1Ki+uzfzlN2az7L+jjnE7+B68EFQjkLr1mbEmI6NnnX8r3k
RkD1COihYP5ReMYucqB9FAdiGIQ2aV28N3TzjIK5Qwu8ROFeTIxS0r8ZDk5y3/WD
WMTHwXPJa0RyolimT5u7doIWmWFn/buZ3soOSWQgHqyrm2pHvuymfBXLOpuWpZgm
SCOdhMfCTw0zARDnCTlu/ntjuWSRmFsBg49UpG/GUKrwhZcs8TDyAARA28m4d3oX
T6actDUVyg3AHk1iKIJhPM2QsI8T5+C3gj1cq2wsNMFTB8TcYIsqiEe8h4Z72NIj
Fp5uUrJl+HcAfe+Z0Dbh8aQ4MG3OS0+nJswiTT21RRBuxP669DrA8ssnT4OVeJ5H
zroQihI4p1jUHGwT0wiTFs7mFgq7zzKupbt0HY/cl7ULjx/z4cDO4XzTTUpC0POv
V+oLLxiePeSeOyST25XTMJ4phyQLVM3cP7kwYxv8p1oIL2Vf6XJs0/dHBmgDOiHk
fvHwWFYhwHfwIp44P83BFCAecwKtf5BhDVxC1dwDHOT1/F1fbYyX9N/B8kqoNVUj
SNR2OgWbSIWBgo2YKI7fpKO7kppR/uvcxaCMmiJKT9qC29Tr9lM3q/C9abvmfT3v
MLY9Uo3T2+T9stL49L0LYYRHVKiuvyNT6guC6BomfzK/5Rso8h28rnC3kO3yufZY
yBZG7VPXBAUQJ5QC2RatCLCY+80PrsB88I3MgwBweFaDUhpQnAln3yD/V3nstu53
R2+sHQMz8btb8BzKZi4G4vNE/2V40TpQtGVivXKpVYHLcDeT0hRNjlUX3jLpHoOR
2iasBQS6ZVRP/RqA+ka/BGibXWoAIbXVt8isfQmMu1xDKNWflaD4rBxHtLGy/dPZ
nEGNJpKWPSSY7o9vRF4jNSTgQM292tUBLtrXeC8IbCcSJYH+9jJWzxVL68tLlFB6
gZCh0eRlhrpYiMZs56QmO0900KxeZC/lcFa/gf4ZqLlgyD+isK9CWP4BNfXXmJnc
2yWgw8vp0gU6jWfryU7Jgzv+50MTn1F0jSPuw+T2PRWF9X0A0GKO5Au8biOuNqoz
fu9GwCDN/iI5miqZ0LzG0QTl2jODJy/5Nv+Hd60QqpKZu2XAfDllfWBgYn957adu
GtwQE6QZPU1a6HoXdhmSF4X75z7HYKGN8d9rDj2J2JUWUdY6taBhSG/p9p2wpDPW
79cFseCu5hJuI2Hf/+qtcVI6ZN1/er/n3lHbMrFQR33+iT0I5f9xnkmccRJ3FkmH
j42+fmNPbgtiumXtLNzBJigZ7x6uQMQtkmXmn17nOqAbFxXoCTpM7Or0b7Ia+Jog
6MW0Nl1dKYGWRwjW0MhnvOkRYYxlxv53fyIXHmWps6aLr/5/C/NT9RDXCAU/OuJy
sUuEAaKh/JNCXvEeNr7xM7iyj74SO0h3dGtYOvzXwqI3VRQvtxb0wfWFN4nvqYcd
wQS5TnrIXD98cwZDCJlC7EEOXobYoOKxWq9lVQ6Ak007lfsb0eLX7wAIDeT20y/E
YVMgaP6nBHFF+eH0qBpaWWuiZJSXNlad8cXXQQHrXmnKQki2jTNFno244VPgLetw
smvPGyAJUxmXZDVX72MDPMphCkO8a3KRxLbWSGDxOWFpPP0Jd7mGabSeU4plJ8/J
byvXRv9JkD9RBmuZqUe2YkSMEvuyefQregp5ovA6kHTWJ6oXCB5xZh1PRAn0a4uU
T3hTHfYOC3pNKgtH8CtWrqaFDK45/v2tZF1+6U/W41EjoF/pK6TGerx9Tq1uA9xl
UJB1UDBTof3sqUsrwhfJgDwV2TqU/azBvixQ4JyBG7xf+mTnWJDzZF6Jmorg2aK0
FI1tUkWl+ZJoVoOdP8wKC3O/Zun9vzjXttqjhp/iA9kOWWW5D8l26nc1+LePj0VS
Usvvz7ylVppj0tKN3GHSWii0ChcFDeD4TOBBBUbADXuO86q4+yt2BYcB4Hrltcvr
UOfCHM6jH8rlEILQm+f2NuhllL28vVbBz1+B4/08kYcHMnBoJNiHk1I9KOhZcAqa
V2DQuKfCFZ1Og1AULuyHnxkzmzKTctjCHBUPAAVoIVbpwA/IWijir7tgKS9me9Mw
UPVdt8OQX6UfqW+ui9bfjakGFflOvgpTVtszuUuIJfC8nO7BjDHBybhUKvmcgqV+
lfbDf0g10BlKjqbC1AsjNPzlsE/T83VNSEqjaLgGpXcefF7SGes11fB2epRDtQuU
etxYBY6coXdgm+Nje3RpZdGNBQDC6wTO+Eu9EyP/EUaiUBraSuoJyKkk0TOSneO2
kqP2I53rNvXLKTwAQFWBII3Mg1ORfxbAKIbAdiLCJhpqvmTBviko0eFhKLQB83ES
aTdZ6uaof5/jd4J+WE7b6qHpRPSiTqftthq+M7BuLNTcdM2s4gq5DJJ1H4p7UyMD
ZH/hj8sKGOpPgGW3kp2vK2O9rovD/ALZulEWC2/sDBBpJxosQsY4z4aQ2kWgKL2b
E9U+6pSVs+x9LxOOfRxV/4OJCRHdeTKTdqXdWuSSUiNIV18gq/AIqiNyqcn2Kz/O
ObnCdCcfTkkcG2XShtUCSkmwQ51V+9NjRko/aaztVJf/0ZF7MTLnQLWzngSsITsJ
ayBp+r582zT6BgquXtXY/AYENtJ6BpCSiH/i/nu2TZfCXjIkEVKZTl0cHZsjCpq4
/xRUZozDqszips2SvvqFc0KZUkYdX/0sxSOpv3X6cu3HmufwNRxMpPxlHOgLmfeK
JW/l8yryBdG3xnmZFYq85amqXe5HO8J6bnO3nKMYwXH//qcGZJPpf5YDhWTL2vV0
OGL8UYL6IwqeU/+U/jU2HCUn/v2bR9YAp3TnE+EMUBB+sk9HQaJ7DpHYp9797Dm3
YZkzyAu8OuzOIwowxgLVZBnIuqpgY0+FDM15fEhkTENch2gJx98ozcT3TbAIYiAm
fxBHSUoGbT0HTTJ6x+MPj9rrH2BKbGRbw9aJzLZIlNTHnvExOVllWbRnpYozOVCS
pdjCB9nM2hYkSUAKjpHQvC6q5WllPB9QrW84Sz+LjMvpFqiyfe/y1PRzsGKb6PD+
35ANTK4kEOuSwcnBQP2ZasBTiYzlF6A2SCvIkP2LKKp6sCHBzUJXrlEoOxlr1tbr
fkt3Rb+fCfMI666Uq3dEfhkaip/CiVmxKBYYL/vJA7vkTu0mwQqkvZh1z2XQ4diZ
ibLsK70yH0Yb7zddkP8nS/ataCMcPMfcefEBkS8W6G9rha5WHO8oYiEKMDzTIZZ9
lsEPcb9XjYf8DYGA9SMTrsJQpy6GO/s5AXGqSOqpZ6Rvop9b8MxBGP2iiVIOy71z
Xuxyo0KC44KknIlgv+9A/Qvd6QjhDwnThxyfuY/ikp7K4TlRKQj1xLb+ctpFKzhQ
iml2NIUzt/JdeLDPpS399Q2wI8PbYBS/N0FRZKKa/YUvxMytShseumRFSSTtYcvP
T9t43Kcpta+90Hnpr9AxC2trS/osJSXUv4ezQ7dP0EAEwniYNtsl69OMEtM2qD71
bgzGpZvvF9k7h6e+CCV+grsh7BVit4j124lWfalM5MgQ/nde3+w0YY75YQt4RG/G
xo0HX91cYVYQZTUT6KMwkm3JQ6Mx3Q40+IODGpfYGBxetaLRihgjyzlOTOYMJCpC
MyRwJ3DgIzbtFqWsiKBkP2ZnzmfFrDAnV5L2EJLF/fJlLSOuNDSZKgTx0dug1Q8r
iQeZkFqIzsEpQT+9L+4pPN7H5yfyTOwvVXLBtFAcivUw4oHFpmrQjBrMvDPWGEyi
gCusb3Sh1yCzB1J3agDy5E/xflUjKJJ2BmlWEMH1phnodP3+gYTCtqq5IPNfovoB
azYG4XN/jWu4jcksiVSBTGLNWb1FQ3IUjgWlXSTb40YZopM1wEBcdazj66RWSBu7
SfRyS1+gMUiOYRPhlTFXeg0Z/ppWZ47lr8PYBeCmob3tlt1HyLczReAo5Ox6yv08
D1mryjCYqi5A/yZlUgijgwwZ/P4XbQQvPZgbyUjmcJtdkv6caLRW2S7ytwM5KVb1
PQshHcWbchrRqvm88+4RBFzI0oPkBGzKgwlqvmT97YSaIAEQ1xpF6CILO4uXfbpB
I6qnU4F02RRrZRh1K3Oa2HcBzTk579Vnw7W5m477cXbAoyW0ukqlVd7T7TJccEsZ
ApQA3jR7+dU6z1PfKe6l9mYcl/F7GWcu9wwN/8uVHqJu8cbSzzUJz84S3vSCZqze
O6o6I78Bd8NQ4lxSTB1R5kuLcoradSQabQVd8oo4YffeJE89ezR4MPKjS9ofD6Zt
7FNtVNc18zgS8Tp8MIwISROvQ5ece+n3gf8YfDfRx5o+SDIq1xXQNpMdP2jttEqx
DsLPrGh2FFZY74oATH2UCqqGqPl0tblFIXWgCthgLfhMCgiNwq9INH3KeRoFsz+n
K6GnwQ1RVf3CbWi6OhdGKDE3KkwvT6gQ4oZ+BnZiF8xwG292UtrlzbzMdcbAMAA3
4MWnEpzi/q2o/VQ5sZ+L/pg7ef6Yh8/WCKctA6oM7q/qtkDt+DI+AZiK4ts3I+T4
cb26wJiLcR18zCYy2wx1O4dkISNFxheYBjEo4qb+1ozvWV6aSOb187lRwuYlW9PV
f8A3tpJLwZ0Zl3GJBR2QhzUTEaGmGvElpiB1sHEWUod5721QXCr9XKLOVgJDiu2l
Z49pPArWti5fWBDNPr68S3O5dXy6eIt+MdLXlTZE5q6oUsH4qmC8WO+pzRpQ4OEz
QMVl1HDHgNCI60C92qfJZAgGXhXOhhmkdP6j1YGzTp7s7hs+eZN2eHhQxWOqgran
75Xr58y1GNFjuP96OmtxzEDQLgDBwBOcnRIa2YkmFIjYTSol+5Nd1vI61jt2XPko
xk7ul6+0fDoB2+SEgsdMM52TdDWTNzvBttkZTFW5wvskyQqmA4zqqvs5J/RahCIu
iU1mWwvZtDvmegv7OsoTnnaJkNFIqWEB5npuAuEceLUdX5wf3VCtH8tFxPT2R8ie
O3/BcllUo6xDSgy11o8RGSOQzzoa5V8/lglExEEJPX9/1Fvg7ZxRIDwUZM9dUQy4
+794X909a31XeB5l2V9tuQdY8eLik/gc6fD9OPsbSt2XRdQsz7hSG1LAVC+UEW1t
68POTXFzu3HcCGHeCfRz0WRkeE8cAfktChklz6ZioKoipLakjtCrlIpUQTgvXSYW
ASOHMMgB4cRGgOIwZJ5Pu6D0KjxGqe6bpBTZU9ok3v3O2beJPSNiQkInVxWGfvBR
LDh4nB1BLtWkKIyi3CdwampInSN0G3MpHIstVgVDB3R57mqUq9cCEXidMnQB7Mta
DBHZ2T0ZZ50BovscOH56w0of2OIP7SzW879DyQPv6r3DL4gpqSEB6fd+MbJ22ja1
0jHFBGy7rJ2fM5gx9rIgbMQfAmOBp70zMAT1of6gOOE/XmvSh7EnPH0UIhmNnwbk
/d6VEFb0z3CRuRkeumY+b8SHO/9V7Xo51F2uulucnLldodO9DzpIvUj93QWj3ARp
xlRIXVpmk5uxrROtU1hBX8you4BWmKlZRmC5Ruzj3qIe/ZgKtnQarcrDH0l36j+6
/yE/XKpUexq6B3AZ1NAajXrt0W9lxz9D7vN5JbZ2fL7lJUi05sLZpNndQJkPlg+H
uzJWHSs3TWQQIQopXFt8QRobH97cFAf8sMoE4GEyY0K5MLkykpZEatMTclgzDHxt
GYCBcTLq2Hyi26fHMpByGWZDZrXQV4Pq4vbPv8Ho9uXiKKMEeOjRExRdWR1GOAtJ
nIQNH7N7E4NfW/yfXVrqZU+MBvq6N1VvtkxoEXyVPlWLhbTMEtP7a+uiWsytDV7r
gU8cQlveCeIwc3buo3Zk4XxOWhxBcYr14XnP6ZuJdf2QsDvvNz8dWDiZfPC+asXJ
hLHJVKmJ3Oy+c1hCH/Q9pjGx5pDQ31N7RYvRAePcsEh2FKdab74nk0MpUftie3Gg
nu/XJVTw36zsFgPhMci/TtCRsRNT3VCj3SkQfgeC/LQXBXormGy8KbOXtT3dLn2T
AqhzyzC1bIMLEBtejVQCFDK+847t9cCRt0p73oYFdDXjqJ/bqckcSh39kJ4Ja8Dq
gdGLsM1qiGkC3WwleWr/+gon8pHVQDmQP3P0f5h5D7vfY0oGt135peF6gVCmj+DV
7wIkHmrBetAGvjyOfzGZnaXgrZKIpZY5JYAa3da+ghht8dX3XkuuogAw4OJJTqP5
7YTOWVg642feoGLd5IJkRHyMzZ+w9bp4Csa4db2Gt6QSi+M2HoJyGC6byxJybLCL
Oh4/2GVIQT0xIXO293UbQfz9SJXiX2vmk3J1aKkserNyjDSZnWTXl0BLd9WHD904
U4q7WX8FXecFjwpc1JAT1Oij5DdXTzpCwl/zGfGRBKZesq99TsLnGF4er09gl2Hk
rVL5cPXQ/oxQ4LtjaGCXQLuV3pOnpyqOgw3wqZUVUGV5YyUNEQJPYCU7RQC9OD0n
gbap7sYSGmnM40WtaTWBK1GOlE6o7QPz8vzZYvoWl3+yDSJD4fH9BSxCF63UKJGI
RizaB3l84ox8ZiotX/Rv8j0xTQhWDQAO1Y6qNq8pDJXy0YKx1Cj/j+w4Ul/8vqu2
SG6PpW7Yo2cbJBlnK6ZhWxz6CUsWYgUGZ664oTF+S8Wrd0WMc4il8CcD3S4xkbo3
K6+LtqxjjAE9rMT8lLdWLFjm4OryPdj1LV7KEcGr7XatWh7DnPzGA8CYMzr+aog4
u7TGiOJnLsq5EIRJNid5eABCW1iYeq3iD4DGw559kLxI+fmz8cD0lLAZXhFIyVVh
7WkrShnnzjiv0lGR3B4PIPoQdJPVRyOQeb5n6qbcs5rROmkAW5w4ed00ekskwgR+
PXSukoQCnm1B/2XdB+OMf2C/YzzKAJ44Y4x0PeutFJAYAsCR/1WrCY67l0/vtOC1
ne/H2tvVWhClcI9WUZ+kBfTFrfDVB5mW5b1xEa0AtmrenGUYe1bengS/v2pUvMZA
s7sYWYnAfWAVZUy0BzaOZU/sAkdVVf4e8qTXQ4c59hmMwTbDNiIOfWMMyf+uviyN
lTmdkFtL3vTkTOEZDK8r+JWzc24uiJ4c+rxcvlpmbdv+gABiGZ1+0DQgvpni3JgZ
esby26AW7r95a0LGMYqKh+2cawgUzBJQhZOC1uQJrDZS3K6tPdrn872q9JwTCAJf
nEmgpfdo+23wsEb0/T012dKjlmrX/LyJR01ZcKzce7HdlqQKKtN9TUHFezUhbMxI
IrptaLxiiliLEEKIF1IZh36qVPKGgGqIX7uvrKKp6uVxpcUdm1B6LgGaNh7cr5IX
NAIuOopGetNX56XgyuilLKHMB2P5nu6OHomzqD6C1dOPSqE7mJlTgXEGoAGVw/0D
Lx7ZAn1lKMwsemCoTr/VEhrHdj5VBqwUzfk7i1jm6c+DmGZqpBiruduger5kW50m
8nItCTL2I3uZ3jNkuWTUWmNcchtAoYO3LlQ4Hs5blDbNgIRw/tVlyAVyIOTqxHkO
eRQcsCgU7qkn1XyPpiTdN5TgwwN+6svUv+XIL26YfBgaRoaRGJ3i1ugm+SNMSMsA
jMbSu4sxh1ejVam0R+XcFE7rNrdYbfIXOcEUb25JbCdQwH8zeOyN5zAV96EpV1dE
hzbgnEzfTDGSoUfLqeCv+Cw/Ciqeb9ODQeWsp01lerIqWfvJeHw0SW718yIDoz2r
LkFTBn2/s9jtvtWZFj52sal+KYCCos1Bz9dmH3Dulp+sWEvWQCIbNwGllOQdHCLG
NTzU8sZhcH2zLuhXfJ+du83M5A+fev61myFRr5qhg2arnBcPWoKZktLS5B0j1toi
WnCL1MH1moQmte+LRRvEgY0EPBb15olmkPczFRny4DncBmFZyfzLU02p59Bi6Ngg
LEFZXltCzlv6hU3Ojf37rAjZDdJrYn0lLkUb6osxWQ3TVhInb3Bm42fF7EuYQC0K
kf230ZIMuyrBD+zQOIqHKie1+QBlSoQbRFC+nqoXFUGgo5Jcf78bZoxzDBLXel/H
D1VbOF1ZdEAPWfG/WKTSVwBWOsGXYwrYJ99eApPMqk2sIuQcVC+64c+tHeMr9duF
gQ+8ND1J+f6Qq9nhjECziR/XZq3Hb1ZyO3E/cqXh4BqVmxYFUjvn3dzKtF2hpzVv
B44vBWo/nh09VZBKjiCMV0Ti3ISadcCDS1CBJss1YLgFIPJ4C4Ff7nchSRvLZ+L7
XW2pJxBffXYjxQ0G8O+FS/d8SSBsyAeHtSPY8QU5cgIG2sb8d3Be7s61nJALMBuM
EKnkaqkxrcmhuorbXxQtv1QiTqvuTQiHy7MRo+7euZ/vCD2iY7wZ2zsWwiqQrPJP
L13sgy9q/1mcOddoTbCT4ntiHcDmHaTGn7z2kSQ6DKe/yEvyfA/Hb4Gug65d7SRd
zVN5mVBQyX1D2p2U2JsYQ2OiSBfeGIEmC9y7aPRvcr3/P/0qUn9US6OyuhHha6Az
ozqb4yEANFgPpPxa6LLklnySEdwccwqIKaSNW8NZWmgnD1hIYbBXq0eFWp7xyoep
tSukNNaFPquA6HlVWnmZYEzGXqB0N9yeLHcvJtp07fJK+EMGP4lrfA703KefBSJ9
kbY6VUB9Bj/gZL1Iykk6yMxgwh/xGEDGZOxLn5g8NZ+Fr2vCYoxGrg7CT2PHYUUC
UPnK/3e1TWq07zufFG9W68bkY0oCiToyfO1f7w5erUo9+VDWvo52Wy8S99bPnMtQ
L8OaV6cjP4l2KL166l8ukz0RlB49tXGSSY0dpgh5Sj7Sq0WeNi3FsvuDXdJQSmQD
MI4QsUcbJbY7F/IQSAx6anHYA+bcE23a7oUTnyL6rw1KNrbbmyjoSoihnJyiebN+
ff61E5EsrCk9qsBPkP/+Dh3ESshLJjK8Rtt4DsCnXHhW20zb6wIXTSXnNDQ/4Dq/
4zmmfkWq/oLJQ08wKAcRHMGGRfoCPem27WHMtbcwB72JUf5iJDgnwArmT4MT9cVS
7jP1AaOHw2UGjx+aine/9grQWrZWtybf6gNPp7WTS5vBbXCK98EgLj6mpObd68ZX
K682bwzuLA//N82MPYtovkGsZZZ7/c4bS8hNlnxaYRc9v+rOKsTUBvty033azr5G
KZUYYYPw5Ik03sKGgWtH3y1iSdr0/Mzvl4iRTtgVMfG3NdZNH70KjhSiXPUgk0TY
y+Jt1KQIjl08n11/+AMmu3/eYGUrfp1GuJlsKGy1dZGXs3cpJc234rtPLoBus1/0
JzIXl0FaVeBWzUK4K6tmMYeWLVK3LeVK2RO6X2WBqKb4VLoEqB3M766y823kYAaG
dJa3wJ8Ffhc0rC+QUa3MqdOoYs4tYDjIgQyk247t7vJK6d6RJLyhC6YreVjlWN6H
lhPDdRL43OG4XTPOdidO2xXmb9R5YLqKoqDBGb+VM4y6RlKivxCfsHuBsit9ZCAw
4eq4/dZ0ICzEQHlL8XKrTeCG5mvHEPj5OZSHCuVV3aoFj4hEu9NlWZIchYzJK34f
4IzHfNCbqQp6n3Zfd1QiAHY9Fl3P00CMJy+1iTAXOySyCEML1Eg2dvqQEfvlPLnx
HaiPLIdpkrJm8ze+rQ8ig2hUpxpuo0fJijpclpxsRKgUIMfackOfhDTIfUFQysp7
lyKUrP6M3U2T30oRoA7Vk9S/6su6x2SEccxTHWjbcexk65MbUoDcorQBX1OKc6/+
D+nwwBVxk0ukS67bZ7gvG3WFQZ5FL8yzTMkH2BgDgPuSb1C8Rtkfy5waVCTu7RSr
QttaFQW2u02f+tXQ18ARueEGSqVdSl9Bu/GzXJOMHFdjRxctPHVBOU2MOu2yK9Ko
Orr3uOh/dkxdPH2EMMjSmjf9kNGGk4wPpIEr0qIMdNEvFX1b7V+a5qk2cMSSBWWm
M75KxHPrV7NuIU0eksknGX+qTVSh46zjM7k4j5pkfbfhi3opdFxnpn2GY39e+sQD
xoLAP6IfeT/KrfhrTtxhM9TOSIvbh5/07flGsx2ZzkkRwob+yrgDpLNiqihPQJuy
ouqcrQe3qKOw9aniLM3d8jp7oajrBzq8MpbUrp1yw79NfiCf12QuorsxzvXGRHlt
WF6YWee63l/idOKRBDLNQdGrRl3caPkC/7u0tY4piejUR0qbyeGebHf3y6Zt+oeK
dQNVh4Y4rgFL1hGliw3aeS/Oy2apir7MmHma1mzpWHH5f3CnbtnK7lF6qoqQxb98
6TGoDVMy+0vBEO/yk0qcWOsEKOw36qPRUJVmDhZ+Tgr938tU26xEU6bCt8lWI0Tc
6ZVCwujQo/gzyYFd+4WKIim4MnyOWf8cXyhxt+DInxC0n9A0LWoIRCeHIP4xuZTq
zbtwcB8+h8PZpkFysIh7+Ckk/JtRddkWdiGhP9OXRhairEc9p8OJOiVjoYn6lBcU
H1t9deEojckqmVH3TGXV2Ne+dQiUj4G8TzGN+vyTpVUy1WqI18R3vvrKz0eIyFHN
sgI6tgOkhfWbZ4YUDIi6ncHB0K0z8PbxBSycuKt2RnSpwifENS9ISiGq5/0ELuNi
33iBVUWBqkrZEe2KmdJGNa8yoGILFgLmmlR8e0Z9ck5IKPb1GU5Vau/tC4QTsPAm
ZDcq6ForX3za2G1vva0KZfJN0m4pnBP0Ysbqh0MJtqZDOln6khRhpN/pbOScTITi
bOcAJPLbviEFpo+3GwTt2PxGXmKr2UFNG1NRXliJ1aUqJ+9wS8NCpcmhs1ZeJ9WW
HNNpuHuaBti6KoBGJh7apawcbgxW7IcKUIDkH8csASCgX4rHE0py5XRSXWdVR1uk
EYugdrMjb/BwZ3HhG3yr0GP9oHqIxZXBc+wypluu2I2Hn69o4TATGS9P881mCFPa
FlS+3e1P1JkGWhwIJgJ3ik8Iqb+QUuqKQAttYcL3KyygPt8EtD3nBCksCw3T52p0
hXiuMfLQ42pR6GWQYOMnyXSPBWTTkMrLDNWq2okQ8FyycIScf5guGARdxCCnXon7
sBXdglJEDM7Qsjo9MPZ35uo9r5OjuyXX2I6IJ86kSDVxxhUcHi6lBofZFAmkXliH
syfCT0Daa/EEq3JAxY5SbQIOqHrcUNQ3pd8wM0A0agY7WXgRGUIJ5Y/qwiOV6dH6
pMjzzW/I9U8pZC/ziFiWcFc7Z6Q1aUbwvcSg3LeUcY24COVYQeAv8xrH7DvGF6KB
BUTWe6O+u8uzkRO2IfSMYNB0s/AOBHkKsOcVXhJoMuhZWY8pJ/gawRR7vEKpQtgH
80/QnNS9ajN+lNNGDpDgRXxnUSyXVQZj2s9oodOdx2D7NhVNf69CFC9+vckUiy7D
1EPqJbSjZ3rfLJ3vveFviN29C3UXQgdbNXtzBXG/8owP3mlV4sYJwW9RDD0AZXbG
2lLgtF6jiy1Iy1o2O6xnLnjK9InqQvl3JR7HldYgiVURlL//ISuLTI4aw1bbhG50
r86iXpIVwLn6qQVRK1eTLjxVpYPUh92ClYUJo8tTc2BSSiFSooHNHf79KEs3ctkS
h6EtXkUP2T9662q7ZeuUjKkF+8cH4nh9eQ1jgsLBdTPjwnlm35UNlbuBvrj+GECZ
K0AoPvQT/6o8SzoirQLKuHVub4eTAhZ9f47VPz9m+WKlR7sQnuVYlbjX8mfVKpPs
Kpt09/p4ERokSD/TJtkRiusCuTcpQXG7liOc7daTBMhsleD57XaxVxGQqbr14vXW
XdplaPQKizHBcNOQtd3ZUckWTpuhKadsNn42dbK5/Iey6ZwXvJcivToQCCPlBzN+
s0xw2iL9K3BNYnYCYc6cFG7zkZFH2GCni9Mt4LbIpSYlLc6YfoAgcEISx24bPul7
6nh6VxE2nLCBzmigzUNLwfG0Ed3Gf7b8MRL1RDov3087Ly0IBAy08nXbhOp180jY
9ZNv0rQlEY8VWD7qaSJT+P4JuCOE0g1Sg3KuzytPOLRnDv9YDhGvjVa4JnJUziVz
4kLeqlvqOl3W5XsOLqR3Z+L2GzeE4+JpQABf9kYI0nRAkCjvzlJrhY8I3tlmwVvB
lyO7tkl+rSFGbt+h9ryzDZF9/DQRsYihQ2lxzNaEpReFc/5I2pJUsEIZsEaVoXXU
ks/WvNOQzok5QpHfpvbl/Rd647dYL7eXuf8RPtXAjI5l8pTQbvJ9hdOlZcY9OM55
za/emeJze9jkAfQtnZXjpaE3HNF4/EH7quRx45wQXa3Peu5lSpzCsd/Uv0im0J1k
G9NBZGmMKXirxN8R80/gc9pZMErSpj3l4QUhzjxGpIyeiY1+wUGW6Ydp1331Af41
G0fnjV5HI/Utw9C/ys9Gr+dfb/cI6XC5spfQ9JeRoQI/Z/sY6aWX7PdReHdwZq1l
csTty3e8Tr6oXuzmIIfQ3Iy1cHkTLGbjY9IbKgTRwrrV84DL6kg0+c4eeZE++Xqc
NUrqI9qWS670mfmfagzD65mXqBeLp4tNrNnH76l12ofLJg/0ZPUhvHAeA7X1xYUZ
iRAm6q0FhSZv99UO+9dAPXYws4BiJqQUGuJI3tob3L9JMiGyW+dk/hSGtFBhlCWF
Wd02EBesuScbM7YoTDIqATAQ7GzXbhL0xDm4X2y1IHe+Zff10wR84MRKPI1EzwDt
p3q/MTm8qPwft3XrVTo79oviq36QOFQywZBhe+7VxSvP43o3JqZsf1smH6VehKtj
wPqJyhuaZDXbrz7FjdrsSettsupw3qsid4xEqURrTBNNCVeeV86AwPor7LAr1o5k
kRqFVhigZSDZ3CWOFy2J5N0/6kkiFIagosHaQmjfUOCpmVzqM2maZm6s4sA8vttO
Wd5iA/rLDoSRbMibivMqkwai40ZqxUULK7dYWkIkFKgO6ihEvhTeWxKuNDM+OyCo
U+dhzbMOjwdmJGzTduW8D8QW88MeU2i8JWc4bWlCrVfF4m9w0zxRKzt43XBPnYH9
9iwaJ+joolY3IUQJXbCG8Cxyl0KM7RArbGX0qws0VX4PuShQ+eYtmDoiFn8BCziO
XPpgUr8sXwDshw0mZ7lqV9+f+odnUgjGf8BY2dmX2UmAW3+Nj9KyrCo/DsIpHR0n
hGBegUkxrsIkEtmu0L4RxobViWsFO6+NGhorBmYSwbP37eUqR8HWtw16uZkPcK1M
F/FHyIrfvep7gsK4tQmaZPP8h7JPxkJj8dASd0EHqxm+Emgjefz3Ixpdk2awxLlh
/y2CXg7hY7wIav20fNg5EckG8kaNh15cPwUY9Ln+PUK6NWRxTfNi2McU6MTYmEzx
xQevbXhP1m+YIpL6EnjUWAPWSlYVsgHxWhCQu2hxUaVxAOd7dp6MtbeDUc1egOig
AGfFSDcoPBUhIgkuXu9Xx9yq205I9/FpsMc+7bDex19ZXRUQNzVuSsrSt0MvE+WK
L+/TY8+oiydZr4N9byaHMDQC5Tu3LKSUxajiiXN2hfLCPPn1oyOUq+sb61uoZN4N
vdU7wLU5mvompLBQY2136dFXZeZjEwuRNO46LTaL+G14c9L3xp7FzVA0iKP7QeCX
AgcqSUHAM0hl9RREGJZ4v9a6WmRmXy4X2BxBtFYVxHkILRv2KBp0QqBj8mnMCOqR
Yw/9tkNRm/uf3JurZqEZbMIzIoJEfISYR2h6OjhY5JtKE6G+xWte6brwjhxdxfAY
jfkWp/yLUu2L3tL6Iukg9fe9+4Y8ni1D2F/aO9lauq7HhF23RC6V1ECXHKQPsk43
A7x2W+fz5NCHDvmKoBRtDBX3fkYtjdGBL8nVvIdGvzr8SoY+I6r6Y4QTJGXr0pKx
wy6+cUiIaaKXLxKvLRjy83eIo5LMosnoVZoeziOufJg7uHpfrrGcs0pg07yBT8U4
3K+ehHWMVJ/Ugn6Ko9BmydZViSGj9UdNF2JEw8m8g6NwwcA1yLduf2yb/A7VyVkk
PtSNsYV9STJSaaQHJ/DyOoPbGiqHvET/23ddGm4NzUa7bKQm2Y3u7HST3qoG1m4R
gAkm9CuEmZyKJd2hUJMAOGxUqSbe5IXuSVRUe3cODB8OEf+iEeHl5KcIyXg+QT9L
0aFs5A5NqaKINF+JPJm7S5fAtVvRXRKApVsrvj3EYv52rFko2dpLJOhGwdHm8B48
Cx0Dvr292SVTju9BqA1e5NtOpughQG5wj+34umUpmi2PQu90xysno6/ri/X0HVqz
Sd1Tyyl1hG0/33nmh4+pExR5VSYcv7Bkq01AhNkGIRTy418kLpCKoNZPZk5ekQzS
gl0tcOraDQp+poVIDOzGwK6Ji86z3p7ZFj5dBmqAiSTW28ZxfcEWM7Vk4ExQjpAJ
zvOKdLroJJULGeiDUULyre5Pi8EnvD0lTcE6CmwSWQO0x9lzaWE50zO1vHN3sKG5
LhoCFERDJAXdAqCSyrzyRk4ikO/r8fqyir4skb0a3pGAMxSNf7qpaXFrqvaBKSTA
r452OFN6jXKU3sKE2fDQO9Ue91Fo29OnUKSTTj6VnUECZTAwjy1bM7YppyM253aV
I8ciWXNS48urPfRW+XCmAtS3aK+CPerKOs22QKNgRaVObvzPP4L4gO39tFAWN6va
r8J1Af8Sn5AJ4VaeR+OWKlicWcwWfX9qEabrWx9hIx+ScRPW6fWeMAghFrt8qFm8
sOUdhv43pXcv9BLl0XWZdZO8KpZpRKIWkUKkAcZFJDEmdgdbKT5XVfTsbBoehYfQ
7xNVg3HC2XWyyCoSElCsx+G2rH9/848ssJ4WhlKOP/GXgpNQqrXcv3Hac7b+ZP8D
NRH8wTyrzf7Yy5kGVQP1M4hDC4r0C6JijSPjJ/o8Llde5x77Ow+95TXiemfRQ+Lv
N7KYWcOMp4Cl3H3mjfFUXwiBJXYc6rKN+WeNIc1YKCrJXvknW+ydpyWqk4sJ7LvK
9xzNolZKJU5UXfLX45vl9MLqpls7n1kpjswOrYGN8DG37g00O5t4nw2y2i59MNpX
WGJb3/VL9ZTfjuxrufjmyboOfrPLmDc6bxMDlCY1N1XZbzywjI+Vmh3ryjmBNR3J
MXEj5WRPjxSwaUsKRi9IkFBh5MKaZ4JQvYX7rX00s6TT7mnzpIHJz7FRw3fxlInb
5w7l7bTWpykfTDmJOqPA06dRb9IetN8C0DY+ge/L/cgKsdIPmo7Rnv9oQKT3hgKU
RGPoG2ev9GFZvhQyD6Qb/HGOy8ROXp0TRXZPI73e9qEusZoPPvvO0o48xGvkHb7S
G5S+QaSw2AIYkW79aOqupSVFKG17GHhtjmpU0g2OXFmcl34V5jqFWDgW6d6V9sMY
kKbGcrrAp0LtWBgkkhDot0lAJe6envfw1MzMEzh/dyv4Zp47mKyumEz4CYGFWxz+
n6JQTIV4by2m709KeWpwfC1Zdu7az4uV8OhjVww9MK1bfi+nbo+WEU4n4pgNsRF+
AcTrzoA4p52jVY7OcfnQVRukbC/Y+NflGACPKuLUh9kg1O4zehUobMEj3QY1UtpA
H6BCrITRwkSOiboi/hjVXHtb1uFwmVdutbFWW5AyBouIKajshhiePvh8X3Er0AqO
kfSgx6UBzbnLcBr2ELn4Rphc4OTa26ebyNkoAop00Fj9fN//2EmSSlUEk6RV7GO4
raB2LSV/K02NIMSP1s8Q/P8zdRvoAq7pYvBAGnp+mWXYoGJjUngXCzz5UqzEj7WM
XJ0w50E/gXzZOS0yD88HPzq5tdfTCuRrvUnXaJ4qffWA4rypLx0GW6YIKI6Zy+hO
g23BAIwt8BcptioCBGchOOd2WUUsAvTxTfVP1IrHL4Mo0c0c+1qooQdpNlA+28Jn
8nM3aJEhwll7pl2rbKqSMU2Kqbw8eXMYWf8dFI2o6wPuw3k/ksxBRv9L/pHQt2Qh
kwGAlSykAS0MkrcWQvmy0kuJOyjcR+S5h3aX7LXCv6qgRxDUiUvUq0Awe6DJQtHB
YXsrUnE6Ow+Uhb9AOHnuUNrkw85s/MpmyS196jeqGSywCgfVKydWbJnCvtRD66lD
PLoRaW8m/gFj56gcKxcIcXRpsZ/QrV0aV623v70XvEl2KzKfSq/whTR1nPcz2daT
wd8XvQpJ0Q2c9TmSs/0VX06ljtvtbGZmhiSTlZQHg1PqJ9qRfWhncA/2CM7y/CDo
CqXP+hLQ9+J/aW1UQLOff09BrdOIbdwbiibOpEyrojzOGSbVa9Qj6ZExNmAWYnOg
O6L/0YtvmJh3/X36PzCooTa5VGFkZKNJpTIcR1h4UziQwL16jpGwDMkNCoBYcdbh
JZKa70rvFiL0OniyQOYNWGmXdxbAQoZz83MNEg5pEDjpb2xS/+TE2sfEbN6UKIsg
KkAZu4QDorucpebSKoPRDk4UxM4FeTXUx+eIOlPxZu1JYi/MvRKJR3TeuyhffBSF
uKLeiF0JnrJqqvoIAj8ZrbuNY552/8C8eiltVOZvSFJXPAd+kOlgj3bzr4QqahzK
eGpK9VHHhiuATi9AfVFBP7TtW/lQQ7155AmZ3vfr6rCjz3V6uIFHMQpJC+jFTt5J
OxcEDzY6iIrQsUlKr2CtO1v6G6g8XlR3jk+Ta2A5KL+AJz1E4JqJtUvJs/aXiN2m
Nzd65+joU/j0rNQ0dH6XnLLE17V534O4SZmXHDzor9upL+W8Hs6y4BgcZ89XSw0R
4U+MTp5GGSLzA9ScRnENKzCyv5jGVB+l+AVRQFHpss5/MvMqAJvY5pzxvWChKHve
+vprfVdJjdmzb3WH7xK/K4HRJfmp1vhJrYLbFj784p7+JaDWYiGn+B7kbUsaJwlX
XGlw6D+yFQyJ4KbjI1tie7+kxwuNv4Jt6niZwN0DJBHDtCo1wx9+QWlKuIkfAy+e
VxoYH/oiXRK4yEGk60pK/c/bkkFdSNtKPNZGheegarPGiYmB3ZZi8lgMkxfKO30W
jaXOUOl/u6a/JHrhVdEMqK9n2g3+lVUBbS2Z0hkcVJkS68BtIEKbqZADEjYGNYdR
BzKQZnx4IzYb8oIPGX19B9HFgyI2Y54qBUmDLGG/zkgrtRGPiZ2Kf6RPJszyCIs0
/oAN8fAhoZnR03xq07RHXQBJ99BmyiXEAORubSNfkcjRjWhLSk9y57y1LG8fwLiy
PRlIiDRnfglDzcvS6/nRFSlJ5AxpWRmc2P9xoMt2QSvPvv41slfVTsdqHfG62TEC
tAgSjAeOhtv57Vv7ryW1ZSPjY14/IfT3eKq1LeGhqVW8KV16Giu6HzvRt7zeSZn4
olqWiV9nhsNXf1Cle/kfZvJ5riczE/LQlL/t0f2Bv8VM7XT44H2iZ7z8MTnNe229
1xgxBC/QTmcT5j3erx6FN+2nCsYUP1jIHlqHUjgox+K8Fi6E8+UWPZWmmHzq9iID
eyhSw+/QpwM3+sLhvc+ozaEoTOpi/6A6WkRLTDZmLJTYmgBVpAqS91hYsdLctbYJ
1N2Yqel/sgLDFJM6pV1DJdMfkmoB/OUT/llZIk2psOdduxZmQsXuIXIoMsADkSB9
ueqNDLFqESD3bLc16xdFwvvXLeGXkMoJlkDlF01A44k9EHBtOSQKWatc5NN9OtHl
iZ7bmuZW1i5ra9AiglYCAoRPbDUZFCwWO/w/EM6Kvkyqa00ElfrJs5ZFc+VrirwX
2wgaJrld32VQ5ygDozTib1wjG8M1YPASf5y8jPEZA7nfyQBTOVXIdAi7cRrbWyJc
RcW44yGt3LhmftQW+diNNSmsQvxpYqAVL4P1FxLBhdSsLf7SBnnuWyeU5NNAxdsA
RGxULr9Yv36GK7Zzaa3vjwgoftTBqdejsLQm+bb2gH2L6sh8ObcZ0sSDIu8N9joE
pnFMYjEFoU/6Rzu7wqtKXabrgenm0Z5fofpJHz+FXnI7A5p/VBcvi5dSuPfI/GdM
M86Rr+Et4UDgue9RIoBxph2o3empqpMAjisgDAAKya937/RVxzbkSUDtvyJdhIHz
XzE7zh2NEnjkN5z0a7vy+zu4p/qCcKvneQ+ts4ZyjtrSiq1qF0d/kwFV3uNruuXJ
JTjL4Kyp5f/WmtJOOh7fyizKvxtn/mLI5EMWbFFa7EC6norhIE3dD5WFZjWXUO8F
AkGf+fhyY7lWH7w2M8C6lOn+njpRRHF5ivER/CcVeIgTgryiskeNbBdEAFbHbc4C
znMiVR1Y7iD4L9pMaZ5akpVWI0IYbWGcoGpXRZySBsd8Tt48ycAx8eL5OwjxkRXR
TGY3CEgOwjBG9Z9V7HFMiEVu5i8/Vsv9pNB9TRMfceFc6eV2jogoWqkwwBiCwUAd
g261kqSANmAF3BAGer+usJWUkUcXCOqV8D6ktDg4I+ZVAHMFDcJ1krOdJKq6JA0x
Jrt8cF+JnkEPQ+7dUFhVGpHFeeRgFmdcwALCd9ag84pmTtuL4CwoPYjvpWsIfVzY
u5LwY1x35yyKypWDwvOvITWjwgnLdNwcSTJHW5yC7mSDYAIEeyH4iivcd+AutnQ6
+uSRl89q29M/cpzUsoBsu+GckIOaWjDcJH7cguRiAk+4bI97V3uXNvQXjdZO8rKP
g+0HEETEsw9mxZHWCTnksm67iFKbJy4vevlV2AwQCn0NZtOFf9y4vLNf8nolSUUd
vVKRKqpA9QT66BhPLFxFqlPwthwRto2B9BhGENmlFPJf2vl0Aqpq7CrGehVAq2w9
lB5RVM957T61s1qG4pv8Tiw6vXdx/gZAJieL2Ce+sO7nYDRYDGDabkA//EusupEn
LXgY9I2hhaWpQeOteW250x6KCw9PSvA68+ijEWa6x1uHCHmUV2kkuSerMfdwBLeD
9AzDCDyI7wllPl21CKwBZW7nI/IEcXav9yEg65Xml+YHuQ1rNhkcna8tW8YWqmu2
crC9hF9Fo0gdvFE1w61LNiRpvOlkfyeieOoyVISsCISzSuFWRnKtnwJKFkIAsGVS
ID16RpjmUMOZPHajPjUm4zTYtBFE2xsapAOIEm9meE5eB5TEJyYV8U+1jqKbFXiN
m9wUhloGuxbuKKRNfYVirdc4fCEbTHuHOXreT7ZmxJjfGGLtVgNFUE+MTlTQVOWQ
oy6xVhhqfKC0Hp2F6Fo6Xp+OX5EtTrll1l2m+dyZldOnB/n/NBpUcD+jNRJn4Z8x
U9vgm5Jg4ElTuYHs2P2KmMzK74Cf7zHdBdgqq2RYo4Ge8aDOeaF3PFoe6aZhbgHt
dPgpR32AJV9LaeBlRRXguhPhh6PFxvi5hrqVmrktuZCcwDV4SGgo/opGrWRt2Fel
af8X1HTaZQO+mNN6kVei5UpYzSweEhyF1eNIW/S0HobojujpUQp75P9U0svaV+/O
lvusJj64sKMrOKQsOTgqwV0DbHS/ZdxNavP4aKncnIaYQ6aXq561iRI+E5jFGu1H
xNsOI+5GaUclaNMO/76abDIg4jTKB5aqPb6PmZWHTHgbjOv0NX/TuNpkUwQKK9Ig
qu9K7yOneKdXGEZBybEmb7fw2wOHaeaODi5xg11NqRnXNUBooZgpBWrb3cNeRhJk
QCzwu+rimM4ek2kVRCGNbyZug7bmc4oY171W1cJeVzA1Si06gXzHZIcRA2SCVvRF
hiDYbGTEBTcByfB03hpPlucLmzm3HmbGSQNJ0/45jMTiqqJqtfAMQ5nNQDQdTuA6
WkH64UW/K8EwoZRE5zvyYHoJFVAWrL8g7SaXfukt80yTHocbj5hbVqOyweuyyoQ2
FUTS3UPAH3DkG7yimW7t6zxmOUi4Q3YPLocy/mjSyrUy25pXGYjxGMiDzFNG9gIj
sC8mKH6V1e+iqOQ/s4YCTW9iAwNRAEj7G0khdgRbAvdsbRQisyHSvyv1wTDdvrTM
TXeNDHO1I5lcCi8k/MhSgjca0YiTmEM9vgx3XUUQpz8ft4uJQYzm5cDJsbta0jdF
0yM0oVe/WTf8wnblokg4/u1tZmOFS6meI4BEbfBSjZ56RHLtlAkvoq4uw+NGEnUB
LzWEyCge5pJDsu962N2yV0KFS53nFKe8REpyjo0Cr5EIJSAsvJiYFmQNxhwtbfSo
EoyRa8CC9w5Lo7Woy45yDfBYdcEZW7oiqzo0NkeV9w60z8HOXxBqK20t18Savgto
7cfZcPU65mBPd04sLiaMv9qH9Hrmsm9MCJp/7GRD+8SK/MFkkz9gvMrRHTMlQBiE
WoYugPib9qWqAsXzSTFvFMvEUaB8oYe050pfQsUUgov3Ad2Kfqn7sD31VjV1aVyr
y+uohIRPBnNxhQNu4Ui+jlhGatC8FrGLV9wM2FbuBIU78KOKAuJfvHPDqIEHu2lb
v+apnBhXyxxdYcE7i6x5fHohPolPnyo3lU7WkqsFhfQqmp/A0qvfz6FamGdFJkz4
czyZCxVM1pGdmXo1CsL4LKZeBnSHuD7OOAfO+442G0WrFhXzoiR1IedkPNjyTG5F
jYetQsSoawbs59S9fGk3+hvU3o7owUfTuE9tRWSlSN1wIf7CWjOxrjZWOZAq7xkK
E2UDKndzYVHK54+XBjO9vg6VmwnSWF20s87mmNmTf1CFBo77yFNx1GR8zja5QqQU
NmNbT/KgxNl073b/BdpxQmrTmf8bCxY1eXUOvFQggXnnT2zxR/1ZralBaHSSs6ZE
Hd7Vrd5ghCeFy3/Kmf6O5a2wczpzP+vIsCwzrdkHxBL/eOODj/8RyZF0V4J6fTxg
6miiwkbmCIZE6hwyJikfhM6aBneTFPOD1BrDUQntH/adLjMIPdWo4YH8hMA2iLkK
0GrCIRtJZ+GvnWHo678J1snFQnFS5R3Esi5t2MmK9BG+W165+l5g7UPuAUQjHnKx
yY9pvxQKmde+aCMKYDpIgk/f5SfwWlZV21zcTqjs8xfVHbrDCvEsrMv6VN2257N/
jfstV8pmbXnBE0vJaGNCDj3yogJXooQ4aa0gFwKV9A7zoT59GFUxhtEVmZPLtZ48
HiO5aByjt45Gnp5a++w8S1adg3vQXEX2UGHoHHnYlEX6bFi1ilLdYThUDQIvYHRF
7ktjeijZ9ItqqTQ3SK7JuXjJd3TEoghh8qSDTYZ+GHvxIf4yDeP/RasIMkReNPwh
cMPR5r98MvEZHMkdmQQwKVLkIq2JDBDz2MtXE7BsCrtfKnwRL31vnsM00IyOt4qN
6l6fn2Bpf4UKot6QuU5mPgi4qgpsnxdIL2UQuPQbDjCVxeKf63E7OrDtmnkktQ80
sb883RsjLShmqiNR7/nhH9mTnXUbI+2tLrjc72DTCOC1Cq5BylSGf4sDbA4RYB7S
nuH6HyZYoNGkevDqdFOUuOmGSK7V5MQrooY0PX3QFDs/J2kik/c/XzK6bXZc8dC2
gfeWevda/IXA9dKDPRc82CKDhIGOoTTCc7B3h3OF1F6h2qYVG3J3Sak5qx4Lx2/1
9HzPHPzGGZzX+fmj7u2KK7je+1myfYadTjPWJrMm8nqdLBEKB0Jf8Bwt1V0Tg0XM
5rImQL8Pt2JnkfJEYPxf+I94Kwt8VA9rpm0MArff3K3OqM/SSs9Wy8o7hQg1q1iq
I9yG0zBX6bLojHaMC/CKD3zVM71Qu0GyX4XbXOnvTq3I4eaj4TN/FQ0QlII9sjB+
mgVprHndxTXcupu0LvNLaLeY3/KDnjqZpsI+d0AM0GrkJdFUr3XS/E3p0AC9lr6i
uFK2paDQRx0CZgkTAEYgAiLMRBPbKq1xQTE3ZytBqVrTtpgIMmfRBqf+uSfdfpro
CHAprXNFOurpePhEPk9o6K2tP79HSNCsFFy66UmQ/MWB+hmF8AZFk4AQMt/CWX4P
sbZC9CnW6ut1lDtYaix35DpuNoHvA9uEkzZrobUFb895EeWmpCf9cstW1Grry9Ng
BGP1G+OppUUIW9lgbd4uH9bCVhT9BLfLLbJKdPrIuqPRK6YGl5q32K4YTtY7P2xi
L3Kq347G+VjXAckAmS+2MWiswmJpPdzzRcISHv28sJ5yBVzLIBxg7pIXbyFp2G9f
MzJA5hysNYP4MUY80kFlcDIIekURcPrQ6XfYw11t9cv/rh586Rjd7qQCtMBf/VEX
LyB8BAgVhFtEF3mkPMLpirrH/y1zuii9EJMI/mC0UPdzssZ9dGMLYhUMel2A1xHT
ElaLeGbblEIxOOajE4USJsSmhJ3mFjIKRCvC9YaYenGAC5hg9bTYX15OZ1e3bDGO
63cWHqeA8XOStzymPXKmAdaG6wxCpiHy6A8GQkHcoASDijLFLxXujdU2ROGx/SM8
GCxmJdXrstG7FMInvPHoD9mA4ShvGoHToFyolzHjcjxdbSHtCUYtWwq2E1B17eOi
fxdeqK1VOR3qlcfx4EGLnMtVt9SEybm+zYv2wThyoWV2GQxjAr8Zk/A5qKpZ2WLw
eSQ5LOZQEVG1wh0HjNRdJ0jZfS3B/gXV9EXQsm+Ed7qgVYqJUou8mSIx7+Xm6J3W
YFQ5PJv1B5HdxTZJ6kUKG4SYcIWlpW7iGTVyTFtkZ8FOWlzYKu4YwdawM4C5xX4G
S/4TbsNSPqvt85yYcR1Oc9qccl3Ornml5VuZPEXqUr/hSLgfNvxwi7sWE2VxEmQn
CJh9tXfK1HgTWwuvlpY3m+EfHLrmI6ho9QHZ+uQsIuX+hfl76gEqDUcnORZbtCY6
vZ3M/zJSM0gVHlNnLpo0N8sDd6jiDhqHxjtJhZ4Ih/fGAn5XDmhey615bBHGW2fh
Lht1B+t05zPtqmWvSyx1Scq1VRChHNoATEefKKgJz5YfmBtvHiVRc2nAzNkvo1P/
K/mYJS8H2VFV6Q3X2qnro2ir5qZUohodxGimvfFb7CumfLupDtX3drgLu5kQxg8s
K8VwsYznnMoi8ZaCK/rVax1f4ppsypGKZ0uIhESpBD3j4dV5XfaFsnslN4yQFqsr
8NQmajVhB9HtBFb4k3+6uuGtuMyDEw9B7fvEtuI4hm8YtGdjR00EEU4UyZX8usmD
tgD2MgaU242HL5BqHdkTZ0x7BKZos27/S1RnzMP/6Q5teGSYITZoLqJLWNLnr85b
KOdhHSf8CwawXZ3z1pG34RcDdpVZZSsy3WaLDmkLXPRj7FHMvESJ/M1awvr/0EGP
S/mP8YXrd6hBVHMmFkaiPRY5t+KmwQP9SHnB04d/D93azUzY3FktmAHJTP/WV20H
71BvWe3wOvKcmyHfomrTH+YBVAioKzt3llvDx0z56Dt7ET4kwp6WBBaodtfJfZfU
Q04QFDPiugiNZ2U+BDhmmYL88qzit9BMNwN/+7QtYRA0wQenLxQPAOYG7skEkZ2j
PbPUwa/aEvjA/N2817HKEqee7AONqlEgA4xV3iQpJQxj6zNoFuG/uBQpOAobH9hA
taGvFzp95sZ/jekDSjuXTMpYtvHcw5B/+3TH1CWSN/BQSKIF8rgELIClVmaMF+Cz
nkNe6CDbx2RaNIW7w8vcrUk6NTrk7BzbbPgEUQujdRGXAvAb253+lwR4aXciQZDb
hgRI9ATWXd0SdfIbZUysM3m2sPAYOVxc/Vd8RZzsauppHIrrMLaa5kFbqYhWaCY6
2RjiqpsO00+YDMgOBOzmr7rBj1/XtDYPME1o8GMA1/PztA/9YXo6B6PwFxWJJaHQ
wNeHbJlkAIH29rPNoUY0vp/mS175Y+pS83lj1cvYEzvzs3jd2OInL7UlE0aSF4rG
pVFKXWlnWTeTjlTf1PhcG9qzBVQrBfXkygmuGvZw0NODcDlALyOW1s6rv/Y1uIiR
mVbN27+IWFNcmTHUJxfFEBBxguCLTtLWWF6R2lYPkg5B+0TI61nJPiqFKIMVaa7Q
bgpGroqcKP3DZt+9lqozj/4l25Z9aSvQ2stl9Xg7ow3GsA5folzXML+OiwUOxmry
Lv7A+tF3R+pXbseBzaEdRYcgPJHEHREVSSajLzlHQEKga1N5q7C2JEp+uRjYaNpb
Ptr6b0527bU59yCFZAaf+OF+eQDs/cwp/5NgAGsrtOOAIVGzZeJvKmZYsgPk20uP
qagNJFWPvIHzDXU9jOPNUsQTu6yHrG4T71X4CYOJ+lM/AwSwExiLJpXEvzyEXwKq
xXJGvOp0f7RoCLZc07v0YtNlZztO+fB8e7ckj5EFKfeDmanmauCB8breNzt3FaP8
gS2/lDOLpDpQWquCE51WacV2eKHb9cQU1VzfiC8bVJfjSxcZTnwsV0z6/O1rWJTR
VCS3S335QRdQj0AluMXN7Uo5t6WhXnemte7WJ55kSpSomQPIH5FeE1mieMt3K3eY
0aol79G/Er7lsRe8ysuKLPj8AxhowUMX0azJcuCRrAyVsR9Q+YafDboJLqNze+M0
DPYf+NMX7OUDxkQEaIAUfiGEC0JnHXs7CNKseJ3mvPHaOY7XKGXWJOm9e0joOzMr
F8MEEYhPk3XQXhTWQOHgEdAT/TzxcytmLYbQIhR2dMVw7mfrnCf3U7LhYF9q2oo8
8OG8Bhd7GyGd6MqhbL7WOuM6ihpDrBeZsWBw/ytBHnWDPEccBRMxTteGGzPX/mDd
e+KL0A/lsz2vFg/P2e/g89nlLdFQGB7J07zTqj32I28UKhy9dJteE8+rO9oQB8er
C/aAT3tQye5EolR6NQ5pVecTNVBBROccUdAHQmYQIyS41UNkNtmtXgv9nqceDUVJ
zp+a/cDOx2DmJQeC5NA6pp4XbqzZ6v32dOE6mzc+9+fG3iw0p4p3MyoAbMS2mG4x
pt4s8vUnAlHC3NOHSq4f1zrtnqA4MCbIi/trgabyR8ISCgRYVfsoUr93oTNB/oAx
ktaBRUYKPu0ORgk0wgMIZKurL7I27S7UfW6dKNLDLaHFLfCh5nUy4v0ICw+g34lZ
cg7ZIhBY+rwoD6MOnPKfDi8Z6jbqE9EBs8/yrpFkT6WKY8WeZ0gm/b0ZNGDom4if
TfcReeKsM06WggwgmDYZtO4wyU6L5JNIjKu3DHokvclvQ8aR3Kzgiq1sU9IU1Lfe
rcrw/8rkwxLim+kqE7cXuBd+XXyLBTyBtw+L5ntiyhQjpkb8ykwpNVsRXvbOqTYg
uAt7lewR6dJzWoEt5RGKIx//+HsDMgbGsFHZCbeEjDnqnV5kbz1hWaBOJLSTX6zl
ch0GYVAO2UpubaaEOGv5YG57JkDYLfeLoYbNSZO26reTFSzyHniHaSgUMNJLf2Vn
bROJENqD0SoNoomBJLcVehVIVmcQvKLxpvI4qrK+yFn++r+dr2DfZq05js9r7vOy
xURP4T9x7TRGd9AEmc0kcs7cS8NxfyNqn+vvRn/rtblH+xV9X0zaDjbVKocFKWlV
B35Qr63rbJCVthW+JIA64g2cDYQCG0Fv54Jy8WCpGCQsuMri2c0V4Ap8MfApiGrm
znG2Z3IiYVX7MMBXncaVBfkfJGGN6lYJtMaDN+MDFAUVBKxYNYUq3e/TGymmsVmA
+v4ZwrfLNEBHVi7Ga6pd43McuKuilG22nDzMmwuOnB68hyh/ywl/VzGVZi0MK2CC
jEZ4qOE7PmKDseMi7acQTfXvxa2GZhpi9pf3ElDMnzAb3mu6WGH2vnybVCuMpfHJ
DueZmhtrGRDe5hL4Ew9jlcfH/MAc/4nukI6T4sngYVQVzHy+gtkjS7CJGhwlrsu3
jpA3Fh3PNssFELxrQHQN/Cj5SGPsxLmtXiQvzuChxa1N87l6q2OD3YtglXRSGnQU
D71uA70li94XIVGzc1ty8+Hdxd0TP2s9Epx5MEGGhf/rFNq9rTRxvqbJ+jzCCda+
pkqwBmhEpp2pxYGhHHP91XSPUrHfkcvMq+EOuMwvi/kUvXNHeowafIXMnVl9dMvI
bmx3cirr4X6ZkmQdLFBAMZT+eWepfs1NUm9cAxpwemxGa3X1ve+dCO2NJ2UyFbY+
ufYAURwy5rVvK+KPbrRUN0ymBec1t2icVdOZwAdW0uxHAnKlADDm1Ii+sPSeDlju
PLPBsgvtwqa9u153iJh2ssIRZ+9mnPgkWe5rFNObgncDHuCDHsbjG2TVwW7KN/SU
AN2Fep7SiOlTjEI45bE3RK2/fehtxIVAVAoI7zmfvQr7ZnlN3bGy45dHvUHamoKf
js1ZFO7kRgDgq/G/1FZZuVahSTqpo32/2OCbk/nX5m/yqbu+dEVmxn8hh04YOq5A
ahi8+f38tOQR7p6kvnPj65MZ0ZpERQWPwgS2m9UyFF23ukY8ra91kpfKEASBIiAj
Cx6G2wmoPiQs7nfWzS58/+PKByUFd6ax53EK3m++7jP9SpCW/tjCCTAEsYqs45zk
i2tIwci57lNPuOwRsT1Ol2Ij/aW1F4pDywXuPcD+VQrabpfNUjriKAdl2p3+dugB
gJhXbX+01vszHbgQpCDsX5LNjoURm0TLUlBtfPOuz118sii5CQvMJRpBsJ3PFzPv
zRUjoflby4y/D3pxGDbVENsJ8kBZMK4bTq/oXr1dNqT3H92WvvUltXYP0mRfkpDh
sYOtd+8JB2HOReu+EJdO7yvch8MwMC4GxG/b+xKVKUuZW8UODZRR/QNGpEBzJVhp
SqTPKiZN/7/VLPmRNmUoPjogivZcD+hjIno4LCKiuGGix26s7S6a005o71cFHD1Z
B/9zFRv5b4OOAEG6w2Q2aDVRQd5XwCCBWiMEWC5r39G0futhmCD87je3DyThFknU
5I7sp5LQl69uwezZ8tilonP72J37s8oiQ0CO5mbL1fztEXMm/SkodLZkEEoeQe2V
Hoijok2RK2m1XvH03b/k9nt9ziwGHywDP9B8tX/GoMqF8Xw2nR4rvuD8HkbzLTHd
DLDoH6btzzdpTWdD18pjXdRScSVfyBeJ0Q4oIsVTb7ZzpqAYemXnnTI2KlKe38bO
ge4bAubLXFBpFdeQPWOI+xv9FQDRABZLE3QeBydhRUbxEemtValsbeoWwmPqJ6vS
91Hg4N4J48oGblGJC01QN/aTfqrgkVjBh3B5wy/yCn6OwXFyoPxfAZGBPGgb2A+p
RewQVmHgvBsTikkc3JqHQSdbU+lDL9GBMeMOtNXpk1cHdRtEOSbGLNe8Qbz+3Sqn
86DwTktS/jVZfp2SM9e6GWt+gpnz1mnvmOleNO3/clrKn8PzeWN99TP0CTmedDBr
WmlNPRiPOwF277kdG5mzH7WTrCbOqJts5TVDS66sc7WK0slDRgGRx91UWwdn+RJp
RS9p9P1bs6YiwQTBq60WRlHy7Ww963SpRTVx6BAjPvW3bvAXOw0lcBv4QctRpaB6
NVm9aKJ7GfxIvwmjf0PXj61FDX2JlqgOB9laLhWsY476SCuH0NboUIrGxcpqj2l8
lCrNNjR6A0HikbIdXl3vq5W0nZG7DfhJ4JKGAvwNzgvO5rdirGoqDNugy9mqfFGd
4bZGR0F1/j2TJSRZnt1/Y8M/iSk8yXsbqo/EdH7YEvmPKnusNwFVyDNKZeqGM0Zd
CDzqwRGkf3JuvBnUCTHMZEAbOdDqmLFIC+w7icd1kVW0TeO+/66tJLFg7/KA71bL
pCxptxwisWURmSCtuzDG1c3TyRX7jEjF03OQH+Il3gIkEnCEnRm4BVlITSAHffdg
GhgIFo8Ba7tvgGHEAcoYi8lSaah2cdpV1fuQcbX/j4BPJrweVcKcTtZMx6iwwglh
9YrYCpGU6snaB6ZNBf0L5uf/QPJVHL+9Ko+lR/aI/B7qz0jwcU0kt4JK97ud/6Eg
7AtA+btSuETU6RVV6/j5lOlmitbvrYItpggqe+MMCxXWppwaq+URlDaLMXbY0EE0
kgfLhKddj+bmti4d/AIKAD6cF1l7bfRdy9JyLXICNQ06h5K+xgl53GLBcbQUJvZh
lSLuMInAvALw9T1QlODWQdntP4GefL2udgHPIjSsAWRxawWqY1a5jlAMvruZBEtB
KJritgvHX9Uf+Jq4Mg0ZhDCuYV8mu3YR06jz/njVL4uuzm+4mi2r4IGwrupj9WcS
qhx/ZvyKDtUnM1KXfGSo1IkOocX5Fe26aIzSatVEM5oq1xqkKpltChbWA+z2/pKT
yDueyu5OvFgTifsLm43Rp3p5gCCm8EJqrc87vYRMtoEFkLGUnJ4gkrIZbOKc79UC
QFNmT6ZzbTWaW8X1t0sxlQMrDQAz7TnEU5SytbWIkc6Rhd/Bs9sSiz9DiHBPuAO7
NEmtjsWWhmdAhqhwC2er3kq+YUGB4yrhJ4z9lavsrM6MpWMPcBISIqpbs8jSq78m
JY8jxnJ1z2gqomx5DIxdl3VbfxaDVMFv+9fKvdJHRCflCECxr/frqDYPIs3abFDS
4pioMtl4bFxJkQWZeVcsmw626GYNyfNxrE3CvlvFWWpoUtf01uvQKA3KIWBtz2cW
+sUoaRSb9ij9vX7pIyZCFUzVX2xbCvzRUpFGJNqYaPTjOKK6JdLAeg7OxSU7ZPdx
DYGKnryhzBLYtJmpd59jRcD95aJEqutVZ0OJfFUDlodrDLJmgxVEWYU7AnqmH3PW
As6ewm5wc52gx0cFZjOMK/yaDGth1n+scdSKh7I+FzPhrBbpeh8FY3TAH9Qckgdd
WulIID79tg9gVJc3KFRUrucx91xjiJw3KGSDZEQ82DFw0HWqKJAXvEPhAWysKq6a
JwFlDCheEuNQBTdikRe9xDbHIcKtLpuC9Db/g25fWHTT2zh+5Nw0mO1z9Va4GpI/
VmWNwWvwXx4QFAtOvM3/+MoWIHSfeeWJpq9TM90yUe8BTSgstqga7kNMTKJhRc98
ZULBrPtYNP8fuORvicN9I18FlyPyDaK1BBDNzipVbsrCWDKCl2AgxhtgBiYxXdga
T5rROLZjxSpe63zTO+rnJqIPqjVHwpWthPXNr8uGWop9fsYGOvXDTei/9qXXibbv
LbqjlYydVknd1LV1DwOFcmVmO+K/qo3dzflwLyB/Ulz5kcTyn8/H/1Bw6v7VHlNW
T60/hSIvO38Q5jmm+7i7WcV/WM8Jeg56BdO70JxnNpxV8dZLm5YzM0PZ1RiTFlAM
4T2BXZV7+GtBUskmXU1qFP04zFh258nrXbZPIxqJnFAkYKigkmgaPOaUqlu9lEkL
VzZK9P/ASsAqfj9ZWCo2XwXq4z0jw6HZXKpGFYfwuybILrZW7Q8EPTB2+54x8aoV
rNp2Lts9sXR4i3U4K1Xj5CwPQ+fsx3HZA27P9L7fuikKPOc+Jyt9hzyecvBHuI0c
3804N/65x1ncEnwYlat5tozTrNjulfBRWfQDHOTM7Kh0bivR4yqY5hFQWaSRyDCF
palGQCHAOMfBGbDBycFn0DdcTsLcMjvZHEzAmQCvIODPJja9HaK+LDTQe8gIUXWv
CvThT7/d+VR/Vztgp6iL6rAgWeqg0lrOTTvi4pPQcHCYTByQ78KdDffYaAs8qfTS
B7FTelff6+HgLlFo4sXzEcOFEYE10OeHcBtvc6lDlPu1EJNXYLNlIeTTnOA3hI8l
BreuoR+3PUqumOVLDu5xgVNR1rKwquBAAu9rTjM1IV89nDiLOMfNubhx9J/YgxI0
Z+ul3N/TZUMcCzLcGJNBRTaBZtgHm6uGCvaIAJfShE4MYHhvi4o4jgr+jbQaU6XS
lQuBw5QiFXu0f+fAl5+5+jH1shN3errsCLmUB5aliID6g3HtABdA0lPTShvOHcT+
/W+xgo9ei3GwXJXv2SQ5AuzhsB1YiZqAj7c8FbHZO9YPC3UHKfOUbaj0d3LAyVQl
KPFz5fz2PIbhqpdy6mk3pmwdCxshJL4TMxvFOmYz4bpyBMNpKYLwQCHAYqYCN4dc
iwQlzj9ktu/sTtdwIZjObgPK1KgudO3r1b2zt7wdvWy/gUnwKEHa8521qBReG+fx
04MN6J6MdMLM9isxmlgWW9DIau8sXJKA1spXfLkNSqtuu238mPC+X5z/94lKH51f
oJtoPGZFzpu8ASdA1Zippxhp7OYDIQ6P3QQWTNteNdRbADnL2iBbRuVNvTgYCdBU
27tLJzxC1mDoL2G0fUP1e36SX0IFQ8z4wlD+5O2bYx9kNdjEdqvYL4iagmNrStu7
X0Jj9sf2pHopxfX7XdA/fMu9dqwjFcTBu71KEFjnq7rEUjgQEdh/OwRsweao6rUy
wy0yjk0QWJukJoFcnqpRwTGHbRCCotEX38VHCYrexP3D8U2zhNCGYhzdqssdsCNL
qkFPQ/7HbBtId9WZRtOKK7HYl0sJzZVEHNWd+7FdwxJST/9LIEc0jWUurXBxJBQ0
oBie1TL975LKfs531xaNG/wkpgHXASPYT1cB9qePka5flmtwBJ0iA2taNAxY0CnE
KlELatnulTwLkdhiZVQUqSPmXYBdyTik3FmYO3xcA7vPtXaIy4EFtKguJQVft22R
1bM10/pxsVYihMu1SQSSem6D2Rm83ca6nfk8p9TXNPpqC+JZBY9ZuvM6oeajp3L/
CHNse13Tz+I2YT7Vegxc2e7S/Qf7sV4oEz/z1MuXrPULqWQghtqMCxKAIF/2AECO
jz/8eAGl6VtaJATDtrSxIv9s/t5VwZsdVxeZNZMR2ctYBDMCP/3rv95fL3HWF9VB
w5eRMtiYnEv8KXahAvJ291hjv6oxuf9hLE2IhDaPKMdUokyTqD7WYv/cWoL8qUWs
QOG1mRUV5CT9dfBKynhiiTagvx4jlkysKQjNJ97B6Z3tYdM3azzRxH6NlGBMyz+7
JUln3rbT2lzuUTz824hNHvOx9wikiO9+7d9m4nL/XwX9JZExYYs5cH2xXBnjxD48
YhHeLfHJIbAXTPlQX9vEwxpDTSC0U8+xk+Ng3yGhiumZRwXBMake1fAw8TOiYcH+
gEgHEGiWrpuiz6GTQcZhzB/Jdm4wX1/UIANlpTsgALr4C6iR4MORM2uwAbJ079pb
z8EI6tVY3zzlxm1QmkDvqAzssj4Igx+6DBslS7XIc93GVoRMNaLoxlQNQNW6Mo/k
f3Q1hTYzcyX7gesU0yQz/IKuVlUCJvdTAVLhHOnjCOTdaPrt9oVSPJrtSIqa3Hdk
aGF2azku4bCLm8/ZtkxMFA8fDv6iduXg/S45H8FI5YSQghuWIFvfQUhIpsfYTeUl
/z7+QxHq48pP44aryqkpOce1lJD9rpJqxFtt2G0PUnj8LI1kDaj0MvByipLSuZtU
oog346VmeK0pJfwQOoHfjdvYECS6Y0wKd/TXhQDcorQZXt16ZLP9iqHbkAR26g32
D1gwBgHfLR7Pj1lLdlr2oMhXVsa6lkBbuj2LUYm0fMAo3P+PrwXa5Mq1zxYbBPv5
wWrgzgfoy9QrG3lA1+awD53BZcv/9qNcgzB2NefWjAzY8GCwcNHMql4Jzd8tJXzJ
EhdPbrrj+bFTkYEc7oOqS+pJQhpPAsxlB7g5cdkOerXSv+MczKrgfVVi4EZYT2xN
6/lHcdCa0aPlH3r2jjYQvP1c4AJY17dmOBqNZzGT3rHswhJ4rXEHN/JNSj49c1X+
m4FjbZc0/RjO9rs3K3S6dZvmGWVUpwXMIQYKmNGOEcXA3NJPlzxOVjl0Tcv2WGIF
VoKE+098SPQT2X2DjGqHUBN9vybzYngICV6yEIKr8lFHzXYm+pKjabU2vnpwZBl+
LpiHOvVxA00j0+Jioz/+V3pOqMRUYzE26q1KCWz3vsZjFXyUuUqDhmD/xTXyBD+B
ncbrbo+6+CeeRiqmt6sUaTzZBk/YFw+ctS5Azz63RNiFQ94zrcTeQi4PLlu/Os8G
YLzP2lo9f5XldAUC4lcY3Bjzyg9YSn+3rhCpmMKFeGVc2AtlXpkOfU1Yj7V1isJc
JEfNZ3lGZBzrXo9RrGngfufIGdyVP1TCzg0WR9yzd1WPyt8cJYhjf+ZjUX0LbUCu
wTyG+Vb/wWOxJFUs+qrV31//4IhB93yN/+l1bnNtiewY3B/n7kpPk5+EOfm5e+PB
xpRa2zhsfzC+2X1ROIspd+q3tLlRtYfJe+SKUnqKTFQCm38bZb47iY81970iiec5
/Ghfb1P4NQpnTJxc46AURdd7d2S44QxoWYa538mkI5uXerK93X4uYXbSWZSpN61l
AzQFdNNcRqcDqpHoeCSv2jASVbLlMN2rO7T3YuZEro1FGFgH/QCcuh79uMLqzH58
WrKMT0i0T377E0vxxZlJgTBUpWLWiN2neDpLLqE6oIMRyCAyMwm6pnieMLMdwHUC
RBczjbdG5Q5ixPh2J9SfqogxzyRVohBhaDagQHaYrbgruEvtwc5bDWoKDXzwDbBQ
JyTkMeSb7v0V1u3WryX7LiG+xJ/AIRwVga1KKQfPV9sT1K59UpRD0AKUYNI0yHPm
9zgh7+ohNn20/MxnO/E5SaKQEMx4aD5ywbWKUelI23QQoz24ortCwQ8ayFqLucHM
44GWzQoYBpqSWiCTPLpOcUGMWsfKNgi/DcNju027dhhg2ReVRgpDE/jrKKCJSluo
mgM1XOH/lmgg9MdLmRNOZQmeWq1ON92AscFYWcw+VTQTZDsyyjaD9wy1OOJwi1Zb
b8Sw7Gg1tn1guED9ruKGFErrKf7ce7E8T2Cd8r2Xxho2kyJVFvde8PYpkkmLL30m
I0ZhBPvbpyM2Rfy3R80ukhSu9SdDBw3ClmXF75NVWvuPoLW492QJww7gXIvf5gk+
Rouy8w2uP8SPkdVN+0K1hhVQeNvVG4NsfpessRGcMPV1LT0AAPjoI4WUuR0XUp/O
IYZ5JhzcpZi1NZrohz8wpRlMd4TuUrW/D8eYGdie8T7pxNgUZeE8pb9GGKP0FaIJ
TR6Cq8krB7GEBNXxZy8V15CGFcL+hjF+DkYvjVRlj7dLfmTWA1hptfNRCL+Y7jEG
fjGsW6l/uC7a/lD1pLDY7RO/gK2bipKYIUXFzATrSAO0gty8J+XWUYEQpKpeFor7
zL4Fr6lfTomFh/p4WF73c5N1bo5QRsvJkufIB+QohvEa8yn43DtN8wM6w5Aa1bCF
Byxslx5APqDMPPBwuXw6TQnTI2XBfoY/P1koRuksJ4QU13wU/vOy5OfOnHa7c42Z
PQ4uX6RPjv3pnXQri/KC3qO1BRVAVDgeDkFq1Uqks8+KYA+B4alC5teULHIMsZqd
CHbCoHOeIvxDh6fGfnEKSyLVd3o33ijp8G8pqivelpZFRzVyZHQdAcf8TuBNafci
sVFfYJ0/PhJNKswTAO4PAkn8SIrom42lSKQAKBzF1iRLgEK0kfNbUysNaWFtCIkS
2m1+KgI2yJe6wx8Ry8Xw2lVlTd6m61vdvN83y2v280wiYK6atIO6jOUYsl4V6jmB
FPHwWQXcA8Ls2FSMQswYFjFYo2fAdxS2/iwUipjvRJZT/zIIOCzitYlt7kWEFAze
jKdAoaXpDoI0zkdNls16lbVeKRO1SitGAlRyUmVzhBB0fac7+uAs00mtDGn5WfDd
yjCEaeVtGbAVuuZO2bDv8Kaw2d0lIL652S2K86G6UFSulE+hkEAySYBC+8LuRE1l
7y7FeOwDJQht0t1gO8xIgyEksng7msaNTz8gP6Yb4pnPsG9HGhPxOJGa997+n+F+
fdQ+odKJgynvPJN66bzqxnMvWe9zj/PrC/JzkFpWZRa7uWvwSMXLVs+8I+FQPC5M
BHXb8t1y5gzU1Dcn0pm1sdNv1b07B+Isn9TfXVbnNRHILoA7Qh6Ex2YG+lh6BpiP
iqCXvtao6LJ9N5sETMadU+RU1O9yBQ0hNoXiiGFYKR328tNJtnHAbcb460prgoqO
UsXRyNH7cF3FwpXsRlcZM5z6ohMYERDGWNM/vvO8tgV3XLqc6VZaWCISlZThUkao
PLqzUEwUbvLIJSxICP9PSjTm8fmLuFstbZfGK795EK5zAktAWXft5SyKxxyz5hQv
yMeQ33Hq3tCq/YzeldF0c5bZ9X3CpXUWz3M9TOAjwt8ZHmdniIfSWxef+oep66+N
pMbMCG6H1omoco22AU6hNAcV5K33B8vGcZvwHDJGHxyQPZ1uI8snOHMOl0GEtjnJ
ijuf8Q0XeVGaX1bIroRmvZ7tm764Lp87BLW2TYgZQcuuB5OwveDkp5KfN8KTFiL2
qrkSJYydXBxMucpoJHkGTaUzQfnxtnYp+5VuXBWME67tIdje7eCiNkBXodbxhXzT
gGF8b7ECP+7cPWz3A52T6HYTH2Lz1vyoyuB+3VXuiLqs7MxPmiHDsTli3DOS6B0i
07Qbkyf1NKa3iQLALI1WfkAvnLIk/DEi6RInhjJe2xBNUilirOVhvRKfVrtFHPQ8
C2TfHYBlO3bM99E6CM/dF7SgLlvD0UYcmBrHA5uVRMqoCf8lgIdrZO+tEAQe1bn1
8GdD8EInDiTZntO04BYnzK4tjXa4z0J9Jj17/9XI3CAixExXuKOjpeE/14lnwPgl
MYxRC2gJ0bPBu64+xcIEmeFBIf17FqVp0X2FLxb6NcizrwDZbjOTODnRCyoPRlcZ
Fb2n7DJn2L5dbA1djPin4WNSgaSziBZJneBO9IGuaLhZm+JMLIXJgBfXnzYuKOBl
QlCAtAf+hSx1ZTOBUQu2uwZFw8OVJkQ/DQhrhT+2wFEREBwHh1aefVgJPw4SVtN7
ey9ZcQfQwy1wa07kKFGXWMPqzc1ugzqeXUFXIvtzAP4KddnKsknnVZZuEiL7t6fS
7XrhPHbT2H/xkWLLCFIp5NQQVGuKcS756DcCXVPJE5KYWu9Lrr7dQ5Sx70e8HnpG
dtTipyeqTUiNuQTeWrNPj1WpZw6g3PjEhR1YOSgZolCLQLw+TA6cFtK69qOzyFsv
DofR3gFRWAs1TdXwvRmnKrWBY3xpZvWCheBx50R3GGdEx2q72YU4CkKNCtltBTLe
cMfdNXGFec2vAPzrROBoq4ZjsNOywYa3BK+aREkGazzOIhPxI9Bb7Ol8Qcjbpw0y
S285aE6E8snRfYtREHnxtN1uytvgPPyyFSmM+7xzSmKV+CRTD2p5Vjbg5ZOZox/O
kKEtcfcg6DSRcNRC652J5vFptlkDfKJx0qr4gdkvL2Cw4jfMO+5UOuVM/7V/N0TJ
IP5YnZKinOiRV3Az4O3nkGGWlDf2ZLbZm6jorudBFNZxb01TLJXZQ/VQ89ULv4dh
qjyh68unk2AWI5NFtDXFThgWhFXs3NEInWWxckOibkxHirHoM6J0TrXwhiLTKgH8
0sNM2kTes0+TJXK6IEQJ0UP/1JRfyWo0ADhz0IrCcUF4M4tlkz2ZAkC2w8jA3sus
Zd4ts/rNYAIAsREMC/s8ezpzjj+W2F2E49XCJHKvrh2SSgm9pB0enHHZxt4tGXIi
duy20h3cye4wcpAnNke85oztIsQ8USoLHDfK5wE9M3GN6VC9rTeaz2+M8kRaFOgi
hgITWIPEeQNILHOYkZ3lhWv7pB4Swqq0SEV/zIDI0NEKZkAd4rLNW2Y65lCVYk+B
C65nW8PQssmUXQVv0cMApqdhLMmzjPkszvSYXlyoXKI6nyLUQBkCpmmzdArgd79K
S/OA3Ccqc7LfaF7BEkGcobYtTBqnJHGkm83tb9nWDRe4Mvs1rEtoIsa4zUhIzFgd
k0TNTF/K+RpZqr3zET961wnebF89s1S6t7U0NkmEVKfvQflm4VwFLXegJHDwG/PE
WEjZFyidDiPstvEOOkYdmNpZJt/ewJQtrEAEj4CtSKOm5qBNzwNbBVgr+6OwFlIr
z6JrWqOys/DxLDDOSL0JJAMwv35eT3alE+hS1Y8NsA2F+4vlSFViaY6dPqvSgP75
vDNVvmJzL5pskgpIbkpY73z+5MayYj7wuKLA3naNETSARJyUqlnYCVZRU2h89CQj
goNSLWyFP41xax3LA7oWbvM+RAq6al3C6tt05p0yvYIOP5r/XKp8ELcbw+G0dLIU
e3phIjAEmH8IQvoQakagdiFjZR/v6i5dxAj5Yd8D9KQrYHLEWBKWfTC7b42DRNmr
YEfurA9rsaRePFSOthd5ByJlEMcdUD7Gfl0KkTdSspdNdiGkYrC+PZ1d8dHi6/7r
DY5TB2XzGsiJ+Rc/ScMuQmNUlUSP/szSvTVHlAZ/F+nsJTeZ99r6yrVG7kzKY2Zj
iqyVmv/W1x7iPuxeK9R9FAxFMUJQl7awaPwWCkBnvUNpVBEyQJamopO/AR6rZdrG
5wbN0ByloIZSYE0Tutnc6dG0M+MCFFPldxNh3ymqrY6KvjCf+OZUemV+YRu0mhit
u55MPG5vBraZmRSHewjns7lP1kmQHq+5Ho3wxsvqsuwXpj73ZMJX7dwnQl2hENrL
jglz1rVCVlkS3vOdENaZoFD+3gkWQQcgzo17DEkmSwjU5Vd/js/zmZy7dR/hcuES
gJh4m/MaEDsVzr/xVIScZnT+FAoFGeUWMytVepGgpgnYiHtGwjoJdfZzcKeajMUG
RYTzGPxnfY3UqBTYy3DN0d4vpAbwlUZqJvZJu9kRZb3bdEmxu20fe/wrLz5GwcB6
6uKdw85cIfdEMconPMFO5UbF/7oax55h8EXqR/5RxCYt/ZZNN96CakXzjU8xlPOO
WgOqsMebkGc8+K0lspsmKsfc22g4tVyCKAl8M9NLXmalgnHyESIezYEojWH+WN0B
A902w1VaGluTtY8BApXhljaPUkY890ptbgyGWFQK9PY0dTZ24uUqOwvqxymwMcS9
ZYCRNrlbxI3mS7f7NJPopmhNBXjGsY/B37D7b9fsg++QszgD0rqmgJByf7FcqiSK
ZOxd/mXD2jjXimlR/hWfAqAWvIta1JnldFO9H2ExcpL9WliTVrg5nkbwcCysJA8j
sEVkY0xvTmkNwZgK5kz+/132pxphH3HZvCztuggZeLdNcW/Y+H5+1ahFbQS5shK7
DxXpJ+jlgVWCVVQMh1eaegcc/cxMkDl4terlrrgTtB3kpREaO4LprudIQ1fWh47U
7xVepQHD06AaAz5LsvJuq1cJlXemtBeotvjOwhN2y15JjzD7mtkyGezvi+7LZibI
h54CYfqp6k5mcz8Fq0HpxcLnCKFnWomiqJhnwf2htA+073yoQR9sY5tdF90W/pD8
oZdVoponLMBzPT4/5isXiPLbPfMDA+3j45gbEUdQtlwml+VwvCoeWQ+Ld8OcuMpI
/sVuy8e1M89/eACA0+iHIb42zQGCfLPyyQo1McC8he3PWslLfF3RUMwfwTyJDSUR
WF3OsMkPVZrSQPGKDl0+uAMxwd5tDV/6WT7sg6cRMKaKPCR/50ECCMLuN8LYacUy
qJVrbQI+oym0FhZm8UlddaaXHJPqkiekTpLvveEj+xCSn28zO/KJl69d3mAgdnD3
0EUjBgeusncqYgx/bpKknWgIvhO25G7IUotQ2lyp99dCv6UsWOkowz1X8EB3I0JL
XdsSG7zZ3dPF9V0fDOVox5DuD/GMLuBHL9lhVxTVxLu95d4XbpMF/TEu/Wmnot3E
Fc8nvwFr7MWsF0vhhDOZrrWnOKOVKlV20Zs94O+CbApm3FJXb6Nq/1Aq+v/n2AuI
B0wFfIl6eDEmdODfEFUg2PYr8MBJn1kBVp0GwB6xL5uAIga+esYHBhI75f76A7gb
7cRrKmWHHUYD9HNNM1nJtU6Rv0L9r5GItjbdYggYdXKg+vpA1Vz6eL+wi4g6ECij
jOSPzIhy5sGPQdzm19k7Q7SS6ZcLOB5fHQ4ty5iVhAr+KACHcXggFJKKGcmKixmZ
PkaSFK0s71u5K/1N9cVDQIAMomf9pURiZF4W29968AhDB0xYxKlfeLfisezNHSnc
agsQpEwQH1BSkdfuyTSPJU2rS8mrxodKoEoeRWAy2clnNijTkwo6umZhtnJF5s4g
EAHGQSRqljhBp6MUQmAz0gdbmqK78PdliHZbOhKRQKFDdyZAYuuHcVj7uMmiNEI0
2fzTsHiBFyhX2erhjZfqqFGr3hShYLrfBXCiYd74q4VUX8DqiYKsDEhv9Np6SzGL
Jr7Y0x6uZqT5JBcjklWHJ943Ni9YrS/MeE+o9wXIw1KnERDebFBJIKA2WJhNLWkv
00sip7OWVVQ7G/0lnkJZrjCV+jTVfmzN+bGAWJtFDe3uUMysHsc1wep78ucyZBIK
e+Yphdh+9OJC3oqpG/IDmw+eDjj4ripOGH/ewdCYpzuMgzuD5J5N2ragB/MUm4jF
yCqt7Hbt+rQmBm4NARHuhDT32P8CoetdaNJwDW45XVZG/1eqtUje+tnlRrq3f1Jx
uahsCqyFAaJieUKS4Cog5UcVF2DSz5wVeH+0bTClqKRgZqZnSnlEtf9sVcVi+j2+
1s+8i17G87XSdan/3CI3k4sOB8Rhgex/wF3rn0YYtjPNJkEwF+9q58O14fWqu+3e
LuHi/BmjyH0GD2iV36tpSdgpjG01nQ21IIX8ZagNUuHq7YgK7m88nN49cKI+7zoD
vVwJTs3ihlDsZ/a5wLpNVUEZCIjCIhsjuv6riiQp/cel1K6CWf9LUVB/eGDSeTcA
wH1mxS6a1zU8smdz/hhXtpoKD9buBkMyxbXxa7wcyZ7I6+a4c1pH4nQIdh4SgK7Y
WkI85wIT7SeTXqGSH/7ACKCrjJ0IusYus5VCwhW7BoqcaeBUqhAtn6j3YSPMk0zg
GzIBb99Ton+wj6/SEKug/IGN4lzi1xTX1uzgS+5wBUigDtBgsKb/7KvKxwRz+NZC
FJyJNt9BbN7jt/y7zhjY4fEB/p/1nAcb5FRmiW2CB3mW35zU5CTzi+tLYJA9paIP
1mnRVOzouDg/XY0pshg9KzrNml/g1dO3Q/VF38aGZnMmDVNj2dd1dqewet/JW0HW
7TypVUZXwisykXScYSCQISGBlPa1OFCsgCTVsYIad7dadodGr+578qpBOoA0U5jP
sZLXNLPtlSOYtSiacX2hfMDPU9sdVOeoNXaf9F539YS0dNM6aVii30Us4BgAF6Da
MVUS1fpM/b9vVsdgZSuuLJRQtMLf2KuOLKlJXWPUo5uPf5OiBXLIyaTKRqiTDniQ
8CgzTQYx/1k4R/d/94fz/KtHUltceEScIOf6gp2P1BdOlIl9cdSI6koKafWgXiVP
wNwsDXmb23EjDMJirDcag3I9IfIxPabWdsEmMXAH3JuDbhkpF8O/jswWguMzIA4u
c3oge5JAWJGaM8hwcJGIy/Jw1DnK9AOWesgI7dL4UtmjMA3snHWPDRnVS9F7L23S
XrlMprpYb7j9VZE0PHC7/HEn5Mt8MtoN1CCcIiM9EfWDK+PGEpbjfEU2FJti47GA
E9wUoudtGQaLMQINfaYWSXKpBTHIHPumedvBtLtNgDyLx1NPM0dzIRXTh9dDIykl
YOIUrzLoSlrMM5WMdlxK0wxMv0wGdcQkf4f3Rrqf9XRqzXLaKjidpx1moPd9cOtD
8NfELP0A7IVWsAAZY8TzZazXOUKu5mDFujQ/nUuJJQKSN/Iz62xeKEBRvBrbis72
kEABUE4NE94/u7NhDFica4ff7tGLFH5ACbVdhfcZWNgGSjji77xiVXzFlwjee/qk
3nJclbQSxGTxiFMN/aCGMOtW0TT2UswYHqzbHRzijzYYRf4txhLaKRp2ZyPqIeW0
yxPPFCSYL/mNcT0w/mOwBzU/+oWLUDJby8RIyWfsB1zH0PkhW1WRZTw96O8YDncP
p3eJRiT2qSrwEVTDDd4WgoEbnR+eGpzDhPy8J9ZX/bFBSmcFead0EarB6GXrOdYc
/tuIoUft71N/pNF84VWcyo/AghebsXID6T6c46GUsamILjwFtVQ/gZlrICPw1PLE
MK9dd4PUs+OfXODaNPcPlIOlWSFdBthMm5fvgTcQQ3OdIne81bSmbHd1SBD10fPq
r+FoNzBW0od/UihYe9YFIVsPUdXGWBjd0xlUfDSj9xkpJColfuTOBLo6xpL5Evku
ec+X7+4/iePWV3n0xYveUAo2THRnIDH+ZyAqYQGq4EbZQ0w58Ogkyv7fCWFYkt06
VUcebIh9K24S2x1Z5jtEco2u9raQ90wJAOuXfrpIqtO5/V3HAq2ElrqneB6ujTUV
rv6gSFni7O36WzP6P5P/NqzSSddxV9VUq86Nhz6voP6eDtpkqRyoRHY3zV3xZ2yR
k9c2HcxXpPY9GxBZnyclnt+tTEQf1t4ho3am8eACRJ1YjgsY/MqdIRFsJnoT4kze
unGURaREpTpC/FK6zrP4ZiFIi8S9sExVubTt4udCsnFqaD8pKDTNzvjL+bOaBgAb
YEqeNKMJ2tPMoiNp+rzwaEvz66ueoyo9DfGBkf9fMmI2xgpZdpDc1XXJbHdQoWfz
LWfODhUg5LVMU+qC4NuOe2ONNW9N5b1IccbklCPmK1uf0AbOL2zXKR9ahSQKit18
wlE8clJxqjIu9m3BMcxbC78iRWBoyLTfjkNI/jrPhxxsbSITCrD3tL9vH5spO3oO
xjXhX/OLqffuojhe1Z0wkkVjKDiDrFySQhNJxQlTGzbLl4Bo8ldKB/XZSXwvfbmq
QjHbOp55NmXQwLVtRU/4nAWKf9wqBzXi2wNhiicqWc3Kit62MiOXCD9beRVw8SG/
I35yikd1a+/BLdABjDyadh7Akia/Qj0RqRlr5tHvMSoStfEHOSJuuEpG/7mYHw3d
EQG+ntmxEB6QfdUDb4iVN15/SVCSVhkahFItQd3/8VWeAQOcdm5cIsgnCC+VmE8A
4RW57Ux0YL5TBjd2RBkD2iTIbAmfA7bH8FJSlGVc2axJ+UZgm83A8OCr4K5G53QW
Z2BEDhJLUBm1iljFBC1MD+gATMa3tyT/IXL7fCMQMXaprgyPpvCHufRZKh9+CQK6
RGv4CQmcdzm/xtfhhdCOlTPgG0nF4H4d98vbyOMxoqN6a07wNIcDs/P/RptG28/r
Kes3+PTMNW2Qz2PecpuH/udvrMkkWgtP+a869fUdsSSqU8zgKqL7MxjiiPcTrLCA
u4Zi9+L/oVZuKzMLHd2P+TbwsKl6dyek/4r5gHvnUQLLVCC5CfP3ZMZqJ9Qc1evl
yPPy0DdSJ9ZLKPvF0/cfEu3sO+sIC3G35jrJGBgUJYDE7KyUqnl2460MfBTNKgYs
awt4cIsf7U9oDrTe4xPX3m0x3I1iEc94hgmeUWWida64gP+7UNdTNjogHnU1lAyc
PvvIaBpqlWVJiN+WXpK9Mw+oQkrUQOA9j9kn7egta3KEv1X5nssGkO8GC/+tRLJ6
gRXh4VWeiwlozql0/ga0a1N5+22rIQUw5e2xKCXHjnbRXYz80tZeDA20hRGLmkKU
C95YICAGWihwzlfLPQ2aMyMmtrnP+d28dB3T7UBw6LKkasGXGWYyRSHu+8PlcTXH
eNiMGME3aX/DGPJb6jGWqv+5JTUmDXuDxrYYfT69WXwdHGNByPfJ0iqwqxQ6Qo/R
ttvzeqJ/yenSTvIBSyxoo2BE3mIi4T7fPxZDoFCF3S4SM5QXcQkhljBRxZWZsFCa
SiMbh9coCmajtOf4/RhPjSQGQIG3qpqafatdkJSuxkT24+vyLgPUMawkGV7tNb9n
r/LIEt9CWBmufwbuDiiV+sHkgciq6726h9Yha6IgVrxUsvgV/uKsCbEomJD/3lLa
awvq/CYmbjimArAoH9QBhLOowpHNWhoRf7Wz/kTm6MpCC8Ylp75iQlbW3XkftmX3
QZykyz4TaIXor7jcAsefwxdrtAiBVHIbLf5FcqNCcUP5JwU/OGdC6A1PxfNJO7Vu
tHvM65r8xUFJlULw+nRnqoi8qwhtoHX3n693C6z573h68B503qdVqntwVxazksEp
xpM0PqK5crA84xriTD4LxC8mj8ALRFZXBiVaeJdP4I1dLmbx5BDQ3qQr2p14kJXw
3594c43GDUALNgzsBbSZ13jhDSHVzgRHRu85f3fSkA/QDTGaBgK/YzQr0z0iBnR1
Nhzj4xo2rELrZFjNL2eSp9W+9Dsq5GEzzAorraEEtE4mXQuo/CqYAbs2EU4OdpsD
zcZ4jI1yIsRpFtIbfhh0b7NnHglDIb5URzqtvkioSfYKMDScpfUyJaaWeb+Hye6E
vfQz2Z8VAbiQ7VEc9dqEq8H58/XQo4dMyjw6ItkJ4poXXZOEVGsMf1++vf2OWVtH
FBC8izPDAMkc2uQuuHwrYn4U3zjddSMydNbpqC35TqAQ4x/uuIFKE5trvos5CU9N
i0LN3LxLDNp6ad3Fnp6XLD4+CE9S/Uxf97rotscuncISNsB+14cHyZgTZPMGuDgJ
8p/pO3g2jF37TuaNkQ2XoqhjeLEayUMRUXpl+cHZLWXmbuaURYaEB0KE8Rvhq0Nf
nSDtwk3KkbqckgtE2agkh/SAvASrYkXEtR/8gtrQvTF1M+/x0jRjhB11eSLVuk48
e3eC9aCiOYvd62p6n5XWeYB0C9PpNOlGy0mnTxHhuf0c5F8wMe8STpaZLkH1mUyi
OprqB5KmMA2bYcqBnvCXrlUSDcPh4vXVuQdXdq/j8ExT7AtAWLoSsZqmgZACV+Lj
ccP0V3sCwhdzokZ+u19Dw0/QZ2xZiMLhPlf1KU7CmMMY08IAWay2FRtjQVyojZdw
uni+fp0GbFyGMjjGQnRhjo3ZhI5w27GArLuv6yDUN2QdtPmjCLgadHFofiszpwgM
sQEVj3elCfrNX3NBLAbkEdmjngwPhnjDBPa5WJ/qfuppLU41qX3SA+d3zcTAkAbp
sly4fEpjSQBh0DXfd4J6yARMUwuMgAy+eAdNEbxf+V3AeAz33LWCOCpoUSLzFqs4
tZ7noTOnklwzEGW2RjwdfiNx+48TojgNGj0EY281Doe44KRarC+i6nG+0zWnu0+/
yjQ2vEiQglukp/8ECAiHKyPeElOhYBtIytMv5FWLmiKQvsnpaLH7522Ek5ywGGhX
4+NXbNEk+z7skFn+P4Tbkur4Ir/80/GTQircmlKq4I10VtfZ6v/vijIDtyJSh1Ib
aoG+BA+TSzGJ+K9wrr6owTm00VO831RAaS8koOJ7j37MTusc2l6LloL6GB+lqCTT
sxy4rV8uglkDDPNmS36xq0BF0TSn8plNZnCRvvW05zevZEbKLnYDY3fNGzK+Yy43
NXD0nx5gUaRedtYkybFf+7QcQZxwzsN5GLtaID9c0kAXcGgP5U7xax2ifUIDATnE
0Ud7j6ZfQqf1Ana291xq0LuMNHJYINC7UF/JjtdEmsfQAfTnFtrl9CtntOnzYn9M
jgwRn8SYXr/XhoCLep5l0fyEPpNZ7KKvOJrymZcPwGAS3xpXeCyLkg5KdwXjGXR2
G7xrj0OmVKv2dhyWezOLXxYdbX42U1Fzd6BvtYLTjIZ7vMSEIctm9sEyrmU7Vzhl
Yyw9z1eCOK09J5XlSAxRq5h7/1qBSAU7eoO+UeO0iT3Lml7FiyzuPqKGL9ihG1/Q
JbJX5S2uqLpqLwikFgdUrCeRxSK17hNMTuUnrDznXJCZOtL8mAzn3iROVUMi9Oa9
UNqYZCt1OxuQK7r40fzv6ZGpvb3dUyRDrvIlbJpAcqz6fG7Swi94bEWgtOZZ9nwv
ZKOhkHOWvjYqH48iHsZBYdz0MSdxf8zmWcvQiGOsSBcLXnm7VCOch1yunlxszXhZ
L5ePHbG3QboxgSJaelbGC3QPo65xjwFxGsLnT/LZknJEHcT99ndDbhhroJ3z9Nw8
jiRowDpFma5i9plLNfiGrS0jQ4fCquE6Uy0g8gggGt5qdE4iwBS7aErBrcTIhS+z
khRNszNR4Hbs90irJ//pGg7VsgLujV54FAcWgfop5vPELkSTbtDvl6fvz8D5k5yV
GQS9Wri24+d1t7GbnFOFjnnzuvKYXtE44bveclPul+18WH4G9SkjHYdEcItuYcF/
OjBztB0AQSLWFl3oaoO0rhiRGWj5Hf0EXUO7kWFpGdAUU4yxIbcAspzCKc13VCKr
nB+lHdPbNlbfnKwXxsicVaFWwti04inpIAfr1+ZP+bfrO85Z4lyerkOy1raGgzdG
tNgODygqGNyAlVMF4PV58qM22FfVRI/82ZqnvX/q4Y6WxSNsXmb2mijhFw9YkEom
k4c3wCDFIqogxAGagsvNK+ZPgGpPHqIMoXbo46FmPcCJO2w0MaWtQX+lbh+/7nnt
BYyw7l26CyJ3pVDnP5EM2N77BML4drTb9+oIfJMKrOTuud/kRk/tbzpSyQI+cWrZ
MjBVsVGnKsc+Asmg9JGdSPVOMf5dIAda/u1wPn8pBghqxBvHhXtD4mTshG8TP3MN
e7tTUupmUur5tTQp9HJmOvCMT2S81Bha6sULR66g5SjcvAzY2VXdY4h4twVN2HPe
eet2QVDr39FVRLMgGg0oRr3vm2ibTGIYyulNo4gJDZIEIJNgosBKPUplpACNRekG
IEcRF28ueWtmEu0tJy+UdaWeu49WxL6WFXGIZBXTl0p3mW0r1M+gmYexkkVaF5+f
PUsn58Nzx7w/GBMluvO6MOuPTwaBSFISpzBGEZRbUrlduhGGUOfKXgXjjXfMGJVG
MSd2sMUXZbkd8XOlH18LW8l4q+PXq2UAp1MQTL6D/wgA/57Yxk6kvq78lCM/JiZ9
rEKmvdTTtvsfILsxtrXDqYt1Ue+Bh57yN8JiLzew+IbWsesop95jfGWseyZG/foC
Ic8nxa2HAoFizAfKaKcmdmnLNVciU9eciEM1O0AxLbygEiB3JBMRk97Q150QIKFK
KBCqMlnd0Ycu9IWjefwTsA/R0DDxUHQN5k5ztoGKVOmM93PK8z8xBFyK05vVyQxd
20VyWn1B83BK8J0n1zwQQaknJMx6Gt4QU+K1gcVATw3AezBUNurPSKwYgG889mp7
uzTIOJ7YU6PyH1Clt5kOPYFOXIzocwTTOWCGNfkA1QH29qATJ0k3jg0WFjA6LLOp
AKFMuVdaSq1sr1aeIfQ9vye47mi6ejGjmbr2s/5ICar4Ce0Tx1/YGPvwUN4GPNnv
EDPZUvvxkr7NFJIhOGKNKCYdDjwcPSkjCml/snwG4G9sFbkicAGd58y/TOIIfNUI
c/W4CzhQpu9ge0qoXBR72GXtppSVCdPw3iOhJXu+oZWPmfcPnoZrvGaA1B5bnyi2
KMuCsUafHAgzX0eBE1q1wNtarjpy4x1nGE7otHDORiGIR41CJDqEobKfMwXz8TTH
0wxGW4M5lpYK5guf4sa50Mo3Gow+xNXPH+CJPGAeoG7IwAuHEEycgb64+X083vl/
9gxu+r6ZmJ01pEUkHM6kaAGtOg6dVneU2JpMoKbOMQ8vpCmVn39/6sbxgLpa4vnv
XRBtj05FB6+xf4bthXigNh18QZbrexrSU11v8SpG2tng4o9AH6fxWhuZ/EKQl70+
WouwLM/0wDGqNHxQ64txDEwopZAsrfZ1Yy7HyAsJaPcAxN/N+hVo0vgoz68ZQvqb
N7M3CxGWegW9RMpPogbmRRi8IAbMewedu7QFrDlwktcD9h9sDGFMd40zG43xh9T4
oKTbINlVi/N5OTF8/z4PXv4EClb9QKsbcKoxUvc8WYFLFx61nx7X4W7hPbF6f1EW
hYkSm5ww3qJrPmL18IE3wOnOe0GLNSgAV1kEnPBYLI1w6EI16WQ5tD0XY/Tqj5Tw
d1f+eOhCxpnnXng/okJNf9YSH/z9GBnzHKFTv34ti6/N8BlzF0+ZbodRoKQt7og2
fjXYT4g5zFMSfg9S1gooihpMlciAhsCuz/NyPV++aeZLLcHD9MZ3Z1v/dmjhYf5y
/8i8PckA58ITuTEW6/qh02aM6tpG8RvFyP/++7C261wdKe7rIxiOr8vib5mdCMht
a2kAtSRnoDCbMoDMqwrpS7mZUWZErL81udOkK4dDh2KmNtmTY4B81UpvHJgVPofB
AMbkwAZbhBt5uPtGJ1ap7I1p1jkUYt3IzpvufNjuAFxGnxk2CQpbfCeQJAsmEt2i
lDhiRRSZHKCsnwU8iShg//Cq3HnnOealS3eBaR7jnI/Kp87n/bHUFFzpFy9Ef/SM
a2FMxm8O5tSNIRfFlURwMrjT5F0eR1zxOOihdYxNLDCli55mVzpxBHIePVurwQcA
drcwT5NbpF2ZdpBOLf1ls2/Icku08ZFUovpSsJoXIOzT8DiyPMHP1d7ry/95B3zW
AYiL8TjWG4wsMN1qeecifH4qnE155VwMTknWoyLygNE1m9t+fEnf6QkkAymjDKX2
pZAmY2bXsNJ6isERrhWCsg9ZuT9R3c1SqiSB6pR/OwaDp9Ci62Sc7PuFneC8Aw2M
1JstPiKLRWsma1O52HlSFExqpm8T9inToTN1/XjoVrTWaj2NczDBn7QiSLrybLmf
iHSSiLjdMrO7l9Cs7vyBXi7MbhSIsD58DdfRm0RXX4UvIcEV4dJHbDUJPMIL6urV
JnpQDF3egqqBcMnObXzqhX3Jqr5FqR+If3Wz9VHwBRXMYJAW3Aae5FgUMBkTc785
KigZBs8W56HvTnTOX2XqfECS1I2yJj0uEyEfZB/lAW6JkxJYC3sZshpGKfYHcOQE
kgrKJ6KJcui0FBlDBAGUboMQrtVBUh2h6YJo8+i3AfG6E2BwBL/1d75W4LjpttO3
WRfHwQA+Mt04lICh9JsARbd4oPKdzb/fGIMLo3QgF3ZNtKsGsOPl08rGtgtpycq0
b/P8D5GlWhVYwgY+DlYmmasAeFzOEdpdYc2WshSl0Z3IBEYnBeS0BFw/TS1vK2vp
xn7oqsVn9hR+yF1mEI1x9kBLJ5wrlI9Yev58m6kkB5bNAXCzrhiTOFHkfxCiNL+G
PIj0ockDFVKWWh45OMAAxYuboOtjZxqt5ibDuWI4oXkTm9rpjHGJdnq3clZm96BO
R/Y2gLye2eevogo4Y/R4vceGzp+tyD6LPL+COSzMn053bmj8MjHEndtwY3BkCjU0
M0u/bbDUmZzGUgHzYId1NnUUMJOyDP7xxcD/TjmzpfvZNtww/Gw/uoedjAxMosDo
UvG7I5+KEGc62zLWxvyo4AfoUZzkWHJjqID2qigj4Z56lz2q0OZXJPYc9tCKuw5U
wCiy8d+U+5l/IiSCeliPqzm88PttUudqyvVtuYYJHX8y2eukq2ugTiaa6/2hkvBP
yo4dF97jag3NfZ3kas+64U90/uFWoflIEtVkftoUvLYZfQpwDfRDvKNsMNJXb6jz
9iTScn4Km/qxBcbf3Z2NyXqo6R46qK2qRIvMfeQ7oahRv8GPrIhPmWOBAJZU31e/
q1O1jsNmZ5rgdVPjliGJa7Br9VkTYbdsBA+BDZuztKmNWQXU9vF95OpPgAXvgpJK
DvL+eL2rW1nmT5MfNy6lc4NH07o5M6l96hHKq1xgnGcY00SKxxnDq9hAOUz9hzZr
BJHeauCGoPXSAwZUY7J5Zbzf9gGhsUBc6S63ZOT9XE7N1cxLlGFPqlWWUIAe+HiH
9oKuc+aoHE51BikXcjG/lrLLJb4vVhkRg8dytpTvvYd7N8bj6fJ/D1PLD1JIYa6q
AIMPOrUJubCkwnm58jottXgbXNvyudDUcQlH4f41sha3vVHZ0ggM5lZC7jj/Ndsb
V8shaQIT7s+8yaqGrfQYhVKfeV9IMPcOeEPNSW/Vv8CaSWPSkdG9GPEoZxGW9X5m
mqb3GtpDWvbLDu+vDYPaKgYnIC1Vz+AgsEJ8+IR+cRhKK13bujH4PHWxrLOEYdOp
QpSLyz09qEWYEipSWgcJPNv1YQwOJn3OuHZ6pRuUGm84X02nHTrGGOCam9WWSPEK
P4sQEpO20cm+ThziTgpA311tvqqH5RD63Shbu1rOKD8viHcHlvPdK+VEc/FbMypw
t2GV+/iha8hTPc3qP6vfxeyzGC0UKjNAeolELknsAZG3IbL2IOj+VyZC8vCldhXC
7jgS6IyR/vuSIb0BeDn+Xwp1oFpJhPO+6j8V4ZtVNRKu3Re7fqJnR0hd0MZBnd6e
oBEUS+KvuJzMlk1XA4plyOJ7OBFI3JPeGoHgmUMfON4Z7eNWssACPla+rbtFWo0U
ENSyoMs6JE7UX/XBIuyQKsIVuQX8W2ORU+E6iHP6NBwu9FPvkxo5cs6oX6UXNvbH
bVqfmqseyc0/3ex0bMVO6x5uDzvYIZuh25ci+6cFoeah5De4ji0S8U1iBlusljj+
T3fLdmL5xZpTEd9BULS+WEvQQmB59IU6iM+mXgHjByfRiClybrxv4LorSj8afsAE
LkY0vHOY1Bq0hjSzlWSAUvSKTVUBuuOjm89tQTvmenlvizFNNMCCQARhRkEnWdHB
pzSlyUmmdr90e+gIyEVd1g0oJ7F6xktfGYPyEafCOnwQfmDA6vKSpntOTAZVK8gd
B5g0gaoXfwI9nB/bE2bMGGIPtMW7vCXb0v9RA1IQVE0u+NwYhhBGrii4zYwRcyx6
zdvZ7jzTY4AKd1hrRFK2faPKljGTdftf9dRQCEiLvzS1ECXSIKzmPEkOEZXu1K0W
vyW5/6FiMFjsGJDliGbh/KF6VVThmh+49/NXlhTXBkNsVMoeV2vy9Nnzx5dRfrI8
LH6LIkL5IM4wW5/UeEkhbM4pc4LP4tnYmgLcLWMekfWMlfL5Qwo2xh1tK0Sg85D6
2UxnlMtyOOOEYF/N2AmLidE5UtiJgTuGmuyAHS4zvq6MEJAOtKsO8OmKcK4A0Cq0
PzptnCpsf1D6WSWGeVb2jh41ZVGeC5ed9+v+4tauDnPG51kgmJ2IBDcIJOBPCdCw
ovbahfhAB3+NFst+BQoGjW7GQbpPV/Grq5jsRagXFYdH8JbFYTEmHjGliXTuRNJb
kNqrs690bbznHzvm69Jvyqbd62ki5fQPV3lo5ZQbSmiN91ciCCueyGU/2eCNIaqv
jMpo+GjjHSglF/MPoLpKUY6Jk6hB+LZ4hYC1xCY7l6y48gnY/M238Hm90WWsXaJ2
7UmeZhzNhTBq/JM9YYwNNT9KY+EiqTiETiVtCFmUjEzeXDaj+A6AKpYy5wkvwL98
ygLKL0GmgeIraZFXhswR6wU0WaMBIKpR1Car8DRqTxj3ALCTIyR3On7SEAHE7Dwl
0nMo7bY8IuvnenF4vFU5WrA/na326EtxdToqmp7XClNKb68xmHdefqRSzkfPmS1K
VEyUPrJVwnctgyTNQjUOrTr4KZJlrpqZZH7SxT4V/bHwt9ViGOldkZrrPi6xxXA+
WxJLdNOx47P3nEkGYv9oQ1Pvlgyf72axrNj4zGp0f6ijPRBvuwzHtBQ5+LaDj/mB
ZAQx+hylCn1gTsfE5EL39v9HO+KiatbfUwDoeVk0hzPv2uZi2T4Eg76wLXcV089P
00PpAiqQzj5GoL4DlkmX2zAt6vT5Qlv2y3Q6R+Z0oBf049aH2rIAP1kgdoPkPwuO
hD5Q9o835DdqBQWMm1bmZNf/gzUYAypsnFVCkgj+oCkQj4dZkQihFzv0HcWj9TMd
scEq/ZJz+T+zTPvXyp3kb0xaaHlR44kJLYDPzx62Vlfrg8es34sfT1CzoSHAfWh1
W96Dbrbjz1mwhlSfnqCVOjcowtu1Twej0C1o+1RR4ecg0LCHhtKnDAMSaxT5FsZo
ZQWiv2Po2POKQlzUOXHFp3jsexbJzTiVwPbZAlLCH0+cY+evNGwpJi/JJJw4ZRBO
DQRGu2dhTHV1SGX781OWZKJBzCXSWCmMShQP2J/A1Oc0iZChCpdJFJHaZVdda4Gn
NPaf/bZ4TOszbyJNFCDHdWb4TReQROgbiHeZcH/k9drmDcbfj+tQGIv1W3EUti5e
ke0zyGw8hGX5bj5Z+0O5S35YgwPJFJRuti04LuhFKrrvVMT5fIq7iY/sluG32kXR
L6VDP8V4Wv70MEGrerySW/TXn3Cq+qMubLIvMjDW13SGpKXQIYsWq34hyWPpXEDH
FsaMbNr/9vvxD5oT7w7CUglGowLA585bPwmnQfUU1xg+pPXDS0I0l5Kz/JIoSbWn
/0wayJH+6cZqD+xbL6qhWlerDsMtiPddVuf7vxMsFRgnHkw82W5posQ4WmUdr4/5
7WeYh8dkMhNLPa14WFA5BULFAIfws1dfaYrn4y/5KJfUp9kem6Q8kQMzFSzVGIRG
m0eY+cpvb3EL4TvQK0LzRoA4EOqNpE2K6Hek+Nvf1sZc0jIyrBnPG2xogTQ6TyUb
Lj7zegZ6fKzS5kRNHuOSHYWS0ZhB4QAIJyPKwtIkfPReF5H2PCU786RVAZ5vkgZR
1JzyWrGkbKE5u0MDMkKfu6NoEr397KMdaPHRP7B0QskMlbSPu36rDPvU7K1shp66
++JZQY5ZlGtYwIqsa9PT6Kdss+tsztQ1ZmupZeGdxDNX1LB1MdlXsH0gIJG360mj
3zFd/qw3484YNsqMTSot35wHlD+ATnEFEi9yvTeLHXPKt1qGrdv8JKFGjlx4hsZj
VUYIf+BzKv2tgBXVAGQPVCK5lWR0ofDNkCUum7M/FqG9oPf+ZwdDzQ9kNfC26wDy
ZcMGWSmR9ZZOhDFSGR4oTJBz/MGjD2C/N5sSUNfaaePLJ1gW5+H5tYX7zXO6qc5e
TTZR8ao3yqOTjh1V3/BY0yWZHxB3PQRDZQHiKsYWGQQHuFaOCTDBCqdE37qnZXga
tep/j1IoDbfnyn/pgXg2+jRU++NjXxWN03YMPRTh126WwH914zACYpVjCsiTPH7D
puWS6ActnnhuvpyKGU4EU84DWI71h11Lzx7+4IFsHVSyae3YpIGEqns27wcLxCnG
lLk8oQQzncXgjnebQzKmTgdxD+/RaG44CC8k/QmPmZWj6BL4aRBHfQLN1lvuiPnR
pGS0IO4wQsVVwaUeuncE+rxSHzuMO1Z1d0HbA9q6ygaNcd0AttD4/k232+Tvoh6y
I0cBgY44pA53kOGmzUo2KIBEU4tdILw8cUidf9oNNfWGgKRL8mAHLZLj9ym/r4ks
tQ0LWFhXKk/ZsJcsz8sP1sSO3ZVmIJbQGTxodv+YrHHuS9UCusBgzIjCi8/bk4D7
vuqrSQue2ga61adMhnkIihC37f3CDs+7nGDAZJ5FDKBorFCTRespiNT5qIsKCXTN
FiQXldhOwPgsfiWXtDUUANT0At0jdy9qM1bT4t5rFFpHocjQ8XJIeI2RfRJWvhvX
lUN/m4csJcRG7vJ3w+fB/FQdRMi6xDWyWXXGlzJ90gGTxF9UxHMY2DcNQorUo+yO
9LmU06m5IgzV1igXISAsWbJ0UTeeNAj9TB7nXzNFQAE5xI3kffzNliImzupmY1Bv
vq9ck5gXaOOv+A1142VmHEL0vxd3dW87VVY6MnCHP6HRmYAOSTTrxpWNdo0SiaaM
Bn0QXtTvN0TMC98II1yTtLaeNJdxz4A1pTe400xaoPFRcqxHgDEZwE3P471XHwKu
xVgDtaDUHQFvz0CDToqbDXXr2+mBfbnYoYtzhX9KFdRz60yBEK1NN6EFbqJMN6TN
oVC9uqdq8aNtIxcckdIWEAa33kDWyzweqO6sEzwyAd84vIlFddYA4X7XZv1nDQWP
cPdmPzTnIqzdNYiGfnNNwco6mXskldCU/Un/S4PlvruoRIM9g1ofnfBq1Uh0XkED
L82Te7wfo1Ph4JLjYv5T/wuG2DeHrI33bxn0+8gg3zMV8vjoZpoOQ9GknhyOevhl
dI/mzpw6OFCadDpZQQpGEOYj7r3AsYPbumPzNY7kyVg1MGvBiF8jV0HceTjRSdvy
21sM3BjT9DM2SXsS1jaiUNNLpBtTW6nUAS4DZ795gFTB1iI0Zq7jt03nS1y/gOU1
TKy84Y7vligpIx2tR9MNgYCw/cuX+yM/YLk7tZh8Y3Fle3gqMuFQHyydzA6KDRah
X2p5dU0pdg+frpyu4Ef16LNTvOOMNC4emmCybcuwk4RK+tZmgtkz9ISYc/t+6BXd
SbdwKVAy/LeoX8k4I7Cf39o2NbGPFgPWq0wpYcrrR448CNHvOjBdcYBzZzqF3lKv
l+spv9u0h3MmIL1turaSNen96S7m8SFJ7KrNDY45zVOgSxTJs0CDxbIZiZitWk7G
edVjneBq4idJZJ28FuCVCQWZUsQ8Ud5GZ4bTTRaoh2ogg5z3RttO+niwgtwkwf9j
6HUdNg0YqEntAEPlwCKeMQ+U0EaX6PxjwlLwUP+xbroBYI8rONcla88Q4GO4R5lW
d44b9YwBjmaxUOb0LcDfZw4hy3N9NQdAwdnksWctpyJnLtw0U2qAKnZ9z6FykaWy
ZkoZ218pUumBnOQqj/4Ix4yM+g1LGBf7N7t4TtYHD7ZF0VEQV8/KQzepUyc7TAFh
30Tx3EukoWP3I8AwitHWi7VURPN8F8GBfDpU9LUB/dxf1TQbDK3CwaFKyDOqj5ml
kTGoNZmpcfQ2dZ5BHb4cMnq+jzmEHdh9Ldfju5npMtr0+ioLceF2+HEzYXWmMHqq
1wsSI7Gb/11Lnyttfd6uDNSYTCPpU/EBT+17It+XFjOK1ybtOFmjZxJ8bRn94uEg
se6Q9VHRSeZ9QexgHegFD68Jqmj5WgT5LFKJe0QOhfDKZOv/uSueLeQZAK/HdijY
/D3M4284lUTRJZRaHVPpDb2BYEsv9Vfc0QSrpp1WXJID6BbFlYYfE8gUycQ2n5fK
WZTnuzG2OW9q7rEgGsdalJ9djG/myze8kKp9zrKcMbhWEIAGLPTodChvdAWNJPkP
E+BKtjtPvRFZb3PKpk6zZijG5neIop9mW5Dxak3MfwIi3dvGs3Q3+ttRR59qwOyQ
kp25ytgSFsQcJHIBd+NJGOxpxcfogcjw/jeVSBrg8dlu3HIyS9LrZjZHz5Bm1ryY
aYc987P+PLN+tdOqGOvC6SaNllL3JLe9XBCeIwnYXlqHEUiBBywvoAroFVxL1aPr
s+wYP3ecT6Im2YtSCPhUDkIR/ulo8TA4fVX1oqbaZVEbgfehEybrJmTWoeaKpRQL
MXK0wYchUL2rI6x2QP1+auWSWAFErIPvq9GekYSmjaiuzBtA1idRATyu4xexR9yL
liVinPz1+5T0lk76l0hi9bJVhwtvE6+iUIcjLPep+lVfiB3P0SRd0kgPendSZMUO
QEmIc2+2khS9pt3TdkMiysLSq6gD5tY4g1xNYEuD4fMPp0f7Km+w0edpGHopq3pF
IVVW3qTgmDu2Hz2qUwHI8RwMjNXI5ndRBpbRs/0dpWnChSrewT5GNFgs40PcFSZK
pWMUDSNJ0M/6kVpdYqoVRRgiUGgcduUvjZX4ev0ZdD3sRjf2VOrlfqmUnan9I5xO
NBT+3wGTs+IQixkmNE217uXAeA2bbU7micMkEkNI4jAvofRODCBsKualHi9V6YMq
SnRH1Dgs1Cg5CdY0uRZVbQSDBeWRAZLuTcoLats/PL/ovW+6cIWhgEVIQOsu6l3r
c+/rptsiSZiUz53rX8ja0fRAyLUZcatHnn6k4yuXwJSxnpnyBPEgNLE16PMzlbwd
izXErGTbBlSU/XS328k7hySxIJX7PGGnS6Vf2xpuYvugtmGoUpvKLNLE15dfj36P
Dlb50dEkV1VpIpcwZf4/BOipRHFlpYeWV/1TYZgNT9IaRUfqQUUFeBvytxqY41mj
vpjsVjU9TyiFQlGoOF69QoB9LtNhIKZCZ4qDeXegtzeNtvJ72OZaZayDK6c0ve3D
xkqRWtcRiIrKm8qTzVQgdqxtBhRjZVXMWiNB1o7vWyu/ztOfgAx2ajBQzYYsPTbn
ItHHTFlM1EoLhduk7UutZHt5SM4Ao9Uw54RpkADJC9McEawFunJaLdxQ6R1ofGYj
uESDwphAChnDIlwVkyQVkyxSQVb86KjjofN1KggWJp0hqoJzq6UX629AeFk+tQUU
bubGajz9T3mgU6QTux4/nGX/P3D6oGH+cy2M7el53eXXo6Kbr41bm2kDmmcDNP8s
WZW1DAOoMiKEK8TCykH2EOVc6nhStxh3VGOdDNK4OrUBxAgfukL+ZCxrjSrGPYfK
Dbef0BJcWUkHw2LBDdjEXQuO12SOf0pZ6dSt1CyKpVJKIZ6OEvFSMPoSarTyI/6C
pEXKa8KCB/YWrdPwvuKWIzvmlwsSqMzb+0JpJXqHKhjffZiMyZs5NXy22kK/z4Zh
ObfAJNuRwIDmNPw0FZVW4SroxTa4NTOL90NH/WC15YinGcHVCPex+JVGU2cAHBpo
//5hl3rtc4R7ke+QeSDBFHu0O/3BQ+D/awS1n9vvLMlv8VC6+lYnzmUvKawE6+gW
lRXUIv6aB3WF/fv+wgFVup6j5B35ChoBUqhX0PP66wbz85Ad2W9SsBrI8KWOhpFP
xWgTEOG5tXzzXkw3HMWWX61fo6tWFViW7PifRMUmtx8QF5KjgmROzYudU0I1PUWg
i9ZFuvky7WqbtQ2h1UdfTRZyBrfrwLcB8/oDDedGueBtU5GdCpOmPkppFq/oSc3r
hBpzHOk9Cht/DT0g4/jR2SWEWIDyHuOl7OEOAaPcxEBzlXZ35YWFKeZlZUyHEINJ
QwV7BLUNKKmtnCeZFqk6T2tsB1Wj+SZ3/4rEbcYVI/94FzggT1nmx0c+iXpZS4AG
axbbqUWx0FGps2ZrMmS6UEkG3e3pHgqGFAke5eXIYyjsIfeePEt84M4xhwjuMx+A
YzIbzN2o8r4RVdN9f1QPfTDKhFGRDmS1CiV7EukvothJuGQyIRPerm82JiFhGKDZ
759Af3upqdGlFzfpDYzq5FYso8CsG1+fYr0KekxxtmwSQJ59PloWHyGPM3tbdz8m
7Z5NJvWfBldFmyjibW8Tri70kJ39lqxv3LVLwLPgfLhOUJbQadRo/3HsFxMRVGFU
EjLdlXscpQDkwO6BHvtjDajuWgk0wze/8+vUEk1z6ZDuCxWtGqQyJN4kUPEvv8cX
pKcMOkLVkyMNmbCdCoyGD2CkfO2Uzq+Bkhm63mx0TZI/smi78NFlrwWpVtbJZbR9
9iCR8r/9Lkjawm6wfVBK7AF+n7D4hcEDunmcwKvxHyv9jo2F5yo5UsavLHJEWkRy
WidgQL+Doj2Vu6w+o08xA3GgGspklLPGNCZ3GnO14q9I7uHLB0Ko8KHFjtJutVbd
XB2vNVr01+gCUzpRtANV0+fjBC8kpg833Zwg9DPlHt0mbxmikVw+JizXskmx06tw
fxHZIiTwFGol/nE12ro/6cCy1sjexFKtsKw5gmv2kJfkYxiVnFP8Wi8mcCkbZTO6
fkhbDq7H+lSWhXAbxhhqzIwyX2AuD5RUiY7WD52nfHOvwq/+zD7fI3zIf2ta69MN
zFrMvYQvYXH2XLP3ShJQcIBnLZO6Y4HZVMlLQrQu2WpOXO5nsW9BRaR1w2VaXxLB
YSzxQvAYft3k1o4E3yEcxdJHY1uVAZHM1NCuA+pO0G8io8lLIoKrUnmbiacqC8KI
Hu0YSTDkMoxScPM2VGDwSXsSRpiLeKDY9m97t5mKbWhchhueRdCSxlbFga5TT1fp
PBwSHk8HSzgL5yH4F6iM6mQR+uMlgyQsp0fEsHKThTh3/RgXAmH6X6hhQtfJFPkv
mRwTceBiL9b91Zxtze3LcLpVdj/0ooj08Fl2N538ctDl0eENB8oVY6VlV2jJmAh9
wZlD7o42h4+wF0BqbNms5yHyGZNYZ3ekLrv8LrWk5Mo/LHOi76AFoRX0ucakS1yr
ePw15AcHtftGCrg2iI3uRz0ptCyhwlTcWG5nxLPtqmciLoQ05apcZa2JSqNFlMR/
EF9HQyEN16p/w86vr3dfCM0L1jA4vDa3WDbWvMxDUBeu3Bnvk28gCG2mtLbRH0Kw
a1dn4OW1GD9ZUNw/MaOIbSjQnrvHyDREPlCvqWecbQCUo4Ex/vSbsu6SU2jHACme
iAPb5NAi7Z8HHp2rAzWM3ewfZOxzb5qStESCM/WUNOSJlE5lz0iUyqKhQ/KpfYu1
LzMJO4Jr8ljCcFFyo1pqJWs91ltV9m7PgvwRPZDQ5JrUfxncSkWggyFHD5oNkuyR
n9izCSazyUBPI02t/qlKLoFtOmaGmC1Ym6L3WHkIMUbMsHjPEwTQOEz0z0pqgNRs
sRfIWWcddCM46grYdapHH8e54eg7zJH/lEPByyAj5THuVHOrKvAKSqUpffvmLVzl
tCiDxB94/1bDkfvKJ34D7PymGf4WrrizMDtisXifKIQp5zcF4N1JIn2T9otdV1hz
WdGvZ92OIgFYMON1Dq5C4Iga5qLCkAHmlVN1H6+bFWgV5ucNbHyAQxjNTkb4yWy3
gYQSn6ga7mnFCuc4h1EwV/WGiYq8qe0MkwCKpDQCHC/P25VgDdoWjqJPJXclEIBw
kd0Z+TwuZyqpq6FGkqMahM+97lUk7MxXn1F27QoWiRTb2/n8migsWZf571kI6bXZ
Lr/d8cFskggEj6oNfFd5c22X/DSdwRpeeNCRcdNbKewsUT7ZVf8WZpORPa7gUTx4
UsApL/g7g9UL8eni9Z+r8G9g3DFkg+ifBYK91auz1CxOqa4nKspjtuo/oaLz/UzB
anzUKZu8GMZzpBnCT1t6EbsZiFnwVrfIEeh77RLWyVMntCcp7bcbbtn+Qv2VNiyx
f8NMDY9uEfO05a/Gpc5U09pD2O/YfruPXrzyIu7rsIEC85T2/Xi5HjjpaOa6Ojpv
8oKbm0gBDijd6G8r6F1VZjjX0z/5VRc7qqGiDM9AwYxhCNxDVsCw10szFZ8sqijs
Wl2z/h2pyWH9dlk7Ehd8CiGDzHV3qP90ZWOQzYtas9n4htOgidbxgBsQimgFhfcO
5w6siKbDAzJSI+N2KCn9GfB4lsAQ/1QlsdnNSItD4qv3iYnEcXJhPhjfseFqLqV7
ZY7J2GOzBhGcvfXEd5aowyIoabPYKzCYNLKxxpORe3pdwDewZQNWKcTluYbIAIf9
9WmXmPo02tCkrbRUXIZzDY8lCEXY77xplGaIaGseR/CZtSmydfZRoNQFK0TrC1cp
b200Nk++LMhwh5NGNZRxuAh2LiZToUG5kM03IR3VwiMRRa2ne9iePZnCh/uFKCRV
Snwc1NVwd9OfJpppwm02DsDyen5JAUMc7Sjwk5tZiQHhU6btKY+Zgq7O2eOMIknW
HEmLrvl1YmYElZHqW16hqKdu1eyTWZpkaxhiG1FOytgAIc/OWdo7tY7/bpjNGD3i
+biYReAY8SJ+L08/quHN0bp29O/SVVwmtbsw2HM0ZaxCsKE7qRbNn9L30gv+716i
tk+8e4wruppSl28rNwD06E4f0PT9LQf2XhwXuxvdvzRNOo0CoLGpFelgbHY7oX4I
Keutaqwqfg36NOHh543V56MASC5bQm8C2nmvPSB21C6siwtJyJul4iFJwXMkpggM
O5+FyT8UC8/PkAUrLv24a+RdiNSJ3EfwzJM0q/1Q9AA9wP6MBPAnOdYQ6dfFB4RE
2KVEx9JxQKIpvIoN5O7lBwq7hEQvVR6MFOgY/CcnGTNeLSf63uzlXAr5agPnb7SO
pVAG+s4lwELdm01RyYeBDyO/fG/XFmdXQGgod/eCbG+dmNxFNOpD2KimZxNYjm7K
PBmNkl87w3+ZbtPmrw6COqR6gqDHcCvNGcYliary+7pb4pkMFWWGWTf5dgc7IoH5
zDUDq1RewjtsG4Rd/5+ouH3WEZ5jRidHlhA+mhOgkOJ69nqfIpS49VnWhQU8lJcA
6zAFW8aXn3c6LIynYaSKP83WCfi+c/5J8SxZU7PyJGz1WkOBCralQV7V4MmIlE5+
MQbcujTJlgbxOTv8ZPZN8n+tLepADlfw1vpTL7w0NmIrAqLYjGy+YOFD108UvcQq
frqDFXn/rIUQm/6atKSdiPDa5ntFG+X5U2G29xIr0mzpesfcdP4JrSifnodnjwTu
VtosK1cL0mUKCgzoKuAJRQWogj2AhwrvB9v7zwR0A3JS7hD4+Fb/MX3W0qoOO5E6
xIynUJ0osT8Cr6tDs+1uxmiMjrBxGH2KCsR+OFd7itTtBl283nMskzm6olGE2HJa
jSZWXbeDxDq3DrHULYFUGYuGyimgP2kcvbj4g5jyQAD/VEGJUBw64iB332T6YiK7
v5ecXcUMsX9k1kdUF3ob0oV56/NZkI5mfyUX0/4UycQad/bQAW/hVcAzt8jg7ZwX
vr2LNX+z8Y17XDaskwu5wc9x7/bTe4GavDCHcP61w2yqXNfE1XUS+u0s/CLs7J8v
b396jqRA2WoQRL5wXf/4xZBDHXADNSLiLSeccjmx6FxHSfgDoccXpA0aBy00O1QM
r+cA4AO6kFM0W3DALq8XvdWUPr5L8oPblcjC3lMj4hwdRCKeshViZNzeuGejJoot
hYFqsueWfOkLnqxuaPHLcy3SXFMHV71ZkGAv5CWyvPPTkp0HyW7qY/li0auY6kfe
BOawW+diac4VnGDZYZynKItd2DCPAmM4HCxdB4gv4Zf0eC6MXUSHD925MBSOIisM
9sjuMetlkGr2Y2rxJfbg0/HHVr02noqWNCz9WqiHxSL/m5yVbDp/E+UaW6MKGONz
LEtg4GwP53WPKO0V+LTVU8OsbYT9jpP6+RGqS4dLGy2nKgw5rpT/s5Jau6qwN+/J
q8UxKP+4LdOZNCiv1xIp29yFs4Db1c5y23yeXsdW/JOSO9FsMI6ir4/s2cpMY/pY
byeuqvSzpOcfngMpQAgZdY57l04B06RSeo0YTAf4hA97b4Tq6sq6wGWpJUMMLHFr
FfzdTDw2KiB9h9SWMeuWuKFEAigmvBwrSsuBH4DKtO0OTYZfPBMvBzrBhN/QIa/C
QBjlR6X+5bG6Q+q3wB77GXrEQG5zG+Teu1Rgqy6t1vb12f5nW6857sndL7/e5tGC
1RKMdsvroCWeW2DnNs6WCVuOUFqFITRPBNp8syjmeNhEmZKvdbpG+lpaoU0N0RMg
NfWTOrNx9JodAiE38YFdh7N0Ke/S9H3btmvJgDmL6N9sMqWR7OMYKqJS8x6u7L6j
Yd5fYVBoLl9DNjnKaNxvH4g1YWrNE9by0Q7pSi7Kpy4MMzW1qLHeRDI2deuqoCG+
2A9sukZD55AydhtRmwum0kGkMRq7wBzaXRNyJgJoBdV+GzvC5zfve8n2bbhXdeaF
tHKIPjQRai42Xd6bKLpvFGpS72Mx3OQuabtV2iLU5vz65kIQKvMTPITY6sGw+eNW
thkHDqa42wJ8TkOpTVZpRE0AZ2an+vEjBeZF5tl2LGd9DK9HKI2kNuIU+rxijW7G
5iAz+xArBVQsiMoFuxLpC7hjkMBOGLezhkMcCvRLsijZmEbaqMOERdPIoOuajwhm
uc66UJTk0tQCmq7dJfceGl0J7dRJvN7wiwh8BXjmmOMtKPWrBqMlX7QI1vBo7ncm
SuEVejajivWR0qG/dSpcH+4hGaGsno8ZXC+iFYCNWX87NymbTLEZwpH4PQe2Fjhz
36YBvudbZ2/VswCtA3c98cM3rdMV9INEOJ5dYj1v5VbV4NMwLpjZWnp4qN/DgFRw
iX4JVZ/m6JrWcO4bMaQUgfIwXwe8rWTeoEhsOlC48JZmIRng1wIVp4D/TYhJ+NEf
AH+jwEMR01TAd8Lddd8Njk7mXUzPlJhJlp2n69u5looHZ+Uka9BlBa/d9Mu4nNL9
6XpPQIvrWrqKflvbrXDk+uQECQrmf4ElOjjfApettY7wWnV/9enKWkGo1+0AyOYy
ghj6fHn21x7AE5bwNmUlPom2eCbO3+VxPerQIoHGWnzj040pRpIBHzHa/rsj1u1h
wiQp0GBF9ZEZNKZj3nK7gHCJR5bleJ9SiutM7pnd27Wfyf+BJwMG8T39IWWm5e0B
6OLuN5UthsgzkV4Qq7IenUg8Eybs3KKTxmwqbcIUqDBbP7V6B+lq86en/CcvJ5FA
Dp+c2DABTm4eF7Bpq/UjeaJ6lAKb/VSOgF8Mi4fp9ua5DusNS6k3nMbMBr0xYx7u
LNlaRX0cbPC51NrxLU7WSSUFHyfWTgx/wDPilNB7kiyHryfEBE3nOA2+cjaEV2Ac
3Fe5JJWGjthCNoBYNI7T0Y/+CZzwd27y3tQpQmNN2IOMj1f/r+YarvMnqfY/8S+0
uzh3voSiTRsP8ozU9iYkn4cUJoJlKChA8WxgpRuQtrn4lnpsnDhAMxl57vt3Sc9n
iOl0U69x8r+0ROGz+h0S5lzK3Enq7+xVvuQPlwMDlbW/6WzkGkQqeMnPJcxNcGBi
/nJPuGIPECYaBStZuEyg9M9T54sjtOeWxJz3SqZ41PlogLlKfnYZH261D5MwI7NQ
X64s7CWf66GXk/k2Vht8/TzlHeCLTTi/6jWofg4sYfia7DjpbC/T2kX45GzCA0DY
vP8YWrCQxwZhkiegAakwWPj15q42lYm0jU5BZvX994cLTvMzFnL7+3ER3AOCebR1
cp+Ngw+O+EfW60jXA8IUZRul3/0pHFDpNM8DUqx4BaNC5CLzZCnKHy5HG1MuKL7D
dWzheXRTNlBSGjgyxmmzj4+r/6u06Qe/aE28gUeJFMWjeVg1l8TBhWeILUQpjpVT
Q4J3Lt5nMFCsJaSiFWF/JW4VZN+kZQkxWzVPVY/Gaqop6XyFqgbKX8Nqlow6X/sy
SwgzIQwwW+C/QRo8BIkLy5aoDsltaGtnpbIexZpHtfgZmBY52eQmecOyYI7BA30f
G+JcZ46e7RYuQ3euPVbSgMTGXXhz/JKVVjIeLDcDWBHecm6vJTYcajBlqlUif/lY
OuceLYc17V8qngpmJrJfo6H2uUUzOmNmDlJrQKvbqoP3Y8rct8IspAN/ZPfvlFQV
H8N7fECpK2ZWGUpHhQrEOnXtCHhoEQu7y4jJuK8z0UZoVCtVAETaTxJY0HHTICsz
r4740SB6CLHoe4Lr1xCTBQ2qtvWwGfSVMLhw7XQhjExA4sr9Qj/RctDUPASmUaMJ
Ywbs+ndv8cz/46NfqsnSg6uKyXTC+/EdDnzXPr2Vdgy7gELMOV/KrQTKw3+z3NNR
MDdQVttPg5lHi97IJUwvIH2RpNVl/9mc9SXcDiN4OTISuCDQTzy5jmYUqZIgso/e
F18GtR6qb1qvh9wprL15at6riRIXmxTG4aFmBKVviv0YRHRadWbKl5GkZD7Bb3kz
JyA/oa9CFCEKI01xYK1z4H/2YnIkjgLxxU38nichPcDl3uhLc83W2lT8Rda83CDd
e7/g0S/dR313k5PDDvDC5cLT0HucDla1RSAdswVvunjulNxVOVByR3BFyQ0YrFv6
RoIQtOobZGKnjczpoLvNVlg1yStNN7rdJ3PxxNmN/fGlRGZtoH2dv6NVS6mPjC0W
lW7unCI7n8I5B9mF1mo/PUJTm853H3ZB7Kw6akhmx55QfhsdWnhAPxeJ4ed1vlUy
bmBzCrGzVFhd+16rjW/bmWn0oyte5fu2gL6n11Bjso2VWGuzDJn91pSzW+Or6YSC
kTGdd3TgqwaFd9FxpcyOR699HSa/iu610CTyCNE6JYEhsA62A94gPYhAQamf3cdU
yQ429j6IUU9udyKdYrYF5w3gN6D3Q1el0tQxmQJF+Za7N65FYe0THDwarjThJLST
Fusq2PdMCvlWKn07xaqgbxJRPuSU5/tbPXH2LUn/jWkxki8nssJPyUlIuwGGPJ65
ipSxCuPXsd4GIeRt3ww83f8cxDI4+RmOLcVUCEcKeMZxN1xD/AP53s15AFvCBJNT
C9boY/ZZGofUTXqyBtWxONCT5qhPTrX0EVRdhXdLWVadWsyK85TzCv4tgEYyjYBs
r6FOiMfq++spYheWgYm0yWrdzcXOGO78YonArkuoc2NcivY8AebcC/jO6ZnLWmJC
aQWggEbtBKFWF5Bw+OopaEJXButEjhGlNs7CpMP8zcGAB7Uw12bhrN5uM37vy1tO
ub4cD9YYCgghMVra2rF9yxETKtm5GutSn1n3KY9/af5LW/7ep6LQ/M7ei4zY1rNM
Cn/Xv6c1RzaJoBQ5DGxVn1u1Csd0QZRDuNgUHOxJDxpeluS2jz2Puj2zPe7CTZuW
+VxW8B5zWGpCKC101pWS6J73FECREbdycXAJDaRY1d42mFCUNFlIW2f3e6DR/KeY
qFVrwYxcRsiRSlpLOk6KewCwNtW26MP5W63qAI+9G9AG6wFOZcvru3QW8hnbdoaj
xnLkDEg8hHXJdmmVpVYeMXEQ7S6Fzqr7te8RgmKWx8XWYB62ThrmIA3T96KJM+Yq
9KVCn47rtTY7DzfuEgZ/Cl+vx0li3f4drwR+LyDMxxRowHpvZKaKKWPoysHzTUo5
qdFPpMyLP3HCgi4fIJUBQRnGlgY5qgApXbOfzr5QKOFtVDiNYQQFfWlJIL+EGyOe
UXi4jT8Nu++Q+JSfV6Wtt48SIrJrq/b82/2wgt5Tk0+/ZAssEOKCnZYEO+sKrNoK
MCAx271Jnjl4YtGlhtbXNOSmPoGk4qtXPvIGxQpjT4Dn8K4sTqUr5/ldMvJCZfN5
VK6eJ70673/V0KqeIqWg66GHMnb6kjX41Yc00c33YqYTwHlk4AlVf2+hsfGjXx6q
b1TxR7bXBrcEKJq+TzdFTqhzzR8IwA3kilTHKsQN5n9BkMnO4JZ/YHKdvdub9LrE
O0JhrbiuM+NDA6wqYhgCT97K2bIbHiLIMosbm3996/9sLUwyylfh3+4iDvtRNC2J
qTZuRPHKaNm9VBq3sZ4gIwa/lfXMFtktqDO/+SgQ4bvKStXwaxhOrkyDpRY6FhGO
qCACgwJTaVt5i+fViBKDRaCZzS7mX6RG1pHJZcPCFBBxa8CcRtb3i/EwRTQlFEwz
IC8VuOULqeqX+E2DKGyaiucdWoAaSDudeCAD2mTus8e/yqhrvbuf2WyCwDWv1AJ3
CjXRQ3XnjTuoDnK5VGZ0lNbzxKtAZgPovI1ABBj+nwnFTPPT4LXJ6M8GfUbTSYf9
qSOvGfS18ro7PZRSJqUTLBSIXJNgcdjZNzNBuUyLtUbi/L6rkojao14oAGrjXIgx
HdzjTvnvkydkuBE6v+nlfYW+HQYftTOccMe37lhNEv1SJDJfV5reCetBXXx5gdlS
s00VKnB8FR+xVCPMjBwzqemw3x4D6jm/R1KP89KQdjxALvIVCTuCk9cI1u/ORPix
0t8i8b2LUgyhDwTSluTBkRgMJU8PL40SfLqwhnWzX6Bny+Y9Ic42TtjSOHIel66O
jipseocVcWeShvw0CdYUKl3a5iA6vEqU/RpAqsyO401Sk6U7SqiC78F8bBnZH7PV
MtFhpW768xG1gdo+ZEWgry9tbKAhCUdD6gC9EeesoIUjcQp+GDsCae2k79WocnTW
yUaab27wAfP0iI15b4+rFAsJ3qU6DNXtEXkneAnn7q2steGmmzjfJy8gqw8jkKwX
jRaFFrHadV2AZOhCccWCmDd0IqQYORFQlsyvAomQlUN1+hGJxRxXUH9kaDckQO0Z
q4X5my5peuC8U6BvJf3r9N3s6zYEU7kYnskFuqtKxu/WF7eXN3qW3PubLDGwtwvG
Vk5i5tvzAtHKcX8z46pCtXssK9Qt6Igg+AfoQuXUVEKd2+QxDYyIRLEos96w52gK
0WQ8i87TD424UGgydCj0jyzX3AQyvUnfx5RDmczLkbV1Kz7YBhhceUayN959jGXd
oz8BzCOYP/obfex+vuOg1v9bcn5KpnEtgeS7Xk3lKaE4N2afqp15My6tCcn/9J3Y
sbH4WSPO1desCjgXXdUdpws0xLNiSjcu/Prhvr+KMgLAAahQbdnjSrsUjJrlG5ai
9eX4JBGRP/UjDp20LA/tFZsGbFBlXoohMeYibQakwcVW6n9ikYSsXAkUf0uhY8pZ
EEG7dwO/WIJdFcCVqOJm4bev8NBeDfTVYyK1szBjzvvbHiJlGbOUgNEinTN4VRFv
0I1FZFi1anvhdXsXF7j1wfM/HNwj6b18lXTF91yOylSM0Dok0duFBRNYWU7cpte+
4AYspB0T2Hke//O/p6DqOgN6TPjW7+5ac2DAY6tJFLmBXUPVhAf5rGbD+BEfcZQq
IPGzxNnAVfrS29W5MXjjiO4d3m5TvYKe8eZl3rQVxRw120ubHZuOp6vB6N3BuDsF
WnJ5Bm4doqo8zJMO1aAi6+FEEnIaVyAAYcXO/ML6rsAHKtdkP2XfP/sd7gaYHYww
sMZ9SAehhE9tL7DokPgWach80FXAH+I/WKuiOoM8VQ4NeBwudKajgHTgsjH9soj3
IE9uecH3AEtfmko3RCySWkG8hupbAUuMEwzPNHhG463hBUCxDu/O1SjqwNAOiHIz
YyQLwJRNgEwZw92VX1Kn7P5jQ1HMWFXgnjeJTeKZrhckIRizI/D+rbjgJgOi2eC4
i9coYngiEtWYuGp/9M5fD/ngkHjay3+JwafW3WhZfNQZ+CqxlAMW9BS6eN7csHlT
7Ds8gWlplVVvZbI1S4I60O9GtqG3W8KwNL3xu14liMyJWagta/24P78vxZ1/HXUu
sZs4UcSJeVfpghNATQO4jvypa7g3aMxNC/wf4TkGz52bt2d2TPif9qYFYhBa+Ho8
mI+Ff0/QoZ9Ib2voankBLjHk8mLkZ0eRtE0A/12wLnLzDZQ+WsOz8nwB9xECEyi5
tkfj48ZFsfi8BdfsJPa29f5Qy/whBzPtOW6LtD4VP4pYUQtnpODPeBjG5Qhd3ua8
5Lt1FCLKjGT/Ps2efI4DKsUTNI9BC1X2gw4R7C+GX/V1oRofk4NHt7lb/wJSnsaN
bPklC8f3Cno8wonfWHC5qucZW/6zTSA/yWyXLz5N2XIu93n+FeWgACTBnoNv2cF3
gHJsNO8xieGRoLT4deecBDr/OT0FEDOWPKN4Kp9WU9f15beVFUE6zipm15gnygwk
qYmuyW8AekDdvRyiEHc13kOpGcLBkQ+yG1hOAB/2LGz9+L+vf0lAU9smdTkTBOvH
7z1fT2QBpWyTVVJJPT/iAEbokrRLUGN7Il7PgVL1wgMS8bmyovAtjOfPyM0Au+Ni
HVA2Ok7mXcoXRvWXg2HjkzIV+4VCIT3AoFCyVao4XIO7Qbn1RH5Oez3sreVPMTu5
rw/Cozt6af5g7NuQk2vTKZLmVFG33ODauo0S55aFCQl7sFkd98JLNawtHtqxB8dq
f6gtmuqT8aeGuo5ADjDf5VVsvQd5Z5X4cgD8lCVHQbY9DX8VotcO5qPkwtXrW+Bk
eA3xLG+MzMmsazyv1ZFV7U1d5Z8fV0n9ICOY24UI4o8278IHM+kEtANaUjjg/XIw
AknGXyOSgo+Sjk6xh7lu61Zx6NMWj4ZfiQNJ0l0+Kl9ES/3YRlDkG9BknwJEBeOh
8Qutj8KLRAZrTvuJ/lYuDgQDM36SMm0MJJLLp14lxZ20wnt2uNmWC4e/GuilUU+b
mVdG1yUdLyEEu6QiIxZJsh25ND6ltgHZdFz4g0WXoD4vGXH3fSJC0IRUaM3LPoie
IfpABQ1Xl5NPY/Ie+3oLmsIKZISQRTjWKGNeISJZX3/V/Zp+0PHEwrGSSRzgG3Zm
GEdwCqGDrpCrvxuCa0SLKQj7cRwzVJkEmxr9alivlMJIKz+2UdqfeUiiv0FRBbWP
i6OBy26oP3O7GcozfESs7NWQNYrtDm0uNNernSCO71dmypAErKK+5ZMRR/9uehqC
jtFo6uceoLrdyNO344TaRUQ5ECb4T/Moduto4nJAC97NQJG4s57TfdYuNYcESBVp
O4/xqjv9S5l8e3/acSEUdSJIOK22PfHmheybeMF5tDVJnXfzo1SB8rsygQjJm1dP
K8FlUNiaahJWcbAPWxv5BwfSFLuOpGBQW73JSaozCT4UlBK8pdh8EZenJ91PEFjE
UcfYLwRqMUUWFq5trb9O3B6SQJr4QMVIa7Qr+sekzYw8jGn01y+NztmCSh/0+NOs
nGuVka+Zulap8u6BdWstM2GT8pBjGGmO9SCf7FndbQ0TvYrGwZBTgpS+38a2uhmG
pxr6PZS1d3BuqlfqrGhl2Xmu3Q4rfLOEO8kS7zDWImu+sYcQI4t3TpXHmY3bYn18
FDY6P9N5NeT9+NL8kTSEGp6Gsqi3fbZaLfFBvZ0GJpPZ70teIV/lAfWydpThmqsD
RIisz5PwjsJghfdTic//LQztV7KWhvvHAwBsZM3lOKatX6O16uJE06YwWCH0w6K/
e34WI3cSgpvl450Qbs2T5p1+p4cKfQ/SaTtrEbyoydAF3hbgzmAiTWli21mUZPFD
KSIlDS/5s6d8Ymp2g1VCjfPnfGvL//B1DEELQzvLd5zxlwNdauokLkSFJr4RNVqw
4PzOF3Z5iEAc0AQPqkNg45iroHT2NbU/xsiBlop4Z6vA6trYNaBe2ISiuY5cb5R1
ii8HfQzDVGkoPhh35g+R+SNCSOMhSjaoEuFAi9A1yyiljTnEeMmOQ6vtKnIEEppw
yJwe616ewkxSzdUAK8Ybax2NJI9UCVRoS89meBHxbRd7bXUY1qK70PFZrbHa7HD2
eAlB1pge9HLA/NdcimuaPeYl2UuwT2NC754yEYi7sev4EMa1hcNhJTxfklEecMP+
OC9hgD1yZj92lwQH6nxyWwqPnU2la2lL6VEfRQNxCNZT8CAjvZRx7B555mUVCqzF
TCRIncl5H6xyXDbiRQJVZxjaHPsTV5ZSq+8z5ZHYCQdfs+giPTptqYK2ezFeshGM
DiyT2q2yBtPACGm5sxAPc2al9yFEKsxvmBlOY/3wSyfLEvSV+CDu1Wu8TIeEUBRC
9wsM/T390h8T6XHGpzMDRVvIiWFhtkQljOZJuFxoMuEgALuxHE/iZp+4hmPElMd9
ZBU6czO8gwxcAmXakWU/tm1GNKAjugTM84Kx5+KN/PVfxP+RNGE6awqox2ny3fZw
1AAj/6n7/Quzq/F3RI2pKRdQN5f/ay3o+F5mFTMmLkiHeErsE8Fbds9e9xY+Tk3G
ZUQthvWojdwqmHFRsczGuHS/hjIDXmn45jSx0e5SKwhHqXTD7r3/dC54QRx9Vw7z
9J2169wkJQ5iK8DiDDeBZb/9TdviW4KMGjb/Z/t+c4WCpqC7ekrfaalUuolacc4P
F+z2KSpUlMWKp3K2e9N2OQ64gjKL6lCgxzr2wtJOblpHX28idNzv2BLSWg7JedHz
8TKWFR955Q1el4zKVqthCxRmnH5wGZ7qOXcBAXbqDKLrxs1jGiZqxIPWuVgSkG9P
55bhzhtgHohvRB/HeF61baeTsYitkArU51si6pH1ZuU1x4Sna6UZr/cpTNkkHNKf
r6IUeIOqJlgQmBbdHD2C+dCPtIAfM3ZzqJlCm469sbrxWvGs+1IyZ+6Cjj+UAU9c
4QkXmh0hT2WLpPfiRRS8Riq7g3cVFufn93AjaGOuEXR/1G6M+MlgbvZturJNIh+x
Jaf16jXuWoTLePhVeBLug9w17JOuIDhlhCmKrAAZDp//WKtNZLpAC4aXPoO+mftv
ITcbxFmsR5vVEOtz46jpMqmGWuZm8MMdGqdcByM733et6g6Q28lUF15JOPKE/buJ
l+Hsp/dujAIyEtMCKHsBEVMnZmsrPZ06m1p+3L2FfK8ciyi0TGvoE6ZEXhUsr9+A
A6lO37wvLqtkCL02DCbiMCres9ep4u91w/L4gwMXiVHuG3grWxBXNgt32mrVKJiN
UMnHV+uiA9eMQv4zwtHCmDPM75I0NMImbN7KY7SpGYibh97EItwaJKesth6i7AuB
ir1teu/YmubPPKBer9ZroAeSZSSdJ0sFPlNp8mP1DNVd0xvBum0fQtwdmA4XDD4L
Bxuiq8ffKHL1u1oyYzl2WL2ipNFltDMI9VgzYv9J96e5FepMVZE5ROZXw4uWy50p
GeWmtLMZ9kTMFYT09aHHPa3oX73dZSqnIDbmCi6VTyLeUeFcU4ZeD3P5LXPgRq2l
9Rr/L3WmOu753j1Eh5vy4SoywEz8VZJPhp+xlVupB8Tyang24nBlsLNBpgCY7lwR
WZqzw2znMVRUKNjFNJ8I+gI+DQ2ZbpQ26QEX8OVT1vi7cJ1FLTKQ8357dtaYkb/F
dJFI3pSvX53PUTG7zsZBaVpBGoaPrkT3ssvuuZ9FiLVvC0+MiCthwSMykDIwrQ79
mdW2rvpACn3IZjzVDwJ3qMNOfeQFCzzNceDuZfY8DKWsVKQkN2EEdapHd/Bz6Ob0
LwYjg327h0aq9wq1ruR6Hjy88rbL9YA7XeBOBdtu5zKvaOSD1ijP8guhFcgL+rkL
z06LOSYl2/aQCZyk/v1Bjiu28XedOp3piezS5GShZJe3ElST6ay4mFQFjADUUTeb
ipabva1mj+vvQ+mMda3ROZT0h1asZ+Mun7SbDKkAxpKhDueBeRvBt+1DMl6K8THQ
spqVj5EkfasVwsbIpzVgc6/0bu0UGECKRZpmlau2vWc1sdouOzBxWFeNuGysbvWk
tx0zR/nvM2r+ITDiVvb21fC3F12D3Q9OlHBo3oAtbpgAQp/emC5NUEkHo+5aYHyK
a8yrBEvQYwVrB33ruO1b7dxWTJNy5+6v5/W4TXJDIlteFdXBco0KvivG9g8QZQsX
/JvtycENN4E7aS5MWXS+l4a0JbIS7S/g/tT2OA5lCnioOBQJEhkE0Ufovk7lja+Q
OTIgubsuodlgK364yZ8xF2bcSZrJK59jr7oquzDSi9aBjD/GW9WpLn+3uECrtWGv
torMU+sopwn9r+xBljbTCD0fXVPu8rqyPKN2uSkJHwD2vQlqG7E/Rk4xthV9R2Dn
FINPGIBPc16h8F0OTQmt2rFmBi1gYEaucdGTmKTbh5M4z4pcshfm9hO3SFWao32O
I9vG5Ye97SqY2hfxosGqOJpeUj3+p2ngXDtwVEXl5UXVOyikVn8dKqcJIV8kgg3d
hT2dNP4chBV2jLLrjqv0EAfBZYA069j8Ht6uVJcZuiD+MiRWBT2vtYQaBxDDI6Sb
gDyWPW0Ha9mOm/zIUGfc3oZrLmyt5plJ297F8VqvEICjN6dNFFOR84pXQxDLRQYx
A5D29nLNXmg2bd/QqtVW10gJ0OXsbk1nsKHQAe3wpkXeXNUnpOKs8ztnqbr1bpuw
M/i6b+LVMwQtbBiDz1u6bqFcyZaOD4viPoS9XYJxZJYYoIEGjWumOErx8cbKyL3E
No+Ry71WQyK8nTsOgcXJLLMrEo0KfxzYut6mYeLz/SqpR7OLOz7+kJ7sowUaxrfM
MnOLRqkhKZKRKLHX4zlU2NqvlqaFEWSlnEFUz39IYo7JhulMgXxmMfS0+yevwzwy
Lf7mTc1bdvVGvYRkgFkfg/0iYm6HeyulOqLM/U2AFIjk6B6ntN89e5Z2lggXYRmb
MEmlS4ooUpiroz0aDjZnv6K7IlxgYBLLL6KWMX4GvpRWBLFJSmvNUNu7BRZX4L76
FNXVDPBNbh5K4zHLeXQfw+96LpOwP80gmQDZkrtE1irWO2KPcSOh/YSzO7ypQfuM
su2bAnWo5lzk7PzaU7uStxRi8luM9Dk3TDAfy5HrrQhTJk6LsvSorXbi4FNB3guI
Wjx3Gjzhg2VOX7164qZ6hmPQyV/sLI2itXOiGnqPr7Or7/uZeSxzozRTuxBXiUwp
T3TCFYtZ0OZfw7qPVjOeNbdP6TyCtLqZG2TRL33hA3Jd54Fg12zGp/sypW4bqq88
FQc0ulwy3fNBK4MOpyWJqK64cAJGOUC6Ry7L1P0qpY1XXv1Vn31B6Jy30SfWmTho
7c8LAAunnfYokL9XlHjXmcxTsSDH3XEcHhh6UeBiktGFYaqHFow+6n3LQQtetqRO
whz4zIHpojCvnAhDAxL9kC4dfaw3INiuHLA78YFeRZJfxSQrYrDAK81Eez9Sal7T
ROFo4vCveyiRBLBYmRPyQozysMVwsg+rNH6JTe3aBSf7s5TboZBCPoIXI5qprdjf
JIs+AauJcKlwbwuvSt/V/pRza+ExRQggdjR6e4UXX5ueJez1CLcm2UafWjHi/TgP
Jy7yftihnhPAQpiSCtALKl/g5E7F0Ft1N5ApYVlyOxGYkNH3t2Re2SaT0JQta5hp
CpBzPDXV9i3ZvCD2INSmVmVirBGpRVC81Wnz7eoAtK6qmOCToQFCC9/ahEQ8zCWD
aoOdXguynG4HIaIL9NZum5jYS4bLoW+GmqJpTdw7AbUgT47CvryKOwpVghWV5KZx
KMFCqYxdrvYd19bRqjvabqTvQA+k1uUR9Jwi1yv4912X+NSmtKd5No8TvDVOibUD
HL0BSa60m2paI0ndNtD6BlVVTlllzbOs/oAsk2LiunesDMXL/QYDimit4+ZjOPzN
t5AM2iDiczfeZmMftXjwhBaK1dx+ciTbPmu25gGxKNPyR+AtevyPbkr53e38MObg
nnPUMrHfCli4rRCpb2n/hmkPyUy3yC+RSaX6kYgJEICHlBWdbrjf8iwSbxBXOxGk
LYVecgWVBq7VJ9nZefSdH8Gg3s355Hj1FAYMYBAHW2aqJXBtB0Ybhh8rOMovqu31
K7b0+dp93Yk6NIrDBHcU1Zy9Hf6vaoI+tJj74gWgC7YaOoJiYhlJq802AG/1//cO
pKnmV2mnBcgablgZHcCZobTRtCX1nkIbtMFHtMPHQeRVHaxtnnjPyndgSr5VcgvH
qHr+XvIGAziAaiuSvDdYC4YNGk10il+1+pcxySB5dyu5hqbV5SzP0qftScbK4/tJ
oHcTeo+zj6kOBSnnUQBKaqnhOESDX/H33iPM1rzqokMq3UBJeFYTEvP8Dg4rGhAk
gurCOLNIw2zH3/aJqMliu+sWX9tSgESX9lY4Btxr56xo34oUenAYfoEQJEnMosm5
hhVh/JGnDheDPYeTZtpheWZmVsjRwPg9Da+cI3adJz4lNkNYoOEf9MaSrf++8Wns
h6sRlG2kEug1g4/fkpubrQliFxjxwNEsk6j6YWeFemRttTgFuS1HT12zwQBiYcy8
S1zRomsY47ZG8L1j3k7vs/B91r7/6k0SpvZyC2sbHU0mZ0SZgD9Z8s2eCj0+V/7H
b8f1xvfF/yGMFVhBJHZlkahc7mQ1/TLexiKZ48GX1r1QJRxu5OojTevBOTv9Q4PD
g9iKAQ5qMrjYxpjFEMr1Q1bW09yusB1Y8zrQnZWlu4y6noQGdxu+69PtxatWYpYq
dc1JcjqmlvIcVgXmnTm0mGfTWQT6UYJz3HNVoFxJm0OAgF1lIUX4GZthVLZAnn/x
RE6nFUuZv52kx7CvTQ19ap+nK7gIpx7lIi2v3QfF6DhYUE3fTDatwuk08Jitr6GG
lu6qLbe6z5BUp+2kOwxVDEEbV41hkCxzwYeAw3zhqlNBVdwIu6YIegPrgHGf5NpQ
HzFFKDXIQUMTIgthn8puhw0r0/v5zVLRJvsyahZE1/+wpq2QlCHNwWLP8Io0X44b
NpZlYJkLa41KZTA9ZGCt/ZgLz3LlaKDC5pst6YoEjMRA+2j3MwtWhk2rEQflUaUn
Hmp0fABhTN/1gukrdAt9DWdEZrl1MavAXPi2ovisYx7I6VJZqw3wwgKswYJ/+myh
rOVPILKYc8bwxatq7xbC/c02nk6DwVKC0OLEs7v/d59kuqZubI62x1utrXkgkC/N
tb44cD+uikS6KHQXCQliSUCUrDlraIK06zvAx1neVo3EilfYU/Z7mMKkAO2mvZEm
N/hKTku1PMjYWh56yoFtYczmH+Rzgwibhivjoupr8V6nOr8X+2wemtM6WTNEz5FR
QVWTPP9iepw2hvTGgEij8+uzckbY/G2YwJjBvQB8oTkI2Yu53I3qbg8zXp246JqD
sHFq9tvBiQ8+CA5X/vCRDxI+IR9yssAClh3HgUKfWsrx8UDuSjkocB6rGBuneu7+
4816saM98v7Tbnn2pDoE3fmUdR0hK189rk4v3c8BbbGZU34uPaSorpObe8g8W6kg
V01Ei+1YXVvDrafQdBAUq1CLlrHPhYjaGmLJ7BgorY9u5+ccFc9iSfb6slqHwe+m
3EcUsHPISozPADrfnsFbMfQV2kmXMFqEMsSlvv1vlD2YypGM/tscG5j6VtcqqJiT
/GV8F1X81gHZXaCfo0IPdIUXMG70CO6ovoWAAu6GjI9rHACCnMHA1JSJ9HkPCoLj
Nc3AbKoL8jyPq2Pglszbn3PAvt6/Kzl/Tjadc7fB/psuplnGKWzKbOwYIi2o02b/
oTocJrOWLUrpcrBmPyCZBUhMuR39mWOf5fMgt7ZqbdE2s0FKZiqXrFlCVJKsis4m
IZYpqU7Ej6x4tsS/7ILk1VR5fFO/uHJb/u7GGfeZzq5usX7A3NcpOTKZyBx1kFGx
mEe67gE3AUI6X2fmIdCntpcW5PextJrwfa/e6hvtTGH8e5j+XZQFQi9QMtOamltW
Sn4HHPAvOIXmyZEpoa7NifQQR4h4uxcx8NTNlhdOfiAKML8wxbQiMzEWFmc5pRy+
yCZQPCFvqtRJUToOCZz4T4tbXwX4XDGI650WalCunTa9Svg6fhlTCY7dd/bzd4bJ
HLyfrZVPiDEtTTUGKDrh/bNwF6TAszwIODTfpL4kFXBPd/sXzpuENDn+PxDW1YGI
Bq6McUNFifwel2mf3jmRmFBBX6GIH2dF59TGt+DkKVcF4eYKG2fVGWSuzdnF5PDA
TeY9cdF63OKpom36TxDT0SqSaUFftM7ys8KdPYKOtZVhcK28DLuDLK6i4bC67fcy
DR4SY/eMEPYm2xAYwDoeJ8e/dr9mXgmWDjnwkpAVxAFm+yRvzaumA1+rxRZo4KQD
PQrMyrKX1JXLSOb3B8ERXpJ+4dnUtXO//QNb8L0R10suc+4LkPFjPtdMPdpAihvJ
qDM/gjI3uhE7fLox6loXzLMJAXYfQfJvMcPjQ3M+zdffoaaqZ5hiI9CSzpgA1Eyy
0OXCiWouPaFxjJS329Ey2T7DUIEDY5TrODKNuUziPA+jhp3dJGn1ujq1HpD/2Q8+
6Pxf6VKmdGOEWTFO6F4tM/xNzHVzwDrY2pGY4dsGeWT0TjgOnzDeGJQQdLxqc07H
X/MX7SNAUQk6hD/f+0G23YX1BFwQP8aFZUQXQwRymlbIL3hend55Dn5hfGVowqeL
53cvb/onHzci+qBu7ZX4D+4AaKJkEgPXJKlewhuvuoKV9xh0hAktiScPeW4NLD0z
uje3FSVchlXHtCpWB3YJlvKQTDRtxQdzt1XcFEj+FsDFCwetGYFRm9wEdIU7ihyG
wnpJKi69wYNq/Y4Va89/P2v7qf0Cx7oy0B/CW0OMWd+gtIQLCjFyEAajpQeDuC1R
4iO9Rt1mH/8LHlrwtMrPh2F6v8AQAQo3KUN3406LcUnuEKfUegoQPPHiiyLq77+D
iV+2Wh/F40vz7Ey6U5N0z2G3NG3ETPszFWAyOZ6QpgKqh70UudKndOQYLX8362Fx
uecX8NFlzA1xLL8km75c4tH/9cQY61mnSOxaFS0SfuWEK89/jg8a+rnR2za/S1VN
DLvl4VMchEHnf5kwLRYF5lMjhJ+lUM6xYpgsNZ5A8vNXa0W8dmAS5kDcITxKrEa1
+CByT96h0o9oxtqkAoPV8/wszsWkaw60bF81dUhOhmG+swMZFx1Bye4BfBO65nCT
rZfJ62lscQKiIwOzxpa20DvEWLTEpz7uJOHO3pl6lRcYjDS8mm4lTi4roFhuowIK
D9aEw+QwC5eq6KmQcKoicOyGK2FKRPAl2IjOygdiKLOUoT2OKiaJC9iwzY6wHRtD
fqm/POgc36+uTFEnPsGntCyf7qNXEZ6NvjS5D8ufdX2cjN+fNDl9XjhYHd0Lmq6d
ouocFWvXyqEt2E5yVf82eg==
`protect END_PROTECTED
