`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xuOGcpKDxdZmDOnbwOKeauqbdkTCPRTrTplPeHS3CTmH/DkhjEJiVZcsWuj/t27C
YvSm2pMsiUXT/GwNPwnyFoytNmj2/lPhgVwNmTSvXTJ6ucf3ojgMY+HOCI55t9JS
h9x1fntLqWQlUBBZ2MycO1EclkW1w/JT9T4eovRu9GcyrJPeKskjvZi3INaiuOn4
MuC55APxe7P/t63TBmZthGVymRiw6svnLd4Vui0B8joeBIwVslnMpWMzXR40GHA5
6q5pr8Ab1XrFaEDA0lkTRqghfS4OLzjrD2bOcqUKHklljZztYvyvkfake7Y76rat
QBde6xnFBbdx6O/v91Nae5QUTb6b4c7Goo+qcz7fotyhDbeQnh1b8bcM8SC+MfZA
XTzLnhFvlN+S/lslNWQi1InvE3Nb6PH9lmQo7Suf7dLDZJb6MQIN8lEOEB1NIhek
9VqhHttX6bQnY4A2NBZiCJX5zt5F9IJAEBkqaHYtKEdGhCn+F3Y7A4N5HueqbAXt
GQWtiRHw/9w6zsEoRWOU4GDpDj0vzRNaHm4ZijcCu7htFU8S6dUZYlt067qDT0fT
COiQ28MFnmEbpGH5g6N6HcDGi2xh0+6X1VuOPHHDPHJdP2mprl5BYWFqUemMlpks
xOHzNEocTeD+JeGUhO7+R6MvCJx/86P0wTSfpbEzFx4T33yWtQGjie9d7y9aaRqj
6mfKK8zqxJTdh2Oemo1xykRF9pshmIAH/b/QY0I6QJ8QEP+xxkUu/HGx56J2jZoo
Gc3/eduwdkxP2LUsZ4TTR4Np7LKgFm1fPbfsGQaMKO46KvdLZbzfUTHLcCe3O2aP
`protect END_PROTECTED
