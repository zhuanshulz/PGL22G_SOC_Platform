`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
27hHFu4nJxDPJSGYlAuUJFqKqIy8e7/MC7wWWcZRu60CIZoui989NB4JX/8HZg/7
pVtzXJgT9AXe8Lqqd3RfWnZPPWDoBm4znNbOlxI6cCaAAGFR29vHF77WbZHz5F9o
46FhmmucZR3e3l34PhdBYPvM4P924E/T4/ayM4Rh1XgI8wfhNK9VGUvpGftNqb7h
BWP9Yh0uqcFeGcjyeCgGH5wOQCLtJUhXN/SOoUy97hQOEyYbxJh4K4Kug/nnsojt
7H5SeXYHOWsQz7P03JHK3OPwfymA/w2Qlu78H7ba3cnpQEUKwLC1/OnK1o0FUdU+
Wx9Tu/EVybGTuJ1iWbUwhC6BOPZlLkQZA8lxpyiJqnefrU5JLd01kBz7aIp98b9Y
CEszACIgTvWwEDTXcU+kgzyN/wFwNHE23gjkyKTU70dkSxaBDv8Xy7Uc6wgq2i70
Jbnb+VJnzD2RgNnncucMM9Jf2ImK4jk5gxVTzXkqEizUl9qyVfXexSiZxWwYf0BJ
E7PfKM8NpOdyNkiBcBW2zKI29qSblXcI8k+EzTpbFXkD8oopH+UauZ3flSpmW8TM
UbrRvpMoZRAQFfrR9xohTA==
`protect END_PROTECTED
