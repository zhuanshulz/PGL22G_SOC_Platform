`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JsIyAvNjTZHW6P7GBsr9aT9kW3KaacImWHl149Q4wuN2S8xvYocgcDUy0nZQKhE0
7xxo2SIAy2Fl7g5LvOlNmu3dM3DDDX22KIgPeI3aWSDJpN54t0i+ItuDtkPMfhRl
J1tWho92SanimUHc7iqevB5zvpW7MXS2ClOKkhfXPSoL+5wVvMHHW96ibxaRtr0U
TvtLhsg9iXde1h3yWxHMmaRNX+PVlGs6MhvlNFdaOFvpvXejnqGSLISPrqIZ+5uc
I789UsOX+md89uS8P2ejyLy2DCzc5aPKpqTKC/JhUMQgF9E42lqDM/AYhAfYSHF+
XJcYKjKJj7SvcKnpSGNDA0Ncyy2/qNpnRrT8chr7xduWkY/O/W+hHofpXHOshpyD
EcFW5ke7pS7M7l9hHFAt3E3razr+5NbKWS+qUYk4Yq0EYjg4d2VT+hYJ/oCn6FTV
3WJAXVX5U1OmsKp0zio4dQ==
`protect END_PROTECTED
