`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d3xciAFUsuBi3FeLnrhrwMRaRwoQi3SyDe/VrJtH8h+t7qKMGjP4vvamxttNcvIy
kZgow6HD4Tk3zDO8yHwFZYyRil5v5nc85Yp9c8uPWrrPnPmqFW3kEizKD0P2tprT
7xhR0zxuIwNywKwAtLyrZ65R29w+/daYqo9uQoZMhRN49FAWjsmZEQUDNfIbmIFb
x7qWkkAsf4E/j0OG8Qvpca7+IbSs8nWDZ5g7vaMV0hEB5gimpXd6MVG4ktdGXVQN
Zyjry2daL72/5XWCaT2qLL5E/bsUFSgVf2VsY9ORPHmJjzM3lPF0/Hb0iA1Ga9dG
q1kvWVWrW/SBwl0bRINjhr7RWgMa9M7UItERecpVKCx28DDmkJQheysdXyuFuTry
8km+/8gySvOElLhKVt6k5oaHj1P41/IgqFLPcTtHehAFWvTCOGkmmrWdVwJeWRp8
qhZCG4y/aGgdawMoLicsTpbIGI2O5EpOXQKH+rVbofpnI2RDwlvHNh0EhtWT3F8V
XXtb3VnKQFke+mabjkcGTD9CCoIzcxApU5zkLWyuLe0ZVMRCohwpv1qToOmSplEK
NoxN35NEy8rpkU6jQiWrmiO9RnvZVM5RYjUV2lVnsx6PdgF8oejt0w/1Odl0KoN5
IjJqlGkf6dIIb8SN7F8Wh2u4m/G8t/v6j6dgjh/8WV0CvrH8Eh942VRMQKN3sBWX
u7hDUYCZF1bfoXHJFH+/LvR24kJnmuxJzUzfaiITAHsDmSvwSWy9b2+MRDkErZzz
nAYzOebR6F4D3XJRDGnZr2MrEEKdMLmE14Z/QYhlkwCfWvt0jf3ou6139QbMsknG
iwYHyneYS+fyhKI/S6yGn2rhRmKVYW1DiMMMg986E2zstVDvyO82YVqk+S9uCmwo
VHtvlKq28maH2FJJ5ujWieIKLSe6HLBhovMQvx89L77lsZzRjQDefaOg2Aa5MnpK
zQzjsp34yY/neoYEUbfD7N9gR9Ru98dqrSo6YtgyZBZwM6eQ8xIeYv4NnR8BhnjU
MOnrAPj6yP83c1a9pHDv3c/lFjBDcf+WPzXNNTqvn+IDe/u0jm28dVh2Jr6sAUN8
+58WX1g0HYM/1P0yiXxSWkXlGGhKWXMmDoATO74xgeteDk5lmUCLeCr+QenmJegM
kJq6UeHZKKhu9FpPJeSaLOf8JUXkzWYxxuuPp4X1b9uIoXRj3uj9Q0cU1Si9lc0i
zYAYYeq2Hgl5xxc/RKG2L//P/RX018AQ+RBowyxH4k0n3JpoZxlZWgugxqGFL0gx
XmBtbZaq18wzLjUUMzHb/JEGxdv4ulXY78OxAafbzpWaWRaehgqt6hM7UnsyER3c
WEIRj5tAwy7EC4Rjt/URWFu5E8WpRUMVhpssC6Bck3JXqnkjIcQFoag70mdc35Cd
mX7+nFiKrxg7f1WROaH2eL92OuWtPJiXx/3XTuRVyanEzEk48fziko2ZoJVUIMe1
YGESPGpSqn49Z9P3stUzjpmbT2uMrAbZVecdz8VanBiijDl6Hl3n/doqUSIk+yMF
KbCQzyrhd8ErIfo7wp/2DL2NPhmSFOK6WnNZe/qCtjnJSDzf8uCA7PK65p0uZizG
tVzPhupOkd6AxsTEVcz9OFofIVQ9tIHr7YlrjJtRzxSVfgAC44Knn7dqk5gDYq36
3qwqA4qhGfOZl8e3bi0CP6xokP4O2/0fA6CddyFOmkw1Xr46ZTejNGu9Ep4fDsqD
NEZZuM/rx/kWwJLfNaeEYa7beKlcXp/uvcvMSKqRlblfnYrxIQX6ZA/vaoSW+x4t
jdrE5rwIePO8yqkTvEMGDaJpIeJC2zm4PpLfaVuDJBL7RZI+S1AI/47am56U6phM
k4aH/ti/ThBElxMadRE8bw+rYvQekrkLudsMMc2dsm26/lSwkm44n1ChKntmIkf1
gW9WgAODZyOAo/0fzFVqJhjibiV+MR6Je8odgeKFEiSqngvtGVbWViqfBdD2+Lru
TyDKjJ1BSPGi0mfViqvWxjCE4lsWYw+iTaem22EEnHANCGx3tgPtVyFVoDw8J8Ev
BPbJi9rHUM1TVT2nFihnwgkutAqMkQSlWTlnynUIpCcUNASXoZ7P/tjrhdd6t+7C
eVYfN+Fijw0CaylPgsRFR/FTzWuyLPwIGAL/ZzM0H8Lqg1cJQIAKqNaPMyNWJVlA
pdw9n3o9JnEkezpdvMeI8cbxa+VmI8gpxs10xBqie8s=
`protect END_PROTECTED
