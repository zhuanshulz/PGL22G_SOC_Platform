`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O1+zZ3F+iCyFRNHwSTkropaoZz0TGc/OSucqoeH7HwhAP/3tCrNnPVgmf8SwBE3T
DX2VjeNPoiwOt9FQ6UPtN/Uh8hsMCfjhdYeiJ9sxDha6qrzoHRG6rUZk5uHJmksH
XJ6PKULMjZCLTcD85z5FXQxxcK5P9GAvUfujXWfUE7QpYM86Fo1k1yCQ01xCjVwT
Zopwrij03HIypdq+kkBP8+ok6ABNWl/ac7xa2xYOo2BQrnUFy5SaudiP11lvVx2E
zxZ0uxsVSVKfpAZ2UbLAGzmbA/5mftwuBYQD8hP2O6OwZLQIHbYrFQdVHdb2XMNe
KIsBJ+x9f3Q8GoiOzH4vMA6YcspqnvMyvKrfKZUjVbtS1/9dPfJvjiBNmF9doeDF
RpkiKhoyWF4oCTLKbGVaBDhd5ACscxwn4RZ5LJzLz35Vju9ZZUiKRcQC6dK41tky
0RWnPihOvu1HKdlqHc9tooHOmWl2dKnduGWal9jjAEXWCb2Vrn+KIUWVuc5RNlGO
PCaTf+1WsqPMkp9lAS5LMA==
`protect END_PROTECTED
