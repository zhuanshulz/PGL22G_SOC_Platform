`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AD6mb5yWhQGdwe0bHhl7NDJVc21pVmtQtFZU3gzB6NF4e1d8mzkJO2r16k3UyqsA
YZuTNPwBd7D4i7WneluCFjoc0S3l4xy+pquYdIHDMqhb+NFJa/xAeIQxZqmLTw3v
phUjYXFlR5ScKopS8EJHdpMYgAHUoELxyC1fNnr6hGqARkAjJ5Iw3NLJjY+Pg3NM
t/cKs0tlXHScvp882ac9qcWP+FES7R21hCXlBZkbTXUQG6Q0rthjWAzrq9Z0Hy81
8xsIUQtBsAI6Wewi3yPYjxhCgX+o7T+17VLYmhemyA8DNOgtKZ64jD1oks0/zxTX
ClkAegvhB/xyYIGpx2kg65UGxoAmzWG+JLMS9Y77KnKajW5sGWDah/mPJ8w5lb6V
vfxu20Iwags9R5Uj3C96UL+KYSQobTbeVZSG7PKXYHVEax4Yt8TXKAUQ9Tdhqxkm
`protect END_PROTECTED
