`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wAPG4/kuEhRUq7Ec8yvkTIhbnrBThHJnNJ7VOmdLKspVlIEgagWAR+9B9yaSOfBt
1DOEwKfDmfETP0o8RZFLdVLZ7xccuLy+dJexXJjlnwFn90S8/x5PRREys+k7URou
3hQ0Cx8t3F0sRM76Z9vtac6Ewje+DHEMUaQb5wq0vPcy8W74oiu7SZOllot6TPeM
Fzau1g5wUlwm380vSPKXxdgcU7SKYDWLvGxgHASBrimdfX9MecySypMlawN63I4l
0CGDKdrCIEAlPF63kG1KnYWLZTHrlIQIKC8PH1Rv9tt7/XtQQpLqCfnRVOH9RYO9
dc3Ji0AIGZTPQFu/pKqPwKml3INwB9LYnfrjQ8OZnX8/f80ZC6F8cbl1HjgEc4DD
izXygh44/XbiRkbEyBXYfU/H9BrUwUIwH/XWhfGbYVl52Z0pQIJq1HymPCRU0qkV
yXjaWLqn6GZuSxkgHktLB6KWRvDEfHelg5/bzDmZisNyDqELK+OyxKdoaVYlAKjA
1J0beMMAs9fC0EJyXUziJfdoityBBFtMeq+nTLRCws4W7Ew2h/puTpk2StBLX3S/
MvbcyWlW+u3lUU2VuozTtQuWHoV5t7Qon3krKw5M60H+GlpBDTsWQP8wNgBOoOmN
+J+VivmwuDnzJWsKgJYMkdYt954MBnjEDnpxv7V2zdJipazZYBh5Yk8/thKoepdZ
VBXBNBmy5VSoIADEhROrWSg/PKVAQ0cV3QAehstzffHVDrdDMeXteyQB18PD2ucy
NBfczo5rV6tvWQmkuiN0QA==
`protect END_PROTECTED
