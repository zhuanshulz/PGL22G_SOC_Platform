`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ShKzy4Y1m6ni7+XEZX42VG8VO/gZkrR/WxXHSimMWYM7iZl9/MzMbhyNisiGmsdk
YQ4DcBbYU5dYh0nYviAAPh4tFEYnQM5iaRzFqvM9rYeuJVdzaj7L1ejWlzdti2Zw
SEEHlWoD+UoEcCk4PhJwRe52gVoMtxfPngMXVpAB3umRRUMNu271G4dqkl6feApT
C4vQRLFmBFn2/ChY8Zo0waDjWSW+EURkgXY6OL/IvUl1h82q7ivS34VM7VdwcguJ
9keLjipksYRZvJ4yDLbi+ZUMTW0umiayEEh8vy1aIgQj6vGvxuT7E8YTC7PIdusQ
MaEdZhm+l93PmUWzpwEyHtov+Vc4kE83HVIV+iq12qAu/ItbZxr0JVvYuh8oJ36S
AwP1aOF3hP3KAnDIkz4WDKvx0vmDcvqy6rlNNpj+L5aVLzHfiLm+heA4zZA6D6PJ
`protect END_PROTECTED
