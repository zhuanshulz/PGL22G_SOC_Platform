`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fKL9MzoKZbZbJAF2nxVeV+F0Ly52JUUXCjRGgfosZtOmiuhdiDFIuHzNZ3yeRiSY
5zId/aJhjYKqz8oeQhKxSRCM2nNyLYPOyE+ho8X3ZFN94F0RoNOi6HFOFN4oDEP3
eGrt0WwRr26MoX0LQkemffO3sNJBOEB5BYb3/jPl8jFyAjWkVj+npwVv6jvQ714E
r309tJHQUMrM2kZ4+rOXxEFZHy5pwLbF/tcNEumljmRUhAi8merlwxzSFr+giFwW
yHTWAp8QVyqTswFH9CV4jar8jQ1pSVWdfec5qkSjSWQXfM+WmMr77wzfWomf/NW0
himEJ5wvE5LXrcrYkpl29e1t/Ms/9lgA4zrgbYvrn50fNKlxKRYKKJA6AkuKPypw
+FBksVnxhpwxyJYlaoXQDauESpIUAA+7fCcxxy+DJL3uENbWZpcyZvX2NwLCKn/C
AVDY+0k/ZdKsb70foNB3XpHos81i0qTiN6GSnzNo1uGPgaJpVEy+DXN7jJfwyJ/5
GTRPuu90DAzHibldAmQtWBIylu0zBAuLgiddgLmo+RYl9/36t9VUi6dy9Z4bTpF5
0rdaLNyYnCxgAnP9TrmNHJO1H8M64vbODSeKdjYKRQVSL4qgX2t/OppEwmtB7w8r
OzzJhfKgylcFIAJleRWUqmJaS+UXXEkBjcV1WVZUGvLPqhnLm7FfQ4HsQNn6nnJP
gf/T1oifnhEjfajYgSG08448wsFsCxgeRhhqkPS52/YsIRDVSYV4f89HN5WpSLVA
nONwRzSN606hLDDVL7Kw0wtZf0uBbEt+lrE0N0eASFIjlzhzBoZQpV7XTOMc4oM2
Ql2G3Apk5fWZgIiTtTqGb1mWbwkoVsOCelXKwBi6MoCD4cbCjz6Fynl4lAMgpgK8
xjXpzDTQ3Z49fdA94Q/8hZAX/SRNxA+n42Gtl1bD1Ze5ly14NK7JTaxeFYqnc6Fg
T44WvJDTYilaxJMWoo48X6x8EKrZib2YpR/T0HeGfony9qM1ym2p/CBTmfbr4zRI
s+xW01LDyxGQ6PDGSe+x81C1enJNnvrXaWOUhak7psnNGQ349vwHuiz/rthD4Rvv
vDknQgJhcR3FhQ6hF/dtbb+zrQK0FbVf4hE2qxcUXvpkd1mRUXtqmm7+Y6ivM1n4
WCSovDFAHBi35csYzq9teyn0CxHf1iY0wwjFx9bXMULyKQROKGP73TNH2kjbagYh
g8E6NJbeUanYIijPNekIvY+hrTXcqeahnA1kkZfTFqhXE43PvVyf+0kZMIU81pYn
/UiE+eXQ0GpdwF6SFk2wfg==
`protect END_PROTECTED
