`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4P7kKHHRaw0X+20PGWq3gFc5TNqpjxKf9cUM5ZxT7Qolmm6R/fsa8OWg8P/blTvK
v+AOuN5JXxZi0GNi/Sd431wqRWSrUdvkab2uqdVWaFOx1DeUrgh1Lp+8J/sBayQ5
IuOtkBFQE4sPnq0N9PUcMu+fVpXXywjwx6dGYeaA85jOpfVYhHwaJ+KULVa348/w
CCvxMWjmWQZGShG3MOFTakusCQieaX+JuoI1ZdWeJrZHZmlNl/pqOBQy0clsYFxZ
gFuj7DU5gmaX9oAjJlZrLgoBva57l5pwozwIp5GUeAC26c91GDZqdtfujd2tJ5o1
z1XcG+RdU9OSTZym2Nyn1NbT1JPlvLx0UEb2Sq0HqVOAk32dcomY+W8vWeauEJ33
tmG3VyHlVRhSbAMYHRineX6ow9EceDBi3cu1/yiDtvm6SUUI0Lw/8WgyQZCW8Jfk
LWlSUrCDfguaBln1KLiPBYMSdyKdx6m4r9eu9efig5wQDNHomkHWch4iCk5WhHAk
4d5OuTcBevr+mazQZC/ldJGg4MLVPT+NDJZKDY7mgg5d8rcP33Fu7J7TQryQ9vWA
vIZPxYdsSHhhsHdZcjKi5w==
`protect END_PROTECTED
