`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q5Ky8xiE+WZ9zC4QcV1izS+Hhzfp6+tMq9Bi6InzGk8BdxK02YhDh8OHlq3fNoZA
oGh6yCJieTLk9N7WSpXpWHr+TVdKnZ59DF6uDJ++FYBws4XdG4drK3MuxVFKcmcP
YQMiIuJ3FY7ncF0JoASs0/FrAh+vk6RLHpYCD8wxiNTdTS+xMDD7PBf33m8pElwv
6J0QBiMCZGlytfwMz5BvEm1xQa97/6xyJAA5rVq2X9lkyqI5uQnEkxOuquvN27GA
tu5ZQ2ljHlsrKAL/lr+qXG7D9+v6lH0ap4rxQYTc61UoqoyZo9a80Q6zuxu6njhL
OnyWvgMVQkRewv7DiSL0AqZWolAJuxEPwUsnNb+ryw/2wZHATr9I216CVGm4yR0i
4EKmbTC3/bFAU3M7KDPWsSHbMvopNyICnTF1StVkj6gbOjy6gVr4HJtyycmDPkzI
P3Ls5XB6I8dk/B07LL+/7iNFsQnDIGI/xhTdc1xNF8P4Oak5beV8mvV/l8FC62eq
jXNJPqxeSVMfo0ffW+k3vBKK5R9xKzeF6csVHTq1EmkYmM8tsQ+4Kjo9Pa/2XOYa
NH8O4J8rwMFdLiQwn9jbUmSSIwTzIE/GQWFZSZ7p+splug+p8gVfF3dK4pcEVepQ
VXD719JdSzF09nra17H2YPgomd7JevcjVFHfbLOa/ZE7Mnv3eGBvUa2n+IDayCr4
HsZR6wQ6JbxzKwm/ZQA9m9HSzWLlzJ/Bxfmb9HWV0fvFAJLRAUmU+C2u4r21M/k+
Jz1r0lM22CQ30F0H7cj83u5CAIwSaB5Npw9too8L2juS8iep+4lRH5j5WR8m8wFr
jAZHNWl2IphU07P05XNA92Tynp7wKgQBbbOQKkVV1B35c73M1e6uwqEoW/wvlm24
aLfNzOBBKMWRdr1OZgNRzfwYBqojvI2462cMqCcczxV1TkT3Zh50R+cPzn0dlyfl
Epl0UY5Z+VmVJ/M9vJWseQ3GnDEksDKObNqHSemr6CRYXb2UJ23CX9LqVlPnCaxz
VMW8+h4YkK4R3nqI6m9tCV5FIn7bL5/GDoC14ZlSQ7cF9dQGf7ZswxGGyeHesK4Q
kHJ6HPL5YhxHPYfoHxECHQbvkTQruQ0kLF6rWSJDjdWKBTN88RAhL2ucqxb+Iwj0
H/CsXU61x5o3J5c8XfMPCF/onPJ0NHijOhHpy5sHdsha3bZq0y3svhUvtxTmet5s
yk6E+86n+08lITvu68GrQkTN3/gk+zoFCeiLJ3+yJ5PtgzxRrXDCJrFsavepLtYq
np6ZN31gPatKT22EQGpR3cOW9MnVzQESNZYcqVvoKElbrvZAgwxH4Uw1fRUxMPJU
BdHbxosaXQKR/cAUo+6+6lIBXFvmiDf9lmf1OcqfW4gziCIKHhL7inUtSpQv75CP
4IESnMAsW7eFxybjtUqj68VRIZixGaIVE2wtmDGm+woIOQAZPO+ZkfKaNm74txig
1GAJhTwZBPKYMgXWO7NPgZ9ADMbzk7PUBNzP1ZOKmJyha5ht8AR0nF9L5b/E6dL4
pkBO7UnVTnlzmULgq0UEApQj7jPsZ9PkmW6dTvq7u/BYp9rI3vpu1VeGRFByBoHf
rdQfb9qCOgqj0djZigHevbx9oI35lgHPd6mGPRwLAqX2it6EK/F9azrlsd7/76HA
dmolF/PiXPz+a5aTVDPnk88XNsLK2AMW4x8mR+RVqzezXjijnp5NWFEXDua+4heF
xXXielgG1ROyal+7FjaDU/qKPlXYN08Hm87A94UmSoIBDi3E98cG3AIG1eE9TEsl
jS8PKovsq+KZFRfjrLyk/a629Jue2DZxssU3ev9klnody3g/Q8Ykj/QLNFR0Vfyq
/r4qkFSA6gHC5sCHrN2bLDbdeU3iYM9urs/B2oXZ3F3JzCjGIAQMt82opPgXx7CJ
WqLM4+y2oJFlZpWqnr14nUlZJKUd3bR7nWYNLEtNpwPDYOpRAD16QuTsMHj6qk8K
/J0giyB3XcCcLEDMZl+ZOzm0RcYXJYCNT33vqRjkAGfI2GBaEuP/DT4K9BkYJ10d
wBrtVKYNFdv20sSNOiswmveAGjEuZ8pktg0HU7S4FBK1lcGYFdUSQPbV7QV37jcn
B4EJ4aNKL1In3NMDx5rC9EZHuReo9vDn8DSG0aRHDsF4FqbiokjDCCd4WSds9xb0
CMien3xQDq7EAJwfGtzkfFL352Qa4NuZjKA4jroCNB7kqHiHuRG8m40eRgppKS4x
CqYpXScDtKadxoOe3N2yghs5IH5qsQu8mtPGLZa5qHjwEv2qUdbPbZA555ENlAVm
vVBY0hKmpPWFNmfZWah+9QeQADXnwYML8WZFIERSBBg46KHqh+b86TFOXk124EJ8
3dDiqhHhYYeTmC2zZwA1WqLxIr+rtH8S9FlB8sBuWPKiWnMTnI2GS45rGiC5f44S
lLTIfvynrHizpcqTn5qnpO/Q02O86TVc1qOL4FyClG5gvDexWhpmYWTpxPQu8rxG
5DZY2ZySvho1LB8lCN1Jl9V3Dvmxa2JiftuvIOkjHs8J+acijKY145FtHWS4ec2b
IxK70sTR0kecvgmYS10KC3K37nEpZ9SNpUeAcISaJSbsC2HGcHx/sAZVk9WC4Gvw
5ULRKzDnL6D/CBHQyqls8bsJfbzDjmfeJsCdd3SQgQw+clCIuvAM2Kw9egsRJs4Q
I+Rj0Fme4KQQAsZSSgO/fpwJY8TECd0JMvfXcazvM4zY7A2jRTt9gRIamropSKmO
ip2+BH4G+RLRh/S5TLA+mSBlBHLLj0I7f6siCvGiwnVtSSm62gcl2cldzfQyQkZT
r2GvyfM8aQ/PLaByfNNYdEpXogM0tdlOn4wcMgemMeppa82hHNrtrxYjBFQPbLDN
YLe5S+aXbJGInttUvRTvFzn48QYy2p2L70UThf1B+UU0Gtwpx1FWz3UUR7Vun0mk
9vhdpnyrV+xLa1g9D1IXq9yf6dD+q4sunIsJOspAzx9UU5Lj0J4ZLF1eTKMHuusM
Y9FsfWhetIIm3hhSxaB5k3QM/cWOK9DinITxPTbbCpL5kBks/MYHlb6dx+FPBoX1
olnVjpQHaq9q36IzcZG5Idw9RpggJKwi/fXc2LmF/UNDts4wSrlxSQLvryL8XBP3
0Q1s6+Yjdli++8hFW0gm6sJn23/kKDGTLhEEMVevO9Tg+WlNeJNl7MJhXjmiqYXl
ohDylkjWiJ3d+5LFtdeUFAcP99fb4ieN1BKRixZx+66oTk4OZw0qnWvRYHHcA5gw
3W4Aue65NYstXwe8bvG6IVi2pzfuPTNuSzVrKD2o018AOKgJG4p/lP1kVv06P30e
uIUn2WMPsraZMg1O67uhil1qrxR/Od0IkejQa74R57OweG2UQtyM6TDrtOj9pOMb
iuesMdzd1xSfAAgI1CVkszKTxTgd95//ZuEvBnODlpAgxfTCyyugKv1x6zmSBveJ
5oWGKsQReB21fu3H655qJpm68yiKBVH8ZXF2SLn1vdZ0mblonnxQtGuI7Jnf2ASw
ceEzVFJlq2/9CFs22R2g+nCTk7CBatltyVNe0eH8hUdHAUktmQO9rPv8oaVyVmt9
wo+w4Ykp/8kmATXhLtYsjx31AIuKu21iLEYLvSBe13ZhDYs7XPFdlpxmt2y+lFxC
MkCGIi6iEACWXldgG06Jz9ZhPGyJJfqoyG2CJ1nLF5U5yxaOABk1z2rMHVrLRXvz
4sOVnfZTsTuRaWlqMWtGdZO7zM8rDA0e1UpiTr0fBrVcG9DxiMOIYaRaAoTnV+9N
q+bmThyWJzncluDocYTVdcxinAnvkkoRkCTqNHw89tjW2o9RQJJ8hARD5ISrRVKP
SJOr7Ezzt7H0mxABZJ1jdY/tqEoEO2vtt+WKn3ZDU4Wt+NwtXwfcmNQK/EzuUNHR
FCHDOEqZMOulB6LucyFIHTs/dWI6AY1dUeaQVT+BAXTmhk1NJW9jlFOoUx3oKPsZ
8sNcbZ6iAioqTosbzeCRG0SK5e7Uo91bTvBw2CEB7X4E80BcQEZGLJEDQspEotYg
Iax6aiNt5pOrl488nYeP7RwvgqB3u/oZfKSQZS42JTtTU84v9DeIGyo4QwVjG9q7
9gthzUdL/1LWqRrPNVU2tfn2ZQbvBh9gEku3J/TWr6eWPyvVtumhD/drhqjSIAxh
rDMsAeRmzDELzL0fT23LJd+8IVKWK2O8UReT0PFT9uaQTwRxDWtNoAP6hQoj7hXU
gANDIUm74+JisxCpE3z3bFszTquXkfKz+OFHPcTanKuLHA8n1OAYkhtU+heBM+xv
hM2JMmMrwgK6E09qRgOF1sHcDjQjumj8QzxTWcufsWjCQ+94SXM++EbtAex3Rx3G
CU+0TWOikz20WbgxUby3tQKG6XmzwGgkV1vo1lVBT6vTRfLC3KaF0dVwvG+X+m0d
Tx2hPHvPyR9dgUNym0QjCXK/VJn+20PzIPquSjpNL0HOYRC9yFT4oOPAToRUAAZD
3n/42+xY4ZLDqeFf5Xe8lPKZCTrTTBsMWbFK9U0AC2kd5xPAwSFPxsSGX1n4G0wD
cXUjHsfPV6EyieK9M+KHVUS+FcxFb+I3tCJMKOUcPmZGEeEImZuldesIe+8CxF1G
qRk0Q1nrqM7pu7NAYhU/zEaAw8zcdt5t5TjnCDgfAN5Urltv7qSPWiRtZzY5xPZ/
tNP8OuISxcIjlgpREzkj8O5C/3CfEhezWGmXV6kS9/5rqtHrF/QoWf+4ADu9wF20
2rq8ylOROMjfEA5svqWhSgWzDUTDtSc1V4SZS2NAurn0gkyW5f9gEZH/MfS+jS/v
H4YqpNedaOZnn2ODonJ+k/Bg4uBEnczg6Mh4h4ACYD1k1KS57bEFoGZbfvpy2EYN
eW7eDfleu23jiiKI92gGaYV3IPKAHqW2Z0JZn44zCJM4DQ7BVuKbInPZ4qrTON2F
Rn4ZrUbx10pcEerXDa++hRhHxYB2Hw+ZLyqRM2lnMxnFfc48hR7OcS2OpsfzyFKe
D+l8H69znDFBM01jQ4GVrTcNtSfcp4mHu8YLjDyMGAio63dxXLvgJIulw1m0MY0o
nsC3UVrGPeqFD8BbsIF+TJbhospzeQBQMsUFDD1cVVJovvrfCKFTZZIuT2ocMVHJ
YCFk9NhaGuhcEk7whbxxlZQYw9+WqCfuTlB0k3mlbJt3Ckgzv8UbvI1Pnr7mR9v6
/beoIJttEN4CX27/KCfLq7JgUa0cF+FB+RS3KM1sl56F1xSgMlmCSDB40P9BT5Oh
lRU9rcA+PNV69PDyczuVFkV+X7MQI0HJQmMzN0s7Vc5f5vwlTPi932vcVJVkd/BP
cupWEkfIGU+osgLvGltZMZOgh1QerAJNaOhuIacaTxh184cses2p6kzvQ5u6j2KA
jMv8JPQbmIzWdmJcNwz5GL+sUOqizLfKibMImAeGOjFluulN6mMwaohqa+Oudi0K
kg42pAwYV01kJnGGx3xKIoQDdupwSSUsqelFZ8qTzvjjRWRkJt+K1bFomc9THRNj
rtsLCYajHIEpUcJYTCiXN2iSIdm4lGlkJMLcvKU9+68Oa9sg3cSfsmsJ9moeqhT2
6oyXHCAMbaWfNago1zIcJk2jw+ZcnUD6UId31LYyVWcSsrt2Kgy+N2RygKTyqAKV
UFT6tNjSEOqhy6yiug7Ypj7d/g3ieJ1eUU6sA3w9TwshA1EoxA0NO7CHweFpL8Z1
qXbCC9by5EXBc8CnbBtRZvvyefq5tOcD+UF0hpMRmXOxTnbpsmX+RQP4lfUmb5WM
ZoL90J2KjWTII+T7ZPU89lFjjDEjFQhdX6TQ2L+MDAvSHY/CKE5BaJC7j3APysLm
+StcjkNon/lNynp1n7UC6SrLebxSqLBz0CkQOrgw5O+A7DFWOOHWO+VPDBHJmYki
pKi0qHRlyq/je71wssHPNPmfz52iII1CeDnMOt1uGMkOWKshyoAU6ympDfe1NtDr
PcbmYCyEwOXYwNwN0nYo1ZqV1vubBOkQ65Kbmubl1NfdrygwQlazKl9PYWCgMG29
/kZmjXZl5iJ0iD0XUayzTZkgPnIJlyvHxXFkQ7gGN9dqaR2eavX59I85ZTGZ6pii
C2RKPExtCPCDJZZXlekJIeQnBx5e6iLe18U60A6l4H9FcRArHOoKt9Rrb7xnqdrl
4LU06x/DKmNai2TtgETGTk3dSXwdWn6SQFFpR1jPxMEnIoMh2NYzWZpzBR10fOxw
5THWgKit8K9vWkrefIOlcfvhLZAI9raE1nUiD0PJLVx71wSax82sYwKCOtESwfAH
SvvSelNQtuccQFB229bRF3HB+5US2PKmQGjNMImrrO0Xz7/ZkXPjXA6CM9KHwbu9
GpzhFACcxWrlYKNFxNUpBW5SV7mZwiIb4oPaCy8Oy+L+aCHuUz+qPRsSnaKL3S6w
soZOFRboRY0ulxq/hr4eMbC7ykfe9UJbF8W+zkAcifvdcX4MJU78CWWg3+mp4iXZ
qBuohRSJqR2IYjD47GcOTWeMyeNxA7wc9TuqTLvJyhCk0Ws12OvUZOOzxNlzoINY
CaGi2nb1NB9v7bm9WS8YJJOCvIWWok8vUAJwn1H4DpIJrkxIQqbUalqOAtqBV+Xq
cipyvdsMelOir91d1GbWv4Qmv15wRfKByGVa29nUWEumwTqHhswMDZq+TgMFDV38
MV+WGx2PEE2QdH29Ny28xkLhL+5kMQL9nLKLsbDRViBQfuABiWWfpK9yig80m+Kr
mELlItx3rf8ozPtCno+1TlaZxGoJQAdIRkZby9dhxd8pFQC4VbjrstS/c8OCAd+1
YaOvHQ+HfWIMZRZRN0T2q/STOYBrtV2HfIeADX0hkEoVFQ+iPj9O2yN1N4VJE3QX
3/QJnCQzULbUBor1XzjbwTcwpGrG87lRCh8PJbMoXpfGHSxj1Wu42Uwj/3vTMcGk
q7K22BgJy5d05+s+StnC4Zdt4Ux7AlR5kUzNiK8sE1/38E053r05KQ3MFlZ4APu9
otfbZpBsD8BiupvgQgldOeb+X/dgJOumjJrdeoOmIeYRhJLEN1+BszGqbeevY4sD
uDr3XkIB1teJntNNjF6TMYYuSulCjRRpRTovbgy/PqmlvDeUyatEpq3QPoS8Lraw
9lRll+uTvrnyWZLnG2zvi44bHxJyARFtD4gTa7szcHmF24KN2yuOIZpToJTbyBCL
sjKMc2dHeFo05qCBWX6cUy5lc2to4chy8Fqb9PKQKBKZs4L398ekTqLCXyR0yjCo
b0xS9hhkxBhW3YPYl1rdiWGwwxdbdESYm+bBGX7ZaC+Szj964tvY4mK1bjO4ZazR
L+L0MttZqm/hwJSYpXhqu2M7N3MhSXSxK+qtgsdJSkyKgHhZug+pUoERH25cH1ih
+WV2ikGeRP94RbhR5BdE0Fx9ciN5nTK0FUoXmypvtnD7TmiPEdaxq3zE5T7nzLxW
fer5dlyXSTk4ZHdlqcKY6qBQXm8WTA+UP7QBzmWtXBszDMLfDOnzy+plauqy7f7K
jGkI7X51OO19TXd6FiBZ3Rij+vrfemeV7MuWMdK+JamZFT7AzhirePiAyTv8AMj7
LTdZK84IoB+KF+F+YgoHjMu38JiVD4SKRRemlPOQauJzxZZam7YcuJ5eoQeAw24O
XMHj9g6kSU77/xpKhcesVfplNVbJkQTVEfGGhb3coTi+PvfUby43w37cLFHq2oJG
wYyrJMF8VZJdoXaUqc3rSc6mgI/4L+j75qW1K7y+UyK/sGuChmllr44//eETYxY+
sIZmDloJAfWV2woVKouSeuhLHHS8HFux8lwx60B49jrqFAdABttp9hyTwhz+BhN2
0T/S4eiqk0mqoijqztEpUjg++ik/ovsqu53Y757rWQQOCZsOWTf+/Rk4PvxLOUrn
2ai+KT2iRFV6mzHJUwq+lrGCc2BG+GnXOD99HmWUl+fAcvlIKOEyVLU08rSUgqmo
lXb3w58EKWmo4MqFZ/FzaFyTXmSlHZoQnLJqlZBEbkAvlci0one0jKyJQYQ02Lcq
GxYdPRU1LLkHyYZDjVS1KR24iuwuJkGL1np+D7N2vmnweFbSodQ0/TwB1dKZVAzP
QcksV6MaFKS+PXxypbK+GqMQD4c88PDJoEIkAi8OuzDHyk9mW0fo5mzRHCmhnbbx
tDKG/EJkk53+Opeha/Er8/c7HD/45cuPySOshntKL00s8NRc8P+6hfIFHH27jwmT
Tkq8vcuNJU3eFk6OpCrgMPeP8czRrmtdXDc6tQ2tNBkiA4p8rgnlg5p7Ebv27TDG
2yxMLkJ+LiDq/ejNHb25TA9MMw3lxL5mLyeJ0GxcvkQLNA9k2PB8+vOUw6EbRfdz
yPkqSzklCjCcZ5WZVIkkqAZKWRk/dwZrIElqTATrdjWmB69L7UNPRAFt2Y0YJ2Ab
sXkY6XewuWHeBA8iPaqkUqJv8CREUlhMMsUcyVKkOC5aIFfftT0YVQzBC4lhbvzu
R3TzN6jhzTG31qC/aIe0hL4/BaMlVSZ34aAdgj8q2ekr8DvZayDWYorO1PeBfNqr
dSt9wHPyBNFgeoxxdlMoZBOdEXvVSDanGaezNhVhlzB3ar0YKimb1ldF0Slq6l75
VNB8X0VG9xUs9NumeR3q4KbcEtHJU1UQ5sdUSUdlU0Mvwa0BVr8aWme93b4q5JPj
Eb60H+7ibKWt2b0fzvq/K+eUHq0L+ma4Vz5JQkunAoZlfNIHAHml6i1nTSdG32ne
7Da0+G1S5ZvmbTOGQCJRLsfYjTIgeAaKznj6zb2KnLZLdo3xYxWHN1h6WhsEoI4+
WwfJ5subhz8R31o9nVgmwHox3Rn7jjjKlLXPIzXEtaok1T03klG4fX8cATuWdONS
A0C9m88CRDQtcPrKoyBgL8mG1wTk29KttjTNQ0RzeY9oJ3D5s5Gz4sFOEtagRfUa
fsYjlLF0IkzseXmxBr9kyFsq3ai/jRtCiMiNI0PpvERle9SM71aujlso/JRejua6
QNXl+dnSUhguNI198E4i40HbupHtlYenJw5ZM3BtvXB/yc9fLAsuES5A/q9BM468
2Fch/ibCA3EtgUIt+GZJ/0IteVfXIYTpngbeGFSJ1n+WVyHEkJN3fu9CjpO3h5qZ
HwMVOl5m6ixDCgcIwv7PN+xN8pLnWzgtngRBDx+0+sxDH7kL53HhHo7aqYL4WIUq
0xUmjyD9LsZEtbXT9cQNlJ8ouQcFuLwpwiaPAF1BS+E=
`protect END_PROTECTED
