`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OYnhnxyxBnVRruCUy4BF33Q2BVFsyMRz54/hTVudjqYmFaGzmza35wXkHQptWy9K
BwulS4x9GHjbhMYEgqn90HMBmRrenkLHDZtiL6HSNd3Fltyi+42J8ZiQOW9mMJYr
4Y0c1DuWt6Uilx9Bg4/JNpl5626zIcotKNIxxZuhJjLF9WCP3OsMo1Irn6u8xVcM
P69+IMjiPCQFoHS3tMmnUFxZjJGKt32YYOXt7uYk9qBozoVw5CVMO3YR9/MnrFt4
e3gMYr4foGQ4fYNw6713V3HoXroOFV/PYml4TbNA7P6j6JW2E1rIDzs3KCaCOw2/
WVGIL9ezS8eu/N/huEfCdlpPJL0E98uO/ImjI/aELggoSmAXNcIb5T7/5dDiS1dv
87HN1IbJg3C+DODP0f76dxDDvfHKZd+0NXSLrfUkGMxLghH7mwwr07xECIq+QQEc
JCsYoUf/a0W6HdqzBlRG1hGokNdhVR+TmihoUvJTBqX1kyRD86u9MMa3mgKss+E3
EoNDiSguNo1IzZViGmj4J8qLWdM9qT/hAdhgdKGSWhY4P7kEk1A3/upKoGPhLXgi
rsi3K6utCMTxMa0URSFksTGHW/nOXz4vZ6S1h6Y9ONzmQdXmiB6n0/qE01XTxmky
`protect END_PROTECTED
