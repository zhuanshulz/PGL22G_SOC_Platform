`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7RC6CiRWupQo2KG6RMa9OJqfjgx7fr5Tw1hO8BslPRnGU+bNNL+2fhOBbk95HT6F
Bpo+pejt8GCCxbEzoEoSEmvPPB3BYF3791hXIdY1Ou7utNV4AMW3cfWFj35dycyW
7ehBoHSsq02ng41dG6TKrKCa4zPCs3qDJ925XHSjjdfmn7aZ7rxDiIlLS3z62s/2
CSaeaZvZwZX86WvOTesRzOFCzIIUnL7DUxGWFzIqwnumvMJBwnfdj6TXjhIugrVm
NsRGXhtYOqZegLJw01EQyV1Etzritf7PvMJ1elcRPd45tkMDeQxVljBZsAYsNJjg
6tArLCydj0/rHmQk1pUIXaIlJZbD5NCKd/aybNtyWgIdzbTU6NeVeJ+ktbQD0m9k
BXVYUv/qRQ9ATHEQsNKTGETWeSzr0Brhf7iQS2Cni/RjbSg0j92Txa5eqBof16z8
VzHCirkUgIA+VsqSbroKEI0jfUecTWO+CmOQWc7+ybLWXuV4xthW8OjepLpppGUy
QGLVZGF3QT9XyNLh+inZdNZzi9W7ge3bqJf9OkqFeTuIzFtoTM5qQCsIHWaNU7fE
U0CLB155bgx8yFNoV2ZWmkb3jtouCES4D4YWQRoiIIzI8Z7CRUJdaC1ErocggkHY
7pQiIqxZ0aTiZ8fIReoic9qwJcVJ6tpQvEP/mqN3WXoCdbtInLtLR6W2aFIE7uI/
vjD6m0hiee3HSQPbnyoD2vwSxF9GAAqaI/TlbDZT82bxmmewLPn9bG45VXoFx2Ia
xloM7DDEDGfODvZAslnyXRgG2WUcT41F+bbu09ytNxepIz+joa1F9AmnbfJe4wBV
3N0vFryh9myDxCbqXkn3vRKy5ps+RWsX4oRp/2BHmOI=
`protect END_PROTECTED
