`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ubd/ToI5v+JUn0Vij7Y6mouvXZFZTItDaFOS261oqgcDJHuTPnZaLfKpwsiRNKdm
2vc1SaVgOOfUhNxF0o6GC0up7FcSy4RoRiBJwS4NQV4gCWxY9qUYrIVS3OKs49pA
UzyxKJgrWI+n2LG+HmYFCc7TmNsbaNIH/s7ZCpsPqYjwws39nmZBvzBG1h18y1qi
mgV6HEdIah2xpvX6BqbMggwhp3a9nyLRD/TjXYHtYF0cJ2sTJPrTwisce0MSk4M1
2J3lvypWFakqNj+hpjxf/kjPAEgeJwvfQjv58lnS9I3xJxvgOQRYQiVc6t4XZt7K
8gfkJG6nyBM5LlAP7azAD+349E94K3C2Icwws+po3Ti3gW2fkvWOVbyAOzya/KLX
/EW2mfucUVYrQR35I2wtCNwMDT39Sr8uaVt2vQmd03AMjiLpa/yAWNdi0mhs7gxM
cacyZ3A5VU3aQARxzMUmrkW1PdUcsVOEXRNOdgCWDG8uzFJxMZlfi1UXz4q9HgCM
P0pXmQommhsUJ7e00/pBrw==
`protect END_PROTECTED
