`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pO3h4dOk1gwxAowTpNio2sRRMkGEAkrf6XRnU0snSnO+2HSgYTTxJrZDIt5wCEyP
HAW9BI/tr8TMLvQdaWLGi+qboYpGp29ae0vs7o4WiO80nEMnmm3EoJZZzfxBClt7
J/3saN+chiefM7uVNP6bL1WEvauSrbSCcdpjQ5t7Wk0spIHsPORBuh+PePyfw8tm
nZz0goybqzaVb1G0cTHhLwTXMcdt4pTZCouIuWu/Lz4VaUTvM1myQOFsurVsPOZt
1P6kvpCXa7D2lhZcxVhMi/uI/NamFD68wJ268v1mG+n/XfGBjh6WbqkWpnviy2Y6
NuiarZl/nr5HiIOgRJH6RtTdxy+oUVMYvsWnD3avA3dQ4sTVsNKQXaPXaH1SPgZj
4yeZ9hYnkywpVmCSTXgraNXIQ6XgXifgGqAasYb/kmc=
`protect END_PROTECTED
