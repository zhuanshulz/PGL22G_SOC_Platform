`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bD68cEDBDM7skV3IWqxHKrnrpvmGoX8mJ74ypNXOnui5RoHmSSdnxLdtMnbzKWjk
nU6yQdXF9EichEtOmWAlu69cM7vFexo+NfvukDJgKdUXzuYBn1Ej7wVmqJur1LBA
2b+ehWH8P0zBO1cXPcT8Bmyc8Bq+XJRfs9uw5XBPWq+JRv4RmWtUlrksvsPq4Sk3
Oez6Sxhl730Jc7PvVxK1qJlnSnAQBa+TEUZ7MXq3GgSgTAdtbDf+DejLzsq6ONzK
cGx1+8P9HLMIVKhPeLs03T7F9g2gBG5tBwfDQ2ijYjiM2Qb1mYQM2A0JOCYshDpW
JEU1l0TyJAUieD8dx4lwzGzip7JbiuJtITSU7unvBONY0FYSeVR4JZaBFVialH7V
yt57vDY4x5FujQw2R+eCCyco9dyXrx2WEZ/fX/4MuMFlZUQBhoeh9XhLJZQsNHeq
la76XJ5owNcPl/aXkhZZIVjX2MV9GsuKrjdD6IPPNp7VsjMI+YNqvOah8yhn7OZm
hZQZQPcCGZFTcolPPeAeo1vt94ayLjJrGwRcDS18K73/AS6VXB2DGluBoeXjz5uN
9NWqXhi3NRVGgyZGZSFODfR9gUL2X1el/YWHDrj3U5kCm57QBCnDsgTUfKDazO2R
gMxiTkQBEQBkl4ACzSLbrdzcJyXSQhv1TvpW1R8z9zvmWQgn3RF8P6L0tRw/inPZ
ABdeZ4oWhh6bMGX9gL2N7tWMP9XE0kQiB0b9Dv8644lMAQHSp9UYOiA0SOHwdps6
onARNDCxLD0vEvS57SAUHcXj75XQv1YQX95dB6siTC3xyvYgh5F4qqska3sIq95n
QS9cKXWv+Ula5f0LNvMpOohlZwjI5Nn+hJFpPZTxXbwiOcrp5LvGVZ96A6mwny8B
80c3Z45EC7dJIZlQlgplJ23yr50OEol5vpRB7cXdL4MbhhminDJ8kwA7C7Jaea9b
ITvmPAbug/I+RLAFNxQeag==
`protect END_PROTECTED
