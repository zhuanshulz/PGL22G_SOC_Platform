`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8jxt3PNoqCo0IoBtIeXHEav9pUrqGQXAogPS4ajZGQcPGTGBtINuEU1ueP1zgbJY
V1w3mFo+Za1bZTQ8jmSx1YFQ17OAfYrL6O8MWac5BYYJCUXFonYOQbzvxl1YgTnN
Y1xNuPlNfhcu0/KbUe16+oLyPYLzyV6ZS9ddXhu2aXQe3al5OpoBnp5F3WMnexA1
mMJbK5ri9/kLSnTlfz3IrHhxZ0xCLG0r68ErQdpbjqEzAm4qFGxnJcURpdB1JPJZ
Tx+iJsNpagIFith5Sz70HZdCrlUc+wCaDZrvAXV+jYCRIQhs2ywAPqvbXbdT//Mb
vYqajyDJUYjDjFQiWByy7IzS/tFLv5skGMT3IPdkKyurAsiOfPKk0nFe4/DawHnx
GRjNucxy2vyuYnrptOFMkw7ubYk/EYWNPg2jubQD0oniNYSuePy7i1HSx+zM6BJz
kveTWt/TO8Nrxlma1KPPP6k7rFRdvvJfWNdKzYraVOjPpbpp5ncc22+GWNm3JoGb
0EQdN5VCuy/P0x+Fy44gJvi5gWotexUrrouXxbXdeTmJSGoSVmrh9Qmk6AryMW9G
f4VKuoz1LvB3AlLv0QgV6mGO4JKn5jXghNgzH9zfcfKPv2z+Ot8O21v9K4ZPj6Qx
I6WqgUDB1XmutvIpjkYfnLGP5rmO/DBDCDstvJU0CPE=
`protect END_PROTECTED
