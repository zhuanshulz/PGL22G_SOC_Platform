`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F/ncA9g8UueeITKC8qFaMLWzGAeuhmpOzs1Vj9bE4mP3inaqDxoXdmuFMnkUiNDZ
NjLqj0gQvjtIEmWP6BOGm4Vej49oC0P3fODfcvbmOUwrvJF/SYOle6yhowCI3AT8
klpi9TeUPF+nf8OKlqnkFjHuBB2jOvxvG+dsfkrDtGyO9ngQvZI3HD4+TzmSLqOY
w1oVSAJ5kiaRNu8Kae8vjRT8rclgL5MUAzf3CuSI7FB4KjQnfXqT9JHEXZhrO7w8
J9OyIpXog6WSV+U8LhUntyec0E4XJusNgrIEi3j7n9eLwOqTo6E9QCtboEqoOaml
zmTGUqlZwYYPlVTopBDiWmAvUKvCvLi5opJF5y/X5cqLAOXruvRg+P+nbdkO+OP5
ugWzXuJurioGEnk+1ibzeEGrKcVoZJ4PHDHf17m3O+R/TT7yEANzLTJFYqcJOEqV
4RfIfe4mEXWrL/cEl1AwR2pAknjTn5CiFYni+vzUEbHkE6UmVDal5Az/TMreeRta
Vi8/CLYR5d1jJY1mN2qB25Dduzz4q/dwW5YgpiB9prqo4bOG/L9zOXh3zCB7zbdd
HMzlrWtJwZ4QRaDWefVSeOKUsI8UGN2JRrWPJ+wkezxuoKahzmOOgvt33oTlMKGU
E7HBk9LWLykGSYEQb4NWAfLSSq02owRj5jk+TCXVhoKTrHCw/yDObQ4Ha5KCEyFU
46BgKhJDyNZCtwFmz4/x7eiK3dUkWwOJIj8FGjC99kx2gOqlT1hhj0MDooJxKNCc
fnM4H242HRSBz7yLxkIkzxJvnPKfeSAs139p65dvDrvVT0HbshxhTyDah5IWWKKi
ZgBra022Bh2EpRCSfR9imI4wcjX+iR6C27xmWCqkWxjqB0CeBo3RgUmSerG8m1tn
XJwpLMAthHkCZL4ssdOQDTXPR+NYzmGnqD7r90dtKXXAqo8ockJeqIG2OILSRJVF
6IR2sR7F6NYUimdAb5OPLC7HBuu2VT72ZVDdClUF5k8rnU4O1mkOBoONSutHRifc
N9Im0SPprY8SyL0PfCwiaoy47x3aHKWtcyOLVy3d6/bGR+FzpS+dMd7JJ7Buc1p/
JkphrRKH9otdLVYlkMGrVZlZgZQq1coaD0IeI3mzmPfStnY7n7KhzJctkvscijdi
+9nzPKgjcd4jKA6oqJUO+vvpmfIQkYCzYqhvU2B6rP7w5vLkgmjcx/iBPeZ4nFlQ
NqdPLVVflOuNI4I0zBgfgIP/ewTPvR58XRk25qzBFnssuEzIo/w9ZaVY7mOzqtcy
4ukKM9QCEuOxgMYe3L7F5YtVj1J/EKwBsnkipRGu+3IRRdZFmGtfFQiimbc4yC/2
aN8SPISJ/VX3jRJQy/RiFApt7ZObp5f47IXdB/Npn2QwvXlGruiuxil0Dsi3kLH5
E72Y8nC6FW6KXXshUpAVaR68McMKo8C9GTY9roy2hAcD+HHMwrJ/Maxqb9i681Qd
xNdJNZKpDmB/X1URhSgiW977DmRFVz3/OdE3+hH+WW1OzR8VliKR3wYgTts2s8TX
O+6x5u62/QLZ+k1OpkSwnJy10f52gD6QwLdDTDFeeY5gmPTkcEEtO6qT1py2GvPV
w8w+kekyjC21fbL8n1UzynV/badJ++kWannCEvxhAc8hYcJUDoeMESODxDBXSCs7
nJVFWmkdKQ22WC4M/gDJk5HahWIf9/7t35VWJZN0Az2VoKekqya4/7cXOEP+CjPy
fRMnUNb38DUWIi5yHzNLErYg71S7GBjyRy8X8i7r8UCGDrGisIuaR7RYDJYNJdIw
jEOxPaSdhC/FmWfL6/wt/3fItUSXtUQ1+/CIxmev16zPTYgz0VfaBfLsras6rhTT
RO5ffrITMhBOVIwRCwn4ahUrna8upb+maHy4VSKrT0cDPGzov3SAk9t1aVTbcMjG
srE22AHSxCjOazba4KV7h3UBht58Hc1c0YznVBBnGpNZs1iVzQ6yDHqdMJQTkFb1
OHaatgYKDsgJIO1TPcY4NPLm3K2RzEarC+AvTYgpQ0eb6akQF2aQtdeWXRJxgpio
AQ0U2jYFh8sGeMeZkLgk2K/V9NzJ+PMZdzEwXTlLvX3ydcVixvil1YD+6Q3qUh3h
8bLVl3dJVFqMWrjS1R77RMgtEAO383puRErrx2lbZ9WjPM/LroSrr5QFL0DIeI3k
FXVa+T+SxZ8IlYqtpeZELDhRKnJJa5dC5hoy4OI31m5zGT5BWBJAAXYzfWJ85xWj
TG3hLrIlmZG3v8nyuP1mejQB78cbgez6w/P02wJ5xkT77VHgnJ3hoC4vqphRP6R9
Rlv9lU8Nm5xIenQ3rUxkMSfgsaWw+vvFgEJkeHHAJflUimpm9VmPQP1BdSZV46Em
H5QULQZRKGOp0HovWuebq3dsCnf/G3uogwpGyhkBDesflDt/2Eo7gLg/nmFlCS/z
+ZxtR6BlosY0/5D499DfGAxIQ/nF9nXNyMMhlxO50o/aVJrqSBoJVyvVRoXXTmbe
wM92Dljd443sNfBYXMUTHY9BrYJH8Eu0cGlwv3/gCq2GHtPJFqVztwtwNWk6rYVl
0VCyXLXHkMGh7LAo7FAgvuMPZaN2lczF+6oAvkcWNzsO15hqb64FCmc1+2WAyztY
uJq+6Xqx+zw6DyX7uxZRd/UE8hu3bNF64snDDq8S9IK/0+QzvVhKM6zl60WNTg+k
xQMO+KVfdv0/NZY5Ddo/SKYJg7kn950rJa+oLeMtvSLCIBblabr6zt29UJlRC3ee
sBvVqg4MjI0+z+hTqQyCju+nAm4WpPD8XAs25VBhb964JPhSCWe7v9SIi12ydvwP
ZGzSRFPA8K2dc4lDVkK1QQBXnmf/SaMkRsCMiE1jzZZosWoVOJZTzXn57sJg50HT
8vBgtbV4pxd2SJhtE4uKpbfKFfTE5fxxMLRcujyu8R8IS+9YUPFbPA1XlX/8kDHf
ED0Jqow9fiu8m5uriCryJ7kvHyJRCwf7QMwmYFe0i4AlJ0LZs2+t+nFU7ng+1OfC
bMn3QLIFVwGlF/xbm/PzXmCRMULG2nmXmQnf0N9Z//uqWljg6gHn3P7noXwtrKax
HHjyPOKxpRABV33tTVie4xJkEi7+f9m3iiz+fCdq1E9EWa5b3PKwGsVcoCo0/uTA
bxy60ZQ2gqJs60GB6gH9dyt2TQto6i5B4tpYT6POV6W/gR/o3J+LIv15axJod3lZ
iWZ58cozZOhDUyyI8KzpE76wwdIWIDpp3MAax9GNLAR6utZ7Vsxp9Fr+BAc2xCVO
4q+K8HnoY/KZmcFW202V2o58MMMEazfrxVioOw2fAekhIOlxw0IQ/6VUz+4Cxmsr
iIjhpj33cvSEAOAbzTVMx1iUgfR9N+nLMmNT1Nlx+n8dQAldyjaJ4ZzsK0FW5kbX
/tkRyimDYrbZJ4xiIlNfsx8RxGul1ec9iY8ilHFf4siPwLGzJ/eoBp1Sp8+hKbM7
4NphXi22cpKbUnaMJNnFExOs+bb37UQo7RO+Jau9HFx0HaXEpCBnORikAqPDFu2C
lTMgDBw6Ez4w8hljj9p/6diTixa/PPvpL6OUQX2ApT3mH2EXFPS+wa+hFjgA/ZGF
c6Etr/6lJlVfVchww+55pKNX58Xw5Ph++0s6GpQ+LnYzePMyanYsanv4ydgztc+2
OUMhBfTmUcbvSRUdzlkONSdbrA/GYPPXw1qfSeEveXHfUEUOUKJP+AAJxUWxDTuG
sJ3dOj4NG0zppy73q4Ug5A+aqABGHRYOuKIc0JvYeHwj1Juc/DlYbnw9097JLnFX
vyAiU3iI7hm5KYX7hwJDBv89WQynKxNpZKjxvDv2mZGQUK3kjkac/tLlaKstHFwd
H3eGkUHebNwRWdVGzTJlnCsQfycIZtSHVM7UX2Wxf5rU2paICdp/D9/f63ncbtGl
awPY9HXLGGddp4TJX4Q3yVULv+tw14+JJ24BIPZtkra+368SBMN5O9mYhwTQ1EId
lQReetmoHaKOHe1aQ4coqd5aT2MTGDX+vfZV8ot2O/JeBgPbArGyKf9YvEUY6Li8
Lok0IQPNIjIiUtsqvfC+8tRqsWA0s3SIOOgaJR7AHtiFijfW1P2k+N+ycvFE3GB6
bP2aKMNBbnrrVBo/R7YWB9JCeh6OMAHCifMY+ayinG8TPU0Ua4DsrAVLpZ2JRnTM
/ZRxRpSkKgo7RJptaLr4i32jzPpQTNR5SgTl/K+QUhfVbNp+0NtjSLGHTs04g01D
b7/3+SwpDtgOwm8I0oG8gWL3XSyhbWNCw3/fl8tMMFNZ12VezmiWq2d5K6suVx02
FMLAlknOlSCpEsCJRI6vigTRkjy93G+VUe8ud1rY/MyxR1q7VSRrniwfiUFzARA8
4OJqDioapZ3Yiivyc5oqsmrbsNxggaGDPJlg8dJ59uxaHRUnnVmNkSQ4JUXj2XEz
ZbSq7wFTZe0pUyiDbBKK6HU9s5FvfRk4Sro07k+etZOzhc8TXFcGUoa0MMddbMPl
Z5IFD/NIbz3ahmNoItfgyXxjCeTz5Kef2jvr6htndEyulwE6Fav5SM7FJnBFIL+d
cajk7nzQyrMZOkAsjUnBpBImpFOaUTVdK9hgJRDFOB6s4gY8nPGHD0o1SzyKsDhr
SXNtsKWLv0/Wz3xpEYRxfVQg57dzILV28+lbG6T8N3qXVjM2pTUfdDnjkOH4xxxo
COgZViDerwo8bC4pz5RwBWf96WXOav3K/iybVhUhncEjQqhuJZUkeuRPz6/hGOXj
mvHqOVaZFmvDs/5wtSE4a+TI50pwzXf/BvKS0nckxLTV10O1fvKlchysBuObYYDF
peOar/fYMg72QKfj2q2WdFOU9RgoQfjYCfyQjUZnw+k0EW4LTwrjWyzra8tDNrk6
i6Py9oKdL9kLknpdocg9b2hfohjCxRCd4zocxXV1mp8Pacp+w05tES/n1IXzNEyH
sYBPfnr5E8No6JTJySWeYFsHXytmrp60Bywbrcp8oxNeGBRMeEHPtEt1Xm8mSAgD
suLmnpgokzZK0jduv9JtyzEeJ9MfcQWU2UdOhfo7sp1gGsc7TXoWe6ekD+LDJOzb
iC8ssadR65U8fxYUF/bdQOdefkhuvflP4prpitn408lCBU0JqbCaF8ux/qUZ94Hw
7gCrYNgBBI6IYaqAUAA9UQ6owYvrhTZe8m4b043BaR48vhQClxYzBib2iFJ4Gdp5
CpLtA/D2oR4bDnBXDuVERPNQ6kYF2M4ma64MNQKjaGAz72yG/bwkXWN7CwyA1Crp
+tUeHB8X/KDu63B8ozG5A2v6ifGJCC5Ryjl/Uw+aHb6YgASpqX7APKArhOUpFJtq
vkpeyN2+R8ktSBTVkk9F+E1oPyGDDZAOUp3vbiWqY2Rj82Km7ofzFscb2vZBnkSA
rvV/UJMdf7mKOoln3icwd68SlamaKIN08P+33sWdVnhxml0NXelhiKo43vNauH3y
MbF5/i7+qXNjPeLzNkJkCWqgm75bc4JdkF57Gmri/v/O3cKb4AJrbs2Onpk7zxeu
MUtE20ZVhJ3W2Hh0ZaaclVALHwLIzvV8/D9TqGUl53RjDVRuA9SQqNs4VNSy9IV5
DeU6dwSzcCQRHStJW+O1BfQyvZr7Ms6R+jjGQQs1/RXOWqtFL4vnEOooRhnJ/xnt
a6Rl3t78KSnfhTbR8Ym1oXxA01rnOuRNdNqLrALooh8rMnBUCsrdFDsCnbpu2eBj
SFQZDQT17E3CgFPswkjIuBJ7+DuWuaJgZxWxWUXeNq3Mx6uIvrjCzEG3AOQ6WnZr
KmxwfqemBTW2m6/V6FTRmiB9veooMqyfm9ccfsftxS08jhoN8oLxOLj5VfVdjK1r
84cRU+EG5D0mF/tylW7gE/mxuY1eZeFPNlbcZzeZ3SzJTuURCFt4GFqSVgZbg4l4
2N0HNlmNXVovIBEJwIxZdM32C5zseG1uvrSxP6LQIkev7tdqPwm5sQ1P2b+eZbda
Tbnbx7ENGYFFGg7WKKsphNVBI9BfAyI5UUD7+6YXXN7SQQ3vLp1r0ZR2eZvSe8Ax
uUfo7KN8DyYqxtNsiXGHnBB8EELPQbB3a4mLekMp7ggKDgZF0MiU2Dv0DF0WxwMr
UnHHGWQK+zDrVVJnz2Do1gkr+lo+830oTRrAO4tHGF9LNphe/gZQlF/GMb2Peh7a
RjrfhFgMJFPy1LJp8jo9L8KxpB6WcoLxZcI7C1tQO/znabGiGX4BXuNE380p5HE/
TxLGB0SYaI2TQnAmi7DO0G+STkLXWR+La0083oV0EObtjGOyZC5QpnaPehMPRSdd
hTddpBvqn1tEytHzJn+h7lWT7x6Ev2uquORAs6tDVFXdmP1DP0l+YMp863O2TYe1
T1tmwnsBCJE0qZrMVyj8sEh7tLYfgY1kh9biTt5IZ2pe90woHNW9oufwI2cBOte4
WegcCkyBccOKmqIeFq4eWnZMKAFGI5Ve583Do5Aik0nQcl61KXMF7ldllgJlg2vK
KbE8FRmuMvtj3tF+mJsliSpU73rElefvlomahAu0/H7eoRfoqLReQQiGaabJY6Zj
MVfdfritVSUySrSdpeCOE3QT++dzPJ2idEs7fzLP0oMnnNoYCW6PGYBTVb2OMKV/
Bj/v3LetOsksSo9YDdOsZ5BLPdVO7IeDlBxxvyuoBfL+tk8FSy3/XGjhDI6bM9S9
YriNHtHcwFdIRHbCo/XaJS4VJV0nenD+m4iJsKWJVhEonB05rLA6Uf6u4pOSP1fh
poLsb6q+Dl1imd1VcK1XXsbrD7LpMgyChEwFD/Jrka67VA8XLh8fAOuoWcVJ5jpN
mDUMsC0pwH3cXjJK/ziYJMnva4HJa0Z9F+GZb8MN3EouckTQS+Rx7BuFvv8KuCCW
1AfLCq3a6saCd3PKBwIO3eKkPwETK6jBzE92V6fbhJYEPqXkiCmsQL/uuZqFcH2j
hLP+HptGuKMGS+b4YxXJe2gguLLHD0HOAyiIIUNvA1IkUoRXtG0iRMdPnWcNw7Yy
`protect END_PROTECTED
