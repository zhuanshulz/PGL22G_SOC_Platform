`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ouHwFFCl6slkq85WqDTC1FPjvXN3jgkz4UER0S2UpCm+wRItuiVO/AIKiPs8QSdW
ms2rOTDHY1ThP+gbpCFbbgnF5jG2XQWrL0n0h3Xbw/VP/Rqo9JuZM+rd1jrclmQE
1Y36nvWMBFmOfRjUs8H14HshVwcNTfvZ0vJmB3wG0+mmqCxvBxByejnB0Oww/oiX
PBcIgkROSLjBZfC3uJXRqtYiVh2hiqWMI/m+wrl3lzQYaPacjqrYYGd1ubVlzBKR
byoK5EW9tLziq0VEP790BOZ/RUe4PF4hg0/3BHzN0m7qGbRvITnJMfNy6qD1MMwk
YLN4THKSLnDgSwD0RuQvGamz9lPCoFWjhxl233QhPrs9Qr8rxHA3TOFtHR98e5jA
XH97y0yThF5PzObBdarYVsyWpfdhXc+GL8FJ7beNcYkKofjmYtCfnKXbf/K6EFC7
SvcRm7XxKu3Ik5D78QZOeY46kgBIS/jJbpLlY8z1KJk32scb2ls7zixZ9B1CWwZL
`protect END_PROTECTED
