`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+akhMThqO6d2vMnmv4DCMTxzfwNV0MNKD7nr0jfPpYAdvrU7UvRH1VM2bwrXgM6O
fFG8YkBZvMgiYH/UVM02cjFtxqDTo7c7A6LJzoawMOXLJgh62zllCYpcNuuV4imh
f9kL9N1+nHSU9MDlNydyorMxnv+waM1WSC+3tzS5kPOGUnvwNLPFymVclnSbKOEg
/3yyx663vLUwZspSVBeatAwZeZGirHh0cNq8e+WhjwPFc1cTV5tj+gGGT1xfJimU
lKI8tXYhQPPUvheTt4d1s1Sx8NT66x8LZvpMm1tQCFDTOjuk0MRvVw2AQ0Przyjs
MjwIh2EoBPfl4gEiE4Y2LbXKAs4sRLdzOAuB6VDHdMmfxg+PkQigNfyvwcnHkaAD
pDKB0gLX+h5GvJ2xQJ04m0wqHJk6myyb/PcKkLzFqda73SjDVQAjA5q//c8Ukwh3
k9gnjq5uKnm2yGXrQedFde5Kp5j/bhUyyTYj7UbJGHsm5BjeocasrAP6IvdC8B2t
qzmzjJKaI2mQ69wyjWzrtYRZhO5K2zFIkbIufhZQDbQkc9wEO5iRU9s9ClAPl3Zf
thvDyp0batt15vZSoNtRvw==
`protect END_PROTECTED
