`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d4EeflusJt/wMWTSQhpJvVj/6uyqcyh+GJif6KzmZHSA135kPBBPIsX0j/a4rbTx
UDFgG9ktLfIqRDnVeZstLLFWWchv9znhj5ohvdSQLFMZefYeeWKC1WcLn0zzV5By
dg7Fo+3B1xFekLoChUm7tWh9aJvCmiLK//0KozuOfeHt7ijgBJoX6nSAeJL51Uda
aj93pecbw2fO2u8T/L7pFQ3tyHI7NclgD14H+EHKmjjTfaqs2n+S3jJBebtF6JKN
172NcvuUzHMUzU8bEy0teLjXtrtn8XJIztXMTbjTXBvqE/EwNjX74H7CNVSWMDmv
1vpMlE03gPgxl6E0nL738Ms2bTmSAXOof+dD75ECbDW7NPu9ivU9VjSAHrfeMcY+
OhoJIf3tQUY6NYgdN4tcfPj4BdN09fpotWDU2mrQ5JdRopXDiouj9oZyLQ3i9Ty9
uJ1wrmG3DPUnPBn4pbcWp+edEeNsHXKGQDW6dP/5PetVUYqcnsRtj1qIjayOVYWt
wl+38rvAq9BNOmfI+kisVyuG3QXvKLyn5DBkoYvIb2I8+BFx1t9dmWyg+RciO3zr
1ZT5ik5c9l30Df8lDKZmzfyDPt/oeJyCOHfZnBfBZMuAZnZmHQGB0Px9fAdru78F
wLw0oDyKK+H++3BER3s1N/zpoBfTKlZQIV4TVyE0BKxgF58HjDXXl+t4yBR2cS/B
hikwZctbckXz8XtGQpJjT/krTTCAdiWnCP2zTiwOHaRKmFB/XOCieDAZyPQfPlNT
4QD/UxR5UC5Pti63zFcCNa59fvg09LA8kUUvvCJt57g=
`protect END_PROTECTED
