`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Soa4KWA4c+Y+XMjdt/fPnz9GRFf9etPsSH1Q+c+r/1eTqdzGBHv+eHfLyD88W2Io
8/Rx2Fvthf1r8JCI5uD6Si71XCgX2Xb503F6bQT+njN4wcCWwex3/xdwfzzPcR8m
q5LG4GncuNTSdgJxP0PERLEqbNMTaNwOBd4UrSO1Yri0W2HLG4iJuvm3yII43Dox
FvmuKuTYuB54z8iI/smSBlfLe6E6BgEomw/jls2eCxiyX4SWainzvbw1hEpJ4O/3
oOgm2b68Gasw6m53c8syktcpaBZO6le8iSnP4SxNQbmKD8qNR5WTdsLFO19NcJOJ
QGlAa6qTSvBOJWedL5Et50Ib9NZwc66NLe9FKO9YyIpAObwchTyB8F3/ZxFO60Il
`protect END_PROTECTED
