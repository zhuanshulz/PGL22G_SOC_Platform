`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qsq0FBUaGoMrUNa+QyNIil/ni4sivonP6E6Zu0+IYQdIn+kgGDx54EoYgeQ/Gmwv
TnyQdGA5HiDcCbAMTwN1mK4kbVxyofzb+fMhvTwpsO5kHmd3Rt4GKyUkY/w3jo8+
7XhpXxTYn/yBWI10YYWjVqqapnLTZm+68mqOn/hYf3lJdUKqKwt14+NcMRQxBcJr
BhYGt4w4tdIFjfgl8R+dJX0pqRgefALNW7LFp9AQGoYjmR7HuK2jd5mwmi8ghNQr
kadeHqKKmbLv7RaBIYbmy3Bog7la70gTvCAbETMxuYmXfYxfNS6hGc9fT5LC9pe5
/b7ZcpUNt3Ul/0rmMvuXr5qWmyVXoAMhjBA80Sx1uOdl7PEGdrMnCLqESKfsSGWY
e5lH7qbFncdJpeS2runRmvW4eV3JMm/RrszqfD7fn5J2NcanjBC/liucvu6wugxQ
4RaqJMRSS85LF+pj2o+dpTKsGMEVoiMYPazk1pbGPkN+4BHc3TIO36emmMKEBjnC
0BTvtI8Xj1Hi6RA8qlb0LgLNAHcWfBEcmuI4e/UlKVQJMGV0peY2Jfvc+l/kKlGn
otx9dpTlUthevsoeN9SBZaMIFndBxQED3Gy4RlksTdpP/l1sKDqsQKJ2wnhExlME
eBBnZZA2z+dfv33KKiChKKPsgWjo1TtvztNwcmDRqpaRTd8ve/3dTmHTueDXzx+K
TatSTo20GobxIhbyauM3GQZUczCypBGoL4HJppumV5EvD9h3F9u6C3tAMxSTeXYR
JGwNI1o8eJp4zvucnTK4lztmdN0GzWcU/C0ygxgYdPQXexht1cG6eINABJJI8Scq
DajqQKoZvFbX7wTqJ5kjWOuczOS1sSjOsE+cd/4owUprL7gfHU8qCEPtDmvTjmgE
CipazKpNJAPVeP/m51Sa9yN2zrNmpp9jlShzTt5fiS8LYpUcONN39uUtrlrdKeVs
qPysc4W9na6HO75Uen8Ney+QERmyWNEWowVZOxmtXq6sjhtwDM4YPexpm4z1yAof
94rLvC+cIRLYti2BzicnicOgux7qUyzMd7rKvbPG3dDhyH7jpTo/H5bgua4CFPsI
H5LTvEQvyyBH8oM6sguNjRMQ4yDIRKS2xSpIDUt7uA+aB4epeohVSQ9cqnWWSyCP
IYN8oNs0BXSSWc4oJSh/VJMeSFpNt8Vcgg0bfXleicr4fGwa2r0LEs/xjZutOTrc
cJzLhjz2aDVwMhZYoqOyIX7A97477vJ4hauk4fQ6h6lS73AxVpUP0RO8TZQzLLlG
TTJEVCztyN2GvoWDHjgNEhFzjUPnx4Og/OFPm4V7QBxnOD8tM0zvK+JQQEXjvNtp
HSYrsaiQgfoc8Ef3VNqcBGoMzIHFcuLZybyyT6TRRCPBsRZIU3N5vZRUrs1Ep9bS
aZpsLGMHMveMPP7Nfbm+E9bR7CbMw5P/lztsENWCETyTdcQ6/LE6P65PgvE01+kE
Z+jYQ2ARv5fJPlywlUveBh88+RmfZohtWWDcg3ZzHHQH6rERsI1tz+zV5E+VeJCa
awqsSeOfyfBmb/otUNZRi1KqmAe/VcoPz0A6yYN69W7dFAPAxC3ASZ0eo3cVkXhV
Wo0CpadJfotc3II9XpyYFkB5oPETlziFskBB7yvnhbKr2E04JUWedofZUrZWa+/t
raShhftUf1ebOcq3xfuth8HYY5qo5avhOEcS/wjPqgT88AxI3+5Kx4Uk8BXA3va1
kH/kprxrxeavjPhtQX3sndcddOsim/AwrwS4lMss5dku8D2OceJj8zIflJsHXTZ6
30fVejKQsGFpmcJz6jAXCrGldlDFba295oUbArPDuZXdkrmoJXwLzq2qn2fjIhg0
JlEqFOUt7rPx6OJwvbzjBxmVBqChUqeM6xODs0dmSxQY7HPSF4eZBtkdpA1QBpcr
rb007+5wPo/09Zs6qQB3YKnKR0L73hnAsySRx+soergfhQovPCVOdkxDwANz1oz7
0+0fYivPFcXkkePa9vMaraf39ceXh3eH/K7V5ezuh9ZNZQLPPsjBZ8PA4E5H2Yzr
YA0qlnAQeef6TjIP9DdpPN0rn9MPwdhR0QnscmnC74kkkiFa4Xn5hEPtWPaVslk5
tyddyL4sI3Ju7jY98kTFTb9gfYi5Phd8dOhup8LOtyUtLpJ6d34oTvfNo59rzdlc
yOT2AC7Xqs6Vcuc0CmiWzNvIKe1PK9thwndGEKj245hnT5G4MPKkSNkpAP83Lbm4
O4mbodgXuYSEcyXV3didK/Uh11LHyTUBupXDm0PE4B/3Uqv9UQS0ZOmkLwVSwMQl
axEnaMZmpGcUPehA2JW4+OtVFv4iqSqhLo2ZMgsnnF/Na7z8rcb+V1GozJIIvq6A
2ZECgGGaCwsjX6bNRJtI5zm04x9rxeSfNsw9Y1OTKzQaI4h3ytLwPGjxCSX0gEx1
olFjV2UIraUiD1Dc9d9TCcXZ+K9yC85Tj4okJWmghR/sUJm4vsoKfRRUqUF5nVKw
j4HOcaKrMzJvuaADOL3F7V7B1ew5dqhWwThtsT8f2SqhPxi+FS4BhIwjUPM7sJVD
c+p5u9RDpk/qgWCIGcZy0cwhmgfdpxB6S133XmIBunmE3p17XnGmlEtCwat1EAzv
zpnzOeZtTsTAkT5zn1PcUK/Q8d7tDPJ0s9GW/8ZkOF0/HdJBoJS/fam3T4/J5m85
Ps/tu3iDtsLBlnn+hmrAP4tGv/KflgBkjTy0kQvzhQ3quOrCJwPfHVm4erf/Q9la
vtKcs2thIT2ZYNUAkAVqGWyCPOysXR/bl+/A9VMi6t1gNzh+kFuqOJTmpm5wd0g0
iFUO256nEno4sx2V6y1cRpRmny2X401glclcyvtWG696L2oiGD0MaNSXgw59Uejd
qPzJinPLhjm/L14colnMtTcu9wyO6KegvZFRMzfa7ciSlyos4+qFIsDokSZUcYI4
bIkN9RFGzfyVbfyZnAhIaZa3ln7rcBXLx8Q8F78YOU6O1zTHJX+MljlSTbMiEQi/
Fr/jKUl8pGmNrraTSbqLxy0xnt5NudoTd+j8r7Kl0Tvn6prGnhsyLwx18xnD4P32
azJrhE2t4zZqY/x3fGifjBWGCMkXAMDjG9Q8n6iBHlOspHr7hFXi34C3owWy96Dn
9cxAKprUEiCEoPdDSDIjZBkxctLKVcK3oLXxAfXvTQnDrsucpV5rUv5rOrQ6W6qU
4kQ3oa22ov8k9e16PKe0AN+IuIKWQ8aAnMdksTfj8L9S5oFPDQmfQsAKlPNHSs4/
XIp1vlrjCPKBQye7Fwr3r8b5S0bTXJfD15c/UJlR/Ib2eauypAYjgzCedZjHOhX9
Ew2Wd5XaAziC1+M/dGZeKBtc6uCzy1t+iEXOeyUvsiX+6IocjNl4sS9hCqK/eE1W
8RlaS2XieP0U8S9aKuAtNVUYofeYcqFzH7is7o1YVCpdDPDTTnnCuYIsfIjt9RU5
PsOJESgAbk7G5KjRJj+2ERVnjc/WDcYEE2IXV+M3DyFhE+vCv2j/NyJ/whW/VHyM
tApxsr2lCC24FFoyOHNj6QWFcaQOkBesyd5M6nGjcOsekcrALg0v58Re5BW7FpAS
DZT2qkLW9ICrqOtFxdqjbKlYECyBvakgo0/s/C/BMFiFu16pjU3N0uWLVqkPplJ2
OVjW2oWdE4mDGOWqZdkF0tXCH47lACu6BLFbKdsyOS471p5FLhcBUUKtqoRh+RxW
PvJ9njEh+VUMEgcMIYUuE98z+tbTGzmvQtw07OKbK4GYN6CMUIoGHD3KqzQB8+9u
UQl1ow344xjeOFXrJC55T5cyus+KYxRUM7FAa9+22FiS0Pg5o/iUfa8htID+3/5w
sr5gVed/NOoNyamB6Ch/Ile9gQNZk7gqlVD3ZEWtpVLEWyQ5r1h7C6huRt6j3HPa
hvYIi560zvJ1WM4Y0PX37NDkV9kAWJhVJTKvrc8NsFe8f/a0e6yaWVlOQtdgAKIa
Rt4NR+xhP1upTjrWyxnzpceTu2jA+r+zD9lrq2zDNNTNrldqnVgD53fcwX/zJw/2
A4unvS+t33oIQIG8gN1Cvb3TTjXwA0s+M4g538W6xVd6ubNQT5Kk35vp5J53joon
9m3K97EBkABdtyOBkCkPZ19enmKxcPcpKenj8vG2FbP+CBi8SJJGe6poqTq+uQt2
v4gDQLiC/X4tzD41saPINZll+9IWeXdAEsAHy9CwzzXvIqzi9xXXAMoJH6kS653H
yfoJembithIAlhVtm9whTULFPCZeNFS9x+t2XIxE2+vhStkTf3WS3kogCI/ugB8O
QkaUyPEEJGtUGPkIJVbkC0sM687xXQ8DOdv3VrLWynFH+1Wp1bqHc2nQjVGej1t4
pKOkoJFCrx51iS0+hzeNt46KeAanfD9jyr8+RkWWxBfmAc/b/p3p4V3T734uY9e+
Y1nPBxTowlcdNBSlyR6GSVq3OpO+tL6wgatIZotw9OVM43yVie/g00rE04PnFpgT
Ap47mVM/u8pvf3hnx/L7679RrkBdtdUxHnC+Ha2PAXIM/Jgpbo9sjJ/q/MI+WMhl
oqNtV3RIxFUwy9gQBTnlkzAQhe08B8v+AwNg/LWCEBD7kzP17Qn2s0Ol0FE2o88Y
dCt+XaDuvdY0PgcDeV5Y6/3fhYYtUC5UboVNFq9wcn2QMxgtrOWwQO2gYaMVlzpQ
K+99EqvH8I0oyKO/irjLP4hYE/m4YnlqKIO015yhthdfQ0/xF+FnZKncUizowe5g
WiRCxFUC3Do6ZUC3oJi+9yzr4+YaRwgLx6JQSyX+DyNUULGn7a8CDwhd58QrPLaJ
LHYFilLerPp7Mr3LgBOzH7GQoK/vu8T5UCjm9Le9Brpi1gjgrVUFmLVyZ68qB7wr
4VQVdt7DuI1GuyVBSFq/944I8ylrpl2K2f6gkzaAhDxjUzj9ON6qBuYRpjfCAuKZ
t96rN/QikOx9kHrTO7C7nIPNkurgW7ozzv9zDQYriAeqydkAsI7TC2XCEOgNFHdJ
V8MgCA8OhEx1WhieTbZTRHHGhEfJeS5yojdtW86eqQwZm6OJ40+tVU249POByEuS
T2eACywpvEVs7GG5YraAnGwloysGFHsIo7ckoCpv9AVrTvupHJ+o6zVgLD6frm9H
l9bHqSh3L3XDlj9AqLIsA0nvCanpszJYv0QsX6z+D5T5KlMvKxnZHbXM4g9yVxwY
aY/fiFOjfopfwgNso+sm4p9JnohVLiNegr/h929nZJw6gjScuYFwpqYhG3WzMgBP
W4JFKG9+UKOpw7Mz0HmOtG9Yx78uZPRQTOBmcqjCf5M/hZ7fdv5dAD5KqRfD/QMX
JLdcNYrU+GZ1cIJEdJHNoXAzN0jeLslQoDyqupiwK65fBkcczFUWFR9RGaUUuQZl
Bu/QEN/R5lIVZM021rs3eh3keREiVUzIQRWFQz0K7obqBP4oDwBMEr+c6pSE2sXG
RU4guqYB8eM4svWvBHccgAiMb5LvDNH8SADgO234BVsNTArF/h1uzHeP7WS/zyqB
DFNxFdTH1r8imZn6MWwK8+X1D3ZhK1c+azUljMHrc1+HEfOZQCsc1wOSmn8nFGvU
bYg2nysO/h0qr/njltJwcIYJDEXbR239gSIPInwizaXa4uft6f03nzA/Or6aOi8W
lltxbqqoeeI0cZLaP7F0IGeIS2jTxvIdz0BP690JF1coEN/ALdPSP+uMUz4VIee6
VC93DR5XPjojQF0O7HgNbkks381hVkTNHbS7/W/HthVv7rxugI4EhMGntFyaGl7N
NN8lP5FAas76NqupcZx/U1WQlmJqRlHTTQfTbD18teTqWP0wswh0BQYUX4fbr2+j
5D8nxq6CBFPF3ti0TMy0o/Bz063tE/FSkgzGQ0+kMwEXhHh+a2dldWQ00ITlRKvk
f6qJLVQC5bxufNIBzOJ585bJExrBLAQgHd5J4DFczNSZerM8I3xkC7FZkFjv1S6x
+vtQ67kZgei67QYhbIQWrOr6dW+ISEo6Z0Hhi99ASPkOukdYWQoQtltdYUTG0u2H
911WH7dc1TEIDdMMdLgQoEZb5wAX9gghG2PIFxJBuiY7FyDYkRlqYSSaQ2IkRMp3
LuLb4ndoAAXuXDnnaSRMrmjUTAX6rYGRq2InK4+FnYHGtoUDVduqcs8ugDICfNvV
J7M2HUoupGhlfw1nlhSyVVTPtMTZMJKN0GA9x8zz/vsbVUbMmNlvauWi/XWy0WDk
9SMi+TljglROwyaDfpBVi5cloLtTunFalXj4BSTK3KC+pwdjxiccs7EMNWfFyXdZ
l9p71mHsprRPCnaDr4TwbFGScnIbMBFA/qFWZL/6FbI9Rrs8Q7+LRss5ZbcVpcUm
CLxVgJpXJ3uVOxZVJFve4/22eA+z2Crpx9W9wXJmeuSqV2McqWLa8jv8A3o/3GFF
ZODLpY8gZqnZHr3wnh4l92QDJWtrZuQkpVgakrqi+p2UGX3TuYh9jalVhK2u1NDo
a27baBjqGhf8l8BjlHe17sFGb92OaA1KAp6UlD87lqSOYbLLy8X63FulWwyzPd8c
3nfXMH8C7Utxrp8d4j+CxqzGJm3vyc8bnCotrHtkXn0b/3gXkGnTtPoBU2Vlqsix
b9ewzipdQbwe4Zpk90Mw9IlLs6Ks5+jF7+dzi/XfONNyPPUXYgnHj9TzZUBJMeLg
T9TrJ4Kg+Vq7wmVuGOQasfzChohLCxdP2cEQ7E+iLxG8+6oAreV7GyIUa1S5mXbu
Rjd5QwzVOfVANsll8TUOAXlthUJeTh7iTyReJkQCJ5jeQVwEAxwAN3Ba7hQWbZr3
XjgnuVSBuKE1sZtR68J2XlGeQPYccFEx+SnZbNg/pK2srJz2Hs+f/MXN/k6v9O4u
t3oZqvP8uH+++8YJUvQrnpHpsvpIqW4oEVEP1dIfaNC794nLENVJvpwRkkOrcn4K
d8u48UOi7ghMQZi0eUTIm461K46mdyVgfSHSvvxHvSuCGNiFe9WE8m97Pxz52FdJ
kESjM0c3MqmtxJKJ7E8N/tMhMW3ISrPhTWDRBFQmbRezEoeclKAqagQ8BmtsnJrQ
o4ZUXrCC7cCxArdSp6HL+0b6XdaX+ZWwDnJvO5+TNvfyHbyf1o+2lzbMRUO98F9q
dqrda1L6AxdXnlgSt/dsHy5CJz37lqXMO7Y3zt5hXid/PdgPi6AuMEpy7qx6fIoH
N+CAzIy3t/DgmX3WotNKqKhXnyC9Xq2nHTX7x47ubFeHrPAmsluEoPmXpttHkYbh
gimJe+RP58im5umS3u/Ik4D/9KTfVbgAWHzid/d+BYmX0F/7LrDbwgz9PJNV6UgA
xedXeXMCV6Te2zBQJQCQH5vrrEkV+joAMRAbUc2xyXtDZKpTRAGthDDwrersvXLF
0cQJAtfcoDFmBfI0X0hIz69UNGoh2EoHKiGLi+GhblOuInc21pehZyGdCZL+prjJ
qvTp4yTfaOwbAUApN6OOeoGlNHN7dzCc0U+u6mNqa9MBFjDvc0xnbGthynwk5Huu
6lyfphQy7ZmPLykzCR4bY9eyWh5uG3YwMbPKqv8sj4C53c2fprmFDR3FqhlTfnRW
H7sPAwGByDLOQBpp00LzTz8rKl3UNFeTcGObg2ESGyASYxJgm9DTzTF0G9wzk/6x
G5Yf6VRevZHkAGdr0gyOf9Dla9rErdooiq+K645sZXjPbkJoNQrz9XwRCOQ76Pke
S67js0vqUev0015nBWfNx0wTWqf+v27lhiBuwKAruAeLzv3s/O0HGvTmgHSxNBYh
LFYi4GGaAQhBeOOOAsGhxURh/NitKjDFJfKaE6l9z8M590DqMex/Wzi87XGP0BM4
SvfRF45lLX+Bt8vwIkJDMnUE8Qt9Pi/ys5660f62ocx7l7E0kEYbdC8o2mIPtd6z
NiWwR9gN1foj0mRyROwdWvDXLnuo9UyysNXGIFekokp7e6lamULK/Nr3FHY+61V7
a+dzHzRxCP35S6w6sM5E5a6qQHGijGP5vWvwgj0KJaI4Euu7vtrC+pKC6g4R7PHh
YZM4803t897JpftCFV+VSwaZKdqi50TrUf3iXMZZHdf+EUrmDo250CkAbDIlzMiZ
tjIArX/qneU8+CISiqlG7elwwroJr7Fqn4w8jJvwg6bUwsJ6mF2ZnL4W+/Lalt0o
1yNw9nAsN0JdXd9REH9do6tk70K2gy+jZi2XxGMJZ7jbgVAloqni3aVwbNH7OeNT
br0M5HKU94ziRA03yXUbQrZWAKREFmAEtR/Cra+Z2U3nx9KFL55pRjcQvCAAAVVG
f6LrWfmL32/IdPZvA6WgbtBhMbRvLabx+DvUaEtSmNsGU5J1xlvEm28jBS66xudU
amYKrsE+MxH7VLuAP4i4ZH5DjcCPmn1lmClzSJNLqFRRiUtQqdKr230SRCVAEgO/
9MzJRexs/+gC3DvaxqBP3rP557CDvAWLmGDLldMT28MCZPzCM2C8PdOOciiuw7kv
zjZWXJtnsYXs3hC6SZ4Ujp+mywnyG+GDqrRvT5QbW45795h/EerMIgWcXUBdcJj4
bET8nid2NQ0mCX0YYn1a8BRbT9jPyP5WZql/Fs8Cxsji3GqO2TI4AoLl2YR4UHTU
Nlge696Z9dPW7cF7KoUbubys7McgmK4siaNVhEU30zKO8ol8hmaFQlgAEmhTjih9
AHUiW9dYgn7SBW5XYJLFiogb7eYAKYWio29ue6sMv5dsgRYm9xFnAOnwJYqXhuDm
gBJC9MzigwCL3S2Nyv9r6tm+vIjLoJUj0CnKQEBB4OXZ0NX6HDBSIzUhtz4l9sHP
Fsx45/v19RNF7g2LhKYEsb02VpHVPO8Ldn9lAvziOLQ8oZ38tSjd0EjqiTyj7QZ3
lz5kyAAHsX50WLXecSJEG5avbiZqkUFuz9DEmcyR+qNX6L0s0HdN1wPYCYQBFXMn
5pTHuW4QIssM5BjNIrVxA3neNL4/pJWPiOtOjpjrPZoUxWIyD8P7ct67aoM0i1g8
9nWt7Yah+QSb9wMwkfn4t08sp83CeilWKmwlFL4kpseM4axPSU+jbS+mKp8W990s
/WDAkkbp3Ld6gMEykPvF79WUdw9ZWci8bOuSDN6W8cxKUML5hKKMFri2SJZo3Ur7
IUsK0qHpXQAJeW0k7qJSjep16FNrIxr/zasiZZ4vWcdDI41dWoLnd1jYfFa3ujZd
hq2sAxDysnc5fufO76acOj9jW7XpX0h07sP8++QcTTerr6IRLuxS2QNxCMpy/sZN
5F7AZV7K8hmsYO8Vqm4NOxoGQjmxmezbZWyYrpK6Mds2PjHJNf6dvZ9aS2m94h35
BD5B/SQCus3JTB09XjLN/VP9k6bBB2+I1BOFi97sfamkmM7himVeai+kCIHaCyRU
rETRO+9CTUMcyCh2wMPaD1rjjKVqo7EOhZLgJgFqNgHZf3hGtdMWRohx0aPzdTPn
NcIucBLujVRBFh4kA92Smo1aNVaiVfy6NcOcUBCAwyVYFgBrkP9sYees9ZWFxve9
HpiE6/jA+E/1SBVDJBuIO705QTibj2s76FAth41M3rDCtA+CS1SsdZwFb5ikuXVG
lJjwoHrTgzp/mw4uz5SBKEB8qXjUKl3udwIu9CoKA5yKYBRP5STkY8HGTolG9MN6
3DBEKXe3ue1/799if2Q/+ikJU4R3Pi7oRCpaQjGftHlhKWvHhAfnytlepF7LtqMN
vyezZlY7aIU+f2V0IXzr3hf95iW65ze3gqq+nGI8jsKcYu6F1q0lvG+5jkCpuB0F
RF5zmGWKBrmivC+QhaICl7rfNzRl+Hior/gT91E2GdaVeOhUohcHUB/QDrl1p9mY
giL5hYuodZ0GCmuXYeW9Yq8ex9EC1iGvbsrpt/zB2G0wtY3zvwIydgq1kWhZ3LA5
T+qW7sXzNlU5m/Txgp5X4Fwm9mDp6DMhPttM7JefNTBAIZOnqUZl2ARlwrOYoGpQ
i3BF5lXb8nhBAWh8RDG96nV3ymJP09W5rhkkT92rRALVL+u4lE8v+3o5hjN+Ussg
XXYf6zoaNqleXEN+51Ch4wyYhOO3Cfem+uT1t9jx06Nyef9QNKi8nnfRTevOmkEj
QKiBBxIs2cp9gH0XpiNuXlnvf7w2QKR5R4jx3F9JigAcqkrI9lNcnigmWBeltFTW
FKGz0ZA7BlBtsSRAQoQy7xNyIow7Ko17J6hpqWh+FBx8Lc63KtB9cJ+MZSno8e2y
c3zk4TaHt+sWnApaSfJKFsDZRMSF87ngkzSBqBJlgx7xlQSPZoNkmmTovhWAJz0A
oZQAVmjjUx82cSGkK8rjS9r259I8Zv1yE6ARynTr/lzW3LCsXEKd/ViHyzN6cteU
po7NPa1Ri4wVpRHWM200lc5zmcsD+fJeHCHdEkCc0NuBnGA3Y9k74Q4PyTYWlJPp
g3zXhBGcPFpkxSKx6L34+6YDNxqU/wULlD+ygkKYSYUot2PqxJ3FCG6hyIKDQnAv
u+NVBuJwodgdHdGpduNrtnE3l6A2gW5hmALzj5pMuYuh/3QBr7JWhUoCknpxh2jH
9FEZ5fJ0V+lJQihqYgOyHBdkAz52mfASwBzpMqE2eVvuVt3DC02nTODE+ijugmmH
7gtKuIlPSaOFwyqaMNGfchCUPEtMuMDKDG54FauFbcHrf5Ue3reFWF6R9ZY/W8Ao
hKV/v1UBVKvp+Qbv7auLGaXmJsEwo+x+uKvv9z+DdP9/dpWz57iy5ewj5YCgySdl
FxsKyrggloVVc+OkNxjwQfyXUqt8uf7aKnWYjcCuHaPgSik/kffARRPEa3GPOhWY
QkR/tc+JFpzd/zUAupLQjrBGHzE+MMepmw7CuDaDWrDhDdjyWz9D72yaaKbZM9Af
r1dLQJ2HLt3wx+mBEQ7TPFUzsSP1ZlyVm5prXoAyQldAEuTmXY+lvrq19GrE/K6i
o3RuQLcoSl1/J1BZxmC7c1gKKT/OeUX5Lodvp4WVEKjxJzpwYCleUqcBZ1V3Aowb
0A+hzgKVwZR/tPO0TD6slQ+bLgRBiR3nqrP0ubClAV3mk2RtyNviK+3zNUrTO8vX
PPVVNqOqrgIiT7u6Y6YnKqmyTWoX4NHbTyLRO1zNYyQTXba+oDRI+iM/LxdYQfIp
EbD1HcHUtluwYQ1H5InR0VPYJYoyYja5HMH2eJJ4T9468bI22PGnLJ8/J2X0JULu
oCFxH2/W6zHHUYAwYuaXOD0cQS9vwJ6vx8v18qYD7DRFgTANhbMkyNsy0WG35ePf
XcQx4e4G8JKJMmdw9zUa606Z17tFR/SNK7yLU5DeMoZYdmLutKE7s6ylc7EYz4K+
Nbu4C6hgspoCZWuwiFNi9TEQip/UGOyMJasBckqTtX2lhK2JV1rpO+/+AQwqB2fR
WaHI8xFQxZBGQc9dxfqYD5WYIDZ+RMbS2XbDU29xJrgev7wPrRIXujaKdU5MsGQq
EvRj5PUlNcv4sVoGFbddhX1P+jRU6i52xVbLVDQTRzI1tFjCVIggD3MhmW+zzyrK
rZt0LU0VGl+CUjBC/E13GP78bmSEOHCrzM2pXwPZGKRSYZdgJedcxZb1qsrITPBY
CYeBRImJnah8njkKsku2CBjHiNfrx5vzlZWU9zxnix464j9v1BybSpc7clR+IeOY
dJiTM2MJ2/cDR9plNzPaCssw2yU1nNk2k0GvCU9p2ZxMM6+9Bd7cVSTtIdJU8sdk
WjZqDW7kK2WGNSSDe1Qf6snGdb7zcH/0MLywinEeB9SXLKkbBRSBpYg4Hf3nomMe
sDhlZM0w5LK0miVTSO9AkPmAgDNO0jdM9bfijnaD3RrQoprEHCeRTyduLSa+QUS9
noi8FaA3NbbDkTtVTiDVu/fWvyr8bPN6HTW8hThyxkhjBKKrjc02BUKgH/EpVP1m
BYBCUG60lWVN2Kr1Y836le5YTCan+spRimhJ/e/umWIUkfXNi4rXdo0HZ2tNEsqv
mCkkNKEy8NeIZ0nEhUaIU+dIdcsHAlLc5C35lddbTWhmd3m6ZGZlj/xuFjZL7ooo
J903KD7jaLngmiaYx/EopmZnunnoEFKFWBWVxbJEkI6cP8BYVsD0XJVBKsSBVbUP
EIa2+wbr0Rg2FHnRW1TnqzuExoRWa/X7entw9udX5A7XmExKYjw/0Aucm4zehAyI
tVpMwSolLH09MDl4yMRkF49Hl/4BYFUG6fdEtO7SShvq9sVFZxuwhAa9LJRspLUu
F4NKsGSPoOCxhjhwRs20K18GKOADnEDAIgcpFeiDjz25l9J9CtAR/rERiLNifNQ4
zZK3AzDUvLGJ/bJu9ovIwdPTd5lSRR0FNh77il26NC7W7acp6QmYJR9vdpnWnVIR
9Z1HKAH6FNbW8FCdlPfxajsWkKqmqaJS1sUIEbWgM68Wr3UWmZ0XxVqOnS9qoHjp
ykUeiBSI7uJ0N1XQVfw7+GerN7hqf0/onrffnNSmGSDwnA2vpRJ9chQTPWFg7rZd
rYZhCNm+LTEA2Fl5vrnaZSPq8z7RkaMAi3jjyJCdPFmAecQljkSzrsa6ttBN1tG6
wAl6ZE2ICU8+hCQOmcTFIUO+CRSUVAnuMpp4Q0U8jeWC6UC1YOJMNekN5k+IjyoR
rS2O2VdCpFY99mMKmffyfmVPR5bOoj5iqCgi6NtipeuIp7JdhQ60X1H5qaDIVOV+
AkYqDtmFxtVqlnBTHscmnQ/XncZFhJ7th67W2v6OJuUKZ5Lf/5lRCX57g6X1Cykr
tgNkr2nDLjQYNCdI+quJeSJx54zcU0KS3EeTnRl2nuoTyTX3ErZcz+esoG2KrKGW
TJ6sGaQFsuL5Msm+uuDInLOGEGR9CkBrgzqwMYmcGZnF6SmlJ/L5xVYQFu5LUdTY
tR/IElszzuVvHwpjE+qHIdxHzQweXytTczg3ECbiLrMPf5Ovx8lxUcNhrvPM+D3g
2Rs9+le9JF7hd1gW8wWUzEC4XSUGa3Xtw8jQahcOer//wbftFR01KPKzr6WLqeZV
YDPwBFpP4ckpV0nL5O2Xa8X4S5ooBzgv3mXBTVfGQRFSzFZ4ZBPXmjfeerFj3aL5
2iJRwJHc7UT3sqFb/K0KOqVZKIXY6Tb+HpWF55PsgHAEowmcb7H4jh1HHDbP/bhk
IYkKZwRS1XM9Fswq5j3jo+hu8+6zAurCl+e6yM/IRrGUa21GB6FzH/tbFwi0fzEs
02eJxZSHUP8rcaJuk63HaF1hSfMQ7nDN+4zuiAKU1Gp7iTCR6Zue9y5i9LZEpxn2
Fass6Flm/atXUE/YKYHuDNdcgrHpwKRaZAlICkmEOQnUdeaNNXLaYWwJCca8a+bK
cAM2k2LhSe97edEjYToG9gPfnPX3A4cITDf9awcMWJ3nNdpFC16qQujfwtC1vQQL
Sxz7GFFCIpFDzCPfexBZ4Apr1Bro0sa5C2LmOdteHPxTdlkiANghXUxO/QxSYCi5
vmmiWemXMgqydU7Q5QRJ1j+sKC2iDzddF8pissMc7J2QDPJmSI0ofOlJ49nLoyD7
VB6R2K2C3VzjtRfuBtkfCa9Mga3W7tq3UPuPjMZ5j643qCLo5ituKsipPnvH7puU
LvUtOoryJIpWbxCj/6FvdvEw1NPVueUipiCOE0QW+X20U8B5Gs4xD7cgI4wECvHB
4yhIdMZsdH9z8yFQ05UhO4KzwaPXuwucu9hwH6kqMTOUKxOKssOxm9oVYa15xtJD
lV7OTL5n0NSmalJQ+/bwNnD54kw/jV6fwqXF/dC4O09o0eTbNVEXvwhgLzFnJbO8
oTKj6e4nW8El8QAf4h6oS8HEhNAzpuoV6WEsk34mhnVSjZGJTDTffrcfiueFdJ/K
HJK25kUCVcbk3IYD3rcGHuJBG2nX3Dx+bL5BJ0ZNiaW5j8k/o3wnvg4PnNJUGg0z
YCMFdi/ZLcizTvxf5HcRvuqWwS+fol7OEfMu1RGid6HHzqPi5u924rP6RT9TGg1+
f48zXK50MURDX66ez0LLQmw0ZyWN5pnp+QMXjjsSG3sgX1ZjSrzP/xfN0s3LCMwA
uvZtv77PIb4ONFc+CCI2cJo8trETAsxm628SLuOZ/pqzAybsqMXhq5SiOW9BL9ll
uR7VoPteQ9e1jjNGC3xQXVVmYn921a+fZMTPaF42pRf6W9P3JyXDvGC9o12KsEMr
Kdtnd69+6uM5Mh6gt11VTvgtjRRYTGCeyUs2F6BYi5MIJzSFXgi2rTPAaSj81IO8
sf6LQDx17ieXGjL7D5WkEFMEVbgBpQynTjlKEgBEwvrLW9r9gTTxskGZnQ3SyX9w
W8U/u5KRVKFe8zZ5O1UtBAU4PYP+SPejChhaZseX2jeCAJwn4Ef5qvksiAntkDk+
fgzQih7qOgKdyuYJmn0J+h3rpHAgHbPGpYDCR2Bp7kku5ropl+VUYct+zYG5GVD/
SxaBg7DHOg0JwSwX4BzjSRny59Og4bAJWLsYWxcHmOrTlp0PYkRxLSkRMKkzPy8G
Zt9M2vidrh0lihoyrf6cZw5/12jHrSLaj+5klVRTjDmk3wiI/bQ97OP1UyDqgzaG
hOE4Zxu2PNEqvHHPBAkYUUxzVuo9rZPixQCdC8RonRz9MYzvUoZXm2dZJhzJnW3W
9kjBdfL8pnm4z6RiipdGOBtCEbYNFz+fW2hU7CGSOBOgInDa4lm1OJrNSug2Y7Jh
b9Oelg+cloeUsE2mAYa+SlgkzBE2p9WiFmtPrWEjpnhiO/qqEbeXH4bGUAJZ40iU
VemR905fQHrZIPrWYORwDdLSP1oDmDcVGzWmIFiLVbgLwHYcNYvOCFFDOX75qc2a
uvTDM2wpuZb4/maRb7z/ZY4cLTttnTg9v0U6/QwErgbbgVt2quPPC6TC5BdE0W4g
b3uoIa22mzxPxjVcXweGzpni3gn1ytV19hT3YNgjYHq1LXCG7TAMG96EfvXtbYuK
OMcONoS6QcHO5gV6QS5P7h8oBJHCxdJ6HxY9lZObD+o8APZUo8T2LyEb7c6EkPJ1
WViRyCQrZhIDDi3D09zjHfNKtco0S9m7mPZAvTdZ29vXmGVpqr+F2anFwxhcSK9C
pDTgB9t3DizWdOJzUDzbP4m6YTHiqu3mx5Tmzg9T6eT60XQ3IAoWmEvzjL+5cgxc
sBUD24BPek/XKOJMORS+pFurmadmYTsgDkktHIjgP5UQVZs/SqeTRbRdzmulaUZQ
6UTueF7XvXkjubysgdqK6UUZMJX1G25JqbhfXlWmh3MTv7Otcm/nvLQfIBQLq5/3
e2SvSp4x+qz1oO8Caq68wLNhssvly5ZsRH+Wvgjfn/i8RAAa/5FegN8x8U+uyAdy
GvxMJgC/l4AX7+7HCbVSWWtMVoNOQSjIYfVs25lUYmL+cACuDEEzI1VljQowXqM4
mJK6L3W2Nv2n3G7LBDu2NYeb3uXPFNBzTeeqO4seBnnAPugE8HgliPTo1SZBOVUw
1215+LHL4NzU4uDzdP9DoUiowyXBIA63yCTP7o/AKAEUPW3kVS8Tah1QE8Hs5z3c
ifm60SXNosKsiaI48z1L6wXLoa9GeM1uTWoEItWstWWzabrb0UKnai3G+UAXWxhT
SsiCXFe9Zx6bWg4k9pkycoPKZ7BcdeL5guHfbfPApxUY7AhcdWy8oU95l4AExtj5
dEiNskyx/xSNJ9AISrwASFwCR1RiUzJJvYBOzW69NTeGGQUJgt9gTBVQvEc3cXmB
VWIUWs/QjVdcRFcqJW1hdxer6VDxu8f1SaBeqqDoSEUdE1pkIMnt6jAXyXYF7+Bq
1udi121U68rlD0BI/ocTY2KhwXpV1L0GXP8SGHbLLEamAXgI3xrGRaH9OpMgVUPx
UXZWR1iYxQuqYUn8T2MvdEyUHCceD/eWZEsh6i85zbsc/XHcJ5gUhIjdGhTknnpT
xutNTtN6+2/sBxrtxbmConHVmsW9Im/Dlf7aXfEo9xo/cCLva1C8/e1tzMlKKLIC
C/9BSK1OXs3zQXSTmZ3U/RAMpRLq36K7XqmREJM+jol3NyryoNN0iq/HuBvtnef1
0dOIFEXEy8caaptmi4CiJb/wkUqI2saXwJ1BzNnVAheHgRGG2NwbnJOjhgMv7vwe
fk4jfme4XWNdpe1dp0+oE7KPRqwtybgmYC5j8xJf+OxskzwCXGH7Nci/4mu5D4mp
1sYXf3kTKLi7NreE1EhZQPdH8qwrobWn3ZlFEaUr+LavdHGpMs3djch2DC5eCCw4
EvGs17C+Prm+nMYlJIUvMyI0IFxvTjhzVnHKWrhjhkXj96POxWLD1ika3uQf9HrV
KAbGJHgVojh2GGFOmrkjljbkr055tD522eP8uNjvtJ4iBz+scmUNbburbquEeNJ2
fXGEDWPAv3MRVIhGeRMLpR8lkidW/MQLHMe8xI2UuN45jY06qmUJlwc6OX/ImKAn
bRntUMVD0frnIWi4InfkAewaxbCjm1VaUlzlvP5OnO5W+5FPd/YXfRzb0ufwpEnL
OMg/QpmLksB95EL6YV9MCDKg4R5r5GfwQSt5rVtGbbpEEXbFwl3kFrmaIzr+uqCM
ZAV6XvlRNy1eCOVFiQXMqv3HS/KHJyR1le/hNJZJf0jHrtYnldnwynmbuiFeMT02
K9tNmtUN4SXQ0y/KnU/g60Faw3bQIqoo7grcOVsoBr2eNFC3JDqI3lJNkRdO/fN2
VxTyyojKzlXzE5T1208kq3SFO867dPaaM6Zh5v7K8+6wbqSwJ3wZXsIv0up30nf9
aoaWW+rMBoTTt/DeLeC0J6IkEdIQItjDj99Ww64Cr0ekeFV0+MjcTASEvgHJyRaw
7X0MgUUP1k3QNAzPTIWvS56WhSvDpQPJbrVvdPTpIJoH3QO8A/R4a/rkszOP0EII
AtqyGiIL1+aFtX1CGkuiHVoieYa30939BdoAD1BvjiaZwT88qlRZvn82Egdn+Y23
flqbz4eoqIAnXpPCWDSMpubd/omVu4pk4QEB5fh/AUcMfRv8mDDbml3FbOroNnSE
ebGrL4czSTHi0Mri/E43LI28b/T4FbupGyaDXyikPi1HIMP3avDo1eyfki4tvLNv
W3nwjqibd5zGOz/kifLAk7T5/iIR6B3pKw3O8cqovzmPSqWXQdKdgs/8ecioKmpR
nnF44KLkJjOiZfwvgu1IqteT1Fh1xXeJyx7aVS+PhDYt/EJDleEJ3bbL6QcRFnzY
YVonDwZZYSS3ISP14uMmaBcqQ+UyWl4bzEc2PyYhCqFGBbbH7C9QkeIlfqqElMp3
9GvQg2oXGh82Qok03oc5F9dkv4Kq3tGZInKs/gmGraG8nmXhV94sOKvmLGK6aYIV
Ohe82No07Fo2w3afersnhWy/TDdzrb65fx4vsD5zGAoh7bTw0zPunH4fLNYmHyV6
wfRl5LJuvfXSbe/b7GLWKT/Xg7CFY5DJHjBLizai40p2p/X1Vsr3o2Jxh5PZvRVW
cAgZ6sGAFYUTIHHgWm4rJsDft2kLDE67hFM7Tuf57+l6095oUoZ4JylTFjPcWRr/
IycR1HUMkrtj1tWQUIaT76NaJyk2efb2BD6ETYnGJIm4nYShqRTy9Eqc2LrpBZIs
RWPvY55+HjaayapzXPyvZIGLvO083kwSdXxmwpe0MnakisAtrLLSxZGWvpcYF+po
r2ZrwSS1UcO+lPbyxIPU4rlP/mkNBiaunJ+TH5G18uJWaY1gcwsPRi94DIVnef99
XQuPPnjMobfVFXFv0IN/p3cTPlAuYO4WUiGyGST1lnBI8pi8HpfZhG+bKRk6bPZ8
pP7iS5MJwafGjGCOIf0lqRefOd8tpWNrW9lzDr4eMYtF5GIJOPzNVnuW+YqDSuis
u7X1QjrtkDAOoZ7O23RtFdUiFM6qcr7TLd2rJNUGjJzZ0LppXHCHlOUryKCwdp2g
auRryNtYH0ii2qU2nzQn5p87E4ogRoPKfw5WQkg4P+6fstOUHlJhY4CdyBkRs7Iu
NqPq0vM2ik9AO/NueIz8Zb2bgItzqsUIH4xwtQJ1VT+ZBsD/XuAJ32EmfMn4KNlp
wJ0FDLHZbQPLCjFb8WeG4agWDuOHYkuJtfvS/gMd0zyHcFpRM4eOeGzq6+5I1WLJ
yX7eZ+YCE8lzcQKtboXaj/M26OvV34GQzO/RFpETg9CjcQFzYDIdkIPDqOYyUEJ9
nwYEDaG72nZ1KniWQ/CQUUOkB12wdmsOb2avHdTkKRIglwsRpBYfQzHA2x97FZQY
io+ICB9ejaeTrPPvW9OOaFAc5JaD4GULuB8CNqvUCQMwEohOrGr4jPp6sjerZQqr
EKZ/LAKdX6Td0+ASP3rwlyC+I+z+AWQ1Jsb6zL18q8yfQYEX0ugEHf4Ki9cmamzE
3GHCE4BGs7t2Yx0VZE8NxmSTWRar7QU+T7/K58AKFKBu2gyEEDgYDmJ9/H7WTYzV
0Hgo0bgOSTYW9ZVxer80rlwtdhDXtemEXE77rE9cELtE6OJSFAK62RLpSOxcLvLx
Gnl+mBv0RNhw6lWl6KdMfLydVHyJnYNMwj+/U/tK67CvUJ+TaFbCLwH3z72dZFSX
xJf56oLMnKas/z1b784OjIrdxFD1ft1p29rGXHU52E2Tzp/68MRUBgW7LUNf2c5g
QGcH868FbXpZYOyYo4Pk5OQXUbxUY6UQENNwrsnuxAXvvBV+5M9hyZWt6TDG6VhQ
uWwaGCDXDztGcdyNjNq0tFGnr2jWeuUXfjvyVt6tVNdx8LcdUL9NLEIqecOCEIoO
hxg4ATIj2NkybIjRf0xhSWk3q6HXsUOSE22fnNo08RZS5Sm5nCqtLAqAjEywpFCj
7vZs07rX0FxXBtQxLokVC+U+YIbWneWw6AgVwrbAwxI7MdEdvTai+08jTUYT3pOZ
di5hAUd3iqHvqOKZcRKRkNramyJwng/jbOqnISKsafyIjKprSbvepAzLxa6v+5G1
VlPSk96WbTnN0PuGL6PK8r9bd55g+Xw1aj+AvfuVGJaO33JXhjLl36fnEuszQejf
zlltDVj4Fk/c5UAmyhVWlOuuCrNHTeNGBK18wh2PkCGSXsakqNovLCUTgNZYLK11
JbWz5dZa5P/KeQMCE/ICPaVTxOEghJdbehKFiRKr4KbS/a3X29Cz3YTdZlVMr7ZM
2+U0o02jH3+KP05s8Ifkwrhr9yA5oPzYf2SjXZw0lAhgebYYoEo4+Con5BHUFHO9
siOuvdzXzpcTmIC/l+hpCP/nebtGOOXV8Q3fpzijS5SZSzYRTAxSAWetaZwAJ/hB
sBagd3sfmardYJlVAqbWJYHO0i1NUMp3NfD1mz/v8nWiYKHF/GZ4hCBWKf+K5c5S
d3y9QOWCciHrIEuvcO0pPie7QSaE7PNlzcBpP/nUcTUoTip4AUn0eV1usKlFZME9
evdM+1xofJS/CdVBWIR9mdie0/6J20ffRd0bDevDI8TAs37Zq5IHqbxztOgUiJHz
vJRshtzfEAoOzl9/pCc66g9UAi1R3RraK/WKYkejW5fmRlXxgkxcQ1RfWqWkIrhI
qwE/gSUotmY/Fo8ueIkjyeCAoNV4bY59PtL8BDqry8LktiPip2rnFsxI2dst/9dy
V1Eb54TUD3XCKnQM7T1I8eKZjR4sESYFTQZWtoJxkVwR0X/Ird4mGb4AWfxKJqaN
e2vIVONLvq17Jn1uvBEbzVbVuHeuGE27ifjkzIa7diden2uA/xbYME29Ec8Urgc6
nsr/Va1JiZsXWhpJTFIKUgnLqsmaKWX9qfZfQpQpGZvwllQsRct1eNLZt5chkRBu
HSsxe1xg4I7T01iuaWutKimp2yA1VdYHoMnPMlCkjCLnXEjb665PTjwjeNFpEaU/
ZB+nFP7hcvJJ8lRb0+IWEYWEYo5SNvwCfEJF8gD8u/un2CK+/FVIKneOLk5W/Wiv
OEKFePgAdxVI3KLfCPmNGd1VVSUgZ3AGyR1X+9+oOBT0i2KmbIY8G9G+c/hIPOyj
ni/ej6CS1bHiyLQ0kJgna7ywXHjRh1QQZwtvznmo6cXHUp/5itX4+z6Q3DufJIRM
TGLOwksuePxNMl5p1bJBDz2PdEbaDyJ3i19Rc1yOXKa0klUG8h2GlHASg73ET1JD
epxnCtpZFz0UW1jxLJ3qLPOljx3fdUD+8jceMIMRWz7KnfVN5nJBtQmNX8kGv4C6
YX0FShkskeQ1a+nMpJ9WkrMtAXYBOPn/5s4OCOq6ImaQ1IO8fENU6iQUeciOB8nb
0dTM2pVm4mNKhc4v0rA/Sl4axFRLlWBy1XJAL18s0jx8jSaLqwkjsin6vBZIhZst
Gr9RxACEsVAHqFdSNRfRcLRo9sy06fcvDTudJr3zGj7CzY+WpdFAE/su+6EiwL7s
rYEOrlWdVpEoJVo920bE88bmuHafAnyejZKp653+fq7METXZVFs5JaDzlmYIcKaB
ApBAIC/fredtUK9k7SdlKiT1byBye33vx7uqH/kQj7c3yd6CXNN9fdjbmmgApnao
fU+/6oyBxT3wAn+cFHZaB/k38qZG9P+yRvmJ7qTrypFVev0dom7GZ/teiNyhyDBS
tbo82ndK8eWrsRXijI6PqW5KAxIbq98SgdCxCmTab3YH+wh2Vq3lPKrXHetKDAix
4r04IXpneTMWwMHm8Qm27ACP6Lk5QI4b9W6VHq02TQetCDgTizwxkNEuOShjxQLM
4hhD7h9+uDnlAAj3oXSqxtYYj7w4HylZoEH/eixZRf2Jgt2P8eR52C6jzYjRSW0N
0K2ynRuM3XkhaCAeGVznIUVn9DyAXGWH0ajpK7wKsVe9yirzVMS6pDAUOHbe3bvn
DDy9cPHV97fj9/ajAj4RXJRH0McjhPP31gdFxYc/aOkvkVbSm4FPTCQfw4doyVwN
BdSkxamA//47DQbJ4x6T6NhtBe/C8YFsIgetiuJSpiZHB2ZTrQ+6ECPLHURiJQX3
DiEZCGDhdvLugp9lZfHJdY59NGf6rfOXuo5exWHVZJiLSEt/Cis0h+XPMX9V7To2
RPjefkaRy3K9/ZoVKitSx+Nej/MtXxIm6bIxy+uI9m/VbO+/2sAWU27USfV8zsBS
ZrFFu2lxSnjMaspwq8XQ+XSHx6V/X7kMQhKpPiYCinkc3WCxX49JKCW5pUHjlQQk
eIPPGijL5o8YEiNRaXjX7h4uWMixAcjB3blTqzkF/RB8S/HF1tJhw7rz48NTvtRS
XTaFNKi4i8HT0gWnjmTwYEF0pIVtiVtNRtIE2wBUqsdrn7OJQn2aHSvDGoVZN7jG
wd48Z7zgY/0djMLmg9tpG5zhNRMNBjKGzuy4xEGOSbPSE2lCrVIXMN+HtPX11yYU
+JgYjKrqy55Cd+cobbAGS4KI1+wUq5etwPG83ubSfUIzadPXsT+woA25/5qJ9bhe
nxg5gTw9NRZ5YzdMlnNcsqYoI/6skmLXLUyyxUDdXmHIz8jVUc2WTW+o61MzdM+y
IwBmwc4zFrKZSYt9QWGVZyfKLtuLTg6C8vS2/xQKwVZhveMh/L0t2q3lj959n+cl
QdRNmpmTafYUCH+AlD8qqAMid1L9f4DpdZBcKDjJwJ4/ZmEI/dxh4tMspXhcqwjI
3vXBQ6t0uCEONm95ow/4PlTxB82XArVrAkFx8ADHpi2cSfIqEJUAqtLXZiudYtmo
V7CwWygiLK5o/3IDN+L76r74F/BxQiLkOcJ4+LkPfgEcTLWgosRJg3pb5jqFzknw
objy0PiYJYQQWATkeYOcVU2SCb6YCEXa1NkFzQlfA1EHcZJs0YU3/ElANTi6DC4s
dNIQcoyBYrIg7roWG4UJXqUlRucFi08acliplpMLfFTCiae9+hhhaDC7Wm2QXBg5
TjmF104mx2BV0Y+l7AqqujmTTblE+C6UNWRgXbkpvrnwQnB/RXKq2eZOLzRVue+D
GLEciRONwR+CAsF/BCbiKt7MEhzwrmt22ETYF7Q6nuCkIlJwUZIHTJWLfCZvKbgx
RHpRlMSQy2tm6sXcK9Ccf+FR5a6WtknbUiInkVInE+jsEeABHWi7xLioI+6i/CkZ
9Q2IiYk5VxJxGuI8wegxD9cPU1nMgVENVpb84Y6dnB0uwDRTmyYyA3qMWTmq1rnR
ssxfFMFsrzNma+roOjtzrNSD/wCYxDB0j/SUmrByGnTbF32/ryI/Kwnp6E38JHn2
8J695suKItvKTPACNxVvpTo9lx8rjk+uokD0eVDOeeip3BD/9C5Fmwgb+2PYNu2f
qGl3iABsuIu5PbaORUrGlnBlqceo6dSY/7M7SSiQx//9UdeJnjbE/zRU7udJcBlm
s5akqiCx+cjfbTcPSWGD4dq9tBLYGotqelagafy/DncZC9ICxMXSQ1cQyQNTU93W
0ThSZKrFo+vkbb/3jYjKcyLUL8VDdFQSvdADl7y5a+Rgc1/uY+I2cGzcVwjGCfm6
QIueoaVXjJfb2Po+BvjuI4wLZJzcnUonLG6EdUGU6hcHSbZRwQVGhcfIDP9hUz/2
ZglCmfuQe3S28wNdn5B8w6CSB1wE21MeJ0O/7odku01GM1wLxCZE6a6pXV2UIL2s
bx4YqJ2ywv2kx7YefIDo+3WpoU5iQA2pLdf2LVAO+eQypISrvXr+owr96FJd8ywS
lQbO5EzD3HZyffHLP8Wt7hjt9n5s4dpe48XQ7T3YJ4n1PhLppioJ75rBMY4/qflw
HGRME+U+dAFmDWv29zH1aiob+Ypc2oV4fYn/X+VuZg1tm9q/tq/6Bm9oY16JC1PT
bgfFoSnAhIbgK4cg9AIdQUs1HhKPNGBCHm6w/uBAHEnBLmJ+QphJMQeq4BocwfZe
2udIPgj/5VpTixoAy9rZvIDKACiE7nyu2PP03HEfcLpP801dk1GS3xEtGpTJz1Zk
vuLRyWfIys28twizvOgSWuwV0+pUxau4Lzw/kwVXFjQHqgaFvMTf6X7hSmbwaEyr
vz6VrVevYWfZzupq+un0BZSvYrtRxwds29CG6eaK9Qd7ZC6cuwJiw5reL5w8ckw+
avKfMZmYNbx0GBjlMJ/8G6T5OzUCG1eXBhR98LO4J7dIcR/252jIO0TtqeMUrfrM
f8f2EjzHzbdB8GdJz25bYY7qNkMUBK4+8PHjRftC+9Al381PQxKG19YCVt66dbik
12hWvh1weXoD+4Y/NmKhEM0b+A6t6tLztshQXopEh7sUiDBhHsu25poyi1Ilonio
ZuqDba36n8FqfDXyomH9lH8WLCcDWhns9NRuQuVCZG1Q3x71XwlpuwjgPX5GOVxk
+fVAJl/nmeeumid7+XOiAxVdHv9dMDU3rJMTkBvqkyxv5wCzbVVcummtsDZICBN9
v7sMUS7Q9NQllXqDAPE79x82v9drm2OLZs85+K6ezR0/9mi2yqc2KmztvJacf4ZD
Tu69YhGOKZQz0IFEquoyEYw9oIvJgVubRgIKdRtbjiQDlBZIvKnv39LiOzH6LZZB
gDQckd+nTRZWhPpuSKr6Qp8zeCWdf1NjcThwgKmVa5dieWZpKqtA7rKbDTgk7/F/
/3zC9Ctr70RotOM6f6w07wPqklwDx5P9JdJ0lGfLpR2aJ2Kb5A28RQVBMOXJqMyw
lh6wtsnrb+Fq7Kaxz+7N/fhpX/v5zogVeapP2cwguwmnMA8GhWaUPL3jZf5T7Ild
gXxPK6mHsrEZ6g72CQKgJP7ko7Xn4pwseEBitHrFPFHVdYctm0CJSHw2Rt+oz8X+
5w8IHYO/y7De1RhHbggKqwxokXUwr2ltgPbOSQ7z1pnfzhhaunkNuSHiz0HRssAX
QGqgiUkbGGRB9JKBc8AjWuYPx2jT8jPl6H1E5qP6gHI8ZXFRqLiO+YcAe0CR6B8G
8YHlDN7Opdo02Tmu/2Z0rGYGNGUzaPz6nOEnmFSyQd55p/5cpA3OCkU/QJZOp2Wr
M3fncRFNkvJjB4RjeXZv+HCGldrU2XWefwSXo3hfvIfxZl6svD6NNKyAAahns1BU
xj4uNcPNBOQHnD/jTHeDsfGpIVoA97iwOzn7MkQLWrHNaddshVE3fDxtsLkPWlY2
mnyS5TB0UXv2cdHGi86jvXdD/2WKA7mHKXDLknmad+CJw79aA2kS1SWuR0jGNe/X
brO3MUd8yv8JgH1RzfMbGE89cHxGVHruLvWiEgTeiLl9jfBRejAbnHrs0c1BagtN
D6tTyxJlJnhWfOQaM9HvBCgeag0fjKtExFcP0W1Xv5iUsrCf7Gx7io/7d48yCDuc
xmPmHWCUueQN+X4I4PXbe94arTZDNmj8kezQQaTy+EgMNS5AfRKFOxOV3C6PW6fC
FJdqlwiwFt8GTbfrtYJlBeVlQ8ifu56jiTAPpHUWBAxkh4s2pCnCW2hqt0b6gZ7Q
EzP+onHoAfULRTOy8+5Bgrf4WcwRQRpzyOlssXLJga5e9ughgR18Nq9SjAD9p9S4
lZjLDch93CZOGhXWlaMwjloQECTiH0v5IiDoBS7dIbKCgfG+cDXGU8xdGoCqUDrx
T2cfmYrnIxs2DgDhmTneCdoQsaFd841QndBDzb+F8bitrTwM8HTeW2JtxNrECPbA
SPVAilInlWiFSlNG+N6ZhmTaeWUDwkcT4B73B6iwNSGINLz9eQ4B323Ue3X+5W57
u34UdhlbngNoAayJzNDJ6biWiU6RClRhjQ2yaPX55nzKQze+zYg1j0IvTQ+kVVEM
FcX5ncX2HDXRtSjrUrd634+c5+QguaDOkSbzv2hIjT2Yje8x0/ydk/xgvGjQXAHs
kYJVvjX0t1KWeRELYrsfoEj1tHKdcMD7slTU05isSy84aFy1ppal19KRlVslUKLE
P43DQJccCU4utfVivTpWlNAYRat3/bUtswmj82Ok4giNsyX2iOC2vm5Vb5Rr48+y
lGaTAnZZKaXHwyjI+T/L+mWM7G5iq9+xYsO/Yhq+nT/cHxFMdxQfYqzGspz5DEKT
P7hkkh54ESsmDttjviO5tRG4QDx2VtWRiMi/no/RvM1AOtGpi1zfvAjn68Mf29n2
lyg0UZEnwrdAVhCzoIQoaLlXy2BlaqjQIj6aHQEA5RlFP8CPVpxQzX0suPEoaDev
9NUskSDz2bBfBHBDCPqYE/aiH3faztC3ZgABo98h2vd4UAOuCgLzayIYGlnakONR
wFIR1kUBxUQFSmRXL0d11oVrEj/ldnbhWq08LCxk3OBoPkmhp9YG/fpiyR7Sn6ps
xWrpziEP7WAid08rYHR4RMPMdRP/HwYK5GhJbS8PhHa0kZNk9rf/EphXKyswhya8
lOg90ZTzOrOyB63FBcQ61CB5IMdL3z6ujRxppICsMa3P4bwDWYJuhBM53IKH1c9z
SWtNxLfC0sXCT44CYzBFUUfc9axjY39z+ed5dGGBzIvUdz9oGfSv+JxBlOPhw4GV
LhyqFnbUDUL47burqhIhYkTkgzUtrfu7sYWS9pj3QkqeVRoI7z+IVHVFin/jc7Kq
kyUgs+ZSBrTLDexebbaha6BOd3mqHpr6sSe1yXgxNtVU3INJ53DYapgm0+ImSEfU
djF6x3h4wqDYIdkfJ0r8avAfKo2ioNeaCK6sIlGFbnxoXtuR++LyxzSgG/X2TF7P
hT3m2KkX7Lx8Ltqnu1KK/PX7W6pHEKM5cZhxQfkHmFMjHhxuMJ/soqEax8BE4XIC
r9B46dPvv9hMvSEK4YxeFz9dMJpBLsgfWKEIQbX9jaNnbYvST5nlyO/iaweQV61Z
Nkb26hXCMNNDSGJU4fTAByFZQUvzHzMamiiq3RZMo+g/zHJpCPZ+s6pzteq0zBqj
+iWX+4saDRep9pzmuQRHW9Y8U0oipz+XEFHwda3lNr6bsr7pJHtX6jCitVpXsZen
xInCCWsokFl1Oz5LhAgYoIfBEJaq3+f43foHH0nihmqwC5Gj6+XCsnt0lOVMVikx
OWMkrNTdsB6/V6lQxj3YUo0oZJB+IFw0o1bbqxk437816RYlVG+mB1DeFZcqqNrp
VvnnGWEQuHqDUM/3mSn+NvH3lE0jx/n48bOc/TR2M/QAnWD3o6uf58htF6KHwXJa
zaPyglOQsFdvOSP45EYmNH49guk29YQt9/ef6NJHXsBLWJN1kFaIWl6Zgjhe4poE
wHJTYlvnT+4YyRO4/+nKKXlnGpoV3gHC1tfQcBIOFhdPCwbCf84nWx8ex3WsUYol
h3oeCzyDb1FszOmH8ex7rtKSHGjjEu4/CiFdXj79W9ccgEo4Jk7Hxdeh1w25Dyqu
62qF9W43SacqHxwqGT7QVSGteNQg7ZCdmSzrM6tdzvThl3Sy9VAPkTBFu30+hcHm
uV/Tg3QmenPEclJis818x97NLB/Mc1TMYRWqqqG0gvd3vxrlOTdOBtbTTS0u1SrU
mYIK8qjMe0XFKpwQjkajFbsGkL31512XPEHdWAVrykEXDEfdQ7d0xRPg4l5I0/XQ
lhbOnuS1SAiVxNtaajWzXfbmAaqdzUU2Oy/8mcTyt0vwDnORINKRerjZ9jT1EUkA
22IdzfqVQi4NzlDjUU4xpufopFvFVxbLtc7fMO7Pb+ciwP9WtOKkzH5xleE94amr
P1Efe3xkQONpLd5pNkqK4pO41DZAU5voMsIjQaTG+PdBiD1YCYt486VruPAlptYv
pVJVayiNREPV844hGVwI7DX1Wu3yHuExvkMkpcQIpSoNVg3SU7xXdjFfUZeYSnr9
sFVg0WpRsgJUdCEXNlPmY+agvPHjEdYA4ziualfELBcplEp07O4mawPYYcEkMEUz
iVQGFkJP+T907PG66K92M26g1xEBmIC4hrNsa0DvEXLifb7Q0+11xYFDbGugaxHQ
OLunFMHtsLwKdIINGCy1iYvO8E7P6WdQ/xw44pr809JvGkQKMSbwWfXxOzRD7wDL
kPJT99TEYIkAHUXnkTSwDJ01KyOL7fF4mmFAx1VVNoJX60qRIlSM+hsBOxIEZRM3
zkHszVxwVxbCxhRcqu2ZyqKCdpwyqjZ5l9uPyv0NUpJhoEMg27oxAFiu8pjTw3er
MSe+sGjsjBKZPIqWrhEFFXw+Y/Vd/82+yX+BO0myhOt7aCx81EcB6efw+eZOAGDF
f+txHbl412R2dRgNZJWeGP6tscTIgpHdKywCf3Zc6T1Pd53fBJAekPntT+67FIJ+
v01N2pwjWtP6F74Fu3HlVm2Njh5feVlYgT1Uq7RYe/L/d0pXPti+i2cKt8MBpccA
NifMLFj8u9/9YPiJXpP1VJU9qwzS6nXVTX6agm4Vf03kD3Mzon6x1MgGyKNgCEaE
rXAbiru4kQtU/8++/yWnMyHTv7epx7LjCGTdoIAgLSfgXaTl5bEfmvKCGpYKY8aH
RC1vcF6/fuGjazSSko0jKr1YVqjPG58dfiqzhNOiwq+pafXP3xBeS/vzuTClpIP0
g4FL8c7sQQtGc3nX2cfF7gcwTshDbFDIBy3H3ySMFtHABy2qHJ5VI71cdCuKqkcW
PblSrPbcYqIxO15mrx4QUaCc+hf5R8VfqGh7My46EovtldwX+/3tlMMALFiSpy7h
WRZmskVAiAikQ2dR91hxS2WMXLCA+NGlgDf6u+AU57AaLDQLeD/xXii831tIVJsm
6IcreL8xPJuqNWRML6q2C/ixPN9kpJZNczik8tu8grE50O66JEgLB+0OmoIS7Qum
djBgtbBSa8NcY65P9OUi/T7Ue71MCH2VbKBsyhRiyl8uDLPwTTFBQ2yu7m5I1aLQ
00at7yhO2np7bPo776ApeDGA0J5DSXRA/Mm9n4oVjnoVzemOOa92vWNEJkRNj90d
RCegI7Sufg402Y79dgViBa+mKAApdBQe/U+/ioF4eVpbyQYe2GFkJey/Gb84wkb3
pP6GBc1LhJ3uFjWspcXP/kwFGtpRzCP3G2rDQBLSLMmtfQxPeDmJk3l+vIGTTBbV
hYdPqgTMuv7fuUpsyQaSKQz4cFIiyOXea6yDkRASn5ufzOGhVy8cGrFLDcRSgNlB
yifYU9bcom+LAyAf4759kuH7bXew86hvaQR6HR2P7cnCcJ6dl0RnyPqN4WOEAII+
huu7Uvoohthe2LvRH1caz1IkcvnP3AUzG5aJo92qNsT8AkKN41oZIGEmxG0B3qG0
hZKsm5VkL21JukdWimClZ4yEecDABEbyFSlUgBVQsGl7+LICRHSLQ5N3ByxaCCHR
T0G72g6QI26BlLQjW6zYim8fBXFK65dFqViRfJUMTrLF9j2/HY0VZusaIzLoDIPA
jbD0SYXBwwo0g3/epggrkYyyj6Db57WzpeBXcPAAdYzI50KDiAi9/5xYRCfCmiYo
mVefZ405MKPBYU2z5jbF4qwQRV4lXipOP8xzyQeBqRTXrweCOvx9u8GO8s9JnxAC
YGCBYj9M1GsWqPztM7rQV4DvcFKJ39/GfxWKpqQHldBhff1plY71LCuVq1V+CJxq
l2wdKF7J4pPTBUOHS67sMyxQdWLDooKzOV5zjw8jZKAf+9GuPBjr/o3itJMfF369
zE+RP/z0C9S7vYrYBuJfNHabJ1AIndJiAnKrgsUgQOmDqsnPnLO3+ZTWgxShSptp
7MY8LHYhPFefB/tCyt+WGMXtXlCAiGX9s/S6K6hhCxynEiyfNDyvQFBHfbVNw9YB
2QJRuaZ7Ml197glHu1jALKXemfQxl/XSalrNUt5YpN1xrvuZh8vd1v+TW+Z6989S
FUAbyRbiaUPlgEP6YEdup50+5ypPVuUosp4XpG4sS9OXELQOJFOKXzc6MTtPuAZN
YQzmzMSE6ELT1OeJTBa6ZNyysKziHqYid2+1FLcOjsHM+IJoVoxcU4ywuSEH6nm3
gPnjFTwFUT2riBqK5AtI5Th5cP+QD1qPqeSAYhEP4DpFB9imrl7sTtvaYV+e6poN
1xL0BxDoo98afmEOYHOllCc0wftN0fgv76KVQawMZOPvqRpvLkS40fsRSZkCROMK
U0TOLkVrbTUsAWFktO/KYI15QwFzhK79Z8/XKEnvzs/wkzveEd1igkg6LuNVrkbq
Unb+36J2LXKeqTgJxAz5knzmKmCuTgCPqqO8KbK1JWRZM/GGoOsCgCSBxNurcn/6
t3qI4ELdH6y5FFl84LDcSS+DRYrbQsfQY/AcJ1QKp5CBALYhp+pfn1IYtEVB2P3u
5+hjMX7oBdVcLp/1u0gU1gewnQ8v42RISaKSfwdaHub9Vge0ShNNxfpe/3stYykF
GDzKbaYjKG+GiXXdkx23TlNfIr2CqL4nrs+uOvPs7VPdJrotFZ4z24M2jowD6S3D
XiIdEgCjVJxtEthf2mMfOWqqzORKi0H5bcGZjDEQV3L4Df33ooGIBuap0w2FUKlV
XvgYi5873weM/WlkvLnQo9QVU+ZhcY0eU6muUC1i/2+JhgNTS47lbjRNFhBRZWIN
nbry2qrRQZVqWXsEKCxMeCR1FuLTq1uuHeqWmxGXKLUfn4nbdcUsazTlaWNP8XCz
FC/WL6MEWUQiWUJagSs6WSCkjsEWvdZZKft8OB6MeWf+cacFGJ1YlczZXYQGbtoA
ngFJcPiHjAZLzhibQn60AeZeH4p0GsntVBIJ9EqRbxHxplUebkpG3+AiGEITbIpC
Az2dm6cq90LdWXrRk5rgrRASAQpuw731u29/pva+UCD+jAZsxXL20i3fAYBnDuZh
piR4xIfnrZrdUbifGPYB0QJsT5AbXk34nOl9btAPvw5gWAYAJN3dDBKYKIIgGwGN
/AMtQiKCVJ62EJD5e23ylCX84zUoqWDTEqnU5cotzp1uxjmHE/rm0UjwCYqELRf8
H6TC/fDx1qNzQPbT4pwxVhh4+jfpQItLOAqxnBc0j2AESGmClihgDJ5SURgPYRtO
NxKWyKGT6+iHQUaGawFSMjVZNLhn3P/TKwz2LCLwvPT1l+CUwMCMZPy9hqb0rBMw
Lq5WcEVkUTVUi58ubRknuoVVk25IJqTS+FLDTeHklNy7KOF7xt+gumJp+Hx8SIWx
BghVjcJIuqVFjn237YHNZfqce7PQkM3hRnGMTa5DuwTm3oFSEXPEIH2oDGbuG5of
fUO6zrVEXKamVWftOzHhLK36vtsD3Aw8+DASijYswpkFHhYKwitFo0YJ+EGf/0jp
LhqeZncCwUk6MyI2eABujPJRcN5yTuNkt/Wzf9WDHWwQVY+QgypiQlQOfRqNyNv7
aV+sJD0zkpb6Nf5stABqyxQlhvFBCvfPSlRWm4+Hy68AFuqOgTNSEfl90Lxg0KNi
IkZ7tgL+jmyNoKOayHXVWGTc6Mxb5zpv0ZbF19d2Qdw0TVcqsOrhyIv/SYoidga4
N2yGcrrcvGkjl1rMew7CvedxyUJr6WluG44674IJ4DK9zLRrQavRL257De8BTyC9
naa9NoMl6v9U57LpNMD1N726IMCeC4wtZX1tU7GKoi+E1fXF9Hj1z4mAgcAt/pVe
LEm/I7Qrm1CN0lP0D5sG/hPwPV3JDaNdbUnvWmIo2ipogvo9Sxq7FfaFFz2i+mYv
t766Jew0aH9+gCKOsY5HVj+CmzAFtLIQWAccXJ0q6GH+lEXTu9+8o8Pzl2JUSrC+
S2H7K3YqbbLae8Ilg6/sRKwZ+FRQeafziSbNJci7U0QvixvP5lIzZMTn3bd41878
TS7W3efiGB3CX6khrGoOfArXoacU0dxKDr6aACqA383WYMS70agGaZuO/tDg7Kml
qvSFOvWP3IbZScp4Y6aiiU/hXFwuS54XhhTPSGLd4Iwvr/YpvG/9CWwSBFrdh3S/
NPLHT7oDroMJMCYXpzSAHCzTRAy8J7fgIbPDhAaLFWRjHim44T3m7kUf8Emqkilj
4xRQjl7ziVi5VJ7gHAQSE3KocPiMu38KB7AiBHIKKYX1QhIWEhfk1xsolxx7irAS
7/G6fgjqe8+pp4kRXhQ4jsHlLmufN+G+qNUuHL+w8xWzxXHqV0Pne+2KTR2LUUfs
01LZW+sS1Askxryh5xa0LfO0WaOEt61nOhKmu59ZTlgjU37dIS2jb5EbWaZ+309R
xlGfyp+tsh3Gj56iRGv/pevtZ8W0e9JkafhRAlr1KynOXjtJCoN8xZBSoFOIhzYF
pBdI/aQ2+rwKJGj3TW5LETUG+KabJ5rbfncb25Xie7dFs5uyjKWx1jkSQt9Uls0i
Nk63oPXiqOzOEJShUTVO8gFVcV3zfC+p82KxMIWolWiVvfC8s3mlqi1jyGg4iDGg
bB9c/S5agf8+eH6pqX46fvlMqDzT/Pc5st2Ong9/rrTw9nMBdm3GccRTIWegLyHh
osfiiLpFMG1vsiqvmmaGrTn2zarfE8UKosYANU8922G7ImRT6lPHdB1ue4jU6yga
RMjo3TTogcX5ZoAYnf5FMEcbKjCimvHEoCDkvcXKvfvK6ZeiSwGigDi8aIPO0kwH
cAMKhdar3olgu/5uZxJBWziJRQYa+vMa2ByJhLFV4w7M1Jlo6TILxizlXtzWMyNc
1WXivTSMRWdzVvbU6K5+cmZnYw6gbzLpW5Imx2Jv7PSm1zlBlx3s2qGv45r3pRu+
jeSPJQsXcD4VUQ9NmJjdKTXfdDr2JRojWczht+pdGf1SSQPSyu0045KeKa/N+Con
BA50vFyfGgs+jLdYTe/STSiJp6HunhgBPnEKMRLKhYd2w7b024z9/toSydfGKugF
f2erMmPBRLsXU9a3sjf/IOQ2mSVoBz9SZLb7JVXGfkVuWClR0av+BlHzuhfzJlx1
5nfNVXtYGSzv2WXI9b1f0tjytRAlBZxBRBZA46PIsobFfseC8Ov754Tti29m0pWf
FNhKXsgOGsWAYd7bPviuRlnHdUqkxcmtEHo6q/wbQvYK81eYeJHSkBMaMlH+LaCa
a+8FuJmSRxr4AKk2vbge+4BcHHg9JIJ1gO8S4dmKFlfnPC7Oe2pdQy6qiYCYuqFJ
rosK4XwRfAYU9d5Kvf/Tnb0oU2XOJiX2GfHZMbYKpZQJX5x3I20laJVFU2NAnlVy
ZzCpfFGqUWsIan3fmc0T6neM/OGPSdA3YfPRgGs6POxKuxDNGwIy5Xw/P0DL9rHh
gcIAJ5YfGJozErGJ9MGG+ZemzMbVvN/W8F2yfERRbV96RkTSNMQEJd5rfivHv/tl
rwfKWc8crk490SunYmjigWna35GNV53Zi0+rANoPS6Bx6Fh4qHH78o3TgvOL2rOi
mnSTGpXBt+t1yFugBEO/ZXFMp4eTk8HJeydnrlzNQNw6DKnNWKUiWhrGqodft+Un
8ky/WkC7VTROrs9YA3XJz8m3sjfBLNk02hLF102pBQv9ITABlnjJvY3AaaE/KgqF
LT+b4KJsPFTo5tKrxsXzKhZ18ZjvCos5WQ5i1QvVXTE6zO4e2dtlcLBg8EIyLEZF
bL/Vs3fdfwaDJHbIB9oJ/0ykwgIM47q2cuMuAwlT+7tF0+yvhgxP0XIfmVEdpC2n
vS8l4NV/qlwZLTjwIx7J6+ZlcpbVTm2E2dTUpG/3t6/9udqrpn6u1tCMw3vwxT2T
u9rcW3nJfpSqAMjhEGHAiEGzRordTOvH1rsYXw4HcroZ/UUHSfq8kP3Ulf0qy+Lp
drsQBKxZFbKYni2GR8xYPZmTU4LvQ1SfmNhjtSbFZMScW8rzcw4z8zIVC0oT2CPZ
7pLOu3OkjsRlwsdkSAEBF3qIYnI9m5F4rd3lEsZdF/QxBJErkStzlXhM5bokH+jg
WOu6nkjz4I4GfehBoeGFJKKTFMXzA91JHWa3Vsf2qL+33TR5CXMEx24OP1ghMy7N
KibVWQqJBmtonrGXn9dSYTrxCTEY60Vn0cinMNa2v9eAdvfa8u+pi5vDaxX30Ueq
Hm10UqXO/r3VRemU868fYpwnCrlxGNCttRby1j+5S3Ik1wHXQ342gXndncp/FEth
FRrv5Htl9wzV8er6INGuV1vexnSPS+8hajHm5nNHLjoqfJygxw2WMoxz0O+A/mY9
S0Jo4M/ZTKw/hQgNli1RUflFlE9O8zS2UzU3GWnXPHbyHXISwgJz0HFTFCwUS07S
ptu6BVX/uhaYt+K2czIBhLQWGtyEgw87hzieTbFzfFsKtsrROuzU9e2xX/FCYm/w
fMeXepPCUq3pDQO0tgFTC+eMRAsQQCpxQDEYI0swOu3jca4Q/xZqmdpWaHAd6O+K
pzNnEkxJ6uouNidSReQ+yjbGJoReiRarHJqaPzdc7VNp9Wdwh+/DCQ0VsgQPitPB
NJ0TcCMEMO5GEUrrBrTr3CMNU/UUUzZtIY3yEMUIzgqoQ1EmgIKoSw6PglUi1g9X
DlpKc8Np8Du7SdsyAxyvnH2inhgQ7tg8U09g6lnsSlyQoMXxxE6dhsdm5o+funam
kOivWbXzKFsHmKcLWGjAcqG14jEwJ8cieGHcbB/5WESoIC9IqrvHeGE3LRnEc1Fa
sISQjRqHJGDzziRmv2q7NlXb/CSXlr/N5N/M5jYhpOzxChSlrWGuKzMiWz8BKSzU
Wd+Enk/nFnNiSLu+mtfA0rTNinLK1R4ml8uMFEKzmuh5/pleAVLBcDrNYzVrCW/S
67KklU489mzApEYY9tFpf8s04Xu0OiYvY9PIOHxv/4DhEoocpLpJh50gQopfZC/w
8K28ejvRYm0xogt6VYbASGFJbXAxblmnkfOPho9N18Fn4cj0ayjvUAQpQizTDn8I
ZIBjnfU0WZOKl4FrRIWatYMh5GqWNAVWyB+mNwNT2u+/uA5+VsXNrhvfPll1kKBG
EPEU3n7JBRCRfNxCjHCGiJkAIcHTCjxwK2/Lne+6KDGtn2qjDsYwEbC2/8hvKYtm
0Pb5fOdFkwPPeLmE6ht0z/gBp+9O44+89aeQYOiwD91+kkKrJ1+wGxx1iP6jeTlL
1XNt/llTnS13Vy2kcbD8sJpi7ph0440IjqbWJ+v9brOeTIrlJXZe79MvyVkJ/HEB
tL6hs+3TQhLP7ENDyLZLhShTM4nIagNpsXS1CnTZlu+78qWpYZNnvTjXvAm7CFgb
dvXTB0TYENL4RmmkGlOJwIoiujyvAZ29jO2fUfoNxykxAjHjrF7b652PoYpj8PqH
iTY5/YPcWXYMMi6wtYma/Gyo7rNGir/PuZzvP+OBkWTh9qh/8W143yZwkhJ/gLwC
lrl/hb/d5DFnxVH4mBKEMyxG96cCK15obDVGzi7iYUBRF6RkWbgewYTCqivseNiM
4u2NX7/8C2BPo7PIUjNEbxwlVXAI/8AoTtGdu5srK860Vm1H5Jv2UjSfNxPDoKxd
DekNrk7vdqhiYCsRJykX3SUTOjUseiWDqh/ut0SGe7K6AVVFznoByEQHUmEoZu4U
7nO5gjqubl7fKd/GopvY2v36zOTGC8Hg9I421rbWV2DC+DhEQNOo+6b+xF4raKpE
iqHHoD92vc8lILVa44si+FhIKprAf5n4RMYMG0oyBrMnxqh89k8kU1Khoz8mragU
dfsMx9gIcJWUiFt4QwBXGJOYAFPfbMYlVnw8QNKDQbRlO69Vr+Nw5MQxuWID4s1C
nLN3B7RVQydF/4dgNYtuLZEaXjhUeW2VNwxeTxfGzkBgbvp7pmaNGIKru/Kuw/Zd
2/oZ/OYgMlhuBymqoJNLzoZu9rTWKCFba/FuoLQPclpM4kCalKSdP+H1KzkGQoc7
MX4FC5WdCJQihMnaQwppk0/9bcnpPAlF+a/yXe/mL4yJ6sBdcC54PkajD6mNslHo
L0XcdXEuv+0PbJLsZSGZRXL5jHhDlIBppRa0JG6dSS0g71/q+sYGDmCMOteCHrko
zhR2ekR/kAAQfHcuFj0WJoEloqpfvT9NCx8qqq2OfDUCUiExtZ6VNIeOoXaCZjns
UpPq78D+0Hx9vTz6X/1tI6ybjQnyHfxTgfi1Z+QxWY0NnI9dJsuzjwbspD2y7KUR
QwQn/uzPccLb30yxVvZL8n8SMAe08yrlLMDE5tqPAlgS3BqKS1zKPX5Xl7kWAUQK
QhF5cTUZYw7G0f1bEcya4OYo72G7pTZugV47ValdL48TUbc6HTBeUBU2F5QXC3N+
62P9nxsU8rvfUPIhAz+Hr8CwdLXrrAGVK7tv/zZHV+YM5yeOzWDnRwqmonZtppHh
7vueT1VXk7By4E79zK8Ra7NdRWmeoTNzrWp84GklPIY9Ett8m8ttQJ9D2eYoC2lw
UVPW9fQhMDQRWgr3BpVfc3Y4uq4SvqxJ0N1lW8p1VARa+N4tAFJjz1PBj5OqrB72
iHIKh1vr4OLkD4nfnPydkMMQhRwZo6i9fmTE8FvQAv89jfvQcHdjb+mFoLNaG94Q
JUbnMT/nrPc1Oj+7MDY7EroERDQQpEziu0xyVSsI80o25WpVByhCuIc8LZiAyvw6
DtdR2gU8150dwpAIhmGdhWNFX/vYSz2upZrqvcWsGb8K6tV4iCjMdeDGU50mXLsJ
YvRfk2qWWnlvGCoXvLoeaRblpymqU8Y7zc8K0xfIYxSIUAWQH4PTi0KW+1zbgXWh
nCQsUQoCYRLwYcJKrLpXaw5PE5R5de23Xz72yws53n4lnlvwI6yQzay9R4T8wu91
dCo2nSkdj49yTBx6FRSgTWC11KjLqP0jCeTLcoUqMZ23jsMhg1x+ugMZonYh9SJA
xy7l48hsbXRCbP7Xq3f4TIYmteStIyKvsvEjQ23RBXXjyCPcut+wkTpJqEXBLth6
f8EF1PbXirqjFsr4LSGOuY1EIL19RsReMnivtlawJLT8aJZJ6Jti0PIv9TaNVbap
twq1zAOAQGzKlMOttjf6HY4h6afHMHlhdrzG0LHWTYjUnPElehfKiU9g86/Ssq1q
02wUtO43nomkqeFkbutJ+ptooa1r91J8HKKx+ZNA6VtCkiliaPeVQth/Nw986Bzh
AH7LGcq3FfSSAeA4e4gernFxfqHvd7zMHk0W6I4vcNaHVs5i1jx5AdIcn1Rk+LDE
BAVaxBQsi12NO3NLY3dLYqoc37IuRv4vTyG3kbtZLagikiHFz++YhAeYaIRapYzo
PXua5/YrX5vwpeTyqqOk7cEeo3ZwwY+Cs9vMtWi6PNGBnOKN/Om5dKI2pof/Lh8/
qTs/Xbh8XGzxRJho5CicqtcSMgY1wu8VNr/CQbh0Ldh6moRZ/jN+3i8mPIZyIyxl
6ZrU6bOuDFQYB3atEk4tiVCSDnNjONnbaAwP3BNT1zgRSNXgTiNBKLC+C/4iw1TQ
6W5hJ30FVY8sh0DTSUCCX+wwUN3KaHqTccu/5DGxue1ns/hv9IDoczmIewUYQ1E7
j65nkZ931/om5Wj5Z+SxYqlTH1FO0F7YmIIIIZwHNMWJmJRFAAfqnfW8DKYEtBM1
ZopAK7HlCkDpymqTiqFzZkjjsLgjPK0TcSDFqE2NozkqmuRbrM4Ri72MqfQpzkB+
TwSzKqQrll20rtMZpDdWz14TeSdPXSpNclXYohjngfaVg3TTYYgn24eYtUpzw18N
b7vTDVyEvWIWFBu4k7WoNFPOoZhoUXt8YRTEzUXIT3+iuejjH9Xjaxj/A/W92Zky
ByU4z0ftxZoJJqJ7SUJqE5D7b+HC+CSocPcf2U5ZARksEe0lYcCaBEDJ1O6wTjEx
BMsU5zp2YSDmA1vFCRFGd5YodW0iVCzyb91wdwufhBNRptoQat/EPxX5QJO3KO7J
z7cCBaXirvlra9FV4Gs5I6NKSn/nsDVzxKWnNZnyt/22qLk66U4GRsD6zuhqI/F7
Z48H7VWa1SF+cPb7R3ZNb79MzQGCE7tP2fqJz8FHoyh1a8iVQ/ab68zasudf9Nya
4YgQubNS7FUga6Os5lmoD7ZK/Hj3r2be3eHGCW8OgIQNCxwFqBVr7PbsMqeL8J++
l+OaViHzdE87iEOAm0uhUmeKer4wZyaOFpdsmAcU5y313YATZnD6DTt9UMgowdgp
p8d0xiAngT5YlAdWqmwUFnYQBZ02PNT1LdthvNONCOpnzfsX8VmWqUngpyQUI9n1
pGY31Mk/UPQ1VXJrBRp3oaeu72MyHmYTj9oDD0rBum5ppTyaCODTtMhv99tos5iq
LOTyps45lZn1lPogFFEH4rL4ru+4VMaGAV0W2HUvty6Tu545b4krXJnref/FlzSa
hmkQTnqTclgBXH/nhP2ZFnPyddv2RyKZbwei42/dzGlvx1qLVJkQXcCRVyd4QilH
k4jdgsBbGl6PEq2UFE3vlA5+9DLDQVhEGActnKvJOb1o8cQHa3R6zeQo2yL095qn
P14qi4FkazDu4i6MYnJ88z/8dEoaKqMdrgNFhMtkk9JJZV/pUQ5v1BXEd7UfAmaR
MJXi+YDrqDcEdgDxr5iL49DIsCEkDJzAT4gAfeeh9ap9XoHYeVBTho352HhrShbG
u61jdCQzsYnCpY//aODe6305OAA8VXGumsPspzLYqH/QarZA12r7PAeZ6RJXNfeL
0w9BYopXVh5ioMufwQa8PVy1sfrbPFMUbc1fdfp44Kb5I93nn3xn2dNCuG32ujO4
ZiABHlmnhzALhXSDg24zsrzzkhIjbaRQBPNibQUUuvYOw0959hMzwWS7Wb21/6/j
Pm9Ma6V2t9KU8mOXw7fkpzBe+GvlRcq7qyRH8EMM8G21xRBMEQAfzkyJLGfDQh21
fS9qz5RYd2lANclNYkSME1WmxYoF0OWC1Y8s7JgmjiqovXI9PJ69Fztd2VbbvrMi
idbSJTNcBj3EL/5ZINnb2R5JlJFHYVxZXkc+OcX0tflYqfWvk6ejYX/zY4AVc96P
BOaXYK8ql1watMlLdUGT8VCaJ5V3/cTfqWSx0BzCWEJQJKpOYytu7ekUn3XzE4ql
/Mt7AFnldoLpXlNWJn0lcFJ1i0GSLL81cyVyQXaVWsWGifkwnBdYnfT18+onrU9e
keQtiK2j/aoNAFu2JIPdACYYg9D9NXZ8Hf83YOYUAX5Oz1Y/Yv3fqcybjAOJ5Ez/
67S3C4DMNJ6drQ/iaEpMDAEhHud1REoJPjFDkK1U74zZwbNcS27T8k8Cw5Vfqtzv
gdK81JQjWzXm0tAdUX6UZ0CwB/B/3zr5MmdBCdiYLDoN/xfn84D0i1iaf+o+Nl5/
DzGrOqJGcO321r+4nSM+3Sm7usBBoDZqo1Wy+TySYZmuiU3vTMtMCcZR+bVnPnOz
s4TwIiwtPzU8oJ52h5ePHSXJ8zjXdDsL1+3nd0z2Yhd6Gv/7cgbNttvQSXj1/NR5
W4plYRE1w71K5Gn44n51VqPQOXX7GkfCUQ5pgGQT6T7cMEU4EwjGlAGMpIajCZ7k
+rjLWNMmBCShcU8MFIdtdjg8vAvtbWpL6bMKO77jvtOTc0mrm9u9mgTnY8shLKtF
+jqW4zdjK10fhjnc0fVNP58zysSQKQJnzexTvunpAtp8KJR9am0Xbt/8jMla64Ro
9xx7QxH9Z2x9XRtd737VwozjphrhedTWi/xw2cemEqr0uoad0YbTrvcK/fwEI0Ma
TEQH/9WzRh3rhZ90Iz9qFwZ7MPe25KFNKj2WJ3uXUCgnlOLqecShLXK55kVJrugO
JMmqssxzCGlvO3emXJpyCXRaLbb8p6yDUkZKte7XpCQbYKkztkPjnZHfSc3kX93+
fC6Nfxs4UlI0GO34yIpwVsuYNqmVrDb+sQez6/DY8YhFYi7Nax9Hbbrcfi72Ad+K
FK5qDezHqLHu+I6qLgUwryewP0A7iNWctumQM0G2bvlZ2+7ZVvvR7aIf/KKUnshi
+hGm/xmvxDYg5XdqTrHEYdqfM4YOFCongCZPtXPVAbqT/m8UW4X5rNIY20duGFN0
q+My3ELijotn8mDx+FpQmfcKHfRFpSsOWzUvT4fqwmx1rCcJvJgtN627Mc6G3SlZ
eosHpv2LWizXbnWxLNzkEnyBy1sWC4KFGlKMly03O7V5jKbBY1OhCcBcvSrdJyHF
zQZSRqvn2iLeNbI8djvdOeytF+9NSiqcvDJk+0KUwdqfqPyu6ZOmli0byPnCt0bA
lOsjaNpuIUQ4qZE71XYujka875zz88pqp93zz9U0U8MrJubph76wKBzqflK2xrks
+OJPhtL9I7ErbIqCe4enTP+VHUaWTE/P89AZV+E3bI1aWgqlxWOnx7NIC2aJBLv8
NXLzuhZixOTz9Nyz5pKSIV7GI5yuiX2m2DbzpPuqT9X4y9ja7smW6Daxwt5nfboY
1KotZR0FUxNk/FBGEadAwSu9epTxdbwzo6aJMFZShxfYB8MijCXY1tRQ4nG6jrOv
+8bCuX1MwOuY8s083jPPzaNpTzSPPO7N8gh179sqPrD2kLG3VvF16qyFTKp2sqrj
mD6n3MC8A9Jj4gMKeCmk+lcyOjymKBlRsDdkLCu8tMZoKLu2eUmQke3b9aOdP0iK
zrxiRzX9ggkJALWHxyPQCZVcXSc2alfbhJUs061Wikv+v3WTr9SQVZtFlbcJKRLz
O5GP98uVO8w2kplyVGZ7cRBKVHm/NW+E9N5m5OdMvFSjDdGAyBKs2Xu80Rt0tgGI
Nx/gVjeJjjHNBfFgwUHQoix8kFeh38ugGhqrUTH/FELvqGPXPkp35aa5t3uQEUiL
OdnsUENMu3VNr2pllUWXAT86KV4VTyVb4xwIxdiagKTqleQ6zSS+37AHXGmQINXK
FfXg0k0wpu36m1AUpanbDaPUCupiGJdrl/je4s75ubyBZGQvPS6gLX2fPYiUVD9Z
y9+xOXRPtJXL5Ywve/Su6lRgTgi+hpVoCu2nqBmrjgbNE2KrHbbTgGVblEcqwHD7
OlYBz2oujOwo/LfuhxWqHP2idsu3vMNeWZTT8H8GDdUrUCnTpiF6ki+3/jZMNdRZ
XX26hznFM9mhjRyvPsm8d+1S42jtFz1u0y8EUvMk8bM3YoQtgbMsCxsF3R9KtIlp
N0JTZjmdSaidSWLf56geRxnsgcOIS0/x9ATq+B0UQEVEJ/MdfhAxzRfTL5lzGxxk
d06FUJg65OGT2e7LrFUtw+By75qXvY8wRvbn/PMp1I4MLbXmWdVtOFZ5gsglWrAk
BXwQ7Z5OTd2ItAqGakW8C2w1Sc9wwGOdBkgZ/IcS9wMVMsL09j+8DiTVCRYwgWRB
EK6r6/BDgt6Pz3QopO4JxWXJkau7bSpu0r6jm4JtqQXldOWRgjd6HYHoVBJLY2Xn
TneNsUZ9hr8OGOLMi6tuNOpOk6nw3pDfca7uBEZCFIVXAunHd8Ai/1ai4XsuN2PF
wkoB8J13V6/h7ybRzqrfSurp1l5w/2opjJ2YaCprtU6vFZ7biLfr5+L9CLbVYzo+
5SCcReK1AcAq1lye+iV/e+Qvfy65K2BLFWOGesqT19EtD8FWBTPT5j02RPA98mJ/
tGPwjxpgG4UKe2bBl6SZbRT0EC+LfTWrHnDqk2CRwMjRbc9WJV5ZOxYwusmNMhLX
4lL5ooT3jK8s/AOyYKFGu3s8tPAvtTkTJH2W3HQJmApY9dKfZtlsPUZ81DiR3fpR
MSuxwAs+stbX/c010sBJFBladVhra+ZGxoesm3ccz11QwikdzpW6HaCm3aELv2mB
JPhpPhKDrhfM5a1Pl5r23iUUwRiyvjPcxnNVA9EvIb0OZTNNZZ29ex9KJXZBh/r3
dJRjytrRrCN1okw+hEjJTEyn4FKODQuLR9UAmh0pZEEzG3vi7TvzGDvdcJ8rHn9J
7vHJR0o8udczdMWbG+bDPGH+MmhS7sAKquictTZvBnSlYUDdwg/frrSsmOqFvt7R
ea1S5JS0XMqkWT/fwF/hjY+eB+Eyu9zZdjtuePhXPYgN+eT1h5CIh2cFCetn6i1f
CELA3KF7dO5ShAepczBwDNx42UsnV1XGpDVzupmv5nvR/+KlGY8gJ9ZmsWOe/cco
xymcLWDFVdbJoXEDVtSIDZszbgQ1ByVysWsoMcji1g1KI3aQnrC/76tgcqDZePn0
BfAJNPS8PUfqcdCk09rddj31Y2LqCK3+X62HpXNLszu7Womqj0FyZJO6HK82FSC3
0VoY4WM0xBY7LImpTR+xq+itp6SlCc5bkB0f3mR4epDi2Rzddj+PBsm7KUpZ0m7D
mqNY1ZWAETCM/YbUl4gAkn+JzpvisbnV0oT+St/mmCc/Y4MlUYFLvGmzfmBXdg8u
U9+ChJPJposXB5tLFU9sQ7UaK6SYhcpR6w6cvmjbpEBytvsIsVgJp6SYykvp+TLx
hk2oH0FMZnCbz6/fF627W5gZlDLx5v9kZAyZuU8j5WE3YvSrBp1ORi1yBniZwtMX
///yaVY0cpRSmQQihbHIVxsQsbeJCRzEWaOV7jAFcQsptistBKF6Hp9ZglEQtSgn
RLcsfcb63rDbAqkKclDRjzdPY706qA51TAWvKgAY0XrKBUbACYEheFsQgt74kyzG
dmI1d8kojuFkEl+cvFP7BUE76hAucSFITv6rkdiRaxWjUOqMg+vCtf5JCc9FvcuU
2Po3xnprfQKmiWXexz1wugOOg/Kgc/URQOGXt8lwfyCtiIrJIEccr+0jaVmcXaHU
lUL2VFuUm95k5powjWBPLgFvyd4sHtcjxsTmus+1nUFqsASkOYMyRvqNGzeF41fO
rgB2FyvETR2SOqZmszuDAe+yvuGd449qbsy6UrMUEIYzgVF9ef2ioHL57IDqg0pd
ZAlmCweFCCFlgB88Iay+Q0EPcpl8LGJs75AAXJGAJzNJJ4pRskLgyajLMi/6YS8H
FPnAuKp1oxFsY3ZX+jm4ZPSO3dvm8zRDMkt1/CoEVCrpW1GFrQOcoYPxx3exwUM7
f3ZY0J9K/UQZp0Bjg+YkNbL/sUC21z7RCM6Kg32Y+lo0BXS78SclmTnO8upPSNKw
Me1+iehaN5UM1QpgVsB8QRH+fEyF+0gCedZ4i8ZHVebTTzbiyu0M4jAo1cfDo68Y
zBd3hiN/LojdzdX3iCvf/Yc1ZGH4UxB2n6IfPMoe6mt3/ENy/I85XK8MpPNzDq4H
tJE5zabSfer1HIdhh2aP6QHyopUNAsUFvIJqU5JX3zYfk1Q9DCoys7ubAfhVnycg
FBsJ+GUOdjHc1OFPezHLMkybSAiuY+07ACJYvAC0q/923pp4tnSRDPZf7T83oSQ6
jLGzssuTH8YYzayIqFOxKWulluPifM8JXW0VNG0+/rzZQHo+ABPoYKmQUSfcKmB3
yxLK7KuNupeECg6S/k7kt/CzTutkbdvj//CgZV9GxMvsMAYqWx4DatcjocehR8Z2
A9BgcyloVOojJ490poCBW+u5rwVL083Z6AGr7RHaauHKRvjXjF2aigvsI0UdEB06
k1hLghtprCGvZZ2Mgb4db90sifDo3qxCYNCUFKWC61cC0Fnv9a5+B1uR6fdhpkSP
/mXKtfVxle+1uk07D7xVx0vq76frawbzP2glQwDl/2aV+l91POI1b6qJCZBpSeiP
7eOurSAK7SuB35qRqY8FnL5SDul/4eudMhnJCX0rUklW1MetD0fF4jTVFdqOYPmx
nvn8IrbjTrwyngbHT4RWgY+4bcUgNbHJXrvZJv6sB3LPijxRPavRqH2fgsmiZwab
l1OWkHv6Y7U1LRenR5CZNl7N2Fk4PqWn9bbew6QdxWlc4j5AUmO0wqgkoTx49Ch/
P9N3tNhkVc5lotfXtui74khKvZbtkIjsocRJRLzy6V6lEr12VEJrZo6+xfS1iWJf
uMPxnj7/D6+pmfbYGIpjml/+L1IUAcHBVtY70R/h8qX1IVxD56lTEW/yNrDdlUph
wKdg2dl48d2Vm4HGa9HTWHYyl1QwjFRZhmBBIlq4grNBC1qF523AahJUnCGG0MG9
wfbqJdeDjOJfIZW7/NFq18GcfgNgcsm1km7Rhsd7TejZXfkWvTFTwbdcaKbo7YGJ
REVlGjeW3CjwMPoS24p5ExN2jrTPejQI37NSPyHBlMcSDgmUvis36h1LCurBIDHn
QiyHaSSEDliMfkGAr/WWyVVmuqaLUXS0UEPLcW57uN2WbkOrvaL73fRlSf9M4P3V
PemIEP3HmSSpV2MDzSM3p6Wkr1k/hnmP/EGe2GqqQxfed0zfkyKDViiEv/QKFi0e
cWvBq7DibWN4VeNl70nf1QU77vVzsayhoSM53pdp2xj4wgDVTkgisrWFRxky578S
cfhPESYq9y+DaWL6ZmJgDlNmGCKYmVtpmM9ybtIYSqWBxy9rIN/dw2EdvdGlVd6E
WkJnJ+sOLYOKQEBpl6EhstQcQGg3XviAxX37YvnN3WuMILvqnkshEdeE04bKQ/Py
oTrHTMGZ9vgQ43u2kb3R6Z+MI2+VCtyjv8TRt2/t3Z8IlIGtNle0hQwwzv8y103V
VWgEQIZ6I6/GuU0o2TKTCR0Mer3CjvWbU8/csAos7QOiPy+GN76jzxK2HCQUBvp7
sjOynJsua0y9eKx4mEQLROrOLE6xh9ms1p/VQwjwgkeXKhCZcfppuD2T/Sr6vJq8
PDidVlNoUtRpdCfPyEoIr9M+S0c42zlx2Du6cZ5GtFxMckeoQEFaDubBRhCWhZv2
oe9ADH8syhXcNfBWKGmFM4Jaz9WSCAey7txWfbMvTqFkG5GNCdlOLnekMgeHphJx
heRSNqdeRdLuNmF9exVKKmTArGA7I7F0zT2rEXP11WPrvlg04I/UvKK0/bbEHL65
vI6mnAWFnnifa38iYQCnZeX6KxVOziGYT22LDpph1FjCuGcp4RwemPMmAAQ5I+ly
u6044I9ENFdTRfKrd4hZU2h76f6aC5Tb+FwU3f9LN1e8S13QgRm7BkSPjeetp8TM
V9bld9NrMHVcrxkrBetfi2VTSFLekoYz+pvfJVaE99K3eGQa/r1nBTbVt1jLPs2K
EkTZRM0tCKQid3fEdG1dC7M6FjdhTfJas/M95+67EsT5dmcAaFM6vH8B6YV24nxL
VqJ5sdUNpgucQ197/ZVoJugD9uUlRb2OYSn52iDOTG4B/JlF+FqQH/wTQ4wapRPN
X7FFtrNbMIvo305Jm+rgXaHuN7Ai9zMU+epUHPkEOysWL0J8/quPsg7NwvPwuLKV
Bt+J/q25iLoR1Nk7jG7W6fr56dbTgmHh6sgfsKnl7JXee8otTK8A727ooMpE9k1x
fTma8Zvza6mmIfBx34EnNAcCznD0MdyJeFysFIruwMk6kKT1f2fweNYnPpxG2SHp
KIniEvVpVMDy+8FaKe/nEhDuzsKtRNw5usnFDYFpS5P6BXaULLK9OwJdvncRCCyy
xqy5hVTE86N/YifWsRxkDH+gYqsV/FaQ28m5foL+jiETiEa5FuTj/slS8+KPCdcp
vTW8nGGv4cTc72jYRwxF44nRwzFL2QVfayy6c94pbvW/I8h/d47NM4NsceTsPd18
Pr8Gr9vKinEUD5PkAgm3T1R9DBfxvvxDdxZ85OcG7SGWqEDF89ixsot0xg3APl0w
TCRYoS7CYjCo/MZ8rbmgmyhsHB23slPB5NUITUvVDLEAed2gu+XkOpi17ztkNpM5
+dQAmAxs+g4YLw9pNCI7B9bBljV2g3QvdkvK2WNPvyOovQVPYaZjGt+J+fXR8rsC
gykDUEWq3MrodPzZWfImmra+PNEzn5IxS/1p5X7Xql7fnedA/elMGc9Poi9JRrXY
0juCp30SIzcZL0bVSnqMwrmdGrTyt9jSMfnpRbPOhKqh5EhyYh9lWwk2k9gDr7ci
GTUIfMNED2QqxG6jH/kDU/IdsH+ZjuZEEBPZBTsYFk953zoYZXIS0pGDz0SYz6RM
mIMD/g5nhFXt0vEjGGDRcpOBxbxHhomrNO43J42GHRDtJAROve+3tI7B9Rbp+kQ5
9R6ml6mwR/AZSsemyOX8AjZ9EOwHrD43b5koR3zN2MtNMOBzUNFkAtcnHOvb/DXh
yHAwSO9EUVwddmo+cRVVosFUby3jl8AgM2VcL2jro62QQa3P1gmAILKnnJdkwaac
5Xp6zS7OR5vZpu1Xc8SPmVapaC1Tm9pgtCtQyyax6El+Hc/x854V3Kjwz1b2uUoJ
Zzo96pD8JF1Tz8J+31z98m715fTQ7Uq5D7TfDxyGGvgmWuTrUTvzzxquE56/HBVO
E/2wBdIOwteouHrFLHl0Bdku9zBSdA3F65KGZL0YPgsp0caVM+cv9cmcxQWVkEGi
xV4QpLKeaJV4k4N2IHac5xvr438Krcf0XiEXRHWq7LsChTAk41q7lS5fDBr6Dvon
VsNsLy1OT3CDIH/j13krNNmhfMkw7HUTHEqoJBQ+IM+bGrYHdhN8ZC0SXqr+dhi0
U3pOPUSAMn2f7TEbQqMnQRCR0wyoXHmRS8ZkjrT36jxk96yuvDSABHJ1NLxqp31N
H9nSsrLzdanllxVByIDTh0uHMOsb07B6lcKaKAC/HVS/RDONaXtzJI77sxwiiZVW
6cpFxz93k1k4eiMNeVEYsuaY2mePfGF2wUkls5/gPiuDwSgfYfPKLkMDt2XgrSEE
Lk7xUx5hifZMT5oHyvFx65UXD2S5JRPtCcb9ic1tRraMepZf03BQXR75bKnNMjAC
E2XelJfuO0PSxpzx63n9jKKBoC0/FO3JAKkIdRSWbzjb1d0mlxbNjs6FbCjn1m5u
O6b61zkzkaegts1PPfgmzxmSlXT1wvVocFX9YHeUrLplWELvjMGgcuAg3giMVyQc
mCrt1+f5QZJXAbMIR/a2rooC/WgaJwGuBEfOkA5RT0VvxWbhrutg00rhlXQjkmrf
S9GIQ4jGOxmJvjcF0LKgAs6ISqYjKwgETkWSClC8nPPyclJw71hPzZF8tmmfonu4
PgaWgziSqUSqMGoaLVdG68/okBqhtlUGJfHeI+ngtSE4w4bQT51VqnWRculDrG7k
FnNZbuKIRctUhPdpAHaSWsgL06O+GU6t190OXhkx0RrDrTxec/0Ef3hebExlgtIt
x7ZFmtfKD/mdo9vo870H3xwEsqPhe7tArAWoVucEHJ0oQHPOw5sTn045is7P6Jav
O1byJjHYmCEabSk/Q1eXalo/j2OwzjvlfzCxicWyVivPiiSbRauB2qVmqcoGWxlS
i0BYKFt8Z1iAXN28RniOW89Gxi5aGpg6WH2ZN1DgqcDLm/rotd9BYQKfg3caK9tY
end6IIY606YBLhhZAeG7OxCbdVRGpQF97wZmAjre+D22KMCPUz6ERaAFJaG08KZ4
G7jEaZeIdtmKK10KuTpKs8BUCo6v9TvilBgJw2aFsY76LB0wsiekQ7caEQgl+Hvb
oLxp9sbNB7/w3p+LaYJXiQET++zZLfXdsYDQ7KLATAxp9mFZ4HUpxelE3xVtTWW3
bYTOK9b81KoTDP+wrm0X/caJQqbO8f3WWOkjvTp+GwY7VggxTPq5dmg7/HWn8/I1
gAmCjcsPIlp4U48wrkpQdX+QScFCQKxO2htNVSNaZOKeTko14LS5L+JP7tSeqbrp
/Q55ZWaW3g4rdaUdiHwfvg59aVjj0cBMpMWh30KRIG5gNR5P3BtQrsLlLaafBRg1
nMq4j1j/14awApu1Z/yQQcrj/VpQePL72T3J5UIucRFTd1N8DauRVExJea9OARCg
qxaqiLFbfkDQQIvyXdm0tbbhKofN6+WI485/W6pu/yd2C5TYVq44EvexRTRIEP4c
pSKgx8dS+xNZAf2g32uWva0dz1qplcxQ3beWnqQOeiee5KnuO9EAkepQm1C+aOR/
7PTiMNbtpxdDsOIL358OopGJZtizNE8f7Kz1KDCvC9lQNrQM6xz6bkkMINZNi0/U
wALj3fi7l7CPzz7tU5C6WStRxUp7cdKPP7jNoLOR+4WQHV//gWxAAmQIf9p+e1jS
YeJeJWRVoLj5IW9lpCjXFzs6krdSgKIIK1HOJSqWaHHu43wMRb1EVVbUvEyDxPO+
rc2NXG6eRhMzc6h4C4qNRBhYC/tB5bt+ytg4g1HOsh2KOXVydfJavB2rjFKqiSXC
cuXOfu7CeIycs2LOvcLuHnAMcQtzMOjzVtVbPheHTTaGBSrjmb3HYyv92+3azcGG
vXDLpDokuadsryjYjzE1FFNZB7Qa7SChkWNoRLEdzHEbUgNeXzeDD0RDTEVHNbRZ
+NbV8DtLH/zC747XXQLrTFubiD0Zd7/z68ySbNuteLfKSOfMC0kYtmwzY/vTrG2S
T36HD4dh33Xjgx28cdQDCnogfWTNjchW1BK6pqUaebneeIKjjS8hFhhTUuo8zTya
BYZy0YvCInAfeKYux4VfrvXVFLxqUZHzYku9Oaqm7ThKWsySWyOh4Sbf8DbWFk2R
euI6BF/8+EzE58B+Y5mO7fUOO5xyOtyojgcPSpqDU+kne4QnbWTi+LJN79wzooQd
RUGEeEtw8hIsvj34QDzvhP98AQ/bUiMICXvJ6YuDKAAYvK8qM9VDi92H0yTxo5np
acFA8clyLTM7PJGEQeAk8g5GjM5SFp2VpMu6JoIH8COLmLdQ74PTB62tY/x1f/+E
YHyFi7bge6exa6RduGDNQ/NVSvw2btw2XZHgSTpPXACbWQvOFagnSvq24Vz4KbtY
E4iy7AhFs9jO7nxmWyqsnWsFbMQ3MtG3pVymuoBJpqqGMhEZu4+uZsgCD7yMs5E1
VYPGMOqPVJ2HneoQc2cHf1bDTL4zR8bKYVRAuverW4oZe1wR/T0M8sKb6osk2e5S
3LgsWIdHr/FQDQXEgP9mdh6zxNIO63ixuDchiEIEg8cPxrSwYlYebZeOCxQ6KojO
YB4YbBe2m3cW9gXj9t8Sws24e4BtgyUuJc48Fez5CvvX1I5EjBAJphAu5F5WX3WX
FV2FDeqdmCWLZaCcfgJMEamTNhdlIjDPCxV6IjuQ0m+5O8ON97bKUdg2A2KHwVAc
AGmsLB/UUop1CQvMHKPHzD8FLHXgxWKNOrZx6C4l2zCFjKfaO2Lpk0wkDInGkGFY
usCgPbPeG9zqsFffy/FtaoTYIXG4s53Z91vKNuGoo1BuiPa8Ki28/JdRLIEvIaQP
+Aa40Nxyibkq/XCcoBq/ynPtGl5KHk6MUapB770npgCOR725B18Q2ZBd3csRY0j+
l4GYcS5SFPCov1tUe3Lb3BmIJj/l53LDzwCQPXjdTqhLXwLAKi0pkzmxZLiRvnzM
10J+lWmcecVZFsSpCgRZT9UHNoCPejt96H2Tbm9UrNi2SBdJ1/zBEvngkW1yJR2M
EZCtBx5soeZAjyVcvoVVOaP/BhQLXtht/Zi5dpTBtrKlfzBnZMP5BfcqIZV4sBbp
9uiub1ruI9rNwtsj6jbZu5v0QfB2mbivcv9yPqjeXV8SX2myvgg8leirxInDiT36
o2vyOuBcoEoiJi7ci5c2HSkTRWcjrVSTkEqQByC8AuCeJcqnudwWLXsYhvJJm6NB
UFrsmqlWhMaAAK98kmJStTNnr4LFlZSgXSExICJhKSh0zSpW7UJUgVRzmBk1MNnG
2BNuWtCSu9MjN0QhlpfmLZdp3KgkO+mlDLzqngdB765AV/6qsfBpHoTzZWctq5P9
/zWzmmoc1gJhBNBKikghH1fo9KK0EoDe+PSCIVhHbgaxZifvdP1gcKV1iRnRcFuV
gz8KKKV38pWvlGbMHyfnYln4hvZDew4QgzNst9nO70Y8IFPDhwWa9jWC+zzP5skr
dXqTDJokhjutbC7siEr/iYacgYWQKeAYTwi1wVlbqQE0dl/1V1oP7hVxW+tn1zWR
K13z8yl/6eL0CjfRcJrHJbHP+IMMQ0Ju7xIVpOEgc/yPTjnfiq39EGnZOFMdlzdE
EskVRFxe8AhNrBF8oDwcS0WXwyusngRBLU15HaTf7/kGoUi5CDI9a3DqkzJQ6jN4
NYsa40w5V9TsUwsZTigvRERS6n4h/kgy8qvOghT6r3SALC/cojn3yueaNhZH5n2u
9Zm8BY5Cs/AW3lSa3Xy1NAOja3As7u4cY0pACc+nZ7J7VuMrIKCGNYIKnV7aq8tJ
6qOdfFZXz6birdNb7dZGdKx+qLsilu1lKgYmwQa+XQrh+U9TMUUqV0iOFfNJ51D7
lTO7egy43ipGSqo4z5434MaNY3Sd9D4UkED9C0UKA+H9mg7wtDfAlgs9nYH1MaP8
e4qxhRFmvR2dh1NmNWg4wFbLImTJw4mqiQK9UkKuy22vqDtRQHnURFarjvBqSnCV
HPkDOdTyV45jPGf2bFYPZMb5xUfZ8MoRPqOtqg8a4d+Pw+lbcjlpW2ZfmXBYAF5I
csob6kf6EDEz2PdJZXVR2O9BQ71b1Pt1NIw0X9TaVxlSkcICGOjWc2oSZMkbS48r
qa5YEeUogJHNHRxNaRZV69j7NQdV5QHi/yhsS6NXJyp+GrOz3HEk03dRWZi6t3zU
Mx4VZLj3WXxK/hg2jEVxDV+vg/nOKN1A/IXyQ9gOAOZEvV+DU5RKQaiVhixCLayn
Zpi7Vh0hhBr8Zk4LT7Osjjgj5MCT5Z2EqePN9ePvIomwXNwGpb8Gulybqajv3E6X
1kBKuJ9sqSyhA6k7wJlXRmwBdYyu5dEUEjJppDmI3zj8xjG2OMZ8Te8YbBOvPgA2
Kuf1p8yWx+84I840qBClPU37aByBa/vXJ4Rlx6EKEDwLM+iN22n7ht32pts6wBqx
zndvZpCknddh871ECIzr4w1yDPjCsOnaQ+EE8RYP6oF1R2S0bZ2ftnQEXOFJx4Fn
Tk6PncbeNZeXEop2X6+nEEKZJJDmahyw2QlDvuXC0fdhz6FD4XkE7IFlbksI+qS7
Rv8OSoy5C+xNANP4hbsdkU0/76sSr1hAistJsagLRhgYrapLBoradV6U7hgTUx9u
IZF9kEIVLVnSgfU/0G3LppPTLciAnfQYUwbE17gSqsts3HYJJK02Kz1YZ53Qo8l4
rCsXPGQPcaMKvAtKR2d1NShFvMySyfdywEdltkIsOOZ1Yfw20Jccnk8zNdM+gE+F
uo0Rt2aGKLZxqnEp+ifMjuUtarOKBbZYIkj6ngL/zTJPFYa9zfNEaomUMkWjGnFf
ZEk6BYYkpR/1sdHIVaL9VvrHDssBxRoTDHmoDzv2rfM50+rZ+Es5KldUeHXPOmir
CicFu6SxnYmPlVnSDZYJ2fopcPB6s0ttHcbRGLsL2cNEsujWsOThi2ek/V1BSwJP
KYK07+KAvtGl6SIh8LT0nuy5YuLv4cxpZ1mTABghfkQv4LexWCVxT60eO4x7FntX
9E9yJMGHdjdYeeysvrD8jXupAx3tFtjbrbWIjKxCNceaIaj61a89106VMyN/cqfA
uSOmANb/D0+8AM2zf2m4yEJNF2erNziDTrxqwILAPnXF/pRr1rufv6ztBNLI2Y3C
M3ufkX8A6TXn0F9e8ecNFJ6HYBAU5KdnlrrUdoqr84eMmQ8MOqTmn79S82fmLriS
REiyg1FRje687oS0xY1T+hQmnR1bnCp1BwAnnB6xnQLesdoEMv/vYcfvimp5YIIS
9WIME90S49bLdU5Q2v4jQfT+Cdh1xpUEsg+QlqfRxFIcrLA/JoQTF1/W2RuVaPq4
ROHVAlFH0lyPnLjxn3x4YVj98tLgN+6ZkfKyB1cmtmHyOYKcK0cM7ZizL72Wl4hS
gsr5jxJCceunvLmx/lXnNLdKtdf6DA1suWhqAxp57VszcVa7UluWvJ1h+ZNFTmXE
ef+ipXkYRmQafJyM0vTP/LTHUCFfDcbNwI/hfJmCUEJiKfVtUW9SY6GYJSjmo0XY
k42SkFOi1Aiu4NnZbBa6PkEGAsJ4P25B7hEkIAGD3SSnPffNEn4o0wHy3qE/orSb
CGEpTGS64WlhAvJgBoF+BhGW/oI+lj4PA4jRMDIim+oQYXSIIzKJlaIM67kggUN5
lrfXFVOxmo6IDmFyXXkBiG5BpzbpvwlNZyctf90i9y45LyOmS5x8BkUoYACsGFkr
TJHj/nEmRuu+7XkANXoyIXLwoCYeQBZWv1EqdNE/i8YuGA2oIBg4sGp9oRDgHaoh
jZFvwXW2ZkSHCPN2+9j43hhEgmuM3Jig2ejpKYTstR0U/6g7rfW3FMgnvy4wPWEd
5chR+gjRKW50i3diGtMnrZLnseZB+BvGF3P3jDW9d2OlxyfAUUDPte2hq8BcYez3
/88LFA3bbd0UCLj8Re3rNIqvMHiuAfeOSBScLqjTDklzAVXcxuUqcP2PN8dh+QFU
08/FprYnPV8kKFMvXTQ+aZ+/YuzQ2R+DY+Oi8h3UWxirYByg2dV2YTVAfhz/d6cz
IflAUKXbhfJiAyr8wO/Bkw5QYFlcI04Hh/b+ztwd406cMHMY8uNDmaQ08m5h4p+7
TEYZNDEPfoli953keCO1I9emRZ8NpxkagZO5LXZ0LRwELHirCweBiETfwjvrr+VX
zsH14g4W5huhAhEu7teODLo3fcr5xApUiuX5qbqW0vl3KKnVFoU/SYg+1LYSZ1oo
ipmBMQhLAc2oHxq51iU0xlU2QfeoTWH9Oj5lO/dOItdKl2BQMQy4rD0bDN+8YFhM
joWfsdyAbwB+GT0AHkGNL2mDYC8YYswJ5Q1Z8jr7kl8PQvcu9WZinun5ZbPWukxD
0sPVimYU8vpGXfjlhKkhGB9nQ87MBqmtiKQpRMoCfxcBBns5PCkIl7dzojCA+eXe
Mtoz2ux4qevb9Ko51ayvCKv2MQIGS8gOApGzg745aZK/AmRUNxyBwwf/CrGbywPy
8y78uRAvacHr2S1bUH0/FNR1hGaklPnSBShYXHPvGWfApE87RUL3e6wTmK+b3MhQ
oKZf8A/o1EZyZQzvcCCB1dA0eSGxzypRbeTCLHKaAVTOwBZfPXmg2ht4YMtTY6P9
Ycec0eUwMwFgU37VJMkg7YYCwlJJx4V0PHJYwin4hSYgAdEhQfU3HlfaIwA4DMqi
j7C9Tqz2XSM8bc3kLAYz2zoCBZY3MbBwruoBevlLdGySUPXMjlXEeG07Ilnnr5KZ
bB9Gb9Q0LU6C9+z2UfxiWSHGv/Ms611tm0PGRsspA2CR6o+LxELFfRwnO66YN+pa
N/bcR7sLoZtE0N6cIVubP6jPc/Gj1S2JhZyqsutiXjEQmt2ToyMnZ5HYsM46AoCR
uJIGqVnKgLrbdsSJS5bLtZD51wmHTBLDTdY8zMd/dppYBEqhFJCfNfiV4pMD4RAN
Iif1NeSMzGw2zIV79eTwSgV7nQshT3Y/2O1Wio74gNed1ocIlMf4bin/T9OOJFPK
ALUzEHOWM+dz2ZSD8t7HhZMfG1aa/dfxragwuEm4Z5nikpWtlX2hpf0biYY7z50S
4l2GlGmOnXsEaymzV33PMHXNFA97jsuuh7ybqxufpW0QHar9CDbncIAxgOPatbFy
7Oc8MsPTHKXF/VHWXsylW7xJzocga1sObCTexWqk9NkeqPy7i2DI/Srbru7HXI3J
bW7rC5BcQ2Z+BmhzWRf450aPbYsUwnvtHxnSy+Ue8L2estisFgiNvS3goi+9ke5D
4TaxnyAPKHd8tytdOhElHAeGG+SRlSnv9M3I90u3jnN5vamLQmav7sYtoDmDKxeO
XwyHVbmO+jX3mxlOGxpbbnl9Z8l83yTLsUYJd7XRJwQ3RAlfU/vWjv/+aUu9Xknt
CeNzeoV0vkxZPvK6HG5E6R3quFYl1NqW+PNov11y7fit5yM30zzhFLHW95qr/EvW
b4hblsqjaVz3kLUgzdhxBmCeAdBGQF006eWZSiN0wxzdAXX5qQQhCOcexN1PqZ7b
OAlCKJfs7pXdXIhED27dQhL2H1vF+f1zNTnV4bqSnuVp4etixvMteDKDJhcp7x0N
WrrGAx5j6oEk9m2I39xGyVnXNJb2HaixxtBl3/eYUA49RRux5F9Drp+IaudHtugk
EN66amBqrXgmXycCfN011knaDhalTZhr/CSmuJ8AI55+uusY2YzIkcsCeWD9FLfV
+Ci9LK3x/2neJN2DKea9YxUucjbDhDtMxSEh8SCDyDefrgj1qCT3fQJTbtaQfBiu
We9hZ8kL5+Zu8K2Wdre8a4QgCaeCE1URVGhVttGmM+G7UyEkxU06V/83rB5uOjMA
8SJPUEGmyLhTSlc0wPQXnAnBo+g/FANLsbF5XUbk5HCL2ozwFoqiHn4epZbQqXSp
yNkvgpK58EXojUrTnwBmoQx380J9I6xMaewbBf/y0uGo7aDYgHymtPS/pGbSthxZ
u1PUii99/FiktaSbKSB/EJgOa/ZcY3TZKW7GTj4s904FyuvudKxmi2wZ8r2DaB8a
/nkSN6KSe0b/xHG9tWSO6AUXsTtc6Ko1OKu1DUnYOVqO2M3h2AKgYgj8eJ41iqKZ
AvJVyv2dqrXq3r2Ccv9V1Vi+BEZtqS6m7TflI2IStLiaTU333Cn1xvf1q0teSvWI
GDXME6oqQekzWesnavAMREDoaCNIfOdhQfVXdLoPVSK+MrSOPDcmVDo3dnuKDRgC
rR/5fhwugfZvkISDWID407Q7sj+GlY9QyvAAS0Km9TZbSk54BSuK4Hdh06LCxH38
BPZbIjq6lPhXxymbp9kZ4dRWHGU+pbjAOU7bprp9eFbDVgfc3YTGcA2ha+Z4w6mw
nU0N0qIXjMa7On06C5m2ies77d1jQAPFbvDOuNwI6h2fVMqicm8rrgqEPFZZmtAt
HKbq+/QbCOjaYtvB8qGDOckWBC4etBh2qGC4hfiPkdh0PDe22a6VUfxhzmD+TB3R
H24yJIUSlD4tXCRC++v/eqxte4/YIIOR0Armrswrk0ShPYEBe1DBuRpY0HIRCWf/
aifLhLUgZ3dhksmEEA5+0tVNOfBp3D6gb9+e0as/AkpdK7Vf58Z5brku5dcTt/Uq
+FILUb5yL1dANs0GIfm3SejSzGEK9HNfy/W049OpvaD3Zvrxtxz1EvIvqOi2d+o2
dyLhf6EydQk7kW0zfbBN1xbZ1GNu+OsGwu8CauPWojQtss709ZAbLj4dzBCgCZBi
VaWc0Z8ZI37DyWV7BULUFG0mMceEp8CifdjIs0Y+xbkj60s6fALavEI1VHP7wXh7
GsGqR3+A2zJ3lE+PKnWUPtBZzNCu48GeNPCixIZWVtlVgE2+qQ+SauDpmbd3R0DX
hopYPnu6G8u4SdKuxuU+pRNwknHA7lR8pF4DucrIOPDh+k+UDAjVMJdQFH5POQhm
aF3HzvRACl9ZaQ8k8NWc1fCQgRjSIyKh5D5tmJAg5RNvBJIIXBml7umqy9/3XykC
0ffeF9CRr68eqqjcf1SY7MDCf16/P97pF64Ll+F0JCq86nk70d5ZlsccA92a0QYc
XumkBhXZnsIk7M+Snbkyo1j69zru4y/QUOMgTnjIiTROyP3piiY38v4PcbS4CGuf
QGfFUCBkE6tFYL1WjRmGu8d0Bq5DcGoRUrGu8MpEDfywFPWiIlxG7fpGx6hEG5he
8XQHhLXoDCKJ7pjqTAjYS4e0JOU9lcKp9DIIkMhZmeaA0PKlJEbF5OJeUiL9xi8S
L9XodfC2gcrwwZXzt2qG+zTdVV0XXf7Y1AY7PKJ0seZ3ftjMDNKa5yYkljdQYbQm
m0a4LG417YBqVnyi2QWqU55sdDn9cLtdrP2Ek4JhfVcR3K425QG5wq7oNnnvWFoR
iDU83Galm4haCBNbeCm1s/Hk5yl+i9ZaAUJr6bgicfrdPLYIhDqPK+1yaT42LMW1
c4K2PzcVCcsyrn42tFyOlUbGBRj8NSSvMhCi3UP9YFQhXnlfX1FT6AhJLsxmoJ6P
BiAT2Xmd/jaHNGgDQZSv1U9ycunByHtsAibNaySLJ0QjUe/jpWAk24xggE+tE0o2
sOnyO9D60w0l0R+EyvhoBSZ3ZpO1zQbo5r6t2jxFPWTXFKss36TJbmfbTAzz4v0u
t2qln2/T03h7G+r5+MLq1HEVxJ9VwBWBBTTkTr8YrDWKtYwLOHgMg5pEGzgVZAJC
sh1NTJFC/PL1iuvkCnM2bGycsx9FvU31jHDJbmwuyvUQKs84BAjY62baCX9oqtJM
/gTT68z0zowrop4fb//MYioEmtDTtNXrnphD4UKsxnYprJvvZDX9Po9kDIDLHpGj
691HMk3u7Q+oCTmd8zJAc74ZPMXoJzYs1cvtk+SQKKFrvI9J6qqqokSSf8fJX56h
dJ3XA+FGeywDJxVNsyVJjxCzyG29haXrv/wm0LXpMYRu5u3xkJWkAiHK/tbeSMk1
wG7Ga71i+CJP4X0SQlqWTzDyXfF3PeosTdsbsbC8oOXC9Q406exhqWVSuwut3oU3
I9KNFmlPh9xLlc4Z8/tJZv+NsgREo+ZGF1BtiMSFQ0EkZE/YHRGwq250l2u8ldsZ
Ip5nEieKeRlQU2uulJJMr5xYH5ZGRTP9u8XnyXasxLTz8pLOTqtoFqYpCECyA/nK
SZDCgk4dvP2hP4NX2f+VHYOFwOXrKuF26qn4EC46j4iZQC9xt4RUNJTGI08yii6P
3COE2aMtC/Sk+N+mwvPHACAZA9GKvhCEEsoGJOP9MGBPA8YaQGim0FY4eN0OV/3N
2L36mCCysK02+cR5qc9cDjdm0E/7+eESxRu/810A9o6barupGasxfstDdYeDTUUH
NumT+nNGWTozs8whnrbolYLyOfCpFfeg1o79SxHbcEKRTBZ59ncD0J+dhF/OhjiC
/PwIaZ8N/0bKpGJkTrqJq9hM9ZG03AD3j5faSLA94SxwaN3axd0OqFnyzNmNcSxo
pwNfqm6TxKWf4zr3CiuYBibiquXeHcjpdj+/cE2vcBfZIHxoaIgHbqaE3u44S8sn
o+o+D4f1eywkzVonqxKbW6+eBsLTPSR7dQ+nb0sFWwXaZlYwFT1BWJLAHCUwppfP
prsd87AtjBU3Z0hsBZrboITSaE+J1MwSWy47aiYktx6OhairoxZ+iakwf+lvOpnW
fDqafJ6qKx+5XPweOl5Q//2aS7EhfPYh+N6Pby6FJZlgct+P1PKl3urNSF+V0AqK
nl+A1AT9PbWAiJmQHwXQKqQeX4i22gCUju6KsHKOJxMg37d0qs6q0++olZCkA4FV
3geqceHGmmJP2dzyiigCQgL007CIBnAoiPrtMzNeNzWrokDUCYY9z4VDLl6aGQgY
wffb/9cH4tXcsYIZdOL6x2mOpplcCV8YlTJwJRZAL4sn+Ia6kJd0IYhg4NJI2WNP
mh0U3czSusYlh1e76lUmoLSodfEpkA2g1Q7MmBf1Tzw90jjIIbjYMbgvUe5NTkBn
YmLuZpRm7wl2TgyN4X6tZI3MB4fqzOegNXBazMGzF/XZ+XRZTbOazfjs7ZxB0qI7
3lWxrR8B+WkFoyYK7GpBDD9xw8DWPne2peTK1W+2QWqqEHhNR8cDWCriMvZGUKE+
AIoQLjuioI4r7mX0ubmNFQOxy8a7jSmu4qvKcC9MKD/x9AmF4AEE5TZACKJDI9NG
bAEPLQw+gM1FFjvXP+JBF6B0zx4nnFIqXw9HX5hf/vYqbpqcQh9bJFWZ9dVZ4ZO1
wD8wx9fhQuZS5popr4KFJ3JpuyAVl2oUzohCvit8HQMoNTge4aQ/R2TdKJz18uLA
bEkqZasrLGp1jyS8sYvV3ZxorgFPEl8NRnaRdykA3Oei4Ko2VwFw5O0DlQko9YJi
wsnQ4ZBJeQqcPrGWIvnVjOvqlz+Nwp4+YmqeN9d0q9TQZg8qMoUApF3KRbfgXW6p
QzpMAB1V0hRkwPEVV+1z8uommnHLPwc3oly26JHRB4zptpno87/noP8CU0c/BVhP
iIoN3RIC8Pm4MUU6B0I2ztw4YwBTkmEbt4zyHvldpMzYP9l4nTGizo/denc0VJOV
PlbhvOb2OO0UwMMjltV9fAWPEIQ0oCN1FjD+sDrVW0E9LBrGSXAXyC6GqjE3LDdA
F848al69s9cJGeaDmc8S6qrOHSeQoyu9t8XKLeQAF1XrjP5SRG9E895L8Wyme50K
dBo0L0VrDWvy0a0sAMfDy4R/Z8Dh2mqOXf9p4X8brgiKfuMa9jSOm/znN4UUievw
89DYXYsdkLPZEwOFMOuua3mKMrrZ188boBlgiY6ctsvhGlMupJ9zuEAIuV7r5lHK
k3Mv9y+ggXf5IHt/SXjY0hVieQ541DgOA4/Fw4K79hyz4uTEz8DMf2BRKw4mG+Gv
P/h6P58zlAg9cVVe+jwNAPIgtL7KujGIASK8PAFtLgXyI/XNaHS/MOauB1/LdOgA
ova7Hz8ZE6Dw/+0uttj8WZUkUuJA2huOKh7l8Ag2QKr2R4gf4TLAqDAX8WnS3LWR
Lnope9XIVT7Ryrd6LXaKpVkHNHC5LHYEgwgU3AKSSUr+tOtgtbZ2hc7a+w0DWyWQ
5UBPAj5PlNCnpFevv43O+r04LN0HcJNjzMJ+fKavAyi3eGp5nTJIk9eX/kmS2SqS
fkKlE97fa8qUrlvD4O40Zoj8AH7zDS7AfiUDtyKuLsxcUDeiZCt+3CV/VEhkjIae
cRALzVcfH/81U8RtEzkp94qd3E3C1Ub4/X8N6cFfbLu7s4wqf9k3NovfelAk2nZn
LSgCSJGlp4jd4/6WvBVNWmQ/yNpA2lWpNyWVNGMD2SzFRX8kQDqmHv4BVYMwn/1/
pNl1wg5kNyPBxM77hc+HgyQpwcMofN/DFg7xsWGah4PqFdxQW45VAT/5WtXouTRu
Gez2ozQwyCzw1uk9gbf7F2erRW+B2IFlKFG1HrHixR990R0LgJf4yi+bxiuzuQr8
16GuSfHtDA6FwwizEYwLp9AxK3DpRorGKF0OBF8gkkj6fuJsQpwi4qoXUSkOTtvZ
+oE+akOoM5f9Vka5jfd9hS0d86/vheczKqhRBypgy32/dS2LoGkhfJs1BlwLBoga
3yPrASMwh9dCGDsvEzxxTdzyTBybRLtVSwNnAwACC+snxKRbkFiyVFixb3RHVmDd
FiDFE6fVxOyNVv/FQbKRnHSbX2Yo6FP3kF0zP2XpTjfJ4f1aWdrqbnsmgr9WeMUo
d0fymiG1spD6VDnigD9wjDhei1ROcFG4Dl28/+S5XStHPeRAxw3xSkmjjk6wMd34
faPESeYOGf0zyZdZOR/aRXKBg+iNmh8uKdCHZfBsiyAoEOMPHyoQsNUFoP6l4C2q
8KipIlXerrGayLnXsMbwSAQhJobPkDipjZI1Okrt+z+AtwIB8+LVrExr0I6w3bKE
Seid9QxdPPBHaJuIGPzsN7QIRgaRxVpKR3N/F5Q+03q4zOdjq8WfK3HKC3tZZJkJ
2+jZdUwLFuAbxT5s3EC6V0wX4wOwQCNSGWwpMzjYtAGYhowttDuYq9TyU/d/+OyZ
EWHvDCP9Y59Usy++DtIzUk4NpODp9ZanjCZEihflKGJS/zS5GDfb8coEvDG31PVA
fUt8XPVi9F5UkJ66UyxyQB4vi/kjOtqhoWQJZvl7BQLojh7BWJrH8btbZjV6BbCX
Q0zJ3Bsmo2/IoiueAlJgpswEvqlnJSfP8OA4iACKW98goYOzsOcWr33SvY8RrT15
z19bOLSjt01tJX+tKOw+yRjD3GXH9i6Odmo18dqFvbQzrha8r84NNDa2FwxUs/kK
T5xowfjeI6G3BByEMK0oaCh/6Ihp1nVub9Jqk44hGEDaO47WBP1aApxuxIscaqTk
YAIKUe2B3kLYXNKFqlVP86M0KPqKySJhgi4l0NTnhLRl4nyXCe9tHzad3nVwsM+3
pec0tt2b6eMZSItXVJnGbECS5yYlvccMYJMqfjMpQoyILyyC4+C6MRyu5fwGPuJz
Vct9b6XByM7g9u9/9Xbur8EStWJ1xnOMlpLaOu354oP6qCaJn+OnvTsc4iytJClF
G2bhbf2dBzgWnwEWWdIeLStaCwhEUQmB0xTXOj9C1vllUoh2brXShVOH77vJoqV7
ro+IkzIhHLt5lrsNTkzo7uK2Ugjr5+bdZCUP9btZEi1hoBMXBjoTaEvm058aiQYe
Zv5jMm7wZ61QP9tSedW5vl9DT4iHbUZYMl4vLylltLl8av4weGDlKcpcNEpPJdk6
i6U8S+sdI1rXXG3zk3FNu6uGakAFBAinCXPhAB4FMqjGaqja2XCAoovO45XpWjL0
V38Z5dXVjxjyIXFdPI/2MVjhImVne6F4Gvzx2kthOjyKzuP/p2BFs2EgI8j4Ybvd
D82775BkdliuTj0QKbIo62PLOmiOJVJAqEkXGeXTfz1bBgYhHlp39ODH9gjM9yC8
kCA26WLOjIWQMplygnux1uZHk1WV8I/p2qQSp79zTsZQ3zLW2x2jHhqhp8UKKkXR
PjrYXdbGYhaJVxfdS3QxnkwLwWTV4cSPMUmbRDs348afORJsAB7Mf31Vt3KrG5y2
Yk/vH6rfVcNVliPeT7cbJGgCk5ph/gBwGz6+OvhWAkbNhI4eyZAvt9C8MRVBBbQI
NU4cuJSmW37Sh055SrK+1pkTKtaCSPO+ZLcRqVkcZcDxo8IaYjsbNsc7gQn4qZs1
xXYa+X7VMqt/aUMoBE0R85Wy8BPvT7dPKXxml3iIvQgVVNid5E1Z+mfjYKeLVpZv
gADhMUZZQGshlYeXOLTcb5NCoWxyF8g+nVzCB/xVO9y09xr2BgB7yty9zMSnE8JB
sabgSssek6ubto8uptG4i2OtXOONMzbNI49zbELP7MKcV3BrB0WDmbGWm00107Jk
heWa3yCCT+3j6dU8Z/+4N4V+Pxdosu+o9mD5IBUElOCaUlAtXoACmxs3M2aVoxoS
XWOiaiS2Gz+CVAad1oWr6JljfNtcaYKliNn3tdn2/AQFRD5EBU8mQ8kwdlIjVLkO
1PAt3UlCWIUXHNxtSF6ZEq3/zK/rGDBaZmgp0t2XeaukFJxbjF7oaDgZkKXpNwkL
LciFAUV+FdQFrq/qzbucsnwXVjXf+sVrAXbechLKFbSlkylhdWSzU9JepadaC0ax
XYrKx8g/6CjCQcoupIPQuieXAy8UVAFVkjC+1ThC6pNMCvCrGuqs28OWrrjnPzC4
kvSiczHngESrUDcqSWvEVEzS1d+wfZcsv7hpq8TEbIznuNoQVRRmmC0hrnnFouf6
Gb/NMzcxOVC2cdYR7zrBHKWuMFsUpLJ/QglOt0CXMv8NExWE3ITVn7o8s+5UHk4W
yqRxjsP25Q0HFPqOnVXzVgHk6w7heRhmawAwsLRN6XE38NAplu6MpPiqsCpCfYuz
TZU4Owufi7ompBcUZJTNmFf+SeWZygX+viRbXADZE+jw014d+8MW6zqtBz0p3mxc
Yg8+Ahdf0+3ECephKwsMWa9nKFFHQ7k1+U6+ObUJJh3X+2Unm3gCbHeBDjpvb+P/
Gvyh52UKSqMEmnCl17kZ4s8vZjyvYNJf4vfHKFUiRcSJ+mAu1Ti94cAz9XElF2be
RsGDOhPHt2PeXLQAJZgza3SkmRN86Xp+PWRe9IYH4v71KBo5f11qcVM7R+NPLwjV
pZVVMnCOtgr9XOsQLRruQIBAKL8d8P1flHAl8mxRCyqIK39PT26Bu2XneZ+6bwgh
tvZrPILQv4S1K3VWIjVZinHnIs8QyAF9vo5Aotyha8m3AbKX6fCaKrvYYivbblQS
sJXj8Crz6eO/rinr89ZKTkeAjtDMKw0g8da4B7Dh0XRtkKEwv5w/eVA2j6UMYUi4
WeDIQ/HWzPQMTdRc6/nhU3F0rc4m7Nq69ipcCCMPrOwnNxZQwtGJxllOfxczKmrm
6fhexeCig+S7KBcPmyuH5wKqIaTGOKCOwETARa1Z38GZzitxWo6SliLOp/WtxCWU
iR79gaxRGvXH294FA7UgWSKp4bjHXcwOffOH1gnhujKifJhPS1K2fQD/ZPk6s4Ho
M5r62QPIfKOVJGYq8vIMg8ozCtuB9Jw7I+MnFN/zeEuZXnPWxh5pPPUx9wNJ15Bm
aZW6RfobAuW8Nad7+EpUV4OhXFPMfa37YIDRBePRsuwkEK/vD9PGmZc3gcAa4nFt
tFnSqJuzEmtuZNidLBUid/arhWNHwHwREzJIvkx67uhRIU/M6REltBpfRvV2quLV
rpLFA4+0RgjB/9Q2aRHliSbpCO3Zi5ybZsltphvkugakNP1XJycYgsojw20rjGWh
+eGNsjYs4iWFEa1uv6umz5uIc9WiL/Bj89I3DtLK1aEb1Oq1j6ht8xE67YWz3nEO
S3kE73AQVYg4kvJQ4dTiSb4aEfLRg1thRB5EtVOMPapfnLfteOcCsKBd8dYFZc1M
u0Zm2gWanG4xn/uKBPYWYKsrvdoJ9KafjIF0S7l5W1eBhXxaavZaEsm+5wLqq3ED
1RVposi4fZOR5acqKES17gSrDYQFObVnaA2q772Fwh4IZZ4RGYWOdTV+a6UFWmlS
BFGbTkLpvVZ7i979g8RUAT6oMUspGelAXBjoeyXuBLxxTNi3KRBcPZ6gDV/NwEh7
HyjOjcijNdNlFEVM4wzfBkl0azajf7EulWsGpJD9BVTPwtSY1L0amISNv++RAqd/
B4tQgsEXXzwF94ydEbsBCdb8AGk1pL9ksHYipUJE+hLgSNPfZ1xHL4KHWig7yM5p
TUOSB8pEjWPsI//N2RyAKL1O15tWb3CaKnmMklqOwtMI8+lPYRjiQvCvleFumDx/
a/gIts/jzFlqWBSbelzvvlKr9ApH3JXQwdFdP7adsQv7afUQEDeWt8G4muyLXr5h
hho+TDgMDn3srM4sJmwCHbGLQcGhKFaeYPXIfsVMSWudub99/LEC7xY+tw3sfGD6
7t/gyVvRhwn+jAA3kDraZhjSqjJhNleata1AQyiBzMwxui47aGCf586EjOYmC+Ml
YYpTw5a3IV2VTSGhbm2+Tf9UgUg4b6fZbt0u+V7u28ifPcxoxZgf/n2ANkhX/xWC
MP0E488xyCDm/PgGZz1w6WvGF0bYpldR8jD155oT5TZ3O+Aln0Il2aIwQWgENzIX
wH9mbJseDiMcXTGY+gwlOZ4rcbizNofZ6zA2ifYmSm+ESI8hMEDQiyyVtoGEy8O9
ADz7naINNwecWr9VWn7HfQcAb20TBxSc+LAM470XVR/H8Gax3Louad9Zalg5lM6S
acRIATQ9NOs6/DqnFDvSYTq9zzzcg7mQazhFTCNdRJU1HwonMh0t+MD3hgToCnSy
tJwo+SyjC2lx9fXYTi0OvPczMjW0PIPUZN1HGRIKdCG83rIxwcBqCSPzLN0bhpuc
IPnSDRCnH/ZeaZOcFO+Q1KtrWN9Kfcy+jrE59mKZzvrtshh86utPj5wij56fKt3g
Ym9TnltjdxiARDOaYd8i13kjdP7lC2r9ZmOiKL9dJJYn/Ezz2MysiBBAMmnVR/Be
xUXTzkL1sMYs7dyQjpitIHLtbU6QK4FmhPauT/ZEesybGfoiqZ4t4gNZgq8Gr4/j
ErZK1gowlj1EqiQ/D0ONEN+fMDmQxc+5zf+b0BIUq7Umy0sGScE7CeTBnt7EgKcy
lNCXVg25Ouvnr8j3JP4YfE9iBn3Q3OsHipmcI/PVi0sKCwyBe8H2J4Smb8lHq0W2
k97RJEtd6NxrK8HQi5Dh2lySLVQO69SodDumLVEzT+43l90r2FugdVb2IrWncbew
AMSpZMtcVXeuILu9QnhOeuUA9/9ig22PSc63/sFcNPqwtZRVdsevWm0NJW+WBNFF
LQPISlTcE2R9pVmvqfFBukhVYbw3RC0GDK8deetMEUt+2dkF2PmT6/IqN7E2hrTE
gbSwlLgc7dXXuIsh+gumKuwWr/xsa7WsFuWK6N7xzzmNOxPyfLGpsx6A5rshgSLV
QwN6v5zTO7gHUEdHAjaAwi9K0GaObpOmjbP28hHMdt6Q+u/lRWk1ti9yq03HEzvE
Y9JDA+FXFrNfaFEJF8YaR78N0utLvxiJjB5EuKvI5UJ41I/6Fi924votU8MAyg4o
w53/PQ02d9wRFYtdLkR2JGlHiFpNbJ0mVAnlh9+zLHrDGlOOP9LaYAX8DGIYwIe1
DglG93Nm5iuibOJAf3VGq4Qv+8TWsCMqbMGBcKSo9zhITBpIOVxtJwRZLcEAmANg
c8mA5EEMr2iAOHBBaDK/z5Dgtvlocmw5mcuzhSl3f/F0h9n3gBop0eeseYHIcTPl
ocopjLF7EKoAah5Mi7ooaZ5LM4zzWNXh/OWh6qrKT3ciBcWVsbI5uj17Ko8tIid2
w4XgBpAns3WqgqjqIyg+kPb1EGw4L/HUzgt09koXSBC62Jpok3pOvX+xfEqkUM7O
GNZJ7ys0l4pQJXWT6dmxY1HDuilEFjvx4fIn46T8IGHUZi7AGEVoyjBmmyyCqzI2
uaFW+jvhXt9RdVpYEcDeHPDxuMuX+DwUTzRYH0Dou+ervglm2Y6Q6pRCvgpreYFU
y4eMiiiH+/IgyqnFfQjXfe1RkqFfIW2SNEIcVfFwGw5Cb+lrklCjvuuTi+jZqX2I
wSlsx5iCv34EhL9MvVBZROA0sarBTQD5mRyBdF7gt/EoO4JueS+UWIsi1VRn7KOr
7HbZIBNoxN1FxRP9C+0Keq1Vtk73nUm9YcNQcwj+CujX5R6+XwU2k7vJaPKSoGaY
Ou45kswelpHxGjggUsd1rVIjf2anquzal0S0nC5PJY0dhQ+oO8oPYHwOdXIgq3WV
BYhwLKBYMdHoKKh7vsLHCFJ9b4wW8cjDiVdvPLYbnSOiflvWe2vRlpdAHFXGAAtP
btn5TdJYmSPTnb3u3QLKArKUi0ikoW3srrFEW0sqjvBgHGDhAFX3dfEe4Deh85UQ
mG0iBB9jnZ8iBh3KW4vWpx7PL+YJSdUXDf8n0m8HEzMWvY1tUIEFkJYLYZhfSCQT
BovPC0tpAg6eU03Q8AwN8IiI1S00C2/4SIqfDjixla3rtH46rYUdJZiLy1aUFLiG
NxesOb5Cpzh1ujwff0V9TPEeb+nLem7/+iRYS1Klep+f6f3G3qHdwH88Bp6VispY
KRmYjnN3uo2AsedZFbGpDZgyAg+l5khyLE8pL07j5v2blWcIUQQnF1RfTRfXLmWy
zbo/N2JzPAa5nGODxiS+Wb62cIAIYHSoaJEDCI0Ff+dUKmO3X8bfCE1CPufMGwH/
7c1JDJ68O1C9veaveiRRagRk7sJObHzzHoYS6zDn70OWmbZdcQzLKJaMJYswVsMS
EDpWiBBwzd/p81aou8F1xQRjnYT1zbcfPose4UBh3nm9R9NJVbr/VpkFcX4tKTkn
fM1qiYs1zSWm+tCBho6neAzyPjhXysvi8y+MYxFogV5R45OY16Mzq32MQO9Fv6bq
h0dS793FCjNsl62x0YTGww78xkCsGPhPFCbwgJfQNEjunQRldgyKOLOOBXRJhIpN
RYnM0tjLysm6Dq7UOnr5RW1trBTfT0aPNvOTwQKS56R0mnqwaipkHdzvQ4Rz+J4t
PFK6Fe4VqeV64YEtEw6BRxad0NW/K5PvSr0pbMsoWR6p0vcn9DnZiETLY17NZlCS
Pf7TMgFLJSRTfHTBm38Xx8ogbQGx1igW1Uay6M9wLpv0iKbouXyBWCwGqyw0WFZt
b49Cw9Zaci69BkxCwzP2azS6w/Jkdl6bG1CEKOymsEgcZAhy+vYS68nfguw6hcFl
Vx/AvGs9jMMQIkAgIBvEL3Dbm+LIMciaPwGpoLtftlC4BH1D2CTkr2TK9VD+09tB
wtNHg9VNIDVjuvAr0emZNY5Ss5jC16sEWofyfMpwM/riVG+mA1hS2bVQdf+bjCE1
JsbHyZPwWwIpMEByA8wIzIDDCcAgwECZx90p1bQLXaN+gtpQlj2t74WTky3bIxeW
2kf2J9VmISCWOX0TD2ywEFVU9vlgeP7si96NGoQBXT0C+LKr7xXpiihkBle1GGDn
NqX96LCHEoRWW+AZqsJg3aVD2tvtgucmrjcusi80XmsM1mZgp/KoPpceVcUM14Vo
A6H/4uXVb/0z1eU1K51LVWpTFHoVRKchsp+oMFrCvanc7Tf2UO1X28+zPsihb7+m
Rw3XAfjQZSF2tSPqHWuezpXC4rhQ+/PzRf31NDyF8k67rdVphwro9OG39pMFem8t
lDBxmZiwUTY4B5E0a79B2fX7Qpds1kyPFm9suaopefp0WN8ulwjQ+tNWpjU4oJIf
BDATPk2MKfs+Jc4AARU7/qRTYasUYv28t0HqIKgZ1OxUV46hHLP1Og9oqizf31cv
d5yh3sRvWgZnERGuv3//RfFnZViKnEtalYXYO3jcEGjSCxl5T7aTaX8QEIauBp9H
02SJi1bUxYXLuWxMg4MJRMbMnimxxMmI/t2ZdDS2D3hO8QxEPXFTlLrljJ+dCrxF
FO/LDPo56A1XlcAEWPwKC7/gWDKX/5uC7ZChbroCgBgpONJxxjuees1LUB1w/RAo
nl2HccHjIEZTiZMqDozmKOaB8vrbh/4xIZY8swd5Slnf6kVEkZhO5VBeb2xcNiEf
i38pQodTbhnq0opOmHrsXDOEhqRM7F+Sgc58/lVf6H2KC0dW0oMadLoHOQ0/aY2K
31pOv8qitv9XgX22BXOKGjxI0XB62B+gCbzaJHV58bKPwxljKLEuB//Bu+PDQExU
gqqdjtJTVhXWru4JnNINF2vXSLp/IFXc8AeXF/M60KhFnfKwpMR3Is4Q/9BrYgKV
UbBHaR0o6ZkNl7ixUpS+1Z6WqH5nBa4AmJxcUgiuYeP+8IJZ6Pvp5UBn9bTGhKyq
BrX2PZ4NcAu/SJIoyFAmzWrzuV1IeLH6sjmvFfK3IrwXsNGX8dLuC4XKqbe6XO1Y
TuFYvRZcCR4fKc4RS6xjBFyD1PnTmpux6fjOciRDReJMtGUq5eFanfTrQPHzuhNl
sCb5Wx+AO0YJGFbofVyONF4CC05KLZ65+PWj9W+lTV8+/bhvjZc+geiOv3WzPUAJ
DtFxUANtwitWpOoAXwz6ylmB4qAVelZUOaN5fq4PZFSXBEF2o1TrA8CHSg2pMMlT
mQCeuILYF0FBHs9imuN4hM9UZ8lkp47PYtAmadZHinSwarH6pzuUG5c7GaPPujCr
A8Qpjta9AVxIkJxQVu7pAnSrjrUS+URpuEbeYxkfvwrDdFshoRitw8DP0kDXQQhI
VQxjv5teDy0qphSNAlyOHt5eKIS85tCwqP+G4Hb4lQlrnVHvyop0jDNyWMvBiT5E
os8wBwmMRIDZsqYh3RlP3DJkQmb9lGyK0YpFZW9ffriq41QNIbBAMwlXg+VGTUT/
V/+rlOF+b7cFedP0dWOfW0lWKdEa4eL/qf51f3yTgWdzZaUPW3Wfa4yO8cQ3lj/j
2nBQKX0zXCwOejKC+nqlth+Ftc0C7vcAU2CU9d+z/USwnQU6SAWEOZ9VsKhpBFjE
SnFCkYkVow7ioOviWQm2JdrEFCSIH2FquckrE8bMusFT5YJZjupIJdZohXkIAjac
ScIF5sSPBOYQR/Gv3w8f3drsj8IiSe5T6mZEjIV0BOgPiRwI3/WAYpL/pmsO3AEp
Lb/BHImhKeRUJU9z1Am04nDMYA7W6G5LKzb/0bsvhVLTiTGCwJzkFTHzi64FUa3B
bpbmDfKocuSG7z8him+5vV/ZcWZVs/oPpiIMHYAIZksCL+ZIJx2fHu/Ax+QGGf5i
syB00rq+EGNC2jp9eALOT9Oqy4DvgQNSESmLBtP81EWx7Fftu7VPr3uYQPZ9ushb
HhLBF9gmOSJtKt3bahD54GK7XurChrjq9ycUPIJM1fcxhyg6CRpxiWLZSssuS8v7
l0y9DtZLLSCVj61LyXQH37MJRQO2l4tPbIno/eQwFmDfEYX+heBHfL4E0dAnifbu
qeY1Y2yq/91pIfa39Bk/LKoZaW+FwIl7VgTLoibDdST8XXISbyo5iwthxCAH9Y4g
xFTzEhMQquQYo/iNZazG8pyONRBJ4zHEnnH4bSOj5aU/UlhdVEwAV6ncpcs706y3
PStNETYUOVK/lqYfimakAKnk++dKAeUpj2Jw7NXLhjzfFQpy7wsvUjCsEq1+imXi
Nb2pj6QdIir9f47Z6g6sXeJ3AxaC8euzJNzMQD1bR/A2Y15+gM8InM9Ff02AoNET
zGnwZVtBYfJ3fNVs4gGsdOl+d43Id4+wrQCrT5Jn+rD3ZuQRW5DD8azuk8MuFlDL
fpKXiwq0O//FwhDEEJpSEbHgrkUqoxtJoB8KP/pFLWLArBY7hFrQS8OwQRsUb09z
qCCEpQ+8R68//15spD0xzOyZr/W/FzjdxRIa6CwFNMGT/zLGx34dwBLcR4YJEnbv
lFmN5+hIVTDVL9U14L0FZ5cj/rSKZl/jNvtt1ZsjU6BHnv2i4R6j8qpjbaZ8OhK3
I7if1nNeBvJhdoY8R9sUYzVMU3kSQgAzcpz1HO2eR4HkKja07KgGRz/dDrQgBsJ/
r+E62NDjM8Fh9KysiHg7bjNF5+1BenYUDl+m9JJ7o1772MgKAec6r/ldY342gDdp
m5bu/9m6GeUlIHRWmArtmhp4bigX3x2E7gCANb9i1dG5M1dTylJkq6TZqu4out+d
hNC4RzYyiupJLIYfEaK7GpxYCTY2iczUUQAqjZTQl1WHvlZlwv9TptzuoyJDl98V
FzJSj3343qSnHmOBFq4R5RBqD385TMCkQXQd5i4yhD8IcK2Jt4qXNsrChLiU7fAs
InTejRpXP2ZxGNCQPMIuvUm/2+wKe4N16POuh0LTlqRJsjFkQha4kFN3qgdCI+Wy
OAKQBYohGzhw5Es86ujNGETupd4CrfORTM1O41JB1Hpd6IC/veuiBgllBtyL5FCV
rm5SYXTHdERLMF/ocP/DvKMkNj1BL7pRr2Odg2SO1B5wu8XqPxYdGamFMn4eRHa5
q60g6so7TnpGbclp+X+ymbf7ammD0tKmT1+CjfaJ0R/2n2LCA6iirCO13lCsVLJJ
ZAMo6ug16TynuWdM3aaKGQYxr/fN+fyvsKVPjAjnHdCl4ANXP0vGrKdbmD46Zcbq
ndCZSST30l274yn/Xs6yt+K9efWcmVZ0d6TS8Su8t5bLEFNZ4Va7AhgTNDZQwthB
xbT+Dow6/Kz/CKjaq/bkgK/XlMKOvHhcns73Quh1bRpmZUsTBveM4Bpw05Kjz1XY
UM4N1fQhK5JaAudTcKx6bxIfk5p8uFWZk3xYmo8StkMeX60Gs5A65BKpcqc5N8Gw
3g1oEwFlA0WMxTj9vPCTrVnQVUPtVodakLD3gA8bXdTRLfZMKTlY54rOO34xAqb8
BmmtWU8rDx/ru7ylcFt3Qp9rRZzcd13FHiFPizwbU/+Dnavg/a2yaZjRvAmJa2Sl
Zw44mxAj7hCuvg2MrNrBe85dzJRixo2MGlEjoTgog3IbPQDsAqhezbEHsSRhV3OD
HjvXy8s9TUh+IeLUjHONvmOuhQRLSbO4b12kjJvv9MLIn6DpkK5O9NTYZ6aDnvde
mjbQcUW0lK0l2MUonURwbT5zw+f33wX6NnefKYrbmycNAY1i85RbQmV3SUGFz7Wf
w+TM+mLylUww9mrSSAk82Pp5rmijfBOraP5oC9sAs0akg6uU3vx/3N31GtqxQwFv
EuE5XHxN40K1EeTn2h5cogCzPjQL7TSwmcnepRQOJjJqwrF2Gh8fuUTR/cbfBAsk
t60zwWOGgPjGVSMCSmfyy1iZSipfm0YFl1CU7UtiSZsaGOoev+Hm6xeIsspt1jJ6
M8S7NIUf5Q7zMP4fUTtH8ncPT0z+Yb1OZ6CJqUxwJATBmVIl5KYmIsE2VZpN1erD
oPyPx79C2gsBnZbFT0xIy4Wbm+ZHersjmJw3vHBdSFZjxDrj6XLdQNeKMJF4r/2B
pkhvvbYTWJgbknhUy5ZSSiTwQKR5bzlJPbL51vMEawEGEuWryOYNWzyuvRQfYrHK
PhrZZaiXpf86eJy1rQtO7s+WZu9svIYgbRach1lHvGi8HoSIjl2qwjfS8hjuhoKw
sVQBBoWcDCCcOezsIRuW6+Wh8xZBbDmtwiFrYnoguV6ZOWoxcex402CreE3pH0cB
/1UCQffpVbpilDUllw+ohizJl3W99jhkud7WXF3b9Vf91F98HMB+u1N21rFoG30E
OK/zDi+aJCDjzUdpsExVhKEB8t7+Rk9Zg8jxUmwdPQIVI2m0maMOsNWbf9s/lJdX
v9h5RMfUs9bKqpn/yG6OMc+5bYgYe5/DwT09YGrrClhHYql0++hRl9t+JN+I7TpG
bGbRB+DCdCf5XNNqGH7wuLMN9ziZ0DAvM4e++006cns+L4N30cOSsVHfqg9XykqZ
4fSmmV6afd4f/WXHoo1hl51hQt6S2aUUOf3mv+Phe8JASvRIWmdSNnbzq79G9nNv
rRZpg5CjkaLNPmaSs9bvy3wpGY32411kTMSyRAtyl836kUQI92DRjzQWbozJMydZ
/1+1rk0IHzRoopKuEnR4PWHYOrIy91rzc3j7DYa4ddjYOj3fY+i9Z+4BTYoVsNmB
3bQ2ec+Ov4se6PmfaikIbT8PuuHNMP7Y75fJNFAHnNOj3rR7CecGzgVlDphtX1sz
p9nzFJJnffqJGtZMY0Ux7YW/r+SrNSz2+krHfv+UPyxFTtglJtrjq06dDKEPp6um
LJfO54LtQ/TVJNgieRuPEW45LQjs6au7abpCvMXESQbBwpNi+pZj3eBtcfvedhuL
0DBiJA0GMC25mRwzwxYr89ykmOx1LjjxscpcwMcu2okbroRVH9UDk0LQN5c6XBZi
4+0YYkAG3xtHb64+FHc99LYMvxWpKoHztWBpJ1BNHUTGq1T/JF2MgUi4lMegmbXJ
Hu6IT+KmB2jyhYBxaDIWldvsIjqV3PBC+BQ85dTtazCCG8whUwsOxrdUGkgJ34yu
OlZfel+f1OrRS1s1OSZtF9IdYAYwswwBERgvtm2CRUPLWvtqeu6ixlgu5HpUZqt0
tNIPMXhKeJs8TcA59nGVxYmsECLj1qKQYyOCs8VqDeiG/KUng7W1T9ZeMx2Q3P7W
m3ZFw7YHDpkAnivKdXhl0Tv7XGJNUwjCMa69ADZHGpHH/jtgUqjq1cXyU6qlSTL7
FxqnONclwqmYmZT3HFnHl8yF4NDm+VROG1bRY8N3mF6qt13V/c0Ej4oGC+bZVXxr
CbHM5noKqHSf8+K1roHloKX4DAGOGCnoksWaVldA0+vxU6SayTlzgH8Z2MPbZvW2
1QXD/tqdODsLC7+dqy4ZNkolMX+VkqRXv6AQdRC8/hCkDE2BouKFIwSex7eWRMA4
9YsgxtVhYAH6o3bNhEaL4UBvw/HopVgIQrYjZQ+oNfGy/oEbc8+C0iv3/wftytTf
AJlFGsCJrUhT292uMyB+hCcG6xwXS13oBOQHUBbjtLcMxXuE4uVtWXFGGaVfKUwj
7LL+RSHTzktR9JaQ1Jfv5X4SC4DksdWu4gMculxU1C2NwxlLJZrcZiyqlBjapx/Z
dABemOBR/4MAp0z6exH2EWeGzzhOlv5LYdDEnlVpZic5Xv8lMfkguMdM0CyQjs9/
IGW+SQDNTY/fuCOJNVRGFEd9Xz02C+9t5R3TB70wk/uAue8ElnZyfdZCF1fkHRzX
jpJcf/tWOYtHJWeC4PRC3a1I3JGMpMApuGzN+jr0Klt6HiAvRjsEiAgF6IHAzL34
FCs8N9esIZme7WyRelVqA7OdyIEn4okfBWzEfy7DMZK+Y8EAzek55YfYn5HPaFLr
gIXJvu1TeCwSyQse5mldKNAhUdRLwRQ1+Lt0+/GxhGmAZl16QfS60Egz+1Tpk5vJ
7sw2EmkhZ1GWtxTBMf4GlKfoC/G4tE4LN0TQttlsqjoRXLiHswJ2Aayuu//8l/qB
pzyMAs1l0869GgS2p8j7jgCXN9eddxW6E5Kk0jR42XyTxJmtL+iXy5XG/ss+oDtX
O5Fw5nwpHFjjIBA1tJEZ2cbJpioxgRpE3yEUUqL4/2j+JAylfysx5vtSZ3IpHgU9
zLssIkXpCd6PUi04Sg98jPRZPBZiC0LR23iFY/WK0I4MdYa0vBJryQak8fHtVc4V
C8Q9FgCZPZyicgijOd8Z9BDW+CJTtlxN2dKaYvDLk0mfHD8THYMPDUf1j5nHPaBZ
a+I8SrYWG+ReHBAbO4TszGg3f8svHBKs7sM8ZFwb1M8K5RWd2VdWFx5iJyCAbHUL
tdWnhHKbcJD+/Q6h486md5+7ApuvSTAAfiQBtvnVfScw/Ug7F5i4BkIBp6SBAJ7U
mGn2SQP6ygxpyHGdnC6VlaijI6p9fAQ5XN12HEIqTjAVvNs6Y/x1QXGVHnWcBML5
3f22xyggjtdh9F3nAzl9GvxFifoOkqIjhNLWONPlH+g76H+lYEep8jBWJb2nzjb/
R/LD2CCrO+vlxsuUralhzcjMLGqVPzmAyDwkvyGwk/0qWAXxyAfsIkHfNp00w2DK
geSkzPpk2JhMEvj38n6jqSU2xIOIsP9b6nu743ECylWsIDEAD9yOVs4rCVsmc/Ju
s2kpo1EoO1Xyl0xbyJNmsH/Hxl7BbJtayIf3OWjwShjCDpL96BoxShqHASBSIxXn
cMhSZiCq5wLNB3a5bi57BfsUL3YFYGrxjMn2Xbi0d+9EeTYxK5hoNZpQU2oVI/3/
jZq/mDS0klD/VqXfHb0kVeUa/8Q4INxAMUTMK4mGj3ws28pSKRhKQ7ZtxQlVtDso
e2fKC37HwShoReBRGJ2t/6z/HF7t0MqtEX1CbwIXcFa5KYx2s3F/JW1OWvtrq3cl
9mQzyJ/HpT7rRXAOxASIxxzB0PJkPMDCV8bmY2b9R31HqnWCBaUNDiYbEkSdg+4e
wL/HzQlZumRfaT3UnvS20/1itXpA9O+Xwm8FdFRHGddEdx3LS9/r5q2oxCmq4juq
7JvJEtyrTe6Ifala6fQx2gOU1j1UCC7YxeHvuIOvBs9q58XEzvcv42y3KuTXLifd
QwBr8KVL2j2wjcNFI50s2U5Kcgc3Aa34sLd+IIJ98k9YX9yiz9mNKw/up9/HPKQ4
N8cnOIuqq1ThmO4szE70QmSiikueG4U+wCdA3JJ1QfHaM1Hqm5ZtJSXCQkvtpvt2
plPiXkM+1+i84VmBo/QclQOM1W273a708BKqzkrgEZzZmBYTNG9qqwDLOoBBNhK6
pi9nnUjfk3UYA9Mb8MDDLq84RJEzk0m3bG0CBsOGuHWs3dPSM1EEsqDea1U6BzBy
NH87wbL6yGk0fYiPVHWY3D9rDDc/sysen2ccfPQBzuN4bnKV3WrQZKbbgIxcvhNw
0y4Sdob8FmzfQVAuA+W66OPiIk/vExR7o5XvUfzbjXYVf1zXzRRw/FEvNoeWE+50
dtCAyUAtPQsoW2b/qmdXeunMtmVHdCHzIwV22T+uatNTjHEkzu4DkxPJ1avE4vHE
5Ltr62nJ4tYYLt0Fl8IPq8NTu0CiCQ1vK/6upwCmImBCRUdSbiHA6pER9VlloOpo
luL0uq6IfdQrxjOHBmUJNAH9Hzd71TML4S93o86jP5cODDMAhl4OVdpfFotejVmt
kH8Ab6+DqdYV9DDz56HSryxrJmrIBjZYhDqAyFCCZ+hj0lrU/TlXOTKFCmk89gFU
iFvUEhr+ZyeOv6S0C+z5+z6ReTWMTn27Gs+pQ7gJJRUxdU2zel4XZkTvTVVQPC5A
Uvlxn+GvJEvSdRAYnkHBuYx4NgvFg7Q9VYxBkd5AYv3MW3bdAPzngnFHUDRA2DtX
tFabA4yL+z/XppNO1vfndg/Ai1TLyixyXwJwA77QTwG6zZhsKMW6GAhHoslKLKuV
JR+2cew9QZibLvfpbYluP3mkpvRP9rM0pLen1LHFJDZVa3yEG7QWUCmieIY5LnZc
cC6tOH5+Zrw5qNgl0A3UzchG2F2wlDxbx9S0jv4JE9SJk13KceGImso2TtpORD8J
Ua6v8+wOFP/gfPWX6UcZZmRhjzvH+9ksVN6s4uUelxxR8jQARs3HHKdzfc3Rhsdq
Vs3Pr355hAKEq73VoPvXFF5VbSxx3QK+cjK+V/R8KUwgtJ7l6IB7iEMc/4BRLCZ9
Bc/MnOc6TEpu6LKzxZ8X7cicl1hMIWvHZ71VpO+VmwcyI6O3LrqhV+BayuRsgy7r
9B4H5fUgAOoXVqjqgdplAyJL0TgP1qEx8BYnB+eS0WPYFl9mFyRQqnF5kWy8pMRN
omTrVwfz2dpSL7aI6iEWtotMNc8cGBTAJp1dxEBwck9u0OBdhl4ZrOUztOLNDvo9
8w9sP4+m8eoGu4ttTAd+DoqzLoq7n1MBN+10OvLQBu98u0wc5f/eUjduSxDsHe7S
m8cJ6XJATtaI6BL8o2vHC+u1+eZr/ub06dbQH12fhhMuMCPrYORdKC9/511YtpXE
ag9JninYAqQ+fkvJuHcpzjUFjdWKM1macPkzVfFC50Ds6yOD6M9daQeZrbHaRBmC
BrzfIknJKqqLQkbobwsv9f5qKbB8IAAnoYnd7DD19AiH5EGxEHktPuSODe/bj9HM
e8x+rfeyqcX8jJZJm8PkuEGNS/KiwM0tJxTwJ7LRgr2nP5BF4Y1TdbPOSFe5Ubzr
t0d14RP+0N/S22lwWJFWLdOOoelzcP3MRqmCk9CMh22puLT74yHfkPOPZ7U0bFjz
zIOsc8+DzmgtEyGcs4IzYppSisLN6/bR3Vhcz9HWQMXV/m4WuJU4oYnOarJUd+uZ
BWz5a0P3SI5mr+ENP8Ook78LLAwPjrxhdU2uuW7249W6qGVDddf+RVOGUTqz+asG
jHJzNENIseYoKse6UhHjMWvyzba+DjvDzdHfR05lqlZFd8H33ALyDRb8c0xEeuFC
xOvUrr4UgpqJEXElnW7PvOX4VdEZa5NSipC2jpHsbjqiOhi6k4L39paeddcmcW5f
AwULap92mb6K5N9EDdo8q2ZMQtXwFr8nKJL8jH6nLqljUyqNQ1C8cyxRd7bTyUi3
85J5MWipzwkTj+DVczFq8KNunjEDJgDjpNWdXtv7BqlEpPXc7HLFx1QYk6vGyrmT
KMcrGSbXn3ZEu3UGM76pdNjD+mcNHij+t7GVCLqT0RfDaLMIop0EthLv3vuZatC6
PlRbwkO4Fj7GnMwh5skSQuWwkX0Wrxo2Nat7yLoovbmn7bJNOaL/c3VdHECuUXB2
0+v/HM1S6FwemENkK52V8ptJAcTkFy2NY/rbI6NzSX8ME9wpAqFhgItResy5giar
YHrAWDSL6L8PPH5QL5MOhN2lE7vKmiMXx/dCKlBoOPlyfn+MIU/ern+3Vx3OECQ5
xm2vBTkiEeBiFIfaWDB5GbAJcY1UZerviTVDOlYx9uXi2g0zxcH2i3lBmh89ecu9
GiDA5RfMUmXUMzX1zd1ELT27vDdx5o8SV2E5Z92QMvTNXFBAy9RgeQXPAXOtiMBZ
ew+KPhut0iPRO3YLTvQQklTfELtEuRsxmBj70+Tg5pOoie3jy17WbcTNP/V/rGp0
7EyuwO/4I+HzNTjwm+++rsxDka/onxD7dOivvgrTAFk0lAebfNeuLb8rlhWQruwC
OjVW6c8GE53Zpuma3bXj1ZG6hQb/thUyOAKHXMaPxkwQKe0a9V+vBEg6O7P/Tbtf
iS1FG2VaPnYotCOchzw/w0mGhKRW7JuypQ97XT0hk2SmyKrOdl6J3ebTZE75rNVW
xCC4Qoxk84EGcpaFhNAXiXP8qMpj9/E0cS3NfrzcDkYeYZCwmw0XCvg1dmFnEonB
R173ZqhbJvjrgTRwZtDSU9fBBvFrlJLYt56UxaDk1dyym6pypeN1JE4oxIJ2m0CR
GXFVi+EGUtvfD+fE6PRjvXQz6RAEea1v0khtQbBr5z4lP5teggFJHWtloxcso+md
u5cplKp9MdhFkp7DWi+g2ciuN5VSxO6qa7rzNl1nKHPezLzO0MO5JNpcF2pyRsSY
EKNjkRlDBj2OnuEFGF0eumMFYuIVKEfpQGHDDAvkOfddY7ezk/GR/NTOQYpYAF54
3p6KRDJvMbFLFRUpyDlHReAily89dCa68RRRGHCjpu8B99rF2ybTQeQx32+62oAC
Tr71RqLV4YMMeEh3b5y854TM/Mi0q9fV07EPMwhdtYEu2jqiSuXO5ogim2MsOBoF
XjGzKZrJglD6Q+q7K2GinZR83bN7uQyPqIvjIUV0o4LZGG6iNxY+ciuYLxzy8Vum
ffH6JhkbQ8LTNB8v4lAvENG8+bMyg3fr28YqqJgE1YIuQz79mPUZ16ezDzDqznGB
gxPd0y4itAWYUcYfs3iNIMJ9xtFPCR8zFvwTKWIRBhGmsoCAQVpSHZYBdftlU1Sv
O8fruqAhwMVqViWcfEVhJP/asMRS2fMQsC1G7EE64JJr2PwtW3bjIXtLJH+v0bXC
D15d+5P80qLiV9eYT3MiZoNXGtE+D5boJyG52ceuSCEk1yW8IVdkJifVsNTAv9r8
DXAn6uFen2KmddK7i5tF67DGKnPK1MNzPmSL2z1ttb8OUz11qTyFdyz62r39TlQy
QE7etwdvbfkLwYASqH3xT1ueZfmttC5HdqdKFr3HA3hW2rGHr1Y2LTocWoPrmq7s
pVW90NuBU5lWIrK/6lHumiDkRgPuG0M3HwhfSzQvGK4TEgXNE6iZCPe574gGvfKG
1ScRu/dnPWTeJydbyottfYab6niv7/5tgkTfpLEV3a7fa8y1iGVAkBEgIWY5chUg
R01fHzSurEIeH10pV5APJ7fZZL+9vc+pmkvLnUQ5RBCYa7R8KTwrNANVy3Eejztn
0IXAcBpfdiXzn60o/tk5NgSBG3WnCyw0UGZELrjs2rDqZO7MjQS1qEMi1EWJ/w6r
lr81L6icjm+iB46D3fiKTpQ9MTswg1vaDPdPjH4ro9xAK22+Mu2Z0osuah/sEwx3
HnNKazk6rBP4FUGLG92J9n0ux5PDUVxqPdhYihcyfJGAEemgnJyHnK6kvH4Cp3+D
4YoKPyxtVuSDGwVifAu/g7hN0NJyeX5bgrhRKvQBIikSO4z1QZCUJztK7Q64qs2n
P3MBUStfoSE7p4xZ+llxxEfc6lSoNvbSQLUSu6vLWnAGMRVZCfnebG8jF0b8afe2
z69Oa7/ohtOqMD2qRpp+7RZVfRoPhyxuRLARwz7i/XpWkmTvvHiGfvbvYtOU4dET
E8XfWX3ECjPB6Nja5B+iZ4t4aJ2nN1U6xMY5T7l1+hqHF49dHyqeck3HsUuwQViM
7rXE2wpK1FPUobpqwD4A+DbKmedO9qVcktL9gW868zhTxSdaaMCRniA2UQejEdI3
pT9Eig0f2A+F+pg43gOwv73MHn0RKgHGVx0zyHJzwLNVC+DXHmLesWiFBy1hWyfA
XZ6yM69f3ymeJhUlzkTiMGj4l9NtcR2xXPllkpHXCbQ/YQM/G1UK82qpsowc5HkG
9x4NmaM/WiNLqBJ5yLq1qznyCPiqkoI2hdKZiM7myo4UCpjk7JiCiloKxkfJDRfK
YjkkcNPZL6xX1QeekAYKpEtH2gfszrioCVPmNMfKZiw9w8a9nNvox19iUjPpNtkJ
B0183PeEQAXp07PjWogBaYP5DIdFKFnJcXxldwiGTnrgqxp4QXiYgs7u1NYxH9z+
gLvAwT8U17hfqO0Ct9cxkRRWcnQ6jfwRK/z4mQtrrA9cOZhxWk2P/wJ8jrAPWpk6
+zcBtYbaDJoyy9TKHb3+ih6n0/ygLdnxsqPiOls3XRQPVirXsamgrWwKCKrl4KIJ
JnYofXm+AEKOcNGxs+bXepaBai91vMipc5kHEtDOHajxeCSwt+pppGbIU+CdDfR/
cdKyP18lraEYNCpo/Ai8m2A3OYv2ylKzuTzuBAeLkUO+E+6Ij/cKnVog2U9eXXmy
BQQw63L2CYwV8h3Fq5q8No53KTJqo33DaJKirBgw+5YwuqgQicM9/MsLTcjxcbky
+8EAfED369Ui7qZOSt9R/353ym1iMp53D1L9907a5Iztg/gVZhX2tnB/7kasiRO1
LrMtRbIDzTtPRrFbzgdnadcEZt8K/1ahmx1Ma4Fggf/hTUGkbJRKB5S5i0ffFlOw
ftHyCzsUnj71AD8xwZzA6wLjnXPu40Fu5zvuMXiEzv8RiffsQ6a0z8wIkqmuiYnr
wR0VsBDAU4kwLNbhGL3YkuR/NBZxOHhZg0TQFlr6p6tA2xnYLww0DQd7W4FSIbd0
js9stt/cAjVROz7JmJ2zuAiMfI2iKFZUaVeDV5oXg94XjNlylDvnN9ScRL0U/3ux
SwXaqT7fIxOUdGoIcHlsPRCTQ8unSj6wrBs4CaItGGcpo/+j67X5pfXmiQyBlkTD
3Y/FIAEVQkSsaeBuEyaIYscPLMxeZ0IuT6HVqnIfkdDr/rLO3Us5WZnkaN4XzxNa
QXt1kTILgVg0AwseChUlJ5hSToJLoUPFWIO3HvEM9wzRUWcvGPE1xjaEyehh0qFN
koa5OyXinpcV6iKwoO9n8YrgB7In+ZiRvLDMTmXMNRH7E/1UkGeCRTFd76a6Dsq7
FsAq7YyATlnfxyhxMfcA/YipgY9f/JG7e0tFNikFZ4JwJNF/pWeUl/WmOR2yN/Ug
r67yb2mdWTY+Tcqi0PulnGgYpxK48XUpWuLNKhO+rHSgWXZNWk1fJvNMi1mu10dL
EGci5TVwuFMwOi+MIVg01inoqvUsUtP5omxvLRHRNwNJRYda+frYSW89uDfBQt3o
0HkeCJESxuD8uPxe+lPzMgj9b2W3/c3ob1VoOnhyikYgY7p3D+pRfaCONZ7NMXms
cNXVuIX2KFyPmyZQ0q34MgLzzGUL6Ns+k5EcKRIdAztgROsr3wXSjElt+8GvfRfU
JkyeTYtsW3+8McY9WnwTQI7vHqTbqafYCGdp2LYOv7cpl3UfIRok5+bTa4Z4sgHO
rCnH8sUQnFFsNgB8jekIfe+b/KS2lc2rjm9SVMBsm6hs5gtwRYmQlLkxT3AoqUij
PV1/RhBt9xT4+V4N/z6ePr3phKfrAArhwe71HDWOjGCoJzUsSvqGc9sAPm0hfqCh
igTVTFP6LX3UDJ4H/IZj6ccjXQzj4wKHGPaqeF+sN/j6wwIL8EqvzE97OAlU/M8Z
N7ywjdfLBSLbUbwUsm8nUPxQLcD6Q+0uvae26357AHyR6S1V9IoqQnCBbMHRJEvn
J/ScvWe8H6gMI3QD0hZU8o6jv/3lY+OtBkjmvudY18+YH3NLLu+3aqyfmlVliMa4
tCgIMOSUJwntJ7mIHmfksri0J/ofawd/bHU+o0eMo1W4IHvmMv/tWWBtgqW7akbi
AA2x6UphymPFfNQBCSXjuXcibkVfjhHDOY4c9Qa8c9L34CLaij0sF+nG5uXMaDQO
S/SuDkNOcuI/flmDhc7WK6uwiP65K5R7n6D9KNgRVKd6+wgUiZ2qjhep0lH2ZRI0
F7Z2NwkCnLC+Ef3FyTpnT3eRJbI8qSlw8/X8Lq0fpQYR2PNUaqlVJTvWrhKMBOdF
SNb2+75jRZwM5MwJE5e7aEwLtOhKhPMwqE858E2kLmICk8sWCG+RHEVr6NKABGpD
4Bx70BfFX0E4yH6JbnvHcs0qfIbrdRoCtvF9bPj7OmGMbzet5ZEPDwTy6gLfB5x/
kWy17xt+dUjU4Go+Qr+PM+pUmbiBGcLYL4DNKzQS6KfGXHN0j2+LxsCm+x+aOp/i
ogy2qMvYOoGXhEGAvdqpP7azxwohqn0J6+0UNFEyAa3D2mCwSEx9mHspKb82GHSn
cEzNuj4n/sLzZTzJKxrWs6pEpuJ6LFoOsZiy0FevxL8NbWTXZw3Sroi5wYZm9Eet
PKJW/3252gdfvoVXWZF8fQTIRgVAN13cE8emCvys17x/7BB6JQLEpgOKVVabMrcb
vYE0NLCjA9khbwh3qETR7xS5SLZ3JS8lUogoVz3j3V/EAZSkglDvRyf8320zH4vo
iXo7EiS/t0TMO1HTHVbjSojy1w4mnysSJobI8idfT2XcS7zSjgbKp0vQxQ37qaX3
f/P8pWbJ8NVzzjmsquO3h21bKQdi0QKWjpXfXriwuC4LPUBvGWq2beGEQUuTzOch
RjEC0ci25oC5zcKyagXQF1zrfXnPylpKzJcHfHvnbzObAeCc8nQ3rR1UVPQuU3lF
+VWPT62eTdc0GxlkdYaGzr089v8XdFCHv6VPAiqLfoOztLovlidILNRj8MBFPhcs
aecDEfZrfALa7bxLXAc0XjGnSDnHjPbYrDoY6aaDShAVcg3qmprlOEfRgsmNa1uc
FhCXxxHQRPRj6eO9tC3yrmUqZIEJzrznAodyJa2OGCJqXFNd8Jh4YUyraqko93DQ
mqFPLpgNgFudP6FaDF3rggd2c833bjcoTC90JH5TpKuMseqP5yyEap2Xei8ggC2o
6QgBVpBwHNTrUbN7q74+bPr9LMcHbpn8gx+aqjlYqllckrQyb3jSonkrSDnMQvZL
bArLnkZ6h94CrLoq7BCpuVu5K2fXHDC7nCbXKoOLVIVQKDTpmPzYUzjShgKAuuvq
rQAwyEGB1fAD2wEYonwNQfHiqEqHq/eHNud4TuzJlY1xdvN1bC2xF3t/KOz/DFPE
CIafhTKHAl2K+R8XXGw+vgaA69p50xyVfrBFHdBqEkTRm6m2DlEmq1yOpuGx17u0
mQZyCrsAhl+TqRdoPGTenU873rrOxHqqtH8QQnxYHjrvZIKPcR/A61XUIEmVb/ZN
Jup2tXvfEcTw9p/mnosy28hB8RDU0+xNkErKAIv/1SWrU1ScQVv3il3jKYrbBOXt
wSQ9qp8uzhrypdnVa+4b2g+mpGwBz9ogHdgMpYH/UEUhFyuIb8WDgXsUGk5HL4ZH
6+pvU7W2l+06qgGKhhxyfITWWHRllj0sW2kJCgEQ7nq+WRnVsmRG2t3fYQqOkJx9
CdLQR0cXOXIFWLF31NJbfrSfZsciZyYf6MFElSG4o8ul2wMDyIWHI5pWe+JhxspJ
IDq16L47GwYZOctwYy5QCk5Yv7pi3emKbsEM4m5PVCeZzigWIISqzkp1BmL/voR2
XcTmnRPU7DkTfWGYrf/5ZuE7JTggr8ocSKohNJ3IO2FAPLcee6pYiPDLXVewlwf9
dJxNc2aHb0cZkLT7PfCFO8Z/5Qn3c0PvqzWAojHHCJcoMsbBceI7FC4XzRyxOR25
z4i7KFlQ2E9f1ddtJpnWzqTfqUV0TK3rVyQ26ZS4OeKm2ufmYgsxPNM6AJFUO4gj
+EFY6EVLTnCwWfUKcED4TG3BgEaTFyx5ZyohKohz3C6w5Mc7BG8X0pYPN8F487VG
tohhvHEb+AfVHzIYDL2JqdYDUlwpVdZdsBEMIolSWmPidBSPhGOQ/GVHFEYaeyZe
Zb7PNHzRxb44J6akK7MWsqQtdZHnisJ86YEQ/krHKzggrK2izR+uU02f2dU6uYIi
XwfEJ2qIyz1fVdzpGLRVu45CUQpOK1gEOCXHydRzakCzmhsAGX+zq/pX5JGI5DDb
HSvwc8byX1QOlK7Xhhe6XbSXSawqLfYCcoTB9VA5Lk4by7jT8zmRz+KtUBgMzqN+
yFQ7zuXsHmuCOWMrmAWWdgW7M3uAATLqnwiiscC8bS8S9BJp7LJSogkaTXsfN0+v
uhvMCKSXyM8o5nAUDUUru/CNDyV0rTsb43Yoe1raAUchIvf9qsI2/KlkzeSjZjdT
FWlbFrKN0SqQNoumzSfcPywDPX6kLaCub2qrEQmMaY1mbdgnGCZweBlAyKfz2XoJ
nHTnvUh2fccnI05ODCjTE9SxLPS5CuqPWA8pZ/UyIlad6pLxerII8/EcymSovqAG
kyFvVRJFeiLQwSj9xrPA18YZe1dqRGNw12L4ZW9a+rNnPUF9ofApMmOGIwRUrvJF
ZyJJLT1cbo+ezTjmBGiRla4u6Co9+S6HKY0szIDQFIcw6nPyYvR5aabBDRTJTH+t
DtihSa0S4hsTG4Um8QK+isRFMS8RUWbmvlxVtXNIi5Cxtl9gBNoKP1/n7qddVUJs
ChKXfEPTaCd1dQ/XoCiht1jmbWQeP5cNiPCv97DpzL6Y6E3GHs6KW1kKFwSntaMk
G4YRVE0NXkN4BqR98frPVhcLXYwIFmtFKvBRxQxADpG+Cpp7kYOPmQFnb5t2FtNF
GgPMfrp2b6tQCgks36j3yIPNd4EWb7ocWtDQTwsea8LiUgyvjN6MFZ1q8cOjk2ue
EjT4tH21MP2B9EZVqi001hWTHcCBbXd4kvJ4G9uA5WO53q80wf6/FfVvEbIqnQOC
PW7k8ZJekUOEPTvXYwdj7HHRoC3qv5pfgW1bx+h9ZP7xkH9/IDR4XCR2+MVyhxcL
1I2mTy6ixHMzcIPuJhky6OOW+wTtE4cf6sXn3t0IUF40aQT+T3GT7YamlPi6kXOU
SqQMZJI9c7hYdsGP5bDnAcHPmMsZzZ/pKi94f/EXDjc3eFrN+uUe5SWTKFPo1OaE
x7bVkhVRv2Rv6MWGOUUiHLb3a6uO/6tVem3Gxm+9Swv1Odu23IOdzVwqQspnItJp
KbolT9LbSgRf/Ys/xUuFQJDULO557BQDwg5dUDUYGLP4pZZx15ywKQVawt0HJblG
hYzmnhAlXDE2WPSpg371id2iOBf0Q1Qht6Ey8BSy38bU6pc2ENwV4MqB1mGcFiL7
crmVPlYyZKgqI07mhkiywEb0tqB+v1gPn822ZxHrlbmhEB0FYRIjxVyRo63aT/H0
6njMkC72RNFOzhoyD1IudyzD3mM3y94iLtbqtWOJuxAFVmEjyoNr1uDyjRLgGao0
co+WsWEBYQVoPVLKHeaPH7SW9DPZLppgG4XHY3UgejzT6o6dy1FMMrzCm4o25eM0
WbLJKjHKULeMYP2+agSufwTyVcKYvE6bNi1QfGnf14Kttm1L3PkWy78Rk8E+HLt3
5FnQejhWfcmoNSo45fr4Ybyj1UQPi4DxvxHBm93155oUA/Kp76QN/cSyczma1x40
zqblypz+rudbLVtynDEe2+WgpwAoidhw1uO+ejgEqxgs4NDKt0jKyQGi+TkqRrn2
AVFpig/sJQwQivL1ZKc6simTUGppHzsdRgSxECChVU5T45Vq+Tt0Ek0c3MQkkpyI
fUETFTEArCB8AV5b1q+OaJgkPAb4lPaZHwIq4VoJXnolTsl7XJHMvA5MwcHXz8YE
XAiNpAEJjjPScxv4fyuCxU0XTPOj+2eolblK3WrXwNOszpNxAafc7LCDfoBvrVMC
BrqWyoPLBoCyt1dLyoNLO23JnuxrxfRPE4bpKyvY9Z6a+B+YZLv3+i0c/x/IRvfo
OTj/jJ86tMgpUfpO9PVzmulaP47MlOTEUHFUdv1ys71WoIBCe4UjvsX8pq6dJUka
qN/jbITEUBDDqiXrcEHYjK86NBvkuMaf72RZTf5RMjG12wspXzwN+COzrkqnGLg4
SYIvlzCBeT1vF/E7Cz9p5CDpVvfFDTzYgY3671+agV+PNRjh8Z0m6hbrcuFgwoqg
OWUyiH4PDxzes0QbXJigO4OdCZp+1/ddir3Mv3jFMTAnHk/cCKAs5ljVUkFudtDF
4JhlJryUvJt9j1vY9aPHYVE3BysDX0Fk0NGjTiSUoww27XDyeAkZPuHwc1JuYNeN
9mbDVrxuM5KvXpp/kI0nUB5fxIOrDCKVUmdOByBzuZYPrt2n65jcznbzyBgzozXn
Vni7oNk3uLkKnjNg7PRF/M6/88FXbGjeBXpUPZIt19Ix8b+jbIsQ+vgEeMhUVm7/
wNEwae2xWFZ7QSe66SZhaen7yTYTY6IQWEtfw9lQM2xtiDmshf+JmsGpgaa8GpQk
7ehbk7HY5C98Ruhd6FpxHssznwOgNjTONtDqXMP0jn9WglO5tlIUcnqFjKz/WAAs
jTdS0IKyIEXhDzE94zRw7YmFkhI8BdjkN7DxFmsJIb6LGvB+20VurO26+R4uUuZN
XJkrZff3zAUG2aYY3Pkr4IwBY/1VbNUrZMwtYXPWWTDTXaszI7sypraCMonsIUsZ
1CNxRcjZpAU/P1cMh30uq6guvm1xgGYhNdkLekktuYLdAohdI/6uc86dWxe90J9a
Pl18InjPrJBjuE5G/wkHrg9LvEhWqy7Z+ZIFSfnneVV878BXsNJ3I9ghhTAwWNa9
WtD+vdw6qrfwLqP2m2g8KVht+RJ+cF+iY0er9e7ms2r+C/fE3NZg4S7rkL230w2d
eHNyr7mAoTqiWefZ4T+YqZ5rsGXzIn0JpSYPBdd1JQBoilNtvWEObvpJ/oIvv+tN
+WcQaCaNJ+FUTph2utV7L0uW+vlFFUWiP5SIDuadadTPYVbPyr4/FM2C3bqyrbn8
E9crS365OojCKd1gXXW/nWQB3JrM2BDsnKA7xBJCxqntd0aw9jkkemw+/gGFqyGL
OQKij4qmq4p81V4hz5qn92Foog2OiZLGzenE1KpLXT4xVngiR7wOZCO+8Kq7/vQk
jpLrpclpNowJJNN3Z9dJ6uqWvEQ5Wqkv/jyFVRfp3deL0lHtY4Gugjg61A5+/SL+
hf0+0r9DtMFbtjUxuQbg7W58jJHMW+eo9HakGDvsl95/4igGpHwWykRsJz40ZYR/
eHmjmKwRa8yzRhNJAOiuGaRQKor13XDQuzSMsfm8k7fkxvisboDPvTQvohCgxsjF
JOtCNIDZ/128ypHAvaXW0z751LAU+FvNxDdcuuq6DrUlAXbkAdhE/v4TMJcVQLxI
vpcGbXve4YAhiGiQ5RL/qF/Bx+vvmu/X5QaaOHFyxqZmjeiYA6dLDC/cBvPlHngP
Nz2Ey1fp3ALmrBFDcdzSe9rjT3TTonHfC5TjQoiPPtJBrczOdDf7QmaoK3GLiltq
y3kvdt0I6Yksv0/UjRietNS8X11EZaqE21liWbu93PEaqTDQefPiJ1NWzBUbPlLq
28d8k6oTKEiseIjtN/PIdA8Ulzq5uGdgGey1z3rWcP5uF5SB35XOCW/xsvJNWqjr
i5tVQf+LlrsuoHUje7u6WfaGuypN6X63GQGJaZcixsa3Vf0RT9Ys2hLYQ6Ml4y1X
in70Vi6o4MlXqDXPsWUH00XZDR+Ll3PchavrLOqehwisRPOcsIY7nvup1qq4aWO9
grnDQ6BX6cdpeCiRS6E+hdGft9hqBiA9jr5cC/CTZdMGt/5+rJhT/MRfBwo+RxlD
EFwuVx1zFd+bwApAUrbyaBproDakMMkqZ3hFwtxyawDO3hnEPEYij5vvjk0Qk+zQ
kjm0HoZFIV+8wTHZwH2z39aWLXm35gUvs6u7G8zcRLQyHqKXTz71qc80T9lOfp7z
joF0VvdmHpx7O7dinyA5Dm+l0w5Milm2SEriuOz05UQVEKvmazu2Ky6Mo0SYMKai
zOKGAecsFIYZl9gCYOMlk97VJM4JkJsAfj/ALisKUrQ3OK24twEnzHpcWRl7umPt
sFhjxYjygpDzNU7js9UhDY4bm0HG6u8m3/1ddTpNKuwelJy6xs05hxFJLOfmQ7/k
paXh12WcGjRcq2ncKJWS6bk44vda9Y6jHVFeCHIDVpqU3I2TGUoxSNdqm1G0ceZO
gQQxUdhdq3HDPd1Bohaw2ZCQRolBVUcX/7WS12S78RJSwEYoKRJSFQUx7/p6kzhS
0PzVTU6NlmtQqlQ7NYH/g7ajJmA78r39DNWRboRJWRLMNWLsRpQeT7Xi89yC2I+K
Ngnwvia5RdldlW2fWxIu0V1lAl7NIPxYBGZpHAGEc0+sEvaIN8tCBW8Rp5Cn7qsx
JiraclxQKXIPWKKmpG7u4C/nazTKLuW6q9GPSbBqM5yWecq5w7cIgIf5Q4W8mQZM
0uF1BeSjP2pV5XNKzg2Ik/PYSGeDdKTNTCZmeGgsIKpCTBBJzZmXxeCO29AChIQK
3aDoC1COM/jesbz8pJpq3PZUpJy46V7lV2BFJBTVAnh51IVctKtaaMiz9L64r8TI
jbcA0oHBVLTHiFYxbGAJA1RDq64GWJOYBoxBE0Q+jRe3o+TpjhbCrd4j4F4PhcKg
HpwstXSzKa3YVuPgC0Hs54fINehLz7dyqruuuewQAQGILJ0Gu9hbPDKzFNvolVjv
0OvNtW3L9oL6jPLmJsFiKecdC0Q+ohWVoUJTApvKiIj/SO1ZG8P9ImGwHABOtRaK
xL3oDGI9MDW/OH7o+6SX6p+1FtBwViNMuuQ9J7tq2y9RLtSxlHlox3WgBZg8SAq0
dYcjDrdSl4bxPV3vD1tLrCaL2C5F3pUDj5y1j2s3dKZsXwPdVRTgeJWMNdi3/ZsI
GP8tQeQ/LPXPgSd3QOSmu0aaho8DAcsEY42OM3QsF9XKFauJzMjsu8wkzTBaF8ap
PbFjUlDJtoll9z6wa9xKZi4LBPzTSCJBVYRsUVT9pEH9X04xw5gR8bkwnw+Fvi3r
ptw1A1NAZ/tXWgvLW0G2ZRr34uGy7nfv33TwTP8G387OGc1JIIZvekgr18lm4jO8
aI8sxLBp2jaBbh06Fav+fS/CKRhHpV/l25guskNAjVb1CrMJkhbs20nqrw/Nbtq1
ldSYLJyZIBK2dAlUnrTRmQAkj9ro/P/owrdvJQVxBKhtWzgmU16RD/S7qh/A65IB
2R8L/u5DaSfom0ZDN3uhGhazMGrw8vyj+F1Dpti0FIq/h1JBvavNaz02qY1ZgBhc
xj185RlwEnHeE7Gsmmivos7t5gy7qf7NyiNOWWowVFgYTSxbH1TQL8DuiQis+n2M
gTYKOK+Pt5lE4VmHk5nVRwAxe4Dlb+aXPzCZxycPcGarh+JVQOAK/M3Xp46r64TO
I3NqpPecGqY9UeS31Mo2RzjpHAnvAotV5JZx1k08g7zQ3DYgTJKE8ZscQjTM+283
VLE2ckwmv23k4rflzyh8cELpZUXQmAhGzoMr1lkUwxNf/YPN2SU/A4da1HcvX6JR
Qw/F77hAM+OXmr7AaAK7NKyAZoNhp1vsvefDi714Kl+pDXAFuEpgxUo9RiXV96cJ
V6CFYCZsJCbtwEx9wKRx1/LzZ1erU5oom/BNQ9MK2m5QDb91Bh3zlIJim1p2pj5/
IuHwcnf1bGEclu4cjchKw0JNHPeATG1xZTg0ofO6BUC1Oz9sBxOAp7O4OqrCZSbq
H8bH7X3ToiR9gtttALlDvBUmYKF5tQfLkHeMbmaTLzWiTcuhDzhRo70QLoEdzhNX
jaZp2O33lWRJHhYskbUQcYdCQ1Q83CMQVD26QxeMWvyhEvoVHF57JGKDYUEfZ5WC
xs9Q1X3J1AmTVqZg+5VSGBde+IBM1vkIt6qqdeops6uvmTwpTCatOWYj8S1ZfqlZ
cvTZM3sTVM6u8maRHhejFle/+OgPGSeoZutuAtWPPa5Ogjk5CkZFcLg54XLt6S4K
yTGhZppjXoA4ZWlUX5smUGlbkCHdzoH+5QcI/8ejQu4AFYuil6G+0GYWbalvcKaq
CTFQ/0hZS2VJFjO+Rku+o1ire9KfSwTtbFNPQVX1/A5Y1OXZx1NM+5jCrSnW/qIh
sksxn5x8AgDmtd4pDoIVjUpIAOKCb038j1yzQb54HcfmJzLu34Uz+Gp2MBlV/cj3
M13hGbyC0gkSS9LKb0nCb80k9BoAoG+mc6ujCzgwCC96LjpNKUvY2nFkSVj4GlIJ
5j+LbntX9aK+tyNe+UXaRZZ0QrT6h0hmza4mO/sIltGNpazp0zscyrfXiuB2O78r
M4Eq7btMZTMwIAf39Foy+SVte2Q+VqmR5Vg5pWltTyjtTgHqaQifper2UTwzrOQ9
EegiE4Wu5USdP0qjajOlXi+3U2tMMwQkgACB6CJP+iljWYFKvdi3TlErdqvR/C+q
BqXA8ffw44kqNoMbNfUPGDguME3+D9Usrusu8PqQNWLnQV2geP8mMmV5hSrt94al
G3Ugmjd5L3t1B6AqEcPGOKrfUpEuphAIyvpHwN8a5Bhk16k5I8afqi6XiDhSf0D9
2oHEjO0ooa1CyzOPBvHeV+naKzpKtEA2PAJAOSD6A2EIvbUveVfymcqs1hMopjav
kBgIQmEqq9Aoj8hjZZ4HFczObhIgICEB+X8YzhwyyKMXFub+Pui63RS/samYFCN0
7I/IQz0qQ9EPn6jRQveBSTSUSJOE0u0khqlWoPDXi047rLNvNoFvemD4r6GV2yTH
hXukzfIeHXFIe03Z41TxM207SxXXnTA625sbbHuRDYOyEg6I0Itj4E7DKSQg1NYg
UIp+P45o5tyJ/eoTBAuLXcLQho5EjbHsfSv6lFCEeW5hwmOYruG4Qs+zsqNgrLWy
m3EHm+73EP7RehswOgt5HaJily06EgBt1bsSAO1WEaCSzdypQZwBfexJodlwt/TD
O97ImM1vJTfJeaK0EjwcmXIcTWfDrXcr05g0XR630Rmmg3jpOerp3xVPvWd5pV/N
1WZzB0VDpltZjRiv6ha9Vwy5xdlq2GzyF3IQwfHf71BryZ6N5U/Ieuanv3JZZ4yw
aAmihzgjJ6jd8Ahk8kjzKN/kwQklKyp8K9YrDO8tVN+b5CAWoc0CGUwV1tpVGhzv
5WgUd5L0V3IN5w+pXKHrrcIn7w8MXIIp3UGzVGIrSI5YvMd8pKdloFdIVjzHANsY
6QUrrfgtdSL8SuWwmkiizwGzvK9xFtlkjmybOuajPPARrnI3VAhKh7W9r/e8D6o7
s7SPy4BtGhRS2Y6YosPGZbG0njG+A7zmueiGAqwh6Noff6T1X4fySuw6bxz40ME+
pxQKw+QA7mbxLWTvdk0Q9seX1hEQ3poeI7ycfVZafEwZQdPfnqZaNc8xGLCeiClQ
/0oOsnqF980uhRqLFy5pkB/8L8HZczuwh5KEZv0NeNmJzcebsRamBBdUkOvlGXvX
hJ7s0GDP4EIkWEkUSB/ajOPQLpTSXN9ca3LXefJv4iHJ+bO8bLjSd4g+PzyECzQC
Tz6bBmdCLP+OWJnm3Zv/gJlF3P9MruPtZT6Kl+sG6PeQbX+MmZ9ge7H905Wn+YMN
caZF9XLjep5j/fj/l/glcjhjy9p7JtMBIEZ37UsJ/fCr1XTZ1KqQyeRe7zAUw9LJ
GFut/ugLKxnXumuH7AnDA/dgxHS9NhzSJXUJYyCBoD7ireeB4afblsoCu0BtU7f6
L10Fu04i+lMdgSGDEtte9aWWHn7UTiBpq77+63wdnvjnrVf9qMjcb0tzFPxqQ9mH
97fx042IaZ+CgeOGKjKHi91hMjHATIPxV+N9bFD/NZnlk89Im5e0BflPUsvC2E+a
eihP3jgU6QDGe5B5WSsJywV2ckL1qMCkfXnRK6lMeEBO4WejmcF60Vs4qU/GB8Vn
95JP2ATHTbS0IeA9vc38kG9acntchc/M2UgT7sfkPJX0qj62mkqhcKpgoy+xVqxX
GV4FfA6QTkTrnn0lPmsSR1bI0nsSWuU2JWpPHBJTqPrMtajaURUJOKt1udl19I2O
M3WWb9/8k7/Cl2eyu79yA/V7W6L7M2YK7qXYkw5ZNIOST1xcM4DKCXmEFWXLZJox
oVXi3zf4N2u1Bq4bRBCW4M4wv6cBMLjEvC3SRT68zUcHzdbyVS0TRMtQMv2p9/2B
PPMxyPywis4GreH2CwrXXl7MK8sYKxfPiyluplzD4U0fV3CsBYQ7iDY4106S0kVB
MK0FB4obZaZxO5estTf8RQ1PhaRM9aX10UA/D8QQFLa0ml089xsfy/Ct56sKWYC8
YbwoZ/YD/3ksEwH2m9qK5XW48LUgKNG94OmSl7F1c5cHa/x3nW9Gl4I+RjgkP6uK
3zgyZ4ztWlnUF74aIUtZ5UyVoP+0R51vmA5/xxmBQnPAUDqBPOhiq9veyhBdfW22
P1Ta2wFJ5iAQAVk9K0ZJeRs0XkhFxvB43a+ByH96vqMgMgsZoV69nttmvWWPyuj5
n/n73ckvXhhNExrIms6x6jvals4xtEfVGJn8A6HiPVv7Z2IKevR2NjmQDKCeatuP
bChXvi5T8SgLd3RgScPzhSVTsC+SWiLcoW5T8nS5+OFIAiEuCtBE4TJo3LVd7k4y
bRNK0Lmc0do7uT4UdMAMsTepQJz7aovb5fTx0SuQQVj1y478qGZJ0+u+iK/AbzIp
EkQ7LZRXgQsP2IkCh1tKJgfc6mIpUx7q/u01LJfhuXNoYVzfCWhzPJtZ8PoKzVsY
7xGesHUuOgncRZ7lasVrsPEzdMqt2O5rl6c2i5Ll6flyYkHh38k6N9aGDtdXIiu2
MKE4XzkyE81S//K1IKeTXPENY8J8USW5+nbjMXbSfL+SWMSWwUOf9wGIAxuV+nqb
TsFofkXDLFO7GvahGrlEhzYucHfX0kkpg2HtHVfO+BTcCQpWlHSKJm8vEVbByr7X
jJDJAts3XovK3tsRz0R2ORbtzVmZGVrvEac3kyBWRPp3y88cgOmE615I/kSgExyC
MGsi5POl3PjQqT0z2BUwzqHEGpF09mi8SKaWgeCC2qV9VzyUapyBk38hh0Ml8F9U
FLpaUG/+vCOsxj0Z7PfS9wUdpkjEPlKePclU9q9Xg0P/ibEaT0gF7bkKA35ZYy0m
tr8M6EpSee1lwnIPWYdX9aVCFjLX6y8gwn3d/WE9eIX38RJj2AiHnCfPz/Lo4SeK
knaVmvpXRUaU3NDd77k5oiO6vTA9iEL6LRoAznFnT2kmGF4Et+zAvS0xi6wiyP+C
bQMoPQqNRgi9usy6BKgZL67HF8AvlxQF5YNHyh8HjTxCR5tXGHhatF+nFau1Uiqp
SeMk7OMX4Z9P4yR47FpkkR0ciNlGvZ8IW60TsEMa3quLKLYQRfbgFlX42+bRt0YM
KqkB245+EowqYP4QDsxnRUkXWDft78gzIusS7gV4S5VSZizcUJxw50XITOrZ3Fv9
LG9lXxvI0rsOJ40OYvmIWe6K8DuTFvWAVPEHA41a+3oc+NKKqgHMbPVNHrTzeQkV
q1QzTlOVp/UIsMqR1Hb3b0BgJ5mIlEd8K/nVs4iatjHq/5qCM/PSIYR0pTmKYnl3
Q6wGquPYDhL6bUOdVGX/XLZiuvlkH/s9R4j+3r2YXICTASLiwJ5dBGhdS2BwkVJk
+inrVC8X9+WwPWgMMO5ZvWt26IcSgDbAZBG/uuUs5El9tHSi54wpjVp+4IrC8ErG
USc0D2FTvkNqsLBw0zPZJSGgGdAuwnjVZ/qdt1ZKTZ6n/J2wqIIFld3a+fBEfrWx
VgowmAee9XUCTgvq+uZKgVBE92mQBkyFWLSMB/dl8jJSJhvhsO0lVdAP07rjPTaC
c6TZHnGG5TlwUenQkwniU6R9KEjPNdHJ132v8V8MdrSPETrF7RGUSOoM/6+q0yXA
z+KlX3fpYFqGQIwX/DQHY32zIWTdQ7BoI50y1Sim6IAT7VtfGOYyxJxqhZg040SN
qsbGiCubZkpP8D9F57OPc5ArhrRjV/qLgx4nKBUh2ROtdsiA0gsV2e6pmzE5DJT6
aLlXgYz9vaMmzl6rSWJQ8aH6BWrDYRGzNBPDQIL14SrKo0OptQMlvW/H+zQySwAl
+RMTmZNzLKca8YlNYZxPuHWIDBbP6hV9GTE4uGSQYMqloZkkKNWthQ+RfVVyLsnm
rm57bxLnQnMTsjzAd1MAdaJQnahCsunt/X/+6+zPtZYSV1R5IAScmY660fUZqlwV
Z0g6Wrc7BtcC2m3JJLF6yjnt/KB+X4HxQJZoicUQJqAXgqXvF3heyYbBYj97vpw5
p3+D4Gmf0jqVEZoU+BEm7JSy+ascx1Jk34z0JwosZnOHe/pgeCEv1yHZOhrSlPpb
ZVHd3nhm05iVz2Ip1J/hCulzxyOnVW3DfFk1l5Fj2YPR72+u1dWmgv8X0mAo/JRI
YzCe1k2eDTdl8UHv6k2DPKTqZ4LSlXwm9erM5Zv2RzW+UHyavgdYpwEq1xlamcmq
hVArpwtLVzC4WuF3nz/6SCq/EQCoKO87ZshyYTLIPaPIkvg1VjbtN9YrZah0qwcb
NI+GSOx/tLeSWvbcuUY2SWJRz3CfiEsHNSBHjrMv8iYj1aO2qpT0t+EHkmweUoeQ
bz0Z3vvxEssDc2kU+8JbshjGi+1HAGzLt3pdWrxQv46Z/o6z7p5M39NkTrFQaLag
nTPoXNFW75xNKboX73lBBDt2tkVjneWmKaDwNLqi+9XNS1StvVYNVVqepQvWVXXG
sYuM4i10Db0GhuuYwNfr0iytdId6SvAD/9lwXRJOhd1nncWsXbAXoKtG9NZYVJ96
8gqleQrixBk8LBQIr1ZiijiWwbkndH7CmEi8y33eT6luAF8kJ2Q/4Q3tdUpNPC+L
yiSVoteXBsBV9Q1e3aTns2najH8ZnLxEqkGqtepCpMBY/ixBWPIpHog1IuQymGpe
Ku8yurM7N2J5sjeNY4T7EhUcV82euudzJtogPodGBYxuMvyRGMZ7wLYONUfoulMS
57s1U4hJiETnQBtO6/kWTaNoCi9+Bwp169QNdgzd163PgR0p95NUMsMmTEvTVB9N
cUhrv24dpBOANT2yxE6fxdJ6QvrTnWNPRNFOGdh0GFmF8/kN7YgNWgyTS2snR62T
n3MLdMvWue5DBC/vxhKQ1lS3VYQTdDFUnCLzqwnNxxhCm/xisOEQWn0m1onXCWab
NCIP9czoMYL+hs7wRH0sCxNbfuqNbjY6VFr1OsusTlfYJgXTXGoGfugySK6vhv/D
rqC+3qhKVlWmg55uTqiIBU/jTKgeLP7sb3aq03zRZut2IREummHQVfE/TcJ50vBc
fXCJo89Uf2pbu7gp/2IoZSuV1a1qowzh1pYtS93sa0Hu+n1kmZVO49CpdIcB9R7c
sqPtuktTMlaOTb9kR0t4EYF7n4SV4pIHQOVuE7IeEOR+pq8le3NZYYR3D9VdqvYO
JAH9krbJ0Ri1/KV9Y4Yg/EBkLfR9WK0PtWBOKnEJBGUq7vVDCdxhm3EP9x7eXgp1
AFiWg4FQsOQt580M6DXotZHhwDRxSx0oFGD7jRN7UIgR6aPIv+HfiHqkft1rvyh1
N2GLy63TXTQr01PzZHpeo4i1c+oxkInfvBXMGLew7uF6OHPszWE1/IXEJ1dDxAG3
7q2bWDcfNyKWOFBDwOJXff8mNOtIlxKH9DY1KRW6N+ugttkcmH1kUimOg9lO3HP7
5ReOrueMaZlj2hjKwzPNB8cYt4VJ/ame2mBF2kpMS6K5gt9BfrfKrm+Xab7ymJUs
/j3sZ1lq7wQpXpDF6e0gxRWGfboj6/5YWlKuVzdSjsckxLLVqwV5GJLzQWXpZvbg
KW7IqgqUzw08cYdN0R79WDUkKVoTCVrM02X0ptp2QuelCgsFQx6W+1d/0HzyGoJj
NTKv6Gbgws+uTlPN3ovdvfMZYOZ034HnaTFajNyiXOZXsDs0hB13YRK531eo7bGT
IIJvMhQpF7FcX/950TMqe7m5Ox8QlTn/kX+YiJIAuhGrfgGMngUZPnX6gUdVS7vs
0XAf5Rxv6j4QEbi2FtPZumrwv/hauEp88oaNkY6wnMQ/WyZtFJp49I34u93K5o7e
tfI524wMW1zIZYe3NqckiFemoE628YCtsAbFujpvArtEiQtY69CZ2Cr5ZXuyCkWe
U4XGvtJkEoXKPzx6Q8sFfioRCNWjBVE8shfGrkseCHeegWlBByQkGw7Q+47fbG0D
DwBm34XmkGLnULNAHjs8uaCwI2yZH/VFPF6+V2gqUPGF5RcCvEBMuc5cxpw4uFeA
2npXIiTcUKO1Q2TD64fRt9F5FgKyAXqHUDg+vlegvhbpZeDK4OPhFfRqalybp04v
gbT3vkHLiyUb+JVdxkqEGEsKBz066L96svD6Dq9Tg55ktq/tAMcONHoMnOZVV7XC
qkyjhlI/BjDennLQu4L9om1u7IY9R1niKJN7eNllZz1tKAmuuKxqsFv9q5duOpsD
8JryzAFmk0RWPq65Cuks8STQiYn91E5NNieBfuQH+UZHp/+Dg8DE6vHs4U8E50wI
+v5iDAVrNT+n6SgPtk7Xb2AGz/bA0No9w+XqmLAxjxX7kPIlqeXeGjYPparea5rf
+pRrAUhcYr+ceC6WoUfpXNUDihtb9ELoRwyKNhPRO1ZdFCCF5GRio0C7tkXn3BIK
CGMgCeSIzV27rVWpUjgOGRNAKcyMUFj+eWUDmn4Lq8fObS5J1eJ+XpJWWVvxY3D0
HaC4/sKMu5Z77W1I6pPWhAVxDFlcQl1LA5XR9/42K0GEikOk6ktoo5FK+adYyulv
Oc5s/UDWv5tNAkzVmifsyViqlzIlf+8qn0y9tA4aD5+pfcWEPmTIJGIqgtaoI453
dJ4lMlgl3+YHFNbhDU4yZb6hScquZ94eQ4y3NAi8Fvey2UQJ8wvHQVIvz16h4G8S
ovowpF/mDBtY9mPdXPg3R+5H0glifda9RhsD0WVKGnu9IAZv8GElXJFfE3pOqSrD
8rLPOw6FvuiqQlhAkljJfvLvLlEhl9pkwNNEyQTAeFJjJb3ZscXfJ/743lmddsxd
ha0NnmaPpp9LSj/7DxLPlvEuZXJl/j1MqeZ1p+CJNjxnEZwBLa/c9yJvXCQPx0Y+
W4hIoEq9TeHpRze8ZR1e3rNTZJwUXkzY8j3UkdVSam+ZXz3r/stGtyhuvVSL1j/c
dpDoM3RgPZtqhRW7QiV9nFdgWyfHz8EATFLe68xaMEVLcc+3IipkL5JafHbAijNg
mwVaE5NqysdG3cs0zB4eth4lds7fDYKZmkdWamQbaHwNeBuYa4MG9TjLE/Afebsu
ZwwswXxlLOZeiuYTUdgo3kuGwjudl+PniXsxVRiNM+EnHCKq1PJCYXv1lSSFpEUs
DLpP0U7RCTrPNM3Oqzb9kl6GBnXl8T6ZnOskqmtXHJfYTOcP05gGUmHb1fy1dO/U
uWFqX82TN6HJ8t0WC66QrOL9TjmNUw1mRKYKA5kTxz9lGDeMDLAWP8jTr1/Ibcm8
7o9GyGkpEECTnrPLYW4k1gXVmFUUM+I8CFwFmncCtjJSAEdZBOm431qBlTM6FW29
/SdInoquekAu6g9kVTkFUZrH/ItVWSMKUg2EPKjPApsK2UXoMH/MUNzYpjDy7ktG
5FFdLaNuvrWKIFoVHWtG3Mwrjp2wuxfqGpRbZYzgFaV/lUiLzgZS3+pyMmnKQtTY
0aVfFdqjNuuaQupKaGuaRLUaGZEbDYzFYqX5IOqCZb9CmLwMyYsYekLqnH6JadXm
TOYtKvxuHrXK35GY022lsdeXw8DDrM7KUIMUFk6rDY8fmcIKPd/s6lTkLeIrnBQD
uMplOujol0zeS36RWtdYBKS13QSaKghjRbLi7ph97URr3Cop3HdKsiNYxLp8hjd7
NIWehX283Y+U/rLIAkawIJ4IOWpcP3so6uEnkyY2lA7RI2FuU/Z+6kVosLqtwl6i
BhK/1tlEW5fm5IzLz6s1NFEhPJSDkRXKjeXwYEOeymCNjl51Y5NRfAQqKbnpz8dl
aspuEk8f3fwZD/CKjnhgIoh593yIlTAu9SzAfscn7+0rLu8xxLX0U5SLsxakBpE4
PpfmXUFH0gJO70BKugnzc1eu8X+/M1J4L5QgfGPo1aX41ntOr5Z5Ab6qJKHWs0f4
77ygIl4PqoRSey4gN3mLAz9vsnxJkybz8ainKScA4wYtHpOngi0sqI2ATKVoCYAK
/16rq462qKIqJbLOpvw6O0PF4u6xVW9idqthrpZhykMVdVPYTQ+uwy2yORSJMIl4
2Ld8CAzDi6HaSo/Kz0BEVXNAvPGRHxSWA5l9FixPMd2WDhg5OsZ3oEAswSO3OV5j
0oiKGRt/SocJ9Qi/XxtDCJC3VJLlZCLB3XPIEyuimWVzhunnWZXQhu/KEu4ZyLzB
vHvt3/avCu4o3cAYPj1BjvxSgFKbAT1qZOs6msecVIWJiSJ2Ryk+NkISPofopaDk
z06Kig3E/3uogONV/jxH7bLFgczx8FiwfgBdxqB/dD1o2n0EEm/YWfAgFFJbs1LD
LiKEKB0rdMf4VNDoa8R8u9YRbysFF2+xewL1Mdsf1NSD4td/v8ZbU41imy/yVLmJ
Uwa/qpc5kKO8vMfP4RWdmq71EKWqW/hAIDi15qVdNfV2iTpl4ZpQlXK+e2WCf6B4
0OPDEP7uaKGD3CqjZ4OEhNED/KalapXdCH2tNOVaJzo6AU4dHJbDXLZ6wpe981AG
x2QLREECx297EWcFwDF9seMhO5amxIU2b1hTUq8ztUbetAmlbWsKQUaThDH/I48o
bb3oDrq++oRgF5iO4u5IemYIsUBVNf7aTdXki2n2ATwbdqVPVPM/3CluXS4mWEkr
ExDwWuOrxsB1PqUOkAgxW8VTf0rWeUYois48PWubbftCR1ntBmBhbQdL+J5brbCP
JS3+iFkTUruwo8XcaLqT/bWq5iXyoULb1dQipmyMm28+rhMEgmRtutNdrCNAihHH
bGiuZdCR8bVqs8Xz3WP8eV4VWJ+01vivsnUtxfmxoiz2csQyTfUBm5YBE6us1nh+
H7rCvn7GIT2IhLhPATDxEYg3L2/yOhRiMKbRKzL458vpeR94un+mERpLcbpv0EVo
Vr2q0PWkXTsgLmjYHWz606ZS66wPR/wSFxP8gMHkby6eIAQOCNyWKL22WdBxg825
isPCBE5v+eM2m8IihWTZxLLVUnNNjWuilyZudkdmMw0YupNj62Yc5p41h/v1WIL4
HZqYmDYMXyYMC20fkX1Ie456n45Ywg9GI+RIaWI5G3zIFRW9K0iSNUkiAN3fakM9
6mbjFod/xp/tGVYZnqDnILFePRMFdLO1a+gF6OBS024gefHGVbt0mh4GMews6Ojl
wWmCKesCyAB9k1v1Cgqg+jlzqtmn2WYf2swGrgO4umSBItnQJBonJqbjIPhDvt0S
tLqet1XGSSsQ29nlcNYD/es9GJZ0veZiMqRtTA2Iqqah3Vm23hqZY++pWw+zElF0
NcwNRW1PE6uc/5UIVtCH4C33N8HMpV8hWXDxJb0VQhdeoO6EKT/iPAnt4RSfTf/U
nREunEYdrD+nhQQ0UaGWat4OVMZ2G/LAoxlo7SXH88d4o8VivKydLzKH81VVgDek
wG2tkTnKDTE+FZolHMys0cAN4FVFC7ESsqpdwbJdRVi+jQ5m7nQV5TPbSPUEFTdz
pLFHjRZe1KgmCI3ZwGVk7xXfkFLf4GuG2IVpOHC2rMLtPKKHffNsEliB/BrKl2+O
0qG6NtNAyANgkWSoEsmpwjRqJQmXr1lCJQLsWYcmzIyQbnI+lhTCObxLPVI+6w/w
U4IzRxpndsuV18KZIguFLzoTqvNbl3CTw3dIpvuzylLEpJcllQhagQWMXIxVktm/
3z+6r/kvSENEPoRPaOHR/JU1QOU+Oe+clZRa/L1by2suLmeA3gHh4VilAPc9BrlJ
fyqEsF6WWRWFQcNKE2jLPJKoaV3ilEkln4ZgimpOyHLf1tpwlTShJPxFVvKY4flD
uhM8DTaYi7texPggxi5a0oRoDhCTRWETUx1jN4n/EmK0QLsGNx7YgRyL7duLQMeE
6zLfuQ7pXaliSP0SX25kc1WMOGi1LaEQcKTaf7Y+BG3KSkCv4SXN/ucu8sB2+gii
vDjXaisQQdveqRY0T4WzUcXE0WbtVlKnRs4Bil/8b4gryiT5YSx3CZVqWIS1Qi1R
AAXcffmNJi3NfhBWFTfmU2I/9UugNctV/4vgU8UEW6v5mISCoysyGT0GF79+T1Zw
HiHVTqqW3nX4SuYDLaj9G5p2Kzp/0Gt90SFKQYsSHhXEm+c2H3n7Ld9qgqRaNHSB
sj1wr7nR8C+48lu9aps4+WR4s9PWTI/npKEmXWgexrjhAJjqTOwRpfjYoRXzJ6Ny
RZx0dhCfu/f0cwAeLdqAxuI69Xopez2yaoQ8EtCSTk6Piv3RGjilY04hPklCRX66
YpYB3SxUFyBxDDnpsKTDppRLviJDhq1IJR6hK3z4SgDeLxXBLKjyOWxPDOD1nsh5
f7/5WlN6KqzQC+OWyxUCpoe7TiObvBUQZGZIh8NKqwbeADDkGgVwKmRNoCCRq14i
d5Us7rY7s0Ni4erSSAojmR5Jy+5Lo8XCG7/yMVwTDGyDWa3MOlB165FxpdaBIEVJ
hZ4933txuGVqvMe6xtozzL5jNywpk/5eCzB6PdWjHuT87k2Cwhbrbu8i9vFGcXtM
o3HV8eX4gyf9G4mKObWdmeqNhE9joXOO1Wsl6koeXfE8S7n8e1P2kBlNIoljzHDH
PndHCaatTUaEQv4nNVi8AUHs5EdYbGJ6p4SI/TN9UGfBlKFpgjggOGeUoXY6Tbhh
dMppjqKloeyu9G8TUMFG3XhwDmN3641G953t17i4JY0BkGqBbiei4mXfPVs+ynU2
m75iOyMs6qD4QlhDiJmUpVSaKDwrI+rHK5I9HwQ1kBNwlFAl4nquUlO+HwXhEwtK
oy/zAJ9YgI+YrYqmS3eI7MUWLwdgOGRH++6im9QjhG3NGfqDij//XCrOxDwD6uzm
GBZs8bJdmz9eDtbt6UIQTKUTiCNrvqu2dXlRHLF318UFc+R0PkSpoOjhfy8CMU6T
R+q5ozJxd+LUwc/Mw7DDfD5c634eDIhb5jbR9Ibz6h4o7/85mhEZx4ENRaH+jitU
r0eVitwemTqCi/4BwNmgncteJxBiSsrQ8+Vpjz1eyzh7CrfPO4ZOG0BZXUQsKWZE
Bv2+lEYGtH0Q7m79Bnt0TgdMsz5n4XyqluURw/6s0oF7zCRgJl7cNEbl6l8EABYb
9s3o23O56PE2C4sRrKisfL6qtnMnkQkKWCZTmMNDT65LtOJm6ik7PUaHWc1dmMf4
ZETj1TEKhgOL3hkMnAIEITMDBfN7OZXsLgqevN37LnxxonXgSvcV8SunwWZXN8Z1
NjUiv/5c1sfJBnDff1eOoQkUZGHQvocXYBYnfWdKRcQUGl2BGgVvUSsTG3YypbRo
VtLM+Nr9IcvBt4o98lJt0z4LSIBXcfQJVilL9898mHMb7PyFVHYM9ba8i1TNRDXo
Fy95eJxiokt+mUNn4/KutEnUOqpZ6qkci3nnm7hh4YF6fk/wI/6V1GW66WsfZwdv
vvvdxv5ir15T/aINupxowG8NLXlpX+4IdcNM1ZIvyPnH4/VM63JPqWpoRC6f212l
5VEtZd1MYwdMuOObgUJpiSH5Q8cA34fP3CQ1nD4KIb0LTPkPReFlnRMnLlWs61Tb
p4/a2v0AYfBYmUESCufkCFbqCKFLFF08Oyl5K2S9wUr1I7K3s4tPk/VKZqCVTFFp
Bjt/8giHDDNSe4T81dEJdtrGE8wdZKqFacgxEx8giaIINJDEHPdfHZ3xqOj0C+xF
Rn1qStn14thZTouj+QO1USHtgMCLexMBA45Y+Q82q2QlLFqn5NI7VurCCWgalTXS
WvROvYYDX0AaV/3plQ4W4FDwTj3iZFWnhMYvmw0a48Q8vw+fYnHi2m7sc/cqenWJ
EQ5IiTcG6r7PkvQS0qhiCKRPJUdNUNqgbH/txtH9LE7S3BVNdQoazV9loFICjmYT
MpUTWJu+B+0Be1MxASVFrSJUkLzRAM9TE9LHAeD4jZemvp1ESSzWIeXk2LLDzv/N
7jMo5fZwITrapMJbgTZrLVNlEJloHr5u9r+rBS9qE4iRCqQbEMXEZubeixkqM/yU
3wMoM7R3A2m1mGee8av41Qx90rPoG6VRyUaOJ/Vxjb41o7uzFLz4lNOmE9xFyiSJ
TRItZvDrtQZFJ1lNjH90TW0dUjZve3yMutWvgoYxqj7Px1E4JmtlYoEjYZ/D9zWB
DU7JP+sei//so6waYa3YzHZ2L2axEL13Ne7UHZsVw0gaUST5NMA8NeBbMpXPlnPI
7SfeSIwr3FSc1TYGK93dchh4ZnarphH70xME4TgQETuvck/SrhCrt8k7Yk6Or0hR
S7aTSKWjeYezbRHGHSSea4sG8AfD5r5Ol8tHFBSSaIGvHl6NGGAJn5pP7Ks+qIaC
jISUqrE3VrVbPB7g6EWqCujETBLizV3UQ8CRlIzV8YEndcfp1iFJ+6T3ufBwGYt5
SBTU+x5HkOhWMKBzzIpzMwvHe3wt8aLlML5Ak+X6AemobjO6/dmc/77ll6BDN50u
hCCq059fFuybG2zCOOnOHlDmCwkb9beVatwoD8SSpxCTa3ChzNKL7vJv50VLcBwE
HqVDAa9X105lZKfI86nL2wnz4XWXCQGPi55yJkAYsxLjUef2sw7WlDQ9ekcSOVpn
bfLUy1c4w5n+hFhMVgd5gLJygfnvXKNm6yOMfhOJRPo3k+/upB0zhRK14ElfsoVy
Ft5eHWTClXX4aBbXTRKxSPR3oeW0w0XMfolHayZdSpbq4L9aqCJWv0DtXWXDJCeX
kdoiSRLaUrXTHjg+V7als2vJyMymNz6bRmBFxIoDZRTrFdPFpKTEgZeoZEppMWQx
pwBCJsI34wlDXzZej8LpGjADiREcTzOU0zxRkiEppEL8Y/awZ1g4doI4DfTj4QnV
XPb5rffHxJiA3BsbcMtmhes85jCD4msVcgwPEGQBtWC+S5wmg1amlJBPZ+WykJmM
aPrvI3kA9qvTotFb7UQrFKvDz3iHWnJVUVX/mUYFY0+YOW7f8bvhUlX74iB67q8k
cjtfrql5rhh9bTUYjR6Nuam5aRJwsDAyREbLWDmV8qzm9+HUjmVhWmgYVhNH6xOH
V0R1jHtxRjRRrTv+I7aRcV59KgHNWwBZAFBCsj3zUWtN1lAyNmczSSnak6vPINsQ
++HEjUvvk5vwwQ4E+kBef5+f29zGTcQol+EltjN2WiKyDrhOxNReFfwuM+2nigPK
BBKhxSUsHLHEVqo0M92wQ4T6TAFb9fuPkLM6ISygOKNRVyBPGNBvmMMJbDHnAIXz
JCWlHN+A4P1wUB0V8UpceXpU5rNM9AU72v8N9ID+1uAl+m7Oi2034dF+fU10kFrP
q+jDiuLnx9ZChorIqtA0CBGsAyx/w6OkoN2dx1kmoypNd2fn7nJIk/jQETvIScSo
x3SQVrUo5zKo0kms6weh//HzaYc9JzmoHodLT8Wl3/qGN/M/680XM5z66VXUk6H7
P9jNFC80za8ScYaTHZDGDNMm5RnqkgyMV3MYE7JTf/shcdvNzLXOOB91BpID01tQ
YWgboEdIUtFe9TYYEyziFU+uwdBCGtBeuJMqc9UzHw1WU6nCMkc13oT+QO7gU+w+
Uuh53PD6sEEXewBu7wS5e/+RJz0yfhQZh+kxZ5oLMpNGaqH/AHWtDW3kwq85Gocl
uRNvzuulJKICK6SrRaOnBXwosIXWNoON4JW3Idh2TvbIJQKt/u1weoFWn6niSlri
ICUHHCu1JO8trMccDN0QvupATSnBdFsPKw4sbScxDEcY6n6vke6sYF7YYQAleJHs
hnSw1/xmDSUHZQNN2TfvhnoXI3brEpZSguw9vi7Yl0N1z4RCptDWgLMVXoDs0I5W
9MDuBR8J8c8wXYloaqpQGXmcTUy5KWBIeVA/LPnwQUqxKE03spfhHi1MckvkRj9E
4Tshurne72hCv2FgV/mJqEG8/nhAGTdw65rmdwktYTmZeUo5oPTwduIW5tZ5h+JZ
yiucqX4ZXmFfr7+Wsc91eWXrnKD7O6mr2fOs8O7583wh2FxQsfZhhX3txPpQ27ZP
dGWCSzGvcczcg5NZobHKN0UlSKEl3W1DUQ5POHEvRMvZ4qQKoOIyygz0cteEWGT0
Y5Zs+no9nLSuSnnHGWIUZhD03bd7RoBI4Y7Um9HFGq5w3BpttIwyk21umqaBdHbq
iV6kbWB6CmEgLctIwQpV3allDIxoufAq06mGL1exu+PzBmAGO8LjsgHSxWBamQkv
HIfhvu/v3SCVxVeku4J79653BIZ/ICrqIh02dVXweW4vQHL+VDkLvkncy79NJERm
n2qNgRwf/l00ensq6HZiJNhW1tt7sR1bP46MXiTEn7iCRieU0nJrz7xP+9kU0nnN
CcnCq45lPsRhEmPnDYW0Ou72rF0GycX7ujlWVDwmVEoxlJhI6BoU2Lqa5WlGnwV7
9JqIbNA19AeQbQV0De5BXrWsSZ2sNGTpHGpOe9VLf8jkWXPrZqy4qoTCtLWUgtPg
wLbByFPMPiCJwkkzQ+AKZ17Jkrr/DjEf8ZFGzs/MC7Cgpm8P4pGpJd0CxBEhmj+w
EtbhXYQ2Q5GhIvFHEKep57G0y2H9AMpoQSINZ971QvT9rEMlm5Rv/H3Q8MjVjg7i
BbT6C8bnoe1LiTg0P46fGtg2PrIJtg3A+hFxoxjM7McZEFBAbO/H/Hm4QTN+qP4b
GI3akxYCsr1g9cM41T8P2i1kUm0nOmt+jyEEgLTIywbxdfXKB+raxFhZbLAO752I
1RhoMizIvqmhAITnjTrdLAepLPTLdk6KlcF+bAcsAC02ms4VmJmWGXojDyPu39+z
pNUdudwJgHS4+Kco1R1JHd6w7nLnWxRalKRg18b/ym2LL22e5Hupt7cqjaAT4gQt
H/DHAmdPwr+MZq04G1SaiEP+YzbTaZQMOpjrAEJXO3d0QGyfTz1qMBpRbjWrX3r9
PVeCz/KbKQjKWOLXkXmfxk2L3MD+Yk9OW37l3oDCyc/kQb1sYO8FsnY1NtC23X3E
b7wmHsYfIjrUM7Rzm75PZLbNlLNPsQ3gkNO9O1xQ8lGp4r+iNa55icTZ8ceIa2vr
p2FnjsOx/+lsUraen0N4sCZJkUb1QgrljtpWPzMZvg7ADcNDyW0pFAXoyIVlbjYK
3agkqQVyrvfgDBCNXbEPWb9zOd4BGsXOCcPy/TaH4A5SLNsLNnqdg7apOJ0vmgN9
f6Vk1zu73W60LBdC0SP2fVzlpDOxHAP4uOf6ZkRuhzv03m/VJIZo6rxDQ/0nY9Wu
etx3oNj2b4WvDuSlYz2dwvovEp6X9hrJus85VzSGlZHR89cntjPmz/bLHs8czRvv
5+7lBAEIJWjq4+5tbj5k3epUnxj+9cAj6YqnRTqCJvLmL/ZIGd9LXYGZ2ZXyi/nC
9g46DKVs1NxBXPr6PtwJOzr+iSBEp3cUbqPw88HW3iVgSXqGZoavI+OFNQ+r+Aje
/leWxbHpsOZYMBomJt2rKEMWrC1VuT/5/KCta6hQVxunfEbOb+Yz0q599LKpkJSc
vymQugyziWFp4E22r7L8BDWJVmrKYFDnW7tq6CjPCaqIGoAKU3LKoGZVXHAGTeYw
9Bkac+b3s2m785yC5wNgsLOX5EBCQsxQ2P16xRxfuERgKR0ENVvYhfLh2OkBiM6t
Hh/Y/Oo8XtW4H0XXetyLyUICyODV3DIM92bgddawAamM3ymlHmJn9LpajdgCNe0w
NqrBX6uGvF7btmsEOrDyx/s8W9Evxn5MDutu5s3sZJXWbl5n3w46wmck4jNltOUJ
dmJjFv58gbReBqbqwE7Y2z6YSFTPrpFbvFRab+IodYdi1JrLwPuIkbpb/84z9W/r
yHTPwopqS/b0CXHaZiDZliizwyj2jZyAAvCSVywjQGWcayRzyB6ds0YtZbvFFfPx
G0e3cpt+0+D83G9qF+6i+BN09+wWfzdgMSv+kLEN/CJa/NvVz4N7uRnUTM50Dpap
H1CE4V9TzvIB/cBqroZlDHh6zr18AUpY2NnV5HWCqE9t+bkua94rf9yG7FeLyBkz
oB3Rt9GnPwlIGznTSjHWaYd/lQL71dpa+bVo2v0EM/8m0ewAkrcMKbpPKjrYKa9g
VSy5oFISpJx70itt5HN7DlTcUTf9GD2Q0AZhHs/dYCGvUpQPxW+eqk0VMzWBYF80
nraQBWQ4sWXbnFP508UgFcaRMTm9eLl2yGhEt46mBs5856BSxOyC581/zcRVwDCS
QQmHCR1Clkx24nOMhI4fBBo8+EA/xIZsQLNGuNUruH4ozGj7iVKGQj8r4xgTqWMQ
76Mr27eo8mfV89LSUmP0UPoV51Gv7yqpgpl/Al7q6l38ARlNyNxUlTgYOG7n+zR0
w8XwGMHf0x5wlhtkeDRA7OZhwk3Vtm5Ph8zPLYC6s5OijSg1EpvuhDee9tedBCTv
k9kURDl2DpmasAsxvFO/ojmg4dtT6K3ieJTQhZ11qOzHzfQf/DR9IJ0d/l3o+wLK
ey08aUUBrjuv6pljZIE1bWv5Dc9otmdKo667wobFRklKI4axC/RY43wmVdXquR8H
epRN3IisHXFl0CMYEvjDc46T4AWyb7SgJvDK8rmENzx9uJXQ1FXNCGLbclUI4Yq2
+rXX8v67K1104JzF4Celf9d8IQkkqd9yN25RVX0T1ATTe+hSgTRyaIRCtOfrAlcC
n/QJYXgp7gayDlElnUWfV37zsBYC72q2o5wuZ77/2gWsGkaqLExclNBL5u9fT1XQ
qwJ7elw2ZArny1zm38XwW/EqQVLsBcfVpdVeVUPMvr/53EGY63Uvy6nKfYq7jqDg
/6layk8jWDRZElIZNGh+cWl68kzS5ev/8LbqPREOF/ZllIvNmDaCqKb+6brU0Rea
S+VCtMb4VdlpQV7J95q/HAhC2eokyARk8OCCg1kE3Pb3Tydo2/eXLPDE70mO3zDo
J1mRa+GjHo/hUVzA8v51K6vRAzLtu8SUxGAmVz7dt8DnAxO8IAiis7dRGZph6iic
jRO+8zzPjh5WBcVwKdlCS1045eTg2TUzjYmkH9/UV2+rzL6RcGyrNCr2qbU+vjGh
kn1JuoThVoFtulbDBFeIWRFcYEiVk5dgo2tU3cSb3dtx4j9Pbycf/zRtMN+WXy/r
uH/OPtkfgIFrB4XxH+trIk+ZYaj5BLCxFth8yHtxqfvbXwI8+foeph334+pn0eu/
w9yzZbuH38m2083D/zU4lBs7jXEoMIVebsQK6sY2PL8u1j1VK5nqvzmTyV4LPT2o
Uas/WfpUfjSGIr6j5+anboXF1FyStaXuwqOD5wiY+TMUoYDPTELChKEMVZm2fi/R
CRj2yjMU5bdGY4HvoHxQO6MIvGP3viihvTMDYbktymVjkbCMt8rKPvAbKN00DrmB
lIINdwyUi6hFvCWd6IfxQQM4/xh/vsIV9WBfSN/6x23JrYIpLj54FGUErtAGQ3II
2cYk9riDlI0A71qwLktjL0ZlifzgRVhrdj8UwhYnx/B7R7hljuJrc6Rk0V+fM9ZL
8Vh2jmfEasb92px8AMSs1QRm+Iq8cS9R72UPevdN7Tb9eNTPQpcW2m/8gT9aQK3+
KEc4kI8XyP+Bb5os2l9sdiWK4DweNfdtXk3OGxF59AAvPMdUe5gDYuJMLyLXdNhJ
VqeLe1u+Ri8lWOGh34Eco5xrT6XzP1ajxL6V5blBu8rhtNSaM+fm5rQlkrYT+BHZ
LGZGwiiW3rTL0CUx8QDisA/WE9sbWTROV86w47u3puzsIsCYtnuWjxYI0rU+ZUq4
xKqwbP//bruPPQ9HBcHqgxB71jcWADkMSNzPWcJFF1ZZCh6+cAV13fN5toPhYC99
ldNuWOov68CXALsSaHNqOCsYMsBSphxGH5up3n3y//ysmHGnC9ykCcQOE0GjxR/2
gGBDi30bGN+0785HYqqvXSqGzRsjDwK6jAGEy3+uL7C9s2ax4AOepQrCSuLELbBN
zAdPTIKgAMvWxmZGeJwCyx+FG1iFWsaNCjYYWQ6x6rGBEg7+tfXD9OhzMP5rKc1t
2zOFzE55NusMHj0kBsfZ5LRN1ieUyydmw/78fip86UQiL0SuYey/aXHDcF4xrOWp
fjcucWv5HwULzfonFLleC/FK1O0k6xu2biUg47J3ZB9yV8kV39c/i/hcnAiZjWpJ
C28vXaLi2yAyfZIadFq/4zKNuDATZHzAcas3hZ6xlja0QviB5MwPqkMUazNaFTYU
CGBnD5+k8o25H/lAigKmLQPsS6z5htqOokQqygKYCHKionlZzZDdUnIzBoJF1x/c
V0/Z2jAdiu8ahy6rm6m9pM7BQu7xnUiXENhQHthoAq9PoSXIgJyosqkIvAcf88Jb
9q5snSI7Ei6JHLy8Z2/k1mfSSqOb726EyyEiO3zo3ndcEx+2fc0MYn32w/Pg1V8c
NiKjuXd0zOmBo55zFzwRIZG8NMJiiQKe848Rv9L9NqFC20YYAczjIWbGC/cOPDP0
pp5PDd2/jyMAm2dwlwURb7ccOsgW4JXb+lBzYvJblTKfmEMnONxHDLPVELX34ThI
rYSYr0qKjIJdzdtuJgD/DiZLa6ZJb6q/4dEjzMuezL4jMKcRJJmfzTe2IQyC8xW1
MediyGvhQexqtOBvKRDUc4mxrpxeZWxb/orJIljrVW0wGMPIok2TYFRgV3EkCzAt
RzPViUs7/04HSovosmuE1pU9w/1Fk3BheyI/0GqXw74FuRVnaBtF3vCrcZvne7L1
4ln3VOKqOkg5gyuDeC4UqjhXOljyLIQty2gOFvi2okWMIUUTjKbHtrwRt4dmSJvj
RA327mL2i3wPXSiwZJO3Z0rQmE37DtJUJvFfFMXAlzpCMHfEUduuf3f4U4z/uW2D
OEd9+2In7Pq3szjoiPyXn+bv/zUTF0Hk+PDccUgVBfir28vm3EQud9tuOCxJtCfA
cdu+VQIn8qeoS7pFgjtm82Y1V/avuVxwNYKD6bAvmJwBUdmjP/h5M9UUPjHHius9
OS/6xsTXeJ64rOapVeLdUU6HVP9E23toht5cXOyXjtFu30sOHGibcak6z39aIbo6
anYgVt02zN/w8bhB2Wspvi49lCX+1y27Iy2J8CWas0gwjbNWiATZH4WpOV9wQagD
0PcC3ksbesiWl/xHkYf98MIbD2PAn1zcTh+5YsF9aaQNSe+qRDGJYJHFsx6Eb3nI
rxjCm1UXqOkRY+Q96HiX0/M5Fpi8uiOX9kABZRCAumB2rogsOjZRxwbNWIZs9lip
vACjo99L+tIagYMFhi+pHEicgZiZomE8P6kRD8ihnhGIJ68M72kSlkOLwlhRcSPS
HLvqiD2GAimmXvHK0E57Oj4n3JFv9TBBynV7jO5dr0LavMwhzOzVdQzBUGNuOV0B
hsglO4iETIMwNF4r66CHhS8NETpXe/vvOHrJRHxne3SnO6g2a6WFRRFkVdImoBIz
u9tSNq81nIdYEgodnvCYkC0KdIwQPf1HT3zmSpCUX//bHbolX3ag1P3qS6zPvb+g
8f/FlEknz9HSjTp4cfepcf9t9fmfO3Gy+o49zWeW/Zv43Z45K/OqZN+Pou44k1T/
sDf3S3dNHLnOz8OJmUJjZGFC46oLi/t3SKXPfDfMJ6TjwGos1jP9abcNB6o/oi3L
wUO79VOTdvlhpC6kNdybftBuAWvWHIJH/VmTrpku0MgBb0su3tajk9VgxrloFG6t
zcXavYY0oMwjb2IyYaNl+e3ciwdIN874yIrxx+hYyPacW/uNGacAVC1bb6tGErce
cSMRYaqjmGuh5XCakrLJkfToPWZU2AJFH86ui8RziClHheITNP5uzfW4gfDsM3uv
OnNW/29vVhlJvk5zeKnEXqpWc2u+mWlZRnlR0w80+CRvH+3xL6CmZzrDaDvwrnUW
ivIvxCUxgaqj35w75JMThcqjS1IXec2L8cy/dxjxX1Y0Q9L617COe8NKrDWj7mzI
e4okKxB5XCieQG46x7HxJhv1KAToRqPzatWuEUMGfPdJfLrvCYW8Sza/PAurHZx0
Qop9ikJkUV0h6Egk0hkZtn+KHFm6YWfxgIcLCyAWP3zEVNswVkdv3erxb6uwbOcb
cyR0mR2qTQJapV2NO78pC0fPIFbGfv1wFqcIZU2PIN+DZlnMFq7A6Jw948dA7036
dnCQ95uf6/CtiKtnoh57h9mNT33ow5pHA5AuQaJzhn05H5x6j1EeWiW5m5PwhWLZ
JZPClPg5CIpFxUHLBb7fFnenQMxN+L9gVfcQ8T1zgqvuLCxGUGYuDDVBgtclMMee
ZBDEfXXGUCwGjzRqQwxz0kjierfObjx8I9ZMuS20lKQKOa0fuhrzLvFDLss4/+7c
HBkAUin6L/QH9lJwQKCm7t6NciY5GDYQIna06uSoShb4DTIw35tLJr0dDyOuLrYE
LPqpbNGWcmynygr7WiVChP8AvcQ4dQkKOgFD9QgNruQBZs9gNHl+GDfc7LCk6AkP
7/+eC2ElaT0s2lH7m/RitHPPaSeu7LgAoYHFMt+0bICFc+LRiHSW0XliG/adHixp
5UcGHwI8aEnje5vPWsR+IvDY5F0rFw6LqRzrP93hU4ut5pcqrnDyeRUkqttfmYGk
sQWQ6zPE4GVDeljGXjntpB1MYEpR67VuYULaaR96VOrMop1GY4ozpcmRZWFiOU5E
euOrDfPD/dL32cyjrDKelLo3+BKEgYTdOFHowlVZYcxIF38o5xyUmJ7LWztG0IzJ
c4ulUvSpPku9GixnXC0gQc0MuQRy19YUaIWnQyrKJSdmjxW2bmfAMDUGtdhIhieO
kvB8btYjXBCfbpy7CdYdlr54+IJIqnSNKJjnLIvwpajGN72RB6JmzzjmrCySBNNm
Z4atIJWc/HtYMXbcMAwIz8655hGeH3MRirZlKul/tZCSc/pTfQTzeg2/+ef+ENfy
V358Vm9hH2uYkEr1kXEAOioKavqa0VYAM6qLK1yMUdpRK5HsP4bfacoHjBzTZW7M
yW6DXI1dGRgbf4Eneiuz9bh8w0HrJByJVRROyDS83ievdZ95aqaZXP9GYH7kHEoy
bN/MMOdzgZAau2SOhYhUdPNIE2FRO+YzR9qOMYnLKDqeOPzh9zn1G+mEAoahVYNJ
VYtveLfEK9VMPNUgoYJxbJYD7HdDZ3l4V5/zcXInbcb1xyiGDDBBwZBuXzWyhuPI
US0h7oGDms3jRAyGxLaR4LxxD38SXd4rRThtYtsxDg2pu6GN3DCF4Ttj4+t4nAxj
MmYpauAADjnKBBvyuZ9z9gdFOw6pL2hKlIquEK7Vkwom4xEB8nisUJa2qkLBpoDT
FC2DTJm6uYe/Ql9kOe3x/JMKQVK2+yAdxxy/wBpexnf/kuKx7WBycZbyk3TAFhY3
xW+nf0QGjDT3fBNqXthM8gsQulyBo2bFpeqGxyFvzy0HtrwJhybWwUINxmlZZTkj
LnqfHHrLW8ueMBqZwIVjcRtPEnxM0KhJt3B7AbpB8Cbxkrbif5mGL7wb0Ca9Dik5
5DJ6/iBIaJmNoiwAqRL3jeN7/cgKLWQhQ8uCdtSXmaL9cae4I2rpOpNaF6cLXADM
R3o9KLlY4/k+FVBdI3wgF1YsLDtoK3/4O/6ckiz2toRcGrv4Zx7QJIwrAAKJQ3RX
cMSlBGpojXSyf0CdsaFSDKQlW5xHYEgdUlVbUJe4xJick9A2QC+AVsU4GOxrmlXz
6J0W2D9rHTRdkJDNlPKwtC2JxtnCJkYNR2oC5mgragcHyjzSnJfeidMICiPCdPwF
MhI4Oa80JGAq056jXvBmzQtCGnx0Fdv1w4KUi4zs67yu3vW/ABzLF/32OvUvq9Nb
T1xnTWyBOgbhyspRM4tX6khb+azyvBol4ZiN+l33FRUIjWcG4lkEvfU6CAY+yord
KzUTmwxrv8vX0EUXnSMYFCmxOQbtOtC5L30NxxBH6sE5GnVSQTAn6Erwj0+8kOT/
yJoju+yZqFgN7l50iMlnnjvgaAtyi58CAiVliOjWa066KQjt41UjtG38bOfWG51B
/yR8nCkvN5EpFyxSv4QYUF9OIVhXbLgx1ObrkQOKe4j6pHyN2gFPyVQczzObltxm
ucijtF0qGxPnFGhlnH5YU8R5UtnWyvgEBvM5thkqc/o4TEqdeCFEaVoTPswkWkAY
5nH1LuxXqqNavG1WIpItIBjgcZ0vqCqrFt0zngJlytbeCHK/O2vJB5+1ky08Xdax
N40kPPrh1TBsUu4NFQBceSVsdoshOmUW0iTxmbT9aDVgww7nyTegb58T53Zos4zH
5ZJZmKz5XesD/02uLPWN2Wrnri9cNDm4Z+uTYkbEbSQSGg9B45sPXlva+/hnETat
nRWjEmB1EGEUVrJJSHfBP9xK/DdnGpedEp85gCz7z+28OMTwsLK0GHOAZ01NUC7F
/ULe1iyyYCLex3QrBNyD7h+DB/pNe3ET9cOKaA1P7zxrA5e+QarjSd+819n4Ux9n
vhf+bOCZAHxVj5OpdWK5hkU2pweaVrw+FL+sVs+ynRGnnIkgTjRWExJ4DqQTe5n5
hMB9hX7PLupWgJ1HP8Gcdw1zNoJgC+vRdcx2RkyQgS+wHmB2KK/c6ex8UVQSIzmn
gPGVn+Tu+f2Kgx1QKS4Hqx9ZZ3XSZZXglS4rUo1p21WOnwr4X/KozSmBHjrBzBci
/zWpgR3B5DVpB9/4UrWi9tO58iDtuB4s7BLVJWIRvoathgaxS4zckxUU3rClaSbV
KmRKgprab2WXvEunuZL/pyJOvUeXB4DrhOIeb5tBWZZDT3YN+6sGA16oG2dMatjQ
EQPaHsX04FuHEb5OopfSG9d5gdAIY+R+WRmKnWXBd78QXnUWItOj1cMyCS1dLurh
kx4+rJiXy6fV8kR/EVE3qzf6a/sNH7iwO8hWC58P9qRwgI2eoo/bM/3yev9LzETu
teE2g1Jdwi3omehk2QOGfbaw8jNcnwkr2TIR8cBM7Hl5NrlfF9r5Z32T0PtOxvFB
9j+NDg9D5mOuDUdZ0BBz7T60Nv2VICH+THa4uSXMJyMBEjywsG75WI8X/At79ZRk
RZVIA4ABg8jwn+cCyjMdRthMEoYV8MJktKoidFgqrGfPE6ZrTSBnvCL/WlshKq9/
2NiwL+tnRiCgDP5b3rwYG3ooZ7uJKJaDOUOCAlN/z2KJa0TW4H4VgAmi17rDULQX
6MDm2Hd/wMZWy8JWueVDMhREQKJSZQs10GMHdEL4+fJ95D1Ju+YKV//JiHZ3BkNH
pt/STDkZYVfzjoDFMJ6dZ8tZc7v1cm7JT5JqhdGsU1ObhXFa3wu+t9vZpPeUd8cZ
wu0+jgaUAh++Vd4AfUhT8OA1NGW0KjVJDSd014h+jHeS0DYP27Lo1AwQVoCiE20H
1Lf/qH4TitQMXarRcRvPUY2z9/Gq0pBrZTitpKgyhgTVPnwTlfpVhQQ8UuthGnIB
xmkWh6vf2zvKjg92LPuzzWah/1x8aHV5kRFOQfkfnWMgmS2v7taLRaxBaOsxicp7
CUVN4OavoQ2b/4mcd0EzKxL1gmRL0ym0OxeRWCSu4SFZEGLQAjb+fWSqtYZiS1m5
IsFkPHAeDekOJLJGUqkHl5XcAmqzEaztPwviTL7qizJFvIsjP/zB/o5Yj3Z31v7X
RkF/tzqXakdOZPxXBHNW5mD8pbMTajQx6JzsRisQc1x4Af32/k2V7LN1hFDJPEjC
mPAqv8HPLiUvxp8z9eSjtysGPkobv+uS+vK0eFpMjYGeEoExjJcsN9kOnkOjDxQv
+I0PP2oWu7IomhuVFvuBGv+eu6ixLuqElCaMVXZ4gcfDyXxlhwgubc2M+XsRH0Lg
eEuViLc2+G4Tf9YJ8ZXdhrn+QQfsq+2mdua4nZVg+xleO/k9sIvw126/Il3breml
TT/CS+yPxUmTphbqlc2BCRdHQkwdPYCozUFFksLUig5W01ZV1OTr2k9BUVvYWbgF
9EFgb5Fd69db1/jwhyB1/29RZxF2lzRoX0gQ+NZBWQ9zcRxgWMfPn2Me//ugutoC
6QQ3PVA9ymd7ZP7EOdrfV3s9zjWHfJryxDdW3P69XwbgT+wk+PuXr/wepDYR2LgT
u8rLicqw9OoMdN7HisxxUwZH/NCCtvwUu6RI7Ws32x0tPLW/FhlBlcvj9A1lONu4
LqKWnuvQtIRZpM6g+7bPACKyS7i3EEp3vTTa1Tj8VwF8fPtwZcbxMwgoKKeQw+U5
djTjIE8+Gw5X2baI6QZZ01ZvqIIyibDweNOqKlyQfnKlglP/NnroCrzoJsFSHy8a
A8cuYe9bg6o6jfipVfh5JBu7llo7gSX/yrhYd6ipfSlZIfC7JUfVSqHCvSeClmPf
0rJjAcwX64axFa+2nRemYfaxmXjUgn001e/1D5KAf42MCBSw2GVXA9zSIT8i1G+D
xj5ieEBpxSVrca96ycbmPW1eBLGSwIRYSaj7ouH4mQm3V81Z/+7V17Y0GmljXFec
+eJAoNP4jI/8g/y0EeRmfvRwYmpbmVlzLVWrYhE49t6z+Gi5c5212WXeg3ptpXY+
OdUwbXHLzb27BoglDvS2EeHuvhrfDMvfYZK/5wYYhyAqR5PlFYquN1/1EKg47l35
tLiZqmEyJ/mLmohfy4gR8/rZEU+HKNSgmdUvaDYILPYucZmQXD3KqVR2vfEJBmaC
aXBY9sdjlOoVqNYnMUpkdLcD7tF+rEI9a5g1z1Rc/tklYNM9jpGAmQyBarGICfef
4FUEZ6Hwbl7HMHf64uxGoj0R0vDN4xqqT9bEWtc6ka4LhLnG0QRnWJA5eJzg9b50
MqfIglKdimmXu1tHj0NF7/AmHw310sJnqA4u+KzGqDr3yo2sX4w2oDuPfS90Z2BE
rD6yarI/JkgBBG6nZnXLZF/a0bc691ildogfQWD9XpmEW/AReprQ9BN3neAEPW8d
VgAGwEoPq6R1DiRQ9kKgbSIpS7thEzkoT89BivXSkSKYNcR9uEIySCyP8DSaPQJg
HVR49c0TNoponG6SMbM7kzxo4Xd3cWkLTMJdIE5Ad4VNtwHQHxTlzL/c+LVsb2YI
jvFxwbk5xlt5ajErhBYxtdtffq8cZSsBzaIpzjGauJqOQ9uOOeTqhkyr9SezxnpX
DoJXuZN5uzID9x9LGfq0WAIIUDcN+wyX33WxVWpdKifBhrHAUXMcYAipdOkFt75O
AXq1fPn0yRlE7LKeSmXVTj1MKeoSAkOXaFjXHmMbRWyM0hg+/d/4BkiF7/psP/zb
dqv0faHXrnJ0c6HwbG0IQ1OUzZ3psbcUXKa8f3ok6JjVnZsroged3eMGX+sQ5NAK
7xqMzpPpi3iRd8VLAKN58nVSaEJpn8xiXDbHhcXZmoWk9QSBOZVkwFul6MtpL1jF
ExmLs+4OcRKyo8GLIoC4u850+XWe2RqX54JMS+gjlo52HSEx7VPMAYtu6bHsxPlc
6g9u3KBFv+p9DW6hLnFC7cXYCSofj35rEvVClyMhmw/RZA7P6XkkVmlLX7Hb//Kq
OOjGIN51qRnql6Sey8CZgbs6IHcua0tTwUqWmO8v3XqQkNKAP32fLAYvGqlarJ35
4bvnDxfHUR9IVv4IIqXH2BkxxqBSC5LgAg7AFTYSlQHtK8qmest8tfBMkz3k3hG4
qt6qXgIh19p11PnPMGzVTt1uiuiFqSW18GxFfD1CjBy7eAtmJzv408iAcQ0jqi/p
jWam0dXt51xBi1pUO9x0SlgwswqdQJ3XyWVVx6sPVvvK4htKny5hplxObDf+lGvC
Di7cP0YrZgT1F7Hp83aQ+JErur7RM+va+3+4ULgDc8VUhT2ljMxxWEHy6qwYtfuX
ACfQqaFCJ8BjHsFCXrZeqwH/AIsrcQe4/pKxCFXDIKJYb57wfXSnvGZgGs/rFOEW
8RLs1K/NnbdAlXqOVbpJGci6WIHV2Mc0mX9EfbDnYIlJihol4P5gl665j7FgpZ4d
jnqE6GZqgpu0B4hYLOvpnruYtuXr2wZ0vGrmWfee+7kkd5ZGYbgXrkIWi2cbdoMP
a7YIa3RH5UCun1LmUnvUPfWomZp0k61olJwa3Dyl4eMeKduXdtbh+e73oCQpbeX0
VONlP7cfv6kLZC7+HmXcfbJnulARbmlWxMspo+I8/jBHa/+Iwqmop5k6GjO1iyxu
BNXkkzaffK20yT19FNAFU/WGoUzsV7dLpgmqPFMJskAlHlGDaiJhsvXoee1UyDy5
zJaCJVhyyV9ZGYoK4FS3bvchkr2IfrFNtXj4vlfuPoJmbkouo98563ofTygi0yu9
gxAeHAESS+xhlXuU+uvaT+lFF2cE5c8g7GiAprY8Mv2xGwIJfKZoqSjkZ08fvbZu
T9p6DOnd+fZnwUwyZKPRRJTqtWbhgW5vRAam94HMX9QlvUNz0O6AuaHoli4hUlfg
0xhh7lUCmgd1UbajBtf8l4x/Ar2wpENFBUP4aVCDYvFd6hG+eZ8dIfzTwyAb1UX0
i+Ws7Nm0bfVHvMzolNlWPW4EYnnqvcNSiw6dDeb7MWw+jhhLVWXH2Z7rAoNa9NDo
o/Nz+0OL4HPaSF/gjoVVVv8ZWZCxrZWyDKZrlzLUaDcX4kvYEFYktLtx9uf9oF4x
ZSzpyj8aiEOA4xUqIbC1KEnvjUcJiMisP7awp5k0555WSUr6SyQ/gKCayys8N5wH
EKYMUIwewhT8TlWO8sTOSltAH0WKfmpkbc3DGQb//1oDYzzY+8lX8vENEXDp0ve2
r+6VMbRK6YC5m4mA/I0EcTuWCfZCdP7JFn9SXW2B5TNKHmhbHwXh8GpRaWetew/1
k9MwikqvbLD+okxma33QKaLZBcI93LlVSkSepUMECkRSWaabNOb/TR6VLLkpAyge
DnLssnmeY9dZnsMRwTsu9Ld0m4ELKmnx2dxSihEOcmVgXvxXmIWgZy5gZgC6E9rS
KkB+G8L2xIZ0y1BP8Eyu6CwnHLLFDlJetJZMY/rg1W04IBd1UC/xYBlldWnawsBj
X9r4qa7iPFJuABqdXeE2pdvh97NED+Vvy17eFg8NDrcRItHXXG8zBAxvCGqdqf+A
51G1ruNQR+9/CV3Cc2+GDbZ0qNWVxEtgY/nU5La3oiSyGZmShrr8jtAQU3Hpd0k9
rb9Qc4Ec5hx9OIl7ha1zw1rQdWEdboNbPm81fbHdjUZZoYmTq0N3xdZJMwiWmx3K
TCAXwj0kRJ+jqjE9wYnQlajuT+/MzGux/Xzc+pLz972FLIVAOUiH/xCBj5/PZRBO
Hp5ii90scphvEUIcdTpayDOSXX6XUPXMB3hM51iL007cpsjDvxAwz41D7I6jme6Q
7UVp2JAMCN0Ob4DEQwKoU8R31+OwC5uYpmCvqqCWUtx3DPkEnAC/dCkR9OvwCbO2
M+/rxqIhGaaX378Q50F7LosEozOMvvFDPpZl4YjrhHQ5DKUqTuEanFXD0Uw91Gjs
dYjf4Tvs3DXv0pFnhI4l4YOOB058QWkJ2X1i20SdVl2Ia/91EN8Jw7IYCzs9XxuX
DO/7PeWNL0EZxGNnmFJpfMe8TMOQzEwcjY81u3Fu7aStRRA0zVfSJk/Ep3pFIBYM
QnXLvAQLXKoEr2/soj/2uClgiCio2HRtQlX56j+a24xBojaNULbGNlGOgVvmSni2
oqMRO1JDj2Snr69KRk1iF8XomBX61mMwp8OfhSSslVCJaG6kdFeorzvv1I5u8U10
5MT5TnP7278D3+yeGXSrLjPzzcNmutlJsUgmfkF3X3recJc+oHOrm00sruzunk9F
B9Ma54eZlBzIni1BlK2cDm5/pjYnPT3nm4Zsx4qakPFWHUMb6NthOHIz+yMXIwDg
4+pXaTSTw9W6TmEdknJxrPv/ds1L2XcT8RZl9jOaMdL06voPz+Ylpy9PYqBGZGqe
7HeiFWDpMZEGruoutEAurCa1wOjumTnqSNdNEM7mdJFB4nnE1w6i+ul0RwaUjnu4
xOtg07m7z7gYiwYwk9UlcEy61SWMWVXgp8YX5/k9yiN4c7bAQeP001NBTJiYy9QW
QXId3lWsdKg0RoSFmXnzv0ZDotuB31HX1mqldM/O/kUUXjENQSskoVEjKs8AapqO
GZSKQ4VqIf9rPA0WTEz9vBk8lRHASQhEMX2wmpIol2oHPsAN4ZIWOkq1XZMkEB3j
X+zA8pPkUalTNFAR2cBZiRWQ+h5dnsZV4xHgyE6Er9e+9irVq+ytoNouFUCPeamC
2mBCUSj/xeaL8WEs3nQLbKjc4gZRGv+yq+GccsNgPGj1eEYi0Qerb26jsx57Xfz8
SsOHCEg4vN9PRcaWmLfDe4PWqyC2HPend+CoXluwbmF6uarUgsO1SGpNAktvvP7A
m3Ti8txTIoouCvXpfGotwZ/voOKr06dzjR4zo51LdzOxMYEAk2xsDCbcyyDhU5M5
cDjulIT8MpRLYcAB7E1oXgpaATe4W+Ww4pkCgZvJsPOm9FREU4+8Wf3Yd7z/DWQn
w4g4jlCPZKNgOv0D6FL47nGY5aftgaUcbH2PqAEO6G8apSPKDSdeOv6U7T++QUJJ
tJ5BGJtbowBt/ChcxV9fY5EYCevvWH+hCln5/FnswZd0F9svkL9ozomfTL+8u/2R
R218gpn9p8t2MXhyxQdCq2tf7zPy5JQCr40CnX3dGpiEgl4G43AaZ0dIUwPr9zi+
UBYk69pw64OhEuPEsOb23PvYQ7Ripewfs5DoathlvtTTeRLhDhabARYJMrNs5n2i
y1M9Q8AoUWOjy3q4l5GNMJouqYob4fm4u80ZpIE9Ac0CrJZIArYC3WFGiHItpj9h
zBE6667Q4Ma+bKaBa2k3MTMpo0qVJIzT3gZ2/bqTisONq7SV7dIKo3fAWmLsEpHX
u+OiomZJ8Y91gNhyqEwTYq2aSB6O7iakjQeOP5Nxc9ma24x3JKyoTUqByRCsFmCq
8v5B2yIo1/ojXpV2zWxJthz0j9G8nnm757Vyw80QfAshzZHbEuV90CYbwU5vnMTJ
As8SuT+9hDJhFpGUglNzIYY4JMylrLnq/JonFYRkYul4DcFgm1DvpasHZHJ42DIt
BGMyVakPzKN2bzmb1lB8fgpV3dAQ84Jt7l5LhwqhyizflrkXz+MbLcqliZJvxpFz
oEsbBFsm4EWpFsYJqIEVl+lX/RHiyTjDDO3obQZQ4jLzMceQtd0Tg1cFrMTdyOI+
KCoYQ26k3ISlXUTHxq9xCJ/qO2yZi/BEiBpru2bFDwLhuKQIp7Lf/Yb9hiYAuRy+
M3Byvh51pQwlo1cULBQE2ZhYlnN638ISYhXsDY73NLk9c0FdFl7zcNdk0d1Ftc40
0RGhOoHrjurElWqtDoQJxMut1OTh9qW86SEOs9jicYevWsjsGWhqXsKH84JqbYCc
ZUcjKXou7U8gzc3/gMjS5PTlUY9/KPwC8y0T6cdZznkeuXVIVDOXpIFEid4SmXXq
Fhwqhsc6b4nRzvPEiaJ263LLfnej6VvMiN2SiQazgjOLEMAp/SFnm0Co71+2U4a9
1vu89r9STdtlcCm98s0g7pmxChh97o9PsYmUp8uOninKqRfG2xp5wzjGKyD/vE+P
pvS1yFxWgmfBIclV/G1dh6W7u3xNH1kiyxIwp+3zDw/NJ3MwRH56uZB6lE6d3Je9
H6C6aTobfGs1rKGaBBjTnd0MmFfiPoOIKpp1brMoKvgZo60NOJVBZwEj+9YhS/VD
/IxJUqgPLkZJzxc146pvzEEGCHq958uxpujHeYxHPmq6idbCTa/98fP7gWpf8SBD
f4itKNjWnMWCu4qdK7sTMVXnTzJgywOOKL2LScDY+agU+6I85gPj++/SJEfLDOQn
h0rHXWOdzBErCPDEEROmOvTLdj3Pj7AhCxTRJoS0zCn5X/91rs9ZM1qL/VEWg85Q
9dJwzSzd5o7FJAVB604MBA6CInlq5kdB4AsEBDXvpwL6pJbnG7O+brbIwFgjp4XQ
yanahPz2gzEPSmUjtYQjKQVO0zoySxMs/ydEWv1/grEvsoEH4S/G0hmx00sFfyGL
L1fQ6fW+TZShnTH7iKqamgwyBSE5ayTaF4slL2csVXvZG/kNU+QcOww2Q/y5GR/X
SlrRlpuSnEko2alau+GzdGi9bNVXpNS0jwHMeuddSyPzOb1Xc5BOGLdm4DaNReoD
NdNwk+7SN+qpeusUp1xcCHXg1uJz6t6kxvv+szYXkWrSbQaYkoU0ah9WTA1DVapD
CSlLlvTFF4UZ9Rxoz1GwdZkuG33Ed20RsQWLUu7oIL+b+eElPlWKLrdReeViqFkh
JNwifJT7VBiIbGq5jgBJrIOk2WGTr82zKb71E4h/1tZovj5AhnfW87IjR+RQYtI9
DxxBOVndNh2BpWe5HxpkvxdIIdAnxL0PBhLmO9ys8Ph4RWbcenZi8Keb2a/A09Wn
yEOc/zs/gQfPkhsD46PGm5Oxs4uxywYXh4VmKXcksTmp97JfV2chdgW71tTSYcf6
gHYfNMYxrrtKBzMLrtPzE/lBuNy1cdbAPjLhu4iBhtsSHvVWIcnZNrsxcIifW9PS
uOD7ZZIyeIjxELKtsUvVesEx+rYBmtT9Vwru/0OP7Z/Hq5Oaqg14R0R7/YhaRWTy
qa8t69qd0dQvAAKAJ7XpwsqWK0xksDXMeuA/Y/HUpEBog4SydHtvFmc+nHg+PHAs
aEfarohFItF4pf0uI9RIC/bCrdgW7m0JqtGmdWW3iEFS69WKKNhnfp8HREoycABj
0Aaw+Zm4oNBgif2nfefcBLiRhiE9QDNkXZC6hOxgWQZSxJRmchPvydkR0FWxOWgT
cYM8ZrfJD6CbS54jdKpiPTD9J98qCTpmfFxdEHj8hiLBrzFc+Y3TYvodFvku74IN
WM6jB+GgW5M/isshzDYFwhH6gvXgMYEhdthvkaBoKpciw/Da49M623iIevjxkCsK
Oe+lgdOnDtNRWYEKQRbGVkNceOazHkLeUddg6MBO8tPE0vfEZUtH1aNpBD6eSOuC
ZdSqTRUALarEOcbEfQC2UtHONs00puWFei73xdb7Df7M2uUi11r/e2qg9SNhJZGq
NjcasfK6rKiN6fenh9s8iIzwFcWPqkgYpefRWi0E3xQyIJDO1uKHTgmAIhMc2GVj
vakDG83TlnX8YVE8lJ3FAM/1nJBFUHu2Fw1SD5/zxgz/Xfm1Stx2ysq5UkYne15r
zNFfe4cPslBmpqtydXgAzVBOpiXNoI9+CkxqGviBLIAkriI/W1CjD7ROCrQnfQCQ
Y/w6uKiZuRyjf5DZMb6DVZ+9C09lQQ0JNrl3WRiAD/PyFwf7f2hae2nDWf0Q4UTa
Mctv0f/bnOeLstuB5+klA4imjUrd8h3qLREjeuDM0PXGtElatzVUEhemzIrDaNiO
orP1YobLrxQ7YymrTx/nPqp7B0acya/Prmgo1YVoXIXLDp9yl/D6l1GiziwMIlIu
gR3evDkpzIG//SdM7gg4K+sw1THHjPR5BDWqdgXNVUF+oF3WvvC2VzRPbMXNoZG6
ezw/HxREMpCmznsTI98c6zztPutauOFiF3N+N+QrNJswmFUTIKPthzcGLNaFX2rZ
yt3rEX+EOENdMK8/Z9qBVzJaCXZE67EMFldCBu9cS/RKiIvvXAicyj0MFXrJU7/j
8mg7HtaFdS9n2VBpVKDMGiyp81EpuDTnQIpEKLfj3gVYn958jP+DSwzcW3/kpg2C
Fkvt6FURKH6Yj7tRqQq3jquJ35dMA0AtRZ1rb6W2JnmkwSw2XdMrmjAX1UzFBHeH
kPd9Fi9E0e/9UxeodhOlAzl/1elWglYT4KeOCTCDZgRgOGyZThiXeMTeVmK6EN6b
dBPa4RZJz9EPyOiNXaSTCTBQ8qQ87shR5TeXG+iDVJTuktL77rap3v48B2NQOczF
aMltrM5A11Tm2yyfpfUhc9yUeRQvuqUAyEqlxN0oDpUQWDPJoGDl2hs5wBp7K6Dt
XOcC4ejCQJsLfwo3ju7dDWBm46KWQf3OHJqsnlWEfG+QRMGGmFxVBTltI17UN4d3
KqOUM4YyNg7B58c2/2UBiOvmWGIApuv7I9OogGfQNDUPhlNN5csYAAXimzA+M4J/
2s9gO0HU3siSAGOXKh8q0Dpm4vo82KuNGogpugmaqy2eygEqKKsztJfEdD381PUj
THrVK14S94TdTgELE6U7FCZyGb4W/0knaomynDO55wyaPN+loK8PecY1FfFOvAci
p9EQhFrwcs/8zAlJ/LnytnHyNk2bU7NHT7GjIYh9tCfGVB80exNzOaIPs+C5DqZ0
2F7tQn7CFSC003jV34IL/bNcOof0U04FIsfXo2subkRhQh/XJvyjanvQzKWA14Gw
+qbH8JUEzvrvdG6a6dYBIiHCD1EwmndlyV2Y39oj6GEYzaVwcnNb70EbsQ4mh544
yESvUVjR1m9Kr2uym8ME9x5Jce62TxiTeWzM/TyRCDRWq86M5ho/RtYYfQDsXbuv
s7/9iez61SvgAAGLfrM/ihUDt2sakaU5ov/oKPwDBfHOBcWNr6SXbodyT8skjNji
/ZYoT0BWn7+EPeIUQAXZ38YvdnNh+jeUxnRPCTnabc7pQZwynJxM1Egf0tPD0eaH
H/5aeIXAF+EO970UVVbQNunp01s+1FCA/gjZYiPoOHAMilDr3hdVL6W33B4dgU4Z
7tq3rED1B8vHENF0V2n3Wf3rRsnX8E26Mljm94Ed5V++b9skISCYv2kPQto83qI2
Ug4IZagUU9dK7bzmwaVDkc/vtV+jl771+E1eTSTpdc+eH0ooVp3TLDzJeM3RCNa3
klAoC1hWuxgnduSlT/ZMatDsrNfZPwBWpYoR+G/14qG9gh80Z0jIyylbxJUVCtMB
TMplRz0qnZEbRMOcVGHnL/9EIJp61RVYYRRR3Z1Pge27WP5GxVdc8JeDe8dEikTw
el6dom39Hj5Wkf1FE2vYNXI5/JdUB4icJT2jO2te/dVliwVRZL4u755MTsQ8SL7C
VXxYVN243UfpRGLM6da1XAxRt/s9t2Dm7VpP28jbOLoe3x21S7fNQBRv2vrvqY1A
phJDXl1/CoUtMrwEfHOuQ1yfuZbiEsgEtncLPYYpRNpqH4LKC6JmNzzqNhJgJFoS
hxppwrV04LvtY7AqbJF/WucgpgCnRdIgGZ1WoFV0h9CUrN1rzlcRcBIWrVfSwnTl
HyHs8HbxPZPSZ9vSXUfoTMUkDQcZdur0ZgU+RM0ff6FAXjUPWVS6MR0JMpOcBxp6
0Mg5PUJ4DKXFEoeZ22eicf1Xn5B6yK2l9Dcxb0wU9MqD0AbcFoikc4Kci7g+pbMW
Pqbf7uz9Xvl0dkHKW52hiyOCyD4ppmXM+Ppe6LFkLSuWC+ksEX2NIJHv7ZFNUH9r
sFQiemTawTwuJY5Cmj2CtJIfKFDHUTgsdtY+Qkd2/payYsrdEHFMQ0WgjW4G2sFU
Ky8Yo9WpyHr6xGH6HhVIWxLJ1gBB3AO3zn65VmIbRMxWJ2SCiQR8qal/p7cBrw23
iZmF40/PK62LKhnD50LT55RNnPH49IKVl2+OQPE+PN/tgulcMZSTLKXN1WE7t2Rt
7CeAdSRpbMp0SI6xCCH8lK2UKzkzHPCzDxo/GOvzGKUkNl9f9WjKpWU6RWq6kBOy
P0gbR0vL9mGvmw/w+ap+zx00v8Mwzv7zNG9SYWA9tzet8px4gIK2oDCSgbp87peE
/vp4j/rSXnvAHJOyIykwaABEnVBJzwhTVTfOktZnsg44V1PSTCwySor/Ix7Vtr8W
LW7A1et2qtXkp4igkSI7cJkwY0SCkhcXh9LO/04dOgneGjKkw7rDb7b2lpwOB+d9
ahdCa4WbRExR2vu9B8UuY+v8OZWzUCbdu0SrlEG3KNJ51yAjDGXydRsBzGzMPSww
ld52xm8W2NMdb0wixhmATv2OeQWWI4qgvljTvYL+pdAXVrYJt3kmTBUhAwkH2zg4
WNKeLaa8HasyuSUi5Aixxf3MoElzJoevJBmYKfuyXwwPhir35qJS7vQ5hUlxaeEg
K/wH45iwvH3gLK9+b6QUlH+Y7stVKcmxkcu855LonxUw2rvPz3TX+tOh34eOey85
hHFSZ6C0G+1kVjQFkpXfDLiRcOFNtuktDfIO5/8d+xQnjaXPCDsqNuBfurr1K3oq
jZ7xsmMdhebl9gB+e+RQc2Xr0XJiub3hHlCrefZSw7NEMFsqpCkbWTiksznhQS8+
mTnWxmTbIBhR+Omnx6UQ9p66US3hk5b+UQvGG0Dq/RKOUzFqHSgzd2bbStwxTDMl
wR3G0qmcpt/7mHSDD8bclpsJ/xkGtfPkdlBT0L5jHsCnCSnM9NnPnJufHzFKU59b
Hpd8+axIQt2s70n2VeHIm2xk/i+3h7IUYLtcZwD+KMjb0G/3kFWRbYa618uFd+Hv
8/DYIM4LZzDBlJQlL7dXnqCyNZ7axindSeGbtP0Kc27OTO68BS84tF/nXxXNx6/T
owzhDVUWFVz37btUjBiXqSBRV2i4dwIa90ebfpKo3bSWsuXF+OvxoTsTUZVWR0U5
r0GR+W1AJmCx/HSY/sFcfouVQ/wZ6d6IMMioA1rcFvpzx8eTuoqsPTU6yZ+yCNUa
d4x41Vvwm+tSE6TBc2es5wrBm6Hta1BnbiTiPtpzbJR1pdgfCMrLSxsW449hJiWO
EMDiTSkL0nyF1fCuEwsNm3eIH8PZwSyi2nD+lDJ2V7pU/QOWEOY+nGgJR+n0OK3r
cJFih7fmS1CH+Z2f18uNvuAo4znaEzp1SOWAvaDdWZjDm7WYOFuFFcAP6bdfNq5M
wn9cNEoDhgmbvIKEGY9sGaLRkBgiK06smgFVcupD2CIyERdaGsj9SexzIknX6CNO
KrFhD02gZPMOyQGO8AcAv+TPzA8CvCQfTYzyJKG4AX2Buc7G4PUkjd0Hc6TRfLAa
aKPf0gCTZIjGKruC19bKafHZwSHq3jpHtDaZx7UWfYgbc1SrGe8zzou0LIb9xg2B
y/8q5x6oX4GTKvLJJUqQtm21BuLGfP7E9xM6RQJBdNFOd2pBU2szxBMfRrZzustT
BWUlBYT16TkFOI+Cov4aQ3qDnmyMfVoXZro2f89nJW7PpLXgSpEfepAGaKj4C15V
mlq92TStuNPe9eaXeqw6HZworyMa71CjocwFkijoxEaghZe7T3P+5BKllAfVuJHu
EcSHU5EMjmJuzqn5ZzpfDJuxERR/aqvlekc0V/xmWAmuk5bbDdFiC6fiQtkglI7m
Yllq48ADV/Vc70KzX967mVqUgkdZm/6qQbSnpfV/w+dHyf95HwFQ9V6K8ersiT5A
pQw/lmMgkiUHFWs/QKmjLPQh1TMzdqIbOUJARRG/vgVn3+M0Xpwi0fPKaT9g3pHx
8thimiutNqu4HEF0XnBdd+8iVKxgxHu/M23zNwvs5mDtsmnRQRMToPEiqS1d5hQm
htoyxwPRZ4iynh16xkUn+qYtXYnIIFhIhz9Lf3UdZJSy8PysDZhaTyuCYGKN+cXY
5lYLACiTnLDA0dQ1XnOCVJtvOgEVZJIdb7wRH2UmQemBRcq3zARQ0ZjPJmQZ+UQM
iRFw2BhWx30DzxCJBRanoWg0amwGeZPKfRyYpkanrTQxmSxBD4qJzPNmZyWccawy
fXUBkbAUjoFthrMhFqj4aFPm0OfRqQ6MH6SOJzfe26rP+3Ts2NhSqeR2myg+w7CH
hsRIeYjpEIuLNUAZh2znSEilHLoCKPNd82GlPQgpIc83lyvZ4Gy8VGBxnIyHJgj0
m7qP9RfGNMEHmITHvm6KmFhBIH2OtkKqFSJxAF5UDwY3MXslUeiLk7wwMWQPVvCo
rg8v1Rzx/uLWF1CGRZ7d1K3VCQODcUlQKZocOLBm9pdgo9tbKeu4uxDb3IaEnbCw
ygDcQN2s/E8mXwzHpiX0Eu43XwpQJ1nSuctRUYm4xQdCoMN0ZgNRfQVBLzMyR2vG
ktY6gmDF6LnztoTRLi5uJz9HDnETr+hwGAox4jU3lRtN6OfQvPHlIjJqeNjRApxX
A/W+eLYdcIYVdK1XTQ/KZMmKWXE/f1r7re4Vk/3Qu6CGRJWZX6/+oRkjDeAxR9Oa
A818pfiVFuKz7I2Mh8UNX1PggTLX+RuQjLsI7B5s+tJs9YQwt+L46+CXxrFM4tQk
/brszBZY29caA7+LpUdgzGEuVAYDzhM6u1Cp7wk+F8CS3X0/SrDHROnm8kYCIOe9
XXr9/QHcKS4Qd5VpHSrCXetVXvh0E0fyRhxFCgXeeRbqL9N6sOl/owyCYG4YdwMB
0q0HvXj0TdoFXn7JNwAJorq5UmrXsYugAnbyrV9WBZUxc94J87Oqv36bWLcctmmi
riHKz0VbSBhBYc2mhWjkZP+5YJ7gRKRZ90DkEKr8j8o2ur1BiJWfYziKrHL8x1QY
MJ2Uj10fM5tcknQ1lxrlTvfiUOHwbg7fM+xhxYQinUqrIKXBYYzyre5ZrOZvzzyp
RlmV31GWgOIRFZ4GIIRZfP0FJkR/93J71AP6wQR3EYH5aRkMEz6+fumNO1dWQRif
EACFzx+V5cNL0QphWDgAIkxdCadMxRhT6YeIECNzXDhPEJHP/x8sVnMCEeBqoqJS
EGiXsGGWOc4OwYvGRS9zY/tVd1t9mLDoS9IcOlN7lN/yQ7wxbxPLTNk3sYcHR2Eo
WWZMoEtK9T+GAn/xTDLTws9p6D+7y837dh4fC98Vj7dgE5ZU/DSRt7YK3b58iytQ
TZWvuAKjiCIyb8KQcRWsxk+/YPTa4eHb4ohHh14GAGCvFMM5gw/uR9MsU7CSZ93s
Cc3k/xyMOXkhOfUep6CE8dlXXvPGJR5MJTaVY2+SufA+UHnrHEZP7bwFe6qaDjqR
+ZT5rz3zvNpiAyQ05/wXd0L21fnRlslhhd90Chaoam7IHgRm2TqvWtYC1D3YXYFb
agCUKMgDxD26USmbwvL1kgKRymkrK5WHYOU5hNmegx8AkU4O2TUJtb+Pu5rrCeiX
iOZ2Yc/d+rN3j+S/UG/1uQqddiYySkGwC8r+Cb7m3vwWy2tQDIUSsgJe5lIrJSOY
Yfyo9nE8H21qKyb3TiywH/euEWiXXEopXd6N2EPRhVEu3Bk/NrXT++7o9SgPtipu
Lc4ZpeBRAbxwjO177q9VgkELaPH25QZ4LeUl/kgUqW4W75C1zriME0ei2V2iqMZE
Bdt2kdg1AZjK2DmUhEz9Gm37FIuy3lMZAVMbrcSb+dY3ReobZpjK1tWJ3bFTdQ+y
lw2iP2WVg7WwTtO/rML2g+Nlyc1Il8mFBZPWzcrNpELjc+XnwKBgfk6t0wnFwLsQ
Ca8iEc+guYrapaKpUBoEjPwT/VRtQAiNg9FXCvyQl90ifzy6SIEQgOLZCNH3S4a5
VwXLl5yHEdFvqlAc4UyoB1dIVnvMpbZiRCRgVlqrCDXVoG1wgEv+YZMlJlLAAzJz
Ufhds1hATZN5ZnQOTppryxHC5Y5fgKbIqzK1H2x56fO0D9XxbuOcwwWl8mNPQoqo
6o4mN+lP45RrqF8W60VmP2l9O9Vu1K9SRDCr9scJGvHFPOVOLt3YL8c9++mdfUTP
uzokA6R8tqUmjORpAAlQxohY20fDC/ycqqwPfNyAXhr5wCWdlQLWEXLH6HytFNNO
fQomQdYfXmPzoOy+z1H9ohsBtuOOKD0WIG8c/d1jcCgl5y/n5Gb2FkdjGfxMdQYH
0TB7345cR/vU6TuhQkcXz0BbldWUqKpK1ADJQRfOJnEumKECzjT3v9D+p1BSOVnD
mNb44sSakrLeIn8Ca8gP2XfWgeIcwzBqmkNvd013naOOhJNO1/aJd56jfQgxlftu
4M6ngk+9HqHJezuwSmulHW8hBGJmKuNhloS0XAU5ieMSriLDzras54FJYQHfx5Hd
6j/SFCDxhTRSIAjarBVZX6ANB8FXL4XM2kugm150ebZyodROXDWVM6SCET/mV0Qg
YOLQr8hX0nLSosr4c5xQPOyYnlVcvf+hdyI5r9Ak4PcC1MQsP7MDIA2vBoDI1t8g
qdR0+hfsagySsqntaZZcbiC4oroUW0RzSnQwq/xdHwSNnwnW9GIPX61Mgr6wRRLU
iwP9DWqZR0VotjETLtt/j8HVvNo6sUksXEwzIVEw5PLS74RZnGAZWpASHbMHTSAp
r6uLA8YUhZNdsP2f6rahAV+VzhieRfxKnTU5mSCf3risC0M3rGEC/hhn8ez1nFr/
Ab+/2M0D3oV5JIXFJA8+u/oJKVOMLN+bJJXjLkv/PRVOtx5jsv6acEIvodkIfZ1C
QkbL9NY+d8KSr96qKdxLjSEE5dyvf6NFVTzeLec0MdDSxfCbiwJxZ+UyKF3u8gRQ
6E9axPr9HytAKVKL0Jdw1PoDEJkSFh+h5R9QWhQy8cu+KJ6D8MEKlrjeC/16Cmyj
pTwtryxynEczqP4xqNCuD/2h51csfsuyai/wUO7VxFFAoBBCIBUsdYopQ1GyrY5u
2VWnQvx/NWPvGIA5gxE9AdOaiWcXbqfbrNF5J4R5GJshk/Es9kLjj0ErEeYsXSTb
zZF+/ujgNSLO1qbHIqv8QhhcAIKZsbgSvW4R9lJXt2oatIcfJV7JsJ8cqXr6oLP1
zB71KloIfRj2Jgcjy56nQ11JYuh42acPHARKczXxDeRL2lM8iv2kdgw5XiDPPCm3
zuyuBc8rrRoJsbtKuoVB/C6aCfdm/NuLwNr1AZnIwBndKcFJpMY7DPcoG8WlOZSM
jzkEetue7yttCIT+M254mM5F/HiUbNykQn3xMMe83b+AD2ZR3MhebT4e+3WD8+D0
9WhLW3nY4Uo7av5FOG/zgK7n3UHzPe9kOApkdEOZWDu18CikI9uIeAd2jhVjgaVd
zhqwlfmHpSqX4VYBz9Vmu9U+tWlswIwYttsp9Bkl/sHWMPSgsiD5f3yeL5dgZRQu
9Grawy9S6wYquI9SIEGSLPyJ1kBGg2f0j+vSok5lvO9KQCP/rML1SsubmhCVstUS
MJ+g8e2ZhvW0zRmOUmWlucu/HVsPKrNGPQ9wAtZE8z4U9A47FAFcgs4HFBYcPvUv
Ne4RPk0qNJUb1rolY8QWLY/Xmw/BuqKUdoMd1e7BfY5TL2i+XEhDXAD66K/x4B0f
7TbiVn5qVIz81jycQVJGET1SiWPOIE+igC1iyOH0AfI/NQxR/7tj0MaBD8oe1OGr
SUwU/+GzCN6Re+J+3RQX8l2pjN5Sw0ktyAGZ8GicAtJPsAy6Y9HOHIh/WzxvGbmf
JtRmNhpjt22QueBsXBNb6/cEYY1Auk6vuumyjO9Wn4oZqM5oVj5s3IuoLrSbQV05
EeVMiiqONMNCbeuIkIRbSHbMiKXj5eJjYV7yjQsHHSbTwGUm58F4RORVP+UQz2ic
p2vmQ9Bsw+wIj7c3rHs9srMFQ7jH12KbuBl70IYJhwSAk3S+lY+EQIaxQDoW0Xex
Ay160z0XwvdCndEXOV5yr7CdSF9yMsHIFeUVtH/x6QisrZNEc3Mcu0oXtQiqsxtK
dL5ZylFrcee7075r9Sp06uTQViDBCsNFrKOtGXURBjn4qJu6gWkOcUK2quX2tnNo
B3nJ61wfWMafeDdvwSRw1iqGyHDQz5DBcl3Yg/UW2SigwchHykt0kmwDFhOp+nF5
MUiYUoBKJnz2dVHd60XO++DsOIrGGwiSZjPiT5BiI0X0g9j0kxn1cFyVlkwKSrW1
P2/Mcb0uORqDkSZfixUmZ93yx4+NmxT7k+fhw8KDaLGPng9d726/Nz25G7CHZrXP
z4w9REcrU1EjkW+TxM+4vU7qlfwVQL4p3n8ZOLeLuzWb+16iSlKv6+0ukNDcv/em
zWEe5t7uPo6L8ZKOPWIkMN8zfH9WBZarW1dFL3EWYlFY5n2hpIWwEOh728XdfLrP
tWoJMMgv/P6mYeC3rc7y92FW+AbEMLwJXJZ/7WKpMsLqcO3BtQTH5XKUOalhNql3
8spTZZNpM5A4qRhtDWCbxRWDQWB07TVLyj1/eQYgnycQw7dJ+J2yIo9DGuY1TSBm
/+ye4t3evo+ac8D1xcDJXE5BCkEytS4I1ojEX6souA+trQAIaY/uvfmvAznuqkNC
FZdW10peEOayPpPkNKN6wc3SxeXtEn53wBWIcHTSzO7GVz2ifjlhxvQ71TQ8QovX
2d7xYNBBk/hz9JMwyHmjoqcTCNKaW/TPYvKqb+oVqm4rWOePnpNAXf0gdGBSCCx/
HyIdyTUtJQM6sN//cmzdsPtablfGXCYzRYf2EEQwl9EC4d60MbfxfIr5E9Is6lF/
7i630HqNmNa62uiOUGbJngyVg3+AvQjBi3Nhc3F5cESzMMT4aGEZ5SOVrAh735vL
oy9KMqEVJFD3ciAdMxvLEKSHALs4cfIKC5i/AP4f7HlTdSgPaoD7tPdVkpe2UpTh
/TipBsVUNpk+syxsxkwcF4WcYdPk/hHe7x393lT6a4Bcw64qgH2KL5vajFLnDQE6
eQCqQ0VsRM3BHDDms30mLwKOI+ufBcV4oQPTsWkoO1o+71DhpnEj7DaZq3z/TnQm
2imJBEERSuFmbyZomEA5CNH5EXFoY6ghsvQYGGvs6wC5X7fknbyw89ObSMWjh+GF
/FK2b03LyKlYsC1XnP7t2iADyqG1923O9w50gE9m6JAlnqyxUqUqSJst8BYAE+dr
ceFXTPhuedPiEipgX7VKI2pQAhy717RSdlknWppQ6SIXwTerudk+vkExAomX2qsn
IZKX6sHOMUIQTAnfM5mdHWkHeyUmwCbg6iUnZlAcLal8JEuSYknhfi/8rQrkvDdp
/uMbfq4a+n+wdQMGeARki/BV6wo32xJ27imeb3bAxljSGrOYo9pqKbTtPdAcQ85+
K/C6fEdhR9oFhvGHvt06Y+Qcb9wwcr95zNynngCZ15BK5fbUZ5Kpr7S6nIAlBxh7
amOryUlZJxcPHKwV6+po7yEYJWEWrh7MTBNzqpUm9ZRXZpzABKp48Z67uV5MyT2R
/vqNOGIyJqjBSKSC9FNyXpik/B5zZx915IiEu8EUBlVIv2Jzsswb0brqaLN+e5/E
3pVc0gX5icjl+i0ixdtJnY6+sJP1yLRhNpPOkr8wOK0Nj9YIEZW99P9tkcVGutrO
N/R3ZlUYIFwKn44iZqeqm8ZiojrPs5aq0KCQ2WmmFERM3Iai5R+UyYrA21S2DVcS
Mc2ldvdUixxSsJwCWiuR3GsyiT5zqWhDIXfvW2eiCKbLzbpDLJcI7Rqf7a/UJwKl
8Ho77RZPFfPra/YQau92M96g9hIMK/Ds2ocqac0Nk48pgmwu6DtN2AhYObZ/3Qz6
K1wxsSOaRSi+eY9dt2KE7TiQOlwuZ1Tc4XIrB0UgCeE54wAsjPYpm7X/UjBU8baG
3XCPLePUeHDBcLHUnhxQmbzUZ2cOxy8sEVmkcwbgDQeQbQbeD5k/3eYkbefFAEvm
urLGwIdxEEM59hStNra7xrFwJ4d4aWx2TwyrJ0nwjGWT8pcsooHxtIq71JD9ZDkE
k/zC/CzDi9ezMSBXQOIOlO9/XoAozdbGuUQMY+GrXO9E+1x/2jh7OIIYW4iJDZ20
YgN6MjZrkGO46n54ZHti5/LhiEB/EqXy+CCDnDrbFuUd0NHHf4jRgh+z0jFPjAqg
L2+K0VsDZZ4RoWGirDjUMhi74+tPp2DjWgR3tcxFfMdLfc2+SHVDyzoRIYonVfrO
eSsb9xUG3DHNhef/3pmrIQl8X2XOW7we8+Xe2n1eBQZD4l8KvVUdfcyGEvgyoh95
BQ3vc9dNq0YKhb7f86EeU2XTR+iTa0+BV/XmnNObqsjAjRMrAWxqvP7sL5Ty1+++
qSdrIVpwe9EyEmOf3QgecWlLtm76hcmcwftjrIx8FlBIbKf/UC3t+sZDAZzfQpr1
/UIjWI5lRqxkBxvfYCpFSTL8d1Nb4T75hhoK6jHgrs5PFJFl0GMt0nExdTRTHzxS
UPYDr4YjTOQXDINdnsmso/f7Y7q+HyNayO0rGS6ZWyLrIClO5E155oDQdkAzE4xb
JdnTOgShbCVlToWdyJ5RAsE4GhIwN+LNSfNAWBNfxl01IZeo28r5VszCPTpQ2Nts
eTbfJ9Z8iiueXG9bpd0Lc2LocUOLDXlv/AHGFA/gM2CZcpWFEQnkpLVDO0WxXy8s
tSPd0v6WvKC4gYJ8zOHZNZSy4SOr5+0fCrmfa2Iy64jy3dh3Hib7sH89RHIugOuX
94Py0FqDWJCkuwlSPfwn5AC9NpZYT7vD3CRYcHbRCNVLdglz2FaOKaxjpwkBWRES
FyzILqqH4MSyRfzbhHd+tn/zM2dkLp5PyBFL+e5oiW8BCgjFTLAyo231UOrHjyvt
E0PTDuGRMMane+QeODcH868J1F7tjVCPFjkxgdy0IFfLi6U0E4ciLOFr7YMQ7mRM
UH9f+u+2JuMUzNb7ozXi2vg/TWNrBN60pVKM1szzCw+362Gsxou2P4O+psk3Z55h
o+KYJuRm1joT7jRZ/cN/9Y6GvPWi9yEwUeLz5PwjfD0ImnBszSlj2rFmBt67lDbP
ARY6G5V8hTOtMo7963jrh9+vPnUZgA1yZACGIVU6un2elD3+/ZiudbWasmUIQuEh
6eZY4tNFALhkWzhDWUcrwUbl07OvZjX7TXT5l76P8dqF7y/lD4aAXKbCb3BgnxkU
P3E+VnTi1ht+omZMLOlsRALNDY9I9alBiqlJJ/z2xf8qUkDdKLxtgSrZ/9uqM45S
5t/Okbt8HZQsQHuF6H8GAaAmkSvHJDn1ez+MAkzYq6AVJpqdy7wIdra7C9CJIpvu
NailxctBfGFnOP/8JlFvb2F7DY2iuojyDDErgNkjtLSWz+sICA0Al85XHCGN2r1U
uHRZh9jX5lHuuaEz8Yi3/hx02YYBOqNfp3own6iLHZ9TelXZhVU4SOQ9VTb07hKC
lBReZlHGfRnb/MMaQeUq2YQApq02Z/GjYWYM7cJBaRjYPBk/uX6H7UAz92O6L+9H
LQy9UOEAJEip9GQYfJ8JJkV2so2Oo17dBbd+HLKPUiAeYAZyprl6HkuzorCMvDjG
2gK2xZElPuELZAzMnvwK7Axfo210L+gvuToOhTn9cb8O6DE+KdW489G7UwgM9VR2
87F+bQAmwEfOD5HOx/XhFNawMW/QTezRKgvgbwmP97ZlbVSPaxiLyXCptvxh0oZE
Hic1A8MEBiJRxVgBy2OTNLcLBv8LJqPpW+xXgY/0AmfU9wkHSruktTrPCgOndfbV
nNFvXrJnGZ9/mQiuAtogmHtclo3ZtPdxEs9/zSp95yAJNxcK86JBOymjgHwVTGQ+
8yC+pwAST69aRlbQOx7bEo6O5FVoNK7/L5yej9XIO9l30W2SdTGM9va93r0PSkCK
7YcLTmvOfwcQjptbmy1Q4YoNpD7otWKZFxQ1Boe0G57wo2iW5DSOyhAmpUMtFPwU
2FauEG0Nwal9J2OX57UFaOoXjbIrmLbE59sioW83TnV7Y1eiYk246xnqN6Xz2z/A
sTZpKyeSCVdBBiXTeV1FP2vpxOijU4V6+pjXVWh28IW67FPy6CJdJdoG8RpNL2hr
hKGWqVp6xnyg4/9KwsFx7sBPLiCNSk9UvA32b5+iQgb8VPKTXsJxHm55/XtMc3uB
CHnO5vjpyz1S/9wBaJLEby/tXgXIeSHLQ9tq6YfZKxqClNJEcalbMjLI3wbN5i04
5obsEcW6+YD8Yj7egIZpvOy6aykn6/J3j5Gcl4AFkik8OE6Gak5jUfXaS2ugW4ON
SQ2yYRvKQxoP2ISZ0RQQDNuvJpAFYWV+U2hLwJjd7GB76/XxSl+IKOxtXbCFJilz
BGM5iwZNwpjhuv10OOfSMiUphDi2OOz/+apUXqElSmCd5at1f+gH3ViapoGbEigu
maSVoIragiVU+Un2XxIIGWOreOeVYbrzOjBkw8iQfuFzyGnFFeS1n/4WLF+bhiIJ
azu8Idg7vRCBxxIsYLWBbn+hZnZhGnSXVyLY9/Y02644v7WBS9+Y1/tEOTcRmPNw
DK9ep/EACfdxQObTJbkmnAn2ScrrozpQ+W3Lw0dGzQPP8jgHgaqSBTZL/X8uvWHp
9dXsQtMKrMyRPdzzq5b60bGYr0ny7jfS4vyc+hEUl2gQtugdXLQ1XY+JDiFx+X+G
+9+jhA6vFMkFPT3THNTKvoGH8Ta4ilhYg5OXqx8rOPOoOYk74lYiYEMrhY/vS7Ig
vUKGTOD0Q7t6z3rAuRaNzj7vjrNpZ7UBmVm3r0Ubr7noSpqhIjPC17NZ45mARLl/
umgiw8JPHYnVo0vhqzLKdHVXhWBk5mHNZwqMyRJ1Mo0AX/ZxerDsISim6R9PXvlw
CMVLLndu/zinuQsvvHbfWIrG3AWYmvt9fL3VvQ1OrLZY+orx8ogpfL/ew6duLXXZ
CBWqlCtTCSTeyyocx5p2XmzZc0eJjcQIdZ3VSSo8BPE6gdwo9bcqDBxM4wmL9Jv0
Q8kLJ8GsMCDdfsvqUk6CcOnjhfGN9nzGEH1ubDqWIFuP+ZhP0Nb0UpJsVfTg8Veg
nILqvDg0G9bUR9bnMxPbNluLUPzW6l6RtLLBPs6PQFSod/LzavLye6cuGAfmP4k8
hFo5i84flie8xsgZ9GAN8w7leVeK8RJwf6AnkVknQMXDAvxsPcnaq+5qjmayxv4O
3WCVIa3XHwPpksbUWnRCo40FfPs41uu+fBQ4BHRgUKB7is0gyYVEf4kubB4kfVWu
ZeAj4atHuv8w6wCiAT5XZEJB/TT8aWuAUs1ggfRT+8F1f2G0slT3pL/kDUmapapE
tLklRDwqMFxu5oGOvih2c3qEJABpPx4vZVJAMPeBOnArxeziAnIfGoblN2sv6u/z
mcF0g/lH5P3BlZHaKvLnI1BjHavp3EUmqNn7jwCV5NhKV1VnZOItHlSsBLTMVjnX
ll9J3EobSNz3sq8N1cv7uLc13t2qfNuziIbajz4QxsemLCntsANbtr5GcZcnZb8K
cZCWFNK3PzUU9zAmYWZTH11BYFwlCIrjIR6XofDvWE4U2ETcC7bZ6Q/sJ5Jhk9KJ
QwP5aTH0IK9fxE02uuSIvv7fNwmE2ob4NJWR6D2QkKjAa1X+rHTuOLIqXW2/AkFM
SgGnUe2ro0/d6ASgH8geNkqg0HdM39fJJaKBMTeUoH0W2WZMfFkJDDIf0Vruiij9
Av02l2402gzSTU4w6NhMPoLtfb5LzqlGAW8+6HoEtnFnwc0+MFRDRrT2gAmtds4J
cLGhb5h8XlZ1IgDeSDUte6fxcuB5rhiG8AEoWlG3L9g1Rbs3STdoY5567ICt6M0c
sNYUhhTUoCOf/NPDcxXrNV5M4S2aCkrczly6w6raO+zCcNAYjTrIddr5ue8l1obJ
jM2qXjEGMaTgnLgslTE8wn5n9MNLKWuzODhZTgRcZ6n7PnMyqTVvo3PEdQC8Z9IE
V53ez41qYQXkwHCfFxPj7J2sDf78kO7RY71lCwFx+RJda2Oq4bB8u5IbX4ZTxVBO
eJS7UGn6vo4pJEKJGYtQP3cnuve6rhWiXkxsXzpQNtwhz2/o+d9jDWupb+UiuRqW
aJj4d/tkcORdESqom5VFiXP7z0dcS5m7MjjTb1liRvy50+yo6vycBED1b759Znfm
JeUwZO6ZyuD1f82dneFeQ/cg0HGRf9mBQ35ji53/6+6TVD5VJQesGw5GUmrer03Z
pzCdRv4HFsSUHMHHkOb6otC2Mly/jeFG7CUJF7+X91vulzRVRzbQWt+x9MCGzJ35
lROyx6JVmMm4zdvICFnwv9OXXnQFfeffddAxHJ35W5GOw8RlvZ27Zoa2tonJyn5L
+kozhDr8RQC0ccW3+vuGFng/J+CJD7rLz33u5gElNvK011AFnhjcIQMe/XCNwlrD
hnoTkpeV2VBUk3Ri97YO5FwP3SYGX6fOa/0HeaO/oi2kpzsovBrluCaVSGhJes50
SiLBL+6ULx+pKw+qcJzCvsHc+bou1iqYo+E36QDr+clccWwueLcTvrbJWuN9PtwY
uff6jO/r5yS8/DFW39m3ppJYBwAHsmCthLx37O0X9ruf5fpMa9PSXtJG33/VjPc5
oOCM8iPQOQIzqv570LLjTbuFvBozD+DTLoIHqaCGZqY9BPveujW0+OykAQyqDq8W
SAEEjeE1qZrU9DLdnAUMWOWs70Q1l9J8Zi7Lf9NsmfLGZfeGHftRpCz6osFbyxDN
E3xybjVkTPhVakCmCwZE9CRb0AhXM+5R4JhqonrkZUxdr0F/jp7FNXAMb4sUElvs
KpLbajCPNZdXgDtptjvUYJymsaA4rEabGAjTu8CDlIzqV44x89xNUQoxwMoZlqxR
7GSIBy0WYt0UK1gL3gMQNQzqnCOn3Hl4Tw0iWKSS1ulZTcao57ySUYIBIddpgm0v
3jFVyQ99az+KL5ANeidE1qAXuASQu/pZnFm8Ll2Nx3kQRouXdU0rOKVB4P9tChs0
ZMUDrmXBq8gWys7MH4VqcbSESZEIIzxtaip5o+R8nonbEXkSi+c9ZiGK6Rbcogbw
OP3ssOzJiM2CYM5o3wKiH9fEaN6SErWZFcJQ1E3vDEjVyi09luukYQJc1BgE1ctu
QqxIJuOXBMwD3GryBpgFpcxvYDg41UxAoRdGnEMhAmfwQiaHR5MhOauPTnoo6/kz
gaQXQfEPNFMMmvVxTDZohbXdkcjJQTmvloLN7Kiv469kgqiRqFBd0yuC5H1ZEtpU
ieZp4q9sn0BK/FS7gz5MZyQpHq5y8nSmYV7dqrAcSZzCwnu4g/6VGSpXTtGyLFfW
jbtkA1cFsqKjDfVllwDDo67fn9UmGjI6xpYAHwlCiCcje9iaHJEG0n+Xxcgi5vJo
kYbfpMJb1osuiAoKyzPc1BfpjXgZEe56hJKcs2f4J6DItVot+r9bpccXnNitVxIo
8frB6eO3b9ZA726dJWlLM7oCM9PriPxj40GAtss94OIcAR7Wg9OLGyJ+MSjcucXi
TmGI3yRB99e959VoxLTCt6Udu3cCZJaoCLvn3TPB+UBsJhuKEKyi0RX9krK0FWzV
7D+OrnYQlzCuTFlyGa88XUv4chqt7wnksk16JYaINNViu5NrId+tYx+IQJEmZV+u
H309bc8BnTwM6mo2xJycZAS4yyKyDKPiv/J4E121wlccbLPf4IONsOxWbZYT3m/e
NdIuRnXva/A1J149Z1asxrh3eRBUgpLd1yfVHiAsUJCDrR3M6KkXkThO+b/DM7cD
OuO+UACK8VLCS8433Dk9umMWKghTySXIBEVDbFrRgLBrg3wp8aZuohKcBZf+/f9I
a/nxHEqK9JyjhB/SHc4ZoxSNWCc3DTnuSAXr2LotFTUFj8wK8luyixAonDd5wcV/
V+gLNpBETB1dCGCbvPN2EFpD0HYIfRgdkHqPOVSM1bcL3D6S5k6HQU7FG8yaGB8p
NCVuda7VNHSEj64QsMbu8Nssnvawm6j9x48F//4C8kpeFzFWq7UFJo5zXQm7KrEB
EzMd/nEf0/PFM06PRbTjaIYYYXh6w+zDiBW4hl2blk/S1HeDK0uoYg9Uu2Qtmqb3
xuGoJD7MIpNRJGb8Oa1Lzs9GO9N6seMYxpIpwHaXkI+Jf1e5P+/3K9vIG48aty64
THYgW3LcKKFC34Nc9L13dXP+F/6OtV3qrF74Uo2u/QRoouY70TIS1ccIais+kVZ7
DUfljr/6z1OJlRQO3A+tDPMqhprmIBoeDrRdK6+dDX1Dcs1lltsRutNm2nVIKclc
+SKYOzVVriLT/3zW6alQn7Y3U/zXnev5f5GuouUZop8zwUl+jtEdXb/rnpwDraEG
BkNIUGMJ+Xbz9iEjotVT8vx4TkPylulqIllOpbZgdzh1HAat2WFORVT3T6oqMCBn
jsrYplM1Ij6ntmjl/6bqyaGBHg39LVIzTj/dS4WpAYncjolMC+mWMFJf4Eb5mRHy
VARKaLrVxOX33Ki+PmpRCyDiperqRm+soYwyIPIUlWhIrbo1xqYzr3aS5odbuUrf
Ckfz0de5lxZyoKecwykkLYvFnSOdD1xdFPbT17rD1u8ffEoyLsMfRzwCzfYSTvrn
7jrzB7wJkNITIqegtor0/0BGYlHD86/ibEbIl5rQ/UkBZveKMJ8bD2DAYWKmrizp
x0WKIP2dWj0Xw5Y68n8srhJsWpfmJuiQfjMx/7Tf5w1lmExCy3Fq51PftAECHyN1
YPLZLqZHfmRQehoN00HF/UZVvQBcex+HfpP/L+Zy3ozbcfoWyy16NjuydRSMp/sV
5LMCY0R5dh0w9pTcwfWoxXzJL0jWHON+vl0enyvwWiBQlW9HATFxTLk1D5gzV+ZU
wec5fYZjCi3fY0WL7cxNz8XrKVrBv7/mSXxKOVMQLzZ4MOmDnPR2XrytJnRcopLH
6mL0i/YNAvLaynmr0gdgLSv5pQ1Ta4rdfAd4HkBiHKcryK9t8hlPsK2QXa/Z/mWT
wbhSl7mkhkuiXr2S951b97oDPl0rU0SIvAvRSOy83MNwzecQ7JXNozUb65hWsZz4
IUUpJtyl8GzfCbUVBT4i2j34BBm7+AAwA47vxQIibAi4Xh5MSJ5DEgTaMWc5pEmo
lNgd7TmruKyMNaXxeZekiRIyIFV9BwggMn0GOR89wEbpUu5REACyxCvOv5xjArKG
i3Z38i1FWFmwfIORbq3nYbKF+Fae29LRoKGHpKg8F7fBgdl1lG0FcpxY30S0fuWb
1gsxeLMo1lSziRS8Byl+Io+75n/QYsdKZtDhdRJVlF7YdWLmxyHMJRM/RfZfVD+E
/T0u5tPlzZZ10fiSTbq7iff/JxOb2gdInIFVh50iTLglbppLtAJKUcvF3r+euAsV
4LJ58DKS5mwUVaajrJciNVOHNVcS0XMZhWDm1bNmqFDViV9LZJ892A9jdMFtYqLV
bTpTsVxuy/bXGkUbXwuhHrmqOfPnmhDvhAcEIkS7Wwk7VfXkB7A6jMg4XLiAx1Gu
egENzwhSs81J5lNfP09aRXJT9UwL8c6r0pjhMnc6BfvCdEI5rO6Q8vyfLml+1XJn
5xy5lP17oJgWG71dt5nEbQuiEXy+SmbBPwVp2EEjdX85xi9GOTmPN02VZ3cQFhx2
TZTHIAetXNRLKfZvbgDrdtIs0FDXSAMPYsKvJSIOCzV/0aa/GZR35IywnTeiLZjE
u1X15sbCaZtLyUxPvBq01QPIclFZBgtcSuqnZA/xnkPypEVG9dlxsotC5jyXZmyl
SHb8cUSLT99wvFI2KCcaAQMPqlAnt5Nu4bFg933RoZxW4IQIKPrORbNsnpANaCCn
5Z3yO3fZnP0vYtaDvTa4nbkCQQWY9Jct2rTU0unC/+tRMacg9ummbuUvR+ekHI/z
am22pnUHVu3DCAUwFCo95YSBjaneLXvdI1hXphiQzigOh0esPSulA9ASlgKSBUKX
mWUbLttrr633Q6zC3/hIOzsvG5XDXMiwSkPk5bolPESWuRJRZOkCPqFWRcbJ3uO6
6TnRyvGDP31A4mKb8QNxsTThZ7dCDfy2dT0WmjCxP/85SG9u8uuTbP7ULP729E0Z
F52wgB/w+Zx8wBZBfpHQLWQgWgOouJU5Ie1787PztlhRl6oVi77IxoT/L4SitWPR
0ISHBLtGfkbVARoLEXiPNZ3V6PuGOrIIcjVRoYwutDTqpMPj9NJX3saZaHs6db2X
UZfr4lhtzs5N7w6MGQU6qag8J8cyH5SFa2vUSL3ZHCDELGYdrQuE/Vo24AhtXvi9
E9NxOXF8a/hfKmy6Bl0VGMyWjfBs7zEbA3XOwl+ONqk3ejKSIJ7MHjKafpYIO1pH
iUmYa3LZoorOab92DApyQusVzx+RIE4TsU/tQLMLq3G6xrIpmu5FMQqu5nHrVbqJ
W2VvF8xGSocqPQYyrFUJvqyKzKqscBR9i6AF9ln+9SDBLlTV2ouc+cRJqCguKO8Z
zC/IBp7z9Nj0jpVdGdhtPoEHjNROMAWWL32w2jARhH2nNzlkoiFFFuyE2LK0c5De
FiXYL5E0anGASwSUeovbidemQjv36O7Nse+gLb6gpAjqzn5YJOv1dydJoBwBFvcK
loAXo/wZHJlGVTon2lepAfyBFoqbKJjLBZcabovZKjijkYtlXfFCf10ppYQp1afZ
MJ9Zf5ZYf7w/LU5EVizKhWaI/PUMeVXMHyLGg6rgR5f+dUpDgQRNnQ0xtpDHdftj
RlIewBSn6oF+pWqGGziIbZjQ9H1uAWiX117KNFHRy17ez24k2iNN+9D4+NipZg9b
u4y0VoQydhPOe2mbdwPurvyoeu3KfgBHl00V/p09t0AfYPlt7ud00BzjCBUPbtJR
u10lS+mw5NAeIkwul9KXOv4J3bFB45m2g0hATYOxZlTJIgfaNPXgNEhZ16mcGwKD
XA1B1KEB1EAORopidglINuKYNyGmRT1giQ8aKLUFBx45/UYPBEKckgEmN48s+hlY
rjjzsKyKvU1Lgqt3ULWEDhkGAp9PeKbqhRJ2wQz1kBj//8oIKeH264NPv7CLMkHv
JBxhEb1ZCdNgZs5usG10DNRJqewx3C8ycfllbUNfY/jSE1JNBbFC02YXYD83jNqE
9vXja2tjaYmwplqc9ImhPPvZOmnAUW9hfAx9X3Bxa1fEW07rpNp67A7xMqP38VS+
cb1DgKxjulv+7vwTMLSCclMLWLxqi/C5TDzBrUFaDRaEap983ZpNW9rAQOhZLOv9
MO1069TKQ+FX/8Zjj65agQCTCRVV6z+JzDu8wjMhEJZLmCucRQZge1L8Ic00Rd2w
dj0YIizraVi/ncFbQzkiP2Sd3OUrjRzQbQ7WfMspBeaNLZRee+vy2iVsDqKVZm04
Em8Y2p119UoMONO/TsJtblli53PxT1Zt81lm8IHPR34szz4jNXIPd6boxTjx2K8E
vfkqONeTxQXoX2jAqH00cdhInpZ6Jq9geqeBkOg72K9ZeKilqCOfFOOZHGESalmG
OVAiSsBvwYAb3t2qsXLW4DOfd09ke8W4hG7Bn4TGNhVIG4cfHJdais2qpiCLwVDc
vcV2AxnmFdjsx2aPUYzbF/rCgs4eQ5yjhCEYer3xHfgz3I/FRsFPVFhcAIdVEWM6
GTv85h7Mox+2EsHp3KS0J0GdHJcNWVAMNDeS0s0slbWA9jRUfisTW2Wz01sVXedm
7TL3x1hnaf3jofGc1IkI70SPQvtzkPMu2mTr0rns2ISiiE9jRspHRqZtJbxfHZI3
ChqSLdFRZg0SOAs3DmES28PPKZ+uSsOUvuer2Map71By6vxefuYWEOLPtFVI4EVe
yzSaGrdDc7NIjXq5R+OVmbZejzCugtJCLBRRh3GU67OzY1jZ8lil274OXarML2Si
gIxLYYUkX9WFEQPDakNGYcXfj6TvxLI6DBCXETXt+kh4gX9rcS2n3lHIkDBl3faf
O0jnWNyVsIlfYSsm7MAzpIbINjGlPxEu96muWt29/icejw9WTbcgrQNtOUlnqImY
LD6so4e25aXn/3Nyv8n2il20/romy1admIZE4NZi9yNkxJrPZXj2w3ujyTPz7ORv
qPq8fGil9xFB/nXxa6uDtKXinEJ/m6tO4OHY+RCWngPL6luD4RdkAOS6RPTrqQzp
iOiq766OKej2+1dBxUqHGxjLi6JR4LcvzqgPeTfUJ346L4IEyyaWAF4yayIxSP7I
y8RHsWlvjyfmbr2VcN3/EpQHwKqvhw48e2fVuQ0waqHTOqfT0SaJzVbhFgyPO3Yg
zZiBtMK09pDWEkph7hRo3T0jrfKgBQMu1O3flvF0c5R1cqjdtpGJxMwvRJz6o0sU
85zHjSMRyfLObBriU/28zIrbL6+U4WNG6ZU/tSSD+L+G12k+4dsfOPMmUKRlnwlV
WqIfi5m9D32+ni1yQXwZm97iAV+3x61rVzUU9lssJXkyG76nyVYR29kGgXDe2YFf
e7gHftAf2+HULbAIWytbZGDYt4FF4bl7kA0FY0KKhqXRnpePvnkUfqYul7QdGGUg
iAoPnY6nH2Yi/pKJ1GyCIE0qsVJerXU+TMrq2x4K1vnwnsso1FNqhN1EB3nXeehS
KY9bZc7blgfD+GDYvnRR2C7no9lS3mKJWftnn7HYmzYa3BSieOc70qESxbWHppEW
0u1IBnaOkE0Hlli70YMVNlDQpIGYP1nCIf6YtGZ8K3RWSdKPYnIGBVGuXskhNs4E
WSwzgWz5z3Clm9NIZgRCvVOF4i0ajlvBPlaIIoVN7I08ryKTN5FDj/Rt7RY1xdYd
EMlcaHmZ5vzLU/gE/80++l8hRx0h4hNjGdjBkBJXnb0OGp8590ESKtpkaaFlityh
0IqjS6q4CzgxPxb4CTXL9Uu69n6IMGOUq5zqAUV7JAl6K3xDocecADHO3D8dDCKM
RjjeAlfmlhPUnlRdgy2D3bYe47tQ1AlCcPvqZA4Ry4qAda/MMVea2ximgIH5zj6g
RsnTpv0VwAZFZeeURasAncTMZJaokADbL4Cj5hzJLVCqILtG1lNeEvuMK48FIKDE
k98agIzKupXLvprKc7sHXRdWN8VMdK2xEC0iUKk/X1CjfTsgnSA1SUT9kjleOXds
gwjiVhFylsGV47uYcPzLWs7ujilPkaeV4zcIrbwTWmq/RJjRDzG8uPmPixPkJNZC
G7SYtNHD+dzdEKNdds6wT1uHg2L2CDrof0OtJrxl8uVHTqdrwGBe1JNjnLh4GzNx
3bheKB2JrG96Uz++BS9vAq95lXCEx1103VixSAuzITr2SACHL7oj2jGR5sPu2EAX
mTG8gO30fZLAVzUMEw5+ZADwcn8fOWJve6PTFIt6YKZK8f2084ISVDqCDb4nvJVf
UQDVpCXmHb6PMJyRM1x1KDUSkDmePqde/z67ovVIPqdNercWGCg9eWgzsNFdyqQL
wmlOX3LKIwYblAcoow0wrPYceOVLIXmXjKA1h2L3EOQA8yl1DCI/6AChydpCQgP3
49p1hm0n9aaebF3cY1aRHMDOP0gOXX4hBTHt9Ak2XGYnO2fjIzHZrYacToEIScTo
V/azMPmuuKrAvi24gVO7egWzS3Rct3j0z7E0OdwmQAtw2YyRuXzYT5Falc0DbmcT
3CqtYTvnGXzI9949p5PYJPESoxySzCRbu/PYo+VXKrb3boy66bp8ZJodEj4/9i7J
iTVJB3QMh3xrjCGWHxQ/Bo9H8vtOXELMDGsmFc+LBn6QhGIj+5xKMPMbbF74d1HF
NyfI0b+bORRQA0Ew9rWLPKzSWUeUZBWtjI0lAFxQE4bRVmwTTeYX9oZU8tvjbhSG
kZ+yoCqk3e2E0UOzSeAngtwj1XePQR4sw4t+jhXPcP0uswzYHsuCAld1TDXhweel
QZvylEfxndltP4274Rzr/pzhVPoIC38HOQOH8xMNE+r9Dop03+MH3AaGMoD6xwpK
feZsy1kuq99nrUFEW2toHM4dmsTHVdX0QUFF0hViDOP0v7/hIvPi8QqiqSKYQWmB
/EuC4z0dQhPH8qScyME0K6bnjr7Rz8cMgKbBSrGTFOzfy5lKqHk28K8LjS/ygcAU
fu5/g/tV79WxWIzZgK2C7eFnU7hJe4Ft74eoFamRrybuVIR8LhqzPIxmlNxdp+ju
4E9EBKxoqPkQOrpOmtCEYAutXLb57IHjQF6Q99/Fv6H+tRP86mInw0vV8iy3hKT8
bV+07bhBXdsIH6RZ5n6t33Bn6DBK26ZlrG1/Dv3zukj9NVJRsSI27GiuMXeCLsiK
Zsaw/o50OS0VyzlHhl72NY1VqGJUKO7nZdL1jvl9o2tZjaETblxPvUWccwpzPOcx
kEyZrkUrz0dRlx3Jvb99N+H+0B/XzvPNk5IL5JbU/29tENk0StldObxtyFd0VFLE
AhzlN4JUGGeikbApCBdDTcOmzs2ZXtYCKdvGKxNTtEzHWLAh/aSySUObbpk5TDZ/
QervH6S+zlmjy6XBVpgj6GUDBu8SAQLVhrdvgDjU/2rq7xg77yjCW5bMu/TnxNz0
lXXW8Ra4PHW9V8yz54fwJD/YWHxDN5Ds19uRec5QAw7PyEJ/tGEqiDvTw/wuVFbm
n7KclhKZ/c9+eHKAl0fI1yiAwpKLOc1YP3kQuzuBAHkxMXY6aOW0N/kgZaF2pidt
4ufwbO51BkgnW+3hUB7zSTQhQDW8OM2O5AM3s8zMf9SeiGQpeHovqFs1i//8uCvz
5gDNpq9TqQUq84Lhs6BePvApXF4r2wOQmt28lCkweH2HsYh3ro7Nn8pSk50Ce9sJ
E13vVwKM4q/U32/+C6lK6bDNXduAqzKy+t9SecXpjZzv7DnxMvcGAtrSv1phTX2q
GC7cnTuIVeIhuIhVQduuXN5BSOb5CspwoQcEQyWQmKFEOSz+62E1H73pqx31Io6z
WouclNLHV5awEtZYpP7kO7Mt0WVr6V0gd+ybtJ5ctNI+d/01A/mHOpItXD6yCjHk
N5pycN1dlDpdNxQKT2KuC7RkjtnO/IglLARYbP4seVXYM6g+2s+T9g8rUBICHJzZ
B6S8we/wmp3da3PpeJTKd/0v6jHSoAXzH8YmW9EWkASeSy1lScGDzjy/CSaC+ZYi
qO2KSHYRJBcGIKUIMjDbDUqShDyCrQm2LK3fTdOSvXAA89iD+TJKbS1XMOejo9ET
Hsv6RiFIrm3hF9jAAIHQW1ibYewANQKyZo3UFgAImp9sN7Q5Vo7+yN7uSJjMC2Cm
vgJ8QN7hOeq4cGU8Ql2u075kMdRICtrkpkdujj6r/XI21AKjMF2CvI7CJU2yIAy0
Nd1z6CAtnihXejDIKkJwV0dFMDugjfPdX9G44sKA/o1zrBzVYE5+nkwCKLPDB96J
W0srl16cmfllldDsR2KdGxwXaVVqCKqrnbME0kLdK/j5fWOzc13Ctx5029VY1gNh
sPGWfmeOufkIfNWSzY8Y+lVWbGvfpAbw02y5Hhq/A4fih1U+K8ECEgQyPfNddNGs
oL2/hAmzfsRGd+/4+ku0zpzWGnmXhv4NORdJQUraHuzVwEmNt18QmkguMWRNCnB6
O3RHHkycaz4d+apx7eIY1xWPZY/C934/5hFFsqu9GHEbiZqVqpwqdx0HBWyxa1YA
ZfCUSKJYcdFwlcpKxkSb8vjwxNZEhxy66AtfNxSIMSi15rA5SmC/WWW45wJzqhRt
tOiAdsCx7DjxVkxrPGFESZDFV3Vtr2TBUmx5ZYT4q6Zbsnd1WdZD719KKAWGsuhg
wIv4MyT6+aJgyWpoXCez87iSgqH+qKJSDoHKSRg+xPbP47IFMkAV/BxHfYAbZqdR
ASgqvQrY3n87533wsmL7Fm7aT4xavMY94Vf8rbtTg5v408okaYVHiOiT0v/lTgzP
6223b3fPmkbPpHSSEvyZzbxE9syUklUwkhAmGTRQZMbODeD4qTRpBqi3KmHT00ra
S2Tsw3L3+4esjTd0nzezW2GD6s0Us305PQy8HlmIegWVZIvuku+q18MmyGrjPV8r
x9238vUsU8AClnnzC41JYXGyfmCs8vxl8O0S+OyZwPOoqq35t5zjCk/3Ee6zW7eh
5okZ/gQVBj7Gw8WbD84GWQ2yZn8B4iqS6cBZTL/ADo5KnohQcmNhlncP/mSunq11
1SAMbUO40ed4PHcvl8vr5xhbXEzN1011aJjAegoCeXlVCQw5RA4CGXRYKA6Nfmhc
9Wy7qUeZgDUtaPNEQHW6dkQtk3Gw8TEuOfhoR16FdU1bN+e7LneZjNymk3aSV+f3
1z81KUcg8W8pAveXyRgYhJqvc+ToWT473Ch8QqJMb/nwQ1pLYHM11DgYr9IGEh4D
fUWNtinSPfD5RktHwLrD7/i0jiU99sY+h69MpqD8DXENqzsMVB6vFq6itP7Wt4wb
GA7YPxwZ3ZaSsE+W8XUnLFerWlKETlhFZKP4lLKazhqZAsCBtaMm6dlau5KWV4Va
FakEoOCp+xsfvXJ0r6rB3XK0fRfv4AB2DV1AeCnLUZvbVYuflnEDrnXn36lt0llr
rugDP5sRSLgF62gKiLbQ9VXuXk45m5bSlE0o9QsY/rVAGRBtYAGXC9i2cFi7hmSB
F+6Dz433zCV9vbc+krCNBP2P6GPX8YJz2g9tyKjXhzHnBrZoIoCEVEdwjBqtTyie
AVeQ/4DNtLKA8C81slRuONvHiD0ucaac7XBPh9u2p4OicI7h3kjd3zmKstZYMW4/
XnrRFKTJi6eTK9qhs1PBad+gG+USRZnEv7LiEbimBaVqH25dRh5ycMcpP+M+wujG
bsrlkWYKRfa8+9BSstWjArSYP3n1XxOunoyjNqOmQqctCSa8Vk83y9wMnk2YPm3n
pexV3Z0NNC9SQnPJ49klqAcZ7QSEjQoXGgfbPP0V0o3m/9h4PkBUkpQPaTW6i087
R/GPD/R2fuWMdVz8Z8hdX3Og32AvTgNDnV3wT8sWtMUkaggyzwHZINoa85I2efFA
SwWOwuyPMmAgodKkZjdLaPjTiiPCU+dY1THTn67naoMIk7Te+upHNkKnscLWrtEy
WZ/5sMgDiFPOVAVuIupa74Dq0nymfjoslTzben4aWcn+6SBIsGg2+s+A3sOB8p/U
BUjJ59w4by25VYatmcIQAYWGSTMNmIXsyYFATiEF+RKP5RrSIvhd5T1h8MM6sD4Y
O/H29sQ7mPjtmqnjWBCAKMuujfsa2Y5wllvEu2EwJ5D0QHfGlpJDTOMDHkBH4Z1J
s5598IRh1BnyGLuE1DRc/Qwss8Bsgyawrr0pnpJJnQPtohT9mS6sgDMzSXMIGIyd
S3OU8PX7UNJOqv5wtCKOuijpWV+ekN8xKn516n2/kxEnKHdrwZQ0oJ62yKBgym21
T01nbBbcsdLpwV+XwILKkeu1KXOcNHYD+pCt0ilz0tyo2Dgrhl+ARBPBOVTeIAMe
nK+DQd1ygEZbOVnQzvdJo9vUHj5izisrVhNpKKonn4dlaPq5ud0i6uqThqkYfznb
d9lcdDtSG/vt1cExi7mcuh7W6XqcBfhruSjK5LP9Jbts+yY00yo53xm74L87AQmU
FtN3M/i1+670ccK9AU38PFYbuKZlE9mp7qCXIMcz7mvJOrnLrpOYfxAwrLs9gWuE
VfqFcMM4yjv+0vSplEy0sIaseOq0uVbsCP2GXIdS19+CDPviVsOgGd2NZvI+9Ia5
eL+VpBpNSaU2F7GSxcp6i9nLoCFuqrW/VWXpex2lkJwVG+koQCwAzizmZWi/qIqT
m99lkkYe/TrUgbs2Bbm+Tl6/LutlRy47a8Ic+NBEqLyEzgGcW+YMiZ+PkTmU2uXe
G67TdrNT2m1v+UsDxaSEPx8mn1k2i3udyeuoI3ljPcrr7FP93qJAIQEAH9tyxPUG
3BnoYY5e4A7avTBnOA7gljI1VZllWfq610elxJg+KvGyV7n4aWs4Q/KeMT9/ktaZ
tIVDNr1FNTtswRnv/CDhd+u2SN5Acn2iTkI3PWrbP+shgThqPgWKH8nfRbmJpsco
8APIBRjHBLAibdpx3L49WHe5sru50fheZ+AZoPXMT56XBuHR6a6IY1Ju06S3D76O
FAcagJ2U+rSIwvtfPYIYCIaJ5ltcEq4i4tuF9RQ9mHPIwS8JXrnyuAqJKq37HG4z
SepaAY/cCLOxyxoX3gnNdsaIhsntQuRVUOdjB6vqw5KfgemG2WuvZw3Tawt4WhHe
ei/iy0hZBM1CjuSx27NIuQaeSg7YmFlPDQTPY2IDNKDWyZwrgwupgFezNPds4Yyg
LH2tu3fZZzFQjoJT6TDobUw8hAIM/rAvNs4n2uBwWonuPd6jsVbpuuSmWRGoSpHN
8fnk3I2F6ERTOZVozewr/XVIhzp0FGSbp06twAumz+ABt749QfB2PsqQOOuhaE1G
9hQ7oGzK/zzhaEWBhC6ytBcS1AwLtgc/8CWlwB87I/lcyy+Xw8hoyEMXuiQF1G0f
Su1HF9N9ImUtkHplsKqP7pErMq2XCBvdkHzj9f6JBx/izS5HS6kPZwWDglTKhmv0
g5IcMmuxl0T9Y+XVlRrbBjsvOMzsK0m4hb1HROKquP5XDt1/CzgVeBYuJ9Oz4IWj
DcZ88YG0fA+adgAcfVLwc38l7kbYsw4kdtyNznwVzltHneQ5WBlt9sUwQccSwdyN
bLa7Ew+iPFja9OXSvKlYDu9g739tiwPo7FC4uQpnr4tVdZh1ZVR4WNsBVYxB4rKo
Z59gbfvvT+KNu88o6QzAOn03jEP1oZu4aXVD1f36/FBMxkG8BVnE4LkplWNWUd7N
b9sUVrvmeCtHAJB8xzFnqs9cWAB4yQQC8lqmrozro+PqGf/fkcjkfyOvqQQzFKih
PWL1QqnT37051nW14Fa76AwdH6GPKARqUMSDtw4jjZZ/eOFQP4FyCmiZ+6tHPTeq
Y2YsS3mAN4Sal5/iV+l1xtPIo1/H2Q8VcOalQswFDx8y9XhpMVSVtM7Oh8cS8VLd
4bY4M0LFvWwwTaGdCs9KV1so5cxsI3IMhsSEnIK0MwAt6iDn6334+Ye1460m6PoQ
xQuf8VsX1808DAu4UUHxLZ925cvMUtjyxguT8tHjvODZNUE8fGkeEkEIGeXvFOKe
LDxMqLU6rNfSVmjasdUTHmpJyKe+eE1YDGbk5ApwTgoOVQrHALjmnVwnEHvyaJ+m
oMsVTOeXk/Wob8o5PUZLlaiO5g8pULiaDQh6zQ0GI6gy0RVc961d9akMUWtyqfk9
LHpGIrgtAhjccUZpUP9gOSB+DOp/EOAuv90arcyNzQA8ZALsj2g9L2+nLEdaG4Cj
JT7VzlHL0mAC8T41H33Lf2I/IZCc5RZDxbXFttL7zgjSnB8tz9mx3ysY90smYyGt
YonX6366cWdAQ8onuyVppbhkEHpFRLfjDxQOcBRcVaf4d3P2RQxFxKoaje6q9QZ7
W4OQXvHJDMshER79uZNUW6I2msdgfNTFNKJiOjwu/YdfITi5ecHiE+wP42e3WeBw
mwKft0VGqTDEslMrYZBi5yLES6jyXBO4NU1W1Awerz6C1MefVCkQ9UhsvwGY2P4+
R3WhXrJJa8l4AilY4H2vkUbbsP7fOXlOzxo6AjCcwGc0ur9LYibfh3ji4GdTyuui
ali/oxI1rR+pJfCtQJAb+6+OXHwf9vkU6Oak9W24VDDSjzq2Z0QK6ZZKaO1+3DqD
vsZoUeyV4a5azeDTxqA4zM8ndBLLpbqQuF2Drs3ptXMeRaBkFtxdEFWpoNuRVaxM
gXDM0k9JAc70CYaZRwW7Txx6zKTDjMjAJda9+GzIieVetBY0hZWjLRwdfj47N4m/
UuUVB0oj0mJqJWRz4cvSZlk7ra7uoqUdaqrJXrebM9/BEWPUN9QLI8ezMq9R7gng
NwcRZgzM95b5Mc1D9BW8uAiE09VSx60cveJbLi6sRz8MOLznkjHhWlPk0/6IrVKG
6678jn28J7pbeOEjgV24j89CysAhFY10cD/nB2+ttreKzgq1NmtXHePbUWIdpjzP
IYpSioj4e4CmKCshkptrZJMovTFi7sYTFclOMbjZffEcezIpAm5eyOp9yxyAy75l
igESM3emzZqywmPZYQJB4Yt8fSY3TSGk9GMGEMP2cHkz6l/1AZ9M8bPM1t6yanSu
uIlprc/zaGKrQzZanb5C+wP23UGTlT50UoSYqnUq5bu3/al9L4oU0Qxq0dItRyNg
CJq2Pt1EJg8AdZyXZJJ8nx3BYZuvg3CWctPgSnLB+3u1gRFFfuarZUp7S5vP74A7
CztKatndw3Pbd+gsraQS9cP/JeLDrZH7sqKyhLj+1v79ftE6VmzmbC1Oz6UemZOK
HdqSVRK2L0E/wpIWsR5t8GW6gvDyuoThUw+3xIXQU8xPEpswye/31fnZ504VSUQz
dHQlJ9YdLSnziifjV3cEm/yXc8BkXrpJPCGu7NPjhxQmlrawboOQUd4bJwsbcKeB
GKN/n/lhjuzb4bbmK81QUX4DXnPzjZB8Rzv4LwpA80BBWjH9oMnfzp0fhbJSYs0N
E8wn1ntmJvnBFIejYhN9hV6yBzTxAsYOZsvvqyw6RAsvLa9zhFCMkQMrrZrVwBut
PUGfrHG7EPv2gIIpofWUcEy2I1AXiJEUDEoEvxFC8ucUVvFA4amX7r4rxqCooHJA
KemfbDtKY8NZqBLRCCC86Qy0I3y5fk0QaF07jaE8QJ05xcJic2Kj7yzldbiMcQUn
bQImqBDebsysKXxFZ1f02IRC5kQ+jsG/SlbMWWE+9wFadyfgGLMF9FEfGhJKF2Pb
tRaB+H76d3yjwXDuunJ8SDKUFsLNno2rjaU6U8d0+CiWT1CAEwUJElcFSjdF2s7p
ivqSjXzmj0OeCVPCbfaiPV6iRwMeEzMJola/G43RkY2BI3y7dKJ4fnOWVUW0uAy8
v4b82hbe1QZ0Ukr63O3Ey8xy1zDbCDA+b5EdJDMaQS22idjyy+MI5ohxeUiuo5nf
rYm0LczwpPRPZEd2iuOBWZEUquIuwaA1pg+jEAkiB6Aw4r3kU2m07o9RcJ15k3dW
mwAo+9k6ezgAFR7NEc4HW5CZVadsmbXbexHVxi2B+u09uVmvIHUk+nX3rP1zGxub
Mgwi7uUgiGaSGuW3n7cdPeLxDalmir9ZsxEZzTob4gO754fFYxuIJ71XG/jpEP9a
Hc7e7/HJv1K+Xzp4RfT+5+dIcyR+HpI1QA6cDauEkGLh4qAQbVIx1VvkSINNz/kL
07/JDhrZKmKdXi6+tRvdTrnMzRJihmIPLfHtj4cwSFsxG0lidz+oNwcgffcCV1T8
4KlVqu8G3X4YxAZB+FYhJ/ODfkOMAdhoj4rlbWD28pcL8sUCwQZNHNPMKRAw+Cgy
2JEf2NZNNWCY29PQaF/z2thodK+gEDKWJnKRl9BAGHB+P05gXJKL2LVKsdFcA2kN
1XTlwB4B3zzVRBWROKK4AvL1kffU9GjNyXnoCkK1jgBnNrI3SOWZ6FyOVWwt+w9F
Re+ggDyQyS+3rNruBx86eV7rGpPixqX6jVtBt8cqIySi5nOwKJl7ZSl1Qt39yUM0
19RFgFzrxUTfNfVbJIRg6pSOB3rV8pQ2Mhbz2snQrAYK3nkznM/H7/iZXSiOAV4i
I76bBrzKwBcu8pTbkIrUNNmi0wifj8b5Gr8AxjiPg+MwZuKr79F1cP2sOPsD+1ug
kBgtDEGXis8PTrK32dqUDTrEz58F63dMoXNKvq1ZWqEs9ttRUAY5ddle2sMcA3WO
uz/cmv8BAr6Ss19xIseTYyDdQ8n0qXQG29uTtxzHvwatOK7KlSBOqshG/tjZEFcT
aluZriyMjB11KC74uConkiJU6iZvy7kVvLwvrtYhcPannuv+UA/KmWC7HVYTndF5
vh53O7nEZzbzASSz5yPN+V8kX30QuQP8n+x40XOW+B6U+lg8l+VaUeoHg3211F23
VkW1/EHpY5a4M3zvxlVuLh+fAe3Tff0Q+VVelsNrofSdFkuGX+fKP6gx8n0aCvsG
oQ3RM5RueI6DOiW2i6Ip6rXniU42Rs6wgSWEz37uWCeummEfxL3Dw/8ztfO7SdKt
8y7zti97DpKfUpGbZ2Q1SkOmSNdDyI20pUlhNfmi0rMLmEVW/geVp0AFm+9Jlt1y
IZHUF+P0ZLTpKalPWiKYSl+OH48re/KND+v0wELy9J1TrqUHCdK2NAs8neB8aKaj
hqYTaI7im0GCRpRPvN1jcTICkZCJYKPW8n7JbDdzplvuzqoLn6hQ/sw2udHNIAoI
4lWeigplANu6rLN89Qkkl5hXnS+H88t8w+F9qCSE0oaIB1Ihg7Ns6yRdBFz/XpUq
+S0TZyOEayoRLmHhU8/A3dqbg8qmfcnPMQW9O0REWlpNTqVNspHwYoAY4LqRpthy
nlGF9qvOOa96HhQPSIKSK7sacJibGyiRW8qxIQLpgcqtruHhSs7FIViOarlXJ0fN
uJPlIptulmSzYF0rDltGBztkYQT2ZSm6G6MNT9yCqGDsYvBdj+VbVn/hKlE5K3Lt
tv4uCkNpGrBlaQlBczz2BmoU4XVzKdfRlT+6V0uD8MusAPpAuE3/6uv12Igwqv7s
61xPKE2+W690S2YGhLOSXd2sKXKMhWHGfcZv3tX2NxOpuYY3/C9E2H8cEQa51Lfm
qytzjPCA9SxyfE+XSkI0lvsIdi9Cf7eDv1ZLeZeGigtNTLKrBYNDycLD835sfUBP
I5BdkK+kAoq9tjDtEiwkupB7RZaorBxiu5137UZdw4Xa4joVEMzoiphs7cWR6nHl
vlQg7rCt48ZCf611faDD32r/aYVMFm6AvH8f7xYXYwWqK14NGgxDZTodHDPORDXV
gyGLOU1dwO2h/Qpa2PLIeTGYN+0ilrwE2sdQ5vO3XQ/qjajcERhxAgefX7dlvDgA
5vZoFU2HgaO9W1cTmJfkIwinTt2RbhwBAzkhDbrhtdAkiW4SoQd3WuckOUeuMSPD
us/5Qc7GLmKUbnAX4mCYVbp1dU9iG75UIb82ZUOJ3nokA0gL54LwaWMwT7ZwFYT4
Lxgu7KtyfAiVf+2S9oFsToco+H7FMUmhg2G5BYz8wvR00vEn446bTIlEOy49XHv/
bvRrfqcaQDecg6IE5YoY5ch02P04MUk9WEVflnqROHRZ7pQ8ZsyEbjbVdah/Tnsf
IHQ0nk8QcZjxPDnKD2tUk4mejWbRVgIdffEPKgRflT/zmVgLpoi42t2xSb6Gx8s/
GSfPLw339KtziOoxRSmTh3ZMLi81FPRs3Vm3kfiySyTMI9CoHOJk97txMb4UkoI7
OnavkETXCZ8hQM61k0S1P0xZvZYYgQkoZrdmDEAtH5q4wB6xz/dYp+x/31cXXNWK
GAAQs/V8j3ME9dDSLNJr8d7bW+hNtX0doV0At+3HgTotAfKBq0K5SgnBw/SvhG6n
a+kzp7u6ru5FwTN7kCtcFMXEZY1DJInNgo7u4us+ZiMNBpcbeHCm4SK6tlD15qUv
Lmkln4MI2GmMB++JN9sv4TyckgAaRedZkfu81mXi+ChTOuGzII074xIC8ermZ0zg
6T5uxy9LcppjXaZac1nj466X5okRBoAhmNgjFYaN9ZcNpXfZ3pJZRc+eCXF4eY8n
UqGi0SEtATlrn8O2+gLItFEhI5eyLB4Kn4hDnlb/Ww/wPh47/fHzdyC061/vRb3x
zpsQMiMM7mj9dN/RWnjl7M2z4zcd6/voirjuzn4nv7vhp8Hwf8DuGzPYJBxLTL1c
3pCk/82huUPQVIF/jrebhNy8L0+oi3x7UhY4OjmwOPGkkKMhm3trgq+k0HUvAudZ
wEVZB6Q967nQSMdLGCy9sQj1e1e9zE28PvV9dfDgbQ59kg85zSVCXn/y2zYD5Oh2
afAy7LV3ye8tu4Ux/UI/Xj8fYokYN58/IJJlv3QaJdcVvCw/mn9BBUaD8iCGOoFI
RSddMhJLXY7NKXwSKTa1KzJR7rZyARnZSaVa7EegG7x84pIIK0NvPrOIcerkLeUH
sEZoWpGF2cEJc4p3tdUjG/p98llwRbK9B49rcuBgSd/3BGULQvdzCVUoOiIPfdsC
zFUlh6ycZ7JdJ9ulIsJYr06yKZAerXACEBW1doLBpZXB3akO5TAR/3od7ykUwDeP
mcYahRfUh3JwHICe21S621yq9b7/3CBIm8Ejp7o3V/X2ckHmBr4043pTGG0unMgy
CRDqU9pQEnRIgBZMMrWMMqFwiI3P5lu8fMNm6vtDfN0QkLfIBFwH6C79NGGZdCL2
ZehrHcwNUiiDdMpZosh8vPxkgDK8NfFWeJqVijZGkVIy0f7fBKhOJ6aaAA4vLq3K
PXWkczwxdRFLqCwrAi7c7zsTFM5sE88TtCscfDZ+7evzOiz6ro2KyJUOCwiBhGT+
Xvp9hnjnYH17zDs8CuDN8J+01Sec8znruVoJgeyUKs6xZ/92P2Kl8VD7ghOxXKjR
ja+Moo0pzX1kAVxiX6v+z3/dI7elJQ+ioYQFJOUwfVTbiEvzx0uoGw7G83fNhr00
Z1dEfXZhzyH1cSEbg69Y1d4TQjmH6UxSF3Me+g8EB45su0jiOV9uKNbfWhAKf51X
HEfcYaAi4bCYT4SVOxJIvZQromTfqMMHXjZWyOFFegIdwVOvQ1WGcfK8ATggnBNF
FP8H7xcayAaSSsd5jDNEKKDUSnNSWCIseiQ4kZK5WY5RJguQUPOyBv5V9jfQ96HE
qN0HyjMH+B8FsSx3V+txoFTECU7FZUorPcbFMWDMkA0/4zq8csl4BB0tCpdWE1uS
+aSAoNCpbRFLoJGKv9hKcfLuAdjPKH1DhtnHQVk3iAHvbntSrtlw40XY8MPCCqL9
gQ4j3kuBhMNkB6DmE3zL5SX9tGdPtRF0gCzOTeS52ylUNNochNiSTJgDib9ZQY29
yH65lUU5t0vYrxnxRJ0pRHejS4TA2skVoRDpPGPHksQRp9ZczIRW86myfd7bH6L6
8ET/3OhFy0O9X5uQCQEDlGJXPjclpC74/5Yr9PV2UxM0M7laaZ0/EPuUZm0KD84L
wxB3nAk7yQ42+5LmW9+pdvtj19lvpO//882Uf0LtfKcYkBcpsPAR3t3YvSQPD77U
2HW6YAUXw4iL63DZVxPYWXAUQCmsT6Nd4zkQM5scuKqi7c2ZPuQWn0KsM0j3O8OL
IX6UeDkWPsK6nj0F2T3f/Nvzeu234rBN+L7A76EcNyV0XjLtwo29YI28qu4OXhWq
P7+SI45d9Dk6FlCMY5qb2B/c/Zf2X9cjBI38GjEThJDHD6LaMJNfCeG0FtkS75jh
3d4hy3U42xu2No1DXGzA4X7eVp8Pr5gZ6g5VFupjRrG29U5xcq8fKCKqRUf0e/6Z
Sc8MtL6XzjHrwQmdSipHXWi0HFB+nws+BvPZWq6WssnTC39PdP1PMnVY8Ipz+QGj
yl3JMOXiETwBrfkZ7sAYUfhM861xunAZ4O2DuLoXXtl4HYX+8eYI886mPyz7831w
xLKMnJe4oGwR0Xi4317/rNnXZfvNCT9mjmi0BSYfCquvqtmvxZy/wpJSZHmLxtsX
A72toLfKW/Sq6o3xy6OQdTOs9e32fYHbsjvlMHmXo1PQyeARAx52MB5aiQuKBMIx
lP+x3EhANtE8HEQjvx0RsIqRWbICVqG9ssIVTusdUgGX0gZU5BZsVAZa7a5iMAmB
IwceYV1nZTFEfkmbttWd+4HYa5Qf2XfCLvdxkSljbwJ0E8WYSxttQOTrOp+DK3hk
1M2RlTuQ6QC8AGlWqQILtwPD+tQgmJ9jPJAN+XsnozLFxCeUpABt6YQCzKljol6K
FwBGzS4wFSA19Mp9sfgxAvy4ebJin3Gl7eJC/qulDNL6NXIHexBl1gxuQ5vtx9aD
+UuK8pqmuFQDZZCWPJCCdkZoPNfzvZiuTqms5okSuyvzhYuJYmftw0NLyDg4axIb
8kdvucsQdQhEWK791exUlkhU20m8q4w/vMb6S4mTUzGxHTz/6Zk7PqaTMXq8lIIt
79BnvPxhHm6BUSTbGKKa9NH4P/+kBvVg+MGF8eBcD4DUVrxuYPv7y47qLz6d1amk
h1+ReH+u7KeXhpm4DVtbPyqQc9YSm4XQkdVeYwcJaN/V7FB2gSduuWxGlu4eK+nk
oy0HwllbKJVqcmrZa8CKrs33w+MLU+bZsv3zYJd9VMAO7MSlUWJno6PL4VjJvXSg
mFcQ+FeV8pICI0bIjMTZt3hI4ntft3TmWcc87bP+PDehU+TrY59z9xphqAzd4OEV
gxju1hp2fqQj/o23KSpF7ZbpfTUNMKOUZeWvZuYYa5R0sOkZ7elolmMckjJKQGle
85o1/aKBJBXrrxrrQyIWS2P1WDcRUREWh7Ds2ZVTkd8fRaBP0Of4TdiIIdzkK9HX
vS/DVUmsa4tOZ+uY8WgiQSuv3HNJoHf7KFkrS5vcjjXPdTLDxhKlR6KUti5WBsOY
TSQYpJKGHB5GI3Uf/ERCes6M6mBO5AfeUYTk7Vs9fH2Q4M8xG7moNWH7/oh632hs
7Kk8PzfzxMLQL3Xj6gR3AAznBhrYwoBBFbIktc3/ujVBg4x0JsLVojf6dS+NOckS
I+iIWJaX8EcEMfXiBihy15ma47UC1bQ9/0kUNcg4TZI+BxLJ5tXZVqjWw9Uct3I8
//FWZSkxStx4R7P0SD2uyZqavZI7+A872RANzk035R4gjX8iWVRnzicOAxXCXy+2
/ZwYhY4L9e5uKcDlGryaMhjVC1LyAKuvzgQEeLs8t5nl1NheyvraJOY158D/fDT7
ZOt577492P7CVypXfBsP6hWXsfgyUT9TwS5ZAiteb4CyoPP1ZMKH8X7ZTBnNnIQp
CkvV8ntTP7lrXTpDo6RlCXQ0lCZFXzhAYYjAhFIQipm+0qlU+mmETf5JBbME78sD
rX+z+X0aYB6Bx6OWh/nPP8pvii/YUlskvSNvZp39ExVQ/CYcN+E+cqusWg1NHnFE
ZyDRO0Ca43Z/gg6PvoOJvWw7PrV4gRCLnRpvPV+FeuVlYvinSBzBU9cQBXnpxCPP
hg8HXVgSQC2F6+LDdD5/QReraZRLatq4CdFZYgdiBhr6OYGhv6XyqCVewxMH/IqJ
42d/4ttZEmPgf4zoXpSO2QLl+jhWDr6Ygj8mCZGsdOem0vWnGeLZE5QMMI6ec1R0
7f20+HxNreyKURvjXKWni/ZIRF5yWTM2lX8nh4IfD6VvY/F2ZW0b4i7ahdNDsugx
V+mKeGVin0eMij0f0/ko9PhZUtKQCk3hJRO37cL/GVZKqDaX3oyQ8Pc1e4y4V3xu
2/bwWM+aMMg3i13ANSrpz2KDQtX0hO/t+Wv3pPt/skCIoIFVG0NJm8lSFg2IXwNJ
0epZ3oYiXfD0RvO07FIg38d2uQUtOgjObuu0rfL+el3jp+2cz9iMC4x5/LyAtHuS
qF1+IujjlwI5CKkGrc7dgDxe9/PS8GuTbFKCtHwXKrJEuitK9Szii38CfmtJYnOV
tZusnpWqqIgh+uH0ZfW5vV20NI4DiUvpYiVuST2UjTNvugIKy7HfSn74GdskVnfW
1xWvCN+uh1xIheyqA3QciuVOesSH88xfr133Ygt25dHAILvcBNYcGjsT4HNFWSOd
t01PZTl9HDeIqRcu3C1zqto5vv41s2ZSSby8Ocbso9guOmZOagvtmbOJhZn9/jf1
KNXqWRT59oL3fYQhs9tYttJqXzJCW2O8uvSvhbQs9ZyqLOglP6cVXDP1WbJtI0Ez
I84oGBWy+6hcU3O+Pfl2ICr2u6Q1c8fyaeTgaaD4QQ396sWFAMTsKjwxJkWs/y5y
MhnHECBUZTziFn6nrE2Pc0gvcHTgVJNr4yKKDVJP2y8GULQpE38XrV/AtmLITmJt
27feRDsW3t37IRTPoaCukKgajoOyDA1jxdjzIKHxSmG1JLC/ZZwN6HHvTT/m5Wym
cc6DYBrR9haABOeoNJ7X6VJE2atj2U/BAD9ZrOFStCnGuca4UXPhgvWMIS66kQUs
ZY1crqSRWiWqtp7dbgRmBGgkYk7qyknvFTFLQVenSwtT8c9Eyo7hHylz8wokdez6
wH2jkP6yRQhryw5eFJ2hqnCHnmd4p4IhOSP0E6hnZQcStcJS1YhMbOxr61cKOZ3g
x2ZLIWNLYBxdzSPTSwC2bh5hCN4Zy6NHntB70WW7g/6xnLleSgFeD9zHEnGwLb1N
wiOO7IJjabiCnt/ogto2gM7zuH/Xs9QMC1PVLigcmHJ3NRY05qs0vyxiFSNt0Bky
s5cWyxrg6wD3cfjPOmzkNwFNB6d2Kv/XtS17qHpay5YJPMXU1OryugZ+1K4RniHB
MwBAutJo9klXojFVl1CjDH74x0CS1Ew1F/YalbVfjcdItJw9ccwtiZd6Jq1nS8UV
edl8djp2z8g6y6vgSDSICV9oMruEEJ9+V9TYJvdWO2I+jKPddYVHktVAK8sFI51G
/2xrPCGM4Dkihttyyb0Kp6rnnrBfW+sc5LYXKLo98v45PpqYHYBhX+7cbq6TvHtV
5/4wKf719r/7D2lEo5evj+RUK2GKz3ciTx9I2pW8B6M/f3z3v8yBAxU60igCiuBQ
VSe+vLNxGtfqb9JGCxLNK78bBxkSP/fY2+iqnrPNTlOHBROwrftquH5IXSA5Ey7d
j3SbNr/iui0w5nnezk3kkxVa5RvKjBssnp8MYMk00MFO+PtlUNQwNKYCs+c2REYl
o5SF/9W400drLru0Z1i/OHTaH4CTS1TL1u1ZFhkrqlznfoKjy0dsBG8CImU+d1Zb
DefnNuiDtdM3PwCLRoADpq1HH+wjcrqlUWYzFvjrbUnkrSqrJB0LyQIGRfkMwBZj
RIw7I9Y7r+hVKg+zNYvWenQZlkstocTT/xA1BISMuKdbidQ/QTRE3iJgsBzaiuJV
IaxVj714FEUYp0T14pL90fxvnu0jpBK+vAdgHbcyepfTKS/cRRuYbU7jz/Lj+luJ
wERqtIxwRriP8XREWGJAFKno1RQQ3DuB+NDiplMCC3YGTvg4x19TqQpVFbJVOv3q
/G4avYho3xKYorZLi5xDzDAWVQJ2Q+XKNnfpd6RPy6hPIQ6Y+Hj5ep8IQ+DqjzPw
n0KCE0Vxx60VeN5PbWRkCyQ7gJS9fwAHK2E0GMVfNanMQEQZtXSgxQSn98iRioF7
Ij3Ebx8mIVnke5WTC0JgdEtzUuFcsdsb7mLX6vG5q/f6eHK3mtdUiiPS54LgME9H
4/6mUwTXedtXxX4091WMUJQUCYdQv0t8xnViZ7NhB7xJ9yhY2YuanWuNjmROJRTn
MRhrP0Q8ePR5e3VZBCEaSrrCoxZA1SfNcpFQVsNh2mQTaGCGkWIEyIeJixgsEVmg
LN5NVzbn+1Yv8Ntgkyf+5ixL7x832DuQ+HpfoxdDan7SHfuWbLij2LywryeQydjL
qaDexboc3QntCbJ1LyC2mM/2dhkw08STh9tlNt47NEuAbfoB1eG31XcqpCid2gEK
Ne4+oAMaSO0InErKl+JOxuUs3kdKSWJC4WxkIHhR4aKyjJB2FX+rq5VzIQxkmB9U
pdkgWMs3gf/q5yfeOUZoWBY9kVre3aFrKuqkJqE9ZJ10l75KvnoFEiEkUmKWR7wx
5SdYDr2ClCUJUv+m29kH7hoUVyCfY0GeY+F1QnPsSxqw89RS2YN8cmTWDJdzn8dD
MbP+M1EbjUVDuiFYt73kpWXbRbZQ+8sL1KGro+tzVyFIBCmFBsZf/I4pSflmXf+j
Tt0QNskemXz7UZWfS33vnFi8izL2qUWe8a78XX2FeGEx8MIwlP+u9B3Bry8Wb+pc
DoNaWiLSkgvw8zGxsmEXF1rqytK+QjKTEXKT5jNqpAUOTpow1+09eGvWJ5x5H7BO
C/GJT3p63jv+BFHs4fOvjfDd8iYcIio17KP5Nd/AKQTExEabOI97zhZuaizI3N+0
lg56xf5RiPwPN9ir8SLPIe0RVyTPHN8jrxDK5zAukRCAIYAVInajM4BRzzzefegc
w7SCp9JSHSf2skiEQcENUl7IMF9Njd3BiU+tCb1Pyth3OPpZCTuh4xPgZQ/92Fkt
pIEayQULsNPonaM1XhgUIl2kmxXvkQkFXRjGowaipsPVSuIXhYQyLeCqL9UrB/wl
6atmoSiv6mtlG4OYqYblGb+WarPA1zy9OFHYJEUCK9oqXmShJXDqnAiXUSoF6yST
cV6QxueOx9QqppxWrZi5QHeKzLw38tZc4j5XQEk+k+CjN7vA5hO/8Yf64c4GC0Bz
4rcOzAFFBxbof5qOUCz7sujVJxbL0PdMu+iPAKnRRZBooF7p5zDodvFlEtRwZNVZ
jmvMdjKYNw5nMBMFY5pvwSU4Yn5eI6VySF4XUKqUSv5b2vbJgHuE+8TfzS2e1787
26bAHOYFcN5phqJe8IvzOEqvJN1A8u/MhIrY17antam4RUMULt9KnhSLuZFUzrw9
sEtLJfcomwt3ySPF47oOXL3IdWn47khOADxJ9PZs5DkaDAKr2kGin2BISV1wN3Nl
iJh98z2OsL/JRySLL4QCWaB+SLIE1FJLTd6FByEukW8F/5KvCfu0ccCaU7tk8EeL
uLudcYiqBcOoGEiE3Gc8Z7U8T9bHYJfbEJLPL8MrCYPQ30ENT3Rnm58NnE1AWOZE
tUbfp43U/FLQeakk7uNEked28yZ6hQkOML73rKiWZrCtThhSwqiQmHELtGCGw8qA
+NtGm9z1DmwnraZSKQtCoh60NgH7J360ZR2Ox/xE29bAQ+oRe89X7Jo0REZfzMWd
X8oTjNx4PH6g8DTBfUCdzIBo2+Mze5MnyVNs86SMvk+OPc03lNTwL/I3q72NYSlv
SWwHfGdI5tnLFByKqLY6qKYCUo2kbaAe/5OzeCePwuf+F3b6IdQyAwub08K+Nau2
A9W0K8Dw+Shoem/8WmLiKU3Nl0hMVXE2pAzlFVZ+5elX38P9urVRXDLvy5OBrQb8
GesCb1tHtpY4B9xvCaQvdyQyKDXUWr++YClZoqNdt9Y6DPm5tc8jUckB/dbMWrQG
fi3HPTw369qWRtw0dxZ2oQMo9SonBK9XIUZd72nDkVTBdYauLJgNachwurNDTeZj
4IaQirHHspy+sv6cWLC6y3rf5+zMEC2fztETk+flMnh59vA4VdhymDeR7Y3zJVli
aOi3B+QsLSIehsL48DkQOMi7BtDxZmRV2ocWYWSj9PHdFAyGtx3OU7D2ItPPpRHa
oSsYVsNV3uP/4sRoZEVPvIh3vVK9REjsFMAiHYsAxs9QCRLvpMnSLlZb4MOBVrzl
5uEl78Ghhdu0ZbiAhLaUDm1wEiUCFNF5RNrBmkIVQxzjN8XPrXqrfCQrBxL4YohM
CMbrkafmj7QRb5uhwnkssisEm8Ckajuf7+FhEon6bXNf3tcda8alguvnbKeu/bwr
leogpK1t43qJ2DsoiWumXcBC+3wllQOMzr2s5tP8VYz0zQGIrQRdebRCvp+X2ztz
iQGYrWkhRYYHLkNb5JKL0yE6/cTrdwHPVmAlmye6b85KP/T+Hx1DVmO8DRgzISnx
AYdqxgoYFA3lNk6ma+PTuwwoPABDMNsTNCHVw7K7ba348Ml+QxGAL+VoPRI2rDVx
slaom8tFJGPnyPYUyx23z2S8X0LGavIIQ9xH9JeTZE/7GrzLaTkJ9uEs37z7yOvy
FtMN97tls8kSKXicD9QYzRFdQjq1xZqHidLl156GhrcRbBD9hkyP2JWysCbUHf76
oXK7ayPj3EinaZeCYNinXeVcNUOSjPvMQWSAXFXnrOUJd8u02SKx/AUcZLT+p2eI
T8j86JlceBynatvo5P170nGEgwUVj6VgoEJMgmX4jmrA6XKhJ1MnXEs2PqJ8GOTk
G0Pw3aKlqnIWC/+zAy99Suqrso/Cr4UJ7wTqeR2FZeLenq54ul08jUVNyuvql1h6
0TZcA+TgV7nrBezHW7/M7t+09xjprO8G6sGzyxOglAAp2lOYS4biEgE17sXTtH0Z
ETmVBUeWQSecU6SqbcgzBsc/lJiy7IrYcX0nhwGNYnzYZMVSoY5BgWgzDW/GcNtD
lwFi5p0Bor5WpsH8xf2vAjBDVOuEqNU4v/MtbuVga2hgmVzW+YaAuDNjKcpihHqc
rwUQUY7aFZjBI7GZZfWBS7eRPiZhCfr/mmlJbMcqcTaEHnR7R1/UgdhUnMq10njD
i5y7fEHCa7wK6ufnHgmu5AMl47yEmWTeNcYppW2XpjRiu8Fw5qEShvtIzTEEE0oz
xsf8vVjbhYxO5yNBINJ4PtbwM83DGY6x874N6jy+X9dujBUbQXoeWLuk+f5UNi/h
qCT6klCvgbXvRX1sQuTo9lDPN8llR9miA9bg9iQGUmHbUlK3LC6rg7AriCdKJZss
UPCV7traGJ6oWebwDqlHxNP6FLqM7QG2k9lhYChelrv5CpZVillXDZUmLz4ceqAZ
fVwdKtMMrbHawgd+RUJ8/r2VQvH/sEh+U3bsQL/K+hdclFI8HwiIri8zjDOMl2n9
+QsUuTIqbjTFmR6dpSdWV/WmlGGgfqcMp+OllB5WLoEaPQValv3MKqP6fHlETDl2
O0u2L0Dsn38hsSx4cdyu7pPnzGFo2ZwQgccg5nzG9DYGXu0VCECLJnLTRYYKA5uh
bdszaM0zeXfxMW2S+TchkYE4Z9oa+WppjfgwqIIqF3gJbCC/6aS+CiKZLF0d48ef
vJuh5pjtYUgChuBkRnmYOUjMF5XzLs918FXaZWOzMTBF8HDX2T1jwoxd3UeUvM6K
xX1kJEREwZ1XcnDKIIQITVwxxCdM0Esa71BqQ00I6VQWEI7RAn4qMxG/ol3I+XP3
Ybhz0uXZDt8mOEp1GVTQbJ2VRg0p+7p4omqShJ46EZAxsmXeuxrIQsDFapvj/80j
6ry/okI+c7kuSVrxBWmIP04riAf3nP/cChzKfsjJFKtRVdWiGL+NL0b200fBzdya
y6Khaj4OG+2PlBGaBkuqplD6HmWS7+L1MDPEfbQmEgohQW3ZWdmzag9TTVD+rJjr
hdvm6sMLZCaHld/Kw6yBAqeGi3pkCHypkC2Ld0jrkcjfAm/SvIlndrNKo6Jr2qne
s3Khm7Hd9le2BDR99PhDEoB3lvG0P+a1cXLsbMULwoQ4ly2NdZXsp03g9lPlqMEY
YTGVRhwK5D0L8/6ZUlB9fM61q4HGViT5P0j485qRMWT/B2euWHA8vZdG6AlcyJMj
rgPLMdCg2smCyzQCW1QoincPxywhBOLjxsxOYVXlGwRTyYLjfpj1wUQz0OsDFB1V
dKpbZNO/gYH9mMPAjFM5TNSsJbi8EfmNKjevphaeGuY5q28QZmVJTMChLe86O8n/
qN+vqok1HOhU1yLiT7iJM7xXs6jQR3A+tviKpDewg5AdL8kN9vFVi7Jt2gvEf1DW
5UpLoV8EvGYhP9c9nehZK92VXNQdj2mankd0e+M/unUGbmUxve8nzd/G/Ag70pC2
Fauca2AgAyn81g+x3hTrDJmxWuPzQQFgpbKR5IugCUlr9p50ceegXDIyEvadvtQu
k5SotAW0kkimcbiD8/L10qRzzJweUVbrI4cgc2cy6NAdqBH8A5PAVhTm34Xe0sAb
v2QcfTxzfdAJ3SwpcXZwoC4BbPoVKTHWpY+wxwEIFHrO9XotWkOVFZueXWKaPCtg
rPR5WiAhDkpW259sgLSdY+m2y8VuvBHrAvrxSxpC71GSPMVWUAeIMyOytGut/xAZ
B7Gu32ztVpKzoRvKIlFR+i8ynJ7j+dkUDcsdWvjohJxQ0ZtfHwsk8s6Hp0iKx80K
xuuSiKuNMoVCF2AYd8mi+D7PqsIvFHh2croBbvmdAYD7vqhaIe6lYB6kMKhKYJ2/
RgpUS+tKFe+6dzDhePpJL1F1thXk9N5MVDnL21b/pbyxG2VjeEf3p51+ScNrtAX4
mdjDsnT46bnug1oOGLHSbuLvYNGZd8bDZLDphiWiZOdKwdnKn/knNemNgd7CFUpf
NJ6YjVWHWP6q+4W9IqA9hZvl7qbgnZGXTxsO/2KQ34izP++k6wWrgRgc1ka0RRU3
UEIGAo15syo0oBMkxSVGfOfDS8TSkG69pMNKjB87JHgUqNordNWKvcn/QzoKIq5T
xLmaw2tlKC4QfxP+uehTHRi2CP/4pBX78h3rHc9cOvK5KBNRYxKqc9+iHUFiFwTf
bQTQHp+O5v1mrPjI7e0LsJnRUF0rkCMosltA0tV37MPLrzFol3hnxfBCpymKUeYX
Bi5OGEckfwPRuO4fLZ7A4zoY9AjnWC46dQW8OALGXgTcX6jhZ+dRZXL1205Cu/JU
22663hqvg4q/4ibZHi8b1ftXcrEB5IdEZDUGpywhJkgwCZcGlXVarpGIbvS1W/4a
9M0Gly5O+4/Qxyw+BFjCcQ6PVZ+JOlHsrxOCuHbFT7nLJxK44HnMQ8VS7lq1xNrH
TsSoIanb0W7dgXETo65QtUJU/8ZjBYtie6zL/tNKyh5hCsoMMpEC0s9CXwAh5RRd
4jFPgtrpeIK4JzCEf0/MpGmHw1efi4pU7hgv4lLyLxnBgkIaNfPqQ1kjGWZgrT2M
fE76CE4rRJYo+o9vM/gDol2pbFq6NQx0J31gNfIvCoYdVvPaGzVc3lTnk8jnc0BS
WiM+5N8/STpvfHrn7T3JqsDmH/dlB6z8v0UYmwbafxtS3WInX89ZLymaAUusVWyK
l/oCrmz7Henpez4MTqHpY+rgNVjqEfKCdjtf0p/pUGVcTqy42Kl7WbcFBAJPAT05
NMWMX5dgS8YPvnVqyOTgUJ1j7K2OHnJz9lc/FAJe31lBclTURStUY041qHJbbf7F
gmhAcFC6IXathAhzw5XCYVvMyrFLK+z0BkubFCLRVgaIFyjdAIKyKmIA6M9U6dWx
skA9QPwap+2KtzqPl3lMgKDa5YrnMm6vKjusT8wuCyRI2B6hNnw+sQ8tvKBXn+sr
pn5oIQyOWzkbvmX/swsr6vqna8vCHH1J4s4cjyrLbYoWgjKZ9+j76z0F24u/1E8N
1cNTmp5w3uH8baV1EGtDNaYbt9svo2vl5NA6vBRHMeV8J8P7LM7rnYBKPBqWdnN4
fmYRdLRBlZac/M5lHjODNtIFZK2t1Uk0PFaJmLxKvnFtg15P12gNi+gU7s18WLTV
jhBhr+QNG6tBJ7raVlzcl0FhoNa5yooCs+okbSsBuWOx6icZdzWTA62u0bR7agd9
tJ2ghGv51rx4lZFulmwvCRMRaeDshE2c8653AIixJVQan7jCF6i5YVQN8YRhTj2X
5J0tYFS6cBH2yGRiZPEyilek6/UrQ7xfp4qEW6ZXkxq+y/Mc2mTicrEBIFV0Xz69
e6BlU+vkDNrovTGMg8OmQH27mVNGXP+UQo15yDt4FYq5Lw+YNQ9mAgs5Ha6msYUG
72LqRtNh90BeBScZUpBbb2Fi9CIf4ngt5kq4yYfWiie0anbjggVFv5nG3zg1ySlr
+9AOk1bAFzwaGjOLiGFSj6PQyiXLpg/j5O5ZjxzxTbVE8VtV+vkHtQLj+B2XcAcf
s/1P1GdHarHSB1Sc5z6mi7UmpqL8Xl8PeVaJmXWayzfzzjulj2MB5/Ri3MXq82YE
HzsY2dIqThiaZBdXjABLhSDPYvVlZ9/u17A/raeDVbQNE5Zd0OWY4yFtZY2YRMx9
HwcagQegUqpi45BvWa0Fx7wxBh7WVtk72pX/U8Ljw3dP1UAnCy7KK6p8CqPVKV0K
sclNo8/buKrtGFCs/ctf/q+LeraH/oWNZdg2vt15uu5skYA3TkGCfaiODrzCDuj1
ZDtmOqk8oHRzT3dV2ACBQc+dAVZu7Apdz+xAASX6nwvJLSxQPha/wW+h3o2VjkUz
1a1y8EvEARUtHTD5OjOXzZNKnyPzNBX0pGspRQTeHpWPQii16sspvw8E9wVlL3sm
ZjaTXtuxGs7Au6tDawxlx94H0r1JyZE0Q1bK3hsfdapLpmIL03A2Kr28QPZTT5wj
TpU2pGFat12fHDz16SXcdhdqstu4yJFIRPHCBfMTVBSQAr2FydsSa/nFiB1SpXIj
yeQ5ZQQwsCkDnd+9CLEpHtLsS18OTTtMYaiPHcu+Sw6zWLKnoo4+dv11oXi6GeXB
Skq3GVa2eMlXVTxoRtmLeO2aE2mSUF9cHh4NntbS78dmGmlIRRYvFgrsuY0Tj0cp
q8Dm6P0OLeUX9LLm1HI2dY23cCMGluapG91QeHJtnhw04fAiCtMcCPtp5QYhiYAX
Q+SmFw0MoocTwGzWEp71IcHtn2Js/ccesFNqz3QIGd9qKYpiwWg256+6aGU9Y6/+
hvhitdN47GP7dXSW4At9V9AA5Cobedx3uNEHAR0XQCt8ysFpJZ4zKnEEZQGUyXHB
sLvqgQTSqaOzf25uebbHUs4c2F8A1y3HjHM8/tifS+JkCUDaZeu/m2UDGSRIaOjn
iMM/JH3fXt0dAx9JuOKMA7dvAPRx9Puk7pg+Df27mAr7AtFPbXmqG83S8Y4QSXdv
hn20prIxjITF3qFdBBBckNedaOD9wCld4N1OXCVE6fbV+asDpct/C5cPNe0E8CJq
pJJNHPAJniaKhyTMEaSyMVzBh44kyjrJtjSocX4UUbGcbufIBJRh+MxmVgs0kzxT
YWZ+g73l/9/f9JlW/HKVULKFSbfanLD1lweBM5VU3+To906JEBEHkolcVtyngO6P
dX4LE4BaicHpzOcEHdhBifGac1uNp6eaiiZI6vNmzDYzfszOy76AJzPzw3i4zlgb
vegrTkkqBDDod1ABIlkxl6cV6aLwhihxSNYKkBNowAkzHjzOzRKLRXXM9GkduLWs
MEF88fQ1BVIWjSFN9v8DBOtFs5JutrIof0cuknY91w9ItasgBtI8Ymgz68ISDKdJ
1Orv6JtXjP+XV1dI/J6h5kEr2OH7VX5jqBPYevOv3UJlVh/cpyJEAyedgknnVZyw
noOSnw0uyNQoqa+HOO0qJnLhq0gdXa8RlF9H9jIJFk7ObedqhyW3jjUoKaFNmNzH
Pwj7zfzvsVcqzeG6nwaTZOX0S3GLRRrILF/6wOdHUUib3uSyRC7LQLXJ6WUxgV5u
D/pwWhPvneUrpM9D01TMUaw8GVSNQaCsqnNQDhs4llrP46h7oEGrPd5uQLqAwOPX
IFOQcL2MapmJs+mt0YXSN2Oh1eEVgFBtX042UGLdYyJx/Qa0xws+jJwWpilJqino
Jl3yPC+8J3pkkPMEJ3N8rQ38fo26ZRElwRmUfEjUejBU/xAEjvQOpnuWxFxcV0XY
bgDf0ybFCJV6xbYRUrTCHL5sRmkmSx7B05EOjx1IXi8PTtB37RIW2Rw5ooqKRRDL
z27jKPNCjjlfpHoIo7SUgYrtnzp/P2T3KxqjyuNkzf22xg1Zq69YMFAEWSzro1Me
AQ9lq14fYZtq9Ctgd98FuPILeSUMCo1X3LuegoKZSw6vss0eaM1kl3aP7jyYHdXX
00Rcx/9Uhu87sMLdon4yny1ldgDrZiLDKy5xcTAXEoa3Nv1DmTCc4XeXkb+RPUQ4
Smb90lMYfCSMApTUO1YE8tZP8CP79yj/rgllFbDGmX8XV08Z5moFo9RhtDbxu2mp
/HevEoqVp+koQANKwaiwOayJRiBV/3Cw7pK9ZqkSocnq7UAXhJIEMVB6m4MlQ7kw
3fBvWRmQkFni+PlLNrYaEglj99Tqm0ppkFR6SSOZbcjLnsnqq+XAgTtwGjUUbS6Z
nBIzlD/eOLAJYIwd5LUzoJR8VL0lMe2Lgf94ZhNAVTTtoEi18ynXgYCOSsqWUV+k
T8f2v1iz4eNBVDtii5TWeLRJn59Q+MBdIQcMHzyNiwiY30/Bs71K9NgDoRE8lIQk
hCBh7GqyM+LdVW/PpCAaKf9dqmHAtqKFamcm8DuSDsaQYgPjuTyYdbs829O/z8dQ
SoQF81qu+z+Z6cOperkSnmgsa1JYgymh/kSnxIMqDUp5n1Ym35c8iaDOc0p3S69h
Kw/F9FHWsD1n62+mDfbQvwroFT1cMz6ZMqpqF3lfZ72NdLDUxtGWRfaGCg1HRTQj
n5j8cYaHwQQNOknnluKbhePPx2LzLZNsWcXmxQKvrqf/YKNYrSO+sdXeQqp4xK3o
kGse+jlWo2V48dkaHhmajbuuJQX/trI6gUoDK0ltv7ALDpxzIn+J+/dEznsTgah4
kFk9vQk9SSVE5uaB21IPeLbVwuZDJLczcRmAJkO2lGFVkBKvnWIwbxJFKsrh3hM6
6ABT85uV22a5GgWpyUEQ7DTw9aGIxcfj1f4NKvPWGp9jP+rDyXMg5YzjgItkpvcD
23CTpBtSMhNbR64v8UF53efCuaC9got3L1HGLLkt/Su72xHm1EDsyPrtTZUqm4++
ZguWvkTe4SnSnK0mp/wCPnQ6MXCiuspbFlQHfRzgaz2JDmUW1MduRp22vyw7yuwA
PFKbIrBYOa1wVeNFZ71YJ8qPbaY1hYttBzJmQvXLOO4A6YPjL2sLg4hiV3vpmjLx
HQw/ebajIiDGTO7PJTQkOuHtwSa0WrfKdi3t6qhSYZh0m7Gpb1CnT/VDGehmLSuY
hnRZ8e+152u/hId1C7NZrfcF4MJEcWndS3GdJbCVFty4c6ks8GmnbLK8rse9TMMh
V+oTd9NCtCG+yfKucBTTdzScG4/iSsxsRnmTi22ctKHB/JZV0vmArj5aFfeZnrqK
HUp2oLQGR9DmWKSxUbyiq6zXkB84dlWFWNRO+mKH9Qf6Mb9tw8qTXDc63m1UtlZ7
v0tNEUqQ3Yiw6crJSncll4brwiJ5wQ7gIfT9gv+w4UB/YqAFBTskm/dTXTW6iabg
Y8MjoqmvpYeG2wQerHii+Ou6LWWOj3RNohGqxV7/7qTduVBPzxna0ffgS4tniMB0
wB4d1/UJBitZGWH0xRbVO0Je+d8LdytyalY6sB8egJFkOZc1bE3Nb0GPo3cesXBg
VLV+xnrZkrJXTrzsq/31nkoTReLHT2KChrqWsf3HKxuvcme4KWifjXkRECV7DpPe
ei7l04nYBQno+e+ZfNKp/mDt8Tz6nT/vgry3Mh6xmcCr2vEqrGCZWUm7Qq/dPylf
tSbOlnMNcYiHDzBwIe33TqLNhttVScJ3d/BQN55lB8zogYlpnbjZd0ibgzhdqagC
7VAro/OOjYN35WgXyf6XWpDUjdtJfYETNIblHhafgfPBhtW1jZaYKj0nByR1IGKj
++ztXQi2b7rsFz1QoOurvgdhsuxx11JNM//38QttRlbx4BQCbt77mNKtAY0qxMTB
/C7OjSULISTGeuu0yjX5nv0tAF3usAcqZNyuvq2u+Vsz4U5r1FWGuSA8srXNlEdI
TWHDFzB6afDBlhGnq5tQ8EZOBZNgGeHC9oxvPmhJNGny7Y4UY1qQ3lvNo4VCfKeR
uvdu+ZU5x4T4y0HHU+ICAhnBJTzPJ3f9B/7GrS1wvwcIyEJHGehMnnO7kcA0YxQx
j6nvrmmxe8d5Ube2o+cGvWWwFFhEtdp2uHUTKhEFajTC/KwQ4DEOjQdW+yZWJglA
lwZIwfd5SgnvRN4eMBN7LZiqAMFjyOgxzCvM7rlhCW5JTN6fl7hhfqf1fl/oZsTz
4uA2/dDYYOTL9im+BAgsSj6jKzV8oKYPfidtLlf5UXJtlz6kB9UySPeTNON4oUUB
nACspdvxstOj7NOR6op9Oq0YGFW4I7Mz2ytNym2hFvUdcUk6l1YoGwEB3FkRDtdj
6hTZkrdmWnEsGcypo5JdMxJUUeWbph07gv9nVv5roZMlhuuMuU3c72aLLaC33tkb
Ouz7/j2hMblAMbWJ9VCyGbCk4G34Z/FfEGmGyxOU51BODyiWtiEvvxBjwvXYkjf4
xi2EkddAm5vntMNANolXUhjQwCn5SC/R9l1+ywa59jOtCSOzgPExcovTtQxKnyqF
ZrpdaVMVatjDvdeS5ltAfS2tjMBcFVvDZ8R9G1EM4gwrynLZimY3xpHGMi4ute5s
1csXkcxdOoz4D6V+Kvn+KVwZ+bH8o/XuVLZoUDvmLslC1z3SRLubd84UY9oS/y/R
FoXXbhFd3CwaL6JHFEM4pTwGS7RYbKG1cCRPDuEVb13rUGslGMA+LOqIZysJUCjN
oGgc4rPnYB0ufks8RNv1StQ7vas7z5zfC3xZN9QIxKS36eqjQjXEr0OKMSQXvuVk
FidtkcWp+j1mjOL+yZm9NLeCSOyPbNsCaqWVYZj2IQAc6leGV+QT92agJTDmZlFv
vuaeocVmlbAItxxtUhxIlPOfKqqylp7krYFX32x12KvT1MnFqTznRvZuH2kTG75O
J4loeTzsstu25B6eRNTKu8vQu2kmnuEeEkemwMF2nbbefBo0n/xCmjSnlxvZJ3CO
YIlpwMmzHt0yEij+j8M6AOne6FL/ezDcx4RL8k02+qGf68m1CKjplNhV2rA84ZiG
uL2PBFE+qu99/EGcLlU0oLfDyo9Y0JaEatts6OY0mr1qhIT/BIsg/dtfxp3zNXcw
Uq7Wo2FY2R6bDBeSHDHo8EirwCgRUcoJaohvzDpWwK+N9tUaYepyKhz+aruL62g5
UZA6vwTROL1oBhLzmQAXj5qfFQEbCxCMkF+VbsAJQW6GTCNQxj+eWVR7Po6w8k3a
WhQ4kNRUVV+7YEVqJO7cUjSJ28n+IAJ6xy/1mSjAPbdJhm47n0lK75eMV7rCKCqS
uyfjQqvU7DgnY6m1Z5px1JyKR8xmD7rvl7l3pv6OlHKPkHHvejYmZ0ZLB79QaVdc
q0xjYWUqyD3BFKRIHZiqlEBB+KfRCguRBBnybvvCzZ8uzJcORcRQrOw/zrxkO6A6
NsonVSBZq0xRIrh7aCQyjv4OQscZb6ngCjYlb6uKRfEff11Yj1iXTtCY5YQTQCRX
RcPvB18LA1/fNMRgS12riL7WrGmhuC0RJxjsd5QzxzPGz4ZUg1dBV4eMc0Sw0Qn9
grP2rUy4F3XUQwehLO2I3LcmUApA95TH9tFVenDTTk1rvqFg7G8hOCOIRnlEFvMm
3f5ulkBEm5WERhkt1gWEkIDI8CXkzEgXTLtzSATDdIrpOyHivox/5xQnXzW7beq/
ncoMIvAUqJSRZVJBYDYhvoqbkKtZhawuoyj58OrvWV3w2S5Bou47Gq0JS2k44fmx
AVXSnDr1Ym8a+MBUN6gI8TICl8JUiKykDxbZjUqdh5KcazhTDwjER0DaOdWJFizX
XHreAaBBPSvX0cwKpJSJlk5o7b19X6K5sYUmAbWDddBwtyNe9UHDnWyFF21iJsD2
fnyP0flcSer/OWvhEj+n5rFPRrLoZ9OxMn1CRbCjP3w7ir5xVPDfPjYarE6zCtbC
crXVmmoqLUJN5at64CmYUq2sZZuZtb4dM+x20ldMjOUcIAdGiUE1xu7myA8XsRjY
RH8/HSRC5LudbV0/nIb0l+UxhN5T/SvACCqtJMmFow0LcDpw1emQcMgG1tKOqUcn
xhiOJPqGAEP44E6JsEU7MgX3ZegFPcKveLXmSS7imh5t2/Rn3iERoM15GmlMCs0i
VUsWjLR3xRZjyJvfNuzfh9BBYicxCaaLQ2dXF3fDZt1lYNm9XoQvFH12AKydwqul
ss1gn9OrM3Aw8oizn5SZkUf2vIXRzvbtCKQhcRtJff2EHrk/noJMo1Gu/u3O3mIF
uFoSivOiuwssWF9ynju2TsXiAJ4TmFRZDuvjGoJzjRsotifRKEC+xA3906XUbmlL
8IbklEQUj5pD19vTH2zg8RL8Sf5z94VEpMzj1i6BWzkVK43qkPRkpZ5XGcGICzXO
xMQT7XfEvjTc6iekgpPCKogTdY5CnlV3deWy0Tf6ZialJhm2iHKlvuTPaBe2LwfE
Ys7mstSeALYcAPcdMFQOdmTdiPyO0wIXoWShW2s+/Wux0n2MHF9XNipFkyHnHbZw
1kPVxvhOWfdueIrdwKcDFN1c/PCo0cVwhgvPRQqZ840mENMqvOFoFHP0XBsb3/Y/
F6pDYwAuAusBn/npnqRQlRuQtweEsMQb4B2fCpRj0pziYZmk1zBKOD+QjLVMB2zl
Kal2qE3jKXvmZJDcWtTYvXTNWcjUTqtM20teoqCVgwnJwTU9YOr3xfgzQ7bJpmlM
MUn05sqCNt15aJmSLVMQrByTf6folWhSDpTyOy5f5S9VTEuEGZz5vvW6tXzr+KML
bz9k6mn/nWZer74AJm7RV6C7jVGA4zH0kqeJBj7SGnQcEuwcYpOeM0J41ZCsALgL
SFEPnyxwVTRoWm7z/C7KyHoy/Eg3KgBAQ2XZX1L51K10n4bzEaYQNy9TYrNTvkus
s7IlFDFb5H67mFEgp1M2TtwrgB1sfgQlX5Bvsl3fqxnZv01kK6spY/oEx+fPq0Rh
ltbDv+/1XoM2msugzzmSV3RkSts9631oAuneWSSrV3lfNd4JRTnz012Rx5jMUxzj
E23auJ2P8tq9NpABys0S6Zcgbf2bnk0TdWTxUVen+qY7gFg0mvRGGGxR50Vymjvm
H216Thlc4uoIwgeTfRD7Nz1KD36/kH80vUU74h/HBwjRDUq2KS37HZzDJKS1CBx3
167VlC0yQ90q4wMqHqkrXBcINoJdteq1ILPl2viyj0WjWDjCGCweTyYRIhC1eZBt
dIbKjeI5JxY8ZTqDZOdtXRhh4vliIVUTG3sW8S6ktsiUPS3/afYwV/wviWLL28Qh
yqqS1PSZrcAN1fstG1eTDriBJp1zudQErsWw6ygyde2eI1VdjxWL5BqluhxhQNRv
kdNrgDfjiCox0UoDSsyZ+6Kyz5sSr9hc/NxQd8uGL54vC/k2Ws8mvwjIgfkrjp05
RF+Fa+GopdIpIbCwTvcrY6ISo1TNy7FjeN81C41OA6J1vG+IR/icg0ZjYdR4ZG1i
JkNFuWig5HedppYyok5ykyHL8cnestojSP0EKL6QNjICEb0/yGByLEjJEdfVUPJH
v9XQe3V1cMUZgxh3LOd42WJJmnqzMbFrV8nxnqj1fX5/18dFDK/1Gf+q4l05IFc1
G9YweBiG+7u0cauDQDj5q5K+euOCK6zyrM9O5k1tw6i/iwULrLSMV64Ml9CNM9ku
GukboOX+S8ystDviJCmGHZJL1cl8XndGRZoJrGiyL35iNtfxIFn72M08GfgBjIaX
UpjTQmy/PF36eMbRrwHG43KSBsGWhRYz46vWpDCTpUyirEZW3PGfA/sIptqZ1aHO
CzUAEMQld1pvNICsW8wuNwSyCMTZ2hg/KO/kTG2jfRTBvFIUwY8oCCN96d2ItK29
yn3sqCjgG3uE0C2jNpgzXnuAytZWg/bHOWIRY1B+sGcEYjbmyiSy7o9QzHwTqqvB
7aGS23I2WT6sqKJ1xFb1F2Fs4cu/u8xQS/lD3LM6ArfPjUS9CVki2A0I7WuA4QJq
fIhDX9vl0XtM0D+U9FkvsE4LadF9d8m3r8SgRvM7ouEEfWk8MwX/uQupwTNHY5WC
jY6QCCdukay+fNsVbbXqFSanmOhhd5ijHSxJ2qQFNwTY8ZTwgT0NhKQnlyLXjEpw
pemI+ABGxgVLkQ9b7iis2neLi6q4jtA51VhafWo0lqullaZpzBf/AQSR++Xyh6/o
n0W68J7gc0z4zBxYGHDA/7uD87gOaV7gQZ5axbeqa5INUiOEHShOIOFsPN0p+yOK
MAX3TvfQ927pJiZ0oej5wFw08x7DTrXspfsZrYj4C0WXNlJS0VFgPNmE+NLtQmUV
zlLiH+pQpHYRnXpDzLLq17wdHN61XbISdUyxYXg5YVA0lUoM1SRCmaJPouT9wjEa
sYXvg4mJlSz4cXyj5MTFpyOZQI+QX7SeT5RlX8iSauqcS7qCq4p2g6jaVuPZWzUz
u59qU0vwEd/3abJtdh+PYaihn5v9p+c/xEogFI3Kkh7hEX0qXfWr3gLo3CN7S6lu
B2LrZHt+MYErkJb4gmKCfPC45/2bYGRPxz1pvz6ep/GleBZRPF1dzgdNysDWURFH
3OmCro0FKugxL1c1HXiok++CV3tCv5k4q10C+S5UypHZxCCgTERCL1a3JZFPc0BW
iqKxPlImjOC5Tv2ozOptirnRDLboWJYOy0x2Vh2C0oRFXvn3+3FMy5Y/459eqkXq
VnGdOh31F+JCZ2eePbSfMqTh99wUKobDW4dw4USUWv1vY9XF4OAFnZPLifsUaPG9
tefUwJMC8XgsedYdiw01YIypghi4u7qnSytOlkvfG5F6dfWzY4+F3ZTWpb/KawnD
XqrEAB2xEloHmcKSzDOoS2JCgxbsHG3GK2XFyJRHtZQJ++b+E60Gp5Po/Qv0F9zR
FzHHHNpXIiZin5kBzk+1lPRUnLRC1L4u6/8U1BjpkwP66VJPznHijhbc4p8J2HEn
CFBxe/jPSDCj7o0FMaWncC68O5H+NTjX3ulaHJngMAbXzGYXvY5fRGzbBKP+AxYa
6zpVXhq/ti0qnRNW66gWWc+3Mit1myibgF41rR41pObil8bWVGp4BcGf4Ct4stFw
erDFHOV3wUVqiCImdBcZsj6p5N0r/IaYPUqJvTTHeOciNtnNMOaZ/d0yEH1WPgwX
VwDAIfIPInHgq7KuhpnfsMXfb3m3G+ZTiiywO6OcXgG1dNuWLv8N/uxx1OP+1BSp
ZQRf3ksXrNJ6/uBuHEL0wvjPaa+JDBTWwIRXnho35NddM0hg/6Rsqxk/S5zXiYhD
ZlyHtQzqEkPr+UHjC90Cj2npu/CnCJRn2nen/98AP6urWlzoiWYYpX7ejaLIPFvW
IA1mYXEThimzklpOo3jpOCxkNJrlHNZU9PxOUpdUGrUVdK8CeuewA9A4ZrXUAJBb
7VstMsBQMmLiq9/8da1RdQf0Xl54lLCHabsO6ztZ5DprkvmQeNhi5s7MviDl0ERy
qX27Q7UlJyRtuqxOKPH9vuJ0cd9IjQitc0jBSn3Vj4MhioXEMfPit5z0oQUxaUQ5
7q4CMY+s4QWf+Cf/Uv5/B3OL+dsn9GcUGt2U0CzCOjv4Gc8tMzb1yUnm80H0m1h0
KjAeueTM4XFKdjzQRwJ2GfaEKEuv7xd7r+arcJbsnP0PC5w8DB7xU0j/Qeqe1yRS
rNLsNv/pYxqX34zmUsDOPgdSS1Y7C4mb6qxVXh/5f8/HOQGRDKYOvvPYjyXKwmZT
Tem8tsYDFmyjHxxIZJrIeGg2s0fmJTNgrhMbP/knARWDabwpaeicB0VEnENvuHFy
rt+S+Qa49dP1oUw1f8dfB6wXLHj+2Slv4N/hxtOmKnYhmCOERtSOZ58ngoby/lbF
Xgsl2il8OY6uxOrpUIdeN5ijscVN5u5SM8cctwcuGgkdKzK1l3qOE0cDVy8JJCxk
kT/b9Sr/0m3YDC9pMXn5AD41uvNPrbAaYHEO9VaVdmRSqQMrRwzfe4lG93/P1QaA
KVXNPj/9moc6ydfFemRdv1aAZdRCKB2u6z+ZuKvedUN+h46/66M8XdUbGPt0oBmt
wd1JDpgVzCfkUSxH/mKsgnFPrPiwYQERRiI8LXUJvgPnWfnPPlNUrNUAtGltZSsr
+De5/iisYdTVvHkd8rPZ7uXyBL1BrRQUKIVOv8uQcNyA7V/AjmeglwtgI32bHy0I
OkrrHVJR61cUk6I/Tpo71juYxpOAOZfdZFdcfeoVRiK+lTjmf+lR/afkCsTAXxmy
xH0M9MIEcFoVR7pgw7QsdyLzOnXzmzNeSTxbdrZUGe+/0JoxQeggAH/iOADzqNg8
V6YYizMsoeSnVV6v1KLl8ynHkWrT0SyS+a0kI7jZqkAnSZd0niNo3vxju3aHLzE0
i9hOGEV1pKRA8jq38hReqXJi7/DvbsHchc8i1sLQm19P+pViIClx4uMTBv+tHl5X
mt7r9VV/L0Tx0sWnVFiGR5os5kgDBCbpQr8BQoBkkmKo2NE2n76LwlHgGva4eVwO
sNrl104Sw8BDPDNs9KcAp5p5jWGBgYFktlRya8crmZUmUIQiwtngBrau5u4FoeG+
JaK9686jpm0QwdByjcSi14nTwof/77moD9NB9TUxV5oeVfOX9fr9/T8SyPNG18/8
f2os+VacZ5TynjT0pz/9EtrMU+9p9CNa7/NV1wFbdVhO1YERoMnAi8BUgmKf3Tsn
ZbiQE32ZM87jQ7KETj+ld/xTrs/LsQemoCq7qbIPZs6Isc2/XfVFnVYIuL1eRHzy
Pyn5MnSPYU47ZXUXQQCefyfyBONmmg3iwbI2MnaS8N6xpNPHu3aaYcMCY1KPzaXE
CrymmDl4Tn9H98T9i9jHn8dk4NYN4jIBBKT7VaP00gEGFFgkbGBi++IQL6YJ5zo9
05xo9fx+jQ5yxW1cesmnNk6xwmbXgjBwcWhQdDoeG45AUpWeZZ/So3HDKsHsoFPr
YOFxQjtIklb67QJRkYLzvys4Qe2iZxYrvsqJmZ9VmrWNQwJ0cjh6NzSjCXOoPCoV
qJ2uMEOazyeuq5Bf3fCxbEUYEmEqbZ+miUA5DfO897+Trw8rBOcdgobAMdiviWuC
XVAqeNlKLWJ+C2lspPON29V13vl8b5947BUdo0moiEmSC2gtf19wG5AYMC54Nu0x
I4dTf/dV71PQjPeVcKcqo3Ajuu7RGRBe9qabjmsETrZChsHTpai7jitFArQBwnrl
jnMaaHrCbC/mymLmQVMijx+9HZTVUTWFcN5HCtOCQgK9A9wCbjK/C7/yTtp0hS/8
LnBJ9aRUGAuovUA7l32ql3yLYMKmjVFEV6PfAvQKSYDOfq/16SMKS86VtllaI7YY
NTlrAbLo1eXgphlw8V5JnuLfOCKv6eNeH5UrkJev4urepM3nh4kZKfe+X4pGEOl2
r+kAQWlv9c2Ffnx2YoWSD1X+S3m2rzDhAApAPT7+l5RE1QhIl2xYOSuJ/YfGB2zY
2Fwqf2YLyUfA6/RVpircUGCP8yD8UZM7LgIa8gVsw7samUSLrgTDre8l80RPGmsl
XfsOeFkO1mJHJ+bkrgxxmxsmTLh9fs5IIMvQRPHodimHReCYRgaqGzK9LSUcPJmT
SZfEv4b9au2QhhA4rMkkEkMW5PA97f+n6YZnWhBxYAkc/sXeRR3UFg0VrwUeKG/8
8opgTx1hmXYzB+1ScuMO4R3cFvPSdQoZYg+TSwjHdS+NOiFc2jC1IwFbLWC16iWd
JC3pHMPiEwifmWgkb5wW4mtR2o3YWaTJqiAPtkLmY2QgbWCxd6Yl11rHt2g0pUJv
EFR3nBpuVeqHLwEzWmrAz0hTQUJ0bGjnEFHv9PAjQmp5zaRy3RSwabVCVmintXao
zOHMdBliDtVld2n4n+gZNNBbqHfd+tNS7uGwGVLMwZDHJBk/yu/ECY6yyQQ7Q4/M
GmyN58NYvfMcQQVnvHzWeNdr0t3Gb2JQ3b/8jKzbXP4bT/knFl9ceCHFnaMGiY7S
gveTpxweh3t/WPHtWU2DOzzTovkt59viqPWV2fEOFAj7EJtuHdTzhSWxr195TzUR
I5VRiizseg/jDwB/k9Duf3kfr9mnIuq6AEwxHSkud8JThUG8U5t2JeYxHwoKYtYQ
CX9xZop+1fTvi/BnSfij3ATdQ6ji3kXcrPJfc0U96ixcXTQP7usO3FaEz6wTzQkp
44bmND4pOuAcVJoVs3blerZS7wvxXrYpoVdql5lYImR0vqTxVd/86uf/+GaiYm88
wZi0ME+Rdo/X8bu5tFAB2ZqLnFLVN5ipJlKZOn6pbEOlGYnvCAnvBvSGkclzbBI4
LPiEKRnu0dpyNfzhQFsxVWni3UN8EyZN2r1NsQR0W0/miYDfJMJ/XZ4ZXhL4Z/GP
TBXMc13x9bRdiWv5t/jFLZWmCU58Fpe2gwYehJEVdcnL+ij8+tptialm6o3oUyjp
QQQrQMyOSq5Bje6hcI+8tLafD6aUeli/lhZevq5zun9BFo1eF/62mYb4PmjKeWFr
NpccP1SqOYHBSK4TlM6JqkmxBwkgcffuzyqwp5itFjB+KdDW6oFLgbHOVKOO7umb
+ACT8d9x/eJNY+O2/pUdaksY1Fedvk+Iv1axku/jjLL57nNs4ZvM9qnJUbmOYxYR
gki1rTFC8aXZtpl3kzWilpSvk9mjeWVQMl+P4XCAisRR4KJWlhKNbQOSdlP+JKrc
bvio2tmExRBd5NvZ3vlUR3pSowJFoT+fHSKvOJgWmme9QNKGGO8Rp/5KekHmztHz
J/YNZ6fKrXGaTty4cEekubYPox+3mQNBgWugzGdr6kFja7bmJNVnky1U6jZ73ddM
QmDp25sSBZH92YvMMuNjU6l2gRVqRa92uHEd7HIzgeleHF0TK+fO+ax1eg/2uvGw
a0XJfKYSO9zjeMmtznnEOa1bDNbN0WXZ+W4z2onc6o8Vg5RvGkIskE/f6DFhLdqk
rAUgELwP5fbz2Cpd5KuO3DqpE0VvCyZ9F8EPYndV0WOzaS4zTWg9RX3YwSgd+s2N
n1Dm8hx7spHb7RoiWVtfHxvxgRbNw4oEMenTfvDxvrr8fUAgyKilWbp8Q2YJgvqo
OWYUgcCDgc4egLvFnHQeQQ1pLkUegXiHXsyqqhKHzakCpxGkdO0xGKdgNKZSbm0W
sq6Xdan9Low8tAuj2z0hyMQPPprH0j9kWOaYoUPiwLJSR46EPwkNCzdv+6DPlQSq
10KwEGlMpTvJKjAtsbK9I43JYUt1Z6i2QU9ZvpiBk3ryTMv6QY40i30UR3LFCyVc
hD6gfYsxWvDovkMBl12TOFKtCxfX27BtU/DLQmAOs2luVjft+kZongjvtX2wHlNx
vKKlPDdk0tFhLzdz6f0kqpt4DAINlPS4xJKg181a+46ylV8HD+R5IHFq9GXm3yon
kPWG29bpB2YlL3ObrYLRmmPSPnHrNBHC2n7ajE0rhpCByHyNoT4GyR/XR60jUfSO
fMkk3mWypF2ghvo77P2EmQGIdRYFFm1/4oLCYohA4NOruYdak5Gxshm1VojH/DrI
SV1hk0m1LDgvA38V64BaBIg7T9+QiJvKRrDPrhjgeOVfFB5lyyJqRYLyobgi+oGL
rnstdS+3N8jbm7cD1nBk2KkxsTnDpL3KvxAE7Fs7aT/mhXNhP2tODS0aolH0VMUw
Ul/ICtFZjXrGCw2ieRiC49WhjTaVNPJ8umut8KBHXpFHomjRikZYyeWn0PEqnrzL
oCWCa6Ji5IEXYj/NMMp9tQfyv0UuvRjE8earzxIqMqjAudXpydQnCWEJ1FvtJdbs
h+ssforSvi/esRJuXglrss78xc70NLVyX+J8lSfBtEKYasKLTIzDLoEz7//F9LIZ
20yktK/n/0yYahdfy5FbVSw3jzn8EOcWtIsG+reQpsPzufxmIBzBalS5eF/cjWfF
XkEnFG+8kiP/nfoYpaxeSOjQREIQvnIRUODoxhJ9gQL22jdaKDszU0gSzpKjywDf
pYp0lZYaS5TNJALq7XJpFX4ldqrq598HzF1RbdfI1A7vEb1dkbNvX4ksJKe6BuX+
iLZtKUPCrJhtmEYIjitC31r++AfkbzlTjKo00pwiIHpq8n0i97ZGGEjnkfq39KD3
Jd1tIO097bZBfYvBRKA75DhVgER/f4qSrKJEUvTyMyV1vkCNnWv2rTsO0v8KH93f
7zmmbX90R8KTDhIm/Xc74PZHNc1LeTnwqNoHKPaBNSpwA6qyaxx+Z8lE7o2U+U/F
uvsS9yb29eA/A83SeAcsvGFm3CUnCzxv2NuGLkwUS3/qzoee6lMh3FgLKCHPvhze
8BRNg0PaEzGKbSGkQcQvMkyke+rntX56Wl7VRY31FryZIeIacbJnMiATrrMa8LuQ
AM4SK64XLfgcJs3MpjtD/UNyMZKjSSH2bVfsvTKpBoh94IosHT51/n7eWINoDUSx
vvgTls67jdkdfgOF/K7EJ8gSc5zXeBkzCAN63TYN/eBHTStaJ5vff/NdcPxp79+w
ZkbLuZTWEqy5WyHIby0FGC0lnUs2Gt9QFhCuouPDPsO2fSTvq4HutgQKKgQ6Gdb7
UdlG6wWutvUggE7rTLEUThJ+BD3gHSwdMSJTGduHW8Qi+58+KPOaxOnjoSyWFQbL
smyZY+rxdlhqZPIODsr5A0uN3tEEJY0rl74A8+z9znOFwRZFF6VrTPLv54tpqhW6
zY+sip8cao7Vx9TG/DOFCNk4yRD4J4IyKy7hplQw8dBvqmCAceGHshp5sMst2gor
RbPYfERSJTXaClJqYlf8gn9F4yfrLKP3W6XMsV3IEEeK9qhK6f/v5XZu3ozYjuid
r2GDdnw8qYQGBIcOs5QD37/1B/MqOiSCkpHg9+xuvk2+P8Hu2cl6nYLwsL8/lar0
n72HoKg2clDtGubGe+jVx41ScMMUowqp7/WXBsiDRFDkDqIidnISSPbcoc8+Yusa
OfRLFe+z0xoaeBPsBKwyjsxHyniaWiwoL6eL7UY14DWecj/uHpDgYGJzO4+dr1Qm
BIiiUy+LkgUo42CTXYrzObHJl54+PMd7soTbbi7Gg91AlTwC/lnfJSsIxlLfFhnU
H9orM0cLJKow2XkhODrdSGUkYs+dLbYcskbi3NWfIUGAObdviU9pElfmYYw2pCYc
O0TLqj7PC6JxnodMErU8dzISgUvrSMSJY/njtf/DFAMkfXNjrFweMFlGr9iBTtkl
WMFlFN/hxcwEiViWiT5mUbOuhKtv4ydWvXWMjlNtgHyLKD4g0tcNa1ZucvZsw+gK
3TrNW4WsbJlhP1yNN6iKuBljBLQe8Dp1ZFCRtbjIR2WhsEKX1rIgLS4tzDf6OY6f
Tr6AuqAyAVePWg/VzIniW8KqmBFtezXGEhbpwIulCftlpLcOUDvBPZUcjwtwOFnT
IMyH5EbGsCejh03ukJDW/KL+0yHaFj9+CjbBwHTFGfSq/nClXPg8GY1doNj5WGST
kbf0Dv+pcDRwH+4G/cFqUrvw19G4DjdBNZPdVjqTI9pQMhPbOdNd/i3RFdRUNwTq
kBFiM0aJCZ2VmIOpS2KInelJKEJ0gU57cj3ReYepfAxpf+L3SecpoiRb4ln6qOmS
Nklm6p26MtTu8+2Lhvu8mYV4eE4mEVIfKqfOVDTngHuGRGO5IEc1hNCBIe9hNB/Q
t3sk1ksXjqOPIHjmpnlda19R6WUrDBqQSu9JacqJTiMyR4BRgGLCCezqXrHNr89O
PfNwsgB8xtvZ7KTNsIbXJ8WzTp5qi3X+9if9z6OCN0Dw+y32bWp0/GkuHjcTO50i
kWIJmOPV/MAtGhBQ8rHVWnXP3I+W3xJaUnedAMGrd68kVQqxx6aBc/4lvArGkbmP
KECrOg6JgPRLHMJ7veyfqDZuD7cUChbOP2+XjWclAVhd+waXtDboQJydNEumnbEE
BLwuznfsFEnQFsNPTC96KZbeyPlg1g4vlLhYNEx1wWXiPhvred1d+TqgoyZpmyFD
MKqZlCvabVnE3LlKYCrwEqcf55pl0WyOQE/k64CzoRWH3QmNcoIENttc03ip6y5P
QpF/Y+OPgkbz8iNvhUunAr9DpaMiZXs1VWQew/031KpG3h8Ol96x3xtW2G8sYRzC
kuH+bBWfelAjKo/39YSKdJ74cFRgyUuR30cz4qESxUn1HJ3vb1aIP8lfjoHTo6gZ
fnNkvKXQG+j/nYs5U1xReiyAF06h0JdQmQ2BAxGE6PVRTiTiXtRCCblnl4jDLSMG
afOm/IIks9Np+7MmcmcvzRkZGaH+soWcTGvOJ9sfmEnCIQToixPzcOMRkpQ4ABQJ
rfB7hxSuFwU3GeM5yDlt9K7j0RS5i14cuLIf9zRFBam2AlAsV8X5jy9WbYAtY1Jd
j3Krlih3dcr86N4Hrxyn7lHVbOnu8OLyNgl3b1G8IcDkfdGS5flX0RB7uGu9fVoG
KybXh/xwkd6VfBoKDShGWVJvDr0YI9J4DeHlwiqmKwiCTiq3yoz/2y6uBSR6W8HP
MPAxXREnLmlX7qch0LU8NjilysquqJK/+FgPhukSbE3vAw3WWRKfAatL7LH5qNQY
KFg5MOL/2Mxn9K+srx2UQdcLP6SAQPBEbhqbv9jD+FXlDNyeUltbMuOwsTR8mo8u
jdvgHJkbIBBX3WwEZ7vL0vfFY0qR0M3vRXaqvYB4HMwaNtTXDNIZBikkGF3vzcvS
8bxRwuBGr7LoGuFRHZJr/nhzNV83pnJe4RiTCMonbRb5b8V59NC0K9kw48/JeI9c
Y+HzpOW7L2Ib7VbFVvaZdPsjFnTiOzP39mq91shc4MFl1xYDJsBYKYrWs3qHrzAh
CkgsydTa4os+RTHQVv7YV+BeN9nwVZbL6q7paLGKbdNRSrD4ZmXx416QpciVbwvJ
7MDFzHSJByJaEVNlxPW2QtNtNN1U5RANMOPNjnNDFgRxXu9rt+CLR/JmIWZPnCb4
IUvdmn/ci9fbRioPQtADB4SIDhHB0hYJx/cq/4WpeD9H3S5FdL6PgmA+vn/Ts+Zh
rlp7JuWBLwMFDCD1jTo12dOdF6Mtv29HKlG+pGNDhtVL/xAZljCrR912GEWD8k0e
vIVF+yLh1z7Ahfw1u6qDwjZNT5ScgiWoVvyQaUAQS9HV+zMyIYhpsB1+8rk7KbcB
u06S/yPpa6mY7yVkaRMD/5E8zROJ5DQslMtIqP7JNAvlRV8EjewKLrIyCOzFIo0Q
J5dKES/7hW5AUjLJP9gqzWVqmlpHwWD7ACAbMYcwdrKy2qe0nXcpq8b4HKzBpKt4
HORZQ9W0rKcvEJiZHC5KS3XFduJc+RwinOlaZuWkszacADos1wOHpSSyxwXFx0uQ
WQ6etVFGiZPN16+JJ1O9FM4V0Dsq9HydsmGUrmIa2JrQKgDqP6SxtAqXwIulowyl
isSDV/bpit0Ti7TSRUqKEn2xJpTV6k74CBHYzR5ieRbbVgz7cCTn8b4TJZLuToGm
FhmCPbX7Lm4qSz5CIsOv8cycM/Dy0qH+LQF0Et4pIMfHxjBSoYHUM76KPh1BzZxT
JKvK3Dx7fWWivf15es5xzTcoPnvOUqDQd/fEbssWL620TKZndVCQ9q7AgAjuzxzO
2bthiuGGyrjHFU36+sTYYAsErmnGofpi1Fcta4MCiHMULce9TbTerZaLQRjuJKlN
v2Gn1nNu8fLLemLbod91Z/q7g4H2JcCTFoIC0l5G+Q5DJKJSxrjcEShe8ewYMM/s
Nhk65HgNGInnE/X1mGG6txayj3m65KgMqXo3TT7nAynM4089qRwkH8zJJx++oJRx
oaSGXimZAKJ7ZHYoBYAg4dtBAWog2SYz7i24sjq8/zjJs/ICKiGausMAhCuhcmTc
dJLUa68s/MbppA2WrtS0tuIL1+/tBlpXptur4WMe7dIPMmdmIdJpiUohak/O/jz4
4F7KPv3c9P1AukvoaRnFwHg/hDaT3x8IW+DTSG/WX18IG7vLkcGfGtLbauqt7AzH
kP7dciN7km9wHYIt3HooBzI5WNnWP4E4O7iTyaWclVP8jf/llBUP3prryI60frYn
f+0Ytk4GnmRQuTFFmeDBz1D4ITLsdeaX1/m1aBTnbrIlrUjDUoUVbFvaRCr3rEMW
2IWUqHx6VDkKbEevSwbrNdJQSiKAT3f8HmLeXe9jiBXRPeGRS/9TGt/XlG6VJklf
bWSDQJ+AhrtNzorBdj4t5T6SNHBWgGGk4IOqFhR3ziGIzbgMPFfewhIHqIozhVHF
MxxJzbE1jt5BCunDOq/sT0oeEqea+CDJjtCX8L1FxNoUzYhBLxhB7dWoFt0eydTP
R0aOEkjjXbAhOBgO5lSNp3D0ptz+25JB4q34iAL/ONrUr50eiMNAIuVZ7IB9dgRj
kgwW3e7iz31xyR5aMeCYQ4AlpEU0QEWYPyNZ5sA/4gIK+5D4RZaNqJmsMe7MRCYM
VEodtoUPwI471kzNu5CmywH0qOa3DlofzYqEkJISVP+6WQfe5Vy7O8AxBJdUM7A+
EOsE7i7b9ac4VVuCCCFcAv+osxl0b5SXrrupoeli9PsbrMmDGbr7drS0pyzkB8oK
ovQAQ83zLiinLsjjemEIhtcH6upfk51RiVPf5VmNEt/vw2Ka0ENt/6Vs65k5iPS2
PZ6rLxOr2+UpwBfL+W2tiGWCwMq97bU7V11TPGxhHRXrijS+aJ9PBfPLtnGzdtfG
oqjlL6Ftf+aCF+4a8B6xXGIkiWHVP4ujA39U0PIgP2ISJqylDAPlaDx39ugN+wd/
N6RDN2D0NjLkt760TxAmuHerg14ogan67pb4fLWW5iPENf+Wmatl3vIJb29Fo308
WBx8+7R/J76zdysOr8aWoQLd6DQ8Z+1qX5NHpzZ3nJ49harTM4KiVavZKzF3ZRyp
prD/W/H+ItsttyOMXyZopc2nvK7lvRAfPaPSeVHkWTGtAKaiIzNpSOd4SwzLVSgR
o6Ju9d+jEaooVeuL780PkaBQnygaUmX2noN3Cl+isRuU4RLyN+USXmua/nnS6qnD
P5r5Yfgt3Ba4D3Mf/uf+BeHk4gUOkI5hFWZZHq1HJQu/gu4d8IUDLrjluY0uEDFz
KC0SgPlU4bFBaXqmfyjaQ2XcN4HDieRwibsT19IFOBTd3ktAvbRxllg9HQf7BLBP
7aifHNusmMThoRjxhQLoZTKLeuciqFWDlTz2/qNR87iU4cST3hVyt7W1gKKIlwsU
zwgtq0AgD2lrp6ikOIBxP+wze3qMB3ioGGtx9uZBkdlQgcpJjUqXP9GMoOgOZrou
nF6m7j4cTYo2sObfvDGlhFKHnjk7Rk4m/ztPczkEAOsX/hmEF/6YMN0nwXYs7i2s
BguTGt1sBEuBBuWF+L/TfTjIQ0e3rdMRMnTPFp5X6dOlrPc8Ies0OkjlsHQNjeiI
rormJ5K7g1FMjKv5RmVBZiSkDMpfGLOjE2yWfpyQh+Nb26frKHuKdX17/HaXeYgm
kW/oGZLmxT+YROp1fjvpyTy38FZQQId47PoW0vn2FeitekilMocyXkIgeLtSSRYo
BPYfZC0tRulIP8GgnVzeFww7/WM5+Wd5lcbx1ke9IzBjqTpmNK0lN94J5yoFywOX
n+t7iFyBVVJjhZuZ/mO1a74wQdN7Ka+MtPRCYOCSAoh+GQZbN4EAC2A9jDQwLXEC
8f3gDdz7eNtyD1cx828DKzBI1NoXkyAz4H6qRpij6LNjkmZWd/0rg6EOA+BO8pnB
6HFKaOevsSLIaVr6YJsz8T5xRmrnencByielB0Hkh+DlCKJpKhIXp0hTpjmOwlGY
gr8Qja0YTI9k8aMHU7dLEsPdjTBBWfpbVc414vqEUlN57jPIyR0DkI2TpvXSq8tg
T0SZJLWV3irgcXnUMhaIpI5oiHoOJqqKzgvnUWPvSK+s/FnATT+nUtvDsf9zDQMi
lCOLjh8mNDUaQzVxzAEHyX1zVhMcKj0ELrDNPPNCay0K7ZkECOI0huZT2KS0bXRw
mhYirk7eCfKaCqd9siXndNzhyAbDZQf0l5EwEob4IGX0RLC+q9qQc0FQgWOGJnDB
ynIzlN99acFLHSqogawKOmY+XONfcuwn2cBAHhiBgHvc6NNu0R0rodo303cpEFZK
NbZEhSyWYrQ2EYZcaZJQVb+JJwSE3XHwI2H8JBiWkZLf6R146JtrfuJH65EbdtQF
vPkS82iKe6q9LyyQ50WbpSGAwoISDy7ncCDIhNZ4KPS30I6KmhvqgROnnwkGBOfi
HVTd8Driyl/tBTaa1ICcciY2FBZtZRBAd1Om5q3PKumMWHFitqOtk0JPP0o1K5ir
6wPmsf5z7ScLMi16mlNzqrzzolXpySso3XQXgrsLMKMX4xKi/NKMpRrr+uQ6eqff
kdSVMGqxdtmgvDNmWRS7qxAZ7TC1L5CZXks+JrpM6bXH2n27XXl8rhZU9oDgxnFV
+SC5fiCJU90zn/8NasTSFe+ROJYxEN0nsdyHns/dZsISIPxa2n+eayBkgYe/6dif
HM+6Uu4PNtczcjzQHAE+dbYDdplZGP1OQ1giA4ol6njhWIQh5wpoD3RD8BjFNP+D
hRMqOo98NI57AnGdceqeb2xfKFVFj8K/FF0a2RLnEnwUDNK31PL65ozzX7J716j7
BSriRupJqGD88NHmDf1m2lr+5Bq32/hL+zosX2qHvq4fE522dMcJLBH9DoFn4K44
cSSKXnFImJUhBPJDRXZmC0u727kWM90rzqvw5TWdOk4oR/FZAuDX5EwhSc5Cx5TB
LK4/4FOHYzHaauBLXsxmQU903+C/z2Pf6WBdJwT8P0FktzuoNR30HGyh5BH3jwa9
1ojEQtfmnzN7QhCEvYH2F4U8NInHSEwkMRiNR8pK5Hc3O8LhnzwayuKKm8dk4TkY
bjpL7yVah+RGVwT/RCm0geChvHz6IwQncaGcdX3rKm/Bdhq46QOJ/H3dLzi0z964
C9NjmS7mwBiV4F07NtLVXtRXg4qWpLi7AG/voc/ZPyAmLrn2TMNeainhwc/ZW9Od
3w3Mis8VQf42k7d65hfLxPiZZgFLBvOBn4KXk87NgigEtRsVKFJTQFrtADKA0mNA
lmH/yrZoCExOv2nxbL/5+ctPYoJuzHHXolzGFdDOYu8hpKxpZuGhFSBhPSiMv8ae
uF9Qptb1IeVCdY4HVGO0WbyaXXagDRQ2u020KeL4PW0XPWvtguEKytrI/Kivkc0l
vONAVXFk8D68b5s32TnzEgSKcQlXKkCeR1fcpPRYbLo9awsiJvAnTSTN+6Dprw5/
B1h3x3fTufBwH2uLuN/ANHeGd+mpMPouiwuwx8wqo1OFNsBCxSc9HZ4qrr892raU
oJf9v1YqNP1R+RoMzHCpGuquUBICnAOV1n4+jNZWoPT2pciImsrL2EAzysSSa2ux
CquN6DdE7aPeAQsQaqHi3CaWmF+VN0CEq7mxtOuRcJbuhtMS7cja4KxCU20h/o/B
jRjrijoGn0rKBYNUyyl1Z4e+0jAjWhU+29gLG+roSaGJjXK7QZg0+OWfoG3rGiiC
wCN7We3q6pZMiEtZ36KWwxPiIe2sNBAY5JIg1DbP1eMY/8qYTeWQMh8arDmy5H/q
co2HOzq5SEJ6m/E2EnJhtdPr4ilWPbn0wgKKwotAmuC/+OizVXdqfsTejyLB7thm
09tLoKzO/R7YstZRJq1gDvxuwKF5ksxhM94CczvS2HvJzpThRUGJgivqw9pKQ2Ui
rmG8QKJBPlkbpa7ufa63LTR4c2F+xgQ5uzP+cryI+LGYZosw3GZUv/TSjz/e6tVE
XKS1ow74qWObcFjteQELPUKe/laa7/XdKDxeQnM78xCsb+J2W6LqxiFs0vVHYiW5
i39kl3JwlTXHFhvNDZ/GGRmdQoafNisPoXslEcXKXy7Ave3Q2pkW+k8MKAp1MZnx
/g/pQRTri1MEcNDYQ0F5wRufjdVcnyrazAAO+bePrIXg1Z1HP/ODQuf6aK2T27oi
8MscU19FYz25JcIAVIQkPGK0W6VA4smZcB0Nvk1hY2UOIOSGZtDA61VZgCURNA9L
kdWAnnH/6iNvkTONvfgICPRu4KBw4hPjbP5Jfud8HLKc2I1v+5dkX8ssYtfmoF3Z
cuDnzzREa16OCfOYwfD0zPrkC1AgXAX3zvz69QdrXvpY6wHVDkUz/DYTt3HW3aar
lcys1dztivsXcy01ZqLc4a0PS0DFCWNT50MgGO/iau7JmxoxRuXHg1pOQflxVm+h
ld8k4xT2rfNt5Q9Ub0BvklfnMYkV4GIkKXqAoOUguKVtET2JEoXibrfRWrzYWlSw
o6dmEfcVRubp07ptRjqnp56qf3FFzz/KySHk7yC+DKri+pzrvSL9RQhCGtsZVubQ
Zh7n7ff3FAv+M5IJVnFODuSNazfyHvQ2RP8u4Dyq1I1nYrBcU8FaKrlZL6ZwQjkf
zxpaU11FirAsWqbz6DL0g4Th7hDgNHZG6UgZg+mFxGXY3iQVyPWlJ8Y+a2AAL52w
UODdjiPwnfby2NFelYws0BMYY4oOxFISawaHIc+ngg8HPxiE/KROslbpMnmsV8jT
IjwijZwsJ+Ezrjh2tppKZ/WN9zAYuXK8SGgdrFdLcjxDD+KpVBzHJmrA1Jz1ktgu
/WFwfNEKVrCH3SvlGZSp2jWFulK8YFGj/DRT7D0/H3oEbbUSotY90QRUC4sa4y6x
cM2KrzjLZTNU/t1lDeaDMWO+pcQaCmkfg1jdILlw2/1Q6Z3AniRmEJ6VvwC0xH+s
btmdLkY91LbeZCo85Sqp7eAEuql5bgjHTliFuwIlOYQ4HhpPfSfE6mBkdRpV0AsN
VRwcpEYAVYOtCqwyxnXcdfP9C5UfvMhtdweJctEJLHKlofIIIpc4u5rMmkQO5Onx
u5ikFecm7qSfFhGfydq58EBDazNBSPtbgTP5obisgNeNjTQ5VtQP26N5ecqBf8m4
zg6g6NilgmqTFc7M07WqrqRzhK4D6zFYWJNrAkydhJtqM37vEjRMfqeq3crUWbMh
wPHGNHUBzjK/7v90lzMpd9tdPRiHwAmK5QNKqmFnjHIsyTKCtKVdUnaCCy9KyQ0O
87nmueVz78WEYiu3hgxQ6AvYNb1cfdXLnzfj+r4rrazlRK4xvKD/IFuYKa6OA3nb
JUpz9/ItzENI0wUQZu/9Qnokp7VwV91lSKYC9AuLEaF3iyFfpP1piDHEspLDXAk7
YmF95hXBXLqyyaXGVpWAPecIHw4KTeuO2u5LmBbpXMaRpy66ud/HwK3W6d5dfERJ
AbwAJAw9tOaRvOT/RH1XNMp2TG/aIT1vYSLYA74UhZsj1rVcR4KSUPhG1AgQ45ZH
g37oWO2pk+CDHni2mgpuCHEOetYoc9feENvpSc0NPpa9On8mJIlsjGg+62HgEpoJ
qT+tTyRBxmxmLkEiztU+Y17P4FoFdxfbmhQVd5NvCwp+0gjEAoEW7nCn6/+tWXut
xaLxR1cRPGl5PRavtoCA/ODDABy0JD5ZIonlCZyPxroicjb9l2cZ6zcny34dZKP6
HVYvXj1REDQzhlC48r8DPCuKgfUKew7MTibhdRSAN8fN0wUb2kUXdrJKY1btXxD6
O6qmnPgfOtH4krgTOLhnGWUYjZ+tsRZj6O1yrZbSRgKEmVX9AR0oq1wDrMtuZ1ep
4285q/2K7JlnKPJ6Bm0FwsNXV0FHUk+R3EAO1VJNPkBb6QfC1zZpWfucr2g56wqe
3Cfn7MtdXbsT+GqCjzbb1tBZKJK9oQNyv7W9gNHGyEFsUYRgteDOnbnvog1bNcHI
plbhEMaBANxJ1N9VPqTnpmOpML2eJANR9i1UmYnyIsAwBZhmPwxbjyWZytu4YOVd
zAGo+0IyGbNwoATrVRXIG3xfM/glc08U44o2tFZyuBImdtsbCBhbk8jur3PgAOfP
za+y6UhQvcL0SLHnPggXwYx6/jwCt4ze3gfqAcOifYgvMA5xedC8L8RCisNegopn
8ek7kQ5Yafnxd4B3/9XpCR4nbRCXD1SsdCnmIp/F9L7y1fwNz9ySkX81EWMeAdPC
mvZBF+dNnCsbf63ho2rjl0qGh/jcSAZUUMhF9GaSPshly01U4fTIYkWkE6a8TNUx
aXvZxc33AJlM/TxanTmaWY6dX0S9EWFguPW26hGJ087LGUEwTamcXWlYAUoMpPLr
4kcG25atzun/LayjgjCMbpdFSAbL8TbSk9/8XwyujUKo261EY/e3x+VftCTwcfIz
c6QDq5Mj7SPTu19H4w9RNDsbPRO0SVbDLDuc2OlnKubFMPFMU/B2pc3n28/ja9s4
u+r05GCGSdl1s1LVTbA40hNMBAg0ndccB5kLoesrzrrc0BlygsRurBYF9u4GAufW
VCGRfIj8+ukIoqzAnh62JJVW9/iWu0t2xWV6l83QAFJAoPLUSAXxD6S9U86dgHdd
k+ZLFRHMdr+bX7Fek+i+dPX7azQ5BydhMvXy61FBU+YSzXpsJDvA7IFmXCNpUspy
t9UBd+2W0f5xT9YtOufMtDI1IkbqpjT5B6ybzyaRwRrPJhfnAKLAcdYTpxxMoGh9
jLbCsNt01qRPsPmv7mGc4RgxUStZ7AEMR7eWTRLZ3sf55a4eMHmPAwppX80lKXMg
PpbFPIFNLYNDcy3XiXzDIBzj5BMwfJPVt4ADtIhpYNA46ptKP6zZUlwCg3Z/CnQy
gSjhSKESXwXc8dwfa11CdkI2tBbGJ7RjT4JTs1/o4BbVDDGwbL+YZGVIHEwBgH8h
rRBAsL6mKD94O62uredK5BSzKFJgW9FPu3OGKvDJ8rkv4OGB1rUmdIA5abOT7djc
gShQg+FP9gHhGSlbVxyrOU5AwClSqjvjOQpWs1/k0cgxwprk6TydkoPHNcs4GFjC
I4KDDIvZN1TgNGHe2NRc9skzYVcKtWBOvmTxv+6BNuZBk5slZzcf2JbP39Kjg3Xj
Y0We0nWQXkaHYcKgsimgQ5Tt94ZKBDP5iliEXXTYEKj9PN6gdBewrDP+2/CQZbYR
l8V01oY4B8CY6MJ8EcBLshVc8IkjZnt6Liivr/TtdOYJ3gsuQKyICFslzHfBbFAd
g78lMJqR4zSVtWXKJ0fDkd5QdM+5Bh1DzPhaG/hj8PjLS3vNoS7caW/K7KY4a8/F
bmAFuIqVzO1pPVfQyiGVYQe4BxUl6QG3cnd1LC2HqkP1NOtulAkRtXCeADUB9Y66
3Yt7TlEux5Q1/V1K1lc0FkKc9Oxr48Ccuc7pSh90Qy+968228bf2HyyH1KH8Kvd4
gGZOJW6/o4E6LcGFP5lzHkTe+asWe4x8jGvZjwADpTS+c18qV3f9TGqrwy624rcl
kJk5bQf7s88OFtHcMjxd+R6ejdswmL7ARXIaFq3h8qVaA9GaTSrTcb9Mwbuh5wYW
YBIOLZk58Q6yRuRBJht3u2H6W7+7LRPz027/7Ep8YEnFVQzk/ojcgY2FKre/CJ2S
5Rwy1P1SRCq0klTaz3iRWS+Fkd2RjOMmRVy1UdmMswwpQqCJUQ6J5y8KTzTCo5j9
18o2pNCbAB35sCdb+DrEBPSx1scmDPCwpb6vzzii09XUiYFSnndvy5B1A5VRTW/e
2LHEELg9RSe1t9UACJe2rLfTMRCgMYe/3Cbo7qD8U0o26Tegp+CoHmeMPHKP6Wky
Amnewe44Ma7vHd4ICAG2SRoMRIOrGwdNO92tHwzkCaVB74CjKWbS5JaRJ/2D9CK9
EuKVPUsUTTgW0nQRVwZhNY06M1lSYqPjgvtJ0sOgKqUmCGDH8mGvAPA0If/7OCN5
t3fUjV6z07+l1wq/CVPAJGXgFpudkF/d1TrK+m1f3HDFRMoYW3bV/FxM6ELAfgIk
qfM6Ox5CAXJAiSGd4rGvUnldDSbzGXBpxh+m98FKQGyH/wL9UIh5BJX3mrUAXFTe
kBBBHZOis3CaqKTBJd0MiSUo/4DeIFty56ui3ABkxc2JgcsI81EiXVSA6jtEVhvf
nr+KA/b54/880EUoJsx27n2FCzh60z8DOHbojJXfQUbwHehkeqa65tkYF9hkmhba
StFUisFi4ULc3R0Z5Li2q0yCgBcNerytZSaLBiC9LT4wWlcyRTdOzyLw2Yywaie4
VoKyNg3tvJf9HaZgakATkrDzhE9rUtfQByeH1pWDKyV2/oZ9h22b+5KQUFq37Wqz
dgGa61Pe4XGirNzWQMvaNmN8Q1Sbf84G92rAS78okGUJPeUGupbTWAq09uft4SuA
SuhawUtsRoOK5yYXaUh73JUx4AV4gZthX3ggHo4/Go9RMkpW3bvb36gXcsi2mZA7
0j7fH79C80bOws8w0i9SSvDCKsJyfkQptXXGxcFvNh5uRqBK0qYLPFrMtw3ywMmb
Kd2v1cTbvUizE4lUbZ7H2rHh+15d7ccS0E3kzl1HN7Q93NjEEYWaLjIQGq0XYz1g
b1th2Hi/mXVn3gu9TUL+9bI0t9q3o9HFBAEnMbd6MhBsBvs+PXj9Ad649wiGvONc
yYyQjLONI+yPHlHGlBaT2R9lp9E40uRTtyZOj0AX8vVlPmPrlR/4fuAFGpMkmn59
C8w0PvQWMG303xucw/VdWHkTo2bCjhFy35+9TrKORswblpE2nYU7JXQLhi0TJcpa
Z6EsYCCVMGjiwob262vCfp3eA0PoeagGU88pbHqi8jmd/Dthm9KRVYxBZ8D537h8
bAPEQIFEHTeJJhnuY2YaY2aUmnWrtDik+NOdUUUhZI+IFbzB/hLl1MLF/Vx/bUEZ
bpbNZ4+vBlHN0OsvayKKrbEdZUnR5onrY93YawUwbPbegTEtf0WJeuvTXUEVvbic
Ga6I19Fn+SdtsyL2Vf5V2Yvhv2skzRVRl5Ix7/ICZW/lGIzLiAacMr7qOlkcreJ1
WbjzpyR8TFkwr6/GzAmX7A9mVpOXFj926gCY3BVpb2ZjaqpQ95zVrTdpC5iyE7Xm
5xrcuRXpkpU7zXdpGaUCJbmIKBr9V3apapsgbmDLbfE9gnZLa/PqmGbzv3q6Qz0o
yexO22GfNiZQm8ERE3QIB3HAzCAw3h9LjOSTBITKDRM36aRmDIwmAcFz7Qn1B8fh
BrRab3VcGTUjv+kOuwKotwMkJ2j/DbCS2DN0qRPteSCZAeU3YHbzTdfPvKwWjbPa
EWWTfxUmcOhtZewxJ40P0toDsWyqBpmaYZcVM6537iKF87XtFfwpQ1w0RvwIu+wq
nT41T6reOEyyE+YhcEFDD/sYx8Ai797zDWRmv1eyIBD6pDewZOiKn1/4Ccj+M5nK
4zpHblfrmDkp/Wv9OXLiqsxSHZZrHxPcvg0nP3m4lw03DxFSihQ6qXSg2TaXJClH
84Uwd1SpulyCX5+JD+EyttBnlixSw6DISOptIOGkMuaGQ92W3A/HT+3N1u5lySPM
toAlc05oREInQbv2X/+nMlqI+m/OkglSeeYBDziKVW5/OZyiD4heUK3mL2oA8S6a
3bo40KKGzapa2OGTX2tgWmErsiNdNwXSMef3+h/kz2Z8ERzKYeTQ82QywINamQhX
MOgFHhIU37mUj+KWUl2fA8hcl0UfvVKIk3S0BclFRSIpULMCA6KqHKuRXypJhgeX
r6wwnnedRvaNuonN63ica2Dbl5OSGzbC2rZ9CeUtF+pxrbPJozaEZ10AajCGZONM
eecMHqL0Fq7mhSuiqcvncwFvNwi+Ru7b3W/7/jghACkLVsBOA3lhdVmGbBOFfWG4
yMnMXSqB1jqyVTNPAq27Nl4s2k9s+X/04t3O/LTN01HMHQODot2CQQbq1vrCKQfP
3TU6weMarZHjtXE5KnyEHLdOjLUxBnbvPBDy/SWA5iSQ68XMlv91ZvsB4WUXZavV
/SBBrbG+xlcyk+IOG3x3UoiDCMdr9ENmZv2eo+1Zw2I2eRLupvd9AWSRrhSFMr56
pOQZ0MQML9K4DbMulg5JVkytQRiFAKXFCY5sDrAIUJ1X3X9e29SFF8t/l6yLjGbZ
/bf5MhOc8nZsVWoLcwectgIPW+jnPsRdAsXe8CHnjNGcEWIeZRGHwYqg4GcQ8ziu
aHKO5kvfiZiPIuFciec/FGzt5RMbeDex4iqC1ZJGxRi61GgmTEUeFD86WD0UMrZ8
8GbXXsXZgu9UaAHsrRofyaijR/Lv8bYQFBJUD8HE/PYd67a30tOXBJ93vezbunqA
BZn+gGjqtdK1e0VuLRCYok/383x+jIp5itjbnsA11ad3fmg0iEb2EUFxhbMf3y0y
Fzb6fplO3j6tvN5YwEzGZOmOmy2boXw8TLZWBrIMSzsLY8eiQDSlQCYxbofK76tU
2Jd4lDUnntPH2Jts4nlNNjHv2FdHpKCPvZg9vHe5hlN8Kj/RiH/tHEI37l6ftQ+D
DuNHn7vEXOTpEozZHTTwslBgvhQyYBozUQIw804RN39Fr08y8Nl5GU99i9fElaiS
2EXXcX96BmUuVYI3w/xNlZkHcVFJoz1dxT4muNfcy5n8C8ns0ZoEFBd0093vfBUi
YhPXiq1SfoTBOBxbYb+Dmqog1anXErNf3Lkwf+fLxJHaOwCKuzqjuLtlKI/anpO0
2aJOXqySYARke5znBjwpgjD0U76lc8ozb+Um5cJpkA4evARiCqE5LJUpVycGPaXY
SKjct/Z/4gqJo+ZvDPRyiV22T9yTduUzhOLWMKyLA2OKhZYv7ju86DR9ecMOgig0
YfjIHciTWuO9/zyTN6QJCsG19gSjxetHt/3IVksfdn3J19SDeEnv5L6Ue9MyzfzV
ATK4+KEYiH3+acx0n0EVfYJf808QfSuOZ5n8FVRm1bF8wAnZF12qoVBKAry8fXUt
i51aZ1i3YZeJB7tc+JaCObQ3lBgH4OrscX20aCk7/e/Gc8xqcNWzCuo4jQqZw+Vc
SovMgIWu2PgQNDLKnY95Q7qr/J4y1WSv2OYCiekLvtIJSd0POfuW5L+o2+tEyIO3
OHJ5EOcHS9XpHgl7bSiPDBz8l/U5l43NpBKmVVQP1o7enLAScxmGhRAW8MjjqAdu
o2xC0JHokeJrXIN/z7k5U8nbChykuRacNlJmITtD3zNWwLrpMrAZwCpc3vy4OJ0w
PXvuJ4TCJcPI9xuGNPYrAI+gs3JaYnZBIpt/BelJ4xNam/JCgq4oTPk7XBstCI5P
DEfQ9NJI2uIpcro0A1PBq2keSrL70PcoabQGx/BZ+yniuGL4iBXhqU0DRyXDPvQi
g5Hg+s1kWGDHepsHmyXyfNECzZkxoDTNWGDfr0Dz3d5X4AvGpWJmi8UiET8t8zBu
JMJd4J/MpH6blFW6tO6A3p6tlf8BuDIJ8wraAN/AqWOs8q+TjN/e1DRQlyG8lDSz
gZpOgT3YGcxAP3mmrDN10m+bgZa99u6VKvTPt47KmXTyEZUFIQfC0T4gTDIOsMkR
lMXigGg00coTTaTTNvF04mi2BWVVlJKSndQOf7neq3Af1Nb7xiZLb0wR0dvj5okh
hNvcWUGjTqxO4WGKpK5B6HsWJUzUv3qkTR1zgeFB2lhQPX12xQ3ZlkNMvhZWCc89
SMkonEAYts/B4/rgDU76FXDnklehr1wAc6DL6j6aDWYmnXk2SV6HHMovIipemnxS
hsLiefEdLBjUO0XVLdkJKal7d2+aOsM4bCs9xlVIAjbXGThQq9AAdoSMIPWt9oCz
P6nUfjYut49W9PGqh/+6z2pVxvBqhJp4F2ae6hxOjZE5dE05U/gzoo9KSx8QlIbD
y5fHrY+oG9VjpicWLziSwDj/HJ6u37WVvvb5JAIPPmMg7LO2dUIhGaDM4EuS07oj
CBxnD3aZOuDLs3x+usYw+Qjc04hhKDof7TtoJiLhocLpZDOv8R9TwCk0LXjdhjYt
qr0oZXXBdXI9gaE61E63RIbdPetTj3qqrc92eKWZ6BBeImwNoqjgv/l6aDi4eFCO
Q7q8/MoYWbwjLrC6zqYLR7Ax4x12SaKS9cKy+ZuAZcWB4HigjvodtyxQhEG53iIV
hvBOEPh+/QbX/VAUC7oGt3ddfl/BmbJCmX89UnVNGexsFlw916meoUWLQjQEcsAU
yZWNxT3bnqDtDECitLanMvmPM0wNZorp1s5JZ/dKCu7r1KOaATSIEwwcXBYy7q+9
P2slNen1/tKvcQ84eKVDNt4GsQTAIiCOav8mNyuzXPXOk/mOHRCcJ+QpqjS82ICh
fHZGHDTnnJpFSb4l8OE+JWHpgLo4ObHehJxf62dfjcPwHBebIP5wcEKPBFMSq7F0
HciCj4i6XDU6DDWrLIHdhJN21iCFoF0veQTBFVB3/8U5+mvXaIBPkq9lr/Fzxqlt
dG7RkPKROdy0bsNCLx2uqYGAjV29CQTM32WagEp9brj+WBWCtYJu+2Fm+3BBKipt
Y5kffFnc0vKYMtijyEC466BE7HleI0CR2FintNyJuyiMtHVWwXRD2ZFaHUOCJe0A
5Myw8M4XVAq3tS3ZJyOB+UT3GzYWKZ2CJ/TL3Rt7sYFFqjUlfjv8fa0gYHBb2TWz
ifuM5+/tk1aNje0DacWJOprDM7QzY924FZMfiI7mtTzqDc7bAKNrLw21k9d7NSI9
nPUEoOT2TbuvFyVJ44hw1vRudW9qbPsRLPhJS8sYHsYjtzthacp5eSaA5rua8lyh
5mbLJtmvApCwn0ob6o9WD+xPddn96xUpSCGY3SBoXxevI2Ova3tkLdLaQODGLLbe
NRo0ddnAlkqtygndPMrmHD2l9wHEPQZP3jO4tUezc/nsEJkOT5Ewlvh1cS6QF5aG
g6VIhc3kYAM7fSVle6/sw7Nbe+yEAGLsYiSr1AIZ9JGPAkBtqVOo3BdthtOJyk8a
8Zb4ozpVEdEC8qwetKzp0UgYhpj+NYrf0NqQHwQG8cE88LZ9cMS9hbbSYT69I7ZE
uwRO2EotKp1u4KotG9IFj9gRvRhKcuxIqLwo9qiO0ZG7mEpDTs8qSEVF3oo0Fpru
BA8jmNO+EDx1bl9t6k+yfQdYyS/YKS5YrN6/TR+XThczGcJpaNSD64z9Bt8f4cXG
umIjkuE2Jg0dpvh4ZaSkC5LVbfymuozX/yFHuNFR08SrQv4UFZAX2LM/2jjdxN56
lYRTE8S66q0dksuQxmtvhs8LOtK2ZfkA/EHIQC2tdf/IGrwN+OQi8swf6u4Xv4PT
nuoMhIoeP6Elacg4IfVcNw/yIum9OKBy74hNHb6dhsnEPTwEfIpCENNY/sTVu60d
ehQj8rQl8owQCSVrIfJhh+wA0qcbxkRiedrUy3q6QOpZandJbhMcfA69PjOaWSWl
gi2Q1dYve1oHmxVtxPr4tz8g1o9k4nx3dSjkS16G7ZAkvR9Rx9kfgEcPUdSh4pO9
dJtvDfJ68DLv20u7JT7gu3/6LNakmb8zVEzAeZbUbermaBCB66TMMakwWSSU2PlR
eVKe5vZwObRwUa2rcFyWwYYGqH3U9NViYKkQFVHpzjgv+2a+DeM8pNsI/50BAif7
1C4UCXL+JWW+8QX7Fudma3lOQVfrkIE6Y55n+EBuVuAwYhf1fgIHyioKquT3wXWx
CkbCFdnDXdGlngagi+/4DwucEQfLCc5kEe4AtUo5aCBO4CSjkxFJAWE0M0Z/WQ2p
dcaTAdC1xNDJFx4HbGuCfTFiyrqg1U0mu3YB50qcER6Y+KhS9e/DiDbQ+V2jr2fG
csOZNdL7HE0+JRYQDf+f0srdYCxgvJJShH7mJtp5VPDEWjrzli67T/oRs0kj4fsX
MmqPtwm7Uu8C80hgYcIQqoXQek762MixXvlswZnwMBq7qk8L3sNExyaqwrcGDd1i
hSQyCLGZspFpE85HHuxkH/ereUxsUpxbFS/XujyuLD3BVnKunhYov892bDJ3HMeq
qpELn0FxwyWv3T21wCQSK4x17bUTGJ2f+AOrHPxxFWGzwYBC1teCTw/S9nHO4wpL
mWIa1YTlWdoyKxSVbCYBiNAb8A2K1qReFx9KGs2csR4B5fK0a+fHYhXp/vYYej6G
EWhZqyNXVLqMteG0h6RC8tgpbkeJMl0ItR08PO83NJt1O3rAD7j4D55xzQDCYKU1
MwPwW9WcMcKhoB6ruoIwLWvvvHhrHPcTj/emWHPccGwb6oc2tphhP+NXd2zrhlal
gaNvsAYAaDonOCxnjhNGgYx8qZbeg8b0VwgWU8mBeJuxWD0YozAd/1E/UUtUFeP5
4/WKtVViXqUEbdmyTA4n+BVh8FR924fTSg+qszePe1sSOVs5C8gLOJvK337rNKiT
reSCU9elUWAWt00AEe+sAZYZ7qREsBVw3tRimyXWqV6/fVwqzSCvUxETHH/z4wCy
wS7XUMQijH+Z3t48Ph+A4lVa2ORsvtFmzd8bWbuzYND8v0aQ+mQHva2FwPzkmeIH
Ih08b1cSaQ0qqZC/fl1NdWEwC8IYSfx2EAYtGHQQqC8UXx+53VqGLJyDN/IJTpT1
lBqr2Ii8I257cY9P2sz9zPzT1NMoyyMcuRRjoDT8sGXfiGciMgMIFJ/173Saef7T
lhn1pzQSPgCRSiNrosc/nksH3+mDTu20KRqmwUeDOsXnObiXUEJOmBfdpUHazeAY
uGxJv5FTvv5j0Xd3fW34E6kq0huN3xECQODGe14EuxnwX/0odhxMOjlv8KAe2uVD
UDM8j+5ST+hR3YRuQeeKOAp5ChX2kXjwmP114xtYPtZs4OiGbK6SW3gl2kMnsYVe
W+40knTHbOuosZMlqcQISmKOiGQzuzT8HzXV5rzLddV33dvEY8xycHHJGn7CkCnY
sIAJR08NFTyocvAk44h79HjgF7gRbg1pcQrA89QkH9kl+uIwxFyAQYLNO7sOoA0Z
yMtd5WDoOzqXber2yd9Zj4gEHmLGl3hRw57+P2p3JLko5gsjW1xq3N5/lc8Uqonv
q48r2CSA1On2TzUbXHgKVwwsJou0NPUVxkzNEGXVbh60zNquFfvfP/dYP9I6DPar
7aIHnWqvV/N5yYxKI0k07pnh/Q/E81WHGa6vobxpwueh8jGpS7R3nl7OmQpMIsWe
A9VUCAp/UqjQWomAMAj6fJiZ2F/4gY5SWdtx8MBbbWXxB4q8Ah4NlIC7LpbqMxyl
y7nw/e0tMg/X3TMHfYqbFt23DdqNh10hw8Zs57xSXbXN48IJNu1nfaQDwOIZocbQ
TQs8G+fNGs1+Pn4P40jlrfjHRQDQ+YADQSAjfcdNsEausaXJkyZ6FEPaiOZl/0jX
sqVgSJXYG/814kx/zIxE5E3ta4bYFcILdW2XueO0VlLVE4qWuaXHne40T62XTlWi
fpMBkjBwVBBPwncWgfpdIgKVeLNJwUEaGNVDGNfdQkLgH2w2y8mim9bnzjaVJ0Nv
yPAjeiJ5tWoAKAtJ1TDqM/AojzMcCLU1yaFhyDlCwve9nge19bLxRXJVPKXt3F1O
EfecQZEEXSjn2zcpByNnORSn88j6GDtZwe1WoL89ilToAmnaHGhUwSGZyw5ke/9B
H31Ri1MJCqeKEJBhhlWQVm8JSvxVVua0pu4jnxIn98XsOkVIbVwedMkKCJsYCBdm
TTWjiArwBXhQCvsF+ZcEI53oRavPn/LyitwHj02CetjFVox4dMzaD9VdnqXQNDO4
aR/i39/CFvQcU4wkE0g7Cx6My3RT8YPHvEwW3IeYt8mcvRI6+/lOGj4p3C0IoJHV
7noM45Tp/CM9jEFuRXoZ/vemaAOKSTW4co5kSs9FTxia4JEl7tmBFRqT1l+M/hfX
nOrdvfOsHl7h92qNpT41cKdqG4zTVoRGNH9L3PF1M73WY+VCeMuDqPNHMXQMjGz/
6oXnAM/9kSgIKWsssqwvwb1hQZc1tDzc+eZnsh3XMIEBEOxoi2gnMLI5aAXRvrh6
eTFDnvGFhkqGeiJoHeBkkYQ6mgAca9gAARjQFMZyQUjUcefcOhqf1iGyWFIdFtt4
fr4J+V6iYZ8tLdzxnCkbgtIoIWqOUWeeWL+jj2tNkIYo+RmKQLrN8szSk65YKVSa
DM/Uc0pY8AtiPdhlPX5DAuodWLJIVeOOOqNFHrUc3ewbELwYk7xn8XucSKOVtVVe
aUaM6zg0Gn7FuUt87FjL7QYyfokzpmajPlcK/LM6PJbeqjX1vGHlK1ZaFW6hrmA/
+LTT3pwsFBNQci5NcNHi0eHL7JgqLCrn8P+RaRtltKMXblgYHeNiG59JkKrksqU4
whMgu/OIVKW7FeulPAV/rqPMnY5xS4pEwjWn+vrFJrPf4ksIWturZ6tm1Z13pf44
f1RI/L90My2DWXNxUIzyUo90EnXZEez9ukzM4LJos+r3hiqwDGC1mJlv0AWHKhEU
2YbNin9aymanrGDR55bjwM2tJBxVzDcEmmSRwXp9R9gF690FBVXsNF+EBBPfJayq
JFqcvF4JIHvGUNq0ZzEhlid4tjvCApDEe/KlmHakEWRX8hkgrCvgJccY6AUJhF1v
801dB9HZ5KHKT0GzOPffMOz0haD2uJkYOTtUYE3ks0HxdKlRG+YBJgLLqEoTpdcU
zairk53+17Xs+awad4tJb2kOSC0oPLPks5YSf5GpTN4ZEur041pFaxG9I9gHBNZU
`protect END_PROTECTED
