`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aia48OoMePkxB1xptTnjqAhF/V77/15b1VLL8m66Uz1r9mgRCGA0t+9TpFIwXFPX
svJyRnSKeE9gKHIhzVjUmgGjECE1OYqJVrU4NeA478lDXi1BcfXa5YZuf6RkV5x/
DeLndRF8SKUUdfqiZ99zUYWoZPd4XoQZWa5LSbXVYSD3Uw7zav5UMP3K368DgqFd
M5WcMVL9yHxcoekOtZkGune18i9OBly5TewvaZi3BLXEHM1Cfwe4VZue0O9lYdlh
GFjapjMWA1aeskrrn1qYWIzv03G5h2tFZjgv57zdoXp3NAh0ad3MvjhpftVj+RLh
2I/isbsYMIaBL2TYNneS1Vc9xECttPGLj5d9XHDgVOnBx4VruI6jN3eixLtzW5hZ
EXCP7FWzY+igNQx1pQPkkOgH8+isTozWQyCFXGxn9vV2KorB5I1+W8rAiC1/K8TJ
mCCjYXKTODAd2a+1dZGsV65hCwxQ8LQINje5Ffi6kwrRQqw7e5NKcTtwFD5n2+vt
KYAA9Tfz1tsLzef2HOnJtkQ26J/9UZkuUTKIFrZoGpsKgXWLHA0enIWyCdlL5jnn
+iENCxiwcAFQ5adAtKMdYO0M22n6H9fIjLg+ZFd5QBsqt5Qlb/uQEGYqheLDij2F
/ug+3xrh7rDmzRKB0UFaQAPdVg0KIvOb0YhOyCKrYNtEVRaOf0eAm8mfLtZ8fHm7
HOrteOzw+ZalLu5B1GL5Ony1oP0JumrlpYvE2rmx6x8gsDHpyrrJZFhRm3ZIuKpv
+65x3UtyS+cePC/uVSvaRUOLdhJQtI6/Lq6QRE3KwOOYeMSeMOvDAQmIxsYDsTyH
BZVbpMce87RdpjedcXgUYH+OIcQls6QxWxvF3roTuxTjb/pBzPgO8Czp/ARDMu0w
Mjg3g6T45XqjdNB/G6H4jALwvCRNtZp99dEez1/rqZEOLrzhGrh9Voq6yxgyPjHy
Cvp9hfyCqkterUltrdn0Tk6uogA9z4ELZPOOS7XwnXbojwCk+1hWHS2doD6WYor1
TejQQ4YForVos4exETIuQ7n5RioxTRQrZ73JbxB2+FUOlFPvggfc3Ny1VNVq7+rA
7xbTm+SAGvTOziTaT7WgGoo3NztgvqDKVOfmGPTZo4AprLi+bRphk6gSTGUSID3t
E0WMELeiuPPDBmMse/dq+7CMRLvH+bNvd6Ba3sBPKTMFEquawOyIEyl59KX4SiSC
FPMSiwc6dNlxeyqMZR6heN09SEPo/bnzfltIXw+ePxZTO3htXTkRTnUGxbDzC9F3
ifZFhgZ2NO8CZAAfeH6sYx3h1A/43zoCVaXEDJeKHg6d5UrOsg1NZP6QssuPx4ng
5ZTwoPszkjxrAsgQyUwujuTukPbO8y1KsqJWYMdFd/ZgOCbO49RuaiwozZH/tLMn
RV/KMF4ld9oD36SGCTbzW702zxzF5l66kQXUN4IhTyGMOkwppigtT7Sbx1rx33Do
pOr7uShfDiGj3VY5MMs+rEZ9Mx1kO2NXM4hUg9Q3h7utJ8UUNpn3L4AHnSA10uHL
PKB038kqEd5fJNBcYxHXxRiJmSBBW9sFx3sy22VlNs0dl/YORr+AXIHfqtZZSc0o
ELgphCK42X3T20In0M9iZ6vIM1AHvUQWepEv2Gd2wjCY1DWs6McX92fPEQsaG6Dw
IPSwaN3Bv8ZlkoZm2biAVqaHAaYQUTH3OH8o298qBTWlfW7H67asQgowGtqsDvv1
XSxVMEk91sA0hQpXkLsIY9Y4esT2dcfnffgmB2Fi0gNGCAkSfhW0tpyY2gHeLrgR
Or1PvelCKlcO+53teirVPX4W/BL+AHPLWz+vVd4vFdZEbpW9igeahetdjxfUzaq/
guNJXkHRquqK1xXn/xgFUWPbXgJOp0S9YkzwNKHGHSgFOVVAfn1nQ3eqjPGbVlfb
NEOV3lotzdZ88LrftTxhEsxyFzX/bPGGa7k0aqEswO5DvKLji1OBbUeAYgKoRHy0
6Biilj5cK7kyR7idZdbQjItEzmzb6FRffKZoy/DRSt2e1/aRmQ+sUb9Vx517jbbM
JlWIMHDXqq+13tEd4IGXfpLUabvLt+wXhQp+ccDkgeVikV7g3janEqjwQ/wSPQg5
/hbY7XyR8ubpuK1Q9D+Zxl/jAiGRxz2sfh+tbRqWZhFTEWmWieo/AbGIV78cBWcc
pvNoMEHxghmjUmgGoqF05ePYh5oo0NodI4vGjCaiRiAyXCP44/m+1Z/nQOkN8QAL
iMZC9IlSpVi4ss+k/NNqzRZX0YQwSvk7xrYFA0UasL+cfDxaIc2/OeR1nAC++0wc
gy8WceRBGP0geKJZMnWyhhagmkXEYfSxLrCy8Ksj1xFzBUQv6b4AfVHSJdNu6c3H
HN4v8TRoXf7V5+nxr4C1go5eXAKHMc8Nala7hYyC+Pt7Roy/TVLNqoY0EPfhHY0M
UaO7A8NvibkZ+l0BTgmXtCbEeG2LYUFC8qd3T7WLTbG2CY+XbbSpFzLZYL5P5wE9
xTKwnHxW9X0A7IuprdVRq8NCzgf7CM/0fTUo5snCMlpSZYpJfyoCdLib8Vy8Jpj6
rEML6uZHTObpdkHjkLc+mdLq4KJNZDJRivy0KgzmfyhDjJTXEHfANrBQEDmNOJ4D
qPyhrvswWNQBjs3jaQXsC446SHAEZXvL0Vp5+yeAEY/yS1RsYPVtmwT0yM08UT9n
I8XRa//5ycBXvLKbxqVlp0N/TYMg+eGe4LKPfEzt1GPPXLl83qvEVa3rUCQw9E89
0q5MkCvkRRm0M32YyUvc9yKGSQNQ7D9XEEuLlvYO2/pyqojxHBfQycSkd7N4nZAD
1tAmVptinu76OAoBWf4d93b67Vi4+qhUUk2QVy//UOzgNuCawmCsDuZX/+FOE3nn
VCRCxDeK/hQUQJiQvm8mM3ILKVmVI4VlJGzisjuu1Ttrm/qUEFTbh6ugwI1ufIFJ
l9kIqJY9FFXZjh+cJXWtr7sk89WDlkyJ6u/ET5Dpak3jX0s93ubWDbaewcZnVWon
ZGwFRTp7uIhLjwgscDPG13x5KhNXHIMvF1gDlQjp9YTC8ndWExif5UtrUoAFkYia
yDTsMgJDkFxgxgveDNXPW1f9qWyJyjW854l5/xbiJ1vQ1/x/olc2JulCdk2pVYn7
J+xPhm/x1ssfaaugqH0gBdvI9BUcYP068lqwawJQ7Jb9N61T6cLQ9f7m/G+yJ6a2
qrehvH2YVHB6KaRpPD1cylaV2k81Hok/GlhzM0UO7Dco+xtFpRWsnJLRN8XXO3qC
VsXRS2nGnw5iVN7einBW7HTZpUf35UGZyqj9hLZaCvz4GWV54iGzzOGuQQjejD7C
1CSL8sCxNIma1iWUTv6AwDYj2fcO/F7jLhDjWjh5GPqBnHRUtjx45VDNKMBhpN+c
apI1Ylxf0h0OzCPq/m+WWgKXXIN9bfyrduvLFSlGkSIGcg5qrJyofM43BOjqZ2Rc
lkDmZAYfGsfiE2OGy/wu4HTpXdH1srjx8ZS4ur08hjNP0y17f+hINmzdqbXePRlx
cI4/CT8jKkA6SiJrX2jzHMo76/ihveOhfDNy6QV5vqewnT9lcCiOkyZOwMXPKkIt
dg9ciS/3pI2hiadvCwJIJFHhptnnnt8NmoenJqFp25V8mKVaxpoemoOFguSR3Wsm
FY8Yh/UUahWx7DXNG+drab0F2/AhAJmoV6a1S59Ntf1qDmqtou/Yrxx/4KNo8BYa
`protect END_PROTECTED
