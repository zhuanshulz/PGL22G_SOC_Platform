`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JBK/Y+jz5uXOgtISx08t6v/ci8g7nm4BjMB940eiagMdOkNdGEcI/6w+vxcjcyep
jFw7VRizhX8AqUriceBWOsTkbtStPYCs/hvPcZwyZwKkHDYb6EzWe989eg2S4gzZ
SxdcGPB6z3lUcf7MHXDof2t8FRZyKJf13eJzS1/ftMiNXYfHoU5P8983enbY7NVq
jSO8XsaYvpeNOlm9L7+jDOQeL4jkH/71YstMb5eAUMYtCCm2jcMvSfkUA1EmreCF
s84Vb3eOJsoFiczRvYJaG5pzSumFDr6IckWBy3Dk67EBawp06vlNm/aw8arG2Pcf
sMPt362DWkxXJBoiIC1fMLj6z9dkaHiGaQ7ZpwqNpZ8EfyuS7WbTFDe1ooy8V+g/
9zmiOdFJC3D7VpV7BuiEIg==
`protect END_PROTECTED
