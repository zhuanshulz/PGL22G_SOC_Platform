`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UgW1P87RjsGuFgl5b6Gsde0ieMSKDaOe9ml39XW3u5J2kgVvjOr0y7WRP5Hhhn2H
SKdDR/L24LTrrewmKNPa2tZDrs2NL5fhjn9/uJAUeHcyejeyXNym/M6owBNLBnFO
OJtQWxlJLfsTBHEONiJ/6+v+jtir9znoHf0X056/bmQWqyYqfAALHPqcL2Bcw7lf
vu2A856guu4ZII1ahEDsns1f64uQ6+1J2osAeWxtRIMuZzeJcIwxqYVljDTFrXQz
iQSkiSgpx2Rbv4FeikFeZFCf25nzc1qL9bB1QOXQgXO11At5OHI3EyqLtQVZTszV
Kg+AEZRU8vQnUISkIGP1LiyTTUuA4Sgw4IERCJVEfR/VedlvMP/wUif7Kt99pu1r
eSBt1VI/jl5bEt461McBNbJm+Ad5S7MGFmT+vllBIwR1x6zoRt9K5iW46p2bq9M+
EAP4Yjc9nvQvu4vqN3z636/QuZQi5YgaBdS0CDbjKq7GW+ImbEIo1ATFvEiHq4ct
buyovNmFIxe2ANi7ZBeu+FZEFSVgYfWgt1zqmC2UwliAjXlAR4/3FbSwuKvvm/hW
NTkjQNnCtUfqP9Jq6SeB7hoxO2zLZmEIDiWZ1lwbTXD8L86VE22b2gvu/XH3hDUk
3xzMOpv8OdKzec//ms+38WAEH3dNWcHY9reXsEwx+b0otuGbT3heHblJvvfIcpen
+QYUGGtHclZUkuwQHQ7ZMpYUPqwza3+mZqy34CuUQG92EWuAR2qWqReKHoQBBUTW
XRviI6TsX2ZXyKun2aWShiwHLK+1OJpJMyIZLGFf1K5SF4iRGCpo9gNFz/C1acOc
CBoD/pMHFNcXCeAOnnwJ/jTKSIS2EPRsEtqfLpRKoG5BujHKQh3ul2x7tt3WgJGb
YDnM2DBYpmS/Zhpejy0YvsNsfA/+qtZdyUlAvzEszMV0FfX9MLLjyFIHRu4nv7u9
e9Zi6aaojaPa/DO1qcWEheEzUz4++uP8/o8HfcVeEmXQ8+5kDWbLNW6SC22uOpmO
oPjLS3rapHZgB3jYF8xiH1vBqsS6EcL0Ud5/7O70PueHdk+7VsK+PNouVPOzrS/e
jx34suwcl+JxksuaiGijg9DT1yvXofsBUdQ0ZRNHUmJ5Gp63pStludweBEguD8mG
xYk+GLMzM7TOkO4I+nO7Bd00DUQ1b+ptN+13ryfcEsk=
`protect END_PROTECTED
