`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PxuUcsEoVS4UKTbnSNmejcAlkpghCSVczflNW2Ir01SRpW/zPa/PCEB/k7eWtNoI
8bT5dhHRt1iz2WoRjsrtRkKvmq2UisS5+9H9IHXjZe7IRF2WWI1giCzO/1lqt4vk
JTrvKiW5P0HGsEYR/opmCfrXu42Ca04KsNg03cXgD9Y5qhKpwI6GPCoUvvH1HDrg
uDOtrUikWgDlW9zleNUy929iM/6YEAfSM544GJZGpgLmwNtHy2UvAcemPDbv/NGb
cFYnuETgGZjcpkpvmKk5hq5zspQnao8Pnhagre+gUDzBkuVPf3Pcf+TxmdGgNy3y
fkO0tk0+ZFlr1yiZPjM7DkNa4xdagulMt0X+3iwfasIKeYbo0ukzEreiP/elOfnD
NcBpjwm8ljS681kZFFo5gbjEr78iIZwibnNdajydr10xdwM3iJvLvSPFUm/AwJZw
4qyD99VBVjt2c+frJ+pUGkhW/cdkBtjdVCxl7y1/Lx0yOVt9xKuoIUC+1XhmfneV
p2tyiO/Uj8KlPtj/T7pCFhZKA7focY5Qv9ycyKb23Iqrmj8joUncxVIrqUMwwPXV
eFMLNNNinzzVtqCBait4A8W6R47jPCTkbTa3TxhXeaofLRQFdFhOLlEkMAw+VKq9
QV/XXyw/8XEgPv6DmSsJjT1XtR2pCrddTavBtMTX4LGBV44+06bDP/nv1eGkhuJY
/4kyIiOun+8xXvDNOr+ZAsKRo4Mo42ZS4tWe+tJbUP1audP+EAPge7NZOhx7bO38
5qlyo6ctxqUsDWRs4W+BrMF1E7g4kZoAT27CPlRbk14M2mYEgI4Eo2Vj2wVbAp+h
HW1oi5hZOLqzfp3u28hIHIQvjXodeEa8jcXFeTYPzVNNqfmBqAxQ7fntsa7ZVVwy
Idp/E5qgI6HKHSuD3OvrUlHP3ME9muOSPDn6UMN/wV1Qzrf0iZhEKbnPq/u3d8gF
UXY8imbh2ezyd6qXTOE0NItQzOu1Ak/9Wfhcg86ayjls4eI9X1I/OPSjRiw6UwTK
1u2upMRRxSDYk+glXUkEWNNmDoEehvJRp9hwx99YghKP52N6n5r7QUdsHMEAukZn
ny8RrpyDuO92FqoNPBxfnBPUUgsKp3vpSbhRSyYvM/oYMmulW+93oycz3X/eDuZy
Se428qxGOwly/g3DztA13RKj+iWRYIz0O0RMQ0rYABsLT6gtRTKZtudwwtEjoz26
n8pxFjHs70FkV7086ojjzfyKhpBAJEbrIiKLZrvENbKhtrI38h7Y6roMon4FhEqF
h4r3PbBOgbhmr6U0llR9eBBf5zFeQ9FUtvCA7PyhFF+wpcKXu8IK8VE3evuzHrLP
kTN6Stv1e816bg0kJV+g8usGh4qvwGejK2yRBNrfQg88E0v1EUe9Qbwzc9UROLX4
fY8h43l7pfQUy6XTA4Rwbn0w7CqmozZykMcGFWN10RGUTsKleYRKnu2HRcnUJUt+
9dlqZbO8ZQQv1xAnjTOdiBAmFjHXba+Cn2CC21fou6lWoDMqUSIejp8JzS4hU82w
LFMwXH1A79q4iJ6fa/JQKAngGB5ciBp4Ebifzwtt7PEAfSXUdEW0V+3WBpPYrlpp
W4i/yhuvlWCoD+Zyp2lSU7CtzeHZ/7mDNLLAa55RaRYAyc+DEzaRV81KvG/pt90g
WPtiS+m3VDX2c1gX7dm3ia2Lxb8VQRjYSwn73gqxT3HACvrgE+NOKc2ymH/Vm8m4
Pm+wR6NwkhLUxD6rkEZTjQ0ezDuYGSwI/XMklbZms/Uwq0yIQilXIJ6IV2ECzdgi
PiJrIXEKN9wvladbTPLwgT1sjf/3TbQgU7AIEGyXONFRpF36jJBLQr+UiKcx/Dmw
nd3UPsg68qNpniC9amhzZKTCRRs9Q6Y/NXO9b0qIAJqSlosfnttlkP6psywPp7zL
J3oAKhJdVZF7wtoWsTyAPiYetELWldl5K+ObU8kqqMLLFLeNb3W9U3E9nVGq/Zc5
mvD2oQsYZCS7yds1D3bITjL2WINdaUtNIb1QNAbMtQi67eqCuv3R3s9upAdpys2Z
s36VPqFYad65Eku5jSE6gITPAn1NokSfJc//hoBN6OpVnF4sHsXyswnG+qv6Qe2h
J+1HDaYC4C9j6iYdPSewpyaDSbS58sV2A0RCVaMZLgI/UqCfyQZbfzD4eNGED4JE
du6MXPWIEWZD/YBr4KYFBqafRYonw4gYAKdzABQP/kAqkzgf9+5sRQdh84OgbSvT
XPUNUZ3w296AOECBCtSlgmKjGqo/aUA+iCAvCAsNR5+eSKQ2wTiWzRjaKMOU48Rw
yEnabyuNtx2I/MVQGdIulAeWfmhd4RYM2wrjlN19J1C4hcOpHkqCZmJlVWYOJkge
lySYD5YsYeM5emXxWIA087Da90oEaUixXFLZkUt7SrW7enEwyu2rnI25/cfJwRGE
jZTntEWRzf5t3RncB540ANusHUwV1W4yQXr3TvR9Jh1iqUwI9CqdspO03HyssA1Y
PFZS+AzLfxvLMxNoSOZq0Y3wA3C82cCdGgfcfcOd9NQiX7/hFor1BMgHhN7Y3Q/o
KXS7OTB5ZJLoSNOYFibWbp3M5QZMaT3bhmTiS4Db3euYWH320eHENzOp8zlf2VyN
qJGULtykYe4FVUtEl5n4TM2k9PCog9xev8+KCAzrYFu86wiw2MO0UKmqVRY9HDKX
/C3PTORZsAcFrFrL5iq5B9YNVUTIblB1DCCy9hLyUFMIUWaHwVLvRwvgEwP6+hP9
sSInRGVZMdKIf5Z2SjTAa0kHZo5cI2r9azScM8Xeoe2A0DYEeFBFF1nJXOIUf81T
6Z0AJ2QoJPhbge2o9W7kilmId7e02+6XVFrsicOnSXF6ngOWYEGbkpedIJztWSNj
W5PDpstHI41Y2AKBjwFo4WIqArFoCu/vkuIKUmgp/DJ6OPXKixnfUR9Ur1heEWT7
GsCnajJdeVuEQxuDB4j8zVvqf7yHEtpbu0n4yWtLxiI1BPqFBBrJu4gCxPrVVRmN
gO9+DuLtKN5S3fVIRuOkrwUshahGYQELolVd9quDThF/bq+aeANzvr04PrvZk6NQ
lzmE2O+uMxJOMAKnn32vKkBnJ2Kb/4DjS7Z8fLulfqvioSqc8rGcTmU6kaEuCbXs
g34ClsdvZ8Dt7k/e1/rq4w59QRAGkpAU2XEV4PQC/QVD3vvKV42WJYzJGBT9qQzZ
r7wi7Vt0rZ0jj8bOFmTEz1dJTNAyTsEl0BxBb3tKoQ1yLyvBS7oo6UMgelMKYbof
vFn3CqalaQgbw+TAst6SzoW0p7fd3MMmY96XX2fqeqVZzIbmXStFS5JFoXRsZI6L
VinFu4kDkil2FHrB/T+9QNHbsJSrIqLGnPM2BE6f/2v43lbasHqD2GUOmXr0OlNy
0oKtuTya3I45I/K0xv66qiuHOx5+COlDe5Sc7HkY595S2+LfN1DZVnDb+t4TE4Cg
cGucXW/18w4WKm/Zue+Oe8tTjja+0HcOGf0Osv2giR+gdJOxiHWYv0TxP+dp7/uq
aEyZbOuT9tqgKmPd5tshCutRJqMoW2wf5YZELFkVkshgluAKU2uNgJGxB5htWyxy
6fIAO/Wp+KpA+0eznwlPIzela+IDARlQiEf+KLtABMXL2m4dqyg6z2W1hM3oM246
S9xgn7zK3+A8/4lp3TlOpgCuzn11tbzpDsa7pblfOYIPBodJPOja+N7l93muXQX4
9YbD700/M6VBHAG6BxwBSxEoLHg92OABgHq+VM1NIWxZyIWCBxunsQOUIR0G401y
r8YQXfk7DD5qK6bRM9ZnqmfJIR/nCMm+5oqNKAomtBzIZRAoBVDbyqcoPu7bfdkA
R5xVeUrQkYS8uYJ30PiPVe5lZ3jfpbI96h4J7WZzgaN2tt2ScCEkHa0uXGh/qdLU
CPv2BiLtobLSuEHd66EaA1ngqyvtmVFwKGMxsiOXmmjIwCo1ZI4f/n4nXo8BkbhR
ZUadJDEGiyiAwhHt10FZuuOoi/DhmDl4xnE11dJ3WDKwGcumQD1QtOlFFykjL/h7
udtfs6/Mk9LklMQkgXrc0OXwZ2Ib95vF2sNZGVxKukLia4cGHauIvKN92d9JBPi3
vQbGy8CuTE3kjLx3YO9mxWfSISufl/6ZOgqv5yjujM0/+nu9MhlanaisDuQHJ+Wl
zT92GpdrJe4cMy47cfj3+LPo2rM7++W19+mSFifRzFxKrsg4h5GxLorzTvNbw3yo
8V29YfEEyQnXnTlBAuuvVg7ZS6Kx4nAdI2qfwERyZrjnhboirhxmQ2Z/NHNlx6hj
HJxkYrR+t6wNM+e7Phe0Dt9FGRG8UcPXqXyFt3mOeFbO9z7CzzU13IyfY6CWZU8l
KLcmn9CUIRlF+1KSRbbUDjJCXYUtX6f5m3BEVR//bZGhURPrwlj9v/t0iYkii/WY
LWPuOpHvU8mF/YnwIgMeOcC4D72X9qTRuVCY3AycRdJc23CX34ouADTegAG+xJGg
fkQ1tAcQEeWWRVNXkBf7dSmk1kEvxFjMXKXazkSP8Smbp7hx/i+PYdQOmksbYeYm
UswFiRGDlu99KGg8alT2TctPNWWAoIEclDXj8WLFlRbhHfvQBuFuyAFHp8eKbmC9
079+zh6zLKEwnWkOvPKwbxY/6QkIQzrnNiTCCMNgCzbHTVjMm2YQt8bUXUZ6Do1S
wWQhz3SkJDYR1wGS0twPuN+R/E5JCztTaqTfs5/WF5Y+0pq+/rmF1qG93mX0Rb3Y
2XAIs8qf28TfoegPpijOrMYwyksydgX08YW8orzIhq3jU8+z7IKpPF9JnqxI3cbn
5jq+spXHuS9rraAs2N7FLf/zlkc0swPp91NLwwcf+aP/Z8/QqvaemFna7QaiLaim
FuYb6zdtGFn6kl3ZRCZ4Akewl58Yxx62A/ehI027ZgM68y4FA+QLqgrMeX0TWRHr
4C5Bh99VcLuJqfny4/vlwmz943CEomSRhfPm4kkSg2c0nbCIQV7+9uONa2E4re9F
sJOtvADGXWXeQWcjoO5ajJRXHNrhfxSFC7PqO8dURya8R16EzE2QQ2AZ/pfJSbLn
TQ6KfgQ8pq1Kq8jLcOHES8kRoiM5gKMUwPELRHksPGkEx2vqIY+R00H1egBA27Du
lLsGek36GH55j0tLbT6FlIc0/CIxU35SO1N9ffdSrCRPU0RtDB+TwKX4h3O3I+Ci
0C6gMxQNSX1Vlvyiexq09R3519Xf9gwajXa0k1b+9dc3qwmVdrj5ffjHSJMOlRAT
j0ZxcJxDkx1CD8htwWHiSM0L4YBBsj9xJVUOHzWa7TMv4uZk6iGu+d/lF59ei5CR
rdrdgOtqkm99jRTxz1TNPhSJqYuu1XdvbD5/xtYzXhedLB51JkmxbleEwKE2tWwi
GCdspF8+lT5FFglGSoLvNj+4/sjB7xKrD/qQPDvTdTikWmZZINbUVgFH1Ntxlcir
qrwSlnVWSEyNXjiZcLcVg7jUKL7hHUMHtHHZ85pD5dyvwOgjs+4PB4oRuEc5rzbA
KvDc89tnV/mJMyBD0l4uIkEjemDdM9PmnSL2R5t/+XJzCsyzteTIPTIkf0EKrXjy
WnblMCFja7LZbx6tXhEOgWpqrOlGhFbShfMCcmsfw/cr/Ki77KLVXhJHXs1VbRZt
BzmXS532+JLNdljLUeRfNczXM2p5q6DlI0k7MAgy51fXtpCkgfxOAjHvTWJBGuv8
lSIePMmzSSLaqEwPTXWtoehmBOZjO8WtT0wj29wqXjmBR4XIvl3bduKjXDHtdu+6
qLeeqY/TdXpUtQRBL3HcO5kd2+cb8+9Hw9xU46ZFNzlS86qGs87gO0WIIr0Y4c8d
Qf4Fx8k9NIZf9uDDs/BeVf3LxRvRbCuSqEJqg2u4Ud89+EfzqZ8Ninbl2v3qHYMa
2j9JvKWTZz1P+MlsbazEJ2GBG3/xzXjpVezfeBSxSkM0uwj6PqJLaBzma27VjbP9
C+ZxNC9WvwseJx4MiVWfmQ8y/S3kwjIh/Z1uz7LtudvbD0KHbik8ER/kDYQFIrig
0tPos9RWvkDM8RlJ+7RJ/9seerNxRKzYBHVPANBxLXIewXTZeKdTedgQTKgq0fRQ
CmFzGAfyj8FBjgJR/p+65qQ4FqozrdaeIryu3o7PCgvYS4/4LcxBocLqG8NH/Okf
ijzJWILmHYAgT6xa6GOE8EcOiTBPQjxjrrj387W+kbR6rDQIXP7k1D5yMGz9K4vY
GIUw8STZ9tmOrxXo5e3ajtitsDUIaidBtUwtibwYJHiQNh9ydHeA6lJ7ZHSG04ld
PfB5mmd/xdYM4ZajYiMr2HDEWR9NoPZMVkpe/5+FiTmq3Umcj/C3DWjHAVvbwIvU
AL4rCDFFIWULHfkaBO0S+u5kV8Xvs/aAUioh3KObgpK+RMHhhTNeJlIuJBOCqXad
IKnHF2cuj0bv0MootvaRQRkFTf9Iw3MrL6vk7Iru0m6m9LHmyLYNQhWOCtk+6xAJ
LMsgrx65WJ3HU7D6pBSBgPZO+jotAp9K3OXr+Sh+3oBbrDL/pABHOF/HEysJznhN
YeA5e4eyJEFQXkyFrEpkT7qf85JO4B50a25NzRmUzXIdAv+o8xwp00MW2QX8sRar
z4fEUyd2oUk0/exMoyiZv752jjVfaNyBcq5ecysx1um7evlbQVphLMALOgo95QE5
UkWWAW3LdzAjMLja5RSTkzirCguooqqYvEgYfen9wbiJqag91Uv8F+kA3tCBOoiI
aN7DMlDg5d3I8tsqEyM7ITjRoUAzyxT+N04xaAekw7o2oHqr8LYmJmbEySi0Ybw+
HVuEBv08IOy0hqdSW+RWVWOO0O4ZCxS0yXpSbJyITmXqisUh8PdtTu0LR2s8Swkc
a5Huchi/333zfTb/dMwFxXnMnLdysjn+t0mXUUuenZ0kYRXdwjRmXHZqNILjvq9B
Nw14bhhLU/TuRByGk6vUjKGkbIwobLWGEja9gmkuxmEzruiCR33In8dsju8bI7TR
XuphN+n2UIWzOTih5CWvcYXvPVvHph4pj9QLNdhKIkMzdioSNSw7QF1w3HzHLdu1
7lzWE3wWjlYG/uZdenGYAl3BeSoTRuoe+IfJQm3i64+/vW6MTj+2kmj117mj7pCc
/W387347TUr6n5T2JHTzfPAYIPJoj83u2XPzQtBx3DCE0HZeCy1Xxk0gfdNFHbR+
jcMGPcoEIqQu/9a/J2NwO7J9OYTbzWRc3VOQY32s1i3y1q2HIkYGCNuKxugr9S5W
ctY+1/A1n76iAC7sn9eDbfXOo3qNXV2bm4vjGwnBSIvhomkEjjeFgdlhG/OKpLvN
Or63V4AIhtWa8GqBU0wIYFkx4uFq2AZew97lLhrNAcAJfV5FP28nBLeHRW9oAnxw
Oj6XvZI8E1WVPoBulUpIEQTDJzIgeXWBdttAX0vAT3KIkLht41LQC5HS18J/+iIK
OxFIiVNMZ3okmGP506F+iuVzyR2hMs3AzifCy3oKQzzGOKaKCbjld/iqkvbyif7X
gwFDqhXHzykLZZ9ermIA4iodh93XiuRmvAVVPbppVjN+3bVo+FjVS45vDPOi1jYN
0/2Ps8qGqsbbo9/UP4iteH7UZw3XM4/9os96rGjP+jnsrZH24n4FEE0uGFvjHfG9
NyxSCbp6PLAGwK57oCG8HsmIFNBfLgDTakaYo3uQyLXpvU5tuNqUerY1ym3Mm4RY
hFMa0d38C4T6XYGsqbOIu/ghWeYk7p6OinPRmuN0sT4oolCECG3v7r5IwCJuFCAX
A9w2JdLU2iSQIv15JCRnzNDia24SE4JegTMtDYA9p11WrHkSYZUUMoZ2H2Q8RnrB
f73PKhdqgkdjCCHvKTQYDfvk4T4Rd5W9gIA/BI/w1CgHo0avp42dV44EYcQ4BT/p
ESvFkyXpNuq9SHIeLfe3KMGQCmesk+oSXJY60GCZhpNRXV6U9B0oB24Bj1Wgk+UL
TxBd8Ts/khdTh0HNoUs8NbQ8BQ+DTCkjy/vKSkNwjP/WkJGIx0PNR9Bu+L+v8fnm
VAJ80ecb9hqIRr8+Lz8cLVxED5xWNqASsMd68Odorg/WsJOX0Zx1Kqc7sRQnhAKa
OqGq84jeYqMKLCqfUsegA4YzRU5l+oswZSinRq3fxChAWSep900+hjG+wbyw4pC5
avsDQUEcTz7gSIsoOnZ1t87TD1ienud9RyopOWeVm/NvbFHAP6BkFveeAqHmq1BW
Tlkz8QhsseRGFqH3VDjBLsxpLlhuhO23Bkn1THK/+ISpYdZo+6QY1tGjm7A2OMVI
oSzaKFv2YM78iSURloDEr5a4Feor9YcVhh9hloVApbBoLNLq6dMDc87KS/nSeIHe
k//IgMmo+wmTC8E/KEUHsiSlUcoXGnDhFDOJAYcq8xhBeQtLPkfKYFm9cz83qe+d
OEPxDbao1mQDDgwTv2V62rMaRFpgXyXtM2pVHKlNWRFMiErhpD98SYxuUbOVN9XE
st+f+OWrh5KfkyobUfzW83K3F8P23X3hS4cJIR6EUytjE9GrJw+ovPaEVgFOawoY
N1FT89tRWm9BJI+abLbbRUGifXxfRcZkpla1PqnSVwBkZ+axmUPDYkScwYeyU3Um
rfQkk2/Ry7IjGhI0EDHw8z20sbX+K1gnkSxl/FTpkQUWB+fs2Tu1GYAusMfeMkbS
fTOQU+3xFpgO+Xxru6TR+HsLcIRJ3gyMTyGa3dz5uJ/+H2SZ4Wect22VFkatgBKM
Q+AfHCfxJncAj6ae2KIKEUhMRVslLlF2w0fZHmN/o6FG5rmgKFbt2nZo60f3RfJe
MEZyHTGmZYyIbAp6B9cYrTQn3BBeG4MTx7b8kU0u25XNXsnUyocmdxTAIGESR08N
0+CY7CqTR9rDtO8jxRW7O2S9HXXYvHMnEl9BQ4QFIJlLy+I+bp+9B6CI2Iqo4Fp8
z0kae3bxRQabJVOotJd1eiUm09WFessGFCekXhYmf0pjxxTlrNXCNgJwPSGDpLIO
NWLet7ZTOHZMzlH6yToKzkD2MtLQCdMG1TUpwr7u1l1Gj6US0pcFf6FUexSmwb7t
1PZhyF2DbznFl816JRnAKB+mTF8r//+kyd6UchS54lZo/F6y3tL74OG1Gl8j95G8
w5BM8Uept61iDUmp92LbEPb3EjbE3dnA4j5BH716pHbGsD/yhIPCxuK+BGfQGdKu
9BFzW2sOcw795yVHKHmPrhXKl2AwEckYt6xvaSsd8uHZMOEaxmJivOx6yTDSlvJq
7u3+JAui7uOXj60HV2/I4/dZyUzRA1klhQLiD+tqV0cytIC26NKo/kCbqKV6buiU
dXT3zIkzVbR3z4sNF9uKmc40D0oliO8jjCg1CEgn5XvHEart6PRkkYX9jYUGzzJe
veibMVUOVS7JhGCEWCk4etzXPNwed1EeEUGGEyOL74q2FF8Bl0/a1PQkL0ulkchO
PuPxjBiuP4ocrUZGr6J6w3lGX6NJheqCIgYh7wfq4Ph5vPCG+ejJS3o4eOl+Kq7F
Np8ZsMXg6zcVUbFnI0LMxMua5wYBa/X3dUsbcxJ1m2gHnzc1A1b+cOWE72oCWXg2
lDKB9KB7NsOyhVV7nTl1Lwgg74k6SGxVRmVVxQYl34XcKcSJUaWihTZcGgj/tf08
VcV9UB9wbkZwyJ1MfjOAHEgbIqwKdip0bRGSwAjOguBOlrLXJoRiBbw8Mo7O7m2h
5/Z4rYdAsfHD/rhn/L3FS/1SzTVQPNw3tJ4oOl6UdPDGuVlJSeo6AVxDIaJnO3dm
fcfeHXq6K5Srh9zthZJit6kKtlhXGnPdJshrdZ8zR/qT8F3WjfInCR9+/zJIEBZ6
1hY364we5cAg4Iyd1+BXBMHn9dzv1/Ox3ENyhExtIcb2IOuI5gQ5kkQfksZFO/go
vhFExj2LVWAWKk8GE4rEtroOOBaDNU9PeA+2nSSc5fep7o3qd012cyugnTQsVAlg
K0imgGFTAX7VKfkC77JGvuAqD9jrJX28kfSmcPYt7kHW058TG+iLjc2PfjgfHeQr
jaMAT8O0KAPiLkeHiNjpSSopWkkw08XQhOi30ISS6P0//ZVzPbBC6/qvE08p+m09
4DV4Mcj5k4Zut6bsQTHRY3fbO+yAOCt+ZknaipOu+ocXtUlZtjLtIkFoezxXZ8a7
ATg4ofN2vWDsn41VrAhcykVSWIy8RoYskbKsH0cbciy+AyQ5BbDy5ivt/HVLtjr8
yr/Hsx2U9P7+q+/umb6IZ6gx9yq6zDLAOsnJ4GsOymJ+gwbdED2E6jhkBlgj95As
VBsBX4kphZ/FjFGSqWAftJQLC08cq+sOTy55v+5pMgoKILuCjib1p4aN7TIzuFMS
DrlzdNbC8ttbCBV0SzLI54j99HZFREQPazMrSehyhphEjsM7K2VFPwQme8MnqUg7
txKsmDtbVw5tKpibVVssLHRv59/osu9bVOGraxJ2fUm4sQSZpoSCaeKjxJj/hLY3
Rlxf4ifUCZWBhOvY4DRM/ZrgxZbYpx9VGdcERtcjlGiQ4QYl1xPjHNC9EyzJobIe
beoWqnTkIGUrcpp7PDc4KojY48fEzsxA6nsvK4Zw65O7bnvAsY99iBV7ENKYxEGn
TgCp+K71bGKYjeD6pxJNvvzE3SnsYxruhijVY6ceGabrfchck+ovTZ8cIFm/T47O
M4n+Io3k5xz8rlo1osFVmXSKYCNWCLP0xo20Wg40iUmn02Ui7OuyjKCc9BXt0Pgc
`protect END_PROTECTED
