`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kHqvlIrYcC+RmexAOJDlR+VjQ1jT6ED+6n6e1rbVczh9DtYUA6L1vx0OP7IY8iyK
OHiKXyx3MeeFhYuMll4Z1TPrkiRz553XZd1Lhb8b79u8ZV3vQwtMf+bPgsXkHt1E
oGUtnxcfcX+MSxVsC1rozlorrUiYB+ULlYZKo7jAyAUMoZAtd/Ei0CnXGhHnzpTG
yKSSABt8be9ecTklr/8kiWm5/Ndqc6gG3oehhasPBm5faI2XYAxmcSXT/wmZcq3Q
TAEwacP2pdNarCq3fXE8K9f7ywVjuiHNlZsl80wfdaZ7+Aq81ApHYw1a1c49mCYA
CN/64QbAAXwtFpf2XxbE4YH4y7fwUBNWv245HqDVdOECFJEnz6kS+Gibt+RBZdVi
Nmaju9AFwuY8do+cRZPmjHyD1x4/vLFUsjBcMN8DAgaKjzxXAy3SGfmqmofPpLoc
j1/qrb932+kFiCb8wnkZqAY2fp/CNlqUQJz9xop0kS523KCjImMJuf9CYWzB21tK
SnQveVXV/IXC9YbH0qi4Z9aF5mIylWyf+YGItJCfzqtsX3rV4RLXP/P3DCq/7Xg9
upUcx+AzQSx5ZJigYT5UYwR+pFPHw6I/zx48ZHKAfzAyx/LPjt1+VdzN8AaXnc0P
TmHBRlzHW5mdQ/gxbqORYWm8YPQslyZisZnDAUd5RUR2dk7krLUKSUOcqiKzYyqF
JlF3IAfQi35FCaI/d+j3Qbi5YUba/Ic21tkQG41LqaqHNKD/7iZM8q94itzbDqZq
bDUp8k6C7WRNakUWbLPdwV+0kR6Zp9O2EpZmpkL5OY6EUSXGCeHATFVTkUO99QGT
cdL04IwIKQzxtXS4t9ZTPL/ZU+blvzpiMrlc4jrunU4pWjAfYAA23+lWEgulj7iN
L3eHHfdap4nAFZeH+Tt7lzhEYRleNLT+HbajezMJLwO4LMjOvc3nFr31n4lxbEiz
tFy35lHxvXcAyvi1muw9DOv0RjJlD4KTwyfG+yjn+Xksq7sb325qO+ktBEvNRufn
oJldAWQqffasMiN3JqhMDCtvQdx+bfcSigmn7pI4JnP5+pR/DUctFxG5NoIybQEk
cdYF4iNat7aJIACztoTsLAYwCnw/4+UMG2J9lchZb07GgXNdhx1J+yHEG8HDBQYI
8YZnJyMFwTeHZbphXbmptiJxpiw+NcKT9pDj3CHxcRTypH0KQjRzNUJqwplIKXoP
exkzj6bwsJsbSAERhUFcpw+/TSniy7U6aTQkRx9Qu2Peol7xmeEIChOvshfJhO7e
U7kFsRKY1wN6DC0gAKQmSTt87JJfZ3LyHUP2UGbAx8x0tJ0mkdS+lv6q+VVmzajS
cDeyJFV6mU3dwKcDcozLzI2/7cn7pwkg17jDH6A5qkvQrJ47lxTZS/I7I3TIU3OW
YviRLMnByEKB472uWVPgnb+GH+ZGk8BPJ6WKBwihGuqLcogysG1pE+FcJ1qqPNcr
xJxvHm0Lep3LyKRW5drRms74rOmfPULtrlCnuUhdJd8=
`protect END_PROTECTED
