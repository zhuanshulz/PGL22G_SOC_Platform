`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PXtH3KwiPYjaif+2V9Yv0KGetBNBzSR4+xvAFPA4agR53X0H8Xu8BecjQzMCCx0c
Dn6NgBgCriEJwpumQqNfhP0hWqVqr5i7dVAjG22b99ynlL7Q0n7QEztJtXBzCd7C
Ea2BElIiDocpkJ7/PwSW5vdlCJbjwQW2VmElcmFqrOWaww8EBlVFJcIB76z3XjRi
jHndQmaBpXrlXe5NK56zGGFtnalyPOl8xUU2Rfj85G1vQD+wkKe7Ok5HlyL3N+km
1wZ0CMJaKRhOJIZ+pqgoM4FH1oFMh8P85iNWeXXAgNBB8dQO0xS49egoyiv/sIbh
1acP42R5Xkl7o8KoDRpLACiAtpsboRt23CNr+yCWd3Hf0l6NgSD6c9MoJ4Ho+sbc
ldXaVmEdVOeM3uB+sdRN0lLvUelDbvwcQXRniiBFpGqIQFkeK9mch+Dd6Qwco+Ab
2MfxGVvXKrsd+LbOmk8IDmsyjc5fHYJQtGFAZgeQzXYqA/5PHYXYuk7DXaY6jwZa
GVOKCb9DqGCRVOjoWKnWj7tYa5jllQNHOByOfg3tYY+aSFdaBA1N7vLuj0zdkb+X
grAQwhkYQNA6PjSSFalpXayTrkgdfoNPGPGwCO0Ey2pNYcDMBJM9rlHe/09Z4P6Z
VCpooLX/ZJbTab+cQVIpK2SBXA8YOKDoDYZYMU5VyQLrZgEt9EZMJTBT1FbjHljd
zA6+U7oI0ZF46QN/1+6Ckq5g0YYUo6QgrOY4LiGB/ilwTH2uV7E4i6y21jokHUtj
fbhlGMp50NQ/WgSFQdEdLoHQxbL6V9OMKag5oC4ZVSL0g8bHBhafY6Kp65gK0Kii
WTbHFLh7IgXxrrWO1kF5eTZso2wGpn1mzcSaRDd8nru34D28nYF5w+EPjF8zudkj
9qvv+h6gpNkP7cnTiXAs3G+XicV17QdhytMcMCZ3O2HQtCvPk7sJ5TKqDOzNoASi
kfF7TlKt4hzT7/d8UKjBt06ssA/HMHdoVxsB01o3RF1fV3sUvQH02KDqzG+yPB5U
d89h02Mffrk+zvUDhybdbqyQpTD0fD20fzLO7NiewcBWkGjUJ4uV0sHnitVRQfHQ
ENEhjzcRdMXuggnACTR3YCsPvXdWrzFHICYhfRa75AldgdqPLuFDrDmZ17hpYbfJ
J6XTfG1UScjoD8JE7W4o+o/fpAK4F5f5CiCj+x/d3wFLP+1GFVNPbJNVK9c9IeT1
JGbOhQFnPyOlcOg5XECAwv4ESQJR+AEdwAQSWUoEWl8MHILBW3jvmz9VwJqfYxyC
udooJGpdmjzmuC6Q4zk7k0vj/zkGKQ5AjEdFWfu+guc+eauc//Tmhf/PzOJMsKWa
Yf8UV5X3mWB1rEWnvDX5fbpfP3NKRCfrmU6Rs4OBq6G5H7Q8NLPWgPCUkLa0dazj
3As7QcGKU8shGd2DZDvFOukRhsE4ORTN05FNYzGrS4jnAhl+vREjcNQ/PbR1ZNUV
gyxdQ/Sid0ELYWRmYm8spYybEM6xoPWqMRd0u8MjRyvnLfVQrW+pdiwSPNuSN1qX
8/e07DgBkIh3zytF3ZwLGhadN+JBifISeREd/vBh0zlln2yvMyJB7DuYl9hjhqLJ
1xfrj50VlpAivGOYXwpWC+z+YdKX4Xsav1ZTYGyl5B/GC/Q3JVonmEd1MCreFYmA
krsxUqwiZp9OLRqHozQZweESuiS45zaHbMewPNbHtZsZOJoZXo/5DkL+gzPR8HH7
tcfBJMBiHllKMBwHWmykmwBXSDyzg9djBuXhSJrnWBwdk+laDKQauGXYZvucexwc
zhHgeBPPKMMNhEzwdJl5hCqhfrSs8V6N/MfGuLG5i1zhs3+4wsfkP5LqrEpheu4h
AcvzuSxiLEcykShuYx3na7MTDw4NReECS2W0AdCt3uUjitCs6nIQW4tILUMlc/vP
aZtgo/6ZI67MNnN+tl6QxK7Wm9eH8hw37dda+c85ra3UV9s1O8qIjYZZiX6Izena
gv1+2NWEuGoH+6W65CwvkWpBXZjXKAKucTpQOkhiXlqiDQKH3V9o10LLKi3vU4/n
hORxbOvAm05vSBNbAwgkhL4bpImQfAl9Yu9+pPXEe5hH5/ZZkqslodpG3fx+U0kw
6xkLHjvf5BYTjjjhRX1uZyABG5w841UUiDaYxrVAcdLBWSLopveAqlCphli/q+p/
4qC9Me1DpKk1hmgy0tHiik9SNeF2Xb5zio3U3mQ8g2Xk0y6GE3pWjY4bnhI3dgZV
xZzkc3clQwmwea4O6lzoHLrI3eDIVegxqSYstVKYz5kQwnsXqcP1N1IrB3N6pDuI
AC48ocIjTupXnyO/5jscYYJIIC1VPvsnefod5ya/ZwTYzsQCyHCstAzX3Bl2Dfos
UzKVp3D7fNcRrwJjDHuOeMphAp70bpdnsqxSp0/nA4VMRoKAAWyIiAxGP3AznBFi
XqJlN5iIFf64SrzXqitGM4nWAqNIRxqbfomzDi/6tuYmtx7IDp69VKIFQ+ycjw+U
iRqm8Q7r6Saq2GDS2SAsG4z2HDG/fwShrUHZX3pFbxryezALqIosy9mdV2vE5psa
G/QtS2oPk+Gswhd4F8e7YWrhyschaJaUQhhRtp4Arg77eq5+/ewQXMwjm+L+iSd6
KDaTfJEWeQ60roJZfcKvmizZby0zuyE16BAmR8zg0hgDyGe9aVS1ddwG4apW5Exj
/X943dlo87MtACyIVmtOpg1yjHILBg1YRW9P9v71X+bbDZ8b4wWBi+NUXv2Ua6q0
TEthavv3nQaz7QSE53d+tvgxpoVpC1wojxE90UNALAXSNGdLe4w3dFbCi//oBUOv
bX38ianrJKTkBemZ6xDg3YPpRg5GF/0wM/arFNtL5gOQ7v20QFxm9tlMUr1Qjrsy
0XNxcaqkWNFjagny8jNBST5D1MY/wosnR0KCYF4h3TzN3BdroTnpWcomg/ruX4cS
1F9y8sfaVqUYiWkBrtVgAlIHjNgs5k0kai9xJb26+pcChvDE0C06wHeL4rL93yQc
OHIHzly4NQ3mWMKe8LH6VvPDNFjdK1Tf2MUDm1X0TxS/LZBFwtbh2h/62MjO6nqq
0ztZrX5oNdXjhxEZMWue7kqyAd9VSM4cgf81wniSRFLRXP2JtBWDYDb/CZwCr4PB
ZSWrpk1d73g5oB3aewZaSDG0FDhp279I5TkcbXFITMqTBWLVUtzcjQP0xy+bS1wz
oTnQXk64Mwjr7I1nWrnTwUTlfJSKPbzK3sGD2rIX9Vw3GkNsDrAFq3jPgjSQrepI
k0ekAFSaz23uGY8Kyk6Dl4z1IHeP/Vt6aL+hfuIm30cdH90FScHbqqEpbTKC1pKj
hVhB4vFsDVyx2zPHCiJOIQVZ8i5hHb7EK/MHWqbKsQqXyF3G5Egovj7b3noqvA82
MB6u8Wkfh9ZSRRHKx1LZjbibcWamUaeXDBstL6czL0FgXv6Yo734AEx4Yh1pB7Kg
wHOj6B081pO3jzADkoTnF8uvlT3fXECMeuphkgldc0ZBeHfqsnjvIgTPl6hJqITb
ZItih4CdXUJm+KylM+8V2fmhcbbuZMd2HDTCA+nvm+toB/W09+OgjF2Z2K0B+kx5
l2eXUPqMk7weJHDrR3nKnXXm/g259BffOOVOfdoPrA7s4PolmoMF+oKfRnBP6kVs
k4C2P/0RGYbmHm+UBe814OFTBjttVOZK824qNF3NknnWIlcVCbXDD3uoc0KOLX2D
q4AgpibKaEdjKeYZseGLkavgIMe7wWWQZVV7NEuE8+mcnKcEVpvJuhY5dKC9rfzb
z1+ZFxYKb5ZCDhqbKvYEoYrJOLs6zr2jzxrUgz6GIuY+9Y+6LdfMBaZO52GwJWIr
eY9nFRLO2r/7reOCDcekUzybi95LgqEnk1qpeO3PwQ5qS6eHtxNS/rTw6Au5ASkR
vNYgxWMXbWVFsEt/p/iGLUu3G1u6gSwF+DovWD9MUm4=
`protect END_PROTECTED
