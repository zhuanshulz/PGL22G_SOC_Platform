`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qOP0sXHIyaeROcMZI1SPxzRSUBNBaublt47aq476ao3OLT8bvl09jOU3Ye1cIJtW
CsK+vcDiZOIsey99neGEsLuZFiDGAmwmFrZyE8Kp8wXcuV9IbNc+GVaEPl1Uy9vk
ThEPTTv0zSq5TVL9xgNuq076iD3J34g/Yxk+qSOLhS3+kho2SYqwff67fNnyebVb
IA0L6qNIGLrY0UrWJ+Ub09jXxz+kOONAmqy0SFpqxyTDNmRwhzSzQrddM5tn3FE1
WD9KAtYROTY6BWuHT4b9xyG9PTHpsDYnRLX958EpT4OnfsKFpkgRjHFhG8KJKyJu
slHmBzoIq/NMeG7UI06N7RC4B/0dXWBY/8egzfR2RB6kdArwEdB016vfSWd45W4k
MVTkwJsiLPFY1rO3Pm6CbN0or/u2l/B8gcqdkgvavvBzhV76Dj1smKg1DkKlNh7r
jNIc2HXwPdDyE6SVynaSJ0GQTQZIVQDdhtzI2CMtICun/gJvSAqrvkdjqXbNlT7Z
VgGFWgzCZYRwGOOEFPEd/NKD7N4SJ8Kd6+q+KJvqDGhb4j/PlBIMWD21O97JUoXY
eeyfClffGFheSx4mvltpgFsxIb5tdzC5UOC34xcdIG39yHzYIa37iAwBbymCnr1l
sNndySTjO+w+Ii4EItgf69xUBJpkUOyJEoN+fs4tVivqN1SCB0ygzIA+3IksE0wF
oVCs/AYmkWNaT5CFlN4jlYmAmn8m5v5Zr6+pgJdLAkRvlf3q9wyLMvmK4y736kgl
K3ifLs8xD3z3MLfcCjos952ARUZqFTpg4eZarotOhJVtLWt1QGY+Zpf2iaUOHYnf
EaqbQFooNKIAKHxrjUGcTEib7zEnC7zuExQ8Xwkuio7czjJWzWElGqwdvsx0Vz3p
FItIvGZojzv99lqbb+DdpKoMTEI7oAonbBL+bWS94oLbHycDK0LYnKxUajYvmxOw
pEQ2C5n7Sv1xD48fVC2T4jv4Cc6aIc3wZjMs1LJpVlN9yiWuI2zAQQsInvZo04fO
xzr8b943u9YlbE8mAJGSjTY5MmoN0E8Ssrgo20fSreN4J7+FTU8MWwkoTAXZqZtB
tfByXrmqW/AERTRBgclByL3hKbxrnykTrDXpg5PdfuGCgZQunfXLHNVVgP15hvSc
GrFLiP5RYGLQu18LqoZsxOEs01WFQhgC5pyDGswLZXFVkawsSmZIzwUEWUbrZecF
ta8lAA2j1HgulByy7NP7nLhy7LbZBkGItlX9jQaiYURDATqB7b8sgfp9fEy/7DHA
VuKmc/8xQrOpifOFxGQH8ibkKJwDQBzk8DkK0zB9dRf2WFK8pJ+btUluJb1is8Pu
65BRoMd/Az6e/zZfAA4w9vzyiz3f09YI/BlLIFR8mTeZ1IDrcnzZvV4Isjou+bvf
oXOyGgWrAllPezS/UYvHK6Dazzck3TFFWWZ2lRUaN7o/LQGvydLSrYbGZRH4TTPk
OgYYF1gAAdogpSvT77SudpdDpk5R0L46+Fss1I5aWi7o2htzwCFqXY3X20Zbr9oQ
Gpi4N6bDaDIMTPkX7lh0mPzIYXPoTtJ62wEOuYUE/YMwcTWA59y2uo6chWliPjbp
jGGgrQIwBgFxyL/dwF1wkPI7mWbCHkN62cSuH9uPkNLzAz0dQMYt5wNTe2IPqvHQ
BuNSHC7U82Tft+aEKp5HVpKAjsa1z9A8oHuw2RZpYeO2F1BNE3olLI7PlQvi9ygB
K+hc7L1mlJoocs2k80/8W0PBGe9C4GsDn4HmGXKOppxbnhlRlZU5OEm9hSGfeu67
t2zbEfaD1h4Ti8r2qIjDGtDMkgqcOAKipfHePUy/q1AVHl2CTJZhX4j9FT+Lycus
rVgXES7HLtC3bASKNO1kl9BJOR+mMV06C6ZghEMxVDzeUCmFERbcUmM5LaQv+w5K
GOs/gPuwe7P79bkh/+ep8ejJaq/1MMEHQtZqpqjvo4RIZAk1hNuJ0XwgzEDDJP/P
PZnMGf6OY+jqY7bgcxvj58pq6fXn245gmrjEcPfeMQM83U1wXEPdwCGMRElGzT6K
yziE+kn+tExzAcNINMldR/6DISfztaJLxSt5nQPdNOK6w4ENqk92cNUfhcyIGjxD
ij9sLAr30AXPFMM2OKTVHHSGEMFAxBpMB1jL9N/WDSNzQDdemyVDJOP10PGXJWOu
wg2R7qNcGCKqxmzXyQHqQWhaRzHk8CmYlGPwMm3LcG/5IUOn4+hDdBGeM+46jwDE
6kf1/QJEhq8UO4GPFVEHNCZ4j624YLNei9Z4ZCDBZ5/N8fUe8wF7P6ARFzoMVHg2
6pTY2VGfpW34VRRKQlfZk5D6VWECvNTmPBADGROK15vvSwsDxp0n1e/5rn1XzjQ3
uavzJzj0eQLsTv1e2FxtTaci0Y6rP9oEbSSb6AmmZquNOr0GQGzHcYEirjvooGej
mcKNvsViAH0vsEVfnWBH9BbRgw/uXi/aPAXPuSNZFUKkUuJ8C+O0padoNvobll/l
ZdyRIlFE6KfEGQbmppXotHwUjujpH35dfXQukUq1IzM4a1bi1en+FrCywUgFzF7x
/9qPuMM/3R29OxSESVvBum4OvcdQRE1zxL3zoEPsqO+4cme0lkLHq7YRaPdAedtF
iGf/76DMJj/ey+V4cBt3GoqJFCGQLCZmW3WtR/1FvUsnOBQnZBfBcgE9La7Ccz/J
hixUrsh6RVUi8hhD6sU1CwBlky9bpHYFS7jWArP/c329a+NyZdbJacxLWImxldSu
XkISJgxRg18LIhyqDUux5jU/0bNEmZ5Cw68OFy0trAjpEV+UQ6P5PkAKrxg4XpaU
97g9KoVGzRGJAzvDkCV27nE/Cl0VfO6suum4nst61uYFJxhdg0RB0WwkjTUdr8V1
RkkfAtiJ1952yMLhKxM7DAv+fYvlGckFxEnGH/sMlsH4RGi5cHgwQkApRgUwOu8U
iwa/k6uGRHi1WxVajXxCvyUz21VsdsS7i7TuKEtDVAgrhWOEEKBuucT23+VGbYyl
QWq6aWq9HXVcjydfppfDaazf/1v+GslBTXKtdrHf5IwddcCv0yIn9HsTIRH6H1nx
gBuUcCKR7NmxElEpBIuyNf0RAr4s2vIEGJ3xFY7xVQEqL84aoQu6Dt6wIJdqnu2/
+gSeN7ISla2dcKUzIeodOwCIBwmaJgHG2/vcq5TdzmCttFjEfdVmmGK5YjyfI+RZ
`protect END_PROTECTED
