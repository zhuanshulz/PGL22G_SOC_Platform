`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RmGt5u3yu2UrCFRbVmsQEdMXTX+W/NPEH0E9m0MgkEXWx7h9VDvu3zV1ptzZAXC7
qeyaaA8BWEXyL/ZzpEE/aFLu6+6/JfQhn6iBF1E8C/dtqf1vE2HV5Enssv6DxaF9
IAPJjSGwz5eM3JA8zz11kR6oKQETMMYiJ0bVZXdz64VPL7EP2oZsh9j/O7kU6mZz
h5A6M1DKn10E/JSLid3QyrDK38CEISJ8E6eskJORDGT6lWP2nxywf9G4p0manXwq
9rTMvV2DofTlkrslSdLLziXf6HbDmnuR2mVJjk1T/Qv1gVZU6zm6KbfZd8F9LFyJ
8+BDYD1EcxG5gkgunodxt8uz+IBfTr55F10TwYnPchmAwObN77dYknxySQQDcq0T
3EKQxJBsoPmJj22HoT/NUbnOZYRIg+LpB96p73GP9SDKwsWmhXiKZpp379oJ+gDg
TMgzUy/xMYg+/Qb/TVew6q0usJE3AnukZT+/9CawUkBNx38R5BA7IV76DSTIfrRr
wBLwPiGGopkEwzy5KI0hjOirFVCzkXXWIdDIA4Aa47axNOs1Q49TfRX6K1mT9mud
joXTu6tL7b+n+HPrFZbK2IOro9M5L0XIyT/vlZhv3mFSsBfowKoNeib2tzY4P2Fu
Xm9gMAyUN61RSlZAGDKygxpfwRgqsRr8z+H5q2urbYHI1hK7sXb3/PdRPIe4aFrt
b1CgRt8xRRYL7HLtyJJR/S8nn6SYRUXLzh0NQH+MIfTt7nDSzjoRjA0QLBAc19tt
dpEoGAEHSfhwUZrvHPb2/RjWqQUAOABFkN2bivyoTe3T6jUHZg4byhmuDhq0jhmE
KGgpSEoE5HMoNP4ckJNB0A==
`protect END_PROTECTED
