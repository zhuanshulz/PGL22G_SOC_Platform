`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zxV1lReqVm4j+gCiAhsAxs7kevRGWt20sTIa1hPSAk+8+hk0e9sOxuKe8rDovZbt
Hg8tx4t8FpLjZ+SEjIkIONxeyLzNc7AWl66qrBEwlrHruZ1JLXkLoYYKPN0HhQUs
n2hcOH9lXDV+M5PK4pbjMyfEzKBoRquPu8pypdgcFfTAbz1N0JJAzCD0uy5+dai3
tlY1HV9gmPVGgYXdgaGQUjpg5hAkUvBkonEr9xvIJADuG4T2b28d1Mc8e73KskZe
afdYqlDKMIjExoCdJY2h6I5ng+UUN2cnN2xBVqQRQtpZurXS7QinR3KbGL9zoEHe
jlUZ2hG/Y51qae91G3/MEQ==
`protect END_PROTECTED
