`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
50MQOtp42SFdXF/BpOecRc4m1yqjdPzSGAeKYxyxh80I5wLy15/BpMWRe1tWFum1
wmVH/u1WyhfqZC7Cn/BSn5MNw6QIDYJRt3spOMFPYCr4mgym+YpWgnbAEDjGOMvF
EQhJBWIZj6JIxjywaknY+5RfKfEj4GLt/KQ4FcLdVHuAJ2i9bjZKgJoszN5+46IP
tpRq1FGu1yKSoW0NrDftRkFHkU2Fx+FQLXCcGP/Ni1UGALmnNWWEa4oujvemMFtk
XEqd5wh8IqfVo7TnHvEg8XNNnynOKx6vxQTWA/dGZgIS5e5vx6oDYicMLLf21bBL
YTpLCcWtCgSEvNtTWXYjhO9d0bwbKhGoKb4upBqdb7iY/pyxLfFSZEfPQFR6ccMl
YfIZ57nW1kRT1BGbUzivZLPq8jFdsxIjBg85vnkxIcIBLUQE+N9KXirSbcsSqkQh
BmfKhHGejJ6ZH635Kzcce/kN1Wb+n+mTtLGKdCaMwT2GAsgRVsmnuIez9HZIXS5R
PY8wEWXB2b+xDjxScQiY1Y/UmLNTkhIV5Rm+rljZX82I3yvM98rDPOrExaBmk5MO
u6zj0XVe9Jfrtfh6RMYiut3Dn/ZMv7MNEvj5F8E2dM4Dt5XyQXIPWQbhx398MsXo
43Z+8kDGzZnT/RszJVE06wFRyP+JALxnL5H6XGcbo5d4sYdB/BuV+JVoPvEP+al3
vLwuDACGTbBX2FCsDsLzyDGcbvwSsobK6XkjttrSHg9LT6pKFi7szc/yjNkOE25F
jkutf9u5I3g4xM92YggO2tvjG8XTGm4Y9Y2i6q65oNTII27lcDtHDpJ3LWvZACOS
fY/ov1pIgwF6ubkhXKI1fU9ePMhcQu/iDyyRXPQRG+CAHZNG6lDchK/EhFCRKnNO
auuMyFaFtBvM+x3lS1rhr5yKeHOPq8/wDBlLVp1v8Ce9+toLLyxuCs9lViOOShmL
4KmYjTbE2fVs0f64ZMUKzAaq3sdrFao9C38iJ34ADYkWUNKxWv7IeX1H7E7D6FHa
qO4KGdmS/SnaLV8UjwvY/oe/YFZdlUGav9VQ+KCRKxSTVNPXPee0lNq5s4a37gTM
jJOmLbxTEI1i75TkW+9MH1AU5KnJlVlnSFptdNnNSk2/cz4r+fpMik7FF5E+DmGs
8XjX+y+VGvToQkbil9ifZqer0ujFUYy4ju5oVkFuKxN+uj+ItFWfkFZobeMr+tIH
lG0TVS4Lb6t8ZjZ5/ZufLYogjOmiUXsE294KhQ1etWxC1jugOsDjRsdbHtyDQhp4
TJgtXz7KluoQu6O3JePeX1TzaiaA4tQUI2K4Pm/DivxhaQUDdFOEfS5NaVeTyFSr
zV75et8+5bZgYF7xrT+kLuIdvGoxD5tvcl+V1OO1JEPeTjM1d7CwT5FUuZjHF0tp
kSgak2IkMuasj+3jhxQjzUMnSJNs35aDL8BqKi0kR92avHdqayfqEY6yPihDaODn
eZtnTCPn/JU4+KSTNCdVSdZVzN+JRz8iPrH4QVfhpENHLpxc5vU+5e2CGxVJTk5F
rCAenjAWajYmsZ6VbzAuslZI23nLfScIecGUk193co+ZcQhebqbaHykW3BrQl2q1
ggfLK257ND/rroC78vP/dbCwADa24p1BdM7JK92iCqPx9nk4I+n7hik2Eca1oIAb
36YfoIq6sKSz/2nn13yEVelviZsVF5UUmG9ncYSrlA6X9MZy2JRzlVOuLzV+n2bK
bqdFMAbd228/nBrcxb4c1dJ1S/DoO08aC8OqnyGGrA+JKohHVoyLBO7YmhDW5vuC
CGrq5FJRoYe9QaPaq68r+gtXleBaWzwL2jA2jmMNs7ok+5p9JDkx8fZVDSFmzrSR
ysqYbh/r5cyStzFaLANfxiHVvO1GRQkyL5WivwiOPW0kEmTjhUILtBRwEUvj32xW
RT5epTKkBqjl8O5Mhk2ISMV549vXwrsBW+230TlG0wzvX86I6lYvJtJshqMNhqnu
Z0Ua98p7fIeK60yTZR2jTRVdFa6Itk3ezrg7zLvfrJIpbYv54/0dbrgCyMha4Nn0
gn2teBuLTeG0zLm/t4wOlPMHDMJjS+o3MkceworYDAXUwmbp4D4TuLsPJfb5qJyH
JXVAcIJy5droLp2TYrfuy+ioOeJ8k9VM8yKDUFjvhsrKY5Xg2D+AXHOCZrgb9Klp
YBzDxaZMFL2g/+m9cc0bAF6x8Su/wYhqaRkfVV2MeP80XnPWVSgsDmG34F2NJfYu
wr9HbgO/rqhALRmtzMlvFqcYVwZO9vCsJIgvDN+tTblBdFHKoh+HJ2SuR64xJ5KC
HozFImm/po7B9pezVFXZC+WISVJe1TGWKYlsXznSDV1vJ/h0JZiKN7mwP3gY4rlP
lhp8UgDDx+zppQRGx5z325gvR9O4+12AWvlajpBa/Lv+PPHSJlapc1XodpVVF+UB
mCHKPIWbDvH6jBU2SBWnh1RQigQ6RMXNnLoTNCtOlF0/YWrUhOBalCdpljnpjjPC
+tuT63aqXsR+aDBnshZVm1I0cVHicuQGA4vVS6X4BYoTqWKnEfiBbI4jKBBfpMCU
8gCM3PcF8BL/Xi5/SlwN6wh1z6EGq5dUYWgUVpwEh3Ugej64dHatl6hbFLEipBGm
K1o279LIZVQx0notpIOrq7g3WG87ufWhLOJwGOVFabFGptDJG7+dlK1Z856TyrOS
j35vqgZqYNOA4VtvyDqbfWLgfxDkHh3RyTZrmSB1yE37ys16+svP6RA0HhKrrDGF
G5SBXYv+xfwymL3OlSwvNkh3nyGYech9u8uHncZE0L2uaFYCq2xlJneiUgSGOskz
tjkjJKcib4hTS0cOAXGADhfNAvNbl+jBLhs5+Mfo2LXeTWiPtkmZRSfwoH4nWx2d
3BhMxe82l60tJjC0L50hvLrBOLhWjW5gHK7cCgg+M9py1bq6ZQQnC3FhrPiXgM7L
1AQ09R0HExKOA1L+OV3kEc5u2rnYd8bu+nxYDq1UwJGVAUU41DXT2d7qLgVkz0Fy
9ZpUToWnS8p+mfIz61v8rzpLzrHg33fc4knvgDRcxQiq0RxlOY9hXW8nOWLg1o7z
MchaPrJD8VEcKJZp6VsQ7rUprqgnpQwtt6sn9RNt5fqMlgzKfAsf0fNUzIra2POo
7gtDTOtQUBMexBn14NZTUvx0K57C4nSnvkIdcdOPLVZfaEXyRFaK4S3bdrG9z62a
uq820uou6FzQOFK/XZCLNYApBHiTFOU4NVU35V+OrBYFtisoGjLYqtoX9f1dvb/5
qSuTBOt1C6V/JGs+LF1VA1REc3RGld0U4kjhVDUtftwCUsIoz9DNMXJV0h39UgMH
I+nP6iPTp49WloIVlJrmWLzcbkTpz96lv8OtNd5CN/LSPyiJZF6DnUds6qj2rRwP
axLp9N3GmEn5Y0v4YvaZtPhc9kBRNdEH4aCYCZavF3FdjjqpyXHR82h7tZ8+Thnz
TPTxXcYZj4kkn1B0nROSpb15y2GlYhBtkjkUp7YXlEEovlFoN+B5JdzqbAMEbxlT
ELM8jcRB8CQ8A8G+T6DTygFRbHTuiI9bdCKJWwbgOF8zAkj6EuA+AP+f/3bHXyWJ
OHeLVz/vvcnm+bcWY4Lo96V7heT4QFE2AWVJCWw3RLOSAfCKKNe1jIH3DHb+qCiE
mtGxzv1X34YUywzBpxFfoPENkdNyiTOOck5rrvH8an9VnfzWYdzECW10NbsoGtV6
J3j2kJ14jUsZwndAQevEgqrTpIeSIjHD6zbc9JLr2k2kObC5wKdDXy7IdQNPeHic
ID17SxVg2FKBwC7nhiEYex42ydYlvNnftwepUphEwbjzNsWvpcC3E1BSIR/BMbcp
JKC9nQjJvW24aN9vkSpy2F1sZvOFKEMYiX+BWlYlmuZDl1XOfjBkgQHDqHdaphMH
vlfqxpYM+YfIbU58mrMvyRKdshNPEtvvQ6M+QllBmH56C+86Vz08Qtl61ebMQkNA
U4RJ+sJtT9+/csEqRs8XWo0OuqkrVAask5wHr/brqX/e0JXdoWC4+n8DOfSclNUr
J/pqPpa+cKOCaBs0rVbdeakmQbnZ2Ce1mGKQVrmvrRLOBetPMgNwEdnt3vP9Iig6
vAkyAvEUhFYJgeN8KjSR6U4Wunvgtx+1T/umA/QakbrUBUTta2M1xzm6BLey4MTC
qwyYwrdCauiccrxgibc4pwmVarmpeq8hOwSnVPcmre010wRWZ9FPTRKlZJg6C4IR
LfqJUSFoNp5l2y9z4yMIIVpZRVstyJAJoR6oVP7g2zCRxYdy2fBNUrw6FXrLrxkN
AGm8V6b6sBEuqXTY6FyZwGAZ6DEnT2cK6hT+aMVefYZZRsJNxGO2nkPCJpf4e8km
THyg73hdQ2bXrt3C8xOcAYi1BM8uglbW1GlNr+YPGv/2JY6KJboJRjym1RheQlPS
cBiqKN2G1lPM6C+j7bDdZKBaCTV1MJhunQTybpdxRlrQLd4Q8R4HBDRdchg5ZltV
8T681v9lQ8Plih603tQZHkyovGa7jX2E+KVdQcmiCkHcA3eje0VlYSR7K4h/0rMr
q6Rz4ZjakH5Y3IccwoqI5bXwmYGYO1ujkD30Rt0fHTICIOZ9dl0/gbKlzOeaSuVJ
St5Y0YyT6uQyKdQl4Jv4FkWIFFh6s71D4Jf2AWJ2QROe1dJEBsK4mJE5FTdW+tvl
YGxnId1mFmPk6yXBZsSOTk8bzRdYx1FI5eH9uJCLuZQCczBl85gsnDoGZBlnyIKy
m0mGwY2WCo9/r8vzY7+9TYUNSA+S0WbjUx370eqjBPN6D7wERWHbw53Jr9TYn4aK
EykPhd+5cOACMqHgUV7wWnrkPFa7CRJIvUO6VuNe2gm1PWMzGIwiIjwRFX33Dq1z
hGYc/nnFIOpNMUVINmitHlsj2m01ckGIrTgx/SBuM/JU1Ddw1kHKbNDv6CMCwrnt
DWUV27ETju9lgFtmkDf6gVL7CUWcxEZlQ/YY72E3G/BHwh6PIZta+nNv3LwwEvkb
01XcQwm6KLFX7G77AAU52QbDXjLS0OfLkI24gyoBVXSikHE/eIM+cf00bgY5idVg
tVRty31I4sNDLPrqFm2RcPVDwYzTsXg7AjmQR9GiOh1GTwrwdsV2ElD//e+IPEge
1+43967rhM/I4ROzJaxu5EWOxk8iS+j2sI9mn3imwuf2WdL/+68g9xT1//oZLHwY
XFQQFxFT4HF76ER2gWVSY70BlKRuqAGTFaSoIkrPj2rXNevwdw8KKWWDi8BrX+Lf
uYomLpEd2GVrFk/Kb/UdpX2NQpbRRcdZOaWGLrbqQv8xyYBVB+2Rqmjy8oYkPelP
tvp3HFO5uHsnF98n4D948crkY0eYDJwIfFgq7t54at0=
`protect END_PROTECTED
