`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Olnm4srNSLD+NtKUH3wO29hmzGwwPnnNnsFuI0J1+SNED8VBDsL17IPz4Hm+6OHT
HwEvj44uVFBuQkI7C3GxPfKnh5Uu/DHyUhkJzYKRHHzMRcotUcMqUdQXBgiUzrNI
TslkjAJsWCL8jlWZTsWcY5ND8PUgmWERMtON40QEthzsEr5V5sCqQ7BqorTtnQnb
NFd8vW3BkJNwahn6K3JnASan+jvdgWklzfFqWUCBSq8q2Kq8kjCPl7doBC8IB1En
glIzGFgEsQacWmx6yC7zCKvewuBsvUJc+ILTK6VxoIng1dPFHSzNjEIXdsBRzLZR
u9Sk4TJKO78SxgPoswbyoiM2JxhWuSp9W65A/8ekbSnnI+9UbKzKPN1y3xxz8Ecg
XxY87X8e8a5EtWl2ObrHbYBJwAhHqBTSS8/ykOF+ZB0=
`protect END_PROTECTED
