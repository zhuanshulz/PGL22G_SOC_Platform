`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
liOEMND1V4JD6RjO3L/Xdtnhkq2dYh+XzWWLMPrflLwYynsO/we9rxxSFMEWJSLg
ds3/jHqYdPi2l3vQIYr9OV9pL2WZCeThK6nD3m9763tfRw+cp3GLyWnupXtUH4+B
lbjBmK1kyGtMLueepOLFeuF7qK385sF/EwNcQQZgzZNi4g1gW5d4+6mwhyF/mno0
mNfKTX5Eo1dZcUswMGVQ/l5DiNJPSJ9yNCQpaNcyJtxdPKWgWrANhcgW+dzSonKY
thgSRWxZOYgeu6oa8b3FBL7RCyw4PmnOOU74gzDkQObn+14rnvJm+YCz3EQgHEgo
aB9aWV/DToBuXMtUUg91Cpggd8dodzb5dNxwxqF1s6zAlLw6Yfjyz5BbexukSLB8
`protect END_PROTECTED
