`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FW+jZeLpTXXcsw8ZFUCy6F7XMPvjgPP/TO0ZqZaRaElp+YSBTPQalON6Fb7C1kf1
xdYCbs1SD1iUVqHOUN2rSe/JyjjE0tQvNIDZk6xJhUsOFLjal/pPLMF5W8bav+r0
O08B1ka6SuNcBNgEW5PXI/wOwubrR4Q4NU074tIPoW9Q+36LsgLeY1xjUlpC3Y1P
eMeZPVsvTUKQBmTBUF5KKLbQ5h3f5FZIKF4RAuy+mSBg3KWdgsD5FOBCKye9DUoi
SpJ44x4lTrfJ/NgSynRRNWiPXit0/N4FAodLpG5NIfltH/+gEQ4fjUw5DCyT5KHy
6x69C3lKQ5bHXe6UJ70vqh7JaYR9dv8emTOIeavc6QcAm3nrzFhOGB3ky6/SYek+
XjhZy90VPMNInF/prx/u7cNnoe09pYscQGtgCm0NVrEUhmoSSVmoM6jJC83GRA5a
D/IoEIqwmQ7i8UUCLNEifhA7+5xjHoSIzKl4+XdvjylTLnc+Qw5AEykXBkaLapyz
N5+2U/teULuB7x602wQDwN03TEWLqZ1GJxzbgaw2w/uaBOrucbjUJkF9OSFog3s8
b4NRXU+4n84hDxtvwdLPf8zGERlSTakyD21viiqP4XprecZidz0TI/16MWiqmOnb
fzs5fg/n5jcahWug6ZR+9kH9QJsljTdzrXNbaegoXqbsU/rBoPv54gw7k+nQqvX1
rTm/RV0rbsRjXBrJRK3szHNvh76gY5uXwVE/HMjyb71KUfFUcTJlPvuFxUNVIJSn
0DhPLJCspERMNx5ic58/PLZUr4VLUPHf5c+CVj1RCTnRTz/gYMqLVPbB1eVOyYaN
OLzzKkXRH3JOpiMXd7x7dXs/hZauyFcHLFxppU2j7a8BCE0vp1ZEZGPO/jGs9fY6
fLNIiXyvQXL4BVzHQuxdb9dS86aZAks+yT6dd6tz90psTq2IgIrP+YcV2FRyXYee
BBPl4UOA/GYtY1cE5QQeeEqmHtGyhj4lNfHY1BYpPXfQCoSS4xVt6+UV5gJHvkdg
8cgzDMSOhn6s38MNR+Og/fvyontVuThV7FSj0qrnPc8ShFHJHwWvXbJ9TpBd6est
/NvCYLrSKRIslkbyVTRtvzhD5sTJXGLoqtUPqDmSmCU7wpZvZQ0sA4ztFKOwReBh
tsEgO7k5I+xDtXNHPvWU4yiHHTWzhOWgwe2SkMm9BUpO0eASKa9j2u41trmruqmq
Le5v7x7+tk9VPeOkOwnIwi9QzVdsSPOQOCr25fl7Ta4X9f7C+MA1SuO+w9RXolHi
Y7RmCkmHSjNFx+HQdK1N2MuQ7M659ZG6oW9PA1U/5HMFRQ/MTfrhW/JwPHOhoo5t
AcaZE6xnMDvqj8Ec/YMHAVUCJGwnAXE7hwt7xo52NL154uCFxILXjC9DGWKskQEq
/7SFVXS3p568M6JIKxE8XbqdZXDB+9hBLjROddnV/YQgE76rKR2jabbJTTW3BKJd
CsWpw5/YBpWsFCLX4xC5pHqGinafzaSXyIa2JRtHeyISJhJPIEFZaawzzRwXmq2c
ruLlDe3g/VBMg3/15Xvfsr5MJDlmFmL9Qqej2aVzXojcbIzTTweNJJZT6V9hessX
OwfE5XZLfG2IFmBXU0tuxovsqOT8SHeAcuY/nqm/ewKFJult1NdcakgUPlQV5+Z1
OeGkfiYFzs8T4Z8UMtiZGA1WyNIZqBL8EmGAfxweAFeFVVG1H6d4hRX0hUewwtht
bRaX6XPor20RovKO1kmcFLt0g0JQDyAAb8fVPvzT2Nkr6LQcf2Olg+IGH5RcOsvT
dAaqoKa2LBqpw2ycgW7uSCga5TlCH+hAcaTTZ71S52L6qgr3ALTDa0LWc7Jpa7rV
yIqwiCfcfVr+4EyK9Z2VXuuo1Rjvn9Y1bmhipUmkgUtjiTftDH9YxTncNfYnoF2/
gA8JSM5mTcbEQaqzgG5oZ3noYzsiZIyZCNRXRNvWIfF5JjkUSsP2UI+25/R8JjfF
lSoNvzTsycNeVD5ges8yNoy71hqv7oEmaiyjcoruCC4wtmk+CHEZ7nv9hP453Waz
VByzuQOTigRIC+WP3DtzyxmAlTORmc+UNPErIIfZqh5WndowGszI9plFq/+5PDbd
SeOmM86DM2nJJvB88u3o9Kqp+tpfiyoAD0f2JOmVaKa1qMU8JW2iDFAB7eGgfHFU
UwSDHHSOw9oZIB/El0UGiRwJap+lKDpccUBAWwJdASdQoJhQG9bBKIsHldtTV9xb
/z1MzrIdG+Zcgw0Ck/Uj7gcTfwpyXHnJ6Wg2Q4eaNuZuZRJRlrjhOfa2BkCBYPAV
nTUbd/bsA+12/8Nti24BkUMBcmTryeiiBfW/Zgt1w/bSCrjJktl3UwCvy6GS+LNu
1scHilhH5tJHj6pjSc8vMkGCUP11EbBG8EPL4JSKpd39h63lwX76pNnAWhoZWOPQ
XdyMYBEZp6bWZc79Uti9A/DVTcuMq6rEryrq1y16Wvj7ffNAq2xp4ZAACT99N5xm
RB0kLOJCP5i+iAIF78I3GTg+sA2mLMa3ucfZhIqqKlv21jPkIOp1gSQjGJ6bDsd3
Q6Eolrg3CaWkxwBcdkJMaMRV97QKRUbi07/2ec30nsS4NcYhAeHPGCt2d9k8/NMp
l2oT25fibGY/wRoPckwKSimdeIdw7lRTmzLW3SnA2nXlINZMpQgIX7OSYx/UJjci
7o6ycAiZ4uI442M4nEFxHedvjIRuP/31BVUhMCxqxpn5wyJcM+Pl32T0NpwvxiHL
RyRBpChVNNGbyc3K4rQ9BGss2R+m9a53izRQ6uSIozZ9C3B9AGOtdKqGITDHivnc
lBvkMfLu37fyI8M144HTRH1LfRGN3BXNIonneT6lpyhOB3G98PJA2em/jvqTOoN7
2VsTeBhfCfF2S1dWe+4gCP/sMUtt1fn51zRhHjNRVIk1f74atCadOvBMZ2Dvs484
SD00IQWGNMdLvMKzsrkWmMKCPSbAqMLEuT5apKYzLlqEOxMu3GP9YUe0fCSprYZh
TlykigKizl4C3/TgmOJp7LxZ3iaEE6DT8vNwPsyfLh3SqhdHZVAjV/IkNGVi33KS
ycMlAZmXflBumfUoZulZcRtS4mnTzHfO1CezaHoAjEQpOiwd9i0mJD6dimjscPXH
eCDsaLqGNIBsySq1Y+K/tKvrpA1MlP28dAuqdVTmngPuGcRsapJAgHT3SQx0PJRz
9BheweXaopL4TyS3/cJY2i+1oLdjUMa2FDYA0KQoW8HqKIQ/NlrqcuRFz954/Au4
ByX5yODm4ZcRY8x//8DmN7kESeOUAcOZTK5WmO2u7il5U8W0Ny0Ou8Ta3rjHxFKS
916IHEwAohSxPYhWyXFXaZtqolWfQYP4cw8+8wHwuPDglCBmClTNMnJg0jt4shU5
ZTDcCNl1Xa9aAvkJekIPGIeXoVLPEiWiTD8OPgiy5xfFTtJRTmOUdNYuicQCN/1Y
A5uvnsIREDWqljkXA5CVOYT93PTOpQqxQ1PP/TlkxKkIxASd/7/Aw1XWKeE/c/gs
/kxosIEO44b5UKwHezNQdw0pDM/AX2ImzpymoCN5RM+3Ar2Ex0dqXrujcVOZHKO+
8vpGjo6gzi7ct/pP6vkpSbCyruFzJDulceti2i0vV5iWjH9JGh6yuwHAluEpx71M
uAGmyc/H6YabUSLRdqNMdz/3xNu+LmSJwCoGz2Ku+Zim00TFdAWhr9DwyuEZz8+5
W81PzKxbbgiNDdEV5Zt64Fm5wsBtc3kAcscpA3aBXB2oy2SynzKxFUkhRVTGPMr9
xcBxrbAQmcGgaVa8e4XO+/jjhTWF9+Gwh+ebNMnZSa5hzG5oG44gIw9QRFOoxMd5
21WB5mPP3KKop4AAlgKGonoEnwa5nm9Pod/BE8fifwbMLnKL7lyw9wVME1gLlPjj
N69N1MDZUGvjCHzV640zNjwuRHj61kooVKQywxliYyOvNT5nkYqQEcvGQcLO52Ah
gMba6Fjr37d87bVaqOrjv9VfLQDWFGMR67FuTRB/mpxSldYmS47graIoV3/VUmdA
2sFlKF9gKZuuKm95ndMsY/9geUu8WeHwcD7TfZ6hTVmIEKE/AXnlWUke7u89/AmM
s2j/kRGBSW48Sdpk7wlmIoFu5W1vSHiuwodcyppq3LG2SsEBGDs2qjy5elR4YKzV
gWJslCE5W6YTnwf6tlAKddigYnNyV9nbcAzglCTFN6thZzX2w5EVnym42Vh7ixBM
TMuLCxf2dw4z1iAYSXRfZg18cU2eF1UroBa0+VHS9BJDhRcDA9jmY0rF8GaFr5tj
sFWxnSJtIpQnYEBXzTYpRnmoXLWsX+fcAcJ24jIuCOCb8PDXXiMBRUXzvBM2v5XR
cpzlhzZLVk2RKc8W9RRAFlkgpUk5QXk6AbnnPtEjCxJbSPCYJLcF9SBIbhIzHG23
jVv3L+Bv1oCPpuK+Um9P3XBkqxIO6G7zKFol1SrGNoc7VnIoiPp/NLsm9y1xSYde
BVfyQbrbLxf+bBz+L2+H7+O99ONqSkk5jge/vPKE0jdWtDxxbWjh92X/rFQkhMya
GE+KrSzfLsFNV3GJtyFDeEFTj4PE0nkaEBqgakqE7f7nikKY2yIbAYPJnx55fM2j
dCq8ja1sINdlr7lGIN2nVnI+bgmIN0xE8JAfnQf9koV20Y4y2sSK/6t2B0JpdT4i
JaGnWjTkSr7w6Fh0F6WZQHSEqzeo4uqOzVb6HVp74sM6i94Ayx38vnw/QYbfPcH2
e22NmGscX/cAOLmKJ94fmz3MQPa5CRXmhbN//kr5GdlFg6TkgElrFS6Icp7K4QMN
3rauilqv6xCX4wBMLNmPNqCLlAdUCJCk6BAn04GldWo1lYLWf78uqaH404hzE1Ko
CEAoQXfS8+I9qS3ZObwd2YZVnHr9HVWfzNBS2a4tG0IVCC/yCAr0AfFTwJcduLv2
W6AkN3Xx1JZIEoR+kjfPEn8xWbN0cZ53ZO7XIruLIijQFfsOdRFLuFUpF5IPd2au
GnlZ4tHN4iKYpWd99XgWmJJQudC1+A7N2hPQL10PrCMW8d4OLTQkqQ/fqXrNjDqm
QdCHcGKnOt/Lwo0EluzjcMDrU5isanJNP15Sj1P2KkhHajJTy+LkRk0HEhpF5Uib
hSFaNgc9zlY5p6VHfFQ0SjmCVfcxp5Qpt8uG8lATTflvkuNX0PzRodAj4oxMA6Dm
kbUWVdT0aRF4IaxZ8Rujeapa/7KCzV9Dublq6G/qGkkuTia+KF3bDWUwT5mOqjIU
asi2ZWgz1nSe4Fd7bvTTNfa4ivDxqFhjdJa/KrT4d40wD7/fVpjjARnEQvlV2MTK
bcGsQRLJcAeY7vKuGL0ZobZtPB30MHKzLSaBbPla9hv/4fhcdsNPurzxizC/mBiU
PrwWUdroAWMc2qkLVhq3hH5nxcC7t6tkk2p2jF6Yf1XwGHt60o1xpPwfvQaFHDEc
msLHs3Msv/tfrHMTjH8yMBLN51VfP+wF/TjCA0xTzTZR37A8LblUsRmRna+45EOB
p2TvR2r36CRNtK0vyB6sZoWuRD0vOQaqTseo8WYHZnhl269s4qIep+oVSC9FlhBB
ZlWS2+uC9rCV54I/AnlQBBGtWLS6wwCPHxa5V9paFwjTiGZN2PZlOeZGd5k/ChuR
v5d86lD7FFFufec1Y4FNJNPQrTvLJ1eoNfELMvhEW+aGyG4T00ekRRrHgfKXFdl0
1quwbAcuXX6yt86GNH633WSCYZSBvoIFvCRJC2EqQyO6gF7xI5LWXLlU314Eqair
1VnH8nmlzskSZB+6lN5zoTTGYpM2SEwU3IHrrg2VsODr6FgiS3ez3i7qHGNiyo9j
kEZj7Exy6qZRc4esL9T4V1erQ6IDaPqjBPMh8MWfHl4t38cssNgum6uMxPict3IC
B/GfsRv0W5a9F/f6aZ9ad4ROxhBc3aN30E02IiU2Fp4Unfh2WwxAdIr9EmWkFl2q
wjwRGfYtMwf11UixuJSmSVYjDCXDGfWBQzXih3WWyHlVXG8xxBJxjIHiNTUdgtto
fPWXMLRsDad5bIx/CU+jUxbX24WLxpZqlJgpgJ4g+OxJh1DidFUhNJZHVaBGngOg
WHAXmPGOtS8GclWtApEcyBB9dARPo9X2tkGH0We3jLnMYeTBigaFr6wHDqn9IF+Z
LNKaczEMy8J5FdWZOLIbNwJj9q8mgf/ATsZmOAbra8rI25bcihaISamaqr8kjU8o
DPmkynbFEwJOaRltaVrjs1CNgSKE0rzeHw+ND7WrjdcYoOkJV3xNorFDjMp8/aQy
JOejcMFJOUYF3zLiKRoFW/WaCmN6an5Kn5Iu6mpwE8q/RRq08vQc6zIvUSw3L2/Z
DmwDyPfO9Lk+qw7hszNusqshYC/axICRMmYy+BwhmSZzjc4zH8IVOZCP8EYKcdrH
hSZn2/iJ+Zg1TMDBjmfrz3O36KuzYfyw0bISn9AzVT8=
`protect END_PROTECTED
