`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FKEtwUqyxp7flbAMYSguOm8x44sBBajaTopoTuECA1P/XjgMx5Tizr/zO5VpVxEV
S8tGNfc/n+zvbXQ30G2WbQJtNyEF9IivbWbgTIeTSpz2QVgDJ5nMQ1MZmODCrFOE
AlJgL2pEC7d36nQ6wufv6o2huO9zhEiUYptIX5Eb0E7tt2UScy3vGchd2Jg52uXo
W/EvT9uojSKpTt2rtE15frchb/yrjDA4Vjf+5sjsu1PRpAFOIsOa3Hsj8nTLqA4E
RwufGZHnjm0A/5g6xcnI+ae1HVuiQGLs141hn2idRT6odn7gpxcK/OC6Ll6bKM0H
6/4pm6oyCY7ghVHWHcTWEWKnJWDVchnCVmVXecGaengINnpNSBj+FCQsmvSSdpV4
GQptttasdg4TCJbcWzzm6UMVeaEW690CWDxLWiOzFElMUyDiFOGTxS2lpCikgPCi
1v+Kk3GExWFAGGbiqtC11V1cLWC45BHz7Fhf+eSW8Ni7DQHi32C0WiZoEKeO5CFZ
ZUyXktXx2Wt/MeqOCGnyBl6Nsn0YZGHwaiYQT1vbG6uAdXIg25xbJpdbBNHvYcw8
GKnnMJ0BWUJEa7g5PRnkTPxyE5HZFsab60F2FujVE/ZEabS3yrdKF3nlYRGwO1FI
NMaYjBZbys9wda1rPWMSlSZacvi8u4dMZwINU2Jg+KuHWEGZh95SCaF+fr9x7yA6
Mhvc6p3k+bq9g1wGNrEedwCUlOp3PTdjWVkeiE+FZnsNLDS8T4JIRQrlLCOQLE+B
8h79vXmR9xkIHR716v+SQufreCskAoYQpMlgbn7cTCRWz1Ib9s41dmLHdFg/1MFv
g00g8HFkfiunIdY6xApWqWWu7XSnNY43rMO23ghBqPpu1FS4+esATSzn5uU0xKHK
fZpYwGh9a7wFjmm4boFT/m8maxJ9ZGLs7m0CQPXTCcELrAnIrNuWPNALJfVD6Hqb
eIe8+aqZpJeHAT7Tn/bL+DqRQWMp78oNVOWInzGK0RSZxGITt1+5SwPIExQkCJmy
Yl9c1spI1ZvEqe+OXltysdifX3EW5fkV68ONqIqGPbBiA6vAU4Zw52zKNGtVyFz8
Bw4aWvGH8y+XINjXFv58ymWnZyfvN4X+9hjUA/ySKmJ8ABYUJdRK7KeGqNXjB6go
XYcVVC7GES+XPPcljQthhbVqUXqa23Q2XqqM1gftg6EoV4ZKtvkCPMA27GtbjpEP
GIsHIVZ68Y7SM/FnJ8Wm2mBkJZJk5d9DdsFnF5lMPMwk8GSrsKc27KqW+Rb3Vuce
GxZbi+usVsmM/UE2F7uEd7ZBTi2qRCY7xRWy1nOYxvW4Ds09eXz3gaaAxRPtJn7E
PTuwzbSKxr+buSGtTW/IIvZFN5zs7tDZeB/13lD2QSvDypeuf4H+Ca9kFcCAYcRQ
m5EaIaH5BeIjuqpsTtLxwbeSM2N63XXigc5f3ysu+yJf+Z68VFK1GaHkJZD8uvGL
sLP48y0rNMpK1WvK8PFGXqNqXACkJAWMPkEFtGC0MCyoxs9ZVM3efunqb3igDZ6y
e/SMYq2Qfze306Js/W/hVF95gMr6Yq5jl4gIrkX1SE5beof19KwCxWRt+DnXbwJ5
XnLoqSP+GbcJUVboZ890Ri+J760e/i8O0vr4Fa2cki5Uwla80pxKaacY3zKX7exq
WOBQRvOH6vCfO+yuW0SkluiZrP8vrqqmGmP0V7fdQB0ruSprrK52XnDJJv3kS8+N
ii1nAJ28WCL1zx7jcUI0ecWG8IbS9v0net2aNqRoCDkSch5A3ThiwlJWYR21+yUt
YMfVDqZGRxOZbMM7JfSmKytxd9Ck58tVqH0Ne17agc2yGavkY08u4ArzLuJaM96u
ma+v6FeIacvY4Secddx5VxGaQtcAPWrDBjmIC4gRnMn5wD+w0mHf9uWdieZuSmA0
0dG7l+YbSKZn6NEaiubSWU9dizZTXkGoZHxzWGUW7gN4zSaoNheKM8Xti6wW1SPW
3/FiBJqBRqVngButMCXvW15lAzAwelr0Zzsp7J2zs7k82kKwZA4aj9miXgc9wJGA
EO34kQ5iiYsT95wZKgIgoCay+4ZDaAWl8Dq3ObedbaBLsStowV0ubKwB2tZfsPTN
eKoOae2t36PPnkLFSXcaHsCydhzDuonVPJtoHOa1pO362S4vybUWcZW1wgU1xxBc
cI58DKf++hKw4qWROfuuLvm4ZBxjTSO7ndo61BGif+0Na5eyVoH1nvgJY9/W2znG
z7uNXzSK7SXenLt0gZQEYNPFXjXguoV5KS1egIMbxnJq56xXJhQJaekRhLyY1ms+
QygAwfOFjlqCpJEPMT6ZyOc0JGHHh6oMOEAqUbM6IwZ+RfkjPrMXcLwI4AjPbj1W
Tgv/wBqHF5538z+kgyXhDoJeMp/8/xporFvQEeHmpUGH9P1ZaOTyF4yP9g9mWZIx
anIiRnc00Q70fR8hT/wjwzt3IYw1b5PnPM/5u17KndOI35ZQk5h6Thmrwjp5YO0V
OBcAKL++fmTgtsGutUA4FeEfl8JOFHFE+BNPOKqIt2ZhuMoUvYgEN0iEQAMm0qZF
6p6g8ObSoqBjxFRwbCcEQ5EPfkoJnQayF+7wzEsYTXNV+XBGmNJsyXVxcZI9gUfa
reJkoLgFMoJoW8pYYX3Ufifad7RKiUCA3/SNAVnrlvsXWlfz5bNgGOjxXTeJ/q2m
4Dpurz7aBqD632eWs/dZNaitnqQLajG9Qt693p6795isRYv5QQNYBoQVUgksenzO
yn1QTV8UvMMLjcATVcOUgBEOzGcK7WE8ifSjhH+TowJxzlPDMSu8ffD5tVnPlCut
hl9IduBWZfuDXSJZ8UQFzrFnkour67/9PvhxPWzoV/JYE1xQtqzmwRuL6HuI/V9u
qwm1uWf1IMOfCVggBwZB80RYNj9PM5lu+cPLb65vUwJvUPXGHVxeu++a5q7o2L3/
adhvcYMGSEjl6lgk7bk0K47ACb3WIjA7s7vsj8Sf1b4uEig5Nh49xjfub/BZ/3U9
dPRN9utBR1BbQW+G2CN1f4MCOmdlvdo8QMcHMYWW+DIalz5x7+PNUfCrGECc2xE0
OI3l5ekUK1NHTperLHt7M+9PQ/erT7P80jps129khzieO05GmUGl3v3SO35cp5dZ
UmbPxyLgqNoltI0BXaKdbOVfm0nKTeV92njVLUxt9UWB/1bdfV/m1Z8ieRKsAQGY
S7yzUiqmsnqIMxE9F+sUX3z4GErp2z+o8lB+biDHF2QGOzYe3Stvjy2CKgEpmqwl
gRtvn9f7jcL01xxfbXx6nz3HfO4uR/sgTt6ALLdWeuhMbG34TEQ+y8CHN2c3onJw
4vIjC1TlEd2OIHwp/mRvPY0uqCyidEC7ICO2cCCh0YXaDqxg/Mvfy8/iwWjfT/gW
4EaYNGVmLT1Z4y/QqXsyHo2yVkeWbXQaeOyzVnCTQlCXZU4I3pKHJMHkxDu62hT4
RRmSWkT1xBliB1fD1GJ7Vv6igpnMHFb48ZFEr4JMhuEUvcxhYqxVHkzBHusXC5bf
j/JELs6ZlWTnODCNU5BBwFEumGWD7xm5fXhO864LRuA5VVwMmPAEaiQekAIB7sDm
DYwuGoF1q+Gc0EjBJeavFnjMacwCmZzE89b3Z8OQJ5ZYE3wqtVFZyew2hbfs03Sq
imPiC8AMfCWdrSC4RXbHLcILT6Ylh0c0sgh8WuFINNQmjCiwBGgXIAdImsS+us24
i4J8grTXmkoXBezwzlu63++4LyTixs6M1Oj+uLfXJ6YOU0TTHgBTN2G0DZsGVgtP
wqj37dohyVIzbFWOaggxuPdgvXWUOVuLrnxE57C1RZ0xMr7K55pAOowrhJZAyjct
MejgiuFu8QfsOzz4Wir98X9hbvDRpzg2ZhoFbjgii2qzfK4crs6yuNvuEngdrate
Uc7o4bUAmjnFNf/fLopMUstrqE/cArODwf+hQrBjxNKU6poKGcMA/KWbfZppehFM
89JR8RShukwRXsX/SO1RwBwKiwKU2eExTwkmbVbfNiEkgFQoWN5fikeZfxyS6doI
GVHDgWcSa1SwlJ9KBLwoIwwUQM33tiDCJT8cbTCOOPfwG9iDjw9+HwwHzZeD9ED7
6Ufo9o40bzS/HKsVsoBIbWmHaTdsDn4p+eMLA6q30s2P4XGPZDx+UdQ/3RCHD5Pw
C8tF41TsjtDZu4mOr4DBe2juJeKowq9LEKlDk4zluOh3Q/K+EHHRZFfgsEJ2Drxv
stNXLnmW4iLl4cL2T9LKJbR7fZYYujtfpUpVy/KMWyzMiE1qCQfgN7HVxEQubIbF
o415E1IumUnVIlLqmK04Lf9UMlV7WGkEJ6wJYcmzbi/9XF+9SGPrHwVW2JkrH6p4
Y6+SCxOZoIccAItAmM/B4RHhbNK8YAtbq2XlNq4l/1QtcdCkOi3Dp4TDwUc87JIQ
Ufdi1VMare7A7qGQ7Y4N0N45CNKNyNIgjwJkboqU/UYlXjDHTGq4mBDco8Y3LK0D
DapXX8LBE6f5FuaLb7uPhoF9hNPgEMhx6gZLD0yLXYqF0MqCkPY4qt4TWQNRdRSh
9kgog3f83dQLTtKTJ85L2kYqwp1YXJ5zXA50S70lvFs9cJHCK+6umLFRV5OhChfw
YW+PFusVoJgNw/gqZwz49ZSPwo92G7CCejBFdbimvo7YfdJi6CILJEiPv0i4I87H
4fM0tzuk8eXFuTCd+34rJGMQZAkLs9hxeu+kP0Os5wtFFs+md8M6B+8AL2HlONwJ
LYmHwef1VPuyUiBdeSZYK8JCcJl4QhaW02zJyO0Hzmbej+Kx1pPMiuHU/MfhT6fP
okPsQLKZdNijXwMQ+e1Z/98hhnolLjBUVSxaZDNRqrBir4hJiIkBY8zUB+4u2Zab
qOtqqx8FC1HeEgrEFdaT1SpJ3f8Sc5Cpl9xrl9pf1nQZ54WDKIBIM+Rnz7eRDF1S
1/MPypx4Eao2IpMwUQJDPI0KH26/NqKzv/W8Bi1qzWWQGC354vyItm78+B+kIzm4
iNfwj7fObthuBZpkhKvLxC6BI1/cwYX2u6upYLgfv4bZzCqXd+pg+Zx8v5aSoEPY
bf196x7KfPAbPvrCNbxcYqGCfHKHmoG3gmYcIvfSz+N8kmeCMJn0s9IeyOwIBSde
h1obfUrYoSsXq3EQM2bFH0HgZxrFgYvS0PCErcdGn+81M/L50MYPM9tr+anjy5Tf
OubK8GuZohjHBGxo3EopaYnY3VOGzIVIwqr1AQu0Ymlk0Zd7ROHimMrSPgiL0TuU
kw3uwTr68KzaeiGuIUn8SN27JsCcv1nJNU71GB257X9/Co+xqZyowpJqLZjwAQyQ
Zt5g7KS/ktk/WTt1ZmdKWwxge62eZjdRfwBGg/fma7s=
`protect END_PROTECTED
