`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/TenaHEEtaV3IXeVSi/u8Y1lnf8hUvSjLorJ0cBLs1dfcnKxRx669MwY1be60iaQ
wjexrcSct0Py4q/7ncuLkhnrCvzQG2LMFOq6DDOSnqE9FHv6exEh6lbOXWugKvLD
RCF2d2Y+x+52XiiVrZfO1jrxW3e4o/PASMid6US9nvmlQF6NQPJND5U41TP9Ufjj
sF1ZqYlpZwxg9Jrf5IhIJZ0iaL2NFBiWp3km83nsWL3VOhDfcjef5tG5ahqzQmMe
pDCoZTKavH6KeAJeNZNjf5rAvyj37I2erYVnZih8Tsk1nP61eJSHES3eB3qpC36g
Skq3JWAFEWemOhcFs7d/yWcIf2LDJUgkcisXK8YOCd7yIHSJmIrK3GnIZC4EAq09
dkMTgMbcNgite9ngk8z17GpXFg89iV9KEJ3dtoSyPGGFNCXP0ZeL9Vwiuw9txU60
u+oyI+HhSYU8MGCgEgUeGEpDFTibzlPUprr/iACL6xR4g12KvWGEAeD/qkrbfj7g
Z0w2i+3E8DQYRe//I79srCaGtBYI/iUH+m845QJlP8TPMJv4ilTynBBWzkbRocFc
qyqLqg1QxMxGGLqyWYHfmEurqYGFgf3NdEKjnDt2CPCYFd82ohHGy9TtLSqQD1kP
IX/ZHJUkj5a6biIWAKVcvdDQm2gH1OMS+jCm3ubUr7XYdOWOZkFg98u8fbcVU/qI
1eONxiDLqnKTcxm8u6+kThQf5FYEF8yujwQLzH/91VwEZC4ZSLps5DPwsyN5hscL
Pvjo2cs18rJ5s1z3bCEPVuhEWjdZwvdVz+bRVq87Foc0eX7TYEBO5rQxhII/Q42H
OaGsxpQWjywk/xFhM/w6i+GkCysdCgI5oYV7/781OKP9w0v/J6+bQY/FgddHERFX
3BWmhgTYTThe8qeE5EIzQ7Fje3Fu8mO6U7wc99fNrK0L2L40Wme5qINctYxIJgDz
620wYier2Qjyz981EeKJECS13AK8SgCRxkk6EVi6ZqcRLK7VO0T94F8Y0Ok8b53g
DbEI3tm39M5eAP3COfRAgYU78e8y6aKnYEjRuw5oZ7LI5KbTPUTQWU3i5baIJ9zh
sqWp8Hu/u643wpIcwShOQvClaQ5uqGQjUS6yHtwZQ4AQiXD6rS0Kewg9y03DsU1y
q5mjlbbgjx7fDGARw5kS38WF9C4pJqt73bUdmOynkcJ7+Dqe59hQDaRzN19bfsJX
GCUFTBDuhtiLyYjQMNUwmYq66/G8VL8dsfoDDUFI6NCZ4FTijMJ4ll5S5aK+4RTY
74KUhOcD+ErNPfcL+Z6yl2pn1xzQlUZ+fZUdAhUV+mAC5yM3Djovo/1GPpNb6f24
MLTuSGvlaCe/SQzxTUz8QZ5PCHh03FXZfwAdnhjQHXoGIe0qHG5ypyvoGZN1E3xl
9TRa2jhYS46wwH0wAhKfTB0ZEYdBCCFPCivAf01fGsP/2/mCCrVTXxt16NyBp1Fi
++txAkAjdS5Xe8ZUUraOFyHm2x6HR8+UOKRXH7OGa4KnI+a/wNg/F3zP6e3mBLBg
fK0lZklH434wTSEhofkz34YfthA005LmkP/uaMgeMNIwcBEBuacdA88bwuy7418/
bzbwGl2ichYqDRWRfspR1elouLx/oAG8fd6kVd85OoBmldSkvimJaWTxax/WOZYU
pR734VUseRMiin1C700zxRIlEwDv4WG2pBTKcggzxgvucCAdeJQuOtHo7XkkdFkQ
xAr3e8FNgc41FasWcQXIItUN+pftfp/dG+w94GgkuekykOnH3w2sHK9CTUpu9bM0
jvxYX2W5NYSV6wvqGBmhINMABxEh3wkFSvRN+LcwT1M3klvubu1dsENPQZCJS+Wr
b4NrGHPY2rDus3lH0UYygXXwLtzgCWv9TyxTLUswNIXqeFCyOwnq30BHWf0qBZvS
sJkCziKBN1mt7TjFnT/9UiL41okvZjaIpuvrl35YMWUcKMgm+TnaroZeEO7JLmv4
wzfMjh1dxzKh1l9ZO8cprq9JDUtF+si710exzQ7AH+8/eRvHBtR6wpL4tXhPahho
WFZkDWD3DBlfld7V7fd0WtukKKKGX5ayaF4P8pbKTx/AuwXEHZra9735hlEdieuD
tRrzKBZEv7KdSnBhYUXVf3t42LrjdFayguX8PF4DRzL9hcyhL4/fKvIKCd0otlzr
fDxlvmJtHLY5xCwVnzFdDDjNm0jxSbggUO6c1Jahz8oPC+B1/+DXrZISW3viSO5Y
TIf2ydEtZO38f44UB08N+18HYScZwQzIjMLbzDiC9l3qzlF7i0okECbSKMUatrM2
kqZc6koB85iQsAwPNywIOM4dUKcoJoqEVybpjS7TUdki3cu6geFvmj5q8c7kJ8Bh
NhX0VvswaVjwI84jAQ9B7kW12+r7Y8RyggTpo9YzMTT13+3ZX9PIsE/ZI5LUnpMZ
aRRcDOcd8vYXao2I81TgDq8/vs8EW4LhTTo8ssA1oSq71bVpKHm4LW4j0HPZ2Zm4
R1ixC7EO850Fu+kkNF45809zfaMO0usq5QBsVxtiY3eGIMDJOP2GHGRDoZRUsizg
albsKdqFzyxft8SkZ9n4rDyTtIbBmF6/L/zeF+HTM9Q/5frwy5I8QSb0WNsyeeBI
2MNK5n2rpscqfh2Nd4YCX2f2ZSeHEnLTHb5vtCQTQcePUpBPIycyt9gjLUuP4TPy
V0c+BYonxZqZ9CalpgRyU6nyeVSwfmCAR1rbmInnjG5duUsgz76PeTQOLoGklLnU
B4zWngeCS0zvTXbt7AidA9laHF4d79puuyOcBRFcyW4zmEQpKD1E9PHwyNNWlipb
dkOe81OoOTm4Bobej3XO/zebA+WYiZ9eUgJ81lB/vDNxToN7Fy6hd+hntra/gu9L
jqdI1acNGlihFzfSY2V/GLL/1q7balI45ULeJbYav5HRS37/LW8FwqCg+gOnGOOc
acXwCw8f4SMLY2h/ue41XQVKZwH+XNKNRUlSrAlceBsG7F43qL4amQdDW29m5IBM
AIQnhHyYE5Wznp5xsatYxw2NYbHRPg9qEfByxPCsmzvMlhfjbZoLCWQ0vXUv/stx
H1qSh5v+8pnl8sWsWUfCKfvc0sYWt2vMInIqFGnFovh+FB2kS4jCMXcAye1oVphE
pIvO2e4gMMpNmwtmAtRsF0mRz5wiAFxkwHe69yJ7oSsKv6Q55QJY2XpTX7mJ45hP
nVKjBLM1++ekBj6US5y/ueKXcVNUFShbMw29NOs9fkV8P0T8+Zx1nN3ygSSATQBG
jyGW2NmfPdeswu3Tbn//eFo8T7kU83lHMHFU5ocCMKbLFXGT9UaNuGL7kvraGEHC
Y/yuJg6Dp+fMxnvUwymijJwQmGyvPkE5ZYiumxp0aEwAtPWA5blsIVaS7fYmUL7c
UEo6h5JeO7VEX/Tz9vEcz0iV02SPb4dAfp9cqzNRz2tavvpuSqmVSUXsMQEjJe6e
xPcp6M0fRfBgxJWRuaavw7Erpe+MaDR4PBbvlws5VW4lutJ9VymGJOU3hUkW03vl
btVQ3/+V5QsOAx6K3ux3Y5WiVMC8mmE6j1a+ktG1TiKksZrnILhZkyddVD0mmQ+b
AJOyLmdaG1qfJL/X/95gzUVko6TbZXiCFTH+KvpbXJpAk01piqBaI4wsS1bWsDJ+
S1gKW7hNfW4j/Rhk/n77y6MoBkmANgjcD1IDqFvB7ZyczBrGoFX8WZUzqaoUcuRT
bqZArmMZDa1yKFYn7ETjMepIeuptC1lNXDRjRIF7biMr7uKYOO7il3R9IGEClt2J
bdRhkP3myb8TQKfPU3W0R6zv6565RjCNgDfJHxxUecmiHwelypNNPnR7tygIZl6r
zV7R+slZCrhc0ij95VsxFn7TEv6uH4XM5UHdXNLCxaqmb7H+XXyn3VtHa8nTdcFk
TtInm6SBZsf32BGAzKIDOjWkIIGNVPCe43MQaHfcuJpE0NAVk0DWX7xTloUl1tKC
+T5vNEaMbv77vY4pBa7iqbkc+kA13TjcnoZKprscoLhX355/SKED0B9bhk+hhZnO
jlkJMWG/SVU72G/pNqAMIwZJsxzScyL5thc1/OWYOCNXlXNEPYdIUHS7cBsfTady
UMOBnd+Ccl9VecmxR0ud285dlQardphPpRgwGWTZDrtE+mquumAk8onxwl5LbbJD
kDbME/poUjRfv9J4JeFfLd2F8A8YOdp9AHYtVwRTX/AJ0LYJBl12z2Eg/JgKOAGC
DiLtv3BAJ201UUd4Q2S8R+QIA6bQMPXqRasuNyq176Ew7EoqDnW1PhEDh0GuD1ZO
hlRRHA7Dm/pwrztq5JLtgAaNU4Acf48mfl3h79fjqmcEiEyUlcPlo6Fg5b2HaTsA
Yp2DqcSn4pMt/GIP0FQjlXnYDJhOE/u6lVP7f7nOs9DL/yVdTuTcmYYYJL3+fSFd
wjBfdU5RSyC3UVyvO48hznubTwWmnB1ld9NY2qjNkWT7k8feuWE0KBcLwEmlOua4
nLLlLryQ1QKA/lvruHAdwcbtg+sZsIQr1+ZrJKGasE8mga7/X7EMz0OEgZm/A7mD
B7jZ+aLcr93J2ZkBrQjPHFr49cTM6IK1RZzSd7ZOlgS8ATaZD2crZGl0kWQrMate
WruBSbJ97MYaTKKA13N7fXKcDkqkxhr19G/TPl83pQpXxWQtV3ve6nJAr4GeGZsN
BzYJQHos+GTEQlEdmJlzcCu+mBMHjXMoFPAaE/ILUDresd7rax+1rJ9ytgVTrtHT
uX/kXQ+tQKOmbjcI2di8jikrE/ohVBwBzUBrPxa0a87FS6Tb3A3elbB0J/cZQ1ZR
nilQjp4c69WqbXfnn2KTYkGJJZeuI4Sld8zeI9DXwLMqU2xm4cgmg3C/l34UXuwd
Kp/wbu4MdP/+HDlVGKOpDi4D9Ljt4iQCqt+FiucVfJh6ESV/JxDHe6FOy/ah4Puw
IZs+ZnVzY8BQDmFfjOUtzBio+Sa3BiyiEPy/P+VF/HYCyDXNpEYU/Zeh+3/yCQII
5wbSUpFEwBbYhjaoAixWE/qe5pKbUJbo+LZGNKZgaHJXI9v3Ci/42wawZyD3DmJn
J6Ti4wtrIq2AGkdkheRqyCl28OmoHt4XXtf6sjFSfxt4iIJQ3skmxNe+imSFV0nz
iQnVVxT4Xi1dFXJQgb8LI3a8QP8ARkuSpPp1OPu4EcKqZWuqStCVDKPKBIZAG/Yy
WoJipj3g0r7xGl9rQ3rgAW4Gh1+jrVjRb02o6fPKoGY/fLczMmtk6zCdve1/KlIn
edt31XxSIx122JVkQqYAA2PwzE+jduEFvXiravdFNOnAucnBRLvvioAo5SVQoS2d
IF8zF+jgcFzV+aX7JGCph2+zFJSdg7jVy8Ugmt1j0OAYQggUhrPuNcfr8fmLrqHP
8FssL/IIERtQJZ2MO6O6SVe+imNugKeewnXxVzgzcyjzmI8qAAco//4nMcVXp0U8
Ez4lHbP9EOLBSaq5Ud9OgfoP8ryQtwlPzKth7Em9RCer7ReQmGUX2/EucrAbUSYT
NgQhp71EltXdGqy6RJpOwgnDurKvs2PokMzBXgHHBXNG9SxdLhUZpUhZ8P0lkrNr
kX+yak0PUBJtaAWU13ak/S0a47/sszMaU4YY7vg4d0C7GmvkfU2+ONofJkITTdRD
Lfw3/W90i/SawUtwYuFcDJgdau4Dn5qb2rUsMsu8dGR8IwgixNwEtnQwDsJsm/Ni
kHIeZbYYYIjxqNsa3OTFLYBBz4/9qsHTwy0A/VDFWDi575YHEKkal5p1IMY0SThw
xU0PSqXTzgk8mQ/KHxzfxOHyxt1EVoSV5+lknaQgwap2bMMIVIpI8ay4xrUNwwbw
6lgY5jTY/CysDwKaOqM9WgMAtlDylkVJzM7NzTz/hJpSk84dKmXmJQs2G96htkm5
B71c10p4XCpHiNbF/xgITTDXB5RLx2LV3GRaJnzcooY42b+zUPD7GLs/61i7LZu6
1VHtbEyngnVBXChAdIrHi4y9pxUh4+VoKYmjg7KgkfMxP/bvhPnCUYADrQCgOSlX
cR8d1FUK1BeaZBvu9qI0qBpFl/F40ofUw7JeWj/oixkv5NFZSk1zG9IIbDtyyHOQ
IX0ogBBaQogTLGh/cpwr+mwFTzS0BBvwAt5QG5zpmzCbRf33ju+0GXBMWIxjR00z
bmVBSSO9OUkSckTjkvQDMdTwWeERCSRa+JRnoDx+RuUOa/1CkfZl3baULrXoWBce
LHxCkwXF0R+r26lrURG1pmOyGihSpHYfmc/Ok+UKdfrQbburc7wNRBzX5G/zIaAA
QUmucl3f6dbUAwyEvE6EZjOH8J+ize5ONeJrlHe1X4FckAzU4wVUG43uSvqxgSPu
T3eTjxJhLyixHQtJndngBAysT3ifc+dv8A0eYh38VJIMLPSZRy4N/bRFo2eKbtom
rjxjybLMBYJ9PGqrV4Xtzw/G36jF8P5hw3ecszub51s9TpmXq+tBw70YmoZraoAv
PCEd015R0nAdwzprmc0kCsrOiEQIxft8rQPoYkYP93uH3GgGT3V6cxeMJz9+cz/1
s/9E9s8beQ+Rfnctvmvmu5uZzWZykM568PMjO82BNPmZxD0nbv5PFCj2G6t1ujvD
oLDNBKVGhoAcomQbGYB3sKZTyZOTQwjRh2tiypQa1yIJGYmttp9fXMAslgZWGrFX
b5LAdF2uGaN4LUZTD0tB/uCr4k0IGu/KRx8KCe+geCRMSvK95zjjV3c6nM9ETpp3
px/h3a1N8844NSrIdmqbKUhdYJa8DNVA4cX4UNTTxFd4RdsFTuaCyvOb04Yc02KJ
H2aUw0em2YCwwYdFFhh/YffiUFgwoy5iRtXKo5yZb+e/oxEv2P20cWJMAqDiv4sx
6gLL3Ny05P5NiBSO3slO7gJ+44FYwkXN8x6+x8Kl3nQjeUIHrHzxI1VxiZz6Q2Lm
ym5e8ylXkB8Ya6DeAZzlLteV5ujOcGQJqf82n3UjftgRgv4exp+28wvo7nLW65P8
VzgztfIYllM7vSlQKsuAGXvmiUpOdVAIMCWHbJgPe2G5SWWjGgc4jYHFamVs+EaD
oHq6vjRi647QI9vW3C4XoDPa4FIUZKhKvwZ+sS2TS7EWQ1fkCJkAi7Ak6Om/g968
xaZr/PxbhaXkhDHlD+jyMRhUHGCZ18nFPoiQa9mc49p71YULuYUESqvDujEREypq
yEeQixw7y0UmPCm049P7DIDWqh6OcXEf11zCeb4vaGbfLaLY0dsWuyFYcLpifJje
SOmotFW+Y/VKgbw6Jz8idHHP2v2ZN4A3e/IGp6TI/LoanscdlEH8rCE/4NH3cO37
rmjkqTTnMvkgxuojs+6k1PIBvATMdEKAHhG40S/U1vgDovwpIr1e18UctRS99ZcM
mOu1Bp0lYK1eYGgYibzW8hkCxBLF2rSzc9e4S5ewdkxlRvSJUaei8OcdBAGn2Uy/
C90m3zO6bftvpJYaUA4pgO9EH4Msb8p2npa9TBqf2xKjX/znW5pzrOA4c+LjQq7x
EK4hfSI3H7Eb3oSMJXIgeMZEaQtywS60RlylhtnDS1ojXf2tt7rPio4rBkjkVTs7
fkUN08GBQjuvRYTJ5R60/EwVZhCnSkW59Elk04AvztFKxZBorSuVgWcKF477ZlDd
uCnvWPCcgE+y0oA84A5YoWl3BYwqHre9S2ep1aIs3WeVPHWyoSvmJTyHTsIi50q2
l6tIG4p0ocbwibqrXrTuE8MJJsPYy9KsmMuOejlIi3IE4LCWSi0PJvPLHzo49cMo
qauqLRN20uOMoWJ6wZXSPzc3CDzBQPDPU18f8/dO+dNsCfOjj6oNL0ormfLmBrBk
/fjDNkRQFuJtxrdaiYY2gdfmspIQ4S38r+oP29UxSP3KWqBuIsU7RWzSYvJ8CFo+
C8eRTFKNv8T+0B7FrFoZaORTE3Zef+V9RVnXzS1iLlLApRtAYYr9leB0DQXEOF2Y
b/iwbUy2IC/tw9o1I9e+D16jX0RMLoXp/ZQENKEx3Z7uGCGrwWms/WNLAnGBRS3k
bCGdsYLJO3s6q8Aj8z01Ir7T/+p0YGBfE0fhvbc4j+ouMsVVlB//oVIOPKEdsdaE
R93zR62EB3B9d0o75587deut5cdgcZIpnb3mJ+xKppe/caufDmhwBPgOQKhBTj+P
PoRnob4B3rJK4hbzfO1FJi9jnjy/FH2Af/vBD8JqwiWUvBqvqwAdqI3XKY1ZdvEG
P7T58ry3Z/SqukHy8r8WtUBiCZI84jm+Btte/+qwfWrBfUDH10L23l2b4RW2gV9M
wo4MGPDM87B7rS08NUUrAobGe9XCbVdlTVHOXy/p/QskfakewkKu7f2KXPTaKF4p
baWEDGlDDKa+fvDLXV6WWExfI3Ogt7sN5XUQaVgKWw+xpnL/4hjGq3AM7m3LqElK
z+Vq1gtS2IycFQj/Yx/AaWwEfk5bliaKjMHIj4+gpr/7WCrto51UACq5o1TadgHA
wj/VHAppSCVZ+lDWJIX4t1i73WZ3VOHLsL245zhdK7lTJzy8izby6iooWo9CJV4b
Rs2lAeqTOPCTtMqKzZBiMTRlC9r6mhR1j/dUKRUSJzO3acK2Xv6E3+fG49aWIVSS
/q2A57TRcxc6U0eMGw7EMUAD+3fXdImbTX3gClzYaWxM1ChUZapdsKXE1o6HHsTR
dAY6ff2gfuLRlpm0BU3wpot/6hP3oWvWQ8j94j5ATkrBSr36XQ71YxTzfWRexdW/
RDVVgJLCOndvyGf6rleHaue0zRnTAKKlasPIUWShyux++7rPmUP6dR82w/qoGmct
lT0X4SkdZXQfC8MAtO6Ey7gZDUzl6Tux8PemHqzIVThaDpcvCdU5mvCYjQc7EJ32
Rwrct/M8/FattIIq+h8b0smPK2PxZCCnuc9U9yVpKYPpxprUGVC4J3nB3Jl4aXNk
2doQIUd7XLZtNgQ86/WAMlN5kZmss7MBAN8Q6DRapFqkChUwTal0aAp7GAjE6f+Y
MGeJeBPTKVpqo5BUvs2xDNn3Mozp0Me+CIxra4W3SQLu2qWvAEZI02tdadjx1ZUA
h1mqsWzrOIFp6sOrloE8odOEYS2+FPhL0Xb/qyacY86RLRILgTW6mIzHXFB8SHae
GEt/wDoRqKPM35yqXjywvEmuvRg39OujzGSJ54EF7QUhLDk5CJAWAia4P9l5Dqec
Et0yvMVdBxnSt+/jZQaQksN8fOTF3RBnFk7/+s7h3KzWSBBhQa05kNEWW2aU+qcQ
sijtlx0TLa8hlApjab/X3bhev7e6HARE9IgGtYG1X7BXJUINO5BmWTBD1vP2nufU
jpme7B4UhXEbNAXW2p+AaORkOJRyXoB1wKLVhS9JC/R6Ug2Flyphyd750ksyhCDd
m4w0E5qvsxiPlUrIiA7rR4cKyBV1u69yb99HJpVmYJTfWb74zGwfbpkcrbXWFz42
TawRvOVFVMsUhx4qluEyfHFD3Is1dYKE07XYqeCcsEl6PmAKow9qZqxkY3nhqrdM
qu1RRJFODwxNrRAqgJhKIYc3zMhC9sKChxVT58zxTMIlcah4z2TE1/759+zusTS+
jKxB+29q3SwT82PobcuzzEAj1A7Ti8RKg8+8MLP5hKxbySd0Adf4HV0eXwHUFMXp
REotUKB6hGWsj10aRo17cGaSnzf8YCsx/PPbg52ITpUi3iQ7CMRt/TrcG00qNoAv
xeoJkxjwYR1S1lQ+8a+k4UQj6qVe+8tz3jpV6r1/opUYCIGRrEgmKZzQ+BuTzbZZ
QrlIr3suwPokNRcKE/89/Ie3VqBIvFGxVkWK9MqONa8KU10QlBpFp2V3BPwu2c7K
e+fVBNKCZ/tkOZcGX9qCEsYwku7GglVUlSWNuB6rGw290qmEyoJPEnFD9h073AwO
re1s2Dk9ZF4ezFkcMSl6xMMiZFoJFFHfUWiQj8NZbN1NsiCBPfJqV8l1mwimA7x3
cKc3u8JJD6dMnBg0tXfG6A/M9evVAB8vaGLAEo2Wu1gyf5fA3zB8f/MS3W3+p9GB
A0IXrnnP6hn8oG+de4BrM3FnSt9EJqyK3+e+SDPYXS02posKwu+pdlJypfZBbJq7
PaZZGxdjxfYy8aqjpB/usnyaEaRRxNkLi6bFYaNNlqFMZBnuccYqwoJm9UFuOBJn
jKtgzaiB3ZDf3yEvpwALgGqIHk0/7dRTgOya34gRZJamRtVWC5w5wFaci7Wi2QGF
lYhnZtdPBAoPCcXD0NhTWwqSRmzBTjFHyIOsEYsP19Dn7Wrp+YLogaKjeMcbzmmp
lJpMhBYRVzeq7HWx0DJUXHoRVukUDshJWwi6pSWVklM7csC/2P0SedqdJNY/jqWW
u6iBAJJdXYhdclqHb51RN8Tw+6PcShMPc8lzqqKes9IK3/35bxfh8cdIVojeQGZQ
AHVQKih1I45ksBY7yq763jMck/hTo4GfLS5JM/otzxWqTHZjWicSnm8BbL+n6OVY
VHaQT4SxN3t0a1FmykvGlDsnsT2nMD9afcibWeJXrBaQHG120+GPmvYDGr9igET9
SAJxOaMFjOHkDb+Uq7s09TFxzCyaty8+D1374MzW13gLBzrcBC0CfV3cNbvWpxOU
lx8j0vNDZz+rrW7+NtCIGNEPdQzR63IJ2VCemaIDdfgxqzdWTQ87SemtUfCTyMUQ
wn8jB5x2KsDXBriSalXDUdgfYcEta9kj/6DHuuO0Nefc8wvqZ4g1y8YjZaJh4fcf
syeKJZcMdF+dzGfkZWoUczOUPCoXm5+0iMZVtHt+ZAH4jVpcakXg+fln3a6i67W6
e3ktbjDoNIFr2PyPyzuhK3oDtz+giuaFHTskii8LfGr25nL0GbND/+71eXAPzNew
wm934ZOU57u2JO/m88bMHV/kAqciMcsbBbZWqcon2KFG+lzD8LGmoF1B+ffXGraW
Tp8AzerZ3DLqb0L7VuC6vD1bQGqaWewImQjHCNruTO+cTo2UCSkhBq97C3WzlOT7
P3GBYwAzT/wgDuffXc5oIElMhWkqaLlByMpqPHodz+IQdWkrsoXYyqAH4VxdIus5
eOl2dhviI0KPtR31/SyhSlKMDj1O2Bq72v5A+zdvhRLaLMeFAg6pH/GTQjezxyux
Bqv8bmcdrEWWEqSCttQVvH2BPk+F1ashMYSGG087tZcmljJEgWCMu1Qh8p+RqUp6
HkRbpQr2rLHYx0PcpKtwwTzaAVHs9A/jvu+Uo58r1l8TMV11Mr1fenJVjH/EETjV
bcNuDWeMUGN//ggyI+Ktq5lzmkyc5exA5A8jIi1wJKwUzCDDZpdYMC52X0GH76m/
DO7I4WYj31mP9mmNWszrjkMEPUzJ4eJJmRupVnEYgICdP2vhuYO//lgGSNUqQ5iz
FWhC219xaXslTWorEIXFRjVqz3SrVvhBkXWDxKABY07fkLcnJsuJ4cxPCwZ8vlPr
DROZYYgNAW7UVs/YZdRNAm7yIyCqwHsOW7CkCes3ca35KOW4O/nkzVCXdKhmyaaj
yMQOGzIcoQhguD4S8EnYqB70XRBvbZFuiwtcyqonea+ldPxvGNA+Gi6TzBuhyifj
5SB+TWDAMWf4GX/t6hPvEJ1QvNClPKnhVe83Jx7WUhkGvE2ZPYwlsHkAVjYeDTh5
hNbhIFoc9QmlB+4PArG6L89blEfAtsg/Mnupx3GgCRfWXPpaPSS8JVbWtmuCa7xo
X/4xM2DsetVAXafvq3GV0o+l/981Pgb8fCRiKlQPh5DGcZtAK+poru/Kx7T5GL5E
vRq/QauJsXT9k4KQqECBl1kMOI/taJjNHb6l5S3JSro7yGq0MNWWnNLzhPxRRQMb
KE5+1oPObL+/dsfihS+qBpl72iq3hcyNOcCaDD6FLU5bUb33zdpG2PWfrE3Mezzd
hfJqNC08oGLl4b8FlhToXx5BBrKBdw2aoD0ALE2TEg9BVPCuwdzIaFDnhmZOl7AW
8tDJfrl3ZKf7FTis3cALtSKo2YM+cqSxuwKfyncWyad2uPAJzBXh+6POTfalQlRv
TjQmYlcw+lqs6698Oweso24qU6NnLhocZowSYO2FYrY2QT8NNptNNP7hEsxmrkJT
ziCRLDM6S+RRvvCBrP7ObHBKKc5XDYmfu90O+KijBN7i9Z8wz53fEbPRGHlLaJDg
bsg41ezVJWxPm/Z9jvlemaxrtWCRgBi+PzsyuJWbXki0trMp+Ykl9av1Fqnkg8zg
EfmyEfCHyozGJaQ1JZZMcMXtj4HV1HLJ0+HsH0rdPshHuDKibky7Jt1owCeGiUZi
mnU73qQImdDXwy6jZgt/0rSEML0D9yT17W3+SxQEyxEPjvr7A9LjxHa5cngxYTWz
tHk6bkytyubKQy7ml3tHLCtevxtHxkm0blNsLjmJah1ibRTQnRn0oEpeOX7cnfAx
GO0RrZ69N+f0OU6Lq2sEY8c6unZ1lhlpkg4qw0lE9lLPnI+uq2t3cl7jKoe7H49A
IxAKLXD8XGGk++WhKhFALoL+k1gPc5cEZ03k3HuTCf5EMCUoXuP+mXq9OiWEFaq6
vmUFLNGXMaKwlZxFG7G65veAAVfIOsSVReDilL6cgCI6unSBhem8IDPmjtRR5/rh
RazTGbRvnobSplQkupsl8jyTeYQKaVGPBz2eTVUmC+Kei13LEy6Fvas9FXDlsJMg
eUzdm/1jrqwjsbQ1QLQN5uwv0EoIdSopJdvDEnu7/x7efAVxgzj0FC2q69WpeGLB
2orNLcvys9E+FbxUQEl4+rADmbxPJvEjKKM8bstSThg9L+uP1NtCqJqUh03pek0f
W6JampIQynDFEPz35GxL6xERJeRXNuo3K5VZioePiE2d6vW/kwuS74Gb1NSUQcoj
mJKQ53zUnwV77oKfZWZZOgBN8tmijOaC3Q+CVM/rurvHXriYz42ORuXQYF8uW0Ig
uklU/S00Nq7UYT6N2abLRcqN7p6rEEO5ceXhQ73Z519EpO2BlAOQE4MvtH6gqfQO
DwmFmiVSBu4UEc8Z0ynY+fOszY9ujOjln+MiHpPnETiBd8wZBteoE2O1CCkvwRMw
aMpw1JranYWBTRA8dfc/XrQuBNzzV9rWInJeviLlq+Rfo5fXnj1KXGP29CFR1Gf0
LEB5p7o2ISMuj+yfU+LvlpFI+nt2TLQUAEH89bRHA4DCQnZhZI11GBuftbEpfIyO
OKOMX5n3V3SYLSVIg2dXL9wGaSFaJ1bfgDyKCCgW17Rbj8g949JE1uPhUU7Z5AIn
2ee3wjidfQSQrvIx7ovtuqx4pfE8nZW2WPxVTLZRQqzyWXvGTqxew2afP3Zho4MF
jOlDIIpS7JwLl/2Kl9T58JpwSzaYa+FKFz2kRXmXJwPhB0osoBnlN0en5LZBIWJA
JyxqAxTFvnG23RdKwf0h13iF8Kl8C9UdQRMMk5zi88Mj4tVEkIGG6o/YYbW5koXK
pjJW/R3NWzBP/oKjJ/XcY57SoBgsdFbYxa9oaBi2H99/OTRIW+t0AxG0q3MZ1zz5
Jw+shQKf2oJ9g9mBdEX7h0/IzoAMGXO4ktD6f1XejyGYgjQ8DUJnFOY7RMevOfho
x6l7E0Sj15A7/v9QTzbQmT8YmTzpy6mObMefPhneH4A/EPcwmSgFtIJ3UxqkDkgM
K7TkCuoZZJNcXgDXMxENGYO976LzOFl9vakR5jvxKbxp+cr2gQNOnNtViWLv/Fwi
lPnY2iYCAK7twceJc0kqpJC9n+r1H28iAbWeE5d7IeztGoVWMOZ+LcvTfe5t75bj
SeT2lq040SFCrVdEszqKPZ5bbP27bY//Kh57I3ddTbXdwdvC201kV7Tt7mrjGpFI
hxS8HYc7coNx6BwTBMg8v0M3iA8EwtEk3lPI2IG91Zi4YhVaetxbJJuIRKj0CMdU
Yx7eqIPYuHZo/QT5GxoUr2GwR70glOyyBsyz9ZRgr8FEKkIbI6EcgJGa6uHb+C7B
4Dj8KefL5Hr4eij1dwtWxxvAH/k6HYKx8807enFX2fJDrOiVATdkSVUOAuCPIYvs
f1Z1Z88YRUqxvhQJ2XJhvwDFUEfsGuVMndm0Mz0Z7hr+ihNtsjtSvCLFhBPNGYyP
G7YYQcV7FsIjAgrHqFlTN6p+eqnC/3RK0rcihVPLpoQ0RTe+IgomruxMUPHSZTUv
/R/Wr8SGBl8D6+SD8VRsT9ODRvpnO2cQLNaDWpsp8a7AFYTvTpfo5U/G79vKNAr0
gPVZlUTnMi6GhNKYhupjD25At/YJ9KcDuc80BVjNHin+h8nu/G1qze2mEuVPPx0t
qkAWlNQo32IfC4D4oIGMaQpiJUlztWVTK6QC15tHHPcnqQ7nX7QTLWx9NZpbp63Y
3xSXw3sDcaxoPPlox1EPvS4ANa+4jrmzC9b99/4mhja/kZfqWEBoNu1JOGC+Ke13
RZVAtHKIWd41DmUNBdVrfUyoot4zxS+nNlgX/mUnL9LDJ6Ekiny85Ew2fAYzQ16Q
0XuMA/rWeEg50KJEvDjeC4pj11jSJD36TcBZf6iaIR29DUjcZqPgSy+42q6DJb8O
Pp4IfduhoeQDkuI4zq+B+St/KRsZoNCWas9I00fejevVRjANezp9qc96/Bm1f0kR
HPRV88iVT179FpQyreWDJj7RBf91tAscnhBnOuWuAC+7w5eoiYNAmvSEwQDnHfR6
4pn1Xx3p7KlhqhaHl+L3gEhevpx2k65B4OX5jks63/Dlqvax2kASGALjfsAueUwZ
5E2DiicMgO7JO09uBytYrxdqRJWor5hropIl3r1+IeCJ3qVzzZnTwUaFtmA7p8rM
ocljgw6oNgUqXYZ6i3VlTQvJZor2CLIEcEpblocNuIxG0eCB6jlwQzulCPUbxKDM
Fl5ggzo+COXDo696GwXiPNjhF2/fiUIwhZO91DYWYIHlFmcXyCsMtPy/QfRkmiuJ
VqInSrSGuXyFkiXLtEHokrWS3t/RnSBP6zJ1gvPN8fBtp2hwT9vO469X3O4jBEOy
ref2oWUoiV6GWeQ004hYsGeCtWYXZw+XV4+atFR9N8AX++F4sukzgumah237ZPsI
2pcUYlS5c7bhXqg69o4Y+Vr/F5giWqP++E28g/q4YPNUTtv6uaqUydLHSCiReuji
xBrhA6riaIIVsOdakYpPc8XFPT8AjsJYEgfcoL5FUteOVmTiSARm4+KgGgR7rDCU
Z9QosryN7KEo5CL4vRcjfyetJvggsAfGIG8+lk2YLAXlv495FFW/RXXEvBqtUxSm
bKum+Sn3oPZqKmzSVjKwLTvZ6YmVOXZMKGtcIoovvCla/fIdG5f8RyzusLwPZOMM
jOIWgXLWhBHa27Jegh4uFicIkcbcFx/Hzo7UwhmlRa8ghhK+/AAY6B+k5SFRqISf
vJ8jV43WDgf0GbF6emAEX2QrziowAkFchoqAwSRVNmg5LDxVx7OxTUSDJpFmTNko
4JhzRSKEeozr5bIDrnRPB/YiMqWRwsBZ0cVs2aDUd4E3OolKMx+M1I7XyWpcJTJS
RP2eqZ4RmUUGzwB/CFLi9AXW0B9M3Ewk9qR8HEDxGirF8X6H/b6mGM76nNg3a6X4
mQUN4F7dqKymqhxgTyg99IuVy17XvbWs1u+AVptROyLXNWIf2hrEvTaHFaOyhUFb
1peTvWNHbk51xevtM2PMfaiPfU0WrSGqdRttwJlCxNNsyr8kniKoKlx1KMmAxNJg
LZyKf7+QmCJL9V51Hruqd07Alc/42pXsHTBHRecNXnFYLtAplD9q6YnMeVMIDBPu
SKZI7/o/KH16w1syHdbCPVHiqX6V6w4+tvC5rhfRf2peKYNSx8tRYUrxrKZniRXr
hwTvGAgUlFXumJecOUkhYw1OgXVg3IqtDZTYzmCVVT0PQGKQJnoOER6FXf/BxPgy
+l2nST3FB7jubKQoJ6ER0j637dGhFgg5ywlTdHPXSFFi4KteVv9LyYfS4t44NZj5
eslLeB5jRBbQ6wCU69CIbpX7vSSyMECB6xLYOA8gCXJ3VEBx48eb3iL8QPtDiei7
0OS/mADRSZGwHMLrDLWGEPJ4shwgxCoFDZSyd3ZkWChqgksSsBBhXUE76g8IZ18T
5q37V4hO+J5unBNf8860pTI7nhTrbUoDlC+2yh7ZaAv0MXo3r1NgxZtHmoy2QS5u
LncSug02r/gCR+fwc0pjQNtf//T9muVxF0imILMG7LfIrEerIaZodB8iPWvBxkJg
IQS0gHTp1zcYDk+gk6I75s7Efk7rLWj46LDYtWQXFabS7VyIFgiISITa/Rx6Ldkf
2MmhU3v+vLW79IQq+uqG7QTfB3/FlsHnJZOVw6oTkfNBetsqGg3+jnn2RaCBrLX9
5IuvKG/eQArRdGakJjTpdoG6eAry6jCOx5DX5CyTH+a+Sn2HDTuQxq16fpcRe/Hd
HMFR1Y1ewPp8lqpWrzcZnuRic6EMhEKXAlk0lmpGWpwwK5SgGa53o8BJT4JlOzn+
DqrbTpINsmy+jdHnLCAL6ER1VuTsQ0li0rkfwWSamSt7Dr+luv35bs6aIMKRycVT
sK8D7815vzUljePG8MsRxYyFAnsguhB59IQGdgEjKwp0aiCad6q0mWvhdmkNtssQ
Ww4BsKcL/I9eQCsB2f/+NAx6ogsb8KuUAIZwBTp18Ieh0t7Nqw95BxY1LcqTl/6q
VOGEmj3SjDiCIzv4rwtKF4bLqMOhign9LJgiwAfZfem4N1+xWhJmQyd5XYhXAnqG
uItpnn/Ni8Rkz/T0HXkiZl3ar/vKq+gPetPHDKtDooQmBBNoVnjGFirYw6YoBYqG
/+Nfhs79tqrRLTiCH2I9FH2mM+Wsi6ZQ323eg3zia5bYzPcfx3X3g+eJBTm1ihn6
6QlPFf5nrMgAI+4NLwo/5heWRQNJlrMfptcs7bfMXPziHeBQ5unxXkMWEiSRjm6Z
zVJNkPRCrIwTaxa9lk4+HJpcL2mE8Pl9pJE1IyrJy7kOl95lC44OlkeOrEiNOUbu
KReD2FBIS3IbFsvDBR2B3+cj2fGZ4YsKvTXyF+KH7ZcOLSRffKHJK3Y+Yx3nXd/u
5PUkA2TNXs0oRy1HNcuwRsVmNxn+Pxx9atlUCYWvczWrh3VasJsvddpWCr5gxzcY
gwX0aLJ5TjLXDP+cFlcOhRkZqCqJP7F2ansKs4drSBolDKT2OKKg213DGWeqG/f3
tOiLUwhVlTcG+x+KsEl+jndzcEU1cVaXYHtpmVqKRW7luw4AZUwMB/GmC3fX91VX
QPjzOY6yU6Zz27/LQxtYP++j45SGIcCnBTYEAaSAn78QVGFRcrnrC308JYAUD7pL
X02+igibEOHeRtf0iA33yQzucsaGd2fBKR+igBDyVw+b+AivJH/rnlWl7dNNqyfc
TL78AUc3Yh5TExKJLo7nEIH74f5JNgY+uX9HjGoaIYG12CJsGeUwB+qSsQSRZi8f
RdBwUtDAsN2Awuzk0WuAfGHeoRoqjOX39QvNdQJ55DGzMVxJihciY+Z5phrP7pNA
4IaUUm4JaqPacW/1iMVIAYkXKCsbuDTIeF46+aKz9P/B6HdGIRRFnq83S8zbfcRf
WLYAkKRy1pmRKi56QvORI3ET7LVzRVetK+Ke1dUgm7zp1fYgI7FvoN2CZlTLuwMe
89yN2Zqvz+vNlcZ15m/YYx51LhefF626zM4JfkEUvFd6kuoWyTQzVV8xpzoFFNso
gkz6MoSoA8vRh7URI39rK8dtzOlp6N/L7Aijuojx0vIIfmDV0GcTXPK0W1TFgZeX
s/rUXshY9EOmYiirHp3fvyw/A+DTR9q+df4DGfXBzZwNf/bpaWm783adAQLQpqAe
cFzqCdOFvqYGJOrkXFCZ4TPE26LoLQIwHM3xdJup2uiv51BG8EsHLy5J3X4DfNKK
x+zzmNJDlbp5cFFDh7ypHJzhBKcMpgEc6k0I8qgj68gsLxauVJp1+9SRDQLB08Tc
7pQx0wRo3yvg1HPLS8lOmLQUFps9t76xWJFCxulxiFPQ74felpQkY13Wtukeb3YY
vh/peBRY6X7EvZTNrnoUoKPXuvL57Gw2UD2WUy3zlz/WpLpdrpfi6a6sFJ6NmiZF
0RIC/la29eYAm0d68OfbTrpMjlE3RI9H6jJv6w9zMb2oRbhtmUk2BGY0qiUI9yUD
UKwsSbitKjkGMFJzqnU3suywAzjATaVoUu1B75h/eDklYKe8VKdRrccKxmGa6lNG
LTMcI/7dJi92kZ3IBlTpiwDuu1cSkii0Ap4GG2rkwF8qvDHTBbJpNyex06jCY6nb
TsoRziWPpWosVCUaJVBWX6cY1EHO7BAS/vSZaZy5+M6Siydg8n8N4cdHio7eaNGD
8xw+yWpAvQQsMpHYst2wscWtWmuLz9HPX5OiENeLJ68SQm0R+Qxp0JKMnFPQvuYd
XqRPAfh3hSNDcitZZjJQbPM5lE6j1ZHLuz5/tSOq9lqllDy1Vvm1JtwYLC+J02Qk
6M/WrmmoY90U8zpP167oSeiRiL62Z1+NBNa37R6xTVupntQtbrgCY6w1x6mLQv5j
dAIOWiJtpbOev6Zr/6Ohn6fENjD9+Fu2Q18tjeZt7zU4aJHHYBUq7eJKWXR35cue
Y3MpDeEusDdWnFQQEMRhI0da/tUKGNOmr4RtXR5TksuhHKhEbpiPydKNvxZz2NPZ
OMS/U5G5BMVLIjCeEgnKfpSt2pfs/EMQa68YiI4XWivoo3uqcDI1lY+PcOX1nJgP
FlDh8ZqRcPuU3bxdaBSL2WFIInnfYkcnQMEkr15AGEk9tvVnsKdafr5kxbLpjTn+
M2rEpNxShSUw6T1dJ+mVuG3RAGrdp7kOWBmlyz+KRLBxL/qtsFFELjhODYWCai/V
hFVt0HsPB3jmrap3Gnw6gPq6WToO+9hX17DmRfW8lN1puoNv53kUnrKjw47+F16K
VwSduEXXd1hV+ecnwLaHqnzFFSKEwCB+qbZmBg4V56UV3ZOIMZKoDs0GcdpggY8S
XeVCBSHlVxyJ4fsirMX4guHYdUHqRUMmRZSS0TPrcuFIq1oGQwHYbF7zez1bA+Hs
99lU+45Vljo+TCkDW4MU3+DcJxTB9j38TD3ojeHF4tnspWfiWtBp50V8wVESVs61
HEUzP5HbXUzzxlYFoN2n9izTD/thuniAvswHD2Xv7/Y12BgxoLH/kN2V3ZKhs/VF
Nq8+t5Q2Ag6XD/ZViKZKCcCPKwY2DTok+AkInKnxF//0S4txHMmfe5YPqF8OWfLm
ueGpB/0aJFXOlJeiIrvwNzBv3j/2RG7+Bc3TTMLa+EnKrb0Y0+6Lgqp2Nv+86Hgr
RwHHRmXOjb0mUjs551ma/T/t1f+fl8q0gYenCiwXB0PZeyDvPP7IaKBJ26wpV/ZK
dXCObMaJ0nw/XY9JyXwTRv1QLbdQ/DdLtbcMj+BZIgG5/bGBIH6O3NIwYsG6KBrG
Hyuif16lq5wgCwOr7hnjDvih/zxCiZxgN+lEHHBg6QUfyYWqc1l8fYo3OGXvYyMw
1ZGhzeRPiLqRrh3a691L52bcABk2I4CGFIn6RRz7gGL5ubfn84hYXjdP4DpAANwW
ai1hRbXeEj2IHaSyn1uGvLjaF78NEDwRyeEkPJc2F1HJ4TTux+HKMsc4JuZVCllM
vB6zMe7R+c+Xm/VPquZGJEEBWcgn+o6jLH6/YIYemcqKdugGOAu2UtGUBmSNF3RX
+I7MMbzvn40mSiBEknZwscrmFHt6KNDUGwPAi4k3HgebdDKlAlRQnf0PtO8USmZt
e5ESu7IOhUOojPvsZ2BHXRxr1le2n+7w33BG+WRSFliMPUmDWNtDKOwRSo13zUi3
4h9ulnWNVUPCvOcwasBMBPEJsNu83mAYnNLHdbxvRATAno22zf/Bk3poatKbLAmR
/Gux7y7vdag5V0x9xuFQCWJQuuRGks3KaSnGnZ/0DDCukbsjj8xFRSrw/5kzNocW
60KIzhd8xIxCuZT8FmbmmkR5ITo2LvzOAufDDhT55F8+3yfiN3PVAl0alhBvbuc1
gcvakNgki4Llxx7pFO6L51Qn7z7lQpjn/ygW1/AC8/JNlM3gRm2MoX97xNNROf1e
ODgD4U6i7RsVPt6HZSRcV1yF2GfHM+l+G2dq+shcCU137vsEnFxkJyio6LB+VW04
iBRkyQwGvWhZM3pdS3Orwhy3etpoNuhRRzddscyklmufM/p6UDd0kfOM8kAa9LNi
JGRYuFsODtiyOqfsh0mFpyFzh0G2g8oZ2rZ3EjVRXeVXyj0SiH4P8D03nSOLnoHz
rcd+zNyTRYbEidI45lgN9eIcL3LsVhtGjz+GDHU3NNQzXWg7GLpXzlM2QFNRzDow
hmA5O5VkOdvMQBj4Z95v+bCQP7wXYiZl3CMUNUs4ZKNe995j5MGwK10iInG7uzxS
TvwP6KTge7f/M3mYH7s2k0BlIRryYyPEmt/dWKTEsTCjEVlFbD2M7OkVf/++KP4p
fBx+Pl4nV5t8kZMfT1cxZUGkJFBjsTdXGOUBMcZckUePy/jH0uvMFMLH0R07jTgf
gYU09NqEKOZRnND1ifWMKJHALLfxpjER7CxxIXuBcPPZW54h3QnUTxrZjr4dvV6I
iGMmnEhJ0pngzwXP/ATnG6p49DexCsqTooWfn8wTz1c4XSbeoDC/HuLJNIvRbaRK
cyUHm/zV4cl22cF88NLN65+RBbS1dup10izHly+hTCM+3YPdu00l3mRdCBSzqB5r
nfI4H5FV6vuZlEiD6qKI1qnqPqDkEO71tOGrVjCSme22zrEdWEoNqVGpS2P0+H/J
WO/HWgWr2Tyyk1JITnT91D+uwWe1RcBSrkkRnqkaAZTltZgALqfXTJvCSQIaqO8X
7u2RBs2DZXs/hDR2ikARO5D6iIRRDGbTglAHgcNOAnQ6s9ovrk2AepykktU7Tjrv
j4QMPobHkkb/yBQFY9fKJIO3nq9NjJ3mYzTINfTnHw74R9z6w1N3ii5zerkAcCgP
uc3/z7IWg1moaLFNB2CVWVWQvwsLak75NJM2MqrqBs1heIFb0RLwV0SUutA8n0lD
f3L0lGHOdEK1Z/2JeaQdA8RRADLYiZ1vBBWh1U/P7WaIk3XH8nlMpktgCX4R9WbV
S49VPOIybj1uq4b/dXy8F/UXDmuGjWvs3xT29uLAuyyJ/9vTC65BsSZOeK7I6WCK
CEfdXYv1le9hCkkbEw6MRezUKtt2LJVWz5aWfCm7C/EfZNuvhoi4NWfMmrQC6WHm
sE6eVM3lcxTEXlJGxWcTpAJstuXJ+LkAHv6cwT+XDtWedsuv7pwIqv5beO/ph1fH
0NK3nvos1QXl6daUH0lswnppbzSWUPhQJC342vARMkMxD+zGiGUyczQ6qvyqK1aW
/VfJRcovifWdwyo/LDvx1TjNhrZomXlEV3+yS6eJleu9vzlsa3QYfbfh99t1+hL1
TD+J2KAZsIlPY46eZPjy3SxzfXWrJzFgeU7LrjODfMYDIGNubEfBVZPJZLij2B/P
To7NhO61+deXovnLx5QwaEC8mecAxkUooKYiBPAfntNDwTG8e3GnBzlliPUHum7t
rLB9GFqNYRARuBmzVsDMRrArBOHY1RxxJUnkAEKBDeooMDebjGVb3Ut0Y2BaAhYR
D0r2bRMPuh+JrkmVRTMvUn1jOgkZ7h5+IEP8crmvNSqTe9RVG5JfjUl81iKJNNzo
cGr7uu5ACMhmVYerou4xc1u/qCjMxkSVnmfziFlzWeVtEqTo4+7Dsc0Qhy5+4BU5
cgxacO1PThgnj/dmyH63PIP4FpNUqOJBrq/bmivTvLBnku3Vf4ln5M7ExTovv7uY
BrYv7OLT/pbAKR2b14SU52St6wSrZUYwiGzQpt4LnXzHqW73KHz55u4u9+IB6p/R
/5nRhLWgh8shW9bQhSmrsChQw/q1d+7J1y4gsqqmOqDGgz4kJuB5SEVcV6RElcSe
GRvrdQx0sFcHK24cRGgA9sG/6QqwAOL/dnaMPAk+jaDIGa4dI8EP/dVPNy332lZD
Encar8EfsJmr6NdR6fsod7VKi/Z+mihJ1FVjmlcbfhITfPFMKQ2wV49xiuIS3ZKf
BUvurKFvwl91EnQJEomkyv6+v2y5liQLQcP3JAc1DgSQykCoeIDpBk81ZLCV4mfj
LoI7HV+CmyvF6sn5mebZmLAGAuXx7+1u1cWzOT+tXeBZagcrgPNRHaGWPEu/X+0L
O3yff7VCc39UBYwFdOyGc9QZBfSD66mckDJd3lhizINWO/ZkAaEVW+0hx+f3IzD8
m/9R14GgWgTugGJFAS6Xvr+fSU1rCqxsoqnFy1r26Ug+Vbk4ZPflC9aMEIa4XYbT
Ui+v3DKHE+PQ3GkmTaCRkN09RZUusvWnkxb6U3RPhhdymuKupf+siH+BaenRLdwm
fqBsuvMx/xaARl+7UmyKCT1MjY1V+yu5WQM8vDkMCAgtwLn3xH3Ti24DNG5XhoA2
fLRnY0bc6oRt+3bQAL5gvVzxxDSIhEUbV+uMIQuzepJRic4qLjnoAQj3m9M0pAJf
aSwrCPQY2hym76+nG5oU9YKELjBJm3nGVB3GOuG/XBgisxgVmBLhS3T1HHe2DHWa
Savo+nXdSwyOOyzzXahfw3YAZZjJaeWvW5Y4VLQG78tIxijHuvotMUeGV3al0Iia
fjJtg747jvgky2zdBKY5lduR1JuRQl8oeGRA2Ch5QNw9LNxhsbs+8FPjAJkpGIQO
Z9L6datbYX6W8q9+FFtyZ0Kdv2c/Ev9WxqsTin4OW7hMgFrvDrgS3bT4YP8ynTxR
tF/7jO+yrkfM1I+H4tRjsUVHyqnph0snL5Gm8ZF5oBGRyrdBf9TGlnWm/ZRNT0nv
OGVVnKxvN9snajTUfeGoha7tlB41FcgY87Xob2EhbX8Dah8IOZm606L9JZoGi1nY
SLSaae6ROylsnndDlrigr5NbWxsaYujN1vlWI1uQMvKliFgE+SyBdWh03gFg5UKI
pCGO6uxazLYWqehvI3mFmyH31AyBw8SYZzmaxpwgvTYj0y6ppeRfk0HEBHZm150L
pmmriADUcfayJJSMwktcT4HW3oTHajGSieXZKlYDIUHLpZl51HUIl710LAfBC5ua
wK3Dg2ohOwG6sI2toS2i2R14CzNCBbzm4ad2Aw6Ib93+5yCXtLlzQjkcBTULisf1
5eo5a+o5yEfwmJ0gpaktVjmvZy3r50qj7X83oyzkkiz0F1iHQqIBjvEbSZLJwLTr
gsberCarkm0lsM8B5b8JL7ECrkzJ5pOyIV+Ov9x+S8fypBmsuGis12hXWe4YL1RR
tVyI0RK0jwMwc3p4NqL+ILkoJn0fWbre2lrJ1LbXbdSl4iw5jLrBvFYSIygw5mBy
brUBRH+c7Dln1incPJF0wLSrNNseBvCBraRTDYM11lxVEe8ZUxyTJknuoqeJgAwF
W5EWbLmVCbk2a5JjCz2DUb3SaVd0iEYoshF6ciDWVxm1FAdTYm2ZCC031ZgpA/4e
D7KzuQJulfH7ldmjjqmGoRLW1xBeKf/jHJt1Ip75EMAxdxlTsn4Q4Jyb6U7bEJ3x
MoUssoOOsQQOMA5W0vfjbwjqlzCBLL38OByrFKkVNFyZw6O7Yru33zN/khGb+5td
aVIAMo6TPiUXRojebMIfHpD0dmMY9cBKvDl3mWpKQTjsV4Wlc6CCKvCnbfuaalCt
m/utX5GVZ2z76TsvbhfIfDScHgLxz0JV24uSoNoFtRlVgU/AMlyzz0qzQJUWtdbi
9J3VcoTG53nex6RD8ecyzpQTCL6m2taMEPLT4s9f6JbvCrsq8tiEWrFr+HkQqso9
at/8432C9q4Rw7pGAcuaLauCkmUvCIluHYInt5ocNxgH6vMXGtWTozWOXpuU3+Cn
riEEhpvqk3l9YrOMwLbFHA+L6N60ObHAMakncMtRswexi+guJfSlzYlKELoLNKuw
nPJJ2waG9If2kEdO9UH5MGZwH0Wja/KFnL1HG6tbuRiWWKNWoAFNW+JXbkFdUCHv
Rs9mBgo5N5ezl1+i89SHSZu7cMcIXouBFbdqhDyN0TQ731lL2POBAQ2T/YU+QYpZ
ahX4UaDuWtvYOwo1VnN/rEgqJHaQQWL+0AVKHxzPSR6cOk8+0YEObgeagQMt8HM5
iKlDk4J9jjMZLAbWZEtkUNRe5tdeVzeNOe6uRZVv4L4hMt2WRHkcdF9z/E5atX8a
yYnuZQUI+0gUUaO0XVN1IrD/F8Psoy/H4FFh8SkopWMBKICpkuvDtPLFWRAR3KkG
VqP5Yd/SqW61u/2zDmu7EUAIaP88/DJchteQnK9Anm2sFt4uEENMGdFCODkvL1+R
58VAaFnbm7SpCwP5x9xArw96HDfddbIKG1OuJghGRNxpmCfKZTzPseXrFYscUYl/
tlVnj9BPv3W1qW8DU3ij5EoGEXIaU2xLTREfxPv6HMXG5BRWyJfgTIwk3Wit9MNE
EaZq/4XWvwJnmzALJCsZz+8+QrEVp7/6fueNVhDFGVcDSawyMHn3ITLiwftE+GVp
rlU+PmGJ3yhxjAIl2De7cVg130qC9ngLaRVnJJQJm3VItFk7FfWPBkpf7gBkvfVA
TGGdc4V+zVOXQnYifTGBXY2QoKtb5pPLWn0ZPW9sVKB6+ZECUqRRFohjABZKmfgG
hZUaFdJIqXbX1HGTHYSf1b+g7xAgNKvFtZPGeX1niuh5HOjN2CABF6td8YLWmlam
XxzssQN+eplZZLiY8rOfBOC3TaOWhl2ILj4RmculXECfl74L8WDO+p7P+Lj1SRJs
K3RuHvKOs7S8jSS8PDlVWTSLQxPhfHnuEl0AUg8gxeBUhf+HceWC4mEeURjDmXu7
3MPsBvJlDnrXmRU5BaG47hYrz6Uq2UDsiorDf/NJF1Aqiq7ZOY04Z5sAfhO7vs1A
UFg9+ezeZhOb9i96bJ9SYB53ImwDUopzwIygv1izYGra5OIjpQDPyu6abu2hO0/h
Th5GC6Qu1ZMlAlMRGLfueZT8PAqd+wUutIlNrQtVMohpv3UjiN8U+vp2dRhXuojz
icEQRda7xqDzKuF3DY6MgzO3/u4EE6YYKaHvkBhjnKGUziybnUjF+Tl4HiERaq6j
1xamWFZyc0q1gV47jf+hfnzmhmllSaG6w2pGSzE8z/3M1r/M2c8q0k8P2xcmDHUU
qOF+ZXPDBH5zxMKe5Y2Tnv2X9yXKND/4n0QpC6Oc0WX2XI6AWYET1LKBXwV2qN0O
01vOpscLCc94+64MQNjqh4TIQT+nb9/LkAln4YwWMlyKZ2dudRp2fD1dNLaixMUx
uMAEw4pYtn7q7iQ1rox5gPRshiazCO5wpbT5EJxjd8vdUPv80z38Im+memalTR2A
Kz9YG1fM84t0vJBIAkvrXtNiIRqCAx+QMLLdzO69/ZYH21NQonyF0u41rS7EKck2
knrkOrF4CjQP6rdNLEKHjsaxD1Q+JPYsmfjDCi9J2j8kxajmweqPIHoc0EVQiHGf
PHKCeqrkYO72NqB6+EFjzGuYIZbIHsPE1jzvoq6IQXgsXL9ru2WF+SDlkLLOedUy
r0Yog/12D+uz1qeg7sak1XXRsMJhrgidCvg4J3JNnrRgFcikBvebXyj5TPy/jobS
xcOtYKxHvkOhlD0PQhUxujxUy24p5CJs7ZFyC8qowO440/xJrswjPO4SO0DUDoRR
AlO35q67n8ZaYx0iJZF8vexG00H8SceWmS1ii6A0/JDqQkVUVfgPAcDJR34Vu0aE
6J+kYYqoDU7a4rQUGFFL8s7zOxqmKdIhLDx3IiF8Gioi2WSllyDJTisVtc45Ss4r
1pb6lYNkXng93j7g5iD7axyPfGTYx22zMMs5MACoosy3HPiIeJJz/ix7DSWCAG4E
Pi/mlOpTMYTsV/S6gm9YpaP0qGGsIxVatevSuCJ28vdubutjec23iPu/abn8o+KI
fcBU4sUIUkWb28bIh//OhxEBnHUAE0BFFE0kU6pChzHHY34IH/JqVTvnqQJxXUbu
bRTfUm7AJ4JISorbV8LaZ5y9aB3kBu4zxfD/AIlyvMBbL5nK2Q4EC8O2Yuf4YuSE
2mQgQmEFauqshnq1E5P8VRDqXSuvR8hHq3oAxXjDO2N+Euy2ozVW7IT+OrIZQMYV
xnfXuhQgPM1JBzAFFWiL4CckKIWK8MYqJ21J/NIX1Fml/wHBG0+UTw5DmAEqYjlZ
oZRM0sdmG5CvaSbnT2O0oVr11fuUuxbPY4AtUgLX8Gq5yMjvY4C7KDkzDz1wHeMy
5lc9kI0jxJXV6FroWse7FpfnuqCz18Q0+tTpdzqySWE+q8yYJtsbeZWkKIENEeog
rBU2s1bYEULZihSScanOKRGBbJF7epzE6ckSitfEy7vT4bN4DwwlSwsOLocUuEXh
kjUT235SnzH4zwCTePOrHpUMs1OpFgUm66VX0DgtHkN5HnoDYiqOOvtJDxXFXo97
aEXkqG7cy8ujFDNid8Elnd68Za2hOZ3+cefwEFvyPKmxFWQvGvdBgjp1lu3Orocu
Q52Hvq/h0sWeuGxSAYR2Pj/sTk3Qm27p+MHAeNCjiAZvA63dfXQcdUxtgFxehWc6
G4FNxG9TBKgXbd8AHSRfOVYaLCHrnF0i0I+x5kbPz1Q5DS7nvgF0dZ5YWUq5cOd3
dnmegxDtjP8QreuqqXxz2Clg2LPm+f6SuhEFXpozJ4MdZuNTHk7yYBQvpXkecIL+
5vhWHKSus1q41/VFz/9YaoqU0CXBxZcmaa2AUEjL+wjUoBQ978bYaAG6P1vNcTY1
0m4wTFzwwnE6KPLJwzjANbH3rVFZkrYBwHEZHZY1Bhk84FRssEffIk3Z2+1dxqTI
jKm2QzjXg+nMVh6pQ8j/D8ZP8ZUd4tHF4taeNarxh0YTOXZsvDztS4ujpGGisEZS
xrBbrHRb/cxQYKMySHddHJnrogWrKhmeEC3IJx0oM8VMwjqAdG7DiKYyP4pniepg
8CgvFsEXrqi2kEVgolN6zfHkCeiMMB1aKWIsw1XnSn+/un0srDg1z/27Ac+v3yXu
Dy/2DvOPkkkY3BamXDHvBJO8QUqTHOegRGl4A0xxTW8gCASE4A8FopYVflaKtclL
5Bfp27UkmxaU4TsyNVtv5OosZ2YU71vdTGRVxFvADA1Y6hRGIF3HT+888lISxggp
e8xpcaBCqH6OKso/debhDEHcrzBrAaYP9HnY1l1CZtG+n4Oy8Xdas/7oZUksZr+I
ACweAPPJxULXe6MeUkYDY20xwAyHHZ52qDRqDBUI9WnQZMrvLONgqjigg+IRMlKH
TVibMpq2eo+hZVpkSEYMCRk5RBVUumVLf/CkvKbTMawFUaD5rUx5vXbjEpTFR/RM
vy76v82t+sR0TxqL7c62gQVvOzhqCdU+Glx/mEMRrHRRXRYjBDxyzQkLsz9KZUtZ
JAuSGG4Ywqqc3++gt3VZtGGUgzdKKEB4mD6OSyt9B1FojT/DmSHTjFmI+M9XiCXF
fJjOa1Fd/IcNsZVwvaS5tl1zXx0iBmKVWKn529k0DJHxekfqceaFVECUT+uz2rTp
IoIPsLJNUQPjOJBwfJxCe4hgMNRQRKKJtRqU1lrLjLw53a3z1hLjjArM/F5+0cLo
9N1BFpm8zMUWLMTDYPyJQYsRHanQyWUmliPumYXThNlzuqZ/o4paxEh0MuseqsKr
4ufA7WelRY1oMJGAb2brg5fI3IAlN+GzJHj2mQcoAaFRdc+HKxMnhilFR/D0pX3t
g0XS+HhKSQklcGCM435OfqpruFfxL81mP9fWI3EXzzoUncrvx7fQ7YIfejMUY83N
6DukuITkwyZbdaHErcbtt/zzSzP86V76+WF4C+dd85UimjM8UmWaHz6HEr6LSH2y
MHP4G/XNTrkQBTmDYaJVhWVb5QwZFR+8yXmiuAm2dDss9tqEBZq0+wfe0wLAx2tC
1fge0L3PGhVwiLxXvjApL4CEDNsPWysE/xx8AEs1lsvcgLU3Dxx0VUKgmbbXMLje
E+rqJ+NWblPZdUh20Q7dLe5zTos0jHa5cNt5SJyQQAp2vqQjs/+D1xvW3y7j3VQx
5ueIdW2Iyu2EdvOC1F6eXEw8zUv4twxoFTCXX0WBFsTYKTlsbRO3/qhzo2Z0v+ko
iC/Jbm+EGM/9/7qCvxckGqnonbpugi+7M8x81T+WUEUU8HklS3z5E6R9UbXPLpbK
QjI9iYJ2Bkj4k0/kmzyotbFAotqrV3Aai7mBr9owyhCVPwnCWrKjzY9wNFZ5N/hc
HaMDaDeKE4YKJyfitPiuE/gDHmKbZnM4jv111lyLlTxo1zPBUPS0/00bF0ip+GUl
MI4r3e3BUvHEbWtzpTG1/fa+PvXraA47TBXZsS69lx/9NZgJILF1UkQ5NQlKdnMB
yO0DMyhNQKPrclhyIHwipET0wjlnTMBkaW0Pa1+AJWCdClhPBAqarLigMQ6ZFT6d
e0lBhzGD60HJ6EOAXDDk5aRAi8FhuuqjjpJ21zd1PMsTFvtq9glkvZc1gC0MWjTU
dkUwC2SMvyZiebWU/qHyOcuk+k8gotZ6fjYfAeEzt9RRwK4PdE7fX6MqfdJKXzwa
WhqiSFlURkCibcXlvL4Csq5oUL7PX94pnefg7PFO8c6Yia7m0F3CbFuYtpVbj5F0
7gYn7lhZiBJHbRFs3iKgInPewtLmRWukgJhnNlZCKaHnU/YsvhGAM+Go3yiCrq3x
bqvwCUMQVHoe3Kmnxz9tv47stx0gmJrM4f8Z16PthXD3WUHvz7mp8D8evcmTsCCN
LcQ6e4huBaZzeqlSfjko6CDl662i0Gt9dCmFU0I+ACXhlkUI4m2lTvJ/KPK+aZHh
fvqWmeef28gagfPI/jQHKnTEFQEL7xkCUokv0XFgft85DfAGa54/WDVELtITadh/
8Zl10shn/GkTW6Kn51n6E8BZdRd2kG4hSUSR2AZPFs1ZdHPMNCUMGGTfDgKvqS8J
KXz+uuFKGtq3ITm/uctaUGpLrHVTvACHeLndSMQToSKlT+DLr2M4ZTcerSQR5+NW
AgkBSQQV+/6/IC4bmVB4Hs3mXhPYKkwh2ipBFzbiAxWTdWVxaTvThdu2iQV1VwJ/
iiM6NXcmzTLSjW5Xk7SRpkk39tmSE8NtZGqjyTIgEJrSCISpVeLobskvHIp6JpY3
bcBjNVI4eozL9kIvI9Q94g9Qk3P7AIkX29oKYY/A08Ihyt1cynlFUWQCG+fnD3gI
Wz8n5V0UWRc6kEWrAn9pvmUeDhMCtrSFlquFSo/Z3hAUCC9MenkJN5iLhbi0gYkk
an0Oudbii9cy+T+RU4en4UkK3FrE/0ubb0swhf00e7RfgSCyQDbplaPSDMLC7B2o
pxbX6WOGaKaFXpESECxAQt7D5gD3NUhcXLNVvU3ZbM89R+VTl9vjhXJp1Kn8xhdF
pBaYXKf8aaN9BWqJaGOW+FXS8K95Ck3J3sooHoHcp/SqPldImaXe1hnaxl0C2Pqg
IKt39OuyCcpyloBLt7adBNekgWQKxe58XDh8FL8xImfxgJwYD16y2SplkZWeLgrR
fkl4he6XlT2wWuab5GXhzgPrQUoA0GCeG5zDlO9stHgYfJcaPK6UTcDNQhWUwSlx
ORmifNkz3IGuhqi7L5U/vcft63DDGnPCO6aqYqOAxg60+GIKPApbw+jQ3YEdrvOJ
31y53P3jzIeX60/ku81DJ2Ah9N8F7wlVnIbW5coAFB9DrID9dQZYLNRoS4WIUTXL
VcfeekFb8HGtpTLaTZl8pgIGSlBVQsu+vSvKOkMu48b6Kn2F1Rar6DLAL6j8qql+
84VLMs5YfTGsDsJi8TL2Cr8LdGV6l6V0ZZ3+VwbzXuTNyxx02o4MI0nn7rqssOP9
3f82THzDzmFe9jF+AJjhmyEu3ejdv4TR9jWqXOxkpcEyUPf0Xgxxhx1UKMOwlg7f
+ACfU5u0/7pV3rQfpx55C1J7kIs/hRo8RV9pHQwRPUaHc4KgTDFGzawhVY82GfUh
LDvqixRaXMTG6gxy1zOPHAL993B0CeTsomjzKZti0rPvJ7xIpEAVjp6fIoctc9W7
isHv6huXHxFF0ZZXLrrPnezdMr8jv6B4vmuuXwhsjbaBf3TPNmG3mirJCyu3ohLl
K6gXGlBK44cDjwY0agO4hcstF1HLIx+5aNq1XG4Ze8jrwHhbT0IWeRAP54G5ewdj
6DW1GLdfTGFo7WKCmovlijoxSRnqsCIOKhXKZA30EIxQGua5zdmXDGujhoX0L1i8
4sjyeBiaKHEE58ogO5xWzEozXqpAyfjUJ00ggElzegCWAUbbf3lYhc8Zv7IcY2i5
2HrM+FKuuQxeeODJ6STUnhICBgJIKXYLAQPpJZSVMlIlVt00pdRsZZWJaTCZfoOw
csJaEsacJhIP0lTutuXIg6zjBz555Atj0WzgIETLKNM3BVc+u42Gobw5S19saj5k
PRGeI+sGyHr5GRboSaj3op9eKjSbHx1pEV47Vx7YicvYRdHA2WxqfdzZrOP59QPK
qS7CKvxUzBNN+H/0kqyj5e/qkmZqaalsrrhNS0OXrdbN83tiYOxtH47hVVmkilkR
vW638v0GFdmtfvVLPMSrIukzNZ+BxcDENHPVO/ST5WOHtgeTWyO0kIIKqtOL/zdP
uO3HG7cerb/pBpr++AS+7sxAFV4nXTk6a/od38WVIHwsp0l8uFlYrfKdPoUDGxOS
yDTXu3B2NYhOVtIDve34Uy6Bx2mvsoNKR6o6JnfDCEnH/PIvZdkXUIT37zQZUmM+
SPgo/5yRHWaJWTvlxjXqL3wwlWTA+lX5SZLjvbv22KLJCpgVS4rO/N9gN5ogPOAj
4OOR6jZfTmY5GukRpJu2CcXiEvaDTj7k1EyMTJ8ZXl8uR2V/Gg42T3Ce50SohafJ
khioJR6vAeOSWnxHW3pSSg/i/4zd2406FAV9gxraVHgu2uvCEUvymxUGa3RdwaCT
tZihLq4q+Q1ip3ToOyUIOOlyGodiNGDZHhArf/SivKSZX6JDHCWUp985YF2ope7T
28fHsxKDPoK+NJtPJP5kaO5iQ1CjoXcd1g2wufRs67vcOct6cyeI3XT6vevJ3ieb
ofmEAj3/oXXpFjxcAd8VmI/JK14NpqmRCCuol5bn5q7GbV+9PZbMY4aVA7okzAyH
OAeRRlJ6s5cQk2M8X0QqSDgixlzC55s43jkwPhMilkJ6gnRVJ8BTc/jTRlqMbwCM
rLxJc0/+xl7LDXc4XuF4GK9r+WfvhqazzhzEwnn8Vpf7EpwMweWpYQu5poIic0zn
pTFMgBKmmH10TSH0XWnrdnzHCY8btT7bN1X/sl9u5465VaV7qRt+uXHGcc8ptbiR
Li6Vi0ySPz5SHQUncWtwFzLRSM+viiPhcVZpMufwjDroIMhGRLySJgqbXKO6KL59
Ecl/eAA8OFn0qIA/712F0G0UUyyt0KyNOzlTlDTvZkwIyyEAMtIVxStrLJJzG7T5
D/XVbxYSMUqZ0bJdUswLcPtO8mqsqi5uef8/b2IcOzw2LU0EusptsYlf4CDHGhGF
2dTXvxBew6yTygErSYqYKNsVaNfHQtHTLRQTilRwS+s+acsBHIi81gMINRJ54nTB
UGo/Op41LfBOVo9D6atNRsWEfCct+XVH0UDH92QfBd9UG9Et8tudN3Pp6QXobW5p
kYSRAUtvJQCA1nCyypgGol24rPRJmpYddHyoyJFjwUqyHYSEf05w0ZMdfKljsMVZ
Ri9PtSqKO3nzykJI7BFA7pN6azRfv/Vz87sq80jGbb9bPMOhUH0CtW91wnw4SsqU
YYtMs0YpObIBcErdoYRdZKHA8kaWzp2ialAI32d5aQEa7i24+wp7Leaso4j/JSFb
5Ni+Wl6uIRts3/pLG68F4LV+qB8QMVxE8mMn1KRlnixe+JTrRWFDO6ip33SJCp0H
bCD3sJPWrgpoJ/inB5iV2+X+HY4bSVcGe+GJQpyunqFxARBgRHsN5eaufIipCtoL
3ZRWDAgMDToOAIgLbyvyuZldS+uuywscD7K8j99Ma9UaoBsfY+PoHTMsl9prcGq/
oS4AQNfdMEmChtY9GcDggBUgdUsf27eh5Fwe8vyIUEGCPdGv8zhzVXVVViI2wIFj
lGnim5T6Kw6u7Xs6CHZqmdsT8wdjcT8bYe2zUBTTXS39xp+24yYN1TkbwMXga1t3
gtc0ne2bLOn0QlTYTEHxZBPpHJBEsb50ElEhxTpMzimpYTu/Of1mC+0I5r7tWXSj
wx4dIzUsSkcbGVR/Vbz30GNSo788Qhm7jg/WznjPhLo1vEDBGAlJLBTUvoUsdJxi
KPz4r0z79k+6CTrhpuRiI+m8jFxW+MYyLY0WdTUwxXWb7B2B0PO5kFPoTwxkzZKS
ZOVS16ViGpXKQCdxuEUegeVK2a+r3axthO2AS3e3y7F3bWq8zijZ/1JHdFiKzpvZ
9x/H9CYOShurw8J+PfsI3xe+iiFD+Jj2sl6PeaBDstWzrCZAchy6RGVOlWWWBi2I
xavvIkpvc9iY6+o9HRlHBy7/dZANrrw7zTxY9UJidZHfg1F9Gulsk2CXiKEaEuy4
siPJk2LsnTwqoA74yPkkz7XWrLSvUk3b/NtBs1EyEnPSur8eg95FyIL5PhU7ifhC
CPajmAw/V79jNK7EDwuZrvuIuPOWIy6uJeADRpI+Box8Uoayy0BWvleAs5QrJQj7
3Oc5jKD8aPl1qMaYOqL9lU/SUwgjjvzXnig3Xb53VeqO8U7u7N6yLSNr/K5eIrC9
HlEmubPfq/ctJcbTSuOvqmoKxriXEpO5J2auIHjqNGCFyTjIgVdyiWIEXN7C60Ca
g2q3wqThFGFVcjH6JhkTLCHvuAReQm9j9jvLCsTItRoyqIioamB6Rrn4BEsfUfcL
9T3LSwrPq1Em+RGNGCQqdk4mLBpRuv49pqV7bOO5ElqprV36a2LoH3sO4sgm3xPg
CbG2FE0vAN7LVUxMIqQbtVq8iEh7a/OJUyFKizj7n9tqCe+4oXiI4SBq3LsYGGlv
TlUwS9neKAnTowfFFPk/79FB/XOF7k5r4z+mipfGY793Uva8Ii3y3Imc7qttu/pW
rykupyNxr8jtF97NVOkgqoghuLF79Nm5lI8ga3o13wIuxkSXK2h8kjJN+1vgWeCD
16AaEisZW5t6NzPOhIJAUflYqoeplSOiRoH7OUGWuAkD2u8XYCQZrS4QbDJzeGmR
Tq5mmjojyRgbM29nXL9K9a1geSJp1nCCZIkmLjWfzTPpwfRW31wRtF3aoCLdy6kF
3hz05hSJ2oii6hzGYZX+AatrIAO92neq38Z6J/4eTeTsTDdvuyz3CV4mAus8brN1
R3Zrx3b0QUDRN7Fc3RBdtn/qECpAJiexOVm84WBBsL5WTVYIUWX4MzvI3PRSuKWN
dQMef3Uk7lFVG499Nr+y6NJrinvBnyauibiAd4O6g9KwVzZcvKzz+Ln1u8lD7cZP
NB/zI/abvZFPkwsiXVNiiwKN9wZ473PXTawdDAy9Bv1dL9hXROcXYJFBAfqMntM/
AfMdPJ+QxLlBKH5G5zQIdSMLw2I4dLur8pYJuUdviwdsjk+zuYiPknpNlJ4DYrC0
EOvpaGM+a1/HcqQbWAnKwi6nid2we93vSQS8ZjkLLvXI9jkY65E4lLq3IG9kMsGF
KKPyvyC3vFPa3D+YLW0nARc2ZXgo171iUZHvZsv377IRaOsdrG7zvwQeNe2RraRy
/zN5i6TqiSgnxha8Ko1+VGCecZC3sLaPBa9Hjil453pInXp3Gpp12Wp+xBM0kIQH
jwaAPSt04gHMVuXhW5evmV5ksyN41amzR256MehMh5Yz0MJjKTw8yU0VwVpPalf+
1scUIYexGSAUrfrFe/TLOS4j9Fg7CMXZ8W6x7/MILVE4O3XkZCjGcBuiwNlj2CuK
/fy5oxlbkpW0dKURSA3RbNM8xj1ikqvm3U+w7/xYzVvuLsHvVFqgngEq6slvjAHC
nCi0VhHEgJHg3YdRTK2LdJNml3ljKHqEPp45A4HoevxEtG7c6kg2kF5Lt8/GoaTa
+basmk/vVGhDEaWJbJfbD3OPThAXZmYdGUN/UMx0X3mJomw+JHnuA6Z1iJoPF8yz
BDdZE4CYtu0adMegE7DbXWWukCQlUTFaMIa9cdmRVs1js2DedjRgRMHVOl7enKzY
q3FjgYZSsVkiLtuuNTQSyZOImZQ9wlybV2vQjzmTPfE4RhUEEFES50mUBdJONnKx
VHcExGjC5Kq5u7KHpHUUoZczOOwrqeCgWQ+hSoa0E4VBicybMqPeaKt5jvpGgqg3
5Ghv4/J89a+MeVWntxvvq9SdUbxSAychTsxzB9XZN2LEwiRoyafuOba25Rw1VoPR
cQdcTXZPgNztNVhJ+jW5jhhRt6gQvSGz1OsuvUFoJ9LARBzQPmMYWbFjQOJZMeU8
at1W4opZ4IDCiYxSn9agw2nKf7/IB4FopZozZJ8m4OFnr+xcEjB6ezeORhA2ONDC
pjeOmr8lphp9j/5YtSUVUwNeAFVOAbeq26fYxZecSGWp2MTevPUoJe9caaKeit7P
+CVngOeymCHt2TBuQRYwx/w1io7YNeOsLR8VmrrLLE1l29Eh6Gzm0YSJqfDyOvCJ
vW/hPRXvd+UquujcGhJWwfQ4XWsGHiKrbgdEe/6vKpJmQaY+WQqOqTq0Wi+JZCju
+BtcxY73LjQIy20MYJOn1e+9TM3J/7xxU+66nrznWS70WEkaHtFDXuw2+tPspklg
gfxxTHHDU/cW/v44xojxDQOmWb13jSVmGSJn18IH7ZJsos2DVV02PD1eRJ5PWOn5
NXiYeL5bgUJ9CLLzBcc6EtlsjaSynwvpbqvNYlTUBVSUKmQTKjfQ9OLHa1JJuYYw
XZ+4Y1VSFTL2RCaMftOJ3V/LLVyXWkCzdsIKbnQ56FxK/7ssNaHAJ92zMyjGjc7R
nu1fl0LDrzUwFOKLvHu3oUobZLny61avMN2YQwdlBnnJ2MOpqNX8IyW5936GS0hQ
MPcIR30YPe84jK/RXOrEaCZoPSTKWl7wanSnNlx4qA5xjMTQQ4m0Zmxy0SXQ7SWm
rhI2K4F1K3ixAfH+VFrSlgNDLP43mqqn9lpi1x9gbtWXTAL1DcJcXpO907hB6Hxx
RGvquqNfQJR9DAMPVVmxkabAHUv4xi0WPI4yGnWB5v33Zv/tMNcpOcOqHUhW1cUR
IuZJW6+0B51/JImYHL86EVBaNip/fX5kE+N2Y0QKIlW6NqKK+GxnQLWVpi7oztyp
NnkvYtYaJEeU3WQl5zQTonyUM3xdDWDdB3Wyqa57pvQwkb5CtCjFu0EA5wLJHxgh
KvyT1arqANDC5SsD/7OYkEGSWlefWxxm+UKhVZ+cfU2emXpGbr+AFNkr6NSbdlnA
YmZG6+oag/MM69Vx+c2WLDGgZzCUAf5Qliqgt4+iUNGOxS9APsIgvpvwu6niUAtp
miNa4swpsV5eQR9bUv9/1xHi8zeVxN14WAYRhDTnolyevwf78bSjdX232b7re/ES
gBNSUkMukn9d8khJrM/OdZVE0dxLXEBB8gMLzi2DPldrfJ5fc4QQPZgtX/PxwgeR
tXDh639s45XkyTyXoUdM30TDqxBFAqH+mzV2dUAmXIU7EC/kcTyYL7TuUaVn5LRp
D//CVgjHgVEeQsFIBCQY1g7rHBHU3akLOX3Ik3WZ0vFxTtfOiYqnTmfjK8+CDI6W
V86mI8vFkUBmVm5HwaEA0uy9cSMK7h8FlNP2jbctziQhB+AtSWBvrGKDZchFUJCR
NqsUensWbqIzUE5Sh0XrORQNk0h00/q2RMSxd5BSnJFV59OvrQUGDwRjBEYnpRgk
aj/BdP/19jof4iqgrFbNrz/Z0r5AbAdAVF9fsQQZMZg2aviwZ6MWdCxjtKVighPy
5CqxNcwAzYcjCfPDmctHcjd3AMJmgZl1l1lAvEKnABX15ZM0/FtB3fBvsSxbi0zF
3Z0Bbb8K1p+6NcwKfswQQ5g2ERhjnkDGyT2ztRFTyay6AksOFeURwZoGxtpdlODz
EgbxmVIWkkuYxXpMj/nf8LSKI5PdLKHNssCF6Lc59J1yR4lruKUPyvmkYaYD6qDM
vLt+rCbpM1z/MYjJvfkNAgIRzk+VHwE+SWMXK/Y1wgnpcnqRmja8fvioHU2evKOH
YEtOUqSR0Q0iFlaQc6MlLZUTTP/dwxWjVKQ9leCYbkFFBDvfrAv59sJaLkS/dpSe
wmReABITiK0NOD8n9rGqUa0ZmY4zMrfJpNkrrBonyEDcQmopmUFRFsZJd6BwMPgk
MZpaAD1yjXLr5PbYscOs1Tw/cs+lvKt9DchGJHZXH/vVzFaXq39epT3y3i/veYL2
lg0ZutI+NRQjts0RDI23jzYv38uDq/tSiCzKqgpnyPrzIzTYr3y+xSgHz62Fl3sP
gGYAGGoRNbyL6nCAPDAoDGJ2TTKj0D+lpWPOS4Sgs35QHBwEvNvAQw9paNL4Rx1p
oMxZxccKzj/QjL92PaIo2roor97aQmT9SG9nefHflkVd6wOfiJWJXxMuE8I16G+Y
jX0LqOECw8PBZlSd9k1cohlZm32k8nndBN+iT1r5MMi5p+mZ7eI4xpjh1GARbd2t
GWdeRDIwIMiP5a6062LM3QYM1Bvmgj1TdF1aStBdkTL8wMyZSt7wJC5+yEXT8BPm
sguy1Dh5RME9SUw6nLUtvZA8WY8vfJXWJD6aW5k5QqxiaTklGheVxMh2e7/2O0+j
JEoWW7pPBMe32NFMYJBlnAu4TUiXCRWB/v5IAu0tbQUcmoASmJGO3k8b5VX+YHBH
xXpqhzmu58fAayYOtOBTvGFwUZPbjOJqnwHTYI8cpp/LEBGufdaaKfLGGfkbWRml
y2wr4sQE80A3wwNXvJXenMptE6ypGwt5KRXaPjUuhBS77hflM7gWQm6JFiLM1slY
0f5KhJPtuy9Tl1z7qPRwIylI0EtqYcCjW+IAMNhA0/bakD5VDbf1WoxAabxdcOc5
+mWrPcDJdgEGjnFrNSGmZeS1KKguG2mgakecClMAHyAgcAVnGgjybbfsa8kpYHUt
Be9d6gTeZJ8uPGYydgVUGq7lU3XBpKU6huOcS0BaevyZCCbHg/738veW4+SuOZO6
gx4XJyX5FVrohokrw6ExiUzTJcKQOMNViy73KOIPuPPxqUXVLBo0yOo3mwzsJeHv
I/jjyHf6nxWhvDH+0MFPMWm9gv6naiMMiKNeWieto8lZt8Telp/Vzbv9VDpAPF1F
I6dtjBNuUh/MHRSjBm+Ymohq0FVkKmlP0FHSMyuLvZOXmLQGni/5oh0hej7LkXMG
ms3KyBUvdpsFkd4BtR900rg2E7vEKhe3CxxpY5br7Afq3HHUYXoG6AqbzQh4kWW1
1/is/0tlp3qfoz+3K/huS3mjSviUBKL2cRB/uhOCEb+D/nDXCiREAV9MG4VLEWm3
1cM2p/q4X8SkweXH1vEatPrcoqnZ5QOl0reOgMR1+7Mwje0y0/lDyvc9SoqOmnE3
GMAtFmWhH0fG8WZ1exLr796KhHNxJYIJTdlvtfqLNwW+RCZQMMt7uFiOzkFjjWEl
40nniWDyvOTmA9a2p+p/WDWEMB8KKhe78DydXFJigjuyPkO9V8/OlSs/dCLKga+9
WeLxJZmu6TL/N2wd9a0DVvn7EnovU0sraXcpdQJA+iIG5zar9ANm8WkaeD6Crz9u
X9y3BttN96S4EdFzLUXKS02odjzt19aP5viNE6ij1Kds4qFs48BIN1rQAiR04dXQ
sBmGHe2sACqhrF5J6OAZnT+etFqZu+riX1hYS5/VfB5zP0uBBeUurW2Uzxwxg06E
FHvB/zRqgboqJixjOE9mq5vr7ALYH4GezrsTD2xvyA12flkzlGCUMpXZQZEhxNbH
xgfQ1vLDP0deM38J55MXWP1LDniPSyz7ChnVa6TtWEcUkhrwSuNoIuHlc0QuuOSa
M3isSotXzmxo/2AtUVNVu8REBgOLP7lY8UENu98RGt/7lrBMrSBiGBV7OYXsWU4D
CzWOaxMgN7U9t6NBMm0M9Ztvs4FAtJ43KjPKy8RhF/EEFyjucG4lvrNhphVFr2Ev
XDBm2jsWsVpJwBwNpE0hncC2gJVbETvuUhafvlnGaOrxGjEYsPecO37KXp0H3qsa
R995je0/74uXEehpplMh7odVVluzWbMKa8Z/hS0/oSnyOjbsNN+eHUW6Jzc673Nn
bDWlg6kUytqyw8AtpaT6KPKn25aJiFZaIL8SVmOQi8vrHrr4EudOQyuyTrqmXeml
ARmYiAKw7/P33zZFiLuOQLJudKXpiLNxqY1kd7n2vv0joIu0/4bNLVmf2NOHOQDx
sl23jGBjmOV3RnFxWEoPEehub3wKjHVSz9w1xxD28CV4Vd7ahy3KQZ6ioJ/2zm2D
lV1NBMMGRI0/JOMH+B/9pAo0CVKfoh4+EPyUF9kJdpurTgu/T1zEq4hRe2hZFa5K
Vg922Y04rSptlExzsmhjcrg/8Rc3hC1zPrVMZrSGVIj561G5i1HN6XNLYDXgN+9p
mOxscqNbHy+cB1rdR4G9ZpkZQt1HOm3nR9mDxiOrk7ZI0CA9hvQGr19qXqTs1r48
xp00ICteRBaPD9YQGb5LpnaaEHp4+s0OrwgK82HukQoRPATN0wyMyd/Z25YplP9L
RpxSnsecSNyKmxN2ALyBUZXLrvR1yz3z1NwAVOKvjFfjWolifVHkYzbJACO1xI7T
UCRFjsYFO5ZL6lNtM1zoQtdLogGW/IJz51Sm+fnmoU733lqddpAipCilNrLqIkYJ
59n8+xXWdi8Yc/xtIU1ndjhxXK0bHZc9YlScqhdRtjQm/D1zJQq2wsZjhd8+TcPh
DLvWewCsbpVTFWgCW0YQXfVzBfLIFA5b+Y5Jj1cUbIpAeSq07ol2BXRD66Hne5kW
HZuRREm38DjYEpm3JGbYrSHVl4Hn8d/ZlF+Gedd9lF8iXY1S74Y4q4JWxp07Fb2b
6QqnVDnP4HmSb1cmeYybbGi7bkF5MzbIZ+3a3F9ZrdNxb6rkEzQwteUwznRR0slA
oi5YHJfKkOwzSJQTEcniqL7c6irBsn+OBdOr7rc8JbnZE2mvR37XG02VVzKNm5E/
SVgCPEsAnncLKdogzlWBw5sbsrMJeEQlN8/GxEWOS4WXnF/bz9gt6A2z0e4SofXC
sUnFNOkfrX0tjyOgj/lYELUcqSJ1pTuT3l2OQqou189X5QQ0pk1JlhXAavbzEoCb
4Fy7DpOvmW4fgJn4FHJmvpC+xDdWFFOe3oAq48Uru6XLUEirGmIBo7Zk1PLA4wCg
Os2CSaAH/W611c2jaM4y85NNKOu8qVC13VV3be2Ks7PTfxRMEI8IoNf/gIbar23+
9t3zHBIbTJO2Ur0y4YisL0tq9Nd4Y/muLDGsdkK/wTyH72rxgxnZdC4XgNCs9GCN
5xbbSvE2CRYJm4otJKQm1eTlAHeF2V0BhklthUfR404gggcD/f9WEHYeLcvJfYbF
lYpe26trXmpJhR/c5U9LR2wdeL5n7bBrsXf09spX0Gp7I2awgK+ccWmlkFVNgKry
tUQp8XdsJiK1PTELOBkKuJCc72lG14SlI2YtM+b07Q/dDtDNM4CUfGBrApJEZj9S
uWCEhlQwRIymVqqTvQ8r6RHQC7lXCy4i53ivXmFkzx/bR4VM8+yVYXKpNs4VYBS0
z/GF4qCsPmDaDxDZ7V0IjPSG0EqI2Eab0NlCMqDtmxry+6kJxvHJyKFMhrhYjDRx
v8NOaB7OlIb5kJfldxoEfwNfJpN51xGf80MvRAGjt151EYuShnq4TCQr9I02znrf
wB4EN6ZgsoN/yR1mMld5ts9geSBHV0YVMe18ht+Jc9NONyzGqMZBj54gmKBnpkVb
fbm4eCLfJu14o3SG6W9igjolhNOQbn0pH2DN4P5OVdBQTaGHfEwKhlw4BZkK8SlQ
Mvx9zszhTAa/5GlZG6gZd0Ajx8fDcLvWL2ydxO9icFOeUeNJ9txUgu4PQrEXyK4L
yRP627JwR8QGieswXfsQsJPOptZ3OoEgxiSjZMInbOIY8Z7H8FG2I7A9F8HRz0f1
YPrSreq1H/mnhtiWSyraLD8pHRqfyCdV7Ih5y3EWocDkI3ru7argDFIWzvLsexti
lI85PF/NYsx8qSy7cMHiECMqiawXaNM/Xb/ecCkpPg9O0acqZX5RdjMchvs8cEH5
gjvyAEidmD1IBx3Luo1eMoYiNJPfThIKKrDKcKfx8GiL6UBMkDdW2oQovCSJBY16
FWT3JiKVzs1EHZnp1OYa3iGh6segLoPEpEE4yA9g2V8IXeQwsBXpj7rx3lwr1JTA
V/nbrXv8u1w/YBT35/twrK/9WATRjB9vd0Tg/phcL2uu8jY/M58MhQYPNhY7Tdnb
qRDqPIVpEDufcgLmduzz4667APag7HmtR8ooGf+bfZBu/X1mBfWwZxhR/kYILs1E
OtgspZTXu+F1bPURH8PKnGXYrxG01BbTIcXlynvIZiy6ngbeR400ywIn9pJCEyca
QXKKMrTBzO5aQ2T5ffhwhVMv5mP3kq+3S3Sjl6NdHRGYfSNdlVhAm0gEaDhW5BPv
2ML5bWLwdig+nvxCq14oJ88lwJJEAHmDI6b5PCuth2uSHJcNMJ7JIxt5nfORjXcn
EhONwGyyzSp11xkROnbqCAIlJe71APjIZxJu7zva5mOJ/65Zao6RV/jI7myyfGLk
0wCBY2yj7buEOb+5264MKswGKnvBeO6G8BzbIsM/YW/LMS5ZKE5inrMdXmit8aq7
T7nhgHyUvHf/ur+pAdT3dIbjiG6+q6DJiCDo+5QPdAG0FEf6PrQ9Fo5e+AIknj11
wCGFVab1UQUo9+82OeqKkjgB0xVyo8vmh11uqx2UBnsGIt6hIi+psvG+kNIepVSQ
1GjN1vlJXu5cq0XKFqC0TIeqDeGJsmb8Bk6m99D2gg+JovJtRdMiemSKosPyZPvE
EnOL4LsjNr5B5+2YF0YSVX4Wero5AyWZiZe2VZxBLlGOyq380cNbD3S94ZZ2OowG
lv6GZ7CHIt31CUrC/hNspp5Ik2huS2tphRgiFNbIB2gpk7X8BI7kITghxb6Y/SmO
JbMtjI3LJTDPVDDwu1s0shOXZ5p3fXD+A6xm0fK/rCZHELB29oBBU0S32lUVrpUh
almIHmcDfJopf6fKPH/VmFUTIC+m1X/JcEJH7hh7EXWx3QXp1A9f92PT6ZnaXhvG
xGz+mzBlARF5ve9QVrt7FAAhHdRPRTgvf/SaATWQU+rKNFifoDfyDwmEXbxsISv9
YF3h7lz54a2XZlUyBnZ+30rZuMtFyiUcW2WXZ50dM95jHY3q6QVxgoIosqzZNZk0
vR9/wF9Nml13WxKb2tA6C/QbLXdi8vrGpRdNkfHaKg7uUMTzkqQ1ql3UW5gKQcc6
XkpeZPP2kA/fpDxa0y6wBzZsZMi9ChC9meXE7zH5zRhQTumOjIqPjX3/AENh7F9s
o1NEFu+QXiKXMMhu/D0/vmwo2P5d/XNX4SSH3HXVeRauQy3pWCXAt/8vEMOIOZtO
lya0Pca/bdWhwLGM2DTbKBfZV/XB4S3HKVyCBmRSUSTiLiPFQ06GaBANEEEnZp1+
UePFdiAW2Ut33zqWELtUvcJFgy2kkfWlaUm2IgwsRbDv13BYcYhBUClIqQ9ptkUz
em4eMSiI0vnYsCLV/yBwC1TZL/bhzYew7kvQnGdz7qNOIDg1mSkcOD/gpl9/30Lg
mElQFzu5RH6hHsCswzSPUqbkqoOwU2tyYEpVUpjjGJEOZcd1C67KEQYFVoASRxEA
AiRLJM990OH61SagHzKv/mKYSl7PUIFipAFAvCxCYu5ZsiA53jSjJkr3xs1LnafN
F8V7TGw3l8I2aFKorzR2/+387Aff4uIWoTJLfhyWaum7lyF0waPv25tF1Mejehcv
4iMqCpVVDsn7YBbFSnzmUBtWoX2NF7z5cdvY6ZCl9I4tP+NBZIE/g9prc7ffedIb
lSk7ERs4UDtosdHj2fMczPOh2Y41WOVA7SsJ883CgZZ9PW25WnyEwb0PEwHCwAaA
6f11VwSRiMePEfF1XtlFhLaJ2q3kOI34iyEjqkiRPZviRIDLQbMi4cwknMR0LuwE
Zy6CVBRBoCC45h1pvuV4Xu8U9DAjIN5MId3S7lirJiMprUIWiQOcZftAgWFOZB6q
R4/o/v3s+AA3lDqxgtoO15IX5Ckhn4tbOItljjpL0p8oK3iNb0wZm/Jhr5ZjdjxJ
VLRutTZ4TWCinwg/R2YJYQEOYgZyAl9pyfSD2oZ+ouaLdf2HWNwUlRC0uoqWGACW
LXjNNEdnGGNEX1UBseuQV/Bpm4KClGQaEVZoZS/85d9V4ue6DpgcayebmObz0ydR
0SCts47rPB1N49+dZW36AOExHFUfyrIrIfApOCjQAn7/UcforsdXBx5sT3BIaKCz
V9HDkFqRmdt5Mq+5kjnUiOCeizQTd8HHHMnhSL5dtQ7wCt7kzhlllXDgpPVjKmCw
Ya5HC+EMUUqIf8GSjbajNIYRY+EJnVGsR1kUuEcy7U8t7YKF+Pz65YAe2IWxWe6U
if7ZJhrJk8/I8N374i7W7rxrPxQbt/9X5HFChxb7RdxHCbfX7CkagXV7JXfJda3G
eMVEzUx30nkwKJy2JL6Ho9247dyjbjB5hCIS/0+WtZLf3EghnstsZSDvOzojRO3n
3nNnmYZddFoYmBzCl0QAyPi00nY/St/B8XjFDZgHa7+4kCcDm3Q6Mrc/6G05fhi/
G2Sqy+uKPH0h1v1aAAjioiQhsmGZ5colDTOfAMgFlDQcrqgPv+0wwhN1cAHud6rZ
tnUKL9bKpFTLlYff3pLr21UpzdgKuDKMiGzyNi2OZZVLc4rGcJCB5E0t3BQQ4luh
gqPgIsFzOfHdtJ3pgdTPeTPBpWTuh2QxoPGT9EaK2LVEaB0THNmQquOMXLknzveI
gHpjZgAjqksH7c0VEDAS6c+Wpm7b4NHgrtZZ390U197iNaeVP0RXwWjbzJVyf8Dv
t1X2IYEX/XN7XildIdUKjNqa80FqUuGvf5cpjEqOVG9nRbtZpyyMcUzQwrd8bYbi
m2Icbjgvjz12s9Jpy05wSBgutsUohTquVlG3D0XGjNlz/kpVcjzZe8nJ+yQRDZb2
6k8c88HrC3sda5NLMxQWi0zIFgV+eYBPg0O1MWOacam6H2Xucq5AhwgVhOMZ4Vp0
osrMpE04xgbMD02IU9tWdacHY21NE8VZRY4llv50jFhrT0S1nbWcnzCY++FZ9ZEW
Lxqlu+U4bgp6GxfDt6FSuAAGG0emE7qToaQBQqBbIVhelViVNWooskX5frdLt1Km
Vp+tsz5n8F5dJURLHp0V0Z8ScnWq/dlFLTIQxQkBOZSfwpMqmoN+d/7RhyKz46lp
bE/fwcANxxpIP7K8Cs3dv22Xr0g4p/NClcAyZTEJrMcK1nZzuzZqZguolUu1FvwL
8VjDfa9U/i7Wd5ArjiBKRaY11cCJsDVzVWOOymyOcz4kcwAsVwfKjK7zOLZ/yGvl
XuW98sAjuiJWJgBM6bT6HuacWFcgrMK4G6cyLXE+tULhOoWOViOzsPUiu9+jASHH
TTmYAiU+BmXf2RhxN/xb5n40/hexs3tobU1SrJ8LKAD0yox53mVqjYlauh2p4LR1
+LLQb0+hoBDypVr+OienDXcKN8CJd6BVngJSNHvfx9nKF67bAzCf/HmL3bELIDuD
cmuSihqU52O0RwzRBrT1TvMOLNI4ux5X1uIHu03Fwqh1qU3RdLYo+jKPd8XICWKG
U7OKvCl3VtvigM6vWx7Bs5wNoy70zbkK6ix1CjOYVHrrGAohAs3x95BRxSHVcpHu
eJEqSlUzCs5fnLfX7XEHsZv0sIhX9cOD3rsw56xnIz1EqRlGVZggvLizSTcbubOP
RalebXvompky41ErZ07vo+wIQlZbbmHpnH770hdXZnjSPLx//ibUI+82pV8VOaz4
S1phxGtOlQn4BM0ZpfMZy+iCbkIMUTf7qva+cuCIIcHIyBRfWQBwHQ1ntXZzrylv
x7iGzZbnS63ARpFrUFsjz/Tg/Nz6e3fs1UW/vuKbyGWAMiBTVZZ6TCotZ3JlE5NI
zcO3Ok3KlAl+CSJCLQZe8xZmv5/B/Ryb5MsnRB+eV5/2Q1V0Firsq11696fcYA3q
/GEaeQmxXGb3FSmQwlfh5tDVRpbzauqSjNzZb87SeHqGag1AEZ/XlTgCOMZp1GBh
pRfXNY2/WkJyJcNCA3JN6yzofgPO1wBR36fbPBNmeKvQlnqG9qJVNe6b0Sm+vhg8
h5O1gy8TFVLVHh2wxyn3yVYnbI9tWUwQJMglPcyhz03BWf9F2p6I3NGGFP2M3Mql
8EyeSe6sVptA9dSHfKkuxcuMV0yl8df964KxJSXBbmlOqAnfxyBqgoCylXNQpq/t
XlC+mmb53jrycaGvCDKR0Ulmo9hMxIZ22ysbFXAAQCtqu51j2x5jIx3+WxYilW0Q
N3gFh9vIdEuauhPZx2z1GRL0HCq+agdq7POl1/zFVYH1IV2Dmk4qRLL33uLcSYpc
vPb65KGgA6Vro350g3+AM/vb3EmdpSudqGcUtswkCUHiCeiDi1Suit90/I4yJ/K7
syCDAtlof1c2NRHReVXV5tLZ1xTNP9FaQ7fjuSbNI/ifB+gIMF07nqk2fQPjSxsM
VPpcozWam/WMnObtKzDFnYdQF2ttK0rtMoaxpktT6QhG/XhZoUeUCdvAiYhZ73mh
qRmD2MAua8afnIZ8BEpeB2+wqU/bfSKKoG/0F238e4xQlrIAP48aXq32Ja00ro33
35yK2Yp1i/R255yxzgTeS/QsAr1koSsLLwaCiJChachHE48j5z5ZfoANHPBSP5dU
fvcRWxHAHPWuJ1hLOZldMw2T8QMen9PaGPwBqWemwDVcCZAT8FpUYgbxLmqdToeb
dp25TOY9LmIHMKFFPhSEhRwFtnr4purtna1eA/5wPn02BDS4mCBgFL/uuWTjGu7E
nb2NHuQW/0wpMgwyz4ozvipK5xGXf5qDJBHlmuxuTEA0Uzz3DpqMdRufJA2+jMCT
UXXbokKvOtT1bIIv6K4schld+0NbnQ6wVlOnZ6d0sMI4e0O6Q1dQPUgHTpZyisXo
uIOA1sVTyVWzADO2LKX0N+dzY2xR6mEQc6HWIBxhl/CG9YMfwFft/aW+xjYHEi+1
LMspzy+SqYn2pQCV9v9BafWslfoNnInaaMoaKCRP/S6IZy+3cyWu7pv2ujMhSq8C
fZXHbAcJGBVIpGTxkumjRavHWET09ggvxxYZkjEH7fbKCKElxVOz1TvS1u4nIxFn
Rw/rLWDY9KCgXleu9/BrNzsXSN4Jq30s3xmLIt0e/TPJE0LofASHfCHQDrTTMm9N
/I4TL0O97GT/DaUF3HF9SNP036nisD/ypS5nvWD+sP4nwkjM+5Q+rCfUWXsMSGSE
pKUpuex+r0NsOMzzpmjudmDsC/Br3GX3t0+/OwzmIJCYTMgwGc/tXj71JoGh7Qmq
K1Z7C7k3u2FAzvg1c5CVaXhoZUwHyz/MWgNh6iPdsioEZCFfdx04AhxFDC4OAUGX
WdoqCH+JrtFbzMrpXNjk9mtRKc6loqvBufuTPyIEsJhQsfuxFZ4PGHcbcgUucTNR
jX1ngGz3M2R+cabIIC0NZ9KBqxhEXYTnAQ1xffuJvyrXKqqmhBP5ey98SHEVKRdr
WUMzy/Qv9TqaNJxtPT6QS2iFxlZSkSm012BkMzVuJn+/bwjuEtGm5FybBFFZjUgo
rcCpprshXHYFbxMjPNxflD7BkrLjbl/FzQu4DVxLT/ane3FAZqtC/r4GyN1k0ymB
QP3pHFnDLy2zOopqr+mYMEG48fNjq/a3Cw4i0Uvn2Osic4lEE2523yhAJ8sDes1k
7w1w7H10mUDyDnxDIxulFUiRdaXGkEprIUr3B4fsDo28nmGyYl1vjy/A6+h/9tad
yOKv2R/eBuP9ZfyzXr4oqxMAFI056xwRHdrry80w755gu5KzHfg+80kLwKZYlj2J
XSWCUIJGLs/Fy+x9ifwOgCU+tbvr/TWXKLF0QsAWbFE7Mvkdl08Yw/OhDWQ34RCQ
c2nEohwhQ/cR4oreeooYvODumKNNu4c2u7DiK9wt9a5I3pwxlXo3VvAXxToNg1Ar
Sawx02q/mCuRVPk4q7WiqposVAs57lVCBgC4azcNKT08D5+BP36pGmVIuT4Ywv3s
t1MOeutXkyY592xvTBDXxrMbHsRPsxgBAcJufm6owWplU3ZTdSmy5nTkdsaQBEBW
KKB7NWMRNGaLUtL3VUaErjdgaFAM9NCjEE9GXJ20v/hGojwiXbMUqpt/PbdkzdkP
lbfYP2kapcQHIK0+WgGkyqrcguEGHa8Z0B3EulTbcP+mOX9xvfo4OHRvv3zPIGFy
FyPgmvK5QkZJqXX4Yi4m7/+0/WCitpZ63UrmbEJ2hRZSYJcccHSrrcW/2+tKGw1A
xiS/6zTW3/twTe1qHdanmsWilv3katmnDCnLStvt8S9/oNwqa14XO8pUgagA45GF
3Qx59xHWVGgzBe9DE+SLGx9AoCX+lzcBDFlaDldIMpUbuXsh5+z8hTIw0PnGbAIH
rG4YaJhZAdxjQEW+UB+2Kfhz9nM3LTCRhRrOQxPZFoFpCCAi3BNhPgSZNqnDTKJ0
T+TZjj/AM8Rncf7PwAAA8ZdwNFEFSiW75rf+sXWwvV8XLDHm/wVB1v1HOOBq2iZ/
4RI0a0jeliVX2OyVW9CwUjIpQUwZLEhUYVi1zFpT6a4QBIGcZJwah2akWOAfxUuf
oQSwgIM1KBKhYEv5NO8eMlh96PunF1EhNlKuTSjjI0tTxl5dBJu/Ida9cRsg+9KO
1PDZa8hUZ7/ZvJYtdpdX5n5rlQSX85uoKB+dKqg4gmi6iqPOlk29hUDQgvr2K0jc
5NgOjkvsLVrraotef9QfXn/dUCemmISqTxtgZFpfw/AbrUjCF+7MoZLO4c1dY6v4
MGO/ICA2k9ZrW6eHMroxMs19PiOhCH7JFgF2LSv7fM0vbIKoBMMn+6D5F33UQz2I
B7LlWq1Byo2zig/j8IGXauNSZJ7hO+SI3XClr3fzq3O6h3piQZeJ2I4KByUpo9bZ
uTCiwHqlXyMGigNRbqRDuuMvetEaAeB5jX9oZJPmjvVlxWTDKMif2WIsdTfEai7f
RE3NVjU41jSnJKRfnoADFaKENl688kJ0OAG54Q+EGdFYn7RG1WqsTzmB5YzRW5Nm
FC9AUK7HuiFS1v2lYVvZyv9zvxS7H2mUxT5sYcmdbbzv3lkb+S1Cq40XGaPHRIQY
BSpMsmpnB019PQv6KCqjAJpLeMejpedIjdXcYijemaQzO44sECz/+t5DVPKYSf6G
fECOFdSVuP3fxikrEToPk+AUpuJAAdpUdbAKSYBMuqufIMzzXwZubrHgYOLz+SIG
4HiBbq1JB8nKq1QvF8KlY4i2JVP0zNM2Xe/V6h1xVJ468a+jFUnIH3luDT5WamhJ
OM62sp4WZydfom0pnUYGpSl+dIT3p1L/nayDAVISBH8gOs6yDmk42yMNzXZcQVPG
1+hY6G94XpqkjhaPQj25DISM2wkSNUNDZ+kl6aLGXIZlOaRxDlKRYDWEHlH7Ijb4
jowuWx3v16tKg48iQRstL1NijRO8dOkpc2sgwJX9nguV/GFKY7Iwi9i+nhTv6DNc
QvTE/J/2M0pHX+rUovBP5VO6ZirpWOZLeZnEyCG4A5lcuUMnQdWib7pGWcZErV4a
vt6iZrQKr6DHI/CZEguqafAN2C5ODZTRKHy2ISYWs7Vxl9cZl+tpaAlwZJgZttTj
G5dvjW5TsbN91ov91vHgI1fAZ+HmW9Qhh7Ck/3WulpnC4sDhF5pXCdtjTiS+yHjw
A1ApC76DM95+lSP0V3zRM5CtpM53P9h13hmvR+ofO9HgwrZUuNWhkEGUbCj9/hXo
0jOD3mTVJ3s5lJZnrY0CMewXCImAaLxoSzxPs8rXwDRPdQpSdz/A/u4eXE7L1pPv
iHbmpp4SoF87MJA2O/B7faYwWVGk4jYGQE7RqxxKgXTb57SceQKIINwc3tEF0pGL
Igt16TY5ND8FibjMELhLAOojUd/cWanIVupwZoL5morNc7zQ9FrpTAv46lwi+TMJ
9Xlxi6T2+gY6qSkCzyTnLRkJzFaTrgdHn7qEEAoEtQ71ajRYZdPbhKXxN6s2OVt5
Cx2lgn8xANNSfEyQSZxU+LzmdDCLD+U6mfta1DVgyHvjA+XskLsL4lV/kpZCI2LP
GvlXnzqvK1lnfEWR+4CGfyHbuGA6oLTWYs/eg4M8NxyV5Usix6xz69CyYWJxkSyq
xYZ1MbVzD7JLydOohlaGqLWkeH4kVTxefWbm1KXtbfTdP1mqAd7Q1DUX1GCiu1uF
1Ho5KQsEWqt9X8lyt3rgkvo1MVjuZY6IqxZ00Iq1+VRZPI0ffUsQ5L4gWxEoHiFZ
7yL4Kk2PUW6V/K+nNNX8Oc3e7Z84H1HxHiS+3MbnnHET4dnw1/hqvtt+NKnVDBRB
D8ZbBgRmZNO/oj4MS/SVHy+CDAmg6qV+AV8WQnqT/Rgu5DQ0a6cI/WZaCAPJfBdP
6GbmS1ALFqJ+1Q01S1VNMItJYAL5pBp41HS0oy+EOUf6Ze5GYS68uA7UNmf6gBm/
owT8BH3pGMxYgZkY93/pu5s3c7TSrVOtih9g2edTeUXVcbrEWtR/JeRdVTdVpOy6
F33XRJrPB+7vGPnxk6d8s4PGouihBpJfrnFwgQR3M1aTbhfUHx16SFPwDgf5ooYh
33miNxuK6yJ6gd/AbLQiNETD7cncIEsVSptIBcye2+gkSaQ937uABCsPxflEhbav
LKMBWVsjkGmy8/yrFzGiZDQ8M8nYvf8Ds29xWH5uwBfhwemSWX0MJNVo/st9kmK0
BnnS8oU/w9bwpGmugRdBzv6yLAULjtLZO24ZgXJxuVDTnw+PG5eJDJZVSTwS598E
BhgoIWLid0GDOIMfX12pjuGy1ND2GThbSDy4+ZQZV6whz4bZFp5gU9NZtZX3XT3E
MwIMKPiPOXlvG+d7CYgo7H5/aprSshhmkOWyeBRzFqQa/EKdakBT9HMRgii78EcT
tdyG9yHpJkU4+KAHidFCP2quIiRc+0ohclaMFgK6iZnqP8p67QVWb834Q1oSWIPg
pdfSaHeWQ/E+PBoBjs0ETcM7dKwzmvJZz6gNK293H25pDRjFguPKR5qkyrOfHQCv
0b1WWTfi4eaKZkOUg5VZboMufEAtqm+08Eezf6G036h4GW6Ha/HicKB9T8eAMAWV
vDvYUPGQ9Ii4/kR0rvoFIeH4T8i99N3DnCciPotUzHOKNuMm+qakoKm4i3tJoiN4
3x1zcGVGRPcgONBfTj/fmXFAXCq6JVcjdLHR0+HxgkA+ScyYA6W81dpaOQQEq7WW
YSptWTd1vaUZLe2AINBYES3K4QT8t0Q6vtKB07Tc6Nv7OZvJ90h0R5AcfCHffZA8
u7tdZy8M0r8Qxs+kHg1YynSLlccGFL+7rJ2hSPrj6a5Lx4XPepCH1WIiAe3ChFrZ
gVmllFXBCO2MD7mGP1GNLKvEGUzEZE8WbGXBbGRMVK+T104e3Uhxe4aVBRVl4x4a
V15RCciuw5opAlvwAfA4PLEags4D44TG3H0LnIiEnLD1ppXWk7ZhxHnXhvaIS9wO
IDpPwiXNdhsUO8jPrgJbqwz7mXvbSK3qQADI1+zmPruoL7UH9dFeBI/2tJIE+Kqq
82bqVQ+lMZ1M/zuohwhKspKizCkz/GeeUgMHZHu0fuAuMry5urlvC/TuG55YSvf3
Wdz47NL7lU/O0rTKRxniZWAzXjE0v/g8LZhGB5tECB2OtyAaLw+1VNEke3JsDIiz
83FiMsyYNX1cSAdYlD3eI5ws4kEgaZAOslBCXhGieLlMW8sYybMu4CMEXryyjZeT
Rf/Ufv3fUGgJJC3QDvR1/toQAuCtml9MKZqJlM5C6oMQkzUe2kXW5SVqLG/qSpry
To5/OOr4SYP3Fmqv2rofN8QtV7SzTx96czg+cbZWs9Dq0nJ6kGY8O1i8G9OXRWg5
Le5Crxzh8hTfQb0yuE7adzoLbwwXuQfD9vZElF4qavZto8LJnVZ5m2n3PLY9UT5A
oglwMxxZ3yXRjsPZsj5XTuAde8FGJ/rsGODGomPBHbXIDD2N0t+R7HLF0nvHmeG9
P1GZC1Co7h7Mt2NXUBYafdGudahkNrzirP8RCG/2Pzroa69FdcAvFeot2L9fgofz
ZWjWi9QHE1s2Mx8nVdxysFFk+BXvyO2gCzZ7ClJjGUnEkHLrr04NRsP9I8rf1k8j
/vDkGbRKb3E5FarYxuhEGDv+vgF1aYwOaqq3AK+vdN1w8oDDyXFOzplq40286zXP
E9JohsXH5NlHsHiaEm1pTH3dBd492k4pGFSYP3HkwZF+rxf4AQYYIl+vZ88OGb/9
CYH98kHCrh/dv60Dwxq6lOEvqr1y2Ogy16D7K/vqrK6BK2TTS3UNHNTqBqcwCUki
1Bzz4VK0tw0FRJsmAiP79A8/a8gIstNXVpTDJW9Ei13ZTN41dJpVBnNKijvX4ktz
CCeKoT/uOBN5+kayXSPDzaPQgwtsD5fdCl3YtmqFvrivRbDeFFTYJDjlNAQ8iF24
jftAvGcfrc2FwzIjTeMuc2o8F6kjvUxMBBOxKt3D/bUbw6PPK+OujmutzX6dehSy
ITlaX2I9W6i7TW120uYR8EqB6d476Gy+7l1n8p5XTZZkLq6tGTfynuVjrRdBYGZy
i71nSJ++0v1urj6E8f9xs6RSCwiqdQZSRHzOALl8N8IVP2pFzYFxb5Dse+kytN+C
Qyr/ihJZyPWW525+qaYMMmt2YN1DuDHf9QHgQUFBLjjfFPfhlZbgDi2lAue605Aw
F6JrTXRg+P3Sr5hjLTFuo600/c2g4tg8Y8sPdrl93G9QIhU+aSq1N6Jum3aAqDjf
NGE7wU4LUjZk3R8TzCECVQNl5It+CIA4MbTgFiE3hbGB9qlAt4hMiBfIxhr21hys
knB+dawtSFA3n2Q/cY+YDuUJaRG1NV60M03p96hvtvcFzITEaJptsNXLnDP4gMGm
wI6PZNHYDbFofOTrvB+NtJezgriCwAfCmucsMZDbpWWqwd8CEihLjQDaTeaVeQel
iKmki4A3X1xq/ZH+PgvCP4bSup4JR6hGAX1dtyXAUyw0wHSK8FSqVDg22HAmcgHH
sbV6jVM1npJ3LwnskH5ZFwiXgc4L9bz3QSixprhrAfSAiQp1RFi9vVEg+olOytdf
waP2fWbwxV/sDey3adC3lt4/tLy0wzv8fkSJyr5xqTV35AUZ9jWjD1rKd/Xch9L5
O9XR+p3WckihU0Uw/VhDIJEf2MVQGSOM+CYTslu5iIZ+XcGKXiAL1LDoy+NPuxi6
PwlYtvj4le1vpvgG4VQRNc2GrrxDWhUSFucAvcsuHPRHlZmUibmjZDbklU6Nfkah
JkZGxHMZr6L9SJpHkyWmzkHmc/EsJ15+/jc9W8lwzt67GhINxycbwkEerzQttmgR
ai7sqjdTg29LS6Ztkf9txU23rdrWDLUkLJOvCv5eRsXAyARMqSiSeb7aBLPIa7vm
jZvj+nIESP35ttsVi4s9usBXcwxot974tLgP8ZOKYpuCq7ZBSDlvbVexda9T5CIO
5a2cnkRYrSkFR4M8zUS8S/cO3vjZVEwAAUPSUiBx+okwL4VYSpkXxIWo8m7DAtyS
3bwWosUTrBbRyNX6tW8cXUx/hDiRnWrjixjevt9vmEFC3bxXzqeTmnF/AtjlgHpx
oqIcckimBufycfRLI26/Ofsor4s0fy8fvgOyO408B6m8itmk5DnGnWfg5f1cepWr
fermFQQYEucU4xOvDM/o7Pqx0H58CntT3dCtIwTLDdo+dDy5Bwo4/Y05KcDhmvSe
9WXzGVBf7jxCatopFn9LA+5ilit4fq35Kk80QO4Occ5PuV2iTRegDUnbHaFmt5a6
tsvwWgd5YSRhps5tt+0rES33pS85HDFMQBtN8fTM4jpxEEDtb6Ca/iwiXvCIKxIS
jcZn1SyY663+eMJ7H379/boahFWC85ir48STQWvA8uDV0FgEZi3SaQuw5ku2c1+4
GIJYXZdsTGRzXGXvZkUF6CEat3FimhLI+qkYrMvpctMtl6VCdb/JjR6ZJo/iZCo+
PL3JhUikCIG1OMliPiTLAnE+BOvqy7tBiIEvspna1qOkvFvyV3ubiqPzAuJ7KTUe
kXNCMuyLq+VzKBzx7XQF+HdHHlZP2Mi7kmypUfXl+kXcIKJKsYLISdrwhUIN3jJv
pA0ymhjZz0PljPg3JUFdTsNMvd+KDgtXqpoh0lkbckpWBUIGf+rjogu/ZnK//LAF
W62bX9fHWIcTIoAbu670E/S4uziXqA+zsDnEJ1cgFkEU/R2ddCvwl08P3lnwi3B0
b7O3MH55T9Q+w0E38NgA4tOuL13FV+s08zyFBchRXpjGa3p5qWCCe/WQJDNIU8qz
R1VLdqH7bndq0GZrSABMrldZU7R8kkc/38gfbuaz92k4LDqaACv3NXfFcPDnyNJD
tq1CnJKQfpx90W0i0/TGxaxS+ohZ+izvHJ7Yo/kxxJ6QeF3auUQPVINdK0jINsg6
9ewEm+6RE/a0wsyc3sm6gglZIeY0sKi3AlC02DhJiZe61sEiaJ6h8DC+P/8mSB+s
c+CrJ2nhfYsO77M1he1DTdNU1OKnb64y2XBVaSIzOjR81qMGjB8YSfyd+ezmkLcm
rHsu4YjL8dJYNpkiMZby3omoqGp5D13zq1n5ldPZJv1ide8Ec0K30F3lrHqowPUg
AsEqOEolu2T+mqcPEA1yhBHzYJj2iFgbjeRl05XDrGNPVyJdZ5QYigsNTiNK5/Ai
BGJRYsH/rcp778oo2EGljIdZQthXD7A++MVo1Z3KPsr9ieDxYqnYv4sPbhM7R8tP
JrtjmE1nNfvKzgEIrnTS7GXKHGV5pNddHiF6dyPMXnIPi7lB9VWqv+rp4imh8v8b
l4bgCaiw/+WxrAawd9jE0YehGi8Q+Yiu8JI9zb/+0PwAHMSpvSrXm6ABc+y+pDS0
ofuNdp+AgQpk3pECoLpDbshhBtciivf6QXvf1/tKPexL+Phr1G8ecCdDwJa2G9oC
jz7Z9v6LGUzcs6klAK13Eli1sBhj/aP6J2stvb97t6s7MmGD6QuW13Ok8xDuGuz+
yqG1/sq6K/aR4UQoAUlHVajKv26ryUD5Iz06wR42CoXsGPHN/VdL4LiwIOuh/H+l
vABoXGSb8NUfwGEty8rUZRbkWeVrg1LY1zpKAaq0jw6vBsfkAve9XL7SeIDS0Lb6
n37iLaIsKt0lsUZ2Esmbd9mBfWbAchdIWFj2RdzZ/pg5RbMQtjdHmyl1C9kbthuu
mIMenWs83CUeHFvkom/GcGcDXQu20cS1vt24p9WTmOuoulNDX5CkQyFG+O3KHciu
eTsJlPr9LttQY3W7fRKzVEwgV3rb0q0OHRdb/a7sHLHKo4IhfDEgXpAXUzZTdx7f
zufe0eA/SIzCiV6De6GXEeihXgjoX6xmw2FjT518rRDPVGgB4xxibnCoY28d6Sm1
r3s2Ohi8jdj/6Pe2Zm3Fl2uKTclSaKOMyTVDaikBP8eRaLLlZI+h2lfLa2jlK8vt
gJyDncrLtRVrjkY//XLJqck+Of7bUHEUYTFkCo4f4KqgAz+UNur4OXB6S3LPGtPJ
nTmIriLVMnGcipPI7ix0m6TeP0lPbBTThKfAc9td2m5w5J47sys/Z8Spp0gTWprm
seaY4snOt95qPo8MPQJ3/F/X4DkQG4szvbKW52qxA4Fan+6B3gCaF9X23+Jrp1DB
3/xr3VsFh4sHhanCHvVT6neJimvmz+m4/xSO30fpw0FPYKX6aC6yBls7YjtX2s5i
wgN+I30wtZ+IuGMofaAXzN+/3rej9b8gJl9yzdza3y1dJlBrZumGRaHtbwX5F1Iz
AqPkcagGOuhg7Q2frPCdz+BJKg8/GuNL/ntEeViF28euAaqjoIYstK3DyrK7oRRi
N2ftEBn0ojfSFrKENMD5QfEhS5hFheRTj2qogJIWujicz1KDKbOPAiEt41n7MjWE
88YE1I/y4dwqZHEkJWdp3yg6n8LkOaAbJgpSiX78LGobxSQNiWeb/giVw4POUpdu
JVptSPiCkru9Bl9nYoUQO8BHEfnpvbCzztVIT1qp1225NlhuusQv9aNdZ1Ciy0rz
ixIQ4LJjie5d8cfbXL4ouvc82ddf/OutfHgigof4KP9AtZFtE12AOiBJa5PcJNoF
JXSeNbAjCMdI0XjniATAqa2IHDc0hmN4CNtkLRy+MX9WUXmNSMU/fjwKqIXFdB9D
dsePE2Sfin1xTAWSZSF34NBnrt5xQMepQzp4pQXCvkMrE4Dr7WbJK2MffI142iiO
JJ3U59SOdo6bsDSMTJpl0CBbf81Zlvys/88ymVzdlaI00MzdRP0MwzLuBCCoX7FI
8bukA0xhy7vmrCwm49xdGRDRZHJJjZx7fW+Bd/Ru+LA46KzCp8AvZYvBBBBEdps0
cm2JrUiPwcvzF+Av650xkCnX7GuvZuaQJVqssu1OIS61X07y5uzpQhsBWTXG7WKl
c9cql65lkMpETnq7y9P0d0XS9csglIqMhrSAQM0UoU1hcsQMtDj1OaYXj0BqDPuG
ITByIy8+dD1PjGPVF5ip5N4rjFMmQ3Woa6Y7aEAz+O4qUDm+wy+9isddg7IF2aAT
yqiZNbpozl9nqJLgsi6tcz/92LBN2GCMNT8ZIGBaduSpton7IQTQL2XaWYZF/5ID
vNv38gHDeL9OnLusifbzstIFRmnoI1yhepfFt4tEiiyazxSs4StRP+3/Hw3yoCcv
WMXyi/nm7D3LOceozVdZwHvAGOpM9Up5fddTqFgR3eyIlSbm/5oRWoGdsuOqAdws
kYxnESXNzA6QGt7uExdKyAZukOaf4J7nZVtibpjlgUXkxhHAAZlwDCkXOzHiIlyc
bZ2UQjmshavGnaFnZ/I20Do9n75O+2SCBgGxUN0atBAVcUKQANjwD8dwzs+ewWqy
SNbiCr82aPC63Lb0UkM71BucHczAGZz7txhCL9Ox/85DRLzCI22aXAERd6t4d6b8
x8ViFhAogkjhHBsLOUcJSsooDMfF4XKubb5yc8lMeeJJ7s6TlPj5U3bxTq5PPYC7
X3tYEyIzeh0YuqETbbXg7ZK08idfpBiwNqCSX+IO8OG/rZOJefjo4njzvoAtbS3w
M9zzJ1Y+oOfxkf62ySa2fS7Lc7La1d3gpIC1vPyXBSVbmIy3VHQ3RPta4OulT3ux
FWv5sGRSGUyJf+1VF0ES0KR1lqaWrfDn7P+8xXeVbV1/33g0yxH7ADcPo+vk/hxX
ff8iMuQ1XHugUOnv40OWrpQAz4IXfdwttZHJEfOCro4retf4TckMl58A3gkLSBtE
uveWOG3BY0UIdz0SGnDW+1UbcfxGTeQ+ibjXik7se1/oI4ou/Z3WLvAnesmgk31z
3TNLcosdwsT19NK8XW3f33YEgR/uDtWvxRwfb6rGRRSAxWrg6nD/BAABlHnVdFUZ
KJrZguYdKg3P4jd5U9MOg1WII3YXHl1c7F34twI6yfMPQxfXS2a67+sIbf4tNJQS
YoGt3axl/zyYmLz9JSLALKz/4l9z/xCW8EvUpIO4Wc0svrHCxKVo550jgU+yS0zL
YscnVEHmPGhcQwgycqDPBNdcEW66YMleOlWw9r1w59ZnZi47P+I1PreR4FNKT6oD
eUmiQ853BY+qDh2lVjx5vJPDBeoLZQRzbfrIkZpv0Ho9SPNKeGIaYfqW3GNxcdaV
F+yl++GIEOVIMMyYjgbR/FBox/PJbC49E+qkC5fFzl0ENEj15l/NSE2rnWyJP/cJ
CsStKeQERQJkhCESHrqKOy3paa8K7omMdQt+lO2pcwAbZ2Cioq4OW8KBoQM53txi
0ARdX0CKMEvV6Ypj3lCg6xAyfANMGb+hjJPAHGP48l03Uc8e1QXDyBcq3J1BZpfy
Zxtnn5kBl1h2GJh1BIKr7Lv2MFyARQ8IT/HQ3yUG4eRTIwL0vewzL43aLP+yHHPG
MjvShYK/leij0tXZf0EfiryGV9RtH3Z+Tn0p9U9rTmx+micmIMDqIKbnmOiCBnRe
dyOjba0eC0UkUEvBqTDnkQLRM76Lhun/1baa/P8Kpg9x4xQkN32ys+KVVykdHQdL
MDnZJXf+/UaHFaKgDvYigzaYs8mH/ApwrezQraMRkXnl+Me1L2bpWrxdLWwPupSV
7UbsAJXv+Ld/w18zbcT0a3gROybQW10XxWYWzFT2amMy4nzyejmlOmFcIhBVDfNN
EIIp5nYEgSKKkTNRdVqXGu3UqC0F8Fv2mLSAUxkuQUfQwUUT0yG67ikagv5tOLD3
vBdjuES+AGleRjWOIFNbZfcpYYLVmlHD0jMYC4MzWRXPF2j1IXH5FjwBolpqw2Yq
PGNOYG8CTP0pk1Gk1+jNF04WDK7FI8rcamUl3QQz17F8Fc5X2+imm4OM+r/eldZ6
AxLFyz0jQGGcnuUX8PKu85lVyZVi+RAT7PJB9TeWhURGfnNFsl2lsCEqQWLx9t26
q7yils2OK/YvZO2SX9yVItqIimyYb+bXV1LeihOOBAIJfbQ/39Zvr8kaLiJ198um
kPMKHRimhtQTOcg3DrY2sDKResPHkZerJd9C2N/17qki4TQvPgapPLYdXnj2mqC3
FClQWIffkfquRPeje51WUmQVCa7ElBQgt/ZaiA11cZF/XamcROn3W0OijBx/L6xU
HXB7x9FctqYTIBhlcpysBugJH5eDJS7ePdGX/0ge/CphTSxFbEacRwo6uhCRttg2
t2Rjql68na5YgPga2r5RKqDFz8mTFCO8c/HY3Rgh5oJc62A8yvQrXuxVnfiCQ60q
NRfgJNL+K2vLGXeOilc2T3m570PDp1vQUNXfBGNUsin4suAwtSHGcWNiHpvNaZBw
v8rh++XFVSGqgsCgo0lci8vkc6f+YqQ0k0oadT9vlZBM/SgwuqJ6Jn9NMTdo8rF8
Km/W7WzUomgklTVCzcYvBekb0WAsEU1vfbrL1Ucw/5EPQC/58Arue0I0mfU6lVwP
oJ28kAzS3rBKP0YFvexQ2B98vBcIVQHGpIxVzyI1MiPfmRAfqgAQDhFKecXmUXpQ
tjX4W5lgE6Q+qJ758zC4lgKE3VgXowht4cjEtoMBkuSmt7vCMOYWrfQwkJq0N267
k9y+oSFOUPthwy7RNqeQVVl4tzZOjJmd960tYsOySY1aBnoJvvERt2TKZSHSy51u
albvDPMZwI3jc9MvKATRi6SFunzw1piTO+9mn7ME7lI/wJk9qtQWb27WdMV2dsxs
q1QcDCkmpQCrGUh6U2cshbtUrza+g9rxBk3VuqrWRbd2V2Wo4GQh3/iqOMhUmw6C
e++XvfXI2yqn1we0p49pkbmcGK/CLnWXmqiF58slHKfqQCcY5ZIRZnySwhDKYiXc
ZEO+qosdYmeYnnu26Lg7wBSNcLbjyHNQH7vYYrGP46fQxADpKFVUnIk0TtNkLsLF
w5JoUJRuYjf9W5P1TrBU/+5/cLErtuRaAv0v63Jp14DoYxxhJgemK/3Ncl5bJxSG
0eUD6S7sYUAeTwNyPAytkszNeyHceKDFkteTvjE8EK+5oOSgxPAt/iqlj5WrQIM6
Tz3CLxywLfWxGufxP/pgzITEomd2aeDJngGeOX76oqQaNtbgRJEjBxmKr6XDaB67
bpcGMU0fhsN+GhOq+8W3wS57rnM4bIG8x0o61DuSXBYLSlyIZIChhciCEIGceLgj
+vxB7ikZY/g5FrxGLrXzox9dk8xMclcIUTHpPG0VyxJRCGFa3EjrPTcg+FMgAt2e
l34qY0tRPTsDAW4+vhWhpoHcIEqrB9rzXZjsHo8xsGs1vUEpetE9sjk0iBhAONh+
IEfSLrrcZXPW+KnZ3dqMMYV8/FYe1LSxTfiJPJ19GNCxOB3KUtd8K5PhAfh3uat/
umWYAQmorOUunoG9L7QS4/ty8u0HJw6sZiRn4LREDCPomuaLYG6+PpQp/WNmQEqy
4+PUINDhv4VnvmTw917maoZjDD9DuPWpJ5y0f9Rk9f6VUT4OfKd5U1A4oufWwCuA
hcdH5xUfoE0d1HJGwZC+GHxKkkSIt6tu06A44yvvu8cNT0IYRoG+gV5Gje90vijN
1gLGpySYkhhFrd5AaDPaGxJ1t9J6nn4KCs5XN2GnGjSU8jXvjD5GVePF+PocP2vw
LyH7mbSyOhLbHLpo5KdezyVOn8Yo/foPOO+taazzqP2K9oYLnepZtWkLT9XOE17M
uAEVEWsEZ7PTc9QCmNnfFikbTvou9y+ph24hHNJ3oBrrm+2vRqKtDSOuuyUk58Qn
joNm8HTltoZUtYHYwhVtxrf5PL0EPZJI+ai1TVQXO0rE3WRPGrZis4ZtOvUeQSqY
Ppj0uHeQI5H7ah79YMVcdYGhgZ71ombhApQBOf/wNyyo+G+BdR1R2DiuYbpgm84U
DN6mStKfRFT9WxA3XIrZtLvjB55ABnCYpyuDa8ITORSN5nffUfABVVmC+8NBql1H
w7L5/Ut+PXSqneLAg0nchviXQ0as/XIrGax6k3WZhCC2aiiU9WKbyotw8piCVkFb
1H1vS1W+rg7OmHZ4za/4qvm/LnsKDfO75RJ/UX35yE45oyRMhF/obof49kPgr6FA
aySq6iFEDPEJE9KWmCKpTL0c1y40YKazVuMlHtDnVhLdFBBsLjLlWsQxS0rWLQPj
O+VduH6pV662qIM4KGkeG/BJN9xBcuCaJpWrKqLuFfE66rYiBF7/uHgi6fxhbc/R
y7m5if7jXO1JWrB+cq6ZYrfgsC6eWn1WP9HWYZFsFRMZxqOz5rg+cQimOlWeGt9K
soaHlk9ey1f6c6CNn1XE9WxkuyMkJs2Dj0dRaVm+84UrsOtfbBS9gLRwKCzkJLGE
zBLkMF7suyaiBpGsRYVr80gYpLXzsCVmA7HqtPWDOqgEzEhJvjw4jEfseWI66zB3
Ry4p7fK96rjAmGcQQr6c1wVLvXgTCAFnFQXDMVjXkhMXgkGHdQFwnFcToxwGSjzp
A/XkbD0UnTjr+LTC7YP93+2nWnxzYMBLhtVnejMmv7s48gfBwJKyNCUc0YdlI1tv
71fN72N6Ij0bKEC9qLxfRGDBUX43v/lp8gbcOXdIuKKnKicUcKgDmjGoHJRs9H//
Ls12PyReaD3TWfx3EvPhPeVbHO7zRyty7N7ZuOi+5vledf/RyKDnGg/ZqQ3ad9pS
HGm9tt0wPPtN1Tt2SeWUz41ROr8Sz0V1g6hGehRxVDWYj0yc8b/jM5HgpTHwIMBR
PN/t+fteKtpiJJv5Je0ZXhlP7QxFg+dHWL3CeXCpVg5R/DeEwMsKS7bBu6pY26St
uID49w3NxMGFPLAm9tNU2/18B8hOEecI6Rpz6mggFuP/lBCNlNdNqkzoqgyEGiZG
rrs9DiAh5veBG+4sTagbBm/qAupJ5GjKmsDwPApDL8GSx3V8r/S7/u3F+CYwoAhC
cUXQrt2DyTnO998jFW9w/YJNvSQex/oQx0V+5md+4mvor33vW5hYKSL/0rgtODuD
KfGwlTtjQx3aNUhAoI8MbK1jHFcUXk6cjOdySNUSeJ0S1dR7UHLK6asL8/IEQzE/
IGGkAsbNrIovJ8t5pzNcMKNO6gCjxRz0m/rWOw6X6HX1pjspAeBQ4dc/SLRFF+Tf
Ju4t/+2s1FhXQm5ydEidEywy3Pqb3e9oHJzjfClokqgF9gjHWm6K2BMt5csCj/Fq
udMvlCb88LMRR5iFlLuZYINjHajggbPE2bvDs2Z1ysdLbhAKuOXZiqlxNcYsMTTN
RPPIfJEUq/3kEYY6wgKIXKFwR8MbHrki0sjooX4FiHAi7fV6wM/Hb+JX450CEbma
6B+eAdlN8wIquYrj1rQ0aqj7/qUVDig9SgElvmlWUY2Ay88KbWePFKigPF4tbnXr
SEpLhos2ckhUAyGeMcaUzSC7BjnEPfZk2rxL7LBAhStgNLTOOkexeERn4GRhSHMm
9NVM3hAeoAc4ieOl7vYVRmKyMpF8RFBc2sAuTnpUsgYx/q+UHOfyjrKyMIdgBtkT
W54fcGQ16/IGHrUQ7Df70WFxgbi7xOZ2ZkwK24lOmPXLJ80aqgcDhi1KLT8uZh1B
cDWqYd/MgjqNK5TYre+epSeeNF6r2JZotRnqPUBG9WaIiBfao1O0BZ9w1O5sGRHQ
laveC8algS2DeDJ27qFcwdRGSFIzGgOI74Cz2YjtNKCYrYj5imCvTe62XGRH1en4
M4mnC/XrIsyOVkeIw03cqmdqfFK8v7V8NyU9dz9b51ErJKzt4olwJApnWUA1tgC1
CrW02hOXe4nnG7YyekfYrjAs2PMTPE09pS2CTw81F5Hcfo8vPXuCzU6OZSwZUO9R
AUXRRuDr3qiW3U9tYEgHkwvE17wtv+IriOa9NLKu2jbaEMwSZSXkKjB67ZsSIYjP
QAhRtHIPp+/6fYcJ0iEuurcZUbXZ/s9HvYnnnCl2nmzxjC7AHXsjGNUnsLTgF1LB
8y+CRgI3sjAtGI2Xys0BSOuJFvKws8OdTOapcWgPAjFsIYwP4c2qRulRRT390832
onuS14GV0ftLBZXE+utQOSbWmUPgJqfbb323c4jt4rX05G6qJcwcGUX83Uxkikgv
KtmzeiqvgUq7YdTtHoh8oRaqTPOsZVOkL+B7PzNDlcruzDv9FMnqOGXjwZP7ODt4
wKD1SDTCrAOOVNofc/RBk5mZ+UXagfD8i5ta/PsaJ46ffFBW5nBXwiDlKEtsXCQz
adbL7l56sQkfaE643QBZJA7uKMIj84O7TQ7LjY5ikq5VQ64xchGMdgBp7hyqlQjX
OD716NC8k6coPhseS5nN/Mnzgw+wBbrIg8YmsvnGNF2ig7pJ0cceOiZFUWtBHLk2
AIWLSRht3qnWJsGbIOq+kvE6e86DWdGyXcD/alXm37yVaaov2jeMQOc/qzaQSgdT
0vVDoBeaPGHQPs5XTTb//VHAORUcbpvho9YEc66M7e7PPr4QO/p48jFAlF8xej28
ZM80ybe9zd3qgiFPDgXG8Sg4rypyurdDElznKDO4M52zc+nTDZQRHV718aCTwMr0
uSZrf4ShS/xWsaZRV+fFii2Rk9J4jMKtKhL9Ng+7c2M2TL/nFZvotqo6b+vYgTR5
nAKZEo4A2u35NOoZ7RgAPPvZw4rbPYfPqxcxC9EjVwFuWim2qguQ4UKBH+ifRd8q
kEUXdh1wMZNttqcDdnfIUw6kphSxiA5M4hOxAEfArET4ksF5Q6O8Vpd+E6SSUXX2
5v9Ga+Kw4Hs/uiGe+FQsuawT0cNwcbayPVC9obh9nAbpp0dAk1u537sTnahrHpUT
eAOYMIEf4QGTrzKmYU7Cd4mteK6JlT3r5GA3i8xM25GqpFNTfRBxH5QfKuGIWaju
8sjho/xnejlC2XOlfhD2RV5t6D8wJMmWnGrpD+/AuKRwu/odymPU7Z8rPDZ0x+5g
KaznbWfyyPKefN5svQW+B/+rIe7fdzTAKcM3lZt3EQUJnb4ajdBxZbY2btLd0O5t
/AAPdcYmwS6u1iWk/t1rYu6mZqCV0ySP9a8BqTHFGkGGKKH52lvfxNq/pQvpq4B8
+UXIESA0jxlTKnwkkU4mc3q3QPr7LYlze0Ny0UM57RyQHfBjhxOa1s3n6BZp33Bv
r5eVD+Ps0t+pGuj5ybBGt53LugNXBakoK38/uF+ER/L3UMdu0lDbvqC37+nPqOOP
n9cyJcqxVSjcA5AWS5kRrVsaWYEuxgnFVA6R7+wC61bYeuM/p45C1r19zE7xHWoz
oOA27klsmIMYO6GfyXFn5POZkjldtePo/datYZpiVFjKGw25L4qthklquF9ewTz3
c9UNIsR26wvtomr5M62wtvNFMS2kDQVY42eTz2BLy343Ii2EkJOAkW5lfMr0JAIl
lW6SMIcw2xBU8XFev9h6NJI/7ElS8KTdm+n3k1EDBy2NH2oA/YyY+f0ljZYb2j64
wZHQ7JGK3YYo1FrqEAlqBnwVQ44EE5ZfBoluvdgOAY59J5jbNVB0mUUacSdUyibh
sqoioKRd6RlINpikevBlsZ+ezb3IDwZb3azxB2J+GeRMiIROV07pLFOzrDGBX7mJ
qnaWuZkMBfLOjFq/G/SYeyQjuck23DpEr3sQ7qyWX6FjNB4K4+IlhbVwvUZ0SuA9
RxSYDmtOk6lhnUIfgcaJO/Fk3/eJop2+XDuUDfNuu0tGLLO7rDxv97EwVIMY19of
vcp0tgXKKdom1ZiDXo+uvy1YIAB/kR7cD1HN1HNMmS+gs3amRxluZdQnsxiPNNDe
rk1cxFmRWNLYjHkftB/vlYMbLYXPGdTTgFpeFyj+3HhJdgnHuI+xoAo4lq9rFgWM
KPpNiXuNGuWqgyQ7ZT98z7tChCgO+hVURvXOvxecPBum1BibnT83e1tLjx24Ueh3
4os94z1y24Plr5UMf9fJYxwJjh2Re53Nym2efb4cH1bjGtQlADiUvtUINeURRTfb
/LZqgDHsnASAeWf25IzIj+c9jab/atrc9GS0KRN+eUkTnF7RR2CGLyqSEC+ZlCyR
BLHDgp0R7lWjiqjtdg/WIt/2Oqx65dbxrFGOP3bwzEuopa3jfkDymgH3lARoKHv2
3BMhNokd88qw4aKmfU252CkO1z4UNYKMRECNSyRWNU2B/g3oqrzlDWyeymgeWGvM
Gt7HZ0ojj1l8DjAqtAfRvEqYTvsd83KH5yEts+Z0hwHahGjaC33Y1tjo1QjpXEDb
PFTrXQQN3Mj3Zrbeh697YECZyOpJfyAU7SRFj0rLPmTbk0ejq0gEwfZbt7s0EEnN
2hbZk+pgN+RPemhUGT803hYIwx6Yu57+9yUJDqQITell254Xpl3QoBsQBIZgEsX3
fCH5VDYtYigjR3nj0ZVmRkPHlhYRcLRGpsmxF/13P79dlL67aEiWVymsQzluyVjC
cCBgPaxbpzvntZNOxXIrBkgLY8llE89zKuVRQiF5mEA3Z0R4yqR69gxHtkCoCTC3
7sm4My+7dzc4sk8391zqB2RNmJrRJC9e8wUiIKmgHamKdBGRwEUXyvju9U0pXN+D
oMqYezeBevorVZhcwd6lkhJauWS/fuTEB1z6XuQ1eIdJjPBzEQj9ICX0yzJH6Exm
6es0bxf53nJ5hogpkU/89GX0a6IiZMdww0YKM2zlNfLjM5raUmc4032DIXaEnPuT
PTICsQpe8YdPOwNWgb6UgYL1oh7KAXL2MsUL5lHgVc+0ZofPd1qBFRyFAPEu3ktO
JEfvz6BoucyC3IBNRsAMy/KxbLy8SpfQz2YtQnVmNCu6rBgpvh4vsKCtaKpR5XOl
VSW3ofb76jQY28fIjK1W4gWsbJ+c72HpE6frSlGlhOlWiUtnXClH0tKtQQzVhIWi
Bn37cK5bWQ5sx0fmvF8q36jSjC9yiDWfUpTmSfJTtyTqWpGB40IoLr55f8Lp5Kk5
I+usjCNgTn3dpQe09m5SfnYRhMYfyYmdf+pXchSIa0VxcgSmIKNQJDrTorB3qSlX
wIIy9cIGQag81Fb2lNgSqy9mTgiREmOMp8sSaXeGkWKiBoVG8PF1FUvXlSfglHca
ABDNFzlYr7bFCyXNczvFk8AFb9TH8PDHBBzBtqFihsiG5cVNl10iifdXNyu+T+pF
0SfsPZmiHUI8T5FG47MQn4XMRiTEyD29JP3hISQ9kiszfwLmJv8MbIN7YbcLjuir
kuxZ3lLrOdb0EtnxcVlFd5bBVu3jrff/NZCdlSY8xjmGYROBqLn8//5/cAtlMV+r
UVkcztWYjsLhUQMKI+JbAoDQPs+0mr5yfgDgzNZMK4Ir9epqxyQ+z1CKRBsqG3Cw
an4I+V1CcEK7nAL9e0v/6hAXVvFhkX5kylnb/m50GBdVJuQ0Qjvn+mAs/W/S+UZc
DBcA9w9jb66JLo4fkh+mNXf+vSlZdMWw0e07wgbhMLyx+tW1lWIfTX4sWBjTQxRi
IHalvpZbUD3iQHEEcNegOLGGeOZqJsBxgJPTNLqx9RDse6dCQBI8jRVZHQFg1E8Z
iM9g3npkDSfto7nNayvWtTJO6jBL6tahtsDgi0kyG0vz8jEf4RZ136pFz1w/fYEV
l1WQI//DREzAvMe1zE7vgtEFePzY/p5iWy3KjNWaWCDcmsLQMCzJrqaKUtyT0otZ
WD8WnlMfx78y4jn5+j06A2kSGpkW8u2l2z9GcxwG3PD2mOdLbb8FVmjy1aiGpYvv
z+ockIC5X8YPyKRO48KoJ2iSdz45vVukYDMr7iSOTL+ZzOwdyKqOu+blAnNvIDMa
SUtozH2Op+asNvw8Hhj6HRs09tHCFgdzrpxQUOnXlsPk9q4suEmBHL8XnMPLS6Bq
rVkUv/cCzUFx7/XVQ6Tm7YghAJ7n51/vQdXrR24OJnxbCplwdekCld14l5eyqdgf
qdWTp0jTJvyijUh2tWw547D/VHuyDASXqIFbOK0HT4YUvR5UUDmGgPtxjiUiJ17u
rjGYxCr1GrFerCnDvmoLLMlgYwQU7X/Pkn/iqgDqdBf/uAHl7NeQW9eteOavkN5N
tLKruRzTzVURso342Tx1mPBXmx7+Itihm/y19rhNJHS/Z/P+k6v5q0Qxz0dSvYaU
liBEgIpAfjWIKGzOsMEwdW2cg+ybPIl7ChRxVg0CIe7fyDe+ksgAx+PtpRD0q9Yy
ZlArgSWlxuy9xee5Shc/qzyrcvzYq5XSg4jpW6trD3w2ZdiYzKbqnGBOKtnTZh/H
vkpfgL07LNss+AuQTnh++weWeAVFGBGjqpmGf6N05PLVALANf0pTZb4Ol0/++Ff3
hlkFQh5aYMVYXyo8Hqpj8ANYKADwAsIz4ltcxvBWW0ryTZ+C5UFFMRBHI9icZ2s6
L9S/IBgEyJPJWxvA0vUmFiXZK1y4NHT2Tu0pyJ0oHgiGZb2asi7hyPRQDsxZrwNj
hS8JH0BBBwxD0Ne3hUH0sxZJczxUQkNMogPQYSmdBTHE7PvLcccKUM37nLhYQtYW
T8XayzoGtvdTACCQyD9Nlrq5LUsCrxF/LfQU08XFlNQfjmBSUjzC76GfI348VZ2Y
cao9wHys7pFXoXSZhdYa0+OFKtU5NpsjHh+QDGkHQaN3lHWBlQy5KjVRWA3d9zju
YFk2cD3HThLmZ/mvxZXcc+1qaWi7+XCsY60jvc/YERzlrohB2ZXvusxtAzJU5/KH
1Pvco8xhupUg/5rAlYyiDSukIhy8tH0Yevy92VvNRuEoDGb26yejHKyNo3J6KaEw
pykX3MTZyy9TeX+3TEYEIa1EO9IWf2JaVNliJHRV68G+UfVGNeCS7RGWgRvslVJz
4woRbJXkqPAhm7aRvHvgfhrHutTd102XmJDFF7rXzimHp2YqAZdnvmhj/P1AfBgO
JcSnv+HY3G6rjRSU2VBWd1LJv3bGp2aII8iwvnYjlteboaWj/AJ3Z/LnMRSxREL2
qetC7LXH56Gpv085Z3uJpF9qkxFcO+XTCJ9Fu+xjrw+0oFoY4df7VWqKpm+csrpg
em80er+UrhqT0XIlA0C5Tm9h2jprC8Hdq/KzguHeUM2wT9GwsUSrBtqZpr9E7eze
TEGjDi9BnANaw7SOlnzMwW1/O0z5yq0INiQzEiYjyTYr9Gr6AQBdh9iuzw7MGBgl
VMcVfy9z9/U8K346nQq/IHahDpg2JH+004pqnRNWFGejOqb6Ld5amHxfOD2EYFDA
bBCuJnCHIiclzJ7Jx4Ejxyziwfh+6S/U+cGNNj9KsMYY6aPaSPvQBs5qWCIcPAp9
WViMs8obMtTI7EcEXFVS0VjroUo2DMtxovYC6eJSKaga6vrv1YIAn+0MiHggz388
9X3qS+/EjusJNqZ995RM8SBYwpC2TykYILpepxyd//gEXPax3lxlqS1XpQDSVITJ
pitYhFJ5RVZhuXLKfN8io55AoaeVkvhDsfw3hKknYdohErRTxFSpovCQDzZ0swBy
BdvHCsnaEF3XkA0Rk07lRhFDdIBoKuO6S8v4I1kNrx8bfyTcsxv3aNq+2J6/xkx4
D7PkoVWxGKFTQndUeNu59TiOrsuuu7oMZOP/PtcMkistaexm2BZ73nHLWK319ON9
4y/Kk1UulTgYND8RBH88dkAZrmb2N6yOgFb6q8PilMvLN3BGDTdPpbrIzQv+R0uO
o9YrYmQwMLI8Cp4CJH7APtcGnmC924RKTUgnQ2IOhANPtA0/rwiHSNPDnkNfKITv
BgxgP3iNwoTZJpXSfRRaTlX+crK1/J83hx7nxHwnmZIzkk3EUVf1ZLCbC+FfZJ5L
FBfrsqKZsF7KXPr+YCTnml/SFBr0cXBCyar9/hF6L1V35crqY/RcHw277rKoV9Kl
kyWhY2zExD5/sXOTzBc0MSlOMvZ/+NZ6soJtKqKWlN/xL/AiR0pHjr0WGp+nIXzL
W+GQr4DTf7Gl8Ehrj4E6AT3yJN6FNf/QkwDxeAJfIYevphvdw2LssfddkE56u8id
0Gxkdnvi6iH+Yo9Q8pRsrds8mto0VAJhlk2mIVx9gPBySUh59Eje5bkN15j1hqOX
9a1E/CkE5VAP26kf48U/bUnf7LU1C5oni+/cFTEU5Ahsls44+rlfQmkiFg9Xfc41
19WPPLwwt38jJ6qfXoWKf7glzaX3Mu7Y6j65LnagVN9bTjDN+y/kna5S9ckFCiq5
RYFpcmiX+SjEE+Y2owxjXIKVgFJ2niyCdaKC8ZBeq5aVBRcI4gjJEimo1Vh810Sf
0DWZ/1Zps5gDAa1G1hrchC6NdYVkAA5jzv3AaYFqzmGDiX8bAbEMvm0wBr4rhjVZ
+sZkrXXtIaDMblBLvxxMfOQwLwh9tLpx24ZAcqXUjSfAGJlBSXwymnLMHg6nYrvv
BRtnmrYT7m3BwX5ZvX0xTGaFXuVFvtyA7QBPWwAXdRRm8F/A91JqkmeVZyFTwVHK
9k6XKUwIaHGi8EBoS01x0evSgS8SJyB6GTRRydCQIQGI+cEBqiEbePDE5nT/Q/E+
5jbfp5x4FEmFA9JzSrXw1G9ouu/FZQ9p60Gmg464ZMEWG9rbsUWrUaIt3pahl6kZ
/lEJhijEQQZqAbKnTX86knBi6r5LSvmxW9JERXhLiwnAtZ5U7Lq+QLnTxVA70PL7
C2zXoygkT336KDiSgW2Vzplt7342rEH4VRO68qPgmOtfKVFrbSRoc/r2N6Vj/yeI
GAPeMXyDU4l53LIEVVLSd6TpTnFLNm8sK4Rz8TKr7SxzlrNM2/1sDw3oVUcdx3+M
HL43eq4tlS7c3+Aub/EjI11J6LHkxLIss51OAw6kkDkhiu8xN7Na2eEID/eYFVeu
92HCPgbdb35S1h5S3ElzgB9yP/tynVZBMWRGUaLKKITUtcagWuQknKHlSYol+PnQ
mg1H9Hk2lDLpuQeBngDhtF0YVa0aUI2GnkoCh5cstFm9JxlQxtb05Vxgbo1wX1Bn
zdkUXfILDy+sf2YF9xeN5CVDXXjySWdyh2Pqlde4yMEDZYnSTZj9ZLdfqYRBFuPQ
VSm6aV0OtDSU5Ygreo2e275Lfl2bUyXVEiG6HIgdPJJIdFycMJt8hMV+ls1lsydj
sJmn/ufiyYBf5Wk+0C4w/kNY6bx7LSVPduSCQGu/Bf+4pTXylxl8iylLQNJtX800
IBmB2V8TA1F1qPe0oKFvgv+5Z32Wd6avV77UzPqBlpSMmnp2m7CuV1EP8UFkenP3
ZVQRtksvs+misbdJiDtYownchgNb+kCMkaM7GViAKgEjKUrkwSeyKH3QlOvvSpiu
1zxmBvDlGcmDTNgvibByOu+A3kLjwVOe7nVsIu7p0v0+8K8jRqGuOIaQ1I0uBTLy
Wd7T278VNyy7ATHagUQ5F2hM6Z6h8i4ToDfY8+fDDUtPQ6LdnzrG6jxSC/k53WPZ
qXIhMIh2n4q7ZRDUv1M1dabuY0gLOm06KTAr4H+aiMgJRc8jnTSyZxIo+YvJzrJP
T0gsqVLmJWTgtmzOwDT5ogG7qW0HFCX1ekavK69SWoSQPPwNIBDGAlA9OsiIw9XJ
T53bZ4jXOIELIYKCp99Ru5I6oYHlgPznEn4NEsFjtRczh4CFPAsU4vyZ0ekrqIGP
EMG4MeL/wEmJRpRE2R7Msa8xqRJ0RAJL46R6Xa4MnMmCLmIFnxKI3G6r1Xb5cwPG
2y0tU8T+lSAS4f3mUQHcLK+3Aa+IiokzBQUPXJf/i+XJPmd7aT49wOWieFEjyBUm
qp4wro1TVEIB8Q0818gP1vyQiabcssnqM66O6Mcuz0Y1bNcPoYK5KaQfhYgEWWHp
zJ9rO16bwv8oPYVmepP+ls15Os7IykLkwlVBEbBgkdMlXcfhq+6Ox6IwA+m+2Vc6
ITXO8BXFwt9LOzGYt2Ne2axlE2ktiHu4oHqB66dM0CHFBLdtxMunVe+ZNZCZUCh6
KnlzFBH1qtqJgkGriD4hnAu4uEX5g7RCwIHXo8HblQqOTS7rFniO9E21mBJJONn8
IH9IDYq+EZxH2KRE0JVwC5adqVGHuw/Obnf4LimDlz25fJdTOacHiA2l5sKMk/hh
D24HgTEF5SLBvvLy+HeYlEvZbjkL0HrnzVF00t1W0zZK1SX9wUY4IqEGdaI36ptB
0DCKLcBMT0f9yJ/WQO6iOe7Z1DbGsnkhhAr1sQAFGRPzn8XU5xVv10QU/rJd0OAX
WneeAGopjrXznWOH3WwC10gxmNbhPQk/ZVMEu1To08OKtV38GJvFU3f0wlCPsFHF
X3VdTgMWF8Hi8uVrBU7oP4cqx47cqOGwFfsthJvBvwb+9DM46iRM0tvZAFN8X4HH
zE+2mdlnU7771HQqHMhiAiXUvr/tCc+kqkkQIDtjG5LNLnRsbCpYIg8+WQ/vfC6W
L/jcXmBPFLaRTggS+kMozpDsVOzrv9gDN17sGSFK1tg0wnW+6Se7LHqPZ6dSx5gy
z8/7zE9FeUEqHQrxGPj0iszukfyu1ZjU9NY1UlJ0oJKx3+D5QK8/yPfMVp1IEW4Y
hbNHjK1qDqNhbwo2+42MrXyZPLRgM1GBNRf6EQeA5WMLS7difYcGT0R5EA0weIXc
fEc+wix2Q/3j8AqqUJk41OojsX4KSqbhORU1SgutcInRHdhP0MHu0x5FHyWJ5o6N
MEM3n5X3opmOV1/V88iT/U71as5jsEZTpQ1K2TyXjByHp+A+3nXLq7sFoGzPJJ46
pjvbbr8ufd5utXzBW/SvBtjtvvx0DGE4Yn3i/k5K0eM3GtrwfQNUhjBBrIdawYzF
8UMwg+zZlPXM3K4Kemo4xrE4QpnGkTIT/kZqQSB7fSGRqAvgZZeohlTSNbXbdv0W
tMDF93WOS8bzM7c7OZHSwVYOkDpHZOgWZZLviA7kCHtPCPz/UL3uut8TwceHgJu5
K/D73TwKQeyPCsmvT8JFLuRix6Klf+Kk0orHINPScVRZlVFMKhUembG9KCYXVv/X
/2E+QaSpbhEdtl5R/AprD45dpSlY0p3HDdOUYTYZ4Wy4iDcvOvpybsBejRn4h4vw
lFttWgfz+SXnc3DR93ETbFhQpEH3xNVqjr8xZVJcsW5ZL2t4mGHUKsypJJXOOnuH
eReEfYxLWONlQ8NKd5n/Gofyl6kDDZVmOimt/r+peWNqAKbS0i3LYB/MbnW8N9NA
oqsz1naw9EA/VprEqaADYCz+z/46N7hiKxu6jjsh/ucG4vTe4q6OBpya9gGVUMNj
OOYsC6mRU4mrSpnklaqs/ncXEimL0VdCbWSkR1uXR5sAGEFpOHtuSz/e1aa2oOiI
sX6+xMXlMUr5G4nzWBmZFY9GuNmZnD6Rx64bX9QaQD5ZvVJcsvmMyAvwTTQQe1T4
3pvafjEpzzh3GQamBahHoDKvDZc056OHIMwxM+uuZjfpMOB7hRxhUp/lKtYJMzon
C2zbqD1ItMiSe1b0RH+dCCJkJ6L6id5yxPNKSEPPv2Bs0XgTHF0WpcbQyWQI8Hp2
4QOzmi0E8DyHX725TMh9lLfjSTsIUNQ8fx39+FF+7ko/kVqHLy7+2PNwV81PLA/r
XCLzMyyOB6jw8IhwH7/OvkWY5I6KrYZ7nxr8VVMdp7TbS7Kk1BCWIqhnOAuYsOAN
HbLw3Pxytu6fABt/5gfm7dOmEL9ZpixKmOPxoMXizAVLlD7G2XBFEF+9Hqwsuftl
XwfdbNDbSaCSoUFePdBC9OnqGd30iLx9ym9cTCE4Syj/lejLPhI8upaJO3B4vs1+
l/x909zcI2vCBRvhBcP/itHvvM+m9ze390X/ZoGzhWah+wKELD5tc4jX0PT8UyT4
0cfvMKXaMkbTI8x6lgXJTSmqIrCCKLhvZRaqeywPRYVJl82NJd9gWVLSE+XxMo+T
OOX5hhBZaAqyth3AQNpdTq9lsqp4BNsE3MMKYH1iCUz92NbUB8l/vhIaF4YauPqn
lOcmmgU4I3Idxm/R23dIwoo0XGZM8/lCn7FHu3petwyMEHhL6Joecmpe1zpSf3+Y
2q+zhQxGXRqHv+yDbyrvmwEYLw2UIzqBWUw6s8gxAGMc60hUHmdQ8+Ou9irKAoT5
ISnexvVn3f+Q1aP3Qo+LWbDu/Js65HcEdfzLsYGkeFZnfpncYMXjj53/wMSfY4At
nTksOhvGKrfTQ8GmubRTsaIIR9NAMXnDPVXDu4x6Uq+zkai9gRKBeSHq8kb2D6f4
tQr7pwPPRAemMEzpRwpsPdOcS2v7iH68pR6E11azZ40PwkpqUcGfyBE+g/1xLSvB
+6RDNlMykrSF6ZQX9WvxNTAZ32isH0SpLqh14WbMVsQ6G8hd+ArTJLsa6EWeoBez
AsAgj2SaST6E2PJGzsOaB6BdqjAjKXuVascsdQnuDbtHI6lEU/jb1a1SC0samG74
BsdZgPolXIq7+K68wikhkJ4g82yNJHIzpuPafDBSfajfYNWB5SIKn6YYzvnSOiRw
7dDLHgo94ZSil0cx9X/oGWHmXwvKyylghNXIe3ocQzlFMCQTT+pEkz7rhwZmX+xs
QJnB386Q3qkIvaDodP7Wpwf9YLfSXZs4gaO+rUdoInlFLXDcJSqw8Ik+DfQeDNpb
micIQdLL/4/mT94HIwDHBALw3cwz+/BShOHu0yS8lHSkdnCq/vwoBsuUkO6kpMQd
aiN7QNEEpC11wi4lzBypWkCC6TaHeacGAQrzBb9r7Nu9xKegudB/AVRvGtIfkssV
eEypTJ5+y5kjnRJ4owiCCEIotSs1cTCElw1pj9x/nbsh8HToSObT3nir2v9E8XHi
FlyeQ/KMeIY2ECC+6ZFDSlewKiCa1hJGV8Kh1U5zOHOTbF4viEyYaU7dayzNN9z+
IkdAVX9gG0g0TtGzQ72Yp7uPplvjY9d47YD2yJBqdPSh3znSYKtRf93aUZcTaJCO
eFHCRKgnRrgT4T/hXCEyJjkrzSOrPABBwpe5XTxs3nxfPwtYpS8J6LKpX1/emkxl
6W9hwu0H/z+Ufsyq9ivhJ3e/ffe6+yfZfNQZZVY3WtWxIbXiLJeLCPbHIahN1TP3
5y7pXeAvb7S9wNjgMZHLVh1Ua/eRfV/meZrZLuQ9vVVg+whVZ5nCHDwYyzzBW1XM
DB+pqeDa9A866g+Ar7FPgqSBMFq6r/RJRTZ+bI+A1jpYa9uHaL7A0hidFIgMRIiG
edYKRrlyms7ENSOw9rk8bEzfqX3gI51jywmzyk9QvWvLOBmrC3hIlSnaUo69E6JE
VVLzB2+nsyWU5E55/2JU30JlPTaKbsEE+2FE7ot8faPVW43xw6WVC+mGSN/rNcEj
Z/55rtm6MLbBzbDhv6YtyRr/3azZjp30ER4EdwgLqfY9oQgeIbke7K3uZzea/AvG
2EgWgqLEupdb/7HKm59X9bUYzFrSm408vF+4lcKLgbC8uK1erBQDDgQZ6UJBZNX8
gOqEoz/FisPVe0+KMQvQNJaHPvKhtT8sOKxbxggEskp9kG3AovA/VYDhXX8YGIMn
0FcIvJedce97lQY/gE67CWMTSbLUF64ClC8wPQkhRFNx8O/VA9mlLwUW5vUpeXFo
m6GTysTtUnS5MBYDFpTo/NNAExV3t4oCzbsKJ30ojWIsN5BF561jF4kCUckNuD3S
sNliHJVQ6OsVb2eTCpYhotDBxPNfWwgtv6qnym7r7vDqDvED0kOnzlmX5W6IQaiD
w4fPN9Crqfqu0QGAd5Aeda28HErN5Na6qdTclYaBcQwAQo4C5eEHiHve/BeBbK8m
z8aZpGadunRQIscGZhlwrKNu+Z056CSZHxtI6sFr1Cjcq9ukKfF0BoZgT50stPuV
wC36KKeqRHYHzn+VRL7VCeBUeAgUh22OL0wUsTuLpeRWGEUeM42jD6DbyuDQGlI2
Ie5TTg8sqXfnDD3xOuAaOB8BdbeKcFVlJxavb6tspTWDrzDCc+zNvkikxJ4ErslD
jgpqcAN1W1SYJjOB/07s/eaQffO8j1K7sen34P/IQu2kkRwwRgKUpz8McpDp3DwJ
Q0T58tXI/3gtss0MWUAxP3AfvUTYcKgD8OK0EPcv7mWiPf/CslVew3PaSjj/ixCN
qQ4ftbO4oPpNX0E/PNohrG6X/KHFnyLyzNFQ7caTSRw32IUUB4wZl/6Ojk7lTKoA
Uc+s7k2ku9elqH7deoo+TJchxSow6HKe492sWOjRcwy9PRiXx2k5Pi0ApssZCe8p
H/3wVlKZRFNQURkP6jM1WOr/gnomk1BRA1JFCXPL3gYgODlTbhLMHkFHxBfqTsSx
W7dugj1BLelxCH7fLLxFZLNnPiP9iRbrZtBjrFkOr8jArlC8reqzPuPKKwwahiqR
sxCLX/QyfSpr7B6u5mjZl0IvXZhlmY3dzJsZqD3Pau7fZYhYDiQhazm9ToHlkNqH
E466OXrR7H2eCfGGT9pRHb+ueQhu1I93eK+aAd3FkqJCXPgrBCD2T5VEBpErBDpn
GlKN8GXBzRp07/tVFeR0RTonhlMghuUW62+4Om1HPM2d1E7aDiIt46m3gdK5gL8/
WhnRHK9OBLmbFRcegd03BCXDuXykjbO8oW3XbkAl3Nan9RZaF0IgbAGG3xqW2cbs
3sHC+SUzhZ8MyadHbFm3LgiePxjFtDcWAG5KV68ja+Gxewqk+kxHL5UOgFbHtAHC
DoLfNxcqdPSE5j0nJCgF9liZC8eiyjHawD9U3yQsDvu6nP77/qC6YISQ4siU6Yuv
8ZL8NlIxQPXjMWv4rwJlEG14MlLpIhdQ+3zk1rCrxyzygAIOE5D0f+Ikz8dZeozU
CvjfswrI4+U/07PvwNRbWrcl7vJNZqBYTLw7APsKnIMTnyD/94KBhnj9UvaNEjtK
0cCKXCP55eHuNTltIzGlc0t5mivgVwmtsfX8P6FLGMtxc67fvGpJP4RFpK4huMmX
x6/oSCMuz6Ykv7i7642aGyLWF9pObdbQiEqQB01Nx6P0bMjMhc34S0WOBeSWN7RW
u5vPJKGmQt2p4gLcc6OEzVDikq5BR2pN6BOhDSeMx6tcPcgcCzHw0D2QAvyY5Atk
Wz9KkLZNugtOip7sHtwI75gEs1miqh1c6dbfOdW6H7uAYfixrZQiizhILmwKO9th
uqE+PQxoFjcWrfwc4mgPn68lLrPA3f0soQ0bYbDmEx8/j21x+0h/kQfTzUJsf677
nN5KZ5YTvsqyyDQGCJ+PdYCoV7DCb3oO46eIrgzhoNYGkM/MiaaW8kjqseZONZD2
v1BdIzDgTDTaVFDjq4hE3BYEB/XDe7Xzd8/XVPPtv4wtWkmd4cqQVlFiFLMtRuOH
zmhfabjnZ3OdItMoIXBygJu9LQg7ROAcd9/vatH7R1212/Kxp9Ck9ROFoHpNBJB+
sX0WH7c1ETbqTy90pmWqxvLOV8vZewkCbdcTgGkDPkxVARrzfyBi16XwMzWAARwS
24YWcWyQf9TqlHNs4tsbAo1tW9DoJFdlH5APsg6cB5itCL3wevLvT1xtoelXkyd4
FqsbE6LdjXt/3gl/BT84tmpZR+xjqwqGlocL3fM8eA9KpxBXJzP6TqiKHh4OVcnJ
f8D0TrjzGWZrS0tsSYBoh6QDXqVtSvOpYMPVvWxD/K269s8XXpliYRH+lrWL2m0i
6tlkb4+22AJ4usR1PCxnARDNRhyGX3wu84xFwst+Ldke/q6sGlsngnHEQVZCs49h
4adZAgqFgke75rRMKKp/aPkCYOl5/CAVTtNPbe/xn670Xpz0bvK2CU7s9SsaEN+s
/TF+ZRdoRXgxtCdsd6YGaqds5Y2OrmAucGEEq82KGWd+wqeQvgt97bkDar0GrnOn
N+anhdVhaJjgc/tKbIYw4ecJa3QFV85NacOlxlwUpB6ysDfGFGF7jm58Ck2GnZPk
0Fk8aCIEgXAECFrwmH8ODLzkkr4fMLy7Tk0KA1+xUfvoS99hMAluE1jijVtQ7OfZ
QTigDMcwK5QnwICE/ZO4RpZ1gZgNLpWNbK8XSIYHVyUn+EONlooR78DJnjfutywi
h7tey3Bh3uwgYp7GlLwkTOzeNv/ET+usOmDEv5YCoeh2wHhroZzNgAN6PGZLcnSF
EiNHgiXX9LIKv3ekyB+rWuC2xrnTsaPGtRNzPD0nRlJ3mCBblEckANZxtAHC7JNS
aSOeI7DrTwEhTu3jU28W8mSVE/Nv8NvjL/+NDyPZHVRX8loHQQRIv9LutBwH5BIg
5eiFzuhn9L/Dqupq8X12/CHD8IETWHrEO0kzk+BWmO03J5saKXSeyxZTHUIxpmuc
yrR9aeyenUEtEf1fW/hHONIafdsEVOCill/VxANhkyHbeK+Pse00gCG7EKsqQ+C/
2aWQIBP4yFK1czbpu0DqAgT9dWMkTt79Us7DvWborIgKtfNC2zG/PzLw3O3VXE0R
sQk9DRG9C2WB6O/B1bLiXd8MUSejQfr2EShI5eUce3NaAlWkYfmCvyfpeSNvweOW
BjZwTgcrXEedi2ZdzJyWmC28C7OzqwISVIA7SAS7aflt4DUCZyqU6cjf0+3iYgH1
IhCV2LzDC/v5UWYFvgyu70qvtJcrT4qtQnmCLAAtHC4c1r81zwGFlzT9j/X/Hml7
SPy3BKEjOI+80zP0N98gLDDlePcgC0/shrpTEG5tC0DPLIVZpS8j+Vn3vhzhnVSq
kxQzDSTdL9GJNhRzV3H74EHlLTCrDlVzhUTDMtmkeAujM1uHVcfFMPbFeuZsIwP8
hcI8pv4PSGqWpbdGyB8rM/4p9Iuubghi3CXpF0Xtn6gCQcAPKMCdto83Jsgw4ctp
qqgfC6gq7w5yWFZf14Dly9Ks1gj810r/yrgcRSqyT74jM6lL8EbFcjRHvwcOh9Ol
zay+ffH42dhiMH8nWYzQomPGn/xOJ8EBBPDo8j4zPA3c7M2VDWHIPUnXc+WVgg/h
1ryVt5J09s0DXtEoLU2fJVQAQ8CatxZEdj2H9Y4Kw5k6o47bs/wB9RP7HA3j/JP6
lydARlh/HirLzrPfPCgcHq2t9eHg9uoG0VIw26Aut0ZJcRF7e9k7lAiOM8aHvU/q
mtFXQKtksPFO4EVn0PB0YWEppr/wxGkY0AxzLwvhDL7xDVIzSDZJdFFykPsvRLT4
qUXQfraoxyqjvHAce4uDTmnVzW4V22UkyxiaybSW71IPB2329OugTeWESqVhA7ZT
Rix7pxrkiKMwofzoMoce6gmC5vQhZ5+YMhC3xhX9nItHFSq1SX1Z4A1YJOKnwjaP
9ZyJJjCqOGho2QrJ4x+ly6wKbXkNbrF69mdFVUuvC6pp0czAaxbexIQSW0J6dS56
EFppyeHJqGZ9TYDoe6PNfReGnze9wilKFVNCs4jlNfZ5Q6MsSXczlocV/v6eG+ey
UgLZUWcOQWXDEs5S4xInPL0TvM18HmMzUxIrTka9pFBg9sZvmoozQWWhHqmGmDT+
m4SkAjNVj7DAWenHIywcQhSPYPeSp+ofCvvh6wSXkJxmknh8CRQy97szZdsLHnjP
iTVDaMLME/FT+1ZgjfvOBLVZ8nK0i3YVXS3wg8+yV08V10dLWP3lAkSIEXcYocsP
s2b952WvLYKHYejar8DLzvxOFoB1X94e3whozB7CbwvWq64oQWT2vIeA35j0RdaD
T59ovnEb88CLutD2UvNc9ee7yz/Rf3zIFdhpUrAede9+8OOxqUrefgMXJIup52K5
cKFeFIMxuMHpD99nITZQkqSg4WUF/gPDDbDAlB2xbEIhKTD41tL+l4A1xhw1Xs8F
YgldkNCxJvhI2sWnVA3FlmsJlTVoRnY9rG/exGg9cMH9+TsrZESRwCICR+ReXcP2
uqk6I5IQO10PKx1p4RgBkaRScNnkV1+Rl1fx314+TgjmOGY0iRDewbfsJGLzrKg7
/6DHwlb9B5XH5JwIR+6T530RnLt+Cx8v96hv8OBv46EDWFv+ThA6o7Hq+BDwCZgP
33KqTyBnvj55s8qN7k8pLfzMaWAnA7byTFo4KetfVsRVq+H2tCiGrJE+HPwVeQlU
ef59G9KDJO6K2sJUPesnIpiGX5QamO/TEWvKoLzqexgSiZWknFEH1k0rpn2YgVJ+
DE+vr8wvp4gN/hmRRCL/k1z+73MAl1u6sUlu0gm4mlS0i0ImiV4CI6zITINYnx4a
nL55ty3EMmmiRJjjOvA/uhhxrlwqhOZU8HlN/4wNciy6YQN1fvJ7JzVpK+rvVusL
X1Kd33lpGmJIPfsMXYEJW+zBY0uqK5Jp7rg3tbTkJf8HtwmGYNAzWzM6F2MdfJ4c
9VIfMOCG55TDB9/a1H/5Ei4jDAAr3IkJJt2vtmQ3lOgydjfdNQGz0k0jSkToolke
0a2/zIvmhgYH29ZJKbSSL67y0nxu0Cq13HMemeV7YXZIopKwWYNIykrSTim+yNBZ
2xM+R5Ex0wWaY5ar0mUGhjxI4qoBjsAm8x+NREI6v7DZQm2QsyRUOQHIW18kAsq1
tybv7cpA7o+mWGP78XLrzA1jqyuTKmOo4695bvgkFqJ6tr8uelayaDmJHfyFskZr
TcKIB8JclvxvVaBcuboFXjSV3JhqqYMDS342AIkG7C7+PNmBpJSa9G9yLPja7g2h
yjCHkPXyKHYx/r78lvddly/6cFfIWxCqfLFQGXjXnfswOMAMedl/3EqIAdTWV1wi
nG1vFPWe2mMA/yAs083Mir77zecTEN27y915NyHkxLdvSFxNl8AOMUXeq3IFzqiV
Jm5np9A6D1+Y3m4YrQPAlEC943ISzmB+a2h5oHvw7CEaH4G9bZR9k2EukT8X2U9a
TsH2e4mrpnvKcMoWKARvgjnYq8xl+GtDa96kPLYMHojAgeZEltsjap7/LG61XUdA
cnzLwibGSAQJyoWfr0tpur6A0/qixb6I0gahIEvD7X5c2wnjA20MnzoMepYmz4ST
LIapPlg54l9z4I8UhcvafHvQ31Xuwg1LTSpOmfNkOAH+L5TUAVH283pPmLfjeA+4
K7Lh5O6DR+711MbuW4VRJWEV9uZmKNttszIFvK9G91xoJKMmtFoSrDxd74NQ0Bxg
PfM27+bNUeTSzO5n9OYfGwuqH+4b7RXx3BJJLCnQpf/hPOII11OpvwLEnmJ27kii
TnTWnHMDrz9k1cbUDSCzpEMj1y1qdiiyHt1ccOs3MMNfdeJAzD3LUA5G36IukaBn
rcGnKoEFPn5L2yXbhJ4VWgsy/VkTUERMj62wCatiBRer97lKXgjpj78PZi/xaQc7
DOMmd9qjTpu1pvPehKZeLsJRP24LVpzqtNxRLQTzXzBZliSBAn6p8bh8lomwRrMK
p2BMsp7KJ6FvN0aXoqror/t/HE05/XOIX+A8n7V5JvarpmZ4ueb7hSmXQqtRUiDN
wLudY1l7omLCo3xTXuOBazTj0Wn7HtSeotoCKm+gYxiWTiuakQXdjk9apADS9qrS
o5MUGojn4KUZI3YnQmBrPMta+ZWOJmE05lH5VJecvT71SZx5jsFjgYuIpBWeUyZv
PJ1MxkW2i4czaREYCyZRh+RZHVPgnSQfnFnUBDtS8yhL4AIMhEEz/N1ABlJvHD5V
tBEO//qpRJVtnel36SzZBZvv+iyv9V6kwaISkul91dyEWXale1ysXcLopkiy9Ba/
/kGBKwLskvVUNY5k8je+R4dQa0xyayExzUcOKw8lb4Fu8zllrSJQrajjqFL7ivuH
kYomHonyPoV4YmqOFdN/2D7KdeYZPi+w3afXUrpC7y7oX33jQpUqSX/rcZWTsAEk
pc+AXhBNbX6m3AABvUg+/0YZru2T17+oiDVUICAHZc14qaXMuBS9vtaU9m9mv5/W
97610RKfxr8Vp7PLAiwwl6FgFvv48EMtVYmkrY2JVvFoH9bs0yXMqD2w3UKECn29
5KMCqTIlF9D+AFq6FcKyyrKOprob5ME4WDWE9OuIPU9LYWz/4e+r1zmyzREN92bj
UK+VaDKfVy/gXJhw3ULtVh/OGnRRwOLmLhgRRvELgOVKVX6YNMBeZwPqIBMoGV9J
aGf+rsavOyChai0DbpoFL71cjuziXf4XdR0KF6kLkqHsd0z7103eLJwo16YBo78u
jjWhu0r0+UIIhizU5vrc2/W6x7+S4rc61ZqEGsNafe2SA+tfN+C1ilTTFC0cDB+J
PvB8PpkucDMbNsB6YZbqpb4LqZB6u99xjLM0WLIIj/bDFoOGouJw/a1oxVojOw2Y
98usomTjWUNDh0m63bkG/JPxMTakXLaJzGIh5l+uD5vA15D3q99xv4ydON2lvtU7
GwblAC5/8eP49I5ZE0Idt6adsQWrALQFUFhaKC6aiV9WUDSR6/dHQLe8z+OrqtSo
oY5lcWcvUB44s0PgRX/6VZrCy13zt0PFCeuWVOUtNNgBXdfUEtv8l8WWBeVyNSmS
URW7yGatlUct3RoE9ydS+oR2fGutCAT+lnzXlbELy76tHgwYG0Sw2tJvVca3J9VC
jXDKAvp/ABfuzM2C7UDxXsaJgdTsNqA4cydZdubM02rfEfJSDqahCNwXSeJay9bJ
n3eJbGoWDL+y9FyrwUqVyP7NNwPDV3IPZkUqKk2vYmt3iRbiMuJhIPbosR8e93rD
vnbOhOJzwSG7bQaxwnxMUZUFUjIkcDwy7tUQoLEqY37qFbxlB8c08/etB5cR5tYE
SshNifNIUxlS5Y5VndoGP/dEGBiaUkTgJbSc/dyIGymF/Tg7D2f6yoZRBHXn6bV1
c9f1QWXq8v5WACf+AJjW/BTeMCu828H+AzlEFWHiCG6kNVfavez8XfnT+eBj4DSm
vx8/I5365wH4lQ8qbkKTsMwU1/wkyiyfL2uVrmJpu9uIjBumXv3ccOVy3vOaf/U+
ISj6UnAZGtr4WC5XJo7Bqxj6av4MNL9Cgfm8glImhrleW8uTJfqz295tpq+cP7Ww
+/+tnJb0VX+b1OvrTOdO1t9IA/bqw7HW/hy04BDdshMd1n3xdUXBiGNnYgoNgZ0y
RrAkPKKLTb7daRiU104G9U9D6VjQ4shAA1s0haHeKy5JC7P9VEvuzY21HNYqtqoW
XUojjhIfjwlQ7dymK5Olzj3SswV8AXhriMwTr31L7IShTGf8bSSheqgUDXt8Tr9s
YIAIoun5fAEX6rwa6C7i+LoOopQ6xXWTu7h4LvWa+j/kdAElOAfyWzRxm5HNNtc8
RqXOLZ7fV35DaRpnrgEi5DDUPKozf5kabrhd18xAKw8Gld1O4peDcxTUFnuaORpQ
t3MYb1aOQb24ioPCxKOfuf9Tey5kYpoyuZI8O1pyLeMAWY656u9BONGcZmoVv0U+
DWj3g7s8vB0tjcmJVT/gBvzW9KsUD3tnyWeqcTaBqb7FYTOqdta7sQ7T4Y9dXLaQ
fB1R+z/pnP3ey7ye2owbPuNGsr+lqiUkfwmBKSnIpZVELcQXy3F6CP6EKdeg4oUH
g6v1hClx53cw7SEIuOFE8HtTX7E14pIgsfx8vO84AHN7beRmu94CD1swl1BUHIsb
KlE4awc/8iGP8MsIMTvjxscPJkoSTvxyJ0P0fyZMBtAtFmF9Rai0wEfAcrXX/j4R
qJhOjQvwVGu0r2doH+qOVJotLwpPunFyrSUOCK7/eARLKiY84nq1MVCvF7bSMHSl
ZYZ6HD3NnlUvEc5RZtSo1nkoUw7eYfEXZLvsHVc+Jq+Bplm4ZqbZ8tZZ/8E/MceW
FD4Wdfbv2OHjoxMyDdtgSI5K+d0kmh8m5YqTgxpk1MFtNeMrhf+QFGFz4BZFS6WW
VQLftq5q/EDovy0Jx5sSmWPZhuixVBL5MMeT8X74o6zIgCMlZ14eSTexPHcx5sdO
zeYFON0lYjindJxAS3/ZdtK3GKJX2++jnXrn0IaHHIiGQj5l6L1+/F+lvsoEmN6w
PBGCpTIODGxI0xuM0ZQ+9sNMMMm8J+EFFql+sFsxdyZPl3YHxdlCglp1MaO4pDKh
uroGskGErgQT2mqeewXhcjT+0s28mi2EDs27qXRKgno1t0LAo90GtRP/EmcPcwWc
TqEwTmKV8VGMyUoMH/VNcpBoO2CvqinpfV11wEukAbcRiOs/kEunpfmvbh2n5s1T
E35VdL5KYyVbmtZp8hnInu6P8Ehl/DfuWXxqFpvtrqpqYR/6UCyfWYljp2+EE/SS
vUPvcxXYWqJ3L+vDo+oCve46ffGSftDtxq90ZhZL8sMMnQzyLvqE2iUjDKxs/doj
nMfcznR42FjxPkR/WwGuZIWcX2u9DEbjGHUQmQMOW6d/jlco5PxG+rHfmMBSlq+b
nv/yqmt9ym9JuG4nHzNsytzqUuQ2QPQmqw+ottKuJMzNhMsZ9ln9zcCG0wHUujn+
J5aoFWJwyKYMRcxQqvMLuy1QlDOi/h/3l5F9DTH9jZeU2D0K/dXtyyIFZ21raD1U
g/9q68i1I8FdAkG6eT4p0bdZN/LqE2zTdWwkpEWR0ZD/fHeCVuJdtjIFtYf/RfEu
Gc47jzuUIbConRptOypRGE4H7BwsQUfrt5RiJfNIzMeXZ1QhBUA68wFv3mOKekmb
uiY4owrLpmAwvl8pzR57oUxroU7IoTE1eVLuHU1Eo/xJCQ/rNe3wjIY4U4VVDVli
8qrUrLX9rtoAxYsMgOczOdvO2i80Q3VZtaKsotoEFlaA+W9UMNf7m6cAwR3i7/Gc
6+EQwsrWRMfLOogY+ygawF13iErgd74z6TN1thvndiQPGau+WylNK59Xbyoq86Ub
0kxFGFeCwNK1SyCp7/RxO+pHgZXrFqeYJLJWctMdPWip0f6ZwF3keTYnZM0Eh9pO
8q/w0YTQw+x+Sn9dg7y2UXDMR9axpkYZDy5rMjLzGazXj/x0pJwY8eZPXuZ/clD0
g5FVwwq2w/n/qsDHBfc19DJ6SbulkcjpsxFznz5+/C96VRLThUHlc4qgotLQ3ZDf
YI3U/1b6a3pXn1rlVqd9OAONOYlThLJkuaEM/ZREANmmt7p/AzfX6XRGmWil3eZb
Z91GC/0F2ejM9i7B4mQd3222LgWEwqbGZRAwrKPQCnmLf+Q2WKsZNBf4WDkaIbtQ
3sGJKdEHNnMDzFsVCfybkmcks9dByae2eR4InKH4AdM26wBEilMk098LbAo5Ixhc
FjuDhL/80VSmzwHeXnN6zUb+C0TldKGC2m0KtekZoJpu8SSCuGNf0We0ByVF6HT5
xT2lHMfHdAoNDQT8LkqdspTPyNQygT0NXuSS9fettRukfABap4WIA3RzjMOqIclC
w8S+7U7koXPQGplDSEu0WS7Yqbr/vY0u86QFvnAE57KgaGbHBOObYDc7iEvzxh31
mMx7+GvncW7vhDZ1S627mFfgs6IvGi3CF+4KAY8DtpHds/UmgYNRd06CoGFBnKWz
RNvUm4uz2Kc/wE1xKxFZMSyedwS3EHS6qdy3A1N7fV3gQjCLucVGNol712zxz5XR
giIwukI5KgRngZmYx8u/lFQGAgyRL5BwHSydhC63t4CPSBcZephfwgTjhIoqrStv
UEYDDt/QREEbomPpcLmuB47NEm1nw4BCNeJUBLNMVK1nJBYmBnS/IQbBXLZBeT8R
tHzKAx+xTyPr2giYkndjj2goBhIN2ZLfQYzLDNB+xnOUkVW9UpfJNlYrEnfHndah
MGnU8UjyxlW0SRNglBB6IoV21wN3skZ9ei6jpLxI3O2wngmcpm6KyEHfLLjNfJjp
QmJghMI40IluZRzFViFib40L6VtfiBosg6kKS4yxjXRvA49S8usM0UZb9YwuN8zt
PyPQEOc36bJ9iChOacaUDknshI02xuO3WIYGJve4JmiVFaLpR4ZF0ISPnL79d1s8
QkllJQLN8m0R/mB6VyA252eSJ4auV256AVKFXsmD+YNrEFUyJVqplZ/TASUW4qk0
3FBGzQuiuxKcDkGs4aYsP7/uuEZpfE64sGuPSkGo/jKA/nkdLUUJ15cqE4H/3whT
mfNMyEtvIb4op1f2eS9HBUHIVtjVV169euX9ipwrHRIqoDqD/nRmlGuOjSrWL7T2
8dNR0NdV63gfZHHkvA+5ZsA4jd85VicSZc324OOguigiR1FL3qlegT1YOJWmbKFo
kcJGG+rfNKYN+bzvx692+Q1oEvEM+X/+WtrWZjb074Dc74n7qIhG5+N53BedfFwR
rP3+K8n2gOW09V6EfWtA89rmkocCM+sih+iVINHGqyv4gO9Sb5zXA9+7VX/2uz7/
nH2qP5W4SIQB8khe3PAwWh1GAVAiu5d2/qyGXBfhLTNuqO+htrfiOZTCXG6WKvE1
kTxhppGwevuZqn8Dcpmj45Qh007yCIJhiwF5173oIBnoY8lS7yu0ixph6WSA3y/S
P/6FLIyRoMngNbUTQLwsuKNC1SNEQXXm34n2+XbtIKCOuCFQhHcHt8VQSTZWPXTD
5saspUOCBXJh7JVFTZm4ozorSIUbVdGQyCbXUNy2e2ftpEaOjffFN1a3qIeg8eSf
BzVXgUWQtpEOuSz7fGei4BH5kSt905WrgHU2FM2b12mnB5ccEGIYtcc7p0q+kFmy
/s6MwhOeXt8WdP2sRFYOKTCFvfGNUZaB8zsfaVWQ+bqnCLN7z1oCqu0vy8xeiZw9
f+qQqHfdWaVWrMoXFziqG/LAPoMu5Bu+9nMAG28lNlYnwNMaSsuvii93AnUaxrG0
jz+ePJ2H/SIB0o3sG6ukXZSMvArB75CLWh+h0szL4OUGnXbJ8I5RIp/vM/sisHwS
lLfllPMn0APxpWbKlOxpiL4Q8Zi6Om7VuYR52iFSzrnQac/MJ/xBWgcZj7pzZb3O
x/vBUdMJVaa8RFeAmYVgydR40P8KX0PqpauzQo2jVTBoH4bW1HRyZf2dWHB2XyCI
6+RyY3TXfD8BdOLeRM9gzfqNO9SxfdIx4L2kLK2bz5JFAveDQSun0PKjalHQ1etK
Jxx6fPxlunoOMKPi66n2MdEqJ6WyNM5U0y1alXPp3Qchre3x90RF5Slm1Y1qJJni
+es5+/cIIibre6zNMAIwUrSrDudKXI6N6B7c1vB35mEjtx2AXftwyqJzgZcN83hN
yzavJXYFV1Q9e2TR+WQ+4boRmaBHJSCpCgHIn/nS0AgZjStSM/Ftk5uw7rZYJv8V
bOEGD02wf00/cY/PiBwW5iRquOdi13I2S5NNJHNPDzKDbuWY4gaekCIYSqEzFj+G
0uHUfNKqFErYbqGI6juEbdd0wyMCIAH6orPM2INnF+11ZofZGku0KnKBq8qbJmbf
/BSHZB0SLGbzKIFY+/Yn8+7snx5qLUz+HpUNa6ylBh/WNUV2JXkKpDIHDvB7UYBB
GN7kZHfwnbTupYqEuAjysQ6zQAGU4QUMSbPn3XoweNaqapc68Z3C/Y2IpsHmTWM3
cAQFCgJ5BnOeigU3MOpHE3wjhlX6bCAqHzZIxqdiRQLHGYfbxN+bLYlbpbNNN6M9
c3n8w10VumoZbE78ImzCGUv+s1R3ik88fkDC/fNvsb7QhXpzpYnogEsBMQHe8Pum
k/bKnjHvq+jTugUcFmN6ZqJqmvgpBP9qP7QcoZBvGo4lseNo82lSqVzvP5wDddHH
ozUW9qxhsz9AnSdnplNJT6c7+9xWnCdAiTAv5ku39iNLKA/X1KJTxtdMHsl36QrK
usXHOIwK7B8n8LjMWb3Jz0z8Jd5rHn9CgQMZPnMpKqHU1nbxOwHUsHfAgu8O63PL
kNwnrInucO0PIXb6/hh5TEWo7JOuH9++WLcc/VT3vJWhevF+p9NcocvUoUn1fvQD
YDLrGleAJlfImg5Jma+WAEirg/o1ml2yOMjXxaOYg4D7pvb+/SgKogSQwVbkoWgi
//SiGqu6JOf8iY7/70JC7+8pU9JsDM0j3BXrwGFX6KIJEmQ8+01ll+vcWS7iGJvp
i6w82mFUDV0LDG8DcfkhpFqI4I4vLEGamcY+KAkineyBlC8EdTOG6G29rnBL518X
0mL/hNqLLk5ys6tdIFnXeHbaWHO85bSCCxAGEsFYS8AREhHT0GDtUSw7YNdh3Xiq
N4TceM7tEGbAdaF6jKnp+e7YrKUCNO4CiOrh78/IpiPV/s7YnylamSpm3/0y+OId
HBqSLcoC0BCsQvH6ZAzbvwmoRGL7jOQp/a1Nfce/A1ub2O2/MEnVqoONbU9qc/3m
5k6hi2xGTNFJWMh/P09a8BhZBp8qAKTkZ/dxSRRFl5pwd3y+pbAJhgb+o79QZxIB
wc9YJS6QGWlN9HsN6FlwFlZvrbmsZ5PGmUx/gLiyemv+7caNbQphKh1Ttg5ChLBD
B7/VJuAJSB3oU34yVfrn+dzWqU7Mmk+/EmNNf2ta6niJFRriyShdE8Kl2BSnNYkh
LBAABtIRFtuSImYVrAH/OmfS5ct4rsH/NWPP17VhsBwH5dxhx2L+iyY8ktqBdZ7r
Hol4hF6mqNc9ohhJKCbnDWae+JCOX/05ktDzN/dUExGfmwdYJRu25l5xu7r0KNpD
KWVKo9kEWa6PFDRfc4vzlhJ2L55aff+LO0gOAlskWF67D8r/aOC9v9qqyR3ykqxX
WFiJB9aUlnDDu9GHf2KAqMANNaYyPVLgoWs99qE2sMmynOYjP+Ka6+PY9a8FGrW4
w33WDF960V+e0kDGCyAxwM6eKqpa8VXm8d75EuFWTPydkGKeBgVCkRtKcHVqY5EV
9C5dcYGjZIAodrm4yl6Z0G2NlJKh1HNZz2tv+3F7N0OKuhhoigP2jCctVIfwc1ui
8maFxv4yU1jNmoky78F0kPX7Q+SPSyPo8b2Y3GL3r+l7nFW/a2Z9qLfX1IT4xL+n
lTZseSIgqHYrKhlLw1rVUMcSAQ/N9tgBzCazIbU+dyQcl03vRo1NgWiv3zYWN/YJ
SM/ZwKa1WZLvr9NkFZxeDqcxx08Fpu0T6xS3BWQRNcddQGDsdIwMnO1JqQxxqYBo
muifTHuuuxkoGvJKUbz4Nqm5YZNEZPP0KDSHk3cDO+fptxw3HEsxKnhvEFAgyOuq
aQlBGrsObWGLxCjo2iZjShJAZ2kQYdiEhdTD0crL/1jg9IaZ9iN9LZA0ov9DLAyw
Fzay76mS369E0Uz+/SEdMyF+nLHQq8zLtHup8uMzpfctbd6IQZ6O69kNHA8RQzI3
BtDtlF3e934XaFKFgRDbIPVxISf05IM3WRH+xKX+QAWw4DaSkIK1Yhi8agSy2GAG
fuAWxhzFETReKgraLhGlZVsAAHMoMEabQvZbVImjaIU1BySg98VolWjWkWixfYZH
/NGer9UKGIa4iwHg3KVhKH5DuzqEYV+gt4sWp4eGYXeLE9Pc3CkKGI35WKqM6yG6
uWqtVR0XHEmNFFE5/SZmGegtpZyTfvahg9ifxp0DVRemP5LAIlpOo4/ugLqoqKwy
wh7bAyiEq/PIeHANx1sQuKBLnNhsNz+1P10CiJQGWiAfbn/gdVL7MWky6Yi6U14T
zrrEAdvhskbCJNTQtD/S53A4Jizr2fQ1gkQYq6xUidfk6dazAsX+iyFfrZVmwNR8
GypyFg3ztUXzNJdVBvh60TNlpyVbQw0Jt1ECHEhRJ/1IUi4QxiltYmzct3g0C8/H
cwHXybxjOijFDW+7H49mffgdMBKCw4E7aBAbiiDGvj32cBis0PaydEnrU9uKefM3
RwHcyQI4ez4akbKBDjNFmql5bSpy9SL5iBlCf9Bvu74exTHor2iRWZDSlTm5ozmF
DHz3gasfRMimEpy7wwO//6Kh/oEJTsvVSm/4DamnApuPm287MwiK6w3Pv7KbHKZ8
w4W+6AvYxiIhAuWy+u83gIwJWnk9IasFFuLO6bxzL67dnvDWn75fldEdX31R3dng
lyxd4puMqpckInvr3ivyST5grzTgYo1k3Tt5bc1ubFcH/PxPggyCNwDyY2UzPc19
NPkyqBbmXOQgtLLLU34u5M6wBRE60BY73kuTMwxehy2rcbLh+JYx4KH2zVtcGKvs
Fw9rG/w090k7HErQybQFJUUD4/RCvTudtzKp2JBZ6XOvOyv37hZ2TjbFyYahjAqR
pvb9l1EgAdQfDFlLf4A81mSrrtbDUk8EZmCVywJu2HfdX3KPVEPPRzLa6M1ClmBW
dGx3yqnszZnyvBm0iJ3mitDyglfEyPv+sF4pWnqeYOj4ZOh6Yx9tsFtV3DoxjYEf
NWFpsCnoEXdth77gbz2R88Pp8Bq9/AIS+23SLa/j5GRlsGzmy4GPZEAxZFz4wlcz
X1XJYzbCooBjg0M8obYWZSM04IM7Xz1LjVx6PeOpyrx1GQnqj8RvUBRGtaPh0znQ
O1KkKNqodMa6EGL4IKmsrEhJ/weH7Y9qLqIH2+QD3M0Oq75Vl2qz8k25kK3kaEpj
Dncdlqbpg407fz4Uf6fdhzyUwoe2wrlXRG4PRJ57xEhB0Ggkk4cYDXCmbwlKIlaE
PsvJBVONhZ5Jveqk1r2LhiKs/5xVgKGrUE01+Y4gURWJjgISSEnsZWu0PLWcYTxx
+cq/TqrmfjlF3pLINp/FyYZqJE7AHlwCziTLNrb8PxVzEXaGWIHwblMzwj++RowR
VHuKIHjBcr0wEQgYRejzbAUVDeQWDG10Tz8udEs/N4MN5vVdq10UgP9lvbAe6v3B
eE+fB+khmH8wyL6cqNCmPxrB1Mwk1wU/430fuQ0tHfdGQDD3WJahtS0TlXg8Rpgk
cH0RCtBLtBa9SZRDbd5CQJoRyXv/G5LGjVGXQ86lcBQnf2/zaTSLxSufwG+xQk/I
ki7HY0l9B69KsMfd+fezqeByITJW+AoHDVeyvBt6+tjnkZMBUXL4yjwov5VFHTIX
ssgZXSnu0zbFTxsewqERi4R2vVYM6E7KHZCBW1yGCmqzrZsMY9XFrlbIq4Sxqj5p
guGWQN+zLliBsXppwN9CcmCR4Bqk7K28zDXPLOxPgQxhqs0OUty+5rBATJ+v/Vkz
c2GS20BONo4iFnmieSz5QErvXF6uTGvNjfeWe22ry69gmGVPGwF60FtJO51EASv3
uOh1Cl0u6FOuIgZo1h/eRFiGHwDpy/AoH1M0A8i3pK9sumY5armE1Zos91ZgjMcz
FMUu3CbvKTNS5WoRfvQnvInz0GXljnWl2TyagLgeNLbs4qQQLoRWUoNjQDp5ZjrQ
DFwdW5/WvM0kxcPigADMQ5i+zS8KeY/Ijfk6Eyfqt6uN+MOgCCItUKQOdb8eIM8r
Ie5O4FHaz+hjof608wBCHjoq/FKoa8yxtoIkSHB35BihMtozti/Q6kL9qK1SqK8H
9hOr+2DPQCdtA/RlxWUm9zyleJaGHWgpO/wtZE+yHAwc1IX39JXgrvMeeItw+jiR
CFW2tEZmaPviYUJu9nFqVi3UEb7T1Mz43zV9+Al14ktgMSLfVpwshtYQjZR/oozc
O0p76DIc+KoThmjD4qJL/nex4+jJV4ZjxzLOUwSByLoVFlfBNLwrNi2zQCFcN3iB
izVWoZ1l06oZDRjo4cdH2DXHXAOjI/0Il8noLn3UXOznLf1SHVS4nOdSaDZrNTO6
p5opXKAxpvKoT1IbWoYDFk4pY7JXAJcRwye6tohmfsrBIrAd9Bg19Ta7HPk4gqzs
6QE45D5rEsjQWQTMI5xgEwSt2CWGSwBxq5+X/Nt+SKdesDowsk0C8KqzBdnllXrv
dDr4IPj92eZ3RogiFg0xeYbrf0Uo6D/qcWUhcP+Hupj1iiAnXp8YelPAvjPFJku2
MLODS5vF5CVAjKseJ32tcQHjGsmTTmM4LQaTBeuL6t16XEsBEabDDoapyqk2LbMI
fu8kk+0hwuVqAkBkK/ktrsSsLGXJDE1Lje/RZRxOS8a4tegQNHTbEFotV8ZjSgZM
wMjj72sV6vI9wi3tHXkaEDICI24zw2xhjLxKoGLuSCAwzF+dxZRl9WhJMghea5n6
9p0Gy5bO6UZ9DS5A+qJ1IMVryXT8rU9UCr7xYFCh8N5OWAnkuRSzHHsN/gNvSZVF
UWh9W6itKay9b04cB4IrHn/vFbFR0Pcuv660zUBTI8QuGjZhjx7evTXSWLZouXRD
83vOjWK1umenKZJLpq0ouGawpzW4cOYrSLJAeQZ/WK0TLwKuqlpv4KBGrZ2UEiGD
oFdzlQlOiKVXwfiYSylOk2EwsQbuwIJuyPp0zgVpzTV4pzhNPw+xf/ScvLPnwMqb
jJZjhyP8EE1XLvRh4VCLxNKBVR7Sy+SI5qUBwvnXkh1FcvJ/KqlXb1Fg3hxb3LUh
SrAcqz1sci4QbhLb1LjZl1VN+XNWPCgMNtwmhIC300RTZk9plrPXsnvE4EyCw7Gi
L+b+XBcGnVpMGIutUQg9H039NWGwkwtgE3fZMjDa2Rodz/AFdphK1A2JmyLLCA7o
JXp3gr22TcgpQCiToZ9LX+vh84apbrbrzv1yA4c2jySRZ1vNTRn9ebEZb2IviZPh
9cR8cXwE3u1t+zo5l2t0Qy6TxNFBlHqne99zOVIY/qG/2JxQlfu4uo11fz0qUVwA
QqDDoqAvRMjPcSr4m5OQ555fsSVgoqjThQZxd12wLr5idBIRmrz7szXK3G73h9mq
ngQBCksyBLHMzd5XFxZuQ6417Bi6LK0C62A1Y5Lmd7gfwPDSh2LFM/mHGwLPkr7k
6yKLAMSaQ9eNXhobJED9oUpwW2KFzy053ZRYeaOlyve3C6HfOKaUWGjU4QCIqjjV
DL3pNgBxOWMpfBQ2ZuirdXxGJDp/hMC9KYA3C+IEbf/P4iGesixWFvJIxEHe2mle
/ektnI/HqtsJxi0gA94FrlEojuKWAEMUJKPD5ztdGMdNb+Jgmw8+6JLuhuhQNA1J
TqQR2yQTxReVmMvzW85xOfwXAiwTyP4qE6kNu+QkKxVH+l/CudZAsysszN063+Ef
WU5WL/NkcjxZ+jAP/D5swc61ezEMALx1VYzhyExcli5bDuW+qAkbvjLQfpRWfz/5
IMEaxgBWBGu6SiumnxSfvHDS61LPB02389kh4gabUhH/HJ8V2IlJyEN3olgFwb1Y
PIQBhjOGoHzjhi7I4Uv4X3TkPtpS899WUJqmSelj2LsWAHjldyAbo5+dBp2MC5CD
oDQDHbk5Q5hZ+ovRw0Tcmlq3RRr1UqSY6jI0FS/GiFJjwvmbZU1nRYeshDpz1MT/
9LBpsRTVaDCzI6tNWHjn9klmVGvKy8lVwqYg5ihfgozLLioq2wfp2IWH1wd9+roO
HM+NloEnyzxyWyo1JMBYRZXOd43FtDaADr3G1FiQDCvEUSBqEbjSt2oKUuxNKPzf
oNjeX6L1WYgVP/EX4gS9nOt6TyKuxAVYwTCqT6wVxMcB5x1UjmVjEfR7gjqUmGo7
sHAOzB890BKIvJsJaj6BJouQ2EWOMoShfCdxy5A88kewT97RYuhYCTvZczzlL0hl
S/sbGtDZbGdVnxSAXFZXanG88WLs3rcy7xlpzaBc+x/m45sBhwHXjOnqOhAzkI+s
bM3Kts2xER50+FOitFBWXcAWnyeTLuUmBlPATasoLORkHZiPJBjPmCLm9FzM4a0e
w+lMjsP7B4wW3chPp+MSMBrXqnzzgCb2NNVJjlJhsuUhtXZsj/b2z+PmAcNVD2HT
6WDjth57ydB7AX1DLjjlFLkVtPxijCTVPowIb53lTOpmfyuw2c9ztrlbxgJ87zTY
fwPtq8nGkoxZ1U1mfN2dJbd5V6OgfPCCZXS7QgHJ55AdwtkpCSALCPiH0SiyPpIh
he9DAxbmBZ43MXUlC1LJjfEpZA8dzVvvkUasnDFYQnvfLBAm8RBSSq2+6AtZ/kxQ
f6cktDyhVivzWo8YgyUjQf5Rkgt3AOeG2srr3arpuqrIJ1eGX+sszy2zWmAV7QJ6
6NQA138mHsCEkmD4vA620B8kxRIp2fJxyVADGr2MlMtV6HPIp2tE5nSTKqLdckHI
bXzaIvtEbdR3EJa3+HH2GsC/oFByUQr3rvR96cepiMD6i/RiyoFT0AovWKPn6/1b
BGZpy/NYgnbGpEAwu1Zt+CtsI5+aF4v81Y1z6oTecPZGmAvoOYQZmXYkwzZc9Hcn
gq5AyzNJGAOxOcmSiYxZLoflBiPgQPubEatHjo6S4RSyhzhbAjDRmq8UE+yscc/Z
mq9AT7R1Sla4VHp0kB/WpbetL7yp3seCBkI9JtB7mV7bFFWHuW1lsseeBWhttOrC
agNZMfXN15pnZMDHos+i0a9s/SO3z5hoAI4nrQlNsO8abEOJkeNy9DWbXWe7zb5o
gCLuE1yulaqDR6x0M6ZADk3raLPUyeH0ld4Wjp3GlAB/mx6VT6vrMQphQb+GzAM9
9Rzr7Lfrq0qL2fXgq40ube4eORF+hYUjhMT6q1saR3Em6yKLwhP97ETOyln4R429
q9hA5ZYqIprzUtZmxYa7SkjP/PsTuKoGH6DT6m3+d0u8ZI/jsEG+OLE7Zo97itDo
oIt23I/H1qO2RG5HWMt6AhVFwRG8LndYvOIpXFaLcl/+nsK5RBvqQc923G1uLOC/
VcZ221fwyjKioopSJY46JW5je5Zw5sstfsKlDmdwZjCrAHddAY25jiNO1xOhYyzd
2OJBvebB/yon+JA9qb8//C5gXL1+PHhBkzMG7bTKBS/LljjdAU2ljyydK1bZeNwf
yqTRpkN/DlcHVD5Fou+CxgYOZUHwrY/VHgET9QnCM33DHfyh9lDhAg3kA9GVzCix
tRUHkh535fYkG+DFSW+HJ8Oin0WE3QtxUQRf1u9Kd3sKcliTzkEWRsOqJ/ivYUep
kEVAcZCpO12gxlcA7mJZ7DkDbRKT8/QC4hYn4UFVIZ2GXoDoeNgYQNI/9LkowC22
kYZlb31Z5g5XL2nuHUWiSsKqQ4BxKli87yvOYAPI7GHHc2qrvhqm3ZJhF9ByeY6B
7yKbQGn+BzajTATvNPh714xQRIJmIv7oqnxrHCB83xdInU1h0seujiFEb9KtLbgs
V3Uo24PlJDQGfKFg4IQJ2O/TqXSxJBC+1NWiRl+PLLep2EEFVLD3fpC1qa1MFVvF
5lH3kZme0FmqWptX5USDAlaVCiNQRKT2wfS9o97L+XMYID02nBvhPg1KVCX8SVCx
oMIB5h85WsT5M6bdCEJLLf+QPekfqMf3w6Ht7RUk+bBVCSeo9RVhXj+6FxciXcQZ
l++lwJ+Fqe2JPDcwv2zllp/22zPmqOdtO9Y16Hsgtw3pjVAzQfxwK/Pfm4+h9tIO
kLwOLKpy0Pr5/M6mmsc/wlLyHhcqfTeoOa9alB2D/1dVb3H1lRRmtNnXxbVp+xUn
lRjX3wcQGpEN1ObitVtVPJkKX7EO5tp5ENgwVJMrpYnHF63a/nDLkcs/Z/m2A9rR
D8M3bfkAqR5DVKixpYAL9sWk/YqJwFwzHgkmnzLYSTdFuc//JLPio3Fd02yFQzMn
771q2pTgZBWFsoNqyQ3pAsLicXPYgs3qEsH2olgljwLMDzQh9vE8EZHQJd8ihnSs
lMoctNhIrITpZd6VFUT25JsnOMO/7/cuicBhJEBw7005+q5BnkCmnmWu/mhsGckn
lhGLoSOPUKwHFIFIT6zH9NxLmsykuBU9WjQHzAxotpoqd3Wf2gMxapaglEMBJ/K7
q70Ota1tioZ/uMbSkdjmdyD/zX8sqFU08biTfjEst0O1Y3QzZj+o2FUoniQekL4G
mUAPs/zd0s8jG0zUpF7n2/pmyq3vYArs/rPCj0+3XZxvvH8V1DmYfkGQ/dt9hzVj
tYwrd7vfBEtqDxokW7A8iS/WB5ewIbYhUBs//uo7++6mGGwBNeHxy/CJ516m4/Ti
dE87PVCD1L59hTSDW6HWKJe3VhjsmqWJdoN9DTWuZqi9uep3rMkrc1LHh3/WbdRK
5KIXulNAECgoiKyiEb/W41SBpvfa1oIpN0woi+DrG4dBpal8iamRHk9Ch8ZHYyjB
vhJKzyOJ64pgSlI15HRyh9nUwPDkTp0gPxErIuvXckonDzl4pQ3H8c93J8B7HOoj
XBTVdfwKq0r4rzfpfk+zSu8vfEqyjMNZKLAKWYRXBMS4X5ZnrbaWRgUyAZ4ut5w8
yNr3EH7R/ZrL/M9OWnUNeSu5LcTGJWhZe+8GYlMv1cPE22Iy4sBPhS6Q+hmWptCq
I4O9bsoFO2KI2qWgZX+aoIlxvB5PUNt/Y0sZmFyzsbgi3FZR6+YdjXO5R7lk3/pL
eGsjQjvCMC2VUDUCr+xIMOwt4bANQZun1to/pL251R3+pqM8ieHZkbEXYW2KDn96
xWxc3xsz32XNYthOZY56zYkIlA0hukHpi50R7zgUIXeAqt4xo2YEwf7cLbVfA0ju
Anc99vvkQcjtSL483RRt8naDd3xcVuIGjHMEDiIJHp4d49Md6nF2XzoyyxNuDTD+
NfE4dve3q144fV7PZ4BXfZ4rnwIwZ0HPVqi3cebJKMKqp0dIe9fwhlErgPrD7vQO
dyfUBnthxe4ObeDCVgjQANiXTNGYREQjpOaLbu400UNM+h1LnG3XBYYSHkxUYZkj
zKZGQ4ZqqLcvnlTsc0cEn7ebU8Qua/fsLCQC8O46a5m+yoP8Upeoaorku7Af8vW9
qMhF7cZPO1A4QH3V7Sl2U9B0ScHGXMGek9qRis51E+3GO16QTig97pvg/ZPajtB4
JR03uMD1zFqdeZFYrgNjG22b3ez9fIhXVt9+pIIpR6Q++GchyxmN+2c3O3niinOy
bxxLlUHsWbNnprabEvSZdD9BkH3hYjiYY+5JZdDjwVXZytRS1i9SdBtnmSqTf2qf
zZT0aNvz777iq8aMPDZAfgyWdzxHX6Y6pzOwz1Om6wUfL1PfrxIXzfGL7Rxf3sVZ
aG0sWTFU+UHMugBuCjzNYjocW+T3nm9wO91FZ+W1GwS4cZsuDF7BOQjxIrcirwVx
gSrbk5ACRFEVS2eMLPBdfhJgqwwstvjqHHhN0v1vmsa9N4DyEgH3510Ox5I/0Vam
bfoXiLZRVzd8vkaeWoKq/Y86ESUUBEWSsCJ5jV4HqJl7PIb953jv1GmGyqxsuqA3
b06Tw+QpN3Q+ekBZRyJx7FOrYFLqhRSwdO9Um4xH5PYnW86WE0Ceeujjho2eZuaU
35FjTUzLtUSyyMvTC4JRPxiwR1F7acMToAcw/+hyOsqZN17Ejn8OT/7KyMzMztt/
YZ93JmBEyPt1LCRF3qIEEgghnPekB9xK0YpmZ8gX02HgfNeEDJ+mGJbI2JEQz9Oq
gtL/z9lyDheRiF3iB5O+D073IojSJxdrutTwN0yoTibDzA+Ur1GqYe8r3Du0rvsC
XTcMpYwW5OJ1UukRD7hMckHt8q2pPu9ed64DxIlElbqGASkDl3vhljxZp75bFOHK
9ihIT2fsm91h6r2ahZFBVQuajXmset1XWTcPP/EssXMC3V6ho2+2RMKge7Us2LsN
N1jlGBsg0aLsPN7mrN692DMKC7sIwcRh2HVysyKeyyP2x56PXT05Dyr7TmXmHVYC
c2dA2hzwwTd+A2SMV9tvlYFHOpgQPs3G71SJUgsrwutAKgCglpA9aUdsyC+nMyeD
+drIIL0meV/FuYMFfloVhwXBbbVN4H0KsTALZ57uphty1SNWuoqM8DF7QDZe8Dre
5cg/I8Adur3mAOdX0JzbnNQHpNrHzsC5AGaXv3w0osBCTJ4kouGe4Q1bYvMlsr0w
s48POY8w8MaNPJJrjb1dBEOuqT4PHBdogvIPEwBMqWxajxWFunFk/VkuurrwgnDJ
k4dlQIrEAvwrq8l3Oxtyk8Yd16P85vFxHuLmQyTLsI4zym9xWzIxbMAHVRilprSe
cxS9VMhug79K0uz+lMELnP05Ww8Jj7DecH1+5rKein7qkagNhlakE9XlhvpV0yRA
T5ESZwS990G17Z03V8QNKB3KOICxEH8RgvlsJfY5p06j0zfdrl95UzAY1TjifXZ5
Po1M7dePOWm6tIoDn5QvmwmksweeHjW3uVCVZTcyDv/8K9Mr+UrbCrKEt/7hQGKh
JTxn6Aeuw/mrP4olRoCSArVJb6hJCLejw2y1QmJ4Xtkvjarl+HvRQWgMPiqFI1VJ
3JEy85HGfYjK1wXglx2Bm6sEbFDLVVR6ZAE6Pdwh8RiKhFfVzo5eDJqJ1b25frdg
wKQAOha363yj9ooUFDbpg1ToaCf1vGqmNPtGFB6POVIaOOiQqcaY0Pr5QO7Acq3t
2cqnfSpqgdkC3/zBHWDd6xxzsn6vyo+gx9izIdkwsqiI0ucCiiKBJ2jpnD8dPQQY
XTgYeCIpssPg4NdXIlRQuyaPLlBs6CFHYko7co+0g0yM0+4q1+NOn4Q5rRFrF2Sg
4zCbJ1GmUGM/OTtYDr3hbKtuw5KXYMMW2s4YDR0vcnERWOqNSnMzD9CuHtYdsH/0
VFTUp32ytk56nQSt8w+6wz8+ZXYYoammTCGfE9DHqibcDAp9i5bOC7MOaEsHP5u5
zKEzvl2zqEDIm7vAVyKnREabM9gCqxUr7uckQUYtaxvMMZSX6bVSsXyLlPUdosRj
4s1sI46vFlgZg6rbhnN1XFb5L9ycgzVmam1BEKoqe3XprpNm425wCrgs6zDW0yko
hJRJdaIYjRqFMYx48mmaFlHAon5cHojhnb5naK0N4OxkkDj2DtgPrvB4Ul53/JgN
KumfN/DbAvsZ+MLiSgTja7HJeJyGs0BfKDfl8N1KhcAErknsNVc7OKTN/F/Z5onB
PKv8/iJK1Z47Pjv8GlF7nDBDomuMSm+e3dTS3SdL2Mtoc9cI6oJpoaKyigYnsEjZ
+5QESHZyZebJhnai6Voe+Hk/nT0mhgTCwIQqYuaM7OCxeGFNetBGf9cHIekdNzWu
1P5OVlI2AO0EHeXhB7uAlouKHvwulSwwc2JHTv3pIxU6owPJ7BAlZL8KdxY2zJz0
S2YWO0uxfpoTwNCY/7hIKlImFrsK4OSOzpNm9wKysugL1tlbG2u0K9Lg6QPUn2Bg
iY6rMxkb2YOO/gPYb4rB//RHZXcy5tpDCq2GrQP9LpDKnocI23RhNmRDaP/sWNB7
XozZ1S/Zw06XlwAMtNKEnHUBL6qZ/MNVYAz9IZTkdUJrqVibvwuQB0KiMogMRCf3
FJ7wxzTn6W62pCVDAW8NtCTw5Q6XDP9N1RBmamITTb6aD6ox9Ky6OHNPg4yU2IGf
iPBXIMSzOaPbE/o6WLnQp6RtZXykgm9DBZ1R0li0wMWd7puodG1yYVii/uzS0yFF
UIwNiVPAyaxkYcz3bL5CHrjI47i7hto1QHr8IFVtrXoFkADru4BiQ/Gcs//JiHmD
iQj/fl4f4V54b38XvFjHxP2s/kGzl/616PAdsOQSpsMNcKF7Fe9TnG8EegQ3lGa9
SMJstNceSyZW8yszdbLfocbVqkx47jXUWqdw94d0AYd/Rdce1vjoH3sU1MUHUmsv
2zs0Npd0FjMXC6kMvnUshTXkQocAQQJ5fHcnixYfvj0T71HAapflOswg0Oo1TA5I
DpHP5ULAtFu6uoySrg44QBFuxtI6rUeOcXZXpbQhNv1RKKf1eApWFTvTGu9w1Xgc
B0QdpXzSmxwdvfrszZTgMKoeHHh1TLYpsh42fwxDTPxj0goK90TYPAR3czTVuQUS
EZA4ovqlgaMmXABgp4rCcw74N4xfOTjrINRRnVAg2Ymp5a0nw3yQDztdvOIiMmfc
q7q5cH8fytxrtipJUwCiKnc7nu3Z7Me2CBr8M3qq6CrYqB7s3+REV08d2LT/SmKj
8m/6ZihWlEbAp5SawLMsjByzAHL3u7V9H/T+7hJfNgKBJJtGuRcAjSi2zOItvTSH
7KLc7FnxvI4okpk29KgyUj/88B28CNNoy0LNz6P/64XcO7Ej+LJqn36y7600LqSj
PupuWypSDF5DR19kqshSNyG5rl6aG8NcYvbhw9UmDS69s+xH8J8q0eihX+SiY9N+
yA1krEjlovxHFpgyTeTvaC1CkfWvdPQCOsK3GeOvf+ayprJHOHammJitwopxMVZM
a83gvEqG/Xdx92Ka3mbX21x514gxkpSkEWz0nQoWFrDT28bfO44hzK3uDlVA5hXA
WJlAdKXczCWETDmA5Z8ZyeiA6Xv4py1S6I9NdYZgAEcTeRhzrvGnDjvCyUv83k+U
d6i3403yJ1gfoMB0vY6s97/LExV/iEcEwvPjUvoGFWKqron9AblNkw+eEcB45/94
O2r+jKjus+AWaGE0x+fk5kTKVUyjzPYS9HbnjF83hvkfkiZkI+MrUvHqEmLP/DRp
q2ql3JtKNk14IEjKkOQLS8RQYqeYfR+i2nb7viaeHgjIjwRbOmf5xm72UDg/ms+I
xp1RC8tVYzexUnJ8T6v/n7C8R9eH9bJ4sgR+YWW9H864i5Pg6/xFF0xGy1482bON
CSoWmrTpvtnc384/BRNAR77x+5oSzkTvQ7OdBuRi0Jnn2a4wd3Rv2Y7SNFlbqBKY
prC44b6RWJ2VqOKfC4hq88RqVCBB+jUgYtAu5JpG1xxfiVqJx1W0NTsoW+DnHGSI
sWwFJ8sss1UMre5npAeIQPZ/tubcexny2fDOc/PaIsTr6AiLXicnqGWtNTHBaQeD
8qPymeMA1AuKGcEEl8iu+HsDdYxDYu/Bk+OtMjzDKqFepEjEoFfTcCCh7RiK0vyf
faueuDVBWi+sZK0eiWL0gadRA95yxXefApRpY4vX8NMJwkU+IUiFaH0M72z6RB1J
UHMaUMtvngbaGbgTLgorQvWfMK64zL+c44C32FlyxS7zHdzmOgYS03+CFSVLsnlM
wJjC0Y6BghmaqT6U1fvfTfghNUD+00WL8LGcIe52NTFVw1Y+2uL8ganJWHudO6/9
FT9jvijJ2Ci2Yr68BpxpKljzkwn/16hanSTcO/eCvJtCHwFynHhGZcW6MuVOHCSI
o9jadTe1TbZeAE4k3Kgdm4ZMRXF4amBXrcj6MuklQTPgF2t3SySf5YUuPU7hLHIT
sSBU9xc4B2eBChPshpYksyysar3cmlKbSuzY6bblJ+jbltNUzuJaLIVRyM63TDtT
tyHwVIvBK0W3XBO2TVeUtfgO0PKRQlcrFX3SK+ViZJJit3QlMxYEW26PIuyObZec
rD28vkZAN3gToZVNITZWS2pe2LpjMsFG2HI1RCEIFcTH0Ytv+7NFPf5sp7Wh7b5c
x7quEvOUBs3weA50I8TC6MPmCgyQvAJHoKOrXZIQ8czePetQwVYZg7LJ/Lee/bse
fpHr8y6LYRxCDsGlwf8BklKv5KtxMKl7o9+viFy8W60wqStxjbUF7/yOq4blzavW
53YLC2A/44G453blV1yx1c/5Ft7EyAml08BHz3vzgt+fak0bQ//jJpdE+7XUQlrN
FE4B6UoBFsCAeIS8E7ZaqQ+Uvx5Jx6xZgiJGXeQ0XDq3fQkTfBaEy1QNnXYmvBr5
vpnRekpYgDEpI8xIP+AKXEJrCCXb6IAWvRm9I/n5D/3EkrMBT3iIYMUEDf5YuAl0
G223i/Edc8mqFSjvdkwEXT5NR2MZ4kARaCo0GfCunu2AdTBGS8tQ8a8MN2fSDTzH
DXP2j5JBRiZlux2Y2ayW6lYXuEHlKY6tBNE5UEE4LpmjdVdUVXUxPUhtI1AXXkRx
CRxdcSZRwJeJom8Ue6zfdmXawUXfxCNHNOIOZ/H/859hlI9r22VYB3FHNwyOBg/g
4hg8rfFdXH/hqTm/AQB4GViXY/I6UCCzkVzGi0aQa7PppQHK5KwQQh4YlxTu0K8U
qIjPomHE6fc6+9Op1FsOPZDq+w3iGdjSd4qV/wr2mBpM2NWEogenTQfXG8GBEo7Y
I/8FT6FrlzKDWbVB2zEljEmcK9+yKhPfALlY7fclgqvmo9p5cHm2rssTbo77HDy/
Zji9lIR6yprFSk/4YyqNvj+0qwkV+/HqF4JbmQumHA4g+ofLBhBENwJAIzf8r9T0
0QFJBCZUHqElS9xNqP9/8V1+EquiGEIwIF+zFdEX1EgSyaVm+iseacRE4agVQ3rw
sVKgsSoI4eooCAqZAID93AT5k5FbekgUOUlS1kQ+uZhj1yQXNu9vLb4tsVDlhPA5
hck8oJ24mENw3loddodvIUfOl4tWA8lKE2Xahbz+Q0etd4KcpkjgJC22/RdWfpDK
w2TJpF2f8vO2FaJqGSMofxbWLt9gt7I/hj7mTeO0RKjJftJXViDgGc3ZPlx4Ss3K
nLhO4a1zWhNBmkNWs1iXmmCMF23HBU+0E3iwIs2hylcis8/hIqziY/xi63bGW+/F
UT1Ap951zrQapAr8LTgweZl4V8XbR4fp83iYfoWZ7AGmSPuD0t1i53UFTtZ0y9K9
5/R42q9tpGp/BiPQayfddgR47V110XYsLL03elRAM1Ercit3Y+fIbaYcire4rVIW
2C9adsyN67IspjEOV8Ag8mOYkf1wPeqAOIp3e28xejswn21RqJDHJRV5Vz8xf81h
a0sM8XtUnDobOTXBEXTb5lE89tT0hFmzbdEuEcjv1BUQoc9+ZruSEfqTZwSbbHHl
jIqKHrT4jCKhaFNwkv0+3ap/xKQfS5a1CzFh/X6d0Ecu6+M/Zohw6oPMAuatIMog
aLU045TXJrBWM2088ikZiE0ruzx2J/Qk5T5RXqAhplr1Kc0G2Npldy4zJCs7TyI0
a/0jwz6E8CFA9Prb72hL48z3YhnasdrRDlkGZUjb0hpMcOIv82EQlpFYDcU6yQiK
/gIIe+yUqXMsxZ4nM0IOWHaOGbcxJxh1hWF6thiPfKZ/krCLtU8HumqLL3ssm6HG
AoruTH14wIoVji4o0M/lN9/KyqGkeAyGoaXwzy4XWUdxMPOSifDWg1WbF1eCE0Ml
iSHyUGgxv+P42aEN4dCJTUvD0hR7VZ1Ku//o7LqCWLsDoPnkYEePmpEGWeocyA6t
Py/6KQxNOe8smQ6U15epGhkNbuADW2R3TKqHmWtVjXHCVdS9d+V51wwBhnNVWqGo
RCWO38Cetrag2/nAaT9XWJZoByhQhIwozGYv2Yf7R3HdDnF/dL4anrbXfxcyjx24
s1kGs61IOfGhtklI314h0Br2Qj2ObskJWMk3YPn79vIqbJReROKdYa45qzWHlqo7
L7mZJAx0eYfFHDWxY8WpmS23cidKciyCX+LZSyNEV9a9g7fOttsHPxZSGcoDK8k1
weA4eGFwX2la83YaNzye1BE+j/lvEkjwTj3lxtJebJY3LFkYv4sP4aaIpasp+Z8N
za1j8M2mRCwPL6S2tqLkte2lfUMBHkNSiPBFSH89fj/MaJ+1WlRSGtpKb8LRBx+f
iqJPlp/6DFtJd0oXZqMe2CpGcN5RXmoqWDvh4LkHuUJSTs0vUJlACHWPjsN6Mcj2
sl1iBLXZLa21FuwB7FLNGmhIeQJO3BesEUYU5wp/oa9FwW/Ruubnd0lvVb+VtMyq
0sCY71LeICjBhvXE42gHFDnspG8kCFdpLMASR1iFUc+XztEEDrvzPS4LE+lm9bWD
IF96T1m5EsgcsNBVPZJGNSTe1Hwt38cC6Pf0q3kHgt+lv9ib2s1RGe3IsoP1dN3z
MFYBw5eOrtYq2feAJzUT+IvU6GrMGMR7CscV5mcR5PU7EILnX70Mo/g20qqLC+AF
SKew36PQS1GtYW4F3UvOqBd9M/darXSejQGDPNubI/MPSCUZf2lS7f1ILfO5lF5Z
wCTPw+TRMHFrZ8du06WxlBzfVDsdVTN9N9DuLFLijwqizUPxrUJHCNsGYRgHdU78
zihJMH3XaaLrp+3N36EkDNSx/Iu71zqdfP/DSJQkF6xBjje/YucSmIip9f/b7RSw
Gbg9YPM+1T9UpqXczWTcE5F0lXEehS8gFw1Zd8v+WWXzFxHV4VXJQpggGGKN1Iq8
ndkvZT+yd7jK6WYE7C/sZToiQ35xzlSQ1CNxe9qnusUAAbQOW8NzLiCf1MgWMZrB
bYCYjq/ovW/UeK73YRhC9SoN4b2JXJ3BtcgXQi1ArqYJOcrj1955zWX9tvrxhjmY
9xO+Lj6dzSvXG2sgKfSsHsPuyby+F6wZeqLq6bw0ylRHDQnETDrT195UDkhZprIy
bZkQSFkWtdJ9bvE91M4TErepKLzWlmcstbWFOJHu1VCMLdaOFNCcoGBaqi62Auuc
KXVkqyotdRXcbGoxq+GoxyzME76HUIRSQbx/8q1PpmvHOncPieLItiT9uLI6fHgf
pTcyRDJucrsMGvYUZS3Ym3w5ijaL1pkNKdFaMswfzx3UiY5viTadQcjoO8IKnVtF
k9v7SUHMTQtLYjLzDu2PhhJMOlojS3p++oC84EmarhpmFpGUdzqhxw415ZIn3ydt
B33EyQixCQ3QuCbNuDDhEujc4KRJBxyyR4YCWgMH1GW46Z62P+2IEEUYTDUBzKx1
28+leCDRRFopLYPWGsuayuwzaEHa5opODUNG6JBFP5MDYvMK1TJ28Qo9ynW7rg5s
ImbX/SajAsYBc0sMQ0KirXA/O9unnSQoAIM0tCeZ+T8NogAJaO4if2+GZbCHwr3M
yxDf0sUwJ//84DZClusNmgVYu6w0xyKslOllwCIzmK/+8bqQs0nn51+kZTw0V+PK
oZmqIQ2za3DZRk+kjAnFwnmkvjWS6VXOTS26jUd1VLdG1xJTCmG4VxdXzQcOrcCA
BHG0Nl2rfh1QFgfEMYAuADnZQm0IZkA9W1Tdg2o2b4Sv7YwU+laffBLrJwUjXQd/
dGKF9njFaCytCrs7QeeBSd/YkTEIBz+D+/knoOVd+SIGJXsxnXV8RXPqWOdyMDwr
F84A4UxDwyZWj/l/Gu/lZpVZDuUCVSmepwHhHLv01nQPjW3VrxxvTVZ5NwMa6f/x
PTTxE8ACjAHeFzdFZQ0CXx8mL1D2dzeaoKvEY15Y7CYZ0J+CRpDuGUgnbiYMdw16
Iy2sZ4gGhWV6IXUYcIe3UfxhhvYwTxZ7eD4gZkQbXspbXAXtOlfdRYdgzkUUgN8h
ZDrW39qdjiQ8mmrwA7Qhyg9WmLvsll8Dtr4wItu+VTLbnR3WOd+N/ILHCDoHhdVe
8WmIrwrKTSKGsmoQnESsWpz1j7PV1NjbXHJtMX1C+ve+aBxEuMAWP0/3d5F1+2fE
iIyKDFMcKJnMpDZ9y7R3u/lF+IzNdhTdARyDQgvn5swzNS6YcwekSCdy14ZvO3tz
P7OcK4Puuft/ls/Ddk+10SEK+xJIuIPK/049xPltMkY+IixwCs4WsTEUfHd21CyJ
HGMh/ZwItxStm1rahL6nRhPy1gWk+Wvdd7+qhwVO14IBpyxtoEkv5UFED/ogAN5F
e9aYGQ1QCS8P0JwzTzZy+I1l7UChF0qni7VffNWtkO459na0TuYLqe6sJVKq+Nfr
1dMMeHJDt5P0xnTMU5eSGxGFHXkl0XNZmQE0lVbGzLR7q6eRRj8hBHuPqL/zZySc
4f0QSXKJ3GIErZ/d2LE+U2XgKe1Yt0nZhpcDMw+N2v+1U7SVBphj//HuohyrXNb9
0HNFYtRRAJ28CdqKZLSgHtqN3qne7UDfBHaGLATRZmb/POJf7/qCGZUpou5J4ucB
sSs3bqbwsjqVuPrgTjhyR9FBqpSyCWZBr4Zv7yPLNGQtgQkzoIXqXFS6yhX+9SzE
x9VhEcSUEOQuPDAKiWrZlS9XX10bNGpk5lqmTUDddJaoJ+hCLIH0Jk/W7OSZEKhL
+NfEKdQoa6L3CBzIE2WPQomLSfEaZc8nFABX3RRr44h2kWIWEf7GRBOCM6Xavgji
pWMNpVJyOgzJgAu332kLKV55EdUlJTXXJW6tjKHHD6erfyk7KJBxNSj9Xwim8gOM
NuiZupnOj3quk/ZmgAGLLng9clpAFiMgt9YY5VM2CXFcuye+s+e/yyRkGEtAXStw
weapG85Iu/OHTiTM1XAulf/qW5K6ybw58Q1W40l7a8NrohdmKi6hdKnWotSELTuE
1HDzLDokRUN7XNvsds5c2AK7Ee27Ec4uphlSceD7xZEvmNDZ6LzC+2qVRJj5bG6p
ITWZN4ho5u5K8zAm0daHYHZ0027DVnrXeODyTqTutU469+lsJ4NgPDmxWTzd++ol
v86AI/c/3OuNM/Er5EPrYAtl9bUeNte0boGtIJNtBrxCBLo+s7PbG6qL0zmsAF7k
ttCepHNOOVvREcO3P0Cu63tKFPSa3+gWj3PEMmq1AUyxjZpz+DRkNd7a+Ildvg1h
ZzqOAZXHjDzI+FfUGHr/s/72v3MwdEOJ4VQU7hMRSFusqWoSVVC1+ZQFezEbOn4H
1tb4L4B5mHN3PFhEvXVlG2hB/W6EbYRX28rl14KZcBUVGqu1oEBAB9YpuTnmkv+f
5iQLAVim7M7znRT+rfEInbqGTw7KJlbBlbkyK77A2rUcWZKDWwq9O84novO86+Zv
WFa8vCr3pHbK3gi8ufmNRh9jdV+1NffqjdUhEb580xygkCx6kmGEDHG0AwsHhlLp
aFyEckUlrNxl5zwq8Jk5MGHbnLeB6ZmVO+pLn7xGkDCnniHjZqz+5tEMql7q4mCv
6UnKq1YBDaMy7lM0kVqIix/cuqA0dJVAI4FDn3BjGA+iBJRfD1naD2JdrAwTVRjy
QwXdRqB7+7nbst/wJXEMuTRMvfP8kyjxEEc9HKdbFBTpqxXRKQApRGpKp51iUGnK
/bZ2pFrvwJ/ntT82OKeShLcZbGrAl2MZ8i3YKNVbWH6TkipRPXCVvk+YS/sr4bzf
tnWDYx+zwyjGLvnKI/gpcdFlAMfgDa026Uju3jgCW92T1NhNwD54S95hv1dyAsJl
D3TcBuYXMcIg6GBLpTEdyWJJLCz3l3ynYg7kE3Vw25Ck13LJpxaqwUHthu2c8GpX
NhX5A52kqJHLWbfsbfjwDFv3MAByeY6Hd1sWcIWN1PcpGHEtbXbUVAZQNcrHpQlc
SO2RX6xR68/sGFTz6z7eU4heun11zwT9USbi/GZPvG5itHCnWRQBHQKnHOQT+uaV
+2B8QTTxZex+x4s2J0o+LSnY14UcSytsopGh8KQS/kiN9LRHsS3qoE7QL4h95/4V
n/mGOFQHJNbP512O57LcrkMo/1y/VU1hL9jdvBPLaoDuawRHFM93AXkiATiBPwul
oZHwH+jsmJAKfUwNdo5QFnJjk4D0X0YNv11j2A+0MKLJgpfZzLH9nu+5Sedim/jR
wb+nYTHkCD9hjlvKIHEi8i19RhC5ypkXVxOQY533wJsQqX+BF0HrIreMZmlNsW3u
QLsMKsJVdd/MZWQl/aOUg3mrjKB/ZkghBNPHVy795l3WXrJQzCd5nU+DHS0omogC
hvFIDYRifjLa0Tj/yqVUrmmFFFv8uIe5IYqSkWN9ynIP4fwybm7dBPtoOHCyazfU
cLvn10xwOIwapTANI2DtLyZ2ekWVz6sxRkYq/zJnP1yhLs/bT8P/fQwB295KjuQH
1Hc5bcyg6Wg9/j7/Qu4QG/6BwjditEZdH8U3vZszaGJC83D0pdHPWWs878g2HGRI
zarrtMK/TVDnDX2MVigpbvpKxeDthn1mKJYp4eo5Z5f+5/+hyJMRlAGKd3/Wjd/E
TZTkVg0p6iNRt1WbgC0W0yfFfVY0hWC7aXykd7zbr/GilXR++v8fXObCEx8GMg6Y
OFNREgsgxRsWIUdRngqqnoYR1wEgjnbJ4Rsip5mLgFqfrhyGRkamfVeBDb9ubCoe
qnbfMsSC8CAD9ajOl4a2pgN6oiNU6X00c3qtefstVK2WqosWxbvWkmeSoehNfbKg
oQGN3ckY9Lt0d33InWJpcuDrUU8kUm9M3bfQeKp31dfwlvo5jYsX/c0wnhbWmBkw
Nj+Fn8N5j79opDDN3rWJ7vHbMBbWBxvccTb8uCNf6SU7HxytFkJIYRea8/RNlvHY
UCB9Zvc0Uo8zT29nJ4MxiKy5zNW5E8F9P8tmH+lEnzNWqvwitT4S1BVKMU+M12wd
xd5gT05/hs1HI+gEor4ch6Gs04vXxiMa2z/6XkRw9MVuYDv3INTxoEGxqg34fGbR
JcpFnPbw7dvybaGZTdwLhcn9yCPxfY0TMje4IByT3Fx+xgs5Xp/SdjyLG9eQOCtr
O5lUG2C0fYrneosdZgHGF2NcR/rEMcDzcgRMP3Puulh1bDPdLtoaHV/1PtmpSjT+
09pyj9xjpFulEd6lcWki8lYlhzHSSuaaW7LCJ5uEm/kxvHf1KJXJgGvuWrxfvplh
NhXWZaKKIgHftv1mek5XluWw9MuN9xVQ8QCrjllondW45GaYDDz7p/BVtOy0p5CB
3/1swU0xvcxOhbDVTykMlftV6NYLQj0RODtFX1TwUuPetCzV5iWGpKBSrPXK7o61
Q09XXnv4LCSD/QA8izDwh4h5amt2zBrv+3oQI2o7JMhNXyv7+xwbwBJz4nFlZNA3
d6jUhwpS6sLRh5E3UpU/TbPcGAx2WqYb+FlshVhme+i9M1uZTC6aTnRnJg9sxAVe
O2Z86VXmBqNiQmuTtQUK6vYj8fzLbI71E3+vjoR6Q7cnYxy6SBnxPYs9KjDh2GdU
6Q3GLxao/olP0VNjVIGJFIxuQ423hPOyBChta8kbS12mWpCVDnJySYFf+oFL40xt
gygiHNmEP/1yGIY1qduW76XLY+MqUMXxAy8N2MPOXKhMij/FKa4SQUQjO/ZbEONr
2ZK+O1TBVu3zgdD4vyNvQgt58U1VK8pXjdmc1Jr6DgE9gqILUBmCzZLBL5kpGk78
U3PWsBHVOmBR5TLIS3chAmuZ37mH9X7VbVdMhHyDLir887L8kyNkOx1lMHbMa6i8
YmJnX4X5KK1FMBhyWJ1Y924YB+Ztx+oL5Ct4272+ur03heXTjcrXu72znWanA14x
POKB4WrIV4vQCYoyG5hfFcgGeWQRFdtX3rXCPYuEGZUF/zfWzmLKVdVwYtcJOV2v
97GF1CeP6VcIHngSt3lysTXRlTvkJoUEubFl3kQSjyuxkXTH1bvIjMb+vRTwcCz/
jjh1Q5BIx72Cz3HsjTmIYEltx0/Hkr8oie9so3leW8yzWhrJ+KBd967jzseIAlLh
IPOXCA2YVNhizAo3SjScEC+HPhBbWTZuAPdY2MQrn2mR117VdJs2jA5fzJOw01cQ
LrBn3lPK+gl4ZCZyBbih7QC7VbtrtBVGnSoGAxc94Wo6BPdtyrWk+UZhqkooF9FH
rqgsk5v8Y6t+lZUAJpE0zwkiD6NX6wJPw8wTCNKyB7iy/LFStBqAfcEY1nr4nYO1
ws3HQcCdFUBEmbTfTiuqMJ+k3Ca+k9nOeSCLVQQmOyCAj3QM1QlRdjdsQtC2/tnw
8KE1IAS/z9CYvgpCYi1whnWDBcm6UwZOQkuAV1EQLbnsUIky0rvxkim5OJQD82cX
ok7f+wpqpw5cK/ecSFakPktliG+m6fTUOLHsB8IDoVL/DnVSDBuRAJgGH+vF0PSP
nijVYAg5eMf69F5pHfzqZM8dQnqyDmPE/zF2nYp4awOs26WkCzy9SLWRiLF+bgiL
5tTissTeAAhHsZcC870sgDM/79RvNETHfyf/R0NVp5zA1OpeT+tFxrHIAaZGKF4l
Rg/dawfiK3TEcEVhOPs7xNIrPRkpDzDinmlbPIkcIZa5LarxtPDFNdI6YmJiaW4a
lCuo1sKodArWCYA1UsKrf5gvwzvZ8yHYN83YwcbNFHwPU3lY7MEXehMXJXZVEKDR
96cJAitSlV+Zh64eNhnBt9lXmCAYB3risJuCpm4lx2EGpqo42aXMHzm6vjmNyqkf
tELH8UwQNyYtuRJ6/2uKaAvXjQh8GV2r3Vum7ntRWxKH/JRc2SbcaO8X0qY2t9JO
Bni8hkJBksduirL2vMruyPaLaE5lh8XHGV3nrgXJTzHVFvRVWLfaGYR2PljJi6DU
mdUVY0/Wa68jx9HN/z1bqFgzY0q2xNSz/wAXWKXBvsDFGuNOc4b8PYhXKHjlkfXm
8eddJ2gx2egeVBvOSDYjEGDxzRaZ3c+DIZbB22ruQwFM8xbt05ZtwKbqZAeE+5q2
uYNw1KBOWulVamFpaIZkdoWYTvl5KbipFSp2+d7xlgWB6PigGqvS3xo0VW98l7SI
cHY7Q4A15mEv+PQzxVmg15LNacWJNwqXhtTkW/0YqSpZxOex1ruxWJ0g7alfzSg6
cXn/a4OLZnD+3xHGVm1G6cgNNnB9KcVR7gUGcqjJRehS03Jjy2up8cvSf9Jrtp08
AYMTYd3zwom6xDEa3DzhkGVdI0G/qfbQbg+pb2r5InTUnqSAADW1hz4JRyP3X3mX
LlCFaXlKZ3t10WAmDsdpjaqhwXq3mS6sFopuAhrKJZEotJlIxTNl2z0k06JNodc1
ox1Ct6fBvvYVsBBh3L02YA/BlwLMp5fqmP43dzQEZMwJk0D6cT1vRbFpDb5sDnV7
ERldxsrhcxgP+jWGMmM9V1Uww4kTEbCUwQR6P3MAnznA+7geKyeOefqvbOHTKp75
Rmgp1e/C2rnPZ/astow42dJlEKzwn1LiUC/y3xg83fXar75LMolhGpKow8GSLSR1
zN34fsty4yiSSeKL2HfeZWaKZyLdH36vhr33MdRtfUnv07Gdy//XI7ODVoZlUB3z
8Q3IqJhyO6MFhe/fn28EBBYTQ+Aq83NGGondwii476ZlEEyYENn8nMTlWeFwlD5H
+sFFHrOniMqckVN+gamg3RrwbLb+I4qWkwXw8Afp5eoODOpIa1bwgZQrrZrX/849
QXxJ40HGI7iXGLuU9o6ayqcA1kZ87AWbSPOuyWawsTC87II9iN6dsShIkNG552OE
5pF4XMosKPy26O8wbjnp6mlC8PAzBNDoQR8ez+X0khYvjwh8EDcAru1M6sGh40wp
m2F/TY+xJFdlyMyn43OMdycO3wfAShAJ7XYdCHwhb69Mobsl9YTfikQg6DCqavot
sqtS/e11C+ljssJQEeniHLx8+rnkLu3F76GpmDtuznob5btbzGgEt6wZGPQpbo5X
iniI7mapl02ptiLnymN01spepglQfdXYL7RJbbrp1GC6mIw6y47yADusCsLgTjWZ
1DIKHYNwhfn+BT0P2eap1vlTxoYQgwI4KiJNUtFJwxp9geoGIQZgxrIKUm6vjECE
u3yyn0pD/+kp2u/+f/QtU0gCK/OIr2pMmAMYM+sPorZroKKiD2JlOVmLDeB4LQSI
vY1vStSLe0ENOOkC0xqKkPlTM50T5kiXb6XPBsnEPZbCRF8KKDDUcl0fCFPmT2+T
sb3NIzV1URIVqpPl7q7RQ22BKL1nZZGCAuqRZgJBCAHwivvWoFui7PgbjPSnfQ2B
jNbrm7koptE4pQPnj4zmPLmv7eiUGZMC4YVkKOfjl4aR3xL90qdmoBM9q6scpGgg
LxoUXv+gl6Y6lhz5wNFeewwdEKQrNmTDWrCHeUT0V2UOFaiXXhFZ9i+XPFLihSBS
spe+0MH0vwsVHCJ4JZT97PYrqLfzQgfNWzfo5Bir7kaaw52SFebp6Ud3Iuzvnmxk
mb6H07r7tuk4Gg/44fD5PmdKhyxgu3yzl5+xntpF8FdQOUfsMx942fjUAF2bnpss
JRnBdgEK+z8BX+zK3iQ/h1UBg8bDZucw+awDvZuCWVcHQw0/n+X0W9tblYbQ9uc2
lAu2kyfKpOCltuV6IHtiXSJJEq9T14cMMlolVKOV07CV9WVqPaSe7AvwrfFSSXPU
23gMyI5V6t7tHSVS/se2AQ+5mPYoCL5lEhzJ5Uz7LhYgeNKd1OwF3qS/lddK5oQZ
jtpW+BY4G8BVGC7o4kC72fS+ZafWtPr/VXxTaH2imXlan3H7Mx5X014PxqGsKF1t
T/K+28v8I52FPY9OZXDg03uKInOZHaj/C69u6/KgV9dr13vnvv1Dn8nZRwj7Lw1U
Q5+FhVVQtMdkMdezlAOtrOJ3EEXhPFMTxiv6E1RTqZD7+bd4UVGK2Wrpk2ygVBA2
mI0uIsdUJitXQMVVzMUMfwRUS0qGecxF3xNMuVDnJMCevfxtgPzvxLvyDAOKB8pE
bG301bb8jJ2DQIhNwmCpqNgJG0GybNnCOGIeDXG7AukCYXekSBS87az7959zRtEj
mwQMzBmWtaOufsPHA5nAj5u/19WiqrGU7uM03478k7B6l+i3iHjtCFP6ayyqO1Gk
qcwB91zjy74geNLg/Zt8LnRAd2SuBhyZDTV52IfGXM6+tn8y/ES8UhVQ4azZ8PYl
0pxS0SLM4aT3zWa7Hr8AbnDWdFGodEC72YrmsqBuF+wajEBVZrXkc3J0FJmPBLky
4hRU/R24sfwsYkp8y3ZZyhk+LS9EaQLAqdaqD/w4tzSh0GPAvHiAJ6p6ejrig2Je
yYOyihdCPfheeunyvsIGUoj6E9GQnIz6S/ePdpldRnMdjyKx3f4a/bVl6dX8bf/O
ujHlsIuhzSkQSqKMy3YO7kR2pGDesiBScvt8lhlEqd8qTAdnkdLAA78/0u7HEOuK
sx4rdfQTOjRt86hJvkxUWnnfr/ACDS1NwUnStJEkf8ULRIYs31iow82aTNtnXHxw
OU6WGwq53X7n8OimHK7wJdS3CQsehDqRFK7BsSISMQC160wEhfxdXVrr5nlOTquw
Y0yBotRRKsKOc9Q+lhzhJ0dxu1K9FgZvy7JYnmo7IlUGB+oTegCsmw1tUHaewh+V
4DMYIa2ePsgbChlsWfSa66/uxRx6P5fyvpjYAaZSKwRropkEqRGGX2jSItgjzgc/
89yxr4q3cI8uvkbf9p/mkeYuFSM2GDQpf828IT8Gowrz7x4I7mvo2lWNMm4SMRU9
5DqQnQGlyV71shGesEC7UjL89EbD6NvWRbwiShx0cpiZSGIdhRxzKJFqnD4ih+Y/
X3rFl/fv4QO5w4l9Fe/D6hgAgTimqX9qsHvRLRtglz15gPznzpXselmrQxw+SPzi
ZHHAVlr2SvRP/wHj5CP8wFq++67uKh7Dnife1EVL2/Orq/cPW0HYzEtEt/L784Kx
aVEOtY7KRzR6m64LDYgii97gxddn9rKQDmy4qO3hJpZTCaExLu9Ai00+HjTrStdg
9I5hjgltg/e6360QF+uVYumn8W2wl6DQSwCC5eZIuXOkdgfOtdaw4hI5PgbHlaBd
36y5uodd8stmOM5okbwuW6w9tPsJ72sj4KALCL+luRTDsRPN+46FwSBPa/ejYKVA
2F+Wfbzig/CW2oWdnvkfg6l1Z7tF/ZxRjeVd1tVcITjrjHmf7Ptta2/J3JkqE2yb
tqW7vGDJV0IqA+nlUjfEeKCniUo7tY/36WVKXR1m9noefhYnTxRZvX5FAJXgCcYh
3fKLp4Su3dlPhWAcqOisGyd3I8vQodDSj4+zXiEyQ1LmD8rMwP3MVT3PEBKwygmX
xV++xhI0/oJZlnqidxaeD+PKUru2pA3ScWRXIBTXETWVqth/iJnv2vSqcN932THf
waGZArA7bkuXwfznys1hdNvuNZ6YVSoDwDmRXOM9lBWgw+kzo3Bb5EgTq/g0cnSZ
rn172fR+92XxLmsie44zWaqWAQJ87EMTkpR0ZbmRm8R2+hjtl4LoqKxCLpSWEvtA
y3bJbAmtvT4Zk7rZNgUxD9DUiLbkVRjcEsv55k4Bs4RPIr+bzqqPLuNfbKLQ0/So
gTpxft5aEIyEFQRiUsspn/3yafKF5bIrKhDfy2kpMdGxkwmDZ9i8l45wiUtUfEFW
ofWlYjHpITvMFAbQJ/CztriJ0AHToZz+w3O1fdi14zm4Ve9qZCR650rNvMc4NjIQ
BNbJS+9L9dpyolVklF0vjJ+co358LpR4Yrp+Z/Lu1ZxsSPVJxOBvWBIVVJ0iemKw
4q5Xt4lg9r5QO7cJFtJ7FA+i+IcmqfFCTZMhJ068+hKKi5hlbVMt4ZcBaQvZryFM
Z6w/GTTh+waxqZnQzZGUXvB/3fIDXkBeOVMYEQxqtWpZY6TMbxY6GUwaV6xORFm7
VHj7WrgReFpZcEy6kclxhXbOmd+8TCwrBLdFB28cPM/mpYOdtPR3hAJVPJPR5PmT
k+HRcZjO6NsPrYeGh0jlcdd4d1rV62A8Cpofy3grskiW4hhQVBtJp9q9JyzaOmv5
n6LFkW6pA+vXpRMPHkxru/xkhadS2ATnJgT1apXv7SybEpT4zcUWs8Nt2hUEt7+z
UIvAWEmXoMmTrEb1MmErJEGwPp4oNvKA4e8X0zJ36JBszysf+EsylzF2xSXdHXyR
tJtT2TROqOBRsG5OoL9YtpShbCzYN32C+28JRBeFFurXhTv/lw/X6vE3oRM895/r
J5kHxOSSKtWg2THfmHJZ+DJQxUlLphSyn1R1nACb3iQDOYO9hOBl4ol6y1SKzfeq
IVTkc/7a3TOT3yMQc6sSNTHFIZa578IlGaWXXrMD3eCxniwDZ5OBAqmm53AA4eiL
+dErEPlCiL9CuuPEBA0T2s5vHaZDxxDSXEcSAmal1qnoNOB5V0ieFfpQLwN89bdV
kXjGaCNANU4eaQf/KWIyApr/uhlcDjnZOIEPljlwozyui3PbwyOThRqClaYoqyHP
JSWk9MSNIv6OQDUA8T61Hv9MfxsMOpFrncEVjNMcVmQ8gOYO48ph46ebMWUFve/2
DCR8uyYX4J4GTMSz3G0e5BMBGwSfQb0xs8C1SlVfSsmFRj+5QRo+3Yfs6258Xo6L
Il32yYC/6AG8pQC5AQVy0wg5JVaPSuUauvivb4f4mskKEaMaJ+LCFhGfofLgK844
JW2H7Prl8FlswSWipu7gDZJITGpDXGvqgJfaSUFI6kGLNwmiWIal851kD9VQEj5K
mpj6kjrSoOV+PXiN2pnjT1sBDTkOw4noMAONdNGxanRN3xgFjaci/NlreYVuUk2C
AUKUckfR/nIRznrThy/+L0vYnerOEh01bLEd1ct8YGtSYR2RddyMf86FdTJFWrZW
78TnZ0bA/lmmk15PmA6iVorSR/GDNXMZNLJgMJ8WfygypVfDqeYVIA4DWJasw0Zw
SMDjWrwlbORe5vvLh3ekH4bp2SEQJaKI6HjsLc17CZojklamkRgA7jOt6Zs0YOne
4tFVXccUVTQnuNjHtPNXAPwfzXMpQpluuwtiIk+nFsDZUidumQFpasFXuWC+bnQl
H73CQ9uM9pCFrHXDF5hd1iSeChstmp1V5Z+RMtQGzSYHN0q9CKdVX2RURAukTP6B
Hn70R3RNDwmO+AiPnkbwA8vKC2PBKFxplNm6BcgLMng9oKCOtzoQbRXLWcYkDZ/o
nEqMuvbNft8bmdCTtPAytTsLcjmjyOqkTylrcHJvaIjcPMTkl8WbzLGi6egraqbJ
0HngvNAkgCkW7w6jvFvXa+3nx6p7nitbWxLwBIKXdDrsjxsiccaY3CkXfryDcfC/
PeXmk63TOINWmc2tHZB3/BwYIOOGQXnlunQGM3uWve9l0KpbJevvnj6ugvelCdD6
Q6Pj8U0/c0ArP9xD3qekO93I5T9c7mZRI+WCRDJbRwemaW2CM//xt4AeGU2LxFHu
XHWs4ft4TBiKSB0xFS99wxRdgLtsI7YF8Cn+ij7J3x9bC5ejPji9nivJ052s/Hhv
CssgziZaq2LVaIZ4Oc0U1zFlEowpcUN3HeYoj9IEfoY3PLofUkx4KRLI2Si3tn70
OoOKwGBTuUxS+13shkJmO+nsrSwzok2rVI+aLJduEgyeuoAU2p6rHG8X4lsEkHAd
lk6zLIG1DQuEsXrNrjenTHwq3fndtQREbHgH+RHURX2LR2r2kM6aaCZIl+ICVXGC
sqwzsow39noy9tIX/CTcMAvIkaJQ6LCryFO1kH/gbcQlXeDMyWPu1Js7kJjPkGBT
rx7BGTPGSuEBOPhBLg5HQYRrgYa7vsjjBtN4ltNMgru77MQyPbsxBP585hgNdgp/
+oKaVrsYU66D/7d+JCNygOFvPdrSvsn3GSrSc0394hMVfrxfh5weqxcn2vLEfQRt
ev1TPYZzwnq0k+wqPjf3DBrmyiPlA8ZSWDcDn8xE4i3NjhQtI8O8T7jSKCpuMpK0
F78QI52KERsoWej16FQwzrFJcUCzFcs8DunSu/7TAiQ96sBZXpkK+VVLrjdy8Hg2
QITEzKMSwnfNz7lO6a+h0etlw9VIfkWY7Pmmjf1aDjyfa1r/IsvkmyDHC9e2VpXc
HO6q2QsWZq3ycnceANhDYh+pHqaDYlN4NZAf/+jFRamsFMQldXWUEE2zwEJHcf63
nQPhBRuADtOra4S5Do6ouCwJArZL3lvs121HcMz9V5JC90xWFCZ21z1vbD1F+iCZ
+FHQQb3jmcfZZ0bRmWnXr9+Lj8gog549ENYugooUYB1Df6OyqFh2hxqwQqprcSVj
48+6KjOf9hqdfgKCU7UwsWvx+lmsqQR0kIFzuZGdlLL2M+C/mXx2C8twWKjOQCmZ
GAOymB4JxzLtkE9J9SEiPLJPaRV8lO16/qnUK5dRT75u8Wgl4Fc5mzem2H5IA7v9
WgfmWxvD1O/IHnfKsGra4BdpnbyztkF5vjJgG+yetdvW/gjqoNLYQsZjQT9U5R6k
UzTCas9pKL8ziBRCNEdUHp2Q+UVUuPxNJ2L61+2NKXB+gXjIAHIBaeJf9OdpG+qG
k+jtirxWaAj7H+Ri3OSWBPX3qwzBuaUmc3pZMn05aVvkcXLZgfzNcmYRxuhLP3m3
+nBvNeOW5/KZeuOgcjfSthio0tJ3D1jvY3wIZr/COEFwmP/i94jWk27m+hN9xX15
BLfeAedA/9pccLnf+mDHKX8kIKSb4m25doEJa5YHf2CzKWjR98ieWsOy1Ueoa57X
HlkedKivYx/FQ/3rNgASpud9n58bfbTYhj8SH6Xenqbt1nFsndmGs/O235YCsduU
Omzue2wfiqmew0gKlCaeIzHMqLro5fqfwdkUSmXxc9cDkhChPlmt0QUi5MY//mSq
03ZyIeRv7Pq4mqnTx12vN7KCBB7NUtJ8BKGpvRbuEO4u3MWQNHb6Iw9GVvaownk7
cUZhgAaPFhsOBKnNkM9TU4kGIteqfMz6MGkfYtz2scjAaFoH9mADA9Oc+vuEf0Y4
mGW9REMzLdy63z5K5Wqq5Ztr8nznvQYN2JSHfQGpvDY1mnk+nDyy3BtX+a1BGZHg
XKmmhMQ73lrwSmjObtXGq0y8fQg09O+jgk4HfYkfxvTQxmow1qmLM+vfKPIXTAME
IPfKraNL1pqR7ZMoKPCgxEcD/A+lV8hMccpaBd5hjKseIXXMQdmq7O0+EyLT8mZf
9SrcXstKMMT4ICu62dFzpy/cl/aedKL7MgTL3VtwPMb7FQo1B5cw91TvZZZfnP4X
kHDCJzjsAN/LV5vwyz3VkzhFc7gZmLESUOWhyscZiBCfcAhhHjNaRLg0lR5C8t32
dOZ/ZVRYPKik8Iz356IhhjNLkMa/QXuGomMB2S++MnvgDFAQ/CE8L3uUjaHawWP1
M+Cws0uwvSH4OYysDjKREHrDkDs1wWzPqwkVNAANcTqYeS3H3iDXwI/x4Q7IjZzN
u4u5JgEd6t/y58twBZoY/R5xfj0ujYhoqqIkmrILd8YAGcgXQEybsYzsI8LwV7jU
cnfHJF0tcJDyhdj+BI3EjkTBirsPlihi66sGj/aWx7OhwbnsSy/PcUmOLhhkbeZ/
k3rBPXeAa6BW3Jq76f347nDcW4sE+hHYxvXGq6O1xopnuJy4ogMqHb5N/C1oRNCq
s8czCg1D42xHUYhLrPZ64833FTQ/ndn9KtKiZFw7B+TeHsAj6+L9lMeXLEanu5NE
wXYssCUcY+p3JScVqucWXhQkEf2csPEvGc/xokLKD5JeLgShLDKrdR6LK/gRsSbH
F2762TjyIgKS1fMQxEVoT4YQ5gU2O7m5y4oGoKW4Tv6i5OgBVrB6705QSHPaDwJ1
DZcyb+YwVvIhvKeLjG/J4SFwDYwlqKP0GQcuye4l7CTc5jmEr8Bztgi0OTQTeeQs
YbCFQPk0d6BcmDYs6V9epMsk//MmjkKV0OGesEl3y2VEZOTk8bMhvdszVXD+uPR7
ggwY8VYP4SAcSlbOIcgoQpwAdv0e9JjplJCLEfXLt7sBtXA/i1gjwTrV6Ie6C9ik
0GoUcO7z5vOzAOVSofvAwbb+Bze1a4MtIYTpVPZsWHxvbKC5sTvU7uxx1fXSMDBT
6AFEoRWg9hzqinSB25+Rhkd/kPE6/xWEH88QDoBFqWrsevAbo/oJVlwd41kqEs+a
0fmCPEjwY81GA/5zFa/BiREiB7fjKVpxQSUNG4W9XBjSq2xsyFATXmpMupzDeIid
r6zUBwueSSpjcv2TzD1J9NG44F3vA+a0XfKTJzdhqfJr2rYB2Zkd4JUl3/VEc4x4
5XQuuOh9oxNbFd3g377XZFr+JBs+F8P0SUZhxGhPqTdg683s7+i01sU6BdqDEmZ6
EpVRZb7UX08c7oxibO42urMU6JB6zMuuU5w2JJ/jk/CR4ORLhyFs+Ao62EqrYbZO
jkBU6Wc9D0JsJilH2+8H2zQ/xdKra1Pem3K5RxakMce9VfO6/bpGSfFUOXsv9cdC
y+4vEE2HQtFlb9o0iWcOZUJFmx6tTyfm8txYWJw7F3h8d/2s3UZ6Hc5t9HBUWwBD
yOE+1g44mtdUZ6PRjEKJdbykBKOIz+URDVB1hVAb1PVgjotLUColwyaUqwgUXLKn
GBnvtwSpirxOaHpLxVzAKEMCVS/aq6U1c3K7O518DWnA8Dfi5jMQnsvpnpLpT4qB
tlFhWpotoXOAtDTLRcgOp3R9yztGCLEna7VUqfbgSEUASAHTXD9a+gq+oOC8h7XW
WISlLSm2h2C58Uf6sxnWpRlrH3doyOtcXOd+6Av/z4NvlwdckgkRfBjPmvWkJ6I2
ymf16hCbpGXOeOluk0Ylq5gDXbdLiwopjgAJqbvsLvotWUQ3eQbw3IAYSU1nRbf3
38I4gUJbgizw3mm0srvClVKf0a3lhE7S98gbnzn0Lxc97pW3AsAHXoST2t5G2rpH
dzKXavLW0Zll5ZBml14jtTWx3POygzJ5nHQ2Yiqa9WW/Y2xlV4oPmcr1RTx86IBw
wsbahWecQhvYscqPR6jZWF5LP8DVTVQR/mMr+A1WEXRPy1XWqNHe6Em3HjimqAo0
+yT16m4YmSs2krmrxDBSWCMmN9klUMkbugmS8TtqClVto2lt7kkinXmfMXmXm/jM
YSXfzIZfizAeqMSDvQiXoshkhRxRJh14kLtseQH0B5Cx2sz2z71k4yXzMVPNzwuR
wCZBGmJi0EbpFA2/g2ao2PF3VkGOGE9sy+2YaT5/ZcC+9XOIPRIFcPlgkJnxBBSq
Td+mttmnhwLvgkY1VUgbZMaF85pyIeeZ/ffcfP6iTiv9GLq+x3mJNivKsFJwOUf5
PDun3lnhjXGFlsL5vDz+8GuNfjoMegDAibIYrwAUnurujaBMDx9b1VIum2zwBaVn
qHL+n5TloZV7gaNM/0vDfEtxXlgr+KS07YJ62EohSclNxuOqxoQ9vLOfQvedMxOy
1skKOo8FORkKvSr2BalsXYK29jLxQIYYsNbNAJdbcINkONyDkjhqcQ0b4G/QDQbh
G11D/dVFr2HdwB7RfNweCVVj7OfjOWXqlM8agVc/SrhpRbiBUipH6FuH7Ejt6XK9
2qnsdglZluUNEeKlNNdx0j6onZJA+mDYFQId/oTRvqtAfoSx0xMUzkYCEF8v/b0Y
5kozKK3kHMYvyCKI35xtX2qUxRn6nmxUsysBkd2dVJem0B6rqm7c8WER1/WhVr3K
GGdpjt0Wrnfy1q6VxQmwbtj4CMA98GQ+OpXV0BlFTm/SFYKqXQ493OmQgY6D0lLl
QPt74+q3bsBu2Xz3MkXl6bpSwQNYr21lzmrBW1XOu/TYkboFovzUykJOMkcrab3P
xLtfuABUeTZCT2+3ZqqHFB8Ug/Ol9Eh23d0YkDGk0wV7bjgNPJf/DpWcbFrlu0rI
OoJEYPF1YKSBgJ10mHjHO0Kf4cxyxt24te0PXn50gifBIRejmWMUe0h1X1MSZaWc
+uznZVsXqUKLBJAB/FLNGIfY9z59dXe60C3lvjtwCj5T28LMVxJQKtl8qIW5B8qn
cpcV9pPSqVFUEhfcw3CUQr8XBQEVne+vtLkIBXwKpbQstpYetnjYpbKR013Oz5tu
K8r5Y5dmpzfEtbaqt6whj3gql/4pbfcIHQyp16AtR+B6iiQgXudiiCVlENGp2ZQN
0Sde/J5LrvAXKFrjdvNhXN/SuKWSdXmHdNhxehZI0gRKkMdrx/mEFmLJkGlM8bJG
A7cgWy6KCG8pto5EqNIoQZUT/K+vCici2F63BVzDwh91t+8hRMK2Z07ahT8SaRLn
4cOLnaSWYMZtykErSJPcJWKATRRMbMcyjxXGRLarbBYnKe3wAsAPW4sFaaukZSl9
QZlxwMYtnj2F64q1EKIlaJlvrQ66UGN1YX6z6d88SgbbOYUWZ8/EfjSf5+pdRWq9
QhdE8QiXvy7XDT404zIX/tv+wgJqxaH3VQjrv+x+CfgEt4TIh4v+tmXK8L7iuZUi
JAHe3h6ougb9Us60kHp+NUZG3bOW2IcmiD1HocVthhoqYRD2TIsLS7SCZz5n+OaC
Hw+uqo7TlCUGnex2BhEiJo7+j3Epam3PQUn3Fw2Qv1D4emUhJGgDARxprIEHcKRo
f4tatP5x1s74jvAo5MxRjAt5rcoEMQ/9y2GcX4T8xFkj/UlYeR1yiwLU7qU2ha7m
j2ImCR1gqp+jPzY5az5RyQ8SCmex5oA+ZDfLxKSRngnHAG4fkPfr1eNoF7RHYIo/
fzB5n1PrSq4Khgp0LFB80DTyj59munjvqzrt/h+l6jmkDS/brL0+tp2YdUOhl4M8
kd1ln3FTnAFjFgICOc5JNOjJ+/X1/dUREsrvAQWJNlkl0lRnGXQpsqrcEc+5L3ci
PqE+ioVAj0AaTvd34WbuHYi72+GdUBzo/r+7RItQJfSgJ9WVul+zr4sEBZa4bNq9
CxXb9e2v6s/1KiofPCIgyGhkPXy2Xr82YPiZ0/bleZTY3Jgf03JLNkt0l5ix3zRE
VW38uHQyB+OLKUM6CGgF0KKHoioGJl+/DEVBcERu6KuekulCb3/MzxzowscweHFz
86zhx6eDpVDTgzldcrS9Agqx/cwX9xoGdoYui4xTwf+SN0uKjHZr75HnVe1aq93E
zBMyvjZaF62VRIY/rt6mt67GIgvIXoTVcXyZLfxz2MWTSJ9YutNfXZj6wmDysi5J
GWTPMIDP4/0jVneWv9C31t/i9G8X7u+18fjcT1QPjM+iO3Y8xdu//15KyRPb/Vcb
7Lc04W3K1ToYfaREfV6PotdRldH+X3MgsstIEtWEeXlQlMdN9FyxXIAS8Lfy8VYa
f/BBRRvwekurpgehkPrM1ICb4iysQFyvcG3WZX0qJ/AEx0FckMfOrBa3bDETfemG
VfhuqhFcQ9Pa+K8jsvc+34S/NfiBOHv9jipFb5p5nnqSoomLYj1jjoK+z5NiBfsI
4b+99pwTWP1KiXH/+gb0NT3cJg03qMV+xRhStA5HBccBFG9T38WjBcnHmcPA/DjF
Ei/va3GJ39weQWX1/g2d8KSP1gQ2FMJmHDo4sCbIJqrx0lwMoNGbD+HOPihutQvi
+RXwKJC9IgTI1sG+rf2Au3KuIteFHNVEMqFMg+TVu3N8XqTCKm+n6Kd7j9BZ36gt
oIlREeidOstXAo/7953BdzOl66Rlo6TfkwIzHOHPeSxSayDaxvM23VgjwmPUwM0d
xAEPyzflf4fHDZ36AsIVoQqzAQ7bKUwQeh33JHKMsH5jRbAgOSo7r7rvs9HamfCB
7PVeMi5+p9t2rOfh/tUUWouGRRKMkEAnqy6IXk4La7FxnIzjRV/UrtbzCoIwHCxa
LRiXE6ALtaatq10adEnCaRtOKrfBbUCvDMpQfS7bu9lGt1mIlxTDPu7C1UtFoZ9p
H/jO62YAEK7+upEIJyxi4jz6yMucFw3VVQdn12nGq312IhKDUmfpt3XkL9riHSbZ
s3neNMgjeooCU0hxT6HlF4z1VksTYiOAIURgWnEfEtvHLabIEcYN0wOo1O6J/hhP
t10EkXAnlOwuRrlUy0Rs/6Sy/7mAYxQfQ3MC7RHf8gOiewC76MgWjNJ2gsQbIjBM
imkQRPUwXLlozG4W9DPY+ErZ3asZ4XjHJf8KMrR5WcAV1bAfL+/rvDsawZ48N0+E
6eviSU5GThbYEZ2eLVUmo5USGCJInyt9VT4/U9e3qhUpaI25GMtQ7rZrOVRjDH70
LgZq04zKHPCBrqGwT4NG55szULJFanyHGA23owIup+PW8SD32B4bfzyUq3+3+YM/
Ag/WL8O0CJl/5aB/VgK9mMDWougD+ZcvgM2zfvn1MQXlGneahK4/GoonMDWpMnTw
RGsPlq43fOPerBouxwRXaTIgS3Uhxpi9ieU36hPPqD8T5mp+xBFSduSSiSQnEHZE
h8aDS03ux0zvspwDc7Q/lXEhPCsTKWPnRAYit7a7M03QoG83KCiExEWvcOaTZ5md
p+3yEXYUXoOnp2S3B/PvKaIqB0ALFriLCoEBhutROEiQORYfZmiP4VhO7SEdYO6t
MwH0JcUrP8K4ihIvNbMAO9AKY2MKgnOh2cjZlBoGyMyM9g13wtPfH9ZB8LtU5gw0
JhVY4Y4UxoVVsuBZcWs415vqIyAdiqzN4bZALNQAyBg5uJHFzdPGFeA3QecxRgJa
tiwK9I3xvIq7bsj1hq16cURRfPn9UpNH6P1CTDVf8KKcPLgAVPdMgAFO5eR1JlWT
0ZhNPNbzuiX6V2gtTroHk2nab0n/ci+BUBW06XN437RkQbsKWMyQ+SiZrAn4N1Jn
hmu6c2qYDyfoHUIfrubw4g4fhah4HR9q3tPcVb9JiSwzSvb6+X9a4E14xULzdgWA
c9VZrAipBZJTKansXlgwpeA1AIF4OoWlZrWVMbv5/aMnDbD6CwQmgPxlD4DOmoKm
B4jt79R3sQDg94Xxeh5EYsHH1K/zXnile8z5JJ0/qUetYgYBYXF3d+64goUaoRLS
IoYu1Qou3BTOPLLfCtLXt9OJMrXclZ7MtgTiGtGyQudIShrr+Jd6sIDvDD23uMp/
8XLK5O/Wz4jE4NhwcpKnOTho9eUGXFRZ0xa6qCXppVnaRK/p5WafyCbvl+Pxqs2n
SUoh/Vlk9dU1HPi4qDNy6QOcz5SdYycZ80eN7MlHqHQjEe/gzpTfuZICIi4BsdbT
KAa5Qy7RQNoB+QkkT7IAAGRS19OPgqZSOhhDLO1lDmDF/k7YDQwKxsbTQe03jhC6
H8PKJBe0eJfEoisiFJMjvzuppKmCqHAuDy+anKdq3gKnCXwe5j9wc7rc1uKK1zgd
HT5dY6Wf/1SnLYEbH4mwdbaRltb02toqtQxZgXWTk6Dv6p5Ant3bb59zSv16g+Eb
3NkdKR4PXyzJapD25IRUCe0UbGW1x4gBfBvCJzvWr4HqGfBdIlm6FTsS9ZLoEErW
lh2tcu3K5Np56HwL2YBz0xC7gSAf17a8dmZ2lqcNt3XALl4wn5kBA5b7XFG+Ihra
aF5KwigUGv2KUzymF/YE5QW/5N2iMBklTplryNWStFZvt/eCCKRkeX8V8QelOFmL
NwUSnSQm6nNxTknkzCvI5Nk4+6vT3NDFC+Oxt8VWISwzCXEicU0wzJEpji4bKLEn
1z7wCQpWoU6uJYyU0OyjQ1yjoevvkthdLylaz7B4fkfIHGwD+s288X9xAstCXIDR
sGoC+hHhpD4YnsW2+nkr0aCs8oZUp9GQ1nGVv1n7i0MRuyhES+4szA5++oWrOfg4
306s8S/sPb/kZuVJTS147bMGgaPrDzpNFRLFb8QIldAlMdfhTHIWCusPJMG/a4sV
CxcgxzzI5teFRwFX2vnrMbIOTWt5hw+68p0wVjc+pAsxbpc5uEP0rFxfaPQ3Azio
qY3Jm9Q6peAtvRX55y3lHh0QhFbSaICB1xn0qwkZGuHFoaVa6McV4xdS6D4OrhTg
T9Q9cYbRo0Y62y02ry8QmAEbVzDHS9rlDgnph9/B+ElwA3uA8Y1n37pBet7M22Sn
wrlFmdDUkYNLu1TJ4GkBxPBZK0cda9jjEbQB4CF6m+D/+atPQ9o2rlBcTFAG0ddo
wgDWifmllGvA4RPXEzOtK38Y5S2mxCA6e8xduqMb65omqsgky8ZyXYIgVbO2Iuq5
S0TIbu4kAOk47RH/vcACO/DXPEUfFLwSbpYWppwQvuL66vVYCByP0rjVgtUAiWJ+
UnRDsaaZ79FwhDpSw3s1WmiXMz7a3vqmMiGMaoC1fBAtfje71ceDdUh1I9VDLNqH
r6wBqpAxwC3X0GlhW+5rAySJrgufMFNheTxZZO57+g3+kBUO+7iIXjasc4ITsnEd
GfxVfmH9Ok66BpKj+cDSxUEQ8y4vaKCmPUjRoMAjTmXVx9tVmIbtlHrELv7SrKhW
Yvn9grQyK+kY1J/YdXOgCpU1qVEsYyOh08nJhj4M7+eIHARnsXqzw/N7fHR+xbnp
PE7TOPxYQgDN8+oxUK7nCWJznTvQCf0eKukEfCT+XwnU1ZQP2sI4AOFPXI6BQtJ/
qSnoPhK/Uo2Vj5nGYm2Dfek+Hrpho+NrOzoDD5vdn9yxjRcZRNJ70k3rEuQq1Tyq
O/pa23122tuecNGflQx4HSQkNTC32UDFWvvxb1yMygE/g+Li+EqApdokUdGG7Za6
nRDwtGQnkiUGggQkg1H7nPsbxRCJ4VJ0bK+LUITgmEz6CAwNRIzgQaDggzQwutTG
UwFPVify0kiIKqOlGjVvt17RB7glQ0Ejorhxq9VztGlmMTry5UnwnmuZntaqylpJ
Ty5ChEvHYhGclSI6v5Dm/S462mI0uEsLDe89ZWCx5AYQVbmENHqDhHVXlXqDu46Y
3mxXdoKo+TLUAvecO8PMOmgO3AgyNtMa51TH5cc174AcULGULw/4VE9aSXqBi1aa
fSMMs3XuC5NGchhiRcfzTCTDOd0Twf/2EudgRUiAN0fypQT0kpRONzjmSUAC9t4O
VY8aeUe0LCI+vFdFJq9TWJsNvo+NdvgMxWsuE2NpMGeZ9vPPA6HShUrJGi97DBus
qb3ulaa4gMJA91Xj46lq3sOJcl8Jg2QIam5tHZ7bq8bpuxbQAXqFPgSvDfaJ3/aV
Q1/Gbaak07+zmCPNLeaYVSRRd8RzRoBoF0qVDpVgDu0Vaa/Ww0WxjgWV6XI1nCLH
ercqRhMeysa0UsGZdgm71CddnAllcANZqjMHiylpYKBm9F7yfNIbyIeudWFbUSE3
GRFvdZrkKaPbBG6zMa5QjuIkeA4z9ODI9hFAVN/qhfzMKkQYdu3ZnbDsNJv7fh1J
XTHZBQVHMuDqtiGx4t9wBvfTsPvpibOPN0puKNM+Dkna8KaG88XJ06cN5BmN2HjL
KDfwz3ZwKVJzPZ37T7Eco6DZvu94wiyKvt7ac7M5c34oHIbqVxVN2iq8IW/GCbYf
C3vGNhFvFStw1rPKxAZeLhSk9JwfLUt+u4q5U3rwIbRPFDal5rQdFaYH4AsOUHre
h57e6R9+g+uQl2rbpZ/7v0TAACRkU89Qs3WuQf77QwBrD5IaYdHjQWe/6MQhQwmj
s73yHsjolfEpE1xkgEt7WfoNb2MRWuDuwjP9aeR/ut5/xXhEaC9LK2hBd+lwr+vu
lKde5385vTkzcij/yu5Hwx5nIlb2ZZG4iUVKQrD8nxLhm/IHJUBsihqKIasmD1hf
4VwQNE9E7n1InxvUkeHpRr+cqA2j1TS4CXHTL+FN+z6qgfcHMj69Hj9PKMv706aG
7XrRLqUYIlLU08dc1E319bDnsnqltbSaQaqHKKkRLLw0NK3Xl7t714lbEN+gxQDP
vaUuuFXdtD7bTj6bcyTeFr04Y0fgiX8z9ojc9d+TQQuDzpPLX/axYFDqhlYpN0D6
uhZXr3ffAXxmB3/ihblJKTMrsyfwPV68m4U/3sLkeqBi53mKmp2U/6OaDJ6XUUhF
LUnWWkQY9eVEWCF3xjnMKmXRfiRI2JE9oPBYNLt3ugv/vLLPMV1zc9MPiqf7OOl5
XYz0XlWCEhvRhWp6TdcoRbIP6xPxL9mJNqPm8xfuQBDl8Y5Ic6CWK0ljmxWxagzw
gd/gv1eif0lE1YKEUIUtP9v166sBLctojxSq4cpk1XzuOBWs446qr7s7Lq4rClQP
B2ksyVh3gIkKtBhxDlsTo60TkGQTkOTlyAehEyhwjxmRIfkWgmg+7g8c9yvdMWTj
Y5zcXkopQfXbzblouqNW3YgV3zru5W5/UtMlF0texdyZo/TG3wgQOPZwWULWiEn4
t6QLMTebaVvpk+FNhNbrtCOxK/atAgYpvnMTJ8a7QCRJhELZOvW9k70mNJA6mBco
ULjNCsx/uvxIFxJchaLq5qrZ7a+B9TnOjUgwvIm/pvsbKuLxiYYdwUEKz0aUsgYP
h84Zo0OPl4DdDp2sOhGFKoyQIkXJSeTP/rAQVoQUI2GHpAsPsI4nsnk+Ljk6Ocbm
Oxp7dQL6l+KvMy/chbmgBkeO8bHrFB+kcnxWOUmd37io1yoqPjIcyB6Ryp8sVtIQ
kRff8MhemWSwV9RrMBQC+TaG+ozdzVT/SPHusoHfhYlVIktySG2uG6haaKtlRquQ
33+xw2Labd+XDH92OmSenoZ5/fdmHOxwKmKHrR9H6fczINvmsAY8G7SelPqoj13j
3I2S/7xakgFToaNzrmJcibGO6dU3cTNDbwW786xJPXxpjhbekMRsjucM2DTmDH22
iqhDZrJG846zJkZjI7q4CX0IM1DCPNyP9eavcVDUWc+Q/0JDU3VsZxWbk9iV2Ggz
PVNx2H9YSGbvdDZO/BTXDRTIPQ+KYfkHPh3/V7JhpzsBIgEv5PTh6W6ND3DffDr0
zu1Iuvz0VQ4w4r3TWRhWU19+KD2G0PaAlGCNRxCxtufKPtWdW2RfMkviJoEDJkL2
61VRBaygJ5SxmcCWlmbb+PVZOrgLCGb1Wk2YTWH1ovKhMtzQI7arnMhz39SZegFG
3xFAqF7FPhuPwNWkQ9EkJ+gcLsoTPM0jf6bIgAapzX67szA/yesUwcolXNw5Ep9u
R4AO5Kn9OFNqD496iLlm+8zNixHpRoIYa7kMm93LXguSjxhp3A7u7EO72RXe2DhT
ESWquoCCGmdmYOo6cq02jYJMMfKGfOVuzZRp5XQ5QJY/N+FLFiU/vPvuApF1S4G1
6awvLxveigHoNZDQHMWyXAZiUiBABITgI7MtRleK7MhUZBpii5MklI6rbXizcsCF
3jrcRLGvPebXlubc04HB2UeMSALye3znt0GvARQCyizaku9BzeZSaZ88LGmj8vA1
1E8ODFV/u9fDBntsWBEe0qNzFGOHDyOGfYKOKEQ4i7AJvU782wkyc2JxjbzKcY2S
PjVjRh06ysuKVpmOyLRYfthrNPiss1gtE86SfTktXhXD/bvLdp1KmUMYDdkJ68YZ
2kdFQHA1Iz3uk1zirvbIqEfR8ClQkAUQkKLrtBy1QA5Q4U5bAv9qBezddstx5KUE
Du4B4KzlSz48f6FaNkudLMPXDQ6A1hMSCn1x0NGh/3bxGfZqJUSUL8bbHPQfQCsq
GxJfTSYCu8BOW4hrsTU6C1SfWZ7qxMuqMHAU7nWdBeqe5uZJhakUxVJDUXVedimZ
z2JJPUZJTFR6jqyz7jn5gUE6TWEll5o3KClpQn6PGp4vqiFOt7ihFm7SyxTVCsmB
9UdgRO01TZIrAV+H1Skzkj/NBBMKz7Wm1KoX2ZSyaEPNUYWTzF0ULjgKcX+ui7CJ
s7dH2JtU0sivRkQlfD66eMPQyMh3KIqbFWd8WoSTOWgX81l6Q5V3wtEo9qSDmuzY
GtmGAw9I/npWlXu1CO46u3Rygq9kHgCSrGMjMktOZHdtyqzDPhNGmrODmmVJGRhE
Z/rISXpFVfkhcvxWzqZf1ApGI8RUMj2oft71WQWNdTVZOnlFEWBMmwpke8Xjw5Ls
8g0ZhsEggA/tK+56iwQtWwxbYGOvL6bbbFeUolD1/c+QE0gg/8gn8zIgkO2bFogs
RFqmUgyZ+n9J6kHrxJlfi6WsHXlSiY2BUulHpUg4N/9Qp1ic+/574prSRXcENz6n
O5wEKI2jwy8Ps1stUukgrePJbggXrluJQxfjQcr9bqDMJ4pCQQ2CQ6yEpihuza89
iKTTnSyH6+H0OmVSayjCu4jhMrNhHWgvg33UnvSdbGnFO7ZGxT2D/0sfgV/i6de/
SWtY8Ph/uFFeF2vB2x6YOtxPqpPM2C2t34Jh284Dy7iMQYKJUPzSzS3Ax5Yi/5MG
0LRJWosLXT20u6N0aWLXke2h+bfWnZRV7ApvDdSQntQYo4/eLyJbkImytk5ThWkI
zs8Lf8+slkL/pKR34VAYMNcfoB+/PYrsS66iLwgXNapgore6yES4THypuphNY73e
+AWD9gsre8xGKat+zmYd5S3NZqb5hJNnqOcasL0sX6Jq7P37OSdAnBhnfYb2n/5t
AU0OH45OvMu9HRM3qejau+hQ7ghKMK/d4eSb1KXUXhdxQ6f1bcwYcrdHhFY5uC9t
T1ugAeg0O+pBwsGQPzJ8EKRJAS6/TeCHqBbZK2JQZLAEUSgAeBvyA5ubATv1MbNy
ygD6J/flT4YAat9RjEf84YQqKHdE4VpOJ8vfcCO4tpVaVwqPta//kRjEIE0J949u
+ttm5fePTyTYFa/FUClRtkJQzobB1O5AzZVRDPRlnti3xQEWcebTTpdIwEI0F9qa
LSC3d4aMFMgCC0auQWkDyeyahNg7nuU0GxlQpO3eAa3tMqWx/53DPuPnIAEsx7uC
y/lCns9Ydj3UV+hVfCx7jk7Z2P3PeLnQzE6+qjDV5xH1GwNgkOqgWTXwdVVaLSIL
p+MzolGSHuBXWALd7h/fNRCQZULFtXT1yxdm64jPmxm5BT3lnsz6fMPwyj49O69S
N+zv/rHIwaOclR6sz724hzxeT2YA9oayEMH6e3ToFoi43SD6A0qJCwHsDIxqyYh2
I/UiXfHakyYTIwj3jPE20fs6W57h/Wjl3nF8/blbltjDxxijmzDOHOkrilvx+skZ
y0nF1fhkaamDOFls7V2HspJqP6FXeySDQDm2BSCdNo2IByM9zU5g1yRhNoHLTu/C
9StUtwjIYx/i/kaDdUJEv3sD5l7BntrriWw7MhJLj1bIJ4VQzkIuKT2oT3jqdZ//
pn4bmaFhFv/W5WGpcUHohgvn82lL2j4sv9h2dRPbxmcTvF+THEGwr1C+IrhfoC2u
MCYymwjkYIJkt44ksO+Qy9cUCkxWquawSXSxnEULlUXFIDp9wz8mo10FiztP7URw
2Q6muV6iAI0XWeMwaZ3TKJXhDarYVE9BqaXiKufWNx5StRyFWO5B1vGcyW8tsRK9
hX+Fd/oMx//LgMh6nChWnLGTeCTzCEvei7s6q/58bbzTW/LCOBWbBAvlYjoeHOcp
Kw0wdyMGW/tKaukVL0VupLo76pJ9DqFKdzrcfMMFDNU4CiSNHRyR/u9InFdP1ma2
jEwBASb+1Clf+loTPNPa/14BYDCLTQyQZJou+v3F4PUw4tuNVnuKhWYt9CxAjLns
Jpm8suvJVgA4J1KghvubJx7EKQNR6VwsXLx2ismsnP4GzpBvek2vimYKzu8gcOXr
Sgxdb74XHURfNnpIpc5UJbuu3HmmuH/ZAVvfpr6NkXPrXJOk0nabyy/pRbALEfQl
GkvjQwHE2Yifs+EGehn3Ccx9dpdVdFMnFA0tOc2jP4MiQMfasLaP1o+PMvBvDGsQ
r3asZQGrFg5R2m0Whe1N93jaZ7h3u32YWZt8IhifNaR8K1jDow5vfAll9O11+wwa
cH5ZeOqRRIw8tbYyX7ZDO6a/OF8vW/oRAIlD5dRLx1fGkC84QWn+765eSQhCadVf
S0F5njOWAh7L9uwqRQgPUsBG+XPpcLPyMK3V2s7Q6Gc3uoL7YzefxfoF1QIvwDHc
7ksxvD+2PBxiGd8Su4CEU1huzu22H1cTulFoBAUIDa7zyOFvdS02lYVAhJNRnecA
2B2heW3S1XalX8eO7EGFvrHcagbfTJ/nCcGi1UotrTEvtfye3qOErAIh/Rphf9df
y8hXySEcys+gWbNXClP7o3Zo0KbpwJyUJiw1ZLBOE1YrIL2z/xMMnvG+FWt8fKnW
m7ICvgT2IY5W7bBZLp/evMMGcIqEzfQ2vUFCsQG3+08O3HjaD3HanwH5qzfokmgc
eIYozd4eyhc9rd6jOqoWF1lAP0qPzaDbrcI4YYkWR1egiTuJBYYMdoB4IukNFxyn
8v0fsTqbrEO+2nlYnjpMreR1aTA1fL7g4/9GH+p1QADOVWvmqPJocGnus8OEATmD
TzUyh/ScWRhznNXwpAR3tUegPX7h7+XOCt+qIC7znhVfZpZY6+ti3UXMXalUyM4h
aXFfZzk0awjPJg8aLQhcFfmQ7gcm886u1pUyIQOm9i0/YRIGTm56DVJFNNTlRCGa
gnTlDPgGyuPcSe7gjRv11pAsTdMdALZ+59Se4ndvQQcm17M53TUdRXaJsI3kTvUD
QomM9qkxPB1oNb0HHuzMNIlpIsCmP6ezyKsWTzHF4rhRN1KtsXoO4O+fr1rJOwuP
F/lqHBLkwpnjaCgubqII+aCVPcFSnVKTNrMNlVptzk7otVoE9amau+Xk1mwQVlMU
knJyzykdItfp0ie5srY8ykmkD+JK/tswdXzak3xWkd1RNHbLFv5cciqmKR9Fb71d
4s2dRxXoyjtMos99OhcjG0P279e+B0LmppufPKnaPNs9px/gt8KohMnTGDjnrnpO
o/9Y4MFZBIQBbusrzCYwFEcG4JDe1GZw1VEUE0NRVvHMi3TzH2aiy6o7RALmnkLc
+KPpFyNOfVd9klGEziGQGFyW+bUjtIDEp0Jm7Fk1KuEgmTVsVD0ZDFPSneu5IS/h
uBtDflcQmFS8IrC/mOW7Eu8B6R/dm9BKWvmvGk4DelP27HcPYKt/QuCwcvnU/Nix
D3uhJojvQFLJ550kP3kfYfxGjMuWh76puZBTF8mPxMziPRUkodiuiInQXf9i9m9y
cxFS0q4kWwuK2SRoTQBvb+iS5SvoTpBF4PNBfr7PHF4wmsTa47Q77pguPIJa0MM/
EonEfaByDcdOVWyBMlKT6tb9A8nFZBHVtYZrnsd5XoqTzC4I+CirfmQoaLP8LClO
MVfIlXiv8K6WwkinlA6kMJm2Z9glXb80fMHMEl7bMooTe7EQaSPAlNWlEOS3h02p
ZSOx2utLqoLHPKEmF5L4fftH54AOG0rYu/OjKjY/JyOU1fP07hAr0K6q2t39HR6j
8pt7RN0b81s3IVJp3JieeQMJemPoXt7nKGKQkg/cK5fWmY5oR6omlDXPYkr1oCa6
4k424oPnBBcnfy59uK6Jzw6mtaWfpuRFOU9JaaV57xk+wyI557747qQ65f9bHe4X
QjvA8PgT44GNyORP8s2dJwkkG/vwtYVc/3D7RMDHY3NogMwblMTqJUAwpHPy1oPq
cudcAajqh2IyJCss0kub0/zlPTNe0rJa5vy8rk1DSR4q94R4c/oKWFjpfxbuPl6O
CW1QzRkH8Onf6d7V7uv/Q98GKqS1tmVRnfFNWY1bSYeW+kfIXfL3AcJyEj3fkyAS
q6YWwu+UwiLW+Lk/dzisxxM9jXrOI74tLf4iN6yeDQicxhO8SS5CAh/6Pn7ehsG9
ANDmxtgxsgKPyfykAy6zEkmIjYwuuu0L2hflKt2u0zUHFKDZz4wyp5SxTbHCdsPK
FOoKX9RnM+CdDvV+W85l/FeCvMj7YcOnlQ6kxEZBqCzTvHW9jQ//IHC9bF+4s4hQ
erbYSGfwKdATbUUxlfHRsKh4XhU9gaR0heHiUtY3gLLyPfDDb30C7wEq60OFnQXA
clgf0GtwqtGWMUfQ1DjXRNkZZDScoqR3vDavntPnHnxKH8xieaJZKJyrCz+ay96i
TnxzJbf8PwZCLCQpjwfOhS/6dYKHa9e/GiCsozIoCbMzHwXs3b0GsmdRnjlDjPZc
GOqqd5YyQlM8GtPbb5u3JmX6RslUG8t2ma0s40odunyO5SHwYTOQi0657d6LzmIy
eQ6npDXZ7kid2tNDgQ//b9OL/cGiGeJzd1DBVKUzDZtr63c0ioMkA5dZxrYnrR1o
t3oKCPhXt7GyV4Iu5kNGruoAAJV22tplSs5Vc426hh06YzQAuAADSaZX13LPjXOK
7jsC3nEXe69PFZ8fEiTCo7G/bQjxgoLk7iyQ5Klfbu4xnuG1czOejHWd520NCZv9
xUOhttePSytodCd/8oa7cRHg/pI6qMNYqH2I4dSDGyW5DFynQ92kuP6hMjcTljvb
hA69/vqtNn/3unUy0uz2dep+adH3B5EHkf0nos+Fa/d6umdNj8Vy/FZ/i0Gpkury
goBj7Xi1X+bOvWAcuDvkL06bM6CeOwuATVhG2Ke3rJJuopv7FmeDYI0CD65HIWzq
L/HhM9TYqAnfp/lkSQJfCgmDN5IO5lUVf4EXPfLM0p/Tl6/qNYzneojn6GM3gPTo
DDxdCRGqpo45TvD6gRX5h7BaMVRjuEsHRLguFYZ6bFJ+rWRmSUgG0NDBrfOLJoXB
pz4OdTjgkwOtNm2Tn3qw08WCP7AdslhNeAjuzHoPRr+0PsfTSd6sYI8qSvJ0UB0P
qvG8D9XR66x33/14wXdVxynzIJOJPFfY7oUc60lDVq9LJKgKwCeH2ftKkIzkKuPy
zeGn4g7se5n2uMZbkA/vxWGMHTi8CSf+7NptFyO42WGNNYq76SPEMaiL6EAJuTxv
+3vL7fCRL7Ow83zeBJNmRpdFdvhSmXDBYl+Ik8Zu1ao45+Jw0sH8NmeWgAFfYORk
1JA6pPWoJpcGT/O4I29qsFaodi/smJY7SYHY+U+EH94QAW9+bj4fVNtpXuId2/AK
MC8zZ2qaxGOajEzagdKqoCH7Yat6qZU66WgvSIYp9tVXfUDtWkLGwSlLMRYZ4JMy
l7DVecq5lMU6KJQOFws89Mykl2I9Uc/xLryf3q4RFW2utIIhLaADXWn9AJoX2A/4
FB9uclXfPmQ5YQ74KdMtDKGwc7B0bjQisa3+h4A3A+yjMcb6VskThjt5K9HdVE+W
0ooJjexo/F1soNrZMBw0Qtx4Uw+O57FIrqpg9xVGy6/ehdCijWqt3FLlrMO8Jxgj
8YXNgL/CLPsUkYtl6MaGenRzpuBcW+KJ+ibLftxEX9R6n7/N4qIKc2uMtbl0QAyW
RXD4v1MqwMdJAZCP3WBBmIZPpXBHOBVNO0PZUwCq1RKGrvb0gEqLjtQZOuX6mIVO
ArudA2zZsNo+13sDEJO046UnCerDhDvXxqUONNaFTxx3BE6q6zRX3gePDONCO2EC
lUSKjjOj9k4gSsxBz0zc+HXuTufSRuFn8CGefb/pzzDEsOPNL7QACmUQPZHuichk
Cty/S7PEK+KmJN9mNgQSMqdfO4Aqc3kKpIYkPHNANEZyCmxigY5hNcth4W+zht/c
ndgussb6lKCxxWB+BUn7SkL8jUhcxhIRhNibJwfvSbbc23HXVw3TL4G2ENNN+bYo
ffCqAWzmWxXsbLMVgfpmcYR1loNj4yNqzSacUxnMnGPglZfbWMdC6sWfl01ohRFG
kqJMqShrOcUX3lT+1t7WMSCZ4UaDfaryfxAuBQFsUnrtljhr/zQB1n/mQzjHWQhY
oKnVx8WVlNc4MdiKbj4KwrKBhybgTQZi+gQGi+f7RssERaB0d26ldSZxjG4Es20M
9wzOhExbsf8XApJBpM+YizbWVmobMh1OExP0BExZzKZYGmbHmstpL11dtThW+aYl
ecB8n5JHs3yUwoodwM4vG+UqL8LmG0bQMRLzGTIwrLIycQciVOfzIvOaLOEmze8y
lwwfBnXxeKqn1W8YV83u7JB3U4f9t3e/J1reiJ5UANtBzul8TL7c2DvItkzmmN5Y
wcQcTaVMz6kwtcjS6dRDSn6MrPCW2yfkAxalY33X5TIFKPPTy6QGnEiJSDMKFszY
Phxp4TuVHzHYYnpkDnmw3PzGl9XP2VOYfOzQDQVyelNnGfiyfDf9P7G0P9aGDz1L
HKFOdY4St73auc03IO7TW6ENbdftPVeFHvqZn7X6K4Id89dm+NAWDKmTxL1oSVUf
Aby9mHn6nMi5Tbc5atSRPf42cErb+g2EfFQdxXa4YqARIDhgB2k1qxx/hQAPQcSp
dCRs5PjnEnS9otOcy+RlaPL0tupJLpxDtHcEpesRSCF7cfcnnAaHxjVizcM8BnZl
2Itzn19PNnjoscsSDwq9k7IEMPIqVfIpjP9zeZQlAlIwlMVnTxYCjQhJwr/B7Gdi
5qJNr0XcYm4yS+ysC5w7U+sAgmGJImT9ezXNFYaMNctTwo12foosky27wLneTMrY
ksX3DvYRIJYUFIxlGRIRdE9vhk5mfehUF5af6PY0JrcFh42TjxAQvQfBL72UTkAb
8FENXITqYMLgT8ShUZ7AnazuPmG2z+blIrVEzzXfD7ivtBushbBdUHSjocRe1wIl
1P236dTi1lqZN/HmGqSXYJEF4dv/7HhVw3OqGpi2nOoMwb+BxAn6D9TWZbpmaAms
Jc1QTQ+bQiftI7YDkMGFAxzru6KpDVsfC+Y8Hid/DTLAOL99M77a/njLElIRy5iD
O5AdM+RxoPSZ8JYgEeNI0UU04hwI2Db9a+88iyz9x1injUArj185+ma3kxftxVL6
UptqdvDGgUzk0EsheZI1BNq2KbfFqBLZmwYo9v2l7XMMU70O79qvRBtjtU1PLf9k
jQTJdzW8rPAc67ArabqKi0VSKdPqKn0890ffUYeBZR5UkOAA/wDj+rrEFr1nNU1h
AVUgxBBLyUuVxEoZfrEYsz4EOOd06X7nA7rcAc6+cmtmgp+9pWNhiv4X6f7+XI+p
ykmcUMj3azlVFPqpCYoPqUdI4GwUUKghF8x6WYsvSJGs7mpWZsFBphswU/0eCTz3
WPuUGIxfWQ4bv+vDdpNvh7mz5ObFpCSSN5JLuyXxUn8DIVh73yd7kerFv6sOn84o
Sv3U64/6IghbxNspOWnRhUppywVQ/LiLo1hjyTGr2hSzcne3Itq/kjmEzO6afJee
ym2JveCUWYCrRFq3m1tEj69MGlQJLyzCCxNbaaP6zy0adjZtWmC2hELtRJV6qQuQ
6nUdDWYBui+TdCbY02rk0LtNVPhsD3VT/EXdQS6qqrhpzFZfrV683BgeoVu4RpVc
MfrR79EnCub97mxO2UIM1gA1zNYVYlrSNhjGvA3iF06iRRlj63I31Xh45zEhqC+W
latB9SokIjTGkbGe1PlBKUJMzTPUzO9WA8by/Knzi+3yMhJ0//5O7pSwD4IpngC5
EbOXKKnM3vgl4z1sd9CFdUcsDlvLuFXkIQORC6VB8UnFhyXt1BZ/7L2/x8o54M9u
CELKmukOUMjtZ4pIZK2KjUvJF1pekM5ZyiEEgAc31Oe/k7mpOs5qOzkdp/zXk6RX
nN/GV4dPCGHRKzUYNjiGkA0l2sWiFkfCIrJTFHAOF7Wgh2LgZlrk0TYgfcr4O1jK
Vk8CLHkjUk5RHlCL8AFR223MSCjCeXDZ/tcd1vm/d7ufdE5fm52KPX15Ivo5w4zM
SXWHkw1Mtpp1oCzZ38uR3sVus8HMq8IkYggLH40g5VNYYkM1stkEP7gEQSkkG+wv
jbtGeTt7wQw43NJKtGD3ME0WXQGBgo2gpVwwvYEoFkYceOLlLM8/uL9YBDZpYXRD
am7KJHnrJeJ0L+YpGMmPJ8kltuAHT0ZuXPc9tSbEKWRVbYYASpr+clOSB3NBSKmv
tlftPHeq7JbOQpZyexERvJKBHm4nN2RZtmqrivGmObgvH54KstqLERSSsBv0rHfB
w/Oi3J0TMvMn1ISZq8Jqtx3AsCH1mZGUXdbEQenRNyukao7pfydEwO4dB2Ck+fl+
a071XwJu7a3eeNBPPyoFdYjZ+/EGahzS7kufCtc9FEvJtCJNu0+v8TtMkTaYiE5A
mM/0Vqm/6MnF0wR4DwjGVVUB9tWfbialEL5LCXBEIiyklaa4AOJMQigvr+/tHOFT
OCxmgs6LWArSgr3bFUFymyum1edT+3ABTF4fLSoj/mMXfC8Z+HLB6c+s9Y81/f46
NTgzhzld5qACM4sOwGsFPqZUWFSLngbJpiGYuC+EYehw02ypSi5XCAg8tWUx6xwM
iXfMDgg1HwT3RQPsY7W1vqJCzOlLksqbBcF09jRcykGd+vG0FPMm1Dg+/mgFxYGG
hcokxjpJAO5kJybhYD9IKKI8s7O4tilHFcY6yxxjkwIdqpgF2kuuu6NEfOMzuRtF
eLKnlLtWzAM/z+LHncdOlvgU8fe7naOXnIkUOKZIwodrBQ6MDhMI7SHH4lgEadZO
+FPM9LZF+KUYiciy56XbrCvz3ShZBDIgPO5lm/J2ADwlZwoM0LbmlX01HzNSByp7
znyTJ92UHg6bOHFozsR2fsxLiHupvJfPHb1gp4SfmY99mBwm/rrwKeZCB8yQfahB
1cI8/epgflShXY5APHZP2RsP4uAJACUK6j4YnTtgK1VRzTUCJEIP5DWdcfSktWOg
jZ3DFHCloBhP06Z/TLF+zqk9DBz7ZxXpnM70T5B+8oZ78+MYTVDEX2BxXjZjIFlK
LaK6wFS5HB+pxbYdNbGmQ4dpoJsostZ0VQ93jLXht/VQT8ElNsnGP7cZ0BH8FCLF
Iy3xCDoTWQWNdn8HJsaRMnCIRFz1yBxOBmVcphW5x8l3f6bcJThDD4rZClXXs99y
MYWs31xIYa6EkC+TtZefOcl34q4kmCoHmvR9KqDWdMSTAQgqayVNvFVFkc13s2SY
m4A2b2SWIKLD0FsqN8I1X9OxqT4x/ZEqCIssg7WDSZpIupQ8+BL2Z3K9iqd87CiT
Q+yG6bY4hwPgTyCmUIqOmmJFzJU9hEljN9hm4TkbY9hEETVfMQK6g7z6R1SNjIrL
z4w2IFWeWY+MKkqRmYGqy4EYA39ZCPF0ujwfb0L4adflFFo2W5bKB7FmX7NM0Avz
NfL1TOujMawbFS7A2TXoslcDRlrjqGP5BL4gk8tpuaK0dQRLbagT4qDVBjqUlBzm
1KJzZxr4XyNrHhb85LUPrMrAnJUFGOqiUjm1mJH5LL45RTZSOh1huqa1T/xzI1TE
Ypzw5NFLhtuS9O85Rgk/DdDVCiP/s1gTQUjDH6VOumbn5V0dK7hTUIzEZbrIDn/N
5WNAylWUMiEMVpa8fugHHskG7NJ2XZznUzD9R6W6KHqlRNUrWimCd4J9jmazM3+l
utCTG1gPh/PqWqB4SThSbXi94JnrT49EnhruXxQjt+TAwE/A7Wu2zYmKzEuuNw7P
T0biN7z9VD50GAqFeBJJIaPdAAKtH3w/HBVkFhF0z9C2Vw2Hn5OEcSZZEzpCmCCT
eir5dnm4Dl+vtodhGQPGcs2xCrZ8ih3/EX0BsMXYQVdnwfSH1TtULD/bxVDOk0JO
5t2Ta2PNpXtqc46+ae24O0afJiBBZHh8/9jNKbY8TQVyvLA+DBKZmKc8/7At4q5j
NNdqxlIesnj3avG9wpdcavXVZWIUX/cuPUXnvEDyLIWCSgeOs7PrcSjTwltW610j
cqfcbsQgjbGDo5THoDsBrBCQvOqHbS6WyfewGD0kWVzAO3WFqlzV00IVRtAL2gxe
moCZTNlkGg0iUuav/1y6n6W6L7sW9vpLmtHREUbGUU8doHV4KkzhQpI2lNYTPhuw
irrnQsBnt2ucAnGc+RBhjIFtZNOKv+U7RoxWxANrsd+vLSByah7y41JcA675vJXS
fZ3cIEsTOOK+Mr5zpEnZqRu7plYuokU6SZfPW0ADYPuhU1ZeyrmP1DHhnZjGxAz0
d8OdZtSDtak3IMRTDCV7bay7KTu1BWwzrW/yNysLNONUAL6vclTLA4+bE7O9Mt3j
HhMmxHhjp/x9mpI32OUjRLWEHiz3FcMrK3G54qfnviz6W4p+U+5jydTU1QH1J1tc
om5YAOBD2XLnsiXiEIS88I5drnHBYt/C8An1MPPzfvD97EwsUKZhXJNVoPDtGA4x
a9y/MGr7GHpu82vg/yaZHKK1ZdLJXVUwAXmLS3Ux6xvfnaxIrpkHDOYsXHvl0hNZ
IbbWTKDwcLXAkGBeNrOmQ+FzIoX65Tsi/UzqvY8Eu4qP930h/fxHa4jpJMu3+npe
RCbK9QeYHMkPb+AhkVbBQL4WjiKZunrMJ8AfkAe1FSbynq2CDEIAB4XVGYVpGljF
47YnFjw69bl7fTzzRRsnoTvEjFIsQaGzNQ+//+W5RziDnmQhIXCIE4BUwWEcoQb2
9lUelj6b+Dfep0//u7clE7jVYqXFpNIvtCIMLf5uQuRyUJXrENM0yb5mk5YXwss+
wuqhnYXsOzXy5k8VcXQ4WOl4DpJCgm9uxNcP4HJalm/0VH2XDJjsnSydSQ1eOdl+
oWkUrl/uLNWlJKVz1a3O8E+CIW/2kntKMBtj9lNnaCiR5eWZ1aekAiyxjoGLVNry
r8QByz8V8xLkSKhjfbyzUu7M49G3R6vvlGbBmcdzSm7KBBoj+4sQ9/Mc+uOp4p0/
Uf7OAuW5qCG8vInWQgdDNKQM2e6T9KlIpg6Pa/8u7FlTym5bd4w9GYPan/+2N8Bn
E6xYH2Wpj1T8wruZwB8gMxNfcsBnKHiId3D8eljBnTkjhTmR7Xb/bh9gnfVLLoch
LNiyOHr8BumS3sPAB+2CvfNs8GNJ2+t1+l73p9pvY1LHPsef3mAKBUcHTk9YBgh1
PfoCfb8Y2eVvWs+WV4xOv8ferxOo9Z0jU6pPi+x3vDUO+sVHWrx9XTrQ9k+dEm3e
4mf40HcdwFdtLL2M5CD2H4FCBuElhgdC6oKjNZvCTQRuwM6oHbD+sRHA5QO3WBlf
/zaMmG+wqlDj5rjhveMX1JlMWeqLLrIpSLCSJFtZGlDa4BL523n89cOUbrna6BBB
JbpBJsN0UluEuRqAaPOehAqnvUWXyVj/oDls2OUq5HBwjfeUPVP8+UtCQpDFAAO+
JO1r09lp/JgRXOtOoRcbWKrMLlJLj/Zg+zzGWOI31mwifvYTDCK/nX4D/ypNt9cn
KpGV+q4earu/YruAlJrMjHPaaki1Hs8KJk4gv9jaIOqQWgKiUIQC4b02Y9dBqOhe
CVco7/svzaXbdZQmggIU3/zRHZv+eFstoodh08IB9UBKNcbmp1IJDVySjRBJcSX4
hGLbFqGLEf/gbwnkV2ZLttVEwpU9euFp8Estvx4loGC6wdV/GAarsA6tmwLyGWtw
QX4ZuNrkkgfSuzhrMyqPc7SGu2eTFodemPdaPoRqDpGryHJXQiz0+S+E+UxQovyY
ysuFWLQLBk68hoq/4Vg7FS+d7MxamtCiEf3NG9AEx1T8fs2DsqdyA1vTVs9kG14e
BvEHKLHHA1HLu15yEeKDmg==
`protect END_PROTECTED
