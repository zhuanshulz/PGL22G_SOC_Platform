`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BRQQaffoBuqK+i37cIQyMgyiFUKmg1atPdZH6lPQs9JgA7n4EvWexNkVRZBxnNDE
NKSwBf6oisYGgJH1rIYj69jVgfFkWISLLP52iIzVQSwH9gGzQ9a+AR6MumZEHBid
vVAcGQp2AOqQq+H32oc2UEYijPsf+jPvuhPV30qHwMmuIPPUZjL3r5ihYA+tFJOU
vSA3/P8yAdwpA1PA96D4C114u6T5FE+7VQHdxS7k1yzyoz3K+2jR0KWPp+N3ZUeR
BtQgccrMvDTWtkuVl9cstjB4/PuRubm1FERxIA+7747UhTqREkEBZx8gNaJzSS5M
rzIV48C5gxUjb6d7G9NGwOp1CA1SOVqs2jV8TSJ1U1GgWvvM3y5A1gN4EvHfX0J7
FABlcdyG8Uwi1OejzNiaHLbm46lqLIfAtZpPXvEF6tEld+iF664lYY03WtqkQtu0
yw46LoLKV8gSy9A44D9x1P1wjCpGRMglb9rmxDhUNBghTD9Zbh8hD6TZzlmLMMW0
u04tz90APnt7kXnubNhE3NGYq/Xmy7nP41lGx+bIzGNyxwf1eCcS3tsdkJdySNyh
I/OWtZ1myx6UXHXQL7ipABJ5+/TFtRXUs2U8+nFTuMxrWdfsBUIfa03eHKwUkw4J
HDJLHTFNDiVdWzr/m/MsVl2SOivQmHM2K7on+B04fR+E7EEGJdD1kuw5wpVdoJkl
Hh3UktEB1d7iNVoXRpFFgiiZFB8qFDsKVsJ9BJ4VXkHUuYECxL8hapc/NIRccClx
OKCsQFUkyrvjeNPXk5QpZC7gV3SRzbwGCdmAQXYu5oTf9wyPMPE9Cp5S6pw/J4xj
Q+bIirwRrJppUwx4s56ZJ0WPsHXUvE6uRiqrtqw9tiUpq1eprVKKQQUv4aKvxNJY
J2F8Nb3yRDwxnLEcVxOLZ/nKbH68G5fOP99F8cyo2PxrjrNpMmuTBWyd1Z0NOAWU
tLTjSNliiSSfK/I1WCZ+Q2RF+Ahdm0w1cowb1JHZZJe7ZDL7XSEbEmZOAqRVqaJI
wEuB/ug+H0SOsc66o7Owbk0aZbVDz5DCTFv8N+77l1GB5CwZd80/2VKHXN+9vu7J
VHA4gq7+yZVLQgc6kBw+emVlW1sNOoYcw6QgOqZiqxbYt99pq/3NKGmek499w6bX
HFT+oxT1Cuy6MtCCpvn5+rUR2O+1Rv4xA5UBuAzeXLTXpkiffxFEvPgE1tPRs3fA
AyY6mzXS/WrL6XTIQCqN7Q==
`protect END_PROTECTED
