`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tV4bdlNx5vEdlzb3P4FICUGxSzEePyYzBh8tFec0CdLa+hMEL2FdrT0/x50STnDk
HJLl3uj36S8EVkHdmPz8jdUkV88ZLR8ABjQgALJ/oHRhyIBlZnK6x3cLXSHUxYqf
M3GEpiK8oqR4Z57avpfX5KMk/xbaSXZGIWGCPwpE4SA4S/PU+/6XmOFXLAiSJYER
uVJNbmKUuvOnt0tyVUNlkw2v1Wcdx22/G6cDmBXzV3AE7fW9Wh8WM22fNekM6IT3
9aKQNhoTBvh46iQH6qK4BD8Akz5QAFZ/slvHnU+/kpoZyb9c1vlcYerI21e9YbM0
odNKewetLqyEyACeidLmGuUaRl5eXfUerWmkO7LxPJCpMrPmcWlsOhzIvhEHQKsZ
gpFaOR2as9Rdx8+R38nrOmNwKqlidvo6IxkaeZyA0M3/Z6icmTNa1knQjNUUSHhJ
yA7eSua34vGvCH2KRLX0kuQvX4OkVMXmYiL5hLhdGyxGnjdxYAqopVUobPmi/8Fm
FF7BY+4Ay7iyYj/UhF79pcVN9htxgJsOb3w6sAoA5U7+7mMYF9ZMcZHJqp76d8ds
npjxooNlQ6nopygNAEWM5HyhuF+B+rDahYGUIt1P8B+bX5yrCF6MZjqRn8EhQL6J
vfoVm0aFW+HPxxToridfwOoLpyC0GJ8RDGBTi/fzM9c8qLkckQ73tYsAMt1Y2Joc
nxNbnwrpX4n+G/rU+5avJJhczUu+B5pEBqIpf9zvgutUxXXZP7lEsfEI6hbIrnZ8
os2cO7Hki0Xl/CfSb52uZVllKsWaXtCfQFyQVI4opc8jp35DAthSkvWXU4NMb5B0
bk8hajsAvhHvPh+C1rWmF/JDISkHKaRNHs92GuxYbStRu5fWk1iCz3lEtLp5Pbs3
YiudQ0+C5EOz3NNHhJyUBHouO7P0HF1FDablNEFpBBKIBLQwMFwUo1lMcqCr38y4
NHDUud8vGF51HTxgBpdPdyWoXDoIoQtF8jzRpxOXFuLx1oF9uIALjKhl78rDfT58
47/aOlQRXqZZw8Z1mjiCzSyIdCZQ4GAIPVXdBKGERAD38mKQ5lbVZz36tR03SWgt
U8xff/fYqNS8BlpIVrGDQy1iN2vN2oS+8mwkam4zVwknAH3ukRx7KGfMpOpQoTwe
F4BE67gp/9b2feHln6lpfnufcFzxED98dgSHylE5kb7ti2y1CVvLV3eVRjxOy+2q
HAnYNYT5D4igeTejZZ0IEUnwMHn/ta/IYO7z8Sf+IqwHTWNNNU6A/XdGR9Urju8Q
x9OVn2iXOzpK5YQj2IJ+c5bTWfnh+E6PlfhDRLBEZcQ=
`protect END_PROTECTED
