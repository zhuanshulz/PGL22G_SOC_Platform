`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uqLzGjlDodMt7thCuHpF+uLP0gZMKB8skE6dj+4FR4EZ5f4XBfI0DcoYn+8qVZU8
hGDf27GdoVLfSnsQlA/5Eemran+hJSRF+uzmxP4bG4XE4C/6FzqbcQWjobNIdTKl
9UflGzNG/WiHwW2QoalDprRYmj6kp5xLC2rf6uIkWHQfEvIGfbiGqnnhtbmYVE1s
qGcV5xzrqF4BU4Pt1OgZLFj/dEjA2AbQjI4cF00YGEVH/HhGAl+VvHj/tnqA9F4R
wwlnJYMy926/Cx6K+XG4TZZp1ontXGjlnqBbsI1Dpji2t2c0beD//PHKz9THpZzB
iHKp3bwxD3Kp6eQNvLH4zwRFQSz4NXi5ORkyrOXNLgetR3RFr9FlETOSkq5pjMT1
JPLlDa4L06BKmXmTME18OJfZJverTmc1Dc4RCHyE9nZ6iDAuaqfi4yvQoQ5zQqrX
KfiqxevO+pqnP6UOzLwpatx2/5szhuEl0/PuHuuyB31E7CsqCvH1yvrqW0ourz1c
3BrF4NhGr1gbV5Z5ZOAgv3qTxUqX+QWll+kYxJSNXmPheKebTG93lA/yMxhey7VS
RwsF/Lhakd1MBrQC2/40mkx/wE9TseUrGUwr3VEl2g6bC2hGLH3thJoV1mvlGNgc
1WucGAcHgUqfltn82AaHWtGrAfzEYC5b3AOmYbPtwtqUAsI8yHNnbV3MV6dQIA7L
wTR1q81AVohxbW8BoQJQ8rHiHTk7DSAwzAcSjzf+fqwj/K3gWRWee7RfRQ3SNSWV
Vch/smqub3avJGPjy1sv2DOFNje7T/O3mYb8QL2zgpq2pjqCQo2xUU+kDRf3+hX/
mbzQ9hUE2JMoTJMxrY1DaSKdvJMq61TsZP98DgyH6BCzdZD0rA2rdoRIl84OHR/i
Fa4Y82lsuvHYFl3vbXkML3cm9D5s/e22xy18Axf/m/rA1+2d7SPPvcnSakh8V/lQ
r8R2P757QubqM+NQw3dSLwYu2fWub+vQMSxrtFIykNy5WSUr91eoyfBRUMgu25xB
eBggaQHqCDl8JJTXDnOECTOPPpceoOVqXNCwpqsY50pOi6yCevhECvsnuvDKrJdX
CoqVS9mi7wQZHR9JIYRtfBWuR2x4scewCfAR5NJHomzfAsx6jFhlBBL/JYuRXmQu
1w7xSZ2ubLngvatuiIlvGrHmrElTp4tqNsaeDMSYAnYpI6rxRNMJz34EHGK+yjnp
zdF1tLX9aLfJ4keCP2eJQSckXk0pVifAmVNvfn52UmaleqZV/xx1kSZeFA4MFAta
j8B3E1gxaoAreG11Zo0CQ1oHR8/GPDutRmIRepRrusKC4wXL1PrlHoFaSnGUOW2T
+x3xGheqjgr1NlAJx8KN+ZiuRBLyqNklvgv2y4DWH0dZ2RK3Cv67OxdU03IhWCoT
XztnxW3hL7yCogdKakqmtTjduBP+FmZbKhqQSAJPGs7a4BcifxtbViK2/KyOuR09
5svIpHS5Dp3KSt7kFWMVaE7Ai+8916JgG6pIrn2/U7d7++Drlh4traQHdhcM4/W8
CWFY6059Fm8h8xSs4d1QBeXjSFPeNMnHjtPU4Ye6jrFgjFE2jQuNiUOERtlEsDZx
24fL8Mw2TxWzfmqJDSm/rRr9brLMSRlb9l1uq99eRifbyfXsitJtB5YPj4RHcwnd
PasbhwwDT8wRFGLgLJ/cLHoEXzQK1nGxBoP+wJM8k+lcxNw8u5YuBdD7eVcJXbcB
xJIW8j7SpXlagAVQ/VGEaRtj4q6bffj1mgszsC3ajGODtDf5h5rzk+8fkKxLUhOp
uLQXwizE2b84KJKrLuEBersCDzHNKYdK9t+W+nT386QO2FIiEhqTALhDdzIqYoxl
MxNH4Od/5vc4qq3y69OllR/s3KXLMrDtbbfCna8hvWJ+yAhJeDBuwObNptvQrGFC
cSgNgWl7DTs9QM4I+7knsSyI9abIUoh4FEjYy7v+4V6VHubwNhFMNTuixVje4ylY
Ny/xDFH3XPzd7avCZ7nmoOh9YF8KJqsp9XF3HRGYWVqn8/eq8FzbS4EqrFEqRMtd
KD4R+xxELi4q2zEgBQWgZYAcCYTVWVnFa3hKURSbHandA2ylca/iadMGmnTTQQAt
eliuuSDE6EkWqEkBcCwtl+nuHULF0Le4tgWj7XYiDzhKrlcsAs/6oTt5pzG4tNSY
miNGU24pXi4hyoWXtsb6oA==
`protect END_PROTECTED
