`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qcnCHcL8AUccIKfDciNgmKOcEqOkQbZbXlhwibGnoFq+sWTJ2mSbX7I2XFXbJozH
yvSxxACrLUrAggRee+scKLF6i7LEhXQEA7Gtx0Uyrehx09O+IDhH60GozRdgbDiK
ydbj2i089YPvfLYhypXu7hy2T++F5hF9CXmH3qnJ7WK63+kUYjJC5AyDQfzwwB9x
5PR9lccNu4fUtWCkccf/HkYuJcsXCtyo5zmsgNgdmmA7o+pIUzS8BF5FwNH9MUmV
tVHFHqplFpo5RC6lFrhRBt9XzBBsipRNfmafFhc1lKP3mLOwJRVKrnzuCph08N3D
MqOD2jcA3rmYve/tM4jpwahQK/rLdyZmxxdpKPYRdYE6V49DgG3JyGgdtHkBmJlW
WiuGA3ovBuhRw/fddYuKpdrJvwH4TOgRJe+VZUf8bu4jrGwF70Uxk1Yun0ergUXu
t09e5QTywKZObBflFWYbRDEyjliyK+qS42wAfWG9dhDgFIaa/e08J4P4F2lEgsfH
JD5HP1bEvD03KAcxEt73M/2eHhO0wE871y1NGcwFZao6r2aqBVyL2LWruAkGHWOx
W++Pb97KpdED1c4wVRqhIy/eGQy8C3ne2nsLeaIGig2KC5tdH9Dj7x4ldKfgiRci
mzGNcxNY12QPaPpKnyUoYmhmEjK5ojWM6qcsjlWJWhS5c+kE5g3Wn59sjiyOKx+H
dPo1xQmkvl7v2DmQm2e146HmmTPLdW6KnyKHMjzSDqAR2cjRLvz2bS64a6niNlId
wS1teQYq7vK2rJ3WwcIrOOktsfkxshl8ZBep4CU9QPMk9+dqR6dRDX1DzP6fw4qF
/6rLNCLkyFs5HY0aaKb4qQDvgaej+UCiGCq3nctqqUSJzwWjbLMSWgsV12G5PEJo
bMJqQ+e8F7StevR996JqNRJH+b2+4LMfFlJ1H0OGAxIN2V/Baw0oI2D1JDy4tvbz
3/S8cIJ4pCGgeiiuIICt7EHaxD70xkfARl2On7tc53piZSMhslxeuRV+hGhHpSjy
QeJjFM8mlP6bOuPOWRr94hCZy9iyaLmczBWaXTVjaRJKgFzL18dZohDtq7wMSVAr
jlbp/FmPHeTlUd/H+UySNj9KIHNoaAkgGYYTWi90TuQQWVTA/x6K7Lh5oNAwTUww
K/eBNeI/kzf6Gu94tNNj3RpXAJ2l7S0CIYnI80fyVdlCNEUMGS3HCHeXLaKpytRV
UaL9b5CWXo1CwddchUuXcaqk6D3giKSeu8V56v9UHP+MkFQhD3ncVJwMml1orJJw
AGuKwZJRuzUUHPg5hSmhg1muPCmvYAXfuSpZQ4osjYi74Y+ns8cBGaapHWjALbt8
tx7dNbcUrd2QnNMQ6p8sKSbXXWHIPnmbDJzZ5pbyt/IP9DC+Te8VKpIYTZBcGe2n
cVjJ61XUTgvh1mIyquq+CToDK/qvgvuUUdBofpcvrfnQmaC61nLmckxBib75D5Au
3R09VMKNzn9bnsta0rrITRTUJflMu/QBes9x3+xuKyh1RIRifcqgFKQg8FC/+wCb
y6bC54KbVHd3QAujJhfDZbqzZQexUR3zBQ8TXrJbCV2F/kYThHuwXpohvGL9m+9Y
ecyyboO+PB1I0/8zFNkogBfALNuauKfTVVPEj+HZnNebOke4SvQvw9SO8zRF/MJn
EWKLMYJXY2h2EyXQwtF0uDOq+Oa1B40HEyPBJZAMoXI9u5nlrnYKDiw1h4ItprRn
rWNiaDNgN2zllnCpnY8UcTIMTPBmB7T0xQKRDcYRmPOxyNdPs0am6ors34Y9bglK
+IlVw0NR/OXSL0YrBntU5Lf7eu72j1gC1nxrPsOWl65BUAvEV3PHazhYlJC0ka4O
Z8/Ke2LaPy+Ej8W918VUXLTlvDNz1YXXDOAoSg49/2wmMQzBVuVtPRYG6Ck8upsX
Z2KHlpG71GP1bmnzg8B/UKKew6eKmnzaWkWcih0UWFqoyIQ0ENjGhJjuk31R2EGJ
s67StND08xqdtYw8xF2JaUoO/IBQsaUFlUeFPfPoZPLc7sX8GRBAaVKLnjN9VWEx
glTRa8FX7PErnrDdSkFdSQ8KM3n82TOz4XKxxsEWvkYQ1jHYlCXHbc/Odfp72Ahn
g0px8VFHe0HmunoHXUz9V6OINCdrwKG936HXpyETbQVQplQ1gZFJkxRUv2kniMp5
kM0Bykx2ML1poLJfA2gfrKj9k3c5otM1x3CuDdaH+LcY0XOdoKp+lulGDAtFDkEW
uV3LvEIIqoSG9tCI3458mbH6lzqk1QyaatRrKhGDaHKkmUMRvAHj8DPLhPaxcvss
JrZir9Qfq7pw1eV7laQvcTRcIHqtFhOngaBzAQ1rVg60hWKzIcC3Lyf/i+DV/nSs
qlGAM8AsHFDHNLeACAyc2+WG40vm7rFrG1jOV2SFsthb53uEqib5BtqxjyOCQPLz
QpiK38e0pv7UCu0NADmLVTKxqVOOCuAgXBPWaynZPvoIqlPmthDo2byYEDkLK9HM
nx/ncwUrz+IuFiFqpl6r1xXVA9EOKJzXGqNk/nf0jzE51vAHX+PUbiQEPzy1Fdoh
j6C3d7WIoLi1hhc6zCVCeCcHsyKzQp7NidXpLPQHqwqD8wXomFlI+vBfluu53yNn
tE9JjVnokBKBKLCOa2+8SmfFw7YODpuagQLMLigSiyDVsswXyAAJFUdrPYLHuPm8
Pcb2DvbqxsmkwRn23O8vAkZx97B5xJ1HFig5OiSiBd1BfSlmHWAe+ZBhvYrInSdi
6QCkbBX0JggQcu0d22QmzGxSMU6JaoRWsXSlTCe+MDDKAOTyrwaJjUmqylejgdAt
iHQAiNs/Je1/hzlm3u2hQmuVl8HUiOVdxVkWS1eVqORSrfPwfbq6pGRnccg0x/SD
a9ROgO/fJnhQcIOGOXDyEzzuLw4UfOvt4hZrlRBwpr/5E37fYiLvUEc8O6MRoSTQ
`protect END_PROTECTED
