`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ijo9jqGRVNHSHjzHP8HwHmRIuep2yAtNp8vZqE5tEMsNts0oFGvsxZhkChSeK+bK
r+GvVic6mLX13vA+8yKdtSc5xONnMnY+hVIHk4ypy4jkHN0s8SwJYhY3jPZ3qs0G
5W9NIvLRczDUXQM5X/gXCd8FliQtKJ2ml0QtZTs7GjzaWnptHNBB2qzwjVAM9kD0
Fhr1q5knJ6bz0xz+8BhbUPZZ5GggfsbCXTLaT8iYT/IO8gOyQUWL3G+yhrNjEJV0
z4wAs0M8HaFyK8BU7b1MsA==
`protect END_PROTECTED
