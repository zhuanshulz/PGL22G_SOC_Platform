`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7VoCmtA1RVXjQKOAbqEMZz6OpD5nCtk/8Wf6gMBlj3O5lpo6fudTX6gfYaYZpulB
6wzk8skoD2TRtk+25kVtgMKHeffTf0tIRa6iJzJntie5ecQaoQN8+vj0stmbB3d5
4drQBCDJdyGZQctIOhCS0DkcUpx8ZbNcR9LFk5AHw0a5+aYO4ivkkqXjAtvZqACR
ZED75t2Jil5JI5T+9tTTEEPsfdngQGKM3As3faxpe+HH6+vGvq9K8IEx8ZUWlyWv
kf77rG3f5JiwVZcLbRAGskoV33W6vJLT7dR+1FHt7kNmjVcVs5IGeWW05cxZGhhL
67Hw1wGm26GtQyqD9rAKOAkaVLPLCziEAOYxOLNE62+CUJPcH+FCv5zoTboHGAxI
UqUQiXS4XP9gR3dHXxa2xTt85O0YHhigD9qeMFnfWunSx7GO2xT+LA0D3i8///Q6
GsH1BnTGRcgcp1uItJBQ2pMSogQ7WQ8ZAe0gZQDxEtRUa4euVV7MJwsTOveGWDH/
Zgr0iWXu6pMmbVGLBh8QjYR3lZqd7uTUqFgqHzbkdocZL+9XRRT5PXffAx26QM69
UJZPQK09mfWmRAlS3o/z6pKiCuD4farIGaFHzp23sl+w7tJWx3qC4ea3kZUi7O0P
ZzdYFYppBcl0CiYFQtd7eBwypLV4gOPcS0NaRXMnRKpjvCGXuGsleTwqTMtmTmfS
Fumt6HsAfASpNCmW8/R/p/2vGgYdyVR2iekWcbl8d+dpKjy+yq/Wlx7zTFiLfDtJ
ivheXJyNfIHqdVhQ6yL2sThJI8EAYui3t+Sm5mQrxSvWGrDKkK8cCnYi5X1aIKum
968kthafb73P4KrovlaQQULk9PTtnkAoxpjTrZ+bFP8=
`protect END_PROTECTED
