`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PjH4xIevfVc/5L3NUzZnC34fcTyJAXcq8sLwKzRC/Htp9K56n5wmiTC92KVTZp7b
eTInbowX8gP8+QKwHIkMeJ1zfkUWJKQDXhdOhyzN+iXHh+i5UX3JZ7qSlfX9rt7I
0PVgoYcUGS47FJiotxCh3DhfrJhAQIc09mfx2JRPEFe1KGV3rH3S3jexvsCcr82X
zkxli4ZcFw80Z4/XV1ioguO0S8LMKO6hNV/rZiWCSJNoyB5uzFvNxNNv8ZDbR+Vo
criUGDysNal9IZbI+gAY5IaZsYsDsaslX0zfnCU16Apvt2uLLZQxZKI6h7JW6v7z
MEOffnyOIDc6zd7BsrX/oLLlXefTsMx3HiWb1Y0CFmi6Bj7rBpdPoBt4eaglcbeg
Wx357dGv9N7vBpkW821HlXFku0g2pXAIJk3vRlvfvdrL1loEY1B9h4R0mzTF4Hk7
viIF4GCmEmpNDHiLDaA6PqLPYEhGh/5wZD6ykEJo6wlnadmUD4144L518JjGEz+j
leLuEgW9pzIYLq75khtrBqkYypEcBqUBmMzWG8t7V4iGMMzHDGiPlW/u1+35WEkN
KPZ6L3Jqyv7zlCy6a7GJxx0OhVJV5dkKaWxHNzn9p5q0ilBrcyK5UpzCbTu5nxNg
7WAxIO1UMT6rGt3p08prpnImm+8/5vdxb5kUOtJLqVzJQMbFnV+ZmHsv5jy4isbH
JzmTfdHda1jLcErrb3X8e9dKnk+Hak3EGAR8XBhcaZESg9uafVC3PMDO9JKeAUcz
p2/tQwC/XygN+aYZi5wMxFyA3ZGYlX50mTZJoEdd9v+cbC7r58OGgdfLqyhkcbgF
riTGvYnhB9CokAD2/F1AS03hkjZo20Aeh5kNw4edfOcFXbXqTnnEIowdjynVGZgV
FFKhDyWrlaIXQ0EYUcG4pFRelGfeezF+5Pw1B+HnqTRoHzzsVl0WqaMHgjQMqZHV
tVqi7PaypM5/w77U/lymFya5T9/bnTKAj8ttnueJYVpvsCshj7OeHsQV9ZHBCt0V
055LeFQGVUgUJhiVgnEyxGnfhofcumdUb3ep0Xuk25iSWhkjeaNW+f4wc50qxKcg
ZR50JErfLrtLRrvtZAcfaVGNcTm84sE3ZL7uOVGCHF8+UcnNPiMO9PsXX50hRcd+
H9gCKxlX5/ELl6DRFfM7iVd6Ti85YfRFpCbAMv18EX0mpRHUH9eZtDirC6SM92OG
tvoAlgC4IR6U8Vs/2McxzZrHOuY4qjDp39PlpWSDsfmOu+gsbtc8jEVt8PgNrLTS
RcG5HpSnxlecynpHmFCSx8f17vrl3A6ELQrN8MA9yxBYMX+o0v+SRzrTtgbbKkyv
F9sDesHVBUJWXXaoJneRGN5TAFtBUDZJKDODnszOIs9JIQk3V71ueBSrXE3NQkfD
hJZoYSRd+zXgRKV14AUlu0xaTSuJTZu67e2bUUCFkokG3ZaH6+TKvx8S7uNoT10L
Jm2dvuIgLFFAZrmt6thUh/3zMfU9KJpCOVtKPwbZ8Ywa6uu4G/jIWLeEqYF03LeX
WgjeOqGl/CgOqy8/yK50FjgTKEbDhJfA77DTz/GDPHMR6JyZdRYyygvboouNG/1a
b+cetW3SoZ7plY/DRbe3ofF6RtokuJREKVU3F6SyfkY=
`protect END_PROTECTED
