`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HFq4HqDjgUaay8DJp7YWVqJC2ynbT3isetgeKhlutmivwJvkckOV4NoNGU+KH3du
VFeSPmQZnL8R8SLi4xIEl95c3ppP6diEmJ8ByAxUGbFwDi7DpweJAYJAu61J8EaM
ICsJ3m9LzJgS+HqTDJcBZcWM50hBPKo9TL0Ma/2/RNhhHnA+SSI37epx0iD5cSyo
hxU85WbelbvZQTNPlM+z0h7oyWGjfzaGVyoKjDDtGa0+uPShD4r77op9vXvW7UMb
h7BQuKYPLmXagPkGyFRf0iS+5zcNBXFncRhi7MrmUSleBpkI4+FlEI+Qu8MVSj5K
JDwLHb2C1t8FhXHe0L2+JHZhaTVimZX5rK+/nto0c5nIGbo9rME6gcy1x7XJxQxU
7MiaM5/UEvKaUU+051Grsj8Ci5hf90xrxM2iifnuM5Z7d1GXqz+jtYEWViDQYoRG
Bbx5wbzfPFFobaKwr418Dn4p6E8+KfmACPhtHOuuhKOhJtkwwVM9fl8eOml+IzwM
ohqqM6UUCckkP+8i/VDsJSeuAQrkEAr5eVnDO9WRGWPPDvEY/FZt5EgIUkXwxIlB
kNpAo+0hnZ6z5Nn8XXhvBezN9QLYma8CyWOhRYt5F9PsSwE7rE7sX60Hrq9rP3vE
CyFCl8xk1HGSanT7VUMmVYPiYz3Bg/Wj4xli9v0zJM8w6nQltqZAYTD8WBdSbpkE
1vtKM6Hu9MychjyT8aHmDVLJcL2VdF5RdUYC19coxjATbkqEr0xWRBFaDCZ+1U5z
SmVT3945FdxFIbMDoN9AQBssJhiNCeLqgaGojBikvu7x0LR0mVeof2lscYcY17ag
3eAv5BFIAEHDkl7gPzwK5IV1jgNespDaMlHVWT9BYxyQOuDqEQdfGLZzvvbASEiv
kdDCAKDEQQcHtadUZl8un4JhoypmXezJKMd+aFfRTv+GPiE9HaFB7SzxMKc1At4V
aKp9LNl7TS3eNh2xzsDxrzOdyqfvJjIXW9h8lTeSBI3BW0RoIarpjbf90MgSxT5i
w6fgJxB7aonG3c9TwbCP8IMQJsqpUNIOKcLbYgmtvs8C9ZokQhx5IpS9qe9PmuMA
gJ9zNybwNEST3cO96DQ+1LABuBqmYx5H9bwJ9Uo6H5FkwwW2/6jBR38NbBOvk5Y4
VoccL3KkqFlIZA9KuJhkYXU0yK4cC1Hr75o6uazdKtUaa8hYRum7aKyBQP1UOW8Y
JIW6IUBJERq3Ue6h66C0v9xbdsP5AsF7CDEjvBqhAqTyI48vi8QPbY0i/XVqMnix
S+SvEgmNpxF624PxOprcEbfat71EQ/8budS9VLgK2LGjhLqfWme9KUrcBmSExvKp
Yn8X/XDwvRTDjVCv2cXrj5j9PhqDHEjx3RiGwsdAAL4pYpC9nTPN3Qp4JaQRPxUD
WNPuGIEzihe4axikRZ1CbE2bjw5Ugxcoc70UFYdqTXhnyj2DkU8Hg1ALhCTLeHDy
1qKUgaWn+m1mVttAFQoI2l1JuPvXJGtrj8d3Hf+3jCIksYIE/PDhba2Z0ZW0f/WZ
sZ9nbeY799av7wYgXBEfrBEvs7XJfgmeh0bytq+UkGS5GiCQ1Yld6z8ff459rXu0
9xojb41MP4QR+YNyDRVmAdGlSnn9q3CE2XH0Ug9/kF0XjoyhmpHmEkVNzThko6Yx
/lmlBFwoSyEMxugCo/Y6hw==
`protect END_PROTECTED
