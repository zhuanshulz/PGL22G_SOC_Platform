`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2aZ7xvZt9L1PZgRrCEFQzcncn+ntwkXxa7tMXn4EmJt61YR2YhQ28utvTG/bFM0V
8pfPcCyhpB/8cWuI4PwSMWTX2B4Cch6nVL9rO/YNfnH5UZpdSn9ws80hvazwfB8l
tvRZlCzh1/d15hhawGgnu+5BiJ5HMJBcEdJuZvGSCiepmp+YFMYJOpXCeupxeGdx
Lr3Nh4LQ0qGp7+E9o0hNW08SfFhq561sHZlsmVX5/0jnY8sq/Vpz2FFX8uNSt7dr
wHcb90vMp5qadVC0K7dA6Es1rIrsgvnx8IoHRy9PdmquNETkhU948l2q08DZriy4
DKjFcJVhr6HRKRqCOSv1gA+jn+y/A9SnTzfEhdAmpSB+Qq6J80U8s35FbRnoG7RG
NRWBTlyGl9NQ1rqqxTNQp7mGZl2UaGjQc2opQTCA7rQ=
`protect END_PROTECTED
