`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l1KwYqtdjveDk+4Z3pyzsV1B0KTIxMSpHWAOH87ax39iFjYDhwc25HqgEVi4Qd88
kQ/ivFUfSfFJdWjgo/EHO/j9KZvsXsBUdyOrnq5fQvKfY98wCFFq/HdKKEoJEjPy
fRCY1JvLn7GGf9fwoRNOcEiA+dRJFGOdKp9n2Sa/qp751k0tXRsnO1YP/Rq66CM5
R+6SZsG66Ha5voubn/Ec8S/LVBhCDE0XC1bPYvELe5yLIxNsccah7s3VzqXtoCA6
ZTr4y/WqY1+MrQMj0QIWU16SNC7A3vfu8kunV+0DRvyXvRIcxJ0c+GoL0Rr8CvYx
XPanUMAXSg1CWNZuK+EkrI2AGvdb0SVY+3+5xAkZcS+lDsFjFPIVAbOOhX/rUT8b
BPNy9LAvkF6NPAeDsxIq6I2n9jY6zIsNHRY27QprS0fCqLh0b3RJTUNmYmnllEFN
FbRhHGR7i1tzI3Rg6dKOnJXsvZCg9gPO5mOzMBcu3kHqYj/lDZ7fw2C7fTOXAwdH
OcmZm6Tm7Dvdr9wB+7aW/e8SwUxNzjvjygbZKhjRdLdh1Dqcfy1At8x/hPNLToMU
YAcRsK3c3mUuSFu6HDioQpwiAl7B3xELLr6SRDO3Xu0HMX5oEAER8eGikS+xOy91
1NiIZeSk1MY6X3Qy5NtnBEDL0MwvzWSDs8bexHzhptZoTiBzjJNOamlkw7zdo7Bh
Ih8JawWm2ToeR8jWKUAofcZFk7KQOJewXnf9QjPjlKaE6RaRclHobGfkvJLQ2/Ss
DDLPpIPcujP0IltHqkbvGShvzOKjWZzmevDmB3nqfgyQxmOyphBeYu4E7Rf4uWEf
QAtpbe/OX2hWUWKGli/y7P/xviysDdB/4PHS3wltmlLa/52Gvl4Q5GOY0jFfcIrj
NFWrNkY0hdBgDZ0YYeQWaq7Q6iy8erFeu5gBh04SsQzwpp0jyzhfOaBIn81tT63Z
9DQcttZP0QMF8c5WtmmU0qwmDmFlvkvsj2gKSyMNjaTW4mckCia9E7UVaSuCFRJp
vAeg7N73PHoGISok9hjlr7Bm0MKoBK+yLqRdRtU45HnlE/KJPNun7YstYQjjnbJb
eZALEY1u3pwD/RnFoMDcqNpBfaT+W/txj7okdY3yCVosNIPVYVuoVT8XoFqo3ST5
HelGcQZANc5pNOTQXrHdRLxwGwfaj9xO20dUqKH51v6qNERVKGeZ7OtLuVhgm6pE
U9nMs37vb/HZ92x22y/cbeM8+Vsu8az99edORgVMEURERm5i4SS1DteGjho+bOzH
MNzHTh7OdhI7ItFFLg+La0TnLnNFPmEY8nsRS0BOBb7BYqBPyl5PnpxhuUoAobm4
oz5575HDKGdhU1YxhkXH0Z9dQdxBax2y81P8bBLKAz1sLAGBBK1Ihuz1JlVnlojk
jZa9JOgsMoC5+r57Ebj0MwRWvUjuufWNxfIad2nsbckItRNQWrCCNSvLZx+THo4b
zkUDMrcMwxJbsRFjgLkIa88HuIUaZGv7tFXtU/c3yobHwJiCv6IBE7xlOinOLUk3
te+JBjR3BgMstpzyKjmDXDFNvgByvzFn78uVyQbmrm2DzANfTEXFo0JIWXOVB6sK
o6GPmNdUnS9QpyB8LdH2wADui9N9rVQTc9r6mzyIa2VzJJoVWG/mB8L4aEm5TYFL
GmADrDI5qWuaH7yO9w/W1eKMsifNwFo2ZXK8OUVC3Yl/0A9b30rhVz/3+ARy1YM1
xpqOWlhkxOIgXUo9eNt1gv8rM7UUQbg0zXDtgzvYNVVLUAOIpFHJcN8D61OVcE7v
6ceuPngptshiTXN2NcscPCCoZ5kdnKp48sJGG5/CSyrp0Yl5mCIy6zNNjjR4T66b
bMBMM32r8ly4YFcbUkPQef8w9vbrT7nlQEC1DisjQc2MWuo1u84VhMrTHzM5nFBp
JyuKCWTHAyEItWMRO97a3dExIcBa5A9GmepUZVBAC9SVc5AN9X1mfkWRSkjG9NrL
VcSuxh4mecSigStElMCC6dDr787eTLah0kmqO2A7sHn+KpixEfSZzRGTYZsELh5m
gvYaBoOkh2VCqjG/nHAr2JrEwXSccZ5cWZ/F0k6YoZUqUGMVGOlMdzmUhTP/URdh
kbqE+V7QrgU1qmxmfq2vYz96nGOhfqIVj1CBG342dtf870KwaRnVLj74L6ssfGa6
dyuj0hNlqHIlUi84dDbEjDG72WKCU/9xlV5oNpOnfhXuhgNSz/pEziOP3pQdsKvP
SLr7s3L/jpPXJIQ988SrzgijwEZp1inku7xS3UsAtyZUXHHe0ykTC7HpcllDjRZ7
cIgVX9VvQtue12Mx9LeXG+WAByJ2w4nIRasvJkp/0z1QiaK3o2GiFNFvSf/dCQoP
3SHtKu8JpwAdJI1UKf6xJg==
`protect END_PROTECTED
