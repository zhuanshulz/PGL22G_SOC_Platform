`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rpv+3bT/JusxpP1U8SM/12mffsQatbtVCfF+m6snAbjWyxajO32T/gtYw5Sh/XEB
3ItXqSaLIMIg3Erd9xZ2flBQQXgLfvvT2CWvX/voNLqrpyyQkw3gvnWoBnGqi5Ek
YzbNk48iBSgyjlGYfpWIdQhu42YO+636uXqh0Nb32C0yYqQaTJVXfTHe+VVrVgw7
M0EHoH4AU03ibFgikm9mk15SJ50oHUbhD7WN1lq05HgtYfmDatPTnijv85P3lvv5
zERHVlrdAXFyTibfn2CG9HNABMBpMvXPF0mdvBRjvL0D81Vs2QdVs574gymiLCfS
WrQEDwxw0BOcOZyzslhJ+eUdUQnDpTUlBJY/z+Hc5MNwD+jaxn2jXkVjnAArebRJ
CSwjIsgdmV9VBMGD+8t0DvalqG0/03YuyjUW/fx0JT6NtPum1Fg6JzHYsYlHgP9Q
3TKUASvnC1Uid8w6+/lglTTF2mi4HIBvH+D6sZv386ygVK59M8HHTPSWZ03p9sz7
qhQzGJeofsJJCKkMswaZsaW90wed/eENB5jiZlHE5xfjcZr31j5qpLLz2CRFzhVi
MzM2ZQvWF0b0kqciJxBmCV04zAHwzVl5iEf0rD3TbonDEpKzzWb3OU9SHRihWWX1
gXwG74JEbgawJ/6lFlad66Q4wbmtMHt6MITUkIv4ql++DCZ3+uzxvP7ZEycIkVHE
cFNItMb9yoYwsNNsN9Zjs3QBxOUEQPqgwhXgDenoeYxksoEBOGV5UGVxWqUy2trH
jZmF52u4hgs+jr648acEkuSSh04V8FhLVj0UDFEPXlJgeoeJWSEZV2QB5YZ9OsEz
O9wibatbsjS5m1FqdUq2/qcugbxEl9qTxeDz+kTf17MZ3Nk2McwthsB6hBzBmkeT
wpSgTxfztytC0FbAzvyzCQtOW1+IOJ+fZm7cxLTvhIRg/39zpF8Trgun6cUSDU75
vxMYmYObxmsAGL4a5wXHIBjTQiZg1wIN96/AcIJJRCav3DGzioZvRt0vTY4cvnfC
BzQ5WhAQ10S6wHhxRoEvnvmqduwWANDiHo1okF7k9VAhTIfCtiVw5itpWRrVNo1e
7HANg1D3Bi7sd0O5rVG1xkxR5w4rmqaRwVaEued4CKpvKiE6bLYqIjWHHFxdO+im
O//AARd1SwPGaWNJ2sptFWCBGxFRNUrc4UdVTOy3Pu84KpHoO6pvsWW5kR6uxAtr
cZ1UlYz2ecAgWGqGHSTK8KjxJN0dneamZnV03y6DwyJXcnQ65jX86a2THA+OZmJb
E8lxUPNuwOKMi7Vxr4uhvxP1S9rpimKO1aA0nq3D8erCjgauwlZMzpsbmPOqqE0n
fALyGEU3/x7wfwA5ch5GHdnfM/wD92iOk+uYWXiyXLhy0tDUvBSwganft2YWz86x
jx1uxd7PQPZvj/FWEZhNlB3AFT5l08tbgBn6afsSAFlNB+3QiP/7Dkmnr2+6h2Xw
H+c/GhlSCgzsJgVoUFZSlQzKCQTHVW04qdJ/ZdiDD6W2wXfi5rPkzi39XZ073PtC
iZ58D/jticI+e3mFmc8Cc+3zqyJEbRDAH4VdBG1L83zOIzMoHuI6NQb0HTO3LRN6
7/a50psOa9JBAklNvlX3lMI2q9Ct5gAaCph3/FKyp7p9VELR3Im7dZTO44dS8p4k
FIUCmF79uyhsXBOd0kheRIoYs/ZAgfxMpaPBAjk2XCRrxp+OVe0AVqXTWVIlWbCe
9gjaoRbN6ZjwpppMh7iEkWNFIlbL4qw4NeczRwJkuDJGE6nfI9rkz5i7gL6BLeDu
06ereMImHbzojnZVZ7KX7rc4q3uS3laPdZcldLifzNMxRQ0hUl/fYYfhuzaIDZY4
Q85w3Vqyl8HBsz8CVV/8XHXv5YuaDMkW5/fBZG5/BZYYjkvjHP6OwSwTJ6X3LLWW
cwl4g6fCqC1RNrapUbutYzuEeRi+kO/TxNoeWyk3qroxuC/LrEHi90LbIZu2tTjc
MaL1N9Cq/MqTcsB9gITjveNaEH6N1JTqfEgPlIiVPFWAM3hIZJzTtPkEusPXkqpq
eTxJJA0qKLeJ6ksMQAwLrSlbPjqO270Hmxfq5znvXdbrWvkKTcDq/L7xzGPD5pzp
/JQAIBEEe0c2TasKmjAdQB0DDke8zBoFUe1VaEUR+WWIwxEtiR2CcIGfaBuIGGyj
RolbMHAqalwI8mnrKbwwqqDd6Olmyeuu/0zhQrzymX38fH8VDNSN9vePzLad8QNF
Y50NTGTpCQ81r6fsqNVezBdVvI8leQ+L5g+gO/WVilH7deFjJ4U7Td9gJEu6QQEh
5bLMG0yERvIH0FA69puXY/3qSub/hW7/rCL0iAxzUpqF1D3uhViNxlsVd14ImQBw
I7HJYKHDlJE6XBP9dVbnhq9YPGj1awmpL2lVdwtKhzw4fS/VQqJKo17xO5M2tmB4
sooxANqqgyGTb+Qb6ZV7HALjo6nzqjK3SR8PkkdcxVjflauIcE+CSoIkSk1sdPXm
dhSkVDBEQooh8N4wp+sjVJ2WMbqzvlHNTS7TWRvtsAw141D1x7IV/rNuEPahXvHV
xhct5X8Wm5JxHC2dtqLDtGpnrzgXW5LCsFmc3j42UodkbRaRiMwso1nc0eklAZ/y
J3kFbgyrUhQa+bwVoarbM7hCmrram1a6dB+ZCfz1/WWIhwyT1+rV3UvoyNgc5v1q
Q5uKjqZNYKIgFqyrgSrH5MeId2mfKG9OSLnh0CzSmoMW+rVzUsrBTFHbl5JgWZj5
KYBwtLgeAJa68hzsD2tfX9BPwQh4Lz2pHQUgxqrdw0szA4JIFGShBGB3+HY0HSWF
dEkUVW1QNwZEOW6lqhyTAqD+BMwfgCzeutNOuvFZnlg7ZE1w/5mSFimN5lUGLkyx
lrsMVJx7PGOrr1C6FSdeG5IEzhs8L1uA/rJTavJRpEcwVbqAEO3T3nIkfwHTs2Fd
u/6+/5HxuibaE1ucDolB5mJw0okwzDNYvtfFhlJEhR1+NpEF+locxXI+PaiJyJkL
0X71SKgUJwvsF2PTyI/oJeWzsDQpgzFSYuGbYyDU+qxKl5C4qCA/VyJxxRjjMbBQ
vuSPCpOtuYYG0rjJr9yCxP117nywCZHoWstCwnTM4An1T2ci+f845fXOqC98V35t
yRd1KUdtm4pMll7WH/gWgd3w/fqkl0/pftiQGOk3i/r93OzgRJAPJBepdRgJb/Rt
mTCHc1h5sJb1wwx+eLqf4nobNtPrvAYhTLf/IlBPm4eOiIPeNkIO2ofdGra2VLoM
N0BoT0zzNhXZ1vLXyS/GhZv2/u5SkhDbSJzL+iKs7L+oFtpbAv6m/1ZkKAfOSGGS
XZBWC0JTmNGdI8N0UAta7BMmGWVaJQl+f0f6TvMOSiF1LIitc8WKQwMW0kU4lfNz
j7VnWDFKVrR3AjkZ5IcGz7/aBr2O8LLt4pnI6KW70nuejfhPeN6O9Ex0I2olRWK+
x/avYxjDuMKd0Tb91Tt0Lnfw/VNPl5SNT7iS6zAWUanZJ6da+2LOSyNvKZ3whSMP
RTcX4CU0kvxq99HVDmkFamUtGkqK1ZhMTYUNRMYKI01ECrq2MXz1rqGvRUBLKWJi
8x9vSfcM0F0gbgCjTE4pNRxZA5Rgaok892L9meHBqjDMz2z6RRiZuTEkKSbaLP4Q
UUOgW0eP8SSAaeIjXugGfee6ek4P4veBzLBZ7/XdslguZsbwLvz26QextVbWI3l6
r8JayZBL4XARbihBo5Z4bvnoSCeuhEBA20x0/BIbpiiFOC0tnG7y8hYo2xf7Li7R
RHQVbwK5JfUGiqgDx72IMy67ikU0uak8U1XM5hntZSfO7i22YMsbADbSpIm9tayX
M7vtlpa1QAsHgzEfd8Un0hazBPUGyTvFuNzSyhG7rmp+zu/MM4Ofk/vHHiu4kao1
IMF7U9cWM5fVz+vF6VARYvlVbPx4rgPV8fNqTfU/4Ir9TldE97phvZlbKfpnhtNo
mMBS9RpdIxGnpZMKMq5To2w9bRZBYwlvCYZrhyt+XdohzkYLqoGeff9vDHExJc7m
xsVxoUKyXY6H7dDdfPO/XrPD9hoWKecChVhBWnKHFsqTkVGMO+gdOz+jyhtye2nd
uny5w04HtHwmesp3h4hJyB3ogEbVpRIH/tk15znYfLsUU5mk95VuKrgngsCZ1LDS
OW+Obw8pQDIp7HjYnHEdYmYx4D9vFiKUQi0dJtr4LycuDA59Q2c66r+kbMHELLay
o62Llazq8tZpOJQrmRFCw8L4XFg2BjMr6sS6TvtjSiV+AqkzCWtKMh+PqPmO13Dr
Dx6wRs4eabqfEECpsQsp7NmkWOAqZZ3VddylYmiL6lSOXrFm1nk/t8EOqCGQaKRY
9aR2amOzpYgUHxVqhJyB5i9KEKNP9YAdeZV7npRIfHDgA16m+0QL1fMeAAkRpw9Z
tv7pqSiEpHKZyS7KpwrlIrKP/9HMdXxyQ1ZzAuwnpoVARCTOZ0mma/HQeWEGrk1W
06CwmYmwQ4QqhahDvskeReDxLRLm+FNyjJNlzYieXEQpdTwbDSqoLuql5O/W1fSe
KC0VEyLJodw3oZTuG/HTOgfk/KVGrc457ZKhxzHnZLCadc450hueTKuX38clpJEj
lx6WRTMZqrjKMHdYHEougVsWeVPU8tf0mUkDmWg3+i+VGt54pvH00GBtD/XRbMR8
kBlZE+Oz27b+pgrDtRty2/VWDX1aA1mwcBcoK3eJbaHYK5GKcevAz393DvmT2XY0
lXoeBYw5tAwRa187AX2jIvibHlyAyBpHkDVUsIMvLZ8sj/JZoukeVfjTCMGUXF6O
90r0kGJ0oIhFT+EcVT1LAbZYNDD7x6pnOTjsp8Au2j9498rfY6wfsqN/xo4TgCjD
vKqX7eA1H7e/MU52y93erdbt06/aTOWdUf3tUQe8BV3+eSoRpoCEn+Q5ZHl3CrwV
I+p+4e51lRhS6SI+s84FGw9pB0+TqHllGJ8bHyLeumpyMhGTZyWLvpdp4Eb6Tl8p
Xpt/M5WGU9GG+497CtfGe+3kAdSOVIzmjiOMu0Fz3G5Q2BrCk+cx9F2cwCDH0Sdg
uXpOge1JBlONRnsf3QsYjHzux7LMTaJxzo3eExkMD/zcHNpTzMkMy36jkJPhW9Kp
H+yqa+OiHZ+8nn+dfY56tKPxDAaDs9XVYInNJ42rY6m0jGTnoYqqXlShgGR/gHW1
sgR3YkkifjFqGe2xUtzsqspBqDuDyWUjbbHHNZXbOnXqam7B08xpos2eKM2rw01c
8ISt27zk0o2EDfubYB/Gi+2jkCl2p3EqdMn/ga1jiBLSsqqaQCnQrfvRBs1ppYOr
UDTJm5R3FOqDKNUkpuE8+kLe5hz7y8/uhXlhumsLSya5Z65NCSwpPRWrjg1Jnd9N
npqlDj8ooM5T3j3wi0Qlt3gNCvauJmx7s4rMXzYSNLBsfEMJeHmn4ZDnvBsuQwqZ
zJR1blx3CE2sFkC8pg5FhiO0JUi7vRFso0slOO2bEqCOfmaAVY1LpEYoWyfUgB1F
G+1yMma7VN6KKYIYUcBDwshPn9e51wXbkhiA+5sy2p5azmc/8q+qSht2xCvZypwK
B1b0MJe5G/hOb49kvcKSttqtcF8EEZhXIxAlQ6+Gw8mg/KMO/kO0R6j+Mgnr0sHP
IumPV6ZoptP6Go6l63dYZUxWggRZfVkT26IbTuvCcFegXSPYX+auoXwpJV/V5qKc
tgg51TYlYxhK8s+QvRCccmseutG717jnNE88PVmjsLipModqhpT3tppgqTqRcUAW
lTTnkk+9PZTKyNa/4lJHDBRCiR1zr3S+3mG0//Lelbz7Y5kPkkYw6Ytq8BcTEG6l
c114fmwZgjlWns/Lv/GzSUjy5KPMhKuD1mrlYkwczJZ2cOb7cJNuf4Gs0/tgM7br
oBSUNgF7htLWvjX8NkbqvuIQtTlN/oeVu9VYfcu5aETNsseZpx1PaE9G/nbfq0lw
PJ8osy1JuSy551AdFYxva5aXFqQ5q1zhTNe4kpo05l2bz/H6OIDsFAPI/f0Q1wzt
p43yhDONQsCUPhlYWpY3F23lMIg9S7HLh5P3XqReV6mMlvTYAbb4YBY/tuVaOvRK
fMB+I/KQOuaNPU/uJhK7JAxf2uHYTMV55Mk5MdGqx442tG+Y9Ub2aZGct00YB64M
olbYHXDVBgJczQ+aVt85bQF0NRIemg4FavGYETpa5PkR5URKDRDp6GAD4gmb2h9H
vHxsuY7Z7wf2EciHmRzw+dOlkvvyn6x0tW8AydPUOOX/CdGvMGkbyG+D5ZvCCyxz
6lTXA2tQ4DOP5do5U3JNsdpVDMCtfuNlsXisHXYCoSid7rTKvDMVCvwpgycys8yX
5rpfYeq8qOaOAq7bGxEEsEVxnqWjZkchmVklBfsgJUh6dQXDIBqnhcc66h4sC+oU
5sNNErKzSsFBl/WlvQUIOBy/SYz8a7OrorcCTsQqjzdkEfB2fHX+X5nK01xA5j9Q
20wGMX8dg9RnprwL+LfMkEWak0h+mar3mAIJBcZ1j9Q2DwkABnlpithyik9aLCOq
O9YpaxnL7OD8EKeXBY1GAdlXhUmla4NkjXEXVIXIHridYhw3vPWs1zdwX0vcwqqK
EDFmDTrQkLyJbRokMHRUOf0qW4+VqYVHQkupzvYqKK+LiQEhqSFMu8aj1nUO8dVc
w9t6W8l/l0qPojFpuRhf9KFnM2UJw8J8hSBLk8haa3wE3vxtXEXTj/kxqklcYwTH
pkj/+1IWWcsXKm29unhjnXmubPsrLq9R+qrS3GGTWkuoSCAhAQtoujBPnDMTufk2
bWD/tI/+uO4MugMw7h876BFypF8ZIn73zt2LiExfLWrEqPnwsdEltyH2grFe6CZ4
LbekJe9Ily+8ctho0meUsl7ZCaxZ3Kl774R2jNTZBoe5aXBckqqkz5IFYVGbnIIV
OxTjWFJa6PXmzbmlLuJSltjYNiSBFW6Nx6uHqAhRyRGNumRNIkynTpVNhoapxPom
+0nuQxAGGg9qZd2hfS64s0oO6aG/5OXYMYy19bAR0wyj3pPMAhJaZrK+YRIcFZ4n
EeXWcQ3pxe4Vy901JP3leyXWLGLUmr/mA1ol/A2mUSWYwbYiWZYeAW8IzaLicCWH
d7okupnZyQdst7poqZLYg4cGMYPuds0WUk7hZUUUORxvL5lGhHgj/TOi8V7Q0M2y
WE4TdbokTQOKOrXQeaALj1BQ5NXvfT51ifaPSd3YRGjLmeLfadvRwIo/FtEZqRWE
NBHD2WGMBzZFGQ88qPOvH+j7DCsXUOpIdIjUzMJnsmuBNbRvKSsOszcnXjh2mGPQ
/cfm9hfe1CUV43W7FdjqCL0Ho6dCk8ujXBSnihr3oy97DBk0XFGvyhedWCqSrRLA
xSEaZQ1dVZOIH6JAKaR2NI/hbE2D4yiiDBOhCLlg84Exk6FaS0jHlzFOMI9ngIYU
tBsWAYlgFIY61ZTdmXM8BWTl4iTa0vb+fjitKxtMPjm/MNBpQrtU+FSBUHL6DmjP
UIY1l9PAQ96zsZK8xxKi0RHqHBk/DN7ATyaeu2ReiIPDrS/524HMnUy/pn+T/UDx
rWEyn78VCE01eHBscU34xs6U1/PBQSQxOU/MBlf0u0bA3nMscj18F/kRXxQA3C16
wfDgSvvTTJifBKNUXelC+RMlK7EzhjuveqCXAP5sec1WK6s7rbfDfs6hbcos/+F/
O1E72ln54kIjGJllMWRTw756bsCBrVBSQ9WmVoClDq2v17FRIXNMd0JM6dSlEzuu
U4z1HadjBy8+5j/zjW0Uw/wvzE4RNJTA+Lne+KTuDiHexPHpw7SsK4Gs1oOZRWx1
LGn5hyDETWhFJSwtRSANghBzPNB+bxIlP050SWDy1e3YoZcNJ23ZcxARF78ba96j
kWK6L6hRZKSDqqIP0DkY4zleLL16A6G7dGBgL7I9u7OquRAqIz6nszrgH9H1FiRP
GwIJgXwIOAcXuxwnkqGHOG8cEtZdf9E5X4XOIUXunV++iTmfumeYZykMpqbOlh+b
RwHZLh9qybl72nVyIPIBWzubbySVAzPaD8O593oaQk9wSqOcFLUMRypfnd0xsmw0
azG6BhUVbRsTSyJl+mVso10t2XgT42PjcUNnHJBx19XnuRZ0KgUa8gYnHBzkCLWA
pUYl1IGSUBpTktxRtnDsWOj2XqV8+/RQgGFQ4S0U1mx2wRklKaKjHRHQqNo6MwF4
oDVA6U1HhiS3XSV2D8Z6QhO+eNUaptcORQ/cA6mh86c7ry7LusKEu50CcH3mELCl
NbN04x3Swg49wTDLtUu7+MzxaFSOUyKo2/b/gnKXlC07yb73GacRT2YJ9L429Bs8
/L5ubHUQKDELFon+ksdF+LKl2fH/tcBgXdqXlNT1EEFe5UXSTu+FQ4GplQhN324Y
1eOBy+Klai6i1aF8luWBDqQ7yqIbrGOiAVs6wPvP5hY2K2u4KJiIOzF9Gz0+wVQf
3G9vWTEnzx15fPTTQglqs9rjwoNLgc13Z9n9+ya0MELUsQDZFRMhFzp3/DZa9sVr
Aj/vbgy7L1QmELJzPBqaTQvNSH2MccyGN3vHEastxt/U83dFWdZ1jWbvBbpFUYGJ
WVrXBEimICZrLO8Qb7KAGLKyUMqpRUF32d4Tm+RhgVN8EtMUVmmlVsSFZ0TTu7hB
6mnkEME8eRG2oDzH0Ew1+pSXbnYNoAahfMSRgH2n3easK14fjJhp37xzaauz7qST
YdOWdbfBBEQdCuhpkEjwJma/2h+18ITGaVuKtnMnAT9LVAR+zja1SMsaX8s4RLR2
xMixt8zt4Z+1qNJAThfSb8/v4R2kAVGj8g5iisfMNMDzVv4qNRTsbAoHI8sG7tI1
zDnEKdgmX3tTblZsfz+DpBKZ2NmhA2Vq13zqFl4S85pZid7ib7ZaSqvP+DdXsahq
M2y027Ntq809Wjuabx6HXQI1Eq+tFskvs7Ymy7BlTTdcPiYhCWv9ZUbJsL8XYs25
ygrfy+xI8Vl0s4nRaJTP6pF9r73oyOhWHW440jvf8V5k/UUKqoGuob3ls+3Ofg5r
/TfaJ8sgU2D7VcFiRDMlluTpii618HXLT5Jnma4b080uMCV0OQwPy+9dDgG7nGgq
9EHX6+dqpZSi5Q7xBCbYqxdH0rMdUU9Jd2JRcjXDVnRjwcAB6EKsBMhg5ryfSpW+
fLl+o5HfSyNThiuWsLhnFFe2PnTWKppvRRG6d2kVWFELUm+fETBcOFrUqviYfSUp
lMWJJTi5J8RAfHk8EDqOkArhV0x/7So/eFxMpZy4kNEebxd453stWEHefBnPdi35
kNSjfryVvWQyny2SlG1cvJSsSAj7yndrt2gbMK4bfZ1aS2gXgrIXDI965bIAD0Mq
ushjP6vrwjKPwycmsu/TJEObD65/j5CcyLhu7zszqBmj6llqNo8I3oRFCxBwKCzl
raRnIqOUE5aBkD5O115YcsdksaX7orRHcNhu7yac+cBlmTBhzb9fCXdd0Edh+0aG
scOd91rdMqDAJzsAfTFeRKKgnwV2+sO73tEAQd+6dN75zQjfltQ+qnxcruolYZoG
9++zi0Lt71nPmkCb41NwJ41CptsFRkoTmb5sQ3ApHMPKtM8VWLezWPeIjbFVzVAc
BTfkeEDLpsIguz+GQDWt9uArJfEvaFcvn5l7SjXtVyW9uWzk4LSM7SaqIUvXwLB7
rjckNbpoUpO7IqAxoDEffRUzdPnVA9bwmoGPz2bj4rRfZXxMtFXcYuyJaqt/iq6x
47b6En3oiIfGmd0L2Dfu+71kIQL0y+jcsVJx6ognSfGFB6c49i21KmrfE2gopm5e
vRIvDSD90VJClkLf6y3J4jTtnjUuSzNLtMG/9C4RqQB136f4HuLVOSjtJSalgAd8
rcgFDHnhz4NeXK/cbLQ4k08r5DF8munGOmIw71H5P5/DrJOIT9ANUw5qkZuilGpz
mDm0ulEdKzY7NzJq6aOvYfIYmi1AGhN/0mG89mblBvkF4c2kCAGbVmLDcvAlzkBP
k3EDzWztwel9a4fdjtphOZOtTXaCVbDXmb3fpOQOj2hs/psAESnSbOYXzSpxHRkc
uzVlp0fe6/OKu7uB59Hn1v+nopGnVWoK5VcVBFROEzgv3HDiNdzfk8N70hAySq+C
UX00rcZ6fvajssVBiJorY8s/y0Rxxy0xZX7WEnidmHtfhaD3dPD7e4asOfOQGcjf
Pqr/SWzmiTbLgChWh3C1PdozoDWemWy8+QTRZqfd3pwodOKWV9zTFX0VVKEF6YA8
hmaT6F2ZZEt/HHRC2j72AX5o05zjc8ENvV1GSj+4YDHTj0BhamEoknD58TAZ/MMf
pA6SmpMRSdQfNhsb5SgNMVs0femg1P9DAYQ7eOzbBpYnhh0gR7p8M2w7L5haCD21
xgIQdrU+DaKmeFyns38lAheLnz25M6XESj4S4YGITfRpdjZoXNKRi2OsF8cm8f0Y
FvKHR0qJg3oDnykXpWGlrrBs3+K8kIZOR20SeVozzGgyBr0SRt7ifXhEgErhwgHb
4u1SKhKQbjVz09EPg2U5ELtDK1GrQVj42sx8XGWuMERaz2j1ex/oGkP28BgXqXmp
LVno68vFp83Lj+A9a9BUFkXM6etPKVNb75auR1YH3WXu3t8oXzg069KbL8yyF4OY
p94phX1blOyU1UerpNFdklqZUPDuxFfdYjbne9c8zz9A8KhNKyHcpyCgVC6FCTd+
CwAL+auek/HLO6SA3FdbrWVxfMtwoc9g+Yl5dIeiZjU4mj0y+APB0bZmG0AixpWl
zmu+jFnY5GmY0J7tZwTu106ShQTJ4ADqhmjFfpA0yh+ctRreMoIrDh0N2+YKriBF
a6X5BovbPteCLDbDN1FQI5f0xb7rJbWsHFbtWPEG9y8ft4EKIf8ObQPJnsIck5Zl
VedKVCAO8+BVvIOvIeDptOKny5x5OUIBskxV0TvwS8F7CbmGyaIVhUnI6p7aLU49
Yj1uhT5pDXmx9MLAkR288lhzF3AiBQzlcAqQmajquaegUG8S+ulrAOQPpSmkVAVH
+/iTqNGp8MAjJ36JdPd3jHfWX9meySaQKX2PpBrmCktlSbvC0FbAfy+mSnSbr9JV
NZ/nnUEWVWZNY7pAoxszfY7z2fqaeXj2qBnv1Z6TyqHNs6TYWaEMkF9XR8jDLeis
nnit/LEB8XEBuNT1P1nbiI/Yrykhrkm98IgbOKP/pvdBVizsafcxM9Ix1RjcRkPW
TMXP1WgJqE1xF0X1dhRGwtPBRasNhpqeB2U+oTq/6B/OcuI4+bLWvZrrtsSEbPZ6
U+Z4GxWjRsZhIWPr1xnw3W6TH/Y2D/9YhvrSecsED/CZrh7LaBRAhn3wHZBZVqsZ
rAbakAdGxQ8TcRrx8XMWPxztyNa1x+EKkbVp+ti1DH06CY66zQyH+5dEmFXO4Ncz
sC5tTnjx2OVOzmRjgJMmoUDwCavZIH+kHiNo4zRtabDkW7KYjl3YbZBHfvxs4yjP
1wHa7oz9rZGWqqZj5qL5FS1jq5YFSgl5ekartRJdqM3eSL3PRGPPaWaXQNpTBXwO
HHvKGX5qyuj0H3eQ/47AJo6p27nNHu9u0kbbP1GD+50o2u7kzKSefB7zY6wEv7Dc
h1AXcAFqrvs+43wrzJuYR8hcvzeoK8Ns8JXeAIwN2tX/ggpvDS16tfq3Y8RxRVAc
TTf8t7HfEtTd9WAmDn1XZuN3yfu/jymIukPR8dTwPIB2hTffCUFK+vYKjCyPhE0w
M9/Kai1uhvIzKQNSzkK2aFsNjy5RhEqUO6Iop5SELp4SudxfzdfwBGArJ8zCsj0k
OYypq4otW6TlKkbh6MZGbka0VhNW3ijp2Of8SWMNIx4/jcp/Z8xzgtQ0QnchfirF
uFAJouL+AOsDRn4RFMjU342LrpdxLk0k4U24fBtphufE8r6LhChPunWAaI1sImD8
Ntfs5ocQW8Xq4/Epa09iMKHvVYJZvfJmHKM+65VBBBRfAehmZzct3P3Tatht6iDS
hbOd5tarCa/U+U3eI68DSF/00JuSH6hGry7dyB+J02QfZ+wzOinDyoghiJ0oqlR4
yDT3tYcohzVKFK9DMr/DOpSy6eALMR7wOwz0h/7uoiK8Jtz73u7CKnzJqiFaZymJ
kKay5mjwENp5n5ccszx6XbAstiycbP0SOy1Urg7uc0vNh1y2KH/na1Qf65ympgPN
ZiKGdkHPUhnIdSCKsRwa+OBEwLXgxIbROx5TjOJEtf73KZmJzRYZDmyICXeVbB0p
jv/zEKUQYts8vwfpcoVi1F/r/WmC0i5bqew5N2+CZqshbhSXYWlL94ypdlJUD1gS
qYwKYc7YCWtakAozY6xGJCW/L6WpaQIJw8YjUI2a0SxuXoxRXLVKkpA+MbOx1cjO
I3Xa12cxLmETytC56kramAAgKIgjDp9yPPK7yzj6Th+wVc924G+NSKgTdX+FHoE+
vOHBs2nfeGEsIeoQg++tsukGg+M0FWc3X8okKklLTQfyFV3OtyF4ciLW/k74sAK5
t5Zlzby/mJ9+Nv7L+5dspQZukbXX5sSx1nuWDcoCD4zUgoZ3KEQDDnFSwsKlC7kw
Kc3WBsuoZ0xPnDJ+E8KuHliGHBua+gfZoYqUww94P88swS1DCm9lB8iD9Ky5Te1c
jjOdmxSOyLNhnlBK2rbaPDgYIkuZiTjrJ5K7FIvwY8HNgHqBR05q82DmhTE2Lxp7
ZE6u+l76+XHgJ2rYFYj/QsD3uHKWyaW9ySmSQOgET9Qbiq2z4ag49zy96cnEkUbV
xCProroISgAeoxDJ4hyXQn4t1l23GNeyAlpkhDs5VYTFmZxYgVxfkdyg1Xn+OnN+
/7feWBm2hI5gsQJkJnjvmng3/9QxLYNQy7ZbiL0fbXBzRLTJ1YnYlERrMAnnOuHs
LrqE8TFk9/e2+4Xf1WUdpJkPVz17sQBC/IU5ex7JY7Lb9zO+y9fh1KblWGat6N3f
TOtYjp8HhLW7MZT+XeZdesx4s3yWtJmnAwrRCXQsjuu27ccVeKuWuByoe2MTwHdW
YMEepCMTu26eMoKM2vnPTXBpZ2IuQzFaxvuzkbnh+ReWG+tHuJXnf1eYFSFEM/92
KDstniE0gA/jEHdV1YXl//GjUA3UvxTva06TburfONw41MBtWj0XnMOHdyXMVLKK
WhSvuRa7ML9KybM1AvHY01m1Mgyfie2kOYwfTjSvjGF6zNPttjjT+3EuGd/JK3iR
5GPVIDBFaQKIpBiMo60r06rejXSZjpJq5jAedKfZS3PtNYmmu/9pXJ54p9ASRwPV
ENXA067A/4jdzjTzr57l5JdyvGWrJQNZ6SDUuuis8LcAfnJmJ4F9kFURDOJ+Ghcx
ZIlMfA1sCaDB35a1AnQVf2o7YdVrmt0aU22mut0achzc/oEzGHYaKt89BHoxn2+k
HmMEs31vgt3x896TTE5D5JgcUMtJ1FIwLvEcJ6BsX6JEJ8bU1hEivpER3FL5pt5T
2RkN1lPLokaMJ1trs2pHAn1jZ9w8tDTeA+8Zh401Ba+54MYLFk3nDdLgeU5/6dtk
PWD7TUp9sKZI+BCtI2djGVnBB4vKY35JVmsiAWNFEZLv0kt9eqhruEnQ0h5iOxYd
p/psEeAKdTMQnIzc7vWJZTlDyPQlzeLNJ3n+o2gsX9123h8ng9QRlext/u3q0pOs
XVHF1cMlpjtV+XFQJ/chUCOWKxLm5xa09Mvlfxyi7keQgl177dPH+mesQt+I2yjW
T0JWvmNB+cgAKCtbowl0JffFjYyiJxvAvN7oCP7hv32hhKU3IrwSes7ufya7W9/g
3Y+cu63aZJ5S5rFAYIPkbzKeuaGpv4MJhxVV4yfUDdysyqnOQJ6CjRNudJuhrPAU
zZN7Kp3Tn1spT0pka3jxuTZDCJat1bCFLdyGlGMlovpUMoNkwSIVuSTbAqONSAcT
v2jt5h+hgV8S9n1iOGcp219GD1NG0/fB55EHz7ZmXxzccuQcnce4iT/rnmBDWZxx
yBEaViAoFPLyY/gXHnIypynU/h+Kg+73ZS1QN1SOMWgoq1snbWdSJA9t4Y39fGyG
k4cBz1sfqLwGlnuDalHBAmlK3Tf0Imk8q+H+Mqo8RWc1e/liLNjVnwPTw/VUwmVD
rMpxXP6o3VLEmWV9a00Ap4qOPHjpe9s80WVAMaVj9vImtgzSepFVzvqZBOUKN03n
DzAuuixPH87WjXVkOPCR3g==
`protect END_PROTECTED
