`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r3tE/qvJFnP7b4X4E32I2FJW60APJJzhtNFyDE1dSbfoeBnROEntWuisNfUxhqNR
0HtrdguLeuSfeIE4x+CM6N3eLx8k/6MEwV/9gDoWUmJ9TwiTtUjAQMfgpw4LKdLh
6FGv1CTRwu/dXw5Qk9AKXfJSDot4jQL6P+wtY9Wbg8M9m33Yf2IDGD+B3TetGsCb
Uf6TPusjbu3r5gsx/PAI1luDXvaW9naMohcTOo83MzPHFdT7m7DKE69xudYqUnVu
A0D3+b6TEyRM3ITwxqlcpog+JdmctYZfrJgUNGidU6x8MZl9Q1FDHC5N1BoTyslc
Mw9xtqU2rEx1ahpbzt6ddhgJ4/9WIPZt88nGe3xRaEwPgoOQRqlJCaI4Bm/9L/FF
WLFwVUS+vWnKQ09Wj/IkcsLpH1RIpxfqlsuh70SMAxhw7RbANmsgr/+mwoQb7Wd/
aU4wEle85iRudETES7AYmstcJd2uxapJgDeDDBofMP8+p/A6CLrMC5CCMeKeyHdg
dHIh/k8KZSaG4u/1khlhBNo+pwlAak30n/I9hbK4lbM=
`protect END_PROTECTED
