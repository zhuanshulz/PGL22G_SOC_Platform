`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6y7+F5Zw0xRGnXMfIW6bN79Byc2kcjzvX0knX9RZlOmyInOOnnQWKhMUzdNvBAeU
neKNuwS61hRv9454om8+pEeA9NJh+YRrjavTLXi2SXOjsBAQydopArw++EIoTcXK
V3HpIeMalREY7HNw8BXbHcsKQHQyRq/DQ1wXXf0xYK6/uSSQEpKdYfVdfx1D5icC
Y/tyFHlBvc7g70/v+FkwDg+t4M/nHa4N1WZUz3sH9hlS/v3usvZPqdLIO9GjX3UO
cuNf8yQKNiNfgV/tm7Ui3jbBBfc2XDWUpXRp+5rr/01FzTrXX9FdLhLMf7sUu23/
bwSchZWdLWeXRKg184sRJJxBtg+O9UwYeZiq6Hcu8+JPPQyDjDRDwZHIgLkz+dPF
scj/dnKotZV9VpuT/NAhKRXOLJzpJnxfMmhS12C//sKxJj5I0IZBbEf48B/NXvMC
jTlKeEB66ZjKNtaCl2EJmYLjRz53F1qeH1L81Fe+9h0KyG5eETkgLWKNlhJfB6Kc
75NznjRxN989w2hw0RK3IT5QQPDBUa4NdEBF6ygjwtMhYzShWdQ7HXJ0ZMRJxfZ1
TbTrK0V9K8GQHUCmDTKf8/UNYI5ieJcJI3aSGf9V7u002CAjNGzAzr8Rh4lgzVp+
orE6Bc/mRSEZYHuJZS/0ZB0SM0SFps5oROKklMYcThEe1ID60ZV7uCF3YcrFpfYB
CInhTq+qKVbDjuOPAABQ8EKGyAoMB9/VDPdYgVBTfZP/IC2yOEp/UEjNGXLk0HEd
WsA8SbrkRqK43XdJ8yi/LYt4tO/F+Qyv32u+GmmGNwmBnEoBrtFumn9wdSh+Gi9x
m+qiGlJifO2bOcwdthhQAD8lQEAYBTqN3AZWpnxcc6Bj6lnY3acc6a/k4WDlIAb2
Fsn//0B6vyx1CoWtCVNkrr8KrtVTvODa1fAqI0lX//uPKFsrE+3VkIoWxVabrT6x
zpRy23SCY7e731M2goGopQXW8Gpr/25OB5VNVL60WG9cTQpNdK/mjxsl3vKhInZ5
R8jzVUnSDbWaNrVdwUlU7XrsTyiOcGNqMwYyQQBV1mVXpU6+ea5qhSTWnboW624F
8AK+84ZJ7byZhiw6I1bvQrNaubGUin31hjkcckMBVrA=
`protect END_PROTECTED
