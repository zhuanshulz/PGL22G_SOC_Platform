`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GBviYyj1YMR9o4cpLDyfSWQZpNaShq75vP8errWyiciecucHEoJqMRlvlHpu7Dwl
WBqiZi7k352T9ZZC0zVE6je8Xt4/gc6ArAFEKht0x/QwTUmFTYh0qosEVu2xF9Z6
I/xBmfGuqzUUeMVbSgKVvqm5DheVCwYorSH9Piy6IWuaWfhxNZN8GniS2NOcPkHY
7u/yAS0Y80jg2PwIz8FFb62qgmEniGgv3mDC1RsGqpec0sjhsQrO/LqG/8KAF7XF
Rab/Hb2ZJQxEzd65wRU7ThyduYnPUWEfnYJR2xxMC/mBfm6SfjDYfXAqbtkbaKTD
oUqjHT9HdGIMAWSGOsAlCBG7WJadR9XWObdiHAXbDbYR/q2DBkUeEQs3G17aSEie
bgDJ0IhsmdZxHg4DWQ8tHvmFhiYdebvugOg63AXduGPAkix5JOsI+dUCABZsJhxV
hINyFn9lvPmiIxhKZJLq1HD9rm3P2d+qmDYCtzY7oTVhsTFSecbcyF/SM67SZF8Q
89ckoouxnEvg52iCjRw1ZBFHi54CBswGjc2uAaZM0R3/vxkHHa85RPE8zKGrxHfU
uRNb8dj1jFpISYhQt5l+j7ezTtj7qfJWwOaGbIBOagkF5gBuh4lTdnn4ZhiKcT8A
GHy9C7knPpFzkA5Y9yd7ymVFpG7Oxohy3l/kAtUY04UZNiAWzljGtKdpAUw/4cSk
z5lhbZhEX3MGzbWNqG9qUH8oSD377b55HgAqcC4PSTOB1xaAVl4iu/MgV+aZPa9f
NE7xSO9YtnWjm/7eY9kpO8nIQrVYqxVcTqkzdE64DQA=
`protect END_PROTECTED
