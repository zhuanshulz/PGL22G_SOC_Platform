`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gVDZGCsHWj0v7NfovN/AriOIIJSKh5eNUUr3g+Q3RfEoOLd1n0yyKyoWUcgN3qGs
ylSwsBUc5yowVxwPRmlKMq8qsnBJ4XonHUKweTlilcrvJaBkTQFbXLYwCQbTmtte
qT17lXXfzQ/kcOMmgeDY/TRegulUullU7yfyqhw+UucJPd1yMK6OKfEVvFhlbxaY
MUUsVS5XXEZy8oR45kr83kz9Vvdr7nHGEeZD3xRUYirGIv8LSSV74lKb6DLj5mqy
c19HqouBR8EG8oQu9Z7UlZauJlgAfZpb+RMKemJ2apDCni+EGeyQ/0JXNv9gdZSa
ZLTzMuZspQUQfLLoKfnJR32HXtLCe98gT5Q0s3k9S9WY5YU1a6QbC2EWWecR+6ci
YpiXZW41/+3q6yI6Ud+et6xMTTSltKvCcnyf+vOO1xrwuqIkGceix8dlj1hOsnKG
2Q7Ni8deqZopt41egq89VvSv2JVus+tlBhNjBQABAcCrk9PXyHkM1hKB5I95V/2i
tGDKR9hbu6enORWzo1rcEZvWA2XgvlyYHlwi8mQtZCo51bMKqvKzlFSTZl8guGx5
ghaf6DTxxbRCSVl7rKsXmqFclpZPoFNRb8nbgN+hj9RBx+7knJckhGJ5hJA3fCLH
BKaXuOt1miIop31hw+Ng3ivI19AlL7oX3CXigmzIGx3yDGPqNgceoa04iElDgs11
LKJ83AUsedYqYNQ8lYQ3HOYxcy5G4MD++QSsT8hsQWs+A3qvEqzKzFf/grn7efEP
n59p1EHZtUcAoFgAx80/OhyuWxDVf3pTkH8eifty3VB89fRlKwON7y4UhqWTf8Hu
WjUeK8dV6eDnqtG3K+CnwceFDk3cYacM5NevVCqfa158SzJ0EvS2iiMejlL7OHG2
dsohULoLUXvPfAWV7KF0G+/A4CgRNFBnvuPOj/AIuFLPta/jlVxmKEhRLM0G5K6d
vzzT18vuBlioJTAO5Z2oN3mn52T5tOl88BF4Kzkd2ZF68DN5sRwXUbw24kGBBpH7
TuxrjqcMMPQ2grGI7Rd1Vq87HPlOn/ly9Tx51rwvEJ3/zf+/CAWJDA4DoK4650ly
46/qxqnPtzd5uJO48YiOFo7uhlHjkSOymChR2XNIjxKeQXhqfywWR9fAs1z4yK0t
IqJmr9zmciT1ZAveypQ0tz2mpZP5HKul6HwUf7N25TdGlyL1Ofj5u917JhX0cEP1
ERaj3rwym2uiEOl9OZrSOhn/ySOUQDX97MNmMZlWG/Bz57Dqdx6UhKHAPCoTYLRx
xuSRKpu5Fh0q8g8gpltGZnvtu2yRmW9C3W/j7T4mkOhYpNKbdTRL+sVH2YQ4hqbL
`protect END_PROTECTED
