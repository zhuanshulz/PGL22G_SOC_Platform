`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qzfYDY7/0vv75agNkzADKf1Vs9yiAdNAgAyICnu2tOG5yQ1bm/V2n0wON4qlYmkI
cwBfhGpRMW8gO0Otu8422lxm2WtbnCz8O+/s614xtMjGYBnuSMWDmtTVhaQeu6Tf
LZDVlXYEqrVO9zPcnR0XaWqQvWWf6h4JrngwpGH+Yn37Tfpcy6NNMl4qdYu84a90
2elQghXFQ/On9IxFDoE5NawAMCM/xvs5vkp0iNmPLP9AA+0Sgo13o490mJnd+SER
VZNUj1/byQ6xgrKvHwAs0cSJbFhHsn/BSLy4JS239N7l4qAXBrkr7JP/WJksKgWH
qFwfIkrm9y6pbhRwVbtLg2bAlpN0GybfpHsT4H/YihcDtV1JXyOr1Sn7GXXk6t4W
XZ4yzi/B/70tcR+UJB5Nao+Zy0CvlwukKupR5ByL1BATHAr9dr+42bxyvgs6bY8T
zIku3Q1rvBN3RF8kQazvTHOy2j1DYWz2pm2toiWUreTcBDAaFWSqG7PfXWFvbcBr
pqBc0gspVJsz9EeYxxlNRpJSqFUex72x9y1Ais6zUxCOPYkJP2WUjabZr4Ccv7Kq
7uZZ7zj1VuThklDdb6mhAvqm/rv/9foTi7/SoGDl4qqxxfClGamz0V1QoOlBaNgC
MKHnuolmi8715DR5SWW+sC03N5t4OLtmZhWmtBg7gb2wpr6MfHLY2ucYWNVwZnQt
q7Bu4o5HNKCDhW0wkri7p7O1RkU4MY4M5lL7ZPiMRcXFteizlJ5T49Qft29+0heb
2g22icP/U7TRk4E0Mfc0UNudoiSYiE9+HJKN49X5jc2UjFf34K6EeHhsPvEE7swg
OSZO7wHYBagtn73hKOg4Jo2TWNu0hEiSIM4DEMVzVBB3vwBxlIrsP72yV2C2j2tJ
+UpO0sSl5amAaEnLeRMptxGB57dz6LqWggcMq5dgsX28uzpDVm/TVfjcSJNuNnZF
hmfj9jI7sgmut03GkTovD0FTuwekEcSZjSE23gupOQAUUrquzDIqtZapt2NrtNFd
VEmoeaDCNS2bSGk0CWt7HvIl7TtxQ1Utll8AmS96yfh/mXG8NCrlRCgX0lDqMhLS
2SLSBjvIDg/oKpSTO8Tl+s5wJzN8ObLjQqPtbPx7AWUFnf80U6Jy4STTEF3Oo6mW
7cQDkJUFEeiEyNs1XkDBdYr785JTcurw2Rl1FviX6GzNvDJ5+RFvf8+qjAesbLyV
ZsPflbmj5JdtJES8Nc3joLuCyk3Tw4tiGvs8oPda2NxvU+zrXwX+zwXsSFZRqonG
4c/w6MpcFfHpdV4tMkZrUzIe4LPEVcnc+MhdM9xXnGImxYj0Gb0D7BBlHpnNVigH
qME4wjRbi6EiZ6Dnmfxjf/dWb/0lM4IWb7LJb3RS5vkd0f7i287eTUvYlPhQLy8P
b7n31TD4IsYiJ0Diacm/dUPEfhw/n9WDeTzgWXDgt1Ze+Or1xRpCQa2eyjJQ9uUF
/m1wyyJmFw5UDtS7tadmNHKkPYNbyM6OwvAut7UPE4cJadrkrIKe2SU2iE2chRmc
kINLuzF3ClkxVfKm0/BFmHHthZ9U+cB/Twj1WGE/3EUQB5HsSYCCMcSi4kI+JdPh
fzGVsYekE9YucPddo9CI0l7djkcOVp/y+Pj2pZiRz3zOazI2AeOD6xsbszu3DtFY
8Q3yxQCbhioWOdDsZmaZloUSn0lnWWFDSYv5uaX3ptg0+aceioOpsmNieuN70QLE
RRkS1Flm8FNbIee54MC9tMId+bPmfZc4L1J7swPwo2jWSpd9+AmxRZoIl4eejddo
nEAgCMOU9EkraZ4nw+oIxrGs1uKvpElmLVkXuIQ7IOvK5PbsmFapsFBNr3M00OxS
AIIZ3H5s9UI2w/wS7VecmUVAXmklb1TpRjZx98iPI2nzO9fXF+50TkviGqxY9a20
4DuoMYRds6/MaAKZWKAiYGPhyfd63BKmRC8NNAjid6dyK+gJb3uQUPQSG8rClEuj
qz5yu3jyX6TH8L4lFPR1t6BVhOgmaZjbP6b1t4BFFWAcUflUveIm9pOyT10UcXxr
6fRb0GLmsExToRtJhte7j7zU5m1NryhPE7HqrB1izOgpGxZpBBGqP4dgL95tHqud
1MlQt/wL5bmntUrkqUwHalq8MA/hlkH4ycuT9Bq54L8S+Fjd+59j3xhoq6spC0P/
HIpdnpjWyDWZ+BGo7Xi36FHK8v9Zi2J5LZQBMNj0q9gOGzSjVQ+iJAcrqKCySaOm
GPgGZqIB9EBzqtQMU7BQz6j4MQ0BN5qtarhE+LVimfy09P9bRxjpALwV/pV9lz5U
dMq2gAijQk3qnKwTm4gYbchE2T/Nc5Ov/yBU6iMKcNOn1dLh3ETkBApkC0d28wEz
dGkQD1Tu0dNe9xZHeF+g/5Jr0cSu1P+gsfxny2DpwztJm+etHlJdrAYRLY/rphYv
DI1CnghKynu9Q73tvlrPmvQJeEwQ3dSiOe1FJayOLHlWXSlZPZVhpGc00xHx6KF1
2jEiookpo2O1Pz601la82/Y8sYOw6zq0DhB2VpOfZWuLhzuW3ALeTWY7Hnt5gjSF
eZmqoWLI/GHnKGzFNKC8OBVgT/NyZvZdNufwEFwopVmvqNdO3KoMcRoApLtJkb3d
z51AZwWWV9POD0pBW3aO+eP2DEn/2ugA4q5M/piynx1YLcNE3lfHzau/nxh8JM5R
X8NebIAk5wcNZC6Ue2x4pN7yaH4WAXejG8wB6mH9/OU=
`protect END_PROTECTED
