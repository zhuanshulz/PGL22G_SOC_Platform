`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zAEpezGLyubFdEnTIvx7uXP079/vtE7qe4qBori1a9XNxZmK8Ir2nTGr6RnFTZvJ
DsUOCetmk+VYvzVvTNUE6gDHLAnjr+MwWiFQQr9oCVEAIn4Cpc1wynLIPiHd74Vj
XdQ38DsySHTxW4AS7GABGWVyxaPPIT6gGJE+CKnyHtBBbZX+bwx+94TNgcTDQzvC
2DLsNHu7TmcGSIIj98+xLKl/sm16kEfU0i8sfVmRWe2WlO8d6kWrfFJaBqGv6j0d
tGcc9GBnihE/3z5ZDP+fgguungjrZRm7aNRDm9InLrO4Hw6bmscbb6u3dEuc+Hdo
h9KvMN6Kux35I5m0dj5ZgSrSttUt6KIMwfKTw6INVsWK23d2paKuNd3ASZKjnl6q
d+D0PJFssjW2w8df4wCrKTnRFZoxYO4xr6bu5z3irgFWSHR9+2qiT5cxt0RgP/lm
TOs04BBUvSS4OxG8eoBjnkPFG02fENNTmoOueCDiQyvEvZdzeL10WILZXUPz78T7
LxyYL55XLs2259aoefiOjjbHHydSby32x0OFg5tGJTFu3f+UplEQL8HGIaBiMc3t
TH4MUmVvZkBGL5bm/SHnII0faBy4Ydur+slTzioOTptcICw4SvEYxCrw2Qt3lXsy
T/CFx92uKPPoxeFd/TpO/oCn0lLhkUxKN/plKgCVjpaadBFCup+M55lY40n0VtKl
D2iWVY3fDKaeFW42GzOq4Eu/XyjxPLCltVP8LQhnIf7+heBtvVW1b/PAJzaQbnhe
EO/lmLC91a9Kmbz5VS4+NBulDWK1ahPDC/d+f/7Rp6eX62PukRyDPgXMYHZkR2x1
bGyxe2F+OpMVltxn8UuVdn8gvODKpRDa5+o43pPoBwiq4Nb665MI5Byvc9swGt/s
CHN5Fvlb69P65r8+btd6yWaHcgr/5SE6fACOsP86sdYO3JAyJgF0peyUfPbZ03MY
Zm2CBCzhKMVvBPwpNGbavQZEMREzrtL07TAxmRGioDgmLCwd0jzy5qxEe2FaNqrE
IzM3pRwlABEOU3rrbjnNoVhxP8ohkLhQjJvtlG2dFU7bJgFH3EfEuD1P/C+sZkv4
Pf7FqzQkQJcQl5zn7kZOekL4B7B2roOhpR7iofw0jBDsIydTxrUWG9dNKy4WLOE7
l9EkUMYCL/dtux3dXGAkjctiqrnK3M1iQtcDEq4YQUxDAAZD+NuKUbgqkfUfWC8W
0cL2NPwC/2zIoJvKOLOkQ6NYyFhNRKSVoMxdaJs2k/wCxTDtQHkzIss83cjNimVp
Fz30pyaM+yCiAeabplXiKI08Qcal9XgAzXm6yrdPwBvTNuzdSa0+9u2pfLe1dKlp
pv5VN+iHwd5+x9HTuSLCGk5bLJ1rb62/kR9lNObiQHJSgvO6VVvAbKEBv/pQVW+1
X51PSaY7FX3LtC+pztOAmgLbW512WVeeA5xMxDOfLSdNNQWUmKx6Me0pC0CqO1tx
5tBs7+29Wm+d7a9yaGfeGFKTiRFA7k1f1IKoRCIiVjQ=
`protect END_PROTECTED
