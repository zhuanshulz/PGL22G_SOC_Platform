`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s1WKPSLEghC6vGb5ISaSWLw0cCyWJ5ZxSnxCJmi6VBvlF4Ie2LnWSkVRp9eflCDJ
cvZkJtd4Sxtlu3+2K8lxID5n58NM+QHahRIBhRPnO//YvcdOfgVxr9fgGrYGayo9
V7kAbjxEIwPYOyjhkghFilo8Qu2Jie7deDrsVH2hIdJckskdmwlfGMP+N5TStYT9
4arh6xJVYRGUJBCUD/Hy/TPmiMzNL/CgKeFUO99d87LJgc5rkVTzK2vODTvwuhMn
g1CwCFEAVJWJry70MBtT0dqnCnj7j21gXvvPtvO+Bs+PkhN4HZ5drCc2LilREPvf
9Nf/ca5W+voHHvP9eGrqV8f8XleBOB5N2Ygf3YH9W7KMegrC0PqocHdKJYm8v/bU
ZeOmmMJiRZrjWbtlrY75wb8wl+VArl8LQbBOMPs7Mmu7R0M23YMJM42VHmtMjyQf
u6PHSk7fE2zkxwP3VXTk0Cti7QiBGoeYTZmahBY1DdOq3gj5s81/koXwg20Q0D5J
ZrBeAha4OTQqNOp4DnmfU09bQSIgRSuWd8MP8sVd8NYv65UtuHxdVEdCGSMsyc+R
IY6PktwVLbS9skJFiV17hse4mEhK9TtIzf0qPZ7DBt3TDdL2j2PZZ9deRVPY+rz7
`protect END_PROTECTED
