`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SUbaV9oDt/h5LsZ80Y/+4tIpPWjvTItsSl921vH5+nul7n36wnpf/TCf2BfdHfmQ
NaZttkmrjw9N0m5jPyZAsJzTyot7vKtcgIZ02iQHfZPOaDZPDhxFoXAyjNA30kxU
MjFSTgAkxNdVOGn8/Bu0qO3kK14LpzimZEcQxE0/IYwlpZfb1YHkK+T/qubUEhGU
KzELKcGcUER6mE9eaTH32f3AZVz+0UPtD+19NADEnurLvftCNFJbpo2065iyeSkO
FkbSWTQkfSq2aPoO/R4m41BpN1xtTE7BSRLoNn9MnzvD39ZTaKwfC/EPWZX9iwTE
s3HNYeQr3JPHV+3idKmb0qh0rC5Sw5Xl9V1lMr6trQTsGSchrqfQwe7a1JwimZCE
SpRe+HupR9wJMr4z3Ei/oMIdNdzCIlRHuiXx3iU+zzQ6i0eEqIUtAe9gMa8lHRIh
cGAPsje3K2VIrFbiZChJXxZ2FGxCsBlLq8KAastVeIAXJkFrw03fThHKK93GNkOn
AMOqJhCW3DFGuzA3Lap2yOjsn1Dop4KyFNqB/8zFhsSwtC/6qEmNfM0U9int9TL4
4uwr6DXBnERyx4+jtLKTCXTqSxEourfKLX+4mpnABsBPPedpwPpPKKpgMCwc1DEg
2/Q7Bj7ZAbBzNIbGRUVHqRZWc2gJV85PloQQA+EIhre2ynEM6DJodfd+9AV8PgEu
0JCNGviH7wSlDFnloLNhPcioWYYgbE5I/krdVmUu+bPWEWUBBlAX4jR55yHOOKHz
Cg7YB2a0IM2WLaXgp3pbq1ct7Af2e9jVBPhVmBGdbWDsd1Oi6Uy4rSgG25W8tHoX
loThq1C3l9Lp/2j18zq3SWpZXzplHQehGJADe5apdErwiYm/DcgD9VmYn6Ekv0wn
48LfV8zoMGbuMfTGGlE8oKuDHW/oDaV8U5TSlZ1p9aYps7VPobdg+DMmt1eAtopj
RSyKCY9v0TMFebHk6HUzAk9hdCRpWTXIpMlnzYgN9Wv/+Zhr3ZQjvAzXlM+Jy9be
F/MGYbkpr4f/ZGD12YRy8xOD7IioEjYECtx6BOYEY2r15Xf10vnpNrJsvvzTLi9T
6JPE9vziWggGGIhZMi+vY233Dr1BkIj4l6l42bTKginP/zbDTS0DJagze7SvGg/p
hn6Mo8XUNev+uFKmyzOzHoe7fElLEM6lw8hASN2/PMXZoKy/xH0Cse7+2aNt1isr
AZjAoYJhEk9K9VPbYpBRO2GWEw6TLX1mzAEagnC4MlvagpFJeG74MBzRoqWuju7S
AZr2ncdV3YZv/iCUkWj/tOSLZZaI53MK7C+p17MwjxIXEQ7rEYPMKTo5+t846q2X
jfPGLZoIey0KFxNF608kWpKe4fgXVpYEWL8iENz9KDW2y2q8Q8ZklQdMgz7yfjEN
vmQ8cwQlg+jLzuuBXqrG9y1PdcxfuXRiMVtO8bQiZ1R/jnPz91ikR5/Jy/X9Eq20
WhkVB/FXcsMLfKAfFOQ6E/2nStvp6oN71/7tN+6SO3gq9TqpXRghW3ml/fF3rsNo
o4S9T2zYkij8850/zpHXCC9QEsVbbsOV6Y/WReL98Wo6CT2xKazJLHzCAgCSePdZ
b2zZjuNYLTwsbU4DhSx73W+Euga3qLHe8R+TIr89h9d26z0CQOWm+P3x/46Wrnch
EyRaFuPb+aWaHKMOQykcTTp7Kw2b4xF8gXvp/8bCrt2v6UVhlykAri2WwuwbqgpB
a8z+ME5TjEH6WsoSPZyrYEC8o3abT2vNBGYpHY+QNQmjfmCTSbu5pp8rlmcqqW4U
RH/l4ruswy7KAB0UGTUX/S6OfKwiQqd6jGxqYjZc/VcZzWxzQjz9/ej+OfzcBuBZ
Zrcp4NO11zPoCVTr2wYS28ohKZUC8FJoKPqbpeVFHT1/TggFaLeRCqfWV2KwV579
b0hjxmrz81AI0RIu5TMbRCOwqfSP5rokam8Td5OokrVVkMyOzWqhlmJCpjCIAlfP
XFQ9JYle3KQMi1KY0Ka+zi5BTuXP8RVJA0+XbBQNu/jNICxKs8q6mRa2Wc3kAg0t
ZQysOzjNDXkra0vbQZAZUmesuM8xL3CmhHMz7Qjs28j+Auz8e5OgmBwIEPrdThtB
jWiZozWLOW0i1iT9oCfe4CFhLeqk8iIHwqL9fm4yzPeDavxCrMP4+l8rXctEZ6Gs
rTEsXwOSNeg+HaTNZmPafxiZe+AAKL2rLoJtoI5YLo0Up5rk2iWGxukwu7VDW9jF
kk+53dBvQWQpYkr9GxYN046S4qq4+NxHxc3SH0WBZLkI+5tIFjyzYhO3RurE6Czv
2Z3gqmfoJ6n1f+DN5s+WmV8p4yOJV8GcZwKbbusF4P2RqZs9rfq8u7bqg7u8dA16
Ua0g3tsIiCgifudfsKOxL+hFn6KkZHb6SdWsu0zH5+BSA/N4GJ3vHD3vH+49TDYM
5gFCuv16mfGsmpCSkWxGgH03y+gB60i9bdOHvGlY0O7rZk7flopbnmtHy1RvDk+n
9Z7+bs49U9VxQgYSh1bqO1Gq9pHVEERayIda4Bej+oRd8FdlyrD13Wz5kHnmVj9v
wXyjfS2RJzI9scHtZqyKp48GYx+eRsziczc9EXUejHkXjS6VroD+FVmKY2V3jmi4
xWFMB1P8sTHpFRiK0Tlihkm5RqQEd2yc8Nzh0oraIvoRc7iBoodsAJieZtUE3Idv
nqd1sR8+wQgFcpjev1OO2shZnUPjBDwaXzp8YKoMedpyPkWO1JLKYALPHIQgHClv
RHtrW6DK8ZOlpKgBvcKW09puJA2imYDoL9g7QjcuDtOJ4NHaLab7VshBuE6V+cLf
KnApHadRnUzKk3FrEsdLwONULyrjN712j4pPqmbHhdvhf2p3H7C8n/O5ypPPNV1Z
hVnbH7JxucPQfzfwks8TtwphdYC1gIhbH+crpWkjPb1ewDGdxYshQeQJEceeT2B0
g8CV4jrMdwFUYOAumX/kND3d2P/bZKEZ8C2V8pykBGb/XXys3nXifLPsNa11i3iN
+J7TJ3WJO6WH7GwxUHQpAgiRxDCK8jms4iCSyjLS0PgeXJ2F3PvG+dHn326hAbBx
20CNYkguFV7BlCVpzcA5rW30wA0pgw5MnGDncT4FHuqyuuFlk0XLrCfElknIESVo
nevinmfIUed4EETzTizFCkvrsxtPpP/CDC4CISr8uZjJZ55RieAlKIwXC2Imtjkd
EmwRy7fM9H9PZnMkNvdLU43AI00JsHd0I679O3CCc5jXG+CQ4aIRef6WVs3NOzUh
iTufTwQlHftIc0RLW9i8aPUGBkTcaGnFaQGZhF+DEVoGiBicZx0pIWwXgnrUSgaG
n3KVTYdCNzHXq6MkWS28/a0XY0jWKYgeSLBwSWaUvv/laXHCPV6R2EZf8ClokteJ
Yu6RY9V9cuegXZ0AoTkH+1ralJn+LNrqmD2EuS0KrEPqmYif2oNNSDsYdszNBHOL
1YZPwBKUMVgjPVwSnGs5Ti8IP1YjV2xAXLaqWsIfUnY8wRGol4KGo5QlyqQGoh2i
fZkA0d7TjkdQ2QyBt5aZqg/X+xJRURib+2eRwRANX0/PXXyfewAHHpEi+QIxVspN
AtRklQcZeG+FU6iLguVY+eKrApB3l5kyTodj9XfkfyyXFYlIm5ypQCtrjKlUlSEF
n+tqKLD6p7sKsqVOHBb4odi8JxEUOjnWaKUCnDMxHw/OwPk1HlxiJ+sMku3sRcTc
r8cG14PpEqFlJXOyhKgy3BIYXXh787LzvwLxJKVY/I7ZVfEj8Lqi1b6A7Sx0ly2i
0GV9ev2iDUpfRgxs43j7/6ZyXap6ghT3qDH7s/7bJp8T5RNWTKMcXfNHXvgUSENn
2eh1lltFp1FkalFzrKfnvRFmdoowNCc4ROvOYR/9xDqhTRPsEu97Vlm1L0E6f6Ml
N/wB0W03Ipr7ixMvcP51tvVBCfEWlOpeM8PGXZaWwgXorAj04V2hW563qXBzX/wZ
bs+KH5e4Tw05r+J5wG9aCbrw9ktxR3Qpg5yPSgOb6IIX29SdSmyPII4CElCHUj6F
ZgM+DDVKepcb/+MIhtrR0AQbfoLrsI8QPBdzPhXTR6Ru7v8+Fvi3L3ykAGKwMEUY
fyfDcU5yJi2uCbZEMKAA4+LeHDKeMl7filV9L+yxzUxkJPdaDF/avMPHTQIRTbZY
Aus6uuA4ScCU1Bye+vPe3sviGJYdDmsGbKs0q2P7NZmwlgmKm3DTu3zCtEa1YrXd
JqyY1Wv5ExMwFOignFWn+ne+rAymoOYxFPxi0lRkjx7l5P8gKPz8XRnMWlPNEe3g
p3y7PhgYjvnrzofv+r8EoYJ439/OBjuims6eHkprfUkdlWJM14/6+N2/lrcs1XaN
HWngvPKwDjqWJ/GoD+g135zqxaXcjXM5BjmsEGIxPuE62Upof8chuFk7xg/I6cbF
us9Afz0KqjWjWucfV//NuUkQXlZRev8bEmbvBg6/Rl+K2UKERf+SG8xDa66KllpT
XTbMvD0cEiqyNOyXfsjebsKHLy3CZ7lFmbx4IeBwa6hURiw5B8rkocWaF9qgNYsL
ScqzULUvuOU2uwZ8+W6yX5PgcU1A+H3xcxSwwyxU9gtExp0s//fUeh7FDfOLwKA3
2Dbk/6evud8yM27Ue1cxcA==
`protect END_PROTECTED
