`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jF4tptWnPS6oRqfjahmUjH5nqsIWZl+UA2izm2WrpBsMhSM7dGufIJ1OtCaw+2Yz
o6xCi8f899Kiwio1qCa2BjOBAL+PDBz5ClG1QoqpNKXCv7eUOLc7AtBqHKuJ70SM
g7ZnpGsVd4cYcLNWSi2rN1zJDl/gAhUYtiYiPTYOyhMJmBgIbr1J+m3zvJB8Y1P1
QG1vb93J0Ps9Koe5Bvu7ld5P35Gmvfo9+zotmo7DMj0LLlSp1yHmAvY3yipy2DEv
5SH1Adi5uKIgaM9apOB7hihHyZ03Pd4pi5MRtODV96EK2ZN5iBpYWOjMHgkTgeZS
7hxxLyMWv/VgARU3g29Yo8nfatkTvf3zWvDqWFLAnEkzK6RF8qSmoCA55N64trfR
nIvVybQtbiQaHXJ90apeI6oNw0Itb6VDfyOecA75BE1RNsxV6mUKcpVR0GAhTJL/
`protect END_PROTECTED
