`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n/Cv188pmNXzzhyAIgtGEuVtu4LC/l++jSeJ8BF6rRvIgHFlZt2KkZr/0MkvcI7p
ZOJAnmqQZYeEa77WMIE9+UG9PVRPpH94Schiu8fMwD50FPgA+fxmGfpT2b0djeEv
ZI1lV0U/jvW1vnRNVjK54nSSqcvMIY27g77T1RMt59BjYqaLSJpOLS1UI20Sgdnv
BIbQiQ/XGxC4XdJrJvyLEQWdVm2ZbgI+E2GzuoGu3RVmI5Cv9RIQCzoa9Fjt6F/1
8qFa+H+Xu0sIUwfyZN/o4kR38WxPrhzTZMC/FNBgE/q2LGUKbbjD4cSGyF3ykiwY
TifI/nfXNIQCupZhvYTY6dZD0BNFKmaKeVxsoGZ7bTNnr/mZ8lcrfL8KVJoA4Ooh
hkn5D29H+63i3sCc0ICvZXwocm+bt058Yz8z1C1Sc2d1xY0RF/c7qXJ0a+ZKp4lQ
sKMQpeew/ABatNFxp5WRkrFR5+DKF/oMEc+APywPGWmfGtA58/mWI0xsvNDj1f9d
65es8csdgs2wx+glLrBOrG9+yQQC7fhb7YWI8ivJTmc/A9ssjIGvHvaUO45EXBA3
6AM4GOkMEKuml8iVDTUAjPP3uN8HFtUqHfjvhQhND3WbpFcudyaxec0XDAimwLvG
8RlBCue1dfznrqlGDpwNkyKAvS8s6LMUl4OBwimRm/sVWNGJERU6qoi3edLFJ99U
tGZQYO7tZuvj0qB4n7Et8hn1kyy2lGUaat+S9So8Qn7rFJ0qXNn3IojY9vAX2ROv
Yq3CATaXT8oCkJyZz4RM5mdxRsBTAtBTPzFiQatRkR7435hMyVbHZYON506bVBeJ
r1IMzw6owGs51bdcPa9OmIY8I+rgeliwiE9blHKfRjyrGtmjZxW0dLbNxKUxx/GJ
aJ+V5B7dp2iRGiaYi1caBO8WLtMFCjr7xoYqv0fS/39oCST3lJKt6dPXSEaObeGb
459sp48sY1IE3W5vj3ON93758LOEtMOKrl0wbFwg9UdcYbkVgZqnjOiInAZ1vqIr
15dfmnskvMVipleCrKQgiLYCuNJVGj4nA2hLHjQUQMhIr+m4ntIzDHb/SMFCehRW
XJvVGy0PqyerrzdP/LJgAtmT3hTbj9mTPQV/tXqQ5AMl0Yp73Xa7wrxlhhzX6INg
wAALgylcNrWB3P3ncRxk+pRAykwbsFczzJFuU/na8LU6PazAwERmaWwhJVRlYKpf
S+GSileSE9r4Dk6AC0pVu1/8iiN8CaFUTg6Fy2aEm2tycaHLSO9r/I+D2zQukldD
Q78zjM3dVHLi77oxXSKS+hWGhqd5pxKLJmKVZ2AhQF6RmkIEcCp/hyQacacTwsFD
zMNI9JCsL3iJ7YHjz4vlLWKHIOYHF5kwmuYdLY0XfM9QhbJHNcM4A/QsyXQXUZWm
WN1bXHu37MwGpgYYV9R327B8IcmRpAgYJm4Y/8q8BCepH/SML3g6OcJyvfce6God
h4WLZmpfitc2q/oS51iqrcVaVZMhuJRW7R+WCvUe8p+7GmC5fJyMn6sjlap4oezo
iJ64n4/R8tKCz/TubfhVb7S+XIejYiueR4umQBawPHrJnGGAVMQUxV77pEdKBekB
CQgLIdsrq1gQ+KcoVQNt3ygo3xOEuw4WlG+793QbtmjLBVxnoxXyeI81f9vfG6gs
EvwbyjhgEgewcICAr4K2Z4hBsYPZRSrLttSwUWrsMglLl180Jxk+MvMR5An/2RoX
nHoN93/5O0+3FODNYSIR6vGQ043K/83r6y34O3wh1nY780QJWzlx9VqbovzUXKCe
pH8ryYCdLhsgWRLXsIcNoREZ4NZN+HLI2kRULx18kqqtMVEDg1W6tzKhca6Rmt0l
gKGg1XcohZz7Ff8uiYgI7+4uSQv29JNrXGOppR7WsfmLVB0vc3qIealdUrGZ+fh5
PXp97JXLILt6vr/u92wUPo4+d0a4Dq+R/wRRcfIeMU8+c4Ff2IiP3Cu67bUIxwXn
V5Z9nFrtKgvBVKPYLMBmYI6n3Ey385fXCLTqV/wO4U9QER0XfdWGCgfklmptePsb
dSLfNgzsf3pEa7ph4FfuQI9W1Rm+q8s4qh9o1J2I+MEUbJ6p9jY7opu2aEC3m1+3
vgBx6g04gsacoRzr0aIHlvHaAtGBeeiJUGRf9kSJxPonRQCYXAnb9IGmN5sIQ859
Wo4CQKXLS6SXS3kvhWd0jr3je+f2GbnZlA2RTfIQYmgstQzhbg/G5wsprBqzzsOD
XdUeSu1sV8sdxq7Gi39YVPRh/IAzF1y4K6SI4x0Dz63bg7YbcuGpBlsY4/uLIvLz
7ScuKlWKJNgOoVurc3fxFUvMlwhahc7r/b5xL4K4YgNpeox+OH4h63H6rTKV6zfB
QGpB8YwYuukB9j0VqNRHWAXh8XKltQXsh/Z09rxZVDJjR2mn1dE/JrWgmN+55JMT
ny3zPBHH99u4rz4avoEB6FoKL7QnDAgWccupUKiLJkfSO4EpTQC6aZ1ZP5Et8r74
zIs4x9MSs0qnMuwE+kxI2HpvEgw1JFQ7OexnHB7z+rlxlqQDBKJzrnD1sdMAdjHq
sQb+c6YJw1gmKkMxhG4ywSrX2am1+ZLp/+5UwJkLtu1tuyqY6kirxt7mwxbSz8za
wFOrU96bsEmA6NMqAbM12hfXUkaXHDLq+r6rUc2s4nSrsctVSCCim3g3CHuksO0u
8QIeiRjk3MhS5zZnJ2CJjjtiqoIfgA7iIGf9hycuGbPidwzquECr37CG4PwCKSwi
Z2qacXMspTLxg4QiioGBe9zGr0T3ZkGQE2OyOqcPN97MYGl8tfGfLWyu0eqthEKf
Fnpltuwn0T13zO+1GSmsKRPin5rhgUlVkM6mvQJIn/K6lOhsFEe1aQj9wYfPUPVK
02cwxSClKPOeCfTis8oPq3ex43lUknv4B54aV1cXSo5nuPvjzY0izRMmAxjs82Zs
/XH5oDDpRebKuqF8Cum1MknLag0lLPy82uMHjUJ1zBUr9Ixcr4mE9302OoIKA3tW
rwyuxZ/D4KTjhywTymH+qA==
`protect END_PROTECTED
