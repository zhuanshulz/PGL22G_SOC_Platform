`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L6OZEAnUu8mFZt05FIf6mljhuwiJ9b7uuxzkuCxcrEVuftj8OkyUfI/gWcuujcFF
l2rgEOGyiIBm2e2j4h5x9vORwSfGJ51FBxMmCK+sFYW+4hk9Gwhtf5DbVpBA6i4w
iyiTYWfRfkt7BZpbTSFMN+YQ0RR3uJgYy2bAMtrc7EI5q/s+88kNKlcplwbVQ3/R
1NHCYrKYQLjtjkFWSRs5dBQL7q3f95R02OfUx0RI6R+7r/Ny74Asu4+W4hFv502W
NHmiIkwn1AWWhB6dOHCRqDbWmeX2HstWQci4W8C2ofjvh5WlPDJL7Rb1xn4++LYs
/Kfc3p6koX5RfCANNSdSSrKubisRGkINFWw0gcr/+Y+IRWBAfQ+fuXi07dvAOU6t
/s+LXoJn4Vx7qTOef2ibsQ==
`protect END_PROTECTED
