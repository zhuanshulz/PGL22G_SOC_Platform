`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cjuvYkaGBKMfD40/+9ehcK2rgDjZdgYbCLSgXzMIMQ/C73kkr6CUaQV0wDNrwTuX
9WjA9vblChyqpJCEe7rVnY7VWZ6kOOsbqYrcIhw1aoa30X0n7itBXCl4tXWRjyM6
Irc3ghXUBh60nla5g/E0wqJMuph/ZD+WrOsXwE89HOYzmm07mcT8eRGR4Dty860Q
FK+Y73xUvqxIDJc+G0cNsJ+FZr9cIwF5fJFrJNNnWy5OoxLlB/lX27o/cilvQtQY
pzc4vxcPQzYt+N9lFnkPdIRvuBPvnYNuuJCNhCoJHv1ph//0+SKDs+xr3rZ9PSxH
dQIcnwma3VDykLdnuxCYJvE7NniKeULxBhXnJN6ONh4g8y9tN9N+juXkrR6JlXUk
7k8Mq/7hjE5Oi0mkmDpBiMY7FTpupqES+LdsltgqOEO/bR0bWfygg6x6XP2wFmPe
rec044Hz1+DST4ehPmj93/6T9zIT2xWGPzvZxXRIZY1G0fH47DYmP1GPALNq45Av
OLltBAr0CCbGeGz4hK4e9TJ5lHO2T/yDJ0n+u/VNsYvcJy5Q/8j9Q+BrDPNNv59f
o3Dp6AFgIhxx4AxoF2XUf8bhvJe4S8efiiVBCv/JagNS/eT8gk4N8zCChOl7HgrY
1ucNbsnB+X5eeniDbLt+uCeqeMkYai4AV/112+Xc3PWNY/j6VBuJJEogdn43zrog
+f2WsI/XZ02O3fl7h2MHUgbo3zCFZw/qoRy8OH/jWMQDswrjAISy/yl+EbKHxvf4
PtLg4PVaUe0LKMz8awJpNboqxHAp3QGh5M0uaCI4WBRAPCAKjfEy6XauiWWOQMaQ
o18t2bgPtFiIu+yzbU95vIX6QbKxEEh1uH0JKZOmwG3r05XrMK18nRH/obHm1RYP
ITnZXKUFr12j5YKGaHGaVmOmpE0Xok9Xv9DX0ticXwiUyReg8Mwvyjmb92PL1Jo6
JA8zfBl2vGyFBvdhvbATzyLol5s4zgpk11x/WfiOvPPPmR3OyyPqhImumbKje/CK
tbxWI1bm9qarAh60B6if0aWcx3Lsj4XBMDj7nbH9tDiDlGIx1AT6OGnETs4r5idB
/fiFphFTtrhNAX1kT/7Azi2mkgUkB+QhtUaimqtWdAdgOFm1H502jlYKXrBEwGqE
la0ZWTGkhsh2bGQqZG91TBX6i0llQ4nfHvOU05woKY+gUgovhmT9JrTbSiy8kTzO
Pgy0HzTy660NbWC43kzXCLMsncc0ObvClZ6C5cGSGIUTfmxTcd7K2SbnrctKUyeR
TrJjAv5XeAFvue8lFTX+k7PTwYdHR+8X35Nol60hPtjoPddo9zArnsY++sEUPkL2
pJ3w9hHpIk74Wv4F2OgOTQ7cTuGa/OodbakEnnJl6+OTcG6w8N0OZwXf8FDAkxeH
CmkXrN+k9vZXwq/07/rjbKeawuCVcF4Wh4axKhN1NiyluYM3+kcLVA0vC+qUG4HK
qO6UMDVwttdrMhMzqWG73TYUNY/RzhPysC9cVBLu+QyzebB0QtKxpNo/H2/kru/9
thAtcpyYX66ZTIVld21aVHsARhtwafK+BD+u6H+qOuKC9OJdEpA2E1IoS1yAopHX
mG6nt/o9Vydydymw2FlaHn32IbnjraXJvZl4EiMFr/y3UbRXxNcT7TSCu5IB6gcl
omjvGsYwYHpOKu/1i8F8vAY1RgXyvCayUVKBzDSxTS5Ltocg6b/dmOrWljCSjwr8
tfzvFV7SVECBqq2hG1N+2EbdpqDXNkloJAhspIG8LJ8CS8ktzxR6gBHv2lZhc93N
x1OJkYMUeutMrpRgvC4chRpQEU5QbAJ/TzeUQMSU37uxRvG9PE/uH9c+LCaYi+VI
f4bGa5MoJ3JM+GJz1McRPp8uxUi/4C2lAjdljcNlpytxQZU6uvi3vW3/6vuvzXrT
9SSHS4ohkWLqrkn0LlONcNLTmzjqhuyC8zGwB2Teu7fAjGzm6c6qaUiY6RwC2Mb3
9eD/8uEkxKQ4qfIklGUrrLx6o/VEf7RPltk7y3BAKVCZ7PIVZaxSDS4Z5mcxntWa
xNTgz61tuZA4Uuf8358d+H3BuhnEcmS+D1YGUm/etjpHpwxwVoSy0gVcYmdYcXSr
bDR1AuE4NNFOM+vUbjtkOPfTcQBpwfEaCl2GSBI71KqjWYyBbp2NcuuFog8UO/Je
COKH0NVrsh1IRF1DoEd4v3ri8eE6q/1xk6pEz/AalUtBdTW6OYzoQvnCv+4ntsK/
o1Dov8QGiivJIiPxV5oneDMmcoqJaHNdjYDPeIG3p5+/imcTDzCfDNA6zMDUCTRO
unJgzJnQVZa/YIgGQyyE8n4vAIpuBrCJtLidfBmN0GwWjCelkVMfRVb+Eys/uNqQ
iJICcm+rJgG0E+3hgNM0MzOgx3TZiqxydOrBcWZm5sERDCvTwq/HtFvpWkyXr48N
HFuTirw/TqytXAwMTJcA/NDAMibu70vWgkkLHYp3GxudtsmWlzcl+tIwWZirDvPq
I3l8Z/zwP52XZ0du6Jip2/JeClc0LTwnHYbVpdCHjJ+gv0keFzhu/N9hNA/yzQ/a
+VJdhJ5BNIDl4eqtpMd+Y//qhcxCytwH4Ak/oVMZ9WU+hcpqT8flaszG8urS9Ugt
9Yg7O8fglk5SwSoJvOb2vWJTNkf5UaxPRXaRgD9OV4BzOGWl27kT528FY+RuYPvn
zOvHswOrqIachCU68NB/7iz2oP4Llrr1TWMV9prmqR1HENPFCKIKgzKEIaSsjSzO
1v1MTGoVm/SPBfqmXW9veeVYfiLMNuIool8004Jk0I9Jmu6z9+SY919FNS07TmsE
XZGW1AXKMcTVJL3pF6LqTnxnzJXj4RIU0THP8XhQWJMSFbvbKElY4V0ovoEVQcPY
uEGhSfdFEJwfIJxBOoPTZuPnbzXbY4Tkw02PUFLiaXkibdByor0/sizd4/4ZRMD1
NestOryZS3Rs4JnfRvm5pbqo0nbNFSa32WG8RYumPfCgHGFmDFiNwgGxuDQuPO0a
sxPz0Ch2UpWn/Znj7Yqczkm/HIsayy1spetR0th29JD5VIPkoIoBhmFTHsku1Voi
pu69hX7A7U35k5V4Nx2C3v0GT/Ray8lulGHxJ76nNNt2g+IaVsx8VaRwT/tf3Vtk
0qQdsRi0ahtb2bHxqN0JCZO356WAiab10qAxA2kpe042MIDJqTuuSnTznzFa2/lv
DN7SafyTJ/0WYnK474PHDpfwzwWRcZtunRWRCZXikanP/18fCWOo/uw6t0Vff+ib
hicwDBJ08LH08Rkb5zaEJfs/mmWcrhUMVxC962Z9p4KcUGKtZtPKbXEDfXrL8Cjy
3bBWuiQCZi1AZJS6zEy0Vxc71Qu9tINFjV+GTyKs7oT/2FsGi3Gi2cIF/E9teIqX
1p9aPBBLtOqYJfxi/GtWBDt1tlPn2pcccfk7N295aaDDgjtsycw7nkgJgePw8vCn
IjRykrHgtvObcgjgDHsOaRFc4yWH1pTn7WWKYMp+b5KQXD3CmaH3DTUVHPyyvqlE
bDJI0ZTcTeBOHA1xgZjegmnMpO4YLASb9u+ps7p1SWcASnxBE+XSEdJBGLVLvczV
x0GJdErAHA+NxuTAel4ZSe0ohsYpaMRf2hLjP0Di4ED/UxiC75ukdZJw26IFRCZT
rDO93Xvlj6xOswi7a3FpTf+CJHGPpRH17Gn3RKLeFB8R5EY4Wx5YclpFvBNPY+e3
IhMHl3ub5E6Sl+VosO/hpkr/P7Qc7w+ApV5UoZTTFPzQUz33bEjmc0CtQMQOO+Ts
dAX3jR5HZKyj52Pn6EGO8Szcko5Voz6euRLlq1ehaw1OhNGY91wBaOoaC+apIezK
wuKw4ojt9bSkb7CPDnX8XIU3d4MuA9eIgotbHUHLWj7rGiFaElUW52IDfwoxZeJ3
dgA1fvxQNBuCulQ9OA7+FrPlpphejfOiGpnyE4mPju7XMT58kI5iWsVQGLMEzoaT
CSxxedQ2/5EGMBfBHIIm1mDXtDKm1CpBX8th52hA2UT0ymK/kwoQ1+OwL/UDrybo
KqzJyeH0EFCvTEIjVZODMU8C/gMkyOqJTGoF1jKMDCx0wFjGdFtsFFUQ82E44GQf
vzNI+OgYNb5Z3a4uWS3fOy7FelZNqtXf0m12Q6bMO3FiXDPv4N66r0gxs3uFbz0y
KaS4769ntyvOlEOaVR7PuliIOM1Fhube6sqoqElcQsi7vC4XmQOnS2pezilShE1K
uAvDhX6rAdnjuwfEu7OlV64Hc+v5OrF0LBvMrDLilb1AMYpUaLre0Z5OavPA/7XV
vHMV1WhKEapcpWq+MMzoqbhEM0jjV0vrfItK2kw7sBU+9H/AP6LjpC4Jg5v+/9Lb
vZqen+Et7h0T5pYDWSXz05Ks4RdSFgWn8LJLx/7JtwKWl2e1uSOGgrwd1TGl+HRq
n3J+GueD9W0eH9dIy3auRGi5DOmsqBWKtwfStoKvSQ+VoARsbTFKiUvmczpGcnZz
Mb/VImbTVDiBQMi6KGnwjHZ/CcGnywiGNxiv3mlr5W+09GHhmf6CWoL9R3lijXcO
tV85T0nNwekOfmrfU8dG7ltBD8Y2EerL76REgj0wEvmjmCkGovks+I4qASNBCSPV
cMQumQov/jWRci3IcmnR3wIA181tj/89SSvIw65Eja+jiXlxgJeP81a4iHPLpYTZ
XD7QOdjN6TTMKWjLKLbTjTQ+RHtBQ6eAgf8oZKdgNz3Nc19O7W+YZwTCbd2cU8C5
JyuG0rgLpYlQfm9Y0spcq/A8YctJ0zS7l7u0DEKegy37diX8yQaOQg6AugxQdhyL
0iOhIPzYajoUmsRNmSF52PacyW69Iho2E/mMEqBudctbZj1vyDMBEnV9Z5jmPS59
WuAFxsVI399ANezq8LBua0Z1XSPfoyNFqL/Ks6E1NBdBgc6O1pnvk3r0WyQ0OqAU
F5ZXWjYGetilvqYm56H05SUkq8aQgLOi6CFYShEZGgmIz18x4BXXEw5iIzUUIcAI
2mlZSPDwEhOqaTSdOjB36TbH0WmKxLCsfRyAJFdbPjKWPEN0dE6vME3cGWxyHBAj
676WNmPLxXgBoY540rCYo8IkCJSPDGCcHcrMwavSKHPKo95vGNVf9N9DFchOHJj3
4uOYmTlKAc00oc8B18evHqZtQA87TTmR+Qp4Wa4IoPo2VezZqqoxQN30M5P+Yp8Z
8+Zq8u/XYptcS8LN4Yn6/IXl5g8eKdbyZwTF8kGqo9VNjrxGVSCwsQfX8vufh7YK
Y6i3yYyy1pBKNRpo+McwZc3Y5PPvyF/D2CupOpljcdrYXlsEH4K783baS3vZYV/7
e9tb0X7wqJw/WF6QEvDCim0Wumq8Y3oNv89i/APigSt4tjqhsNZ+6jferMiLltJF
SL5zVUtTeg8LjdI1u8+gPw4GzE4BZG+AMqzc1iXZov18XVaP5fp2QG/agHoxmK0L
SMi48FqmopO3h2BcdV/QmU6QBhS27O1IOyMxl+fhcavP1HwLcwejdT9FI3rka4iu
rc/+MzxjrTDsfrl78vairolJDv565/f2dDgTLyH2TgN/ejV4BJo6urvSEhlPi8Kb
Qv/znv/p8vOoK48HQiYzH3qEKgZAH8LWhpsKh31q2kiL+sHD49doXKKtlbGosdmB
ZklG8AmNn+Tm47RTzBqAHLoNpeJUFkKvFVd1uCP+lyLKWEq6pL9RyHBPyFp4lxi5
QAhXcnvqBnESTFpMshshM94zxxXVRK5z6aP99L45aiVpXNVlzE1rFcp3Q4ToW1JI
NcRBqkANmTCQIEDf08KLx4NY0ZRckuePMp2klycD7YwTh8FnL3saAUV6cbk9Eq51
GkimR9uZUf9P+uCrZ5awEW5MIVLGS5FN0eJZ7xr7OFh6+kbH8JfDVHSILV3XAgCf
EaxPRiTzOj+8W6iqwFcj2KW4BCqJqk+wasG4VzONanaE4XBk/FHRsEXXvxNpCSgq
3xZ1Hn4bJR6naip1zNHtSgi+YjbgixYf+a2zUxZZeTnqj6g4Z6j1TmvL1vW24mb7
8JgqBhuVjgvXdc2Vsj0l9poGtgFilf2DBbWSs4aihZJecf5dCdU0tnBHnWW9N3kH
BITywxVp2okgcZfe9kOZQtSDZ42p5Sl8yf7cFirQhrKLmIE3FuVUbnrJV+MX3CUG
SJx8kFQtaE/wR+EzNTE911YbmmUMuAC30m/F0OznY78Aib2/hMkBdyxYtSwNMpIv
TBrMmC/CqI3WKS4VodiSDFzEUWHD8CKnDw2CEerLTBHGyiy9qrOR1I2zxY/T2p0G
fY/KueVbtJJdPWtwjyjUHdIxE6zarmgUdSOjsOmkrBoCYOYCgPACSiWR1CZR/++b
IDgDBFLm1eFBLLT4FedbH3a3KFECYKCxQG48TqqDJvPpIzN5qT1sF+N5lOptyENz
4KBgakU/nBH8JdwRCb09iLPNP2wjp1eoD66XkBSjNn9AEr2Up/fB+wRHxhoxgw+g
mVKcWEMRArld2+6Y6JLhf8LdP2ySXlHdWWk95V/8jFBbuyMplOYEsZo/JjsfQLmt
GCFmF8tE9cB9KnnYzQfat6f4jsaF7nNSQDA5YBhZ7Ye2bp1SXxkBP+pmChRDJRXZ
dGVPqGyVhkFgZ8hEkLp/2MsNMTi+3HnHxyNm0IU5RqMX0fpjB6E5WitShaqcicQF
PuNLF24L7+G/2StTKmmxeUJUCTS1xeArqjoVecXdbjv+EnIes9wUs7JOa2dmEZ3+
fNtMBvFuI8mV/iDTO5fC1+VVuzJZcvL6emzoI1m9r7XxP3EqOJsKDC8/bIYeLKic
gaG+f4f3vwURQ2YO8XEROxP6tCjfXpIKJVdYDXm+ltBAX9A+wvppg/+lmB0tqTMG
1WbDLwHuSlrRnY3b0E36Ubo43CpBkqChKwHO6kTA3MAEscuHvrp3e0DRDauMrqnU
oQ7Gz8+dcRpy1vyRFp2sW+yBcpsMCwgtUjSfKyudsH9CP29GOAA88RwA13Nwprub
TK4fZxULZlN6J1jtqAdtixCT5wQzQvCtPp5LjTwA2lWA1BnyaKhs2BRN5USQjJSK
0lPEeY2ziyUSheyXdLxCbt2Mndkix7RGHgamC5vcO2OR+t+JCRfJU+WtMflL/npW
PARSA1fZy9lzvyLtE0FK0TSemTfQoE2768ejMhkGl7PMkejkP8y5llOJpGuXLXjv
Y6VafGNE0KLkCq012i/jhyjyxhhrYimAJiVhaK3Vf/m8seAYS3IfGHzaRuRephwR
Ran8ZSnFJM/HxqMjNXPnGV3/SXjRS3A2QnmCUN2FmCIxxqMKIcVVeRxCYDoIUECU
W2NttjWZ9yOnBVUGJ+6eRRGa0ycCzJ32NADk21nKDHujgXQDwZKlUkV6meZcW1nq
RS98dSmikdcV3tcqELrV5IB4/1v+qbagVp9FjAnMgJzg2oOiMXt5c6e0z7llISDg
3rjAPOT0yl5EauPVSAGaHqmr9WxAvkkM0nX71mNLtLEq8Cl8FvK29qVqrmKeGR1Q
26mTOKC/nKgM+lB57RauOGZtvRc7O8tApSO6hUycEJsb0to7XZ7By+S8F+M9UHtq
TCLgu5PQWOIANNIIBjDnCuVDKwvbcBIPIdBGKbiNIKmlSq3pEYsnUuxA9btSrV/j
K+c5o/3d25IzyXsuPO/ObSoeiaGLfIyaPt779Sk5iyYWzUTR3Jn+IUhWEf32PpO6
EPEth0+TO6ypt1QxwwF1K/yrzBmZ2GajBgeYyOJ7+d3aUIRr34l+QjgfNJ35Vbsu
ykX0fFcrCGZsITmq3ROnsLXRFLiFpcs1+/gz3T34ZxXkDKFozfa3jS3CiUcn0M27
Nusg9aAv5uk0SpzCPpgILm/fUaxEovMEQRXHny3GOAo=
`protect END_PROTECTED
