`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FVFEJ1cVPnr4wlJv8Spp6LtAhE5tOiUSJunH6SHa7x8Z9T0y9Gc3356VgUcQyeuR
azxvDus/LYM5oTTKNUulGwktd1OhypiiDsyGQBoHyyN4cjI0NRr4VWqQdAbcYPJH
5cbtsG17ciKOhkO02vvmxsdrWkXZmhNLMnznl5hHtLpdpEgbfuIJWyIkoKg89B+n
9WNFIPk+J2FMGN5mYrHaBZdvE/x3cpy4jh+NcaypVg4y91doApZGfHM2U/H4r/Mc
RHRQ8NrGRREGwmFJeleZDg9/uus9XO0iAPboZDHTfjW/iNK8nMUrmJZQ7ivu5xgE
R/HVvIXkmoM1b9mnTY/mrosK0tUyA+zIL9+3YsqHVvDq4UxygUU0BfrFdsyxstzZ
aU3H16qJKqOk9Lk51DLXua31zudUp74TG94cXhBTma6gTI8tlkk91D7wfgP0AJdh
Uffd+m+q8q0to26SFAXHvXfRZzS7Yy5kCZKyPbWzZLvJcUhcosWNQDWOX/h9t32b
TYLzU64caf0dv3Ca9AlWFpgZhV5YwmIQjJ7w5oU8Mir01EGtLz8g0JG+HMKI0bpD
2U3bNrosAZqPGxgyVP/0gCkmxIpYT2hh9MYoF5bg3xKksIhnDCAYjLGChcws1YO1
/uiB2cas3c54UnxU8mNXj4vZcHEK450KcbYdZqH1B/wARYNkye3+fF8fE/D4YY12
i6DiNFodhQUcSgUYtYjK62a0Nepbuith9jmSrNNS2KowMFXI4eXpLhl9hwPBmlSH
`protect END_PROTECTED
