`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UnSWdnONFLDy6zP8kqMYMfttYv3yueNnOV6x7wFEjkpZrxK4d8yehQayV4RTsefP
u7yCAZ9AcNSnhXgCQbM/LC3GIC7FtlqNkSdbKvX10SguzvoWsmHgnERdV4GOyzfO
u+03ZsiO/YCcchUNnVjg/9tevLbS+hR3LUVCTbGDzSRR5nmthpyxR5jup2r6E1eF
hUl+3KUK/bGkWtZqDJAKIE0EQ8vSroK2DJsect4vO7M4LRMShYWQYsy1ymOmdclV
W1ptsnj3EqVupkj9XdqcFfhaZ1a+8ypRLTWwPYafKu+n2jPexvwKAo2oC65vQzY0
PZqW/6ldsx93VF02piYCuLoOHBOVOGTlPtbntD8+ah3xRqnP5Vng2jMZCci0QQ3K
/wzhkXmoqJQz0sH7XroSYBhgvFl1gB1/DsoOQaLQb+NVVWx3zj80RvYdqOneSOFB
L7uuK5jy7hZncwAOgT1wfphBtFY/YnEizUsDqhX6EwwO2o+uwo8m9kuwu2V7J9nz
Tj1eWFRTXJVSpCj/EfpmraeGacsqIfer1pYB//tURb5YlHLwG2WXHmWa3Gt4UAsG
JdE5WPwwNIM8ElUtJs68DUNkQCWoEOAeXSDzvvVS3f9sfKS7VqSjfrsc0I57MOJX
u1H54qjWAD8x/mSpnbHv3+vAgfRIk33ADXjNO9JxrvEtYsB/QhHpwY6GUf2MI3/g
0lu7Nr2awa3GY5ZUnlu7A4zHrENGWTJd/MbhPNeV45UFwZdTUkJ6Rt0H8ltOSsie
Y5YVcVHguVPKhg0ojYwwrfUhIh4QRSVKoAF45nRSdBy6HofmlQMc2HljXachO+d2
pv8jflcExaYFoNzKX2wSsvpg24dbt/3q2dZA1ybDcWbvKelBl5AdSkp0JnFF6Noc
pfkw+NOH2KYB6WlwwkhxnzaRivhR9gzdrM4VfSZgskOJuQHs3BeDzE2BjTjSZ+Ox
HqCEjZ01u7+bx2iHQLV4ceSaRfR62lFz292GnxzOjX0Wr5MI/gn27BA9QtaitwYR
QpTILlOGSjy6sI2qA19fjduFUd0yviigdbHuZafa/q9jhOEnoiURKDUrfTy6Gezu
x05cabY/G8EMHz3s65XMnZXiGPDsqZaxbsZLPrgC7MPqZl6esD/Ln7pit1u3Y6n+
SjUfZizWyFSYHKjUpxHFYyVct/Gepy7rOv5MQh8nHT+/JtC00XGiBFuEONpVWHxH
8genVWwPuE7OAPCVdWxy1lq6G8mVPyXYgawiJqB/3q3vjm6XTjY7BzApCFHFocza
Y/g9NNWWDb7U7/DlYIisz/22YFRRlX58mt6C6PyijGfDdUkxxEsHjW92RTZbnro3
D3Hx0FnR2S+L2KFtkKRNqO1BEEWeloG2peH4VvZpAJ30KYaNu0WQ1OZyCSWZkdn6
SeKJBRBPtp1Vq4EJ+6SWl4bi7qwS6SolsOG9lsqj8RU/jYvagwiHj8KTeIRBPaAA
TJYmfSpXwUwNtrQ6s0YE+n0sV5CpgPuZKWrxt/lI4zZLCj2iSRZHW/2KizHvqBJ8
EqYPsSbPO8EPFffK1fUm2HY8s4nfNq/3NJOfzv5jGMEy/uxegptPRWfNCAbq/uKW
dZa8GfrYdXqCqCIzajuvhJWkgLncGseXmwp0SCpqZghebvjxQFGpyHY/mvakQMek
3HNUNM7iDAuiDpH/j2t7kZCBAeIwwzNeq1F0sjnEd6KQGBetsuYzMcPZDZrqQPQa
yBNKZnxROmt15M3SRaqzuRQ+lJHaOefmVl9J8cAtnoeXp/qvMQgE2MkW2ZvIV4Kp
1f9tI3KXSwrg3GjyeIQLw2FXBGVDWh8lJqaEuS5fYL7xCgm+/9lBsmsceedhnRlq
QdYwmckBYirZf2EhRiD5yByzFlbaemq/z03RIlrlGi4kSx1hEHadws+O+O2K5HDZ
qBAdEPzOK3rtmkj3xlu4544cXucxyhBDIRF4frbvoNeGfs+BgXSnUFzcqYJNlNFJ
T3t5R5hW8AnsVc9D7LKKueO8WakfhOM2+7cvnU9fJOmtzOlammExCJzwh22gOgx+
VXWwCUFk1n8mAAKs7weJKc+uB/6UaWPzPOAJSsSz/LbDV36E1tFLxLxwW5b36pG7
ndrFb/OGr6pcSQf+mQxAUxEwyW6X/d+Te2/DFFMFw1EfAKhu2rSOZMUln9yee2rs
KrU1kl/g8C/9jvd3x8NQQdGC2SaU+kqUmKpvnvvHClMzzMFs45Tcgfd5YhKjo0Xd
wuwVY7pnKBvfWOEzB/yF/i0oSNaoWtPEeR3dnC9XrrAm7F1AxgqC/D3vnrdBvESY
u/ye5bsLSs8KAeK1D5zrK40+ckl8xQFsNVTPwypHMQr2RqHgkpI93v720Ij5bf71
hmIFNdAXZrtV0bNAIh8+g02UiBFwQbWlkJLy4pm2zZeK6WU4SclpOMNM5w4b4Olh
PyUDtL57KDgSeFxCqLPKsusupcY9zubnc652kwZmMWIOQXJ6gF5alyyUbbzQbAN4
AxHazBvVl9zuSWdl8BvTluqVP/6aq3QTqZ6tIjnHyuA0XPwEGxtykQWRRnbpCRt5
TxMKd9Nj/bwjURkbh3GNdbtXoDl2C3Qz8MMb6aK1+T82l7k/dZ6/QNg67RZtm56r
LR14BqTSDQqM7awaqtoIOSbJLRcaHm7VIfQf51+ElKdGNJVGtEeRyNJqD8jWkWxO
wuH4Z1Orp6JuIszHmy+6N28hW7lLoF8iUqNGvV8kPBLLzXeIN6docKBH+UyHGwO2
rcP62nZROXUlbN1Trjwsk8Vg16WbHK1XhhOfvZLuETvFJAGOegwTr8LRIbc/tIfq
B0w6RJgsP2grDD3LgPgzTPVQSYaVQvTJ/oOdCEuTjD2HaOvI+8rQv+i75OX1CHDT
uegnkwzWaMRypaNYD9VDPc/BpZL/c8NZDcsjc9Gr2ZQRWjXLyY3EED4BfyKw3es7
wC1nWBuSZO2/J3uJJWx7EZuf6FKsgkP5Bvwe6NkBkTTizuQu1uouJofBZeb8V8xk
78YTLFlhQR7YjAhqtooaN8pGWVoD+62147llVxyur3g31nDFeTQrpuWku2Y8kpGg
umx1R/fplX5sHyCnhiTRvMVff1asfp94UsEQbGoYYAkdT2OXoEUBEC16jO1dsVpv
RXvIff6rN2YrOYXYDhrMGjxQap9Fh32v80E+lxzs8IpsqdejgWkgWvE086NbHT5i
BQzVJkSJsQHAbbhiqXli+AOGfebRUSpc+Dq5uWUoVluzy2qWYDXFNdjU6dDu/TQN
avMh7c3akPFFSQCEhu1AAClFg9OcEdypWhaKAh3l9aHCamYQqpLA7GarN7X+MLN0
tV20PJXVSIicX2kVvcW0lrbjt6u9NKiPaLkllvkEiJmIGID8bCbxEwVj9+4ZuxTc
wa6CzFSUcNziNwPnKI6ZYlh2Xi17QX1lSETgyKunDZZL8VU+MYSz/wpjbkcBKJIu
poHn06CD60jbK931Ht1iwYkFU9JyXvzuKJewcDb3dx52MSPdLbaQ+Z6tT7TakgaV
BIWVQwF+ozdBnUfhQGFGIQN+KgVcndrf3eBjUWbNyqrPWY+FP2zL8nURRa0W4gVO
wWOWAHLsk7+LJIEDMIP2+5w7T0FdH8McKrZ3hUB3sDhf/1qtAT/J1G3MkstYZVBd
yO80/qpc3W1XK+VFLLXdza6oeysgUQsz6TyjHszsW0OFDK1e+AfjcyjGsKQ3KLl9
46iXGC9n7amKCVVXlCWedtXX4tGTZZ4ldCTI1laVSmYuPrj9VWvVb+91UoOCBv8d
3ZDB65FlAa4Qor4MgdVV0M9I71UdvUMWwZVXnrYJ+EDw96AFLwMYGihA8HCASUfR
UNw7A4FYnPqCap/i+oMNievf0gCY1QidqhzGU4hw2tkVtTMGHov/t6tvzWIAwo0U
SlzvaMRV/ZT6Oubtji0zhb8IlI3Pz1+MWl3qDQ4rwX3/m0hrE40UEhCl0xMWvCbE
5IeDa8mhg07XhSAXlY9bXYap1/rkO9A0u8aHaHFyRBI8EJ0xeqvUIkbPmvtmKIb5
GbmPuABSZdYVF8uJQXv5I0xKfxLkoZAbqlilXIpP3XO//KaedzrJQn67F+Fl6fOO
4MncMFmDJPGjxNOpVbCaLtiLbGqopay6g2EYqxqKIOPCPBBByVPvfUC82pLHWBzy
S6FODyiN1ke0+gIeKYMXGqSBPKC0cR16i6+8+lbJSUxWPxEPFJUxx70lmLshn3ne
EcGZMaCeO/JVr5kahp58FfhEZONWhTb3Cy4WQlz3Uv+eBS/5N2WRTf8aeaaOAZ9G
LdTtNpIY9W4IPlXUMUzdB5FHkCeOBqcUdlKOO7ZuNnsvXBfiU2DPr7O5M0oKKyJQ
KaEJZMbSMVT5Wj4KAERJvC/a89OvkLRS4Vsp9XIBLwgJcXOZ2WTC8kOEzhMbkqzt
r80no764trRdf42uNG4QIy7d6iqgvNRhGMeD6tlRyB4uJrqka9keDIeCMAtKeDF6
sbc20ihpH2Q/UFn6Ic0zuZo5JFvmUJtAogJ8PXKoeKHY7HTtFeJFQrWVwc6pSjH1
SIQ9wrSvBJV+1m1O36wjbpcgfWSfagyykMFeHzyIaqUZWVlYOgqg8VwIaAL+R/g0
qPWbXJ/5Jf42EIzBLG608hBDgwEqG2ZBLt9Pe2RolLc+u9LVNi2qzdGgUuSJqCTo
0i0eIn6Gmyb0a+zq15TlfZf89qGOdZT2lnXzjGwaVdmfZbOM1OISQe73fVWKwDSQ
JmboG8GPTF4fOKHbC75e79bY4zFEvZQLbu4mdwuCbAoNDsWvi95NXqg5Ikv3Mvcp
lqN8Q+VBkX8tWugBnCImaL5V+k2GaqVBANcRQnsQxLCRx3IVxJQBX05E/MiXJPXv
exgO7E6QMZqFzWpncXjo8zqm+ylI1I3KeAeZZ6FuueOja2fzmsY2bxSqbptKWQLV
WkhMxSxt+yg72vDcIbWQI1A1+cEDWaz3sEfYfh5kwT4Mb4wMJiX8EgPC5qNSBNeB
iPTO4RW8CRGKB4SVHzSWxkJzfpyAzYdqRw7/MuWTxUnTJspocRwvhXYxm/Z/pJNv
3rl2KAtwlJpN/Ja/vyKmfyUvr9FFV0Ak+sM1noVuo0W+neH6CVX2KP8TlEn/U2sf
Tp83HccSi8VVC3ne//U+8IkMMlFEny14kZpwMNFeTnHTxB6haE/6kiO3T2XVyY2/
Z/3eW3z7XdAUlbNxREN0M0NGQSje/d92Ut6N1WjOpYnzdYn/Oz28jw6Kc5Ip/W8o
B/xUQdWcCV+jRC62VXwDF7TVSqsGU1BJt66KkPqCLNapekflxTKP/SIp2hvfs6jf
9OcQtmNaITcZ0ZJQGB0YUeBto9ijEZIdLe68DVBtKL/a77Ky7Ltf5mE1sG3otGMG
ukSK6pljESvRF03fxErg866ScATVS9wrotr1e4n0pQORgS14NKVr7V20cVV7k4pU
G5iDRCtMuZWlTlq7ufq2oA7y9/IUlCDE+3e8zHiLLBgfJnLITwCbkly9X15x1Rvv
D7RK3zfcMLO/ulTvmjaTNQL7+wGlVPD9Wsn4RRLz/2cW6/vYHEQAoCFPqOvgeoBN
tCg3/TZ8SpIIK/H97QFj8dCz7NqyyxocPanW9feCex0Fh6FfA4OXYTO4ZZ/PGLTB
sDOFiAzZ3TKOSEQS9WqczGddh2xvykDA9OS82Fl9yuy0xLj4ZGEjlIvwfvOviHYP
CShteIX0xuKIIx30xkled5RA1DQw73AUqzdvmcL8YA951jERXN05wiZarTc+jeOy
hrmHPfEfA3UVUTuoOogmVNcX95Ryi4ltLMocti0tfvhoKoDBzAiMZA5xPkwMGp4V
kT/uiP2vtoX8L0Ztv6SBrYrYl6WZMEsTOGOKYSQeU7kcrIkFndfD/ZmZH1RQEOBU
6nkcaFoQapY0W7LoPQWZNCna9Mk3KClXlcFyD3/D5w0=
`protect END_PROTECTED
