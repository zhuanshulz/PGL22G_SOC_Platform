`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7r+b/HZRD0JN37z1aeTV7l8nsRnFO1BknSFhj9uw4K+/REgkPFIJDVgdEy6bRxly
1P0mWE3aTPiA+Gnqv52R0Bfe/H+qn7m6c5yjQxMsPn8ZNqm5svaOf2iw1ppo0edE
2nE7n8q2PtOh6gkiEa7ucaGecWFfb2JicbFANidg3OCghcaUxNS0OcWS5+eAeW5p
ldx4YWFG5BcisYbWKO3IPO360v0+hEe4V+Tan7rpRPMG99ZLn8mtvmGQu+1Vnu/3
UG9g00my1sga+hb84LPaWtd4v0B23xqI48E6LoAIk0pV+038JjnAxujsVqTRxHVG
oPV8ot9OIsoScSbTFtmzjGtoSNvFWWFzQ4/vwG2kv/12V2qwzjhbLmvfVvyidWQd
gyWyz+8Hz77VvIWecssq1606pP/wJBVwGqdqje/4z1mlhzHQLL9EvgwWTojd2PCX
ARa453jyMDL8M+wXSdTKozMZhpDb31cMQiCNVLTeNFnJzxiF7n3NbAzmCrCz5IIt
WRFFR70XwKIjNSIvTNx1yypNR9CfNEj6cB+N4pMgZhkbfEK1rP5/u3E6huFmBm+c
FewmttBVjAzMxquliH1ha4Jh5zHAXl2DrLU8V+IBo0/72rHMyf+579Nyoam2L2mq
GZvlVXGQBcC/yGE02YLAVaCcrLfu6LerM2HdFDTat2CizOymEmb2xvZvq2GXoJVh
GGIRunyH7t4+jmnPIz3d/BL19A9Sprf7Pa6Twmvq9uAr5Bkt08UsonjtaYCkzI7R
g8QVpLP3kwplVsEwNoN0ytlzkSI5WE/in2u8xXMUxaCHQSA89pWyQ0UYIEXhaLIC
hYqfi/ClP00MEVJ5aTWGS9IWVd6iZGq6sQvqalTam8xHkbyp95M43AuiTFwXQw3O
gowrCQBX+BJRNzYL5AtX6zm1Gi2UtRZllQNOR+CKvETx6sQ1Ab4CKF12roJYK13U
k2DDLwgDoiKRxl7i82fUp/tyEU6MFqybua+vmVna9poq+F8zbTfQyfIpmAqb8f7y
TvXwi6+kwmlF9wcoGi98Bi28XGaJ1Z7wXZIWEeT5khgZ9YbpNPYyThtxpEJEvAWO
5qGLVMUY5qjVJX3VPhpay/AHVGSJ3dEzoRDoXGXlphljZlZhczxmI/FQbfSVj55U
4swOu6GnkYZ6mXExy2BtLELv8azlUJ8ohClkYniY8aoeeh+UERhuIRikPpInY+zf
jnvczaSjQtgGYvDsTnVCE3jgcfSHh4Fk8GCD0a5pZXhUIq+ZiezG8F0EKXvA51Xs
I7Dfoix0xUAEnOLWyPWsM9JgdT8jvcInVA52j4Z7t8GtF2O2Q1/YhpbbYFn+EUJc
`protect END_PROTECTED
