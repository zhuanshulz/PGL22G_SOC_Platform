`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uRTYVaTq0hJTB2XYjMbboaxPiRRUuCoq1wUtAEqmKOVaP3jJEu+PGIKCL8ziBc0R
37XScGCty/0JcNp9UY3DOOxMB2PU3a0RrNOFszJLOC/bCq8SK4EzbeRzu/WMjwy0
VzRBg0mqt+PjeGzN93tuoc4S7giTjsfv3zsxO4K5kO6zwnthpAXrHQESl0UV0Aie
y2myQd+sZkv0q9y2FImUh8p4DCLb50D5ICfuZKvb4TmweZcu2GEj9WShSBn4XE86
cr0UBr8c83IRSpvGwLj/wx8NqdxgVCm5QJI/D6PLs7qdqS9NO83FC3+LgIPP6WIB
/sC5vQ6SF9IuO++CFzIzyUxs1ix/esvLgV49H4Vb2NGqlb+5X82ZmY+3GjpEx+GM
VjdL8ycBYs1FI10L0x6mEjX5iU5/zonjVOudZK+3B2XZPwOjpED4JO2+o+QRWELo
H14Pe6zuIhMDl1cVrFHTPpHr2ygX7Umi6nE9EuXVWFoIerLaE1R9R3G49rEKYRHG
DSuRB095xD1v7/4nFI31UlDHcgU2tlbfNbvovfcODTlKEuzhgBf/MqPW+gH1WmYz
0ZGUDICWFCLzjm1MppDK0djPOkJZYLb+ut3M4TCp8KO4r19BcToHEtXuD/Zb/gYT
OJgDoiCeNflxRqLa8JleynJhSwg/HrGCR3OXCEwzbyBA0is7tI7f9dkrEl0yqn9b
ybukXpcMiiJEpTlOErmBjmxjkTdShCQGONj+5XKyHRdJvZTaMObSTVVuUyGU6QGA
KI78vQRZk2xJyBLQMs+RfCPvj1mzVUlUirVCPW73l/GgkOK2ftxndQHYTA+FmHDB
XLt4EzMhNVnQzReaGRxGg9Bu5VkV7W8ZqEWEjmOkYXee8haf3zUCoVtB+Xv21Xs1
awrECINF/26xNEFnIhpVQaekfoBhzNZA+7ksI0aIEUOyHp7fSme4F5LWWAb3WOlF
cF/LjavPSAZlNquY3jzI6e2KtA6lZYiZaDm7CJ191h39HNC8g940V8Pv/aTZUMOq
9P4oU4uUHsKYbksvuy9UWSNLSS83EWD/2i7uzq6nbogWat6U1ZG7ewa7HQ6qHR6M
t/EK48bHSq2wVne3ZhC33xsEKqV2fZyyQUo6oH3U8vMDPnbvSoyjziuPI0XHWIzy
l/U0TEPWmxB+R6FigFKk83rzfFdkY4N+MDWjl7gkFcTIYQDbOSwDFKDifoiwWGIJ
7a4kQS6xbZ+NH7+rSZfniadOPx8ir06UV0i3VR8RzfBicFa18W/MXYTNlZBTFzpu
h7RWcCkdBLGVnjJp21B4zfuuAq8W1W+V/5T+zlSd0QjYNFdE7aC+HDSW2yGb0UOb
6Xe22imEYh0jUgk2cJh/O0lxNFv2IN2Snm2Ha+v+IEnswnsstdq8XHTBL9fg/btO
CiHcBaOTbe8GmK3bPYBj/ZvtMeWD/RGwxmX+YhLb5M49ZbKXBGuAC3ddMrs2KE8e
pGGR3rjs0Jkd669ejuz3yH3QhTTRsGF2vYPemUMD769eNqBg7M++3Kw/YL56Ohwp
AHaf9JzU+ViZB+mXgVfL0JX8YUTm0on7+sF0ns8hRVXpbedYyCjykBfwJ9mtrrsy
1gJt6ob8L07F+apZizpeZ18yuPrpUFwWf/nvLHJLrgQqp8TQKsxw5gnpI35qX10s
oT7VRake7VQXiQUjQfxNhHqb4lBIAJQCVlE9sCeuJOf1422pAUFKp1fIAZ/87AFP
l3fwz02GZqYZOLlGy5JAD6ehlQk//Y2YsWKCcmqyg+66uwe9otEBw5Ishnw1mgaK
+VU/HqC6Q+Favh7AOcn133VeHMbrRkiStDRrNkGbAr/G1a4c2u8g4DWIntR5MiCi
OQ3jBnpnEz3cVk3N3HHje9ihHufKaH4GxvoyHWH23cqI50+ZTx1jl0IWH1KhE+75
JNoR6ZpsBD/zCS8PAcveHMYNKI18SkT//M/Zx0Un1zTmg9CiIQEfql9LDPFycBhT
7OMpNB9br0b2pexnUGwJ519bv8wLEBkFZulxXXpKxOl/uuf1tfBa7ASlv4887JQm
4HYycOsIXhzCrlyB5FyHgleIa71O7qoclza4ISFEWttHcvFhqNSzS8yxd0YUl2tp
OeZDHewmhzz4sRKSdsrMTazl/U4S+rc+kZmd5O5QS9Z6RLELcEB1W8J2IpNvQhD4
RmKy9NsBP2iPjfOssRixA/hNPFxXeIIBOzBUaTiWkB2SC1n1bTCpnNEsvxZzyMQ4
aelpD73M4SyEo0TvurG/BGBhkM3//1Z0D5wEYy9onhEMAJrGYKbjAEx1kzd16g5C
Q5/KEV5v22vc2ShEYW4oMN+lLcpVO3ozwqdN7Icchf/RJdBkq7DBrteHi15w+eDC
33EMCaD8tlpeWSjMQ8N22byS1u0ExdvPQePFtE6O6wzWTHDoaWMH7A2k7yivia9s
ZzqNXetsExGxXFrml4zgbCWlySzbjmh0lP9KqeEHltl487Ew7WhEUPhf2U0Kkkwy
1KhxLQyKQcxhfTAH1Se9f1mLLSEFb7pWRlD0ibrLzmsRETDJfsXbhB5WeQVqMdW4
MOFZ86lW5PRsGiix3hmt3n2xqJrX0pIi6aq0onLuyOaLlLbWhsHIMPTT7cC7mb+V
06YC1bMvwNCM4yJKmHkRbKD8pMaEFoMTJPxNuNqhauDaoBWsAD14CQSRcUFwr626
1Pk0DkakOencz/Js2IFqIjHwZvMtLlNdqNfJcJNujomyufTCAq0fkiDRaj5lscOF
XgdsUlrArue9TiQqjyTCwbCNFot/RtnD/1K1leyKYKd8DqJcOHQ4F26jp6xUKe3r
fxVQrzAjRAjKPNQDLQ2TohC+l3yyOetXZZ4/Rdyv+wGaxWRSMoZFG++4F+EwwOPH
j1Vf2nZ3QSE6TKVFVkSQDgBQuUeHYJObGjDRpK+NsrBilCZsSWRg7MxkewFLctgm
aqWfNTbHRe5vzJOOKKQVUWwJYj6z909M86GDINR0tpJW0VnFKh7xkFf3HigY2Nkt
kx+4q/hKezTcL/pVmkEwdAlDNGZzp9FuWOLR/w/vYJM382pMDX8W4Ek1GJnzmw1i
4+o4IYYNQZuMsSSwHyn0HbVWAMqyG/ypdZtqMr8luTxoBxkZq+/lIMsoqKVjVaVV
OwMC+wGAyEVT2ULt7talKj+kmHjLLfaoHUKHad2gLaNL/84TdrHKv21Jt05VxrM/
ZyKgLeKWWJodBl69PZ0ry9vacPPgcgy/fUdU6PAQWMg=
`protect END_PROTECTED
