`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vIkHqwjgsH8Otp6mQ2Jx0/fCMXdEdqfT20xaw4NN3EpDgVHNmQOM7GsT9O/Hs/Yw
rLaksiF1VLNbPluPukmTL8Awa/Y8zNNUM+Fr6mlvkUx6Hm0kvL4N15LzJ22HHPHa
bXlYEYZ27Sf+2B2h8m6RGSJtj//hD8cVPxLCAohL8iDxm1MDQczBPVdNWFQHpB17
Cle143Ne44W4OE2YdRkJYFxHbx3EMJqUWu0708NqnP6TNSqbver/3va9bvwmcJiu
SeXLiVUkt68Q5/JPO6ZGBA0TnpOHAiw2Dl4d8jjTgZphg9R7hgu4kvcm+tfVFC7j
s9PvbRyP79LM5eBcH9q1zi6vso+dlvEANLMwFUt/yJos5IVzOuAhHiUZ1J4WdLI+
0UmvBB6GndpRXUqski2BBHOetogVgKyU5Z4KRpC9hnlpXtZJQKgC3VywEzpP484E
PyLtstjJtOJXxiGu1X+Mby/6cQH4D9jtD/r4iHZfD97TFLt1GBRjZAW2AzIY786/
uHtwgvIZtBHDXIWwCcvDQQ==
`protect END_PROTECTED
