`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JA9JPIqXr5ijUrdNjMmBeNc/g/qOqcavLfnV1f83TgpJlwAY9MRgC5fznPzye3x2
Tq/a88vHefhfxuvd9d968oHeamSGIkRt/elyUaE0x/sYboXW1+JPIYRrsXaE1XHS
cT5a0qiPvKWHb7HMI0XtnZgdnfbJfHpXsyBhUplW3zkiPlGVZ1eZCsfjlHBPSOrp
bnWkyECMoat2eL0Ng6GqpYb16kK2dCuij5k5fZam8fXB6YtqgFwO0zdFW3np+glL
8YBijpIWVKoWUY+g6zedtc3VH2NBuORAeyop92tuwWINs2EnfAN+dmebyyDTcWnK
ZOILR/0QQVo+iQaWgpCpMo1w8f/P+5RueJbeUN8Dgz7ekIlx3KQeRweGUxvY/U7Q
m9Sz65ahoTZIPl6GiIa3BDe1QvkONK+BsZ7IAgLUFMw2vKb6gYJ2tu6BPAuNRvEE
fGurwVDMlN0DXLFTqm2KvsEk8K3jfYxs2xWojha/ueyH+zlFokVyH7Cbyw0Mp7t+
q/osXx0LV5G3h7LOOsfARotnWwr0L7iGWnlVynHX8pL8l+VwgQx/nvGxaIM6xBA5
J40ckHGmOQ7icassGcuEYyO4Mn6as15vukomNGhkF2/KejnNvQ7rjeA8zTOVM4YE
m62kEa7IT51isQOwwY42VZkroqImDLHf1NMYWKTq8aREUyJYYqnmLbyVVLmX1ED7
L52C5QChPmL9vKPoGwFqmhiBz5EF3sN3IhpbFAc1EQSW0stAg8MiD8sFEgEem72a
+Un4z8oiCa2CD+fFf+HIkwQLHUsyF92GrMvS+3sLnIcX/CjW3UTD44dhjvI+hRF1
DtG78jrZn9J28az/tFRvDG3hQuC4u5Z2kfal0eiU0UPnUbT2U9LwseLknKHNivSy
LirP25xdOKSBLEtB7xieofeACdLRX3DHlzWoWrRogyG9B72Tn2naX0H1cYMe6y19
5w0buWauJ9HvROzzUrFXew9j7X26O7tF4EWujoJZz/jt5/j971a2dvydf+7PcEz5
GwgutrqySNh4lryFnbkMH1lO12YMR9awiBI4LVvlfBc5awHaDLxiP3FBHu/OnkMZ
kU26drQthDq2FGqoqXAfYRFvszISg1pJWsoHle9D39rqUbc0Bp4uLthM+zdsd6gq
xyXyOp/abL3Mb+Bo66spW1KVHE4zDDSe1AVjaWmaTxnkBSVJ63w8IyuTcx++3LyB
wokIG4Pqbnl+u3ULMPMJcvsIYDyCyBJL2xnpLSTNH+M+fxIyLFOOT69dXNgU4ynt
HXYDw8dNP+oK/4/YBha+ByVrKIwRk4IXTsuWOYVBJBK6EANbuIPtY7s2KgEReCoM
pA2+4KLpyttrA57HMTEEn45VfeDt9wiuEonpqLCYUkdwpWP1eolWwKI/QGiGLNg2
dntAGk4T4hr8Dz/9LgS2ZK10lCfac5prZljk0bU0KrlIm9lvG6FUO9EyFY/sn99J
FHExfrE8kW5wO3Z31CARk6hoJgMeH3H5+LXFIqpynzMDRNU7+PKEI1T7VU58irkK
4dji4GX8kOBjRXOql/w0zWwnChgtAcPEc5kS73p7WRM8O3owmuVN4p6RbMqNu1db
EVZUteav448fP3HDH96HfRxv8mQvpLGv5bw3XVUtCWdv9Cz0WIho/3Sg7x6jCni9
XvrIqBrfVfnWt35xhPWfaiMi8f7K5lqw43yNNA/tXh1vun8I2H6mlAe+7Bggyx4x
SS2WeioyT2vOy+KoCsxg+UMlCSB5spUhAuufB3fnNt37gtZ0zwDhBuxk6Q0spHy/
0r7MK4Ayl74y0NW10ywbcCfuY3+9l7o/Kuorr+EjPkuqP4QW9lUDfEG6wq24aMgZ
kGhIX5H0dEBEc2oSXN+/VmxRgp8mOxjRjewl7w57+e5s2DpEfb2WU/1bOfJpNGDZ
lQI4UT6Pi3MJHsUksDgEg1FQ/yDUkqJIqxOcVMCFw2Xoat//4QyDMuypmqhE12kT
2S2yoDFA/c5q9ihP9Z76byeawoNkmFQunOKS3xOO3facCvilkQkkpUDUZ8Q3HxOq
tpJZW/ryOdm8rficNlbrGkRjOe1NQquXnIYUAqAwvXdpjUjA/JbFmV6hhmpH19Yz
Z5vaHLBtcZIFjVXr5GkOXWvGHzXki4CtMubkMjLoD2OSHoNPY64GkvsaRTmsNcQB
EcHIyKdou66EoBc1ZSfYtHecPYD8ZPOgqG4lrA5KywyQbExSDzgdRhe0FFdoRCUG
W1B0isydaUc2wh9zk3s2ab+L1+WgY6+HSvhmhfZlJSag5I6+PYWlKsHhcc0xobdx
Uc1NIpgFV+iqlu/wF4ZXDn6zKduEYzz+5dO73oLtgwiA0MOzBY1qCDkews7UxjDx
M8TI6uD5dRte/l0d8jQjggKD2ROHDKyYDNSCJqWswpbJadAF4dUp8pF0/TSXPC89
n9vaNDn2FiqMxRkzVnTWYMU4cnwQoNP99HlhNLJstpFFlcBFLpdCZfDdLG/5KSpX
guEeORSAXP/QWd3T9adMo1nTeAM3aDhcWsIwJMzJ9DwWU0HhjOWt133fcp6pqjWt
+NmFttlBYgTcFPg1g8QMH/58M8Ybk8gEhhYgIJLzO9hMV+7V4DSV6Re2P3+OxQIY
o6JnqMjO2j2HONgARvLnDapTpMhSeqDnjccYr9CgR892aIeuMKl07ydwlZFd7mDY
BBBPtj6nCIGDyGboNY75wwoiyz8Z4NzSf8k0dZyKZj0C2WmSLjxIxG0DAnXVKf6d
5sRnGOXet/RxTN0wnue3gJm5ZWcJzWaJx7io5sK3YerRBRx0VK+Xd+fUCwzI6Xl0
3CTMcFNR/19lvmz/2xpPeHvqDfDlMUauMd5Mw3cRTzY1XTyoaz2o8IqnYxsNicg8
xVi9snb1Q/ZTLA5644v0OMt9+DHBPhJMvul13gRMX5G32jktI7yH1yjmDWUMWOCA
mo2o0t7wRDf54k0Qj6RvcYAF16hKUFzNvpkR9Ci6xj18FsUwErynWH8gdEdnm3lG
m6faAkGTVxAOdDqIFc+Dgg2E36xfvIIuU6GPBMVdwer86j9U0DXbA3Ommab/UhOY
0Qu9evLPbio8ZZWtG4N21xfEb5qnJVz/c3ZdCLErW4nqiKkFpz1QFikNJ7uFyGtK
a2fw2qfrWnmR7WN30DczJtftPLf4p6jqSBtA8ai9rEBxxwS1PQdeX7qlbxvxM++1
jLjXlwwC/QLwXraDWFdZIaz0CuzLlXhfVJi3yAmYLAYlKp184FyxUajDkfSz1Xid
q3Ha2Kv8Qq/uLqrjdjNwDlEt5UJZvzkIHTbuLfQpr3cle+AZZCec4qz8wBuhuasJ
r4RPgvsoTE+lXm0R23XXJcW8p1aMAw8cbnpZQcfuqEg/NYkfKrX9DhbQnrJhC0Q5
1Qnk6uSIXry9NDM8Xm7whPHtolEPEguH5BhlrJfMlAp/idjPZp4QH9JNjeQmkBtS
BUdN09XO2TTPEPjSoKBPv/nKxFyk9hCAMLX63c79KEtVLCZHQasFqEYAbIOHdrtd
FewyqDuK1vaXFeBtgcOKp7hsWmUgYnTLAaAiXgMaouRybwuI9/sL8g2PB+jiyhe+
OPnFiJqSCmhU2qv0vqXgiBrlIrZN31xt+tATifHynweft4KLzHo3kOiBtpkL0W3n
86wg17b6tV5QDLJbRs43FVeJVJ+cIY2r8X3+jvnePnRjDMHPidRIRxe9pYAu6KK+
ITgniDGE0/00t8UoFMa3xGGUl4A0P53WzhWZF4+nXxJWD+57GSplJpnL5VEHtbP0
5bO7zsOrkvqYcpm9Z7xsjrV6lYb/Htfip80B3vtF6lGNGUpEbSm9uqxC/8VSvi60
34LVwOYJDFcMMvJwvwQ1nACdIhvTuud0hGQyeIDpBftCTkhl34CixL9AgTiAQmfb
X52plLFc5ww3woYSUl3XkmiQB1TgshhZzXvmZGb9zkQf3eSgkPwdD+y5lw8XL7bZ
q5PJU4qIoyz9eRa/spzD2qerH1gNzenEJpq3fzV6MmcXanuw5NE9MTdEA9X3ip0F
nFgKLsA7/2We5xXNNLkhEmR01Tgd4312gbrLwPUZjfsclda/nqiTHyHW2w9TWK4H
8LJ6K9ovlMFOjquwxzRIWoRmtwYMsaggFwlvPAs4zH04100HJECx9CBzOz+dX+Y/
Yh4ENzo684gtSnQ3p40DOwVKx3l2IkR/N6bXB5TIXiTnTnZZT0658aoeV0J+6J8/
6m9fICra7vngG1sO9aKjIX6ZO4+Ppsifp4t+TtxE00mcQcILXnSX5PRYdLrDUfiS
nC4y6wkwLBrFagTWc7WUGBELO0TuZEeVul6Y8cncaTmHl58ZPrS4mlLrjYIK74Uw
Wzz0INmwTpATxrPyDat5/l8Un/yQ3jXh36JIR9RqGEBqm8hZBgHNzmqRLtu0Griu
m03wr1p9lJHCDOEHlJd+KmoTQwtJmpXK9psFFvUP3T1JtBPW0+gT+0a+Mmk6yglv
CoV7nP4ypfW5HxbV+r1I32PkBVMYW4XbdkoyHubJEnDXE8897wNDJEOOJHyQafND
hTZWP/Qla+YVuO6GJ5BC4IF67c/SXaRJQmPAx9co8ENIyIOdsIruVIifJJMDucgw
8u7n56fPED3KCjXVMFGNYuUH8/lFSyN2P0pXDgVfjtMAOFyZOsDIK4uxG0cbAeSO
YFP/gJ+gIOj/mhk3UsFP7T/1lOA9TSTRjlsy9iRUFUPpjyl2KVhzwT4LNyEn1+Ez
DG/u4rzoem5VjMYjUeIiybn6+A7IZef7WOfE5BHNxZfuD0hrfYTcHc6Eu9dqUmlG
djIEzoPV46X9DIOcDSv0fTGvSmZDjm4xIfMTAfla1zi/fu3ru9J5g9ToXQM9dd0f
pVYruUBsOj/OiMNwwg9kVPA6+q23h07oRQYnO6I8jDA9kyWPEHg/MvsiYb7F1aae
OV1wRS7CWH4kWrEjxrFsPZmfYc0PL0ISACCfEJGFbEGKZxNamrnt4Rnvgtnak3ZY
jyJjm86Y2geSPNSBaB1ktntnaM+MnpXNSqYY19J5VhL3k88xxKHOlBgTGPIANVJQ
iYefix06v8lFyKDOsU1a4QudiDT+tnPmNuljbv9gu2Vz5gnoeS2p5mUZaTRS/ojY
52WNWuPvZOpoDhKwJdumvZKHTC07sOTj3nazltfDRUmeJaTU5oAloU6rUMSQF65z
4ObAp6+isK0b9kkoSfEBJLs2LRp8itKRjM6EmiradosFnzRoS2soe8VY4e/g2ioA
nSaNttZEfrH8WXPc7R1KrzvsuZhX9DOyZERp28Dj5uamqvwjklhmYZUcENVj6GHq
7H/x4IqrDEFbOOXCepBZd7RojHpKeeQILb7riNrFLDtVtPivMr5O06JVbHD/TP7A
g7vnrr8mAY1UYsi3I/s13bRlmInIff3LaQxHGe8ZO0pXCXDUypVw/Vjd7J0ATQ4W
e2/SBsibyHsHV2zs6ahiVbMs+iH2/VcMy1Qlo2T/77lWXwFpFOWrpDFydkauFR6g
hTO8KWaS4HbUfYV5/rAQ1hen2AhtQAF3f+eVjqgJHde4EjJpoRkrpvTbkYV4/mou
/oIDIO9EYnlTbPqTojDV/vDEypBq7puGfANJuVwFFUxaVeRsRTd2dhfVbsSi42fZ
idxAedLjh21cx+Bf6+jLbRxUAekJhBZiGLJ8Br+EteA6jFbuNW5k+jUu2EmxbYQI
CEX6siJCA1K1cszUVq9aWItqd3qD3XK9UqchtNwEWtFGSGBoajnL7TQ3pqGypiOq
/KaVVS/Mdy9xlNouNRPGg8ITscD1/vZvnIYiKIRi3K5EM+qvE9unWEXhTo3AkJ/A
GsGQtTmOLfV9WZccSx148ms64vCuc7xCXEFBvtg2yaYsAI2yDE0YcsSCgb1CHViB
xKg24XulGnNGlp3ILDubZ185G5eSg1EOaz2CXIkpvod0LFl7rRP3XJ+cc4QKbEpu
X0M6LJ4Y3eG0aLJKeTui7PJriWKqcuwEScpPjUTx/8XXbx9hCS90MUUfP0vJmVVc
JyVoGKiiABA7utcvpWrz3rMgUjpc/UAuPzSwEUczrkz0RQWpvdVeE44zN6LItpKn
Lw1H7Jr7GX3qAaLpMDfbpEjH1vP4d4jTF3/MSXG43HMRBtJssfFjoi0za4GmmBm7
8nPYsiL1j/Aa9prDiGjyOY6xM7nUxp18HjU9ZFMdxnXlGBQt4FmcFSWFUHfwXlov
TmMnQd9WxbHcQ/npxLs9SB8Sm1QgeXzljxR/86YN+8Keszpusjg2ruHpnsx5dlQq
FVOdBO290v6MHgVXZOkxDdZ4+jnIXeSaavVcZHZWd4l2fXHMN0YQshfReYGMz1VX
Vs+HPU8Q8R1leFxN1IGxrC+R0imM62mzLjho0S8Z7Yq5RRsRCmZtGs/L17w59BUV
nDoZ2dsNaf5yv80Jsjt8qA+kImMIaUylC0sMNzIkgC9+9ILnKPp+NFf10VYyST7D
eOkSQQotdv/iKstpFSrqY2Gt4uY6WOh16KVS2hnQxQe7wx9ssyfSmtaT04UQwnan
t1cSmLpwdMw1eY0v9AtfpBRXmYheQPpK2oFgIFODtMDPj1qsEloSWzVxnC82PjIM
gLZOuGFzZvXLPCH2hF4BaIiCY1Uo+vAInnflmLNv5E+raVOSTAhPX2qKG1pxj19X
4t53ik3R8zzMYmznEp1LE2Jf2iX8fo9eHY+J+urNhWnO8Oi0xQ5LBBX34gnWFhMC
qvYWErHZeTclkGGe8yrJnclBKRIBFVDxJt5GcmvdYzEj6u2ZGrKEzCdc2njhX6Me
YjjyWhem58/kFyYllQdNDe+/Oy9Ce2k0+ZLrJR/nbay3+2/yLPxfhs5PnPSbjMhF
epHVmXIYSuxbcmp3XgGqKkSdiGRPVq6psOVHtPm4QT9IAnYHaWwjZijn6ug9Y4ox
gQluYpR1brAUmk7aDnSvTIYCN+PXq01naKMt9IQ2XfHrlYRCHmxmPg8rXi6xBgTB
N5K8eD/AWNyYBQFIpHCa2ooe5fv+IBt319BWuzRWtbw4A6GbzenAFxCVnJFoMN+L
g+oRs0h4ZCTCWAtO9wRGnRdtxHbY/TsJiQe3XA7OJSvAcyaV97izfc9XbNVjf4CT
T/fD9lXw/pdk1bkbwXwTBHXPTnaxxxSRw9ffoT5brdsC6n1IE+42PjvoVG8ushgl
S4kuxFwK+aBCqvh2x/b0afrLZeUNb6S8MldcDihKZ2p1AK2gHjzzfO6HI9jfE3WS
emqOHiWJ5+ITbOAguQZ21+bpdRW+RbeMIFO7lCMa979Aou4H42wNvx2fp6PS3G4m
Ykvh5THX0KPQisvi3xkRouTO57Nyv3+Gx0sVmckcNd/CPbKsjLDsnUzMuUbd+Pht
CPaRefvdp/r0DS5pwXgvN20SiE1fL08hwgROFjxeNEHpuizpMFOJD+RnpEZXRXEw
WOSPL+KTI7Zh8U8DQFtERboQt24UpukGOKUJMbpNPAUjfdkPv8oLNBPmkcnkSrZP
+Yj04w8nPti0injlbYz/tdq86ADuBNqqbzeyW2S99riJClP0flt205aTq46MwVI1
+HGboFw4wGTnwK5yceIFLmvHFtZGA990uFIb3LfQRWNjCrKYwKlmsixphMY/ZjP0
m44zDOPszX8fqOrSdAmLGPsJt7a3mc/6w9g9sTg97FOc+6GVA3X4LSdEzTW74ve7
QuKOOQd9h1d8QQiBDJ7mreYUkv9MASOwmTTJUrLG51QBas5mbo7Lnsv6vo5eeSpP
IVdcKPlQEaXWjOq/6jZX4ukqsMKFH925hTpUTTmKKyKWet/h7nzgyCs2PSLEyLa0
1qDseNchbo9ppJzVok00SKu/BoOn57dHpA71N4KeuW6ZmRkKHtlZV2+qiFYuuRqr
9mKYziFjR0cxKXXaS617urX750pNDNwBzwUgOLsJRMvCqynsWG8SpmU3lomWDnPE
25mlem6p2vkLo1LRP59Xlm1YDWj/ZYWCMnM6ju5xDNA1CJP5f8dLyU7ClScsRnmY
xol61qnO9J1r2BClqflxU1XZmEqWiRCz2z1PRWTrE9/7/E0ONdHwtDWxBSMf5i8d
rt69+7VHXsDQkJuKRx4LajsZAV8JAKdOdURexcJM/HzmoZh/zo/x1d9cfoFxawgR
Iuv1/h7kgoRO1mz2pz82T3UMidfXasV06NZegPY0k8QsZSMHgmeM3nJGU8xURyFQ
qGwc3sGX5Kyo4opadNdPAUxp5+WCwAwdvxgLlnHuwE/Wyi9P7wpYypWoZYlCpRuM
92SoIsT9F5ViqSF85E+VkpNR1ZQ5beah9l0gD6nuAsIlUc55fOVqsAmpe0IhqgLe
uBB7ZsjT/dThV9bz7uBpWVR0sHGCkwGLGwd6ItOe/WgDqmrxFXmx1DW/u5eLNK5F
zT1aXRTST9hNqJ3HfUgHSsKA7O1DlV6DwazHOd0UicPbuPclQZo4uRnunkSgelht
EIV47YbiozC2nhcuAl77Ipf0ZwooXOsbN1yN8yP6rg6lpRm04sAL8wBabyyeIgDr
az50Xt7dgM29cIiSY1ifChkcxXcBC8lZj41nxo7rcFyKfTFFS10otkepmeXj4Xcn
47ew3QnVeX50cN5aoXuvPYGSc4B8/SZIJbZa0TbQho2PpvH+/DObRt0y4zZXD9Kd
GViFnjVmBQOwct8oOFC3yvRgfsBBxbmP6sIfJoucOztguRq8QhCJ9BYnIeQN9r3G
epLcbsxqXTACgimljBsaAgLOQz9kZGjRhfaDMi5OzX95OBJSk+NSEU3MS3S5wryv
hJ69CrVJnQBSHje/MEpVVYSvr43qbuR4gEBUICr2Ze5eM9x04Yz8SYp70vkn/LKT
s3hlKhgPoKpoU+fFWzCzrF1GPf7zSMVePokMS/ptjjOqmM6Af6FjsQbDiNbOUr7N
xpeETgjkOldf52VmSiaTMgWAt3oNAwm2gY70JuMmKh5X/C21K3BXvKhVTLksyfdB
29E1e8V4pVc40nSiqKXXR/GLYzcpHlLcSepd8bujnoQf6J0Wisl8rjS8Eba2Rleg
d0/e6cuotFjq4QpESA4KusU89x3kN6lFbdIBvim6NWgwSCUnFUuaM+fpjh2uDCAT
xkyAI7pv6G5mJAFg1cR9HzSVzJlbTqAJBT0YDcLaE5lukzypNlHjiDjdqJLylZnO
t2MQRS/UifNVYec3PTFV623rgxWKcPcgZUhG5KFIBVZP3pGa1U6eIdtXlPX6Ocko
ml9uoyne8SJSwLHzRkALO517W0P5Z1GcqFLtAeE9NqyRlhQLfWaQnU6tjPIn0MJR
ssZFzmEwoLrd591qnFdfNfnN9pF6XqyIoUo/TXEt+3/57Po2hCDCNzB0FDTR5NJE
jq2Hj+OW18fwLQazIEOvZg7cxmAyt8mGL6gW12/8EJPpHJpbxo1y/7oMBNY79aHV
9jbW0nxX2nJdaLQSSN/lIYmR3rdHQL7pFK+C8hhfLpC063S+XNf2q/+WTOQaZSEM
GvrPlFrdf7bNT5SsDlIQQKdO4lhQPERzz9mSWTEEHhgkSzH3M1CJahhkDamKAsQZ
GRFr1RW55xESzpP8BBefVHcqPDa3sX2Py8X5qDB2v2jet98tyJPqYCWDvuBDZKbR
/dHFp3XLKLPpB/RrxZsxCx2R9ASJAiE3dus1uTxbbG143ib3CLkFhNwjzyhpZBd5
mpb1RVAZ1X3v3Xqt+ikNVOp4Qdnv7UyhYbPEvAkZ9OZS1WFRsafYPanMvUhjhe7c
1F+NGnyJG03RfwNEXN7kyAWmzAUaEYCCdAShMoejBYYQt1RFntPf+FSAZJtZ4wYt
FKF7DiYB5Ht8KCRlZyH8fZ28V3kDKdOGvORd3XacDQa2VCuAETGIo0UKLpUb1DuZ
HaV01IfuS28/k1eFXKMvaX9zBDUBZDaBxAv09Ve5WAWaBy6N+H1FhV1/kpTHl51t
o0JM0VDW5Xlrmr+HWC9dONeo1PW3S6O12+byq15LgxVUb89lh5ixOCuBw7A3DjEh
DFMVMgYY+lLxso0byAtyIh54PPyRjjhKzTbh8IoWFXs9hSgja1KMNZzkCcVaLZ1B
f5L7akGc3w4hLgQ4IaVTFw==
`protect END_PROTECTED
