`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oSYXm57We6naPUN9svYLMAo1WAdl112jYQAZloYg7XPGFRSSzS2zS4ddvU7cAS84
nhmOzFIQQJ/AWC0+YgiKq7vy1ohqN0kmNWBkCKoMxafwmGEYvLqFqFNZnGhCcEdk
f5yQls5Ae3TsOcT+0Kt0hnVMOctJo1vwyd483657SbzPlJMpTSgYOMqCIMNpeh49
zQdoDU1X7Y80IX9j2gnS7ZCiCiF1TQzjlwprHI2tSnpRSEV1fH39zp6FYqlVQjEb
K+I9DO9cDdl9tx0glBjZxZaf8HVNB+L6Qw6JdxYjDbrs8ua35UyLQSVY0zSTUgWF
Bihn1bdTQSwZRLuiXVk1e60ygGa2NQexuxnfcTaiIgt70lasqRamTJKe7tZmtmei
JqVWzv2w3+kGj6tUgHCeQ1KHB2cc0ByJex0/qfnaV73Hin9LQwGvmPXHW5Xcc7EW
fskxF+u3COWAjWrRobZZhMUR/FjzYAGK5wFenrp3J/PuOotN2OZzGtVhDTa9yNO5
ISvlCdBpDmEZNyaqoSfBYyvhIrRdEZfX/6/anXHu9P5pA8damaebcVazMnxLkkfp
820BWHVYtz6yWAEqRwOD8RZW50g5DCJiKINsl7RMznOH4vUCy1TJn9QzWfNBFtMH
DTs/Yhc7Dbw0wIj5gC8OZu6cm0LFwZRYT0lkxV8H33S7ZjzqfhXdC2Sw/CvYL2zf
zJOg+mTHsNWANF0w9YeUbJum1qOADu3RqmJjH27j2UCKeDHOaU3SZcLengyjBngt
WfDB1mlnWPCiwCVrZEN0AStPjCjqPTStzjcdzYC7Teh15GKg1sXhQ2y5IM1iNZMD
SAvLo5t9wHfCee3Rmt5LXUkPZBbjy4LFMw1EHKM5fildkMaswk1/Za4+bFLT8V/5
0CUlaVa4fRkfi89Rv/rkxfJcpYM7YFR92bUXfJzL34f64RSAI9UMJJhra/NxP828
jgov41Fhf9FdfQhlLC2wM3Ic5Oyqgem7ozHn4aBm+llOlHCAZgusSqerGgUAYYJS
4YqgnVBItF/Gg/9b2i3c3VW/y9YgtkBOUilj1RxzlDSTpYAmHF+kBGGVA9hVPeZO
/A4RsbWrEl+8iSCkttB9pu9S9caoC1vEU3fiGGrdcOzBd50dWzAhYZo5xJp7IuCn
XLtihMn6g1xionm/vSbN8z+dHYJBKcOldwQYKnruk7iiw1f/q5oSEFXCfWInVPUc
LXn07tDM08gjRr11OxSWFz2zkOfIYUIzvKcYYUzJ0H2+TAkCfGmhf0Jwu3hUqJDl
fC6f5g0EGUi4a5Q7iQVvip/9ciLZqFd85IK1BZMnmuuwm63odpcsmTstpAWa5BSU
qNk76CjGRXe0tnmBc0x4OABzZr4ti/EmvTIu9zkoK+QkKIbhlBmdJw5BOSaPOOD0
dUX3DPXddJoSk385fYaGwl6z9fBOgTPAYZspbH2E7Zo3PN5NSdAqE//VvXuJ1cP3
YCb389FiqL8l4KF06GjiaOtJts0M/+hZCP3qBuuf+EOY/G8C7D98SBouNUthBRuT
RTXbVtAtCTbNQUmSBQ2noRLsJOnU65Vrr+/9hTN9rakR696Q0+neuzLidwI+kyI9
knTRChZeFoDsoy+cMfN06rcwZiPJkIAKT0jGAl98RHu0L/aumc65m36Fpk8sMY1k
8BPFUuuA16yKHsvxXmrSG4FjLZaSj9U7sUrsSJ2Av11wTAOs0TUGUIgQPo4dZjtM
kSLZD4bxl5FTFh5EzK1sqTT9S/zqs4f3Io9VIpqmSZWLbPNM2ictCcXnn5Z9bZu9
Ym47DUuxKDQpahi7cf7Qlw==
`protect END_PROTECTED
