`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
67FpW44uR2nRfNnClw5GIzaXDbJr1KO2KPcxYdpSYXneUpCwJuayOV/mAOWWSNat
fuoCRX3sa1YGBseGLe0cFW0bNn68muZz3BNvhiVypTO7kJH+RniLrvvvAqBgvnAY
WDLNBUdlJXZO5NW4B11IgVaAtuQIpfuW7rHDN2BfFZsHEEug3TtwhoBBUttym8EF
hU6+eX4Qg+vOGljMAYDgo0KCNpKyrfwR95mi+UOHLFDF7wpNEDqnd/qToDhkEViV
A+pz6B7rRnoc4fB+Jg9opRHojQZUzb2Zk8A+4qxBbnAunsXY4Rwd0/A9XRyOsAAG
XDvaDF2bCiGMcBnXvBF0Q/qPxuw2LGZnExs4j0+9S4t2f+tCuh3WwhYmmaIhAZdU
6EFmBJF4jYSCSWAdrFM6r1bVU/TGiMwNx7ndGXJwx9NQ/nnHF8TwFqFyT3BElEYk
1FxUPrSxTERFpmBQxKoWefDYI6Z5+H33/tVcydeEqX1HkYeK4kb9AiNoX1ZaNujZ
MG+zQnYxPtSc3UEiDZ+3qOnDmjZmAb/KzzfapixYArMNXIuDImWBD6ADU4haIDbR
0Fg5GHNkft+X9bXW156BC9/+3cRXaap4C0SuNptX9NYEjggU8Bo66Aw6M2Ta7909
jjhWtMHcnpzKjvQ8zUvumVEE0VBlVUJoU9Qs3pHDoS1+O8DbbETQgogclasWHrXg
enksqovsn0E4Q6sM7JR5Srv2g6ucpULQ4mpJRMU7fNmVUW2rFyf3+Hr93pPW9vU3
`protect END_PROTECTED
