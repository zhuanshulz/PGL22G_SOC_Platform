`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q4x8tiwH4EvEkwoQYtFjR9XTJ8xzmpKOnldDlOrKfIoe+18hSWsPYPz8Ci+960T2
oCTLaWavpc0+701OrNXgCcFwMYgiY7Mfx9koK5DOCmFT4cEc1pC7oaCHqNBEBNPy
dgs6IQ+6GZhjP4W3jFMkFeqnmaggv2h/yBIoukwABvlf4769uFCTls/FKLWDDwyq
RaTgja8vWLRwEiT4wOnEt+xwRd5hLOj3KBlxGe8CopB0C0jP8P4oH1cwtD7f43yc
KzLiyYV8MwgcQSbS8XxJptpuA9VfLu0jAzNGumg2uGQvRGV833Zof1gWhR6WKiQf
pmDpjWGpnmRoYSo9/lyXUIG/Ys1Vy1CguINhhfzObVRfisVwMzmKKmzoubF/tOBK
F2QrgX+WDbkf+dj07k6Emgxmh3vL3MOig4GtyHPFD7hZTYcrzUNiV7QNZQ/E2YRJ
HdnGdJqQer4tPfzoADCkBJvI8yS+V3sh1pIud0X+rF9OErcbpbn5R9yaGu9cOjE4
OqXMm3VeI82UWt1KQZZyGVq+TrQWMD6CB4ePuTlNR3Y9i2uMdBc8r2UfXejq8HAA
y9P+Mpe6jO1xdvxGU+yeiqmXwy0GdimQ1LnyPi1wDgjvZTyTKDkV7pbBTy9GIpse
AcZpRrO3g3C3NwM/hQpq6x7KuGbl3ANPeehShFPpYcXX4JvT8sBdg26Jl1U+bp5o
d9QfnS2WFMx9SSntSgTGnDNxD5hY8ZIzvF0AUQgcams2SVjLczG+A1TgttUWdGP5
57ToIDRcLzjLkZPKgIZLAy+AywtSWhrdfej1+t22QdgMyNETCjLIaIMjW1rNjVZw
DO8xEES8ruIzbbVAbaYGrdTJ5EYq0cYnZ0caw1hd4ptIaNXHPU9X0M/KGueIS+SN
Ec1F0kPDkrdnzPQq9ATrgRk9XQEXtiJB7D5c5SKT+pUw/VMEmZ8lFPSyjsVY1TWV
Jzx9aTGy0qq1ROs+H8Poj21rU1q1vJmDU2IP4abZWOsBLbZ3eWR7rm2p6jON7Z9X
VGU/X2xHLN8lW6rIE2Bohx6vpJnKPUm5c2KJqrIEuTckHe92U+/VwCv5UFg36f89
Z80yigLrMhMEmRUYoxnLLhB3YV/72kX0ihTbvJ9yvzGhmVc74OGD39RCl1W9tQkN
C0wkFiPRHYcZ+0uIfKlEhYtx887AIQFoaoIgDldyIhcVsmQLOYQEuRF5fRyhTkpv
bgUfJ/eZHZKFZSjMr+pxTSfd7V8Ca7ACF8jhKSYT7v3KRUxSDi21dO/4dpPf5B64
`protect END_PROTECTED
