`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XGeGRef0ZjraFJoFRqtxDm7U7O8Z2eICNIzP5x/dakMlAdlp2BX2IY6ZxgLe3qlf
96YSIgBF9o1PWjvRvb59RbC6OtC61Rd1vxoo43wjytak4QuQQyjNwSBleJYxVt6D
dtYfiDIr8HHpyPpBbaDMuuIKXVpTe5E6s57zMhpd7PWq/vvi02if4y7SnLICwWmU
7URMNz7VT7v6N/uOrhM9qo/6PL6P0yBJSSkD+Rded48dI4Lh+9Bc2qxb8PNFRS66
5UyVD3U9/+j+MnAPfcREl/uwoyVZyzoCaJYnBhayUgPyhqn2DgLNq3vJkt8JDvay
SH/X7f8gGGF3d624FDh57AdlHA1EDccPF3Gr+LGPNgSgCliEDY068nEIgX7K6183
C0HZkDFJZ/BL3oSdajHFSqGa15gi308xSAZvWVYxj18WQzfzGw+l2Wn0wS0eN1ZP
+kAU5Pt517FDCsyV3pGr62/ssS4PDH+leDEUrut40yf1uf0wcpiHDoAW13K6gdxW
CLuGrrvBADr6omQetS2D3wPQtC5rtEdGzXsgx4PVHDOknpzsJaWM9Namf0kBYeTy
QLwxJ/+epAsY0AWH0XrmuOeJHPxPOhwh8Fub6M7jCKw46xs7XPavY1B0+2Zg+prT
POYJ1Kwfxh71jOAc6PZrJuddvu29IeprE0Apz6F/BSEvbCoeuV1U7JOKAyvkrUYQ
+KM+/AQOoi084peKBgh1cQ3f/7csoSzIwxXFgmzcll0fks8hF6t111uhn7IYAxBx
B1OUJFfxvqRvtoxvu9IaTWaGr20OcEnfhl1y2s5OiF/hBhkzAq7XNZ7Wwqd06/zA
WT/Ri8ecBRp5wibWJyIft3uDbWdCRBoCQ7xB+RLJXTwqwIkpbIcsLPqJ9MmYCqXC
C66SU0KAFlZzxxebWm5vJUthsvbQQpbPySdpMRoGtMiygTa/kh8jtzqX94AlnqY4
O3GNvdWndNJEQiQNQ1BjvjQ+fswnx1lEhcGOTWRH/nzGcX11ittK2qypWWMp0ME3
pMulN6NPTiZOhtspv+0304Olitz3nVgwjbGfpp7zRWozWnNkzHvQ6gxEF44SyaRN
NOpA8ZTPFCCpLJNXDONl0r3tRyFyLMRe/xTJOjUk2MHsWeXzEKQI9Gy3Iw23uezd
fF+HdhQPXnmyuoUMEI4PTHm3mTvUcufBi5Dtkdy4fZSJMWzVVkCNCANyDijw4bdD
O27ICgOkRNwLI3fAGc1AWfM37h4E8uWpo2FXY6nqhzytawzdVxreU287KBYq0lA0
MnC5U0ae4etz5jccDDYDpjHNCWLlxwYMHoID/tBoOS/VeMYenjwZZXS79Ux3QfnO
9AVtJq87/uP65rcZDQgAl50tBu49P8kfRnXh3Rd1ZsPZDKjT0IAYcelPy0FFL4O8
2pCJHvJa4zsPTPcsMKdGI+JQ/trm273B5qaYjy65dkLfACg7seL/IlY7fv0wvOt9
8qrfbvOVk4cu+kg1OGlgOiRU9ygHuqeZiXv8jWoACRWc2/6b6MNPmEbHcRrrgZ/N
RgDfbxg9CYudgkff/b7w86kH/3lg7T6YYPDzvdOKOSvSPy1nAF/QxuqWuJ6f3zSP
KVITKcQ3il6bKTg/6C+BUwt1ysRo3DW2Wx2z8z4jwGF4U+IFtKkvG6gbBr7jR2/H
`protect END_PROTECTED
