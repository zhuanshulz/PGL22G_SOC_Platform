`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J0+0L3IGdW8Ah09Guwr3EaGHfPox2tbyLX6UQhUGOkD/Ia7W+1JByqXxeJDGO8Ya
2VqahAtef/ePZiJ1tgQdo0WaoV9Z8+glrgga8Ryuaoy+Vx+7re8v66748aJWN8B/
b5UkUMQSUKURLGvczrORPxUi+sgKGyxL5b87dPF/FYNoz2Py1+V1cJ9pvzcWBfFR
fDITe209uNCbrD0iwYCF2V5QdDN90oc3IPgMwMHDYDgpuO+sciNC3nF8bY5c+GZc
gPWbhDwQjy9W2VqqTkRtP/qk04oFcPMlYcgOFciT0wMfczlNmL9l+e6WmK/nOxwh
YYXAlSOyn76QKgIYsJMMvyG3Rpd2woLjnVqXseqDZnjNWAqH9ApehllLBp8Cocmo
blftEvtKAkhpjv0DhUUORm4Uoc0aaf7eC5uGUfDmbqX7uDzBTnDVq13qNBVCgdGz
bRS/z7nF5PWLvPShRoe2hE9/uSScn9cYCUjnPsJHYsgSV1li7votZ5+g4UEQ1RZw
6zODYI1VL4b7B5/P4nrFvttKIlOdd7uYEQ79eUZihzD418/U+AWriLDR+J2beLwC
98Kat0+lEj26F1irNueMza64ZozjKFDDY0rsS5RJmdKMb9sNCU9eLuCI2CrZbBnS
z14hrzkD+WAlDZKddvPCk6/7FDobmskbVKoHKIkmgJQmV8pBR94Q2p2fBR3x4GiO
Qcn9ebIxa0m89cz8f3rcSRfNMMVy2KwBpQdXoeXsiy67TjcsG0DjrZu7D+n6FERX
nQL2BBDPG5C58JPHR8AqkHDtlnpJBMJsoPLnc1asziROLjp1Q6qjRFDyZRCikGOE
CZXqzlsDRrWsFmBt/tz2CYRoCfRARedToi78n7AiR0UaUaSbL/x4YtahOD60fynI
UBZSfXD6BJLkkzX9ASwEJDqebqYnYvrMeaF3T7etc8dgZpRyU5oKwMFsK7xzI+3C
WtK2PA+GtnozCTcYShyWzQVcw6lJyu5A5iomNQeNk8k=
`protect END_PROTECTED
