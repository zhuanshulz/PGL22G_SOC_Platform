`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XEifErRtVlS1Ts6WApIlyUe2nx90y1u//xUDYMqTKKBnVbaBxSiFY7wvO+RBi1w3
d4sYLfEfqMdZaadAVKYv4z76Zb9h7H5pEwPiYi5grH9mbuAXNShJaRaBIWKnxvS0
Q16rKhsxpoKpmvovToNj24sUfbl5WETi8mfYD8V4WPjowvIF8u72g7kdMvE/KleL
LAMG2NLXOkrrCHzv00S2mQm1WFJLaOsBBFPZJoAOhYmdJ5gAgRJ522zX8vUEGJeX
iHAFtadFtyKTrdEXy/MEL2UO52WrNGrT1UjhokZl1FQnoCpZ38o1s1fPaxnVXmmU
E+hIUbqmT/owb1uB6busEQZishfXOYUmnMtQ9VWqlv2kSJKHk3LEk4Fe0nW6Uxql
Y/PSDJljlZyY0BiuwbMUtmMbHjJGSOS/R+D384GIbjjXOalCwgXSWYyyFzXJTFzf
J4iVSYx184SpeVil0sK8vfAb7s4RImPt1MWH7Ikcy2/SorQ3pq5UIr9CMQY9dYNs
lLW1QjEP7YQ7XXzfn9rqNBxWRNauNwEW4nSvD2cbmel6WwOnFz2TjH09g5hBbdsH
ztKtUtACfebiaKR7zDaPcUsVJABjDSFO9bWT1CAtJVINGxWt1IDlyeUMMrtz98XU
MNnmVzpVLdCTXel9gOQBcsF0OQL3+QqZ6/WRYcFaw1n16fRAfiBIDu7iksf0x5mG
CtE3vevAtjRgJlbCnAcnH/4BMIsvbDCr2CI2xIJFGgdJhrhmM6dTFlHmKM6H4TrN
pV2yiA+PX0N2gleKLf3pZdZq/ujmB/TWc8o70Rd+PsF5G110Cp0gaSW8vXB2sqz1
OR4yFmaXdVLeDfkO1CIc0A==
`protect END_PROTECTED
