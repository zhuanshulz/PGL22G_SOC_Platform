`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2QdUXCZRjgMnLdTeYgSh7LyZ7xIG5u5Fn+wNfWxJtxJSFDlG9JOwy1hIf0G7ycrL
wgNCzBlsKk4Vdrl8QSe+n40YnvS2XgqFV+eAb9zJqfSVbgEYT7S5EcsRvfN4xXgN
kLZW83Hr2aHluh47/7OL9KNsZ5e/m+Z8qlC9mpzilplTAQ1w2M5iIe2369RCOsLt
/2Ig6v0W3TJYxtmjKEEExrYxk5d7dikjzLuISSsSUtc18T+b0nu+X/uJzKPPycn9
ViqNaq0+uSewie8oYwuhl2il4jl1KYlEsK8/MO2KEdY0wHA5vRCks/GFg9wYgTAs
tiw3muv7g+RODwd8vkCA2zpEGpNCaeUEuSJJplXkdzS9WjtxQYqto/PgwinId4bW
Q2BmnZ9R1KM+4bfR3JrP9rkfndIWo4eN0Mx+Q3VkDK2yaZXgoy7ZHWXyDPRq6K11
t06XlPuqFlaLiLmDn/9+QNj7eGtpFH1qQ5i4m5dF1flH0FS0iOPwwdT5kVOgAdIv
oUBeHsStoUB/hoZ85Nlh1gXVkjCEFlyOXMOSdxJDEFyZ3brVnxyxQHkeY1liR29l
`protect END_PROTECTED
