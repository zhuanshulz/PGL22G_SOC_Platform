`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5euoBnTaBjWn+exaKXygcCnyNcPW9KzAMxl/3ixKvPTqQy5YTBieHcTrUpdS8znp
J7481r1iREbNadRD/uNwqx1859ub66uF0mTxAx5fNzn3EOZ2DTC8nb22PMO+Py5t
jdDMfGJsAXpZoYOj1lLFIk4ch2KFm8REPEfyrIb3n/FprZqb4oiPfRSlT0cYo57q
kotkSpSNtF4uBMoXjWVl54FiZaVwkCkj2SXtIO28xhhBVnCUQaoVVNIXHyPDQwOV
GQq0zKLiMsWFx3ROerStdhqVjwQaApGr2ytVIOg7Ngg91/tT/1C1xzDHSgtRK7s6
vJlvVVjxbTraFgdaNbRgTeLmIiWd+kt0GRUUVo8D8T5LmD/jYYssOFjicOjA5Ill
ZXxTUDFlkfsLSd0+0x0dPiq9yOECUpjSRj1Yll5svObXgvYgJtQvukeXUZgG7mtl
MHSMw85XyaNULXVtS5r15S44pm95rENJPlE/4xUPzgV+xXymXhK183Jr364ykg48
DHNy+KcElrH6NiJe/pJ0ztu+4wrFZ6U0ePf6f4/lxgdiqLcN60nlvn1kVWok8TQk
BVeZ2eMvn5ANuPZvz4tmjsrh2k2r/3tPIvf0HF4c96eMQ3zC0NfpGCqGMYe74Md9
wFDJ1RQjYh8ibZ8GSfAjx4xNRZhI/+yIck2aP9lRK+eGYZbGV8wTS+cKHJZR6wRX
BdGlLcv3pmyruO5Tb31+I+DkU4xbL9UrSDN4cv6NSdg765/sdnVYiGx53ULZ2RXK
rt7Ny7pXnZwA9cmvCAPWKmiXxL3+tcd22IqxCs8E6ElE90sajknfYxs18IqapmnD
6Af+J+7qh+5Ttm4eQv9ZROz5WsKdLwgpiUuqftVaGATluway0tuCZ/41liJNe3dQ
Qzmkxw4zShdS/5w6GDaTrbLjkWJxh2WkGdR8ApkROxR0JZfGU1afSG/Vxewpt07V
uVjq7fTcMaMVnLTEL5JoMjNu8RohhM+yQJcRY2W0IUWLTtPiPHaD5QAQxQXmZcDr
gL+VyMRvRFFj69by+731KcfAQJyasQsBopAkCQJmOlkvt4v/aAPhiRs6yRsVhiVU
+Juw1WEQ+6zSPL57BOJHioIQwngj8foM2KBzIpr0Kc9P66k33YDGlVHLAiY/8ob4
wYtXQR2vfnuiOONTiBYT5qgHNBROPNyS4itsdCR1n3LNhHB9/mMXpLneYSfSgUDu
hX0RnB/v62tEwqKC50oF6WY2qjJMIa4gAGYI3KkcGgomMTYfQ/RF7S4y8ZrrXEkv
J9hpTKnGTe1unSyFm9HEPbD1tfyfDqsBGIvWB9xDFhae06c22mmMVuXM0a9uMDkj
dOkaiJYvKglvFsHPqlpg65cX4w44wm1LD621WgvplUbNkmeaq9qKUY3AauETPeU7
Xqy9Ek9ttuRQDNZ8Um+IVw1uBvD58jtqDuaOp7W4/MnlS45SsUkNziPMm+WOftYX
DkPR4MzZY1SXtCPCNWzTDSpI52uFcch9yhggdNnodWMxj6DF8KbCOMG650H4xS5W
4ac/W8JBOrbyTGT+lFkZX/0uHtW68wIfdj1vvB6hrPOCqgErJFAwbaj0lw2Cj2r4
eABtgHrJulIcZfaP1+UHiXXxToVcGwGaADFluLrhzZxdLq5fVPXEOCXNcri9l1cD
6aIxzaeywZ1I7gvH4I/shtziA2rkpdj6fikwLv4SPIDX6ISdxbzsNGBreWtIQ2UN
dhNCpz85iiyUCdZGO5j9aEl80638AnESZZyOnOlkYxBlf/cL75xReWQMV3hTfMIN
LpL9nU1weOuXeWRsfR9zgn/CiO+KFtqiVEKKcah/OQPGExYwb9xrwgFwNKSQc8q4
2kiPdaO3weictZRQ7v3aSuXeulULSXJAKxeaO+15PdLCPiMdIeRIHRMMrqd9pe2o
COlOu5dsJHjBy43mNLdqV4h2I3V+BueATBD6Ad60YQpfAFWrG/JMQ/SdSPqT5GUI
BKORaCJFPDKxwFK3M9/6AokRbyCxMU1sq/XjUOYUJg9qgHE48zI583vvW3XlCuFY
SxzFg45fOm7dZcA5vPA9/g==
`protect END_PROTECTED
