`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AWuYmEWqLGAC5d61FXPTreEoqGB+bg4Gi+TuxjOkI5Pq1LHXukHoL6xErIbs4ZEX
DPfjrKI/7w5m0fQ465uyZWTplJBMDWKzN6zLMG0aodHwR9hFEVhgZizwOBp9K80T
ogDh60IVK154IY7GYadHBHxOP4h4YexE09sXPmi8YQux+xfUkT/PIBYRdKAKroJL
36tAFUgcqcVdZgGRHdEZ9QLIYazP+zbfcwBHFc+EnxkZpOj+B3hhdLpv4FojREmK
VclpXO8Znlbpa17B0dfBGqWPc+8Bd/FnhaTXYyH6/E6jfFgOeGDo9a+oYKb9d+6X
KytO1bvTSD6c3EhsP5mi34NDbVKK8AosYfX3H758/NyFIgTlEZ9b05QgzoDrpC/0
j2YLgBEC6Pr6aukjMTHFvOja57YvtZawCkP1RPXo1S+SdZuktGCD3RcWSG58Bz5z
pCtzSONAeXOlglCBnNzjDjZzGfvuclUCTshSkhxDvf8LosCRkq6ghBe+6EwXzJDY
dquU2g34VsRJV5wkVG8aTT3ryCEwypabbXzTEeK/DbGYmQapkEERldzO2dTeo+F2
J7/PSMEdRJRVOCFkVlJGvBMexLsy5ajnQULK4U0F2tXIlEMxy82h8p9Pw9MnithA
gcEjsua84XluzFkE3zEV2yZkn9FVqqo21QHsPY51Fo2K/tV++FG2hrJfMf+rxf+2
90fzyN3rV1kx8mXB5pWKbO9FztqkyVVAlB+VRh0YU1Mik3as4Q0CgfFtT6575lIU
BXUIS8odjJqFr/obZgSkb4il8TTp79XFEvJCbtUdJbSBVvfuptBVx1zeeRX0e+Mx
SVVpEnRKlW3h0427gD5eGlwinSWT6j3doqgKHqHsihTQ5zrDdVHBiqeOQeTeoW0U
cGyhq0DPGDZ69QgziPoZPrAyaR6B0V9oR/qEbTJqeOy4ZlPifvr3Oiw5kTCKcshi
8YQmW6FnYkipXhJIq0g+hxOo0YISBGKMmtNO1QL0ytNxbMbIWdgiug3f464oxipN
uTHSv00L2hFYHXW40ffvNg1CH99SrPmUtFS4wTWKLbeVDQCIGxc7Bo+NTcdPX67j
FskVwitBctnhlluBIqI1zOXtVNAc1Iw39peEL/iL5lcrFa3a/fFG7fx+zVOYeGoS
n/hArSh9WieIfvsW7kYtgzH33E/bWMsAWiV1dabmD9/5oRWlC63QtNjtKOt3FIm4
lGES4ZUu3nXDo52ycayeLRrC9hRLbiN4bn0txFdDo/vifE1nuM+kGOave8RrEryA
rA59ajnlbnhagUReUtb8hIwsFFfgH/YQAL7NZ9E09vxNYQzqqBB5XvYRQVnhqfnH
pQunRuPY5JbPoSthXm1D4o3dpK2POqsUEacjbHJrEsV6SLSWuzgPbvBMdCZrbH23
C1jHuUed1JVmf3YOgOIPOBhATacbp/aQosdMPzJJrEqcqeTQNxscC55Rj6TeNBhV
Z04XOcMMci1wjbaVQhXIHTlm7ayXf5ep4zAsBEG/ntlZLUHQnpizZrQRjFd62PS1
PA9OhW8n7ufL/QDhHyzbm7BM2UMHPp0wx2HGIhgckn5LPIqBVhyTr7AUKLzbg3X3
8zYXsfzShNPZqTzxAU1EzBY6Ou0f2+y8vLzzNSWn1GHtERSHr0eOIG1vpD4v0LI0
MRpjAKzuH1zeq7iVnkFSIdjdAyjQaaftdgBr0SRiSgfxz0wwCp/aUDMSb3uggcCM
/G4/kSZRKJki8jhyU0izpvRB+1ovEUpZQchAsIayGjxpbwf864AzVVFMIpt7uOZe
CK58DFZkNojH5KMrbx0Y6FStOmfxxJHm5K9hm4E9guPNxfGHlXyghPdOjbA40upN
SNKRT/7WtRiQO4eDfIa9t8y+lKCpZGeF2xxEtIk7p6td2zCtn4Xot4+asZOL/QkV
pYeVF8xm0Q/Vc+ZrMZhO8m6wENDYBIUvrI8cW5PM/Cr2cGAAABAOaxPjm9qxcmzx
PfZXXHBrPW+Mdy9neQrYbsgRWg27xbh+IV+vaHNdq5djVp1l39AA14hY9NRNE6lc
yHRqVSDFM1omMw00qbsPM1TrqPL/R+1YpvqfUUVguOyI9KDTrldVCUMadGBETsUd
rAB7GKBG/7fD36JQn2PtWu0I/EG74ReQbPcvv7gIRBvkR9rHvQACZ7uZ1r51KMNO
KbcU1kG2u5mBnD7Vmnbn72Su7LreSVzG67J3OFSf07fia71d8mRO0UGPP1n3IICo
1CKe/xRjFBfHY9PfhnAKmX2YZDpbDzdcuLIdS34yO1dHsE39/IX/W278SoAd4iEK
wIdWI6R2xQtl3T+IMYTKNJnkr5tMnNoTIHaOFX2pGH0y2PKWlgDzeNNmuN6FgC65
OCu82XM7BGi6HYh2XnQm903w6VYhL40JLDOCUmkezM40f4Q2MruZgFtOnyXjXkY5
NIcUrvyzcUoT680U1jSo6qNINo8cY2AkR/DfEhDcwpsQqBoENk0hGP2CTtFpOseX
SOkGpvhUsTS/UnvRrJh/WdachQOYtbnuKv5q6FXH4WTjfTVdqVHcY4LHMxTonr7V
F4g5pViA4CGf2UsaLIinOlUnz/b8HdtPfXTfnTQYwBw9baZCFveqOVktlHx9HFaM
QuBqyYcb4zkeJ1vJYicy/ECQK+JVDmHbQtGVeQ/h9ni7+TvKkit5D/qXjaHGRZn4
nEkjUQElSBSUCzPhB5FIV7vXv8WOMlSkBs/UNLKGdX28q6FmrG7oE/6RFaoi8kQb
cfxSEDZMKM+HELlKZEIXTLZux+KtAiK3sSgRLISs1g98UPV4cgrRjtlAKESmit9Z
k7YYHCZXeLN1frG8NSV6WLCYEqn5zg4T2qW36oLrUn1fIzBkyOwMmM4uCtxJ2kwo
37TsukKTO7thQzxwo10FS4Bladuei0/OIT9pF5j3LiaS6/kDHiC9T14VkaE8squz
NcSw6vPTi5AJ1fgvWgQ7mEJNfuKMLcVkTXQGVlvMoZO4aoXMf64Za6ZJTcOsfxaO
4Usq5LiKg3ayEWsG4gtTL8QBVYhsBlF48LEyzkkWoelJ8oGXk6PGmFFEb2dAjr8y
mcL8LeAfEip7c6RaNijdDwXbTrcKvPLJ5M4LQpeEAIX1sFek6XssaykAyHZtCj8y
VwKHubIRnfOkYOeXyP8khFJfDwSSrv8D3ZXoPWKi5mO+9YOaGpfgZprDVfJLh/Yr
o1eyddwxfjyh3+wRcny/Rutbok6frc6tm9q8aiZuPQKC5SxM/84xSXZb+GWk3bqo
llZ/glNFkYr+UOIAQ7WWXNki+TtdsHFpEpSpyjin4/EmYF9ertWiXGOTjk+1po/G
9RcDIbvRM9CfAkp/rn+h7oxl2k/WLqXkqUZqUXXSOraevmy+TS8M1l/5yPMzjpCM
L54AexXC/3yoXcSV+DZjafYkEbwWyRlaSo5YAUNSLAUZqyq1vLmhdXh7fUWKDWXr
wo6DjZ7K6iPvRYBn7vsph9GepQ6ah98VYCimagpGOQwfkDFSXujhvSJM+s4kZe8Q
Xnrj9rGC45H6dUgcmLmdSU+wtKphY+JRODlwVLsTcDPsfGDirHe9HW6qQnDuPkXB
pop+43YSgUMwKX+Nmg3QqmijBHk4efAg0RROzaylZqm6MD4OLjRwIe7HhygJV5Qa
ysy1K9IwfNE1rDsvx+SwfLVoRzNSAwcSpxaJ3C5JaTnY3kTTI0mQfXNtdbbow0PQ
SixItho6rifYBoujGaMdIOn7KBvRnXbhYezQ3a0I0qRTux9BXNqHEGIqt+z4MEer
k80DW+uUhw0Mcx83kpkteI5/zMp2x2y+t11d6gvjYoNmg2Db8cALzfx7YNh1Ug4l
kZnrD5nqE1cB3SQhyUgVCPevNTmI+20wT7pEPEkpToSJ+5PDLgR0wHqMIGy6v62i
SBErtTR2JcDMC2LcJWS2/N/CnlKQKdOUyti6Moi6/5PRVG9u6ha7uHJefghNU/01
UsFGVG8QOEsAojA7m9gMnemUPxkZ4HAiroE3KsobMmgaRlBRjQfd8GA7MHC8u5KF
wXq37V5Xpuk+b6QhoUi6vLvE6TnxYBhR54y4aq7J/FdSagHvPEo02aDwIJjLbNNN
riH2DqXu6Kc+VMXt8EYchBQns6Lhk+Rf00Fz8qqC2DTCfQvYtHqzb8dvG0kE9DXm
irUVUtcSdMKItFz+jexARMFvwK8gaoXh+zRFAzDy734DFpZDBMYomOTALdDtXk8e
5y6GgJ63Wm1Hx7NQKEwlU0zVWiAWkr+cGIEjqyMOnoVsHj/y6UloZw5Iuu/P+Q2I
DUBWZTTh7qmw9CbU1DaEQscPEzPu4H0OzMENfxWbGNBLawZm3hVPJOy/JjXYIZ3j
v5VEGFO+70Iy7GaAb2DiD+O04xJD/em3TedXd4WGxaLmVYMJorqUuNZrXMpkQhZD
U4OMv0KWFTmFarm/TIIhwL4WWuH7be/ae7Q5x7d6//mkuv7gm8zP+/KR6+lHesot
f2TqrCBM9huODs1rkgXuR/O4aLgZUJRejKxslCQry7o8JPVEykbZalZy44D6LEjt
/VvFSEMYdiOe+Pyz1+DxaUER9fO4Xegl84/7MyLI7IbSjLRLiv+L0IzGvBGRrzU4
E/uQYT+7kqHuZ6YuNOltmcsfvo8kB9iSKJbvhWVBQa+Q1cI9jIgEyvj1tcfJm7nG
qs4ubOq0ryRbXuODZMRtDPxwLWBNj3O2A42mCVHg16SmI/FRYIN86lfii9tZgA9U
jfeAdr/93cG+Y6AWKSKffx5DeXb2AmKVwWBOaDPyfIVjKfOtP1vnqNUKswj1CXBV
gqyPktBaSUoYSWAKfbE1tTVrFFWi6nKaSRK/HMduKxkEVb4NRihd6U54HGhJAGVJ
iZ2P8gNauljxXs1ixhyHbngLoPdA2033J0NeKdZiIsRYhpfZwIBgSZfB/+9gR461
RnUBFgDVOAh7xbINqvytaKF5Pjmjc4hGe1Tp6ZmLUIR6myLq2lHJ3Y5JHzLfeKBh
7mJNk/ZZqd6ZfdKHCboE73U76Wcldv0Hap4EgYZT22uFFd0BI1oERsJq8S//7HZU
HzEILNhGlvZ3Yj0q9mmCD2HZSZDaEUMu/Gg5oOj5RuhOt4exyHcONxfJjXEH/9yi
cf99KcEFH5rAMq5AuljXNgeHfL8tZm7Zes4b9usYpka5ncx5dXEJELgqXdX9kGfQ
spwsl1BQty+XMOJLlI9WvK0NHH/uNNx8f6sWLCVjfIVu3gCTFqqvx5o+4Ae5aa9g
9TnepuqWOA+3NhAcoBxJTT9Uz1jWYTfO0HTLNbET94aYgl/sjGIbdzT1FgsRbtkz
X4A/XfS95wfyaq4fxSvoIro3Lk5me2U0JrjKOmD9KlEH2UK/SJ5k/axaq4HNf65k
Hq9cN7FFQes3xNJ29iFkqqz+QkHpP0ySuIvmNmeufu81rTl5anfD7/qffIHh4u8F
fobT5ItZyRbUKfbDcLpBrJCsEiaOwLWshwAuVxqrbgGl8pIamybIW4s8bUKWmkKW
PIOY+0NWlC4aIHf2es6TSCxldCge859st7U14Q3GlfyrvRps502py5v65pTPHUam
0eDoz23H/vOrDai2ETwouVf0whwGuLawa5bdAZTirNkWZQSIzsR6A1WnJnSHwYEG
YQExx1ktrB2GxWVbChY0wOZhJ5Swua1ryqi8Ibph7nZRRDrxFVF1xaH8nYQb/dDa
95Uag8OTFAvNK/NfxRjIbtd/xMtdT7uMcWlT9knr+VRfEUQ20rOgvk+LakLDDzWx
mU7a2NScBPhWzG5idst9jlmt/7uHeL5cfWJI9A1an2M4gvnhdUApm/QHpJybNUzW
PX6L+3RC3m010M9QIvZS+TmjCENnRp+q9oFZlCCtYx3oQ+rUccJHbN9a0EUuzmB9
saOOaFCbcaaRp1g6zEDddRwTV8vSxuj1uykqS/Hipe6zT77WDYkStK5Gx0ymaSEr
mhJHcjmm4hNZUXGl4snRJtmRoxNbUgDJ7ic3ZJmRY0Jr6hSNoMFj/2W4N39YVFws
TDxzvrPxAzFakM53c8ZS86M6Z48stnbIfyXDPa3K2DE+syrBVun40qraUGNSwlRx
i907ZCtPTc3ur8A7pnYJljkp+6POLBreGZyNyrut6zQQRbjXFSxyVqcW/BYSHavp
NIgPGUbFhoyXNh0UK+kDNPJ4VT06Yjs9N4tDFkKvf0y4tZActggUVVhQmKR2tYcD
psaXvEQnoa4hYsHejHuTVM7S8O6O1sNoBadwCops42mGg5ALFesb6ESMfMcFRzqd
uXFWFfSKyBZY+HBvh3/1anV0uPdhGp+YD2/i+Dz2Q4iepEd0O0D/l1ul6jK3sLZm
s4iJCijMliPBjV2AXptBJRHpeb3hmBs+vks3OxPNGuloHldvQ0z/xAdc+CUM/yBW
+s/gSKhALEnJHKH+9aFrzNkkApYwGbAzGxakkgD/YDTm3iYInSMjnXRErIAnYukE
KESl+NzmUV/CADmsNhi/csZA21MXKcbkrutRCUO1JPJ9OWpRnuS5qmnhhdTMFvgc
D5TKzvzshuZoOGfFl5EOkZdwR/qj0QbPWY41NfcVr1rD74gdSUdqZ9hgU5Fxufda
02dDXGQMFe//tK+NvUtYJZUFxfHmb9/3GYQuFmTEQiqdj9sbHQJ7VZcamPHdxSzT
dT8YVRwLZNb33KdHmgYCk4WlKrFJv/MUOKSJ6d/r0t7h/JfwQETLHfku7Rgdw6KU
ypGlhm/ZHibcBADMVv/s/9UBDVUIIMfofgFp9XgQ4J4bSjdkxLOetKGsVusuStFT
3WMQpOblyPJzt6hPQUQ+lE1HtotUS4KD+Zx2JoOuCr4enWQteFmciGW7YqyFbtGX
vWrbl5T04fiiBgUfLxTSZMjCcNTftZ9wGqT+pK/2BNBZwi4M0bCsQ/muGK7FN0fq
I8B5WJdBdVkqJyTxt1UHVIASP1BqSkv+J9XDPGPWiBDyaps9gkCcL1p3SNheEndN
+FZvLpbkxSnW9YhtP7wVlt3RWpw60Soj3nhoXcJ8DmiqJhzOjux5VxZBNFxqkkAQ
AGjYeepwhIAmaIwW6RgLZMp9eK+uVvQneL/0ungZB0xckUoR9ejyBd49uCvBXFVk
cwzcWB6ZUONgsiHD9WIMy17j2fzLRVE69qCr6VuUcfsT23TwlD+ihshOdl+CPdmp
T5JK7Ik3EpV3Y06uuMeIx0Y2wLNSok1UwmaKMvyaHX0Jy4KK4RneRvTjneR3HxAt
92Kso1p0tqxsVbUX0OY3zJco+srOvU3E+Mj4bztn2Z3civkuf2ZCNEqf8aaOg5hd
GvkiP+lwQp2TpI4c7IrBCcRgbKkm52ECb0vfa8MS7jGHxpF0pk53rZ922TzwiZ7d
zX3m7fr1jPHV7VHLRradqBNS0NaHH+Ypq4WRobH5JXUUY3DyYTg5R0cvOi3vYQtq
htc+rUjHQwmY8u+LRhBtUld0rgjpmrS4rqLzzTmYJV6PEY2AXAecfDMlvQXz/rWj
77f5cqHDTWcZj4jcUzKlLFd6WQd2EVmOgANZw/A4mKsxibId+LQ6CxdHCXN3chLX
zVSbhdP4vyUhmrBfreVB5YClIwGLZexjwblfWLtmBVtl0J8fv8cbizVOptMh2iPo
AMlTEfzqJPm5yVL6fIZBcXF543o/lCX5qDxhFLz8vAoMVRcd4+TR2nRkjJbhXSpQ
E5mbeiFEUZzolSFYFxki8DyAzNbzBDWKtAKezg+nGlb2xpat+3ZEdobXwM98X2xU
vftQkLUBOG0/fWNcvv/KA22+X3VrK31zizNWfWe5RQ1gxzU8SKINkv2X5YWciZZ2
uLnUJEgBuqMahhLRX7EXwBfpkxpgIZAqOYfqC47qI1MsJivEW1GJR2/YFf1qcrOA
Kq0BKp/SQ+gt+t1sovZyW3wxE7ITKJJewVeSfV4ZPa2Lh1lHK6aAu7zyFnFUGvs2
vs5rjXbjsjzSEhxvD5r519wZcjY3KnHi72KZnrQyg2mVlwM6tyRj9+brFO4NEWHT
cVzTJFAZxZ9FFn+eUg07NLEhqj01Zx6iWq43LUED03xi6MnvNIwLzUMwPgDhoVdG
n/yWERKr4D3LR9cjhvb9fnj5bnXEbfXj4PbXAU8YW0no7TCS1Uol8/qvy2nEbdmF
pfgBdjkJQ5PryVQIRNf39EK1eKjE5R7Q7vVRPSCcpX4jMFg0KH8O9/nlruwnBiY/
Msspk5eyeQZbwIXma0H/iFpauB+MavO8WaAD9Z6UDW+0mMz3dzuxZ01koHnGW6Oj
hPti9YL4zeB76CL7Nm0DC4Lvg10zj8gEGWWLhdUxaOfEysd6CdcA7M3QPdGwlucY
Cio8732vK0ajTZKLpUlzlx27JeXSmxoJ0WbcsN0jTmJhdcrh0N46wnAI4LmXzzRa
`protect END_PROTECTED
