`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zjSZGzZ/7qV+x1JLZ1pISW+1LS5Ef/1h3szQMGEDmeahlM8X9R/nyNCQGKcec1V0
dBhuRuuoO9vpjmHNvO2sOUpQSDIVME3Php36qv2uSXAJEw3ToeW8Xty4TXgVuNLH
Si+u1F6u6Z0ofxdSSRkvsrnv73/gN0WagBThLOjhxDB1xAD2UZdicOsArcBVcZqb
aU9rTURgdYFoczoj9Z3UqqcJVPHnSW4spCklL62NfxsUI5V7zcl8bT+EJxawZYbU
Q8OMVQNmgxbkxyIg18RqeKZHZnSk54a0X9p+yspPg6NgUgZ7YkbvGVDrVpD5Bi/+
5/lRNuyIwtsXu+Qqgn/c20Vi3RrApx0f7DGFVUk21oDoCuaL9KgNeN7cMKdnp4y1
4+oHxKO18s9x5JH+/gcopErP18b66p2vauXEI4TaS8WcUQBdJrr/tb1Q5PJRyptI
YhYHgH6rTTcmhMQc6d/zwHkH6Hk29ldIUu/meefQzT1tHdTMoBZTztM1UTC/DmKf
UDQZGOuBy3hQzKMIgppripD2cLi3wgojdds8fQs/IH2A0qW2sOX2Xfrg5aur2may
8fumfn7fM33QB5fP1lZ7weZ+hfclc/xD80ZZucK/KhNnPC4nRHgZq6BNAZRficjM
N+ayAPRE6z1WChlSw1Hq2ZNlSoQ9NlNQl/j8NadnBZKmOq+D/0xbpyYtWJEPsfHN
+1zUnC2+eALOAoFz3WgsZl7KU4ouIfqP3zO9iZxjVpCX9KZrmnGp1b/kzDRTzkJp
jEIdI7T965nBMD/wjPJjEKowHwfiXql1g0/yPRm/O3PWrKJ6WH4FZOwD/ikBJ4lG
107CiQsTfSSte2JMqpKj9UAlL03DULyNkfETZGn4muIKNcWp7YB46eg9OsfUICza
PC5i7PDQ2NXB9yAx14jr3kfyYaVt2mX5UzGPaBWEiMmq5JvHiZwf1P+2NLqN8rRF
NQoOi+/hntMc4Vh2uaMtsZosyOTY9OTQiykyAnhF6yfAs5/P1PWDvOXZRWT30PRM
GBTaQAVd0xYGtHtBHeLynrXBviwnXojcAQ6AdCAcYS9OhT0e8wGD/q1o/V7j7rPw
/m3Lzi7CbaXLh08fnejC4/F0hxvAvmyH222upFPAy+nTMFHoAgHGSHodsdfZBf5W
`protect END_PROTECTED
