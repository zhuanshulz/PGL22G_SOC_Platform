`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EdU+disomzaeCTHsXMkvUbPA+vqgS7kjTVoUB6m6wZxphTrkOTqWNSZxfpSdBXxs
x10y0pke07XjS7B4GOBthEFFjr62j5AtTNNyVDUWf+dRtqSapK/IncJGn8n5B69h
iUDD/Y1Y1Gab27SlBhLQXyxRVeqI7nyxmzCny2WRTedOQTGiHnkEKuJoT3rFJcOu
PmUkOcUnga22wnoB9rwShi0VYplCGZsP6oC69Beod5MDO8uK+BUPBNRu6DddNrdH
ZoOhcwQOfamQ6OmAn+/Qkzt1NfoIoYuSZOPiHaL1quNoNJqiym/Nt3L9OIZEojh6
ECv7nSKN0lkYJUCQvI3ltFDGkuJn36FMLhvbJ636x/VlAmiPVivEh/rVzbgv1d0T
7a0syRzUwER5IDAEugmnnVg6/mgFrhr89wL1E/tvJlFsSwAKmMIWbHYYM6KL96S2
G94fvVBnqpryIIQ/NPhq71hLPS+GA8LIQ9U1SawwQUz5gk6bDLw4crK6e/Bc39dh
XZQK6Ku6S8lbHh6jiqBZD6+pIgfCYW0fojqweH5zAbLfrtL9CU28qrtUeSZmM6Ct
GGZjyT0cCb9lG7Xsk3lDPRDQjzj+/ebk7UyilpXFvu+gdOThFqLIfeYmg/bNwWgx
TdWNdAdsZpv/dddnhYhzhWoGWIp7q3wzJmvbv7fLus59lukNeqZjUWv4BH7VEd81
N/EntV6yyFGNIK0dTXum5iuXI8EfimVFgRYU+G6aLKcIznsIXlx2ySy4fhrakaPM
BiOxdGpeGT20Y9auZaHq4ov8eZ8ThpcVuevWiSjPl/3giJjgPmYH3ReDVhTfX88U
5zIzAurcmU29fOUSycxFQ07fe3bDzmkPISyaMAShhIoOr3cvr9Xe7bywObepPmAt
nesPVD1kLn0fNKMMVS7kL+tnAOJiKSfntVv1sa5vA1UEDMl/secCYQ7DtHGaPg2L
P6YxIMCEDSG9WlCpOvo1MA==
`protect END_PROTECTED
