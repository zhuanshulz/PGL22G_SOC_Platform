`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jee05LErlZZaTxU4SaimZiPiAD4WqYARiFnoc/+Ay18x2ciGfIVh1GKutXh2zy6V
0tkNfpmZj/yb1LljuQYPCJw/93PagPFEaekt+Kx4FLw8X6idrUlYc/aXT3MUhZmz
uuEgy0IKcGG1dueaEcSw+3GWCzBWAzTDCm4nypr1e42dBGn4AJbXa4tA85Cx5OjA
LK+8RIeXQ8Cu0w1/HrOqlzvUOjuzl4UNTfvD01V7RnJGRJiRDea3ybsOtNQ2cePw
QedPJMS9ju0EZPgPjWJhaaNbCTgEObmVEwBsky7h3FEGrrNjcK15UuCe4ZFTo2ZB
Urz853unSPdyGHYf3bpSzRYfb0pje/rt7OK2y3WN6rV/q5RAOZDle12WstZwKZp1
Sk2cpZ5BXpNmxjHkdT76za3ORIoE8pG0bjKjSgoUeq1lYfetVfkAXk4k/ohKzhSU
39tlCnlMoTAtTx0g0dPJAvVw7YwG1s31oiEGfVUNh1E5hJ1jg0aEfGpePVy+WqTA
8i7ifJ+HhYIlImEcaLYeYXPhc/0wbnfHeq+z+gREhkQmVWQGEdD1bAS/cnVR7zRM
paNgl75JjH/EhDs6cgZTA0/GMY7U0x5fpRjSwlJSRJpPnppfbKtzRvAm+E6YGXXR
w2WZSTKClkhXtuWFytGoqo4lrjajGcsMpoJShdoFbbAZ0taAYUiQqPMc5S5pf1zK
BgsB8U5LYSaXe903HKVYVsOX7GkNvBw55g2Q7t5Al6RDsEvlY6iksn1Ui9BBfoUl
eZgmS79vWvi6At+evaTjEZdV5CzIN3jNcpndSoUf19b1yL+r06OgJ3eZgjke6O9U
jT57pKQYP0q2ai+G88+AHVsrEFbEMV8CtiZlfyGO0Qf47Of/lC6av1eNxjtGmcFf
HR9oYaNuR/zmltBN8R2uebUfuWPjkIDJMo9mUJjVzB5dGRy+rpVoh+xnFDP6vrVa
JFDHdeiXFT6t36LZlYf27KM+jIfw4zvrOMdg41vJotHcdsI5eF1JP8EWpD/LGqBD
Q4GQ0QyJ2iFKWWj1jDo0XCu0IT2K3c89nR36w56IYL1AbX0kRYwenTSNO6TIor1N
QCS4pP3flBPHpnn+C5pxwfj2Dkrb4P6RkzlvsIuTRVOWPenJIcdztT3+9FpJr5Mx
ILvnWH9ZCOSNd1MDuuKmCqLbBxMp5mLt85dNNrpAB3alCjw8z3Xcl9cKLZqybQLU
hoCCykWrn2psajkPNV7CzA==
`protect END_PROTECTED
