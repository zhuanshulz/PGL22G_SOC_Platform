`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KWmC0MNu6aPvwbAWKwl2e0vNvik3Pea13INlGAJeAjqBa1r8q+TuJS7f01OacQQ0
5ZgKUaaP2WwG5N8/UoKJD0iMTVKGH0FSoWeL7+yIZlG3vsnolzlJv4QFyR5jy5Oe
XX1NtLlztbRoc+Zi1YqIxugEq/OoOc0VSCRSvAdo5GyXSwKA+oTilDv/ABWNYQr6
DuNNqqwvfyc/A/qrhh6pCpl1rRWmKS+zzKdKf1sZLWjT0SoM+Y6BhcQnktrMxEFb
MM6akqDb2GbQjfo3gBrmBaRaoTDnpW5pYvFjvK99kMN24uF3dJYZxqh19okgZ5nZ
1467nrwEXHr7+1GYGUm01HvIwtvWeJGkKlyW4/eO8Gi8r53NcQqdyS40Du+CRyXP
jy5wxeq18+YUW9/IbkciEg==
`protect END_PROTECTED
