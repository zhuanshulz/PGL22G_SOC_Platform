`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
doIcFMkjQch6J9S78QpByn7TSfPSU3EYq4ZuCnSPNQK1KvWGhjtSc7IzLXH0HFt6
UXSxoJiQDO5RVrOOyqm1cGStgyDBSMOQOV+0rZtsz+raa1+JzEnKBedUaei06PxB
YH76WzBU13qY7ARZxW3uIIAiPHj/jPQKW/4TiTK16HR7jqSNJanOMZS76uWffWeu
U6XLIHIsYT/SsuIeM3TlFu6vnsCX4X7IY6odhmSvJIIG/e7m+VyuAJZkj1U5LxWH
zHK2/Yg8mARB+t2/aCYJMWeArHrpuv82/nxr5i/zHZkxiPk4G1mFJDx8s4EjikMt
1Xy0inQxFkxlitSXBbgxTMkw3Ghr5//OWmGa3xOTc5nX0GMgeU+PcYme+sH7thRz
3D2QcS7KIwLgeKxAKtFkDVYK1i3wROfiTmZcKioZSaG6h/XM91uju+IX6gZdLbMC
0Wz8nAOEkEXgbF7lUk6Aq4PtLlj2xp+aI93o+NUFgAo=
`protect END_PROTECTED
