`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jAs7wv7jtDQLk20COG9aN1PJuaRbOx30ua9jKePrDSlmWyvUvdb3WwFnbDmR64Fh
u8V2igJ6ResEIAkJvWhHDngaZW6mP82+ktj6LWUCusXZTf4EoKuQ0IO7yGw3C2cC
alb9Lo1UEx7YlKwfd1AbfcyzzBV2p1exEZM9rqEzQZPB8CBzNm+iN5bG3ITvNsyH
QdRRIqn1kCto/7kaCyywTzfxaaBPF2beSYwzHBwsZmuwZieVLYBzMiThHGCGpebl
Kexir7+7C2FY4AZqZeZfc2UtwPiQRmYHrdsDdz6V0ycyPnCfZbiqgG55LFmJ8FOi
Wuqo4pkqsVd4HhZG9gSWAxHDyJVssNpn4Bl3eMm9K6GE6SiJ5gIVnUccMA/anDj0
zflW12OjcdXazQpMIrCTbJjesO86rQxqD0i4nwiUnlFV1CyCrqzs0tVhmvBr/wwL
2a6xt7+q3H2FctwUSDdBwdys4UcTU2CIYhYIlTc2hr4dFda//fiOlUwT71t6POYp
t95U/eqU5GiNVSqynLhgNOtFvD1XY56rLRTn4yb18T7wtrwd/XdXwElElKgC2kHP
NvnQKu2pr1bJATAei6kbP3dFCQCatyxDqez3T8i5PB+xUGo8xjGqbrxmN4ampzP6
T7eqFbChSaADzOZrYBtOhScxyW1+YCj5/rGJFlB2hqDHNT+5wLpc492uGYimIYN9
AH/VW2QTUAKDcFfMf5HRuxupxrRjAAUUfH11f11T5L6Tp9ufDMFmiQ3TkT+XTO8b
/5QITrKHQXW+/OE+PKA4CswjEyNBbTgAMIS4Z1SbqyrsG0UmwD6vM/B8FWUw4aok
aIuv1QIzSDTbE5MARXjwdGA4GN5nRpiEv7n8Ts9KIDCftOucoiFwh8ccw3VJz5Dq
Z9qfXW5Saib7GRy5u1UbuzrwL1SQ9U9LL8UYn7wjqIHTHB5VTpfJtx9iSDAb9pv5
Hq2f8Pp8l3S6okagPqGCmom1hFHrK0AKdDMDjHZFXQQ7O3So0RRhMcQ+STk3gTbt
FUhfStwsdyyZRY8TQc3l1GF81zKTMXjCfx3s279scoB2++PPUY0oEJGXdk1QHuGD
ZXYzx9MwXYNrHfFl15Ept9inO1/aixQj5RXPTyqZzdRqK61zOv4R3piQWP5A1jl0
kBN26cdkeFOOypPwrmRjfEvLOE6Gjb9FPS7Q/K6Q0sHjtRUZzYSv4Gb9r0eMhBio
CcLKIGWAEfPSq6Aptp8ddHcLGB+JBsl14aYuvuVW/kYHzZYyQ9NMREeyfiGJ2jhn
02SdF3eMxVbzLkMvZnpGASThMU9+F0jKQvTfJR1BKDFHDeLrF4CElBQbqgZtNcqB
8x7lk9/w0HTM0wjzkXr+aPbV0o1vmhKQFzTPND9Nn1FpHCf34EmBTLKVE7moEkaH
YWYiJLq5W2gRxbum0ecI5btk+czVyup5j2i0U/xn/sPK6OzqKLnPSkj9AWgAF9Fq
+ZT47P7WF0YvOpL4UOmfq5uAEfL9RvOaF4XEBvEY3i7ZWvPcsZWCV9A2Opqah4T7
MfJF2H5c8f1AFUfemzeuurJUIHRHst2yQ1elqRT4j4yZeo3KuK2okv5Is92NZGgJ
FocjKf2j/Q2OP5nTKGAdH/n+DiTwNAKcp4qI80/YVeEmDQp2ZXUx+/WfkATSMKgO
xPgmmWqXu4/Pvj7+Im5iUF+CX1Fdu+zMted3TNRNfMDO5mux3WRm1q8k9tO/Q8s2
KjWlzDUwYQfOeA5HkvMEY8t+I2E1IH3iiuBTYYWCwcuuhcennepiITVbFEHTx+zM
SkvXPp5NOpHMd0SqJvIR0xguuwolOd+c5z9jtkUAoEavaDkK/6vsJWewveXSstls
woezSbFJYr7C/O/3cSl5ncDIU/K5/lKU27vas0CSbEBZiDnlHTnQk3VOC+gCsQzD
XsyQES1Qjzj76vQqXJ9nolFAVEfqc3vvSd0fy/yN8S7s2NPk/8E27c/RSy6RuQgO
AX7uvVPorQC5RgCBspoajpEaNttJ6DXimiKbuhrmjij/hQxQzJrO1WLcHuszQDCw
KF2HsBjqS8bxSKMDJO6FFGag/nRBixp/qePMVTlCjOc/DowRNa0ONmvgMWn1M72k
POB28e+pEi1PeIcMBpcJfcHih0dLK2Ht5K4/YAjJsLEeaUc4cqfTxwWqMLR0oGSy
tsH6flcpjPI8gN5yewrPOJh0LFyzdTCpScX6SQw5lc4utRe3S7g8xj78j8VSRcYj
+PVWUkYRM9orCvsy59sKwYRrUFDxDM1tWPW9kV9zmLFgMQ1i0C8bDfrYxAU6+DfC
7p/0eE+XiLuxdY3M2ZYJv5Fsbc10WF9HpDANP8jO9AtRfvuoqFepapM/oMUnpoi+
Vnu4HkC52yk8Fpydrr+7rKIwBXDh57Fodv9U2uA1jAILpupSTBT0NXHRfVRbWqFU
fwm6T6c7g8V+g+hYdMzTmGLWhxDOVNmshkpncOp2osjCTTuMFsar8/D1bWOjo1q1
e+5ekJNCHb5VKZVbfmfNq0TGjW9VGyqun+ftU0d9raPPDPWXbDzCUYRYX2Yiudop
i4K/yzaNiZ2Wbgq2ISeN6aW0VkEWfo4WlS0htPB/Xc2Yo3JAZ0HG6ou4LPJOy4C1
6ypxMCa3OD2YAZjp2mUKvFeWUTtNTn34/dXbnE6a0ZAr0XyjKqrWbBIAtGG9YbI4
2c2Hp660KYZ1gIt7rR/FEfr2KyZDZAZg1MB2GZZIruey8HiUxOgyqjnS2RmGnMOW
e/bH5ZP9mNLg0zc40cm1JYO5WldZs3QMoHHF//oiRqorYbrIWChGa90hUOeWVXr8
LdFEU+GcCNq2WhK/uL5DH3IfGCbDRsZtAHYgiYauIP+HrWGk2nYqwaQGYZnBV8hu
ucVLyHAlw26sH6o7BoLTDAEK7fZthq1lOwLkOChzTtzqibF47DfNw70GIxkFqx8r
Df7OJpjWctgFkoNG8GZCnyua8b9rh8+ybTvP+c1DvCv7DnK3pnkRLW+UpwMYp+DX
GOnhqkR7kWL/X81192DH+5rAYALkndc9Swgd2TB936odE//akw6aZAVMTXYYuOf5
Z+k+tExR7dWtOMFsHLPbQOdMrmk8dgQYo2hFSyKdDJnwwYyCIT6UfOS88MxWPlVL
mbKEL36wKdEiRgNgyAVMochupWpw8sXx2Cu/iKTFCNSaYmFWlMIikshzgnQGAWK1
kzGOgcx6n4uvLRF70e7D/p+Vu9a7LI7Md1v08YSTmLLsgd/zlX9Y8/kkaVBB1ORo
NwiF+FP9fSu6bmKvN/mbcsuwA3Gq9DZ94ywjy14x8WfDYcfMTP1EUFhP7wdkUHS2
/lbY35XMr+WzuxySrRZMGVqUybdBU4VqU2qt1Kl5gBbYvdGaezeA3EbnbfthGSvt
E5LfqL2nXNQgOwRWZnwu3Lpp2+hv22EBGEfO3wCqLbAANumOqMfj/34CYVrU0scf
IElKg7b5uihEO1Kr+8yUFlQBzSURte1KVprz7BJC7TKnOEcqtJNGKs8I21OeSCAr
Ww8fAccrk+3OOmEPgqHr9jGDyaOy72OqK2YOG/9xRIdYcUBPyKeXrXlPfhz7sOCK
NLbcgCzkdv9wqqm+xN+f7OzVa1DQl1/1hns/cEtMWq8RNjdzl0RsTTv8pE/KtVf+
hVZ93KyNmQnM5aVgirCDVcG4oJofVC8GahN6T2uQCGBYz7UwmMChNmU9Ytu9nHlD
XsTzrIqyIuKmM7Ay8yOIdfTU4+wWc/+HNGHqbVJ2OzHjeNSUvgIgrFDxz9/gH27T
B/BgvbRXWisDy8Sx1m9B2x19Q8nU+G/7r4j7v8bD1SiApENbWedsSs47NPDkrQoe
NMQMbMEU7aeUBLuU5aygLMeXwqr0clHatBgYVEIyIegy6WVkOJJIbAdWBY/lE03m
ctpoDJUBIHmgvCw7Z/1/nsMK4ITxOKCKd9CJtPFiwWZ1FYDyrq96nRXs05jjcJdb
26rHmRraIA930NOEEj0w+Bl6cO35HAQAWsuogCBN4uk45I94ioj9PE+MURAdkEno
JNgPcpUOvVqm2H5GqtMRWs3aCzYVfn5lAn0/7DoQ+k+13+NFWgT92SYRsGhk8FiZ
/NzDDIuR5oBrAHY27+4M4P/st/ruxAHqI28jsje7NY3EMN3SJ+LqvEZgY/z/b9EJ
/8WXpv7ps7SGTAiZ9SHaU3wZeChUNebCt0T++mslwv3Bov0EigNNZW+H0c6gl2DD
5u0Tn3PwYGyQqx7YDEYS0j1tn4WrWTF0gqKbc0aCxOCum7116oRT/bRL7hdiD7tC
11CjTQVJDNnm427unxdXRVVVZ0PVIHAEtioelbqYf1TA4b7N9rZoffOE4S6e0Zdy
/hZUiptsKkhX9+f0VfSoU6Eajiu2oRALjVS0ApIRnnLyGXq+TkVxnvZglTAdCtc0
b9WK/dJGUQGdpnLBlAX1pVOrMTICLED1++4gkkAmpnSjZCa+9bK2H34IHqZCRYqL
dLtF6Ls5DsDiRQ42yO/cMTEO+aF+kPVzFu+xZCgmyy0C1ITU1wgt1aLoDAC4LuBs
fusFnHxFrZdVo1KQ7cciEaUwyEKSThdroMjasGA5jeQnygXEb/nV46ucivfWufGA
p1oguj/NAQd/fILJ+sNFccpozvUHt/rOVLUmZ0tKkWou0JlgxXAxpFJxrhdxS3Ot
Lfml6wwJ2gkKJfQUhoMMl3h5laZJFRHhXHHC7MYaNsQbsZqzB5RK3WwAXXsQY4cL
`protect END_PROTECTED
