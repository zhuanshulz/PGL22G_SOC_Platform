`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aNlxtN4xF4G4CSh+P1lOWIyvDHZySgBqnjqtQvRhJ3dkN/iU4t+POxfmTsO/8+T1
oeli2Vu6C/n8ChucLCSWbMZfE/2ySygfGDSqpI/7X1GslFVwuPtgxPKLq8gSiAq4
fvUpUMFX1uh5psNpI1oDL8aQbrKg3YIh1Rw8+4BYWAyszpBOhfzaJ5Lnkkx/dxNT
06nNvEr0fjUqe2ILB/tA9LxHHy0XbxneLmh79J5Jb/JpPk7Xm6Wj3KhZG8gnrWhu
6RDbp6xtr+RRO/uXpn96TylDvH0c30uM2eo8fQjqBDMdRK0mqKwS7WdvwRbsoGZc
ANk/OSl0O0rjqCZEJNYjdFyxV7PjJLtZ+xo/wl2LXBl4elHBgrC9EnhlAiKPclg+
5uZ+9/DcfXD32hUCAopa0+LE+jfTxuDn9Hka74Hfg4PQ1w/rP9XSXM5EbXPIu6Iw
DBurGb3LofHLtUyjG2pkOLYJ6CQ/JWb5pnnxcoEh9A4cDZnOQTLhnTGQZ/7WiEsk
BGe5Jgq9oarUJ+zfRwcmpgINgLLPuvrmiGkDd/ToX2Ig3OOFMc9QaUe1M8GcLx6i
5GZzml0k280n1ZdgBreOGtPsJVsVDO7isGSRglugbRqxqYOfFl5jibFSf85xSE1T
ycFoiQ8/BE2IQyot+h/Q4pPNGz0saMiYsRAgIcl2GnQlIZAUnD/VqyQXLpt4Q0w4
MAfKUrHkBzDA49fi7EzerIl5y7Z2B9TDXcf0kHBjN7vu63fI1JYpDxHrRyoRb0xD
9jKPqDKSkVukchDzcHj7VcJLu8OySa/gBFvDYL8FxAG33PDgBMefmXeg75WTKYsP
Eafe2ouznDF5Cu1sz2t+o9bfc/l6MvMoYuvj7kwElBs=
`protect END_PROTECTED
