`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eRdxpr7M2TDYomShgyIve1J+u2jjO0qrOLcx7fwPRMylAbK9H27B2AO3cQYrr1Gk
auBtUqdxezOd8wgx4SqhTyhkQNFXTIf4wSYTELeykfj16/i6RPqmMEEBzz3uD52U
pPT/6TUoJQKnaTv4WAPU3MafFHJvJzD+sBRap6vVWKNNgNG2kmvelU2+apBeYfGt
yt7ETYBm6h2cxmwc8hWUERaej3rltqD0Y0AVx4WcfAi9m7U3wnMoXdd9FGG2GlVH
uxZgAfSg19kCQFUAfEndTfa13R44R2NQMNRmW1Dg7vseRelSC8sgLOoXGOtAMTcs
bEw2b/QEX8kDkgT22+ugWxAE74MlE1gTch3zWvZZ0Qw=
`protect END_PROTECTED
