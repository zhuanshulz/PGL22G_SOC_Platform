`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0VLGS6zpSAOWgqrWSaXOMsgZQ+pZfCT4T/jLqV7wVgOjpujUh7NFPrVi6nWu821I
toejRcVnMSSXqwSlvZMFvtcf/3VFKQRyybvmLv6b8jk5lmgqwW6G+lq/mJ5VzHUo
fi2ZcOK8hZShVOMOEz1/ybE5F24fUh7IupEoaG73pnz1IIlqgDJFys897YdHQPbS
NAFVuzp8AmD6YqYdMYn2XzuFXQIb7B0M7eAO04HFdSeYDfwiAE5IRb/696qAYZ5N
VLazxs1xOzkUeT7vnNNp/mpg3Xmuhe9yW3V1gOpsK1isnKL7hhSssaIm2eiw3AEx
iMGJzq4FJiwexFEdckygIdtM2MV7hiR3AttG3byE0wzqFR3kzVXRF+Ik1TqcHi/1
GVAhZ6p0BtUns6D3+MeWPwIKODykHainYcQPANCHF9KHngFscrhauAgRKbUbiIII
+W2wjjejrngHFmntCK3mBDAH1HCCEwGXGdHb3YnY+HRhHhGhh4V18mOgfChE2b9D
4554R8tJtUjROf0ZLzJR5ZLAsf2at1trpuG750ozzgueBv9ezUhMb5vNCH+7rCZP
2hmo3VqgwvfTnCZygd3B2LwFdG0n3LBJVAlSExxdRLkDShDJHnIhKd1gDhxHAHxm
+JzYGayS3upZRpP5IJQc1aNvWMVGZl61z76HT+dqZfQry+/AHHgdF/rLVtU2wPHc
rSvTmx57lKzt4Rp2cvIazL8dIsd7FK85Emt7dzuipZ+UNoMr4eYZnBbsQEVbUM2S
WlyQ6P0bAKlpUDF1fnXUR7e8+z6UY+IedZhhrmwxpgimWgIKIG2fbnv284knyZFO
73/Rozex6eK2lw08pb2oEpqMirV+H7rwtHu+bfgyBgqPM4R7bVDUrgUQiQnnyH1a
tKAtziG57Gdr4pi5HMQJzI8/4jHNYg95dgTwuB96iNsfbpkIHrT3m/G+OAEKexs1
hdjD+JwCV4nb/luDD4PztfQ98yFhfeDuF3PJeYOf7It93NC9ADdKM+16TC0kWFdk
keyo/hIwGbNz9vQXEOw3BuDsjmd4HtAGrY9KWMoeoNlbSBesVbUyqAHoLTm4dVmJ
NLJRtBdwiwhY5OcRucFLcIseptJt4NcPs9n1teZXHie3cy1oUYqCk6tcTM0DMOaK
J+zdBXLOUD8yUCLs7asTnNpIf9n/Z0bR9YrDg31Z6298en5Sv+FTyfmBEho9yRP/
YrHlaNP7bHU3i/As8nCZLA5xnG8SNBRImPrkkJab4duliLD7biON95ZX37NKNN8h
b8Lfh04OXgw/lEMKTF+I1Ro535o/S1e03s38ebJOfNETiiTrIQvydExjLOrV25d1
iVyyyFG2tz2gOabWPIpYU2yD0wjlmvE9v///PO7lAiuMlwkV1eVuX1VOBqMQhgs4
Zm0Ko6MUwq/mYFl96OoSG+fRj9TsQJnBA/s36kpL9L1NgSAOverTvoHXnUO5u862
MDcaDlpSBME98nIQEADlmNDX1X6iGGnEwHZCF84kROen/d5zLKp32q2c4FYTNwaU
uIdpKDLJVEnxUVdt/b477kyug8bPNVtP/ORlS9ivOvCfGgGtW9Zoz3977ercOuzr
vANgMg4dxGWmY+TpBCK64BliNhKsyCgL+GRr5gfYYG/x6n4hB6FeJKSIjWYQdw85
UoPkU0a1oF5JLwovEHPEwGOgRgSMKPdKWJcGQvEaulIFlDHvwFcWAylbTzjFCe+E
wk3IgYtLU5Vn0/ogFwnNiWObiyDJ6HhvQfZFvgSXkYRw5+14zyRwCN5tkNWLuHG7
zHdgD+2IqEpYvv5kBSB5D5pojKvJ7vUqFOrPIkJhUGSgjCthIOxF+1/tzXD5Yjx+
2MHfnm7QQicSeX0mgvZSsDKwEN1i/Rshz/NRC411zqX3yddiPxwWutCAZcUEYVFj
tME9NjhexdAncS8p0vf3EtZDY52dVnAOT3MN63CO5yWbUDf5N/C4s6fyoNCgDoaA
IxgkKpy5bi938Hj0S9FtOvHKdxAffFU7rCmKnxHwZKRUdf1OahixLmlZeJmg2snj
+j+zU+mIdEdewK9JqKDyzo/NaEegaZBBhUETv5U/3JemD927Xaj0+oXZxAhdOjFF
PzK2KLzvFeZT3ufsar4p0kng8UiAtR80wK4xaHSztcruzi3vFeDtEFBZEKJsTslt
G9ZOuIalmWf6uacVMw24AV2xtYZIdW0/h64eCXN1AVlEGFCJutOrctYiqPRUxTtL
Sj/pzibB9uNAXYKVX15IrEsxtOecxHT4sC50GbGgBXQ=
`protect END_PROTECTED
