`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qFhWvjAX7MHc2X1NhTBvYnX29MjYvNIdn30JPeuTlO2YCdzHqa8M55Qx2sbAkCnV
skLRB0I+4W1zuPSBO9bPKK4PRxrXrSuF4Yw+OfGjIZedm+KKg7nDm+dIZYt5DQ3n
5RorMEwdwete6w1AKFYOwrApoLpfv3iBzLmDQMCSa7XX3A3q8opVQDhcLjYfAKA6
FdUaory+XWN6mfPgBOE5aJNAl8DjVMS/a0d3NrVMcINrOoUptf5tFdAuuCz3Ymt/
KwwjO1Bum75gh14Y2a4tu2lGsCOOhUk0ZyGNT2dWmiOFbLO44a7A9RH0OexzkGUp
p/9t6td7ybREf/nArfaWLMt6oEqHxL2dd05b0qa59b4/Tf1PmUajbgleT1V5eKD8
udkawr9ksN3Z9A5sBg//+rNDQJLVV1cgTtwqz3MGRek2F1PLH9Xuitoq7d16+W4a
76/vkAlE6ppE5yxSq8ZC4DSxkShjZFGF86sfQIF6ce9nOsoA2Y3e15kgW36btbdl
NyHE6uS58BJjqLjuFX/uextFv3Eb6LzUIP17iW2LdkmBU5qscXF3QfeUc9X+qH9u
W5vsVzDZdNIQwaKCRMIHgwfiLPBBG0vhhD7D6IJpQ1J3bUkGrIHjmwjgq2XEUrXW
LaneR9U9cR4J8VO22VUZ+8OYx6+ZDfZmwJvV7eJCMIPlxv7DgK6lPeRGnSO6pdOY
8RFDaXV+EOR9guPtLqDjsj41a/QpZB/1RiFTzgMHW2IGTYcKA3BCyNlMpaS7R4K2
5l4g8InShKX+Vqhz2TGRww2bBAAMDQ+GDynzL1sWx/dro7MOtgfI++FYNGE9T1hU
Dh5M7uNvtf8dsbPzbKviSCT52Q2zb6gQu/XDaPwvb87PZGfjqSiV/mgYR86gSeSk
X575Eeos3hsvog9/RpW46hl5aTyUUL9D7PmYrndHukqHjyYCQDE1a0TF7E0csk8R
D4kVk7djHid6pBWSTy9vh03vI4t8cnS3rUCbLadtV5CSGvedM6ay3Lq0Im/QFiSY
4PdskbUlt0mYpqUYXDUE051ni6E7NaDgTc3JlG9di8BBVYTayFqJ6GU7kqyEIXVW
uprnAOUPslu5UIpMpLG3grj2maXKULk9TbBkOAZJBklkpiA3d3I7JRxF/vNxA0r2
S2FaNLHJ+5V94/UBch8mtw==
`protect END_PROTECTED
