`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FbQ5mkmmf9kA1nghkocpXNBMZZLP5dwXm3DTREeaPnnuA05biSBJJx8Jw+Wjowja
xExpHh+71SlRzN8JeXmwcFi+tep1NMpnoRcM+0ncL7ctadpNEQuSi8ENyqji4afN
SefDMLwTXC1CbFbPLWmRLkTKY0iYujFLcZnxko0riVzYxQrK6ARL65JaGykQk2WM
E0C0t6c8Fba3croA4zcRWefc5CSuXh/Fg55MBopGxEsaoid/IHeEOsg+ZlmHjYWH
DJa5IDEp9Cb2TQy0tuL7zMQtdeFR1fjuNNlcYnt99UM8twQ3rSxMqYwUuJ1IXQe8
xXA16OHJNydZHnKqbvMyn7o0CEYXl8s/hquyLVmmJrhYFaFgkJ2p9I+F+WFv/AOo
PjaByNh/5aHaTVc1sM3KT7hmT+DTAwrkgJF9pvqxEeyGHzuRI0rMewH6c6rLV7j9
56fLutGMxGywXZ9d5E2gh3HZLCHX5lX34JCjAJN7HMXk2qkosfhrDKk8KzthMezb
o+PRkI2LFzGfJiE4iEpKz9zPS2Sxli1j4zulDbD+zWKqj9iUkrPR0QobkVOaLHum
WKJzVHZMkkAKzN2TsmFdt+8a4AfeCk376yEMdvze2w724WFLb8SJVW3/loijBQZu
XBFZU7yATXmFKwC3KZav5aHIF8ZAT2ZdSEpZJJCGWWpfEEdjL+oDYEbZ2Grgqsaf
3gHfV26IevNujui1at0z16DPU9Ush2V3pT7oTY2afupFs9EhKcBN6kYE+01l1C8R
eGg2Yv8XL8r+GpXdqrb5caXoX4d6NHgVy7Gsmmx17VHzl/zIOUFwxz0IfrFsWy0B
yrF63qTh0zBmD5TXHLDo61QTQYGUYNHOpkOrdP55ryHlOD6Kkt4fbDh+KS3jEJq4
xWFYQ1hkv4P1+pP9HHsCD4Q7YTHwaYhcqlfUvAFJ9glg5NMxQ/JMT/LUXb+9mNfU
4FPtfaYtxHmQFv0GxAShXfMSuuOhVdNsnz3hJFKaRf8Q27jH6osjDT4VtLxOGj6t
oFJka+TbLhZwHf9CkRflWVl9TQ3Ut2ZaNFD6U23cVU6YjLePV/2oBmJopakFoJco
rBWhRWVuq7lc1taACF9voY1i8lCyKJmB/Q3+c+H3DYkNyMTCLv1OTXNJc1Mbju2r
OnIktGXsjsaF49zC20iOKbsnpG/sAT2apKHK0em1Bk2Lzz10UCyqJut8PpRJQenm
VJjHhunPMw0mnkG8R1H+D0q9cWlclG7sch1Q27PscuFiuOzwU077k6pX3r/xBUfn
VoJ4GjjFQpcvQJTsWoDxu0h2Kk9CQ70d009vivUzunQT+Nux6bOLsEqlAKUfx7yF
3q2cIvQp5WkEurq1uk8x0ku89wWYcq0ZZG9ovT9+AxrciBt28X6GW/3kfyMU/Bhj
OIPiSwJKLpm9vQBLr3cZsijkBLraRYX0NESzmQlutS0qcoivRcDsriC3nycTyiQd
Qu3hXS0VO7KPWg/yDtF/lK8Vwa79KNO3ivRJrsr7BHB3t3CaDbs/kF6vBElpTxM3
nosXV/2TFle37ViWL/JuPWX8ymEu14VNU89z8fq+MLXJMnR6PpX9F+9srDxvrCV/
r5nfB0hWbRbZro5qgaYvkPSXd7ttAF4idWjwfQGLHsEKM794fgdCoVsdG/k1PExT
88YY4Bb+Lvs0fBXANBCBudwxQQSWpW9Ev82O9UsBnyXFyfmopS1SBD4YgbBptxgu
zZ3CseVjpCqy+aqe9b9q6MRhHmbsPQi3oTbRDWxnvKHCHqYXokjXyrs1A2VYRMYa
ZMmWqI4DkdEkYv28XkoLh5+GEWElcYfmjpJ6Le8shQsdiKuCqDT4XpBFQhvujhzU
Mx6rRGgYkHGAfGegMYc6gtuJd9ahcRWyUKNC16fjx/IijEJ1v3wd0tFnf4B3PSAm
8W39PIZQa+yP03MunVeEtxRb/5cYdEMNIZk7bXuVQmZ4oiwDLjp7MCCC7dOf+nFN
0VE0BPItbWWiH7OpxtDp61jXmmxUC06ZbYnTvZPmxKiV6tvbTiZt5KqDvhKUlvGQ
KU9XslkIvKHs2u1P1e7amUIMSuPGdhbWnkpIkOaFZmThs5NdiNoWd7dEKD0eRYPp
1iOChxaIzmHaPbaS8zEhVx4hCrAED9lFiiS18LMlY+E/Xc4eoq6uRmEvPWKnaftF
azGNQHGcLkDYT+ZtuFghbpS/4BgbPhi6aS4+voagRN02oeCYYnFh8JcxnMM6GrNG
xxOFJOFlEqX8X4gtTC40r+gJiWcFewyaSmWjOEa7OL/Vr60m8qkAuRaZZtlA+5nA
vh6BddJIVXc8YSaL4U5Vxr3rHxU0/2NiLvKavxEaZ0XRYLsye52CtDRDnMJgzeHY
AcaNXVVTkRUxp+X3C5NgaMUPJI6DVsB58O8saw5gybT6UkLOj9olimaINoM9p5Ha
bEyIy8EmdwUG20/4DDQhVQJ+87CRyIT/IebRvICjaSPnIsmxtVuAYQYOmOTDSzcQ
pA1RJcUqvpZ41grKkX4WhM9t0qtPBYC56w9OzUgaFbUVxJCvAAcXAt+koiverxdp
odVhZ3W8wWMaY+h/LwP8t2Bdjx9X0Iw4YeP67DHTeMeSVOR5yVQL72DqH9JwTuTA
0fzsrCJQm7M3+SIh1yIlNCxCFToZuiqKug2dnX36wwNsoItQbTEoaYxc+wuHPB7v
vB8d5Y9uMS8oh/HgI1iNbzP8kgY20otJU0DBTSlElYch3AVA1DTK0FDHJw9/ePC8
qiYdYl4l+KrRFehIYswJo3PBCf/cPem46uCZ+GNZ/4yPrWoU4mWr0hb1N/T9Ykym
v4QhNJsiq8WJZDPweiwmDrAo9aLx57TCSmGd+jz5bBfP1c1ljKOYXeZjIQf20HFe
B/fUcvyXY6fNuvIfaPNJPIiFdw2xAES53Rj73GDLB2ySpwMXp8yaR90VFVgYVdTA
Nnj1TLn0tWq8jgFDpegkfpcilnv+m2m1Y+8+M8eF6aUzYyLqbDbF0eS22ZIJSjgL
bmbCJ0YQDdogy5kNXHgTNGLX7BkEnTmuerSBky6BGcywO1aECHsQ5cON/MMOZnll
Tm8z0lXHxiAJ604KtCz+8IVZrYrWCrkoSEZgptUNpFCu/GlA43DXfyJF6HT9YaiB
S4TU9RV1b5Fw/kXEb/FXCMld2+C3Sva0SHZlyCnWKqyY1RsRsiFQYiKaplp+7czm
Ic90xX1PU24ovGRWahoTRkkckhvl03rzEX7bMAvTFOGKVnfxEAyxSw0IILgAdAnz
BRhty+qPNi+hpew265uXJwBh6hsV5JJANq+0JO7F+8T6BJIgg1ltyF2L25MoASQr
ssMaoA2cggVyhOqACvNI4uH5RZey8RhziBF37QB/5JVhUraouf/rbkyOadpTqbW8
nqwcoxxUPnPPbAgwYCWaVbT1lgIzjffR0tj0bs54bUf9jk44Pzk/65P/1ajro3NV
TcFpQelEhPXcV63CiTRbb2lqPAQzI/OnRn/bUIxBTufCRzE6UPske+9VrU2HvZJH
fTAkSO+EM8IlcY+IY0LP5mKKk/zMfkQh5KDNUSD6UAPhnlyWMCCtRTPX571nJYh2
OVLsA99VZvgIuDRg/BOzd7mn26YqXUrkcQEFQXyYRY/wHZss+REBqWvMkg1h+Ns8
3KemjMQ4TFxFbQmp7mJqm7zg46qtAQnj/1aR0H6cqltOm9DQueJARWm2t9KDcm9N
TfY29AY2+bjIBk4lR4Lvz3+tHHwLCgRvZDPSHlGsDXhXBd1NDZtmUSBKyWAgSFd5
DAQ3q7f8/eB7lJl06tWBxUO59bA4xbdAYqxt/sKDAL2s9jbvgZr6NyfBFOsoypZz
k9oAlU1mIMSQkDLayx0yuLOxtNkw65GVM8ZTO4nP7HrT5Cmd8o/Fbgrnwsuv/zY5
Dzj0Z3QtO27qK63Whu1yfx9IOaBeJsSnAJNLd64gf7827LMai5/4rRhEQZzPFqOI
+HywYAz1SaKSY4F4VOfClgb/G7YeMmkZSgbpZpxnEOAIhXBy/NiK7x/W3FTl0EFp
JtlUC0jQXXNE8CdEpa0CfkA3mJyj4188A8uFGWaY58+vF4ww4oLLSzxblpwuH6/k
TnNBqTN2lg6lOXM0FyUZUPqc6qfRJP8qqs+OU7c0n3PlIxtce8iBSj5T0XHrnYUi
FZJUO6GLS/ku01eejgkj1oZY/tHSpn0fyPxxi4Y6lHyw+f2cX1TOWd8wClr8iIoD
sYc+60epnrsx6Uga/GGcIWaFpqrStJyesRnjDkG2YkDyhUftwItpWst8fjZvnlKy
Z9xaayVw2iGewIV7M3GVfDOfo98Q7Spinl8xOqfINRnRUbmFAFKZOJqHMJUwhGO8
WmbS+3HkNzUpHWqg4gU8zE/zGcPBPj5y1DJzKwVMvpnutM1GfePou7vse3VEOfe/
PrpJA57dw9IxQy/kk57lMulcdEKMwp2WXkLKRAjL9UTgvLHn0BQZPQvh3xUW4m/0
A1y02wF8xwppXWC89N5wHcpyUQ/PbPUA+6iRsEWGrH4pqzQa6rAAuTD5rxVdV5c6
R8btf75QsnBKbPU9FdpLKq+vDpnMUR1eIHVjokKH1lZ51RGpDoirlcPdKRPuAfQR
/rgjLstp764aKQToVx/Bx+Peop5vwxSNWYjT4X6ZUjIcVwlkJdtUqjfNHIknUkrR
wPX7hVzq6cRjWYLaog3MXxeZjZ2aKXYqmlC9K/HbD8FtHYEzwBJC7Pa5HriY6FzM
cXKMq4I/uEsTAcrS3UsrPubPX8CUtOg+YSEgL+AzDyMd1AgrkgYatGGo6oqvtKhs
tmLXqJXSVA96urMkt7pMfsLRbX/g2Y4KFNivvHjYJ7MwG3mu7Up444A5w/uDMJox
qwI1I/byA/+2dd2GLfo8qM00MN2b0rBUoPLUHxTuLkKJGPvC9Xo3CF+ums3+xyiL
wmaw8KPAA78ll+VNR99GVW9g1RxCLCC/sTloemdxj4idmn2NCplTgXKlHr6CGbzh
wBZjIDFsdmzme+z/DLaTUGzPVLitXD0q3cRQK5kXwEopM++fVrreC4Dnrn+uoEDU
nAO7bR8mp1i5uzPmBHKgABrNvR10Yw5IPOX10Up4q6NKmBzgtKH226n6jQz9F5EN
r2H5eFVbBVoxcz8j9GSHFSvOwfJRvTRWLVLBb3WQGnYpOHG6Ns57JXDYO1X/ufuE
nw+1x/rs+l8TjA0nMesHZnpqt/53CNzWF3IcCnBZJvzkM/8+7zGu0FuwGmHGiksZ
QRPboDv+pUXY4xguJnFq8wJwbslpcUxC/m0O4RWhvQPUpdnC15mAXD0W+Chmkaz7
VteOQuouwr7d8/fvuk5DITHNkmxIWDyyy6auulLgBDg+EfZCWsZfqWx6/1aiUsVm
23XFqYicODJss3nazvbNDx4fPAp57E8ohZ14zCki29ZhCRVRyj2V19KtuBGJ2knZ
DYFZiTlT24JiuF4JjV4bwCjz0QcYx/2vb3cPIpMUCma6BTWhZoMGKrpXLylfpswP
/VPVe/DXGpMqxny03OQY2yVMQfEOtOqI5RPhaNjTbp1QHLOMpaeff7lOKkBFL92j
tk76oK+JsgSowBR4dNWStJqrGjEgfztwZU8KFmjGWW7oDsjEFyVkWYnfXoxj363f
krs4ZXCHoyT+5HWpHx/9QXaULryJmuhE9iySP1KaCynXhMYU3b6Jz2DjminBVon+
IcMOYS6TRGZXekPeyLwreXOj2RW0RppVGBGqdGUiB1KQjWyhKxOrAnf3X5l43lNF
Z+e1RU0PSUwOdv5KQZZnf1LOBU1SqiMiPSBUlwTLggjIW8opRilYISl9qFrOFl5f
jnJzNnFRbgLsU4ZrWXYdnCqlbnK0XDVnY8/GY9VlVI/bojjH72UxEpwaR2s4d0/z
k3VeURknbrnhpbqXaqj76jExJ2bZIfC31JXsVTvn5L1L/jAMj3DEumoTx+q6mXRt
2MkwNUvs7WuZ6PTdv3U4Fujg84RuMY2MNAKxh/LS3es12PkHc9avWNfe0Jf0R5Vw
duobY99HmOIgddhK4MAlcHpOzNBrMWm3QyfWDHr45vwq57nVbBwvqdJmqQ70XDr+
Dq5mPlZ926WYCieTdzdhp1uOuh+Ua3QTm4VBSYYY3/f6Rlf0wLjEaeOkK7n93KQg
BNdjQa7vhcjUlfO4QQ6mM0TcTJVei0EaS9KDGjtsiHuBAS39+kT1qry4bpjsE72A
89Jw7Y9TX7aRG/BADxdDN8AvAeuHFa60CHPJu6h03/59U6SeAHwsI40aWW8ZQdud
4S1/KTsHYYI/+EfkHkM2hLkWcHIYi0yXzEqgVUw7YAXhoJVP7wHN19ga/K/eMC8s
g6kiovnK4BVIh141zJa3QqoanJpp++kmbPwaop2p9jycAbYnnEK6fng+4+fXanuu
PvYm33lBYt4IFlJXL1IlJz8iP1fY/qvSo+t43KQm/UAX1vsXPVuK4KrqqX2rTUpH
mIzUb5gnI86r3NvLCJjXYloVwlQjrfGwBxg50vy1vUjTen8qPLwrDrmQuge+W1Co
vdmcatrxyTC4RAiuAt3Td7W3lCS5akHT5eRaa+i3XIRdRYmDLMRQZcUY8MUQNKVZ
3yI/VjusJICMD6rjXyKPCEIcTTxFNTKNGTqldtixU+zuiUvRD/TuS0IJTRaXARMC
OY8Oj+OaW0B94pObikH/1igTr97eyy5Z/KlgOYwP/AgOUfGZ/2oQC1SA6qR+WYU5
lk8R781hq4tqfxCdSXcA6L/i3WYLc0iDI7LBwSR5psPuFzhMxGAf+kFpksUI4U+O
NxfyTraJBJwLwlxJ4SRXEbhTB1ZJfwSrLxpbCZ6VSKWhE+JwazV0PzXQVF6vmCsn
O1mVY8tGQwigyRD8xKsxV6GvO28uGZFhdcqzEMzUk8yQ2zDlppPv0cX9NWI99llf
ANYD8BQj5Sn4scrq+o+5TqluI+XkjEeHlAo1/AAcXp7/tzPkAY14oMoliN4gdsdh
DzVgZpqdPAi4NhHrOXEpvzFrCpgeWFi5TC7ggvcw25J5zk9QTViPNvPQqdVx7yee
asxQftGcREmnVtZ/36hwOPyrYBwNFgZ4gZ3985SNKiP7ICmHQNYEdoDrvSO8ZJCV
mXqHQIPvTzb8dgw/8zwGka+BsfHeC2yth0Xi/AF01cCpfcDiG7dgCTZ4j3Fk8B0J
pRqO0XK9vRJ0yZORzEwUV26CHjbecgdxnBviXmd79A3auxumBg5Izb6l6wljDGRr
dB9/IcwKzNyRyNiGQ22qyQ32k9rDfry7OyZWzLE2T6XHP4YJ6BdrzCGQWeQci3Jt
LozrvrGLKcHfTQNgp2nRdyDpJLqG5B5dxTQ8WsBKqvsu5vecx/t3Sc0h0Z0DcB4m
`protect END_PROTECTED
