`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
diS8h2nvHKbD+tfGP9UnOjjlKJUpAbpny0uiMTvy45LhLvt9voqRku7i5Ckxi1Ky
KVYco46a9rzRNOjKBt1VZTXhil6OMibc9oDnkQbawAbECJ2cwXmh/In+djfLC3qh
B5TMotX2NWGa14tTE+XIR/e8TUSozPWrkp4+RC0J/zFL/y4xZQfi8VVxdwwz/mya
/7OCuog6V+Ch3NTx4mR1yOLvDH3R0xVR/rbp5T4IhWsheJO8XWLdtU565Te+ciQ1
k5BQ5nSpE7SjNwfw4PycYYAWz8n2euu6rEuzHO9E2wAQ4VTez0rO1MS95f4VnO0F
+2I4KkxcnF1v2mw7HZbDlDmoCjI+3GITxxeMrBtx0fTirArMDuqgCsTd+seugCqt
t59QhYsw9VpGPl1X/lKwFXXNZBsSdzJNSGHMm353FpEvDSTyjgzhGioTpjK3/nWH
3ow47Je+I30rNWfxRVhqcpV6bpgouLvRFaDWAbhf5cHqdB3SafNE5+crB2G9F2Fe
uWMUV6ZuH/C+q5Q5ZhbtGbiuwrPpIzwCSf5h4BhmlOBX0dzHrDj2BB0vOh1b4WMW
tL3HBuLJhNZp7POz4wWW3shITyUB86+zxa/qfHa3KC83dL/QYqjveHEqEmeTn8SI
JX/CslGrTYpP2GbX4sFFIZnuSUM7YvUoWQvQqVH3LSGdUOzsu6WbGtqunKaEsIRd
agWYi7Qs3ddEKCOJqxBNKAgfouOY3mDB+F2ndVbpkMp4AzT24uKOcVh+MAaFslkY
Yl8OaL3buEWo4ycnkWFPHDk5aBYhNJwMWn0BerbHIgjIxNiShh8cM70PH7gxNjqC
eC/eN9CzleJNPGT55vDNQ3kwW4YTnfv536fYmYUCuNyf26xPlqRKNczWF4Ndk/vl
8dfnOMjJ43vUTrvMFmH+wEhNtQvYkybS1fBPWgvTUO1gIbrjrUWxfSKdxfNvo3nl
xs0PY83BlskpJqOATkBrcAh/+VJNSH13sSTWZFWtqh/u0NUIQ0z5rWBH94G7OSLb
mqyfIpU0VgJhXfE5MRVt0/0L9rGmQLcQSzY3cmqVdvXsru5Ty2hxM+vfirmcH64r
ORQyTx/nSo3vc18OPJe1Qa89c5V8p/k3ETY8IuUYvzsrGf+UI0ybtlLVRsc8jc2T
8SQercdlQdwx4XxrhgSf1vrrSeTo64GxlUCx7rMmPysHEg0Xuf2bN67RKIAzVsaI
vaRkvZKaThDktTfZ1MlyW9UJSN5fkPpw36nTlsGHMv5rck1+NoiiKKoXimiTqlW8
8BlSg0/HhCWauuWB/zJH5aW23nRogQ1C+kwqV3JO4eJmYJJoRIwE14JnFxHkl+mH
xmbTMnq9q9ZbDbB73qoD6M/akgk1GVtd2Rpigev6Oup0/gr/ekOedor7hIEMbiEl
DEAM/nqHOI7ITiLmouzy6TEaC0aC50MPwdfYVOn4Iu0M+7vdSykYURSYau5dD1ib
1DLAqeSsKgRqgloMOXTJDl5r3Stz9+1QI9lQ/V6kRl0VWuK8RRI3u72B7F1+4uxd
UsjwuceTVdmpa/gvyYIrGf87Gty14re1h95jiNQmhV6l+1yJiQ/R+cL7gM5Zvr+X
bYB2JX7qBZnRc+teXu5Ut+O/QkOCU9J0MfBvfyIEcoBHAFzgRMcTqD5DjUK9wOim
MANVbFiE6YjsjOtATkGZfsOOe7U8haahrOM0aIhXKAM01MsT1O+VRw6L+GzJ0Phq
cQSMdXCgE3rrH5ftxaeFNIVVBXXIeaL2Oar/UrgKN6c=
`protect END_PROTECTED
