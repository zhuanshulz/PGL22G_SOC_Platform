`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pVss7oooNSbPV6eIuPo8lVKgjaeDQetoFDNUm89vIOir/8jpGpQbh9HdhIqWhRw5
A/yWfuHzv9em1swM/CcbNQ0x1m4uw3VynwXGyH58fFKtcvxEs7DvI5VBKke8BPVw
aBesV5sL3ronnRLaP5HjXeA0D7r4MC/pG+48kGVVG4puu0ld5ft9WBJ2Fna34CDQ
tyFOqeYAD0P4mC9NxzgcrZAI/hxxW0uCOmvHfJoOZUHLjLKiyVcB00CVdnrjMAA4
fmWQOVaRoT4+ek78/XVjoQSAiZH63DDKUNVcXCiz5nEQOYEj2PZ60MYk8ekpI0du
jyn44w7XNxlZC6qGV7Vkpim40Qm3vUJpLZwx/PmpXdHB5UugpO/jSYEnBRbAFqWh
wK3sQSdIQ+26zC/GGE0MxaclEu9hYz5ZDf0pJ6E0ghcF11fRflbJIqy8IpR+KVAy
iKYR4Ce/hsk3otn1lu0SaPHC9EGGCOK2zt7w7XOC3S2SaeBHUbRttf6ve4lCMUIW
zTkUcAiJu0jvE5H55YoeOMLe2K8pf3oCEN5ZYaIMEx3yfa2viB2lEEEAG/rgbQOE
`protect END_PROTECTED
