`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ejamHm5yWhCmMIg7LQ8bFfzdl6obXvukyx5AcYUJrmlbmSsmXuwbfZrIjNGGNIgt
hfOOJowdZocWYEdqbkwNmJFYpxhFJAeboZykT/QnDF1NH4j85sAmNVi+W62TWJCK
yQdqhTahAv55j9PVVhJVBELebYbDTFq9syLTYmODcQ6atwKeq72L7Oi4UAk9aJlp
e67ggs8BfNvP1mHzD7RQASfMtDfGhuMoX9IrCL//7aYzEGzO943plfpM13kK7uYR
q5mUdggW1+QcKFCT0ktgykrUL6a28jZjIV3lg73vBLVCg9mDCpRksjdDhMH7k1Mb
FlrlBz9xZTdtdw0UReiV4wgmQjn2/NHgLRrphkKu6m7kilUlyMdAC2POuUfR2O2M
J3fJRgn8fDiuAvR1En7rxB262R1I6Vt/3e+zJxnOTUrVzTpcI7/qnVYdFAmBRz6y
9waD8dikn/+v9IjNoNs/oC1xjim8ufl6OIfLWIoNvvR7RhaRrFs0bjJ39OFG4tyL
7vlZumKk3bA3+Qr/1vbVNNFGO9QRvJwMt28tFFctvZ56pIIDOBSXu5lqOisKk7O5
s/kys5OklPJmdsdQ2b0a4fPhT0uCm45ppVg1Ydk4ZxCarj38Pvauu2OWS5NxW6wx
HpMm+3z7NH6cGC1rrJRCFKarpk6rFHt5ogOBnOiIvXXuDyLREYYWnhmYXcPKib6w
FFRAVfUNy3ZkzmtHWXN86lirRXScz9jKZLQKURbisAq2nCe1SNMQzJ5+70XK5JQD
0SZoLygZRlueLymbVqB44F0Oi2CR+7SbRUv0/6XNHQbabG24DnrT9JIXvVSQ6ZCa
6mS06G2BkJhX5VN6p2jf+YOKtcHg6MfE+4NXV/pU5uZC9Ei4hPZ97xvmGAE4moy2
crXEmU0OpRqCJTOzsV9EujgkLqSi0qb5O7JpgudbepNFSo2eAeRk2dWObZe/jT1c
PUDNA7tB3WAiev3+DI0FjoxxgWR0kJH+KEuZtaXdwmxFG8eANySyBruEWSQAHHJ+
pL1yhw+Vk+JcA9iJrUn7CrzEW2HWh0FiuX6sjN/zjToZiQY1xxe0xb/8hUOeFNGc
GwCXYmBm5W99dpYBtvQTphzgjzyuFs6OEXWRXR4SecnWvjjeAe1okQiXeIJLmBvp
gpnp1MP9vsifHras3IWCseFDbbdpU6ipq6i4GfNMcXs7/J9po8FgKfCWsJ47VF0a
dz+20d4aePsouHgx+TAHrATbfJCDGDZkJRd50SCtAVeSlTXgbB+QD+NcIp8JgY9g
Uku1Ihkp1XpvN4fYCyN0+cI1oI9xDzlGsrWpQMU+rTy+55wc076ueJQhdCi9H0w+
inuctqzJQL1XiHLWprYOqbM86u6VdjCe9tV7Cd5Poq0TTPinlFAYWWjRrtfn6OXM
M6Oc7UzauxHdd1dKEvhRm0B5f6KCZY5YFcqB37ZVewtgM5oLmyYWGLXJ9TFBH5A9
9yJ46jsKO4Z9uv4MXkcE0dszR4YQcPnGb90T3RB+Rz09hsEwrrle5hgph9CbZPgO
SSJgosgbHxCYTwtxKyq2IobM2xWsAb7t0FiKfsYMubpAQvh6Du6JNvAmNv0SSXr6
VWDmyFyxjRyO9fE/z1sbiMd5CSF6cqJESfe/N1T3ArjSnKOPDye4aLLc9wUQUHo5
gbqGPS9WihEQsYhPKR7XZ1GEfH+XlMBnSvwA09YO8cHGPF3XGC7wBHlHtT3WCL51
qfnoZwGZYMS3AWi2NGSaRg0koYij0KXuEWCCSnjBtdQQY9Q51LFcPk/r9EwPfHiB
fPysyEUmc6yiHMVTHb+/42e4xLxvzcASBKISZdnsKA35IgTw6zo4hhKBcvzEJdFO
vXeQrIcoJyWka9O4lWllmW7XaeV/+DwBsHGjBoa5U44+5Rozy438himZ59c6yl21
xooVRQsi5cNXr+JlAKIDZ6sa5Wcdy1n60o/Dmzj5bMcPfW3IvXuPAiA43JdKASOf
NtZxkkJaQdpgAOpptmF01mbE2/BWuOydEjPKBob78bRPuMiy++fhQRdaHtmcLn7G
geKPH+ssMl+xXogo6UnWcTrTV2ieoZaUHjtS9EA6wxDjnGXE84QjynjYdSI6USZ/
HFnBf8FSWw5/aa4R/Y7abSqGcVs+X8DWGa7oUWISgFknvtLPihwCa7KvnG2oq45x
g9G9FBNvl/OoXCcwrE5LKyeTl2r8aXNWwSjdo5xyG7BhfzufO7gNQ1SVbdC8NJz1
`protect END_PROTECTED
