`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O1ksQnZsOE44S7wGQChrMwjb29TenqiAeuIbV8m2qS/Z1LRL467ewdBcWdoaikD4
m5ltRTk+ccGbK6zEDfgLIugjL1H5UeB5SV0cCEaMDI0N2yYbuXpOTwtXqgrMmqjg
uQKJGqHbr6w2wcGLBMwKdgPwMGFbEt6NAHahxwgQRcisMSHGvnB/cb6lnwFIV9Tt
Dz0CTqvV6B8yLb9TsFqG+VrMZI2hdEf6uoFqJJArRQmIKjz2u5VTQkyx4Fu/l/86
dTkNvOyOFZm7vCiteAw6F2s5g88vdcENme5bprHNkWz0flzmYlIzZk7zc7gZ7ye4
WPDeLed01dRV61IDU/DOGtlyqTQgHdMkfo5U0W6GDBGuWk5q4gWWYab+8MqIJaAy
OelsegjGPjfs6tYy6+wV72KpBi8qhuBBH37Pxc+HyWmeT6JCsPfmcNQdBBFK1Nk9
`protect END_PROTECTED
