`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/a9bZMbcCTARRQoPPYc44Z/wWib0Xw2/gptrBG7yiZNkde/WNfPGl0pVCeCB2flL
t6TVejCsBzRNTz1kYwEHqXwouuHXix72rxhokAssO6VeR3BDGfZnGkyKEvLihXBp
IzWEgxwV1pEOoMLPpAWpy+icEVcLobxYot/JQe5/xxnqhphW5ANe1ZWmtvBRUl92
L6bzbvEY+/03aXGilj07Y4UQFZoNZk/WN6Mre9DX8meX/QyXgI+esYv7oLxpej+6
mVXFDClKuxOYp7ekcS5z0ceyhKyCDt5UdR523EN9yOacK1eM8GZIAQydocIbzCoO
LHmCi7Zdnyv/yaNaILpatF6foO/5TT1qtIcSmE/rcC1W8HkNRpv6BkkYdi7X0kIZ
14AA7DEMBxyN2w6ZHG52+K4OGxCJGqKLIDjES4adwCb3aphj2v4HTM8FgPhMCLkD
k//tZvoAo7PtgFYt0f6YsjTZfObI1RXDYxnLXDpTvkq+JYUz3uQdfOfxhxiPF4VL
2Rs5xy/1xb7NwTKxWlDeppp2IwgCAXOqcWAhbAl/+7VGwkQMtQ+RNbp6amu/zceQ
n5t0/7sWZYyF6jWoSxMgHg==
`protect END_PROTECTED
