`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nm+n2PUbs1Wy9DhKVRQvCS5t0u1iHhVc4cJ9WePQ13XBbwu0uZ+Q8xw9QpjcwTEZ
C/LFtw4/tGEKj2CjeeDifEz+lq6MnKowM7fPpnZ+k/hzw7XQ4xWxekVBKSREPnjm
UN4t7I5xCnDUrPW2YL3xmoCJ41zcg716cjNizNpmrHoauRRzz1NqKOrKT9Fh+5zh
GSV2KqEEZtcUYU9DDchts3RWAVqdDq3a4e0lavvTTal0iasddGLKhhDU6pmhw3AY
kGHbAJIVZ1uDFyjxrRcqCoS9K359ZIuOn5IXfIBe2ynPDdlp60/o56j5iwvk33pa
cQY2zeves6g41wQqWt+PrdRCYw7xXNrXKo5Utma1ejxYD+yKGGgWoIsIuVbpK2XP
TttSVL8mgmnjUQoWM+mNU0jTwQN3uEfzcIcFQ+96Unz1qHfYW/2ZYMFIhp74hA5Q
`protect END_PROTECTED
