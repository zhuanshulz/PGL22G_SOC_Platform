`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4OD9JVS06oKgzKutC74gnO1PgfaiA6jbPBSUMAxrgm6/Ux4eSsVCU+399kJP+ll6
+nh28sAW9ZKUBgCvrE9K8bB2CFSCanzZtpDpJmhDw/6jT2DUqY3XZhr3vg6gVa+3
DUGf8L0TKNeatQoV4ziwWalyhmyIUeVbwn/fbVlm1cdfFevnjoP4c0Iv3X1bR3Bc
9jh6bYwqCATVtHfy9hgnyYlXIDc4bdFE5HZKJulwwwIvfVyB44kS5NhIMN06kpAR
UTbrWd+eihPT6iJ66t6PxhmrLdYEeOD3n9Lqae31Ya0nM9IqDHkp3ayn2ebp1/GW
Kc21KwvwpjfVsBfZ5OkFF+Amwzm4HL/HTbNxcyR3MxQmIZpCgsLOITHBqan3KwLd
snKxoTmaf28ghFzYjM9ee9z6J8mcFPqI1YKiwfmmGcKjf8h/7PuWIFQI08UKOi4s
8wdTUlH8Oo02SV8erJOExGnh2d/TiOqgCVwdYKj4e7ZOvxomX+izc+mt4AOy2m1z
DL2mhWwQukHFN9oEITBH3WMtv5NxLOJE+p3ehKLISRI4dnKRCswuCSolQoccnrlv
QrX1L6FuWS05Jsr5l1n8LNb2AVlqYRvUxO0DZcaHgJY=
`protect END_PROTECTED
