`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OFuiH7l1UVBaImQ2xwuMatO/pdi0tp4JPG45FBzMsRZ3BhLHHtIJodSS5qVRtz2y
PSRFBY9XnoYkJTC0we2Quqqiwy2Hb1sX09BjH4ow4yojvLZ4tCM69CGW9bUqcJGA
PcKQzjGIpvwvlGrKfA+fe+TWKRtgQBuAC6k+rhkCdGQvHK+w3phqDq7rQmRpEyt4
Ok7dAkiyNtU1+eBIe7JN7kkgrm72ADB2F9KKF/oZIewT0dTDMOkC/BCHMiHx0lIL
ELr4M4VQzoHkqJl983WfhZ1+gq/7bjX1JHhFr1NY+67nmJH8hPm3+6NYLa9EiT09
I9qWxtfM0ZuSL6SZijuc7ORxyOJIhf2sz/O1nlltmEnLex/HAnM0q8Fx4KqPus+t
A0Z2Ksq4FZ8/hLrV2Vr2fA==
`protect END_PROTECTED
