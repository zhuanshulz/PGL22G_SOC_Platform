`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PmPmI6q9iV60kjZotX3LZ8U7cUxkMer9TyjZXLOHvso+eFhObRGWEvaGQDeG7pq5
q7MmLexIWf06mUv0AykI+4FEZszyaEzs2YWQJAjMM/6OCgR/LpE0Z3v0Vkba8/zv
w7uRqkvauz+B4P2M6Ry9SfQ3V/vqIRsc9kMqeIcAk4GyiDeLOEwlo5EjFImRUaRH
j/VK5fpdRc+MELXOuSAaZsZmLKcvFNE51TmsIKoL4zqBvazC7CF2IKO/OEdOBnPo
QtEZAcMoUr55bS24E2jzJEovJYK1OVy4BKgEfkfCW5cu6COUIeGKtSp9OLDVLzYS
yca1V5MyDYzRtXAd10va9ulqm5ukhSJIuUMOR4CQcZSNSO7RhDydqfYrnOek+O3x
4MYdaPN+3NQ5BK6xH2sPBsE3TQdGVsQvdbQaF/Khc4KzzftUPyDKeOWmgw6NClyh
E0B+bnu1ffADgPD88MgKpA==
`protect END_PROTECTED
