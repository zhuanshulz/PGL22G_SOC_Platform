`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iwpRrtN944fHS8tn4AHUr3sLvQfu4xGfnBT9u+N+Fd9Zv/sRmgQh6I4PM6dkUf3q
HLFwCZMSOuYTPzzm1UjVptWOsUAveKglRL7ehH+yDuB65f+N8PDl104nZiowTzqO
+xFbM1t1oSSQO+o5mDEo8NoP+/6ynBkYBaFbXqJ/mYbcptbSqxFwMkmmGv3EeFya
BjnU7AKnhtLDQTX22m0ya5zZFrE82muUwSP5N7WM32OERfTJdCMYYSqiR67sH3/W
MZSxiOtpcKyUJgNyq+87DSwh8wQHZhdaIR9u6iDL7b9O5aGPdUkXkIfNZV7T3Z7g
941NZSZY0cJT2m3oEWHyRYY+37wK4sAdB3h+EanX9qs3a/oMoebqJmHtk4uOhM1A
AowGy3MvROLhbiTP4Gp0q9JtMIyiO+jhrY6M0yt/0NJ+8+O6d5Bxi7X7320QXYjh
/fjjd/6Eeb/xMxin947nmLPpCIDK7qEHxQXWIkmLi1LOgAAmyNcd76xLPZKVjs9Q
26jyPZwpQzDSgKJukq+yLi/BNfnkzqQJzVL9qby2nAi1d41mAO4owwZlY6j1ztuo
YJDzGkX9/FlnTz1nQF0CU27gqRDHiv5HsZ2AdV4cIVb1BH2961Dq5R3LYyQpS81K
KUMW21ftcJNKNkqde+GFf/b6UMuDEW211sfYxcIVUaDQrfqtPd20hw+GlATUGlNx
/WYnDYggl9gmuOlZi2AoMZKDRpoVeT0fxAqsMLbgsNoeC/lzN1S0OBPPK3tvE7Re
5aB+L862p7egO65/koZp/XuCAGI33vL0XiYye0FiW7JC3WAM4RvVPymHl6cEQ3At
QGpGCXEmgnTMBpt+hdXysJglxszERoe/x3mKfL/zGAmdCDOQ+Qa3lKCcZW22AAhI
h/nn4IByFtEFdU36haJPLjhgKICCNz2XpIuYhfqbcrgKjdoDfvZd+BtCiULqoJZ+
SZk5jDCLz23EtGz2nR9xnP2nJokOk4O/360s1I8s1m7d3oCeJyBunYB16TOYa5+a
PjS+fawR8HEViEkzaJmOWMJx3vN9afkd9dukz6v38kVH7mhMarzka67dk3zIJ1ra
1CfkN/n+1RpZk26It9wlTSpTd7LmnouCXJ66bbBAoRztQ9aagkgarcl1I+pmgR2n
OuRH8KPTdkejcqV9DqtlCh8q3wbz5UJHKjgE3yg0amRVslsXH0zepZB5rgIk0338
mF1t5dF2KEI+qL5u3UEpuxLZsOpssUdk7tYaQkiTsfIkgJddOT98/I7bQcDWPMMk
YZw0Pn79NtgFnwqIN9Nppd1rMvY86wmsCfQX9QlOPGnKfllXa+t4QAXRisbn5VcE
by5gY1Hsr1ysEkdvVjBXAoP9hBf0/EuMgi9azDmGcTel6BQiHeSPLKomiGFBxslr
Pe7Iwk7nVemhZnmP/v5bIOQsn/q1k1qte3gyfiv/1XHn4TxtTeaCJXmq+ZR8avzE
TrdAXXS39rBmuhf7q6BFK5Uoa9s8Dy/2mBh/pa4wbqJAeiovhsvKOWE3xpTjJIbA
VMLD+Jsi/FSFgj2yc44h3N/By4JOFP6EtlFOnwHBTtSIaNhS7yP8f5AdE9HdAXG7
6aVzZLjmqevOMNpyQXqtCfrGVoPUFyCDDYltARPgBTXSOPQv9nzCjgpm8MKgzHkt
GsspmdLP+p7JN7MBnQDqRf7/ONorE0dJKEhbaeNsnSGks4IFeYK7aLQ++MA1AO3k
PT6EkRoSqEBdAGNz0cNsmcpItwPKrTiYly+H2aFlBKn3rvOzQBjNK+b5epDl7FVD
wDAHg62nlKmJPPgWhF0rEvqJUQ7VDgK7AgEjxKNh4TzyQpvMz9vd5ghSQj3iaBDC
mGrdAILUxS4ZJV0mtfDj/shEan49m7ewlgK34u1JXLURpb2LbMaE+C2AX5IEIflw
EKtnRGY3aEJ0/rspQNB262Lw6WOhNNEBkJb02uMiSsbOaPeAv/gp7ZyTg3FsnPrx
M56N6FLYnPiNBAHYGfe1w+V95blfvobU0N0PHMLs8z2Ni7o+XTPKYAYL5DsP6yBK
crsJ9cKgeIJz+uuMpTiYGiUTRGfo+skxaY7jNpVN3fOUFz/awWqVhmlgUxG4BmoZ
h9m1PEHzMTBf2P8e8c2nki+bLhf2y83IGcbXvuTU3xY724dBE8hceo69KGitVTp+
sXAD7YEPK5y+GzehxuMEJlXI+BDtge+5snjMcMP5r6AgQlL5uRcdlNcHJm8mQ9RE
ASnCABp45+WseuKEhFE1UFwcDvSQMXS4yauwXCDuzRph0yG+T/iA6nyyBObdEB8V
cgxTrcQbap7e+lY9RZCeyvqyhLwdrUU0H0AZ4LzPDeRcq9RV9dAdG03jWcogvPOM
76c2IKXHVA7wxfxY0f/JqagIJUw6VKXB01y2oc8iLfOmuaT2fFKf6PK91e2dZZXQ
s75xEZCpKW+QvbqoBpEknJXOVygRZ0f/N9sYgm7xQY3OJlJjumDueLPNb0sMEVns
zBPqcdnmlAGt8ZPanwSq3Tx1DXHTAEeePloXAMr48lwjqFbvKx4eyEpN8SOsPChs
KytC1KMN7eagxrERaZwVDKA6zlwf6SpQRl0Hkqv/knrI9dvnOuO4yuc/6kPcJq+v
PCuwkwioXyIcHnUl5XFnc+3i/pddejRZStNTskhOE/BAg2Xtfib0K2s9w2roNfx9
Zha4Tm9mH0N7k3ynUtkISCB5ZMe4xidAydCNe1k3kPKQR2sOqJLt2lheDg+1W/YJ
bifPxqol35iGaJLvDpAbJAW5KSblcKAJIg62OUIE8mjk0O2oTRC6kXzm95IS06xg
ARh1ZUenwmLJYgAMuNWmDsaEhhJDxtWVtkoIyTs+yZxDy/NHEif9eM7mo40xPZNE
Ov2dvxmIE+qmirF45Kf8MpBB9I6y0VSb/gXeqKG1+/u/tMZ0Dhg/a9i6lq+xQhYv
rbcsgwE9azBkDJo5Ww9vFZoLJRuBbfu1gZ/4UM6JYxxMslvq7ZWn/I8OKLbZ6lgC
8+v/Nz+rtC/TDDJYSconqX0LHKXZuLpt+4FbdlrNxVCr2crzXINlIIikgYuokF4M
sh7QfSJ4O5XdfO8UtRUwy5aPqCQPbc7xvJ6RUIKkCVymO2QNevdcl8b1MId+lJBK
NVNY45QmJ3Brhq4BTm6xde+976Iq0rqB4pXXnK2Ru5PFepBZ3lmqZPzVDCUuszNJ
O/wWTJDjnEixIqEe3yHkhfn8zeVD1RoENqOmLSTNkqpu+IFtP+PL6Erg2st08CX2
u7Ca33mi0I2QSUad1KZfHHCdQIOTuiMNyJezqsyD8RD4cgY90Enj9gjDZB4R1sKw
oqCG03oZIsVqi5JQbnj+fadrNir6U3xxjpQGPlN7LVQCazML01BIShMvC5p0cXkO
8KYQbvZqN/BzXePr93Oid0VNT7ZPCI78ShAkjzVFU9+ls2Fy8giQvNm2ffJnysD5
1cBrSAof9G/LghEFrlO++ZmpP0SiyjMrosYMovPG4VkhpgCVJksAsn7oUvhTZCHB
ioX50vMioU5raceBunKeB5CNiZKO1SVnY4KDetO4lvUZwChb1LnGKy0dBHo9v9T0
wBcx8n07yV88etvHtq/GrwXP88RY8OQRxUTGIb4hvKMn5KQltq1I8hPGDPGf2zc3
ugasXVVHNy3QarDINFd/J3pzw2t6qM9dgq1Mq9yHWWqp3Nj/Afd+lgZrGxG5ur5I
mQNc3LmGJKJpT6QolQkIbO5BxJMEes8tfqGNN7dmCrZtuIJJu+MweOuh9fg2NlLY
ae+wXk69Eb/0e/oLICIrqsj3T5nyxKJ1krtGrU6BYiJPYZhoulW5/jADomltV/7x
duaIWJ+1vcAAqobltWI/F4yf+Q4eyb1q/HpOsKQ42TvVCLgwTEfBUe60YjDnSMdh
mfDz4ilf5gJh+4bZoPnjkdxmD26NV+GcXCVaPvNhitwtlWxXcazbDlRoMDto/p7K
2vISidMwGUzh7pblyjyTbmy2MXwHcWwKG6MleufPEJPIXm+JRWG53TkerCL7Q7NX
8KYvIlwAYXywqhdGx/muMjK6/GbtGXMvT6DiXbqbjaUII9xW55/a0vIwNrFPTCiD
7QykLPYATXZENRo+liTPXpDjJE6eKFGT6xCxH/TvfyOrn4x4KCBghsMDfvZxqkoR
EkVkxqWESXwy+CeF5pwbcR2cjsSjzZudE2x4U8emrZU53SwM7H6laBCk7Sb7MJwh
KXQufLRa79s4YEjGqCWYr0TIlp/rj7hljyUh1kQx2e2pdk1DCPYH8MTuv+3ITfPw
vtLSEI+Ewbp76yzM6Pz50pbyM7DhqBUR3rpTxRreqtlp5uqOyn3x+jWj05dq0PEI
qcAHqT7flSwOISMfpswe+lEBOgOBhUqXN+ioHG4wU2pZNS+TO0Wq19XGgc40+Tf7
hrjPLP3v1jamWdHLOfEwQMNpFwDcdGH+HTWIrmVYOAceM4htfF2vDfg1Ah5KWEy4
VeYunldV8FDxpsE1lTx2q2zLK0MO8oVc6GPBrZ+14IfDcrjw2RSKy0saInmsKZcG
NZ2ryrhyIzTJ5lx+N6Dm5NleEH/Qgxb7Sm9cN2+ZkIeJXUa7/Pt7Y9Mn1cymg3+M
1bHbhAfZwp+5PJ6wNl2YZZIbrpVAO9e1Enlc+Lp5FCsnxlGfiiYvSI6TjB9emyck
ucop+B0sLvlA6VRgrBW7Tw2ztn+wBSmicbUybiCl+8KBFAmcLWFFGxNRh1HiTo20
XNQMgBUpRvxGIECJOnrcNLNVtDtgwx1ZIiRVkd2oDt/hWa6HD6+cGx+s/FAYlFEx
zDVixRGV6qs/u+K0OEXVxvX8oUBTwKvX426s3L8P2o5OJrHnFc18U64wVH7dCrrf
UVr1qLk4zqiY7BnaLyS2xBmZDfgJaocafeEX1wqu0G1mhFSXYcQU9x8JKShmHNEh
Hs4oebpPI64mMbB7NkTgTT2aH3apEg7yJFJHZAlYtSHYw0AUN0pqC4b/x9uhNa3C
o0X1h46/z95KGxh8Nnk3+g0abwiIUGEwCkwHbVk+Cv84Vx5AXeoou32o8dE3d3Vk
Uyizo7tN8gnD5hj445WRNB5TeBoerwg/+yLiwIR57bCdbeiVbf0uafqkhsEp5JYm
GCooo4scKmxFbrQf+ny6uTDXmTcV1G8rNCV2EKy/n4As9uNYtKVHA3CFwem3Manl
4AMHYali1WOWaITP8HrkTxXzNgj4sod+3W0oqqj9pK5mI5ieSU2MS9hbcikRrX/2
/hKqOCqtpo/N1XdkGgcC3VVg4AoY2V7GFDYr1FE8Elk0mvFyRPLfs2FIL0W9Cjp+
TPlqtQoTx0B8Zdp912EfuFUIA6AJ2p+mqxqC5PBUPPgR7IU8r8HGY7XZqshaLav7
s0o6ET9iYkTIz2eKVkDLcGAid3FozML+xs8NBZnwkgGucoYAvQGwJDwsAaCAWfK2
Q2AKu3hZr+pvBUlO72qTKsDNO++4ntEDqtpje9BZNiTxv3fOgWWdufRNezc7lV5v
E4gYitYmH2u3iImtWcCU958CdSbsccFSofPQyplRoMIIVZ5bvcY+rnjaxK720XMw
H9P65QRzMbtxKOkCA07lnsSYIf4GRZdxRR3KAosmUEYBogBdsZThJrG+jUoYmy+s
WuHsqevK0Chemu3UegbHG2KBQn+eW9PlqUY5hJMrrqoMYPVMOHfTFpMUiXR1RC51
n+6Na2t6V/NewfVzFTP2axI8tjD1DFQXbYy55s4bmTur1/kMAwl2ig57qMIkbLBe
bg53PTmKZqQZ1dXEdLaTPDx17hqhRyx31wBe78fb7b0zbo2YqpKq53gs9vBOcsca
ZAbQBS0BvGOiwCFcZpK6GtY2Vm5rnSrpEZ0o/XbkxEeFTpAxQApIwXguYWtoFMeR
2ZJCAn975ntJIcBkJ5bZ4ul/xLBW9WuzX9PVluIQKMUMhl+8elz5zuv/nRlJoTzm
Wl3z/wCdvVj1gXB1FTd1Baqbi8gMDgwXyk0EYgKRfbKmXIRo1eSVpbPCXx7aF/U1
+Oa2Jt5MEBGSdTo9+CLPmkw5bGkfqRaRnOIClb3YryDobm0toOSxsg/vRWhrSDb6
NmfUfAjasUuc6twQwzzLaW3HoR8JIOqSGk67o2n/4Dgpjk8F7P9RfusY9ZW3HLE2
8lfGh95ZxigqI9+aqka9yDeXET845d9pYF5jZUVZBftKXG2PrxNBCeBEMMylfR87
cXI6hAQba5hVaAtpEjr7Ca4/CGtY62DZSqNWePwcVbcaH8q1DGaqjxHI+Py+vuhM
6Pnb8EFv+rHXcoCTmxX7AdlOqSBzWkFiF4WDrt9VD14SnkrN/ISbciwiSwsOGdBC
n7IgYBsMjC/rQiomW1brhhgu0x7N+0UlZo8oGwyUkWN2lQoNCW6vIJhLwdVJPpyH
AuTaApkHOyJRFTiQCSjl/W0xv9cLetB15TVGv9aUzu0fwNdKjLYTQvh8LnjJAMtl
wOPV+H8vXuZN4y3xlWZAW/X+2l5SzW0xiPDdtmVDFwCoBdqC3BtNt0g/qbA+U9Vd
6WMVP4kGGikbKOSzJj+889vO2MgYbSMZgHtHDCQB9TBP/wswrcWCu4XaI9TziPME
4IRshnmWnVmbe3riyfixQFlHxfVUQUJHMSPTJSuvddZDzufa3lSOhxFH1gZYPomU
TqKkDR+pPkuRJGiIY2nh/RqSRtc7Gd0OmSS7J/xmevYYQoP8pT5JumsapdbGdwu7
tJBtqSw6mJZXDKwVAwPEEI+KbL14Jxvt2AyvFDiLuQhyFh+OGpZZiB7QqD66fdYR
c7PEFxHt7jGPLzBYfegRCZGKKJYDABV3a6+3+dexg9mJEmT94kNdAcDfGlsGpIa3
nFkrbNdrSAon89IQNGH7Hv5blQJQzpdlLou/VZkelF2ZQFG+6T0kUEZP71+vm1Mw
zCZS9X/wSTpss+iIIoMFjmSTqL3qJ5OvuUkBf9MxjEwdm6h2VquuGoke0Om1XJka
OHs5H9AV+amlU1gLz0T7a7JutGEHHXWJz0QSfdC175P8eYWdHvAQcsCUDYdbMnq6
GWfTgPmFlj980TSO4zIChwVF/DJgVUbaIrZm5VfqpAkc3ZxNKfcaI/Qf5bEipegZ
Q2LrBwG3L6VPKL8I4ewns1pn8jvpK+voUKGYvX31CvPO2UH9OgKwkpk3Lpyw2ZbO
TWbyM6oDOH//mVItROjscW5tZDMmDqIwGzUL3+zKAAGvOm6s9hRvFevOPTWcJxso
7QkiQf/AtZy8lkXvGe6YlctQZUYkFV9cJjzbnBw4QcOmfAahlG46gph8Je3MXXAH
cs22HmkfkSNl5HtPc8RG9SknBdEp8YINKjDT9Wv5t4gdDytwmBAtYb0UFMf/4YFK
g5YvBEiEUl/u+KWvV044Ncva6XRQEUkDZKZ6ab30aNQ2OxVerfVumMUuuZxT2C++
OwbNiooz86eAlAnkyK1rI10GfjLtMY1hXuhNgFyJHN89qnZtM053MRtHoloE/qFV
rvHOcyGMhrUTlEjWZTFI2zAjcK6gFPwnWl2nzDdov8AtLP3wWmXlYV7xjiKQdjQA
9ANuiqmaAvl9O77EehFFqq4mtYZM5LnJ6fUeyPY5ENZ/VbNxCs6iRqQ5EF7Ht43e
nR9BdAvtDigffNmoroEy1CQ4PZDyPQyfATMp6sk/nyjEfoRggN0z8wZNO4HqO8hA
nnmILotLbn8kVB3+y9UsNZsrxaO8HZtcbHtz3dgmgtX26Qcd8qNwx5XOFK8gl2re
I5lHdYRjTp2L+lF0lFh3a5oJ5HasF0NjTdjLAcwfQLxIPddcYZ8oiZ1d3EyqloEO
ylZxnPptG4p51KWwIeglOGR/Jjpb/eQZW9j5L/AVZef4G0nOpO5tO8+FxZrxLpU/
B4nIfSIegZuh/D+XcvsrxBlHHXz1t8itbCOXC9ShCx1kgEBG3WZuk2qmdvB7eIXK
2KXiIBR6LslY6SMzF5bstEUk7dHntyrg6Kl3jyxL6kvhnZLoQrb4SgaqL3swCGTQ
GMQKZBJkZug9b9OYpQ/ZYw07sIHIOduuQBYJhNcHsT0BIwC/yL4Z2Oukl09mBqN3
KfZFUH5MUgsLM/xhFTN8BT7ZBhl+5n/z8mxAyd+8PKgBJyuCMso6yNMqSztexXIN
KXqAsq5WNdr7iSCcb6dexwJXNNs0SjhveiOhtFge7IwBNMlyKicb9hyR76Dlv/dS
RVCU5WgGccr7UXBgHR5F2XKt8gq9OWKh9zFVtIWo4xjHsxpjuzVry/cqGg5Hl+QU
d4InTXozcpSHnQj+Zofdxhpjp+CRISOCAiQF+va0ifZWq+8ljcNuO7ZVT5XwctkL
t+SjLaa5D4pCODG4slgn7LuxuQpHVQxz3YipEWvJshWzWtRYqUB7dzw1yW1lWgxv
owBeJDeY08HlsGEi2KrNkWgwDQiv3lbv8zoNWktoyMx5g45W209ayc9sCrBrKo1I
FlDT0MXT7fyL+S+vZvBGMui68USPGeeLVzpnHf5yR3Dol33lZMLxsIgN1satGIDd
LxrvpRJ8DGEScnxge0N3ZTFyZdCKWnyTMl/4aR76Uh7dxhlB66KKwWIR/IHBOZKj
OD+1mKcUqF7EnVjs77u2upWRV//lBflecu9hrUm3ymXz5CTYax3Gx9X67NF4pizE
K9+JkEAvkSn8Ak48DainOs42Jj23Z2yQLmYtBxutt+a/kjruXj4MYHKRnEJtYdp/
b8JdBTa5bzjb03dhIUIVVNNI2kM48GwkdD4UfDg8t749BqkL8WM+12tJST1PvQUN
52HntnkUQJUuxU0RzttzD01cdperOUDsbe7O3Vtsu6MtThsnv+4XtLCIISzE2QXd
xVvOSYOJJRbBljgCzHux80EuURXJzneJfk72j3sjpXSHFMrOXyCQj5d56QjS6DH9
MO9ygbeSduGQBPADGsyvfvwTGZDDab4YwyGtnu3ge/9CNM3BX3AUnxDyLEeLK621
idP5hRl5KfDwoqPMjrr+D6kxg1R0KElebduNwvNqDl3NmHu8hIMjUG5APX79Smnz
smNuNPtFeDKLj4WA8REJQ8InQDkwqb1K2arB556FvT9e4ivDQ6Q+BALQXj9kd3qB
nqTHWqZFyoxVQzXvKoonYMlt0XAzzTooZt5zY8WVGJ92tVc6oI3/Mll2/Afxef45
ea2Ibl+GV5bDl6Hix8fGsvWnyJQ4mggSn6b9KmvPs+RUE/FAlBEA04P/woDnDLM+
3hjGfi96pUZOHBOq1CYs/YQUrhLweGFrF90+vmag8IYy8zFqvjtvckmFPfb/1S/u
uVMRLnIX3Mtf0LXwL4zt3GuNHZ1s19IP8JwJPYDKR7PSIv7iw3vIvrOklZ+MVyWf
ynKb6mPjekbpM23+WO0SJ4B1xvRoSNnHzj33kcoX1v+BM+vkQ/OE0smZLoeuOPFv
IDt4jHvQsDplkL/3nGRzCr/MXaE+fRH0RQzgujqrBslQHcRiPyKQfVrTgCDavfxS
R3k5VRsEMjkPt547Hb5nxDY+spBC0GZLRY2dKv1vjUC87S7/4CL73aCcAQJ/LfJB
4D4RJS2bqgaLqdNa1h/MiqlnqByuxOV+C6S8GE2nElG13bkSL63WoZluO8DiFlPH
yuF9vvUzhE0KH4sVG7etgMkvUl1kWz4FKL1RrD9m8V6FAaaxfbSI7iswGV6BoGIQ
HY5HNVFEhJiYSZZa4CKCoRM6DfFGHcCjk4xhUeBQ34rOCEcKpnRfTeYkJZ33bGO0
edFIbp7SJ8QcyHuJm49TdHPN0jYclUEusEikKIPqTt/j55mfwJmX1eqQdsEVR14B
MTy0Duv82ojaBO7DVYIQJZlA1qMwVfkRg3E3CFrgOJxtvIqlK28qrKNxAd7jdvL1
mIMT5KeBpC2/4+g0UB9iYI+bqiMJ/l5mh7hKT4II4b/fdDwJFd24elQi22QOXp4u
gu6oeCsHoMqz7NrBXXsEo07No8E8GfeLGEfx3NKkdDFLkYhgluCIzDPL1jydxFHy
2MBOKuf8/qQULx3e77dP9G7wRB+GL/+ruPWaJi5PBQqcDN5VMYr2OmZkrbC6p5n1
mTECRMCvPzSJM39zCi6LI5rdYqgDR50ogLMPO2eqFvezy3TOsXzafIHNP2PantWX
4D8EpVWtHQGSgCcJBokH093kXTQ2O3sHBZ/CWsd9R98YdGFlHC+wJ+wb4DjrVcuy
eedFtdxmoPzMhIKx1hn0OmZsxim7dPYphiVFwVxN/cX1z2Wf4KlgBwefHX5lsXoJ
SxI20YiF9WlTKqQ6HvEAurRipSmgKwLRY3t/ajfN5WkALmJw/Wii1Abbg3BDRNaS
hmN446P/GYeup38mQBbr7LXl5yFjRZDwywiLBriXDIb2FMugwEJGyfkc9UTDpm5Q
/h7U+f47WadinLMg1RBQJ7oNmrBEswgaUM5nv0uOX+XjRc/s6n68RdFgQkwpN2Pb
//6EUXEB2ZPA5x2CHFjnQOj9MF6Ayh6Qs8qzTRyQEzpSjMTW66RBS6R90c5tV5EO
lVJhC1mvTmzWMfBx0ZgbGNadRNJlToK0r2AENfe1sg+aw+diE/2dGmWjsDjFNOyG
qGt0yuzVWq9VQ/eerw/zA3Y16U5hqUwzloi/n91vE3K/IqU6UrO/XqBDmiZAUjYO
MyG++W1kvXCM/RCwOUcxGdN2cSTFMZIOO67IB1/NZyIzpbw0Dq1gDfMvE6a49Jg6
sJyPR2gG4/zSXMl00Qlkd9HGgw27FX3We/VFPDhvxMsItiBKQx5L7uJI9K42OAuu
RhxMxq19GYxw5+fThiozfDi6xuMJ6AKgA9l5l24HOHRQKvu5/2ACQ6yXx1XGe508
XG4C0xo3RfE31ZerNj3OoLpu3RujoB8zSJwrS7bV4JHzc/VHgg5tcI3khCvr9mVF
vE3EQcEncCJBoB+TVb3EbA0uO93HNbcbS0Ih8GlyLGfm3jqv6G3PpnMbpJZOQELQ
0bZlPLakGCvy2OeUxkSdPJBu4/VKIVgR/fH2HYjTQ9YDEY6kYCdtYSH/YFl44xnn
RYtAYECBuPOS9sa/9ZIXM4IrQ8Mg3ZljIPktE9V0cJbKhPsz3TFkehiDK8EhA4OG
GnGNA7B1/7Ey1Gy1JDSL32BPTwrbopTq4MdnY2Iip3hFmPINR8UdwBdFWonLZIO2
L/bi7pcyV+q2QBb/TYXdtEksK3LlS5M1dzngfgcgeeMJd6rosGZFNtbXLgSkNtdj
GvR4EOx7y2iXe5N1cTKY+8VEXWG1ye0Fr48Boa+rwLWcWnm+6TFrF6g6xhSIWbDg
kkSHxkJg/Txrgm5XnLNxANwvz5E1JQRjfP1wK7wBZzXTtrwwEO9SeHTdFpQAgoe7
pUJdHLpuKIqfLGqpKisxmDjlinsaXjgfECZoSEJeC3H0oq1y8Z2guOTobniVWTJ4
WnJncOonmflW9otnR0y+orTmhKUlA20ZSz9QEzGRXuNNbMMj/AF3kKmdfc+fBNwD
D6iU9ElSNwH34PUzfDHmQjKnLdbxS7eVKAtuLS82GYo/lLb8ltOhpETCTdW3KArO
u7oVQTbCZ2vNlKgvVUerxXQKJk1dKhobkA02nnB4DSCfX559fGHB1OgfRvNVL7+x
Vig2GaON1uwboHjScQrstAPK4nfliLtpSHWJeMO7qWtf8+HcRoYKLatJviY5C13a
OoJ8W+ZKvD5POAXAuxmQM8+u/sdcpTkPvlY975NKIuQKSoTTbrkpPhtAiVkMN5VV
N2eyi6q7etage80DGa3U2+jQQZ725X/vJeIXhIsL6RaWLrNvJgLu174ycANxuWw0
JiPK7HqRhh5WABW9k8ZGN0VEXIAUQ988ostxk4f+J+G2iLTz0t30VNlSpihXEX+k
AC2RaRyMiQksUPYwV57MAAtU3Co5vQNBD3zo9t3J9oD6gU6ZlItlcfjXMXtmK/qS
ftsV19wrK17l2121xskOrkptx/v+AA6Y3WLdAkDTDI0+oI3D6Yticnh+ccAGwFSg
IcdqQvW8H4q5/i64HuMtD+V3S2baqTWOOcVuDSbcyiTl33qYAerc0ooBss983lY7
Wi7Pq6h/1iBhtJKoEkGMf51CPzuYg6iZDmEj2cr4mVOyNHMzLOok/VRwGQi+oKUt
gDVotaBkDie3jnEA+Md5W65yGtFsKWY3ZtgC4JG8v6QOUwZuq0gV4C7W9okyZ6pz
MgVzpuFioTshysBDO8ZFmcUaAZBXuGcO9qVFYMkPbmwn5H8P2tp8nDB/mxauRKZt
A6//3itf5YA48c60NW7mgFaWCtoV0xaAauS+wY0y786D5TmnR+MvpYsxEnZomBux
oRlVc3YeBietbr6OdUyquwHWf4cJwGpoNnGlERiLXxJaptq+IDb+hOLPLSMFHtC5
kfk0fMLTEuWgTAlh/VVnp1DVcs6veKO1kcw4INByLKvcRHVtvK9OBKpdAtZk9Y2l
h2FH/dSFa+EK/XFJOpSOIXlAxcaqqtecvmMCS6KWirh1D8+IUbTvWPvQPQawYEF0
r7BMRklWmAVpisl5Qcge6CzMuX63bfHcuoh61GM+ZpzR/q+ESd2hkiSRqDXGLarO
xsJwEnTXRHxS8KQpdGIViOEvmkypAzvV7pQxsqHQAkTwiPWqUWYmd71V+Zb7sPT0
2qYaNq2vsVxhloMKmB5kA98kNt9JKlr0fMsvze1eWJV7BfEfbMIAAyJHGemmcF+0
XGQuAm1EgJCffoq+ixH7WLilIzthiJ01O7m5LoiQc0zLMf62NsLvROSPJLkaeOJD
+9ADJTebRtZeEbkAasyqlnNu9aGVJEHQBN8ZG5qKDhhEp7lsr+AEoyjXe8m92pLb
eTIjurzGrH+V76MSuu2GJhHcxsiZxP7cNinaGfi5DTVrGqBo2bBoeCc2UNRHLPNR
lKi24MnXFL9rDcHwXav4exNQo0oH35K5lT5mQUbDyiGfiery0dEoahBNu+09Hg5g
Luu52jMWowgiFL7csdfzDpUrnndc9Ja/6/bBe0zDVFlfJn2F72EkUB9q/cU4gD4z
/cKmjFJjMWlzlM6KXVQ2EZkxwnkspPxaK1HxBBI3r5dyevwaLPiZhxa9g/wyuuEn
ZYmkzLgH8ONrKKQAwgsm+tf1l+Cn+5VPubz3m09U/9ikFVE5LQ4fiA5VwiYKFFxy
5U2nPY+ZCFUZv2aqxvYRu+apl4kYMmsV5lEMFmYEH62DMw/VreYiK4xBUeWeTWuC
IuIghUXJjbtq/B1Vsk844ExVvfD3lF/PeeXKRu9XgzkSilN08ch1o5NOge91mf3D
gkzSySPNhB9x1f98TYFs3IKC8NLF5ewx7qff2G8ZKDGCfKoqUriA5cHIVA4f+bIR
hlj7Zmyjupwti17P3XtAs4hEzpb9kObEXHZU1ejz6i2u5mpQbCULKjsxULA3rlf/
LvWVzPGsq1U8/XIJOQUfoMs3IN1Ejdbk+PPeDXdUpGGfLhBg+4KW4BXi5JF1uTqR
ipkG1XfWRr7x89U35EMklPkbITWHg5Kqed8/Ryb6h14GxprlRXglf4B37u8qHk85
HRaz81Blf2evKnze0lxZctgp96aIELfWX+wbrOIuBbDqvQgU561ZbQH0DmRNBmY0
WVINUR23lkhoNtp1fWW5UDcBtLkfwojUl2zpncPs3mGlgG3wM/LiLZnqXFRAZjGn
Q5JlXtNDS9an8VKD7LHV/8h6OrxTYzMprleaRZJ5/bEAY0KDVXYmRBx5Qy3Iv2zV
/AEqZZDf0+Y9VpU7HICQpMOkRXDYQDVJAZ9PtaSTiF/6mBgU8/j7XjiurWoTeNxt
pJF5rFkVmeFBxjaecIONnO3odIIv0MQj0py6D9POBzYJal/MFWxxknBzbYCcy5Mn
qQl+kgTe/pR4UWvWO26ti60cA88N7WKA/nwiBcC3T+z5g3RUN+wZXW265h10V0N7
5hmDp0MjKmvcwwZISJkYABkNVCKun03gr9TtIKreQqf+ggHb4WSm605/Y/nUsa5R
Phhx9FFv5vEeAsQvcyZfIL4GvmqaBCXykOeKdIazUyusS9p++vPmYoCAOewq7hzv
Zy+oh3hmMRYhW/tORJOvYmkcExvYzsn7tk3PKCqRImUGA/FaJ4LPROjFA/LFWBtG
nZuWsGSxkKRZVQgPdA+hqVx+m/KxlOKcf7/8l+vLj4A71eCo9nMD1DS99MgOQGvf
Dd7xi0YwwypulEnrJPaVJxrvPpBxPva1d+/Mv2BOHA9/WMNPAOM7G9ZRIZoGjn6t
eFQCjj8NxkGc7IDMjbaUWizxNokMTWQZDSW1nqtygs0iphHJAabNIpvq7ubDZfa6
zOduNXR73QR/PG7ABL2Zbz7ih+khNxR01ALxwyKT4WUUx0cq8wFIpIPcUVXiVzIo
ji7n3M4SoFcNcdee9/SWPLDWBgWSCGRBhlysIjK5tjihRtCN1X9SWlKOu+oUoCHi
XKSlfo1EG8KYJFRWK461TZ36CX96dRkQajCrebo3I7fwDZOag3qooSeai6kfIFPc
wCFhn4BIdDXMhbiQtnhgEicO9sJgvtZwCbFekJvPfqdlOS5t+CwpnHu6BOP0B5Tv
a//q8LaUhKeBomRyrgS6Mh7A0Jg11H4STMCX9ZdHXvU4nUyYTE+FCMCPesVf98sr
E3Saak053DDoCHgUfBBx83iD89dzYiVxF5OSHsUfzWtDAUy2Vj88ry3bTC19eobc
QbGpFnjovygFkWLTZoor+hsf9zzjC79Gy5DjNM6Cw8c1ycKlJ4pZlMh3CYZanggp
cagGybGal/7knWyiaxVO4KC3vUUiUhBxQQemUl13awe5TLeIWv/YNu94QqkWTchw
0DTZWMQQDSgkRTp3Tw0t3WpOg5b82eGKqDWJLEqhJOr7qO4TAqu+TZ0TEO6/msVu
0MZBBe5viv9bgth2QXvaMcjmJAU9pwIaDxlQNyFzWW+NDkE5DbnKw5I9dDRSqde5
uyAjhmmM8IYHtFuJM+mf+kRgrouOQmUnwQnzDua3+yXQLb/hKAbuZ1aese7uj0/7
mwM6gvxwjcVG5PeGVNUSzlyCt1MCtlZRAnPUxls2Q26o5SW2mW+yYi6dJ4vK7PzM
bpGEI012Oier3LscCIwAQMEykNbfufTNjcoKWj/Ep1f3stRhtP2Whgq0WnWJDN1k
yP7iHl4Ax4WKYrdyk3q7SPWrO4q4zFoXUfNe5Ze53Ux4HQwwW1wftZL3BbY6HAyH
iheteRtJWdDpmbzGISXEVbUpAe87uM+Kbm9ek/+qQoAkS4p3m+7LuwX/nsPghWyx
4YUJCkZvlGDllH4oKo0mvnL+KfHBEZS4TZvqcZIadJmylxoT2sK+7+e1QYWi0t28
OOvwv+iZL+aTLFzKEGhSUpUT0OE8t2W2OS4ziTBdAvgfqc7Osur0VfS2K21PDzvF
mSD2/vkFDGxJGPy9qgdAT8RGUd1xexZbCHrseYSYi6ATCfSvDRrrGVoA7QHTKDgD
l594wQXP1add381pDQ+OEHZcpLOibM3FmvMwOaLs32EShXOim8aD1E9yiOPqZ03G
tC35FpArCbxFMHGjyppRcJ/VUVrw/zyDDni7/dylmfFoJnef0pEeOtM3OX9J03Cd
YBv1VD8bJs0RR+vEaZkmPhTycijQ6XtU2ajTVkevwHjZPlqRs226Xl0D5cxWE3Ow
r/k767nIwSE70Sy2pSapvBigM5nWg1lD0tSzEvePmfosg8fI7qfuH5uFx4Vec5az
6hXRlzgxi2W9dc8dzJ0P816j0KhKziytOqoBxFXSYp3cgerRbV/2kVzY6wsdN0jh
YbIqsGzyrwEsb2NOhfy4fmJQj3W83PNBhjM+jJGxKVES/LugdkNS5P6AKEJijamt
qnwGNlWN+rl2nHky53v9fViGEsCighTwZCfE7ejEpB70ovVI18ArpBDPelMTPU+d
jNJ4drPnN2om57Kpd0PAPFByH3oaiu+TUUNsAD15e3/m7lVwgZwYpYSAb4WqvGrH
28IIkJvjiYLY73AqG3OOCQMW5TXTBTkZabSpapRV8A4pAIhm0kOvCQFBJSVDheI4
wijjosbxJmBhI2UYF64YmLSYUaGV5nTmagEdH7uWRBKW0Hjyr6Q2uRqoBt0SDaIU
tmUNoLq/cvdCxEr+zuAai6Adf/MnvrT8OzyI7zt6Eb7fkN5F4S+bOng9O74nVj4G
fS/P2KbJ0dww0CSUCnlbh7XthErbrak2VAJrLngZrwWkw+7keo99gA9eKi1aMwAc
Z5sNmY+BCU+1LswWtjF5J0+vJDP1nnB3ehx+4qaY5mIY5HdiloFs0enuFo0PNZqi
LIFQuPJW0Y9UZn3+poLphYSmmxKK1vVy6O3eoHU4hg3oyAfMB0lEF60UjCWg6oRF
sHtjliNqh3T1QLzxYbKZA8MB6OBjTM6QwiPLKTamz2rd9DQnW34o2wRv9OnHMe3F
iOCWFaUXwUWJefV6xDzC4KRF+SV6lG2cIiwKfANt6JtGEky08z/aYAUVWeGCPJFY
tvb7HEHW5/k5GrhnVDb8OzutC9GkHZzijd+NYL5R8WZJyOihM5rJyf3JDnGTH8i/
SyBCpltg8UVH7AcYE7OKmUt89TH8NQMwupZaaqjFJ9KSZnqx4qOMULyULLUGWtxz
w/i8uwub+LVn9v2T75xUu5zD3wyibTRSQeGMRHdE3JBKwJEKkwa8lQ6w2G8jk+wu
3/CUFx+vWkg2a3PlQC5Z7dhsgboYR4g+DMv2O6zBpzEavvT8a0a9/Bl5HOJGPgeR
kUoIusJb10DsleI1Kvjsm3Jw3futvHVM7HBCNXqzu9DZ5zkOn6sZa0H//QfkhbOz
Mx0j2ryLa0l3T5h6uOl36Hagdfjb0tYq3N4AgzABEHzPziT4JPShQF0kWB7H0CWD
HH7g8ebOT0FXA+8yiabZ17M0WcP2+wTs2KzKNDh3sj7mnQb02xjAKTr8Xe03lcyM
BMfqDXHPSNqUTV9xjqL4qKsxOz9qNWUQsngWSt1R7eEZ32SdVc0pzayfGlK9eeZ+
xBbcsmTnDB+B8IpqAv23Uw1ZGJ3Y7VVdmHjRerAKkt/xSbXAhvKM7jBc7fNGG5Hl
7HQ0g/kN1BToGbMKegcJiRJHgSIHBGK6M1aut6mA1Ka3Jbr/kboVyrTcvgSmg0PZ
kCDkuTVtCgm89676Sxwd8DDE8d9i1jLLBuy/f6eWSINPITLOUC0FAUE5ojCw83li
qV3ITs7c1FvVdW5iT/3jiuDCZmSOr8MaF+6DyLXVPLi28FwHBLe3DD/EvI6hcGL/
Yigp+sgAVYQ/ryz9izjpkmSHYwTh5dVDG74NA0YZ6OY9azefP7a6/CVTVL1DG4gr
6VnHsmwT2b5mLxsbguVFsoHyFQFGzXVB8K3FncDu7sr+gON9SleWTgHHtEwGRDTX
HQNTaPqFwZhHSBeR+NUKUTzGYrFzRlNzz46EiCcWndkZtx3n+pTppDRyrRAXvfGH
gU3wo4xHY/Qlsy5dzim58RU3/XOuyPS94xwkJTEES+jKLcIFsHCvCFV8ElIyQEIR
zLQWWD+/HQb3dYQgX9NnPcvRxrK/yGIK3vbrAntOEJMi7x/k0aNyuKoeJpu08SSc
O0dx4hbIuCAOcw3+oo5fcSVUrCtFTX1nSjGKUhtrxzUIk6Gxa84XXMKY2LYSDf8q
6bryFLWPPd+pBviFfFwv/kUQql917DMBJoEPpo/fjpq3WcWiqA5ew4Aw5Yrseqna
JNRF6/WWmIekWag4HExZw0UQnfsD7QK1gFKDak2h3nTTXNVCkSGnzfnl/CbQoXyg
HaAw38ruCpI6ABhUjvaaVimhhUWzjaJl0w1OCgR2xSgwSXtvrtAgR+qFyy1Rvr0X
6vS9yiYiVQaUL8ahHPFxYIdOmIqWsTCGLkxmgOpVZHkTg3aOblw6dFLN7ZDlPZgJ
LdJwl7AfVCC3r4WC5GzmPPAxLwQ430ahjcZb4w281EslVJT/7Sc4QVrLuqPvksY8
h7hQLwomTBfrdO0aEYy430FhvpAsJ1QcIoRWN1dn13upLufM/yZAxIiBSWyWLL51
QnvBwl5wak+jYKZ0k9RnGg==
`protect END_PROTECTED
