`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4lqXP/XnVQslyKOaANIowkDyCmpRSjFo1nOW1h5RxDJzEJDocJ2ZoG9nS/+7LuNF
HqggMsJpNivaMnrsuBZuDG/UxdWtsJQUbMMF+Z1A7d3XYK/SZ+SZfm17HroTETvq
gFmYC5LWbfAlXcDl2YatlCpZDXQ//gdCHbpUWqjGJt4n9+Sg/R2qHq+rEv97v1wG
EiqDOtNP/1VyaTK+sU9ZaIhgqItj85Pl0v7fRzf+zGpJcbeYTgv8E7A7BJtte0uy
d0V0sZmScJtmTC8HnLAuFt+G5qVEO0UnHKEtEUJqtSsi/8l1+FjkB78s0YtLXvPH
3GEl4AwbQg3dhrLarnrrffW+vuQYl9/35lmVfL6SHR/9pJVs894rXj7iqYvuXFUh
rsoepg8i2Xk/V4mNUvII4Nz8i6LDq5PAp1k9MAZzX1MkaaNNHJQEebBndvOAGUPT
Vm4ua4miFkK1dFv7Py3a90uhK8UyRdDxZYGqB3ymdWXzFIBGgA6mQV0A+yQUjsCA
o4RIaEJQWNg9+qlS2DaC1tP6BLMN5jWeJM+mW+BWGobp1hBP2NwXbjGFRAyqVwHv
Ve1B6TPVIZhnxaHUoZOfnd3yKGoFL1Cif5pVp5Qw9q0xdKwLVUN489G7Em3Jzq4M
zGL7VWsU/DyYZr62LhHwcLoettxcdebbRjXIlVLhbmlDQLbfjWEUoQakinF4pv/1
/lbp7UlpJK7R76+ngs4MeaZ8rxJYlRe+U7Zqi2rwgHA3CLhvrU4M8VFq/CEQh/Cw
5tNQZat//7KtlPT3+CGvYOYqIPjjiwYLAbk1eHOWKPO36l31lJoTMjmKCdTDfgVC
kSBZrW/i9w0FsZwNiuTHohLVUnAhUjPsCmLffw60A2HirZqQtoXADAoeHTo+BjPE
gnIa6K8unK/m+fd0UoNTaqvzmBpCfuWqTztSYW2rZBrDWX26YBREi8oDZg26U9zv
7SWOBZ89w5xNhNNEQG8Cn2At+P08dTG7Z7ekrh5rvJDr6fr0dnpoAhBP+4UjY2hm
KEcRNf2oWmb4x1GhUTBnxf3fhsdaByR/hPdlgpCxPnqBASJVs8QoddajgUU8oT3i
jqSY3sr3b9Vt4r8fa++ao9qP10M8XBJYyggs7YlPQStsWboOwDeB1J9oLbtsTd3+
DHEDIsCH69SZUU3w/TV+rEeglKJWKvEADHRk3bj2esnXwAJI/liKOHPazkxC5Zpo
psrT47Da642JcGoEgL+WNkRbiu+6RI9cC3+2AOkb2AVOzuqqdMk2yYRPvAeUMsph
j9hxlX3+sk3EChQXoltWSWKtxRXmO9gD/5ZuKhQm+OR557XUC3d7H+9OyGvzuXPO
6ExeJVC7xYLJMxgdSa4HFXTRV8HUNiIx1rULahEAN573SA1PS5GLqZRxS2sVUXOg
2kqenPlZqFvtzngmq6Qi60256XtOCObrDf/gF4okY3gigCc/RnZRh7GLPWoKRknA
vLfsqRVGK8SABR59dF4NmpyWUBSoRS2CJHHtx+jY8CXL15cZphCwEKB7Bo4FkgEP
MsHIJRW3CZtLCI9gvc28G81YKvbe1B05EU7rXZDIouiLXb6O5exY23yGAGHW+yhl
vv0ocG2NNtczkUwyglvBgS7Zjh/d+nss8HssVsqidgWtzjZDUi+N5pOmm7kqtPV3
g6ZEq1MneDh31TfPlmjdpwtfQAygKyrBuJh92lO6Q9Y8CJUeY5T4AQ3mwNVwqXoE
en/XuDGGqoNiNg3hq/FV0cQsg90IBJ2vzoSlf6u0FECadVLOtLFV53rdBrxCtayS
tCkr5tkPd5mhXK0zXg3I1SmFfncKdGt3tPVbUOlNCqgKy7TEsbVeemVVJv/SjsG8
ggO9XUCZUbtQGtfMrRs3LOisjQLGkAb93MkTkj6pHaJ0gN3EzWHxS6gooXP//Vpl
Y1ooL3itktUNXOFEAI5mG47ViFOfLT58tC/yYWo1r6Ecv/m9GeX40NVokHOcY2jm
g+doH0Zgc6fBtmkhyaAyMfgDGrbllXMIdwWPahPB7JBwPltxZTilI0V9fMm2MZnh
CD8e+134M5yJErWts+cDn/faoo9EDkBJfK/RReawbDVznavhKDyr2f0VGD44fijI
`protect END_PROTECTED
