`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oHKY3mku6qA17dhwoyzfn4XvsaOVbFQsBc2puYY8S3a4xKANCw2aksbT9/bKNhNi
QbN7BZhqbpiXQjRE7+Jt5LXbuXmW4g5lm2le86dDlUy3/17MjRxOpqQ9k6UdiSEF
4CrZdzi8vIrKfG099etde15rdY9url316mhQ5c1q4soJ8SDz+5RvP9NOEr7yhgaE
TWVBAiDe8UVSJvd5t48CDSxYFhlLm9h9WiCqzd5UXwc+jLzHm3RIUF+m2lhTGJWc
sMkPm0Q01ITSjmBcZ29U05dsG+XlcSQ7ws/cP2MfoMpMD1fOWX6+XYP0017V0ThN
rl04c6kApBdKEgUyQXbL/UQC10TxQTMCb+ldoC+WN/+ibF75Q3ogHPtxsNJsdFVT
O+VMqIx5UkulYJbMm54iXyOz1aOnmtmXKv+m20l1Y3ph/X3mjx1THhvjgqZ57i8M
EiqB6Np9jgIVbK/ZDe2o6SCdK+BPsCEBN7SsPxhnZon4zDpAMVaL1wjOZMMZKQk9
JqrJeUS9DqZX4lM59m4hAkcgvEcct/XJH84AhvDNfYGZxs28HWz3Xe9up4bU0KWz
vhKmTU7YxAibB3nvNfwH2ZtcsRiS5L9VhyXwLhN9FJVFRyJyNUAg5ZtwGKdI/CIg
8eXv4PhZZom2lr8uciGnHMp1FwwGEpD3hpqDdcr8cRB5Eqg2LNUvcaoFjtMk+tXL
kBx2qtIUlCXJ6X47J5jToZyQh0WeJNK5gQL99GU6wBgbUFOOq5G60yvPtyuZ/Hhu
MMGLxnzTFPOpyZFXDoy+9KEQ1HKUHCC6+hIu09NMeaYMRb9EqqEXrsLNx/RTnhL1
yZiDoFqgcZTKjXV8Qqe809MjkiLW191XjQnnJtOVnJSZo41pB2GF5bEBCnbWRhT0
ph7xVTK1wtirjvn8wxAcc2Bc6dxY8QBwEl5w2Oux4BMAoogkxOVe2lTjP8UXl9Sq
OIEOsAH6HyDMwzOiZIdZ3TN1UrtVMh6mBlNU2QMMAJXFcwRrPquwYnOcB3lmXfHq
w0HaxuYkJftQ3F9Ln4Ynd3apHEZP6XHvNtjU0ej5SC5JmZVRneLwr3qAaJaO9FcE
A4o433yuy75DL3bXFW32bEUyEiPO7XAVEgLN+B/99S86MY7yeaItteKzWf22sFIu
VTr4SHMHSK135KsgeZtqTqgThpauTxRkoJuNk7rjGqg2+/YZIQTwUJi0cjVyLyoO
llKmFcrb5a2xMofUTB8wH3x6nJObLp/vzAnZbHUrAg9lhT+7exFhpuF/yB4gLn4G
RzDUkGp3a1OLJKcDzRC0EK9SeX6NmXsNKuaUibCBToTPzoLiKcXYtQF2SrGt9m5J
AAFQfDgzghReBPiY9Mc/RlnVujm67196dvABHu9vrtDgUk9oInq8Wb5hd4qsrASq
GfWnza5m6JdnX/SktLEtDcZwnwr9PU0sIVCpKHOQo+q9rX5Ka11VI0w5vD3c/5NQ
eO79lAbpYLzYreS4d6ng/OutZ+kLT1RbSWWKJgkwbHiVzrK0a+Ug3+y2VMCADh67
UkMHrWYUhgH7TXgOoeS1lT/USOi4IXydwoyn7IW4JuL8qElyLiIZfbvUPL2gENk2
nr7giId0l3Y62QD86WNnNLGmU0ia7oQYnyU8xkNNaAvJuRS5TekJbXopqTKYkh+Z
Cralmb76UtgWj0gkQL28/3GVoSZoSpxWZYWTPzZf4c6nOGXUftLosYcAApsygGXa
Z9qPoHCehYMoxBQIkimnGin3HqB7xYUB8IbDdI9bIIJ3K8z0QPwUbLQCcfDTeIr6
JYuZGjZ6TabPN4oJt100yncxLkH/i5zvh4TTXJSrKTSFQyfRynPzHFbAn6Xh3Nxm
SA/nvsBTltOWW14GpK9T5ATXG2BRYiS/uPChoivrg3vzatESvJ2HQSEc5dxuPbsj
N4Xp2OjeLTanz0dnItcEWFkefqljumQ2Qwo7Qibe4A5dR6nSGGud9Hz2m17BSAP5
vIz5DvJDX8tEPCQgGCwb3OXpK+zAiNaNC7qisa1KQxtAU3uyq3mGpF3OTpqsbEpy
aXsm4PRlvdHw4UUWyG3aSdGDM1JJUaQGyBDoLrNvD6S0YwcVOkD5nLPiHCXh8US5
QTrA+Fc/T7bLAmwhYNIS6fF86rv9Vq6WZryhw4qRH/MOShwnj4AVwwlHYMEAEHg1
+6qyIG4Ew6343rxSI7/ZrsjvfGS0lQl4P1/QbzXAECRm5rAEMGrKQwqj7KnKSnUA
/Fd2gWJiDG2tXoXbUXFNJgg16UeX9+M7x93ZALtlHLyKJPsoVTbPF0I+Q9rgmzdz
Y5UOwsP+HRRcBuEGc4giVqrsET1Bx9x/kJuXaxa0WYMgTCcGkD0+9kPHhUxTVHd5
x3ayA34ORdZ+viz28GecxuwoXGZimyAaCyZZ1X1Rn9w80UP8uVVruu8dcWZ1alER
yFJ4urfADo6MSbj8A0uxsuHqvRq/2eHRMAzk1WkmUN/n4JLFmpBm5N29BI6HHKor
1qU5EoQZft/dK3zmNClVP8Nhwx+pnKTH1SCvp2FcQKAUKuoxSLRXzPcH0gKVh+9N
BZecNyGw/cHQSJt8jVpdysSLMWvF2Pc6XVVLMfDuHjQuNS3iZsMgqVfVFYR0UQUx
c4Qnb2UJ+Sq10DJ5EbqbgDXdd23YH/q9oAt0NMIYk8+2VOMKG03FihkBjQgfFadb
nGM+2ZLG3fnFqVNXFM1txghXJGlM9A3AKcK6mF7dPr0W7hsdD0xCpzZBJMsmOpxs
fyXOJQUTF5GEQ2m0L/8mhluaNuxjGMn8B9QRduNheeSC1mnuq1ZVsMliOqMHq8up
eBvU13+UOtf4kCyRnt19X9y89hgTrGvf593H8s9j8rKMRAPqOPrC7gIk6xl/HKg0
lttIxm8r+/uw/pGnvnvOX22H3PfAOfYGbBLFrX1d76f+/cuRwhGS4sNpt2OgOmM0
7ODFbv2qnKOXMo9TpQjZUCrKrbw4KLi6X4NlWj605OkC4Fzof/Ai0fgThlhoAvTx
U988kW2fvaLh5wFsVBD6j4aYVFnDpn69cLzX0dmdlja6vpsdKagBn2jzOYDgUXn2
YXWR/GWRWXr1R3+EGJR/IIGO/RUUA2g4mphPLlJcBbsfA74E69JAELezNfM/ahmF
EOYZGwJSLryt8qeqs3/5TEhDw3GDKvI3YsEy/FQDU1+FnOmxD+vURFUUrRKAGdBT
e50710lMZNsfLdNHOMPFXAi7eGe2r3bgXe8evSEP+IxuC84gWdVojx+WqisC8EE9
JAB1oxLqUtD1EIMKTBUx2/whJzUeiL7pF4vkeY9QQ/RVZPnmLLQU3oUu0cFvAjgI
w8TkiJ5OxvXCcH9q69FGcJ2z8ezX6lQXvrxStszFJLb4VvJZWwccTxjTa4VSoYs8
I2anjcK1bFzBmBnjBDb1HMwlP/aijQ2hGwRgVTGqjOVJg45GWw5dNGfvLJk6wG3y
Cx+EkM9/9g333V8RjXv9E3OOA5IGB8foELYkzPw99Srr82usdz1fOSePzzzE8sf4
qrAUVyDwhaZABKK9GbeClyDnmmPj0ca4zH9im3ve6Ik91LNplRKQKRKb3LwK9Do3
V1K0ELB/ZFyGBAYckjEvI770BecAz6Tgf6Vf+t3G5U4vjlVpD19YWRqtcuwNM05c
xFZvR3oZKn2QPoc27gaCCPgvzyBBeAwftA80dtoAfKXCEJwcMksHwH29sjH6GZLU
p8qsrAfIfjklHzrdTtYVkKlFx4rQuhk+o374a7SmD3BUx+VMiTlYDo02iWBxT+5M
pvPCAdolxKhibnYHCuDAwwt7Xzmipn8wOub8SXPztmnFw1HjKwsL1aJQMgz5rfHU
nI1hvbqCPaQOYTx26XxtiLgM1bxPdj4yv2HV8xO3UjzwygrqrqHORasGu27admSf
GfcblEdMWwkkXfVqBMRzT3bevAMFJfVXXBQq2dhnZFyYZp+n65bBrGporG8JhqmP
EKFCLBrxf1NH6uFTUlK25DCvgiD3KvICXI7lkmJttem7DhF6ZO0Srmw0A1I+2IHj
ULRFtT2yTsYA92MFG7NrZnQ5dg2XDkt+62SnU9fbqIJRHcI3/g2IEAh+kXOaI5vA
KVIN6PNdjjJQs5/eMz0dneQUGQ9Ue4X+6CmqqexRBUNxo78l5WHvhuXvjlejgVge
cRwQHdcs2UwlVMiKrEZmNh4sqblgDiAYZyxTuNW9apRGr0xWYRqUqGAvkL/qiU3P
wwzXv5i9Bqlb4PjWwi8NWtzhwlHCVtAmhsYQ4pRL4dgWGPUvw9Ar0KuZAsxmDVKm
dWPZpdBprZfWcB+MNTYClP5P3glrwmgniX12IKp6vWIu0qPH4BJdUbm0BvcnPk3x
Iln+yOU6PtxpBGrZ2pI4t4fnOcTPmvt+mOYCvsg7KdpT1DWa9NhiNpbAcDJSjH49
2q7Zx1wdCNgbwwTkRUOuMt8/LftVbW0WfJDWOzCOEbFhhTdh9ROSwwEQ9tKq5zcD
uEsuwObUavWEPoXNjtIeqcHY95Djaha2MDZwfIxmeeL4xm4gkf5u7FUH8MRQ+5fd
mnNgaHHgbcw48Gb6F6HYpprk4piLHgONPLp7hlzXj5OIlR2FWA5rIBfSJDWP5Zif
JPv2UyKLzGC5yApqyx7QKqMefaSfqWNjpumMqBEi5j/0FbDadHFiXJ3LtaTs3i1a
ORLKvvcY2TpN0nHvU/gpi3QZERivg+O71TSfbUo630X7nlugPbpt2M4cGzsGzg9I
aIVmYJ4crG1QHJuzpNsNupg8/9NKnaVo3We96eym3ahtVkvZ5FVkqfo2bTtRCTbt
/Whs75znoEN6miyzeAFN6QLAAg7evoA40kmDzUVH2FjxSb2sB8poduX4RjkuZ7Wu
92e60L+Ztxtf89Ntcj8FyXdKd9lMvYO63+44JnzcU+sqieH6Wb3EiKNjs/8A4fN/
eXhUKahJJUpRlTl56ObnxQU2LDHWPA8SEYvM16yk3zxUffIqV+UEN7Z8YiF/xs9f
fH81fODWvf3Kke3nNjEi3jqc4D+I2WyqlPXo3gGHyHqPm0m2QyJOCvyk0W1zIVrg
GQyOZnvbxAH09XPjVciBtyZQZVHH5wUaUhhU7r8srSJd4uADpp8PqK+SPq0tXExO
D4xyurfKpe5DNVACu6SQaW8eJNeA1+x7tC3DLOTS8n3JG1pdFn2WHtkasMMOjaE3
7/600jIe3FVI8HwAIWNpvfWIX+/EH+EqP4F9XP3YvWTnNJXwIgw048IBeoY83ww+
2Ict0CEh6Wil4wDyviohOJUbfwYg0rwfGaiQs1NC0cGnsBiWSgNH5W3tOejC5u9j
jno+8bKdwHOPdQ64vutP4iShken9g3Fydy8C8Y/qC0jC34ePNTlMrtin0WkYN/qX
T6eSvu94A6yOqVwOH2wiCSTSsl2XGUZg0bfQ7kquz4usNavgjptoCjn4xfcfSU8f
ho4Ixn6t6651nUy730o36geae8YEBK075vU96COHbcGN6jtcWfkARMbG8DUyr+CL
PvwyfJg5qYeXHDoKP/UhmcjPSXgHNECMi3rUDvlmNWFTLKyegRkpk1nlK9z/xBT1
5Lh6NnXUMZHykcC7jUn3jfoWmmGAI9el8BrloYEljLlvqBwZgA9K1+fyAJf9wbr7
Yffr9WKm9fSbmFWH3nxLdNHMG8MZomlLd0UPeodc/m2YwUa2ByrhdcXaktxWfnCV
066Doubj/ExU+ElPMMMqt0NmXWt2RN315Xa7gP5l/O65VFzfSAZuNKj5Otrx4YnT
SOFhHV5sRd4hvAyp8rKZfyRk5tF3/wrlzsae/wyz0j/74c+UfwyJ61gzZfj0Atv/
5Wcr5unSzHxwpEI4AEepk+5Gqa+p8BbqvOtAG8qurN4gOKqWEtcwRHtZ38of0gds
iEqgt6ONR4HYr4tYKqMHeNOHutwe5cOJu6TzcMI7z6LKCLhndMTIh2VbGTphdqQQ
uV5rwC3MfDHRtaMSbh2iE0LyGklrOebc/nAm9pgrzGmWvwoHQuqwC5j1H8HiQA+h
n4YrTdrJlur924gH7Sr+RyakbzkDnwGj/r/elvVeLHEvrP4bUn4zZxvdILjGtfvZ
kR0cQAPrY1YFaKKWQHJr089HmCkcLosasG+T0q7x4h1JB/uGoj+e0z6WRKB9ULeF
ues/wb8m+j+WvkBdT3jPeBGqpRi3OWrtUvQx3zkoXMO7xxOFoOw4nms5I5ypDdFx
Pjha6FRxovMGzRzf4yWhO7EJjWmjlIXhQX1puTEWG/SRVC9SdWzbpX4s5d5BWxpL
TbX/WDEd0aWgXqaYnW+uDpYo+KGSMv9rdZsTtCp9UVrX9dlU1PQok7z0K39vRu+i
8BxH8nSgcL35duj/bmYnvIhe+lf10oyB+/mPhOZb4i+vdpp7wquVolOEFpm7/Pw+
lqMVxL/HNPlRMERDnoH831WFK09SUVorV2p89z/R5OB1ObQyH6M+hCp1WsqLyy4R
FmQEGn69dIdrj6CvD1hfVUEuMEi1yTLVQRlOFTpPsvhwWo9kf/8nR9aPzk4jyIgD
4KbawVM4m6kxtb4M+3dykw2me0l43nas+Iee+QRKW4uAKe4OJkBlfU0WCLwtqhOM
dZEmKRXsFR0cb5zZfkfhVDCJ8dCZkwYuPVFYJCxwC/BqzO4My+KQMi0IlSWvvuNp
K/yzSO0uy3A1UfElLu9EGrD8gOYNrfv1uIIWhQNRXpli5MUOGTmlxTlawCvizqys
En5UZ2RlUgaImtl+U82vPmiZBDkrmFSPuwgxB4OeptN3GFDIgCdwkKEbdC4ihaMB
mStX2phGdYJDDoPvaQwKe05khMQIQ4rc8Cmp1lhY7euTk1Q0l12lJvW/v+Rcivsi
VuvLYynSssZtWX7eQWEUlq76u2a1cz80lWB7+pcB+gM8m7zj82PD3oI4cp49r699
0wJz8JAqBqjxd42rQuLzPVHogowEi2QDxw/sjkRBydlvarebhD1t/efoeSXXrd37
ZiU0x3IgHksk2noax2W4DHWsS5/EJEr4eK7o6xvLhHktTNTNHihNAg+LodrEv7Gv
cxicOKcjdps/FKinzoFxPkT1Ufaf21fyKfMtL6tOFT4xoMUBSvCZolCMxRN4rSzF
+VPTEcuWDIX98I5uxPcWqPKdXESGKSKO1j5yVfNj6Wls7/c718//P9c8lxXlKV0d
26fUOsehIUTw0EoJ6sUmy3qxw3PRhQW2rY9qHcU+j99ZNwGRduDCqbxHL2rOGb57
3j0BFJ4lzGaHfuRmyKP7i0iXxr21oZSlZuMEc2BLzdblQXzdkn9dLNyrTbOfJJWr
fcWaGixQAVGfXbVH/Pmc/5Byq7AquaPcJPJ7HvTxHjvVmo3AXjOdWCElZXFbo1b2
zafkaNsj2EakKm2WYzUONELl5sNQG3dozU+fdr4i/t7CMBonDgaq/iiANrHRotpj
qfuSPfxCxE7Dy62xBn42PQhInCcUkwUt15oGVh38ANHIK9nuxileFDz6qk3GJsdN
XAyS6inmID6ktrjPzKcMmdSh15zB3fQvdNqySpe0OeGmOvjs9C7qMxsQWEkDe5zc
A0lfroYm8s/3jjkEZgg6c+9uq2IEhsXFmmOl2zhUXz9DhQgc544oC+6cdHAp22la
50K+r3PVc1ahgSnmazs0qomNl+1gqVSukugLDC9ShkxCJTVbVG1Y3jb5wiohg5+5
TDDVbkT5YCWMCA7m7e6LpqvjGuOxkUWXtFQOuFyYdE7kzEW0DRsGsG8O2nDA0IPm
YElOCTrhsINAixG74hECx1Sc1g4RjHgLywrIf58iZu+1fP39lIEtzQ1/cZKzYAh+
PNkUq8fTGQQW3GE196HVVqJQEhySj05S1K+KNz1Apm2nRCh2mE2b/ME+O7lxUa49
bITgoH7ort85iu07094UPBRkkW98U9iNs6Z0f2dNag3ZZ+Pn8VHzy8dGyt45DZt8
H5QiG612oA20MALV7A/5x4z+AVF6rnP7IPlOuwItQEhg4P2O4q5eyBJPSRdFi5WL
CKQZdrnUHWFb4tM1p0UX7PcHga0oslVfLA4XmNE/CuyS2EBcg+Sovcum2kSGr/0U
ifFCVs170K9/5/+B+xMPa1UKC1X9ZF5Z99I0KAA/ZSs3ZCVLDmUffctGbh8b89fp
sNRN0X1hubDOVis40Jf0qhxzZdgxi0072iI/0lsE0Zy3YYs2bIkG7Zu4/+8aJZv2
Khi4By41YO81IGn+BxsTpxxvf93eNxODiY5xOIbnqyVp2grcTz8O/MZbmf6Z/UiM
tv7x9Y/ThT5jTzj35hLEkBVVvSQX/xJO1mKTuYQ5//eoS/DGBGU4JuzkGooTrYoC
4iFy82RnCxo/4/rm54qrNM9eZwLWxc51hciNElk9Hko/DtRTD1/Hu0q3et/5tyNV
HeOGWy3y0aqcTLgwfLiKPJeXbTJrQIoaqxOFeYa3cl24qwYF663PTaph/3EQvpRO
Mxtzn3T0qETBz748psMwrJwKDj0NXeOYMn6m9k/zORcL3UHhO9BWQx2zgT4afRqM
K9JDSOTWeNTQSM7M+NICqmUi2/1PwZMJZlwDm5SySxUUALztapKxMvl955Q78iF8
vzXC3YBo9xINV+69MP3m+sbB844jB2Kir63SckOTafVvX8O3uPtcvC5ZNVHN0Eg5
1x2Q9wTTCaQqv0Kc6l9naMu4RJSppMocA7oEpJoPH43nXsI8WqxHZa+3xykk3mNZ
mu14MZX83UnLApE0sJT3hPFWRLSno/h1KaVZiBs/7Y2lCInIJmqNs9FjoojB2yNH
vIawH9dS64HsudH5/YqU89jJ/UCJgTcFlcNe4TwgVO6vfD9HPNiiRvSoh5wS3bLb
/Xut7wfDRVGnS6YWCLMLNBPrdnmv0S5SeJnyQYAMGEFjpdIffn8qRBnHoSXiAtW9
7F+e1xezc7uCM3h/ZEd03UrvlnqmEsI2H+yvaLo1dm2nmibiptmDOtDvODYlXVg6
rA+xprZRIKogieBSDPfPAunm1VvWknKud9jUObXQKCAvnuS8OKyNc4U8ZpnAe0wP
Of+KOmyQaaA/so+84wqKxychh+Xfdq0CzQ/lqVB1QUhh/yNHFJmimJS9bfazea0o
k0TXIfiyTTjPgHDfW/pN9ehK4IW1pEvVKIg3fmhum5qPRkQmBpYmLzynIcdN06o0
vMiUdj8IA8bs3B50aMUD6UV5HyFcZRFzCwjWMtsukJvX65ALBMaIQ9om09TSoHop
VIPdxYQVbdQbc4LHcUoDEWl7/zfnR915RbXAYYc10dtGI7omowlGx8jxnNCc+FrT
/T02WfVNTohbMUHk3ozhiOK3i0dHRH/x/ffI16dd6/SRpIKdzIpI3UgYZePW5kOA
1wgnCDJ43eBpJkJzrydqBT7ijPpFrZPGXpCrjGRjYlgb0xawXlz6btmk9FM3O30F
Ga4elfyPglLr+erjhYRFcTtxG9Y9py4EUzOchRxyYGJlU4SILc2WlkDTCn54p4Ay
vdFGQhDvcXHIXDl/9JVhF2/fIapd+7JCYsRa8Ti3xndKn7gUA2EgqbWq7epVU/ag
W60mUHRVpI2tu0ij/qE/NGBPvXT1CHlFH0NvCk8JvLJpJpSJ/KdEY0Gm02mnfE7t
N7AYpXF/F1WAJwv6siEDWLy0BV/4MjJX0XLVoF85HaMDinvWl5iMKY04L7XC3F4l
0jn3pf0fbcpJpjPpB4lVx7EHF98On5XM8ee2q5zVhnEE/ZxaHY24ZE7FtEMEnQEC
ndE1eYxisJufsUgk0zjdeWCKQ4+utDzTAZ4zZCBS9jiehb+rntaVUkWw2ndK8pEA
LTLuTGKS5ZIaOV2dTEDu+/8sr0OcYPmCbwUSULsLddXkdJuIU6BaF4GzTrRu1u9M
yK9O7G1HEvG1XnIJp2aU8HBI/LaP9JN4uQl76mbrERUTUuCYwhUtK/z43q02n6lQ
jqY9ACIdjw3tVABBw4qMYrLfS5FM2rb6TJd9zf+qlaGlm2nN2es6EkMxm9sXLcLD
ri/UC1NOVlgzS7Eg9qw/wCWEqI0Os5ovwEUwlm8Hzg4NwjJCcaBppQ+W7GNScN10
uP1HEBQWmvp01uofcksmisvFheYoKdapKyoQa0TThenmC5kqjWr9ConZfC+IV6xD
vUK9HuxVY2v1Hgn1aNvffo7ZbcU6f8Yjk7/sEqkVN6OJdq1ZhSN0Nv2ndbhWqz8w
KN3uT8ZN7fcfFvJv4sUPlXG5n0MGrZyS+atylz1TGzvTicPGmk0lmkm67WK8H7I+
cZSz/PATDU7JO8ucj+sgAcDQ/6Ht+dlkcqRdVTjMXBcH5fY6HLWLjPp4kMJYM2PC
eQ9SW+K40jmyOOlLBWaNiTzZ3bjd7ThlS5Ye8Z/9SikDlYlAzprcINI5f3huc0tS
YNdAfcDgTq1m3FDvaCXrRcIVChU6M/lvnrGLr6FCtCjUWwUFViD1eg3VU15ZdOyw
k8/8XHqa+mmc1e00V3ovglSQr53UvdUneIikl8NhsYNmhNkOTDD4dkc0n9p172d5
Rc1U9UT5zfJSAzxPimxk6Xo5I3BxG2amQaBYFUnXMZngPRAlThTV3Rh2zeihhfSR
OPZRsp6Mz4v0Aw+DpSrTJK+l2cudnddvAVVNuHjy1RLeIjqYOk0phWuGikpcUCyU
bR2KL8Vm9B2s5Wph/BHR7FytB1d4/6PM1yuAVzZ/QIei0aRXRF1zqSUIMaPJcUKY
lcJ30/0hMf4XBRXnnBSZtoIUo9m0BVoTMxJfG9zZDSqCUJHgE+XV9mnpIChW2+bh
pjcW90oPnrV2D4BxonsQ5COIscYuKa1a/zbUNDNuGGXJbBS+Q7culGpC6vVWppAl
GehwGr6ujeDNjL/bC1WEkEJWwOH7UW+AvimtesEFN/+oB9SNZE7qIwFiHTluQ2fb
S+vfTmhbJSptsPf0e/3BiwphJu7rldAvYPZSjU9CHFR7lqiaexXwHvcgDDSc3FQC
SDwyHX4pZO0V6DxkaCFsxTZXA36bZG9CFuy9O/Dn6xfzmvuWLPwPHt7Noh4ZWVZJ
bfCXGv3eMN+LvMeHnKDu1QDRBft/pEOvQBe37yYmRvFg4+9VkkDTZwDd+Z1aippq
xxKO5J+V77T3POvPzLQRVoYqh4C4ec8mZsxZj90AazhTutJzWJBCJoMgVgMXBi3X
k/gKXeV9poJR2DcRNxeIN8PDD0sr8Bd6Lgta5/l7VWYFIA8//oK1JR0rlyl51wn6
VO5dJMv5GqOYnyuPfsLrYw+VL7tGYHGX2taG9k+P1psffICu1HfBkL051p1OfBZy
OiR9JH9afy4lokp8BxyYj/dNdWFC3PvUqfvVp9Rsq36gNIPwYIBU2kNhjbIrgQme
aG5JOswlK4jJEXGWiIZ3JRLUn5raQwhYz2USPWDONJpC5F+AtyuxK/T9vDNKeFIi
rT76JRbu9fbFbl/Qn+4XROxa8QFkeE9uIaEBmP64pkkN0Wmk5CBrDvVIxe7P+cQr
Dqs8dD4LGG0XQV7wf9LJrhIYvYz9+cg9fmqTXY5SXl4eLIAlHNA4q4MSujOEN7nS
OLbn83knW0Ls81o/Vf1Scm0En7WRV1XWUlKV8YK1zTWjDADw7wFm5KlGlf2FyLhL
y/yNQv5HUU0+Lxg9H3M0lH3ejQvcQXNxSFTlAU6Vsy5dtkl1U+7Ys7wyWg7NSaxt
BXgxH1sgyCFp4DY+awOxg7qgeg0ovk3spa+CsXnxm55Ci6rdEkRGewBvfs5ekou2
gwr4QYWGojjK4ueMecCaWUAieRRArHAwczC9FOJWwZjQObCBULH4qk881aRvLxS7
MDWn2TaDb7Njez8+wXkE6noakKLBXyL03M4X7oX5IjbyLSXFUAI/umxvDk1w8UTD
EVdZ+c8zikL1IQuWlwFS3rs2KjiRTyod2X4fkXit80ejNaN2Pb2hIne9N8IlPmdg
EvTjOHRBD1cFb08dZ0BWtwPiW+MI6g69ADx/08AqHog/0hVQmdvCxlQihkVZE5QF
PMYd2AAMpKIZ+x4fMftEf8GbZhEgkdiU1olmIrn36LL3t35t3X2aUD/kLkLtY79n
SuS2sKb9R7ZYWLxzvNUDrbR0UZ1RG4VxK1WHrX9gBr4g13E78vS9UE1McOZQZFb6
IubRJUpSnI2tcxnY1Bjv/WTGUj5yQraR35txXxkHfcr6fvotZh4n6j8u7piQldX2
ZYyFXnZvtbwKTr87iPJgWQzfyj8Kt0lPkz6sKolQ+9c+LdioDGk65fgAkabbWr8U
4He28GVpTjEK27IhdiAwYDaR+xYGJqAuutbWZot2FM7XoHac2bNSwrP6B6Q5/l0J
igTV4BTQlq42ftZWhBk6lcwX/Vh2iAKm55mImx2zZeWgNj6a+i3x5TYpzz9dJu4W
7MaNyytwcZeXc+qzLcMgLO5AGIdzmqSLQFZaEK+ypJIMs7aTUBzoey9Tf3LCJFOU
tALe38lzbcnUV12ui/1UYkF9Em/B4sb7I+hOCueltYqpqcZudp9A1/Jt4g4CqUvy
Wl1HcVhgdWOBOPRPprXG6gVls+e7nV3c8pi3sr2v7p2bAk/84rFChRKVsQeYrSRj
ejld/+P0CHVPgk41/7ThM3VRXomE3lsCoEjs0gcPWodK3WHkM2fpr6+jxJLkcAa0
WDiSoCBefiV3ZBjheYyWkNsRNLag1l2UhxiL/hoRcWl4U6JdCa6HQ8GQuIxpCC0H
LHg10aacqgV4T9OhTQMyH7GSwGAN+QAck3NXXsulyxEJ0NNABVS4UFeoO2kTKV9g
h1Dz9jOwT5H5K3EGhZIzeVGqQm8pnQzEJg/mDwobNHV6p6j2uqPnMT6TpNqXosT+
0OyJUx3yStIuDANeR6vcmxzorokZ+TVraaFVNR5BN89zGOTppfwc5ERoyuCnbr73
7ihzuKVb0vHckggfXdTkSliYlRV6LQPz0nL53lXPpuFEzZeJjBfVymIquWOj9HP8
ulOoi9TF+u4KPSdvzlbbxOV2Cx5RUom+DCnW6S8UTWp+jFsk8Dwq0Da0qK3039Fs
MJwbqL3/+Q4hDjl3vTLyuWKDfd2IbIGCeh6L/M5O7YuM2O7DY+zrIEUPWqA7jxjB
rqc/VzSfJoIhtyh1WRCLqeAGAkQ3q2i5mCCsRFOqesxDEVawdR45AknZhJyE1afL
LoRSoNmFVyQi02yywwxfhIO8t0ZjIe4GE7mI/Nj/ZNcJ3dlJSgsvy7bwYbvczPK9
nDaPjM289zSDvM1zJxoc/xgYfENtLF/MDQ49BI8+zcaEVbfibdSm4JTL3npgRDDv
lMmlRE7K1EPE/1fINq/9VPJpitP9rHmcfs8W0x+FVuDN/em1R6DSCzApVrxUPb9U
IwdLeIHV2T3thpQ3XfornmcY5U6KpbDEmeT2ukn5saZsvEp/qPnipFksSx1pQMAV
jjWSqQ6m8/gQWTEpPaWg54nNa19zpZvbrtpGf2Jg3JpAeiMXwXYsqa1rpmxuDfLT
UQPP3mZzvumljX7aYDzQO6NeY0KTG8njHY06FPY0T+oEjAyuBOXKJm18Uu2vBwOo
9eBUDHU+F5IIyxDPLrW0E+PtNi66OlgJi51yzw8HuHRsl1awoqrQ7vkCRj/hX3fE
73TDZkID3epCgL39jyZlga9tD5g5Dkvn4SMJESkUAytHURqvflpeiQGbA9WdiwP9
uMUQCGJhG4UALhEpbatK7bWAM09jG8ULTG/DAZasmP48mrvHR+CYvSXhtJN/d55p
LFQJ76ULushfr4ab50BtdplU0OMkWlyeitNPfRUzQ7CZv0v0APHmU4TL6iyeHeV8
YlQ1Mo+8xXsp7oBIkpnNsj8j3HueJP8d24iBnDVm2GdMZrXER33pn/YGY58Zn6Yb
F/HKdOR9u+2vzCmqtbhX9/KzWYYcZzPeyMms+cqvYgzlb0jXLxJY/kVEWlRzs40Z
W1ddVvZ/2NWoGBBIBF/oQyv9xvGVupkzV2boYockItjNX0k+ETtKseeqqy3wNHf/
uEr9dSgjzQgsmgBKGfQDUizyyxb8tPuZAlrJHYhY4lumUGMxxO/jzd8tomDAxQWV
3snGMQY+zBQOlJaZutDIwtZvfOYF9WqFmdMEf0XgJFP++Ezq88RDjoWlDzVrWkE2
qDjGnzQRkQ5eAoVv1lDWp0hoM4g9yTPCH/lxVAFuZS5fDbqxKTY9KRo6hljVTnle
bYDdfIMqTKzR7i28w+o7UUOvSZOcc4zC4TxSrTttKeNef0y9rldISvVU/MqerLcR
US2pjh/gK3g51L4HGgadkf6pvqBnJTdbkqsB12sETDXr8DIeQd4Q6dW2ycYKHcGB
wRResvDVxWNs1EqKAxgRlegTnff9DrMxg6rF9iriKlPICAQYfTYWIAs3oZXXMipQ
vTgJzg6dZPdwj0/CuFU9irI7D8FbOIV/uVgnyhjj1/cTIXtx1OGMQirT8txjhSsR
zUP/GpQlIdaMahueU1p8t0bx//GuwGDDrn3744y/IFWunPGpWlS3ZMbigJC6mOy1
tmtD/LdbpKTolGmdWGaevbO6DEkTJPQ/MXU4rk/StNNeta2BU+lI+mvTzzIReyKg
7PWmSZXqElLTGkqY4gCExdE/CZVP7nTfRhsZ129yOsvsjz8gOkDaaEY9ElXwJOxI
w3AbzULDqxTSv98r1HnvkHr2bYqoGwsupxd7I8pTLVZh1wnHxjDFaoIrf5xxk1sz
Co/OwPXEBubCP3uOwwPka6Oyaos0LFxmtut7v8rF2A6LIXT1oEYsWlzI/d0uOvzr
8+Gr/Glb5OQCe6PBpyE41P8kd4HA5GME7cvx9fM6NQKK293r70Vu7KevtV5Xs6zO
2m5mqeEbQ+OpTuUCrMc4AMLL0lvCap+E6ctM9PJ0mVNPiWkCSy+ybdym4SpOxBxk
M2Xw3+iuK6wBuv5mammnWvpz3QSe4IrXibg/RVr6W++y+CoaCizQHsjrjkFt11XZ
9nZUVKEH+bcbwa8+3ZP/sezrQilJn845pCFVsBfMdvQROc+lFOJS9ybq37r97RHL
t2DKXsxKyeBEGMYBps9yWortZSfhset+E7r13/C8i8Pe8rrOxAOTWdI62VkW1Jqy
diF/Yp5e2+rMSuiCuUhc9Hk1pivI+hfIi553JYTwd7k6Ik0GMkV6m0WYN1cJ3Xsp
KF8wPLbYUZaOdPjKiDH4H6KadivaqtWK38O9ni7SQqRljMUeKQv1uBq0SPuQSjzu
F9Gzep59z9KZxOS5iy9N7ivwswq5U/i/Qs4N9/rdxOwLURqYXf6crhw/KiZC2G75
mAYjJp3yjcVepg9bWuCHmtebJpFSyxt9tBmGAoofyDxuzuYG5nYv6FvQw40H/xyy
nyo8s32pHx9uZr2FCq2jvzmPL//2GdaZ2c74KC4S+xZ5i9xrdPMCoEiRdnDY+BZk
2CUniY1V7zyJNkgv+AqPOyJ0G4zsdTxZwESKmDfcwi/Jghy782JGQNbIG/soKNWn
ucFbJVPqAqY3hsWDFbdxVYeVH4S9Y3TJyeStVCTm+r5NyuZEg6XK0dT8iENa7exO
Z336Zw6BazCzC2rqeBz5eg+AkeEKrxT4vtyPd042ldzhWIATxMz5gBBlCYeiR/nt
kry/HBpBMEz4VUORBZ/q4w45MXBvGieZjv5SYr64qRdEBYwGI5ITMNISq9rjhjTc
GZnVDXzKakFPV6XO7nq/MiqRufajhCT24vnaHrwh9XtUb+zNXuP69EWTIdxt009F
RozYW/31XOCXESVrDG15hlopnF1+N6XiTaBSRYL5zieCS2mMtuQGAKkHQFMk9wPw
ufYkfff8YiuNCfkY3P5SL/5jvL4o+GQNlAi4URJjZRoIuRYjh9gdOxmNTKLn19i/
nPtLegWMtnmz5DBahDkk2JMluaZRSEC4z5fz9cXkOUjj/Bt1qhFKSWYUBX1PpaW2
xbAjNVrTN6702bNy83GGZocX8INu/mHKFEJLQeNyUtXys4z4qaxttsL6kBOVuVbe
1WK7PVXGtYFMafjSLqoHBqbTpgOvO4TD7OjwXABhhyjdxzKJ1aa3spPdJzb181iK
6UIWVJwSpVU0lk0D5MqAylWsRB96E6quu4lTuOeN2fr/WxV6FdInhTHtXCTla9Qq
LFt7/okApd9v5EGKVHqFsOxdQLj/Emp4CmYfv8fPwIvuvG1DcIHA6Frdc7n9qUMw
ZQSpQpWSInRT3td2aCmNVax6yVPbbLNDzoOFvVgXLCZNRIohOEyUh3/DaknW1Ltn
tERf/sT3DtLsUfbhmzNDYar0ObD6CjVgAKNapYizqlIvTIdhqKLAj2DL0yO1Mv8n
pAvVnLs8aCXgklxUoXHPbMGZlivUFInE9Wb+jU/M5rpcb/7rr1Qkb9nXuOqbAxWo
aWFg4uemJbq99IskZNaINbhTiZpLoG9J+s+7DArHqfE0V6Of5zGJRz76Epdx2KOD
sVkMfCGBHvoMJPYHwpbYarzK9dFkvFtQqLn/vn7WA+/w31kpmpQMEIep/LKV6Ooy
TYro/w6LbN8Q9Vv9L2ug8ti/AmglWy4gLLLareAXSE/439lWvki2ugiFaTcj1bbC
x/2HlXgYOElfFSC1Pffa1P/CEj+gg87i9ZnvO2NToMuEdH/Gu/sD3jjo4w2Ngw4R
l+30uNKHonPckFpCTU5xIhIsbeNnDBR7OzXYXJ+/kpA15I/HtLZzO/eWhCzLQ78r
mC0o346hHvRJFJuM//wik3A3IA0bhJ9mjZ2f99g4wbuDexQUPHOWhgWtPRHotFWU
RqStRUH9jugLI7PZlewslrAKs16gGfo5FJuyvNh7I1lL4pAastf8j4YqmeYqTb5e
DBxeTRmKNCkZ165blZR5Cmakjynld+LRAca2lHgopW7xOxPprdJHj6tKJxXYiYqk
pCY1QCSgHayDH62We1ntPj7LUcf8vdOmHyfzWz1TEgnJjtemTP0HxIaLyuUYrLgP
OnOYPWj0OK4VT8bnMZT5YPPR98IzBdy8nySvflZZe9PqoOs57saOclHDGEr4QUNA
2ypOo0VXjQljOzULeHHtiQEoiL6CPgsfkdaIv03MBprHWzG+ZqCYPyCTAOut0ADB
GT9JmmdSUgyDHFhHiegVa849jkMqFIDiT2xaLf0AF4XdAyl5dkjsqxv/8IJGua8R
e6Yv2edssWpyPxz4qr3/+0mDL67pha4WX63faLm9KakLJFqoyk3p+7PHsuSHuq2S
Vb83Z91SZCl0TH5h5hAQKENUi+/G67lhkda62g0bTAWDzqjo85Bhkb+IT/5PPHld
0tmNCHchdPVBjLBLnCSvpTh0XAVpo4Ev5CAVIgQgWQf9iRoCt9iNjIbsZHXtSeM3
E5qNOJKBHX6qXMoaIjVFVENH53l1OjwquVmixzB/Wikc5Ldp8HHy0Ao/NOAGbaGb
6N2SasjQFKPLQOHRSO/bsRbF7OXLc5xLPr9x7WWAlSdm3OOWleXf1dwkozUCrvPp
FwovHfnJ5ikA9xms+3NYKWvuXJk3VfuMeA8hWz89aH1adAy/49sDEC5QQ7weXxkJ
O49yXZSUcGJz1121CR8RhGx93gCWUH5Fg7EUx3KrgAp2r7KylNgxn9+MZCUq3vyM
YPG87ueKrNywII/WhMNuzYr24QWOb0GWBiH59PNyLXtzSE6Kr4pzi9opknS/LvV8
jl1WAp+dZTlu0fvRFSYzqX5fOhJztBy5OTRzn9ZSrPD34JHu1yPiCt6Xozzf1V9n
su/M9lc9qDDdkp9/Goal+LAeT8hLVCpyYKr5RiZZ9IK8F8xq6zVVyma2t5vRc1d7
7bUvyIrLGbJkGuRICBO4e9eXSXocS6zioy3IO9HXDi1gEx9f7QVOLp9OdxdiVISw
jUSb6LOZCgZyXoUYk8la3/1WWqog/nCInvpk20/ND7KJ1B8p+So79XovQhFdWqa+
yMucvC2V25Gp2d1hFupxrOozWNhTHMfWMT55LDtSpl4OvRFQs7TrtxcuMMvjl+z+
6IeL7oJKuIB9EaFll7iZQbziwOJx65LmtKernmeLvnxO44N93KwcPWlk6B/Sm2cz
d57/wPbzfjtlMESALWfVvmWZMGHUGeqP71p3GxHgdEH4MWNUSvo5Qx7QBOFwOk/3
TV0eF2Dn38KpOwkuR8sZT7m8z1RA+9T8neYNhV+VHKEeYSiXy32p6n9FQ8aUWoyP
2GwJB2ZRkrijKctzeGgw6NP9fzWobZ9cuAYtsSdtotpBsHYoHUIqmcEeeICmImbo
X88uHrnDXSz+Ijs2bbMrhhz5vY18Ikkbp41sUpcYqOaT9ML7HzWG37W1MHfed9X5
nSDefvPiU1lIpOh2klLVH7Ijps4RVtRMnJXI2sPyMB5h/HU+Jx5TGkVV6M5Jit1V
ZtwPVRk/7rTPUMQTpT6VoZRoeDtm+OOCEeiR626b4B5skhCW7PkKriHs3UlLDQO/
U6tncxrlCGYrjGIiH2J9KpoWkZ+v3hGEpNunhpkwHRi8N9940u8CeBiEhtrNQH09
KAHe//un70HIIkrb+mVhUSJGZqFbI4ngDtupsfgMazCNkRiN8mxxHbPX2aBRxo4p
o9PNzRJoBR9C+ee7LvxYJDS8APrfTDbHacX9La2kd8TsD788j9mibxTjU0xN2JD/
yHaRgc5aYhjnXy1JohznCP4+OEh8hH6f7+7NbtF70zXIe6dJDMQXvLJrdQ+Utup1
HBvSwDDI6Xb+SpxIoWxPv9YjyGkfiU1JOf6M8QDzo+BNwKHU0+oLnqiBRb9A9eE0
eRFct2eOHM0X2tHRCUkwSNXgrErM/G74WrwXyp7i+9I3WzQWvt4cXw28FBHaGe2L
oBTWw2eAA5hdN2hkDCBTGsR0zORaeo7s4LX7kIWzGYdzpv7jtEYA+ntXuz8VB0Th
rxRNK8LBqDvSXqFNu159MtLewUW8wVLz1wUUhSuPoKh2ufQzLeGTSkfzDUJNOMap
dDDzpIt1KzHlNaPGsQ8aYqxuqMCZfh25nk8A0l18y7Wc2adNq7k90yMuzkOjND18
gC4Qzb/X5YvRjmlJ9umpWgLonxAUtLtm6TU2qnbnNgZ3GBZ/vzjETvvZfv4+Mc+j
NAMv+ypKjMD+hT7ruhpcs4tJlAAAO9wvushsr67ui9FYlroRoinRl+P6XWn8oLY6
rz+b8PyQzaeFMHckWtF1U1X5VsX8j0em+fbSoqy00bS4XroVwYwNNix/Pl9O5Pyt
fC5FfqE8C4b9YfVA6D+AmOKStUwcHW7tTra/rWz3dhf0jdLdv+SfQkfPzVZuWFRJ
IA5s/w+EOZadV1qorRk+2uWo4Rk71eK0MR17ToiLpBSvcrL4opqJUjI6HcXJiRL6
uqMnuWOBteF30RRg2aE7RZh/8blQv3EMDYy4eLaCiTeE/LgIdkEmWj3GJ9CHhUrm
MwA32nR0Nasq5DSq301bKroIQQQVNFnH9bWV5/CRiJk28khN+qlTeKX0NxSgIeNp
rnHlDu+RzyaFLpwsTeVnJnyDh8MhSxhKLq1EZdBJVaUw/o2DUpyaXYsB4NtoV3y9
XtTT+sdebxLmnBmXqmvNZORbxa5Tc9AM0E20ePWSKHEUBEZFfsOcfRQlV4aVISVf
tSBb8r3Da58TGhmoPOpC/MhDdmHPB/OFJA/zAzC8RmCK8lZVKfKDG7kc9JAZ/fXR
UHGMNVJv5ompjOXe76PyG7XOhQZ8wHnSP4KXl/QjMi+2iJ8fLoECHyo0iC+9kHUg
kuYRIChIIJZdy9fe/ElqnQQAzpb/4mJqzi089XhBGiWrCFHAfVGbzc35roqfNPP4
Orx62eLi1U4SLm1cPPb5BjyD5Cebwcd4+SvQtP56WdU8/LtaCKuYmvaxTrRFfp4I
nzkX38fF+1tMiZ5Hww6WCBCGwrjY6PqtTX5NTOeZ31xDent3QZhBoiuWstDZ1NG8
9spOOnd+RLCyYdKyViKPrHWYAkZB55JXFlJBtwB+vsDvdamwbebYnzK3OZsNR+gg
QIviQ0lfSRN3sEXFL7mBsT73gZHF3f1zdfezXPqwNehcFG3sbwpVY6KQWjs8Ga4P
7mLBB3PTDNN08+ocBjd4mn91kMKtGqELpCaOfqUcqUZ3r6hLKLiqrH6OK3+trAA9
s77VTOkznaPW1o9HF9t8GrT1UWWEp+2xeKonGRRL+7RRrj9fpa5fXAPrIvOgn45l
0V6A6d8yhwsjKirT81/1vrwkV1UUB334pY9FRbSNSGy99CUPnRqLdAAFfX+CCqNe
3xG96IJfFDJYj8lfN5T7EKUU7uccKH82E6ZJy8xDSIJRl194uVIDvSVes8wUoqGt
MwLxhvjpWasC6dMGyEdalfF7kEopBSFv4lyNw1fj5xBVHIPZb+5G4db3onrT7s0U
UGCTuxCnavbefd8jJIrNqVW+FirjAN1mtg7sM5yHbprQ0gMAiLK3aOmCCNvdmS5w
i+YDQAQxPMJh2pw67DTM5v1pyC+1eNzSOyxCR3MSXXLZeXyPcj9J80z+eZ3M7UuV
8Od9HoVwemmzdhxDULnNmD1XxYBog82Cfpl8I30xOtVXq1mXd5TzZsIr6Ud+KDQc
ZmD5yAQZcgCOFnPvIVOoafFOPdtVjoTn0C/ap/8REtE1/99+Pnu/qVJY4Yy/0gWG
MJBor+7H8c+0gPByY+xlVqoNCBUlw7vy7Gc7sb4xjJ95X704XhX6ZxX3GopcscRw
VE6baHSYCNrBqeNSrCJ8K4Ed35qoTt/zGm+rAIZNiCtmIMFhP3hjprPrWeH+pga9
Jnf0HtyGwuNnImYcIVG/V1iZjeCn+f76w0ziXiT/XLTLic3dJ0hllJtgjokPNaqD
tNQU5maezUntVyZwzqaRFBrg6ZEkJam+DNrTWG6lpboe+W1Q5t0DGZcee3zpjYfa
8Yn3mfU/Y+ggOgwyhnrFSgT6yRUVSS4wYozravGhgkzdtbk48Ok31klyUZG0PD0v
ToFDVZtj9xvToG65sz/lHTTEJbM+Fw7aNtpKNZcIoEAfG4euuLzCTABZZ3KvzAKv
581qRfrMSXdnOJNtIlE+xxL5dXWJVwyIwgf7O4VJ78KZvBq7AqLYsV/IX1itjy2x
H5Jp2sEbqsk3THfcUj3PKgHW+vnrcVOSYmj8/1Vk0Q+R2rZZIowwrHYzpfdGsNhS
eT4vmN/YBznL0GU5oHmMz/alNpyN1iMfIK5awLPyUEb4E2eIggxASmTn1B94SA5/
yoW2OgA1E9YRcPGHqczTOSTWI00dGjn+TVAyVZB8DGC/tesghcdY/Y++M4yw78v0
B7tA4avezsTvJwnY0J6sXxBuhyNY7+GOTsnPcRt0HYz2ftbyixtndn+CWorHYEpS
PWKGj9SgMVlHWOtmA3zcYb8ONkx/LeHvJq1NBfHjaLM6sgKGfflKtG5kh31TSBL+
dW2J5O5PjKatpRBjA6OsyDekCjIk0dZ8VLz207nAqTWpT6/TijN/MoiVJESbFdyB
mQWcGLXtSlDJ1b5ORzAAMolZX0HOWTH7wsEMVJrXxwfXH03Ph+zg56X4+AILk8LU
qeqWX5KZH1jxDlul3woGmg81x2oXrdzDrJjV+AtrEBO2PO1TV/3vGZKoGqcFIJdM
YbdE8yc/dhlwjBkNKvD5fPhPxyZH4ROmYba2nyo7jhwEsFpqPiQgNBhFjmrdrFe5
BmB3WaDz4XH45aVRxg1Dydfv6oXqTuIpBqxy45FTtsojAR6P+rp7mArkWkx+W5B4
NzoAaG3PEikvpUF96z0sRfJdyelfK+1ItjC7/vg1V/QcxdGrpf+tvoLsT3/8xIeL
4KyLGliAUvL40Nf1qKfqO3rTHgZTHzm0DtMSHT10IDKufRtMTKep//ZA/nIKjeAb
Gah31gAQi1ewYKvKaql2iVTueHtPO98GJps9LrolfIasAf6GukQBmJaY0/4X84o5
4FEUEqF67DMEXfTW5Ud3JnVomEJi3sNJNdoQ8O4cYWFs8sBwDaNEnltZIJXSjxhu
JmwYjkQiSeB07wYe/VlszBv4DHlpmVIMNLFE2I36sIveA0oomk26mz3Z3E2vgyQa
FWMl3A1r9dwjPHyfLIZzc4vCJDppa1TkmgQaThfzA7MeY1aIiAL4FCMKmcExDOUo
Q3b5Ga0je5xQVlxKvaa8245w3g3iyx5uRRWzXUNx+Z6FkUw9F33S8Wqm//MBGyLq
svqtkU04QnOGBjY9U/d6flTNLM5DwV5LYlIk3j06WKN8Lari+7oR0RchGuoFbECj
CdDox6FWyPY5q6RoVZmDrguIMRz3P+JuQlW0RA6S7mQX0mrAav7rTuZ8kgoFJvKs
9II6VNBBJ9cgIweyuZ0ZI5Nq0LDnvEIVPN+B/3Zq5xSUY6Iy9nF1GBVetpKl41LL
ULVWSUud7Do7ppQvEU6km5h8TuTKZSKFQfDg5qiVdFZLd32Ol9Op3jyM/qBluOuQ
s5zw9ZYEBQZxK/OyfDLP0aN+lDHw8+RbgdjbQR4ArjO/OAVqieBOkDhZPkjoXroX
u0azR6hb82tF5wEebfooXBHF5cNfPpZNHSlyP4wDgect8O3+Ut+mOM57vFzY9tOt
r337GSgjQNYHqaWHhtTEXcYLBNQE4cS9+/WnTTNs4Z48NvJjaZ5E0m1g9us+Qi2n
ZHDt5YdYdoqpDVgVOf7NYNAiU+xOy/UhjrlhsAfoM+/P/3VC1fbbYBU2yN6M0Gps
8LjowBYvWjgXy+fqEbooPNo+pD/1ZyGTxXpxw+eDjBgPpSde92oiDJYgudM8Z0Jv
n7kB38TrFdjSjEHOleoIeRaL68JMTGVebN8KI6oWNXOwNikAqHnI8kRtyJF6JGef
UfpbPzOCfF+hLahDsgpPgcfTdvPK8lOXaclKfUcWOVsaudAGN3hkK/hVL6HzCUHg
hidaCQph7RvLac+dXq+EKDboJ0ht5HAhDtG7tb6sKOLV/bMyX2pDwWJf1eck5rKZ
4mwk2YGp59rq4H7G1oVsgOGT4ncQGbOi1hwQZsVYz2Kt/+tjgsO92Vb+hz5QmPJk
joyPUgoFi7ax3nRQ1UzVRSF36X4EwRtW9oUhVxwFRgX3EMSyKDcghcQZtbc+igNx
qX736G5x2RcWwgUuOmnDmm6lc05XayeEZir4JZZzdoOUKWlvSOTEMPKYLdgUDgyE
p4yGaFxQVHAXswzqMWiawUw4PYFTi+jTz4nqAZGTAsGyPVQ9s5bwVRu6DUxc1vVT
jRHR1/nNGd7Ptm5zuibGkd0HA9EMBGHcqINKUXz8pVl7Hqx/ZHuAJ2FvJ9nY+JZg
ceN+Oo6bALKL4OZWCSmUtVzVKatJSb98gTSKG3cS4muXJLCkp373gRQl+487ECmy
0RJs8g2LVVPEeRQcqr4ClBPa1H9aF71QU9aA0oLiFkZy+7RofbEwtRqiLO1881gB
Ro8jyVxjAtKA4STaHp09KHZdByQlGuUamePfD0BJKRo87gYvTcW5nWa8jV4TEVhI
3ceUKrCIkC4CPLm0F63DP9I51jN2mc1r8rHzzOuTbGAGYNaHvjbCSATOqYrO1WgU
mQu9CiyIEg389D5ZZf2zSXBuUu2HrWv0zzuIysHYiEpXGwwKZhfFgMUZxEdROQgH
fkCzEkwhecmA1Ccyau9Xa2fl7SaCpoeRx+Yb7LGfHkEWylyeSQlmQw0AXObEkbrb
hh6Q3TgkQr0ths8cUhRlIqC2Jtovt6kl9myPs+FDpQUvKNC69BYy2HDrcHpwe877
IonWpTDKdmFjWsM7VvxHE3bO9tuWuM0F/3TfeRwMn0b8PJPKkKabuuO7KsV9oOhJ
mAuzoEsvjf13sTTf3jtBGPGuOOdTnp0qNd61CHD2Jf7QXvohPYPeN2P2GajpjGSr
+2wlnxNUDRfabZn3XccTP3IfwcNTELbXrIESPdA0tcarV9gZAaIUpwbtzfV5ufsP
QlWB09Oe0A+mRCfJ8sG/hX/Luz2ONxlqO1zMT8ThDocMeUURIuOgZhDcd1/EMx13
6AYBaJBzh956UJxPPtBjX1xdmTXL30Dx7/Yawwav/zkBjqmW2l2M7Vbjcrqd3K9y
wV/kKBSYbRFaCkfiPP+iqGKpSxFdlDWETeCnm8dYKWwE9/Y6EmB0dmnycZ01BWSi
b2WKZ63e6SdCJRC7jTxxjiC+t6VbcecIyUcnb6plPdDQ3hXaRA+PFGQhJR/lekiV
OKcjs3FJpPMcI7o7yFrqJJeTT4s+5agbRtfDbxYFsRr1zS1eNMwjlxdUruFWkpfs
6g1f9wzaFisrowE6C/0LL6f6v4o7dHFDb71Pl+rjTXW6vBwXk3+yZ3t5D2pPWgOT
n7VozN2F4uBDq4KlR7cMHT1Ps8PV+LOwOIGaUlcKyFaaGnr0WiePt+PnzYr6A+Hn
pleshXtILc6xsM4U4lTczypjYSskn1Hf76bNU2PyPTbfEtOOcmNDDVmFN8hUIHae
gDRb9R0HWamUbRHRMbvXxW2bHVix/kVeV4C5qKaDMrswvtdwO2SyQeiV99oBU6kI
paiKR3JCGTMEt3x7QBeQKzoEk6n2HP3qnoGBTHlgje+6mq7VPNqRg0FmZTJAtJE/
W8YmWjNcrp7r0LwLT3jNsZSx8zgsq5jxBYMvFjAdYivtF3EtyGqJHiRBJiyYJWtd
M4OMsC3hrziohoTPlLfBSCUGcQC/r3UfjbYM1r19Fbr4tUDo7D/bitrSK5talKia
A9U/3cxHSJh7PWr50sLs3sVbSVCJlOZkH+boqpiDGs6iFO/amGNEhwfYzQ464SPn
PMOoo7CzgxAamati4sqcq54J0xSdDZF2Mch31b/U/YHQ5wcR7hJ27pDnudozAtvo
2fVRQdYSudQxY9Afxlc/AgKAKRsB1l9qEUQ+X/QMelQ9i9c1rGFkG7EIh9HRjXXm
j2ATR5Wq71LGgZSk9Zvw/E+im/x4sepUztgYw+gP5EBJUsxRQWOh0ntKocLekjL2
dCJDW4tvB45DQ4N1lJBMQxMvltlBymtXRrr8fw8u6hz6Qqip1zQBlamL32X3RV04
WVBzGE5FGiVPR+/q/CYtYGxXMGnleaC0DdilbCGG1DcQmojjejsHXO8tRDRbscB8
ZYxW23U/7hCQVtdVAQbSWHBTlndzOG88pSxwrV/f+YpRgnWpZMixgnljmuhgerir
wAs+lQMcLQFNlEscG9Hsh4Clc+a2LDpOxrO6TgF2kAv+q0W5pddK18O3FsY5XZ6P
1kCgB1QgRst7bBpUM0UdRjlWLz2alb4ggjLRcTidxZylxKgTAFAz5n6wkBSaO2A1
fWh+C/yd+Ndd0yp+niExi0fBa+RtblsUKjNz1X8qDMkhuvlIFunLCAxUgpfSiHnc
/p7Z5LBAm+Zh8vnq/85yzzZNaC1GF+jBOe1v+A1nByt9uQPh96RlKq+WkkR0LIyb
AN4mB46UTlN9ciJDIvBfnV7xK79Mqp89eXyhoRtUJUDJ0CM4/fdtS5NADKHgUH2R
5UuluTDIoLyxQL2L19LiSSv/ionBGf6yw0zGhRE8apYG57euiFLbHzHslLKc4aOj
H0EO+bGtzWJAUjE9aSzFXVxj4Phx6kyBMiCYWbPUW/45zEn1tGNV2e5bJy2zXaYE
a9jH2K2L0vj3BZWZKN3yMX5jsres0KwkI62ipxhrpQq/lgyDhk/Bj4w2qOl7DQY3
sAmu6vqkIt0BER6p0KNXrqoA3jxusjByPGmNMxPv8zrgVCtcz89iSJgRwMasnb0z
Wt+wCr3sFaU75MlvU4qKXE5MjkDhq3XcHU42oMgTnSZ8rRxJQuiBiGLA0LH5tHrF
l/FqQGVhxZ03t41H5mKSUtocfMBgSnk9mRxg4mvlTQ5rObq3jfE+bFXwsUs9CMfx
U1I8ed3J3QSALy8SZEPGmtQcZGEvSRkgl3hONq6MABRcnyOt6n5FQTTxWWQSypkd
h/67Y8sEqa/6KuegRmT/pdG/2KfeO9yne0b4F1io/f+bQAqmLKygPY5rf4omcSQj
0ABpADdPGwdp/wPX3cZ8Q9ge1vqSpG5pkUPRTgwYV4Ne0QNCX7bHDS2fdMzkS9JJ
J08QlCVoD/+t9ICRNuYLcLvrLWQ/Ol+johEvOgG2QjLupzMsBKJYkUjNCCOnyzvf
eaH6nTiPNSO+wA9Oj9PlTuXE0usk9v7G/eJ53n/JWfkbx8dUns+FZ3WQBvWF4g82
WOqTPAGDicpJPg01nj1D6rcS9pB1p0CzkGf4ipgzxpt56gGTJ2k94rH10mMx7NWI
PJGng25Xiu5L9XVvNGkUSIqQ6C6BTlkCFdj80MVkUi3AhgcZrvuFOzBSeGt1dEUU
zQSLawYgLycAS9WJzfpwvYtRsbUmToXoXedSspDkD85eW8+JLgpQeXq+7pjRyrYE
hukECn/js67TcTDJYEeWFCaDu6K1L03mrbnaUC/cGL/KLoFKMKucfrGEINaLf7eR
E4HJgTZJP6Mrt2m7xmiLpShZWDPHGzh4488aK9FKJCrOkycb9dA71d+k5PrW4h7B
KjCou0cHIWe1uoTxtVRiVi0k50n9DRPzI6Ca+LoJDVJmSNvhXU/x0q6/O6cceRgR
DwBvowQH7U2gydj7/y1teGjvy6X/j7flspSZ0ZJGuxMpi4wAsRcDoo6V2o1BIRa/
7XoPXwWTwGobZXbKwkX4bYs18blh+51Ux1Mxt+vkhHJZxPrEWVvJY42QeMMzviFx
O93HV1JWfnm6t2pq5qFtCMRTL9HDiPmYls/rTfB8nVo2WYD27tWOdo1GCReoIzrO
JArkkPfDEgR1lMCw+I7zeS2novEHA3QVAqtA60R4wrTTpPtU3IeLwUKxEVR4fo7H
yQJWxmQUxdGQ7Ncfpmwwvek1EgdqbA+I/T8zU+AndQRjB+8pomF/NxtPJH4Fewn2
Qvkw6osqZvhq8O4UngHxoCqsZxoMZHe7w9OH6yqeMrLW3yppcEysWYJolb9Dl/Ae
1Kkf0aJzLNAJRupsozEMhBwXK6d8Vw9/an33p9wKx/NJzVNQOgMlbNNuk0EEVj74
YLSDTT9FmQL3Bd5iiejPizA6NiCWZ7EHABnHfevG6Vo+DegfrsgZGAfxS/oBDR64
7egdygaoAzchQ8Qsbq9n/c8+FoziG8MhayjdckcmecdAWQ4E9nSy8SyzFQUkB9Di
y17IMu8tP6urjsd+OX6pjmYjvaTA685+sB/B+3XedkT0a1btmZfGqZR7BQM8CZpC
u4ez+WeyBdbCjidOyCcj2nLFvRa3JbGRWD9CHqfZTtXbMnI5g4v1mIto/ktSDKiv
+ovs9v5KMLmI7m/wL3C1uMeHr3QD8pvGwLRFweZUvxzzKg9ctDtx6S0iY6pY4qS4
XPer7CSJmchXbSnxJqopwHvR610uzqF43UgFCk2eThg4D8lTlvYCNstsgvHkl0n/
N0MZN05gbmPZnAhDArNBFHwUpkKPrio4ATYM8ovOoQ/+d58dmTVl1PFVUaJ08g1f
SlNLhL4U35GuKpEFK4sYPZtpTaFjZQOLQl5CbP22ZGykIOPUIFloC3AL0xbYhdRF
TP48HkxcRvamuJI5ODGc3knbaddQTM6zXCYTSjsf6w1poqIV04NiubFt4EC4svwb
O1X2Gzdf3z5qvpPVweeiRK/+V1oa61vKgyiDS7oTNFuJjiepGbNYvdtSgq0zDCFY
+jU41v6p22dm8XlDrN84jidkvBeTPqCT7DncgZlNBQaG/6vFTAK85N3m7NnwlQ7x
C1l6AXJzsE8F5o7dFJUtaXj3Pd6QKF7bdmvRh+JCTy4ncumnySdTdstQg6K41Kfx
M9brzG302Llg/J75IUU6P0Cosr7S8ZX4/8g5It5WHjLUgKvehQFb5lDgAaLs4Hrz
xGVEfwhq5/LCSBB2f2PFtgJwkBeiWucKMsxpU9TR+3GUsmHyn1y0xGZxW2D3wI/R
BqsGfly7YAn2iws9ZtvoCfqMHe901PjLqGE0JIJ9q/BC+CvA/NNtkTpyn1S/pkO/
9CNpdAeEUjTobkY6/nP5mv9o6F7Kru/todi3THwlnKePl3QO7H7tNlPN1sXofewm
t3ECqpjIxn8Aphozc7QvreQ82FxBO9ziddgR4l2cOl8gF34AJdJAzz5O9J0zASvX
Nt+07FmRP5MA75BxJ7gIS9857UsqCmbWAeuDYxh40btVhUu07UK+LJuYJk9JQMV9
R8AT38JwKGx61YFGIOA63y8aZwR/fxAoJapEXANHDNtqIvnfh0jMSo/EFBeHqcYA
NRphZtGpXA0fSj+ONe2ZsFVbpBvQPzFDadaPco1Svx6x55hgCtsLOcD05KHmvXOj
ZznsknVbPLkO2GXfOu6+CFI5Vao61/MVjAk3azLm5YEUqhAuq2XrhI3n6vub7ZuZ
gGYKYVXFlzmRFIJrtLKt9VfqPcBYaRAEX8Tvajrx3JPp71mRGNgtQYxwFm1c+eFM
c1rmvGdZcUNZ81tZGEnsTRnpLRUnTEHGmQ7Shf0hiXxl63t/tuLVMvKuWZjhdh5P
ppW9qPIrmsLc5ds0y39R+p5YqZvRuQNoESP76nOH3vHzcWMn65s20yHEcbTMxfHZ
fanBTLfWRsw1gmgST/1OwaQogMcZDEljaPAOY/W3Q/heF1KG96fmC7TzGCEifUU1
ma6mbGdkyqY3JCBcNJjxa7LdDKmVnKmfee1XNN7aGFqm1POSWnorYP1lOKtTU2jM
DH6CISNs8msgMxtdyhTlqdzsln8jhiowcAhPi1+yIXXEyc+SgJFx2eJmutClwzNH
J9VeOJ+EIRPlUOqWYDYKeW/jrteTPMLREuXE6jBoLCvMZBIADOn1YhxdMbxTqJ9s
i9Egb9mGxlFqqyOI4ccowStX7XYyQvbY2l12F1VYOT49tbh/O9YHN+FEVHjw7AFh
9hslJkgSF2isg40aO8T94oJsQ2PdoQh7TynEsJaZzgWHCka8akgdzIsECjYIf5AM
b8E4MMpJKFNgvead1DCNNxnwkrK+T2Suymf/zA0Ayq0KRmfqA9PANlSTxbS+MKBj
u4MkE36RYS4QQw3FmQyWzD87ia/DIYE+H9BANZ6eE1wIi+v8Fi+L0WCgTweMdq7T
Hk2VA5KZ/CIRva+PtvmPpolPciTzJrTQ7b7FFzCp8/w1m9Hp2AfTQwg+iIGk7a1Q
2HzIfGmIr29qKYq4r3BGxt1v8R7ZvlLjSswpWDHcMHjtALqjDgNqiQnFhmpnr2Kd
ubpEgdH6XRJT7FJdDbRRcxhf1cjypxNk76/O2N4J0/Ooy9RdU75ImPJBIZ9ow37C
MpbImbVV+8xn4TPJNPJqPeqC/gKGH+jPn8CetmzCXeqx8LPGLrS0xb60Q4/FJsNm
kjrt2QdjrOGiQ6SoU6Xo0SZ/aDG7hcPbQWoyVnOsZf9pf4gZYZy9FPEYlcx93uR5
JqLq82OezlW2wppmvCOrlBILqyuSCjx5O0kuInw8GHAmYZpfyFqwV6CsB+drmfpI
iti5X3IvYPvCNpCUnSj8/tMy6R3OmjdeF8XfT9nvnE1YmByJZX+eaTKRdw9XZsbB
n34pKmHm/l3w86oOv+zkFwHn7RfoYsolFpx2fC2AzeIrbYmTX534IX0FzewsjoAr
d+gETj6SuKW14mcveQy1pIsRHre4DfSjxYWAH+fjMT/34e/grcUP59GZv25OAZ1V
stiFtaQngs48bosiG/sNZif5Tc1flZHc9RDXwe5DBpq7rI8v7+XmaM0m2XdHwQEE
TgxHI2HXSGNJWtDYcCBTroWqqtE9JrM3krhYBffa0cYK6l13qpOnBbp/p9CgFmzO
dYzNg3RwAa2tW2jMAIzMyNI+T7Kng/6/G9d5QOe9/+dMR/Y8GEQd4IW1L6Lnrjbt
kHHWOz8JhA5HrNbft9ZXJ+IPaiIERt4ee3o7wZPno7//hmugcgq1LUHMB6UQQ2V/
bxT+3DJj2HTlVrnohkQIEX96YZqSJBp03dXDDie+FXi02wr1GmSCrVTaPy4j8TqP
gm17sPhyBXUip4iGAMDtbrU1gvlwEhOELORoF4PkitJDsTvi57I1qSBNoumc495B
/rXrT92gyAEdvp1xMziXQ9TWS6yV2V4Ao40OdB6wKHfS8rcAwSYnDm3UveQiVJs4
8cD54/x/EDj38EeVSXZleBf/fDjCYZmsCh/gQiTbtpo0awLoW8Z5tJLHQNEbzeI3
dQfU2nhAy3rptYYYrM4dk55q1dEvi9Y9jV2VLq4ouWLliGuIU/rXGFHHt9awHxjk
3aXbuIRXiUH5zqSiKUXcFcqiBVmBMI3+qvlrR42UKcTln3ctal7oLRCvtL7zuy3C
ozyI+qtKnCivBXFziCDR5vHP5DVxrLtM2lJ1xvcFXMjX3zIo+jzgG6UWkgZzs5xa
+8HLUY2WJBb6vF5CNEXTrzfowpLpRmsCKVk7qUxGTWvx6xFSi78ypoqyjVCOmKWW
1uJmdf9j4CoYPRLOINQmvo2WCBhlCV8XVPag8W5yVvqf4nKoXOh3HYQjSkzLn1EV
FHFlebrfuBPvOTPBvmREoXaXfyChFhZpyLNk3qAUXdeccyP8pR4OdHFC56BcZmH0
J/7I5w82AdhfbY3lX+7G2xNuYiofSQhUJ0if44ZrF65n+nlq2G9pTKufTtAwVDcY
PTR86LXrq76/QN8x6TcgrSuS4FdhlGr/MI1fMmVi/Ubgo/It+3UJI2o8483TSkkt
sg70jOxA8y9SsKfXRzlzlrnnAN7c1J079lxFi1L0B4lwPZHB+y4WCsW32FTikN7l
P10+0MbCGsIzarCCnu4jLQmylQ7Rhj2zu6orZJd/9l3haQBOPY2kN/z9MqbvsKRx
UehYnpglRZkM3QJOcAkIVOR6SQLDgvn/8Ewu/NCmA+e9Xboy5DXLkH3K1CmRmBlT
1fLdeu1NPauW1sfkwPHKsuA1JguM+QxX3QgvTKE5KywMn6axXRFIbQl5Y7f57Eiv
ATmXQ/b/2VLbruxWsv5/PamU5fwo7XobyvO6Pd7bcmg4zL5USa/DF7MIvPrIPg1i
LAZTVPeLIDkjGwYrfgxlQHQRqR5xhcklmVJiiLAyCsqXhTfEtkJs1QH9r1rJ3QlW
5Cy94SsfTC4BOM4uRXmc/4Kb2YxRjnCN+uq9NtsOEB/L1fkJB9QtCaf6h2ZOhx37
baG3tx/2rXTvAVOKGTJl9XfabdpNzT3kFNSAEqLap/9kOYhzcCoxKTRf0xfhNx3f
jEvf7oed46EP/64E0Vziqg2slpidplJmDcK9mUgIEhjUldKgJC792wEFFYoEakqM
0Fz5Z4gZnC299E5+YdZ7J/14ZGcz2n5SSjEbaqtNux3MNmQ/F2M4kLiokzyM9eZh
PG4K1CaGGAUUxc9Tqff+eie1+lRKD9VWA/5Czk+LdPmnyHikzE2WsXIAX2oaN/Ig
kAicfmd4XJBOcM0G8NSBvCk+PZYlqAJNWvmMp2Jo7IAR37y4c7A1JAb9Tt/n3U4r
EVhIerB7c81g17sE+w2jxfDpzee+gan6Wov9Os1VnUw3u3iQB1ucsMUb1ERNyuaN
6e2cuBHZlvNXZ1eCsabODbmro82CoDmFz08B7ccWYzqvnQodVBjchF9rWEropxMp
bUNOsFBaa/HgSY6uh2glq1/mOp/J7tB0BBCwTiy0iYwFqfxKNVFbDT6QMiE/wFRg
ozyljxRMe6VlQJC6LlhbBp1pgbSFDlIU85o4Pm7pq8rHWhOcYYzBhIlNpLM0C3NE
WqLF2F1u0vRIMxXwKk5Hd8eUB57mZodCQHBWp6zd0zR1H+sFDS4Xe1lkwnnD4LX2
cYTb5aq7r5RMtCPfQEq1+fRnVSvcncJTILBGlwxpgAh+Dy608RgdVe2JO7sGfeID
z+QzZyMU3JINwS4QvEVOQCEcXOGB1XBLqjyKwSGJU+gaxCQfc39DBa6+toPlJr0N
i3Xuk+QZfMNnoFeFh/k/OeMknDTP4r2pYMVKie2r6y88YqXRHFTtbwN3jmV7imrr
gHwHabtfDrlMuxYmiMjjAGApaFoLogLQlh36nrTYQxGpFkvgWNRGj/C25X24fTiA
Obk64xqyqiIyJJt78R9jPzOAsRe2/Tia9yXbAAPfQAy/r8BnoMDvt2DqP5L2oxDA
AL8sf0BqxgZMg1NJ+wYbpBj6Y/CO8A0POUXaq/UsCex1/K8dXW1bZxCYnHUJwgyA
LAe5RJlIOySaIITdiAJsxj4R+K9ECTjuPohtkRjI2D4VyBsoE2tSqDXTnJwtTp3n
L6F2tfz26357rHdAkyR6jcJIiVnSF9aOiNooIvKCKTxSZUJkN+4NmzFWkfObMMnY
5Ke4T1kj6M1iJoamfBYQT1TKiVn+dMRUj3off+IqkpZe6Dls+OkY8lkOsPW9o9BR
Fm9CnCNwYUf/Ac6W67l1/+7X9OJHMfuumy8uxe7YmhWjaVahm62FCDrRHXNsKv50
u1OClV0Sv6JRgXvOxRLuCtjwYNp3Kgt4mJ2kkYI2k/fcTpjyyH1VgBBvEX/jrWj5
2KkFkYMlU952OpbwKkRCWTc419NlU4BI1RtgL8c9wk1N0gNa4lWfPxA1Gq7wPj9j
HSUAr6wmFrwV38JxhLuzMtcrfNBt7nSLAcvYj7YpZ0IAflzCBqnaKY0QThDFZLmt
mzrFp2pij/t2TJQdwDORHkst7hp2zzutFIw4sO26JazwJre4+FYd/vwIAslTcDaL
KzDCZjeoU1Nec0k5pVE8O9j2IvE49LPIMJKJjd5VmqX4D/Sf2a44YioipJGMMqff
fV2cc8ayfzyM4fk2rDuJC4GT0PBn5z10vC6lrb4E5cLOzkEi8nt8fopAu6AJojiR
0g4h/kjxHkAPxus4HpFYNBw+GiOz4ZjSBUDXY6erVl2K3jxYjtqXZD3p+0IohXEt
zs+S5V+SJqVfwxo1KxnOa7U7hCX6JZmvyFuBT3sVcV9JSgq6io8+0MSwENnaRD1g
MtSB0RKgPyT9HHZ4LLUL0mjyZrQG0ekEmvdmDJKjj8tpZgGTdnpXlhj8ZbsLBYJ0
AZGnVsnKMl4yXpJP5qBbVM5VXY/GexE92CTr+kWi+Ov4vlvMeKTQe6yh/8WzKb0p
xkIJpFi0FePUpQRyr//Ye5JZtgt/pjDfBMsr3TyyWCGOG4+dn3oX1Pk2bFcw0cxJ
rjq2LhjmCoLxSszl5x7D40z692VgDGwW5H+pc0l7pEUjfDmwohk9kv9gHFoXtCTm
xP2VzzLigQkLkf08+d0vWbsh48+LSf3DgQn/MxcMvPegdSseSIezlySgHErxlsaR
SZJPeTOUcsBJLNiiLYIkDvTVb+Der37AWbpq8Ov4ZkIrX8Jby29BheNaZ7RbUgwO
Du0LPBYpAU4DIvG8lf66rMUZgNAWiasEQcdVJOryDbvlSX1a0MqBGXcrtAUd61cK
+6ysylkT99awDdYjZNxqm8NolOu3eO1lsQKFuFb2I8xzPpPAPQwYoS0Bz9/beQnS
bjCLaWxNBAITN+iQfnsK/tMfBB0TbRjoBRnKFNKqXTjsurd+b3x83XtCrKzcK9at
3lLuPr7aXBE6wijCfrAGIRLyRo9XijEZ3ZelKJzuamRIQHk+ziEQBHJC0rfKru4Z
AZi9SOkHbGhFOCTDk9GO+eMieYocE3GDCUIKdXyKsA0bXTNOMNGplJrB5Fah3cff
jbitznDisa+G80yIm5ikGxv7dXgw5ToMSPnBgwXv/kWEG9FNji/Nugc5RS38GRrU
MWW50mVrepghD/8LANgFATa+SoHX72+HH2iqWD3K91OlWiZmY0KcYJMcrMzm+mV3
U76TGqyHP8oT1imA79fElTi4enKAmUfi2qJMFsVGm2mTmQq6YjmtRg7W0I4JQidm
3M8u5fM3sxRdxaWBqocw2EIsuAvsGe0IYqXbZ6q74QvTOmONZ3WfwykUExV5EWkC
0CEYiFzcEnocmmWCahhN9/XWs0yZ5riF1hhhYJTTRw29auaQ/ynRj5ngBA37MQfv
docsbVxolx4s+3ZX3TslMAW4uK1F62zp7ogzhcSyzf8u1B6Wj2Mci+ed3lZWeQ88
epBTxLmR7S3fXkzxX5tiGP5Ls13WbOM/2EDRYVEp0KtDdpPowo071uGF+k2HzHeO
ye9YtKduiHF7xAEPDfaS2WbJARWRi2gSOWz/ZEOsoo8M33ML+tie+fXi8SBkk+WY
zyTvvrK3UMMnW0zWNe9nxERVo93UtEJlBxvihiviPS818xi1SwPipKk6iR+oMUtp
a/0VCgrMFyH80FTimATzxfVDcSuR8W1Zfq0h3t5MHj9jeTG75jaLhjE/qcptyuKs
BGBxEZXuK0R2vTh1OmJjeXU+shpHiONxihpnzYRB+8l0O7P0jeFD8pXzzP/MJ+VW
1/HqQ5G38uwv0nB18EoY9Pia0ZShrUCv5aqB7cGf1CmE/aN4p1nejpikWFdxc61u
Q+hbg8/U8eCN6EJkCGiddSePZvz2ONesPZmAotyi2UONj0mJ8BYOVkasPWZ+U6gP
L6Knq+65AYTLQLNxuLmAjpGRKh1yv6D/iJcpwMlVSK0CfiYmJ/PUJNH4Zvd/HcSm
bWQp9TlNOVC6L/WNis5hYst+NYaXXCfw+sdyysQbvMDn7ai3AqWscD74c43Gc7Ms
WJkNtSC9/zSk1UD3qoGFwTTw1QipR6dvcPOU6JU/cGFzeO22HZyA6JeMlqBv+uRx
9BUBqUeOoKgqci4Qf/Pa1Oxcf/OyvBwuG0SOseIfvXay8HDCReCINdmB9ab63Uk4
2ewkCIAP344KZ3KHlx5SoJMpKzUULVGnIJ2WF2QupiCPP7fhgkuvIT5Fwi9ufkef
wgA3qSsVoUS0t5ppbCSHnOe5932L2tqqskorTGxNuEOBq95+lCZ3U931wv1qziph
D2KtbyaWn5wsQUcXHMHcjAaDSKQmFfhYZFUuVF0HRN0VTu3u6/s5tAy3vzxaaymK
LfURq5/qH9MGsa3iKdOfn9IGVE6AbhJK9wGkbfZyjwx5jXdlvObcULCHtc+kaqlB
Zalvz1YGMaBL7UsP8aNyAuiU2pSNH0rmbaSdqKwC8GbMuivKiatmYznqPqY5/4nt
xzIuMgSgq+Il0bEZPTGb5f74YI2pVQtuh3BSMvjqBmH1qciXyE9YVi8bri8WcSr0
yThh6aUWJDwYNAP0EZEodpSTnE3/C6ogL1ooxIjrhfA5x2aW8G3nipSe95SuedlZ
9K9YLoGckkYF7Legp5aREMYW6EA95etAVXVBY41Aa4BYYQ6XrJsZWVCmfBJNL+Z8
+q0CDKhQn2AYB+i3jcp6sriutWz51JTcwz623ROfOk53LWlE78cIZwNxO4XGABZu
6Kz5MJ5y5RKB6dypRjEumJ54qJ23Ji5ZFxRpWvP8kXtWC01VJlsUtPZ02fpQyLfW
KlQoQYnRDDzTY1ZWBdkLeqx5Ki/Y9rZfeLqWUqkmzvoGg9zpUgi9PftpMoN5+4o0
Gnaz9VTNN0yOZYQUYCzKLcAp9JAW6j92h3rIUV8bBjDHbA4sdhaavVsaRfJ5gcE8
VC0CSpUO3/hBYIZYIEaL4gCwItv7TDhyEWBUReB41eY4xcdOy0wyd+tT4fHE65ji
5ObM/6Bt4vX5DOqAd+XHDUTu6VhX2TauAazCfNLhT9+aPqcif9Y2sBOVqGA48z4Q
+SKQsED8JFhCUJzZrcuiQ9hLQokRgfloEQyI2lCESEHUqSadgn53skRXXPncvENm
8Nvxtz6NAUOfAI/8M2/xNT6+u9NcZL1rCNvCPoC3/r4o/9RMs95gQtAvFMe/DF4Y
ARzNOpw+pzAaMpscLlxzRLgMlwFeKlnXhwPUq2UkUVHDFhUS2G1aC+lg7nWf7g6w
56W+seKYWMLdvyhCLVoK+c3e8Sf5xd1LyJba5XCoCPI0UbvYlw3OmuTvrLPSBOQF
zg/nsQ2nfilflcnYn0d4LfWtuk9fBXoSue5o72VK08RkcFtwAXTwl74ux4FLGwh2
8Ln2B3PnXlCOvUgv76fZ40m+IIQoo1SP+XL/uOHZHe5i/c8hqQCxuB3+c0KbjxcP
/ut5O+VFKadYUjanZJXAnZiK6CA+dQku5VT8kGyL8diwirZGESOmQpEFF8sc6PBL
sFKm6zSolI9all/daSz/je7uw+SaqXtbYtdT+VZt01Ayij6C7guQVnK6g6cGQxYY
d0ptjgUlxRAtW6liohxGRcBme4+N8m+Infp3yy0fKoU1yKXlSxI04gbP+XFE4M+B
zbAcIURTxXzviQvfOQSrMGuvtfMXI9J2qqsQxT+XfRoEwcIpEtD3i77nUKN+x2/y
9qKcUy0Q6/OmlYbqSrG0dQ+Rl4y9xrhuYS2LecUQTl0Rw4IqFzsYF85uQ93Lw8Xa
7LXRQmloMJz94tNp/rRE6+49vfdkKXofE089WBS00EP7zD+bnwkN2F1ykk1763N7
gNrsuXKhaGeEyFn4neK2sltToTGUdXl+iRjOH4Xsp/QTL9jYkubxIRVQLjXSCwFO
Lj5BghlP9135F4Q7MP2PtDyZq8F5hefycSWWA5WSUfF8Wv6Nk2dnh22bdYFODEWK
lZGsmiczJ7g/RWmG3OJNmqcC0IWGmYk9mLJI+t8sPL7C95Z3MgnmTmPPLDX4SxNc
MwsX54UuV7OsPW5i50+jBMLs4pSnPSALOT5/IXXmq4QZE4eLn6OwuWxaHbkVGryT
FiMbWtriSUJVhxF3k65z7GNUDTRccvbTYsw8MyVNwvXvm5/nNZfues586MhZLC2V
Timg1DsJ01CWBvRH7BAJM6C2h9eFIahXMxts5Wlbbgfav67qkK7CydDJ4hdzRofv
i3gUUwYpCwT+MDsjEKY5bqytVF80Z3cOgtNAmtoUCQi5hbyhAp6nRuo3/ohOqQns
0ut/UQE9962bgZpCKkCL1fFFipb1OFo9lyKyePczpORrCrg1OPAkMyINDwwnbd9t
D088C2dBt3VwjAskqMdsFe5U7Q7zIx+AB4Ks32SFdeOUbskEDM7M6W5AcmzrA/KY
dzjO+RzTjqwewcoUTK/VkZ2fr0Zh/8EBUZW1kDW+v45dFE9vUvwYi3Dvfr/qTMiI
SjROYjGC3R7nxw/Zi0jpHuz1++Ht4r8/XfUuI2NOmFIshIwLbtOfheXjB6pdYrUe
IkgfLieM7mT70hG98MNBoB864+uLqOPZK+SdguPlYtkCm5guRSTJ0ZOOqLBfXxZA
ZTsAttx1jVYR3zmCZsdD4yHOEnkX2QdZgPHei7a//8wYE6WKbxQKlibBJ4XE4vQl
VQCfc4ccPy3LW2X6nU+QW6koKWUkx+/l40+ezYRnCPHjo9sxNCDSu4N9h7U3Eo6P
/VTiq0aq8Tpf9Rn6Kx1+5nuYZsH8uX9SWmsaZTrfZOxtUNdyTlG9h6tUN00dHdwP
h0l36mcFY+7iIjCAX8MdCpS0O9pdFPSdZAx5RNvQsKiKMUEmWPnlECIMGg2iQ8vr
nTSGdlxqwgIfYJnIWzdkTBzw7TChyoFUNFrFuSHrPSTut4+VXCRZe5nBl8mxAlaW
HT+r6T8EsNKeRZnDVd+3Rh7xwCX42P8v4MaMHTL0+s6pt+09TSTzf+SEkaAA8e8b
mQbB8BLavqeTbDxfeBjJx5kvVoCW9epuOvreGS9c20rL73WM75AcHO20nFaajfkQ
r4RfqrTb2yuyNnl69FuLs2FQjZKrwmv9lqOcHJ2AvPm5+Y91Cf6eCGtTHgGbplZT
lsgVvVY5f5bEaCxJPIUlRcs2Y4lWrjf1uA/lfXKV1cYBYEH6GrB4IQ0t82WpQu3Q
6Rop5qYMmKWXBl9B9k0lSUBpYjnXWxNNz0W7PbxMLmkFZPna56UL/HH3DY6a7/46
AXjv1ziZ7Yl8U5a37+OkaZIcmrygmPc5svqICh4tw3qTZbLD6WjUR4YFR3n6rUjn
JWk7MHjoXXfi9EFp7DlFW5OsdDu/igsGl02zscLXWTF7Mw/RLHD2J/VWDIJA35uy
vpkKCJAKv9VMLS49aHCH9iu/BTvIpuNfzjW7MJUVVX8P9N6Z+C4IrM6EkPaoiCv+
UM8o2hf5Ho72CEbB2lD9sSykmqnF1wDudvAEqoyPc2TEkrlbPGWRFsvT+j23/R8y
P1TspdIbFFu2Fd2dM/rXXA0eDml3A3aftuRNnO3r6T6oo3ZFxWodpsObYDnUl3PB
lBlpRuWeqS/j0aJpRXO0lVw2Oz+q4PQVkySazsysPnw4cpXJShdGGTrwgMNDVXFX
NjHDjAeF2dlhE5c8OnVnHFzhex0meeKl/waH15DUcu32B2pSg9lavBme+yJ9f7sW
msfXHCJlIQnIURoJJeDXX3VfuDKgy5rEP0TcMX2xg8OumEOyuethQMV2ZY0OhkQZ
fpvyEN6qUkvp6HEE9DZXffe2cnaB0Yb+9rdY7mvVSlVbtgkApug5rDHoQO+Y/S/f
LBIxpmh5iAvi6lP36qufapgBsLO19VH1G2y4GWW+FdtRg4PBmNozejlmtKr7BzQS
CoJPntkOfAPYgYtQTBQF4C/3B+m3ro0MCO2UVHb2Z4juqSkOPtiLfB4ml3/i/GuG
V3s3zCpfoaJTfyczqOopp5EEJPLPG67ycHiQTuS7ktJPyZxDF2SwQ4C1a5iiOf6R
YQU7Ki/dviZ2f+rXxRpCFWvfHrhfSCCwZjvmcq/tpGt2Pq2iYyQxEneIAZF7xqvi
OGnTDMOSv4WOMm9fsjz2XUdjb5pRgfnPG7gj/EAl8Z6qA1s1VJbHHCmNn7EwHZcz
ivUGsDE2Cs+5ZLSCTiCimyzflyac3zI5rKKQa8WKA66YLA8cpX3A0RYDmJ5YBPYk
6FfLhPZid6lYxJmbttoaVm+ZtNl2kI7mBX1eAG2RV6wS/NRHYZwWTzLgtOswLoGa
RqCCtPmqzQJEBmcAbF4Q7Rd7HE9IywSZ+XPIbfTfQJdy7SsZbZZAeLPTZQmPpCWy
01rDMqVeYSb7KAVHkcTeGQ7rhtgiN2hPUb7B9sccK92kV9fnokAnO2r7tiY6F1Vl
Dp1tRkFaqCIM5yTJ0m2vFsioAD4cEooBuIiAyuEWXhEZeKBmxWkrhAk4MkpL1Cum
9tdtiNEft2HHDGQTFGld2YDorbgZT2X/uyQAsav3rvye60FIO13tLwhHoHj3AwIa
E7WCVn98MEUY5QXqHwEWXDfOA0JiEIwXn7Q3RNzQRUJajtaCJhclRglFXh2FVHzd
I0zMUrKS1u6k4djjHp8BAQDoXFr5VA1tKjFDFzEJnKs+Q2pyVyIDsaXB7exyeHmB
8BDDfu9csWJEUSsRxXrvEq5/1KDqNOwLU/ye8MdPGU3hMpeYsJfLV5fmhZ5vT+nu
x7AUaNOHwbROSLXDq0dkwodf81pNURsd43oRUoNQaK6/tc3eu3CgEr9/BmmTz2da
CCco83oaw1kPhXhmo7ZcQzVR6lJ8hhwpwlzAO+aESC474oQPZDaJ4LKBdG2wvS4p
v8W2zb2UPe+edx9l1Ag9Q8hIFyHLClnErCIn4Hcjmxd5znTmtPCFxCc4mycxBbc5
VG6OUIrpJmiYgCofulw+2QTA3Tpn9n9CLhI9nZzCr8sqz2tJ6awEDPC86ji64Q56
YN2qvT6OtR8YVBBzcrA1vO/MSJWLvkXvb2bSIagxMne8a0QmV62YZNMfBAfJmIds
H5GM6JRAxy8qYNMuIIdM/ZzM+Y7DR9z3fIqNQeCIJ3SQHOeYMx9bYuJxMNjmgmU9
uD+h+um9aQt5hbvnxZykOt90UpkFckltko3eXgXWUCdKOFcI4JC7LEPXPYgbROlL
oJANoSTaHV8daLUQd9SCY3a6U2JT0nHXtpdywlHstnRRERctwIEHVaRSW9Di6w1V
3hmf6ITyJFHGsY2JJDyXdJsg1lUl+v3NRX6FWms+3T7zNVZjDRD0sAGK/Fj8kjXj
0FFiiFOrWxf6T0fAyISc7akXy1NiRaAfHnOwsoL/y8CYY40Er4oHh0eJFiTuQ8jY
e5RZH6id9XMilGRGROXLzy+mbFrJenaXC6TfE1fChPgPd8HidEx5q6Q+HDdV7sMU
TSdp64OWg6EJaTCtSUgearcZatmMhZeyM+OPLFl1halKWqV2UijeOua2f1lE2r9J
XUF2JGWii+vgcraZciLpoMxqtLVErS+e3Ynlsf4KE+8gaek2gK/kOsKYWc3xGzgZ
KrOdOsD95n7yEzmQHqfXFJ9TnF8SHZpFJb3YauYQxRhaRBckEo/3+gBwrYxDp/fU
fcVCy+tbDUZqEUA5/Xvpxl/zh+m4hQ2W7GgA4ZVOg22zCkCQAy3j7qrU+myiIzAu
1CXwx+cvU41ZiB/DTZgHrzrvBNbQwfFKnzSw4I3frBErabNHlxyPrhwSzaI5fRfX
3Bx/BaxiWX2eCAtasCBda8F+rxc4jfdYr9gNuQ4Oqd/Z51Tl4QX9dLB8FqaPiEq+
8H82c44kLFUvxQUUnR3Eut8Fhp2Tk51znJNqDJWN6ZUiR1K4AEjjWV4lHrYcoi60
UWJ5BKFMnM3VLNF2/zDvfNexvioBiINK/G1tcCCfpx1ji36Yc3+RhZW6bUufnW5J
eDptK0l10B+qHJZfDcZp+X+YvKPhghxlQhGGc7S7GQrcxlYgYq7tQYQDqzz9GPnx
sZinXYE2PoYlkiFkF8KtK0pB30RUSwAfEercrSvUEo0x/6Kih+lKkcZLKojmuQCw
3S0RO/VHQVQfG+8ignRcZQqzRa7H/hqjl7u5Pi6Q+IndfvIFTLakVh3NRNKZ5RVU
kNAOyi6G5abBH6rE5PtMJaL/oOx/1+5Du/vK0VBRdvPIYeTYSpK8wrU8Cd3HbkGk
nn1IiwOaMjYLJmeWgMqo6N2WGNzRuBlQaKbF88nW/svl3ofQkm9UXodEPZ7Xr3Zm
iNsO/LxZnxMz/Imdqlva2SHe7ndROlv8CpApC/qUTfa0ZhECzpLqnGDRHGS/RVC4
dj2hk7ArJeFuPKUS8txHaB/m1TT6oru18koiSkL8XbuUFmhpSDhhoyr46TfkrnZj
l3oqh00tqoA9C29ivOFfFkfTBQ8xsIFe/7NahlZ8CBscryeKIKU+y9wgNCrKzkOy
CIyNeRYUv+hKbQipeb2xtwgs9LlKqDHs+g8AlOll/Lm3UV9JSnvyIcfVaNbQMt6H
OlMXmGKV/AY+i61MmwOv+3tq2iJZACxJbeJ6jaMyy3qq6KG4IkyBabODdj5IsiKn
t3Z3lWtOL5NXPW24cTL7LuucVw7K+amLLwX9gUbp3mf//cn4Rw7/TfUb+6GcjHmg
xoL3HuN5IMuE9fwZjde+nVAFsB+bTQAmJtfg7568dOXUIySi0j2gSlNV8EAZrlxR
hnGGTBh7pEq1k0/0ZHl0Pd5FONHkgEvEOkZ2n5bGET+VHRwMpGoPVGxoixB+DQ5O
5gGwLFMfD+Q2brqAanREmg4tK5L8W1X8yti7YAnX6Nh/9eNCN14H8HuZ+Iyh5CpZ
VneOJvf5gbEzY5UtOq1bf/AqqvhhzZtIbss9jkY5NuJn1+SqWonq00kGyMhcXBck
dLIB/MObO8wo5doP8fwfXiH2JNTVeUyI+aJrX294PyWhML/V8DHcmSTfeHSlQo6N
iYgNOCbbqerTLrK7ikJDeY5IfFfs/unr2Zz34LLLrUfdWtKsFmTXqlImxMQXIBiN
o7Dn/S7UmBp5PFicgwwVpj2L0zk7v23+2ovOeTFxMugtyBWAUAQPMbxYCmR8NNDU
SMcflPNGP2i7jOG8VZu0OKLOhaQYyZ0hqw4s1Y5CosgFMzwS85jTP/gznabpzbEu
EJIWj6WOLH+4Wj00vI+EJ6/FNSmRe2ilTUIBBjVYcJMcrwxDeYCeaRfq/Ffp7su4
q6fqneyXlwVAPwG4EQvb34ZcTW9m3wy1y4l1xdcQJ2GB1Kc3pthb9w4EJ6jGGggm
71m6CNsF/Ela8jlCYI4j66lX+q6ToEOUUhMqHGcBWflXNh4+zNl0IczCWsCuX2xK
jhufaq3W7mqFKtrJKUbBAoDqAeX8POOgs7+cFRP7qzJY0iSkc8hTodgeR9BxyIJA
RXf9WhLFT62V0487+pzs5or4gzH1Av/ySkJ+L01W6Cu3O3EDpceub0UuDUrzASG0
i6M2tJflSnpVgYSXcqaGkbTJ3hWBVb9lZSmXRxkmK7WfFU4mjTNQx+3sQkVosVid
CW1PLa+FQbg027iXqxcCYlJIlVOWnd4SHhsreV5MZjw8ggjlEpD2lqWL/sg+Ae9y
NGttL/d3RcTBwUHmq2anvXXICwMaqjAor5DJcyBllORJ7Towg1IyU3C3dunn5/0T
jSf+lZQjxV1CGjDkJ01frEor7lBDJi0D4zF5N51S5OZgLtFmoaMW94jPyppJ8qbt
oGpHt/YlSB8kJm8lTbsfCFd0L4iSm19oqFta1/e4A9YL9RjyUtizJze5+vFJfnWr
Af48xHo+eJgpTas+BahMHqfuFPqNNNL8JBmmnlhniZYLg5FjvETu1btvB31RYwES
W+9kOK9ZQEOgr1B3jsduG2PdyQssHYIiDgoRf83ONq1c42VXK6bJUtKy409URcS/
GPqzXqA/BU+z2M/3zH6kb0sS8V39s9lVCkZHNuPKK/acvzOVYBY4VTG0QN3FPKLO
Usq/XYZroSRX1QjTQy/K4fv0fcvtuiW/KLHbTOdR6/kxfE7VvibgML0BeZkv3A08
2DueH5gE4yvnAaa6TncoQxXEZNltlqqTt+vninibWVFfx6+2iazEU3ZBedFdAPCt
aTSjakayPJslpJCx1KNEH4mTlzk6hzDWXSpmK1G1w//bNtRBlq7/Ks41T33gG5ZF
T/1TyBo7UohStF7nlOp/FNaIKD3NBDTs4HAqjaSeRfhsSMMHwPt8Z8iSNWj/34M5
ynCzzP8/vAiE7RmhNzPr372Ah+2EtGkWROp6xaBnflpuKfFmGwhD6tryDW/T7y/N
c1c5tNpXLXnJIo+a0D/qRismyIK3bJmkZg0TB71/u4uwDf7RRuN28oPtN5fDHWQW
DkaZsbBHDnEYus/4r+hpHdpp5qs8o2F+6KB5le2A5kJKAXvMQ0gjgdkAZiTazdH0
wWy6z4BLbt4ULEraIyVJQnixmBu3RgKSzF/sAgQfHiQy8vrUywq9OSrRSmDjbKjK
VCDD8gDONawWT2cqKNY50Cv/1ypZrGEdCVK5FEemXX7v04SwpGHNeBPkazwk95Le
qei8S4BeFNqkm24CqxNbzXOYb2wYksQwmVNenOObvzjD9dWQUHK+92urhQ+VdKLX
3eV5TxGKGp+lA6YjdynbF1lzKUe0q1K2vi0LW6wijS/Fvs4hRv7NuEesmzdK/Mb/
0O9F1TZ3nIvZTc4w3/sgE3sR3Fd8oDMiQd2Hh/w4Yrdela41HRvnM9aBBAR/zKLY
Ia4DMXNaXcZqPFEgoklfM8y5ZCRHlRJaAdcKHhktumJc9ZgyL1rRz4PPbs13p5H8
PBWe6buZ4iGREsRQz7iSGtT3F335uAtkP+28W45z4ikmz+1cx6bOLYMt0f8qiUY3
vD7EajeZWmYs1uRBvM4QoNyQYdWPEaSJO9rVhgLrliSqXPCNNcS+pdByD+fBobo5
YjX8FWAKTD0NmgGZP5GPPQHAV4+LcCXA9r7xxS/tDUem5gAkij7/8Bj+3xJTkEN5
8AbhzfnRrHm+dhmDb8NQFj/f4yQazTmGGBzEvDWETGcBCpO3v13XUxNQNjzgfat8
5jGVXU8ztI5dcEESIPZa96lLqATiC+b/woCK5K5Stn/VuhbJyyiVwQkPibYT19G1
VJ2JM6ybnm58MgrKj6PryMA2sITgxe2iEIx1uFU2eKcI6TTooEEo1ixWzgdZ6WFi
T3P2jqdtDZxiAjkxSHToPdAfgkp8Gtz7hz1ZIaqcAYhhxGupaECjBlMYNmizOig6
wak84lJcZSy9HNoEJjphfFv7lsF/PT7zASul1Gv4Os2o/4FGdxLeGQjX/+QKBIaj
BkWm5JLZgRMrnPOD1LScakfMHEHA+ZT+feKzOllxPUC4bhOIOkUBPGwLGKpZhx7n
BekW38OehwSGBYYtj5QXXPxqH8Wc/+CxyTaHDCpFVKlK/3ZPUAzG1VVQ/fd01e6C
/Tga6BuGxDAwVwbNPmiiD8CaWVmZqKoTqbrN0uoIeC2N8ZKn/shR7bRdEFAy7chH
A1IVvPNMjEBNBEzozk3g7x3B0QrLpGSYjxob9uSWLzFT4/LiEZF3I08KoLXXhokz
fXMYOK7nMt/MHR/8PmGkgude7PnTNFfs7tVRJ854kNamBaXScRE68io0zzynE/EQ
G2hn7+d09XaGk9C2o/Zkd5a8InybCKIg+3B9pb2e4FAyWkSqEhje26Myn6Ggpepl
uqSvtFsQsnlWusPq/L+bHHuOtRvtLR16JV9paSxXYhLw8fCcxxzkQiVG1HgUN2Hc
CJ8qk2ZeYJfDBGvYTvtM00wHdIonPw74odBdx4Yb1H1Fg5vthogE7o5MHMypNIJe
xbkFIMWq4YOSua0ATbBfVPk3gILsaJlkq2wS/sMzGMiKrSk4Ot2r0JgVvvDI3UL1
PuhTd6506aJbUvRNJWAIQtqtUJ4EDGxuT7oBy1IpK2Ww+gsnLe0TrSTm2Izg8r9e
ijoKVEE9eJpDoyjZ/Ey6yEQd3HzxPkf+yIaVdgK2A1lBVMMy8rGjCkWft1SLxnc/
eW79gCx5FHZ7Yws40IbdtmgjDoPAid+Ii7I4vB1mjlTph/RmZ9g/OivvHII1b7HL
4EIJFHvRI0KA/obCcitrwBL+xnuvY8wSGWP3qUQM0ATOewenaFsRlrjEBBX6hbph
yzVXU0zPnFJqA2jujFpzAhcPEcinW931nlS0597Q3XgwNaQ+4gLhZRGdjknTF50Q
3EuCu7F1ADOeq9c0P9u98KmkkhP18U6H+6QsQDBUc/ZX8E/jmaWlYazQpqZxFaFp
OrLM08IMTzZmIRgIkIXJQGIPx87dWExPQF35ltkX4ncIbpf/RO4wQuoLTuipxCv7
JzdldXX95PaLiXeIVccffUuU3gqa4FT5N38EpYY+sHOouAb57DY4vcWa1dFCblyf
d9Ss44nZ8esQIhlF1rKLL0R738zfLNlVRGYpQ/hKp2rles/PO/XlHCRaXUGEesRM
cSRsAvUP+4CTYIlQVPCks80UF//iYZJwXOPGNzn8DbjEBvxzibEBAJAXw/BN/E6L
iMDRBcpzli/rt3zHWx5Z6iwSThK2qvexbf+QR5BJ3bTLvaSD2Ov0GlpDHc/IyU3J
LweFzWjukNHYlqd/DryWtqt8tsYsBM7QSSWpRAQP8phidLUUiuylS//sxzW+qeHJ
WTjl4lkyLBkcBd6lR7KU27BgOTDVuCiyl1UtuvvpR+vrinbuC6L0O6mCDnOTqurh
TfJWlxnCjTpPy+OuOxz8AqDfmT1z209x9WFDVn6ChrKLbC0vySTeLL1XwlPx2LMV
Eeb8xN2lBH1wo3X9hHASc8TZutl+jbWnRm0pfNltgjBEHDAdCuf1J8QO8r+QE9Pl
QTx19Wxpf0PqltZGg2XadEDNpkbOl2qXoegLOzfjll1NV4FU4uSb2d43q6cB1x3k
6/WMuIuOvq7YDkDN5DHiLcfJGhU5fykH82e79a+M/dPUIKzvchrcd5ISvB+FtqXS
czLarbyVEyDeWXn2KFH52rm6N3Vk1zuhqEs96dm4hFU8pLk5QwodHJjpMaTOOUH+
Ww7HyaBA9cfx9PNEJFlQRRTenkS2M4JModNeRC25WzjnJ5GcE25GdETxSRDXrQxz
ro9WtnjKQj1crkQqhsX5j0VnLdYjUSeXL+g2ernnNs2vebqKJET7+gEQHGbxnrVU
lgeELdz05OLAxh5Y+FD68QGPQcBZuvxKsIydwVNXYKHDG3S76HIYx1G2duKVL5s5
VcG/ONKMVJ+QMrnmXZtVMEfcL8TOuXGugMHBeXf6etrWHPrp5Q8Cg1VTxuexfJ44
a/miwxFHstBAdGHCWmqNTwLWbHXIzlv4AYAmGxq/V0Ghp3Xofz0nURwygMqk0u3C
em5C0rDTnYAQ0eyS9YIGVhYB8RfD2teb5HkcH88PqTf3GxCL6egfw5NMETS59FFG
7A3dE9V/FISGdkZG0AkS4wXJY+qbKOFzib1IGf4GdqovzIx2Tr3ILaHliDRUZHrQ
K3DX+iJ7l9Qputy7Az5EqKZ4tZitNsr5nYXcO2QPzamMD7Ly+6p61mZQEnya+r02
EWIU5eM7gwbWvqJ0hg2/o88TwNE5mLn0/qjcXoMtjBenQ9mUz4HKLPqPzcKpE1Dg
KPUkvp40aJM+Wl2iKS4t4CB+I9uS7t2wwjAb8YVAZu96DxTvN5mF3t5e90WfN1l+
ebKNM6sRP1WL2hVZyyLJZ1J56cO/2QHgpMJP9AedP3eOlCkVfz4zGpNKdhI7U2Fw
1AdTdsBqyhm+PNPFluPrxfKET3eBjr2NgB9OHrKaHvIc7YvxUQJx2kG5bMG3+0SI
KZNePacjF8Ya8OIPpDid0ju18J9dl9CWCp70SkNwu8HvFx+qL/h5qRLc/p8yzo2n
GYjHz1WzVEBAKN2svizd7KINwGofh5Pmu8qcTLdt4mKkerjeivmHTpv8y6YurxAa
Mg4eohUba1eMX1PXTA+O8/AseNqHvZdZ2KrDfs1UXnhpBnIArvzqrHVkPNVvSxhF
OvA8SBv2F2TAAXEInVUsw44wYwAF03DN0ztUYqP5/u/ga/X9yiP7xShH4xDFfmFf
NSL7YPFXKn+UWChtfC5mO7JdUApgmfx+dzWiF/ef1NIwPylPfWPIeLItqo9zv5G7
fwU0h/oeeLLdeLTah8PY0jUrfJ/A7S8tQ6T/pjwV/WucpLdUDDmDg1LqDbqJwehm
ievzGO8+fqzU8uGNBke/f5HzQEWRULpd2ErPQ9JOZN8NL/9v+AADtrXpVWHNKLwy
cHek86cFbaerEmWIKHKUnQV6K/7jP9DBGsSwuLPIxR/a/FW0/I2cK6FeLfZLheQ+
eOrSFdcGREn1iJNDpidrb3oOa+T8p6FxRxqzxz24c3bDDzJNf7NlWmB1Tnljhuan
qbZ6JYgRH7cK4O9kaab3oGE/wOA73CWd30IR9mH+/LcNLvGaSCeb3MkrNkkU6We0
uDOnA2zsfgLI7yakVWDzTPCkunpFwgEZ5oonHcG856WdGec5cAKZ5oNZ73e1skGR
ftwLRPeZ8VuslVKA1jWXMGjIyJBMcck/w///zobbRmlzxuHO7jYOZR/Mn8vu/edM
tDghBs0SL4sl+TFqLNfNk3R6pBIbPfS0YNy4pRBL/MBXjIaDfZUnHjlDLskUn8cr
b86NzQOqq4YX9MnpvKpNNPg+frKzNQIlGZqoUzDyjjsG0ti4TcfRm8Urq/etKg0B
B14GY+YA5gXnzq84bD3WW43ZvndN0iHbWAHCxoP2BZAWJ233uwxAppkANg2JlPuf
HOhg+dxU6YHdfhO0hcFdlCXgV2YqQullCdJUG/Ozcj1yGDJUWYAfSQgOqfhIygl6
/5iDXyiNTWINUnMY+bSnu8sH08o5moaqfDc8PYcZOsaa1ID3yB/9uNzUZLHDbRbj
/VYVQbshP5+/tIhaWDW/5ULvSw3ORWq7Yc89y9S8hB92YGEIrPyBenUlk7OAvo4y
0RWYpm/8WmGtKFU0tg0RkQ7eRVPTIbUuU/hrErV+XXm5LfI6KHaWjGbKVSKwuDt3
JgAbhQvGrvENpV65WWHVLBzFqk0vxXloukIW0TwcD+Kwl/pG79y5wV2z+0MjM6g1
yKP6GsixWh/ml0IL6tNrWG54aGqaAn500eyPxvcQIrH/srRS5Ee39j8fYC9g5f96
1XZz50Q6pcxIETcni1SShWPpYdFOvLzFnrkWljOkFimUI2D+R3fyYwZbSrmRvGGt
EmsdjAulJoGHHNLhZYG18y0+vxrbUmi5kJsKHxjkhpjHAT68FKLBP8TVDP2eUDja
C2QvsolAGFPp0dnMJu9FNR7k7eSPup0M5FvWvV25jKuicf9ELDLGKmFiI3Cp6obd
P4JSaYYFkQaKNe9v2W7j5y3Sslmzsj/CP1O2KHvIf43KixWXYBbV50KBnHHLtlJ1
m1xYK4hOXCwQKHUI1v83REErx7mnduIc0rT3k6lODblXex3lv3UGarS4V1mglgjX
h0kHduD0w9DzYFBToTl8WRRLJJZJPHx/tvD9LkFpK4JWVVEEsruvhsyUkPTR9DCC
37SylsmAX9JqqkX/nn0CABM7sGW4IUmIPCK2FxOSxqZkTaKkVa7R0J4peXNjdz/j
elUFADTpVl6Lln4jU0iqGG1QloqF5doV22Oe+Igxsy6r4R+w2OJxm1j9lX5oosjG
vJqrf+Kgq1BxmiWCqOk23Nn8rIQLoL28fxA4DEDtuMJdSbiPy7ziTshtiJhyy0An
ZrRvJJzojhs//WFNq/XG48khhXZOAMCmZrfCqI+0/YVTgnXPHcFBVpJpVvSeoouu
Xm/BWiPDOBJBXNucGPPTrX7fnxWF25vPOaFCjFrwqGWnkhL3RDq++oySc6s123ge
dT3mZIh7b/+9uhcSx7Y/Ei282DNTQoi+hvq6Y3+TLAdxktj3CY6WU8GCfEpAFB6k
qdq8gHJ92tJrXsM9NP5L2f4DTygE+hYxR0ZJUb06dvwTfpxp1f+aqvEuoGYq7MxT
RuIsraQQoV+as6/ZzJDAbsegSE8xyhZctJgmGZ4Bb7jCB0VhyhBVBJWe5rMaF471
eB77rHnwRLRp7QVhpuS03YYq/sYwqrWi29uyII+C/c6sDroZukHDEw+ezmUctfIw
c6iXBikMypIypKQu91DY5VJp4xvsBDkVoHc61fwfH2jUAVy3kCmGTwVbqSRzn8Mf
i62mgftFPEfsRn9Z6Dko4UWf/IvKjfbRSOvQTXnXMke1UKxNZoaDH58VGefe5lGz
2hXuAuldBWdjl8aqJTK5DfqrvXwF5hl+t1QvZNYFdT14bMMHnyzSkct43j+/BLX6
1vevDQ/VcpDzNnDK758XufaV32j+3/a40ZfLnHpclDiw7SK7rjiJSktclwd9kyIc
KWjLydnMNml6EfyRgqygkuF7QqYrWYuHyMhTd1X5Bw+cq30ZfPaQlXx2eH7P9WOa
agygjfRYR+yBX39IKlDWhN5MeNriWmOvjMExwaVGltVnss4rtW5Yj6ZvB20qmP2n
TENPJ+jty1daArhF0pFpgEq32vjP0kPdpJVetH2RZGqtd2REXftlg5XGaFScNGS6
0evsNs32opsv5uNA+zOWTWljIzL9stbpuI1Q0saw26FqG2lj+rgwnUr07zG1exW6
/uiXj19pKxL6bI/EXUp3j+hvA39gHI+g0FqbUpIZ4GoqNOvv7/uIyib/hXfOZRij
Wyphx9g+Qt93cIcXJSv9TaVwxT74zisnObmphmBrleo1KHSJ+9cFdaFQfpgADSFS
ezrRzmGKSf+Q0qUqI8saE09dWgsBl1plrV42MXY11QrqUENZYnzpq59f2G4OT6FO
upudBa6Z1vtuIGmqBnyDhtXcLTT039TLs6NWSYGDDDvo4em8nTck3bLTWfu1yxNC
ThWmGdEXsYJhxK0Ayrs5Pvc0ulJo1gII3/bprql7JnhXDVdAggggWf87WWKm+CWl
jtXw18U8WcyEfID+TP2clB00nF6S5ZK/aTE/h4EWx4kZugVOBzwZ5weBnVGcZJ+O
FqOpPgbL3S8EJs1yYbn3CQYYt+ZJHunlfqiWfdEBOSJHdGVE/qec1GUeR6A2b590
awoWqS1Q+7dKGSrZeCt4EQz9XYK+mnOkdvsP8sHqgdFOKScfwc0+iLwupQe0Dk6u
OBB5S3apaNaHRgQv/X6JwYpCKH1SXmDEEP+DNI3sz/B6UZs3e9QgC1eZl0SatEcn
bnx1rqGqkmFXEPpSwjvUQRU4XHailwOXsIfSqVkRF7CSWd4uzDpUVKVrQWcee6E/
RooDwEzhcPqAX1pJqMQIYeaIoREAVqZFvMYsSRqjmygjQkWdxK7rzNGTt+57Uf8k
EwZ72x7Q9H1o6bFUKWCBKZqHwK3MmV1lWyC3tkoUM5vwRaolnQtiPhGPtWLEvD7w
PRqySnrUGQ4hiauZkh10iBw2NBfZRoIWvwNJMpIsdQjoivL9i/d80PadmwGCwdKs
hvnUyMaOn97UHKGrBo97VhyoyYOei+VHnMOAduavdWRxI8iHIc9HTiJK3xFSKSqS
17e2rKxCvp0SoYi1p+fq5IYYiye2xcqZRroflmYQRJXJuFiBPlnEIvoCNT59p4VJ
qcLtaHu9aBdmXNgXQkGp7yj68T+Oina8pixew47O5oSgJvspDpUqzVvEXrkOcK3l
2AQTT+aOUM/g7jabDUYxsSt/mXFnEbNKqOCBs8uZyqJP7mg4W2VA3q5mW2c2G6Zc
DDlu3JP8bzkJtQdwQf5o68qMMjwrSInf3PXlIjDV8zYn1pis+aBV8oaqxsOZeM55
09az05DgzCrZJibRvtcOmxRnCsAMfSoPocWofmvj54KEm+Etp26py3DMXGcMSHst
x6BSCQky5JyBJuCNxcNm3pKuCoWvJUONFrHM3oGt0vp4uu49VSnhcsNQwnvYALuq
q17oc/X0NYRjv+1vjEJFjRiteK8ts3lEv3zPOtGKne87g+AdbnJBk77/LH5aGMIR
FBW7AE6MkBQ7T4En6m0kaCc6+AOQXaPin+Rv5Kzp1ZP1yp7hiSof1BhJes4xHg56
1PGviVTjPMJn7hkUX3HqaHWTCsKF9wGVr4TFF4lagnzVe/c696jwR1ZyfDcHKdmR
lEecnQVR+3JuKAq3QCgTLvvgC746+HJu7YvXc3iTqPPnk/yvTwP0SjuiPjJ3njIi
olnova7H5rZRcd56QRykmNgsxrrdXJUVf96jCdB6yuS7Wa9KgcdJRyiADD+zDmld
cpMl2YPcL+ML7Cii0zGwNDP1PYARcxCbfqd/xbsvYVa8/szcnd9hAteiC9GoyYhe
TpW7LNo5MH3mChigApXNTAC0ec5X/CXG3+FUMFcEkOkqCB5rxAaK0QU216IdKLby
CChxsbhvdH++Vu7xO6tKZktWsN+1pxKB5gzeh5u0SElHODD1kXsnNOlseoMYkfzp
nvVpZnX4wYIV5X1C9DTUGh1PANPlaUuC886p9Yb4x2iF5R63iAIeQI14M5HIK7i2
t8KTN3vepxfxVOIURzKeaH5G5lmrjOMaDLqU170OlDPH3Q5lPjZLFx+0lcZCUThF
LjSwywQYYKja9o4n+BJBu0NNKoG1QpZdUM1il0JCgjImVwdWxnelHhN7hMLuBpgH
yjUi7cT97hoctP878ZEGc5GVeO5DZ5wlsZ/TyoqNMetP06Ph0gEKOx//WUhJ1gJa
vLHapa8e3NVUG8CzoovuQp8Z/hxcXT7bjNVlZu6L2j0A/taSud2Zgc+t7Uyt8J1a
Td/cwHRjdUQGwjcBcUyOBCb28vmFdsu+uoyTPeDaaOtdze8SW0XKydP3MfXnJuEE
JT78CcZlsstwhw5tKU5MaEFjT//SH78a+pTfpf0WB5+rzkoHqoM/zwSINjZC7ktF
Dr0sFup3vFJHqHFKbEeJ0iDh8MpquhLqHqQDQGABLq/Rs/wQJYckf7lb/A0o1MYF
zwcfhtuiV2e0DMuKIgZdavm8EdoNIleuWvKGQcOqWEW4bMiya5zUyH8skTgzYd+2
UhAver54OPO8s3iWYfKQlqc41L+JePWC7wmiqVoZNMZdqss9OAmw13rGeFk/DEM+
Ap0AApYtUDlaZOQktJXyBcuiBE8yUmntoGy73nqr0Mc8hsJRTf/gKBVJVGrdJeX5
dpTN34qooUoNHiL6r/Mtwm9xK+ONJlm5DtOdhhr+P+8FMFrTdEL6wtXSYmTufPjt
UI7aKmq9h2yOUNH8NnySiWkV8PQAnC8PLq1ieUkOXjTJPbtIChSGtamsiT1pGD5E
carlaXcO1mYjejT6QjNVMYcd6nZ7x4YF41cSHzC8e/OAA93MICq5hJ/boc3Gmmog
OPmnJgxn6skIfkxVZ/mu+q657FT1bdwNokiE43cAgzrqXOFBljkEieVd3yz/HBO5
49FzlmjaLloOJIHFmnD6jFJyCrBoeZIPFviTcoa4XJkPuBhLU45c2TaKeWQRqJsG
LfeEhMWwDQ6Oo7h4ZT0tJfAH+Izgcc46wEqXK7NNZ0MAe/DIorBMXXZE8eUmO0iU
j0hoTRMUo0lWFwbr8XJO+AGBF18DjC9kODUMYoS6l67Ukqx1neHmY6D79XfijPtT
sLk1SuJwW03qpDK83ltRv1blObna8ou5DS3hy1M9ZNJDMXeXaTofT8FB0Q0r8i8n
CpZ8wmhkCz5vk/Y6WI9FjNYT4ALV1B2Ndgy1vjfN9qncnXMkhhluFHygjv8eqPWH
jRvKrPzyzN9Pe2w4DtUbhLjIav9+vfwOtWzllih/S9dAh2NphDaoiB1Y8GdcMOA5
14F4MyrcaW9cBsFiVbeaZN+vSZnWh4hkYhe7J8g6R2Fc7DVhn3upTQ2YpWA/OXBp
WZ7PTtO9Zk1+/EoWgE3OdlsNtThqSq3bQW1r9fi+l9cuk0BA2pXoClQRZcTWwyad
P/DS18Wv4O0laUYqf3WQUFSXpHjJOF4Va3ERyFYFs3FeCzd7yUDw19ADE1G+uoXy
oE2Zk7fhny3zGpL/fHG8oPdjHAx0NyFU88QzSt1BEwSWDJRPz59sdddctK0OnvZU
fbIOpoYp2GQAfw58HTGq1Kc5mPy5ohPKTyxhAywrwwlTZ/BQKxUB/msYO3DWyJxO
vHCVYDkjys6ZLrPIqoFS3GkXw7nfSAY68ZpokXZOo8enc+HfWNlM5QNt2zsV79a7
YeurFlilFN+sD9Ir7+SPBaR1WljdZ0UUjAh/XLA775KTOkzY2+J9ZJWyxVo/N0cd
FpNKk4p5X/hbDZ36ykWpHQy0UHOkcS0rjqXC9c7Uo+fQjFyp2veMMabVO9GO6pYb
03CwYVKD1d6gELARfw3u2P1O3BZlB4+n+v7SIN8Q+/AwVsL0vBHtPbobCZ2tf8EO
a4or5gA2P3fHAsWD1c9kigVbWC73g8l8Tb0NV1xG1wnGVLtHJbNBz9xNicruTYG2
CprkEkghpPnpjDBM9ltDcCc139OczPeiXaLjsMidLHFXz1IvXyXliOWNME7bzaul
8h000Ze7y92nxeYoo8pA6EXgAPIItS3vjU64uymmrI9CgHHKyAhvrf9VcbLR7OMs
ibodK7hYB22EnBDrc2S3NH2DNajpXAu/CLpBtmVo1j9vigJQiXrwc5VuEBuinmkW
fbDNq7577aYKTIxh9Rh1bdzmhOEoK+KzyMWAW546w5ICmeQbwphvW8JUj771mvdx
jY0m8eCrGp0ftu9W6JdLZzOMvTNDgiTtDRF1nnABypkmT7uMAV8PSCdJjkxEx6F9
pSyKhA0QSzna61bMaS8rlWgkZx7iy9c5XX+zu5e+L2YeJIcPHudqYWuWie1rR0nS
aN571S6umHJe7DSALkQncN1oNeulXb+FWF4N8G+XW4v9eMYF35JRHcB/om3t6eOq
1WBBM2hXeHp01CAP0cRovUZfIhvqNxm3K6Cr3dDIC9PUD/oXS1c+AT4jIjlDrvwm
mYIJjb5b2FqiKxdLKqzYkql3G0zRyW1mZ4fWt75yz0D2QQh51A5hr/nkCZInm4J+
nbSJK6JF7US6aHjVTmR1ECG6ZdgnmiNDWutkJtvnNGISETAnu4I9L7KNHDKdXwLy
rOPnDVDu3ms509dvGZxdo6R5/0AcQj5L6aRp+gLzzfHTBiwSyU8RE9m7BnZLDU7X
UZSwiZDE8ax1E9yZ8T2audCyCJA1Q2XxzJ7JZb1eoHpMkcLxIRtcQkMj8QzBvf+P
cRuw75Cg3MMtoi6DDlTYC2x9r/56Mxelh3NHZTOWlljALyD61YYpTjGc8bNXiAL3
5jldHFKTCRcF/OWfzHGOkhDI8IS4Yc6beF6kJkv9ivCnAe7E0Xw6FKiXPAsBNc/G
8v+nKpDSRKt1RGgXpat6NBAEct9pe4U3g7gYRdtx66lJVH065yKg6lPgh/EsGdr0
CqMUF4Q4JYWt4CWYMTGUh7LVGzjZ+0FETvJTCE4y+hzbwdi22MYfQnd+ltssSAqi
xaBa1edZ02GLh1lkUn4w1XYRYEz0TaeYX0inxUj1n6bAfgM+9wj6L7rLbH+mINCE
FkkV7su0piOItYpFmIanPeZRNy1d1V7dRF/eDt8m4eDJKndDBciyCIWByh9OuKZb
62eGGiyC/nW7ulj0z789cG1mXLuVjUADkiNW/jPQs9tQiVNuiM8VMywxCd3tb52g
dQvepi9FyG2xOIa9bodsgmbdU2Lu+yTTrxLr4MKnwH4u2TS/xGusk2eHj75vdbZy
QCTxYwGb4/zUIZ6MJjNtTvM197W/c6OibLpnlwvO49Qy7IK+hnUHEujQaFw7+o0s
lE9nQVIFCA2jEcE6Wjko0ltjOuH4ofLLpDG8+2hHulq+PENhkqCX4koOkXetc6iP
TgtF/ggLIk/mFz4gFOmFqVmZxcFktWLuVke046sG2Q6ruw8mnANgqRNVsqJVesmf
8wapwtpE/rofwjl0r5wqtwqrgPUnO4yu8pLN0ie2bFEB+V+j9rSi12xLBJZJRprP
DIYZYfnXPtzhWGwOLjqxAg6mlwDVJRo0qFrgpK8LggIqo5ErbFUE0tQTJnQFZcUk
SNOpf4FXYCaJJtWwqLmHVDKSXIuCL/fiVQeFsQjOIgBgysM5EiK+kvyghAXuOX5e
baEkZlyJ5kNmwqdtPfXDf8qNNX0RoPZkty71s0g96sFLTtxWSnM1ua0Tl/KKSF0g
ApqI5eDAKMqJSbWZulcXEW/BzytPEo6KRy1A342WxwIGKcmx9hg0evaS30bH6HJ+
uZ+Qj0jFzoPptAgLmYiqxkFzS1LW1q+eGQ7w66EocYpSxOv87pAbMvD32Dd9XIFY
P5mnrSf0/Aylu/o8UqsxUG1hL42ux/AMgb1N/6tll3VCrgGfmqqP6kO3T6BPRLns
GM8DNsLVT0zPuhN/GgSUR1WiBy49kYTfrl1GNxSXcyRl2VTMFiCzlipDE1Lpk7qJ
33FpiNNKlKyJWVnv+8xtyoPbwo0goEfqveMcF/gKyy42dZhJFmok0Z8QiqwK0Yo5
sdRKEXN4EWYwlT1qQqUuB6BocMO+fI9NeKQU7bKTqOqKWtx9RvRjVszf8NHtStaY
iy+ZpFJrw3EioIak/igMN9xrp05sJnLo/G/hBQxDor2pXZLmo5YamJoFGBj3+CTZ
IJp/p0QX8SxrZy99YhHgdkZrjcPVCoHRKWoNbz3drJioe8RvShYoZu1PYErFqF1/
0B721R925aF4ICUlG88GubuZRjQHcxM6V+bnjsKVVnncSvS93WI7GaWJvGhZOV9x
TTkQAz9G1Ro6WhJHstEX+fEZ0tTY+2MWHT8OcJO2N4O1NR/Srjjhge0fVTnCmfB0
LgjipOzZR9P6clFW0ebpsOnY1+2Shm46276bL1E2sY3xal39QAZRAUY7Uupo7YEn
oWrbIId2VTGFygJP41k3uLQPibDPEyKTHyrbNkmMfcBh57liMnfcQ6eF7hiRuu4N
TPlZi3vVk32KDRq+OCt3gw0Fj3t0TDoT1iQeUspiHYKyEdKc3U8O9Ugk0JAawK2E
h24xaDJKECZ14TiV2YLnynpVjedEs8yPxyCgXPE8VJ86PQrdxCUL8QOray5ue22G
sm4aIHynFInfnruU2P5+M13dJTDvoQbP6CQ51AK6G9u8KXpyjZctiZCM9/My6JBn
dcFVVoio5tQ3cOLF9Z9qqMxgzgEnmAyipYhPfjwj+Dr5lvPC3c/0l89UFmsqahz2
xj9g3zbhe+aNPaTalaW5rypt/3JWCgApyomOOLaONyZ9rlX0mFp2QqIyQ0hKfI4b
sgZKkV1cH4JCDMWA+lddqdMbtAnRoxe/ir6iZ+zzxu/fUB4Db4zanxQcT/HvGKLn
DorgjmEcoHKE7xI/Bnly47zw2v6Z1X8ZRqEHVaQW1QdDaoMijAbpCvVILZOFLsKE
ECQijhBTtDl0ojVLjWyZlwn13xszPNnxnGIjBpUb3HKi13vRbU4+jOUUeSE3axqu
60J8GRb4UuIW7JLZjBZ/LdfFjxNFXgd3JllT+fN9XVy7AWVhZS8aptXNuyzgBLNR
4fnpYUT3CtBN1RVXdvqOGemx+9WQx4Jzpw6lJnSmA71mo/OcXcBShW/k/mQrG8JX
pf+eamjQfxkc+zuhVrsiAK/w4O30xJ+4bdoLT+YUZf3MFePEWPU1jnqroDIIorJO
C+6Q67hj2jExGzdrarfYSaSGiHFOYBrd2O0paGenR48zDIbrQZOfn5HjBM+h8jEL
5Lo+l9EIvKG6fRFRjdq8NWiZrftyZwtimG9bqb/iAlIb1eA8a0dz1ye6MINhJKgy
sOM8uhQTliMpXkU0kJ3VbtM/HfL97gXbGeVeynC8M63c0hD7hGBbo5M9wuveSaU9
P9pWPRlHKZcGfKgEVrkqLRRyWPYsdHAMdTxy+DK2DdXwtAFNKs9uS7nHmqioVqk6
rQKgx/uLdG5tFakVOJjGLaQkq+hTxLxUCdAFB9D5XtK+Dnfb0B/CEu9L8ToqmY0C
LetunQO8u45v1MLoOiXGf23Xeg0zWw0JLjh++Nn4N78Am2LldxRuwH9I2NUTaqY4
4Ssmyq/2n39EMpiD8mucu702taxyeWkeiL3xBGSKDjq/C41Fx2SE6Lw0XB0Pd+vL
Lt0lLKkuA/dFTRvnXda77iVz/U0vHrzOp8H8lXuiooc7mFLroHg6dU96aMd3IVLb
XDN+BFTNi9dG8wslJRNPFJbwd1DWj9INFthf+NNafE3DoP1qgLu0veLaMV+cNXH2
mOib3Fp/NuTOvbiv/xfbJrbzQXpzJuHBtu5h4x1xW0PeJz2GE3IFd/UoTXIQVf15
ttdE1vdFTXEsif+OYqJ/fWhH2ycY8866FlrsNk1Dt0HuplETRbTN8hTP90b8Hoy6
7Uz2cRpsKC7IGTp9wQIS2umwKdJApr89pCp6+wOlanyzgciwAA9x6nEQ990yvapU
Dm5HUAZk2DDItApEddddwAfjbQJRVsjTPozOFi3ZF6l6RNKBMg035tlgoVYfnLMS
eJL7T/Vz6r6zbhcnaXhk+tXaNVl0MMEPz5iUkoyy9OrfzVrttH4nslLoTqzdWeEW
YdpuKUundr8d6By2Q6YM3/Anzd64WWTQZNkv0QxE7jJ+iss+UWFDUH1oh56wxgTf
vg8O/+Sq3BhUISqtVopf75KsDZ3ZbyxJUG9FYInOCKKNmfpZNeGbNWOEfh7HOSIm
sMcfYRnAaH5vn+zxdSPdfpbirsI+J0p8JZ58DrZjuW1RqZunJH3JKRoy5LnBbo0W
S8CFVx7XTuxb0EifHvCw+F6MChj52RKUW8qMRYfEhQ7jDP8fAV3uo9B+Xw3Jb4XG
AV1eRMG23GMDMXPcNypl3WUXfvEW7Ee2z1ibQgn5/iNoXkoef2Px/D2VPpn4Kl0x
frW5ko9dGiH43aSia4o1+y0w/6bHcOiYuJIuagUgJJia/ik1xMeLez7se2ETreCU
98PIl4KhCH7aGUwQ2zWv1LuLehUopBs3UibcjshcowRwtROa5CqsbGR3Rwfgi/tQ
OS/2wfJIZB4Wdm6tWH85L3z6X8BEZaKCdHYkAZB98+d8uXHYgcHZ04w+pr7jGHb3
QzWzNaaoP6CqoAU1qtSoZRHZxndO4O/dy2oTf4neHUxQ96ZToxWLNAMaW7flsKui
j/7j3NCcC04BOcTbHJViuFi2XeH/Lj7KV3PEDHwh1OLkQ7Oo5IEcqqKjVXNazGN+
kZi6IgvISHg5n1yTHQBBgtzCG9FqUKJKuDVnCXXSRwIKv52GxJhE0a7pp4hSRNfQ
dKti31QBRw+CKruOqywzmYGN5Q1QC/m5RhMlvH+bVG1+hE8lylMW5S6k/EMfD/ZE
6kjgY4MNvveseU6ij2dSTNyUBReLZRu+O0hca60nS4WtQGbHEO/vsRMBy7lcq8JM
EaG1va3GgzAjsqonAXDu+OMP1lXVy5o8ic8buQUsTr3xAZpzuX24VihC37ejKAnG
vqicntLVrqmAu2NPaHhR18mImNSkYlbn0EZYwuMnFCAufMwHinGR0ZyXzhcSfuhP
2oF1jV1+c3uMnF4n+UI6c+e/pn01STPmjBy0nMtn8Y9tmIlGijh7GdfpoIfqK0Ak
dcnluM/h7sVmIT6Yew0MrIGZAJVLFPxorEOTiRx5svO4M0HP5nLAv0yU9W71bFeS
ZYxHdP67XKQXXQyYbyaqRjEDNpe7cVdORC7feNY64U2X2eWlB+eOfQ4PeI3uNFXN
0Ubmq54LM+kgmjVlel4C0KpzePb/XMoAXQd+9Wd3ZF0IXALJuqTCZaV0fYvp4txr
YHvgebqytQcsC/zwQAgloNJOiTabF7nHbCfL2PQs3AXURgFbyLSgBLqqf8fxp/Te
rqF/CWWSi2ibCeOy1wTyWWO81jrEDPVRQqLbvgmNdoSQBDPvWWTQoobK1ox5dRQC
vxulaThmbAjWSRUPyQFQz3TwOPGGhdZY8p1aunTcM31F7tATXbPOC00dQg12iml6
21iZZIIDhLMoyQDYzuE2bARZ6xi1CRPGSVpzXpzl6QicSZH5k9ZVwLsUjJxeK7ps
+iNXtgFPJuVUQx/YAffOA1IA1J0mJfnqQGw+DsA75VDMU6emKa+mT7N7Ga0mGHOT
TLLYAzGSg2BFnfTQL/6MIFgwagk91s3eiKLObH3qrZ6BS5E+WEDEk3WqQSETAVPh
zWSlbzGDzaQNdcJPo1y68IulyDZXJcrJHsHy05RJRmAyy5hhjlvP4o1ngb6R2Zy0
ehE0Hxo2XlC3+HG4Ra1K/sN8xzbEfDt8yyhylRXsnEh9Pn06Lv5DpSrHrzR0O5eH
9FqiE3mMONWsj/GZQ0N3CebOlxkCRJRHm3Q5UsnQBmFxLANCz73JhiZTFngxPfW2
rUz2mBRJwhzwIk/TWqAqYOMyvV8Ur5wGmN07pozCI8GuQfMDGrPiWeUIRbxax8Mv
AIaPomv1yWD/Q4Zr7zy8a/gWlomJSCy1iJKqP9yboGguC5ttpmvSHp9pEnmgeKQw
cjjg1PHrhPR5shXcuQur8fubcWbhrDqa9W1/PBYfIkO1eMJ5v0CQ5mDWPBJvK3IM
Eo2RMt8Wz285DqrQUjOc6opK5GV1tw3bhowwJVAgHr0R0dRsISFcbTHuGtByrxLu
ZSUrAqOcUuEaXtup3wcPxyhD2xXaoCBx5xDPhPzvMTdo1ApuHTA8eHJU+LJcFpu9
DsP5/LvxFfUlt3joKl49DyAkmcroeeKRrQINq8WnxV/cE3MVVXbRkICaXjbS+fwL
aJAUE5Ch2czOiRKTNN+HrTwtHGKWfwnlHelmurYikvy85hjsAfAIRFWL1N1tvu+L
aphjXBdahqZ8gKgHHGlpNP56R70QnQfRPTme6m+9Hj7Dqq0ueEAOjgUkz6VBaAj3
X2rJKMCl1c9dRkTjKCTje28ylPQkJWYx2PgGHncFzdsddshzc3XiXjeX18oInLUK
dghIWIIgO18YO0SG2cHfnfxdpO9XxxlubZ8W4m1qGSC/T0ym00Fu2ztroYHtVmcC
0g0OT+bor+kHIR0ijDg+n9yhy7nAIbPdotPVC/KjosurhohG7frgvz2ODVdchZ5C
Rhj9bC2nFA5f5ft26CCgewUbY33ndNaBxDhYaS9ryL5xvz4H4fOTQLvvJ2ZEXQLI
1OinRtPAjoIH6E1vLjX0MBNfu8kZqg9hcbzJAUg1twebZyiJ+Wg+m0L2GLqKVgG3
DIeraCS4OdS7BBCcsqAsuJWOwNIdgWe4gNmVsTBgKYPSPxuFRsGzz08BzGgYvx6I
cEfGjU21C5xqD8mQ60mVrgpUc2rio0S6QT+iAig8CY313moiG72zCANWBO2NmjhH
pGn4eN5sZtRi0QVz5x3vTSV4t0CP417bE6Jt0lP8WLAy74nbZnvUIODofesD6Pw0
MuuTF6VaAc6WZ57ljFQZ9wfYVHiNmr6IRqm7vHxdwhhHzlwcal2ANTNldY/RU4w6
IxuM8cydlW3EgR3K8n1rDFA7WgqTxuSdc5S6FyPpGNsG20mbyET29v5dqxpkzSVY
/JDRon2N3+XV+ANbJqwazAfaFYcyLU8cfA8i+hgOJAqGEuL6ViUnddlvjFBmfEcG
z8j7NFfojP+0U4w+9/93MJFccCEVobAuplmoLZLqnQPbY5U+fsv8u4610VD13guG
aHTkrw0CpCWj0v07WlH+IVGxLMJtdzHwAjvnRQYqpbIYgUKhPARXBqhl4je67567
+dca78ydgHvM4OiXeKpR44GNhxFFzxkgjB9MF9pD732AUg/SIz4WrJO2pzjzI//V
kayeTb9uy8ij2hWInHI4PF2QnAeopuvyI8U/pQNV8o6nAT3vZUwj6qEHw+HYjPh8
fxTMfxNi2fk29G6oylrPOi1nsunOU86S1ZSO1oM266vq8k++OhleRVDnOYIwuUFg
wXtEzFJBud4S3P5AdjXvW4OilrQCsnJ9hr8YhoWD8oB4pxRUMGztXi6MJ0HaEk3T
hkkpeIuSwFA2ezltePikNGDZfYFzawjhhuUga8aRzA8l1mo1p5WvjxcK+OX0KsTs
PKw1EX6lCGyNQWEKQcbQ1DnFBIyWxMGTW2SDDvpabupphefah8J8nLAeJApB1YkD
Y1GIXJAFjW1SWYoqENyzQUdNC6u1nUIHsZkhKOpVO1UOzXMWK5b96vwCvnMskJMz
A0n1JXLffhLTbKIbNGBh1NmW3ReWGVNhNVL8v1Ah266GfJdASPNDFDwidXlo5G4o
HTGqD7zcAxZd2Um1fjYv9WrqlydJ/Ig02tZvuQYQJq96mcdHK32YI8Q7BmUhBLW+
tMG8V/JhSHPL8eGB3O8/PWW6eHwy/8oBRxMQe1d/NMNygDBQqyfQiRdIJQJbnTPW
O2kaGnUkaYF0GtjJT7q69wofvTHAqqiWq/el7ROf49oBeVmtlJHFmIsWoGnVyumu
SVvJ2EcgMchjaeRdxngouAJqltwd7W9fchVg6cqmcOL0/ksWPVTSfczRBTfJqNDY
SLfAbucZebOKk6PvMNev2BAqpMHuY9uxe1XL+Gm2XQb6fkfl1zHBx7Udk2dXnPY+
qmTPrxJzcNkTo+XZuvmupkU1nJHsihXfnJgBUmblaMvJ43yU97COBDQC+wjrcWc7
Nv21p/n5uiMEBP0N8xIl8hz0hzDa8b8739Fkh5RKTobAhDd7C5glAsChn3nTuMT6
laVxtmrfBs+F2YCp+Em+i5s2w2252GWVxj9e1iLMkPtb8JjIzorJ4cWJaCoaO0Ff
5YBzSL+fKaRjVsrcB1Wc5/JV4kKM7/wRfTjoh6GbFfNGfNWv2+oOCsU/yqZdPDvG
Ezljna2PEl/6GjpEOLc3g5e72Oi9kngrGm5ZXpzWsceb1/Sxg/xCYxaS7h/8uwhc
iHYVfN+OvlbRjyrQpPFujhLGl1pum8O6uMgDuMY63K0YUZPyWjuTnFjvwmnOyeNX
oL4GfaPfdKVM+fXIK0CYrG4KCl4RXxccrDq+VMmXRbpp8KDZsfNDL/ssnxBL8Tlj
zbXKSBWBeBPxuzk8l/69PP7OJPZTJbL3CzPZ2rBFIr71toH13FsF92lBbCD2Iapp
JBZuqwc/NwHRoDbKpMdorUe2DM+ixxTBCY/UCBuBUAk5GmemOXuGL7LT2V21bMkL
05jbFAIRf0wps9V1nqo4qnpCsVJAL719nC8xvRIl3Xlw3+pSx6oSkIft1bDwYQ5R
JietKK4IJeg3OfA3TwvoLd7CUeQB/GAicSk3gdE5OFy7Rj6htqaPnwwjhBhdlLe5
sUneMGpENVlIIczz69nwj49HZvD4pWw2PrtG4r7AIY/IW+JjbXUphjy6ibZzf1Tg
SP6euvLU8XsWFxwidthG9xv6u+AhNb8BPG8+dDkU8gAzER7e2DIgoSo+ITAvFg42
7NYx/0QfwNmeAY/J0XwsYuj4T0+DHk+C6AxBtjrn0jZv7zFS04d7MKO1mhb78hWa
juAJP11aFEuRZ/P5vAdzdQVSo5ygY2bLZgwrPvZrwrWa+C2fQiMkTYQuXuL7cZk1
Ck3C6c2nsak9/mYPzFv2EpZVZkISsD95e9a1c0eV65199BLeNZqRnKlDXb/I6YiC
dyFP2GQdVhIJtJQsRDCZ9FBTEM4IHl3XMAdoTt4Qd5fPS+uwUYXCUmI+hZsR4R+T
s4O2Lws9+DcSdlj2+t09eHh/sLhgbYroeCFowwaZ4eZaRSSuzg/RMrSKGS3sFQhs
akOxSqwQvAbtNir4KO8J1cay8kCm3aaQbxy1FwD4/NH1dZe/YRD4XKYywwodnhbU
Bgl4zYHMMFkKFXtRsbKVYNjoHu/xm7b9Ydy/zzJ7PDuQR94nTGaiiVExrVYWUWPC
HoE6vzKKHe5kviCWwujlRFD/wbGL9cI81VDgUh2tDh8823WNrR6Z3VfhQoQFUXVp
869diflmxCWSVSLX3JBlH5gwsdiAFsxpxVWiR0aAxJKIFDXTrRqEhEbYApwzXUgH
1R0Bf7lNdO7gObpy52e3aS5eOqDETvNMFO8425cNCgWDMqBMzxNB1Zp9Ai3A5Nso
zdLvWCT9RF2f3A5JGnmU1zm0ENQD1MzmrFAyPZdMe4MMKaLWAP5C/u7y5LS7XiOV
VHgawIm9wmp3myhA3IxVaH9kWKYh0JfFQ32XEgBPzxLBXITJuhhZ4fd2DbCKmdhg
CRCbjQ1cV5gfuVa/5HVccQXHOi3yMvd8UBAQd+CYu+Em9OQj8QTkbfw5qGPLrhZc
RHugKmFryQfX+FQec+ehKhqQk+NrYEdaJD4L108Rms6lGjHKMuaBNUEk4kGZ35w+
y2DxmfkAIAP4QELz9MAeQ9h4B4DWTW/gBTHdHMit9yzfykSt6XFy10l9h46h2KaV
LQ/mbVduJ5z4JrJNY/pWRYjYqLSj9yLqB9obvAI61eArOowOI65oOepqvLE44E7i
muC1K2llOVuYqahykU1LrLkY3s/GuBJjZ/RGQYvRMNQzm4uSGimz5WTrfaHhJcgO
PhIZy1mGHOZ3n/M27K465uQrbHwFVYEoBKSo5aNV38/O0yn0Zc/Metu+XMn3nSkh
Rp5mnQSZqQ3pj2at/XKv3gQQqpJOV0Z8XkYaa2iV2eM3oENySSFP2YOHq+Qjkk32
LqmEg5RpLr/sTtA7ckn3RUSDnE1WFyYMYKNWnFoD0o/AisZVslOXMmgkRU7gnQKu
MwziOFCSsBnMQzGKNTwZ7WDKr9nd+DPKZqeQZae/UCYr9goL+VzCf+JlMM66Qz1B
8yY+lgOUbll/iT2uqjdehdKV3BCM4T9VVagXhADZ3MOL+evTbOSmgBZn8VGE8NPn
Gc1JVs2ecOT9EojcDH6JUnFAPkikmmQONlFHiMw0teYvbrB3cBoMvc9ZXNi4f3qK
YWu2oOWf+fenwTnm/kN2oIo8S5a5R0+jGjydGD7l6KXbz9v7ZzNLBYFN6lzquAMn
ucUcNrJJI0Dqrq+f5aGboU6rx2GOiSbDqmOMv0vhjWriX+k68B6J3hS0hle3gxVk
dRwL5SqiCEe7st8BwvLLEtWLKzxmQMRPMEYnc7Q3WRnyD3zqUZ64UFvR5aTPbLAU
JBH4c/ILVSjPAqhNhwG5/fZJtQH8v1Gv8t7/7h5BJ3WwoeypC5CnU8oKE6t5cXVn
z036POzA6racEgtxhFaRcdziQM3DuYFXYwWEPqn6ObRvSof2sXI/SAY79Klah2hd
+1vdAHZKtw3qQaad7qwUj8UY+9QoGmk3eu2Lq4Quq3HZ+OkVkoRYYI+Y97H+NMOQ
rL0bYyQ7u554raXc30d9nkqIRapU9RX1bM3FaoguZnwHDEGrACMIvJtA+eyANPNm
yfKc84a5EinGQLDrx3hoZHpGvCqDCVmzPHycfdkxz8X8XgPg7Df9Cef5z0UxxHqG
Yh5ivMbjv7qyFex9vi8U3KcaPa9MxqvhEeHawOQhtnFX/40bOy1JHsdkoHSQ8jHj
2UQEeq3LriEv1sT6fz9sVzhO9GTaNbjH0udjuaUlo5nTC89uNNTMVznNhqSQ7oB6
5qWbCr98PAHdfU6h2fp0G4XOLNXHYh4uuTdENtAUjKQBCS9LBNAadvTZzmHrt6OT
dqtjmoI8tHJ33qbQfe71KPW0sNHuVe4uqN/YJzOgE4NDssteeFfoeYCYVUaHK89g
TO78FLm88PdL8yWK3IpdnNHwOcQkXLCt56z+y4j7XcUWd63v0Kk8HUpKuPoHDhRG
EUGn8pUD9AdgzXYlD6/IuHDJ3uFAIXYe+5vXmjOYGwmDIp4ArQvP9QdB0vWfERfs
ZNQg3oVNQaXkT91l/t/95Hfh7GdaCJSNieBloMk8fnq0vw2u1RzjHvb7FivMg9si
5jMXWXefzacVWZ7Rt4jiqynYi2dCiG91YSvDSGdqSwqUzXQaKNgTDpsDz9f6HQ+R
mkx2ev1cxkmf8HKUGLCq0ION6QOxJY7tAW3MOICCK8hh4G8Aynhn0z64ROmY8oSM
ZgK0nvez45a2Z6fOGI+GyvATY+kTsNM1aKaU/Lm5zx3lp4u01bmT5L7EFBTnon5U
Q64+aPK2D5c5A0GKdzKsQ/NMIzS0dgC6WqNs9bP0VtyOpoVp8oqdoBRLcyle9a2Z
Y9Kn+uZpZOKIHFi6Xo3F8pgeKEO1i1NRP1WSxzWi5hcPBVfwu/3E61Lhpyu+2FJ4
imyyTmgK2pkGPdV0wX3ItDL8jQtmHT8Cc/Y99HFzl1d5waweevdCuWMyIP0is3zq
WlbZoIeyuFulV6i2qetibnKf+v7a1UfZBnG3dYQA0O1TUFb4AJj1wpwSu96EPliu
8S8vj821+3XR+mOUm0rb0tx/6NQM9/UnWaFh7jK0Z9k6JQxDhJP89ug9z/W1k21E
HyFcaUUMR4SppBQQ9P0vq/+1eMNh9lQQuch/5YH8oR3PGjcHq+FqtQQk3euwWFrI
9aDG4xEs3mYVb/mZ8pIwh4DzU3qPC4LTTr5EZLf58coYoR0gbauuY28nlwByWSJY
yzRthMvcNqslz2y64EdciTEtFPE5kBxisWLDtyBAEBBkxTZMHxWMDfZmuixLS14I
OU/tCRz715JDdFaBt3zxwX2HUAPKXW915pFFoYVx7mDC4/e78ThUS4IaojkxB+8q
nu+46B742QSFbaxjOZYRidMcljeZLeTSjUyCO8fj6fdLMS36HJzYwLa8SaPSx4Tv
cfXa6mJFwtDf6UrnUc5nALZf/YdOOM/iLCtkunSwJPYdKQ9ee+RDbavwo6C6mK3r
BFDOt8DAYT8rzSEb4/KRblFh4GLacp0K5R9dV13e3zAKg7f60z4XPzt45xk/hO8n
GPbji5s9ygebUSEK2lhJ3nj6spwkpGS5JPQ+7d08uRoklMHsAYwZSmmqj9y/t/ot
qAGE74M48QzcZrAafZhRY0bfJwNAOxs7W26vyBaQctrKFScs4tVnsNzd+5QpDVkf
Q3hZbyGpXHBjE7CWsvQSqDQXS+YOuIXaqbChGP58+jG/M0AbRTHP/7XPFhlPPl52
HNkWgme7UwRRFDnfHG111PhPvqFCUtzsgtVe5AtZCZdzRp0yqvSmV+zJHMmQ5jzM
VQFMW48UKf9O3q755uJnX0uZvMOSoMrsjP1JYVvAzYztBJIXyENaFQJIJWqekeiD
1Dq0zdh32oU5Gz4SL4YoTrP9fQqjwNlFqG1PfbZOJzgx7AOy3J/Avdsej+/9koM+
2Q7EJieiaMEpGiHovsP+1KCAH8YjxOEbXELAuv2q/l+yiYmYXjy3o+C5cW5K/lXv
j6pUw6R9UzNTAZeEcsbgEewtyKgSYyymPzvP3ODX7solRgbK+OJ41mH7wzL1tAjf
+fAUwYPRcGMx2ciEKepkIeO7FOTY9HUwAIHgyVjoRipR9HBXiTJBl87FrQdgnlEj
ZsaTWZhcacK1z0uYNwnbZRcoszFjGvm0OisxpBIO2wIgmGnkWyyHekKzb+BC0l0P
fbf/qKhhgHubAmjlWV8jL3xGXWvse5qcAXGqzINYwB6UR5tFnpK0LlvilUsxM6FH
Sp4ilBECw1MJUV5A08nsLD/+JPGyIUYr1HOKicyDWxmlZdAlEWYs50Mk5FE2HLZ/
RuuSzZmRHLo2T8/l59zU0yBjbYiCuJpnacm3WPJxBaaDiagy8e+My8p2SHxAr3ld
jGXcsVhzEBZahGAQNRrqN8bAOMs2HunyYuvQDOdAVY2BemGBjCKr1fEx1ICC+o/8
XjX4ecOf0D+Lva9jgEIIisTx9jxwFEct2D97ChfcZPUgML0+ppuGQx6KYl2Li4iM
kGq7emXWy8sZ2gxSA+9SfNupYCm4hReWn1khV4ts+lbJBOdewQl0LWy6oHb0ex2X
DZixDtiB1jhgL+kKh5pawCd+kYfVpUiukBJku9162Tbi+/q6Rtli/iBTDfkKRU2g
QfaXw0Qivz/FH/rDkCk4PqNq1yiiQ0Xld2SFpJC6latMP4WxT6WaOpy3FQkhxyKu
1X1tmx0lCKP1CCbPmeeBNcrznNsyh1Z58OehVumP1aYawcSXZu+oaohfEIt8xx9d
Ze/hNuwMgVhqyhIO0VSh6gDJOT122MikJs1X7iOjO+aPicoisPqbfgLovonGXyaX
pOg3TcBrcchht0NsLwmkqudzq4PWc4eMaURSFrIuXtLvPMD69PMMs+5hAbeDuqaG
Bg5wPC/4s8u0JYXc6WHsFRX46ia34OLuwzs2LSfrjjjn0Pw3yZeuVOjCeSfOnBC0
a1AA3U1Ey336lKwqVtY64aqb9lpR5wLqX1/PJLiRg4fg7tMeLw+4GCAog1GUOEQT
GGaG+TcOcEnSQRYyGVNVU2N8MNHXzEpX08nud701976t3eKW7w4kVX5A2e6vpt4N
tLnBMjY6J/2AUl6XghH0zNbp5+JujDDbv55YBrFtsf6U5GWp3lGtHGHyhg7Sb+YJ
0TZpS+cRxnav+LeZ8T21s6bjQOoJGNX6uOHYD242ejh6wrTEJa+bG2h6U5WLnHnm
7SGKFcUJUhem7rysbIFD5L+6fc1NuetHA0SCnDk3CAUEi3xzKUqUz5wUB9bM4VX8
NrhqOyIiBKNWcNRgYJXBw3qVFS681vhzSkcTtcXWlWvVctr7pwku0BTThKa/3TD3
dIORiztVYLP/tOZjkzL72gvhdb/jPRYnrBKePjpsF0tsk9YkdjHIy/mB82CTGvIR
PN+uRj8yzJChqJcDQ+/qhDRzcISq+qBkRYQ+vwOSEZ1r5AVmznP87En3E6SvV1hq
jToCnpkxQA5euy34QagDYA+hlymcGUDn4OnVqneFKat47eKhTSCy3hVMZglDn8BE
6p4LiMNtqO9a+8zIVpBeiuGvOcnqAXwfBayA8hzZQuJYhHze0ip9IkNn+QQkLP2/
Ft4uGIxum/T/RGf53Nv7CHn9/I7ECSqRicqwPdTmmfBKp9N9kaxIDxbrM9ReDtps
mTwvRVHi5I0E9+X3yRCZDlknsRWGLn5Xz0M/NBmx1pwuQf03MpbKsw3wU/pxOX8i
yjXUHK+lavuKOx4j97qDyiGTP/sG5TBRJKZG2B1I7I+2qN0rnITjBXMa5Fd59WoU
N9tNls/AOMjT3vOtDrHl6YnTN/xyxaxUEcxAQ+n/H/DgrBjGYGrT/TtKx/RxuYbK
AiAhryQsjmFoUj2U3byWxuwMVx2oe1a70qCYviYx6AY/es6XdEDFGxQdrG7z06i4
iX/BL8YEyO9r2cbn4KzLgyjclTNiiZ0QbJ49PnGOGPyvHcq0lv8cKBzvP//vbl3w
mWIfLaCC36PT49Sq+xpDpKxst+uUyum0rFTlIF3xv6OCWxXf6A3pcFLK1vUHC+PX
pPq1B+akxxunG5mQVx3TjUG1YaV39i4ExvfC5+rSZoHj1LR7NfArrqvG+lK0CY5r
pNLPy30jYPHz8vtRnnO/tgXQXTuL7gNe32h6fQZhfxVHk3HlZovXL+89RgRfIkgq
pRlT4V584BbhA3j6ApDDjku1C9abTXdQDdfnOZSdE2iVt5Dz2GiGkfy1r6dYLYDI
pnLYl6dwjIn5ny3/BMONWIpUbeX+5JdLO2QG2JOsvE/zh7m9LgE/0VArHkvmrGFG
jtihJ/veYY/vfdXwSn8AUm7nByRtnZE5+B5SgYW0WlNLOlFJudx/0TAf8d/Hqi0Q
n+tyIGvSoPQcBH6YUAfnGlBdVhwLeEepLXb6lhhd45iT/J1Hd4FfqvOkYDZ9QSs8
p+G5ND7rjiB5QbjT3eouBfJzziKJmsEN24k8GFPs5wyXjfuyCc0/hWCGy5TlCzDN
Zh6HgnVoR1/eBYOF8/wMPPDYFsVqDDmG4jQJPEfX7LE0aP9+mf4dR1s9nVOoUXCP
u8nwBt/ndheeUPCSDpyOMg3xzJFePDQUwu6Wqezc6AlVezTwlL/X+Db8BZ3K5Rpi
xalMl3ay6YUxBkYyA2yssa/ThDT6ZuLgMvWWByRFOSjUqNhXqCw34zm6QdADpIHT
fqZYkamjxAmgcQx2cOLx1bK5Wkp3zMdik5QmGnmcRZm4Q880WCe/hcmXoCBsn8qZ
bA91JgLozCetxl5i1Co6AzwFlliqlt/8TnuLxbUB7kHfdSwW5VcpVIb2R4KSJ/PR
sdpDUPRZ1j5pJgCQ2+XTteS2f8Vo1Qvmb5U9/Fgc5qhQ0M/ZWh7GpfB6LAfQL7Xn
hDVaPSUsAnjDMdLK0CFrJMBDjOLu8FjwAzrynqaCO0H+w2BUD3yRYveq+lw9R657
3Ogi2RjymGoujuXzqdkPNxVjP1iaNnr3amzOhfT4eLBsfJ9iUPdAiwKNj/xoYUF+
ihXU1ssRvXgLJW86mx07upYd+O9U1y9NHhnYBFz4MM5/PPspuFmYGXPYtqnW4gVo
EgVX5r+wGrCBlSvBLgSV3P1fj+Y1nKrowY4Kw4U9I4QFtxW0tQz96IYKeQxO3Y/1
su+ftwJj5H4aVupagJimvScYWBIfZAfV+lIRMQlYZNJXPLBuayNHtdpdvp4nsykW
Ru8pCtylcoX7fvL2nIjsHjMmfP/ZBCxiiuD8KNsNyL4KjRzpTCxXEHPm0X/79uT2
vgLjvo09UKoU0snD2UC/293NNGnw6jNTStyWnSpEHc2aLetmV1nOvza6ijoKDku1
ZabQe+XW4fTvQonjZ+73PK4FEnsudVHXNJwUqG53YSQeGbUlGLcZ5CK1HpmmqYAs
xZPi9Kqa4Eoo0lPcmxsO9R/rlwN+3lv0WV9VwunbImG8DEdb4FMbolyRwyqKei3R
XJMORiFUmgFApSApmWZK0E2AYF87T3Jpmace3Qi6UbXHyCKg0XMgUB5lGlvbwpDN
+WHRnJpVLNs0h3pb0XLWnXRhKgq1HdoMIvsu25A+80uLSB8sLBF2DcUlJKbBsYkT
4TjjhITEyDDcCc0ATOZ38wcKKtRlgaaw2Dxh3moz60ZXwlYj+Q0biCMmYdmrB14u
Ikq4rcF7m90qzotwCj50v1MX+wACI/yTvqghyAWqgbuTtw1Z1u7Q+VUYahdka/E3
wXWiVfTOozhTmQvE68WsBtuqb3ev7hsmNh+e4tS4H9NNIRBpTGyIaDJ+XvZjq9Aq
bvTYZlEx7ECqAKGdnbg10jpFKJKbuqN3VSCWKEP7JRskv/FybRTgBPgO1FxfavzH
zwwKScin3p19D4Cw7RnSIRRZOBcK0oDAdALu9bMLRJZS62kZLwGCFwmLiEcNHcCX
BvMYUZdRnV/Xu/xQpVbQ1S6YxDhGoiZkXxbx0lg/F1vvqtX1lScfzERD3/P/Wz7L
itGJdFGlJR+36PEQweNrgbe34aYZwqRIjIu9r36YZlMNVDU5mAvblj6mu2kWxB3F
8Rv19kTqA0DPnmI0gKdsyGbLuwn5XtnYX3OhCNMdZJ2UiH7EoZwytXfsddLnc8mc
dn+BLuE9cSVRUKAU6XfTHUAtIP9uGZIhtHAuUgqnqoqox1WImr/Zg/tbHoeDwBaU
AdeVHCOzBy3NCXFLAYpfD9et986D/CtnpnLpHqVB/hGYYptqEwSurjlTmQv8KN3a
KJu0d9q4vGHn8MKgwUAos9fPfihxEIx8e6OZExdHl3aI7WBs6kpYQrieKv5/ePNr
/ojIxs4i/BE/0NBphOFvRbuQTcBmHEt1evv0P/WuzdVtI/RaTmfqtYNnHB7RfoS/
qsJLSOHixFI0NWlbQvYrSnXvDSHSqr2xEdQQ8E0fK6RtpbGddlS/wOPvUB6tjJZm
mwpwitpoex/QePsCPK5quqNuWnGDRP92gZLnfz+EavkQ+J376Y9MrdAhHSPVXC87
XPEsLwE80n4AeFt7ni+tx0EtDvPbkLSrAfxQHASt3VGmI4Wg7ZW+hkEEGo+NeEvq
UojgwpsdinLq4oovjokng26bhcaI3JRtCildp1qj9ZECn04/PTEHw+RKfJGo77yF
f0QHPrwMc73dpy11AVtH42CfGlPONgr1XUyg/dC+5CyqmdVXojYwzcPgyZ6/FxQd
D9UoLB93XUKK7rHzBsE0IkFkt4UJx2GOxHJzB82YTX/Dr6tZhf+v0bqQyInCQJzV
155OX4wms9SCUCSOfFXSZK5bC/kOcHPpuRh41v/Mw7ifGdNXE8yvOSL+uwPOKeGY
HqWGLsN8iIU8jKS6GN0DiI9WLnwLmWQazzGGmsmPGWHP8oVrC/lpCzhZgnESgBi5
1zuaSyzptixvuVc91XYNBBFLsh9r9vPTyc/fyHkgoWfmywAntV9R6Q6UcOSaHN9Z
80e44axR975OVigFXwlARClhtfAgGWlkFeOaRMtgSFhnC7hFK/GFiaNhvRqhnz4h
j1y3VG0qhh1YGe+EdwTyMttTzr5qZav8MaUhfJPelCV2HwIAtb9oqOtqZig19Or5
jtbWfgg3N0Evbs2xYpoIx4rl5Zo8Ji+MOOxXNfqu9naAsa7rf41aCrVK7axa+ukX
bHIjzSAev+KncRZ9bdLdtUY6LUNLfwbqeSx1h6K8j7jpuba0t9+32sqzLsKshb0D
ZI0fw2531oT1n/JJIuXtC4lBFdiPwAB8dp96WgjjOFSWghrIXU/bA5TN3uWrPn7i
T6TDk1TnGXP78m/iA1gtI0vBtCiBfTElW/hlB3c+L+jGcZLqzulQub1rDsWPdTDW
2llWCc/8mLgChcoQsVeFytN2fYgRVkpcax5PuIUJdnpUhP9h4lAlNHXTm2QZ0Ojv
EnLjI2SHhGT4My1LFepWTOzAJM+nXwtEq3MnMJ+DLiaEZAEOseZgOhJ2eGV70f0t
Y+C4iewjb5u9j+tnOa+AkVW/B/LrBlojGO4B7XVbp+XKSV0Cw+KFs+LHmHuz34LQ
tnGwv0JzROfu+f0vyU9GkN7h8XpjfPxF+u3InIrev5/Atg56mAupvf/UupTeKNEu
QQIS+Bhrbzob6kdZVIfnTJF74lgavs16Q1oNjXWHTGyx7G2KnlWSwHDdVs85zQl3
JE0KoJLBOJzmzCZUKPTOGuw3lOY/9blzIUSW6U5ptJgm9nVgrmNTnmnbvIaTHDYp
yavU0UJvqZinJ6DwbLHjdtRIsW3DP672KSxdmpc/yTqiqvv2FrwvRm4h0LwrB/ze
UNw02NcPcy9W0ggJ7NqnFM4H6TOytDROYvKM44kuWZpM67dk6g5E1SfQB5rZT1yy
l09KcKYCpoovR4Juc8gKq2swaeQvgjM/a6uJgFBE3DseMdqo5gCPSpuTF9muz1ER
sVbxUpUxiyC31n1VAKGJ7D6B7SkdxrgpRjTnT9Mx/y1fztst3L0ygJWSzM9LLA3G
Wsx7b+Ef1ild8Rdr69wQiCN+LUh7PxKSvx/upGwE7eEiX+lpIAe823a+vHDXxZ51
M/nSlR7Y4Km9Tr4/ZmDpcAs/XGXTa1rNlGV3Oejyj4wNzqRJp7JsjmHuMSYvda11
mQdTiB+STVVRXpaTMrn8xsA3s9l1D/Bk1l0OHkPYfB4ycta/BWrZOiE9/aEM6FwG
tL1Nr5xG/aH1NQSEhnna3HbpOJgpu7W/rdenaFEj1zok/9kQWzoIbgWia0tQO3ht
VsZXagxbwdHOKgMlYrNbueMldFQ0K6gF87zCxOWkMudzis2JRPsuQd6kRSnAFovR
5/vbj8hx72O5PP0WKNkZFl7A7Xy7giXC6iPBjILnfQD52eZs2tqV3NgoqdKlPhJr
jjKUyzbSfUN8jdxiX+wrfGAGfi81/22gUuliw4ragCUZOiLtV7rY09Z9d1zLZ+jq
sE4L/NAlZaTro/TvztjVGK90EJSVPZMZziwKA496Zo6Oa5CiTPN5/XxBTBALL7oq
sMY9c7FbIBFidq/bGOQneA/QLTRksTXBPlq6mpgdflLP+czgwa2KWGmsDnisr9Tw
1OvTIuFxDAK6NKGUGs+GAELhYX2SIRL+eZSnDs8MUQcAA3I1VqOg4hnLTUn9FLIv
k48y6gS4MClzIdbSvdP7tDqxJohMt2bjc5Oj2Qj1L9L5fwxkwtouC7TygedpiV4D
a8om5P/VJLgfEt7+ZtuHyzJnm2CGj4i64DNm19GLrd/0jAFZqMXW2pI9P1UoUk22
9tUeHElQUlkYT7eaUSMCR/RVBqdcl3f0r/oBXHbpXLXoqOI9BZBuoaYL9RKR77e/
Rxi+Qq0jRJbx9dnIq+1TTTAs92NHTQnBUHI9vq02CgcNzLjoiT5v7B4xm/pALoi6
ZdtIR00Q9w0BY4OfuSGSj1rPeQC+03rYrS0X6FrkkgED59QuWFn0VdijFxtAhxUg
G1frDg2vLyl6DIXv4V9YwUZFKInBuT66aGHVal1hggrFBMnU3XmTyfoLo7KQgnOj
AiVIXrRKk7LEEnpR0ErpN42CUHgc1qkY84D5PDsDq7cGTGNyCTSFa9pvq+LB72C8
P6CAV+KClpF4bFU69Wqk1GnPSevH6Mjj35BFVtCOaYUz3zq9l1wNxkbtFVTM2Nlv
i3aBYQhgoqaZGu0Ysd4rUMzih20EZawsJuWCa8jdsRnclkU2s5+M0Vlas55OPk0P
iL8KCUIVDiQ1rmbRf7H6us/2K1x4liIfcxlinbpbMUInC6BJlfnF1g+SG5fHX07K
z7HJlivN9KwC697jzV9jqAwCJXcvxoHuR4lMS/CgNmZemtOXdJJcHveVpIi17krv
V0YmP/X9n80Z+zEKQmY0M85SsjqeNoImKy/kmzAHE1432dmI8Na8awLtn9l94+aD
hY/PIvA/QBLuO2TWK9tDApFnB5WwZiGdmphRzx+MB24FsqS3FL9ZtqgoMQlJOlQH
GeMsjdKyg2ZTc6jUwXzZCyRFLbEhyAyGklaJHxI/O7heV41kdHlUQjP7LLleF8nm
lETcyckMBBSwe4EzM422RkByuEa4HfeX9aS67So1NTLcr6g7OGoSWIRP4w6Ekk+N
mGG8KDAOMRS6yU0y1CpACcejIXNZVkz/PbjHELt8hDS5gtce/9UIZqf/Biy96hTT
iZQDYLhlL8MVmAyQ0QFaKk5etgHvNQRhkFlPq0S3q60JYYbeXn03wHNrKgKX3F0h
YFcZLEsuzl8jbERIyBr5Qs1OfMKMv67quRI+ZnatERFT/1OUZc1J9TYLCUsZwogE
4kIEf6Vd+1lYeLSFzZeI7L3FlGBlHVUgIXCg2vZGqoTLTjoSVnNxqlslMt0I+hlQ
DZuwLt9SnCEB97TAIBFAAJP/UdSOLg60+HGYuGtggsS/R4Z0N946DoLPIlgJGnWn
IzXjc5iYOKldje6h3tkr9xC8qDKhyhy3TraFJLit9/qyB18aOkgWgY43/zHbj7Oo
wa7GCG/GHpKk6HhYVivQ7ZCXighyJwMGnxWsUwiuVd8Q+m8TjkY7c/UjPesYjmZR
G2LhqERZVJgIRcxLcHHg1BmzGBg8Q1FtEIpQfDRWjqOrG7hD/CFnH8d3CISY3x3U
web4rhK6l9GQ94p66i7vOf9/TcCRRom7EZ3gSEC9Q3VVtXsBSjRhJl7TiIMsCAZz
WnQroupZdeHQzPdMOh51LTgLeYoHisFbw3+WgcdygCt46WzgymyC/nDBOc5CKhup
cCj9pNNk8Rf/Ox7CH1SBwmxPn8zjWXGOcll9pVJWJtV2ft/nF9tItf6N2nFvveq2
j2c3QmsldWPpvwOPpX4Pzeuyluu2RIso/y0PxVReDoe6k0CDes1Kjjy4ARPaK7QF
QhBE5aBkGGJu6LuQwW9ID6C4mjM13WcKDFdqCywWfay5wPmVjmaRGe7iL/Sqhx5k
CcsHqsbaGYqx5sj3X2axR3pY08MKgg34IcxXL7Jq/nIORs7Iklgo+2Cv8NAf5JFR
1lNyCKbN9epCdU3I6oSRwuUaPMAoA4g+9RmHgXBy3H6pSEBlq5FLY2Y7Tity1UcF
T4RoWCmK3nv/goU1EC9IgBMmKohVxAY6NUwOJrMRWDVOYcAPoQ+AEgxNMaUIUUtF
NIwjXPSraocf/nlq90KMl8AMzHKkp81u3hG0nj5hC36FqEmOPnsnPstZ/b+8dU8r
KU5VDH5oOk1QHbGK16ujgmDplbNzsoWBYsCz0+7jKFNmxAdtAbWbTkJn3j8VUTik
AD8PLJoyne6seKppgqYq0siw/7976bV1cghg379gf7UUeIVpRnK33CbUGP5eUjNX
3pA3V99tEEYWkbPld6OTOEhI2Yns/pNXc8/JafWR2327SUqUO0K/P0JWj93Ry2ez
fghu9wCztWe9aM8GAK2anwCLsbriYhQDTOeQMC8JTsu1vcJdtkspSJhWBozlLEaT
dQo+gDAQ1BTD2P4br1Q3qpAIZBPonI0mQEwYrW85C2ZfM0XSh7CecY9c0obepYho
joBQ9oAOlfIjC8pkN1gU0tcVPsXf4Fzyunt2+GhIpPo0BYZvIMezmr1L7suMXhqy
zY3/uoGOg/nHKJXomorKep80k2Zqq1UK+3ow2yRR7kkQIMk3m5hoT3CjNdnux6ND
latHN7jqYek6cffJMFKMeW7U3W5FgeR86BDnnC5270bwqGaITM0X+mC3WrYDCsGr
3CuN9mTa8kH7y8iSq529SeU9LSkOQLiSA6LXt/mHy/lHKM4Vq+vQxUl+Z/q0tXtx
xcXJQkN/DIok4Y0fJ94KhJOEp07JWkC20cPDmeKG0mlcyXkX9NnCqBcgQSnXwH9f
NO7Z+PciHbk9AbWQDd+Dap+RY17vTgAZC3C1b+TdjoJzk2HtXOlP90UtcYTmWR5N
+4clfHtfI7FRfQvE5ruq/d0PlexqHe1oDNHRMeo+9snrMuZMPj35QaWti/bpDUby
9+FdblmLxHsGrvUGQy0BiqyYG5vrG9GmnVI6JiH/z77tXxDTt+Gl+DIJRB6orHGJ
C4PhPjrUxiyWk8egLSOspb26IHvsbPTLfwP8wXeO+zsg2lPNVezF+bVz1Eeqh8yr
N5Huo6Rkb3pXWwaL4pA1JVVKok5zV1HfPJb15DfhRVkiBtsGeYsalUVA0Qy8/X7V
PM+3YPHWmlanGizJbmW7EAJ3N9h1iIIvv7TX/SF2jDorrs8Rxqf/GKUlTDxeHOG+
UWLnmUdWPsRM+D4cy+F4CzVPAISGXQKGGC6zUFBzBSnTiLQd9RPpBIJColjfSUTJ
Gvyh3lQg24GjvBrjROPL5P+b+JxfcjVmP9+eLS4GaC8HF3kkdp8Jk9uNo0ShLL5T
A6gJRASV6sldv6QBg5lp/gODhc2a0toYMe53aZliBPIlSMmNwC7rdeen3sTNeGSa
dCqgaTl9mRQPm2XaZ3CAgQHMXmbRKFdaEoMSR0+FFNkvb8vSg6rJW7/keWMO5DjH
HKyYyUpnY4N00YGQoZNWC/APxVXuJNWbSqgop27VydbBZM7/xfULv8/rs3ubvyhS
HQDA4XGf6NQSifT673Jbq9L1bACFaW7oEz0v7sFBwpdwPx6QwcnMHW5pDQMT0vD1
yOt3XN/LqajJ8YRAsNpI3+xdVEyKwX8B+j1M3VcezeLEgC3vWGeBABz1BgVQ639M
byOcN4wt/+Qo7znSKYu/7o8wjnuR/MfzQIKpA/dD7iFlfk57ghmxfarqsPOYkBD0
l9SOtcxftRpf0bTto1LNABtaoOcCWZ/SVihCaN+wTVKkwZ1XxFXlfLy8opClHQPb
2ODcWTEKMR48pzX7toamwtcCE+Seg91AMMzURCj9NKQQ6jzquZt8N2QSLBbWQQV1
6np6e9x8ZSMblArDDoWSeVaoZxVph53Bt7kVpA9ASiKtXNtYqgvu9s1lyrWe0NoO
nVuz3VLpnnyFkrPUIXhKmqHvTUSdwWpC/9J50nP6TzMyMFM4qHt1/tPORSALHFAe
05wlVMUI93o0UEYhOdk1tL+96TKqvDNUwa+am2v0SOxsvAB+ISgWd5w5H738vysO
0+THmjtS730KwbbCpnpjPHS4S2FzyJawEgK7hgFXuPbKeC14hHZ31kuSxKN8/jlY
C2cpQ067n7C9bEqaK7g+PkanKgZjazyXfOcvWHfAamJXbrc8rvED6DzTNt+mdGtI
veq3lls10T+kRXRXBDfNxVNZco8V/xyB/EGr42z6V9i0kD/PUoOSz2xOhRMS4dY9
bMot4/6HJScl5GMc8tZ0p0EuHOAs3xaa7PHyBSXGlrMzzG9oa1f6ZxGqLQLY2som
+BP48u7Uyfksq2UmtmSYrk7aqI7aDQg1KxS1BCM94Q2f6vJNeWVLxpUTw4ZTPkNn
a4ClIxXOy8GsDWMuaH5Z2TjBNk6OJpFFlk5tk1djqLP3R+FN/i7TKnQzM9eBzNM/
ZgjGJSjiDJQh3xSuM8emV7OFXDKVfnTOJbq7on1xMVP7el6us52IQXu7RlcHrqX4
y/wQtrLSNxRBuLJZ8i9WLRfv/q2QXy9ceRJOk1JV09mgirDiPH+P+QjEQ3CZVIBg
fV4Za9xTaHcPsBZWHUcXW7VW2cai1FekJHW84Hg6CIDof0vlYg3sTW25/ejWfdK9
mkebjjP4XcpIlhksxGsFW4/rsjOaRJFPmde+vqxtGNcJRmDnf869UWYBfRhNZ8Vi
z3+QYfheNjsqtGMRxjsRa09ZAdGbp5SmDuejH0k1Z3m5m/Rd9T4NSLxx1lMZz0sL
GHsy9qvCtrP7pO/Uso5LhxU03Sjcy6kgwSiYqAabXbJ7Ln7eICknYOn4Bg2YfJT8
7TkOPAKJJAj4v9iqWDs1Kmdzea/LsiS7hqKnsNZf/RL8agGQn0vOd6GJwenJG4VU
apokSIHWT28bZnRN9tFd0DbTUEOEXHDaQCnzA0q9InvRZOYBe0/dKr849zynDMom
H/qJp7hqj4m9kbrTqYNGMk+FyOntJztzwNiSdMuzpGS4yE0qSm5DL3ebkBfqNygi
aXHlmYVhtiuDwn8uJYzQC5mi2OGvakRuFSfFDHyvPM/5boa1w0WCosNpX7Ii4w+g
h1gD6O4GOKz5w9Qfm5NGo27EvoGFTsCPnwTCUxk8pWcp7WDubxHs9fxweiK3r+Oc
GAFI4qzXUSt56CARQywcqC3G37IJ4WGUiGipDoDhvYZwOdOzCR5PJaK8sEVtYe/E
bvBewiX8PYXHegg/nPTuIjeAIV7oDkcc93bg2xB96cggtcjHJUK3txzJ8cW7elWI
aSXANyLCr0LI3Kya1xXRKpT43FPDBXoVyCr041TWZQ8i9MgGiZXk6yLxaqxwaof7
o4FrdluXpBUlKotbL2l55EgBvtTQQeiVbLI3NmUHoI80EAj0DtAxoZinTmX2u9sN
aG48X7mm7I1XSKIm+mUn4e7Wast6uQeas3Tok6nMfInyBNOmOISPjM05j/Wk8x2/
2wzPdfHTCfWWyTV+w/ukbW0JqrzRM37dSPuUkkaNxy10prP179MObfMA51QUvU4t
0F/jikUC2h9yq7BX+sUOyLBGMoBl9aOAUSBJIPv43C4OHeHZm1CB5Met0tNDzmEr
qSTR56hySlEMiuTwrvp1UERd5JzPDKS1YtF+ywJiXr/JQEpM+nzBAXZHEZnUB0hQ
U4Cw8aKBWWmMB9WocF6cQFx5iXGDndO9L+cgP3HsxdBduw5gnA1QBdX9ZPk8eU1O
cFZ930yeYukyozhDRnhPDot0k0ht8DFfNSwx47cchpv1py7s/ApaNdi5BzZyIUTR
sMq4QZZIxmXV0n7+h/egXyGix6MYDWN01q9UP0VRLp99JaCZVVNotBlWMpHxQhVu
PWtNIslNjPlTFvnSqUiGfEqmkLbyqiwnwd3jpIVgQiKsmVVp2PPy4eXu4Rz93XAf
rgRFvXWLN8WlLwd+bIQG7bthkq8VSYIGBB9FCTdNrM0HS+MzNQ4fKXVZujPu1hMN
6XVulcooOrmQM31FzP3Yx2dHg/3kthPwcKuL/KZIYF5xft4vbLYfibZ2XekICpWq
O61J9GhFZPUvEjBRj1Oeuck5nKnRvbznvGqg7jiafTlT1c2SVpikGTKyGl7yMzEb
Qtudtd9lY9vmWPf6gdw+86P6CoU2AptHNZQ3j7xgpLLySeh1Q3LpuJb9R4diTKUE
gmUHcqJe6+lU8tj+zl/4WaqYqqlv+9hTDxkL6lAi05pUPGKR/63V9HOx1fNCk7ur
85xtInSpzrBS5MOFFesvdmZzp0vmV8Y/GdWVM4zE+8tD0eDYv8WofSllroZZwEzg
1JKxVPYVd1XUOGtIjZrKTjGZuMgCKDsZCCjPVre9qtlVHM1k81Pl77QAgbWrcl2J
Su0IUSRCOA4cI3beZ4glm2jFYDLCvp2dr/zKkmlSacF+3K3gMPbpZE6a2RcDrug0
fdV7jdrwYkIXMvrIr8jYA06RkCNQ+ASKPgLai8RfSRQomlfOTLQ2o/pHBkmF45MR
xrxz4QUReFRYw6lcFDOPht/Zwy4g01YaQ5gRbvSgdYcHDHq5NyhtLu4pOUw+BvZs
qeDsDoNqkwss10yP8TyWRJFAzmY/VtPk30k7QTN/4QCcPTP1dzzFKBhpL/Ny/d1/
KmygGhppQH1z0RLn/aEaT8cP7KGv0ZgS7Hfi6bZKXo5NnIxoa8MREomXRp15oLGS
Z7qSlt4H9bKyq6/jCPJ7RD+6tpknHavrpTbjewS/LDwdk6pjO/cS6wS5o84KHCfI
SMz4bz7C5mwYz/ILdOCPuc9Fyn4NRAm34DpF0oiUYxnQ7Mu/SDamjcP3AhAYP6rW
AluWNStDNI4Qb47saS6FL4aebXCXSNVgE6m4qryujrnsh5muONfIRh4/B34A2F/L
2oZ5ekWzB3qPAlYM8IslVGPgd6eBglzWwmq/7cKTceeyc8k2guUssejOQPdxy3Io
KDaV2cJopHkf67y2n34RKgVCX8abxosTiFJTyFgztLrKUJiWG4zdZVeCZtyKUZLm
bFncQKWuLbgo/6BnbYTpz/jyVTKMGvNU+nc2q/cBdPRz1Zo+xye4SxLV4rmT6sLr
alGpG9RuY8PCCCbC6WYvKOQvHcbjjbFW/4kn/QI4q5Li772KMZikMNHQV9UwU6Qv
VGdAvIogdepolCuVySiCduVivJ2R1/ShRYQsBUgsPZtWqzMn8xkfiNMVawsAKBkV
iwwJfLPvxGOpe7Zfws5FMRt3VQ9JLGjRw55lf59j6aFDMFbRQutgTeirHZvg9oJC
/XfG57hSt4z4mupW/rPhg3xrzY4udAmzeagkQKjr5P8LTZ815Flq4LNAymgEeBSu
Yqb+gQ7KGxwlOxTla134i7iU0kF7iBlmYnUFKRFV+ea8DWJH67DJZitUhgcvVN8k
SQ1jx+Sof9MMKH+Pr3wnHmtY4RpKMg3cZU+QzCj0j6mb3/ON64og6lh4lsz1M2Fp
dUNLf9LfbZSf5AaIqV+IrZ8ADmP+AeHnCosIA3h6QMOe1oRvx8QUV7Fr3YCycNtX
zmvi4sglIdwsdMPhwIUlqaeIzqhmaHTa0o9bHwHb8y/dYJ1XDWvZRNFMbPbl3Jt1
wMwyguKMrOCVfdmriS60B2cwTmZ+0om7w3an9tAI4PwoXRxuveC64Br78SJ5bzQy
HHqiP+KB3XLgWrUHwOinUMVQ0EXPSlL7THigwxf87LjRyXPJV/eJRTnBxePfBVd2
FC9+5+F66GOxMQB9TYOOj7VXpWBbQz41Zj+HV1GxZqxgExcy4qK1+blgcDm8BYVW
g3+i/7ZNbnPDRmH9Aifdof+aQSRl9yCLc8LhyZqEi2+OrTBr1lSSOiAPI4lav3hG
nd9fIjwrwnqpeO8YPaf4ASfGQycad22uPc7JNizBZ/6Kf8VIdrglCOm3jzwgsaAL
6QdW4PlpuPK687hKBXp068jt8JMwm3PUyHECUh7DVJGK2mDliOmZidoyFYqofGSg
0Bq7tPRxqctvhsPSWi9+ZDFGab053Tusc3DcbfVyFfzB8sk/ag+kxCwV2qHTisrt
CyeaP/0D8wGQ3NzYMV2zsTYiHsLNmQuBNXYxCyvsNf/UnPPTPrlF1B9it/glALDf
GpbvZFN8sWXwx4/GweNCSn0UlW4JYKMxWZshbkluS3zTLJl7O8ozi609PXuqyGAB
RKMC3/1YIT8/riysdXGALFGeP+NGuHuuICIhMOzLKmd8Uf1bZeHJXCgMXeoXcI8P
YLaUIwy987EvL6Lu/Z6Nxo5IboW5G1i/DqGlLC80ZWkisxpOda/gjkYQLTO5f92r
o4IWvALaQe7IbHrkRchpUe4NXgNkEUijXqPL1tPL9Y2Vba+IJYkJH++l8xbWm5CI
nuVdIPQDh9GOWuy6uZfuGtNwGMffvqKBeCIqyyXK8NX1hjLB4G03nDWBH24hvR6g
L+ctEk50EmlE4CybvqfrV6cXsdZO7dMM4kv90DGl7PeUA0A6pouDa6ZIvKbmFo97
TkQ5GCCf0cDID7Zy4t4Fmk8ni5HcJ1uHccqzYbL8TJXGp7V4lI4xfndfQZ/RPqkm
00gBB5l0XpkWLeTRXnUyugJ5BzNNS/Wjn6CnxMoBBIKfs/xRaTtUj03fQyRwAbC+
sw9hqLuPGiK5Q+uj391QEHT2lw1wyHwG1QZUaaWzOen6lG8q+64SK2r+b+kBtzj/
lXlcdz98wcqgkywNYeGazu7L93bnUPadyLMOXAji/KXuEm6oUFncPDde548Stf9r
5hxCFhlDpUxFNTaxFbug+6x3v5opDuZX1PpKU0weoTS9Ml3o43+pxY0mkMMAY1Nh
HBpMB9ldiY6xOwTc+z8KEtqwUd+Uj4m3cFj1Em2u7LRmpwACi08WIDcVxTeSEl9I
ST9Q8360p7v6M5AtfssIlNEUx7BRhpoA0leMSbxLC/OPzHNwQ4j90Vb5RV5FW/e7
TK38LRk2Sl4wgeZuxtSCyh1qOEhtbuFPbJ47TlLgu8mCQml/3IsMvk5TIfw4ZIGN
1GCND/LE9Rs6hofcJWz6mm9qyaj4WRdcHEcZFvjOmK0zv2lGnInzsGUActRFKm4c
/jVv9Kx9Nxb/zm1IPNLrqgFgT72jmzudBV96ngm48iDMLx4d/4NCFVV3A93s7Gpn
JEsU4RrWGr08Kv/xy/QF+XBZ3AfHPzH0YV4446acSRRPm38FKR+E1G35uaH9HBgv
9s5eWVc67/a052OCzO1EopfRjTzg5+uJXuhc4tmL+S4I5hn6dMYifcwzPRwDiX7f
Ka7agnIovUTebuz294B95fONlLrtNO27KFcywiz4YPKDP70hX0Htb4xe0wMe3Fef
EF/pRrOZ3ahTONsSdeZx4V/LhesKLNCtvUf2MHy2+eS24UaD6zeLG8LqiZ847HvU
nTHSnBFgGb3xQm28MCW8HBWQImPr7fWujZGNdYKq9NfVLh7vflzJqXMHE4vLdyoo
d+vFYQhFZeYiXea6Ino5yjUuY1hnBrKkL++INyqvStzUbwpmHMPoUwuBMSizqaVm
OPVAOPIY9yeL39Ar0yhYc8+9k5JoczBVc5THfsw4Ap/rWtyZKYWDq5hH1U51RqbR
tjC0yzhCzkOWLvAN4SDJAvrrcl7NZxNKcZleBnGHAOeQ6IURhsZPIMjvu7jrlpgc
rIis8dAXkfTHEv/iio+xtdyV+w2Lx7yHeDNd/zkCNJyFJIDnnpHoe8i/uEleOhqt
h/uw5DOznlz6rWbhUZuYRtFbAgUT4bKlguX0cdrcXadiSmA26PdfD2fUVZfTnHSu
Mr1rOf5d4Hn1zCR1cNKjBPwyYL+HDiZzJjQxT2xR8mn57Gs03vv2oOetiOI0gKxM
w782XFdejxwI/vRqjEb+4Ys3KW29cDkNpBzjecSFdWFH10O5jtNDpsRqTwo4a5gh
EGtT4namlkP+zuVf6fOHpciBMZY2pF6ATVoktU+aCtwOnkmsR1ER3HFSTZrx4ROJ
Rr5JN+R9/GXt5SdpCo5+Z+VvvKFCyqx6TKJZQkjlboFLSriRkkRWF6zybmFWGDlD
pMzDI6GX1B2PB7wkHiWX0tBm9sco6wqjUp9iE4ixIAHFSjZPF2i6oa4nlzqGg4u+
KFv+DpZPeIR6uWb/tEe7p/bjCY96QmqRZZu1OC96RY+D+Q/CHENDCGtkPT5nPHp7
1iKcb9/fpu9p5Z788o5mkpXG2su0QNqNRQwFle2kddAqvYq86U7vT1wDKlnfCNDh
qtMOE/qoijIdZxQEuffWQ0mJDgyNnyvqW1GjwQJ3N9mxLiRKrZp82pYocNqZA4iK
u/3QO72a8K7Xicmrf8pGXHzSTDxX9a+TeDKGyTh7QZ/4wWoc36wuvvVhfjptRSpM
Sn4YDHICdlMMgNvpIZuCfRiDNjkT3/ljqpN/SK9iSYTu8oZjl3LKZbovg37BSsOO
V6LO+CqjXnwpXfeFuylW7mdB+njfaen1Ntw+qiLdr4Cp6hm3u9dr5lfbfmU2j5WH
DgreAp4w9yNDJt/SiXzKKOW7uw5TPmqwq8JMOlax8oWO5OsK1JxSnqhiHtUU8UEL
VyAwwVbs0wnNeiJfTBOmTzGmKi5ydSzPNS7fPUXcsK34cIGInp4oIHTdiMKrCUYG
ussJw4urLKiHb592S+0WqAlcmJ40KzHSkOxP/8VQP1CD4GL4j+i+YXI2XsRumqku
wPhN8ua0H14p1DMCk1hJMlsNp44pBG981nVWeSZhy2AoTR6FUYHfYQ7P8zrTujcZ
B6RLxwlBGVuht6zvFejOZMhgL7u2VdqYSE08QbQ0Ye6NmDNHq0SM6VkbuJEhO9+J
gjMHT/pOrgPK6HfFIVtR2Acp9t08WsvejpY4TVSbgFTNKmzIgNeWkAmwHQKa3nXj
uIoLsVrUqQD4bFi+Q/QRCaDu2VE2kiVA2qahZoU2Lftn552xbok5kiM2xhI+OUfn
2ueK0XGZA32JZ5CawpgTw7XYoU34vhEzz2w/0Ih/sCixbyXVLSWaG64I++ApFJ6h
eu+AgMuFxJGs+B6WUK4hPB/ID5hv0eGjGpheqSmVlWLtDU466AZ1sQm5zM04a0N3
ih6bkyv5c6LOG2d0tXmqJ8KDP6590P0/3SofNvRKRQECkFMlfNa6IFiC6/kFHl3G
Xd7GH//icpchFkCKep9Co5OODrQd7FU9cxFVVhSOXEIGMmrsk679cFCoWM0dV+WJ
FNTt4lNHjBZLnxi4SuwYvLWr+ce83fHuVCPT/BHxq8V1nbA3fEec5sEZOmy/vJ5M
/6CkhZgcQiay/5hq9xEyCuSq5ej20R/rkPKMZRKfKUurcLAm/Na4RBKAA6m9ZVLb
VRXWf0kUicd49PF/4wp3Un2Gky/yCo15vc9nbjn4nHbsJgkmq9BV3N1CzNW9ju7t
XxAYp0JvTqhr0aklOyYQ6TDIwBYNoBWx5UY874uluT7EBTtpUMcLIKMgHCPJgc2D
1aNdB+LiHVl4eEsvqge2SorBwBy7zhbxf1GYI5wHJGJkurtcoHa363/Pi4rNdtWP
3bLzA/DMVN8tniuuagxz4aI/fomz1LV4JoYzHOyhpjWg3Fyjx6leY4PZaIQGnY/m
6YwtxGzsDQVeC+gcii4hIwucCSlnNAbei18lwj2bDdHhzfCgLYgJwRNbBXvVd/uu
JtrC/iDR7FRSCCs78hJV3COIC23uXvm70aW1cg85iLiVLV4+Br4/tZ3S2F4CrPeS
7J+S36X2j1nsVO/f8ljCgP0qfQfmV8tQHPozgQs/Y8tNeRD+Qp9itzDc665CW5GR
cM+xMcC3xfhl6G9MjQFr8tz4CxI39CzBnlbx5hetPYgI2YacKFAO52dsZotW4U7X
SBxDP6s8PgtVIPsyZKnQIj/HntJnygbeQi76ZKwZCsjiG5WrSZ+x8RRLIZpNT1xs
a2GOUmyTApn9waqSoLxmt0oQcwbdPSXjjCp5sZ1QIsL933d24rxl/3pFPz3iuPKW
+pWJvXTmRdm6y2V5DK6bfFt07fny2GZdaRT+6d5/avqX5GNbs2XPNIeq78eOruTU
4bVFfniiMQZK99p+S8BYmGgQymVTW1creZeUYApNtNZwxu4CEQkZ746dz0Uy5Oe6
QcOF3UHsVhPQ6S8FVXOFHufszfgYDBop9oMgcPIKMyTAdgCulhHkVgcxAETJyLwA
xjzSgge0zvlpKp0hF/aFImuBFvh+237VGOXenXRGSHl0z2OcWS/DYM7f3H21st4g
SbOuBK2QIcWcZT3jrljdMSP7eNPjboAxvo+HBXLDuot1KhKOIvTRzDGa4rzg6gf1
MeagM7lZS6ASKwtbZPFbAXvc8g58oorFNjqOWZuHZce5wt7CQlVasb9nxpFCaQHC
kXs0UjOPhhnlo2z+/z5CoTYwk2+kCnhv/ZJ6Mud8H63w5Z9m/vF/E1nf33X09otb
4Vru4IzuDVT8couDUyZ223QvFLQ1kZSUCMgo8skwPo3Lx2yLG7LoT3ZoBLpne9b9
uwdLm1910He52mXKJRwJq3X1xao2UxVxQQPzMkh+yP+DQx+o3960tshwTaBcZXIl
lIsvCGqPFx+M6dQeH+Nv/DmeYFXqtGug5NDNjeiS5K6j/41E9Yuhlafy9xWinL4U
GXptKVe8IGTGzk808O/HRfH/IVVYFEUDNqN1pRhCCwEUKrLj17V5lwhosE6AMszW
HLsIVtPwtigz9Yy5pfwmI6H3qfrhjcCPFIuIazjft3JOcy6l+1VHhl8ppmw8sZ69
kW6YAguB8peP6ki9fLlJfotLvMFHmPDvAwo/j3e770CvO0Y+KO6Vq/6DBMwmW42v
GkNZqQQUesN6pCe/p3WlwkV90Tms5ulFwCllRNANpTIoYjr76u+1Ppe+gX/TPLep
giFnDHtfJfYswhcTTQDyiSpOSFlvDjFB15byKYMT9GAjdmP94cQLU6N0W8rO12KJ
3gdfP2Z4x+bmUJxOfgDWzygTAN3GT8V9PLEiIzhsVvyXq59q9Jlqtz0nvBKm6D0M
je59m2et3Nkgu+cPWU/0rSCm+UoBIEzR7iNYEJsmoy6wQcB7ICax0HoGvxMtACcF
fhlu6KWgE2AzBj/ONum4qO0BUKhdBWgmvRzRNsQBNV0OfHwtFDFb6c47HY9gcGIS
YEe2wTOhLcqC0D7jaVOH4RdDyU6ittjhrgQ3cmX6oJC/AxwWchWOlpylgHVgpPGv
75IhF5ugmfHfk9ZSbzYcHfk/r1Ko0jmc7rziB2f+dUQ+pv6apzGh43jV4Bcf/jou
Eg5OLg1fbF9Z3cM7b+ycCFnCVsDLP4qme13hjqTfiY+h6ufL983WSYziIRfO7K0i
juB4gLfCMXS8QwaFkFjpaa6n65LshwrX+/Z+paPU2Q2SXYbCtoevYIVvjW31RoiL
aKjTwFlXEuSs847OyYIDMZwXik2z9Ucpa0aRhQ9qMnuI1wbLrjCWGYANGsPv6rjo
0veDsbp2sWlOc40J1RiMAiXhtWBvW3xvXtsf3E80lSPFuiysdtDHWSlcZ4wo0l+E
cb1O84H2eSs7NimVGRMe0llpIFoG2WPW83o1b9USeKy+yXytlWuPS6PEbKsSZzNi
UYBRWUffNilyCJbZ299QKFxy5W0U8fIP3/H/zT+T+0XMJvcoVO/onK1axGuicWOn
f4TKxJ/rjSuPdBXUX7QbLWMwogbir9ce33xGJVddMY+kyxD7Munc7mttYIrTggTx
WnqpGuZCd0l00h6hOFf8oZE9GTu45MsG8e6shRBjS9e5GSwM6xDsOz8MtkRRlADi
O2sxnJgoZxkqf5SGGqI4GZU1W+wU4TLUVPT4KeOx3hFO/gRhY3d5CxU/D7bcSZhR
gCVMhztnvPh4N9Lv8ZFvDhKQj7gzGtE9/5+f6clSGttv9hXq2VLMozAXWjWQzcmy
iZoQjMW7VLhaZ8lP/PbJwcH/0roHJq++xk76jDC4g3EIc7Yz76n9tDnZk9O54qd1
+O8e6/3AmGNmyCyR9ZaT9Qax+HUhmVIBi1uLfb8M4sF1g24Xo88hQKcQBsMOYI4Y
FMGZNI8y1FdGyiwMjbJcaPAIhheIeF1tgJ77Y82X3i+mgyyq2bflXUX+pc9McyPO
Zc0pYAhagT/5ktQ7CcUaLrQN/5VrTbV+jixBLq/0EySAk6BzED0NIqoRcrE5sJmp
KLw8VvfggwzcaYTuA24bxNx2vZeo/fp9j1pBrKPTCI2ImdVp9ol9tvYD1tzZmMbI
q5n6GcnlhBPO6jcDcW4KoKMiZl4iFiDf9/Z0AaR9X/Ou4v1VH6kLPhktibaEOWyP
BTUM0VxhmzgIWWSzm+3qQon65QHYMjZanhHvv6594BWrdeZV+bjYenMynUzprjpE
tm4vGPWjXXPpgRyoAxZ35UB4ZvvdDG4O4u06Ks3l6Usm3qBtVvCnC9WOMKRyOWyI
WGUWtuDQQ+m+Jj90AaqJ0Tp2HR0o3kLc8z44/hRv2SkPs5MMS1hmIUdjyUIT8hkb
SwSRYNnxm4XDI6rwr7F3WbZurZxJWcZaMosXKfwW2tzMIMahdDA/xTSXc+tmLD8L
R/8tMX6/0JA64WhOubIGP/+Nqms0lB1zi8Vn0cSGYusZI6NNB1pXGxCm/Xrazdcr
alm08lxUnXb8bUq7Jy7zwhzdKsYS1kWP029Xp5T1P9jecXnhrc3Xfrwws9y0MxzL
EibKBOHHN4B+W1MvPpC0V1VdoYj39PRdL0UB1hNZn7mkZpHAQuVBPk4RF87061UG
gJ5qDuhYAxaVsQJ1ychWO1369MaCx3GPN8V08cHK4SAmEnwpPy81dgkeu+iIfXqy
z8Q23YgZxTjpXZ7tsF8mPPVYu72px3J6QXEZaL+p6qNstn+sCDHjEgpoqBY/xKS8
QLVoMDXvxrxHz0tFXFbi/u/mV9HyIEVeFUmh2TfRNnxR2c/YYgFIqJtaGiNT0Azf
ETtE3XD6dF3Ycflnn7p7ZX5Dr8chLLxYQquJk/0/w6UKw2RYfmLI9gX9fBQyZCsj
5YR9n11FWS+I++ypOhanJWoiFAQYdWP3DGEf8A3+7IZr9fK5/Nj/kwNaexMpEtj5
o531HCJSc1p/ngpneTMwZN3B0cHcfJRw9gmdvYqShnw3MPTiK3kFsFwNGAHiZL3f
kkIgcNQS9EJUVEW6gZGIbtMSR3kREf8EcbtDe7ItfvpFtzungSuzCdGX6gelYCc1
WqHuPQpkEQ9RrkA+QrHlWMFUcAV6S4ePfxo0/RV0F4u7BS15ZXsQiQfg9gOSNFKy
z8TwKODXfSOlB3LngO3ymzfQLixfW1ddYYaTaGZ0lfDwOFcF8it6ESnE61wvOjwz
vFVe+uPi7k13CLrJeWh1pRg68v5qZ6MHN0cL8N+ZGp8IPiZgmb6tvF5EDIhk31WI
JTCZzZ4nKConpI9MvZkSs11H4+EWSJuggOX5yIMAzGgSG7yEBnOrxSEEbWEIvM45
BqyVfCj7KLop8vEFybnK23NN1X9+9VDhJig6giuJcVVcjeFx/O+MXZzn0+vxxk5N
bBeiEjio2DQD6KBdpVeVAhHQHlhndSw41ixJj3xKMg8TRTjCKzQP4UveH0Iw6IEb
mbm7fzOqiSqlD35mqK15BdKw3CxMCJo8dlzpEFahkcM8Yb8Gs1cS+3CtILdo5vxz
bMXxBW/Jk0OnUzjVnxGSNmkXqEuOC7cCia0cWn1h+Pszk9mG8ounimr8hUIgfinR
12oOWPscf4kWckE7dDoGSdHPHjH/Lr1WQvkr8sBxWSXCZ4eWY8JXob4yMfEkk5Lc
IQ57M1n9sgrSATMgf0MJxfVpDxeYko3Ek6eLRQ6EXoJxNgJV2Jk1yHhAXDSqx0N5
PoBwL6TJF5c1+SrhontnqMapfn7tIAbtb50M4lvLaSvegYsXxv3A48Ls4h06i3cL
SrTpX5/jdiJqK6MGo7wvy+UWer3o9mkfwQw4my2cHyT4fsph+4G4eOaWovhJLiPq
fGirReHZ7wSc2w02vjoKt6zeFl+2JcyV7fGbTx1+Gjg9DrBEhe4mBmmsODhemrMe
8PjmeSCKhbdqofOrTQnLv7+aD1NNh2SRalrXpNhUltmhSfQH+BXTGNlj/AuRjS8i
3Yt+8X98EB6VeAWzg42nrvOO9vPIJUux1+KSzLcDem28tTn+ASOk/lCrjx7MuZOx
98qAddMkKM2SUBL5wFyPsTrt3u6pRz2vvfGv9lPK9uWudu5oorVYOEsVYN5qnrnz
tqXdiwkgPGV9KeDFqK43/DUJhF1yqY43h/t4nwEVUKFccOWjNhadzhm+mwpCfbxT
8VbPSzB/Y7TlKTE3T72T9eePKmIyhtxOsMKdY4K3ZiwKrFHB9gkuvotNjO07/z51
JQ3rPYL+6q4MoJyNAYI2xKvqE5/LLAsE7f581u05cqlRx+CEfa9z52v0YzWNcwIN
4keREwHHM3hqOqXU+54h0y4wNe1rKqPUxwlBnhtdV0su7TFVLzH0DHQDx2nFHOeN
AlvX2op41SMyrobccYFAPnFMmUv5dKXNlwf7HK58W7qHEyIb/AvZMVQx3WigaHle
7vgPn66VtJ4dwZR9SaEEJg5wA6JhfqgT3z91u3Kb00DaQzpg2rsGv8yokJqGv1KI
s2NFezBPvga++yU6obbnE27y2tNh7eJSaxxCYn1VYIDC1eCjscpV4MGJ22ke5ld7
wOIqY/N8JYb5kf/Xbk52OvBX9hNJWST7bIZtkXwIjif6uofbkUjbOxrJsGn1nQVG
qU832zQGUiVwaIGv3sVv9CF4jMbtitsGlvjugYDdUK4k1A1hRwXoC76/psfhTovI
uux2fcxpbEc/oE3xVmYRTlGRMsy0LxpZ04ja/mg6gIukYAgU0yRywdW4VaXvekl+
gcqsFaRrVUtCfj8BJUxUGZgM5yaF+ujfOOEAyn8wupDIv4e3dXKZ662EZFay0rTi
/MelucUWMfmnOQX+NMiy/MK1ocd10SkwzJfMqQSto32P4GvxF6/YaWhiN/jumW7S
obq2DLusVGXUZG+tMi1hrXtsrRnc8ldSNPZ6i6GU1P64k4thWXUzpMBQHD2OURIm
pRTFYQ83qfxQJtCv/prm4BBtRHxHsCjXkbd9ByeJWMbA2LtDewZqKGsbVEF7vp+i
gMmE1bDjVoBxlWMmGVW3Y9VMoX7n03sxtShvBUXmMbEZONDi0h23/7Y80dcD0VBM
mjV6GYAZBPNQkL3tU+LkdhOWSPmv13PKdRTxhcJzZEUpo7NHPuYqsikOosZXsi/8
dZkgWY0FXGHa3QUAb/2ZJgy85q9vSqqs383HW9zPLC2QAf9GcleWkgzNN3XNjVsl
FzXv918X3N3n/INubPHMvo0WlX2uG1bjZFsK+5KpEXkaT1FjUa0Ns1gtpFAudjUA
ZEN8eZ/APLfVvG1zwRB9Ul74ivATaQHJozWb1naz9RbwnaX6ZUS5ozn0MBNeEwKr
GeO5v6D/MQ0Dl5gZcHVdtnUTGXwLqnGm0gZLS4Yys9KCz/lSzpbkWF2opEtIKphF
f66SVJ7UgfrsOoehguXbYyOTUugTnElVTh7v57V9LsfMobNtmazrjwGSnUfqc5jd
90p0gxcwOG6z9Odjib/nlgYoQWpUTXo6XDMMCgjcsb9ljDZ0Z5s8bbGEqwdM5Lwt
LGDt22u383voZAUQt9uvE7G7mQ9Xkmx0+n787UMYfyUb2UrwXhPaCvOm0WAkY/DL
onWJnbwPe3yRhJUlQfI3O10d2I4e1cFfmsd5PWyaObXHAOEpd/VNcKKFXleaFm5o
QZmMt3VDe+uew+M4qTcs3pjNOjblQ7rsYdyNpQ9AKk0V+IUhL42Dfj44EmJc7DPH
750GYNIYx6j1yJZH0xSpQHt5Iuyq59jJRgzPQ0xb/nWLEyDW8mxe9wXqhZmfu3QO
7W/6vIsPJMiI42APLPX4NP2/xlqtx4XZo21KMhhjcWHqcXewjI26/i48NB2qP9S7
vB4KWPk0V5uj1MQ0ekKHDkudj/JLhFTY/Nrbc0dXsb9MdD5VxCaVwnTKDDabRAHw
6IjubkCrYuZj5WZYdg7tka4r5O5dCiKnDlWjkKOHTF63EKT7p4NbifoWDAvpE57Z
SJu/qbGvQBkSrBxCmiT1qwMGblFCZe5BwFnzIwvrKs1/01A6YMknVKwzU2dcp3B7
jWKNwJG6fHE/Ic+DspTe0Rio7Oc24+LZtqUyeM3YN+gLhl8l+HShFWtL16eYx8MD
aarrAr9upeHd+y6e+ou/kyCLAqJFdaHPAuC7+tGzwTF3AIuu+3zzUhNwtjYX0yBP
To17EzOoFE67tC5VW+4Tzz1dUOZIU7tOrbBVTcGfOx89y8VqOF8NlRUZtDoicwX7
LrvuO0TpBD3GPQfsoGuMT9DcO4K9E4FS4Uq5ZO/7D93fG8VO/oR7fiWFhfeXAM/A
G5KYgEdroid0G7K2n+/jG4tMgLYAReBV2UfKd5lVH1sENirigDEIDEzLver95bF2
nX/ddjwoq+x6oyIEdGayzh7m+3sIQFxgLzt0IDgfLmjnRPPraMboQTwUDRozjOHF
NCJYiNZJ8npkKL+QLM9gkRh7uDVrdKnX8VHa49GEZRp2lfka8ly+3W81KS0gK8KA
HZdCQXDy4P8yYRQCxlUoi2GzQfWKhdOvm9vA2pvzh0qB/ESNP1iKb9U+/UxtxlNi
BJa06BFUV2/OL1rhbdGba4Y2gdugiC6BR9t1shTASjp1F0ZW9rHhIblzct06aQci
joBc4nphd3Of/Kasa/c/PUCRs83Pvoi8xNrl7aF9Y+DxIlwlZsgZN827dQ0v/V6j
CBijOYK9RYKf6el3HnjRwAwgK2aHZeZ3onobB3IqazbIzEEV//8KkqaNXQoQJaP2
PJZQiFhIppah5LJaOpdpFY3u+V1Tm5QPdK13r4VfsgD9vqIUXpqucWwUQmsearK7
LH635TjlksIvKUDldl4rQ3DZojVdou954NPOfza8sXCgWykBWhEAkgkIh0Vias49
Zkzi9ROwvnFKO2hv1o5y7pMvo8u14jcf7+OavsEzRtkpIAT5A51Z0IUoYVDAa3P0
QOxJGlczu7Oj0MGnybVtYIZSsppzRxReU53cVmgp+/f08pxRLYQWUbXZWcPKiI+M
RMl8qy9vjsvR5bl5ukdVlnIAIAQGtuUhAdD2yKf9HrLXekfsvuYa4QhLCSAtT1/t
J5iL1GcKC2oVUIdyMUrdxc3QestiraVMtIgVvgO0iaOknRCyHk9c201gVHrvLgGS
OnMIdP8CsIbsb+N/rnzk02uQQrYilGn6ijhE9bf4bBg0pMtDrAEvY3faDtBNz819
YG62Oljr38Q4OlZZ9mgWOLA3xE++qPDz+j6c1agd2fn9bAWUy/yF4jH0ymauo7Vo
zewhXKqKz/28qjbY5bLHE2garg59Huaws0VW5Vp/MQl0Rn+cvgnJgOUo3INasA/U
aqdxYY/9ad1bIIOyZDtgdkRKOV6COHnl36zztW5aUoK4W4Qy7tor/RsnHhPX8FiR
dnOfQB5+omv2aSzEtEKXQ2wSXDBcm6OqR0Ksn3T16PLtS6ArmN+EW9WmAzVfdqot
MDJAH2cr0ESpoL2rHmjzv8SISc8zvL9PDpyNJ3EoEpGuLkxVwsV+8Vb960wtnPBa
vEyHYPFw6Nsz7CUNb1yN/iM2LeNjhSpwx9K9/4bMeQDH9YHicqj+ZaG4Xzo8RwH3
Y2ES/lSN/itsvJ6k6hKEKhIJg22NwjFGj5IPRxGe/aF+tkEa2rOpzNDH+U+Sd55P
LLa2ZLr8bFK4/EVJAOIM/bXVTAN0uLrNiMjJBKmMQigfu4l9+YfvsIBEb/utqYCs
y/ZVrryl6p0IVIGKQVn+BoWyQZpJbVlMTUGFi1prQFfbl1SuB55jEs3VjEx/wnkB
G05pyCp+iQTAQPIL76J7qBp4HdwON9pExinK5xWiL76sZOB2+N0b9qZWwt0XaF8h
xiRXeJ8KBS68EXVgAfKt2iQXsiHKap5Z/VPa02fybaZWIPCwzo/x0hRGOGXt/BQL
Gbd8yhdDpR1dIz2DtR8mGGSULAM1+UiENch9yhlM5UwSpeL30AfPZcskIX81AG0T
Q4lLx6HwywQs1BcZfcmLIGqUDFNh/FJjEYvyBM0x8xz6jaxfxdO5BhY6uDItzY4k
7Yf+gaBjRLrmxAuz9Q6yY6GeEsTH4zDaiQvi8E5/42ESgGoapJWGE+99Y8mP0hmx
oxwDccUqP/j2ufgKXAlN9qRPGD/W9MJWBOI0LPIwNOYMNBt9uTdUNrcdgeSV2p9E
QOQyjboWGooPyvS9y2MIsooKgYdSJ1AIxaO4ZqAEwEiUMT4zJDbYlx5BxH0/C94z
ZT+Jkap50fjXp2rbmx21kXROS6vloDf66qBiON5edZXBGVipVQodmwIBmZPjRrnX
WHZil1pturh/yxFXW4O6Jc2Qc6JRep/m/VmQlJ3u2pTLMuP7/vuloIv6erjHUqTp
g5MNvXM4hpe7WWgMsQR6806gFV2InMU+WsEMm7TdeTtYtbXmZ5M2nnxj3wciD+XD
FS3VFlRFDf6gKJ60FE0CVdRSQxyX3/ufXKZnIG1sct/ivUXfnpVjhX/uFabGC5FA
mQhlC8zqZ34AW2aYSUBbc5l+W+DxQWvkjjYVMmTflP0HAIssmMf5UI8uNXsqAueS
JQhbi5nLHL3wsE8usUclzdZP0iimxpSRWFRx+3pHiXQShnKmXRjgWL3zvtRD/J1i
JPPwUursVaWzrkoAtbWbueGjwTz8bDEVtU8yRPs4AWhdeiNN4ciqv9r588FKs2F1
bhVTwaomMd4i3gLgRFgece/+fsOxYa/Q8nFPpOA9oIrzn4BcA3lxSXgn3td9DJBz
bzLBLPWoEe44rRkxk//TaCNhf3r5hf1HKNug8/SBx2SxZc2Szqq6G9hQiLtDUiYH
ZUdNl53s3pmNcdJaT0dHNboQuDD4pIpn5uR9n6CatYbdp+Srbukp6gdo4l/8sIY/
VXJVlknhR6QR1yYfHtD82cprrFnbwqojS2cP8up3ucwcMT0hhNW5c3qyFQwiiaXx
HzwrV+Xmp9Gq+DbYbHNyYDLNhGtRlrFFk3T4zr8wRnUPnfNYiuoITX3K2GZa9Yv6
klJKCpUSb3AYaxEHOm0aXSGjuswk5/tA5ElCV5BxaOTUyK1Kz/rLN3Izl8lslZIZ
UYAJx6KyvqOB6ufQ+LHcwMz8bF9mAf/Xb3qI2NLgaOkOjJChGnUKBNeR57o5ICpQ
OUrghdKnaAnIvdHB7/cTs8iEzDHjuSjPQ7CLG4zUB/yxn26TVY7VeAZiNfHPVPXd
hBcIDwN5/jeGPmVXufimSSdQtocU4jVFkWMO06J1lW0yO6rkqRGHs2lc86aeeFFY
DsTVvtniBuZYE2VI5gRadkKnLRiO7HsQRqH0Rkwh+9cd9K6fzrImlNg5StWeMD/z
FJko7RdOrOKSkSURoYHkS7ld3DV6PQvSvBrbEAVHBuHm+EayXKkONZGm2C112NhG
JuLTnxkooi9Tj7SajEwgWoZ99KspVzuBucoS3Mgq1udrUs/Mm8h0zJAsP5acbdGy
JZQXuijgqac/TQRiQ2foYAdG5rPwdDmxAIdMkrEt2cbTWsnr17AoTk4NSZ9EbGXd
io1i7G18Izu/Mdg8gLI84h5sJEy3ODcMWgciITOfDKOMjJsGOKESEb1S+XtWgP6K
sJhVmPHm+VKT/oaaiEBkxeHJ1yfoKf7i3EJ6iBQBkt6rWzwcBqJJMLPJUhvaTCbd
kwnt8zAjx/IM7sdsRXlU+pNqGikFHiGGIG04LjwcB5HV+2ur/cxlQdxGwr8Uf3IX
BGYvMzXyoqaj4O6P3lZETKnJ+e6qGbTl4871g/OcUOxmg5BZUY6rT3oDFUq1pSCB
rjRQEMmplqInXBwX+vX+gXm1f4t6p4nf2+CgyHD0UNIest7trecTss+tU8PFLgAX
EJdqvZhnQScWmcJFDV8q/fZHVr0mBuDa++TVM7f3CA6u/pjCv726z2AJvqqPHKoc
PViAjCS5WsX0yS1skX9KXvAweg731GoH2lKuR8Wav7HYJpWHJRSOe5XWWhzdbNUH
r4V0EtZ8s2G62TXG75x0kSNQ19LaTJF2i7pD8hIiz+MYpLA17WYc5IUwx0GViOWf
nuZp6U4t86S3GRvvrgv/U8xl6dL9C3aweg85fVcOibOBxrsdcWjjz61GZxhwNJnl
yFZ/Jo/ZfCIFF86zn98kvxmPjOdETY3oOCRRy2ZiKnMf5dXppXNpadtFAZzQyXM/
DHt0DPvkcOFmKAce7+YCaTMe3udlK6gzcvp+00o4ZwP/Fzu21Q4YGR+I/zwk/R+W
yg2L1Zxgm2ku23IpNllR7J8ha/cdAOoH1+Zj5zymZ9PzLZuCuNMgdc1hINPTvC6B
EeXqmLvcPKeGekGnL39FpjYEfOgncK7/i+rDNuWbspdf3LM6gfajJMR85wq7t+v9
C6uZm1Lu+PxRnGzdiQVIC9YxvPH1c5IczUxsve0KaDtSjiibshJHg1qVTrG6Aq9l
CZjvAje8pyPhcB1T32t8rag/39lnWfN/T4dElhmgMvYcuZxGVvq7jrwF6r3L7i5c
IkyjcMcidZ4QuSN1U+9qkyoeyfr6rg9FaGOynEH272wPr9nQMtvV8ZRGnQm6XBzE
Jxds2puvoKJgd1m+mSfPnknbnfv3JjzFQrrzsFLculusoPYDe+JFXboK816h7fge
V8L0J8WDMS8J5EolpMJkAnCBM/jfL+NqovEx0DqR+ryWRpTzWaY8qAiYIxUmiNul
doY2a9mcIHNYm22e3/Z/Dk5qAe48cFaMnnjmuiSs4W92SVFhaIqiaadLJwUfx85F
ZFMWPoFzx4GXZhDMae0BLgKb6AcH5MLdLQnSGebByIiT6Ei8g0X+eVUO1X8KsEm7
yiKV7yqxmaLgyUvxIm+GDHtAADIIrvSmW8AJOu+BucDdBsMOAbIQxqD6DZmOGEPk
9Ok5Uzs4WE5tpP373nphBLOt/VF3B3le6AVXuC0MXRu6SQDdcwrfE+bBgl1ei5UF
3ylXEs/1JWJFFpYG6zOXgfiPnOUuuXGEngSsu2+bBt/mmO1dyJYFwNmWqziNQDiC
YH4cSskU6M6qyCHpINhHEi8k+zd7B2LR7EhFlkSueXJsl7udEmfDrXgBvfd/F7bT
otu8/eqBhEkRdmuJHxMGd8c2ewr5HVfgss4dbg/y1Y5R7DMSTObBb3ft7Ke/s4NM
/yNo0MTevmvXmsSFLzYbK7crlPtLuA3XtlEZaJ/0CYik48EMm7nzGQh/M5A6BfaC
rY0KiBkKU8YKrpSe/t4/iUQXkE1mTjadf1zCSvEYWtKiU6v0oqCB1zHp5Nlh66yG
HU7VyHuKz1rLqFXhKJ8Y5EQsQtoQbgYr55ivRgEMgFeSy9Afu6U/S7TGqBn9e6Lj
S6i5ymvrIsTF9YnNoBZ9UsuBe9d1UsflXoES+DtdyH0MFG+ylGGeQzySTOZgtKq2
OY2Zq0iZSC9O9DjQP5Usy4Xdys5tOj+6J+dPcR0tMkuQAESmIjzzrdyw4DbGOGJK
G9khFpnE7OZkDZT5SX+yH8WY6ebt7K86jzlbrBqO3g40ASwNNHJqt2QDdVcb4/GQ
02m1k7OCehEOEz8jyjMoyeVwIKwyVC9s3FAGhlimde2BkZSv7RZ2Kcw2JliMnk/t
Db1RM+XYaattc9xEDl4Z9m5YbNy0R8gqKaNzZ8dIO6j3Tk/dbyDP0mTbbCWFIE/V
+27gsR2NAnpz12oD/7IfkVuCHh/CgzGtrgLel6TIRJYvPr0t/btfVcwkXSVXdR4m
nDUILurLDhZeHPqYVmPYZUG3mkSdT4qnFpo1CiVjCZ9mXEAe1y48J+gph8/OgY8v
JlXkbId23BIZZzGGa/yc5x5sYRQQK27xTmz4bAtX+3zLwm3nQarj+1CEupHtLVT4
0B7aWgPIE8DIbiE4k65zj96floIbn3imCqxBHf0+9VzHFctDke1HGFEaNRaYNlPS
Q/IW9MZ8znCj5Ksvz0UmMIOSyVCuiO654R3x3TwI2fZiCYYg3az/KTwo6FkqOojA
UnVO/NOogGk4cLteyeJdIL2esnwANlP0UNQHs8SKA/YlE8qUUvUvA/652hi6CS0n
wPmyLuqChZSCpDqriY4Mdb7MyKQfEPPQVsn1SVYBQTqrwicBeLT0D81TFdpnIKPn
STKcImJH6BNv7h4Tfrz+WWM+JuXG7CkQRjMDK+lL3VOWQCWUkhdLme3L6gN9Z44c
or6zcYr19+B5h1/H7BIz195z69Zy32gGscBZmqkcZeRFw00RoMtMZ2PnRZcLkipV
1sw8qVOeZGCk/TZAjRlnxsP+J+gctYkw9yDG6lZ6y6GlegjPGf79nAKcnyxSEuKA
vZLiq2ixuF6RLkFpwAMsXHR0ZByjq/ueFKXHQ8gbALlI1xu+6ejX8NDQavEreQAN
HSpnZnB+WowbZfYSDra+V0yxUKGwLF5B6k9pb5SrvMd3cCCCJEqEem1beBYzx4P6
/elT/WQx9I0ONCxps8/NbGWGgKL389SI2CSX95IhdG+jx/TxtuoV1Lt/KvMhkETc
Q3WyBH9EJnl7yRRqK0Kiqko/FbZKwe0bkUSvUcEqqTaWZe9oFwLUeIMjgeQ6WQc5
a4bxRekwKrxH+LjtqkdScSID4tmopysWwrifWnLKyi2Hfoo5OOSalNTW16OZYK29
zSR89EryeTqs/GpXWvmLI16vvf5GF+C7yKIAaXKWqmZNddunlwosXTh7ykvy6RPu
lKO8JJPv5nwBn2uv2uon45naEkyXlKnt8PXnE1m4ARDCwXZchQiYKYNOjrYH5zFf
QrQTlKRI3BB5URdoX4C1HClYXd37eUp7vX6msVydSK91+NTPGPdvz3YX1mUCUWcX
EfKq5JOIi7X2I7m8rlFBvq7HkQK7xR/SGjJB7Ssortl8TuToLGaxmgOGfU7EMVX8
lyfgHrtJ7/tCIjPN39EqIj/fvhK3G1jqg/D4A7b6y5ktum0EFIdXhPjOp/I8EWnM
5ctUFgJrZEFKagtqEhAty056uEUQCW0ds7VKWhZEOirIDPJgCtg3xngrdrexlYFR
KUbhYpZfwFBqwWB1x9JGZM0BfKsweCwSUcosDxyD0fE1ewLMo2fcg3EE02WZzCvk
q2a331CJYZXek4nwEN9jJXW1bbWRY/ZNPcmidUWyFHL6UmZBkMrSfaYgQlvHceGh
tWm1Dkb4D86hfV5KyEhLckWJhFV1GDu5l1w5POy+cqv3gJYPutEelaRBaeHarsO6
TMI7gT+uOqyaNfAhN+M2OvG9MBO4+i0KM2sIjZx7dJWJP4x15tRYfs6T1zWpGgkj
B+z1WQYQoCCCSBI6cRJV1ePdcXr+9WiUA/lX8lR5IYhNyOJgepzky93c//EWuOyl
ckCmMY0wIO2ha2UhiDumien22kOOZQbPXROZEnxXvBZMsViIx8EJCSZbp6KdPHhq
NjTmqQhiJnEjyEk86vzt2+Nu5KOHEXRpEbtTeX3dRxG5n5FdLBJBz5gKrsaTpZTu
2cFIRtI2lCHZjKg6O8H+p56vCvAF4jvjcWQ6t+qfuW7PZSeFoJG7/3cVxR5tibLx
jlB4i6JShdGQo2IXm1IG1PJ1veuGMITL8/z0sKqD/1mAfQb5gwMw+m3GN/LfjxuC
Gl6kjZu0YbIdzbkUflcKMXlSVX2NI3NnRUXIDewvN0xRXcod0/r70r5nNWtqTQ/a
+9s+rO/dPmtXqhu0CeGCGITwJFSlmjbQhHBLH42Y4yuPT4LtXAIiCOtMExV11M5R
8+3d1fYGCgJbfLl2y3/PGAoqxHf4Mfc2MNqkmOnVNKMenoM2uQqqdz4uK8MoZDhd
dyMkd8g7EP2opE/bjfaRlRlxlytpR3Ws25ChKvxCerYZV98pkTVP0fRMnErKva3j
lGMRvjCnHoMllipOOKgmpYRZVDuR8rjS7LNgZtsr1bHjgyfaub0fFEff64q8YTis
Ab0SQOWe3+GKxNDcykClNK+t/Q2XxYQTnHOJze4WnYDkT85rUZNN4y+VsHpaig5g
0pTBaT3f/AnbJqrXd7Uzv20ljDeEcrNIDTkByKvE4GhnAfuU6JAeQRg74vQ/gY+l
krNWdBPkISplF+umATCM1jCTmEkDH00vn6jwhafJ3VfvvCsav4icuH/Dj7sIp16C
Uc40pgQjHtIgc/rNPL5bVIardkZaILOyOwHj4McS4/dXoDimb0HsHydnvG77cKpa
e/REmbhMFSV4DUKaIyvofWHZeBBCk76WuQnt0VpuhxlupENElF/W9BoIchBxLoiw
UNSUHJXJ2FOf6FhyLGcrK+yaxeQaWoCseH0/oBptP3uwD3u/qee0lBSWxcf2sQbF
OQL0LUKT3opBzGCscSOf2PuBhN8SoKuaENGUzh/1U/xb5BcYonWwKRR10lPic06w
Fz0cSv0mrQ+NupO4OrRfreeX5vR8yPW8nuuv4hHA3I7V+HkSDTVtc3pQpnZvX3Zn
pq0DYIH9yXTVpc1BErT1Jx0J7iPjxpyvgce/cfdtV7WljwDC9lt+3uMEeEOBx9Yr
G4BysngD1L0YyflPVLkMDwlhCQ+tVa8e8cE5LG2rpRrw2X3jat90qpLUR/ivtBSl
D1wobAKnhwqFAiFXy64nOJlVKaF63tBGLoER+gXbVx4sW890qt6BhzZKpJK2YGsq
6GloTloUO2LpRlAKFWQPscuzDuIFpUCIqqoKy0j53mR2JmNGELD+PKL46ti1K8Ze
OFxBT7cyizJC6xEr3jGKcgKbUaDxFd2iMh+6oQJn9KhGBA1cyD9eqxu5ebq4Nndq
ZTaQD5xd2qWmBdcW9mkssiDawOyTzCb4ScQbnxPW57BWfiYl4RN44BpAGEaiZdx6
OD/J4oDKIob9Fdtjp2nGM1EsLOEj7CcPGIsd9ctRsDksiSCL7NxXbF6oX4K/wxgj
jH+/Urggz6l9fIK9r1SW4FMBi8PzKZT58uyYkes+ho9B6i8G7f5+yOstD9vV26u3
9un03oLmrqaa59+Mfc1A6qXXUgwAyJzuSKrfJiUm/JPTrgVNMUYojqyA48LHr6tD
G2EussNYKs6qrlNwC8Nrwxp2NAksH5wOea1XSAHSs7mnN435JTsZyGfzEGHtCJ8i
nmKZWz4Z2Lzs35RgiCgWJ7N5YvRqM2Nda+fTrYukmVoppxGoA/cMMCydiVzMK4zJ
j+AcUjX+l27v0mlSTxZkLpVcjR7R69nWCgaSQtd/upQ7LGBADpJZ3KThd64hx7fK
90rbb4RPyvfUKSyjiYGZ7PoQwHNN2Hyf2BcHucWH1+c9elGHMnmxkLrE/BxzxBHk
Dtm/g8g+L4q7V9Xt22XbGyOCpbvTMSLe9SZDz5PcknCMgu+D7ZeCqSnOxFCPSOVI
MChG7iZFCXcQZSuiIiJpZ3ir35kVaIBagDglEtxcTWawhibMREctQKqS8411RCRL
d8amyI1DQFwvJ3p1BRSzcXaRex5h4VB0YfyqHjXuIuyztHDcnKGFQyKzM/zD2MEF
YeFR8rgYry2SYVqqPqpeEj2HCTFGV5zVopmYhdKIJyu9n1gRt8XmFIxmdAOChn5Z
rWKgCYKfpTWQRTS4vVk55iCxmGC95jJyQXvQbLjHclSGMe4sQ1ts/o0iuzHbTfXa
1219NHjAwelQJfUZjbpLEUQdhI3UdSHzFWrE+fJ9SW6bxQs1WGqGdcLw8pmoshXx
lUtzc/cFGHUpamj57WcoAWvysgCvmiijUPinK+T3E8vG/VeWzXjzziWv+0Fnce4C
iBo3osVdw25eTnAmk7m1T1iMzQKjFDsoQMKTLjdiZeeFIgYxx1qrMGsHDPTFZmqG
Zlo9fe3zVSwcrAXtFbLL49IFSLj7RSzlhnXOfedckR65hnuhWkmGr2gUafZgbsCl
3mz44Ni+skJjWUL/FvnfOBH6GWm6L5KHyxFKft/FNtBTd84Q/OTNgeyIoIrmu0UE
JQAD1ttGX0izVmAKo6fkyjibbxrQ2yy9pBp9ceGwMRKWNWDlwCfj7qnO63/5HtgK
lY4Mw5MNQHhSDH0s6YjH7WdWDVOrq4Ip1B6HpJVjB6GkT5BHf4c3WwZG+tG9yGS0
KGtZO+PmfHHu8jr4CfAF1366tkofhBUEkxmvKDCUjqnixVLVlMC06YxhzQY9pYVH
3oCKGslL8IcEq+sEskGFjyqgr8GoEZFzCsIVYc9lKmXRPswtjaFzVu305Vu7u0uI
bVqbXK3+HfYJ7ZlsIdW6XTNZZvbwoKQJw2Wbz88xfWXB7rZrVY2SBGRNFOT4o9pm
70ZqnLPKYD1eM8vp+eCORooEmH+hl1XLSuXuoam58HGIopBKMe2iXrceactvTipa
NiwZ6CLA4XIoux2UXiqIP4gaSRxYJjCVzc1j9RcpoA+8f4FQ3FOXMk/LoopPndat
29zegG9+gm+5qekQkRq6iE3obJq3SGjSMfszEJthFHhxlDjWv/qkBb79C8GCWYhg
D/Zrt2Ba0379GKLupKnIDAwORVq2X3ADxWwmURoC9rx+yss9JprW39eylWRM9Drz
+QfyhbImU5zY2hMniltAjSnq/It53wIwcUMqpnv1drX6NLEi5ocm6CAvjxvyTljT
jTAM0Ha4E4VRLDGFu1uAXyPg1Ina/6/nODdbGXkjUacpRXiipd8G6yTkU+QvT6fA
G4xy7EsrDjeW/sIAzNtEBkSW2Fd41Xf4yseETTKnKk27E8MXyGxiK1bpsmiBSrpV
7Hn6fUgWPQjRYVH1awaVz2aARBGfxskB48ssaREQvEdelr/RJjbm2t/ch2awLOrm
Pmau+wpvBhajdnuI5je04O6zkhd2NCV2YQtgN3tM31wyfCFrBx0Dxxa/CNdoGQnV
5tjVsf296slrwTA1Xayh0vQVQNgKhJp9CQjxFaFhjf7n5Dq6X/uySudRZGB5NF6l
3NQpBq/D7cWTumOa4EuSZqw3rZLdu6c0BzJgeTTmKDQ5yzKhQqigiRtaZfU/64Zm
NaWDUAXV1rUm01tsCFAqUakeHuxsrpOCwdVX9PafwzlE0h3ICBc8jJWrYceySx2I
ZjP4MpEoNYI9s72ALlSPYjiv2UgxouZo9c5Lm78GnG5lOrksnWtvtFESzjOTc5zC
CJhCEazYI8lqQIIfFyRo4juWfCEUFPRrCqHlNAF/Dptiu2F7ecclvh8qgkUtAegL
ZMZ1urfb/gGyLbsfFug/E1+ga82oBq4sf5xNCxEucNLhr7iVF15G1TRlSuqez/gi
mwxoSBu6FlwZOOUfEYt+N9B8KVxfXx0FFw66zwj1nUymSG4b5EoCI5j/V0Ayhdn/
dM+xH3cy76OFOJo4UYa+Aww8FhaFJG1CA6fN8Dj+iK2lmO9TfTmuSa0RQgjjSuZQ
jaJAIH9Qdg0X+mmj8qJ0FzPktPth6njwy7PqruccLGjbvVn5VGHOsYGcsRUURven
9s6MB/G6lLySZtxUzs/I1fYUHayLi2+huolrWwt/lda+4DioHqFY7IhXFhIOkkpR
aFgpurXrdEhkn9hq/7nGbAN2bEWZ1W9ZTUr6fwSp2kXFXd4OFLQ0nZuCMoJk6zQC
erjttmdhZEp3e/bLEYwx7N5LcL4b43HdunCRRpmTc0MCaTNKqgIzhWnBJar8bSG9
QQLTLWvk6qfTnnQJ3Rxd9lgA7YV28kByFWFONanSKAT6s09OlBKiDOTH39J5PEbr
AWqjcrXK4jZGPntKFHm/uC0joqrkEkDU+ApoqLwf9GghW4RyQno48buzYof3vg0l
Vatb4Tcv89eQDXqHnxSRWw3VsqTZZF6Bnl9qDY306+dB4Jxj3YRhDcQyi9i2yMyV
dRTocbP2nft8+fkugLzlb8aN1bfL/ksWX6sL81+/HBqc7pehNCqNTetTuHGekTP0
d75dUfNGVsoQibcNZiKJYldd6Oq6O6b0k39uU4bwfewSMS8609bGk0Ro7UkpkmQs
lOGxbVBkTdo5vpSpWsxm6GqIkCGsi48xrjM3S9vajjKZNo8Nut91KwCykQVQanzX
3RE+KZ8RH0DvLb9VO4ptF8Ci5EtHu8Uz+h/yTqBjAzA1FE25urX9xceBfHDiPSG6
UJmGq9PiIwO0TXqcginES8SqyXddoEt14l/jn7eUuqhfGh08ij5/55f5l/N4G1G7
oAkNC1rBagQjGbVa/QRr5v4dkEtJwfEm3lYMmIBfWMN6+aq9tUk126pkLCCX375h
U5YN9mT9KkX4l70Vn1wITNtsaxm83kXljTQJRM9tbSlyfXV5WX2MKtbC4c6dgpql
6BCbnASam8iQgUSSOSGes5WvLM5tWTcBrUrFVzIR8Qqh7j174ppbqYnMWS8SSWoH
nruC/INrMDsmxmVQ4tujaGMFOdyvl5qA7FkMuW+foV7MMHWeofsJkXaavU/+dYw3
kAlDLi4mZyd9HkVt7IL4e4W1XFnCXU9ULGO6JusNt/IS8V6iTawpLL3skByE/HSh
Ptr+guUp2MFmOUSxWB/kJ+0jPj+Y54ZG3ywZPdjK5uu/PV7XNKxtfYEO+bqwigvh
yfawmRDY05pkQIQzSjvpt/GlxrdcbGwtW0I1bKPChE0EDoY8U6jYxJimDLw8rOOI
kWT9dee5wmyXyNG5NqSxIoppmfuwCNgXfSp+3xmHG9xfzT4SHw7F5m4GuckzGtom
OmldVXbTOSvCqtNbSC8bBlWMvIo2umCXCocPTkGw6bBukh3UGCYMJcV/3+rsjF0Y
2aEu7wVEPfXOT3QC9tp0U10ZfIuO1n3AtSLr07CZSxRGag/cfcmZpLCh/pZijVLp
IV4aneRHaEzLwgRXWUhNxzXSe6FhsnxrYi56ZuXARA3e2y9teaqO2Qi2aV+a+1Cj
mCflTHPydD873wme1uE8ex6jp9VF1nmwpbZG16U+dIv03pTfDXijKWrewTsczSZ3
OcI88ir+Ay+pdxzrL/n+kLkmGefnIZEroRqqZRELfhxNFwBesLuqrR4N6fvD4fTW
sqeewrqgJ4LSYfqguYjFqRFAOUngxYRd4J3l9WBnl1A4hwzx61qK71RqSEkCJ+CL
B0H12hvtZ2olb0Q1SVe73NGMv/Uad23lMCEEUyl/EkiuherA3xjhBSiSHYVuz2Gh
IQsqwCIvktIPGp0+G2MS2R7XwUge0CJ/iPAOqaKEzeU5g2geYsZd3MpmLry13Os4
0vpMRQrUHDkB94TaOniZnxXivubgzWHlACm2aPggL1+38gVnx11jCmjRTw4RhX8n
TcwfV73rWHcDmWUo2QcdiRDHMxIjUFBV3ERnQOF2mtcmcqd9WW+6DnZA4Ss8Ob4e
IqSOJJNNrkHSjXdmMyjX5bNrYVOLkyWOvAtkinNrK7rV088o3VhcLtm4aS8hC4/U
SlrnRmJBK3dtqFrJDtpxH7hexwNK0iKNbcPtbdpUja1odixFl1r/cx/lN8+7DCos
CxwRoU5GVs732wf0+8J0eefK/6Q3ZpsozmPsXCS34PvNMEUGKm4Hv5rNbSMi32Pa
805XbelognXk7jEcBAB43m9casu3P2q5hdetpwVZ7GiTJwHxzI/PdUfpgYWmQJhq
VlA7AVvXV0EUne4dNuFkKMmkPbmfiMXcbZ7Xb6b25TMZz9NFecgZKrohHNHSJCxr
cVkfG0TM5tC9X99jfl9lGWE6Q96w0N6CaBT/hpf3+0DFAXOBNPYc08gz9YQtRJCS
oP016gKKedxeQX3ElgGq6+Ou4mknb2VSKsiy0TqMVBsl418Uj/13AZ1AwaHxN3Pu
y1g5pu1A/1DgClGe361XE9wJ+6AmqN9+gHZu5Wx0VHCXNOQgEYAH8Ye3UcFSp0ug
K7FbxdSKMDsTUr7cibaNoGZ9HGw9X4m7FLMVfEP9JILGExVAmbCSh6kmpNXUwAxn
ralu6ka/po0FZHUm1ZjPsfSnLpPM+sNsk9jv/0zJCn18lzFOKkgteE2/jk8chtWu
S2ZUt+5F8kh47yQVaRJYP+GK/FgD1qd9swOpB7AoBfDj4Sltv9qmhTgyJX1zECht
3kP2hzOsRyPmvVY6rD5zRnIc574aIVhu2xNQXksMAHxpNEr+OjvAGMtMr7xAlpvW
LhXgyTA2gg24gS9eYtkHcsMyAUpztymM1heTCws4Jh22apfNHrdkVfbnqMqxpsFA
mlHyMWiEj7sdzPkMaUdqGFx1XDBcccOCP2a8AnwQ3kVq0gdmCFSpSTqpXTVOd9GS
VHwp4HXjYW6yQLacCwGfwlEuGcXjH0Ba1SephrBbwq6oMsbgQWeHuYqQ5cISNFSF
NAlfkfhSaIisT3f9RWPp79fN2fFQGzQ1Mu3jb6GvblL+DKjm0oFsF+qhjpTAxLaQ
S/UgnHjVffztTRY/ylLAzF02G6HbTm4YYbf7V7V8tdY2eBH0wegs988GdP3t0T/7
zoqsCsBqXL2irH2dOGLNFnPgSP03vmoyTxVgBeAP7xPwlQqr99um41APhjkoM8I+
WPHcA/GYEOkOpv9/14jJjttJOsZAnwULUsD//BNSwuAZv6GO7wtIoLoztvranYnZ
HNHxTkoH5EzdkT3y/o2+MVi3p2SPIybqq2TEfRW5nwmt+ALJqo6VB6UlW/j3zyK3
1Edq5EWRfTphoNb5M0mauc13jOkFR8CC47Xs7/ff1Oh9/tSvkbK0zj+0eqBKFENe
aSxxOQg6+Z96yxi1AWc6m60Bm+tOhH+vyx5EExAfE1ozFMvxxeDWV6RU7q9og2K7
NW5ACUecUeEl9ryTWZQ/A4QEyZ+87GpFLxeAHmstsMSyEnBrflUPI3A8Bs6dCgwC
gmQW6V7MJ6Fzw3GpuWXnkE873RU/1MvzxrJ1CSeMn11jjZe+gl6zmDbjJc9XC45f
zHdNw1zET5+CXBiCKQHhFC/UPpNJxUg9zgfJY83wFupTvVS/abxZzcZaDyQJUskp
ve/BlAOKfy8gq+m2pytjqkZl78eFBX9qk1s3c/Ig4G0gQvSrS+mMVZFWIgNlyl3T
5cSw5OH8yiM7xcv5Agelzyk+BaHgKb+gmA/rfhqdy60ETTPWM3HYBAjVGCWxhnfl
r/aHDm0RNUowrrQDpTyTdgxAO1ez5lKcOGNjb89MvQimFwazkq9KuCipvVjYgSK4
xkNCsBfEaHK7QUaOnMSlfmhmcIANsxYHdfc3SdYkza+LR3TuNQwyuESfnX1i+zvg
NmPbci28Xj+svkUr1OQg2nNyjos4brOciCO7xUiqgavwt/3ZudldIZZ8YyPqZvd1
sgUm6H+DDap7HomAqhW/owqnZRNs5fo+ZYg/Hm+vxuP3IjZvl8mw5ZZdiwYAtzrQ
O0EzbuWteIbODp2aNP4LBC1Rmx2vpLr4n/5BCNNJ3iaC6a+zy32yn7okocgmXg/f
9kvgXAUk1TASgyZ3u2uqLorem6NnZ4apMrJvjsc+C3zuBQW2/Z1FMN3gzP5aQvoP
ZNMLvaeYU4DfYah+zBdomIXxF6vQRr4PJSLz9uDc/zcCgNc2/2htbA4VdqYnYLjD
OXS1EKVFfolokwpb9dZz9u6r1xMPO+Dx9Xv71TgITxWmD1DMTbLVX2YSSTtgjM07
QSvrKuWXaiA0ySLMH10QI3XDbcDXBLB9Fc7zCp4EGH4CfXo6j9ewKbaCitUOVTV1
+JGOGcfzmSDHnyjltPj/bGTlDJ/iXfZlE1dtB7kgsJu7/tXMR/1sehxQT0+vXd5A
38ukxlS0YaEurlb+Y7NZZ2+eDgNMUcr5BtlJZxOlYyOQDt6etWPMeCXyPznpCZjf
XemA8qW6qwY6//WbIvB7l3ThiCac1CO8OnaUd8HAaNo/qCb4FgSFqJtTlkJto613
VBSHDCS3VtJkAxtjvPUlaa4bIRHGNG4ZyYpo2wK5XHY9b1ZgpNDEtBBYw1GDU2Mh
JDI0g4ynZQCLz0j1AmTOKgrSjvsMEYwRNQ7pxXdtlKJ83GXgeQV4KbsHAPVQg0UW
adnWQUOnqwOVFnGCzJpmv9JDgdPzLwDumvHCy/YmTdaSrExPvJvk5fddE6j6C+XP
+1o+fiKTYGYYpazqC9LZeRqYHtw0yTdSq74E6eF/QR+x/Z5G7MuhnUDO1JaIB1m+
LOOBBLl+NkBl7zfrTRW84C4jAcU3w1ItCAdl6deWeLuYaedlCDE04r5+/Bk61uZ6
4WA+bEOhfI3/1raZaFZNV+kiFa1AAGf0mG8EWpeBui9NEdbnF9XWfwy5xCMER3FF
BirTkpflGyo5JNGnidmPpVvv5GGFRFIIK/kl++B9Wdo419ZLuD1sd/ZqVM310BhI
2DMNRl6nBz39N4ojDJ48zMrSZsQ8H18dow2vWpKuJhneh9OcXhETtlxF6+wVweji
sVmV51MtGbiw1+A4wSAd9jhx45FknU2SfswLceBVaT1v0vD3r4+9g0AoFpHKxQ0x
sdVMhT4wAvgo7qaU+As4UVgxo49LYYQfYDb4Oj/Ocp4lbipQNmFlFJ1JyqN4UPL9
z428HKffrAMuDoC6OSMsecNjm8Q57se5FiZn0lDI7kHD18/9rZOsZqO7ItiFvwEq
eucG7sBiI+ENdsgz1z1aG54KtChVkPP4bFabtzBuUaBWHTT4IB1v5rEJRSdBwAzl
dpz1Z9VemIUVjNOnxFRl5jFlJXQ7HPW+AvrsB7ko26wjfQlXBj2J17rhdix8Dth9
2nSjy1MCpmQRDsTtZSJmJxkSpJ1zs0mAmrXI/Ff9a8whEVRYJe+aiRq28I9x1mLc
4zw7EgOeijL2waBYKzUx4AVlWbTiQkpxxbYGA9wVJ2kzHCWOGNTxUeLvXUXJZZw8
ZPo2Bw4/2yuX2RB04o9bwiqWMNp1uaNetkCSZLVhfigF07hg0QhIIKXzcZVi/NJF
+qGVUBxqcPTaAjwcGerLByhwTeWR6TrXv6uxcwfMpLt9abCcGvQsH8o96fPe9cvJ
VRXHdiN/jlW6QU6aqC3s9V8WfWo/KHFTrgTX3IdBg9MBtHbsP+cUGWaqJOzv+hay
ryH4q8vEEf8oWsZSakH4V6L2+vJ/EARA90wYzfpyVihoyxiFoybNvSHG/Ktgr7nH
NZN97AvIbmo9T7lPVjKtXBf9LXpzHjIdjmoNCbbJNzJ7X1oQPtasqH5NG40t6QhZ
EpepD9XyzxLuV6vZ3H6yrem92Kz2x0DFz0BzXwycG7ZW/Ne84YcxzIla0HqOg1PG
y950Hp1Zo49s4iAl1KZxXG4R8VYVUeEDcB3JMRgEj54Lnd3CkWv1irSrgP5TYRas
GrLD6zQc94SMDstfEznzdLDOb9xjoOLBygo8G1MPaK3onIUobR1A9aRA5pRfOuZW
+ia0mgg1Mtt85VfyusSxXn/nYe1zSE7UG57ix7VLGkPQLzQm3k7F8GNyemicbAL2
3iBbKNu1lqo/xti1gSV6tqhLYCV+j0bKB6zKJkRxf6LPHsZJgan6vmKrB1825Xhl
Vcr83QVrTK95foQFqZbM/zjX4oytEnxmEg+eAGl3imHbN/5uW6PcqH/q4lbvismc
//SFHON0oPKbpab/P40U9qslVVYxvnkhvQhZVcZnH04su5Il78VUzAEeg7zmM5Fw
CCY4t9X4+fjTKnQUOVnForE95EAX2HO9BJeMoQi6FYeUun+uH8mrdDEws9d4b4Lm
4Gz64B6kLByVUciNcMioQZYqviSOaeaYqvGvFgdk2byLJlIxbzppiGsD4i6fo3Jo
BV37uW/0KsXg9Jo0jNZfrNrMAx5d9Hjul7Y/7HNAas//nzD2sAj5v4XtFI5wc5u9
8sR/H3CxQGL6thsRtjoaMzP6WJN9KoY15SDAMmNwyQXRw1mlSY/zax4U3m9muBbT
ALF/xlG0kY4dF/o26kff8aKY7BxaxbDnmC6rwnZvz+uxpdLeDVkyButlwg1Uh1b4
DY6wa7bApox+B3dmjerKodN462m15lrNreEkMtGxPUqYIyKEiIsT72CtH/INsVMd
soszhN7aZ3yfhHoyvFRbMzSreQSr1yZcytUcJ+sFcbNcOXlFos+C9AEHYoA/btxA
F1OHdF3lj3e+k6bIdZYZzzouTnu6ZVLpHOEhrpDS1Js1jvO8Znvh1mMJkoxiELXo
zkvwNdEwLGK93qyvwm/yeAqXauQtmRh7XPfAoKj2RxaeVSZ3YkJbhyA7Kp/f6Aw6
jvkkJiAow8lqDCXqgDw3Nbgnz4KfohUXi/RiTwqEc6mNkQGB1RWxpuknUs877kdt
9D/+CKYR/IQFWkNW9IRR4zynFvUhGV1rS1iFiebHkIplc06rRB8cv8fNJ8U08Fyj
d8+iW7oCzVjmOKy5w1Wn+jVwHGzH0gypt2kJ6IEd9RQbGK48octvV6vfN/T6wTQx
jo/0rjrohPqrTRW4JtFHmjnFHxxRN9wlwl6t1ZUObzJaBB4gnztqrUHPMWjyjdcW
YRksoSm8Yo5/g/I41CBTv9Q6LgEA3kXQfguh42w7gY9MFh03PXvElIEHwfRK43Wp
XCKjaScnnM6q4xSR4/4qfO9KqZuc3wUKLosnv7sipbyfPDOG0b0NiQ48LY9RRC0z
YOC3nTWAz46Lc0ti3JmDTCQmx0bOwRUU8L5gy7QfQbW7Jlgv9B4p4aL4eWurzHeY
1qUQftLg34cDF0Ke9uy1Eab9syycKxhedFeoxS/vT62XAut4vBpIdT03pEeexBk+
I+6EMwY+Fk7t6Ta8rV0XlKM0Qqim9Z8h/vcIhzv6O/Qh784rmLaL1xSG4KqC2Sr5
xIG3nr7KlYJLzIme2HfqBfcjtwQARaotiPDA4socfZQQYlAHYhq+bdowGyeQKRt8
alnc8PYQArWrQHyqTyYjokiGsa267HOhSgurOTdN+fp65xVZz3bQRzKZKdAcMOW9
CbUsqY4GD+ESjlGvC73pECK+sObidT/wQklXfYcqCWO6VZW99z3WPu+UlqhuPoGN
fALrVEOuMPheoICJlvPXvU50eko04thbjeRTDxHQcjzpwExe8uj3pWYzZ/rKKTrv
N0UlzrEwQ1GVpTs0S8RvZODibbXPYGtjzOvwPb++hVNRIt/7Zn9p1P7LO2XTiP5i
RbidV38q0t1/szlgSlnsOG0eTG740BjoCNMbzJXZiYHGv5kuYhw+edF4mscDkxDr
AVqkR828qTGsHjX49WEeyYnUaE6D/o2ujmX7O4Vx6piwspUZ89C5080AtH0b3GhO
ec5XOL+zyDpY/AeSU7oezbNiftyZYfHGDxvH5kiu/oT063OqOkx/IGFcqTZEd7PW
lgKjZHlrobTFTnXr8n1LJhPe5mX/PkZsAu0Kln+3Le8o+qTANoSARRYNzQJjgVNi
dgwZMGutUBGtR7yME9ytIHT1lDCuOccBwKPu6WUxpdrK7fLBcNYyEZzT9hQpfUbM
QIF2EwPFyMtMrS7Qwdt64QdvhDRfR7qVSjNFM84F/EdIxuEDptQCV0KLZoI3NBoq
vcYbnRLdUGtlAPK3i2ClP2ohNgHwGajEtP4rDJKDZsLoPciRKc1euAqN8RqcksDO
96LJfNCLq6C0vemvsP8OQnhgQbfMBioPRPNyy/8fzPZVe2n7oGOBu+WFFVTW0Adp
wcQIo3rgkBj2SH+kx3owwWmIfYUc3t/eqlo3H+4HkhbAsMtXCQuVgv7Jni2q8OIc
U2vMUTWO4PsP86mD4F3kQmf6DL3P6/yKUeicFzodCGMTaObgmbu2z9u1mLuGokWb
ijI86wHWMHWIQFz5j1eP4uxd2Nt8nLdLztVhA6mYMla9Y1iw7k3OuSl+yWO1L7bU
RYkW1wby5gwUy/gjwwBM2G9zgqz7MADDewuxPG2lin1oTcwuI5ql1mIMG9zeCz4L
7HJDn2ZmyT9SeLrr936PKV7PYhtFDsgBjnhS2SRHG31aHFBPXbmKlcRKCuKH+ecl
BN2w7H/N7KvSZfWcAQBZAwnIcJQmHFe+LGYz0cnQdoByPC2p9E94HhIrOu2GrVDA
3L476lPYL9bo2iloqBrVls3RcA6Hkv+THRXZQ7fmUXKAirpnqi6MvXm+yecKAXIG
Eti1qo7Y23pGY+aFJkG3oMifk9wcwr2i2l/H0/jzbUwaqlZ20y1FVBPMbA189sL2
zQIUqUeCANM47r3WrqvrWXiDGEAiSyeTE5SpiRR+NiXEX9OOQ3exuhjv1rnvvUJL
t1B76NkcsEwf7ykrlDqSmf9HBqRWYxcqPgB3wF32sLlTY+oHHbA92cECIJ1WFx5U
SW1npXj2lU7fbMTqfSm/viYBX1th3jCUhM9WTyaQwBV/KWaosgPqOFlpTGaazZ60
ICOgtXkffZ8DFrVeARaRpatEMOpafM2m97Sgq0+N+Xdr2AtPReLjzOiWhlZ0gDuC
tjRIcCVojhblNlNaN/ElfTCXANOzJiiOMy+KQTIHd9wFQVr1JBRAlF6nEUbP0to5
HT3UUdAriBxjPT+9lCXkHN/WRfJ5pt8XgHoOrHqHper9fMC/uL4fk5YFYzRgN1wV
1oO+rJQLZRXLWyFxuMdghWNdMeTxRD4LSuk4eJTNkGA7rNrar9YImj8atwfx6cME
RiwnmXq+/1H9hcBefHIZbHhF10EYMI4QWNYvOsZHZH4ZYU8YrWfpmyJyGbyoKF7m
YQSOtE130GxSdKNA1hHWMK8OMK8R1Yzd/TurFKzjltbtAX0K0KU6sPioAduFtyUz
uYns5uDwFzAsOa4yj94AvppRBEILjApyk8MGHep4GuAhaYmNSbnPBG3Ty0jnvf15
cpDdkU2TQNiWgKfhImJI2pSN9U28FlBHBlXv1Yo/ryw0a6lr2JKXuU7om+DmM5nG
xOJwyZ7BCWAWcFyWjV3qCzXufJ7Y+HucdRZzNtViQMMMpmj/IgYfeFDtOjt03XS/
LvLSmtCd3qFRVlSGtGJ3jAfn96vcailwP/bJiWRr7TX5cNPFwHHajV/ObpDdhZfL
FLfRS5rkZHQ34yCL6KFb6GdbvYWiy0mw3tZ2jpnqgMjh7nZOWvg8aFCf18qkhUQP
7l6q7kxGq4afn84v3skQQGQuSHIvVb/t4Klm95vXQ5pFJFe+B3iPnJp9OQWSlRT0
u9l/JTjTY3EzCwwBOI7BcmtJr/JmN3cg22lsqll5hSBiiQ5hcbilzzpkk1OybKu2
Dn1Y7WM01gm48afi8el1MsupZ6AC/6+AQ7soUtTTuNPCILCkLQuHPBWGPWuN7tZt
upbsqrMegbrW4vsZTtzXhX/PFGSAMysft1peRqzbEYmVmldeRTdl9kW8AVDzmjgt
DljEatFJ6yEdYpBRwP8oXmJWO71wNJDE1X2CMmnNGzMgIv1m7o4VYSjJ4mLFoK2l
NRe4rCObVJs50WRJ/cSIu+RNSLP1d7dnzopkGE0al6a8rhSPhnFfRsttDXfTOJPM
Vwk/46hhD1cz2Xxs+NIUirFrLqpWh20FY8i3nWldX+zz2dg8FB2kfXOODQfQTEHs
cgBMiDU1+DjwX0nfeMUGyNwJygT84miCLnT13FDLQD8D1/es0BLflZQ0ueM3Em3t
pZm3zwOj/nHDdwvJMmbojNyJFMIDJzkzE1I6SPibrl1J4NKNOWxqkCHwjkUEjv7F
ebyyDBqYIABBYb+q/gPB09JGglQnnVNwyPCGAL/BxcZ197lOTzf4XSeKyWieMerX
yp2P4EsmxE0cw35HgHT4c91EGelZaaNlnJ1KU+W3IPORGDTRE4Zu6/bdZHVB55PB
i1Nz7is5u7jRo69qZVg61Q3T+W8mHhdInM3k0Lqan1IdHUBy61TO7rP47eA5Waa2
fyjtJvH98Kdna9Hx9d5+vQVE9h5MtHQzW/qVs1yArOzDIjWwGFUZzU7bJKFxKWQD
G/RX4hzKdIHymku8j6wwG72E/rFRcBCYM95WyW3LHLK3MsYmWMRpN7Ym6mpN94dD
VJB2SFDwoQ7DbM76KfFUk2PrmYCPrpODz3aOZvGULYB2Bb/qxh4+f78YpMoxYoY8
nABt3qD3mr88FXLM+bqhfFT+mF/sj1QKKXY+O+zDf5Rr4ilnQSsIcAtNhTHGLlud
Pqf6KMfXAItXqyBtq6+vS+NgS/MqPlBkbOMfnHTmeOw14jLTYJVcFiLXbObe1riD
Pvq2hUpWFayPjdvZQUdlvVvEhnCPSuVLAPlyj8NqNQqGkbiBh4Yn0KBGZ/L3AX3b
Uw6zRztOJtIshgtxpF63+JwKsDhIB5mqk/0D2hlGswMAmU29i3suBCtxcd4GH6KE
2qC6o7/VmsFm73vKpvOZ/TRkG6FZaT69iZZNfrHqx6lFX+YsjG1MtQ8TzpoPTKG8
5+Pu8AweYo54FVDBRuT21oBox+cCIt0YQLAZPicyvPMr0EIS0F4YLdKpyyvJzn4I
D3EauN0hjrjm+4/0PHcvgmxoS3+PIyskbBHdIuYZfwBXiXgmpwTXwhGssfKS+kvr
P1iDeyY22qvOLO6YVYQe95VqLNStTw31QuDPHbG4p0vamzqlti/+O6Nh7/rJN0b+
wXumb4pvTcWgp63ch9Ky3k4TFdURyZE0scmuvr7eQZWMOLBeUpVoASNc0E1nQcEu
smRgG+TVwDEdGYZJ+Rt9W3vpWxiwa/i2j9WJ+1x3HWCPmRDJnMIiCR66VCTYRvw8
MrOTLIV/VOySBD5ZweCLU4PoRMsTtLwMObOHTWRNBDFTCxJT6aRuIrzge0g94aud
WFJKWxqsn9QuGECRbm+CpqkXeh4wGy+COe+NdGZHpVZSJ+KQMVPc4mEWfgprIcMQ
FEaQ/++BkLyWy/vXBhWmXWPmxYQoGMnu4LiKxv8+vB7WjPhYn0rj+cFD2DA804mT
cWgmuJ31H3vyOd2hZjqkO6VOq2mtvLpi9gaWgDT1mF48vi+sG3Jhgy2oxPqEKCuq
blk3XIVWuuy09UkIMV97exi8wkemoy+T6HSgJSKUGKJAtxhDgDGIAD7BDU4MkxV1
GSOpdS8br37qlkQjMJJYldsegewANsYMpuEjewb5UFAvcGjv9UEaSHwYdjK7471S
t7nH8jijIzvi5luyNc8c+JGM7sOYTJ6Cd1mtEPRIsoazw4spY0/5idHs+9dsMZ56
v3i0AlD7IaBbg0hNscEM6hZ3ZzcWfzi57k9YBDYz9+Y+kuZxZItA9E/4de3Jz0X5
UEeZTljIjoQwwDDWLAwh6XnjSix1TvR926OTp9AFIUqsAVc3zJNJdw+BpnF1LyBC
LGrnCRVyU9bGix/t27SGjGzzZqbXZdr/1n91etypk2QsPNsiLUskwol2tczmgo6G
9hAdyDp1c/MhwARnDll80yCDpi5L9dSNja8nByBDqH6hgogk1HIClJRdstvLphkx
3YsWqDM7UanfnG4t/+tZiuu+6SIYsP8m1I/tRxwAWmKZUeWGF5Et9yowfN20IT+Q
Jz1vw1tNSBFih7URkRUYZOH1PGIFFr1efRXoruJAUnibBs+7UvkqDfrCYJ1hzJJC
2mUDgP5HlDJ+NnZxplXn9s/uvmaJlf/zKmzf8BeRkCb9aYwLxpNm4gv6lXwHuuRV
vcPlAKYGM1aORwK6aKjqHQH6yeq0xUm9293eFoqON6xHQb0znhdnpC75Vf8xTkEa
FYn/E8bD9ZgrBcZsMY14jL1pcZb10jAD7WHArWnLN4b4TEvOEaj8Znnv0wR6wEHD
oOoFf8uwIJ2BGcO9XXZfXX/7f59mWiUNabfcwMaHpa/F3vymCZezs+eGM2YCsYOx
0Eoc6aqdosnf4ca4S1veXn6H5cJCn9YOXSkjLPW2AvcMNKkVdgmieEpraEwULjnC
Cw1Z+9XtYmgTEBYWStKxrx/+QvnQkWklTB6JTjnGi4RfsegUbwY1ejDt9r1vVCHA
bA4GLrwq/V0Iulu4h2YftrgSIRcg0t6YIAZNmcECHQopZzmoWX+/O70s92IiKk1N
G4mpdoSQzNXZW6Ed16yMMygFIHFNDDvvg5UsUjdaib4V0Yqs0ufffuFDWN0xBdVZ
R1MdTCN8WIi1w7BQOyuRHBrWPixdkVLRUpZGE8r9fH55RxmchfOFxrDGYLmoY7hc
LIAWN1h+Gsb0r5bbOgFvlhp8oZYWpRN9+RPEQBCsm9o+PbVpHe7iPeulun+UDokL
IDS/MckroJ3CHYnkdi2kAQSCb/nBPOOpUpYeaPA4GDLGoE0+erAgJIKuzEKaKAPN
ifNSJZzoqzxhOCpFDsCFDYsUzHx1zUWWVFswVZYLs3LtWTmweu1hs/K7CHXl1rCy
YnbKGHeh12TPXfcPKkUFqIgqU5ZRPbMPopH9Af7f4KTXNjDl8sDs5/p+JUbJzcMG
Ot8Uqp++fqvyO0IM7jzUtlxUPazDnG0fyPnzNT5YkETLTRIQLT8zWYP2Vr3oC0c4
jm/45duUN7VdZUCfZdD8KVdIq/u9DPeHrZtjklODWxtTNa8b0GJuDHvKLWxbXfSp
AqbW63Y5+EYCVknaqpAapswwN2y/I7HbmOI4+nDXfN15Pu3vW3/RTv6u0IjeURXS
Wmvt6pZd7YFowMu/JHVA44sXm79pQuhSDZ4P1PBKfWNFufhii2RgFfaNlOP/eV7T
PlSzbmWg+Poy8+Dxc4p8Ibew8X1tH90WgPCVGh4a34WlkHD5i6A+Epr8k7W1mghG
t5ol5aHrJlK56ZjLgCPyY+EVI1awLEg+adzw29q4WsGXzhpBDyRC1Omea/KWxeWS
iEamw427OgTxyLS3i2UtcVJQlI2DQkp4n5+xWPb5O9pEFB2vHBxIlb1xE1pB9+V7
5SS2GANPRasW5xdhtJt/JWifHBvglDmElwqJlidtSbtslJhlJZ4Kj4qdy/HGhcB9
mj/+W3/+aCg+8XBJJGqoxTLD5Tk6y3+IHaALbqTYVNm6a+6RXiTI19F0QvOzoYIt
W2SY2VuibH2V0+A0AwcOkmbv8cRvbcTHIbCLpcQYkjqCyon6F1Sa1LuiK+4K0AB3
tjQM2rOY+JpV9Mlll0OFVlP0X3wjA/3Tcdrj6cLIXPpwDHnFWCVFcjD3Z9JkNLTv
eh6KU+R21DWb6VFAm0UwR26vUgaY5xxEhbaxNLOEwJr3uSI9F6VTWnlwku6XfNME
cPecKqYr+4cNAqTTluWcx3Z6Peloe7wTG2lKz8LChLCSt7qyGD9SC0iaipEqI7Mx
/aM9y1WL0mcHNeu5kVs5A1Pvh0t7K29hM9fq5AlzFZU/XZ7xgTwD0xE9/4KFaH+O
+VyUA5XcXTvU1ktRiVnxx9iKHyRi3YFzTNzUiqGREHakfI8RIYC5T3V2uF19pERc
Ie7IWk+gh6d8uw6So5vL/Yg6blAOojTcAkIZFGtaDD4tS+n0Sv7Se/2ENN6Iimy4
16YCwVtgkE3EJrXsf4mghoLCmCEr4F4y2b41l9z6SVz6yBHiR7Q/2yAijmYup5uF
pdSrE0e1KLsrEo8kFccQl4RxzwD8bX91JLjMrxZ4UlOWRsZY6X6hi2Y0zMhkXXDt
+YaRfTQVG+QMoCxWa4Yjp6S2CMfRIYpYcldMozVUQDe+wfQuWN1XQsHdZozCqRCL
lpdMib3MTs+Zd7voWp72YnKDH0OjXjylsLWK/ToOUi3lWwIxD9gkVezL69uq9bhc
g5Qs0URKuOFXKiumVTOO1C+wFdQJdC8YAiriGU13ttnhbYKLF6o3h8afsvq+4mZw
SQqPcSDnD737vC6ClsvRudqxRZa5V0d9glpQxXfaAWOk4jmpQZV1+yB0/uicYvix
5hR4SFaGd3AieG23BPyucNNlYBQkfmdEuZA3nsaJ6PWAP2LZEz4LOK0rul69rFDD
VWIrUF1o0pnBadPxjJCQJXaHLM1/I0HMe6h0S7ZlVY1A2gXcW1IfHe1ZWnXG1kBD
w/kl8YbU3iguv7nNmrFZKz0pevoThiQyJM+cdJGY7cwXEMdvb7ehrbGak3WI43+e
QZTAZrlazxLEkGKkPg20inqS36lqHVlk4IJOif1jC9oOA7Dmg8EYWnE0U0nzUunl
C8H9giJCFE7zmRzMLvnPEbFgRkMM311qgBze3rLCpwcSY7X0SjCTrRk2ltDb+07R
xZJadCtZkaC87xCiMje6N7W7xVu35c50EyKJOQBRaJRr5MN0VU21m/mRv6deUgmH
VnDLrf38WzNDKwP42tf3fS/FNVPVmYK9AM2jAcwuaWhN5hpYUe7irvDXhAhltm59
sXsg/vfnS1w17at1xONKBXpoCylJMD+WRBB2N2zBSmtnhMKh55CY37YMEfdr5y1x
LS6lloYnrk2IDBZJ0aFeN0vwuU0dV2g6AzhdzJfgIh83jjmt/dLZuhbeLk/lVO6R
PSKFlOCw/rwnBlDpn6ZCDEd2aROkHmwLiGHMS4YyOew96CaonK9n3ZlcsXeCkM1u
qFKc8Y5oc2Kb3+8M+MVYpzzDImD2+tR0KDtw4Id4DYASBYdv23qrD0aQPnGvS3ma
lP0SB3oLclZDUbJ1TTpm1uQrb5xT/I8Y6mIlq2FBxyEqX9qg8ZFnyCTk9PHvLX3o
hsTVyBazrexb9AfVDQnE3GDe99z3N/fq/6Ct4t2enY0qsDmX3t3Ip/URMPdhAM2k
yAMDcErt7s0XBz8NujShbua0zM/18azLe9TMBWiIMLsgNWgn0piMa1GMZ46SIcYp
1H4UhrPRv3fDVEE6sxC/j7p/fvp2kx7YFukuS7JMeLxjiQCm06jG8/G6BiyVEESH
CSyimaIs3SYLkU2pGdgBAueSyUqZvzSSuACobr1xTg1BJxTGzFeJzwIu79WFIBjV
VNk+Lr6vbXrazloZvg2U1LM/Fv+O2tIf8A0QUrNnjjhvbwDZfY2OZ4hNspY7qqO2
LdTurCI25+RM702XNFkDF3GHZpRyaqeKAtJhjaUH/VvfJXhJjlKnzsz1yS/gUWlV
baMIRP+TV58ML1jQhTb+V6RKcW+YY2LSI4HU9MbOxodsqa50wrLo2ytQ9dyp2qE1
ykfe5Bg37wBhGsy1OEeEO7eWYiTvnRWaL2O/WVWQPmHktGLIcH4TKO3SDqgEPAte
2yrgoY3PcR6g9KECP1NZfqqq6aNzUn6bpOE6G0HGcaXCNFsNyUxZwv/PU+oYJVRX
W8DgziyUZQ4Y2FdPZBdcgPK9N+uPEDREw+cxP+kdnJkxTgSAYMcB0XEReBy+sLGS
Vb0Tlpe5LRWazMSnE22fZ543hzzWNyw/TJUd2nOIPA17l/aGvzQwmeXOLo/m1EZ0
CKBJ8OhWzN3K7JdItT/BBebLghseinmCBJ7hzltfIN1CbBeqzVpHoW5pZsMCzYYG
4Ax4RLYnUwg8e/bXq7mFSlNk2rLghy6H3EOMIzLy4rNjEk5nCSkdzzO6MHrau6hv
uuBEr4joaZAxoowKwTvGTe4JAJtYs4daqNHoTXGc3UWR2MppVFJ4q9fKallBGU9C
qWUDrX2/GGlzt461HG31kr46GVJo+bjivEel7jhFBVgq01Fvtm8gV8OvYb36srnO
NMZOcUjbOY0BuGH8YzTnbMEXiZCmgZVosEvd87x5qs5BNVaZjOBn3m8sv7vuIfeY
HyZSstFEMiWCZHyAELl4iMsaGdmATNcBJTSODVuvRboZT1Y8lF5fT6qYT4oQ2C9i
IDsxvHSkZskHt8zTonaHUCUeNgPe/AeQKg5Nq1dSz9w2OmZjbJXzPW6Z1Et6fexj
V3F8onr0s3Mncv03CZ+aU22or0iy5e3lrIE/gG1OyFzkV7NmqRNEuFmVMwBV820o
ciGjuU1C3FQQ23oApOArpOcX3oBfh53GyHiCDIU9nVflMUmJzv/sXCNI/VxIPf16
XQPsgIfI7zv/2e83P9xsyt4dYyxk/2IeKFXsT4kaBii+rnewYVYfe7fGnGaqwaaM
16msptMTQd4JSa8oL5KSUjBpmOY6gA/oBtohw995DUKTARRgwAu02KocKMfh9yBn
WKXOXwVgT3TGLItcWIR7Eb3iSM3PYB+RRQaYJIT29frrwXmrLNvlsSXulaWJ4MHv
O1D36bgvVtGyIgASGGCG3mKd12WhaXBxw0H7kmsi03cxE5KaDPkyoXsXUTzYChnR
mHPGi+Eo7SmNHNrUt5B8Kw3JlVnZZogIhsjmM6VEJu4+RwQkRxW0IOC1zq18+Mlf
SG9zl0hZrDPiKwrtogJolsMCzO6uDQ0EiF7n5jofsZcGjPwBWF9S6kc9ba2FNoNU
UZATqk4H/SIbLOkrx1PepSlheoX1ozQeJHlmFS26kM6R0G2KmKKdiUvrAZHyy3ir
1Aqgh0f67mZ4ITQcduY+au2SvS0rgST3S41EgicFURCBtXQo6JoLloHen1UcJM4C
hDWDhjASdIBQrJw5dVeBmCKiCK5/OCWKpLZqiOTpWDCginf3AExSrORSCw3IleVK
oBkvB2c29QZFrDBjucoyZQm0+vauBVLo0iYw8ro6v8T2nB/c96FddK1PZ567eu4r
xU0UyJQumDqJBFyax2DvZeOxVIYn76b4qKQS38P2+jlpQzwhPibdCv9bw7bjE9Me
4DXfiIyJAp99HcHlNF/jQyh6K/Th6t4i+bGCQ5mnFiMbkI1q6XILzonXbka2OA7o
MPi5qBhb/cF6z90w3oRzHg1XXdgMlq7tA1EAQBu0V92LaY+LWFwSGN4ZLqtz50tN
s6WeawR5fPHleFQ+vxfdDYy00L2kvegI9lvXD85T/6cwBggVkXTyXCjKEiUUIyul
N+smQaW7+guec1qmHrRqT1z7Q46ECkLGmGA6gZMK74rnLPgfYj3A6R7OGPHNPTEv
BSzPW5/zbfIYDpdzzkKURieZVF+aw13NsRs9Sjl9HsQgJXV85tzy0Jtr0dEBbW8Z
xwtITdJo4ZVRDk8JIbkklkBb/Q3x/E4QwywCw8r7njLJwvWNFlRv56Zv51cyToE9
vWUyxewkdtsmCxzaxU3SKpyZ6HqxVQJu3NaeWDmMVznyoiJQ3uiz65mTE2JfhwJb
MEpk/F2/x4k6FoDFAEFhibQPlbkFeGLuh+KedrjexBD1rWe5obAtUqxr9TgNDXXG
zpoRitvDLMZIMrASRTUpx9iY1f13vgaTxgcQXgP7/do34BGtuzSWKF5SA0YnGVyr
q6+yHcvVyHB83VpunhptDzA+y/IeajTEwH3t+7OXWt1nxt5lAALmoGncpOyOaj2H
7Hh41hOYQmxm4m0d998wQndNkJjkuYsxALaSx2fzJIrdyKhh26pO2EvNIk+t5Q56
fbqKM9cWD4vlOjVUjrj/8e27x01QHUylpUpkmRxgx4e/R45Vv0+eN1wm0XR8xGiK
B7aC+MtswqoQzXaEe7MZRtJ+CnBmP2ViD0ySRQTCodXgjmRV5OunupoXABwcwnzy
Z4yl37BXT8ilBTiAoHceuVQt7JC5SQV4TPQKjZDVgfTD9ItRrYukdUoVAm/UFN+f
FjzhxMdjjtMSGLRAarTjMthnMW4VItqpLWHQRi9+Q2yXYZ0On6wUkE7ffBI7S2/6
VYEbOczhgidHbsRuTFAZEojrZWCE4FmUG/AWRM9ATSB9J9ixGk9EZHU6vHoaKPls
jAWaWaLFlvCmgg1flw7XYL6Y6Qe8gglK/y6MYE9Tnjp9bV/aTCIj4om2P3pALEdh
9BUFjljYFH2RvEbU6L89YYC94jfMUJE66tmGcKLr1lfNXfncGJ7GPsj2Q3rnS1CE
eshWLBypAQPOYzW1EzD0GgXHmbzCio0vkw1q5wQv+92s0C5u6F2SYH4Avg2fV26a
T31Enf8J3b02P0aCzwukGvPh/4WYSutkblA+RA+RWqUjxC3H7vrM6tiQ9OJlGti/
3MsrZ3vxDKkd9xjz6C0Br5pyHEYhGBUrhnZLIvj1luX+aqPsRPfOLE8EtbTRpB3c
XoOYfzug20ot281o9vQjI/1dgBPOW1CxeNV8M/4tezw7nakkNZUZIM0TbsJ7/FAu
I5LRcIlkpqAxwekerza0BVYyLrLRy0SMQKrKKZJekbLKQwjgSIczThbRW2li/E/W
YXI7D7cjmMBvkZr2/VOlat5LGXe8CIvfSFs46DgnlAtpn7nkHKItRY2D8jRxYCg8
vzTJXXjJ3RP4NkFPLjM1baU3HJC2lsbx4AxyA36q24LSEyVJFxcVbnkiLPxck6U5
sSZ0ugJj3xj8NKQf3jAhnpINvxV5cPF6MFqqnjKYQH0mmKxOthL4SPV5phNkVQy1
v2Luu/y+mTvOP9nIvDggKRigEGaHoKMJIesNy28tHqXID5AJuiay8G+WZcAOD2Wt
ZlOmTtGRH+hrdMbh8pbW9eSK6gmVLHywGdchJTkdq+6WFi7qftRNAHq8hKPVxcPA
j5dQwFlIMO7xneM11Yewa7CLmQKotWD+KGe4XF8hkzEpaYuugP97I9S0cd+ixpUP
Y+YABu2LOcg/vhaWRiujVBfNCVZyrtohRmQVzsMG0R2bmy/Fw3l4rZG+ve6p6/Z3
QP5H3hNnylcEO9uq9/KxOG26oxrsrJKsFRVAik5nE3oxxo7UdKw2/HpnxjgG4suS
/ZEKAgCdeHj+kaJjSS2NZ/uSoEdqKJ6mVb3Mzg41A1tOKKL0LOhxJJfgit1hYec9
mES4GlvBMZ1wh68IRcRCWM7L04FKCReSDowqboo9nkG86gn+fWizFbTuTbAmNmDL
Uvz5344oDXK7FGLzIlAwiY1vSJL0LvGviIhaVf6zKCZScaNF2k+8kFvDUhcYfAef
iGhfZvbVOLnp2m9ywdgISpkemWMv2RxWliVfHE0/7QerQYBJAHX34KI0wfKS4teg
bR+0Fq53V00Qb/XvaM4y0nGmE2Ul1YA1TCQQJVug2exSQMdkqDVSAVQgHkTdMty7
hUM4BWdSi9Boq2tUdj1TEJfiOP669Fq5N5yMBv95mboAY9iOPbF8kZgNIHD09TW8
EdJLief4xRJEcLD4kiq7e2tH38Qm9LduelHR5khC4/mSbO9u4ZrzRs+0/CqKQBAK
8mnbfYuGJLhKVWhFti0m+bbaXhCu12LTI2WnNMu1IkzXMwtV1MF0Lc5+JEJzsmVQ
j2a/ngMzzBRKe2y/9rOpnIeXMc3m3Hd2E0lapCoBBxcTTP+QAJgDa7KwAYjwq0r3
jU7BnFflgamzeVG8EM1EIwkbVfvWhJzCAIERxGttvJB19eifqz1NcW69cSzd+tdc
ra8D6xRw0UF1aeApCONcEKyKNnJXWX3OucAW5lozoR+VLM4+7/IRyKFbH2W651Rt
dZph67o2VkMJeUJ0d1v3rCoRVtODnf66MefqHJD2MdPaWoWO0bTO5ZjLS+JTIUqS
hCwZ92o/QJJ3GRzjtW6ptLSsTzbNGDhi/012YV6eeL3tFHRyRwU6yCR6vXvjaBkX
g3Y8RBMmxlbU19yPLdyWDEJQoOzsx40cy5ncT6xDENBOJT0jvBXcmCtSLy1oVvCH
cXSrculYYqV54XBrj6F03PrJ2DaHOEQgIoE8F8ORfbbYVR35fyZa7cwTE8DrOXyf
ZlqcMZCCgjOn89W1O7Y53eOaC37HjNt7fh+EsqKMEEFZ7Eg1KFSoVPDMcTnZ3ReI
6Q1IussSpYtmDGxJyM2bOlNDHjk1giqQ3b/TCFdk0s1+a+0r7+2lbu9N0lPaqF9x
H3UuoMaU1lCE4TKIw8OoRXePr1FoWLqlHGDioGxBtXZy3nomk5inMCAn76H3OtIv
OgdJjEdOnQA0cndkRm43sarKXXpZ5hs76+Zc7EaVzKbGjZK2H6P0gL12mB09uc+M
BDzyeIoF0hP6rE7bjG+VYM+Xq6QKeamH5e88YEJLxgcoUAcYSKedI694W/e65v3N
RFkSeBjSl+o36AvRiNqxkP/qD9VxJFWHIy6/IxnlciMf95v+mwICIKQOlrn/W9le
lXJ99WimWZ2TuGZya4TAMJ5k4NyJU5qS3BNfiIkaEb4nH2QItlGaS7xrVtH9pUgo
a8W2WOAQy/vLabAhxHKUyQ6+t74ryqKX1z9FsrFZ8jDzCmYAbfhkRzbiVs1NMloY
n24sO+a+nW7c0EPcQWJir6dOzGlepTvego/JgVO4w4EAAFJGuh30lh+tc5Mk83y6
cfHW4AhFZaS5NXH8DMMoIjxUa87RsHoyQeRRpuahE3eMv09Dbvk33iJkDAlKsxym
uGQQbQKH1GKC4bFnwH9+LdtmNs78/9Hkl1eLfziZnNryM9U969QBguQcX6rD1hwl
OCEjGCuOT69VxdEGhLnGX2nVw4V9iyg5U+JI2SpSjmhoQ74Yh6BdLrkTGY0Glsxk
WWoxdwzjVOi1oZiZ5umvBfHmcNH4h6m+scHkbpamFAVXV1ZBVpNkcUMZObAINzX1
mjqNQUT84B3tPrA9b3JD2HNZidDJIIhgJLmViL9CCSu9HKNpnKaEJRiLXlOcaOPB
nBEW4tKZjRMRMTZFxrOoZifN83G0+xM+XlVQjqDUCtlxeOaRzmhcKDaoq5RvhXM2
kHaFnPKJgip70gnP2L8Ckyy35Czorss3wqZ0sRZuKgWhLCF8HJZxvgIlpGRH6RUT
g5eb93/vusARwAqAkRNGWK7gMLbT3NIJYmUviC0eobR+y00Xz26NeHfxLdOvY9BF
XnueaDzMgYCvpa11k9zj54taJm8t16bMfQrPyhKHP0RzrsDyVSp0SrGrtDoiS3uT
vPQ/sP/QJWWJzZmTSYdCpkQPKM4FoQbnCRuzzRjPE3iJlbahcfEpdBa95NL/UA+Z
fq5TGnYXfqdLyYyQ9WX43QW0lWx1RrLMzEdECjZUkNy9gtUdm8CTZCXJv2ewf/Sk
WfZyghpZAVjKJuPY2h7nmAnPGT6kl+35nZfEGD2vhF4wT1wyRSllBZ2IrxTlqa34
uncZSy/XxFxzrAaVZR9kQl8lKVkGwbpXw+8c/SdKg2dwsteAJmwaSU/w2LT0B/ir
G/xaCb0auy1aaqtN1vwcz1s2n6JP+W9BTxtklUaAWD21bluinMT2s6a9+maDcI4f
KkVMxHyuCUs66Uc4Xa4e74FzB5xKRvtVpg061JYPCGbCFhPb15XqjtxwtrRnthjT
tnMncc5q5Sond2L4NP5t75OF2Nad9bJ2jZ1woKdOdxWFXE6MGQbNIE/jHYZANV2p
fZAjSSdnIHh57/A8VcOr8ABxd2mDqtQqYCFaDU8pJGgJCMBIzKNs1MjnDYPWaYYh
Yin1p2P8OnEby/Vh1HeF8zTnAKUZGsgzUv4zuJxqunGB2GkKRrA0CUMvTULC3dvh
5/og52OgHbuY5559L5g+o0CCYJoNgs80JdSFFT/p+EkIwnt98idmBYG5bloNIhzq
TtpQYbwvCNY9YYnYIYuLWY8+GTrVMSaEQenfeQ1+5qKg5lDhy/t2EHMZmcLLGSNN
2PvmpbBfKzyu51nZUZiJz03+2bkyJNkx4DgQvHyJL9o+No69qXYzp7Q7ksXeZ2je
CBVbHtovAYGo26WnRdn5KFA2xuZhN+A+f5E9BM2KMhCpkgEkoyzCeK1YK+3d8Qp6
ZG83YRMYTfc8sQIYEHjB+eiLfcZ+LC4srOQ/gV8tokdHX92DIQC2hNBqAySWn6lT
zyc6C7J2Q9U+9PdYlxATrQnYnswVTXZOIvwhiT+KwgNkDo/K9SPrYoBckzlL8vxB
LsiiD5Gp9u9KSwQqcKoJpZDMkw0NHtOmqieUVUydHcRE6Ij3fHtmrgIUbWsiBDX4
FKPIgOlniz6uExiMAFzBYKuK/TtG1cy9wrs5jy2c45N+SJ/dN/4F4QCaaSb4ZuIi
tDeHMFL2sLwo6KZrkKC91kknVh8Fnat4+n3YXEUk8/4R85XvEuVlM8poWiryNB8l
HRfnUs8TW+h6YU70sRtctHPoWiFRDGXuW8Vzj75BqrCeeI9aIbmpMDxwXGiXLh7a
exZEwr+YfxOBnZYz/PqDOwwg+wL5kea8UypbfK4ThOmvzGML1ttXgv2O2i72lEGn
U/kADMqzNmznSMKl3fSIhb/R3/cAztth0SRwcKmFwu6id+x1XK6fBD7e5UPVRFUC
IyNMxGDT3tcprV2JomF+0ULeuPXf6fczb/t0958YHY6qM43HnGiM/Nz5/kgJr1kh
VS+9JBGPIxHqu+HheP4dyldIlrGIXl7vwofOv9OpDDqSOC2PLCzWU5R1OgnBNxQi
/gNdJk22fN2ReOdjwekF1FDET8Drlrd2D5ZTl0HK5YpAnxvWywlqHGBHyJPg7hv4
FI4IkLcO0qk05t/kEN+IFEwIdqN2lAITqQfN7q+u4M/J4Z0TdyxEORsjb0aNbUuN
zP0Hh0OdTadohDC0b5DmxNkrEheVQhn4cHKL7l7m383S9stEqpZbUGybMWJLcezH
bfMdzqINbt9edIs52O+DZ3pZXnGHbINMwptV50mpMUrxLLex9QLAgRw05Gg5XezY
cQqjRarfyJ3KpeDh8Nyzi4mnpKSxOvTokYZ8kz2Iis8FujeYRF6xY9aL8EeZ6zrE
j7B6j7U+TOSMs01f/FCvdONEUlLDRKat/zuUVaryNw2K2nJ6sGnP/LWbpp5HpV9q
X2Jcfnpn4YzrnfX6i/goiiPHy1YK8vnhCTDbbsZ3SwnqPUAgUWvhhsxJq3xREt4F
D/txzma2RoKX4khlVYn0zHVo7FwCVbF0HCDHwcbLuFpYw7huEI/BFsvCChBWChUy
3lZItjnhugAAqgW/HNNUYbQig1VOov/tyIo6nC9n6bvMHzyh1JkhZI2YT5UnjfTG
LZ/HTnHAkxYvfFpSBk2G3wmB/YzYs5vj3dwgG9+qaK6JZbolwb8X1kLg0NwTFJJW
iZtBmX/lc6SCY0LxMXlrK8wUf+gsj8ZVtrylgeolgCuR7eujal7L5RM7HlEjN5AM
oRHCA/NN0+1JOoZbbht5HTwrTlGF1bSoNCrvaddROwkiMzA7t4+aOW4iyVlIZZs9
BcnnOiBiU8fDSC9tCJqDDi0/ZddU9eteDoYQdW9jDqMtTAiOdxhgGYvXrmUNkQm4
n6mm/1F1WeQHsoJu9a09XDrZY4ZK2N+OYHbvD9wS9+iNdgGBzvgMDTfKz8EeYP34
3fZNwIj5pgwWsaTe1nACfkKecuFeUZxjsJ3eUvEth2UUb/jauemjBD560Px8G1kn
KWlTVmCbO8oohXeFQWXhLWAWeFQZHRjHpDuh1WLiuYF+23Cpl9v6MQCaeBI1a4GS
39D6glsC7KKQhtOslOpJVdIWBZ/u3UBmISASaRM2OugGR0VwfJrphLkMSzjzrkkd
0xubazdpKYcWKL5wP7Ce6W8Vo7LVYWVX+L6vNNSFaCorn9giwF7V3ELPGhdXDCbG
sosYhpFPjmCE5lLaOFj8FMt/eOWDKqbI9VTMLUGxIVbK0SeNmReVIhfA7U8Ah89a
GdD3b+WpA/sv28L+vfcOsEuCneLUhgRNdDmp26X8scffT0YmmtoogYIzyS8jJ1OB
oLiTK/kaviLYvCX9qBtWRj0S0pSQ/BypEbwCxHlYAXTAyFgSW4GDgOv8NjV2nry7
75Xn4AiQ2HFNHABNJlfjq4P5KnLYGxK3SGK3DtkZcf4j69Rm1Si7aUrnLoyDxHH2
qSjaHwpJ4g81qMoyWaGtVn2cBV/Lepidhr88gE7VjvYSs67SLUIhcREKWMgRils3
Jkx3zapGJ2rm1h0JBUstlqC62xvcRtKxuWNxiKob1PklXcJOXiGrVuiXEi4thGW8
kBHlRDmm2qtpxnpWAmHBN+wXwYoesIwmLgLvCHT3IBiqC0TkeK8V8RBf1Fz6Hskg
8L+eF+yv/CRLKPuRM9zz28i/Lj0KttAMsHhjsP/0fN5/sdH1mvtiEbJM9mL5TEn8
egYjEZW6eWOEIqrroHxxiSiYm31EWZdDUl1U69tG1bat1qVwpPWp8NcE4wWBIKsK
BWYWDdFzsQJcAXp6qJVfBdESoTagGxYOE+7+E/B65vMTBgY24EkosniE9KVGQjkM
Vd6Nfel2epYCQ2ylkl5z9trbIEXQc0HDlyDXumwH1AP4NzXVSj/L+Hc32q5ZpJzz
DOCSsXzNq8gEpfj/EjEZ6+73lfcdWgRm1heGim0HQa/GA4wQEWuVW8TFm2egBp1y
xuXniPam6NqEngLKAber0XEoJdy10D62JUfuh46tWYzJkkaHW3NfDy3U7HicAunt
jbllww4uKOdafp9sBaMU9KSBSPmpvHjttYKB84R2c+6zCdVXPjwDEcArdsUNbW9D
FAGuYVkx0EFep5yEKPYVF0I2Zqjwrz7o7f5e4OcIykqpU6HHKCc4USjMdUe68tuU
9Bze/OX8jk5JtzFRA9mdk6d9HWEGTtDbQupq6lGgnuCnHVRowvrIBkiKTyP2ZVcp
ojiVWxleAloAiaLUx0u3jR6miid+mTk82UE7VZToRwoz2IqFryL+zlWSyqB7MC6a
DhtWYlDLkaMmNuik7rVquAuZ0Sgl0bECu1x2KQb0AbbnqXfZkKwGvEzWPcULNRmA
x7IzcgpsiXjUORI6k+ziM4Jv7XRORWUdr+Dd7ZC/O/O6iDOMluhzKHtLH72X8vtH
mm7gKGHtI5syQGlFfEaaBJashHs+6+3A8bhkWB2EK2R1bNmWh09kOahKWz7PM+Fw
FfpQGPX4mnO5TXdO2s9ZHEjGEK34d94l9leM2SWpFCrM5kG62qPgOtbe1OgQy4yP
lgw68zcNQmspdHkqDaJqcWBHxUsmaLfC0fC9a/zQelFFLJqTw5tVDgXlI8QoTiaV
8Fmdp+5j9LGwi93ehF3cor5n6n2qhn6VFAeHOqlxX9dopT4pWd8kgewB86kulbPK
/g2vrIY71S1fy1WlrOREPoZbTjQLrtXVNSZ5JrJduFgOcWkUsJg8P1Ob6JTgA+32
2y5dvxZHxF4Ycks8UHOC4wEw6tlOcQAJh4arcwQjh5P/nPXIe50FsiFDmYBibKwX
0bUAVYueCnZ2Fu11z1WXgfiH7/7NVbW1BBf1iH3vx5ygw4frZhsmU5JFkfkGyV5+
Je3A9qDdS2QMETxqIeTThu8M8M4stoEngwT5eh9cgACd9vERUbkuicpRMSXP2fWw
hDeihN38jfHM4VgxF0oZhVO+DVaQvAjdCqGP+c81yTqsjY3MvBlBwcWVoWpuwn0B
beuJSe4l/XYzdOHyg4Pue+VcDNjhXLH2hCNvMIhDRJ+zzASdQBLJoTNQN3E8Yr1x
FStVHFIJ7BsXrUcVjCCGKmpiYPk4tkyIDYNwY2A802qucBrFKctyLyHNozuC+GLV
YR0plOQlGPrBL+SCbVZTS8eEYv8ygUFDqQUT++WQuDs4kbHME283szy/E4EWtSVT
9TZr2aCojjE0F+KoCSY8ucUBVaxrT0Ecm0rcVyjCq8kUITxA1mf32oqpS5cOXlSV
4k8/P4BFoLqfqByCZoEaJog+9mIH0SC90tcl3goDpmjiga2VPB3jkATABfKgrt2r
eCrNHM5hVpAYkZcRx7usSkRrNCDlJbAPcHDQo6L4AsPzYKyqFkzNFjb8ra3oMfMh
9/yUuyFt+3nwWCNACH6SSoksQkvDMrl1qT6qgb0q6RrXUw3dAFYR+FJ6FtDvT29Y
7jSw6vUX4FsI1iGldxGApPEjc/woDOswDHflOQcKb9oRAX1U2vYduoLhat5D+O0U
z7knStxho0AeDLVv7elBmrUNmb261HWasUKyrMx7JjZf9QfK22oPAkAXqxJHB/cF
x37Uj4SK6KsYYpqsQP4r4Z/qgM1qgvIlTcNn29rhEvLSrQU9f9Z8BJySxSPKWeVj
B1EvGeGwVL9youASYB4Bs+LsAfkVnWP2tikfJA5/sdoQTiTLVFbNK0+gvs521olp
pQIZCCemGBROWsHFtO1C2vuAyAVM/9xSDvh1itZsFpCO1AIY9woNv4mwjL7nVZ8u
c0PyP+yyddtuLjyM3A2y3kFeUCO2seFksF1HTIyDl1YOv9z1wETKn63JqXjxmYun
uQBLZ7z6HnP5X+2gtf0W5zKLTFETWIalOyA1oLFUOM+GidoyopNPnhvipwENkEQf
THYNFNWCHE8QLif7cvQon7NjPU6FOMdpwT0Q10XwRlD6mBIRiXUhNShpgySuqUWP
PXwPBFXdyaGQ5GkMognd6Edvr0Eq789vsRlkETPiE0VZuhwf80+V4UZOriMb5Dl0
bHIOwAnMXxF2zBbMMxTKlQXv2fxDQVfQmBjqEddLA+rLa6boV25BDWbrI6e9037a
Hh/ApLHEvmmf8RzAO1vpby1SuGHfDADPP4qte5SZL9H6ImUd1+R50El4esav9K4p
o9/aAinl7va9ScUcXOf1ohpHxMIXlmggpE0vyoK2anSp/swber5pjrT1Qb/bx1v/
S0I/4ZxbdSLzSPsK1KFBWXrfQgXVFkJrc7S56HTL+YG+znG7+3euQ4MH7gxBgwCB
O6d8dJoY7NMFu9QSsK4gN3Jn5FDEAVN7Fy4r2Mcj/jdE1ucfLwTKb2LVpMx27Buc
ZEb+dlsep+KcuFcP+7nGQZw/dHkBOegZ+earWmC8rEmfzVtxVwWQ6ARV3waMb70o
BQY8J/wrRfWiFd05ywdWajNw3us9D9dy4Siw+kbPw57NPIUhUV8guK1OeQRF+WFd
HsgMt1cMc09b6t6h8GQESV1JenqoihNkf7GQuRQQFbmjoGQSXFl5urv/ly7AK4i6
LqJ6Zk451leUu1vbHgHJ+AflS/gV46xzlMSg2XuJHU/bdbsOHrd3+YrJzwziIzP0
cac2gckGBXERldE2+afcxTkqVjswN0/r+wF5YSv8EkV7j7Vsiws0IgeMqe2ivYyD
b8Z9FggtCc4/zzkkw2X5yUbzpu5UgtRasqgA3iw6pZtUCx2dXqGs3YmibC/G3kT5
nlzFil0LIYnmoXsIwtoMNnT+3DX0HgjkckF1ILIP6OmWgvPE9BDE6PgYUUpaN5ZS
35MSowcGo1MWvI/2hYwW6+/AM3YjejMg2LWQPPxmB2YPgBZ5+jLL92a5fFssdSka
tM4Bg0mTMT9OBziqjF+dyC4yDDJv8kcHAeTSCmSYI7lmA0CyhobuWfmf+rT1ZYXw
6agejlhoDCj4WLcV5wnDL/4Kx7R2gTMglDxjPl+PCkW/zEnyH+urWZfgT8ifzJgP
7OIo5U/GvL6N+67pPk2lk2cEfIG0c90wX1L/ySzmEtEncKOQc7wpj/DTJFnzvxqp
si5qtFMqoYg4KrXmNYMaG4gaKzYEnQMKzZE12npKwShQVqIgjN7XpCeoJ6TbgOcE
tCa4Vki+XcFK9r/VtfXM6VCtCOu5D86B516Dj2mCPVaXJCLnWA5MQRQyfe9opLEV
kOyG5p436aZgoe1K/IljyNAON0QMCGRDkVtdTzmlFX0vGIHasPizpKFPWD/UwPFE
OXwcusXFQUUNuaG3+CDDjaiRhQjkmNeY5gPkfgo3kVlUHZ9tooAvWMRLqi3/i/Ux
pL/byQOCYv0k4BzDEyw1x1SqLGUCvwnQhRq+w//GOLV2U9VxKJT5J6j4gn+l/C7s
3Hg09vVIy6nkcY33obTd6ZpEpCg9V6motJSr5ClF32N5MAU+69T9t+VXDW3cnbjK
nMxSPaLCzZ3oAyFgvdwr/0k0XHRXyNdweG6q9c3/QmZaYpaly4bQnC/Kk3HkVXEz
v83it8Ay5uYw+qyTAOxUMjx+zKuO8CSnoQQRoa0T966rcTdFz+rgX2qFRTiSqCN9
aTzvujCEuZ1wIxFNEatsdN2D6S+fBtAwC5PsgplTouSzC06D0sGYPpn0+qoFYOP0
FtGQh+Ruog65oTzwdwSWPreheQyFliPkdVjaNMGp9OEnmNJN3k2O7q+W0w/PpDPn
x5q7bG7hR4iYs5IyXPataVeMNVDVPq+a8vJKw8pgUf/Pt8eI1aSUy9MfF1/mGaQM
qC+kUWKbgLg5W2jsFHAkzFHCF5snAq0SYc08ZJQp9DIAxpOFqH3eANCfUjHAiGdy
hckVXRsIDiTOQZh2LFMySSVOxwqq9TaV+oudJevc06o1c+/AuR/I9mh05mq/RTIW
Dz0nqj7PWbqSMjEJhCtmo7Et1M3xevpDXW5EsSc9KP/9HLVuUoH9Gbkq11TPq3BF
Gvnje7VlMGOXBQ19GJOoWP/xhPhcqLHi/VqfNMbtxf8TWbAgwCD64/s/2g/GmjwU
E8OVLYOU1zMJkyjQhiDeDjqKOWAnv+zm4bOeFIMghH9ToCbYWqQZHmMnWTMPWcDC
GgIFp3Kt3DCE3aL6Lz5mtdDHMJmVFhrs9ztd0jLdB9X79CijsU1oyPayW3ZgCabn
TvPAUC2O5ng3jycuaCwYCFmg/HGychOcfeeJM5MMFSFxq2tU4w8P3bCxI4USYgir
h3m5Owlg4GECZpKMDUu5y5fIMmTdIWnLLnR9UYml+gfh548uHPOjgxbvBpgnqrjt
no7KVbfd+CK9Y0KrMbRD1GSbT9eZBPZDXdCjFXzAU5NFiBuRKmJZN3ZtHXbGF5Gi
kcHbnrpgOI4XJV3WOepPRW2vYrFE3noAhcU3yyHy1noif/BNLL59EIoeT78CO6E0
44gATO/GCQAYYYJeiXptkoQh4q3r0WtaOC5kxBfnmH+u4MpMOxgaoLlYGCgZH2rT
8pzbx0egW82Y1VNF9O/PIOfoS1j5zQ5dusWaitWtzZocKSQXNDkeCKjSZEvHzs+J
xoKxB7ZP/wQj2cnNSyD2Lay8sRaG1LR0+/JBoIPslbLk7zDkhjt4GaPdfhn5sxhZ
zUH37PIZk0wUGDThyuLacWXnmlwzxv4AoaB7w22G7nGerO98gJ3t6GOD5H2X+j+U
DeMTE3NCnRZPEnsx4vDQGU2jel0v72CR4TljjScHGq2qPv687vhf+/QAKcwKunJv
wPJvEr/xRp2+zKEJVoW9/kdkSVhX7/ENrdA2NzTWFuNFCnBKuU7gE3fXBTCjJLXl
WgAUlhqbgo30TH55Pia0M7YyGjKXYEwD6n74alnvoBR7SGITMtImdnhXWud4JD5x
3tvtJOarOwy1fy2QHm1p2jnHKYZ+GQbzjFxg7fGhdF+XGgT8v+GgosaS6lXNaJXT
+K0oz6mp/+0ap4rHmIOzJVynd2bITll3oP6nk09iiXUiDeSFYrEbZyb7yGlTdCH1
4/xe2/grLoR8fjLpPNDC5tfGmSZXo7o6yNo+rkmgM/SpfTwqEsrkDXj1h5CtYcKw
rhOZpNMEB8dwyIR5+Nxc6uJIH7pb6cMGK4bv4VGb1ukWrFmVukAenZ7XQwmGgdaj
oIKoOy+4TAwbh3bVlvlylfgGyhlZuo1H4jg2GgUcG9SJaXng34yZ93nX4DVBY6UW
yHgYcR5d59FxvVg6mKoVmbSZ2vZcASsRu2TxftcouDK8W68mjsOUnG1NJe0i/a1F
xWKVc1mpdfd8FKFEYxXwy6cnhHq8YZajiZ74Vzilk4mVrTcw09z0mOOel4It/NNm
K061DQCzpiUAQqDD2l/6xnQKfQJoekJ1bp/dAJP81ObdbEv/yBNiNl/SGP7EUV3M
dcbwLL9gmRr9NaUFYO2sh5NXmC25I+6jfm53LD3FZe14yH+yd0y8SQOqz7jxq8BX
ctcqMIePjoKTC1peMjYC7xYJsQHyJusrde34+NVa4eGjU4cR74RsK7FjN+l5TXhN
KHznZPE5CIlhCyOZkHR3B0W/o6l2LgsqNQ2vf/4SJ7AmnKjkQEkA/YTQbSgjunPp
2/MEgmgYQFKZcSvs9IXt3S9s7dGAjEJwITyY7ti4NmzGFKwppC7V+4HvZuKcuFnl
Gl2b8AUyI0bHB3xTh/PnQsDeTjwfesTgjm1veCEoDv+iEuMd+v/vR9KqbFaXHXOj
ELB/cMmOXPs0BtwOWZ603WOCFODeKhk2l41E9XEWnB3PznzroIxc2b3pYRDIfe4L
qRTOdBWk35GmjhMfuCg8fjhnQjomq5iUvGYzH9nVNnszmZXh1gbOW/vyuuGf59yG
QKm1GPr2/To9/YVrOHRNT7aQqAyVB89NHLxL7iOHBv5SSgZYPOCEYjjIJhPQ0JJZ
FfEQPOCnKQM7EjnAXLx9EtYUPDs5PSMj8m+DI92Upw0gjxkQwRPgU/anFNjqxcC8
oM55Et/i5CJVMJ7Z3QsLcWMkXcWCwuGSgQEIMur85dfj9ExRYYEDBzC7dElPxrfs
/sAKGrbmGjumLnlvAICMw9+kUyR5OZ5wZB/2OnVVLgIMkVCQSKd99zLgOgzXXDHD
K6GmSDaYKhb84U78izwUaeaEEYbSuwoqMM3QjVyipKsqYRD+FZUon5Q2p6QvBJ68
d0lwMNyVC15XPmVt26cPL+BxhsxGBVajvKiqaLILLAkn2mexq82Tds5oVF91LGMU
DM09xgUQAZ76gYlUQShdDlF3nImnGuxEny+tsmlysSqsHsvnl++6ioX0qNfKzYiO
MhusSpqMfWUvQcTbsgNpa99QW+Awum6yMEpIYctYJsxPwtahRggGFQmplID7o9jt
FBAGKUc3JuthAGGnI/fOzP18g5VfdPp3tRJ5GSyJ0gEjlcExh1XcYTBP1HxZwLY+
KQCSj9TfOkaVd8BmaHLrDFnI2X44/ZPC9Rs0frzd33XoKZbWUbm0GFWkT0JYxVyz
OMDPttvKEuAhwap6eW8zZO6ne+8mb9TkCcYVY5jKrUhNLR6Jda7elj4tmHi0rzTS
SD5OSsS7euH0EnE2g3usf3WfBqnah1weOnRZabp0b5AvEj4oWtB8HSKF5DkWIP5W
wgyHLNYNWmRgvXi85FdTM2EejkCFcoW+nVJ2639hOEVFAOPxyoPdoxoHXigVdnIs
9FjHlDSr3ChXcwtfF7d+wjhku/wZ8bZ53Su/CAOSkJGHmWoex4z3BVQncRJayZjg
V9Du24uxw+/j2bbTI6g7L37nJwpzRQwDP6h0DQngwPZ/lK1RLZa6YhEvW6L42sDT
6TO8/UEEXuyUdyYMz4Yav5FLEol3QsbDygiUXlADPuSqS/WhqGzJzWkxO5MjRhCU
V5BLkuyDVjvmIurdNhtOkDHRpDxrld9D/AG6Z36OBGwifCh31ooiYUrz3YRjI+iM
/CbfE26RqAYGhntWoM5w3fyEs0lJZb/x1BpZSkCNuCR0uZg+ICxyJN92Vr6CnxJM
SZ3/ErzrMywSagcY5WEMZd8+eiYySP8whBmax/HlsO8YEniSkm3wyRKNiQzuXVWg
llVo5eBNsYuPlhN8VVFAv9koi2Z3EG1LNPX/lrYiESPX8qGhizEkCrUXwS3hb7Fi
s7ixikDFXS0Y3qmv1mQt43AvbBj6cDAWVFb+tW7WWHX46Rp9+SzsyCa4NBQNndjP
Oq85CTZXE4yU6+AS6BW0orH63qHi3mOEzwx+fYacA/AcOwmVTjnflP16CLuwkAKC
Jg0JdNonxUrKO22o9RxkRn/ER5oUU5m1TYzg5ee4y3LH0Cp0Jq2lQXf5dLxKq6dG
/tnQjlR9gtJSXNXHRUAUucMEz0zdIL9EJ7ytEP+/6kmx1dh2yZ0LKfByBlQG2Jgw
xbzEUhqHK/CXKt3GM6xIPo/UXp8xXYcVJPlpFOQYh0ztoe/8bfKXxxM8OzSoBQWI
eNZOTmR5eAah2lqEzX1C9gOj7YI/ABwq6Fx8DSCEGAQ00j3RSfM1MTkKBtfVAiFx
LnNCM7L85RScYLzbNjhZojO5k/fnnlgeh1jtf/G1b+xPMoXuqRTE/w3ivEmF1eFa
mkTgVh2GY7qLa7etSNOPS2NoolLAId6EYHaGxW5kBu4lGk5UsdBq9ojaTq9BVKz5
NSTjtpxoiaGSGp92JedkMRa9XefnMI2zTZJrRNv5hN1o+gwanFiLOSjgFJjCwLOG
KxoNk++UNSmK1mVezSrUJ+2SdVaCA1LLkZ5EkgFqdjqVE6BIl1vpD2a3OmdJ+M9L
TW7w/Oxo55nA3Cl5UWbcm0acnvPKURaDJ4brjl2J9cZT7iYjuCN2GS+OaECWQu51
0BxDreaEmhgYw00XVLA7gkFaymxdqoNZ1c+svAN0dBtbinsY+ZG+I4OW5CXTxOqD
iO6KgiU0zQQK0hX8ZASaSANdT2eDWcEPWAfDsgoBCUM0DGOO+epJfqJZWx7Bxyi9
rEvqKwKWDfyQoTBwgZGiNl9JmM5ufIQiAmA8PSgfdzPwkRc6dLrcYG4fMDLWHz/f
yPQbHh13f6jVXxEbd1VGK5qNiQZGLIHvRHdk8XY0WuD/bXMhJTuuD+dRqfJjxudS
ZsH5aw0qcigHv8NJNUxMq15aAUtsBZ8IUo70Xc+QwhXi2M6FcP8yhagB2C9/6wdU
rk1T9Yj0slF2s2K0C4ahHWxr/bC3liw31BDPhHdzaHjdtGbGgKs0S/eAA9u/DlkS
w6cEnkubSVWUgAYHGx5t11teuxGc0WT1kfOPfpfzigBzwSaWkGNzJLA9YXbd9MU9
DP7TFAs9RJ3u5fKOECo2BMHSmsVRrq1jPqyioGUUfeKWaLopDHx8MEMes/2g/lFS
RE48fjSsQheSksZvuYG0TNVS0hDrNIBqP8mx1D2GD3/PgEG6PFuJborG2t3JEkP6
Dj9R87YKzPjsE3kv90RRhAxVtB1bsPCNjt2hOtHVmgssjBkm9etQ1B0JDS9dWEsj
/Zw2o8G++DbuDhA7IkiuZUYz+JLZWwhzGeNa7JL9Q6ruMYMI6H9JLLcL9F9IHWN+
sbLwkOwVPPfY+fO/7zz0C7q5QT1St8bYtHEES4RW2xiGoNb6We2Pv+NK5JMYo4vf
tQeejBRRWKpqdKlpdJoF9PJDcTosB1gorJJdpcWPqaEfLPNZxBrbgaIuaUmWEHMZ
o8pDuje6HLp6gZfLKHddHA8JK+JnxMaAtHfPWcAgqHghHJdFz0NGY02L+CSwDxIn
a7eUT/3QkOeyyAIlwLF2rt2/aAk9g7tgP/J2thRBtvYwpNN2HKr9kWgSDnOPUDRc
3BkXGNaqP8TgG7Gw3HMDShl4UCtra3i93kGLuGGo+oU8EtybgEKDMWns/NJPlK0f
O/TXzbAWJOgdZs3wVv0ZsKe4Rl0TmdFV2S21r/g5JflVQcJ7GIjb9O1cWVVmhqWB
XHH7s058oHd4aMbwpcOuYDexrZOaaeTysG9Rn2oZQ50vcVqhqvqav1ac+DxddKs7
JXrUUrM9Pkw/Jn2ggz/agWrUGkqyEfTp4i4nLD3LP+sd1Bau8nhT5O86OK0MRYQK
BwG87ddLMHdDIx34KSmWbUU4bpFMu/26PUne9QbOkXqjjpsribcmTfjCeHB4ITZB
Bdz57dF30KabkpvVMzsg9ohFOVj4WFB20ZBcJLg7KcVb2quD5Djxefjqs+Ov81w5
+3jI/3gUk4Xn6se9vN2jZxsZ/8VMHijOxa3LZR3bEMLqdtXObxGa6gLQ7f2Hoqm0
ObSTi6Wo9JpCIta72UdxMZXbjPb38iAdX2ob0TS2ufHR2lslmJ1nfq8R0C762C/d
p3Rc5oAznKtmGPDpUK4AJCSqtAWNZ1KZF12F2AvW5ykMG/1JMt2mLgwSn/v8uLjm
LMgQZq1rIoTW5xuang60QEKxKYgp0IeBEIeIFu8GKXrk+MbROvK8UT5fjwi7CboO
lhh/xfUVrmV3WwxyYyqN07a9+JLf9kQQ/p1ZUkf9TjRQgkrvwvkE6ZHxctcoqFGf
vKRl1TbHZB0RRImigfLQVImZ+bMe9iveLhM9HOcyWAyGoTAH98vArlsHAktgbgD4
09VHaJKSbHCekqCY6VjJCEqTSMK9pGjjfHqs7pjXOUTZHKitGEc5EmZBZxjGviB6
MMAwhIi7K6nt/lThWBBWf9jvHv1hIKGnbjrjboI4A8P9lefba2pqzD9/QMbVnDrj
unQdPZ/M6LWzAs+qtnuf2S7I8O+CgxlR4v7gfULnsSqzooKiuh4osdlUk/ii1f47
Gp8FKQdE9i1DeGqTu/72BmMKl/712ilX4DRgyHuUg2hOMAIq0oWn2bGzi/Va65hn
RUDoI4JZr0AcL3bTbNJtoWZXLBf+rpjTIvui6IXo9txzfGg19x1wysuruGXGaJIY
lc5FwsBBfF8hsYGcmk8Z36jkkTxKBqKMcsDUueP1q3jT0nnVrUR/V9e3IkEBRJkN
N8ZsIlqTKgrdUZZSxLO9H7hJlGPLab3zONEERTNu8PAOzomq/ySjskBgo1e1hdfa
HZwTm8EMzaxOcSAP0hoR9gQt80rTtkJ3RxbwoGpAEDF1DvECiBEb2/xMgUQR8sg7
xWkUK9RN4yU4NOzMFEAitSktwnP7j2YH0wvwDw8CB9DxO5LehrWETq8zxJhYShlG
C5puSCVIOHOZ51iBG4MY1rw91gjEixDV47OI0FbEg/Xv2ckU0AcUOQMpbE5bQ84B
VrEWBedLLJzaSpZnmNdiV6RdrfXqzFAFzbVKfC+bMPL8bIvVB4oBylpfSgqiZY03
5o0R7CYsh0KYbK/KD5PZLPwc/aOVbiNkIzwYWEYKMDsL3dtm6ury1+oCB06Ztgqg
Yfe0YpdKz6H6UfGK0aQCTdykNAwRuWlLlG3gDE9ZKoTjoci8QN0ZMmF7/xfO8mem
huWFZm8LDhoU6KfadnaZx1IQ48Aht4YJyhobZJf3eYDXPGtRv/JH+rwNSCDlmidZ
Kzi4ehMVQDSBFn+mL4RK7JbiLZnKSx5JhrWe7pmPcqfzD3494/ZyplCpQi0EHh9q
AbN3Qvbwsgc/1VNirPcXHs4ocVGqhin8JC4psGdbzE1w0+CsTtKA1JU8ZMQCb2Q0
J2kK0TH3xaFDL17gImzz1V565zSrXElmdZHcKL+5Zt8+eWPrK/60aOsksgG6L+n1
uZleHbi5+pW0D2FuiG/fYWS74dfYa1myeS1L5kID5wa85/LvVlTyuHrzN5wFr0NJ
SQFjY9gHXzmYRfEs9xkMnxDrHGC1S+4b7af/zKWCOcYcnwF5QYS5YFl4DdMpDSzE
nFabqWcwzEizXwIxbnobV8IpztpOlEabv5Ur0WfQb3T3M/vvBWMZKTALpTqgKNhw
zpYEWWc7HIBMZllSmgTfm/YWa0KH3JUU45pcRKCzedPEecglYdMtxA2eF5BjPUqn
mvwBoYK7k1QexzDut/zvR6tfuIIBNkjX4ASmzA1/rsW7ixHMnXIgI8nJ8asRm9eA
bsEdrCnQUSEKeGdvRUzTN37XOp+WdYAKjudn5A5ovc3VLAcZT/vOSvpQT5BlW6hI
r7QETasODIJgmGgg56TWg0XNDCk0XVXeyVAaw3RW/RmmwUiYKmv5mvsSlTVsb34j
6qyypKu9DUUIEM92WEOYSFsGKF8uVDKqR2KPHYgrZLayVvrJy/pxIexlGyDn/y6A
G6QbiwQHowdMzdz4YEtigdPnIUSwbTv5WKKhGKSvI6/SK76qmnwXygxvi3oHnWcn
MaVZs70fcUeh8gwifoLgeE96muBPHrGpgg1KdRw6JRnj4VnQCgmfji82CLDMirML
92iiNbJX5qPcq5lH45amTluu2CU3fbXB3ge9v5f7iCHofUcU2ZmoM4+Nxdvt+orj
rIY1HbZz2pA/0R0AKHWX3PBNNhUFMIFRUAETm778fYONtiN02SPYJjpYEZ8A2VA3
bYxJYjhfKhphQoR48Q1v0FWxcYIlMqKyCbaX9l26ib0wP7EEVLZmxHyL2Vrmo7bX
kCNoTqDq3plVdLx3AQoSkE2s+BeUTlKyXzMkKgMKEtdOKbLQauX4aWc6z4WhWhf+
xTf5s7wOtIB/M6Auv8Er6uKz0dzSgioDdIWCKJW33EhwKYvPeY3i2qlDscVEfi0J
FDBF3nvB+ZQaCC+By2IoBj4ymY2UScpKnipCuGVmAJhp9dSaue0MskVPme0266u+
mityO4ZNTc8HWajnLCEcDguW4f8JOZqrgSdKSXODEkO/lg5lUwbj6TuxiGfybTRz
KFD2h2LRusOoVfHYf1Rw8YDfTwKQh+nMnqBMMqz5WP8bmPq7JbP4R+HPWRDlHxI/
UGGXucM7G/bce0zp6nKcoKclmUX9wR7VX8BtFq6Q2AspLJImf1D2GvElnb39nsz9
Ov9jki85r7NszZ1hMwjkahZje5qsuUdDPBgm2mxLNVS92QehW7cPEBHuaNlka8jn
rmobGmAWfV+s8huOSMzEn4EsRscXN15Mi09rWRHKLrDgue/qtshF1LQdOuQyMjsI
0JowvjMrZui4RjSm/TYf+MNUGoC/nFoAri5++JYUsYRmRTbbOBsnGI9UMhrMUb8a
D5I0R/9xD2Mg3AjGwpDKoRURCpYMzPoAR02LECHrNcCe/BYIOlzuyCp8caKWAUif
co+g6XLD0r7zUG5yszkZST3/JCNlf/8M9BsRDQGlkhICEn4QndgUoB09yzj1wXdH
5eQimiLYPYFllebHNsE4zZ1kyIocc3ncBeoa7pIhzFWYCPkblrqvRQLQRpfZ0U1y
d3tofGX2zO77otuzV5iX9sMdpbFLOuJi2RLrojZt8YNk/BTPtnsovn9PQEtF+/vI
hfzBpVNbzHdqiZ9qzugISHWTCXa59k+TYbNRIcsSZwOlXakVp4KeViysZ3gyWeUe
Wsp0kq+fOS8yapomVPrslKq4o9bGiQHrfCphzvjEp+tNZxeH1zWY6GnsPA1qgwKZ
a3MfjhtoutRUBobExpK+vSePutgtmweYHTGJqJYnrUSU6BKybdf/FiogbsUzsa1C
M4VF3In4H4OdMhSIZNW8jQv6j89KeVzLq+YVjGC3KDJyX8qW6XexFqXTnh5DvLCN
oEv1KNRXBK4EOOMgkrPHiSM6aN8TY/pE2HQ8O5o86oBlSwJudd4FThIEVveY+paV
4DK/tJqsC8zodgOQ0hPiBhY1kGmdclmLDSz4vW7ogms4S5l1KQcouc045h52ZFiZ
H3qNrl/bzQANFQeh5BqKwToiBYJ/vmdNZL6MqDej22d1ZCo66SZ576Bvt14Swwpt
1O7oKrY3LO/MM9RfEiViu+FPJ9Rvb5DhGQQrsU1dqtDI3ruCw0L5VOQCOcaF5+Ay
I2l8kYDB9nC7eW5YfSAj2cDadbmOvkdTndiDIm3MU+Uumx4Ca7Vxe1G2Fcr+Q0Md
OS9VBCZMufUdHIf/wmHoeBMDuz7Be3VsGA52XrHZAmQJBxg/l3stxny9K8Ianlgc
KbEZk3gw2GWZ9PSQCQVFJSJD3XgBPCTc4JTqmD0KrtNJYT2MIRH/IHkdZWr07Ebw
wKb9I7DfxHDPTGdaGT32eC233phnfyeZdMwISaqfV6o5vCmAdhjhcKu+j78vl1vR
k6ZmSwnU2DAXU0eoEhPTnOsggaM7KK2zu3+RfsBt0mG9SJ1rGeJnpgz8JTiyZEkf
x8grlW7/EMEFhbELcOefl/+CxxIEi3g5mMa9rnaDg4gWTGrFtNsacv9Ky2FRwdvT
urFPLXhYBTufCPX9KJwMIH3Db5WJkyooVW+1EHfPBSHShxyz0a8KF8eQsDUGuv16
CRMcl11cQ2VInU496yMDP6gobv2D+yq8PTa14jQjEz+naaCeBNC4xbXGs7EoPn62
kaUOI0h7eEIWLFf81phpE2sZPtytWAtEYoFYNsjKplMHZftTOVG4YQ/erWlOaxMK
e3I1mgKxRErCmeBC9zgh79kP/Cr3ejng8KUAjRtmgGoX5tZo3qsijHdO9smvPdyV
hR3pxVKpYkf4t5sLaKx6Q+kwS2D3S6IhI1lwnQAayrYDfD5j45eg2djn76I58rXu
tTR8/cWCKs9piLqO16ob6w2u/yJTJR+4ZzLrkk+ytfePQz0esHfkKaZxNo1Tj9Qf
4zgnKefI8QXMWi3STGbwJ79NefNUoPEZX7J7g2iT/tF5wh2n8G/t6eYDp9JBAnRR
+eNDTmJTiuwm6sWiWpbhxYsx6QzYYED7e1MGjJ2XBk2+SNutVWcJ+CwV6bCEEL6f
oGrMoX70qJgrgRoQzqU5EV1w8Iq4t8gQAzjrUW/mjxvPSrZRd/gerdyJSs/oEbZR
IhrKW67wgP/9hrAoiolw3tZf00zVw8Gum3x+rbEWyMg7KUqDL7ZWgx8mV8havHrL
l3n0HGyPDM2QlN+1KdapQPZ2KICQAje2QUIhUq64QPbxOf4zIQnMOeDAaQiUplVj
9X3if8+igIEDUmP0Q1hi4gfpqarNljfXFKtv8J1EBO2NHIIyr/swtQodEadQxMHS
k1SX18aivrK0JMVSwH0d70kAr47YvcrW9fhMqjOv/spbdRgujWu91cMr4yUN8wQb
WKBMUmemAWELM3XyWrkGA6EG9QYlyq1baOlk+JzG5Qo7c0hlUIWqHEh36xgr4M4Y
znvZIgEqdt8Dc1qQ1tkCJRvMJKVDCtV26r8nv9R+19JnL47Lv8lPnXqUMcVs/dlE
5cBs7jeW+anwRc3JiREYhcuJ5KvAZjkkbvtKmslyuXNAQKNfTPNuPYQ+UmYqrHPx
CbZmAtim/Mj7H+ioPtrG/M9VaEYxBac2YBXcaXuY401bV5kjWshHUy165dhfrib8
3Vgl6ijXggx+knwQIFoC+lvKmi8thlQdHeQ+e+oo6weEFWTEv0/lk3b91gPSiPv0
6IWV3p6i/E5ytqfk+YDNei1XmCTB8eeCUgHYu3q/1hQovOnhJHZ+2HFx+rU8sM+w
i8e8HQ019F3ZC2ztMG54tBL/mfSVds/b7riZzORjJYsPHACDgs7RtE6eq62oBGY5
tDa/hkWYrBTq5kqCSXTz12VEnlaWdb8vJfhomrT7IdQ/t8yAHWJBEhJWPtiXGUhW
mmVwPPOkxV0/RbbfZwgBEtYEXreyXUzNtXHuLYu8Nif91NTptV2W4vpIjAcZG9F9
daoYdhSGa44RVRPkTRsr2PBItc/HNPyZPnAaUX/VmyOyxDlDuAuHzHKy+wAEqgFy
0fUpqV/9JWDe8YcblLVrWpYxKAbxi1geK2xM1iZwrcM7zR14m34wRN+4223FBbN5
tQn/jRv4BGtXtMHDFKHSHeuA6BbjAUJkO13gfYGwvfyix1G4/kLWAPk5QtdtdpXv
bXi2GYFGOFl53t5UI2//YKSJ9uNVPBtcIfBWrRfzSEcIRRjCMQ6Q2pU0BGYpPO9x
TXCw6aTbYsFyO0WA2LlSTSOxL5iHJ3tazVkAR6f5wM0rzUt3WBjLoRVFVMJQGkmc
FsmMarunUMRvWlJi2gWc6SlUGgXN38LhFNjvk755VRPidcWy9+EepLcxAssxbvcR
N3BCamjo4xtxdHldeDXy5Bth/Y+o6Bstn2mOz7XJwxbum08ntUwA8yUiOlWhFE3t
8ce0T6wQp4EPvZuG6wW8J3g5s+2+0W05WKrKj9vyTCr7n2fqXu4cwQOA73obvsrw
8Wv9rbRNfdUgJR40n/dQenZDksFL92BmrmZVovbIR+wDe4GM243kbqqmsQUF+qNq
smF8i+xYdoX5FA8JD6sFx/ID0d/2QRdvotPzQDXJEKSu/IOkX9dQINvacDG+ltOY
fQZoT2DjJ5ajcF3zx9fEJN55Owqj9gzQp9v/LGEy57vpWiBcX8EBbD/Lq20Ik8tl
OaaROxKBPCgxZpAXhH2Zs/QRU06bSO3MhoJEPJj89+WuY3WCXQ/giNIwp85FQo9U
5D12bL0EwR9aZNbdo0+42fkAtnxQALMJEBJnLryMU2bZ9e5OL3KY0PElNVDwZfbU
OhNGI1EA4TEZ4jINQv+u5zyivKAHlcW/YVreMzS5//UADPVQ9ISz8TWKVU6wmOP3
Xgjqft8RWhN2BgvBr3qzoy7PWWtNw1z3nGh8S76Ebe7XCyhNrLofUvtJQ77QC2t6
+cZ0ujkXE6lWWaZfFFlIZSYVOU6uhRSoWzY1waU3fr0ExdICWT3TshEskteWigTj
6fkx1J/6BguUwPm3hQPWEKQu0K+50zBAsoQKUOR6CQ91KOXqOR7prY5DT4khSDfZ
E3YYcTfeShQUVoCNOrkFBVwhm3sbZMkLa9vCWa33Qs9gFqqhjAyXSzDsFc6HRU+w
0/0La0E46Xb3X92NH8/nk+ngqkjPliNnxI7ZAJUih9Y1EWMbmDD+lcvuXFmBcWOa
uj0g0AicE2WLboHxn20PujAV7UZyH0KHdDa/l22PZmmOdhJRLgB4Dv52fXKuOOJm
O2iqhalvWvRztNgPsQwbwV6cDljSXUs4dx+G4isD9I/TPnJQChNjHFGbYx1pkjTQ
lxWkiwIV06EGv6C1RJ5tAz9D2KAS8ZzrQuJhiUvpbkW3KkUCwoCZ93OHfxb9AkAg
3ODrGvCwgzhK36IAuk0iNEsRWeKBNUzW6KKf6oUumM5XzhZ4FqaN6qb8jmLrpIoc
hQHe+KOMMYnR6sJLe/Ct1tZj4xP+uF76hP42olQPV3Yh2OAvgywCyyJjR/FDwU1V
Z7r+f+4NfWl9t9V85JCzUQlpIep3wGW2wlRlUZQmIHscd9jfZqeo2OX+YqxgzIzc
Ad2fhD7Tf6vsYgmOqLzt2QaQ4Y8h6IdOlomT6B/GFlYwXP0c7EV+/CT5salW7Zs6
/HserP45KcdCzEZaDtubgn5P/ZkO8QCReH6nu8GYQdvqGKWx5nVlfx3b7jZHM8g/
jSpda5Pdwvuo7guurBE+GbrbJyG0666LN2xoBbTts9CdjqL+dnesumZbGV7QpP6q
Pc3R3pzrserMDcHPHv3nugiDrgl8LPitMO3Vnt4lR7NDjuJCAjAzbxqXE7CqXl8O
sC8unZcORZ8TFvxm6KtbPrP8hug/Xwqo72TIdu/Ro1t9Ohg3pvI9J8q56yxSqt/9
Mckmwj1UIjP5+xGkW4WjpTXPXBI7bP7iUI1tI3PGr9UHy+2qvUv4sfHTfM4icmb2
dg7GF9CSiAtkHoG2nL6KXkZFejYIxb1WbNI6BprzF1ELHGn9Sn4g4ioxPRrI3Tf/
Jj/Uvtpq1Du9cruy62r94zxrPYGqlciuWEgJGaVSR1IRafBMP5tHIlfHF3fFM6A8
InP55z7TshfFCX+QxABG8R4P+WPGvhj2GQ8NrFsKQ6/gmkRu/I54bPCPQWJgwwW0
RJoTgqVznmBqYeiE9e3BfH3/NzkHdYVJUdAZhhRa3sQNdgeOu+L66BryxgXfkSsE
tIj4wOKjW8bhvVzFSefe3eQun3n1M6vV64aLq6Bkse8sKjWIypUb/dZrQcQFGFXW
rIuJ4r6zBbcV5mMX6NzbGcxWrB4b7F90YVjGEPdWmc8f4GIs9doqcRPB1dcuP2yb
vqr0TCDJGKSH9pMuK9zTu/4bOPBNWCq1CJGynigDMaasx/qaOMDN1J4hKRyrDfAM
EpXTv8NG9urKmCVwrMa+IJLWy8OsJXvsDLo9R81sZHXDpnkUIrrq4aUzY4WNUw7z
wgYF8RQPoR4NXF9Ikc70/DTB+DIEI8xPIMQD2LKjuKWuzfNFHXupEElbRdlGykmZ
qQoYt9cayq/+x1tGN9l6gZH02+zEzY2ab49/NP3oUtpvMNQvxlrqUMSD15aEzqua
2HXmN6Z2LDAkZjOs54dxW1UOUweCndGetfxX+kFHaJS3p2Y36R3oBbjzBC2gTQtM
QN/WKkHfAVSdXc/ZyE0drfRmQJrU5ksPsNwItp8ontVss3aUfNtXNGa2cI6qtPSp
RIeWawj2UXgFvvtpr+datcXLc9Gt9ztuM3VaGnUVhtjdUXEaadxRjpccwJbIxObk
7IbuyFImw15SNVXVniH7Tc8bl5P5cLqcx0AYyLqXT5JVEOt1WFwszIUH+9+a0RCw
45jHv/DqwPVFDYFr8oTjgxsZcLxvszRzmgjH831rEo3f6bU+ozrLyPtCf4IeG6//
/DnmZUnywBO8mJq4Munv3/uz/5CWTGGn5WtfCelZo1VLA5wVD+9rWI5OQ0pYBQdP
K0MRPPdVPJWOA+wBSzOii4ouELVa7YMnBs0eDUCm/6lC3+/TXV5BIii3YjRK/889
cSqJTYDJXmOScB7/GL/t2Whf+BkzEoVXuBhJldIioasLomKk06de+sTUns00mefc
Pphtl8Umg4gNc1WX7pfgJPYEEuY9DcrJDkz2rPMOgpkOEi1niRm9fm/GjGVkD2XM
pLOodRDmTlg0L5cJYeZmIsPC1UgPQ1Ah9Kp2gL0ZM1QBr56EbH6clQ4IdXFAGnLH
ELtDJMu6APpIEiAYmLg/ol5UOFufXiO+FbTFkHyM4AxxFazEkpTOxQy7IXsKS8SH
r4BnXxyFw7ptj30UFZF4oM9pPqinnfPXt+GD9FaOsDP4jb118VxEyffbFeezav3T
Dwj5rA2UazVeBCuGTf25v3XSeaekzUSdjXFVJyv+d/6yWBvCuLHW9cRDL6JDDCHV
xDXDSDOGUYtw5irZUb/mv7ieQm2HIzIlQ78sBcLPWHtZ4NTI+NmXSrUCDB/NhWy/
Z/tqjI2Zt44kKs1AO2PAPSOTKNH6HI1AbxjXVQ00xyUb96pm9bWt8ZMYFLhK8rG9
KcdZL2I+L1A0Zdn5H4a4yE0KkR4ALRWLPINWUfb6tDZghfCjiL1acs7ceC5tvfks
IHtl7aLLKPykUMBNSikuts1+G04myPrpyN4IYWyfOg14PTw40OrcxhWc865kHVUA
zuI5M0i+O0/84S777jck9KVBY4Bcu7EAq87iElxBeMdPSNb8u17TEvO39cMYORrU
VFNK9NAjuRWDr3p9rQBZKz9d6ytbfQ1Db4mlitH+yR6sbpxqPF5DXWyiv2DFBOhF
PnwnkkUJzWy018BCTmG3nbNn3OzWWBVj6xcvTwowlMaxDEPIqLrK2usnmDkSIjkR
pfR09eQrbita+vV3UNU6aw6W3f9fESmOzdKX7hhb+Y9hAZStI4QAtsxTaigxSR7R
MHK45ZLhEv5rzaccqdKUnKUvmpGw75QT0NYF8V5yLwsv965mI3faBqB6x2shnj9l
rCb1En0Jp5Uoxc7R3X/lq3luUpFzuPDgM1TG7H4boAmYXd5q3I1aAjBDbUKRFW/j
TdjYc48UUBrYme3SS8dg9/lumG810emZd6RDy5z87Eui4f3ZQFmUa1kIaexuM2CH
NBMjlSfitL4nlHTFuOfpe3MfuXBTxjClD8FmWAq1UjRry0QCugGDQxZ4HOnMFDxi
+SrZPtp5e207jMoUkzPOkxZpMu5DJnkrxUF1krgnjXRil5rp3dCUjhE79Ccc4r5I
ya/lVBr7TO4UMv3NR7MpIgELsYx5sqahFNfyAklgdF+6YdEg0wiVsiQj49olUsMH
Fhpa5W87dejsj9p4nkRpMlFD4tJ1rf6U9eXnx+NfW+HxDc9SdIvO9AXVfst93O4j
cO2D6+8cYuFGIkRL7TD68OOHozhy/zsozWkgCw6W/j4KN8BwRD8m26aSvYATCN3c
gj+cj26dOBvACoLWdjiLage21XKPLxr3817c1J0bWmb8/lztgJ2G5K2pzJ7QXAyC
UiDKSr96dZ3oXt2vqEdd1m8wqokPIEM0lsQvOJpsqQRhQBbY/mwWhLFHRD9o6gSB
eOpq6dKOLUfZp0MCn1nmOZ4GhIHwcvgRNyl77uuUnaNQdLA2CwMk9ELyEXHWH8Jy
VQsnFoMHq0mjDDnGZLuUX4GooJZjd1Y+owgW8DnmCLk1G84Ued97q6Kf/mcEyyGb
f1Bwe+86193ofi1kf2Fnns6ZQc/XR0IFGXhkI4JZegGHA18IhMEf8vMnyC4P3IgZ
lt+h22b+Qziv4j6jYuKU6byr6Fs86Q3MIBRxGYGIJtlR3ADzjZFNUdSE3dNb9JGA
NxPKeBlTe5pYdTXPxXMmC5Gn4LQPJFhvkjWFe+YdIJdo0/76qdYyks12vf3sr5cD
I0akMVprmvigi2ZyijTVi1daBLxoKmm2leXcRo0Wf51zw+E8HXBQVgtnMbyI9QSf
xwVcMfehg7MqVmlCVlptBdTzGmyz6RGDjMrEFX7yNOgPgVuQrF/TU7aXruqQFmih
XBXPQYzvOFvfiZhPiBMliRDYq2T1gBtXxC9Jf1KrdsgmNvyR2ryCM/NJ/MMpZuZA
QBw9IB8PnwHdwLd19I9Vp4HnmLYaiirkrOYIuDtZilgEwaCkJwp/4C3y9q4GIYzz
zGf4x6Yg0qMZDvPYmJE0H457WYbpK34dMOCaZVeuf/8YgEbTZVN03SUIqFWREzQd
ScDTIy0znE8pXmUVxbFyqGkSsHA5qa9yv9aGo23Fu+sw+ALpkmSGL2e6RUihixlG
xIaVJdmiu6o4GqrRbmSPvGSNVypq0jN2qemvHQlNZRgKBarp20ZihfeZ52E0tzcw
IAtdje6+F5qwUT+pD87BMxU3U2+jBJ2Vd5lbCpTTkTAoVIMJRz7HydyEKtbcs+vY
peDvISP9S905Hi+I6HSyfRYLQFmXdonAi5eZoNKDdrqMw82uRQwItpXZ1NK1dBP0
xVzjWfCbbEbkbPNcKQacdsHaMwYhBb6NUWxgQQbYYlUI9nH27G62EtafOAcJmccr
rkCWEqXVQnCBT8lJj/Elyok8Oqv2Pdnk6Sn+PinJnLXcDPN/4VM+3xPoNaweQYer
Li5sqizA/T9EmU8oiivEn5BBlgimGwz25pKGr+VlzxxF1cUMlalwnW9omOi6jEdE
74o6EqbsoD8u2NVF4bsVA0mzMQYxSqf2+6/DMuEHMCOJZ03+b5dGWbYfo95n27sQ
GRHgbT0ZFE7Q8YSz+gzpNKatbRkBnETNNnFDrVNXqdQ+dj78iWpvgVNatCejWCD1
aKTw4wFqmh4sjUSJHYM/ekk7LWt4vQxDTgPjeU5IQ01atlX4AUlNxVftn2218G7r
YoeeOAkYNFY17ZJZXgdvPBMxzxx5yvkB0OlO+ghpc/nnbjnzO1xb8fy6suyFuTzF
0gPr9xsGOMOHdRF7stOPg5rHbVNEUvW6HBEhfWyOZFBEyJAOk1c5hwppKAyz8+FN
FaKWwdfiyfG7zt8mwDJkrCthSZeGkxPvYkZCGeIcUOjqHEEjNMyqH04Mg8c/E5iT
wcH8P85pR6UzUlN0rJMZ1T3Q8QQAzU9ImfkUMDmAczJY7HJrMoGaoKAUGTvbZzW/
8HM4VaC/z2ESuz+4Knoo9t5GxLKDRY6P1yuygkcf4Svmt+5AG3sSdPHyQfkkPbM8
Jy20H6HTDS5htVaKfOrWBFvXyEBZpnWtELVoO3Ubv7yuTNSlfnDXj6MnT60qayaU
wAt+JLqFtNQVky8As0ESql8ZU/GzKmOgAhY7iBFMaAIZ+R5M/Ji7BNT6JmzKsTqs
chGXU1aF2shDsmqIRALP7ipomJCu5Qd+4UevjaT065IhKsN06SgnL/wde7t4Pr+7
xHwMpoDenGrZRuO5h/aXFahLXOCSBeyjmTaUiYhn8Y42CRsXsY8vi2S/UbfNrNQX
AdiEj1YyQ61X5xXTT29kZBR39MEMcpNIYfmFiGDbc5PAyTqMM23M8mukt5mhHo6v
7hDIhkcWEzZvctPHB3nPdxNLZV1XSX5LbQQPOnv8VjftuhbWrcKbTSRfPSfGDS8P
ycvlSSmS4cbpghPbddH5qHOydX98YKaRv0YC1KUy9IHFLdTg15VVrkZoKbIZracp
TGhI/T3bJ4n6SeqLSu5zHWK/rjLTQP5EZJbjvihOWyVOniaitW5/U2wTkZnMk2vw
w5qYjvQ5nZ6UrTCnkRP16WezTKZ1LHI3w6bBdA3bjSYmNvdo5HtMY58mkOw6buuC
P4IbLi4OqvYTIlO7FrJec0zjF/8lddJBA9XET2rDapZi6Sqs9MpMQrCvRUzZOICq
W2QcdkL1wyI3/Xx/KtC310un9cVI37hDJVhdwUzkoehdFc8z7y+OQs0EP+1EK8ic
KlXayIVEHHlZsROkEuQYyG+X8zA8mSvMqDyzh5BVv3zMlFbmbBgfGxwJrBnHn/Ma
tGlttmaN6tnoSrejCjiGFTAbWQ6bBThcD4KEVprJAQ4EzHjaeY5oPNa5iOVDozKM
LWAUiCw+c79fOzQj/ZjWINrrJXB62G3obQWwh/jPW+7ud38fSmCVjsrHCrUxc4l1
cHl5pBTfGBfBwwcSRTzthPqhbnXAVlyY4CMjd1j46+xlRq54KgNOVjTcYS01OUSQ
4SyJvj/O6z7eCZv3g+BJ3B2M7Vnll6WKWq1fX83T0KttilOVpp2bddweL2GIVv3G
LuOxTPeKrFNGhdWSEgf9Xv+nTyTmEsV9lIW62dK2wupq4RTgDBt4PGNglGX+JFKC
ZbXOemyt//gG7LHyuO8V2KrNEPPTEyuAcvg8ipMF4Gv+Oq1zzYXUZ+1bsJwEtOf1
gmP03XOISxFOz67Tej5FLKLckD+thWMDbfW6AVlvS9DP0/0jNlz5amNiliaxEAjC
vsuvp8PcfGo69YOOoLso9qpq1DGmREEUk5NwpHO40u3p2dBXIJAdDB3qOm5SmrbY
84kth9KRC/mGnuPU2Y+X+cPd/oOibu8SzVh+FiG2WfOgLUNQaDr0FypMgDiR7yQW
jHHrJt4kiaRbfkKXUNguR1weyZN9+Y+AAlPwPYtlvmigWrW37N3gQy3u6ryoweAo
aB3E2XEToGqEHOsOXd0OZJPDIMYnK3coHXkUqlhsXpa1XgvrmgVOZgwEo12IWhXb
MqX8rPyop3UHnv+lzv46o6+ePgUx6GXIAYz4c8D0ElIso5ZFCTMwrpPzEo3ph1Db
n/H+l7GBDsMw2tLSULlnDW4LzIlKINLaKE6eEJRkzLL1G1L6XQR2S8GqmkTAXZ3X
F91A9nttoT2Z9m9QzdlAF+cnLtpG5hdV89sHp/iw4xUq5ieG2uEsMwrT9lPmjmB7
o5lO7R9b5+1m7zeiftGn78hsHJe0tDto22IAeK6XshOg+wqoMPOo+4L8Ew6tZxOP
HyjFhSVQf6U8Y0h3/XMZaXCDaB2omSTuIqr9H+tBUEyT62UdkgzovIDtos5rgj49
VvXLoflCCIDSPIdWQ3C1WmmoOiykgXfP/sqVQD3dGeaM56S0SYzY80tSy8yZdS8/
V4oTej4llGysmSZkT8CmByN4CaVTE4JK1luTA4aC0I9ew2ALgbwl7JT8vNvxYBwV
8g9hwLHYJlcMotamI+ZVsc3DsMMtIFFKsGNXbVIqY+mRirw5+HgkA3O6KWqEmpt6
slgXd0SVqMIIPURTykA5N4tnAexrleI8fG5poSRXy8OVum+sJE46+BahkWuWD7JY
TItS/15KSXlZy9VSb9Flc/eYl9klkFDMNDh9ya7iPBI1StDxWmS/+cbuGSpWSX7C
T1mmGrnR9CLE8q8MYab/3C8JZS8SXuXjCqHiDgrnNwhj78Omcq9ubDDQkAhYfTaY
llRSI0//vtUXx/sYLsp1p6Qg3+icGJZcX/0Rk2n+skvAt4bWNzrUZUeARMuXt4Qt
TvriGM7sxXAwB7vfkbOu/LpMb+Q9+B0KOljcF3B3Y2X3UAM4hTLn02KpApIo92bz
XxOOgAMDu7sBXvToJKBqbxfapWIOC2rWnHMM19V68Rr1y2Hv13XnIOO7x0hp+3an
YIOJth8Pzr8TBhGbesUlbH0YEXHxQiF+qQ9dB6dUfpK0rNXShKwa6zRncA0jxIjt
pOef9Dna48+X2Fgcv6YWn7cJu2OUEdTMWBOU0SXKoYkeuN/ErOKA6MXaiZg3AfcE
CvTrg5HSiroO9sXAQW5P+JM7Sz6jZV05G4ePb8XFyZaYpzV4qeeJnlr3dDlfZ1Ny
i3o7lkMC8yTZ617N61J8ZEPU3RUnZM7wAqpkhlDd2wbjGX7fVHYtQNYlj3x3Ur1L
giJrzTHWTpR+D1q+C7StZN78/bSDBMZgSwZ2IMSXg4j+inL9tfhA0mObtMRh68EO
eUIPe3NgdClLwdN896g8Vsz22rFZgbdhEEwZ5bZwfJUmcOOaOeySZzuLFMUZY4W6
ohge5w3FWCuX/5WAghLw7819RBRzkd1TH42jaFpJ1qlYj0o8eTfiI39LMPg8xZC1
x/2GieCVZA/DNKFDPji50t2IMgr8y5hUhUYmOlalV8BwuUw1ywEhRmBSP3gErWHV
lF8nbwMsWI204LKaW6igtWpA/R1yInAUAd/v/nhUIbSdwZZy732W8DeYo4J1gweG
cwUWBxODZaDDRLyS5bOOEuDMXeqMlUNnIQpi87EBIwXJBqTohtSUk8siGr4R8NZj
dPUe/WrcLowRt9CEj+5rb2KvNKWtxfmnJpxbJ5Mhxbw3ETbJvyL+Su78IB2qYPfF
YtjRGgcSftDJlG1J9c7v3NX++LCa7OXawPphyUYAIU/0gTgzf7o5gfgkfa6Isi3+
X76Sab+BTTKHk8XOS594ddebDTSqDW13t6KNELyPoSetpa+5gAvFsWwafWFvbswt
BsDb3pfd/1eVaHTY/Pg4ba4tZ8RSs11+UEsm4mwZM6+SLRSIE2WUkhu4ZTSBv4ZT
YnwazSL+22Uh8va3ThZHqUpXvhnP3mDHmqfKQ/tMQQrJ1UToZVwvlIhqQ7GuyrPV
ECCA4DkAfSaWr+9T3Ej+7mrw+ED4+u36VLAHr2rhNIcfn+iyh/mH03F4fmMWX6q0
xblaqhPHXwNnA8JT/zpvJJjpQXXqOVsfL5xCOeXmTU7KTxoNh78T2m2Cafan024D
j6WcdgTyKrnWxuC5RgnfNe9rvS0MXTWISUgL+cBJ10O2o4f7Yc8gALxncmJTWLl/
FrDzT3TrGbDu857KQVovrNV/fe3tPHo6VZ9YiysR75Ym0sOtI9BvDM5DbvUelnmE
mRD/Kc5nEIsI16ZQ6Kv1mzc5BmqIaXGZ1mWajOo/bRCESa0kFXiz17+P6C01SpLi
hxgACij+a95uhhirrYeDrpusYGfB88nMF4pbnsFyZkM9RDyZUVMBqXrqqZaGOrYU
Gq8KlLSzHSHF/RQ9SWw1lbsXfdcik/IMVYW78StiyuPRruqsirM34vRadKFHkIGO
9Df9+wYgNa89gpYZ+UsTiHofIAiXqY/KyPWb1SxsIJKs78+6SofWiCKLqQ9I2/bN
dUPOVVYLghQzn52EpCD9O3hO/rzzr3ttd68M2EwO7SUIyihcfP0zSLNty4w+YDKM
6zCsXbQXn6f4Eg2oeNT3xEn+MjtIo9IWAjEJ+MyGLOQ/dN8DcqHo6ZWT8GNuB9CG
CqLXmKeetK4pSslBrtKKy3589d+m+12eF+BNMUJ8JYMJqH7wI28Z2RE+9uIGJB3y
pTnZ7eknb0pJ4AcQCAt3hCRPsuxF/m0QbWAV1k/AphHOxdbFIAghFqyDAdIpKUcz
/NFcR/O/qHmdfbfJvIYM2/+waYboFGR219uR7ggmofaR55kjrAh4uWQ2uwVaMrnw
3T3RrjrSoqC04RxozDXBTqXWm6wRCquwBrJ97jLQvJ6B1M/un1OOHbUZ1uRnyiRJ
p8UNBY9SvbEDhi0nA6SUOq6hU7aSCpLMAG57ZpUO9WawhzJkSp+UhpQFJoBKGO+y
gNLWpT09U2kYrSzufahaS/WqQDv3Q35lNgRZUNNUS8RIhk+Gfwk60/1hLUknqoH0
oXPZLVzgbEkTtRs/ucmrfI1XTF5/VWgUNQDQ7Pbf+Ylx3RZwKjHt6BwgdF2ao4SY
Pf0u/tDLe+zzmsnTP4+RnzoMJcQdbH1gPghHZLwLHfr8dG8suht9cK/NWJnfACJD
3stKFTaOoIHJW7WVkJnHgdnmj/fOPQz50Fy7/8dtcl5cawM5GCcAeksED2zGlRjt
J+0Vd2mfiRWxLXv6fPN2948rGuLbWsGnhlvPhL1qOBqt4OO4h5+o+jWxN+GVxE1b
nWgHTY60vm0cPbpdukHmgkkK+YK9Lp4aVkWcZHaRCge20PuMfcwFQye6uRGr3QyP
si5YvwQs9J7V4mGLu+XggiL1vITaUTPdQydbJvzGGn0Pp3YZ1Ph8dKSI9J5Id8PW
je+HELxN6hEty/iHIFjYa96NmIi94/cWVzMXSR2DvyXVEb/X+bzpcWlNuUWLG/Qc
FnxHtrBBEY+d9Qnd89ZN7sCOjHvdfnRXeLJQRnqYDUU1HHZtuJ16yzYvcgSu29ML
aBpC7GayP2ovcJqWHZh6rqDmkv+GFeDWl2lBp9TMf+dAP3BNrxLMjI/62M6z8t1n
yLZ5DkGA84sHlgi6hbp3U/mUv/mAY5lAwKOlpy+1daPVnotQdJzNGzH7zKK30HfG
F2rD6FC9GF10F4VoiJ99JJoyVTd+Brl7SdPRrCzHVU8OgSq7A7bGQWavktuV2GPB
u3CP8velf9rAP9AME1ZwCYOE5EUa0m/eW45Xu7aix3P+ERuRF7VFY5Qn0F2PjH10
HJxjiakQek1o2bgnKB5t5H1bH1IlG7RAUDTvw7Q7DqejW5go2K/zXtkVWTo9QDvK
N6mIp9sOnqVwJhkkBEVMCsqQKMHVWdZ8TDZO9Tfl50aTykj7Sh2OwpZYdzHD9IAh
3jFjBWLAbthQMy1mj331z1D52qq0ZAmEhMLB/siaBLotV0Z0x3UXtYmGoF9C9wg/
8RFsm0cFRwbPiXpEXjLuGK7etCJ0urwCKe1pS/FXxm5S7h9eBGpa+t8S7HwKayuF
4EGvwYVrDAr/ejReCLDL3UP3SSn09t4xTpu08Zm1nnYt8hFkIcNmDdxMmf834q17
tEUPzrekG4voPKG70GyhEH+hl59IFCwVhpLiJ8zA2CZaqVsHiDdxAtm0Clk16ntA
ufu3ec/xT40gn3tBJyP/Q1NOOhoI6y2CZWlcYvWJcSUdMTVlT2200yS+FstXuyS9
tlNXLEc7MzqXwwTightmCzamdh5ijMvkuQ8Wgn4MwsyYxsBPtyp/dfydhvqOaDNt
3njIh6TJzl7LH6/6nnOu9WPef/gmPwpF5SKNFp3/nb2fPtddRP4GCe+hT0tCp4oi
kHVv0Kdo9wqhQOdYr9vcAoTJiukQzNZuc4wkJKFgxghgSQVkgItcDIeU9/facCYI
YsHCJKEGBGdx2rGA4/4IeA+Vot4OEAIdJRztXg5XnhwKBL+Y/kOqQo8DY2zOUgN9
4JUBgs0hmwMrGY/MCU7msUPzZigDnhX7FMuPLCg9pPOo9Q+xbcw2EPzHx06YXp1h
L86dBr9hkkQ6E8AxX0Q4Re5SwDnBytPfaiZ/dqj2I3zTHDSzzU4gPX7gg8ptdXpQ
ngm1DRPRozcz7uY2Me0zJ5Tat+a2dbI0Ig6hN7fEKbCBDeZXcAeebGnAcNpj6qeH
HMF6f184jBG/HS4rsVcGUPoNFY/g9Po+JcXbeEUXKJ+1chxJ+y6KGLzKlZWM74wB
pDdNx0CU1qvLnbpkbN1+/g1/UZ8rocAaNGwEAVfO8ywwkli+tkl6UThMGsi8IILU
uk7KCMyyY1+vzzGtARx01Pr6KJ8XLsLyNDq+y9I9MzXRvLOCTXMPdUPdS9qONQsx
44PaLkRWAgcmatRjw2qrMR0SnhzgtMcvYqK1fjKBhOohFhke7Nq3w/toztpndaEm
gT0CuzBqMWcrv0RxKslb2BqNQceE38nPfdOjl3P29JSEIRPJr70DZfopRZXlTAi0
wSvt+6BbQMbQ93z13oushVU3VH/Vi9MEM2scUZV+YpKQQBQ83/iSijBRQiIFRfNl
70sFB5eKuAV9C5SRBJfs0joxcb917nY6i9iD7h6TKlbgVadXgIsk7kFaosM4sU6s
hjIntAiG4mqI5WIbCqg0yAb5WWUmVG9O8tg2jXcqrpKCguUG29uafgqwehEiJeJT
axg3A7fwxP41Q4rRRns+8U1z9PKEB7yhZWqEIzS0+PD3Un9bJpvZdcIwBc/jaFIr
w33Jxgml5f2mtI4potPpSvJ17IAoiz/QXOXIOI5vidT9mRKs+y1lpzqb7BQRNtIG
x5B7AIlobycvy/eBAS4KeAKnCNakidxat5gBPvA9lYUWsX1ZIgFWRttTi5MPIBIN
SyWMfEyT2zBfgErG4ayvmwRhdKje6Y+Bntk/jhyU8Xh+3Y0cNwKw8SKuV7fTs6jv
ImuWK1dfnfRocuBLLvlzJY17x4xLzvIE/alMsvBTpNocOnkiGz3W+6PNAVl7AP0N
WG4YxeyeD27r8HrqP87N86+pP+XXoypbt5X1/fh09+59/pbpMoCMzP1v3djR8wIS
5kPyjpVvev7YKonZ4hClmMhJp2+SXmxpvcCQAFCOFjElSCvLGoWR9T9XHoqAQi3i
XARcXjB7oLIsxG7UBMc0tckFzg6VOL6nOyBDYL7/rSwFcdZW++XdpJjNYnzVBG9P
7CgxwKD9LQnEazOmW5nrafd0qThhFy9Rh54rt+WvBV7QfmNczno0usaMSHl7SPql
V1gMVCQ51AD/kaN6SokKBASGkHzQMYGBCn21jSmC7Khued8a2/o0zaIGvtPSp0tB
sU1+/NyJjnQFm6PnHtNhUXlqarhU+M2/dPThAbozpocDsIyJiyO0duYfNr7a8nd9
bsqXZr0ECBBj1CznR/r8plupjIFpCNLX4pll9i7pKh2NjV0x6/1uUyDgH41RsUeG
4u/6yiGei8xt7RlVjYn5fpUlIeZAuuIpaGeDXIXyjeNU9oRdjMwgBrDoC9otOZBG
gQM72OdTcooGkVfKG8BdZBYQJLz7DVibqJzFYTcvxOB0zf3uWJUUmVDuPwtd8/HX
WDIHUHoxU0I22vYi/Ytyb2yK59guww/ikgq3lpuOt3k/B9W/Mqmdldde0lh+VJ/Y
DM8dao28NMcaGCvIv0c87M0TOCQIbge66lD+8PnsT7TXp6DFm8K3wZvshel1APcs
G0LeVGatJSWcOH9TzHSNGsWrXraNF6ZMC2WSRAKkaTzyNI7N9NUpLAme15NjZJFD
FrXqcV+MPQMM9OdV/jn2JuRVvD8/mAwE8MLd12nffuZMvClAu/C7JsWS0UOVT6p5
KaHzJhpwYzH59+/sfPLPdkwsW6Mr05sI1aMZUShpIiOWZOOEC6Y6fGnCV7LkAXyw
FzyHwnfN1akCvw1uX95Nf/5AsKfK2GuTi4w76XOyRdLMhBa+wYFHNcXBJlCjFoa2
YETRBF/qoLgnxVnE5OmebAsMIwHordDgG++MBkw/DpK5qRWosctGqn1Mfu3iZA21
7V9gQT9sOmLqBIfVdBYr50VQnFZcB6k+/Z0BjQ2+SfQfDTqP97KXzYKi27VaC/v7
KrIvZ2k28XglZxfjkB0sZ1KyfkqM6GzOK2slZmT/zTGtvfvAmyrP6MH6UuYgQOlD
4LTPEmbkf/kGPrf8BpjKGABR0bc/ecY4r9HPsb7wJWPiub6fIBjVmVhZAl9JiJiK
x70Q0BKnUsD84tHB6JaI/g6oRTwOgeezVrXM/suLdFFRDWJwEIB51AxjnCPIZcd1
IoQ+PvCvYWq2YnAEFuc6oUmn87J/cmPM6dYHaVlU4bAOI82n1R4ekD0t2sL26WTp
KIttWzDMKENR+TK8R44zm7W40+HG0BfU7NSw3z71iuN8bLIrYlzfI//oTE4fL5FD
dBuZfFnRBwYOndq7VqH9aqeDIx1SDZEdI8XuQQow/KR3uh02yUsxOet/gZmmXHJf
1Hf8JgBHXgmhrFbQRa/S0CDBTd8ad55pIWf+UGu98RUx+fRr9BdUUjsLcGCd4Gi2
inssv3BFnHSoKgw8G5yl2HVQ8D3yxD2BTX4LT91XKwftihb2Vkpz2SA9rGDAMzUo
B1dKJH27vQP92fc930qwAVgoGToP11QlPH9geJZuoC7NMRabf1AmMKdRdyWPU4Cj
jWd4dfxmsVd/PCqH0ON65TIvJc9j/NWUUI7T90QE0zDwdSJoVr2sNChaayQdWK1U
yhYcarKoOiqNPXwVBv3ZxKp3vnL6h7lIfDq2CIK5KWphp6h5XqYzvucz2s0Aw3sM
l/lcqZGPHhFrAqNggpmf6vfS3Vi4VlnDtdygV7gYSOb7q7i7+JvEJCaOe4w5keSW
zqF6fNd50pqTbzMIqbsmWtIMeC+jcFS9er3QnzFttVpVFJ/K+KiUEY3+L421dlhH
ajkbEUJniOZfwgk7hsoR31oY5+kGWmS1iCn9+D1VaIAUuqQbpsgOlZWjvC0axy6W
l8FFJyGJ2HfUWtjKMa8KcizEmsGdztWn51IWq/SBIlDTowx3mJu4K/PochbfJoZa
wBA5M8TvC8KeaTxrgf4N024v7Nj+dDOWECNkNn5YJicPSdsURtp+t4UnQDXe4N6N
W1yKUmAcYAfcq3S2AtrY1R5U95+vaDQDwEurFrsM1Vn6x3tVL2mkl6Q9YRqKADhe
/vkrpNP/t7f/q23CedsSFX+N4dqdYc0WC/rI9dW9wXHrXuN/W35lINodgNJ8pApt
0PoajehqZF+f73EwfIBI9Jz2ngVVoNZPaDSgTapzr83XLSI8EtcwfPMPxNpRiGww
xrV9f3EmCSGxoWpqqGuBuUeQNkR7ZZspnChm4DySXMIcAFk9oynCIDShkTuuzeEB
b3KPMmsCBTCHBcvmIZWiY6ovOXa7CSJcl8ElCogDPc/QlPlVJa6Jq0iY2/Soveca
QctsXuYAAc4HEnQv2De1U91Ug4jZ3QrrHBWSW+Ma/pBxONsO5KZkgPsgKM2vt8bX
UbXqZlmCqssRlus47UbbMkGWbyRdekork+mwuajKl/Vl3vNV8UTunGayg9yYo1c/
YkIujwhXpNd/mDSod8OozkA9g8uo6YcMGAtEgoM1C/3LWrrcdUMtwM8R8e9ytSaH
IntipAv3CCjAR1LHbqqNRhxilVL3HFW/Rum3oapne1uVIhChoQefPgetazoIstIy
zD8a+Rrpy4jpxmsJbyDux9naWcHmkP110oJCUct9BMYw1/LZpatqjyW+7dyaxZzL
qF0k5wDl6/3GZ+8pio1QJPbTFfghfB8ddLOaq4O0FIqckOu/R6s1fNog/bv+y2lB
/heCwk+3jzlINenj4lUL9D1jOAcqSQCVJjXfNKBb4KLCPRewviP/vPwrVefhnslG
++mp7zgRYXa6a9zJC6QCMmjf+tbnG3ooZn6xbknsNNPqeI7ZrCXFmsz7yPzVChxO
qwgR3m2m5q5bMCmHoSfh+7DRX1/6Aez4zs+9u6hW5fxnDji2rqMO2C6vqnGH8TUQ
F6JJs0eOmC1Oy2Tmad8jzlec2FoR/G28SGvUHWYGT74VnId6MkPsJF6Yo1QXMHex
x9ySlZDvwqhCOjip3m44+dHjEoD6Taeqx/p5mNXXc1ltlGi5kcDJwp3aS6Uhkngd
DrEqzIo2RupjXngwANrTG16yvjNTL4HR2MVYbJz5daUF+bU54krHbX77pbsYigMR
DABzYn3b7D88qB9sDJjQUMIxf3wbalIYwGWppFplVj9/3U+BCCRNa3lPyEjQU5SZ
Yth5CZ4K9b0OywsWEt+mCV1ENsL08E0HI2sPTT7AlnvjBSrqdowlKn4pE2Sl8Arn
eqF7wLYKZOILQXIpeFlM2NzLjZ9a5bVs8YyFzr9OV1lMu1HeQ1TJEYyUEjiPa437
0RQZcWbvB/KuPfI+Uj/Vjv5ztS7a2sv5tbbzwwtWzfXdta7KSHcaQ0oLTzetT5qW
M70c3j7RLUxjn/HKB+g4JlB7voyWdmXtm8ngxE23lap7FEUZkxqTBnhPO5lIh4+4
0IN9ULH8F73QjHiU8FRqjFLXoJL/np7uZKayf/CG7MsFZoqw1i+GLNw9JkCiu7uB
cxcy8oXUIhnoyAnim9E05lwJRPokOfc6r2Bog40xfDhK9ASQjztGqb8oE0imsMds
uqrAemM6dc1ToCxSuNTfVan26p5Ct5OtJmCFsPeQ3heJJMtPa4ijHrU7vt3ybwyh
0CpIkNQlxxF8LV6LQvmI0aTrPndYhDNryUz4dody1Tf56Kby1aHb3njPVQjoySkS
u9xkqDxNJ5dQTUVeczr7m+aC4rOyI9iA/oP+o9k00vfcMx3kSi2vLKU8CNwspGzg
X8KcSSKXoZrzRpyIyhviKGQSuSwsnBm+iYk/DTh3Ry9n7MIjfoT/JfLZPKaiPkKi
Gw18Ch0So3LGaWkQMWDbIUbD+3IDx4U9ySRIuFiyBhws0k8yQZkmG2KBo5lbxIep
AFjwySmWEwoAutZMgO7DO2yHYj9SZBwa3ShfJGjuVXLmJavEPyjXTEey4pVAjLUh
cDigbEay3v2LqHstMYb+4tOg/YfOdrz9phg85D5rYYcsK0PLitsdWI7qLe51Am6T
/xasBLGc61yJ/eRnu5ZsvCXBUZx9Fag23NorndU9Ajt9HIJ4dOlDhuA/nwFoHwPu
yoy/ZLPwo09x2qKG+Qnu4uixWAIJlb89i3oVMNeHZYaR3hI10PyFIvyE+e8YE+EV
EwyfQEeGBsah0lpDoHoSZlQOy86YZlVSk+ryGV8qIKgFvNhWi+IgogM8czTjUFQh
2hbUGLqwdY9YaHXEfiIL74VguJ4AdwuD0kLtFbsNnAkjM0wXGegPGsxw67Aj8yh9
MFRJ8vfpDoQb+jbIoK03OQCyglF80N2xHcY7PQr0Agn7Xjb3+BelaOlikhEXFYD+
HAfROGoBpQHeFg83+wJuJbAzahE6QzDK8Yy1JCxU9RMGXcyUy0pHhozgRsJ7EJzv
khi872vLAjWjW9/iaP4aMc3yfctVvRs/rnySiq0taJY+AP5QjhAHA+i+grSJ+2pX
BmJ4eG8MJf27sLMtYKu24d/xJUPAUcJVY642x+vobmZcK2Zvt7stjeYBz/2usvSg
m8o2eYgVlZjHlPC6p8i152rePb0v+Wa6iH1pCWP9JrFT/vsOKdYkqPwp4VDVLpVq
2pvBQUAs4Qq7fcDuFTQMuLFP6YOm7fIIodVmEJ580CjUg9nrpnnYjmYA+DWQAwFl
+eJPvi2AJzB6xYTDthxhEtweSJBA/oJ5pkWyeh9F3YNQ5h42MWzDdVdg6w2hZBOG
8/9X1+3I1Gtrw0/PTfQrBlgohACnOvZpGbUO2eyjtBCBa5BiR9M+Zvnz4dgAx6Ve
LyzREyJfmyqHMqjvdenjVn8sG3KjXLz9Wdy2QjkKlrFKLQ6eSJFXraoILdXd5sza
YOh6aKWUrIuFy5BbQXP29s23Mu68yWGQIko7+2qLPe0QASPLbU0E889EqYj8M68I
pQU9AkPrbmdp1HlCsCzfPbR5x/MKe9eUfIF+RGy6y6subZETX+uNBBM+Wkwc2mOO
G0QVlqN+ahB18dqNoiYhhmRRt4frHmD0SbA2COhj8NBpthcq7OZ2PmYb9HQnNCJg
o+uT2AlJ3rfFz1E+L0l9tG0ZqTKKOXXgo4ICCFAqn2Pan6KoWkC3KGofBiZCTTju
bOvhqbMbM7P2a9X5hRZbUzDxAu/bOQtM3MGV/oetIwYK0A8eoIyrFsUquF9O5NLY
V2RnWOBezBLd+ANEl8le+eZgaxKumESU2SFF+Lf6rO7n1scHH2RggU/1xEXi0IQ1
N7USKLjNJbK/EshQp6diXtje+ZlxBbTDY1tYqtEw2JeKgFSEhYZioHzb1Awpva9h
iPug6Dhbjcq08AvgxqYRFf/fW4dHx3gWlow69ST+U/Qeu/FlBnI3cNWVib2LpogK
zTPvl4NBVfnw+e9MNlmGJyTRIgFl6dDG1E2EzSVUbdbtXH9T9BKO/To5DcJnKZyi
z2AprvIn38WV5Lfa/fJ/fRVe63gTdzRpKMKpBt+zzY7/3km1bpyrjP5BySPoUPqL
XF+K3ZWbxCB6Wp+uPWEGxG2b7Zak2N+ZMgfXgNYKp6mIH9d7+211tiXPaTfndBrF
0+xjkpiXIHARrcpvTOjuY2RigOQwYpI1EpdhzJAkt4QGhfMF3UBXM+3ah9k7MDqg
jo+YBAePlibFFag8FuEH/XuUsdwJLTluYYFJ8Aavy6WGTZ08xCrcqJ8LPnSL+E7G
m4zlzjB6jxtx6okhD/MqiboqNwqGqWokQnLXDtXDj/mMjAJoY3ptm8Xt7ETiEOpS
JcZmVmXf7o/+L8LX1picMpJvit3GqrKgxcgtlKsvF9r/NhfteLj5yRAQtKJM2FFm
1ox7+Ut9CTqs0wloh+oSmNjK4H7ZCwg1bZ1Ewl033XJPu4deGisSIew8Hi/eKuru
v/spT+B58/aCB1xChLClmQxIrN2wVE29MwXQMDEudocfMQC6UfAK4yOd5zF+em6c
L9QM01PnkTZ5e4TgZv1b5fCbLUYEQOKfLkkh3e3Mwk0vHaoUqYZ0aavqREYr9EGa
4pXcXXe6xAeyXKN1Uuz+4KI9HG2KOtARNdtKrnj/4Ei548nMjh1Esj16OMF02GlW
VwmT6Fiz2O/jWwt5DjPLnjY73JxZEjMUEvA8h3/51T9P7zkONL7Y3PL5XhXsAwW8
1+oTfkcJf06FMBeveDndl1jLZA0HRLWGUI0in1hualXl+VApirH/vVIhHDBQecJu
X3aMfCjlmoSPylcSU6HJUe35iuNuF3cC3w1P7OW08g3PvB1pPdNr3LOnc1zUan6o
yqUDNg9G/KFcIx+f6fvvP9jUX4PD9rGCEqe3bQqxj1gqDf+kHZkzAnzgr9698UY+
e12dkxkvDw6hgKftkwjugvBnsIB0GUdXPKjqLgbA7pjSQPrZqDCE2npy4TtfO63C
m4vsZZT4NXgAvdivi6342kQItlyYZqHgEegKxy4xLPFStjw4VTcnzNJn0QOIz2Z6
mNbBWo/0HqdZsfMcmCtwJAbid9r/NDH//Ii8RHEZlJfp9xI4k+KnyblmdFyYSNe0
2GT/G6OpEl6aiP0ANdGOnBo9aAvgg7yqHLigqxknFjTHpKTy9Cb+DS2elMmO/AFj
SlmREmm/GqEtM34AmmDwVtdC4v8ekdOk78hHZC45AbZDvFCmOKtog2aOMWGVBlgF
OLBKabmrjNjb//O2HYHL+jRTQ5RG25d0Rqm9DtwxHxPLKKyp5vpddEm2zVOB8VoP
H9Sto6U5I8yttMnERm+s6nBi35U1/9lWKzkJNRd0SGW3LBYldRj0vzh2N6ukk4Ee
kXsceJ4/mjd1NenF2038CI4GEZZ5IqNrj0PTWaxpQuVlL/0rSN83j1k88qOeASyb
xjs1cKCGbHgGhM3w8rwaL1AygjP2AzVgMzN9PoE2B/+g1eOnu05pEjz+kYihJYd/
Os+0Yfb/4ajK8bUqmBgLL2QpoLR+YxoAhGt6UzdtafQTbs9JT2NN1Ft4hr7M4XA8
0eE0ARloER6SYoVGG3//wTTRH4kjVr67xlVJ46U0pFnT14eExFImnhhmOBSumvU9
m6m40Qx8Bm0Wfp/j66Ulq4nwyelfoGJxEbnG+mQxKMu0AV/FTrQ8u1d+Bi5Qqup1
ARN2leEjkJ41JNzLWxA5cZ21uOMC0Cqj1YkDGSqAltKBKBvqKK3fBoBEvOC8M20z
LfDMCt5ngP+RjzPsT7dp83iGeLtSP5HRrAdFf+V4K4upkLAKTGkM0ajVvbbr/wIq
uRMAhjGjl6w4cXqL/5jDLGEojLYqf90xQaE6nHIl6s3G8nngvyPvnbZ05alG/UI1
6u9ineb5CRjOEdsui99fYXbDQQjwi/RCRWQt9gtV937TYMDmnm6LHfCogJ2FOOKK
c+Fh07hAxqZAhPX7KcBu8HeeNISCI/BmjkD6A8nufdGzOpuOWnjVyd9s/zUBCM9c
l3DrbX+dU8N7NX8uW9MUUb7yoPGFasuVEtRHrPhLnNaQUj+qe2sXnPTiVlJ+z5bo
mklYDijAtZ9nFwt5EI8KMXvw0Ge3l8D5bHkHNAwp6QGzh8Tpd6CwadO6/UrO5/Ux
BpjtmdVew1jMVfdZkm+2yck/QVQh+2eOmsAxjSRBOoOocFTvE+D6O6KI5YW6EdYx
/Qm1dAVi+WB7+uJ5SZLWKST4GphdVu7E/saDjPgAykND9/2MHKnllGxv7Hr02LHo
yCQRpE7KRcLxQ2RgiXNVTV4Umrrtxh4ASFBkd1vK+5XJDMqtNhhYuXifeKTF3OdE
B1utf0gMbOADVMHnDlcloXGSzZ8C8up6yFfLWQYP/YdjHL7KByU53nY0Qi805RcP
ONHJfeupfCB3tYh8RpUjrtL0pQOLoDVH0ooZKggu9hZknh5JeMTZOGPNul81OZUV
jmdUljnl87SjOmMmSkLao+h7/mIBHqC5wJ4Xq2k3r1yqDrdh0upCNTf65shV1qwo
pV2AVyoOu1gYObC5xFWkWvyV1/NEmypWmUzQvf3YvgPrP1VMCKE8Qw+4W9EIwI79
qrCKM4hvmZkGXGOZEH+Fsg1iNMeoCFxS8grToI/i+SUomkhVClBEQ2I4HB69GFUM
B/uhLJNq9Ryj5X0Wcu8rf/hUmb7ZdVgCHT+g59nFnuMSJL/BsjomryNFWA6PRqfI
LTrBvXi6hh225NgUigPouFY5yKvLVSYqULo9XXC1aGCiii8RNDQi/RN0GwgxLYQV
QKzBDyUP5r9BnNqQgill3OOTk8F652yC088vZnzbR2OIySpPqhjAChn5wOFQdriJ
avxK85cnx21nHMTWLqC/6f7jabRUgtNuo5CglRuZH6yBdOoPHQ2cMVRkqD/vRoGM
wTP1YmuE0Zhx7R3azDAN+TWzwhCTEoxHvXYETFHpfVNOU2BszlYa1nV8UEmlnijo
/wqBBa/7ay24qbX6wxg9fWbDID0Zc3yb/reS9wljmFWictXrehoSEsthzXey8KKA
Ln4Il2L7JaqITf19qb7JoMwlKuh/H5cxehrl0P1S/D0k93Jpr5gggg0g24qx/Ns8
tQCaaGm97/ETAK3CtqEk6DLHV8jtMN8MoW4m3fJ+GhTUZMfrrla8pMIFcD8O79Eg
VgJ7qNnkeNnfufQrF2mona08ahA9LTmAdiXdB2hDAMQM8ITUYp5ZftOOiinzGV8Y
W1eQvhsi8rarYYu3825EN2Lf1OQaFY4CHF+DRZK7AMKUl0Dj0l3CkeQoHVpAkwzz
yIDOrCCu4ci5czvk8JAyU2ct9UaxQTDkyXWolxwewOM4IpiNqrHx8EXr0z+858kB
SOdoxLMrBZx2xLXP4IvdP2zhNgEWFRngSa6kbOmJXKINbh94BcpBfAyAGB5kx5eY
0po73LQ8k5OjMyJEl4XsCB+pbOkC0jFi88k1jnAJI9fUcIj+9Gn9Ab/8ZxuH+yyd
zipDGzP6YTbBMmjTp5648w86x1WW3NTbm7g9+xFrdsh26P9VDLKcfTasNqcEyFlK
3x31k1VPr3qfvslRhGNbjg4+1L8q+F7ZG0Q0Udegrg+nxkb5536l9AZ8CU5WuLW1
lG2Xx3tmzZxGteNMRmuerwsvd6hb1oaTZyLBDEcgMcQpvI9nvl1XK7mQBVRxkU7g
lV26qQZNTDZFFQKW82PNPBTCa60lyA3SP79eBa2V5wBCW0vobzVCANft9ivJZozE
7EYpsj71Jw2aYFHx353hOSnkz9r3tfc0OQCcIUfvJ5XhNVNnVjYQ+zYP9jL8be55
xxWl6EdepE0GtcND8r6NmBwREsP0EfdgA3jFh/IlMN6tc6WO7OnCzJpObcgzXv5Y
zlvQyk9ooi/AkqTyXAL4NBpmAsKcdUnZTyCGq8UxyPN4/PAOOm61NJgZty6T5IPi
x4DUpxLiBXLHShwhvvjFhb3aNKS3PpvgjUutN3twAhXD7B+cOtTcYEeByASXX51g
EKQ9+ZO/vuJkFqxd1t955OFfcUw+r+aizHIu/jQXl4rGwtxTuKf4QBe5uAk0Mtwp
Z3kH3gtAzmbbPeFDGBr5AkHRQQVSrwqISZuVbEAadP0/QEdtS5cQHpIFX3pvRkxN
yJvaocfKgYrmiBYwvXfQ13T+W9WWl1Kr12w73475hQ3fOK/9aJ4PN2TWo6gS6Tm1
3EYakZW3Prhnp5c+q2YI0Hi2rfg+se2uhxkYSg+BayPBkUZf+bphsfNmC3gzaYfi
1jJreW97Qj0nrmAupz6nnbbfAuyKZwQ8sO3y9tP0L3bktyBc1MYN+V0cpycTm//L
+/SX7zhMkQkiA1SPNSybKKE6nP+dAQKyWhVQ0c5IQfNcnO1X+3DY5+M/n3AO91sb
oZBPONz3aPHS5+9wGEW5mzAUJbQXE+N6b08e0sI976+7bDeuhhZt/z1xf4qR2Efi
WnjE6GUlMD4tvwkkr0bML6YcdYMPpGjqUL4Z+u0Qjd4YnkrcuqZvd2g7NrbuTw1e
UEo0pKr3DNuJ1Ex9dO4bWtDL4OIMbHWuADrMQkwpM5okzazpWBWzBnE+a0PjUwBr
QoQIlYhJVjBV+JY42im0Gtzu29xHeglif24X/cnFK8rtKMuGgOXCPVbq+FuLP6Fu
5JowwpA937FtuOQfpCpKPAApKrKSqQ/RbAOEER//mGVcl6ZNS2ro8lB3T+DSl15V
HlNMxDlt5Lrefxi55aVlOll9Z3eZFAQiztIAEME/Y2OThi5nyiM4d9kDbpiJAEZ5
BX58z6fs24UAQG3esv4QDP0rXvCtXZ0euRluZ1hIfv6KyO6QZhdk8rXMnE0F+uIc
uHxcu0LZmpwzlPz2+2n4xXilbcmuXTCkTIEEIfZ61i7XKaR+b4/87qLlQToLXUhf
DQyk1HbJtLOlFKaXdxw/xWaVZHLq1NPYAJj/J5SlT+lC2Jb+p3q/a9XjdVKRpQVF
DcBN8Z70DM/eg2kAqOQp2YlhHh3esviRcy8HbTH1zvZZoVVHwgqXAc/8DFLOIwqe
Ch0NC7AdJ8UUgnSpewVSvqdr6WNXBUA6la3cfEUiBwCq2rh/t5z7j5Ifu+1tkyTx
O9MMLoH21MRV+xV17Z41Eqq6rDNJbvRLyxGGx5qKfr1iJdS3Q7aE3PaWMvajUW/m
XWXOzuiLF5Lmxq8OHVQNP8tOZ1GG5DqzAdgxHZR7M5QqvJjt7D0kOPRLg9D/Au+h
YVHd/DhRk6lrVXrTEYHrFl1gB0Bgq3gAiXqM6A2U4l5sxzgxoUk50CT1VVZAlEZh
KhAzkeam+ldOcU3NccRUxgLdyobBTyM/TSWdoq6pi8fJrNESls1Ky1hsivEKE1b8
DmKYsJSCN6jkqJMGQNTOObdnz+puGtq0k9DXr1GGx7FppA1C5wig94COSUXj1KTr
B8NsNY58NJRPmIpnltL+DFLR4q88QYKuHdlgU1yuetoM/2i177WE2vw4XMwM5fBi
eAuSTUaI7AamAo0O0yWy3YlApNr3/3xvixgXCGJJv8IJ7U0kHqgLfwAONJO3nHmn
QztlZVOJayEgUD6cYzdMKrz6J3vaeGqfVkAYBhKEpwGhd6++JJs6pCOMAT/xrX9i
hKt13IsVx2byTeCqKCbzgBqZEbl4Nsp57yv78MHOgxS7hzJDK50gVbyOliWm0LkL
bsBKXTGmtVEW+mam62AzvO+5TFxQNlnsToxftVVin1lWciyzlLwt44aIJnos52Xr
mFygaLLM3QB6VXAtYHEDt1PRlwL0v7XW1MiuP041xp1qAD7eLaLZmBRNLZesNgCv
yV5PLguxWxaawr/go5PEo+ODfvux3O3y9UkjJgN2MLWZTBtBYu0GM5vEoBlzaIoK
dXSKSGhf4rG18BUGx1t9mgcwmK968tK4mCdkwuVfWdjSNc2SoMVIhiexW9lWn8+K
ZZI9uVXOQ4YpcTJ3EUHzD/QziUKg4KZsJPKyCAYTVo/lJpbPFSkNl50rkQi2tYPr
xgw1ixytJhdQO6SRnHP5girocyWytNaV6ocXbHAuVG/11Qw6IIKEw48uVxGreBWv
vJ7IOC2edwQRo/YHBQ4KpjnbsNn5Kctow0+oxNReczu2HAZP0VDsrwk679/vVC28
ipMxGvrZyFZ4NK/OLNyRwQdPPQEJ/b6QP3WJtM1BgnZvrQzzqExGVpTa3nEI8svp
Z2ADwcLSF05gO7JTEdPZiAz5om+9M5EblfoArapu5XIOLn75oqZG6EQSdnom1JbC
3n0mZV4zzO+HwEMMfnAAp0wvTvb5GrjL48jIWtfGo7ulirEMrKTt7WdtiNE6xvsR
nD6nCxV8gG5IgzLpC48k3Hf+wANRNg7sAn15TDARVNEnGMlRkP9EGTzk9/vnb4jO
rSQVa1OSFoGzxEFyHZPwIH1R5pBgE/XhNKVFZ0fcfHFpdhJcK+zkhciq34cgDOSG
p3JqTLp2U2ESsZZ9ERFPejBFsJ5K3YT/9UNK2Icwh4xoYOW1++Y3MwymQPcVJbMm
gEM3Eyzh1RYmjuXhYY8XvIOpRNNn23dwAI11/7WWlUqfVhAZsPiF1wjXz2OEXfln
mTQlyNvwvbclmaYPcEHBLMH89mgvtivV7+mnzUGh8mCMS8FHqIvUslidBO8/ekAC
U3zARYs1Rufkwd8fEzxYUa7PFf56bnRTUGVwHPqGwtWJKmMUclPyPcK/ID41xQd8
SKouRStxso29EWc4I175aYwzCtAWV7xcNBYuzKKAxKvfJGs1exNWexvLAHUpicfy
KJbReVYEqbkE5iqOG0o1/FqxLgSrkl8MURzTW7u4ALEPTPYThVqmOt/RLQBv6Wpm
1Gulv6NH7psHwas9mAVgWbJBzImblCsVsGIS8ZCn7gzJjcV5t2aptrrbQZHmqfdj
zispo97mgkRjCi9qcvMUVTLpa4/rgTy1Oo+qjnEdBnkKBAjaBJOFxGwm59NPC5a6
+pB70UxK7IpBCIWAD6ln1S7SvxogNp0GwERScG0FJOBdgzNCkXjfvvuRC+G7fJpZ
1WEP+afOHfEpqCiKFjvcYuLHhcz5prFLz0qiTdHZqAsJZbHq+9ABlU8/IiMuKJj9
qOCEHu1e75JQxHtnQic2qZ65aiwk/6tGldC2wFXXRdbBA9aUa0t93Jlmr5O0Yk/t
q0GLtQTVMjhYxY1QNyZka8utpoOx6k7Jfj7D4BUkuoonqRHbcMscJsUzVbo+UMG7
ZHzQAE+32GFSvlpumDxsDbzESJnsyf7Y/PQCZJilXNLWgiJpxfTVzwJiO2A5lk1V
iX5Tj88htVgwXxeUA1Bbqv2SRWMRYrs421VAsWXqqBDxyVye4u5ZpyC45+4WBoje
wXr47daFCfsfiCATjV4CbIOoxD78pIGSav4aK1/aM+c1e8Z6ClUxo2F2gXguMfaJ
lVuVN0jjNeSuI/1o8hbiZjsu5TsPiiCyNqklDJV5pb/GFqy+k3D81kCAJTt+MzYw
1wIJ9HhMxy42/go/S7JS1f7zvCttCepCf326M81DuCHLraALWULxajObvHxdmXPN
i0/U1l0syhxIsI/AQX8/edbl51Zy5J066J79U2DRLB7NAVWNW0E8dI4kRKEfE9bn
XKxh2e2RbyxZLvVLgeVNabrjEmsp3fKPgNZ7FGIYm58/hzOt4/fu+mQjzlQWwbWz
jXvyQd5frAyW2YjRJib6XP6uENhT3hi+UpsG8GUaej9m/d8IzmiKsCvPQ0PSZlE2
4gX42D40Z/DDLSoKQKwzLcCkyOLh/fXcgvgsrVEmXUAtb3ntZImvVtPHuC2Uooea
zKaUU4uIIB2hqS7ySdUl4q6MsToqh9r6Mqtx473c2+MSDHi+brBSVdnzlZ5CNcqO
inJrJ0uTA9qWG/ld78bepuK8fagWyWlu+WPfcA8/ulRzjpxZbSCQBgMKNz4wyenW
6ONo309iIL19fp517QlBkBPB+QdXawlTIeOlcZD6pf02Vq1g4SLQhsf/tJaruwbB
X3e/3KThylqEeHuzxdCygANayu+I5vkvNrCio89nm4tNe51Y6rgm9CvBSFaiq6d1
AtBZmWr+pmB+jbO5EakmPj0Tu1ZmMqnHUISut8fGVZXtY1np2333xQP5wm1W8lNf
x9B09yJYn4vnnWu3kFrOnEBS80tzHFvMljVJg+I2VNN7SN06G6+UmJekknDqJnjG
qx1ZoeOz9gpBXXb6FDYkVmgg3GlEjEXoCluWZu+WPO6k81gIALRMh4hfaB8+DIBn
aeSDbUOwaXQqOeHSdLjvOemm7j10mQBH7hNytjqUc3Zww3rdkyBCxqYjt71yxDjZ
QmDb4SYGgLW/1+CbC7LSEabhuebi6Y8KEOThepdj7t7f2gA7l6/Pt56RSDG47P70
yb6kD1pEBdZEAXQ1Y9vHkg3QeJXwhChrjMfu5JtQTWl4DWSFCJKLmtCJpTfuNICl
7eiIpx7mTa89VzVH1mVJSHYz4+JOSRhOYTPNsRbLNP/8f450u6kK1Is+BoC8nvCy
bR1IsAYyoiWq+3XZhj7+Ga0T2Uf+bYLE0ks2qLsNEgi7tlWWjuZjf+wuxiT5AsXz
bFWnVIop7hSd8JFQwT82AD0yXZ8Y7kiDQusN2zrbcxNm2TcBymjCBUnx/At8XFQP
6AxlVZIbADoRR+OM/P+YrLPFRtCiak288im0p6UsOOTNs785ROppAfFymLlUrA2t
3cP3wndOdKwA7kmUBJo5I53zOPyW+qOdj4XVCR/4QJq+MzCEKwkwqJJPBHosmWdc
XOgKg/kvjql2PfV5NVb/Wgmd78/QioqQK7488E+tS3qBbdth2twrfKi4c8CiPmjF
r+F4R6/vwwyQi2s2FBHjzbGkUDncMEtUG38eQTmoaoiwQQlP8/6QF2VRPcwG09Qf
fxKAZqSXl+28C9N4KOqGOmRmqyLD0oNwLemQk+sAuJ94+JNAIkMamRYh+Dk6Mt/+
ZGOeq3p2Rk8GPW26rLVsQPN7hwcpKZRgJFlooqfqIAHAQY5IQvn7Y9I4W7OzXWvE
qKMx//DUdZOfcjgrd8NLfcUrdywbQM1Xc0OmPsfu94hfTXYL4jn/cxJYhET3Crq3
IaeTZxj+koCxuKDqI9bo79FAAAyUvGtZ5Tg89yYMarR0w5QP5XQ77FD4E89AApzm
z1YZgVgu830WzNmAYBAWzD8oXTjr8WPbPVa4+ijIaOgv1rM4Uiubb/2759EI+aG3
faAd9Mk7qFWuq4vsW/dHoWza+C5+uuGFQ87LYxdIJy0ToHGqcZOXdELjPYl1apuN
zOIt7Rc2U/fjlHJdm106V3TDFLRaEo9bg9X1N1sT9doAymhQObGOD/oLNaL+YeF8
M2PsBaZG8QhEUtFYyohMh4UtfUA8WizyS2okBqVWXNgLGciHgP4+F0Rt1s5rI2Ar
U8YSA1q3/ZtQ1lFg8ddX/zCsHBzaJIH7NI/MCz2q7ySIcGxAi8lOWX09+Zp6ScZY
ybC1B7U8ZiG9SeK+NfH0ypRUqm/OOW7T0GFjCVVlKA3a7RVqm9liuYE+ZrMjfCFi
Q4S01XMhV1qLIfKrTuaaeRXE6gDhHFLlo7hvkDzfPZOsLQiNe7X2yitROv11sEvK
eos6pn8m5gVJai96ol5jG+u6d65j7aL80e5lqH7tyv/KQZCel9O2F9LN4uvTkZNP
tOEwnlDTvmnHG5CfpHdbto7exFYuaDMvwsz7y5vOc5GNCKAB1TlY4V92ZcOutLwJ
e+5ZEOrzR5FSiGW7rPLoAKxgkVNqvN4yV+go8uXsLXC4Sa/GJVA+6Lr+l3lLE4Pc
Yr++jV7gQ1qATzzXyYxBrxTWiMSP1R9ihTqMKHEbHklUHHkQyX7d/bjhis7FpjRR
oPMqAc8xCef+6K2grugO7S0m3+GTmSqvoe4yNKIv11xlkR6B+x8I2iOQJ4NS6Ymz
6hKHc6cAEg+puwVd+pq80u5Or5F+dhePLIJzt8xj3BFdsUJvIvfTL36S+0TDwVgF
Hg/0bSYpsdY9nKrf7OUmjMfNHFjvJFOu9I+Barp6PZy6ckLOOk7OybEBCTT6r/0B
xqYat1PZrykvQ3MN9j1pGh2Ew08dyWwy6j5ZdJPTPS3z6gdGT+cpZVYOU488Cugz
faklpeN3DCoGNr9GZPVd1bM6vNuXSf1pkPdMlc+1n3XggxyXldujUYz595SXo/z2
UJkV94tqYfkHu3ur4PHZnb+IQ137OqLkYKejhP6y7drEB2cj24ySBoBfjiSX4q22
0nREg6Dx5R94h11H7mEhOe4ZktbGYg+IpilwVK/Y34EzY0DBt09p9mWiEPmIQIpo
YbgUQ/ZpdbNPLo/vLOBYL/GR4u4wBY9Ssrjs05Bkoaqw5d5S+gQg3AXs15suj3HJ
b5qxHAgBNuGspJkf7GU7CaljE550WWhcYlrFwtEMECg7NzFPcK1oi1HTJc/72yT3
AQkJPXhA0De7eQO0WHzAt4uOZGBmRM3/KsX0ingibmqGj/w2sFlkFGUUjxfJrrPd
mzn5cjmVVTJnkJyMaExg0SHCVHTi7yKTRrGl7x5K+imUxF+UaRb16dnNr4qlZngq
qfLIA6OCFjsh9KGeW4qBWJTGA9WbS6u4np9IJfJgiFw62ZBgn1BCbR8NXr4IDtIN
34YAfjUDazjKvcI+tvRxP1Ofr2LKHLXmGuDeE2TDYeQbQ7f3KDDNEkPXwI8GQsZQ
WNt8dbvZbXap7SddESRBOr6Vv8REaudd7K8OSO1pz1PBv2nf8xAn8/iKsEyPUA98
IO23oxQTPdwB5CvGUdJs3bvElcpEHhtbOcp8HTlxDiGYDXivplG7xeb6qX33clHs
e0ujm1RwbFfoX18K8OV33spVbHnl7qmhyBUEXOlLf4xvbz/UPgs1YngGQZrdIM3d
ib+UJSn5suS1eW41Ut3XPKgOTY3HrD6NvIt53sAqUMI4WhfT65XUU/zoRGE7pMbW
Tkr9sNTFL74rjpWJBCp9BmwWHp2ccBfYwzD4hzEGfqQ3TfsTKkSbK4ej273anm7W
kmD8C4fjIRcqP46ssktcPVkkxIfbD+OoDto6r+5VFYW55FjNh0t4wcMoIaUVXb5Y
onYCy7CSjXKIl8kr6uINIfwJ2fM34WnX7NtXc3jE0mm1yuGafn5rAhSuCflPa/ds
+WdJC4Yj47UfRDKhpVy4CCNr4UClI3h0g1/XbVilFFNfUOkoJUgYI6DhR+rVYIte
ADUFQXbgTKIqPTjG52g92Zb+X78WZ/t/+4f+LFIcJi23LENkU7zT7f9jYXIAMXjR
8DJoKDDVCYswsLB8sA72ehYFpBAoPPiz5vTAVf5Lv0m21rX/3J++W8b8P3Ur4tXw
qwiwHVhpdD8YHZ4UrxYc0aYEw+3b0AbB0z31DNH/kwGcrsC9dvCjQ591bmU0Eoqt
XjsnCtecUeafVvHYWUXw3ru1OeaCGiauuH8Re4LGzZFk295AqMFZXISt2lyz5f5Q
9IgAjqqoMZeJK2X9ZjoPx+WEM8yBTvMqw+t+GcJhgQjkUotXhaC3208HE6KU1pcs
JsL8dCbXS3HonyLvD5iSkJt8hgmVbyNeLkp5Au01s4vqmUEJeh5jzbMBofL2ufcC
sGvOs+fqO4fvtlxtl6cRLoBea/b3SlSXdTeFkikMIuCw769Aoe3/ArHSYcnfNG2b
Qt9Dy1I6aNgz/dAA3cJIzec7WRYtZN87+BY/cTgK6pm06ISkxIbZqsyOE1gJrBSK
Bb7JoYhLh28aVi+j4s+qfMo53dcDUHRllbP/1ftzZq5lcSXkGlZxztd+dykgDtWu
B/81LObSBNSfFE2yz+RjQr0hRloodZlQfXjpmWy1EgLzSaTpbuc7/8waW/xVGvHo
iFLuZEllcr/ZVumMGzA5HTFXtCPp+6EqyGwFPAjor1KPxgTbjo6ZtDozvFbdAVig
8PXkXeufw311cJva5EQSlKtxY/4AIqYJk/Em7BGzu7G9klCskVGgSRypT7owLTmY
Fy+eS84sYHIJLQ050Hv32CFCczsW8hgc0jaThbI9HcbNEgw+q0qpBNZDB0cFk3E6
Rd9XxVPlH1am2eoyHEoG32oi5LyrRFny/x5B+SjB1HwJSKfcmav0YiEQGmViVOBl
b58TY0IDYN5PX125ryaeTYxs57p2aLTXQeblAuNShdb4pgXE0rddiRK3Wj98Bo7d
PlTtfHXPiNbj6S70NiPRR1LqlAeyNFU+G3thrbOgBJqUjJHXSImr6jqJbHOKraDw
x8gJKTIgo/C2BlnlKfPzLKEftLoIQ3fu02sDcTGNh+p93W69jT0cREi+DywZ5gYd
R6uhQXgzhP9JL1r9tz7SC0w5fxdnRGicTAs/zOki2RSmn+SyfAuI7PzPRzbUM3F3
CHZQjKFhiXqM8ePPWxTYXUyp4py+KG/K7Ng5F3U2naJJPwEPNypMXHkJcDd18QNl
BG1auQOMt+UnI4wKXtZYtEkMgmm5bdxcow7g8CjKk/yhPYC47BTYgCb8Ha7HOD29
6A9ckfsT5QxGsSouEQFpyKB1D+doH5JqFKIYVkaeA8RmxeGB1EHiti4t4Jt5wzqk
luYnztsavBYIpXFqS0dL+aXARXtBpNsZz7aB7gEW0Ahq/JwbyvhcU7dx3TtM4i8l
azIUradzae7cZrTDYs0w5fCnvtpfxS8wg8JMhyJ5ywNXCfHRWal65YxIwu800K/J
wCAHv2AtxNpes2BBOA2NC5T+/R/VYbmC1XKwlCaVBskIyb5uxH5Pc6oJyY249pYU
UtL44S0Q5b/3Uyu0JMX2hlIF4nq+cXvN6o2TLJ3ykMsU6Z6vGryo5ExiO4qmhJj2
cTwbG3BrykQJU7xcGbnBf37AquZVF8nEvjkBJGrIHQfLKlUsIFDkIp3mp9fS8zmi
WNwSpMX9W4d8mCtfeQdmfDTAER9zjSwZWMqrF+Y2zc3l+gjtLuMDbV8+yuPsd3U/
5oHmTAbOU6Ym9wAMyY4W5dgj51eU5xhsKQ6i0auTzoHAmY4DkDrFcKm67i/94BZh
iOCZxusvyLnpB/icldZM0VAmT6PwIRtLgPrSuBq/ehu8chQN+D9GpngAa27LDtOf
O8muplzT+j7NEVgcYx0wskwv/Ea5dmq/ZcYYXnD+MU0qy8uwkXcBtvkE4YLyTzhS
iWkhNIjBrP4hT8QHUFe/O+wGK4ZQfnkzae0S5jqjA4s87pa6OyJmz9iAVZ+y8/1r
1or+4o5/p7NG+HhVYsmtEkdad46zkThS6nJSvrVd4oTcFOiSJml7AUqEl5S43ck9
CT0NN5/MZpxSNPQrfoBlZ0+PbngeqLnsmnxKGY3G3ftVRpd13tewk9NvZsvktXkq
07Gj5l/2t+eaKIzgCydKQAh8DshcK2Sbg0aCKlfffWlcZtzVaoIQWPAyw0/ptGF4
VfRDa6m1Rlrip15xeS7QFsebgwjZnJvEqoImnb7e9cnLEOEKZX+yNA3lzkn/WU39
dMrcq0lgXgmtu6Gbi90qeitcywk24aE8xxJi4q7GOe/InKfdE/oplMEcPHPWCBQU
DJnrvHa39y92ZCfr+lliDFVNp3Q2R0D5UUHEPjESqdSGDUp9Pa0L+SIAGUnR+VXD
lF/C50tkSqKdui1a/cwBorTXp7jhC162nB7XEm75e+Pl4zoFHcCldj1i1bZetUIC
L97u9XjX4Tfy5qJdjJcDS7G10mVPP4o4YyKmvuj3VcGE6sUAxxTZG+RaBLjPzuZ0
emfNN17rhr7Vwr5v9vYRUdTRF1bhDfue+tR+Zs2Nu9IHqjGQ7DW9SF4p+LTBJ8yt
Mh3cdOUKlA7yy3fQL4uUYDZm03z9pTzF1lOu3Kg822zwG5L4BxEtI4ZHr1A9X2qj
HCTfs+pP57m4wJNzDbZsQeY3ak4xLIMe36aJ0i4Y1fA54LtSU+mWqCpaH/+PRXlZ
fk9i4mLPOexEYPynaFmHvsw69+ogN/fxNaOJVDyUjvKhRKEtAAOjMQN5AmtU01ge
UPSN1454jZpmy6DGKH+T5OoImvbWgtduyhfoogyWzTZ1ThOwux3sZsdznm3Q6DFp
UOOUhWMaOXzKfKOEvgJjWinkraGJ8Z0Q7FlZ3EGJ5EMWqp6gQUodbtQlLOT2ndZd
U2ss26Kk5ixnBOLDWS64O+oL4BXv7hWsXlGWfXLtmE/tJ7sfqpuAE1GOXE+ksNRc
uCyDnEVlbtUVUGuJjfn7mNhk6StS4aGwM2mZm3tFKmReH6kT0ZNfuKlKxnkKvo5R
v3jY7NkFDeDPitApXTkKkUTZQAvmILBDABcqbzZij4FKOXvv8svjQl8GxytPNtqJ
DeRnuJume6JOU7I4kROTIAWexvx2yFh34AI+7+ZhENPrs2T6hCgAq266p3Iy39pi
t5OdsF1BSe+FMY+G8GGm7VLUoEN9s1U3SY/N0Fd+RD4eeKUkEUuMWqy6UZjHlOBc
4f1YZV5ws7Mg5eklq9yoHkNOrYAi1Sf9AxWB6uq7lptQPoDiH0WDwCZ4SOwDPJt/
k0HmuEG5xL8/9pV/geft9EtvWY1KisjWrOR0GIJtS3yZqyxRQ5VHPG7fmg+F5BEZ
ILvGAIzVnkXploUSPl2cl2k91jWUPEteOu/WFINwoRCjGhu85wHCfIo5Vu6BAHcb
6yyL+z1kEsvJYnzrGs8hgxK+cPOittIdbAlr2FKGBr2+QuPLPffyUfcBb877OC4K
bHXQdBVSW1bgdrYKdmqR3sx1cXrPGpTqQGixtXPWVvD7RhYXoeLSA5MgEkMvWVWy
2saKYC5M2zDnAW2rz68BXHvDBrQe3N2MVP4SzCfa4o0TLqig9+cSMVtP9fwYeoFU
ZYkvwCH4URpxAiaCA4Lxjk8R1QWk5aCAnzyuPqVXlgYCCI6oKkfFbnA2dH8bV0X/
2mRbB+jlWHQHsr8b5E/GPACId1w9Jd1dFi7PRcbDygFBoL0kQEolr9pwFGzBf6rO
6w/XIXSzJCcB2U+LzCFfJgHxZucrPg2eDgVbHgMRC1FinigAsbd3mgnmZh50HRPF
y6amYsycOyxm4D8bIpAPJTXF1GRIo2cb2b19tOvL2uvzb6IIkMN9RB/ZmDma0mK3
78v7+key1zia7FQDwHiTzft8bWCBKbCNXOHB/ZzBYGzn0qnuk2P4tCqWJQ4UuZii
tASRenSZvr5dGiTK93sf76+kDQ4C1YOvxfDU4/WsIU614C6NJpTWwEG/qHww4cAL
2BBvqUDov0WkDyi953txkltwYLFOaiQQDa5uVdX0ayIkdMIWGfLj7y/eoZd9v6Uk
mWZGA8wrRWhg0yLYoZuuf5iD9m9J5p4UtS+Ve4aV/U/UN4tLsrXp2eluf4Exxz1e
Zia2u3GpWkwPgmUzj2wCIQ59u8E9aaoJpFYQ+rTNIwwWXtKOhL8Sa46PWsnBcM9Y
eX6Y/7EzfE3Y3tmZOIp/BoJCZLsfAOynMPJivzCn+f27JAJS8vOBJAh3PPE/e8IY
+hwiDldmPiKlw3ci2EQ39QL9iVEZYj24GCuKfSDFiLPJ3V9FVvWGnLi2YEzj91AO
vwavx4ls02JdIFbWC+mn0kI05LGOJU2tqyZCKP5JIv2hBZj9/FoyPTvmIAKzmKUA
OHI/ONJtXXK1mErTaHs6z/OHNDoI8+g0+KZ6CqUOgQsfPOnOVyIjj2KPKVriSxHD
y8n2CoxOQZzMmbPr9HJf5j54b+iJdsEJay89916sdga+zuEhhGK4nVCbdmy+Pzy9
V8VV/h4E4dAt0gNNMgrhLLsk5qOE8idEMev1ROvNYZel1lGyELmqIy3ngESDtGbC
RkgvaydUCWPzGQeP5Fyf9hssbeomdN1M44v5p+scgN1xmV76UOyw+CDNy2rjZR55
amcivxo+07IFZ2S0GOwEwlaAtnPSdKvCe/0rvk92aO606Pa4xflOBkyRhLDEWSQ9
L0rEypZ4qLGgulwUOFxJP0esLdooV5SjmVmWq7QRqRgpffmUXlmx45P/cmZMrR4K
xuj0qHKbLKIZyqOMPoig9ZgeL6T5qkp49BCux0YpGNyRju0omoUx2okXsqdDzRsr
xoxhSWbKvLctn5uFnYhKXfls0UM2GbjlWqApCFVa8WmcDrg87Xigb93oAHCQCeM9
/fvnG0LXKMNfjR29y+tWEPHF9parqJtchWpL2jFJ3eDpK8p4L2h0erwUevp2tTU2
aNTYPFLvVZCWq+mVKsnBnc2dJ7aLFy9bZZQa6SdWALFHCNNxCQp2ZdgLrtWwWBhy
wp9sqTZxMouixmbea4QWkDr4/0EvgNIvWVeb7maZFaPxIO8e0JrFTEC6hwHYzLS4
XHkDgbt3AeK+KV4m1gFTswau5/JfmeD/FPw8xQz1CB56O76cnEXGF7jbpmq7skB8
BRIaYLTi79H+PK/x7eDzwajLq9PT08ruzMe7rlbYCQIbuKwZifjdisE61PfUrB8+
9c0Rjs/QVSIsFrhFZnH16C/8fxMwj5K4ap6k7I1x/IZvGtIELTP1/QztBbPZs4KU
Swq/thKuh/4BPDnV4vtFx2O+FioSHX9qwCld8HiGq9ISkoEeYuFTGKQS4Bsd9gO1
bGJ9uAmdzt8fqVAMK3BnQOyY/tIeJbEWIAUJlR350e3cJrJfJmAz+J+jyMzpNu+Z
XWRSNt1f/wMq3XBP79hmDETfSPxFR4LrdaIDTnfwbpGVVl6ecAz8OtYVCYAxDPF1
B4AhVDwcZfszY9aaJUMwrPdy2MiQfy1rVkx1OMymqduwl8mVBPavMdbQoevVwG7l
Pf1iOR4oUMkHbKDwFXUS9booHeO1UrKvmeEP2jhEDOOKz6ctxZ71wf3gPzetcfTR
7G4p2oR3zDcDAkIEQ6ZEq3tfJ8L2Fd3fjNYleuSIyxzD8lpqaOUuRF6+gH3BTuRt
Z5vRzKgCWWAyYuM+S0/b9q3J2QUiyepJHUhVSVkg27rk7zQuCABPIDXRcywDbajG
faE8wLM57U987mVxfX4+K/5OxrRMi6TVCAFwwdGSIIH3z2CFUjMRmzRuyIEFuwpZ
0eGvVou0zuV0oJCuL6ugJEqKoYNn1Xf88QHVzvvBrDW5lr9raeiMDH4bKwy2g74q
JHH5SK0dqT1Cjoy5yEH2A9qU2yoBl+PhqQ1cpsJGytxb20tNug/hC66mauJPqEkb
+A4gY9tpb3h8PMr7etkXWvwiBU/e8Wg31F9lhkg+IPWy5W2SoqtHeeqa8lDmm6BE
IjaaT/bXQUwzXJGt/n8ozKidSgF5Lav2/8Hn7KpPsIJQPXcUD4R1mCHmFQjWSv2U
LZFjcgeX8cqDfZ5lLT3afV22e+f4HTlxsocofxuIBB1KOZ2ySQtfXhD9+GPHJIfv
Dvq9bRLsN3fWUUNRnGyF8RwMlp+44qsltbt5ZtQklQPkPna+JZDTmwhGj49QY9kl
CgsFZEgPnXYEv5wVRB3hqQQNeC5uUbZgWPpCNDzxoGZT1IY7AEDhTBAiMZIcDQgD
lEBJiJQFeXd4/PBLvDT/XqyZ1s0UuikVq4JRVVW6j+FzdsmM23wyEFdT1kxqAioY
alVOJik9Edzha1EjzuqCtBZXBPe4cY9UhsSCYUlIH9I7QnImEZ5JGuyEyiYFbrJ8
Dq/v87xZJLI9YSVDJyqMrYBf/Ha4I2iMiJYXxIeMb5eJQirebH2SYShucjZnMu+V
TXlWznHsZMOLvqHgO6CJWSqBns/nuX/Kq91K6PblXgbCtLnjm+CCkqJM4KKvaL0d
yvsKMxFLUBW9ZA8u4fPNdDQ3XuJ3hw94Hj1GBx/a1tZ+idcqE/+9JgDtE+CM6niT
lCGos31CKUR4xTKNUutFYdzwONwlSdhyvNDf8EXnMNagQovpjl3jjrTOesQSEgSt
g3YFZtjCoS2sYdl/xckMlDOWTLnKZvuc65Nkjl7VZsNPyAdOaGV8IDszy0UxXaf0
oPgOTzd3es7my3cshzj725c+ulonc+w9V6OrHDqsAQDeo8iF8nIWia8Glb8EIxvw
6WCJMdP/ilBH6oUDlxo0SaKsAW2Q3OR1WU0kwWuHvR8JG3lDYQDwKpz+VHYybG5n
NSOx+8qd9iV0YHmArKWytLBCO4HKhYGB3z1dtAaGUHwj85PX+/Aa88yTV2YpNYfe
1HPPZJ3XwZdEJHHQToQ4s++WwfB8IJV2SOGrd5OefEuTsHd1peLlN9yLFPK8MmNc
3xH1oCYEMS17uyUxsv+rTyNPQIvxJkR6RFM5Q9LpQQPJLvPNM2fTzrEgq1MNeIM7
HBCJKm/08yguesQWTyD/RL5/3Ld8aEfvNXxTt7KuzOduPQ0Mr3j9IEMTC5TCE+H1
mNoFBgqhppq/Uj9/pK/5j8FfNSSo+LmhLctwv6AUhxfmBPqS0GKFEuDCGnICOeLH
gpwkQ/Tj6P2lhy+JldaN3Xk0iaSEojaNQCi6lSnR5VBjumBiwGB8lFhLu9VBQ6J/
kUhO6e4BT7idlDPUSNdse8PXM6yqs1dvId1L3CcB0wMqfWMXb01ZHwsuFVbFfoTa
ivbZYbioQlZNhVrX4r0JNFvTwgB51niQLcJ3XMNUQ2qKTkASiqhHOao5zmarc8aZ
GSeXp4qXkTQA+mnpaxE8vUI+wWgMehZCohxVM863qOy1bolIprHL7QFS5xHrQ+cM
acceq1QX0DRGb/7OL9BPgAVg15fvze8wEsqDLDjESo3dzPnXUnSqHwGKm4qAKpiq
ca84HZ6eukk2UNfajRfptBjYOugeHrcso5u8yGtmPnC3/B7Iv0VyFChGMY+yohkq
8fP5nm1ZpVGcm9fM3j0Rq8P8isqhdlCvd0B/AWB0y0Cl6/0wcKMRI8dokDbwqqzH
8lBj7Zhjs56E+L/LxeCVdK468x6G/qcKZe1zaoOyvoX5me9tFojNrimNvsTlIjk+
imB+6ylwLS++5hCUd0IxYXZdc9RmpUUbftZyP+iAfj98uO8nz085DYP23vwqW/X5
sGcwdxvueZD09Af5W37BsfnFvSHeGzHsZVyeQMfZy1dzcIySVm6uulmNXcAXVset
3KoyX8gq1iVaZMrDACJgJBzg0Mt+s+heW/NMIcat6m/r2Ej3qYgCA9Z4WQkBRRy4
R0O3X8MiS7/tpDeAO3IOv8W08oAdorEY3F3G3qsNPGbxBliG8CehaWMBDqC9wSkx
lMiD4QWQyTMzoW5QoA8QXvPPh4JuHCWLHqwN4yFOvaC0LWZz0KGUtqng5EI5lRyO
GqWlMFbCRtl1FkgnvGw9mPwFssJa29zK1nVobuFn0LMW0SIMijU4QRUdHRFxkNWY
8ODWWjKCvbUfMFywXJ8r+DgEj4X7y/4fUp1ijvEsRGg73oVK94kQxf7G/KMNfu8S
uSBgxIgAZFNP4JyZfCsM3vtjfJnl31T4McEy9kZsbRc2Td2K8CRLmEjyXbLkYLto
UeJTt5bWfo0gqe3WBrcpgsqHNEEPBnHmhHwYknTWj9GenBqaDfgWjCswnQsOHSG2
5XpwB/4JOK6AhQSC1RUa/HvsBGYZ7BUH3AtC9tVFuhhfTOcvncXCwrQVudZvoxp0
FdT7s930Q2TyydPVQZ+X85ynWfjzohmw7P+j82kv1iz2U3EzXqjQJT4LT3S/9NFq
QYZ+/5oaKocbQGGwXsf4ofSltawprbogSKnPAfVL8Z2GPQZPdUXLF1/ovmsFSxGp
y+BjIYRCxiz4/BRBJQlVkITmM6RmA+OyJpTcNx4RqTxfCV7jDv9gt9XIE/91G30q
32er57Tqv+V37nVfHlosHozmgxvQpRZ73UmfpURG56bYYWAtplTBTBuL0wZ6b81f
3n07Hz94dUWZqJ69dfYPFsLNCkRJJ93JZSzJWTkgnh4FaXnw+AiRgC/Ucr7OEAcI
Wqb/Sa5k6O+ZbBOKpNfs7X7ctduqhOjJDuBX3LzXUTn0yLSMqQqF2vyA5bSsRo3H
RJSv03QME6csiIRqgwTl9p4kbbwzdKHfqkHHwY6Aes1n8xqNocA0M7WXYJsrjm0j
019xB//rxIZxMBVh6eoooKwEDpuXIVCPITrrAEHgj++z7ECzpDr3yHxwwEHYrVB8
dvdWRRuu7/yy5mdLixo10/0x7pE6pfdn/oMyfmTX9cK3jhsEHnf3pTws3hSOjjgH
v0FXKtlZSiLV6ARfnTPB+8jbkt6Cx7gSFJZncIbdVl0/DzCxhQBdiURICb5m1zxG
yFn9TvpXPF1zaf1M8n7w1mu7xaYwtOYckvbzOHIOzAiu2RMJW+CSiCs8t5V43C4u
Y0smbzhYbBI7OFG7MEepfcoodX8BS5dJ5Dn8StaeBj0=
`protect END_PROTECTED
