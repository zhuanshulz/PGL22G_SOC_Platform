`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gUHrOnlyjnNPokWAn/Q9DRPKXp6d5AVVTZpg7GFSKXTjzUWBPB9Rze0Y+BCQjVwI
JsHBYXeCqaxKpBiBu8MUG85lfpHkwEHZr7Fi3gRdI0KtDLFcpx6qsNsZUeLHYBsa
XYx8dMR5yFIR1q6E6qdHnetEeEYAcQtbPT8D5IsvZmOILvZh341jtv5T/YiRI1hb
pZNR5W5qXfPt1egPPvW8+Esgb0A3dKj7wcMjAlnnHd/fDFGBIoFQJWWnEq+7HsvO
h12gPyGm5KcKEIT+JTNg3BsYap/w3hWjHiRyctIsiRfOO8jqKzDqWYGInH0RAbar
+chMAUCmS5Yabe7q47G5Yxlzr9Zxkv0Pxcx7nPldaukdMJRkiLg/w5FL3C0Asb9a
KImYEGvq9pYYmxrx+yy3IBCUK3JZVcsNNYmQMQYFSJJPncL281jenJ/QzRKjXfM0
Nljt4xO4YMQF+PzaC5Npy8o/aMRnFkfb7fbyCOUEm/Ajs18VVGb7G/8jc/KZywmP
XgpGeHyYeG7yQCkQfqxaPWc4ZOiwCd/cA3xIS1T/TkHbrfTiYaZJWIiU8Wd83DeP
`protect END_PROTECTED
