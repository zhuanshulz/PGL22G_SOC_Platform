`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JeN5Vn14fuuJvdY6jY6RNiLQdlKk8PMCycUZeZwv6c8Eec+TN4wJ+oaQdVUYfDTI
XjUsQlJu1mfUCJj7aFQnSiGh77LVg3FDUKffU8VCnpSTEwGAKCCcF4E4cCnmbR/C
7h69sePZrHF2GYfClKKlVt3ihLuIk42DKEu8FzQWYqEcIU43pxWWp/92s1ffpyZZ
QXkPYXQu1EIEmAlKTooiZuiW9cZ5nLbT7pHyhAr3dm9lVN4+L1nSnb9nPJiKwtHA
1SSnyiRDEqrAEy7I6iSXguX2GSxCu74+RvAJrg3rcTLWXsjrwkejI1pi49JtZkYE
l/z9E+vif2U789J8iE4pHjb50KfpV6pQRmlm4M/HzNujqGls715YDiDgCPX8v7I7
AK2fXimAJsVkO5t1smJJEuE7YIEj8z3TLQtJ2C/aZ1T04e5VoAPCPORDe+vS0CQG
//m8BSIQiblKsdTcPpbYYARnKMqZ2xbj5DDe6fuRaHI61gYNddGzEys+QC0KzDuI
9D13C59vwJfahH/RQyzaPXURLf2JzxF+7XSYvsxiDvDsF527YQmteAa0J1J/AMBK
tmQueJUkQC8MvH6i7tlBJ83ScuL7nYi49OOZUBWV+FwnhQkdvFk8w/X/x5Dq4WYq
/cBPg75KFXG76q8IF8Y1AeLZIsvg6c9XczypSb2qvAX2PHtyEqDu3j00zs4BdLCq
c4erFqo/1PCFEdAzZwNASN0RlWqOy/KSVTKn+KkFrsKEzUZ0uHQ28EPoaBLcajsq
Bd7HbtD5ULoLSWbiAYozIuiOScVcIY9JCL02KjWb4UHDW2RTPWQ9wiD7b9Y++P5K
6G/nmOuKvWmr7HJVgh2BRQexjLqXc1x3T+BUmPlq42ds+4HIGRZu9YWNXBUZa+Xt
aOpozXYXZRfhnmFwnLXhDR6FF3xvIlJDrFmi8yaU1jhhEWSOrHjW3ezUv1cRqzgU
CMvD9AXchWbvix3ZemtLVI6xo8d7pjKOSEOQU6c0FBTXh44C7zSPa3akO0Hp3HDc
kZ+SFAeOyTK4Lwct0d3hMpb//oIrUNhneAVJzQY+8UINA04R7iJiH/X1A/jCKEIk
XT+UqDXgsVSAPXM3l6FLB7XQE1F0qWZyVk+h6HS1vQMzpfBzEMugHtIueRQCAUG6
nyeHleGng5v51Ygp/vE3S2yePRWcpYv6CD/FscnDdMyIjfwLuKTIZpSUbw5CYjpC
e9NsFAMG65IjsZiPz3Of5ZTIjR8iHTdyxgRXuva18559k5gV03QvU5sdQvzAy+y5
NEBINEF/Vf7LFAQGO8T9TNspKnpMYIaDE/mHpy94ZO2VMWRQpdVv2/ez+gsG2psb
qxONd4DSaGJQcbEf8cjFp0JKYJqpi7Al6SBoo6kaYOAfS4oHGqDBdD9qqdEqNozq
PHIY3a5qgyohgGP6yA5+57En8+qvRVUuoPCyMeiYCLgSPnAJuOtlp3acilWy0Pnv
4d8gbVcpTBsZNaivutnJCsOBMq/3j03p8MjMimWrcpI3NbCiIc248TtEexCvQtFy
SrLbWk/5U0A4v/EziTdQHuVIr/JCw+0tce+x/eFLjTNT6sOn7+ffiwO3GXjVuDlk
20csm14eZnHKiPkbfTL5gJ0BEtz20YWJRakYvKy+Vgb1MXJgqIT3mMWJ+BDo9MJQ
s9D0EsTjI2tIUu/Oedlq8a5eGIYi7O3czMR09duvbbqy5AeAA/MArBCOCViAdVC4
3ByoekjiNod3vmq3hEnkgqhvNHeIg5LRWWv8+rR50AW86RqNCAKmZv2yNqVDjVR6
xRbzHn4Z/Jy34u8+X+1gV9tOny83obsCQ7TEzQ9ROv8AULn/W0tDZf12g0ioUkkR
LwlLqWz3E69yhoBmO749rf2FG7ST7HslrNvlEWy06yItjG+TbquiSkjtL6Tu5GAB
9WBQrQvslALhSgqynqvLpeYDXQydLrXLSbp19xCeeRP3C/eAdeeXDAEyhTf8x4I+
u2rSKwtdPyYx7Cd5ngcN3c2OVZ1bEbZ1UNpYSbOhYYTwt8gLDoPaiZG++utoKdKn
zfRoXFZ7oB08HRSLco74uQ2o2yKmn6t92i6b+0Z59TlgnCJeUfyxKD8N9ysI0Vo2
iZJPuqkIu59UVYaol6qpvVR9PMzrnlilocbFrUGEVaqNSiKNXDCIBQJj2kMj3P4j
D7zKOsCxWQanaxyXOM8MjmKO8HE3xXaAppgdDrZFcxnaGY00ujwTLe/N9dGKgJLU
KrLRDv2x2/eANu9evs0bmvhj8iCZa14VNrlgaEJ+5fobspKgXvUpXX0K5Qe1izBo
IVwRzxzKKkvOdvre64A6xUgG0I3iHsjbZPQTT8Acon2+BKMje9FDXrHrs1dgFIWl
igW7pXhJdqq64UyXZ9w4/KTuEoz3IxmbQ8lQm7Xv7OvhCvjtMJGiYN3lr0uV/YEJ
HqxfKYxMy0SMWAigF67bgc0UhJUb2YvZ9UBYynjFx8wLQTpD8C397VPjf2zwhB7z
3X05Td1wGtP+sOwwuzIsrJ8sIg/dxMJ6RuRs7p0k/6Kk9zgu7v95ob7vU/G8PPeK
TMwXfOKG1volJ/GKievJwhwvIg8ggmIQYobdmJNVI1oJXbFgtKFR/xKP22Fu864G
H4stpbkyFJPjDv+/q3Qw7uBGyZQiLbfj9EdSFy3axwwvHy4Qcjxp69y0alu7iCfQ
3piA7cCAW8Jktq6qkG8QeUgpofSYrY8scN2VoRUP9wviITnrGqCd5arsQ3S/Edfx
oetrMDrWVR4KH4QR5pQIT0T08qdX8BcWfwe30rsEhfnolUBOirbSvvnzcO2zkLq1
/36Npx6R58An3eSAzRLPq1tiiiaM0+Rv/JKG4ZehyNnOx5vPI5AsN/d8uLJqkOiY
83rnftLQqW9w0p2fR0mna9ILTHr/6fZUMAXmb3KPUqeewEXgl4cxmaaUE+wBoE3i
TJkGKCihLzKBB4xtMQ7MyA07JrmWYLApKOm6vSvYHALBMNDhfqkbJWpEINk5t9sw
SrNx5/mYopeT9ir0BuhFiCTVaM7fScwdnzG8xnrwwqX+fEk0avqmVoaSnV5dQi5d
DokwpzaBiSElnrwHnN4SknAeAY9Nvkl3VEKo0PQsv5+R+f4KLmxz31D7z2Jaulyd
B7uh9sLdjayORTh48E+1PKM50mZ6JR41A3Aw9xFOEReY3C/+zRzL95rAWXhWDdZu
z7Qv4jKWEu5mmSoPJwWicnG3rPIqoNEunnwVBz851B8rzOZMRNqZ2URBVrf3BaS7
ZJLCSDZZQQxbdhblrMMn8m4nCvJL0OWSTqOlLK5Piso7tqVyrPcyPZ6po5rbhNcj
c5SfqKQBfjh/kZjWTYFk9EuGUf5fZhCwUzszbhA6z84I3hsTINjh+OLgvP1pnJ5c
4RFBmE03ViJsM9SHi8fVltibEhyv/Y4Ww8b0X/MVdKhk1d/mDBnYQiT3eR+Zm2QJ
VOaQulda7ixp/yqMby5CZN9XnMbzBzBe/iIqS2KGBdL4GXMMxWFVM8m5hgej5TFr
Q6L+hWGmu7euAMjUlcXEdlw4LTiKUfqIkDSb88GElQ7LcMy5GS4vii7Zqyc1ynnY
1ShNm8+EuEppAfiPVasdgeNT47HWrk73MXvkr/zZ/lP8whDtVufVtdiDljbB2KHv
cHl9kvsq9eurH81feO0sjDpS9R7gLXT0N8afrdyVNe1gL5i5n7wq62IfZJKRKn/9
5AXLkyO3QvWVfndCpyOYcq9IPdB/xEMQhWlMM9c7XqtfieTjtCQhTl3gyYJUa2Gt
bxCjZXJKbFPAq9lC2IaysJGHzddn1XJPsa6tWqG7QqEaisOAb8fHq+9S/Yh22AFx
zZzFhgZvaAjJSnX7ZG4q2c4uDI0p+qkbcCSNNr0Fjlr5k9rAXMvGqUJWI6tcr327
3xhzhcVVZGjH1kE+5AO5bz8F3g9GYtvIjtuhV6M0Azga4gslr4PLJR817eIkIGTz
z5VfVTjSRaXDdHQOGCFiDv0HK/fZnsECtDBdX0irWFdm6frJHuz1rBEWdw4T/KG4
3WkSCSNoGDyFwWeFI/g0mO4qPCDbZ8tYiXc/4xoBZ4jaFET4kgziBQ4jP0UDMyXH
Cd69lKxjdtyt2/LMTGdzC2BxIdIdKVu/0UZCDXHWHdBA8KHJ8zOAVzR16Ks3LDfz
piekz+7wQcOYqreaG4Ivu8SMTBrdB6HmypZrGIpXFthAk7fGpm6XtuJaySrMuT41
WTieYaMqAysgdNAGdpen9ZCCKziBtnJytLzco+psRvgAk+y1zyb+uhywE+Hhs3aW
Qxwp79X+5nnNGWFPZ+0XZsWFL2NVe3ckGypEkNXoqBFZXFydy3wN8bCuFFxrBLD9
t0tn9JTiCHU6BrLzIL1MvkO+os+4HoLA9o8xb6NHQC6MAsT8ljlHvsltVoFckvPm
oIwp3ZQdWdZaCihZXa7gnnxiXj1OwUK3j5rtHx4wOWpMBpb0u+VKeqWA0NUAvN2J
e+/26DuO0Yth9yE9crgP82Xk0p72O2l6BXasdbsorey+r1pP6BdF56b6XRSmIKG3
MtbXWY4Dd8YGGoAXNpPhbi82TwxDCvjiPfZeFVxznsXejNU/c5xIK7Wn8xzPPgfx
xWPBNItFVXhLFLIGzTyeQXNR3FPCjWoZdmrDGbMqfS/zu3R9zEEycZmXWh0TH9ku
bcwlKqGRwRooO8KZPdH7s1Z/pE1q+hnrwR8zqCdQzZEoRfSwAOmVjqziRTeH2CEE
tZ76Dc4/YCfUKSNR9ASYpCORNc74bUrY4bA2iPw66hR9xQOo7sG6chr8c5L5hPLP
QytKyVzfJkr2EvkyZuqv/hAMSAovVmlJAx9eYDFGxH0077fOPFE/hsQLVcHlEfWk
AnZxhaCjKVEE00B3uhM4YpvKhxFIsei7mOciT/ZRy1AaUDSa5lQjooVotXNi6dE0
79bTtZlqIYEmzVH7My+0CS8HzRSMimPMkulSnUxLpV2Hvl/BQ0RJQEwp7UwO0zNI
9aRdur9I2lyK8Xyrr9gQ2FEKPNhJWVOYbMbm1pKxxRAdmtqcnBSCeWKK9eFW5a3d
U/6989g+s3xoJyLekfCN3YOANO5jLJF+U9FwdDrZDsXlP7KH5gCWC/fNfX8tt+83
whFfS3yEVkz2XahYroAgJeFWgv3lFAARrfcSpZHxnrwaGd8RltBQ4yZKiaC6/oty
nU7EEKCK1p1pNevPNRFaq/kleTBcSf1u8mJ+/z6RRWFoMXZvdBID09ioflTLXXQG
h+x49lCGKi85ji754devAgJH5gwH1knARBt6Ccsp1tP5xuaCKsUFP6oFGGBtw8Gd
k+vCtG7Yy7CTqf85Ovl/Io3xyy80XVNDLSZxEnAFi2yPk38ScEYoWtRXUzpskMMY
PsY53Vc1ogKlyEvc4KQRKHxXYTlWtlCtNOOI8A42IfoUo9B1TBy63ZXKCGBs8hFz
/GVVIfBhVdzmwmcq7P3ulh8tpMNRD4WXZmD+realuuCa3UzncvK7t/uahVXnbJuU
49HMr2sr4Bw/xEjeBOV6l93fmtjNCQRf8KzfvZfZLC/3gy40EFZssNsghFGe/Wnz
+v3AdYYbuiU6Ayu+PNmvV9rJUuwiK3GjD2Hi+wGIlMLlDy9rqKmUgwd+2P2cTX/C
tG81xDG+AbSez1eyQtW0I8+35NPDd2e9r8HpcL/5Q+RXAOIHjqhpCNyUHz80EPKM
WSTtZeFjNqpMzvOJ5orVbdEPHu3vvUP9KakYVqxvRzv3wb5pLNDXO093l4RSTOtV
5fRORzP+eWzRAScSEMrVmYwI7deY0i0iKFfXpmmqAUwi6pXZVch+IOgjfFLJChPI
C1ku8IRtLXdv/N5F2O0Fu8/jqCIklFEE61dDAC32wewF/wlY2/gB3sSOEkzZdDF/
3PjNnCy14n7kGl1+C4pRs/arlT5uWmn3TlyYcXcNKaP2t4tY6+eH5G8WNpTKHg/e
6AdqraU8rv+NTU7MGPM6K2fmu9UUc2egg8+5y5fWVmwDITk5vtB2TQ3wikeSgsgS
EpjCMZCsQCH9WbGCa11FS414D47ivnTHr2yiXVMJlQKHEAn/sU6TE36QzZcRgLer
YwRS6zqqk3ygmYEvBktN3ccvWa8SlJOQhDTAXIAnv0QLAC1E1n2b0WERg0VNHlv4
zX+1wPT+Vck1LlQcmJfveKkBgQd7H1WgZqFATpkuNR3dvm1u0arWGlFZWoDDZDyc
4LnQZ+KOvzNy8Oww3tug+BTedSytFDoNQAcOc/AXJ2VXyVorQF44Z5Lk1M2hmt3T
/MiNoBTY2CwrDzMEbDGyoDZ/8Glkux0Cwo266F8Vyjrfc33ceMauDJiOayaAbncV
A0nSemddwD/NyQzxEe03dKrL2Ha/Cv2B4TYTSR5tuUBZkeMbu9dq/dFchgEwDOXo
C/y902Bq73FBcYwucDixRH9Jfady9kinsQbDjbxvWFAPLvD84PB2jThxXwpKoBb2
niEwXPx+T/lYb3WeY63vK0SGAcMqsXMj49AtWRy7/sgMG+0JvTA4Kz6aJGbkKq9R
1H61N1tIfwigoEZVFx6sOYrKu2Gg6p9HTC/YruRW09RvgXuOYbOHRHGgMgAnZDju
HVWshsJUrMxKEJKhCxH0+Hs3naMtz7h07mj235k2U76mWVrGzok8qwoGpGBS0XoK
36lglZhupnXYpkM9161R49OdgmK7dd/aUlrRdRzmmpuygminR9JwEq2kps+KTS92
tpIYbdEr10j0it0WeOxRal8McN++sjoj2HNXf9V56VuAqyJXsJnwY09YgRyU3gZI
iX/1Dv0eZOdc4z+7N48dTz7v3H9MmGSApy4y6crPyMsbaoPzAqSw0amHpf09vETt
lJdC+Q80RX3AW5Phds8wpiPl8doJgXfjKrwyXo7bBU0oSVkoiEH76g+HFNyh5cHp
L27r140D+CsxCtu+nVrlD/GTyp2+ypC9LqSgnLkNbQ1WKUKEdzwuUHmw9yYexnVy
7Vpx/IsvtIMlqmxfhEbQ4Syd2NaY4BvMj6xJl6/1lnoX5Irc0xJKPaXU6NdRyPRa
OQq8mb3uAq0BGj5ngfwUgNYkViX+VxILNJd5w5d+xTfiVh4JVrj60+q+5J/MGh5W
aMMY8zJr0HCMmm2r1M/4p0c/2YzC/xyvNyA3u53HtpGqjg0Ljca0XuPD5dfCTJZs
SL9oin7dp0oUKnWj1BPVLHnZgJjbWELKhhg0ZP7sjXGLS/8Oz00u52K1iCg+VkAD
j7W2iRlGX3dj0c1n+0JoPabzUEU1IVoBBH7uKsWl9OZB4aNeMTyyrCNOVzTKMCCs
sCr2L+0Z8jgfX3ODLBUM607gosFdgZNPWsEbaM2VOkVjlRcxpSJjALGJAPo2t1R8
8mvv5NBteCVN2NiP3D+JO/c3mIsJ+w2xOi+Q5S4GAnbe/KUZv9cyz+DxfBr1sdnU
9ThKcwuCuvbFc8tZyoqj5M5MBYDo/P7srI2ZkUXUDx3Suqd6qQvkVmkMha+WRsOz
Fyd9nMWooEyN6dBexPL4L5BTAlcV78boQGuLi4AQ15sgIcqQyLiCAasC9e5dK+m2
YBQGD8O3ZUYX5C5aYOH5jFyDZAxpOtKpUAZ48ymKrf/Bib1ntk3bMPgxt9EucYd3
wyhL9g+KOuKTnOxl7lJaAxioDkAIHVRszcBZxzSUk6X82SXNEK5OTAeH7oQNFut2
I8Oye0dvfiqE/ZhN2w3VCcuzDkiB2AlnHZB7dF+7jF6RbFT+ScluRh53BdugWjw0
JrJjF0gfZPXr/z9MLqYPhQ==
`protect END_PROTECTED
