`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B9FyDistql+UqVVQIt9byUxjGHCnMk0gxl7E7pcp1UKZnagI0EkKWM5SyyxQGcQG
by1ZKOPvHISwtGTaQn5yLTkY8u1wX6TA5e4CLWPtIsavw0CKbyM+S421EtXF7xZm
Xn9CpI0+eosutPWTWLxlvUAJuWvaw5js5dhSEd524oq3uZfV4zkb/p23s2XLOoRG
p68O3Yr+WY++WaXuCLg/T0kJqbfPNCe+pDkqcXYyO279x5iF2/7S8YolFWGy4ceK
Qe2W5pcITsUIX3vHx6ws+A==
`protect END_PROTECTED
