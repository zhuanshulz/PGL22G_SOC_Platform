`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LdrVGWIL2ncBdKsCm3ll7507nvLoU6cd6TxvhQE4aDUf7Kv5SSyvHkh36/0yxf/4
Fbus2RGJvE/P2tsfUdiTpHlpMxTwMsicDMvykAAjEjUHlYHduh6XuAfiEb0Sr8NY
Hkqn8zLnO4anXvwkMbpnDIFC9ilyhuZfZwKaUXuWb021LhjbVgquenlv3lga8ECd
dw4ZxmQJKAzOhd5Ud2g/eZ+M2F0wO1gXMrova5DTEGkThGwfpiIOqvOxAMCysjFO
RCLmkWFk/Oi9OGvzP6LLolQclijpMVBt1ENq5z2HyU2hu/M4OwqMoqSr7vSdQ9nL
ILipUkEgE/lc71MfWRWSoVdtBHuOg3yE9iDJJYL70+V1bntsRrW2XSlTD6/t7JRn
cGpjmS+iqW/q/06SePdQkFUVV3l8n5/ICDUht/F7Xdf83OSfYCy9BY4nCzqv8QyP
gvOq2KO0jz7F6BDSn+5KiNPL0DOrDzMWmFjOEQXMKlVv+/w85wt1WFY5u+J+877K
u7iYN22vvfGEM8NQ43MV50G0MRqUjewvgsFfKubZ0fi7tGRBPSakKFVT2Ws+7Fjt
G6XN2XoffFyNChyMBYrqOa1d5EQBZALmHvLdflssOHfWi2G9xPMIfRL4DVdkNmiT
9niwkzDfrO6OswMTyHI2u4+U4YlqgpWe1hngR4tbZ/LJGw68AnLgMittXGcckp58
d+Yt9LvrsPz0kSxEu9y9v4v634OGEmLm/x9eisgNpSh3deRvHbk7skOaBsYu1ySw
UabHFgP/xQEZFWNnEvjIenqAfe8T7gau1Vg0B2rze4v6ddppGG2msTtLz46TlStH
j0UAF++1WkvC4nUvt7dU5zjRoS28uRYPRy0hunT/uHckk1MZhaJZUNAeLDVRTgS6
LgkATsth6di4DhVI5L1nmpH7z40aAW+l+rs8vHyeu6rlV6/uf7+v7Bfz83PaYUfT
J7yrMDxvJ6q5owu7D4t48sUh2ZR2x+doFzyd+uUNl4fb5PMiMTPHhWNBv1NMR8Sd
cpfmcRoBuGxML+jcodecC6NFihDii35Nq3wjsAjcZXs21y7JkSu/of3SMjPTCInk
ILliNRktAvJQKSwMXzfem2yth2w+bXZs5T3jXMLG41JGTefdCcy9zAZHZsNK94A2
y+WPjUy6M8g/GDP81qKQdqUNFkJ5VQ6vDFD9dqzZZ/gutPoaRovnN8+7nO0o2qOh
RtypBk0L/UogzzXxaIHEHgPE9KDpyLVYstanbsbtpuvTybQk/UsbgXH9TsRAgYpA
p/T432zLvxTBjoQZHX19eTSgzUzN9gnSlEdizUSEKWMGiubbzq8qTf+q5G1IT7GD
7bCDKIL5FBvdC5gBX+bLFRjnj14ZUVTH5HdmRTOfzLFZSeigGUqS8jkGW9uzYMKO
u9DXmf3HWc6NuioiKa9dQTa7Ttz+1FvZWAPFsvS++kC2CaKo+NYA5AgpBSqr0PME
Q0kIdfawfmcDXhwMI9n+Exl2OoH5TP0Uf9IL23kznqpUAGA8LJHCCPyxxHUo2+bE
yG/nD60+YKZigHOCUiuEilD2kvTKLREXkozAHClUsKk4RRvIPUJ8rr4sEGReQYfN
HcML12XYUuTAtuAkdSM+AnQYEaqQTLKeXT7LPJHWlJHiZewJw6nZ5VWcjoREre/7
pSbuKs1KsvycFijx4OPBpAvYJGnXxJMLxdXRCjC5A3YlgEm5XZA/qy5cvgRXFhEp
PkWQb7sp0BzoKIfin3U6yVL1G5wFrXnXSopTGK3tNMAuqrNd3tO7BaA+NcJ6XrEw
DafjwZTKlY6REG2sUL9ZpU2Xjoz9JeUCMYXIGLsDrowQFUEVLU17JoGgw9sE1Hx6
hgccVUdvkOsL/uU7FyT8p/vzTkmmSy/mYqA0XaLKFSnv+qg16gwutp/qA6dGb6nl
xneFFL3ci2nmqJD/MU1Uey0KNMKldyTnYZ0Gy1dTAfM9nD7Dn7t2VPl+6Ja7iaB/
s1zDlJQyGwNFHwEmSUtpmAELX4Acoo6Xvx6vhZuekbYknsUCPlS8ewh3lPMr8Gyk
dF5YmJXtIpwXDVqpQBkZlp+VxHAeUWb5B0JLyEYuJ1gfsy5M83NX+HK+P84lBYYn
MsL595xPp6H2nMSgBynhp4lunYKvntECcdHjYBf2LgHApQ2gg9+nsw0bhBgFgPiM
ZmJc9vj0RFjSdlQxLJhLu1CeOp8QhQ51VOsKpsdUEmwJEXtrSzJeFcmn6KfwTFFp
b4zX4Sh6DoQ7W6WQgv+TtpIyHZEw7DgdVTfsMxBlbnC6rupuA6Ax7i6vqJy/MBc3
AtVyxPxQRsknO5oO82RDxaQX+oKnKCIk9koqEJzbn1dJ0qQdjcMw/BtzAs45VMoG
kU7MgoBZmFBU/nrYFH08BNBeKSEtPCqrF5imC+sRRbHDLXDr0wyrlisvVfxBWOEG
rX2Fe2S2BoW/L2KmIeozSKJrJxnjySBfrPeRk4p2ycKNULZcP3Px6noZDTc33VBJ
ND8NtqjOFFWwYyPpaWENevEyOsnwYxC7AmJPQMlxbmRtufrUatYEMH98mPNp10io
cBo0mDxCyjy4DKfdCBodvLCwav6p0bK6QIEEdgITkIxhQOBWC/wWY+zzMAD0xded
+il5pKZ3H53lIpTaL5W2TYoi06zt6OvyfVEk0I9OFebnIyCPD5xTC7sUCWFxdfjO
kDH49QdvXiCd8zDph1p0Hhg3X1DLJVur2o9SddzdH98XsKa2dQ+9BTMh0110xtN7
XkutyNa6ePM3NAFYO5G2VkP1VhAJWT09WFeZfF0eerKlopamvcbzNiYaBfmVGMLq
5bqizG2iZACs+rWtEsOt1W1vSqwUuJDzXrobDZt26vsJMtOxFrSxHKL8IdeocKGs
GvdaTzLY7BgthGJJAss9DUGVFhMEX/zWOk8sPt8mlmAjDqsZ3bKggwB+xEUq9Za1
eNz2LceCZAe46enbVuez0ax5ul2EkunMruV7Ao0rnaOTvzi0v1LQ5Nt5hGVSLImS
YH5lIQfxGviNDP1mHBk6MR1O/1aR12KLYlRrA/P7t5zypHCv4MqY/UjsuZH9yLOa
WFQJjCI+wuQi1F893oLXERdMTKYSuAvRcBnYctjsAl7DWmWZL91PhEPpNHdkh7H9
yitJB4A6TF3o78a62liJqLHm2jRPjTZE4b0Pg2JS0uQ03NXkbV7zliBP8qaPFwUo
3/zWj0Y39T+POoBPaFtxZHoutAg5MGlfhCNfuVwvdOQyoPCp+I+R3zk8E2Eu8un1
xYilVv4d0tZ2P1LpWVhoBCnKmwo6PqhUrWUJfC04BMJQx001H3OXtaMnj+8Z+8Cc
1xqlr7JpPmsu0zyph2RNDXP6ymQdSDq03BVWMqb3BvUsAv2ybQTb9KIMAHhiKiP+
AeTzJNllPN6PObc0iirnA35ZIrOByrko3uC954GaC72xu/bbNoCDCOCQ+dkxARwA
TnIGs5UCW7CIcUx1dPQmSJ7uYpMPceEGef52c7rzg9xQrWzpDYdMyeKEhiWnNfLB
zvOPPQwAfX0egslnAyTyq4qRrFpu/MqsJsVdwywtPG7SnvOXluWRr9VuLNJScnfS
WildpYZR+A3wU+LPo7bnkz7M53DXkTI8DU8ROxtLyN8HR0NIwHCyPJZ3/rSJc51a
XV7EEfm9dLCINc/heXAUsG9m3F8OJcfMA3qLukuNQm1gox0oo4xO3cyXcpmnq9pj
7Riils4DGhWePRe3JGMDxaXn/duqcL0WOHDGwVgJrGKk3cFIoJ8LpK3gy+BIs0/T
ByvarAzKs6ZTzMJg5w6/7nSGcC3p0PLloKRZcLKvmg8dAel9uB/cI6s32tYHrE7J
OhbjBBw6N1OFYz1mW+E4lk5INY1ok6Ik80dHpunIsPxX+D0D6IUNJz8RL/WvPGG5
AinYu/j3LKkQfqZ+FKlPa7+B98AvBTX+AND1K2BpBL4ft30wiVyR06rBmIjyLZ5Z
OkhL/M1OjXsz0WNpnnFGGCBbVqalX8icpY5z9NLJooC+94JICUE3IclKRmVJXOR5
Su+1NEZiIUku+HBf0l7z0JfLKt84rXlsDWie0nHV16rAFGOB8fLdH4b6oKD3eaf6
ZorpH3OqHpqeUnsN5n3/j4FshErBQCIkAF3egqKG0XtLjpSKP/hqEFyp7/A5EL+Y
UdAOUom68C8xjM3TNd1cbQVvvZKgl5Pav+DX6K7RbyYpES4D1k4aDqyyTtpP/Qay
dbzNyw6fl1y4mj+SYg/yivCgPdihIxfDFUF1abXyNYf6NvKQOn9gfvacBu2N20vo
qSp7aqBJXzTGcJX1/X3JA4pSUnFCBRtWguHNe5pDR4vZSIs7owXL2UVMX/CzfL6X
reV8Ge2k5KY3VIMV3x6YHq8YLH6/dnFIPnB1s+mRC8p6VgUmd2DCZuWNNu93CbZU
2+UapLbxRqakKcrNJIz/tg==
`protect END_PROTECTED
