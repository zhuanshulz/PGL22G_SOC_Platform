`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OqTIFtSkLASGysClPScO+zNj+Rz/kSsn+u/UIB/R+zEGyzvKHjpJQ6mSibcAOoPm
nR6gkpQYoTieAIAkB/rK6vlGQ5QT8Mz9AqsIh0y4IsdC/UW7dlOoliZKPLFxEZ5Q
Ss3NJqbmPndMhUXLYW4sH4NHqbpQPI800l1AQ4Ygw3SyVtRIYewlIA4swt7mx/7E
VrQwKinjF72kZtOn8RVKX4ae4sCOvn6OgIQ8JWIsLnPFhLF9U3DMwBMeLmTKBv09
zrvQghi6mwL91v/t+j+DyzwFLTSIlYYn2/g/yvZjW9sJEMK2LUBCop/efd9uvEPW
RjNRGBVfRVYP5PGC7YIRitnm5fETdJzLmyMh6kbbE4SgC5//QJY8lFtaaVZUq+8u
qiMeMUmFZA69QIHq7y2Q6yDf+0mGgHulO3rCCo0z/7bI3dumfPrOQQ3VcnUgRHsW
Gn9qFgfTPxBFC1tb09k/pjEpsDD+4eJt8UUroWQajhoMaR1ImFgFXfDq2jLYOEDN
7JZ3SScyQCMXG1QeMjxUceKkbl3zT0qJT5YJwEQCSqpo1XUTdUgz37GgbOUj6M0S
/gpDPmdKUX+1+JThe2/BXq5hMyKjDu9SBq5XzkUuGAqX+3Y9Va85a8ZPsWL2o4fY
yDTj7xlePBEEpqGtpzi8zlQ+srzmrEXUjia7VrGb4Y2o5IX3C1b/kEH8fylwW9tW
M+MXIKW3f4Uj/N1DMLmJ5iNJ6sDca6dGSJzTxzxzel6FID2nFqb/CVm8tx94QcOX
SDsH6jCwhRBnpcAYNZIiwz6FGmLeBjKK7z59vEnecmM+Vbz78YP/YXi7m+TdmO2E
5+3NvNQ6zhT8p8ylmtOjeFfeiYcWDaPTd1xpEDmta0JIkBbW/3YMgNnSuUj4/xgO
oM8Up5FmiOZ5hbkcEMf0OQ==
`protect END_PROTECTED
