`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q96hq1N6i6odBL/uavr6LeQZ5TIM7ZMWESOGCd8S+2MgHqItOM9V9Sj6E020gaaJ
H72jHnh6s4eLCseq1TFdha3L41EOXPBRYTMRw9N9znIsHdRewGWpDK3ObOoCzDB9
ZID/Deg9nyxBicb8CUKjxZNe7JttgUyX1ToMT7+Zwuu7oLLPGQpEqAStHCV3CUgx
MQo6Va+HrdLf1YFQwRrZSX8HA32G9luzPkbD+G/YKBoqmmY0hY0z02oHMznSZ6M/
3k2k2DsJPeWVWoEmAEbB6IhY90T9Bv2NZhJOVXKfYxfXyvYnhh7PL2bYomJY+Aqn
BRBsgfSXUSA/A+G7okge+uosJ0C/7RjDFRAxruef+YYNsQ9S6vZBI09yG+sp2U+Z
ZRiUUxUmR+B6iEqhSjA0yzeeQh8+3kmCmg5UjwoV27m+tZkItvNxKEChRZqy2uic
QFufpfHyAbVQweSzY/roRj0d1jMnZBKPAmTPuqI7aPUwqgf8daliuHLB5Ei0CUPF
fUGqM4ULXKUMr6D9c77DQnlqnMwrxZrDMhilyMi6M33QEhIxyrjBldP0op2PgeOH
UaTQB5PsyqcnR8LKaUblySURzGZay7kF1t6MnaiJfKlpGHnOppEBvR6wR1ysT1Af
xbSYXrn56ZA37C6sEG+WB4GRm2CbGWBWjN/APzvX4FroxsEBM6kijqW5QL1bcHGd
kTK5cvyHWBSZ8MEw12cd645LMQt/Zj5hYR5pagFjP3T7GUh3D2XDNLUT228yNuNh
VMYMt/ZGU36aaiMpNnR5NdUxNzkZjD8vlcigevxnPZJpgHA7JniS8dObcw7oDlNj
ETFDi6j88F3SoE3FX4Y4qZHoznAjESTot4F90jZrTZ4ZXAUhONjpGK74HskGHDID
U8DS/Xv1T0Z+znpCyDOutY0YLRw5NtkkiNynz4yyjrR/cMU+p+9SVLBv9jsR0HUU
SRjCJpmHPeZbXCppHCtnxgQWsYxB6XVrpt9Wu4jKkGv9mWUMNLU78h4DhjWSknWQ
ZaE61i1Cg8XmocSuPDNB2s38JeGkp3ZFGU/VxH3fz9z+XwUCgQz1GoXMoIByQ3z4
Um2gJxpT+/NEDmHACvrketzQChermBCum3S4CkIj+BOwPi6vbqZkiZNjDm7oKXMQ
FVo2AK0pd3m+tFWkf7VXOUWswclskpW/wpUgxR9m8r/XXfju17OLVaKwwg5q0bmp
`protect END_PROTECTED
