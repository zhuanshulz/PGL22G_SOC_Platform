`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JxOO7iEx8rvRLkvUYtF0tvOqGZKJwMdLRfZoncYI0uHaEPvue/z2voDr1I90Pm2Q
KgWlmZTe//Hc14d1/N77aQ4msE5zYR8lk2AHU67OqE0Th2tzh8+hcwSc2rC9SK/M
UEZCxALu1VymUTKpLow83edjPiuewOhQmLKDrmcfBYKw81ouJDI0FXFeadXtukPU
xhUZeOirIQx9P4X3K5df9j8DJsuTGfmEMHCtzH6DZFhhtEcKtcxzA7pA1+TApCpo
7NiH41YQgHWA9PdPXQotA+XCTuYwqnYX6eXU6EZ1wYOvZOlyw43yRabU5Vk0C5NY
vnCBNxwAQOBh3rOb8GuL800DL1BNRrBcekY7OgTb/f1szvL6dy8Mwkx/xHZ/mnca
cgebB8NRdbwJe8UacUnNSTcRbIOitl2bsb33GHG/Nr5L6z/kOhhm50oB4o7ewrNn
VnO5Y4YLdpZ1yL7Vn9EhLAqW9Md9eeG2g4TWFcUxeNmSIC4F2ilHVaIPKn64h696
YmCdpzGyAs/5Fbv6HT3hGliex+Z6W2Atq4APBWtK7oOOEswSmwX0e1B4t3sCiD8C
a2M7QdlkQf/8SAerd44zVdh8HiYnstl1oH+vmhHRhmjKgKWqH1maxWoZboz1Yr0A
Pd6bWo7dZvOykoMrKei4BG0lwmBsAs6r0kYfDRFIcN2/HoowHyygRPSnfIVmqTU9
0DSOif3oHdB5xJtu3RFBX8BgcOUmlIrA0xlHlZPSaPEx6rqqpdXK5P7LKohxq3Iz
zJTKdi/xNPrs0/nzeU52kbmM81t8irYw6tCU1LoLvMCQw18gkmH8YsQQwjkhrQh8
Y/ZLpP5cKztEHarw0zjHiGV9lMufA1tWRyNRL+43GuZ+7mSEeKVzhnygSXuj2eea
GGalc6oX6x4f4veph1VCv4C79BOkJavu/MhihwJUvpT01v5/7G99LCpAfZ6Kfnrq
k1irNtGNyTl+vg8rf5bvh6VSztNg3hn5AAf2/8OJdvjdYT1sOAeQqtLW+TWjJUSF
`protect END_PROTECTED
