`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aQWaqxAMfju395dyguXUMcSChwyKFbJ/0inXbBOSmOKLtbeZHl9vxTpO7+NmDIeO
1vBaRgXE7nrpLImtC0m1p9WVC/HomYgL/VKkTWFUc3XoEJ3VnMAt/CCOn5B8qqSd
ohouYEfEF5Oz4Uqoh/DFXodVf5kECXM0EEui5sEWNG4VRQcYJLivE0I7tL27ptvu
Spo+Jixickm70zQ0Qt9eapAt3VxXF9o34Zz/eZV3d80FopYBh5q8c1WOkC0had6d
Js1GmXtwkcxOyooKzvfPgDoPBnfBDdRdxBFEKnSxgBhCqHmfhu0WzBrgbM+ry/gV
IOtxZoDwX9Bq2Ddko8PPy3d7kWM7sbgrJmI5ZVU7XQZC0TY9SmXuB/IBWXYJqeEa
lKrtGR6ojtq2N/KUIVKdeimRTS09q2X/0WsNaM6WUBR0J1yzYFEn46+O4IMcD7+t
GOPd8P+1EGuPJnTUTUhbbMnuhcst2DK/iMFQzOMJu5PAkZaVt5+p7f7fyEatRbv0
YzhGpfvqEnhpgEUtTTvsU/jzMX8u6cpd9afQTnMs56G6FrRavmHbOYp0Zr9+YfX9
jqJJmVARRGKI7OSq7ArMMw0uWiv/pLV1khYUO80Ch1XeauG4EGQerkK1ZzGjuE5m
u535hW06F63BrM5uIJSLmtYWVPX1+FzVkXzCa3XcgC7jhMDkkqSB5rza0yf2D5V+
tZWexpEIScpfG7a5lbuRBzODFOLjvEYPUM53vRVRzNDL31d06UJxot5umQ5pUv31
ZzgC5s/sLTFuZnxFAt4jzj7A8+6ZXJu1UJ98KlVkSu0a9rDf6skk2eFX6AM1FjwS
GuQiLAYjQ7xhcYM2pgFfaE0POlUre8VWrDJ4DRGdGGxVg/iNllhSp8H1gPrvM7fP
M0Nj+ytLhUF9PIhEHwUS/yputr7A7GHU1wvhPGh8ionzEn4g0yiCtS6Qg5z0gNK1
QRipjFrKa9xaG6f2G66/fNUcHDzKxGlRXy3ggg+7BNT3gWzEFVLcCV7UWOl+ZvEH
syW0aOT6FGGRscnaRo/VGrd7przJ2vz9bTgX//AzKOYQLmN3XRd/SXVFi6xCnW+x
ALCRMOoRbhoUkSNPUrQT2u4fj/Kg43b8jO2wPGxmM6shAgrlU7WUkjb2G0vAoY5T
DagkmJditeZOF1HXXlfePdtEQW44bYy7LIZebf6tAXsiVQ/GrEXKHK4LN4MrbAr2
G2WSFHmWYPlRQmtrxBu6hn9nZeReJTdwzsywFFEFQjELVg8siBbZaRY+Ud5QBqfr
lMzaks7BvR11H1Ydv5x3ehsK/d/7n6Nei+iCCssAMIlMFwKby5LUTtJm9glYy0/+
B4wZyWuGrdhqFPTtXsH5mpjkYEksCpPf9ywlMTueAJR88dMC6cs/a7Rg6AOrYNKa
9meCeii4+4MLdtcsz+E8n6ZhoPju3wrQOV5kzz95RIboV57zl3LQ+uKwvhYF9esX
h05sG4ClgehZtjiLrZSIO2btfmwB2rdilC36LFuD+8/lPsAPLYe/x5l5dAYfrpWX
8perVXS+lFgpVOA7S/LBSG7BMINhAfNN/fgLYbUIp7RqaCHUd8A8SUIgicUxzYqY
Kjuo/fCi3/mAliSzVsKNlNr22a+ICnYvKrnOQmjY5BsxZmQWEvoOIfv+egSyP8Ui
etAwehqMACVG7geZpsBXTMqBJRfw9xSXkRmo2DJ0y+4Rg5KANvCGwrDe894gjKoU
xTZnNQ1lxKgt3VOQNtHUhXJCfDCPRg0G9gri9uNwx/aM7JAFqlu5Ueff0LfdMZ86
HyqIhkwnjArT2hgyVugAK6x7J8Ks8hD9n5Bh1irrhbqXuYvU5KvTZC5mrnny4zDC
9DURTXVBV5JBKcGlYPXHVnGmXMgQKFx0agr9fvSoGFfZo1m3I+bNRWjTJJAy2OAV
lZPi3um69plodOkw8LsN5rRxHIPctFAfZwh1CA6C6OKlszZZ/mrgEiuVoK4Gie64
nAzxIpvercSFZbIoTzBezh61lS3i/ELEJY2zVFC7htAUuYl7ved4lwinOmGjQBYX
nyRF2TIO2NyXilVVJqKYjsz80x7rRs+cWf6K0WUVcgVjxHFQPsX/1ZxZg0uQVaIo
2y3mr5z2lXWteoSLLXxPfJMPqRWyy8lWbsJ3eippX5sRr8fd7TWz4o6wkXO55w5J
nHbR+a7+c8P/Xxr4PPD/1ns9e1gcmmohOgI62EZ9t2gmU8jLWIyqOccc0zC1pjCr
8ZZFV1CWh/TBoI9Il7VDjCyiRG90pFf1xEZdvjv77FvF5wmMntf4srA1I4tkRRoD
XwMVUwxWemnenpW39hgnjvg9z0Tnyf/y1WSv+35Aqq7pvsNbn3JDQgeYhS40tRtz
fD2inNstR35JKGfRCz3Ww7yQQv9KtKzrKDppbHWP1z/zUVgTE8hYUJ8oWHbsL3Dv
wez/QUAE4WaBtUb8KyeETzBHi6s2LYmoFJaTDje/JCLyouFCoUraNuDLPHEg5VR/
3H9xt7jeTbp0O7hc2K/TosaSbSDZibv5MoUhkvuk4LntWl5SY212f7fkgW4sL0tc
MP7qNfoQNrEizbdFxqLpetrFt2JIxnKlZb6pXXZha0bgxwyLJHs+5L4BdBoSQzt6
Z7XSlns/oQ9FFKX6YY46wLuiz0OeVrAWx5zpKyS522gkuq/Pw5njdBMt9/2sAIlq
4jta7JWvSADxw4mHXnApEQ+AVjDrjCuH0FuLmohjdczsi0lDsR3pKvlbOR4TJg/a
Fb8viDbn103UXtrwHmu104RIfXr/xM+XmWjndr8tdjk=
`protect END_PROTECTED
