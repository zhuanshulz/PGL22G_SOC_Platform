`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k0nsf3FSX/U5rWKSLsRY1ux3osa6OGljKTxXxTttCWuq8H1k8lfHTfn4qLBYexJK
B80Hrr1LAjSe1/kcykxS7paWp7RBBTRCLPg79e+utgImypzMKS8snLP+VbPrE9sa
wf72ujvd+rCFUHid1nfDe5/tCbYeapSvAD4dnc1lyIdzhogALQUcXqEGyvJnrEqC
ywUFdxLCXRBacShS+inzXYtjvX1jNKWFmf2KYbN+a3xNYOo61XRAO/yPryhd9xeI
ZcmKE9FaLOcx7ffgTya2rLJJRnEXdzx+12Oyd/BCzOsUuHAO8JuNBIDTg3Rdo3hy
JFGPUrNtGFmuOTY3BQ2+EXjON++0fiFeZJw4UpnMS346Kbc5T80UcuFvGbvJcNnP
P8S5rQyzmNqrbWBMGAoBWjgTExQpZ5WxzE/QvjZum+KB+hzb1QDoIMZYVA2IdvbV
UQiUH1rhP/hZ6vVopTtmLWR7YlDz+mrTSKe5KgT5eTi79pIcuws9GmdGQUWp944c
UyU8gl40eDyYmgpYdOdsqCQgVvdBWHLeNnneh4IGnj24o+520ISsRhUM10+/KjgT
e+CpZweGCwQnvkhGUqSkoJXXbCpdIw2OFOcxwDT8Lzfod0BfYZBXEzhynBgw6IPB
yBjzRov0t+uKnrhF7U57iCQwIfXRnvv08bYYS/r5Or7pUQAfLEZIbwlPaMr4aDO1
3D53NlG4jsS97hpUeoCsSN2UjQURJscML5oP+6Pe0LNbPWWbxWLWxThj8aCgtfb4
GfrAPflAHyE3K0Vob0m44+ws3ybHvtDJSPEAWIyFHmgg6OmLQq+DWCkNUlVn5dh3
RFAEDGZXw6bjrYb9BITtCqBB87uKWyTKKEDSqkJEtwI=
`protect END_PROTECTED
