`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q85BVJhZhrcWCwkg4psiZgnHPVJlCtau8jz8+4WAiQWaSD0RYVRXH2N7x2b5poXW
/0HDIo2CcYnC7vwXT/YYB2vzdIPOJAIcTuv8JkBJUXe0rOUe+62KyaKiXk2Y3fJZ
dhbCaefZ2krcucq1fyE9F5BZ9WLTOoD63u2/kq5DAtsLLb+4jAvXH5ePZ/Gjr/Cu
T3y0Ip3GiJzmef72c0NMCVt8qIa1EhgVDZLQ0j0t+Zt6FHDJMiHlk1TJOWlM0Qrq
6UU/rpqkXbsgTHLoKId70VkczsL/Wg0AC8G3P7+AB/O+k5HaU0sgkKiFH/CN0o31
RwF4k1gG9PTEC9qJ5jJF+oDkpq5nGsKYt3D4wB9lWyniDZokzQW6HWdYLroDebN+
73dyR8BtJXKHtvjmVAGYkTz8c3n+W/FXcmQC9EGfri7HY5ANpVnqJab3RcwX40QQ
5FCqaeFItpmGcqUSGHBjBBKLW5+UgFHSSrbdx5txT9VIoO3VW/zPCMRYytw+k+Jv
0PRS9s4em1QF98/Dzm6ugQEYgmhIgwmrVOavWFcXSlKWOYBey0dXWWqweGAMls82
pnac0FCxsM1lth0nLc17Lu6yS1UxjbAQxzxNE/gmxM8Cb2+TAbNsoveJD2xDPUao
FnxJZq75F4Q0dkUoXiYaroKN1mzInwZcxH7vqdgf67ZUKKCbv/UL6P7kiQOQJu2z
u2sG601dlIR3mTnLld+evpRKV8qftx6t0m+RAcEdrbuwMteES4SjUp8VNKs0nKKo
g3751EgWM6b70rel2AtTeMDRBBiUwRVi3GjrtmspsXLqbnFf+QNkAeH5BTncD5aK
KUSBlAHs17HOMeZSHU/6j7McpMwYfjXYMTjPdndjTqHbaZjUxRbMcH2a9Hs6tRKm
nZ259qJFCx7Bq+CssdS8t+rdZ3X57SXp/sx57Q1A3bE9yj0SXwo3oYbzbMV/+m41
YmOU9fm4gUEm67aXH/ib14Dbw2TX201MEBJiygJ5ITmQGvCRCgLhkI6spJwfcCjD
5xMLgCVSKOlFc2zkOsE7ThOBpBFDwwiE1lVtqXJe7dxKY3SYziM+LvBl4OGhAok9
HBpuMY7Xz8KVdLTL1jSXZATbjHw9jadmfAAf4U4fbVTw50Wms36Do2fwojZxYEZH
N3bxbN2mGLuzXciBoTFb50AL+LS51cmup3ZJMTv1OCNwnp2ZaPaszpMQatrio75+
jJKoLH1tcdzc9Sk9nayvFNxdfP1W0yhnnh6VeY+8K2ALH/F0T+zZcgKk6AlWf+6h
/9bfqQKdRCrwvPpcIqL6QNev5wea7lzpcFm8cIxXLgsoYc47KAM4FRr2oEtO/U1Q
GkwUkvyHdDeC4DxavK0xZJOHwkReT3KFf+8rQpwMO96LJ39xVjEAFSoPWa2qoB9v
sOnor7zOfRLtuDJGstRROhC/ewD1FeUB1nKFKMQKvTKZEQWUxqWpqh64TctNWO4n
Kh7VbTZ0153+AbpR3URuMr90pD+QvYZvpjt6xP8fDtMdBEKzKnLYZopbMSDa1DXh
gRRcQR2FQPCc4IUD5W0eJy7PpQF+fN7e1KbEGjgN7b9DEnf2x7tkwT32Gegecmd1
3Koe5Udr0e+VLRT69SQtE2U/a+ba2LqSRGmwKTAWslKixG/4hw1/1meF6QzqPHbD
AUsGS5rT9JZzSGmEsV4bMCROCaTPf9emrS5/e1aU2S/ob0KEFw5znKE2Zqhz8MFB
4KPhOGZFdFTqDWONbN2llIOTRUDRjJ4DairGnzJsia7SXl9U9PZOpCXliK0clPoe
aLyucoaoK0VLtYltGJVDm8ktrUz1J0Q+PsyLnN5CiLIQm66K0kAyTPOKouB67jzt
/NMhhXzmEWDkpLWrGB/MFs8loxn+ufO4JqaGeHAWIMR51cvNXiEGo++p0T/81mGk
mpVDVxDJltNI5orKZaR8m4+utvSQbhy9/q07UFVEChGqkO24ro7mI5yJxo/7VXTI
z5ooCvMFm5u0WuKP7Fm5BPoCETqgm3miZUW8biAeRcXm0NFGN14anfAm4H+/53SJ
iiSM8uyRFj+ybXcJZLud2/sk7nWA3NnmJgQ4j/a6vjrOJmVwyDIQnkxZYxRbLj7l
UO+o2njN5lE1lwyDE41LXpG8/WBxs+lwRRyZJzNBOfhyySlP0LcbbD/9/EHUkYbr
0H3siSLD+JBwcqEUeeoyXvzhAkxQOiUIWRsY6SzMYbP7F5fhokyCLwUre01Qln31
9GRSedfmvk9kMCBA4rkN1RmA5JUtFaPPZCZreCmWNTJKivXFiGFryIanfgZlP+gj
zs5+5k0piR6ua/ybpv1RHPwqfQc8Aem8SXpiI+eourR6n48zS31kMAfXmkQbgIUE
aA5rlRsZlCHL9DeMsVsVXAwFcckhImsZnsWu0qFQ0MaTUJcX9ERiOtACD8t1NQqI
08GTQY853CWP1AHW3+wv9C4m1uoZc8vo8F5QIfr8wqacg8lx+TQwYh1Xzzn9LnNf
Ij8ffB++/6oMLR5EddIrmUoXQhCD1LPikmcNt01CGuxJdPOUCyI3wmUHf0wtsavY
AoKL8yMxe/6isfa3CYoRulTO5BskZYCf9Q/2PBalZ1jwzTM+JvWx/IXN+g7yLNrt
1kDkN8f+TlEiAuX9JQ7qFfeHNtIRHM8zJlHzMzIMpdgT3S/OWF0AmbGeJNu6op2U
DkqpBD+shxJ86eE+ob57B6kLau+i1dIcTHopAuZ8vYkc8lf0DGxjzhxF6EMp7vZE
/1Gk+7X3F4GOrTAsDPIwtYsEqybesKb0w9DSMmNcqKTXG4I6hKgN67E+fXqT3sCG
ZjOCqp+x9OFpaUYVQRwh8w==
`protect END_PROTECTED
