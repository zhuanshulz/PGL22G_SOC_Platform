`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oH3gN7Nihy/vxkXeq7DWwhqmuWiZ0EWIrRlqvQ3mRbpc9TajmfQz3z3f/nbKzLkH
oru1VNR4Qje5qEUS+5/vaY1G9vFbI5ZD1NovHCsW1TPpN6HoMyJcB8W2S18V2MEe
RTPKwt0Dq4WU7mvo/TyNq4J6RiR9sjPBLjvd8SYZ3anf0nn05BNPyDQCHSIYKRwA
Q2QTkTABe9fbr5o1Q8FiPTarsFQRmYfZexMpAqH8ip72U/RWDroBV1VO7zbGgd6n
9G1UqouUg31qjfICvfR0SEhIm6xJojhs70dUiYOTl6rFiKrb1XsaQTP/Azu1WYlj
8aqyaEdz+3YYUll0xDd1fx17pXF7mZ7s8Q2ICzMmFikIhf3WcL6Ha19Uu1q3jlC5
x+k3k21IAZh+WcBrPpqPGW4Tr8HU5D8axF2IKpoK5wUTDDfBoPau3Yoa4D9iXl9H
3z1cLBYqI2lL3Qchg+y/l27Sl+7TeBUOw0ywGvfUF+9x6mZ72l6iexTrVamtVN8j
lw20BT5/XboxsJ+cytd5QqmPySFrEJGvt79+qE0tjezohASx+x9Oyr8/eEbWCH0v
HRGnUPb6/R+Tgyg8/dH2bSdGLCqTEZEj0QLoz2l4rH6m6D4m2wIGZIEIgInBH3z2
FvyWfqQbUnFv5tZE+jYx7hbj/f8uZt/Nha0+rodZYxULG3phrcF+C49EbN1aw1t9
`protect END_PROTECTED
