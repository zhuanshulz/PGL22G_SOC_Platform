`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hpCLc1S0cKjmm8cnPUr1oA9J0sRK2ne0IkcuXVnSzl1DGfGw6XP9ZinImY87PzJp
rlkEZPWftxRcw9rC/mGXm2pyCZOTHXSTSRSq7Gu2TYz1yy9zn5UUXWCjEFsLDZ/+
U7anTDb9arEAgnnjMIGaDb23P6IeqCTkglYGeIP3lxbPNrgncJr0vBsvfmmptgQF
MMcydGp8hgZPQQY860H5KERtGzHH3QAML5cJDON39Y/7V8DZjHArNzf7y8fSfRkY
jr63DOtV1o5iD1TIAkV+UV8nMbtQz0ML5YUGwGheL5beN2/EqwAFdrwg2NCsPyHV
rsS3qSkwQx2Tm0u9UUDSbZRdcV634wp+0h4J7Keqyjv3pImw1ckpF8eIsX7LVsHJ
ZobadyDFss1f1WREEeqWJ6MZsP1xvu+E4OcKzEy8c6XT4hiMqTQHJqYvOs19IPrw
16gxqdMvuZWEAbUVLixKkruNdD76KIpCwJjCOL/Mg92obOzxWk3ADi7bAk/J8VCk
vL3HKzVWVIpQU1wQuTAFDSgVXI4atsSBCPjTb2W+R7fpHTLORbInYhtaoysVR+7h
gA4pMBkLjgR1lr261S0ijVbGeeIhcf1p7t8/J19zmV6J/VVhf6hiqTzJZEie+WDE
conjZW5o6k8B70dBBKJijbVvTxmiBK7JIp7p087b7so=
`protect END_PROTECTED
