`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r+zm96FvhHdqNczOyyjYgAtfodXAfcE1JAVHhATEuUGWLPf5ChNqqm6t7H2/HQMV
TngYm2vFDgKxN8fZ6Cm0wcLIfbvnvRvTcX1HqAVshvrqbZswFdkGbskz6M8OkXUI
TJAS6+QzQsqXIPT6z8CFe5437I97n+fRzyzgxSLY1heQvoJ1TwCL2zGsGIfh4aUE
CjrwNjGprdpuQJGLdU9NHa0PMM2lgSlw/aWTWLZ6zHPiBnBbjgCelplWesYN9IvL
OpAyX8mLB9w88nynahPKW6eOXz2UomoBMMkpLX8dKPyiHvfOsjWeHU0RndmlByXX
1bL6KAQeP7AGdMl29nr3yhSOIWcpxzIpXNu2EjzxoHVAzGXC+IpdBSuR7nappkQn
`protect END_PROTECTED
