`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V4GXWdIZwfFPyCTXan6waYQn0QXHpwLn7D/FavceN5gajG5YKgL+7yVkJqguaYVk
De3OIdlc6L6+td2p6FBEaXP1OcclQdw5PMHvQcQJDMij6pg35jpJTnefn86k/OFH
FcN0Iuob12BDTbNDoBPIVLIXA0vGOQXg89pCzpSlxyPp1wYhuG/ur1aVK2906QHy
PWsDojpZRozB5Xrd97cQHZ/SF6vnO+mvLuOgJA18vbGz93Vrd2LSEPqz3nbOmuqN
fjat/jXc+QFDKaWpXtNc3t7JXriAk9UKBCFMnrq/nxyXLaOqgtotcOql2gzJbShn
If7VdM/2ji2UNvVrlkK5rKZOgg8ubDGhpWkBC/R+EeO6bhb5VXNNNPjvtAxXz7Be
iru3Q7/G33QZOS9DN496VWG8VEIEyFy3R6n3AkqUTvTuj8sTbOikOov8VtaUuTmE
JZIFGNCZSubay2iMFdt69Lfl8caswt5V/CrGe9VpFQNvu3NIMOmUqc6My3xJSJ47
nobuBLtox4ahRgmM8YehFX4SCtCQbMJMZ+GF6JvMRiBiDjuRFnh6ymAjXhElp1Z1
c6W0182g825M8qHqbEHjQcIt3jZ9fcrDMORQlttUCtuYzVRGlldrO3fnvVrXND36
zOkoE0BXcVKFZtYCNjDeAWKOEzFVvr9UgVWoAbAEIV3XEi81J2rOGnNDd9/KSH9p
gA1IVH71ixEK/UDVtUHgS0bwLS7e3YH95gHBj00yNehwB6AzNXbphfOMrQowmbnG
iEWV65+/cEVyWHi3ob/EgW/Qul3AhCQ+4h4QzeWQoNgesJz8/A8fWGUUwWVRtSYU
ADF1YqIflYelBmCsho7ZotyyF3E+fzwQuC6AFWRMNCawied4NOIjoc7IVLdUT/Wp
I9HQ6PDXhaMJEMpr6af7erqKjHF2IiYVxNhyb2IndX57bjV477W5mDG9LX4FgmGt
PUHcrhe7m5biK7n9yYnluS66qmLVQN0DmidN5y2Zo6OlzMys2KBOMYgKWqqGWB06
DLQLqDY4jx/ooFrExtE/an4733GGiFVRFxthIgtDY2TuI+qp0BHVJ9n4U/1wgKYj
RTqu3bqcqxyNHNpCE9YPL8mcGzpi4Pb8QvJFAsLc5f1KZtqkSRF11ZbI5fPpVgDM
Gd+LMNWUTiHTtngTmpBjxo/xs36iYFLAZH6fUMpfdc8Dmtg2tG02tAXqk/CNDmb6
gPrAWFE4Bmyq1C5bGH55Q8ufdFg/iqmE+cd3JKnatUyvTBWtjSn9dMYAcY/vXvOr
y+YRhI9NbS3E6JNmvw0wpxGZdnhyPfgGd/pIVjssNvjWZTFPGT9Z7bMj2v6EiLhr
TRCckrxMl/gao5jquPvfYeE9davcwRM3UcQwZ8R8iGdqrIayYQ/6WFRnUk7gvK6B
4DPZHRwz0sJk/IdJfPKscQ3B4hWaVFaEkk4Z947dg4rUjyPbzLW6tGg/9ntHb6oN
`protect END_PROTECTED
