`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HpGqD97up+FlP8nw/cWA6ALDTDx8kqY2yUDxZ6qtXA80KTb957Sh9MpvFHyOvW2D
qex9TYTVRXiYfaqxHONMLX4xJgx1qjyGXCUztjkNGkdBaya5U+xeGW4Qdiphlijw
ljK0JifVipde7tL/dJqUjATTlhliVGYCOd/+i+TwubIlWYf7/AYULIx59Vw9Vmx1
9LRTq5o/onLZ7m0yrZfapGXZfJzx6kOXzgM3zwCgGfddW1yEAQfauWePo8tlWX9p
LfSV5By8nbKzFhNPoAUJEMQ0ZmmVAjGrow4pP3/5Pz0Y4lfyeLus6s8liIcDJD8p
uf8r2u2G2h4QhXFHHKOuyuPRtZs3GFq7E1nWOmP7OlKeSgNTdNsxrw3+zZMAcuzh
qiyyi69JhSpFF9KUDgaavSL84OT5Rspnibo5EH6doCd8c+FSsbBCqAb2zbJyaU3V
d/BgQm0nBnFJco8pmomt0E0bkKj8Hj9LS8BLb2CM60zgKMGn2HlAohh9adUGGul/
gsir2FUKJLozMPcn6G8+yKYiyx76B0nudIPRRgv6P6/Itrc2HJV0xZaTZveTgWTV
uO/UnSfDpiZmbRTjQUB77OjZtMyNbDvMiaug5gdpEsb+LLDyO2tav0I8u3NeF3mV
D9dncJQYmAO5/C8yc34vzMWgSFPemQP2HmXmFf9BfjYXARy8JNdwBBGZLmiE6oB0
0vzbnu6p2KCOOLo87NHLDsOsFxB8rC2wT+awuU7VlsnlaWFP1tSBiJjJYrO14eFn
O50mwBeRFSSVvKoxYa3unjyHorStrc3Fz3KM7aib5taEGy8O7aFZbhI7niIY/eex
rr3x9HdyghnGINn66YVc/4mTUwrQbFawbzVTyme8eq7ukr6Tdc6/gCQDxoMkAQCD
kgYMg1SgEyy6DINqJtNYHqSf8MobF4gz793CcckCECF4utixZ4PfhttrJt346AhT
NMbCrJcXjm3wGes0LKCW9tpEGvlrnGGPw7DkHL+SlZ5CSWxwzJ70h2UW/02Ql5Qs
tJnnXd2egpSPh2oczHIfcFIf4nhT2z76IWfViTfuKSvhE3whHsR8ROeYAlrx4Q/T
h85WostGdhNSP8COhOv7NDk7xDhchy6P05m77bhJrwq+Ot1Zq1KAk+htK+QS38Hg
0nEDC39Ju5HvyJ+EJvptxnpmeb3ZpRTzjaJS2AwtD0lW5PDvNecYKRgbmwJBI9nQ
CwvHYn6oh35ADqiuJepARV+l/GWTj55tWCerBj2Mv/NlThSLKkus62ZW8PLCvk+3
vt8DYjP37uESMQGMQRXqckWBKjMsvBsDWkMpXhwDZIfYN8dcpKZPNTu8b+VoIHqM
62nMTcx9SGCBZ+eqp+lYnpoZworNmWyTL/YFDZd5Zb+UYk2S4xVgWSXqw+N/uR8d
2tX1P/bxrRoOP9Kxf238sCzmylxET55VADUAajUeBskiLx3SEkVhYOCGojMLNG9A
E4ssHNl5ja4qZynGuKJ801EL5768/MCzbB3C3//Km/RIDg+7oJvBnyT12ApikrcU
slGbhVpCJ23iRwT5/2/UMbXna9WbBXvyhtnJXvWBIB7vq3xByUyu/VMsriMdL/qK
qWTQ1h07GA6WYG3syuVfMrjliNVP+K/YTKTE2d3mRXSf2LZy6RoHReOrbYXgJzLI
oUTBmnBjAJRCpWjU6U6pFhsdRzZItY/IHXAKBarMfKfPIgchmNw0ITavQB+QiU5C
iQlhmhSMoe90hQY0kyGmLpJ6Fj5oDtCkNvQfOy3ffvkseS8SDvoA1AmJGzj1Itnt
`protect END_PROTECTED
