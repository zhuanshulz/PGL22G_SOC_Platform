`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xioPpVG/17574Pm6fnq4PY33aqw3An6Pn8RISpT+0BceRnqsOEQTqh0MGZA2P2pn
jhm7fv8l3jVo1wqZBEH/Ez3mWYppALmqImXZaVHrsZboENkOfdkegdncnkZquzIg
xYogMIW+BvGk1DnWxQoYyTfJzTtBV/ws59E/xcEXn0gJz99GXwplG9mpDwOvsFNt
yadjYGmC76pLbe1+s/vxRoJNxk8saLcreNF6/UH7f4+AoPdiweE+LfCy4OGcWoVc
ehC9fbkmhfowtLY/VpMgXqh+MMLPBGmTKN9hgyHUk+NL8SOUUORS5L1IMZtF1s/B
MhfWZrlC/IrglG33nr1QemfyzBkTpUiIbKtdFhXuyeo+UKe4rvDgQ8JsJpgZ97BJ
Oa6AAZkcqfgYODIxluxi1sA4+azSddiH2TQHVmrT+zCOXlgCmXXAwkVxnvMgBTQ8
RvZitPx8tUeiWo32iTo7bkmUj5bTq00Mt2Os7+GPQYuwQFdEwKaHG12IOzwnqZsT
Rz+sRn8RnaDaY4woTrQjx2MbdMZ9BR+Rlb4LNKc5sET2QfIrahvPBP4+hd9wdBL+
uuGnL2rKNDV3QOkMHVkCVkc9gaJyX5RKLP0Ua0lgOd4+xSU4i8MOq2bLynE1Jd3y
3eMepZw2WlH6pnGrCC+E3Hg0bPAllW2oDtK3sj1Aui4yckr3EgwrzaGie4t2Whay
SsM3GLN0pQ1fW1JR7A+/ZHs+2ZzK8nN7tN9Pk8eBMNWNT2175l/To8Jyvd2Dyrgj
O+kuS/W4XVo0BZ5LkcPLol/1mz8/OzdkGgeUFc4r9n5+24Jm/o4kWtamYf4FNVKJ
M7CSM1xVaXCAOqm/Kws1bdRJWxPn3UqgDXcbhsxZviZA94epP4M5ZW7KFJ/JqFYe
Q0/WGk5EA9FSZ4ylWrvV4O8esAzXBRw57C8ycZVj0hUqiY3AIqDr67V4kEv6/iQk
sO5F6v00kCVGyMqfha1gQw==
`protect END_PROTECTED
