`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0gWga42fspPcDbx8JiD3nJtLIyfdIyOdUFoNC3+oSF+6/BtFIH/gS8l4ydjjHn2f
o6CPcGoR5DTgkQDMhMM6jQ720Hr0i7Gw3sU3F80LJ+cCCXj8tzb2K3zM6bCH7B7V
39Aw0sUCYOZ1O/3m3UhT1AcBfeRAQaiPtyMOdUmZxy4LZJ+GjGsOAKRcDaJmfULf
F0/1WftgvTWhAWIPLTr5QktIAL2dsDGE1Ip5vm1ElatMO3xqsd+15Yj/fcKd+zn6
LJNYNy4vT2ebMNJm8oOZMNDvzSerZ6cl6QN5j/EL8ZGHoPPAW9w5IDanuXZJzPBU
vPBmgyxkHM9co7hgpHNTd1XGcNEleRGN2MxsAHcGRZLhFzQlOf1tyhhfZhWzBEXZ
G1TmOC+caw60qbLBY+yVg2q/2YLzapftQWeYiCVRBIsnp7kpm5dJRn1fodGdMM2s
PU1EvDOnSyPteAIlpIdMl0oiRqDS1CrWNARfniFt+haubRrOsKz9MSCkN/sqjMll
yM/b8msuwR8YHziKIw32ZqLyI13YG8M/r7XtTPzZ6wYvrkaqWWz9Swf9CI+gniyG
j718rZaKcbzlEaHTH4OsY806wqb69aOsNZ7lF/Fi/Li99HAMid8gaKfHahf/Egh8
wjIezAfllFJ5rDYx4heSLTOytgOS50EQ0/4ffC2XiZAWeVRazqVtaYFdqQycLnME
XOFP0RcW1bWEnNdQ6MICrCoSVJ1EfccRoqDx/V6jJsG5rbgr0Of6fbycVhfNQXCc
eFUt9id8BtM04dyfNnMOWgn5coo6Kpfm7f9kk9jyGLdEi+JW7+vWXzad2JhxTKgr
Rggo8Kpv7Fc4ZSN9Gu6L/OvRLUvmWU4pg2osv9kWIT2slsKtZfrhfh9Wn5vU6+HQ
8CSqBFdItCSk93dAlMmOMmcrl6EtUys8w9Vked2MhPJ1etv81pcKCMWdZNaQRl0K
Yz6wGr7LFCOORXUyKsirIx2xG4cg7hGCWzkf/rN0ktWC82C3sdguXllmfELW4kz1
o0O4VJr1bfM2L3FQXQoMQ81p10pOG2I+czbEIXessRVFZ7a+wg6yfodSgziabSVu
rwnqdG1oyenRHKhmdCXw9hiyoCaet4VEksRUZNWqr23A9g3OrqOFHPazc1mgywZ5
Q3f6uZy4P2K7bErlliW9goM/VovzjehNY+43GqW2mdeGnXheG6Bi2Z6PYxCY1CXs
`protect END_PROTECTED
