`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FIcVYxgog5zexm0v62r1zWOHubscjXJ/uB3IpWmg9mEtNEKUucvGGSkMKATkeb96
Xyg8ojnTvXsoW+WeQph1yFPq+n1GfuXMJnsYKMhmEN54ApS0OzZ+Ss6ZskNqRowG
UBHA5wpulYQj4BloEOoVAmDR84MFkaKCgbWg4wBKMfCVAJAF3HbqdLyzIPE81ejD
nRTjOelD6I9fbhNZu0fHHDYIytVt8RA++W8DgL+ejxFpV82ZUxZJslrtSzHWJ0lS
y8MEqTqnuIz/rh2FzUqHcw2AXui0Yd011RWnoiiat/sRVB0AGdlneBjMpXUAi2OA
f7WcjBWlC6fIUrlx2P7V9osQDPEMdo9UZeFVzCA1tYiw4uohKmdIMXmUyx1gG4gn
uKBObQ0JQiAkAxypCqGZSHGbdOePRDg3UrR+8C40eoLvhqebH82qd6TjS0O7C/3G
WOotkOi2ktO9rsypeZ/IHMlXMVUIb8Dan53BXRI2SieeZdSkQJEQhVmxkFo7jvI1
9dee3iHoSu+QqZC5rVSpz+O9aAi6Oy68j5x8PqpB2Gaj+vEHq3cKfeZhWwMZLLy4
3rYM37atJnjCYpvFazmB5OSvNEKdzwC95XXYfq1gQIEVKTXeDbE6YDTQGAmwqN+L
78YICqzyWM22Wr91xkm9R4sKhO2QRDCFRr7Av8YS5GV+ivaFx3WS2/xBhpAb+E6Z
XNMvMotjX6zN8qElQ7mDoB3IVWqFXkYK46d11nra8jL6QZCiaA4CnaSLE57rNSgU
zRizt1WaupNGg/zJ0aF42F2V7n0KePKTEy4W7lUzUG14Yysdpt/eOpukX2uzRjwY
xOupujsRcJJ1et2HyAMyPBbE6Do3RsoRSLgv3oaifXIKSR2RHr8Sh1RVSCm54Kjx
/9QcQRz2hBu7+ptsJMzngf0v3lI7DFlzcmuNG2Fo8R1AwWuzmmO58CxrdK0i36JF
UgOKH+fR7IkNXYl/jk2rM2jklsdph+zcmQZTBqEOxmn+AHPz9LLNiDziLoAVM6wC
jiGV+m56gulMfySl2bjOIev96hO7iNNgnYJHGyXEb5jaQ791x7HLJYXJbdlfIGnf
z+Xrpd7nBGakwn87d8TzACvnucmuHLSEtbz+2LY84cWUjkobL32nKmL8kI9jDNks
1gMFWSX0ZrCCw2sbI0O8XQ3hVea7f6Pe57fL1VQGpnH5oF1YiEXRBH+DmUYknQ2h
+DbXllZjGey8vEHHYWfdnPJe0hW0ab1QjZwdUZluqNiraDmRIpmBnBPC6QsugOxO
vaQibUNdV9Xeg4Orl/YDBrJVhz/WzDw1Sa4I/tkCdh+HocruDKd4aE8U7N/Yl6Ef
CcDeXcwfbRVL3y/9Rh6psiluUuMRwKs4GHs+xZuZmX4XMN8Wicma5BZA/Mym/G7L
DlvReFQaHxP0PGlTYKT68WfhzW4tbsd/6poaRFhXWL8ANniPWerQSyePFWE2+nIM
X+NrP/ZwpBy9nzqzpwN4w9bHfUjMRqvg/1QykFStJbZYnNUwgwosiXWUtuB5sWBw
uJEEb/4+dSBFUUcPNwMgsrqSzI26CrQi8x/ZM0j3GIKsbHU93MFG0aNztvj9kPr4
KMNEEWr6Ry8Y40K/avMPTG+S8LBmu44BGh4nWRhuYdp6MRlFbmNkJi6uDSEhPD1y
N5vW0V2y/fQQQiP3nfnr837YyEdMAuEiDJlQ1j84IhHQuJPE06XkbombSqd+qVCj
irofNa6yrgNshyed8l39EBEJ9ij4NsHTSYwjRHagebrHtTOWpmro9sg1Z3FJ32xh
ud7A6H+bRpXzT6e1s3bADbm+kZx9bs1wP+SRyuzlwGnOEjoaaTfT9PJlIY/wdGGL
4qVuSNMgjXBQTeYANEJOMUrcNEDcNhVN+OImkoIKO2hnQ23pJOKUkFI2qT4AWzca
a245n/z3+Bxx0DOZTHwgsM56hoPLnLlOPrSN5F3bYlR1RFuFTLv+BytFSM4D1bMv
ZhWe1t98hJ8/R9XmMJUGM+2dX/TCxQOwmwTiSblkw085rGFFswHMzOaSYO5PcgiH
dsCI+q1ue7ENIy+m1lwbVJHI+od93kJSqA7GgUb8eL/5FoutR2857d+5X8Pjfbry
83HtmN4ZEYfA72L9YfRvWMyJcJbYm0LaJ8ieobmI2jv+9t1qtXh1wzAh0oaP6DPi
WvRAzpcevqeYmqdIixwetPLPhMYVYpondV1lmAIHpChmwlPr3yL1O11XMXmlJg/+
JZww6rI55q2Vb4hM4c7AfEc1DnmpxGTZT9pSYzM+n0G5ZZTfh5fCe7iohj2bFAPE
5zlto9Arbr3mpcC+vpi8Lw2uL1zVFP2OR92bXrE1NdoIHotE3bC+rfl1Oq3khNsm
HGDo0T9t0XURihkYa0so/iwuRPp1Nqo6nlTo83LM3Dgdw9nnN+nKLgKFJfaCEzo8
X+UHiXVHA0xANvi0o5HYXZwlJiWR4V4zLGv8g3hfLfqMI50Fi3wV4YcBKW/vwr97
S+Czkqkye4a+/xEDA42eCCjgtiQuG3ahapppKUlfGSS9mpEaB6QkgCqWnj0VEnuw
AVhjFHmqOf8qj4/mSRJ6xY41PG6fPIhLfJ212o5ryA4TK2WPcfEWYG6x0kWvFovZ
FSdcnOwKbvIs17bpIXABgn+qFs9LlkkhGwT4SJ/yFWhglueaJf+Pc1p8mpjRWS+/
x+TLx673ZzLZh7+rL2bgFYYHAAuwTnBZs+pl/gkdiXlROJxL0NBCum1rWJaSUh0V
0LNcgJ/sPOFdhhTZG9XjPbHfjeLQa25aFcgq9QUoT2UtAfCJMAiCMF1XdKtF+JIE
G6PcNo7YcBX9AANHmMYJy0Nch8JCrrWbdY8VPaa7B+RSoHZqrstvgzODxAwjpSqV
OfHSW7vuyTFmRRkR6ilsi+R35GdAH++PUxik08gCshBjvieH6pYD4cVgzIKV61sV
zrc1Ad8AemdkhQW+vVkwVf5y1h0eMi9Or/QrjUmOoQaG5HXVZXFL7LVsYAKDk5SD
08HTFvJYy5Vn90jmoy1CbfMzTP272PBiXfEOE44ZukNHZvPWqIqrEtWpR1ObqUYv
KIwE6oiB4cVRMOON9YG4MYOjHRIezkPFCL7WhMHuiWFlegBvo8plcniph1S0fsye
jfMYAA4YPf0lgipVN0GFIaKkcdCHTgW0ZXn85jcD/8UsSxYi5wluxDaDalBdvJ3H
jxQSDoQLTeoR+G01Zh644x4veNWEKnNaLWUMyKfhM6MI23a0rzJVbFQm07h4gknf
mGe6mOAx5fVji4MpNT+3+JswQz32KOJfW9JoV5aWfjRIK1j7GvTNJi3FozvECfKQ
s6jb//QIi9hijP67UsVU/u9HBcrvKUk42w7Z+d0UyXNkC/jLZc5et0/mfjbW61lh
1pS0zcGxuooHICNV0Jzz7yfJLjgX6kt0zfjQp5RMR6TP+yBh+ADzyYpB0H+GpNGV
5mL4MRYP9H0B2jTsnFQfzXVdqtgRo6zo/zhoeSKNxx+2YJ1NXFeLi2fRZw2S46jR
obwz4Sl2O03aoZt8UNL14rKo27PBMEqhQKoWW5HafAwCE4utPHrdGrTqBk9fSD4H
myjDP6VmoKkDTXpIdxg96lIGAPgKhftpG9VAQMvCmreKjqMhn/WALqfnm/WoyUwP
pFWLSyT+R9PC1HIywigG3rhq7FnMcMl2BuCf/H/pm0IglPW/dT7Gkc0uEkTnPTqa
kUZK9FhzYLOD3NLnwanuLgCch5r+KGvtJ+DERoqNmyUr64visScH0W8Aobv/zy3d
OzltSGF/hcruq9DmZDzzgO4DFO0vKjrd6AVR42JAbLCb/PBPpvuZCz8ra6oFMKvx
gcDUR0AbTAtdFImfX7AlNYn7Gol1QVKRR3+2MXpigMFtJFT4E9nNmtdm/uZsmJh6
L1XsQRuCyhk5c7c1THA/g0PyVf1gdzNGp3JiHBSqNUZSQEURrbsnX61nTXZvLY10
pa0KHWJFsHhPe0n5gs8Yx/m9lZ4kqfW/DUsfbe94J7XJDESjl/PSEVqHu9w43JyS
XZ9A7VdXIWiWhQJ6Q+GW5yX6rHc/WjWW8GjdzCXhHnp+SB30h7dfUt19x6cH4Y5f
Y2fVyGJrhkD7td1giQpruN7k0FwO4NUeqRRnJ0iKVtRRK3r5qN/EUUREcd147PE5
ZsIze0OIgwZrqqL2rzJCHr53DJQqaQcgT76YCLuH3ocxJwWKa/lNK0S4ojmSqnA7
kv2mRPB0wivqMHRLxnKvUhGczDx7vdUx6hcn9Y32DDVt6gcso3MXzeGRTBA2LiYJ
vQCzaze/c7sP3hBADVoviDeGTsvImp8ouDZEbn7iGdVtWEkEnUFEpqm9Iokd/54d
kH/dazl85gunSM7J8F/vbCRWsShjCtaafXP2HkNFbkFmOOZ70a7yNwUCsXmhcOzo
UGc6S7DoWLjUiUciVLNRwwDxUQNUV9LAzLpEu/wN1kDe/81EdlZaIZk8wq8fkfXh
8xrs05eDGFfiYEtQS9+IFph8St25vhZrSEppZkPjUwRg0YeNLrD/iUqKhtjMYKBk
g5gtZPAIFQkg7k2rqtwoPZiHc+zlYwU1HTHroaNwi70Xzccv+MrZhly7db0mX38j
3dZThxvXLPSXssG/mGxz4GyEdbxR6ZFN2WKAq0re7jthjc0a8y35PV/P9A3fMSJV
jF9hnwR2y5MA2y/AbvOC28UtknGsslDvRR90fSIX4bfUIKRJ2Bl3nKTSj/Knr6Lt
PDbR7CxMR935hq/XWZMwznwXfhBMLMf8rcYf9yl6HUcwBg06FFG3TUKrEd7vZkFi
Hxy13aEiIpZ87cM7kDVEh1B0WCKLXGChMQgTDzZQAg7lZ5PIU8oXfyBGbQJW8S9A
Jm11KD1OuBqt94YuGYgxwl+Ljfmi/Rn3PzXeHUzpzndq91O720drUX3XPCLPIOOR
aKzysbZRwAY+0fvbRNo8cZVwhdKAx4/TcLHlyzvkS46uPL7bM7kd9Ca95sQJS6GT
up8UeLwTQ3f/joDhjE2K+qmM6gCCUWGdsEj5B8Snl5We26fCt0jQ3ggK0QrcFgGt
NcCWr0cpUjGAwc8g82QgA10a+5vKsMWGXvS4aFyIMs23fkUKOMt7RCW47ShUhvYC
26ai5G6gSkSH8hcTZ/Yxe1XC2+1cByFpXP+dU+DYK+D4ldCMRw8eQG1yyiafJNZA
1t2qD5IWYh8LB3vJrUKgH4eqJ5K2E1GYapD5FxTayEcydTruywVla1KIwBXNvMNk
wOKddYvZQeBhwVuCTNs/BZ0G5Q7/NgNCttWxoNAwW9BgNUAtaifj4HhDT+iIZr46
eDmPqQUaKMmM9EKZ86IoA7i6R8/3cD0xS6ZRFpKqOA4qr10WesffaQGvQED9CXnM
+C+GDhecdiNet8pr6QOMsJZz9KEHckr8JHK0cJbZavI29sSsprC/OrnTltbTlUbc
Na/q3nngvsbvzoo+hynMzC97O7+X21BflJav7Qw0bGl4lhzCz7eoaxMHbdoynPxk
QKVhO4Mry3tk5fv7YCuikadLr08K1R32A0DPw0061DqcXIMBOFzFrbxGHjqLVWr+
FZUDXGiLq+22ylVpefXO/06r4ZIpbgXV5qSLpE8CNb5GuLU4hpi8J5Iei8r/4YeV
qvjugSSJcgNRX8pHG5KzqqdlMPSe8+UznxY0C4Vr9MnRfhDEcZkQEmq+zAx9cbbA
CWzHRJdvxwxn3glfdy49fZnAuhX3/nRF5/G5I5b3y33cWWzsHeY6VgFzTEpTfpHM
EIu5zj9ZjMDIBAQqX3T3c+9NHml9PH2zodFFRM2GRxv4RWHc7EJYplfUITYer8ij
peUMXjaRbUwwbA2IMTpteWXVbEwRDlOJlmYpQs7W32D0Q8jjM6u3UJS1nSShjiBx
ot5QOeDawv+9wzuNBCB7uDPhE9zrn5xXE4lTMw44XAtIvxEozgs3TlWIv4IpjFdE
10YwSU/g30XhAfMibLpMp+yXCtwfgnC5ywzRaBdC1Ma41oXGyRr+z7586NFzFudM
P/mdmxTxr719gfIteiAODfDQa9q1xg0RgeFNVsI3GBrU4Yu3aPFBN2jDAttwDfFe
Wb0tvmuUEDImnydP6pZuibhWjoCT4ZVmmU3zZO9f0DMbmYuBTcNAgTgYSbxR0wfA
PUsisgbLj702QoUWpAGzBMVBZXBYhSyusc6B0YwCwEG+Cg4S4Si9jxmPFwxA1EC9
oiOVt4NNpZGsef76DfK8NxYJbED59Iv+MMO/WzBU6XHmO4MIsJinyuTJOa3fF4Cn
w2wX4+gpcDgpkp5LN/sMKTNyHNksAMm3bFCsQYl74RAC3BKhgomcYOms0JlulMQJ
FdR2j12asz1SJkLdhO8g5oBMJQV2Ld+ADisgMJGur5aL92Xf0zPVnBSQm+ngWkAc
Ys0ZecqMAbUmkcxgAH91cO2Prt+3xqHEJEFTfViWKux4hZ4kr6pkMblXOft5k/ue
eN4jNIKaOYiZAqRCl5llPTfc1ahCkqrkFGVPyO4oTbnvN9jfkCzVb38Si7617UuJ
IHzdfVYFEIrX6B6g8LAIHrhZAQOrDACYMXeRHCXVITIhQZlzKWBKYWMc+xpWTqDi
WfySfV5kwW1AkTicETIjAxwTXiPE+KtX894WGX2sENBnOX+ZW47Pe0Y9E8VqqXn6
pWEWwOO3YJilf1iOxZpa99hHKOzz1M5dxxJT81LAs7ZTVS2xjooX6kxwxa63GfMa
Nwki29zJyIapYXD7kqosCriD+A43HSqmLLc/V85sUJOPv/oVpF+6ZN6TgITJcc60
aZJmO77wOIKvZtdgNT39nVIH6sQ8NszuVYj+SmKYZNTdOdbzaAHecrEMCNKQpbpS
chhJ+5EjDqS7v/QpufL85iIqnIamxl6jw3ivuIwTRNCWorvw1w6VbTzOrluP1L/p
BlvjvdK3i0pez+D5e2IHNzrLZqTg3QZ9jZZBWrCdUsW0vHgrOJlVhJLA4g4qhRpv
M4eNSdAfRwyjSsGxok7D8MkFYr1JETep/BIo/of+eWisgj9JqUQc767VJenCRvql
UQcbAZ6SuQX8wokyRWgPkb5ZrFI+llYUM/gdI6E7Kr3XUN24JizeO1z8Dn10NRwk
hqwHeaibaJWCe5KBiqEVORyUVQAACV/zaR0rLKeRj+89d4Dgf+P3bdt2XNt0QlOW
aHCbfEeA1KhjdWHKQpz9jUAKvlZrAAP5pn+/2XTbarS6cpy1f0ZxZprTWdV7VoIw
W7/aI+jWpYNV8TniKeai4AfRlQThCL3Aj103B3mFFZBFdli5GO/fJJ30/bMR3JEW
h7+5ZuBjFIpUrYZXxNHFu7ijMi/Zkhy3uz+eNdgydAUHgy+6AAYc32MBxJP4UaJA
ivIpOmjO1+Q+fC9iZJ2+28+12UEYSjFLyZYcsRiChhZhYdE+iz8A7/UxUWWuv1+y
RXCkf0IDjPotzcoMoyMe73f0l4J7MDzYF15mwZzHaYlwVgFx+Y/4loD9Wu0ZuQvG
ByIjOdn7jaSyl/s9nLgnDgelJNnRDvOEI9QTqOwqGS2hgkvBnzg9AecXTc/dKzX1
+PALgg9bn8VLUS33vDnTLeHWoznLBUguOrfJGFEZy9ziIp7PStxMlooUfcLbWn1M
Cy0L690Js0kydh4+RZF2m4JqfGRemrXGbO6/+dL1T16mAPBpAMJS7K75nnBh2O1W
3cQIvtDwInWO6r6fyEbnioR2TZHqdJUxo1B9iTzZIMyWHioTPPStxFvlq+VyW2Aw
zOgORlNyp9my8iF8wd/MLh2wCKDLAdQP360SxqI5wAz73biTy2iDODSnBxMQnFrr
pcFzR3Q/k7F7hebNTPxUjMooy8NthnGGgAoFkyLD98CvblyHf/hBgSkqnEo4MApw
2HtFnpwT7nqlBxam5vWgrhjWH/o8QEGW2qdvyH3xwVSA2x5BlKgJSLQFKswD8sS2
zKJP5kFdI/Td125onmVIAf43D8PG5hJz+0BLO+AizbbhOnwp5j/rQgYGZ02+BJ4E
f9gnWp4dyDgM7F3OodL8VZYXDJuGCch+HND23Dm4v4pOmEAMEvccuYl0Tsws59Ub
Zaar57um5azK0ulBaLUYShqRyekHCOKJgqQYM7SQ/+E0H8ZqwHlTcl8P1hgr9NRE
HENnqfLtU2mFU9caHJIWyu7orcHNAIhzU869JpCFrwmCUG7kVeqLal1dXYx03AwX
Av+DwL4hTQSQDzGAPQ4kwDRSPxBC9gAMZY1eVDrvMJ/tyZ6sEIfB4NPJ+FJnKuc4
wrpTZRhwat5pFKTsOB+61x4+tpw9wz5epm3RMEBws7cPpz5f0SfUohvFSEHou9Ge
B7MsKyvOmsk0oZ2wIbhbxx/YM6QQ+rBqeRGqT8sXkDSCdt+XYu9o+FvMvSmq1Bu2
RrL9PDddaF1tz9wqultR/oXzILTOr0+u5uytdEX16NOt21A4pUoy9pXND2pYRMFV
qW2qkiaWxwU+uJkjIrCn3KaB5HBJjErzdY+p/e5XEJ1ZGrknnf2DsYNtEpAsTwge
`protect END_PROTECTED
