`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/a707QjXIqlsrAhCxv4lD4fIxqloHpv4vIySmYnHEGVowrBrCUt8U5CwtAK3Ebqe
RvSU+mxQD5T1jtnGIKtDI/c5mBtn7tnP5b+YBUklfft6Q643q6B4pyxmpiOiPEna
VYB0xZcSbtoXa9I0U6W2Shl3nJx4iwIrDyjCsUF3Q5gRxgty+BYRQnJiIpTyDr7i
f8daAKlXZgxJ2KlRBUa/BtzBs+ZOcRVcELUasWtSZUPLOA0S9QmVprkEWVv03lP7
96mkOBAAAS7i5r4K2+TUaJtjF0RHR6IrQ/iMUp6PgZA5iP8bwaBKss3oEk8gVtab
jXVvl6jR52HyAhId66ERlBgcSVw3LPt6bpV5K6Pofm83hRTsIn3mbW5a4DRPO7a5
`protect END_PROTECTED
