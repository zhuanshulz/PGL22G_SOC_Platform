`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EcX4TrDkhVvvlgmAoBJtwd7OT9uzRcaz4450nXIi2HlzXDB8tS22+SOB6C9OKsV1
Mt80KhuLPxrEgWOrWwVyQBkabuxMQ20TQoO1u2q9aKQYzXxInpYNJM7PBbmdG4yp
zscZu+0+pATB0/Hu8SzEuGbdgQ2k47yR0nZcB9eKCUZnWJriGSPtjz9uriNVCFZZ
jjUtNHLfQuPYekMW3MgstgfWNlHFUd0Py6/ldzRdtS0v/12fkvVqWMyiJf3tLJzM
J8tw7KyvKFpvrFS0uf3IG0jb+YEiVkehDVJKeKdYHWO6QDVnanRyqcbGwsvqYhjA
2NWA9GZyUCm0z+Sj3/nny0eh9z/CURmyqSu8cI1ACK3joH+rIl7IO7XmUQ6/2/s0
4PN0l9RLusJRST5RjZq36S6CYz1gknldzICOP+XN50wyhr7hbrwhOHjyw14CARCH
cJO6MX3+ah2KoUPk9ddrDmmdVZVFHaRmGZ8FnX+QznWkubDWA7C22xdYsbVM/SKC
1fEf/FpLdpF4CVuGhf0/fHfyY09t+4/BI62lo47Lv/2jd+Pi32eYJGs4r6Hg7Oqj
LEu6eSNNVEa2oJjAOkwG8qWNwhPoZd0GZSuvtc0clxmRVlxpUNQMvsY1cPmd6ihJ
xMsaW02IgOnPUZihqlnQZAgfSq+C7MRsdfHNRet1vAQy4U3cQ99hTzM4uykbr5a+
AfaZG4A+fCRRTJoPZG6jw1QwZSMai4mCqJFptCNmvqjvTd5E6Y5NiTiFLpkeKrUS
VqkiyfPJgpT2pooMXnqQ23pGHcj0xv1HVmfR0Ke449iXBwafTQWkocEEghFkjzem
9sJKazy6pYOjTI3naCpC9KjzxYYS7R5588m9HG1aTibP3TpKmCDksomxwhXNHUgI
oV0/BkKnY5Z8EUK+jG7ljViTT9ctOWG8Mi5nQQRD1+U=
`protect END_PROTECTED
