`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DLK8jzn2Qxr//g318nxVZn5Tq4RKiGxcCiARk9h0tMxVH/zy5RVC54H7yWrcR4PS
vAd+hUc/oTXZh7nNPSVgqFS7+HeBJBfsWuBxx+YRWZNlCWprhry/l6+1N+E8JNs0
YRyphvBy2QmDYLPYSHjjc9YcyWdmdrKMuWg64opLbPft/Le04ZRY8coPgtSMEaep
f0AyRw8S+xmuMPPcyw5jtrfU9R508kT8k3sZfplGuBNQR8fKwbIteVf0n1ZPl4fu
yQ4jVNBmxzyzbA+LNa2u6/S5XUIRYRyzeIjQBG6Um/eN665p65tgXNUSgKnYlutB
tWV8F31/uwQz3GQ7DcRHVU0kuRWpCihWJdtv8bhlzZiKmiZYRInRF3BUlNGCTQ2E
NQ1Z7xdpgZuIFvCmaS4HTH7O7HHvc1JOHg7BCyYpioituRBX6t/OuqkRSBC7jntv
DvpNszL88tMWU8wIfi+TB1B5cIsAC3dtOSmcFOrgu+ulwbe4RRRaxH3nKFxyVC9I
ABA+XGpQahPiLDb2oAOfPOAR24BDffjGfgoztufhWrk=
`protect END_PROTECTED
