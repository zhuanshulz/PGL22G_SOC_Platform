`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wGy+cybVsNED1BDqYA5XrfUgjBSTeaZD7v0ci6rMeYg5ZjXh1kSMXe/1qP6vuM3J
wmqeYlUQD/cJS+o+34oA2D7h914eumIW5nn/xGTXhMqBkLbHVIPDu2p5ElhL+ynG
QuzmXSk2+DvvOkhTxbvhKruraDA01wDu2PFeEQbzGRLoVzfk1VX6qBS8ik0wmta7
qXSfAHd4YWmUEnPfs0T6NBpwi+N3slb5vKrHD30894PzU+Ev2rdP7bWDAGRtPjEv
D+LjbIU5SjkQ6q2bLhEJSslsYdKvcGnRL2Og6wodg+J3aYe168ZdNt19alACjcjr
`protect END_PROTECTED
