`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LkDc/EYEjlyuWwQq0Bv+qN1n9uu8TH+zXgVXiu3MTIdFiyvuzU28Dc6UhfimM83c
vRfMbVtizG5INnUh8fxxPNXTUkQHwoSKabLwYK7xv7443MSGUfC2H7ZVhjwaW5iP
YbHeFa/82E+G9mCSM7vwuuT8buUcWuwubtIxDWGBtlqbmwvWSTDdQxqWJvCBzrdc
CKqaQe8odpZ0MR+9a431stBG6aZPcXYcN+8xKfElEoStMPinTvc3lG+84jqo6LRb
sNUYWpuSk4u+GRi3AxOr4nCPHHJhdZkJmgMvhR8DGKv+jv+jrGXqzzbjmzOVq4Go
zzSKZ0Tw5O2zCZMT6GLBihBbSt5XKgxcHA4O9thiVZksne+p3OZuuVTPYg9Y5rex
dBhKEfN/QKuqDRvXPHWebEBWo6Xga5R0My5zC8fLdsu+EzAV5qYVHXn7mRnbIQ0Y
KXZ1wyMZCOijL5i9QX5IPMO/Epl9CZBWy69VqEntERX2qQygZR7Dq9vtPlMJWY2W
eR+dVnyr1TH2xJAqDX6gfAsFgGy+h0qoknLs++tMIPPQmC+xD3uXyA9XW2qjRytN
HYPp1fBS0zgWT57n3sZ0q19xILfQ3ymjOhzk+HYp9nrW66tyE/7vIH0YN6ek/YFt
YdHo7ZBXESiPcQ/UM379CXV4zq270Jxt5jadZ0YKN2UzwlT2iGj5PqUgBZB8PON8
SK2DtXeFO6zLxCqeLoAFTsCF2/IN2El9Xni4E7lqrT9A5TfIvfikdtJVj1QPOa03
qriRu3b4HDg44svjx7ro5HWpna9gz1wctidy4SYSC5z0XCUaaz/IJwVc3oUHJH6n
oJvY3sz1RWNihmcsRetJZUI5+lExEmrskuxrZmiUZTHmg9eJK58bWx/lWdZ3/8Ud
`protect END_PROTECTED
