`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tCXHi5uddffOOBJ8XyrK7cVmMcqCVpIIiURmlVciQ70LGQCXitOfr2PBdG251BGc
N1FdZfj3brBeOQhVvf43qAW8Jj3tr57SumYAbKkREoTrYf3L5Zj+5JYOiW/Wv9C1
LsleQEBhPaVdqVpDdmav6w02N/oLwuZvSAg2wXvcA3oS/8mq130zFMyd6RVAmER1
bT2YzUoC96pZkR08ngArqcfmzvvIV4MaT8tNe/iwbgnDJApzyltz4daogDdcG8mC
`protect END_PROTECTED
