`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vtZfTsbLB4F7c6n2hAJyk+T1Z6gpA5uNyVamAGG9PSfHTHb4Jpekd8FuTumeUBme
qzQW3SPrLGSjHmAVdpIHHy4kWN+T0xgtbKjcpE9L+fhA4/d/JXHLAIo8iJ3aYOfb
ZMx7HVi6Z6PWnUdsFjGgEfbOPEEU7LRKjqpcFA9nwb/JsJvAVhvp2JRioJKn3VIA
s659AFz+QV/Cb6AmAuWseXlJkSosNqGBqMp/oWx4VUpKW3Lwy2bBpkx1/7F2XxfS
qS+K4LuLOk9zYV8yA4fFvRrq+LeRrruAOtIhUhXyAPOwE1M3+ufjOa8tk4EGEQ+e
jxLuPtUWgUZLfCd0BPcBcugR5MzncbP9gvlEORKbXDapslp2fE6p12vwb9wRXUzx
ngXoVdu0f+WvO7lrp1bGdedxoL7OR+49x3ciIMCg3voXlSlyFolYxWc2D8XHRG+b
EZF/GxXHYWgWCzITbpDiH1rx3MqRHvCh2DYCkIKdqewMssP5u/SnYPNrUo5WjQrj
Qxf6rTUZS2xqZPzvltK3GxOxce/Ao53YZki03ihezDqn3d/xp2x2jqTqO8EdEPpe
2w6MGX0QZaGL3pd54v8mR0cVgc6seolCMmzTNrnRV0Z1eABoag4vRRGTwDKa6vWg
3LHX0Ip09EKlRgCGSKSL06YnTEuvSwLOqIGDy0XuAeL89P0e0YUP4VCWBIvyWqyl
6+fTh7WZDJiEKmMeUA4UZ9J4cFl9rWVfvgHxFAvBuwk0rJjvSP1JCm7CtTgD9oL6
9RCY3DtLNrqzuH60+G/hi1er0ZpEH/bsupx8M93EpY2v/iPxbSIzOmiOmtYHM3e0
NA6Qj2sdNyN4p89aoACR8jFFoctxozuGDuXyMQRCUtbDAzS/9WzSHByzL8YkCIYy
qMDAtfLPck36bnGQy709YyIW9uz4R+/kgICDXJ9CchkPrgJ+hIgShV6qM66on1LD
yMfVjIpRv2sfqC9wy1FfMandNED1zhXN73Nmlk4hb1cTXUc5uKwfX7wCyZFAiTK8
feJ+Z/oViXgTVocPiRLY5oBrTmlmLHIOAbfuhKNksleJ7bZXq2XN196VZbJIufqH
q2zHHJkeB6HqAPRW79w3Bhv9Mh80dz9EQDlDI3ZGbqoXUoZzq1lwkm3PSOoy+oKF
nlxyzrr9L7o89Olt2AzWTebEOoepWexq5a1UvkzpcSRoDvrhONGNTpKdvGqGGmOx
IYHzLwbvTl3HJchOs/V/sj5TscIZhiqj/EQO+j3OglRrRloELwy836UN8vi/Q5Ym
/hf2mHW3oxUU7mtL0cZf4EQz/LfAz7aaGq+J3JGE9f1/HhXVUewCcvbaGoHQRHDS
LnghH5qg+G8ODDNtGwokFy4DmtudYd5Ms6/tILG9NUzdWQmUE0FJr4ZflUSaJf12
k9ASXG3MsiR1sfTzZlXXaXvp1Mjw+sVZ/9mOW+achgEBn93WudG4Wdi1epdiHvjU
wTj52kMZN7hpF0AjcMxJEBdi35w7E6BI0Hrf6aIDuUM7jVoekmbLOaFlaV8XtGaw
1sA+Ri3Fe5Z85RxPi10en7tegBz/MBCer76ru8v7/VQU2ICRbbUaaAKmcZMpmGqf
60dcBFSjnXc0/n0W1nAFapbZus8xCVYSWV7cUfGiPtkg+s7Fywa44L4sLN2+acGC
BHjNW3CbRI+3Dqr6zawvYaV4Q4IMZRa0fFOn6sJRPVQrrplXSGKUp9AUYh9LLRUk
6Thu27YmXd3VuoOkA+IkewcFfSX9hM4maCY5MrpjK5J00WX51ecLemONY31+pIWi
DNF/iExiaEeAXUHvTF62HQ/dI3OpPm+VlwzR1Sg9/zeSrJS5UrWcOldh/fRhYVJv
XmSsjN36GIvVlxwovvKGInPoyRYOYxw8hJx1sFFAS1E=
`protect END_PROTECTED
