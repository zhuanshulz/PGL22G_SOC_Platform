`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YipRuDtnA+a33li9MKPFqOJ2ISwyIFwcfwf/aVVjBkLISWmuQsvS+ozc+dL+Ou0W
UqvoKfdSsFblT7xlP69ILNJYHSWuLKjMxqzwofP5jx/LwHDnbO8SsFfuwKy+gs8U
izcMW2k0f6XAqh5u8TgILaPv0oQXdtVmUct0ahjqu5PMTvtsWnRke/1MFpc/QTEZ
GEg9ThYBk3/t5Rl+LAOQX3J7lOLPGiegVuQ8JtZrwwQDmRN1U2vvA73SYBM0DU3h
15gXhq0TYFsF2tSmGI50leWRqfH65azcPjKgqvtAl0amxw1Vg6kugEa4h4GXTMYG
IGfSeN8pyJJlOHa4TxqmHbeWc6y0G3+ww4D4voB/gOO6++XfesnvpjgUzT1713fg
y70WXp7jT5DAAmIxO2IFY45se+HRb3q27p8vjE8Up7K8RnMG2+0M41Tjz901Tvcw
1R2zTq9xFUFYHnzt+V2loRokv5MVwn0V0VMGpMp/0nMPgnTr2VXyUY6K02H5ARWX
iXDQXUJEOVX2y/45BrynSleWqYSSAQA4sQzwvMmmGQTNdECAjYUsyzwZXbgzvDEW
PDMD49nTihoRaDXPa9epv+Fulbxfsm31TCCMA7Nr0DhiQah6XcOiIR0BCP52SDeC
E76Y6MjHoHnL34mqLD0iIp+kYlzsFjPdTVJfeF0ajWalqY+X+FKjBTVuslnMtxxl
6TCVL9cbA6aA7NdrfyqkSziLRd5Arn3PbLQQYMs9YcpmhLOmcl4GO2SLJpZskTMR
qrltibGtKIMIxaXNbXbOKex31juiH/2nMgrT6bfmHwM8Au06Laq4hqzljlKsm52h
57LBQEHIExb1hfEtZe7jXQu/bpUiaPYjt1KoMJPb8ijVjS03nwqezvGulT1TOu+H
vJTjRfKlQwlE0vx7QWzLTZ+/GxakYMpKDgoxdcn738kAYvcMVNJe1tSQgFEhDMgK
BEseYKCG6g8+LIx5LcliSw==
`protect END_PROTECTED
