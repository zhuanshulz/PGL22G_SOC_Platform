`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EXb3Kd2ZFh24cLOP+kGBKxbYrp9NT3eXkQ0PKTQ73F9kWen7lDFowrF9L/JPalNm
kslpoI7IP/rczaySbiJn4yhx6ycvtag3W9jnfJvfN1z0/ZdLNbIHUh53HCb2y6Os
avJcHdVbzWba9rVeGSE3RE3+Ju7ZNHga5nE9Iq1iDY5Y4mRoIsCCXxzfP3dGGOEW
ug3f1+20jQIOijb4MbSXFmBJ056dFN1Rp0POHJ3x3Y2c61yDt+xfZzL4ftZNIQe/
d+aefQDf+I5pkpslpPe5sRzTteBouImqlS/wP16IMZG3OCW3F+1IKsPGyhi/xjla
59CUHDPK0a4WijBWi5pWjkWnQLfitdjF+3ZnDOURNRhB7TQ2WKbj695XJsUX2JgW
KawqowIV49wbK/USSetou0ScHMvxNQDl58OcBV51DWe1ZLXqXNIligs2l9LpjpI9
OfaBK6ykOnrSHmJPuHnvk7cZLoUJCGJ3gxugdruBAgF9Zb5EpwZJ1Ngv69SXGPdo
5pHBiakwO/dVj1N9JS7ZVX/KXOM0iiZg5GEiFaNtouNpIzkzYuEBivGfBhDDcHg7
/wXKJGEUfCDzRcUK2OV2SFotED4F4V1KNTjHBpP3PBqG2kJCa8MQZu3Iwwq4EfCE
qwv8Ypb+iolBUKTOsnJZXGDXkLDWS99SO9sNtChTa3Tj6+31WEczXnhs1X2Kof6t
IJuav1P7fK3+Q88PUwXR7OmALAlw1+xHgRCmjv9rkOSYCjVc73t6/WmCoOeGWOMM
+tK6pCt8OZIXQNNM98b3iep9xpfWPGKC6QM4b3zkrN6edZfAY6Q0U1i4sE2g9VEJ
euPlad6a/RuZr2vRnIErgwIsRjGeq0hPp6z2lBMnI5843Duv54H3YoTLfcm0wAD+
1PIXdRgejSGY9JOwts+cYJ91y5aTAIkVM8gJ+4cSf/WBsEtAwE4ZPIdZ+x18sxZF
kswhBzOySfRmLLZYZLWEm/w2nw7lYbx2pj1enREa5l9ZHzb0BCCn2TqOn9440J+K
nRbcZnE0I8kxvuekaHeNcJsqmAWTK8JBQM4S5tkZmN81uiju3fmbSaz2HM+pl7y0
w6ncFiVbNty9K6B6zJjO0eeuMYPFANVPIzzlGMv9zsNTltzUcCDs3abb3Xo0m24r
OWn1SCk3caLqIftFioflFQ8xo2vgcIWzV3c3nGBiPY2r4db8mf4eoFbMLBNcL335
4hHO/w2OdN3L95iB7ymWFSa05czdr1IRwrqCP11lHrwFU4xNzKoJiVVZF7ybalEb
PmCj/gbDk+ENXbCbGblQRt09IRSRTFYycRFjO3gjA3TWLN3SPHzcAGQSGfLv04gh
II3D9Qae/heE0781BXBb2KAmRurmMlr8Q/T86srvq5hRUVgb674nQ3lPvlR9yc5e
Y64CY+Jgshc6sU93AeiRDeock3aWt6DEA7N1uHHNKW8GjX79UcAxYOKzNYbE/0Wr
refwH2cwxHZ5UQxIGB824LgVXbvXNSyDxM6f+ErOIsAMG2Ro7izt8Y3aWxnMvflJ
ppm6iBhWGhW96Ygy4W8rSjRFkyr/zWHV7yAxuW6ne3sJm58/Z7XQWwlKKiAfKAfk
hKTouwJqprupHVpgwr4ZGNPGcwr8ybfaK+/zxk72K5dbQ9G1Qa9LYoHd06kltBuf
cm7uYwM7C0xHtpvBzV3t35b29silZLdVBKnDPb5ZqTCamgRwUjrTr2YHG3RGOglw
WoiQm4VSdTOKswtznqdbRhTNj6Vewsn0ZcTA2K7klilNvALfK5CfIzA/IGDwfN8T
ErZj7B9rp3ppnlOK9Zbu0B7uMl7ZtV4YwYXUQj4kbTbvakjWFe99VOR1OsYXhowj
om5wqGRWVuW+a1y1UpT00uSRU9B8O9pbw24XsP7WuNczPfkrLGvJo24IczzUa1nX
3PoE5aKk0jFn6rMpN1QK21j6zomi0TW98Y6PY3aYC2i8x9RQKl5RpES16N5ItlRd
zSOOHR/01fNQjDdZyY3FiC0Jll0eQzOrgTh5ayABLZYG5c67zZ7x5WNLO76jswZT
6xJg6gixB9kxMqunrM2J7lIy8qFbs71xWCMKWUkRFpooLuGStAxBuE90EZu5cLuk
j1lGcP3Hjqnez1bIEPbJ18BEPulcOHFp100ZB0sh28M8vLIslxhfKOz4pnyCB+ri
p4Dc5FR8mxl6awYjKdAC1MkWtO4NQSB4nEQixwAdS653d7ZLGj9B8FQMHIQoqH3Z
/KP+KX+aVGKqasRNhcoqfzyenY0OTJ77Y8qVuE1cXLdgmXW2bxMk3DW4AjkM2lBQ
WiFzErdbS9JhpwHpipbURzbswRk7mDGRbRE2hZ3E4fwNZ4ZznrCvqcHIF7Rs7Qwo
yqXX+7FXklhcoebBnl2czk9ZbpoMVgIf8rEOZS8OoDEIZ6FFcuxWUHYYUZq95VHi
Ayv7tdlMhn5GtLw4hfGxaUHhzyrgxZzWfG3tGKHDU4vxiILRA4afvjaMLbGZZZDd
2qcqvaZ2paisjKgeT66nUF4UJ42gvr59wKl68HIRmuVBmgp9gEjziVr+9PMFoDbx
Gs2CmnJ24q41fK/ezCa6g9xCXlUdeixspik2p/WvltYGftv1m6K3sxa14qM+elfp
3KOUQj4Uh4GwWIOBS08R1HT/RFPzvCDSxWTk3jeILW8muRK3KTz2/r3zbULhfGaH
j1DSH2dU2mcZ2AxIQyDqrx44Wuxl7Eg3jNme8nY/TS3YldXDOeARx1/f2JXzIajY
oPKmxKRjq3d01TX3wf4cjSto/fYQ19mjBN3G9AciYcr7USfNIhoY89LGSPyJQXmB
ZjiV+DeuK+BJHnclGqAkKEN2XCErS9OWSGEs0FuqjafTCyZ3X2RClvIxE9jejqX8
q8ooZ70fcip4UulNZs9Bv820GJAIR0ojgD31ZExQ8CcUt6jX4WJQKE+MiE6h1T3g
05G9usW9qoPxObduXobNV6wEj2qI6e/VaCHto5VcqixWbdkR5Tpo1Heqn5qRm2MC
jG8j65wz+VxXSUDvx6ihDM62TkhaWmI8Rc4UO5LyA/r3siPNg0w7osFooaDfQ4+M
BSE9AV/Pi3+jLF8UTe2keQUY8AMIpflZf29U+FS2WB66ulN4tT9RnWfODTDwptlv
INWtO2e6EfcXM2tUqBakeCFby88qaVeTdSjlKPm5AVtuX4ps6CSiBMFwa3SB1+iG
7ZpA05fUUbdybEP5j4drZfgKkjPF9EPm5aLTiomdE2wbtglc5vgutPvgSwD95yHA
RXbL5DI1DV+RqB3jDxNCyZJGzSb7/thZrM229c+wV0W2hX6pG21mGf/4CBDunogg
T/j3qbEYBnTsnfloge73JuNM2fdY0nJo/ihnjpOkFNpTWDs2nU2PzSJxGQ23M5Dr
9S/d7X9BTjxVwEO1HgIgHfmskCNO12qJFE1kyUQhJ8lRuchzJKJpEMAAEIepiMpc
yaL3kmA4PVCowgC/yo+Isj0S9DO+yWuHRywpRVTD9yn8tQWXrY2sMMhSr62mdy6T
DJr08IzKuH3qsW2wBYL3GQHtMM/LBgKJyF5rj58QIjZ909DUL+iE8BKmvZhzKAwq
9EA23twBLJ8IOlzcZogCkeL/NnOmH84+0gCfiXL5E8Lk+3w5fHIC7/NyjN4TBbqc
l9xLp4Un/+nyANfcHCrEgnc82E7vTGLnf0MVYM+lPF9KgnPHmiGF7vppZpNyYg6u
ldk9s9BMH+7GMbVRJ/CBa7dUWn9Q1GLKMoetlrerCWy4quN1oauLnSgEoq/xzKyD
5Hw/bVKrubKkg+kKNvr/eTJ2hC9k9vud/x4d/BFd97YrOxM1aQUFkkywOKxIJ/iM
sYVWy0DxNuuh7nmpHv4mxAAWZFye41qjk0VkMi8Y3jKQtg5xsLDxBqzcD9TIczXj
dSAViZp6XSdVkz0GtDGZKLLPqQzqe9o2K8n/TBQpB0WBsVWEHB8BQIk1uppzeogA
15yS5xpAj1sXOu+sWjo/YYcGlJyBjzim2wSQhHUMxcMr8i+k6VQj1k0PishOi997
3hgZQD66d3bPh2yPtWEeYaOSZrrtaZRcZEPxJbr+0E1idSmDmRf5VjHEaoRhyDzE
QWLr3Lnso2OuzN4UDSa1ygJ8HdxhyzVTZdPxyH4KENE3vdXN24MjWmFGZa9uajZC
jLcIJoqI6ce7RVCaadO7Ihkn77sdVcwu9fLC/rxz1wXt7BSF/vwdCq81hLrzeBmU
HMXE9VlFP3oTmjImekkQNCgzT78aYkVYgaahIqGO9aHDXucnB+2qG9wEFJ8/qUsO
B1p1vpuSMP3x2b2+W+HnLrjMJf/utMB6cDZnUSB02kLz5N1uOyLLbkK/HuDN4zkM
Zyh5Bi/l5ftWCRb+5eCcy7K+Z/ocrTmZcWsuJZxxu8Q+t4lMwqvKzszhIh18vO2e
O7YTdi5aW7EF6mYXpxKDHgSg7/E1G6TM5Mt2tKcAiCK4d1tAsl3bQjBKVLDXzuHk
nxbwqsEap5x1Toa6IRjgG0AQDD1v3R3uEq9B2qBzFpRV4UUBJI01zpUvuxLffCLW
PrCINS38YWEYQOidB+iX3MEUFvLnkAf5QUoySV5DGjSz39rhwF4m1nIu3UYa1bzt
imOCQD+NKpbPluBSYaQ3D/0UKvxirWRUxzahGwKt31uNwDG/fX35H8Gp5z3ucQ6T
8/Qr/zKV+Zw9bx5y6Hr736brxD3Qs0bltgGD7txypoQ7IJ56BiKv7igVFOfQU5QF
qpPROT639CK+4YcFCxXntm10LtfxKgvksHCvXIETE4zIPXVRd/fps45Zkcofn0V6
l9HQSG8U9FfkzttSvVURMrXyGlOMS2Q3WmYX8YgazpXhVByOV9/xqHUiQ1dtIY5/
fr/xsCsLQLM9rQtE1fXIyEKOtJo4tCdWVSUCxjOgldAoO38wbCQ+k4eAV5xRP6Mv
ZTANNneB7Hdq2IQdIq73zcdwH26+O4zKdzHWeUgt2ObxwCgbSaKBtvxUDrZxykaI
r1gT/g8DAHYG9i05yNb8fptfmX94IFew8QfIHwnPARrYq+K6sHbkRlv8LrBa/kZn
4LCLXMxSuRYvdp6EJBJqQBWKpjHuR6NRDRMxi1FawwXSbjEMZ8wf6zbwwFDnYZ3w
Ub1wIY0i7125DM7SwdK5sjM3jU8r7GYwdKDXnr/SMKjYXsQovYMR2uCPJxSiOkGJ
jmpvdFPd2v6CpzRCKZTLlhPyjWqQdp7RY4yMuhtI+pQnLc9AunBtM4V2cYllL3VW
C1NlJ5EVEKW8LcUyRHmCKQiBDwU//565St/hDN2jW7e/2YzD6Olxh65wDJeJlG2n
0cdDtZXpMj/pTAgWSCExbRKRsxBKJB954RJiX3gogoRRWFtCkgcPEdxeKLEYhThA
gdqT+zl6oSB5LB2mF0BMPl/pBcSULN+YYDrpsmYqxYkH19jz1lMKJso6WUk87CFk
PljTCLXbdss7ZZGyKbdOGNIwqUYWhcUpmOQnSooaB2d1cHNsUGZAOgVxiIFQ3fpf
EVX5vSZldgGeAkWlxseygbtNw7h/IIApJj8zn2/eFMIHToH8OFwZebY1LyCKFmIk
cCsKHNwccn5614SrnRdeKHvHdn0cVa6oVCdHEQvrIdHGbWinO9yc7yB1hJAXoa0T
Eeg28T+pt6JLlSUPkMReasMi/qGaskxtyoFLTs88p56EQCRfLuaWYw4TZztL4zf3
jO58Gr8sHKUwihznjgbdjqkx+RDhr1wRhXv4md7bC8FHPd1Btu5E24qO56xStpgT
Kp52j87qTrFzEHK75m0XGNOlR8gI8bguAXu96ISV2nj8Kb30TcxsabKJP1CJeJ28
FP66MmtpI+y/10NrRlGrVnlvPeTjsWp6Mr8J/W+362TNYhU9jdLLrEszk958RH7m
0MT3mR68MWlGKgpcq9PHSxafO3KoywHh6pkmJuz7G7Qz97gEdiijAz+gWMwG5o+i
5uS88BRaegI24mVT9hZUxNgWngF2CYn+k5KwEPwBJpnOydyLOZJU03osyIvvHF1i
T6s4sztFAGr8Vf4geV70uX8jd24FLb+lceb9+Kbrv9s27YTgHxXZXdOYdY3cak3+
rhtWRTERQRz2NogGrS4B74oycDgrhEfag72sP2CrpEQdIh5hkwlHYjhNHbaAsSzw
h3nM1CMb3I/6Ys0ryQx3eCSofHH8c83BHA0ybBIOHPZaTsbUJ1j+wCtHrAf4QeCf
XHfmBCM4HnmD0dSBhTMrzQSZPMTLRnvqoZaKXypE/7bUHhhP9m7DQflS2abjFAPZ
LkUko0EFGhf5Rus8tP2UsvNGbwcZIsb0MrXPoiOwZzLoEcGcJYqWDXIQXO8gP/N4
QvIRpEmQku0KmKj877baWp138rQMXTtCW8+UK8alB81zpXA4Aiph8z3JBG3payRL
WfJ7o3mZC5O+lfRHtQtaFEniznrbc17SBIiZnh7vb5DCozLOv85507MuuPAOqNpy
d+ma/DQImaCAZh2WxHeap3NhI+q61CwupuGuyzpyRo8PEYXa3XieS8DT1eY0Zy2I
TU9lfBKHetYrgYK2pqZ5VwaGV+33O8KTW4MXeBZ8lkFv02WJnUoKNzB35PLiR5yi
Jl8ErZlpVo/osYT5DnZn6XQh0d6hiX2hmc2cnAU3Ch0zqnEZbq97a0nIrmp0H196
n0p29jxQ/aoxNs6gS+Ris3IFAa97VhTdNEUwdEMTClrNwXkmsxxZ7kN/rI7d6OqM
zX6X/jpQtNCxqg4sN1Ejg52kep5quy0mxeloLTlI166QThkCDLCX1bsC7uCnwsq1
6Lm3dm6eKeHWrApamX53vi91aNWPb/qjC6sCIHxx9sW8FC2M2602Q3Tvfl0i59pC
uAuqojxPkjpS/joU/M6IC8MDW+I4mG6385ml86EJDk8iSU3emLpFfyI+LGn991wi
ICz4grGqpo3r4SP3LpnYNw==
`protect END_PROTECTED
