`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XFgyH7iDXpecgAfbjklBvPmaok+HkGsgighEbDQfF63mSKcu38pHiHtDKTdj5KS0
99ZYEyaqTk5bGJlaitVtwd+EWqJTGaCNVSim/darS5o/OaxKJZ62BkGJGIqDOHys
wTrp+wiEkbTyhCq7EBtrmttRLr8IUfLN6IU9N5g4sX5YgeYDiYW9teXNmF61L47Y
TVOwLhgFA+WO5zVTPx+7Qv5xxR2SfdBaUaXUHjWejPrd+XHH4XgMS+kjwn5gxeRH
iHyVXONpzsjitCRhvGXHB6BBxT8F0Ip9AkVod9m8/GVpk7dh23N7877tnw4KT0xr
+A5LuDhdxAyNKOxcVlztlYbIwRU09B0ZukWaJqFQ9OpvEXl0/xklj6nasdnjd55n
kDnNR4n4Y9LqCBwBjMvWm3p4C7ZvNjeyLc0c1vhTulgKcxpWPcNMXpOJh6EWUqVj
V3JgYsoyc63IQo6qipEExkhEtIn9Nvs1AuTLEPvFZufOsG+Knxit5DKrKr7An5VQ
wRRZw9SeulxmlYPrv6wMw3wIHyhcuMmcb8odN0lI4m0Sx9NC5YoLy1pxBt5RdNFO
uKQqXQ7XeiclkYhfZ2bvQTZrM5A0B5+FiQEIV/FJi0SUwRocERvDSn8u5LVHEPxW
M0BMeepp8oLgd3YS8OBBMccrU2+Ee5jRT7TOGxEoMLqUIFmsgMCVmQI0Em2yamJ8
n+fe3FYZJviiJsetYtwpIBeSY+LROb5s/cYPrgt6FrSyB9nwARA5RYSNLnXOhWvr
TIhXl6W57wpDprAwEKv3md3RwuNHzLMOYp09P8GvdXERTc9dFUXjFeuozfZTbfdR
rN0igWjvoRxI9UeT4M4gFxA2x8xI7d3RfiqGSe4Axu9aD4nTCAFcl0O7S2zX42bE
RkVoUU3NfZkdfJ/l1kEr5KbVxWOx54un7hIDx1iaVJr1Si/PC99UuYXnGZJxM4mS
MNUuNkTlGK6kXno1nW6ytTyph9gdBYDXsDBw9Z1CwEnCVMZat2Rp11qKefUekvvB
Xd0vZjsHvsQ+CkrgWtbF3tNPbdHrVwBPbpm9sl3VonE0EVH0NekXFLDPFtZJN7FM
OuRNN7l32sSLlNLmGb8/t11+5lfiwJzqnKUld9Jo/I0rMm94DIsgYEpgwCTsPGGz
vPpTZPo4Mud9DqNy7NpH53J7YOTIySZ1l2LOEQ+/72v33cCVG+zVr1dyrGz6xCeg
CIu8kFpVKqiBmpJgsiJ6Y+xh/kaFXIQ5/VzwAif1kzorq92YOLiSNXVuQflo8Ca6
YlvBMh7gwO10Sp8OpETpdN5HOjgklFovhbFf9vol44zDYn+27BAXrtUGiMAwG5tq
UOtTnmUIQ/3R6i3/vDqzjPx3yg8yJ92r8eXE3lHDt+YlLxdWLMFItrCqQXa4K1FC
lYBd9ylkcz0WWMhY1Y7oagXB3g0n3/hNdd77SeZwNyGUAhS/PU7dB5zjOW2t5Lwz
7I7lHhC7t8AaHqgeE1riNRf/iGB6Ogb802vf72OdIYqK8Jvsff1IQJFGgr+svFo0
tMnKzcf+LRKbiIuSbO+1iX9kxQ4Qb9DTwW5SSZE4zUcGcgyhc4IMcV7Cdw4IiIR8
cis4YsqEOHbVbgeXTauRHQ3a6/lcsw5H97J6VLZgGr9jRbSRCUV2KrEJSWaQY2B2
IIKVQ99bsLSOhll6EmALbRXopJ4GbVnLQZB7Bd+jmLAcYSAy7gC/8h6lMVPALTvP
vzWaM3jEaJ1vYanixHLreEEFVa7k63XxI8EvZX/Bv53G+1jJgehGoBEHybg2bGAi
xEsfmFBJpufLkUcYB9Gbz9usCFrtmcPNtAdXDgkkOWVDmmIGghnkFOintc+tkjQN
`protect END_PROTECTED
