`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kHQTcwb+MOYobfdFj0Wx5Bu+0xq8co7B7vzz0jGLSefhQiEgNm/z2/W+/MRtJxaN
p0Xtj888m5OyzSpNQ/PDTFWUwmLsBiw/zNj9idhvCGBuBSWxRp4peSqhy2FytMQ6
wWbZCTrIEMa9teAmIwtA96Pf8SY6O2C20i+Zw9tMekeJtV72ac8/Drfvfhec2evg
oBoBkxntjatJaQY6ygzZdX1c6bHzGAzy5zjJmaD4J0UmlxLD08Bf0+WJRcoK1KxW
VyFyd/neA5E0qBwTUXQpkwb+pjxkrsOWSbCUt2jJaX73XA4EKU8wZGiCbS5irb9R
2rImZNFkbMjLVeFdlSglmwZqHdzPzHfMj/40AsJfVUw=
`protect END_PROTECTED
