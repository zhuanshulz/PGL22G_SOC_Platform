`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v1UpLuDH4jUIDavKgf8QBlxm4gGBReBTe0nSMaCkFYeMipMN92sgugTik9pbDpcD
icDlwyAmZMwAM0QwuVB448SGJPJHZheqdEREMVROFWBeEyuQ/d5t7nyXvnl44p7d
DghLxCUPzUHRPr8LS/GFPJqTeX2X0a2fL84NXx3sGNIX4a+XhM/N9azC6u8Pfpt2
ZinfUAOmaPW+zAWMfpLgQB+UO4Aj7k0GuHK4OdT7JoYovpG5bs+xBMtizdUk0O1X
TTPkrAKI9p9mrB0KaxGm6sTWHaIbo3/2ssfpBbUYgcNw63yQ8IzxXZezhnoKbQ0L
Rupp2beiQNBfFuOCchHpBPBg8TxS6LOPeh98+TuNC4+3dbR4BMnlNYu46VRqRTVc
w4mW73lwa7bcgVfAWb9gMjuN2WDlf7hPSfh97XFk/uiJskYAotOjo2yfNCxWKrRq
EkGxPQyTsrL5Z5/CiGBcQ5REqjmEX0vh3jDb79x/u6Px0kipboZfalWeUzVBGAfj
yvGJRdSYFNcYWJgOxi6KHPJ0IA1kc0SAmNBpllwfS+VYS2H67Q5cf+I1dHD29alX
TUchUdN7FW1CIv+83kNdTkpfyGl9lO/Dp2LrPgJQxk6sdEtLXEz50tIpmPJWAvNI
+ggYjpB55Mt/A41lOvq5huQ1WuK0tPDpDcGqkICeffzxwApbHXcH7XF1A5Yyr505
jzZUCwCklnkOtieWAlnnmgFiJutn5pZ2DSRBY6WJnjpAQVaorOMRw3abMho0NHuo
5CapVQwcEi+HRvGtlHZH3YJW3c5qHxl4cklrf9dSYdmrB9XBvj7YSU6R8Unk5iXD
MWcvg322x6RI2AUJJrvho9hSnjAxagaoVQ7myZY/0Uljg0+61VuuvS/8CNDSHJLs
jgUc9Zy64zAxDdlfdSULZHDiwNFf27octp+X+Jey9C6YnlFWCdINpvXhhkSVrF6f
w2IKaCoCvYP/14XfjAW+5I66VNFb1bAfUezB/XmPaWs954Ptgap0MNNA6I67Wicj
oRDu8zBcwJ9I8XtzS9LRKGiLCcd9kfXYdgJDIbxugAdk619WH6LC5YYbFI54vuVc
V0P5gJlC4eO8bpGM09WgHWYFoEli/OnApscZjwlohbRBnHXXepqokrVCtYQlb84I
1kyB7kngxMxQaMrOqxVhWNPe3dFX3R/jwnBOsube1F9rD9lWdTyW7JUFbh8Oh/N0
s+LloSqkB7v0yS4AWSJP1Qou0jvYVDSXj7DYek0Xg79dfRKDAK28MgAGm8JsPRcy
0JS9y5ZpJSOuuOeygqNvm5i0CHjvCuDUyRIs+f2fscw6UwpLnM4VUye9Y4145tSs
WDaSaTnXFnq81SQK+FtdO9OKTBXyDGpT4aislUg5a8rHimzSmDczYcDOfphV7/gE
VCfGa1wWBOZKGulhXzYm7FCScoFhDPjnMPTRM/5kwb68Yvlv2OZtjwaWEm4yQCr2
1E7lfG2v+lB2bFhizFJWCNEQkTaxk1BMb4uDhuOSjQi11TE+d7OOwCwTPCdOIeUp
GbjYGeVGu001UDqiCvIYuAGsFXlzm/ByQ+Mx8VNM7DcbggEFqZzlrZL/2yudcbZs
vZcIC/EjTd+O1z8QHwll+HTlsUHglnpB4EZpsWICCeLXir2MvIKIme/iNNyy+xqf
vKMiV9r7y7zR41hqbyc1QrWLlqje4n+U7oclS494xsNCMeYOc6xsojKuxkE1c55s
E5sBJVLCgJn39DndJf9FSxtEt/MY+qrdXjEfkGmw7uEz1HzboedBYWRsbbKyN/Ih
pQNs/8x/Z+kbXGgdFXbPBtHt9CnBYWrueg/dF2r9RDTXU50Zn87wXcDDnjbgcaga
Ta7ueu17V/+8uiRPHkeyx70OUGJ/fKBP1tfbTrvobo8IhCNxDVIm0alctKR1bTQo
f9onRJJHAE5T8DMHD923nIvfgLFpgX7tIryQZPlDAeroxyAEwfWBz7l9XzzhaAw7
ycRwvfB3wsQIlXfXnr9QZYE2FAXBbkUvrn06r6cfhTUJnVjzOV3GQ931K674dqR2
o8utuC3/hGjRYvK2LMeA6KeOyDAAg/3yklTkYdPhmVtEHe+/3VMPC6v1vdBKpXrO
CO4d0mhHJpE8RSDNZL5dEj9/moeoppRrQsFymnWhOVwXQjbOwKn3LDkIMmrl59+9
Fy9wjzn7WmqqoAgwLXuxYsGQB/uHN2NI9Cwu3g5rHv99NUfOeYRetncu2S8ouM7f
jZ6Icb93KX4fYhknJvUWLvwaSIE4S2xZpXzSC0MqemA=
`protect END_PROTECTED
