`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XTUctboD99U813vNSsV37qI5CsNtxfr2s6HgXwMsG+x6MSXNu5xmotDhRdEaf8SB
zgLIN4T1aO4STz/Z+WAyV/gl1GFMMBELJB9pacs9g2Z2BJipNhkgE+fkVQgAOmJq
rr7vlDnzp/1FsOE7ThltpWnOp4HPHXye/uNMe4ZCL4QJgHlhnc5WKYG1uQSVLHsr
Zh6tbBDYpR1GYg8MrJO+5ijg8vCCB0syXdHHjUzmKJL+deu5t4gdm6l1q7qekE/Y
xCWR5/g4BGa1qaQo8aOlFQEnWUrl4YrzZ3M3c5vkbJo4PimuwW1MMSpuaznQDyPs
6ucHpQnE7gjbe0Jiq8ChqW4q5mqp0ntiBbLIBe1P00xeUXN6iP8bGAJkmUzUUetG
KWGZoGdSAOGAHu+UU28L/QqCJKPx5d3Fav4rT9buxb29iCWGssKzicqM/qLmElIs
PCZwhMH2+321QarBz3U8dh3xDNmUFfi21wAzgq4OTpv/fO6hhvjr+un5Ykd9yJLq
Ac+u+sR+JCcSyPwdlwfLgGSq1sg2oeuzXXxx7qYCLQPOwmC/WbYEUf+1YeFT5odf
rlO9WL/BvJI97K5fohWTIs65g3KspZMx31eLo1h0rX8f+0xBDZLRul8M94foH3ar
+2tfIVCr7TAG33GeGEMQmUzsJqN8oAGgWUDOHt14PF4wpkLwdWLTcz+T4PtUqd0W
ftt2TOwYIT5RQeH+NXWxsc49N9SBdsjKk+is46gVCLjYTe/l0jyHEGV7ylN9WlJb
XhCTTEYD1q8e6JCHmrn17BnsoPKJYdabYZznX2I+Hu7ccv+BGddReyuwdsfOjQqG
qSDqTx2ZIhbT2s0FFGN7tvqW5XjNJduDq4a4H2YZqdItr9i4YomcBHVjud4ezaFC
7osF16o1qv5VTQwUsQLpFDG4G/JqX6BlDvSUqJ1ier4ti81in3z/17LZAz686Xq8
lFlRsgsA64pI98ZBACBnUxgaLwTpRSoxs6hCMy7JEd3+gjmTy5H39lINIp8FdL58
wI+l2Eyl8jSqHGw8UMfLqgERRmiht3dmMUXzHOFF/MLoroJ1aL1bbsKlOjZiBrRH
ugsi6F76OGRNwPRqnbBgOF9bjtaB6NK443O6LJhlO42t/8qmHeTlYwcwrWu4E1Iv
OC8op7YPHXUcP6Tvd1Lk/TFV9Fl/tkgIllHJvMSsv0CQRsoCJQ8I0JJ9ZVbfpATH
+lcMugLLupCopSjAzAUpi/mGgjAtH3DSL0EPajuo2mE6udoXdaxS3cwt1wEYGi6c
/0mgFfXUiORd6sOQvJ/ecN7/m42rnogx8XoAbzRc0jKAZHc6XEmeC7+Y7D1zxCQz
CFj7wF0LRvDSA3ZADWVPczx4W1TBgDJgUnX9edse+Qll+gBX8TlWKBym0XsbIUNo
CRIQmhmhnpR29jtR3bkh49GtK4sO+sTomHfpNpNww2qxDCn6/zEOhZ8Eu0qmoDF0
xKs+ZGrWj7lofB2nvx09DvhA/sfjMmLXaMWkLerulsfKSBa/dyDdQDRsRD4uwCSq
Hhaz4KPOdo1Qwg/cCuytWso+Z0EIN4oEVlwzqqHDDj3/+y+xNpB+bDfCgOJRGunk
GnfwTUIgSyFE1XOi/A0/fJMYWGbE3nEa6HutJuX56Ve6ccW+2YKss7emZg1qCTWT
Ay0iv7E5l3CRZMEeNSd0HCQBHvgsXRCD5DT4L52G7okXH3QDli/mwwPPJJb3Lg3K
LOFQRAre7qAQhW0EwigCcJGcnVn6Uwe8AaNElRukAnYfpinqIZiqqZIo+S4jm5Jm
cbNvDYJl+/jm++V3XYt/EBYqdhga0I77IyZYIC73bPFISl9FD2xRAgJsxPG503VR
1Tt4yT0k4Zb6uXwJ9uehkXeBNfcCDJ0fpYCc3iFRxVwIh2VYSEPyA1mVh+59WyGa
xJzYaJWtY9v4Aed3DWcE3p1sDn4GHpXR6m1vEJUBRk8PzpXcBYhjVCTSEg6w9/Yw
2cKxOgYoZhLWLKz3G9JX9wcnoThxRfGjYCFJl6oVzxSqS/Z8lI4PiP/gm1hw+k7T
ngEHcBrjTXCMcymSNJejPapjEoiR0EpBarGEjqn87sbUvZvawMItvshu0A+hv3XT
2e6d4+VwgmKMaE86K+31Aewj7kyf+7Jai0AVMJva57VvubimglzSkTVdkJ+qUbNz
RrTLA8BqWbFdK7zLpr4ggO0KQTVXrknmigfkuTfbpdsLmjwIpkv4DrEuHQ3KE3rS
oimO+mN+OFrS54fK5TDAej7bDFMqRjhOgJvhLbphvdP/nYxnTQtC1OK9FZXI+aRP
nQXNIFgUcWDu59Z+4NP4jQ/s2c5TGsIHv1B4MyPpRBD7sAzthkd29gz+S7tGeew7
ZiOFtgI0Ko4IPQ095KBBLKg7UY260gtXKR+OBK2krNxFoZRninNkV5awIWrikmfe
CVDBb8J3keFJc6iCwX8P+rinOChJcsnQu6L4EdPb3fLu3VlL+KzrRSrKo4XlgKfj
oi2A/OLudjDkXl2IfurO+5QmgrcZb/xxriUcQE9AKbvIfU/G+E0epw/OqDrhvu4p
G6pFIwd2mVNI5XAe1lQB2O9F44Lzp1nl5nC87LH8441ORV84XqXWCtOSyF1fdaEL
zO9QMR6+o4mQbehnuY2Ep93Nf/OKX+dIgi3n+uV2HUUhLX8LG+HX+sdEEgXF/Mvc
JVpjE3XqLVBfMjYF8VfLUT6A3AMmhZA1UxsL9dJpCrfhyJOHSFYi1NEWkORZ2ywA
KcUtQL9QHmTX5Ot7p9ZhS/Iq0pCNTu+tjREwuhQ9aJ06G3/ZnpR78Xo74zzf27IA
7VBRAD2gpscJ2H7xJ9aVbskPIXqYJT1dW1qXoVC+cQLv5t62k8A3ut33fU3s13iY
gKd2CoBgLWSNGKY0OFhlC+DWbNBOTSxKbxGNA84wfXh+vmiur0dq38EfO975rWVU
0yRw4j1zlkM4x4E8mOymJKOId+IBNFyFSQRMMdCWADtkNDqeUdLrDEbY0BJLIUvg
LgUdTYthPm5mokvCxXkmwzGRF5LkpM/RrYx98fEIUIlYfFyL+j2lSakEw0yjkwWe
bNLXlAV+p/2814+R0gniv6p9iTqolo0CJUcy70axYWRUAX0O4h9pZO+6+f0Tohsl
ndTfd/oJoEJJ7aOnXaIlQ2EgEEkcrnMz2hx9X4kvtEQTWkL/AIRAmzmAcFqsrN5m
Z7iR1DAqtRyreMqkdHUJH48FhED0G8K41ECdPmzT6iSmqqjXa+qHtnffG9yJ4QGq
wsXzUzfoULTnoaobV/mALVuHlmI1HgGZNwiTSZwfzyi5e1GDeYZbMitwmwy7ScSM
OQtFXGjD4fYCL5Dp+BvlEvyVaOM39/Mec8MB81nGy+NvAuwiTdb3us1KgZ5vlt31
7ndBF8nTGIIb98m7FGaF54HuBRkb8AGKa2Ep30IOd/9q3oDTDrxoUcA/8Ezr6eZ/
daodkQlO7tRnzCiAPyCX3b0P0dHFbd6WiTsB+jIDa5GPqp844Ef+E/dEioVth4Jk
vLZJ26f7SstEhwFuHsgfhJzRWWtAzbG1nT1ak6xQsGYM0uZuB/C3dcnmNt15C1z1
mMTIEhr9o+YYFDAIpMlD7GEroy6sonj5jJTFdDjbK1VUHwWsvPNV9ZK5NIwKzq7G
M0vti1pqbVshELfHG0josj2a9wsXL5iWN4hxXa4F6czfiLiW+cglx/9Xj6oDrLbl
u2iZAcj3afyGbcu30uiR9043i5gzLwT0Q2WqbunoLxbUBKJ3cruvsIpDmoxLkW/x
A7mPQJHKe9mIAM8f4vHAYxQS41OokBr26j0QpQOiGE80qQsRD9Z7GEDz55Ynt5FN
96ym3bnF1IRB2/mEu7Yg1hpbC9aB14p9OPjjbnjPZiXlC/OsXNd9FlL78sdShvQX
PBuhEsPST885AHeDfF0+vpA0VsgojBaER9hog/lyafsBLgqR9M+euA61SmO1JcY4
SEAGKfqxjtHPKPkYSliokXpBW1Dwi+Dm9W2DmhqXwbrcV3z8OdwmLP3fnV4FztJl
4BZ2IARU8T075VPcGVfyj1QYbBM8pP81eaXt9wA3mPGxsgXM17Q9oB+/W9bFN4Vf
rIDHRmN7SyzDz09v4KSoeR7pkmNyFnGSRw/HjnmsdwYgnmy6J7knFacWPi/Hub8+
y+qUJybLqRYoWkh4D5lLQqEZxg26UdVzSspcFMc+4G//RZFbz9TQVVf57u5XPH/x
k/T0//distc/3HivCzu20MZXwr3ihcrkkTncz6mRYCQ9xm5wYlbS2pkUYbNPfsio
j5fDGt7y6uzl/JlHjVerbrUX+jWKQoXJ7GcnHacZC/aBNyX56gXDxzMKQRtl+3QQ
dhF6Zo8bIGJWPZjAMJ0YjMij0L8BmjDD4zx09QgzFcJvzBNDjllw7Y/XN7oI2ktg
C+arNFsiMMs0D++VlHULxCtMU58EAWCTr9fWVxZ2mKDdq3piewWqY04SjnrfA3m4
kTkcO6UC/LvL2nMNgrcUtNmGH8fGa/WUbgoTRpKyCAc8cuuW6HzfZOa1cnowkJlU
RUEhQ0znUtkO/cZw6CA8+haGCLtC2nwS47MwTxIrESDgWjsOARGVJ1aGswtpfSnZ
SdMvDCtA6RLIaMVSFs6aPuPKk2RVCfWcDOZqifLyDdvVMlvbct3JbSsxfDb+ZbVR
`protect END_PROTECTED
