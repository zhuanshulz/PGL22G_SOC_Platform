`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1TNhKOxa1ta07G78RE4mIoNo0kAPPvDkBPC/lVOkHfAVJJ66jr+k37i6noDBgX36
sDDa+QyeMv9DkeebcXbdf6NvTcjDIwdlqeu1m/y2g5uggEmMQEXr73EbZy5xF3Pe
X33LvUNGqTordUjJY/dyScr3I1m+eJyMVyEchHCVj2tBbZVT1AEUHLT86SLFMqhn
6c012h82QtCldFgJCdyj9ghdKCdpRcObYuUjXnSj4GA7ES6QfPrujBL+Aaz1FknD
qKWihA0l1F4JzU0oi2fUE22K0QcRGEES9SBrYrJGTv3cOaPwh1nV9CpQQZ9Gk+pn
amxiUjK2eACbzvM+hv0KeET12GLXNniLf4JGASqdaPrj+Km7eYutCURALxvzOfo2
XpDK8dI0RkD1to9gwp9YmiMx138yMyNNPyB5yglKWnZIe7+ovviepT78LKjgTQp3
xunKtkhV7hJnW+OKK4RwwEhdFlvk/++RbIQuE4pTwLe1fVw2OKBEOUNo8n7t9mEu
SadwmOAHrkT1P6uKw6Rvr74jb4/QBHT8AEWpdSiUHid7SjZ//Ih3dKA46Keu/9LJ
a+ZmdBEkzfyfEbRZe2wDzw/Ra/5edXVjk/bAenZX9GKgCdfBXR2KkZhOP4YXQneW
6gR7yR7hNu31sxOzWGzEtQ==
`protect END_PROTECTED
