`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BbuKD/idaFt4p81hDPZ/XMgzHxIVZVy15BBAfGH627iKxDKN4CdmcCJynJ649yi9
+KR6ZOR6QMBdvlOpp6QYaNPilqiudpeZVVOgWdzfx7jFmjY6zkpQgUBtdcEmCXyZ
oXpI6eL+RjO1AhHVXNVWMaZv3aee9G7Pu8q+CvQ4Eqs9iKiZjCAlW6Gp99wDw8dn
A3qgTxIT5mJaFiSLQ6hPhe6lFx5fiXJH32KPwSo1vc0ArhgWJaJw63K2eAPUEoKS
UPkeLmNqZCqjzIPVKoaEFMhmLENLSnLnCLSYIo2TvNU55gcuYOqgC2Jdt50L062V
hzmPHVS7hRqGTT1yG2afYuVieitd4mkNGdX5TO1k0iBUxIRULW3h8NM7gZzPZXFT
jTrhrdVl7LYHNrohU8wCIFFeMpuuHgfbBktQB0Wn6dyOU64jttXJm3zYVCsjAMuk
xSj80dFvsILhXRTkUHK91RE1Z8D7vBliPARgsgK9Uf6pWZkXyLc8CDEF9liPnt5D
RzzJ5h3uo48MRwPes43LoeVuY8sBve4nPq3i4PYS8wlTCpgTsAwUQOi7NuGSs+Z1
`protect END_PROTECTED
