`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EVtpF+3qfngYSoGRbrPuWXRt5+FT152oE+bbBh5Cabgpf1lhnyvy1FYS8/4o+FzW
O2behMtmxGII1J5P1cWrFAEft9HD8mSCbeOgcNykNbi3E/4TVWjlEoVsqII/BVsB
SEAiYY6OvLeWa8x3hlxl85TAj1ehmPe9n6lSutnu53/s2Ucfs1niqs9TONduEkmO
RGaverSpD2BeORSsX2md7lbj02mXg9xG1lwrHZ11lKAv4gvm92QvtkiNtT2D/gkq
BCLf3dIJ2U3SeJgWbHQu4y8lC6+G4cL2ZL/zlNx518KW4b+k0K9XJ0gLs/wcCMcE
uS1APowtVqP1uhP3lUMDFpbx9HpPpNcnKixKIuZ3xSZXHD8Y4G7O/3V3ryDzzGzT
UatnpquzqBfvJjvddtki3RaP0w3lpf8RYSIMnsS1HHeR0llLIsEg8NABFRaS9lDf
QlhFgMJOYuuRRZiEG2RWy0Q2C10Wao/bESkxRmOAyMVA2yilIIG/HzZRhx5iRrpt
7/k67wBmIv7tjIBCwXYSxiLe1joNJBWirdq9tHWzKJ6HcHlIRlTUJPB23n2yk18s
dUOJiLMTvjoCqhdx/BSeEP59p/ClyDrGsPh8e+vXaS5Aq/doS5ptfI7yt4A+MKJ0
8ePXDhC25s19kFswaAXTu5tp58f9G4EevP0sl4rbu2fLpL9IZUKseymDsYxnZ8ys
Xa0IcaHb8seE/ewPqHnEgZ3qTZekx7Ot+rbAHCTs1GlFGVgSfCKXlVJ7qKX517R9
80ErKIddktCjT0favlWL8sDKGmo7A5ys4e6qT9VXTYPDARZPrdxPp9xMTkKIycLs
MkcZNbbVPecWJQw7bwXP/Y5Pn5ycXpa7uiO6eSDgg118oaQ4Vm8ZaERcwK3dESg4
DhB5HJXSkBvTnnT8CjvAVHZdNjJQB7TvbSpus/zAUu6WaWlODRKNk9q+Lqu7kWp4
JA0NEqOOYlLW4spfYrntBZ2AOcNJ7u3Gcx/mXkz5mFUDBxe8I3dNvoHUjc2ZCr1v
I34AAE1ZRM02bI7JBzlmfunQj9vagfkK2FEf0nP+FsthSrAMP1yAoxHTgMyQZfLj
OSFwOQR9jcJ8LhHjgAnsmUUZvhcax+I1QjNrXymuc4Wpm+RlpENtAVQZcSgyuVlu
LTKRF2yu8wyh0XPFoCf2KUIpT+Md4dao6BIxI20WDIeUhiWuyIVnOx/sI/+3RSMU
rs8+VHPLq5KDf7bM3xXCj5cyNHMi2P/nA72CgRNF5nYSNZKCHgDZzQrH8xb0FLRT
i3l7Szb7LqanJVv6k2i4+Ke1ywtlLSkPI1dNR79E0JpznINaDpgdLG54DdXpE/af
Vy8VoA2MJGQlwD9sFQObrI2/dd7XkCztRu52Qzk9vG2CIDa1vMRd7gni2/JT5I58
kksbqRg87e80vlN7oL5dimBYR8Raeh9gLORDb1gc4Pi7PadLrsjMTHmGZEWrQ4xO
t0EvvL/WNkNGaiO91dlhXGJXkKMMW3PNsE4SWNcIp7RdTm5edmeWOPb+U3FECmnW
T6OAQFNK4N4rZSvmuD6KXg==
`protect END_PROTECTED
