`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LPCeZmoSDWbsINkqgEjZ7aqBSrkJAwQTkhOZ9CbE+oM80e8IbMFLDJA7QJ7yFW94
irvoBVqW2Veent+9tziGiIz5bdedyEMIbmheHWkyL+vZcNjyf5dqzA8VUOgBmhzl
JKLt8AUJFee8xjp9RcQaepOIxEtXdZnDdUx8zQOmQl3IOD7phLVVpcdS4uzk19F3
gQnBMIbHiSjN2vgAP7y3VjfuNYL2bEXbSg0oP2xBSLbo7yFz4wHRWJReG/Vd1ps1
vYJJwvjJ/sNEsiI+fJES4dx1tDF/mju4n53+S4LMyDlHv9LW8lRa5p/OoMhnvX28
G4SXyk35ktvGGu4GAQyfpoDhbhqRf51pKc9x4hnjaChfqn9OLaIFu299zAv4czSw
UIhfiGBoBjAOKY6fbbHpLDuWon6nUJBUQe55ryf7C5Onzydcvfa8t01NBd+UzaWa
/lyCHq2X6NXApJzKrKdGySlb4DHqcKR9FykOSWWdNpw9/GWEQdCWvfwZ73kyXIc5
zosrDWMNnesRbKPu8BriepQdakS/1lJttR/NCdGoMBn5/CmWGF85dvVNuVRbmHSg
1rX77Y3XwYy7zJaYQD67hA==
`protect END_PROTECTED
