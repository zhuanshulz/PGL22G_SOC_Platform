`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
22nGZSzhKYpQ1JNrgR50tQ6mZmnp7J67M5K6p0cvZkTxClD5ukyJLdARrDXRxACA
xlRFS+4c8AhTSuSX0uCQhTIHCNV1UrriR2R/ZoPxUmRlBPUfxrMHZv7lKb9Uyn83
Aim1vO7LGlUj0vtUmOQwn4XeJwaFEyB2KHLEiiNaq48whal0AZu+ZBay6kC8RaoE
OVL5TWPSQ5DuuYkN5sHp00EoQmQvFAM99ZXDGOxugM6ec2VkpXLAyTHWWB192VzD
eLx4JsA77jMVi5tbbawAdptfR+/gL+HCwxyjCCrzNNo7rXzj7C80WfRhmHn+Gpki
jTQIvud2ZPCXBGwL9ZzBLVZTFtN7n0ohPGBFFHSjAysKUxsXRkQ4dgKLU7piRNas
UpeKJmDEXzWblsiV5HRXiBxmwb09r0OhsPmaAetN8nK2RCBFui3wopi6QnoEaNAD
cO7VoSVUuxVVEcrQw1aPvNlvj36V1S2Mg1cuL84NUavoql8kfX8C2j4E80//ISOw
DbgfbIz/+3+FmuSUlUgTSvAJwGpMWNfy4JuE9s7vdPqn1uw1n1izpPqDf0o8szB8
WB7F/TBr5VlRLuYbcvFTZK1mrhM0/zRHtg8jlhs2rZG2D9uconU4l1f7dMB96hiq
Cdqcaf4CYdvFQYxZYSHJIJo6P7fRfnk6yHaM9I3nzi5zC+dQWXkVe84gXGKtDsfs
mmpA/4qjv0599lUUd/5F4sIiJgLaeItrGuh8e7aAoYF0y43ifQ4enbODX/DzuLg/
FPda/hpjCahjWvX8ZRU+QOJdHhEI6USPqWuLY3SNpVlyVDCK4HMuCxRY7DQ1lI9Q
xryKEop8nuna/bGcQqYyOFjsFQAF/cM6jeJXwd+2myJfzuuSgtzRxqNJ5hra4Wcr
QwEM+sm/R3Cb8Ew2OaEmcn9CYvO6n1d+A9r8ds5E6oDdiav5kd+QUME1I50GI8q8
6WJVU1vxuvXy8TlbyjsAepxuequjPLktaYPa2gt+Vl/l4y8sgrOBUQ33edX+yy92
1hxPg6b1IVGRFjt5uXg6So+93q8t34EJjGSzmgNn0acqB2E/ZW/8cbl7mfw+5Pbg
6J/f0hf4z4UfwCgg5L17pLaGX8dUOVBx/XCi98NTpHDkDDQWV/MDFEs4Pg6xl6CU
zEZMz1d+FixTGjYscqQ/WvFop7egeO+h2UqPjaXptVYM/+lmput7wY2vZt4LqC+L
`protect END_PROTECTED
