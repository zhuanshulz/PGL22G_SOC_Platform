`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WzoLOpQGqUQVTAywenRqpHoKRfw3Y5QYx0NCuah2EexylFyvw1mFwf/A0IAX4y7k
kIewEuXpLGdueGbArbaogEZTToA2Ic7KTFM0a/ipbpmQ4jDKaWpZqG5ZWzrhd8Mu
Mq43ZtusmGmdxXefpuDAM0zgdivlzQ02F2s1Rqjgpfc2PUpzmYavewaWDS5VKKia
crB1iL3dsvJ5Sl7oXWsPwTBFj+IWZpd87d+ybwgUpYxtv+UdlP9Uf6ffdINv552N
KVcbr266NYJg5BecX/R8uwFCyz1c7rvUb5njfRphGwFqq56Sjc/pukrK4xxm7i5b
lrcS7MOMlNMwcvzvFbBfSrtDecE66mK3BlTgnf76gmWsc16k+5jh2IvUtOMWQQVw
7jl3sKfR6PJB3xFfagoSEdStSwX1P/hRv/M+ZlhyKzGImJBqHtDf8bUaKX26FiDm
yCnUIWoslc954sCINBvZuL18tzTGWfW8j5Nz2fWmuzPmBV/6QRy++a0Krhzi7ij8
2/dAHO9O7nJ91yguPw/CBxR3W0AY5VQJUu6V5LTY3PWv7AkX1MyIxTVatUMAPHfL
oGldnyy8HipfhifxlbMkPXMhM8Uus/gxllS80SHWtEvysjmqx7PPDQ3+bZDJDIak
cJr5Ivt0BFXqB8Fw+HbNkizfuTOqN2ap4jWeYgpsBkMJWCa7DCkD8Sigpc8d8yvG
9DcbMiIb4piSm9O1Ppb79cc9ijZxaGSN4BhgJgAGk7yB28+gQjjCgOPkWX850ZwZ
DPxtscMcmSC1+i4U++aorIt1SklEpBkTTnzxGUi02nly1jnSZ1CB0XVJ3Z3Y8WUM
hlvAoI3r7hqdoW04+3VpIjbUBgGA9k2LfNrU/6pBJngky3/3KgaTBoST5DIvo2O0
z11fiO5vn/ODhzUL2vwIUsbjudM41ZhbuWG07mzqimZ4kgpe1J11dyCOPRWiqBDz
DpIKpXv+R9Z7UfgxoOnOQii0z9LiOJBN1mC42jXJC/TddmvukBel+tc7IKti5VQs
mBpyev6HYq67eO2klqKzY5cajJAfSmnPM3A8RBecnmxW7IFQ2nlF2hWX4Iao8zAp
MJ1boWzpdmqF+Exd6Sw/9Tswkeivc21/GZh9+IPNWzJHg+LLVFT/ULsy2jDMLXU6
WiVPp/QVRazkBR97RCwtLhdxS3cJfMEPVQ6OA2PQ5d2I1G+oVoEb8VfPnOHAcK44
fRAn7MtpMtlu2/1mNkMh6hs517sESyqP3iMo+1zlXyzT5R3fYUcsKsGunGhUs6W+
GWtiYLJ80z4Y47eBVZ8czrjN8i2r+Wk2zBD14jcXRSLW5lcasysHPCeZ29B2Lv91
PvkgNhAUJ7rXnYCz1NFy2etEQbo2tHOMv97WaR+JwNzQQOR6YnquUrmbHJwebL+i
1fhlP1Pb8iN4xtDsK1H0WaIgcnIzIcdd17dO+yHxbsCkDnO/0FA7QLhQdPgH5PiP
KGupZ4w1RWtow6nRaNm4SwiyuYkR1tnWiiu71bkZwquvXJwcN5dbyVfdZoCJjDHt
Rna6g5jXzjFfV/CRynExJOaR0DTUNbiExplVo3k414LkAl4hFr24WC6QFZEvMn0E
f4JURjSsM7cyNlvkR/st5Wmrc/iTTvanU+KJYWkGcNM1BpRv9UYxhdbE7iF/KhGs
rr2AttmimIqIR5V/Endz1AVHun99bGeKa9bR/IwxfQLiBqQXFRs/B6ZPPULihkwI
EyI84Kt47swhQb5LkwP+9PgxdEBcP5r12C8IFMWj10bQizKvkuoo5qFpSQ6wvy8J
GtPTGLUWlpiX2T6u0pvM3aeccgya/97LhdtXGlPL4WNOaIVMn/rPWuBRgeiVPP7D
g9V25BL8yXWI1kz2tAM0OTNn3UBZOQ6Cpjy0sBk6i3M4QAJxIKozAiEVDdeV8Yn3
UMQSMpumBqJJktSqVDGuhOxEXBGJNfeEqJxfpQWVEn6Sw82sznN7Pd9wyhhmWtd/
2XhGnkLu/a9BODBFLiW2zcKYlGS6B5mi6wPD2ABHRyTma4z9xafETuEPzqrAMjQx
prsePhYDqtBEUfQwWEUsDL7qLlmkGOykk/uUIqFwaK6Lll6wnz+9QBvI72n9ddgj
eUIWstF6iqnaKLjh8uC8B+WfJevYwkkr6jeKVTaxHG3UrnYuDzhOPQOvm++oqNlG
dT+aZEtCNr9PvHID/kdE5HOx6PQPugtxraajlSp1Ap1w0lPLBY8aRkxT430p/2+v
gEcAGPelczYHHq1hwr3sH+PFZ34+o6Ai6Oa7XD+cw0QgpqIlG5eOwXFDgMFLvRwi
GVC0bvBPfuS2WSUsFBHSVZXEyuJCwzpmz6Zi3d7mY/L7kwq5SYyqcebKHNvP1jgu
mfkKWW9n8ySqoQDD4A6kUyTYXZQe6Xm6x/6ksDVqNJw=
`protect END_PROTECTED
