`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qy4cQDJzrMY5Az4KRQxff8l9hAzMNcH+4CygkmppOSObRsNsqyH5rJHyDpcwr6xc
VmvQpiS9Ws1LtXDbChQCEKO81e0HmeK/Saw8DeXh9jYc09h5Dgq9GePDT3XhqvX/
+9K5ADefZJr3oVJZ2s6ZZWbbaFvPe3UnYe1/OI40E/3HX5nvv600Peib/r24bcsi
pVFa/YlhnrqX0iwTRGoFzspK+eQrDVnZW5buv5b/WJCA6TEGtJIZ6JrEU13fVUjU
NV7oQDwWezn9J2lzPrhqv/DcmMQsS4R98NiM2LTKzJu9r1a6BoJO+81akE9COG8q
6qGYeOuqG9rvl8q2XXhvMNbfnHnZQLKTRuY8MHdHIMncJsDnVfceNhsSKH9nc0Qc
lo8XFs/+4Uy9+A+aS/GrY3i9suyKVIK7Fxs6z9NXEQA=
`protect END_PROTECTED
