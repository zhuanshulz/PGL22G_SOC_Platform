`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hbpkjemoyLhUvf23A8BRpB6it1fzitxJSqy9qSeKSj3CeUK0ZjxTILlQtT3r7e++
zRg1gJTPHCsLp7q79q/DFDE/igrAvXozmm25drLEnp/cGIovcKzbiG7C6AO5+047
hxwBI3lf81be2e5EsfWsZbJGPiPEH43/3u/pBfJxVvRzUxZr1Yqw/QB5GI7P3W2E
kRUJE3ZjUQ7YgVvyCQC9gsm6EM87e6xcmnBjEw+1LGt4iws9pr7M4YyTBpVyH3X8
hkHpsLG3K6P6kJ4Rf52IH9SpVnEDnkrXwoRqq7tFbKrss2SJj3F8DgpwUoaVA7lb
0A32nDvzrAYfGegkTXedKA7hFMoj5hqPIeFptmOyVnBowVZIO7+35pmmiNoFxU10
AqNepvW9frCpKgIveUC11R9zTwg0VEnAIGO5H1QHr2wrWFbrf2F2JjnqzPzu04r/
kqQRPNDG0e90nMjElWNbpzADu2SQfcI2AFGbGqT9ZGhNn3DANL0mM5MQrvvhCMNl
DcXJ/K86GUBQ8UACCcs74UOhsy20zfzzZ7PnrXLMnpjA+LIfHzTKb4alnR3vx6w2
wqQR8XHuEdYtuKE4BPLMCN6taI5qTwJtrLTHbTtH3yV2ejNZqWYJd6LkFIlBPRpc
gBT3lYG900YMF+63BYEm//yBjSpjFNtxeLkT9HXDKtrjOEmDvqmKC8P7LafD4mTX
o1z8Lt1MHh6p30k0BmMijj1flj1SFrmwsrTF0nBH0oG/jM8sHisH2GP+aGqMbWnu
QRZ45uCEozdW9ZhjB5QqO+7gyRdEwFSZQ0g5dlNuekKp5J8Sn00wEbC7KzPmK8k0
9KZvyVuH4H9NuwfJY6V/4BzurPIGcWF48OtRnHNkkPSOy+zUdzNF0J9RfwWmQ0ei
EmlyVIfqasayPiJxMcNF44a+fQ3hnXlRZIgzRed82/aq/QZv2HdinCaVLNRjlZ9i
IxehJxhzFQyKoPBS2IY8lnblgPtWDhzZyIleROCKGXq+AdSiT9UlTg5+Rs4TZH8S
BWJew8gOLJYJCV7LqAkP6J+lR2Uu+TLzqIFreQ6PGc1qL/JfQUiVUkUDghCzImPK
k1JrOksIaD9SN1lyhXn0+VCIATVhsXH08R/9U//Uxo36BqeJboy+VUA9ZOEqCbH9
MeKzz2IqyrFPlYkZjPvtxSziaPSVmdhHvWY5QmpSa2pwbIOcLWP9RqxOaP03vH6E
byCDkBFkHUHGSfPY0MJxLfFTm2AJTVg8MWwXiIrV6Ajl3Uu+JpfMULleIN90xO+1
jFxkUDF3RD+GVpMHZi0q1gzEIzgm2fcBG9PM0qA+jFKUA4BjBTQx4VMKcHMI+duA
oKynoQ76ImiW9nvBQEA6CmncwTu3O6Fy4EinAGRmiK6ynyZHTALejyuM/LVar+rc
lTXtPMmmVDsy/ZVBXlowQkI8ds0Zi7dy7ke83FC2ElmhRNJhfZA2efUHfspJ8nsG
FpSU8pCFUMC9qZVM9cBDLiHsZtfEvTRNRp8aTOMhLQMvLdjV0GeMwo3i3iTUj2Jy
8b07UMsdmGkdOmyAkcl4XOmHhlE8QzoZQ83bX+FChGqBSOiFQ9G8+BpGtTZnvvGD
4B/CPidKKV5f+mTbPCFXQn3yCCZXO37P0Cmfx+AI6h+qKukISToDHalW0ZfqliVa
sPFEhIQRRgm6ievnheMbZmWS/P1mp6boWeKszXAJH52EodZSp6pKIwNYZ5VqoW4I
jKWHmmNp4ExNFGVBmc6pIBUaXcFCC6Fx0M6UH7HwTnG7i6t5o6x8R6CI3JYL3XIq
zI60GhKJIIITGa+wmyOGl8EqppMBbtaDNUhYm5RkqQ4cZDv3vtU7OYoofEJWjpo4
oGb7uNkXwmE+uhR3FRiy2QSmCxd+unq6avvfKpc725EHg1+CMgPWmPNak6SUZ3Fg
fx1JPpv6WKBm4QA75bOJf+CzhfPJoxEwa6qx7c/LXEHsHtWa0O6XU4t7jp/2Aurm
3nJqr+5YW4ACyF8Lejp4MsLlkx3DdSBA6nhQ2IjC2XJ/TaCpjiDZlcgkBD6u4S8v
UrVG6Uv3nk8fk93F2Jcjlp005nh3OfS9lKAt4xxknSHkZDd9IMcVfohkBg0Iyat4
tEg2SWge6bjWIST5p9/1V3p+LcEZETCoZxa6glfv17BThFJn4koU4vuNb/BhKQfN
Wli8/qj7qQiovKRxbaBUXiS5HzvUCud5/bxXz2fc2oLtR3abdvUnomXXWvUCKif+
ubRp3EqPwCS2tzsyGN01O7OOh3cZLJNKo8AV6YF4PoTEdeSoYGiweRuW8+12gmu+
KDQs9Hh+2E2+y2Dtd/HxQWj4K3K02uiP/d5Rhz8+2uj/pb9zevtYG0k0YIYAbGhH
DXwYXUXLvrShIxzSbOszqoChTNAG2EKG4YBSiQhg5MT8Odbj3LS2fqGKmyQiTQBR
aWcbHG3GaOV/S26TpnPbbG9E0yhVrb1rRBVYcoVTS2qcSZV+7LrSAvZeioqzdTsq
IWr8LXWQT9PVs4vSUjsHoTN7niS0sbCYjuLEx4zK8QoWE6jyy+4RH0bOV9eVNx/T
UZMWwOs7eJF6/ObS+3rfx/HhwNJ1sU5+BOlThJhQ/R+3/kjm0Wqz69OF6zhXN7eR
+PN0vdZkUJZsaK17ieAu5Y4cCRcIKcpMPZgBG9ZDIZ6InIJ4TA2btcPfQEDNA6l3
JUQQ2DCaeYXrQyOuRaBItD+DpSBcyl2zBcDLgrFrGAb9akry8RER0Sjz0HfIpmZS
srWFNGo7TnrCGMLZJm3JkWAu4WJdLkSVbFjAQ7ANTazhbYM6dcVkDkjjFzsrJWdk
Vl+rqMIwfXNVhhgfW0ai1Q9UkecOf4fz7NB8Z0oA6cYND8envJIlUgYwQbw0acce
L7Ceu/lWTq+jePkKhvTdMH0FeCQkc4lxK63JRvEijYz8lnGNc1/YzltHj2tEN0ZB
FZ8wDL2vkmNdWl5OaZ7R04k8B0UQO0JPnd22jtJWtnWpCev684v6+/LKrQSHSwsj
o/PhtRZJukohilLcRyuJrofAOrECqcl62qbOdSh2FhpNp9MZrBJvLcxRWvU6EW2e
BkqKuZUBtmyGAjz6LNBIwkHcNq/m8DB+JkuQ0D1Z7crUr4QNvZVEH38TtkEmz2dw
0ZQeIzMeql11S23BKueb7frs0sjVdGLpdtDHxfjKczxMwMaajpvq0sHVBBbaL6DW
35/EJ+sm0oaBEJ1omddGcqg3B710wwP80qnrbcKvO2B7LfOhDDAVl+7fgsfeFHgi
SPllZxqx25g18KaZW6YTCcQRqMj/Attt+2GUslrdx2DRSrpdMXLgpQA0M3P0B0UW
AyYXkd6IbYirIgFScv6Flyu7Sq67cdtvkdHL83HL+cSPsgZe9P/FLFh0/FZamDTo
cBTsM5+KG4nZDlWxayUlFZzpmbBSL+CWQjSLepZm2DKmURKdVyNqoX7Z3OsOPgLP
9Rt1apHh7FGMXyRGSgicG/Bfj/6qamczEJcPRAwSS6iOIXuzJ+mRnIjhdnrAdeKO
pXsm+oP82DTzUUEbeFcJh+wZGOk1gbtaxzsqQqdPYOxA/Lkpq4uRJSmjtJ+gO0Pt
wC8dNcCHhT6gdEhUKF/NfR0pmwd4k9i9yf0Ujzb9ecun6+r4VN8b8el4Hgp3v0fe
2oLBr8D8sHmEIOUoxAxxC8Owx0gj/IFiawRr4kjNZbj5U8/Kds8LjOHIBXBtv/Zn
V+XNVAQhwUi5MiAvttKOR6RZiJR4maQWXVXU6l/ECndtxOjpkRRxV13Z3/YNHIY/
dPIoA20iuKkYm9BE0HlS16TVx5mI3J7Q4hoYuzA/9QaqWMPxOzm5KBl/OMdkjSMe
muDVNn37LJAlefuoIseuC+MEF1TM8xKjPBgvpHy27o/jtdZspcCeb81dOd6bLyQ+
PbBEPi+vKmHHJQjJ5akit91zWjBD7+7jt0Jbe1NbkMQU54xmH/68lSP5Ta2tNy0T
m4DosMhZKjiBwY8sZt8FTS4aMppjvV2UlMTVKJ2w/y+vrC4OplJthG6t3aQIzIHE
ozPR6miMBTicWVvPn6gB7SscnMj+dUdjJVpywpFyhYfMB44LvIPI6Yd2LvAJb4vZ
El75G1vWyGTRSxsaZGgPObFEQnb8zatdI9JIDbQgJCe2nzUReCqtiPUcQ6HUNgCV
hnCTQTBE6ZVgbwoGXeeRIp4thC6QctLgWMsSh50U/oR63m7tlFLon38ywUfyk7Hk
G+fhe6zIeT+x7XJzc9yUvUXegxQxpgDN0VDozFRqFjGNNPdGfCGCM0rFPPHM+9n1
Y647kKfdUnp0ojIEDbnFHkbMFEZVUH+sqpAD/RULjID2lnkk21EDdpkEsUFHkjjP
oeQrQYeCeLjag+elB0Aue2Egg0VPC/o48U2ukUaZ2/cxy7Zrhh1ULAIocrjX8NEg
FXwM1O7u94dpoa5VIKbC9I8dcNg/UXScZpUV4fEP01AMxBVMZueDr0cgCCxFAob6
G+hS//IBwoDZUIwXr2kzzRTvTbJ79h4WPbElhKpCy8FG15FzL5+S9OSM3QlJeb1k
Xlz9gtP1xIBY4WngNdZPAaUtaEVnT/sJS+1sc73r7BNU/UuHhbmbIOf/32Vp2GAN
bvgpzQQKQuwMqCIAx5Y0spNt+LU5sDuWxaNnxUHF80M9vVe2cBmGR2AS/idotmRN
ZxdcyhFbn91li/ZvuWu76Qbro1NEcJGB7S2i4orUCyZg1/8j65pPIbDbrKf/c0UT
x2GsNbyjc6I0QCmquHIEIHOzt+Z+WTuCZdwScRkmKIho2IjN6P7p12iYJNmspcub
tC2ydiGsI/XUPCPZei3iTB+Clcw5JM2koJzUaWuUYXT+w42m3B6XXYe1j0+K+DfG
O9BEB/NyVG2Ukk3tPDcOhPRHogNHS5/wxGuGoNYCg0Yj7LdQ9uJJd4ULPN3e3nTo
LWOSo8c8rdHO9riOARkZec4xB8z26k4rYWrQDu3bpKDW6Wyu4Q1c19Q36Ctg/RAh
ddedTu8XAsY1FebF1eXuoZxrNgo29whOaq3TeDYooBsxdSuwqcV/kaByuZcwQQKm
7b2QlGo+Aq7rV590jk3FS1VIZAvH2UTDpWzBj+jOcBLgO5DHF3Yt6JfJNs+DUVtm
WZ0eDj2kw6N8gtha++fPRHztB9KQUrzLTpKTohtKiDBYE7yQ9Zw7CGB8yquUZqJY
qGlK92etg2A/qVWz0UW1N6ADBnOseNk+Gop0iFKtyD6x4TCsPuhGXox65pOS9Nsg
kwwnfKl1GFFs4XNoNEJIkaBJgL6v3XQ2/PANEYrLLEnVRKtEN8BwAOKYHEHUHiMZ
Roi3/h4CZ27koC0hUdCPaiQm5hl5f1Vol75ETKCII5szX36O0k7Ge7DtoXxLle0R
eQQnHI72wKP3KHHBYtGx4O/QrMkiDHwcTqzYeAVdsl7xXyGiLhVL8GnYzLJJgb+H
pYiruagEM2E81EBzwr/vTq8U0yOaNhEpSO9m2X3omnUrE7kBc2o5WUhkGwR0FK4E
NlzbehyA/i4HW5lBI5kYpvOu5dcYdlM31+molRnJZeZUQRZfR5kcXjxZpthtqELD
zhulAeuE01vtLLXmMhii1pq93TOJrg0BnFjSocUsaqKrwew/ESu7t9Z7t7VJ+ZXk
0P5MrKXmxWUZgb9wrixBknseYdNg7D+W45DW62WBVs95vy5E/8+pofaM1UvSgUk9
LrBe/YAXJzFcUlcgCF3VYiYVRjU5JeSzAW1hCG+IE8a5fBT/OPf+aM1BjCgQVYQ3
TGWI28bmkpabJJEFimr0yI5OrRGmbRD4X0WQ8UC7Wi6gX/W3L2oMVMp98W2DKJLJ
1zFgF36gSQGn29jxKkQk+3GaAaNocCMYTUm5XbRL6TA3FzNrhXOjrzu2mlhmYb86
QT+lv/4oFk9GbX7RDTs7rSxrW4nH62sKTWpk+GFAbArF9xkk7QJgMX2yeQABBmUC
PW2SC/tLdMwuinFkEwIJUaRAexPz/pt+6NYfOAfZzI2jgeTW2ArwuOf8HVL0EO3n
7uBKVaVjmscJjOoEucrpEtDMxsh/v/LG4hwYDhb5uLWqOrwtGyO9ACRHbmGLxZsH
vTuHWM2D9NgASYGbKhzP0C5aBgl6oz3+chSaQUZrGCUB93dnxl2ED9dv7uR2O/o/
6uKVcgSdxK7L3P6GAuCP83Qcaa79Dc8uxQ0l+1p4pRqgEMUvYjACt9BUuuTJS/ZQ
zJwdiFfwGZOd7smr5DfH/RSngd9t0IH4np/ykpNl35Qxg4YjpD2RiJyL9Ez5TmjG
jHbE5XRuMW+TzHTsY+VeB16qNOrepOA7vnkK1fWIfJCbNQzPn/CQLtNkNzTs39EW
lQVaS4yy9jinlSAEWAx7llECtQkpwpuYkiZ8xHDAEHLGp6VaJZkaPKXiROaXuRds
ptVmv7m5AtTCaorXUYIG145vZlF0Xh2UoGG7fD0+DWoCH6f52Hek1bi3Te4wesed
mHZbNcHXsbuV8F8r9jOZMEkTdyuKJYvzOUCHrEhe5+UZyDTRWLhkBcowA67Gd6b4
Qt+SKNxFVfLLtPnRLgf8RC50o2J6+ZPjjeP2bJArMA9+RSC+VU8cNgjNbZFfuvWI
Ccixrd1318r7P+nT60HQf+nhBmP92EUs4oAEkI0VnoaV+830X2p1JyD6oQW9UOKW
QIeMF8WXyxfeh9qj0I6+rV8KZlpTegU9BFIEWU9Lsvt59urnXZtWpUxP/p87+GnV
KEJ9Fwvpl9hHDQrCj4rVI2nudXKTeNEJO3QdHefQrg/cII0Uks6yZWLxunyjTqVk
Wcos/GowFkrzQ+Nrzg3Ily/URQsJQpo+k8zY+rvQ7YpZFGdsq01bSp228ztB6tPF
AywDMgbZnaKAIV19JOF7JyqDCHc+/KzpTIrtAz4EVE6yb0ZVEjcLpNZQpOG1D+FN
njS60xSS1K+/S6JGHsToxHRmm4I9n9zW1xKsrVUE9jHsAKuc6JvFJvBolVLpx8bf
RpcvrEn5e/8lpGOxRRZFTTFhaRUvycTqyBURA7y5qa0OYTAP5P1S27G+EjzbPNBv
R8j8pUH1Bm9Fk9amMdlxuEZhNvoLqfYrIUDAlfOvbpHdHglbm0QuRCnX3/wIYf3J
r+WEXFB+Mceot27Ol7myBo6NsfhzZEf1/nm3NVhdnn6js7ThGzLzlxubjkMyNMba
9f+b6uD2+5afqGyP+/e2bKPJx8nTg/6zpSZ/wcZlTQXO484+MRT8kKLcOcEtBi9A
nAH+4WjEsK0wyOZESk45i6M3AITVdfrSBwkgoEU+yfchIN3gZEsWpHeyrMwt4iqn
9mRfTlg1LEr/7xPz8dN2xHErPCuqwGoUMxx5osfKJfFo5LD14vhqdD3e0zUOpbQs
BPPSDS7GHdQEg62lxxPuPk6Coa2aGd7bq5sWY8dmY30UCywJisRm9eYCnBCZHsKN
Gts/zZu7H1QjxODMyKkknSEMYChgU9W7qmc2jwUH/SxUWDvFiST7e5kuXZ7L6pOd
4aR0XGNJlo+OrTqofB6bc/gXImT/Ocpd/340cBlfmc9xufUeSjQFfvUZVfcruSya
nrX9ahEXaHzC9ZWnc3ATjQkxBgLxwiWJXOZC7+m+AXmdKD5Gpw+ZuKa246JlGACp
EO0zD4Opt/wl7C/7VlfvFEFujjSf2VzFi7vweqFutbDS5MJ0JV3JgymoJ4BHvMhp
uEqbJD8Lzvflq9Qi+GFJYL9z2YvC382jkZHiwRy6ThmcdeScurm3B+QDqIR8Eeub
8VUUeIIli2/lVm1pPsegULiKR3Sxf8LOuglsXQtU71txeWhhxWRNX2wg7IDg0vmP
mcrvwEIjIqwcBLoc2noxfkkjrVPSjGWngqGeIIxVzXexQkLxEede0DZAWliKEEpF
Kf0y/iPOcDD3KhCB/72jDg035PEDpx60a8D2CbR+lxm0QKQFPnIAfhLIHXvn0uAQ
Jyv6l8k/V8uyQYauR+0+Xu8rYvmAvUwpQCRKNE8g9c/rvrZrrs6erqwXX99ujWY1
XrS2tjQnZcQVHsQlh0q6vUSPnivKDTif1Gu/j96QetZXCU16EJLPXPP996XTXV0x
+bFzcDEv0hhnkNvD8RK83CfRDycn9i9BrcRQ3LFdIEGB+DvWOFQuiCfRmVj2kpKB
heZxlT5frtgnWC3NASGsaIf5SupwHaGNw1HWZyklHNJFZ7dbIN5E6INE2gKSa2hy
u+/zLc/+Qw1FvsCkss7qP9hl1mFa6Ay8l5z80IS8j7AxJlvrOgFwEvqZChtrbco6
TdiWoTvepMrRKaLH7L45qTLXG2x57BmkHWb23KbW9AcAIXUkG2IFxVqtiY/dTs5q
DWwW1xseXt9zyGGLU5dRwrEBILS1ZSTqg8g3EaUhbzp2KfII1gisXVZGg63+qb1O
EYZXMPDljSrE3EvH6w9kaBbVIMMWz3UnT5QdnpFa7JL+mwU/KHHSJct9cIsg9LdP
cqsEgmz8tsp86EVUWI3vNu/zRZ8QqKUQACUj5X8bX/ucWiBTiklAOp+WF6kUFX7q
fIRA9icnkf+vb1jz9U2yI9VMoZdVp9qFPM/lbdYoFynBhkKy5hkB5wuvl80CTbFg
mUjG1A9JPw4e0gYXJsytZVOd6CHaj+FbXdudr0hPN8q+Z1NM67TC2tRbvrATpV6b
FCh2MkY2U4gpHaQbHQm3GUdGJezGYpvZSVAAeT1yuKBMze+PH3QAyCjuoS0S7YEC
OZbTlyo5eKtVFfPJ/3nwT0aQkZbL0IOpXZKscm2/Apc4KguKVb7zvEyG2kXsiOU7
Eq7l9rY+OEEdHvuaP4cOybUOuN23k0kvGfU4CT977Ng=
`protect END_PROTECTED
