`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FmB/yPWodcv2RDkljrfRcT29EzPYm6FGEht1NG2aQcTdVa0iQPym8HIg+7wayoV4
Apmwu0Mx1C2921tFGIi59xTbfmSsKXAyD39LZqiqsWuXAt6UE2yFUmMID2H4NMBN
qIyGlPZtp5Rb/LE4+Hxw520AC1FUpmATPrj1zoNIxNIfys5Oq4UBXR3ukBHYtrX/
KLeGcU+sCRm4/ny494YoOfTe1ej/jBpX7z66TNujIk6SVUjNFeQNV9tyxjx1zSpK
BKOd1WB1DRmUvmu6K8n5Q8sMdmQP3Z18qN88oqlqaZp0CTy8Tv34NXQjYBc4EBK5
1q6oE6YdZBVY+FQmlAZiGrLXXxBujASfH9K+9tONyhgJ3ovxCxettJq7Kl1fkDFW
vndt/VttGzoGQ1+jkfwTnOLAIgjBih2jmRB8mbREQQXwGF4OP1ii6IkB3ZMj0bJR
9h5MLcbdcBNEE/Gd3nvCZ48A84KpRVFQUxt9BaQo6NYr6Q+JNfwUXikQpa/MfHmK
kp9PxXV0ZAlkg58Ab6R16msoLiXryNLE1z7CqzBYsvoR8+NB2ak9n3j4Fl7PD2Kv
nsY+Noy+yFrmC8CibzAGCiktLNZlOF3jnS+KiNHs3eMCy9050Ou6pkErIUWcr+4F
w/Xrno1UP79s5/RHnDNiXcB8Drp1kX8HsZ5gCYVCyxczWaa69ueJJE+hf/D9cUaq
KbdRuSrl2ekTgiuwT3D3K+x41jsRWf+dTwGOtpOf+wI7CVFUiUCrq0ZKDi5IOomg
Bq6tTY7FcuifBdQmn2+ndf350n5B7O8dy/h94d+LWz96DBN413WxGEO0FzMXG9up
i6/5N390uxemB+U8VsedNdTU2V6dGrzZxZjEHUQ355ksKIjMor24aRJUXKxkEYjf
SZNHUFuJDV0PD2L8OhIvFdNpSLviO2qqD3O5bJI0B7iSUZGKZVt0xdEnwEOcOYMD
EywdXRJNzPRfA1tT7v8seoTlT3KQT1jp2sB5AMSGXoGV/NXGlqW07T6jSwnKP9B/
7l5UMrT5dI6JAutm0VZcWxyU9o3QtNBtZfwXuA8IjmumaOZPPbtEFtFoY5ItGoPY
Z80sALsh8DwRW59fc+zjWk5iMWDJlqcamFXRhNPN8YsimLp/93/wZargBQPoIvBm
YPIqwLPK8x8zGLv0FxaeUQotETsTZeSjkd6Nwg/FCjANW0jWgBZ2Wf10C25WfxHE
tN8C9w1cpzxj0nYmtpmtwunmkIO3o3QZZFS5vurQCX/RV25uc/A6JdxJZl+dgF+Z
cMJsy6RbgEQl+azeB4eFEfAO2pst+FKNydR/Zimi1SOfeufYf5jbpEVnFNhtQa/Q
dwUzknwjZoX0QZPPNw6SUCT0NtUtaR235+zUVmWtHMzMMV7pcfvjBpj//s05wUzA
MqrW1afpuInKWKDYZZwaBz7gBE/6cxxZqAjpigLJIFUxOPDK5hZG5xMXnFZD0DHu
Qv6C1O+iL3RYpgBU+0QsOUMvPh/vXGDBUCz6vxBSF7sRxwE4Gciyx7Mm2GJkSSfR
q938rWlWz9VvgNVbRsjqFETgm/9gAx3fFPMOwMlSsV75hrvzk9cb9IavnHQHKhX+
MFQ9dmi5v9VfWC2tx7WKLo/jKkLP4lHMt1WqhDhWqxpbejrKf6jSa713dTqBarD4
A4Oux3yuhPUAa5zAWiRTWJbcC6Re5ScWwMKStRdSBqqqNhCYuQJNZRRBJwQ6ntlX
vc7Tnr3nyt8Rn/J0W1Mq4UXbMYDLI+aGdm/D/Q8n3cxbEtIV45Ug0V8ChwHag/gz
md14rImQ8s68LzECnwY63vaLnUGg8gcMFVhtaTUM1L0t8zzjA2suzuL8vsnFCdJp
teFAaZKmlSjV8MijlkFEWpd3dC5e5WxJS1cZjEHPdpauq5x388qmk6SVhTwQ3fuS
VIArU1n3WLWdpa1HKedykk4UNw8InURoMiOrElaD/paWMFWyfJyRXdWJHGp+t5KJ
nqIcY+vejPs2cfiL5ZyDtJJWfRyEBbI7hcJYvu5VwJ6Gk2x8U7lYHFbHXRcwnc71
FLoU1K6ijGhrQZuTFvF00ueCuvXPo5XsiNEodFNZiq7HSA0k3U6nLCze4FJw8wJs
WYhedv8mNMRIfSiIyEeuxdzC+7+WP8BeBX1WjMjX3xcuoEho9NyCE/ocFvwpqn7p
0yn2JbIjAxncpXZNuPhtBz0hqnKnPCluK+7ITG6IiHczvzBqsYw6q+cki82x4YHj
976NC2k9n8Ih5gy1rXMXeeDbb2T5n5HKpOVqlH542+EznR7LJz3Bz2SYyshQlHa5
QdQUXxZVJJ8A1G+OUhSS/SsA2cbMUflKJChz52YdwFK10t/w/iloANHm3p3Ai+9x
jshelVB98znyjpfsqszOYQiYpyisFCSpLvZ7SiuR7pBNwYJrcN6/JShdGUcjikA0
MbJzQmI6H4If8uM0uwdomvSj96luOUzBEZ2ov4kdYu8j+51sE7nmL+Z+sV11Xvwc
1LKpf/tZ/HipGrEp/LADRMdSJApJ0G8x1qqCYsEkl65/wul9nbTGclsGp3AyeQF7
Itdm6Itv39WpOfZnqoyBGpU8QEmmIDL8giRe3cUsXlhZftOjLLHexiotAOGyEnm9
qTr00O5hzy3I75GjA42A34CLEtr44wvMj62uZsCBB2k3RqJdGAhiVgAtitHUyate
Xxgy3VG6XbvHKn4tTukrqK3bwkkqwZ05zZ+gOoxd9tnRniE4q8hw+tHT015T7gXL
1RL0nrHdLH1g1LE9eMKX1Ut421rgVE7YYntoKXG2dB+HvP5w5XPRk5WWGz1hukRp
vuGIHUIIKXc4j7t+1Ilw9XRJjdXaqZvrg+W+NpgOZ+6itDRGxLEwfDOxr6Gyn6T1
QNydx84GDyopGW+DUqOCcbZUzeqjUAUnb2SuES5lVvUwPhaSQcyFfprEtR59np0l
kA0+qTTnSGAi5LsHp+hvA0cysRBzDaUB2w2UjGmNYS0PNFIUI1wmGNfVIg8tB1wR
nDgK/qmALAdnDovkgb1Z+ZBwARt5K6BOKZGHzMdbaa/fSyM+7gJ/p77VsETpQu3D
nfO6U89AwKefAD8ERxRgwHMVFYX9p4iSJ1UkGmX1ph+1G+fqgA3/Rj1upVBQ/jZK
ESTU/o/Qfrr08B4QXs+CPn3Fd+MwCMOYXksJof20vMN4uRX+95rEifkpANf1pVAN
7TohRcI9LktUHHrvC7VCRyVs3Kztt2rF1itx4oMuyMLIFwMHcf9LxI5VDULiCsTG
TvqSgO6X6vBWcj/ZIFI6oGHOTZrL1tAKBaopQQCqLuE5o7oqZbgzLzkjCt5WkLnr
9AiAWISwWsyudNDCLwEniyAjNLtFiqyz8KQU9DL0sX/bPZFAGzhn9Kpltrtzo5Ps
wC7ehy6OKd4BgrVNWnGCxdFOic2ZAGvtWAPwbcWEY3T8KwvMbz+PDWNj0qfw7QLD
JGZH4yncGizPc7Bok9L5MMxPr+LoA1CGF6+0O/4lbNpl+JnalqStr04moPxdUWXT
4YHBOLrrRguvmohCZpp5fglYEndBw/g94gIci4yAcENUdM+OlTM11qd8BRMzppzz
kHE0zfmf7xSfst3EJ+wLCxXJt46hBrzGB6FZDxlLwwfhnyF2QlICdVP+TY0Hbwt/
zS8/tAfFHfwXc1MQy9buTRLD3cdbppnxkcAQMuaVOUUYnCAWwv9Lzc2XJn8wupQ8
peOZj8Z7fvejjILLTymUbB0jYGONydeNST4d+MgZRxx72/ulmM9aj7cp/aLfOacg
m0ji5zjxReiKBJMq9nQR96ulsfmXbBMVs0KqjdMSGgy6INq6wZqkHoxBJzItYvXE
Ma3bXxj4dUYED03YsWL2po7qV/BcRk4cTVApIWScnYHqAIUNTAbwH8QISCu8viTV
aYjbqJ2qefijN3KFD20TZ2xLet37yKpJuzwS9S71/Jz/ysBrTPAbWiCqEWgh4CT6
0HrpT39705nEuSUcd18j1tqvGK6qEcBRoHe1EJDD/Y8Y5HsYShvaFYZMUlHJn4hg
kCD/sJRrcNIhWhF+GQqwUxxgptssn0vGOENta6qqjeapiAe22vKnTOUh0uOZsHVR
o92cs/T40gNFzk+qC3PLZ6LV3oMJRvH+NZNRIA32x0x+1QYOJxmd6PumfXL20Zfv
72zdxDlS495fg0JYTtkTc2NhrVT5w3SLFNFPYhIM99FfKRj9dbVqZZSuQie4lucV
aNPaWQQOJzBYCeyQIIp9skYirImUc+51Xs1q6SrZHBfCgA2dPA3sg4dK46cyTusi
yBirpIjohqOb2rbn5x259ByMrJt8aQH/b0DAfHIXBMimKgR4JfROW/ee5A8pxRPt
hvp9ZCiUVl1IzYoBe1eMKeWJOK1EI3Te3U13I0Z6EfBZTlh7/Qr87IZR5mNrAf1x
cl5XOdib8bmC4YTL6JFCrmlOcGZ6TgUZ1XksVLDtVoFwGEpyM5mMXUWh2sipYpt/
kOj/NPKd6ghhwH6FwB+Zvc7OA6qcL0lxn/XReQw3MuGnjFwYUCgFvnkZUlEWzlX3
Q2nPM7FGmVlxsnqBIFB25Ie5peqVgv9mJY0/iKE4dYy+b25alb9X5qePyS5GWK60
OioN56QAXYSpHknAi4T5tnjOkq1uWp6wLyIwrWQ73cW76vZhnOTovNiGtovDqgDy
7jq2pLWyjQdJ94R/TGf9pu8wSFkeOyG5p4AmRsjwXDklTQO/upzDWSP2T5h0y8Wv
ADithsjsOrEzYfC6sito/PPOWKRpscUHz/VOWSbzP334uCmTdICe/S+yiNPq38Tn
gY6DeCa1fhqxUbLC6hGqRXv1IxRDeSXR7PFi4j1h1k+v2jjQpPH4SfB4w7l2J62G
//gCyPMHVeEvEKohJIibpTZSQHKZqRrd5ryfvJw+KaNlJ14nG8mjH+bkglKJcSkk
8vd+lxwF4bdxVL6SDbbq07G7cASc7SxEpv7OzMt3bI9yFenngreDN4wgGSrPtj0y
B3BBdX1EN1bI9Er7ncupl7rVhE9PuMu2aQ7hisjOWBnEV5VRp/4kE9faM1xet8T1
mB08oAUe57zuaktqqg9kWnN37X77jqAic43tNTdGzZ7UXGPLryQXKeb4m+dJN6/Y
dBRSO5lEZ0MQ/GrZEfExglFB2K0ld2kowOIJ7TbyJuhkSv41JAewLgMuXNS0yLP5
a7Cd8s7WTaBGTLZa4v8gnfHENEt+j8F66Uai+DUrkc7ysHD9ZXOdBR5h/n8pq+uW
HKS8FlolkArEAhacOYDt0mzZNLXEkDKfOV0i1F3Anr49lJz0Ro2juZbjVboth/zD
hk0eASmA2+C9pY4ht6iCyXA1UsVmQCGb46+JoJOxfETfUt93EO6GgDi38aMgKyxh
i6G5Ed9t5lVnKy08GAD7FYBSKitN6Ci9Pb2bVfa/vTrqyb/d76fWaQ16CUUUhZVH
fkc3aKP9WXwqqX1vS+4tOziCB95TfqyAeDWNp6iG3YMFuB8B6zMYTnxlF67dQ4tv
zJH0wJZqTKAQuYpWcZWvgtxmnPmNeYtMct1TCIhf5uF6bFGFifkqLySRqSDLIKF/
E/YvcbJwWAQR2zwZeagEoeqhIeESWI4kuzllfGK0E8JBHEv+IWQLtBFwiojEMNrC
/sRdqTHvd2VrBSr+s4sonBfsoY0CQ3I23N21SOIoFxlBsNQ74f2JeX01KVIunpKJ
/D70SqlEf0SXgzBmyAHwsmUT+2cqg1YQDIwxoS8hyFReOFiaEq6dstUns+zuhxgl
`protect END_PROTECTED
