`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l99vl4U1yGwSotRF34v55JCU/LpkOJt6aP66OjCLU2HPDWE4p7aCcBd9Yzy5kmUx
SEkyl+nzxy/WgFmYeu2h1sA/ZvoNQXQkxkvRiqUXfTRl4KWhBetCDfZLebLmRKWS
N8fH7WkZb9SuXhzxAuEPLuMZEukb0ai8vICTS/N2NAbFR2nmLGHVXzx5kYZAyCZK
S/rNYGUBVMUW3tMJDu0lGXe6vCxE0caC85nYzTrBSY5RFAGTPmacDPAZLn6uvLQj
5n9Sh/RqosqRTka5HKqM/NCpYfPBg4VLC+CXmC+rg1iZZK2JBvPWiuEF+OtvJvvA
VYhsT4L5U1jVVIqjjpgkq6F3mqoynHz7LCKhJzBsOgR+tvIP2qIFwY44VWeq5OCx
L//BAlU2LICntQ18WOeqRHTvnPnGBDBRPpB9a0w2x/MtHNPRwXKucjQyBI2F2aOo
zdkigwhMrhN0jpiTBcCQyA==
`protect END_PROTECTED
