`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nEl6hRuS0Rl8+WieHsXzycnvphiva7D9xc5KToPhoimLCtWooqbkP2Ih+clLJOAh
XPr3Yqw57WwaEeZLYvLpE9f4zfqEG+7rfqPctsABh6Uxw5objVfsy5Ud8DLWAQ8b
dfT2oVlK12PgKxJA9hTxQKHjPte+/Oq3pSxov8QQdE29JU+MVfSM/8K7iXhp0avt
DTpKEJ7JThrdZP08+szkjk5n45GjnXvE1wsclpO9gaX3fkW83mlbsbqo0ppQhCzI
Y+eKd4c1Ef5v0YpSz82utIpHODJ07U+Dd5xfvi7fDh7vr9sgDJF9xEebwrpsbFfu
BiKfubr35/o/RJQLJCjVRG1BDzKTyods6lpLHe74tHVUijXuZR/91m87sat8MlvJ
Lb8L1plqijnsrCAGkJDFlmwQjeSFeJwWZrUnc/GaUtFbRzcBIoG05EUIIotxDzbm
UB7E/9+i8xz6ud7cLYfa+gV5O/LYGoiW8Cn/RekV33PklMfhGK0iOg8JuHH5Dr5j
/iM8Xt7l6JbCRq+Swr3UaCMWlyGwJMYLF/rCYR9E+XuiiqUwMrr+Xvyw2rCDq7Kk
GBEuJjU3dNJsaqJYasxM+xWtTAcr+GR7oWcWWPhd1UlsMm/sYorzuPJnuhMOxoJT
+SG3pRUMCUGMZauOYRLcJQBAcuOAktt1ZE7OAv8riF4TFHAHJPeAAsZU3YBHzII9
voYkxuYtwf9QTFsSKl35I2Xrywjx7feypymGNV5B9+VWAEi4/nViApwLbF+nJP5y
Fh/g/mqAKjOoMLRzrZuOalo4eMWyWw+V2oyJWKrJJxWXWLCyQvhTJ4uovXY7D7Cw
RTLZ7hZMAz/j7RVkzr83Kaf2hQTM+F6E5VPlpoYKpv+B91zRmh9kDdvSxipZPeuw
9bgoxOdF7Wcs+fX80JXYAAmKRH6FqlkkEOopYLMbMpw6uun10efZur901L4Mh/4L
PBOJ69HrgP9xDWT3y0lP0e38WDMZ//VZP+dZrCsq5IMMtiDQ18CHd3nLuW9H5QVg
cBoVivlo7S0k2OH7jTiN7pmj4JlL5Tf9IeaUD62Oz1CaPmnvdScWkTRMhqdUHDey
OvSZ1nBAwrc7JyfyHwWBz46NWhrcCH5nr/ctDWJTPCSDtPyv/zslQLebqZ9s5u97
B0jyF2xdW2pYpsy1PubgPNK162ysFUMSlw5JtcifQuVm8nZGm0SoUD2SF9sZX1+N
LrS2yqaRnKY/+NSR1HlK8jV6lvxEfP1eKoMeiO+4EZ2ThMOozs0g7PFJ+5RGoCqw
YpZVv/040F00LvobioBPdm8sOcFADI0HWF+ACvyI4MbkwtOqhBMUlis7t06DfZv6
WWg9hrx2138zj8BnIqzbnkoTO9yl6M71rDgIUf6wxm+ypzqNVocmOKyBXBbWsRo1
JkbUFXkXFldMquALnxYV/kzH5izlW/wxjmUxqLuW4WVX80ImwsDGRp0UFZ6kA9BA
kLUv3YIWuU4AET3VfwAgVdlEV5HlGRON/Xliri5wAKW1zp+PPqukgP7GNYZpkhhD
gBy1Mv3RFE096YyTFHGpuy1zuq+6pWi7Jc/wlyw+HjU89YBT7mqJu3u3ZriE8I/n
GQZtD6OoriS54MNHv6HcFXK+ZraUrDXCtbAfLzt2Gzs2c61pdjO12xi7tiFa4EEv
Dq6wRP6n3cSn1ZqEBZ6wbrZDW/LQTuANkrJT2FdgSwzOldB6wbvqu48iiW1NWfnP
oP63JVJtiWzPlWjxdG1Sntzd3iTuT0dQfPdE+/pfbBWWYNuyg276LxuItLQu1OHn
KBwTaUugZtowSmgXTM1PtuUvwLyAol2F31mBsEkrgSVc+fRIXCdr5nta7WZnck6C
jEH4EOac7+JlpEZVo3joPCMCRTtTBO2cvkQfZVkiFqRswmjXJlkhMZ591h8E3QsL
Rax55ncnxKdNnABJbfp9FMx7Cdqec1h+is38sIscZNII/yurpB042RYokNZ+1blP
tZITTPCC2Psm6OYbP6BK36u9fGPEx7sU03pCLHdwJRprgxZw6mTGoMBjZEYIb+b5
YW4zCsWzTO53mwE299qR+BAzS8jloZye68HSAsgsBMvnmJEezlbR2/T3JETVbT/t
IVFbDtXuyOzFKceESbOufcvp9yKqXuWDegtGNNLd+xQp7R6nFdbXPqKl6arE6Vu4
HVaYI5QH7Hzv3PkQjkJeJn3gZR6lvkiQyWSiGh807ro4bVCZbkvURduNbp8McGwL
W7ULFjeXJPG//99l8gH2Q3qNqn6hJChHxl5QSvU1J5fLQrf+r1/EozWVrg+izrm/
ypyzvkr9rmYeQh39i9CZqw7QwHs5d8Ray6pabnOq8h48PDTdDP968vTdZ6f/T99r
9RWx6Cm7pwZPlNC1yqSKatklV89Bbxp6fZg/c+6/UBODy35he2x9Wvpj9LkSRw5R
+sz7NrznzUfmzrQGUXRGxjxVXaXyche7+Uq1o8qciinxg8KAnNEl8+dCgYrKczQP
ForxZJltXjpKDbxzE9E08oU75Br+q0O/AUX64Q9+ug0XBYglbt54jRKkOMOTTp7K
YYyD1RG/5htut2A/+yCEyizkFxwwMhwwB64Uzhi/XzVVrJxV/zOLmjwJoUiBsVqf
cX6RHdFLWcs3mbVBJ7S9SRyZZxf9eqaHplakVaup/QVrRCxLtZPkkGGv5s1tuFRn
ThPNn4v1sh4Do4C/LQIB9wR+HBx3zZP3GoqjewZuEogzDIPKWVmf+/0z7BhnXS7D
hx1LXwLAI0M8LoVOKD4se1otC5/BCk9SMUDQiRpAzznKQsf55Bu0Wq2NqPWSLrT5
4xDsyjxmjl2NFpZWtn6aTGQKZho/juA9rWbnUsSFvyElnzeMoSrmRD8kSYjPR314
48yX0dTHFVH5e+cWYA2kRzHHsXVT7C3LogZl/mgIjey+UBwXKv0SxNVWQphMOlmP
WoLs+Dqsh/T5bywolwIieuXf9r9AaGXSMM+jQ0t6sDAvKHfRKlup9VgKT55WRJQz
8E3vs/LGuK5wMt/uddyk6dajTneGsvvG+NaIme50vYoaHXWn1aFE4Z9KuoT4HDay
kTPu1C8Et8qNAirV11bhhyNjcLcLsrEN5Sfbw95y7a+A4DJolsnea/BudyfIii8m
+0S6K82B3w/TJaulWWHW6LYgdntCLc49TbEL/xbIKSwaL7duuM+z5QjuNWZdjy4L
58UUnzmMnbRkkqljNAMIPD2CHQNpM5NjvX6o3j2npe+3+tE2w5UDlQGqXDWtmwxI
ZBw0efcrNut+bX/fUFKsH8M1EfvaEI1aVkOPm7d5Rpxfvs8drPH3O2nQ/9FIcyAE
Pjc1ZvuXpEnwM6hB8Is0HuZilI3jWdWDLPkV+OKCpHoQNBx8Hq0WyLxTUIVMTyss
hFYiM7jJ7l6UL+OTluxcLzyZ7LI+igxwyzJWiXp7yVWw7b8PVQvAoCrMLOLlr/sH
G4XnCErHP/h01Eyw36+Z0g4k96kYeBERlMLIPVOjFoii9MGyEiSG+l8w2Q8yKPIl
M5OJdyajDFabcQcwxU2iSSouD5M6Tip1oAdlAEdDLrHNJ7uVy3bsIg6+JLr7ItOO
0DXwsq76GD7CfKLBmA7gVpHKojCjRVcxSfvjSmLEydLDDHwAtLHxdHKsn7q+yOe0
BvFkj0PP16jBoGDNGlExEmzThFx1y7yxDmk1E37NMcLmy5EmvOaMvxlaY3v/hq9m
4DPpfEC9sg6IWXgqIaypRf0ShBd4Z5/Nrq+79p+4sYpTU2KSvGfheNozm5eUN8uA
PVlTrwwAKGaU+VX10KtZxkzEiubmM4Co1Mi70aqzfZE96VVoBw2lzCjA46FG00ES
TDY979PrIiJTc/he2zxgupjYAGByRhR0CoBiNc3LU7koVUlyvqkMW2hvZqmN0myw
Io6kp2L4EHsm/oLVOjTzU/dnkcdfQvtV2qRnbwSertG8RE5eBYUuEvhVw4Mzljdh
JxfaMbBDYhwhWJbOybd8ea6epdoPiJcG3D+pcZP+WhsNe4Sun9EteG4Ylt1JUtXN
Ly4ZNrmp3sAr+V2JwEmPje5Ra4QYYuIibKcNDPfAKA6uPTD5wR38/DdWiDMq0ylF
0Q3iNZM0aIvtC/xhgIdSOs1yuA8aSHOgdPx9sYlnOoVbp6ASdD7kSuWS1G5yLymG
zNLVAUpuds5TGnWS21j/gR9nTtaEcoho9CL708Xc0lQQY5Jt8A+4hY/3wCKf52v8
UVqE1I5EEB6e/9kFeADSiU3W0vTvqrPHKsbZk/j58DcfyGVRjBijDYJOExbCRLEz
NeJH1EdUoH5WsF2PCW8ECesUZqHBQT33tyJN2UDn4XxDFN3h1tr9TgPgyYTYxWW1
6E1Ers/qfRHtynqQ7hisNis3g1Br6wN+HpMR5Pj3J6QLPDLp5th07ZIn5wSVclCw
34uL80zhHQwWfXEEedUyDoMNGR29FI6EQnnMOB19inNmpcMvfrPVmAtZe4bD0RPZ
UwxF1eWh4OA5di/5TyklAi+UaAtoxRTh4IYMaFj55lnaTSwfMEP4eTLoY337A0pm
Qq/DxetDNUSnp0RmSRS2qtgx+3daaqzXYil6tn9yE4Sh3pxieczKW+8iSEogL8LN
myU5PpMGJZasHWLdZm64OARN7D0CjCvKsb6cy97nWogt0G6IeoebZ/lbjSYfX4JC
KaNKRTauGcT9wFghZhLQ6NJtFSfmNgKdoEh6Rgk+RRCjwc4xNAGZExTCGg/6mVm9
8w2y+DHPoRJ7ON3d+oQ1eAmxL3fjzXDBLwSEOkWD8DSy8ZfNM1KXE6wNzy4WJHIw
CH4XVIKSwm8J7tHntRkffhxNvqRydI+IXIfNvVCSE6x9rfL+CPibNRmsIz72i+LH
E6lLLmZ4YpZMaBlSdK9fvzc2/hZNFPshLrE+C3mn77rCD8386JizlpjpycUli+8Z
1a3CKRUdURnNeXzN872YBWN9MMBV2U/rvg1wfji5P5bDYeFjjW1rs7NwtdrRiaTW
b99BFWo4jD76BWfmNZb2A6gKJjeHHXTwH8xaSWWbIP7CYb7yFjdg+ZzSTgKumHbz
pASYu/33HqsAJgCnZ6MaVIHq7e4q4xCTLWZtZN2p2sz5jcxDI6uDvfJEN6Tf9Jji
Lt5bHct49E1qzkfuUa/5eE10LE+ErFztq2EPUav13oCNB1SZDvlDQzv01w7fVrOb
VEu87KDruF0hFovT2m9IZBZ1GlEXExvPJYfyJPMotYYyYG7Un/5k1L9VKWn/C8iq
v9cS2AtY2quoMVXn2U7BfEDd2k3PIreGWHYQGH0qoCphBc5efPVOTRnMYihKAas6
fvpSfpTRXqVI2SqZ3hzgl65auc/satmH3T6mjtDP21DB8NtsKlHXk/PoNvIi1Qrp
L/O8MEyCNGSTgYECLccba7DwM64ELa1KRQBBuW3u7BKT9fWcKVeIhE6c5kZdpQ8u
HAsxV/JRmuHw4j/hBqDuclVit4DtXnL4hHgMtwL/M1XdPvj8TcPMMUruS61xmRKC
2MQQqeicnPJxMk8tQPCINu7bL/hH8KJCRzWwewJG+0i0jZ2GQ+9fo+EXYUVHMSf2
`protect END_PROTECTED
