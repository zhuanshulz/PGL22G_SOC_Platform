`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DwXVt9FmDQFEP3re6mCHKeAiwEjsu3epL1A4+p2TZu/qY7XqmD33YbY7GVEA7dQY
4lZL/aqamJ7dmx/xaRvjraplSxUKA+N5fLDn1r1J73w/ejbNP6oD+zXa5+m7Ev2y
Sbo6TPocfPPkPm7WKvXzvv7izeAaTF7UiQ4j1dhw0UCtIdOMe5Y1LxsjcKnNLOJY
svRkRMqKq+fz0IrKryzpSnQw5H5rNq7UBVdp0rpNg8ZtE5ap6PiXCEIi+ua2DUes
rS4Q+PffXPsy3mYqTtHTFbXdBDsSE18TAYgmhOyZselmMIl5mSQIeAlsWgvu5fps
Zx3OsqWFmSynr90syaycPGU52AoDnWWO3LpkpLXQs+73x4ldROjriCjU9UoMXn7C
UFVeNKbc1sdo+VofF8iiJtpIbpadxrtCQ/FjAWhsIuVTHGEG8Xjw17PQ6D0utZ3/
pwwqZJQJNL3RcUV6SVuFLsVgFkt6pcsOr0WLKWUB0C4VkRDDxWCFKO6OPvQAuTC+
PzfzmWwkcwr47FtoLYahHCwmEp+2dwVCZD+vUa+a+Owg2r8Zhzc6M766QJJf3RF2
xjmBcTHOr52bMlLDS3Bt9bqNd2aSzQkbrkN3M/r2LfEHWolXjfc5zO4buqpOKtT5
fZnm67tApgKb5V6aUDe33kfSNXdr7jDIfjrM6+7a/I266hjyilNlcTgGk+WZxbiT
sdZoQ4jqVLmeq4HFEaGY803w+OSjO9HycxDQte0LUC8kfCvP+eTwBmHb6+Q9hkJ9
eWRXR9HJdcaZrFbhbHn1tYqmOQSS/OrNxtgLKpUiBHut2JDzS8v+D9rYxyDeOz6h
ZGNbaWT4iTKzfWidilQeXd547LqxH9AXY3/PMjGeSVUj2VVV21835wixuVOOGPUx
/NGHrIPpFH6rXcJK12J5o6ya/A1ibyWTursm1Ta0fKRzeIgv5VsrlF0ihafBLDl7
PmcvKbeUNZyN42JeZvLzoM06jiqEYmMhRrTjhcyDhUuNaGCXrzExCqs6piA67teL
fTEvPT+6NmaK1VW/z3U1OPpAziZfTWhatW+wMAjxymEQUQ4GGbuijS7K7okqEoa5
K96r9o8+Fh+WZSTKommkLu2NBKFSJ2/hk5iEYqafg+s4w4vjYe0XNvj85gBiMBc5
X8MfodubHLVaw+UaWeA5Ple9Lj4UuokZBLo0t1ga6gHv03U7vJWiHbJwnjh2R4p9
VvKT08ZVHGPcyfgek4WSnw==
`protect END_PROTECTED
