`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U8Ici6ZKkTyvOcjseJrKfxvm3q0K1JTOG/cbDm5pyNIKOCdk9br9UlDT2M8Iv6ie
xfH65X3YQytArLmSIeCNcUTwzNViUb/DSj2fX7X4OtVMD/GrKo0m0koEpW9n79E1
38+T6oGkgB4huc0JEnwwbbPtz9APnZEsNiYG6yQuMLiu3Tq6Q+mgQDUGDwUQ6RxE
a7qSVZLyo1/6nhgcdgwyRZDzBbIrkFWZAIwH7DWynaK4C1LTfl4dM6W48X2MqSBo
hOuXo+hu9e6o7+FdSPdOQJMKchfmF35u0xRwmojD1xfKCZJ8UR6fDxUsHKgnbdR7
Eyq/6mUiu8iIzWhOdzSAYOV/SDP50QeSHXZ4USwmguahD4jJck6EEeiC6OIxO0Bu
8r14/XF9mlyVFF4VMSHCVydAmYUtg93NUgu8oxjdcQ/ylSD3OqaKCjiWmWdujHIA
RAQE3ATuB9wtDU/RQGOL4Lk3hOGBAliz3ZuJ0bhu8zW8DKia9qWaM3KqJmffqoUD
3CtrBPZomXAZte45zdZt17MqocuGvtEBflMSOB+ZaOEO0pb66yXxPibG7rSs7J/M
klMglQUU7oaHQrQrDuOXDrwrWnJJA363lpGqjE1kAGcooVD5e14IzvHy2s/7bBBf
JLqlL/l7Oet6qR9jxOywh4aXxavPCVEUCrhGxYWG8KsWIPRDI8Hu+ES0cw/Wha0o
jwx4VKblWKdB91keCO9XO1hqagn12xR5A+KAAnm+v0iRiznl7QD5qAmvwQ4kArFP
hGBy8fZSgsM9qfHAhTJOchpwDNO4yOWN70gax9upuQijyDrhUPGBKd7P2I6VH75W
IAwKqX6L+9JFKe2J6gwg7ZQ1G3wDhHGTcVWSo5O341UfXREODq4/gMzIQ2wpx8RW
8/S3TbmvzLJfunDvAZqAF9U5z8GWIkIRYiQhIBd4eJJd7kH6zyBn/XTW5fdBTzuv
Hz52WCf9Y1NjhKLuY7PQLFugepaGXrFNSxh6XOD4Gp5veiE/OE0nzgrJ1f7dDLZq
ehMskuWlMs7RD54t9eQYYb5lxYiQmoT1klIypHF3NEfLgvYEkO8X1YocKsGOmhKK
eHAABaksOUKmJcsN7BxObaKAKDDj03Uw/1K86997NyvAR33xRP0U2ZKGsViE7fZe
8Pss3oUx794lOAVWv4ptjy7+0li8DdkVdyE7PUR7xLanqxvzawRcKOWVCAoz95uX
iu0i3mXeGg0+qzNpRBiDqZ6P8mF0Vv2gBrrgYMAzgRTW3iO3xK1XAjyGG465gG5Q
D9vhEaWO8i3KNisiu9TObXgfKo8VFx0iUaWCZnvaY7/z93FZsexkBUM5JftFTTLc
LsRcCwnqOwcCpg8M96nJ3GzdoFW1mbtxchkvc6hfUw7JbohGsp220vAs8TZTWSwd
`protect END_PROTECTED
