`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bKOmOdOHc4pdUzV2Tu9a3ZxaNI/nl5i+bBaeFJ2Ggfd7ACWzZS6Lj4IwxNRxUKoT
Z8LNQzyaZxqkyjPpf+U35LhDwlZ84J8VV63kSJ3qrI2e+TrzJymaUiMJy7rF9eEa
JO6LQXNTYlwMSmHgTquntKlBsCa0ZLKJ79IzmlIFZcZj5jaN9u8R1glkqZmKV6AU
28qa2sn4mypDCrLw6XaZaYl3aPcBv7sSIskug8SELcqkWjrsMyPDq+AuLG4TcV82
/HAOHW31T0fkbV7J/GsJ9+pAjpa5Bv19erkQVbcwy1JtcVscK7Djx+kYOXuqA8W7
Tli9zyy6W6xKF0FcucEh1TAZ4YuaWXl5ZqLxVIRpwcwHr4Q+sddKMKxUucgIOqV3
`protect END_PROTECTED
