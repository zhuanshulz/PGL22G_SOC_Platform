`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5/ImOkM9wC76s20eb8LugJ70gOJrJbCtHPtlnBQdPxBd/l4dvuvSk1iPND57RGKT
9UkkQRwNwQ9qfAJMOgo4oPq01Fbw9hogxmzTSu+sKvKqrwMwuVZp0qpwZ2XfJ0Ir
5Vpu9wGtIA6TJdSwVAUMYSHbbgs6b/qnUwK+UnAmP5GJ907wHkS52zlq3PROe9VC
8p+nDFoaiLLJ0cRbNYAxJRlBRVIhNPDzh6u1ES9r/yR3yT9r7F3c0PvBVzJDbfJW
HEW5lQ80vQJkwou1/a/2keJJYEH+EwcCYzEREHCgCscwOFJIeRl/0ecpfZWRSjai
Y9tJb+uMUOefZhceaav4txoRg+Ayx3CdYS7BUt7y67LnN8pFCAKgkSKkqcYMhkXT
xc5DZ4zbI/zalkiF0b2q2VNhoZyBad/2HZkvoaGsab/vwiyCCsP/pTRcah9tv8r+
uUsqteR5Z3K6YglF4GroWLfFtVM0cW0txrPld3FpmL2cwFVCJRdWiPOOfCTj/peT
l0CKEFXRGxVjR8z7pqar2+ttWgfudjoVDpCEnDtW6evJxmuJZBaM8qEyT1NFmQX/
eeAIEGwnV1K96RQi6/JdDHJncMF5CgGow5yqEb45RfNnw1NFcedotq/AO74ud+9u
VcpHI7ZrZBtbfrduY50Zm60/CePOR1in5Vw/k73MIxiLSEYdqRFIvndObItpiPIp
49TaM0U7LcuaehTix5Xp5voPfDBIdN3tPtzXkXuP0v1jge0zotWgAuY01ZWKV3qo
LZnwhizjoLetV+1yd3ANlwgZJU33KmCmHiQQzW/xkNgHDAwX85pJEg3OXnb7y/iU
IfADTZIJ3euPCgARpEpml4HCalxD7HWCpU+QDdbuUZZqb8jQgnLgGlLElpoOztU1
O78abJW20Fs3qe0Du4sINOBth7LlFJqs36nViud6JMoxsCMaFzUMAnCRgq+8aWiQ
vgVawngHql0bTkCq1xqB4Q==
`protect END_PROTECTED
