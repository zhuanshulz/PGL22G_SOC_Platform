`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uAERwXNUQp2cB1QSQdXccAuD+GkcfahEu6+X0+6eccNDE/VXEpaEOpxCHwR1yVl3
6HF1Im7QNuyJluwlCNuBAXUDEC7jBZIsgaB1XoXVwl7YtfDAENjvAz55Z0/Hkx9a
Ej6I33mjPA/YoKNYQDKmOU4hC41VTC8ODgi/rl/BHSwMOwYsm1xIHD1sMMzxEM/Y
gD1LtW4tRr3y1ywW4mC0+I9HCGBfIbx2V9Ltd42BqhH1T05H9hGKdimz4Ns/ixAX
T/4SxqOd0xQ9l9Z7Yzkc7/8bp0o6erLl+p7RxonIqrOSM8Tlr5IHG55BaQ8qhD9O
4dP+B4gCPgM4UOnyH29PKDNMI9ghKs7wlSHvHoK5KV0M2WzEjg2MZ+WaEw6yenYn
F/f/9QITov2vQlOSkCtQXCwFIZCBBZIUPSwUKsVFAAjxt3+QHRvN+tBG6GYPfMSn
4vcrluJEV5kGEcw48YOGsAz3C9UOTOWXsoeg102gs+C1zm8lIoMj2tGz8lKokyfR
AYYqKMR/zNfTvPK9s70buZ9EgeDrI1Fi5D3GtxEY3/L/nNxUWcGXdyGhPu0iLK7X
lVWz5NFxqwqRclUQVXwPlu/EidaPBtXeKqCPsBcAfFGlWxfA1yYb+GhJCXKtAVro
1qpxFtK4dIGKcCnaMqGNzjYARHqS+VKGGKpbaYmzDOM7XFr0T+zdSeNQW/LbvZlB
LjrcUoYJoNrBNC8Qal+A/NJsauSJxaN6nhLYUVEfiSUODKVogUytDgCw96o20f6Y
kmlf3FMTsdgTWDml5IXZU9lVLHCCoJl+h3tgu3OavosUGoOjHpJi+7h1bo297cYB
4ey9Y/eU7HPZpSKCzQ/V69BnkVQXKcYIWnhuIdmKL9p2npxURksxGN88qPRQ1xf2
jdiqZ39UUpWqvlK/E4nqJJXMxZ2aw1a6C95EBgKZo5inCTNdq/AOXIXWkGcG4Qbq
WuGofsCzeQLW7ZhG19+a2lODJgNhaib6p9o0G5onmS9uyV5bWdW3UtF9JvAQ7w75
7/Nz+GewSfKvV45vJJZOlYXpfwuYkS9P92Xm53BfjAHnr2GAjAjv+LZ0MOLLc6sh
UCjPSW7MtI2LU/PqpT1Scxc+kf2iImjiW7HuE5wLK9DVaAeIsRl1olubMd8jTMYK
bnhnL8PBtQZGGBKnG1NVIi1hwCpOKDb7j4Hd/GXzCzXuSOM/jdXA50apvBixJgsb
MRzagi2yfC4GSqlCLCTWCuhVj0MZmwCDU8wNEcglWJCoIBQoa6uMcqJ8TVNdgWY/
xhB2tKbzQXCGbuPK1aYQCMtZtUGo/6zA/iPE8VmHrYZ58IkoOZWq2t4RDLj1873r
UEVFdqn+oRw5vCPrYHeMSsRrb5J8sVmpeEJuDWfmknHf61QpP5164gs44QIHvhuK
1nQFqn5abDrPR+OPbqE1F5PSLT4B0pjyewtq61hIc41nLWlzrC791m2yh/sMR9bj
B39bci0kJQiB4ZTwf1eU3K0KN91ybDQKOXdjU6KnSWSCJz4fVmKy9ZNMiTw0OOOv
JN6DQvXScpOF5t4jacF7rUYa9OfHrkzvdYNqScCFaoa/JGhO/xeLU3cq/1qOzxk1
8YpNy1+5/pshrTJUVu9nhwlQh5p/2UxQMa+NgxNoyBL5U4kB6Jzxt+XthQeUsQ1C
Kaeg4+wZLJ3cGrulAM5WqiHjtKHNCIdLLLhveCUpa5n4u3VcKKPPsoTowIgsh2gy
7P8fhv24CgeWxa0NCdW+UV7KXN1oYJoBpWQKERKcjuFWESUeGhGkfm/mOfaQNwJZ
t1tZ9J2pivpwYempiCtkGVJSAD6Ky6d+w/gQT20RKmJvDDbhw5b5gCuRP3CIc7En
y1TTHGTaFRWytdV62q1IY4YHr2hI4gy1IcB5i9bxZDPjDbcaqQv2Bj+7e5xpSE5X
aL3zC5Km/cETpoP2krHb5fuRIcoV1Z//stKrWMJHFqYQn+Dxtx3igA/UNV0mB9Hy
oSGRUPdoOz8tVBLh2hdVlH0KOujaTod4tW/DMvF3kVzgl5DK+6C/v5aXLi26vsHr
JEnsGyy4F0OPrYf3XrgqrDZ5xVtX5YCe2VMCoVd/8WXB0HNIKMRNlnjgCKHHEYPz
VoZX4WplyBw6kmf5ERvnjESFt7Z3RQ389PF5rm7eo7YLODngKaNua8q6vjZvi3KJ
loQx9BpBTaRIUcH6UwWwyqbWb9lR9u+48E9SUExV62jRin2sCOo7r0m2qUHGWJwg
o63hRYZEawNlpHb6xiJRBnvuE1SrxK5AAWhPUOHC7rdOAfK3cPzSu+CHY1UgE3Gc
WLvEr9+7Mcb5v+PXOf9EhuReCpvvyhlQ8Rt0N3U0QnwqBZG8PWBb9J0hblRKrBR5
v0dpaPQuqw6mnFUmzKAPwU4ZVsQTB6Bogm5dtF9klsh/GHBQYiCDUkYlbrfP+Pa/
lpepJpj0DuevP1A/XMzOgemseozWAU3DrZK5L/T3wD3r9LPoGOaYUK59m88R6zln
WPkEcqVHmvHAwnIuatvGBEgaX/dvMviWzIL+WuoCT7FFL/yZHMlb9sLhIbFUQIaP
pdZo0zKcps+jfTnntCy4k/b/7A6OBboogxvp6Grw/j4/xF3nN11KaZhWF8tRfmPm
QMhCTwyqlEUnBU+JvaSMLYOAjL+tk0j+o2Qo8w9qWAOhvLTE03cJy8T/mItfbf0F
0VaD3BgGS5Bx7DYYWC2kZdbfocdhlXbnmlbOZpbgJhIF5PKkLVmd4jwmSI0A9LM5
2lRQZXQLtyBeBYYKMFnl7Z5ZOo6tY0Mp/lylRuT6PLKmiPgYaYaCz0R5W56QBxIk
HLdh+hb30mX44mZYgCh33UwhXaHZasMTg9vKy3NRHF3zQPM0mQkSGzRSvRPQhEhO
kaDnVSHnwWY8bWzZjhm/SQ==
`protect END_PROTECTED
