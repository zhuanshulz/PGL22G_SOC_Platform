`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mE1rDyZRdtvb42yUb5ZgvBTf0rwDAqn470Uyrfu6WRm7rWK8U/PrUdj7H8uQ7r4u
39S7VLG9Cio4kRXLzipZBhMCea2CSqWa9nndmDC0x70sv7UJLDl568ZBVzWUpO1m
PL1JosCEZPZJsijbRhUOPDVOPaJRTsR/9zSGqIS08mQtABoRE7uGygred3IoU7mP
3odOXvCZ1t6M8lvr4KwhzO+HArhl1L6v5CpSmzQ7Ye+z7B3rHYD9WlAlhTadmQ7Q
a1to5Q+Ki7WA6V3jxFfvrb9+6/0v+oMgOOmAL9tOYksbB/Xm/EG49KsNxwsO84JJ
v/8Y/J04LHK6o9ew/4Z9y7I4kAVoA604EYRx8SuWXSlCzlqNISLUVVihGpObiwnV
MzOdiPBNUdXZbnhRqBFJgP3uDQgyKTfY7guA5uvd+d+fAtxINmX0BPi+LpBj1ZCa
U7e663t5xvOzUjkdqFP1L27q6+wI85o6PFFPyT406jNm3VXzBpfTN+mTID1j7mb4
I3CltgeLpX/bIqG5kLvzAFKtyxIuf+g7J7p+tmGsWsfZxZjlJeQGo2ik8POZrpib
UDLduv/TSXZWzlauJhurwVF5KZO+D/cmYW5labZ3DrHvGq/9s5U7t1OxQyK9aTb1
iscnLbkzWwk6hvFTMfOH9lapwv7cpOQn/oiWziOOkfTbD/YPw3oi+7ekWzZ2ytnQ
BenbstUQCPJ19VyKufwit9cwyK5AFwoNgkswVKob8visEUjZG5JL2aYCffJBmhOJ
buYtuG8cbJ0yT5gZ7YwXfzdz5o6TeND4zXSoHnW2oR3e+X/Ldw8/t1Cj6XtvIPpv
JjYfsG3EMeBxrWLzwnm+OF7A6edNbLNrTvT0nTZ7VZMJwEABi5lfzFA6bMFRPXY7
Uk3Vx58t00/aHERuu9dHWBMmGXS/jLSCYSeKyIiGM0xSKvqcscwqlE78E0geTjPh
gujQ7VGwBcHmhanLEb3U5pWuC7RBpkf+0lhysUcfsCdYgjIgt0KHJHKmiuun0uer
aPrs30AUBbtxmD7lNdS7gAOdbXsbY+3IyyFuOZ2Et82tqqgwHzxvxlkhBOdwZGnV
ontA5pGmKF8XuvkU3OrNilvw0e4yTGAK5RVAtoGbo40wYmcIxXEwMG6NwUNQ7K2x
rynxNt6Ts5My1HwkZzguV3uyFypN5G7Ar48xOpCj5XUmNlZgRMLULMSz84k7fYWq
GOix7GwbV0ITwXzXGVtedEUZQWbSw/zQt0SIj5yZJZxDLlwzER9DFWsG58FIMO9G
z5pEGEAWpE2d83RFbzuXJxCJaM8KqLypoEIKnLkU3a5RNQH1NuLzkr8vT7tmB/gK
ms7AXZ0Y5nxi6/sBh1gR7EH8I8Yg3SjX6EkGHv99ujckn7pHNNeShxGRJZT1COIZ
7cVi3rXko7YC0fPhQeqO/VKWhbUI65lk8URnLUBH7f+31rgb3X5y5Bx3+WlEnpdY
fw0vjHVbnbab+xnvaFL7cstsYL33GHSZ4n3y7ZyEfTc0LdKDyhycEHrjICno7KB1
tR715WlBzV4Jf1kBOo5zGOn1wN2QuZ5x7UPT8n3hln2UER8g6HhuXcPD+9CLnqLa
q7XSWSOSRxjDIrH3TF52BY/XuBRN529Yz93zrelShOiDlVKweXZAb/AoRX9zVQYi
uOlsE5GoinczoBChs5XSXJQF27EGfTeLWYEO2xeAkXH4z0fMNWRH7krqPsgiZY29
RD0TJxKtVUXg7zm6q/DnmiT+3icgu9eCPd7HTQKdnHZ8Joosd531aqQmooHTQHtW
bRdqU3g5D0iots2KpjBIr5j759yeMdrw7DggM42G1NsmWhpjKZaWMOWRcHFhBppz
HPw2B+eMvVBXOBuoRchRZs5J+DHCWqRh0KNEHOyMflqMa1U5YOE/yVqVjR6+HbG2
BLQD7tlcpSGg3Gs+x7COpMUNaPe5aHA8kCUTm/8YuGXByfsWVPtjn8chPS0W5Dsi
Pay4MOOQXXZ/b6g/tT1jkC6OOBAiTcJPzsZsgxL+rK9gnhV5vSwMvhZezksFoF+d
MJwOdMOPACZIs4FSwpLKv+fOYXaS1WmoyLZlID3zg6NvgfUZUbAq5ePYpv0fGgko
VG0351ey6+EjwjJZH+Pr5uQe/CYnQst0Tk30RZ/ntm+RiiQsuvnrr2vjLMF9W4++
YkIWHpVreb2ctiyGEa0EsORZEBTvAoP7Ych+tdAX++XJx62oyYHOwc9KvUy0uMN6
izq7lqylCkESqPodLre6+IEqe6MBSti6vr6kNg8z3CC1nfrpsPyloP770zoYm5BE
sjqpMUDZlgpjAnel8HdfF3YKn7L2M7eKE+CXnPeX8hLYss/tVc9dLTs7IQj6dA1u
eYSn/UB0w9BifGbfPKGAovDJZSeLCwLdD7Z+CZpWfpa8agU64va9NH0YFuDJavi2
F+pTTYJv+2IDVfzKaGMfWet9Lm/fl85jJwqNzw5MFN0/fWZfWBuBhGRbcFRxu32O
7/IlbZxAKjapPyuG58yKNW2/AvED1hj/570KO1LGYbfmeamidazBScmHOi1IJErJ
dWVEuLjCfGfGdUpm2FCK/iEhmIPF6sNHWzsYegvwZtEzA+UOPdgz0elBZ5N+M15G
S+3AdvfmdSrQiasSVo1tsTqjiGazxE933ulq8qMNDaLraJ00Ha/gjMvRe1R+WKfD
sR2naFFZuHnwTrcbjfFgLN0WQSKckvRGGnSpGsAizoKhADmWfbQG0+kisq7UlENV
upceZOQwDyvsEuJw/HfJ++5tYH9iAWx8l/d8tlADJo2ZQGUk0Z/Nb89ZYAq717J+
Mo581v76yhNl4USHpc+/1w==
`protect END_PROTECTED
