`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lLIMvlDkJzp5esarF0cklNdrxGLrN+UgQDm7c+wDBzbXGjg1wsOIXL/VcCZDPSbW
s3BOeuGW49ofWogRg45T8R7MpHDVil43njeoIvcmG4pFE1TF16jPUir4i2hKdpP3
p7djZs8VNsbzHRsRLllDfmwqwUfHV9Tsx2iAluMCRtof3UyK86xH1qfBTVAWTYpr
/r2tgncj95T5rnAYYlLn/ZQWjJokeb8eP+1HT2uKLMBFYcAVf5gVoKMJC85IJlB2
u2lYqqHBUyKmBZZ6lnMgjfKkryKJRuMy0xbRjHaLgjUCSzamm3BMIMf43N1v7oLM
G67B0KWwUEtrnbAH1lI66QzRXwVz28bd7Wa1qU66Y0c/31ZircJGKyeZ0FA9uG/o
RoFKchhEuE6X6t47znznNg==
`protect END_PROTECTED
