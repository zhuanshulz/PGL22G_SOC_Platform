`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WyAZn8oKlIbuYzlCCRQcZwlwetOoNumWSPfa9ekxPEobdxoChZe1HOjmsIj5wjVk
Akw1Iz0mtTqQC4LACPtza0dk7S5tslY/DXblkCya8n29l79Vntdl6LiOgt4ZCKYo
1cKMwuVfZmv+jNvv7DSgqb6bXxIBDN0mCziIrFV7AmhZFBF9fMgS/vRLhUJBuw95
WbMyl+xg3w8fTHFRc8wpx2t42StTFzcNti+zXu4KAOngWcyKdwRHW3v53ODahImm
3zHlactqml2AgcQkQy1kB6t4LKvlJt4zvBoDoxMk6Bkn4mW/35htYHeTrLAa91Op
LOFd5mX5QsuTqaHBe5elUMNNjgAE/JQh6ZedUwK0k30QHO5po31VtjxTu0LctQIN
cRWVmjTNoR2sPs71porh1Tt2J9eXfDpmVJQ8fEQ+fa8zdftZN1k6lR4dbtlKALvX
5IjYyDJGoJFjIs3ahfEcWSHEgNEKfNn8bc7pwdjugWx6pOqJZjt+eS+IR8jplhHv
847eXNfxCDsRke1xWFPFyRbfEiiFC2xodaBrO2z0yxMAmmxZhrP1FafM9wwJGk56
T2gli02wCP3q87xIQKgRR4kyDzSqjeX7MC/L6pCNkDz0PFE1ncB0Vs2X9cLA1rm/
i7nQBkWXL6PcJyKQy21tYq3m8xZBEljihx0Wcuq2J8+KD3riVgnNspZrqEpKwrjW
rsIQlg5xq4vg6K7kv119Wau5ElrgmjKv+ObOuuoji7bAtP72yaVB3SCtChNvzi2j
aVFwV9ttfDo0Uq+Hj1O4FDDzNt726Ws3D7t8iv1e/mwEhepsG8/06Rk8ilpXYhY+
WR2Zsub0idkO+CuccLP+1PBnagtsZJWzamVxy5oiNf8scSIYgyfN5E0yHk+UvpSM
mldc5dTyuMNaCnQttJlIM3AS2n60OMP4MRQYoO3bYHwPxZ0cV8jTQxdQyIvIsVK9
tGa1Ar8dRNLVIvvcrKpkk+97tlzl8ADygTD71f2l/k8CoNct7gQkhjApF34kzqQf
7COBDrWnVrcklS4ZZS4bQz3xa/1ndbn84WPwLdhGBgU=
`protect END_PROTECTED
