`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8n74HjLhQ817YdO4y9wW4kkDPvwukqpxIzjgGGQodJpCUi89g9zod66p0JXPfFlW
X3YDd/w7BP4HBTi+/IKNuKqcz+HrBIcd25ik6XHGc/7rm+L7KJVQH5MqNzhkq05m
nR8b+0WdakpMYBnjaYmciKHxoKpO2JcH0jGyK0ejEf5tjqevey+dPAj1iRyRry6h
d7iFpaihW5U+nFgqPt+G9oHsnai84RCvry6GpLtyhdBABNkyP+5wbrKYVXICFQk7
jFk40CkOOd7nPN9ss/QCQ9fZJ2s41nI7GokdBdGH0/X2gtxPZYjfDbksnsrVKTbr
8BwvYQicFNrk/WWbhatQUBNCIX1eoQ7Ohro8zIcw2cA=
`protect END_PROTECTED
