`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V6RIvJBqizhTJbhWusRXC4L9rlyJnDcKDZId4tRXM/MzOCAaqOA+1qehLm6dMTvK
L3v2L1OXYFAh8Mnac758p799opMk983i829N+cp1ryzEA+zgWYnBNax5WHMLUNTa
N6wull0xOC0JU+39RqfCrxY+X/jCjqfivb0RT/yXzxsTJ2+KSjNPU9ZrtWZVQOuV
z/O7C+NMAQmiKg88aQOFhLOQcxNzLViET+bPznDB/9Zt0Mf1wuXYmFpQr6x+Jo7g
oBy8iqdCMgkW6MALUmW+FSkV8kWwo2e8L6VU3yRXNBBskyfewJtLzDI+Zdh50P59
Nnv0p/TesB+dEDwR8TmwYT4meB5uo8TJ4aAa8DrRrOKwir+qEAF84p530GOWKq6y
afNtEebrhQnAhDeE49aCt1azLPtJaJ3dUy91EFbGTsDMIfn0dXttE2rqBS/jzeHQ
TGYKEadNNWi79+2b74v5Cd6f9IEpUBp1xjXAz17zUzGrN/tHqFyfOm/hu/3oeKVZ
+QYKykvfqPeVIg/GXTD3dAl6dU/0OGDEC0HmvHqPjmLkeds2nKR9Cca7727HpF/z
2WsHFUXnKk0sdwspJaDcXNvnVNU5yNtAf7xOLribNCu/1WBZ2UmgL6WM89dLAsPc
X9IdAxVHPrx8H44OyPXqu8+34Mc/O0JIxBEM56/Ty3spSP8uMahKVbDmgOfbbsKn
MriuYr0j2e9fNOG05ii00nI4h4Shhbo7XT8vk/UmeDsxXenX+agFsvDWdD0OLcR4
3X76rf/nz/PsvSQthQrvKqotM8xzRd6CHYWhZ1pQdctAY4YiEOMa6XxLAF1AULRq
BwPdmgjuixLJKnoUahRFaUDVupPIx2n0PfUVn9BxcfMaAz1IE/Umrp7FPmHMVuf/
BWf6Bk75rz5DEznm9UkTEEj13q33J/adQGuQtU/wHLI4kCaxsjMmx/hqTBL4srey
`protect END_PROTECTED
