`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pWbM57XYIwN3wp7SYSvPDfacUvh4QBhiWLSVqyZUI+1UON6HIedHaIFncd2B4a8C
rUXG1/l2gxhpuTc6phG2LsfVuAvjEQsve92LqkSR4GxUG7IPdJDMZskTXq3PzbJ1
mDeimEE2gDxdSEYZsmSmYB7OfRba+71jBl0n8VtecG+o7YmoBVnmxjlxn1Kh+Pi1
p4yV9aBFulUkfmZnHX4lDZ/3Z+iUFui1HWueNcg4Zai57GFwWpXX9bInjuuta172
jb58M42lT7GJIBe+M/8+tiiVaqSS+Jr8IIz3XSD22QslXrx7Jd6CYhXc9IE9XA8l
iKzN7NjzjblCeJfVaMIHXC0dSTlIXDTC2XG+JGw/YibzfV3VS8LSGhpjD4542pGy
65V/yv2kRbFqeo9/gM9/ppe9ftEM9GHRlIHWj0qXGu5Bwkz/mKfu46ogdmMt4sfH
9WaNaQ9xIdu+mktY/wKdOw6Z0Ur8xUtkIPIJm61MidzJzVxBCC9XIFME2hHdHZRE
JOzmHmRu9Pe/eCCAbdeDNg==
`protect END_PROTECTED
