`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XxIDU9X68BIB+uGvqTs1HHhcdhfO/AubLjSU/ov5xYNCwNW8Y6fVjeIo3o4weQeA
iATc9Dz916sLW97biJDziWUg4ScIFZFgJwA08wo7vgnGVCCLFPd3FSi8jr8fX5j+
HsEjasd8BUDgSkbYdqVMnL3K6Y1qtaa131GOHHuBhKrDWa3EX9jvB2SiIcR1VGd/
Yss/5IzjaSaO/cZIge7dTTtIX4GH7+e6QkXmHi5jCCjnFPMs+jeMH/RwC9Xq/Tgw
Rdwtnlom00XKY0DWx9Qp4TuSxKtC4hHubiYbdy656PE5173XhkDv+fThFX6TFnvx
z+WVzT1gizVO4g+E7ZDQhveKoBJSRsrdgMOSgF3yf9Fnh8ZcfZZ0IkQEQ3gZXJoz
xRYm7i29OMGhuBXk6lu+28zownoZ+VRzSRKmGkzhC8uuOEHHDjPImHkwge+JrPLT
8eWpn8E1d/B9ufPm4JRBuuYUhChkJz+BcRJ1tLNOrgGty4VDChzab3kwHoWXZJg2
MZL7Mf/24gI+mB87tKatqyf6VqJyj+TMAS3GZ+YV+N6R+xJf6QNPuPjpBWj7J8rb
HIin73Fb1ddDgfO2bWhGln83rPbJLGbZG+cgs6tes5n1f9FwRL7QHUUb4oObAfNw
UAw8rLRjz3UztzK9+Z8ZeILd2yLgryy5avfVInBbF/m0YqKIvnFp6ZnQ0QqBCjvG
U66by0RBOMXW9JlkBSZeIZ39SiNvqwOiGHl3tC/uYoqb++bQsvFdhgQNvGUHRPGO
uoizQyQUueHasVanpsKVEVCTMKVY6hXDlDLAS1Yr2rnEexiAfqMsdKE3cxaTPhWJ
g+8CzmJrbod2TGtPUL/tfNC6Ij52l4wfX+mVFzVT2wqpm0SSADD3PNxr5TBzUGjh
MlQtPJGtO+BlB++HQRy1cbRS0bUI8BF8jPYBvyHu6WG2WbBre3JNc7VM4nAohkhu
THXbARUO/Sb6MlrctufGfvHDOura2nO87HHr9RqD6dw5Nd/fi4U03c5mYC8z5/ov
99m7oG4Xntl3cyF4EwuGC6tpZt0yVBx9FQtVS9r5eCUExNmaFH4uUqfGfNdbaL6G
U7RSPkGaGahex46duTZ/s83VoeHgl5spg8skGoVQrnQp9Zim6iIcxfxJirmJLmuc
FIylJZKixL1d/CCbt2VXM2+EZpzaR+j/lGGAnQAobkwEQjGwQcTSpD9GAI8zSw8U
JBNLDT1b75n9cn8d2YhrwPUTXs6wMdbTWoVaYKcPy1ebH0prnBveaEO3AaGt4jAG
xG+07Iosl4zHN02jzU1AWl2UlVdmn+jlwyJCB5BVguEUfO9Ojj52H4aVKM/1jCs/
NkVWDrJ/QP2XedPFduv3JaWu+YOLKqrr8++9pOf2oA+hXaQe5CiJC+Yyr267hOV8
+aYXAAtn8gEPezMJXz7Vc27JeO+EMMp/79IUYCzCFmQt3wJ4VVmFrE48j2rSRFEO
UxDvt9eKf3VxwEPMHiQkyK1r1j0D4N+A/75VY5XbKT1vIEV+RWOIVmPMkdY2iXiY
cioAFN7Wz+WoU4ODqlGZjlG2jfo40tlb2ciG+CrXVKepTbVZyCDjyGy7+zefA+iG
PnI15Kc9B1z/1ov8y3BTyluhqy07EJ6th/w8wKSsaqGsGyddhxaoWsbvyPnDrUlW
S9KeKANE7boJ8v3HWfrf9bU9mnAtHWdKilMzESGLpM36cKU2/SkxAyBfFbolTdHg
GDbzA/SlmAa01wa6+PTcqIuBieu4QKo/MYolFAABsZQ8caiMxUh1xWUCTALpjfjJ
l99Pggo/g636h4LlACyeAYkNJy7G58PFVyx3OEtknrxYrDcN1O/+ULNLnmXEhjQx
aJZq60epbkgSX6i0JSRt7FkAdqu+lnTP4RQky18rtNEwbz5thUZ85TPkregFhxZX
uWvZhfeXom58i9zh1UA7usDbb7oAf/qwZnxGaVbdSksUJtDzueU0cpvUF3MPWFsI
XOHPhEkF6J3u/+Uv9woRQ6P8/NGE2bdKsnm8oWbRsESeSFbln1FyG7GYX4qkqtgv
QcwgDRYPWjLtPsl7MNjXaIQL2hpccTR3RyfGfzGBptw6XH2o4bNnE5QcKRqx7lMw
3z9ICt8Yyq0xo6QfohCgpVmip6hIViyif+1bzbBp78vRm8dhLFjysy8gFc0kxAc5
liL04kzJPvbcb8TWNhhWPMS9pVYqzDg37MmGTQxeDGIBMFfbFLAtFdXVuwV5/YdR
SImXofTLSvgVtmboLSURJ29h8nwo9mT4Yam6H9WXFmKThZ+G0JKOiajxXZWBNA46
JqtpMa4tPvpA4EnEvSTH2gsQl00+vmZZh0ZBNstD8GpcG7pf/rx6Dn3WUy0eD3Gi
0WXCa8XG5LFpVmAxoweH8rZ/eLNAXVNuMlxhOgoZjVVPF58V/5AYfo9Q1RPz3Tu1
CGfQA7FLOLd0HWJqLrguYA3xkdsaFbLr0Vv+Bcf+t7vmsBCok/+IeE/Z6a4IEZV+
DegJyW1c79UmB7uus3RXJsnMam0EgkEKf7jvP8W4LIjNRlf1cMMrP3q4LJgB/hxR
Zr1Wngtjoao1LxyLt8wsbLM95WVGSnDX73NIfC36d+QbLgj7S+mRz3yow6bb22Uy
ijXvaNdWv6AJ1zp71/MxQpekm1f63jzvo7GexYr8OftNMYxJB96bH2ayc95ItU+M
YkiM6eWSBxtvxCnRPIZ/j3Vwo+3H7tLG2IJFdPmlHja4k9xMQkJSezpiPPAsb1oh
8kkj3gPz+39Z0nTGX57/GV5yGfqb0QUBTRJ3wAH0/OUL4Vgkd+dHiVvyrDH1xGV9
qyf03tvTDQmsI1hTtV+o07K2pwAD1StyIqj2Hg8nlj6DL+WTjfeexDu7O+6/khSx
gAJf1qE3F+GUpy2Vw8XMuURzeYYxWgcbURGU9xraC+UF1+YFcWPBfsnB2or6mQXW
`protect END_PROTECTED
