`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tkc/hzOGukP9rNdgno+KaxXqZF2/xo/k0Mqos7dZIQ/zNLN2tQLjTIJQpxLvl6UK
0n8i9IGlYapSTYeR1A8AYbEiWgXGVNQfZJ0xx8ky/EcHMMATYOx4+dF8cauh9dRA
K35lar0CeJHk/loCV+bZxm1SEUbMP2N4tZQV3nH+pAZ92LdCT6MkzGWK0Jgfg3Rw
SPXfapuK1GiXsNlJ/d9h6TQAMjMwRU7/UReGFOH6xQ4HNUynsjlsfkHEMZ8nN0Lb
6mEUbqNeoMLDYhgKfPg6ZHXW0Mmh0cy7ohpkDL3+jsiUUzd4Wcas7YaMktPvOqmD
ixb8oXRXMXQBz+zs3iMglWwXWpWQYzMTZBgmNGh5DnUSWaW/wn5kroy5Km/WGlzg
hc3YrWpGsSEUAI5sf5xpfmPuNfObpKhCAtg9zYl5cSZntTUSY/A4JQMYjQs2IXLW
AIWrZTnkh/17LxYGrTMa7QSHWZJHboLmqucx4Jrs8+jHETiywwj3NIvEE4BaL7m+
3ElDaKxzvbgpfeJBLaDAW0YGd4c8GjymCpKIWoMAqyQu4TpRLGyg2izjLgDYtVd4
9X1IChmjfdIO9E5JmIwkxsw41sIsiDk5uCFRiiQ057HtA2qCbLV5WpgLxIVwHJXO
7KE922dvFYgsgujKHxjxgo0Z8vcx84zOIkYFPsrFrMqGHd4C74M1m58xEZe2KnQp
Lb6Wkr8dfom/KZi/FbEpHDZoIy2GV8V0MF6eY87sfs7U9ANfcObsLr/41xpwt9fs
aKCMXtq1bKpyJ8JbAk2p+EMpMqwnMA9YErBL7D8D3Vd20w1KAHaNBQjKHrAFOoVI
Nsq9CFrn8l64vlLxyEiReIv3JDXQI2TmvzebCeSn9kjDBg6hFdO83k820SUrgE7L
xdG1GeACD9pAhA1qjtSfk7Z8PK4ZxR0MUaka/QiHvwLXkVEmyw28o1FPrk0oR/7j
GKTANzZkImB8Sq6XxUJpu75Rk3NO6w31j5yzNgX0I59PxovkI7XgNrTB1UeI1Boe
dUuTZ+XbmK80rquyecObv618Sv88D7NACV3SAtyifqIpES0if3jCQV16RdwA6I8o
9D+iHZDM8u068O3FzOP9GfjFgO1Vn3hFVoyf7oWuHjV5gQYoa3j8lzYIaH9zvLNM
oQhIWda2XEvfbn7gcWgkOe2fXVnNLrWRR+VknCpICi2AqQq2HvfdP3qRH06Ns4+A
CacPj5DS/Mgd5sl019ExnEiw7nNVPoX21CbuQHfINzhnFYffLNZTgbSyGKWQdmM+
jJbYj7v9K6uCTcZNkzcJ1qy1niHPsDQos3jGuXW5f9Rvjf23MCJzygnhBVsw88wc
UACLF5trHwGOAVKBJxWOqlGNR2CER8mSR3Oo2hAiiUG5TjFSP9aaY9UwI4gbr2XY
sONwz/xREY8L96dYjXn4rRp9pdPi37Ie1kvj6Uf+vrSBXBtCBnsiAN2XZiRMHpT/
CPt3SvwVH8cMoD65vwGpfFFwPACKsl+xcG1Mtbn7kKoT+mtgFtcgWVkAMQQlsskB
MhGjoLRo2UYpYllGj/h1jqzDhTBKLmpPRDaVGPStse24xC0s8MuMBgE+A4UvTy2Q
4XYa1nf4dkfGmQSFoorjgInshksoocGGCXhZ41PgMEuh79Gv25GZeKMTKrpYYVRt
Ii1dcRgAudnmdiyIH/MV6FDRtwTDjomEXeey3M2/G9yrFI5vHBwQ1kVSgZlQbHUk
NYBenpX0IpZAUAZUy4h+poH5+3JYnFgJWjbsKnv1EeYB5vOwh8pLsg2dqlfODWC8
QtN8v30H8Ce1MWiqQgjcn9A3lti7Br2qV7COQcIAYSLgfH8lVvmvhaQLWDVr3B4I
nWCKftEgumccXJNtq8Z7Z8Zo0yB5EDjnWdGTLTIPVJW0LNab7GOt2zkQg/nKuF+i
jUBfPKO6uH0om4GN5RoUK5+GpSBCXGqzf5HoySvRRqIXFDkhhp4OUEA//ixW9jl2
HKKpwl/WOytYmqMkJOICPze7aTe6WB+My2dPgEewckohtUpGnvM3VrrizyCqSiF7
rWrrT49Ia4we3hb9XKhzSNVtOC1jO79NMyB9pN3KUDon4BW4R9yOR00XSacJuNwd
TUCYTNlsbJRj5beTwyhuq5wPWD8UGRMwh8Xfa/OsSx6O/727o5y1Ixc7h/VvXbF2
V+hKjIHD4vQwyHFVXT5FQVTCJRgevqHZFyXhwG9NlKvvN/6JEefMnzclLFFbXnGz
RG/zHGD2VGMO+3WGzr2xFBvNQG1f2c32Sm7jbBvtjDiPdSB8jeXSgtbprFe4o0jR
xD+xJePl4aWRr3bs1fiwiBB4okp4TOo8/DbDATCTC1i2uTlaY8VPaj/lOo7355Nj
DwNrIXCL/++U6hOJ+GRO4BejDEm+egcWv38PVNy5sj5a4Lld9RUWkgqsPuwAsBlK
VSUtAufWJJ8Yzq+GTIIyxo8SfR0K/tAfeFnzP5OCPDuYnZj6y7E1Gy9V3x0jM36M
gwScYG3LGWLI3rzy3nB87GZwb2mVQTu0P+bjmSIa44U00qH2nEibEdN8bXNlfs8f
Ovv5BoD1Bsl+Nv4yQwQXIIMvyfKXCepL3I/jVi8vZAdYYaY4Y7vdqhh1ZGMB2NFC
C16xgH48LpUwBmp9nT1Cd0W/MGiROeiDvQXTWZRhjSc8MC38EWn+V4QxNtx+gUaA
dUeL/gfgz4acN7JbQwCtvF8AQVYY0guQEHaMxnctuBpUaJ8YrOSLyhWFWVOqqt5+
Oklvfg8SkZYjpa8As6/gunF/qJilIK9jXq2yXeoITMTyCdFpjYvcgqq32nwtgjab
XvaLGB1lkymMMBmxvfnB4UxKNLnN/JlRhYM5q1euXidFEp89qxyY+NSGARC3BDEP
mPSN6hx1OptZh8ZWWCBlhv0/p64PWFZ0Ub/6ElKsv6KjRGpSHLm8emctEsrpQMAt
MNxXoavRyM9+gfzOcd0XJ9+tKSRKlbK0aDGJC4T46fJjIr3X7lATHG8ql96SXuXV
kUiLXPuvr1j13l3VXinkVuEWGFO7IauTUO59j5oqGKwoaBuz9CVvmJuuQtwVCdur
ZlK+TTGkfwkckeChhyH0O+MgKkQIgiaenzpf/HOOtjaN8ICvNWBn+el74jJHTKfZ
FDeLmKMn6gKYnCDiF88j9UVwGdghpL7O+qgeBI+8OAGN05RAfVfXeXg8eaQ2QqA9
SWHz0aB/J6eNzaziuPvksBA4WIhVB2ueCHQ0/EIqny3Sb/LmQitQ2eiCqfyt4oI+
fRH1ctvlSTG38hKfXwi7koVtlyMll1rbmdrWuCLEKE0jNs1XqXunn+t4TlkoRJKh
TqcdR6JcB1nzQpUWeqCbY/Wz9V5ocY5CdBGm6rx2GirR2BNkmEmMwWO/SIwCjoFK
9Hipw9mxFsgkcD9B5ZCbw3kfNWvekSjeKpH307Y261J+o+AGCZ2TaV7a+2WGVWQA
MrTSmNzWESUF5umFwPfSXdwP+gdTMRbKjlgQNp0kSaHe/PqGVPvd5s8/l6JndbNv
pD+mq1ZH24blak6MTepl5743r+WC9DMOIyAGSMtn44oWhN3weKqb5ZU0dYow5eye
fAqTUwi3pWPSBeaY1R9AgdVq5v1C0FhU1MPO6/R04v7D96qq9G0IF+cA2V6syLu4
nMqgpuuL6LuaQQc8ON6AUwmGhvvRZnB8y7dvoT3C6vycQQv+GOujyXQk8M8Fl4G2
og51YFZUQxUD3zPqZ/ckJ8bcqsY3mgDA5/RVkO5acg4Jt8EnVEPYn3wn5XSMFimZ
m2Gqq7O47ehH31mSJTYY0FgFL+HAqwU9YX5S+sl65AYGXLBXJUJwY2ViM0y+Wcav
42H4dklGMeTqLLp4CpDnW+GA2cx9h4W4Fdoc4vaurIaYogznWXXE75g1/MBx0iE6
cVG+mh0nSq2xBNOHXwDlc4lVh5/XjSl9P7JTM02jGV3G7gN/5TrL990TiLiS2ybw
mv2s3BUjtbmU5AspEHZ+BucFkJIDm1q9F/jGCXoq4/+dq667z74KaYItKT1hWfrs
zFtOLTbbF8CQK6Kr2I+4XUH79OBIyi0WSzfPTJtgJyvVkTx99B/LTu5KYnbyHFtm
9xdr+B+mnvdpJLAYxmrj49N+3wlIIXxGRnjYuOxReeLyawc+5/93hB1FabSViKrM
+j9d571tslCqvREddA/XNaNoqBFWcyqskbFdoumVrWe/GJ+m2tiBBwnMlG638i2H
/j4/SM8u59W3YUlHOwAuzilhQltgAJTX0NBATCnKA7ARMsHXweuMCj9yYJ2FkcAc
ie9utshUscgBycDmTqcQrjyBLtRU7wvxibPVI3BfAQolEMTlfufihu4lYpbkQ8jT
YfMNlGr/a4EPvQVtE4ynEQ73x4eHnH+jliXcNbqIN/obsb/wVF7BHatKIdm8tMRi
ZPgW3lCz+SpjY3SGzkgS5ow6E91lERwnNEN2k0EkCCSRBCw6WHfo0MuVKuD6y4K0
zcBY2DG2Uu3scAf0f/qd2xzTfQCiWkbIKe8BU29FDnsAo69mlwhDqOI4LqJajJqG
RZkf6uLPPE+PYBkRNov2/r+52Qks/WiY6xRrE5s9f1v1aAIS5+UIsemWXJ5wDzx1
McqUduzUgScFNLTIZLKQ14IyBymVVLN3ufI7ffCrGJktj6o7YvI3XeWIM9zJoBrV
3Vno+BU35i5nPOHvGvKPLW3i8DxlVKZJfhVEyK56K10bGPDi5BX/e5rJVkHgiLXU
zuI5ALhIqwsl9nNymNEjvs2gOZkYQHwCLGT0OVFvdGnMR/vvDZQP+ca5ymyyYBF7
vSV4xsRrtYxhWfaBS97Fwt2QetKFrQ1fmE0Xj8b0/1L9hNQfrszLe8eE95CJKcrU
OnBtcqvGYm5H8TSeACS3oKbUgoTGLzGS/aHlAhw2P6Em/s/irhn3fXiBQMj7g215
AMjgwOsAL2Sq6gPz0/ZGLES5I2WlcP3B+naVDR6lyRcSIvsmMgEL2Sa4+NbWu7vz
2WgGNZm78NYvGcmWSrBrOIKsqJuz+CIf5zQEA4dyvyLyFMrm66kNq/J4rxZJlDPC
uv7XI/8dAZvWDsjftPsc8ihbEnGmEMP8gSZqImsPusSPC9LYJP8OyWw0VmqeFX0l
UWAvndWfMNzt54VGb/A4ZOzndag3JksZacpqRSTgssVrHhF1OU2cGGLZ/JWw8WBo
E9wYCGxEZIOe9FUpOjDB2Q45dbbzLzMkJcmLhuQvhBKf4gcwAB6ymH3Cpw3OHv2n
PnYRgH0OKRxJCB7SR8rBi3S2UexJQsyP9UyqKAzk7kgyq7r0IDVO2RNkIxI8agZQ
uVXNaVx6XlO6Hezklsp5HEpqZ90PvrtHE1H3giOs/Uf5+15QeIh28MLnH4k/vUmW
END/iGmb2Swq5qvMrlOt2YDU9KkOxI/iI9vyzIVk6HO6xktevGbUt3TKsKQ9DcOT
xNytrqsoUd8PcEv1fJih0EDsdhDgRIOkNDIKEvJ0fbCNAJHA5b/VFC30Opu/3T40
py8bCtUyqWn1wAPCDeilOYeznRf0eYB6uZ1A68vN0aq2zwFWimuDweaxVTKriz2W
Meva15nnYMEn4+VcN8z5YC40xapFtfeBhJXulKyDROi4rZbnhR3nSjqwOLbTbAwn
PDPxwazDvGTz2oRSjWk+5tWi8QQ/BgmKIsAdjbL3ylCSNHVG40eyg7mgOzBI+JZQ
KCXWoK+C9E8ae2k7b1YLDJVyBKE+lS3KjoG5L4VQkSZ5wogtku9pY+6nTjI6zjqq
haQQwe7gFFpscjKcfnugp7ABEdoLQ0HPhOUf5rlfNkOaNb/KhwyE3xTQHeqxzSS0
Ng+ihttyxazaAeAbtjCM/pycQNb7ppBL6QCu8cnW4rxXQWFy5llQRYG793zPLw3J
fCqN6i/KOSH2jnv6uKiUg/71D9akXf9N/amMprJR5bEUPNyxH7AqF4OOfK7xjIJ8
fOMqiityvxlJePqzqce0iDeSCXG+YajmLR4OXyNOMUNN8euNkMUwlYo6d3p03cTh
W+7BDERKdpQWa9Kj5iK9imb2TcuqzhaDFelPsUYs4sxnorLTbVIdGZ9eYQjnpDcc
GI2Vgqm1OtRMy8prbbc4KKjp4wf+fUgiLF0i6gDisMsAS36jc3nSddWghXqyZ7Ol
YEUZTLMyaQB1kpUqLHPWlJJBe++sU0hO8H5UaIrgXow0kAYH5DVnhSO8BQt3PkA6
setoOox9ztUtLd8ODZgzCa8tDodWMf3RJlXMbQoGfLLwNSojFAElKdo3eOXU/QKW
PR7/d83MVDsuyKjYtuW+7TjMQsVlBgO7WlrRlM1Xwh603wVFOjTqAwZ0mztXF5fj
+6+faw3bwQF4h92JyjFS2vm7NHD+WYve2Q/E+aZ4QwWiGOcY9Qqsa0O1IVbCXo2j
rLVW8mzokvET4gw33Hloqg1WbCt7oYFSOUA0SWF7txKAwNSHnWDJMAnxDbkP+0+V
1Hnn5HiVHk/52BOqx5QF5C7UgdjKRlJPSlk455Say2Z93LkvY/3E30D4WHAZoTPX
ArU00T06KIbvTRCLUZWFdXSQZka91FibPpeb4g9pVpl1qjCNxkQpPnOhwoXrJz0M
bwA7XfSOEhaKNUlw58Sodr7XKuJ7HJ2fc5ummaMfyDEzkIXe9xOKjq2Y4lkP8Bv+
98uVLvC6T8/x/NnGwb2Yz8JJBJ7A6HKUWo4rCXyAnFxxxt95BwcqDtQ1MSd1gRne
XDhndewLFg1WpcGhARLKVRDzXTzXx6HCocHGHSmOWZdVVCHgbEPqNYdF6fESZTF/
6xy/PgGkpQdyUfU7r7KikAxcrBo2f0dd1frieoJUz5Q4XXM+UXd6y9Iydl532x99
jRM7TZG1+DxzSNSAb9LPKMkAljNkwlEqlVUGzZS6aJGyvKaepA5M/vpjdojIyxtn
7vWHliJSkI0D6NhiYbz885/qjUGKhCZ6OYPfSymCP2+pSWmLBNbxUQvX5UR94DkZ
Oqp2DKWo85srD/Z5Ot/lTj/5Q+PefdTqkqU8AM2cmtAzVHgG5qK49nD0MiAymVz8
IM7CMCsMZHlQbWAiH4vX8e3Tr3qVcrKtbe9/d0Nx+JuIhVr5QHQEQMSqglFISFyc
pAFeyxj2qK9YkVJ/mCeP6Ba35aWzwPB2O8ADvOHNpi/ZtOXTTNiU3ozBRq7t3mAV
5RFHhUWRwu9r9nIMWBIwfa5NH/wMpZN2bFny7LcTBdkvwnL6u3Px0IIiqLC7XFg0
tNG/AM0iU7eD51y2pm2GW87HsEvemUAf+8I1egRyPrV2fVUkzIJ0JmwwyQaoXsXP
CQ/a9GZorjUTAJY//6wR9bCo2DNoSQnny8hYReXN6to1xi/Y/fadqyOuXleOd8dP
1yp+9B1do0mcwXRG2cNnG/zOJb7L8Ck7C117R4xv+GTf4cMZw1kVb5X1FlyjgewY
9WcgqszFB2WzwBtVekYGJ+zhVRjs5pH6yqqPeij2rE8hJ46m3Zrl2Vcg5jZ1SlpQ
eMThIzCAuAevt3zUJPHX3nhErrRqAN+7bl2Lfi45+FbWDvAiFPp3nCVUyh89Wi0N
/O582p+Sz8JkNqED5p54do1UTF+DGvAhUAVcc4lK57B0BfDXJKcmPU008Wm1cHNH
ts9uHN3gRZX6A1LZYaL98M3h0tmebU+p6I1PqZb7+WAFsH4axq6iEWMcmssVWXoM
TiJH6bNSVSYTiaKODVIbTuuJ9jPki/ppc50NPndoGYupW/oYX7okwk+YZmlc+THr
z5e5xINwgq+7sfCcvXmV3Jrby69frLC64rIbrjFOIkESO9M+J/Z8W5aeEzjNoL7N
hdP34bnNdDSoFhslkf/zAiGOgUZudhRUvKzxvx6N1Ye338pMdSco4po2Q251EcIP
XuilXjzOe+vU/bRm4t6zsAoi5oIpNKxLU1KuRSxDrwKVvNb0/d8atnCIxyFFSoEh
zu6tcmi8k/RkOdJzWtLQwBbPTMgKgWxUkoltus9Ho5BF44k4w2s6iIew28lJx7rl
x6jOx5PJ15Ex9cmuS/iY5LUjCXVZCV06MZYyFEVTeQm7P4KRbUT0WPmQZo9Lr+eo
kr9rgSStswSkM3Z2dXCsQnkrYf3f33MzmM1n6Of28wnEBs3tWuPdzXB77j4TYy9w
Zo4OKDpzA4kob63ORr4Cmee7L76UcVAt+RBGM06Yl63rlUVw13bjWc3sM9euEMad
cFq+jEFSOqd5t32ekte8qjNTeG7q8q8CUf0A0h6ZQ4nQ1dnNiiJUHe8PxKY5tNMM
CjyVtGpn5C+K6QfjNseMv/6Do839kXUyvOHmQTgENZrpD3h/Kusujgjn2ce/Ghi8
pU9sZ3QIeJZ+xuyLJCIgSIA6j5goA3hI7i/+Vy8HsGC4XNBpeKMIr7KzA6RRaxAy
UVAqO8fS4tlt567XD3fcoAxbfe4q6HWNlt23D5pOT9ao2c5ooQnz1q7rWZHXYjHX
EvZieelYscnuDSe7rtm7Ij/ll9yGE7NlyFq5jXmPZ09NrjpmLA5wdgexUZqZzBAx
qCd7ZQEv6hi8l1JO7SKr5OdDWvulIwWQdKVsG6O5PzFSlVAPh6eJ6SHvOmzRdsX1
DnCEY3+Nv0iZ7+PRuUAJL9meTcsqNWlS8PyRBHYFFU+7Muk3VAgZF7UsESCaU35E
RgqLwy+bqfkc5nIuc6qJVqM1mjSZWxD96QKnKYaINdkQV5glOzzgIcqLnJq0nzX/
HPc8IvNCyRMVVHxihlp4mEGb1AKeBlapT1uJFW7KQUstNzj3IzSw7XI6oCDGvfQk
PW6cxrh1hPyKnrFIxzQJguqfrQ7PAkVAd30NTI7W4DI7Q4i2iZVKvz5QFKueqvJz
T5pb9m2ucec0raZ/KAO175yGybLyY6oLgkeCbQbEDnsRjS7Ft+tzwngR6MmzhFCf
KtPvWBgKG21CIZ1QxpGLvdNil7i/LhlbbxuDDMPGhjQbvBztLWOtXh6Ky+xLeFvF
TH246PpU9IhBIOiiUjMlkr8gcy4DJYADSOg6Z6XtmvfW6Tf0iyg+8RaxcITHmbUW
zdXQ2sh7NCq3qeJq//qTzWp1hIJohGsXZuBJah1lQ1r5vDNT23ledXX4/PV7j7qc
1+zc7ealJKNFrTNbCmv/EYpC6F+SbdJcncoZmyEqyULHB/9YRMLdU/qwMTfZXiry
uEJ055XDJapQRodl7TKBXP2ub6TRUfLACcDU/LIctEs2zrVHt31iPO2rIgNnsANS
BRJW0nSLQIVt4qoGOsDsMCWDrjLPQxB/96koFuPqURwNuXUFF4rW2RViLPzhkMCZ
rmHtGxrb/74KwgqoKrhzZzByNdEz6seN0s75cwxun6JZOY4C2Zws9jtvdA2TxuB8
gL9kp6GD/liq3oBzLeTY+BtQoRXt3H/REv3InN9jc/wrsrqy7OnEpw3zkwL9hkgg
g/+rNhC8fwc0C7D4epgNUF7mutenrfKZbF2VanR+Dg8UaWYr6dUuonvOW36BAbSG
hD8/YKM7cijmPwTsAr1rn0yFrO/+3WN/3Z3JtjTOo0JjiO0in9o5/36qgBDTzPoO
VpfuRPtpir6NTBIAlJ1doG5B6hxJHCTuGmeY1nYf76u1sdIEJKIy9NGMVNDMfST/
eU8lgPu1NtCrVf/ChuHs4mpd1IN8xkbByLJtWXSQswXGBZTztofV1EYtBbPCP5/F
HjrAXR291jCttfT/ExbDNt5sfDPvl/XtdmR6/SbI0mFBN18nnFaWOAdCQmjKGJJZ
WV6PdXHTFu+DEwJ98TyWJKQ2NRd3iT9FmKNJtVEUe4pqYUtcQuNrpbziDrNesZ6a
i52RzjxT3v25MdTXwQSkUciUSXxwCUGER+bcg3OEozdHc/5HNww5Qe1FBCaO6bgb
gSiuuJEPDsjgYzkaJ8m8XaoCmsjs+wGpAi5QWixOaRdLRtFPl5HkcwDnZta/VY8B
TnYwssMq/3Ey+mexHXTsGd7fiq59MwWFDrpQXYwuEF7j8Yj1z07hYaUaleSWfCY6
MtQzyeBBI+2Vt088vLQgs+8kOJq1OESlDD9YXT9cP+wOw/9yFj02g0gdxeuaKtzj
jP3wfgwKPGrDYN6n4WE65PvNqhG54GnIZSEYpcHNIsPpw38IQ1F5EBjGWeEyy9XH
S5+8K6pf6hERPJV3BFv0PZdy4sU2LZw1KHnlAGij4YK2BYIuI0DUKtLRpoDD/oCs
tCySF+hZQk5CB/2CvJ2vcTBoxFWam/meBWe4apYD9TvRQri6ULUuEc65lfYSi8MX
k8LKma2Z44MBkKfW6tuoastjAmm3uaNArbrG5G2bb6A0uhpM3KCw8GaX6vl0xuM/
1u2ciGJwZ/vba+tfhKYHM/cg6VlY6ylrS3koTWQKgSCnqX4mHjASzwCnPmSIAeDE
/6AqgwM59O+qvTDp9AG0rTe0GGcJZB2Pnlw18m1s+VaAY2JsiAkINM6HAadGCVTH
mPceOZ4MwUHqtM+/zyLOG/L+pSn//tLZ8/NNoTOlHYAy/N9SfIzqFS6KNuPv8opY
2xGT7KA20PNU//N1omKkNiiKY6QCzooeU0iTF1/ivC+3wdkKPGFXyi8pYobhbC9s
4kXKx9FLpEfYUhuslE2SbU6+9E/W8Njy4t8ps3cQsUJQmkOFQdYE7oFy9obT8kr7
5cqVx2la63aXboP6LWqP7aoC4vtRtF5uPoVWEJbCR1IA7/o3yLKIqzLh0aNDBSfb
eE2z1l8+vtodd8uCZCiRAM4d7IhQ52oJuLXY/WqQcfjZWX7CuPllpk/3cHy5z24W
DjZ/S6f6fgl09+C9K4Te4Atex/v8tUL0fr/f1shu1kQHXTVJnzuUohkEMQ9o+ZYi
0S0vtKDWV9mipOkB4xLdOLEHXzCUxJ5YlfRuM092zQ4NKbfnJqmWOh2gQFY17Bve
6nrHHhpMG3j1Oi8mHXf6WFigppG3exRCEEMSY7EWGwOc1F3gCxXF9yHitu9tDdVD
xOfbbLw1Mi0k2LCoZYhNyvIzr4rPiDQ5dr8MYq3Lcxmwlk8xcPs9vBQkxPZZsp5s
0h1T/uo+u0AnwLXWfBMCLlsy2H4A4potOkacJadI0+ZQpzY2JRB4lTJjW3MN7owN
31Sr7yoOvqnn90f+oFm8a56CV02C2zSfrF9PNPAx33TpOAlnM9fTt7Hqn27TDAhK
JfDWrOCLo3y+u3VHvR5U0tC+A80fngJMe81FdSIg7uAFb7QyM6HRG2hhzqecRPON
aXJVva0cwMoOvzmHO2idzIFHch1o32jXM3A1cTVsXo535AC/uzvOls6E1booUgfw
Xr2YIjbP77yRpuXa2CnD/Eyg+wz/Z3LP5XM80GnnD/SCMo9ixB7csQGJmsHEYZze
al7za3Ma/Phxy/WyzmXZdSEuOtF77ylrdamPGWPiZ7uQI1P9Al5QyyvlJiGIigoz
lSw3bGgLhHhzHCm53zjaYXa+1m7eAdVcYIEBc/3DoW4sGhDP2EuSPJVScliWSw5+
OFRx+3Ho5jO73wr1lAjQrSc4ID/r/cfa2LLj0XDIlLuBn0Ct+Ptq/sU+sOuZfsOZ
3C0kvFggFAhbYqrYk2o4d979+/3NtKmHjC98HkX2v279PhcUnzyomNp1K6RkFa21
tTJBLDtFH02uti2PPB+5MT0rQtLceM03pbAgB6QNTyQgMthwXXPu9ADymWnrARH0
UM9d67eDZF37P1Oc8NNgxxJW/BEhqX485jztfa0y6VeJN4eYX2W5LkGp/dlBuEbp
IbA3gHrLty54BkzBpo78ui095LLQZsccSFaP8qT6JiMH6EZcBflHT1fWjJ7/ABsS
zyFW4dKoCo4XelNA9GiX1B06Bp5VCe6/tDX/zaF7WZPFlyqDWF9fACNagiZEq4r9
ueLJME0NW3yebuEKZD47Grxrr6Ofi5U1ZyhSF/XYapTQLpJUs6kpfFgU6nwj+eby
yFJJq6ZvSNvzSg8DREfTV7lu46RT9hCkbzpCz1AtpZiFR+YMjEOQhhAZqvH3dhZZ
haM4R9WpqhBoCkVKOVWEr8buVoknJOOkQja7Ps2WUNgkWxl9GkiaJ6cw4e/0HB6H
doNcKt/tmnRwjDV85T0+3UZaseTyA2m7Cf5E51Hl6YSxFNNjD/J4YmNflXCDtxuh
rXSm5ypkKCcx2xP8QqHSmaRi5ZuOgfDxcGSMythWnM7TiW3M5dfXVftSfTRKpbhb
mphhi/lKBtPT8k+Nyw3PEqBGgZkUSwKf7D3bg8b8Nb5mvfiAZBqc0sq7GzCPC7gw
AYHlMPBEZaBf8eP1WNBTfoT+YNTRg0P+hvoUpPjOWdCUDRata3tFDj/1FWFybPUE
oss0BK6s/qxfPy3vXKgt4yeBOKQWUxWzgDLKHrZqv5U4AoY+uEBUO33nG9TzzyaO
fvEhx2oHjnIJJ3SYMhJR/zTK0FrdpZOuGEBA+E3XpZCpbzqsbWCiMK77h/uVyeu2
X2ENYMv1meK60RTS+A2QtMoendYj5sSEYgteKrdUgKyXiJM79DnGVVkWc+JF/dpL
r/rzG2WoIfA+S+JlMKPHMp+RXqA1B+ue3JcD+2pDj4sYC5+KfSLLVtvCyVr7gG+S
h1PxYLeDMNL1a8p0lbuhbpQI8NNekM7rNTF53f2BQhnf0+e016lL9qqenfUKC0Go
XRnYbvCLAiBmur4U2TEF0qo1BlTfgjuLKs7JyJxuswGLFkvSZRAVoemqqikOsciV
vqftBRBhQucs7QWHP1gBxrd6u9bhA0RAx7Xst7BefFmqCRfCIPDi4xWVQ9fw0dNn
tgG2iol5r+6Nm3wJFXAZxkemRGcHj7j4VdU9n/ZOd0kRcVr+VunLvuelpXfaQQwQ
yhp7+C5w2Q6g2HoOnhH2/CyDTGQXI1X4uSdrXCNoQkA6FtMIel5L+mlLe0aTFasF
VLeB6t7f94LqIfefgUaji5Mm4e74wuj5HG0TtiD76NTnXQljdsDUcVlQ68zl1gHF
0QiznnLTmBv23SLYJael2r36hTMXbasx+XLNs0b+0QuOvST2AKXknFr5F+y6npzu
WJqIkBCMTQm+Fn2xYqxRzGtiJcRNE7gKWhB2Nl0CuxwNcBIjaiDEIvyIkbaRFDdz
YRD93qDGmLmvplRBTeAB7imjJy/iqG3ucqx5pRcmJ3353GXFxULiwptujy9jrgNI
WwF6ENZxNxD0lb8wS+/gugZWd/lojQycFPaCTBJLf0C4ZhY1e8pfw4+P8bR8BOfY
Y0fIVrx4ju281DEngWqFOlxu0u1DtZQcih/jIjsUsWCEBfLD2dZMyNeLL8nKf6ky
qc0jn8K8jfRcXQ14psMv9fFp6SmhdkSIrAvZssaWcylfWltoBDICFnY/P0nD06nv
siVIzHvQv+A6o5jYUk7h3fVIBisvxFmiWgNe7BPZlu/8p1LJc7KRv3hIYf8dGu6i
OKrA0l4A8+OYp8MmcXUzO1S6kX2uFJjasgyMWAcLmOojwP0sxaCZY8c6Y0iH7Iao
2ghwdsR0+tBS1tmf91q5xBIwZpX3U4H2peDgrUdjbgJU0Mdi/DNz+VCOF+Q0ih/C
SpU/XHKXj6v7t/GkORwaadbJJT983OZtsk5oCkHAzErfVoInw8WGj8pF1vT5FoLV
R9YvUjj/leyrXv+/w8JqeIqbgQLIaEwE0vImYHkdkvgLfjQP/KtHbAPi/tV+hvnl
PsO0LFJXDjlkG5ewaqTiPX+5y/gOGVDzsxCizebGetHNAMVXPw7wnc1AP+XxIPY3
0opjZZIk7iKuXJnJfFBuJEoLBNdOSLPRamZwSLxV/urhYQUu13fcHuNeZC0ofhHz
UHqZo+a8CE1sKd3Du4hItKwqpG+3eYfUuLiBBDp8fom5ttZIRBLXp7BqLnk2B9i2
LfGQIRo6JA3xvivqrbXXraK8QKIYZHA/rb2hRi22HnQbByWCnArE0mhMtHKuHHxH
eqCMrTyMstfBIxVs3tEZrtLbstlXrlJ/EUa2D6iWHm04aFDKMqQVDIzAf94/KiPu
ycRfm2SJ0EPMeQ8H6WFdIh5CN2tzMsPZi8sTmQWI/tj1ZOxNsNz5N+NH8QBX51EI
Bycz3qnZK+KkZNceQZMHGzrHmn5dlncqn5VlU9KyI+jyggPtlxaGPWXNdzbNTVu+
IGdZ0DZEHSfmfyicPI5Okrf5ZWQY8k7pBV2ORwxqQ/fEreCIPXX2koJu+NDniCm+
pRioyz6DkbUx9TdeAJM0UUXpC0hWXgBoIE24R/YJM5HaJKkymkDzc6B8Dj5Pi6eF
tFj95kDuNrm8pkTzjYIcRkp49kfT3fFSnhdlwqvvz1jMkgM6OU9MKPu++GeB+e9V
9maIwgWDg9G3bb27tZhpnWSZw5Qc1MeKaIPOva+uuxohCi7UjS+cmB9OmS/SnAZd
pJLQgObepRGqMJ6OU2PelN4WCWDRxr8V7Q3DSr/4kuMuVTxM7uTE9ThpNTEvcEz7
FSaj7+aLXP7uueo6VrtWbO6lxtb62gbzIJRPZki1WdacTfUkKaAmJssazoPeH/OD
GeUfuDzOowAkVfL9syjt1ms4uBR8SPHZ8hiPGGwvbiAC8OelO2h00q3RmSnOomJd
LSqY7Jl60eVCOJJHvaZaIwnINawZ67LTPbrIBlOcIwdeD6GosY8Bg1HfU8SYlq8A
U0KdPP4bE0ER3pJmLpriz6NiYb+olQYkB5782dyOcx6zdGZJm7eUNPG4RdYMin42
lNleF6PPnuggDSjJU9ldfenyhR9Jci4OZ1HJbEiWDFyxF0ntG55HzROQaxXehNYv
WyQfvg/XcK4GpAS59gdguHFF7q+FLaFaETHcj4UR/1lkhJ9h/UOJFyrJTjJSoj6j
15rcHEo+weYwx1Hv1WMQid8iPFA0pte6KujMBhYaEIQvpihNKiAegRoDMLNt7AO6
uO39KNvkhDsfDDOqdzKUrG+AgB/fDSsSCXAwVnNIq50U6iBslizSvpNJUzY0D6D7
9YDApUXS2BQk2O8AjP3LQfX7HmyeTb4JFnsXZq5h2x1DsccBzdEnMlD1eMkwcOtL
jTl5Ej/0QxsND0Kp7cO+c/zZdazGDfPXkRDgKazAIEASpha/R7lRvG32Y/04bwoD
APUhHvIc3xQEpMFsVimm0oCOR7B/oFtOg8sjTsZGjOHoOBOk+vDB0JNoa0uEWUw8
4tZEOv4KmVyBWhIsujAuCd1HqEmamLT0q5EV/bXUu2NDOFSPDO83M70prLtcSR0q
HNWqrmb4znQ4NVbLxNvBn9ZA2J3cE7FDOc86ZWs4JmxAXjSh5dnf1EHZc4gIjfXS
4GWWI+wuS2W+fGeRfHpv4bodErt2HfJApCn2cQWpHiSkDwhsFmNaGY3p4TLIOYB0
oaM5F2xrnsOEUlJ2n9oP1FDG260xVi9VJO2uQueYIlJ/moohxncsgm1qC+5l/5UT
KihUuZpmnEn8Yl57eB6uHFznPd7LCk1iXJto+Rs36+ovnsUSvnUqe/aBEDiqa3d2
LXQS5UBRjwrt+Y/uo6qgqacpmzDqhrNjDgnCajZTlBXDSJZveOVIHCdlUYSzbstB
SI6UE35o7Gdmq0/FLMdEQ5OFhnLfkEaxg/BrCHCp1QeROcN7hxL23DYxU5D89Uxn
foYJxP/6j58t+mGMEezX/rt9nedFZ1w/UOGlmKNWPNWYLgjytx4067rVhRKGnZt9
IimA26G1Ms3dmyhEoMUJvshzJRJiTbkDoJuzdhMyyeGYTmcABBRrsrgYqUROzDez
3iDeTs33INtdNYNKy7cfIZXfI8KcXM5Fx7eTxZDlBV/9cGzRwWg1OZ+3DE9h/UoF
XPmQeA6G8Iagx6PdpdPKuRbYtoMTVMxbHaDbV1vv+tKJJBsWcMe7ZNVpzRT3B/eZ
6+5Q4h1yPplT5++0bksVRoGwTl/k5XW3DTvkob21AiyOXs4csft23721Kux7OdIG
8eQGSjTu5bivxqyeFmVo5TAQhEyeLg+I3mKQDnqj/hcOHkjc1Gy7PD52v/vdoc2A
82NJZq6NhMncvJo5nL0r4wxB72HW2UbxUYPWyNep10nTD8ZuUzc/mfnZjIIgHjVK
9lGIuA+4W1yb4TQg098u8DOBybG4ZwQzcFq5z9tyGVTdsXY0MPSLizDqjMEy7Jvo
+gv/6df8jIpeuJGHMu9SY4ch0JVUFuOw0cRW3s6/NBNlnMV45tdxPbL3vWzELFbJ
3K15ehJLKE4MiNDstj7IPT+BgiteG1t6V5zKB6IEbtBpu/FI9TNFXXFRfJBxYzjt
smizJNl261gSYUaOow/NqO0PA2IVMBsBLr5JT26OidRzOD35a9wBxFkD/NETo6gC
pMMTyqh+Ejmw/3EuFRZLFqL8ZbHKQsWUzINCenABuOzo//kYRuPMFSqz9yoGdbt/
2+I2YQmK8zApgh03eIi/LYPCW8NfhM7Xu9N54lmZHeBpdLSw+Qj8EkTOS0/ikAkZ
zySBMIdBRmI102fyhipAfMPInl09N2+f59PKj6sUhKDdIa6D38X251f1pKqHYm6E
CqFUy3N1gVWC8ETp0926XboHd/JtOy4D9cRsfIhNVzOvL/3CMoW6HI7Sm57L8Spo
mA2tLmgKJgrCyqQEG6BulQIsXnZnp6+Ssru+7MCpr4q0FGLeZ57rNv5/SDi4oUr2
i2qmmotuhOOzfxL+o5TlzVzHIuMncuIjkkq1IA+BPb/9CrzDi2qpKbN/yrsXeY/a
GAm0ezfAf8ereOaQWEsvncfrlVG0YLRNSMT1q5e5UofX822gHg5+/GT8o2iAREHf
eQerPWvhQ6W2CZUKiPKUV6PiOivQ6YlorlJU/zA2mjoBwyweQJJeT+dMjyiQZpYu
CbM+l5WXufohh5QlR8gLez7NxvlzN1IBrE8HRSwo+LmxNEIWHEHRt+0VTBZrpGvQ
pENoNDdZpwczIJHcKPnWgnCr/8Y93jKBlGwZ1utZ0h7+vJikXVUV9VlFLhOkIq58
YHzQi2Kh1ml+1XGbhQpjbPvnRXc4eMByAWhjk9Q4ar3bKnXWjXaQ2YeWJDnYorCZ
tcMQ25wfI83Y0JhoC+XjNtzwfZxad/QSZBImXbszby+yAliDhNZ2J/BdV/PVn4m9
yF9V9HIURDsEV/UniftmvqCJr5vvQAp+AhSF2B9e9bDatj4EJde3dG+mBlJ3aI2k
ZWzsTwBCel0/uuj4K3Pux7a5ZChLGF676fZ7mrSTtobFMtkEusDPJ4roN+g/VXIW
ecZE9HPU2tlZSbb50czS76+YQncjoVPYAFdE0Nw4cdYRqWB6JihYBeOmsKndvgNU
hKyTmY8QVwYaNREN0GAGzoUmwrZ+APvL6MdSVFKZ+bS8yUyMKSIRMFSxhi3gLNfS
kh/GnZ6OPr+2sQf6GX67KLW30CxQU03TVvK0oG1OwaGWbvqxphQl4UiJRdMEbqXa
BnYplYa0+fqO0U3KGCUjal/AO1rwQzcAuFt8ITCua/+IKaIh8TsQN/SmwDNbO8hX
1mvLVpVcG9eLjLzKX1nb3+kbplQKPzOUnC1tDC9K/9EuaRzG8ymZVMnagpFpWpy3
GixLSdwCRz/fSYu1PtKN1bNkU+6cLzj+99/2mg6kwIWEygBAGf7ACXesisPqJlem
tdFjBwzIogmKwMxXXkQkCrW5SMwsNYy6I/1JE6zC+ovhfM2M9hkv/Zz5rCCZnFW1
Zr+0HBJcGwpNNaxHnpJ6A8oW+v0IvRwgSjufpcSbYqMrm53gwIvSRBHkeGFirTX5
ulrEzdln6yq6Msxn7uPuh1MMIc7wX6fHm7Jh7euSact/2Y9a2cznnVNp5Rl0suXt
Y8xXZexOE+nmSCZ5dAQ6VtlUzg5MoM3EpdVRzfdm92q1TbqzmkBSWyOtzHD1qaPA
wpzzkmpMo83O+BQBOVF3r3AbV6pD93wtEaFgcSBP+gZscqinlvD2VcPf0isegBS5
RV59I5qaCkphWwyjozdgzi/i86rheff/rFkRQRT5OtpTD6RpiVpxL6/AyvkR8VW8
Y20Gzs5lsYQwAlbR2LLgp76llxzx1vJ5KaS+SuuG6zNHIa3FEPCBV3Y0JZ5UGDj+
z6j1lM0hOiBxbYv93Z6QLvTnpiYBgRXP9SBBWe9GP9aDg8tCupVdqcs9y1kparUH
cHjcxok3AtHNFNy6cCr8D97i4zkO33i1MBSLsit39lqq7XaF0PuPDeuUU6Tln5aj
Y3FGfNNwA42S4nJPKzGdHmO82VsL3cAMg/KOFtcwwE+OLz1EawimYO34lfyjer3A
AujAt8Rb4Txd7yxi0RQOx06D5rHesnWHrV1pi5fKgO0EDn7UKtgj8mBj1sXBK6C6
/anF7zQaAq3VEfgK+vuVF9L1715XU77hID6yeJHOarQoRLMpWrzKplYdJZPzmtnj
Wh90tLUnB1QBK1CICKpH+e/XQgwmlyoYcZopnl0O/SOpGVVfBbUyBng0duUaUPIg
dW0+nnfIIs5EBfY3O+16o1ECZTr3Ls9qEBAE880g4alo6O+RpBFdGDLN4uWvK64H
jHIHyIXUwyObt4Sr1i99GnDyuYA9GKIoWjLBDvXkwJcXmHNNYXz1GargYiCQciI9
D+CZIRY42yaHnqMmBSeJACqp9mB08pZLbkMWVoNA3iELO3Q9aASzQPmVxr3zlbmK
aGPqevmxxc2R0bBoO3gWbou9RB3vfwW3CZnCTiEO5oh0EyPbuMAyA/0zBLTnHBuF
rb2WtWM9i9rL2ncSo580cg+SkcuB10bv1hZKBYxmyeRQdslfQiAdKra91AlvA0qw
wkV/QsGo+OnN2V6OXxZpJTzmQrAI8V3mzKhPQ5lENstzViHaDDjCyhNt0hsYBLaI
Ww+wC96/Qhql3B31usxGuADm29XMBmqknRJ1No/HMD9x2g/wH6B3EhLiX2B2SZ8C
HIY7T0ZUO8f+ALUO7zVoeidUbqhqUaMdrOd9dko4r0zM8KR7ans7tISrFgVW4sRb
gr/yBWQfNGoS+KevV3TTcuTkaayvIpdzvCHN/vCbFWWVJhm0cricf90Y3ECZpo3N
kFrCOggPiRHUB2zDTQKrqmBEcGTJ3RhpK6wFM8qJGmL7Pob0MUXSlmUbVclGAL/w
HKquFNYZoQq5eIn2hiM+1bZiv5efjdOPyRMzs3KeihRlPbAl2qC/9CEJ8j8ZBuhf
usilfJX6Pn0Abgc5ksYRgOqEN8uJ4T8k5re0tfi3JFAcLe4Tv9ZReP/sNgNst8ql
NIEX8eKacS9eCweWOd/1tQx6gTWK04xpsPpAq+fEhr/1ltprilTOcm2wGbOLAURU
X2U0lvwcYIkq8MQDNwtDuz7IfHUIqrZO9JD4bl2jsysEX2CqGYc6FiRc+xbbH2oQ
9opLB8Srv9wUT+W6ZOmux7bLROBSrha64J+4WH2RVmI3Jt7DDwNGKhvogjNVGTn1
nQBq+NemErnIm7iDFjIwfDvEL9NJwi8HjxXVIQxxhUjs1J8JeeKTUancpymUcOeW
j/ecqi5CE/nA1pcuUyp+0fF+2q4gDSr2ZaRyRhNHLJa4aHBTKqTnsSrPQuZD9+VT
yio42DAD4K55kRo5rwJKTWliPeI7hUlqPSPNDBaPbXvsmoBQljcRJsZaf+LSu3BU
8UgosLOAe2Voj4RL3/JnRQjlUQOBqwPoVLPlpc9MRyhHkpSpcveSDtcIUGPlNjF6
labDEwJYWUeCluhB9XEBJIgNFjW000BKMRKEhAnm1mGK88iJm/ijbWukqrme3mqe
j08OcKjHgC5crgw39bv6bTbJzyzKrEJFqyFZAJy0G2CPAYjXITW2drGveaEjYg+h
wLN9NqTGZa2Vi4juo9rIBiAVF6FsMNkHAmJ8LzPrudIbbAa2AMWRqBhty2DDAG0K
EUVnPDvy5SMSZ+QNSRxFtT1CEBe+FoI89HjmTbwyhy1w3veCr3bpot42l9qbj/cH
Qhm1e9auAqqNAKgkJt7Pp2djnYLwotEY0YPVRxVpN885AIn+vpQdTt2A8cl13q68
Mw7CoofdoozzdnorDApYXfTGM6ePPBbVjSqqTPyPsiaB+kSGs0XIAh5anJJAGN7F
acCWwl+ABoosAmGsz2Vvw1fvWvSBMvy92xk8Vv54FBUc2Xmra5Jo+5gJAi+fVb6t
maqnTEBuhC5ney4+8wiMg4za4WtEHcLsZWlEpt/BgKI+8ygHkig0AEA8HUuKNuJ8
KlD5Z76OOGqiN8v9P3v08FEIE+wfBz0wO3Gmxm9l6duOXe5LMm72d2qvdudJWMfn
WOZJ4Y2LqNaFxqfJN0iafzgwlkZeVsIL2psY/S2c/9GbBm5cbVsdHsIcvleI4JSL
q2OCyDYxotgz2c3MaxkZFldYcJSt6mNsJ5Wsi6DKkyvAxtXgnOOYNQ7zUIMbxzcj
LPKTLQGE3+7r+pDEyTeYQ0iLC3gNY5hPLNwpNeRe+PckXe3eHW7zAHEeFDw8i1Tf
Fr0vOQG5kY5thIWQjoZ9mHsCpk5EfrZb/yjuN3+uvpwyCwPLQ6rAXNefZCKSIjkE
I2PmGkcSVTEQhYH9JFRh2PoDxO2WIkRaiZ/AoJjPN/B/0wD/QooaqF2HmjgJMqhE
tte4tIbD/idIrPP41qwy2DjGf2+YbMnPlbyFWDXFzA5iFHWvsM6gXN1LmyHi9IS9
dIgmRY7IDLxOiT6Ew+FGNjHIJ0P7ROSNCLn6UyxmTmfaUHE3ogAlU9WY2HupzRgj
Ldfh8L0XTfg0tf6vVUbYWYV4aw73KJDEhhGH3oqE4LtZySOOvUTtQmYd5Zux0Abg
Nt6INfcIVhJ01bfLyYkHmtS7+tBvKFzS0Kczvbte3FGgYUxn0tmQZ/r6V+jKXi2N
HsK20Hu7GEK72r2WRD+27ynNMqA1ZVqmI++UTnhHVpP4W/xtzLiYDn53s0FcDOKV
lw4zPSCJjTGsG7lgx0SiekrjkLeZbE5yoCR2SG6uV9LD5xR4TStrr0Wrno7knTfG
UdnEtnDFYoyjApT0atuaLgOAG75fSIf+IR7G0hDEwLt+Bk83EFLzgRw4+NU+5TFM
5BHFX342dOWyPFJ06oTzlB5DZ2/CcYzVjyOI1j/qbcuLNzg+r1fnWY24Vw4HrbzT
nnMadDZLN60mjEH39BLnXCrjwnvRrjshDqrDgPKi2rKrvqc09iFYUpIKH7Ed3fyG
ATGMLl+6m8WFIHUiWepbiBekiUbahFl7fSNpsojIN/a/g1D1pvEdwn7eFgXvwEru
Jz4SWuprpGwF7YmuvRsLfWtkzgZgYGxUJJAi8sB8X3YqQkUSOHM7FtdDLCCdEAg6
3+aLN7P0/fzjmhv6vQ00LQs+If4uo5Ae5m7gePFW9X4VOBYhsus/PP3QEDHcb3JE
bQ0UsqccfQL3qWB6RKWtBLw2QRpVZjhZ1OEAJ+8UcNJ3FIaeVXsEHLJcfIsEwJzs
He252dQEzjtvN/ZmsWHPWWfRl19W0oLVAdU1TQ1qYFgEOclz0auMaR5zV9Lg7X8k
geOAEX091bjB6sndhxrYds3wYHNh9a6sGgec0V0zU71+HHm0zluSnZ5v8hP7teXD
w1VSowX5NIdw3H0Bpx+C8s+qL70INIXu6eker29GatZTYrJ00loX28UVGoXVMRZ6
H0JfAO3NEqsvFcTWN1zD4LzfLAmP7lIVI0M1XKKSgn5GEG/nI2QSCX96p7Z5O/og
qKpHiyTS+5eiG3e7oXaGXy3I9dHvQyVdzxybsGvguB+3yZs4Rg/8Jl3YH2oL9A6A
meJWvOke+1/vL8q6/AETC2FWtxZDCajSqH+fZfyCMqPOqE8I2AtJPltuyHq4+LrQ
EVMvzzu0Or+TGPKMmapReMHrYUapjhcWeDK6mHK3kjdqfVX3KQmdzNIQ9+h44iIq
kPPYFwrmLG9S4wpVnHq+gd3aZOgZusmqmm5I6Ci0YhZEaVd60OK8JKzcCQDey5d6
mQIHEjeoGyjOSUCzfJYImDFWZj6Q8QsGr/Vhsd4VmsG6MXh6ZNcSOI29dDyGxf4Z
rM1wjpZi5tTvZ0I27cjscwmk0Sms5Fyut/LatxdYmp5RcjH+zQK8QaAUgRnb0jZP
+ljywZaoeI+EtlYXl3EBQQhgGdOzvVop0MwAleyBLI0rie5C1PqEMrkk24AbjEsm
uKObGzb1KNx1fHtOO63QR6g35GKZCYMKqAXenLH/YM4rY/0o2jhCtlF0JivDpvhe
SXVcs+cM1VkbDv9k1dG3uTmoed/escD0Sli72PkvPH/RB4Lp46M79xLSl/q21VIy
5qSwGehWda5xLehvZms71+DULKzUj7imOYVN3r3jJV50Mo5YMZMxTt31IKw7UmbM
+UseQxb5+duq5IMvSZlF0Q9Qd+PLcdYDLCwGLCJjoSSYlyRpMBZOEw4M7sN2Is80
zI2ROsoDpC2gwnL4by3e6wDJvuNemjGpkazGRrllP4Zp2kSGBFnNgPd6qLCToUj8
GC2LadiOy/VVHj4hfqqFIDP6LTZ1dLwBq1jNva3EJ6qYGOEnfN/f9r71R53g9jG4
4lmYZvihAbxhCLtQXVQONvn5H9Z/Rekx1fzJRUk527/oDKY7pRtNKAACP0OtmWey
dAM1PP73NFysV6Kz+aCqcCZiACY/lDmtIFDOUYPhgkR+Dd/j3pqXtK/zS7YtSeLI
iiRFKxvB6970aic/lsy7G5oSFs67HBKqtfAX+YcfeW9m7XlTm3SZoHoNoJcjISW1
HjSUSqRjeJ09Zv++VVYuOqe7RXPZms9hKNrlxkwCry2oCMv91vR9kynam/N+j78p
OV2cl6mHgQUB0t+vjEuj06A0VnDFN/TWBogPDPX0C0jXTdBupZrXhC19fy9viu/8
sKCHTlpjZ/DDvAZYWTEnqQhtcxgN+qd6R+/rMh+T0Pj3l9cFGpHh7xV793SOfx+X
dpvd3tP5+8sk3gTM1pI4inJkYIW0o6L8EhajOrv57JWOmDvA8QYEg5heOTW48fbU
WEGYAqa6j1PGdNNt57ngdqJL5Pb7TGcSmupuBPvjYsOkyttB6xx0DUhr9EF24zQ6
GvR9kCXbg6y+UpRuq3EYTFxvTfzUcbm6ZYLiypjk3rgvc7KKNOwPRXLDhW+RHb2S
qmxoHFVGMQ/YiOPRM3mmFdTkTwB+K9o7q2Iy+/KSBpAH7G/aD9Dw9pBsj5iDJ/2b
LGgM9OKnpbHf61zmAgweHE5jIlLPX372dB6wQ7ghB3/YqmEGU1mP+IHkhLZo9tQI
gFtfvFFvG8Zx8JlAFuJ7bJwqxZasli9+UXwE7REJ+5PAXnyHLj56jx8JFDtn710w
M6QG2xfALFapC0clVR3BhE3DhFQIQDYwhtWMNFNKBGGYA9fj98UkyBsFvesfjtAK
8HY6WY4Q0SzbuvrkQKSWuDilvv8uOuwjCPNBRy27wTa3N1R61wCkEheaIh/bXuMN
sjQCBaByRtgUOiV/waUUkw==
`protect END_PROTECTED
