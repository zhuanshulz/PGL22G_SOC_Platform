`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z3YEwtffgsy5v9hxcCRpvpnKU0Qk1J6Ar1KjXgG76cCUBfEd+LfijKjnYZd/UFXG
HYDjzuMnB9aKDnIKiqlv56DZ+JvGo1KhT9spex0vsqjQG46/MumqQarX9ur2ceKO
chEt47yMIwY6XKVoQYDnghDbL5QpHCkl7rYiUtWE9pBlCLyjAoSuH3XPoU87v8XT
BAC9eHe6v47JCHcIYbZFzZQSjLcKyQaCkNEzKrsrdyPcmG1Ez2FOglg1l8uhwY3C
ZNdCMvxeXjBngYv6x2LOCvuqC9jNsl9PnWi5O//YHXq24e0bRqVaB/8eZZaIDNCW
GaUAlefTBDknG/iTWi9KLDLCVDYigKA8QLtJRWwy0hpJSeDg02HbWaFwmqnd3TH8
J4KyxiU3T5Lyo1dWa45MjgCF0PuxyfpdC5kzOrFflKYBcqXzCllkfdCKr8WXsUTS
vaxNiWIs/62OX9t+qvyY4X50P9feWUUDP2/jiWPvZrvUVkmlybLyJj7X99e+/sXo
JrWtokqJFCKTa9YDVcaFgxVpyZStYGhoYeQAbxWmbuaGKSDchOG3veis4YEeXOBP
KngZJsB2gZ6RTRbWu3RfU5OyVQ7dkJTqpuxUfuCczyOR2OYak9K7oBiY3VB0+aWb
38hN2r2JYvi5cL3sA35Anrmn2sIMu8c6Gp4WUBfTjsQnQ3pUOXsm8rUotcowN+fz
oGNuz9RvsZ7o98Fi7v9jT3RAYXi4ubd3+RnvqFg064v95O7TaZhVOPyuxI32NcoU
CYHRzl3oYYaC588SohH0RC95rFacd8CUjkYnvVhk4jtIJYBEy4ERt5bd4pDcs7Eo
doo8+gvCqgwh9jxOdYS6lH8gtrMvZHL92pZ6kqGp7PkVoqgWlvUfc8hPEGe+oF4I
VqreqFrhjutSN3syJVHZR5pqwKCg1HrKdsAo1YpS9d11Z4e08hXZu/m0lPqlIzQE
KqUlzj8YXE9Fzmm+BOn1tntimy9KmFfjusGlTtUXgucVSZICyKQc7hCGyMR8Ljjd
BwYIss7GbcYv8TMMy3nEaafEg7P2nUwYoi6iPujiTm2qVWOUmogkEEntHfVInE/c
/2zfgpPuTyYOgTNStGJQA3hKRdniXh4OH/RHoziwVcyKzxBdBfMd69s1wEh9p3vp
p4PJ0IvTDuHFnXJBHMB00Qb/N/YWUoSWpvrJzubOLuKj/wvVDlpQewDc0DI7upX3
yqWDv5d1rT4nZreDT2aMEZ3IzC29WRPBjsw3FLAvpLJxRKs6VB8z9LYM984PAgwe
R4QvQR0CWk8igZRfC7tt4oW7hRijMAA8wDXxI8DbhXunPqWuaH/sbkPAxVjHkNT3
n3ylez/177bNK3EXzdXNsZbxSL6x8+PCT5JQe8yYYa88N80txOdofzNomiTFL3iT
Thb3JHatEi23b7YvHYLoOp7WFR/ZGxCybvIVw2l9D/dQ7qAVRoY6ABFcZF1hZZhx
vye2C+fo0bfXYx9bneI6LYWEBr1AXxnfj6pAPSHnFqGHDP/HfjYQoeKeGSJssHHZ
FPTWe4M2x/Ks1Biwi56Zr4oKfuSONjFPFsxDQIT5IH/LtAUHWmlGSjOP8A0O7aR4
pQos8VGYtzFSsFuqamyr796UBMVWMg+ejMQzVC3L4K2YcZYRlxGmlYT5nUatBkKu
`protect END_PROTECTED
