`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R34fbxLZn8vifs7jrJrG8tCPE+SNIMSbnKxxHcqU30VaUUsC+FrsocjuJ7cVPWUj
UWhb41uqki3yRkeE8Uz7tkgCj/IFaccZST7BtuE+/hJjz/aIN+YffGiGorEftoGc
Dgn9udX8WwfEFosL6Gkskuw0+uxSAD7dZEqyl9yzR1lNXQIdYCOhUzlmZ8GGnOKK
ShGWsS+ZYB6f8a8nI0gJEKzqK4UwCtwqY1hjxj/UrGw3PTq5po+wFzliMA9uLkjj
pHvPejjII1KhEhPcs1tMCTiB8CBZ+DdUmdY0tcs1pwWjxPbbq661SauydMjTk2l4
duaaCKN4k6jH/ulP0wYaipZ25D3pmU4w045WU5eC1zKVAJ5Ob2YmjevmvPIigVI3
sE2da1WfMofR36i8bXBOFg==
`protect END_PROTECTED
