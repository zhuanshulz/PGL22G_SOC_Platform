`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DOE+9EKMZz3b/DaeJtADQ8PCGq8gaxlAZiiCK4o+2+Jv/ZezLHOg49eUvPPhC4jL
2k65Vz3Yjzi4j+8F8Gd3yTm6zoBktyy9gs8LFjg0kdoIWn3cA3CNwEUTHUlastEw
irEs0wt7LV+XO5h3FWLdPJOem4Su/uEPTmzMqiXgkk0JZWYGerZQ/q0+vMJDXdRw
3blfBwEgVERHQK3DF+OhqW6NSyymQ73xx2CA+1OxEwCyJ2bKvzy/2EjeBBiY8sD3
O+Snmqk/8SMXbCiytrUboM+sm9m5JCFm0xWsAt1f7mUiFoLPQ3Onq2RiGPE8xFmU
QWM14UN9HtdbmrDZn0oUo6qcgJIxmz7MG/tCkA9/WXblogQuz6HJvsULkUq15y9l
Pr2ZSCRpAMUj4f68TD4eM3Wk6WpjaXFLLB9wRzc1hEsvn3HkQZxj4azyHKSfdecV
x/yVb6QotwnbOX4k/vD6uuXhf5PBVTG/pKRyYns9GnenzlqUg03WBgO1m483kkW+
GMa19hQ7FYZfGEYA3EmFTt8Wj2ACui7U5HzFfySZebcWN7FND6+xB0TwuvcB0bAC
MDdksxBRK10GwJupP0hRy6AeVNVvkqOGnclCto4TRY81koyiUArxM8d+y21mevyq
cfnKV/8vWIBx6jw21fgMi6qZztIDxzzfWxQYNQSMjBBD1Cm28XY8295LqmTspij4
ZZGvWeNrvWUMaqR8LBg9rjknKLdcRA0paY42LL7RjXG3ATyyGVV0+5tWLFecMOF/
Fe0hXxEs9E510/al6PwRIzeEibDhbmNzBnkt0tSpfc3BNay4VzFl8ePvyXn7RLy4
EoSJkxg16C2tXGbGVipozuursplJYyx0LT1I2RwJmwdFtGHrq9QFTZ1Ac+mpvHX+
ls71v5gy/5r0YV/oXJwfARCUezAF0hv/ds0DXMd4FlO6o1ja8FNBrsfilKpExSUE
v0EKF4Da68zmmGr/FUvKc5dXg/xqddFtgS3LrWQmeCrALQxvtXR/kqJggyG0zYwq
epI+rVAdLON6cCVjKL1avTPIuAw77GLOx3vUNwfLewo5oLp9N2XjUWgIXjlNFoXy
EOtO/tehRMoO2p0MK0X3ilZaX4hcEGwBq5zCE/tggGsf7+ZuQcbdQjIawj5Tahto
u/pUHgcijQMlnLmILr8ahXnhikyfDCHAI4BleVaZ2vyHWwzQd1R8hPlyu2rPSJet
N4Fw97VYaOuVJpA900vB5bvKrLQx4IZBJ7kQgKTBkkRDl1CwOaS8t8S94mMh2EFV
GIRpOgs4mG5k/ZuesNF0llg2fRf1ucnw6AgF4l+D2t1KWCzXMYA5/6Y5cyVhcdhc
5jwkTYpvi99wvnMDOpHAomCn0BNdY2EtySnV2tD20sSsxRjW17ozXvmHJ4xVzIHz
EV1Uroo4hF0vR09x9HJr8avN8DaNI6xJlAlNP34QyJwpcAkwsi7L0yr+tEljh+8w
DTJh/9wrxt6a9+lBLA9Cwj0z6B2OONsVBJQuOPGXdndsv017FO3q0cdKSAz+kRn7
jBAJ1b90ge574HQ5mL8rIBdZ9ihe6ZYsaTdCzJU0pjjRB32fI6ka78HUOHa5UhZz
u9kEk8S0kbWzdnzHW5DgcIoa0iNrdrcvrLyWmAWEt4OjqsluiKeMcNk5+UR8QCgk
zUAgJD6ZwAlUEZ6hvVM37Z2Ej3/FXCQ/aQjuAKWGLjpglx9a/wQ7hGghd2oq3sD9
+poioB0K07jR4cNLjfHSI5rGWJ2v3Xo8DT9U9FOg1McsKTDmUwBt4KQ+QoNLYzns
5lm/O9boV61yPpg5L1M/awAt9eVaeSYiYJ5TR8Z36YoXyFqLf245Uyr6GyY4kXYt
laoTP5CWGOKDCDnR4xJv3BSKtLDoEbI+SosslShKvXjbphHO9OnS3lkjGIfAA0fz
SLb9vn0qy1r/wOXyIxDR49tZQO8H9QvZU0UPVQgHwatLnCJO26NQ9qUcU5SP6ozl
`protect END_PROTECTED
