`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
myOawRM4v7HhJWg3IcJI8k/3pfC2dxcxPEqB+YD8HNvgfPXBxwDxsM479Gs1z37A
qR542cPey8q1G8m5vWCVOzKXjJNNITzAE+aO66dIw642Qkqm+0XW5aUD26ov10DD
F/5gaHtbAtv4shgzCBv4h5JVwV6sQjoNhuQWLy/YlvTv/pTD5qJjKSip3EeQoCgJ
rzTRimsFj8SUjod3qn6gpNsAQm1DPZ8fonWWR+Lo13GGENNhirwZu6qCMsLT3Uv+
NdIzcOLQS0lfn+m1/TYEoij21iohJXINKlu0TM7RlcxDqmMtgrNPdK6Z7iugvRXj
Ie84qikpfODP7+vjX6DIskCR3T5avT3QJODzrKYwSVqx9tjYMulHKWOdyCaYDb5t
rW69dzfmp7sR9RGiLib/tpil1iHemiHwYPNjwjaHTzfDJdu+Lp5WgTxOWvc6hKJq
cXK58bPPvESHJw9w3ny7XHSoolPb94j8PjJB3OW6UlFl0/Q4sSy7wkL4R9iSQdG5
8gnBlIk34XPZbRHBVRMRaI9Z3gchwwXn2kFYi9p0vjm4uDg3Uv8GtI4nrdbWte6R
zF47qvcw/UQJe/r/oUbLO+AUsSflaLqJBM/3iqSQl7jVfvjbFOi5iY1ERS677ols
eBkPv3iqVbwsrbXvAmkekam73xMrPP++ChaRxhmlQAwYE/Aeip8Sr9jlB4T0RBM/
KIr1lDKv0GEl2nvfJRXMWOetsE15wSGqGIEbjrGvDqEWUWvogyujT5Z3dcIgdWR/
j+t35So7GV5WV63PS/2R3EnmIblbDEptXKeuhTc5dnggntGC9L0WQ20OTEEIHiQV
/eQq31HciTG/8fVQ4PtbWRrLnUGldREcnRCrNifRggjkYS9IwzGHB/aX3imOOd9m
N+w2I2DTSDYjgUHHpYcOmSMhV4mjJn5MEgJjvLjDHHdENtRT43IHY8SuoGPrQqWu
irMbpe5A60caqx3LzbuGOEYh8Pl/BDNqToEq/9MwRvDvRkEkdDfEtTqY6FM1Ng8E
fbC/mXV+DXF4Fg8qVdY3jFL5Xcxkdgu/2+W6CbiDbdAys2D+Ag/UMy/grPOS8Lby
HQ1aR9esCCCBYoVhLTfueYaRNvRxwFx+61wUM6WftA9/NIJT88et9Bqc08FFEHz2
gFC+B6LyKwzPsisuzM5lNlbNy0ytKGScJCBrNFOXjRnAM3isS79cvYhxuGl/wxo8
bJA2AZsdIpCmfz1Z7QMs8gfqjNOKyVEN/yCQMU1tCvKxLEoyuSZcuYjhVUi6TeBw
yAiEDOFJWJEKFXCRww810EWoSihvfnUYubnpx9nvMtS4OvVAv0/sCLkKF6DJed+T
OsV37/TCmxzFi174g62crFMXsEBniHZxzqkFtYFuug2PZW2nRT21+DDwrJK2mTkS
9qaugTrsHAhOruWIZrqnD/XUrVaG7f53HF6uJ6MtuyDoytbpXt10ezl/xoRHVUjR
CKspvjA4KE3gTXQJvNlSgbGdxxTFAGoRDQHUN/tgJjhe166320WHhpCA7QBG705W
ijw9RrXQQPMiiE+Eb3r9LtADT2cs9JPtMwYNxF5P5TPpHXqHb7jeTrP+c2jEr3y4
xO8t9CaJJbFT5J9rLgmdRSbFhk8LxSgSGSOoujE6hQv8oXdyUPOPASG7tSsTIsCk
pOuj4V4VFAoiMImUoZg8Wt3SPOjUIAKwh8OrsYj4zI37sLSn1YVk9JsHw9rqH4os
hFLfuqlAmm7t3zP5SaRMUVkkQ9USB5hwT2z3YWY3MgQB7A3oLdPusVRfTGrSJ7yi
uqUH6Vh9poehELgSAhOOnvZoQ77GAOU37lFiU4PAozD0e3mwHobKDm5GMxurFcs/
jgH7bzUSRz49anar/Ag58GZm/NsNx9d10RdFeDz5ntmJzfyxN5WYkwqkntIiEDVp
gKGnOQ9CqrQAlksyS+cIjZFo4Umdydd75mTM+qdM38kAl+kqbuYr5rJmgVtxUDFc
UQZBXeRXjDGcgGV3Pu/RPfITbFAEgeAzDEdfIbeHjV7hiB0RfdFb2OzsPxC4lHEo
LWgfpoUfbp1vuHHjdDQp5gwkjXjO8CEQSXTSFQebpfYgwlKN5sDI8X/yjmb/nmRI
NfCPR56+NHj6YZpiUW93GwFZfxJ92iS3boGRInDIg0+WnL4J+Hu6iY9/hjuw/aPT
Y8LvdoKye87g3eCGMHpaFwZXFx7veXSLl854l1hUAn6PJFnKaz1VpP0vuT8Ajq5h
iswDf6baE36/jixsA/nPmypujQ0x36AuUBMF+uh88r/5MLoe3mVAc6bF52fUsHIK
r1wCCfCFpAEHiBFBAyOj5MzJEo6ezvTEDUw0c7u7MojJ9oCf/CROfcubnIlTuT73
Gbfz6Xs5TtTT1CaX5PrDRxGkoUt79u9ifjOcwE2UoP2DVsocKgltj00qpE/9XQsa
FH4e5HJ/JUngK0nuOhqv/M0wKwWFaJqvPuWn/p/tOlQF3g1j4P3pf+pOe58t7cxa
Xigxrtr0rN5N8TdGzzOXrfhTLJe2K+e4uAGDV6EDjY4nliWCX4MRlNNFZOktiBCp
GUf02cZaoFUNK8T0yYXYm2hEtlSTlAdlSk1J7b3tTiCgxqS9v8gHFRjxHZ+DqaMV
Kw5uUt2VpU9y7TsZ5I7uS+29hpVNPKvAs4/FlGgHLVMT+xsjW3ZcPOrL3Nwj4Ohs
Q3KxtzG3bLsm3J/Kf9HbPprPU/GGf1Qp3pApul3jK5VqPmZYu2seXvN2kVafAIVs
3kOL/CdHC9w15mhQdLautRheD92N266v58D3mZGia1NSC3AgbDXgA7ylSKEa2yqr
7YhVBjdfw1FfhGE2aLX/YNJ62Ktm/y1lx6hh4+s2t2NYHVEuBSoXn6LnhpsV5Nw8
KWZ9hIWIWUzJzxbFO5g5+sDUBb/JeD56opmoqjVJiZzAeh/G/+oondWm55CAoU1+
fT42fFjzpPkVFf7Q0cg5/D6fKDSn7t/T9MR2NzXKo3m+7nbRgMuV0vN1xISh1Ffq
+gMrF8VqglQG7/tziw5bNBq8W7f8tPXfVuRE5OezZou6tWIdLsG5FVxfQVGQYJRt
tAsWpmUuPHvstQ5HKJS+JF0nFV4bVX0IY2QUZiv3mygKxFXq3rCQWu40+42VmSEx
B71mLH6JtGdKmVfhfNAJdBTs8zZjgluZPHmnA82/RcsoYJnWKFefY5fbBmXb6se9
Lmjvmubtzg5xNwi10PyXVpXf3inmBvfZB3+kFdvSgaU30hMiinnBNdfuIUaeOybX
IVLdJ1p9+KLuXGWukJNekRobX5hgYoAVgWqUuK3ltkruPbACaUJBGAhcF2AHRNNa
/ZXfA+X0zZ/QnDcUFh2IWGELmaAFSLeFOkSBWn/0Vf4aGBHNJnV5T5m/xvF5ktlf
Rqa6z/o22T2PbzE6GZ8dmhGGtYG9+jY2/Mz9yDLGvfSVcqMkB2nlXy3dGQnuuIod
4dxpuAEL/TmeaBFh6+XwAByVA2tkbLy6Wp+iRE80FuaPsaT5/aODhUBkrv3n+UzR
ASc/mMbtdt6dsxhuUmovtv7qfOUR1ienzA0uTOIgRYA+4FmYD8LRKNDXgWFKIqzW
9wAdPhFaCepNFYv6iFcNNfnSCukmdL1QIN0uP2M1yIrt4ewruBL7Fp/Q+T1zpJ+B
nNpI2OGknkp+3QfWYVOAeUyJwxEIY7vz/qYxqCgHNvV2e2isV2/eqJ+G6f3N5wat
nMTrMq1OFofxLOn3v4L2ffGzm6GuVar8iS0BwEBiV41mdI4MixbTx7OKjasTKhtK
zgN/gABxF37tBm4+dQSjRXN0+sKOkaal4AXmqjz30p15MWxbo4foBgn2vCWvUI14
QErGo3kKe1qFkU4YPcNN+4r1FqdXIcIwCNPlvl5OCq7l8Ox+qbU8zM8XO6TBE28o
rOGLIZHOCl0MqQ53ZUsAhA1yD1TosIzMrFjQhviRVzWE55DmLQuwf0aNN/EVIyGi
YlCY95HFLN6ncJWuQrF3KeupLNRgQ4oCnhoWkg1YHsRrtUXS/kU0dM5HlcS8nkcA
8ekx8UFlE2ZXFbZHklXxzxa1JT82LNfGCnyMosVfD0S+58u2sXLapS+akQ+lnTkO
ULK+F73bN6q7V6v4IEQxt4QDODBjDqY31qq0S5m9oJ3A6M1ETF9e/CWNO657jR98
dhqgCfpR3LtYb6W5+kChGCwl+7H/FP7A+i0Kq9v14KR57azBPuESy9/MlZFSBKmt
IjCKa3nkU6eRypaB9naVtXHcwrX3uPoj0Ne2zSSgMe+d7aO7UWOl1fHfm8DAKiCB
CPDJiu9USauitp76Ln6wkBOJAkAe9EPVOeYm2nJcZmUsAxvh/nh9TCtN3RXmKwQ5
YTbo6gQZcoeAYVte6BNdA7nYOJIRLAehS7PuChHt+3QYeZy7y5wYN1HYRM9+dAn/
w37q+jnSE6/XJXfM9lBDvlbleFUUlhnMUlhRb+CVAPdV5PcTbFkV758S0hrZsKdS
cWTsY9qy7DMPvipmGTCRIZ1JNcKtu/4sRvlDPQEaBpwtGr2IA+w3DiH6fcqPHz0u
JeVM6fbYvdUHPnPRas0TESLNnXvNkn5KfkfUJtSUH8z5//LgGcVgMfyXMu4gWjyw
LDHk+sUjyAN8bh0z22iDdas+iM3QAQy+fE210OCabonGIZS5oDuWCmkxxEf/4NxP
NVnJQaKI59xA95Bi0YwacgO5pkMs3vP4xUrGn52AIM6WIDvoFTGxbSQmDNWEVb6V
4PO3d7Z2LM2w3uyVu/TaqcYtFGDxFuvEyMMRXf/TaWURf8goFDDCHodYRahQEfb+
c1u4IEgU45wR64V/7l3PvPVfqJHXQpZXnA/ASEWVRU5+RGbUKDrD1dn5ZhAw/iD9
0n8PfgCWck7lE3NuAQlVEQz9Oe0bxaAbacRLVcnJdzl3UWcAfD9itn2nHa9FBaHk
1ccOpdD2hpsEc8XTfQsieKUhI2TdMEyWXuZSu3UzVvhCscu9UxorMeWTizl7rDkN
sncobr6qWpQKZq5NHFf7nDnYZeRVLcuEpi/I6hHu25WzrOGfzW7zULOQmSFpxeU5
oQMEVQzKgNwzDUfuZkSf7dDlTzrYVyOFzTyHoAxVas9rq5+de7WFkikIrUm2lWGO
4G6aWTj/kfK7mfwHCbHdBm75F1WzcnAYVSc/O//TwlKvQ/cQt8JKLVGFXMnOdsRL
F1kXstMbXqWwIaZBlKJxL45OfHr+CvfXVwGAHTVlMkYS4h2R9MM8/1KvARHXuPdb
S0+CS/Ul3T+Z//PfZcflbDGHFJvG8i+YClGiBV2eRxGH8lXHSFrri0oJVkaTAKjG
ZHMElFgMAuFGxkHqUvH1HP86aBTKfEPL+xTjojqElJSma9JMwFtrJwkH1HuEa+s3
lskhjEusQVDSK85m2H+JgOU7rl0JHMtMPye184FYjupbDtefAqlv6e0v9/DVomX6
voQzpm6chCZMkzhYIGy/R9KvZNisE+yN+urUZpLz4VoheauB+sNiEATNV9s5vdBk
Pi5towanPmpHh3aJ5PEeLGcDDZgjteFmJ9nBbU+f+Fu36U2SrNiXMyKWRscAFqYD
/hYjb6AdLij5e/YQHDCilBHRpPNZqiZXnjhvCIDC5cdnLbnOqZIPc03vQRgwNuUu
iX94kJbOydQ5obzl3yHd10l6r2vWgvF9J4n0gR2TqcSDdy7Z2u0bdYzPY4hdpLDo
dy5jECm+/MAuXCCIdIkpJDEK0jMnIlBMrk/qhjd3meMBW515Z+vDAQ4BbsTgCM/G
+6kOnRFheOnkfxeKSILUruCqCXwz6IEWvsCrgV7LjfZ+Zf6aw3HKpijRlpxZHDWb
KpsesYwJyxRWrfe+nZFKj3IARTlRw8Xm8BxJH43ksMVWyQiS6iuYrp3Axg1d+CjZ
Hbr11RHmR4fQ1I6pqZQFsjdbKzkyKFFqQ8qB5c0X8b1lNVtkrO+8+pcXdNFn9gVT
5W8pZ5+Ey7VWgki7qj71gZjO27yOOOCJ1dlPqDvmHZOuY0JBpVsgIg58NcfK5L7B
z4HOe+TX1TUUAZ1rcrJVs/vKjYeMBbll5dt/RvXrgwRKjdk7Nq0oi5banXt1qd7f
Lf5ztJDmq+iZ+nulZnLb2/ZU+I2+/3AzX4Y/5cLv5C1LLxDRHKHUhj8mmGyPkv2r
`protect END_PROTECTED
