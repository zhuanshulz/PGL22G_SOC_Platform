`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vEeo+1VdbnmN+UO1O7uF8HvRlkyfN5o4E9BTJRUovai7d3ti0hbQYI1olKcrpUvF
PisfpYpu3861ug2VVbqq9kws7peFQ62Ku512k2P5JiuUdhotkIgd6rOBQhpBz9mW
r1xIRaUOakKi9c7uB1TbPkTmHQdk8A/el4CMvZ2VJFrZoLcrvQcqMW6xC7WAOXdY
C8NFtPDcXryD6ad0L7wTGX/3qNB2awBbkj2FCqxA0DC9v+mntDN1iiGEGmwNh+hJ
fUe9DGjtWxpgMg98qK0WpioZgyh1pOlsyTYsxaqFZaMguMRIzR+7NbEci+iGATAY
8YMA+t6z9HpftictBb2yoCu2urLMv73fLGs5ScQVn+f6QOh+6FPIQiqP/FsYu79u
M1EonvH0eMBHSHRn9VTtfVe1WgaV+gcErfPm4M8XIqbefQBnx6H1KsAFGUst5feT
aqsVXO2OI+I1RhwGKPWefH+ED5loVekG4ezVvpxOMwYfYSHHkUne5Yl23rvB/qiw
jNvJK/8wcf2UVme7Z528/iM5cMVr/JGUMHtFpVu+ma+o9uHw1JEOPJiS8owJQBT3
U/2dq3pecY6DwseZyPSVOyZFK9i1GjQUgWzB1AHzSX7zZIMvGcP9+hR4Cbykn8vO
XJYZ7LeCjuP8E8ShBL6/RA==
`protect END_PROTECTED
