`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8I4kGLAY0jVo5dA5pCxh3EhUT3Iw9/fT67tz/PRxSaO7nGlnW+/VSSSNCKwgNMro
NHhZo5YX5pBSmJ0rqX7St/x8o8KZ3GItzZOQId8FqhbEAZ/thkXzcutTDuU3XfKf
zHugpVhUtGbDcwFk+YDSf0kBa3DfkcjZY8wnALubB7ez1kRf1rYCBgMwoRgMKI4j
KX9RbDQLN2o6dSn+pWijWTx1Fi3qE7rN/FQ/qQl5fVDLaVUEFBf5fDBSihjysWti
o5H7EyqfuE+MR8R/FQCoI4ySg153ai0pSzmmNr46eLAi089i1MC8t8prb93FuWVQ
mFkTK0bvZ/C2xLX8VjinZyl017jEkxeGcV9ZArLh/Ycb86kX/oB698LCIZEFmO5m
OQtOpy5VK00+45CxoGdmcFzDwiXEEF+omyHUCJAj85O0rGY39sdfCFUWTUdE9L0P
qkEDgc7eCg6SQkWmBqh9BoaVa69aRwi3nwX/xLeUcRaaNoLdwwtHbC4u3H2VM6L5
ugLdLkj5Yk4AtthTd5dQoMtRLe/1IOGCh3niiwSNWczB5ZRvbeoO/arAM8V3WllY
hx1SbGNbmbUd4S6KMCgmlJpZCFcI6YRNuKnsIsZXpxXnCtEfgv22UXPgy10O1Tkq
Rm3nAWctS3aMnKliXSFCsytXDJlwEAZflTjzY9Q4v8jUmHUgFAEiFvGv5wHZtXM9
+07GKgvDUdexK5gHPF+jqfE8XxUs3YQU4aqVScFHKp0cjH8M7yorJdUrXCqQ6mfo
z4TJs81B17kWnj1dVplmAskVfTlxuFIdVdTcGsxvH3lhNOMCJCUZzKqOZwXSR9lf
m7dcZotnGIUNIneg5qz3la3DCoEbBML1nll237zDSAmjpkdaotyqnNH1KG+jIqmT
LQNqbdfgrwA+gEYu6KYrfAO831CbMTV8NcSyPh1NjTPDl+uvcX9Dfr5IOSe20obF
kBUGZdeh2VhjCMgbPQnuXcQsBQQg1g+Z4yw1ccFNVXXn3xrmi+uAFNGHo8Dc1Lkb
NDvjghkxLbbJ0ZeWtaAG19ZQLTOmuQinS8skev0rdDg6B5/4CbwcRfWsYmP0zU+w
gdFxMysquaYBjqrdmge3Jw5Tg6sr7tk73Y3kqlFIMOEUVnnAeSEkkcNp4u7v8J+v
aqD67hbRfvZouoDiHVk5wo4y2vlWiynQEvBUxyyYQsoPpcp3k8Y4X4WP9ucRGwAz
HLvCf572e9uZOaeMFp+j39gu4z0XdWcOvv826j7ju77meHQstLyOhw9Jy+qKx/G2
zhmzN6iI7ipK5eYVs+thDpyys/lYkZu7URfmu+ipWSVVHfyOElovLxMs5Dj2Gxfa
B5Y9XsKFkSRR14xwlITqjXamYB9a4XeJ48Oa6sunYJa53/F72IgugxGjfOgfbpn5
ZkLD9SM4jUU9GUdw8cy72mvjXyQ4IZZlV2rQDb6KAGA36badJF3PnbOhyZ0k0ibO
/Y6Glj/Wo0sjhScDlBa4TVgNKb4faT9kkF6ievDzy5nw90Ygk6Tj0sHNTRll+SL3
6W9x8UHuf/NrAASusnLwbI1GamqEO+7KnO/77ShtFiXxq3/Mg187ymPfc5HV1Oxv
YNWRMvSvvQND/WiGejJ69fO30syAprhHh5AHCqzibc0PrWvXV/+xMdhRBvdYk9X0
JSrMRscUsktGdxbZYTpsQZGWTXbXM3hYKv+sOtnSiHorp2svktMYjZyJBdqfOgbS
hA8NOERzqmwDx8Q1fkdmZZ3KAcI1zbyXpj+AIosVCMsSiL6o5lUuXC5TGq44LDoQ
6omY75w2oFue1/dy3E5I/WaL0avEKP1FXloRdrCNym31UmO6wYW5nf9wAAvxP0kw
AeKTEi5/jPjXxSmA5dlZ+BjXtZeW+BhOjacHmSx6ro5NYIboCLg4uEFRqK7sDd7K
gSn6C/oN9fc4VhaV0roS8JFsJaxm0K8rooKoq6V9Vm8wPPNgFaznwZz43n4h+4gC
qPr+nPmdzAKFNRwNNdmiAUpFbaGu28mV8oP4I3CQfkA4fEjNHhLPmPsn1gfztC0R
sbPjOXAzD2Rsyqwpi1fWaPlrT5JUfk/IBautskrPfR9fzF7NdKoagrQbAbexO2he
DqPFi8A0gPbFDg6EyOxbP20Zh+hnsXvulZJKHyIMeTZkCARh+tSaVoGY27f6WOI1
zuLhbXV2EZTWq57ciQUlaGCslmA8/i3B9n8cP/JmFKsJ0lJ0IH9sjVOW9aYGoFGF
rpS6hq/u+Yq5Bp6KnE4B8rAqVUHUDlrMpE7A4vrWZl+dVSpCLkDkAIKj1y4meA2J
Y5nIGHkEtr1x2go3Fk0Fr5PqWkR0vXJizBgSZFePi21/PTedvg/H5ifMjwJMpLJk
55mtJS7bWTLWpoQh56uKP354n60eTj/YOFBzMJFLWawNfjgCxV32ZljRmL2vB0ei
sj0grv3acHbCxFlPp2Au1M0ELL+kYJ4Fiwq0r4PFgdsTfPXTlpzcqvdls1PcfyHp
LhHhUn21HmPe8fppOkBmoC1mQ4YFzl8T00tu8s55tiNHs4LlZYD52VExyPRjeqWB
s/h3PwYXygWLWN4Ks9+C9Yq5xipSw8/CdXPQ9OQaKSmOu0++IC12fnR/3VD5wT/v
RWRSvR+FwG2ofnkLXHm4jS/heuJofejc4ILLXhWd84YScfNw7qymSwwCiXFguTE3
jEhaW4VGaLyN0oxvrf+qQtcccbiZtZVK9MpqSshtLBm+lcciu+lzzrz8lMyaLk1o
Ly0TW09pobR98E9k5FbZAR44nVnsJeTjD8mumBf1ftKjf1+zkRXQ9JBmBHT9Pexf
p7kBSn+pw1w5HhRbw8aRLqrXBdKXX9hAIF5gtRV5pXRrL2FnPBR9cSsit6ZEyHnK
1l9vMa1BvVJ0jpbDRRQbPds7qqq7Zx3e6lnAA/OHF16D0U+GgsqBX2BVgm+ehIk5
0flO8LOFt1yrknzxN7rkM4xQOgeEssY+EIOr8n4BaKHFkcWQEhxrAVhLNbQpbO6j
IOreGWlnOfbF+qQWL7n6X9fVtODFpY5E1LS6EmoW8wGZjpmdyajywp2fQWM/uPF7
I105FRmki7jId3W1hdiXIVbpWwrMyOuapxiEvVSAwAvCWPl+/kQpAg0No1ma468P
VHieR5q02hvMjFYax6qWh+bV8JegNw0WmdNoFbyRHfixvPMybrrh7LZNxY/Xslc8
o2gZ1TGExmXOZjpyHBjnRr6mgpK9yTq0II8fO3xRDvPUjNncBvGmad8FxSdvyzE0
t9bv2J+Et771lURxS6q/L/1leKNxVHnpDy9eUFlIoxL+98abS3mOaeEMygdpd99i
TeNkYBEVNgq1AzfUlPR/WJKYEN695C5VQNQ3PBZJBifM/iI8S5O3JwJ0D1Agarnp
uUOtfnXd6Ttj+eIoQacW77coe9uWUEKBcoEBCS+qUwykfiooBQNO2gFTF71bJH6K
ismo9mR6CXX+If4orbsWxU3olKb3uFkLPdJWojKhZEROEghmdpJaqlcoZ7FOaYWH
CuOtYvpdlyJaAMU8c4mVdQGSyXuxalApvpgF+As+C93YYItn7eOcNw5xw4Vq8sZF
2hhUFhXg9TpzJfQN4RGXhryx8XyQjvZYD1VPr7Y2kKpOyqJO4BiIDdIJHHJTA4G3
btVR3HwVCdaJyy0UG5H/+2FFQv2U9VooR7f6v4kRVox30WVEDQKnMA9z9V3hzY2X
diZaYbz1MbJ0HC9W8WNFRr3PMmTw15ReMc3JRRPvB6qk/2/vhB+QEPkXoeLMWLJy
XtMx0wkO8WRulK3xXJozNOvvfjLFsFUnvoNeEwHdBhqc364r7Jv/yPxjr7gJyOsA
Vbc2vCfE26J97tkwfiJRBXj0uOiYfEDo8FJt16r8KuH6wyagkcKr4NT0oEQ48h81
lwCI9xBvDiy69ht0jYIwL7SOaHMFz3lRloufPao3qzws1x6g8txd7dJwIPZez0WQ
sidvdZ3Q8/1Sz9AvkDVd7nIkURWESYxOsg4uM0bZAhY8VGRtfyzB8RzAPzyXCqt9
kJw70yAnWU2gf1m9gX8H8pqoCPK/f2iZucqb7rtbr9GEj4ualsQfi7CwupdAJA7s
iJXhLX5CAZXDgrnYakPijwzcOHFsdv1i7SAQizPyWb1KLuUeR5IxWBZysIJSVC6T
ivv05K4+MSFVd/a2VuwgMwHz9cBmv9UM5If9HWhE7NAA/HmOoMMM6hhRmVnhb30h
XCpsjI6Bvl3pJuv0a7SgPGyUzrUkOOHV+voAf28MRzIJnv+7zYzPLfM0DmW7OWz3
xe40WEAn0hxmU7MJwdPmDJ/4hyNsGXF7x6GgNtPKKdH1mhNWUswKuxRk5qT8g960
o9tSnW7/Ua/AGUwI765CoqehG8V0bSgbZGOQVopuyK640+19NjnLks4VA9F5jioF
GJ5+Q64MziJSXewjiHADgjWBjQ+U0jFvY/tGC3cMOcxr5Z70OUOPq/ImJ/6Bu1qP
0uv/9JgXM6pmjxsrX444FelotW9EkKdQ6cz5cmR1/Pb9gG4R56U3e43W98/I2psO
nCxCfW5sadVvY6NwZP9sP4uUxAlDgjGjB3/lJ7KA/QE3mJM44t4TY4AQZy/M1CfY
FJtw5wrRNCkideY/1Q8LabagUTo9G8hISFJNjKUR9LUlMIVHPBhPFXhn1WYYr20f
pwnJLYbl3l3Rkg11eP1oR2ntBP2uuZpDzNz5BTIifNcXEW0uK9KNAV9UJSeN7qsC
3kI9J5tx5FimAV/EnliBom5xrPtSg0AcgKjcPpaK+4gFsZSwPeQKfgqfNO8s6Xwp
QAWkD6Nz0ZVNajuuC8lEfeB1VPfleHqiOBtRUI0Cbo1jDGQnXaBWEsxZ8dKk4dzN
JeB3WMOTy7TV36ymEx3RCuHCcrY5rBAkbLYOHz08oqB3Sc6ofpQTnvG7kDu0OZ/5
AtTln5ozIj5nLWSNSvPQkA==
`protect END_PROTECTED
