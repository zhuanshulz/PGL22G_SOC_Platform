`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YQ5kYU4apCIpxYYNzmWns0Sp2He33Oe82b+C3gHhfvm6noR/T4kCLXgOCbMXmA9C
uZ6YX1HuYcGnAD+GcGZK4O1jYwj1Bmm5o9nWavvtvmv9jODzwx+4FU2Qn0Ixrgkl
kDjjXgz6G1kCQQRM4nQTtkL/z3mmX+7BWbPAl8vwbBo4uwycpg/NJa9ugSb+xFCw
rSxxbUmYnTSFl47HdSnh+zjzmonthEo9IR41OsTE642z/fFdESQx0JXpKtmiPBCu
VJNXewMEELejlt4tW+L9CpQWOsD7m60FU/IToMznMUdvQe2Mgr9uyrhKoBrcTkaZ
P/uwUGQcUFDoALZmy6dbyBRpzxtGlbQlDAiihUYWL0S80569QJJ/k4hrKa+Ajbpz
Y0vdeZNOZziIm11rEDpA0NmDibPTJ/9eG4x0nonvQlKD3T2XUgBBpBk/74xQMzxD
l5USjfQtkxd0mgJVGfinnjh2GNdLKQYCCudZEGrch5MT56U76Wt+CVk28EgJG+Ma
u6c7jf/LENl814anqV4IK0KVmIvqONOxxPARAxvP+/XzVJDGv6F/eLVuoPJIRQFY
f8bZq4XAeRSynC0gw1knUMlEhMM3lkDcEq1CKt5k+8WV4siwZlRRtVSeoDOGI2W7
2TT7bS86FbeNTbIb7zKGde5yimM96xKP6eHwqLQQ4VVHQQi/UQ/NNQDKIwcqnVaN
l1wFj+1R9eethEAWmK+Damu7bETcmnRWXOq+FVhhrg64qGlVsQZPBTteLvVUGfVA
vxGdjQv/PIY+RExEyET8sFfoeKL9+zSxFONUSNALwPQEvAw/0w1pr0Xm/R6N7J/t
yRAMnvcu+XXNSMuh1evU0g==
`protect END_PROTECTED
