`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AJNOC/Spbh4bf3ctwhGqpHbS8fwCT1cMVQTsc/o03VpmzJJYGAlsnqxUuoM3asdI
nZjON+WJKw7InHMtdB2dyXBG3Vr4okAhqZ+tUHAd8zjC6or8vFqz8u9BK25vODDy
KKYPASlgoVaynZZ+IwrRia/RmULwY2VLpIV7VeddEfrvp6IBRX0SwICy0KvfG8bU
CIIGd2fJCLR17nfPoBjpXbCQ18dhw+l1Ru5Lt2AV7+Q8Ep5Q1ekHJL2R7xbuCLXB
sldDwmDuj7YacDTQSWWj68wFeR4RFz77/OivKnZnFwCYtx2APKUM8615Va7J8epn
pyOt5NkLVLjj3byykJmMnP5XQP6Ou/RTt79IN5jiuKsLmHpDC5KsNyXtW5CY9axP
LrYWKaF1MWbkK4KmrSMVSHQe7DNWwZcx0BYu2Mi4us+Ms4MeRhko2/SaX8rgcUhG
7gwWv86h8qCZDvQ+iZUARnu+OmwzonzMtwMvrh5dnz4RTIljK0OnJPp5QHzfBAE6
dWdSjHNw0ZVSDQzeZTv6JW9lGHHvfjLVHemoQrL/gOssXt5tXquYx3XolywiHOa+
ZBSBHel2tfywCi5a1rfsqQNQ890xp6+44EN+6t71Q87qsaL0lq+n0paFMR6HdD4I
KHSi93K/VfdUq8S3POHXnnMEhu9lcGx0VrYFVRACyfZLaf0xLiPSPi+u6jN0LhqW
tPuGMANkxZkf4V1yoX6PYaRxNsIT49E/AXEwJfUJoE5dkStQBinANrUBmLWxqTeM
h00gBJKedSSAP/xTlY+Q1PmMv05UiyxXBQec/IA7DB5LunX/szozjEezGdLfQzto
BepTCxsHvMlD51oiVrQJ7M793d6Nk6M/4OY/rvkTC41KDwJ847tmv/4XiuuU+p1h
Tki3aK3khXA/KCOqUB4Y+Wt/S51IHFgiL0qy65yeb6IjDNEhpQ3Oz6/afPnk64kw
i77YS3ompC0RcVK7ststTqwg88luRRM6jfvtV23uv2HrQ6QivNWLrmfY/PedFHcS
0c+9taqF8xv9erm4nTRRtoY8PIcnZnu32UMFu6t/ZaFC9N7uoz+MuiPjGmLVExnk
XCL8mVoVLd1ehWB1XJLwmH41lyeC6IyBwvnc+peyFQnmllu4rWbVGduplzO1BEo8
d8eMXsOSBYOjCCESHY9bvWTBucy34/Cmc+6nhr/KWvp4wHbXD2h5+dA42LaqvlDn
ZWuwaRe2Grf+KiS8hpgReAIEsCCT2GgZSIbmQObByT4ExcKEaWMgL5mzXHkaG9gt
qHmhll1LtqoUdzygzUuXCkLVVXE8PGvR4fKq2LAeI+LTR9gCB3AADuqEKsyrWif3
MwafeBFbro1BhG3kLH2BBQzT86F9XHVsJgkVRym/FB74grpkvvbKdteg7DWm65Ku
tFfbB0mEx9WYYUygp2BuQWztVScP5KS1N2yxsRav8Jvlo9FwtHGQGnHzyuFxbf3g
`protect END_PROTECTED
