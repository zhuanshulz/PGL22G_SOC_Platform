`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3L69XH7Yl4oFlusunJ1U59zbSnZJ0hiuQarVRS0qh8fij3fTILCNykr6rQwrQwWA
uPzH38/CKBBucuKzI1M7aG6hn/yoqwQa1kNFfG59dho6SnPvqanvUvoqpXcQKVFc
JbJLeplssR11lsoymLfADliKLxc2/lreToGpg4pcef2t3CEbnR28DzbwSKEYItI2
Wz9CfRSWn1B8bw4mD2oz+qTdVJ/Bn6cFnjouJjxPz8wbisoEtiRz4qDTZWiqY9//
nNIYl/1dJcLnxuGy/06cCatqGmt0XI3r8TfA7u0m/zlru9IckFCAceadsS3GbpPd
7BnjV6ZFyhAeR9/OQkHZA7sIVgXHq6nXnGmnaJ2s4muJ0pwgv7H2mze1LUTyhUPG
Bpu029Kty+cfgFpdqQk34axGl+V6Dus+RozMVum7n6v8We3GCu9x87INTAc8x2bt
6hYFRWkKQmepDTNqD4a3P5SlRwgZ534pL/pYv0K93s1bEEzxQoDvN4drNzE4lz2I
ZwTikCLA0jvTzGVRM9QzwiFb3qTHlWBIpmWHVAOWtroDBMwOnpc+a81tUSFoWkih
Q2NAV8e7/P8EjLbdaruvEbj/lesQKnbEwhOJbRnPMALdxM728qmmwiJsDGLEmnDi
HHKDXgPpKQ3qov8onUU8kIyHWOINsnL89tJMG9/pelUwqb0y+3p4Yj6R47yRoD+S
mX/bh+8I6JQ4317gtCX4WN6qDHiYrWYc7yqLcuJL1+cxYGeP18yJaCWCJqNi3R1c
IL0NFVbKnzmqdKTV22iRgLE34ZfJIHwpmtp4E29IdI8CQsb9tiP8u0mryK2ovJu7
RiyrC+S2XPDPWCTfaePK4Fl816bt6anu4GVGIrpBvDSLu7yjNXhxpDh5PkmUU8rh
7d2wFl5tXjVGCZeHG6aG5OMFbynygGaZ8SFnBrFTkAD0+yjitfgNA+hU2553iaNn
qnLsZxiIguFFtMLcZDAc92eYhm5AnbkaMFG0mok2I42mvHkmM6fYqioxYNuNv2Av
gZ5UFtdidCbq5kYsPCrJcxovYaMCLobERx1ufxe350z/oEMDO7vXoF3fejlE2/bB
HE4pOilx6MS8yWKLwVZDNNRhLEU6Ztw44dhS6Lun40Mw3Z8riLv7r6C/YS23SqHw
TJu8zn2QgbE7Kam5xEHs5Av+zRSs46UqkRIGoecpYg3ExMWQQ+MkeDQGuYnf3Eis
BfFt4lfPMTYuiJpi/beJ20QlLBFeQW7y6V3aBRWm4HYGu4uvnEsqvLbhglyiNTsB
7gxf2ruNfChwnxAq5qO3QIFudlqd9UgqExz9JUDxjVeVC4HucNmkIqwCKP6DH7jE
um9T5yTNPUq24HnsZ5R9M7JMUWEL9+fyxX1RkMql+eWP1YWcqCSKqADA+v9SPWf7
fcf06Vlz9fXDgA4Kesdff9sACcz/C6PzkUgjZWbonbtqQ+hQgYwYWe0k2ITXTWQq
yczhkDbQR+KH85OUa9zgosi9uEAuNlRDWGpUsBNQHoDBIoNJr97jhz8Rhze9hwEu
0zVCCTA028b058dfzGVXyMZ+LC7VXY5XsM5tC3U/1vVRjN2ctxNmBzwLRhxZRgZZ
eItMkdGgEIxRfzc3PnEM4tY9ul8XWIT719p2dHEni4A6B6YcGHSFu0QuFaLuuxFc
VT7by1StlLOxmH2znwImT6f+D3R3PvwjUmqQXdwIe5sZLMkzQBpPz1ifJqWZ4DFS
CBKE0B4uf7Pbm0lsWLyYxH+vyutRVMRRAK9rt3hRVF81b8nAqlCFWsksgrcwADez
/8z71BcB+t9zL4W3RqzJjurXBz7N5lxYTVzzbXzCTFc30HRTaFwzmfHC6QgCO6lq
1WDsepKbLZTCfZFpdqvGScNZoNl7tEYbIZVTd0awE1p61T2n062qWe+qhn+JSeg4
QKGA8aL/4IdeQAGkk0y54tC8NWLVDS4NiiSzCwZ977j/WyyV2BNqhWiAVt1zSMhx
fJBfWhUoYC9wwhVvZ3p6KrRyPo0D5iZa8HS/6VY9adDJj16it4aSTA9fb2KfjY5+
CJQObRg4tMuGzmah1dqv60U6uZb/thhs1AFiFeCkyo04lrtT+cawTKtto+Vp1O2t
26QD0OdCB3DEmhmF754wgL2rkTmIF6W1dlTLydCFChTSJzgYBzK+JUmprQ543Rh2
FotFM4YoC3u7LW1/xtrDr0Rc+BcVK8oobSMv3Za5R80vWr3K6Tg0XlauqO/BEqF2
cDScgwVgOfHT5vYtwP6m3vANXPHB4WDUcKouaPvLptJbt7aJWTB46f6CI0m40Tdg
KwGjg2vbpKriBe/QmrSMpEQlOkz0FX5aZe6ZMdT7iJKxDHriH7VbGT25zYyuh0Et
VYoQVD99nRizqLgabx+thra6CTvx+7bxguYYKHoh1yROlch9hMed/4fyUeRx9umw
r2TTE8y7d57vSwYtGVUeSDL9hgfziVzE6iAkkUyJyFcJdK6LXWjcsITXGfMv5Ua9
gpB6zeZfF9UJuTFIcX1EmZOwCEky52vBvDylF/pFiOzFRlxd463w6Ky2/C+iwQqi
NN37gZQgAdqUZxLbNN80nsTaPXnuEOpI+opCwmQYVyqXm7igDn1zn6DgKcjjiRus
/fsKGtFG2WWZUvt/3h+XWgnmleaHI6Bvxfk5uleXP3OdNQtUDZ4zPsN6i8DaKhRD
LTx3CRVfuW0AnFAzLRtJYbUbTLV/78J9D4l14TWx08zThDrvBMgKH7JrMNWbAz/E
OcOAY7c0ktJNm0OOk7kSZzhpU3Zxp+jl8vOzk/9am3M5GyVKnmYQhY5MnYpgYU5Y
Wq0J3iGIwu6YAzmcm6EBwDw/iK1+yBYtGDZa3eIHisaBFR2hvp7p+iouS5LE+Lkf
w/sHXTNCzwqN0mBpxrD2AxWAQG/1sIQTcE9qXu5i0HB0SWzQJHFnIvOBk5s4zYp/
Ep4PYnmQzELfzkru5BfFJhZXrkMZ8VbZG5P9iW6FYfxzIehh+pE3nHzmzDapiNHD
ZOwTqxWuz0dop5CMAWHDiNB9ZNGlq/R3ornRLAfQjxXY+JEtJ9Y+koQ1eBJWUrkO
lSokb4ZMbauQhHq/1iEl98fxwPkKjQzI1TtVHZ8DrSc=
`protect END_PROTECTED
