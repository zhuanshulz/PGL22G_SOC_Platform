`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/zrWjC0F4IQTerfojhKhVZUHNerPAlRs2hKVCE8lWIRXOjytf6bZaDNibQHhlYx1
g7oJAxwegdu8SSTQJXIJqV5zEllv6L1ZoqxRIh2NReu05UlYq2JMOwbd6GphRCkr
Zy6m/7IFcsVVd7NzXL9dWzNMzSyeINB7BFH9v0SNhDtWd0NB4LdR18R0vKgPnpGI
HByjodw7xCbg+FTedovJweFadrbRr061Bj4AAN5T2Sq36CKbX5hw71nIQ1S+RyJ4
JiHl5JRsQGkf77tB/SY2KXLcr7VaobZGUrS/YJynbKZEsMUW5PjLW6qvWPgYjHDP
Yn6MqzpxyqxrZjiPVLgC+G2VojhCfkV67V7P7LNUbeuUYp8CeifA+M+/M8uSbidi
dMHyYrweKy1psQZJktcyX27JS97jBqv/tpi69egu7ITuXV/b4pj/whssAsGFFSRv
tF+zwU/HA6p2sXigUrZlCgTz9OVSS/ja9eMR2oLHObmVmmro/dMI4+GYAAb1sGbR
aiegvQaIk0qpooyM2+cp8S6Fl/6Ly1dOBeGc00uzRFKXVOILgDSeDzJ4lNDzrFM2
r8e03AEq8Aai/ZZxkntQjA==
`protect END_PROTECTED
