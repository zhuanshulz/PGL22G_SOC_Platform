`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xbzscwlJM4CEjTZ35hc7T0E+jfE/n3wbbgZr3QndTG3ybQORMkXmXDk3Bc8krqQJ
BHStCeMWvfHJorW1kB+ONi3X/rnjieJzunvBgAt/jgOgR1FqI47WSZaYcjIjMJHt
UuewGG+joF7Pm7PAaBIATTfu7UID0tIFN4ikDg81nbGBINEVnWQgTdVdb43Re3Ub
eGdsRUpxiKTcLJfdZIs2WerH3XnXHHHV8yhSQCn/vXnht+tU4q0o/fciXYunCFFE
L+gRP9MrS0i4H9OtNNZ3LqZ9OTsoB5snw5hsUss2yihoOfvPFMPYIXFinQtX8Fiy
/IoyJr5o/9PQuC2xu6BheL0Moiy6fdIkviGFr6Owk0i+0q7tRJyFnyx9KbS8Kolz
osIxkcrWCDmxlHLP5UeJhC7sQLhVVQHYOhI8hLLd34oxQAbj6UmiAxWOL4Wq8ySt
hadH1sAeQp4zsAeW/0AoYvElNcPyR43drcmUEnjx7rFiR5ehoHffCoB92r/s4jvQ
LWjvhW2szVG78U4Xve3ajV9SvEXZmpwl3PtdkMcEw9oPKUPlkBTInKUudwuvIJt1
HRhmIizl9nyffzS86OjVra/V4Zo5Zrs5VMAqJwwCZoIAtGxRgpy8d2pI9pgAgARM
lxGfr1+ChzWs3WRij8OftJsFUqqRpBqoCOiT2E72GRv4d1HgHG7B+xOx7AG+yU/b
6+LogJiunT/jJVx3ydnLqD9SGWqn62CMHA28Cbq9TKigktmbesAcJusdHMhcym2R
KB2tXCmrccBO03LBq0Fc012ZRg/7zzqCfV0h/xAzj4DXpGsKfVyYI5BRJk/uRxdP
rb0yH2YfMO1vbdq6e6t1hT0/319WRz0ExbjFwNKwrBnaDdSHyTdPqgKInWKDlOAB
AeNhrSdUSV6lfVUaPxJ/f7hYHdWGOnwzXL0LGFGuvMV8uXTmUkPzs/RphruVze2Y
FgFkx/kpmujIM3pt6AJduq6aU6sw5j6a/Ih5RyBZ8r7mvtjxLDqvQEs64/dPYF3S
`protect END_PROTECTED
