`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IEzwhBhYwHmeQ7gXv7jLDzxGlH1tWK/C/ZrEHEa2d/IQnR6f0hfWV015iUvcS6Xk
Oo7Hye1RWxxJ7gdiQHQyUYocCz/+2+rOWmixPC4MkoVZnbe+3l2w51CIetGJytog
7M6zbHUuW8xiXngbl5I9LEA3JQFqelMPPeEbtNFaXj3pbV+Pb2Nn3iNJgIh0Z2oe
VKQm79sBUz3/lqA/bUvaHS/QyekbNsp4xaGsa2/39kg+nirhFtpQ0Mv14Igoh9aV
yaNps2jGEGHEMk3g64unGsQTfl4TqCrU6xx/u89x0rraGxbQqhahAIeGZM1sYOfC
xm0fFPGPU3LK9zro3T6m5JlHei5MIZAkyYbuvLhP2F+L5NcpohbPI+JrUASqpJfR
ztFOiGMDghKyLZfuLWyzQMsfFI8pjQSvC27QCEch/+Zf/ZrUDMPrMpni3l5hkKan
+KtGRgtbCPJvokxB6hZ8wuGKdqZ09JldM1i7rzH10URJ2T1G/eGZcW+H2ENshg7L
NUSNAqoCeuvTTXPtqVfP5JKiD131NGr2JOoy9svA3DGE62moz9KEsfUD66jKpuTW
`protect END_PROTECTED
