`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1tdt8/YojB4e8yV71jxvPccYznl6FGRPX4MYmBHzinKE6mKo666wGzG7ECgjo3kx
cVHcMw0FYp+1/fk6WWMcgp4tOx1Zartp+Ma1QqABkEz739rDQ5WKdK5sd3p8xpVA
b8VWx1yKYzePvDoEXwRSKu2SHglciCuoemA20RtrThDwl3CLUJBssvLCwUJiCxJn
Vcv+L1lJdgIeLZ2ZIYJWvJhWfy7B0f8EOZI6Pyksz1qArIKpTWUnqRT6VxVSwDKj
wfwoCtDwYFHbEBxgUwTYANkaXgj5ahWAWE7teG3FepErcW1R38WrKcw+rqUju/ld
/KtKoGKW86SkWOEox6SVKQV5/apk3IbF4+LW4puHQs/tH4WLvWN9F0x+WG/0cgQE
K4sb7C2JTqB8NjoWzpDq2NVmNK8LvAKHOZPasVMr8gCb6EtmcCp4wjtelzzwv8sb
0Dp9H/Q0vClpN5JmqzyIN7Y2Zj3BhU8Z3McCoB/+rlFuq0ytolSmgT7NY4pXxoEZ
lmxveH1sItXEBF9UTcpvhjtpTCRUuGoOWo7Dx04UUUoz+E86XtyCW+oKpQM31xzT
gYTAnW7z71qdQVOXBU73Rwr9N9ANZ60P04Umse/W15rmWKRvCiRdn3rksvqvKLS/
63MHPR0auLbdZKtC0rJLcLb4aGXDQqJazibsr/NnPS9zzNMMlPABSFHTZbP43tKn
c8E3KSgect8u6B2ZdWd279Yg93fCXUI+Fa6HlfnhB2LmpVfoACpO71wAyV3qtmDw
HKis4MWzqndUR1Bquz1f1sG5lgUFRb84wjXIRrXf1Qg4lXtKz6PzRP4ng/JI0LAn
zV/0YdHlvZsF/xm9tntxyVYJvHDKo3xi6wVDFioLryw7L9Vc2ixX8bD7bBLHt9lm
2Y0P4Z3DW4hoqXF/doy4vg7vOEBmzrE+kyJEHXnStgNKugKPdE9FpkLqLIxpy3Nl
LrHYmASFCltCYw3G4EMUqldUXdTeOqK5HWemSm+s6mGhWOEc66234DrgZTdREF1M
UN/zjbhCoLb80cRcBWtzXpjmvrluiBMf5R/p26SjYfUTFi/gVIEgJWzCBs2GQewU
m422sMNgZ8+iUMKb7PxUv5rmgALU0uUHX7Jbkwd+vILUaQdxMVF3kClkpyhvPnCX
SjcPxF5POoKmqhEzVpJ6/I5bBB8+phMSkq+w+vYJALGiF0wSMYkD9SgE2AlnRdVH
LYutasq+q8EPtlhCRobA8eD2llz9DWESQqz2lyM4fiRAZvbTFVBqsrKXDlEfSzj/
cuQrbnHBCZY8P45eZiuyIKlX1F9mjE5G0RyoKZzRyMuWH/tySAzUEU760bil/mqU
Ek1Dw4FnH9jk12P76+xZe7lvCgumef5yCvm7u4ge7l1MgU7vJ9Qx91yd+0fq4r9T
9om28c3ojLCX+hltnpMrZXkIk5MRg/CP+0gkEd3xzU0c6aijlf/RygZNKJ/CEpIJ
Wb0HnEO8f8dhv1AGYcKM3OyIftD0vckVCBkJghUm03fBF0Su/43H6pDFYlb69Fme
fxwzjbdcLWbb9WqK47I2Nee2NndpLq9UFrBZm2c3l03MiAjCohPyK8zoCtD1u4My
dKI2m5fM/Op1/clDDlLPQHr2X1xb3mO/lrj/NNgDG1QuorhvOOWvJ00U++jTcnKb
Dby07wNMNU/lLBBfu3izROgqnGSZIcmFNl2qbeCfyfQPnXYFbqa9jcrSZaCxSoW8
lje4b57m0Yk31eu4MKrEuiZgYVMp1PQ85/mDJj+AvkNmCWq9RcDqY1M/z31wwklG
BV4QX12NqTljnSa5FYVCTZGrim7m5sjKaDZHkXftfpOOcp6PvI5+A4NnN7K143hP
DEBudHRbZlXup4EBxTbnm16Fn8rYm084PocKqvBYjzCb96jJcBnkrxivdsEVRxXt
C33rOud0JN5/v1KpwAv8DfjOpxAUYqUzy9bvh7O09jti81ywYAOCbl/nG/OKlks/
BX8UYYnSB0UpZ7I3u1aKraVT33ihYPRESYk4AALvXKEPU6qFX6ZMPcyeISa8HZcR
CVrM53XenYids/KcbaAx2JalhsIMNJfeKpd/TeZU2+ugY3UZnY1QN+xIIsZaJT5j
2HmH7lgDy8g2DfBThvjeOfUJ2Cq/+SeSz4NkcV/vqTpJ79jkHyAsfsz7rRzePLBs
GeNrx/7YVn+fvK5A9Qw9LtzKd1wgBbdjMZiQZQRevy3//dwcTmlAYvcC3ZXNZPj2
8g1eCcbrYJuWRGhMvT1pi0/XJf/YHMyzZkugyKKqf/CbdQZuoysVnK8nBYfiL2RO
5wpbiG8h5c57JocZzOnKq63ScFgnWCVKMM8T11PGFacJjhdFV/6okdELgRB3VVtU
BwWdoZSmNUG6NWcGP3KNXcY8w1+zlNdeIw7cNgnwHqHVZ3xKu1Tf2awIpCykL3TO
17O64LGm2HLQzYVWiA9aBgMcdpknCJiP7iIh5menIUCNiDakfXb0YnWAKegAhsIp
2j2kUtZC+yEgP2ClkdCQDz3Tg6hp6GqFQX5ydkq1aWjEnvLaacrC5vGr+U6/fHJk
b2CZ7APTyww94mqe3KiO18h2nBjinb/2MqAxdmd4BwaA3yTi3aMzufsFrRVMSKdG
PmOFLjqgciWZIuW7Rt12DeQVCyAj+AHYXACHBc88LL5/7wy7cMADcFaAj76YeSJ/
LHW2ffG4wTwDpTzqnDjfhGeUe5aGNDUw04FhlYTpNwAGK4MDh+x2INMHQkOyZBby
oa5f4DO0ryQYHVQtVDRZ+mrimaEqsM2GrqT9a0SaYkjkJlzdr7D9Pd6GshRtvrmi
iuQsxM4yV2a2xSzWZCnH+miELMvZtrzajEP6Yh8e6T6x7eUvZVDJ4MC9hUe0ErD2
79vKbeWi4QX0eFkk9GL1/yDYVqDpfOJpYmsTq+H+FkKBdnGlU3/5aKptMVC8hCEW
rTEV0SkJplSj9UZd0etUVoHVSNg28WBJ/gWwaJORj9Mu2r2zh+ZV2Kq7nbXoXazC
ZXy0tXlololm+zhkbMnA4dEnQ0wPku9lLnWdFCFxJ5dkdWcdhviuAyeRTQprkIEn
JjZ55Rs89GWAbR61j08ITWqZ5ZiyYaTI0IcExjnzMG7Io8xyJ7OvG8uYH1CqzsT5
vBT73E4kZkwyY43FA3NQqGpnSIeI681jfekuAIqkyFsJ70DzIcrHdQSj710Tkb9L
q30V0GX63P91mxMmtIikHetWEQQAyZtwyqPYhwDOH/qd4E4x9JRqYKaOBZkU7FJq
svGSkjcqxjy2CyLB9bqTbpF53BcKslxvrlY75lRttaK3EHvKgSYknUhP12g5HpZo
S+9sFAWvagw1Ge7TTfxeZ8+Vqtl9UXpSmbOQyrBn9onHnmSuv4x+hoMXxBkHdI9B
DGRtac1oApQxZDVEOl26FDVXPWCzJmKo7zpCJ/IMw42Ge8NRUkj+VuunhxYZ4NDh
xWgK6EIsvFXn7VepS0GlQLP9kI17Em6ZZvpEhNkwrbtV1pKSMyK+6FAotfVwbKfV
dpZcUoKEOej9L/UTDXZTno+RkCWzjuy12khEWxOThbRR8jr+ATag5+K1PtJhcc3d
2i7ZSpibjzT7ZwfFLe747Ype34/qlxFlCopO8+JZRAMB2BhZE7Q9C7+FoNTzwpwg
XuR2RM5bZfuXp535OWp63oRULj579V5Jco3Bm1PPdfZsCiPhF3r++SKeN0HnVWIu
pOJoj4tlRpTZkQyF7oZYfgibGEjFHf/i2tf8l1PMmULRrdlaHhiYhKk/cGhmTZ2x
FHLqjIC9hVd2/HUBix782Xl28G0uxP1viM6l84OdgYM261yAklQBxgkE8vx9kS/F
jpuX3AvnPxJMYCT/p3yWmCVCIHJsAQzpUlP3ZJEWYXmQaqyEF1nqZ3nDxSDgPebD
RbfnjpRnbcgVMGIFigt71gFfu6yVMVRpY17KJznxFh3bFpPDjiU2ia1MaPhEqe5d
pp61eoxD9hEE/hYU1+PSR+/CQ6j/7LKEKlpG7Cs1920=
`protect END_PROTECTED
