`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ujW4ewHAynojr/tlC2pjSo3+QwNLzR8Bv9vQXmW6KSCYs9sFVBJhQ+4lA5cNFATe
fIfQn1A3z1VdwjVav/y4pB0WtCG/7eWY0VJJDL0lDKiN45SoROip7C9s70dVAghR
mWaGb3GEDMK6bDiiaNafNRHaCjP6PHzhHZGdNPDAoDvGDTzclmX09cNPMd7rgW6h
dyHS4pTEo3f7vqTKYQkwB2STA1UY2S3b/KaaOH+MRv7gNfP9SOOYAIx+0D7PQKhr
AFrXB6N11SFtu7mB56sY36Jef1fu4Cu1YJhZvApzYkSOllEd0LAl9NfJEuSmOt8s
+Q4j1e7rOKxxvbxvsaZsMWMZim+y0liDvB9fVXyd13ZZ2iIfK4cPETJU+dOYCtTo
Iahhe8t0PGExDYNzQFNIvaOMii0DafMIASKBkDylfF4siJ+eBKAA4+fod9vqjVVS
/JATgacmtGkEm8z1AaXnFfPQPfdDGv/3IoLbjlmL7S0l6kIBrX9lZC1G8NJnAgRo
RVYtRNwcnJyK5+TY3omoEJjPbZrE7ZjSL4jHlICjT2zuHV4xwrWbphbLRjV2ZmIT
vsxqRTk1CiVBYyr2O1rvb6U+Ngxj2064LZIy8PIzmgM3w0cTEFmSZrGisFn86UX0
HdIHWOhQid41nkipkUBI9QUfwD1MXM18Mm/SyyGnW2RmOJehHDTFoz7gV1mW2pye
Ab8T893pAt/JzLMdNFKbfhrjTNEzKDxvVS3924yiOmNpTjqWOgOlaHcKUwuf84dQ
s0zwY6d8os0TwnYC2fSTvttsl5HlAsGrO499Fdc2KQLfsfoChCXSCF0XjS3/7koo
TQ/zz2lolpVYMh9aU7XVfuRr+XqUUsPHpg0cciCH96vNJRnkOafe63OtyD9dnu9O
YDxf6kS9TGadmF79MuSp7L89nhuu65sbTsg+qkyB12dEHcOS1pXXtZEOQtN6h9oR
bjhNOs3x1o7uQXOMiInhdwtTE+tb/acv9C7lwUNU6LtZOgqHlL670Nt768j0Kqcz
ffPrJPm4lXeM/6u5Ew+PbNFB4seIyRZPObuCdhT2XF4kHXpcexRwve3VFRxtnsXZ
TtqK3gVbEXzE9/e1N8jZLzTeG2Nr0zcnj0Bg3iL3SqWKTQZd9Vend/zSI6p+I+Br
riSIfH+FgLKMrKY/kKFOFOCppteFsJppcxgRxMldeXGeS5npap9boAz6GFTxqMKS
oolXXCcBxbaIpatkRek/FHL1XCbSR6dHu4dn6GsZG0SM95doavnkk2x0oY32RExX
UaOC/PF5gqztO+ekke1vhPoD86mMcfLCSezP0VeoJwwPtzRtqrsBrVyq2hD7OxOg
905EQyRoG2ArtreoVVcbWg6cj1BhKI5q8G8QJ9Q+sCYQJkiDy1PzEarS6TSkGACk
mxGygkzeS5t1NRw377FAI4dCpLhSXdmL47fyhB25P2RVm7pjIQKHOnzSy+dJV5w/
xT4i5lY9MXkjXmZOf9+NE0k+jxIPsLGATT5FXh6vN7WQYyO3sahkfABkMOFJ090O
4dnCsPhgzgLi6hM8wEWL//+LYUq86oQgGwvIfsNYZEFgiUAXl/lpTqSCLIpp/D4y
lnSAzo4h1ti2Aque9kpQzYrVPghJkD1rtSNexC8QntMRZO98hD+70B4WPTgVRsE6
e3ZnjLU3gdT8gZPYTeLoxASbKzPq+5pzMRf6ZkJJHVb5fy2a8P+/w4UPKicGGJPn
XnDvy7MFMreza4c6wyEeu11jyXxdEL+owtV3oP34MCzbqetbwJbXgcJdj7QU+xQR
Cx9bzVUTV/NgSxZBT66tGo4gox9XJDk9O7IF97BoNZEKIl2EVkMhyxZwSRtzPamW
vr8Yb8aMVn4AvepOjvTV0EesY/uqTmjnoaT2SP0XbIcNg7IbwJm6hDFig+qVe0rh
a4GEJQ5Qvg+hRu17M2qOr6i3hzC6+jMg+qVa/XZ/pUnjMq+7eESQ0ACJfhnhxTJz
YPUrcStpFXe2R4HXUOtZptZTfXgkQfbgvGdwC4GCACloNlKeWnUIv2W3uxOGeQKi
25OqHbmKzY8/Lziaaet6Cjpr3LPjLZpclQ0yBRm9CV6Dmv5eDH0PRj5HkqF63Lg9
2PFuygne2i1MKd+5ekURv7sGK6M9PGC5eHwFD0Q1OPAa8ol+rRr1G5QxyCJQPRb8
rbTKX2gs8jWvwVhg7O9Yr4pApvoiGpBARd1xNykvPgemne1P7adwMODi+z7YSPmH
DQMS3rUB/v36OwCDBLztgMa+mgnLK1JC1KPhofGyVVm3n6FNezT/Zy7aZsPofnYB
6RdQ54vQpDboMcbC0uAy0KyJ4F2lE2JHaOTKy/zvNlaECPJOkuubQ4jUZoaqOWjr
CgvEVt9AK/m3gtP1OLjiBMqO6K8n38c4Zzxq0FUw+BIv7bZX+hBUyWJcJyPFZ5dq
Sjf4SsvMIZeTP05tOgpnBx2++G0C72Hv5NH7s69wwujtFFPMYzFHL4momQIdDQ9b
JrUVJ5PUiQU63lj/Lg6ZZCrDTuCwxfjUaAJUeT0mwvKUO9SnT22E9RaXJ1tawei8
4x+CM3XlSahkYXeGFf72rFfyZyvel9seshcXadG/DnHyFv86yW/bOVkmwPfoqsmh
H19oM/VxSNxm0U4trPWB297DbrXJy/BFosRazc7j/TTLsTwUM9kC8LJL+GhYzZwL
CxxPyVVocV69QDBfe5sw1vtzhqq6pyeVY2Vj9FQOzoxKyyXJ/dnWuLa3wfzXpFAJ
jOnEw+bOG9B5tdGIL7PYcneby+wTjmSn6R6IACaQ8wQquPeRbSu0lmuiWwsfbmfI
YaaeIVPrSlLWMT3yHGwdSo6NLWUI1L4BBfLHRsAaOP8krRpl+6K48QEoJ0Ktfy3q
4WGEoiGlKGsIGcQsl3BLy1zbxrsjK3W3Yf9LDZGWofoD/1yg/EDtQnrIhBljU3+x
WmQarpSe6tG9mJ2XwPGlS8Yl0lIvhf+hdSFjPoKrdJ3vPbBWJjCEym6m7W2+DqC+
SWRIAMNeA9XbtKMVbLvglEHurCG95ZqYRCdV20APpYSNUzHrwzV5ACwD0wcCNbgh
ODDH1k2Z7h/B+pgGlSxuovcPV0kcWzX81wVcEavKpSiN8IUR8qk1BOpZlw5rYsWz
3kxf85/Dz8FvuaTJqDlzAisr+6B5AFpSRBFY/2xQUs09KNHQ4bwH7llNJqxX3LRZ
yvB4Q/KEvmiSX7XetnctDO5GYsFQRiIOHEl3TuSUlpSSnWOjld3loPLqZfIy6zGs
hn3XueURewe1qsnnMamE6m9LVk/BiB7j8UL/X4xBueaP43+wNySyaXE9dCJQN18b
LkSsyI11RGG+QYinZCmzdyPrVuwHXZKwrpdUVXmhpIcL2eXc2ovp+Q4ZRnBOPgAd
bLouCI2Bs7US4x3cYOUHY1slJ7tczXQjkDQ9dPTSZkrt8Sr58nwclzM49DDdPSWv
BezXyZFnuQ6PBAkOO5tRYzCUNaKyvMQFnidKwSBKM5VWHn34unfUbQKYcYKpiYS2
WYvEJlq9OlWcsq6Jimm9jIYHLmjAuEUppFW54a3t7V4q6b1lXajPtPJuqsHtjdU+
zTcvykZjFzslAteNiq6Whht9WJzbGPEuXijWGfbHiiuGM6BBwIzYx3OQ4L2/P31x
Ro/3YFMBqiRQ/uZpWRKQ4DKbHVnLGrB12nRFtkpPEhmvC6oiXSZxDn3QZxaFR9cw
PjydITvzPYuynUZqHh/o8Z/6HAWJbnvyb+krXCHnhif6b9Tj9cE0QmNIuSwtekYx
To9cfacmRxKopNjNTyrnMw2Tnlv+BTvKSaCLZlc9ePIlFaOzR9NvlvJtozn19l8l
tKdTCpgamg1YsL2P3SqQbE9DvoHYAmTyGq53I6P26SZsK679xFedR6Rq95+zGuNI
S7pM2X202gxfF4ev3ZBr4ibNLK4w6l83JTVynnF711jIhGjM7olvDLr5IauYTH3F
t8FMH0/rsWMgWEs1theXX60osbOO365uv3/Li+BqYVVUMYgQWUnevHB8JxVM3Ef7
E3MaTRtTl1qccLP1rwqpG16ExI2UJ6yI3e2gQ3RFtgPuTDBOMm75jfYimcE2uDoI
bolJaQrxy9W+BuEgaB/q0qLZP9vSD2oxMVFhlDVMeoHDcO9RweEEFyTJ+ZTipWJA
/Z3637Tbeho9TJIu20uyXvJ5ZMXo5rpWbQeGwss6XL64bcf8fl7Wrj/VEq+lA+ZY
9xNwLgczQJoQiaeARBMRa1i12j+vRycTOpcUBLe2jUA4vdtPTTKSSWvzwzjydfl4
CNtArF9M7ks8Qs5l5O0hjJus7RFtEDpU2KkBS5oCwMfmlLGZQXYSXfOWO+69mVCa
zYJfzswGFLS6S2YW1VGk21MFnOVSsk/X64X4VO8bL/4A357QlJxU4lEHMyVhvvri
Q/MpANMkdW5j6e6xRgFD5xVxxg3Oha/RwPghjPrXBs5L0sLbfolf5hYgokLbBX/b
1BRkYmQfqmlWclOpLdWGMK8YHdSPEJYHnheF3vA+FFWcwNz6RnAec/YSZJS4/Ezq
lVBGj+ewhct8KJxIv5jOsoP3awh0BKISBSJpFuOeBO/Q5fpRbSBKAx1RiujDYY92
ojUi0S0xN0v0jslj+TVHXG7nbg0HQd4KbmKIscajzESohX7QUJcWXXwbDphlMVyH
tuz2Xa9f8nVra9SJim1Yk/h/fLhIdpTG4+keGkHHslEkltPmkZPY2EuJ2/ApuyFd
j7Kyt+yJW+ZDd7O/MN/0pMlxUmfRyvCm/puXMonbaDYcWkF5PSZI4lYq6JmateqU
YF2A4/PnkivrBKZMiljij5g50DED3t8r1iFYu7c7/1PJ8gNNL3Iq26vsjFCPSIAr
mVuUDCgnc/zxpCi+lBcyLN4nn9u+5/6adFZKNj2NRrKucuwNPt/sSdtn2NfUoeym
3piJfpmqt+XZ0biOt0iO6SMvvFVw7hrdWGM5IKf6vvS2qv7SEXbPxlsBD72JPwG2
tIo6HNBMFKaacjDapSPybQRBtLyI7tynmwlM+dhg/Y8lS7CN9mrzvKudjVAe9sKO
4zudAbGR+Ju81zDUb8YOBabERXiKKe9Dbjk4yUxC0sn7EA79UKjHzErDyPmmjVTV
nud1PHfpbybRQkS2nzXzM79haASIdhuZNxpUFEHdejpmhVwfT0puz+wmuUbr05p3
cAnBRGiG2Td8sIgamyjERnmdkkLlhigQ2DESUbRGPDXvIG2YjJEzw5oSmCRDaZ/M
OPr1zamDBdgr/bmqLWhR4a4pZb95g0MI3VW3AQ8I4ncGesI6G2J6RtluYP7WFIkp
s1s4SeTPleWk8lFpb6IRVNfftFdOdnzUg9S3DRNvOfON7XF2/vR2RqwOTpLfg8sY
pa/69bGmT51nJ0nAe5eFYqlrIPw3Y7hKBygBfK5+M4+hSUyEPVypmWRKIWG5QD1W
/qeuiwP03+C0QigHIipv/K8/x5BuXkG3hM59bWSYg6jvrM5xxs+wotojYEU76cXM
tOGsuWFNNtO+B946M/4vFLPeX8dRA+YCIPFvH0Cv8q5Mz2SunZ9+/zWLiY1FMXd/
lBWrBZm6AYQieyelMRwtuwzxs1PjcrkvTrxWmEjtvY0b1IFC6LOMQz/kbHpRkvIP
2wvzL9gxL3YHhUF8rwXW/YqsmykbCU+l0g+fkjVbCQkWLH1/s8Xt+S1ZGV6SRHkf
izxwnhR6pqtgwdI1n0XBSXlSDdtL5SG1mIXvrk5cmHENFNdz17Da9vetjWR8Jnc8
dwYu15rXzhtBmAG1NhEQgr54mL+FRpThjfZeIcbKmyq05nV2VBfCk+6F2vcheAn9
NxcnH7qYDGE0+O1MDZrkdez6GxrpFEZMjvDsyddi5Eao/BGcWSSLt3RgXEiZ2p44
rZ+5HxS9Aixsm203MgpON8coILs+7bd2gQK57dTsknI/L10Z5kyp2zP00KzYPsFc
2+qymOYTgTQT7DfgZpdh+WB6SxbPayr7jjgdGOQ00b4r/FLKQJiUrDakF2zN4KJK
OL7IePtRWBlSuWhzJUJl8yFgrB6UHDZ9qQ58jRrUGrZJa73ZnGjk1ZzT9EmTlJVy
zmQ3l4h+K4/tBUS0YDRH7J0QUGlvgviHUWx+j8R4ihYO3R71YxIe4zlEkwMHjFfA
v4z/e8eoHe+ShEFChhlSUOc6CsCWwBLD9XVl0MKoG1zri0mSwHHXnA+wbXJ0rcKs
x1WKUe/FUvZYsEWkO+nHicsDzrCV9Iwh2Cj5uiQWV+zbSVwVnb3uA/znxbFwGG5U
poOwc/zfF70HCnvuM22E4EuWIDfGxQBHWzMAb3T88XN3PMvq2CIvFIOBqBW+ig/w
eDoyrXD64/mGbGkDc/hngKxoe1C3p9FtYoeVG2qcpAau2L+2EaLtdWsIIspiZtCX
8zzrGH3oBpoeKScZ6oPe57JNqXNi6xpBfQt9ThqKj+YFENw3N76EBxwhBs6LnFEZ
8mapvnlpF1d9tzozkbEGXL8qCSjApScCoHbQxikD47UHvWh5yrQGdb0TXeK4gI7O
UzqWz97+LrPoEnsUva79x/QQQTscW33wM4nmkrQhP24eEHbgwwCvcSHTQ5MGlX3f
ZtzdD4l7SkgjMyxK+bE0IM3giJfrt4vv7HgoTip1OcfilFIi6b52ID5OeX2yRk/Q
gXGFKzpS/aIhuOWvd0CTmuGMo4F4wHw+VqPqmyFFT2vSph2kuRy/IJbLh9EohR9S
xzMwOAteF4b37ByvvnnM7P3Buw8VUsYSftv0Hb2cw8t42un+P6mDMb5XamrZEA8i
f5JGyDoSZuJZdAt8eUYejcuRa33npG3OYsJJvgllwdtWrzPXj1G+AcK1Ci1wozMp
+srZvikyaXu9crBffwkr/hi5DLCH7OxNro9oypWJQ9jcjlRItERZsa5iDnnzUG8T
+n4Qc1wDJRm2CxhExNYIwhu2LBNs5oztgKb+aml6W72yX6TZdbzPhVrT3IKjRoTx
2u3kXdkjknKNg2lthSF/inbmEMSseNYYg9Qa9O1PxAzuVZPWbCQwrNb8Uie1U5tg
/TuYjjmbxuLdwOzFkvKtvB+aLc09N2ZGe8oE5lpD9vmdLDyW+/Iku9+dXt4p6+zj
TJIVcbanQGBeuV/pesQBIGIjED4++5g5vGn7dQUJ8VnH+zfa+nA0r5y5CNx+0fIw
h16BY6VM2XFONSpVdYEEFCM2fA29LZuU2DXcnrM3MqtHoxZKm3tskFAG8kuhJdQw
tb7aY2tE4qgRiRnxqBAdykwt6inK2xAvKt1A7TsPxcTLZQvcT+NJOWYyJDC64qTn
8ODKrMLkfd4sonWIm3JsFj0YdoCQs9Pt3gjXtzk0iyeF1ae1TCn3bktVIXiA0noP
WhdvKMCxdZtHaAYYUmf/61HJHqIFgiGGqE6R0MI1/WFCr44xD9vmOivyUM5RoeE1
/Oq3PF290NnzeSSQauhumQA3FiWGHEnar04Bk8OHD0onjLgZ4Ee2s8LG5/Hbb5G3
LUPIzOpZ46Krp2msMm+S/f1bJ8L7XVKZVOzSeyAce026Y7M3/H0DJo9KrGfBLy3n
M7r2vnzrr/5S7Gqei6m7ZzaHTZ0bMHS0YyyblPInYhw/yzAnx/8SXVGWRa43vGW9
eR4BLibd/mVMI++aPLjcaRtUtRpYmxYXw6+FBq0hvvlOn7ws7oPgzI9moivYtmhY
0hEgz5NbGtlpffw6C95JmRrCBhc6KJFVU73bXjGpdXCWOje8CAS/+Uk7Td3s3HsL
vhCYucGitg0ppp/Pf4K7nAK1MoDRfYElx8AvogXwloXKKMZJXhr3flCWxqCARMap
EM61kzS+tMEJ9AgSJ6U4uQrfVaJ2Bbfh2bCj4+DGfm20hisWkhOPKa4nF23RCeog
3/skW+Q6ckCCrMGMLeUtmL349AVonbw/CYaVoyL8VuTyR8uFVbrB9TwufvTwQM0A
UjxfjcO6OuDmX6A2EEa/YIwLM8qYjd21XRm8cdAPTHaYmIWCPfocCmSnJQQvs8qj
Epg1vU7GFPrwbcZLfsiPyFN6HD60pthXVP55r/Y1zRA98xBYprwZUGMCoXJRJL6a
BXarMek0vuq8mKSYQDGanTuvjjGc/g+16eGoQX8oja4mCGnTunCwZlAbF5kgN99p
oG6RUhsFmLcUyKL/0n0ZRr5DPvdH+53gxvr9WAcx0Td3sYFTGK2x8saSPTEilYT1
wfYrIxGRbS7T/2jnierNy0aWvFsBWrd4W3dbUqrXjRIDCaAVNQWszSczRcxytvzl
+Zh2Xgf0JJsSzEUFJAgfEavdrrZkyRAGQsbX3lYDBKiFbf1mR58ZoibxXEk90sm4
Hzuei/qedWQOroefZJhwhKFWXH3hE5HwM9ub4FpZwjot4cldS/obKRZ6FPPVXwcy
5XdNNbQvFbkVcBqPhDZywefE5pvKuP78ukan9tL31t8/KT5/KLkR8cM9aVseL2am
DXB6vR0SxaBBmW1CRqqaiXZ3DszFcp3vBEmaxMbJiZtDD+kJU1tI+Uvf19mMzfQk
WhtcofdexY+MfPdcnc/JqkzyugV2pGCxeqwLiURmMxr5nMFWGEAY3UBFnpX7KH7w
MJQQ0v+mAbu/d3H5+OLR7EL3B0cXbNEiT5AD77sXBG0k22XX+mONCWdMm0PM2rUF
JhXBSygvRWTFxEgNXgSXvwcL01riY/rWCzF+BXAJqBqhAxiqSOPDpGQ7dvbDYKpv
4rAOmAO4LURCOtBdDf5rrlXeIgy/Gdsl9BjQa8zsiRcoVIrbnykT4wa79hRAt3aP
dv8FuotXSZrtyZJBMzh1/P3ToBWypnERFdCXVvWKUFmzGqILRzCXoxlbyKgntGpV
ssdTZWK1pQhqCSoIzIyxb1MqLJg5TQQ6GwU2rYduJ7feufQ856YYJqp4OZ+PuG7H
7yiN7mwQbByoji5/Cw47G7iwipstcxONAihmlE+CEFKDy7Vndk4mB+RvFNOfnKOX
D3L+EIWttHP76KOv8JAJ9j6NQrzH+4YYkutb+5aSw+I4v83/4kYB95XRwiv6Z1ZR
S/2F7KX4s/uBSSRKxMzvh2jXBUIU59NonbxdRzh6Dn1NEhKU7jGMF70vM5MFpm6i
5OzTVFZEb1ymgOFE50/U9o9nhESMOe2K671cril4EMMtLGhIWwcElL1vteg9aCg5
Ely4EjPRAISuPX9N7dhmNzkZd/XvqFZMuxz3NrMjF7dBwOM5gH/e/d6VkYJG3yuu
11CrzMfzfTxGMZea0zMoTTkKv+0Et5roK/Dx8sXjR7aF2zBVY+NRM3XOFz8BXnAj
SkPrLfe3t7LB3fw3FmbaG59CeapWKq09UTmNSuxAKTtqOUSdlx287Xnn8Zfj3YI8
Ah7GjoZjALGn5JY+7fZN4401rsvHJmhISX7AkyF/zZT1JjYgs5jOrRZnZrDVStP3
tKh7iRoWXQkijG6Y38MApUX1KzviWEOA1PS0g6Wl1jdWYsH6lYxlrLUjBamfYtgL
ZjR8wybNIDgiAZnOH+3JPRfRf5mVVm3s8/Nk0thm58uGkh8BIeXnKTOYWY1l+MQh
egdXv3WE9tfES2duzqdgeGhDpWSLhghCS8YyIZJFglPjRMlQh8W7Xtcwnx0eaGtO
DGQZq2geVAeF3ygdcOGakGtcTl0PcXjUlEgg6dw7WT2vRwFj2GQL3QDqc2zG/1O3
sRc5lUywa+uwlgT1/dH/Uwg0BHxoovDNfn0/C6fq4JkTUXrUvsCu71nyC+qFUtaN
MGjzb0Pm2gBG3JP1OEN1kffRwTc9J6WmaILcr9Bb8bZHRFLKkBbbc58UzTay4JKg
ghFY8l4xQiIgtMcF27YWsj6wbP8r6zBlj5+YA3lhQw8NWY+TRitUeTkuCoLpzmFi
UqmiujPx1ClJ7F17WZwWCiZq/IG7kd+3eJTlE9iWORYKnTwqXG2s8mULsro3b8t7
B9DJlBN//J9KEhEokir/wgPamzvR9/m46Q8JDTPFrAy5HCOFY0vKzmabaDLTBiGd
IZS/LlnRWEbMrnvIl3+wbcFRvKAl7NHaoonyEN1w9S3aWPctZoJoTxjrCcfz2b1e
j7SWVBQ1cqJY/ryFipnXwt07wWt9vg+T+HsRMLUh/VZKq9WdG9lB30FhqWUJm+WC
aswSdWpPB6zUk9sSdonDLwcLV+TpTlh3SrJNPRP+umms+BHd+ZGzp/Mc6tMWL1ag
CuV7ca+jV0N67B36JR460ay8GMio3l8BL51i/qd5rjtOMMgL3NR2fDyvtl0+dhLm
Tgqthly/iBTq4fo5xmH34n/vDor1YAQeQ9+YY4XqixxUwSBKq56fTg5O0nb41tvZ
YHQLEkXUXd2zwMtcXGGkBvLiuDcGwjhMRwg7y9rJ/JGh+OAS3M1cM9LmkZwX9x16
aVWn4xbGX2mWAXlw4P5kwSLls/9kPLWXxM5BQBz3RVoruvpvwklHHS32h51JyViL
VeFL+ThhML1r596mNhOP6TUQL+KZvSSHQ/OYL1a5dWCvlT+bDWnyROtiqm2NO4KV
l2Ucg59VTlRKrvw8jusMBerU1Flxzm0QUCBkjRDu0bwEsyKSuiYntBtMobca6m0f
ya+D6ArX5Wx/0OtdSrP+/87zfTfWnTUAJX1VHJ8jkhIEvP8tv2g28qwacDqoLikQ
DNUlxyWVvm9lWXwZgc/s3/seNnC0YhRtF0G7ZyNe7EOtO2UoyOzTyIn6M50Fka6c
oYbZFBha0to2tzLEYiQoXSZ4d4wKvIQSWCVjLMaueN7eHORgxXRyHHxVA4KDymBx
aXGnmll5TR7aP0HSbKetI/OruWkKaFVv1pvPS7fJiZ6daLRPkQ4nhKj+A6Iwa1iL
B8rzFKzOhmfBvZbIDkKOxglXxDHir6xiGGXKkVVOw6RIrZ9z83bsFKkcpOCuijg8
ZYV9IH7tcbIiS6wmhJxM/1+8IlnW/Ib9Bc7XclXd5RZsZgZpbeL+1MzLyOaDbqJG
bhuBuFe2f2msvfBzJz5K491uk2N3f5kETonILDz+EBoS1h3xu+dmLsfw6XmKbKOj
6FX0doIZ0+Yb+coNoyPFVO2pwDdCvyOzPkVJ6/+sBbBC1IgFweA47u0x90fXajmy
wDdzwRGWZNzY/GEG3g3WE8/IYpBz6gjV/FqPY5kuAsSHSvZlKVNLCp7JOXsXA7U6
Ha0nCBUA8KH+V0yBtyvnzNz/p4CGqQ2jnMlWXNxQvCXIiVfGfcYiC4glZO7bNA2+
pGqI5Eg4chwRNkPuEGlON5pBYNb36AdTKZdmhlohjETd4uwgjHEVJNVMHJLKLxQd
qjAn4x+XHK9OQa0G8AUAhgqn8dRgDHh1mXl5hchJGwPgwHb0dGjclJDKFCvlvZfa
jogEG8d+Xw+3Uwq4RIMq/N6nuuIk+wPDio9WbPa+goSD9cFzyEVheCKRBAVLO+Kt
wmAWDq2TVbK2diQwQNeWVkqPvYD0sBk0M+kWZZtftHgsFCZNmXrEdh4hA8IKZPal
x4A01nFbFzToTXHZjdTIBq87M7BPBkTthwvcUntDCO76ZoXfrLeJ+aRsaFf8uyZb
4kK0xoc3JndLO7naILazW71XsMkYWEZnJKhO762lArT3tGpHB5qP9jGWaB8as3+n
pjICWJV2dvWfTkBXGKZPgVc3Bqbu5DU/HOw9oQOwbntWzsoo9vLL/aje9B9ZvdFD
1c3BNrYqtTLuKL0wvAdUM6KoI676swTob/bxZTeyCDYlwNyiV9vEKZ+ivqKSVklP
S49Qnpz7w0dDTFmXVxpNtaLznphD3/xemugH+Z2pPZdKVgHy0FkJ6/cd0AS1dMO5
uuZK2nOGgiCVKYlW0Qgg1BKeL8M7nu5OOm358U537nvJwk2RKNXvcer0mzidzYzl
2HM1JvuV2ByB388o/ZhKTDjwQhG0Rw/PLCw1MXyejkRjxQmI+JaL0cW4vClTUlPX
Ag9MnIqR1EBNUJTllMpEfiGxzZbifkO16U0F6iyNoCurjt7YcEketlQTJBbC49Tn
GN7emNQEZajLE9CxAU6/tKuwmgLvGaQGCGLJfbTs4BAAO0492eWm2a6G5F0xKkkB
McILX8XNU4tUOQ17TMWjvx694w4Vi8+088XtbemiuZMvqKNjybloE92OJA0Qjefy
Rb3KJmNma2ruqaIbAS64v9BHZXd1JeohrbgwyUiuNqV9YdkOOGSaQnwMH/09Pf19
76OobDp2YzrNxvZmOGI9jWYe/lEM3MfixkeybLiVG4vWJrIEcvFn8b1HrWtZiuMp
R9Axa70C1S2Af9MK6+AhgByeAapbkVXqF64Je2Vcut+rRh4tq5ik/Y4ThRw90Kl+
uJQgGbWGeuHg/qzMnC0j5GG4fZ7p8lOZncd0Rh/fRM5PnUu3TxaJig7h9hJzynQs
6G/Zf86p5Osqpm400XfHUI0LAckxd0TxPFJmBFmcb+azP0mvKij8NBAEwK3okkxH
90gCr+sLbHHkGuXBWn9C39OecbhWkI5D7BuhAuHpZtvyxtP18hjDBbAHhx/LUkEa
y8i/AiDD79biSMHAeci0egXTpc2TI0p8bOh9x9+7FJAa1f8XQ17PoeGTwRzm66nh
qnSsQqQTidazk/A4P8j67p2qR1AO9TmsYxL6OQqRXXx6N0SlN6igjVtRbFp/zCby
sO8SBOpSSk7mEdJoneJEN+W0x4p6/84qa8qpg8eKzE7/1ritJIwEkG091YBw6tla
7IOaH7O/wlmSCd5T+4uKjYK5ME2B1jwbQFmAjiBS4L7LcKhHIl+IYE1SspnYZDGz
U2wCGJmQmyR/L/0eoP3+lzXMFGvx3rGg/Deqc7zeFC9skvgr7JWAemIlsABD/VDB
EMqJJqU6SS/AquhnHPHs3DwNhm5+V0D42K2CmWDDS9mOmXAMCsfbBh+5/Cqdj26L
HaIGHyjmK7gRCrJcBifyAboyiiq4ddAu4DPhpEv1JrW6ZNNR7XlGjILODDMfzcZB
XL4kGN3g4I4QuNMskQMqJ5hXSXzsGOLOmjGIGUdoEFkCrU5uuHIoZ3MZ/1Todqff
DQrPLQ4UN3udB/rqqgCaS9k78zLRm9/+f9LC6Nn4mHZxjNimB2jTC1uWd/k1PUES
RttB4ytPoSGxmggXfQUo8sy5W2BwUjKpEJNOjgcsf9RulOKcF/yMYXOVxFbZjIXP
JoCYDtuKn32vxOmwVSP5JlAFWeug/Cn3/LhbjAKC1BRtbZR28fVnCnIBkkmq+5sp
oUmxSxr6vUmvE0b3CqnUrSWujtYMxG3LsOpM3amekUM/v38klJenJ7AHhKt4kQjK
8d2I8eRk6nyCGNkUzR2cmo6dcFF/OisHaNqR9G5vtX3jEeUHeiW1y2tJJGoqyXXY
vfhnaOnIVQqJaGmYUqGtv6719yB7wOMgWJijX8U4sWGMtpWvVBmwHZh+zn12fggv
728iHAKljOtyXuxXN43croDhW8uSiRIPLr9INYg2z2bAfJWF8mwX0eDqA6Rxp3NA
Ih8nO80Bjkn0Lkfw5K9UmgXLv5SGXRNxBH13FffS9u0E55G4P9HQb4tl1yIRhkG6
nAUbyOoqPbTfqLzrH/FQKWc2UFPdjjZZCEOAXwSFc0Y6Rxo2adEcO2R16VRLQulY
UY1YME9kmzsMDcu8DAnGgU3JKBnLHPMS1dbvwYoCD1U0rGq3At9RHrMKhcUmwVsd
LiqcLJqyo3g7ZaKXB6F2Sy481pjYNCzLx9N+wB7aMkNpvWdDkC9BZKSlwh9xS/08
Nj1bfowRy9Atnf2AgqjOsPtnrF16pYrymP1tH/qwxks5MFs4+K+VxpLopGaHdGcH
GtAZcbetCZXjcLnHiB5GFrqDLKuBXh2rm5lIhz6VlhzgEc3C9DiSzgKmGBWGfZrq
/iT+114RbfuPeQHu5Cz7AmoOjc66o2oTeLd+adIjf85+coHEh5Q7o82AuILiRmRS
wK407vccZk612PSuZW/Cl9AqkyEIoxNLvPEsevNqA74+AVW7rkGWOKFBR46x6yQP
+WnqZCZ7gMbQehr8V72jgPuKKtlzTzPvxbqdjUFS2WKGBm9+fh6mc8y8OsOKVxHA
PCI1lbz6mW3Knz3Twgpgp/inOKtFDxrmywEJ1fhmnkZAmIOl+tQzk5vIeVa1VlKC
rlWMyscHu7GBJ8gzKIMg8nH8VfR2ssSewk3I63cfx86K7nE1WlBIBGW3xvwtkNl5
BS5bBN8AJoEd9KGqTcucyWPQcaCuy/DNvcMIRsKFob0dncMwxFE/26P4xZfeXUAM
M4z0R2L6pyKf5cc3t+sGgQDbh76StfsnimCzqE3YLsgWygWNC4LDIKF1glJXpKSC
Fqkb/HzPskdwOltFfTZEyDOYBvfQx9lLDPuOdriljyhaOaD2owPXnOlVo1z/wK4z
3OWUDcZeEbvhibk6f1I8oznZBXMwC/T0ET56vat8liY7e84zyaSVy0GL0wgpvAuO
yn2QaMzrYSIzOMBDIoMqhcXPxaK8P+/NnpZu5FEmqhOKNO2KvHXPHSkvi8IfsCcl
nqZvXeOElSNL8sQo/vHZilafZKaWCXgZdMdry5xwxiKY1qo8hndSlyN9WPj7+kHR
scT6lHGEA0qoB+FJLIBseHf52Ie1VRZozBfmDZsGYSLvSU3QBoczqIAec/F32krg
iIxcPXmvvNiH7mIvWrDz5p/E+tK32F6baaPx8G6WqJy2h6k8SLlBcVzJpmeI4Hzh
lkRXI8O3rQXi2fL6Bg8CWgzhyt5DllRMO/DBq+b6Yy6T+fJT6hcxXGKSuq/rLLtb
5eIeSxtqE53k+FjG5EswnGE0EKEpTZ93LId1zAtT3L8FvUAHeZshuCKTNKFeJuFu
HxOQJnHpeDj2cTAUEKrB8PTK3i2p8Dw2nx6QuKiMpTAGnvVDQ/cfZ7bWq3IKueTb
RFSEau2f8mdsFi/lFj71CWZgV3Zl1eIbvSuzzmSxKD0w2rulC0Wg1FDHmLEXHFJI
LYz4QEppxDCdr7aNM9aM8mXAXBeaZFcIwrwY30OzCm21fdHTaC0h+HMAYL3aoeei
6kOOUQ7BadBlTE54ZJ9bigI/plpA/aj0GJkCqTLmgiJbrJ9KmsWO9fn8Y40PlnnL
pYcVFog+Jn9b2Fczt1Sk42+FepR3LFZDRGbTH80QZRXFbdbb/ej123sztvFGn/ub
g1TXzUmQQeMsBVATWzFj5Y8E6FAcV0JFPzwZ/oMGllqAxMAod//TEXUZdgFgnVNi
eph1KG6/6HdRfX7uyuttid2o2uiS+r66vKgF1k2p8Vx0cLtebPfRIqEvNIg3Jw0e
Mwza8jx/xO+zyk1SoJ8PI7dh0F/cMa2EBQP3smvGGASJFG9szhUyeyq3bYI+1yU8
rY8BaF4eIyH3voxv+un/lmTk6L3Eqs2obpkrcpvSqAxxx7f6tge//K5w4IpEQqY5
EN8+5ezret2WLgPVP0985NyzSqSW4qGoE8E4k8ofBaMpyfv6IJ2Y5CZlHvdQYsKt
6h8P1QKdgLpckuVe+BNPy55gCK7qroldHVXOOZBBRBSPNEzu2V704BUSeQGD/zik
oBIp4PbwMNW5IVyvanTDvzou12TIxXcb+Cl66O2jBENHCGbKq36Wjz+PiNqiMJBh
m6qhO4X8afXyXDzt1wpkxjD9U49jBUP172NRl2MHQljhnzjy9lDh/h3oUXHgFj5o
oSF2P3pjl3pg5CdeLIuLOra65UuMu7/AKJd0fTnZWl0tZ0N7o0y6Ux6bLdbNEPuZ
OxQzePzRy7ry9+FgKQFxxTOFFV+aqslWzAGRmw73udHnHeUtrZt1vgDigl9MqQg6
Qw5GpQxzfFXHpNPzVP+3cOYj8GqA66OycrONxyL2YqcCjLVp7yTS+HxYAsR0UFtx
DIKVNTXOGTbW3nSAaA/2QHZ0MC0YWsW/j8k03AoUSjKTxn0yq+h0JD+hDvSGoHUt
KEFAvQNIzxuh0OjHgBNAZmIJ50Ao2691lV/upGTvjUV/4s2rQnhRRbB+QN9gY6jP
kk3N0e/SUh5rpUyVj1BeMzMXDs47OCFq/l7/E5heg0HjvY9NlXPDuIMmwxl5N+8F
zy/oKZ7HfT7bEJkFS7Zrud8/7eZNuiOSI2cmZr/80aijB0OE3Pb2Tqv3ZaSd+417
aXhb/+b3mqV/5x4C0eeyfkfJ3Tspva9ucoFxcLb7vsqxV2zAehBGDurf21T1CacJ
FstTgM0Z7PqZn/YPX/HL80vvzuE9V4T9cEI5Pnx7Re59jWuLJZApGSaTQqMWw3zF
MJppVOYrcgW1/gcAuwxN6nW1ClcKX/NNpbT2/PiQvb4ySa+CRFhgTaz/7R6gD2qo
EyxN6e4ksDHHZ43/cjj9QCKBOD682o7et6MtH+tObQ1JgvW6XiEkaR+mC+IQ3svp
y9i94OVu+QAGoXxbiarjfbvJ2SxAq1Y/wbMkfz0vaJFPCbJcRjibrshTtZhFpTNv
SE5+evtTqxvJHWDjQauLl8aajyUHg9tZj/qp+h91pVK7Ds+DAzTfkoXw6lxKJmJN
SH7wGWYXFOEZVIRBUeubJI1kTlzOpJcKuLVqP/5sG3gaDFYzhUBijt9mxneTOT8l
ro4ytLjJlhpXjNP0wlsA2Jkpl1wZ2tAsOLDDlwcwx6OK7XygDjpF6ec5U+8rAc7w
p8wmdGD0YKEQtIaJKdLukq7mmg7wLArtyYH+n388w1iH67SHtG5Ykd7ftIE40t1a
XjC8Pu+UqdRZxzQYaGnltKHUFQYQPDM6D/VQ1XMGlv3EIUQ3telNXwrN7HgbMnkZ
xc01KzmWhaUHe4UxjTNhnaOTdkqIR6S1JWPDTJLuWdPf3io44W04BDMZYg4XqWnE
wVSR3jazVnN3bHd/iZ00zFbZZf/Hr+WFwYileDdfpB6mJAhqyjquupxB0WDz2MzR
mWft7LTykXix2KOheujwdh0Zth+T+KN/2n6HCtaFBiG9QMmGUHY7VSdZRRbM3Lgi
u3BUKun2kNabN9g84l9vB3IxYYz0PAIt62kT4HdQP6UB52/zpwYZJ/XVo8wVjpXo
yxoyo0MM+WuKcJNNUQIDqwT3QIdoNY0//zG14ypQmf4nzTJFJC/dijaD0sKm6xhs
sSRS/zNyEDqvSpFfq0Oz8mljl2RodLVamBgDTwVtX88sfq8A+md7NawSkqbNBY2V
BcrWiZmvT6NUs7JpUjymRUM6LjSwe3eDdy4u0BmARDrZD88yYTbbnKxoEcZaa6kj
XTGOLQ7AY3ZMpy3TdRbd64xXyMzLKVvX1+2nzqhNWrhka26DgwjrlYY5laiNUbab
eg4rrEGZeA46bmSW3UcV+iH13s8WBzQanZk1eQB2yX4jtV4dnEbcCbaOoQKHBJ1u
DuaMRoe4NXAjI+lHtmMmjPvp2qYvTkHMVcqXkDn0AXOMZH2Aei/c6u9VC9rOe1qF
G1XKe9QgOjOOg5PPQnUU+F8A5t59kgXLqUY49KSk6eRV4gHq72QajLzW3x7ZZV5t
4F9wwn3q5pypHN95RomVfvlSvWjLfsOJCOSY8TnwtXLsTKcRCstqXK4KCKPo8mVq
kIdeBBAfXo+4YSJd0nccdAm2lCZswLrRvbuh/pyPujJjfGpfy/2AI/1fuyZUKJt0
F6fCX64WDVl75z+KabHXV2b43Ama/co1opksXb8/2hhusDQIaG5qnicMZTStz8ot
XULYLlUK5F//AUZ753yx3GDWR2SI5RAMKwfiiCtIrCJ2d2bjxrn1vrKegDt1QeqM
8aKk3DsbGha3+eFCc3ntu5mGrocflY4EJS3W59yDnD0KDxl65gwZ6zrr0pe5ktUj
RfCYtrnrPt8xYtAgr9zYvED0JYGGRKM9y6goTaCLQizC/YeM8SBnWHiNFXBAoj5E
1rjhMLh+BFdZr1lpJkKObABtyAK7Qsczbl9+IrIJpg4JcmohlYeQBg4HR+6Covr4
NsRaDcHN2edl8iA3xzqNHy8j5oj8Nl6FbmOqHrY8vv3xdk4HtPRybMYXNic4NAaY
Pn4qqlW82gwki3+gxhP7gX89eBKLDnS6wSKhv7an0akVewY2u24XDfJTNMSJhY6W
dC88U25I/gXNvXm8dw+VdsZi0MPTBJevOjKfrXtzFx7xUGUEv5oNiWbXV2ibNj1z
Fa53J7kBLvBcTD6zgKX+juWGXJq10VW7PzOsgENPhrHT8v6Tnli6RBbIRf9WJN6w
oqiXKJDsLww6KAb+d+s3e20vosWaONxUu55zAsbMLYxUT53KNweoCfdAGU4uuPy6
ZO6lMm8lAwWQc+jdaIii0vhpN82dDd6aeEs9lQB5C73R5rWw0UxaXHdgarIn6qqR
JhvMG14Ok8kvGNdobMddabPOIj9KjuydmO9IA5ZY+O5xNsdcNEitKU14AnCXbsPN
hnEa4rkxGEvQOAyQzbItNV/FmaqSojuDKmgTAkkKjKxywDjCkYUD3uPNumhr7X/w
v3inIQwE6CnSFCSEzRTefDs2GumYt+V01ctXTs5hjwMexXXoIF6ija4vF6fBQtfW
T45OOXyvuxOkVTg80seoulP584nwWK7UTh8nhfR5eHyhj9NwefvmJNiMO2f/FFBi
XSqrnaITL5cjc7hosvN+EBLcieEyWgRvu227a+Qib68QWxI7BYSoToYzJlik1SfY
rMPSUMlCQJvJWnM10sfGXXiJhjhocpqFUUUwkMDeWX00CiAwkXFUdniTSOzG5pJD
0gb0i7gwluWRVKEqJcHMVzNcdo2b9nWXvHJnrRqOcce+vRpVgenV1S88tw2MzHhk
V8WcTuiH1coARUUGnhyQXHseTW8XGmaZ/Py9qXkKynGgEu5rn5g+TgnBmFCoeglR
4sw2++mFIUiXw3VTVN0JUOeC5mljqAbZC4mUhfv5Q9mMvAJsENYEqcxJNzw7NRaS
LF/pqw+fdOoqHuYZB7mn1X8TZwe/WbG29p+FS68TO3QcXtO+IlwbGaayDbOAb9ea
FgN+G2n4cpmsiAVTQI2DGsGUlPeeGpYWdaL32ePmmQlyHB6ZWlt95xnyB+PXzU4Y
v8zU4/c7d8feerx2uBrk5uHBIpwmq44zfxEFvVBEG17WVlZBUqcgKiSnBeJS5gg0
BX+4dEN0WPCsNkEhnqv6WOm0MH8oM1FPcf2ieMUrMmDfWPXm/7igiNAky1nNbVpR
2Z/vFGqT2WUhFAWcMkDlcyMtnIYCxTgmkPtlQnQRd9Ts6WztDzFGLyYaTd9MAbrF
aF4nBSYx/bhWwZ9TjJgZJiZB2oHnzCKcIJ4CmDdYdKFwhSeWUK5M83HpVvnlCfai
YNNkJDXl90G3sEt4yoiHidnYyUTPjzDnd9H/VU9n8mzOp9gUsxmloNGWzomsX2hc
j23qMAjU9l2DI6/gc11WH4dVxg0QKZierx+gIpuOroaAoMJBUn8tJpR50lpDzNxH
xdBLg1T9BM3GcToVhWl/KD6E107CiFpBGT2IiEbVyy9k/KrErroBKoWkCpo0fzj2
2KQR9hpIaKfATbOHx/8/WJWDfBe1XZ3b+XuWSicAy8l9J2L8jZ9MtOBX1jAq7Z98
7Z7Fxo+vgzoKvmQg9+hrs6KzbVQTtinYBGTo6ml8jf9mxfz3TbrWRRlaYaGw+3//
k54lGW0CEVaU9JEzJASyFMETnuTm6pNUuT2x8QwWwMzEZPcrgfxkdM+/kYPDrXtq
5jSV1OsbAEW0wWbR9QCbApHOLav2X4pcvx4f8Uy73ZBDPAdjMOHtdXxGgkzE5SAk
gY2BeS1lttyaSBdH5XDDLfrGr/7CEhNc3SfYIvbkNAvq+jYNeXpK/qBDrz8RXotY
NY6ZER323PJ8OblpD4rIN61ZctDPTotDQg4elrfpoFfF7v06oXaaf8jXI4ZhCVn0
1yrxjqb1dji4FlleaeoABGWXZJ1atTdlJJyFIvkU74Ewj3QctKojrQlvUx+ydLFG
3HwVY/I3NMF/eRxrptjdJeXLyaEq/a85oWkzFz7SIXa5MvhTnh7RqoIGb3ML1uX9
`protect END_PROTECTED
