`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tlVk72dxrtDu0xR/SUwB4amDGZZfdpcFqpOhv1WaxudX73pxTq7XRzDEIzXcaJ76
x9msMKR6yCcbqJOYEzmBiTdUMpG5p/KocEGAYfhSnDchIHJihwps+LV+k/50ObZm
OPvJtJGBjM/lq5RBfsy9GJ/8kPh+8bguc4A2wv22VSPt2/ykxxu9MuXv9GvVw9o6
TrnXSV6BwTKD9ezpBAMs+FYCM6C3mE7jzwba+Tp4FIm6U/Fknedpa7kF+x6+cfvK
XFGgwauMUna9foaxPDpOppIDMBq5Lvt3x+630Uc8EfGdB4HhWuIw+w4cl043gATE
HbTCI0PeVSeZBEEUiQobrlFdK/RQy/pvhGbLRLHHnE6Y+Ro2XGSP3PaQ25P/qCuR
0UY3OaxlhzMdfRpMTe0afcqpDTFYweAY9u2yBcxGWtuoe1fT2v8pbwpVubuhp4ej
SCwRtybGf705grwqchsGMNk+3JziYEOwtAUEZlEwgxxJyxel4ABW/sHjGJytkf9s
zXWPtJ0T0oKL++aPpCo65Gqm0+3rbPrA+3ariWoMIy9UsLfsIrr/9h0wZSKOZzmt
wdbDYfULCul7r/dtvCtD2OgTA0dvqMwqRbhTKB2bBXAewEVO50wbzFOmtK1g8AdW
wyExBh/nuDdsFfgFS3DIyGlWriXSFb17cVDL4xbFo7ptbWOL9RVxsT/Kb+beTiaO
d0U716lMUWHdnedh15NQF9xq7VVqH050i0dGrfvKT6Wq0fhPkIwJI3PWYOvBQqeK
9megkfdyhiBKRrKPMvPCbQcMB6DOFlNAezWvgt+VnRP0s8wCoCbTAyv4GC52YD0V
zaE0/lUIcq1asDcEYAJ9ea1ZWzZeHvqz+7TTfyCZk142/IbGqAv0DuLdIA1MSx4S
b4uOSzMxi4buLF6LMKKlp3DIINr7crnFhEbUV+arWJ9ru+k3EISa6JxwyO0vccNN
Rtm7e8HkxRRxyzTU5XR5YnH5tUin2ZSL8RQPrDSwgk5e3+OenUZ9dTdRMOi7oU/z
pv31jQQ4e/YUEy6yQVthAnUhQp+rtQ2WomZ4pPDLKMDte3hVV5orq1dA+mTiZYFU
W9OfMO4qHbrH1ns5ATIxwAmG9zcYVuGQj7/CbbQ/IzkLuD9MnFn0P1kEn/HsXzdI
Lx92rfSOL3j5gBeoRyjjoj5zTJUBBTuHbvT/WO6raOEFWGu2Icl7gSzHDsvGEOym
p2G7eASATEScwG/mmHGzGj8tdE4bn1RCAa5rpN6toUlJ7UOi7dY2bv245nednMew
YKbYUyTm3xx++HkHAQynP9nz9x2lONUOequv3b3ATqAoPhOjMkc+7ocpREtxTYBB
tEfFMw4UDkwn6MThz8q9o6wW7Uj7f8MsDpDQlcaVogWKm5V8VOE5CeaOzqTBx1aI
blpWY3YASPPw5TlmbSFikA0B9krbicFDq5mOLC7jbor4UwbPYEBxu0ZfIFu5Tuvz
6Cd8Xp66mkMsYI5TGGtldMVyuPaaVxOZntS+ie5ta5sh4C834XkTJeMcf72dNBx/
FoyK6Pl+2QP6SLJpKKHYM7j8umGy6N0R8IqOgI1qxAOF9ipUPR0Yr/d0mUtz7j/m
RwFBq+bNIuCF/jVT1lh04gHnX3vyU10+Oc5JwEEaPJm6gcKtTw3xVLx4Ia9/JFI0
TM9eY04nbz3bgLqvLW5iRv5D10XS6yGBJUu/m8fuMT04q50/lie7T+1JY2zWr6Yy
51pYYKbT7HmoxWjujgpdXDX1tJ0/BONkCWbRQGRG+P2LUJnZul1G/WM3L8Cf6Vfw
1mFbYUgBLaxngxjNd/2WBsnzzNvgldD3TKwhcMFksibjqKk/wArqSJf8Xi9z7Ajl
Z4nXWbZjPgL8FasIMjHKQ8kqtVK+9h+uslJwuDUnvD6t4E1zcJgU1c46gLWYVosA
w9RkFdtcTwnBAQ3BPXJxvbE5tltiPh70oOsRz9n5oOR/POaNXrSMpimfj1QDIlWp
NZMpfrDUZzuK7pXcfCRI5lYsdgtK4AU8+EuWruJkV6+bThrnE8XSyRb9NX9L9dZI
bxeDORSZMHWY3Z7dh47MJ6dOEsPcVoitEPfzAC6taMtegDxslqkhJFGj7g+Qe+qJ
08UKJPd+9/iiERf+jwapsUL5iwrGxtacI4djuQuFg5VPsm1KTA9Ga+8T7d5y4CgA
razzajk5i2VVsHB4pMCJ02Wg9rRaeL9NNQ3PoSo1GDiknFOZayMgMJtUpiKQn2K4
0PF9hZdXw7Ai5o+sc2liDts5vbKnHcvBFwGJLokgJwgWkPPCr21rPH9qlvCufwcl
MCufE6qcmwvYDMq886tJzjzU2BQDi34jJCwkm9712mRLvJ57M5A5x1PlMujm8MSD
6NFXNim5IEPm/ER8k+X7aoWQgRwuxttdylVT7yU2AapMUb3Xcx0YFFoFQVppnEw2
eAQYZ5XhigoRhqiU3+FI/opoDyDmc0NvGdKaec0YwEDP212XkbBDkB8+3RzFuEAi
X0FQolgoufZaFKK7GaRjAa3Cn4NGESvF4xvN+7rQjhoLkFCwtXn41xG4I7Z5l0ME
JbUhe5b0Nt9Ol0n/pVqRMl73ZPKUTVQCxhUe+LB2Cgc2JmkYAwmXvyvFnTykPWos
gauul+cmuOoFE9BFUE//3BTGbkul5/xl6fo1adPJL2MMfVPrnK82XnP/cc0zQ4Zp
TGcwQn0KB2hlQC3hmddPduHgxnvhM7m6tKp6tInSOMVdYFQ547h0DodctT0OGM7r
08c+KO7kF2q6CoIqKXVtO6Pxen3CCpEJPSyVx7jWp3+uNRnydu0PQm4WdGvMiHCG
8URnwYTevyYIibs9MzxZ3HbTxLhxhE2WvjsmHHhLWzBFcG4CpQHa1/rWSbu8Osum
sStmAZaBxpx1n5U/UtpvF5D2zdDPtgq7d4fYUK5PcmunRGJdSU7Wg6WgOIJ5g0D7
Rhtwec4gBVsLKZRPkiFUj3sLAIAA6cgGvUI0TL3swIp2RT/ci8nLXhPzGzCR1Pqj
wTnRdAoPUJSXkUNY5iarAoT3n0N7onsrKi6VX8Y2hVZ0j/OjhYB3Mkq84wCJ/exj
SMFA6e6ncG4qWkNGP/PWZISmEQKt++FeZLZbi+gKAkddI1cUV7D/G5+5mUh4SbFy
zrfqfY/IlUqVvYE8ZyvE9yoJzoWKQnoozIF7s0HQFYmjHeR7AY0eneXIhyBvHe5g
JCqMyVQE3ebQLjyOkZqi1tvR/MLywTlr+E9ntIJwt2gY6/BSvb0uNTYbNCujvHQ9
cV08cTU8mrfv86yUd42ml47/J8KgYjOdaBDh2By7POSewqt4PxmzG8HgK06zVlij
4Z76ZRG/asg1M93GHS9oOuvGXRhNCWlWgbbE/0nC3HLx4I+/Xqwo8c8/KI40ZdST
nZejRZg42UpWwFgd+Cc8MZV7Ifb1e90fZ8vNgmiMIdKrPBBBD3hYTCxWRej5K4O6
XvMLvEYMvEh1kRLXHcXWIAAQRXCFPMQdLX3JbEKLiEjkr7xnWLBwnKCDhxdza80r
bjhlMUpoUebjafJsPFvkNp0H4G28WI657wyTUid82dbHpFMi+CwhFznFhs+j8E/p
G6MhZ9RjoeIVuCXUrkEOqpLEkQhHJCgXCsG4XGwUT+8gLOe5PzU+zdFmo9fopb+C
YsJtwnHpzFJdTvskPyI4G/2gdCfpahtleGI/iuejOzxWgC+3DvHA5zz2fZ8zVB0d
4mkwouWc19Zl0ik3zYg+J7puyu4Z9kXtZXIb3SMRqiVWA7Q5RUZjmOjEqXbvlZ/A
yJ5RNJGCDcCvT+qA/nvnSnN7d/Gq7G0K1FglgTKhVHXuYvyeOdJ4UlDuefjnSwA6
`protect END_PROTECTED
