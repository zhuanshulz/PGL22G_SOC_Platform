`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LQNRWIxjW3+MHmLRcQCoV9HtbyV/idRVhV8ElTPuPVzCc36e9xspQdoyd1oCnwhv
5zky9IoVB6eVR3WouIHI3wrFk4NoYi2T9ODCn4uhCWh9KfwxzGbllyPLc+zZ0+vF
EI+BPvDMw2mWKJCUqYil3NpQny81kQbRqNlu+SUekLa7Z+2ZJOmH3E6DJZo8Fxw4
CVhQD7zwB+n+wa/LHZkY5q+sk3NQA93c//xadaKiIbiXFZbE91orV7x0BQXx/hLq
4cq1d9CJS+MSRpumGLlvgUzmxTnXxp8LliCMBrrCHydtA66Bd/xZlfMzl32FyFYl
sDvYyakfmhivEIoGFQ+hDgxz4gQ9Pb95n9QVpYYtajzKB6wvxbUI5tCJ9rW9Senj
SWMUMbuMQjjRGscHMy1JoU/fQbhi9FLn85EYu9C8OAHQSjGBLfGswSeK4W5z7pF5
BM+X9bISwJp7yqhqPBypsLnDvEW7IEJ2FJtRy33gLtYwS7kNAWv1id1KEEnyYHMm
oZi/e+DuqjTr7GC0gcN81iLoB/vIpdItE34pSMGMDc+0yQR6RbpZgS0Z2ffp6d1v
ofecqawEvCF4JnVcuz5F3XDtKlj8pKxF8cnAqAXN9ICuzTEXLBsoELcyWY1lzO+6
m8aFCAFzwnQZe9RFBtI+D1Cc1Q3qAFVfGC+NkWShwwmhuayFev/RPbxn3IPZL93X
tq0+isdCVx64t7hWzeLec0Vc2XYpDPqJFP4SWBfR+BE=
`protect END_PROTECTED
