`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OynwksZxLVDkLxM3rdMhUj8R2AJHiwbw/fD9fka6oJGHCR0r/92mWMCHvpM4WYVc
4yvZyc3ie983K94d1ua2j1tXU1KnFMgzNwCrIgJk5fAbKh5gOkT8BLB5frsUOJ1v
1VyCSP0CAW+QHarlBdAvRSgEMgqW5srtOW0M5BZDahf3o533nGmdQd4xzcSVIUYS
D7z5fGzxV/6RQKCpoeQu+9p9seQYFS4d6zB6TFkzzLVx3nVKJ1T2XU2kUa6Vl+Kr
f0eusfLO/OuhFxjw3GIZDsSZbxyCzrshCqGiLAtzB6M24VKbMkyyg9T/mSc4agiT
lz410TxFOt7xVnLy3q+wwyy8HRxM0lNUczGQlU+jzSHXeMYxrndaXEmTOzU4QWlx
W4RuzP7pToPj96PvnCH5ro3XZeJf4eiyTTxbvBqOMjS+LdKBXgPELZQY1QQgICmV
gLwa25A2r0ZTNmAobyuQ5OqpvHp9ps6xsmiyBl6JHdRMKt+Yn91zQ2nbl4KYKESd
rKn00u59HxYj0wJZie5aaO0jrtWw/4Xbf7xAHsl+8+Q=
`protect END_PROTECTED
