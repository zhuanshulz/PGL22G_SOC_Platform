`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Lf0kmkzssukM30qCxS9y59KyGZGUGwVLoGdXeEprPDKhbkhd9wHCl6/aKvsfogD/
AbgMI3AJauPkKM9svFdahIhjOQAQgMAOYChF36EDZv6olFWE1ATWlD89nCj6ziZl
S65alhs89r4v1YsG2Czi2ENj55n19TUzSnFz+KLIypQQun5bo2EYWCyStR8p2pH/
eIjmXwz0VPdqxSHvvX9z+0SRKnG+p67lwO61bvqNfvkUHv4k8TGNd1imuarhvYh8
b28iPjy1Q5uLqJx+JU/sIza59zP47erhiRQuBVqjUEiYZNqNzlLienyfd7BwHZ8E
0aMIS6zFmVQdE5zeSLn143ANm3VqV6xNDiSR+rjycfnoqkTOC0COstVRpTk4UdV6
OqqcJADZqiusrhutnWZqDiECKkLL4TDoLKUnRK1EnXEvVx9x8NCxm2LSCB8HYWXZ
mUZldbpwy5ubtnXTAhqF9vg/L80RM+NceaSxGgCErgEQqXFQe/x06avCRtzYEPD0
FkAJUab9bWOZYq79TFZf17wfRCWY8zL8qtViMQuS9My+wf9RYR9/sSgAwU6QBwaV
tBUoLZKC19ni7bSH5f+3R95NFBrNnn6Hj6hkrS6IwP0bwPwUFn5GjvvV9H5aHgbr
DkEqxBGgFsCQz+tkBTBdPK9dBX6wJ8Jl1Nu6cGx5D5O2cWuSlPwTCp2KOB+5Va6y
SjIQmTawWJYqMqpb3tcOa3gLWA/DeKgPbWXgYpGFsUN0sBPHsf3F5FEYRHX9nS+i
sS0QDhZn60JpP4aLRbZKn1WwWdkHbWuDYhi/xuCppcrrllWO8opWokx18UW5bkay
qN2PjXSKyB52d2jvbr473rP0Uv6+F+Ff+cqMMWZtZjg=
`protect END_PROTECTED
