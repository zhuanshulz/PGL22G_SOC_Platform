`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
npLW3RUlSPIRfH7fCrgn/WxGOo+/umq8waRKzAKjkg7VYh/m5Tx8ZltxZiYImXEN
kzj0rDlKaqmnu9oj8MCTnRNlDflGuRwuZJgcE7L9/ZlEE8ZocQ2UCmaxxYe8GMfP
rSsbbaY1mYMpjo61abik+LBQ9KfLBMJxDHUemZOLpNXonw9b1/JP20lWjCe2YtCW
B43rhDI93fIqEbFneXCTNp7igcasIXKZ9iIEXgXaZZljPG7fJwiQaLmMKaP6oy8V
lsIOD7QyGcKmmOPn1auEKPcym/kdec3l0WBjf+ZY9qSN6OuWGyRFt4DcDJPI7YQ/
x0oUOBaQL1YP/a+LQEp9Tg3rqpNfO+3IusfC9lWqgp+o8MlwJjwsythzt4Vgyu65
M/bLliac104NdOiTpQ6V6pPXOg/UhCOpUS7d1SUHdKQshWJ1YYrI9ecYyPFrk6q7
qjuhwJgESOzvMki+iw8dIps8/LRqBspNx0KS+6gzZzYVW3FA2yYUq9C+OhS0OrF3
`protect END_PROTECTED
