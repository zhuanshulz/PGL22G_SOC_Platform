`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3Cb/1s0CfgmGTrRVpkeDXuWHDg39xy/47yVosE82dNsUIZehUJxofwaM8WEdXrv/
VqqkiPlsSiBBk2WP+QLQX5KSDUAg34p1umbA2ipUub8JhoBqYRLvHrjjyU4Vweit
GjNiLV85DgaGM6jBwv72nb+/dwqxQUEF3uNCbBLQDby7Rpk2szZfPot47uSpenF/
gXMzTNkO5wgTS4EYRmAebgCXGmCxoB9MbgW4PXsscXfnTbX8VD/q3fx+WZ3wzKJk
k/R0Ya6GxcGAxDh5Nl5OpOhVO0HL4ElfxgUPe7jwtJVwf9ARUgkO+gkZYtqD83M0
+3gh/ZfQ0MOIYLzF0bKYBifJiCNRmJNtBuWPUxHAVcGZ+gwA3DAg+mfNu95Ry5yq
lgRx7oGYLHkUbuakG1J6Fwz7nv9xtlK1RE56hubxv3+N2HanOVVAvz37Olp/lTvx
8+I3W4UzKBZ3G+xxCj2185XgxzpB6XKtlLf85g1hAzR6Wp2qJ7/OosOCDSZaGJEv
4k/Dfnupry4nEmjRuNKCMMWDZu6Rm7g32vB4sb5gpbQUKBDJNTFDB1B9U83fsKxA
3S9Q/3bglvbDA7kFffs4+Ryyr3KLZ8U5HfDNM8n1LmSqiUmVwICLG2Xc7UMJJ9aL
3Dmj9+0hiI/CPfZISS55PXaG11fjcBdjgzvwnP4QkuMGC1b14UNh6ovq+kFmCy6A
asTARLzDzFIBp3rsML4iRg/tjN4FQuOi8g5jHtAMpmhU065w/GPLABT1hMriKGSe
imF6Q1/h8Fryr0uKKoBHJvgtm9qxsKIn2bp7uSjxSoMXhzl8AETs5KyeCc4r2LlQ
nuqI9y8s4cwrfPQISnlMGSjQ0347K/7TZ0+ahPVGQeZw5IQIj5UbVbskM+Wf7vSO
cw0V3DhOhsJpcrVseTqt0d/IxYVwtRFw6hecXdh058eDkeyfS3d5XQxEfqHbMw8d
RdwiH6w5eGLRu2sWtS6kscr05dfN+eY1cLFciCyo9C+He+zjuT0pThv8w5vwPR+C
c7VRHRVISu/uWX7OvZ2Adjx6wrBphWM3j0cHzxFapSO/rjYHvW50o2KjD7N2Iqa9
R3bL8Foucj9MJvjnuAL6ZdKgH1UgWk6EFp4fa10jKq4=
`protect END_PROTECTED
