`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qc5wvMVCg7eiZ5s5sUA7DYYS7GBqEy6OI2P705mV8DH73ZPQ67IOMW2eDDsEz585
mn+dGVt0XGkUXgnD/k17u75ztfrSMYudMfjMmFHnqBUAkooKLJfU/h3SkEkgY9CU
a1PdSrHxTcPzHEDDeE+TfxsNVbZ2uIi66pB2fPnz6KyAFQgvZGo4HBEIhZH7j9Ha
Z9n1E18wSJk+PWaf4DRQxHnN3sboT8v560ZlKQCPNRbBzyi2gtZNCgOYJBy1grzO
ImSunpNcmoZmypDaVDnmuW2wob7MsHquus99sZwrkEdHMAdidoqzslUf/nPrQ5y6
EtwlNTTOc4xs+8yzVyJ4BPpHb6EikVWoM40cxiVGSRY2HzWyM3Q0kcDLElRaVsg8
IuqdfXVGlPCjULC0C9b+QTsfGXDFDweeNKt0BqbWiGTsPHiZiv18yQvZ046oaoyz
/R1cX+80Px9LetKmfJQXYYeWGbmJu5KmTZvU4FkSPfMeCtE5dCIdNOzW4tU3FnYQ
RXy4waFnJ5GSQVtFf/QBaQIgb02ilLGYPMvhO9aYfGDnef2n2zazjvU9xJ6z1/NA
9wA90U19U4AkVaPeP0QlkDHe/x/NbvT+3mRA9AkSLlthlDNqOJyw75ZaUTNDNxlk
61Lu/7LAftkgJZi47wkUjhvZH/KRmPKa3eDd5fGa0OTgEgu9oFFV4XLHEn55m2RL
iQ78QhqnrJN85CkUz0LrSHFHZrZXQohuU+8cWOpBAc6Ffzq6dh7t9xi5NALCLHlo
HpR3AoZrDqv0/ivBMo6VmP8DXJT7KyFxG6ldMSD0Zt2yWIvtbi2u4H9GYSJ2zagR
j2VRt0eqbBAc+Bifbv54vudkAHocOW2KTU3XdE5x0Xo1BHpYbt/X3Usmg3XOo6ff
tbuPIuKXDNGrOgiz0dHGnFb249WVl87KxxFCrVbl02PFltYop1f++b9OcVVhnuDZ
MAwCBbaFkgnqqtV8xm/ZHsQYHLCE7N9EXiAznAkfs5rEpTccGymNze3xf6/YpzP+
wvEIp0Zf+IXnL3d1paTqtgO24XlP+dF5xHekY/ljqdA+d3KzJ7gCt98OLoUj2/iq
nk4734EWmzIIv4QWKdOyorFPX4HDNl3jHHh/g+0dudeE6brW6dXccRrzJGXQdDJR
lMtg1E8qF7kCUz0zSUTVFTg2ryya0wO3I7gtd5Y/AMyp5ymjp3DiwBw0w9jZ4f+Y
Y+hh+ShMx0KMFh+KHmKwxlwOPGnoKvw8NUIonfBcnfgBEXDpxVSyWcNCVxlIbtAl
M1mkyHlfnvGzFgANODrELHasl379K/JuriIexAA8j3OxjYmxfSO3+uY2LeCD2Eyo
IKix+PYopGQ/Wet/MIsk/qtUi0FcbS+jiesb+PsE+6r7bZLKsW6tRK3drQfWPCBe
hdISUCLQI+emmrpl2/dO3wGY1tsLvhTOK0U2jdjmfjWX3tw92YdxEQydp+pOxAWQ
RhTbHQ+3nNfy+qPxIqRnga9n4CtScGQH/z/K+Oo0wVsulgC106wVoLckQ7DHwEk+
kXiJKQuXV+dt68BMW0OUZio+RyrEvC77W7ysszidk73MS7bHR7lH7ZHlBKX7J71o
AmBgUFcFsOjOTxLn4Xxo5xbcHZpAnsWjRaacpz+yCD/5yA6ZE3dfeBxQxGxU4Nt/
YNEAyG0Cd4bhk6zuyukxGIuY4IBTkS3OtxGfk/U8U9yIMXGrb/2zsrQ5G4PzzZi5
UedUfqDcMmT1z/WLNJBH0JOPPfgHDLF96pF4skymE5wbqmcDDFpHHEscRvUAAkV4
XYkF3OFLvEyH3IuV7Yb8dk/4xAnqUpXDWCPzxs03sF1ez+I6onV8H3eamUHx0JzM
OPKghXFHzIBcSkQn+aIo3id9cxWDl91u4ktG9ECclQnJWjp4wjQJVnUxDbeMPYmR
G/wI9fzxl5Bjex9947sCBsTD7bxTBdenSLXS7T7yKXRysARNEUAQSDbVRv1C0f1D
UqP9hYbnSFBnQH+6ozmlJZJibJyBI0D3slKRpn/+jSYCGqoiGdoDzuGjBl7tY2oL
lveUPsUbBybze5/xfcl1nLgtFQEkIe57WNmnwQlcYDP73MphHCX1eLBRGmkc72A0
IuZ+i4LdmpBa83HriT4+4P68yptXoqVy1TzJLcxc1Ji4ycN99PrmSbVPIMkXADYc
70KD08sntiVbSzVLyjwG4n0XuyqtxWeFVZYv9Odl1R28CGcTKdWI5hwIbniZj3Ys
+ZvVUPe/Qp0NF/GrYmt3RLOmq2ce87nI11ZDv5SdbKjuzx5VjODmul9Lq2afOREB
IIdno3hVH/o9f9keXpX0QUORKP9MQ3nyonEafVEpLIOZJ4pQ4dCr4R/HhyKa7KwL
PFHpIorEEIZUGieAgtfoSp1Dw59E4f7ogScKbjb8g2lKSkXzAa8ml1yoGjMaBxWa
D6AixwRaxAF4DoMXbbO7REnIUBZKGvfSqK9jNE3FabU1M/PVvfexT3ybV3PY7iF6
N/Qohkn/J1miKcgkc2WF48rXC0IntyGdLkegshfMN/E6j5EO/RWxYVvdDRAMdtKN
/eLLkI1XXnnNnV6EPAbd+HJOpPLAMY0oQL3qMLzetuXUkN+JD+KkjXY7PYy8NmoA
t8IvJdedgg+t83Ss8gIwsRdrjHS9e9t144sa1uxlUlL4e2CLUMM9x7mztoHHewC8
FELQSpTXc60G5wIYVAm4lPeO+hResEgMR8eupfq+F/0kr5UJnFy+5KuTHxJaZkE6
60jUXnQ4VfOtoDnknKsliJnsnza+tGa4q548ltvJeebIYCJHuxmYwn/zAC7+MffE
7Pno7IrUhZ1HNbRmJjdPR6cQhq10KqKHKIONh9awJETKU8TN3bdTmUZCntQ3vaL2
YLaz688dUQ2UaOiLXyzOqkhKja6GA3Zb3ZzVDbkd6X5nCiwfn+bd12xWs7J1EgOw
2TIqpRZP6ar+zMozNbvc9Hvn2hIVMrspiPKdUKn29Y96JRSPf4V2eW/vUW9lkw7H
fB1NPHSCI0lg4I/QW+HHAZq8Yd4tCB4SowZb3XBpUyl63bpEe9oDyWmQ0Q1IRy9U
NmsER0nrf2t5EAQ6WsEYO4K8gW4/TzaHkstko/J8Af1VAKbGmx8r06Ry01d4GkEp
Ls8/WyftMabKPpUH8BA1sZxQqTwVcPMtRJb5HuADhdWQDJYlMEC2160BdDggY4SO
g0ggVHi6rPhH7S1M0AQzsfKdXhtjkd7IoEWW2xC2Qud0dJylNWK7VZhS7+To7uf7
iEZTmyZKSN7VsmQa6Xr0bvJGc0rQ92OHgXb/943jTwX4usDeze83OGsRKUtHftNH
5T6vjCPJs0iOk+zVX7ax5O+n5btfQU4AD2R+qwrDiDbQiBFx4SQKwzogHFwQjlAw
hWit2/pITYE1HtGFo78NZVrY1fvYUgzpTO/o8G07iohpEbFyZpucl30hdndhA5qW
6+Z8dLCvyp64telkFcFOooQ5tY2B0KX5qyAOR7WrM6Y1iQtKQsdY9nfBPnO4W4RW
tjbYohQyaQWcI5XZejnuyJyrR42gjoIoaF4pbhVyW+rNqr8QH+b3+DILLEac+PhJ
5n3g1aTJzg3TbTdi2+828LZVOXbBSt7/KTeBYjX6NfcxDOb08Zud3EGWygz+ZKdR
fxbAu4W713w4B7+PQG5nGO6OSReOYasHh9Bg7XwmfqC56Y6l4xqi6hwNFOGfPGi3
JJxQ9FXE4H1lLwDjT0JgTy1goufLQOvDw1X2uIOfKfkkvBoN+a3GniimbGxv4gug
SJvOeHrPUMMTKwm4poIRvlVQb9pDwwwVjpY1SJuo1/hsCIJt+dV57vzo2egArh/0
q9ttH3K8/sxKkN9Fxfy5fnLF+hwxXCzeLKzr0R9f4xZ8rJAdkWc4YxRhAnfNWzR+
DArcAQRhivRyIpw1tAQkKmttRkFhHSrOZ+N+R4YxAtJwnwCX64XJYO6Nidxuq24s
Ba4FCU44od6RGOHdJb1jqkZYJRpgSo9Ys1I2GhyFxdO+DT/Ct6dqR9r7L4AP17ft
5ob4YaCI/oQfxQAvXjU73fBJgoAfELnTveIUYFYurM0sMebp5a03WrB/csWG1usJ
uKYyqGL5BwXtV4HhFzrcSM3RB4OagbOaZ9Ed3SagsOhXmfiexY6eFAJuxI0RUBvY
cAa5VYkRQQYf6xLenFpy4aYelJF6ju7JORYl/np3pQnaDrT2bCEMVeZtmICvMnRH
613nHjEID8mGzvWmY+kvdAi4ONxHe+vTDY3SIV3G6ZMiuTGOui6tFpn1uav7buRD
GQKBAJJZRwVthhoi4+/9xY5VxHN1R045GYezFJ9zG1GTX002HBlQ0boU+BH2FuIA
dC+neup/WvsMKmZv3cGLAZEX9PVpsySNCTWCu25KZXnHsPcRFeY/2pgno+x8YWiW
m9TiKmppA3x77mhY7XcBWAXE5eVDc/z+WQV/sgd9ePOpNV1b5m5JEY781TM2OLUD
n3f7cj4Xqhl8XVYEzfzutHY3Wc6kOcNHFRldMEN7QVlZ7cR1NR3Dpwjc1eM/LNfp
kWLHNtBqF5zgUUDB3fkATEvPGHLUO8szkVbQvYHGe6Tz57hBPF3itWP7iCMuYvrl
2WLwYngQdhhYd4MyyzJ3sj97JpRpEii9u+lvhsSJFM+Zmszjz4SXWSpLEv7ZIq+K
t/KNHwOdccri/OfU9iy0m22yaBEIScADQDpvAM0qBMdl+PKyDZfoxM1L/XKjMCnv
j9+gUptPmej8ObjlKtF8Pj1RV7xYNUfSc1/45jFgGfNKP/aaQsfaf9MmianyzcIW
7IPg4ZsMdI/FN0io7OHS12rmO6kmDSXhJDl/G6Yfoq027btY36OJNmIP2oUEPHC+
SUUWg3NSV9MTNOjhzk9Ood++Uz2kZ2JVOck9lpvBz0oGGl0grnRJn+ct51EfkoVG
yYHszVdZzBebf0JXb1mL63t6NhNjSj2IiQqIIVKn4jJk8Niz0d42tetxYTFV2MKA
ICzsUZZ9sb5W+38eJBmpiFaQG1WEExtwrCXdysvX2YQ7rhskz7KiNHjGKMm8t7RF
3FEw+GALkMKsYFetdHeqSYCkhfcOTy7HtavBHAByO+UbW88cdK+1DkBv6vaNpNwK
8UAA/3E6umh5/0NYCFdyoLbU5SyyrSWHh32sQpgAWfm2oeQ1FhxlQdVa0MGvV3Zf
6AiMqgL9gnnHZduZoW4bZqjvmSpWOu5KKO1dj0NiUmFloLwKikfjJLrzHO2NElfJ
XlDDJszmu1/dPKeY1VZnBqBgGpSTHfoK17Zg610sRkxZq/5IbZXgghCf8TVRhfHr
ETzi+S6BORJl+1I4ulSZksSHzdhX9Jt34KNeExq/YI4G/NTMyOF+x7O5EhHHZ8xN
a9hDDiAgCQOJsnErIMFjM6Z72UJ9jWeYhBqk312YQP5vmCy2TiFc1jh97rVSxT5j
StF/O+zyzFPEb/JiqukdoRKJ9GwPloXP7Z17RqeNdWVaTIrPuAdDW1RKB8C+1Ig2
PmCrd0d635CxCD0+dQtLEqbHjfupjgv6n+nOa53oMBjbnd+Kd35XhJe0KCdcB9qv
Y8f6IN3X6bbfGEnjKet0+WR0u/yh8igVPIju/ihbbFR4kX5BKUWMhhgZyd7Itr6Y
Nm4P1ul4ZmyP7hsi7ETwIm9ZVOkO+M4Uvy4rI+oynQMganic/APEYDT7jRbES4Y2
5fx0GFt+p0oFBIUVsfHJo4gtpLuFD90xHVg6FiPYfIGHUQhSwNCmFoK2r+fgptuJ
7LW1gfjJLDbNiAh4CHWw0fRvHxj11Hde/Ki5ePHOKIAfc8tRC1rPAf6FeoxzZD/E
71TRpCGR9ZF+b2gyGvXwu7ocEbgUBou2DYHJFznWDA56yiIuRUSY+1cIi4KxrelJ
Ll8oLX1X07bhpITINVq9OKu7MNREZP/PkpJMnHufS9TXS6zBIEpQWDA3C9m/LQA1
2VDSyJdnrYY61FxwpDBye9TnEsD/4zvhLooFDTRU/z9Z5pv9glBNwXDRjVgZYMjn
pMTMizB0huFxI4EyeszXc0Sj7mNxi+/SnXO/KYj2VCIS3BkOwATaO7Oc6UNP7wJy
wkgR5oGvQPgRY4PpScQf2w3H6WuSyln9ljTKB+ri4EB1RG7s4Oq2UgPaFuQszMtO
F2Vcbd0E1WWX5+u4x5r+rCBnFoIKeMC1s58r1BSMbdNHR7Xi1jpFx86xeOGpIBYP
5fG9Wm2lGL5/2wo8QKOMuCYT3RKiIoNGPAHNsTGRBwWTeEBubP6sJJse98/orn6u
q9zGGpxUQXvkMvcYfdkoIf0euiv6ro+KkMDk39OCQ5Zsu0+K45A1euDUE8BQF6Wb
WE1PzLOD9NN0HeJW67w3S6hKxUfmolvvCSb/MYw8F1YB6ngjW6N60y9bVXa9/z42
6g6mk0iYGSq7MdEfvlUbp6cyxnujOytCZjkhL5E3J13gALghlzL0g+6IeJkTGugp
SvKU48Bk0rqr7D2eqp5pkQP9+tBST6m759zebycHd7WwhFrBp+mUcrVF+eeVBCsa
9up61C+fSYnzyhsyrkJV73pyl5HEIjHuUVgtSAtOalAHDe5jmf5OQmrTLIN/dWZZ
j2qdEq7IJOdhO/bAJyQCLQYGD8wNtEYfrA4KPRaYJ9n/KiTOf664poadoYwkS19W
g1cMSBkfGXPCyIGI775Yy/DVnf9hK9jmm4q3og/YRmvQrlhx+kojSjkSmfoojg3j
POHTQ/QJ8TXGwj6zP4ciyOjnynF/yQkLlzqmyZPnX+Ve5uea5mpcyZ65rdnu2NF8
cli9n+jszcQ1almLh2Porh/x5bPV6IIBdeClekrIZX1ZRxuBzOwfPjLVQ7PheW2t
Lb2zfoo5gBKOvYTnySOw8ZSJiY7/kANTJxQdnI23W91QN88gsoChILhSvKX/wbWp
uqtmydJPDqWmvDqpNKJvuytz5t/OZ6vg4vVxke9yt6KCoE7UB9EcaC+Pf1EBkgcl
Rrtp2CRh2XsrrAfl1/owtTk6FVMfIl1dYEa2Wg7Eakbh/mf6GGU0Z+jCtq7ly1Ov
Ln7YYPcDJjHK7fjV7HGm1rfEtq2p4GQ9+5qYnTlAGO452/qxl8VQDjbe+eT8aKuB
VCzeYint7mSOBvewHfu0xZzzwn7oLYPXA8lkj0YviUsie8N6iMmpw75M48sCuBoI
70dYs9i/hBwkLf0gw7Nl5wobz+BXdSfLnP428+Qlqr6ZPI/N5ZFY50ofOtlxrfPo
igNG1lno8Jrbk1dg26l6CSATO3PBMygyL1hQeRnJNGWlnhuBNgsW69iUTX4bCoxg
bWcE0XmTr+pmbUUCXnzG3J8qWrLJrdSl1ISRgoIBQsEWksfqJgvWaAiqWtuHpuqL
5Ut3QUe64s5cv2XF63swVCAD1RnPu9hg7PN0QAEF53M1UkO1Or832Es/wO+ELiYa
ZDNzzdkVizyaD68HJu2EK63kMch2PRsPPfCCz9oUMAKmngxXXbRSz8i7ZHXc/B1R
hFHOJJdofbri/gpr9TGl8TDZAenGuF7F4sy5g8dtgsrWksytDWQ5GNl6y7/7KU0w
UTDASWTk5aPfFkyOqNzVjkUKfU2O0ZvoajmtLiRkvEMA+abY5TnBfHcvbjolvYCA
YwtFANUeKcrs9lhsBvVGKNdyYD/AwPMDtICRyb7+Q4Pc8xH84GFwhmDV0jaKe8Xn
EQnnprYqG08a3QzFFAgdy50QWFlfqDgWx3Mx4DF0K5YLzSWjKP+JfE4OSo3178x8
y19oFaI4zD7+vvo9wHQOt+GjwWKbEm0dl7K3EIGR8gPKAAx+NA7tlFyU/DWtr136
RYtfGv2PBgS3B+BjIJCbMI+ry5hFVWX9zUAyVxxsCo9iQw6dshdURKhWWi6fn7jT
ozdDZZF/XuU+J5yysChHRi1Y6KABdzcVFUEDFrKQUNo5raHhPyjrESJscNrL/crW
WMzxl8x7UM2A1dJf6wLqmyL+YC8cGjNqyfsNh+O/+HJdUThnVRwqIYu2mcErqU6S
H0D3gsqQuYK6vbdzEp8bCPGiCoyDj7cQfx8/3FejXCkTjwq73w//5GjFdejespMo
dJWsB5GK7KfmEV1bkqbsOHXaqb64yIjcQyG56qhcvayDuA/8D4uSnok2ANXhWEAd
xZLvZVDdX+nAXX9FcndOXEQCCv2rZ9/rxbycbKmznUDB0UU8BpDlxOyT4MI9hywZ
GdCYFXTWtIWWWzRp2mwnU16iAy3rcqWp9onIG+NVzF2TeZS1MbQGqNGH2U++WUOH
eabJaG2qDG+R7YId4+eHuHSTA/iVcclCuXxJg1KbSogb3Hmm12MhJtEkV8moYWRH
8EJnXB4h/LxYCS4JBd82alr7uJBtOmdNeysuMyLENBPykLmywSzcaXLthQoVSeN+
RJULX50RKhM/E1DbstBZKG3SpcpscckPE44MaQPj4myxp+JszJ2jEBqQis+P6sHn
SaDV6DUn1w/vBzx7X3A/Y4PvKlYZx5e8p2BtjWt5AJAOA0yMviOj4YaEvQpToHU7
p2hjUrJW6sUcKPcV8lwhoPZ0bAdSbwWdZZq6W8OKktgj506GSZZITzsghdAfAhOo
ptcB4qVLhlbA673x79CWBJufzJFKYHSQEH2bylzJEclgonceOpwTsNcwaX/BUeem
nSdPkNdtGrI712CoFBeLNfSJa8lTmbzPvRsxrahSHONffiep05nOhT+EsnPt9T6l
c8ttLhiEGdwieclKe3V8z6HpduzSa0U9qFrYAp1YTpQ3s7h2J9pTygpw/cefJM2x
stAIbMDinRticSRonC58WevLevfSXOMSG5vqom0teko=
`protect END_PROTECTED
