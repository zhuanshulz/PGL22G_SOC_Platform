`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aX3yeZXoS6wvXjroqtFGjpGwUWRHIaDziVtqNuWSTEcNva/7e0vMQRPMGkaZwLs9
MENt+HR12HMdxXn3GYXmbSPtM6Yjbbf6ArrF0bQb5NjN0WjHfRhv+hGirKVrP6DY
ORKviMcn5o4rYso2HkL1DBykDitN++M8qHMmPg75CJTOJ7lv791Poj95rOY9x8K0
SAzMqqn9g5DVsTuAHhEjLoD/CXa1rOW6aOBEJQalYKD7aMDSoSUIiuuBU2Zn2JgS
pux8XUjpbBFz/A000gUq3fUCYVPDNaZUevVKCAiy7RSwjCsEQ0asmwETJnndz1KE
6W87/7S4yakwTseqgItgjzqdVZ45m5ysgcpF5N7kCmJUHZKLQVr4qjY7smOyUVg7
pVzkXfio01Ah5HSXQOwMRZ9pkp5qjsj9juMIoZqAYiFbdblCp+XiRbJoJOPMC55I
uoktOD4a9Rx7/lsGvi6GPQ==
`protect END_PROTECTED
