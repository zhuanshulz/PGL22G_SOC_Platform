`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FZ3XIzVqS00kc7S0VRXmREnv79z6L3kkFqG/3agHUARBmM8aG38sx1Ebnb1ICUNe
PeC/yTGxk5AdOfTroRFkBl1KuNdjlT1UyH4jXdkgObl2DtK1iU4xYKicklMhmNgG
a2rc7ccmkY2aXpSn0YUWEGXtScHJ2AyC6oVOkjHWrbTaRaOEuF9El+A5YpRIu9io
6zmuCLHf/EALfirsAw2sN/y5iuFP1wiAihFdTHmJOU7f0XY55Xxz2+qsF9NhOEuu
Qz0H2zyIo7IL/DP1TA8a8QR+8BBTUSb6pt2m3olSQYYcl2vlf7HOpe5l/EkWQjel
8gU7EX1/xhiPHDrKZEepaBZlPzHL+sbfjnUaZyDHr13k4E2ojIdvfTCfAAr7TApF
w7vMw3ThsVpCW5UcgoQQs0ldQq5yrAgh3CLhQEGv6rVXvJeLb2JCHFoX8+Ssz8x/
iqgPKPxS2i3JGHY48xxPXImn9UCVHj4WO47F8PXDHG5WMYztR4tnEdeyedRSTUPm
IxhZXfFaDi43XZecUd1oMRO1acOG8k0goYA4CT+AXUcLzOJ6/AQwurKYEcxacN2y
SiavpbcEelhyA80o/GCRJL0cP6nE/Eatbc5ynaBi9pxD6xZiRafek/uAPmYh0Ar5
7u2WClCB0jIxzV5zAqHx0O2bAzm6H7bj+X0R4glJ4rmmU3rfUZ5IVcBv8b2nEcsp
Xsft6DuB3quYPkTqWazUTPaVvLQcV8k6OvOXvmKA+FPi3taOx1hZsbQZ+cpHfkZB
HGih3/TbG/KPUC7djPZgfTTi/BWwziH6KuPcIn9IeLTkDz8N/C/h3yjlL4gVCHFN
SmoiUV6IUC+g6KOsDv5sG2N8dDiCHbtuzC3yC2YsU35wY8Ubw+d6ly6dw48xFA9D
OccpDWcHlHIzs7GTio83thmpS2Dd8416BcNrXBZ7zDe9UrZTp+iJqX9FXaOj6Gcb
w5GpBL/+HOxMFKQI0Flc3hD8Gq4JFUOjfNDJZ1xEBX90EJ0Qr5w+rHzBznW/DYRa
i4fzJHyiDO+nzq9Xr6xBrxDKtjmIWg7W7JZX5L8vOGgRu142bED2dI7GmWMHmwli
VKl87IvPiAjeVyW6HR5D3pRydiM6dvLML5qz/nRT1E9MiR0+KUcxdmt7J/ohHrVF
/lyOJY3X0ERnmxlffVBPOI6+RKMJUzwnCMM/ua9am+Ph3J+N0bZTIxIghRpafJRG
mV5xwCEq1Tg5YJGRpYMQ4Z8afjLvAoeWDprxbZjWfeiwD+VT1DEJWNy/x4ubsjTI
pvHK/4klNbT1DBNLdKJgdDY7G1w6N4L+mwP4Kh2D2iamjVRgl42uBffzZLLEBbYS
jUWjLk6vLehPjy6soPhaUa81omH4pF3tQ3MBThjDBdApFDyTEvgjbowAWO4XJTl5
1KviNXdUv8Lhrjo9MKKkXhi68QOWFPZn/jc2pP4l4GtlawzmkKkD9UqQlyZa7FDJ
mdS1S6QXn/U+C9fXKuTPo1dkRdo+HIZDvHRuXTXDEYaP0+Ev4NfnIx1P9sFDhO4d
+OMrqKt2Wa8vsYLggoilvYuUF0d2wCiPxO88sPwnpAEu6bNgpZyUbWOmKf/ZSxfP
Ig0jL14t+tu99ZzfBpaRC2952Fqw/gc5hQ5xsVybM9xx0YQAGrJMo7hQDVtLR+3a
bkWwe7OQ0uf1L8KU8KtgUZaC4QaKQ6YE40c71Xjtusz92SjJtiO7OqFSrRqoPfE8
F6rnHXFVWKp0acyMpMvzorpwfSKM5H9aETF4RxYJFQKzQrNAL9hEFSKH1RpL46O3
9GmGudzT8d10xmifJmGjdlPTQwZ3FoSLDrzbPKy9/8A04iPLCThi8NT8lfRQQlK4
n2GdjHVD71Jzni4E+xNfjKCDHMrcqo9qrn8aZI7bSjpmFrAcZouIom8w3RSCUjm8
fl82GJBpb3wu9AwTQMx+GF/a2dJUcJiIZg4Pfp6i3s+LgIUteuuAo0p1YB6fa/+8
9saURxlQSyS9WVrQBcO6NlPyy0pL6tZs4imOG6rfqGvixQeDsfHuJPih+8OinkRs
MyWnSFEXcWcD8x39eFGce1mZIK9vgk0ty3XWtQK18n8+lDAyZXjAh1U9i5lw7ouj
nFgNIwS/M2KwaqUIIqbqhUzCz+mrJDkMpeHZGVfQNaqy6pNFoy5QCe8KWgdPFjV2
cYirK4ToTrslO/LmoQSVb8Jqz8/dbN7/lC8GRRGYV8rsZYuXiHNfQGZ2VqsS4bH5
OWO05znPQ98iOO0JWYPVWrVZbEZOGstmFc13gfk+LIfw4049eKXioiuBl2WNxSs7
QeUwzo/0HHq3TTR3dJuyqFlvqUVbDgq1odaJhejThjEliUNJXLpQVK0N+xNMsMwB
K+czW3ZNY2tBssBtXSU2AJUX2RuT7rPq8VZdW/iVeHp6gwdvDZGTlqWjzXWQWhTW
X4Wuy2L8Py1PbukS4K6Yyl8cfjL3U6Gfd3xx5wXWjZgellOwa2Km52WnlK6/Fo74
rsQi7iv8+otiEzrth+eOI7RATLuTKc4WPDabEiVrRtgaAeBzgwDSdvpqaRY/EblK
uhOGvspT4IxtecG0VBujHbnovGqNhm0dW76W3AJu4m3bPUX6+pEieWR3kdhIWE2L
w0GpA57nICyty3gJkmLveHPJ7RouAR17JcjbfBM6Y3B4y3g1Pp+2OMGd560cO7Uc
VQ6wAhbQtq5eWcVtEwtROlaDpAuHQ7bQIFFVdOdoHR0xDyJJBygvrYWENZReihx+
oHXjg1u57sy+LiongWwIx26sFfr96Fqom8DdulE0+jbHQ4lPo2152gLecKQE4cKf
PNrwmRzjKBKFwejjZlqMT+mLzZG/vQcr5LE9saAR5KFpYDyYOJYQz16uL3YQb4KC
EpNrTeOjgny8wJ9kRLucb0Qb/LA2sQK1/VUlS/78vVjoIYLU1CCH7ILHd/OqRub9
IKsJFgZmaa0Q2ilnGtEJ+e2edxREYtRS9vT/+XG/W5XkNTv2McN0U741bn8fVEqm
BKMd2scagjbtIM2Gg2na329JFqBFrL6yeOzS0Ad0hLNnZ65v4+SrcyVdjRluIOsI
jUV+rQPxXVZh2yjuPPBd3jTIGjax2Zu0B5Z7a1043bPI9kBxGh2uXyoEYVbbWnnS
dGhJY8l8Ly5xzh0ws7uD2FLT0cPramNdzARihDSxBKsNo0U2/4yl2Zg6NG9cAy1s
rx5CHXIDYMddLthjJYqD5LDSp+6p1PPJoNxrma1Gbsqs35WZm5ne6q19iLv5hlSi
fu4XW20lv/vuf8SHxNtUgTAiQ+5CWdOmZhZE7xiywHDNoZieF1urIBxT/2Vk1CMH
`protect END_PROTECTED
