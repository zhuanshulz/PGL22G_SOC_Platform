`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ftvku/N6djzyH334+0X958sm2o6n82itOLK0sCydI+b1AcEQin1ZkrtfbR7X0nXs
5Ynrr71G9EbTtaDAu1aobUckTHcuesWIk7le68yTVIfoe9jXpRrFz61kZ+Fmg+O8
OcZLy0X7sEdil+KA07HqCRXdQrVn+GUNYBidfPZ8EiHhUMtXiTL/qvPmKKhmyrBW
ATIESwX3KXptUYHyT/slf2r1cB/5EHLBwr/gcAGjslPPozF+kW7bsvDu04TNOw4i
fmXycVAtNX1BQwXkQ/lbnVG+msFEA/RWCPdQmGQWs3OyLEwL28klnnZ4+DqC7WR1
qr0uLQvuny2dI0DHCP0v7cPaS/riEXfC+9PARbHfehy67tc+wtuxIKGTQq8q9H89
eSlwSeVvi/mph8inEiM+TsSXGZS9NFWn/DlbP0x/ae3+OItIQXc5VjsBT8l2l8ga
E+vVTB6AO+hPOkPuMYXlPqCvplXQifY4ArBKpT3jjjbsF/d1wxzslFIThvfott7Y
W67IROBUqGkRPY5uRDF8I80lSSRtx1ftOBdgvDiBNRB+/Ok2ui2kA3v5P8LLJV1N
PT/nfEktmk9iywjvK4abYwZJfORTGCugFxvAKZ3nF/VdldNvjG9GfkhQ6uMWwjBY
Q3wAab8JxuwMta+NAAjXtvrmECu47cc39xcyWtObpf3J0e0xMRIN160K1QdJgIMy
t6jtWF92y9KBmHYDpYgXe9tw2AwhJkrm37ZdkhVz6ZfQogZYA97D9sAo2wzFC8a0
t+3IzVfx8yMC0b9fRFC9C/1ztGx+nVrsIhaCAUNfGFVpFCw7eSadnHVyzkyZKLmq
6UVKhYk243E5g3ijmw0QSOmbeOHFr4RZ9HDbMXqto6k=
`protect END_PROTECTED
