`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w6SPkKVFtGG904FxQ+t2qQJEQlGUoh6f+vvbHi0Gzhq/nF5ihW3hWcrolY3IZ4YY
mPOveS/fP6sva0v2xUMxFdw8tw1MWizXkg2PpihkTlSkwM8FfJWjt0iv5WSnYU0w
344yUSVtd2STNXj7zpAoS3lGqxFGRWoFGCDJdI6s7pCTpBCF8/TVPY6U9XoKlakE
OCwkMiEBXoXJQX2r2gHU+cMbHfoDLForhKf6gABYFfs1YKw2VhhpD/RgSA1i5wX7
qFMGmyLBQ55R1ae0BX4mtK8YMcFI6I1Yx8l3jaIVwIgDKaoHWmXQ3jG1ckNyF/Nj
Bd1p/ImUFDGtU13s7y4EBO4ryq2RfcFLxzBMV9JLUqdlgYH7Lw9SSXKZK/YP9Qro
pu6K323emD6Ds2otxZn2OH2UUxbRSkfOGaOAUSXVta7EDVhZ87TYMQ29vPciVeJj
1pV5XHHjXLrdr8hAk3qGO1beMG8vu7GJLuq41I/tkf3jyaa3UxCN93KoA2gQEUvc
vhgx5+5IUDXPSqC2XUTJrI8qxQ80Ixq3agKScKnkkhZMuBE8GxkBDUKYdKp48XBo
j52RBtFwYeSQKxuV/H4L5xpgBu1GDUD2xQFosGtHpIvLV9kOXZH4Tzb204hlaDRN
8cSoruZmgo3M+H1+9log5G1Qx3irdWzmp+SDQG91FmFn8fIaeEDCvZJeN8uO/M3V
iC5z9RK/jq3aik6Elr+CA5OC0PBy62SfvJQAIvDXTmKuESDCT7eZnuPq2SabfG3D
BCkRT23CZe4ZD4BVwlEKXkN+k+2QZagKrS0YNo62j5h2l+O8og1yGjOPToTxmh1W
3h7eT2h773YE7SDXNDBcUXYSTrtpxsvi4ecgR0uPQ7uxn2LOdxRMvypLtVxGh9kH
sBKkFWsuM9GRvPGmaIsdS0ZeF5UVJJ/qupOJaWDqNjy5bc3Arq7iHX4Dm3O2BoVR
pHiP/1I+qDH+TtSYsK/PNAax2IqKr8S+hQzBfcjFlfyXrI5FS6pdP1OX/7ZbnyKJ
ldnqAwCK89n78xHffhWdf9VUfGW2ASo+M31xfhWMG79oS7KOxBfMtfvWNSpyy7ZS
A0YN1BumkDDbStN2v45GXZEt6/CiTgUfzcvLD4X7h6ZSnw0f3GxjDWPuYgxQb42X
KahPsF98XHZnfMBzXUype7sE4g+9wO7QqFEVXJqRjS/hSMSRy4aMWHdmLfH+yvZ7
thSby114h3Bq7+zcqwtiTWJYbmYiq/vpOqeNBnAqHDb9lclwTDJBQY1N4SqD71k0
/jcruiZbmc4qo4xOlQ1J/w==
`protect END_PROTECTED
