`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EE6oCuHWMmz/R5Tljjdn44FO2x9R0GSTtSsSSKoHdeZmxRT321Sz96K6fdh5q1Nd
YgEvH66UMyalnZNsXyIlz8osAc1/vjdFPNNU/XM1yGMlQPovtDNl0T+Ddc87u3UR
B78j2Lb1eZu3+PMvOBaf8ev8FGTFfmtRqs5ixBPZlZAhwljxBqufSGup/EaOL7fI
1ed0qAP2zEPqrj02rA6Qs8m0Bosi2YzPkwREywLyuQ4of0INhxTD/Oon1K0xFLwT
VlxU2Fp/XBgY5kNqLYIlHbNWJ7YPGFnPwi7EOBlsAs6ZAB7vIbKO7yLfp9j1c6CG
D1mgTEdie2Fv+S3s2xVEImQ7LQbS5LsgooNW5h2u3JWiAydHxqELAjy1JclXM6NT
nezt028UMWVoI7GqO3LuQHToT8qvqv3Rmhn0sfVD4bdVfSudPJzM/OX+QckDpGNG
4R16bUqUqSkK2XaIbMVdCBbiCln2NMO77Uo2e7vccyx3hFAWUrc3tzGIdy71xsPt
QJVbc/N41PfZ19CtUG217X0gOuq54JcQri9jNWJA0L40o9vjeo09g5z2tRf4HMvd
QOHwnVyK7auGNuu7k4gUXEafcXMYv1y8PvTyYgVlT2F0Dp2XpZhPWUXJdTHa0urd
TfXfXoQXWt3p4li2W+rF9GTO+FVc51Qx+ynks7Cwnsex7tc4WXDJL/Kn9UsuAIc3
4Vl1y2Bie7CdwCJdOSMxH64H5cOFdRlNItJszNrJKOdO/Wz3mor3OzuTcYiv7xNV
5CGYpdNDCAMQeUzHgLlCWHjkirxNZ48r4FDBXYvLWzI16bkFlwNqWzOpm48dsEZD
`protect END_PROTECTED
