`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vNiY7CBxe30h7Gt8iLSsGUGAWqHmCiclNlh8aUxQZm2kyiToGiY3pzYRZwMRohGx
wMByUlz3knTi73HDB2sV32AQ3SnF21bYZfyjLWboXFRNC76SaswXcGlGw66LT+6m
kPFlHWrnczU3x1p3E6MVbdKQ9tMDmjjDGr+keMp/or5MvFq/k0XapM3xRJYKJrv2
pqcOCP44YKhCKMRyumaJCJoxyGWCeTzl4wFbcAtmlbeCdFGUkQZX0aEikdR9Uxwp
aCykGuPu7CC+TFbYCccmWwtXpuyD2RyZALUMeF5DwkXD6i+unm+CTUda9CrI9UpI
NNEIJ9rzAZbI6b4a6MpfeFVG9Ik/Am8KoTiGfIbUq+sOMp+SeGavg30Hp8Y0ZPcT
go+TJgldsmbD1q9iO6BLPHorNI30IZZV4QIVlnjwytGlBq0Zk6YfyWEgny6jxf3l
4pPz+WlzwhA/IvRFBL1zcVBw9VwSDvWU1ChMOJoj9D+Jcj0S0PgWn0/MkbHnagpa
CRU2n62tnfYy9eQGyZolr0xNaBo7S3czpsfPsvaNcrRLyV8vCHQRTZaGfHoJZOaZ
GVIwQc7WE/BBRZs8wHmAH++/29f0aB7hosbQ1lxtu9PjIlhZST6t01PMtcLOsguA
Uu3p0Azl7ArtGuRAZMdzczQRB7l1OS2ckExyHcSmkDQN0RHehlBMOHFG6C2HFM4c
w59P13aLzR3u443tnQ3Ybz+3hTzR+Cn+4JkFOXcw54mjGGlMPPaiLi8vDcDwAehY
80/nYBfBGATb3LGWwx79Pb/yojja9k3PcPzDfTOm0J6FoqWx2qPLFX9Tt8CM4/Zg
FC9/uqtqYsBI9rX2gyIKtKQohrEy1Nm/+hSOBHRztSwocvuGbrDlIoQE5WbK15L/
ICOQmnPHV8vp/MHQqKtuSCnoPO8UyVX5iZxcTjDti3Unzbv5GDnb0Xd681XpFjFA
6fCjpN+oONk37W4ciFu01VZIN8h8NkTFfTOm3bkFDNPA28uR4j34/URSBJj2g34i
X63ZD+Nfw8DAOGJDBVgbzwjYZKVmXriFo5JMDwdYeSqLY2YHI//HyqreKzfYbJY9
JPJTy5pbpn2ZkmZEos9Zlb/wddcVfm4WgAuOXq5MJf+V+HL1Q1vFkg1IpDkO01Oh
/4EPKu5ARQFL1hPjnJIhuZ26KbqxupPTAzEQibKBhE7qs2zoFvdngT1P+17Z6AP2
szZ3xhtfTwkKJndCfxAJ5yZFycF/IagdCB4dP49N6OgiMVYz0dlxwu748wjBlddz
JKK47avzOOoZWcAWUFdQIhemHSiNDeagbI6C0Zl1tTL0iWaAni9WLgl/S/hCuLjK
JfS/hcf7h/aJmyKTtV5Re55guE525rbmrj61q/hyioc=
`protect END_PROTECTED
