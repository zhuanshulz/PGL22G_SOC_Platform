`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jepqCNF2oP+0e0bEj9kMnBFQ+SqwllIjkCX97I54TnJCELedp9wA0PIO/FejYBRQ
scucR2/x+Qy5RIsJGHaOqok+zc7V1sci8PSBG53z4FPsWosqJFWqkStxObWUTgM+
a06nbiOzpQHYthR9W4khm1inIrJ7FvzYUpXMOwdDdtKhruH0xriab84JMqEisTx3
KEn0cMcD91kUhY3AqCjyiz5ELigq4VwjfpYYx12JiqdkedKBZgapQaZT2pIOHpp6
+gQlPO8fgOTA9Igt0/NdiF1I2S6ik9iv3KPAiZoSeA7B/Bt50topdQUW5V2fBi7F
43ZSrfRsBuu+TYkrSYhN7cEbpU7cAYvonN25pgcy/t0RzTE0zNm+qGlYRn1R1+t8
JSA76nZO7CsQqSZxv0pRKILXw78ANAjOQ+ueGA7Lmw4ia4AdBzAc5vXveLi5pEp7
PurFGOrIjlYstAZBeSK+dVSyYLBJMCFvBoxb6vKVInI+UwTdb8pgrNkWXPj9YnkC
iqgaAVwwR02gibXOvf3YqSwBqrUoiM6u2LMSINgpBQFb83CpjUWJ6BB4xWr8tB6J
hlGsy49RBVPF10657JBnHMVveNKluKwXFki1KhET9x9ZN0t/WG2XVcp1C4fLvzWz
EIpozxv/SL+eEgzcqQPUq/6ESJCmIOsmvKD7vS1uX/I=
`protect END_PROTECTED
