`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6C4quiW67tLf47N8NqxeZbfOS1QUisiK8RuEoO4Z3dS/wuthidgkF/ewdCHAZz+9
ore+rEwkPISul6emGkdAqvKPKRqU3URc0MLYJXOB0kDXdhF7Oxum8ffYJ73kvM6Q
WUM8UNGvsCTf0Nl3Y4EMDG7vlSSkoHx9nus+HO9hlaXnL4kEeW//DvnKk0GtQ0F6
EEBkYFHbugL3b/6eczFJ6gniSJbf34nzyRyhvUF609MBNA6ryzr/fzS7pn5GKQwA
x3D0g41bYyqdxJhb+ET0OepoBMuQBMr1txZQ9Cr2cd2OK+2fpuRvYA3i/ZaMDxSP
E1PJSnFTbyoJD8DpejypM0U2zXB4Trtrkz7ItJajpM3TNw3VBAuxeyHjBHg09G+Q
6jFpJ/rzRKJIlGRQ+Tmq8fwJc56TZ/MNxCK0bszb5P2hSwY3VTyJ20bOA+FROPRQ
`protect END_PROTECTED
