`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0pf2+Lk5GbVF/w9LfzKoZ0EMcnnHVq+F2z3I4gy+PTmHoUJVz8OtGI9HaumGqL4W
9GYJlQnjwXCIyK96c22AcCG26z6u4R/QVMv5N7VC3ka3dPUEiOb9YPLEQ46ouU0n
6NCqf1Xef98oWyQ8WwP8j+hQeD9+jm1wU2T6hH0tzIP4VwyECDhP2ZnkV8lhw757
oy1esMibMbqFFzS/oODngGdbKgkYVRObSmkEl1alYngK9IMbcDYhD1Y+zaBCt0tc
8MADRo5MVsJ18jCUQ/xrmZ2urALJH759wiiIkkjO5+SiOsi3p71hpnPqrRDJxw2C
nx5mvMJcYa/qDT2HzXK6xesQ7LeDsgkIpylhuPmEU92q85RwbKkrurpe51in0pJA
kM8plVhe9Yb2Ha1sNJ/y3fjgWkUcSlKoiSE48ZvVGofBywWIHVbNwst0BUdd3zhZ
M+cnVInkOzjcUhoSUiQAm4RtHmHmOfvIQQLk3ufoUydHRdgrPD/rUm1HFZmvZfTn
1E42Mj36aoRPcrDxS/dvBHMXS/1yt7Co3yKQmWvjVWtPlVs00Gr0NpchWBjmFJOo
+l42eIfOCeKU/hwA5StIL0dRNQzz27EFM79MpcKNGzuILuP5z0QXhBJfyoQDAgXv
1I78GSecn4J0FATg96yO+2XGEBr0/22bN4FnRcqAZFHWt88WqcCeiamY5gbrK/A8
gY3lu+NkDsGuggEedQhfzKME29SWmDPMixBcFjOTgtAMGNGoPeADaPNmm2MoKev9
WpiQDdOkK8zRcfBBsRCBD1hI2FlCMK/EnIyce3xv2t8w8+GYBNm6u8e9lY2DeH1i
aY0kqevROFYZqc82zx/VNETfx5q2vxgN84Jhqd89dzhJEwqKkYO2UnSkBLCUgJ0d
P4NwN0SwAb9wYNBqWUxQqJpzOONthfvmdT3ZjAkWM56JxSTC+MQmR/XFgE27whcU
goAbOKDwAowEfhLrbPH+cVnJTFLToZdLZ7I0gwERCE3VLyDefuLlShyOOMnlgSdA
tbwT8yhKyUOJfZ3Lyanr5xcomzHiZHwoCHDxsZL8ih2A9Q11V8zz1fezIaiiX/qa
fasr9wNmbCHCHOvMX9R1hJsGFlOeCPSTtuhVdUJNUIu32SdyG3Rk3MS5cIFR1MN7
zXn5nB6BJpKty/yr4Npk0KVaGJwlkIgceVPU9pEJR2RxnD/ftKh2ZN62hJv+GOEe
Zx0SGm/68md22Y5EPfccx1tb8SO4nRzkIBEI3cJbIJVChfW74cc6/IAx5K/5HG3D
gxVtmE1ePl6bUH0yTGm9meyrVk2UBCHBKdsMBdsi+GqbUKiBhYpUPqI2PjxjA4wG
wMVzOVr2m0doDO1DiV2xxwYi0WtEzD0wmg88SmFqmDjoDprQmrImzy9/3bFJ9kGa
lH9pDy29QTExN2WhhLEvWJx9IC9hYRP/q9Cq45zTSPrtGShc0n219vxDHinKQxgP
HYb29tcqXYD9zR2KUGMkCdXUG1wH0gpV8bSMTMvxd83kYKjJYTmYcyz5kj1aqx6z
sigFyd94rMRlXdnZC92alh97OmIKwcj3i8C46/I5apSQ1jkTVltFBz4kDz9qVoc7
gRFyE7lhKXaoGA0kl9r1US5DcO4iCOp1rYg8RoBKm6FJB2DINksJ5xMdV/N7yLW3
zviLlUiOpj2WtI/3j5WjKDOvYbw7aXHhH8yXwtz1t5IBNN2dMcmA32YoJ3WbDXZy
1CbIzfjZ5SHpBwxtP9OvV4WXo5y1B7fbX++egJ3WrOYoCLQ48gU086uOhNOGcGsu
ha9BOBnI3JxEE+R7iKwIMqaEneSdDeEHH9M7o31iYuT1iuwhsqbsPnwQbJqt1yuL
wxvzbMC7EZ5tkcSuQiyy6J4Nnidg7irFho6hLIC4bq461/wmfJNrbbzhdg+aOpLZ
+5SWXmjFEWFAAB4qxzUdSpiwZnZmjx7zGV9ON96MTBI056uqDlNLmYKCA+4QLOpB
q0mih6GPHyTJT2bk1qSgVgZW6aYqCQf+xrqUZlyv8H9vjGPYt6bhdunEumUfJcUd
VkWTL8z9xAwic3GtpMFmTejaLDQS9YFFoBhb/Cm8uFbAhMX54AG2/iPQN7++SQgd
M6O/9VBMgSUiAzOgWgcXiITB8SICTvuQJPz/P205ppvkhNVlCEbegjbHMMnHbiG8
mQtSm/DOqCLOX58528fO6U0MBgpVhQ91VBSVAktdHGrrabjT3Qy7NBjTO/SC3IZi
/3LeEOa9Y629m31qwv9dVW7y/zwJjpeBShKUo6xY4F66vRGXX5N78h/1mlSVH4ez
kHNYaG2fQAAquzDp2cm44TbAN8nt2QLYIpgStiaYetjYDWeFYyOOogBXa96G7bg2
y+wESNV5ho7SQJqGYxKSk2m3kwCSp9Zlnpn2hFg9x7w=
`protect END_PROTECTED
