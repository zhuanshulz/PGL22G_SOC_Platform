`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K3VeinN9b+Q8AjsPy7HT3DBWthL73uQOC1ZVaEmvblds7K4xF22emnPYWLt7LCJJ
xPBhE3oXDT6KvPSMj3JbnzCOySlojj8TzXbjP2JMm1Pth1W5SSRT5fMS+QzhM2fg
2BXFwRGQQmuWmTY/Wj5NQnwOadUjRy1X96Xp9zalom9IWjBaILH/RipM+MspuYZO
MZj1KbF0+NBFIvyw2u0aykWEr+U6NWlhzAtB4WiEGIeiUKKUNF3BJXjaiK3t0XPs
r/hRczoFjjdsFEBUjdfr1sFwTF9F7RWhfEej71SyX6ZBVCASlueDE1kyLW38yz3n
AgkK0o3Q2ZvSBJdtazbjG4hfmIo3Tnc0J7UM0+si9J9a+ml4HoNmzvVdkcWHwxUb
2SI+SjF/CjXdG55YmMI3O+NKJ5JGCE3WeOOijU9qESFkBdxZz/f6faKggF8ykUdy
pL/mHttgZppgCZS+JlmuzgP925DmTGTri6un1mreUMZKHuqDraNMgf0f9+Htn2++
cXScXWxilnWv75jfRpn8gEJhOEUyDps0MEWUP8rhra/EJlmtmhIbn/Ez51Vh4V+p
DAfLuknC8+pZ6/haO9gw7B0SvWXSXkTEMooP83unV1bw1YneWEFuVmoyyVaGdgNK
CdenHJK06cEPilR04e95M0OClwxBQjZxI1qQFpW8rzeuN9eBFwaROUgd0iyI/wmd
GvJX4nfcAc+cYW4wRaAIbxW0FpW3euYIZkkUw0N7msrUmqG1Wx5sZR/yzzerTDqj
P/6qX4G2mCvJlhWXW0zpbmXBkLdP5JoONArGGi0U7/XBaKUsAZDpTJxh/RlMvUrX
R/a6BAJ3+fOBErtG25otANll2NSXe280A9lWPlIfc1c8VnUoNFxpnsyZB/mL5I7t
`protect END_PROTECTED
