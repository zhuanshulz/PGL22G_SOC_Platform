`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n+tFAIAjimbFM0g/IIPFozusAATeM8P57uGNwQqgYIqCNCtncZQ3DyYtCChEOKRw
CZzUMXLmf1NEumXCzA9jk2LleoRQ7h+o0y4YdZvwUdxCOrgAHGMbCDl0Iia/jocc
+IFM7BfurEJquXDX+IG+aPUw1WteV0dYVa/5ujRU47Ncr0FU9umVXXXxCkX0RBrw
kIrQ0YVeVhC3bY9M2aRFC5qKcBSwFQzf0h0ZgGLb0ZAaVGBh4dTVCzWbJQOzr+d/
iv2mImw6gSDk+sIj1zi64A9l2A+vr8oY3CV9RT4xHkohRddGRSElb/qsj9mH9ZI+
DyGAJyo1O1MGT4WoEGDOo+FAvlA7hX8L+UeeudSmjuF7c/WRi+9tnax7ssPHNNsi
kh8gB6xzcwtpnQ//pZ6SOnIK683YxsuW0MYcgfeV13mxtZtKbKp8RkORgEU78jLb
IsZo0gBGixyq9so92DjQYyZhQY0ly4q6YNc/fzCOOwSWZD9pWmB7lmzjiRquXwz+
4cwSJCMDm2bMtQO9dVYlF9gc1IPcnGq9rTS1LZxNCNj74sQuTw76CNjLoDEB0x6u
SxFUZfEDr0/Pkm1PZAR99vF299x2nTaLBaPUrbkcAIKJ1ZI9rMX/2UHsK/SL3fzK
BbC95JN43CZXyGk6rKB7U/8oPBky0EcprOQgpUikWnw1lAsJmq2TndD8m4822dZq
g3aosXFSpmQKrrKuPtwWOFMklRh3o8exsd1MM18tJNg69iGt1TXrgoJT7Ez7Fjtt
`protect END_PROTECTED
