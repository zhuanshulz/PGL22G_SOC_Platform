`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Pr4w3IAptEiidFdFgQ6jWlGwqWQBVTUR4DnQ/RrM5WY8miLW3tU8NX6EFZG3XaV3
qMGGFRPhmbQRXiBUTqw2xRXi/juY37MCDvyWS4yPhBoIVmetxOJxgeAWvqzHA7D6
DiHvmmsAb3B24iR5p84XZDYZlVyY4YwamNF+FSzmXFVNSpzuvgME9IBpQdfRjqwI
F92uve5fJ8pw/Ew0cVDi4YYkLcRjL/V3LeHAhSAX7yvn1k7RUosZJ4QCLOuJcJrX
5YjN5r6Rsih7ncsUU8VpRL/LuPoSpZEsA/Sso7a9evt7tkGBiAIF28vJ5ga2MKT5
0tji7XnTUviJXiFHmX+yYzxfldPQXnphNijvMEMKrcRz5UcOyJMFfIVP+ZaPKPJ2
b2WpGtfs9+7qpI1jIuwx5Bf9AUtD2N7wPNAQQ2xDCt0k1PdE1RLk3OcUDoK79LYV
wuzRgpWY8NajXuqJj1QH2I6Qp+ta+GesLBl7Ud0CVRdVfLvStNumMxeIAkIj62of
ZGMvuLSSDurOe2GO7alOTMvpqM1nj98qFrlN2PqP4zoOq8ZYDpF5C7+Ar8qymcbO
WA5ViEkO0PjgnLdad6VxXXsNn9aYQ1K3j5F34yDxViuQVhLujw0blWrOp7n26n73
qVUvov8Mo1jfnxPRitBaq/MO/ZpNzGtoQfvBxsaLLHS85Dj/ZoZHKRwo2a5vZNg2
`protect END_PROTECTED
