`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y/FiXo9Biv6cehraEANSxrzEiu1MwQfieBDDIq71FjsoEHf76FGbUcyuEiCL8bXW
vWpWL/0NN3YpZhUrOjsPeGhLY5EvZbXOZGXCZ5XthQKK1cxzXOMVKuAzKoDm8xt5
GxVzk51ybebpJf0mPIgR98+RVDUSvyVSUwYNG669c4NlkU460+f+ygZUwORGP0hx
QFAcqoGU3jW7PFmLLqmG4CQrQ2EP+TvzXHTfaCTj1flcqv1iLXD2Ic9Q9EueGvIb
LcXb2xzCe7ZPbfBs1Yi36ix7VZc7VNgk7Bf66M3Mw09oLBAW2ul+0L3r+7IFcebP
a5x/1tOl4tk1/xWsysbGoDNmUGDJmo4sUEWDug/bf0C6A+QOxviOLF8HwsoJQgCT
jlBi4uoUPxtrkiwU3uRKpJZow49DLFZw9KbpP4HjS7/Z3hmKamlEFs44pGBNKlKP
vQDrJgwkabsCPi4Zlq0sHJCEhCioySdUG3CY+LlBpAtqjqoyjR/FI7zYx7acG6ES
mjpS0xJKjkmqKzhk9nx/LqevW2JrZUD3kJbOv3WYLT7wRfhMIHlWguk3E0ow1N11
yxZhsoIlBFB5s7fgefN3iU9JuK0sljWd94lTuVCNSrPRXA3sD98EdSyEBXBA1T5H
LZ0vTUyagnGRp6biBL9SDx3FNJvnkA2OHPCuukTjjakGrmSWnJkpovpwi8XQKLzb
Y6dXMGhdE7YESMO6yq9/D0+v+M1RgOfIJXuRVvwlh3P0XSLlUT7Zg2sZtuaZveHb
bEsYcSH4NSvVmUl2nLsdZ4bZu/5t2UsiIz91oR+vxTUjEjGUbq/obWq7vcv39Dsk
gSFzU5ztSTxBZaVsNH0NcOGETeIC85gx3bVDBy7jL6umo5WGHpj3iDDY0xgFsHe4
T2BD6OxYXc/xZVgDqDfG32iDovSlj3ELUDdFPFgJiEPSfXmZwdqO1SYSnFiiqlFc
qRBKGrHxJsIt0tymVqmD+NJRrA5RJSEkMpiBgJfcoXCdPplDQCoCw3WyH1XRAXSz
49i4FkqWDlQtL9S+jzfzpw/DxIv/DWEE5aHvFeH4l1BcP+wfTDuJrcjhsGbRpUSI
quDrURVodmzrQdINmUKjuL9w1QvG+oaTSu3p13y58jJ7K8BQC/OVpan0rG61u16X
NMIA4PCndfR/0K1uDXm9Xe42WeMcf0ELE9KA2E45JU7qeG808bAiPFIoFWioicNX
vBd2VV56YPRBlEQ7sKvUxAFQSwNGI5i9U8o3wmPxgvPv8ZIcPJUjX39id/5wSC21
T/d4iolnswoERq1Yn8bOjw7/uUuwkXPPZRXiyayb0USLHTCE9JsAND/XXmtb9lHH
kHirkNvcgsR4c4oy7ddxaezhaLT41AhLrvD2+TtTosyiyeM1F8ZYLf3+ONe3AdRt
Rz5sp2UJo8subgODdYoC5B4NKmCwZ+9yHXLW9kGkKWSbAYDS4k9ZFX6Ayuj0Aj8f
6aw9FmggjJuDNur+cwcTIg5+FDJFNrH6COD8gJc7CtIOla2t7EGG1vDH6yn7MJoi
Vjl8ns3wiRfa+/wBPxk+eiJ+ONKqdhJCDzKbXwayVlAuFkzj2p7asOMRFIDpKFZ/
ZAPAOsAImmG1P4ytA0ODG3Gr+Jfk8TG1gnaRYJ8lV9bFb76XWanriltSa/vwYPPU
/dP5nSex+AxJiXmeUKDeuIVEO6ysNmrgVoJvvINDsnpMndNU0eWJ7Q3hLyFWdnL3
Q4vB5C9SRBwWo1tiv1tsJjia7oD0m1u8kkp8HTsk+sc/t8+rz90aSr1O0JRQ5+0N
KkvkflOuTVME5BszbWueQ0y15k93FGxYfrDSncUI7q/MGfOpV5qVDGOR8deG/LiA
bfrG6WF6sqMZe1kV5YjGBGwmxE6nJgwNo35KtfFdAMkJs69jP2S+p0DOso5BlTiD
YzmjYBKQqv5sK9EWpa8d124YkEz7Zphz8cvu4sjZAVvAtt3WZ1FqLhtan4m4WFYw
ecHtOU0nYCit1pI2fVajA8fLb61+L3IKgL+g3vjj0IKhUvQjHtfs4rePQbuQqkOR
jEVVP/n0tkcLDW2U3sjL1pXwPLB8wSdR/BYm6EneZYPXK2g7lDW6NIB+Mk4x8mkW
zO6pGoRY0130LVkkdfmTKTLd9nRFn+71+ZTLrTr+z6p52bKjNkVXlUo9uHsWSs/k
hQD2WA+hXq2tcj+5oA02HWlriIsuV887VJ16/hb+hmI/35HFn2eSGPk2bSYztKIZ
`protect END_PROTECTED
