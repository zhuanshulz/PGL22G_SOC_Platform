`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5CUUw2PKC9mLPlpqV4v9fvD6CFUfawV6uoSCst8fwAnXYt3woD17VZG4LWlzLgua
+JRTqxEXUhwV+9u1x/lB8DqKMgZ93f3g+RwewKio+Y0KkC15o8WYtBLkJ3dpg4Nk
3J/CW58MB/KOKEqI4NYcab61eBTOOaB7BGxodQIZINapElYSqDOzatzVPBwbhTd5
81A7xAgnWmsr7gZXKuPPlvEstpUJP/WAPA2uD/30FrmZqz48jeYAgr/FF303tIXe
ZJ3rSQ/+8khy+1tkyztl+qkwBMVIZG9jvz1XypDOia4I0j2eHYzDF7VPyOAalVNW
2XrYFvR/n29TIrolSevciCyQL7sakn7V74SRhfLYF36xx2ipZDe3OpicfVm9mNch
d31BnQHtE/Z4KSqv1hXQVUYYVHxj1TDXGDcMRlnLKuyEMcGQ4SN6/3c108S0y98w
D8VmF1+/56YTgea5t4ED3vRqSFBZUltudMFfsd1uFaIN0FSvmH16iAQgI5B3TPmA
wLNrMFQR/LJ98x+SuFutvTU/1pKSbBJvMsvCzwPUoa8Goo6ZQaB1zm3tcXhx1wde
rviZSYsujif9s1t5rHUnowcnaqx/O7h0CmrlgR4P94ZDXupA7G4C1+x1N+wvRrTm
AfWG6u5RQ7/i6HalpOQKP63Y/N1Scy1CB7vKwkxSYBSHgPZwPu3HYTjR65lo7ihb
wYQD4VVN6nwtzMLrKusCCCkbnPsXJmC6IBH6W+7iajw=
`protect END_PROTECTED
