`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m/TpYFwNSh7EU3KZwLMLAueP8j+0XkXwSzk3SbqT6Dqw9eiXtmPvXMLGeL9suJCA
ZSPoQ83gnXo2S3pZB/9PATiuny/oPMm1e1O4qeUpBn1b35Xjp33tSmJQFFRD9KM8
DdUDqpyBMnULPbdV4lGow1KGy+q17vQWFPxbJX6yYPJbSZ9bjPM32BUlYMhBVZ4T
no3IEcLiyRQmBdkuq0EWDE593H6Js/5GM05/Jogdh/zt2z/6q3dTlnhl82pBYVxg
KuNspzjDq8jlV5eyuLwqRQT2ZnBQ3Vtvj0FvmfCY8PDZBj7Z5FiiYFBr7DqmERNG
U4XdghCNtS5eLDqF0pG0Zgl0/ga36R/n+2PgxGVVfYlRVo+Yz5XGBmqz4PooLFKr
sKvAzlVBwULAJvJmGSn9pyah9eQuL5zEwYElno2Pw0ynyx6QP1XGVYBo43d0OPHs
c7Tw0mSgsT3sxo7Wa56t7QohX9pkaYNLcnAhYkgqHYSsupFpFzwBjsKPO6t4QV5o
MKbz45vSKIDdC7ZpsXnNiZAHKOkLzAPjSkvCsAGme11FrUgsE7jp0jG7cEMXwg8Z
vl6acaEcU2rrkaet5pkWd4aaP4jvkcfgF4l0ABYr2Np4jon+n6E/USDpX0Gf623e
pvpsmv2sVa7xT1JBG5dYTuIT/oO60FeVay928XP4yR4mGTYSZsq05j7bTtwkh68a
RAMBejOIK5wFBjhRQiNdCYJbOwp9U1WhWJMPYSDaAbFV/AvXQHer98Go/2KOMb3M
GnkNAxUX8ktq+6/SE1OdROKNZMaMqJVQW+ac68HhhOHijkLsdtsTa/s3gy4rIAsj
bUSMlSJ+HfB3IEOoeRNnbqDAFhw3mNL8NasVImGKrhqKsX6pN+tfZuM0iiR+J6o4
H/3ivuiWRNkFE2jWJ8Ny1aIOLjAkFuHxTaveYOV5XMFUhGUkYc/uPvvF0Q1E83MS
VIVNwAIyiDUhSLw/+RcNwrNOzva1ElcooUqK9dyTR6ULkojRJ3YJfzjdIYQFKq9M
ICf2kMtSvaJDdELMCWQYWWft+p1QJAI6VAoMSI8YJqk3YPSMOou+Tui8Fvmj2clt
BVk1BCa4KmQ7Jp9q1svTsUECmGHPXKyJI/6CRNn+pSHqcvDIZiBX+RzpDdJVvMdw
HS4lIIZTh6FDXqmKnrS7l1zD78+kU+Tp0rXCkjt+GeyTpIkeYV8E1+227H3jHIVT
tV9vTElldZaZta9NX/q484L4SqIlRkiHN4kQcsOStouyzpqoniyOk3xtL2lrxysg
4eh1yrDcLFCWV0C93TvcVs0nih39xnyWkzymaDnOXwE+CGNJfPqunBtaBVDlskJQ
`protect END_PROTECTED
