`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7Y8B43iYKLLpscpCM0JVI99UCGOJ3fzmeAg1ccEk8+PzGUbEVMVOk1lu/v9L6GQa
tTqhu+kPvH2DMruSq+NX0YgIFsGfB1KgOHQEyIlp1iUmcxOLahKBIgqc3KFSb7sa
jxpz71L/uCgdvhGMyxLR4zRCQMBfUjvLF8gHpySQMEIjZARiKPYJYweCyb1TqBCS
uiEsawR3eUpYNj+qTz6M8OvVHKjk3rpshU8t+NCD+bXt22WGf0NUfZ2lmoWJWxjI
5R1Y8tKortTYZ/IX8PuodSRzjR+wcqRhGpqq9ebcfz+xf7Q/9/0wln/KJEBN5PDv
fLkv/mm7Nrpf/14erC65SwlPuIkZW8tT6t0oE+tghbwGKeDbuF5rLeY6rwWDA+6C
fsCKfopFwUo2qHt1s6jaaPV/fXlDK6gDcmnu/ShVtCqrTNOIkjF5sJ+EP/AsvmB0
3nilJckPK2cu5o9YUk1KGr8DVbM9Bcwcv4k5v876OBEy/nSbHqiU11gPKUYm4WEM
J24y25ETPuMbaCmlcLQzfGfyxFD8GHc3caizjTD4mLRT0v+ORVubRGRiRMd3ziMO
klkbTtbxZtklLM7t4BvAUg==
`protect END_PROTECTED
