`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tW84DInkzJf66XMaGeKmUZ1Yco43b/4R+vDXzyn3ye9XQLsEP1NCE83itzHB8rhH
G2AqvM8RVoqr1CTsKXkhNOdv2c654oynnSFfIqB0RJ2yKmzVSIAV0pPPQh0Yt/Zy
5+OmTZjDcDV4yW5F8nsYu1Fm0hOxE2ZFUJLWcVBokCdLzsabXeogcy6K+XJw6nyT
+HFOyP7D9izeCrwFyWLznNHWRN9I1JFp3FE9vYfutoPEetZtwm4RkufPaN4xI5u3
rZ8pv/3M/zw9ORI+7r2dvp5xkXGA/rFq2iALSY+OiDRu6jJqzYIMU39wXzrYNtsI
UXJblWKinAw/YzuB+lGnideUiB/SJCDNP14x1352RpuQ/5nheexw3ZxqKeGOY3tX
aYq7IMB1RPF2q63w6Nmcrr3Yt273RVpYA84LrRRMlVdBGl/ol6OTcDJbl6zkDAnK
vBT/1io9XwD+LElniIfYNEDER0XN/F6hWSJzmdtUGkeK6C0K7fmNPsjB57O3WyiH
upa7sNgr/rMI2Bnk4uENHiYF+LbG/osYClmEguusl8ccTnWvI7n0vL6n5KsIL0En
sBZHyz3sOMNkQ1tWeW4BfOPal0w0opLI5VZ7o60ylWyaOW0trCZ761HPi2ljxuOy
`protect END_PROTECTED
