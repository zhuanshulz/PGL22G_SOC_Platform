`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mSwQJxJpUzJd6/H0paHcIgJz6XJnjLBbPRNMG3RldEZCe+z2rrQGt31pREVkMhne
M2PyFnCCiFpXWxd5IZSoUAZ21FlYqUusbj3FXLqa9Mom2HPTzmIMJGyTrLo9mOHb
8Ve4zBBo0PIAmH2J1qJOiG7I2+oUYhbpFcXN2taGkobh+AgrsPra5aqfNQl4ODba
bNo0G/jf6qhC+VK+6NCnx4KCTXSg+md9OL9882SAozPm8HmUKcRNXRyDQ10saovp
vkdrIlxxhcul9F0wh8MvdjTXAQCyCVnw8yfQV4ynhNMNFxsmErOIF5QgAvFUWUmV
MN1xhXXn8n55Kh5zmfVLNPefmfTBMs9YsBWHYtG0GMu+XAu9U1tAxf2ITV6Likx2
MAkRU/yS3LDKLGu7+KnuRXVfHscjz19hJbKqplp4K1KVQBvCiypCr5hgb05V3UzS
jt6+Vh0jUNmMioxTmmkrLNs/Vk2A/BzHKdpKz9w/5maUwGTNzgtJF5+U+lATBcmX
/JqvoJU8Vvn4gULj29viUIWhgFCo+AaT6hoIOmPmOJoxRI5IVrU+eR5Ts7Q8iGxW
Tv9n/ViADKgIjuUFgk7lSsyZTWSSAuqXk46ey8wbdgPAe0ld81dc89f3TghOG6Uf
RjdS6YpwdSW67NnodQgvf7eANj/Yy8iqfaoNm3jfwmwoOa+SaH1XsRFa2Pwe8jJW
NQwXNplSlwASLRxdwRLGvHVIe5O8iny3CTB7jU1ULWrkfECROj6KBKDtiUvsZT1M
PUbPdeeTn+k4t6ZHATtHw4o5FTXsmf4FGGGTChubNeU5Qr8t/iqJJ5cjTX7MISLL
KvFQwqvfWJynhchnfHH2Z9/seBgqRIIY3R3VO/WetgI4cMF3K8Z+duM6XBnwNdTI
nLT+wYX5zDuiaoAMcYFJhARMGC0S1rENz5XxI1wEIeXwSAHep7cQyM6cQWY+qRJs
jhtR/2xa5Y2e2oJEr1+bMJtFHgNwOInD9dBJX4CMdO1RoSrQlExs58VWFmXnMweO
tnuN0Vb8+txSmlBTT2qTO5kyd2Y4V11rQRCMT65L1NSTNmXJaZUPYmGjqX/Y4u01
Jsn4yNPnjlSNNMjGL7koyVi5jH61Rz2k2zYzZx1ZJ6vtnOE37TZ0Dt3CvTJYw/je
z2FmJew8xIK7Z1KsUrRGPH7ubqWqrtRYGgpUn6BNq3bVCnkIkYf1EMQDrhHKhRVc
xXWybyQ7o4A6w0JSHqlbucyLu3fYpCdUdKSeKZMkFFLPaSJW8vQzosj93SkiVCk+
YuIh8a0d9Rp9yGYSddcxotwPVSYpiEBFa+QgWjAlh1KHPEurG9AgzEcrMIzgpII/
hpIdEPIMYrV6tUlfZeNE08xJkTPSyzPgA0Tdlqe1Liwb9TnaVmrmn33yz7VLo6ka
LmXBZE9wmKpvhGKhVpY/O4MeXL0u0ZAgvwptVgh0jeSugW+gBScyTLF4MSgFhoDR
kYc1/Uy4qWIbyOhaqOseEbRGZjsG1yYthILaDqIOVDvIHMlBOuayd8bCuarDyeKM
lqwJbUSuim5NaeT+3sMtjA+EKwDCKmcObIxc9qop6MmwItSNpaYLFTttL0LQ6ku4
6ismbOyMKTXXQgO5N3cyjbgqg9ar25DnM+W9+gynmhsnCQbttEAtwGB7XYk/pVvI
dA6mFy59aVpM4uyhmaoaEDTIZP3VVm2VmhETUlPfI8vU4I6rIarZlBUAfoP4Ybsa
Qyo1jkk+WfUcv4h06oAdPcpQIJOa4n/kHBoiQqUvSPF/SKD9iM2Dtr6nVM8wOpp3
y6ny3stmCBVExvts8dEiSnyXe8Ndt2WinVl4piVVCh16GJAeXRZExFPbNvWpl6V6
7disDB6WCMq2pyes0HjPDOKA+EBFObkJ9PrKCUQMK2X26ONm1ETdQQ6D6/lyyTUi
yjVKDiGzo4Gda9egyoIjWJhtuBAGojCXU1gFZLp361sY2+uSHci2+mPE23HA0Dvi
lUw30NE3h15okpuH7jOe9+ZPl7t4V4ZdHdbrcSKjshZTvkq5TrhclPfaa3iZFHNw
CQz2bu6bv9J0xB1/sAaH/hUFAJvJ2L7e0YKyjCow51nO37UCMcDdu0lS9BLcn5p9
cgFJaG9cvnRKPTTpw4ZI+7IMNwBOzWLVHLuvOyv1G5NWDC2dEtFQ+KokKavndzgb
tkz+A19mRgY0q0UrBPg8bZTPUvUaom44aE8OUdtzNN8H2zMkjsT8BHLIsZPNdAnN
OA+wTUw/SrGej85lhoAllkltBMfQ4Y/c7ixrNp3lWgNwQy5nadWRdSa+m1XSbwVX
OS1nQ5ZBmhttlmCEVR9cru1RkTFwEKhlEOuZnARVL7hgqKcN+haM1caSeqC5mOLQ
MNcYrvTwiCurU3uKhbPwS/Vd8LXQXrYE0UH81tfVjWzrQxZeb5aInoKgoQmk6fKd
AFSVGdTfzEaD5qMJnboO/2hX4STfIkJZ15mxVDw2f1w5MymIXQDXj7r+nNCWbziW
fvjh64BDWSEuiT2Jo8iPpm5ipp9o+nrfw1EgaPaa6KnF3F3tpHoKDd1wHTM02r1+
AiChmMls8skQ90fJQLx6oQwzvXsjM2g9IaLxijJQMTwJ9zv3zOobu6HlQKClgZvZ
ylGhz+PBrywPdRUFQ2ytcF3JVEUlkB0b0VPMWQpcf18Jc6cI7UlStQkj/9v50rh3
dTj1HYE6g0ugGLn8lKu+Jo9fTQm2jWFDtLyidG7qErsUnqCEGPVw/09XbL4GuyzK
ELVU5g4YQbmJrqSDoUJ8afDvT9V4iOU9GgEGtCpmNeTol57iBx7driyu0cnyd7px
QYcRQ6OLzPa9U+Tb83j/Su3DtGvCy9fhfsblkY6H6I1CHD/m0NA6fKQjUUV6t5jb
t4Yn7ciX2rI/DO28jcdPUv6IPz7i/silTjJuSFOw2mtqrk72mAywA9BshF0MWiAC
adClUNfvre6Ho/LVR57MUMP6tdLYtKwQplghUf7QR3H7a5FCree16MRylvKzcy8v
SKa8iy4b2/f/DxJ3O2z/xmGrvBGvwUHlZuJAqGb7pyPZ/oAiPoLGRf3EajCTmr5P
UBcVuh3Uxpw6IRqbkP8khg1bP6wFkeis0thgc2AlYpFKBgtxHOgg3/KN+0U79bZh
5F98aodWkw6wwaQI+Aig77lWJd+XE2PtmkRM/57GaYadhLQJT5LDC1GlIym0/+jx
Fb5BSKROYI48Zx7gi5B+U9bRoU7z1ee3UzBQ+MUgzcZhCHaSdUhGRU1FjE6cpGU7
1D7f2ae1Hrd39kSc1+HeQQTbnesSeQ5gmYCadTdghHJUhTW7QueD61nxxyJcMV5Y
ahOiw+UzR7siM3a9a5NAV8HJEy7mygPMhID/rI8m5qjwaBLf3PTvmCn/ToAvz09Z
nqVaI5JVpA51RHVIEEecmnRpUwwTfqas6RcgQRi0lp9tZAFzECrRcw8DVjF7b1DT
aMfu3WyxJdlXwXMDjMvFrScIzRr/gQ8PqvrhgQmPHlrC47jVi8WDNJgpRT53Fafr
MMWarBW6E20BPlO0aYd4bDpc0QdFR2+7u/sPDXocKwVtbwgh2PYikMtaN4jK19Rg
TAMQYkUHvhM5v0odzMeqNNQFtEekMcUZU9pKcNrlZKGEQ2H3VBTAo3J0Ra1/gS6O
szZd1LNIuzFqxje9zQcZAtUxQbIIZITtGysjLgcCjySig0TFhoNfPuw9R2Q1cQBr
9GC3iGwlvIbXttWxZoq/iel0iY2pzf1VW9XkYqKi188naS7JhjIokSbYbkBdWEm1
Yfdm72gGZzDIjdpPEYyvIk0/aYG+ZJZzQ1Ro9P5+wiXzqIOoGe2K+H1A6NJYts/3
gMJlUqaRnxchkJ9DBj7YDK9wm7i20y+uaQ8wFjYHN/FOZvGLbjczBxMvW9TAKNhD
qFVQSSoRglednDhNYWZoF2hAVGINMMOQuylzg7fTZjarugjJjgSSo9xjxJbMoolP
Ko3VhKfu2anL5uYC2XuEJO1Jq+9rt7MQxK3YWqxQGI4mfvJSOX/IxCcBmBObFOpJ
mI4Dsv2UxRdxGjTUEW2/PmI4aSy9D3lfJB7mmACUxQZg/qVLpuC+u2ZajDQU55m5
6YEcjSybaGrkrSHQ4MRN3PB7m8Vp436GfpSIhVzOoFsj3HdD5/W1+Keu4qF9SsJP
fhJppTdow/dq4tqLC5l83GOACry6vIuByreA3t0eqquD0YLDwqsRyWYP/NQpbO4E
g3pWyMSGXkGfj+2GHvYHZiwoYwMmWQueAV0cxQDI7MmPwE3WHy13F4fe5rTzF9pU
/TaZ4HUrO84nZGY+AcQZBBXez9lhbYqUo1OBhHYAwr/Ort+E1w1CGyboqxF37UpP
LviGW5KyOdZ/p/NoCjmBcVp57mQU50DHlcEXp92gQqQZ/yzeyB4JtoO9IJDPeAcm
eJ5+LHUBGU98vzbmc0s8wdGmKGf+j5B2E9J6rQU8aMJf0jcalH6dbLkdAc3A6JWe
D4yhnnelGrF0rw0CrRDSduh6Ja5Tjge7DAadv5Y91LhRga4tvdLIqWDrznSI1Vle
6ZvYsV3V19rOsqix3QaWDFO9k6I3+J41vQIBs21/Um3smMIGiiUEEFCd8Xs73mwe
yrUZXWOVuaf7WdkJm+noLeUd2Xoe1Hw9nvXihWQUqMafNqr+YIkkMZr6xCdWh2Zj
MzlRkT7gJLH/sp0b1LO4D5XflvtAfL2TjGqMNk2RIait0Pkm8dXTodlhhLFc7TB7
JxCEMsAqNW56yHVCJRDzUTRXq1FgPMb0jmlZd0ozyZvmj8u0mPuMeZ978ASJNuHO
jlFMOFBOM72qWLWJ2lXWaxaC4SGjlNamYoJKn/+bMpcalKLTxhpBWh7mX8wsAw6j
7OLgRORSDW0hJCxkHjSGYi0YZG7BtmS+OB3cPNWAfawBR/fJ5vDI6kxYDy/Md7zE
SM8M/xCXjoUEj0/PwzXohtJ9GVPDfh/lR4s0xvwh/xDBDG5MnXeGzJ9hNry0x5VM
zoNcOjcEUYWnYEoLlEzwVg3I+yztlYAmsmMYhEFrM+d1IiKTKWxFgKyt5PV02/3J
l/+8tQgoEyVYuLr/Lutt0EswNlCRSPTdxNv1xdoTr3fZR65/FHClKSqO15ZodjX6
i/3TVVSWUgdZSWUMGIOyy+GpfpoBKzyPrCUiuGGluxVDWEnbgiWBknPxl8MLQbhD
aPB9UqrjPADIiBi18CrybNqrOti1xvDJ171vXE4FPyUoxq6UeirbTVPIsXEXZqp2
FDqNdahuZNRkQsMiCL13f2KTyp6D5LBWMUhYeYi7tD8odsftQ1n4hCD+uK6N7lkj
g4P08nlgr8NNz94zmKimsiwMW3uQhpQpTUyTcRmWFYnudO3YxLQlQjeG/drmcIDS
0yD/MdRBBedZpczp5v98kFRnJKtcwIaNo8rKp4xSY1nrtl7JDqdwIIV0U130uugE
4Q0REpwIIMDQ8AlmReUUAWK4+aSyBFaBCAiCOVM8yIZeC5EfDmFIxVi0kA00tbAA
kLdYOcRdfgVP2iz9dnXgu2fJDii9QAFiQU2sH6oORPp1smRLNwwPdIgY4Q2efOBX
F7ch0PIRlnkiG3ewACSFyPWyFx/0Qv5rWHo3IChrRbSidCJLyJaM/rSgfShJ8soz
mPP+GWo+KsAfCe3cyyvkhfyNVOHL8E/HEBLXz692uuuCYvoHTQByJwn7lRU2bcX9
B8hVAUJyYgjT6faWMlT9qDP48zlf58+VZIL72JxpF+YdpaQCjJ4J5OzQ71L/dFlD
4iFoLb2gA4QJbfddGQWrQKRHoFoFgyzCbIYD9n0csVBi2eiWp9dtgpuRA+CahoLK
B9nikRbyXFtOvbI+54e15tHnVe1kc+dp8cE6HJz6m5C9SrvLS4k1oJLL74qVhU9z
0vDCX/1cN7GJ2ZmnYMCCW/bUqeU1YIuhUSEC1laxi0yS3Z6nTKeOsqqld/qJfBlp
9yhITyqH4y/27Wj433czKRr6nOQeNRSEh2y9CoCvUQJneVPXXNOQC2w8Vy9g6tRL
yFdHEoHkQMovE4Anc4voe+QW3vdPXtiZTHrvgkGsA/UDsLaEcL7ZW9P8ynnA8+3x
Y23aO5qZ5PAjdpJ2kLAEENWJObOy01CJ5xxC1j9L8zlM/ui7C7M811IOZq6WREBq
ktzyeg3e28r9jGVl2jYdAL/vA3bl3hcu+7BOew0aweuDgpSJ9FqOZp+MIjAYYnHd
0izlRfm7GfJ9N49N5xFsWhPhTT+l06NkCQV/zljDbW4dmdD8jSwuLv1qpI7w/e1I
yjJrZWKupCLIseabJhx36sVxkjA7zjdjzsIbc0BiEeQgkflD9bOmtXzm40+9km2Z
l87nv2YGe3Dx1+8F3k0GaYZUYF5h/1t8C43DzNr0XeuyNGWHY5a1m4rixFlqf6wk
ZrPSu5K6+MMENS8DHE+13Dk/EgOYJeOJFF1rK3RKbCm2EP8wtFTCdEHshblctiiO
peHedJUB3U0jtXZ4WhdLHVl3don4Svm8n/q5ojC8Cf4HwbPA8ZtoghYsEXbOVoX0
aqv2XjMZ2nfR6LdLPjSGea1OLU6TJMwN0A+kSQOCHoF+ld81KSPiATvR7MXG8Jrx
mTY4T5UKyhfFByhfVKL3zsaGto8Rym7YAP1cncLdkyF59Vf3hwxw8pWXPykpZw5e
+gNM12tvRO7qy1p2nYMVTZOm/uo7IldwpGgEpFw9soNLx3vaBjAvqOYQqrJZ+ax/
XvpSm3MHshAGPEViCiCTQTvaKzFzESpvpf89JAvpaZRAlX800xp7cN1fAW3PKRXM
qqvdqnuhbSPIczioXiz7t66FtndqIGwv3cCe3k1SrWoyHwS5owzF8oROi81lbb7Z
EF2TFZBn2gbbQZvkdqD0tnAQLJE9S876HOi16MJE5cF0gjuddeUZsszTmecM139+
RYmAnkxbUEG7e36UwKthN97gzjgMwNzapAi1qfjb1e1S9v04wQaBiTXUDhUzbMBY
f95XTEGTIZLJTEl45+XGUp89HG1DszCA1d5bu8T/n44HdAsrjNp9m5YjsxoicVkx
b8llD6TlWpacjxU0Nuc9z80FrAMj9AraozAWXeDldLPwNqOyOJfKZlhk9QCkfgLo
aVzUOD6pr2UvzdprbEyXTeFvxg6SbS8ptaaz4gUb95UDBnolH0MVkls1PtkjXWfl
+Ql9EkDdImGo7hyFunVKyOSDE//j7yMLmVYBVluuCuFscJMP9YBrENm8fewtTjue
Ry42IUn2MK2Fpc9i4xi7s0MW/3XSRjIZsu/2KcRbQgpMJ8IR6sz9UiTT+tU3Q09v
460A4WlGHIVAmygxo0M5trwyvwEwysYHZ4VJF6P6PBDpBcxNYzylo1jRbUZEpGA6
TtbFtke7Q0i1JP7W53N3HHLIPis5uwjKdkG77112cmcKbw3mtU1SVKCH3PKkRDyE
ih+FcDSYHJnRjBIY2EuLVusVKfS1Xx/agQnnAvv8mbYdtx6CWnWnPniPtHYq4fS0
XbGdA/OTlKyKNAb49YLO6ScVCxq7F2RnJY0mDAeFaNEsHvADSugNwPs62A7pTpep
xIhChoLlmBn0ZUiVZQS4fsg/krZY0SrzmPBBJC//EBoYUi2JngKU30M3+prKroVx
1ANLb1ZB4RGu1BNE1lnXaOv/BmyBZEyunc7i4/m5PyudVt5FWwJH7KgdqTuRn8DP
9xvZ4zFCw4ov/UqcE8jBkoboo/E0lfxeHxPOrH04Dw44VREdZzV7O+l7yTMiMI0f
TonaFBijrWv/aYiwWS4qmRqZLAQdAM9kfThtOMC91ii67f6FgjYLZg0MO4mbDuno
L7lX9gsvYE+FMkEpUhOBM0/dHWbNYJrvIFG4d2B4KqGFJXVtGutPGngVhhnOX8y9
O6s9x9HfHUfVpsCnSMGMB7C/8m1e/UKwPlVYxCzWtVvSDG5QuZgEf6024NRij+Rh
We61XFl5CmCskqgxoKh5mcNaGsQxQVZh6j0TcfX/1rtUhUTBDFXOECOG8AZJa/Eo
a8wowR8gmOgJe7mdNIAIqPUpROr0CwoLPzleE7xPMDXDT5Q1LRVjI4WT+VgFGdqg
9Xfh/pcT2dlaKWGZngEun3F425a3ryF0CMY1uQ6KYmJYx67PB6WLsFs2TGn4iKi2
T9PeWOQPcjf9w8mSAHZJu5sfeEiHVJ6UySw8cXdTPVYerWlMex6ILinf0CxT7iYJ
ql8/028v/KWpbYh2EYoDEPvuZEdXgDjgwZxJIbKAUt1PzHM0HvPuXBZWVhHT7d8v
BzkoTnUJ9BcsIvXVmxuDgokS6shFZBhMJwN+6drK5pDZPmbDGCA29pamtKaWoQTa
m363KKB7T8E37tsHuLKC2PJwXgCd9ggAO/mhMRdenaCpVs7CryidEMWpBrMMU3h6
7bdg1A8uNOHLo1KPw7xTWJlwzaR2onSwdhzHKxMpdM/kyxUgTv9oe6DoAfD2NtVG
7060aIVSd2yrDw3JAb/Ox070vb4ALjPsqtLTH8uEn75FX2LRzfSJDiqbmE19enrn
`protect END_PROTECTED
