`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hntURt98YhyTd/GKS4KfaWfBhW8Ia4jJWu/Ygi1bsouH4r7kYcFES7GZr+T1FDFt
obAWmVh81m1SWouZ88gO2KV6kKR60A3xuqyh9+01DTR2ZDG6P3IoN85GpfmtLj4Z
Cgv0hYCHJCDX67Z7mK1BCAHP7iZrI/yzEGVx9uGzOZiSudlekn4RLd6qFloMUVOE
tVVhD7hiF/5BxlKa/92bAPcWOQXCkx1euwQMpOLxGvPyzWe48YGXGWAqhIIN3+5V
7jCJCyb8azthDCypIQ8Z5mkIAGSxOF7wyGgGlrvwqT5J+svIX+ftS1ohkqa9pi0i
SZmCm9QczaDRmYNx4L9yuA==
`protect END_PROTECTED
