`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6b608x70iGZsatUlBVwjDlbWftx6tC4UCaMX7sDhhaoS1xTX+9AUjsmB+KTl21ZX
zblkePyiGl85tY68289FtJkID70oPq6BsbJ4f3BZjpFz1P7kXxWxXEFEI4rPp6nP
jC69fWwdiCO1jAV60Zl0XOjDmY5EAUCWu9O5+b9ktVNwQb7wBmikiYPTlP+Wl7F9
hsaw1J01aeU19b14FrnnUsuJw2X9S/xQhM2nssrghHInBQGKC3e6pyt2jj/Jq70C
gRvHgRzcCqS8LUHp9snwd6Z0+MrpcQ2AJFHyvrDJI8KBsOZcLXBhl5+kKhWbLV9t
Mv51hM2ztca0Wp0Joov3Oc7FHvNGFv0DH/j8Ak//HVyDvvDunc62DmQgjsjoSnWF
iBjFnFBALb58szlsW0/mNbGO3fxFez5b97CyuvMdibZouvURqiSpi9Ng3CbEi9Hk
yIYcqz7aAqxg511s5BIEySt5wgY38+wmSXlZtOvj5fEnSHa+j7js5FWDroGZKsTV
QtkzNrncj1y4Be6W3eCONCQEcwFsdO6ZxXl26LUInZjobsxiWwOdR5uY0bn1TN6A
KqFDWiVB0h9g49qU0mY+QzCFd3iSVDud/bnEgGmqsPr+H7ohzpktP6OTRsj331t7
ojsQYG1/9MK/rhPIoztj51Xct7hzKPu6ax40FdKNu8xVRFe+f0GtC/Xl1WCEn39z
iq8l42xoQcYAVG9Em9O32CzpWGxjx9Mwaf/meiFlA8w9D3p0ewG1ZDF7WrVLDwOE
KPi6eC3mZg9zLgwEQEWDINQl9i3ibAdiOqHbXXmiUSdYFSJR6LNSWpH3+UxXXC25
noy4j0TX2uRAH98onk3/sqjReJzz7lzXBpEcc/IRuS8=
`protect END_PROTECTED
