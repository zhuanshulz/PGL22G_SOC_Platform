`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h7TND5ZZIj1kKV5yYmuVyciMezoPG2J547w7sA5TB6pjym89/1OVXNcR0bb4xHPs
cMJUgrTSgLvPg1ni9y+0EF1uzSGsslQxTujZDUloEtSdffiKf7+GgLIeKGBe5PCJ
lDi07aXgv8sbzX1lZ1KwY7uZSd1z9lJJeVSf7N05ahGYQXlPPLnU7iOxCa1v/eQh
G+GC5Asjugk6ZZJW1UbWiQlxksprHAnM7/8HeMQ0hd2zotRKXPaGWXLqivTAs5tR
Phg7WFQRHlF5NbqD6AJlrkwO1gqaxyMr6jEX7zR8P1l3g354ocLz5NQLq5pQIvXG
IiZdFGEUzGOf88/dO2eARD1sXsrXboeW9ruFBwjdwncnrDUnyRT3fsrdMAnJCgU3
6yf2yKTt4uZh7Z6v7YAstZ3OV5oRakI0nwZKV5+kn0FHey905p/bOaqm4rh9xycc
vGeMkGexFhB/6hDi4MTCd+zUgt23guP31CAHOTKWr66qHWB2bDiBiHuYsUecgQw0
N6iYrw21uXCsVq1PuiVW/hzyUqb6c0RL+08h0TugvkWkp4QHpKemfDkG77dRCxs7
LprQ6RRiTLPuqojMk5impzYeNtScgc0qmdmn3gB0X25rvculC3RdDUT2lhNydtd6
rKmueNzo0viE8femFerz58vIISQrb7YDgYprBBXGlOjEjFd4aNa0icF7/hKKwbrz
E7YOenCz9BrPCo3jaNjWxmrbBTWjPTR5XMTRGZmZlYZjGnOOaJCKg5T9/hVZh47n
D6PzHB0Iqa0X9+9Srps955bH6nwTAhgbXtIBnLG513mKU6ygX3EsvqSY4Pk4gf8e
BfKFkW/waVtrT3+lRQyKp03J+HQk/L3TM7TLn10JEiUwMsUn56tDx52rOuNHcNjy
31fpiDbzByW7gt32vwpPsMn+O8IRF5F6dYEr9gRryOEm/s4vWMv/64SkiGCzLK3t
82XEYm5gI6qIpOVCJKHzj3fE0u05JrlDEA1rq3Iwk8WXdkq/WQwOXPUx2n5cEuCs
2LHUETlzRQQXCJadksl6ZlBQa0p+ew5CGDrj/zJ67MqwseJIWddkw2Hwpurtl13V
J3RqViQj/Vn1lxiGnPBnZgJyd0z2mVEPuVXw5C6Brny0O2mYPXCzBSzSAXFV9Ez2
PIkRa/vQk0gzFocsqcYPVEzmN5p59q01kQ/Q8y+wXWXg/0mwC3zmjtG4yD9CtrV2
Gsjq8LXp8vJw/jbF9qBmljmx+BSUFnyJCwkpraasb4L5R+ChbvBTPt8+hF8KiriU
FqYipCvsYljUtOiE3ds365XgWvzM8fHHqACN81RcRtT2JsXuyfeoKjg2qFXiE4Zc
SMnEtFEEV50izyE5q7Czpe2ZPq9qE7vHI9fYticsPij7cPSCxix99dlvzdZCXOLS
FgpliQvGRn15mLCtkYeE6eKLoEd192H6/w26k5t+D0+0RwGRPogCoi60h5MWy3yV
Fi5zakMfH5eB0VNQPn22zcQhGbXWD+oF49BdQWPSe0GqrjHYSljkiRX3A26ZXu/2
APK9kOYlUVPGjCRdN6/TsmSzIvf1Tnl5xqobsG6B8cbacLj7QdAmmuS3K3f22wwz
On0CUZv4Co79J0OhsndKtjFrtaS71NuvJytUM13h9b+h1WPpbNgT6lEkjOr9sKo5
Cy9CvCKxMs+MEI9n3z398lSBFXph5zyNrqW2G4r3B3v45Gg1HJ5LUo5GLXkfxXXe
QCJp3JYrTlgWEp4rwpN946T8WoW3ZQpte1xNccmsTvtLTiZIWZ/jMIZPQS4ffPDG
dDz4npnNRzNZbtfowdIWpY8OBneXrHw0hiUz7u+kxIL59LcHnc8FssQnBy7mHTAk
hAMW+++YIuwamVpB9FGgz24EuS7dKnur8m5NWSfCFtwJ4Js4sujHuP2RTfx0yYCV
Ho9FhzU9VjXYGgXtCQw6U5r3riMJR2GSFBUchTXpQHcTnGb6QBYJt4xdfBRQwEhP
d3FbS6RT1Xvqsf5/XpfyycU+HC/VYVz+2Fnw62MOZDbgH75tNJ1iuiKq+TbvZOhD
q3eCbWnc+L2tR4MlyugWfvtRpgPrByy2FQw8wOzofNRrCXvaYIHkqrD+0Yufj0Ia
DMSuAAWSANstg51/RVZvFHDRyVpDEJ4AfGJka8EBCQjtln1jlaw1h+vmhge7tNyg
YxGVJwDqhpC2sWdv6Zw6Pqw6Qi3E9jN/0ttWEm83BVD602uVeaqRVDnIsF2dzFGl
cQcf6JRlxoEus6E0PtW2M4QmxVaK+uq34BMfczFEET4DQqNXKa9MD5QPAia1njmK
OSxIM1O97t9Zn+snkm+c9IQ8w0ewoXEd50yXSEfPuPS4Lj6wEKUuFekfuwfD64ua
mBj0KINTNGfBmQAM4qhRlJRg4psw+ihzrqNeaNzI/50=
`protect END_PROTECTED
