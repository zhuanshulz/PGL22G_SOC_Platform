`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NIPgFHQ1dWPhZb86LrG2FJtz1hKqg3YAzNlpuwAf7tzifLz0V5w3Kwvi2y3eAFjZ
efvCXQ0Z1USU785aAlHAx4bShS+gsDeBu/82Hw2uxXm7epSnHPTWJDZcYwZkxxUa
vfL1J3OP/PnBIeGdFPJW200fRkkncbw0Py4qL5cBpZk363vzqPpOWezv7UzPKdcE
m7sOVKcvb6pWQHiU/wvXp4/rTO0mWyQMIcEl7z8EHWFpCMJlWqkBUm8HYve5SU7f
veQncXW9Cqnwm32/rUwyM+wR4/5Sqgl+K6cVTxgOetD/9LHEpLy9QCoRFCVaFI/r
gMbGO6bqUrNTYmPEGRAg7JgYjMvhEguBAL6aj1sy80mwSaJ0gZE1kPT5SBodHJWn
0i9OaMzN46E+HheXVvO2OSuQq6qnpYzui+amPTnQD1dwpYPMpI5lg3+9kj3W3f8/
rCS/nTrHzCniL/oL8DuCSNqmqnfJrOLpXv9CAiuB76UZFdgltvJfBjE07wF2KZHJ
hr7XmPHLNByR7ZwCUFfPDxUA6UyFOz34Z0IdrVhNw6Uyr7vkXQ7e6zHzW/tCEK3s
43U1BBGgMHOY5ni6x+W5rUVlC8IQzsv2+FUoQluKS0QAt73g2qCDf2WoxqEbqJKA
qgmDHld/KgZRWiYTlOidns09n+O0+9Dt2vcoGNeO/cEL8HHk31IqPJAVKySncke8
qxMzMrhMORZrP2BlcK2+9P+kjdeHQe3y5aeLb0wyYojsoEmzKuGtGWIhCMdvBccg
oSl+iStq/nMbc6ug1ztaXI71jDzIjepUHnJd4BRqmJNv/pqcU2ml1Iqg0zo9pn0J
rUt6bRj56Xu8agfVAjsgrYvwkqv3a5+lSdnYzyP/ZpkuDMocotCWP324/cNW2gcD
kabJTcKqbk+F9+1jaq5CXo64df4GLmQVCOZw4rqemqbWlVw3kS5xmQ23u5cxrbug
NRO8q5K7eW6v/GX7MWGhDz8Y6m1vRshf6rJG7YGqMkeGqLXqhLeimQhygIzKMxMy
ka3QNp7W2zhVrNyht8pQXhHVzbTgUO7gxOJR7H461Iex0RPtmTfEh7VOAyQ6pqwR
76czeEGDl0N/Z+KF5sH+1xkmu0RHwqgzls5OjHanMpWhinidNkAnWnZPPY8xle46
XMTi+sLKsiVaccs7lGMJGdtFXtn7TOnQ3jy9B/aoZSJFxp+225I6ujh6ue4OZJab
gqyMcnEIm8q8IzuNKHPrgsGmD8pKliOCWzW8KEitUbh/ap+xJPyWYqfEG72oxaTs
zxDIkGcZ5iCKwoMsHIowX4eyN+Lyc81UvE+9mQHqx6udoZa9TiurnJEZDlMCKxtc
`protect END_PROTECTED
