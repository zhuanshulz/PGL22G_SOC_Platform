`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LmyUiMp/sSyBals1xRj6NVSaQwZiE9LlGNHT0gAfWxhDoa5zE7KBZkz/a/S77y/P
QMBkSVTXOAqXr3UaGB+haCmV89ZU0pOLEJ20As//X8/XntxHmnxt6evprBu7uYM7
af5L9BQf7F69sIqYTpMgSeEjyS65IthsvjnoMj//qeZgXSbVaaw5ifG663CbodlO
G5yW4EWPRzhiAqR6AdRIIhffPVv9m3XzhcsM1gnVY2JVqF0wxUwWTinoZft++yEf
tmiayDd7oaRD2nyQndCNWdPrmRLy4/dtAaxB2QqQYrFgwTV48AE6mjqY1wz9GuQX
tPH+fasrWTZrJBXM06JqVkexXwBELqZZ/2Z1ql0P9yaF/rzW4yhVKByvZkogmKpB
WkzUaG1pHuYAaJY6jCJb1c1IqGBUAyG1rwjur2tSTImYBU132fLAfR8snMLMfrsJ
dlApwCoS2cKUxJr6/add9dBq3dOWak7qEhcE3Wi9a7lDOZZKmgbtpTKXfgEF08iZ
fIreWGl9zVms7CzPP1DvyarPzJ5QvcuEhOhNXnNiW9sJJ3sTrzwjlo+BvwTZcrdR
/WrPDB4QBoS8dwhqXYkKf1l/jM3FoXR1xBpdOjEyy3VUW1bRA1qX/qtyY8GJHjrJ
Q8dGLeAoKDgfneB/7hITmJJ7otHKtAfwxHceodyKezinmvlaFlImrMOR4puR7ClU
ESWATCJOAAWaxxzTEmhxRkgCoWMgNtuGlibN2iOP2cQ3u8bCTekDX1XRFSmfQHcJ
dN36gnqM1OJvlQWZhxQcsSPMIEHYr5VS5Ff/gwunSI10WFOfW4JS35wxZiM9Jj6p
5FMEniGyx7X5D5PFKnZlHgsV/7ld9o/JQhMvLJRy44UdCVGJ4hyftKhvATYmzEVS
9J9BGWml5WnrbfpKl13+HJLU9GaZs1hYpE5AsY100W+5aPfG8noRL1xRnpFWMf24
3Bz1eZGQRc2JAXx6abUk1arUuTiWti4QPTMhHviRfibaNQY4SzrKkOO2FJBd5rVD
qYUFeW5PpKvZ0WuitPcPJAKK0vHto1VxnGQXitMEAz4ho2wi1mFNqIayEnAYZrET
SMU2UyfNyHtUFtUZpdCBgk+WVhkLYA3fvcZA7TfE101lSlxJ6WLmqb1wVMcVmgsl
874s1wOPxYQvRKtg4LgGT/MuqzqKm/LnZJ0yEkzRy5x0tT0Wv0pg3jGoYWdwrS+K
6yDUioYKY/VsQntZzN/Qz9d7AEwGh5txk8hVQsfPqiyiO8Je4xk//AuxdPOXDx/4
NdmSp0duiA8jyxDCSjTNvtEoKW/WRyK/MMRNnqG23FaqFBuN4II7uDkzxBD9tO9y
rWAlRnsAYynnU8oRXD/LPdK/3VdDU89eRqdx2p6NEqe+/+eqc0mAFSE+dnUu7j9s
i2RMHUfod+AdGvMDQw9PCI3fl5K3qypBtzP6nxwujia0xaDsnXaKdyPOrcgIG9KP
+0o6rj8mQ/EbOIGqWUGkgUMwuVWldTNM+P2omb6ytGz+yn0fCMpOwS7y1MxoCEhv
CYDh9JjrKTfVzmu2apiboDmm675m5177A8iF1BS2Ur1qJUNMbe9LX0P7LrAaQIfd
eFOYEVrIpQAgsCJZxakMyiYE/WzHJLjGzzovYaLWW3hcmbTtsaYAh3Vt+UcrngdI
9vGfGGqyQXK+VieuJN4Dlf6YIcC1TDuZ6OazvEvtXmcEqfbnnGpDyqtRvdXQtmnx
5Xn1ld5bEnGPAeG9f9d+6+w/BiYNl5sxBJiH1EAyjTNSFro1dIgE+Q7csRf4XFPD
IvmY6aGx6ge5OXxtGms9ohDFRgqdWv6UHg7COsqpL35t8FFOYAqFH8pzyaZ50pu+
dMm8vtMW3/oi9RMKIp+VmA0IuW9GXAH8EUkRQtAOYl+1j4AFv+hyLsTcr00tFinS
1Fcwou3H6I0f4PtLiQO67oqmspGY71WPz+svOwybT+Q0xzXHa87+WrsmRlxubXmo
+AtoP3s5AFBTeXpQjhHp5FNL7iM7BlFjBhP1C9xx5mJ4g7+DbqF9/VfycBXEAS2f
H4Y0DN35BpYKKncBegpBxTX7fAYGIkin7lasiQxtQAWw8Hd/RkFI81AJ3DTdGCzk
I/6s5y2OI5OnHteLBPr5cSnlOc2kZl6RXiPzdQ0h8/MGFM/+5jcmtBNDWecp3dk8
JpYnThW7VdHbpUZmo1qjLEA3o9Vm0xKW58u/AxyIkbJ1MLfEZzcXhJ2me5lGvIDH
q7wksDCDLHhMId7y3XTKrgTkcOVYMDhfDLmwB3eJK4+tqu9DIuFOU6MPZHIEKDZC
/BgcUJoqgRm8/tZ++fiEc5HYOLNbSzq6GkKsPzOhR4OVPKVthhX5+bywCTVq8aZ3
EYyVla61WBbwIplwQFAFx2zWL0gBUxXjJz8sjyVQYRs4350G9AnCYil2FkgSUCNA
cfux9hI/KGy9GLCLILtf3bUWrC2iIKiK+QXHHPzsRESqErywR2lHgwWgPeyscWq1
/0d4mMKnjmlFiY9ERW5XGNXdIr8B+i6N5vaxcnsbYTCsfyN2vS+vMhX0lK6gfIhd
WgemugshWGzwRjA+vM6T5yOTdu+vVyK88ZGjS4wpdB3BVBGbxLeYax8dQHuZN26i
9oGbOExCk11wBexYDCxwBDyqiRxOcq5aqjg+cOxI6bHn2hPmsRlR+kDnzMZO/kB4
x2hvchZbNnXcFY+11uQbG8PO64aWDdpWDj1u4VIx2+gyaM5Yxz1GLRhfrordQ6L5
n9rAoWnEJ2UExn6WT/eKFYXKpD+cKIFOA50IInO/FsW8Z3+gGzQXZlziTO/Rl+4H
m1iTxEKN9gbiCl91C37Vo1F/tnfm0TcBDfuVgWvKQbCI6wbcRcWYAsTQrPdrPf3v
QO3xTt64SXy8rpeA6vDzaspX9T9EESOPwxMkmhktayaOlyMTXDpqzin17mOhULhC
REKgMqDS6eCL2MQqa2USYaHtwhU0LM8KfJa7x2XzZxZP6E1+tByK6chsGT7IdQxD
3AWXPCNGbd15r/mHTPREMGwhBmXJrDILC6DyN3gHLghaqOPXZIo3+qvH2AXFGv7T
fmicS6xRwYbePjSO/7NCS1F7owUoNqYk3iYRd/QIpMxAkJxze6cBXfbIIsoqZvRD
SY9caQn9kqX5tEjvJDw1GJUx/5xFzEKIgmXzM4Fs5rn4tAMOJuX9LCvggBUs8A6V
Y7OtkzUFXXaOZsJNvB+Ce1PKWc9EYCDL1raHdHsWHT7IUJ/YkhCe147iyjERiHoe
XY35qpAzSyvOI2gwUYVvK2jMjH7n6j2+NA/B8wOGGiwCcgdjc7HW/6lN3PhdgD8Q
aeKTb+ioqZHUQNirTFZr6+nUNmZJ2ZFPtiXNkDLEn12afo9Ff2PhJJr7UzFmMtJq
YDM4WcF+2wfq26RG2u9aVcCz0G2IQqePbxC1oSywNSC3A4eIJylIjmDUXMW9LTjE
aInx/Azly1mPNsW8MhbCZL3ATMnhGJae3fYE7+aH7iGOnVW/gTbGgj7FEWRDSyAH
6htyS0g9YMg8nbu5HT1VfEM2dYQ13FWqyHNJH6J/BpOUNx+su3/A9x3JTpai76vr
oniPyT5/YJqM2OMdHkfxdXD3IlUhUSb5XZKNwh9y7uRP7K4dn7s8CYRf1Ikiid+Q
+57ZWZNC2eAvQTKw40dsKlTRHusxRgvJLMD/QYG6YU3UFTrRSayZPKTQzG7WR439
prP+YsFB/3ksM0ZFftNQfRiRM+zQ6rdRG1tL0OQl7yNJYUhDioFxHp/gNxtioGOR
O/U5FMvSpFaYPZXI1IbD9gdxWHj2sagcuF8VBzZxYPxCdX8QHRAMnqx+9QEsCWBx
ObPRepkVU4gdbMkiLxCRBanoO3Drz3Xe2SIoIqk9NYh9We13JDSlT1rI53vIKLaS
KinlWxsKkEQmYUuV3k/FiHIQT2KuMXAr4DP9kFK5nXt2/G0vrUG+itisc3o8gUzg
LeAPgg56ONwuG8suxuE4DHPI7xHT+N9gyReO2bc1c5gv6Vxn0cx2QpZJjZnZaYXf
ywUbpjrJN55X0arVTn1MyusdookhQ/jJhlrmErt1GXOBCOLI3tXgkDxhLWk72dBs
LCv6LY2LeNDxbyLWKuu89TskrlDm1v5+LWe7Iwni8FGppUfhoX9EA4x3IePSpKCY
pojUYquYyMbyxowtrgGgb77VmgWXAfC/O8mfqurhboph6Z/1IWBtMQpKvWIVFIXS
xdNFviaVI1iMX1VT/0r4wAqJAtuqV+goy5bIq+8JOLlPJdce2VDs2Utn52DZt0Dg
H5hFHaP6u0A4CqCpRSp6UFrPswyBzC/QU158SG+EfrmrTIDjei5Tv+JKC7ghjEpL
vXBgXVADw7qW3XZcv4hHOntKZ2ctq71e3Zx6jRC3WPdUsy7LpgD/oKnho+dvaPJn
/D8lcdAicNN+bZKjefcNAaWUKu892ofYaedKFTCSQTqHAw7snnb0xF9RJmF0tlTx
b/RFovVtebyvwBEuQYrYoFepCFgVfbCQZmu8VJqdIN6P8T0X661YQfhgWsGqpZb9
si/cvyvwAWILzFdsB438CpMZuyQIMf+mW87GVvbmABoF4DawdFJe28Pjfl7Z4uvC
72q3LP4IGk396Ou2iXROy7UB31TAuNIHaoLt1LX/7EoF2aR0bwEf6AW/sep7sK1J
N1xj5cPXW5L1BRPWaqKoYtT9n3xHeWHwvgUDrdDvdUFoTTbiUDnJfvgrV+GcP3P+
GMptRaDU+ESip3DAGb2iXp4DzJKv0idenYqbBjo5X/CYfdNuE6XsWZ42Mtgh9IST
hiTRP47BMgR/LCyCc1xpGDWzk4HaFOFJorswo6/nHiNYSdDJnkVVLKabHXdW+Ej6
Zf+5n4RURAlJOXbjLeE8Xs9QDVHT3fPLp0HZpgZGFtpCHQdiHvkmYFtdmIwK8tnc
QJJwSq+wljj0yOGBxCJVyhxhd3vh8CNydmeZnbQLl3a9ZWxvMKta9/shaKRPEnHJ
n27vKch0o/+kb5ED0aoMSP3k+ErDIQ38105cXXUVtw2cZ7tzg+TiYpRdWGKBpPo7
Olh4a0DGkEwWHfXsK16PK/LDE0C41x63VzzhT4CTkKigsNkSy+kf7nLHDbtqtxBN
jdNrBcVLkZvY8Twxo2cpEnjoM9p8nNQGO2tKnhWwJw0Wq5lUs5bgGBQEbWsFhY7v
rzBzk3UUapkFKP1YgOEBIGQGyHs53vuDMYM1mcNFFvM5TZLgfRQeauVysv/n71GR
ONEaA9Y7ZWGsj8utT7c/PWI7mw+uER9RAS3C34IpYMC4muvizHShenf/HRKE9Fjz
fa2DdspxBQcrxHSKgSh3TyTXtIjJCgjwdJ5sC2sY58b3BpAT/kGZ33Om11E+GyJe
qXSijO2bcrN2kV97snA8vyZwNwbIGqF+A9AB9Rk67H26/RN+CRl8NQf91XfIjd5y
OVkzK7c31Cj6HUFTNM/QaMm4XsbRV+XZ0VK4vv7DvSLmfkCOkVqVbxypoiIpM/Uq
36calcCDvU5qJlmrNvLPgjw7m6f/NSE/yRB2jnDmGSSuAp1QYEd2u4VwQCYm0kts
RWkTcG8tqU2rJpfLP4DoDREfmyAig9JFwSGYqVBism8Q+Wd32VI2Rgzli8P+xgmT
xS+KA0jaW9IvXMYonH1SGa6H5urL0LO7cmHW6tZVsNyzb96ht2FiPMrw/KEqWnhh
/xiT+I1ZHoyXDHjKxkX1GcXdXyXp/gBiZ4KgJIiEkZiIu7D1IOjNSt4NDSbwKzq2
14OagfYw6XqFMGt04ela/LWW8rPf0ZoXaDIxcWOGI5UeOHUO6RRSzzwKS9MJybG/
82qXk22M4VZmMSJVmTXX+yMbUQwxZtTlZAb9U7zuKCMutsI6MARQ2nATU0bYKx8W
tKXUpxVqq9YMv4FBNE0bESO1EO3Jh0n4ZK30Dp/5wAcrNeZuftLDoACg3ZghiBH5
ZnGrUz1pR7Y5qrdV13Kuj1V0IrPcshMa8aYDFgvdGv5Z7uBIEF46Ss0pvCD8xnYI
rYu8q9QBOVKIbmmz1VVV9p9nUjUE2SWEqubNo6udgmeCDl9JGAcIOdpVkurEDIm1
sWOTCUfxXeI1wGeOgv4vCmZdPIBTD/Wxnm7AWcyshZzK+QigE09XkvqfaCE1GfuR
Id1LhVj7YhNfPIsWIPvMvABAsdIvlttjMXOtkdzvR7NynsVkZFh4EG2I3RiI3rxK
EGZhQr5/DxFULYXWzRgK4/9tFroowThAHxzZzgit+6f02pXBiGq9Dyh8QVSHoc2z
hL460nkeKNJ7fWSuYWxOald/GLcX9L0+t/xMXhPoLL4cuq4UJCK4FpIK9gqY3k5f
OiTnLtactN/l92et82MTurFmd6c81F7MxdJZgSX61BCGhC6C2JP/WbEjRc7tYGAU
aopkVel70MO+Mxyc46aGld/qun4bKGOiOuOb20eou9a0quLFIFw8wCl8Uu9cpLLw
w3ppbmXNmvF6/8XC8q3tkN+sKvZ6jde0leEH9fkmT2zs53y3sg6UliEq6n6mH/hk
V1dBPCnE4ih8W9GwSnPn4HauNeJw2lUR1dajt2x6edKMCVc/+KyElfxk/BWGozEt
5WE1Rv5UA13Q22Hy32JV6f9SgJUNbqR/DzbuTV/GZdBfD9n5wySTNOGxm/8mFJRY
Mex6/iQP6R3LnGKrd1LaybtO1SlCgyGaMVGR5758hYjrASZUq3VRV4/BqjUPSRyL
9uZx5aHrtq4yKpM9o2gocAfqJJRueh9zUmXImqQI/B3CBuKWnSM2vATcTeTt87Dv
jNxy4r0+ZA44U3VS6ashAwOh9LRT8eepp2miYMxbtU/ElBOoihq3zV3DLv6JzO/l
1XID+AhvOLCnGl3C6xDZpDJunTNEJFBWdyZzHi2VrklIrivozgrQG3XbZGbIpJh6
DuJHOJvisxhLViq98hKeHX3S/ME80DXDXZ5+UFRwkUg9UmTZv1i/wQtjiG5YvsXV
ovVXrazSk/pb0Z9PpmcicRXL06ozltBwMsw/lPNiamHRTMm9FdFtmYVvEUq8NBtt
Iujx2dP9IuyxVnvgncmEFSCmB1TJTagmCdRzCU2P3x9/T+wgdD+yckEsdVcXWEZO
U/JXVpL8XJlI/T5ecuDT8SJeAGajV/30+JFfXH9SxMDBaUBw1WwN2mY9sZsUDKiF
sFAMLZYnEpdoHqgWkCRKhlB7zvHf+NbRR6j/4pxgyINxW2Jn/WTZn/Obd586ImVG
wMrRxjMOJQAo2k38sUbeHIGh0oKXnxOLxlmFxG+t4/FthN85YXi7mZBLY75vqzuV
Sv1sdV165oDOe1qdXmfktw==
`protect END_PROTECTED
