`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WggvC1QgRYhKrBReuRBhuDEVqWZV4ca6VCiAYymUM6kM4qZCYSBed0NOHvenf2AR
rfql1e7n4mcrrK/akacpwL9FkiFzblyEVr94EfnPOn7gRI+i7FlxuNuMpAMKaMFY
HL0t2rO3kK64HuooX83HS8YIbOqIlVBtdJzhIwdx2XfbshqRTdeQ8RmOQJxn2Svq
b6UcLbgUR/6t0zehpp+0HqmY+rQVAgKcKJOyAN8jviizCzrbaeF5eN7vBpjGD1EV
41eLDlE0t9PR3p3wlgRP0EU3i4qS86b3sai+8/d/WGBipACozA+wAvvQo8uAGvtG
RJ96QOnrVmtiadJ9eKL4AvkuRfd/HlyjUz2ArV2u6F3bk0+tPT4/4QFqE1cr+Biq
nwfHSA64C1ADAtKvJBZfyTbgm/MJioaoCllL48xy4pkzxq/Ii3jfzxAAzMpYhJdy
d7dzSxiklkyLdZALsuSOq8d0jgSitUyvQT86HqoAly5QcA7fnjRVxeme5zPEX1mM
Fraozx3CgQUV8lKXTz9DbbxvH4v9NJgUZxN4/T88k0q3JOhvrxNSbb+qRpDY58Ot
ToSAiORikA8dHyWyfG1PGqLPVKhx1YOirTYeFVmtsG0werN+DQWIdfRZOq16uTZX
Edf7GFupFJNMPluq++Yjg8kZY8gVcTvF/Pz7QFcXEQ9xUaFybAz6OMf1QpOlmBZq
EVUhSJicWlVvsjE8KJcJkz3W+m1zN/tevjeqPKF+elFp6q8ipZp+wFkFrmpjn73K
+1x1n2IfCY3mRBRpU8f4K0WM4JmuH3rTmHTIBSguGWhxU6vCF2NWMU1RTsW6WnDf
n37hmvxAUCME8ThJHJKd11VkMftyZ1y0Ys/KCN0gNjTwF+f5+LlB8u/LJczGVzag
BUH2XWp2FZQZCR6d8HPgVBmGtP1hbVAewTLj8I193DYueQ/UK8fLV+0f4fPH7ZZR
0v6EW4tylKmKs4+f45dyrwY0+ncBkCb5XzIt48EEwSWYUtq0Xd07tQ8DCSa2EevI
MlkY+htEExFER+mGr6NVXaAcy4AHF9/7CkQnxNQqdi/4WbeRze8uzFHdc8lUPGGq
ok/lsXJWfMto9YKElsxH47EY1DSJRP3C1DZWMdFBF6G9Td+laWNACzDsg6mSlRXx
TBVCoPhL9zMLkibZMSryZ0dwbYmSQCpHYhfc+GIW9Ol2ogDkjrUF9jvM21ruf2dY
zXqBOjilsJrndtx9V3bJkF/D7IX0hDGZ6sPMY1WT4wdHiRJFkXHkcpXcIRuGl5qG
O++Gq9PYB0S2uLy0mnqrVty0kfD8G2MsGntaHKWebh9Tgp6NsT4LUZ/3+NhSGzr0
KaTvVQbAWB7SWMg/FpAHpR1EyNlO3hn6ZJ8Mpl4MeRGhMk40Pg+QvghJi1hx4Djo
MUECQ3GyQaQKNuU6fXP5Wn1NuO90kAcvhVJ18FcM/vq+d7i5KU6xPf+EsNf8xlim
QVLhAF2d/Q9Jy3YOBBg9P7PyJY5nmERSsdufRa5Uu45Xz4FchRAgMkXZlN+NzfO7
y9c46l6wKMiyJ15oT2q5u8mg6x496RG83Zg3eZRi/k6OASyJbgd1tFGagg47F7nN
fkc0wFziEC/dRT1S9k7jY+/YMDyXWsa1K/i/PtuOk8Ulro+kCKr9t3LieO3cxDel
N8XL0PKTLj31AVEmFs9CZomMv42EQku06cD0uIDWbr+FgWdFf1OSwzDL3JErOcei
GevhbQDDoKZjnPoDZIUZOPswWNfK2+3/F+1TKIYUtKz71BJ0zjaBpBltWyJ5/zEX
R0G4y6bH+bO/FeayE6R/7GrGPNnpdp1KNMwJIW503LTUZJDrVxpPsg+fnHq0ppOd
g6gllxz+jpZk2YR3lxb9zlbhLfXxxX48ShPH+FubQj5UGZFG0ddP8teHY5dulDnT
Gg7YvQTq23U4+e2hko3ANuz4QLzikT1RRsEBYwHFy9/n6UJ8WaLMMU5ms3lRMr5m
8KZZvdUS8D9rcbwJ5atmTe+QA2w58hQ5VOlO2j9fsG2uvFx8QjzB4b+iTypgFtSk
hB8xoKpBUf6cX3RUU+ipOHXSI5TLGsEzGrLY3md0YXhpYOuYmdIs/Qgq99FGqYeb
OSxkHkHXqaxZV2wJ6v5sKwBSNwRl6nV6FWIubqDLBcPdSN14cdpRRoq2u0a0Y8cV
bVUH5DyLdLP3arD/nG3CoOdXlKLsrLyYDRYTHWnDrP6OPbjRw07uuLOAbAlvBOIc
nkFjAljxa0mswYDW6BneKVxftmeG1KK1IE7BszmTkTIK6H15oiIItplNOmjsM3ln
qwoXXhrIKMBrNQwXOMK4olLqHGGEcpQvt8XPU+CBS95Aclr+63v5hrJ+10VFQdKj
VfqlIPneSsH6Y090VYzAyfhwOzXcBPFQyN7nhJTGCubDvmL7/Jcgo94xxadEd6d7
Eh2LlDQjdnqeCKYEADWSaBxy5z3TO4vsTULjiX685GcXi4lbJwBG4uBEmMfZA8M0
ZkSE+oXtaBM+oqtq0CtrVRWErY8H0mMGLCoD6yRFG+t6eBEeSFn+d3/PMZahErKv
nksOdlmmESpoLc7GQ5edWNyNWREokFWBI+NTVXBLl+jfroyPsPbCHJ2bdq10HUej
RSbjkd680Vs1AhiSBTNMAPwW1M8JhIw4/qyoAE1eJwG3bcY8iHsz4C8NZ2+Wv/9i
ck75Lxnmk/2AcKb6DsIbZ7zEgu9rC+BIAhWTLNUB1ViZls79hBddPJ1WOhR6UKXS
auYRK8PH8WCfAk5rDtJnEps8BWZ2yn8RUm8r1LwLfTIiudK9hUHupEtwP4K68yU4
rvtt2I9Pv+wagFrpTLM2j3RQhKVXcQ0/bUJl6DzoiswJI50jZJ6quanXbTORtCex
j3s276902rGBarIWVqKUpciWg4pwloYuiVRAQWyy/FyyCIjPunBNQ2Nji0U1EkbR
Qur6qd6WzO4p10W9w6kDiNMZTflAajYoJwqpe2mpxiyx/f859FDsQSxrW/TGYLjm
FUK0Y6+rUNebhlIliSOktQnEoEjoXSg4rEDKMfdtFITf1eDGne+D+fDCkOPe8tNd
HPWGSp8R9NRIeUZhnHsF1bC4NeoCnZr/iZkPbPX6WX5UURQyLFKmC2/g8F9B3+Kj
BvMt9uCRuyqNLQoeTdsUvtUbeq5vE5fA70/xWka1nDGpfs2glz42AzVniOw6740q
Gc9H6R43cg3To+wYnTFs5s4BeeZCX9jhRwxaNHefVePNUv3I1R9XPIxiwLOTmrrH
gDIWFZhFYKEjDLWZGtNBvFiu3pcMZvQeBitk83GfuQHgOYYDqxCH2k0YEnSRN4X5
JbQLYuTK6EUIAmj19N9DXTAhsGDPJQ5xoM5TIhckipER9vZwsxVkQ4wJps6aclM/
OzxfPePBEomXm9eSE4j6q76IHNH1CRkDNFsSzO7tDQ3dCYKbkUGZiMaQ4ndX73lg
D9whyNuhyi+KUs2GVPt+PO7kZ2NIjqGj7vAvIsrRn8yHnb0b/gU5haHs97J8vuhJ
QWvIxuoVRDQ/4tyWMDzuP7uEHnf8FS256LgN3IMUD2v0atONti6JRREimDJqRyBi
Rl4cPmlfMnDDrt/ZOfr99OT9ekf/P3KhdHVEiBhvUx3+LLkwTgKDaPnQqfV3g7sJ
4tsyZPkkOLNZgLKI54ReJJfO9iE2F6U2Exliqsl/8ZMhTDrNmYbO+skRFv5130a8
KeGCoLnqp1vxMbhCq48qEOABaSXIEeCOeywsw3/luGDaw6fQUUYp2DGlsMwjuCFH
HpV3E7Z1j453qYzA3QjGFAYHfD4vYlklCVb+vgWiMUQnJp4Kpn1zdd9/K+y8oSd/
iFcpg7EcSAAOOSMXSkkugD5SkiANuYf3nkfAVrHZ55kRWSwFXlnHlPbYrNh0BXi/
1sKASrTTJK4KNbHFhWFuLoxDUhcI1iYw9QWuuaqoTRJzSWL7it3fMdjApimVstA5
xGVO+ha9IjpXvBJ/VVaLzaGndNQFsLdWiBiKpuD6qGM+oE/D/I+MeZ6ReWQZiMNu
gF8p7JXMZs7FRLKH2nBT79HFUHE4iFVPdtq0zsnNVqYTw+t0qCmcL9UsrqRxDsL7
nM+s2vSYIuM7F7oUi0aaxfomOFLzx6LCu99OaT1cNknW0QtesPs5QH7QDHac5uCq
kZNDHi1gu1Fekh8+JbiYKTlBfevv+t+THULL6syKlzNXzqblAkL2l5aJoP3VncoD
qb9m0eVUQXdS+n6+i+w5++lkGM7TXTfmfyJiYfGS6EAV3UbdYtN6JGIhd/QDitG+
Ci1XsK38wpifTN8Onz3iFvD0dIzPQm4rEmelhcQ5Y1fkZkrYUUJiF2KoY0XppZFU
`protect END_PROTECTED
