`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rp70lVQ8AaJ6t0bV/L0vbiNcXMY+pyhFsuupnvKY/5S60850SsiR0oHjN568V5zb
illdYs7tYPbkOMsFoASoao65rVozqDhY7ch8xcJLa2C76t/uE10PSIuula+xpG8d
hLlXyzoMJiwzLpX69d9uDa04/amt+5/C8Wk5vBvFycJ7uwlI8fWon0jXDNVzR/0U
vrKV/QvaPwO583XDmX0Mi23jx2fTkyOhq2lbhVC/5qGoOFKWSHAqaqAbpD/5/iHa
dw401t7XM7SH+tFMonrUreR0vWUCt1xGwKV994vpK/fFSCPb2OOnVgLKu/dhvd47
1vXXo5myEeQTLq46Q/ragZkOeNzCyrbkJJ2M1R3PhcwHMJxB54q50BGsT6u8Wmde
+huWhCPPebqm3G5BzJhyxv0waLjqMFLrbqvco/k+rv+0aiugkl0DeX5gzDQ5u9eJ
mhyb/gxIsiSrSLIAHRK7oTxNjNh4bTgxJuMZA9RMTQxwAz43hSExLWCm26eEO2WN
kMiifmA6hjU3I1vwuIe4E9SP7IVkX1NnwnEso1dilqbbjism5tuMmVA7LfUQAzY/
SVJcc8sy1S4DOx37WL7ptiC0N19WocxxAz6fPKTGY/syKyNUTNiQM6PsYb+uA1Da
t/CiJxZHfTcbMNqlbfG9kw==
`protect END_PROTECTED
