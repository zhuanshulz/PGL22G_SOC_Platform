`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nBst6gwmzWV/Tn5b+OquXkdVzCOHA0yZLvl62ELWZMlzF16U7WOo0dUpPez1MbXU
qAZploSCQOnGHZnxU2/hsXDX8b0IbLJBWbfIvW69iO45gQAJxiIFtSorjqkP3N8/
8smlDtD6ALmfBgYnrz8Z8LEqtpRxJi0MfTMnUD6xEI3La971Pe5ZZDw/qvTyc37x
HipSSEC/4rX/acoT6K1aAm6vsNKaSZKLEcWGzoOpK0fRr85PGZ+fxUJC2N0Xe2A/
kJu+dWNVMQQ0yenr4wLS0YXN1kQjkosxt3BFYntPG0WSpYlfStnRe77zWliFqUxE
HxbuID6aJT1nbKZSsxT/GeyqYWaP1ZrW6tbA0WVZdJsVf1iPP3R4gPSxzk3WcnLg
IkU7qxxCUELm5m/MIrCPjdSMYV1aNwBSuNIbRVLJMSfSGV1o1Bye6yGVieFargw9
3O01YVzg8hGtA5WMK1pbsZGVWjiyKuqPSsPf/pCBRJoyFrfMast7S/1yF09RCw3p
KjRvt+40wBQgum9PfWmH9doRmoFC5kCb11XmBwhREHZluUCp4CJf7mvDqNAd65Fv
0LAfPJD8uK0KIa0ic/bPavFmgTZ98TMHFjUsdA+8NCeIupTJPrtOsKRl71eKYOm9
IKMOstf9uCMQzbqYf4z1NJXENxpCLvM8BuLUdjNHo2f1hAWRdU4XLwW+epXimjU/
kacaEfHAhWWAvfm8Spny0wBQzqcTaAH+lLLfqv86BnwSzWt+lKwzKDQbPc45Fl84
tp7XUr2JDSM93eOrww0WPUHzvtE/t89rZg+2Cbw9EDWPUVhAqDZboTkS+91XhFuK
Sywzv0w9/TIngJGFke01NDSJOZ+WQDzKP6eC4QQ4jhXFF6bpXZb1GOrIbIjsDT+H
TktiWKyyULaB+DzKsB5nN+0cG0UiY2cZ16D6zckFMpyg8ac6DBihH6UVVWqa4b1g
6QY0cibWnnOMLlj8Qq/nFHXLirQaFSrMjLhM/HBv4FbjJ4egmcTaUJOlkRZKkR3U
uipKnHrz9xwqnQ7MJvAYxfStviiW8Kf8RShoPte2/EvK9r4oOcdUnZjHAKnMJrwf
2RwlRBQphyg3yKqse7MwR2QE597PiKEJjxwqg7VWgMYjK+Hl1m7jGFaQy39udsQa
mAD7P8ul0FlSnavBFaUrQJEJqQJBKFkPsF2E2NUT9us=
`protect END_PROTECTED
