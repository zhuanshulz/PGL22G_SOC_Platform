`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RQBIiivSar5YkuDXcro9GPjPxq75a+jxyKvi7MSFbsvNAtB8Dtj85jDLtyiypyUc
YmGIQHrHTdQydXUrP3kCN6sQcJcy0JqVsqAaOVzHjcps4pwtfjEBs+zshB5deCnV
b7oV94qX2B3NyJjQxvdUQc+Rah/BsqBpNLDx4ktYsdL81Vf8egTDpxkI2VB4dcPh
Br0Dy5FHWFNR06E4Y7lgn66uxTmtduSzBtmetslyFi3oI1rYoa8xx6x+WEHSUuKe
uGFbTfzqjezMDuNtbHSKzT+rDWQ5cetJSF4dw9q+PrQftr/u8fZtGvGYZy3ezJVq
u/lnF6qyts1yYdIdkhCDUcwjKx62/rkFjXm4ugel74N3uE89Maow4SNm6XFVxXd8
Bo5QH3EteEv/1VEQmZwY5IHY25RwGuYSvZbj0tWp5nWWwZHi5f/pWCUg8dq0aypf
tyH86KcMzu7HtflP9bA8riL9NyDlF+RGK7KNUeD6nmFdPqrC6OZQIb3SOi2CV5C1
zeThj9zj49Rg2iAfWlDoE44ycDXpF09by6httJeFILe508i58pWFpFm3FEJpFesg
OIzVvjpyaXUAaXnr/tVaqFFH4fitNJboN8TftVCLM5jY0XNriaGdSrJ0TlcInQ1p
uOqTNmfSRodXN40CtBak1qwNYX1dY0L7A7Nt450eBqhkkiOe2KX3ITB74beycGWA
Lm/BR/tRvuP5Wp62rRIzOZT1AnWFaum0KXd8INlMJLQfFg7berbl7FyJyZjtPtcT
tc9sA63XuR3GsfoW4Eigm+ATzcfocAl1q/Zs5GzI+3aItK4Ykog9OqbuMB+Pvc9M
KP9ycONyGo/Sb8eqFWQE7ExSMEZ4+5b8g9S1vuzOIf4iv5uVufEtzD8tgkl5W3xn
shG+vRKgDiJXdqVFb5cnaEXtx3JFYmtuFKRwC3o37aBLY6WhjEyh54+zWcnGpq8l
WoPmPVzlxwV0T+2Vsuw4Q3/IdsRYvFbagAhC7vumoi8aJhvA6aBxhYxRR7fGQGg+
odyx9YXNX3UI11K073BtjKj4i94FifbCURRDRC5+N+nXBBxu8m4A4CWQjMN3ywBi
OyuwET/Mo8GYrZ+ZkQdMvi4Y4qZGZx4Q/lVCrIEXDTFshGklZ9v1C0lxC5h11Mm9
KJomtW7l5NmFaXBpg7s8d0l6gD4V5gvNPmFfUPESEbSosKCYxkBC2BJwGevWePGx
OXcU3J6xyrrnI1Kq1L735kc4JOQ7XsrLx1JcvnS2lpavZDwz8qqplex0OIDDZ/Aw
DNuKG+WHkYFLobCt2K/pPoqVArG47uAP2aTqgfKvO4goeKEIyQHtyyvvSAWNbNIk
ryALgL17k41wGZkw+cjXPpV/YSI+cE04mQwVNH6ohdPIZAio3xyrVC5T4ReJmJG5
YFzZv/vwiCq17gvW258YQ04Abw6xM69+QBWl55KKaxOAyw8cR5w+ApUm6UBR1e/P
sZ150xHlLKfqfXQ+/bRU0isEBQV8NW9NYkPZ9BNKqSmvcJHUg+432dHOGBb8rpGu
hjW2F5O2t9fN/Ym9SizQalnmx4uj/+YUI3BvQlT2FfBSIYL17jBtWDF0E7LzSY7I
Ixmk4pKPbdBIyHdWD3ZivML8jsgC6yK/o9ZsUGrBTf0mOM2BydJE4o4VQtP2sioL
Z55uom934dp1129qPfM+Mqrq2gxJuDC5Dt2po7iclzX0HFobIr5PYdKthZLrC7Ba
Pt8RnyhJutDmWJ9s0aUZig8FvteSuqF8R6BoDEDn2a7VxyR4wcVgreyF83YNGiQr
+ALvhtHc7MIwX6e3nQChTN3gmS59zgWswfvghgEEwnxxuPowN4wk7cfPKTM34xjB
wJxjoEHa1U19i9YPf2ET/spAFd4+7Fzdhsxim3wWviqgKKymfXvHqn8ZNOhtEwDO
Mx/SI/agCdmCs1RK034QpavKTISzl7v6qjfjit48R04N6NCgmqpZHgeUlS9CrH8a
4Z1oi9c4GmaL5DzEeWgaC4Kywt/Zml57zLTjKTUydrTdR7BIAZhY0WjRNqBySAQu
qjgWkmAfBkmgWM745Y0W1tAhAq4+waxLL8u1lhYIjFP2orZX9uABKgDCGOJBRJD+
SbI6drDG1zlNaFb67N5lFNbXcsWxi6dlrh3i8SILqn+ui0d2+rfOXlL5dbIhHHNt
qYqybvRPOZ2AzcPyK2FwiLVkg74H36YQKlpj5K4TSFH17GmBhBvigvG5kZ0RFCI7
1PSby72Ty4AQVktcQoLNse8ZOw1e7Ze7pEex332tPpIhTO20mMYs/8kfsNSiROeL
C/rkaxnNxmxrrWH+NTSfW+7A1eGAXPssOnKe+JkDQQUyJHmGKS0nRIDvro2ihmaJ
1Uj6I5LZ+nT5n9wQRNFV74tN427U0rjAqtNR729tYHC5qWUY5vgBpGFb5grEttTO
k/Up4rpSV5htMMhv/BXrFvgZ95mN4EzKdI/WRJaIHfNH6i99rpukBxB+u7QzF8ws
O9Yj6ANTMEju/Oytu370UkSsL1TVSrkCulTRo5J+HuRZa2P+2ivhFDNCFGe+ovZZ
W3V8bKrV8RKKPmJJ/4gldIB4GKVOEYbferUUgfIuo62lK4mhVsbKsvlG5f8yBaq/
c7NSCPBnXLFoKuxBUYEhhBBUjY6iv+qLsaJVjEIZmFCoCQ1sjpTgexDN9wKQIvKB
j5Y+QDMymvDQstiuKvsBbC5sQhl6gAJ2Ps5kCOzAUcf3kSkTSzk/CUt3+m3uNLuU
B/eXm2ZbESmbVY6+7nmeX5MwXY+HoGc3WTvbJHiNP2+cd9UH662q7SYuSteh3jT6
Fiqx2cD/ro8KG4lna3kH7CeSNHmAkAfikmnt89qm1bj7aZNJKqxfO2gQl0hSUNpt
fZ1B8x7jG8hYdpGuCCMXXCTIxKrW/Ck/4Stu37T8W3HtsuK5euFONY3azOk+D6Tw
maCnEh5NaEjhGSwT5jVocqpHnBzBr0mXN/JUrDBRg1geo6CwYSyVEV6GXh/DcbZ8
K3bl8qnLcgR7TqRhxcDPItrRxP2hEdjI1raehvQUBN2lo516xoYWIg1KAIhUP4Vk
nzNibPoRKMmwgphTEG0nXgu+4Jxi0aJLfl4EOJ1ojoHmW+7rI8bsVfg6ZyaBE0iq
mWzrTaE3ztCf0KK8qvIlMMgxPwZH7+wbMb7QAwub2ctwbaMJNVF24u1SJIWgjt5x
TZqipLS682wt9/9SIz89tyyLl/92yQWUYYg6FmSnYRUZsQY01Cu8C09lQdtKTln1
Ra2dtxaQzdsN4L0jCKLgTpcT+zzc/PpeBIRx2pNhW9uCOcOMnd1dzvzMtMI9WuXH
H6eaTW/5cq6zVUDZQusCCQbZS4DvCgZyDCDkv+0vZoUBYmMjCDticz25Gr+U8PAb
UmJfuKKpfjd/uXDNnXHx+CNwj+NOMMhZ8Dw+NfNDSzfcRf+cNwxgPUp2gPV+Re7J
z6RiYsbJbCjHM27wJJVlneHfgLCDNUm0nm0v1ZXfCYcjgYiLNxZk7Y0RMcfM9YBj
kBRkepV8leJchXT6Xd6FemNR/X38uIvFCpdpco0Gnn6RugyMKOMyCkzdHBaBUWHd
HcMQNpGaHNPERttjIrHypXKbGtwNbb8+saDKosHcUMzxSv4p67jqul0MqQ0PsfLd
BEStz/0cipDHK+xc34H0Eb8R0gU+qqR2uCq5y0c/ZY6TAFBpw53AvVaiK9kz5QoY
Y1vZQi4YvACvHDLluF/EU92bMlNqfQXCmfLhH726vYhNhWfueewSAjVIxkkYsWiO
WtCV8vy4A1P21ZtU+8t+lpoBfnSDBVZ4IfQdSGwR7xcsc9Darle/OeJnyn0XW5QX
pDjZ3A/Ib8lYbY67jCMDadTQC2dHV7gdaTHNoZg5Q8fuX6sWaLCUVw1EjHUewhF2
ipr+ja9MVVcHBP3ncDTlD8DEqbqbXGHjCPJxrXOOKNjZ0k+QnkTUzjlX10Nc437s
cAojZ1SrpH9T1Y/0jBharzwYRgfJX5pGFayLO6SXP7I40vlWIWDkuAT/rpUZUfXL
cePBYOMg0MNRCEn2mJW6cN6cluBFegR1MynUTiqRArB6vamP5Z5cq/U7DZqY5Qig
T7mr8qFjGyAEfBjS5JXzgKGcNwUihK9sCvSzOTAcAlDSm/YXbk0CJnPBwzZU5iNX
0zyYZb0PUipYHKMWEGzy8LRUsTtbp6fYGM0BOO2N2MshcrYd+5joEtEqPegHAiDq
PhVjjwzS7eQ4+G0xc9I8vI/zLjZ82GQ2tFGM25OFtjZm2lpjcVgrfRWi/Vppr19a
98x6Rqf+1sFjQZpqWwh0EVyPeDAPwDXwQn8NraG0hHnB/IBbTLVwVJ4JZqWrGBVf
i+Kqtb9uex00At8IaJytfJ3QklWT6tkngoVCsiSl8Og56JO35zeZq8ptshL5I9Wa
JXNWThWZBpK0gih8DuPHDNzBDtF0/hWf1yLfF6kGKikRKMSW2wh5qeOUBPwZoeHx
W853LNGSCARtYerRHC60+2sYhNIrFpmnk0Gt3bA1EOgFkexgzfnkIvBm4Pumo70w
Qcq8D/PsDRw8RJ0SLLitcC7dToZFfM+XXpEI5Niev/VNDuh6Lf1GEqhodpVcjY43
Uh+T7qCChoximbqhz18keWZwlnmW+HHLIYwq3zmATjcaIg0vDkw668EPQZHkOFmK
vAQqGyezlJhRggZJekVaVMShQqquOj92w1CDXDBhtwg9jfj1UxUYZG6P5vSJU2sr
IV2QFmEMa/VT/OshhqLBcwQLHWwfslwUrDllN8SnJhiO2Gox+LtXfxipdNFAKll7
YGMU6Sii2o0qSiS+7FQ6DOKETtFp+/a5QfSO/5jzri0nFjJlARSzzaiex0Ys6c/K
iWo50fLM+t9CxzQT/d97Rs8I5dszckfeS+m9Xq7JxR+bQJ7VGKqWm3/iE1xFCHKB
dL/iz1oKJ99giPt6TF2vGHWBgzoCHq35kHGekBMgUD66OG6gFQKQTLGFMAE7OliG
hKKEXnpKKzPXPn/328ugKdCdnBULw1OPYUQlgaBPCW7Bk7KLhXkayQtT3+ah6Ga6
Kgcz2YCBEhLSA3rFQd8dY+MU2nsWOzlayrSJ15HlCOWJledCe+1KNfVyIdibOPKB
hwm4PwFxhRGWUfjvGdmhLvs9wFzjpFFgJ1SJU3xAGk6pBCak5vWvbAb0G4UMpQLW
UunhveVzPpuuUbp/93OmnltL9CAbmptx/ekkhAJloro9N3utoyrfnwCBV0claTm3
G5od/dCpGd0wrlbvgXmQUZTT3DBXbBdw/ZTwknV2nYuAusFpe3o+Xksd19FIOB/D
J+sIkHmqAv8Nae+b2PkKgV/ZEBK6NXmi4ncFdgUJ0PGOlq7EDzhHmWbxTEAoXW1/
n0KpxcEs4KPDgM45/6F7Bdwn0OqfSpko8JH5F13DwlymqaH9vzaXTeTn61kbqHiK
iV4tKYpYSCSS4++eCVXjHJhgA+PU3j+kHGjJFwttymnzxFLvTCDj2O8KkTCj/+5w
zPSkuLF5+7Cr0UtYAEhJLLnuI/0gASa/eTsDrtQWERi0nqlm9d2K2UVcS4YOihoS
7aS3YijjojfUq8jiUp8e/TW6casTlJfFUJo5RkieEISVQFUwLXoO9GxX457KOb0B
FMzqzem6H2bkepm3yZISyzkAbDkxjs6kFBI0tcoS0inBTzFolbYG29B51PxHBQUb
RJyes4G7i/XnnDmLYBTirJZTMH2Q5lyzwmbauSy6doPsxFDN58ijt07dwqwJu98Z
emuJkrpBOSvzuhUQUOgBl55EYb0JxLZF7CKLDmoL+Vvf81JnyVxRwOhlXcXun/On
0pB5/HLXVKezPL7azo3kUV45H/yTLYW3LPXR3bP/vN9J5MBoFtyPCc0FaOCNae61
1C+lmXmwxiuCYUgA+2vZGqELgXYtbcuo7gtaKH5yG6vU/PnpGrJX9x2jjfODtFfu
MSyW/3bP+YycLx2hWl7k7XcBxctbMZYVV7JQGsMVuYMRx+ldGq5QAEM570ND3GGc
xG+e9jckTmfRqk4tkLE5JyKFg4ntg33m560A1LkZwbILCuV7JqUr2x4jFA9Hckto
8LEfQqc2bE4gf/2+O0vk9MA5rFHaRvjdxb/FrF/T0Yla+CRsaFoqBGLS3yKm0IyX
DsfZMUrVeyuolRmE2EmX72PF2zHktIGZsOb+4UTNS4P1hQ6rgajg0MlrY1waZI9Q
zn8zzi9/uCG4hFeXKfZWz5fBELLrDDBvkiVWK2Fuc2DMi2tz1qI3fYpuOHIqVok6
RFoISvk+PQTngS4QKuoK7ZADvHvuSNJUGxDMmwGV2KHThIIINzuVeDZ7gVpjq77a
ZkqX1eK1OTIr27kmqe3qSItFq1tsgPHxDhsYTasxO0OF4pcyWDqIocSudTEqbhbm
XDWsZvG8nLT4gYB9ii/NBUCtV4TMLtLLyi8ZmPB3FxGROu4Gw5M1FOzCIucANrrC
WewwAfdnJWCAqMqehYUvxfj/mVUGlqAl1UK/aDIQWpAtCch0OAN1OmueV8Xd0DqB
LF6td02JAWPoIAIpR6+NHpcByJ3AVzNGRZDHdt2XxrXLOV6CD2nT8lrT4rMDJAIz
mL3RfRC9WlLw6c3pmV5Drs3eiyHvSSgZOW4Lv+1qpAJ9Gn5e2ELfNdZLzaYPbOXF
8C6TkKSfMh7x1Ruh3Uiz/Gn0xGEaLyhpPxCTSJdG3aQJSA/Ppi5ar50UKG9gJHsg
7gEb8leiiCPhu63qjPdtuVaAM1bJKm6LVQ3pY3zvhDxU2sm04emuJdFTbcJqJ2uv
CKi09ApZbyA72fMOR5GozGhe6KwRg0ywq8os4cVhcI7Q9wLAnsDXs64YS7cK229C
1HbyYOt09zErdcppXiMMyOpfArCjctiQIVeG5nKK5ybhmKAE+Lw9nXvfZNvTs27A
GcZuAdffuL7cawmBk8MkJwb/Usj4SsU6NvR7FUJw61UVx6H02htyjD07iEMkF2d9
L/O4PzuLTB35mUrSKD5unYOCQr8LqDgg4VbIpd8PsJ4ugwNO5CHUX5uj/3qh0CTK
CJTDljrHUKRwXCXPabjYUSKOQwY1CP8AAoH/QPzeNintIaTXqcHgcpgXE2+De1oU
tBQpKThGT7qkRAJhDEFOoWt0EZDQBnFrdoRGDmlsGTR43Dl3nDa1NAUrtG9p4AvO
BdmQI3lMC/HEgFkkaSP942QWUhJDtngvBGziyIxN8lFKsIvaxtjMeR5tLkoUyYq9
Pa2n8gW6lxIR2AQsaHupP73z+M8U59uy38JP60QNO2xeKPyDDOhcAMHrtC1PSz8m
ETRuSVVSHBsnfyrVMzl2ZaWHnOBiX9MwUI7DlT+UJrl6xa6d2oqiurIyC6Xo+q9l
rvnJkyY9RSLHoO7rdkI8q9/OEnFCQ5g/qfsX4SyMHeCqgaX9jNvOjPO9IAA0vq5u
1HW4Pon6PB73wxSnuAfWJU1NcSqlHnmupkfdjCY19TJK8E9ZKvvb2P39m79Hdzu4
E7X2NDwg+y4LiA/F/DnHeBpIUHiyNusyhH8iGUchGCxMuQfgLfuiIxqt0iAOZCsw
y/zDyQMxu+sZpzRWf9MAc6Td2ek66s/mbHtvbPXSTJB2sIJ2odaDmfF5KbGmaKVr
Mpw+hfM89CoYy+03uckV4dAwyoskAdFH6f7+qx7u5y5GgWbketPUz1r4nemejvnH
yiCWkQfoVMvg5TVN5t/95no43ga4PR9yzEMC7U+UkFcVQ41+47l4q/3sKa20xaim
6dr0uRWtYPwWnVmKhk7r8X1tBcGnmz0lekFF0UMYusfkIM4sWqB8q0S2mF4FyhaN
20seUEwp3810sWnN/Qr1hSt8Pmr7D9bmDdIY7JX3UQNijJjwUnsq09oh7EzGEU6u
PWZ+Gt2YwEPt0texGUya5KcEsJaDZFisgkJxE3qHrGt91tthod+dUtl8dnlpfznl
8xCsbWYBj0qy2IckkIw6p9FQ5OZYOYRVIz+hl5tgDd3Z6kFGNf8ZBJ7Ij1oV4G+j
VByp9uj/vXlXt9u3Xsrig6RPholqeeZo67tUZ/PhQYSOyT1RPLlGRmaz3R6BzCEG
P/SQz2f34WTvPBXh41QdA+U2C9rms6MWEYSxIwsVcOOwl22s37i84Nbgic2F4lAj
F7YVrrzfDEGHFrlzONj80ESZe6oucInbXQrFj5CyAz5ZIA9fanf6avZ6YGy521S0
DymlKP4LEY0UdyLURJ/Dj7ujLYJQ6Kivs+DSJx+976LeRa+VBb9nOs71XM18v1HH
UElr6S3LP66lYesrBZ46Vs5ardYuvJte2gSUDonjF3GnwhczJRKecVN4y0EYjPIG
UAmD76rBMTzmO/LnFL1VAAuaV09tvL4DHv5LyoC7ZBQqywpwlu26CVm/AgUkfgBM
KWlVTkCCRhculuMc+l1zW0wvG2EMzGgZvhjHZ6pOlb0pherV8Wu2iRLu71NxANCY
wMdothUiFWNo3lApRVPWNtNl7Yumyt21R4eJXMjzD0p2/wp37NTpw3OQHfnz5u7R
QnkQw0qDippR0SbM4tsVx7SxQD3r+n1LscM71duTwM4YLL7g7rBhPdIQeYIdGt2m
bMSjUdYi6qLN+sPyyN5R84ZBshfY3qVzMuy1XOoxn1Is4n7+OPlwcIGKnx5pjd2O
f/yxO0Zis3gij0F5maK6DC+Uc4iEFPI4cKAIWIAPkdzclvuKfpFHJUoX4Z2WszTN
Liw//FCz6TqqtwKYmkRcsc5v76cxFxPRD65hf3tc7iZzk3fL40hlp+eUynMOzj75
AsUVLTJbWO6xE1DiSCQzIFfJQuH53Yz2jlkkR33Z51Arr8KtAtqDwkUcrM3JNGYJ
19WwnPzhA4yo/Wzn3abEQIzq6Dtu50/Oc7oTlG+9TywgTkFfs0CM4IdueroNmgPJ
bj/+4gzv5IJ6iqf1Z75uZLSsH4TjhW+G0u2rDuqC1s72c8qtCjQKLy/j1oSCXQba
RrWyILneMsMM3bTRxP9FjASeb7qXfNopaIZ+eBzkhe38T+kCv+754ceTCozLFZM+
2eLg1+lSSMIqDqzgKM/XBzYtcdARuCfnCO6c8Q7S+Yaj1bkjxW5YH1fLGkp3UAQ0
Zkl7SRAIr7hl/mH5BeXUxuC5+pB/HmC8WyZmTLs1JxLCCqgHbqFPcEainK0L6sbf
pfMm8X3PuEXWrf5Xh53PR5GmhpQHE+4lGT44Q/NQ3muC5Lgix5qfocrCS2oc14up
KSUxix/lg3fI9Vro2vO340LXzWkvj9fgkmDrgL35wKV/qSfKEfZ6vmrtGnTJG3Kv
lZnGBzppT7/WxaUBR2BvPvAGUprdTFCfR1lJBvb7c4mgTY00tAYfll5EEqR+V+kb
cX4VtePsb+rIcDMUwtBeODEu0SfgVc8AaCm4r/ibxgoLWUbjS7tGblhwp+A5VnJJ
F22wTmuhchk/D0r0PTr1W+1NlcGuXSX5X2Jj/JGKA0/VpSouyesDGVSmwLqj3tcp
Pc5HsEMlFliVv5BAK40l6Cnsq/MUZoV0kzo6sL1wQJGU5ahK7cRMkC91+F8oOj1q
PG3dIw4tBDZVUe0+w2zRvf2NU6b3n7ZmjdNUwXVzi8Ld1JsrN1Afaro9gfsBfVgl
LHU2HDveu9mr+/XoHowyeER6EG3W0lUNoTU2SDAwD9Rr3oUc3jGot4smm14kn6F9
wxjn50hRzk+xwm2HsgKIRK1ECIx/Xs1YxMjibKKGELZWBebPgZHFU2DNs1WrioIB
jh1BNGDX7FVhNQc3cjSl+5uF+Oi1BrJZGEB+8eI1nIQhyacLt6ggsOXotZYEgirC
fJpncjGhdQwbmCr20wloo7nB8CSfznVkGTfg8qZnaMREgmN6VjA6Nj1IiPWJdIfP
kJd4kx/Gb2L+f4cgEAFVsuKx6XHayk5ra4vyguvQvHm75UHe43kVTyhBcBUXgVXE
k5M1fYv3GExBSvHw6vU4fSAM2wi7MRxr4LjAvHRiKxKNDtlB8dvVOwNo08XVcto9
dWpePvwp4s4CH/rDLsO4ScRCjdA4a/TIdhgXA9dBQ65NenYhmte5BmdOxCEXOGzw
9Zoqx0WzDPGgOBIm/pYQ7CEig70J9mIq6a4lkhvABNV+BjvEaRwKxhP5pCdqiLjZ
VsOiJE7u9d+uGkeugEahwzvEbRbKU1Qk2VSw0NkJOdNJs9r8QgBJ2WR7DdDPsWjx
CMWIq5A/81FFf5sunKWWrtcoON1M4hOv4yJmCVJ2XudFJSv6WnxsSH6X17yd/v6E
QL8Ci4TK6TpruhP5mOHqfGiG+H0cPKsVwoFH5qkRw7F/slmgt2NZqurypHASFv87
wb2dyAkqCAEaxha9LDOwYPAnukXw7CcRMtkNFi0PIhhUZHLMVaJ4UYV9N7KNEpak
DXsgvroCZ7MKxWmeKB2nD702sbbBt2ciNofGhXTIWSHr1Re9Xgq8nLyouKA0omf+
T++IDuJqf6cQwHm15wk71d9/lps8gfYi8Ga8Qf3mWuMDM64Qso90RC0s1K9a525C
Hoe6NbC++FuJM6xoM+f5RhpxFQxUmZOoOFYML2QT6Twt53INyAfzGhzuskp/2FQd
/idKD5g86EYtMtVaKAVKtYvVgzlBVHQlpqVTRVkg4ow1TsbVAQxjFoDvnmXy22FZ
0B07uMYJRhOUSx8qNXHP+Q==
`protect END_PROTECTED
