`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PGuvBuFJUM3Fy9mwk18lfCgADi2oFYVnDq9Cs3nuSN0oKzwWIjKAsFfL2zoTIRFN
TEwhNz7CJGZUJ9dX5LiTXr5zD9IHXKQ1odjUvfod+5CZjdXism7Psil4KqpcQfvE
hELvDytK/0IGIr6CR6qsWSIizwrGdlXlLQ5NSdrzZUhe7TyvGQyAWMtmNojmckLW
tQjTAq+rQHzl4ORkUaEVPBwWZCq7XfqVFll7w+0y10eJ3qo3BmZGaj09tHMKKvgQ
tbuKNkRy0rj+Zbq14Gn6qbUyo6PWBqUnrVOBJ5IvYFlAKwmFR7EDgxg3MNTdKHwO
BJNUCdOJecDDKMJQ7CmysOkF/kEtgPG49fyYr275CrmWuDYBvsadL0WXB2B65V7k
jOrRyEnrCu5qN/CDwgMVQs++jPyV/YkzVskJvSgn5dRh129ZVU9KqZPusaCUWcQK
0r2VfRyYthMPuTyTvctTgNyjhGYlQR0C9i0FR7SnBSyDs/z/E5R4GfjeOKUMP9gm
3AKb8JTwc4PR4cG4carf//Dbevs2zZUTyPw0w0sHLzSR7TjEqp468tcPnWYFVhg8
egl2YYHBvhOyV8EeFeszTZ2FxyBrPrgfA+e1fwJGI62PYVuy7XSyzmeLFNViiksr
lxehyFTwAjYhSlbV83mEAuOiDo2gFTr3SKG5xws+U7kLHFB/v6UkDGYhR/ISTANH
svcy37nYmE/q7RtF1R5n/yCP9//p4hD+iOy+nOSuJD16C2mF6A5iryKfLUvt6Y15
8jPrRPg613xXuguiR5VscXxipAL6Dvxi8rs8Bonl5RIYubrgOSqf4Hts25g2JPzU
KqBKDoyRx0vvn01bE60+MaNfOpR9qacntFViE53v7pYqVWjJY3M12tJNrZ3Nab02
EQuhY6ejvnTjXVglQUZHNNR1E5yTbwg4SZxbFDCbYEy1UZQQFqxBedlK4GWwM/9j
bousiN6hivKWQ45g3pg1o8z1+l7oNo0ud4jZKO0UhTx/iyF5dMyIkPuIO1jDAYXJ
QnHEWXxNteSwvbt/AT8GiZy15fra42mEfG3N/XgvOWANX+FE5UMOXsb22EUEeb4/
Wx43IC6u0lQRldQgRPhzkriQWAzbdIVfer1RjW4T+oAL9+eq9cpqX9c0WksdyPdp
uRj895oLpDmWwLjKPTECIWGOTEm6QZ0d4l17YqeqF6JmHORksXhjVS/KcIyE/vT1
19fj8UURJmgKsdOE+w8Hdfq0pqLwmtB62cQzbIOV9AHj/LWwBVoTAyFd1kQLltBI
2DavBsCVxK7OWy7huH2fjxdkUEcILZEUAwu264mbJUoe0cjwKlKvahrjaFCx2ZiT
wjF3dVDPndge16Sex12au+em6ooQPcrGQdkV+APY9a+PDEfGwdXkjAwEr95WF6lE
2rqd/baJt+rUQzsDftNGD+4RQFRznAaI5jeO88wmInwX/d/p/XsQf3BC15eGRJlT
9Xkl4T/kz9nAXBXO7BA9vRJXReFcHI4rcXsVmxJMnoCKx5XdmlUJgCW2/5DLZr64
1RW80cX6DclEh6ME8BoBZh2lL6q/D2hWUmACFC5gSX35H6++POYbOLpDAlkHnrgY
2EGegGaSAZ3cqs8K5TVTKI98Yy1KwmkVdHKtw45RPIXhbANAkeiAaQJqrTSpzGdJ
ZET3z2orX6jRHQkB6eqgdZLsenIwrxcnyIedh9FTXf7uqFMlHefUMFwWm/aC0y9Z
hWm5Fqb41LbvvcPzRltymDwAng+PK9RzqegF/yQjfTC4Ks6lEiWHuoYb3bFqCYnB
PxoxJM7oHBiXI5zid6hm/VkqElfQHNis3vYsXcUcW6Q2Ap+jKh4KESM0Scq+JneL
BqGiW+Y0xo+vaaAjalVEYZluliixhje8c6UYFgd/zF4i20bbcLlWmNmuPH+ec22U
hXorZ0TNLyIOVN6czbyx4F1Q0fDEOfOXRVHXwle/z9fiP+eNewDBmL+dl24q53VE
UsY6+DjLLIIkZUJ39W0YUWarPXR037Lp92vc6qRCpzlSqqtsGDi/QRoO1pN/kX4v
VnNs7RQ4J/VfoppQcMRrGNwwvjBJZtjGeoIgzwhBRXYOmPuPE1KEiEpDh1WX19H7
oxMLqPWOrhwC1kR6VzOPBcj2C/sdGY45OQxVaia60f/vO0WXYEmsYDBRCcgRpRFv
bpbQRkHZB5DKMslNz8HY8KvcVTZW0nMI16kbunsEGZW9nu3RlhV8NOEcUS4zm99m
l6PPIzRth+fOOWlDgTj15TyVxqpMFYULXEHoZKonMX7CvfE8t6LHKG8EqJCrwjMW
ifh/GQ57rZ0DNFH1RJ7zio1HcqXRz308sqJ6sZF0b1JOGwvoEkt6IaM1jNZSvEje
RO4UHHZ+gNfw5tvhLoalYSu8BtbSH+nrsZHcvZlbO0Ki64ZfFVyDRkGsXVWjiIp2
MYLLOdhUJOIEHAyC/NxBTq+w7qv8ZucvcbnDqgEE18+7h8LKXH6jSI7B3+Hjj9fy
8uQ+uoeijZ/pJ6BRtNn6HN0xHYDA2rKJiSSoaRpTP8Ta8i/Xbsdpsd4G/Dhltdco
6xaA37xGUBg3/MLn6XzPfEIXspCSPxGr5R3LfkKQVAWBvCmAWZJUJ4etZRRGLj9r
AyoYaA74dKYEZm/sPj8DH8rStJ5lNUTFkA/enmv1mq6xqNhHZUrmiNmquK1h5JD0
A9Mp/t5mEbP6kmVyq6g++ubml2Twvwq4SGcGlbJoCGMjLQ1eHUrNGsVo96KrAVPu
g5xJGCqRA+wwBVUKxlnn5Il1StZ34joz629AUy6WpBSxpPEDtFNZ9VEpaDo56fzK
261UTkNLejX80zmTlpWyzgRgzF1blsYsPb3wmoqdAKy60Q5ewtXGxPOjK13nQBUn
c5LXT55p0g5a0iroMpxouHeuCThz4nmnZhw1Nz+LEb8vaidJZCUhQcYM6sdBC/CC
1tXAfi0yZexfZiQxw4Gc680QWag2oKbprcyhS2iuyBDYITVj5oLOVl89RDnVMCss
XXyNpLB8HKK6HivBRWKOtMxTiGZ4Xv7HGXQ16xA6/iI331uO9O9oSDJYEaqmdr1T
ab23xgjt7v/uZiV74z3NQcJwyd7CZevjQ6GBHBlc2uL42Mf3fvzHdabssU9h1Emt
MB7s/OMWo6PZPw8F10VfK+uJzga/KR/lGMT7dgThrnrhErmZwi1zAKCZsi7s/+jh
fGDFCp3XoLd6mPjcEirDrtYwrGJ3ETnZvVeEMPQK8p6oXJcNv33Hx7kUSM7tMXYf
pZzKeBD0QUyr/YmO69uO1yuU42JIO86kK1BkFNrE3uyxo9IKBTsmNXb5oFJp990D
Zk9DHfGEc+h0sB1OZTshg79N7WUmPSImYhMeG+3QBwTVLqkTNshhCJhyx8S2hVrA
2K8ihoxLkp2csSRbUg6UqvWtIb7oyEt/RIfXqXmOWGdQ8mb/H3AyKsa69/A5HIEA
QCzKrgmfXBDI5Hj8O2AFJLtlujz93jz5cceqP6up+VY+qoQ0umcFILSkW4N28pGx
NAWw+v6ECrbkJt/Aa8GZrPMJz+CmGE/0PU8k73kukSgxeb7SKPUV2kTmENgd99JH
A5hBSwJxZ4l4U0w/4KBIE5GtOE15GU64IXzxxPBgLyQPerZ78b5yTBR5tHJvtTbq
`protect END_PROTECTED
