`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RDjW1sOlEf+Dp2ti3Go91FBi1rSOHU1WZOebo0BMRmFHv/FjzfTwcDU/2TI8ZaSi
EjxUzWJPxYgF5LFz4NEW2zgQeOikEDYQPT4a4NOL76GzYDr4bRow0bs6qn2dIu0Q
TtU9kbH3sdxg1vvtMcga4KgV+9+IU+ClPeeNA3VUooN1y7Zh3uH+w6kAqVNck2Rb
5MlvH/6nswMSXovS6wR/bYJephQggwQWOvY9tW0tYOC+uagU3dhlf1mnLAmZ9SRR
55BZLkXai+98G1fKXqIEwaH3uARXQjG4pqaEKm5upQyXCGy53IX6JBgWhhZH/SIt
hlIZlr5AicurjZ/3Tm4uymHoFM9HgBuM7LG0yGUlx3Zu2DqGxDOwZ4cgPvYga6OH
M7sL77jCVudEfHd3gJ6uvJNc+H440xjBGUlTCB+EqFt6R9lqGXN0t7JG1Eex9f5J
4R9tZcL4m8twcH7SzySKeBl6sFcJOh+/m5ql/kqVHz6LDahyztHKx0y0fWBJmUvO
eqNNHut7KH6JDGCXSVE3rfBAIh4eAKzkXTA7K7nj37WfZRitqGXUlMw17C8z+ZeI
zF8C6W1xAVA8hdp45SktM7tugGAEjTq6TiYs0rBHyUZj/Fd+5kXQ9ChU276Zo4fX
`protect END_PROTECTED
