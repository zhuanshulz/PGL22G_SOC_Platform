`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BpL5JZHkzvKVypAmR9wNXQE1OKlLC+/DPSfXg57SSyR331a19UJo6rdjB/QE3aOo
7yIh543Iv/4H7WEbeiafWDz8VfWojprEC2/0FzbU859XNaVxm14t6afwiykm//C+
0UKjlcaWpiWSMyK5SNc1/ZGjkSuKWuoOzGrzhogZpEIjFSjOCJ9n2rTBnXa4gr5C
6gU81Jo576BetMIILNp/mhLsBC3OsVtzgiIydVwHzs6FHWcqDLrn2Vl/+6PHPgjD
Vr23rrFV3GuZ3tiFrVaLynaIdkfSTM7ck12NfbXnkwiCQgeDft5/ZVqZk49dvhSb
zQioJ7exXEgOFhcJogvYQLKA0BrdSjvuwSYKF2cXtyFcobDbEWZrBwUaSzcoXVqI
2o6hunpX0zShIqs0ZgIGH7Ko2hQgkDgabAJA/pWyngHft0UwFUN3OCwXt0uAH0yF
1FERykyeT27XDY5iiF4tfppD1kRjL3CA1CCqG8blW28QZ04saRVTzPTozN2nop6s
00ktR43M73zKduBrSBOAArQ+1p8lldeQ0N3edvzLm/Vx/JkEx9URfLXkXTP6HnWx
iO0lacIHJihFib1A8VIIo/AL7bCevdlX7fy2jn14AaFITFiTi4hFAVRoA/8T9z2S
g3t+dws7RvQaXwSLWVfKrtCge4y9RpeMQFpZoBN9lkhdK1xD6PHyNPWfD35YZ1sh
DpZMpGrlu1YO9ChoxGZOTzuQDbGErD8I3jw8jUbwrHK0i+l3QEsE8QPUq1IPgfrh
evk1rOu+aYRJhSe2wQZ2HvG+7BClrUwCqaXyYTV/bQvx9BZ8Co2qnB46OeqW6pTt
T/pw20c0secXRf3R4bIipPNq/Lf8rs6ySbiPUIql+Npwybk3kF3c9DvHBK8eIRZi
KJdQGxMCfm8EY7HWU9A6IzoriXN39fKmsn90AZslgu8=
`protect END_PROTECTED
