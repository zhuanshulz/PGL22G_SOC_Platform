`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/hMl8n14S6PxXZAB2b6nU2Ud7jKoL4Ct0fa6Es7EPK3oJsM+c1EyHnH+yo0HdJD4
EOiqVJq81FvOV2tdJ5eWNOB8waac5vrCglg11bObmlphHizY02SHZY1R67JGYot0
p5J3mEAADpLDf36Z0/pQMqJMwHJfFMf4zaxONHKMSij2LbHFtJGMALNeOIK1g513
eJvYOQqbpvrbrUK1ad7ZFf2ZWvepOBOePZUr8+K6aZjlq6D/Qc0J2y9Q2CMtzrpR
sBlelwMq3jyLlQGCzKZe0drh1p706urc40UTzif8TnX+P1WVa48N4cnPHYI3mZJT
66pBsa5cOVltJSvb0KBHjhNShByrKoxFUqXOyp1dTwz1HFIzizyYpqQGAbOuj9DQ
zEWeYosolssyYPJrHOHozDe1rAPLfBiQSGd2goBOQEp6Xym9Fc/Y1hMOFuMoJVWw
zPJ2tt1RQKzBOCYV5rEwMHNFMWFGMXpH8wHVGP8GEjorcvppRXpq7zEfElLU/ELy
kVHQWKn22vGVzAa0TAoE752n2Zj+nU9tLgnh5wrtL4Ds0teE0Hp2tnN4VsDqLNcW
AsrLb8uch9v5T3jFQC7MCHtwyE6umgndW8GmKGy+PjYQDFcka3/qbeHghSOeEmRD
idvoHDk1rClzfB1l2wLJiA==
`protect END_PROTECTED
