`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7Ayp46hMcCEsd35vPOlCrs8JufKTMDT7vX0kq7Soe3zsrhwwcCfV1CG8Vkqpvslj
GoLY8hq9iVfeMOi92E2XIxHEQkr28BO/fY+i3nSr/QoRHubi80ezGJGggDWhIOfO
s+4ngrTbPPkLByZ8V92SY6PxkVau3N+n/knmf/GFzMjpdIxmJt5iRpHmjedx/J6F
8csVC69s9LmF16LQCaTsDWcEfm8yK0BREyDLuSWLk6+ExTmgsvnI+TNVf74WquP9
JEm4Gu0oeGF38emcpTxE/sfR1OI8HtyUW2kzXe/LKnfmz5Nkp4Brb3pthM7bjfZ+
Fcfmax6dAFIQ3+MJcw3tlzv0jKlJlcLOabVsnF0k9gQBEB5bI9Qwi0Q2Iiagr++I
riWa/9B7MN0BXujUIlya3ngImSVMWEkbloUdbhV1r/DPVD3fKmLd7/8GAK7ag6I6
ffahOCYT72gpvj25AelUe6BAcdQGsDbJwjw2g3oaw/b2PfheGaFVVriLbpW61lfD
2miSsjbkj65Cout1D++iELIk8fO6ZM325Pk9YowFmRDofv0N/GHi3FU4+b3RFNXI
+5R0Kg1kmT0b0Azs7s0LrPkPgshzKQ8YeiN9p7FlwcQFjtnEK5SgqU2UOCOgNUMz
7iRRgX9ZnzgsYqiFLDPGIrc1TE2v1loECwRMKrLCBO/lgExbZNKw+tT4vdGUXNth
U+BSQOyVJzQ/aeGjBvEXdkXdeEYTQwKcQ9q8Gj0XI2+qsnWUAq+TnMtejaQXbDV4
AbsZZsics5TmNo8P0eO3c2MtKqH7jgU+833eS07k5ZFILJjceonGcNvuI/MeccuB
YX+PZm66Ix9aOFBXpOjR6ZR7YPO9GycuJRplbqgeaJVasdVbBKhQJmORUMntmJCY
nBCHX3YhNFRxAuH4rxgvUs4bQS2gq2deW7A5MCplgc/Tu8qIREEkzp5lYE3ENy6L
Bcb3d7Sq3pb/mI09I9TtMjzI2JxelH2YVRerLnikFwy88dvc9wi37LsTKYk23syS
V1z0cpFWkQTawwybwZgqhF49Nnkb4AW9Z2t2ER6xm+PpXOXgcmK+Fr56UdrW9AOQ
8dekPy+ez0YcHooKvD1FC5HllIyh///0OjPno+2Xdseifxd3XQadj4tQ330nLa9W
uf4Uq87vALb2WpbrIJNNTlHOp4bj2NCDfeRGGKuYSqPeSNGKqQr5uFXUfk6VbGKE
MSZG9LcyI8fMuH7ujiMFDxiHt2m/7kjhx1LbVjFmkTOWH5qXHrrZlgYnFYssKbDQ
bb2jIfINXeJe/UhiqrhenqQ6naNhR4bSNnkEI12grFDyZGXmmRNQeSSVCHOirppl
8SvPRYgvvhw5hhXkyyn0I4cxEsiRIX8jgGMnXQwWAAU7YAWlLZmCZ9EWtWWd+qUu
x6FuOkItd7GuZdy5JS2xM/53RigcoDSqxsmmpRPTE5pPSxFT2gFHijBKS34IMDar
U9aM0dzMTdByL2S6c/Kj+oRSlgxAvTx8qUsAs5nzm3LFXGVByicl3CG2FOHV1+Hp
gWpbfB5YKxbgI1dc0L8juG+Zpb02gNB14f4OvJs28/xQ1PRzmVbE47Zb26kqKIyB
LLcmZXaaUcs47MgwyODS1lJcgXp35tVA7j5AwxfG60fLEHT314Bs6AVIArD8xeAi
JHF4gY80Q9SbTLQiNhfRb6XAnZcmpilK2BPB+Df+DP3jH7G7s32S4x5PFHQ+rgwH
`protect END_PROTECTED
