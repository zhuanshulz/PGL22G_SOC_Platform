`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WMfm4B2CaZD00GvzkD//U9qTdVPtTXAWCpm3t9EeU95kXmQZqmFRCa2wLaI3+pn9
OQbOw4Npj8sxlsDo4CI93X+66Clp2M1BnjjQx3iPl50UbfGN4m5H74quptIC6bSP
tM2AySmGp4BOUjmWfXwZZMPAJAmq4OQ7iHovPbAuKBmw+o+2nKQZ8jdJ78OPb0qb
tYc7Q1z9TMQBNob3GulO4CqPUaC/st9VwWWlzzgcYgvfCbUrBz24qItMRmyLBG6D
CB7qKnFLFbk1BV587lPZH1H03EiF5hgntVITrrguorHNl3i8a0kzlbT5HSAUC5s3
cAfQ+1kO2zfNQiE/Xvv4loya+120Vz2gq4KeVMvqfPWVL/l8A4hE1pylyhQ+UGRq
il1Hze5IXx+qhgZM8Zw1J/Gbx9ryN+PjjcDKxiiocdalkKt9aTb9dOG6d9j8yO5y
Qx1Cgufn34dLJqj6DMI2dxbxgmX2B422xEhwsLwZewuRoWzgynO1M5X6bcuc7hKw
fged68YqbXerkFBBdcclA1FA1guOop4cCjvMdJBbpXYLTccmmzEYGMZzekGCQqSj
IOFTI+sNYYx8U9eXYTq4+6s+O6OrgIrGQTMVdECTRg77PiHbeohKcXSssBCWtEcf
s4as3VcvnQ8YXqJ2o9U49UuO1uA8ziiT84kTPARTnMqS+uIOx8HTLesUgea8/+Qk
+6MfHtAeNGxiEpJatCtnCdOrKccXw2ZSpnidWASioSAbB7afAnXwuHW9fX7AbcA9
qfVNf1fzhiQ4oWU+PRISVDsUEHe6Rep+eAtK0eAHtkNq5baTUJFpY4gbxCt6t00L
v8jTgDoGIbrh2ucB+HTmjQ==
`protect END_PROTECTED
