`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OTqni1MdKgMoakX4yYRpwkPd7a53jwxChIrAEu41PjL7FNgFZYvTV8SrpIy3x8qW
GDo4CqdfGjdzQf0qIYn8ATHRHs8iCxzNH6Idl7bGeP/21uW5VPYpvvkZs4dfA/KD
Wpjt6yMBeWcYpm0d30K2gIbIXha4Y+sY9R5Qj9MpPPbg1+2w+3a45WJG8ANUh/52
CUUQXZncTsf2Ye+uS13DHEktKr6Lp7rwdXuXDmIjN3ziQ3qjhIbY94BsC85+QhLx
2VYPr5bnQfclOcKzP6uz2C20u2T8O0PolXdzXEqd7wWnxv4fWnOHWTyOIl4xzK3B
JB1uTaA6Xx+i/pqVanN1mOZXtA7rqLq7Gi5c0U/vDn0iLvvI7Hn+DHPmWiQol6rU
rywzwITwmuchAswW4f5lSkCzmEAFhKOSN6A1zvpv4AwLfCykpxlXQg9362DlpkS6
q0ZkKi9rpRMJB+tKkpEkJGMS6dW+u4ufixrnf2PJnHRGbOZlEGi5ng0csHNElL60
4ZIgv4nqTQkWMhvysijtizLhQ3IFAFgP3BTH/mV0mNbi2wSAzKmdHa8ToXlmVxsJ
1XCnMXTIM1xlTWShJBTjkyajJoUQzeolZ2rG32jMMcPDXF64/sQQpHCQWb/GihbD
mgMq0hx16RXHTxkhY8GVF0n9yOeGQEyDyWakijtY7/iNC+KvMtA7o9v8OWqI9Zdw
w9QpfsGnYz3Osqz3bGQ5zFyLZHUIx89E8KLgSo9gN3h4seTJ6VYbVuWiK0gv368b
rmRXRTwugKZEA28/8EnoyxH527ycG7iwX4lxNT18EfUE5HBOaCEEt/dCzh4f0hiV
WRvDxITU34yPQXXNhukeIMlEhPaJFYt3hfneKn8hFmnxtxJsHX8Jj/I/Mx3d3aAi
n/N4XR8alM024iZKtc85R+zFpmsrMndzI0uyBRQ3RbFxlOInWI5td8CVli9pI/8/
fVNdyT5ARLJv/ETL/VoRUZkDIF0zTpFQOGOd0zKXH2AujcZTOWlUf3iikC+8PFZV
DyZqvU2G2IQaR5iOZgIhLLIv/N1jWNiluqyAa61fAscwv9vE9P9qv/IG7qiMHTa0
Va6aFzAKv8JTR06Ffag7sS9ZQC2BrXcey4/q3ePMo/kfF/jAg/6qRjVugfPA29MK
3DvmxcKsGAv46XVF2cgladcuVE+gr8nOxBOu5/kJ3EWJg3BdFiXMT9U7sDQeNFOx
IrugX3b+w1ypgl5xQW5zwVPbuLWoaG1Zw+K01gNsI35xhbrL3jceqDwVrcfiBXAX
G62+eVQc10MoKTKcu2FLtawOdxXaKfXCj37hAjvvI+h6xoN/ThX+eE2FjTrfiE3+
e9KRhqgLET99CHrIzpNdkhuAxUmXsQC4b4TBIvtkjj/e9wI1+vXVTL+Nw7lxHRVc
AUteEFZiBJ9QfiZ76x8SbBmbAZEjWhLEjgnfIDG2Vfye31oqPhTpNSl1BEn4Mnc3
E/jGu2GZy6wyG/jLTd+3nfaiVKYoVBmTYfAWbGTp9XVBJVjpDfNBWqdliBaH4Qll
QWoqS8zy/SCjYB7NozK1vzhRaagMWvjEQ4tzV5ol6YFSNqK9/VRSR8/AYt/od4CA
EocUUi5MGCxk7dVRFtpxOovqyueLnaZXKJifONXfTzsnXeM87ymQdvdgnA60Cfp8
RYWcKjaHXTbhQK90l/mcBrdpyfCnKQ+CwcTTTXrs7yYECNArI5rM3jZus8qT3+Ux
SCRpH1dpFlBIH36aZ5ufdhb78wCsKrGozx7g30GvWexAGW7Dhf/Lgopr4TNWg0n2
ysyNlb25eirJqGk2+WQ/a7iESwd8mpKkdyWt78HmKKGD31H2RX/8yfQFgn52MTHZ
31pt1WPzfAclAAUIvvKJz8reVtepQCcnK5nQe78YbkxDQVma0ZdScOEIneLPFTwh
VG+lU5+WB0Dyr1UZBeVBBv2Ow3Tv42o7BdmHGMOv2IN886vxzOg63fmSmq3OoWci
uvjArrDwXBkwt64JVares1Yie/D0aKoZjRIoGm8msEmY2bHvw0x3TVcoKruVsezL
RgjSYVKjjKF/vQh67OY/ErwO/FXYADeQkpvDlBpEuUjLRkkYIPGzsXOhZ7Vj+owu
EDqAX7AVTzpUU0pWggkGrwO7mq9x01Dr67BAMZMzNMnsVi+CPj/lBAzin5O0r+lT
a9M4S2O/Z2tt/L9TSPgYCn2ECFKFprDqFh64gmnqrT4XtA1ZwVpAU2Om2Q9aAI31
QujxrqKUru1Jx7uqB1jT2bSIh69BDvMVvIfMv6pXtiZGGvvhtF5NuBBX1n6NMNTz
ZDY+bW/RBUaVEALPnqtf5QWuj9mrBJJuY2+sbKd0uCDiGMSO2wj3tpCed3snfrRa
2K4Q3KLthaFpbHX/oGlGZRpblsnnSgRDjPh8TD2cZZGLAYBe3+aEvrpIWmNFmYuo
nqO4BeltEHMyjoeIPhJiXltyQ5nS9Js5GpRgLBhv6Sg9EJ2GGLCdcdbnN4PLNuPS
eJNe52WUNl0unRn0jpMJ0zrG7e0zjjePVXvhrtnEn1BLoIhZHRgp5yISeaoOuduW
qPBjqK82o59c5EYuOZ7VJq+hY/RbQsumgP5QjfuY7/h/se3uBmBKJjF3MR1Ag143
t/cLqruzd3/KicaSP6Xnfv79KakOZwL2FKU8SVWBL56LJ6nH+2Myxdi00Jo6OZDo
cN9bF39HF1yEYbg/AruSxa9nrkU+RyyWxHk9LuI0mgbg07Qpi9MctB3QW5PObety
Lsf5prphplMqzXz52eXKyKq/eXs6whQkIKd111OyPJHRuvkvtqVoebjWCNDHRvDy
RUngF8K/NR39hSGJr1EZhuzlRFH+nFFwwMrL2TPeuiwfBAy1Ilmh0J0feat3WggC
3xHRKGE3F3ieXrXfU+N7FKsz2neveEb5mhrliMcpKp8XUf6EshOUTBNGwXJfE9ey
mVMFDKR+rESEiagovtli8nI7mVQIyq6MXfC1UzQIO6+ovv9jN5ueIOCrfb4XqNrG
23VfhV7jSEyD7etEO2ywaoJK2CjHm36q6caVeV09JMqv9ugY7INfW0AmaDY7xvXN
QUt8EQ4bqqgQ2gRxfOy3Mmcw8gmMGTKnhWcl9QqeYjGDTc8I+N5N4CC52nhmMLiM
DqSyPJL7tl8ZThphgsq5AqxZ4bu/5VTePDw8x0Nb51IHA2G3/BG4V/yALVGPt560
tlAPE4LlYIFaBIBGoIQ1qFPHipCeSUn0FgcfCsmKdNGsfDQkOSuPsxqeM1BA7Jf5
+wTExBD8/AiCdBUGasYOcOA8VJ//9U6OUOfUqfangA1lzoe3AOzZR8Ras6WDexpC
9qk3Ijc4B4muf8+ZrFfVNFaGFZqqj3AK0VemRkg7qgcDzh5YpLFehNnuMoOMy4b2
pXk/KBRu//9ERr7D6O1z6KtG93t01xg1p87t2nlPnDfWpgPqnLPjZt11KC+4vwRH
rOu9R3tkG3ekclh5R1dCME3kNaHCEFtEH80UmOQim5OoSXv+ppGAMTG6PDyFyFuG
iz1rlkBwvrUzdo7dK8k/yMObCfmHHQpErQMI/M3UFY9wfDOjFFlGH/9UYiYaYzdT
NuN2tcjb3evDsFnUPvP5N8oHdVMwc2YQKXmNVkGPCQmsXtm8jIOGHzpAzF9dWCph
FIHu7odK+/7HeNHOIV6vAG9Gi5M3+VEtrcCQyym/6Dn1543bjKRsfleSxP6saCdH
ZmrdQYYAUIuUdBAI8+SNd7+K4+zoZx+J3kH1PPgjPwXsrnebFMZ0qAcAZGcdgvrw
Leq37edSvkFSzTLk/iAvpztZ1UOKfl9pJ0iSfLnu6Yfvosn4BvGSgzOwUobINVqv
JCjKi+R+oCLZipez6KxHuxiDJKSehUEzZAj3SWzeinIBJPLxyTiJpGTbkgrhzw5t
QaiTa9/YP2hunhPgWy1R4U+AnR/pbsSZjCXd/yXziBx+9UyEoo1faOSkCZQgqOM9
1BUBxXQoGxlKzH22mnHB+65dLYp99gF5N5I+HtBOPIgVaW1HWI61726kJyFtGbHu
v6NqKizrHoGBW85cCqMCHym68WBeC//fCADcfdc55nIrNaqOTZSu5KXIYzsZ3TtI
lvffl6xUinrLnl8Qbw0kQoxKNeAmcn6ARgmmYfyO87+kmBOt/54AQmBafAOoX+wu
Dd7omq5CrFJqjzoVv9QjQAPUIXGbKCKq0ucJHjfqR1eSkeeQr+wW6UO/pf2R9Uer
kZ9M/s3HOew7aM0XO6I3b9YFBh5KZvpO3KKCWApDxa4XzOaow28yncleg6ZH1QaL
/Jb6Iqc2TWoaaKxNcay9jm+S7EWYA9K6/MZgsUGGm0mh+oSS44OsE2CH21D/FVwy
y/qQEjtQ9BnFKRhC8AVp0oFlkvfcbAAzo+n5EVlzeQVR0dXz10fhfyFSBW7gcacU
BtnuSM+Gymq8Ye9dftPcUyZ8R4y/wBfEYbPL9TQcau7yexPOowjfuOm5Q1tRNOJx
svVVnhRDc9VoUOXkcHv5iT2qUc+8tZcyqWW6s5oy/sNp72r74g0+8TQBrPZ02hsd
XlWayZNrqij8u8M1RhPUWtl27EvXrnyP0i9QCwWk9VypsnVzsnZVuOJq20yQFtv3
iZjeAqSNJ8BSKLxJ4rA7xhBdMweAasXTXEAClLXA5VthQcPmNzbWFQdqt0sC5nYn
Q5wykhe54WvGT1SfcyrMiz2aaEfy9PlWh/kIBma4PlvgYoV5lrR4KBBS0ztaPOyP
MZSw03xahAqlLCYxO1AheJIU7Cu/maxnIau9YfbqfMRmr5050kRIZuse7h+AC8hU
IW2osbRIVhlRO8p5UXMKOfWgBFVl86/PrInhvfv2j5+essC/g7sgPg23AURo4Or1
V9iqU+263qOZT4aKb3TBdaJgMgUFRRIzqfdYyUn4bkUuJG5knH9OogHahGhSK6KZ
gy0d1C3EM8C0LwPNrWxDu0o9rTThHP8u3eaz97WwJtO4Y/bE4Ni4ftwrIUb9tqEI
otDRqNiOnOSkxBy7BktTS/84UOI2nq5lXqmU241jJb4Zpc9wJMV8dKEXlA8LcMi9
x3tKYYfFx1UoZcQ5XcqLAkkw7rkMA/hmKSlV+kVI6unx9N4jkt+Kt/8kxmq2wXIs
KXkVxjx/TAwGVwCuG21RH38CK5znLU6KZqN8AEbxn2yW9hAWx299WlqGuvIxKjzQ
duvRD1bDOdP/H3bDchfbxV+HV01zSJbOIf2jVTsa8BlUtFU08EFxIvNIhH1egJxy
NFb/GDfjS+yU6XZu/r8fGKAXjkDtoxf1nFDUPjZAcaYPKFw6aLzOiof5eRMDkAtE
qCnsWOlFX1tPCz/bwdiC/g2EIYrzS6vrxC7acs8NAA4Xnt7Ujma30dIrpqGXhkHI
vabHV6i60p4fT0bLx3dOQt6TOsvbI+lu/MZRlxhg4Smk7UFWb+j/ZYkaWC8Vzkf6
mlx85sjOORyhJS6ncOlMQa7VyCDv5C4yLlHsUH9lcoUDJdQ/rwPx0G/1e8XCDoy8
hfCND7nfKnD/eBpNyVD/3Q1dp/mzeP7zAmzDMWbahpo9gmzC5DLL74klRXByoY9q
O6f3jmg2ptc+XPttaUQBEJPJB4B2E6SL2pW7Sghf87qsy/c09fJ6P/B6HirHeg7O
9OqrR3ha+a+hGnS+ZJLxCJSsxfmPRgfurWXnIRSJBH8onaAPShGzNj7+FxXomoF0
BDFVTFM7/azVYb8JgaennnlnKQ055H6XkEJkrHK47FZgGv5AOXta3QAHRI9EyVf8
ngyy94LsGNpcfedhNC+S8aIkg8mNailA3NdE2yuY36Ukfhmw/l2gGHMHQG6D6xvx
AWJZNqehgzEJ9Qk+HIY1R2sf4EBs/cux0qBZhZinzYHHs81UdfjxkPT59cIlbhG3
Tqc0OskFXKi6yTIgkGEluUvEF7489PNW8jLz3ReQb6MZ/TRAgSPCMMw6fOH3OnaM
WFkujrJvIXWqDl13HJ+LWLnrh3cYDYR1RKs2BZJNhvHi2pcuiJYmqSzYhUGegneM
w2sLJQ29ISFnxnouNV1MhtL4J1jtP4D1HKbk9gEx9T5K8YKP1aPll0iF/+QYD6PF
41cpZEJ+onNaGeAm9PR2s11YprsNchQVh7izRt6LqpV9pcGrmWYnvKxyQ3eURWqI
QJd1O35bAwMs/Rx2P3CXtyITRJ5o9lJnuss7LZEgNZnw0g0oqRqLCXJe4kgWVP9R
JSzNdZf+ClwkT/lxNkoWjIMSHp+gr+EaaioOPhOdEI8pbzH0U+cqMBGrt/7hA3zu
tl2axNZ0fWWvE9RiXkCK0EZFv03DvIrrWMCWxkvkKADHViHiomMtV520XswxAcz2
Ah3xbcqYehfK0KBch1IVfu+CBmJVcCC8ZdAsS+CU/lrjNsDZyNEi67nnFZQQ4Vwd
XBS+xaXnClNGCBQ9qVX3UM2HNBIIb13tjd07Ph+2cw0I/rdGBiYazYl/+C84GPcP
Posjfale0f/hkMNUNTinmY+JU5lTU+gZPGbKs0mnvk+AN/a6RM0NGMQ+9n3d9/1C
PLqkrVoM3limHNKNZ9I+0SNcf3WfNJ9bAawNibCPAZEDOMSUzKW8C9V2opYjWJAU
eQOAPeYecp/1KEY8WJvGVv8e2KOBoATLsSQ7iyMvmrdoVoqOOdL4zzHWaPYbULty
xqKiOZBfWRZSJq77jsKFOnXYcnxy4nnUgGYd6JeQmFkT4ZBFVbkbbysBu2MyIlzs
u/wScuBuQNj5N2pxg39UymGdLXpjBYRlB57TkMDvzzusXp05XrKru896rj17egiV
18g7N45IWdDvsyvm8Ra8UsSyJVkwsa1M5y4HQYPpfoLJVnrp+KOQeIwwkYlePmXO
zFYosVYr0aH1gzBff9KZjtiByJc3kSeySlXfWvStlONAKvn56bgvxD40QkV3c7K7
FEyqtXQwP9Y3Jo/Vd6UXZCQh8iL63fUtN3yqy6IddZ6L3dbMFQHLs90vHW5xO3Ze
9o+ZKEBxiYF5a60Fxxojc+zbvvJlsvgI2uhiQ/ikDDmDqrEkGW1yQuCy/dkZpO0n
5qtEXy7o8XBbJiDEK8njyLyHcOdFB4cbqugA45YwW10Cqo7RYJJRDFY3z4Vo0AoC
mrPmDKRGEzGdsqdJSvY85jnbpv2Skz9k7T34g6TKJC2+AlnKd/g6bT5zL4xRLQNO
oNSSpXswMcasvQDFCLjRhhOLdBiIYobjAPKTAAjMjn75GJZYV50lJM5+Mv4zp1Zj
jRpG4VjUpd6/zXqlU4+vydjbusDzJ8tir37EpjRpSGY6D8DhDvexk3Gr97Ws3Og2
Vt+op5D0YhLVGyUeJQ8QVsQlq0pT8E2jFVoGaqQIaMuqznPwV6Q7K506wciNrdR+
6ppGjE5/ytO4pcQpxz8yR+sHPhaKX08dDIUJhiAS1jH8Ank3YfcoRasvIIipP3gM
WnS+6VFv2OydOFkzkvtGuduIENJUenutMHWxv54G5iZeLf+4OFAv2YXwPQGeovew
raZD+sAeiEvtghffyH+BYxWsy0lgmshr5JQre2Ykpgm3FmqKzNynIUXu8vBB/pm1
JCbzK3j6c3V4sgOKNoJ8yGfMlv/4k8dZj//cqgFhpik1KsZHScpx9bGGWfIAbMFa
wMa4AhQzAAsjEk8o25mJpW+bhs9pw3WgZG+mx0Fe941Jw/o+iiNFR5nFkfrykC3D
/Q9IlQdZw9wZcAV/W6HXXKOaWog45fPz3GZPTMPT2ytx/466mUgcK/S8WDn0gKKM
1JeNlyQ+SAAMeYHaUM/8/2pQ/OLo83sfrEbFjqyBMt0DjRUuUPLKVNnZxtk+ul8+
kbRlrYjs//yQae1Y3ZPskgUPOe2IEhQNP9Wffh3z7eUkeDg9w8rASYQ18pV0gsnz
JK3XBtj6FC8i9Ju12v3hj7EZpuIwkZfG0pvc2ekn/vRDQI5cvj45b38APDbv8npp
g45YLyVf9l53ngYFTQQ36d57sLprlQY1UXGQgbIQlvmgOZaPVAcxdrFQmApKwtlG
s7m/cwhnEbdpyMsHyJbxnjWAMxBGfZzlrSCdbghfZ0B9N6Oi7ZdUKYYzA7BkHloy
`protect END_PROTECTED
