`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MDxeCM/i4dPdPy2NKYGSWy2iqAG/P3AINXnd2ahSwhKdefVkwXYdINAQZFYksPFK
gDv/xOuslzGF5S/tXjwvG+CYRmcS8Q2L1pWdk+x2dtnD+aWNw+EPNfvaZJlNa9Lb
k1Z2vtL6DY9buhbAR6yYWyhsnY4UqarKRtdGqMct0SfNEvPF/dSCjiA9iw5gf35n
tsbWZ9A7O8DgrBO8xwlD5IJZg7yyqYBEKpEKY93c5NlndbYufaZjiAI8D7IAMsYh
ePzypqAcKYuagAFJiXr3JvsbFHN+P20dPjaw7WV+pXPnnSrrS+Vczdr/uv0zseLK
Tit+tnx32enBVpmDNLEfG5yIOEs2h1myLzNQc+db/YHejs9xxmCya5fqiw+USRAA
7/2uNXyzsjv54A62KZv3elCU4imwwmbKzWSnLIu05SPX5YqQTbOnUtylerC8mCRa
HWqT3A5pzHoauhb4lvnlf5YnL/tGEdeAFdc1N6Fof3TA7m1bgMx7Wp8CDfnIVXKL
Pf+Uqr6TcI0M33aedC2uwmbuYSLHbv/tMAA4R9RLf9HBnS4CAkEbYN3LKEusqZhH
2rm4K8UoHiMdjKu2sdSf723UL90snLECZtpN8OVqj0jplPR6kOXn6BrB09I1eUIG
VM3AGKU8s8f4xSxHXYM9AT5Vspzwvo3LVA00evRv7gXZzw7YN6gCITGq3fdGSngB
ma11CkNFVO43mJit9Rmr1uaeKNk61FUzhZ5ZbJSPLOvzH0m68x6bSJqlpDm1FiDU
eBVBTmTwKsTw7M3iJGZDIkXfMm0x5asxhZF66GI3w+IsMDF4hgNoqMdLZZlioceE
zJ18FsSuMXWDJHhsWxTU/DtxjRRXEEtbn6TK7+ugYdEJlk8a/WUUV7+4pYKUUoX1
Rh6sTI8iawW36TBxek54+IxpKlOxTnvC3pK80tPr1CBA3PSiXjxa3jaJQYwESbVJ
xuoqzCNiq3yvvGMwiXe0kQvCRjDjB+I0XsAQxgZGrrKQC6nz414U12cu7puxIdW7
ai3SPeApavtkLp/1HRYvuFFxxJuIbSUBXZB08VQNIRw/JtitiPnvuyVy/1hEFcWe
03EcgxrTErC5HEkO03m6f0cm1kO9uwSzG3NlwSKvMkPJCRKOGJLrrwKVlG5NUEju
9Svst1heX3XFr0FEDDR0tBtiGif+482OHMlLezFF0hp/jihhut4l0i65ZZYc4aft
ajxP7mTF4p8HuTOEhyXxQuWh8ibWbJTqKEz2BQklkHMBi43Qqq7xyEV5sawOnq1z
aXoQXkgAFvSsh1Ivkohwdu/lj7DSwRq6TdNr6K8Q8pKJTeLmqbJJODNlbwhu5S4V
FyDI4e2b07vwvY5MtL6NzxkCIIXLzqINn/QYAvZM8vuAS07bqdaTB03UdCKOVRZ7
7KDVagzQVFvx5pSGpTJ2MbNkuWBLGEFUsYWnlha01ZDhcLj2Hp0Q9HWBzdLWNuth
7e2SIMyd0KpglE6NeHoZ9v51OV4bgNsuKpwpaMHE4aDbz+Gp7/3lFwpWJRo8XJU5
4XJw0z3ihAWLvxSB5ObUBhFjeWTUvgSWDl98eb/MLGv2RhY4a6rATG5ZnjzW/5JQ
RUWuoOOQPspvHOm0tkr5XPWZnlzQreUQwJ/NUJ4W0B57+Te42brsY2roF7iG8XS0
DVhvBjHtWhkT2BAjdF7d8Tl2EWfNYq1w8KjIWd0O8QDHbFB2c0PdrE8/55f9n87k
t5pmTC3vtJTAVyhmxjIx6W0fS55wkXbPEj5bS18SwqkSKHxeqd8o/yDVSpQXW7Cm
9GbPs3ndUaVH1GuaCocJcEZtTTHYEVJSeF16oOsHoNPkStv6N+HmrXRzrAcL5Lfp
/2YS/VxEz6kBeJGKZZIRzFn1lxJTvBiykglpq7NZ+ECGTfqH44fpo49mxbKXI+33
DsdD9Cwb3ULfg1FgsgMEMLYy8S06ckhDYdP0sfnv5BytKVi2avhOyxCA6v/9PY5J
B06/xflg6KdIR9p+1168Xuxuj9S8OMUPMfp5fUK0hraSi0mFX4DKfZ5hg9BKjEog
TSVQM4GYLHZzlVYQOe2kzUfZ3saXXUaBUB5Sp0gkfQWr0BFv/EDReyOCwoXa7GLE
yprfb9XZRnmmOPG6UOilcVjMv5VgmYnRBpRawpJKiVdEAF20clFVfYGS9vnmlCM4
ZSGIfCE7px6MFvoL5klDz8plxPjU8X7n7gOMeziE5sMxUgj8cq5V6cNgEjD7PLpI
eEuBangPOi2uXgaRJwV/KNT+OhsC7WEhBLCv2tJwcE26dUR6ojhJc81yIzN+7EKL
PdjrO0IE7GovFlFx7NT6J5hoG/O+5wNLEzCjC1XMbvh5066G5NFTF+aQxMlIA+fa
3j5MPQiZCWut1N3enjrdwCY4tnrmj7uKjD6B0QB3GLLMzaJNeiEJeOkfcGsEbXdU
uYWOrs0o8TsFGDyP4hIEygq1IJlkyWvEOexsZz6LuOnEA82MOE19FxUVw59W2cYY
EV2cHIbOB9XFLEeAKa29atdSQaCLAxdtc+AqRl7ekbSfNwqXWNgmWMgeKNaynNYv
tZ2dd4XFBR9nkMFi+VyUbPzrhT539VxdqoqlcGFV4cxYOW2n9+beNYhZIOnVpdjx
kJN8HKzY/2+QUAR8sDrczZBRxIdGDmRBtMW8+gLovNEvGrvu9s/ety+TCBpqAOkR
XW17Ji2bugtFIolgbgsoi8iR/IXMQQ7MccjGbfAl6YoOJcPfuw1360KT5/yAfe15
pr5uLUOAe+moxDpkwAZ89RUgAFAlWRLIKo5asF4bTCN1FgZxTDY+mH9S0Qb+mnsp
bTLdB26HUviae7vbeWtH3TB5f09j1YMuHBZZPOZoSLl90Ww9Pri+vOu8UIFpl3MJ
fG38XyoyTo5SUIkoIwiXnn+iA2ikxbpl0VIOFBzgx44XxtKH2fta9OcYWIWOhpFr
OGoDwEdjcZs9QeH58lNW2MWisU3kWHlT00wjVHmYAH1U9TqL6M3aGcKT2kE+t+Ch
MgyTQUX/AFERkxsqOtgUaVHRnZkVEk4+qeutm+C/uBWkGQBCw8bzLzWqae043Oxu
KxFsczX8vz11if5q1fjSx0qjDCE6KAs8DT6ROGL2YdoyqtwsHgqri1Mc2gll+LZ7
kTwzTLnWV+I4xYXBAtjPimD6MDewp1pbnxsQg/lVfRHcHL56iaoe3D7WCjaBevgB
s0OcabCwV/mMQNuWt5qXyXbHAy4hKPE66xoBrHUke7FN5jjJqUqzMxPLIUO4IAhZ
UGvQ+Qrs3LlIhSB623S82btLNX3hjDunxpWo1GBiMXZf4qHqf24gjktJGAIaMbDn
vsbVvzMSA7u56sqg4f+8DBvBqban6KagKHUIoz+SF25KcVtK3BrLSxaTSJ6sM3rV
c5YPHEOVANaQPSWKme6vJld9YxIr+lyVZy2xof+lJZI0ACKy6Tqe/6sjxiriAG5Z
pIA0xCUe07+JvxmzkT8iAKtjOwvm8Tgby737Ezg6jTltcmyhgTS1Ja67uKMQXrBg
2rZ8lhwOpZUKgBPGYMAQaZI47+HwgQLT0gGkrETa4dR9BNx0F/EuNE4DibzCPHYp
TzUB1KkJ0gD1jq3ZHVIpUCllzd450M93T4WHMJFWmSzKZ1/olt1H/F/olXxnzohR
xMLkr1AJU01f/oRuzGxiZAgi9mp91REqwC7u1cjnkHdRzCJ3OTvXigefhoQulI6k
F3HoM9rYRMEZ+v+Nj7jJ2CLhW8y0VlUgnwOBCG/ZMqM=
`protect END_PROTECTED
