`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ICcS8cppjbI+tP6ZwXcx8qKjHTBuu6jczxo9FV2rmNJzZ2Ln9teMNIYM7reOqIA+
EfUu7JDwf8b0oEiRIbDSDtNVZXcy/qurJyj/oXBY8ERfFehJkEdjZjL/blYHYqzp
fy+Juj/zo6dAK2Jw5lZ/TXIvoxs1HlWeNDTz6DoATXSELpje/Ni4ylcfeFDZuLuV
vh0cRmJND0iw+ZhxuyqwU04PDZmBQra6Zjalwo/42RfbDqU8zfo14/z3WRQL3y6+
M9CqGY+sejUv5tPRzQtkSQvf3DB6tQVPPEkJIlJMLBv/rISzm06mQa/cNnmoaS/p
cbl73+VRZ5czmjt+OlFyeWhjWT2ZAI+Nnm8J9KIWct5eT7Xy00seuzzb9pcV+DFz
cMG5ONLZkJ1nLXa7ZrSPMtm3cjcW/jtLBvPu7hszUA7G90mYFJ99nUk6vb37Pvi5
aOP47NEG4HOVNTY2gfhuJCuvaDJKx5nifxxJ/Ni2paJPm4CwpY9lIG6ONjwAwAJg
25Ey+yYKPt+iiA0uJgwLqoxGX4hWKc77T2Zsvs/V54WxlhzZ7IzXFS8YB936jSTg
xhQaedLGH27cPyV4hao+O5B5hM0Wg3qxKAyylid2cPBQRYa6Ww0SoJStoMGOhw+d
lKasy90CVyHeSnJZq83pU6ajtUn5dzCVRJBKDG9MjJfY/0YAdeCPSkC8X/ZKxHGQ
cge0Urg/Ps83Cjy4/yS5US+X7eP1PPIAB02qx70sfLzAsqIq/YKR22qKFiLhcsvj
Yn8rzz+sjiY83sq5te9sCd2F+0cJK/15QySVDHv8WBpiOIf87LOHPD1bwDghzGp1
nJeE6CTBMM9zMEKBOD0fmCxwI9va4T6mii93zuuvuP16K9EZcoJHqZptNjXtxyIv
UoJWhIrKae4CRh02X/g+A73Y5qfwZhU9LKYBuh4NGHR0P6bmBPkQ3dUHqB5R+R48
aTfSwUAtIhu50SOjeg874B+DLbT+Qz35pCT19Q/cVjlC6aIfe6nMSN4Erqgg2XNS
cxuRfsp6906K/6Dza0lpQEvhpHsaxMNn6LQyWzk99hl1wgdgnb8zT5OCeR6BsIzT
/HhC/HdPADBucqJxs5BoZdnLm0kFjL3+ePWT8YcacKXFoTBMmAHSeEvPNBajiPEM
ypMUOcID7r+w+IszeCxPudjuXFz82qHX+1nYYaAaMCbTeaOstY505FKQZG3AmnKt
YaFyrI/GrHq/xbnQrGokNUMsBl1ISWiB9FMqdNEFEk1QY4hDh4rgnXZg2RAWEoWx
OrDZUUpQISkUFSxShU3cPR0RCDcf4vdVGc6yANZVgUyE9T29lj/O7sgyMu/TziL+
GmnlXxTiwQp95MtxIGlh7LinrC/MvRQuWFMC+TciEY8E3BSUsDDYlChp3k05Lkho
dt+NPTHjR2ejdENt81XGhObMKgguDYYmWP1hwRJ8fhpHclIZJNIJDe34H/y3GlYo
Ojha31vvW35WVc2O06Kta/oEyuzxF+5TBzL6ypgShGn7JXFnkmkL3aspoYiE3ycH
A7syf9I8u0+hskvof86QotNAxbEG/6TovR79svnRvEGaXOS+de2ENJLs0lja37z7
07mUyv/mzJwWJ8/fCC10lkNHkE2CHdk3hLEx9EMF7tnIPzlz+lsJnLVLc/cbSHN/
lp5mYLeTOOh61FJc+4ah1CWk75UtJ5PX7uF6jPYMNoq1vJ4ZSz/qRDwg59b/D3z6
RSnvYctjmc/jueM8jGsicroQjRQvgvogYCItSDBp8nRpDUSbkxTAqujQ3vncHhBI
JGzu3bwEE/3NkvAkujKY+wFB6wfbucQe1A4vnWghg82IN5XeVBez4PDQ+fLaahNW
a/7b5KY4aZa7APJKYHeKmfnC66hhS0/WbToDFzUEIbqjLyxrSWt1FDrSfiGwPL4T
EOTXoAT3EWQmUIVoI+B3f9iJxVdyXHymCsSdkxL6SZhP9iMWlo3FG/Np3m2kbQhy
orf6Jszf4mOUpu3sv5ja/B5VHsKzTyZITdKNlxU8rQM/zzISYmkrmQ9udIPXZ9gP
Dnagaj8STTpU2vT+q1G29S54S9RAiPlE5vxtFgEXWTKcAEPCxO6dwK0kvm7amxsJ
SuDfNeuateW24vgeBvBSKKryJRdtYIxZJNvZWh04PPlgLW06PlL0gG4IqONlWmWj
DB96WYxpBELkiSRKOLK8tqiC/WtnIHF3ea7N0ScTihKZ9auGXp9Qnkz9CuM1p6tJ
XDGdPwHlW0oFd+Zl6aeLetZuVVRq5TXGIxFKBvq8uP6WnzxO5iiKMkygrlK+XJq0
/SE+ManAijo7kU1a4lqNQ0pD5nK92V7ofmryAYrHfXpKI5e4sJe1JKwiSN/frI0F
vdYcf0BRst+PdyRTePOiZAsHLmYzQI5gqiJPUqvuphQ/nR8u6YcNX7xcbXpdGKjm
ua34w4JuRJsjEXFvqOTCxHE/PlwDBGmdbxT3sz/qHk9QA/7wQgBCp4ggT3LziYGl
JUKt5SMnroV6U3a5Wb5gG7aeZdeesNsmc9VYCZSx/TpWbZeOg8pC5lBTAY+HQGsd
eEze2qEX61Fn+c4SJr7gX0+Pw+9xoyAA4JCJHxLG1ge2NJs93w/tGiutPSR/+Q4v
702eJDVV3WWeXvOjV6N+twWc5YqJY6brwe0d2D1f+L8=
`protect END_PROTECTED
