`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GqHYfHF8fl8bZAd/bn77PJOseUR33lqpK7QILdxa9g+5TO1qOizHlLoL63qdCJ7/
tyZ06ivBGUf6/gOMYVW/ojYARNpfD1GoPQpzlYs9uQPTWAcRnEwdyQTZoQp/XslD
Xrbpa3CqLSlO1vDBMrDa12c31vjiIfo90pyy0ECMa6T22hCc6ILdlax1PPZWAsGp
lWlnzFjTD/EhoGftta7az0N/1DWPTMaXgiOdLbrufNediXC1jYzDwLfFQp2XWv8M
BxKHiaNrW2zX3JfcV+KWm9UgKLRNqOVGVbMymSvLbtUybGbEa5M6PCZHno5CAQOg
9tvQCWgQqtSIgu82cX/LXu9ar+cebz57BFjuiDAN2P4+RjDjYHdnB8bx3pJHER8e
4TSgfKTiktmACb4SuTcskgO7Q3MlI1QVvjZ3wILlUnwI2W3oTCqKJzXptLlR4aeo
LqR+e0x1pyIlSsAXph+Fj4tHJOKp115M12C5Of8/c8Y8EUvp/rwRboWybzoLcUkt
4FQ7VdCCL7QFMjBUEf7r4L7BA54BTKjrBdH00Bo5vTkYYD6+ZWXBWd5ADa7g2wdh
1nN+v6sDYoTyao9+xOYNJPEb8ptjYOvz4DnxXqgRHs4q2OvrkcL7Z2vlwQpnhcf4
qQG/yVP3H7VkJRyjahmpWmpHkjlGGTQ5/7QUrpjvlPn1Bcwsp0lHhm0BLRC4TmxL
h5ZMo4ehc0uSNnjGE16tyNTFWHNcXM5z8tY40aKR+pVHZZhooY89lF43xHKyMwR/
SfPsPfzsk7Atw2ZCbUcKIz7qfTDGORhSxn7IEvMzs92A9fs1Aa0dIrgfIYSArD+R
SxySQH7h8pf9ft2pyydPV1XMJ61wV2h3OrNO8YcuB2MOH75gOFuxd5mWNQrndpdK
hhbV2wVWAYWndfYVncRTdalYxeWdpWCPM5IQLBluuNN61gPixaZqa79qFZntr+7B
kKanc/Rjx4wu0kZd75WnzAmr5hop5GAZdTH5J4J/o3zdYvMZtRzkMSC0+ZhTaz6L
2RZXn3D3pIiwR1a9+2PZZ++Pem7WqijYGnqWUy0Mh/lqxEk/pLc8RofhU394AZYI
OQgJizZac5Imgm6zPmUxMEGMN7TkqHLqECQAbRxhlEnL3KUaheI1nyqhSDvFITop
g94ndu6AwRzv4hwM+KUQRFS4EcE6oxLwdA54CtE5M72FSaJpaYs+qtI88pE+DW4U
D26nkOXImBItcVrzjSs197ukGYfuoiXHDRitwLUS7MUlKBYqkWkZWARj9BmKSLgO
8JUVNuzq75qGvYOArhGrdzi37oBcUIL4+G1dtjw0xYeafPU/oWMdi6mCHGefYQo5
CsqdM4OqJb5BxplqKgEzVfa9+nkofNQy4P2LlqchIScKglBOLqR9KIYtQtc1nIUL
3AV+lDZFgRhO1HBqFyGIuyhzDDutHXwq3hrIqw2ov9rqw+AyX+v0h2ygaXvFdKmp
JQaHLF0SR65Kmd5pEg1n5zHDSBUCZSbnMnf+dMbVaL8g31PP7y5+hVh+q25WgKRX
5xJtPEz9qH1N2wcFVyh3vM2sKkfZL4GV+KQAkWFClqAXnSulEVI4z3IhqEV6s4wb
cSNTQfXNHhGCyAf9214h9CMnUpoXm43AkAzF6GPUdOb9Z7lNLB22ttR/aPx/nO/E
KPRwN071J2QlPOC55ZxhmqMczIB5+qfrbQznjOx4ODkYESoP76vrUWFHQe9tMixa
jJCRX8NhPmFqKynIOntbOkiCrFbJk0V/DhE6WSE5W6fYCmQwXHom3SM0qem7fzcf
Oz3dZdNvHJ0aSBk6cOnGFGQ3scAIrl6wcbBHCAi98fWNANinanpY0+A04+DHczBD
PMUMdyYOW4VcyXNh1Vo41mfE1qTRkSE2HIxSbSrKa2HpbBdCnbfgTrKDotO2YZDX
VEC3Xzb2Rh9lJyAbFaAeXXrBb6gqEAZsQO+VBKyZLXwjNhvmN2m1RwNaf10SJdVZ
h6ybGUBUSgDTAWZsbGmB5ublZY5ctxlPD0KhbnGPuD6B68RigLr1VInMfcSB0Kzi
ye3t6HiyC88hObv9LnRqLp+JLizwjZce43FiFvJiZwRxWrCUAHcqLS7Wt+Ldt3J7
mX5zfbFrshl9k6F7jIrQaKyigkHEErUQxUrnm0FFMs4PSvopMqHI+RoMqOHMYHuV
2OdXmR/KLaXqOq+3QnLjjg==
`protect END_PROTECTED
