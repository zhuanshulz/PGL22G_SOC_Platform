`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nqGHm0If1Nx8dv5Qu7lq88YKyio48/tMHs4fHcdaGNznQWZgTJugalQKr+Bqvvgw
Y1zKQl+1vQHcNMAfdLT2xjOoMOGZFkfIPhpa8TDbbtmfQpMrV3OSoAcZusv3xwaw
xGt767trrWEr6BOAd1WZJliqGklYMsaz/a4Tju29o9ZxooQEA/q9sjm49FkA+Ymn
EwqUQSCMYLbKKkDVB6yjRIVg2G0RAggp8TYBdFqmjW2gBxvcny1OR6ZmREEpHrgk
++26xWf44u2OKQkvQ6t4F+CFI1rntXEsJpY9/2Tyyl9YAic0PnMEbexatKxPSgmM
SxJ+97myYd9aUEUuHB3FkXTrqqjGb0wKsjSIxnAXJDsVpP7ye1WVianMbgx1qaXO
3Efex9Nt32Fu4lg5np9JxgQvh9FMVYcsWszUxbaFOhfwtEFiKcQRkD7xKw4NF6l/
Jlqc849tA4K2b/gw4Bg6Y0Ygi1yI0/bDa5ADMcwj/lhXyHbJktk+KEzamqpYD2um
v6KZUjXMdANYq1VH6Aa/hFm6AuIrh+nhGzVBI9A0TLtG8VsParZA4+JUeRGeyMyc
2JFNdsjgsmP6jygCiG9w+aU+DDgP4a0J2n/WwzcCUVaWOzVjHcetYQ4YVnL9sinG
T8CQIxnIp7kVCxUlp2nxw9beKxwnqG4Hl8uMvndheh2pt6IUSwAtQSGyH7ZuSdUQ
/xJ2rBLNV5wgiU6CMog4/nJj8FoRNCM9pwDfB5f5OEYif6ajl+wqZZIT/n3L0IcC
cMz75DbACmoKaM5Wlv1rhgHvYzTTdTiA/i5FeqAi52pTet54ZUTSTankUF4MvhOn
GULVj2nMZEAeV7jlfbb6LmEWMHo4S6ZaqFoNPccl4T0C76HwNSgaZRRMV5Bk+HFt
3Mzbr31SBhMFRq1lLz0t7X9EaQsg0jS+hwNR9h82HEczfDEKKmDeNBA1DH49bz3o
ObDMa6NkHrab0mPCb40RSk0YKyNc87UHBmQtMO78lQTf8vkf3St+LxyVTsJKEd5k
cLWNFZordTCePH5I6GMNGIEqd1QC5TJiqBJLs8SUEpaeaOwEq5iQmGf7G7tUuN0u
lsf+fTDtshM3SUf9QmP+a8lcB+b0HJE5nBWmRx1r474u7b6HQbqWCfscgEEQpUGd
pH6GbrGgYPkiH2KDA+bU4fB2Fcnx/OiZ7GQTWpAehVzQkOjrQat46LIG5LFOYGgp
Z3LfwD8+RxT1qXvZA5/70mZYrjNtA6z9kbSnoKXUKaCdocC0yZFPbj7+EZpRhQHU
e05s8dkYpP46n6QUEN//WMnUezewY9YlDgkIRAjUe0lG7ytA5nY2Igrq4gUYZdB3
8ylRjxPA8B6B2jkkYhj89dyZObtenKSJ06d1Td3SSrallPVg00l1bn461nXLm+ZJ
44OhSNLpL5TDuMau6jvZ0bZXISsJ9uQTYCGw7mTjY0BUb3LSE5FbBQDmRt3nD5xs
c+KSxnHBN+YIc3ab+CIDx5qOSvpL14DWWVc5bKnvuEB4Ih+/mEJ608wNTVgxghAT
jyj4fwUdpTGvLM8pWp2WWn+y2Av1VsnOKsN0+WlxAKQYpeFInkQYpFMscMbcralD
DAa6SXPi+H/JH+GVjBWDfqC1KvQFW05JRmUIpiWINgKQcmU/SlA4l7LSK/HopHMh
kWNqkDtBthyDKwi4q0lgiEvxaRE8O6jz3IES1mJY2uJNj1IXEEzKyAsTgqTzGBm9
x2jl894l9hCRIzxeMChd1V6KvS1Ca76JvrpbeU/CXgRmMgnEDDXVdDkeTPTJmodK
RJx6FwXlY7C8qICnRR2+fgS2JgdMZqfBBYnFTeOc/b/fS2rHfVGiyAbpY9vT512K
SkoJjJOGZCESSmvRugYb/+6j7YlUCCYll4PrGfX0deelzJtHalcevZNDQzo1LgJS
CQOA5bNEsHI/q/HzxaG7Szc8CdeKPGLZnyZavrjft9cfQy6pFyboA2wKrJpQ1yd0
DxcEBY9ezUklFfIUjHD+/bsQY2RWqA0NF9DHtOLB9jhHBbqkqkCIW2T59AsdCSdU
/WODv4MZd1J03qll2c0exf7tWMzcugOeBDBzbmZHEFEZ9NufNHKp6LmsCjij6rCl
K1iKsoKXfvPVfw9rBYn1BAkHTYf+yS38iKSI4MNp77SZExC6Bx4+O2vRttD1/S9Q
4NtcjD5o6QGfeyNiAjVdLawFuvecNwEASsnVpWinTF7JXvunHW5D6qDOIIdbzhA7
9Z/wfhaoM4a2y+dg7ui8fh8/dZFZZW+vE4R+ZoVp7ymZ81dWyFXO0A2QNBIUTWn8
Sa/WjjR61dxr22NxV0EUYnyCbBG2wZSR/XTGDqqMZjvgATj3ocDL3M9NZ6lrlJ9T
sg82vFmOobG0EWETSyMd7WJCj1bk0DGR+ArGrX7Mk0KTUJUi3aKUWhCpc/CjkaJM
19I7pe6eSUBa08AoiNlWmZbQQvU68UyJqg37Ker/wfntT4Y69amyq/dkYOiy8Rla
x0tUmRjyLLgUtuAXIVFgaAMAAOjEZB9neiy0E+UbRdjGAWclu67SLzEaiPUmw8d3
AbSWblGoOknFLYkrFmE9P2DNNdYx5Qj4ZAULKHXw+kLydMQetDC1dQlUm1ssSCKe
A61VyEAU21bmm1o4E49rsuHGfqYLo0qEIXyuNtw0agVBtio/KNYGlRAVXB6Q1PxA
Ns4UIE7L2Eryre36f1gDAIizapmAfPaQM06qgjIG5bYCoe+rkSqbRqQWGPvAVCV8
GG2ZlpAXLevZnNBoOIUM2GD07rByh5R466ydu1cEwWXmyyDb/bnrRwLpf+Ay6Rt8
FES87UTshs9OdtPt+7RTvPXfjuP5mQDmGl+bmGqRCMVASMYZNumoxtxfb2pvDbxL
IshQu34m9D10C5c5+AHSkdPsZwKDeNUTYb8rLn+s+gg/0/GfEsEIUGOkNtl5EaYE
Vb1yxLTU0cbbQ3Uv6hCQ1qZcVbaWl/e2EVv6dOe9rYTMVeJ+GPuXU8cU2MA2Y/hr
hT1XQTNJ8TRvKh/Y8Bbt+XLbhWTkpDVvDCLitbr0mqmeL3ouTl/bJq9WC9bAb9Xy
B3/cWAEYr7ZhSTaMV8F7i9+VWjKVk2p+DKIci4adAgB7vqYUNcuKWXtb4IHJHlfS
EpkbAYiRwWVZaea5CJ5MATBCLJMwsrzgniJVjSL3EgCOo+S7NMgo4xzxdPMzu1a7
hILWUjsblgUjVG8Or8umEJhdHeHFXqRkxFcHtNM56v1O14VyVQMVURoWLTmqNQw6
LGa8WP0aH8KYi9S1uKwpV83r5nI5Ow/sxobGDkd2xHtxamP+UwAsetjRC8GuzExn
m88Lyv7PM+32Y80EVYUIRt//PKB2D6z3lBHZFLelkiWr5PWMdYCWuwLAkSl+yBfj
ALn8cJLnWyr1KAY9ZOlcVjwhBuM9uQYMr9AAe6mrYnbfr57wnCO9oBGHwcpiG5Ya
Dg/hZWXrWMWWVB5bDDuHy6kl3WDZ5tdzahBFN6/2eIPOpuVLmbkWs+YP8lSwJSYW
/rPdeJnIL2j/IKYC45jRWL2iZFb5qurrqC3LosNsWAngS4IADt+1xxnRQLDvyidP
zH9UsZvjzJcm1tbih0C/OYXyjZWg7WY13vY1t7BFseHh75CPueiH+VQSniaC2hkV
Ce605K5N/qaYyNjCNxrG6bKR7+KSiqQjq7/XO7OApLTRYVEeSUon0sa6xz7oARg0
V5YzyM8XGkWDzt4xawGN4GHfAGMJkDDyhfue7W0NBYEqDcWJvFaQHCjkOmq/CmyU
9tg0FuudeprkZCngXAZfA6xZDr8VWbkPIrQEfjH1GMt3ur5gdm0Wr9iaRPmI9d8E
Ba1bQS72M1ME0XRuCUppVuF/VC6rQEV7UqnabSw0Al4tr9iNp9GR6NKbvL4oMz+O
3pFx+vQn6acMcHrtb6m8lFM1BBR0l5R2KJAHP2nrtxmXQQF25LHrFf1Ueelp+9uR
R2rSNwqAAUAPR4SzGn2cOgFAIDs6XbiC5c9rBsXDIH5JUMAe5VaGTenSdamybvMP
ZjVAMcIz/3lH0nqzF+bEq36jjlAWxW5h4VLw9zqPvbmuWhLrcojqLIJ7m89O/VKt
2wJGqWp8RtGVY1ZygCaHTPWFtZb7fqnCJwiadc+t5we23idc3IC3kRAvLnlYJTrq
2hq6Ykf+SR4q4RxxLbwMARySqtLytTi/dsAekRn7r5WWrj/Cl6XqCV3vcVnwJ0CP
ndWUvVjo8tc4NPnoEU53zAe2UNNwPxJtOGflTF1Q0K5GH8pvPBAe/gr7rQL7K5fj
yWLLDDyRRLjwmCZsvdku/6vGXIh7Una7KgK7pz8OncrYiW1rw/LqNaAMEOwpJosD
ERTbrDahCb7I91JB1QzJax1zGt38fP9WbARopG6Q6lBYu1JjJtMEbv73vSfxvmKG
6Qym+U6kd79Ipf7O/Q66ZN4I9LQU9JTDC+6wXs9z8YxGP1sZQwDX4V25NJyYWavD
yr5p1iiA49UyjxHM9Tgwg2ZrigWfoiUWqM9OV9QFkf9F+Wu3mIiSE9tSftMmslsr
klvHBnRQLvMs97CK0Q6E5v3GgRS+C7F9WJI2mk6coPEIVP9sQZcrhBqXso2t2SV0
cLew3vmjfBu0QoFTP1UHVdJclrmXCdxMhrPZTCet8WvM3y9A77I2/pwvHfKfTun5
hFJd+Fqd+A9UpfEWeh6+liM3PdWOGCcpJUSCH/ssPXRP+bEzpsB7jvcPdsAjrxWu
omzXdUfkbloISCaZbcjDQOzmCccWQVa8wAP1DKuFy79unHr+0WT9L0ynYcMlHd4B
cKndPV2sbou1XfLzCFAH+CQw0eF8ycXvuP4y/BOtpFfFqtPY+ReFszYIAyVvD6eg
V0a9S7dJmzhVlyvRM2QWk68acs7O2Lp9nwBxHDTFGhwvk4X3CEGB3lpbgduUIy7D
stfeO79faWIlpUGRlMSVmm5oxUG/NgQFXxdagpyJQ1KduU8T2AnB1vsuzJZL6sxk
CMVCB3Dk5kxDf3bSBg0ClaxDehP/zhEGub3GyLYgwkXzVTBiVJxnUGl8LHPenRzG
xLARzrf8YMPPlpTGg4cTi+0CJGSMqfO102IQc9ntO0uuruX33Mbxs46391fA3reN
rbgtDJFwbTdKro8BknpMcOnE3rHKQaP3AVjw+K05pqW1kS7zVy47kGN9AhrZf0iT
68jFBYmq7vTPRaJ7/u912mxG/QzvOehFazXHNkDoh7M5NDsExXyzDFAht7myNM2w
g+f9boulb6ARXrshdhS/K0UcAMFMjm85hi5zoRZN7BoyTEIrXpP2yEwFlfUVvGph
VAszxuA8tEeXnzU6NGbXS98krupA3Ms8w2mQKO/oGegz/FUnLAPVdqlHB7lY0BGC
6lZDmfSVi0tgrf9MEZbgjRHn9aJbuAIKnwNboUFmXQYNBUzuXsJndInhBj1CO2hD
LoY4W7JvAg71TZ0vJyS0tCOVwJ7CV7JuKy0hSSbng5X/zwfclWB7RNF+rWtrhgnj
7yzL/rSjXQI9xeh0BP8UR4qBdqqZ70oZVSOycBr1/YC3hOMS/P56RC7szOCPtYb7
g9AdrCLuH7TZCs/nM/nzaRvl6g8g2UWwBXSaWAC+84ZNRbQXt+89fWlkBRiDlKlc
Swno9qQmhsqOs81OUaWzyX19IoZs+xWURFsMHyrPTtcxvVgSJjZye7SvJ3kyQydq
VaK2UavfXXwFiWg+dm4fIG+CvMfK5Ua5Q8bl9DgkQ0rQJblNxi18T1doxd7YId/E
DXrGX2M3WK/LyDVKryZQS3o2LHFxiLnqvBxl+WKQEJS2CwYD7Ib4pI42NMXNWwRM
gLveAD/B5kJzOBY8zStN+LQVkRX/UsF19FfINNrmgUWdbDeG2A/BMTEPZ+/uiS0P
spIMydXw8F4BcVqa3gNtiweA5B9cBxa8GyvnuHUiu6OybuUjRj+pzYkcjjvLb0hX
Jcgg4D3p+UiSLWNVXYZZCxWN2Amc67+ssuJRj/+lRX2LTCmicgNsxsXPOdW21d0Y
TG9sy5z6+FfUQCgAMNPoooNz5miLOGdMXkIRohT6RBUISQYIhJJKJPcdFN5pSgAY
N8TOLKY7ZOJ+qDblzSNzhq6wR7a70ukVkJJbfQcGwsaCpioWh1rizoAx98FYOF/7
8z5XI02rh7iTOkU/YMc57M1MSK/4d1TmFa4z/rSt35vkDi4X5v9j6FacMXVmZzty
kTi70mNEXSxCzdQRw0tyERU+1FILf6/O6xXPpPDPgXEUZQOlFNKRcUv5wvv/iKqT
ZOpWd1RJc4fuUWYapL9WzD7w0laONQV3rwfpO/strQHGR2hOIaTfAzpE4bjQuJLB
5syOs6MEwya86hPeR5W07XbFp4jAR1my8WNe9dJxFrC5xdA73k4Yu6gqcC/j715a
JLn2p5d7MWT2VdWe5lCBwc2DJfjheDvMAyB/aNqmFnZkm4gsb9owuPTfQu3o+Aep
5uqawvR/Seri5ABDORNtVdNrTZ/21c01VGxSztNnNVDNWhcdjgEG1y7qJcp1QBkV
x4DWcAZWFRuKxk0+cfPDZPtrY3A5GNVUp4pplAgYU9T3Ba+27/Wx7DauwsKqPu03
kZeLroU87BntMr/FkOz2qZdK1aE1GQZ+lgRGON0mLkwwKmvasBST3BQskDpRNSFf
6Hl0DPkIDC0+TgTEr5SKpwS8zZyCXTM+89BiiZ1eqGJ7neyYoDt5s7x4LxMR8/qR
TurxTJBTECmrnZ+VDWqS10Y5sJxVb1voum8ssuqd5tnZgn9EvcSmY3Hs2eEQdrGp
1DCkKZE/lg0FCLCms/7ti5y/gYpWEeBdWPf+ZwYjaRuHw3gJdYeLHWhusAClpGVl
DMYumKM//RhduiyFbrETMqyXlhkd3v+U9/jkyMO7E4UMYTJO2LLbUiSu7A9oxHGy
kAaYUA0tFcSgV2PLA4a3u+S2Xd3UuSlR1rV9aiG8jr68GtV6SoG2NfisR51FR8J9
tGwQ8uSL3GRM8RXThn/rI3nsvOO/7SLggCfX2uycdCI=
`protect END_PROTECTED
