library verilog;
use verilog.vl_types.all;
entity ipsl_hmic_h_phy_io_v1_1 is
    generic(
        DQS_GATE_LOOP   : string  := "TRUE";
        R_EXTEND        : string  := "FALSE";
        CORE_CLK_SEL    : vl_logic := Hi0;
        TEST_PATTERN2   : vl_logic_vector(31 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        TEST_PATTERN3   : vl_logic_vector(31 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        T200US          : integer := 54000;
        MR0_DDR3        : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0);
        MR1_DDR3        : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        MR2_DDR3        : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        MR3_DDR3        : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        MR_DDR2         : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        EMR1_DDR2       : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        EMR2_DDR2       : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        EMR3_DDR2       : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        MR_LPDDR        : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1);
        EMR_LPDDR       : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        TMRD            : integer := 0;
        TMOD            : integer := 0;
        TZQINIT         : integer := 0;
        TXPR            : integer := 0;
        TRP             : integer := 0;
        TRFC            : integer := 0;
        WL_EN           : string  := "FALSE";
        DDR_TYPE        : string  := "DDR3";
        DATA_WIDTH      : string  := "16BIT";
        DQS_GATE_MODE   : vl_logic_vector(1 downto 0) := (Hi0, Hi0);
        WRDATA_PATH_ADJ : string  := "FALSE";
        CTRL_PATH_ADJ   : string  := "FALSE";
        WL_MAX_STEP     : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        WL_MAX_CHECK    : vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        MAN_WRLVL_DQS_L : string  := "FALSE";
        MAN_WRLVL_DQS_H : string  := "FALSE";
        WL_CTRL_L       : vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        WL_CTRL_H       : vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        INIT_READ_CLK_CTRL: vl_logic_vector(1 downto 0) := (Hi0, Hi0);
        INIT_READ_CLK_CTRL_H: vl_logic_vector(1 downto 0) := (Hi0, Hi0);
        INIT_SLIP_STEP  : vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi0);
        INIT_SLIP_STEP_H: vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi0);
        FORCE_READ_CLK_CTRL_L: string  := "FALSE";
        FORCE_READ_CLK_CTRL_H: string  := "FALSE";
        STOP_WITH_ERROR : string  := "TRUE";
        DQGT_DEBUG      : vl_logic := Hi0;
        WRITE_DEBUG     : vl_logic := Hi0;
        RDEL_ADJ_MAX_RANG: vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        MIN_DQSI_WIN    : vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi0);
        INIT_SAMP_POSITION: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        INIT_SAMP_POSITION_H: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        FORCE_SAMP_POSITION_L: string  := "FALSE";
        FORCE_SAMP_POSITION_H: string  := "FALSE";
        RDEL_RD_CNT     : vl_logic_vector(18 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        T400NS          : integer := 0;
        T_LPDDR         : vl_logic_vector(8 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        REF_CNT         : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        APB_VLD         : string  := "FALSE";
        TEST_PATTERN1   : vl_logic_vector(127 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        TRAIN_RST_TYPE  : string  := "FALSE";
        TXS             : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        WL_SETTING      : vl_logic := Hi1;
        WCLK_DEL_SEL    : vl_logic := Hi0;
        INIT_WRLVL_STEP_L: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        INIT_WRLVL_STEP_H: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0)
    );
    port(
        srb_core_clk    : in     vl_logic;
        pll_clk         : in     vl_logic;
        ioclk_div       : out    vl_logic;
        pclk            : in     vl_logic;
        preset          : in     vl_logic;
        paddr           : in     vl_logic_vector(11 downto 0);
        pwdata          : in     vl_logic_vector(31 downto 0);
        pwrite          : in     vl_logic;
        penable         : in     vl_logic;
        psel            : in     vl_logic;
        pready          : out    vl_logic;
        prdata          : out    vl_logic_vector(31 downto 0);
        srb_dqs_rst     : in     vl_logic;
        ddrphy_update_type: in     vl_logic_vector(1 downto 0);
        ddrphy_update_comp_val_l: in     vl_logic_vector(1 downto 0);
        ddrphy_update_comp_dir_l: in     vl_logic;
        ddrphy_update_comp_val_h: in     vl_logic_vector(1 downto 0);
        ddrphy_update_comp_dir_h: in     vl_logic;
        ddrphy_rst      : in     vl_logic;
        ddrphy_rst_req  : out    vl_logic;
        ddrphy_rst_ack  : in     vl_logic;
        ddrphy_update   : in     vl_logic;
        ddrphy_update_done: out    vl_logic;
        dll_update_ack  : in     vl_logic;
        srb_rst_dll     : in     vl_logic;
        dll_update_n    : in     vl_logic;
        dll_step_copy   : out    vl_logic_vector(7 downto 0);
        srb_dll_freeze  : in     vl_logic;
        srb_iol_rst     : in     vl_logic;
        srb_dqs_rst_training: in     vl_logic;
        dll_update_req  : out    vl_logic;
        dfi_error       : out    vl_logic;
        dfi_error_info  : out    vl_logic_vector(2 downto 0);
        dfi_rddata      : out    vl_logic_vector(63 downto 0);
        dfi_rddata_valid: out    vl_logic_vector(3 downto 0);
        dfi_ctrlupd_ack : out    vl_logic;
        dfi_init_complete: out    vl_logic;
        dfi_phyupd_req  : out    vl_logic;
        dfi_phyupd_type : out    vl_logic_vector(1 downto 0);
        dfi_lp_ack      : out    vl_logic;
        dfi_address     : in     vl_logic_vector(31 downto 0);
        dfi_bank        : in     vl_logic_vector(5 downto 0);
        dfi_cas_n       : in     vl_logic_vector(1 downto 0);
        dfi_ras_n       : in     vl_logic_vector(1 downto 0);
        dfi_we_n        : in     vl_logic_vector(1 downto 0);
        dfi_cke         : in     vl_logic_vector(1 downto 0);
        dfi_cs          : in     vl_logic_vector(1 downto 0);
        dfi_odt         : in     vl_logic_vector(1 downto 0);
        dfi_reset_n     : in     vl_logic_vector(1 downto 0);
        dfi_wrdata      : in     vl_logic_vector(63 downto 0);
        dfi_wrdata_mask : in     vl_logic_vector(7 downto 0);
        dfi_wrdata_en   : in     vl_logic_vector(3 downto 0);
        dfi_rddata_en   : in     vl_logic_vector(3 downto 0);
        dfi_ctrlupd_req : in     vl_logic;
        dfi_dram_clk_disable: in     vl_logic;
        dfi_init_start  : in     vl_logic;
        dfi_frequency   : in     vl_logic_vector(4 downto 0);
        dfi_phyupd_ack  : in     vl_logic;
        dfi_lp_req      : in     vl_logic;
        dfi_lp_wakeup   : in     vl_logic_vector(3 downto 0);
        pad_loop_in     : in     vl_logic;
        pad_loop_in_h   : in     vl_logic;
        pad_rstn_ch0    : out    vl_logic;
        pad_ddr_clk_w   : out    vl_logic;
        pad_ddr_clkn_w  : out    vl_logic;
        pad_csn_ch0     : out    vl_logic;
        pad_addr_ch0    : out    vl_logic_vector(15 downto 0);
        pad_dq_ch0      : inout  vl_logic_vector(15 downto 0);
        pad_dqs_ch0     : inout  vl_logic_vector(1 downto 0);
        pad_dqsn_ch0    : inout  vl_logic_vector(1 downto 0);
        pad_dm_rdqs_ch0 : out    vl_logic_vector(1 downto 0);
        pad_cke_ch0     : out    vl_logic;
        pad_odt_ch0     : out    vl_logic;
        pad_rasn_ch0    : out    vl_logic;
        pad_casn_ch0    : out    vl_logic;
        pad_wen_ch0     : out    vl_logic;
        pad_ba_ch0      : out    vl_logic_vector(2 downto 0);
        pad_loop_out    : out    vl_logic;
        pad_loop_out_h  : out    vl_logic;
        dll_lock        : out    vl_logic;
        srb_ioclkdiv_rstn: in     vl_logic;
        dqs_drift_l     : out    vl_logic_vector(1 downto 0);
        dqs_drift_h     : out    vl_logic_vector(1 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of DQS_GATE_LOOP : constant is 1;
    attribute mti_svvh_generic_type of R_EXTEND : constant is 1;
    attribute mti_svvh_generic_type of CORE_CLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of TEST_PATTERN2 : constant is 2;
    attribute mti_svvh_generic_type of TEST_PATTERN3 : constant is 2;
    attribute mti_svvh_generic_type of T200US : constant is 2;
    attribute mti_svvh_generic_type of MR0_DDR3 : constant is 2;
    attribute mti_svvh_generic_type of MR1_DDR3 : constant is 2;
    attribute mti_svvh_generic_type of MR2_DDR3 : constant is 2;
    attribute mti_svvh_generic_type of MR3_DDR3 : constant is 2;
    attribute mti_svvh_generic_type of MR_DDR2 : constant is 2;
    attribute mti_svvh_generic_type of EMR1_DDR2 : constant is 2;
    attribute mti_svvh_generic_type of EMR2_DDR2 : constant is 2;
    attribute mti_svvh_generic_type of EMR3_DDR2 : constant is 2;
    attribute mti_svvh_generic_type of MR_LPDDR : constant is 2;
    attribute mti_svvh_generic_type of EMR_LPDDR : constant is 2;
    attribute mti_svvh_generic_type of TMRD : constant is 2;
    attribute mti_svvh_generic_type of TMOD : constant is 2;
    attribute mti_svvh_generic_type of TZQINIT : constant is 2;
    attribute mti_svvh_generic_type of TXPR : constant is 2;
    attribute mti_svvh_generic_type of TRP : constant is 2;
    attribute mti_svvh_generic_type of TRFC : constant is 2;
    attribute mti_svvh_generic_type of WL_EN : constant is 1;
    attribute mti_svvh_generic_type of DDR_TYPE : constant is 1;
    attribute mti_svvh_generic_type of DATA_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of DQS_GATE_MODE : constant is 2;
    attribute mti_svvh_generic_type of WRDATA_PATH_ADJ : constant is 1;
    attribute mti_svvh_generic_type of CTRL_PATH_ADJ : constant is 1;
    attribute mti_svvh_generic_type of WL_MAX_STEP : constant is 2;
    attribute mti_svvh_generic_type of WL_MAX_CHECK : constant is 2;
    attribute mti_svvh_generic_type of MAN_WRLVL_DQS_L : constant is 1;
    attribute mti_svvh_generic_type of MAN_WRLVL_DQS_H : constant is 1;
    attribute mti_svvh_generic_type of WL_CTRL_L : constant is 2;
    attribute mti_svvh_generic_type of WL_CTRL_H : constant is 2;
    attribute mti_svvh_generic_type of INIT_READ_CLK_CTRL : constant is 2;
    attribute mti_svvh_generic_type of INIT_READ_CLK_CTRL_H : constant is 2;
    attribute mti_svvh_generic_type of INIT_SLIP_STEP : constant is 2;
    attribute mti_svvh_generic_type of INIT_SLIP_STEP_H : constant is 2;
    attribute mti_svvh_generic_type of FORCE_READ_CLK_CTRL_L : constant is 1;
    attribute mti_svvh_generic_type of FORCE_READ_CLK_CTRL_H : constant is 1;
    attribute mti_svvh_generic_type of STOP_WITH_ERROR : constant is 1;
    attribute mti_svvh_generic_type of DQGT_DEBUG : constant is 1;
    attribute mti_svvh_generic_type of WRITE_DEBUG : constant is 1;
    attribute mti_svvh_generic_type of RDEL_ADJ_MAX_RANG : constant is 2;
    attribute mti_svvh_generic_type of MIN_DQSI_WIN : constant is 2;
    attribute mti_svvh_generic_type of INIT_SAMP_POSITION : constant is 2;
    attribute mti_svvh_generic_type of INIT_SAMP_POSITION_H : constant is 2;
    attribute mti_svvh_generic_type of FORCE_SAMP_POSITION_L : constant is 1;
    attribute mti_svvh_generic_type of FORCE_SAMP_POSITION_H : constant is 1;
    attribute mti_svvh_generic_type of RDEL_RD_CNT : constant is 2;
    attribute mti_svvh_generic_type of T400NS : constant is 2;
    attribute mti_svvh_generic_type of T_LPDDR : constant is 2;
    attribute mti_svvh_generic_type of REF_CNT : constant is 2;
    attribute mti_svvh_generic_type of APB_VLD : constant is 1;
    attribute mti_svvh_generic_type of TEST_PATTERN1 : constant is 2;
    attribute mti_svvh_generic_type of TRAIN_RST_TYPE : constant is 1;
    attribute mti_svvh_generic_type of TXS : constant is 2;
    attribute mti_svvh_generic_type of WL_SETTING : constant is 1;
    attribute mti_svvh_generic_type of WCLK_DEL_SEL : constant is 1;
    attribute mti_svvh_generic_type of INIT_WRLVL_STEP_L : constant is 2;
    attribute mti_svvh_generic_type of INIT_WRLVL_STEP_H : constant is 2;
end ipsl_hmic_h_phy_io_v1_1;
