`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dgDqLmra7yjc7A09HBv8jTWc+hwQ6ITXdJ+PaXnw3NX3VhqA0o9+dWgl21Ulfmxm
dFu8fre1QIod0q9gMbj/SfBtljKYsQh4x6xvPQqKyZahrW00a2IdPpOkMP8+7ZGN
TYI+mw4BlOKlPi3OX+QMxD8c6hbReGLu7iepXF8w1p4HyF7y0ClJfJNyet6L4hIn
gfZmswV53ghvnYe0tP+tqnTavHUl1A9O9G+nq9qnWJDK7afc1TDzeRbZqQ7MgAC+
H2C7/LEuIH0uW2/gnZz+R8Eqc6kiDcMMcxSAzLKgN5ZkHox6BLYD+8VKCPGucJ/n
k6eHPBSHeUZgiAm++B9JltHMbyNKQP9e0T3Vo5Rho7ctoqbsJkz8oVuzC1Zcd26R
B32IVfnNPHBeRq4o47PjaQ==
`protect END_PROTECTED
