`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NpDNPDNmSROXPKKwMXoIqVqIRYPFQ9Ei553wppnCkrT8eOo/B7ptmqeM9Dwy7i9Z
PkPtSzNcvokZHN3u/8KG9JCQABXzAMZDkKP2VaO0ohAWc/8NNsjDzgURRCxwHz5v
2CP0i8dlS+6zK8pqBuOyOPGmkwuPppWvFxBk3IepjY7GySvdxk04PnhQVJ7PgRXM
04F/nUd15tpZSLhoyCJDUjXWkiWFn4aiS09s9l8SmZqPukt0va8h+sF3vHC5fRNI
eDhIW94bLs0DnBTHw8QP9EfBUkDUywGj+v416wWegZF3Asv2d/DBl3JsNsoqwhzq
npkj63QSolOMkwTWxH8xwrhTj33/cUH2fFE+/un/9HdQD1GTL9Gkg7ZYAUwY/SBk
YSsJK7T1DH1vZqfANeY8NFnnDSXbaRyZU+9cmrabyyWQJC3m2ZEOLzIkonHCRXjE
jaUMUbC0VrZPT2O/0Xw6xYVjZ/UZCEM4YbPwoY5eXlXYtqLvYu1doQXXf825DGIV
rvVpbaBk4uxITfni6xPRnPclL/eGZGpXCOaRVKaPg0EMMzF4ldAR3VXmo43XKKSR
TO0+MItBoCXtEftOqxgR+ghyGPFMyX6PNd8BSx4DZgddkx8RDNXLC5HcMy4SoJJf
QUbgn/4EuF7YLgHDbI5fEtnD2OHt+KinMBEVOG4ImfnzLRdGnB0IYGF+NB37cdkH
yal/KDkG+YDGpaFk0i05i5LF8anQh5vvTwVCbXFLkyqzz7ENLCbTCCdHCBuC0/hD
TWt47+uPMT2LPxW8VcQzmQSELehZCuaheoMxLsjaCEdQ2qIKzo7Xje8b6xhcIaic
wY2n5NjZLW92Cz1oGUbjMnMycwk/dheCebUbjS2l/26TKPTrk0+icAq5B4ncyTXy
1hqBekXdrg4fOb1S45IqFXSafCBjURcNP/SJtCMmG51pyfXwmkcl2jFA3K+Tp1GN
OZ428293m+Tk77C0aRhIgQced1X/OBuiBZ4UTcwl6dalLQ+1zqASVfL7FsdRoiDE
6h0Q8EzNcaDbqUAx+36aPGoBc4UECi8GjkfGZof73SbWKd8Skr1Rn+dumjjIQYD9
zgsMMdCLpmJNh61+1VdzCG4j/7dp/4UNXcZIZjRxLCVqwPl99vf21Yjia5CjadUl
mioxv816lBKVeaYmJ4JTxecPyaVQLMwqsTgmg93B0k6pD14aDxBKu8lYmtgMfBHM
dGsNaGur+w0mDhyluOzQQgnfTAcHORZ4bB7mNCA3XZQNrvC34tRpM55nFiPtP3ww
bajLgIt72ooVexrkTj2xqxBAnB7TnMDy8C7r/bQzVsSGj1aAEx3ZJ21xXsNMch6Q
VJh3cqLi2hH2odsTZ2ZVtnegcax4vzOmM2OPYw9Lq6MevY5/z/odmI5sW1DdiQJs
ldooXqSJD/qd6fo7QGEx7E+Zriva2B8jaFAU8pZWuCI5auMbF9J9Me3ltVEVyx3x
AnPcOWclwyLv+Kwu8OZYRwE7I2f6KKACa9qeR4fw2NM5e3tpbQGRseBQ1K/MiMAu
ASmCObEubYsKBbuVfs6IytrQvDoBtaJMh5lRywPV6irgCwWhG/2b1uHcCyT99AlZ
AcHbcAXxpI0ShLW1OuOVgZZFnJcrn7DyUbPsbRRIO2ujcVkFZHadmuC4e7Q4nu4a
M77ZW+Wjnt6/iqVPcZEUfXWWDq9T5l3PDUMFG92ERuaQvBpPKOGH8TWwT8BnOYmJ
ZJ16WrI+0FznEpBogXGiFZzEQleZogQS6T2uOdse2Vjo8sUmTFJXXXVJdP9S9AR+
0yb7IVHZDixlko3DEL/vIj/zgHwddiApBRRTwk0YZDb55BWBbsCFn5AbyYnSApGs
gcv8d/EnxXVE69WSMRY3jzm2IGjD4Mg5uan6LDcw2v72ri0KWj3l/PUwy3uzKE4+
qI8fBBOskFFWaK/P296QEyqUFMAhkX3XPidm6/Kmdj4LXWL9/ntg87+K7Flb5yfX
B2V1CzkQ7rt3VSUtgXWI+tnjhmhfU1zOFIYxDJc+QeC5kN0KAmBAhBeOnuvGH706
6nuO1Cj7NqpVKd+J1azdPtnDOf5AqJUJ1Bk8Gcc1YZFiFXue1mYHnHj8dVazuwff
x1CtBx1C8fwvONQEFjajCeIM4pHK+Bhn00K98lf8eBYA41OAam62lXqINtYQgVQ0
4HVMmbgWRDr2EnTgjtr5x36GXwAYj7e02JniRW5y3VMckjSb0Yd/h7NNGvRCREMd
8biMWIaw5k/uukqzvEVWUcZ2Za2eGRfr58fjWBepXUv2u60+q7aidcAS525YxARm
Xyaf3wF5al8+GAdFjhxgCNcWsHYVy7OhCpERPQsNdhvG6Uyq5m3tvtvIZpokbThh
5JTV6OMyijVve+kKnSdxX6tatT8OnDX2umlT2ULeCdEhkGZNvrtxay+n/B2F/MbC
32subQBZvnRthRJFSpJDcDOCvXpv8S0odsKPS/9ikCwpyia1ey4hFO1Zhm7wfcwh
Kt+NaTFwsNB+K1cYt9r4hQR3mfnJkUyb1cFRZHhlYBr0aiLopwcieT0RPMu8x99I
QaN8qBfAb5uNorIKwoWFBmHYDy2pr3ZplmYRqt+1o+MBudWVd5Yk5o76hXEu8Xvg
h/4UNeXD19gRFZm4AnYRE0uamgbOR6uemPTF++zvC98nb9F6aBknUlsgYvJ1LjPv
cQ9V45ulzZqKLJ6GCV/HhR6uJrDTDdP4TO+Z2C3T+ze7FruEMmRiA60ypzIKFf8/
3XrovyYjkh3d8lc2zSVlReZYFeCfRtSrlefqc0UnOWx6rSk2kDj2GXlCF8HaHDz+
75x29oMH+KNW7Q1hoalMrb/elpJOR3z64FTAL/u8BJJJzAa9X8upd0nAcQ7s2A6+
6JhROVVq98hV9+MjSy0t+Rsb6EGRGsyR/VToVJfc0N06PPaaNAUxRiwevLjx5dJ4
rI1WcLB8pf8AkWcx0vtUs37CHDtiG5Ko9pgYD5pV3zTnb72IxZXGRygxR6DSJr+X
/suJZ5Wr3rBqbGiUREkP/ojsj+hU3FzMu1rj0mTrN46OJElxkOuuYZsSOEGn+BbK
GziQVE3M2A4JVdT0qeOV7CsfEX83GNMo4e9c7S2eUynewnYkR4nKSblbl6BnjZtI
A/eCm1O/oGrLlF10IzhxtZhJD99E4Onm++BbUrgnnalNO5qJs4fPO57nH9dbAGDa
k99Oth1uxUZ+eDR/z/0IAKxacvXrwUUwHTgMI7V6GYG9KO4oViHxGO1c5YpdGCwT
4/1C1FT8BCQRoD4i0BbFNmsOijdFEKXx3ogwCd4XehpSfnhmCNMI2xnCiRyM8IFc
MB8B8sxdQH5Pb4mBEACjeI6cKKmP8YlcqvuArlQevcn/GyotEhW4X26BCW5G3T5c
Cuws2K42K69AdMch57LsDj0GZeNEqK7qBp4eDmkB8KQOQvFrjimaU273ApaWQhRs
cYgoOccD3rv9/Rtnbc4txKovLJ+6hKk4TYYZIFoZIlJGtfRNZSnzXpV5+U7eZm2l
W4+o+tS3RC7zdCvNAzyPKp2Spv93uP0KM825S2YVB2CpfT3RU1orOryykJkT+wOJ
Ry2ppX33JGoVmi1icTYOcgkMBy03F7NfxO/AEczLqNA8ykpAIDEKMpeDyxk5AZLb
pNc+Ta/uO9vOw2SQmu5KB0lWtCDLW/S79XrEjdPnJH0I9S3XdIAbvisg1Nle5lcS
N4E5YmbuY80UCaAHZKhyLIqjiI7tAo1gyC23/bCADrvRVI14h+nByiyQJqiNpMVy
bHgAlxjfFtav6pNT+RImTXIcErFe6RIVTnvKd/RejOwVII/a6rgcXv+eFZT4ncEn
j8OhUjvSEpve1s7/PsDbKlFKhHI3Ol6c0ULAdgfNs9bXcZpED/rlKjcvRLwRsx5v
4xOdjyxWrxXfRZKOklZtXwjO2vdOgQQdcFHC85ydFMbwPeiwhsLJy6af7SH+mgl9
BbhlvsEm85dy67Fn76oe6/cwziHM8CifzHANUzEO2peE4L5SLM2cwbMVZGHjLuDO
EihLwxpGuIoqN0GsFoosKGI2wovYHu+lxtyCx1kND6Qqx4OldnLj5/C7dIc8ImMp
vFClw6gmqrsU9BQK+PBc4Thdmaqx9LQ8Uiy1RRDByvm/cZJ6vz4z1Rgimv7jhyRI
xIQTlcSL6xqRxpkT8mzolydqTpo2EPyNcwotUwN15gwiJLRiy2cGHIVgKz/Mdve6
6L7eDhy/fOU1FZulupKipMZy/JCMDS9gydMa2/sEa+0OxZbDxdx9qgq43jjjlA+4
XyspQCmPmXozIqPI2JtNpssVqOQR3n8jylrJMKqSFHRkMU8nG2Nx82mOAbgx/wea
E8zYTAjybcOgZj5dK5pyIubnxvK5xOo/K5auzc20WH+TcjQMSYHYn8NX8AekArg1
Y0lSIdjPrfHoE/J4ScOPjvDdu26ORHBHDu/k6X0IVx84SofGg7TTFXOzwjpXza8m
bECgn/f+OuBAN+qjz2PTBCwu3eLs0K80ut1DGcXBdSUrF+/H5mTTvMBU6PD3BnQd
fUGlbiszk7anBp4NRYhnNVm0s1UML0yxnJCKa1LPp0kIVXwxO0CcafsUA/drmyRy
DLjNkhFhrjFtIHXIKpL81fUsM5y5t7Flr7VXFVJm+cXfWUMEQtlOC/UHPlJ2Pp/u
nujrZJ5kdwHrvZz4q2Snnp3AC+PsmtewLwV8ZTAB/wpdrwdcKbZi33/vjJier06f
0g2wKiRdeC18RNwIFbnVmOjJ27Y9+8PaRvNyP6SY5nK7GZ1fdIiS/mXZAP8mYWm+
g5xiasDa3m3Lu9+nDteB45m3Q9qS/vARNw+yKBZ5NAbJB+h5MsEkCvlaUS3i+Re5
k30w0ZuByvKGbD5i1959KhXEBrBFp+c3dMjejting4mILp2OMXbDSlUDAC7v7m+f
fDl3mQlgPatc8SXLUeYXo1v5v9vqagQOu9IlafuMO3A0vvgKt50N9p4Rx8LHtKpA
cwKiJaYMxQmUuPXmwKvqkM45moYoJP9nVPnlrXN2M/tRqMaI3c6H3JJlTRB87DT4
EfgU+cAMTvFcHmb+4h2+XsaNXFCTQv33CWA9NgW5QtdDlyLvq97glCQLTWTpARFg
CcLiurZaEP6HuTBxSKwg52m0EI65+R+n5FAmlPs7UN9G5I5A9A4jS+Z4AlIuRfgW
lxkVXgEBY+/swVNXtEilMEmzbIF99pgA64v7o7gSbBegw2Bmt1+oaMZ/tZ91iIcn
XuOVFEevX8fXBDAyTq2ue3ePVIjLHa2ZZqzJCPEuZlmTbMlIh/RDpai8RcMQ1AEP
VWc17aGKCmlceZz7XUB/EAy3ClYyG04a1guhapPXaGgX7aDmHhQak0F0dXL46CzY
n/QnuK8bPrjiz5GdyIXeu6qUvybPVX0dGVknRpXpsqdXahq9xVx2qKgDZPvJwyNP
vdy4lDLqQ7VzXb5/QSQyT3FGSrg9HKOIJJBNB84QStg3h802giRZ8dlGbvOeDCwm
5+h7EuAHuEboOI0bb7A5bsK+zoSx6cF3Vc/v533yoQBLp5okbSr/7iz98xl9CyWJ
+8i9abUGDOoIbKFafq++uRetWRM8+zQ5/PGeblWNM3Fz3LMqZc72HmMm+EN4CORk
sh31K0tJM4OXGH7nfVIjdex5/XFsGXbAr+hnvM3Ji9xMjmqip1X0Kb0GXlTgxlKO
R98TrNIAbjVh9zeE7yPkEHwsOi1Msa8Upp1VsHQqJhrJnk0LRKg9mQBwFPhkY58N
lhEhaUwmyTLfr1fNsHETDoir2skZT8bw/0W2razwcJqvAx2Adzzks1jNhhMIEp/a
yZtwocU5nfoPN9XyA1abgsw2vPfyBNyxFG7MOVHiGDzL9WPDZmDVAZJ6FFuRTy0g
ocjWG1WNbu8lLQL9r6O+UP9kdd/jwPobZO8aJ830nSSaaYUs0wrkQAhwvs/EA6dc
BtlSSu5FZjbGw0fJabvyUxnZ22UlayYhVx5PkjYEVcwJ3KWfmtUzbGtprV0tvCsP
O8HPhOvGRFEdfgLk2X1k7e8dqTT/ldjwXNBhiFoMIJJicogVg+Po7S44HCZMV4mp
K23L/Hpy+BqJV3axmBR01Y9Yvyf6W+OTRc/fS3Ahw6Nynh8ypRf/CFqwqqIVhhjO
UIg6bNTeajMH+ZrAu7/RC5b+O4MLncA7ciaNFigEKOzesjTWWymokwV0IM6GI08w
TFrIU2NN6s9uqYnVL67sBRjnn9itmHeiobAP5y86y3Ax23zPcq4oohRONh27PBkf
9O/XAWx1LhZN4BWj4hqjqRIt9S1fFgkRY5bpzRWSCXcaT38kVgvD3Bl85XCVz9pF
pI9rGUxFNbrZ6X4xAA+h70bzN4Cym+W+QUmGEAmG4OGHVTOzcCkU+Z1Wb7TARnbC
5hhbmr3YrtiAfHjRAqf/QMTUAR2eDAOOkCmMQtpqb19AmglPxcTSpHW8dd+dVyP6
AEO0R3Ua9ZzetptdOC8f2SiC0P9o41kW3ChBhysVs9t+EOduuR3WjPbofmucDQqM
Dxr6UiD3P51pW+so2ho8GhylhXgTZEyRvb6/0Z33qy0INP7JLa/D9qDMa7iCu6DC
KFUSycfqJqcBG0XGC0TA19Hu1jgh8dnZtD+y8eT5Tin3Cq3InsOqTduVKiiy6f0b
H2XTQRuHFiRzRB2Bt3OYSrEKmFrBcMXpk+chqF48j8ZPZxVVbO5R40djA7zJKmva
wgf9HzA/XRyAa7npxpQCcZzBguy+FVraju0GHurzTPNSfH6P/ZUA/SRf2NWTW66H
ezpcYibJEry++MZZkZsvauLB9NL6kI8BrJWRXiR5+O+YsUT2ju269YDdbqqZZyuE
jwD238gfQGPD1d1+PPK9ryyPedLiQo3hhTGw9pxk/00kJMR4ZzjTODXnknhVzGff
siY5yEM7mdCkKKW/ve3fbVdIFs9kgiMmZwque4/BBcV5BcsIItq8oOIUGQiRjMCB
vttgXwu8+OziuxBWzknylTI5aLZiugk3Rs9RwOq9FG6kt3Jm1Shs965I9+CXYBzV
mnmyx/vzzpmzAAAzV+bsgVD4HwmWj6j6N4GjzC8+WXfk6zcE0c2ieVWHlr5wosmQ
8GNlOfUjjufP3ZSphss3XX1c0sVmpSGcCArEaPyMvzZ/4UYuylWFff4ePZ0eJfld
G6ciYeKLWltL2/DDFrkiCOYcIveFUM2Xj4XYRF+N9I85w1zak/g+nS5swFBB1e+q
w9+Yrl7uYFjsIj5YILdwBZKVauDFBh8GsJxZKfbAUoZEYWtl9PSbdzoCOmdMtgIE
zeJ+7HqC77fTwOPy/shN5YWDHS10iofpfQr3491Mc5OXvljUfsa4KBiXuHaNui9Z
3b/kq1Vc13A9SbvPUHO5QgH6t0eH76rRa/vFYQShJm5LcuNevK9z53puRyreRP3r
YYEn6LaelC/eDW7POhJLnPASDwv9uav4zP+XY/XxSvKKl13JVclwVNwYRAO5Cupf
rD00AMiYL2putWGn5Q6mp4TU0Gt5mQKRgAF3m5NvugAPQ74KoMzMKstYCDMyXJTJ
ufTw+Qtrdn67rgud4rqbfzBmjHku7zmBNSJJZHhRnu4CD2w/H5mcULPnrO/dfvua
2eIgx+/ra18Bu0nEnQBcoGHa/UR/Yvik/NzJmT1FfInQZ0obFgPrBU/boUMMdIVn
T2hU1V1tsp1p8KvhesSSXWBRST2HkECKYg9zSsr5CQcBpd8sQu1AR1KzRtnzXS8n
ujGMFEPEwltO8NpMIScBsHZ5nHdnvFWwAtO45o7ZqBMdhKV0ctyAan0Cpfb7gYVf
hmkehX195aJi98xoblCXZrOi6jGb17KY2Dpo8RFLFj7KLMDjVhqmjGIp7x+ZzsZ6
giEOo5HfayZFO0Dmul8Xaf5Uvcxi0vqaozI+musoIsdPGcbKYNVeX9xa3d6dvryz
iZWue0rk54J38qG127RcDqOQIShldt1zRev5/viPdnGXljo1Q7e1Hgp1ArNqviZV
+kNwQfVictlNXSZ1fBOVc6wucjcsR3TC8Z1c4Ffm8ow9S4p9vAhORgvFPHBSnJkp
nV17wzEgTCMPAAMRyKaMaLqYaqNN/VCCsfTLtUnk+i+PYFY7wIv2rKnzibsq8opb
PH2zvJQCMZRFRVVoCIl6XyybjgZSmc0799bV3/wr1HiKpTVbycgnWI9Rhrx75KAr
9rVQs3+o+6ZEbeIUEg+sCmxfyZERxrjN+uIKPm6FGewKQaAfjEP9pRUaDfcE9fXa
Tef8m1wTCs26/PQNvZ26g1CF3RsUMN4dwMrK13X+t9/6asBmn9SKuOeFEDJD+y/O
4353y+Sb092I7D6SDRSCKJAv553i24iVTbwsuNB81Rlne77suKP5G+Niis5m6Dkr
dTH8bxX0QARNJS4UgtARaEbXIWm2Yx0Lyoj4d5SlcAJxnwV6t+LR5KSNgmJYEvQ/
1dVkNGhfQ6OdbvXsmJeFtOamM1SBTQsgQJcEcwX69yRfNY3n0RTzTQUGUrkIuWKT
PkB1PFzvlVTyi4Xyns3kwHHxo5NkV6JJagNwHodtREKLIibP8Wx+yu/Ns7YlQeuk
Z4Vq2GkZWeyDNG+GROrzt8pl+t/1CbjsUUq9HLqDd5jPCbNhehGr9PkO7pzWG9C/
2GWcP1U+EqLlh/K5t+eLxRX30EKAy4H8DktXn6D+VNN1vot4Wo2fp0GTrvjH4R0N
EKwaZQqflbtzQ5C2VLHVW1EaUxH+afUtxnh2d9Tgra66330vGkrBA1YqGOL+thtO
adv6a0slin/gRsnm5uTWT92v2PQF1SZi/hUnNT/UEzKvoB8KIWnrBbPIKwJc3X81
+B2Afw22YfegN3RKm+NMZWM5puiTaRN4tNTk1x01T6ZeZjHNww48IKwU2IpaOyNT
TuFKUuII7lreHE+AkleOyh6UYvbovGBNqASxok/vlW6gtG2ITI80lp0c0yoYqybZ
IFBOc8P5IOdUGHQMOMsGY3soEUb00DAO6rP4xfLlb+5FNTWFoSUchGWBWT8EYBdo
iay9CgjUMtuF12atjU8SLkmmKnOr5+pd9ASmgc8bCtLmKkU1wU7ik2k/0a9oBYDS
DdJ9GlpBX+tBPlnEeuFRAA==
`protect END_PROTECTED
