`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xl/N1BvX+Rq/bmtcFDEPfkTDjytGIIGlfvhhqZmRUg6ODE+rXpEXDi58tB7dLbBR
AY8yzAVO+kBFnn1h55dKiwsSzbd5YXPPXdz0FplfZIfhhrgjLWl/ZQb+c1q9zKDA
bl9DdKUq4GjnIQZ9npZ7Cft05usGpsdKPFdZLDE+HF/e2okbJ4d7fucEIUSMnIAq
Aq/a22VsPzV1bi218s/9/qk3qCkQfQ4B6YjLUl+eS3VWY8XGkp2qitt8MBhcDowC
1GVIsPiuxHaKq0dInWfbgzczbO98s1iDQo/QXWvlmVZ29L33G4Ged9Vd+PISFiQp
dZwOhoqimZw3Z09zxJCOW2lhoMj1ZsSE/pdWHlPdAh1rg51s8IUN1TXjqHDv2Sqk
/CZrFgzf8p6mLx9TkhhabrWuodncyS1br2glI2E/V1bZMVpjqno7cUsBbQh6dLh7
lqswGX+mpXuTCfUSZ+M9h0nlHG5qmwJfFkO3z85qNcBhYgkaHKszsZgAdFi+7puz
WnyhMMOFCUlvfyeerJ2vSTtNzJ1EPUPLrByOBGvXWr45HpwpFdpU2nx1voLJGMcj
W/dO0NRpYzZkVzrL3pGR+S7KnPXznRs2fIQJBKHT6ACsAgmyTwoI0co0Nif0MCmn
4FiIH2tbnEUmBQlHHamERKaw/mW92AVMGTzk6Hw8ed565uzc4f/t0UVSZXkMlSg3
+JiN24d1tCB7fbadAxSLF/+pqAFnkqdq8VLlYgJvXo29sdcFIzvH7n1ZXbyR9mxE
4c39cgZGJPq8LT2q+83Z1B4wVQa/G0p/TQcN39YlUJCH1vlsKGptUk/FhlrJ+y+y
j8zpBZChHWJwI4itzfGsqNyDegkt6DZrW1qZ5J96UZVuy9GTN+wKERA9aMMNvR+/
2v67keoCPunHIolg0G/39LNqZMVe0M6OLdgUNqB41rr21FLSPEVowxs3xMo0iUqJ
V3MjOHly+/dx21PfXmJCMssRmAkduk+cpPn1EvX5LcQlQUnU39QkZB6eOnvqazNO
BwCNpciliK0LyRe6SvsUBcJU7uIElDWrGq6dKHlOdQto7EpoxlvaQBJNtGyp7Kp6
tO8MQCWhxaPlsTjn3i6U5m10ASz9p67Tv7dfo8fjRoUSMv+mfLsXDnqbPzgXYG88
6fcE6NpP8dVorQLPmdKeLnB8lw7jUsIDNE+voMbhP5xckP3ikpkzy6SZrPXNNQaj
RZ10q4aYrORzue++oF0DWJ96w8YgxfEkJTqbTIfZXqyt9acDIEe9yEo/+7jRnGNT
MCQDSI8BSYev2QsiEG/K5CmjKtxYnIFfgxffBTMDHCPhnE9y02oQVvi+tQ300h2t
3R/7hksDd7rQ+JEenylKagpZMhW70vDEnLHbxUjdts27g1B2qzJjnHw7knbZN7Pk
wOiqJt8kLX5Tves8Kw7xpk3WPfYzCT5ysuk6i42XlETR75V9oR8n/vnXlSVgrNTA
M6cWO5OUYkez7DGjmTOslR6U+BygdiCVwlLwc2tLyCTDGXCIzjwHthD2GckFzHHM
q7+MYZ9/r7oZWg+JCU+My9bKWcBdhfYcNN3MHNPiX84xUxIpuVfKba6DC9P3fHyU
kPp7Q+TtC/qpa8fT8jRXuM3DM6P8Eg0iigQYHVHzz9yrWi/kLvcRVG/93hi9h7hR
fPebAdmOvaAn1zsBQJOenNHNAj2edAv5l7rPKeIsj0Qlx6wuwAXoesnbvyqzUEyw
SmY6dCV3zPu5hq56FPa0zaDL2LxvK830VUh64MvHFKMQ9tx79w4LuaORisE0xzIk
WPwbx/GiInkBudfhvfniyRM0Dbt51mjsQW5xTsfuK8TOnqFBJU4K6SrxXzOR67Zv
0qIUnktplhMrSOBy8VFag/QAY3yCWc4K2Fv2sx9RduItp7IWROUz/07cILxOSUCY
Hr4k7ZaLCIch7koGH72do6PEpWaKkyr3Yn0C74/nrbFWC2i6mONWQD395qWYDtw6
UhaEFTEFMNHHmkXDsABMIDNDAxBVB0jg5Bg0RImVxbACp/V+jwjnij79fGzJ/yqD
BQRXAN6hBTmQ6lL3pSfX4REZm0+yMjG62pc43BQzZz15fZdE+Qo3nubPYTEG6hg2
WJG561MDmOWQB7FeQOFlHEOP0jLdab2BRTwslqSQ0rMBI8i46fI4H/IJzC4zLkfI
HGhiITFvmXB5j+QYbWroPX62nqNNX9JSRHgFHfP3m4xko44NEeuHxdoIcJqRPCsC
7w+7QIENHi1IiDKzZ3mpIg4ZX4l9KHfJ7z73pgmxI5bRbG+dv7ib/VDOw3v9Ert7
KxRrS5uoYFsAmVNz3cysCpo/ZYmsc5wR1GXBZRraoXjMDSRYNoK7U5WjxgqE7YRK
DvbrUhNG+Z0mEa4jxxVv5nP4n2bgIPtTG8569EhH4wXEt9WTgNmBvUPqdjeAmGuJ
nDuzV0nKaVTc5oG4mvwb0D4eKpZpkNbHDrcJIL42JGjdaQpq8SJZqX0P53BqhGPT
KtO2rS3rimcr2Km8lD6G7ENwRf90goTvASq37bvo+6NPEvskxru4EdZRbw6VXnhu
7hU7APdIcbUX3LSw4zAb9zvHz5ftp4g3NX79QylObyPm5fUkRzmZdwMpfChB7bxz
EHlO0MuIxWcPA3CEGVCfaYGTOonXOtBBrVOAHrEzuZBc4q8YsVyUDM4StiqAy5Lr
oMrkcRrYeWbgrLGd+B0Rchkw3KOD946E9ckEtEpXfxIjV7fx4+104fPtpraCg+dN
ikM0j/NNcSBzfEV6xEdjPJjdjWkWOo3oMBtkDH7drtIFAPBuEZtpuCTfDMrlFco6
EiiIgV0O7SiAg/yv4Ntnw77MFPuGCabBVhR1Xfh3uHF6vFzLIcBFvMJ/X3VrVFt/
teR2QUl2kHHK3Ld27edZ9k6CQAVLMIFS0z7I8MYmJ6B7estHqbXqaBG/apgQgD/Q
YTSeBFZpGA6bQAQwU2cOuapstLHs7bsh8Y87FaJnXNGrX7jHQWS1SmhKzBRwg23F
AZUfhXwtAy+18TGx1KAHxgYWQqqpJ6KArgMKONXYmywt9t6bw8GhGh2RxDIKTJke
sexsdX8tUcla5P9kxIoUGWN6Xb2geDAMpP9YeDpMw6ZhTuyT5wiGn2oZTwAxMCqm
xMAeVDgx05NceN3oDePREM4mpVF3T+rjZ6xQjKFcfDKlG/Hjq+NVhAT/en0MWYnV
/ib7IAvEI9PQJW6YMngFWGyCGmuaYvH/PIxWAB0hxJoWLKyvqrZpHgksnU96KbN7
hxLpLZrWNuje9ywASDNcXm2KVayfoXf2doAmAGJ9C4p1wRSsj/ltf6v9I+2nlkgc
42vlCuyXvEfcuWTps7Yr2JgyEZgcThr6q6hxl6/O4kmBeqGWZ/2epgaB0shzZoTF
Q+fNrX1cY/0mbsdLbo1ddIoEOQGauMSR6LTNpE3vOyp10B8TAevO2oZXLce/A1tE
b2cOzh+KMurV/56zbJHuCqFhskp5erTUPAwTsxvzr4heOgSWhMPSI9IsT1XHrhG6
WsVRcWCEaZIemGRiyop2JTzxX0dWo7svISTaV15099iavJ1nrBPq7IMrEKoLSoKv
R0wpcBzp7zxN4vUT+R1IwN7Qjr3BqoDsDRVFlHnsi3iLzuzXOQDmbiCNIPBwKZ6i
/OSUG0pR5AOt4u6ljFu9iXhKcxm1CUrTdTxEqHwVTc0i7pyfir9WVCwfoArYjWA8
u37wQNy/EVScN5u6Anh+gtf8ZnGgb5TawzAyMHnOguw6lWTvelO+aaab5fbDY9AM
p010DeSweVfHZ7PGnC1JRQS4OZUMwsaTZZm6K6Xd1WqFZqdPEky4l4uBWm0ob59V
xiE5587tV6Hu8AGoMri+1ISWFg4McfJACM40NVnG7Kawllp7T6iDKyFdUHaAl6N7
lxPPbXmXrkDvoWFr3Vs07eG2Zq5rRJZXw0jdwg4qVDI/t3usBxa19bLx15K7Ss4U
9rPLU1HvyHGg6VbHrGOA+2JnWAFVhVwmq9EZVjAhIMxgZGhl+vy06YLbRJDg59XH
ObJIZA4o0QGkudVL3ko/yNBkSqcLSjyT9RSisy3/8ljKu1XyRTyg5ggdKoOjVhku
mUwwsLmlqsgeA/yz9XoFdeeChengfjsDOra8w1gEdlwAcxvS3jMgWSuD67HmLSCq
CjjNXeY9WV9VIbpZmAIl5u1FMI/wWUT+JGj6sUCVhuogvaMvZB6ntTtLtLWa30sH
O0Rdrr3so8rWzPaUipQchrzgBZwsKqdSBiEZGjhrnEW9FbxC4QP3yeXlDLo8lc8M
7raZ2AuDIb0WwZd2hBh514S2jDSBh3CfdFKQbCRYCEoLdrCcc2SG5r5wHypiDOE+
qBay3j/U2XWgsL9eFaGr39MW+5yWogtuX/GfBxW2LaDKYM5HYaHvV8jkqTFVL+Sy
2pQq8+oCPUrnfGdadjtxr3tRGYYsK9kuxSB0igAR8uwS4cDA2fpiFkwToPhkOZve
uPq1WhsMNIvJOyR5Z1teTzv4lFnHogeEYVTDuJgbg5TPwZcFUsqQXfD0stXG75N9
MF/EASg7M3tw94bRugDwH4SgnaKZpwykXt6Iz+VOK4Pus0h95lpOvNybr5aiIBiv
lMskPT0EhUpR8tbHGe1TxRisUld4/SjH21N+Oyyoqw4Z60ycuKl54SHJS6UXAhUa
vjcV1Qxe2BDEqX3bhcqR6ZYBgWhiTOGyWYB2c09cl40l8tS6pZDhfdaOV8UIWOQS
qotDpGIsHplLXjGJl2xVG9B7NPV6xGtUl+uyHeQ7PO0lh8UcP9eB/kmc12Yfni4L
yVKu5rSqqaPSJScFxDUCfokL6CxDmBV4SIDWtQzrittu68XFleB0AySlApPoalc8
WWW2g82f+QpyVbolj1zpg6/ws6QtRaYSXRxO7MdB+5FjbjA60Cf8+pKVUIQCnebk
zvXY90ckiUauc/USSO6zbxANhg+GQkH2/OFm5dkXeIwNthm1pWMdhpVmCTwMhV99
avl9NPiipbZt84FS8eQ64yxDi5wpBdrA/NGMsNOfJQP3v37sQmX2iOFGX2uJj4J2
LMcP9pKpOfXAbN6WvOazWAubbdAAP6ukqfEGc/SYSOo2FlgL9w0hpLdYYYZmq7uG
o4pD/oACgiPBwa6lDox6xvY18tGnmcJQ8ZdniCJuypGqz7J6cn0eIz98GXNZrZN4
51AZNznnzUuYY25aynML2plhBonh6mdZ5G/76pj4fTLvSXakuSayHREE9iYGzCzG
16d5ztcsWyC26SC/IzwXVti5TVXgw84LpAeryqQFVSn0lx3QHHiuLWqkJQGqfEHL
Glyr0xEgIJEpvHfS+qpp2ucSYKwL3claTtGy5hDiRtVAj3vXvtNxdXen+TdnBcQH
FhMLuxr4Ksb8Y/uDZwzBDdyMlhRyzC5Bes0krR29cx2+Sw45kWYiTcEDlnRDAtQD
cemgNgb6v0vhnp0qH0SbT3QAtTwqYteCeBGUjnAIFIKPi/iZ9bewJTwhR13I+JoX
ihC1bz7HFmNKREd4cOEBjXSVSFgmGbjomXrsb1uSzhPh0Z5u2FH4aRxH8xb1YivJ
FkyNIWO6oFay5Z15kAsh56SNLx8ehVIEQImdYU1QPWYes6tPLvFT0rZWNT1JoNSD
YWAbVtU9nFcD6UOvDMCP0pbC7lpK07iJfZnZnNjrXnH/1L9wyEteV4bJN1hRr7Ly
SD3ybfZIEQm4ZWyNq3X7eOT1AEOvlXQmpf2Qh4u/xoej4LgdlsIbc6Q93fgEI8+2
XD2NwhVU+eibBqS/hRk/g7Eeye6BwFL5yHxa+jHArfE2HCRWucza8E167JWM8ine
p7HnQtNgxtHTEQSR0tnMM9NixprHvlBL/qopa3KEmaHFJDRgNs404n80LtUPC4vZ
9zRT0TAoxW5pgp4gWnmP25VRaqJ97/DedppsDz2NosbOre2ZhmN0w5B9ZUWV8ki3
ZEN8TtNeyvi9zVflM3nIh2Ykv+oV3wMZIkgldcvrRpL2dnal6C9q96JDaYtM6a9G
i6MlNREenzVsIytB74oSLDQvn5wx8Kk6sffFuxVz3UNuk8Gbz/w2MOluLJLiao8h
+sLrE9g5+Brbyb03FtnUjq1cqShl++VP/ZUVnBLe4VNTOL1sUb5NUC/D12w1QRYM
iHAY+HpNTFDrs97AdPuZY/uK2DD04sbhYtXjTqkU53HPTqa6NkSKgfttjUHcGt24
kcN/alZ3YHh3F+lwuWZRx8Gn5hq1X4hpkI/eMGRK/e/hjHsYvy41Sc2b2LDNLKT7
p2maYiU3Ja1Vf9olrKh0r0z9IzWkHiWONpZAQRJipxoGS9/yCVUpC+cgLTwHWpFk
2Dxk51yUhtLuqlyX9u65wm/K+UCxl4jNV9PShEsaG5wUf18CBU12pyYf9aZceotv
yweqwfsyQMcv2aq0YTIj+DDmdYMiOgpkvIW9lwqPv9QyCYbSGzBO8D3OaYlI0flY
RfSs2q3g7dpjuZj50sPpuqvr95fmQBpdOZx5XnbB33JIpOPElVlz/XwMaWrW5Dwr
1CHQDfMZMyoHdJYtFz4HwvE32AucOfPVWGbbA3/22EbYXRFS3ghoqvZTOsrCk06d
p3ePjKsbsfKS+yPqan2OEuPuAYIHoVCfZKENlXjjbc00pvs7yak+hCAvYS5RZRW/
VnsAhMq+xYW1WYkT0fzC985RJ3Qdlr/4mrO0D8wQDN19OPJJjZaSmngyvGf7u8ov
gdyVbD2+UvGbZAxXp6/gDhHgKlFZZPyHESO1o5/NCzIVBOulwpMfj37RTJUrziRS
iWslG2Y119dQ2p68CI4agH8neOlC8TyH8Usf6NCU9us=
`protect END_PROTECTED
