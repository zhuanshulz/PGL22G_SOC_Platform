`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t73+mY88jImxMOzl97g5fV4mrmyfV25SJSWs9BU5ccZyRkQPRiJl4z75EuDZeWxW
4c88dpl+hZwctVzNcQ3S+MAp4w/cldYpf7m/wCYWikrOxQZkbU7+SZ+cf97SS7lY
6mi/Q/Eau09XXP9nARWSET4Z9K4aGEiz4vc5KUcrOoFgEoxDj1xIlvB194zfIfyS
GEf09PvZwYlVbUg3KDvYBa7kq7ABYKo5lo2hA5Ersv6jV8cFNCkPqpW5YtNS/O5q
q7RpIuzrhECLx80CRKwMK+DF7FcqMwCmbkMC7uiD/6ckE0pRdL8ePMcAoEOaVYyg
a4K9wboSvL5+x92vetEUpA==
`protect END_PROTECTED
