`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7mUqZ/mTQ48MHuTjM7vktoHHx4Y/lKm9tG+R+gZ8URMBCVp/xjlDfZB+7OZdHzfm
k5I6cBfpZgEugjPGQUEgKaJPAs6LEVFqs9qjMbKFur8ZhI8ECIUugWQviv4/yYTl
jzyo65Ee8M7E8aKYZvSUqEWzH4t1znvA4Ux6Q2K8dCtl7pn2P5QfwT+MEa/EJulO
DIEfBu0E8JFOG48xaB0AOU7UKzuy3+GG6chq8f2kAuQq4kr1oY2mbHW0Y954YWfS
G+bc9wSnFhZycu1zMvDCvTBRcPxmNU3qUn93RKxT1zmtzU8YoS8IklKay+85N8eQ
Hn9FqQUPlLadYUpyorUESkVjzIcXohyZasHOFFUBAJOS5jYzVndgXLxJsKlhwi1M
um2bfabxtLLuxf3kCZ6D49ckd2Qv8H5JL2ngf2AyrrIDLn9IdUlK/Mwn48cOmnT+
Q/aCx90ovCBxUrQdQhe5yCkMB0TkzJR7wsxKNoWhvgwEp+h20O//fqAuPt8L+psI
UuLJCBOOLD8J9EeZ8pVL5gar499foX+VkZrUYWb5XzQcNRJkEBOK0JMcoTnVG3N1
oNO/XGoZM/0C6Gv7/3x3PaKAGEpS+dnBi5kdRIbTWjUb31e0YAWKQ/vgrM2Vlt9P
kGl7MvxNFrbL+rqCsuHT4sCSqrnBidIhdxWBlofdd5N1Ag6/SCgbhgX04gwnvYkK
7k1FtLt16GJlQ/iQpIR+LAZCXb85SSJwfnIBHrz/PG+JxzGn41qCMRxmtDJvLcV1
HpDzSYtoX/U1l5z5gkFbjvHcYHczF98HGkeqAXj/2+PKZmn0mmXnM46Sr6/Bk3Ff
rcPpRtdkfPnNCZ2n+rkJ40kBdWpoPq9CfFtrhq3PxcGP1RJgXyNj0iQnj48/NntT
k2zvAfWrDCtWY6ToMlVcO9lXlMfp/FHZ03cesDM0lA/S9zxRPLMK9hLWRjENt88p
hOPXscgOXdoQ5XCBN4ah8ANwLE9WOl5JHhVAsUt3yhvkH/kvSaVbnsC21pgDjG86
g7ClJA3aH0IlUUhKYhEipBgn29f2/hiWUny05Uz/VKlY0vR2YXm8eRJEQN5csTNi
XS6fvqYsLIzWHwdW8/8XydlBK8xH7LiwuEZh1AwXLRomk+YTEvQ5BN+lKcfQp3qG
lzAc8b8ytmo3NNx9dzYDczWh95IXmOoPsGQLyZ4l3AHFALNPMsd8NJ8P3wcY0YSt
Nh2e8QjYYabRDNutlf992cSi5fMgZ0rPMr1h/aFbKDC89+MhDEnEO3Y8KCtfh8CR
Myn11+2YLxKFX4fN4bCf9tdPqC8lN7r4l42nfQnpSER4rRgAXTTkXtkyqklqmjTV
paU4xCKd7EuWfxfW41qKdJ1EyuNvysJ3an1uscuztAjH1/o4d6TEgMaUMyml5pbb
oq8AudLB674oHphgaHcCQeXNIVhmINebITGmu3gDSkSAacsOnH0GUsbNHfZlpQf0
TWSTGkmwD0QdP+h1fEYZhXs7YkUKqnc1QlvGYIh7Nq2AHtaSdb75GI58uwVMdRjs
y3EYna9oBmMPhLi2DREshAZihh3P6IeutExcGt1Fes22p3GjfdIRZtYRNuRQtF3c
exnaVVq3gJL9oRPtr34oY7VYxQWRGOPeYbSwOqjNt1FDBDbLuyRkmHg2uddNwT8H
c2fI9lM2Pa0ASEZH89dQwgub4gWmBS4GI87vdJVij2Iu/fM5vCvra3veOEXsE5gQ
uV5D/kF5H+M01qEgtLGUMwmHuISGeeunZe3nXVm49s3dd+sr1Bz3gfVOzFZZFgnO
jIAa/EF1TkOGb7CoFonC7m9kwVtRkrHh+uCC9C9IEwqORz9k5QxcsWICj4Mh4jvs
GXMRy2JjRh+lPhvnPcHBZ2xkcB1Agzum0zYCytRMsact0gcQNyhjeOdcI+dL4gIW
6lPLVf1MkZBDKte1nUr0tFA+k2uhVNsoGTbXlx78SE7RJWKPRJeiC0v1mweD0ka6
1zy9c3qy4qwlN4rGPJkUlRKus1YgthJ0SiQdYS61kESQSHdPS6zfh5+C4mGkXfJP
96OX1uVizuzg2j3BpuqzQycOGKhbB/iBiQXVvm5hUEwwwZdNP3pd+RWinSjEYXoK
P9wBxU3v6FxvUR8P1jFvR9jgPF44PNPbOzMlVWBgb65xAWck9Trx9OdEdbGy1aTJ
gdUMitdvFTNtETG9pk6SWqa/bh6qkiTVSrUk+9/tUfBF5SydRD/4WQkaAKefmZQJ
HGhkktCqilB7HcL13cY7CjqDQa0S8YdkG5ZP63LdlGUbBobKlQEoDtL5KqvYfiY9
DWSL4ns+nhofmLqBjRhEzqINT2k7pV+invYJ6QRJHBhE6sY7oMDIC0sBd4f+lHYu
NPqwO7i4KlPlCR1X6yHYvJIvfXJh9wOQBelLyEPFmF9JrFubfax+G6wpOEM4P78t
sze2vaIzM52g2LlT6QayrOowsJUA2QPnieYLwp75wnaOFX0uHse2i91/GCw/dawn
r4zIxE8Jaj1Q0dcl31I1uF7aLBMmRDFkTd8uzIaIdFk9cyKJxa3YdQBwU+gvjGG4
/r5vV5xoEDZAh4oEcAr42WiP6DgajMeSiGRiVZcu8V63oTa0xSOi5DAIyaUFkIHZ
`protect END_PROTECTED
