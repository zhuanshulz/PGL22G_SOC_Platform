`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V6khHKYbWXwUj5pTCI5kgfUw67zgqtqt31/dpsjhesAW7/P1vfiyIUscqkg6W4Ei
bDT0s76gIliHpU/MxkixYv0UVzIB/rWDu7Bo8II3G9/Z78mdkF5vH+7F+2HvO8Uc
1BoUeYmbmEFKHiLuFa4wkCEBFiF9TTQKufpHLNC2u+WPwrmOgrj5VyRZKZlmVuKq
aOX2N8LSsDPoYEz6PwH4erDjQ7tPw+u3LJyKRXc2b7QL1UVgpINLDt0phPZI6yVF
I8sLgUP2OKcYCYAmcbT9+DSIuYJAbHlYFAgo+itnhZ8lMh5AULrcAVuGUBbd0Pd5
H0fmSaYr9zNtzW+bnwiZtsZrF8RuWlLjUxKLxKkZaSvTy50hRqiwch8lylm6feB7
NUCatQStbuKJfx8f9fh4sw==
`protect END_PROTECTED
