`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s5r0rxuK/NRASjWqsyu9Oeub90BYAyjV1kupCl89zCyZgLUh+Y6omUMgRSbVCAAI
0GE1Pw9xt2o16Q2HVIB2G9n0ZZ2xUjg/y36aPdk9rHZ6703aNIQcvFhKSH+GVUaw
MQHTscG7dMm0yH6kXGGzuy3Up7M4zWRjeS5L9ES1zmy7o4HGsg3A4FkeNiEoq+yf
FXmTTEQlg79D/ikw+T7NWZtzE5dBb2k8O1gJ5uJU10rUBQMXNqF7i2h27YBRh1Ou
0bRvYCvSxlkiKPol3Oyuh9wk8h3oc7oH8iuNKTnGlf1+SIgcwmgAsziyQtjXex8o
xrLy78IG/HwVMEHf+XO8C5CWS6kxju45uuX55bDSGogtb+y8qKU8VYUR8M4iUQ0o
UT8n3bfLVVJCBZ6tWvFHJxCt549RBUUECqtOVBhr2zRVrCHBiA0BQmqxOJ8Vdlvh
Vpz3zWUK4Mn3CUywKZ+HMcR5Si4vS6zwLcNA0YjkLmOLJcVw9i6P9OsN28FkJ2+E
Mx4qzWgldZg37PH5ut8zby0gyA63+3i9oIoAMTQfZaAuWJh+F5BzYJLQ6fr2/R6N
3O9QTiJdgXV90iYrOBaZn29df9ZSo5x3MkdmVqz07OreGeyfwoXf7n3NO8mzWG+G
70OXoPZBDHcv5X+JBdCg3231luFbUWWXiSHTStxgh+Ukn0dhUEYagBOOjv2b+fzd
wUqBeMLnY1JKGU6siZwYYbcP5+jJCknpovg88MrBNJ/DXarmuLb/IgqKxOmgg6gd
23dgrUMnqjzOkJV0VNjJZsgu3hYs0HXkNGJCsXR2SECq4WwdeCxg+1RDYz3E4naZ
txtILlhw4q1kJmtlyz8TPU8Um7nSmrCzEtljiC1OZtTmGAWWuL6zg3bvOtqKH7me
h23VdfqYCsQBD08ERB1WRytRW28e+5G+msh6r1KD28MMahW/3S0qQzk0JbfGG8I/
b5S2HOP/V3wjS6vjkgyRGNJqkeKT5M1g4CcxDuwsr35/coZi+fpbdOubTavX9BxM
pEsU1PXOevqDKMcRjYKZ++5o8xHdjwkuAHPMcfYbCTOmKn0BDMMzFcbEzkAD4fPQ
OWmlz+YNQc3imWh3JEk2aBhuPercdPpkzDoLHsnt1caLrR8fDEJEcYfcNFpapyq9
y5Gk/8PXH5Y5/7d1WMxhchNp0oS531dcyNSy3YGXY4u/yZkN91AE4shpR8vTibPG
aykFFze15YWYSMV8PXaydjHOg5sqDqmVp6SQVfJ57+1qN2xpnyntdqMnFj99C4at
SPYL7bKYs8BOoqIOTqz26Jrc5pyAH+duTGpDV3DVbarwrgIKisrdcl6mwtwgItTq
F+2bnAFyBMSj85OFmfHjP1Ov9MuPFP7rTV3FczqeY5vw4MYK/MNs9JAAb062hlV4
RdSeKprPcsFjC9sRUd+T2s8Q0bd+VZTmCs04sapvH91+cvk3TwckE2qjiWEVgLQt
`protect END_PROTECTED
