`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gwTQGPKb5e+BI4tplKdNp3ZxXv9snyo9GY6C1a/XwIZXD8fV5SWuuu0JE1yMOYBS
DTgDC7EOHgXOObd+ZXtVaXg03oj8JJdbY669Tc2Iq72eM1d4HV1qjMSNUzEgaRiL
CI/wKCoUNswvXs8xY4Ay6UxZ3wgzu9YDxPU7x+6X6Pl639YV9/P7WqUmDMJsuVZI
9BRLkQS8yxjvWYheJAyqlHfNplRChFVfteY+05Tp64s4UyNlm+WE3Ctoabo7KslG
/N1bIq3wosgrTL1WqJTzfEwBZNDJ40PGRyBRv1ZDYkaj7KAPmrX9YpsCVbHHkPEg
wUgXTdEuTSgIhqEf+3bA9R6W74Ut2h4xYiKVlFnDKr1HeZKX3zvi38+mdZX8IUb/
QQWi2Hqp8DvRTXwaN9ZSYajMbL9gX/4l4zURIVTJrBpMAbDTIqCKBJ8eRVWVeV28
9n6dFW4KezadWYQbAoRlpkHExXCNmC2YOMqXwOwD1YYzZsdw0zj8WMvdE6bjm89a
bISFzgS4HPVNjgYPGvygDpsuwb9HX/hR+IVzeXYQtnTRuReXnoe5d4/PoEgPX05M
uctRZpGsQDaw95bRIBppqsjqr2TaSH0kqTcU8I+d8g2PuU9+JEehaq0wN45T4yLm
k4pM/0L33+NRGywhUeMllELhrJ9guJIE1glbUGVNAcNdc6pkSXq8k7EEt/kejMDW
UhHJzpDJIok9blHBlpARxDhi2fGnsL0FCbGbs0yKfHvYhGAGuPJ8aXHOIYctNxU/
abbKKYuVAlq7yZ7bIk6a7XUuUGYe9F+EsA0X1Bf3xnELm0WQKtcvwle6YnNyaSzj
4vnrYw3SM7Y099QRIITn1eXKpEClPquDGNRRni/V2QxjBa3ZQdp/PYY3wCjBanF1
WFsTa6svKIS0NHCQlb9QJfGjiT0pHQqb03W0bMuBgtF9cZoN5TokkhRqVySUjfXZ
ACvNTJLGdDSmph74Mnrjgw==
`protect END_PROTECTED
