`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C3rW14v8aJB9KqiQFeoS5jfQP7ePEdwv/QncxFwJFKSeJH/ywI1hZDxrK1lDVT5R
H9mo/gIkDhcuK1bM+80cMU2dXv3SUYUzW/XZ0FpRwtn4JSSvEJCQvVSrVz7xC+Zf
6oSEpJabyXqv0erSOFMylO0fH5KuDeEo6de0TldqV7koRygcoL27Kjm1Hv1e2waz
AM6Pw7UjmuI66TcGTEkjgaZivbfE+yrPYcs+Wnl5Vkv+rYLWu2AkwOJytaqz0wTI
KE9ef49xShziZ8WwhRv8PJGFnXman9h0HNDSfKduHfC116Rbx92cCp7cnjBunEyX
WXG6xPa4eVsQ/FTdDQ4VthdZBH1SikPS2ff1KQOxnj152wImo5RFjBFgPIBr2r6G
aLzc3pye9T3VoRY/1h74ejrN2HNlyZPYeH+rXVIg0Etvm59TX0w9Q1/y8AwBmnZX
+N9aBhvdExU/RoUvfQoawrH03w0Ep44QaeJgpyfJ0XOl840jnQ+076uyxmag0BPO
bpu9wjn9daNaz7drQ8II3sFP+YRxqS9N40bnrm3Clh65ZAwhmDHNc6P28TgqFQIP
v8+JkKYAZqrf/K4ZhISWC0F+Z4JpXrtEBl1snkuoEfy9kJbZzj1kDH/OgczfDrgA
NECfyp+ogOWxgAuNSjgTetlQDAJQV4ZSSPB5Y38z0LrF5N8WBeAK11t6NkVnrOuo
uX64mh4TK1Bh1VurHKR57uUVoD+r2jyRz1jrGL0dLjEZN3l36znUM34apWMfwiea
2vwQGQRYw3geIjqcdjRxRBst0MBkJLnYwp2ViFvmle+2H9jvyiVRS7vexa+fWHBh
/isiAhezFW/twXJKAM4ODx+V9Shbz6lU82AytF2ze5SHvcxxDeD5f9iTq60SVDvu
MZ9Q56gqGk6L4kWY3mK23Sh6IZfUsTaH25HWogkK+g2wcFWBX+s/HQKLBLiCxmFC
x223CsFTLKNiRmZ1LwnQxVStFF3gi3Cj7zbOZObJrtHMUQMWMghWXr8/UdRPtcni
/QB0RE2PsDen5RKEga4xVQ==
`protect END_PROTECTED
