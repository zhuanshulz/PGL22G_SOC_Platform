`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VPpQOgVdEqEq02Aaq5iSeR3xC4esd7b5SYUiQprUgYy+oi/81S0kw/L9Wsyy2QYT
dhtYbTSHY/4PAdIHF+3/l7SgmpbP8Pn6oVjMSGU6mHudeHVdt38UPTmBcQW61NAA
8R0TnGrKyLT5sM9ZExzQTNaJUv2S654Lxbx2kap0I/N6N9g+9RDZANwv0CeDhyBl
YQYMrCSnKuO5ekxUJacbuw78yID87+QICN9E+piQGuW16MP9RFp9Es/L4LSX0+wS
nRg/U66ofjTdgPctZB+6fPknlfZW6iPYlb5gijKiFHZT8P4G7UTNiAHdn6mbRh3b
rkYGuy5ecRfsQ1XMmH9xIdci+N+w6S10lai7le5o2rqatULEtpsFX+kH4XO8iDzO
a9qm+CSSAxc2FCugl90PMi0LwpcE5nmTBZjeKj52uTBBudTQGKzxj2BG9UWgo0Ps
CGx/x0unNBNNtFwS0H7IwbU3XvmisPWydsMaS8Ehahgxd5d514byjmEif5PZWOlI
1bjy4VnJmlW5Nqyg5OKaFojoFQnZfin32cXLsEIfRbhiyPzjCrQMpCUeZE3XWhl9
6BLi+X8z/KtYHCUiCKbLTKfjidp+mIh684DwN6rEM8+oB6PRHXbuC+g1VgsdiO6U
Y8ezzMIWxiYTayxlW9yUKQmXa5DLr8jgoC1x0z05h9Np2TVBaaRmjlr2d/Ysp5SZ
d11TwE/OqAzp0Vatx4Va3xNmrywzWcpcv/IcbPj4C8di7fbSavFh3FblVM6af4+X
0eovugUIgROd2PcsXbT3QFTzte0C9Dzx8UyRzMC9ASiTMumfepxOXe563dheORGj
oJdyojXnl68tzJVZz/HZ3ksY0flFUXusciycDa72JN21xKBv900hByCzkqEzSy1m
xeC/DJ32EFZnRnPLnum2QCvBg2yZuoD7CXWFeFuKnYptYz1aidon+0RXp/zCArhp
ZryNQqUEbRAmaX+hcwTbAUGCLyrWYOI0/wK3A0kSlNuZkPWMWfdtHB5goUcsl+nz
5tvVBLV4KLaly+nmbF4cgQQM/Mc7BrTsG6jiXGw9hyEsJFwMlLYA/JokQywK6gA7
nPhWkK7P69UCxsDhv0tgADnxMu0sop4FgybbQIKMZnXW7q6C4z9EHJ0RytfRffJQ
PKg9D8JwSMOv/Mviybl3YR4TFbzdCIqYKruc6FStEUMDx+NU/w3i3AFur6Vre1um
VbKIGPSjGbx7h2K40EG4qRvfaf0DiWivbPtY/700rh0ppr0NRpHqgLdplAa5e1Pp
1JMkDidblWgBm5dfp28xXwJvdvWxrxTsbZsk5KcdGZZFin2XbgIyC+/Ww/8Kr8bN
5XDykV1X+lzrx68dMG3oU4TXwXEl8rH9P09DIPkZOuSc3YFOuY6CMFiD42d4GHFj
ogSxB2jMc6G80j43z71reNghkkaPuLwtJb2prCVznOpEWrRZHVQ6osTrrU+xyH1/
U7S65pfnsA73hReJ/IJmIDq7AxSV6zk0ZB9VKEjV5TZxGlP0MM/A8A8odNljZq8Q
Eib6teq6M//FEA8PJWPb7bB1vXYh/XpGaEqb91sEnKl1aKWiiACKJDkPsUVefYwD
8uIndpPKXLbLU0k8EMbCR/gVTK7ug2Z3lFZqxcqyOAT338ZKRLafQf2FM2TX2WxK
p/pu77mnsJxvNdCn2uXxcwYxB/ku5CxLse4jrp+DS/fiYaHtlEOvs/hvHper7chb
UgxOFpOudG0a5mNnu6wRIIBpJDwGl5ylXvvOiwx2r0gdLklI/hdAoiSR/Qgrv1y8
1zEiK6B1GpgZWy/sMu78VcBEc7Ps/GDdMeilXDQo9f+mWJ544aRRE+NhTt3QpplC
DkB/gXmufscduX0uaTZqBCyXXqxGJCrDZFULVEyVwO6yQK8EE+Ie4WUPyERJI4A1
RfgRQ6089y5WItmzkI7+MYjqpzET89TkqP4hJZ4M20HWMUS6mCBNXVQ11VDznFrQ
Y4Li5mESY9NmEMhqLUxaXQ8XsWNh4/l3VUjycNmrBp7wYkm11mdUC78mS4tofTah
AFHtQIiRQyYTU1wNAq2OBeaNuNhsA9ee6CC3bUSw3AB4HETi6OP1fzOPV5QYN2eh
gCBPA+pU8RCK1xx+bvJfRC+wKScd+afJ/Y9KKDVDokm9EeFf9SF0UVE+wgqK0dcg
cSAQ/CzYjNVXICGAISvd7td9cTcth5OI3aaqcJFgIN3IyMAesxjrw2PllQ+hKTBe
Ul3kcKE24fDfR/nWLp/ZcQIsXImDlHL1+Hjg/GoMt+m2RkC5qhdsjkeYWaCyM0qu
YG1ZisrX5gfG6FI2EZCOhKBXiI9Y78dGJTiC/TkY2eh2th0DHagDDQ6ux6hBkThN
3GyJPYqgGfmvpu8Neo3mBwHrch0yAOUBnunFfENPKNPKm75NwVkjIXEJBQ9uWm+I
suiQ0984xFTnczczNmKP5YgFj/wUoE3kCWoxC0sJSZv/ozCI5uR62oko6S1ZD+sv
tekm26BRyOCL9x9VAokExQSijT1Eejtt20r+Tfxcu60+mZBZdyvksv8V4QmhCWC7
GbzJ+42wQjSwe+0OU1Dk+QxSFyFxrhvq8bVznm31kJk7YoWwVdl6qMr0v7/GwaMW
Xw2+0rGZniPMNbUi2Fi+DnElz9UsF5IRPmLtRce4xRkfUocsHzdJGh/uztYNIj2g
8Ro8SywNRKb4EoRo3ugUyiAxRcyoxjgcB7+kyLiiENiRUMql+J6J1hH16NMfAC8N
LnhHbzIkIm/tU3y1Q5A/4+4TInFu9MkIxeAOG7CfX9fQUzf6YI24oJAWHEEYBhxn
Dch44Z0G0h2JRos8vdifkg==
`protect END_PROTECTED
