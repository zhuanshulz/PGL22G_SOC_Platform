`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y4sGdXzoALfkH8XnZb0jvhMSohR5ctKaVcpRmWi8qZuByQ7+YytuOEwxKSTteclb
uc/TmK3PebCE2WSowgSfnyBSGebyIkE0VKkDmL5+KCXyPS7745tvrhqm6j4muYJB
mmj+9MA7t2A5FJH8VyDu3q6FIqX6eho7k1K0isTnefnQcvTbUOsit9WulvI+Z2q4
2brQg3t8fPQ/Q5f4lyOGdhjG+M69DPXyK6eaM/GqSRnvcC0F1PheJz5Hdd6kbtlR
weisHN5whDiTH+fDxKhT5JlXP/fdR2D2XEuZl4wa9Sv07GIIpWSIuLD+b2eatNN8
MrXSbOmnBgJ8HRiV8mLfmfRedaJsTFEThyAfO0h1fVQ3OYLvtZZe9bVT2g73s2//
0bf4zvf4LBtEK3F4vvJj4l5GeVfV9jLbqncT4+v+HoDoGt4QWB9qItr90BqvFkbc
JUJJtwyD0DP3a3AvDRNsdk0wDn8OubjUGbed/F5pQMzIJE4dnOtlAB9DqZgBI4XG
k31KT+7DnsN7kB3WHpy0RTEgfAx4yLeivu3fZBKgAZl0fpK5OpyunTJF8JlJPTIk
sYTwz7ULUZjCrHjF4cWGKvAQwYZ9jtsioe3ZrmjorX7RzlrbHlF/j2r7Py4tCqUJ
dZRu50M07mUdsqnZgIZgJyP/cFTRoGbe8dCZ31CawWnIW02Y2gPnfhhNW99FMmvR
yAQ3/RvtJAbBNTfdtEqlwGhbG/OEsM9zAiL5PfaFEsRpXeROelDn901f4Dr17E8S
mC0Kxb0uOFZPpan43HdTp+jBokwwyPS6iLaA0bpyJEKrC+z2onnWGhE3nds4Di7i
Pm10UVCoCfy3NA/vTCs7tNJtGmyAzm/VqbyCvz0mII8=
`protect END_PROTECTED
