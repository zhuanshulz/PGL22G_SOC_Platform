`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e5sKu+gS+js+VpAW/CE8Ro9GVtjZRhxej+nbW2LjguacLieQ7eCuG/YheK/AlNIS
rId/N65q7cyup2tqi8MfxemugdVy3wTl6TgsOWV4wgC1t6Ua8CwmvTIVvNB4WJ4Z
jSERNJ3iXUUdUc3yjTVNAMg3YHGz9cE7LNmIh2pZ0VsDYO/p+jX6lKboBtadk9Pn
larCvKFiuMi13FgKjDgatcdqE96HakDG2FxhmMn3VjsP28zwYHiK6EqVyqi7OtDY
ro45RK3PZVBLk2zXnCi18ZCPpm5dC5pW+GVqd3z/iHJe2vu4U0ARHMZjMVP0wmBR
cPHFt3S9aQNAtJ0r+DYIsrFZa2uIPLiyJkkfrw90jLOORbg1Q5ml6UKTlbzuu/35
xKN65tbmwQP/iBXJA1ov95uHj+MSVvev1nvfwMQPdXgwdTY1XLYdw9loyg52hWcy
dOf5gLV2w653U1llrPcK7+dCBvhw2p5HvPMxTI46EI7bsU7li+JaYiufa/LS4N7+
yHZWpg6Rys0Pw0/KnwrsF7n91bMBVHl3geFCsHAQUgprhDoPzqdoUwL/dBSShERo
MssRrmz0cBIxUMLiJhrelyfxLlTWFWSi3YbWp8UYg7P2AqTuTqsj/pW2dnD2YmcJ
atsoVOaAvqhoOTOFDMkl6TGML/XT79sDB0aQw5HHhfbtu1KAK8fdAy3hU5J0YgWa
tj1Bos2j5+bpDSAYx7f49MvComEYZZXQ8xfR3E9Q3u5zQ5cJlPC2E9JGzdr3/IWk
DVv7i+Ob9hYQUERdEf4/kxzdvM7yi87V5JrqZgleDeqSc6sT+6vNPc+C6asxdN+n
oej/1dkeffzUoUrBIWIWI50Eip9H3Sh+aOpQrqaWtjpiF9eqnmf3a6hkw+dCf4bd
y4RddoH6EBbf2lF9cnMgUw==
`protect END_PROTECTED
