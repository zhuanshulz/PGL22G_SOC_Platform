`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
absAIzaokctCXZU4swWtnHnOfZMK2rmJVUhIWwyGLOgfxqTT8iCWZFnUKzoCk4hC
J6JE5CZJqvMuhPpbTZVXH6n90xUIWlwDynkG0cvqaB+HbRHoBetjJIFJ0E8wTDkP
2mMk2T4gKzt/o07RD6fXwHHXlg2FBSMY+pmBJ4jp4bTBVkToZaLBocIy4/vKIriv
gnbD50p9/QwvHKMjrpwSr8k5MtPw7dxEVohO7Ckv/CMPTE0vEtdkDkMcbDnZay8J
O6RLp1e4Ca5hmtP5byV9ZKQL4qkfiEXCRoV0xq1W2TR9W0alfmrznwsqLNreoY1N
YslzwHdKCyeYWt1iSRpq9e7ZzXiEnRlR+FRmnBbiOre5FGnhErOYSZVKAoGTqn0/
C1FuuoF/+KvzJWZOYWYjm99H9ek5cNShQM7Jt336i/DAQyKnas7kkKtmRCpSb6Zq
M4QfO3KPfpPKJqVy1ZfyiMDBWAXGOOnIkjonKijvSc6eNnnlhDmSnZbJHJVGpOnl
SHXWbhhzU4obKGp0yhMONaz4Ayb3Sfg+8AoAPt1Rc0sTzZLmnSCPbMbSZoP+aNK1
7I96ydVKaJ/pV+X/RYdpUk5CL9pKaaAXUmgPPxmU/Oi0iwSBYd0f+CQOrcrtHZTV
xL2xO2901/GGY8sgSPyA0gyfWvlGftvCLPg+mD/kWAcLLiVLc0o3aWb9IAffOrDi
Yd3NHIAhXIB42dL+mNRZy69RxYcKr3aUkSiazyBpzvI=
`protect END_PROTECTED
