`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xjsqa4TiTDF+PFepxi5/mIsSUMoGn0YOPvK0LbcnSGLhjEoBtTdD99651aCFgCbr
2bgxc0a4Sn+HHQIRGsCYE0UX/ezVKMGnry7Xu6jDp7YFhaSqw/momKisVBn/8Mwc
nVDZWQd6oqSDabsQeXsDoscvmoB8zdmmhXBfU1kpCfW+X3wQmWFsBqYbsPoF9TQn
fshIQzzQp6xMUz6HC6HsfCEY/QNHMZ4lX7Kqqvg1SulI0UT5a0bLCyDCDtyVWLDU
im4SVYY2VqmGvKKp+N0fNZ4rQFUisOgB6Wt3gGH6mubCpZKyBDijwN1dpSYYawWv
xSACEylb59Q3geixqy9Bj9V/bEdzNtY3zs4GWxVDlEl/XqVnEvRno02YDrN3rD3C
UbnYp/16PbaLQdx5iGaZDbEhHBhJJvCYArML8B3R9t16o5Ax8wOfsF//S3wH9dLZ
+h8DnzJjTAAUCRbLBd9slV+ag/TTPGcte2uXG3HVm2GiHw+Pws9Xw4SSp4UvRuPi
5ZRGhzNJ4ht52/xx1feqFbw29FczTfeFGtBXjXxNCM5KxlY5ekw8epBeGeViqitK
Ag8SLn7HkpgJhPNbIHAgqxwUYUFO6lGrgz+XjCrn4mi6xwRlHvKH03ceKOzn5bT9
Nx/ooFQw/J+Bfnj9PDGQ4pfSJUFbEI47X8GPbZtb9XEIdjII6/1vak/c+kAmmZtY
AGNrX9/sxB3WTc8VU+gJXMravrAB/l9rOi6/2RBs4a4c6qWVeNKKhcj3XemxxUln
QOxxXFozK5IL0NzIruqnNKpxzXGCxcQ055QVdzqcpUtIKY2sDilLBCxHlOb0/MgQ
DO0mR0ktYRMiG2FeM+iv1xVXyzGVTFpzd+JWvvNGXfJCScD0lfjyZmoXEfRj6RlZ
2nIrpJbRGb4RFR4mJbkgKOixKC5RVGN1UQGZPcI1PlMrYvbg7no7JMMpJU4aBS42
ELTYl3N+o3YLl6vO++1oILPqyblP4bejjbghNOHiy7qbaFuWHQHxnDZnhrG4YJUe
AoDCNkmKyZ5JhcA/2UfX19G4Nm/6Z+jJOy+ZAM2V7W1W2hzndGsN4sS8C2EhfgaM
eU4Q5MZcyW6S5TUj6utJijEGr8BifycsmiuxtLH3SGBtPElD2RFk3J69O5RkdbBT
mioQa8oTvVzu4vAkhbtUIOCdQhkOhjY6F7HWpvMjgMZZl/zTi6nLSruXB7gi9D3n
bAl3C1B1z8znsCzy1Q84cY7apOy3mEX0tyZuErHz848QCPgAkjbZGea3EL9CNxm7
JsbGoPSk88k3eejp71Gnig0Zk3jwXaAfvVIEQxZtOIzBz0R+L+DQ1nJxC7Dm82MS
MWEVbNBVpQKGtoaBpNoKQe/wMNXxh7HyXMTSUVjQ6Ni/CbzXR1PtAF9BOqXBF8Zt
bvuinfVsh3zFW2sd3piDwswdyP1m8TuVRYHKVyoP7HH8n3IrzhEVD6VTh72Msoer
mPoBv9ryEmaCIIeRtpWHE/L0FCGIECROYLQNd8toQSn4BQ/XbKCpO5HCtugNbTlt
8ae52yGFGU346LA9/4tiSJCr8HvyGn0b+D8mZJMfnMeZIMPAsskD74AgnhaUmcgF
VBrFfDq5LH6NdPSydRd4PDAV8TpxOPuA45FiSMaKwH4=
`protect END_PROTECTED
