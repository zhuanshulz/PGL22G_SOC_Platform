`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FcbTl8asIGXnJKT2cKViGumUI9zjWzgU0fsDWR9jtsp8UkgGzYmhnxDZM1WwdxBe
BUt/Q0WiV85IJO7hLFVTEV+ajOyuFQ4qoalr/kb6pMB+UQRLyaLSM5Y2fk1S/nGV
/PfU1WH5RyA0q3VC03uTXGmhPsDmZ7zpqkE6PDn+QfEKVby26ktT+bmk/06MNzLS
QYa3w7V5xaKIe4lqmSj74S/oiUXg9tjJVlauVvsA0cSejorXJhtK39z8Oj3p2jaf
SrL0t3ktkP02KJo8hfF94g9KRhh5OacJrmqJuogBnw7mHO6vJ6eXUNJqqNgTPOSV
bSQ01rt9gnFu9gC2A+V3WSXK84egpMtdF+cvSRoH1aY8X/Y5qt3C0rKW2UusBAVX
TNaYAIw7UBHFhSaR0HjMLU07PpzpKNxRefqcp70NMZehy/rLvlOWgzfKtoDWiYpA
o2tFX/FqeLJP3pjI9VGbqkfCpOjqjUYDCylEVX71JGnzj1EvsCdP3NPaTZu6OS9I
ZZCuWXb4AjyFnhJeO0LIbXIz1PBsHolQYEi4AvnJHMPqTTsLSv9wVtovkuGDuMQr
jnKkJlulnvaUdAWkZntg1LVADj2GVmqNdqdOBIuyuBPLwowPf+lkAv1H8iAjCC41
oXAzDLzis2xHZ8mIQn0osjCrMV8/IHfEXYkvGC4v4Ba3ZemWaPZEOCh/f320HyoP
tlHKG1zXTC44nTSBEoiu1uHycJfnDt6AtOd6u10T7grErIgcJo4yoJmLXWm4/HXw
BJRfskXhyct89wjk/2KgZbIV6SjUkBqpGVHu9y1Mv4kulDonSyo3nDBV+EcfhAyd
6IFK4uibpyiyYgMxq9zrFkXsQbC0Uirh/7P5qJ2czQ56SCH37wT3f3oRCcV//4O4
EOnCqMh8mqFd6r9qemuJufElXUuylvpecyDmzTQ2cBikujnnVrOF6Xv8ZyF+3A9X
AFGvv8dCV/S0m99pN9E8YoJUrox5yVMP6+8z6CzqMlmJJUdxsFW+uAA5ciSseDZQ
RiQuqxb3QEnVwaBzYX+6aNyKvkdwpWi/eFECgF/JK8vXrq7k5wp7hlx8xZTe3cs3
/DR1kr5Bh0aWr+bnZ3RZ2B/EBJNGXhyJxGPruqGbYf0dMb86wAi05aXY5svx/UcQ
iRlw9eCU2bAIgSSsRym+5fuFFm/7cjbeUo7dkRNWYQ7ca/i0u47i+qaQjccgsMQn
NL0+SEYSYkR68VnJFrua0umhFiplbayPTWEgjTJP+0RHr8u121bsJdUMyP3bk/e9
Z+76kJ5ZfutsZ4OExXNwQ6gH6YZyQbKJXef1lDI9l2ieiF8SBaulMObisTfJ5yGA
eIgm+Ix1/6X+9h8UjN95tfzEhyS37zAmqXI/+HEyCYe83FtOB6hgcNd1bWjAm3gR
R9W9vWSiftmBim4YUWhnsRvTgxlCeVcaHJwYlw0ADb7UueY0ELGveEMAY0wVvA0T
Y4MVovb/LUcjZMYc569JXOUb/sLZcNp51lKtF3qiYs6X3pEUIEYSUtm+eMuuwwau
DedYBNKwMrQUv4+ocObDGjRdU6pIxsO1f9w1FEQGJYkYbdI5saUzwY8s66gOOVtW
HOGcGOnUVV0PAnvWIgkQyBcGl/5I89jSLNn2EyCVZEOnVCqRbb5QJnHbqSZ4apEj
EvzzNLCiMsWYFjNEhnBOpryPLRy1HdzzOTmT3ODHzG5AsfrdmjbiBs7aANmp82vn
iN/7qgcKmNsvW37/EgeWgwc2xpPAOWQ0YQlN0GihXKM3BcDBluUIM+LWIe2w2oWK
hZ714e7NXU3YSSajCnYEzW2ZglojKZ1YgH5B9AzOeGY=
`protect END_PROTECTED
