`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M5nQV5aq3kJSJ6NNgI1uvCEs41YhVhWE4Dy1jDtN3g/kG5hiISj+NNEqAy/QV8Fx
JsWhhtt4rRpOufoTPgDSU+k3dX+PkKBlNGIZ2B2kCLpvxRV8p7yiiV0OWJwbF2ft
hu3rn1T+FNEz2JShOIK89qVZFpmPbmHFNxMmIFrC6rWDGr0Grp0JbZ2m7r9JOMN8
dt2NJxXhcSNZOMacC/6t2Znqlg0+aqLA5t7ox+wVfYvLG/xKYAjkmzL90fcg0rD+
iNI4+5tadWxv5NPys8MA3lmoO4vRQbXljoOoBVHRbSmyWCc60Q4Kk0P83ZYdgosv
KrIED+yN/TNo6XkJNVVtATeNTHVKXaQsL0/Hp7CpPmvPJBfWPSRX8gnLGVQxPnQ4
zMRUzppWO4UIvLEJINLWXrfbH34wyqQpyGzy2YkOaVK0s2EI97uSQUgrLCjKRhLC
GONQDAU5hv8Ew/UEHnwbt7EfBo711E/8kkkXOQx32ZV5J7Dzlt/MU9kty9Lf12Mg
lXs3f5dbsM/Qsi8i1bwgXq0JcHIy9oY/OkojtJZeWkgM6YDkZYqnOQkQoE/fhSVG
`protect END_PROTECTED
