`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pXxKmx3zv243EaTeUuSG1a/eTbDdWuAb99pGRBee+SsjZv2006XPWFJhMPMjS2MZ
6OV7StrQmLOUwNE59aTFZlTTTjWfHHASUZWohmOSniv6AFDkp1/UL2Kb/7A9w5jK
tfDduUpuuDRlbJXzEnfOeBH0153YJwnFzT2+KcuaQj99rftEdNYY6lljLte1ENMJ
HCmpdjlIRHI3/DyzLKmhsTEMrL+5RK6Q9sjrst+OLkW6r9KU9dPbt7O9Cq2eK5P4
wCdCygtOic78yPy50sm7EwPeJ0yZuc24/ajV3JgzQxTlH0JK5CgIJX4RbO9rrauI
Kl5QT61OEQhdIqQzoIKT3lDGxv2Wc5ylEg+NIKA66EIHqPWOOfkfyzSa/RnRKNBT
WPmC18nk9lP1XfLgC+SuM7nliU7LTNXXxbeXwW/KNHv4K9r7kz/TWABaxdxVv8CP
lEsM0z9VwYXz4curewcFAwoxnqVtt6biZU+oWQyPGpLth+rhu7PV28qFyCEu4vi8
v+wpHEQAjLQH7RUJOj2FXMABIgtcC+bVu1+JDNcX1DE/Bww1JfUuNBCO+GqtF58F
mWxeg5Zg1BXq7UYx5OBD1O+6/4q6ObhfdfJtS8q/GrXjg3H52xQj00Gj3OBgN/gC
nBn3FEYEj2vctWp7TC+kGZX6CQSmflDRRNZGENLOfDvGUgW3rIpd9ie3msKMmY2b
TtZXH5YpwKtgh93xN7yOA/twCa7FweLNfTEpSNo7YXbTXC8wpq0Gv5JQ5dKucuxD
5IWnT85cLJCkKKWeD+lOM/NAXJGtfbZbyS23S0HvKcV3sVsA2x5mCoN72JOljQzU
CUcHa3A339BcdMj5BijjzN0+ap99T3qNIqR+843G9szKKUxsi1mdLHF610vZv/U3
EIMOVDF07IeX765v1EJLE4yGfjvD43eFhSDKxwZO52Ucj4CroYJe14gdX9BjVjbW
edxWfLBgQXNpu/FDaAMYP6GCDk4qnI9KQWEnRQySBA6nAzAkyFbQMLnkERS3aW9C
mxIwisJ3tAQrdEbAQJnosg==
`protect END_PROTECTED
