library verilog;
use verilog.vl_types.all;
entity V_OSC_E4 is
    port(
        CLKOUT          : out    vl_logic;
        EN_N            : in     vl_logic
    );
end V_OSC_E4;
