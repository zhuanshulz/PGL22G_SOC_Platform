`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p08wEHlkmNzbFVLD6yQvzw6Pl+ITVw2lsOnbenPW6BENDkwrcFfq0L3J/W0HvYHi
7V9s/993R7loSEUTcrjUJdalJpyzc/sudfOZU6hNgp4+UXt68KAvd/Y2zsBFfmnb
FdYl+9BSoPpPcYwHiWfG0F0v/w/V+wBE7DFD4Y4cwo2kBAGxXjp8Plhtc4v+avth
/OJEr9E+IqAdtdr3webNOxeCb0wEaHTaR5uzGmclOrTzBILWczE31tTGm4nxhAIG
SRJymkw66L7iaYj8gPzVOCLGByN+QUfFljANXBTodghM2xkhEuu2iFhIpWnu2T+Z
vJQ7pNQqG0yZXpD51YFycqUzwqJOtuuKuwBK6E7dYwsUb5RUWfyO+5Nv2HkWjEOW
Gxe51k8UrG9l7JN6Wp5oPd/rbnJ4t60nVSnKS0/qhVhE+3RwhawKkvgJr++judCU
Ywbkhodk2aw5zR0fyBxp7QMunxFqbgwOspXK+1HKIBrJT0yhqOD/Ygz3peBwh9Dk
0Shb49m6vaS+vxUgXeRO3YdJ0dU25WtZ0P8dE5e0tIIpDWOpfLA5hmKpVIKvjHDQ
zWiL8m3wDiAxg5mYe4kOwHCBSoHy4TBEd58BULxDBJew3zl36SXd3zo2zY9JlB3b
yoeXDRJzMFjIGG0GmN8/8px5noacLSzN8v9cdRaKbPDqS1m3BOfkU6G8K5IOQz6a
sBPXnfE6zazby7LE2y4L0gZCmO3Jwse3qw0WMcZWv5O9CuSziIl7LJNQ/P+d0Igz
XM1q+ZmqDMUiNygzKXW4Am4/9gZnJ7VnhuM6SLrL1Jw=
`protect END_PROTECTED
