`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mpQBH4x/kJ5FItafpiYbFRnF/uYb1dlXR7tYSgxBAG0QL+tbr8MhwuB7FYgw1gXt
/akEycWQskooOCRfb5sU3Bv+l97P5wXZ/dA2ScN3BA3sXnJ/sbZd6PbLQDwya0j0
TIzuhUTBdnNEkplEsV7/mDhT3Ymmb8mmUz0pceC+DBeDDUXIwElEjNwn/3HPKJO4
7uWf9UBGHCgbZvlsjsvBPvo9J8rY4gCZnSQeqR9Wisc8UZUQUyYc5/HUBHoeRnTZ
QIZvxQObmLECKsW17JjQs3TMS0ZCgtPbcRT1dthTWLhlyDv/wvZ75Olgl+VdGYdM
iaFI+WKb7Gdv4V1ktDkpLNIrSUlgiee8rG7ZFH9/+JlX9TaU9occK4xBhrzcFpNb
w+/6dySo21DsojxmKE1apzynjR/pV2lMTcPWdSM6m3tpFqiazlYNSnFnHD5lMS3T
mKJO0TH57ToziLeki/ijxxv4POOicRkTFa4gKc5TSNLPEYSp8W8HOvqG2/ukoW0f
w45AXeC9p2670s97Zh9ga4G+Wxp0pMG9XPR62cwpjIA6FXiUuorc5dAstt0A5Qt5
N3PNtVFLHUEeRSE1cFlH0rG6CJ9gLaLTAHj+yhLU0sNpJcqvUVG0YdQO/FGr32Tx
mxv4WUM1lGoEE4ClnwskU+oPijCeWPe/6Hd0LGLGjASx1mqGHQW5l3i30F0vsESU
hQ8cHhdbYy7vIIyX4m0LaKdPCcbR/Geo3auXCboraHD96QB5K0wSYXpnbtjvXkLk
yxv9UX9sDXzQrk9PNfv2QRACPHT4/kxviCoJselDw5x4zEdcR+mwbO+L32cVVfAB
Y62+yNjpGzFxUrnHMJtyng==
`protect END_PROTECTED
