`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RPPKP6Hf5kzg/r+FXRkqRi8FmdCrL7mW+1OJjWOsCxpVEqmbX6QG3GgW6yr6jROy
YMcRcQ5QyUpZiFXORvHr9TjRAuQ/bdSJPE1uhm4qqeINkYliWUvKxmmbAhbQN9D/
kmV42ebRu0oz49xfKrb1WYSTt9/SN0W5op+EXWTd5wxmwq84ajiHZ4XOfiRlgWxj
MU+IxjANfYXt9JRVhFF9wZHd9Z8K/jU/v/SF6U1j2KzvEFQwBoWypVpBZB53s5sP
jrw3sf98yB6RHCFitlKryOhpK4fvgTUEQD/H5NKeEthvZqN2J3Xzr6pBX93Kj2l/
+t7iBCt11YTCuQVh8U4xqfTxsFnGnVdJspVM61ib2wqdGSDfQpXbIIfv1wyl502X
EqJUd23p8ZLhjhkAG3K7OX3LMpanLlvOa2ESoGey1e0G580OTrYabaoZPvQ89iyp
Ie96h7Dj2WgpHU8I8qJ+Qtjf03S/8sDCbbwm2e0lA+t3zHcUhunf2pTKHgQz/hFb
D9whzDoFr87c6xoiAKvhAikR2QiLDBnjoHf7/j7Z6xtmJPZyN0pjCJgaAhSQe2da
WPyu/kQ3hocT6VA0VEadb/Bp4wxoTrUR90aK4rajM+kZmzRJxrfhwb8giBgHbXvP
cHHnWaN9z59yck4E9hhtngqiQ8qt85pTqaElmTdIp1yzgURP8enl5CrOJWa8P0fB
onfhZpFCEd7XFuQxDfqHIuskhIJwv0yOVZlWTme+g10uyED6O1uHezVwGkzXlC3n
pr9c9nKbd24DNMIWYtAxErs10at35qb6tL+s734nvMl+nW0SwSaIL6WcepbleZuP
yqGivYaa54iD60f4moGaSb+VhfNgkRE+tdqKWdqQRVCI3PdmMa24tOYcelICXWE6
eEkGEfgR3kKBTttZUEsL8zj83jFX/YygHhFuQrrvA0HFJcUyNjPvWZvey/7yX1Vs
hCa1G38lmRqKik5Q8FWgU2Rgn/C+u01hSdb4zZ3lfumZ6gGDCuDQBb0lhItgqW31
Rc+pUtrv2SQLE20UdBX5hOp/+bV1i9D5aWH73/kxL7QWobjBBJOe9TLJHl/d7tgl
Lc4QxV5Cw38MKvVXNZ5ysVfD7BpnFvb5a5WBC2t33Tr6JylVLf3XAC2lOcoMESKw
fHjd8+GiS0zX6MlDh8HbfV9TdAyBY9ifx1OWyamfw8bUWKOcHWTpOPjVW9lq6bst
f15Ft2mVsxBXO2JKAU26k8FI74bV9uIADJxc6hsJT6UjnAuv+sBmS3TI9zMrxrux
owtlIxxxnpGlF9EABquYYR3LtL59Zw5AALcbMtU6N7UxgkwdemcpfcpOIqXpNliG
aR7LZSm+nQreRC2C9vYMTTNDyQzmAltfjX8RDHnrzejnHaCJ88QXYMak+tO58MNa
CYaCcFdWVZ8vXJ6AGFHeVf1QF74TZCwAdsRac5IQGwhfAoCai+tBvXTjrx89myiK
EkRDGUjkB6Wu4jj6/Eq/UBBkwv6/Tf8otlXYvVvoLxQknbJjHjhtZSTPhVB0DEW4
ZL6zJbmlLDeMEjC690jusB8y5whDuiat33eNQfzOiW3eVfipLe7UTixs5ijfZ3xo
1c+6nrPa4tLVz6H5HNB1OjiACKlHXbFVDyjwWHVz5c7w6sqWUG0q8lAynVvtMirI
FC8XEnodTKtHmi6fuufv6N1LHM07sOmeWx4kDUVF3q6IvMYkSq6Lj+ee9xyz/0CM
Ee/XWoEU5xKNEYneV8+uLSbUok6UsaqZq5oxuQowD9MGv/wO0fQ7uWJVgo0LOYhS
WpG3TygdB+2Dqqrl9gZi+5Gyqp0xZP/mf6vP1okJDYPJnzx0KV/bVcmSjsvuiLn1
A0rFqubaVY2jQ3JBCiiJ6UuSbRaM95yH77lfYxsRtRpGC5xU48FB/SZiE/6kpFLh
HMojxxb29g5M2trqCTIAFYeofq+h2kGAl4hO/2eLWqXKtio6ZSgDqOKw/bi2FY06
nKfgbvj6Q+RPJArRsEMs45gA8DGHe+jfFT4YyyXf5Sq+U7cQ31vq8Def/O2nR9H5
Olcb2u7XWARARndlr/5blLApD5Im7pgh2wlhsXsxzQJkLr5lIFPLu7uGN395B2Eg
wzz7KaGDm9eW/lJZh1R/sEzJR8zHnfWmtzJYTWUiR3PZ4+oSMtoUdOHjVZJ7zDGj
rFMOXP1/hkYF0nI72oFgea+jtmDs2K0Ud+9N+/e4m6qkn6/uV5osX/NeEEF5S8DM
jzqs+ngVDNU3GpMjihNbo/9FWyCsSMl05Tg3unoIQEAPSntu4r5PwHz/nZ7hY8gj
agpK2HUMelVIkuo89Dq9tc0xPibktUQbDZivCNsG9DRWUcbe1Yu7x7Hq3siyQmNM
`protect END_PROTECTED
