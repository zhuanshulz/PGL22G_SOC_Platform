library verilog;
use verilog.vl_types.all;
entity V_APM_MULT9 is
    generic(
        GRS_EN          : string  := "TRUE";
        SYNC_RST        : string  := "FALSE";
        INREG_EN        : string  := "FALSE";
        PREREG_EN       : string  := "FALSE";
        MULTREG_EN      : string  := "FALSE";
        POSTREG_EN      : string  := "FALSE";
        USED_PREADD     : string  := "FALSE";
        USED_POSTADD    : string  := "FALSE";
        USED_ACC        : string  := "FALSE";
        POSTADD_INPUT_ORDER: string  := "CPI_MULT";
        DYN_INIT_EN     : string  := "FALSE";
        SINIT_VALUE     : integer := 0;
        OVERFLOW_MASK   : integer := 0;
        PATTERN         : integer := 0;
        MASKPAT         : integer := 0
    );
    port(
        CLK             : in     vl_logic;
        CE              : in     vl_logic;
        RST             : in     vl_logic;
        A_SIGNED        : in     vl_logic;
        B_SIGNED        : in     vl_logic;
        C_SIGNED        : in     vl_logic;
        A               : in     vl_logic_vector(8 downto 0);
        B               : in     vl_logic_vector(8 downto 0);
        C               : in     vl_logic_vector(7 downto 0);
        P               : out    vl_logic_vector(31 downto 0);
        PRE_ADDSUB      : in     vl_logic;
        POST_ADDSUB     : in     vl_logic;
        CPI_SIGNED      : in     vl_logic;
        CPO_SIGNED      : out    vl_logic;
        CPI             : in     vl_logic_vector(31 downto 0);
        CPO             : out    vl_logic_vector(31 downto 0);
        RELOAD          : in     vl_logic;
        ACC_ADDSUB      : in     vl_logic;
        DINIT_VALUE     : in     vl_logic_vector(31 downto 0);
        OVER            : out    vl_logic;
        UNDER           : out    vl_logic;
        EQZ             : out    vl_logic;
        EQZM            : out    vl_logic;
        EQOM            : out    vl_logic;
        EQPAT           : out    vl_logic;
        EQPATN          : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of GRS_EN : constant is 1;
    attribute mti_svvh_generic_type of SYNC_RST : constant is 1;
    attribute mti_svvh_generic_type of INREG_EN : constant is 1;
    attribute mti_svvh_generic_type of PREREG_EN : constant is 1;
    attribute mti_svvh_generic_type of MULTREG_EN : constant is 1;
    attribute mti_svvh_generic_type of POSTREG_EN : constant is 1;
    attribute mti_svvh_generic_type of USED_PREADD : constant is 1;
    attribute mti_svvh_generic_type of USED_POSTADD : constant is 1;
    attribute mti_svvh_generic_type of USED_ACC : constant is 1;
    attribute mti_svvh_generic_type of POSTADD_INPUT_ORDER : constant is 1;
    attribute mti_svvh_generic_type of DYN_INIT_EN : constant is 1;
    attribute mti_svvh_generic_type of SINIT_VALUE : constant is 1;
    attribute mti_svvh_generic_type of OVERFLOW_MASK : constant is 1;
    attribute mti_svvh_generic_type of PATTERN : constant is 1;
    attribute mti_svvh_generic_type of MASKPAT : constant is 1;
end V_APM_MULT9;
