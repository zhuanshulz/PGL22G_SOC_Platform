`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kqY4rEZdnCBq8m3VFXDnTdjc7+zdYIdVVIGy3D86QzhLp6n+19Ne5wJ/9PwvokC2
tJbQvh5dZYTfLBh+Fnerq7kWwvPlLk10Rpu10ZbnfOvOTy2ScYTrKLo3xV7xY/2o
jnSKZX5qAdPW6EYiV166hrdMJIgY9XnmHcweQ1IpqHy1cc5XpLPulZaHNrrniKcM
dHzQerCKaJI9vaaB2sRGVOIreUHx4pOU7/UeCAzvJWpt/045dJ0fRfzuq8viemcJ
ZcOMUSaTu80p1/vlFVb8yeK+yaS6n0D1WbMH2mO7Nc9DkIYbuSUnpydTyVzhMhA7
SF5VUqMkLcAncmfSWsCTuZudpypeir+zh9GKbF+jZoFXXIOcFczpIF1c9cb1SDPf
S0W3o2VpUZhVoxFm7E9Y0ivRe4iliJARMevWtPZVrM8ovSdS7Uip0I43uW0PGRAS
et4J4eXqLOaDjlihwHdBsdHiOxEA92CL8B3KKmmuzWYkpAnZLjH7TiVBvUknQT4v
iE4TuqNieQkA/drL1Bepf8TDRVy154GUgwDBGxEBGm/nUTuOUbasqdgRMYReRbGf
SF1SxzluFlOrhz46/1an6J7l7ZmUdx8auLgEbDM3jf58MqLjRs7UJrNrjL4l3xRS
H25xE5E5Fbjv8k8yPSNEgQ/iu7uaIyfQebontswiG9uy9s3wWx+MANWtmOxxUx00
eskiYn3No20qBIA4EiKBk4cwCo30IfMn0l5PmSFGQ9wm3DDperUs/AFTzMMnEkyf
Jcc9jzmb4bNu8e73rTihBZzu6OkJcKzm6jqCEmc5p3SQJhVlFITQTwF5UzKD3TJw
BZ7rEYsISTAt96jYdxXhw37ahlCQvJHMx48DN/z+FpZ6X8LFb1o39YvrPYg5NRnY
DSY9p8CjcPeHbThIA9usfOjPOux98qcjEq2TwYhXqyUP7WkAn44hqqO1+SLJedEe
23hc8bKe6Fobzgb4hmjoa+eCVdvWf4c0on8gfdwzU3pzx+xAY3o3OWsp6Lm+WXSy
wOnBtDiSChdg0/8wQvAfsY3XPKTJWX9sLcDEVtIc9XCLeiJinn1+Y2N1VxXTpdUJ
YoVpeA1unCy2PuCg1fnBPabvYWLdNkJx88JZTk0N3UH1/K3OOiXYAKGcRvKzVqtJ
NOo5ZiLXKZL9Rb3cGN8W4W1C9NdU0QWZp4V4VPqicmc03wniyOkrz/eU2YQr+7j7
P7OysgRBZyLmI+twgooCoD76uTRxPd+iUHLIRR3KdR6ee1hse4G9Zr0mbdrrPBka
WhDu65Hgrb0rZji8ftGtbGtDUcVrbDGD7hN9ubWFIHl48WJJ7NKGG6sR5M3JxZEw
lmvVkpyuqh7IExcpUsMqMu+wNe6g4Prbcsu17DkwSQJZFbxhWqkBnUjuLnPV+qtZ
5pEPxY5uYC9vgyh6x1eVXZJEA8yx13MMfL9Tjnpo/k2t2a/nz7c3SzcQNOoKy4jp
1/u3LLLzLXnenRZa9cOH6t+D5aHEyw8lL8Giq/Zxyc9GWtYBFN1WEDdrbm4GTYrr
r9fqRIwk39trG38+bdv4fiuyCJ64uPnMA+AGfqe+5D0tu3Y/30uZ3Sn7b+jI2to9
1ImmZd263wStyUkSdyabxNx3Lq6AtfVymQlGYNyh4/WpctpIMLO7JWa93XoRcBhr
ypVAdEOzsqllbQZlwTQmeZ9ZkDNqIIKZK3YVMp+UYZDaGcFWEC7/1ANctajeILX6
IwJdcUZwLzg+jmc1S0XJ/fax8h0GCPvhcMKFLD9ShqGrOg68RMuT+mjU0V4jJgJm
iJJGMoZe0ksHh5r2VO8eleJwUXFRLHwH7uYPDEmw1g6vU/OKJbGhTjSUMb2SXNeK
YgTKKojtqXY/QiaMnjhwRdhNnHSlDzyzNa55oqNrjm6ADmuPbbozMosXUFHGRIU9
4SrzJ+En58gxezlC8wEPlCEzXWDwu6YMLCgyuRQIGvWHprX1hLHHA6zPy6ss4W0o
cjGWukwd1tT044j41SqBSqRevhgSS224huKcdGC48h1zPftPXII2WGHxIbWnDWOd
uFc+KTk/Fb/13B8vhah+QxMwT6qK7qnihZ1M/WQ5n9nonD5GIo/gNTelAOHJlvBs
JYNHDqzhcbKB5wP19LYEzVxUEb7RQYYI9wsHK2KtKWxpdwq1EL/mkgVbvLdEW24/
U07yCepa5qlJ39El+W39VpxbDjBLF2qbqt8Tt23uZ/Xxbi2LJORxv19Zk0/j2rS5
PPGO+YAoYP5BHn3B2Zgf19pXkezqVWd2Mwh8Q81rn9mrzYOO3dO5yrKxWm525c4i
tC32+h5ksuFS1KjLSBYm6VxPnq8CzzDcEZ/CDcnf0s+tYA264PwN6qQLIXAorsZb
Ki4icMd8cVcNd5wsjK3s5Lp6yVkRdlv4raOaxc68KE80tdh/NSw852ey7cE2J1t0
VTla4k7cUUy2cVwB4Z5p64vQeQD9sHfwevPS0DuEN+GgMBBYw/NyxBjkA/9ahNym
Gi1YsJLzAdE+f6LiNNqXRhLFvfecy7yaItAqtRAKbwrolwSXA+kxOkvLudjNfwVZ
QE/QuEdBi11fRE3gT2bYLnRurcQ8VddYQMDAAZN5oE5ltrbsmf56l/Fxj1VpU2aC
70/YhFTc7DIrhIzBHN7JdfqeHMSsseLLxLFSkmpp0W8EuyMnDONi4+t9t5rdL9Z6
qnJj8xJdo40cUeUkJhGjJRw5/6Cwckd6sf8KKFG5xfT/OY/aSjHRcm+z1EKiyZ5x
CQapdZnzGnvj878997GWtYj+kEquQuKzfu458rbpa3CcXT0g63/GGTQ3VYWREXYE
0TC9ZOSzUBjWuu/sWNDIqd83FEbV2cQXV/qC+6O/SO/KeB3PFn6MSFLTe8YiF9N4
2S4KV0zW8MPLHIEvzYTh1fMDnL1WV3M+apRCE++nSTT9qfhbPOPVrOfkT9EmqH19
PZt0WBZOVjIfnivnzp5aZ5wVUSocyNnftKUP7LPrZ1Rnb6upbP3hmYM/DekT4ZxP
EW9rG9pPAwIqYK/sUmpAUn+cuFXJyCh9DgZtXhFvJRybRgD4wTYOLMY104poeuok
sEK6EkFBoFDBrb3KFMziUpgDWZyQhZ3bYmM4wAUprRSsebbtiaGlS105yHI8DPkX
P966/0oRESM2xmAchdl2SVsYr2vkxW6VAe0p7y9Op7JAq2ObEBT/SADLWQZ5FA0k
tId0n2lq8EfoIcRSwnfUYdxSq3hyBLKOeIBF/yyfXbYrnFztxrXqpTgVpsEeAD3o
a1dS+Mh42e+j5MmXwDIIdi9CgDWNmskI11Yn8cC6TBY9OuNHUZqWF6V3nWHoiEuw
r6xpUis+RXhWFMq14oANgwWEnEJJfKlswSj4SP0YTCst+aR31JBwj1Kx64w7FiHg
gGIzolxc/8tUPP8UScEFfu5p7pSlgxRrUVFb2H4DXnKOML91aKLikkxJYHnOTaaw
bgUU1DuGr/ZevJpDtp/PnXByGVpLPCRwBf3z57B7XgJWn/6vy+MzTievk2mKUG11
k7T3eByvuMM7kFqAJXcRQh0Ox/ZX7uwEQGRSJeISE392jU+4sXq7rjA76ZWO1m5e
7RR/1cC7vVrqROfTHUQX+3mdG1W2rvhv+VlEgXNOMb/n79pVQqwlJKip9vd6cvwp
nY4YcXi6ZLSzYOS7ILfq7vQ38HDSgLRs6wYD2ICe6ExBZ1iQgUXM1BXyRp4vGFdL
TUFCbfT78p4E4khRdmjRnuhc1eisqAL8aWMDMFz2RMlyN8fbptj3lfPaCaeSlNfM
3sjaibHZc9byNHm8mhhT9sP2RUOz0sklB1qjFHgKyLnVfgBDM4AiaWy3dAgfD2BE
5/vMx7XKmr0rX9rYGyy29uTREEhfHBul3IwpOmODbtY2d2VpRdh6Kdj+RflpPQQS
Ez+AYDDEmVw9kjMSYjXIQPuNAJ1K5t/cDF9O2V4T/3qDRnds8iDccXgiKXE0Fix3
CpI1rzwyXk+FpbWhEMNiznzne74/om9hzu99LJaQmMMiD7ECpPftoSR7uIGuDf9h
0MQlWPr9ABqROOPUylzlMqk2eBS3eduo2e6CxW0l85kbDJe0Dmw10mK/lFI9DyIq
OBdwPRiY+55tUGGuX73WAE5mZ0A8RIQdWj1EDPsgA6/WXptEQYcId9VfVGx7H08O
UYZ9lvvG1bIAq3ENZxMexfLRa5QqqoGxahT+LvVkGgZZM6PvvJNy7mXM9FxglLz1
1lkX33/XwVX6+wxMStESieAUXzMmhYn1Va39oaB7daEccY1rFxv5MsuVpaERsHzg
RSfaxMufIuqqQjbUD8aTaa9xvWc1ozMX1586eNzJOSCAT6JesrrwIS9GXB/+dNBs
yygXatUibGGCw8pQJ9UE1P4lNaGzFhqS0Y6P+4SHdxMPiHhWd0iJs/6a1BnKxbK2
B+3owR/yEpoKODfkt3d+fDjKK9ZWX0LvE9QZJOWkpctFM0FQUZKvZ9VTNWQcHVs7
Q0uSp1BlXfW7zk7Qr6BS4Bnf7IUmhn7mGIWTy++agzfMKoFzryaLROw8iBmCqWSe
78RmtkEpCKlKIC4XTfXyGYg2dhiGzGWIJkvmr5BtZ720/t7HC7NZUhDBgK+sY83a
mTZV0AM2X2OlBuWh8pUC5XtaJIIYSxmrtPqiX0vMJ/Npgd2GAiuL4Uvp+A0391HW
OIL55iPSKCVESxbzIwzQ6OdKImNvOKwVamyBKOjxDt3qbM45SKVwnqpJr4nfwZNv
1YXaIplDu1Re0TKc1d65HqgNOH8UAEokeCC5CTcvKI7GhtuUPG1sge+CfN7KxLZN
nu2m8z0XsOpLwnt7HYPMqg5BWBmAaRcd0E5Sg3/+QqtHKNo0bRsPGW9+pOII+Ipc
CRbCxqIhIPYWIOXsbAVK9nkCzIZV1ArR/txxs8v4oGSZX8TRRWsMG3N5Axl+r627
/1ECs0Ksk9v4cJv3/ASipWy/4XtcWJQtSgLHKfLmMWugVsKLWj4pd0wY+RklkMrs
++Trl+zczA8Stm41MqyPZc/TgDq3s74XI9Hy33i2mcdddcNom0kbPlyDOM/hqZQf
2q2X9OigfQt5I5efnbVPrNfFLRaz4Xh4NbR+LIcsh4DsfOZXdhXR8bHJup8hCBrn
/2JPiZF3SO6MTZttMmuF2zw1ilD1Bom7TKQMmhCpzpwbKV0/IuXpRbCOzs7ogyFv
ldH70Q1kq+KLs+AikQErmdekN9LF94F5V2H1mHlWdGr7FpWhi30e+SK6F99jk2Yu
ucsaQNYKE/9VPhX15bxHgUh+vldjyDBCKZ0ZHVjDrb/SMQHn2XAACJpbM4VsZkzW
Nz77pwfI6LKmUvWrtnC+JMjOixcWKyRxM06zOKcotatpgA/1lgMsHBOKHA0umdOY
jPbTsKZHWvPtzERAp4gJ+No3ly5j6eigLzsZiPl0Hc+X21mXpTXNt9kEfIEhguDL
hCk01Nlu+df0WUmYryc91fn5KX8fdGndbiuL75Q/XYBtWQnhfwaUtEbUuh0EBIAF
w/zE4nP8sRoUXaVAp/9tFMGQT5yhTb8I6P2uZnz014tYe3rI4jeSfJxgz8O06hBd
I4RN0+xRCYE57A9IRqJ40g5JdFx+xv8LvCv94jdhyR3ECfFmE1/xgpUfw0NFBb/1
tRQ1QV2KhwYVAuV2drmbspYPaTaUnFkLd+CnIN70Ey22WEf9gTvozX7R0k9XdjQW
E5etEAScrBDgjECj2FK++jiqHnS/1iUti7z4T2S29PTytC3XwLT/5uXmLKvmE87m
m/ABbirIXe0CSSJpZE1+/IkChBODNHGRbTzw3MctcbL0P0kK3ybs4NxDn8TIccYQ
WunvMPbnNZi9+rzEo2g9tOJeH84opUoBv6pt/uDwKNEgWEK8lMBErh+TLN2GXdca
fcyM2qFHlnvr5rsXV+E3lIELUOotvYVHIDpjKN9kwjLPR+97CTe5oD6/clvDPDkO
2XTNg1WlvRnFuZVQeA16e4eZ+EcFxUzJ4e2OB4PGfZyoH4XKDa4vVRNvC9Oewlok
px2o7oZWxt7U591tuRAzNreKqWgQHYHdcnqnNBlEEYDG9XOwSPJhBPLJ+/ox8X8J
s8kP3NJqZvaYKPcsdsUCbxISQnV0itobz9n7Snt9khUGnKgb9CMR9gKH9d5YdDyL
6JsahsETgnSVqrIvotHrLnYBFS6W2QxKoEtHQV7YDxfW5ZxlVZQKVLLJ9TpqH4zg
NheoAO3fCb+syLn39FHIM8jfxhenmyj1fi5rJ1qaamJrc5hoC7uEr6pvUr9ssRHj
IaJVmgCaFzdlrmwSdO6aaFd/Xd2+aFWAKbgtamN5zlqHgsBI5Bn8UZmu37QlAiqF
aw6LrR9IJVxvPoz74xoADK64kCoILzOp1GRKDxpdMuD2OwU9f4OxlB3G5yVn0mVE
ZbCupbP+OO8DxtbXorzB/VfIGr90Wzc8N0sH405Qu27Wits0adiAxzvUMReZhZfQ
SP/kKDgLM6wtEDU/B4FArVkWZsI+LDjwPDjuOAPbSddxHMc16zEplHfsWhAjuk+E
S2WwE3uSM8RI5UZ4Mp2ydvYujMOjl+98iI2EVlACBunqI3YgI0LX30CP/a2rt2TQ
+VgLFzvQXspBVAIqV0n12vgwXXkPKOATQoaQzgpuoIpJ6ociaOWxoFRC9hLse0ok
sMdF6NbffhI8a0Zuqm6L+5ilHQFGi9JgjnsvKw8pkdjQefHXRmIJYHXosfSTRAUW
pD7M91iFFnvjveeozmn7BEaFsxdtYAdy5O5rgs9EZzL7pfl+yBrO34HJYYDv0VTZ
1DBQcyhbHaPKioq9Asb4EgtUVsUMHT5Sk2jntzB1I//M+7+aPPOMGTYsQVHaMGDi
4e5SlWkLMIvudzhXWsmNZKOWV5Zskqi6wVTvgQa2G0ZmGwoF8GKHSopNEif4pPsn
BKxdImns9fuCYOteFshMeyI6tcj/SAsBdsCbG6BqeSEStVi6nMUu/AfeEGHpsZ7u
qMRtzGRJB1uoZ2kkZHxXgAxLjZuJ1DqMDk6st1459GqLqdhLqxYiYz6MvkABRhDI
9N+0O5nAEvAjnaGwaWwsVYC9JIuehMvWI4KhF6vkgYmhpKGNDGKw5ujBSG150Gnv
60Y1zMNnXEkm0vzBbbdhh63K7Q5TpXeDfV0S7tWI/X/AQVAoXDgwzbpn0tIYTQCw
Ae1JrxRvBl5TDa5Wj7Cbe6UbonAMZdx7wRl2ZmKY3iKszj8Rx95NZLAvak9VZlHk
QDtkDNV5rhqMXfFtp+jf+GsL2wNIUZNAwIqbF88ZhH+WAVdz1yOzOd/alWmz2JuF
e5gdMtid7XK7+8YZgwW/SXfILvhUA+25y+NT3XVUxF1BF/Kc4AvO0Q7sT3KzcBYM
wY3g1hQ1o2zgpJVEvWFvWuxymVbo+5aqDIV/FoB+UIYuNmUbFwGA6B5VRB/W8I/D
dipQNmOVI2zUVZeMHZcqgXSpuBNnEioGwnSuI8cL4vK0FfHilEtTwo8E6liLi2Xz
RwQvvepH/hwp/SMjdU67/u3LicPzgbRXCKSX3lgGSIwLvJs+Y+tO/yGx/gzxJFcb
cpmam9qxhr0zEk2eem0wHfv1n7AnZLzpjsHoFMTmcfZLmgzfu0rffXypvA/Fect0
Fw9WGfpxuKp7vN3WCzSUX7Hu18q+iKeS6RLykcRd+ROmNzwTfgQRQDvLv/EOBXWF
0Ri0qpZju4pPzFZTi2ZkQZtyVoyMWrjmsU6gCPbIhCwmDNiFXwLEoD0nSpeyzpU5
jc2y3N1HK4YXUPPdiU/i6GGLvvd5SK5ZooCKoeyxX5XHqU+NmwaqvPbh1/BUKina
ySg2/9Th7P59H+cCjzLZ3d009xwJtSY73/Dr3jkwahNmxf5yRn4gv8u5qR5vY6tw
zwQs7OG6tLfPUBtgTZ4t9Yf8/l1ZAn0QfuBzv2CBUwTc9D6zPOteSesCsSowGIkP
onmXF9THEzeip1R2yRQyVYTRTMX+Jxbc0jCyfHBS3PWHdLBHFDLKX6n1iaaTs6vE
C8VGtMJGSpZqBgplOTjcIiVH3ZIuGxrZLkw2NlwU4je/ZBMs9jjjbeNvvO/5xysm
95TNbq9JEu9I55AXa3112br6NDgnuT0nOC42WUOO6OqR2gnJt5a0tU/lWQUQmB9b
96KEWED8HHWk1ID6SwGfcjl2oqiWc00Faiga+dF+jaoOCwS6cF+CyDLRo4XtGmbT
j0ZdN+YguL8xzPKvtvKXbxAlKLXvrMzbv7mjV1sAduSBXhIu55AKM/E+RInjKNoF
20RhnuiwfpEMAcEkYva6Fa0FtTUhJx6vcDF67RymE2SmpYkgDITk7SMH3m5ah8pN
QDHyjQMnXgcgr4/9HPpfXMDpQcQIwUIYUKqbx8PgOigw/0wa+EtkdIyqaV2lG0vy
Wp/XxnEpsJDWvZr2XC2SNdGvqeHY+LA+Y4Y8adrMSoEeWrRN6tmRJdG94YBN0Zga
/Kq++zMm7V5K9l6VI9qhT+rwLouAbOLreamjL9EM89yKjZs4m+sr238AbbvztaC8
BuJRtfX9or47mAQadBFjFl9AI+kTKoMD/X+BMPpXXAt9OFLC+gJt1tqp+9/k0EmM
xeGN2oB83NNzG8FoIzQ+1vu2zyOD4oBm/yAH2gP0eZMlqHADWS1dezp+YzelC++Z
5HB5pZgrxilSJysnqRITWZaMz7wlvqgBkLR4gyCwyn0447E71ir9iUNhEOSMjNa5
0MrhR365GuKE0GlurLfAS8MQdQavIfmXzrRMpbXkIJeaUK7UL6W/9CBWz+0BcVs8
EybVoIsTBQjcekKjNtkCQ3Ywv+Pr5V6DCj8YFmF6KlR/zIweJG21SSNrjJpp52fz
ch0QW2UX06BkQ5V2iv0Q4ApiY8E7xAndYIVKcUCy13diATmk6GXJ0FS+l18hZbph
nPHtaEm1nwkp/skgDaTr1b+x05LzPNc7uhV/es9H5MuaKGAVNyWh+WB/A2jSomm4
WvevCv7WL8iJVDUl/WaWHivjvFXkl/WMKEt1MM5uP2O4d1LYy6hA8p/syyhRH+S5
Sn7cKiZ63o/RRX7WNkN6g/RIAt8JALpHCosX5o97vewEiLoIgFgTgHbHDG/BJryL
UnDwzR9AKOgxIL9NtrRfQdZP18xRdIRfrRoCGTcxS/8KXeKdTOmOFuDZAeRPQmwd
835POiL2W3MGMm0tb/K+LRV91qSYxlnIPKGbPLm51AzwXz7LKC4fvzmhhrd4iuwN
TPwH9sJPircwDcVF0w+WpYGA0+8/M3hzUsEz9YLNCZu3CF0nYfLzFrJY9xFCsHNu
Yr40XlsQKn9GSMwGPWD/phQ3sVrZ0Q+afCLuwxbYepRfclRl8KGU+lA2haMdzW5N
pykDALhRhqJPz+lv0u6bgM8BeJ0nfBnaqDKjWZbFtzZmDoP8YIb3kDc7mxXsMS+j
QQv125LMGkiiPp9HjlFFqoTPmYk14L29nARYwPhB4Hhk0la187GokKCYKn2C2+TQ
8GXcZ35Eupjp4RLoSx0Z2kHw3RRlfsHpZukyCvAigLuespBwtCPBrC6yTWRoI5Vj
lR+0ZEo3xcphFcF1IPxX4lVNiQGaZ1usHzY6bvw+UCRD+rYqaF2Zl03Jb3SGao9q
3gbSqtC16rkn9nvjpWvEp++ydq9IGKuLsVkaMwh0Q/p2o//QxVFqSAgCnvwE5Tpp
+jdBdo9hbRvmqsaqp8nWw1ttDEbaNtN2mXwIP0jEWxLv8Vbk2TQPs5PG004kGxR/
vN+xl55V8sy2nZbQJn/9iVo1q/u5sqMD9YQ+eqrU5SxRuLy400h+VgFAjKWq/7sA
5gzUMBoDAhdN0yFuiFiBuNyQGiT9rdOGpN7OSKz6LnNmT+60XKHN5yrsABEtm0I1
q/rnDxqfdyncqzLcAL1gGUJFh7uVkFTs/YjURNoDg4Er2DZrLNNTJ3o/uUuhMaKl
ykbyZzcArOne/EnBPl3EFMmK9u3KadTK+df5eKtmsIJnrtGWecYsYfZ2MThxzBuA
Htw/hSyUeZDEZi7ZtJ3WxI6QHW2IaUJ5PPoUO8s55h3raWwIqSQ7dp2JZWursBSb
3UmehAPXII5KiYSFv8H38CfTF1SzATsAf/kyznymnO0xzK4bXem6JtDcySw+uV5S
ZAOBrQfR29KE1OFacjN61CMK1dBkxn9rarg9WnhDrpGkHYq64B0QrarmBJH3BfHN
kS3/ItXMrj3rsMCMyDWWNQYtSh1vyO6Y7fxiDOUY8JZEW/2VKIK2oZwuTIiIYBnR
07df7tnIUCoF5rpKwDfYy/Xs/lSmf5w/7feb26JSgTQm0FAyGrni2LoT6BaileVI
b8sJBu63qZBbATjpAkWIoARPhpnpGSsk1TRoZN9hu7PTxDjhoWlilzLHbqIRb/J2
xeUsjhMDgY3DEE1YIvPqk+R3pETmFEvTkoVhj22aH+HFOmH0ATWe2OllvWIm99DM
bSdce0vPwiMoRUB90i+qp3IkSY9FCDyVr/umDNNhy3aXz9Z6OPfalHK6aeIO0y5e
RUZ1eiwV4bztJxyVrgDwUnNtVf0bMvQArXP4Hxevcsc3eUM26i5soY0srA8oWV/e
LEG2274c93Rd90jPXgwiiCN+6pUdrN4rIezbnNq+yUE9iXor++GznHRMGSXK5sLk
dIkP29/2GNZanIBJT47P1XLsIzaDVlrBEI+9bJj0c01wafIc5PnUH95qaFP8d+tL
eHpJslvzO4diqHY7gxVJSSbAe/s8z1PvkqG/aTmgsdP/3uf8GNONyYBGWDIsBMtz
b83A8QkbeBEtnGTsgtqYRiMJbwlRtQDrXBX6TVpZE5wf7ff/sUUlC75vmfqy5D8F
Y7UaGB2M39m0F16+D/IZE4o67K67mAOVtU4Uk/lSM0UuuI09ACHXRPWkmxlQJVqH
L/2w2EMwL3YpqOU7MtEN2Gstk8DpOgArlhF+QSGbjTAOPt8aJTWpN5Xkuv6vFlQ6
vhdoYAomNctkyaur0/yWUm/XmOIOoFZvOTxrTxtAJZZGhY7jn6cyl7yx9ykA8uZa
vhXKDRXf2Gt5CXOBAwQ/73EGS7a/0K5QW1y96XMfHDqelFnOvbBH5lVWMlBLKkdX
5+ZS1Rn8PPliUBQ8lkIi+Zy2jCIIaCFiZ4Qb0Huzp6KVHlH1oB8BHqm2UDi46MM9
QLxanycvr9alw8kZEIjPbaZzFRbQVlqdxWkaldetPztP3ooOi4VVUJsNxjS4v7VM
BAg3pbgFICf2X6dhYir7APf0F9fwPSDdbHn3ppeTUHq9mLXBJslwXeYf/MTiarSP
VrT+SBk0IJxf9TYjgJg0PV0tzzcqRqGcaQ5Lto8VnVM01ZcjbcdXdaRxu5DjMvmi
aeQ49LLzjOwAx+snxd3vQAHdobhuMjhrBEsq6fchzeTjGZEOPSdE2Sy9/0iRl8+R
umnGV2i0DDdbTHDDNuboL5m2TrAZN1eLeTiQ7zUqcNS5A9WVE7KkvcuEkqcYfjg/
+z0halMmeV73iJv6yws2ABxLGEsU+hWQQ02OLug9VBd3wxInY0eKZc3OQBks4C/9
LQqS0z2XBN22o52HBiQOgbLmPUGkOK0CkO6vOh9pGUP8p1BlDm0qiXZ6WavoUn9E
OzQ2JocEMO/LzPwrMQpFOTlOld/JLl7RyWjQcvBsjPwQp16mT46wXHBM/ZlR343d
x/qDtnd5UJ3zM+EOwh2abJdk9iBP5+VinodNdSabaqrFFoCrm/aPmjorPSX5TcS3
X0NLIhyn6BGXUTu3LTcevdaR0LbecQuNFLVJAVzTM9SazZS/oADzK5fJVUqFjyk/
X9nq+taOQ30EAMJc8j3NQFl5FwRD5CkrwFFHDxYgH5077lQQEWEKNU9PRDitnsRc
td+sW7eVAUfhO8Rz30fJHy/TqaSUTQKCk58QIe0mYRxRQtFizhTZ83khV1Bdu2lt
4h8x1u9fqZcG36SbslrDT4aXi85LmVxubunHQJRz7Ys1seouIQJx2Br/I+kXVvht
bp/1VGpUpoFkfn8FxUJXsx/KKkRgRTzGAx0/LtlROCsE3dYXeiR7d6b5k/HSq77H
URegEt8FVth75VNLgk9Rn4cewwcDt84JUy5lGgU+kTHMblyzOUc3dx3G7fzIUbpg
7If5rgQHXTrPvhyGg2LpYRFQJKdOHjo/JhzHbLt/Cv4uoboWO06ogYOR1GmIIoQT
AcOJGhoU1N169sTjH59X3T0P88ogd/I/JTyUjroCp8H1gH2H2Kt/TucX6RUrnTBz
e60Qk5yDXXstgEP2W3CLfZYLWkeErFYVmck/54X0NUKA2wmnJ7K+rY+Z+lwv6OmS
c6cYF/FtJuIkCsDgydanhA48advxgM0VN/Y/yeJ3eEQ/Uos/poJ0U+YJJTr9UVnc
7SfHfu1eOLb27DRm8g0ryvTjrv0foaXpw6kpF8c/WuiTGGuajC9WMBGAIerWcxpg
UH/kgfrz9Yp9htLHThu9j9kRvIUiDv5gcJdBXbA7eHOajKA8JOcSRJRa3UpdvwZH
pk5CNPp/YIwuGoHy2foHBFVfQwEq1w9rODLVzb1j+0pTWAJYuVrPAjQSEB2o/osU
BbsQbAiwobnfJqCsvHr2ihTGEgR4pinPxVgvuzxRvc4btc9xSWmWK9QNK2ik19ss
hYcqjQWucAXuXSqt3OzmS2S+2oeIfL+JjjT/otu7WqZ/UueOy2RfUgBGTLSKloDn
6Z/GSGDOyjO4+c2kudJ7o81nU1jrTKW021JngQrMLAX0p9obYcFQttuMzc4ql0DJ
fpOs4ujQcd5dea0dScv1m49aYpTThnSWHXbdDDNrdn8q0ZDxjVU6FQKFxIfGrBvG
fQWtSVq/CFxJ89ozKRpIlZH+jbO5l/kp/8TpoSGXXpmbf4SP5X1yTQMV2BRx2Dbh
qXkITkwA0WiEQ03KtzWE09cX2S518TWNhOqdO8Dhd88TaWgRvJd2QsazGlxGYg9U
faFKlIFQBVFqi8e47Rl/4unX3u4hpFtxZkCSbTknMa7tAiChQpGu7CNI7mfuJwRZ
V2vNeo44CbLq+dGvYfFtOqYwzd8oCn8/ABCFB/WzXX14Pxn3BZpwX9zHhH+Iuwre
6WVa0QZNYdm1pQHJJS3bl8hGBuPfdnDsYVaQ2Ep3RSu2cS3ZrBwFkatKX4of+Ifw
j76OrM6zvKYToCzfqzeVhR3uAe19tOS9r0z4E8t2A9PwD41OOyX25fcBWprbCKX1
mleay5wr42UxCVAS8Y6mzZ5L0xgZh9h450eJNHkvwyhXFxNA2NrQ4wtHZoGFVUT8
zcjoQlO74psE9hkEIz8zHLnH9UYVpNJjuW0+lAtSJXYyZ0qa4IrvE42jDumK3y0O
1dFwkr4X5GHBBAFnpZUMGJk8tObwUNlH/ZyD7jtgol/ufqB7VZaAlabPml1sZbgR
92i1FaruO+x7fXob0lmL3ekycTYeBBzzP6AM51cflRdMUhbQhAn0WAtR2X57MZQE
z4xcikBfTqKm3AYGUgyLLkI8NwFoPje2U/QciWMEpyGSHBRic0wjzPy6DKZf1WlY
GVX2l+kf3dISrmJHRUiTqmw6RoPo2SyemkhS7iF9ZkyolM5sxTAyWQMdT0fBDFCd
TiCty76H1nR9I1Anwd+92qsUIkEfyySb4+qkEwIU/YeydQVYjs2KkxH34HWeGuA2
yZLpCVWIGRFPi0IkKiMBrLLaPPpX/SECdOABcxX7D4rr8kmYazqWn5x9n/d7dJGR
WNpug7jI88RFTNtw97M3252Jp8v/DWJDXKwxexFWg6f7LnhXAU+SkALodNprnTHl
kQsF6ran2pgqb6npLQVTPqvRFC2iy0kyzSt1MXSsqgdyu9CVuEdTriaXeD9CdorW
GmOvuYrUQthzbxwdBDfE9HN3uHzfhP+KBrWh4XygtRr60QdI7fj65gH1R78y3VwM
0zsvcDEVgodyQrpgphHo1vRoxmyp+mhDcOGCX1DvVj6rlDute89OPn5PNV8lMATT
SkhxO0UdaNr5yy2SGAnlHjZXhNfixgOsJopFrQJnaoixCwlXaH3XlYO/TbjQL7W0
JD+CVfU9M+PxWMoX/aJjAFZABHOQIWdWFwtAjPm1D7CgaWDS+aMZRNb77MEBlj33
ooGmGlFUIcudrC+9cesdL4UHwCwKT0VqTPLXswmL4Gc0j5Vtb7HStUWYafGJMsDq
1O92JgGAx93bJWcLK6d8TeXVPlVY7n6ZuWAn76WSoh5BAl2puO3ZZe3s81Yx0HCe
zNV9LIvoPTko1eiCd5Q4ImSbdSy5I2/fP0WE5RN64sjjhCzFsnSa/MIdPy9KSY21
Hlm2SqiAZae7RVjUg8IzsKraLQiFOfgzJyUwaljjlNkfRYxZx+KL9YXhVXkR+F2A
gmGLbaoZbHtQ35xxOmqJkLzAtOZJ6YTPL+lUTGLI1jjBLFzmNsTxaOIKfNFRW24Y
h+MRjwFA4KaV/BY+moBA9KlEOrr4CmkepHcncRw3/4Zn4geEg41T4gCt/CqOdTs4
tB+eewYe2VqNV2A+OfV27hgaVh8gE7RdNRZyFx0uq+kARNKdsCtHjQ8EO20Jk9/7
1ooHXVXh6781xFjZNuxE5qLdhvd8eLq4Sy0wbsdv+ejW3h5lOhs0GFKW6oFDZBN6
AMLzPbnruHQLzmLoStiN1bEbdTa0OuiNJ8SAh8d97h3ZJ+9C6dw0fWFuxLPTdpaX
zloM6Y9tCJKBY+UPhJUV3esaL26jM6g34/ENSIwmB86fmsIjej11RX6wjNR5wo5z
7jtHJQf1HgsFLqt22+7pF06wxAbBUYOyEwwK7fg1CgjhEpWIfmI4PA3WBY7hzELz
SRsmg/CrS7WxSSr9xolP1W3aex71B4rJIbr4huve/OwIG5dzutNg1sfWsRXUZlPp
SW5gj09K4z1Vmab8uhEfbguZkRAOJCFFMvCRlC9ZtBHqP3yXDbSLe2mqze1CVx4q
B8UrqSKjsHsMacwsTMIqytZO0hsbmsf2rQFGbR4D776Jw60DsfGB/G6fO1wCz+co
/dsdLsPbt8AUzWfHnes57oN/0Pzq6hBus7ThYvSj2oHVS19oqV1Sg253ajofweMy
NuOKkhnJs4W0UPKy6EBeCAQiRJqen3uYpAWbP47ForX7kQNrDistHdFOc6GpwqxY
s67cEfJk2cXZuLKNMEgt3P7YMRW2q4J6tAOFy5KsKWNbUb6rW0XYmiARJuGl4iGH
NTuqq6uXL4KmBaQbhNITI/nuHylXaf5Za3xAuNgf5VUSqYIHmiSOuYkuYFA8z7X8
+9n4dois8hErqqCgaSFWckUQhydzrblOTLqm6RAw8IogGvz/76IpUGBzd+OdRf0p
vZytwoEpr17JpQWRUemuHMPUkvOcLRpgxhuq3mRTJbxXVNn2zOQSG1P2QLatlul/
gt4fiMZTcD7K6JRRTyQ6VTo7XZ8F+BVT56n9yGIwzydYorQJ4rr8Z1injifD04fZ
anqrswBIxqQp09dZz1W8/RAM2O7VopZJThTdFOua2aX1OgRmXzLu+qpQYWJiXjmT
Ae+diFh4A4lIcZIllN74vv4+8yawuZkFjIlqCbePUuvxJLb2fCx+kAvLFQKO+oFe
GV6LxFerb/+hv1c0d/XB/F0fhOnpNNPu8XRt5s2c/vJgJoGO3rXISZsBQmvWlS+w
flkH2Cj9I2qaRjwVlKomcO8poZ3ZLKKuLjvirL5wFBrE8RsTkd9Qzg/OWrFTgscr
XiRkzclZPEA8wDydh6guKM4T3tesruWjRV82q2jTKBFmdxpZNENvvjgtYRyCy+bH
1tPH3CBgsCArhIlrRC1Df3AHTItp9HlE2hfTvFdFqnSfbpzhF0z8MGZ5dom3V4jE
N0bMc2XPIHN1SVC/PgpWa+Vhs544eeIafHdi3VpUMwDpiAgQn2VARMqbUW1JCCEW
13bsIr7B+ZSvCeEd/vIHbZwEUnlxEWfsXCAow4fd7YkK61MV+XhFo1SPkswTZBeB
v7gw6mqU/o5wO4wPnwjmo0NZiG9scn3BVEpx8h23VlBedsYRyULy2AQgJ1qpq1/H
8BSnAAJiEqhQs2MEdREN8CoB8daU4j58AxF02NwmxvelNHapd4ZgokOT1oBu6dXb
afFpW/YyyWs2MZetpW2kQL5Y+620+WN8rGaypJOKYi+o6lQuQb5uC8FzQLInd2cA
o9zKE1tX5Pe61LbCRtQxKCERSoYjB0a3SGEvisxT6todSvjC5I9dJU4SHFi0gsgA
QcMQZNowgco9GlL3g9RQgyUDYxb3OF/IWHC/yhXZDi3e6qGAYdzLCsWeyJ7Udyxi
/eVgUlm4UMpmyOFj7GCLdijOj+SRsjUDJu5wuqikurf8v6G2jOWhBZfylMJImnvg
X2I3zAheB+mEMqLI1IjWlYSFAA0P81JI7/nVpujfIvlzEP4o2P7sxLKQjaenwSuq
x1LCtkjn7uHE/L0f4F7ZtAL0lHmFqYLFdmM7wRRuZa5GZIVnXKV8NuGZAB4kzlRK
Ky3yhtRYaEKtLmSuiXCDTrQoyJURiOyF0TMdxaFfKea2kSOx8ePnoI1e0lu9FQ9E
p4ZGfOa3U7aAFd5kgYkUBSXwhJlQTCFS6tBpgkhCmOR2B2OLr8U0jQEmZjBJqzVl
Z77E8n4TjjPYIiIw2z7+w+Ay/7HNw6nptZnLoTmmqKh3iDYSrIFW6ayBHB/jnKCO
MCQTTVh7g1LMFMi1Ezw6Iuqm48dz0ToXd0hjk+gqoQ+4OjW6ng3+nyPKu9SCg+zW
Wq4SIFzMMTcXTgIywcYgIb3LJd0Jxbo//fCk4MmBj2fmIDN3rv6q+su1wlcAZMbo
YNugmosL1IRyfl+gQFz3lNqlrKlCidvfGmngg1bPxZwVCcVJ+YU8x98FWmWPIP03
OO4fz8Bi587vWIcIdrMEUkz35mlWWQfmManTVSuRZff3IBeMJ4rJs9r3lZma+ny2
lRJaC2ENhqzVwvlByOOIOcMMVjB8rVhS7Au355zyuxX70kWZuU4n3ghbrCR89KoO
wVADH7JfBe1LEtmBnokg5I5KifahMh8KhMtL8o5T8ANbfcUrCq2YzXDrGi1faguZ
9bC0zJZ6KvxazwwpO3qH8GNERsVf5qwyDBdu7AhYFUE7VaGajmTE/ICi4uzgIvZl
gQNkFjWO+HRVFQpI0bvSEh+lUsttBPUXut+URp++4sLpjY7T+roD9xhuVJsxlS4v
2GAC+KLRGwOrH0DZUFkRN2/Hm9YQV67+D/gN/v9WWBlJ10MiWIYLNLVzHZokTC5c
LGZTSjCvRD/YHGDnuOoGtOQC1AUTGOXVM/Ij0fpX1Kc13etcizNlMILAY9ACMQNa
YAmeKVy/9948Z8uL6pc0CdIFaew0gxPjrXGdaLSdVr4T/h2vgJlmPoco2ms1o/Jq
uvAAypt8wVVgozQ3TpA2Q1DZCY1v5N3Regf0NQHfUVxQjXzJHZE+6TE7GQQcqdW0
4APSDvvN76jnCPjmdlf6P7MCBhQ05GgaCkQxf8S0JhbzrfE+R2uEyPTL8XbB3liS
RVmrJN6s32Q1WXm21cB13bXcJs7aeMZgt2vpkQsvC7FDDoo0l0AvCjmV/jj0uoqe
H5qQraIm1oH/9e4x/2EX3wYRDP/piES2nwwfKaOhDtSiVgcBQqTeenDAKl2uSbIU
pXQIPzlxRcEIejbZIoWmzPH9bGKXfyLK0schVWvEKHecDL8n360R45bEuayjYyQ9
R7F20TaNdlPPE6s2iPdcQLQZDOxQsAtGs6K8sKHDy/Gp6ONL1iT815PFQNqz+Fio
wkl0E66vVyJCsNksJzOaCY00o+uyHd7mW6XL7fc2voPnJ8XgYSjzZmoJmrnhu+HE
Endo/WTHZag+o4d0hDfOjCfZ7m/HI0hdUt3w2rGcUWPKwfI8f+0XmV/B3OhL2wdX
P4kikB0cZ8xecYa0AHijnneRhkHrjl6fpc6fb6zkvXSqa5ndUsLA2qiDcmfuUuLZ
nTiOu/kyHW6ZHXFIHT2g5b7VWWbXgYcEzHD/PHjjPgD2R3xufupIxrC9CKpTLd9T
7MomramagulZqpXHZXvnkBiBrUccJGsnoFmcTZcnu7Oyh+LT0nawCtXhDmcNZ+Ow
8YlqfEa28bmw4IGoE//EMCz1PXjeuPpsyq+tckwjtUrIsnvEKWORBaM/IShhyHH6
EuGxDDXk0ej7aPu7vrb+96RjhTDQVr0xfwM5n6XJmy7zJ3A0qupgZEy26mm2XhZr
ajg76I8r92z/PWqPmDx4hfd691Np/9GNS3Haxnj3dEsZkikv+swyXvKnBUcwMtVl
0shRt5DJTn3OMd7CGXO2bK5ITyyPxU8YF7XzevXzX4RqCCaQmySHkMeRTtj163pX
rRW9Ny95KfaLNlmMWP/YJIMih+RCz1PbnNAmo+O37P8qz2wDctUFqgbDlcFmuCDq
96Z9CCGFb34tCrl4H4vq+32XsPgC6miecmRJWH6ibPviu6IcSS6vFfd87A5e5KAL
ff7mMIxP08Tss7+bJ9qscpppb0CMIPIgW9JjVioKEgae1jCY/rGIanbKgNlt8X1o
3uJ6E83w6az7VQxtvQs0zSlTxkuBMx/GI1IUnWuGUK6rEQ0+V/BsZuu48gUtsaER
H/N9ImPOjxCyP4d2qCeGbsxqpnlGcY8FkJyW724HTn9hyzFAInpg4lOcuy3uK9tP
hjH0lcIc4FGj6GoFCIUEC42Be1DUTQxuGnEenOPcalBY9lAHCWt24P4Da2bQLA3K
Aog1kA8CRP9QfUIGuBo/ZWl6tWD5nHScr9MXY5TbzQ+auVq24X2rfcfxaqgWQ3Zp
oMKBzQwypJXBCY0rOssFFYoEvHXsRegfITRWfjixzbR+3klQQ6yn1ed2RUEbGWNP
eV/yc/FPNTeJH+vnfHgY+uAEEVUgHJfORLvrfXIKtLfZW68Xuv7CnADLLvHXF9NJ
ZuOvXHgQfzJ6bNJN/H13kl4VTj9OabobmPz7gNiPQmV1BpU6btBpE+xh54SvqNlq
cHYy1vLVI9ZZq6pVgajmycIuxTPtZDPb8VX9wyAqAY/+jw4j8B7715oZr5toVs2Q
2siP4tpZQVwLtolxlZyawk+AyIJgH2MknZ1WeGw1fIIoYDc5GCWMpy3ciAxxT9nO
fy7idWi45J+gz464PcPmHgRvD7R1DYekBjwNQZMtwJzlGcUPitB0We/FO3GFIF4/
O3PG1r73cIN7VDqSnidfIO45+CzCRZhS8mab2Si0hLDZMdry7wEuc6l02wY03aDg
dMh1a+5NF6xmV1H2da9dJN/U5bwo79S9C09DPIt8EqEeIYNk7f1RaROQGpkvKCp3
h8/kf3z8t0/4E9FuMuCj2KnryUYvtCXLq69Kh3sb7+13XI1/N5LRtEl6B/ktnPba
z9bO4UrtMF7B34kBxm2vgKm4mi3Ffe+s3rjMkIgSLeLD/S3n2XOpaLHJ9jCJ/m82
wLWbe316JCCnH/K6WXF5kNkJXlTOFVx7Lgmh4rfayFfgxzda7hjSruJ8SCxz+3+K
FljXqtrkg4TFaSQnd69d6edUxtUz31EMbFrMCHrWdSXGPwQ8zfLE26TnejfhPfpO
IuQ9KYhhEOqyHLCyYISo94aiCcLfHeun1yhLqMWiVdY3/fukavo3FzMD5rOeXGF6
tWxQn9Ayr+Da56nAYCNGOsHQBveB11RlX87NLB/rihHUpeBIQsGstgM1JwxkgYmo
RxpFhhcvkNhVC6LWz7kdmURK/TGvVc756k0xuZY7/tizHdOAyohZwgIQh3zm1kas
sTRdkxbDgFY1Wxf+dUFZfhy2S06h9clFjXVP9gUbMPGb2OtJFyiYw/GVALqV6IHo
TvFUWbDp7Fe38T6MVyK+IKE6nMjXyJhsPwh4YevlrqD/O6SSvot+3EUCawy6imAb
olKmIyHYxuCBeuaPyD8nZ8cj/0R+nqn5F3C7GNT9dEguKZxPKeufM3bwxLy3Foix
Ac0vmDsq4LZbGbcyS1cNhc1IVdYFRzEgJQOGLTSkLDCZ0fOcLGU4yM90e4eALw4q
KA1whiL4PmYR74C/2yylqbzCKwhQFh33IvEODPZ1zF+wwHtSTiPIOpTK4foRFeuU
2j0CVm5PKX3/Zkjog3QHbCpG7xrxb7uvmmv3H2qfcB87jamg3uSKjmJUxiUcEx57
5TMzaZICH7dIG4Xfqi+oeQ/xGBCiMFHzMVaMwUiZ+ze4Vryd/qQpNL+u3so4vtuI
jaCA6uRsS/56Q1CeoSWtGk8houc98dPpelrcb4SN6wERZ4pGqRsL1ZlOO60tExpF
P1GE7zjdZ/l2X1/qj0sSugpFEGVF8Dn98ldAJFodsnAkrlGtxgxuqecleheFmLvr
r8zrJdl8X5tE1+AW5+MBPtvh+sG6qKNMNq2A5df69DHmSDE4Nqw6v3Scd6fVNUov
ktrb84GHBuaCDIDAWjtrxPazxnXCIPF6WPzwp3xAK+k8UtLRbppHPz/gCmpF4KGN
dRfjlu5WzTbKIxYVhPDxIfAC4kVuYYu2iAWwzsGUuOea8LskINV2pzjxsAaxVss/
SK8EfF02CKeVHLJy5zOX37E8Cn9UF/e+gZ+efwITOPvRyRlTLoeNnbHZnNfZEilc
uLSoGDUfecWTnRZxcZr0WvG5IGp7L4joYr6XbAU6GlOK3bHxy5Cy/SWhsvOiGj9y
B+g4C8jegAf4Yap2SRXnAM47B2l+ScomjNNq7Ribx1u+oXBhps1BqOww2I87vOg+
Xd6LbDqvZ4faOElzkbIF2zuyTcw0CuJnZTtWOlUmsb3dE2oRtDZj7sGc9L2+lDx8
nRxgbNtsCCsLqH7SOfNnI7OWFgU5pGPX5PECydx+uZImWXJvrKdMYIbn5E2JdQvR
R8vuuorAnUqNo5GNsjd3m1mE9hdzlJnRTDomQdXL0haaBg7pIQhkCrq1KUpXaHi/
4M4vKL7HP7QGY7OV+9UOTuoM1nYChnGjkDvbzqCi2ew4/fWPJ7BIIbvZHngq+q4Q
p7wDSfEFAZsmpTQWkb3l2O5xiB9KAsZwomwTMvqpAFuxULFd4vbBofw6TLfUtyDp
mSNbAFPa8nweRT8I/3DQXK/MrTYGlnrOuY3m6lvvNOLk9tUAmwh3m1TybC5K37xz
EIo3q1NdiWEHW6aC/JY1Sl8gnMwRQy5aiFxSt8CGZx1HAajCEf/UZ92GbJjxfA+h
lnEbdp6DTX2GcQd4pJNsjyD9x/1sgyC6UQBn964igKtRFjNeY/jHOCr/FxC//ut/
8kvzc8U6v2R5xJIHIsxAZoXZwCLlN2dBVxLd9S+IQ/qvlu/iszeSGG5Q3phaFGKh
rxkjmCiuNf/xxIKnbS+nUDwDTPTb4irwh41wBAdZUagjz4uOoL9WumDCwSJ/9JnZ
s2G6Pql1J/yPUdMdFITRYTR2AWX3ShWr4eVvhK2pxd73Ttcbeirn6t+Au2oAIXbZ
oxf7Jy4pbwtoASCzGSnWntuDSDPrt+7b1UcYRB4PSgtU7nh92YXM0G+DshAJxsQ1
7Evo+EOMuUus221YcRA3zd0HxNzqNWPCu+bjj6bBctDRtbUnGmfsg2XavtCQS5Hs
v+DR0kmHc1TE8GW3MiRRAHOorww/ibXa+ccrWttAtQ/jNgI8w35rUTu1dVhCTDWd
C6ycKufxqcR4rqa2NCYqNkAr/kMAIOBJp2DYpYeH40ndoD5ayg3CeaHXo8We1kkd
OniHUQq3UGnlibakWN3UwhTZpAZR/JTJTFSMd83O+tKtVy6ZhTAG9Zv83OM12FCI
fRO/5NYzUqGbyZ7GMBKM1f3bzgdmnRRI8mOR817mdYD1lmlHjOEzEEU7CAOM+l/5
CXeE26e7WeMX07beghN4YL7b6KPlqWCOJWQlLIPQoFt2h1hRb7lXlHKP1hYfysjJ
rx2naF1pPjwhuAdfQq9MayBbCoejJyy42CYa9RmZ7ZT50oj34i22Wl1Xz4g922zZ
QQs08BS28F6A+r/EYJVIh2mqAORM+PZrWVIf0VCgZfqGS2kXJTfv5fVelvus4Ebs
mxRc75bPyMR73yfR9gjZMcdwslEkvIOkMEBAkVvRAEVBOk9kqMGTYvOSEo38jP+Y
EmcKgKfnHF4DUoFFqvDAIntKn9FkRCo3mfRhdphQcbPxxwaV/SV0D57AMtEiBEgt
eJ782zlA09JusvzIhPcr0D/wBB9fFBOuMKxXAaPILu1EzkIJcIX7LP8ZmALsLNJC
rTfiOzzILAneOk8Cnmofe8fGSrgHBKlAeOk+7O1yUjkl3rAMrbTYEqSspvznDf3l
qb0pDLp+6fvUY/QF15ChlBr3bXk4Jjs8Fb6EwO/Q2zCX9hlwJsh2dm1mutfCuBIK
dD7yljt0yCsyWgjlk3cS9ft/Kixc1Jr8q+exw1hWny/7diMSJe9WKV9Oftxn+r1i
0OMNFKEHdJvR/PcWj1SCH/lZzf91L+CCDSctQPnXRVt428ewy8+4XCFYFmzjZm94
y9tdhDWjE0VfV13TErAhKMemvfkKDdPBPqzSXTGfkYLUBI7PJk5hAUWocXtbkyFN
hNFGlpFfBbwsGEvmsV95s4FG7+Zrb3nqDyNxaMoccPby5bws6A07FvdPG+aHYXPd
mlVrFpP+vyQKvZ/+vNpMP670FDZ2+Q+mjyuVTYXk4gRI879eLa3AFDdxWnKC59Up
L+RUKCS3Q6dffj/OtvvmaXLEKZYLvDF3Y+8Zt6EuTihCTI+wYimxLFJCX/hjFlpx
kNu111imLQRzCumSX/CkU5Z19liQDjiX3oEq3b9LReDyEHqBJshh2yC8S/z2e4Ka
TJgfGNR2nFvlVtbUUby2rR8X5ZfrmqDvQqNd2dr8Me/StsH2vA8saO3zzoEmevkv
hKHs9abUrQBoHfBwyGXOHbGJw7fWEbK5CluyRdaBfz7WNYpG0DfsxF5KsqBFJ9y6
zCUO/KC3lSccOeGNut8rWbvY3vqcB/TI1Ho88qjl+/z1ilfBpoLfux9tzJ5/hM87
gTaMsd9BxyZULbIZluTg71i8EhDCsZTfevYFZJvzVSDIq8lRQqNvg7V6L6VQlT4z
3cccudnaDVCHYUz3bkeYtuFOLzFOHnsDr57gb4sitT5Au7CUCBWooiOsZF4D28mS
PrM0utNEZ04JOLv5w3w8xZ/09fh5L4g75a28NcAUpEkAkHfWTbiaECdWYsnrVG9M
6HEyCj2Wn7KstxzCPIh49cUD4zBLIRjJS0u7asJ6PuKBIzAG1+jlN+KWAqpPK1kc
3ifJpWkTqaPnqG3YNRldFz6vc5NVoZBalzHk0iF51AfzFtZQFoJb5jOKC1pfAe/F
Eso+fwwE9gdczSpBfmWOMQLYwz2UmLjdMxK8na9RRv2L9mm8ezWeXvebVUcBRuoV
ZPdFCOrCVubIAQc7XmKhsMZ1qzyyKLQ1oLZ0CGxqlVhfutTMex/r4ZG0NeekrsSG
By2O32i4GeXMigRfyfc1kG4bajsKQB11E8BlYVoCSXqm943yz2W/A/dlB9NF5d5n
5tOieoxc+/MWOWRn3AJ+T0UDQ1BatX8rhvmnuI2F+A4o+1aIiwK91DAN05GVZul/
PyUBRqPbB+RcxUB38rpQPdSio8P+5JkTZbNY9Aj3MpqM4K0z9y7Lydeug6pyxVET
tBSR2s3jsN1deMcfW5Ot65aUMJYZx1yYCDGLqFautDBrdPGlSWmh8Zj2x1KOV6us
3Magrf8WQ6Lqyb2kWHIodHAGiPJLOnNtgBdK90AnkYKH6rr3jgLzSMNpvEMc1Mrx
wXbryRF6j8qnX92JxMnw+1rhfjuPReAtEoLC7frrdaJ2zFwmqpg743D3hTFZj81l
lyEJ0pGVQdauxwhTBPaqDkr+vc17Qh/P2F/LaW086YqNYVZJJ9MgQycWueN6nl3K
n+Qdg3L6mM3YLGxk68evxZ+EdwwgLdLdiD7Eq8XUu1EE19qKYuv93+emGnZ/6WyE
04m1Lj3Lv06F/FiQ/Ky9NmGmvKHHk01QuZ2Hs4PaFWBUN6F2VlRxqOA9ELQFrbQW
ISQ/+AkXvhXYAkwHRmha1STmPiT6/8Rb+6gyFPLisR2PcPWPTrn7tYebkcHi2ySo
+OBU/AKJZjabZL+nRev0ZC3C2jXNrzMV0M38P6Rt3+A1XWNZj7/s9Vrqm8tAKzn0
KZDQ76edB/MtJdilPePpAfnedc1CkechNT0Z4EttqmBbI3FqT58ciPI21CCKp4qC
nvXl21ljdBDJit44q1WR2GR9vaMbR7Z1l/Vbg7g5NuMYJHCHqz5ZOdnj58rKQQhL
HEqPudyTgaCsTw+EcIKARVUHJctncEU2fLl5os/meZoktZlSCvdSDmJ2WGBvMuKa
BEMgW+z04/teKFh6vxBtQvCGA2ptYhvsPvyz5ORe6OzUmu17RGyIEUBfbfj9vpjb
2Y53js8tRAH22LefYcOCbpKzXj3k9zU06QLDZgE+teHdL/Gvn8YRpCGyxLPhMSJP
ID9f7qCVtoMCfjQdyop3sihFKOGVCOTJNsqvA8R94KxJFXmqWWaeCIAZ/2GHHttb
Bd4CGdx4KwkQ/7Cy6/L34vd3RuGQw02ChnrJxmrqJbLmRkAfIfJh5ydy+VQ/myUW
mmR1J1UxPzWFc0NPwV9nlfHTbYPcbmO6oKywvZW8DCaov98RGTLj0cFMOX8ArsGF
TSZX2OJXbMYiz8P0B2EvPlspmAaz4FDtcgY6eyVwJuMVqBtn70v+GJkThfjwzxll
ObX+dqtNcMrU9RPUVp84Q68At2CaahZpVzcrt5O+ZgNVvCZiTXxF2NLXd0DfX7kP
yHOv/wnpz8kTEI3qSnbxfO6rQgDx4cs8Y1Puej854CZNwCNEVQDYdWCe6pa8SqiG
CkfqXri4XYJfGZH8ckNtrge9+DHfFXJJoMAnFfseegKfm1jlS239RctTh5nEpr2d
qfviLtYIR36aciYkEqZeYwW5wl5lazaU/V6nfOqSrd8Icsa43LZuuMtLiE7OIaSV
+RhuNoM+3WtNOr5gD9OqYxQ9Nq4+qFVvgKsO3c+SMDBqnUK0hUW8TaQyAc5hrddL
3/NefCMQkGgSpKCaIMlqgNFxsqfniapH8thqgW8nyrVvFRZMC/8KBF1jkffO2UGy
0X+20Wx1uOd7lZZSXASbYzZdY9UNFZDvY8hmtcQdACmEIXBr6qSHdNFDCDVD6oui
I0Symzzz5FUmdYUEGkOgf/sfDgkf0GHSSiiALSaFhV8RbUaHIwCDGMnfRCXlDHEO
neQx/FjfXJhCZsve1drdAD9W1W0c6X95iCy8AB91MXiHi7S3qY+hbfUV2y1rxnbk
D4Pohahf/ZyNKOXJS+MGo0oJs26OI7tScHTmTCbTWNYFC7y9ggVcck61emPCPXUk
ppfQY0WUinUq8pPZ39DGL/SMy/PzpsE4/736Zvww3IQUKffsmtr6PEYfu3ADx7hi
Sz8FDgXqJZf1P0+0L/ODIOqsqOlOM5RxxQ+QW81/kC+G+mmYnZFovc31Z3+mu91O
qQ/FX24JAFcU8PPREt0623oBs2kYSy6vVC7ZXcvsi9GQrqXLZqCS1WrzvceTr3vP
mATxjMfeH/raRO6QyTBzOHQ8/Wm5f3pwQIvcL2PLQm9LhB0EvpvXnF6P13X6YX0q
468cGEBkKSbiC/71619h4LW/vSbrUiCobMGNM98oi7RKvu2G3z1ktWrsL9CCFVW4
I1zNeLVkCswAM3uTP+ixNK2Zqv7Fx9Lk+KKzI039aaTyU7tZAx6m6Fp7MRUMVO2N
qIyKcWYXV69GauSLeKmE3xvYFwN/GBDwLHS6YG6ges45E2zgY6eboeogpwd2uY9o
DRF8XONC5WBGcATlmiwNpcOWBDv4hYINx/aCEShSYYjNhFsCRLfZe8MEO8ARjS20
CG+/AwcIf/Bp0ACbWh5BVtSSwoLALI0eQeG9WQgs6J4Ct2bDtgdy+sQUQa1reqEh
raZTuUEgqHD3GIL8gb4Yg8LYvc1O/vHdzL7C4Cez1GsSVKSmRIO4Uo6TTHWR7mtM
+suR18wbYdZPErYfiQqPK9SZRnDEjMJmV6scSVVrOqUx7OiaM+AIkBeoUP8793zk
AxavBMLKGkMHqN0fjbs6J1WcXTfnwNRdBYYHOxl0mjX+O+XBGuauLAQeK3yDV9mk
C0XH/sbNVtN0QyeFUw3B712S8ukN/fbfzCjyadxZWm7XcOoYokzSoV7GQ2kHCQg5
bXDlwrCh/dV3XrhbzVCH4508nFDUd0rTndknTt39cNhQFn846pIU8Owef4amRMg1
9WoyxOSD8D1583R4VQ1T8Q994FoPJfkIzq95kS7MeP0+Jplbpu9ktK4PjXrG7mrH
ZjewsZcpv0s4ZFuyI0TyaK0TPQhIPDaD3bA9717vwvTARtm0+Toera2Q+1Dm9yP+
H6i0X1rmu+M3S03d9LjVqFetSpxrdLbjamxBh4qgiDD2jhsNYgsDCU35iETHkVPy
ihyvKYI6yMvWaTMwkFp9oOxQcHCnOV4bbCKqjND1CTi5e5wlhqBKXR5hYuHUt0pQ
KOVBZtYNUWN8cZRymENTcgL9oGED0gQJp+AfKeoe+WPwnpKsqaPdsiXxiPDCHwSr
u076qFtRnQ5wHi6iuGhpb9/e4T+RAY+gM2oyh3SW/TFiAwmkwDBkh0dVfr5hcfIb
M/X3Ap/rhweiBqwGr6L+BZbgRbK9h3+udRe0bS3rvbAT0rX5Fg0XKWS5/vagYfhF
8PbKlQtpXXqAUlBsHCWObhKN03sfRGJTqTkdb2VWd4g7LxYNp2DAwDHxfUYLPoe3
5wkY20bIJQ4moqib+IwIO+HK0xd4OEa4agp7oB36cxIrdU7SdPovlUWdYeapvFXX
7DySSrZQ59iVAnDv5SSF+OaJowEhS4BnTzEkY69Jx8PSf4ZzU0IcqjaUQcNL/Q0S
ERY0SEq80OgsMmEXuKqjaTXGLg5GDDOphqR1ckmseMEsHhwy2pvpjk3LAqs1AP+x
xHeogaCGKYnQOVtDkNHq58R1Bqz+F+xMIrkm7dlHxik1mn3Gc2ANigCHZkK6/soi
UxSzqSx9/K00uF23uH8yhY6QDFdzgFIwUzpk0l+3cw+r9rGWtVmhN9rE4sJuotjU
msW7CS26x/g7bWbhpDbHa/GsSc3YiSRr0NF8qEuRLTYIR3l6j7yiTKy540tD7fOe
S5Q2CpG96QoyofLQTcGMK9Dc2h3gLOGcCR/KlapFCA0LKrzGMWgWYGTv5eQb8HIn
w7LvmuNBO9ANad4RD95lTFrXUfat5CKEPunw6lctb/wB0NSlX1cPEBAaP8IB/BRb
gkwW6b7KEeBQsbigvtQJ03mLkH5tnEtqjghB3TYGJs8PQYUFfs+Dq7QmqyiJQPrP
mA39CDnyBlnf3x/DbhlHU045Q+RyehE1w6Iav7b7jJWtLufLD792C1yBezj/gqqR
azw2LMtCfe5YF6qglKIR1SAW476L/dA9NDIxmQMjhTcKnFjGpvJSx4Un/OwFnZ7B
FXnmls59oU3PPETmkcl10fPq6+NI7+/4ZcyvAZpAiItmPIkGrSM4F9M06C912zoQ
ZKuPAOKj6d2bTlypgDGM9GHJ3dVAh+OU3xCdmRkLVMUfoLmWBRPoSDQX3ANBZisB
QTDqkV9fdaRZUlYB5iERZ7pJUuFGe1RghDrLrUW6MzdOcB7j5uIfXXUGBhDDAMJ3
35koZ5y8lc3etsv7DJzjGXCfDzhY9GSsuJEFGD6K/vPOVKK2OrVb+tD+7c2BLIMP
Q0lFdoIyyKKtYDW8iSKIVh/23tm39e4KgOYwoLgyHxjwqZ2x/m/9h31uZOhAvvn8
bqq7EKgTR7Xv2gQQyJPtIxSBV6qSnjWpD2HxUY+XGw+xRYJ+l4D7mex0wbaHLQnc
vJ7rI8kzJDun0+iSGWXt30Khh2fUR/eo96fF6FVMaA88npu4lGjLQomjiLvjALL5
ggrwak2txB9Wq0oMYXslINNtw/vUh0IBtdO8L5xio8UBReJn5aOsVy/zhvDtBTdH
hJckhVhp/N4d6zZWxNTmg413JAgZudvFeDpvQ28BylQlmbYNZxQwRmno8NxBNV5m
/esvTH388Q43a+QtgnOieuketpOSWst29bH80Z9L5hcqXdFS6sEJkhHw0+OHzVwh
5MiBeGPuEeVTbQhXAGR1dTeyzBzJkvxFBuY0zd+JAUPr9HWBHohMuYQ2ECBNRiz9
aZcZTye1O/BD6wYIgF9e3MfyVNPm+Uo7DHMYbHKOgBSuHjd3WupdyTsN0uhsPnvO
mP314iuOBAz/08e+TiiYlE10hEG3EyfVEA6gM1142LNggqBVgmOHDjq6Ltti/uWL
uM2TjRT88a1KoD0JX6+APPgh86B2fqNsqcM57X26zO0xavhDqWKCt8+tPY7oYPrw
ko6pRyqXsc//y+z/C5NhyLGxkLlX2NE+iu1d2AV5g0C/Gh20qB78cOEwCqka86aB
mxZw26NFRatqvVJ7oFb22cwh5AZiCu5Jie/bXyKLX8qB4xikdRZ+0GAP2VU/UwDA
2pspvwg+9vZo4e67+Wjm0SSp8cYnUCxcSN4VKSwxAelVUYOX96nCzDvRGj8XLKZr
Iwvev/BvcbVfgK6mZzcJidydJzSD299MSuq+d5m1TcNAkw5aIHEx9FBghUNHeUYQ
bbdWR4FReNwjTQuzPg2ZzxHr0zNMTXx5HdlGicQu/AGBoTNQ0xgHPpugec5knT6P
/eOkHQRiAlrn1y3gqEHm5wRGzqRS7n7c62mLHZV6JPyLB72ANRaFXuMpYGdoC80M
mLpcEeI0wnNvVh/OpZhzH2AQW+Q68MnnIIpPlFOjRxz1MSJdd5FX/+xeYE1jI1/L
/QMD187UOUhJd0PKg02fclWEWGgPlEDAPa28YVFRdHwWtas00LsYFGGGPW7Svwr/
2zgKKU/p8YUqTnrsLOzXHOI2tKP9gVo6bstKjIcWSjViOEA7qtam/HOLhYGsEwPB
4ehY0sX0kpO+1B4WSNezWc9drvUa/j7JIMMfTnPRQx+Xo8mfVwsU06iuJ+CCOIPU
XyWQU1NOZhMO91LauQkzzh68fS+ZAQ5ywH5yzerd2aOI4+lLFVn6icUMjpdeRtOJ
7pqtld7kONIDJrOxypj/Iti5jttiRfDLER3BxQa6P6pHpQjuMeH5ndXwB+1I6rGZ
iZVYDS7Ecl0Li8QJvyYeP1OEh0SS6uVvYqvAr7g1L1r+/09cYUNarMtFUuVpMSEX
dAqTjf+VDF70s8kQwhbnYM5goW8oruWL4x4T4ArJocEtAZVutbiu0JRRtQCfeEWF
alKycEcE4dkEK3j59klk5CTiExDAbuuB2c16tf5Ok/H5gljwegyhGXM403VJlRnC
WIaA5tSB1T0W7pau6I4RSTVhIek7w0Azn1FZK0CNCxQEU1WkaO+CT5GV1jJSsBTj
4qR4DICfmI0RG/s1fIJj+SutC9aDWpxERMyoBZIlwmArqg2YBmq4r4N7LisophDr
Al8SEs1HC1xzkaJfLiQoT+qNsCNX3UNs5ZMzvj0uRff7UAk6obNHVEvgQD/3dRPA
jowv3UQUJlwEedw8Ux4vxrZdAlqpy/r19NVDB0n/r+8oKFcmXlwb5bEOCQYzvGlm
JI+PL7TWFvfrhD/WrwrP7Vk/EtoVeNtZX3DxG8Rjy3iJGK8dkEpXviHof84N+yB0
cHmTIyOg1SVXj+rIy0LxKitjhWXOgfqd6dXUQjMS4oKfyiP14JH7il5Pv/CSD90n
Mf5IGjyVFNJ5EjIPWu9m3g17bmVttohvv0hhbRTsrEbjzG5VTEOh6lRJdDU9U9pv
NGofqllTGsRKxCpxW1xHhF2MoseUHBk/vGWHorc+cRlA0OHyarN6EH0/n9l+WQzS
6ikrHYWkHfiU5Rqd12vlb0BFvAg8QB1XzoeiFR6TUgAf8MRTvuPiqDrUTW2ocWyx
0UFn/C2ZaLCNX2rAL0rbvC0IP0ZB53V+KKuqJVjUNLKZekceyttoahcgkm+rKq3H
TWTA95afebpDrbMTQo8IqCrzQMWPZby8GX72NccCKKEhc43EkZmB6dV+MaoQh0oK
AnPYPmhd03qj0atG3ZPoBSqzOSJS8rXf/0KMHJ34Ccc16PE3/OsqL3d0+svrS2p9
UyYGKJfWVeP3lQAD4tKtUFeJc05fuXIoeIcz5CV9R9nzCktvjm0LK14FASD3mWrQ
t/e+mMIp3Fef/6dEM8AYillVHipshJO1idSsDtvZZWIxmVlqjewFMoGaoV+5elkK
O/QXeaAEiOFLpTQNP+1BjRPOdBlaq1cJUkcSYOxTw77jE00B8ULRmmoi70fiNx8R
LjaDkxuNX390N8KChWln4DTMzNYzrF3WZ8N+bLo2evs/zQAfjBPo9SA3S7UER6VN
W8VWIXRgUp1qFEwixivxF/TCKs/xZo05gEtuiacX1LyLJoeq11WRZxnOdyxQ4uCM
3tIWi2taMr1fAXReDUqW6t8acEPc2iA5XnMMH8CEF36nd4FXfNfla2pagp76DqBm
jI/Yd1yGsT+3vgYEdzYssw40uBTGV5x5G0dpkLbtHjSctDCSc3zfITKpR+yam9a0
hbpl4oxpoCPOP3zebnVjlz/ilBUglVt+dBVP3d6v3wI80Cc9LtNt0K3TXXH4/ss1
nkGd79H53IQbw1l22bnXR5xmrG06YNRmL9zUY2YRHX2toEz+urm16ZtB9h6LSBGn
5CMGMKie7swv5ZuXktV0L5ZgJ7eVaxKAR+3RW/0fkAs8DsYSdOqT7+zFmULa+iPn
RRUVXAwoNsymrFBMfgAF5LtINz6KEYcTTiWLUGxnSKEPrx0YYWhhWFBHQMTxQ2KA
MZrBQ3tteN4svLxEf7rd2hAufvvxWfsv31OlHSwyxahixwPAJF9QBF/26z7H1yjH
xgiQx+Ycldm62ffAv3lUUlXHSucL82k11w/cOrzXyCx8mmSKpPZ2pEcK9WFvwUDu
9cYh3DiPZ6Co/uUQDEYmN4cq445ynJrnkPUORmSdiWl7gu7ll3yShYxuqGFjlUCd
M7mhWrdGi8zlUIpWUro8Jj5W00K3kkbERa7H8zyzsGFAZ4WWkvSdZCkCluzKCMfp
+bYG8bbspDSp/ibxIF392nVchAMCXVUPkGjTEnVcG7bznn3nlAlnITZOhkkujPST
/y/iH6jCmCkioboHI48W/SpqnwSRlhXTvu9A1RDWgfSgr8zsa4Lhb19GXcYOEOXM
z05q5YJkS2P6Y+QNPUdWODsNIdPImdMIiPflFRaG73+lnETNAkBrO5UFuU71idh3
KR6n9ogVwMq395cywYoprApABOw3AoywX5bS4P29Dz2FlbLzrK464XwW/uXwgL5o
iUiFJNa/DAdu6MeqyK+/l5HT4MswsCGeQR4s95NiN5yGnKFdFELYf+E+nil+EKlo
1zbaLOL99PDeacLc9qT4/sA7bbIqhNd9dKCbb3VHTc7xdam7o3IUjx/sI4zN6/n2
NSskhehjTeshBCjm10/lFS/DPvBXLnTl2Jq0l5cMy79EjTZ5bnuNe3UJ0Zoxwv8y
DQX00u52aHVKQixCQzsR+y6ZK+GryHki9HKOjwSrvI3ruIOWzJ4u2RZ0MfyefaA1
i7b4SYvEjv3gvxCKqqi/Yti96kzpQIFtuIPvSXQBNm2uafqasmMkvShBKcnu7lzy
PTo73Eb2jTxdI3IzRFMBNfA2YCxqTHm8vfCXv6DFBjfmJ/L+N0KHbwLm9DHaIzkp
U0DPvmcvmLkw0mLT7mYau7kaIvFo00TAYV1lN6Hetdp+apHeSGkvJq6//6JgyO3J
u6J/7IcLaXbaYpUE9LxbOUEPXc9AVbgRE+8Jr+DqW3dM4esQJeGua5QykFf+eDnR
kXeY3+6lL6XUssho2da6B4tb64AfSOxvH4cAOIQjfT8WeaAnzIooBQDsGyYBsu0i
YAjaGxj+UyU1HX8gMt4zjfWzGAIMX195+tDsj7H/A5ZRU8QkS9gunF1D5QhD4zr7
TCbVwwULQQUlCTvAASzpj3+7Go8VcL7P2sibTSqEJDv9at9TVdICm3V5FxVM7m6E
SOg98IcFPMgXZvq+ibdvm+1cdxnJ/I9WHBLnQcbF1zBptTBIVQPPEG+EnoUbXoLV
W1/uO9GEz+JUgZ293Ay+tj/E9vLxUawzymzhKg9i1eb0kMKAWdJc4BWPgWzLTRCx
a6kwLq/xAfHbU2PFi/qLfPch4b4kWwCycf8obqC+1N4bZys2DOwAn8eXeEAVWiDR
bwPg4Hu1Nm6nLy14CZa8OyIggLYabwdNd1zMS6Ty7elpz6dpCVfcYsY3CKWKqPGD
gOiDOtA0FQFcSBa155hhgdYNRdX8EFCOQ5qkSXsorXfTo4jKUGhA1+oTEuqUo3ZN
l+Ll62OMCfS3NOhV/l2Q6zQIqzAM/aqo+rq1m3TYem3FZoqps6F4cIIzxzzbo3E1
GseAAC8NIN5ar++51Q0af8J5Oq1XDjiDIAzQF5/4ENP4AIoV0WzGolGQHEhPmSBm
rbcmCXu1wZfe8rilUXbr0VxVoydEQtO2BBbtcTKXEqlnzDMk5RePc5g666BRKei0
f0wOW46FeJjc1Dvvtc1JDeSoy+/4LWxcsAcphEuKLl81gQ2Tyq6bP10oNTEtBkf5
9Tow5E1z+6RjsglTPGF/oRVWHU0a4CwFGMIJ1YVFn/pZTo1mgjb95hvZZwyyJ8f8
vr5wGsKZ7AZ8bh688B3V/nsWrTs4SGbCHiYGnzcGn6W4+AM3o4Yc0mOFJtKmB+3c
An7OCvjAzfztvtSH8Rd5caUHeko9ZJSJJesYeDbvrK0Di93k3UNKEraLuoZ8gaX3
XnTrtqBa+/wLMdzREerS8cXwZjoo24fCl2pNpKHUGpkGkaZKCq15tTAkkq2kY8t1
ZhirtrsQlz6UCpry5rQR2inixpKfJCOgxpHUzyqv8tiI5hzeLGxnehEa0dO5Yyw/
TJTDr+zsKLrIN45WUQfIozFqkqfoim9CinBJTaEfir4H1KijdM3H/71mQ157+/XT
jlqCJ0nB0Gj/4a2hjOsm6RaVnmDwdzR+4Qpd1z1SS6/0S9o4rQW48Mwzu9JlJO1I
Bbd/sDEKl1EfqCgUmnQyTzaNdLRDI6o4mPHYs1XBCzI88WOoEEac2YZVSFLkqylW
SVf4X1jts3feMaWOet1MmcCTXRRVc/9KYl5jaDTNvlFdANpwGUcEZz9dIMznA4Oq
yB3aoyFyEjYQj0yBCJkdZ+FOyktD/bcM4NpjlkiPbbtl5WYoyygGJDV0+JcgwzpV
MTuKKRTCmcO1heF13ojIeg6CZzB01v3G5xPjKfK1DbgA0t6oFS8RnsZHTFKjrVVU
7pwU775N12ejHNdi6Yc35nQbdn/REz3nuTcRhTPR8GmxZxzBMupLWmkfJrz+k+7i
bdKrUt/g945c1284x/JW6ugIeNaMt9g59PASRIoQRPMTnIRW7ILhy0/RYIIfRH3e
/gLtNF8rz6dwVYTWgvCctA1cn9/NvRtYEEZIceL8muVAnRqUmMvdEWMw4Nawmszx
DKwwgjTZJaA45nBBspSaGEooQbLyWsPCFzIltYumW7T5XkP/bYNNis+5c4o62KvR
mXwILOddXWAJZm/SICjFibwYxRDoWiDSBf/aF5zHtRB7p3Nu06pphbda/hKWEZ3u
YGGBLl+2bXPJd+zRVVzk/O2J54hglbK6r7llHX7X6+Hlsr+fFQdxeY8EuicwxQhF
SE6RbjDhNJusgJgXlYeLdQebKdT3Gy7pA/bRhRz1EyrsNFqeb3SH+Lp/yeTyzU3L
idS3TUPPsRTZ67E75W32VT1mOFtJy3ElR5E4BP80644Ei293hxvJNb9dno1Q6wxW
1JzSMrzfcMiMeIfY2TLS8FkT4wXARs/7G5mg9/0vUsO8Pxgo8fQieR9mjAcgvuoQ
UYauIOBgj5iu14WEVRAfqhs8KfPvSRE8VMfM6PEpGjdMEZm4jnx4eA2LMxg+BmD7
Pw1bRja4+Wi2n02W1p0TPCRkWbgy87K+OrjjCmIrt5hgTsCoRwyiPv5PhBsQ5yOl
2KypoHhJLtiCBSTg7VeUF1PzRLzA+mIGRSTupJv0StznPlWVjjfTDU2DxmeACHZK
IPz19Zmsv9X8Tm2IkrMRjMeYQ9qI3lvmbFNoMZILOlyCu/+YVj6YR7IBxZZBfFIj
UAg2K7NENbm1IbsPSAksng7UapKwlBQW3alv/HGaHloFQYcebbj3z0R8f5kSxhll
ECAWPOuSFrqG1vviF64DgrMNGewkxovhvVhTaDeKdUljgBp0CoWK1JUOJmEuSMVu
MaF41PiP9+bxgpT8GQYNWP+2moK5LeU7+ORiHgx7TYmH0jyLnzFsU0YcMWO9MS+a
WSGJ5Bo7XiVcnzmAXgQU3PyemHx49hdlYrFYI7Lvw+TuaDOG+4QY3Lo+rhmKjs0h
9F/gO5VrIhZWk/SEZ66CnfpqOfVenF938y9D87vS8cS661T5S+p9XwcaSnPnev/1
2hVEl/Ks9gedZoOxahBVhev08zuZsJlQj/kNAfWVNe2KvidQEbnjMojGQQjrTHoI
9QZzxsPvep2+77jrj6xnc1i58DtLhUa/GWa+rnhmxWDiA9p8LiKEObmAc83sNt8Y
ZvZ9Z7LReukwaGIa6zU5XGKzB2mzeYmUHqPK+PXz5rKLYgezPfhg1xUT/0cahgLQ
9wZejJQ8UM60dZwHLIMoNiMQjR8ag5160jeDUDQ2XjoFZDFyCoXx4aryUfbRmWG+
5BBkdZKPdRgqPe9WE2m5g9QhSyRO5qzM/BMGXzp+1XeukI5Naoqa6+rGqTMy/lTE
5C1AFLl23G7/DEl+YmvXcVnAUlEV5+FO+6x5Bmtw5D8bJFcpptSGMjx/bVyr7XJt
fI/ZrlTsC3w9zlCGhLd+TYGpDZWJf/gSzWFSv+iXGDMOU2+MrGrngx2PjNiy90tO
abbYr8UQvKhpiZHP6noSKQIAezdBbpxRjSJCY7upHV0u8/wPGBiC3GZeOGWeCDme
AM8vQ7jLxfiYaK8OuXKK4noKycZOIDPPeQRfjUYrO8ikjyRuJsSQxQgQZuAkPMY5
Fu29QGnDm0luJ9YuL3Lq6wvcJBBzLuP2r3Bj1/aL4BegnQY4zr7la2MYc7Qvmwe+
heazpjlXgOdNQ4Njk2eXRjz5hyns/NWtAJb3avuJGbUA/RBDJkRrt4krW9PiF9qf
pd/Ji/y28vsNoUFG28zUmg3Sr17YhRsxK7RSseUmbM3/cWXGi5Rcx6cbvEZ+Eq/2
7LW9G6WyXp+auI8aMSjEkhRGER82s5vPhsPn8pYU6iqsFPhoaF2DYero3h3QrX2y
2erelT6l80EkIkwCuhKGh8tXpE40ZGQ8s5JOLjMFYk5gaCz6rCGTJvU48QvJahrF
20sQYlm/mHOdmFrUIVmgBTW9rUILyuPB7bYiNXj7yPv5QKRksinclOplTDk83U0h
/PjPjBhe5f1AvhdLOCRk66zSo1ebQJPvjwQZeDVXZ5XzIwzH9qSTJH9mud9uSlj1
6WxpF3Na4vminyC0sIeyKYGejM5wLTYnXaGXSbobb96xzH+ohXjobzFXgIgobnTU
Xh2FvsLmyg+ln/qgrV402aJKqa/81qnScJsggCSmMDyiHSqHfKfSrX/99XAKM9Ay
HA1Z6s1Ht2O2/VwczLI6ytIizPjLMaf0nHY7mwl32VtIARDR02NOSvH7X0Hdvxp+
g1XwFZ3x6yibbhfQSesLphF0ceA95b6uH/vJVmABub2AMc7mtl4So49yveEba5df
BT7RtGNzZuVfnpl55xiQ28VPQR+TNFCrbixHhqz1U1D5rsPNmkRSfl154Weuovzc
ddtJVxpX6Tt5AGVsqT+whJnzlaKSPiQe4Kc2WYytxsQ9pBrrFyA9G571iWyajzyi
P9F5f8AupCCCIsqbhd5aynRBZdw7Epb/LkxBuxdlV+Eurpb0o8HuNXXJnGOJmYTq
JQr94X3nJAPRd2zOlz+0zMCVzReTcfmvkmrams9uo8B+tcSSMnfzQ0qv0ekozB9o
iuS/jKZebDFrSEJsUgUmWMi4VWe/qAF/zhJOx0xHYMtXgBDFj/W9/f1m42l9JDtx
kGzK61Rc2G7PYFMVhM5QD2YFpRHJoRQnpb3wntgOvefc/FCOSljRwkXS+dKL2XSR
B+QNGV1krABm88jZar9r5afGEHgeXcz+s5zpHl7MN5aUx3+xbtGoIxCRXbk5pfuR
n/3c7Q05zZ8RQzg9BA+Qj+6jUmOHeJS4eXq12DteC6bq8b7rqms3JBwvWVnGszrw
Jnl7bU/0emm43qfmDK+OzRS2mMf6/XGjIklBrpPyc3bKqs9FSL/pQRPjoifd4KHp
TjZN2j8giZYuRJa6ROQFx2TQgTyGeaXvnrU9hFxLpPEtYtqHNP+bvigvEyYXKRM2
2lx8wdbEqtbdJL6gzzh1IGmjjnwxVbRvopmpG9VhoKL/YcwX4O3Hvo1sey8GVijI
IvuVVSibBmp+a4PbbNnBK7sAGqs2Pg3us/lG+UXIOmk224+6gQtFqbk2tOiBCL0w
b7vEByO3dpCEzYi/ZT3pRIdC8ajPQMs8Xjjkw5EdCWriCNBFQY2tRQnfNaFiW0ra
0+62Nv8L3Q3lKXtXvVXdQanf009pRFqA7shf/bqTFVYODk7WHyGfIu4juNovK2D3
sCYYhvWm34TAt1wWaxrKdpnJUWnXacxE+x/xbs2JmPbH66tTwwOST/xVJvWK2471
CgJ3rEq8bOJXhsD9OjMlRQ2lPiAYqoIFhtsAE2eNo/nEmYJPpvZ1YV/bWzcvxre8
fOa+1Z14/XKMSjBUzTYlzLa2/ApyTcS5pRMNz+h2+vcHUYMqGOCjb5FwfkIo6DHz
T0x0oV4Tnkba4l0e8GeW2jrxMvtwwrUlm8AyJlgWqCT+kzLSVQbxSxX0AP9DuK5/
k6WaaoL0uZuIsVkrTec3u3yk3Olni9YjjR4tM3AKDgHODbu4lTGVY9wtGViZpXzL
ONmc5VgO7O/U96g86neGEW/hTKC2IuBhpkrNTcqzDp6C85kCyUIkzP9+0QpNYyh3
scszOK+Y/su6kCO9pnR5AXcHsDf56EMWqQX1a2DFGp6mMknivxlNQIU2P3n8zAnS
+d78tJjA7ijtB2isOG5mcLZe3pJpLQb1fKMKSp1WGp2DnGYxcPQb3bl4qRNKGjAn
D0bk+4vPzMe2FpUAm1trJ7oifMV3Ww1r+NHH2VUq1C4aTdZfFIT55pBEGN16t1S4
9whBIL4vaKe1r7ep+rUzEmCDC6zOAY/TIbsYY79NflU9EIpvRFqghMEN/Ed+wSeW
QJH7n7gHm3+uyiA5EPzGfy3GXv0Wa3vNdJbKSwLYEt5+tMGVCot+ol/JV5A+Tl04
PWTz0Jgyj7wzKaorAx5QUSn8Jas/mIcOA6xxzz2z/fjR44SXON4opjeDNhjWat3C
XuIhjrki+rGXax86xRWUtpEtJw97CkyIFcLy57BdbBWRwj667rBJBZswVo6qFsBS
rmTxFIiDKu6sarp4cVQiby2lu1tooQRUO/8DnfnoUPRqpd+lyzmLrLQzpiSoYme8
AnF4tHqcvbTqJhtonIFo6f03h+/RVd2xzN8u66aFnx67o3pNAzpdOqc/ovm5yBLA
iKS/yqJM+vQb5NZvE55FAlegbXmos2RbNqkIHxyF19Vo6zWtNVoaOdzDne0BsNC+
UOxTZMrJqd+mMIdPzoaxHw5M8a+THqtCafQVPRb8yKe+fCSGF+iybvvyqSBc4j5q
rd2UxwrgqvdfSKL7LI+6xooFkZYXn9E7q5y6qeXEIjs3GrCRprisGcuZOmvj9tjM
VMtunca6RtAeSdA3S9cnS+oCMutRuGJbRl5SiDIMaDWycw/mKZwyX7CNj/8xwSTf
+R0W1zXcO3qQrNmLxZoVEX2G110zt1X+oULyf91lGWfxr03DQo2P11D4xkFPRMID
XhEN6lDkSHXJubptiGMtvwoBRSaiReNWEblYaM4ua0unzB91pTZ11GaAr6IzGNbX
U6DV52CbDf+Xj3XTMUP6b6GbUPgNMdR1MgxK51WkYFQLRcYPdbsOc79j8trOpy6O
qQoOvW9Ai+7JZmgmaGRmFUyb7OSb0VLR4hAi12/Gg71oFAAeK/ADnPFfbABIQKBB
389fhGe+unneJ8+ZtA5WWNuL5+SJkNtfr7YSCI9CQMB1VGIeS6tAaNOAl1llsKuj
cKDdcqVrlApb4FA4FSDP6HfSD/u5iBLzF0CmYwbnNJA/X+MDbQYOu5vJ3zRYE28o
XTKSCserHLC55fNyRJUebMwU0OLZmvpZmsq8BxzMpIsP/XDaZKnwJ/eo+TYZg/JE
hJtKJLgzFSuUqK1zr8m3CC6KLAn5gYwDPRQJ3a0ZGYjbkjwoG3Py5qTb9QVI7dOP
FZ8I6s8PE13tm6R1KpPRTHtv7yaUoRog1FaWeptkRpHk7RynUEvUKzUb2bSsz/zz
FeuiFOCKJq4A+Hsd5o89DoedR5dM6FPNfSVJkp8u6s4xCHbx8b+HbXrIqHknSEtV
rVRf0nTOJbrsS9PPB1jCMyLbCnCS/5BaOStYOnoc0G4VWaCzu+kcuxsEB3McGqep
kKunoISGzVgJw7LF0v3iPsr2vZ02dRdGE9ZVPer9zDSwgUnMuaGfWvubzFrn+Gow
ms+5+uSXrijJ/a032j7E3rLbJIPqWSfJXVIenkXIZpLLuGYuSqLLZhxO6POTz0pH
mtRV6KwfL4iE4d68Gx8pskoeciebqVgsWd/khiQDbrLpsgdzRJWGKrT+lYsqsXqr
cbMdoJnDTP3brP2fv2nuRKnwQXdqZ7RWGuTmIGypGBEmmc5TphUMlcZX9845H6j3
HdyjOuM75lF6WlQ9Ui5ebcaHaUCGsxS6PT+UH+pyW51Y5CZs1pSdECktBqG+U3MX
zRMfDmbmxbgqhhoOusSCRCr7rWNvAZ625Gb8evB125duga0mNtsQlJgjiH0CcKtL
kruhy9I26HuNjVBolgmqwMLIKKwsILAVsfNl5DfN5HWBlhxzfJKh6ooe+AiuGp6r
E/do408dk+q6azVfeXhh2o5YdZ0Vi8Ah7AvsyZrl3xQobPAGCzrUMpksLpMDJYki
+bUoePl6XgKiMVIbwiIbG6S2BGF+JVD4BVekm07vH3bS9vipNERkKzfVOe1UMeif
U7HerUPc4bh6SR+6NWRQTioHClpKgHObePBlYrnPXQjZ9mHAyqIwk3Y8Fekfag3g
K9dJ6qUziyLdn3FI3ICH7SOw2Vq7BZNBWHvbxlRWDlZI3c8YOod2qTrO3TKiu1dZ
7CXsqkGPQP/aLb39BTFMoEqzAqbogEXVtNgu1Bj55nTP+589td8r6Zav6IiyI/Lp
ob5mklfiNAYL2HGX5s95t7HsvuWhf4WEyXvRrhkkd68DcmW/LB+BjKrETP4TT1Um
jWyeARYehYx6r/6xoL+dS0vS81j4EmFV82QLKhzD3fxYBIXmhVkVVYkhoNbcp8za
Rs9ViRuZFD8AwBI1umTEzRyn8d/dqvm/G8NsgCmMnJGkCF40QTmkljePuvteqaO3
HJ6LNkWIXKrpWJq2S2OD3dOQOlIi922fESebZajN9PYAa/gNcMTEJmXVvQ1U5phD
91IAZcUtXN1KcEhVkkEug8AbfWlG82XQD3e7tf8zYWYs+LqlBvduW2hxxgFcxjTb
raX4axceQikWodLdFzgY28+/uB3bG/SR7L2an0gSeTVsXnEIB4zFY2OraKFkpjuf
JlcfW8URKSean475G1FckidzzbAp09DrSy2bCafO2+2DgQQEEU+x+Oz7+cymh6cs
DlzsBJpqvcisOZ3/1VpJ3i9J1980dEMOj6AZR7Q+8XUOM80MpeKG9RuZE3DgMKHB
BClQr10bBOYJ1aaY4TEUmbjollCzPRLhvoif3tuw7yyPuyPeSph/MdDm4n0bl6w9
AkbhjD73HSaI/u1TvAJ0EGPGmRfml0IwgIX0FleqfOjfx91ZqMXk9KBLr3H99eWK
1G93eZqEwq+q5UsofKgsTHvHMnwAGGNBgx32b6CkPhxAOj8MqKy5yGpCvsPRUS2Z
wGWc9WswHnl/9On1tVq4njbvEHsPKROP6U0dXqxY3HjGsOSyEBrIKSN/7Ph9qm7G
Y2FnQIjYsFENNQhL23SVW1HdO/xpEjrri4WS7LKyDH69/BOtQqgAabVmEDMFSEdd
tf+2bYH2XcGZBbEQdF7cWH/iHozYzq28+peeusJKdIiUwlhvLBHhsQDTmwaW1ITI
LoQ4jkkxER1bmvv2KZ+dGdYNMajOtc1p3J1XpbrPWJcEu63WGUlVJ5WxXkGNJHxC
meTp6qDeOMC/9BnqLbIHylYzFxTucLsfzGfcWzxjn/psf/LI7TR4D0sea5hEcmfw
QM5zDSqNqSMo665wTVSZAxusytDUqgQ5T1HVfnLy2xZSb7QS/+x+zbX45lPL3q8H
81e+dcd4UxWVd3gbUQjwksO+7fn4dcFe//33aXZubDWgW0f4IpWhIs9zPDyovbjh
Yl3CY74pSJmE8L7okfTADCb69kvcxmVyrEw5IzXoTddO1K+6vNfh95mFHyDldeCR
iZPZbvoSSwxxpbhbfJlW71W4/aZRxdesZXtOKvVxFXwbYlxzcvIRay6c1H+46DtO
wMqtC+PVFUFckh+YZt3Gg0qEkwktA5g2srs4M6Gi2rAgRem1Y4bUVmD2shp1cnxR
C/ZRqjLd6W+MlGgcUgHH9W09YfE9z4vTqy0Pe7j7Vr85YR4j570om3ufU4IE1oil
nT5S00GVAYAsmK5zq/vmc06wSQvL8K+UebfN0NH1R9W54qNrf69TmkZjBtP0EHKk
bqen/jExd/1EgLIW9+gZiHaJbpOMdYAHU7CW39TMd9E4HIHpuHfmWC5nEIAD0d9p
ij7Qor5kcGI0afyjLAq2KOAB1CRjwCGRhofv/5PZQfGKSc2pO/NgqxYPWU/jQnJJ
FiqFqn+rSMABmPiG2MJHoPmfBACHpzPdoVdaGFmJ3KmFT80n+dAxj6wyzb0h2Yq/
FMuobrY4DvyWtxXv96sCorK/m3WTmg3M09zY+EIt7SqZPbs7tfkd28wi3nUQy//o
TRlugVWxGGoQpn272DyrAydAvcisvFjXmWpvjqLYKG2lXX41cdCKEdq3fDs6cm3P
Cu3w/UejqaMdx/3JLdKALv51jzbWrqH+NIC/JLJmNXWrggbmOsDFBBvBWPlVsY2n
uxKg1Jv+4SR4DVg6Oj2MN+GYsx6gYjfPEu6ffSXDX9fT1sIuj3I2VGH33MVPuNY2
LMoOHCOaoAtGfxCj2y8IfrTz2AojfWnTjFbm4rd6N+Rhz+ZhxFumZXo5S8KyfhbA
yOWyvNpza4frocGTZkD93M006TlL7ruWDyVMaUAwYP6FlOPg2nuRa0RLSNOnxYs5
47URzfr5l3a5yTOW8L+OaQWwfYUjgpde1LExRti7A34/61MCOJCSeC6y6VG9ELR9
PrMEChBfpPZQTGIcfEAmSb6QLWzQu+u1R1gE0muWdiuO5ptr9/IMxpI15OvVrjaa
UXPSIgppDA/2eSyUQfIU+fDMJ5+2dnX+v9VxtoywAw7i+UJGInix5j751pmZ7YnW
XuO6mkocG49GYk9C8rTPrAp/3W3s9V/y0GxJ99NV1mNtRtx8AlxUj+ZEApqcMkHW
UFnagulTzJKw9Cya09ddvMVtDTtW8JBfvb2lBhjixwUZfTm+4eRYHjXKr+sqF6OQ
f9hpyTA+QguwjbVZqqBk9L4/dr/Dtbd8tZCNOFqbOmk3TlvtJuDYhLoumiHau5l6
XA+HaWNAIm8Y+IaP+nWWRXYz9r4y4D0FodDEnur1CP6t0wB789VKK7cxy33vAWxJ
SumO8WL4seD7ZifemT1rV0Me82jh6B6NA44Lllpsu1EW4KpbD1FnJgDjxUZo1nm5
Y2OPq4XHZDqaJ4/LNx9FRMFXFgtOA6hokz0U9/hAFt3y5JxqPMy9B3xxEQY+3ghT
6sGzijhasuK4UqnmeR8jn72AlmIi99q6xyQWRf6P7m6VTwZ1ERz5YyUXDdrcY2ew
CqIz07LS5X1IcDZ17rlXcYS4/IDYA3v2oIa3LAANanXg9Ii5k3Z88zdhv7pGIbay
m+eW2YNFHzYKrqzKarM8dNaVq0i25oI01MjRWnKpEkjkn35GP2mR1ZkeNeoQWTmO
34ExH2qpCHdCddfsVUBR0bNN9r4fhCppf1S96NPN6vB7YPV9rbxGbqGMKJaeISys
lchvah0OU9SFgwV54ynFksdS1h4XrVIex0EMMiMfa2lGLyim3SJk7kCVKv4usgIm
7zqOA3Nlv3KbMjzEZxB2ZRKcS4ZG6+Ddgyz+hrCOzNFEbYKqs8rdSvIJKxlim/9v
IrupL61+UUD7vvrOncbX2LeaGyiBxMwBikMQW1SUTxgvn44nzndwWjBTLPWD9iQJ
eDG08IPXgBVCFqbMJOgPixYr1Fx3hehNn5Foae7BwJGez0ZDtGu1UEUnAVAlOCdr
7pr6n+1elxbE39QsU4KzCbufDS/KuQKYyEi3lHzxXyxMJTn/8nl2loPb5g5bJUOz
imAFoA1vpAOMpa7BJrryFOvIXazQkpsRw03IAwTWFJahWihc/GlDcSXZO4zgD1/H
EWd3HqUQd18fixHHcluEGpQtJr3bWYpa8+pSeb1ZyNDB28/R3+dO0e8HqNk9o+ST
0ehi41yXTQ3gYpobdVMFavsubG3/Ensqu7kI+BSrgovKpqoCOsHo3yTVKXbPMQ4y
woFwd5Y5PBmQWbmJKW88J1kkGsWDE3eCqgkTPujdyXydx8JypU7VVSPdYPVQryKt
GrHYof7WFCGkVPjFSWoQzBRqRTahDKwKmeY6+yFmlD1TiMJzlSbSG4TGbUrl3gUt
YVPyA+8Bo+SyzQGg/2GA0e8pFmFovzakoYeyVHoI0zJ5phvCnBd0dM/P3OZvG6s7
IXvYbA0aMMNhygSYvwmW3sOKrFmfic+accesOo8rhokujsRslD0nqMV3m9p68Ul+
+wbD4sPg+3GHrORIG5aWHDZUuY7EJ0fQ2Jj2OPNk9iUCetU1bC2Kbol7obQGWY1W
fmrSmJGTssibnjlkx7jyRZL2+zZpBUorME2LpbbjbqdKw+Wkx8GYUSFJ3O1ZtEha
KXDc70LWY7l17GiwiYV80TlM2Nx2jpRtEtM8GyjgyJcX74j2LXTBsTsIIfCgNmZj
1UPLsGW7Eh6MwCKhJGQLc52lXQb20+YKdMsNdnzaVOtpvYK9AdEEADJgfdeOczLC
5dqBnDkoCWA+HNuD0/pt7Lu8A73nXgM3xBjBuSqLS2c1oiQhOab4W/jX+SuzRKMl
R5YitUACSyQbvP1l+XGtPf0OLQ6jDD8uI3dhyRB+EH0Oifw8Y8Ym5W377e0iUZuX
NfcCF1SXjNlhlhyUNn1/Z5EhK+RUHCspoyW6BCmYcwwngtyhGCjnXFwqoZhPu0YQ
OvrmdMmu+8q2lHmhEfeLIhd21h65xb0fYBe2qNZphbwVyUTGF6H4cUWVrwllHKU4
LEsYnjDwYUx7x6QWpvfKKjkb9U1XYfSGL00sZIf2NtWgfUO1CVstn+XwdCl3Abix
2Q0Hm1MGE9FY3mua4oYLQekq/WApdAMyyXe7AkQ9aGEcyIk4Y/v1OnLArIS85Jfz
qZLEisjw+XjZ4OTtbjUX1SRHzeLp5ZlaWx/Ixreg2zUPQKfPZas5BF7NffjZFsL7
SGsY2gG7PDPA1ZiQJD7eEU/2irK/1xdy+0S0QheJLtiPtDmlpxzSQKbp6fGMSwjF
PM4vbW3WxRS/W/brT17gwVRnMt/mk1U1w7S2UoHIrdn/fuxI2YEaUkOK0cSvvmNm
IygQzXehQQX4oH8orE1AMICsf/tch7IrtBjmwAQkbN6zF12oF5HyrXIbqPObeIq+
qfBMpRUICtQn33KsOLlXynnyHubAwBjaJrs5YQ3529lgP/W8n9ip8ya1EbN4fV88
DEQ6qIrKuzh2sBOtCioFnt3zGv9yLD0IthtfPl/a2tbLi9Gpuuqu29KlgRRLLo6E
O9L38yO0oU9D2ArAKzNdqykA869UbUZUu08VR79cbNaLIMOlkjkzuDnK7e+ngOR5
iD0pwnUgdqB5dPJHwqfXZ3pM3R2lpHQdmfrUFPARJqxw2U0UsEbsgZZ0jl9jju1n
bEpaQxgU/6XyXeoDO7gxOO0+Ed3i15rM6uBpxWdFbGAFOoR57iYM34R11dtvAKN9
Xc7oMOcIMKAqQcFtFJJO6mXohj2eDV9r0BfuEY+5zYMi2VMhAbFi6miFGuXqZuFo
b5IPF6/+sWZLwfD/QpAeF1zDsnOD4HFJ3ssunH5deqZR92xNHvt9HzFgDIdj26r8
aEUtDtbWENlqou6JyGlDrn/jAmhsCtiBXDGPQJY5Zv8FNdWCyLQ73FDiduYaRcET
KuDnDfwlUtdq+DV8bwPPf2BA7qIjoWEQev3SUknCaPNlRI/rkY/LgN6IiBg6HpwW
KnS7UyaTkIqFYZmUgqLH09YWIfUv7zzaQQIyin5TS23Cd4TpieuCzYcyJfdmK5gV
fc5nb99YdPEGgv6FlcJVRMc9ruB8qbZK/AifxJKJ7nWaiavCeLBSb/OjRbZGj+zq
iUClRr3QfpX5SByo3qTRUW9bRlunPSk6GAtUaI65ZhyYUPNXqHbpw6yaIdlqV1Mx
EgCVNSJYqMTUKZKvb/QL1VFvJHTV9Q8Vwe3wHqQ5EXuNNW+3N+owjLWJxxLf2WkD
214o/cF+YBe0W8iKxxHVHQMaMTMkEHU7fbwVbKEb9VsDUMD4g1vFlSpWEL09wam0
EcHlFp0U6Wy/jMTayMXh+UisB6rtsbzmX63Klosgm9KO1CEN0lZF+UsKxzAiC5Vw
AfAlB8nrXoyuuj5E1gDIL0wk86zKF8Dvy+TmznTfYoPopSxJ7ha7ogzggCWVAoNY
8t5Njc4ZAeVwRHjJY6cZ/FegNO7W+rQirqfQWqFIW83de6PNrzW6NsgejfL6JKZ3
S/TjrWhBHG5y/6tlQ7Ro3ET2+nHKQatFSI+Nu46cIUCKUITL29M3pVDQP+vyZJmC
pypBV2njTvOKNelh/gsdThRBnp6R5/KAPV+f4+WqFpxCdwsaQvyxMjQzxjVJhKtV
oJCa2dJcPrc530QG6X4dB5kV3MzyKdaS/i4D/xnrYRule7rIu1qNz4sn5x12UmCS
Pvf2AdAF/ggWwFdWlV+vNbEkO0yS2q0hULn8KUNqQFMFCiy3zHCw67iEIZIDT39O
UhcVgcgsEx3iFlBaKtX5TGJJSj14HsY0OP+UGf7z4KWyjlHneBZPS129mSAwSvcj
oJYg8rycu5AcFLnq5PzA9YDnDnAHmlOZL5rNWokaoKCWFg9iLuPSJzf4VxudLfWE
rg89RUheqRcSTQ4aFoD5GJWG24JM41SfP9zzE1OxZTIIuDJgbPDDR+Qf13JZD3uI
TyWXlPBFQI85F8/Kik1kIguuw+Nu9HcyzvhMpGwMSLuorU/pelF7lnliB4GGoqlL
eGSrKOeQE3rWzDyH+bblFZ5IhIkO8Y8IYupQv7TODblErVjqEiP2d3KascqlXYCx
yQfsP7OrrIwM21K218qYMJET5FNCwA0k1LAEyzfcy5yOXg4QqyTqt4kQ3a3Yg1pR
eVG/5kJEIWuV3nual2iSQbhNcHJdlAO1RGe34sS+ObRmlUafhT7auOI6ax32vOXD
W7RePpHx1kS8mcyPK8adr0JLDDtGeoPX128+EOJWM5L35BYUjCYdH1ZoznlSlKfS
l1lJhlsGe73L2y0k+ekNIFaaRRZCZPivLbvUVyQC2Dhtpezxfy4vpFSGEMW7x0ZU
kayCLsUDto7qiaruK/1/hJU0pIDPZ7dRKJgpZAKAd+jx6JOUEgYNqBimk2LreRzU
JMAxI9ouEQT2EqbAMgjjmODcvhdHIW4DO43grwdHUgXJAJ+3yhoiI0XkZvNuxi+f
rmV2P3AMIF5XGHP7zcOWuTlQcLEQwBi4zgtPcgjGCerL2ZlFqoVv6j2tnzJo8+8z
XtS6ukhpGeyJj9IldptoLvJlVQoT6JOdpdmUFJkegpC1vfZm07E7CCmlHUw0DABS
94G14YLRrMWkn7cO7zl0FhCqz37ZCvCoJupLWQTclOUW89/SqgnZWCW+OJR4tzox
ZeyGgCLfrESr3hdsPcwxyYQL8u4q7nUQ16t6ucQLRNX44PluByH/wjAHmiLq5/8o
o4IG6bUpSlra8qO1WnjPf72r2BVZ1w+4BGiuJAUnu3aOhEJqr0Asv920jBbObdHm
mmyMXDNbR66UIbJ0czbl+7JHO7Q2KRew4h5VgUg85v9ajMZfSkBXvcqCsTfX4tdb
aY4lOZVpksoxSEmT0HsOnPRVdlOvgnPL4PvxtqQ4C1JoIMME4L4ex50sRTJireJc
+d4Sx39mpEHnnrdD67GxV6FITzmwzdL04YyqdvMHkr6Gc9N9EdW3OI+aSTljhR8F
U6vQm8uqr2VKMw5+DTZOUlWnHFljh3EQ9S5I4OCiuw18hhtM1xbzLCsAnc33pySH
LKEpalDQzu8Q/XcLLErzHizA+z+g1iVEb5GxLtbD/Qd8+LOQenDUpsQSgID5vm86
Yxk2nYww51I3GOLAbJegJNIIpw46MTuPlsC+Jz8ylG1HMj6KMTzzZpNBM1cdy3UR
Nkot9a0gUEXeA4hDf4lE1cPALGfiROyZ65DW1MWzqAAD0OFFzQB8Mt0bhF1pSGbA
vPqehzE+xeIWMTDaPhQuaveYfSFjrafPFUSl6O6YS801Ab7+VxdVWrjk5B820OT/
xU3lI2XJRJBQbLRuoQ1Qbi4t1o/VKrJ8FqVpcKCdjxAgYFVnzJ/W/+dRcKkZYrQe
CEO6ptyqHmDjzMl2iCLw14+524XAy/urEvn+5Eu0TyaMmzse2RWuHv1bOhCYAlNw
llFxSFk5TCiIe86XOIFh40OOs/TWyuxHdpjkZMRCYW1X82MbiGNrG6hGrxYgo33v
i2La5RYoQSJMVQNFty9tFXxI4d1Duse5Ve3yOGdOVkxgo5+TbavjYxxhmzxt0Rwr
ylO/OnxO7Ds4n5uxPEJbngDr4mGGCFuKy+uarcJPPurMeeWNnbYf4FW1cX/oUWMw
tTJ/vaUrPQJJpz+Owi1X6CcMCiCc2b2USXAsU7GeKGdBw6s2cd+8DlxQiiRCZdFu
yLqgv2kbcsWe7xmuvDYbqoG1p+obHuC1G8fzk/xpqlhf9TvzsnMQnNXJksarBV0u
VzQsR5xFkfJkwrySoP+azJf778Zd5JRsG/NJO+Mc6+klCSYVIzPMknJinK7bFfXY
g4s5e9CVN6k0+Zjs58/XvE4kOV65XaoG8xVkS2ywhInrC5uvqCXmX8A+iTARs/FY
DX/6m7dbLPU7rOn1pcPwOAg9t25XtcmchIVQ5w2upcLGR8++p7FVt4NvCK8bJMIC
kUzyBfHbbCPs70SPVClMZg5eS0Ked1g638DadX9Qgys/gsOu+K5LU3j/CAex3TQZ
TlBxdTqMIQjWOo2Vf6mIUfO6oVn1lOZgKz6G/mddOccPaVdReFCc15P5DVXeTkCc
9/FkhJeDENTzAPn6iLh6C0LmW5RsI9ONZk0nwU+igIKr9QQJWpxxRK63zZ8fY7rz
r6o1/I6rt+hhkLJNxbzNiO7taKWcn/GqWp3aR8M8SVsMFVLyBuKbLNM2Jl3+5oRK
fCPkKoJLHa5Hi/nubXT45Z/QfwyaB6q/n4I/3R6zWPO6j6GFsnLIVxtEt5Km4f+D
CeOWby59GX63Qw55u+Do0tHAgtF7pQmiWcj8yHjlGl7hUiTOsGcq72MQB+Ammp0/
zX4VkBsWjcqI8QtlxoKBC+JxRKAwb2QMya8NFymkB5YGkXhep3VZ/t9nwLPnMEUL
I6e+sG853bkMToh8LhSvg3BuHUx+TDYdFv8QsqGefVfXM8upxzGwhD2XY25DqEh5
XYtylgW1ogGQSpzkHEmVJSB5Hl0/mLr5zyjN6QUyduIkfpB74kXy/6W9aLeu0kn1
yGZ3wGFBRN7/XbQzkRz3AKmtYSiK2grez4gn+T2Abtv3sWUuq0MZuJqD8+qhahlP
kcck8d/DBhhdjTMUqVXFyxIBkcrBxOX4kc2lcaS2FA8+ckmLnTrIUmo9KMKqq0d7
+nErLsrxGQn2lWzZdhYp7AOIrMhqIe6T4SWoWfJxnY8b4U+dVmy1W6QNPJsfUcMm
EX8PUNAXhVvFPLjAVbGVVtcwH/q9dX/Nns09IhGuOjmObrSmVtkC05D7S1XFvPnI
QpnFdm1euGNYmQv+yeGXtJ39CnIfcgxq5ZU2ErI3XKKBYIE31tlVL+ck3B4wWdvW
51xZwQmPqn/BpGyb1v/gq13diSJasWf/ugsv5CdPAxmotHLUzL+mI4cwxDbTUor1
kkBgxThUmd4+ndVRUhaq1u0UgnBpoDxWBjAEGBVm3WLPztJCUYrhpW7DTrXdztAV
R7z9W4w4G0dNzAxqMr0eVu9XfQhWRNJkwwLo+M08aYquflR+GzNFoNj8NlW2KjvG
FWRUW6I9toC5/npUVcgDLYmqV9nBWFExiNBuGVshjzz6Y2CnA/dAdCwtMD2ChHb6
9JxI8SixIjdUJhN1ZY8q4InFaiAuDaMqhVA/aXYDJDZFFrzqg1OYo1jVJQbvADon
TZcLTPc5UbjnBkLKSfVdUUDOAHbbQPgdk+6QAhFNKabSDgykEq2lCFtb3x8TnHBc
7Ois56tvrhSDMdu8+P6KGu++uVa6li22NW7NGyCwjLJlKZTvcQR41sfnHYxzxTfg
dfbJo6CwcZ773j2b9gDfskg1hSN+dmshRNNFNXl8nIewd0srTLPeeFRTBKJFBGOW
s5VOyJYVhr41ohJNyTFgYqUP5ERNlGuBP1mUgczZrtqMsXmTjAClh1RZ2iBY2dfK
CwQzpzcvsVh2Xn49Eg5W48TVs5E0iGlVQ5KQb7i50BkZGcq30UHdaX9TXby2enrl
Vi/+nsIRQehEPWbmjp1tTrwgSwR6o9Jo/hNZVi5rZaPibqExA4SNb4nq7BAT690b
LmafgfZQkCG5Rk2wBDaBQR9IkIFSO7QAR/dAcLj9KVHsWVb2TPzznihWHdSQQM2s
X014fxzk2w4BmyYJ/ZMbmv1vgwrQaxtMhSPDfw+6K0mMb9y4rhVBPByswtg5c0c2
yL2lKjVM6sgLYjLnRZ+SF9VBrk5aVTWJVAfQ93b1ZPnXfN87/7OgVOw7NAYAHduz
gJXOIEuf8ohxSXdumRG4bolaWpPlJYCyhmU02R/OI/0K3RSoPJFYQddtunk7jyxb
N/6ErneCNFNheXnZPmIj/PWuAmJjijAhXqYfesTjGEjcPvCRucL34TsXzrMrmKxo
5JnYsLZ762fgmma5ZUmUAD8rRupjR1BqcY9n6I/8kGja0vJRoQ4ZMKOYynP8b+0b
HeMkQGfbhG5/stqXsumT5LeWBx+P4uX/SzkL6nd4RVyICD+lrXtbp83IPIb4ZP8m
P6deCPq0/M9bMnmSSf5/YhoHuADnB0N3OFO31lXZYY1dB8OKLJU/oQGpqfqj8tZy
TWMMNcD4hqzEwWVvdTG2R3AnvOvVpcHXtqWGJQEpDlXmJKUxwZmvBdBDPm6OgAIw
vg9gg21NE1elJW6Qe0gQjYbV0RAVcs5SJwDPJ8ftjD6W6lgKtVKM/wwkFxBf5QRJ
0Rs9ALy9RSGhdAJC+4Vf2N0meKXR0P2XdZmisuFBVJdYWhJwzNme/Wxm3rMhi7Xq
HR2zv8TOA5V596Dt3QdNBi8acF7go33CQ16dwA3xik28WnZ+B4kb00JymOc4jqLF
sBVPXFIFB4w5Gq7yOL1YueUUqb7/n2qEVPsLECPpXG0Qd/JQ/zetKCaU8F7osgJ0
M5HkU045p/0/TWwURzh4jYmUlqmppZas8Ex+rfO47IY8Zr2RaGo9G9p31hDYAeHR
2xQlzTl9vmgShwSBwSzeWNuERYno/fLnWWy/86CQfW99Ttn+hlFoqrAxAd0nug23
zKkDPPRkvMJVIKm5nE2DepDO5IbBYHidUTWU/8jjfOjPqkWyr/nNe73MEdV5itxY
LY3ZxuZjMM3Mixdw/7s1YxTPUI0+HZYPEiEIwIkk0yvFQjUGVODkqTA6lfacpDiW
7nTp3MnuRzymxymzln7XRFgpTtIgBkoJiNW5m8SSNy6eXqQNBkyqEPPvqwf2RApf
cWW+463Nrd4tohwWtweaiX22WrTWDxA2ejk/PJHZBPXAfkLkOhnOUtUuDre7SkxZ
CcjcVcOauiYnAjOmuH14QOUodF5B0uIKND35xsmVaAAG1yGmaXQs60Re2IPX6pve
qLEQJoA4l7mOjntWVM9oA4scLm1M58GNLeKRDIv+kZ+jUUbIGhbgdqswU5n50Izk
M+NbRKmZBclb1Xf+FetpaYBtDC9xHxj7qgYYl6EGvFdRj5UaapWK/6m6yPqY98Zd
ni4G38hlPrc/q4Ejg47YsozOeXj7/2vmppq+V37PNh9CvhZTU0KFpOwx6dADnYXz
2l1r1sauSRXKTrljUxAsecFzeEch1a1DAO9kQJpPxmKIDamcE+QH17j7mQYfCf5J
kStl1Lk5+wbinrcTryz2rIDaCQSEBcOqOzoC127fIaGZXgPxSzJ/ffuNuOjpDzkU
I+SHS5cXt75gOc1N9mjEL6E1nRsCFX+KHAd2E1sGyHs0YSlnVGFTOghzhmMyvYjY
wrEejqXjUX4avlXv8RY9g7QNyPrnGlXMH9jTtfZruoQitgaIUhDmup1DWG3vhSHq
uUcettpZ8rsEGor4WNgSZwdz8LLRjS1KsiPOH43GUqNp+o7st/5RcWkSzyIkBUC9
DmCggYC/y1gc4R7Qs9FFG1pZuEvoyUKZ3LnH/YNh9ipyTma6EzRAhaqVXHRNdjj9
WWayDRhbuZCS7xo88HaxMQsKJR8Lo2kaYyN5fiGctPxblGN8Y9CeEJr5Dovhtuu7
hfn6wccl6XuZrIlXL1AbSiJC9xNxxSo07PO8kJxTXbTohTIIDbU8ZIwYGHXVnFRF
fz9qV6664BOS8pomGcwBBaTh/OBMrbLt8td/+556nvsd2MOPXJq5VupwgBDE9Xdm
vZNkF2I+GYuQiZ0o1nkV0nyNNyDBQiLC57y4RXt27DYBp7R3EgksM6rSF7zjDGTo
LrLbQj5qhbw1lw5lLCHmU3478p5GZr+YcN9mFYLSRA9QB8r6+W8vJbh+T0jFzhTJ
/WjtzJMmBuY4Qg3t7wSeRIgIlshDfcTuDEIAyffil+t7w9O4L2ssjR1CwOspQNbQ
mZm0x8HFmCQl5GgUcI1UIfpDTFSPGhy2PXXaow1+v3YMLWPXMX1AKw8kkzEUvBID
PFv/pJWLZFAkU1nvK4oUehNRel+twMbssdq8RSE7QwgdJINtPGVyQCJ66YWwlINY
1y5fK/bKBQSzMfqKsNpwrVlUVm3fQwrZDlSO+GU4uGGRjQUxiqzRsqVGqw60osv6
7CA8RbkhDQyCPlJuk+/o10UUK5vtqQN1Fd+c6VO/ZuCwi0tZbTENlH0UKez1Vz/v
jaVWTfGHT3zNdR0D+SmUIvmp06AtzbaavpcKsu0hweJaHvywB7Kz/UURw4pFVpO7
ZOEsghaWVuT6tTAXwt9gmclQrQ8lH1PbeJJ7CwanFfjpiVkfKenk0kFgyWWQ7W5V
37SryyMe8XSavMDy4w9bWeWqcwYmfxpne7yq7zD1pfDoQkcmvR/IvrdsJfs61FIE
p0OyBcnUd9rR8j/4ebcbROiQCPQ1gwz3+5nEnCUS0yGOoLTtblwJlvJfHSNaBH4U
v1I/SlgfzbpFLfjwzl9GyxUBxRZAwlk4HTt/lCA2mCutW5WQEA6gN5y0oceIez9v
HTcGQft9v3e2j2u1YYLuyvp/b7b+h65Il09pDxLCDaaK2HD/kkF+zY4POIUTFZee
bKZLAkatDK1D1J79J1F5stE5bGbZrqSAIgMO0mtYN3o3h5uLupGZaNlvwpL90N6v
kwPB050or3evrV7ePh0yjijqms3zfKgir1suKQGjhO6TWTSZ9CvjDGF0Hmt+brUB
Md+OIjU9Zbfkzm/d5+EPmCcSx0dHafYXrP2sqDZn5yM47Dt5KTT/fPYdARMaTf8S
kfqxY7JTs9tUS+pVcXjKIqWoGqrXtI7vq2A0BhcUcxiVGxQind87WdjXwIrsFYRS
Ivb2TqP501464pnZCk2YtNZ+FIc1V1qubiNlsb7Qrp1OVjkGs8vUBwv58r3EwdWH
E/SYg3w+3jLUxbI3BGDJ1mA28YOYSijLNC10z6IwJXbYmTPobqlmydqbQlqbHZ+4
sADTujqtPw5GSS0oKRUtiBM90P8EAxc1DXTw5zO1UQ+8EGKbDLWkpcHVeYGsOiwU
+bGUh3Q+5I3e9ewl8Oe4aGFEmnUvrwKL9Iy4bVTugum0/aiXO5AMmus/OeEF4SrL
HVKW85fNR+pbpeX0a0ARJThCfmjBFYoYlMNGZr2sEMW4PnthVmWXYIgj4VF0j9an
D3w0O03Nvqyq2dJKCHcf2rB8mojoLCv00XrL7tvw1Y5UvpYqs+bk3FcYzXFPXwwJ
yusgQXinmpauBOoPDf3KI42spli+GtLTSG62kTasEjwJxQFmNwsSVdlKT+h4RcnL
WpuhMtLftDN5CRF5Vkv/FnkSbEoHgfSvjAUXdqiiBH04CuE4F2Ift5QBhQ/x0b+B
B6Vd2A3IiOgW9JE9z6Y4Chw/0tgRblsUFfaqIGzcY4l4RiUuBKTUuYhGe3bDWbSG
HSug++v6CYfC0+My/KZr/ZOkqO7TvzvzOtPkR2/TUps5J5zauaGjAkOLRnSDCJM/
amY9CeUwkm+opm3EA0UPkLWOTkT2wPaIf/jbcJlprqBQxU9raUr5O2Fb6zvkwmrl
UF9xbym2SPfP8bLvqA+C+AJxh8kQeQxuEtH7UXeNF4GSZyvRIynZ8Yf9b6l9YJJy
+OxDwfB1F/UYq5cZKdnHN3OQMZQzGZTyKJkaUGQwYyvbHw1/YjyPiPGC6KSm70yN
s19c2BSCbGFW+1zUnbZR/YdV9GscthjH5QVRJxrBc7JXV2p1kvED+6C4ppNFrNLP
Hj2vvcvDoLzpKUNvy6V63wMimb5rqiFIhNioeIgAc4ZGe3lXSwQyp2wH2v3X/wSp
s3uW3XK+kT7vAdv6z1vtzNfgcqfH/2vBwBZ1mJqSNrrdj884GZ79bmGtpKE+3CGE
4Qorfu6eGVVF0Ab7jm4gV1E4hDSWR6E6zJPiVVSN24QTE/doJPVMS0F+/HTN3a3o
PrhPqAZdSIGpcteR/d7We6KAwwdvAN1K4f/TVt0DVvK909qqrNUYHZqDvQH6nVDl
h9D/ozJ9f7NJ7syY7a4HM+AkXNv0vZbejlUZD2xNUahYZxOy2mitbiXBpTreI1H2
rf1njbpJQPllZGix423rLzu2HixFXRSgQFnEUMNg9o+OaPJGE5p0PZBO2+hAUn+E
l8u+7gbp6CrjdLX2i1ohxAh8yCzlqS5kIn+/sRoHLOW2WrXfB79DVzju7n8hJx19
0y5jPbltbNY1gkx1DLuSyvcLebappi7zP7VZlzHwZVSXgN+sRdJWesaRA/Bb0AmV
nlE1jA44ZlnOZP5JFKNRdgk3gY3u8Bdd1gO4OpKI2EKiYlLs8luh/kEnlMMM9i6T
1Lt9IohfQmGajfT3M43rbdmo1eF+mtsijgCkrEH6M1Llq02vDTmwgiHd72fmPol2
f+J6AH8Orldb7i8XbRX7dFzmTGi+wJgAcAgsXm63N3Y+BdqY1AWAsHu6lp5iYSWA
crfjP8EIQ3bj0I39ppoTO7N3RcYdt/9im67xVE4lpXm2qGQ87WwBk7oaetdMY19n
YULMgvC+0pbbnwp2gWWMw9kaeayiGbf+yvEBuzP6+QTKcpgMPWYTDpRA0mHSoQ9y
Zz/Aep2E3CAKiU23Btr1qq4AolJgh83zf8nw5f6iPt6yTwwYEEXTtrkkiC/zr2fX
/9+OdZTK9jp8YuDr1fPXnhZ3zdYBcU5PtEL8D+g/o8r4obzxplsIQ2G6o3FOOAUA
ww/D6Se5j7709TI47N4UFzi0ys7UvwxuxyLE1vXH2iZ0+IFrIX6vluFhECQbjGYS
gt2N79FtI3IpTC8TFq0bk9DgsOCtN5MnZ+a7iFCZFRPgtPkumuiAMFIhIrwnO7B8
w2XfkjugdqjCbomgElkN1gyqvgwTJ5eMJYk9mr/MIWMq7JaMacbvApQa9Pe5eiTp
H3soPvh3PVLAVZSi8cK4W7NU9Vv+/UF1P7HMGhLcaPWlz6FvR4aGtgk6qR1kJzN6
tcsakkj5mOEIDqPW/L/ahQA+ExNjURztkryXEHwlRkxIahz9uAyAaAB2QkwtZyqD
gjm2W/xvnSgiw9b75jhfsramQ9LzTNJjGrNPq5ts76lMVTeqSszR/8Bd4TqD7hFE
+39JmZ847pkacRsNgg+5jIGimEsSpiXLoR+K1fVAWoJvrngXJCMaPlNS2SEUZnd5
oVS6iTOtHjZHkezqVQDe+7Lx/7tLr4q9CHhHEWe6dCGPHCMOXFHT81Wx/sl5U7So
/e0rRRdcb4AYLvxiYWbmJ0/MfW7QsngnJbgVvWzT8r+iEUibFvc3iz3wOGbY8u3U
gvnZ7Oo9wmNmoeAknFKHzIJUA8ll4tYbbOdr7MNSvDRsJBqhii5zVBqobnq3cb4T
X4bOSSwYB0FNzPK9Z63vxFkJ5fOC1gYfncKf1RjEV2xR3z5lN/r8UGpOm3QVZzza
5m+5tR38+go+SgmMRertHnYEHPevXUYp0t3O05sUQHxmEWluyAZZY61wr6W8im6E
M03mqkK+UqjMAVpWYr0tHjSWu3NVr18alcxiC6gLJUBKOAYJ/9T1mWAQjEV3D3w+
RtVXhNcvVPUf8sLQbzgCwDkVofgchKgwNnRG0RrHyTp/+P/DvIJfEygzdPF2M0zR
jpIqqCrLtghFvFTvX71S7ei7K4FFez+P+Hhx4jhMCHb7hgRwD/VpXFj2i6TsO09W
eCUaf+HbpGD7QLqknWD/CeNocr4grQd1oxaOjH+3Z6GU5dO/4obnWqsi3Qsm+iwI
lt8YKtXoujquUfDnuw4twsEgM17vkdeJo7kxmO8myRmINVaSZplxvXCYg+PJOv2T
nDxNF/M1NxLKOf52gzU+G4+2BN1Bs7n7EwxlQ9jHjMgsUyj3ooq1frwiuQVc5Ufo
yv7cFoxRCATIFE6PojFDxtnJeKyPYTaJNIazSp4cRmIlz8YUjXY8MuvULHUH7EGg
Ub8YYcCGDaYvo+QPqnsoA/ITMaVDZsnkZLx9IdLXwzetZ1Ux0ObaXwTOa0zreJ8h
xUQGVxjfbeVmRb2/tPTjWjtN649F04yA7twXFBUz4kme2agmX9l2CHnjmaULz6MR
BZZz4XKn8fUcuC43KVQT4oPAPANyuKF6v7Pe13L5gGG3XeeKheaTSg3ZYUcKhqjs
iCVmBnBWyieozidwSJcs7/LQExSduxitgjfsDKUDCSuTxx9RllRqzE9BPwD7Ja7b
goSeMYuDkJHrQ4j1vFVR+lyFMGn5uQO8FOEZFb1Ro8VHucS6Q+q+AtVGM4zWE5/5
6lMzf+bPGAS5yKUu9BkEgUNlzOVZXCKiOH8qnodRxgud/AjjnzEFqu9kAfg5i1C6
xf/QbXtujVqZdsYjlWJ/opmoKYPW1YK1q4gU3ttAMrfynDN051P25+Lx4O1vbNJP
Vx6BWKbuAKlBn3CXkVs+D8S8xvRCJppQJQ9GQ2zJSFuy1l/6tKAaGF1Jic1kRC/D
eJSeoQkH0kx6j8vWZ0W1PehoazOTA0IYTZURbL+DCcw6k2vOH+jhcv9XYtRnSpj6
OgorZo2kxohureUKlirq4hLyZ87piS48NK/kjp0Y4YjTmTokJqO/zVv4GvOkBpYb
VYNUk3pyp7vEQlEQXNT9nA7np+YuPwzyrCWTrvMSoqGIPr5ITKAYXBjXkJUxvh+g
UC/NxCDWXIaQvn1aB2rWWffRSbRcZDrzTWdmcmDl23V76KvfpsonhjYXAODz0V7B
mnei/RJqME3SDSjoyedZQV0GMAUrSZkJvS4U8mkiSowRU6k1kDqkednJuFxd4Jz4
EY92ZRNpSHMEd9gWaOVdwSLW0XIRsjIMZn6MWffkLbt8VBTGSaFtR+rpbew92uOk
tgv8EQhj561oHg+skn+ADKR7z1A+zVCtrb9e/fLoP1ML+1yjYXlmR2or45KgdxIJ
TI13XW+aCBLILsfihb9bEM2tsbkdTvkeCaIyOqjxn4344q1n2/GStOFWus2xx6fl
EueJW/Le6PrNVwoOmJ0R6q9Cs6aOpnCXg3arpi5xd3suousESicvaZvazLIUjplv
JGpnjmnp13vSzyFxNJUnkFnNwr7F757fQj9rB4lORvBkDJgGAXcgaSMx/cxSaoFg
MLBE9v5/zcfLJotiRaLbBBIThOzd5lr66bo7s/jVDeSc5wsSuqQXAVwNyIe/hsIy
q4kwwMeHlJS9fqRMj/Z4sPDDQTszUrIZdhVfxqv23KkNKSwTg4jVdlY57moOHOxQ
jzGC+9uWJB/ZdojFlwKPWTbkPwFGGyvzUjLP133+geiRTZLFpLZahmvlZ5yKessv
/PvlWxm90k5y4sm4fDqme7q3Z/mT75WNeqxkSBQZmM5BFzOINw6u5nAhH+IjukhV
9KhdoLmXbLSFoH5/0dPHnPfx73+ytcZmjZafzjp9htwzLAY5rmZVvQWQnDRYPUQQ
+Jhm452m1/0452zCGz92w+mLBub3ky/WfQD9OCMgGabpnFRKFnf8sIaC+wNtQMNR
VW24PxbNB/gowTMkALez+cWZqWnm8cosHxemeCUYdDd9GCdt5BQMPFJYFt61lVYM
Mc5y7+JazTHrMplPvu67cxT3MKpr5VMJQyVIzphYsP5uM+G52DiGGFUn2RIts6vA
mXJLWc5UmQ3+zNOTxvWpnvZsekLk19YWZ2AFaKHL+68WRcl2/2kRVpW7FAOiIIUA
fmygKr0NtXmlCSPJI97sc/7WuGhXfKQ8RffMp8h6lh+OK/PkuQw+cyBD8gRD2mJ2
O48CeufIE/OlSv4Dry4YXv4CJ0nTiLP6ahWRzSlRSU5u2wqCFU4Cfj49y1XQwFhQ
eTDKNrY5eP5/wu144w54kize7AxdwaK5RwuP/V3dwdug/v1o18imUDAfBGYRpO8c
PQfRSwI9hCz+/e3j/goPOCkQw8RjaHTWsDKBMIePI+t/XNmpy4Z8EY6EY3hIxeuI
N/JeUyTCXQGCkbNhb0fq6Ms6r/fKCbxBJ2pmKuSZ8WgoNss9Vhi2p0uZTF6l9Qh1
JjEe81SsJqfOEJe0YlSmSeBB05Jmkca5YIwJAxLkC1T/xLiiDl/5NzzZh/MZSgI+
VArFH1S1r2hcRYdJHlOv2JXTfIdqM5ARxaPu+cjQf3BR5FZoDiZdTA3CQK7/LDgz
aPQbBqkQbZhepr+Ll2Ig3xjQpnP/vz4dnQBBaK6SWfj7sBA++6rENEg4iYsJWgul
2BvKNuWDSYwlLkGJBj1oeujZqEyj/TJtqb8YdnKs0zgdYbgC0YmXdzri55OQ9xV2
2HG0EUrG1DtbCOZ0V7rtsBhqHsrpljvfvbq0jo417zHWkpi1rVC/WETEGuM9yCe1
nrkMgjCeRrclBlnV321cj1iz8wQnaRV1dit5gk77QX9w32R4ax4khb36C16fBoYN
ONr0nt+P9kyM4nc/JLBcoPZ6V9Zu7C0ussv/MivUgmSi8mgKunqtiYCZeOznSsT2
Z/brfdAM616wsW+v6mWI27nF1pCF0roxMetcgjl9inNi8DgOy6szlteMusHxduBp
TQASx4EF67524kk0iJWqJE3lhRs3uIvelJcfhCrbIK849WMjL+Vfe07DZJjGHlvq
bpK9CV2deKxOwsUl+CqioDhE9hK99rjvVa8Xob/BAm4mRIfEj5nWpzkEHFi6JC6/
jrNwwfNl+M0+yPeF8T/azfo6pvdDYZsYJulb+tQ4oTI+hYcmpDajg9CbrdMb/qnH
HXaNf2OlEAR8j31xUwSv3PSVjEXA54RmNnfT57WKQOnJaZoYKUGKZfGv3yRiR3NM
qeTQgMoeIe3/hXwYCF1evmgHhreoI2xy7Xfoa6hpbx+NE9vqaEF5XhTpROW0SNDq
amLsSfQpWm/lLTK+BQ+iodf6PbajJH737Bqa6gqY90ApZP85eHNzDdNoxMMADxzU
A3gxEH/ZfrFrV5j2O34qRjqbU32rHVU90hGrWHXrDr0IGMbdhczRdL+T6nUMCA1B
CmkgHjYhlW9EPwR5GDYJzRzPw35RdJWhygA/w/sm+9SnnmJHaYV0Q0ZUExH5TvGP
jm1dIVy0rd7/8ckikFxTKvXtFoZurRjwmU2ZRtMYwJbond6zfYKSXMkEzm2WMWYA
jnUOxkc9YxkMa5n3zyLJUrj+XGw2ohlk8uxT8CcZhqsZe4Ws1VjVahBFRzxY9Ni7
nTnS3dwAE8miQJItv7F7PitGz48ao0N6kgC6iFJcFzfUhTTMC2CU/DGmn2RHKxGI
5ttkXqn3wLMbkdHpfyP+ZF2OqcK2HJSVLWRx4ZvWQKpIXJDj7DLLGk1h00whJbmO
rNnPrt/Q35/mXGS8woTIUKBAt98HUzjpV9faD0n2E2WHxo8BCLhsfvoUnBV3nxe1
12UdAhj1snTvdWq8eVXkon6HEL5iTvxGHCjZ2O5qIjGTDw/scf3l071/TQUaA++s
w95gJNxJs/WjyGAAsz/YbrNVg1og1ghfTE27g14Exu5k0WsD+tJq1MNQALoo7FVu
BdT5VKoUXS4wakN5sGr8V1rIndJJ7sBqmh3rkp769ZmPqlj+kThByHldwCgpg7Es
kcz0TeW4PPQhqXxipJHfoAsLSlJ2di00YuCn99SfvWrcR8NcX0/2FQurQaqaEVmg
VJAowP6VMdkS8HmKAigQWz2Ocf2172O/B/lvTq4k5dvSp97L6TpIbAqI0d2JvIEM
zBHMHLpwqgmNg6F7srtfgC8q+Gok897kS3XZX75FyEfQpLSMy7Khx9AXPtC/5/T2
cSjYteVehKMO8KnFugeDypsOjxeYmmeiZ/ql8+St4EyhCYrI6O7mTe9YW987LXhy
kJOaoYQ0UqiLDm/RoNNnLMbNPcYgoHIW78O/VAAJrOomwMcVqFALgWhsisa0bc05
BjgJi9jYGwNCze077I3ZfXcKOEPrFCKDC082lwxkMU97T3CyAxXYdSjQYZ8qG7LH
FCWoywYk60bzJxyaX9yaC4T0PDvcNYhvLjzd8RDQA+jceFchDFcWDevLLzEOhFif
i+Rh94lAbQE8XBgzReDtWPwZq/fVzzr+X95KQS+VGhAqiXdTNHH3Xh3ETCvoET9x
myMs1iBVRgam0vEPfWA/Mu5dRlcKOrN3R1iMAWGoJNdiIvgzbeAy87WxIiCiqpvz
7tBUOxKJ4LZjvnI8aAkeFU4IskvYg6agrbJnDhL/OkKD1T1PP9R7m5FkqG4SDFtd
Js3iVh2bQ1kQSjhTFLwMeqXXJec7VGCrxB7q+6QoL+P/KdfIQtP5msrngDsxMqFr
hTDtKBP59EOxV+UbbEf2XPyj41OnsG7csxsEAg1xFYHonsm8BtdnBtfs/5sH0n1k
36pJ2y3NolycDjqkmpydFKypW0Ha+IAUvlZygyUYi5jhs3LrWXL1cag7XEa7582N
zjeFyMuDRcMzIzN4j8/CDphBLkelUiSHc/Ow3hW1Tkl9E3Ye7501+AAaFBOyDEbb
0GerL/DogOubkTZx85LmDiBCflreJUFcMJQywepBxDmXJS424HbO0xc1Q78V2+o2
woGXXcUtLwISBCrsd09cVEqaeB470euJULtrN6v+H8SJuqwE2tEOP/X4ExalZ+hW
5Y9rTBNQp4UNPneiLz+FgG1utPjFjJap/oKtCaC+v639yN/7lm+m0tA19pVjBAah
YFGEw5VZH+Qtu1i1ZK6uURSpN+URTuwrJ8FXR8XX4FD/j4Y2JElAyOOOakq7Jyhn
6+TC8iNj6h0J3qjmgX9owav8sS0j6t4LviGMMbv/sIZow/3tGqOVRMfycRX90JFF
v3m4DfZxDsux8X09xxSB2IEB7VIen5qLZ4AU9RJi7JeG4ixMDFO4mZbQG+MKG557
JcGcyWFXOhg451+anwta3vPsrQghcDxXnE555UCTuZOM1PLM8bWejxoIFie7PYaT
ohG3ejHoFj+vNqSR2oCUl3fcBNKA1GI3GfPQUhYdkS2YrZaRdKZYai93ZjeXYR6h
4J4AC34BgE/CHSijbxzwwchR7Pl6CoHUr5a/UXTOZfnZJ31582aaLiFGkmjaCdw/
0HzxOgqLkHLXqRUCGDIUvDWwq/KBW4jYDJuKmRMc7blbprdA3KDY7ovA0d4Ric9J
gJdWusGjgL9xVBXll4nlsIaKdQEC8pqqxoUVwpdqXRxRIFsJdNltYzMGkVjC6ABu
BfxWmXtAv9gfxrTWc6EfEGingaefx1iggAvEPbbG8kMetDOrd/WP3l92g7GNpjnY
qJYE9KkIxGQmh0fhhdzj44M5TTYFJd/4JY/2O8o2j3qL8uxthuKM6LFX3qMmvs5k
gjaXLXcrbVO0jIfCfF1KUM9NY6R54zr17t7h4TTKqWIYHQHOWXwDdqifEPcoNnaU
h6RhJP4/wFnYF0j9iH1zSiLDYRDUrxaEWDnBJ8O6dYioRHwYYRCMHYY7C4RmWA/A
qnRCyRVGh0DqZiuImIiTUGC60pTAkPw0YcjSRD+xOybE9wH3JclA4DzlTEfGA3J/
F+7R5kQGcvRflE79lJpgnF9ettQQnsZwKN6oat0Fggl5wvOJqQfO6cDvU9PiymXx
VPLqjREBTNeDyYxma6Zb1fYXfD29CWYt5JeftANw03gpiSacscaA4JUdwkv7wLrg
3oGEHz3v6iGYaBCEicnotZhdR6FW4E8TntDG4RxZc4rvTvjjd5iiJJ+PL0+aT+jx
R4XQEKE5N82MZxZqlZGrP0V7AJS4jv0SHh8Mv2NrX/XGuDF2mrkwlu+1jLff1seB
YPi2ObDHrfGIlwqdLl7EiWwozuuuhwNrp376CWcU9emvD9eLVvHCfrdOoVo0LFiB
c9blkN9bZqFQ66YVAHSIddoMB6L4FrKdzaqLYY6CuDMQgnPJD+6cY7HTK2ZkDM6W
5bpwbOGKRXU9HDey6l65DY5Z3IfepsvQZI0mRLKsD0n2X/IRAFcsFGSw3cPV2UVk
wdZsNCgHwVFrPB6ZrTjTiQzgPwcgTdyhx8oTSDVWigfgcEEvADMXE2VTRZnAGhHS
wQC/jCoBc4dD7aY93J8Qj5vsCkI97SzJjQCIQ5Iy52a0UFMKmWEhFyoukeTn/htZ
KdWo4TQelGLRMY5ObOJ3AyNBjkvSM3ZRczoBXUT6s4fq/o+eDV5yZdD4pA+zGfr/
zX1HnrGf4mxM3BWn/bdpYESaGb0e/v+iRiXofuWqbA6GO6OsIIESt0OocjGVYysJ
dabI+7y8MnYOFm99NY7Zd7jwBMijVFupaT0upMPqqCXe7mUSYIRBIEaWRWf/Swx/
YX5k+S7MuUL9YDzX13QDmsfisjmny5ick9S3qsZzzL9abobahv9c6UapQ3t58iZU
NRkRknLVZX2IBy5w6yKbJ2MaaRD9sfQ836JLC8nAZ7oIpRYyMMdhMLL4QDfs/Sn3
1WsNjX+qh3k128WXISFYreEdgZb3VKbqOw8KHNul3D3feEVNfkdsZdS9X7x7CIdF
oZdsllb2lGd5I+BjEPYfSUtIcGgZ7kJOXu4dkixdT1kev1TLam90fvGnm8pS1u+V
cZANMrtEDyA9UoqgPO1UsPgaR6+JnW3eEXVP9f7bUFyUBeMT0dRn9xt4g9zHs8rM
88NCE0UzlXccGFmuog3yf1sT72K9jBraGoIHA8jtrwue/xtr5WhmD1MFtC2tKI4f
tSera/v9tkfkyp1iRbGkgH+krAASRKLCeptuDk+HMJvvxihGlUulhXvowRQVUfA6
EQBnfo/4uCvMsHNuBbTZzvS8ypf8H1XlchV3AqScj+aNePj3LP/T7jPx/GP7MDhm
+4X2YXjDQQI2FJW6ubssKSwH7hkGJqhX1ChPu+XkROK7CKkdg3D7Bl0BJdn8gStV
wDmeskmHhfNyI5k41E+3U07a/y3AuIEcoot29Hcfuk/kJVnZqUCgbakTsvNQvTwr
4Nl7pPZhTVtI8II9q3dWl3WiR6yk93j8aFF6wpBJLRW6EOQ2QDTQd/MIZouMFHM0
dtz5zNAfgaTA8ZKjS+Qfs2VriuBw96/0lb3EWmjBEiKyzZFvhXu8WGAzga+ixzli
JPbWvdelZrOA8xl9Sj25HzC+SlCfeUUwpw7S6eQsHAYhI6B/1TeB26sOijC+c7FF
rlbNDSDMsbY0ipQZg86J1LDg2C5T4cNwHh2Zp0shJ52UnmBxXjV7Py/k0yMsuBnA
5cqHgaTv918MjT0eAKm2ejNThpoqEgbtr5oBtWNDFwVdP60UDRohtgTYtA1x90bF
FL32a4jCTjdeP/8s+DaRUA90kQKeCOOywJI2ZxZlDkM8BrcfubYMybnklO0YfuNo
ZUukqcppoJRLtMsxe4mNrjaiVQBS6xfOK6z7dlmPQ4ZPyMAstMh69+MZ/HzqQIs6
hwXFT6en+eTHCuGxYfuN6IRnJdZj2mEe/++h6CPoeyzVEet7U0k596Dxv3uxqXpW
zXSSsRgBQRwohXdLr4iTqnJ20DLUWqeEm4zdvBlCyfDy61YaTi7AtgVmYp6R5IMq
BPMRYq3xObiQAOCW0JR7J1zgaXKeB0HGpzm6Hh0bBbN/UgrdVJG9qWkgTiS1dvMd
RIBF/5d2LqR+7m0kEZvLuOmN9S4/bHaSd715hc4EJj38xN+rNH37opkcLLeKsNUe
0yuYzj+ia2BnsD2fTHHtp8H3C2yz4skAG4MaUzXA96oYJNmcuJuWJDbtlFI4fZpd
tj89EhjDHShzmxo+XAH5FOw1sYEaUMYv0xbDjsu3PLl36uRWfvMwuhgTkhtZtP9l
x1fNfxojaPRNlMVK7qN6XSvTix7bLLTx5RZbO0SlG3uG5sr5wyVHw+6YJXLWWa3n
PWZdQAJOnw05YaZgeHAFGcTxqlf/lj4M20ujlnOp9oE1KbgVOzM7Ov1q4po2lmWU
8HpoXGlYH+YqB6s/qzZ+ZHiyeQ5rZ0MZwDe/EuNK5BV4XH6xKnXNxyRNNB6upgs7
zsEO22nEvkZd39ogAd+LaFsS9lMjcJUgRyjFYj1PrIHV+zB+njpIm2/Em55gUrao
npjzi7mBngANhIYSuYM0DUSYiT/tXuOgrpLR2V9bKlt6sJPilc0LNu/7gWkz7Bau
YL7gaQqfeYK5+5IGmA/XxeNZc6Ye243g2Hu4PlsuTfnLKbO4GNhMxrqu4Ohb1+dn
+z9B/Bu+qHeg3knWW0UQKCU376L0S8bdSSHDa+VZuULFdsmdVD8jbnWHXtcieRem
JkiW/X94sUDyYGTw2SZFAz8XB12tnYVQ1juiMThAc++E10Fvm/26h9ivIT1+SwFF
8gXCwoY+B0yWFrDHEKrYtsS8OgankdHlyk+1X2gAcCH/eA0HOIO9wIy2P9DHmM4o
GCaG9YW0kvwd6/Bd/YbMx9opk4l4wNP4l8CA2XPYPDQYjeETDDlAF5cpEeN/ZX5+
sbYxr2hpwKnslBlNUy1p/wFd0PcF+GTVYIvFe5wdaJVSs1nn/B+xDD24rhlMZyIn
drk2UL4R7/24zu+DbEmYbxwKc5+XGpv35Z1RVxupbfKR51jTgs9MdmrQySCfRFn9
ztcYQigkNvhOckv5RSEGT/3xqduaGc2JVTp37w/oyohZ2+twCwTv5/kfHqwKraDi
GZ/Mdzsm0iMa9ZwOhc5/pE2EkwnoL0NDorVvFUEJQIn6NwiAL4vHDwxKpFSaQINy
mZ87uUH00rxrE+6hmKOS/JnNieeqmcqkYAnXvnI47GG7hpajq4OByTAtbRlGXdru
d6rxvvfruyjWXMXnGGOPGnBULkqaoQeBdBV8Ip7MdlEpsHwXjV4QeMF8roj8uMZf
L5c3p11Jj5eakH/DBpKouhcO5g8BHCnGOyiNVAnv2edJ5I7K+vUE16HyWVRqZyPr
zw8Y1TKOV0KxWBUcQMIQWecRRz/jPIYh5TdFfus0AQGFIOl+nsleEeC9wpeDqgpZ
HQJ2hXHYZKVcKBoLcDj9T/V1AG7Uu339VuVcI9TbZasSrXgcCB7y9zGmbrhXoAr7
klPlspl5HemmR1v/hne6UF3tra94rQcdtILqajjcrf7i0/sR4Dmid7fEkeBMX6DE
IvEIG4lR7K5YWrZd0T8LMnxXDAgbpaJ8mh1qn2b6uoXVvC81774D0jJjrCBxZmU7
iRPeyJ/+1/dvSZvveg0VFs8SowjUEAuE3CA0lJDmJp3RW1bH4F1Lnb+122w3jTfD
PcSXQTfCqan3G8YEp8hL7etxNtZ6Dzea3GWEPvf3XnSZ8RhLXcP+6LcdPEr9XLk2
8RdHmrGlZeKDlWBzS4TjrtINOlMhpIEX/znECGtnPcvJiyQefSGQ7gYdKbFW2gy5
fFRW/61ypbTRqxpbSDhf5VXfQ5RwAGk2rlzUwLC0XGCmkeCbyITHoHsUcI7U07bV
phZjAKAVhx7q4Rws5B7sC2rupWdGioeNL+aZsGPpJWUhtF8qdrMMaTeL2jy3xlPo
P47aqH4e7gzb1NAdsZ+xjX3Ii2ZrdKx5NSSgpnhfq/FF+skU8nvjS7b6eHedkPyV
u0uVXHgkMneSVFSINnxNEO+J3rTZaJ9jPd0gp7PsV5cJoW+g71MDS6q+FJRFFE+x
XJz3Fdx0b9MSexDe7XnbLcqGir5N74SXsteFOz9VVV/Oh04QPPuLwNFYWXHYbv3K
u9gDql3PCBeQG1E16aEUqN476UiUy6FQdzAT26DcqM2Erm4+Z2QH54/wYCFnrqkM
I0+oOP0aAwe4keZPlbZFJm3ezkO//DiZ4YFE9uwa41uRzUVT9HbRv+Dx8sDhuwsd
wTEwAcvNN/gwNk55hegv0VUenitEUsosybrqtZWbCMz+Je+NZPNvSeBe9FbT+u11
oFSPx4Flj9/jAVuaOTutIdiWGJXeARV53eiA4/0bH+JjSFC4rKFR70udzBxquqCn
/AmJBiJwuqEVh8wICxkW1rDpnUqt3i1zINr6xrr762jl524TyVfKvUWo7OzpzgSR
gMuPGt1cwbPmEmNCIAMyl3/GeaM4DbqdlKYuBvcZb9hXJfCAXBKyBBVDpmXUOZGI
Fn0yb/VRffHFZmY2xus4PCnwHp39At1WXLxOtLmgi8lRsU8ypqP32ehvK6Xj4ciQ
EnYeGV5JxNFakVR5abpajR5kVFmu+q1iEd5F+v+4JTpQcAdXExhDck9zxBa1aeGP
FnkeRelTptO8kGATO3kGGSqzxLTk9Gk85RHnDp+8ADjjCbHX0gGEcZ+Ymo9jGxy7
IcuvoZ6OaxLguY9qPVervX5FIVxF3Wc+towHbaOQekhm1tEisP8ax39ci//iFECy
REiQ/8NQzFD8YQ7I+uwwH0ywRbR4CpS7zHwzBjTfSfHwEnXXl1TZtv0RR5igMtrx
PmAazXCQBKHhvbJj97xXU5+T30wQ/UXuMMKuJKsHo+0KxpCoXvBF49Akl6Muo5TC
iNaeZc9H078Tvo5+I3cRUdG2Y49qGEbNxomCg6SHTCNdrs5MPjzK50bjcEiqhZYQ
H1jUF1NYpcxncell4YDqZ3xkFzjpqEP1I3OGWHPya8PiAELlfmRa78A15N9WqDSX
hDF1Y8koUME6qJt+MlLtFDEMNVTX3Gysj+yh2RjpStpwiQh/Cr7SM5vvoyyc65fV
GLlQZiNIW3fKNiozzSlJa/aOduqj8B3aKgl+6bytXwUNWPgHxEZFKHFiCIGiNzAh
6s/C4uMWTfvUlhrjAGa+DSKUpu9TpwJ2Nt0Flo3nXQ7pwnVzu8Xke8MdU7MK/2dU
xQPfGXu3leCzi+QLTvuGQrT/2J2SP26PKGqHWWFu1cdMs4cyghOj3Tfzbve4Ak7I
lwR6JmfU2pGLKsCwBB8B9uniWDH6cAkc6ph0DwAESt/EFPr8F50loEyLjG8/tLh6
aMUi+7fqa2sKt4jbbDatjGzpLqIXtiWIO+5aV0zpU6AOp0T1wQCJMgct2psdQiuL
7coMpiVYwxZZZNHg355PV6Qc05wZKYiY86YYlnuMCHLZ/M6fV5pShJaJ7P646SJt
tQZLkCFdC7iq12zMLL5dkN1DxzC/1ZxpxFB75NXqWO8vBnyDUXKB5xYbjVSxMzCI
AkbOlYogDr/iGpTuXKAJhd56C+4LOjMZTlazYaUY5KGuptqjUFdYw3xD7LuP2Tn0
GYBuBfFTsQhCmfBKD5YI7nwbcCyvgBoas4iGsMn85lETzaGMVBqbdAO8NGsg/Mm2
6K0+yNmNy+Z9Y9Xi9VkE/qhhEXWMnXTqAzwCNz4d03XW9ITVJMoJB44YiRUUrZvJ
PoSbjF77aiUpFiEJu4YBxKZrX5nEFet3eVEW95S0J2X0bV0J1Oc1ebARwAS9HKDl
BTV4zh3d7qd9lWX9rTJjWw8XW+CwcO0SWJG8W6Q/nudNVxrMRp1yZT4HcEDZta/u
YvaKD6xL2VWyxK6aGoK4vpBcPaIwH2Bufx/bGNKOjamsKnoEG/odiSnqhe15s1zh
QedWPtGnRr4P6tKjS6Y4jDaIRYDMB9E0BfmL6qjvgnovlLCtY78eCb+31YZ7M/tu
Fj1KB6KASZQC3J4hE7FIose0Zf0MrE9/7QTqew8Sjff/HpWQGB1XUx4jVVeQhw4C
VqA8ooq32okGU/vZFoGW33CH1TF0X4yHlT5Mf7+PLkwBOS4udM+O9BfmgPU/5xwN
yepLYL2zNz9r8s8FmXvpw3TjfCbe0r73FzM1jWtZLsR00aniC5JqhblEMEroZDDD
O+mxbSxtGwnbMbr1HMY4EzQjisD00vK2U74+ZEILH2KAcfn6epm0KUxwxFmpTaJ1
lEVsztT3u52BNyTMbnQ+aEfH3X9am+vYdc+dm0/xU2jm7NmYUSgfvFJjqsUqUygM
0XS0zd55FM5wcJBPQzTdhIaTViggLSlJ2iob26CqclFY52Mik8w77xxBEKQV+9jy
IyRb5b32VIfltTDFPzGmRAuYCA+C/qJHGe/So0PZRTwoj0yX7C8+nahYW/8CXS5E
5TQmdlRbFU/vngILMkJ5hRA711yXbgu2C0plnaYDX20sJdX3VMd3R6w7YJJcBIKB
2Csa2XMapJViiykeMApvJWTqYdbR26ULb9CXjZ2NaoyLEvwmCBs66iUtbTjG8Fip
AglqYVeAGTxCvWvoWIXO1r9Hwm2q0QR0ACOx1BGwhobUHP8E29+WMWWjkqQ0AbXK
06YdxMxRSnuiSBOfgWQhThg1u/HHsPOWXcyRgILnUxD0RCsd2RU+tERysIZoEz7V
M//DrmCRPxhe0o2nx+6hvFQymrxjcpPsh4e7TiMXBKd4BGkSjNgWDF3FZ6h7pZ44
qyMQUyc2QGpkHJos8MK0xIp6xZl2DkacffoLECcXlPdKLqgQHQ7F+bhnuwUCYs+r
Eqz2q65TTEPjMqzPdSQ9bUS4mc5jEHTw43WryPR1dXNnaxCER2Rqz1aeHt9gS895
HZFxNWuYNd/kMPsr/z07R3TccrKK9g4HGJH3S4HUsH/3NuBOPTuRLc4dZ5CjCgD/
x1yicvSmcBq2Ppv3JT/8UnbbXH+Ll/9EavRVFsoxJFeahSQxLFi8qJZO3I/CjfQF
9SR3QjIg9rcpqP/IvMtSWekibFUFBDwvxEgNfcIamgR6jGwdEf2nL9CKnxYWzHKn
JQZvsdCmPsE04tS/YpMmPl6XyETjrcVDJp2KBeEvsldJdbWHd0uRjtiMi0qKek/s
N5oo7RPnkzYAkLzW1PKIOQErUeyyq6xGD5iSlEr2D1cwMLlJfdD09QU+NtzMVtC7
pKNLYI26zC+kzejhl7P7+EFVf3lB/Ofhdi2Fw/lqmnbtB2lNfMjH1M59cXB5XIOV
nJwOItV5Ln9Lh5WAYdII3w4RprgIb4Jb9tkZDQu2SLepwB1X53lSHisPOuN3gVj9
STFmlksn6fGLKekSIFbh6B9Xwi3qINh8H6LGk3wQSMdY8xFZlHMdeK1VS8aqAy7C
9+ptCWuFzJUdQigiqicWDgMuKoO/71lCD5NZLSYWsUP+A5Oc46ScLX9ExlO6KC1e
P6i4bDRP6fiSJDQ2Fat0ELNuh4QIcGnRB+1EG/K645BYiNEa97yJpBAOBgDHvCJa
GMdsc5jCiE+Nxw7WDb4kgvJhYWXBqPoA+QapiXrVIz81bgdQW4IAWNKcZ86fqJz6
VHonKieLk6tHl3GpRMjCPq9AU6ti8imJO24DxtVv9KrIN3RXBl4lGD4LuOyJKvh+
KapOYEKrhuiafX6qAwDwPIHgFYo35OCG5jNrWkXgb1TPXog3aipNFyiUGVJC9njY
gGlu6TUWcIhJ0rwfIBAnWD+pKQ2nZWCsIxMr5hUiK8E1KTAgXSxl+lISZNspVqyh
hF8gyGZaex8HPIsXJg3quSvhJATpnPunG/16C8QJMGH84V/UnidXSbGR1qYyT39h
uQZqorxVK5PCz64HTRnDkjXV0ZtX5R2Q10ue+t3oFIfeogepfNyR7ACGtfBwP/+J
XYUd0/UoKIxHzMlG7v34i98jtbEIhQpV+5gvzjLqax8AA033eqpxcxW5vM6N6WY/
1DgJ9PJe/uafxgb6UfWLR8mkFfaSXjC3eSTV6qddWiJc0y7zOWaE3jauZofN147f
lALRcCevIrPnJoPbDG7X2xvEsm6DlodyJrFxfRa0dGeRffxDeupul2ea4KWusTLn
q7tiV1ij584AR3O4+KMO+9dhmL6BqavVgtyY8F/JXKX9LYk0wioP6JiGX9SGg3Aw
7GmHaEl212vrMNRJOhZLB+vF7QXTU4vGfYhC6+jViWbgUiigt0w25KFUxee1LBYK
ruQFtlGxXVcncLP+YnjtKNytTLm1/m0dXvFQ2gMi6kGSJYyHCTRVXhIpTzVtyfMb
u706eoh0qhZICcqgQlutPtoos3YE/8J2NHPgPqX/ZR3ebBPpUGW1xO8HYjWjlUUB
l6YVDAAbgzPbkSVK+Knr0nn0e766xKWchdiaF7lfa9SmPYgviFVF+AxMEiFIyT/z
+MkbltGss8MmhEl3cRdAtkl6vhxta93RwXu9EvHcnb1x8zZRVwjMwhE/Ydn84xsw
OQd4rWLWDOVSO6WVDyoic8KeH94j1n0ZdmI51iznv/9B3q0STaYsoFyAW3x/43z9
ByAv2RK9/a8zJ6y8PbOn6u1Gbh68XMW38Av7G/2k/BpX5MNjnMYaORxL2OPbxy2G
Qysij+bacQCC8hL4osUhhIjDYegB2y74Ay6tkGlZM2hwh6wh2o8Q9MI7z+fdYNaN
ytntBVwejHYUEmWWwCtEj7aQU7ZKIkUgszB/60jSpIOYC6gZbNqaW8ouRkI6oQIU
Q0sr9ZZa1Jv8PThJcAH9DVpxKQseTLWhJlu3mhzOttzO9rgLWa2jbptC8Cq3IHJB
eQcA/fQmrsZWAXRG8tMCpRAIqQgidTAp+8dJtGAt5vkzpYY4ypWHZJCpP2f7nDUj
TnJAZat7Ulv2cuczPcfayZKcjAh/3cXU/OmI9zVkWjZ2TuvWVXtGcsLBeuWaLjGk
HpSoD7iccO7E7Ox73PM65o2cJTBtQ/r1vO5QQZPCm5yXZLtoyU8SSp1hkaJoFIb3
q3Vbu68oaSXGdeQ/aRNu+7/yeymqKk7bJbtYk9VbD474LdD8YNwv4SWcP63EVS4w
tdYtzyeJfOoLPu5BVh6F3USNbBlbrcLipzmJEKwVt5GgH7ghVdNkRjBktF1zXFnT
GPYD3f0EdiCsA9vkew8cnk62CQc0yWgUXff+OFrdtBUTtnCADbSFTQBEV+4sBDR1
GT7UUyflLI7PeJvrg5QuYTi0m1zAiypz7yboctzyVnCryppVWoLYPURGnmQar2Gk
dIJxUr+C9XRJlaRsweKBjWKrpNwxVy64GAxZUG/BqyS0qxZtPQBNoIj3aWu1GbOR
1hCRG7kiB6DHfIBs0782eNoN+eG/yHxnflrvjW8kvioQ7LPBXSi2h7jHyk943RAA
sbDqIqSUkY8sNEh8iN6ua7OXYWuhbWDc4VJmlmg4ttGpI8/pWdQGEcZ14kAWwpnm
rMPzJWmHYs9JhIcxBW01vEiiUqvfpk3+CGrtV/nBSjhjEo4geC0OYWaLz3WBBzZZ
DCArUJTnXjdkvzYHx1/gheSkHt2J5uHqZCW+N6ylNoS2+W7MU9uM6FA6RQUyRt8N
SwDpy1GGWkXo5G7NUxxOyUc+7UbBxJZ8WYPM8CyIFFdauULjmnvuP/IP9JdtjYM7
8mS9CYh7muLej+lYQyKytlm92R0qgP6hAvFa5k4fHwxX5o4nBrhoW8ODiiQwOD5m
oMdKbgFJPGy+ZPAvVHZSHE8V+XqG5istyeRhqzL/XzM+TGjaEq2CnFR+MyF1qXgB
80z6skuj6JjIODkQQipVTJDFv1TeJHT8i0rxS7V/556aGhNBaecG7KMLEoSq5x0z
Xn9jSd5n+lbpMXq3MVigjURo+x8Ib97pWXvqGkcbZlgp9UkhqzrloWZS1Dd4PYAT
C0MQYrWTvkrq7G769Ew61w94zE1ykhFBgBUyZKxpS9Y1PFes/X//Wd/JMvx/j2Eh
KppOxTZAPKkb9O20FWo9hZMdAL/2jqIz4e/2pYLK+jD6/0GJVZ1ApVLrQoPim93N
oi0Gp1CUrcvT3QQMhS8ZsFvA2pX6EPVeNiTlCA3pcTgd/7HDh5lworfFkMuyiaU1
N+8IneTZxYn0VCpmb1UaBJJR/oHK1OqTs7hvnrBxnDca3QTZlmb5ptRfi1ANzt+5
nVeiBkIk8PZzSIRwhoFgn+OJhNjQ0E7fNAYSeK7xm7WTzSYslOQdNAzy0vHdM0+f
pxM7YC1YqFRPOADoJVlYH1mq5GEkmpbb0yUOChc9b1fbZr8WvueOONF6eQT525NJ
1HzxEoIYUWPqnQdzDC2YHCvbXwAVTz7fNrTz3WMSm8FQYYmjz96kVQ5XovQ6gphL
wF1cClPAqGIIp9jJwSEPA52a4t72APM60MOsaeleFkjQksOEuH+wHA2KdigpTPKV
1R+9HdEWFPbG3nzibgJR6V6qh+K8aFGqhOBKDUDkXc1ofuyxmd/MsmVkZLLHALLP
5PDfUvXVi0+yif+Nq/dMf+m/jyD9cf9J+ZVbCSedAnQJaZ36pHkhyFU/fP6dN4QV
Bid195+IseBS9q39SVcJc1i7PAnvsys/xrt14DeNouJrbXsj2nRnUkeN0IVxR+dZ
56EV3QakD6HYfMOaMUV1ODlyoZ+jtDqalh0ofGNkx4cX4oH3rCMi/eFKkklNGYAs
9tEpIS0Vrw/OyMR3aQru7q2pSWYwvHYh/SPGj8r5/Z+ksQ0PLni+6IGTMZPec6Nd
IFgFx2WJUda64o9UvmOqBpldypzbwvaSN7CKx0sc90J/GFZewq/xXqiq6txgaONy
AroE5ySnRYk45R3hAqlAhQXFTprjvqPI/0YXcnBHAUtCxwR6RZNweZOefCsvX1ZX
+49hgUevXwUSBNIpWNPkbI7VBVHeDmKO3jOvFTPvBZAJEdGPHqrgYMeILvK3EkXe
QZhbZ1Qa7/Cwqg4usPTnPCgJqfagTDdCHnRoQHuIdQFpA+6YACvw0c5Q/a6M74DF
528OQRzPSchDjqX1AXSBPmc6x48WYrgacIqQaEeiuEq90MpfaaeKsao5pcK7qP9N
Ih00wNTbqKHkqRrNHKsQCehl6/rTEEorgErCHXr2Zn2haxoZfn7LrYoMEvJZUzrl
78Goovnw3hzEM8DJ46S8teh9GuXy1KkfH570aW8sRMDWd9l1lVfWZaBNZ94yD881
q4jGuk06y5rXmzGCKJ9ID7f89WDZYKZpgZBuDF62xOvzJVHJcx4TdFWFXkfTL2BU
Mat/qCIdsvIWZu55eqYlJ9XGmZwFWDAXoRqVJRWgUVsiZ2DVUtMRwuTJLLjmwk5y
+h/qMY+KaUbFbC2cjNJld12ymt+zUJID1nOhHFFkSR+QS7eRwpUo9hN+e14Sl9PV
iVRokYpQO8XIn7T+KQ7Iz9gG/5p+m8GXFtAri8cNT0Au81lY0tKkA2rkuG/rzmIg
NQuv1KcARnN54lasGYsNMUbSYKJSeaJqORGCbA1mSpOXljqYQ4HVdeOND5+9gV6C
5blALJdTtpWPNhRZRBbRlgNoefN1qAF0KZIyAtTt/EjxteZBAeF4Vq1RFTmoAzpE
HtEzsnF1Uww/dD7xDomxU5LOX9FBW9kuAOLLELI6vSQzrpuzPaMJDyiYjlaaua7M
+kyH/llj/39lwUjQdV6vxnJWCmiS0gGLklenpLASYgiSTkTsUYYxlF1/FzcT7RyZ
zG4RLn+ssVlsYlJTDjQYJO+G1uvWh4E55jwEIuOIOKkgcOPveC64D3pdIZwnmtvs
VW3doMj9rCTpthEtaYpKBtL2ennpSEujfidLfDiO11ocBz5R9mXrfSq/Za9X/pXw
/RiSJLrEvbYcMI39HEEKuv10KmvypzoHPFCrXlxsEe3FEEwyFJlKoazFWnL9ZszO
ZZ/FeFEaR61FvDmbqx1QvZI/nw1nP3LB2/g3CrCMxyl7wQyofKhh5hZdDrhaTvpg
Cwqo0NFzy2H3qqNkfMo0S/DxXp6bj0LHErZAlwO9RTPTrJxt2M/Hi/2q1BdngmbE
VCLs7euqk2VdB6ZFbwf58AQGYMEdrPrzQ4EhrA+W7hEbYI5KZ4hi895vM1kEvz7U
CLRsRvfwbVoLRKYGKEqTJnyDoSP3Xvem+GS0F8waaWfYYsbr0neGkExJoAZZ0M3/
tPgNyMVIlnQ2vTLDMqIWKslWm636IUEZZIYS/2RvEk33e576sztjKU7b9dYQuf1l
EAzoaHMsc/oXB2xTMtkdtfPUZuX9Xz5DRTY/qGcYC+FZuzgPiV3JR8MCOe6rlLmj
vH/6CvHtFJVvo3LDL3sDlw1uTLwowiYwLKcMZ+6x+dlKukJMHbBqcE28Ng1QyvzB
SI1ypZAK1oLeQWOh0kL1nSfPromQSdvDhNvWSI1s273iMPV9v8spv276ACeRagDd
+yVNSiKinpoz4HMiPRypW/bgo4hGR1q6QjfKIWf6p9oNpqZb9cUpb6xgVjvhQJhc
zqpE++pxhFCEeH6jvWcQgGIMzr12QqrcIvJPV3EVKEM+ZhdGFKsH6iPeuzPj2HM/
kzvxcmaVblr5VOLdNzgtUL2Dr+EbUaUfBszgb/1xT/M4Y5ECCgj+MwEwgUqqsjZm
Vzmmdl5xHdDbytLKSKAPbj4g7nIO0rMoSXEGEd8F1Llk9DkNdlvehjoQXh5wdSkq
AGZzujYQXF4StPB0Ig7VdnK9ThM6SrsKdNhlrFmXEquQg3086/yAc4mPY8vlg1fq
aJlx/Misaiuo0yaChafKjNZO4wsd5cPJ48U23HTbZO5alkbquYluYeOoGZveBXhY
/inbbD941lZCbk9Ukhce5+mt0gdqNvkNQhI7ExWiVhOaii2rddascaD4G6efbW40
ts9sKjbls1aF7ZIovFrntbz2d55MkotkwHMrJOJQen1yUhRIEQ4cW9xo6HCa8NJb
o0lzlco8YDYYGMsQUIX3RHHzZ8FFh/pziJSkzUzhLaNQW924PXtcaUB0jmQc9n55
44yacBE6NddF7pOEn1e+YVOmnmSIaFe42WaRuoq3wm07vTLykl6WuXnsOtgaLxuC
ZpU0WNI/beJbwapqoxvaKtE0+NTxR2xY70rx9j2mP52piOkQeYlyb4idXBDdqA2p
sKJwsphiQP8wPOTUD9WNGBaC3qCiEFUL4Mv0paWTpirpK8ldjMSvQutx1H53X5Sh
1IabjeFZ420Rts9/b8ZczaDj1W/pBh+hJCvsXbTCujjMKfmc2m2tCBSZGwZ8yor1
7GBiBzI1U5Y9l6yT9LP7zE9nW0sdTEO0UA5MQAlrFfkeczAvhGN43eW+Nt4QZsqZ
9MQTvVVt4rertT8jtUwU6412xDCUobTDVxCRkukjp0WNfhw6e2puph+k0cWbdX/6
+bQ6CSN+ex8Qc10mw5BLctjlyZYai3D+4FzZUBbArwXTURhLB8yabv25J9FMGNIc
c2z4LAz18zqaeFQv4rHqEQTPWt1cL9d94SHyPWdjC8awfLcHR9I1+p01Hne/IW59
KJFXabgzw/RqhCssS8DURyGf/ERyInP7NOE5DZdpOllHRb8HEN2/rAGsYjNEBFaw
rIHcmO9uI+ToL7gG4eGv/P8kJBCW6AbkD9eGtgyrsupWr4vnpcHx0xgzNHwqmbuY
/nnMCv7XVlPpx8gEtmzMGLZomN7P2A5QUed07u5ySlFfJilIwKf5Rge+L0MQKGsu
xjPQtqIAts3D4PuXXWG5D5y85uzUBuF9381Pk/bClrkxIrcaWKa2wT/+yf0P1toZ
eYaJVIb4hMaPBc9J12+KHDOmoKUVsPVcZNZQfB7I3/K05Xf5I7y5VK7v6kBT4XF0
UbO7CMMc1PheCSah5RTy9p5H/rHUn9X4TXGuS1/AztnGkrwV+7g8cNzx8H1fuByn
QwDtbvmbVsQRNiHlIfahwhOOgY5cMCiL+Hvn3L/RC+ZAIXRSxuOfxz8SOBOzQcN/
zZQOCMv9rAErS2LVEVLV1JIipqZ//2a0NBuAcg/2mG+OkFyfFVsyJyn6SeJzbFjV
7oCgI/6sP4v+tfPu57BlUHk4MEEtDOR1MPjjQ8fGnVg53rCqGdD7PVKJePXmS7e4
oX64vmH7plHECG7FiQFT6YrQ5Q6aqWd+soVtKvAzQr5O4HeUJJ4dek4PRP4V5V2S
q7Ygc3c8CtiJwMLg0GA+aZglojq5hMjPgzuiTi0EpuhF/moRBg5zT8WxN2hJW58o
+6AFa1A29Eeuyt7yWC709cYF3wALxar+eXnGe5dtB+bhKI0jy8GSsAnBcdE+ixy2
aA0TKARU6vuLy2nXLRsB6KJUZw//1dlgVU26ukaLyzqWbVDIFDHQW/uMhmklumzj
HZqJVV95vUTH6zMH4Lucsr7LNow4+waMKHUF8NZjcd5cXxIqqDoxQ4mZ+kcu6UFj
w6DFA6S+URfZssWGEeATKg1pPLfq0vnlIlwdFvXr5WySHLB00ezPMvDchJAcJq06
YxFZFj1um0EQoFz8w2xOOrvcrinK+6wtRNKG7PozTqrFKqV5M8GrlRRFGr42tMjh
olso/rlcR/CN0JSVYHmf6shD3s9iHy/Ai+Ahi+Vv8BExHzFH6rhDWI0OuexH+HJo
RYkSGH+K9V8KFvYZd7EXuVCJ7kE5S1xgvVjp7hjCo0hyMCz+ZdJffIiNslOeSJO1
kiPp5xirSd/6/WcjjLtdZzPD0dSFg9cCTY2J8PiI5rPpppLgOVavnRBYQrgkPQi8
ws+qncIcx94uT16wjj1lWKQaw3Ryy5NIefYbnWwzD8ipZVQQq3B24OnxHVkF03NX
I0uMX2KVMqM4XbtcPaqI7N70MA4CrOh+2OYJ90qhZ4SNFOIVHVW5f51rEiIOJbBK
m5pgXlpq3kH+yTyEv5bUFmilIZqqZM00LTsqCaF1gy5PdRjAjK9C7SOKOv+vBHfz
vRTLo8Q9bpBwIb3uTCJHEuBlPxCmoxJhpH7CB4u9rBf08SEH019jacX06jgE0Oze
5aWt16BEeogpQ2GZqyifUwp8sn+arJSbpH3/nVcSU1lhlQMDwVAKmeTwQ/TCBHir
6/u8X4H78ZF6xOQZE0yY4EXB5M8WkvAJtH99mUX2KK4kQzCnJTPsM++v1dFHBr5K
Ui6UUVmvVjYhK6Qcl/7pdgbRH44P4qPBtslrLb46Xn3eWe0agjqIegSy/fr0/s43
cf99V9LEyBJ+ijCgCW4pFEoBsRyLuhCA8c0d1HJMFSyWA18Smbc2VHStyLZVNPQ4
7kx1c7lpiQ58Rf0qrUeRGSnDRYCmuBMdsSzlAANmWtcD/0KYviGm0l9nGMQvJWGP
0gRDpoyINDD6P203ddJ7oclQQQYB6ZfVvOvvyc+7g4Q1mDlSXygn0+5+FB7yeMLN
4tupqnu5kBn7xAZT/Tw7c5f7QYejNe7lStftmhdz50RzQhozpCAuspoPdKKvmece
ZLUM48WMiWIqeQqLyEm/QGCRk4R3ly0b5H5qZxmgcKOaODMsqtQ+yin5lZvrn17K
rF60s581hziOXpMzHVFt9Tlx7ToqGL0rJZOyzk+Q1bbMvWIk8cgphAT7Vleoi3+V
tJjFelK4KQ76vG3xjAhVAirBDfqEKzwIXk/7Kxbd1Id9hVl2Ce27wXzjGOZf+XzO
4YtHBBFzfSqsocxO+LVPlBCFOxlEtNVi3P7I65Me+wod21nVtBws3mGQ6m6XnpXz
sy/tt7mBvGrt4qqCZ5zQR4WnXfuEaX94zYvlMZyJUNG5ASTgN0p1dn8y9HewG0lx
IvdrI9cb73Rz+wJSDI78A4cHCWMJetHYgLiCPwwFZD7DRyhTyaXMqlAv/NN2R5jL
BGhaGINXSSyjwWZkj4NamWqg5CjvORg2R1f+7VV1kU7weycMGCswEUGNdqoNwEak
VHb0LOYdWLk4o89q5M0g6QvxMzrCrWuPJaEGfLZkjqev78s2F/R1p5E/Pdm6nfde
Mprlxsjo+CnGMITC9YMhYCe4sy/7N4SrC75QEnI63F7Tr0Z7tc6MJeN78SA7NiVa
b1rTQcR+8bB55dQMrvCYJvDAA5hHHaiBJVLJve+TVC4S4hkfC5B+Osf9t3SNls1+
e3XwoNI/qDffaeaje7ciQZmU7tJ3u+1H4i7qYoiWphiKRsL9y5a08PUPyAHJAF9r
5s7UtufGQOaci8qJPr6i3NHEzY2mOwgTT8xH6LPrytuZQp1d5iab9uwGU7Ams59j
0jhN0k7TCNA0MdWFtRd/r7ce8Q1n9qhgW0wDSXbxXcY8oeuEP/XBTsx5b5w3wZZY
WvfN/I/5VoBfkYKy9JI5Us5LTNa92VsFCLWhIa0fCBwScNwhHaVFJ9wYR9INIOCX
EzGWRA5K7hyjkQCj9X0XmU8q8dnWplVePOMW/W3XBGnVa4p2bAHY2GkVFDc4HD1Q
MXa9/wwL9y6A/CjhHdJy1mVNyhG5/K473aIQ9ZpxmEa/nT02b8Ye/VjKCw8+tijw
2GOP9EDRM2WXASA2FfaSi1lIUTFXbgO5TP9Vd6r4dlBUpH/+rdHNgfkTodV5guoh
Cl2Vh/LFarVBWqfc2gArqa7OA7UQvmiimtVlHCnFrY6iGX/BLo1I86A/gRp6956x
BOM/03/hH7mdCJIzdmIgdcLT2FMVMWIqX83ZwISx+1LcS6RK6/8G/f3hByBQ2xoy
6gEeFvXn6CCFEfHksEq3J0igNQ0QJ0patNJRDKvlMUBriaylLFv1/ykQCoNtqzZz
tm9xmyCseXBJktMoCbk1ixuy2IOZJt85oYTcubpmi40wkCyxPH6jzmGMXsaZdwGI
O0fOsLUPvRwmZAD5VDr8KFZ1UNEn3+ltWsmUEfqdAL5sFcq8UOsYvwT7ANTfG+iu
XYI9/1Jnm2Y6JBp6x71YqTj9vGX1I4J0YCMiSizx+Ld6AnGIOJ0ozwIZFq1w9L74
RzRWKE3WlxGKu5Pk73KNnoxFxp2FXzuJD2OnxgFNWacWIaI/F8HWwEFGYX3AJOFM
H0Fc2ibolTawpCS1XCWIOw4nKxsmc1TuAsHqAGN4grTOqqD56FY11aIcrvD5IJIU
Y+uhQjgNBWWiAStDRsgvvdmgsdYAnyrHV0iALXqVCQO/JS/YRradtk5ooU6y2thh
5FTmS6Ucq8cYujC6L2eXC1l94HNGVwWYNbXLBAawjDu/QXHWSn4lEFUemm+5ZutN
r0UTbPZGDPKSRX3Cx3UEbLxhsbQ3C3rRy3UGAeRFtHE0nrYRvmcGLiOOmhS6vwyJ
9CDYE4r8QwbRGe6EXjWDG8xoYNkyrPZ1Tz8h0g/NG/SVrtYnXR72CJfYyxaEvEk2
Zz3Hg83ty5qx9gywC9GwU1lQSxSZ7qhuc5nPHV7YQuFPueEqzpyu5FrtD5TZbuJv
YfTbi5olFsLm1EuU7YFC5nv+2aKx1LzYZUFwLcYKjxz7YdoOM/ezlAGyGKGOJ1aL
MAX0ypokhcmj3n5XVqZ/ZC/WuK8Ch2RIj6pYNIknnJMNGmu9vhrPkHIgY34CeEdv
61ujK9FX35xeeXvydOTTwDYccypR6FZpI2I1yp813gD2rohu6Kf5WoyOmVA3SHOA
Pp9bv+qQufknyEKKjB+mv1L8Cqwm408o8q4OZ4KX2+Nll07GQ/73MkMJsCnflr/+
GaEE4ZuJ62OPGWwr5OniDQgOcaAr3mNIF14+Td52hdZqjsgOVe1bYImHUwwC5cyv
bO4nPEGt074cUTmndzx3rRFlOJLrJ8L9CONDqJ+RDtYU1pA0NxKXpZfBUSfjowMD
ecfSz6ROBLzlEilBkS+iE07sUP8Ih2ukNEVQ6Mjh8IrpMAcvyFQCuFekGIidJR81
So2v0Sikp2w4zThoR0lq9Uo+S5Vd6fA5KnOfyyzZ4IH7ibvtHz7XNo+M3iAT0P1Z
dL0Xm3IanjTF2cE7D6NBz0Bw14rTCBdINYZx4YDpF1B9z5gdWDsLjpCg3ly4QWbc
T6Xd8mOmL/HkoRhN76I9olnSb3M6LTHrX7TrNIZxyhLkxncNpH/oJ8EdqX44z39U
uFnum6YBbCYS5Uot7GymvsTkYL9dpgoHqrWO1kZ+z9YKH9Mp+f6G+uYzQNNRCzI5
nEnwAtCu/ppHUW3Gt99DYFqY7S8sRxY8zTsePSAJgnZDlqRs0D6ro/AiCPODA389
z8Svnyu5VcRjxanrdhHFksVHuCpMP60L9SiJ0MHb3RInOQ1qg3hN3SGTlMXDYqdi
QBXc0+dGYDeNsEBzzFkdq3PRCqkuflN2QzV78bVqUVzoqSXds8mUoYeYwgI1gsQQ
IJAnu4FblgSGD9/waNVF2i+4sfVW6pzwm+iYPPtEjmy3gDoGVTShDQ390LKc8C4B
J1UtsuOtQgE3pmVhWYKPjHeVsqIAZpDHwPv5ykvEKO0z93xHRh9k5CZUiLdrA2b2
Bfc9fTPc41vAPYcitS7k/BvvNXf8pEEjWOSqStXmIpfHDCpijEMLGnRqvUUQAJoi
5SZVsTreTtT1e4UEevuqbjHMGkDk4hl5ZTwXr0hBX+dpUxrCn3fu13l9Jqe3XwsM
itqXAROGxsYkXrZcwlrdCpvacPEV/d0RVzZQh+2zTL2Umb62uw74EkpA6ysepko5
oDjTperLo27GM3HAVHw/FyHJMsMFMU0WhH5yQD9MCU6uth3EDdQ2nb/krJkfoSK2
XhFhrZapEDDsBe9GCtVuyhNE7DbqQ+3TQbGkBgRVVyTJSfsQRrNfsbS1YNNYEvP/
iEAnSoltrcCxPBryX/SqJ0HvgQcvrqwsUIbZUf4f2eq1tSV+f/zrRfSlejJpxXGd
vSd/arZSZj7eO5utyXofhpBil8T1z61T/DktGS8bRv5YQak+J4IfIaHY9ufE42bS
Y+7MbR912CR1/dvJwsZAvhUtMuHQeHzM3zqYA2JRLBoJrfjYQZ4mEh2J2dSYkHjs
UAC7f6yih/TJYzwAgvghd8XA57xcjAknhcnbAFKTsYa0IrMXtSAjtR/cwkJzfF4q
O8LMq8Ayng3qvPyxypeVKFE84Ur63jr+ZJrXr6XdJYaRfQtHcDkDhEMIXGkgC2RM
xghcxPSh9ef4FN0J/68pmyf5/xm9W8mqTPSVQt98dq+ht/6dUaRz3eK1C1LbUQnu
JMV58iVCxamwggYT+LaI6e1ORxMJnK9gNwUO7kmIOvLrIzZrwWU4LBrhAm48vC3j
MLs6NQtiwf3V1zL5Kod8OBAOoxxKvMLebG0e8nyxTPYGH8mq2S7qVsKaEqhzXdW9
vwhShnkFyKsjIQICSRVcPaRQ+X60dq5pqr3aVi9Clyq0NMMJmiUXatq5SwTcoB4L
4KP9LjtPxoziCHpaOlC7Qq6z/7Oi5wTL70YwfnVact9y751KTiQdRrrOHYMhO6C6
xMIhIfj7nmDO4laXioGnhdu1MrFOm542fGYfWYisgiBiPoTtpjQU/6FzMezdzgxy
bpMZUWigx5YqU5XrBfItTVWqQ6LoF+xUimDGYoJUSkT8msV9Emo4q5johXuQ0rWx
rlE7W4VwnXXFusgJFKp0NqM4n2gobNryxB1GaKLWeyNYWqISJW9ukow5SiBArNMb
fWaAdaEE0gU3vyP1jkLT7zmg6LCvMrpX3nH3cC+5/6BKfAceB0jAYO59TauyQPA0
9lkjXkKF4pW/CwsUpl4RO4qKPmtq3i36PXb3myQoO1S75PvDu0j/Z8rbr7A69iB8
WnuyZjaVCNqHkVUbzTmabiQzK2O2ZUMc18kyhV0m79UAt1AsgtYnNucZUpGlCyeY
OCFwYTSIdWGMLKcj/lwNUh0sECSSj8TB0wjyjuffOJp2DPF17p4OIZiFNlRwQsN0
RESCH6i6vWSaEYF0JDkT4lcplt+WXLX3sYvjGpaa3mjJVUmTwTZerLncWbEILWT4
vOVSct7R9wUEh3LeRHsLTCVIjVZDZmJbdin+6ub4K3mDWPrAe6QEFdMX61Wd1x9T
P6g4Z98/yYVoqeULPXYCtWqaRMgVFFdn1dYjOOrn1hMmEJiTFjBO+WvfD6NH+QYv
CTywvAHxg+oysnsggwB+R0rMEjptwBHYtV0Ms4sPPtW12wvKhX7+kOrEs++//7iM
Ci9blOFc9TlgGzepMaBaM/AjvP+ckHBzZjnO4hAOnPkBMfGOfag/YnFS0IueRY7f
JJ5Dtnl9Yld6TCtQ+TSM3lMmDpzLwWfngkZCh86xeHOCQxIy96P9MlsF/Q98hgf5
fZukpq9InjpgjbNbNhGm6CX9th8otEHTlTTXapac2VOsiL20fNWVb1MSjiXve3cP
3/rn1R7bJKBFtz5AI5+ZS0qFhxK0RIcLmGN5i00cQZyPwzXSzwsRCLMWOlQ8GCCD
YLI3WQ/1LHRGdY4qQCQdX2Pc9YyVdZZtUMybWrXylrzB3KZHeoPqglUuJ75lDc4l
Q1kjgrpzIcwsDM30QcqVDVDuanP6rTVFFgwI4AbU4hY19o8WMFXfBtCw2qLECy/g
XSYRICSiBipGhyH1olOwj/KjsE0JhPqPMYLr0xO2gemmkpCb6ivOTZwJReIolB+b
f2fRS7FzlypmAXFwvzIBryFTy3wn6J9eECdk/Ld0TXECGvEDwgwwoSokRtQtr0/2
UqpQ3KfP4WJqLDo3pcWtX5QZGidX9mgtC9tkmo7Hz/VMaZWFYMb3or37p1nwj+s4
AAEVArAAbetrgdkLPvWz8aIWtHWRPCXPVrmYmyyHNy6tdUaUMQvGEH/rv4xgicQU
ao9fhH2GtiFFVJH6BHGoFvIcbCA1jHsrMuKv+w9A4om+0157jpFegUMBChPFZFit
HiiBNMmZDZaRtG+LIndEWApGL2MMVD9ApDEdYxnONSIwkaBwWCqS9NMRwVmywHl9
+GXSz1eAWZVTCiNz0naYbb2SbCbnNqtGVYT+VV4NEvjkuCvtzCd4XrRq4Nm8FohU
fNs8sr3wD8LAj0NHyfStDh7W2NyCxsudfyUdJuKTTL2MpWaVXV+J8oPNOvUG6Lm9
6SgwIXbKLAHRowZf8V2TDbCqEjC4T7QT8yLemuymGgojcaKS+dwE9KG7qcvEq/Kp
A6x9vhIT+PAd5VTCHNKyOFP8y7C2GhC/1HZafIbFYOp7edms5nW3NYNKdkx2STEr
m0jRedc+0gbAD2BLfOmDOCJZCkjQpr9WpegOn1A8BxPBxT4mhDahtkU11vQyF9L1
ZMtn3U9nFRpyQdPZcRSK1QBh7OfRP/FWQOLhaLqJ8FdBn6NffV/OUTGZW7jW4RJY
9DF5dpENi7evWEOkZPjHwAA1JtHzkGY630OTHWgaCPo8XmcPeQGkAppV/GoD+q8A
pTIuf4M0pq7Mw4CjjfXebb1JjwlcEamI2K3McGHDUCsrJcj+AThW7CdkUPgCbq4+
d8GAj7OqKVBziPhpyk0YKV2BkaOqHTwEFf9EKvCHeTWOyk67eUl995jFtu+XjJFj
xYyMxJ3wgowBYGzYsess9pa1YRh9x6xdxONQcBsMzchiHIDzcWz4H6WWut5Hd+0W
prDvuDOR+6kWGrcFytc4Mj77k8JymKLWg0oAtrk8QKo7aloeL0qVOgwtgl1UdRxU
5isdOOM0bPPqm/UGNnHYvnIwNS5/P9KuOD/2cbqLZSgpS+IJmY00vp2vL6xr3wTY
k0T2HlxZoyd9mdAVlEUuRgQ1F7nNJiPeM3rVN8tP5DtBkp0no+SUA6Uq9LOtrcIT
UMNVKRY8axFU+YFReSk88A0R9/Cbyb9/yh5mGB5u50mQzX2EmkufdxqNA5MXe6aJ
5dgsPUYo8DHshQxq2ajN857vhxrXJyN2oSaJ7eSYALEpIyQ3F1bQ88KG9WTznSmN
bOoWolIotax6EEm4LENta0lFjutnhJltsHtYvaiFGKXtJNc9wDlQI18edDJirreZ
ID+t8wmzL/JnNviq+FqdLi6sW9X9hMbHzw9oaJU4E2AGH/CU9ZOw/J2o66/n9pYk
hUao584RjA9tKha07JDL4zA7vS3EYeao7gfPnpMg0bw06Cs+6E4J5Tkfh/KKqDmd
wHnVSveQR5w6Mtw59goNyBQHUGCdOo3XmMVKtA3VSH0aYNIr9pD40epEQSwJoWmd
1Cl+D+/5TvpQgVMZ+NXVWWDWo3jKAUV6df/skbP69SeGMFnHiFq6hDjgGE6UslXD
1HR2uldDl3mmI+I5W/+w0xThx0Gq9ju50qB2miKrRu0vtaY2/mQHu3Fy+WmdaqY1
VAOu/IgcPFI+6UVMf3nYTKp6oNWCLnWu1dGAi+1uuUdey5VFBR3M3H4pRu0xznAb
nGRYmFsn1ExBUJerLhhlwwTWg2xeL8F1FT20JI2iUOd/V2GrXeC4AsdsXLip8Lgx
ddcc5IgDJ1ke19Ic4/zCRLi79y78TLgATARETcnrBrrscSBHXR07lpLAUlSHkCDv
bJMn4wB12t6PHBmHq4G0vv8Bb+vCwDxdL8qw2LdQUDb6cnNcmdKVqh8sKRGRrESR
LeyJkpy/pWuR4TzKnTxr5tLDmNzsLN5kH1vyh3PmtmO/rwaSzLwXp1eE0bX0Ajh8
QLMjLFsvF48a1OgJy/ZOGoaRvm2/HXDbf0e1ovvOnKB6wl/pUaRMN3Ro66Fhj96C
JebB/vCeQC4oU3epbsRWgRiVoKhgE0ScSG/CU9d17iMvFaviyFNXbbVd+7ZwckJ9
5g3UFJAuDc0Cwho4d69N53h1olVlYQBIejMYBRAH6B9pOpLZ1M09OBDdB6D3CBpT
WZSoUJKBeGbXCkPIutpdyfcX7zafW302SqdvchqIsWfzAsmRFg0R6N98Li7yLmhu
IdMxLI0e9vrLUUYVCYD3NQcWPnjI1LpmsI7SPzot8jNiGh6sOnvhu4JdUUFzSEdP
4OKhWCUfbRGZsYoQhkTa7No7Nnzd7w89cAnLuO9h/Q+i5dfT8fJWHFQjJX4xgbTR
vbe9Yvz001x+iovBczRxjkFolZnDc13m3KU751GrN42Rn3mP+xPChSAzTMuuP4KE
lBbEdC/KWk+WB9Za0piVGEc3KHA2QI/mOv+PGAiBcla/+3G74SywSXSfVZibKojV
S/yMD37VJfjFiiyPsBGCyPA7X3M0TgPu1OLoyV7LdaXwu/BIywT3t5umFR8gcPYH
ghOplxws33DhoEopl87ZDTMU0ET4ZVlizhsc5q5cSu41KDSFaIjg9WR+cUNXeWfZ
ZMyY6R9uG+K3wFjdtSI5uG2LkZH6cHx0W4IOvyZvI6OqkDw5bx+Ej6whC7O23FeR
cNUWOsX/TDQA4fiobFwH9TEkExRWpM0sodwr5FpIWPS+PO8dmlAwurtQUGWu0Bne
FLmadEJYYPRF0GCfDQ2JBGIoW76MdQQfe/bZQgI1M2dhFvaZOJdFGjV4vFak8fAK
TwtyaX13j4Vtex5Xr0dgioaSFqNQ40UpXrc8BiBfh85iKBCe20oGcYgTY5nluBZS
gAmsx9k3Xz4XVaUTe23uY81bY8RRAtlW++mvwdDz8pthsWq63ls+fK10R0MkWuea
f+JBE88WKA7k1Z6s9MY1a6Ox9mVL2/b96vl6uPjEApZd0z2cWKYTpUZqgwk8TUQ0
xN1OyxGfSgIStSqEom3yYDHj9GDXTuNx0v7hevG5BFv/mbtoRd31IOcbXOH2e/bf
5VzF69GgIf/+ye6b3EMxxdxhukHtiSRmHgR12yIvYpLupTUKzhU8Yj78cYChay05
Vyn4nkhpPmJI6IAvTHdY6YC9ozmD8JLDLpPrl/Jf+OIUq5+KbXw3PmVGVRq23+Hf
F/DP7cy9unba/WekdIqA6mgEO3N26PhU+yOOG40h7rGsEvOFkWLWAR0+QYwpn6P9
kosYiooV5Dw9OWWDPuJAbUI6Qremc+ijrWyS3q/vwIC4GZutudgc0LkMvIGUbGZ3
H/3UUsnJVD4kB9yzL0KTHEmNlAjFCNxW9UYLDqyyrxpmXVzB6ONOSeFUD/vvNDf2
TALq+EW3FmMOj3lt2SZMurEity7mTx14SbNEMOV6J10q48KcCssVuMt1Hg3exltw
lJLHLSTE9RSjxAAbyBUVRGnV/90FF7wJGp/efEVFPSzjxND91454qDlpEZzq8TPW
6lY/XWSpWJJB9BaXgX+J1AE/DFadCjr4mV+veo4jE7lIjcvdmEODVTM9x5iIBFRQ
l5Wfb489AznzgJ3QOn7pq+cmWg/QAbWKxJ2Sax4cqADxEvUh0mfhIi6Clhls7Gcc
hGmUZ8Zn2eJVrXWIM5Ni+CVz4fDevgEIQogcC4381Un8SDwHOCSYmwrF63ryLkgS
GzDOATlLS25KAu3Ft34XughHiRpxf0/UCyik2sjEigqlkdGUc04wVyCo0W5EWUDm
aT83qUVGHV1UBMxqhmT447z+TiFVZfn8zW46nveZx65CwIL53/BwSVQasEwSMVGL
yxl3gpf6sTOjYo+VAL79lA/T7KSAgj0J8cSJ/fyPDK/OlMdRqn9qmTfjHMnlf+1P
pD3LeyKNoB0rjP+YONGqJmDWIqnD4APnpg5kwMPdBpmur3LK/iBwlPgqukZRjgOn
NBWPlVhj0Pij7128P1ZLfI1ZloVmXXBrpMoih+k7vd8owBbaibbzDAu2zVxPMbh0
R0brZzzugrXeaJ9Z7XrmyET27LgBXyawBEVaD5FxPyDXU7OSocVaqLd2xm43ly8C
11yb42POijodZk1Ywa2b52c8xdLIJGCsUohHrYlIaX0ZqN+PizadA0BDo46y4wGd
YLbH660tJN1tihLPB45Bxv/0/poMIJPbHlLiY1gMDItz1eqm8G8XtS5gBcFrBqu1
k/+V8AzUDGBWIJIEiDa3rzRdbyeX+NZL+i6SY/BPwklQ1QDGNfFpJ2zNWwygyqnU
tn+6B12WBEJyKE+cglwAwBYIkjlYeDPVRfSonfpRqSSpocVt4q7Z5s8vbmrVnWCD
8Kjb3PYZDAt8+KhbUvpsiQwMWongfkXWCPxg2CpGpTiendh1jYEss2wWh9PUBW/l
Cv/3L1FaXd5slVjgKmqi3kpLftdaNw/JEmIL2IDay81yIRdIFUzhSmqdAkfDbpzc
oC5NE5tqROs8HjOvQBNIdfmfh88/yjITuety3NQAJeMkw79JI9Xhk/46dtL+Q/yN
CUSbST/F9IdwPbUuOdZad1TT39XVQO+nPQM3C4Pf2t3zzGN88TMs4QRPLaO88J8l
vnVAu/Q6SwSEluxRNYcD7k2UgFcMMH34S87QClcAM2xFRAvjH0jiTsyqxGgkmudQ
C9ejZ9Rq5w8A4iDPleps9j9YoLZJfz9p9spXAJWgkDTnZwEJg4KDCKgrLmTYDp4W
At3taauLwY2zvtBwEaOWp5nsZ4v3sYynML8aKtbLDcretoIU1h5+YTvdJnoa2rCS
MnQmpis5KkXQBuPDCiSItNpKDb2SEghtNZghJFlRG14SjGL5vKeo3r2YV4r9lqE1
+Ai38kJNLH/GBsy5gqv+dHOBDsJdwUZFEqsPWBxhoNxmQdFlEpPN3BlckIreQRCb
S9GRfQYjZVxrGQkoMT+J3/egYH83NFXAfUdCj9u6kSjWbMZy4fBbDs52Kv3MkJRe
vR8ZaxGavYQr2hkmGp5jmWY0TocEwI3BY4DlSXiEq1QZcDwER6s4KHUZVXifU3kp
c6hRgtcjLRiulk2biR9YXCcKvk2pkB8y7v69mmgP4U5izn0A91zpYbUPeZl1l7+M
amjkF8BUr389+AGjOhY8Igrxqf/ptWC9qYPcsXxWZFLsHpdWpJEoGg8e6sswAOiW
Fnvd1InHyNgz/yEBItLNtQwNwrX5bxHbYK+3HFyvNL/9pyVFh7cY0XuvZ+U2tixu
mVFn9R2GlccEbO8LOl1FBinMHl+9iEGUhZfgmhsKwRDrT1mm+98p95tYRMnwfL0+
PtDR65Q4/pGUP7WnzcG8qRJJbaxNpubtHl0PFHTLp3WPFwDBcWYpbQXuWQZ+VMxa
A0/nOYlsXJSAoQ0wZJrUpoFnx65OHntShpys/VG4Y1pmsGEdvVY3qpmb1FdgDAit
X0T+kZih43fIwjlplbaJDZw29fu6H58qi/hX62dXOaKijVbRUXXhyXvv7fv7NeOX
PJIQr4uAC5K59tEKCISuMkFMNghT8uwYZkgSGNG0+dkwIrEsJrrp0UPdbmGC0p00
3dJzJNGykd2Kist+JM/6v9/P0QfEJae+by/POEVH7Iqfm4JL9QahBqxDuc+0+Y4x
l0T6gMO1JJRcboDheUGUW/Jx+RkiZ4S6KEQh/ttthJkF6RUVaHg1ujlu6EgRJP4I
PxLGjdpCNbNHELIbocqT5MwKhv9+6A78lebawu2oznmLt2D0UdXxA9XD6IKmT5Jv
ZRWXSyh6FTZgrOjGRe+ix9Ea+p6Gfqv99jSCCCAnaqznS9F4zpc+kAoeYprxJUGZ
lYfg4LmyZysznt0aIdznL7IOiO+GOgqKRJDT8TNos0rZ/lZHjj6USRDRVo0pSOTc
76efsPo8egvNIs9IuYpgv5VPu8l6ljehbqycBnygTE8g/8yUKH0ntiIKgB4bICTJ
OlrkbGUnWmoh+oPJGtW7NVkyMYqzQlKbPGY/gOB3UENTnkBCYwF7kvZTV0zWy0yM
ybdT579Ow3L7WkNe2nx3setEnOrjtjslLHckPOB/DhrHctLcfVltnWE3NDoumkh7
BJ0XQ2bkNqwLdRRcQtRjm1GP3fzhDWNXY2Sbyp//Cf6Y2Fh6ulkMphvQHCVhEaCp
WFSR7bWG5LFFcBZJn8EJH2dR/99+omy8MtoFUlaZA0SKpL14OqZCMn03NI7P8NO5
6oSoWT6ytR5+EpqFNrSyp6++kevbKon+ynZ/V8a6ziiG7PkzqbqqnM3zwV959okx
ivC03dU+58arJ0jXoDGPs5KnPJ/2Gf13dwahv7wTW1rtEFVEvROndvMhKv8r/N3y
vnrAcZVpqPgyWcoBpLihjoWvPBFvLBWfkA9llG/q2SNyUmWrGUEywD2vvk7bgI3D
eESq31LtDyaYKHO05PjPpFvIGbOLlINnGLugwGDB17+hBFQYh9L9h2qTloUYuv3n
TCw3/1aNg2gpuc4tij0HSSvRAG7NtJU5crukY3z93zqpxv79E1HgbalQFqkvDArb
fGe0EQgKWLVftT9HUqJOYH2u4oFegrLODVOBZd2sjVL4D3qQrdBjdKrfixt3JUSH
98cb0RKkKrA+A8P+dg/hmMmwu4Rp74DtjbqyiWErTXdosdc4OHyTyR24xILgRnfv
v7XrZpmqmYA0wYq02be70fXm6TTDKRVUB3RapO00i6MuVoaq3d0bjKW/sFHmotOZ
B+Z0bjJE8TsU9j5+U9OMHjTp6AeWY2ZMf3y7WA8SGNj0Q4ztua1CRdkE/b6bYGbn
UUv5A6eyTanxFwl41naPRIzHfuqpWQsHDJGcEkYqR9wSKXa+Hw7st7ItMljBWoRX
BmG/7ZQLZ7o04tBBb2QK8kI+A9l6v0yP8TLinZhronlFZXpD4HBCu3cVzraWPqRb
Uef+YMOspdimU11CdyTn0Wr7HqWzBMemeh96j3omwqcjvDZRutcGbTbxzR/4gj9Y
rIFSl+cgHVK/lM7+WZh+WHANqLMbYIfTeya60SBakGMX8ORKmup4Lywrx7YwoUq2
BuaCZm2fQFxmkzQ/JB+J/wt6Acpr/zsOlU1JT0QbsWHw3N1guyAAXV24YSdaLAP+
Z+BTHPrRR+mvHJnf7K6bTGJskIyqzGn9HQkGdm0mosw1GZTkV5yDJbNo60YAe6bJ
q6K0/UE+KcW6Tu1/9ct0VZnmGPDqjCFj4eBi/OYKn+fPB6EXDDAuReHg76uhLb2V
TTeY5RX3PqVU/sx5Mg8McdLs4ToHm1MAfwMwKoe8/e2/JSEJBGMSvGmdweJEyyMh
mqcTCKOUuInpBt5Jpxvgb5wbMY8HzS4iJ8y4ut5neJBTMz7PC4An5JFTnSetmaqH
2FXBp82ZATjjsJ9KI15c0H8VDqXCLj7cGFXbksBWO9VjJcvKxMjaDf4e+JX0p72i
hHSKx7coMQQ056vMQu49nnLpmKjw2x44IehbCxgvFN7y0lRbCqoOAT+pHQW14gpI
p+5lMzquXrTGyoQZk4R5/F2RErXDdnLLwhhlccjJ3CQGgcQR7CGDwpEblD7SGC8J
4805YUcm+hB8c76GijNtmdwjcXSCGUXTNPk60FGq+OCbigYfTIcLFPWZJ/recEXz
SAhOiUmHeTmz6z8FoAHLWFmp2ieYhXV89Ps8U8ZwYAcnQS0FmrWo1vzCv5wFkgoY
FxkpdSiHzn8dSSKzRECPbOCQ9L/L+BFH7SxIxl/YfzhfBrLUL5Rmw6YpT8UJ0AXW
DBzl6MEpvPGSnielQhTJdv1O1eC7Shk15IJXvgTgPfU745d59ETPMOs/uJKq5Qxv
/JgDUEavyUzDNiDRcytXwXoPjffJlvKlIwCUpf1kfEbGx9LVbr5PLqYXowcXEhjE
dRKtsaue8WAe8w7HjX5XOG/IR+2UapzUBNYojWqxTjS6zeENSIuNYmPGpKhjb4GC
deczJUS8sDU3901+KBf0tZVdr6+hnb+npf/Fbyr1ilf+eKkvpC1cw7efQmBlX4M9
OfYXbS6DL57VteBxmU3iAP485ASQiACH+vzlINdiep8CUW6k4kjJ0U02m7G3h9JI
QeCJD+zsZmauaEQ7FMIdvE+gr6L5ElqrvNQTSJ/WBN9RuXZstd6SDWx5xI6g3u6y
gN5f2adYVpb1uYcj5Gl/k44JBVdXBg0yd4Mmo4JVqZWxn9pf11VKfwsiF3saoQBn
wiqPm3Gv/cHVGJu/IWpUdOq2RvTw/JhUs1sefhEgUmCqWmjyR1UVBlkitHbyNnTT
klyuXCgfBXMDO3xnXgtHampD3SL/BTImz95GZyi0IF2crAoqmezlwVFZ+8qpAHGI
1TQThTq6bw24C9ALeLqgoDMXnfmlU3rXEXOQsmvpQrMgPTEoTAxVJRj3UifW5RYQ
5C+8ZWk7xPJctZr4yksmryxFCjITTkTEA4PK6TNg3MtE4+18Xcor6JhUqPjxq0Wl
CP8wa5vf8FBaHitGZxsFrYCxDri127oHdj9/Kg3PQFN9y3vAYmjH4SSPYM4029qh
urBGfS3E1nFALoZsiefJEyT4v6T5TVD8cXXu8Zvo6up2iBti+CxCZrIfXv2fUqjD
o4+8qfE6i3rgvRf29OpOJ3EJU+6p9e/k2RlybIck/tcIYQjmWP4v1Usw9sufPvTS
RJ8VqeHGM6IF26ByGq4T7+5NSb5Fe/oXNUdD3Hr6GDLq17YP7CG2VAu8YMZMtJHi
g8QEmRU2UicKydTSf5e1wbb3v8RHqIvL3QdUJFbpGjIDMpNht3qDi0hdldYtMPIm
7LME9oWHfUNVN2T/lNEsPLNV3c1RYQO88ExWFzdSa5YNRH8cKNiBvWYB7ROa4LZ6
lzF4ukJX347IG7bWCsAf3yVZU1ejT7/1NNSHOGi1rJ70XFyTeePJelYZN9q38ygJ
C4Wrp3rXtrtI9+lTJZ/xOc4kjlnjuM65OaOw1244xroV0Ogjp/m9RdiVlKOdojBH
/shYH6y+6XpPldxE+QP9/7r+cFrDoGhrob/J9tLqbpteIsdCG4R94WMKgW6R+0f0
AH7qVW0dXV0AW2bP42G5ogyGEAGmt/9vvAY54OftlM3zXrHDvBiSsLhUv7ivObgI
DTlxSByeRjhWNHcMiVdPvRSuiWES1FroJv54K2y5z7NbUstdLDutV0JwLwpEMqhT
M/rH+EUsuzW2X9T/WXYIrafadeXuL5m1nom0nf1BnIKfZUEucQweKPElUa3cVJbJ
mvj9FNxRfHtTox3R69X4qortkQlLPDt9rmYbpUUKAPBdfZrQ6G+U1ykAZWpv20/S
O+7UG5QZ6hwWdMiodO+ExLY/icbhRJo4LoEADXCviTGTPxmEIbGYvZSVND1i1pjx
ejIiKoNX5aKj4188E5d/LC43MwkTvOph7kN09wg8NbzO1OstVD0xn93yzHUwsobY
vXJ7Kj+B7n8CorDunsnXXoaiNFRUR2drViPkTOJKhpFNiqDcbshQlUNuOaVZS2hU
dSVYeQr6onNTMmXffgskMhChe2SbVRZF7q6ePNZR82kc83D2q9Zt5UNooNEQE7Oj
fEck+BHhS+m3v5nZATrM8QNUCdato/vfmd75sui9L2xZTZlrW1dV8JMaI0t9Q0ad
8pFwcmA8DxOLaNKGkUDpLxBi3/88mUCJP/OqrypDUgLFPAqDigqSmJcJdlTcnSzk
oFfm1QmuLKsMBPXDVlJWy2NfPKx82wrhiZ2Xn37WcR5Ypc2zBMVolA8fXvKwbeWZ
+J6KH1kBqeKvqTk0m8lNPJW2pReopFc4Wtb9JOmyYcFRq5ngVxytNOKSBrXk8xjS
JmG5RWbta4eVdZpiQlzpGulsLjAnq9acBLM4sVwvLj6Wc8josLN45PIFsXhFj+9f
hzW3X5vo/bY+0dpaJUSPcxPZAB0tocNNUeyxBu91Mi1xr5/8a19yDWmiXUhByii6
bMQQa3jTlXeeS4IgcYVpS+NXvWegYYaWREIhnTmSzbuC9yV1PoiXeTgD/WYMqe61
11UhutyUMaoT4vB3KZzKe9l9mUI/G+yDd7AQ1dSNBCcPj5RFCsXm4NjLV+ShkTYK
XHB8PD0bUEUvaFFFJowSnqiqbAKtDBYtLIP2EseEQp00lcnDje40qD7mL9U7wsCQ
hh6wUl3PDLrfB3SOd6V2cDSQ/Fv0CijkcBMifxyTdJxTmdOXfpsAkEi6IzR0aKu2
SoeqzcQvjRQriiaPyqGxHTOiOCk0fWObQt2JEkD5m2kClVHI0lkNaJDg/dmk41vJ
l0NHF2nEFlRoyRhmZxRSlKOMaqvQtEdChSH7Ufsjkx0KaqdhR8BAMGPRWC1AhpQw
Jt6jA6qewgGpEqoIbtzwFXYnsKnustioNp+pIiflNK6XSfi3y8tUkUBYdJq1GMyO
DceMU4x2IrjkLDlI2RY06MdwhRR/b/lkV0Yaa87tMPEn4StSgViIs0nUJkwqIpPH
c/9QZkIrTithpqnXa6+Rs+yLAIjn/Ja9L7uPYy8+4sZdsiiUPycZsbtWqVEFGcpa
BEVpVuk89oJX/fje0mhA7aQod2ZM6rW5/++rv1CrqQ6uEtZb7kt+NqdCwOo21yL8
JdPZgvwT1CL7Dgky1meRvpdBgcobgr/I+BLZyWRVBBn7TGSEeFlctJe6Ue1yzgmY
famtHafQ1uNiIiorZ4+jgvJATzqI/hgzhWTJMauv+3OeowQ/SlxinHmAWTtINcsy
ISqt58pV5fRmD5wk5SYJb3MJlde62cCUFqtvf6ekVrp6FyO/wpuKN84zHL2XU4+p
FlqLesyQREnjOlzMebaKlE8JMdt17PLA23yL6r52VsXf/YoBgyPDl/ewnnjk8gxA
6IuiWj1knJZ11vAJ/C717byXTTR0v3g/9HyFuEeYkmlA+wN2jVDkVcU8lyNY8N3f
xwdwRyKeMrSG1HEKTw8Q1f1CQ/IUR8GP03OyPF3d9y1OgGMuDSQoeTKNrC6yGu8r
EoxU3aQpngZHSeGAv7sIWiVPVG8kWBEDLg5aHfBQv2am0UQ9rmPdRPZHFY9pZLgB
k4EjuGvl1h4ygB2MbHGOmRPBBb9A7c6/rBxoo78IWv41QH8BLBFnvV494d9bjV2u
DMXuzkL7Nfx/gZhQKBJ9t5dmIRCrpAEuqr4QvUVX/o2zbeiTAKprPWSQ20J6/W8H
nR/dmJ2xW/H7r07A0oXCwMdtN25gRAbVDz9HtAON5fCpl1ACGHAsZxTf9/8RdMKR
+jdp00JCo1YoqI0G7CEcgbUsy5Kftaj8izMihhKozuYTPRUWVOxuvsHuKF4p0dip
0a8mmF7xOCfq0t80SN0uPPen0al/nA9GrYBfalIVcKkZUtSrHdFwvbIbUs5J353X
2r1udE3jbtlo9swwhnVyaQyZj3/QibCL07mv34nvw7G1NSJputv8c+LOENQbJSMz
Fvj6g1zVOSwyXw1UvlFzORGgtR+iy2dpf04GA/vZCGx29XAlPKNCHOJ44gyMXzaa
soKOpApnDVVI9jh+7V8fIGRZXH8x/NAt4vuEFOmnVR+q/PuoMT+JWc64AdCH1fNc
LIgUx7Z8ujuQArubDh/ZQj145n5FFztQa6FZw3+XUInaylfXimilVHEWzZVhTtxY
+fvQBzRh1JJzlCMBTrCFMvzPgfyzEo23YfUpo6zW0P2CCJkmCk1kqB08JzxdDeCQ
TgFGx8XSxIb7eo0c04WXMNsOnzS0KdX+EKM6nbhpnld6Zofm4m9i7p4/C1M6EVVe
YvD4RBC+95YNWi7EYMH5IiQxyXop9YQqKoql2xWVH7r/aUNh5U2d2pgeReuqTn2X
FG3xYCnwBmjnym8hOvudv+P9t4OpOVb1DIZ1uJ8QKhZtpVnstnHUXaUJcy7IJEg5
J8fJKu0c1DLqw3ZOKlHnuNKhuzrq2QODP1NYDFMOuFGRkigaxeBqmE1cisSiEek2
4pMTN8mOYgvDCa53RynEwsBU/2uNwj6sbSpiW3C1twPQ0gDDG1iPiuLfGsaQ7ggt
8rtbH94xW1xl2xhBjmolXAC+OcUjkPL6dsvG5bJSkLxmIeDkM4cm9f02QqrXGIln
Wxj3fFM/JU3XNl3f1biqAK8gRHBI68QJPa3KwYc1YiERED9ti2qjxJWTcI4Mm4HO
jCnWBGAibQCwmlanec/t/JWqZbKtVCLxJ1A4c7H/nf8KRMsZl/zrNErQt0fDSPZg
ATswlcNZVPinwU/OiLt+zRCLlWI5HoOYAZ5STB/VOxD8qWc4sJOAQjTu69j1rDOs
eAHUGM33lw1U4yH8Z0hblMnaY4riyr1RWG9g9zl1RiqePCbh5Wb7tIn2YNIBZUzZ
3jA/VA72nG8vS/4bZfWUq86Y5I41o2No3+faCMTU/lFz1qIoTUBqt2vKqpCcZUcj
eit0pCS/Trd565cYzinxMfzasv4hqWuN9nE1XymVdd7r+C9uWv34cSgYzZMed3DQ
sPHT3usUgGDqSVXFFx5/1Z8HIdx+7GxcDvUat8s5gwtGoVbYsq78fQIyPmlT2jNB
wJgZO3+Nod4SOS+3zSZv+zITVKDdETvMcbiakSbZFRGQcGslxPVz2ATMHw7KGA1W
ZovsshracbZh0ZXrQB8uAQsKerbZaX6pZnUrvFj8E8VBO+4wfgWB1zY4pp5f1aT+
JjKHEY3bQgnIbcgbu5wAkrlespSnSqxskFCduv0eD26yoNdpiuG0ibYIXUZ3pJzy
38uF247oEhblrvypFdxLAP4F8MbElSLA6SVBzRVrCxTbjsyqwC3NgvNzHZ1b8k3y
m7hB2cmZhZk+VaoGaiqbi+tPSwUtMo8rfIRVcZy/d2FXIli4uJS9tNw7OC3hN9mI
7x1adveRF0j4aWhL7yIXxaigmeSt7RjheWBjvUyLAcx/nz7iNkKl0Iw4W1px+aOO
BYcL8D4HdupQArtabUiTMwLwcdcQ4wDzxHKSKVuKBeSVx+e6U0Fz2kL1eF57fB/0
CSQfeh1k2j4ZFGAxTbsNiMf3IaJvlu2P2H+zUdWZbtiCqNAxRioW0tI5EeWXNkPo
FNpSUMPD6lsFc1Ix1DKaU5SB1v14gWTl5RxzH5BS4LiMb8Nrju4EOV3R/8LitV/K
tlr1z8cHc9Y2LbQhwIRA/I0vf6elpiYDFeBqO+PACmlGFk837schFzeLMqaWjaRt
XDrGSg/4XrrUmZ5BpYu1xZY3CaqpQYpmlMwNfPvVkIdfdsvtKtgvkYrE1qC1gg2D
Wry3R3rXnBO4xPTfnBnHdY+MLMkP/BwfgkGMU7nfU8fLMW+BJFkeKRKY8JQ+KPUV
wG7e+Bn20S1aTRbpcjD6oy/TgXivont4lzrKowmGhH5WxM5VkccQQLEJKccUBpgZ
IHjTIeJdHZTbOpQidxr78sMBkl7bLFgjhK10AgCTHr8CEfCxaz5ScV48zJISdnkp
8AGRUvuF1OQA9Ln4GCxhxqRmI0l1xp7KOxpQJPa9BAV6AVOtE74hx0MtHt87KkfO
nVCVWh2h4ZnhmMYrgejG/5C0bG+ws50E/Jd0jzCh3E+iXgO7btvmb4hGHvUoVG3N
bk/uM7/BNtCdhFO36Yz/0Bev0XyC3vG9ZuF891wbpM/491IztLLB/8dJX7kIFNFD
qgHPb7ZntvwG9uaZR9Bk9ad/CwUYRuY3CzdciEVqzovzogpWNknICprSLUXRI9Gz
76/OwplybN4MQvZMWU2R3s17qEXmXBKsqWtGWsYNFJDYoHwRFTfGCSvo54B9hasP
rYP+WfAphsx1OetUDqUsPWNaodEDnVJUa7A3I1XODhJ0BM6g+IttgG5a4tl80Tia
7I/ThHYOfeMrzAk07Mlt823vGwq8s6SVtbODHLzG0ZACzVBqm/Vb8Cxg/d3N83ml
DRQR2/4Ob1e4KaYZFUoSmYMbE591iC8kPWhDSwcc8eJxQuJXhVCDKU4cf3NlunWp
Nl4tKbcGW/myLdDBzEWySOgljPHQMLb8G2DhUeKyHvmlCp2QlG+3+C5W+WotgqiB
Aotlv8WIhkavSBvUPwUnWatHTRgGwN7lVVadepzeKl+3DKIxo/rlCeI48BPqXNbG
hxUJNSNa62bZXEF0IGBQHiGx3qmWkS7UvGhoP0XCDHltXw+j3ENHNrxdTyombb4u
iUmdp8r00STsZcQL7MmAr069FEtftOq0WaWrmP0J5dznezNNnMmGfEzfddQaaPM0
t6yNHNMEk2lgKegHzyV6ieE2iEUTgA6/lbOwJpXmTDY8ZTZoiUiKw2K5MrHQrqlA
HwvDqVDhwUdsnROHxfajzygenW4xdNQatX4ns87Z3my1yjxcnqKnXCxgiUAq4kBH
FCWKntXooTFywCQaL4PBTXkWe+zK5AuYbKfASbrHhcXiv9ofAQz4FQvFSMNyYOcq
5Ay6sIEnrxQXKzdN1rDvVo2pTKPyTSFO5hsPA2QfkFSRmrhFtPVv+P2JV0e8GOKS
GwvAJ9LvKACtPE2neosE5QfZNaepP+6J6oplO5+MUp2F0ud4zYxxToMcfr/KZxHf
McnBMzXuvOjOIBgYzur19YDVIEOW5xZQyzYbirUI8dPzrMCg3UushJ7rYtpKltwx
s2MIwpLSC9DwPFrcBwvbCvuBLH8yS0etoYLy1fPn9qzfxai88xnEkct1zI9+OXxf
zF2moKKJMeqKqk/gJamJJ1A8H3VcMkEcIRZi0rgroi/QgtSLNoirFjVg4LLFfmWO
/FyPX5dP2iDRDvkh7GC8uvUR51hObjpctjMI8KtilMBCMw9nGMe7U1kBIA6qw9Yg
YGzj4yq+sZXv9RoPBW37H70wCsDitb5VmmwvPZHbGgjPNIuyHHEURTBjVwmqIn5+
iKgY9fAepwSuPDr/bT9s+OBmYPQFCaY7JYt3hfme9jewrbitj4YJ8BpgbEKsMfeu
Fhzkf0/52UQBHsYe/28/2qD26wE69WTLo2LhsAzrOjt6z5+TSjp6hq2nCerhh+u5
7AzggJ6vSpEvq+1P5Wt6kSvxcsasHXb7IT6tPErvZNOHJB0dWl2bpIWp9Ns2VLTN
jd/FJrX8oFTuSsc6uMWdbS6tWpG3Bd7Lu2fC6HEgm6MUog++AmqRE4kLd8kgF5ya
D5eGXwArnli0cZ0RHgN6T86LFtHotO2nWaj8KRIQYjRP5Pa/1Or9j4+QYcLjSxJB
c2XXiX4Ne6qpEPByXd7EIL5u74CAqCM0AN8FzX/BQINDz8McKnM4wk44XlKV7bXL
qxvnvTdAAyz1Ye+tl5O8Krt7sJDZ+cTf4cOhi60jBpbYaGYWIUs5ONcuFp1S57rX
2+B43JjwdyvuN94BFOXZajBeKkVQixidUAFc5R0EsUv4BHBTrsZn6VNNLaeoTzYd
qW+4r9koVfunE5nDk5zyOq1+VJmXP9wGT3+gLyYuylkxUJRcrLIJ+UJG97j6ucb4
y2+Qmh3T1E02JS7vnugSCn2h5J+69ClTDafsHTexb6ly2PbL1bCStgGAREdvU43B
rjeGHNb7Qbn9DCWUd60oPnxLYQ7l9tEoPR3l0EPUedDM6Y+Q3WZ0yXL6f2CyZ3Ax
JPTc8C6eu+xYZKF+LcV90ZaIHGe5oZtxbmuM+VIaIpvfnD1RlaJpmwRm+VVCvkeb
VhLR9kHUvjr2CXrjxSHUnPBoYq4bShFdtprHWvsrL6Lpgq4Zmps7CpuAYvQ00srl
BZpDXNGM2nfJz9vzGolW7JERhkN9PJc/9km8hYFkDrHcaH4k/Z7vb13K4WIeIlBb
KPZ3DqWxvN5ymkiIYMOqkSviDN/qEohoEQL/3aWpglrU/fX0NSJJjp4KeJmvI+LD
PPOPMc3JObeCcm0Y4i1UF69Fuczglu7bWDJ6vVjkR43IF6Y1nmbvvHLUdiAsw/+K
vUhE2VsbPwQksVYBIMAEz+CcT9lYTWaueoGrBBrtNJYCNYvvzC8cUTfAx+ZRetRT
EW+U8oJsdpsWdBsMfMzFb451R6GUSuWEx/F8U4R21wRkLaNNrMs+ndF7jxHvRf+q
G9++eDDZjLURxUuS2BDPmSMUmukoVOYDGXfP82ZqfMx2ZXvZszopJSrwqmrntedp
BowJGqrCWB7v+jFN4nvCY1CkPHCQ/dJ4Rg94reprXrsqDkEfNtwHfLfCHkj+aAqW
4X0FQwbzUNm1UR+e05C87fZa7eXzHCXXQlaJF4AU+D62KWihAvOkdyPBj+eI4zPQ
U2ooX6hsDVoDmSV392rYExan4qrbKSKPUTq+h6iCWrqm10O+2rcf2wsVxkhRmMd3
dedkCETyhqzK83/UUWIEIhMPvVvwr6rgXM7TSVSx+Y051M2K7K9XRjM0xKk3OaCQ
1KANlGxbssYmo3wbY2q98zSr3+DVKjv+Y7nzt6504Ezi0W+rlWZGdLdBsWts1Tbh
XGNSOQbOuTKMoe8rRku8t354TlXaAvZjMn0XaUzkUi3j741DHF/+qAvM+gdsGTIJ
Xi9xpjUpMU6574NlsA54tCxpK8V/KQOQwTRjdQ1vOb/gqpX4bSmOfFPg29o5TivU
UAhz8IudwemUZwijnuRp9RjiF5CNOSdBFuMRLX1LItDktpsbb7PJqW3YIdjn7mwt
32Y03ok8I7/FFMVaFGimx4Rew4v/y1+l1AD8CUs+dZJSOI9zHJooXjjQNoTP6JFw
bMs6y+49nYustVZM4lYNK3AmWgCxgPKqRAu5GPvVK+QpxLWHKnzQeD/ZBe1m+fzu
cJEux1qTIUh7lGr5eZ9d/MV4/lDkvaWtupXcy64NUloQzB6tKUe8rLWKZW4i/Tnb
Oc6RO4xl6gzx4j5hhIVeKJmKJvoChSztSpjZ97lpV8jMQbJjlQ3QDlEw4s5oxVu0
ppaYXdLnJw3/p50jS7WbsQ2+0y3wlFXAL4cbPlhnEzK+FXgeSRyrPlhQx1657/Yx
4LRsZvb0iizFF2RKRpWIdqFf8rqId/X0YgRzco8FnxaZcpQGJJ3YqZnHdJVPrXeD
baovOrK6l8mIwz6PJtWMkw==
`protect END_PROTECTED
