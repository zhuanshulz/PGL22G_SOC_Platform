`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
83WEzg8l/5Oa7ukzAqNBFjLQEYOGpLnPXqCA98KwaEbplnEeSmOaw3dvaRqWHKXR
1O818EToeNChyaywo+Wba+6C/UbSQG8/sU2jgIpW26UywFMmu6T6LVV8OtiCM1DZ
fjvbMGjfYVidwoqemMKv2+rH5FwzR8RnA01JIVBeXUMJbbu+j/uUnm2F59BaobCk
kx6xBaTyRITs/5EzRSS2M1+dmkrpAomJZzZjvWHAgRDfH4KndNQVFRFrywJp0KBz
hTAkPZQ92asHqSKJt+d42ycUlesk/6Mj0BHW5ys3F0YYBGHlto2kzQuyKugVE67Y
4sSDT+Rdahj/YKKBZcJHfpaDhdDRCT9jZFl9M4Aqg84HKyZ5Ve8wb9G0+dcJSYRb
tcjhAxnm4vjpXUTpTcxI0BAOi2ShBMDbPu24zQiZt/ZSdkJhE57RnS8V0a6WNbnQ
`protect END_PROTECTED
