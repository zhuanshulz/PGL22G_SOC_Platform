`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7dxVkROnYP7Q9opclH4yxYLqoStsqF9JNCzSWs1+gXFFJqHnhRLn5W/1s36rnXW1
TOrYcvdcE54w1CsABqnALue5TFHxGw3FUQ2w71q1nm0MJbATKTfk32IjCyFVtj6U
63N2ak2h02bVzgZOoBf0Mztta8RCuqaJ51PJXhnXZm9+ITW9wuw3TS0Im2BV5Eyu
Ic9utpL/NkEUL6RzC4ZhSsTgl7cudykrgQjhm6xhHbYHjL2ycr6A5rzOfQMd4msp
Hv/k5Yey9VXFUwOowT/c8CsZX0tKUGbN/N55tIc5BjGxjcUeK0W6LpZb1Uk8Bgxx
8KE8Fncr9oiiMD6AVxD1KmAkg7rviuDoYLbPtcfoL1hTIgPDKeJQ5ErX8nHZGoNk
ThsU8impnPDN++zetDqhiZbOEy1euJ5ybE+rbWn56/wZkOuyRz+5Hm1BdlSOjr2u
JZpUHg7T1jbQKKOyl2Xhj/dhf1yo6tMo57wUINQflZIRkQYDCgW3Ui1EuUwoUPLQ
M6gTPzC7lOCGw6bF22HZZtz6GZUT8FhqYdYf5/XP+HeayDCB9d/5g6s7DjkSxbrH
i0ZHVJn2dSp/kvsCR4hiurM8ECHOCk7CpFrNHn4ZlrOsMnh6gAN98H1q+MUpW7Hf
0uNMbDrOaaqK6lHAatPTMiDLsC4l6v2BUC2QyWLq+AejGwNtYgJv54GCYzMOPql4
2igsZENfbvrLdVz/5dmk13nsOZ/QrDG5EJkqfA0HDKk2/eKwmWZPZg0wdsMMdvrE
1cwtQ9nnTvGDV6uxELwn0nGkzVMjIHfj0cXJZBZGMHaKZe/ioc/EGqNDT3+84rHm
HYV362qb7zAFWTi8kk4z4X9VnSGDXLwIDROlDLLLwS8kxOyQ3H7AjntpUVqV/V72
bSm4UZz0aqPcDsxuO7dc1/ikx6O1pyHb9hzty/u2XiHeBSY4v9wD/PknaXMYkVvZ
h0WKaAabWZyYfzDtQTEE1dwpXJwdX5E6EWffybhnNVIRrgHZMSPIdO/hO8vy+kFU
wr1OlZQiganbQd6g0xGeVcKQqXfQ8Bso0zdZze4Y66/a4Sio3pElNotdsApUS1Vs
`protect END_PROTECTED
