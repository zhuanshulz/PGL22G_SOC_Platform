`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TlMekCrpW9uJNjrc2DzTVyWXHoVrqqVsB651BYdWRUh/I7trs2bxXH0MAAWJlLht
h4MvHQrBZR9eZsLeegGFEDM623lgFThBBvbCjSm5K27atUbPSW0zCmOBpmx5Y+Ns
zQqX5mVCfQ3GeW2boPYS+0F3135rXZoSpcTx23wteUzsTh2tGj6YjwcQzKphclxo
OyRTmGywzPuzD92dtjPLrN29qkwVDwsBGcAOAolTpafO85bCqeFnIO77TmZTbNLy
xs0dpaWYvcBXYZeBWgIut8Ip3SSkfz35PE0srndtteANfhLnN9YNKEoHGXEtDAZZ
g38uouSBt/6jODdWc3N3DyhQ1j70qqqZXwl/8q4EfhDJJlbrRee3t0xQtR12sRrM
gXXR/CInwCVzOA30ZS22/oC62/AG3DkLr9IfptWx81CkFaVml67Q2q2svq5VqWiw
x2aXBWBsIoH7dpcci3liBCO6hfJcSNJFrtGtoaiy6tz8wqMZy5J3sJ+DFVUNbm2o
dqpBOFsiNjrDYfHKAxvDDKjU0BW8Ki/M9vIvxjPe32kigR5QbUHVcTujqhFWPNG2
pk2m9VeI2ugNL18pEoS5WClYxKzlxfhZvM8mCS+OsSjrE0B0k20Z9q1O6cOyv0my
4L8iJP0xufKm0YUWMJniJzLpTaK1hYHMS6EVbCbxX7bGLbLoMVhbVOvwWUKf5XF5
PKU/zFt6+RphBFZRwbslkw89yIsM1rojFP6304YoXGSDJQk3tinM+dd3lEb26Nyx
Y7ybxUidYZ9xyev9fdJKnECEFg6A0f6wWN2Qp6YcGzqbx14HDysWNotpOIDaOIh3
`protect END_PROTECTED
