`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xdczztv1fAGNiyAtR895yDG/6NXVvGAKzgJ8A8Vp/DnUQyx8EC/GVn3oS2uUY4Qa
QacPq4RIbtaN5pN3wLLGVd3SDZWHfuY5HNMyiPZxOcqOUcb2RpMTOupXXdoSDfwg
RjbwAavo9oZ+KncsPKYQT8dY0B1DfVT5JcelKsrOSvlsQd86uD9RIirc5asDgbHu
6cGPBNJOwCSVsTIMk6M7uy0r0/BkFdAY/A2CzXyghtTuMoO7uG3Pvyl3f/KVZt+m
84ndOZ/bYCWAQyhz6W7dXoznxPUXslCvj+x5JIgiati3MMX3Bl/7o/JVTJbbygxg
CDc1AdWHmqFee6E+5fprDGJgnXM5gLX1pNmpXXJ8YjuNAXZPCIP/W33a+zujZV6f
we/RdKNZKNvUcDKt0CUsvxiFlfJBxzbxXEZppsfF+KkqQiDCQYvekZFIBB2DhZm2
S1FbjQANCMGyyc1HtoElHivmDzN3LZKdk2bBRoe+Yb2OwnfjLoGDEO6ZPWPadOv1
nlqkcpIXrYwsyq0NMpk0iNTm0o+1rSVYT7kN9cz5WMQ=
`protect END_PROTECTED
