`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wCHGkB9u/oP7ur/U2qg4zVtvU7ocTwzx3Y2RgJbexSwGTUxkqj2+mParUsBhZLSm
LphP3L8IRc0p0vq+d6DBjPUf1Wgl9c7FisjPadhC51dxOatdeDOuEJEso/gb4d4P
ab8JrFCGCl+u3U7JMK71E6C9iVs/bVZL21agsg0/59RkfwsPE3M5/MFjV9k5m07T
a+HeVUth1wKqYS9FjuhPvDnmGTgxaY4r6A1gvWCouAjvwOy2YyLhrhXjT2BpkzbZ
i8ai3K7jQlWgrz78QK81m3ZoheLwtArK/03sQkD2jNmJMkjq8smGBFPrS3cASi3v
9SgAgtVjkJdtMEyN4EnZeu8bGPWIVu2pM7jmgZ7vLS/QH0oe7LQjK5WYHNJ1Pt7A
BNZIF5ikqgv4MNYxVD1uNad6RewcxsTBTuWcCO5m+bYyC7ouQa3REipfUxbuVDU0
`protect END_PROTECTED
