`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qYhvBFjE3Z9qMLvCLyWi8vkFu72dzCpvRKrzGInr0j9XZwPJjNONjXpyYbPPYMA9
O7RFfjLfwizl2C1n6v0FQ16CQKeCvl46U3KA6w4zZzXY2YvS2GTLmF8cju1/q1/B
rR0W9Pfg2s93He0c8Xu6Xr6KJUxsbqpM2ksTaC4cfVmY9VhSJJctrMyd6Fm2HWol
8q3HGE8tOwNxQQZ9vP5mSrzb03jSg7yyamta5HExnLV5amuAM39iIXpoC/G9RURb
bFfpkSkjVWbHvY3DBQKV/YzipFxTu9N0EYsJCiQTrrBjqXFUph1rhGBzuwj946rq
DhpfjtDIUDvoqSwht0in7LrxWdJZ4E4Ilyw5Dx2ru86O8FJh+T9q3inS6qLyrTkU
1suGyvenP4+Nk8d3oqLBLB//dSRzcV2S1pvUMoXiim0aOu9075pDXQFMbPbKFvxU
LezoQsYM5Mns/uncYHDoxOXhbbR7cDiMVmpaVHu1RL6xj4hulFlqE0a71+zYcCxk
AOV+ItrPpV4YurmnKhHCyNHm2nENP2TySZKB0d3bqQKC3Gnzu6toMv94BgZ+XfNq
4OzGcZM/1rv5rON0Q5OyGnCI8TMUwzgLelmDpP8K3RqyOqo7eY5mrMmHgTYcIP9f
sVywKHASP1W7Cc0Az0WYLb80WBsCtX95Mj1WKO7rxHCdUtEOsYAmWjOcnq3/J8hD
7o9JUWoT2DqWB3IuMm5AtAxVjK3jT5BYVOqh3ztxga7+a+TOS7zwOrWO5hsSWPV7
6x0mQo8PtKCeFupWKAUrt9G/IFl6Cw2qdLXZ46vVVAWezJcC7kvG5d/qlGL9E5mw
rUtafFWsknZteJotC5tqiaXw8Qfo4N+hK7NGKvMow2V1z4XyfUdBLBm00q1exT9Y
cnaHlxkUttha8U0AW8rIbvT8bH2WUVWqzKsKPBNLTS0uAYK8WVbxhIaHQ3kWmVeV
Fujoq6KSWIA7I5bX2gEk+8VY2gAWtDeYAlQJXY+OIBWg14Rf8NTzSrrVlALtI/Zb
M8ytoxvbZntnMM0U8nVSxVeHVLkiJfunjax9T1hTpNN+fwOT1kf+xffx4SsfcVo/
EFPV5bXSa2CBct8XoHJ83EX+xoESnE99Luf+JpX+8/6igchmAESRd1izLxxK4Q6y
4Q7k1mUOwBZ0sodiwOYJeHMXiW6g9WNahFWh753SVeYteL8XkzTvTilQtW+oEgiH
n9p1NAZeANIcqZ9aeIjHWW1g4o/LAu9sJD45guIOthO2y8zTIQrjVVnma1h8+XHN
zrEzqpAyaV0t4aNDSmHOuPZZDyIJvFkOAce/kyOU2f03pOwyq8aEUk84vWCSq/yi
uub48uOodf5+P+KLOejlkT52soP+Foj+IRMgNfzQHmDRuM+DPmyNRYtnVwRy8ewv
fE8wb+dULX/C/oHwy6rAM+8wE9htXH/pVma1/r+miJXjt/To3nU28p/UWAi/p8C2
P3C/yDh+gW98dxZKJ3okfvYxHAxvYGcq+zUoveJJejiShJ0BN+L+1X5mz+/SeobM
`protect END_PROTECTED
