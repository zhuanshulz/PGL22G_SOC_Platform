`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ONUDA7hmAqSLaRBWDg1P5c5szDgsijV2mYeZYb8JzBOqUf+8L3FmgCHsiKQdA3En
epcpbJBErmnz3wXhEJXB+GNje5E4cYzQ/EKLpMIsdydwwY6cVaCRXEk+bCcSni0w
8hyhM8+ymRR23IIc2RRA7ZsbyVVWlC++gppcxxxYtg0HL5pIITOMFsEEyUmbZBhK
S8OnbMwE1cVY+s1pvTRwGChIXadWTF4Ismx+pYa3wk9Z090rb77ipFz1siW8PW3G
+KJnbfTn4KAtE2XCdHhTVdte0XfeF0EE7USdTZ3+IkdhNkQ1BRd8u8qsy90HtGHw
54YiynwIOVJ9bJduL9qH8j24JSMMxcLe3fEuIUxq9hY=
`protect END_PROTECTED
