`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zzKBpMfK0Z1v1DemKgYEIyX9uE6tWFJcF4D2aBwtxN7N6EwKhz/jGSOyZp+Hig2B
DJHHzMQCjwBPca4K7alRLwoOAYbvGhsjIa4wyNUrx+kakjVpUVEViuazTaHmDOqc
cEAJVRUAnEHXJc3WnH2NeD2LmGNrJ5bK82AdyjUtAYSaAIiDHouSAEFE2+cCp5uc
9z1JM4XoBIAR+bQNVn4k32Vsy48vIcTiV6P1z+F8OvAlUzJgeYATeOorI3qO2Fq2
3Gobjw9tXRDpIVfe3nkdaA==
`protect END_PROTECTED
