`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z9G9ldSv0weTtEULifntCnpCbv6VDlRhon9jMM4n+nFOr402Mtdu8HCo2WYJuI+8
StFMgAq8w9RQB9h1pYyFIN8rROWcBxxYOQEpCO6r2tN4Kkx3rQ2G7NXRsGqFqhik
t4udQ8KCW7XfOxixNlq4G7St2Degav8L05IynLFNiqJLscgLcsfWlYiWBpmsQvg/
HKsnm4VFlJG3TvOOS5YzXABQglA9bihD0WF/kahxRbsqCOyAin0xxnhKukfXogy1
fAsQ01z+UhHuw6ubmRrMH3e+Hx0EcS/LA4QIWnC4qqBd1WjqEGQt33bC/rIFP1/4
DJ7Oq4/1GY+fg/UqqzlZwkk4SAsohxqm4nzExe/cr1tDyAigPsKSEQR6aMnKaDaN
JWKQ2WkZyNqycWb78M9YPqgzh7B+pmOXRi7qFuYPzDmG9GP6vUSCRoX3zx1yG7PR
+pb8GDulH7t69tMBNhMk0sRXvHh83vpe5+kZcLVvNDikIu33hLg/tPt2k6LQGh6w
/YfSglWhtmSKbmS81ismrB3NCi1SuIWPYD5AoNHFPNbAe/6ohDMY1DYxdi8S4Oyq
uioSjsu7UO7f5hYqrCd8s87Myo7kitLq3PNj2io5RLmk6yju93rS4Ipx1pxopKPo
QIuzbFkmGePf1ElGnfsTIG4jNOSOA/PA4y/BaRy/ggB4IaITCPhwt/L1OmLQ2fgL
7WTm4WSXTHoDGX63al29mx6VKbA5fDCn9bx0Uq5b5j7fDJScZ2HmF8bHSb8iIYDh
O+dQ5fiHTy6um2yq/6H+q7e+YH48gF25b7aur+CjpSw176GahJRyR1aPxxLnMFpb
bMXuKZed4qutQiYbnstbN7wW+4jax/PtQtCaI9Hz7575wHkE4gMp9wMAxKgMr5Mp
a+97vBmEHJhz4H46eitcakkHcWYEe5jEvH/298MpOKqX4kB+DIoFBmugJ6uq6lvq
8sxl9HnVbr3DrCMDhoNKRz/l17FVDTKslZiyn4C+HYGG4ZXFoxQI3Jt/G4PtAK0W
Z241qkmV9cWOF0rm8Zb26PMo7+jcW1mpCfdkwP/lVlUOLJmzotbyl7GWfb02nWtc
ayumvDbDu6wdllh8uDFr8joaFCjHMIJk3u37i6G56pjK1agrLrTKujAYlFS0LN4X
RbiC/B7psHkpfc2d6sz3IGYUaqV/8uD/GfEGzwXoNiVm9/9wg+QNosERFYXl4/PW
IMsjV6cMoJc3VvPkf7biMuSG0hovGKLz0cq4vyf+b6/wCH0+iP5Gk5D7Hkxy97Q7
pgNTnojkfw2L+HOO67Ss4ZMhprwDTVlhrJtBrL0gAKJqi4H9Ejoue1OZhdWu1PA8
T9H6g0rDItLS09EkWEPD1ugWft3W0inuxxNeYfsnBXqwmrnzwP+O4KQfbgF9t8fM
/VE16lglWwXoKP0lmB14zpUrUkoO4oacSeHUSn02mxFCEEtZwhExq/hAuVgzUPO2
UKS37KHWyOqlEM7GJWFNNU1oG5IVJ2uJO7N/qqLKcl1636/3kSmbeOgvuvklmfyV
18rtc9WIDo46J//x2TGYeXwt30U7FYTmAsyFnVkUk25F2g+Paj5iKqd7Y2pZGeSk
qF4hm5O5Elc4dzf9C4yRR6PEvaepEvGSG06sC7fr069IZKcPEh5SYCBRrjU9kpys
FW7/jGFdM3wfUa0VyBDNKw==
`protect END_PROTECTED
