`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A8mZo9FE98c0HGK/c3CyPQoG+/yg25imc0fLKEuD0x/ap5bjpao9D/rV/tDYo9hq
1aFo/p6qCPiASSXqTqkYhvhdZixGmIuoDilS+p7HI9K4rSzdn0kD0ZUqSqs81Eq3
r/ca2UkKZVp0IU/WUBNe8hhxMi6O2cclVNC8n7n84RsiktGJt5pXceVUKSwVZ+j0
cSdlrbEKwLC4/pQ6fl/dU/wJD5hV4Gp8F7YVoV+57Cz6WvGIYVp25RH5QjZfRl/M
RnLsmGbqJYHi5w3yEOFPkydqkEGFmqUfHU+aYT2sntXeAcrgKgSZnfcX/oTtx3ce
bEFs49WZlUIo3V8e18HgTRu3lPA9WoimdEANX/cW00r5VN4wkSCRvfl0vp0de8Rz
0p/BeBS7I97IYUcphK+QN1dN8sveAgL/SiVqMip1dBbvoNz1jax890XXzJH8RwqT
XCCQz0XiP1wf9cCuvrLRftfIuGKc+3HBjiqFBkft3PYZjClFW5GGcengTM1ESrd6
ikWOHQQnC25y4QeoeZ/kA08MZOkrfCIIuEvSBe/WseFBTCR2OsxH3o2yIoVQ/d4x
As6EafaG1P89uZassccNPFVdjla5HaK4UYOc4F4CkNrTfJ2FHiCYJLU/0LO24J7v
pE7VNAP8bcOnvFDEEv0NaDEEwzgIThLWW1EZ9WaWHBcZh78Af6wPunWhxMUksXy9
an/8kfxohMZYe6Zn/P190HvQ0n0znuuRFxqaGCtP596+rYKYdPracIHuFe+th56T
RT2dz+N4LE2RgUVSClhM+T70UEXVe2y4Ho3JiBAg+zS5I6Vy1ro0rA19u6hrXVyq
Q3BKatY3aEFTGMzeF5UEiaYNp5YSALoQ/9Fvfhwisi99HsXaVKn0WPng+iA1YRjJ
sOyQCNKprbtjxK6GGF31HRntKD3yQvJISVtkjiZRZpT+ItJe2tcEPO9L0AGosqMu
QSVSZ6f8MRrUACfdmel/9no/RfqjHEipxmOaMV9oe1ltsgWT2l+po0MyGx4N3We3
LBJc8H9Oe1YLJXNPvFh3EuHTRkIE+R8fzMasLwR1Jnm/N4rpe97xPE/QtcxC8tuF
zBAm8Bp+yKXsmwEM+HmjkgCNUxUAcg2Ii76rN9IKR9b/MPiCFla0JLIQltgctGDG
eSWjCpmLC4ZVAdwccpdW+djRZy8Sh/5eKEeYwGsZAqrLock5bieSU5blWyN2s8AE
PdInPyNa4yrZl+zV/COMxQOhwEH0/AqMhn9+DcEqkPMzn+HezLOMKm/expMqHB2+
tUY+rwVfyVP6I4uARwgGbkmuSERqv/6ZrdjnyoIW6vQPIRnMbH2mzGSUaOHZj9x0
LEa/5zZMesrfuX9okOJRbOtRkWPbx1khx4zI3Z8IZoAm+NiVCAnYBxc1VOlpMOk7
NDAIkhaeKi5rLmweaeWvqXEVsyn7X6xMTfYJn52bA4pNviEy3ZMf89SqVmjcbtch
YO68CMafe4w7nDoIAKbq62K0enbcHX+T6DG1S64Z8GDS1evNqMvM+uyNrdA0Jxld
z9wKzGPkvjmw3bN8cIBGW6kjsg6i814hDyhDJ+yYaXindsY9K7x5bTStM0I2PyB4
Y5RbKYg3HITXdiW00yEN9Hyp2p2riBM5Qo/wzcXnYmWNHgQ8Y9rJiaJ7HqjxgUCu
7vgZxAW+WUbpIjz2LxC1JNyKnuRLd+EPkVOv2wZh2zARRoT/ZpLABSl6VhQx9ou/
UNxETOxIe9mglqeh0TBZalIqz5uV0P83GIiDg0pYyEp3D1O0zPwtDvfA+N5vG1uh
uReAGkUbxoatkFap18uHJwLAMixXctaXCE11FMWm5AublSv47PHJVA/3aL8YqG5E
2t39yEvvSAG1HkidUIknuWKrFha5hM0j5FJJbBQORzlpfLUim5ad1SaU0iPoxvPN
1i9f8Qh63quY4d3pf0NYyH9/T9hZONby//ZLNcrR8WJD+6trxtfWRk82eGUqDcOK
JYQ4EIrtd2qArWH/H87yEpqWO9YKpPbRMlQZeYRg/ml5txkUhekTx+abFJLvM2YU
/m+94C9grCT+i4oANE2PpRShkxwqtE4Bv0UMcU7MtJso3bfvoPTRHymhjjNPlg8T
aniaiOc6lzIDbDxI8Mse1m/+scgtRhPy0es9o95qL3yiYJ4d+cXo5NKT/B+Kqzaw
8DYJlMyC0la+p1tWiTFy+qOiKwvnUrkMusomQJcu0quYzMVF+rmD57CMmAEj157i
Nt6VZpNyCZXPHb15f6m5i8f5FFu4YWU7lNfS5zxC88xM+uR2es3iMkNGhxvD6uM0
wftBfN7myHgUOnvqDhWn9SjS5ZeUKSXzdOtv6B6Hr1wOlrzXw5YSI2uncLVZNP3E
D5+FtgI4xRMVOYvPpzF6orn3iebBkG5f5qRrO+EIq9c4UTGR0U76IHW90N2jG3KS
fXF544NVzEonezezAaAPOS8VFeNJeOHfrdgR0SExn/tgmcRyFVOL45sqLeX/j/S+
W9Xqld0vhDBBi1ArjCC6dBtAGlwk3BmfKt348qLofvIV3MHPuQimDtaSbglGC5Hd
ZijabdklSf6lsOnvPfzV6WQEUIh52h3GUcpe9rqBvn70+bDgeDdBF2JrGRgGTyMd
lAOctUoXjd6pqwrGL5ZvxdRswrRyT0+oltgwF7+I8w0YWCYV41iC/E1aYtzqI8wN
kiG2kw0rArcYWP8q6G/oFg8Hfp2w9VM5jkTYxyeiALAZ/wSMr9nOTpxCFDz2U1zP
8jxpDaV19iZsz9m+trKqYWdB3o7TZi0N/kMxMTdV71gPXz99sBRVrBDG3rOTPaEl
ooFIQ3Ozcr9REdZEjzt2JcSDR0sdK+AFhnH9xnQ2nKUeGQTqTY/LhOSr3R5+guGy
ChtVsbYk/Npe9K97FHvQnmyZ3qNt9JhmH9S1RFqkTAmGbPJ/yYzOq5VuXVUa75rt
Fv1AAneua0N0IcqmeRqT6Ov0mkA4oFPRlvjFVFRKaxOnsh94IHK4VzBMto65GiuL
mIghvp+0on998K2x5eoaS9NQfxOErj+bwTaPVy2GVqD5fb/vzdjFVrNgn42GEsIM
zmgydXTl0v1dvCaRE0lIf/ObLUxZ0O3JCK8MxIHZR5Hvnf+nQQ3SkZdMqJNYDSVQ
MonWyQR7sU08CvMIJ5JQI3GcRLTbn+I6ZPgU1VLcmiaKj0rIQRNBSL2wwIyg17pQ
C3apTSGNwGVSsysFMW1F7t6oVxPwxuQ+06+wjV19FC2xaJjw6/KVvI/2XcLYx5mj
g9OlYaKYMl5KNs70Nn3Ns82b8Rae4apRtmxL8nbHoygJiCOjav1JXiwdw6crsXC/
FvOsGUYZU3683VixwOIPCv9+UOiP4OdOmqxUN0M0p8eRulzA++T5U9E1KVGRT4/U
rwSq6mpu1PaIbJtt9FMteDOHgyHvVW4oR1rXxjM98UZL4F9cJatqOt3A6d+OJHxu
+UPBFdalx1prr+vjhwWueeiXx8ljJPaSxg+LrOgH/Uqb/OwRA/p9SJIUNKhR9F7X
GJnYwXkEyk2VDlgPjO+qCtI+xe9eAeQNOt1UpKJCg6JEY4dj53V43BZHi2v0ca3k
sJOmIjsq/qoWdCFD4nxvyI+FfV+ZzSR8+78OerlxdjRsr/qQZIQmWCFSOtLA8sKJ
wC4NORz6mhrieqvagSNVq/3bWJOF3lHNM7IWgj5AbXlUW2hcGHhxt1ujoC5zkm7y
Pc+vJ5bsx8+DvZJoU+oBfdDknwVuDDudQw5ZrxKMMWQR6DI9O9H6zowYlxz4eS++
SBpH7v/3FMP7W+ETHl4/qZEdohqKkce7geq4UmCGXV9KpFbkYQ7BpQcLDufX5wHW
Ks7RZw6G0eNy1iMqslSpcKNfSYNbNBVOAr9bq8rNUDQcs/L/1M75XJaGZK9f7YUK
XkOxOnH8PaERQ+MoHKXu8LzBfPgQGqlDGVznVIak7TQId1UQFa/Xxu/+UIHnG/Pf
OdH13gAr8DEdmrrIJ7hIJhc3tF0rXJIr/2jPWdvbZV7mgVeK8Nrb2btaL0xeoGbH
vmaH1ggKbptS2Mv+dn72uO579B/9a1FSfBtJKhD1Uh26kJ492t+4MD+qTmzMdD+F
a5FzauYI0h7ycwyeWytDpL9NjOr1aMAgYDeXGjTq8NSuYsWldu5AZS+nksVIFHi9
PchnfdpLnLA5/YcjuP8eR5R2Gsr6M9fHdUgyGbYzhStSGQhHHXLKZdGXtKeWu+up
m3AkM/axJjjQWQYMzmeRCtEb/YTuoeN9x2FXIYj1GSkt0roleR2tGlh+GKLztsjk
9ckM2Xvrl+Q/ebn98erzWDITA0W8N0cK0tIIRI0re6N9/LMoBJ/KAPCeyl0dF/Tx
kX5KNQRVFeioLYRSYHSpdAHcMRZXpeamkvV8AGLhfCndWN6QXjt2xqRoQNqIT6GB
PBSI8P45GtJ6q3vKRcrJjg==
`protect END_PROTECTED
