`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MAztmpL7lGPYq8qbsqUj+szXuVigi6Y7y4p5aqv6vONjHiBJtL1rq5h4rHguktku
jTESt8iRt9V63WjY7i2Ga7rUgw6J79/7zVU0HD2T/tYMwjPDYs+QydtkXtW/tjd0
DaAGsdNVtAJiHDIP5aGKyCK/aGk/w4gOb37wYH6lb0MH6m5F6H6bLknYzcBqN+Vl
UJNo4dIElpY2ooJsTJ3BV9MX9S1Y+sdxcbK+AafsjSrXnHwewd3gf0lrAmmH0mJM
2mWD3cv1W6KAOQvwqye4OImibBM2I7P5T3h0erNw6ChjYXD4GwYOnPdTDyOCckP8
hdmOPvpc66QyaytYIpEp7vHeCNfF+XsLclCpT9wn8lYyeY0DW/E7iSFgM/g19Mj4
bZIIz4B+tfNmXuVnKEgc3869XolPv2rMtfh3GYYarub3S/Q9Dgnvw/duX+P9h6tV
bSUCffWvXUzZ/PN6f29qdAfRilco9/DZXWCaHLoXrrpZ8z58eVo/w7S8jHRK3cjP
`protect END_PROTECTED
