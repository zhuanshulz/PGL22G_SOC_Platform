`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
unaHX4rH4yh7Rx7TzvFvkBsX3AzpG7F1wC9S9PcOzrdzMRR8BzRwftzdwztCLrOv
q/HdTP2oySaCpkahRu22WS2ZttiCkrWM/wuOwsQcDVSqYXVYKf6QngCjEWPZ4xrR
/C7R2zQu7yuYuWzpqfdXgb6Dh0QvNn1N/0Hd0hvfZWDswu8jFUno9JEND8c+tb2e
vrq1Z57QWO8KkZUkspga2RgVUT3uyIcjqKT31/qcDS4Mgh7TBfCyPH5d8JomQDgE
KyWfUtMWN+gsmI3vm9rM6Cvk0++iX4NFCM+8uh1+v2E3f9jrASeYf2tjNMG0o3J0
gqI2WOKFzNLQ09wqrjeI6BVpYWjxSWRmQBuZ8MoHmfj/ie3bgl9tkhGh2e+0AmZg
0h8Pf7eWsN+Ve+q3BPdahM6xjm1AsiXR279Ha4JkkjFYc0BS0qs/i5nMPWwxAKXb
zNI+5Ka63Zr2hRQgrNcIppA+9dlpLq7NpAEiA3MpeMj3TR5SKWSJefPc52RXfTTb
+0iNN6zVefo4scn0kZ0w5WDmJ+4E0J9kISp5ntu6xLSXFAn49X2fBCvaLqxOXar+
NDytVx2hXmY7BqljpfUa67NZw9KMaAOz+SGnwShcSgb+In01rLo75DP/znW0HxiP
V9+fcG/VnOEgOgkPv/aC4+3FuYXrsA4b8hKmc+68l2hn6ri8Y9CoWCNt7zEmpFiu
nqR1R54Nj6LLqjp/qS5gLpGj3If2ge/aajgQLaCUCCFTuI0vkrNNpsVybprZ00l0
pkUgUEKaP4Bek7YLPpA0bWg0SHaNhSJHSeLHsQNajf9A9cEJoW/VylY+KlsYKfQC
tHs7SLO10UTS5yl9jEIq8T/ZSX7bUaPVL47Tjzbv3gsjaJ9BRWlzAgZzFDGrKapi
lp1wiV1ReszEypjmdXVobR8suGflLlQAW/h7h+KVWAuFo/MaArM+xYjyD4BZhhBI
szUkxnwLVV1exCggdDqjutNzGG8NcbEhCSrdDZYZiMqPtgdOSEgwyhzzuacF8r3m
6Zm/uJ2U7nmO2VC3T/HcWBiJteZdnL6MhGTaSHCgOy1PCc03E8huyyRkUDyyor2C
EEH4rvw/+yPqQnbSzxtvWDZS8X0pTqOtyPMRVM7UpDIsI4sbNyABEv9ffd/wL2MF
Ov04j36tQEWjlTZ3W40DT/PuPFNq+P6c8CxIeabgzGmhm9FeGLpqSPSkoYwjBKJl
QFFvKeRbjrkEClDuijGPyIe21BoQGvyngrIIt8AdGK8VxiZuBW9PF5a+7U5mFYG1
ptpYfuQu3PtcUqeai0LC1lVHz0YSw43EKaoAWGEy4eunbk4LWrHw0CtN6X10QfYy
GyOQMIXP/1QF7ZpyuaN5pU5QuXKivi0FHMOWNs793QwUH8Tc/VJ9IIj1H3k7pIOe
ICcNQmS5R+A2TdIWCOxUIL0j+gomjDilG9UMrwt3Cf29xkSPmfhCXILIvlGAu0SM
0bJP0QXSZ+u1eN/5iDoG3jqy3zvNDywAV5KOUn5KhOIkhaHbgL5X6+8doRpW+oQr
r5eJPQnct0RsdyagdbEu02tZOF70/3dPY50YuQxBZZRlyRxkWPpA/iY4XpV6rkv+
k2g0zoTuJYqL7LFGFZB+gM90ye8FGDg8i8FX93/eNMYJW9zIXNF3oCbWPm3gVfW6
1FRSCqtbbnj3Jt0f4HjxJ3kIm9a6Pb0Pzz84pesuDxYAnfe7zhsL95VooSUkgMsp
KkYrLQaAh7XRwQ33Pvq+wi6Vs9pUqGPi2MAlU4si9ABl+3gN+VChkBOqDSJkLx0j
20MoJqdXiCT5I7j/J5P7ONXaCOO0kgqMHvKMGT7adzU=
`protect END_PROTECTED
