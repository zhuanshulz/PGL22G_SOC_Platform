`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cJJwLSouCVwPcmryZnM5IsKBWo59/mP0YsGVCe1aynMF1l4QYY1JDr3GiPTI0TRs
Xils0CtEQpO4CNMkIySFfuw0xVavMuNuXfuNl3zBkHSEQe7OTpFHPBEZpl5hi62H
joSCI4noHx4lEPna5vVZxYnZp0wOUgOvNmMape1Q1X89PT5BZG4XgJPuup6/bnaM
d8dzj+7uCZsEeRVQ8g4f6ur/tF0OMZg+gAM7eCD76YR8YgiX98GiUR9vxmPTlq3/
HVikIYmVhWA9yPfFuR93ZgHBlerY5S5hN7tJ9g72mcd35Zpc1np9lmGPmIL0cxLi
CSsbae/QxvKqxR37Z4Fj6bVTlDI7VHFcD3lbUYpyqblxczECuMYTMXhRTcWFP33a
08jrq8uFFtwWIsWdAtHTOYlHzmixx1JUTk9AmOvzt5w=
`protect END_PROTECTED
