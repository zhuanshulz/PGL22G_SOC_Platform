`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GW3/HfFqOZ6Tls1minm8qQterWmnTmmpJ+5uhd7hHkQLOWokcMwaOuxDWv7XvxCK
EYdPQjlSlZ1hfqfyHOXcPeGu58SJdqczbeNnu3qgwkEdkOv+oHEcsYg++iKXAzb3
7sa1jFfVKCTA7dx0ag4LNU0E3SumieY7jLu5J+OzNgdfOCFR09iuj8ZQSrqPv2Mq
Qk3uoKX4qEWVz6m5JOXW04xxbwLccKc+d/BYAcYZq8Ebvm6k+EI2NEZ3Gu2nj/PK
qg8gDJ75Gp3k1VdjyIiQQfIFcpufG2EWjIM4IloSH9CnvjIvTgQzTRY9QcfckKCy
+5W+x2kikfBMQs+FiBRQUW/r1ySE8jSHmBUD8FbN7QQUTYo7dtoLh3F8miZDYQxd
/Y3bQ+cmajXFzxujuA3HTfIIWa01EvlXFb4ny9sa6DAbIXvV15QMgAZv3Wp8AhD7
QKJSpox1onf9Xzg19Os9pYh4MkvBpEqdWaob2j9Ka5y/etSMrNaKlEQiwpNohup2
evfLXEPxmaj4b47O23df+9xsRgzGKjzHSE/FYuBJ8jlCkcpfWUO+cv7dZOyVmpHX
pCZonk5H+nuGK4KNQMI9wOdHTG4bZHzb9SSWfrH2o01hqIsxP+csk7iC1KMYtCFJ
QKnPYhZlRoppFHVnFWZ7TB1P/x0xFZCCcKJVHaYzbfzWMz8VAZHRZkImjqzx6WJw
yeNOlSRkiA1zUKUGoXemgju/EUYUXbLnYimhrcLv6aNqb/+L7TIURGE1rVgIEVAz
SmRApyTXPwSO+2k3pAcZLeC+iSMRO3DtsdJdj8nj8HK5HW03f62tV9FAcyrKkujy
Qt84obLhqpfiL9H2yfoUNY9logi46EebREyhQYT3CZq2U09vJIVFcVJ5s2GEE6Wz
NWiXD1tSWydTOq3Q1XVdKafMtYTJAaxezdKTLUUOsJFBAVyZydiCqZ+OUhXBtVW5
adwrMb2T5YzMo4ZQKHpSNVGDrAiFw/qBTZmqdlpNkARv1W0njU9u8cqmIrJuq/R5
ogpwRExoOJEr4WeUV0yzrpxgHau7a/D31C10D1ujwG+X/vIe2U1T61GWimxxePl9
pN/CrDoWMmsv8NaMlh8x8h/7XP1a1v7YNcD7/acsWxXIp5tii8CMKHrbOb8uYgBq
nJ+MW8mkIDcQ7CO3cpfLnrxa6ULGzvTDdKusxF+9UGW4fduvesj+y+qlGdt+fRBX
OoWok5Vtvphre3NEWX+CdkjAzqxvfDAKilofHW85X0mnc9uhzNsQJpRyF2sZupzN
gpyd3b8HO62pVZSx/fankLW7WIJ6IV9azk3qPTAnj/D6tiFGlYN8i2grbpyTbAS6
l8lw3m8pX1Nkjpph1by408pRjK8XfyRQ8htzprCd66me2tPPGJQVW2M1ZjSn5wHV
2/pZTAHwslIvJTxv7Fq2ToBOR1Et9P3H2YRLndTOphZbaMgStnoaZYj4Z5frQOKJ
Ux6iX81Kbb2S65F109KLSE9/g9K3oU4QL82t2KVEPDdboNxNgiq5rFrqRydOg1Se
lqoa0vbZBOX8whhHFo7wnH7QVNCayFyKfRAIwwD5T5Ol4QS14zrKYmzTpQMr8avI
Gp/iCgmTyPt5fc6tjeQfLT/bN7a0+4Si2sWv53MxV/xpFP9BdtJSLun/fdxqG4Oh
afMCljsTkAr8FstkCsho8kw2k24IN56cJoNTuEWHEZ06bvDH073g6LcrwCwSlNpd
UeN3/tWKY+Uz0h/VAUSIrq6bnxLWJU1tFMgrEyDf5DqteINYaz/BCfFhXunrwwBy
20AwCsatCjYuff/qJinPHyg74gUns9+oCI0n2/yHMLo4BaGQlF12Fb3KUvrHHqV8
lMYJPganZm/uF+4/IZqVGayNQaDNoSzKwKIJ4+UMybBIhnMF7ONvAjRixQbXu+fP
mpreXpEvRDJz+REnLlnEsTf+ke33lx5RqN3llVzSNFqsrJY3/O+kSxv51McW1KLa
2PHLIsxwHDjmbv/d9g/iwMpuHvwqx7Y9wS3Sie3wg9nfoG77XmzRpcvesyl1DInR
IE3sgtLVU+fRc7dljV/+vN5kvCFt1N9Z+pu4owb+/snia0fL8OW/hlBmo7aG1cLY
MIyF/GAlCNtYKskiEK6KaNH31wI5HEKqrszN58KPFyNodpcqnHq0Yxs+NFRW3hvU
hf/r0q5vwLz49Xs2+Amu+ab9ZH9vR7UsdIV/j+pXwMerpXK4aY3JF3QcFZiuL/df
M9RqvU2sbzgclrtcAHAlwWqYOZJgcfG+b9QPgoIkmwpxZORxwUFybawFAJC4SDpm
/tDsqtTN9G0YYrAwPeHjxTnolD5kq0kC5pBAdc2UyhGxyK6RFkyvCVtPAmaUe+HW
dioPD2hUmcNwv1TNLj/Kut/SBH4GUYNp8XcPtbEmmMbiFyEtkjZ5v+c7ybnlCu6B
pxs+PFZ8IGNOu7HclPQoGyXqjH5sA/R8DnjVHrYVXF6th0GJcYr0SmPrktFkrXc8
8iHRArPMivCU+XqUIiBj+jBg+wmN5XnH31o/ku+kbLJxrAQa8j1X59x5x0vG23Wc
aEjQu84mF1wy+dhoph3mYf2o/0rrJnnnlHxQWkP2Nnm4RHdZ+g2oQ6U6kGMg4hAg
XY2bkzUo1H4Kr+3ymephqaw+fMh3REbDmpmGSwy4C/iRxNjVyv2WlPqWMFx+nqAC
tUWaDj+DUApdYu0f/gi1WPwXZOwX3LDaocIHP9yCw8wlNrM+3GskIlviybQsnA02
d8TwLcojSRM9Vms0JI8omuVpVliWjdOh8YAga07hkFfM4+zJQ+GGNE1rS4UBQtCN
41pavBV614DaJgPQlQkSY1DgJ3XcbwqcEptq/Zw+ewZIpfIuSMZhtVgGipQp/c24
WHaASzXYUARDjMjQYoHEb++BYzTKHmWwVG9FS20HHw9KCJdMCz5R6MPsyVR4INh2
++C3YjUHQXph/O4CoSHeEtyMkUI7XLCOhkE5TOEJr1QPPbMnvOuBrIl14xZm5PLf
xU/KsqFq6KlCCTD+WfQwUzOXWdHalSBuAw7CXhZUqcqxYQyLa1Y6JOaRRoShFwCS
6AJBOi9FBbwQqarmR/Tg+rZby8/VJAya5pwi8Nl8FeBuqw2gx6HIW0Rpz/9fjsW3
nXguWMDprikfFvp0SBuzo911CKRbw8nQXRvz/JmEREBmxm6NG+hsMutAK+SA/f2D
QwVV0zeFkyZfHVsnEZnvmC9QJm2q3j4mm7mjDS5eaQQrHDRDALjT5UyoQUc8UKJi
iwgfHU8LXPt9aPKI5YVo+YRLi7bSHHJqfJYL7JKDIuwESS6w159C/778TIvRaMtR
ccWHyg42jgqjGceJ7sD0G6nDrUBKxb6KHzyQzHK1hbbs8tvwmYIj9iM+ncs4hAm4
1A6vfBv0a0gQ9877XWWbHYzYb6qHT0x++c2sxZS9Sl+vYy8t4GyBy49hGXNdF2rE
NhfUGd0mLBmsJFmkh/9htkCD68U1vT6rbR/25VcB7cK0enbYMw8AZaBECJTcHyug
`protect END_PROTECTED
