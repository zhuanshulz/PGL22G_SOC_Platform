`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M+8MlkIOL/5uCCungyZ6kFbawNCs/23lI8KdLrg8FDumTpgD3OBldDxVfMGhFfls
yQK67qQBYiWO9QX1BaFBJii7rvxrfxIqACFWx6EO/fW5VK/JwhsY80DPi0ta6Z4w
G6pxDf6mIswKLvl19hFE4QS15ITlFpfghJK2IbyfprHhMRXvJGGfBo+X5wHH1RnA
Y85bZEq1bbKK7zPfLa3gwxTRLQj1MT1698mj++CbH/zhd3iVck7TpliTAj2yqMuW
FprWfBm8O6DwDpNeVH3n0dqYc8IVfmoJY1rl7PIJp7ea3Xyzu2CePsF+HacuqlG1
gHDVgyVboNnH0HhXXi/BRzxtFTEUIJwDSAF2awxkzr1KRjc/7GmBfFcOeylEqtYt
cP3XJzG+Gs/e1Zihiuc3FItGQktsRxi/ce6G6JfWkpORleVfpvVZbH5KYGZEZms7
ShsSa2DB7tIiS69aa3tpKTBvzlzwYx9fE3A0Dw59cOJIORpBV9+PgqDERb6nCacW
0JmbOJs54/fvt7F4UHiZIEIUBDs977e66mTS6LwfIxr4hyBZxZ6z1XGIqR4TzysQ
hBG+ayKiEFt0XOv2XJkMDcbnDRisEAx7sg5VhYVtxC52L4HYZ8Ev4BDYrGIRrBg6
QpkBanZNBATcjJOp2ap1hdgSmpcjWahUg/n63QqX9A6TuXbuAov8xZWVGqKkVVBd
61xspNiHExXb2wtownJ/PLl9afxYJYkHl64iV6VN6pkSOCMPZeMvuBpGl5g28nlO
K/SqURhcKzvAekd9o145fHsY4SdlsgR5pQsNjzeGqxGdqELQ4vBnfM/wasi9unl0
zN1c/S7BwEZflpulvUE2jmPuwDbJ9Qcq0nrZ2FkiHKoX11gwCFb1aCuOKR4P+NqS
FpZXjsKrH6C+GK9bwoosWVuVYhIEISK+tA626NAnZKxFZpEVF2/1F15P3EiygxGf
a9OOz4C6dQW7Z+X9cND0vIwsCLc7tidJP/LMXK0UUihuG6TraYr2FcqvQbUNnRiv
nAEJsdZZUOZVssgO5brXZiQiGRA1QS+m90b6Py9ULXFoQ5CJKL2mszzroFMgMdEw
Bw/lv8i1TztRzLioIkoBZPMzlOnPtwFyAOVl64oHK7js2mG+dsGbMQW/IhDSQDmg
KN+gqdYHPx7fKCwcgLcPgabfB56sW5X8VP8bRMtsz/xREwEvA0PdK6tiEAWR+Qk3
jtjhG0inKGsoyQobDmM6dVIvRs91ohnW9bQr0XaHgs5VEHz3ty0WwcytPPcEnL7P
3+yb9A9yuaiXDhJCWUxG9ztLDMyZUg6Hxq7HtfSV4z4p1MXiB4CwpFsG9ZnZFhB0
5bS8D9b2mLKKUDqXYJ8OcYPpkOTb7chhpVUX4fpaWfjP0yRpiSMN1zGm2Qd1/LB3
IkzqnLoeoi8bQg8/k5YMJfDBz/qrm2NrBStQJbW0gKtOqxgY4pTdzwFVHbk9ll47
U6X+yeDxW/No4NxZ32rnQ09xq83SUKgJUCggBCGbc+jRRkhpQdh2yhdhyPAWCs+Y
NyG3vk7AT5q5uJSyZ0CeA9OUT8zVJ8hp2bJrxZrsx88d0garB9MiqWMr1zmrXbYJ
ReuMd0cg+5eQynK9dok4I1jKVIJ/kvn3yBx1zZTyWMwe2Kscyomtgw0E5VF2j9Ft
4OcHSe76/ZkdykkrWotG29jmFienX6GOTVom/Hg3UXnuN8/RC0iotg+TOzPxD+WN
LHnRw0PZGg9FGsX2QfsTyNHmu4NjaUdowZJ4cDgXaWKMQNVWZR9iczhbkL5IiTGZ
rYz1uHxOIaqJF2u3a7etEA==
`protect END_PROTECTED
