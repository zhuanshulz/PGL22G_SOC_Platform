`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hp3d+lSW9yA79k9XbDFg+dsR7uJmBQNzNdwhrI/z0KxjWAu6XhpWzBTGGuG1fhqt
pU1LNq0cVgYzvsxG93aepUzHex+PQnS9fb4J7eHNVR1ZStVUsiC7t63ZENxbHZMO
G+u1ub+TCFtHe/z7ifYYlyb83d99RSSefI0wIxxDgRU4gle4mzBR1inCTh+6pJt7
w1cj6mbr5u3Uo5AEZHvMnGR0EQzvIGoPATt8eqgEDojw+E2E4Sw2ivbZ0CiQR845
GZSSqng1XAJob2A/gyQiu0synv7Z/xkuVmuNeuiOz4Jt1QirVNDwvRmaE+C9XQM7
OKYzM4m6G/b7HWNyMreY9OOFHVWw1JRq9yeJX96tY47RG7Jx9xS9g1XKpManHCIj
7Ht0tFq4uMcRojbK77ZKXPyrdPAHiw/z+4dypu8jcf8HwqTTVuNRiF5xMoHKSWX9
kjN4haGo3PHfp+ro/OUx/6u8pW/656fXexPDoxpUcfeCEW0eGdrgt/5fe/FoA2KH
YiZRAyB40dm5mIE+LM6Oa8/bVDw5KH0zw3K2TzwzLkuXvAOBb4ucjIlGfROP7YZN
VBVZ7nFwx16glgPTXhHtAjPdbOVeP+MWSAFGdGgS1o5XsS4as7rvM0TIVGZLwoKW
Cs+o0CG5b9WkKAGaSFpFvZ2Gad1vvyy5f7DsT6uj+NivJwe9yCkj5VsSL6VEYyem
GEmgLCzl/akqvab1DWz0ndwmRDXWi2hvBFS4Ko3mjoJS2jz6LyLlT5nlpbobjvQB
gPvvtSZOvP6uElMWVmPDvIu4DLNXxXOWZ6hcEYKpmwVSh8SsmmFslx26ZJy/uMVg
7nWNVALBg7f9+mp4gZs34WR5KbIJVjGepGFiB/6DUZ/P2mgEAKb2DyG9OCy6JpEg
VuKzAwyODm9xfA+ytKtaLKcMWrwBpK8Lo+1TuwSsG/n1SdZXT0+Nz2ta98uGC1vy
bxOkceBe4SY3/i4baP9alnj3N7/I/y+D2ebVmubF2lZodGWm83qiHbriXIfzE9LJ
Lwl5mnP0THXwMaUiUwekzbXYhSAZNg8dmG6qg2KXUKe3fYdPDKNJkQ647LV94Xt7
a7RnuYlRI00wHrX+KDRqgZmO6XwUW/Cdfw8uuYMAy808ZEFzWal4RsJjK7pMVQaB
uRrhSqd/J5gErawHhVECMA==
`protect END_PROTECTED
