`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XrOlNdQTrGZWY1p7aevYVP1WKoSk7wQf26DezrdSBUS/6i7DiqhoupgDGFQiZqSK
cx+gS9BsM0348VbhbysJ7XsMxNdWcLvYxH7i/r02i70I3TfwtQiKmju30h6dy90C
rAoq7hg9QaYfNwh1GGlThO2ErkKvgGZt/Fv2RbZ6KdqLwVpKgB2bhHy/+LMc3CMY
0HuYfxYC11n6xmmPlKeLuHWMBjqp3uQUJYdRAtQZ+7vBSC4YYLPqFLHrVUb3vhyY
7QZeuOqnd5ND4AbfxJybnmWrYpOdEiXCLoigCmBKEvNKTeQ/akuI4LHGFN/SpXNm
0E8YoBmea3+/TyenNt1aF7TFrHvUnkPsY+P5sFQBeu8Cy9flL7yDJBCxfzq/54Eo
us99PcXiQC48E49qNQRZ3qBo9Xsst/BUWF0Rj01Ux50TP+tTLF37krekcNLDuUf7
Tx1mM3ynNaNafRG7FsEvDzlg5Ls/jNFdv9IEnvyhOdecN+sBtXl2cZ0VXse9Pb+z
tMVj8OcG8pJ4GoCwOJWFUNhdC/Nme1QYU/MMd1UjlqusEWTk/TLQ+Box/tPz40Af
HUVo0aZSLDYupcQJ1GHLe5oiL9OButhgACXeRkYy7AkDPhx4somc3+J+Xyq2dqM7
QMYBy6wfMGLJ5YCAWmlHnj/7DEYrYPl3WZXKuBnxzsR1Q816iqpzUKg4Ft+C3fT0
bhVKgKoRDxjEMYvXxH3z6xH6aGHf9G11Xgs3TqPP3DEdsbGZnUFjVVPf2uJkRh+g
FTIdVDGqpd81+Ks/ZP9rAw==
`protect END_PROTECTED
