`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RZSfAWmuiFh2GE2Nfiu6j75z65pjc3aVLXtPl4NmrPDNtncQW5cqel4hGfleNdeH
oa0GB3Nq1+oOUP1TkZEMPx62mq1Vf7cWJsagbaHyjqHsNHfGOgfn2KqxG1GRBEVz
OwcimUKM5JmvDB5KndN4OyPObJwkw2mNlnZ42+FkUJkMIBnnEDBtjhdNf7zKxiHy
HL17GrCSp2SQl6tZ5JId6JOU7D661ciFq8oEMD3cpHCsuuIw8bvITHW14VQ5tPcP
c+irGC65frLEzmryQht1ujcFBPbWfR9QIMfjXH4dK57m/0qXiX21DQMFb4VCE0OG
TGK7z9QtRy5A9dpTmw+sQz6yzxOESSCdF0YErAYzPPCVE8/EUkfn8viHgt5e8cbc
Lex9RhwFJBWgfZWe8MTrl18qPjiYINBVvmW36bFQmRoIXH7kD5lnkXvggtdySPES
0ZpwR6N+qYY3aIdINLLKecMFWK5amADDNzpPmPgKBVt/ntbQNVyFDFge93BPm9hj
oVy+9dFIZYVP74RH0XkYayCo6AuElqexH73gzICAdzw1h784y426WXPSdMf42S+B
21M136byz1VaqJag0GcWjIUTY3KV8/mk/vbRQjb0nG7Pk6r/V3eVmrsJcuIRrnHv
3JL9/Gs5qTUPadWkggvopqpAzdjbRqkfBxKNO3yjEX1kHgOKL173HiBnbNnpsKAe
`protect END_PROTECTED
