`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A/TssfcBQE/0q762RCYWSbnc13wIztz1qbMn6W3YIdqP8XCr1z910TnevGhW8oJH
VcfmdY3U96D7uHkh8SKA1+lSRcwcyTZYnZ9AjllsBU8svbF6ZTJy2TqfARB8Re+R
5IJacpYKpBV2aRLr44oWkeNHL6c4DRexJFMQW5g5pxveaBreyGwdSIrJjxsam25D
6/F2AhdZ9QpgQCQpjHBnnDgPPX6uRSlGhoA1l0o6aauBF0Ry3HOALhLbFm9x90oA
78DRd0eGVIJtDCkc5zGd2WhL2gketmfWvPJfCmP8AzX+2u3x5w9ifW2BRXadAblB
ixh/aG+xz2Eu3xw4P/a20oP3IE+pU1tIMapJMKNCSM137L4eF+8kGz0msPfwGGXJ
MH4/nBugVYt6BVOr4MYUbcaAqzkxSo9WDTxEDkYLzP4VPFSfpNy+wRrVcaYtb096
hzXlEAublJAquBFggI+ROuC15XnIOKvb3IpWA/An+Nf/IDKfHSvv/aAb62rcOkuJ
2wmUHAgMAVG+sX6qpjK5kQWihFrr2m1Qbz2XVfMQ3WZo+C5Q7X/7gRaAc9Seud9s
F4kbI3hZaRKgklDo16xAlteLW9TV1tN5atyiZ0ULHuollCdflIJQdNPFaV0jv5KJ
`protect END_PROTECTED
