`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gn8cb7fGeJj2jMQ+csqMElm7fbZJOjlcRsDtDcAYPiWXJERe4jipl9mg4wiUPtdd
Z9VntHH1YsgqgN+CuW1/BhBGPFmp+HpyYTCd62jIs3Tvlbjke7mIbZEfbzMQ6hdn
WzB0rOh9mPt8h6i8ExFLymyBaSxjDW4+O8oRWzjsNrzMVPdBvoiCXMGG6lNsX90v
6oGA1f5WKJ+b71+bDc3tGztJbsoQ6Wf/XrasTVu6D5i8jId8/0vr/X7MTPlpxcSv
Jp63XIwKsXHGWkrZRBtcmbieNFjY8BJuJXik4Z0Vpa+k2sMNsRURcp8OlMAOX8/N
rQcQ1q2UmF4TE2Rwytr6aQtCiCbCZKqX1jcGT2LqTx3QrR332rH2nrRl62IrUgPG
`protect END_PROTECTED
