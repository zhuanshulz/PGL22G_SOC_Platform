`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/zBW0RJgffiHedeKoNAVKhvd1oYYJcK4l911VvnA9GATlhZye1g2b9G6RRvnJPZB
YC2EixR8REmq9WyrAG1CLzuCSiTNEpqdh87WRdsWLha1Sb4NFOzPbx0EC9yboEd/
o2qpeUFi6eGIBMrelmEe22CjSBwR3tPgBXZRsatTZqSjxjrQCoBWflalKn1p5STb
2T9e37w/t0Is4KdSung1WZY3fBXslXRnwF5O4wBudPBpHjgKhz5kUtUS8FlNBWmP
YyvhZdfHRFfv49OeZwcE+IK4vSvDrbol3KwXcepWY9uUu01HtNBmMg2x1I0VKYBv
25mnO+KvPRxY1RgCBt8Y7MYxiNWjX9K3ekENEquT3hqWmWRM1t7jDZMeUOIvML6O
EKyjt7We2mAFv3hJ0G57hA==
`protect END_PROTECTED
