`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W7Iz8vP8ok44evBWEdvOK1jFwuXkJfm/9lTe7Gy2+f3wmTmcecYm6kjh07r50Ul8
7JcGX37Y5B/qoeRNa5QwCMbz3sLGWdrtoYiTK1Nh3pQfPwnxiUggFlJTfaNMCha6
kqvER1v1OUlyAXC1hF63bKj0PneafKCbYsX4NuPztX2YhwzBhkTAS6EvOaZX3BUH
b47Xiot88NhJYEhFswybJG3vUy2FrVtK6AviDxxjW3vIrHLG6xcdXWkW1sJJuG2h
SjyaFlaFVamYCS6fFLLEu+VEwf5euDdpRObauHGfxTCOA8IdKmMJ1fsMhON035aX
N/W+MlNKNMVMkoX79wFN6mroWwHFcF7YuDq7KDEMJfNp3NEIPL35XUQ/ZWoHA0t7
EJvwmVZJN4IP5TqV0WPqOeyiGyR2ofxiB2VnMc1l0DC3Uq8SC2y8fXsWhpg6he1A
ZDJJwLfciPX0uydr7bQWgmtUOq2epm2aarCVU/FRHT+mkZp3HahAQILShdQis/QL
c9DrKcsmHm1Ln5IxxXl2zN60ubiXwd+1kkecc+7E5Np3XnrJsAsh+J8tkzmQVjfe
9fB2tMpsXQuWS5VcEBL618WEfe3CeB3AckQ/NqVi2jpxZl4tOH1xNkZIWwAjCWwP
anOCfhnJpNIANOJwgrQ13FotvldScEZCf9I7R45I8ikafnjMCE4+BNyuXb2Y40ba
BW8/5jJK4EB98VDkCpIRcjS8Ni9Xeby3T1qk+5b+4N8k3HwbPhVeaLEkIiSkbj+k
ydWKtW1xkYr1imOBseEupNdfoXxCej1hfIJUCjl/IrVlNtg19kFl+Bm/nbgukDgH
mXeCHgx7b+UjGID9qveojY5W+vuIsZzn+2smQYj0LHAyUHZFkc9A55e+2VSlzaOK
lxFeHvmAPKvnVfo/hE/IOyuT+F3nPIhX15NVdmaneAAcbwBmoAYTxDBMfzyDHGd2
CqDgShzbzlGseO7p3dk0UacROslti1+gjN0Rt7lvD6FU4mWF9b+dfouSRZGnbVE6
1y66DjYIPQwkX+edDw6FsOYJob5tReriY2MtLORLeLg=
`protect END_PROTECTED
