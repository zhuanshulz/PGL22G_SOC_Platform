`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mie08jXosL2ZOal7XFl738qy57FJ0dxpE6oSuhrRFjbJCpx+etEO3std51T6qSN+
xAp7OTKKCdIBb/WBeCQpVz1Y+Aa0JHqHacICM4KzL/xEbgGDBiU5MD55HX5f4kVl
7ocBKkoC6RNL1lUQ658OiOWiPn7XSeT9ViOO7gl10F/MWed6yE/dS3cmFEnBJ9AC
md8+FOJgmk5t2egEX/eFR4+OrIW3yfWO8Rc7i4BsPyYHaPIxvWB6rWgvj8pPAoBB
XPyOTrYRKVduWW7QdSnHOq+SWFE+0p8c7czBFrZeLm0xc3uaCqk8Kdj0I79G+b8d
+kV0zn3bnNEwfnbq1wjCXVvKe8kvRZRsNN7An5OgbXy618zg5Pri6JyTOcvSvYOS
pIV1cjY5KelrR5s0itWHv2KfWLRewz1CBz7JS76Q8Y9EvxZfGf1fmy3GcOn58Ors
jwSstFpgC1m9ysigSsRzvcRBIuQ2u7uw88Z7070O8XTu48bcjsMd/GvGKKfpUdJ9
Qx8HuYZAt9nSOTB+Pyvrbl0Fs+UrXFXpdvCOzJuCu/pKgnVKivnHxfh6ZTHSi0wr
EUlMuRsIPFazZsNo3u1uPw==
`protect END_PROTECTED
