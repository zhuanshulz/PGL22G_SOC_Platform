`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8W0A7h8VYXAP5ungFOjq4rLK9Wizatd9ODtYCp04jfaoMQV286EERgWfTsxNO7Ew
F9ZIBJhRYXBReHMdn43CFBInd+IYVKq/rgTQBJXLDuXdq+C4Y+syui8nzbpBo7ww
H19dS46YyJCaOMlugECihAF0MOQI6lj8sgi3EV0mfnn97nsROxq70NHkjl+9gmYr
5A+NU84shN0q0CVoPB82ot+KiMMWRSy3mCGXjIgP6VXGoUuxB7hNnvOhG3LK006N
lsfcOG+NDe18pthqG4gXsgQLA6WHW5f59BEVFcHwkEhn3L84Z3Cqws+NtXnakHN2
PGowqsieqMRTzjPbq0j+DvIKCqIPA3p06B27dDHsgvzt8CkY026nriyrsiQBaOrr
dXn9NX5v8+8MgU2kITKEM+iuW/tT7FiKqNErDEc9yK9/FWSNgKI38pn0l2/E4a9J
`protect END_PROTECTED
