`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pScwc1kJ7MKwgYQfm9hmjV0m2aw06r+b0nD8F7oytbU+5NHMXLjxxPFx8SEegLV3
1hPfpPNNXwEsglyH18I59HoXlG9AG0ync1bdvQbtjewQUwljDY9rW7tUcsSAozi0
YEOr+PV+cFLBwg3Lfo85GnyF8ayqvX1CFPYNesif6YqhwG5SOj2jNpc10nvA6wxl
MRD4WtZvv5yplDDw3lUcvRVT3okCBNv+sKPiT0Yx0Wn8VkIEDszSydlsmb2989et
FK0uyQYHogaILewAKR1oys6U+GvLrGRajbhWQKJ/APUMYTpdZ+nqL7Z+lpuTW/o1
XuVciMXTeSuOMj5j48tvR4AaKnnJP9j9V/Q5JWAFzElET5gz8rrdpo4zaIP228xx
G1D6upwatJ73DCntNgIDttOgB9W/Pvq7n1XI7sRgcI+LxcePrTKz6Zm/IIaMkLZE
TovCEO5l2G5zfDa6d2l1OFKXL5hZD1MX9zjSjbn0i7TOM+JdsY4yO+rYPHzIHdnQ
0SoVyL69AmgDlxNJGivkKQ==
`protect END_PROTECTED
