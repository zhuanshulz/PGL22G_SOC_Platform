`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PHAPCuHhBKpQYfM4frWcJ8/MeacKnbJzoNQfPZCbNCjQmsjHtG+EUmaATy1SShl2
qjS0Ovw3m+p93e0swZi/3wNnM4E+k8l0IMWx//MTaKiZQumfCkjXF48WiSiyjO1I
K1ACTYloBg4+QYjiYQpHQTZwYcIFwl9gdhAWxm+UJaTzryCP9Xmc0XXj31r4uge0
yftBOxnS//1+1Bg6AkU5KjS4talq2i4eCQqxbm9VdxzbH7bi8strAsub2Ko2xeJi
rAqM7PjafGiVtSssKcYlt3+y0+Qp7R3lhSld4RzjBJC+ycK2zUqkMHPvKqVJIwzs
rZw5NHgyudgUD85pwiReTw==
`protect END_PROTECTED
