`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jK4eACoj+NVQOO/lq5fff9PUvCjkzIsxXmLjocDCAnFcGBIJfxZ60EVQJP1S8Cpf
FvItGkYWMoMAGZ6qMmfhwKYQkaouEUZJm4c+qRVN6Mh/fLkV+qVhvsSWrobVAclp
MZuhmFK2aImuB+aOWZlgvt/l3gEnemQcGU9msdTHKucQxBe2cQfL3gysIUd4Hq+6
BZ5VZclDA7BJV/x0zYQ6iJH6CLUj+iV1hqHK6OTB4DsYqSyH+8YgP2liC7QWfh1v
omF/h8thHmJ6vgSDJ/ECCGUllwA99HWxjybj1JStN89AA3YaNvro+r6z59dvItRc
tqjNj5zM5+TbiC9bElf+wt/uf0IQozcGH2hQkhK2BGA7MEV5DBk5c1i3uLGGh/RN
t3w1LC60+VQrZKbtqp6hmtPoiRuPQs+AloUg9IHqH5Nyd4f84ol0qMLa4F1Tmi/c
tcCKUQsU9QLftp8J55dXmrQLvXUH5w0WVonpYQFt813mrBGn2v6G9cLN9Lo6TeK/
ag4ValNoBqb4moRXsQk1Sz42VA0gQ8QFdtJLX/P+Z498Q+T+wQHFw6C0jJn3Vugq
uqXwvm+VRJieTyY9dXiTSGiIYA5WXGx1yDv6V4w3C2S3FO6/DwZlQlb/2kwxrcIF
ec3kiSUEsgYxvPmZtpq4KiwG53D/1Jx2YO8qQmYukSOCxrfS5fUZFY0cs2rDCBCI
gC92lpIE2XjIQm3p5LIp7pa9G/RMzJESk9YCzak2YkvVRZFkQbcDTmDKKlzfWk01
jsZQNMs2I6HbKv6UBoActGgyGIOWvgo2q99/Q4X2VrwUMerAYSvKTDnXgKWuKgbI
AKQdBBgtRUt+IPAJesJNF2dyi+Oa5cgB7GkT85zrmVHhaPIRF2ZdxPFjLuVa9P0F
uJ6TZAvczHCCMOkF/LHr1y8N8KsQzllNT1RvjIVSwioqZiM/GY1Bkv0zZNitE6fk
+ArUjOIDckeoJcmrVPS4LFBmiB55oQO8FROyAg0G6qktKs0gQx8gvAegmyjBgKJB
H/oaak6gfjtwU5/9FPOfrYL0bjcdnA1Lw7VYSRIQqqKA4AZVyF6gjxp9gY9bddE6
DT3zR2SXs5ab0frepYL3qgOwtBf3bTbe/x75vPpr0tOGBBzrjdBFmsRXvMHKaomO
BH3XabsrTwPHln75zqJiGNQ0p1miL1C6IQunyBNDYRmDfwQFY38d/9tWmS0YP/fb
OYCtGb2uei0sNSl4xglkVQHHgRf7EGBD/gFwuaHanwBZkAnRI6cUqmVaHrkfQ+Ka
T6t3coIU2sQz/YfqgVND0U6bePmqKse9b9r1zDlMzrXcSSvuqkqogDg+bm/axCrp
nrzf1qrNlZKjnRtgsM3PMVQNRtk5W04q29BMjXeiRl8USe96/hMXnR5+vfwjs1AL
iNvnl3mqdMsj3741I6hLw3P82xP6y9xPuyEsnlodY9A6JUw68SN/bI35Gvi9BqfT
6U7j5CLkBgrHhOffcGTInykw9acacUulBEIB63nayyn8YOnSWAxdwTZFLyRnlg4Y
78s2bDIQ8PglBcoYFSJZ5n2Q2ac92k3Gda80W9DD9FiEG8myzMCVypylQjLVBHp8
VNgqqA+r9K/Kl/rg8yJAMX045wQxN/8pcPpAI5P8m/lCUMsrXo1KPE2nIudZzNk6
1KRTvRCdrBTl+n0M58k2C3WPMDTNmH9NZFEt4ljg6cOHZYYhAlb4ZBvGeBYYaYHc
L71LqkGoyK5zmcteoEe0a/mxVw8F1EexKHuwXnjxFa+mQT7OylyThORcpLSnkQI0
ETGeAxmJAiuD/xE15JsrQpN6lQZTDUPMPp7D5ftnEFnqo8znGui6qr8BtYuo4Bmz
BNIfA1VfGChaeDMThU8K5DsKVjQV3lNh8oGhaqu2NFyhVfImh7XUuzQZ1Qf3nx52
wYehynm8WIDOh5Kyxyxd6piEOD8bxODI8V3Ci88LnccVBzr7UeU4RekqZyjXB1Gl
O4u7EeuuMb5pALS1aquQIC0Qoh3kCiXRpgaNNmc8A85VjcyrjzR4kYc22StNaHnW
rSACe8PUkpyFvFPgS+VxNg6Xhiws+QEARH7edcNnf27ZVwFnbUEtmUfFEe7Rs5Le
nOJJgmzAGlx+xeEhf5987935T5P4uOtlvkFhXGzL08KdXSbT1gIhAmz7JKCdvH+b
F6OhJUGn+AyPyllHcn3/iS7tkWhWBu1yRzhQjLSz4Y53KntT7kspiISsCU8yhqke
XaXCGWxMuNnBeN5VX+EWW6GoX5tMJbBCIFhsZoDTFmXvOLAZ2V3SqfnU+kBBLS+q
tds5WvJWWOscnUKS8wdLJnVbCdE147Ty/mH55AVsvWUE0SSsItB12Ul+L8WHgfTW
gLlwev7cGy4SpRsCF+2R/sEegkvrldxp6pKY7dOrsIdyBWb8qCfl4xOwoe31lbAm
XeaoVptXX9gxelVm5HMEWBpHi02LVPN2JBeoOtaG5I4psWkLi17AQRjFdjSWtvEP
QzoUTBpVxBNsbt2bymsp50EbAxj9Em3VWE6IyWTK34iGq8YVvUCiYwG5/FHdkTFC
52xrRirhwxASgK8TO3orD9b2m5MciQtnhSd6cVGAAYWEtLqxBMc4++BVVcoaVqi/
AZOnku3NzCp4CdIlwES6W3fXdJlPgbEzZMyIAccgQdTtxXEunrp7kMD/Vdn32uzd
5e2mUq0BbpBcyjpigDPaaqfCGZAloil3SJBqq+qwouMYNSbhEknVnoxM90aCI8lO
ONAcTedR5m/R2ll+8DpiHUOiy6IKu1ORWUFX/nb8gWgUnlVBkB/GG5NaAZ8CD0XM
+PTMxxMWG1VTFt3xPR5ie247i1v7pDRxOBdUcka5ranc8AuAaP/8EDIl8U7VM53d
B+LWNgc8y2g8esraRpbwz6UPvxbu7r/4QESxR8e+UOf2/v89DWjyGWYYBSxCpx9n
aqvH+z6NQJtOwzbAGkgrjif5uLTCmatWHQF/IoAs8F/bAqEYeFWPTAPKLxxsSP7a
K+J9re6NlhC4AwSY33tg7J13yggCyAQeA/QBchDVjKUgoJ8/ovutD052Mf9WDdmO
ghI0BkrSjKve/Jnuub94G6kw9pZ1ZHp7bO0IsMMa6/SiFC213X530O24OD1YJu/1
EbqnZEcpkznXgHzOl7avTinZp823QGgcXK4kXCBl6oqMC6pB+29Rg3oBE7vhKhBM
8Hk7SrOWRJvK9SGPKefnomViDyUakFdlWz/4RjacmxEL7qDOLat8SBDu74DWLw9t
ltrZ0mRdshMKUwDiFvqq600baS9zty9CVHPXR/eD6uRQOldcljhnh7qg7bZLx8xu
fcTyjn2BEP8ixnuEjCoIwtWBLGIjsBK2496PAoXt4LqVJHW/E3WIm6FHZiSR2BgL
/y/hxTg/abc/1e7zU+Us8xQjos/QbZX1uS0yHBw/T4I=
`protect END_PROTECTED
