`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s8/eCQVQ3zBuQdEZgnNuCP4w1e09kzwbpkHJl8RLtrfFo9bfeiqf7K/KhiqEPtCd
eqmrknoj4va0cSLQv618YreeHCbk7ohEX//plK2ydEpbvNwwMbYLcejwkvxBEyjm
Ki+6iEU2QR0XUv48YQBsCl1lXdsriK9rAFxC3manBiQ2h0vdKwxxMZQGwwXl1sR7
5OdaMGIEw3moKqlmZJzLSJztfmd/j4BZkh46Pnr2He469f88M2DrLDK5MFGcX9gm
YjYT/mJRO+aT/sXWVN3/hpSPYNPS1BEv0RYbYFH0Cm+h6Cl167GO5qim7SpojUE4
SBjgfE4sY4a136+n5mrhHqlNiOoTzTXRFL4ym4iC8Tb20JaxffiC0u5wHCSOmUX5
YmUOucfenGGP4hxpVihI3MJu/9aJ2TKfkS1TmVw/Nnhaz3V5mQr5mMF8ktY9Nyus
IakSgguPrOZgxQwOZfZwx+T9eUdqVkXfb08IVn2vNotyyfR21B0Lv38yKotPkX11
XsOdDkI8ALDNky93vtMkwlMPuOxmwj2lpDc2qGXsejNsrqX1T3+wPB4krGgRw0gN
+hCB0iAUPJUTIG1+xwTEfCkr24OEk9lVb7+B3h07vn5j4OCGneKq7iVp/61udjtY
oNwASW9BSRtGxzUXlZagpqhvYJVVmB3GMipigqTUMHx95Tcn6bagE7a6uoNycgcQ
yyQougf5qu8mbvc+RfW878wxiOE/GG3c5QUXkowJ5koGEDz8mGI3Z6DbAMa5u3y5
oIDo48xQBHi//0y+byMuGy61Awv3JW8HeJ+sQ7WFJ26Ic3uoMYjiyIR8O+uIiNzw
6FCmGlW/T2SpHGcgn9aKiniYgOYOv/pvfUVXQ3pbVbSRoIeSut6iwR7r9DOaxfw6
IlOnQu4+dwN9cdGYWc8tp+vpdSA9DAnMMnvjOwnwGTQTw2t2NDu6R5B17l06Lnmo
IDrCo5/SLhoRfwXE9xhidfGPKHEcQJCZ7DYxyCENkTluhWw9sQRCdoHgmj2zXTfE
JO+REYcf/3v/D5vDRfDlcl2w0th1v39pAzDcwEa1bL2aBJBfLhooRfazhUzCm3hp
66oMSRpyCCxK05BowpDxuChsUb7/dArAf7jkjzTWq++E6L0QvXrElVUg/TN3l0bB
cQzBkm+XLDAiFwNouKF+tzUs9sn8Q7ps9arEpn4MhsQFQpEfZ3vFWVcJbgc2djpt
uEm5gYma9LGX3vo9IMFj6X01a07wJo75yC1cRe+QVUSoFs2C22+LTVV8YIGeJWP3
y7KWMLo98hCVa4Vn1zSqNwNLfMpTUPTPpkjvH9Kn8fjLPmM5LQGEW0eaONH1l5AN
3JvsZbS8ejbHk3md6wma3dcguZz5jTfN83VOqEnP62Kkc9L/9AMej5QitdoLg02r
010ReV3d/d04uvoU4Us5KhD3dhvcC2zCu9DIRNJZ+uhtAH9Jn4KUJq4RMCheeTzG
+X4ICN6d8a0BpcskEnvIFE43tigQprB2QKfJo2QZS7lP7O1FoPCJP946NWjmsHKq
xdJjS/fzhnn3p4eswOoQDf9zorqwOEmsROddCoS26dfDSGYRSIySzIrSgZjktH/w
TggZDQnA8Vcl5LrQ/ttf3r5Btv6OLlSizQICdOJNAZLhg5BdHg2MsViFPwDCY/u0
0SmMbq0uH/OzGsyjSqe1J6k3okZlUGDn0cWE9HmjY6rU5ldurlPBG8zg/qyZ+LNN
bjCaXsPYh3lPu8+OnstIIA==
`protect END_PROTECTED
