`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ELQDqyAWtL22pSDZHtGIQVJBzEkQAHfdZUs7nX/vfzCePtkc0D+4SkGzxvPkhzhb
ShgRQ0HJvf7NKpcBXDKq124Lh9WukskxQFRxoX8NnA7vzDXQVdzTZjomNOKxiMjl
7ElRkShgjoYTcZet6GSjrZz2S0aHeMubYzeYjFk2LKFc1qA8QOWqUFCaY8RPZg/0
5eYIFFJnU4qI/5ygAgS90jjr42DeAzBkEW//gxc8azdeMWczpy4FN0Pho2Z8iM60
G03/MESxdhGLI9cHyJCNO9JbY3i+78xRtYrH2C382nL7lO8B++fp411tFQ1fHsyg
zQT/vLDvcABJYHHDCKenv0UoD9DZ7BVWe+SvG3duS5VIhq0JHWZyeA2fq1GehRdR
wMhXRPDHKd45x4JPi3TBHLGH+Xsp4T86QvJschquVXo2MVeAM4hV3M8jZbLl2y81
rATtfRGpQ1keyE7w1FMfkzbxr8E4ofA8E8smiE5QbBWkLwl6/sre2/1VdqA+OfMz
EcGgsUAMaeIOFAHQ+1Xfib6rHYLiqwKjGFnoc4jbxgJd3MgRsjFtb0CCFhLn5mb8
RuaEkDGiW3IFXJilzi0vzQmPKIWwWKRhk1ApwCWnu0tViLrtVKn2MeWPtK2GERWg
d245xvDqYNZNQ5em9ZIxp7qBj2VziRl7M24U3iJ6foTGHSu3JvjIhfve0vK7Z272
7qdj7QHPWpzbUHbpcVdqrwpZX6BJXKbDgrGqarmT9dAuRaWJ3raDKZpR1EsOJqsj
fbFQD+PabDTvVziplceOG0VaVrulGDv5Yx8W76ErgOZ+Ar/a60295pPmBKLo9I7i
uEJtYIQzQGBrrwiGnw5N0zxtNaFG+764XibftnWw8aAI2386lNhRhxF7/8EGIoC6
XT0kxyw4CfeTezKaQzQFjuCXWeItWMdP//FbvsU1coGiT/RF3OgJKgQ24WarNVX0
6KINPmGez+lbBOBhqU5zs39/OlxHzSx9bNu6XNlO6xeS71JqsmyXr52age6l8QGY
kZMwVLoSBoQCUZVNefwBoYK3l7DiCMSP7t+jLwP/A3hbcQgx+THgdR7TL+SSsnse
7BPNUP/gVP71UIEd2rTbWXQoMOayTs3eIwBzVUwe67HQiYm6aH6Iu/2cEU7VN44r
YqMg+RIJc3w3x0voz6VYThsH5EFVYjFjFuSEcHG9mko8sc3u2xDEmsyucoSCQVbi
DnRCMsQvLv5lKlnAguFutHm1a+TDELR1N1eY5b3bdX7YNHDNPneQ5m9vNC9l3eT5
dzsfeYv28LFn3VEy61z6iqEG1rUvtZlhjGSjWu1+CVDFiEx3CnR+BCzyvVhX1uNL
zB9jgPu00DP7KsuHQHk/SLDmwG06cVOZ14UItNsaSrGqaCaapwm9KTjhjJOSLmYi
JJny1apK9gzWfdphYh41x3BlU8FjRsWHQVRf2H24PlVmB3zpGwA9wd7IWovWxZ7b
yRJGEZQgnJ0GXwKGq8u5F8hp5Owg3WkcJw6S1pM5fmmXym60JhXPKHpEamul33gP
lWYNCM2dF2QiZh6En23pqXmnkU7OuqbU86UVCwuvY8iXK8tuu2vNJRDoelDK40fH
XLr6XKEwpAUwkffQ73vHXzF8k2doIuOaep9Z7247SGwykeixaZrsiSjJSPeKm0Yz
B+C8w2LIiJVpdFzQ5C+lVv2cTmTpw1Ct+uU9LQwR7VKYXcmAy7wPdMMD51VYqZWJ
Tu33yOBoY7I9Ls/ZK7CWnMpbaLbSM0i9G7e/Nm9CMvPp7eVwa+yUvXvZvCKEfAkO
`protect END_PROTECTED
