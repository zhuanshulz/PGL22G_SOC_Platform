`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cQi3qubi/IIXRHjH9ZD5kNbVvGyxehSfNFkJXXi3BfXWPhANol0ZL9MxxrgFK6H1
AMXOdxj3p93BYf6XAEduFc3wGdmx1rclSWa4Z6zjklsEnSF3wUZdrPkEmy3PCwTO
Z1lwhCUIy20VtxZ+WND/7cel7r+vuxdFJsFx4qYJvOXnq3We320emNqJfJODT5HE
frXPYg0ny2et42Whagwu/F2rU9DlgyeVILp7biPAlfcA8UP9ckbNUUMK5a7KWwIF
+tB50QXiIqiA6HiYhIBcltLZhTDdA3XiL33rfQmwIQsID85oCJD0XNCMwJjReuuW
3N+JEwJ897Q/SlS0RmrNEGr7IsOH7DaCrXjDTuku77UIH8f8GkZBi26S8apt6Ipq
swqxO++VI/2wa6KzM1Pwe5gH2HDVgSf9nCRzCArCZDbCk6zwNGXQTVRDmOcRruL6
EyQ2h2gflMxg/tTX5lqhlPE32kkbmzLrY+yewy43n7i6lkRx8XYTz9Er384VN4ku
hIIbKVUXrIuWfiMi5CYKRH7ddrXFRT0Vr+qWtn12OOfButHVKxI6tjOywdcKgBRT
Nqqu55JCAgqhBA5delFKf7lR0gd38oYK5Hw74OSGWEYXWb0XrQCQtOV0lrPUvq+g
ylZyrgCy/UBGE0pCH20n/OTZXY4G8Rvtbpvt7dqhzsoVNF+Zk/mL5RyCgjwiFbhe
n3SmnZY90WOXrZ03R7/nXhwkDb54uKQG3uUg5k87p6+yVOteXGpPJDzdT7Zd461U
UM3smBvCQOkctS3I3mXqNwlQSvMkaqx3/c8rWitpxUJz4TRODUD4Ny1Q1myHpOW2
zEnCYMp0EKNrRZvzPRfVTLjLk0mhsLTXN8Lmj9yxJLHunaT6KE+OcoPaG6QAqk0v
3iTBg+rgAAc52wLaRfZ7Oj4ARgirptA+pH3+YNo0UMeYurttoZigZ96L6ay0ymNS
ll9mZXkxgQeL+g7u+dHQfXg87HX35c/1lgPoWUwNrtQVcaHSqEORchPDFSRt84rl
uVVpotdnQ+0h5jo/0gk5K/rH72FaUuiRumysTfPDNuGlYJWz6nA1lgKhJXzBVFD7
5tRNjw7tx718YdBZ6EZliEsYwkOxOx9RHeHMsIfxkdO+XLiLgoHkf1Qown1voG7P
`protect END_PROTECTED
