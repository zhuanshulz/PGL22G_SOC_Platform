`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0Bj1C/pZob9Qs9fJcwShsR6wkpLnCyT4nhGgRpd+i4QCZWnVl055kj+M02+hVAu8
Ms1rwyPA0jfD8CZxk+0eFFaWQaK6MS5zUCBHo50vQpxGMmuvfkLJGd5jezyiA1Ba
izP8iqEUAk3MNV/BABwqYSWeYY4iCRbSvVU47oPa0prjJ/4SBuvRq6B37kn7JZ/J
gX3lElSKS/wSnmM0yCPFrF93o68Eh2N022eTzIUxsSDwKVpw31cxn326Fu/GdwUI
R5ZNZbslcwZ6C93IjWVfUFZ3NJemTWfWTsbeUD4FHvweK6NerOdHLGY+twkk55zA
PEN+V5/Yf0ActyU3fz3I4cg8fSqgdLEnI57CIxF6Edwbwqu+1qR57cI/JkhE+r73
ZmhgYc8y8i/r8GrU47eSuDCAjgFehuFTyEzfu7iQM8/P+4G4UrzLwOiBVk9uQnCh
sQqyInpNbIE4jFzyjsEvP4KqbWmXpgQ513WMC34afFXnO4BSyit6EoPtqKbF53VS
Z5ijd+bgDJJnVlrAX3R2A+uBzP2xiqMfLZm+tH/dFZp0FaxP1me6Eel4f/eI/VuF
Xqybd5C/EvWy6z5uPf8bfy/vpjA72wTXIVPeSR5afyeAAVPM/grWkQ6z0AnQ2HIf
kbgahVqgjOGhYwgqkSM/04xsLbVFxQeAbFvm1zjUQeWFoSzD86quDfsvC5t3odY3
096nK1GrXY8yVN4uHCq2kxCoh7H44I2DmjUK9jvW0qy86x4h5EdZ37PK9TDoPj16
WHk909Uw6Df+M6aDGLfj4DBWjWma+CAaJAlTfZ9PaaU1N7vsstVhK0w8wIl0M+xW
kNWKHZwO+98f3TeZxuEPg77CIQzxA6RATRX9nldXvJil0AIUYIypBxOCL1kbe1Y3
AaZ6HJk4JSP2mx7sQW8sQXnqNc9bRQSZ9yJy14moONdr2Nl+5R64ojgfh2CMuMhW
IoXnzE7LEmNZ0JW0L4diXdYEiYdkeBEu6EosVEOGn1wXae5vmxBFab7G/LVlcJkp
jm+oRQZphJ/v5MMtWH4eSBXz3/SE5kDbz9+2c+sPQnFNAr4KJLx59VL+diPDYmx5
XLaC16hb1ytAOxF4DaVPyuxhLoLfCzQLG2BO8+Cjh2JyNXtCA4qgHCcUiCJkZlKO
V8fCnrR/cIiF9Njc3AR1dVX/EHDzfMsNiOQ08x0g+/QYWTxFJRD5YkpDcrE8OkLV
TVrIYDy1qtVihHIddbn90OkwYpqYtoWERhyCbENvr2A6BrWFgUiBxNtl6F8Yj9a6
7zRnKMi6Re7e0gi8ipzC27N0DegeURqIpWjKiGGgPIKIWyTLC/kfcnJG90YqLuCl
+4FKQTOlVeCS2+FSSpeVFWtTo2pzuUDJC9J2TtCMml+vbpzXPD9/6p9kyuAMGcOH
t7Qd28QrxuujPAPZanTioqnnNjxogI6qGhOO60Gv4wQTeKjKZ9P2T2JKbBfQRPOX
dHGzpcRSJOYb5xI/lNUqfowFxPWEm3jLVnNEVc5+WCPznkdnjXteY9F2y/GjDE1i
uZ23TmPMom25EyZI2DUq/JxIMMHeufXh8cu1AcWpV+RLvjDDxK3CvbMA52EDM1e4
+rRmUAXulKgMpQnjvvFuU2SpEdTyiezxi6DOD0eCXgv5CHgbxzhNOJwfZoAZAENc
we6gR8BMr5s8orLplf2yvi/6hw+czoADhYlYrf7gM/vOlotMT5j48COOM2wPeP8k
DqVOfUMCY1exqZf2p3uEEom41DAqS6CZ5vOKHjBA7bqt94kI6QEAKMi1d3JvS+Hh
NiAKp9ZpFncs4zdhQZlk7A==
`protect END_PROTECTED
