`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2/AzBR7LIYJ3QEX1zo3qay9QpDuNQfsnWumNCo21gThobucJmBfiNjmWervqnlKB
bflZwpR28huPP/ctv42jKFuJRlxUi1r8FZ6/CqRxkCw3Sj5PXZ3yHRDzul46bY4V
Rm3Y7IZaqwzQDempt1v9rNDTHOXYmZzKIDyMeXbzE8skMlkXec9NAGRPHEQfk3pd
qVcq+ZY8K5CeVWaP2HC8ytyC+Yh6rRUNQBs86EOWxr9d84o7bhAihHe5R5MsWryb
LQBa6vXkp4DlCUXSR71X2YSQjJFGlqVlIMZ4XsWAt/G4R+pRYJBPw+ebjKjV5vW+
HavfmJrA/+311VYFkoZDeWO+hlPyBzkIfRO1cmOnsunYp9uck1DwXvtkTu9PbNcu
77PXuhTg+KNIET/jK+2QOnhbUEFF7M47ORi4eAeJ9aLQWd9CXL+hdIe8H20CELg9
BZmBo8p7FJxWuP9HzmNs7P1P9b33Bgt9QzW0s+Pzu/eVNFi9xwrgXKoP39CNu0Fr
FCo/9duQyRg2RgkahSBayvFqalGeICSYOCoQOA35PedefGmdUfiTNNGBMM0A2/QT
O09lHdjNaXxtplhcuFt0UQHAAiGMwvfuHSb8Nn6v/HMzw0DwvOMscdg3q0CrqgFV
59tagYD3ttziJ/CxZY/54nJIEhfPbgoi/TswNVQCDFPM8mZlUBvz6xMsWjwu5iCO
Out13YRkHgDa98E9AJkAyMFS/EF0Db0UNzm5Kz+gmrgEBovVrWEoMaRVI9lc51qv
hCDbuETG7S8T0hCNecerAuezvI/Km4trhXhAcmYFQ+gjptKr0/5E/z1wxOhrCbIu
uHiMkvq1+4r2SwBFn4n0rWFtFLjcLWtMKgzd3YOpamUpx5qLyYKSYNIXistDUV+p
aw+++JCcsTHo7Vv8/Gjk8LLbmqcNnTzmRW0RcCYTI5w9zN6Bx5nx/vkjmF64SxhA
suY7SDw2qXQOPveFaPzIL+VRswCe+cqc1MouAIxzcNPMRTOVvu6IHfVrHf9NZrjj
wKuoELRzz2w6956j9Pvg8aE5XVLOYo8ECTUs+ckerC52vQJSCG8YeM4WtGJftRcq
s0AOyt96/z63IGyJb6mk9cUDhOZXJR0AZGHOfbMeNaAHi85mGGZlvppeMRnzTjlA
lhq/kCP3V9xJd1tujFgIimmJ48+F7SSZ5Bv3mUjoLYS5TMJzmIk05t0I+f/2Tc83
jFPVRXXGrfD+a779MZuwOpu84owFac5IF0FM44FQeeS9sTJ3STfgDuOBMUx5NGgA
Raj7Us2tpvK92bekkWdhNnv/Hv1AyJUYPtXjNHXddE5nedMgMzAXS8K8wjU6e0Kd
23t95OpW/Oo1SRqfjlwTR7/2cj+CWLAzgfWm8XP8IEXv2RIEdu1ryr0A5neIGqQm
wa/tvPdt+Kj8hC06wSvJtyBGB6/USbxwwyB2r0ylCnan/0LIdrZghB93lvJFELbn
ZatvbTR42cw5udO85IAV17Jkngxu5V332rmzii3GRcrAQwAQ0bwYIWrW/TEzWNJQ
L8gQRb0p85/+VNrLD6S/fkL4J1BbgwMqzpzkzg5X40Thcl+t+ACPTJlBqEk1B9CE
sXjCR7wW1X/A5SQC4O1Bcb+0Kbi7704zZTf4JPJI0iep+lRNNmG3EZnTlH4mUCML
8kC/KH9nXxByDIuCmd58a7Fe/r6XnI+8xWYSdvj7rHIU/03VKlsmurYznTBY6LL/
QaFXVz0cszG8yDOC3GUukxWKI/uDI8otKxvu25YYF0NlpWTGlBixnLt53vMOnXQV
dbJO3H1xzcXqzhqpA66qXG7Jgc+vEQX84EenjoOR0ZuQVVt77+c242QC/H7Fv1RF
nf1NTmC8w8UhcI2B11w8Bb9GkpkKW9huhNHVnuQqDTMQYlfJmbV+4S5sNGGkFSM8
fev+A9o4/8OAJUY6FQQdB0wk3Ruq+G05aejAebgjDSA=
`protect END_PROTECTED
