`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d8/zbYTqQYSFrNl394BfLIHL57NypT/HrqOfyIuegNLleqRlVWmI4iv7y+ng84Du
+di/NzrR4gUNZpQlfu7fQ+SDvL8qhGmWL4LXO7ksj7CFHBk842ocUYmVXh7vhXW/
3GyrfCLHfsoe/xgztr8JX8nveEHXi0GbrNIyNHetbogW/veeGlQQ+Bx/YZc+Q5Qk
CBh9jBL4sT+UFFTLBkIth4ecNMt0rF85pvQPkYjwIZONEol8Cnpbn3tdX/E9VASM
EC+z62CjOwJw7gPHvDK8cyG9R/GWjD8GAmkYhCUjeCpHbUDhREhgGJazL6MT8uMX
HOEmkQwG+4aq9B53oVnrqrmKjyB+xhdk/c51YaRKbsfxUaZGnXIbDnzR/mc3PSp/
8+c17RG2sw2URdrlL3jOXY0xS5SWUaNXk4XSk+MGOgkQB4kh1ak1xQIJqNgMd4kK
ThBuiI3sYFP3SjIBU44AMKg+ylllAIYAE+qjMXkjyzD7xcbO23Nqi03G3Drs/lGe
Iut0MwkubNKJf7NqoAKWp3wvSj7Y8sjau+DBhbli09BNCpntT1sGJUqgURb9I8CF
8SuM4KentA0BSWaftOwEy++bB/9xjog2Ao+/ueFjTCLYP5QDyWyLcNip6mg4myTE
/3RzfUhcifxDrcTWrg6+EDm2KRlgpNJ/QJwCOWmv38PTehMf+zEw8025f29NcxeP
PkvXLStJiMDq7AVbXyBphTX5/LrKB/RPZ7fI8ig+7W0=
`protect END_PROTECTED
