`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7xY9AvDaYtaCk36pHGW0SKjvnMN1NzW7qNUMh/oF8rIq3XBPucUiBX+Bq5wgKPfY
Yd/3qi15EifC+meLnRMS4ETZz1Ke4AyXgK1nunIDhyTlbpnLJbDlczv1/TmWOPYZ
a3uANLVs35WrsADacIM+KGT8yD0tpy0vcSvyKJVu7f0/QqRre6b22NNjC0CoQlHt
DclA9897Jnh0qqUtE1XgXzQZ8HtakT41K58NgBnZjdtT0gkKOy1YSDmd51zfmvYL
aELPYtFzf9rX5w+szGyd18V0FzmZ1NbYkVIJkbLOI42hX+66o2UXKRUus0aEWYIa
2FSVDTSHuaW7Zo5MePvWPQ==
`protect END_PROTECTED
