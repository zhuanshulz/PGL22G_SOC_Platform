`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DpQUU7HUweQH1zfh1EXdzFGCWTSxeXOlpqPpO6DYkvmGrOpvpsgVeLmLc7qoIcU8
watmNqQwK7yV+uNd0x/cHZ1UNkFbg4OeaFb4k8V8F2grEaX8yflmxBzi0+iKRhE3
AIVj+pR95ontByw5Od/1FpBiNfPuZ9m7LSh3/rmQZQHqWCIrzKLudTf2CkBvetfU
F1iyaiEVpqlOkDwiv0lD/LVEmL85uwzq9iwluAsIQg6rsoE3g/5HrAs9bV0hGigf
POnFdccnC9LlyfEp4SBa2a7Lp789/2m4fxucOVbcDctxhc5mY94oeuCndN+KdzYv
FxbosBjTugGKLEZpxV7wLN5XdSC5bZVDfFB6NeUe4T1zH3pk+dzzrbO7nVaXXBSH
VOUcwfFY1iQZ7b8Jy3a2MumLYoZvQnu+wblDKxRcBR9vjgpSqr39j6k8kgq4v/8P
CMTuI4NK5Og5qkE1dUy3OkbvTfZKKaYSCJ5lL7SniTjbon352hBUmsQAUifhvrGB
urcG6jL89Hr3dqu8GZWIRR5T22nMDGvE7TN+WefHPo7DE/Kkwrtq2Vx3UIWiXMA0
0etFcTyO4QDLw3yRijhEtakLAJgmVKbwYZpnAyxkahCBgHBKkJIOqiknA5kf1rKk
3cUSrqNt5LAOhm2Lrbn+g2AzCVnYzoFxnu9yChy2wgtCnctaYE5RbXQqREUW4lpc
Hvsu71dzJaagaDmSyWlk6UER+LE3iR+uEaRvbCcvMMZvXsBtLHE4j19AIdvbc9Tl
MW+odtNFyN3ESIu271xn9J/ZRaMcPznRl7y/rjCOdE6piZU0prgScmaMcy3EUhKc
VUxcUjSCBoO55Ww0XJxn9fpcS6bQGaubVdnt9BC+mSPB6+O7IfYGBIF9gpu82JL0
JOx/7/SoUP75USoZnP/Zt2py3BJpNd11mz9nzWiHkyy1ri/UNygq/qDfwyN/0Xhm
P4xxAFDKyln1QjHNYAlAncau7yRuc0FOygJt6Hu3Lrw3yC4pqHL/Z51OBlR22CVX
SBKuDlnVFvZLoofE67l8AXCEFyCq+lc80mhtk8muFPAv2DwcQGFHx3efYp3UWYFv
hCUI8YIfFJlH55c6f+LRFC0/ORA52Xt37eT3C9wRItpr/VExQ8nTo8mWSG1YlEop
j/8zXRKGOUBg7URMZ0r8Nsy50zQCU4RrD5vIz2I53zEEnoLuPXgVOR3faBvNQbNC
tRwxLOdNQB7vThgbl/gyQQ/YxjvzgnN9YoLBiFedx0gpoBflMmT4KcTWMbqrapPE
lH7MfQWrUdvgWO7StNuEw0aMpQfnlN2XEnbnzKVYgTDu8858DcNuTQ31UF+w0RBN
LMptsDO67QC69UOw7kRIDvlhM4hWcT3laQ5knZJuzyfzHPxRviYE7W4fEFUz/RZf
7v4nvc+qEO7cI6uYQGU+Uo7aKlVbOqH3HsOCwdCwfKZF8Orvw8ekrXQ+y4j6M0Fs
8nUXxP1mFpVna9OaLJz+rWABHiGWxa598xlX70uDYl5B2cKfZ5B/AfN6cisgQYUq
qm/QD+osfVAHOKk1cdbK0lvuIaeF/97z6FtzfSpxriwf9000clABEJb2NUQPDTEE
Qfdqwvt2WzHbElYgnA2g6IJphI2+s+KYUgSSeO8mTG94Yk8ydtHFK+FQe6e+XG0K
2iqETyZyPOzFMQFYtg2O5ha394avC3t5xZclpmbMHKJ+c0RlJqENGkgNmirK0itD
hTkSJLnLbyU7irxjpVvd9sulrz2D/njhm909PSYRhTQQnWiti+zLaor2ZUDtvgTi
3HEHLErW9Tq0pYkDwbv7An9t7xc//gSlkFDuBGoHlUtJCmdFtpqch5yrxpdgc0ef
ikDm5P6NIGJHh9hb/5LQvTSnBs0XmtX5fCh97v0PRGKifEnlxyR71uG4TqGedddS
v8BNAG5H/mwntZCvs0Gg6UPeeoMKxDeDfrKPvnLsxMMSO3ZYbeR0+H5rf9XlrQ+6
/kha9NKwK6xMGA4iwGmMDsfGc8nz/+mwzWOD5NnY8LkUktdhvzJEn0uI1nXCZr6i
k+Lk3oDkJya3qdTZebRkjagfI9f5I9LNn5q1M9cfxcAO3RF6Huu8cytecS1GKD1q
TEvGpW+gnLRpupAVTayXWdFIXqALRJDcybkIJbrRFyVFsbkgXg7mRLNL8tm77fEz
EDBeo/pvAUZnIAWdFeu3t0rTxtHcE5cwM2PKAqrBPG2TSCop0RIMCVkEP7hJLbbp
nNTdfPWNzetjt+AdU7QZckEQ6SS+kV7OiaHUvvJ6V2+LfHnWYKBdnVBL8dP46Iv4
CLADo98xJ9UPIYMhjB0rJ+uSJo1H4McKXhYee7Xpo9Jc4AbzI7aER51IBtzHsX4O
84xa5eyP27x2jVCv6H9PuhOrkLpk7+evG4i+XrYGziKUHg6RF+Cn4bxmI9oC5b1G
6YefQZjmZTcwS7ALiruAJAebeoSsm9j4WEcymfz46nBdGJU5xPtBxU87+056rDl8
5Qb768TOCQnqHZQs9UDXlr1yPQnmFOn4ZgSRINZy/h0TNunPmcLqHv9Dj/vGMhxu
P5/OhloVlm/bg/wjA8MpNW8gPL2+HNTbUAjW1IbvyBvvpW8kk2v+iNB9gixbFSyS
ioibUNO4oCliiXkooJCGTB04ZjkhnDKEzXwdNHHAg4/902YzYoargVBWnq+RUvGm
FkSUnnh79Ofl7f02G/UO/g7ltA+aCm/2MvpogL+OKADDh0+klIJu3fKkHYXAymI9
keak1oUeifWp3/MaAAs/81+m7JO9mK8gqjOHaJgWN9Q6kjXd10DLyhrGOwKk3pWf
dK974UyMKNG1bQ8kyZpMqDvcXwatN0mkzsX3QcGT+OV3koYt0yLPDGkSAfvRSvte
zC2d8t225qO53DJa7lkiotzNadqtAHWzLQu6s4stiJLXt5EluPQjRCPeV0+T5HCL
vjUBaLekAVoAYlLmXe2NwbrPWyed8m17Nk9c9dkjppSKaJWyi4gfgv4J/45kvEVK
HsoCeOm7BHV6d/ldkR1SNQlgZ0MDqLBGo7O7TToShqHmFhIp2ldY+RuutiVxMSqT
ri7jgZRYpQp4rU+41X2SmG5Mbl/zrwpgsxBA679uT0UbAIujOeCHUdippELVS9Os
flZN+f/VqJ3ocOmveZmgkRq5nuNqk7UruGltR0jhLABR3QLZBHbG+hqug4QmCh/L
My1qA38X/ebVVQo6bMB7XLpuvYVUc70Sy+CuMPdDLx75IxaNqlRMK+j/0FNaMwl/
cAQxsgV0qYFvrax6LXi3fFhn6lOd7tbYPYFGwE4+v0rSEqVtLKECwfZ0Xpsumt0b
f9SuG1GLL5e11A0fDl8uF76/9drW5Zd4kYB5wtXHy3yJpCfRFn1w5XzVn7WMVf05
A9tbbHd0RXhADRltf7ziV3YrOHAAC89RMk7Kdvl3qZziVtFVKHT0Uh2uB2Eeo6Rv
Acn2W1oNuzGUm2LwHyCBcDrABoKQmpXk2opXN2EEIr9JZJ2DVjNjh7Sg+XNjTue4
0k0RAB0aKWczd3gYZzGOkLjC3L6RXGwBGO2LOqHKk6BnYuZjUZ2ZC9okWRIC0kkW
xFlF2IhVgKGSm7oKrtsvXJ7gM7f+sN3pba7dvznsYvfJyktD1r2miNafnH/QL4Dr
ZBFmCul6xZu4ApNJHA/AU51U58begShBy+oCl8gS35polGcoKyS72bNQCN77tOfZ
sTsleyNDWKwu6EIX1WH7TynB0hjHKxPgmK9J0WQ0JbWSV3AIu20bpQbg0kfIsp8l
devH8bLV25kaYEUVdXLQF1eutR+ZgCdTZkCKbdCwNdTRpvFtXtWpyS1fb5kEALVx
PdF0pyhJFjB9ELn25NN+FAdSk2Hjhq8eSJQShE2nduWFRM6UscXz9rI0hxPmn2NJ
/jF5rFuo0ms0S773FAiiTshTNmiJnNay8rYZzdA27oQWYn4QclqMtQFFLIaYpc8s
ZN8/GTXKVGD3QmmiyLJUxgN9QarJ/gjv5VqsSsTISlFSoNKIDhxpvORRyRRBnNKQ
6Fz8GHsE7uyB3lcmJCNGS6kEBjUOaMvZ4LAI/49hA6pvO0jRbdHlhO5kV/+XY1ey
2IpnMov+WwdDUUvmicI/lcIBmkYiq/V8+a/YOGtupiU=
`protect END_PROTECTED
