`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6uP1LlTnEb7QQVoowEAV42L87Dn7Pl2Eyujbf/oq0j7t72nGCSvZ/aQQntJFsn4k
JtHyD98OzKnNW5qa2tzn6WXSFMbXtPhCtXcUBb2rQ2C1rwgBEjgdIwTvPd4KpjXH
Kdm0/ZYVyQB2As95lliT7oOSI84oDz08+Uny1G9BqpuLeN3uofwdsAfyQbpiA44q
Y1K9Mm8bQ9dQIUIbhfnt10QCADsQ0ZNGGBJ2DvypHvBb7IakYopP9C3SDxyfOdNz
mhsCMYXxZhgkTuGQpLUsZX2NlYyuzHzcn0IhE9baQZEk3MKb8fT+pJ7bn9Gyf8as
pJAKcv4dHxgTUuHOob5edixxv2VceUWkQjYhKXFB1z85v2jk/OrsPNwBFzPE8t44
PulogzcXCGPXiSC3snHQ0JeyI08fkI8hOloDKHxLdo7Rp0429Cx7wsngk62CqPgH
AOnDFlOdy8BzX+TCijbeYRXSFon6xDLp2TbPt2fnG1E9BHypSqDLBw9S4nYUfFM2
96WfPGyY/nKwMinc3nilr8zvdYI1uFSMo3bMnbnbnH8DNj/M4fcDNky/Ir4j33Hl
iCzU8rjyzALuUqESEivxuWxeb72ySlEGI7E2ezHfPxtP7kSYMrbeZm0Gsnjwhfhf
L4jBexbHsrOlfxNHVE8vgRp4xvk1DXlwYGMOTq5Z5n11M36L9HFn7334ucLEr/1X
BozYPqAsCIkxIgCTa8k2Ytv44+6ziMK1eZJ9O6SNaE8g0gbC+EoxLbotRX/7Jx9x
A5oOPh7FaCmE6SOafBLoGx5hhsP7LZ8yodKSieBzfsA=
`protect END_PROTECTED
