`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aw4BLxsiF+o1LaRxAFnxBSYgmmM/dB+aAOR9Ux1OZQx00NclGv8OyWc3UBSr/U0b
irVR5uplFD/wJOLrMHJiuABuru/J7P6bo2p6u0OGI7GqUoztXUvghbdlObGkGWAg
ETKvgjDIHnkgPxZPm3Erf5s2cs+Ar4Qop7vzaw0Os69Yk6yy5ogGxbcaAEo+rM1B
f7M42lDyqgAzBkvwg2eHBhwUWvCFXXoO9O/VRjnAgmJM679TodiSjpJnYvX2c89t
ZpnGHM/5CXs06VQ1VC2hn9RZtsmAudDS/b6ikuK0bEKG2okNzWodsXV0j3ytOCKP
Yh11u9TFxjfDxf2UX4rrIZ0uZZuVuDbiFvHky+yOzulq98OE6ijVOIZbfCY/4e6Q
Fply46w0s+blhalUaF7ObFG34HtlZHlb4fi6lbQJxhGu9wl1VQ29UlRs9PxRPsv0
uiinKudZGLkWMrCTOOD0O8WwI2sscgRcGqH4W/NqSEFyyvpXrptzijKQEZVnQJuI
CymCEnZvOSIWNSzubrRgikFFWAV7Xv0K5anB1tl4zfvZJNRRWQdskOoDU1wEfy8z
slNvmP4vBoRn3VxV66UUypL6X3KDkRj9pgrydN1awJtfnzQzOKhQf8kVhr3w8ASh
nF/C6dFSUCvzhIadieEsrGrJydkgtUY1cjELL19NXQugkTlJo8uKwwFz+0HwzG+w
tTHc9kdGeLTdmEzBYqmTT/EpBfq3qItgBiLpurE13CTyK7+l5EnSPdEVSHRxG5Zn
ChgVFHGip+gwdvr4+8T0teni9RlgnwGUrBuovuxZlihCAKh7MPS/Di+EIYsY2J6C
jB5NK4wj3JJzljD+vcmNQRBR1ZL50qRuP9P2kEVLqzrNQkECjwFxLm1xdb8Xy7bQ
uOXa/aT2OphRO4vZklY+nLWgeHiHlAupBvMs/hh8NjNJdPmH4IAKrpdoDngp6ShQ
SNgkGhnVGVkbsrB49K6h0fl0vDIjZS/HQlpIRnV22PNf4jeO8GecQnWY73G/c8fO
rieLcx/6CKtzvRe6K+IFCiq1R6hxA+hjgX96V48/bsHK7SDBVrFZ8KufOMdHHil4
DPySmVS06OUmC+3NLgJRz0ZystT4V5BvIRPCcNo/qrbAuonWZl5zudxYGXSwCljv
SAyg1M3xctSoDJzebkuwZvF3Q8JsHa+tQGwXKpP37moOk4WdR8s+3JXF9ujVURi2
jzkrCn86XzfU7hJYfBoN2rY8xIjHZBT6eqVBBxfAyIJWUCOt6UGe44bj+0ruwQue
LxlHm35q1wvyPgBH/Czzxc5cvayS+Or4YtpfuXVokupEWSrhAs96Ccd31DtKNqf6
vTH9fZuehGsSNy2j5+hdKaWX2O5wDyaYovfdcKOjn8mDs0vNhpItwbZrcL4gmUq6
glvdceee6cUjfwyBsIBws98pRYibYZewXe1R3ctWE0iqW9JKFKyIxJXErsnsDUG5
4pQJlr6pFnp6cU1OdMS9/hGEmWYm8HpF3r2k94jsIbmq/F0dPvgXTM8iCBRhy8sS
wLCeDX3Q9sqlEiO7ZDKEEC+haRvoCzL6KhWTnjf/R9aCTMnFW4xyUCM7TgMPLU9w
zAaPsG0IfRix0fBn8Aztpo5JcBpjiHWvDXhysoDy4460XO29wa7y5QxJhytMWXYn
Ir1HxJR70AlzgAlG437KNYYp+uKGlGk2Df/MRYyRJaacGHO91t7Yny+1hjjOkm+k
MEbcmlKQyDCVPa8xmZsqkFhK1Vmy5Z8CnxNEdApuw9lkqfIrYyO1xxnuzQwBCX47
nktnUd4TTa4IlkXKixiVAP2qrYuU/PuaJPCoaW8mgOOzeFCdphXc/o+layZTrVXZ
BhsF6W/gDiZ0YBAy+CfZ0vHNUmEbd+jdO4OCJEfVX2qJuuflsdQK0ffql6hCZzmS
pjF9tnauuTXhwP6U1wvp1BHOSiCHbB/WtisFeA6LZQpkuf+u7DVSTWi9t/gi7tC/
8oDY9DFMi+qWYiox47bEoC2yRRH1ohkYjPUCkeIUCvQl/76snbje+1grM01vmOyj
x3yn5iRzFebD0EXgghEcHHrKey9B3ucqkLkF01zztKDWhWHV2CDEEn0SVAcFfLge
VthkCOwWpNHyHgz0eHwGtr7tPxluLIn663NHIPjQ1KYdXKVe1m3URltiKh75chTF
WJHOJJQkwRH+TRdHaqVo76jaEmn9ea+xXNdKQbhyK27pwLRx1icui+uCFu88NFVu
4ofTVGN3U0rjVjO79v3Z6NTLqKKhbDJjzFM5mcSS4UjHTPfjr2qSrsgohaqR8fIP
9lz8chOFdAKdDbYAWLb9JaAfatEcMDthhlRInfKlaZ5F3ZWzRy0LzpqT1t71oGmW
eG/JEI1n7EGhbaLl6QXHzcStq0ys1jfkXVNWISRw0j9BjhP976L7hKABmyBpFRJ6
p6aTofz0kTfPmoGG3Bb42cuw0/V379esM1bR0mZA+p6gYPgtuKzrEpfr9X0DTQ3n
tOlr9blAn5ym5yX45YwHsgwHn25ENU1Ut6k4PGESaI2/PPL/DhrRwgiO+IZ2H974
BF2xmEFDaayydFdnkwUO7hf/h+4rTS89PXDeiUqZdf8QdcMsmOTYmd7OLeF/IGHe
OFu3eOuY2wpLbdjIBgDxL6xWpJYsEwhA3Sn/Yk4CT5gDf/MB/5xdafl2uOqGxSGn
J0OiSqVZ5i1E4n6+Sm/c306785bUHWP756BAHuzleSRCTHMvdnqHPUKxehd/huNo
7krw93vciqGZCPxCjWBUAMm6wInKBvlxJSuGGrVgLUhsaafAN2rv49pU6zX+1rCS
MyjMwv7JkpH5cFrbmkKXG7UzLJI9cQmTF+KKmbwu2NS52KhX4QCcStqI0dtb5Gfx
X+1D9SAA1QZEojIVrPW/nigW6SMDAO9n1cIQhGhmSxMxZj795HHh2bTDwWygqwSU
JC68qBiLAC6btb1Rm7wjmMkdV12v/3IwPU4bTo7tGmOECJ0QilhdrKTXkPmLCJy9
TigA5C5CnD2CscSV74UswCjOE02lxILSGUVefXS+tG5OS/zRt/XY1WTRrYFMfF0A
q+o3z2DsKzSruSIa4AX0EnD4sAff6Sx+U7qZJwiDWbkFzXIVed9Ns69f7oUAWWRu
orSDS+Pme0mSWDspwsMO7aluQYt4ymjNf/OaxQU50dKemWyhzRPgRpz3hvReCDP9
4DCVDA+G6RKx4fnO0A7p13DDLSylV+1P90JKVYiMU6GyvynNK1s4RXhH5NK6+Lgw
e4YPhFSi/MCk6Pkns6QmeCqz2uMkHtaRPhe+DT54PKQLh+fd7lCBPKA+m7iUFkVw
o5n/P8kPj2YTGfYoP8wWX/qrwVjQ6AalanNtIdnTbyF/JZW8Wv2Z5iaMFdfe+XaH
qTkDwBYs6HE8No91uhqdP58L5OBabIfVVwFwZRMzVQilBym4NP3UAA3XWcAgUreQ
Jo43iIRoqhw5q9gYHEMLrJ9HaquatWNrN+OeuQmUSlUfWADH1W9gXZS3YwazhFy2
CHO1zmdQbaeMeYQxViYyqpr2w1hlzDwVSMklSR09zaI+c96zaLgbNwOtgiq2kje9
EKT+N5CKIXVQTiVKfsOmDxxL207y3KXnUP6t0XJRtirdNAF/y/pnfxj6u9LF3QFX
lTW04RgAxRrUx5VF4jWYA7yO8kj7wnCc/61LioNWEP6NTw9sRrCq6YqGzhJzkKNx
R0zFxzs5nY1ypMjENjCDdz8DixNGjvQV3pZvqsKZX1tQPSHYyY6TzWAFEXth+k3r
JUOXWynJaH0fK3Qp02MGL2cvcnGN9F8YrTvh/jDi3YvrsjGKG54rKi839TMu4tTi
k/Vob6K9WEdsGSCNfX6HafwA17SODtaDMNPRBUC3ZVpN9zvhVbdCnTPmls4hicwP
9pripRN5ytS/6ygsJxf561kSZVnKGpCSJUfX+NCMVxsXTshKTSbt3Hi8xt4HFg7K
wE1TGD5GgQyN647KyF2qpyna7i+WiGX8t3SejuiMis3Ks39ifx2qXstqHf/S0bEw
TqVzkX881POJVGgDHeoUA6ut3SxddTThu2X0H62A/VG3UB4JcVf5f8PNnIbfL7vR
wb8gUVvPHFqp3lW383TUjKBAMavXk/DbQmdbrCJX6Y7EA//j56eEh47dQEIltK4x
zX4i4V9jFuL6MrncaZAIiar85xrI4GTFwnYWMCaq9u1NZ1hDME4wQUrHfQdr8hDq
syql5sSzs7Y5CPT48P1+oJSk98NPCUCJyDCjXNxhjJQAhYBb548g2uNIAsYjPlxj
fncQ902sYTMr7NvBm/pweozUcNb3Ynwt9/SapYcrPQ3tOgrpsgie70k1upoaFPyh
L8Yct93hwbTOAQwGx0YxDkwCEGZcyqB1cySPygdEYnEIbd6Bh2uVACHqoJA3zMr8
t+nfe46buiBINzNnt/Kl+8kyUFx7SqKIZn9Xg8D5t3M8MW1gA+qTYohKAcafxD0P
ug+j5CYVyjBca4yC2nKaLfxPsm4rUoRMKWq5tSOrCQH0/qebSOz6HpomyAyB8HGb
kn8NDC3bIJa3xVjp+etQUQmomQ8Uo5dCzKAuo8EPbp4S3rbMzZHnnGolpufZjMrV
N3BkSP5bq/P7c5jOy0ErDF8u0gaNS6qfhnMz71tr037aExxmgjclq0OFNorT2oIA
96yYDsfM1YIRN0ZcyIeOcu1ykwjQdBjcvmeAqmVRpSPrndlpdxzmPyT0aE+3ZC5/
EBceiI9cC5tqmJpLriTe3RmQmmG2yLtIGVF6DHKdB45XNJMM+T5MEpYmMy/ZdOLi
nKrHO1W4p6PiYIpLjeA1vAlGe+5MsNg8nIuMdluLEPtu2OfK/dhEbnb1z1E3h7pd
nqKX9w4w+J3of1pKXCWb/7yT8CLHKrSW35VK1YUdcO2YD8bx8t60Uog4XxDe2J+1
FO4esgwxuaxJofnnXdHeRNBFc+L5wbnSEElnv2T8bM6GKAE3m3LUFhyCi/TWzKHR
RsuLEylwvS8rmJLoxrac8UYb+fA1o4/vAUoADJw4oWz03L/ReEm2+1UkIDaCI8oY
/uklyychdSdQg1uoaMCBEvl6SoNnk2I7fEtMnyQGaJaMcGlozogBxYy/o+ThsNFG
FuwKdFv+f7lAk5bRPNSU/w0G//ghSbAilzlB0vIPqQcYBMhwD1OnpWB/4avPRT4m
EsEsvVaLdDSBdp3+nvx5UEweCv5WfBV+BeUQYIWUHXhH54onV7xCkaxX0nbBe8Cf
tFoXLnFmr1LtJdsZG5j4kTRrDlj/8wH7647FXnI4fyYo+SxtJC/umD3istHxMbsy
+qG0Fd4vZA74AkUYVTM0ZH+gSbAXRaoBa5HKhlmOiwRN6VybamOS4ekw/azxlSQP
Nn93nkQz9gexCM4sEkc5s7x+LYCNLVRidZEhTba3BajgACzypoiTTw5pEq0/pxJn
LqOopq4OA41hMeYkYpSA3bWfKW79wHdr2idV4msJN+uA3QBwK9j43YOgal52O5h+
VajEuCxJ59zmHeIEPm1TNA7dbTUhn53e80uvJGOpOEVDwAqZyBF43sWa/dVmeGq8
cCYuhDDWg/cKS96oUgJloQRwOWpwvwspjKtWwHkqMZTvPQChoZxM2bBpyeowhU4R
OGE83GvS0bDyF2rae0VD1wkU0buTbWoxgdnCmRGDMsWRcLhFg4O15qCwfgsDlidK
Oorvl89gDtK7rnb2lZQeeCj6lWQH3ZKhayhHbvxjnIiJScUC7WCjQNvdLWvNteh5
MZyrYZXzRjGmAFn/6YrOLK3cr/3WWrvKZFBe/GiePmj5sfohQOUXI64Wa2rJHNI2
FdBZI2bqC23Nhyx99E1PhLQsXfmv6AaE3vYSY15sBUWxbxZ7JDuyRe4TyZR5rYJd
2h9JqPC7hzFJ/SzT2gus0kUsTEGbSQG0ieCW9zbEqAxVzTcftR5h9O8jIpj+TWAJ
lnZYrlYX8OjkZd+aukyDV1vQbjy5QHMo+v9qcS/JjE1ao7Q9N2Xg2118nj5MqenO
+DFfY+UmuWotyOyePV3QzM5rINLbrjRh0JXf68VXWqphN8iYbDVxF82ACyCk6f+b
Iy/JuW0wuRoKTu3YoZ5KyCMwUSaAg5zkWXcZdtZ8ZoZbPuwoxku9mdo4WiEDZrOl
HcKTR8pVQn9jYSdZ2N31WjgCl3rt+QFZ7Su4o3JABCFIkmQovjb71rQyDaOSPN4r
ZH05dtRCzzTXcQKRoXW73teJfzEiW3Wuh5pxnvARqEoda2UKZQNujAqVMV2ts28M
AceG0b1oY/VDbrajKnNi4DNUsT7FH5EEIZlVDxKNLGquWnbj6m5OlUsfQEDzyac7
fmwpQ+Y1gtR1JP2YSnJejksajGmdRE9L8C+mtamf/hpjAahOpcJg/zDX1pYLBJSJ
FS32bih01xF/NcHVb0BIwMTTWuL5a62EIaIp5ujJQ4M=
`protect END_PROTECTED
