`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qRmVIvQP3G0fAKd26yK+dQEtKhHk3YByJ+RtRIuIK0aa1HRUIzDFmidlibl/8aNb
9evDXPyTbGpDanR33gwlqdDD0fwmAy5a0CV5ENJvKSf+uoKiWBY7jfaYF3tdNPnl
bu4K9kVG8qxo0JDbOaNc8/w5WGzGBQuMlBw8+TeJTBg542F2rbeH3WdhCYkFNhQN
1GAarxkrJBVT9ymB9xcuQeHfMTrgQxJ4fc5V6ciswY1VYvULQtlrTTh8zpdw6ZIX
+DVojWUzx66BRcKPlsYePZ5m5eUA3g2oRMln2w+1wrugIjgJOmaFyvj2lo7luTPn
i8wf21Ud56hdBHiCgjuqV5pZAnKeuz55mh2YU8s4oPKSgNtYrrq2yM7WvVt4UW7+
At5ZV50ZIwl/iiH7ZDUrZOAiHPXtoUIRufD/CCUDlpFpYdyDCtTe7I4iCjB9iRUG
`protect END_PROTECTED
