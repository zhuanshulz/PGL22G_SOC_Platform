`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6IA9vm+WKmQngtrCFWIHaT5WA7qM0VeIKfPJpnC/J57mZ0JeYqQtrJj1FuGCUMPL
p5pvuPAnRa9akCQxAi1cfeygEBXPNpHNwjXl6c9/QTK/u1iuIE7HNUfGMH5MudMl
E1HWg3wkWvWqgx4m3tBxsBqjf8ShVHQzFTmRtLkGTmqH4Q7pczZxoGg230H8v4bU
dKf4GQfNxFC3Xe4TRWx7Xmz4xvRYhrZDcEEdUoXB2IwimqtLErXRtTPxTyYZosnA
C1B4PE/3gPivpivTThynyhNbhOxgEISN0zuYM0SD5ecvgW5hTFZnP/WhaKnKAh11
mD5er8hSAVcYlkz8W6HAVME3/XNazAcltCkSib1ELscvuGUugdcc9tqho1jA18Ba
VoDryF8EOGD369F7rGsuBg5SskQLauRobopN5mo1Dgpqpab663d+TdqvnrVKNgHu
`protect END_PROTECTED
