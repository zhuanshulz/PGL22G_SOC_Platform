`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MYN8UqlrDWAaMkP72nGVz/DvO1FuaETfI/VmV5aA3W0LvuRLKm+pNx1XUB+ZEP7t
0+WZqOvoDFypf8y2FBAbN8+/7nZ4WPqm66C4fAVP3Qu89Ce1zjIzB+m5lCqiSS7L
GkFeaLaMhVEmbREwOrzNz77YUgEztNgd88d6m4Am6moBooqb6w1r2NNsBGBkFArt
OwL1Iy49be7ysb7SGyeG0QIfo5QHG3Uh5a6Hm+t5sLGtnImOcbSuE0y9wO7gx8Or
/LBa8us8OElvl3wgu7OgwgUsJeo898yy1/1MiS98M6vUQkT5mkhUFUBNMqJHMFId
xIYwr7pbEFisSK2V4Hw4EFhT+JNVSsBjffYttqZ+4uPr7c0U1mTqfCKeHnzVpZis
wlBZeQYHSvRTAlKIG6D495/1EXkVWvCQproR6UWzxTV0XCcsN/aqHkcBaonKKsTW
zEpL/Bu4ftPNTiv41Zk2rOfYHS2zEe5/kRWmveDa6CKsjccV4S37YlR/+Qk7W9Gf
X4SwtE82dhuPF8ctqk558KwCgyw44nRtcGS5r8j6vgANpZDay2nOEyvzYj8LzEYZ
fSPgSlnEW9Auu0N3gVX/0w==
`protect END_PROTECTED
