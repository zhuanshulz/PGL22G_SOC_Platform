`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5VVOdqigCMcbwGXikB15Ep9JWSWVSQptsZf6YJ/JWgUpZjDfj/4K9H610AVlPjgt
lplO5I9xP2nBwwsBS+J868rGxWdL3rtNnvgh+tScSqiJsojNHgVE54UGes1RvVy6
vrFgQDpkmn3cUX0UIB71EY4NLhFoaSqZMS5CI5xcJWABsYjaDQC5wOGCBEoE3V75
VPD0qiEak2RkxuGzkiJ+Pm68kMr0usmvKrwhii0yN4t1f6HeUpvSoJztVGBsGW62
QikrsQyZhwilJMgTy2a52PVn/3l8GVoA3vWpSr3Vq7gFeKzvbvCPapcrBnlkvyKd
W3yWza7wYhtLWADp1XXGuZUJKCj39GuHCo1mKLCtkDjovMR8CUXqp5nclL0EhYI3
NW12l29sOwt0bUcEMgFtPHNK4FZkZ5OD9vMNLUIbjsFuBapdlwimF9G5AXaZYZNn
A4a9AZKKZbWdWn0MwUyV/Tmdoe8MkNAGbKzQW36ZQorQTp2mWZf/UbcJEurA2tEH
X2tpyGMdYcHF1XQ1LI00Ovn4ug2K/xFyWVn6NgEtSZp4qMb64Tws1sm7HtFP6jZC
+ho0lOm9wVb0uOWw7Zy0a8wweXiO6gpJcDby+xsiReR2OAVDq59Yqa0ajoKGaOan
59rbZrVdbQqIaRF4mdhjmdRR1QEENa28tTQvin7ZrLryc6owSUnQlGSopiUR2XFH
xKXe+tWD2fD2Db9rGNGkvIf4sOv2E13ADZTYycLsyCI9wugF5FpKcQSvTuT0UMlo
aI8VtN6+jBbxfN1/7H7th77IKBwZWP+y+2OJR53h2paYPCmo8WcX0AUhWG1wVbbr
fWGHtnkutUM7U4rRz9Xn77kPZD/v+kKAFXb7MTOFeY/I1AKUnwn6KmUAI8TI8mth
wl5XCQLU2u6Z8MR+nM1+494WtwVu4heyquSVPqKFHc+hjTjZWj/4Y1Sazl4j9Mdk
00x3t9UdsxayDMkCZ4xzB+8Pc7Cec/KgSpfEuyiFQx3ivg6W7qVOpEmkGn3sSNz8
jlYkLfMCzuGTUWldDqXrm+SxQUHa4FOSlrC087p+pVDajuTniotFEu4B3dKTyjtQ
KXAU6n9HzIEtuwUlbz5A1kTqb6k56jkMZXGarSUclt0tAHMjHChD3MBxQefDgliz
CzpDIy/DZNtQba+lYHLbEzBQVXOP3mbVNCS4TATqGlKLmehc0ivOoh9C1xhGRNwB
Gh3e6OHr1StTEzoKtW1LLvrC+JZij7FeV2kC/H4pe1+Eat2VW8mXxzkLNt2AmSV+
VYi2fAG69F7/MrmDBie8Txlnn+dXtdewwPaOD8HvQz5Lwx75re7zBrCaBkPyIXJC
QxqyhANOuAbl0MOxnkVM7zSFsNgDqbtQzBuf2pBVt4RrvL3YQWAFctDpmn4o9Ze5
1C/MXUOBYIpcSWsbEfQ9BbBd1r2PnY78xvD16gwBE+bblas39fIIZYYrUGseVa+a
z80TBmoo18fiZcwpY0MHSTxx18JheA24kDcv0kVOVQhd/9khb3Eyh1mGhqr1MRz/
ukp4OKg4j8RidtNsHyhcsT6SSkUopm0b3hr/edMiSDg/+R0AJg7NafaUnjlHxjpi
blrVLStW+Xqkxq9nM8ReacWDUKlP36suejh+XXlEdtzeeBDj26JkrjWFLTpA1t8y
inPt0IReci92RqluIKdRdhpa+8ZFVRs9Swbr+SmsPmqbLqAz3K7uf9bYoLtcZKtA
dC9/RhLIRXg5bUyQMYh8DzeOhMIgZ2++eW+xHUSxmGQi4SmT5hIZNyOF7BUjTgdz
bsmCKFZFJDix646o/x87KNhg9tApFwZ36t1LiMBgJWC9VCl/4S4Hjl8I1wAGsoA3
9geiS1HftvvMdKrlJvZr7ZneWpzIvFW180IERZchNFmcap0pRIuimTY54qIjgBT5
gwvJRLURHZT6pPfXd1EFeWaDoPBsOG/oP9delOLr0xYOUcCMknW0ItFRxNZbyh0U
uCrhN5qkjxxdVc7bdpJ1OueQ2KfVkGr219n8PJGAfRvzHWDkrZCM+gBZ7NKFkBpQ
rqmIHQHfT3zcprVmNVLnDtIi/sJi3Wkh70ZRbFMjr1isgm4O97Ryfj+MCmhPGcHH
DVduogP1BKTH64wFkT1Gmb4Y3wxpuxyE3lKbwoYtjW/aTgHSTiC+a50TL77B9Ysr
Mwf0+UTpttt73/1DcIsxIe2NMUIXHkvjq4npRo5TGXwCapJxAzuxaJ51rtJBN2A1
wT4o0BDfhK4y12dzwbUGpCahXXkKa6GnQV60/TTX/8xMEuI8qt2S3PPrmCMu5D1R
XkYyyC8I4e/8GpkNvvlrz3v3Vm8D0IIXzhFo/zb1ZbmXB2YFM0W+8Vz0D1TOC9AU
Mpk4sRb0pBjcDEbXogjzWWVT87pTr00R8tiUE1TRKvXV8mHv0SbstluCpG3agldK
vVGMsbKuI8OFE60/6ZKY43lQ0YCSrm9xfD+PYEgFJYPS4l4dquMyIkdPZ4fWXHaG
EiRNGIarC1wMcG7P2S29PS10HJMTo3sRhVc+EY6YxGg=
`protect END_PROTECTED
