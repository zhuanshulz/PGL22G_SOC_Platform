`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nVDclvMZWjIs5Ojwf84kB/Q6hB2K8kIHgR+YZ938+c5x3nVha/LeWeWU4bkrpU1p
dPq7rqABWdoEEK826/9Aj/gWlS+z5YBP9XquPIFqJQQZsPqpBU+HrY3rdUBtGJfD
DOoHzkNFzdF2Ec9jDT0mhqRsA3gVsAsp9RjAJ3z2FdmfN3lcTir7H5FuM22ZCkUA
2Lqxj1Ntz/XDLOulHNRmiWPL6UZkQPm5Ex71wbO0ooZBHiIw60tKTSzt1k/9eh1Q
EIj0iWuQXJzxM5Myp5knJB8aG+A4ZhXGauR2YJyPnG2pEUEaMwLPkisZscDQJXWw
fo/m+0KOzhZQA2KGg2et787qEh920Y8VVF5eipTYxLNMi7vi3jC3hLJ2MdfRhVDF
cByprB3kqcV/2x80EwnBSe0F9dCr7wD7wGgOqee2IL5zofHQKminLvmvU8MhHqOM
z63Wvfm3HmNuQ5yjA4MP+paIU+5b38DsZgoXyzTtifHCYltiSXx0Mab+AY+/NxVv
v1xawfMHBAjjtcJMaZg0LOuDS49fYdGQMxXeCPvyss2TCmPk2dGah7qwBfqqrXT2
+gS7Xffc8+2lKhuz2Dq1rZNVwkUVrW9hZtDEUP7/c9xXFb3oa0FDQqv18WDAjE0N
hWAiMYoU3s+CLNk1SImc4Bu/q0XLeMcz2aAD1mTjsA2M9vVxgwkULev1HoIQT+Kb
sPjHA0H1oypwyCcIXLqjBHbzwxMech6MUYdMUkMuV/f4HiWi+jlQ8k6Ss0ycOobI
KQcSw/l2a0tMV6upOVwyYvSSUkXdaH6RmM0vebllQ9mM9NrZNJJTClSVXVTxdXsm
ktfkcTkFVOmvRyq9dWSMXnn4b4jopmMWjGLAvKD5WJ8z+SaTVXSFfQxo2hkRR2S2
xxtxRgFFgs6txj49BNR2UTduKmQOz2tInAYUQMcPlVQTo9eLU/FnuMr01iw+xxmr
V5GNc/Up4AWu6ladP1wIHp6+p/I+PB7h5LOSQuxKD2U0BE2Y3OTrGJB1yDwXdwH3
qpIms/WLQPw1B2dVklEKXlLse5+hupWXTt8d4aNoEtmvt3WCfE6kPxDP2Xz1lm3y
+/wODMW+1mGoSydrmhvjSl3cYxIRE/xMdvS78QxkYPAV1HDhd55IlY94fzyZKbKU
gGGiXxvqERxlJ7VNJPE/fwZ2DG1kSWC65Cq4WJ/ktNIhKTu8UYMzg22GDjZY+tGm
XCwJKaUdv28FfUguHNRqzomsAeNV7r8wRzciuX3wOnsI7/IF/ILKeVd6RM+4shGG
5Iv19hiw9W6V6RNcA78pdBBsi97FaomhpVWSTvA+vjJnrm2H35SQXFhhpf4tRkgP
CQL9nIuiYcKNcll/kT4fCif7tUfv++Kror9oPBDMVaIKqUlmNxsN9jxdBNBgSUfL
XYmLuWhRoQi6CEf5Tqrr7GTMhdSHf9yvbe/wjLQbf4nOkjPHy24AdLnJQHSYV3s8
Y51NVh2tRvYqJkZ4ATdqSLqxcLFymppVqjDF8BUjAPX85BOdrEF6jWmf3ArIrXJP
DuZ0F+O5X3puPzHfyUf/dFoAr03l/6yd87OYmAAciyH+oq6YHebeqsM2yEH7m9bK
Ny/yZrLEvFDZSkajQ0U6crCE5s2XGKDCJ02HK2hzOzaD2aOESBTwxD48dCW33mnJ
Da1cF+jhDAQqnS5hje3mNfkrKE38gQCsZdhhTCLZKdXkdRoDGlGwUqC01H07r5WL
4jfrfAQAa0oIdTwXEAFntDQCECjp3tKIwupJ3XgW1rWw7RrzHkiGhzffMm1dXL6Q
EAFMtn+O/yuEmMTz/Qy2rzBta1xXIe5oVaEwtZQCinXF9g2CHKkvPbtnLwkL/mih
hbvfNB1e/Hrn9CLzd3QRVti3KU6w2YVbDqZXjbX6IOlCJ5c0jgUQ+0wvKKwuEZS3
ypNZBlE/7+4EY8CYVLkwuw==
`protect END_PROTECTED
