`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EefrCbumKEVI6x/hSG63W1Kj8ETN54gTzeFI8TZJILf8au5o01tJ58a8UZkWZIIo
Ja9NZvMeE5Duj5eZY6F8vxEf0bQa/398Y5Ko7h4cb3OHecCxeYMzkRc8vIVsuIWQ
iET+F/MFpSY26C3LzaN60JvZI396jV3Kwc2QxtpVGqaCaud66O4EpQQ9J/s+x8VU
P7WIJMp2V3K0eSdcFgFupDDZXEsIYINJ6IkJjkb1/Slrz3TJCu+YeXpBKRQTCIIr
HwZ0n7WUaNVdLIegZaGlbhg4o2KbSyH8PxIVBpp/aqARuLw1QEkEASjISCmd88Rp
I7qMrP6OcPlCF9b54OH1Rx8Ec3I9214KmCcD7otnfy8dN6OGNroMED68OX4/WAz+
7cEXOOI/kue4TBE89OiK15TiYBf/MDUtj+L9Kl6WXFO9hNoVBSri19n9b6sx//XC
8AtTqaI9gk8k48Pp9sDT6bPOymFaqw6RZAV4g7WffBqiK4pz0cJ7fpqtE+gPL873
itk0r+FDVMYjqa795BGiA8Z+9jOULJi4xA3OCK2BV/3QVEfkR21vE++YWyFAIzMQ
gUGuPloO9vtqrvt6OY8vPWZUAnHb1hSLGA7W/pKZhMq1RmrF+iTt5Ls/jLWH6EFz
IAVmL/GZTUsumLwgYFQN0hsj7AnB1hXsk5YZfrHdt19yl+3LqotQzTf92Uom/dFT
siLgWFZuOnYCetaFgTIH9NrVioclkoTpPzPdA2Ga1wxXIbXFWOQHBjjU/mBQQFkh
5BDT4j13A5fOAyQkCHwDJoYDUacd0xY7KWFH0FYydIDpcVNm7683NrhqgAbwrjA0
v97v6q6tUMpYWzvL4YR5qkFfwhutFPnec+StirydUv5TlcYBovDB1oi03G8xU1s2
mTCj50Prv4aLT+mrakQYO3a9ZVWGupuUmNaLVAEBhIIqermJC2TgTXDW2eSYgK59
OQTrwCjhBumaMKZ0sDyMaJ5yScL2xVPZtsWMbmsrPkIhvEqMpZx8nm/jL1K85/51
9RDgp1CpkhBmb8+gGi4eKQyyHO3otSATSzAX4BCgY5SreW4xVBMieklmu0uqQ7RW
+hESnBjX4d8G4bCzWf+Woqv6kDaNn+gLq5iawV188HGFUi5h2BBxZY/2mJRLHAWo
v12ut/T+uIfqwQQQt0VF54ztNk5Z+qkia6zrMGP4CO+nDbWR/uEvAHydMEQ6Ein7
78w7KQwAXCYv1snMiycLXDsPwnvddjo4tzEmBtUiP8A=
`protect END_PROTECTED
