`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ha914QmNUVhXYerVq6cUKovbdysGfIvyJ9E6Ihi9IHTxP74rNmDoPcZksmpG2hka
V0NUR2xWGEdfRqLu3OTPurswokFLvlcsAJ5UfQPBulR1UB9CjI6rVkYcH9gDqMY4
qKB3b+n9RQTx2m7JD9y1GL2lBxuluGYnElYca3XpX2xLE6wmxXJGfk2FwGlePxZn
6/BUewEDzJL/GENb7aq4EHE8auTc3IlhZ4EIOci43dZtMkgq8byGgO6HodZRAwio
xN82MgUTo3Kuxh2sefp1y0CsMj4V+NE3WiTFqb7+Wh+PLf5hi4hKzSm5Ft08/MnU
GCiYqxlWD8bhv29DFK5lk/kOi/0CmGljOs8V3uokmkfIN9nN8FNdd4LhQ3AW0S+s
/Ycg27o6ax52zY+Z4qHcy1QQp64HqTQSRHFH48x+Tq3KD0zOB+v3EwPOBwrH9XxZ
ooy9zR/f1rHr4Akj5Ng4Ck/DN1HF3I1I+xqPywc0jsMyvSLr8nOf73qGuJFu5dkG
yT6LhRWRfdryG167mmyFYw==
`protect END_PROTECTED
