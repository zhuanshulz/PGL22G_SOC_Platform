`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z/mhvdFUii1FckN7SKO+T9lVxUV1iLGofG9eF9WWZPAJzMgUGbd0eHSpiv+H/Bit
7U0QXmR3rjvPrsdWSt037qnQjDLk6LWIOtd/wtiIPvB2uxcOZNhXwGefY90OM9Nu
73+xWlAfMDgUrs65/nQL+pbwlu7osd/zhoSNISVizNkQX7fNP9SiMJyWCvFVW/19
20jLOYJ1avrF58rgtBA4Psq7R9+nkhaVKWRbG1cwsvoYvrPfeilNwjFVyWNJyxRW
BfImj7rTKMtg7bd/We1amEmgDw8R7j5XZK6evJLwMk4ByOzZEiMKek+PRIs5eh9b
+fBLUzd6eibukJKx2uw/FC7aSeB0+tSJ0kCzhsO+iLm9wio4x8JtCegOiRLggesm
/aCVYeeNX0AW7RvQyCmAmdTE3/RxTlUAzVsf+XxY2EAKIEjLyI/dUMaok07Z8G3H
YkGfAzOpzEuW3SjzGKQmDWijrzus+JX78HFubQikALxBpgZGWW9GJflhoMhHj9xn
ezU/WuYOpbs3ebtX7USCr7MV+KuOIJ4YKtZE8H0xyVsRns0ovOEso6Ikzk/Zh3g9
b2rvBCBsINd9/Q0NDUnt11xp4cqGjPBQWOx12DPaOgmZI9nXOKZm0wnVMnGkzfmX
ZprbRfffMc1thjPkR2p/bw==
`protect END_PROTECTED
