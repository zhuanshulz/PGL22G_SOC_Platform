`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+XB9LjSS8fPoE6TuvWDwLRPcwV8EgoNb/HgbGIW2YUX61YLDYcRcp2sOCax7hBBS
ui7CHPPnQ3QWhdgA2C2M477nIMSHNVwSn8HgAwK5YIF4Mn3HeYqLhlof0Bhy6no+
Upc/2wHIQqvU7gzqDgVlPItCe8ae7T1f8j1qn9zzL98vlhpgOTUve2uxhEJ3XvAN
vJLwQD3gWdoyiTUsq9eYWHukwBGirkz2uydqScswyocmhywDNpO8xlWn+tnc5SNh
OkpMeOj/PilBv/79lEAVvbbDTyPyf9twNKsgpjXGLhdpVTDWJtm/R3e+77FZB2/d
+61Rlc3nPktlr+SpfmwVNIwyIKb88iDDoeC+Rb0mFFTJwbF/jAdU0IIJAiJYT+Hd
NlF8fkTFPtEvGa4mZtyDfO9NMRlKhDinrARWbr8CX9MgNTEB0/1hXX1HNrsoSfTK
x5W0tTlRXWtqGyHMbZanjMMEzKES3GOspNzOxcugHZNZX+bZiQFjHtpfB/1BM/T4
dAbhq9S6oo/kN88Kak8ZOz1r54udLSkTC3utUKIki4dhkZYdMco2d8uHQqeg9gFt
LL8JRewSz+f9OAk/Qzqlv85grogvhWmB1XsenTYO5Qb0BYQsQFd1EaO/UYz4f7dv
lj80Mio+DTnk2DnUcePGTZy4eMkoui6D77f8TV1jMANKx1+oYlbl7b/k1n+76LYc
Gc7JONflrBk6jTNEVAWUXO3lOjDEJSvpgnTL731Qi3BwIgID+i4mM5JIK/xA6rhf
D7W7vHKPbXeDe32hrje8f0Ea3ztYgquqTsljJ7e5KriHmqCiwYyUNfrz/7voi/uT
6i6aKIBuIiBzmkGwSxSxl56AqVcbfOzX46/MdrX885YRLgznhRUinAI4WBnSJjSt
MQy1SCGNSFWJLDg1LRyIrZNGdL3BsBaO9sj+D3q2RtWdkiZyJ7TC35h1TCsw6Kax
Sc3sPnme1nktUHMKKMVSxeVv0CT/uz0+NMQX/J5UYgZjGl/0bmYw5f0eIp8N39Mn
/pflGGfbxiPI4THic2Oo+anB1amt8ULTXVR91CDO94E=
`protect END_PROTECTED
