`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2IHaLC8f7/RdWvC5WmxcQtv/X9WQbIrdLOpJLgkG2I6jecGhsbie45hvRWewVEY4
kTx45w/J0keZj5jUvYbTy+CON+pqXVUXVPPC+EIUuJoYJ/toItBbOBGsU+BDuIpw
lkD8Fs7qGJUCUZsmli4bg30M7TwibPTG8SKCbeaywwHzJZRlFMyQcm5ZTDDy/V8r
rYc9zhAf8WrvzD4R8Xx8eBLJmPUqglLfkbFtxNEE/cVuHR+ecAH5/unC8mSO0ASu
Fu48UVCB4HNfZinzE32c4cUVpNsp7L5vh1/g5vdN7p2s8BBR7byPE5gEvdbk+G3Q
EIYHNe2F4KMc1CPxQ9g33aE3pH7b0elzIVNZhgynVkdsI75GsJJDo21KQlFdaSKp
TD+kAARpnlIIfWhhcfHsPyoteiWEkcTnonOLKHzS7XXuqots27qXfmfXfFGQi4tu
+woQCo3gmnzK1Cr09fIIa0S0qEW1PynIIJyZetdmFOZs6AIfDs7CFF9Yq/t8ijth
5+eczyONLleG4ETxlBpKGbfdDLUS9xhebWH3QsAsmz93S+t2RjrzFMEtgrGzFz/w
dOocL7hYRSCn/2APpRP0Pd0VeVqscUIwtRD7LOCgwYW5fCQiNFMSAh5emrsUeq5m
vlWSYvtjiMXniYwJIGBuJ0w2ic7KPxPna6Yraw4fRzxvOSdCXzBLeqYdJJY45XTR
GYKe1PNt+44LqvcYMMfTLknKGI8b5tvv0Liz3ARmNrj8g7vSrH1B7euG+6vGVMJX
G2oV1Q6FdqeiHnWGiBXzM5PViAEJ2D8AVXAunt9rsLxRDuJLYMWqk91uEg0veWWR
gbYsfo+khrDtxM/qU9mTug4mPmH26Utm4RskV3QrjJK575sO81f9/TKZSX5gvp6B
cW+bn+auc5x+oVUc1wSZo83Tn7DghNViGg1/zJLRLzseATr2DrsYX6sLd5RNrg3o
kjsOL3PYRWGr1ZOeuX+Oc0jCseOY9UqTIXD9IDbDIcIV1wcwEash+ZvaVblNNjwS
gVvRLH3Hvu+vTWpTQLwKVOOPgGOXRo2WvcQ8ZIcivEHxEcHoaCnuwMg5HTQlJTiD
CovpuIQCkQNb4B8faKa41c6aRS5seUu7MQ4VZ4UIM2Udtg52812J85mfzQOLd577
M6fZI0r2vr4PrAeG6nCJiGZbtFUAeXts/FbT8TgzuSrVgKe0hGP7+2764HAYGpWH
f/P9GdS1YmvHdUqfqhEJPw6zQ7yIKqyC6eagDx/lMLkf8ao2lMktSycP46ec/qhu
vg3y4fhAs9Jzm13ueeGB+8QReCXhdHjqg+vZ+xuCmoaN+b8zY2kBelpABVjQuZ6d
BtUGoE5F44/pOTOCbblF3NA8gajs0VMkuwoHtqYpJj8R7LUggXcmYm+9EYtHNksl
xLcc3bCk6KfNmiTwd9+zDQ5kG78T6J6hBu5chY1wLz8cvN/aoHc5eKGvCrMxs27Z
KUb5K7epX+WpdI/62rKqxWU8HD/X5vmf3WRJsqLaqoE6CSwxXUN9h3UrymVuCNnE
gAg4WsPT02GVDHaESWy5e4ph8Fgmk2tU7KT+pP+GCdXlcnJEBOMfOAwf6XWSTeR/
/Kb2jbj6vrtObCb0w+oIjvTbSKcHCpGfFxrAh7Jzz5r1ms+yzdEy9rISc+CLaW0z
/Xuqa/fdwOLfN0tDB0L4w1ewozWUTQ/h9JCUHUdg0WMOU2BpAySs+ybXDNrQMh/Q
vPOXcpzqWvrOp4rfXn8ZFjyBSFOKNQyYIsD/NL99XMYTvhV9sODCMTnvzChgOmeo
JX3BcrmMU21WsNNGO1USJzHogCOc5SiMHMi7/F72KsZj8JyvUZauAZHtiXDTKSwO
FIf8swlBrblxEi93UcTrM9M5spDC22Ox2NUUq74xy4rEBpBMooU/51Oc+v5zIL92
LrArHAe9gvO/X6XjuT1rdX/xpKjBNOY3tI4EoQNAH5kH7Txv1+Iy0a8VBW4IcPq3
AskcltnvnW+04B28MLzE1OLTk8/vR16yfAEQV5xoxdNjwkYveN+pF3P50FOLwDOq
y7+o6V0PZMZTSjnlZybvn5thdH81DEJLHbQvtrnrunrSvUbiYK2fKe2p11TdZhC5
vPj7H2KZNEB7Mboml6amjivgtBX9F0U4ecONMH0Bt1or7Fx2KmtVaSX5CK7jF6/a
3Z9xJCVH6HkP+1BfX3Ds98Biq4PsFW3v7FEV5UyhCWPCTe+3U2zjir201sdxYPzt
D7b0EWUTYzG5sxOGsU6tHQry5r/Xrc9GuXVfuCp3I6WHbCNkm9Bv8gErtxm1zrDq
8cxal6RCkHhuxcDsfJFfcjqKn2TydcqVYVTDNJRjdBLwe2wkt+BUiYAwvMFcrdqg
jrycIAsxO1K8Dh/M0oFhjAtCSNetoBpt6jYVxIBlPJPdw+EoskP91wTR70wScY7s
gmpzIIgfAUCEh+HyT9pWXF349Yk5HTXFusiXT/IlnNK6d8Y85iTnb2g6Ut9bQ8Z7
LINtwX/yeknSWz/bRry5mOvmypcz7p1Ya0NsMQSMqp+9aJGjGdYMGjcGBxzjxUu/
xy0fnBgusYFSMmLfMnoy9wiMK+gfcqJeRxSQj/1ZexXqlFjdnjIdEoVmgTrEsShX
rnMuSkWCAtvteGoUIAzgDe6Ntyl8JhgXt+hDkYEqMUbB2VB6SydbFpn3MVHw0iop
ZvGlS32vEhtaMwbnsy391yfeu8SnMrWF35xX0h++ex4IwX4PcxHsP1DP7xy27Owt
jk+bX0xy3NZS0vY4lLabJMSeYHKjt77RKz4sSUW5hht+cZredgNKrBe5FzWMWirp
F3x2ngeW9Oi8AptoiiAcfjcbJZAlHgg+9/sQLoWEjbrpwJGPxZaZTSVbCXYAxiHD
gxJPdo1whHvAed5VBZxlYht+gCQ9XSY7ZeeDcZQFM1ha7nwe2G1o17NIbimdi0Xp
Pc/QL2ZIhvj5sj9Z07Eh0slf56fFSMAMsiWOXjis/YoOjeh/UWLeGZ/HNDe+2xnQ
5o6AARx7r889c3jHBeSoeQaw/KgQwB58Tixv1AvKotr0BYEB9ucaZodbU+GFu8xU
gkKRCfG1ASlsFiFRo874ceoKS20iB+cGPKeENINCYl6RCvQ1CeDfnkADtnweKaNQ
j78roCNDy3hhqsVzbe7VM2q0fogkWI380OZW7BOOaSE3K0PmCrJc1xo60txjROjn
SfgjrvYRcCFq3D3uUZ6BS2S1iPDtHPEGeuySLP8eD5oSzJSHPBMYSq4rem6Mr6LM
ZFg0xU7u+RDkiJPzlYtbGUVdrd/+Ki5WYBmG8fUEs+BkX/AwwyMwnw8KZqWhxFsS
T3XcCPYBKSVLhed0Va1eJfUn12DCJUF3/i+gGbmtpWI7aOrc0WU6Co2pfX/cHXSy
woCXJRJA1vIr5Knfwg0g2DPtF5agTSLb+r0UbIqJMKjULcvxStqgDcEnySM/1P5T
moDqVlAa/18bkUOQCLkNs/GK7Um/VvOiXajOQ2buuFQMpOjKGhlgyxRkeY15ZQNV
sNmSQXED6P7qzHzVwVh6zooD99faHTa38wzHLgV9fCkl0paYO8r8pv31beQ8t+in
6fcN+4+aw2E/6hteJEUhP4QMXE1W7lnoqq587ArjW6IaACsnnZSksrNNiD2rDFcx
fEqj8BF1MzoEiaHm/pHD1VOehRNwMHXLBan3e2YHv9jdSqMfamhZ5EQJKThpPRg6
WuDldIwvOl1uly5cqim9OF8rmee7pu7wFypkUA2ebPt6hM6j77b+0NPW1V96mtAf
GZ2v2ic4y5CkTDQLUuX2JZAmzbI/AkHm2VKz0qEl3wwTGFc3JavY/JVe5ubyZZXt
oDk3fsdfRdaf0msfTfSx9dTYjKAJBCiuzE5wt59zVF+NW62cZCRmwihWLYZUepbB
esXjRcHfXDYQUIiZqRVmTInhCpt4bi7zIs9uMd3jh6yoO952j0AMWrPZk/oyfzqH
4kGOmdYo43/204TOcu2rULUIRPI0kIoxsWFM7dGuxjfe03GBcg2miWTZOESotY8m
wWzqM36suHfNj486+AsORKJLm7HBMr3AQFJ2PkAX/4ThF15AfRGwkm+VL6HImGKg
i3YC5XISQS5s/wVZa2nag+GpHRjQNTzPo5lf2yvJPb7A7mxytuXx3hZ43wXaMlei
O0SNkLCYktsHFpbUdZiEom0C5ZOvuzVhUIDoZ893Y9gCbc/kUebqch2QL5o1j4fh
mTX8EKdbo9scdgSZs0zZHxcofqZXaoHYqvnMV3g8IcGKN1s56El+/oxYwV4VZnxD
euZcKCryDysWy0MqzX+GwaIKkzKHQrEMD1DhR0CEoAjE70DIlgLtUB8xAdTZQChD
PiPIFq/ipsBeNvineML9p+Bta3MTaIUkChMIBe8xpYCYc8545uoc9J8pzj+wMK/+
vwfxq0RNT/16nt/5wCc8GpKwRQfpv3Cx1cm0QL/09XJiNOBVdN10sjp/ZMxYqKwN
KFNNgECvVA1jCIt720hhxpE8SYw00NVVag4sm4adAP2AQyweTEPa1zrgqQjLNBsX
fLT5zBdoxwgHi5Cnt/r3sA==
`protect END_PROTECTED
