`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NOwS6BMNJQgSFcY2hZ6o6miPnv2gOsvM/eUKsgx5n5I38JKvFmpQRkEjVaD0lFw3
aPLYYFBV/8Df4Azr7F2pGWFmKGwWDnyyP4Xu/Pzv5AaS5lRtxheaa7OkmtppgK/w
KPyJyhAzqtI3tm0eUrtqcPtn9l1GYA0wFV0rv5A52bLk0dQ6gArFYwTN58Cn1EAZ
Gj3q33d3tAWEmabVG77N1pZFSyBY67SLjB68MKiZZgly+s/czbNQplfD/lL9BgUm
VUnWNab2zu4+5nI+S/Mwfflnb8zahKzzo2opCkGKM8Or+2I+QsGrNfKKfnXz3e13
NCk7VccQcZ1mHGsV4yNw4dM/TGHhvD9IX+LxUi8vMS1DK05CGqutSDO2tkTYmkPT
itGfIR37ayO1XhXlUdsaSrZ9VRUIJ+/CA/mWEllK+FskZuBHmXwEJncSuL/B8g+/
jV6JidnnzZ2svjaiR6QR3jNrfooNHzSVcz/mCWowlxGNOvdLHBWw9xBM/cSmab+v
faibUoR16uERoPx9kldSl52ju4XGesaFxNhEhHx4idEcBfoNxRcDvNGaOuCN5sCI
sV030w76cGmXqo3k4xnr75OW5xfEgd0hSNNlcZpjVIeI1JrcFh5IwlOPgvfdogty
5K6Fnk33hTLsJ/JIko2DI4rnS2jPmOl0fL8F42vLGN8mXgjN2gpJ9asX1LB28YUm
+GisQoBTlM06XCSMhlyAhl3WYUPV0qNbvOfrohkyHvCx2hybGH/R2W0Y8h456c5o
`protect END_PROTECTED
