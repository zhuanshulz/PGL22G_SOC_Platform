`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OcmtS7dLm3BPNrUobh/ufBgZ+haLkWmWm993WlEfSxs00kakw1MUXDDT3XBNzqlD
QLB8RZifzIE8daCY5VIDTrTrgAuAdLCxk4Rm6M7tQ5l2AwWDFHY97p+Qe8rxdpDA
wcPfZJIN0HdZsaZTdh4RzqmmS0A3uZr7PBVng7x67vLgmQFAntcNK4zMlk7oYCYQ
hswxgL7JvHyXlYsm0+X4+hIp5n5ymiF69DxS5HMn4enMgOON9J8cHWAqWtfop5PP
6af3/Th3BNuD1wdXNjbhesHgpbXHt0IWCiu9aGL51QvZVPXewloACdXhZ9f7835l
5UV+6fA4hrKenmwAJe+Mc5Oz/iwBMnbCUXte6a7y3A1+v/G1lu8P/Tz/pNklvgfF
DNdyDp5F6RxBIv69AdR9+cZgBPi9lkqhAan1QeSPW1yEIH4sXkp1Dq5f5xQsh6y2
VSnS67NZGufGWpPpKXq2eCfX9e5a0ZpcKrIMkjK7ukSI0S3NiekQRP2tdecUIn4F
nEItFEtvNk+Z4GuNE81oxnMfyMT1PJr3sZHFQ2gYqtckBcgx/PW6YWMLH/vHxQ9N
Rinq6pdROVU3/WgnxIbhJw==
`protect END_PROTECTED
