`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QzFjLbWK2cuJ5/MP1MufPoKTRYD27j/2eiX0F7DJCJcfrl8bzB7wQMRFSD4Nv3Ut
2aLQ6/lHyrgM34/Y5+2yESprCisgxbgtHtboGzcDJ/InZHyzeQLgWyKxpYCg3pix
1Ej14XLzo1UshNCvZuj+/MGYMsZkWvdqwTSEixy/zk+htLQZdx227+HW+7HjhBxm
wDTpHWE2c0HrwAGnnDlj92LkG0lPCxgljpKmFjDHNKa1cHACk+dDIh77IgWADAPX
f47+2/oQW3KyX1jLsOo24Sex0eLEs3GNOY+ROK5/XYO40HmEG9wxdEm/eW3zv94j
gIbaOfWkDmUjbhD8bIdG3jVtYGXvw9/17G1mZhOPi36yieijBhTGaIpU9xkvXX3J
R6Ta75B7fbz2xCnSEUjT4AcqumN0XATe++MPzzq+/xTx4+cvIe3bbsXFG9NmF2mC
fDWpuQFgdyWFgrPuuyQ68lHuCWpglNu4xdg3QttdmWHb9UZWBBePHHgy5hkTxJQC
sxUTAAe3KlysvASetPf7Seg9llNbyACWxOYL1o0VM6r+pofptCFKO4uRMw/PnnP9
Yv/UgfEdPQr5KdlHUyC6utQYTfkWib8tOfDD7+E0agBRhdm3H+nCd5x4GkyrARdP
ES3zdRSwP+NIonpltoT6p0kS6dT/oDatYBubESqhKiext4JrnWQsWeGkug+CW+hf
bBQ1f88tamkoHLhfxU219ZjOSvYbxal3EbyiLznNY50=
`protect END_PROTECTED
