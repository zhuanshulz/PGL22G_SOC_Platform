`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5S9ukHdhyKNTnGLi8DMuIZ4NPl4ob0kSQdC89KYOuXGuWf5ta9JnKPQbSlu4TOXL
ZetnmuL/+6gnN+x5MEAeOfTKRKN8OQqpvENh0wN1xHt0CQ0o79sCCHaKWIr5rbEK
yZr6hxA/BG/8O6DvAFyPxCEPPT9EmJDwda1fuvThidS4BhFyzx1M+VzMk/eB7our
ogUdV28+iEDplmjWPWKVk1FdRaUu4neIWW9Ejz3GWU5fhWa+XUwi0jauArtiSSB2
nUuIZeSh4bP44huyxDwtpGbQPFLJJD2gMhOYsvqWMeWxpyXZHRF9vMJOi2+GhcPn
C6BnyhrnAtWUQTbKhuNaS/f4K09mGfxlkoAfN+JQrxLLNdnQZe0qPtcXF+yTsLWy
Vj5LPgXP2oLy6+8zwiYt+IEeo04NrhTo2zNCHZaOW6u0klIL2fc44u++12zndTz3
lVi9ziXLCMe4dB7ebPO0d5mVvUejoDGWNzdb27PfZD9QPqm/tMZoLPhepWafeJga
vEK9q0tn0rsceqwzymQqp7uoDrFB0KhKqjmHBo/2njhCSkDnaQQI376Y5HEskAJ1
luXWcMb+8IEN02Bv80NI4A8JA0OtPmwQZLYoi34DYSa7VtFxYm2XihANEBAMQNKZ
NcceuacF+aOVEoyIRvVl+5othRws9Wh/Aq9dqukk2FP5tSuA2wQ2tC2hz96XpFhI
NRMocxEFtbiJRJHxDFH8ZujEXaZNlS2OrTehl5JETqJp683UzYPh/91AEkvLOcml
bx1Gl5I581kbXmUbat/RLJIplcETdl6LhhhT97IQiO1+84lRl4QxYGTHf6xTm4xI
OU8ITofhynF8WNeuuFJhkY1tj6FkVFvbOlM1I1Jgg/jrdzqPYNmet4v9os3EXDup
NTIaSQDNXFFU3pKXMR3fXDxXGlpmf5lD48AwTCF95Ow0U1qCKXMCl/6/rBKMjq/k
NzwCCEtqHEnRP8mVzPzSK8XzwAaBdjHEsRNThMJ56ZchHE0LRueDZcNb3ZOZJLEl
E1a6UZQKN0UqZ8laDxqGZz2DJs3OGFMiAshvHUUqMimirnq/SmpMrE/mvWzMYIxL
2VbB+c5Uk6V8pRIBwIkvieudEeqkGZy8Xz/lyxQj6Rn5G6RF/rNMM7LTN+H1T8HP
IFELtDkCPx6Y22iXjhFsz/MAsvfrgzjtXteTLoWQQfU=
`protect END_PROTECTED
