`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H5An4ynPluqXju0YTpH1XKfNTtkgOphQnHCAPjHpia/g1aE3kfdL/HcTzA6UlYn7
pxq1+cAafhczXfwtrjQ6SpYftvJMvPMCdkUR5Svvff3AFbgtOJ0p7gQKLJTLGt42
nKXZ/GJO2ShxBQOxTsjL/sPIRPX70chcoPLimHIS695Bnc59WMDYW4wOJHh2xF5T
ealPjm8CrPyD7hcfSF9sby1R9e5G5t/bG4aOEKX4LR4sRy+pm1G7IlctFnae+qlk
Wdo7IZRo6gEPOhtyORalgkgHfhdLT2J+YC8IGseNLNkDue+1qmkc5HigBJRuQQvq
vNWp+THmwOc2Q3JQiYTSF3ETq9vVCx4XFSkzw0ge1yNgLOyzNlrjU5tgl8F0ycUK
LhvGCAOuq3tgcAcDHd8nUC+fbWhNLS7z6j4o18lzLTUy3I6W+but5AqRm3JxwBYa
63+MjoIpXbMNSRcdnY5gY58ynrxb0uOcdwqdCIft0eBA+PrzMz9WqAgm9K0/UsMd
FtuCcwuIDWoy/RUHVy5DmQ5LVnPn6jf9WTrtaU6BEabzV6SBrvX8KhFjjVADcPU7
pjQWa723vRn7sDncbzKhJId3Px2QqdyVPCdRSgR73oBB6/YHXEg7RSCvo2PXxcwg
Vx95100VPL4XOBLntkLr/PTzBzxy4FMGKgnJ/kQcBu0djOdIn6M8xn9FLqxtstBr
rj7HiafzuSf84VY8B+x/TI6RW+QB0g7t2F4UELngdWvbCNfCVcrzhnvHxI2ES1wr
M8B3DyVOaGee8rrVTKK3hcMlyJwiXB4Sw9Iz3MCVA4SMLptiBjw/6PBeoEZBFL1P
AIDolbkEMQO5hF8lakrfZh+Hd7GIbTvGpX3WiXkZd6910cWwXR4IS1k3cFLm4LcU
5+l7QXDaoGBK+PZXcC6jm6+KYeLc3pbcx9lbOmuO2XuBJN4a8Hs+PD4RXMs79zyb
Ve+C/vSWafalkSfJJSSia8wtYUzA+WAwhb5FEQYHZ0EsmyrGSI7R1RywTlW8zXEY
yXRvLYjF3XbBqGK6Q8obWNn0gCk048v6byCtTzMK636heJtkY7aew8Uqvcx+A6+q
If4nbgEus4qhsE8hlmzVyPE65QSMB84STuHAt1tzJesC6D2q9z2jaz1lX5v32FkL
ObMUSEXuhyyTyFglyETFc1yYjWmJE9UomdCBRlzF7QChUrnbqZz7OAzV9jqbalDe
g0YkbqGeQwXzA/VvkBB+xj0DoPG9yq9ECghoTW26ngI=
`protect END_PROTECTED
