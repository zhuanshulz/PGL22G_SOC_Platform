`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WUiXnQ7hwtGsRvE74rw4iaRPa+ui6yPinoFDGWx5uHhNBY7AKl7VF3qyYb9qKjMH
O0cDOAHMOS4oDtHqZHsmhUSuV4fxuuHV4hmINx8d/kXbJgPxwMp7UOSReuWYOy5s
/Ue3XJSSto+nnb50yPfmbP5Oher0xUto48lXE/eOj0AAC02MU0T6AsCCHDTEq1iG
K9fmyB+AyNQ0F+trP8ha3fHjuK8jxI5vs1oZe3WxNck/Z9gVP+/j6h7nYWkWrCrb
UPW9zbU1EBfSMJ5iYnfkXx2d6mmEgxUtyJ6CWeVUTNLb8qzoE/C+dXt62qCo7TOz
8ACEc5mbbKqN7zUJrc7jkQ==
`protect END_PROTECTED
