`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hfevE7nCzxugPiuHhClZR2dQ7Hfx66QUNd7eKQzFwHfp4fpu7A+cH5LnfIHIAPlo
pX/011F+joKdpZn8+5esezfrdVR07UqxZQFg400gQu/G6yhiNzLWfUfT3jWnEJdG
0U2U0ruxQFvlnF0z8ZsSWqXaEYaX+CKBeUo6bwaQMEiQSsHkZsLGHXBNs/fu+nXB
Lspb5z/ST9vT0tiQfvvbKwCiFR7spC9CjaXEjBMKWLHOFskzhHVUugEbWU8zPD0o
WEHa8PwBFVf49OhjgcMcnQK1NftLMa6BGAzfKjXvY5Zgh7+QlODQZvOwTrVfbBZZ
fwLuL+RzmRixGyYFnAEZBUAwnlft7sFX6JefOkrd73lFeKUbRSYFMOs86nUuL/7p
/jJD8pa3elxGI5gPhGPi1J+iuyV9mR2dcMNLGw4Q6fjbWr4edP06CGq2ApfDX1ZQ
hlZscZiTgkNbwvqo55Nj9ZMxZII0N5K35cJDTNEnF0Px3wddCUzrtPvsojeBFgu0
Ta27QLm3yPdHHl6eY7RISHWHCJRnh0Ri7O8Gapmuw7oiLDFgtMVK5SbRsTQ3dCqJ
ks0/idnm2a/ukemWBjfxL3V760KhWQTtJxlFcJWetLJw+bE1sJsK11/NFxtZPuIm
cpoHb+A6DXX8qbpGtFxLtqRutMpyt1XmhiA+SubF5BVGES8JZOwvIDK/e/wR3e9u
KlAi4giPn4+jUvjCFK55J1knD9wX0zAhOhdbTSBsVRqGpnVspieg8l8UmEP7hjxe
6BFS6DLwgaAbfgNrg4mSqjfvGvJ26wHT8rSREHyiBjr/PAk2eURUxrUiiju5penA
Ld+sTm/MxwIuKLF5rAjZOacD/tc7u2yoIyLMW6zVnShzefDVZ9MAFVqbamUMtiJP
6NX2tIpXzAMpIJXig/ZUCg==
`protect END_PROTECTED
