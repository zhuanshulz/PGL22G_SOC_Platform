`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h5qCMRx7SeDzNIyDDPYE3etii3NnkZpJU5zFCAtyrtK2KemqATyU1cPxL0CF57DV
a8QF+k8YQ3V8qQTSQdBZ+3AAulygsSK/9nShl7lImvgxX4ZSrsZPy9j6rn7XQdO2
yJhPBzW0E8Go99qX8OcSo82QS/2yPu3Ad2hryIHDnx+bBuX2iWQKKO/jikvTCbZt
hCv06SbHzUEmxk1RLx4zjSHm3lmG01v7XaFUfil0tKtKDPruvuTvepATSuvhwWtk
TR1h1HpnuwC+vDZF3qvbyevSjdJoQBEPL48JC28v7c7TuE3pVOOwm4Eqjg8k2Yk9
Tcf9YcWKvxHbgva0ufPps77NpLRoC8tzRvbo9Vnbr6ySfU9j324rC1K1BpwfqN0I
49FIEfihfn1vfCaXPHGR8doiNQ33UgoMrW6shx7YFm+RaqeqciG1J1EMQ5t5Hfk7
/ZSgf3RBFGXrH6WL6EP1sat7eJGFR43gE8mUSim5g7oyP7HBn5JUeyFQPtJAd9TM
1X6sQEw9EWVHQjp4QAELUXv7dQ6R6sLS5LWekeld794Gwz0/sIOrQPYcZ9zIbrhI
evphzjm1UM6nMwpd05zd67mq25bmdIxZlnl0acd3cKlkt86HjIGfylfoYRdUt/Sp
C3hC/xMOdrDPclMTZJHyUaUAUoos5UEf32LngMpFetTax124JSOiqhzI2Ronx9vV
ZgQxUYmQu1/LGuWYprSTH+ZVgZcRkLY+wLG4o4sagMQe/rLGULb+OIBtbhuqycEM
WOvw/qnUlTNVcc6tz8pA4J9Flv4qif1qy7blmy2Hwg3cgwrEIQHURXL0xMnrnbYQ
2ABREXMFDvPSwS8YpCqSxMA1F+AWIi2NBiZgchefjbUg+ZkVR9gip1byhT+e7WmQ
WwNzy71F2zu5JVtnk5+tGUlUtOIPhXv1ScO6xFkHvOakrCaAzTKsDdFrRMNYs8YB
oFO4PY4+7yC3XqP7C1dbLbfUjAnu6fYrqmc0mf9nrOovneEA1kM7ddJzp3u+SWeD
b7n/ICwvEzKI76OyYbqWQy3xuq4VoRVXhyxdpWhwcw8qoeAX3VCcg6bJL7SSVH1b
7Wa+Qxh9lPPHJf+OemE6xMe1T/IUT5FX+yLW4oXPfrZQvvJO4Utwf09lX3MIVt70
Odza4e1y9Kmx9EBvVZoG6E31ezN651vqn/2L8sGKsAh1g7fdGYHgwc28mfGlQIh4
TpkDlIZ4/NpNK5gOvNDCM3HUAN44isba/omFdoqRVDcrZNGjn4z48nYw8xbXT30A
b6d/wHhubla5AffrhWqaXMJDnG4cAmrHtTAeAS3vQWMbjIxj+HZmt2fhOS4F8SoQ
Pcqdg3WozG/F2DJ3OMPpvYh6yFMPbyCUKrpLRXXjfyF3SjSYNmgmm7d/B9CRjbTy
h+lGcK/AMac1hnrniGngVQpDNbhGC8rjWy9wcFoL3vryiVhaYYQh4G+duWIdcQYT
reOusMELjviu/tY4TY3YDC0q3KUcOx4tIlS3r/BN7vVDp6aW/5OKSrMw/Jpv+xJh
bG70yc4DQ73xRhA2UHhyHeRZIrxTmmkHEIwLoSPx7aVhl4gwuu6AFVxN72xOBlo/
QyNobvnIPd9HbdBgENKXTjb1hN8Zo4aMl+kv9urVGeWYW6+1gDDV2sxt+D5xwALv
aIU+myPxtmVMjX6pe6VLeWnyYdPF5lCXGumyJGXvJto979YEaD48lluw7WkKazuH
FODZ/wZ1eDvSNR6ggsaOecIN+XRQdG/kU6vPQE6P06H92LVPggByRw1bKuLlVBed
7kW001KuRELb20x8Nv9IPbLhfBsMvu2BQRYEgeyHjFYys8AzwoCoEaKaAW2vqU+s
emuVkYIUK3EFiY+aWOVkhLML/X0ZmrUZxY2VoNdFqW/JB6+Bwcw69MDEGcr7nGmW
ZGe1JpS4T/hLRKKFYpKEedugirDAuggYe5qG32qQJKXSp4W5Pax8hZrsoMavegQ6
zScPBXlKAb9taQQTiZ695N93Tnnio1b3qE5ZVgeeMh4kE2a7IUrn3bovpfdQYPsG
44bNCWQ2O+PQy8GTyaKONRVVHxYsgVs9wZvnLZrZP7nRbFODKAl0PRm9R1ncNOss
AQzUVmQDEwZwOQctPK9RW3Sxr+INkT3KnyxsoPCJAO+G+/oW8cNVyLCIQ6y3Fua9
oypplPMyR9hWTk3dF9un8d7tIl+4di3viczzff4QwNM+HhLacr5d6k5unHDHCtvW
aUERmUFDuXhEmVHksA4YXkIf85aG/PqniSDjNnkC0TDt1bCJbsDf4nCrKmkRrTWS
AsELsNr6qwi2wjYzVuq6fI42wAv0HlJQzw62DnZd9dAhVoVK/vMYvJQEc5MDToIO
Xf7S8MTAlLApxxbRR4bHOo43uwtduUYZkzQRivE2unx4D8FmLJG+Mrwqx4C7sOyd
MR1DB8Ejwmwo7GjFF5F7LqiflEoh7P8ZdK59YjcvZfcb9CBhK79AZhavmEXSthfY
5lYeWGaCPwadkdcupBSXQ1HdQYqyGtIOdWwxD3coZy1EUwF9vdxTfgtLm4GBE9tc
k2DvWUTPvQC7ML0a6PseN2W8DACh98Oy492mH4mz4ZJJSeXz1whaSXwq9QVTKDDb
j6Ymr+95scmTwHs3+JxMuAmF87+Pjo6syKO+LoLLliYuwjaSHh6z/9LQVphNE6W5
4cWLtOBsj0aTOqCNJeyK7sENt9KJaPC4cr7+ZMCpYGpYNFp66kvu4lajnGGsnpEw
vG5ZoXIzo+/5UnouK+RBIOAmxDd51DPupL7OeDRLPUVN/itbiTq0eXVXBwCd2jV8
Y3tLSvCbmuR6XA84ED3ci56U68qDrkDzfV+8ISqtewFtZ5YHI6hvddG0/ToNvuUZ
3cT63lzfD6g5l0Dp+WvckTmsgZJlR5JLLsGY42SPa6vXaNqu9LrfQsstaMhXPYQ1
WjMPz0VMURPvdujgUzMxtKC0R75iP1VEtZfq7435fO8+Zk54rGm7/49vGzOts5AH
1pYQ+jEYEPZU95liM6Xv0U71IqYo5onz5B1sYTIRYP/ehApGypS+1gBgsJXpEBvu
KXA9y1Pxo8AG6RTd9gXUdS17BzQKgbbmPEMgSQj5AywUfjCXkwrAkPDiV7qgfhFU
ayryKKYHGEOPY9c9twnumqXXIjPxKW5D0a3ofN9uSyot4YQekN7orf8rhRXqPTMX
/gKHwKiWgg6mM0GInVCuo3B2u1dpx3b+pB9667WoiJ8f/5Q0mlmtdglZ7/Zh70jt
JDVDFHHBRDB1A6iij6oXMPIIZjsYvW+DEKVComg6fIl2TnCLQeAen6cl/uFKxf2x
O3xGk5sZxr9MPuN0SziFPkTObwl+541jqihyYtjlkRaFfb6Xm6Qgao9a8YrIOE4f
m8SX3D1+kN26qkIwS+PS9SsYVvzQePrT19e3IGRiz9+bbhX/VcyhS4f3ITIyz066
MQkrW+97dBhJpuOOfPH/dKBJxEapAIqlSIGvfdy30DzHFV14asBFmbij2I6ZWcBx
ODNpDd//laH+a7sz7+5jHxCr7kBJATWbHodIev5O87JwjnfoPzLqnnkpGdaM5g2p
DzMOxaD+0L6IkbeOwwgIJXyeGvHoxFY7qGbFwm6e5nW2IYYQ+YIEaSMRwt7+O8wv
J9mDw0mO374TcYs9DHObenKQTPcUiVKQJzIxKwK+/P7e4ydP6JwtIKuj79v0Rlsv
/+jqGw9h+6vwGeg/toVlAiz8B1htDJE1AbL7LDXGp97LQ1fTeuOQuuLbLT6R0DGX
AnwPQMdg9Snq0KtoJ1fyBGGNO6jr359SLB+lVfXqS7DqJJK5rayVL1+q1I5aGWVm
+D4Go5BcU/c7l1XY9Nubq2txqw0reuMgIpoXA4ydyq37ZjLwdRAJLSmNLd4Tm2tU
VNIMPax0mEagfj1pwyn6AYA3ZF5/1YLmu3w82IS2hbv1yjWYYNunR7M8qwm2QYBz
TCI9yK1ko2J+vTNww8t5kQJmpnn9JhKcnTxHneqqJDTklGysKRcQpVGH27voQOfF
xpedbDoKs2JGbNzFV6oARekH3F4qbQ+pWAtzpXNEPGlZEbVy6IrX3wQBuAbgiKs5
5CmgUJ3BiJ6X+IMfgc46rYZLjKHjIOW2NMv16Lwrz5bWLIbGWoxDI0EWtf11s4Hx
q5cPiIYHMp4NyjTA3n0mAKXE2xfeseVnNZam+PRBHgRjDk2AkxA7wKPKyQyI1YC4
zVqt21YyP2qXo27oyatIEhBx5FuAjG6prsXnJIfSgZ+bwbcKDw5QAXHcN8vdZ6XT
cJFnGotwCWI4kDzih45Uv3Ys2DxdLpbUaH5FK2Ud1rIp7KBu4bVtTfPPLBgsj8jw
W8RH5KXwUHCNfTRilSNEMp1f6fmcLGrm7P2TE5OR8GObNj3TjzObM/qaRgcG3Gcj
RH8QDy36mYukE0G2DGaYfQHHlFbKrfMkCdAQ2VgrTDEJ6mijQn1vQmRPR0yk2yeR
6YobdgeS0/z5Ty4CXIF3ri9kb7fF/lSX/Vr/OuIc5KLImhOwM5Iu5gFErkkDIOfC
h+jrHilFITV9iff7U9vhbRYB58WxDHprILFdIR4Fw3AEiQl8GFs4vQcz8ENu9DiZ
PHiqCZ36VSeZ/T14+BXNGplrNYyeYDAVjpwLyz51a3f9pqlxDBnLgycTEllie6ms
PJMy8bPkP1KnLbyxt8R6Gxt8o+j9poFmOOu9mDDsmW2rImHCvZGru16v4JByogCf
Z6uR77t5hXNiO71w/6gTNUCoCBBjdey4P2OzexjR9/ZZjrxn/DzFqmiW4oqQahRB
0/KyXzHG5jmFdIG4h7wJANY6Ic0+xjEYAv6QYjY3zBd0YB+b6qtJtT+m6H8JLFOC
jMpjYsY6vYJVeKMv/oAexUfeiJnZfyZBvsSnIbWC5fDvzrVjt7S39vSMEvdlz+g0
awD14zncXiLeFi3z705H/0H7RCRIAJ9WcPz7Z4mSu3vsemsoXQzcnsFavfRYASR3
bI5y5QaUya70bNTvNDSjKP1M0NQRoKBA+pu39eQ+UxnTyQieBtkU3HYVibtn/jaI
keX4O5I+vtyQcrIzZ73niy/IBhqN7JDiKeWVowq+q/lY+BssBT4Rha/6dJI9HRWQ
4UHE7B14Ri8XK8aNl470r+cxNnaG3TusuqDVy+quTa2/NVpLSNr2o3ouD5rqdVO7
4EzaxUv4ApE76Ofvj7y7MigQ3izpw+++jVin+JFQeuDQmF73Euj8460Zev3tXQYV
t/X69M/SOvJ1+47EK4/qauIyBhqywM3G/hsS0sll4z+cHfh+xxgdMaWni4yan3Jh
NjzAiIs8gq3+rG6HCVobk6lFK4bIhjVnpVpk1zjm/IlmhUa2Ytb08q7npwvVaT9z
fm/YzfeJuoUBCaLszGCskCRrbiT/esT6OaDoWDH8KpdWJLDgWux6OELH9lkPCanP
xprwVaUPJhZXK26FUGV/nz28g0nfpisJv66N2aSUKCxz5KGVHpUGsEKasR31oYba
jo3f4asNWKlKDOP90mYdZWLbgBmweKU8eNEJiyX7iEvhhR3Y1W5HfD5agdKUlabf
AvYYICx860wSSKIUD85tIDpTBz2XhelOydY6KlCg0LQCZsKEyD/an1xrolBS3xLk
0DAd6ZiSiU/qOBw0jO3oyby5h38v+3YJJam9+AihCnrLeItDcn9U/ItByv+Wj9mx
Vr88lyHmBHq7Ccg0GmrDnzzCzdmbbD2su1xGvQBwi23g0a+6JwNnBjvoN3oxkTIM
e7//O2cDrBc2m1YOk+hAN0ia0Fdw0rqhJJO96pRlrRUmiLVKi8Rz+cTAr0znKYII
UZWCY7AC2U1u7liY+8ZnYglEK89eMT5D0kq7eQrH21VquoWzxQ3y0d0h3Nz6IIPI
rvXyQ/fclpf7lqGE8fMlyJSoraApmw3uct0Ty1n5MEDcdrk+0i4oIxHnQ2MwISvG
NfWo60D5rkk4O1cNtzqugVcUOBMov7ppW9+MCm3sfOScJBPwyWJsWK3fEU2i1gtp
xIa5M3mKE/lzBv48Zw5PO3WyvQ9PDkeRnp58w2KQe0WNXZjDsGKTYaXu1Uttgs0E
dEFUKEmuz4RkIdQA4ODWblj+RxeYQtZVneCPxSagQEG70fOzP1Lyv+JVxNnAzGkT
zPcpTtNjbRgs0HBy2mIEkB6qXI0VmYYH1Av35Kprv6lyJ8NoDAUuFYM7TkCtXYJW
1Tnpm0PP3kIdP63Gk4u9V0wC/bTdZhFveEsmKWJqTQBuhXmTd97fG/+u0S1DmbKO
0y15hlqx6E16PqmZzl0YxPI9tsRIbTF9gIX5lerIXrT+aoEPCK+hRhd/YZPdac3C
toxLdYt/ah5SzmvhD+hm5XM2DXE2FubCz8bR6PUDEc4fth33xcBeZgyg/SWjfgwL
xIzdPdBE7wvUvyzQzMl8dntdXaQm70zoQa5hw7jE4euNe9xNxn7elPC3IN3bmTC5
mIMXex06yg/hjiOtegiVSiHGaHkRpq3HmuhB+VtC7bEY5jGrrRyVCvyv+i9L66Ng
E7Q1T/f6pQ6aZauoYLEFx/hd0u2Y9YINvMZ2lMoF5OCJh0bpaHAK+MvIHmPuJlHX
8Q758Chk6v2KRlvLPvT0DqvTyRUiL/gzkY8JjrLN+CyGpxl9Zu8mRfo4b8DwzfnP
u5TWpLFz5OaQ94Ok0e3sJtWrnWIMm6womr9/Tjs8xvAlDaCgZMWwioUTtD55N3s2
qFA48anUqS1ZGCX5WvRirJt8M6xyNPJ9eCZDCyMUhklAId8q09pb6W7uEd75IEKx
K6RkyE1dXkyrgbaaN8GGBUkcF97BrMMeDUK6a/Lh7F7aF7Nu4KDp7j5Zg+oeZI9v
wl0O9JwgWFgw8fCgu2++Yyoh6w13E2S/elPXYXjH7fBysZFKH7zADG6Rw0AeMOmC
SEP4JcE/3w6MLp65pHF5a9YW37n14X1MfdXbjl+3ouDaYZY2ITSMS1G9dfHhhW/h
CzHKtk0gwZwR3nKQlc6AVxcAq472JowFV8GQVfeQMBqA054eq50afExmXIdfAgTS
Q0L5KiEwCp31YMlyowQ5ZLdLovY8SCKblZ8BDL+zTpLAzTbRtTVn9I9i/to9Y1wf
4dWb60rodZPIqq7uNZMjM8u4kkanAk3nZUpwIyVgaLX8DFFg5HS3afQBG6c/O+SN
aSxo3SwOJR3Po95KQksH7CBizjcs0d1xHmFSY7liQMp//CEnxmZmkdmhZECH1cYs
YOKGwzP3e3FWPSt5R4rEh15WrGigmw7xOtntwow4UJi8oljw2o+/6s5KiLfBNZ5I
CCOisv4ivsIJJ9LByxHL3DWN8sT8GJdsrkXVxnxBqkpa1kH2MKxfl/GAzxdSarYY
DzHuFoSIGfnKz0hUB604cir09bwLwh9yDfcur/VqaxvQRm80+2jTLKmEz1G73SPF
RF2euLghot0MI+Ql1rIn87Nk0ZL/WCiPQdEspuFLK5We+hwJ0EoIDhi0jM9WFiiy
lbEckPcAcF3Mmqgk4monbrDbVa8aMS83TQHjP837QkLCDMtc5pP2MHcGj2WLfpIz
sK0wvF91tLlBaGEUg3xODl7Fv0E69pnYTN6x9NracKN7PRG/hEBNv4lI543DZLSz
KxnE+javg22I7ga8Hu2wwLUszS6I4MUpQtkwmcf0VrTKJRWnv2KyR7KDMgWXiUKu
wkfrF/vEN1iq+GIwg8hfhNB/X2nVDc18ymDm7JfLALCj3Ntg4c5On0epEgdyhgXU
zO+lEsOJdQlOlpYblNfVqfnoJIZ+ckwRhTZLX1U+zPv1ZoLFhfKfi7+wmVWujy0C
G52+ZTvgcLd0LasdwDOQ0M6n3znC4866960+7qLVJ8BDS1DvN3U47kUBYU4qPhJm
uVx9Unm36rhOx6yBgQUH83XYdDJT+h6Gbyg9wNyLwAqCt9CQkgn7HmiZXKJKNQGE
oUAq9/Z8MggEHFa5pGdyziZHCHxPdAut1heKOZofAwuSYfIVgXeQKodlUpOZ90u3
1649gUtK70rQwIrZSXEBZjVEdE4xun5ddn0rMx6CZZZHb7M++SQgB9GUTWVX/JCd
IhrxROUZXwyxF4kzmZT0RnDEH61LqTLnnCPOgvfVkp3AjLkKYwNLv3SlRHUtOc/f
UHfd9BrOKMkhQ9w5VW+v5JKsCyafKNATo3855PJCKe4hfPhZsTjjVP2aKUBeOeql
XOcJHE1Ixf/tUz8ZwYxtNlkCrks0lpik5FkuC0xDziFDQnazD0yu3dcR+6IzzxM3
gFeIuHi/coEH29fds+gf5kZSjCMpHeufZmSOBpAZ7wcBbKyOUgktmfV0vEUN02LR
hsnHo1TBy9gB6GUcnzgaU47yfZ2xQcoOYfbdjaz6KM0=
`protect END_PROTECTED
