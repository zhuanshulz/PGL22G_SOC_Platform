`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HXzsoIU34c4WLheeRvsLaIgc4HtEfknOKtZjYLzF82M1CiJKgKqvXNC6jbQMKqHE
z4JlrtEpywg4bsPqn37YIp761+1efTaZEX3rQ5rZAQaY0FVu7fwYkbvEfYt06zqu
dKCweFgRGuJV3bEVNq0Rlo+FvA0GhFvIG2esI4RvIEDRSDVNEtUogDq/S9/ETv/h
Qqq4OaTQpAdxaI2zO77bipGeIFY+PdWO13fQQ4Zyx0+x4DcXSwftbtF9VG9GF9Gf
GVE1wNiOJrFcy8VchfJiSBIwXRPWVYaQhT7gKwFJjFbgbXQ9rkUEAMnwYFB0qLz4
aF2fanEn6IsMYsJuvOMbZtVP3Vp66ih0a+dnvzO0MWPUtiiduE8grS0DOirhryfN
YUBw8zCpI3mJwmEk6MPhgoYWH7QnpImftcrNd6M2u30KLDzS7WtIxGwe6mjiPv+a
PqlouR1YzsEFa6wSecSXin/kfggcTEgjksL5h9pDtjKdKfXCHsq39mFM43QcP24a
jfutkVwd8GPmLUSHWhjdopd5ePu0ok8hE9UQML7VqnjzNpMAZ82ELYXtzsBChOVi
`protect END_PROTECTED
