`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A4OlOZU7qdgTjdVkl+NDvgxj5MKBIarleqOrvgvNT5VymblayjYFRR09ziHL2P2p
W+Py3/CQtop5zCvAR5BCu96xVjMf5NukJF5MyNCxfC2yiaHpCuRxW83R3d+qoGwD
tQCcoNhygmmowsrea5gKoVcV12Y9NfObpN7Crho7WWxIODdtNfthPkVuswxe16dr
tt3ixjPGcI4zv9Dxj53Rgdl8RTQEyc9ARE9yFsA5UieuodVbCMh1Zv1EHEAAZi2x
mN8IZp2mRXQ347z0tsQNe7tf5SfbqplhRPf1V5T3Chrjz6cnP1TEBt6iwQte+X3T
202SRIaMkEDFvhiNQp9HOch3KFnTEwTmTllY7aKj9yOk+jGXqHsyCuevvJ8NROI9
0+XMQgcaPrcCHfHmVF04mRE+fl/Yf7x54N2MZxVGjWeIi3srqajd8KbLbU5s6p63
JXwTlSVDuo5cDbCtSWB1CuNJj/rX3eJqF5UL36BT73VFz9RjxNWu71OJ13Ok0oxQ
Z++76OiRsJb2GPT0bBDPeXyJ5I+2/LgY+xgAJNvxnfB8ywuYjd6Em9mjPbHT7fwy
xgDFCaigBo4rYBUjoy646Q==
`protect END_PROTECTED
