`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hKNag+TySEwSkfxni4YlafDmike+uDD2F3kDEJdyeDGsCsQtgjaYhtK7n/Bpr3I/
gsL4TkF1p36PpObEhAvuHMEgeqFSqxGOkkOOTRqipFwOw+1yabP00zU9qUVJuL2P
pig4YU88E3DSb8HRSSAuq/Kjm/NoxV1h10wuJecjGASxGmZG8TXRD0ro7yNQsZOO
2H6jqJxH/TX0nEswZpe/oRO6IiiLfjhIMrMZnY3fx+YaT9SvJugQ61ilhC6nnGic
++a+vMb4Wtf3hCGStyC7gM/S7U0dXCtFYGf2R7le2SVYvkG+qQ75CF1idTDRwnK0
f1usCUVzjFqxUdJ5+27l4KFcblTLLVb3ZbPkaK3YHezbsVQao2Qlu4cyUAHGjdTE
zcqbhIXz8yaXaSkJg7zzJoTVt13f7o+uxJOv8ZKqS+gb3IoTMypgSJthuekaa0Nr
s6FRySHaaaZtoqnfZUt7RQBV+3TyOdiywK5N8/kT4Iq4KMH/N9ccQCYP5lcn4rlj
rUmj1POpwabDLsJkMZiS0LLC5hl7T3RMSwTxBRcFQ5KrVpqee9GJL1jH41AcXtOc
KeK7oWeIcV5+rlZWo/q+KIiWfmR0mwrAOwp2MsxQl5n07qm/yM/jJihQWcRGVAzp
`protect END_PROTECTED
