`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PperPNUFzAPh5NocxF8OF2MEOjc4I7JlQFA7aqKmzshNkrT28xtFmWZUIXpdz21A
hZ3TTUnVY9d0s/qullHJUztES1Z527uC/S6Mt14Cvs9uzlVoEjtgST58Pdnf4uwj
zcbP/XNyfXlCZU3aEnQKZXRG9EnS7s8DDEWdQ38KbF2o0ZdhFeJBGyLC+NMdSQDu
/HsmEfmjUgOJlo2jK6RVFD2RiJqYwb6f59yxPcoW5Gf9v4h0l5ptZlMaQindUSLa
rG6uUXvF5GvlxGvLVAMT0t71GpPsigrmrSZPAh2chpjQNDchUzfxbz75oQE+sEtX
H09JSwm38WfenF12S8N5yZsmi5VaLhc1xKEm6dOcpdMiv9mSuEm8zhdc3poj7Stv
TI+N+1HucQa0uv2StcNwJh3+VYURVqk5Xlg7ukw9PDq8JSA6vwkvlNR/jl9fZywf
oXZZlBQmM9KC1LacIrt/+cB3af5w81SK9WfwWGgfpUlQxuEijskSGzyEaQdr4EAu
v83xxLyRd8rnNvkuOOLFaJZ82ug8YAvyv1zYWOVDAMbta1goJOT66Dvk50ndxjCt
GB5BXVo6SUtz1y8alTpFWDPVc/NHEaKBRS+N3+kZOxwhBw16Lr0CK6Du1Fm+3hVm
EIe/UHULkWzgmUXB8gknRsUMqsyo8dO6+EDRu9/Yhzp7SL6BVhXULq8hobqm5hJM
9DR/ClkUtQuKvB085rmx03J75Jv9wJZDhcjWlPsQ5cR49/9X1bmkS/z8ls5olrt5
9wncFvccfneSfzxR5Twz0uHqkAZAL/QVKx8b4Hm3QMceVagQfnC5v8OkXDLohgYq
Up68oJyk8RPa5BzTaBGzL2ZmNhDjiajb90eKq4kYFzHCFjXd2/h+8lPgI00NgU/M
Y9n3fbM2zVS+iWc1pOY4ICgXWTyoPwUq+FOMWgVp9OBhcBZYaYGEY2m9PeJMY9xb
b0EfLJSCyJL/O+mbqnN9ATDQxzDbaeNRuhvAgrmEZB/VJvS1srOFExZJHFNTyDik
qNdYMoikUewKS1UFpZ9N1djy8HegWnsMm5eZGTOZFZpeX9TXWvmy9g8AjB+HABAw
ytXDIwjHm3ys3PtU+YLP9gGfJYYYTlFPLmVtb01zi33IasKrOSBoV2LmNMSPlqZl
3cE9tO7sUMClYQggtitWWvz5E8pyfIeiK41DIUOyww8emnpJN22RqSIswTENNlcZ
wt7m0MmTFli4AmgAcF0aFCWSTDSXeXAJbmm7oYqFQ9M5E+pswXpInoQun0CiKuWa
hYwODGVfv3YmhnZ65KCgADkNQ9D8aqml2Xcg5KqHOvOskcIGFLMDV4Yw1EdGnYYh
/w5BFE002SXB/ENS2QP0sus/5hoYRoe7vNMutmytVJ/iUyOtBtQ9VJ+m6gUDlJpQ
VITfTRpQuaM+AL1cOMY0lK+vZgbN5RX9bOES2ahYGnyqF+22MF6P9YTx1mMcnQyK
jvSqu2fYcnAJ9l3mC0xuKNYkW51lNU25zst2QCTXKCwF1ZA+9UP67vHgBf/5VHtT
kCB1ECJc1GcYj3xwpEZHNMMA2+BMyDEDMTvO7FT3qACj3KobHrs56is3ayWXcHQF
2WdW3Sz1MbzoGGk+IoLQvBFInNYmLBf889eMluaguaYKjVQtdOcP2QuXxUPK12I2
v2al2ynK/fQdM3iD3D5E2CuJO6vNPN0E6wr6SINgdyvJEwVEjh2fQsBXb41dCaja
5o54LyCQYlgs0jtF1gp7g4ZeixTvRVyj+tXh1JCPgJZuoAkRgdPL62HyJuJElYhL
X7lnV1uK+jheGXfdAkwXKmFcwcaF/i9NoMkDOHMFd+5hBfPaNoRQFc64tR1P0suY
/YLOGKqMUrEQeixdlAcazPd9TI9wiP3WMrimis677PNePZBL5KfGhZ3qdFK2wakC
9ZSbMJKPw64yKmWi9okIqvCXkVCTQZr8G5epIWZv+TgrX093aGIkpu7Cu39ntYKw
0C2U676Uo0e8MhFhLi1n4gWSvVcHhbPHJ8LeGP0Hce0uR3+wbae3paL9pl8MMnnB
APiYffliXRelKdB95i2A/wyz8Pfl1TOVKQZT7tQhnxXkTJPGKfLjmFVZlAkyxBx5
2c8SoQuoI4DvwOaoGXwZuQ6MY8g7EFtrFcUF9kvWoQUxQC9ji4+VOu/4iPY5OriS
/lkCAoBkff2cMcLxxdN3+mIE8qqZLYk0J0Rb4INyM9dz0lwGOpJUkS+PhYFSuzhL
/9LhJDpHYmSGDrnzKUvZ15kklPIpy1tmseLCibMZmmo=
`protect END_PROTECTED
