`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3x/mrWQ4CNIsN7NAamxuOQoylzqbXHn4VvHKmtXqe4HyurKyFor2KKmJeuJxSHOh
wdzv62D+25IZocfqbrRBbbJvB9VCXIxe+ND3nuKg0zXt1s7s5i1ggrG4Lj+Oqqqz
9GHK2HGIlTHbqL46A9xtXlAQzh6fpVRyWCg6jNMe+n1ddZXXDvoqiyUVF9forp4P
RpF7fqQpGDDOoFhkfZ25+NNtYAPPN00weFvXE+7HXg3BD+kHj3m5rAQq0mwuZ+YK
a696bRpgbWPvpgFQ8wQUHE0zLwNEFrTnT8nqwyOsX+vDrBpLsmzi8kEzlja+i8jm
YFMN8sVl2bJmAyJUpMuyP9Cu+NC2yryBNkjZ7vGuYGvHJN3ZpAFWqZkSt6IFM82c
EpnVxfhbquQOTpzdOOchra0oUoNlcOoXpYElJegjf5ozef0rsijOtDZIafCNQZqn
NO/wgc7hwVO2+Q4nwCjCtPj9F2L28U6h2AYHpmQeps9LGiy2hzCCD6pS9fyy36Uw
uPP6GNeBY6GHjZrVGenkq9NPaf1W5waYqW6YzKH7OP4mUzAps/BaX9Fx358poOTd
`protect END_PROTECTED
