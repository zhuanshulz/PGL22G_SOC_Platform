`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ru4eMZI6Qm7MnQRhSMEFoIyRY5o6a/YS9TH+ngHyec1cS0mEVshaXPZnYlcXHsBP
gNKM70eckVnNdAmjysN0xXeZaOYNUfPynHw+bqmBNdXeYcISrIcdT9BMrk1FhBK4
iqcR4sVR46us+ppFGtXR+13M2ixbDljY/sHocDG+CWJ8Ez8Y1mc8ba+d2Dw+WpmT
MJ0uWWOtEmzsHRDgCXgksKktKNaDWvoKT3DjWg0ro97b5yNEIy/yWOSdm3cZiURX
7usG6pFQIjVz7Y/27BKZStlnomVYrGsTcXBGZ83fgdqPVSd9FpdvdumFzRF8lZKq
IDueuAkDSSHYFy3mXFCwHs5J3n37SeEB5ElidBUsrDeYgfdz0xlO+r1V+CNNuruV
0uiZrmElnxPBQciMkxcGWCvw2KUZRdQW09olOTueUbd3R+dw6ZQOvfIcGaAF01eL
mTVR6YggUDRwjnlqaoIK0wbqWn+V7zxVvO4Q6egNPGuxcu5f1Oolr7BWTQbx6rBn
gV2LeG2z2CyyDieP++abMJaR/EnCLvi6hIqbdNkTuZGLwiUgW9fQNGGIiivCgqcV
3scgtvwJ+/oOU6JJfYa1n7VEZz3ZAYxuM5P0bimTldTP5LIULndXGk6Vo2Km6h8F
yulj/Dq3f7LA4OOni0eoTsQ6ZU9WWKUdg/NbNpGkw1SaWrdwv6yENtHrl5oCIBpm
iOPIJavlmuXpV+1zN7r4GPHVXlCfrllN+bFy3nDdBxUgoMTpCjdT7fOo3MeVrSBr
PxW1N/S1y50RysrdQVh1wLI7+Bnh7H+duJgvtXDqn6Dp6WQyFM7TqG3yN39rEBkZ
MAxFjo8AEPpPFS3oxMsSaEt6CQC1gG7t1bEv/39Flo6JF4yWOgiiaRbP4uSGrehR
ma4ntPmsFdEN3pdkkbA1y4uzgSKQOoijVfXt/ldkZckhTTqwmt84ZPKX2KGY5mFY
3gh6fgj422IOOQyYu942UZ6jkwgkUIes2LOAor1GcmSJmZfJIILAvoMHDRauner8
HjLhMEtIACzOLQWUNxY6kIZCl3OtDIYLmpEyWdq6+qrxkedNz1IrvV35Jxf5OQud
h+sHj29MLhOHpw2NJxYyXiYfb/IGBZ4xA9yZkAQe03nafGgo2wSnjgo27ZZn4xcB
/PuNThsvnfYEqRgUbUxX+/SD/X4/TxXb28QPnkGr5mE7U41m1AM0jMn4yde2AZF6
a9gZZYTL+bUzaqngZ7mAST71515V8Mc9b+B3CEKpzdAELfwe7n+t14hDqtscSrI9
hY+b+5IjBgGkmqXbX03kTlGKUIW+SBaKs9wdnXTEVYTgVippTqMQZrrE/ibuCITO
pz4UhCpNhQG+UB7pM5NGT7PnQRpUYUErP5B+G7hS9HwSt/LDyum6L7BTPI3P5Suc
NrXmE2vF7xt0v9XowwXj0riIg0u7vQ5pQuHKrtM+Aw4ZDe5BGP1ypmt4fq1CT5jr
k3vpfQ1TLX615iaOwfgutQIPngxKL87n1JAiqiwhZJRbtXDh57jwkB4y/dZfrQzJ
RoN+xJYIZ3cP1vL6bSAU/cMZIUs5PAdvCyika1GRq3iA12oCVNC58FxL5LAJuytY
/PkXrABYBHq17QG1xq1gQg==
`protect END_PROTECTED
