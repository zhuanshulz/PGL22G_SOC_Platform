`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dhA/J+JY2D+UvrmDMC7A6i4eGb9gGRwN7L9jzzcqYUXiNKNeowa6CwGEMSQxhYTw
JoLy8s/JLLQn52x6UAdq7Yh3xwEYLrEwaiWKu+joSPuuJoJgBp6rH7P6rdC5PS8L
XakEL5ua1D7JSA8F7JAxlBfqRqwozRG7CulR9xFD+Uld9rXz1mVvriHGX9RSr4fY
+4DNYYklDzNsJ6lxBfVEIFUnQcfwTDg3T28uxW7hQzB30Wdrft+CZSTsUsSlqczT
KSWhNE5zi3RrzHJo0vB1ElQpePv4cpsPt1bC2TA1D3Q8vE/pa4XJrfOmeZfIiL4V
RQpv8MuObVH6E/uHHYMS8KzG9dtalDQQBMhqZGZW7O0amNIBfoef+UEdeMVGNrY6
sDEKdzYu3xppVzigvOFIHFFQwT5P6iIUjWNOW8iTQTqA+KFEujp9nClsEje90XwY
33hdWJDeINbCzE5QY/xLpnQc9zCEnuu6TU6pgHt/paDDg85H50v/Z6akFdOE700j
wD3TFkmSvPyFaRP/dNpO1MaqIVL5yXvG2I5QpJWmZ+8LwGYGDRA+3Roz2jBCLcvn
m2KzbujzFyjljLQL1hnZgTQuG/Q9eR4/0kjCpaEtl9glcJ+JWv4ntVz3Q8/JYR0A
S0z8AlU8oAJSp3c9QUDs/t6hKx6dBHlhDr5si0Uo9NO08zxHvDFGvxhBIsAes2Vy
UfWyU3eU7qfmB9s9TjTN7etZllaMXXoVSePf28sRffXh754oP4+OE0bS0C84QqAC
BE8f0WTp8ryI/XQC34Prg3OY8x7mM4r0cbIAZCx89WNVUYPAR9bE/s25Arw6hbsZ
xTXa7C4fs/CAqUdNJMpix5HgJ3iVqKbdRZ0eFI8uKyt+d1oGUhIqPQSHn0LyHYOC
LDS6Cj7XIuy0hH3YxrNgQLJyVhUj5q6ZQeVjBt/y8kGRo7UbTXy4kiLVQBmAOLF7
bYGH35coaakNgU2RSpWOCp7DAvIcHs2JUyEiys++i+PNIkSR0Lb/v3ha6zL1bYIu
+XlgDBZx9GgMr0itGcCrSHxdgba2aNGyLpIPPP3rXEuGr8Qd+Dh8nf7q/V6eUbOR
3Xa2RkxN15c0pt3jqQRthvoIL2GpHguy8ZeUJnzLD9lGdbF0Owl4FQV3vlYfzWHQ
ltcuLRW58ZAo1bkHJx3/jwDQ0A1s/IKm9HNqn4tn/2WkVdkXXOglmqMuziFBefAE
OpIQ9Js+2eEwIAbT6Kj6vOLnIqAK/i8GvxUK67y9h5YQNh+9P+w7GtEMDp/ScQ0+
YdjBUwmFc44K6iCXmH8J9Df4+K+PK8qXYvHrMH36zaZVb/FgKnRcl30obnNFLKox
TjQKEm1cyd5CNcas0mm75f1IhZ4aZlW2CEVpteHqMpKY5/SbV+JvdcEihFPd6faB
`protect END_PROTECTED
