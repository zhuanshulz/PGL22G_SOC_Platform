`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XfCoo5gUwRm7ioqqGO9akonm9+emQc1u4S4LZ83aTXclgHzp0N2HAiWqnXUnm5U8
htGjKc/Xg/J8y3RGBCAkT9i3213iTdws7UJdcWHZib0dSjFBpgTkOUFmGnwyb1CV
mX6SgD+UzqUeXJ2gGXnEd6ey+ucXokH1JFmF66tWYYhGpmokNji2/Qn2V1hjX8E7
qkl4kYlrPhcO3+2/dMzHA2Hp+uRZPuYu8Yf7MaHd/HZ6qQ5BDdypbwcsusZgaLTB
f1H+ZGSgQ/f1ttd/abnqVe1IPf/N3ficSSDoL8c+Vy+sew5sTx/5R2uXlp67nimy
aAbhPxvSx1oq6azNfK4DLL6KQurt4zvVCfUFE7xUxGi4UuxeLV/ucfY+dRUCo4uE
cc1WstKM4dO6Td1LV0UnojvpOwAn1iZhvcWKTa757oREAUFjLQpHSF8l/6ffJX59
qRLDxFQdDFtvT1bXRsdkmg0JmWvkCSn05XRswD9J71jJs++3Ue6uEeGHbvsLpVKa
u/OoCVnJUHykAn7lmizgXlQVsRueGbMBkitMtMVbLJZ1o5eA6iA0my8CZYRbDQzh
S8159JD61C0CNu89tpCm59rrWVE5HVN8cAS+7+IqYFQqtHWP7C415JYC5tzC7lyN
IzZOdgAAic0h97OhrXivTXeCzphPIBm3eIaahPQvzBsm4B7nrKP7j0d++K8pYgw/
a1caVymIJe/SjHNjcdPfzI4olMyjbztPqlFJM6es5B8BlVI3kd9islOVKiIWTd6t
Y4MSX1tYVZAww0L9cBz4wXl7JhBUg5WKi8LEebj9H2DPbP3pVmCYSxKZtuFzYHxg
oun2p2FQrS/uuhFoXADLj58EP2CxlKhsqRHHb5LiDrFpzlSWH8OcwaAMgoK2I2yH
VfiLP/U27ClS5I0wkZPE6FQ402B7pcCBVBP1EJVqWqO9cW1IaRFuw30EhvxIihnx
LYlLsimUrGI+sCcVQ4PvJhptGNDDppZ/WAxzzshqtuwegqN+eKNK/0PlhB7TM829
VGkHZxGsfBIZR4ryojybcl1Jz5fJ9Uv61HvV0SKZcPTmLpeeIEaspb6jKpZtN4ys
9dsVBdf6q6m6oF/zq0Qm1QWvKz6aJH6DTQGxLdCZiGgR60U9ZMQmt28efS4gT5P2
LLaVUd7xS8Fwpx/wVm6pUpILAcTq0Ss6WaBDjJNFv79Q04GNwXGgRmJdID8OVJMs
1npynHbWc1qaXycj6fhnXaXOjDNTFtfjneYyOA7+c//FtrEgT0rH+YXFS5t5O7dN
13eZsvPmJ3JRXOnx5+97PxYAouwLn2kDBNSwZMNeZFxvGi420PVkpoiK6wS7SVqM
3QoSNpzVG6GkI3PJIzptZMQZA1LX/FNbzv1sqGa2zW1BmvNSMD+MBzJKAYgJ6kGg
sRbrMtZnuvFzzIn6y+ilDDED1oAWdDGZKjjAgTwW4kyoU4rd8LVgrksHSBcT7Z5D
QZ3z5YZ0S9E2ncK82ouWpl84KcuOV3tSE33Xcf2FRC0+MHFNrTsnCHEzGFc0oHpR
ni1C4yynIEQEPZEfcv87JtodDGCdCGEhSsYvjSs6bpj+4qf3QZ3pvI4EMpO8mVcZ
/3XEG2/4ut5Shn3QCmUq0kuNlAAXmioLiDQ2IwAmMKcQTt4nmqjzOTFhOhUSVbQ/
9W4bfe2pYZlIpStdUyP+KwcflqrNWdNnVnJyMAvwFlbDFPGbXUX3lFEt5oxOBXpQ
SNn+ZtiG9OD4j+KY18OugeJmEl0mPOVMVB5xI1SaktdAzON6V9OCcWMUTWXLAs0K
CBWuvLlUgj25JMz1m2RdQqfeybwtilcBqG/Qj3R2EUEgRweEkjjZAxSnjAIwKM5R
jqwqba+T3tKOqZ49RXbB8OsmEytzlpc+ufa+3cTvbbXVolmI+v9dMFpvOddYHv9y
tIYpyH24PCXNXmYThI3zKu+fK9HxTWNFMCZKcqKQcBbXJJsZrhelkRcpoVXI8dWA
JvLtYjftc+4aZuuXJgUjtK90qHl5QjVCN36ZMaDV0Xh9/KOwr5IGulAYSe72eEHg
OTlkiXxv/8O71QnsTUM2HXIaml5vdjU6vOFnYI7tfu1wIXVm6Wdl+oL6cIzUWDdf
U9vPrs8mGhMDLsKkJ34X+yncZTkJXVVPP7JwOrGhHTxuBkadtvl9Dk/ykTyC7hgD
YGJpAFEgz7y1eUq5iNQwZOQhEjWOyYa7DW57M55bIS53pFDUpGMHedzXVuDY8/gE
xv8obefnvYwJo19w0L2n0E+2t5RYrhjoprV01O/6LpIhlod1RRf4xzxQkA2G+9uV
PD2nku51b0oEqI2dIBre7Yrgn86s+yjuGq0FEOOjRAxjAhW8Kj0yQ+9QhCIPG/5w
a0xggn0CvTwrZMXKGWUYN/bKoHjk1Da8Xni4Q39upmRF06zsCTSJurDv7VtkRkWt
JrZ/TgxGWBYFy7JD+LUhNyxIo5DSZ/wfiz/Lhw9LQK16xsJwQyDUr/HuHRPprOMO
4usCBz5g6ze6OTKzMUPJI/kqyW/5vW6eeyqXyv9SdDKevKLVyOPM7wKJNKXalWxH
KvlhgaYefDkykpwejDGJeQcznxwMZbSoyYn1GrpQE1kFqWo/7AluGdjbnxjgQaBy
4JnJuIH5FI9qU8j45UJXSR1Vg21cIsXsaIyji4iYAqP3z4eREs7i2r5SvROCdol6
QZsm97ZWGSv/KeTCsksBl6MSDIOeFG/VqtPi4ycJC0V+YpT7Wx+JCnmzoTK+9mgT
jaDPOij9sdLcyazE5LRfl/xQmA9krjnzzf1R065wG6a2Px4DIx0hxDNXei1VJN5p
pjFUjMUlXOeLHBN95AwRJh2i9S7SrXJKdvaw8PKLd6pLvReeBdC5GdT/iQjxeIFz
JevrEJZcAU8aOUTdAN2nZp/sF1d7miTHIdkrT+KIgGGilJEk6NzGLDNJofHmR+8w
vEiaqwDXKcny8oGZXeAt9XL4r7JVcxniLs7JZ2n1liKPaVQK+dbyWUnEW3jp0q6e
AWK2A90fQSj6uHpYaSV5//tlzwFzDXD7MBnmeJ5GiCu4kPrjyiaXrC9P2BPnd6qY
OOZWyw4JiMPzLVDh/MfmDrT0ckzCNUzs5ZE37plW3NCia4AChXrANkAevjvVdFNv
rgg6vIP0GupZyC48q3Pu0Al/XGMlnmfw+BGsUfpImcPVM/d6htTFOyDU+7roID36
NEWLDEOn8R+3CVgxO2e7ZI6OwWgyjd6cCI02YUL5LXievNIPgTxfy9xB9kpM6Giv
RAwUv0nM52B/KUopZXyYtWjeZ9DLmMep7qMFF+h6sByoNAgFC71HD/0x5e2dpIF5
goNznO774NzuMY0W2St1s3LP+hJJD91tFbc53fG+9D/wXOy9iOLZ7VJ2bUv6rrtQ
5YBEqKSZXeGbJD0cViBO0321uSvq8yKgGJKwnuXWW5E/7tWuFP7gDtGnphm2Nfi6
EEpArDfKnx9/VhaUPAzaqiTUXtGIxtqn1gd/w1U/LVgmBKuWZoMLYeQYhRTuTISV
a/NaTNHRPldDlYN6zmAwRZaD6ZMKjamKWpvMNYh3Puwo1QqP7H9KvXEyFarNzXFk
StfMo0OFnFCqBqDaiqWqWNNd4eiFkX4nSkZWYQaiD9/6lIZwJpUUysZwUk6/zAor
pbusE1kR3O3k2gK/8aouFDjGWUgxbIXywniFTykyI6cfVgJjCm+XzgQPe9xVw8P3
dziIdaMJiKW7r/9AoqSSY+yH1s+ERrA1ReLmwWk8k9uSFbvSiUIdFY429FMUYnBc
RiENqt407P3NJcNFHVBlAW4U35wVg+BjwSq51qLMVtiMivfk11z84VgzGkiEIFjc
6v7eea140wPj4WnpNfkJQvR64TWsFYpz/ITCFUgUp5KdkxwxmTNsIhZrjiU+Huw8
/iMDSMcER+gv29SiUKwZdbTKGGM2AR0BgxDWWnDCBFPC5UYxiTGxE6mBcOUS2NVc
gBKTzUB2rxpD5P14Az61zxoJYU6coZCS2eG5BzoEwsyv+wKXcQLqYguo/n/BYyV+
dc1qd/b/xT1bGIZC7AJQYFvMnE/VJU2unmt4jhO069j1wm/YadvQ/1453ZL3TmJx
J8xcbM80pZCVPDB7hsfyULIsTUNKGfoiKgYAO6WDuz8jcyVKbkf7WJu/Gdf/UOl5
FUqrvGhqvuPrWzFE815dQpmZSycHq51mO5QBqGrAAmPL1XF4Rph724r/doLsfj6x
BN+HWvslD1QKRXVJwKq33To7wTWN3UNnFZOPE55QjkK3W503Bl5Wx0we6eGH6X/J
eLv82ZQLhdbmq1TtJPk4OWyp1hhppAKZTha892r5e8PT8yIfz8xFDQbcqXBE+P8R
0iiTKjNdoG8pK8gbta7uvnL2Yp/+USoFucWPBe47NGPwZlhCn8asRbdrBCFzkQ7m
kjeIloAMgZ6u10BVSFokixNGwI9u3M2WomGRe07Ly/c5t3r8Vs0qvdjTL/So+dmF
TquXaFf1pqWXV5XF6x6RLutFPz9SQ7brZBQ6C2aHJ8l1k8Ehin61k9yIw9ekORPG
8za3m+jGOJGTNzl9FF2kPf/DSamDPGFItracPNiN6gP7wL3wz/E/W71tFS0U8Y3B
BN3TOOrURptAetXbqyiY3ZG+BllOlD4BLw9j3YK+n0KSbA9sgppZvUTA0Ufg07Cx
5gfJoUeBXKD9NelCtim+l1j+ZrkYmRprjx70qEv4zG3DMarb+Yaob6X7QafLzyTy
oLvMNH+Meu1pcfeMqBfM8CqLazpGsgCQfMP2hSFSYFjXql/QNY2P6uDkU3Lxm6Kb
fKcQB95AKXrVcgt7L3dIqcsNYWjrlQopC7BnqtJWBRDbkAySCQcWnsX1H1R1G+aN
K/V9M13ImBxLbDcw7hVi2u4X7aaYZvaSeIoWzPzygr+BtACL0hT0CFYyb8Q/89Cp
FdiaT5iO0UkCyLwDy5RL9jPUI4fZ1Epp9v5DAvWyovMYXN767JeHhnpNVvPqU2sm
EeIxYKHxXNVRyKaexmRKmxfRhoveHDJhatN7jw2vzrqYbhMOshc/Qnk5CEgu+GFf
omNlmweMJUCbySu0miBuNFHSSS0DzFSe82VPPuDfb8W5V854Ogih9PK2n+9HAMn2
godwe4C16eYbTgPOJc/81P4IHgy8kzyXRrhJCYPp5Q0TRWzkYQLZnjveYuU5wbZ9
eodsLk2TM0MrMVT+lTU5RxWIXQW0kMwXriwIpo/rid8PjJsn4hRcP3ab5AcOgnKQ
2o8RUuqnSTlzEQkA43a320u1LpFsriiSrG5eWgXEbmOjvUKC1FXc7ex0Djw2Wpe1
9p8eYYoK9Xyx2g+CKBHXL1hGQbjMwIxhm5831+KO5PQO5kWI0syzMV26w0517BNy
QIFmm1FAAri+/YeePiB4BESFLF2Dpl+7lhaSax4yPAkLhPmhOJaIrUb6OGm0TM3r
9pvMOmJ5Q7wyFss92GGPotnKqY5f4U6waIVl6rN47ewIQQepinApQUiCQ0t0C/OM
i4eOqPw8wCHy3tAFL8pRS/hZ4nQ0ES5Bgz5O6NFKYudS59o5GK5N6hx/3WNFlFBR
Wu45HmFtCN+NZufnOjdM8OaUM4Ro+8w11j/dMTMu1pPqmgtDmfM6A14Olv8Ws1ZZ
UtQPmi05Q5dYCIzScuxV1flDfOZOqWjD9k3z2MgS4zQPuCpp4CjFLz7QA9To6veo
o0cKb5Mv7wJlbygGW9FPDM1Bn4fvbdpAvTN6EyzixeUgy/glL6e5FeVrMLtr3PoG
AG3sAogfZiCgVk173LwVP3TdKqQUdIcIbonX5TbYzcgKHVSTMXMQfh/DOMhrY1I7
8o7ZerIzUx+cR4NipWZJu3Tr/DSuDeq5qlZ6n3xPqmjawcENP356jNt4+qQeCjao
n1PvblGmTUNdnH4kdFIN1YAfBFvbZSA4H2raHzdT1aVNuGLrDOUbVDmCV1qqkw2x
vx13ymAqqGHKvpZ1H53i03mgnuWsAyGXAJ6kaDON0cxmwS/X+Tbhc3xFg6S2rLL0
ZoCTglTYgA2Lpqhf3xNGoOIQ69VwlSrctkk43LutpGKX6k2FZtKyc0cNtKeJq+Fu
jG9Nrv5v9TCCIiht/n0KausObX0opDdOM5uzJ8yeaL9RxFamEsKk5fkoC9X9iQcd
A5/cwz+VcVxmTidY2oaUa0u1M4ECYCvlHH4lF5WjqRT07YJwUiycY8fk4JIzN/4M
VW+7El5w1B890KD/Tglocp2xP01iOxbdFOW+IFF/oEbV5f2T0Xox4HGi1A1Jv5Rb
8tIwu8V2BUoBjuelzfvfWVajtpFewymUZXcZ3psaEuC/wo7MpIyqMMMwYPM6KFY1
YIMOpz8ztRGDgSjEcih2Q1qPs9EucuO1pzVmQKQN6wERbJ00CdfBnVwTC2w0jbPO
XvcV0f+Fqt+jhQA1Kfj/2uFHj8XUW5eHXqkxAbL/x8dtmzIjCPjeyO2pV07q1V+c
XzfcbvY5tuB3Njdf5AYwLSPC5PObL1Q105/nVBvvQ+XZu5kL/NR0/jtonjinA3/P
ZSFMsPVYcnUk96fyhXJvIPbvv8wH5LQzgjFFpaLiP3MpmrWUJJ4GxVeyQuoSYRsB
dumEUtEKtallCn7maRjlnmryKtFqtFfCBZLeLjVHbwtMf3wKswLekED7h4aHkIrG
aITkO/cjU+LheGTTvG/f42VM4vj3QjzapDeN/IvjvhyoNVs1d9WIQ3di4xZWm8TP
OmdukSIEAUMVL2Rv3gEkuUqL7bfiFszq8wg/TgRu5TjgaRiJNW9L8RBdta7wFkFr
0m8kHtZ/4Sovam7d0H1oSOCSRGxy1iUDgFIOiCcHAyrDLiEjxyQlN7Q66daSKVFG
r557ViYlAUcTKMGLlbXHiqweT0RpRtfPkkzGT9HKtMFzybqlj2l0EgWNnme3eO2l
6918UB9R8ekaQ8wJu+WFtHt+KUkCTnUOAhSgtmsVQyo1/6+FraUvbVKJ3NGX0EmK
UoJZGlC+MmOU81kGl4l9DZayMChyaA2UFrhGSwd41w9b7vvsl+CQxckRfEecsSAq
iWY4UO5BkgEtv4NoMDsYIUEtOGLbgyaIHvvLd5WJhbhZHxcqmvOQdNsP6PAzn+c9
WCsYSR1MqmOUKzU9x9RS4hSQ5zUxkkDdHdQAQX1jgSzpGsXw4z1AsCK7s+rUslKR
2l6T0DKQ5kbvO2f6CUSWt9i8WjXzC/xUNMBJ8m6UouaKO0v8MeDhOR3aSGf7V/zt
8f/fNKOfjHookqXU5dHCix/FCa4Dt4J09yyXMcBYQ5+INLdHXYvUWMmGyKQMeesJ
ifOltgxjKF5GmNrVeKDUENRHrG1W5K0aXiNzVBOn1UueXITKWqvIOAYC4oAKJPHp
WkxcaG4LuT93OZm6yjDZ9xGLN630brZ+l2e1BpbJwLtlXW+hgeGOjnLJvD33RzzA
/dD39YnUq55HlUctvKTrKDGVkMcTUVVnw8EdC3XTF2qCfc1QsjHxla0Sf3c1cjSR
wy9y/gPP/nCW5137Qwg4kqD2V4alalYR1+0B+PTYsZGzaA36LoPZ6XClLrQT0lCK
CZECCZdqilL0MDWp41AkuviDvFdSUoucq43rCwNABinsfDBR+RfRTS+QxxHseuil
8lM3HroNqmtMFIQU6oR6QeSimS2+NBBrC/FttqllXBppXZ1PK1P3CVaP+zbX8/WZ
beXpbuAi6AS1QirIQHkGPBmHIEX/IkXjosgisnaQRJP/hmSCIlIUvi89UsWk7ChN
/YCh97M2aN8iSYb4uTorfvKdoc7DflXz2iG7THWPHiyurk2g7FnfI4fblsrZqKlT
rRwRo9Si4J5g8InrOrs82yCcrB0hPITcFsVWFjR06U73ruVsmG+uSmzlm+dCtsz6
qY7bps65h3CjRmgBAtLV/ZNwri/yJeKJQ7xKIm476usP+glMC+eSGbHrowdMhidy
+zXrEIfEwd8BnJdQ2Go3tKDfcRfha5F5j5sp4FSjl7C91MmuLP8i0PbgKh2lXmiK
IU+50uJYZH4xvt6LrxGFUJqKEYukT/Gbekv3YPL19WSdtGf8hdXU3on3VvX2i1vx
Wyt7sXED72PrFnMTZgfYacdWLe0fCjNrOIoLG+z+SRlCTqzWFbGIhnTLlvk0VwZD
Gy55vouIPp0EWKOrlGmbnlpXT4wD6LldqEEc3Y5f5FrWmZmfkeQ6Ihk1Ox/4I4zZ
8NQAVnmnlYfkY6UPYAL3CyvYhN42b3ItvRBw+XOdOIurZ6lZvb5eLaBqOX9H0CE6
lA6Y/ghkfXMXKb2KV8pYvpnsOTb6lfRh6r9wnO/jfEVNbfTXA4QNGkF9x/tY5SSN
javxuq9m8or2b9EDpoiWCdIZx12EYuAPPZ6dKZCAK6quHPKUkm3pKggvBWhcVJau
GFey54FhoB10Z7slWRmjAQM27oaMPzsJPrPUMvdedcprWTEb1ou1Xrf2XmZ8coSg
s8YpjiWewbJ2t0FNN2HUx1DOZY0eLTlfd0KZOHkHrPOTaw1nd2RTgxJpHEXMOCZH
gf37p8HS9Ebfainub/X/xgWUBlK3IjqwU49ozY/XFbe0ZxD+jMDindok6zG3O7ht
/RuKIhcvrPxVvNSwXd4Sikvc56j8AGla/5uAn5iwBiiLkueSPvaMmRxIeGXMqVj+
QngfPOtuEmmiXg3eCC9z+R70SOS2WQSveZ6B+vSeyIoMatVEAWFZYhhe3KX8c0CG
b0nclu7MzIf3b+643eJcdCxSuW98qXvArq0NXHdL3VIwzHa7b8ojm1Lnv2WjyV14
ijLQ2jbHEhhSJ5sKCrtyqMraX7GGTJZp+Sv120KvnzIzhJKCx1ywr9sT9V5H5VpG
97i+TQqZnEeqNcI+ovskkT3geuxiSnLSQ8eK1SK/MCSeV7p9srb9yKdsich6dXVG
oscalQHJ8BH1DFPa9ykZ1PkdHD5nMbz3WRl2eZ+RpmohuU4By59tddYJdVpajEjm
kOa7lxGjlfH3ZEfmUILpFGgyYCcS1hX0TyAwFqeb46nYZIT0r+SMmlv9iaEiNMdr
L4wMImX4dPaW6Pgukm41H2diPcIV2S8p9cXPfQadt1FvbiwxOf8G5tUJ9P0I7cSA
iDS9rhQrdrcvTtQmCpCN5a3YAJ1BChJ3QsYM6pedoXcGHOXKvpLrPi3yfP0Pk/+M
a4eY4SySje5FNyRFp8prOQCHYjXvG7PfUo/aGBWA2/mk+SZ7Gq8o5d1ALVWk3nrr
ftira7plWknuv/m8PbZP/dZAqVRb8J2EsVx/E3c52Y6CAUFA8tcgV+HhHBpe4VOg
L1HZ5l4/fI4bYwpjN+GsVWM0zn7BwN4/6R8c6unttGVCwoOCUlIfg/f1LFTftZyS
1eMekGK/KDcS4HUu5QAHOQSOe6Uj4UT2rjs35LJSq6xYcKIBy1kdh3C6a0SRWPDv
MkAXDiyjkf9zHG6Y4Ofx30Q+19vCxnxJhzWWlhmfVflAsRHPwVm17/atMfpyGbnn
wkTZm3EX7tQFBueyqIwr6y3AHSOLJvt/Q5vG2xWjUrQScK3PxVYPfRHr1P/hhUzF
ydB3ZpeAxg9dWBUz/iUSXMzUpmeuM4ek2m+xooqBqmR8z63OUhBAzkia2N5+66RW
/ejLGuDZo6JmBhOQH81CV55J6/5/y+WP6UC+ntAkbv2Mr3qDmR/rUri0VDIcai/s
pO4eXj9+ciMFNcO5Mx3TnUBmyyPDBpicUdElzkhL4HFy33vfxnNqR+XwfVCDF8IP
oo/+/48ncpYpfUTuuvdw/CEOQ3GlXrl3ysKv+mbCZ1pocksRCT4/jaX18S9gWjf3
HCsOdNh2sk4jLYQBV/aFWr00klLSQwfAxKdlFV+rv9RRoUezl0+w6vEsaXg2g4Ut
WmVD31eG5SbeCfwSwKPYIG3n63z+oQ5h+9gDtq8cq9A4ddBfJYmkgSKyxfnvf3Og
AlBVSTN9C5EjOPFabrXESrAeIKELXdRcS7K11Q77cnM13sOiAEpxVGHZa3/HaaEU
RJ340QCqBZWGSl0lbwZso0/VPHp1pc/B+TYftZBybzfSIiGtRSwsdCIE4PijPpMx
DbZlI3WDZILuvNUI2BmUOTrB69bodM3SzbwPqQs2jWWTgqkl+LcRdAaDVvQi6PKI
1kS93KhYxnTSa0ZTaCxh4WyfyCcK86ZY/FTTRrI80waDH5xlzIv7xw6/j72vv84N
xuyZEaeOt05KoPKUMtrrTPlz1+K2E1T7k73jIlG+kF3DfmG8Ku4dxJtyBp9kxVHj
i8wjBc3TVXfqvM3/nuZr/YivyUSS+fzCJqvsAQldWx4FRebpv5aUN10Meccf7xjR
VTcdV5DfP2UYz7XZBW8Uemu3fLQh+7Nvi+2FHemsr/npeqAsNUn3kgdAfmoe3rqV
AHlnHCd/IQyrnl03KCqxDqjGb3HeOglaWewLN8l0PSEFgumsOQg988c9KmvrHCJ7
j1mYA1uqvDNsIHZEPge6RG0iR6IOjOU3lw6r2Gwz5bpYUhkD/NjI64j3zLXraUYZ
c36pimanPLxHp4AZ39CHFhwJYAJqfQITsa5Sh7UtNgEJNv9ZMxi3O9JM7GSLJeOt
/y4XCXNTy8TaTqGY2vKEak9H4yt7SgaNmnf6AUAEHP4+SES+PiGmgvRu30U0uu/+
t1xTj1prFpNtcuF2BBNYDWYxFyKXa3E4g39/Ise8EHAl0kwMc19R/eZXBn6pxXue
9BwuW4WQTD4npRF3k1teSwoWUFfwlPVwGUXl5e4ppei85OHx2PeJ4JlH1Ksv2L26
lA+EF7WHFJFIypiF+KUrlJB8CApfiPtXFfKkEtRfPLq1g/DVelXObV7+kAVKOE0o
budRigANRAm6ogaKFZnXssCmf1idehbKfHnPVLBMjRCQH7mNX/Ec6+LVlrIliNjM
vlOoYJx/CmC1GG6Hn5aQbzo3sqodGsiX3XjxHU0Bnwfum+mE0vcg1MbyVp8A2AH+
ojPoOU5DX8ypHAqUv3zj06n6b7fjd/8na+itE+piw1Q0piSFWvKOe2ATEJuaG3b8
RfjdT2FRJ99mEvM4jbT/e0LEFjTlubyiHsxNORHa2GPzGdaTv4WgmG74E1MM+QID
OnGzJ92K4OrTfgUP2NIiWApgcB9QVQJE+eSH64Bn3ZXnsJNXqxi85F6qGtalkwaR
zVplokMB/1kfgU1TilePmdrkXM2RQptVA+UzKWPwTMMlmymg5IIKHbe9GFlJet8H
ompMlBFCdUFNqBAGXiTJM+h4f13WoybL4lvVAANPyKzRfeYMZY/zHF421KqV0Dd/
mFkZpjTtR2aQ8bjDWXrGiA3HHF5H9QG0a4x2KapEqjAtYT4Z6H9FdH5iXIbd6cRX
enSi7JLhqxwjREraM3scIkEsP+kg9UlNtsOeOeNwD9YBi4+0EsJp4ulQmM1+sLOD
mpkoOZ088SiSh1Uv386Djg1z2J+NwYNh3deRR9XozVS1KaXW9zxmCYvBSOMMdgYY
J1dRdJoDFGq6xB7cxe5If21z2kCiMLqOxkDkf6XN3mLRysl+tWiTCWeSktvZI2P8
AX7h9QP/GrRvP/Pq827wb1YMkR0GOfG6KPdUEQzfggBgnNmTempeK5/N3atmMncE
Qysk09BY/dhZoNlNJUPl0FUb4xcTbpDmnhVnorygux3nR88Ha9q67q4+ohy9qASD
MMlG1KDkjTklXnAoSN29a0LCSXIi+LIHGloNZqi+8yKzqAv4BEAO4GAvb8bi4vLE
36XDXPk0yd+RFVZNXCTAcJEO1r6hqO6aJiO4i6CeV2tRivhsAqj9BVcpzeCvtMPh
gVc/j9XcsjWag/oMnIynvnaI/Yx0AnMksmrkmM2oXzD4DXW9iNBO6D2orwd9mi5X
izoVpok+uFwtcv1p9vqQYyWGOYhlje/wcWtthqjxcvN4GTp1JMT3vN97rSozHeFV
MV+K95EfbgFWpbyZom5YP7nJ+WLVAJEo2a6EVRPGRJdMFEsJAT2uE/r7KWo4qD0Z
1OC3lzrQbuosMxWV5n6QS0jtfzEJiz8RLewKFD4EvXzjiUNzzT5KdiVEa2zRGLFh
LKLYnEheHw3SzLTO8+vFd1oiRdwCTdTirs7yBSIMDpnWtOJTQEyNonjRYnhEKY/1
XX6hTSFwdrdUDq8LwYISVhwDu1cWvicT3BAFaa5Xc3l1xqLcWd4Glq+LUJ7VuPNv
AZZE9+4lCWpm6sFXzdqDjNbTeytyMMCrfL9m7agPXk+5dK2bBHFFXgc0MY2rwPcY
5/knbEjVAl/2V85WSbo6JzBgw2gPn8iIssAigdlJHNHGKGyay83d/cCvj91BtWYr
N95yl6GemaKPkxvlAz50RE7ueFRf/3ApPKMIwTIRzzUvKifrww7pT+uG6FndWVI7
38paHj/0KwoaBN2rxF88dwrn1r1pUBpMFgoBGPIpMRIkoQ6CYwG4500Px17yAy0v
BU3dABXCbZpXeydf7SO1gFAAIb5DRGkbtCXfmz6X3jdq2oGOaUniOOsBOdqeAnwH
4/P+tIEQonm9t8axkvl1Ix3zkMe+RHCTWUGAijtqrnNUf91HFXGAGczUieJYrgiZ
zWtVOPjJdPn0+pvnvohAdChsaCUmVyyDeJG/ys60mc8cbaHIq2ShjjZTDvB1ModP
JKIUxuDOwhmLqVw6PLPvQgOY3hCfXdHrcgkdacTsmgzWy6q6DnZZflQRCcIKdClk
tEwd0Q1db4IjQNaqC29LCK0Laj8rbsQRuTtj6DZAsYseepTbguAHXLmKiYCQXD8M
PrbcYl8oddYN+B3O65nF6q17fzQ9deJ5oyu6cSXuNAlTCwQxuXHqrQ9VgFy0bzd2
xgwnvXOdn8VFxe87l8XUoGuPMkOYtZ7BEAZdORgkkAnbDmZK1K1lSBGnYZwkmWQv
3ox1bsoluP9fuGxxvyXzSYVdI1atM4fEJ2wN3ziZPKUvv1cNJeyk+R66FYHZK0om
Hbm2JcXkSAKa4f37WfgO5An1NUDCbmTZwKpdAVfdSdxPN1OXJIoFditxGQroHfRu
DZ0umRR2zSDV1lQ2F5jid4nSNsHRLG/jXDDs2HNbC0isFH+y6SbdNcib2fSJac4Z
4ukH5FqBB55SIPylxblEoajRCLIp8/e8FXRPxguAh8/qaksLI57+9efvSPOR6BFh
1TltSKVolRWVWQ1vsxogwcs5pyBiRWFmkFLxwzTuSe9fr1FA5XQjd9GUEA79YZfS
f1BJNUbsf7D0zevOYbDhAXrGvTbZeBOWJKQozB0LZ7wYBRkHl2+pVriUy12jeKpG
zHG7En8VFzIb3cvitYUiSn3FWJ+jxJTJVOLSor9gLnaVzEGih8TXt08JLVDi8ftW
D5gkY3sh7z06CCYvY8Tchjn2F92UWo9X3E2j/QWbBrK1Z6A+ur1qnEzUf1abQ8GT
D1bkaiidMNijPoiNmKMTzkexF/vtObKnV8FwcTesO/xYeVQDAEeROQN5/5R9q0Lp
SEemUkkAuQO5+CBZw5vW9fXaw03A/rrXgHENF/OWZ1g=
`protect END_PROTECTED
