`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Cf03xtgXWgYqoEa3W0FFjnxUXKObjo9eSevoxf8roXRKhqt4T76xU6s2XonuLBXX
rbQK71jlB7Ji48EK1HtFrPyrW/lnWlld5MZ7ZE1jk2iKiZWRRcn+qODieC9pN3ir
O6tqPIMWiSajILdphQUNxzwdg0SdYhbSZMt//mgNyhsIR5GVAIee8Xs8mumMIE9q
NgeYooq/0gja+nid/Z4SoNmFNFEeQ7jnhPgZbPjbedL+NTNfIsldtBvUdQaAC2Zm
3DXyf8pXFVgZZenZjbenJKBBpfDllNBZD4ZIKxFa4Vddy4615s1Cte6DIIcyaH7q
3uRUX9fzIDzMkmVwNYwI0rNvWErLRdzsVVkXY3dQWOKjOWocSkJfAULzgVDO+DHx
ZcG0pLYYMZK3ouiA4vzlb0zV7lV2PuM3ocPpfiLrqYHX0LKk7W33ImcY+gsmUIqH
TLaeA9BGmOUL8hXics9bpe76UIgGXVJvSh6o6kdMXuta83prlgIKsybHLGwckl4V
ktqFFvelN0WTqrf8crHRiA==
`protect END_PROTECTED
