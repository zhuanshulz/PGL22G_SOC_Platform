`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ofalS7xAmHxTY2sdCcWP1ZmwntPTO/i82fgHG+ijICVAPh24ikwuOfkH6Z7OZhr8
VGyRZz2CweBlCYDsQbAKxvEEEJfmBQhcSJwZEQepy6LKhIYx5lvIeOWK+DjgJiGY
7IRQvO+TKeiFcpwc7xv84Y634KX962SCpsqqgGNt2TJHW6Lk+VjMJtjeM/pauBkT
900OgFnM9aPRd7RDOy2sRswBJdVEW57fC7HfE1gFB0i87wmN6GMqZXvBCEeKe0C1
MNcU8F8XWrxZxmi172K3gMEFcIBDHsy7XUvAITvQ8ZmuhZYxKEXUcZBHLSQg5VbJ
+lgE6Hy/8KxjfdJafwAP8GM8wCunHdso2XipirC6fcytReD2F8EimJZO/3d1E67t
AgKcBubIYoUtK9bEeHlhcgPf2NDTM79y/NDiTVCeSzkE8hZrnAnWj6Xsh7sWIFLB
bh3eie0Zq4ZRgMfvtwfcbLQfg6yPs177gGg5Q1tRkdKT5rEFeXY4bTGkHo0jqC+9
M/mmnrLiUWmDoug+Ej9sJ4rrLJapzCB1FH71mgl9k0ZV9JYQ2oABH9cmMJZqR3zp
Sy0PIR7AXAGTtjU7ofwpgASgFjmxz1wZLpAjQHlV8/C+1FyvDWmmO8Yy73V99+UQ
zK1FDm1teZWxljB8VikttAQ7i8DJEQ6UI+5DcI4rnsPgRugvCuw3pSHd7sEFuzBz
H4ngE5BnxqYG1yvG542geKLzQVRrVROwiR1OxxMjVzrb1Gl46pTd5cHzOnc1SGSi
tuLXYz3qUzTReKcWaIrgXNhC4ag35MkGQ5odZDiOpYS2diYag6/ISCFUEInOyzlL
hsupHgbQeJZBVSVid3zsDVJT/1uUZE1izOP/DgXo/qv+Sv8v1PtlDQ1Nm5rfqFE9
Ouo0MIxPlUgZNvtUsqUCAaWbsPEZbWNz8Xjwxov1UvrfnqQgwCpKchOtona+4nO3
limHJWzpNJ6lgeNLMViSa3h5Bt64LcC1s7D1p7VdFie/tKxJQae1l8GVDrIQzefH
R4XatCHwZLyjVI6VMoK4AgPuNAhXj260fZSvFeg4GUYy6k+TZDwJ+KzmDcUnJ3wt
N4OyNnR413ojPPm70mN7PaVlzI2SEGGcXDoZbvF/gPurmlxgo2mdZpNzR881K6lE
SFCBuw2Ihju9IKgyHjVX9RWBqyvB2LH91fqHHaTHrRilUwV2TcEFfR0eTK2Ye0mq
vPkddXE6qYa7VMbs05dgCsN2LGRP66LG1L2vYSR9r4nyd5KKBmiTtfRwGCWh2yu1
3Eu+Emltppu5rJFfnhKT/TZTSBnINRH7Oow8RLD6RlvfVimhvrEmtiMZbAFcDk5g
hkpqSY+07y+8J0I9XnAHL2EPy41tB3plu49hXRM8pyNBpq/dpt4thi3GdPVqGojl
gcaseCMHh+sFJT1iRCF7ymtXMqRRxW4QDuNHIdcKMYQCD6hHaMlRWqkGPdOMfAnr
hpLBqQW5dazyXOVWDRX+b/ffbZB4R52HEeQaqyUC2KQ=
`protect END_PROTECTED
