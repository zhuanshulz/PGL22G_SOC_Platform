`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nO/0jQpUjgzAuMclbw1RxVPJLBndFre0cABRSDfAWKAi2Scqlm07v1XhVBYVGm+h
tcavJWQHaSYRAiCVrTWOtz2Nmu8gTbgdjUUEMOHjh2XBZVXzIQgNjEAozUzMsoHA
vmpSzKJhNUm3dopfAyhk8TdvjXcGXmj2Ef0DCObpG/wSPf04Qr6Z2fyOQ5rXWCGt
aAmTdxLkVQSAZIcjebum019XXAvpqSAw4sdHb+oJvOULq3ydgZSVuazTOBAH+cht
RGAvcGppTbwcV6Qm2qkKu8s6F56ArWlVAJNWJa3YB2OAp9lj8+Iyjrq9pp2JIeGi
V5smuelPYKqnBFfvuwALdN2HTaBzOWM8LCjpFXlsAHu3znDeSxAZ98a4Ju5xA34n
s84+oH2IkAyqFBXfQZTJC9zYfIU0DPElw9AR1ce88R9nCmcKUvR2iPU1ecLfN0ij
f0EzoN19WI6a3PaRitWApXu7MDZW7jXr3irAzb9HK4CZTy7qQtuWwf9SYYAq5Kpb
cIHa1fABT0D8RXICQUYff8nj3A4o43734aD/T4jbG0IG4ah9kTb4RShw/OlS8Veo
pfVTp6zRYDZ1fZtGKno9MAW9oUVrEWCiv4nxnZxBArvVrFwaohmJ7bTFPr3e2obk
dSiljBo04yt6p1T1nUThrPjotVrOtReytnhhc71gjrqqy9Z95RcZ2/QlLRvsqqhL
WGWAP0wbdADjgtm6LQFJIQoRCdIEx9+kSobyM7Yd7QbvKsqdeS8WlDQ73/IbRRkZ
iA30AknOnclfbW7OWec+3Uvx0jagFCMRyInUlmNR22o8DyhOcIRSYE8p9keVc4Xf
yczxRP82rbpw+niDrpTM/Kg2Muk0MDxvK1jF8GTsw9LHVBQXqvNJEvEm6vHhAsAV
fwDpGePCV/FbCoiTsagq/WS0uE3i289Z4h4wZ2t2KgZkBQcRljdOOYZrrZIqzc/3
IZbMmKEj2NI4lN0LZIuq8lT1WYg6R5GX7DoxA5IKsFfjFCuvzo/Tsj7Nz/Hbd0dO
DnxR/nfFYqPGvQNR9jLLRghX6wB/CNmCXnJaZnrPRRcu0vBkQSYOzX/lX3AzQ7hR
JP98DHma1jETzk/qDgEMcxYJc2Blo0lzI3Qqb42LqsFGkAv+VOGQ17+YP/Tv5x8u
dUChoga4oLC1ymGARqi/B6S+JRw523gwzCKcVwT05cjCg3NtPOvhc1zyJR7ChQs4
7CMNMn6c5XR+qxHCn94iNyVb99e3NoW4zTPT3ij4YLPkE8XLubyU6XMYVKJIYWM1
sh2PwHmWp1VakGH0nx0/T5+Z/VYE0w4sEBerfctIF8EsVIPFqmo9RszxiJGhaLtg
9PbxVwwo95KAXFiIytjzFSwLIZR1MM82/VKqbOhi+YciwH6oEIZXbGbiUXk+yQuj
BJQ79jaDunrcmQrBlI5uZxISHay94gV4Hf5nbd92e/Ugg9vkWzq9zOlhC7xo5f75
p4LT6p3XYwFcbLf/kk3X5tZNOJpeoZzJiw/Jq1buRlgTmfJTRwAU5TNcPtxwiZ0W
Pw1E5wmhQ4xJaZeXn5qBwv1hIRc5/LFYj+FD6QrkbHDJA6oDkS2uxnzgWXpaeQ7D
s3KLJZvJWmwihEa43XxzRrX1VEHRPsJRDYrjgWcaMlLctrl8Aj85v9x6u5o/zkRz
Q/F7zPD2meLIzKN/1JZ65GxEwtck79ko/n/DLwBJo1RcjGb2OlXyEijQqe5a16HA
IZnHJgTGEy8E1rUDP+tX4JDZb8scluU0g6jUBLBqiCC6w19mwOrox3t8OYORItv8
RuvzL5/1lrP9iA79BjSZvoLTB0aTEaSd5cnca+PFRJDiRD+17qt7CzWooCSfm+hX
7bDeMD7L6YzlLcEhU0wV4X1T1TloN3GIKUyiPwyUiNgZM0HHb1dhD2cKjCm/jnkC
Gz+7L441LW7mPKs4bt5yCfgRoPg2oqjfLktSRB/YX9zXn7Po9aa5yu6irwd34GT8
14KPHsLmjFFqW4pOCZfXMc3jzRGgyU6ufY8YwsnHoev/YFzuu4lu0SNZtGYcsYEG
OJ4M3yccI4MN5ooTJs1hbtwl67JDlIslXszoRl3XjKUMtimgr8OWChScqMBhuxMs
ThTCSQlpij2DKRnOfQWlcEsVaooRpJ4AQsGWArLbta8+/gWPlUZGB8jFQr9P27wP
i9Oql1SyKrSrgoMujYD5SI0FtRSmyAhICScY1KhmXU22kxPNmOZxtet/H+MYARro
RCfA3h9wdbVrzixZ8/lIRy4Gv0UEf6LH7Awxbi4eEbylB1jaDf9TubusRSBuHHeC
abFpCd4yxvYnijE8RocWkh7qpYgA/TaHeiz+AwVkVFiUOWY2s9F95cSxa6KrYCSv
J/Ae3h3jqaO1dE8MJQ/aZeAIIA94intP7SQ1uELmghj9E/O+vRpg20Zt7H6rDsdO
qe/axOaKPybL7zEBij04CxQLKB06/3IxyrUGr6Bl+RWm7DO2oQVgPnMVU5M7DxFl
DR+Z8lYD+qwjiaI7p0gIchSGOU+TkqbiYCtmxOxGOFNweBqfDOaFyobXY26gyebD
R1KtZELWFUQElaaGp339b/OrNi1boWO17R7lQIfuACh1P4xfrkwpDCJjdH4VNrTT
`protect END_PROTECTED
