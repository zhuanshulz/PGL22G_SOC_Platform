`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jW1djgOv13oFchTT/oxiVT6IWcFDp05U4+y9fz/SGmWYsABZHcihceVJtg8t4Pen
fompsPShBZX8X/bQDe69885IIgQjH6jagJOJ/CtbAfc4XmqINevXg2h3FIu5yl8q
RajbqIbINQgWrkr6TrULIYi9gIg0t9XjWTgP7HU6eSE4Jb/5KoT6EwgKrtzwrjyN
6KkowOr7SsoLp1hmCffoLjByK1FnQbblAcLubD7vKVcOsUx14Exyr3t0uXMSprQ0
objn/0Zv1HQmNE3lpNfWg34EMkRHi3nSCD8bnVlzomDeymDZGPRll/HIoD8pINB2
jMpxrc7s+icWDNmK01NaOaV82yszd1vHvmjB9wGc0M2FDoLSlVfjWONMPFro8JRK
zAB+D++fwMT7UmfklZA0PQgFySw9RZry6tvH0jYiVLLRM6zJDCsE20R0dz5KrpjJ
5CFh5ooKLWXuW0w9R9WSU0LnauwI8LpKuX/UI4y/QHI1grEdH+Rjm8KHcMzkb/F6
9wvgnctV2vTZSyVXqnoJRU5qZlAUPR/i+svGsU0BNU8dCkP18XyV2wfYDK3zb66V
RVPOiJqGPNdYYexq3ZeTkGhHr5UDfehyY/EfF7979fG33xlWRTxPqfDvFocwWeMC
V+FKFWV7+9bs6RuaafRl7+7NBXEoRyPj78ARY5Lf6q0oFaLpqm2qhbVCPvaBwe25
RkRxyUjFqXS2OVOBhyEhs0uPx+z8hUD2fgIls60k+b0=
`protect END_PROTECTED
