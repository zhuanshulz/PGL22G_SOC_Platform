`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MHzjJOFaEvkI9w2dFrd7KmMJW9lRSTelH6yu7V0M3nX4kqx8Y2pRH8ywwOxfRGNp
axxbZiztW/gYJUqEm/LAnVK/RQXtHRaeifUXP017Mjmj7HUYVWoixp2Ipz+50oS9
8ZMp00yG/O8HrQJEVd8C8hJ0+DJVosHCJxMy1ZdLcY6A2/DgfTd6ixwXTD5ViDSd
h9mpGZLIMgqB0MGnjcCn90mzRXgm6ZXZOQvf5PwHgLRoyYvpPMV4XtI5+mUb7IMY
3ODtHggCQYqz1GHnzIIMRvkiBBxbTctCPkie6gKRvegc8wcBGByMY6gChvzdz1f/
l1i92OYOtO8Ji7fOPbpYm9lOKvKwJKi6DduFLRALGjQiNC4cFI6Nvh5Ki20PMkV5
C01tkzNNAfz9XNt0/tsMGzGp5gvqmnRWKzQT9tNQ35tLkOyPWbeL3+rJMjGggvyM
g7t/ThfPwbrSVOuvLuZu9J1OYjup1ZlLr6cyUO5+1vybN3P01214vn7n+TupyoMN
9wnkCmB0bHljfVIyl98BKUMf+V18Gy0m2B+t7bdg9auvLo2sOBzOFk55yyIJpzot
umukiJnngPElrtOsq/I0k5mPoHbSLIFcZpGxXbLRyx+ulEIgJrfzfo4H7YwFVfwo
`protect END_PROTECTED
