`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fxJ7pLcsldUywwBl/lH56SCWsJSUpDCAB/WsnFGerkbohLW1YrrncUQqe9tGwJ19
8HgrzD+uMpVKu0d5Hh1W5x8GYJaosBVL6+avR2HAzBWCtAbJwUPRzz6F6XxHJ1+o
cHGtHsJ3Q/N2ZOBdFUXPbPMKqFYXVd40yJsNCLwh5GRNw/l5lI3cLVa0lZQbj9vp
L9NF6ezsJUPKPl4762PO6GFsCwIx3znMy9sPoq1a3LzU54GofEAIldjO+PwujKbP
bfIM0MkaPwVzOvl/qyJnFtV/5aq7CX8l0XdoCRl3UAzOejT4lQGOIEcyGUKQ1D2e
wn8pSOJARP9INeDZPj4Xk+YciEJ15a2omHZml6eRLWGg7c3e3lh2i7loY7unFV/h
04auREv0RB0GqJWYFDcMAMaRnTUNrO17NFQ6ptHniZvQsNGe4B8x9362eSAOaqs4
Wv8o7T5VXBE85lz3EKZc4Unhb46burl/XK2UYyTb776+lKll+OjiGAQ3xOq096Hm
w6RrpwoyB/g2uhXXtTu7+kc1SbDRiDLe+jqjxJfqFvxIPZl6e/R0r3lwiY7ezQpV
8WLAtNdZfJpqJverLcOnbJVSnHZtecX/PSbxjH5e5J5PsM2QweSHLTWZYO44q+EQ
t+6TT+HLq0oeW/VF75dk5hZreSYEd4nUPaOzy1lrqZDtSX2YCJZWtZUegMpZO0Hl
IZle5iCqSL1kpgD9cWetappdH83VjkE2fVXHMF4tJ9CtbXR+WbdGGXPEmtXqzUN3
yCtN8LkL0TsOVU93u0aJNccxFPEdXzuwQhy2Pjsfs5GgiczsKBPcNErOgscadX+z
BP8SaJO0aLo9eHhHP/TBbC4ZLQk6NCOXIOfFLKOcNU9T+IGg3xCwhkIU+0xuhbWM
5kAnn/HYQ7SuvufHWDozCyEXN3x1jrZq5LSR3yLfwJlYwXL97nKPpPIptEgFESOF
XhJrjtmF69IO5bc7ZVwG3uVyKPs8OyI0Jjh32TEqaEi+LDYr0oKb85ahsIGAzfqb
T7pZqHyvfczGHn1DRirZZtBS8Yiez2rIcikStjNtZSHY+m/XvbDxrIhli1GDwGzo
z5d0WpJyiljssDfic1wv5n11Kr0yqofFz66ojevhawrilQRCcvO8hvdKFV1eM3Ew
WmqKI7tX0H8Wq6KplMqEgtBa9ZiB0BOyKBmh9QAkHBKnsbvgkv9ou+6toZz+QQou
rffjF10lIzezN5jUnFyhL2AobdI7pOeKuLnaQge5EpbgTaqXsKM77Ll3S67zum6J
+Suw04C5X0uZkrKI77EvZJC5T2OycJsW3QmiOMagJdDtLHV2E8AxA839QAJgJmcN
dj2avJITcDfjbxuPAhCoMZ9GaB+58oHS+wPEY/vQlcPo6P4Xoip3T5paMfR6mL1K
ke50DSOD+1GCBO7wchfwjY/rrvbDiAICaP2KfgW7aVAiQL93/y+t+N4PAHufBfSP
QulN9H+bpyBSlfpOsSVqHr5vfn8mvg9iJ+M6jrLuZXoNQVZ80uBRzgGPfr+UlI9g
Bn5R/vEy1GH3pbVoNIgTKL3r30GPLJGm2LwyngcFQC0nmLeiTWJOq+crT5fsq2BM
NELiXyyrf8JxN8lNOvTkDwQGHy2G23cmjPrnP+aVM6etta2Xzo0jml+vfUH0HimF
ZFmuf2Issuk19/Q4T8uKoXoQesxMoZmRtHiq/iXNVkwgHroUyc8JUNayCquhgeL6
0M3ULAoxWhCagmKjn3w8hl6G50s/shsPVSOvvnUZxc+ZwZ/gflQW8sUpVv7VcNbd
eKD8JRG6q1VAZCxV1Ca7QAawjIPaPad5+iOhQyqMAKafh3SIGgrDtFJqywzWdqhe
coh1SvM0Q1CQHo4QFvyHLZ7zLcBL+vjBhwWby4RvomTdX4NLOCrFLkc1qA/Nfdio
2Z62i408OBPHjujTXi7TrloJ1RiIw5nXw23rHPSI0cDCJ3hq1BDIfNRFz/8CqBAZ
aAVnX7uovNS9CN2Oh748dcyLC4jy3AH0QdDO87c2gFOlOx62n/kCLk1KsaBN1Uhc
flpEFvbXF9AlOtEZcGeJfWU5wSmzTubBd/WP8UeN8BZEhtdPqM7rrY5BKRS8oqKC
xHlii2cHNnsxXfYjUenoH0Q0fQ8zzlpgSiU3zmbwlFk8KDPbkKSWPrwF3KZKWQvM
pNtF3nx1koT7dj4Fbzjg817NWn3bPn8L3iLsB7tItg3yfuk6sF1q+i3UM4C9RYhx
y9/HXSuWTQUPuF2CFClZujJfQqWg7MJniDfgIUWsQwFbxuWb3JAghKeB/d/gsxmu
LInSH/6qHz5YdTgPu17do3GoOQV2Cjlf6sbgeAsnhJXi/BkZMqRkcgu4wn84XQ0o
TWqzdBFzznAbL+JH9vdAUZS0uQn7+u1hRfRDxu2oabEe7onB2aZVcKz7wtcMCMIZ
sRdiAdVkdPiKuHnikXSbsLm+HRShk5SaME1Gqyo/JESQBH0qlA9oyyUWPeZ+FC/S
0n08Xw4KW/vGnnxdTRfkZh4rh5oTcyU9im3h4xA1vYpq1TOY5Jyr69vwuzw+1mL1
Xrl2Rs7CeIyDgiKbuaVAZnHBDZfGrp785RE43r7gJL2D6z3YfMbclcuNRhuWUb/H
yYImLwJyjf1ZgWF1lHMtPvIMZ9xEnHl5zFcjcDVJ6xXcI2LHE/os5OrgBPBkl0N+
aWAt0Api+hdkYPKRhQWMLDDqkYgrAM6JY0WFKEMayf2+HOAaUFUyPyC2GLGwYpdd
vTbpquozD81+2xk5K97A1vsaG4tdgEWO4WU06lj8QmPwOLamlMSsUscRFGsrfFFG
ozr12/0VKnlHvMz6y4zaO8LGNHW5NRbrmh99jO5qN1upZEHL+ZuigWIXBg/cz3b6
OPwnj79CCLrMPnQLNAbUo5bpYg8Yi3qMKj0hqk1eQ4gyI0f3W0LtWrMI3uV1Qi5l
K/S/FCl2R2+6zJLQe+n9uhhd6/Kgk3shQPmoYSD5ct0jPScsSnfLsR6U0iW47Q85
jSrozbfUfcIx99YEwabc7pyVcB1huAX9ut+IHc1tzJNpYH1lNOq8Z94eW+FJMznK
AozfygLhwGpiH49WxgzCNvRS4Mro6TzVEdJz92iJjv6QMyOoKJcJR3bYJfIXCG6X
Nxq93vUh1w+xo66iOPQENMo77IlnbBR0odfoOS/Xj4tig47zRNEOMLE1DrWmOd8D
cbJXxfWirSg/9l0QklcAZBrmNI/C9rkyS8RELaZ5pAKhW0GOOOr+dvpeiGAyW7lm
Pvu+FkqyzJ84nFv6Ewpxmq/bs+hP6ZrZWOTZUF3B3L7LBXou6NGV7sKCeI12Pdzo
BmUCrrWAUBEkR4TCBuMPzOfeE/ODTS7WTehp6Vd2TqjdsdmxqOllcaN8Qa+k3SIe
6ub4RitaX4WNwPef+ZaddijbLhxY1OkHpwHhQ4xABZBJxg0oOvSY5ckVl/rUHVNV
CndU5Pqt1oDdNrwHOZcPgYJxwUMoanrljhPndYBqiaemYW1/day160EYmvLkjr7P
BF5o7QH6rrUhHP5jsSjEcYcJY0gm0dxwzCBvtJJjQv6beJnXbXnda1OT7rU96U3M
YASmYbRZKGGtHXAzUHSWOjpgShluKXZEBLPTCfvjvwzXwsxgowmkVio0WcoT9OaE
77jzGEl80ssy0TufiyDFh+k2BjNYZubOSnD3N7o4iXGxHVfbAKzQ9Dz9IFLy+10I
aFcMqfg1Zl0lU/oT1m3aAC0FBGxBZfvmjUpc3k//xNJ7+SLGsMDH9mgX+c4XvdXn
A/7H2osp9k6/knQyA6p52z93o/5e39616mAxzawuVje7mO/OUsdaP1KLxKQQw0rb
kPp5bJ9HJJctAFfg0hYEydx6U55PKG1/3+GtnKGhxQC2GcfHq3HQ0qM9E7fnc+9v
xv6/b8lOEqMCEx2FixG8c+WGUwGtPl1EMOO46sNhQf4GnUjkmenOBZwd6OdhpVHe
XFanyJworroyxw440ARoKK4HOK4ZMtPRbp2v269E8ya8+ubP9rcnQk+WwtLEFVlw
7BMnHHo/5A5lRLOywm2bjw2p/zfL9q2UpdTISojO+nsPz+mfwo+vdNW2/LdjTjGG
0WIA/IGNJddvTC4+jR5SxY+cabzVPjbEr7S0xlMKSmpd+PW0jGRx8FQrRY9xFQ/8
NJf/ik9IreR//c9g1iPlGFOphqFKTlSRMohLxNCF+Xfht9QPElwMAjA0y5oHEUDh
K+QNiglbUkyeBrPYGN2ARb4CR2wVKxurUXCN66isiyKqCcnb/buVOh9aEJjaXkqk
Yt0FRBxjCS0Z5i5zZQ0cbT+OrjUXkG9Vk/THLFfK0AtcD7PnBabbrLNw/Xq9QSct
5rFoLMOYfdiTHPrLQMb3u0OsmCYZP05GgGtcVF2mwT2cm29S8uiIa2vn3dXXLADV
HnycHO8SOgiI0IDMiLd6FLMIf26d0YzXT+mqAm7vtmyYh/XfiTQU/d5waDZHJnQN
LQgdHpMdJ+1QMPsQtPej63GXWDH4vgI6iCP8uNmEHTu+UdJ8TJyJNnGIhkIvZqWl
dapLQuZFK1jYM9dQGKBzdSfOsj0fjs6MiyVpz7YVJH+piLFS7QE5XZcWjqX6Hj2f
ygOwBRXYCmlkh9L5MG36cWd0R0n331PiecGL0gERtX11zKMs/ouazW1wuT3fsjMC
y5HMiaet9mVxXMZjP1rRu01NJvrG4qqb9EozWUMWOLkEKb7pgmBYdTJuHY0VpsVN
/ikP3XROSBMue54TMvJ3qRitDFpzB297q8cH0MbODG9P0DkDCdvJsLcc1UITRHfK
jKnKO+iGVe8rpus0ghFA4kmY0voD4CZMt9MTsHUYBDhnQ/0e+zqraPaXB1YgOOHQ
GImTYX3PQKei6XJMJtZFkUD1OK0vs9l75hU5S45u+Xx92ezFjNzoENLQHtMNV/12
KLCxuJTwy+bQa0omrHWiee44V6bbuGC8GFUACYrdJrEgBbkBq97ZcJUDCrTRsyLZ
vfi9Be4OMThVoeHlRonXGPJmTXk4zFuNf3Y3dgnqiYNUs0tgyw4t+ceFsXdY9PkA
4zQci0KXB91niVPPXqovdHL9GsNKzTSScUUlOSlPScV8uOUEQplDJmljD47UNdmm
cvP0FEncnSfLPUOMffOpYrPEshYX9dnkklqk4Dupuq8TKetvL+Xh9gERowRXBwca
XarT/8hfYOlrIoRsTWvHvYhwCwde3zanFrNed8T1Id89+tgYoXbh2rOU6OXhTpPz
+H94xqreUglFisR4K1f+K4Ij2oNxbabczjWIhlYQx1w5axn5p/H1ZRXY7ryVYl1R
GfAi2GueaqEoyd2c7A/jX2pgx9ym6gME/Kdwc3L+Z7Nfak81Ng2RWmO5JgJQcEoG
e16hb/iGQMymEkKaEE9rn1RngOjcbymqTXPmbFegtf413PbuQKMJdEMUIoLwRQAd
8CLKrGaMC14BxhOJVSc6S0ugA95ttlZUNAqscLX+bL1o5FduouEk+sNE5d5woVlI
SfpgeXrI1sWXL/5fe1iVU+fqJGymLHDL2Ge1iQq6odRgjLI7yx7t2YkF+AQqhdy+
gIxpihmr7pPDO5RPgrDO7WTjpUzL5UkEJLScGTUi2bvpt2RjJxGh3UQ/42NlavaU
lxxNtXx6NIBXM6aVgWzhqwfhR9MO6yfrtNesO2xebr55a3srcSwulBezQhXYusGT
6ekkcH7egBRpJhDzTmmIBJXIen/B2Nib3i1Be2mMvXjBDKjwR+J01GPe9qdFxXZY
iVkpNq6xVYCZ7Wre26ZWTYyjXxLh6XCowPbmS/kC3BrNmwKXVfJGC8iuSRZjoFAg
2t8j0/65uDBVEHOz0ObHgeyrX0p6StBRxYnTmRt4i4z56hwZxzpFHIEzfWRmzl3V
zgE/q7N3fVqurkmDsE9sDvMSZi7pJq6CpT9v3MzP1zCUgMe1k1Gfvz801UEa+osf
l/qdIxRK1Y/0SyZhN7pXCUgYgt5mFmn6uJzHapW9jRUnDo6gQ6gZ1vZ5XgdbffGt
PEk+Q6XzFlhRADa5cNVJ2yTtpqo0kSIbSuE07NldRxPxVebhAWktszzLHsnguyz3
6mfvHK/33kE5oGGnVs8RaqwQNPeAXlN5KCNfDKHDs4YetDtHW4Os73AjiQ0Z5WmN
0GhMO2ylCHKicDXAI9HwsQ8RtEC4HgOPtVjSe/YoBMDgumu3inojfLO9/3N7W+ov
5FeRGKy1nHelWqDtCpkU+zjnKXOzehv4ohWw3SUPsgLsoK16jB0o5p2PupSiavZo
83BtL1ElIMXFN7lxF9dLAOV88VS9fxF8h3pTDhgEVYqS41OdBVrtQU6GyoCvWXXZ
T5CiD444B1G9WGlBDLyHln9E8gGG0jJ0eZ+6fEpaQBkHm1LCRFm12vawBfaZa6IG
JFDVXne5BloLbBgBy+s2DrWQa3S0cXpx50QRPaKGrhL5fr/aSMWfJvqLIYiPT16+
LrEIeAubVesSfQqlhPzKRars2CaOr3fymZOcm4/Q+b3evPAVTwmqJQWcpjsbRTKb
6vFdMJiwN8stJ/4hih18XbHJ8qMr6zeRxCtH0mIlsVnGzdh1sldxKnt/SxjdimY0
ncfEqH2W/iqP/qiDKsaBEayWU8r/EElN08wJzhsQJynGp0d7cgmozOUs8CHk9n8o
IFXUbwBHgAAT0W32UUCBkvBQ0fDzkWtl6gVW5FoMNck377iPWyTHt7rh6ueR/63T
RCCV3kqFfBsY5NXEpGNfnIwpQJpzHjteJjUzahsdDdfi1JceQ5ms8wgsVkTTzxRS
qiaq/7H6CjZCtGc+gK8vALNyHasGceQbD8lqqiF7oa8jNZwcV5Fu2LO3bgb81rii
6ApOa5aAAMl5UQFBk9AzZ4BfA2ssbGWweNxNT/gj8BD+5XM3AqaXaWUmpJezARar
adb3xbpWdUupMzeuQxbgkixDj4K64TAwBiAgdkzq9ndxZwzS+F8hk2Os23PRRGd2
qsk8Gwh1k8Hyr8x0+FsqginVbETK6OMgWwuiS6z+xF5rz7Iwaf7XlnG+0YB8T3G+
BUJ9YPEx+RkINBt4KgJHTUS+36UHsfj5zp4vzcuf7J561uczyER1qHxVrhT1yj2b
bX8k47a44vBKmceXfcps7bWzCADNypJTsYJd+tmc9nQzU3qzREtVEbPth++7v6LT
p6UpiUvN1Wg6nwOVPQH5WUvOY9/s/eltpWo0bTAkGN9j211tpKa4+0yAVPQFdruz
P1x42lvK4RxXpishpZADbppBErHwQsFtc7KkddXx7STXks+IcPjUGeYgwKj++Epo
1KDDhT4ZoMBclenBLA8EBPBROR5JXmUMub/xqnDDjKWWKA9acm8b3eEvXa2KYcY6
1pmWJU1hwM01Sk1eWHmxyfyHa5F0sW3Trt/9j7MTS2YFOeFhQcGw3tCsfzyufnO3
ZBpTiIHkva+dMc04U0LjVvVpnbFTNJhsAzBZi5PhLMt98QxucOmhCJNGfDvetSED
S6uOUq/+J63KcYqOkNDvraSV/3i4ce5Hafk2yeYMRPPufTobFA3yP2f1+xcyrVFN
KVT/EVAhNmoqDciPTo3FsF3LoH3LumUg4WpFX7XbMB1wkKNDUPyszt+c5rTSpi+7
joMynYErZQIPdiqQHyteRLGliMEmFOM/EoG/4TOb+E//oV0Dzw6yBGSjI+Apb5io
BJcvTABNVAjoD8X4KlxGveO3RWv83RFGACuzSl+w1NjLpfxFIdtsaaTCN/ai9e7K
7O1WgnP5MPI1eXVb1+YVImZueIELv8JxE0MCHQJddlehBFLT5rTTk5fOYH1/u5GC
zTOc1z70lHsbLPspLR5Fe/F64HhvShEEGYbAMCARNKz0vUU5wkhvk0MEcNXJH3iN
TlWR3Y169jcWSHekT/YLtRcrMtegEwzCRsQtn7w40Pmb86EekR3R+ya050Yp1RQr
xH/HUQqLU34Ey93R6awNbZygH23Az3rhakdN0NJ3qTJZBFFx9xrWrA44Ca7EVwLI
OtqEfi2cLWBAtozEhv27YnkeRBbN1G/OPLC1vo2k7zkNrlj2oL9y9YMTa1P0Dkx1
wxrrUzTqsgWFMMO8RvqwTkM/7a58xctb1snWqPuUNHwWGlKxg5dk5Np97XcFGiSI
F0Oy4NtppIQOgmUophRmHBASa8ZpXECNlbAiQkpdk89Tub1AzldzpkKSBWnS3Ew6
SKROG84A3GQdqCwcV274+RuWr6KEBWjvXjKMjgqFhX0UKz1y9uAXkpq/dX+ZegnY
WRlyi2/6KRB4GstBJZpxbOH291RppQt43b/pr3XxA6K23SHsZL3YBvx+XAh2+vF5
oESyBHcqngIa84rSsrUbGbQZQtXHc4DK2sllGYYDIOgoLGeAlCxQpeFDNl/sIgMa
qbCEgVma9+B4dhkXXItMg2WFKk84R+E5wv0GUvMbuDf2HfKFQOgLVzTVfGTpGqvc
A+ZwS68g/J0/giYT4slJQ01ihdcHlJo51eQ4K8jbXT2EEnd3MUtA/VGEQfu0H9qN
39hXgcyMm58CLACR1ZEAcEnLpf4C/5u382nY5WNYVWenUlkclxyZZXbrbqemfBn4
FU7m+b5Bqrm7TwjD3fvrDCO6B3mSHpa41qQueiFjuJORbg6beglyBR4ejAugr82C
T0cOdmLRCwjjHKQO1a9JSeTArxmsIcHNhVafpT04tbbdrRYL3DG2yO1kh8PJutvx
iSpVOlKauw+gt0CFA86JHxBDTD2gyY1TSaonNdnn0haDts+bPy3gF/MbiFBq5+BH
CeOrJjnFaHRieTij9s6B16FNP9gGkRxPeEFskwgwMFilb+dgVPSdcGaWnBQYFu30
VMeKSOiV8Man8MZyhr12QvPRoKWFRQE0+X1ZcGrDlK0fhKoDJ/HNJq9Je8R4sQ41
UvXIDBKJYiThteJduqlqwln8wTcU0YP7gmKc1Q3MTZAAEyf3nUSag9/Ck1rPSzS6
j6dQaGi7ez85i3kWfK+abMwthVqlxN1ckGtl2/gxQlJ5AgmjgrxUmNcxuzjHv1XD
P3LwkZBmlFah7n2CVphvNguAHLvP6v3qztRNFYZR3Wz6+2ChS2OgmHoG+QL0pQf9
E6lB+/0L3iG5xlAF9Dk4+sm9UNWS5HpvgHM0FZxNNLhn3LE462lDVOFjBP09s63X
B2xdaC3WGmxJotq8OFMDq1dffziEXQevg/3sPikPchmn50/ywSSl22ffGsluMBZ0
jxWVuyu0Fkk3yYCqoWvrEBMuIg17bLN2evt7+cUkoN8T6xdT7XoWOr+Bd4qsCNys
J5m9K6cs/SdUZfEEg0psuigmtu3hkTzdZJpC6+MNnv6xNZtgU5Nc75wINrhFwCbd
TdZvqBwkV6giU1emt/AT4HF6Dgu4KkVuNA90ChhSn3UliydFyw/gARKytiTSTI5F
aX3q1fNA3TFEw8tbqSOMh1QebRnseTsi65IV2OoJzhH9nphrc3GrAvfGZA/K0Gy0
qAH7Th1T/JKesqskJgk898KXj5d1aGXblBWX1VoMHVGWgt1bhb3nAv3sg3gRIdBM
+ffQ1th9SACEjBaLUCaJNrURMl+94U/+4PpVPSO6E9hyLFAdKipqQ8/243s1BEqz
VlOPiCdYB97vUyF4jooXkJ6KnzPrAn3+kkZqRTAR0Uvq7IpWiWL1yLBfCseQ+Lva
EVVMnhj7cWp2BWEpHej7ApqMgkrahjdoN3IEh+XsfckHA8FSwESCWHLnq7YZZJ6Y
VsCj2NPiCMZBBd4ySyiGRY7YAoWU6kqNnS/uUq7dCfQwRoYkX1WXhznIfaqHo7ge
++kTJhgHnM4EaAKswE4k+T61VUJRFBkNeLzv2zhuylzOkVj6u4iZZHppFxwo9XQi
1AOY4rhqT1JZGld99BJDNoCz4Gu1RdJ5VbW+V7J977J6n38gc8F3cOhzHBEApesY
jSu9bA3HrrXi0byirW7gsxeT0Bzbci01PwLZ/wKhMXFsgAJmO4THO+ajr14t6XNB
nZM1oo5YvkqD9yNxdnHwpO7S9hEqLLOgfX66qFQkySfcRf2A+8rSjvC2fecmn+uT
b95EvCZ0cLG9pFpVM2sxkOwFxaM7bJVPbxL2UeqWdz0L1hswe0wJ1+ir1XFbUCeN
hKMk7QDydZAFSBy+b4SeoHMrhbLdfDBYzsPtxLLbHf9o6Enqxkj41PdmsBmS8z+/
i1kNJ+llUru80vTXwobp6rE+mbDCkzmdKieODOa81WAVW4WrSPJFwrOrGp0sqeox
RsDL8u7AN2rAe9tMf2snQZM74XjPxYjsJHHYi4cwyqgchQdzTQoFXiOEAhtiqUkI
Aad/KLJxwogI14ElPjYOl1QZZS6h4VPZXtR0wCtBR2Rmd+DFlZh3OOvpLzGj0m9m
OzUKTVaCuykky6Dc++M7Ojzcsr6tzsjYdz4BYD/gojiX0faWVOBiVdZuuq+OIOQ7
Dec4XhixiG6Qn6Oh+7BqI306H5t+eomdpMJipRI9zUUt8XJU4NuG+VGliLdsofiO
72zk3C8NKp6QAWbpJrr23Y7PmbDMOtUW00Wygvpgt//neF6wzPyYvP2tK+MBIRfT
jyraGTw2IHUjgSvYruPQwa5S4OKjux7JsqJ6yQHXV0+Pk+8DAHhStG/7cVfYAIpZ
c7t/XjWwccWV0DMDNozLzIkG+ErAruZP8RhcTaQpabYgKvFfp0HuCODFCGhdVwhu
lHm0eA2cbozledXrzXxhsYEEHthPh+9/U2e71Jg8vnNy53xumfFbSl6VlpIeaRLz
vugxPk3atp3JpKNAs7bKF3+/ZM+/rTgYzLZm/uYjVNiG32gZU6jpY87PQ8GOnVuZ
5IPGkLzchh0e5Q2pRp+nBi5oHL5D2hdic3UgvH3DLO8/fIqHhuHLa5EptK5n05y2
S/Hv92ZMVukoMIfJ56vqGx7Og4d0R42TMBkaLcsnOGXVLVKco9aAPzFDl/MbqaPJ
AQRvLVAj5lyrg3jZqoqd9nSKZfoYfeuEreIiQCKPxdkDlMfnYBjUMm20Y7xOi39M
KJaVUzz+Zcvn5QDAy9QwYMNaJDz3MU2xscgcmtMAy88vm+6OTClTimtfncn5RejC
y2/xAK+h5SBuUI02VAkMkwDANoXcJtDwwuA+R18Tgz5tRLyBsH1VeKg1zc+mmw4H
ak1+4j/P5lYzvO4CY4Iuq1qXgH7fX4WUdq58aEhpO2FX2QrH5+6bCSD6A6ddmbrA
TG9StIThj6ukOsFrkAGPz68bfFYmzMrlBi2U3DGPsCeF584H+LbD3q3BbTGQ80y/
KnYXx8AsMcvlG2eWYeIZ0gqSo/fFh0aN+oqod5rZlP4yk9WK3pUPZ3hNBnpkyR6F
EopzNXRUOPEMCXjdnjt8ihjthTmgQMmhrLM1jwlGdxL44V2YIZ5SdoMQ2jXn2EAR
UOZ1RtqKAqCsZCZZI7bpcD/SRxe6xn2vkhhtsjW7vkjoooBZlaHGXs7gG7JRczce
j2hkGGPti39EBzw92/pNC0amF9vbib8WEZzc2ZRhbT4xSvnloHLWLagTUUaJKwqN
ho/gXszH9k4pMO0sb9C/AQk4+xWJU43XtCOnuxkR/NX5Xq1fbqwmnt2VUd13xJI6
crc1ORWDKu64Y8K7pfXNrc+7Bc/wabJ+RPueR0+ARiBh+3RkoUSwZWOpElBfp31L
a8RV2mVYLMx0X+huwrVEEDKQ5HXBQ41yoME7Sqr7j/wjIHflQ8/+VOEJhryKQY4B
gX7PooKiVvF5TvRX5GLdPy+HFGn76p2oFjFcuX0hmVqm8LL8Dn8PuEoTGe8+BqYo
/O67JbkrXoDdw3JmeMziqGOpz80EIShJn5G1k1SBo/UBHzfEnBUei2Q8H27mx+XQ
H1vyQ+8PMRXrtJFkISdV9ooZKBRqmTBpwlfqk12c0JxAtu518z2e5vfpDDKxWMcp
Oc/8hu/bXlHjesiEYkxkYhv6W7xm4W4ItfLZzv4oTdn28HhD3S1Fc8bLA4B7Ht2e
xWbgiUuMh+m7bqwbHDTZPKzgC0vVHjKf9N+IW/2GfBgXrR6kVdaFYKnrQgx+h3zn
wG0RHgrwqSSU6/oaHnWZGxHsY7By0nZHs6GCUjOPVY6EzDJy19jafRaG5QD/GeuQ
aE7f+voyRljfz9NQ2cbNpn/2ZxiUf/4DNZWEiSbT48fBQ1VreWJNfa6J21LxeuDk
Z6t6Kj7FRtW388icjlahPmAO2wElvEMDOzbY6fhW0T1y9qpY7qpo5HhEsrNpkB0v
xioyEvDkJCv3De8rHvODVjaGkQJs1mwjqytZxgb1L9IYCpxE8VMJ1mvCLcBAV1BO
gRB4wC2z9URHb8V4ks4WzoLLelR58drZEJm/Pm0A1U7v+D5Y/OCygkMug75F+6eY
h/4xsgWO5hFWjtzLTzXo+11pADJO6hLwxne6UUlj2tusKug+laPlShGNSP9JciG1
zjZshWLsBRtZtuFbAXYQuwCaTVCzuARb0aP14eXjLxspxvrpdjUqzdvH/bCiZpPl
z5nBd4FMvQsSoNIdRs0LdeL7J0/mleXdKuSVMW1UnjwRxCgzw1Gx9LoXG0lFWmV4
bCzGQp3gug0KXmjSBA9G8GJUC4GslenC5q6tt8PByqXRlPyqzlrj34yBNuHCAXmv
3zAMTpknTBT+cK8jymfC2CWNeQpg8xqg1ToVw0LOe9RIdJy7YzCrfdbNYjhDSSis
0TGWqNObRGDpoZ1h+AVy4cblPQPOCbWmfJ4xTSOoGn29bxr06RZoT4lWT6HYFFD7
BZvYTh/vYRJsZ39DMDDziXH4ER62URydTK5ajNiyW+uQRuzmVliUwegoFGu2SZiF
ZkxVPoMUQoltcnT2iROkZCY+886/b0n4RPkBiOXRA+nFpsxqUfiDcCGBkJIqEgT5
jc9bY0KkIaPPPu+7/2YF4Nqy0+E0ZFRYeXytom/sAoqQCKWFB87IlzCySA+4Nme3
lyoE3W4dcdIkWAR9Q4nmY0VQefRAQX8WDCFZbEo3jIQyOZwGM7JafTFXt/BjgMiJ
GurwbGqI2LcUtF7eM9Vllqb5M2k9LVka3wsYPq4t7e7NIbriex2F1UuPWT/Kyj7Y
1owl3waf4t5GkJekPRDK7nSDD3KLaiyeifR5zroJUKdBOV3JCjqXgvA3/GUgZXZt
fPDCqOStQoCoTGHimEjB3mMOZ3vybVW+tZ5xNcKcZrijHHEohJ5FkVFbc14WENEX
fQ1PphEKFOONMcjDUIlTsoRGKMeO+p0yuzo/Ht9hXP2+wNoetos2EUzEoPSFd3mr
LNakAlsFOyDGdwXVLPbXDAfFGe/0NLs5TcqFMsiesGSpi28lKBrNnuJJdwPdJZV8
S7ExUwdcwOu5XSRIRKcDvUtmMv3ofQV/AC8C1Zt6Fk6VLv4t6Pq1pUQgJZRDO7H1
5osNnFTLN0s5IhR36on4AlcK7OogfNoYtbQa7cKB+9+4w5A1Z9nCob36uYKLrJwQ
n3+RF9Xh3Vq+7MtGvw4E4bnWmpabrkwywVfs9LDwDy5ZnefSiqz+VXLyR+okCAqW
SWkhbYD4UHtBRdeCqX8AuNtpXngXLMbSmNO/5Yo4aNFon08If1uZly4oZ1D++ebz
oIM4LK04fjojSmhNY4N8nrvlc+za5NkbzkURBqVkthywp1pyQ4kvBZXgRhleKryZ
8QzbuAo3gNnVKBVLoWxGlMBdegJnY7/LNMRUgOQSQ5+1yQG8vgbhUbCs69MvrdQ/
o/Mht9RypFcDivrpQOszvMeMFsxRDyaGrG7BuWuIws2tdXziz0YOh/tjYvRik0Q/
r7vPB21YfD15Oh9+V/MGeQ1z8ZXJkhwyT/h6W9GQAYaeDVOc3cecEsJmRVyxSokF
YIwjyJjxzf9+HUMkGXL8R4+py9D9hOIm3SWowkROt9tfED9AYnV1NCjfc3IlqRpE
8SAXlE5afsRJBvxygun1BwJpt8NNaSEhHjuVtlXTWq8kxly3eoJm7X8XgUMCeNRn
puXwb/S1p13aSce/uKSFI99rbdM2//YKwA2DS/uHel9o/A6v1xhm/joTvWsvzRVb
yt8DMgAFTQv+zsXnFnLIDRhV1gd/d+bzkwxH4ZxQk2sS80W+1YEfnbTNer9FqQ1s
qB4L+fVkYOjccQLDyJR9VzmRQLb4n1GrtM6WQrLJ9RfPTv+fHhKTgUfs++H2TTUT
dNVC5Tst6tvAgp0WiuLtK+sYnIT0uIAG7DvaeAaCjlf6F5w0Yf+DSRi5YilzInjb
T8INwHNMJUOzp/qO25W7V2GlLYoICB/t3E/YtH6NIDA0IibGeMY99ICK/h3Ea8w/
GNybdKkjJV4PjVRA65J+jfv6nlKeh5sdN5XvJhC5Yi9zNFRyt9djkKOLwdSXAxJH
gBkQ/b+dFdJiPmEFPiNF8KyTMJRAz16c2qrCdNXvBpHek7qkTh5prarkt+mGbQcs
1I1USB5gqblTtdtlh9gsl8Kg4U+v5aYzCF8bZznaZWtJW0JRhcnruv8VtOhrtHBB
hgATkAVbnbtiIJl1e2xQ6AO+uJ/kZ07ZdurKW8VX/8RifpBCkTGKh3qwm7+rUUyv
T0Gsf3/nfMpQYOrLYLtqU92DCkm67hcAMYZ3zHVzeNVyMzSkF/qLHPQQ3yvE22aH
ftVmlJ6FK3kTyqI8fBBa93m9x9CGz4C9qkQqnY2cHltyBP+uJ8dtoiI12o7c/qlV
lWrOBm9+GBBGH/5VcV1m6Wy3UKOdTesh26MDED3RtUkr3vcTDo79p/c5ALNFEjnK
IVyWNl0jeiPspiZYLeJyencZ/wfV7tyWtKfCKC5ZFdAz7TbHv2HxXzTZoz3Hd/Ws
24q7uaXpocEE/10ibocaIVBp8LJ/lGM5db+aiDmZo0duuZF15k6ZayCD6f1XhDk+
6AVCN/b9U14jrcT9aIIqr6kO5+oWXeepJ7fJ7PXz/uM0AvBHJiqLrW/zw3Tcx26c
JNSpZsOoOCi/LLTOcyea8UWy/SD8vh2R1SboeIPwBT+m3bY8zf6XJy9JS197e1dP
l8+9sUxYS0TkWsKwvcto98Qrg//S8pbIiXcq0uU8aVS+1SAi7Sz459eiO7kS6vNe
CgtJFDkEhsUMPIAide04wtTFnKQZiqCZKfc0wGNCrOlNAj6jYHKXJkEpsr9kGMsN
sUqFS7ZTLFvzkxe41ztWDRAKAqngzr9Rj+R7pmGTns7ajXSQJqoKcs3Oc54CN1hA
hmOY+GZbRw/dGx3Ytl2P9yoH7f8njNvDl5oONiC5zxv9vFy4jIShGkMJBxd1cWry
GNbBgCupptXUfNxgHBnAbFPjpzWzZemXuh+RvdoVpXaJsNeCoYqpv8qeSK3ZNQsO
kwE/jbvJwV+xbfpHqS5i22ghKAARTsBcTkN0YdBCoXQj0lGc32uQ/99oxZu+GD0c
CuP9oTBwUizFj63ZTQV09z0szcR+9dkNo0Ce3bJHwL4D+P7uVqD+ugSTiNYx2rSB
A0LbWrktlMqhq4D0hPUp1DyXMvBsp8n9nAx0vTNSXMt0sHU4LlHfU3KtyP8zlLYf
4fsGUE1aacYyhNoROHXp1PVJSKu+cJOjzQQC4oNnQqH9JsSnEL5ZldK7Ky57csQ8
fmGQc9eqDCFCKIGJxu1XTL09ODl4j4ue2IIqNijvk5WdPvT5WAbKTUy0tT7FHMKZ
zxVlwwzh5BHyd3qYxnXlWXodiPK43XKE8ZE0OHKOLZGUsPEUBN8qjBVzdbZdw+Us
uSuIocGbwpjKn3vVJWxZfZx3vnUXDqd5jkKD6dr5e2x85wfQ4lT0pvs8x4z+dNZe
0BXnvtldxlsWOwNqdfw153W0zDt3Gp+M5B4E3XvzR0Gh+DBGGPBGUvywIWV1EVuK
8FymhAWaZkKCaxRxnn9sji6nvGyCXz71HhUQ+i859i59k6VMJ2yzzFILP51hiSvX
RSwFJlAcOhWoej/hpWivYtskaRlpmEvvK0/E2qXAROYf/eyFe2Xx6PmQGp7hmKtm
t8U0pUAK3d/5hW5hxLuRu9atqnrPcySD+nqhrrh+2+oakEJJp0+4lNUefn8ICCPu
DaVEFmEUjaS8Um+RQ3rM26bs0NLGB2UuV537NqPlDvMR/uNoGyBgPCC1J4GIBpIw
esor4GVbOr7+j73eg1gmpLenUvYm+xNzavcjR90/nLi32kfDYJN+UdyaY3nh76mW
2Rkwh/vS6RUGgZVnQPhYiTzfAi8KK7EEfBOu8FB243NeuKM3FBrKs5jtcndEgVpg
XnONN70VWasC8P2UPooiY73lW4+Nq2BfOGW/1C5tm69MXfSWJh0xkxGE6NzAynGj
a5IKr2m/GpAXIiP8ytxF6afJRxAz4UrQHIBpW+NpMEyUhVL08mYc7vM4yE0Jn/H/
6L5ii7DBpTsAYXCQfmEnaJRjtS6FUZzo7Wf6K+vo4GharJexRC/I+J6UVz8Xa9MP
96L+b+vuWoqWoPj79cdFFmJB2H2Osxstq9N4qZqTKF1Am9E+B5kZ9Xu9RDWmBDHV
j+Sn/VTX3Do+uXBljIK+X8QbubOKfD3iEf7NKkUM1BI2YcKRip/R/o6tN4rqSkTs
ItG0fCllcSIggtaFVcb8Uh93/c4vjw57Tb71qESFkhxXwJopuvYzCfuJL7vBjUEb
qEJNuGVBtKcw/o2V2Ndk99eIaypcqEgBmTLMLQMDhfMV4wgRYOV+js8912AN9+ag
RbFRz3JxtZUwdwuDpGme+4JDqCIJ5bGHjv6VTsDdozWhJksnACuYcffKkFLvB014
3d6WT4NXcnFAq3EUkhjhnIgpyOvsSNA/tUwPNofBHWRFLeFc8rwLpVOw/KWoPUDq
q7CEsbY9FKB8fuNqXxt5Z5VW2/9Ru7dFkdmoihV/tDdGoY+vDTXZPzzQ7WVKPVMs
uT/FNlYY3vaGtuzF+K4OpVWqg88vzc4SoFy5KX4BG5HFAEYyar3a7eoEk/zIbddx
k4I59bosdxm+BMXKYjPN4Iq1fiV7jr+imAhDxIcpris5dlWWUj7GKfvJuUeEp3y4
oOWk/4bv1gBUpycoKrvHIIkvqH0WCb1rh6gfhofR+B2mSsq6lzMarC0mMEqj3jsl
PTD3zU7juaJ2kmt0W8FDxtUUPP/DVQMyvbL9gSyAzRB46lXCZBbmx4832v1c0vjj
tbG6R+O1UA0TC9Ix+bRGyrFN5FTcKVkvACD3Lx4oMOP7l0C3EjlSVAazt8ln9JXH
2prb2PrPmAZv0H5kzJZTapQAdsT7t+DynVFko7UDw2c33NChTNN7mvOdRdFSFcv2
TNMbCDku0qv/KeQ0WFKYFpQQ/ml59RVYIonZA+16mh3npLoDa7Yvgs6OX+ElwUoc
RvnZdAUpa8AUWVEGJbU5y1alu3vJj+/C9Y0kemgMWBNfNo/3wvs+b23EyvlalpgO
HAagD9hlR811lI2Dgwj8HJnZv6hDHTL0ylUhFTJ54czpzdfGrHt9P5eIyCqypSqK
26xfdOzoDrXu2oFdmgUzF+R8BPC+Yw61DGwjH//IXjmJCGsSZH+fadzRLEVbouwQ
vKBX7ZIUucZj8Xd0GTExfJCbM/Zo2Ojaj5m8/kvqBX3W1FjTQyGPMvOR3bCrv1Xy
Lw50G+6bnfR9c+4YlZPVCCblx5MsW7Igj9HnGif/vKlINpxMjd5HfCwDmzCZwcJL
cHmntD8/LRaOMRS9SSGUZhBaymIZiMNxK07T51SJQXNLfOt4nMWeArsI+3TWqe3r
SwkLa4BXYKz2kCp2U/oOIiB6RN1nlcTM42TiDXc8I3oB+XzmjqmOwCCv4ZNr9F87
lbqY+LA+DcvoEmcu5TIk56L9bvGD94rw79qshRFmY6QNp/7+wvQN4I7Aw1SPhzjF
M0hUQ1h2ZpSP/5F8xEEWRE0iwz+BjgrL5h+gPU2QKH7JBetEuX9fqYgzlgUCrXK2
fkk2g2SrA7Ceh5ztKmmezpMZxrAJnGaZzp8t8VizGGWE4OWRV7BxFG7F/8nXKICo
dm15CGVMaSIS4Q5nBHQd5XUBPVfbMzw8Dw3qU+S0fBOyDxELx+yC0doqYY3oLUxN
2B0nH1bspSsaJFuC7BpP4NY6KI2eG+Fcw3WovrhG0bOfQN/CnggrxeT4YwZlengu
HTKaLiI+XZ7TJtoE6WHpo41lDrH9zj7gR8N7fhqP0QtXVa7NCMKG6wJ14YHcPEHo
poAuWX9GtnXlIgVH2n7NdFDeQ8zmshxEIQsfJxhS7vCWh9xqJLr6lgS+sGHlrjeJ
EF+NCnqOa3CgFXZ07QnEWPEmHWzitPAj8xuyPwQXXfaeMWNmaYdC9cQ71Qs5tzxn
gSXQTkgQG8kaw7A8Hwo8fwJzELk4aZUlCpBfJgWwap6g1KXTbJAERX1UrrxCJP41
+n38ICzQWAsLu5DcKmW9ytTShY1L9BPUk8WHG80gL265R5mbxjAj8R+HB8cOFjE3
1WxURDdVOXYBMMxmR3enMQ010Evj6Mr2iQeSt0rnxeNVwSACSQ7xHf46ytzal41Z
VK1dkY39/fbIiLse7DBm2+QJdhsc4nr1Is3Zh2bRLfNA8fxJAtB3c7F/uvqXGDh1
3MqgxKRZNFBh8cFHe/Ilc0QVgSZa6jZzdR6VFYB2XuQY6NKOnQ00IN7Cp6sCen8Z
9kGKgc1KU8XUqGD+AlFfuIdziqKv+HKYdnhtu6zdwjrGcALjVdjjj6Wo0RFMdfCD
LefhO/AX91IN5//FAqUAn6v5YOswmtHLThwYfMF0kl+ZSD7HxAmq24ZCEg3zEYFj
9xeSxm/H2vsorz95nT3dLXmyM4tGMVsw26oDaOY1gCQdmgAXAbiMFlOS5knzDvkg
09WT92vUBmHcmAuBQhjzCsfc3eBG/XP4SIFQthBWcxy8lXOXIgDy0j1TmGBlZ4Yx
sAfc0LSVxMVfmEnDmiQmIQHIYzp1SJpZatkbnO6Nc+VAfgDebT5CJIcnnNrZDrb9
Iyxz6ddfU+H4WtJ4N2Hz2FoLIsD2ipHWrtZwRZC1hySQnRfmQlMMkg3a9Y6733NP
fdWDqH0dWSyam0NkYkGSaR4khQt5YjkgCbDWP250M46aaN51ARCTigBGqjxqgWt0
LBsAQgFHoPKC4J3TqQVXVtLn81SP8xbhXB22KP242FdrJAcpKy24R06eIL9NnqeD
fjW8Vw+KpJuZLvpmUWWtGutOmWcpQ23Vgve7G3Egrr/K/KHFmrr0AVkK4nK9fDFI
MAUUopu9kq7Y4veNvl5bpuzR9NXzkYIfhO6YdwH/213YsBFMpugEABjc5SRW1qWE
Hu1IAFBfzyVqdcGFchMCa87U8u6BUQ264CXCHqC38aPLLB2TSRQvAQpgRq1xGlyU
MxEC5DB0w8h7kLHYWH2XNs/mNPmbUiV5FdUrAG0lTjZmpGoxDuak5cGWQCcWy0uM
Ct/WXze2ddVYM4TbIJEU8VGfJ+Kb6kDgqL/GQKlcW4rbHggASKSaJCKwVpy8DAXM
P6bSNTPhj7VolBE87Ry2b4UkJoqz/v5FpCayAbvbcaq8ku2XMqjaOGACY0vcfHH9
ZNIpAot4Qf9/Dgh57pHPcBI2iYAjRfidWa6Tkqxg9dc/F3WKtDBUfONmz8xrTZcT
DM8QTQFAgg6kMrR5/hntGGsYgUaLD70U/moAD8P6XEWucxLSajh5B+4UywQTQrUw
7fRRw6NAA9Ot74XpjgtO2xboKshmpJRE0Ti34gLYxtfHVLUVhl7zTSXPUGmG6v7Y
fiXWv88pEocwYjlesjmDJxEPb3vIsQI4IgWSHZ67/5li6gc+fHVM+zWFfRdtx+RQ
6Z+hq4KUTJpjTm74o3pHWWQsGDXFdvJZsap5vXmAwwL5k3WmQsW/Q1kWjfVvJ8QW
rtZYdHuXxlbgMY8mk6a9fCCxiEGzdBb8y+OS6uZ127DcLSaicUyGAw0XvK8fJFCG
95T5ley9BlMYBuWwHIswpsNIMG7cz2e8Fhxw0Fta4kFRMr6F78L1KquF5oBWQayU
A8m4u4Y92bMOh9y979WbeZJ/Go8Eb3+pNTwgnEIm7kceaobU+duBzmS9LEcXB0wD
dTxC9cBPNQ3L/DMu3DGrxCQ4hzmvnVgi4YFY//dGCNE+/qXTKihmC3+7MJsTbuRo
3JlghGsJdJC6+ZOJ6Lp11TZ0TuwbS8BE4jWLHYY2ipO+bdRI+hbhDCVTY+URQV3H
w+KXBasVcM5ZTvSmA30K7b0GDbrLMhhVeh8O1czlaFvnDHoX2+t420Y8lVwLRAyF
M/G3WhZ5uOb5DeLYQOPnJNweKvsxjdd93TapAfaLbm/yTeai0x7M/lZ03ACJI1IU
ymDY3gq0/Et/bYZoAooXLrR+Y1uDsarHMyRa7W9G962IJjz5UczXmG5j9JqLuFXq
cI8a63k/Uuvfx2mO2ex/uF4bIRri/Rxp0k5d5zn7o5eWMBTRlBtjIsoSiJK37AaJ
YpFzk+rVyHVG4M1L0M6GmtwREjbrupm+aAVfSj3c53THR28nZkcIVEOmCm7EJ2Ph
ea53t2pFQkmSt4uKkObPpurnGsPItcJJc1ux3ci85TWtywRLk9ZPF7b7i5Qeqfpf
wCF37f3y0oj/auUQcn1jCZ2Yl2Pb6Rp5yIPG8eIgHmKiHNvkURT+lwkiv6EjyElP
v8ZZ4Qadjp+qzmRl/KmUCwqDHu9fKv561KYuUF8tl623+bfBPa10T/dF3Kcw7vtG
Bg4GixJR4/5t+dyn0C2cfVsVDM/Kw1GbT29XQSdQW3rraicuPUYG2+JX8kfRQ8qY
RMLLizk/sY7mqnMNtrcgpwSMitI+j4Jh1khJETld2aZdU0pvlf8eKX9NxMhxsFyk
bo4nFG0d3zm5p4wJQgEq9hF3U4e49uvO4Tfd0LysocWQgn5av/Jjj1vnUXdUVrd5
Ulp0O71AJ6udWWYa+Wk7YSC2wcv99Q6g8ZJ6iL8hNyxkV+UPzOTClw3kQbqPccG0
hnURpHK9omwtPse5LatPwAGP4eJilLLP1oFy1Fv3FHP+FgHsAGsM5XBBMPBqB0xi
K7iH3Lj5DfKMvG2rM/8qiKdADJ+76tbADKHP2RZOvj94BS2bBGD7Rn0qiwM0U+xh
OOs6P0LHiwRkzrycn+whUxd2XJlppaEnOWZxHq6f9bsHhuYxqx7TILxpwVqisQwH
Nsoswhre1qvN+UUeerHWz0gYffZraa5hy+muO3eHtAhWI0BpSmdN5eDVnWnWGObx
H7eC6Jj0972JP+QYalo//jzN1FAz5aG2Nyeao9eHgeBw10MKSW+ik+6qpHuqRcGA
5LiF1j3XHs1bKccIMFRuMsqp/8h7R+ZPkURNwxBj6qnVyw7xzKK5JlLU4dvW2l1f
yoxN6Xl0eoqVlMbQE51kUbOcOV7x2I2wXpIo4VdyVmkju+G9s/7XjSzpkbfl7ieQ
gmvXQH0CCRqe53Exe/ix+AqWB06TeTjgwSb2+hIGHS8UsxLT7nLSKVuE85SnVeoQ
eSiK6F1JMOIAq4Z+CxNeLJZMvaBoKLj/iYMHxBNVqPDFQziqutTGbaXR8kkjBx7J
B0cYyfMVsHPeF7qOf/CZaZ8A+mKavn7w/224Y/S+2zLfxb/N26GQkLx704v7U+oO
DD0WYcOkiLOWGmWu7254vmiyF42ih6/awO5IFMp+yzQPzZcUW/L7CbVIYuSxaUJB
I04V0gWe4mjwAAfGo7tiQkcjtik74vUCf7TfD8fAxmTp2LyKxFAUcjEFAXOtdW2U
k9XSKmG7Ma70SAZeBsL/RP14RBNzfFDgx+55822OnC5CLlA9nW2DYJaWTGKBdGfJ
SXE6ERtqz8xsNzTU3gu1f9ZDGDWPGUiCzrxxlHigT5slkqpr54jX2VqBPEmh534/
mLn6LY2SkEWVsJx338cX7GXeoQrfNifXnJCl/Z6XvlSjJqx5Fh0jhk/GEJ5U9awv
lwFxHyEb1d6T9WTT8FoChw38ZrPh39rQGl03Jlcw/ZnPsM3FnRTWgTMhokCedf8v
5Mef9CJ9GWhLMSFN2QCAui/y/q4dHeRPLd67eVX5KUZd3duiuKWLN0l6CRGXo9tf
oFoOOuFEd74ozwjMPsghgd13EygbhUnB+cq17oqasSsGmgzOHFOF6iZDJBJib/Od
YaMWgGSKYTtYF3HUEd4CosF/leZyVrwejaFVFHF2wTO4jfby2JIXyAXKSz8qkRs9
WSvpg5oIAug6m53zXCsxRFKkFmVxioqngZanbB9IS7C6KGcCAWz3O/nz7+4FU0c9
NjUwzdDX1bZPV+AnKn/DLLWuZHTGmFVHmYKaK7lpAWCFYWqTM9Zuff1nOfD/PtMs
6EXidRUXaNo1+CFwCIMTcZBO4t4SVOb/3RMOlE6ym8+PSlUSX/PsLaHRDfS/but2
mesKanXYD2wVOEW/fc8pROblmk9RDylA9sGq4QfNyqmLomrzOkjuXdiX1hztDvFC
coYNtbL7D3U78vK3TJJp5aCGeK5FTWiPRHGyUbluks17xX+4rpkX00Sk5tYJasM1
kntOAKcKcpFP80KkYr3sftVoa+SxtgFRivsGHAZyHGDm/Iid8BiCwmsUo60ZqveE
r2yUxBCGZj1CwRy2tf7wO0fBVTLgGI6A6r/NLQvAZWWdfhmVZbFqJQiDq/a5q+jr
m39cbYx+QbRHqNq8reQC4bVDQ/8i25ojns94Hfe7GURp73Jd0HHBmp4g707rGAl3
gM8tLLkpbw/7EevX6iuT8DlKQBWWUKQI6Kzne3qBAgHyOuMFP4Z2iQQLNHbnZSGC
YLWeLBbIs8NtFT+oahodoSPUQ5/X8Q+cyKh19KaDcspTuDal1uXoha5+c6DU2CaB
ZRTEBg1hsp3/L0OEpZg4uqRKv5XHcwjmsHKanQoRkkzGCOExIe+DKNyHryXq4J8i
brVHfIAb7y3q6VODjUc/b9ymBCuGZE8QwaLr26APE1zSxRHPF8HXs7x3bwrKRN1k
JDx8uPMtWScClxU0GfjfgF+otZ+7H2ZbNGxGu0YVxijAcJ4fT2TSzrVol3X6FTTF
VmG6UfVkYO775nP2hOLMjXggeBdpmAvxlv9Ie1XIIpBpbdtkUCErib59bhuknKFu
XOZjiAHaTR3URdRiQt1PSr4XbqhY2FObws5U0mJQweyVFDRhs6mLXn8Ch7OL5PTT
9a6zRSy1W00uJxPUthz5N0zALWj0sOJsnuqlIvqUChNpAIAaMd4CNNAxToJ4D2yJ
3QVlPLrnCkrI3btxtsJH2I4zfaOqzx+n6J7xrECa6vsUXQdbj1r8NmX6xUWSuUuS
9lFsO+RZKhg6INyWvUU6ptZABQZXPpLm+Tpbmzea/bjkn1nRdfiI4K1DoAVqGXxH
3OiDaO7LMhOOSsbO11eW44NQTHsZno3HCI2OBVbsLYxt1M8yzoHKr2EYiSlTM1V+
uikRGPGLze24iADA2as43sQ0AD2YSRDoFdqyzF7CJlCQPo7pMQH94tI/FSVGkcQe
d2gj8Iv8qwwzXLpdjUu0v9W7DonbKHPmjM6fSuimKmbJdpPkRy1hmy31bG813Fbz
mfguySLX2pbIfSu/Fq9SAUQYdpVY2Xstj3uT+djJXNDUvpFO2AIRh88hMEqsjFsY
TeEzX1WEYNBw9ZT6WC1DRlrmcIZ9DaPQfOJkzbrpXUwMzmf+8pYlPGmFqGuJyzH4
mZTKZVRcOkU4R28SqP0V6datHodSZ/J8w8yvvADrtg0skOgPBLeIQ6psmYmv41uX
RFYwjIbE8q4tMxiPc8k02a53Pdqe5ULHJTYcJtyjmxBGYqjBa16AXJ6N6t8Id/1t
QeyN8uXBlcTJODvQxiONn/wUkd+teAEebogFSwgzL3GH6AXz6qXdxPzkl4pnBUdY
vilGZss80wuDyPma4aQ++IbIOa0ruIu0HI3iXwIDkFu1J2wiqEMkvZ+Pz8R7+wm7
QYBzkzTgdqyXU4ufLpZmfrL5QKUvwC/sQTt55GokUppmwjuKklfZpf8q0xXtBhqD
dGyC7sGUM/Zo4AUxlwwjMTaIwLmQtR01cJAZsMCMJRWSovd9OXq17T3QQFh9kWqp
9HNGXoE4pd+19+ujX4TABPkTTs3RpmnIwYPFO5d89Z75J+vzzl/JOfuL0SKtzNdu
5+UqMIS2Pa5GEozw+SMtQyyigNyAwv47Tv+86TJWSU6q7q/Tj0GnTkprz4RYojyw
GtNDiGtAn/5QoL5akcNbhUFyXtQ6vr1dboMJBkPttuYc/GtWTAjpzujmYl9pMqdc
xM17vg6LeVN0QBrUXjUFY4n1/H1TUf5iDEvL+NuaHQCRipe2C1AlLipstFRWcvf0
DaVk5ecmhv0YlNw9JpEJ7fRetJXtXw9xi+L30afn4gc8bAmg1sQEFlFayI4V/9oi
vTanM9r0o9ogeAOc53zGgvtA8YvRbderIvJeGo+tYRe4V3p8+PtHPEUJCaMdxyi0
mW7i7tBgPExzGtvwMi4ta4w6pxqI1jMZqQHufE2oFv1MvTD9bJsRrInBOuZTNCF6
6O+l/Zp45bbiPzJDk3zBLYfURswsamoQ9PSCWoEmv4cO7Qqzs65M1rF+Fsnhk864
KhIKrZjxpDQyYt0TKj6F/GIAxZbmufnBHWKJB3YgQZ4U2VflTWDm/Kzx8sy45iOL
XWOMJASRzY6Wjj7RHdJDuBVVjUdT2/VMgw6IhlhPFIo0IBl/ryX4Su42vEguVsbW
jY+ZpS+qltQeECL5px3L7z8HC2asHsoVt0T1mlgZ0vDD0QOmv88NsyJ8ct4U/pr6
cij+Ljfo5680WyYRNyC5U8vCkQyRSaHtzmJjwMCQOEvRtT5idW5PP5IV7xl30bzs
GNi9S9sfSURzfnSGZcP9EndHnbqomb+iG04C96jqFP2rGo16MPXyrQr60kcpPXjE
AdD/1WLFoLkJo8IbwOpEMbJ6tnvnnGjk51zuoJsh21Gg2QC5u9LYcH0pVeQAPhz0
d9q5lgScgNd/qXcptxrMKgJBK+vOCuwzv8ic0sFtbbynZmQxoqpccOqzTicsBbop
mBU51zl6E9E62WpUE8XjFnW2SoXU7wjV1kdlLX7NRdhvBagcpZexwoJArB6bdDDV
Bky3AuIJzH9KWKD/VqBcK7XfJC08yR0P0nh4ORfbTbjYsddGjKNl3wfCG6j3pVIy
yEr9xCf2UGCw422kmP+09LLYSMPWwY8nFqzB5biAwlUeyTlVv/QeqvL5AIX8Tenc
AWGJDI1HzUsmiu6OXH3o9qBnn907Z1xnXjQuYg+tD9kxWFTwj2rnudkhv0Zdnk5b
bmAOLuc7+OESUmVqm0UorspijrxCcY52IxXXQAZ4piI2bnzyg9b/dU5DkrzXv2oc
jOgs7dAAAqgfZT/1myP/pS26j6MuEA3MyfqAP3Sra/O/RmxHH50NYjswI1fwZf2V
s2Suwn504r9W+xX5ktNI1ux+vw1JOLeHUm7JPWfwX886JzP15gBl4b5nZeeY+S3q
zvyCzPpJ90DonPiHFhvmvhJaJwb3qagb1ZAzMRd+ohq7W10hmnGWPpE/zK6DC9S2
oj0N94j4uk6nh5jE5dvyFMFV6upw/iFqDaSY00t6EooyJ2eIwa1tlfoRdCVyqa/e
TpdeRqLs93//9ZX9tPLJWZYJvn1utbHqnQwksWmY/1fqfqu3DwR/0wf2iel8sJW2
fW/guPP0oAg+TkW1/ZtFM/dak9QPxukkvg562gzfP8RSoBy3S7C2mshEG0DMWuSi
uBexRl/EEaBjf7AyP4VAWitP3wsLWpW+3zbvfevBldy02e8IwHTpgPHHvu/wekkY
slJcEi3qMfs1BP1v5yRhksvVEXzVfwOA8jVbbp9bA2J/QR71OcGaS7jR/B6e2E1H
LuKUH2JGLVhqAq+EgepXcZAO3NVFzPmpCR9OCQzfnrKp3j512WzJHUzMM33pL+Oy
jiMS/MtF+tAvcfEmEE/Vb2qxwIeeNJ2k97vkWGoJ45Np5lwLFM3l6tWHn76J7OZE
sRMWgxY9R2rg88lLWi7poMpXutPEOEW8Plf4CpsrnQOF/9uVodKCLXvsz0xJZ2v4
tJFdPM4vOPcECxVPRRn9tzbfRC1lu+vIFT+jHWwej1hk4VqLRiMtESQ2np1oXRDa
AvUv1vXY7MuX5oafzyP6y6C45AFhanypvlUOvLRZAJQBttAf4lXXzlKG6pZjLigC
46mj8PN3kzADrTaxGZWEqALvS3TBtV8AnqxVeBA0ywab2ET5GfV1XDQjcKYh/icX
lRIt7RcrwfYfkbrC5BUCSISF0dFYABWicUPU7MbkcfA52YFO+ZLqmCsEDlifG7fb
7mSOkfPEyAIKt1I8PjpzG9Y9AcjZSgiaECjSHbE1SqVqkYKjtwG89WKcRqyvxqRU
vQSFeaDHsDeCBOmo6/BP982GSSunmGxiQj0azHj587giH8Xj1nXPzdVP9evqyn6k
qatoSqpG3855jiOkCcibxXTYndiPVZKQQ9wO4Q553oja3JYs/xVZwdM/SBziNluR
R6tu8XZEpmxLDKm3kcDTq7ea894aV9Daqan20lWWUUCe+JFZLJs7C0niCRje7elt
qy9hOM/iAEmb3VhdCtDxsROPJiXuHc8log2D1bpeU7rlLy1+3dSs1VQOQk726UgP
j/nRYkrylHm7dQ2kBjhkBtLmvIz0UMWb4obZOqaY+VnGUY0e3oYzv0W4uXbQ3FZY
zbx4JE4NQVS+qtWNLabGW3jVmdCBFS+GU0+zYJM+eRqvqd7U39gQxkeoHXe319H8
c8vsnRQupf+0slZyKgqB8B8RU4nSVzWY6ctZg4zIo8GeFUZcAU5WlsdKDqskE3kw
207cego8rXPNnnfzWxIdfNJs2GmXhXp893aVCgb3nnr1wwiABp6Nekb0YotqPjeH
IZpB9eLQT/dgMkD7ueLegWrKfEF6Yk39EA3xWK6uImZHVX3hOiaViMHZ7iCJQUFW
/s/0QjXZMxsqZqHaul9CHpQA06lf14yKiOazVW2DGvKgG0cS2Fz6PV/+sPKG0QRj
Z5ysGVhwHwo2AF2B5WYUIuZxrlb1iWmPqFoaIDiDIci4EcSLJTi3qB+iencmiGUs
VVMj26czBzx9PMVspH78x57kKMz02n9bmpP0gDS8414nUtMgvwE8vgSfTmy9Ecnc
UZmny0LvaowT5WlownsZScJWs7garddHs+ADT9BZbHSuIna1y905luWuuq5CiRTu
tY7xUqevxePaObXzBIyE5GVn8Uor8pANGjkvA00OyxJHxGpevWOS1Wu1aTplpaoO
ZOgJpv7PZISR0XAY5JFb2L3aULEczNLTxNrnKCoXPouWzd5W8es1DWgYvl9EnEj/
WftOh+sLgVJw+U4YoFDMBZOhfSLkhwIg2joToNer2pTc2ULculMZKBLifitrknHx
w7pxrVDBUYF5D1v2hr8pWoXBJqJ1pdnGnpxQ4QYVvqSZswiLT21wXDOqW1bKgsrd
70oe2KfB+ZK/JHyUnsrxvn2u6l7ACfr2Dt4Qgc5mM5UFVKbcXKNSyE2IB4PFYzk3
+YG8jE/4kyty9sBl/tsAVpLQ0WSiHsgtySma69NOYc5xim0OFsD+gTeoI4o4xlbY
NmcZdVYe2TFhPRWDLsDRl+en1gXObfNZBl99muzBuOWh0bxk28RdjOCZ6vrrLT4w
hs5S19Jpn2MDPQ3GsyHGf88Mkstxe9AFL4NmTPkmJy0D8iViKK3svvxyvY+0qTiw
n06ZUv3H+SubBqIizRqL+TAeHTlmftb44Xfne8H2kvWd0gTTrwYaWsx8m2Kdk5ZC
7xSO0+Kfq8DaMwwG8RO79cpeyUKRaXLKVkU455PWjJDLkI9lNfKRnQlAmp42WP0E
FX7hKPuyTfxg4Y6HEw/2Tj3rImh9xl7j3tbf66BXnxWiD7/tOAqkFaVU+wD+1Sha
7xRzwm1G1E+diGTrJQzNVEptYmQ3nmGxGoZJ/X8Ioz1ZVyaxemCo5YlhqoWZ43bl
c0hCOc9dUknim49h/4uJsr0Ax2Lo1GPiD9+UPbnzsYqDjWxeggZ5Y1EXCsUhGs3K
ObiL7CEvs9Usm2bOJGvjIF3kHv6PhPrMNSf7m56b+mVQOg83wzPiAA+VXCQTrSQc
165hyR22MwUZ0qX6N4GUunyMYdACw5y3nDUgk4DwLLzBu5NLAUKXhspicuH59IIR
7Ix4Fl4wSikI8SaZ4TrlVwLg2qToLXUt8chDP7yJuPRZdL1mFlZp34HOIQc6kP3Q
iI4e8hwoSroqmi78/xDevk8xY3qxwdPncV1zYO48+rz95PGW46jJdYM/QaazYFfv
pezRid1fCm8y3aDQ6hGQ9/KVyZzLpkRRBIqPCjgpgzGzzVkijqXXhOsQ85Xh56ta
eJVsWgYPoYMhTvN2b5V+GEBc6IyWO1dR+uEDFgDHCgZ4X84XDbT8xB1/l3cl8ZKp
heWycz3p/htuYOL5Z6c5rUFFefiFwj5mKE/EMbv4j1AxFHmWdZ1zTSqNMr1W59Xl
HhjFENiXFrkoRydYm9sFaYDR0UdeQMm0au+7OqOZIUC9VK1u8qDMNF1d8ujObw/i
x16RyOCxMdOQthXu6WzurEYm4uLPpOdl11K6B7W1L25dq4QGAFCPOreWIvbXL3Wh
VMjfdPhYdQNFVIzyw06XI0eNJFF3XLeyOJvyjd8epE+R21f1xGffopsKaF2t9Wyk
3KEGTiIpPdPqolRbC195nVOdCaZaVRPiyEqOslz2A861T6CvIz/RwpHoV0KcotgF
/yGUZMrvVPuEJZikhDx0czAh2uAsG0qqMqiyhkv+0k4YLumfUe8wYDXvoJO/ZREX
yY2Vsdjfugkl2HEk+4qcKu0mjt7E6yO6rO6HJ9LKsHYqLKRpfNgxBVdu777fZOup
k3tQSeQcghCs52pwJOvEmBf8L1UozK44G3fgjR4CCMqpsHD78cAM513mDfTvYVrd
89TsWbRjEGYWi8Es04Ka3DH5qjhrZtSKlbCbTdR976GsLOORXJVT8YVrcQbAZRnT
RqprCiRM48D2iTx+tHM+GZ4QKxMVO4DpqzGsIBLDynVVBWGCiTIcSv5a9KpfODDA
4cBhzU/F7b9cYbe56OsI5Ad+OSuPIjTI/RNSmb29CTJ3yRGWpkaB/Q3byms4OJn5
+e54tOn0z+SWxMdGv0sAvQF9+5vaL1vMYBKrMfppFWcBgUHoXVmPVp0OZ9AEBFM/
z8FtpwWV57FBuNKqMtrYyRQaU0es0/BtnZRZTpI82I5+k4KDI27DEI8aDvk3tiu0
R007Cs/rYAQmAhV4ECFKX3MKtrA7A3ACfbBgDLFCLwdNbSibq5d2WSWwaz/PIAyq
T0siDd0xPpNW1gzLfpBlKsgte1AoQ0gGgPiXHfAqh5wOaOCH1Wwj/N5lwM5dS1bb
90yWpdDUerKO/mJIlVDBdmCwHaKJh1AdYUdzFZKAcnHYK3woAoI4cJGQQudZg3x+
kDbGS2xznOTGA/c2E+Yc3RCYohwYv2KFdHbyWdiAboHcSIEoWQGORw9mAkpSnlXN
28UVUJiaqr5kYLLKOG3v+yyqA4vGT9cQhxWOe8JHRo+2esao/4tYQ+bDlg2KyN4y
XzZ95sdyPoShtJOPwUvUKeBIbhfLoh8VR2P+oLT/1uS2/X8LAUNAPcfeJr4Xv/vC
jxvQNLgHh10CJHhmFOh81YbiWd0iySqGj/bfLbu+jH0ipw2Z4ipEX6Ympljm6ljG
haghSNJSIiKG1HnH2gPWOh4r/6p0Nj9OazqN2j3+mjuGu1MUGBroVSrf5U3w4Xl4
ijMBSf8Y6jEYSNi+Ic3Ji569D6VEx5yZBja1wwG5e/rt4ce+KHl/YE/nfoJczXOW
SrYyVSCgLYYfhi4VKE9D4FOpePrPOr+54gR9aEXVPmvgbTBeza6ZVLIMVq8+Q5jn
P1kShrqmeC0SOhyJSeDDU3Ye06P16n4E4jOgP5IaNNXDKxGLtqdvoU+CldaVC9Tb
YznC+PP1QkDfXkpr/oErhwNNGEPFrZJcFLmBUcOh4rhV8l/gBmoknGr2tdsegZxO
cSYedNsL5Gzu5cg2vh/YbiynxCWauJ/duC4ZNLA1ssymn3qZIgC9XGkrFhlnDqaq
6yW67UfYBimKgvWkXqqiMc3GFJAmlAI3mJH8QbVC19Hq3wDrvdkac5r3e7vieXCu
Kcgoh8RTZam8Nb2ejmnANYWEPF3xV1PakV6Tnd0xKAMtO2owqir2yregGpLYoha6
piOjvSJnvC4UsktZAVOgbSiEeTq2J1TyG6agf6nifkZvJbgMFZ/HQiGTj7zU5S1U
TbqKq8El2aPfNeqdAhEojMXt60jC2RzodQAgso3eUInbAyJSL1At5TCnDncyX31W
lVqiLTs7MgNkspDVtl25k/G37NFMLR/sEIc+dj5+lq2CaKabQbyX2H7GAs+fYf01
Db3eof1UR46z6u4fED5l0Qamqm6vyz7bITGdt5zWfVmopa2LkWandl4k7ctE/F0/
z8d7XoBA6PAFQpijvgQi3cOezATIVoRwObNX0tj+RZHtHL1Ap9FgDvildcE1OfpR
zGRc4GK1mCmgEVWfDqc9f+rDpx9NfL33GRLFuJf0RNeBE1pDchHEs0Dpo7kVObCZ
Ne4DG/M/l7ponqj4UliEoJ6PWs7uNl8nVo5SlJYWO5zv272ZFU6i8Yn/kO1tKEAe
PpQACu/y/Rq5CQyrEsjvUl3UEy2jVstsoycK2nM4CXm0xokkP58cKePAq4WAwBv7
idei5Tkdbxf2SJRQ/GG9S0Dz5zO72joFufFLnZ4ZVSxu2qXdLajMRAmjvVKo1gvd
LDroZ7cMujTSwZPz+vWHb3aiAP1Y+DHBAgr2h0EIVoAFlC1ngyXHVahwnHCJsP9S
gZN3c36UzHknesDW73PcPnp6RyEHSHd9jKlHRx52jwPljQmq/YAXBXIxOJ8POew3
X/PDX2Upf27KwljQhWJFknD3IIuUWbBBVfHCOALx/DLifySgFtMFkWr9uYa1jWXn
CN8xNG70LHqEKjtN02LAHqt2dXJs+m35wfHppJH0cuv72K0FeyxdA9HQInod6Ph0
5ReMH8v5388FBmKk5JADSaXfsESVMxU/NUwVySEAsmtP1d2FmwtdSuX7zdtMPyQi
53IBE6yvbEbX8Z00iUZL8yDAbZLKIkB3ciciSFWgtQOPYAPpksmzKZNq9RNGdm1u
mZzeRY+txA+i9/hV6ABE0kHONAMIkq+JrmWzoHuSZFU0gyC5AU2jMBz8Bvyf4vr3
yHUEBksxZCCpVK2XKxfAQhEhjpLjhCH+vNPoCIdhv5EhEyrqwRD4Pm/cSmWU1TrO
IpScF9y4i2lNxNcqjyRA6t3EZ3N2QoJ7qk9vtiIefQEvMMf9dsuRDJaB4WIBZMvX
72fEkY7PqBIjlo5878wNxJjMIDknoDK130wkmXLX+peqmLckciA9dOtWN2+duPoU
aSdzcJS9wvjpn2ERNJ72tqC2Yn0ZH893S9rAeu5zr46GOO19yx0qYBUrVVXIzn/R
MP+RPjiBmIv5mUxZRvpU840jtNbh7+yg68AOiBhLjeWNLjFocthapU1IMnd0m2RI
dHPtinjw/4YPBAicseALSMaTI4iL5uRLyAVkN1f0OvnWAtLSCwIqmMNPY54yXhrS
64fBvVI28R6Qr/KDlGXmAf/T2ajG/HJFRl3fFdkX14xQDw3QiOUNpS1X3a/NvwMx
IZSysjHwalKTqtKlDCiKEMbTnwYjk0AJWffZif9mXskpA8ZooTsE4XppNaA6stxl
j9g0zc/DysbUB/nNXqXdGsqYVoesMZdsdbDu/9uPDvswkoifvnHqFhe2qhZEwKF6
yo8128bwNAcDnpawJtpXj08cjTo4RBaLykEGQq3XuXfYEI0ViiAI8H0FtQz+B/NZ
+Ehc/OJlqOKASblkLiYNS+S8FcTtG8LnJwi3Mpowk26f3ycZrugUOn1KDYSWpErL
soeNDSYbAFspTRD6vB+U0QUGlX+5HeQ7qoX90LRfe4YFRcyunPUWY1pHjhcRI2GX
PoC/5guR7oFn7Y04Cck8WAJm3yVJYpy3UqtkYuIw9m0HFtWlVqLMvl7z1OYz41vJ
LpyDWEnPpL2k5dWcIqjCwO6ADZPfkNddkqTwj5knXJuIyPzeGeu7LCZGunNCytf8
94hQnike+9E+RncAsoKVD0M+FUemSBq+tbies6HtM98Em5MAjgyRUuz6kGiUwdb2
rgqihYwF9L9j+cfwxswLCvuKOOdmVaKlm4ex1oNL5hblZ4QZjWrhCC3bkVhOEYA4
kvYu+KDVIP84AscVOAtHpuYUDFH9eLDvTd+LHc4GfKLOC4qZzV4tpELRN9WgLdhe
sRbm8SaaJiN8rmaMjk/3Cd1mWaNy4kl+OgLBkYE9gt+YraLEMufVktqH49q0nBqc
FBZHFMa8G9sBJMriLFvoSBoZ2GC0aRBRqmcyXIJLMfl0FjCX5u2VJvc/u94IzN18
/nPYz69kA8LQWvxzBpSL8t+rhsRxh79nkmD7HkYR/TooqUG7jRfSrIeQXtpvVb3Z
CtqaQhxK3wBFibrhQMQeMdZgCo3db3l1qe/c6ab29l5B2omJv5TfsZXg2/g4OMN5
Q4FtrS4kkXpK+J1bugBCA79tYsjBuQXpfmKdW0lj9Q36p05Kpg3CAUkOMtAdLs5S
n6Xwqhqe64YtVNK7JBUNrD24wQ66+KAjAZE/gWgfMeQjjRd3Wq6pRgDgN50LJbhf
Jq99hnelCPNocer/yvDO1Yel7kaWr8wCh7skTYCn5kem17nHu1QSNosTHJZPQVKs
drVX63i/T+29Gp6CLiNuIV73Dj39H2qOcYIFp1iihsu2NUhVTZGoiYbrMfPdHoac
knvZW/7Vn4RCvq20r6ziuwU439XezobynyvPTrOQ1vVytHvTtg3VdDup1NjstJhr
ko9IDkPNlV9djEVPdsjadkgt0xLWFpfvDtHNduqt9oyZxQ/2ie9D0MiNk0pCyB38
YRLaZus+srsuSXSah6do0CF+jir6TL2ZyUBktnwpHGYOjemQINhIVLS86OtRLf4c
CF9kjI2Xc1BB1l3nCy72n+EkyPAu3ncWzOTBUiBPcbswxLWtvDFb77uegFtHxClf
izvcHyHM6oO7izbFvwDIIX1SJja00/c7XamU5bFM0SBFa5gygn0Val0UB769VFN2
u6Q4g0IrjRK7Q1jHscWNuuzmY8c0+BSWM6zHvYbSQtD3c/HWpm3lSqAHyd5qfqp+
CQaXJwVH7oB3jvsLSUeFMfO59jjc8o/l1yxDAw6g3xvnL3i+Fwt2+4tHIF1+SwBP
pqxmQ1yNWxqi90oKCPd5gKKxPrXS2vt5rVnQMLwyMJmjcQuybjkvZ4hfS25+A7+i
BfThPEZax2zDSKQMuoCd9Ul5AhN3DZ8q94c0neQ2c/ePxV2UGZMM7DfvPiWEP5DZ
AjWGzZwBN4G/XZpjxjqnHHbBynPX2fNGAmNTGLkkeHXsBQC73kulGUo/B0LStW+R
4ZoXTzi0J49LoGEd4jBTteCNO2mqy1rx++8vjA/HQ57tp/ThlZVfF8LWqozXWZzR
IKYlrKWyNkfacjpXU5//SBEH78FfOS8pXqUdD1kArDuD9cCffiUmbMc687JcsN9/
Z0m8m/dt39FstKNCJOQc5GYhH9H/rwDduz0nK9WbD4PW+MDv49N3pbstBpqUYvyR
SkpbJPzX79fXCD8uv4rv6W4GQovD0xFA4AVJHG89yA5ftxiRN/Ja/pFClWm08iPz
J0miCdC28LUja9w9OUcR6caJDdfFYrm1gfz+aO8LfgceB8tW1mRPSlIXTxs2ZM49
c0I4fsBAXFHHLqmFDhXJWBxwtfzrFRFQC9C3LjZvH4IqSYiT/xFFLbgOYxCBi5XW
jbcDgbyHrQ/E6QpD+kks2w9uLDPfcPK0s+cMzebIfQ5eDtz5w7MLYgkitX+TfTLW
hzPMcu089N3LimzzDEs7WbO4+9qdeKvqLEvJYvoUP6znvEBtO1RgAT3O+iJkiw10
g2mxx45hGtAfor8pYTeaNsKHKYc1hYXBonkHDwQIr+kWGobW34LiWhtIeV0ItYQm
toesP9WvTwiaXfE3viZWr+uEBs+UKxBD+TAIRjWhjRJWMMdEJd/2Gugr3p8j79+i
CoCGdIYvmPOje9n4gdOYfu9g1ZQ2oWTzFnVQ7/EB1RIR95ImEsd7doKNgN0467EU
CtPueXiaLMj1rvZtWoQTU2rpLHNH43uKh4528aItWC+tLs4y5vUOUHYrYsB4bLV/
FVzC2r2TQe0KGlQ/IqTIdpZ+6xcx4MjwBAju366coe0tXLysmS6M9Ls9ggW3snfq
tVRNcT9x3BErxClzcgXx3BnmSxd6cusp4ULh+0vqTID7mkpO85x0ZA0RFqZupexQ
BlejJCUq2tRM32VHSKEBynHSrb7NT7wP4UA+kYXNv0QFLDdaXvdPIHN2go4/iea+
6llwQ+g6z1s+dDLqNmycx+UIqBItOUOWTHcRjIcSIhM8zoEovjuGjq17sMZnAht9
pxko6k4pxjze4SD9246PYDTg0YbZt7X6NBrGtRn4qc0BcKlY0iIyIpCNxrtgrffm
Qd44CI6ORissg1HbO3sxvaHrLiwQKT4NNyX37FNJkj3XFgCPZDw89JmbMWCQj8dK
3+L5Wv66zh4QEaxMj3ZPJUD47w1M85SVvVvUdgc+o/ZI7SoVHTHKDu0q89Pkd/C3
Atayo7EyqTke4l7TAX5lD70w+GV0S9ETw42SJbmq+IoPJJM1JDFGn3wzsZ3u4a8N
692S7CtKutAthRwbgmD93ItUWytGKxjHXQAhDpyk0N0Q5ubdIcTvOPcyh9CG9M0U
eM25FOvJTXUbLPseKfgn3V8cbosmJD8WpohI4kiQt9RD7LE/dl2cB5atpw3+MSQ3
dIvICMqucYyjRuy0uDaqd7x3qXoopS5l1H77WoXyGrMM5+y/N+1E5waPCL6D2kbw
6n/RwKFR6pbRPHpFMu4WRaSay3sNouNaR7EVIxV13iYIu0cx5bXfhVSGxjTWQbCz
CVwWrm9b3gHh/PfGz9pU2NcNw9yobOinB7JjKGjsqq80zg2w27CvpJkP4ZgQVFW9
GP0AytrzbCRmm4Zh7AG6N2k+JPyHuORx7xfl7y72x1liOZX8zUiewpqu5wxBXDgQ
5V+uKJ0LMzogKUh6Rl/9smDc6x3lO6jwDIuS0ha5hYPjM6NZ9ZGLoXvGJxbbWsCb
Ijv+86/haZTlI21uvvEntJEVyYGuSR0vsVeFjVFgNPloXpFff7lorzL3vHo9wW1u
ayDpIeuT+8Uwsm/bIPHs1PTAB9WMvM11NZ1+sEx3k3+/Irn2ayxHIAX2K3q2MkIp
KqGWv+AG6wTBFUdI81SKgxipBeymQbew5FsUpVUiKbR6Gi7fR+RwUl5+F05lva3S
JlN8uMu8Q9R+P+SiJtmJAlNeE48LIT8UUnYhHiGh/ZaFS1wScTZdKYGPNBQVbhZr
V6rOcOf1NAtuavNpt5BJ4xnbbMs13uYFXdfK7QJM3rXcVhOgvUpvtUxICbtdYoRC
RKnzk3CDY3k57eQQQ/wAfItTBXo1UyMMNVQPDMk7e7QBTqoFabWpOE3JRQjPHCoD
VDYgP3HhFPOG5qwNDCBv9Fqy2EP988XuiOVygou3FOKFmb+uMPgexY8k8hnVcAej
05gI2vXvxvSzUwrCYuFrL7SI8awblHjRmlLP6pf9dnFEwzMYBlne2MEABsp7bhiE
g5E1lom7ghvyj8ydF94+0T9KxAXwebrRezrp1R3roWGAR5ZyYs1ZJ93nrSorM4Ry
cOW9aAVeLcgEdYJNIUy5tJuijQoBTIxLrcSLN/A1H0idUOfw0gxPSpDa/2o6qvCs
UZpjw0BM0w1XYHy9uRkF1WRW8xAlkVcmxvhG+m9UGrZ2CasKxXgw6Abcr3tuXd5a
PQUFZaOq05wL+pUqzQhJIOdKeCN++SXaEYAUDowiGEJFhnATKHIma3TgIbP3eiFO
HF05/rzYOA/ud7sZD9TsbDXMF8pFcR2JQmYav4RNgpwmXCAiVlluqMmEL9++r24j
tjTEvnmznVprpzgEhO//b2JnRMQ52wdpzT6VQ/8BuT74rbGdSyrqn2Wz8f9+XA8o
D5DyCDkd6g2AT8k2AwvZqhpZ1T1k/ODqU/CHlkOSc8mhPEeGrt6xYHCH7OZdPkyU
QB7OAx+NrSgsgvEjOuOvIA338cfqNb2OL/2XuRSLISM2NBcdQYq++BTYE53/yFLJ
U86TSsp4e9P85EXJ9AmZn8/k7U5VOFHHZzzxE2Tu4i8boLMNPVWFhI6Ha+Lr3RSO
TZa1ZjC4zYrnA9w1OAN9ihrdJy6oJsHlaQFLlFYTKqXldySgUmoqBRz4GK0e0XBZ
BPu0MVtVzO4CashCuspeP/q23pFNhdv2TlpP/vVfNlmpkHrQPD7R9UqMvnUq9ale
Ekn4jQiYZqj1803wWQLMGKfJcfvFZ+8ib4xOhRC1/ks08tQy6XmtO7aPetXWj+ez
QyYDAXkGozXAc/MTAhnNSNSqDnrw9xV0sWP61Gkb8BvMTTdw17FNnPAdhsm0wQiJ
DTfgNXx2FhCnuobp6udZsoLawYOR9LX54S6pXdkdtx058Ww0KoHN8635vqR5evz7
mrV/Xb9epos0c6+gsYHeUHv/GKjpMbijVnjuQsuEYBnQmVlFMiBurzgEy7VFweR9
WhAzVDqh56Rb74fCgSJvMnYrRKuIcBZiYLAlgRwbIr8r0WNe6FSVsUxiEP5O/JIA
qLOMSQULPUjJRF9VS+GAgZwOGibAwzM4H7UZ9mpu7CJdZ8WxDhtHlzAaLjvkfzsm
wPa9/fNbwpGp5uF2M48oMkWjkQfm2EaSDEsRZmmAztAqr1nXdK94nDEtuICvqJhR
d/wat9h62C4q50N0T4YalnxPtPlp4pJVmvKijBe3nI8JNA+x7CBpHRg0JNISjFau
OMVJ5/yRIwUZc+hM1Dd/XaPrFjQQ16duyOj95MXjUCG78sb6b/FIq5+4aRi7tpHl
IsAS77E6IR5XBsKBJv21GRwtxwYzN6e0+fDsEW3tIdurFjKB1rXDDV4rGhzoMtBV
CXQZ8pf04nkXiP12qwMay6yokY5HCQoWqHP9xrX2K26IWfcl8uQYUFZCpLEZWtMq
5LW7BVBYTRO1wb3d27ri76Nnb0mhPQ231xuynqNod4HFZSZ3A8iDDyKfw6YS/JvJ
K6De7uwhsGLBIWixTquxyunIP3/+h5EpCC9HZlGjZEC8GJf5Jhkh/j1VVE/cczns
fk0JC00yPv4p5lwrFOd4ecP8FagJCU7//U1PEAD89d8B2aPe9ziFc5N09by7nbmk
sMD+w6JvXMychIDOqR1rHr1OtJPth14+pwF2Pe+QGCn1V/zmp5EBUq+zKMLmywCG
gemZT0i1ROZhYrkWpwtmCXDFhdxkj7f5GUQ6PrqFQPczrfPbzld7hKpudwqsoENe
bRffVSG91Fzom3p3hS1OCxraZ+dtDkunAQp5UixbQPTbEN74991Xs5S/FVwh8TuQ
QuGbhk2/PFJPS4BJFAHHr/hyhuYraIE46kS8OU0nIrkopX+EYAE5SenkUgu3TdS6
3OhewqKFOJB4lgafxWELoWyNiT9z/biMFJzcbjbvR2Xv3xKiisghKPdqp3LKLW8B
FWBAhkXr36gBpYjGBellTBVKCtUoEzzoTJZgirCpymGP6gU6z8VN0sq6ALcBYtLL
w8dG6j85z8T2ntDLZ+a4E1Mqe0rnrDTpV5o/DjFZX4jq5O8sfpdRJ7AG5N0QMB3M
bHCYEkl1VsDs9sOVaEYeOzqxjxBTVUXLwhMjOl8TEnJyuu6dWexXGdCBp5Psmx68
VgDH6wHCC/jTrbSN9EZiqu1nYPXm/XqyTTar2fjKGAsdPr87pal5xGyn/0B/1LzE
LB+3m6buJRMp0ImYeqCfKJE3MNUWSUXpLOoB0Fyo+4XY0JOJFexC65+BLDHCPFb6
ZKJwIRDT9UlMVeApgnEvKHI9hCPg04VUsNhS1eJ9MEoWSmBSnTeNx5eoKFzL4x9m
AmnXDg2yimrrWICIV328IyQNvIEbyXny6PA3WkqhSuMuxGWHTohD6IXywB3qhbLu
5WgTZpqvi++l3FKi5eo3FwFHtG8DZy4HbbBkIG0syVrPobu5E0cCblrUOf5kl6fz
zl9MGst91bgX6foVh5mvQUvDztfM5ILgsqzROAxNBOfSOSOEctRvuwCrCi/hMxyb
rbduQdSa+QTdQxPd0N14x/Qre3Wze2gNtvqAR1qDHS9+NaiU8GZT7v8O+l730sGb
5S42ZJiBG0+ji+UqsvjHdf7HnTpDalr9KJ6mM8A9jP1Y3dAblzY7dNQESd2hl7Ex
Y7GvAnhxgnI3x6ZeQLDzCPHaBDwmVeDDLVWVfKuhaXzOqx7UuTpmn7X1EpbzleDL
PKbECdtLUgcuu/JUW3Sl8v1TqsZQWXXt8BJEFcjnxm2xfvPWKzm7BmXEg0L1Jh0H
znb4UlEnc7CXcSVYcxrOj9kZc+jVDIprQvlSoGgwOQeLooA5NPHQBr4sSXij6+s9
g2UCZcvhINopX5vDINEuWRU84Mj6GY7ozOqCDiamqbVaNXaw+8tB4Z87h8DA9smv
5VkGkWyLBtnPRXgb9ualIdo+RSZOus674hU44h0BoCPyRlyERVA/4k46d0MD5c8Z
S+xErWS/L+M1xdQAXlgvlD2m/zEHTmn5U+1/7t7wfXPDeVwPTTe97V94sk8lODwL
3inQijRrYH5VMqtmQKDHyx/9Ej6zz8yRS+gFKkQG4KpYglGN/rFP3MvpVd5rlVgk
mMAPJrdnENS3WjYRucGGHJUZvtEVBN0MLbwSNp5nNnSqE3mDq2Qu5L/RbZN0Jbmk
2pExkRJvXU94a/B62YvybiDTeWIgautMHBXUgzbr7GkJilBHKyR13UiUUsubG8eL
nD96mEULRWbGv06zUX5ZnOxCYaMJsG9KgEBjzQEec+r1SdLi0XcuXU41ngyuRA40
qvErR2paVQHjtkqn4ymcwQSeeJFcuERKWvemibSVblLJPrAuWSmuO9wlRl98Kcnv
mGAhhR/Zms/NyZa+Km3bjokV6T5SCm2d8Nd73z/lgQup/XED01NF+hNu76xiBr6E
oK1hpTPhHr0zINk0W0m+ZEPohJcwYt5bVtPmx9pJac+0Q1rh24enAG/n0Fsxe9Wc
bWAfQANlYMxah/nov1KmrIIredh0lFXIxYPOB7/GSNzuFzaeHfUVE2Cf7UPJ/BKQ
/XDecibzTYLfKvWdEMDB00L4zMjdwTIYCWJBGcEvAWukmV0oE7l58+f/61pWiKsf
9GXIJAzrJ6MUGW0aZHZbiMhjI8qHwGPrRPSfHDUXg/malmdq0m06KcK1yeY0gIwy
GdmG79Lnq3hWg02S/fehWnvsVQWNkXWxkzAKstw4mS/uKLDU6aGVbFjcmyKcY6Z5
gKM1lZKG2iYH0Ol80hRtn/HwfFFKaa3/oaDz9pWvDZ5Be3mVh2aV2c1TuD4cVJ7J
oT8WjDNlNqcMZVbsFZf8/vrJ0/poutGZ5nwXEmPLal7+w3h9o9V7Eb3eHcffIG+d
hb3fnrST4lVZm7k61QIORjSbjrIy/vXub/2w0mvBBclSp2DkpRPvYjA60yUwqkgo
7CLNaPJ5hYF8B/6MpwuE8niF30zdb0zk7KPSp7NTTGY9/TYqL2tji9231xxYUhrc
e2gaGD0HrkpVInE9wmVYd7W5vBwFccda3vqG+9KNkjtvU//1Cluyumw18Vu9TPRh
BhpaqpTbOjkUCgablV6luR/8R/5j1gN+OOBQpElL/vg4EK7peV+Pj3PdD0Tb6pdT
HP3FY+DvBu4I0ZDGY5Kc0KasziksueSgQSqJ0+m/0cg3jqdnmyMGFTq3TbTQbu4P
6OvRYgl76kGeNluvsW2BkMt1lMHfziSUKmIILuLheGlt3B0mGhUFJorgMexJKvI5
yPEyZH/VW9EOJl2qBmbVPqYZDdKgjLG5BZZD80rJpy9KCchuLYArsZbb9A9xIPhi
pKgJZtk0haNHBz2wq1tNRo6dF0fgMkFwZY8T1BnCzqf6JOTd4Z2VE4WmidX96Twq
lHF7lTaPbx2k7pxBuw9naOoExOM9ahZ4CCAztqW4n86jAiG8RgwrYujd867nvAB0
2ua+rxrEoLzscpvQPkWE/RCdQ262OpZCl79QpD32YdKjPp/F5uaQTrInsyAgcDBx
6oXqG01PZjGaOmR7OeA/ID4vB4J8asFLgbm7stJX5ONYz/q7UKJhsMNMUOzIzG4U
gd5FiW+xp9CQ5fOd2VeiM1037bGnk18WTn9QR7o4JmeeawYOq3GvTHXuSL4sIeiR
rz3CLfKzrcpnWaq+NB3ZUGkdoJ9qM1V4Lztf+WTNkUJiuouAVYK5XZR+tj7L9lYt
6rkHmuydfzm0P66WZNvRe6uNMNpwRtpNTcCy8YAjWRFEnw4S0caFK9LokZUAhAnl
nF23u4cs5QuEWooZgeeIaP9q4vF4lb7RQ4FVyWhsRp9nXRbq8aEOVeNZun5kM4E/
x3i2/Hvho51h3n/h4jVWRpSS9bGOdBfiScZZtjWPkNay9stoGVzdTDOqksvCfzhL
TkReFZPdVgRSkwFWlKnuaPBj7NUfv5Iv2cjPy1mJiX0r7QmVyDLcgxAGUOY8hhZO
aHEaBMYVbDHGyjqqpaA1b4qFh7pKjDMSaUZTEmFQj16DFOlsVme/lMrh9fwE3cc6
JSwmWSTtDx7yGHpSo0/Ychm6jAdsqkOBIpAJ353+bt+Hm1dp7KU5XYEgQgfnr9zq
YYcAZJnIqJ1z0EfSvOBuuc1UVMH/kXyPaq+YNlUe/Q/o7LphdPwRuUKftZtuVoaJ
svI84+4uXADQXES12LKxsow24jhsetDKGjGCFWJ3RiNRU8ZrJgBdWzzLom9f9TIY
3I0NRFNqbr/6z4S4bcRhPlVRw0dtTon9G+wsb68m4d5OR+ZFhje3i2IFu7pXRmab
1Ih7xLK1WVsYC/x6/+ZYFkptDrmoaJRhE+um+slaw1c4+CxC5wPljKX/s2JDrI7M
aQBVDJ+ubfyXEtqN5urqWI2U39iMQpWQVskS2emjWS1Ftedq8BhoaqJ39wLl6MOV
ooBO4pbb2qHWzqaaWREzfvsqWnhi2j5KDTzk5Q8QtmvlNXXc3A3sLthdfYncqSGM
zBuhTTPGT5ZSlpmHUOEWQvAU6hhnz/n3VGAYQsXlGwUyInDwJF4YWGVtYW8VIO2w
sBGGttYwRmIsFEDsbZp8W0DiU8wOUsnwnMPWaLIaOmmhYBbtVid0bNNa3fIZKahM
PlfQbbJpiPnNFShWLmwRLFO5mRuDFbYOBJcEIbzb7pOtCsAmPT1lmGiMON7I4zNQ
/eYi5A6sBAHCzDNZn9gHYXQmBQoqR20sY/PUFD+0XcWI56SreslU733fe5LNv4kJ
bYCcshdsJd8ZTCL0ODd74hVb5W/YXwEhpgNUievWMd2GzSdv5N4iUm9U3xZc8LHR
qzgPU1lxuA8Cq3PorxUYOZ+mnC2dbwFVWfFFKdLolEiYolvGylpyzM8dc6kDS5PS
mGbVOY0bcNmP4r9IUKU2K1d5ts7RHjEElyJJ9fqa+8tPNIx2/AeuZx8obkT+2cDK
mXT4iNPJBBBE136KZnbMb8R3ZZ7hp9zt9rXTSAs0BGyvyJVW1C/xocUBwRuSqjvt
q/fpOlCODuE+jPgq/L83b7LLyCSekwOahLxz6wytPC+c/oCpy1A6XugegPpWW0Rd
pMGS6xc+7dcOt0qlF1N5LZU27TBDcdMix4jCG5rLtsNnOzOp1ptcT+cEfP6sgMny
sY/CKHkWDAlMSl6YDYreKhtV1g4lWlpXD0Yy3aiHM9rX42P/MpR8V/PG/Mt7Rq/r
9duFHpQFaH93NHhPx9IlJHftSRxOko+UXg33o19CWnn++byTNxEdXCPF0FCnF5oa
G/5UV/+fUfTA2p4Gv7OBCy13p2RmO7C2zAS1iI6OiHn0OcrsaJBHd+8dHI7sHJ2z
45nCwA8KIk8Jscd1qXA+fWEdmiN6nf7pJW/SAutYLYIk9Q1hLJvY/8ViNaNkRGHZ
rGDtGZNfSbpFDwa7zlGmEY/Lx6vNhNVvA6YX80IxnAYdfjB4CemRdBwqD7PphV7B
AV/28zq3U+qM3hsh/uc3xUMutzhPvujfM4wqJFJNAtY6nCTYOYcUODeFEhmZwCH0
P8eVw7g556BV4tsgrAjRC09SqJNztfebyAZqCxKWX0Ll6ndte9IOSEZM5Y2HuK90
5HiP9x9CoKOPCpQj+whbxmy7JIfR3NPt8ULvCRIX79xeF1aV/iauUhC+i2P6Nb4C
aeubBmVJSm0875hXsn0fF83yqPDwvJOUzMAPqsE36KXg5y8/Ltl1zyBEjAzpxbYz
JLnJCX4k5mRg+d5GSEKufKWPH9dbCUmhSp3I/yU6hPyZk+30IOCSIzNKpfEAO8y3
aSOtoESeNEb8Top4LmsebXLNh/+EyuLN0WBJT7gCjMszeRdwBg5HMT5u6eeLqalU
GplUdNH8fz98bJQ6rRal48oCsISCedCE+KoY1uD7Ibt+9c0Vo/6fCPAIiaW2W580
nz5RLVpjuUyDsBY77bywLCglWFxeSU96jM9MRAkPevziBBT77qxN94hv2hMQYopA
/iGJU86d/a5ZFahYFz8xxCl9bprQ7Sn4xk0XKuScFk55K+Qv7G8Qn9xgw+zLLAQV
dttdVuLL+tgJ167fhHIpKATdapYMGP7zFRuHwj7bTm0ditFOU7ND0kg2EPNAf7GO
zR6+R2yOb9bwjzYlgZvfhcsmEJ9DshuWdanbFIOxMPOqGqKyYAQC5znAkH3yrx/V
mugJJ3kEkN9CgEXWvyx7cGf4AiWtY41KsOlXJMUm0OKL2grm2JtuCylnEWoY6OXK
bLV9aKpruUqsAkMeceg1iblJ1MebDYin0PjeIxwwfkKusEZUPqrcQCv4QM6MLGo/
zjJmhz02TsWeBAlh8ByWbYOy+Bolao7dW7LdyageHBVchp0Lj5HU+xAlya8KtzMq
3p7pctW7OO6FC+AtfbdPBlcoIdHvpcuxMFBqDaxEREyha6vQPyG19s6oA1/bUOVQ
4QO43Z22VfvNCYIAnSM/kxZLuE0FZ4bUWexq1wrlX8JwXrBctlChadFVLJzbXvxR
rbLhw4lKqyrP1nSBC1y9zzFSNnpoblr/REXk4B93ghtZj8x/CqLvC3VSLiiT7BZC
ou/o6OIpnXPc4jLX0pwpibDTbwCxlY6uI9AVDM5S5M8rpP/tb64EPgfUe0N10sm6
Og8O8TuANGhd7TrlX4kaO2VivTcPK7X3u7+9hsjvsW0ecnZUB3+v5TGdAzvrvREB
GUHXgc3Q/l0XnQFfEUpKvNmQafF2kooK53uHdvG34faNe7Ox1wB6lG/xn7jCj+c3
j5lh3RndSt+xj2sV62h2Y9DBPUWFOhpPXwup1Jqowt2rkfXaKCbnUVFeOyLgvMVr
1B3KIyXRaCHu188DqiFAjHld0+AC1mlihEG/YM4+rd/uqcTuaKA9XdyUb/KGmY3Z
Vg9zCD2THjQcZaZbPPWB33xZ2+beZwjEPGaEuXIhgE8p2NXc/NEoLkinFgtatbzu
G8/3uSmJ942Rc/JwPLGcPaCeMClsLgyCHRHlu2iT5K9mV7HoPyj5+7UudDF8NqHj
zqy9o07Lx7Cq1TN/IU5UAHIxUNgQOeIBchBZ1sdHISvAk+5EHyRT+MUmA7hMOeYf
1vam3cBL9tYLNAe8mS8v87Xv3eFSfzkAmXVDXY2EpyHCkSpfY0Gyf5fu1rwGvD0I
m1z0aQeTmVV+w1QtN7DXka8rEMoazbE1LSwOTEM6rfI9473ME5GbdxS4oNvVfIjK
/EwUPjvmu1bFR5G/1kSNCJJ4Is8fwBqfdEOqiYwHazP/dE1iOBqLYgscK1z5yz6F
q33YUnO69yKbw4jM8dwncZR8xC2pAAG4rBP+Yf0rZHZsqRhEnEkqlPl+s1zEsmvX
72sdD30CquN3IV0+qgMp/KIz7NCSMYhcrKH+esJQQdWZ42oPAtF6/dzk67KDyUho
mwXQlHt9yiScpq6a/JK4e+hAE+4pfWKlVPgfpT5UzCocElGUqFjC0DWG+aMXfgtJ
Pfq8P0WCjgV0NX8AFMO/yobdqfOb45iQjOETFYkUhC9+hh7FsgeU0mdTPLtwTo7n
Pc3/Y6hgld0qnPKoOqlZopoJVH2Vkt4djuGc0Fg2XPGHIobp4UKr+CsdaI4ybZNH
DsCxkwS7BLaNjZiKOYjZ3zp5Wj0sqDiXn6tYLv5fNNrogbhrsn30MClgcVZnBw6M
x8JbWbSQYoFaHsyzwxlCyt6NiirIvfPyxTKCHCOTplC84gBP29zvkGa2f9GcNvEx
80yWXGO8fIbYQ+mNdk4ebhERC1IyyAM/awr/f5uO3nENtlVTRoJq2zGuxeING7/9
1YIsFV4+bCVkp6Y6w/AcN+dugTVBxBZVR+HkXDlVK4pX3KhBpEqwFUu29xrtNUe9
pB1dmhAMNwleQ6wY54FYvSUUt5nCyFCAIEAiyhrKtLqaMy9yCj/f8S5UCctKZIm2
1IFOV0R2a0I3hvxUIvrV/3c8fo/XZgk7U+h3ocawHzJCvtJ9YgVxel0zPaoYwkuq
5MtLDeFwjvyUW46XyiQfYZKs5EsWOTEavolq5eXCqZcHVrz5Td1hka3fZNCbCcZ9
Q3rH0X1g/6DRthD50EBViJONf03Nkca4oac2KuxjnuCZE0/WZHaGOAPXyUgeufys
+AiwTfUxB3jP2CclqQyn4un1Nu0Dec3cE6t22GG058LR75qFjJuSgXHd8/3/f3N/
tPVg+mUweh0Z4nHPbhKdHDpLqjmZktobS9pPv23+aljway3nnuFCRi6mfDhu0TyM
6JJjKgBB/ogqUA7wG4vl7Bt1MIN1chB5CIVHwpBVV2lwtnMeQ5USwkZGYvuEDvAS
xpNHpp7JskQ19JztgOwtrxnytQ0QkU4g/ZCZIiSWheaEjvJf68bfs7ba+hvA1Dqs
UZjmP55gBVIOmc/1Hc9aZQbp5aCNvRQJ/O8GTXj6XMTJN6lF+DL3m71tJ2PIvelV
WxT4x/XB6Gtf525TMcs47pNi5Jh2TPbGpNSpbRNKO6wxhv+ySh4CcHzbretXEMAl
vI2Ukha8qtUOjFj885ZBMeSxJPG+qkQX1Qz/B/aI6wfqex/NP1C11OiZLhhr7/Oe
9ilNk+crPSMRVN2gZxlxI3XjPj3tBPjxpD7f+lU5Qboit1+r22EPibJP3oJCVZEZ
xTyA4PMPdAUPuac1aw2sD/8t4VRT3BZnbZfkVVTpwS4m4dIIQMi4Zjy3Rslez4c9
yk4QmlGHnrZ1orLwMCxITPXS0wvYx3DAscjMB043758BmAlk4fEKv1hFy5b3tqhu
W+DfyRHzOD/ijsZT3nkqEuHTwUTesTrIoBmFtnLA+q97C7IXktN5IdYu/61YVPdI
scUBDaS9Rd8U4iYoI3mrv15INc3GWxrdaxUTV54gBsHpq9NuTjlezZnUKlmDhnVj
i4aDbE9PNq/nHdfi9oCu7oHvv2FV/IV0vgMQlU7LILN7t+TOUjisRDmB6CNeN1Sz
7DnYHOIFgJ4qTgx8pVtE7mb9gzdxEesgaDfNeYbTDFwwy1Gky0P0Dr6Cs1GqIJhO
PuS+KBozhuQk4UFr+5J2UdQZiauynOW8hEDnxRBCE/TAdYQpz0/0EMmHiAHxUzxL
rfmMiSE+tXooltIFzAowgPKpPDS350ima6cZtCsUfq4GTE/jG860F+xkIIrExKi9
rQJWk9kQVdzj7KOTM+vHbhjeqCEigrvLcxPBTW64esgQGjJQA3Xdzql3zSMw+HXc
Syd+o/8oRHUUpgiO0Abp0TGQ8Sy7t1b0SWJEuFirPN6f8/UPBhA//zJm6+QHg+tX
3ujQojrkaDSa2BR35nAnQYPsoDNB3Xf4uD5VLxLV5OftodUEnqJH4uiuH90yfcly
nsRT4L5e3ENbsrJOWDfa2liluWrLC10lAXdy9sFHjJZKucRN+BrJGJaogMcTRn79
D9IO8k4Mhd3TSiKs3Izvubf37yqfdKUNpmKITBGdjj6icyVKCoLXFJUOh238eCaE
tv1JfbK9kPQCL4KcDDSSbQ1VU5kyMCF5P8PkdjKsyO2HBiaqv17Xv84IA4JEkm+Y
XfSq2VVLgzRmngDwMIFlcSFJRFYsDRwdVsLhu66DfAnD4KlhL2rduWxnTPXFoak1
In6S/2pe7ER4NLbPmUNGf0iveb7HQ6Bs7K+dtpLxjfpD4HuJQUeWEQn12O5ZqE+p
AjHGfGFmwMEDrqIZoVOHc/C86C96JI1nkKFYdIHGA7KfBl5N2fi6A8HzB3k8Y2yA
4EY2WsbA8TFLL5pu8kX6yINnkX7+2TYDPxGwkbK4klNNeftbLKnEYonMRkRu/ZnG
RtGbag52r4j+huwX/+jPpMywZFXWiatuqUWhZMtoz2oHkDMIIIyagqF9ITIZOqhO
hJBAap/d6kQLVng44c63Efmw8Krc+mk9RufEFF4zokGldQkq2SPEyPGpi3FQGbV9
akrY+8aeBsGqWlTTIRTMYQsZOG2tkyH1OE1kQT1bE2PZROFRUSc/n92V8YgowGc5
CdP4hglwrhKjjik0KlsFEqgMVo5C6RRYKqnkl4WfrkKusvN9dijizbj9h4sQ/PI/
rYqWsEqlXTnOpb6hYzgGNyDYuv6mkKA2kyUw6YOJqvgDDA5cbtKuvSccDRv4DrwI
dl8fnxzM3Y7unEmVvJZJSef8XzLNCRL7ZIUp/lficHZC7TgKZ/JFWXx5sxdoXrRO
Th1xuRcZeuJIdwJA4koWcaNkSwPon/+2JbUpp8Uln3vc/+sP1UgLpgEYRQRjlzhn
lA8V6yEwhcYb9zE1+v91aaS9V5EnkK2d6B7weiaEBEUePxs44jSTHw71gVyk2BOE
P+Cq25BbjTY7rvgP+rJYLGndBPCbYRDuouNh9QceCIV+7SbfuEHZLXTxgvZy6NEZ
IZwE3nw/BsaiLqTng7ZsUQCWAi3dR94AzYIjUeJVvXzpmWvkvmfezo3PDHg4MDm+
BpTEUR1/9xfdXudmRv3oMSPW+77XbNfefj4AVDpMZ5TN8jZGKsxKBjvlGlO53WFm
lXE0LZZMfT9HMiBre5/761fEQ2mrSlJL+8q797AxFgS09W4PkT8A95PQ8uG5HH08
CtdabQQAsUCWWgQJTTOV42daxvrL+iJCLba5DTFL0AXTlBu1EF7rIQavgRy+mpgK
sfqIL3j+qdFBoI29LHpQHdL3UOwsJUf/N+sOa5HugqzxyCmEl5KwFUsH/+t+vbly
fuiPCHyFhx5JmowYrowLt5e+OhnwojwFNn8ihDMNTOuoHLO1YNw7GxYEXS43cYLB
0dwprwj1vJFcNxqCjJ7DArftfev0Doz88aTa+GeclqBwNJ3xf0G6RrdYJ4hgIKv7
2ZIxjK/gp83fNj4ltkw4uBSedH9K5uTTF7rDe0Ajuhr5bplUOOb/TCOUTNUshN2u
/CAk1GSVn+ofFp5VGYf4zNqrtSCRrm25Uy+d9xpoJzG3z9bfYYG01nenFccirrou
zbXvPEEuK39N/l348QbbuJH+AEgivwAKlJ6lL6+Q1wMISUbIJfScm019qGttH+28
Q+wP75TcVYopoYQ+X3ylzcMguNPMCfCbfO2Zbqee3oy5HKIvji744jGqg2gyKqyu
W45EeUn46PI0D42TxTJSD2taupNQOAp/S/mXNFd9qQ8D8H2Imy6XB6D6UiSR3WD2
zOrBqdZuXKFL887NLdnWZXAE6cyYKF9aogPac3NmvUyXct6o0IV5nNEgkxE75ssI
QHhtnCf1rlcDPC3k0Jhs9qC8NyeGE5+VyrufZQQ7a0lxLvqyEriR1mZGwNrVAp8P
8lYzdGVO2/1szc5KBtJnUhHeCFCSeFf0RSRrGeW4BPoNO5OwPY+v8X5irdhTY2DV
mLA+d7UILFyYWlrC2ZcjAVGjY618wdQ0r8jhZadJYiRxqmNulGcICZEkVOMrK3yE
ZCVshGelKRCAX7mOCgD/9bGlfyBAlGH0vz1vC/Bo8UHhLR0Hb2dEUUoPmuZ7kNNU
bcUg/YWYZppL/rjPByrUn0E59Yb6CsxCTuRyfQczBiadeqtxTLejkdKnMP2vXOOM
nJzK6NJtq4BAdQSXTaci+2E5QSIVzVska9kw8FcDDmzjdRvNrzAWHM4lm21Rc3TE
RCYTqY87b3+zVF0/yywowToDc0UgAAK41XFTtmoCoLxbPNuBuzm7lr70IcrHjuF2
ks9s749PubS9t62XAhLaJtuu2IgkLQ/o2XxgI9RO8DIqZeHBrRxlzoPG13/yw1po
2i3pML1EX66b+qbI4DcHYeJ9Aa84RXU4FcqR+VQ8x4GyOnab3JuCiMLgxmIjViLj
Tw1sMykg6kJXgU/vlpIHlt94Dm/Zlkt/m8YpmVrb1Mkn+DLOy1EMecXDnorXzD6H
w7VfpGvwRSqxFYffFQusiHV2vzNOyelLCb2XV4aI7Tqk520i4/Rm7eAb4tkz0V7h
e4hrs00BRhvVJFsh6suRMv6ipzIpnkzZYVyH2l7y//9HCZpb+RK27shO/+SMUDzO
nt1vC8QeFr/KZ3CLlopSMwaMz9K9GW1viZ4sR5IQMowiDQ0fI7AU1lJRjMEli0/Y
rJnf5gapdjXcBEdyaov0Jz3lDimmLp/Ejf6EEg45QliJXJpptkyXm/rY4IxeFz+5
xktRl8hXRh3iPvktMQAldpzgXEyalvqjWkmYblpTeKE+IynR8IGOs4WibUjmk61k
Z12kK1EgzrpfXHd0e3Uyy5pwG5fW5IPFpbf0oZ5nBJIvJaY28yUqcUeSKA3Lj1uf
ZydxxoSdLujxIYbu3lL4LfsXHPQFedg8SO+47badKBKrOd7KUUS+63oM+DK0r/Vo
QNTEikrwtAgsHVe8hj1UeHfe75OjJiKMxlqlMsSGGZVh6jPre8kOu77bu7fajc9p
els9HSQzknM9LnDLVqlEIcDfiF5Qv0kpm6sI7fYnLHIWw5jGq04oSAF+KX5VNEiK
bsFisrZzOVZ0gIhkyl/X2uKZdSCS5g7SO2EAVOsOCUvjqYiSQbQ1nzs7JWGXSIyw
Ag7IkPrmgR9NT/TUnOEiVgFGcM5Uz4b/xPYW7I5rhHgmVyjfNMvGGLvMg2AWtbsQ
hfTVTzl0fo9yE0KV0Y7ZM9w2xlBRBRplJJ6SWQNDQuxF/iFwhnLxXgoO9xsA3Hdx
URDWxUxhqv84w+y2OUp4CywFQvjOTBszFChJayiM5tVfp/HIWFSXpgWTn87i2uBH
MrCMVqQBPIk+jT0sDYzj6gMRVsAw0XSD7lzO9iOKBa02NgOCh5Zp0PVhosOBiX7Y
c7ihTL0BGwFdA5trJMqmfgjVJbpjh3OFNAJHkqUntASmxJdoTAm59bVYmy0/IGyO
Z9g+QWSDVHiLgfbfc+yB0ZLTX1lD8KCTl5kI/DMSrD5XWe3jfe1ISs7XG8w2gvsk
qthGsswm+GCWEE0fqDqO1LAKhjHs0Pfgxcx13H8AaU1CbrX+sFEsT7SCRZt7X9+x
7+wRjoTNhvXY9rPUTdNET0FCu+kH+CObxFIrR9aEq9GJiqqpkw/+uV+GpIm71V+G
O1J8jmU7n4XS7c94ZiQH40BUAW9c6r05LRLpEqMoLET0KA2h9SdZKdDlQNtqYqNj
nS66fVoB5Fy5keriQ/lSgqg0iz30iJEfSr5Fcxqh8hDh81iFq8CUJc5UEjcPBBQN
lRYu8wtV+mDJkDzAhfdcMEwSJNRh1v/0qyacKHO86OCCf727arkSu+YjqaS6BQzu
ivtGn4dRXFcTePjCuMpozmVRm6wFUA83Cdjbr+kQcXdH7tuIj5jbRiR97UF2V8pZ
H5bzX1Er/AQ8oIfz4v+A0ngVoWJJPolEgtNmvC1Z9o1YCcage5TdTy2QAvAJPMvk
ZaT/tVhoOWvZKL77dc/ERuNREMxT5KhHLY1fP1b9xcQcSoFhu+tzU7HESl5peIMi
uJVtfzXTodcDMc56KKb8x/Vy2QqiLXKJp+WowNlLKHrzzRQQLd6qCOODtQFk8dpj
SWosWKmAeAjN69nlaNzdqy19lV4rKYFnb5RDoDVlCcvI3C5XnwzqttGbyYHPgK8x
Ea5IdvkCe6ioXabp7QZrVqqyv0OLT3tGWJDKibfzQBtj/wOqb1sUqVfMjOz2nTi/
0mVIPzzZXglXmw90FKaPqJkuA5ITCNwG4zls+a9Tfm1QjT100Wp35uCJ8pgLEHoO
pD4x1adHWfq8A0oOU3UIZ4SikmApWWP6/gBG58QwQfyvpN6owr614s/a50VXllrc
a6yfdE01K1QynE5W63yQBmFbqpFqSzMb2J/WR9aE4nojxSgNtvInzRPYinxfeKt3
AIBymGGShA2/BlbAm+wVU+N+gY162C8X3pGGJexz9+1Bj6OiAXTDtuppkDf2FzDG
J3dn7GMj708geYj3sxZbHkbKJELCbHunKMLEBCD1E9jMzWl9hOcGQvQlbmVfniQ8
tUtqoEmXTwi7vHjPQl6AAK/A9bONowv5Yisl/484XF73+AFBquLTR4Ta/qhoPsdn
adGBiHUzAFGrzR5q7vcUxh86OjwNCLkJJ/tSkGXXMGIKCof3btqxsDeCYJk3HJS5
sOb9CR8Bet03bS04L8XOsiWkaJRkLdBp+FBjmAS9d4dz87ynpMGaXgY02BRc8Zvm
oy4cpN5Ibn3eUccGcTTlZEDu67XSt8NqvEm5mtwWdepCOJBEOC6mT/NmsAqg64YE
Kl/uVQCEuzsgcdsxb1IkjGfNs07yimtxuSaPoFawrlEqs1LTJLB4kKRbNntaVumM
rsXDGcLPPoBoppByM9/KNzbeBey/5cVa2x5K0LhjTn7ceZWkFCxgUauhdKjOJnzb
qPyT4GzsMqTV7mJa0+CZZLSV8HdWW/I62t+sSukc2onC/82xKX51duCVnb2gWgpC
xPvYr/6WAZNUH/vUq1mb4YIwn/NXkIERaXYTGxsNhWJqj/7GLpaEotdLf1sK0uV0
YxblYtg233FWnJdgMJscaLqw5n5T50zgL+NkFhW20Rkm3zI4Ng6cCssIS6tC3Fil
LJtOOp/9IKwMrIjrVaa3WFfHVFWCmvX6bl+JsMph0sFYMl97WTVPe0NpGztoZ8+r
0250J1fgfRERmSOMLApUiKubPLJGyrHWM3FkJ+MAW7IIic2nHaMlhVtQW0KBmfzN
5l7HofhFT3FpiIlQE0ANVDFeqiFG6K8ImSz4f4mwmo+8mAn1UfZAMQKkTnZzAHjK
SkSulFhZTiP3goNtruPeYy32ZBhLI2D1rfRR9ivRaRQhTRzH5eOw5/KmhjjaUl+8
K5+NGYUU2oWnArwHpYv+heHSJ1VtkXbrNWngSvqIHBb5uLGv5JMvWT2yGm04YSeJ
k9n9NxYIOdDvJoufqH45X1C9im+11wHreACJy6doBiaV/7hRebiXpYTnLNvWSIeL
1RP8XYQPACdJFMARP3U1D8vA0TOtOR8gSioxaGo8zBbyyWHAgfhe2BlqORjqPAiK
0lJUkdPe8E7A9419EblpoYOvtkfCE+twtD6VGK28ylaynqBpFrFunjURO4CntKJy
guLUy+6iwz+17tRUoUavZv/cJb540SeRGGC9D+i2Fn887jUYKtEWWFs+9RtTbwZB
u3QwAuDythcqxH6G2ySIeX2a0puxakdPQs98f036qM7Dc2zCU+k7FZX38gB9pZwh
LkZm4hZiCZZN8qxqMPVITbho/jNyMkBQSu0QXN8vehmqnKl+as+BhTd3iZfQcL+r
1f8Az75oCvETMKtg5X1BriyhYW3DkJFFWS5th+d3QXPTdAiUJ1YRagK629NCk4th
idfXzV15NMAysSjfucjRT8Fb17jeKjOUJM1i2W1o77yliZMgR3LWG417Rvid2qfq
3Ejknv95XwFlrBWy9gD0apAwDTKfctQys4lMEZv2Af5JtbL6EBk6UzLGVkFXLaej
ptszAz+UGom7uYfjZmk5RJOkGzwEfd6mEVI+kIsNWG5kg1TJSZmb86E068nEZg+z
WH2/WJU3bB1laW1XHLhPBV+zFdXxCWFXCTNzbCD/c6oWYqNgF2FmuSim4h24n4FL
CeKCprohjqzdwB/4zMUK3Yyzn/dO0WKXVY+SUGyKU7ndnnXMZOn39NmSa6IrolwB
lLp1QaOWOzADtpLXVpRNrR0+JUgI1JWbZJQUtrXLF6s/Bc0KGurbkWAPBG0wfWYO
onj0IWvxPY7Qx14vomK9SQ1bPyRFkwX287yg8kosu+lxsgSg+ryBZnqw3rXH7Xkm
auhCqoS3io315Bx1SjNA40VJiLQyelBvMlz+xPKvWQSGHdiYpFxWxIQQt9omu6V/
HLV3ZHm5M5qIv/t3c3QrwoUrGb+lJJ+sv+zrFh0Wz38Dw+sFdF/PR/cl29orFQvT
2rVlXmB9LLW7EVi4JeZG+Inbp7glUF9upixRFoT7bBAxcxvIbLYjFqsv2te2qDTh
s4L9XKsbukl2pLT5gbHiRDUdrj8QtaQomObA28ej/QM1TaKf78AdZBotGuuHE3D8
K8J8BEjDtbdIlBSbdhhDjC30ZLEVY+9jmG20OZQlKlAiLGjol/AX0bbdXJZM4C9a
g+L00z448zu2tIMDZwnzXFqLMSK6SXgFJrSZ/ZLw0/5HP2V/aHSp+ztg1I17kUJw
O9AxwaIpfDYk7VotrGPHvVGmk7YLzelTv1Lj/ayjk7RZyeWn2+xucNBd63Ko+VDH
IUZvVWs5MT0chr69/As44bHYXArmh9Ob7sW93x0Hw7Ew71dTCKLtKolwVk19gk5c
4B9GMo+/bSMJULghC+Ypif0QGX6/W5S4pJj8qio8N+lDiEJpcFy/57Pdat5CHH2q
3qqQSPkTwoqddlzyRfbjgFd9tttzkompXlcWh1Od8l3r9HS+UBZWbqpk9YHHASJQ
gWYtim1cPdI9gTZiwRjhwby+CZeaS/Dy1TW+EsTT1HigHjj/UKZyeCFpf8b/aHyX
jI1FRzApe4l2JJc1ua25sgWZd522R/L7mAQSu48VbgOzz2/S14jIvDvRaZvPoHv/
gdxR3VbOe4IvWRJNUnP/bt9IXT4yACH0d1YBS8guAyyyiI0bOor8/wiOa3WyfE9F
akA0iFkdk3SU7hFXntjHM5+7VG8oT/5+iEqb5QeNGX5wO5cWsg8yLsdAFzS00gy7
+eDQu3uImABW3b+WgBNX9aVyh8N6ko1Rmf/adXQhGL4GzNFG5E5UcGWVQDlEUVxz
0PqXuUHh3e8EB1CD907Yx33QoTuh9nhCfC549BsRybgdcQ6/r0U8swz7qbiBGdFE
XwhMt7i6/ciR2TiG8OpzVYS2cO3PEfur/5tlkGFG5qtOvSD62raTjVw1qt7MeWhH
MgCM+wQwJ1uUawaSOhzwplCAxTfZM9P8RsGt55Dhb+TrjLee4C1YbP6cCqJg7zt6
bra8P2XcAMiF/O2mcPaJYOa71I23I1ZWDOThGZuF6m0lhlGp/fMUkmFeoMTtA3m5
oWh0/laoukJNDT5E90/TSVW++uo1zB2YoRdM8HeErHEoqlTGiOA1i0isvpXNb9T9
aSPFpuKxnMhqt4Y9NRWcs0xw26u+fcCov83/9nYyfuxh/vN4rlrDY9bN2E6MvXAf
uVo93TKUIi4FQmYbjG5qdBclj/AKX5/ebo5w8AVl7VnSLSy1BtFdE76XddNNfgyx
xM0N8R8OIl0KEPEvvZAC6r6rl/w8Sp5N670833I8c61nitaXlEIru0/HdtsbDIhQ
tzcVSVriVsunbO+Ghxm1YgPXZa+RWYrxfya1N2pP5yNd5OMkYbUmcNyOoO/Pz9LL
Np9m6j2kjRIN6eVWrD6Kx2lBA8yzk6TULLDODHf05oWmAJin977kyYZudCpW/MtB
KB0i29NbCXy6L2EUbtx1+1EP2bGr+IOGmXItBRBNS4+Zcmrl2gUHWB2hCgNjC1rH
nPEAcCP9epNz+IREnzC0mcaR9C6ZL95o31vA/daL2ci8nit1Z4VzoU3j184cEeyq
ZATh96tIDnL7VGQ3xESQMLAGMVynt3laF896I7DqrNElzuyt3vexkuSZbV4Ww3Mn
BQx+Oizq2ISaYILs2bP5lM1yQDKw5BOT/T+Xfp+qlF8TETTb9xvose/2sdq9tL6F
fA0v3ZyVYgTSl0KQolKrlV81i+ux3n9TOk+vG9TjlCmZLS6t65PGuWZHJzH8Et1e
BdMi3h69YCO12dvYWM36xoLx4brFXWrJoVrjYQ3/UJKpZDgyPhwnfwSzqabdbRAK
pQuOB4XmP3liU4msG3I5HixAVP4ffuSV88aHCs3ERCySf1uB73RR9Qj/Tishyq0H
bO3sLFYY8Ym3RuLhh10+ItPC8LBd3OPY5gEH+Zsfuukf/TbT4O91LioR7EhwNXcG
q4f6ndnvUPHttFoklf00IDpDRbVeFLdy4YWFfCN9IIzteXnfvhPCOWncV1Bo41rP
yKLBwdWv+uAsexQlCcZcQ0OFdO0VMVmpnYBTGsKSGfTOCZtSL20u5unE7EXueLNj
Kx9gsNB5vqt7ny1EOAmfemcq5009AsX2immLohCZ5oiJ2EBKAcedqpAGEGBi302m
YeSB+hZIISHIhB9616hGsEuQuj8dBJ0OUrsPUWasnArmPy1qB05lzoabQqQg0ALK
4EHkpAmrUMNb5ZEZ56Qnvd11jauu0IyGxfWvIJIci6RHAAonHBF7R+lCZErbRm57
XAFA23Z39qonh5Wlt0ktuszdqzi3Q27u3mbizeIB8vlVWcCPgSPdyuhQJVlIAjJB
V/gm35q9GDIZqlJ15o6H20hONRZtOKQa2OyEST33JwfEDIG011qsdPskQQHBChDC
KYA2BnIkUOKkNnRikUUxIYfVbpx6UHecjEq3CxmZpPrj0Ts066DdKWc5I+66K/EK
fDMFtvQPt6jPeaIMviSfNAT+0kZvBMOcnURz3sUdZjxdWRkeKfO+VSGruZZ4KGTK
BrexoWLlUPGUwLZ/jEduLfEwLQABT9/zbilVbUu2I4F5CdGvHEwzX5GkDKgQ8LcK
vrlVS/g/nkBFWJ1Kc8ggbewl8ect+pgj9AIM9ry5yZNjX638KlDohjsXYSVbCzqB
4dT8zMAuNnxa3+aSovRCJednXsLsA1+O01G1R3lkipCug2bU22hVJJMcWeMrS1Dq
zVXHKx+lLh29ONAhHzyU1dEFpxzG+noCGNosY34Sf37xLGTN0GCa4NuA0KamFRk8
n5kXHdjPprrQlAFErqZEqmOD92eqQCN08IjnFWfzYSEAnzHWUjSFAbf+oPKf3bNn
8x3o1WeGeOnfL11j5tbZkZuf+3xIo+am3XvqKFs5qcBOpM6tjSUz6y7b5Sr6qFp9
Yh4Rc3NVv3/Ucb7dnD88IKGhAGc1eDj8eBaBv0DQUTh8VACs1QdUs+wRl/Txr1Le
b71AGTsTaIzDj/PrsePBOeGTmABmeg7WcZilW1j11xCEUCp8IiwPaNEeGblopzL4
3yX9UpXtWF5kozosewUZj10Z6TkHVcrkZwwg4FtbVPBB/dHrHA2/f2U6oHVG3pGP
EeRT16/cRGE5N+5PPkGyY9EUEDTOfELaksOIudFI2GWbwvKgOlcYC5eo9BS+axnD
huQGBXxvpfHiSt39gxhS8mGrxyT1LdUQHO685n64d0WTZ/05fyzKLbpdzjHfuQOf
mnl0YZmOeWZRadD4roSPQh1X4023rvhPXiisIbFiBLidRK2MF29YUfnzMBdHnNj7
+DtMxXWZlkxovThlVI7SBmxPCyzqRa18+pqx3mUWKJfddH+ReSLb+CGdO0ziogA0
4AFxa4UvBEyix9yC/3sX4/DYbxaRa+7TUEoRcfMiHZMjWc7okQhtKKpZwLT6ZHUz
Quk8+rrfH5gY5A9BVadwfDwQGHnWCih/6koR83LOY09Yi5wb3w++nz/30AJNciWX
m81L/fdWGzGtICwPX/lvYUkswGsirxLz6VGEO538sre5LGYg996sSKtB1rkayCJm
8VDN4R32eBQTHsFwqZ1VJFZJjZHEPKNgcm2KGxs1Ag2h8Jgx+/QzPI2ijJhNeOJs
f7oIPQq0od3kKKkpj5HBch0dyGgmZMiX+IAFAqyUy2J71zAE3MarN5P1OaLOahSo
XkyPhYa+HU86ki6BgKvFgKRY34kXlB8UwoMDSLQHhzvx3sB3nlB8mqL/AGu1c4s1
WYCSTMX5Gtf3yE3l8ljt82c2nvMunSAEulaBf7fBh05Md89scbGdUBhaBJEqKbzu
F429vrOD1ji/tvUTBEiCA5uK0wnrLsmzc/TVCmhIsjDuAYD9kdJ9fpAdFK8YHTZe
3fJOfAsT0k4w4nctps4sjW3vQM4m34ExMDhdafmeksHa7c1uV5Xt7iPLUKenOuVQ
Bhkl4eiUb6fH9ToSgdHWoTYgFnrEcxlfKDhW2hJQXki67ZdQDsZ3+5Cw1AaLK+Gd
vZOFcN16/yu9TC2PZAR5B3ID479xjMyEaJWO8vRXqDn5mUvoKymFBRYLXdf108DR
fLZb1oRyq997cB9/V850mPqekkI6jILd/wX1kPqZMZcm9KAGTwa+Qg/gvxNtcwOB
QysfIQjVP87JHULvF/wgkxmNAF1T9KwzTZp7vz4C4E2jjBkJWz+mwkBv8n0tyyJ8
lpSCpw9dZPPebR6KHAUTjJR9DHmjBV10UnAwDlwqbma6tja4HuUllTG7uYzLljOK
ds0lY9uqLQd3DL7mnObgolWzYULqZTqplXO+EuVWpHstApyXLhLWc2Azkd2t2l+A
tuRp+2P3oirkhWzahT3dzrg9vodrDfUylwhd9/0YOrfQDIDqixtNAnzPyFBEJann
73yOKwbkdR+e6klWvmr8n1YfcXaLXTkAdzwP4jWqHUHJ8gNVIEBarcQmCxlr8Ah3
XPtjDaEiHaxll5LcJykzTpEzOr0G1tjr+vQNBb+EYALjpHiBt7fQqFA9C+OFHm08
RAoI4lLb115bsBsEiJYTtUt0TQIGACMFmo8XY0FGaaPUMGw4dNLUlTZT+RULCHwQ
0QHmIc5Wty7YOArsIyGiv0T5TfGKTTkmPFZ4EB5q8CrlBm0GAqmhpoFA7SWgumaC
gLGTehPxi0hJdb9jEt/juMiIpJTpSMobn9FG23qdyQ3/gJSE5eWyeRUm551fKdu7
to5gL+dQA2XL4ZVDg8njuynCrTPbtwLKPseyIt0f3WVwjQTDYQ5VIGiWwzKh3bvK
TlvyK9AWc15r4sXrsKNzHs0QO6yrJNicjsHWtgBrLpHpSjlv+9Z8nmFoShQSYugS
2ptfuPT6lMMf/AJjsJMw6qxbgv2dA16CfLh/p/YJIFE/kLJ1ox0X7K5AYJqBFku2
w2xq5wU9IW5uyWQnnaWuULkf5uPHL9PKYKte2JdX/kSaRDpqY6QB3uwAqFPo42g5
M+K7wJLBB7kz2KnA9gYZykBHx7+Q06GbqIfZH78VXx72JdcXBIXjkq4oPAhmKmZY
NXFBiwUQwYt0Uwtmaahtc4WEEAxaw+04lJ3eaYZQQlmEqm0v+lq0CbqjfBbuJ2EN
P5MRRPbaLD4PX84Y9mF31hXRwKzVSEuatF+3fanqDfGpPwoD5Dfyt4Dlfhbr5G1B
Fq0IWVdPViXvJBTLJmElSixCMqW8NKYnbSYqcqaF8OLfKzfaXJVGuL5Xp/i3yLGY
j1NU48CTLjEtO/Fo3PRrcL9k3vIVqgUI7ba4zDIHrsiE9maMqx9DwIHozVC2sptU
gM+uHMnzDWDZ0wVd3d6pO30oBO48rPxwSe6Jek8k+pbhR/sh1wh4SkenTdfrZ5gY
HQ/160A/tpjef9UGpRYU5NvYro4v7sJMly8BFGAbHOYt669kuU32XfPT0IK/w1Xf
tfOL3irJ7q7f7NEfuiggLr4pi/Nca9BszohAvAvjB+/XzOIw3moy+3LZ9NfHnPWS
gXgeWiv3t4xVxLrPSOllO29m3UI/D33AJ4+H6Vr9HZO9ZVlTWV8MY4CPO8Ml7ggJ
BN1IyVa2LYaEsStMVPVX33VAmYsoHXU265LOrvSXMHxsV8EWPNj1oTy18HeZHxMR
Rqhyt6esaHj+KZh7p9xGMqnU5GfINA+JbNSZpofN2X4zbl2+Jk2QqDWD3PO8onXm
N7YZNSV8wBTxLkquhB69yp5PJyzQGd8JzJf2n8eFwsDk8YFm+DlXZay+xBOhofIg
E7GxNzBjdgLSZX9du9EFcA1wnDOHgHbl24K0pQGEYq3Kza4HzUfgGJyuiSnTRTOe
Q6eCLb9iatpRE9ZpS76zaSlG4WSh6Y9t4xK6A+pwyR7Zo07xOo0hTZgPJOk7udAg
XActbrSPFQR5/RG/I59IJhEVYdTjsRfJhMslUA3ppCMrFheYdqxiTDwC6mhuZqDF
ZAaE91sy5BXhaNjv6EgqFgXWcESqCl4A9u0q5SzaTVNUiSWrHzfN76WA9atTf2Xp
sdddldf2jzsOb90OiWDntXx/kLK7YY1DJiHKHS3Ic8HAjh0aBgSMwzdpxh8Iyjfj
p1jsmsEr90BQutmg59s/MyOpmDJKdhfsIY2bZfGirWjMCUr3n4mLMUxLpG65uFGU
61VlIHKkyrF+YA0yAvoBx0laHPcO6PB08sil8uzdlkmrruWNIR9PZICrgON72l7L
IGH2Zk8EStGuAnLDrzFybQL0R0tXDEy2y4LN+RhXRyFY6BZfsDaobVYTbOUbxXcU
zpW7lIJRHpnINvTEOmhclQlHdKU32f+P4HTjqJVCPgDOqkR4X8gX1Pmer9L9bJ+z
ZxF9Jt9kdcNphiR9oTT8qzko3cSglYE9YITZVNU11JxhGwyDjBH4xZ6wj4WaZYX/
q00y9ysZUv0b6hT/5TeFL9lXVaHhuQfnVZkwG96Oz5QAU4HH7q7Pnn2IG3rnOQmH
rebJyM3RUW+bvVheYf864A9RI34d5LZaushRkTNQBW5whqXGuZHdl+D/MNVs6NDT
x18bRbdkCmhR9K5fWh0QehqtZQFABSJW7qYi9khFF7TerPADwXNGN8DQXJzLA7BK
4CdQQ/XApG9ct+Xe2+IZxExldZzYNxOBp/hEXJySrYTxBCxnp+5dhXvMl4RrWo6v
O023tnabB73AjFPDe2dfsiMM/6RZg3J6tYWQ2aYToUevYd3Ztj+0REr18s/3d12A
9ck8Ot1CnxjKFI4NC054mYE40yi81IQvq97rUip0gtOBI2lZgJ6d5exS3Q4AVMuA
kKIQvVZ4M+IBUbG4yFFinsdc6Du/op2BJfSCisp5t8TExmpL8oRYivXxz0o4clQx
mTfJNG71E6HuE8SE4mc0d+yZqKEufnxeg3M2wm9+L00+MqPDY6MF+zJBJJBdav6y
ZziJGSxSO+f43+UB9GZok6enUGrunZGtBAEl8i0YE5euEqqXgWYJ1a3J4+pTDD90
BD9ezmgoU4YtD69KumU7+/su8HlIQ0TRoh70VUiIZsB5cJ6PF1A/V9jmpC18MKWn
cqYLne+FhCnBb4NJoguiQQtAw/gr7vhUl1qxk/YoB4XYI2WjQibCung9CmUeFgOl
z+aLhWJ8JVWQEDqx73O2VEwUop92qSycfQWnHNF9U107Bv6MJ3/dNqy52lBc++zs
vGlw5Mg4fjLbaBu7R8ZvpxfUomz4koQ7HcBZTmxdpHY8cGwx9R+enTqzk2EmNveg
+giPWr+qO6T81Oc+kaNrQZRRIPo3qCFOO+ZRt4NTHAU65gF3yH31oUhiQOaonkF6
CzvjdP5HyE+8RaN5uQ+HRX+0HoVKs8ZyhhAF08AwpZqxD4WN6yonWdgWl6pSREC+
RkZ/IXPG8KNpxCDqiWoTsCDllcIEwjICS+whqyZDL/gGY8lLvnq96WMfc0U4/78q
IxxfDai5c2afQKK21rGtVSNMuV+7BCsHHS1FAciYaAOaMiIT7j+LkkLEhAhysJ6B
2z6zGnKUKCARJ1u3NdXZ72qYUyPRDbxycsYmYmLoG7ysBaBWs4RqH7SCoplq2XUn
H1Tr0hkTFaYmFCiGQ7udanVSC4AxKZKlgfNpCyVz853rSo0atSBpIQ4V3uPHtHIY
s3qxkw+RCUWeDiobns2Z6mvKFDYDP9gEQttDY1NeE+RqcqhsBRHRZzM+da4pyQyY
PJntXVOIhOjsyhXCSsUm7ZgsyW/ilcIqEguEk8Hvy7Ji+KFBd86dCpRkeg3/FWJo
yU6piXLDkCil84NOeL0h+GcpGigkhOzYU8Ige8baYOiObyoR6deG8R8vFM9bkZp7
srA+FbKwUbs8fvImRkTWkFThAg0BmnvJ61vYkK3UGVCVUKfW5js+45eVFjPguR1O
imDJvAgPTOw7EbXJ3ntuP6uBanVkQFhkTpGQsCA+Mkzdhpe/TQK+t4sVPvc/6jBo
sMBoZYf3/yO4tmzR9bvF1GmANsc23jloNyKcG/Lwggd6meiW5rCMhqF9sQyHq5rM
VJ/okOVNMM3WdUzfyV19ldR0JCCkdfx4/xR2hFDODxkSue1+AM6nNHQn8HNxEPqe
JgMhbjSfFdnNIpDSizuXZ0J45xTuvxE1P8690jKYO2s0DimC/5H/wHs7yFGQzKVR
2+9R1CkvG1KxWOaZuqc1PvxdCF6rTO5m6v1qxMgPy0aIR0/HTpofAX6CQirLwSVu
iUfQ8qICcDsnJqUIvV9RzJeqy90yIM1K+vwPONlV+DnX1FUdpNJuhkJJWs590A4t
e6dW/CQ0pnkEjszQlDF8cHg2RPjbYH6HstGohbXWskZDpNjxCPX7wW0KddKY8T88
g9wiEPODUkHHumOWgPj7BA3iOquEGwnW948p+I60SM4S3JkNLQkxzdQWb/HDtLon
0QtWAMJe0TsTBsmlZNj8ee4E6jXr6XTmuy8HWz4qqCKFneVH0JEf1SEm5gIXN9oV
+53ax8AFihXV2yCMLhASuhE4a/O4lhy91WltURV39LKKdRx6v1DRmC8xhEBrXfUo
QS/HrWBhQK2O5YcVoJ262v55Iq76CLCvzkk+JSx2UGFAPTiUhZ8ukYvXo182mHbd
F+sxGJ6xCHMcywSzDzQDxDBvvhklmFpeOCQcu3uh24Z3rOlzJJiYQqf8xZZbgAnh
WyNAH+1/XaNdHVF22yoSI85IFSlIjOqcT9++AfHu1jpBrVXWNJ9T8U5ParPlt4ay
xv7bjE+7kMKl7+BWZo2DfCf5JhTyOETAKx0QBh0kxGyvVS5AXrzmCj/1RmPt0CXZ
+YXF94tVorqtXSVlNq63wG3weU4/xfjnZQobXJuJ/dibI4IQvdtVNCcLmqG7JQun
4T0EDGVJs6K/8DJaqUzAYrxHsKJjTdRfBvUsL4SpBI4YZSAjFqt/woNkAcTG4Kzz
vnW45Naku2h0sLhgDep/gvH6kPsl69m5MPsQyE9XVJsZl4Erqgc35ecU8sNUCfsw
aKo7iklWNKXOWUloDzV9Cnu2U2YwhvvzLpSCi+8JUXWfTVfsuMvxbwAogLmBwrcW
s0kvw9FxXbGVSOlRsl7tPGp5WjDpb38hbv8ZD4+8gRCGErUb5W7rkXYxivtinEL6
dYZf9xhn1Dh1HteCWT6UJgwwAHaDYQUbaBvu52FmVoo6gpadQUsdSMykMiCUVN+h
LufvMOWkoZmsGOLi/epzH66BErmp3AKVYyzAyFNgh9kTAJeR73UQC/1P8qtEaZmS
bcCXbUZ7ohW44NdBelELReTqxiYiH1u7LUB0/hDshLqt3KnEh22npMe1HgL0wRoG
aGp530wke+fAdFK5JqpG9XfeguXI0/BBQt7sCsQv/90akLxf6gde4Q+reidBMFHm
h5xxO5zngCDQpTAaNEYNsrvCHeNjxK8+bmYLRY7B/yGHsD5FexPGR6AUTO8TSs67
NDsJSQ4jxr9Ui6edgNEibjaDKtRzfyw4wfl3qDjnHlNW2/Lu2S2Bg/E4YABBG67Y
iPYs6K/y7Tq5hlq+c3CUfKVpY11xfNS0qgS9vxbmXUIxOs218BN2Fxaaqo/PlYcU
ZlL5Mg5156++AhRwO2k3bUD0H4EimIUuFcdNZOHgbcb8Sf7oHRjUgbNtyNVIEU6v
kYLn16WaxKRP23/T1d1y7IZpyGtjfar4ZHpF5+tTbc1PYAXuzeMCZfvPbR1oUCWQ
uhLDFjEI2YIa2ZkjxATd8/0juwyf7jIJGNq23tkCr4jfohEWWRXf2pxqubwqdQm1
DNksfb8Dd8CCY4ceFA/EEzvuN01/olR+DUOnmz66PKhx1m3QosxugG5PuWrY5TgW
EDP0FwZXlnOuE53hkSDohTgkBLlk2XqGYIYXHP4yDofbpMZk78sZ3nzgNiu9pwEZ
pyCv4WJKrOiyw70jebZ4vJGocupo7npTF364uFsJWrft8jomo5FnGmvUAzHnB+iy
m7eNOe8BR00uxmW6RLSuYnWK5JuNxiSON6rsRViIIwaou2F4ytlYd45g93Qyo3Rf
RfGD0BWi0ftdPp+jNjvpEJ8uLXbnjFFXaOJbsWKkJamAei8BUH1ivLQ+2cD1uksE
B87RtJiwcNdDhPHQ9yP2MtEUYdYchRc4BoHx5q57bewbVul7OY22DagkZyjcbBgu
5M583PCJAeKN+QdwmlCyNsXk+IfdE2OtyS3Cjc+xJClZQE5V/53gct8QyQF/az8F
AQHSN1EklT/SDuVdOwpXYlzLRvYlR16hc2buZb9HIYhkNV27OFH880TcEPPfuvzB
VhgF7UaVONg/wgxD/sOf3GmOYin3Dx/29EMOJyHKsXr74pbskA1GgWeQDyDiplR5
m9lPDeHpxWX7YhhHa2zgNGpPMDKPo+m/fTz3E5g4OuB0ou7ElZ2VBmmyO8Potwlm
+JAF5O0KBUS19H8S8/z5QsUc0mxHvtUaHk+srceROXkt2tFeqwFuO2ndd14BxO9a
dSbRSc951DNhOY8ADx4qNOIMgyVpP3wzmUdxbwfbaoEbrxi4CnmT/K2hOW0XaNzo
T1P8ao3LahAAIa1glKpLn2guLsi4XlLLSgCcSCC6uGhjPL+9Dbx+iTpmI3IUgA81
q2gpjj1zObAPLB3+6HFpdT78WF2cqkFUXJH8aFMBPZgbcREwLgqKex/CGqJclWz7
ZWwDQZPozCAkeQg4zW7V34FNNn9FjWizyRVL0N3eb1DM7Knx3JCQVxffnP2QRMfK
2kI2b67cjrr6otXpmxy6o8J9MTIv6PvAHdckDUNydHTQYipDyh+jUd5uGxs9suw1
hU/7im969XG1vTwKzvaTh9KMb7jHPTIzco7FWtnpOAAQOj3WwtzcYz78lVoJF/WA
IW1cRjKOv5b59VPWWsoiVdbw/aRyvKwm+QAy0B/T2fWvZ4YjLWnn+Kx3F7I0U+Z0
sGpA3qJ3Zr7wk1QDtf4AD5w10+tg6x2RVZynPXDK4K023ZSnT1H9CQDtmfFg2G4W
fRhzFuw9lxqNSDRRM0+WQgn8sVH+EV6ALlDo3kkKfkI/MwakXYatErT1iqb6RAjB
2HmRR3DSk+03vyCoqU8aMLYowk5HgR4JApsQIfDm0rnDmjokSAFl1zRGoOvg7Ndl
n0YLKpMTxiJ3s1/zpaqIg+GPbBu37fyC0ph1/bI5xKjkmAoVhyYPgtcWC/DzwhJA
NfvgB0rCzp1IMcv/mrrDotbD5/+CJpnoy5Vle5T45B030d3u4yIOeF9E8MYaBQCO
potCUi9jE3j0VfNHQNphsazPvf1oGXyE+G/1FPx4hg5ciBf8v2yWZXk/s6Ih/bfP
vzrRC8ZR+s59VdR20atX7gYPZd8nIJYo4g8/a0ZdV4i8sRP3qLaTlhZDSNeQ1S/U
0YHstiNa86ZGK4KJeVafc/DjZJUSqH4NjMJl9mSX8YDWlmO/sNT5ghufRMugmCvF
Q2Zu4pLmtYchUDcjSUucDspmQE1+/CIg8T3pwpQL/SoUivGNrst3JKCXZsibyeBC
Ad47IjKZ5AS0pUWECURW1KwoYcehK92dWoo7sBW58Kft/T0KG/7HFlAIHWHCRQlO
qoKlmS8/oujqnl4u8NAzJYBDKTDbqytpS//4v2vXF5ia1sfIJuTNCBqrOzTrVWSo
G0D1qRJlL5JHp3WTDSL7PF2guQt2Qxqns6s9rLgnXfkWi5w3KfOzm/jCQgKRhkIK
4/Bpif6mIGPhfdWXwvYgObbvDNVnZhL8Maj8jAYnj3Zk1fT2mOnnGDnHp+9OieQ9
0h3d4yEQnG9yYXV4iFFZEEhdo9Y4QGFJkiWrgk+5GmnZMmWx/72MxM5dgfbd5gHx
92ZuWhSSekUq7TJpR836IiRbrEBIjMmQ250U1Au9HFt5hE9gpD0c3TJlQfGvFyfw
gx8y6r2xPpcs8Zdf/LJK0Stfxiw5s/ElVTsH9BjVsUqkIeZ5ruRf5UPwm9GFMZ2H
r/H1hUzgMBPoBFQOVhUuZwm3fr6ZAu13htePz3JIvj++dvSn/HurN0UZbhMHIA4R
iqBacODocHibaTUDbM8W404w0vgqN1/8/OO15frJCc3TjztDFhnCMDS9hbRrV4zD
1G8/ejEurYSu5iVkyZ/GhE4qkuYsuR0fE16lXUzchxBh1DLGmwMd+7MdMwCzlNOi
MobuIfXOsdTUk5R/E7nZNLkgUfHVk0TMt9gw3Ar7FrFPUDxdmuPH8CpxwD4/obaa
57v+x46o48T2XP2BnuP7mfu9JhDpmspWT2sRbfmFe6f0N+pW9l8emlVhgF0mRchD
aqT35QcF694XCP/a8Zi715uxafEjORf1E+wSz4l8AnPAC7xtLJ9dh9D5TtncMbsk
32m2kSbHIb1+78cP/nI9RRSN+0OCoujVyq0JdxEeMnWVMZFmc2BEb5cGYvG1EiWw
H34WYBL5JSc1809KQJ8boai9VVegheA6QVm/QTvzbZiKHXg/Axk0RCZTs6rOomC4
n4twTgYy/Zp9FE5Eiu/VgL7itaURIy8fuqFm0OCE03Op9/iWAE4Itmbl/nUR73Sh
TpxSdC082a6tGjmU1YTHb62kcjbdTJh7Mb2hqotiR1YTVJzATL6Ak8mTSxiNiKLX
Bgn8HVzpNPUag8Dyzg67vc0z1+O/Lh0SlpbaDbN/lBqKuHY49QbIxv3lDSVkl5+G
wZyk39wiCBDYXZFqxBJWjDTROk03DWOrEtlEU9qG1VAigVNF2T9dsV2UbS3wU+W3
IjF4IJcC9xplFLQe7bVRuFyoqErYl9E2NP9eeIHX7zTLKmd/xt+QgSymvqssq1zp
k3M+ZUAaCzF7HBrMl/rg+8a5gDinw5yGrWtFqQT5WYN4rV01erf5Yy/wsA7C1EG1
vTS89+fPdd+TRSOK0phhMsaCollX1IBHEdffnJbnAIL1DnZrBdgYUp1eRhrYWlIn
nyOYExVmyMOQozk/ylzQ3P4U+113E731No57o6yGF4XrBiZWxPD2qphrB7iUoA6X
t5ooae+4oBTmdDkVRqOhHjRVBYpzoJalNMIaFmni39GbBfQ52OVjIx54wO5NUsO5
/omF/4N8V8KGfyI1ev49a59FhlqthyycZTla914uqyrzzL6yc4cQ3JnlGTqbxdLR
St/cwgfcfBsksDIBC6+qDcxrlao7f3vakgXUKU1vNIwgKa152Ib61/iwGCS97pxi
TWCZh6ZCmBJts0VX+W+W3JBPZ2Su6yioCj0CLG5MbUbOfyoa1Q5HoLGjtNUU5Hp/
JsGqL2FFK+HTq+dxRltmJB35Rz1RSGo6uWXhTEEfub82fyg9iec3hjZ4Joybrg+V
vUmmSGGrpk+5L43/OqI3wFOJCahpJJcso0i6+EgNjfVZIhxO0NlTtiQOy5qlf54c
KKO7G8d230DUPa7roMIlVZlDd9lxSd7svqOkkcHh63cs7YHpEiGCz2DG0zA+xsQb
n1E8QM5cBEVZ0XM3H0r5aP1wd1oe1tgEt1awUzzm9eoQ5dikVlZ1jHhZ2ASV80eZ
xic7urTK8Jbv9OT03vsMcm8FvbGjM0bdvmEMqyc0qAzp3MqS6/Zwx1iE2d1d+KPX
xSsxBeMW+CHqKqCg9W8zDUWAahU/xoRbCNrfN+CZL/RHWrgC76BoCwZ6DF69AatQ
OKWG1eIphGw3cBBR1YwJ675uawBGCBtQeVauO9ty4qLGVH95rqJmVZb4hpzo5sF1
oV4zIbK1gGRQCiTYwxkFo4yn/0GGGjQ9Wi3mykdZgk2igxu+y377ENe61WqIyhGT
hGqeZbCrJAVcqt4OUT4qp3rsTikE78Byb9dA6DIZFcFkDbmUkpuPoKU1wQd8MTeM
oMh8x9Sx/ZDMhNTB7tfOWh5UBefZre2hMR1KYjjCYIA1acdFyGz0Ko7KXNeHKP8h
E7/bkisdu/0wIbQ+sQ6I+rjVGZQhkDPTKTzUijw0nlTPHHZWae5XBAyKeG6WJ6WP
UvutI+qLWB1sRmDp4xBzLIKJ35A/9xLHH+5Gn7oHyRNEtdjhSIpC+qae5GARw2Np
xF3K6TIqsQAr+2zX71zjWItoL3H9hQaHA8+NL2yGPRbMm+CNlTUKdK1qR3l99NuD
NP5TguI2hUVNqZEs04eDBzQH8rT/sYcBmRTM18DYvdpMTUQFxz/Mn/L4qhIPrvgn
W8hPKp2PFYjRiaeCIjKj1KH90jdYJZsPTufW9P9DVTkdt7/DyIOHDWCH+DirFIWS
s69BY6chm7OlZ+NvLGhgKTsutMvDs/t0LW2a1bfaiFOE0wsLVYmISpKwUb2es5g+
+9z2TJkeTNj6ISfprYYmt1MzzjIUmnMHhR5CIhGyYZePt222VumDl0FFQAEWdMGI
RaHraanxmVS8TFRyJop/PtKjcze6yn90IRuL9EGGI7prfvqWzvd1XTdRto8zqEXa
1Rc0moN/ilUjYkDj+AMXpb7mH4wisoNPVHyvkjY3i2puckC5uik3HFJfBhUxFoMV
d0SSSoOv7g5hilUUFdcHH857B5XDbBuJxKdaSrf2vidkqXLRfpaStok6mCgvRu+d
NnPf1E9lC91vrafqSunpR27dUzgxCIf4tNfAWv+DCeydiZPi9/n3xEKzVH1QRLMS
fm46OPuDXkj4sYGAqPF6XcCFTkVpUYmVYjXkcz6WS5u9GYTpWHZus4TQbQq94CQ1
Nlmk4AR+MXtfsqX3KtOQGvd1Zd7RTM35Tc2cyLRv74bCMzskxzmvDHX9eZwY4/5V
OYo/2TpsApcYqD4e/ofD7ceCQkIeZaY71JTNNbOXDttbiSk7/6h5FWvEJlqZ5Ktk
KZCUw+ABBwoZ5e4g14FirVAtOZtnIJ0xMqz1rC0F1Kv9CD3dtcQ/NhMEtJf09r+N
IDMqMZleNmd74NKmjEnzMaVfDhw2cCcwBby2A6qVa8AOnU2WylN99q6bByWyeH/a
gMCl3GYW/iLje3KFBa7GdkOIB+6zTk7kg++u7qHMoYs6qJDfFRcyijm4NMT0/eRb
QHgGtAIUfRhwkRshE9/qaAdrW1p+Zny4lWB6ztpe4eTwDcbRzmyKeAWdCmo4exoA
hLoyvW7pyHSD3Z+wqu8zE6F1OJ4nKgy/mxkT0JZn79UlmqfeZ7X2nT3COFoPR7Hb
M++xtDoc7cIcCBYPzyFeC/hn4lW4giEATgmM9vm7FfCX/VT6NvtyNLpNegxetdIj
oL4pHwMFHfF+tmZJwUNFAEzuGgamHA1pRQV8+TorOR6GxIEEwSaYQCjl13QoaKey
0ouKnwavIMFUmtVWAvgX81vjdOboQSsuiv5sOW0AL6g4xKfNNP3B4MFfyzomhiyF
KT9xclA+TZAUORRFjz2Jm75cif9PXvSokF690N5Y8CocJtgRZ4OpbQD74dFAQRcI
WtxIPoSF12cuc8LTXmMuYfzH0GKeMb+uzCAZgfZbGMnXP8JqQb+tUh3xeFet8PHO
pHIV5U3WzQRK8aaSD0vWBMsy5aVu207KI8Mj/A2mWSjFKUD1ovvzu33tji1nuV28
xwlqsgoCWJpOWOb3MxXxsRHKokH6IXAiWAbE60pHbUc0L+khD2r+cGHX/Joo2+oO
yu4PW/syGQbTj+ZSn3r9JRJAL+YzVAyysdBdcBw79zntFRglvQAvUtqbFb9ommKq
NSwZw/Q6pTBxqwA0q0HE4r+I8RbTZOIPwvpfQVZ5hscj8RmgJMB1OkyCOX47leGe
A6ZZgqpBDKwTq/xbB59uBiAU1UWzUItCzIo8mRPn9ndyWwFpwuiby9YQG604j0gQ
w3u0wH21aCTikN2A68TEbww2ObK3gilfIey8PtyEkZczTWpWuHmOxjZHqDTwvyym
PY9LvaPIvkNALbb8E4m4acofex9qBnLyKBzP94ZYJypjN3RSS+9plSSSznwKEmXv
u4HBTOySL4vIzuZf6cvQvLfBKwOCEZ2XsFqLp/6SpAKxE8dAdrSyg45oouqcgkog
X5DRsbjiOhAKRS0+6kYeF4Rr8xluYz+qLOd4+qCUDrBwC1j80Bv4FkiFny1AMUnY
7w2VnDcfy/TS9D+b5Sp3BuTNP3OcLl/zfjdSTC2Al//2odlnwJvxIOxgtwG2+A8E
FZkB+HEwW+4zCsoyjyTrAW7wTRP9BCA5cqpG5DoLnZTGqxCJwTjZanW2333Ilb+m
a8GM3YJKTJSMYVmTimJYY+GyoDSL5ISEvHcOzQ+KXiWYHbvVjZyCHv4rz9C+qNQA
0a2Ww80VTPt8S6gNRp+ObL75MYSUlXA5P4nYwrYvJSqBxgd4DHhyNJioFFbEotLq
548LKKFjf8WdSmyVojUuOcscUOeTpcToBOgPcZRaKFkFZJ7OvG31eUBxn1yvJ4x1
i1GhizTO0MIVSWhsl28riPRRdm5dsn2IuS6ueF5tie7IGhAZwHJ9wqRj7SY01YXu
gecXQF3xqGOk0bTzYshoH64bsrlzSSzhnhTFLElInENKOA+gSRhgxGMr3hAGXTg2
JXPzIBOPPZl9gNU+ZZDmY7WwNzyhBgiGOkHY5h4H77nqNrXIa3D2L6IQToDYmHrw
lWI99AE6m2mO07f/WertcKvrS1iKlajrNCWZ4BZyCRaduytkbwS1ApM1tIvfWfUn
fEQA4gTFDw5pt/qbvBbpqp5TvtHFI8ZzfEX+v/HOcWMgks2UOSylZ8SoMNnRWKv0
W2d+s3JQvt2ejBWfK9vmpdchvBm5Ywx3LYMhgNXdxBoupEWl2dttwN0ej+2a1sp6
UdUiBStVi6ZhAXtM/3ssHS5uVzy4FDHFPmNYVUkcgcb+YA1fj4IErWVLGRg5EUKb
u4/souzMEGZsTBvKqixjk2nNfa7jFookpNblWAMGgUHbJpaY/i1gxfP2j2nSDvzt
meI+OUPbilyLpuTRhMm/b5nsTx4Sl99ZCdtlf7pk7MFhEZGc9EZfIY8+C7tptAEw
qnM6Hot2TsR1sOqCXG8g6F3O1zN3BoN4+stiLJxlfNJLzz5O/KeymFUqfyvFEkC5
H4AcjIx96++uCT1E1jmWaEIGzVhujbNFmFfDUwG0nPlFMxH2ZAjLk85pBdxqIYcp
0yoX7ui6QfwkhvS8QlHK28Y+OxkNHsNvrH0EKbt77LMKC3ol1zoXd8XSZ0k+uW1q
tzPfbFpkHtWARRcEyLUC89MUcWzkJbO5DCF8SUaBKYOkXAF6hmxbJrOoGHv4GSXW
Hdvt8AAQuXvo/U86YKF0R6gTpb84WP+EtwFiaqXj+Nd/Jrk2aisdyP/ff+VZREJE
iZv4vQ0PnvTte3FVd6ksGTH3S3T9oGadvW8e9se/i3OhbsHmW9Xtopsb9qzdnFfk
O73DY7pKTZoatpIjN4X7gNmgv5G7/GVrfb+hhNAQ6k9Kczs0TLx+l2+gvL7geM1W
CQJgW+5H9Lf1JSTh67SGGS3duXzzK4/DDAa2T9RdSS+wAY7WXgkbyGpvxafB6Nk1
LVjhF8U5GBt55e6YIm8t683RHlizeiuIVP+p6S/jKjMLqF750gL8Rtu4jh195NfT
eO/dFmUSvqKw0tULt2pjcIGvWt1tjew6gh4YfyD1iyz8wzXJAsUM35RTXseEtcGf
7T5FrrU8M3QtpDoJCx3Kk4kynhp8Wqvx56u4uQY8QwkoEFAJv70vkdINfx5f+RsY
2LltcRsBXrezgLrkdrkRRYpGB4poBApk54qd3Qz+nSiBGSd1V6L/0oAFZwJJ9rX6
NTUfuPmu96x0Nql5kNYKgD1T44shvK+X8hF1GT4+wtVbNJKeUF+06WXLKUEvRiU9
EQuumuiBilIuFvRnWnb0AFfhn1/Lftrp91k1e69doVm/Sc5MN3LRXNAhQGZRTb58
/SjaWXupxBGz8wAn1PBxsIbIvGkADov1rucge9UItxoAa5iWVBtpeqLfs5AxjysB
SAA5GoTChqpk2ZGZqaeYrWu//H6Znh3KP1eJvI0d4uTSmFklBkSHvW3ZNyLdN06a
lbz2lKrFQaX1T35R2eVqAwO5M8phbzVEMM3zh6zBNkW6Auiw3/qTpdFIXQafx7jS
BzGllXUpZ3yLoU5puGdB5DhVdyv61mP4NL0Cq/FIDHIyuR8xzAzHeitpGz7x+HBN
cGX8pJSwaR/13XAfEG+POACexxXMSxlzC58E8XH2LLajhBgySYwJuFsyEqoyy4VI
O3knWGfEHJOqub05u1jD/FGU7owfgE66Nr+j095nj6hqW1mUNTBimSFvjyD9kS0p
4qdwiaUj99Bj87/+GP63gK0Z89jcM+Wr52H6Vc8FCiy9tru/dojyUDnRG3qQT0Uv
VCgLVin9unBEHgFAzJwhXQHqHlkg6Ym3ayTJ6OZUBocqNcHzqijvDWBZ23VLPi5l
6OSs80ehZTuEYwbDu/QA8Sydy6EZZakkj9Ims2IlHXD94Ys1CAQsMCvNVBfEs73k
DIB3pbAl1L+ZkZPqWKd5tlJPAcydykoCMA+Q0HANQOtiy+7c8fCv9jyFre1+5DRR
kY7ofBBeyW1X9N5WIm1fIHPeP0fS7zLm9D5SSVafonJlV8N88Jc94vWnEAVeSp+2
DaNFyql/hfziG5iG+4/nl5JvCp1E1OPunAWj1YVDZ16AnandUgv8RdCIwM5yeQ/u
8pzbhJ8x3s6EcKyD2Es9MKciiOjc7PnSfRJTI0/I9zgsPlyJ0HS+BZ+LSsyJsqjx
zXfhlS6NLQUWOz0TO7/SeWw8jptl2qt7OIwMtxaq4VWadyt+707GbTAXvPf6fP9m
xUzEfYEWsjDnU0c2wgWiXFW9wTX2SyzLRbdmG7OUBqodYccGPEu29SxLA/zhhyRo
WBb5/6PRDi6netVoW8NC439xXodidh2FtUMFyRFGf31Tb46JsS2oOG9vLfK/Ct3Y
6+dWjahHmAd6+xJhOHvynU4jiKAjx43E+h+cjcLo5dLL6/1APqPu4jqGd8fBL/c3
LSpVIrS4PGqM6DHRpAaYKXss+49xK/YLTXLEsfN1+uMfHeSqESo3tTtmIlEWsOUn
+3L1SS0NnXQqd4ElP0QVYxwuPmTV7fpt1qMkqJBZdCdqXYXp/M9rDowPMmihgBsj
GU8LBIEH8MHYg+3/o7CEr++LmOpEpOWHz48kHxDoU79Gus9LeD2Co99SCL7PxXNc
3uxXwBZfsvKBYNOGplsctYneAN7CWghJWa6ktQdAWrJePc/rEO1ehHZSmsVx50HD
4aaI8jYjlD4hZgP7Z0iZf7gHYRwAKHZ6rTcvU2S5vkG/S/1UfUK2q0udnDC8Ta7l
TI5XBrybEWMOOTf2rYBtkn8wpRyIY33s0zxe5UZrMYl7RLDGhcK0r4yEWdWdHoCW
zpc2ayNX1if0VbZ5QRcALBczDo3HybY5juJV0ZtyvPa8TTFQXHN8zVNnxtrz63XW
sXrb6Pi9Iv7tCl9HDrblWszp582v0KQmmOlsUg/3wD4LSuQ/SiD7+ZamEvFMzeJF
hp5muMyXUcSbiyuoCNs4wH0KSyv6wmrZMzxGJGAciQTLrK0uqLRv3A+L/VcwKd1l
Lp1fyM5sdevwlbi+BgDoUV+z5QwAY0VDcq0wMYxlhRDbAi+AdrFG0TSWgA8BP0/T
kF7VVXzLEcX03edTNrK5/yGWpgmAowcpeInaqL368/69JPAfhclYw4KOdcqamYjH
WORCrqLbIP+yIg1xieEJhWAwNKVWmIrnRAUvnAU/D/MD8JmG138uED6NIsl8DJhR
G4FJsfht2UKuPJ7uAlQxo8iNZVOEkjU4pLvs/TEZFQjC9W+ysf5hTGPPmI+WWZ5O
HSya2P59r28p/GABJKyu503PoFSSJUUg3Lw1DzrOebJhLbp1I6c+kl9dmATWSZXI
5htu3ZjkrXM87lRdf0GUlkX+GZT3dsUjkPlHyp4UvbSRDVVaXq8uzEBw6MYgO41o
vaj32h1NqudJKyUDxQm4E80H9cAmeoXasvjMUySvdsMd6KXbOGN96Kry7GpuGCKL
f1m7xB0lnGGO0f6TPJXTzDW2+P6pBmNDRVVqmr1mHzvVIJrdfdvIN4KmDJkqY8Rh
p829NlhuxbRKUQrUg+GLxrkGaB3v8gWB3LaDIxSj9gDYPpL4YmjvdxNjmwcPNmyS
nMTfysVUHSmO75SnQGmdtw6XaqGh1UJau9dzPFueBvZpv7E1ntPihL5SOXZhDwwK
5UgpOJlSar1ZnlBEoP/tIBcuR8qBAnfGtTRr552+2hK3Q6Yuz8ChwLj8Sg+UWuiz
M4cENvvBOv17xVOVKLQZIeMBpnDHowKtZnE9xEwDcgxIFL7XUManeAirDy3cDhRS
YcLUhHcHfCdkQDu80vBUz21rBQDLnHIyY/YUR12BPGVbKFmxvkc5iaVFrZV3B65H
pcQSTKU6fDDXQ2GIho3K5M0UFraV4v+6LeEFgsB+9hK6hQKZajKEgLV1+7DJwG5X
Cnkx2lQYrDQ475eO0DghvI0IYPcjUAd/G0N87DaQBcJwfVwnOHc2ZENcN88THwTF
z3ShCAC6WzbCV7qJfHoQ7KkE1HXySJLK+IwHXTPF5ltBnS3b3l+Ts1cEO6tgKE0U
ePQtxUr8WoIHzu9yhMQp3KSsXHZZAR/IQuzOLtulC/lv3U6KKaOVSVjQU9+i4Cxk
YxgfK0zgPAC2BTYj0vrAWaspa2Y2PuFpCFL4LeUJ1NptNtWANd9ZzExCYxXW/PKz
CN+2PCMS+W5Bcm+r92wQ/B3hbRnVliZQWrVRwNXB2YTwReyRdias3bcLWjSvcfuI
P6x4rTCcyL/GzCvbHYfqXFgIZZymJfiKRkfJM4OPe9KqKCK1a8C/QXiWe+rAcABi
20kNGaHeIbBMuHcEHRsj2fBl41gbRLX4fVcZIGQx5vSRHXatSx2PMDPi5aTjh3Nv
aNtQ1+sQ4cfCNzM3O2A/ujym50pb2J3Qsya+PBdcunH3SqZ9Yh3xx+U8tEK4jI8Z
CVyWL5ufuOavRk4uLfeZQwealHIY+BUvIJOFGHcyt3yyn+d4tVEsSHIyaCy0WMHo
4OrCGHCOO+YL+Q9s0vRz0bXSrhay5BqO1vl6UKout3AzY6zMb6LGUICHxYL4tUUd
u4KvzJ/4r55FAyed9FmsUvVOqfFsmhVg6jbQBCIATfTQ3OzpRVaxBiOj59KUZrdZ
8ZRl6rHUWObXqyUSYEMoQ/0jMpRLHiIZFb1yfVg6rl8sm6OJ+K70oD1idSJyk5ch
U91mABMPhFSLyEm3AmfmQA08P1mXfsKAZWpGFQ2MN1r1DyFH+JeeFpIeol5i3YDt
+CcugEV52s+rfSiHWPcALUN3XcHmcRJXGY19XjZjbNcojHLOYHpE3oJVuGBv3+sp
gSrExZjnUI53uhJEU/Ins/Y+U3oJnu2mvOz/hPb+z7usthmdbKAnSzOmRcecTZ64
b4L7MCasyS7bHgfTPl8/TRHx6w++tTbcTNTJwTzCd8FBEz+oQaYBLDHAHz6gjLWf
hgTwDZvwEDLSXw5GxR6ppNmdJUjhHJjDPRcvczkwZ0UCDf1hGjbN5hOSvzi0OkSp
Z6UrnfVvld/mH6DbkydipZF4PYmfPrXRurhgzlBxZzVe7MrirRbOu9datQtK8pAF
2bQlytkMDfZHq7IjVSQqes2kMYKcUpE5yRn8Dws4Wz+reH3LZWw7xppD/rHmENFf
n9J2IvGu/U9yiaiZ9H+u1zQ8/Q4tCWdjFANvqHOuUVfTO2c0bS8NgBIMotsqPgu6
2Po7lKnXIAk8XV3EjsSMLK1AAnQW2VWskCcWzRsI7mh32HVgb6t9M8n40IZ8zGap
qf0tUlE1lmeoWUDjT2QCSFpEydnDbL+mClMjBc3oZGKS+1iwiJjDGDGiJVDYjgH2
wpEBqfwe9QP5zX2dHt8TQ18XhBODLsW5kMFlirE64ePxlC7JJCto0CRFOxxZD6tu
vqUaSAxbd7kBnVpmylss7NpqwAXB55JHbd2ipaqFn8j9oj4KZ2E9riWyQ2Yp6/i4
ZylrXoL5JjU0uZABXf/ztVxaq2C8nLw1UVbToDMTjeUrxDWiBjaY8HFQmU9uxDz+
R/WleC9tQDvFLZfUhvFyC+NHNJw5E9/wklBqIA5m7dqn94AVbdVghsdAF+LNLSCJ
7RWSYM50y7Y/cwSk5Cyjk5QnKEQdH6Xym11Al6sHp+7V4Rbwwv4HrGMAqL4Gtyj5
yYU8pwcVTdNU1b08PpU3SrnewBqvESAR51fSI8CgWRf1RHjyEBnpHMwP4EE2bBxT
0522HnTLToYiCffvv2X0AhUKts4kshHLraUrwTbpvaOonKsmFitix9e0tiBuYaT2
BQ3UMHKrDUrF7eLg4uIsGA8HmrrW45S5BQQX9ZvZFgc8UYq8tIBn5ZDPz3Y8M+Lo
uKNa/cl7Lykd/ewZHA6W2jNrczVVEiquWVOIUhcadvRi8VO0TZhccS7e5JlPrzw7
w9QhFI1dZk/0tNMlGPRNNW2FKNyklvCGbMtdocuyoX1FopCQM/k8lT7iD0jHV7pz
GDWj6NG/wgbx29VXSPrFcfPIdWwrwtfYKqfVCGOOT3AAwWYGkgg5iMYChX13HZb4
BP3yrEY14yg5XjiiB7HYjMVSdshDHkZUvyIs78EiVCsJ8osBNXfKMAJ6Y1H7mi3N
Ymft+vKNlp9SXAlgkYB58hmDEC8U+fewb1vbvVDSsn78d+MJBC9Q8Q9uqjzavwlA
9S/M+ZGNQ96/FMkfg/F+kFSNGNo4DTcLjb1r4x78d4tf7Z6P46Ts2bmI3MrGzYlH
hkijiraUEQtuLy096LUjSFnUQVqpFKg03Rphqb3xiUetOd1NKsUH19KtnkI3dwmy
3jd8GcTEzrM5Mn5mmBNYckshfrzUA8I9Lsgesdlp0kvBYChslIuAxq33coqDww8M
V+BcIYhD4PJeppWtD+U3FPr/j74jmLnexqY26hcJRSnqLZgyc2aoe4PZ0HkVNH7F
ECxZUO3pIjLVb96hEZu3S9VGHcY5N6JIR7x042QoBbOAWg60Kcl+OAJSWTV4ZPUn
zdbag071HGsNFNl9d6tRk6BXUdt4vdfjzIxnW3D47z+rpmsIiyEChTObX33ZsCbW
St3uJA9sudpg+mf3ie5K15i81yZyW2GgEHljCDyzc2+xLaKsPcrB8sGJvbyw2Ge+
AA37oZp36wRUT/XxkhZgX5KEXV1HwUxsgmxxNcU7LfGvCMJn6W4FSAUcYU1B3ODu
VGz0+cM+aFWGoFjuaxF4ctSF4fjTgMb1ub9MH/POFIdzY5yNqL8Ze2ndoeKIWbHx
SeFpyjS9O5j78NeGjkU77uIwgGdbrmY2leVwd/ZeygqIdOv/csOd+t58LQTx2xsN
9xf93GqI4pPPE9czMfeowMj2R5DQlRw1idZCfA2dD2ERk+165wCwk7qrv+FIRDsT
ppKm5GdMY7sv9scJBqwBAJNNOVsVC3AvNzWM/74Lr8zZWcvEjt3vLyZJyfchgnpn
j7pWqniWzOccu6T+IpEiIovFwUEG4C1+boeSQGZmt08Fmn8Dx0dGalCbEWy8o1eN
hGQLcOgcNqHO/tRhCl3GalbVyQlgc/Hz/51XGYdQXhXh2hjy98iE4hc/AMyNAtP2
27mO5QBQqRNXqYDnnwwoqy4m62/agRL7ue3DUL+QA98zbNPJsty4gDAxMF2Ib8hP
a5SdLT5uZcIw94p3voWlfdXw0OcP84VHsN7tLdYD/zyx2mm1wczaZdNkrKJBZY9S
QFrOjpyCbdc/nklbvBM8Zb/fmhsybt0phtxn9xREj8Jk3tRDv39XwCpt+3/C91IU
BF4kulEYJKIBOAZhyh/dmR1lO2GidRpDzD2C0i6Ug7KOSnY9rKkIK3N2nNc5ltZV
Gr1Ep0+IjXQKdH15NnlHhPde/yJl0T955Me6WZW98QHC8jb3qo6rwrtHP2WCepiW
1anh5mvXerWUgK+YBGbpCRFSc6fTOdi0H7a3uwfn45FaGXzumTzctTV3oeAUXKu+
ctmR8hgqHILoywnHvfUNZB5iUTIgZpCj8MBpkmfQ0zxIeujU4yUDUmRWGXdPUiAv
zv8kYkaULFWLvTR2Dbf+eWluqsXqw9QdOa3s8xpSyX3TLKuwnUjcPONudLVcICwr
iuZLODpznZiSz7XpWX25LquiTRptWH6VKPE17xslGfzVsqobp/HH1BxIPe8tjsUr
+EMWEHEDwYOEZycNvqk+NYuWMTddarVRvb4jpwMRaLm8/9C3wZArTVXEmWnYdK8J
Rr0uLpSR9Hwb1gMV1UaSGDKtjBgn5WKBM9ejBOHt7+PS89FU9Ej8QNBe+9zR6QX/
pS5X3DZzngmDswKDqBww0YwDUhZpOv4GIMxYjl1MmuDEvi+IHnw+0yHfNFSJrZ38
IiEJbrH1af3K/rHb9QdrMQV5n8SQFMEVvTizo7f4YJznOVD0MCxW0miXWr7eZAoR
smjvcFKodK6PKZG0xMq8Z0AspLzbRJ/RWvr0EF1pZ7QEsMZ8KA8UE1uwHNlamq2S
ke/iu9SPK2cXIkA2Uh2w+hOGsTjtObV3jKqYIC2Loa2WxKgSyL9BMrkSoYBQY19K
ANLfx4ZoP3IReVBvtyx1n5lhfA3HYjq42y/mPICIIhjJm5bc6BhRMk+x+r0YHnei
oR1ui2mZj629oWZBhrhEk/0BOlctzaAT7KTUXHqfF/9f6WlQy4sHm5aW0+A/62v4
06O8lazZ2TuJy6tLClinEwh432CIFeJWwg4ou+44Rnpi8Q6VyCw11UyY80oDsZDR
GWPZBw1d9g6oqjsEKYxkWc98ljxJr8Khi4mycflR15WuHkzaJehLYejVfDrMNDAQ
2yJywbH+l7nNpjhZM2hWzK0o4GEb/I84HI6Pj2fT4tQWLlAKQaRQZSVIHdjFcZ+K
Y1XiqEveB1JCYvXPzLK5sCg47XAG6lCNBENERfc8VFBU8rwIWeoz3hvsQA4anvl5
1YHajK4XFB/PYlr6Oc4LlBh+J0RVY+xK4Qa4TQGETIoNQvJLV3w0W9cL+n2s9mZT
5RHmDQqVa8auCgXM0GjSASd2TAmk6+Sx/jlpWdF5IMOezqI6K3xPevIkxwmkkFYD
wt3AML+UeLej9B6rlXz/40ZktAKSokArwxg5+ffWTVxLgJUYm7GYRMB/oN+pdkss
Nt8Eo9bP3G4cBrOBUB4P1ZVL44bceUyQGAWSam/s5zEpOIE5FerCtr/jZ0holdhV
fFsRGTTgv+LQZAnmNcIaoqf7ziJ6FF9BhplfMS3aRAK+2bGJ/AIkMwm0XWxUGKlI
OQL2wgbXLL8BlfqANYOfNnt2jvjK9yDPIAb0WfQxSYp3jmvFTF2rX35UQil3GAxI
0HS4b+aUg8dvSF8xD/xkEuhsARA90NsS2s8jXvV93o3bbqY4ODDrcFB7BdZlOLCY
pyvPTVwXLUsrXaqsTwe9zAoobrNqr3ubUBy4LTMZYk9TQ102zn+WS45yJvfgiG2Y
22eXaahGhlMve/kX5fqu21McIVDIHAUoL2p9aq8TNBzwZGK7fEtRqQAwp76bgDh1
s1mb2w+tc4qSpDuYEKNWcRfnk9w7dqCjMPVZAbOKJROs53KKQtz7jHocwnFibESc
+nUI+YJu7APLzM7psMrHRA2p2VtoYEYpB31mzFeN9QkA5lES7yBUkUxWm3w55jhh
emE4xOvEcrs7/5wETJsPdOAOeJOuzkLbQnHcSq/lrEbeRPqPSvXaI0/v8/2vdmPB
lMM2YfxnFCtcZDacyobz2YH8G4bQWzM6UrnaVLV1TeK24/kf4RpVv9jgIK4ZKgeI
PoDC70EKdwRRHS8WtVZ/dkVtjpdOZYGtR3GDBQL7b0szoupHMO3f/7deQkEK+T1n
2Sa6vh9JtrykUD4nkdyTJ1SFwniSHYf8EWbW4FnwALp1gE6cIuTmAhoDTrV8Zjmd
Jp5/gapM1nij68PQsOl7QRco1CqKCsp+tUtVmIT5wwF2Bfm9Cbgaw5dgqirWf1VR
Gdt2tGOt3JM2yiwOws7nAmOJoWDpbpHr4y2/zAoqBqc6v6bhsv4DEN/io998maUu
RquQDhbuE3XkkAdxnXdBHMGGVZF6Nf7wDUrLTYmq1jJE9kQ1QurdymdAT3zweOTH
Re0jk5+0CFgiNmA4gDOMtXcIlY+bNvdTpY8ckmK0j6uT6uccpeINXmFrKtgv2rKo
hLXtowvDE92z7/QZh2AQlkQkmpToNx/H9ZxHkgAUu9wokF4YuEXKgmvSbRnPrQhx
XrtrMaJPw8WgZP7ute8AwoMBUciDJkwfJK4M4MSRkKVsh4gRGrND5KqfGpJp6cXQ
14M/NQgA1gfXR/b0Rtv+N7tHodTG8jXBUL60yGqShzSd6HOVFczOvnBfE5x8HbA6
Ri6iuGP1uH0pXUSAwMjqTtxe2YXwRJZOCI1rN67PcHYa41x5e9gVzX7JyK4FhzJR
e4vHzylX/J3UTezU6RVfnymJHY+sN1PtYoo2GT/fHxtTgXpjouu+5JpyWlluRejI
jRDQseP/NVVHr492Y8BNeBCdUemS2vn69t+IO8dv+A0WTJ4iIWgFDPZT4UtH2wWw
2L7M1ccssovFnVqWSZX9qMAYi9upgs9hwU9/c1I3OiNaw8nllzqGVcuVxbIxVjWE
YrHuyk32YTFPy2xAu90h2HCWqYzToueI7c1P+QixVVAWL8KDA5TG3UUR3VDPDHxi
a59qHubuwKxwNAcfHD2evc0XRN6YW1C868umoSQ2smCgXtVagqOfgF1LsRoKkPqF
WGutFkO3LNVPMNBo1V/o+SWLKuuqBRaxLNi3oYCmLFmfj92nGHyg366gbnBcghVL
M3+mPP6TLtUuJgqTSJyzXO152MmmcTcI7T0THJjaFFY3N5a8A5faZJRTCVSDLaTV
2OhPbhHQEbEbttQdDCTiRcsEXbxHYAl9pukvf4CHE/gw2ZicNxCdIShbuvMlTJZ0
y5XzBu48VcUfZ+KyRfQLSkNJT2Jw7fXZkHvcSLE1D0Fl7GCjhtreVpND7bjo0Cbi
CJBzcysTrgt/2YZs/fiMyp4QEGNQS/1qG/uHC2xshlELTAnIqjaOkm9wOlMJEk84
JkZ+QuM2Dsxt1tEo/fIHbJGwbGK5c4qY7tajZimSTnlHj6MPLqmFXiWpcdM3Ac+I
c++sAfz3qoLHv7D7Z0AzCRmRAiuIwPMI12cgyCyA6N7zGqWyqfhZLPBNolCYsCGJ
QOLqzv5Stn1qWHhHp2LtySMbpqKed4ac4+ZKD8/Z7Sp7vC84cb6N3EeBj9fcm2E0
Mi6b9Q68rbf1mpqRcJ3brGDZcoouP6rJyqiSMpXUgU7qRWSVRyb6Ddm2ivl8M8qC
Ou3wsY+BMe/WXSj+1fM1lHzhs9x6rAVGO07btxPlrU6lXDhridfNYVmcWs6MZwto
y2lYB42GrO4p9ZdYHOGDGIjv/04lluWufwr3DSnLfEnlcq30742EZ9I5Xmw6cSOY
9WObE4mVorDFYkQcfISoNDDf+x8SspD+sZlHIg54fMK2aj3y12pkG1tDvX2ZySbW
Qf/MO3vHcY8wCGcSZGfzEuGj2G9AKJsMMt8ZvjivMpjZbMJ/XrjrCXuFNmznKd6v
Kx425/r3BFz9v5xoTmdpQH4hIUXUc6YhtojolTVr9QJiwm6XFc+fYlEoxqCDNbkb
yH+ykGh+mOMig+muLimaODzlKgSoSUtSFvtqEI+aR9YryaZqNMY3MEFBnVoDp04S
W/77PoSScbO1V0CjjkZrGv5s/WiAe89qsQe9U0BYVpA8gPLmHsoLODG6XM18uvXg
YrNz2FW7qqDx5XptYgnIXBvpe4Anu1DxrQoeCcEP1wt4ewTANClMBQ6fQmqaq2GF
TOi1/z6ZsoNsiKvaMj1odM+48ic365Aa81JVfb4KnEBYwD8ndpc0wfYo0w83aWui
rKE6Cj+8ScUE+ONNd/eF0hWhHjFFu4asW1Zj5I7QVlmcSW1fk7uvdpesds4zyGVM
d6jsAXlN05fS5UntYODtkcSYFTXKDLaRpd/2PKPbzCZNSHkSR0ZtNmIJeUmKRJ3o
HAnqclBzw8B2MjSwzbmbgL3FG6Ftaoz/ngTluIbpph9ew+kICz5Sjj1ib51vMml1
j80kpvSAJXKOZ31nQW8O1pzvGFzwJIbkmnu7F0JujmIiaKo7jU61uAPJ9BpZ2Xwx
zNxbhZkupnG/GoqQ4bY9owqVbNA6Viz9rb+O9nfERfqEYdoYYAvykCUahiKEJjl1
UuWc9Qe2PCV3QZ/57NeYpe4hifhysRuqKNdLoqinXnEOW0gBeiKAe1EykJzhkLGX
UOgHKz4og3CJNWw4qd0Jn1wYAPpUtVfxjs6pOQUDebjwIuJLzfcaKGIw8pJWLej9
shKfMTOGmiYEC9dcioOYMTNlbvwPgbOhuGyhO4y5xRoqa44FlcutBaEdJZ6XI7VO
uCura13Wb34QkrVHp6DxnOL/0jd9T6gJCy5AY2UG92CCvYFdzzzr3QiaD7nOoA3H
PMCAViLI7QY6WUzTY4r5puuCnLLeObDMn5U4SYBt7PyNgK6r/kVVKokec0JrQw2b
3H3K4b9Ni9Hrp5WErxDTAnC7sqgxz4COgG3CtEegU8x2hxZgSKCXArspGkWiahSM
ed6nmwK6spE0TpNFzqCrpyTAZlDMN4hC+LjDofQAAEpxlqyYg7cO5Ubk53nP3MQy
lUl14mniT1SlQnHL9YJ8bIxD8+NvJ1GVgggy6hclTLFi8MR0CqXEXKagEUd5IZrX
fpTV2mEDgVsnwKjVdlvf4QuBSgk5AGO+JbGBFBO7jdwJJq4odqMhOPBkfV+0zZTk
W3ll8LZfNXOG+uSPyoE5INUKqPMxns2VB9P/kRY75B8TDjYkqrhCtYu/qNsvCU4d
H3FPGHRySLI23jBYEHpJmtXZY4pDI6902GnaRdwUTJDvuer9RzHnLP+qrmEvqgog
UYUUF2a5aWZGKQDK+nMcjXGKuxxf6VLDP7/lyJ21ZPg2/9wUEYRHKUuKnbfX/wjU
6M+Th4fzixAhBnCzCzfKUkxzwcaaV8VEzgrRmAzDasyScs8YM/NV7E+YvFecnR0Y
pWxF6Q9TmwRAIteeBIWwWvecASNlPn8SeBWdZ+lE/Geyf7jx4z0RqE06ey1oquIx
aVwvfwNthzYl6RnwehrgBRBvzZzHgf5sN11HNzmpHNwFY0gpW5UfCmoaKPQEkXHS
ia9navtHG3WQHDnVdnGrAt5BoMrQT7y7xbmZbeACTa+MN1VcG7X5TJUW+mZQCrQ9
ruCxu847T6i1bdTWjOAH3HVgdeBmtnG3KEn2Y/AP+z2sS3LBbIoFgMUY1L0gC2PU
Ij1YvSHDBc4Odlei0Zx7flNohovS1xfhBI8EsHqgY8HstzipP2+Dw7NeJbQDpwYl
rT3n83MgwYo2CXYcpsa22OLl8AFctDevu5DIldsKDLMVXD9opUlgGlC6cm7/Zvhj
hIPYn2yf/MzZ1RDBdhMlZA7OaXGYbNMxFsEILIPm4IRKQZDNwLx1wzt5SiXuyP/B
DSOT+F/feaoqt8HzOlG/nmU/ADIYcSXbHJoaF76TT5NmS3qJMioYH+u6g4QyS+gS
6l/GotVLxKbp8kwUpuvIQ0L/WOHD2X3UqTEzGhOpF05sU5ryYrEpMkq/+Z9x5RNt
rnPw4Pg1c8tIPXs0MzshXKReKfCRIUcGjdK9hV5OxfMVWNmFa0fohjCVwd4irYPi
DXkNHXzY3X0wL5Fp2LsCwzw9b2qm2xP+eVApo+nP5mMKqJ31DNnpF4i0/kGTVa2J
rwuwvOW9R9AjM0q4lfol4KHQhXuMeusLfY+zLWOEp1uf3d1j6fonNR4NhuPnC84O
8qNPdPq6Mdtvu0LtWnP0XVly58HWrYFVY5fJB9OIxAMGVL6ySdvnZNVhPwdOufDl
ylppntsyTiotHMYrW3CE3hN+HPLkQFMSavTMdys4auLvChPe7iKuNCd7Qmh5HUpH
EppeU0pL8l+fyKsj2NQXlHiofrRHnXL0ALDAEFXoRWliNZWixa4EUMBnTJ+Z3Sxn
QMpTJe4WiD8e09txwAUiU3S55zLwOTWkQBIIKMnk8fgBAbcTW9f4x12yXptLJvRI
yHfIGCz8TnEwJepIvBft7S7dXaHFSSBTBER4GhJ7l3ZFdxK3ePQMcQb35MXnRvG6
xHpnHVpB7+PQosmaQHHBFK53OK7b8yUkH3pqtj1BRC1sF6ob2uPjNU6lD3beEuTI
XaOSM5vA4BDWYopcKCMkbR9rh6iYRyoRLlrW3BTrk+aLNbFV7/ahQkJjCIppINFA
aX9ZtEzvBddQp/ZLrK9Lkuui0aSzz0imox3FQTkV030zkheJedoFWTa+1Ut19lys
XLSrpI+5NDUt9RElbjQKdlTpRt8PiYxXTt4WkvglQ+Qy4dC5DmbM2TQFMxAR1LIq
JCvdqRta8Ceyoq7gfN+GdV2/kSIhr9JDKWxEcvTfH3ozBu+AORifAfJuF5tSX0VP
tz+P+jhWmPw5n/teW4SKoO4bxN9uOIac+ZWzgmDFt+/YOuxlChuwGByUzNzrZJQF
az3xFzvxb4ImwV1bCPduFdAcDkfz+ZJ5JLrQXGYhKn1WPgufikUsLVNATctWuLHn
GfsyVYtdtVpHR5+pfWVVqec3DNdIjbb1wQBTptnPUfQVTaWlTlEh5QfErW/DpAiB
sqMJbuyxBLmUJpT2W4jhumsCZ+GTnuCFelZAYSZhYB5IT3Qkfn7UPR3sc3AmvZB1
I3jn8pWvwtk/5WK1kHupOkBqfl3SRy9bbR6pwuzAt+ldgrt7Fni3jgcZvmUnPQQ5
My6EOT7dBZloQQIWypnRJV/Nlo8TNtsHbHbo5VmAnPHNxsgGiK6Jd/zvL7lPRYim
ats/jaMLPDnD36C/vQAwR3PFiL+9ej+jH1Gcm+aotX7u6cfHD1SGS9U8t8W9oF7z
gB8VcjAIDJ0LYjStaadlUeGCJHgE2FhVwQCPsyeZ3oDXaAWrVTJblOarqxhVHVDa
BHjN3KokN3wExYXamVh5hzWJn7bW9lrO2NKuZC7ij9tQt1LTHrcqANQ9tAuJV1tw
RHzEckL6Ywyq+qZZ5MtPclSuOYdjbUTlYfFQIRm6y2LSX6iMJ0c+WD6205yGFejn
qnVNmPm5rzscbr6x1AEbZp5HvJ1L0OVULrDQyNJbRFrvGNyxFTR2H5Dm/CQvCAsc
IjjCdkHmyB40+JZhNOgL7xEOdpaDYnPJVp2B5/Hw5IwKe87eqbOXOfWOH9pZnZ3w
DtLc2abuoY/U47Erj6vxq2x9b4regvI/2AxB0JEc9QUcpbYjNLhjdSc7Uf0oIofO
cKeE3GsqM+fW/oL6jDZnw4F8Nl+OdV33SL4FRsg1di4Fpak/CC2UfRQRlvOUB6Sz
TNPIdeoVzZ4OnIvMHYhhqxwdxjOFOlC1N1AXiLxTsKudakPMPgjbgwWzvjtQglIB
HqEc6KKlULJ84L1oF4fhEg1rukYGGNcWWOpkOYO7675tJFQW/P5EFTe+nJNrcZTw
uFbUfgy4XTqpkRARbt+8NE+UXpwDEv5b8ikjFcnyvC+7BKBMYbfVNHd0KY10HOMs
OnIDyKWE8K0Yj/V/QpcJbkCSwII5nasnf+7lKz72wlYUQRyWNBo8Mq4hJbG01mSj
C9dGdigAEIltzDTc612BWlVWzOfiHR6SATZZKC1YLmkcS5tMmJ0x+3vSJwYDfbQI
QhRrYGTPW7Rjra+aI/DeP3bL+n/DxvJFAWFD0yNcfhpPiS6YlWE6ZJ9v00FbWut4
w+ekz7Bi7ZEm/EAAzIvfpMw905V8eyA+W5D56ln9SzbCnJAznTuuQrMiKAAgLPsm
bDCwG+KJaYAvu0JHgz0/9nkn5ZoJ5sYDiEZCEbqManP82fJMvuquoTD67N1UhYOS
PQsfILu32aoRLc0oqPVKCKuLjhVkifknjgMAnHKpnuRopHTGQJei7krV1iZeZqHD
7LL25o2ztab+lX3aBq+88mdKiWBVfkpJO3JriqZStZfQJBsKk7GFfqUfvEcDL/YG
ohry6PYfHt53PA/ddSeOmGwbtz5qxXUk6pLKjjpCTzAoACr1u11PmzoADbyku0vf
3PWQjRA7uFCN7XNscVfR2cfiBurbFZrWXpl5kQNNnsIugoFsbjXcc6Odh0DcswNG
dWnj/vVIFKY3jdjzz/QaGSJ2Nq/0/fD70cXc66THdLK07cDfvtGP/D24mmDfe7kf
BIrUyrGgfKgBQ03vgWAidvktxal/Ij7/+ECLT589h31pxVWJBR2c3o8JV9lV3rp6
pG0wGRQqe3xJ5DrKoS7Ue7jFnlDJJZ0cpxxULxS3EY6KkG3+DW4rR5BnTmBZztvF
TTtYcPsIhBqiw2PhkkKL7kxvWasz+AihJDpmqPVslRcOD5nkpPUmaycz+ys+QiFl
2eLtY2HVZxDXUxvLAfq8rpFML8gXhotnEuRrjIjV/2JqPSIMPxHT0PAQwzh9w49q
u51hhTrJfzrPn0UdZwp1d2XBhKdHsintrIAJlU1Yp7Hu9RNm5nBf+53spFx/58rr
P0iMYd3eQsAX7Bh/+VZIZsb6yBA/0jZpucZ2uJI3ep1TUNKGRHQwr3lyRWd3+AtE
OcYadeli81ZABo7MzC1FUNUWoHTrAEHZULz6bKK86FgKisD+qXL0GjA12i6PtUPi
fBe66fTPPjric3LSdAq9f7czlfNovZA+66tahEz52xk5Q/jnDuDMjsC6/lsvJ2SW
w5jBqlQez+QSrUKiiXz7ffnQMpANE/EY4cN2s1629d4DnDHwJdqZEK7HgXG9T3uF
AsRYt7iNjUM8hQygYlx98xTCc8IX7HHP9tCi2PF7ioYuzpWXdWeC+VTRqwWnahsj
o5E06LA2KGXl2sfL+tfPrQecCMKL0DOJw0Dy9D1Su+LHlgfnV17k+nEaJZvN3q/O
v9xrcJhZForvOSu4zFd5UWZphxsxZFrRk3G7JJnvABxFjGbNGzQ/zXJlTFHDMcoD
xbLmpBABUsp2RC8x4zrlUm00TR8jxOFurgjpyXgoekfj5DJ1vAalX0FfCmJHT0N3
WjonkQXVVIaYGzq0v27eEiJjYHxAh70PI5sjEqRKzdyK6FfLhHPJ0wtoqq6Dvz9a
ngFkTnIIHlbw47y6CoJgsK6n5z11OjRsjY4V57XL1z2Hs7Cfb1vXNSW911gvsEW4
fu7QebFG/+ebKlJgXgjeDcdZNzCqKMXae9ytFvBOjTxmfJ1ddQlHG8DiJGJoKEMD
lwOXnx506QahDZfkmor4ZJ1YYneqpNNFFsYieiKUS9W/dhqDPE/WDXQdGf5C40tA
CzSZIMal2ghiUwptvpIq934CN/i5DaWIjLIZCDtVriwBe1Lago8wu0zEi/3hOj9c
RftVIxx6d4Nn/T4mIwfKK+lf+GqJpL8d+Fsp6Jh8ITzPtuRQkv0a1oWx365ryoIN
RRleqKclxDS0EbjgisJ8W83EIl1P+IEW98ALj4b/BB2ySfHsijR9egjiqpQniER1
WY4PbbMxQw+dy5RR4ZPwOAa+VXXBAY+aO5scCO9doFxlGA7Ch/mBsWzkBfjycG5t
WauhF0jZ8Tt+HpWd8sjFfJgdzmRcfVQKVS0Bu/mLg3WaJdMsm7e2E/6b9ADKStDq
fbkr3pHWXbfq5M4n/U+iAwsMN3jraDbfrgEipm9OuhkdWYS9eILlxQKPRJQ5FSZP
Q9DQpbwUNW9QPTb/Q4hLWIEcZtRGu57g2yX0Cx+tIYWnMGhOaQs5W0YfBbIBlhgP
i7magqRRS75JuKyZp+Dj/mt3taJAyz7xs1zrUw9UQX2aEP/pm3WBN4aMWNEzr3hw
JJgiS1Y+ZJ3HQEZyD8FMRYisxJKqIsUtOaExmlECguBpFcmfa1QimCEYX6QT/rhh
jQlm/X6zAoHYh4WIAR60zvX5nEfPCgyqAvcgEQbFGmmaS7VWUbcJhsjFF+ua6q0l
VAbKhv86ahS5EeRVAgOok/3iSC9waljAgx8TrcnhNOYJ9Oq2pKjCmVuNrR/yBeY/
/Y/jESuKPzU+0DyZXXMUmepa1H9UtjEy/rM4e+qhk2qWerMaG+PiCRMUWHGDth4u
VVL+sEe9TXgsA+EMuRvWjuKyIoCOJk/R/4zAArrBl8+h238l/jxYrXSkI4u7YWPr
LY9VWUh3mqNkP/GvYVdMjYaUZPb6OoTMpePgKLslzdy+fHHcJoKiiuoUm0MD2op5
D5AM4M2U0BbKuQlyDz/IwXMexGFas33gfd0RfIkVoNBRxsiVueWHGvznSktqcp5W
5zEvMlX80ihWnBwyYZ8r0PdVq0i49SBxYeqxnfjwWnSBlR1sDzR4GlCq6f6K6D6L
0u2W1gHuMaLkg97npefp0CcRY8glGKsBKNK+N6fYhgxfYbIGoEPgyUJOyc0p8qM2
Yx1fDXdZsPaIH/8dnwlb32bkSIjTNh0DKPnMtyS6Mq+POqxXhGrJheE75kKbPSHx
BQtAOUNZ91B/KFC5SoUXMkVsg2hibqRmCdC9VhEE/bfNg6+Vcw+f9dNcR1YNkBFw
fLJOOD+S0UFmmJdOCt9I3qDjJ3r+YRNv4K+9qOLJp9Lukvg2Aa+npp3frKwnOQZM
5+G2WF+JjXrjUieumU6bFaSmerjuYJcFIVT6Ttsm0phL+2oHn3M6ja4r/KlA9/ri
z7oQshZMq8Ys+I2w3UIo5qBlyQAK4LLSWyrQqvj7iA6O5jE2LuRHe5DmhEHSAB9X
4gH9EKjdup1hSpiMUjAvlE4Q0d1XZp7ywoHemjeHF5HzUUcCQJrPtknjK2hzP0zs
tJSUaAQkv0//wHv91bspoEJbgcoGon1lHPAI63+MjEjFwwh/l7B+iSQJYinmOcKA
WrCq3qE05ZrOHmPWzyDB8LX7w0S8lJ6pekJ0dgMFehhXSxfYcyEg9+fNQrDtZ6Kf
r9bVMAIoZYbHU6KSf0ol6K7udXsPJUu5myJa2zgQbXIiuAG0Ge5N3N4qJ/aPMTxI
JuL5OpbDK5jhoJDkkQjL0zs+LWp4cqX0Cjbo4HvxksXEh0e0nu3JDYJLifpRv0lN
AZO9QaNt+z/I5Wftnn5vvVNw0mGKYwmZy7wM9sgRPltK1MytuNSVFATPkSQuPgry
bf6Rm0o04jQhA9FRLWyVaMxKWTe3fpRGZR8ppHa+I8AiKWE8gUNPy6x3m52Cd3ab
PUaumR7lTRFtpr8L0clb+pzhnfEMST2oLSH3cRbpta5vtcXVC3NOruQKGizOtHwu
UrZVcKV//E+4aarLMYqPrUE0rCnKbBXoW7cDqWFPZskXUoGCDCAvlYHUgh+QOTe6
2uo5DYEKcMfDopZrSG+qBwJp79fbILJ8MpUykFpDc+S0UMCzPGxMuOTuuQ9oY/eZ
8ZH6Dcjk4y/YK0hkHomFY3diOwEUr2cZywp10jkN6AiJ6Br1wMIiQlVaqR9aW1zF
AGRMMOvuBGRvYSffjCKAFFnY2YZHg4+kaniRyoxXg77HR3wdKwMli5s0MffRKEj7
Ucj1mxUPZfxQA0dI5m2sdPp5KrP5Q3ITwILOpDG/I66nYZ6CZKADJC5u/kF6LoSj
jpLN4dbbqJ5ci28YTjgNXYffS8TgQdR/Q7Y7FihhxkAb94OQHe1dBtCNCYm0hL27
q7t/5zovJwKMLGj3XoOOiGoUdujAjV8/LZJ3Z2lqXjfO3yoXppoXvUFq7t5Js22y
V9oeLloNECG6L7TzF/qp3NYLTTprzIsEeqvgNAUwwEPz+hhFxfTmbJIvqfMUjpG1
mq+j8cwwIoEkngOgc0ia0g02n2jN+vVAvU+Yk40KbTxcmQ1D0ZqlSLUnDf0lXt63
JEIcHC9bmhmRqIRbCZv5O78LZhE4jMookQXD9235HkR03SN7o6mqSW38i2ZZbN31
bx47CEPDj+agth8TujbEg3E8u1Fozcr5UsHXRmjIWTHVAXg+7zQaxSAzYleCGyOy
/4zUdwfO3QPYkZMQ4u/m7WOVVU7tumO3aiI24P7zJHdPXadMvv36zoFjq1006N3S
2mUrTZl9+BAhPBi24bmcBig8C9EgHx5DMS/Afld03UMf0KiN4O7ofCPzsBQbuDWa
7qJX3AL8NKd9Z06DcoF7PrnPES2cQLhY84ObTicbLZ7Drd5hJn7dg6PbRIr9QdKX
p/WPzmwAj/iDz1f9CGK2y0z0x5QFFK4g4rxqRCk3FW+1KRsT8BSixR4KAMiabZJX
LpWjLoN/w7TPnO2BdpNKr2uiN5NqtYTJ271zt4brSo7OU9mrHY4e0LfiHOg1Yv/v
mjpZ9S63uAGXpsf3dBfXfiCTwmoJ2enQNlRVGzwLa7XBLoem+XSwCE4P7+1Lkop9
NwO1TMXd26bWJCfG/VvXXYRFgQar5j6r3B+ojv3/rmKogVoiMwSj5K9dm8CgiuoG
AhfURsA+1kHSGbJVzDB8jNDyVA3IR67tI3gnVgXInmLzFUhKskHNsLnhJJqWmZpX
hX1AZwVo/W9anMHt5OPO4hzZklsPgGDAt4T2gbBslAsPTedVO+CN4BA1fBQDvxp4
37e8ehvZpzw4cCtw3zzLXoub4Ghmh4T57SLyFgaAu/0VHmBxkWkKD9yVkj7i4SHB
pd5iL6IyD22jf5druabv0R6d5q+zO9cjZzF7ONCYGao6hKKiaZJ4JKFfrwgighUa
KIOJkk/7+HYfF4YXqWHsHzniiG90nd2G6h8I932N5pt3bUTdn6nCd5VuDJirKzvb
CgPyn+z/EWhQNk81sfSFbaCykw32XGtFfZGiXXnNV7MDbhWyzJ2cvdufxEBQxP8l
wMwK9BQjFzh9L33+UdKCQFkS4Zb6nizdCBLq6RU9TGaCWE19G30Y6CBQbCBBTc0L
BgzJCMHbX+K61l38wCSMmvGeR0iMlTsaaRjgdgIzbyRhgS7DFHXmAZmL2aznZ+fL
aPsPneTFDjwZp1zLkhDA49kmCDT3pfnjDjDCjXIQL5+r1azznSuakex3YPcN/OmD
Pa2u9VYEWXcH3H+L8rZXqtiuCZdlbOBPWZ3I37AwY1ZaHW3UiunVcLZVAx0ICftu
soNj5LkUhnVqUHDJFV6m9c3SHvGfH7JoWYxsEN8MNpW5KiqlF7okdmgkeN4sohsR
tkT2hnY5xzbYlfgaI/df3H5zwqDlQxUpHwz/tY+Bo2Gh10U6LYB5wHd/pmSrSdRK
sRdk3+7i6Qrl/tIBquJAkiVvM4Z7UwTu9nPztQPoVbXKrU2rnkctBBQrkP8SXEVx
ruFvhKcFPOHnyiz8PI9cKL6e6xCiQrlTCY2IK0Q0+VOtu725p+9jd0PAYysFVkBD
dUnwwLTcIOETK9kekXVcNLL912NhYQk1vlxIeT60XqSdHkMccuStAkqjqvHbWEsP
cD69ZUNl4A2/LtLfLxaXuSt55pNWzPV0PgT6yKSWoN/h9z5T7LaWFZ23ahlv3KxC
zghulTjlpomW9rTC8EnpWVC9GHVJL0AbmoiFE6IPzK0xW1ujyfD51KNg5r/5kcAV
G5x7zbzyYxN6eJC9jkZQQy8jVz+cWYVMsvp+pMy9ejKX5jKOkzZUKLR7OMAqGWFZ
ggXygOCCmlU9aTs3CiBvEOAbUQVfoY30OipXnm0Q7nktPIQ5BorppwDk3KbGKI3l
f5dLphaNCx0Dx3TZBMI9ZUVCKEczl3glo05Wz7QHGHdimskawTZCZKqJDoyDm4E0
HubD1Fysy+dQsZF5hYOjpm+KfC6r3JvOceG96sZ3okSoj9NsLWGtCG3aIE9b0jRh
Q51GDrNZ2KNQR4nOkiXISKlnCmU+0AdYNtePTHkG4MkzRXJQr8vstzlAv+amYHbT
gqC4GDKJKpXGlibvblum8rWya6UHb4sC3HvcarBXOrgaxmcKtxEB8h71ii5kxLg3
upgBRdhYW4VjcVd4vvmj+enFcEGC9HWqza1aw/VZVBRk726JMzIs5VgEaTlpFV72
R+aD2MIS2HsjSIRNClsIf4ok5pEAh+1BhjQyh+FMRVk4ORRJ1/73Phd8nv+q7ELp
sv/x2+KykJIOdyNX6CiQu+0jxnB70h8+WOgT88qKdSk7mnmcJV8ssVkbL95jnzXV
ESBRJaINDCbsMB+Kiob0PZWS5f8l5bFRTX2R8w4sxwHRDKIoleGUKkp4Amc6CuMb
A9c4250k+yM8Hwzr9NZAWW6H06mHazMyOo9qa3k76K/RpzrsJV0agZV80yQPYi+J
tGBdDWFiBJEMs1ruPzwhWOHvx/NQ6iTOHqsqx9pxNjPgrr++vI3rAvQVVfGGuqAe
dwp5Zs+/YI1lIThjXCWGAAl82M2WoVuSTuLj2p42nPTUqU9N+eCz90ryHTgjALaI
1yeCs5l5I5o049KfMWsgKil/Ift17wWGkeEMLRYCXhH5h6Y7nrH03hqyQC7Tz75B
/vmhbeW7qVn277IANPU+2GY1BfShTfcJRbZPRA1Or2rS5cp73eI/nMgLoAH/0ArP
4cDHbomXuTDgP+i/fnNDlenkb3/d2XnYsHAIzaPP5xC+NTRHKRR6h167sKtoneaH
NnGzSbnVK5C08luxRbRZ8ko77OunRiWGqTpRWArlAtaIkpqzTvH/Tn2E0bCyXOHA
BnGTLqeq/pVhFcONr0dUalomlKT3FFAtvt02KIH5gZZU6KcRENUBFj8ZxSIn7YW6
jVFfsPAala4eIxmwVU2NJW/AlJxY5ql8QkE76DjD6sEEcqU03Gyj5kJX0mhY6Ado
5nO5ojuJMtsEI8SlShYc2GHQSlc6aLZk53oUjSnMppJ9PxMQ0zDUds6Cxt7XPqV1
iRPLsaLKPoW4x/DZCbOwoTQUcUfBX1ov2GpkpSmkscUihWYNz1y1Tn2PgKhAHxgg
CZSFnKBdRZeSk6YhqPeHfmun1mo5piKESfmrzg5NoXEdLgQDOVs1CLXqLqJosJdL
zDxoFQZhd5cN7fZreKLdSbzK7XetUG6yC3Y3JarTIiTcP8rPbwDIHGeP9WfibGrl
xOl1ChiL42ny81wIAiprGXWzChpokC/p8HeJKtfMYeArx/99SI0wBiZr8jo00VeT
36Kp1aIKlZ01zPs+cV8fQ08JyFzXkZRXTRa7knrFC2iTR90rRK8KEkF9zxr5p48h
N5GVJfehrZ4pgWddB4CPYDAjm6hPvux41weU/VfFM57vQBBRM3bJ5+XA/96xSbI0
lZ6gUCl899noI7fSPE80fvtdbwFvch4LwGf/qYNnmfghGFMBvOWla7kcleMMgILU
HjhTWpd8geecVcnaoVJV3imTm76uDrbpgvcyICskuuFp3OzcusuI0+3eNT2LdJtl
8CwtMSJ9zK3Wz+ucbKybjUfeaIDEJoszg1DJ3H3pufDKpbR1RvY0ri1BIAjqDAJ5
QB8jeklqrr0b+7mD3ZkJWgfzRy8ckYrmI0G9ZP+HsdrrC7Mh6DfB0AoH5OT47T7q
CpII1kFLGUta6ZKLkad9bAiF/TAdRl3kKpbPYwzaemf4UycIdFzHuRYw0DmMdf99
OHYZpuS+rjj7MjOUEBFwtmfXy/o19mDk40I4hAuyYiZZnm54zst552oIi1tVPyp+
ZmUX4Iti7DVIKK2CLj/hYxOaWwWKbdEAc9dy2+IK+O7ayF08PILUpVaHzybibyPz
g1/YVHp2Hef07gvonuZvmV5Bba69BOQP48Ij25LIIwcJfsvIWWoFkQLy+wnVn2LF
KwuMdaMXYEPVI0OF48Y5z5RIX2glFXkepmkXC+gABdC2Lpt2kRQHNgq5RgdTrpVf
z/Uk7lQ51i39n7UoYsHaXUhUG3mZs+MGarpCI17bZzeIGzoNjQCLm1WW1eXDLNiP
eqIyR4iA8smlKS+O/yZOmU0Xlg6zVFr3wrUvabo7ZKeGcu0YaTzNukXPTxHcvsXy
ex8XkI5ZqQkRkKqdR7ze9z0nhtb9y/s1AvsRA8Tz4jguIj2PqOiuHy5KtbRFHPOP
QGNhKZalpKavmXKcpnufIb+xMt+OfISDjQEeCOpBktnIBCsSlvFxfLaeLXAcHOhB
Iqvynnn8uvirMEhJZlEHinAtH8g7KkM+57HGAGZkXrQE6qSXW9t6EnsLudexRR9l
jcxitCXGI9SjKC81c20PpGc23QKHvgAeUWoV0e4+94Fi+ixRFPhghJNk5k9UPF+n
32dxTuijuzNlMiakR217Xn2SJaCHI5vYq4MRQOgRojWnG84m0mPi+7OePDnyWflX
THqjWfFgyFbyl487GNQ4U7f2h45so4Z1LKqvFGEr0wakYZA0KydJGO6aneNN3Hj9
6u1PaDZBSwZaypxNFQLWVgyPLNkpSY6kXGj635j5/F0tnNyjCRz33aWPnBOrcAiA
Y6P/TnLco9d84xs+jTNTHcqOPzr64+hxg1r531uol0UD3+IdNyFJVc0j8G9K/gdi
fPAt2I0avlcS3deEYtYmMEHXaH/LfLV9mWkflGMaYJx71N0+mtStMj9pjFRJdeyS
+1fIvPkONpGjUFKawguf1kKqKJvzPfMwcOP3JOK8OISm1ahTovxeL0qzA4TbdxmB
ICX8LdvwuwlYMP+b0P+o8WdqDWW30iYk7cxrg3ttXPjooWfL7iaeTwgL+Eql+Yz/
L/1tiQWWJxDk3LD2pg8Cdz8qXuyaJb6TzlRb+hNodw9VXjzcPAVukJOip/yrae7t
HkSRcgnn302MMHN6qHLI6qRJjesP86rDGcUCaWzMK+SpX4+7XPacMP75oXGTmOQr
C+sg3Ty7WvfOP163/s3+yOrxXpTrx20wMlgqAPlkTuE1JBHms88udbLRCfTW2apH
M8QrI8R7xwr99IG9C+zJwP63KA9eQ5IB0MkVlks3YafvnVR7mVU7iBkDx7Igz+VY
9ubTup89xvRX7Il5KxYaGxsuyh48SENqc20JuShcPFrl40ugLQZtrXFQ77rVArUP
3k/r9+fUDjElpQEtRBbGCu4cyr/e9SYGIX/Hy/MoRjOzmVYtDEQKMKbIe/BeAjZK
IpH97/65KFTVLgE9CBSvnTfVBHXiaxHNwY1rmWCKoDt134pfTk9nC2oNrPdZz8MB
VMew6LwWTPMu0qc2EypVpnY9l8i5zhEZ3t8i8jTlMnNMayqX0DrVXWklBqXCmaXs
Q3soWDX/i4tNmvLNftIkwQ1Au9yCT0SHZdARFucdjiclIsWpnkMLiFaecAGoCUIM
b/M/T7RJg6XNcoAXY3bW0T0EnHxtDVw8UsEoDted8y+Z811NHRru+6TT59VDD0Ml
dPbXTOh97Lnty9jQLXG10yNcQ/od5S7W4dJf6SoFOrJxOLcV5yd3SbGs1xqfhOJA
+i+DD7GSZlwNM5VzJeJVSPE6l1/IavHgGbRFKVLVwouGltZvqAFy38JngS2cYjh+
MlhanuMPLgWZR729bEquv7UrHj3UAJ5eiOGHJ5qsSjONLxXEanr5vdcKPmLl1ZvT
iXlcr4CfibqKEoNQmUcY4dM3yWeWke0mqS8vS8ItzECVhQLMOyDX2h0njydfCSJb
zXeqOqli7ZhX22QRVrDvU/7qjSgTstfag5ashACHGAE4iaKDrxxs5PhX/OaR04O+
6Cdl9CncvAwyh1be4++ER9/vl6QsQNGzXc7OO6t81MymAWGLtrtmiFCJZhKl6EDs
kTER2BlU+JOEZV08CmqdAJW9kdyzjonQ60aDxWxczPoMNm1uMsO5Jh8cnD6FwnFH
12Tc9wF3qgEDhbp+TCrOMGZVc6YNZ/9mMdv46sDJBpO2t+FQnCx9S2+A8KwLTEKn
JWNuHoUIGjGv5cArh7gZ9LQqQ9H1fJ/qvrg++JNdBBG34TEA6p+W8rAxgNK6wnko
1NpXwj9UVRXoFVvUvkqwBNrrlVcRfxHPSBZUVC5ZXFwTTnm2z+hqA/HddvdbZfj/
EtifsrtQ3k2/wxBjz7gUohIe2Hxe5irElhdwIO6ZZpmsZBiY3U/b0xzcsIT6F1Cz
kI7Pr2JBxAEl82Whq88UVrPDp2EmpdC3LV3VsUw1MxWRIf4wfQa9BYA6JwDdxDUP
d/FnqGG/sl3+pCAieEn/e2+/rj+tMNLipF/BI+cNBUgqfk8d4Ke6iGgo0ucVEGK6
PjXkBqdiQinMWSMU4FKpZEG85sAJb9YiCqhIypFRiMyKntYTurGptj+E/jtDAjiT
lzZe3qX/mE8e2CMJbsj1sR4he/tkAsz7tH3xLLLOQX28yUXvDSR6OXdI3RE8Qfwh
sYPl1sqsclDw7XZQldaPjTRFnB6RX8nTUyMjBD0BE77XPDAn24iPIpORec1t7FVk
4RPNf0BIfHk9LTfrQvdHRKuIohtbMiq76n7LP+NIe/FVy4oLQhVJtyffoIHDlmlU
C72T725kq5+lIKGJRiPMz/scDrVIhv8/vV3NlCEqWuwHCcFs+eTNlqijpHIRlB4z
LUvS/ijGd9BuHni+4sVLUO37seD8Tfe9nknu/5xzKkEx9gQVX7c/BIh++7uj7Fh/
2wwVz+pU0ufr51IOPxylrYfj9Ph9qprOqH5hFR3gBsXMFNGJ/qtlKwbKGPdfNteu
fafgSHrbggrB8ubEaEja6ftUkN5KVqU6TMPU0N2haGQMLT++pY2PBhn67PuYDRaM
iTATut5sZgHHE8blWImqOkE9uTEGLRVK2Xp4pJNtByevAV6w0fpKveXVA/+58p6t
6oUmJO3ozSyFD10NwpAeFNtMhb1uBS83OmQKMmoRX7xaAluAt+WnnZzkJRblrx7z
wpWyOKNyAkMxvxFxxnmvSA9fEjOZtVQNK8s/60BQMq076npeoRMz1fc5IO25iBQG
eZJi4MHNw7mWNa97afYajjE0NTZ7hbd1GG+O8OnIrYyDLN5/hbhnOajPHS9mSsev
jg7pHbeacQkrOURl0a1ZuEWYdd3l4R+Nj3K0IAuvcq11hM+qyW0ruyR8v9LK0oCm
qEpUdxzip1pdvz7FcBD/+r5i6044jrBFgCMULer9P6CZlVIUGR7HYdFEAWYJBGeY
/BCU9n1szRqM8GhvN1xi2psEDvGCOdu8phP6mZos9C05j35IeWQInx5bNxJzzg1l
Nv0gDQejnCMd7YcUhY6thXShwpRcpMMufWahDJt+iDxs70jDSgEeqnfSbmXygrgU
pDx3tOirVwwDXNUxMZWD8F77caCvS2SygUWbsv1/7TZ/4WpDFCouMViX0ohcl1NS
q/qIEONX/VDfMFZ0ebEp5UMbDDRxj4Z2TVfwv/M2bUBazSDpVSc+9bmyYtCK3MJy
fDUZqDpAeWJbZKhTIFSShQp0DCm6N9lEE8Ow6ppiXt0HcMdQUMJ0/brs/47LL1lz
Oe3AM23J1KOAIo4lPnPSMzzp48fHFdB9irP0do3r0QsSGfuJmdY21i2aaBWOq5m1
BEKsHWZ7429BqfcDPq2LGNkyC+sck9C2EdeQyy+5foCnH6ixxgwLAEi1J0armuG+
aGDBjkP+5tr3Ly1r7+a2V40dEII5x5y0hRV/ohnYsmRN2DIqf33vDdWp951OlUJa
f36hB/mN2dUuMqbVgHXZrqGqikc9quEP11knm5RjXCalVzF5tRcBWVNIEmQqB7L1
ewo9iCQ2+MhA5oa/gFGHCKi+aT1XdzIFT1hUPlWVYg1FF52MXZ4AGpWkp9xcA8/P
gjB9a34McnQkwporvxbYC8nStSP76R4uBZYF6XSwZKTmOdcMP9yLL2nH3M/NCraH
iAvw2sDef9fCmLYuJPCugAugS7NitUqIAgt0gOj0Socw89VReBF4HkNiRbFuLBem
48KWGUJgEWJ1oFm1WJ8AOpJMC1YVKLe15yM80CEz6KRscfHqgqSK8yL6AHZYlyH4
cjsZ5aE0E2H7WywfRCuDopmr6e+s1Yf35KLYZCTHnzl+S6wp+B5WJjg1pgGtgEZt
KVMMwi8n+cNJSnp6oQkhDTmp1M7caxT8eri8uUXgxwd3PLahgMKNiR9BLx0hylWx
6ApwPQDkzn4/rVa78/RBiMt9q4WkE463ha0k1dYoJdOVLsOABalkq5etL5LkKggw
KgxchF3V51QFhrsS/C2XlNiBRN0yeJJ24a84cLYjUFFbluDul08JYSZ9N007Q4P1
rRwqNrWsEZEUEmvT9fqJHOXzHiBREaA4M4ZHvFNeOyTFMQer5zzBGPE6LxVh0gYf
nULHawjwkqhVVjT1Ji8KXsT71yiLwFnJHatX4t+LxefBhInS3r+ENEwHxCyCURgP
7UZXIIoqSFEi8pRqE3efhZPSIywCD9ihcQgmvlr/l4tOFHwykxhoNk00lSSDtJo3
I9s9IdbpWdGdPt+VEvl6OH2nMePWDYHPOMiU+ZcbQ5PCNL1usRzSkVS6tqHx3nvb
UCIrrPlmlYwGe4RO/aa53EnEjZpDu4DLSNhesc297f+AC0zUFns0lttlbO6U/HRx
NsaHHyl3WBy79TPBc627769N6SYpTB6zNTzGAr46h9yQv0fxhPoBqFCqMbgP9oz9
g231W8WeOjJMkReXHqVYriiRKzmwEnUXM5JQbXuRCbV8E00UddMRbXaneK2DQ720
olkVtlN2rXtFCoMksii9tKbv581ZC1JCC5fH2h99KzAPUeMpqS0ql+y2gKoo6air
sgiG2Pts12EEGMG986aydFExFrkg7nkQxXxvxxZ7ApP1FtZAY86XlRmoEMRtx2h+
MEsGeQdC4Ml7nnqYGULCIYlmbbIvbiSf7YH97G1PAyt3rvWIjbInM6zgLqFrcmeE
5NZeaDCJfxOxuUnRjAXoSE5K9w7Lt0rYdVtqi4bDPZI/ldMs7tviINfMypCPAsl0
5Qg9lP5cGd03hKMkTu14Iv2yE9td3mW85Grnmy9by/jYLfLFQ6XsOm+Vx8Hnamii
+asCB7MBBeglavChTAZtRR33/IN+oQmvEk2exfWoQyh9slJUqhUrWImEuOjx7+Pg
szJakSrbgketCR6m82IgvfWuqmKS/JZ7WgbWqVL8d0N+dbJ5hmDh1HOKMHJjjdoM
miTnrBqNXAApdYtJFtHlLO+zpjQNJ+hTiePoRVZMT7pNfBFDF+DpMwaWFfdIK7nw
YsUNjL6AHySDHklw9gJp5BBS/lLCsd3uxmYyJ3WcmxCGT4r2mkYKEPs8eHBZjHGy
whfJqfV+JR5NT1wfbf86C2tS53scK3WeS3RG3zpPLMnelAxSGIBQJjnabFXpR4IC
7QZaxfuy6pKhbjDaGGDVfEURyDYavXsGpSuP73L7hIuY/HSNWvkUWm2qeeX6tIfB
fuPZ79Lxgxja+InApSpv8wVOWYStGY/PdSKyc7pBhasXsLi26BEAylekJ5rJRAdG
JXnYRZxR8PVTbozy5PLhxeB4EvzrM1sA5+a82vuOobNnlVA3yMtydlPDP6Dblrkl
fVH4WkvchvjcM3j/QRyCzBj8BEbh6nwFWoPJlbJf9mP4uuQTvNpQdkNQVZNsCOX+
S09SyL3oSaaEyBrh3dcYt/X+/uZ764SV7XWTP39mTSZX72f0VklU1N5OtdUcOl+t
4wcqVpg7upqjODBlEYGRV+aLFBPGlVsWdD2UmuDOTRPy2r88WmKkQRT0yrm4cMIa
U0uV67H0InOB5k10L0D6oDJqCwlk9G0JinOTapFYXZhP+c+X3rIhP9PWUwvsAo50
XNVCQ/GfsGfVUo8WULYKCo89QmEJ+rjCW73Bpj5tOAc+l9w8SyIeWkKljDAKTXFf
9t5ywL4jSvcuzQDULA6yfG1PrEJ12On58RSSgBgiiTfVAVvsOm4VWFWVmPe9Trik
akKCYQo6Zf/ovIsALbBU90SxDqQNFZImLZr5asSBorFHxcW/SPQT5Gb01VO3fDbV
0Pg4XSRAn2iKOPVidC1IEnSEh+ZNLlTvg9nP1te2GCQbD77wBxonQExLd7EUBYAJ
xGNES0PpIDlkyN8H7gLbREuDB43LOHVZMWjqbfqXqoFtpFXz/AIaEFhJSqsKognF
HTi4wsKBs6Byg8B4aoDuoO3MHouL86vBsLSJHKtiffdfu7zidDZQ0wK7Xg8MKR/4
m7A2ATYGg4y95Fjb5NSF3CA43+WmYE3fGTUZ+a8+GGccIs1+i1aEiKUoZRP9y8P6
fsIn8P1tQ9QHX/UNILGz2TbdggMNj4YEDDtSXHxt3q6MsKlqpmwc7ngNmQyA853f
FT57ixjRLd3Nn3Q+EwpCiM9oBs41V9Sqqqfzo8YO+s0opQswKXjCjYc67lcIIbtT
JIyZnaR/RLE/DfEGJFzt5IMhPpalFuaACZKm4olPBXea6yqmmuHfqBU0TtX7oLWZ
JrqzVfYdYrQukETQQFBs3u3BOBP1zwZ0LYWBXYv0WmJJrIZhnZCuTSzYgrzmvs8N
FRLKwazZvdYd+sTthE1A7OFg3Nx9+p50PlYo0i6GY/ffwtLhGnapYkQEq/utan3v
FxnIBlnk0eB2JtNdOKKVxyD+VZG1SXB7mPIr4TREVHJPu45vX8vE5y6hlW34HEbq
ddpFuAvzG3zNc+48/0Shc9rGhv5tmTzlw+zkponE5vYxwvR4pGuhOXxn7Hlnjvwn
AR2P1q3f094TygOXiZS0rUYrEd0a/4ayZGnPAHB3hgdmmOFtADuKeDpDo+nMIn2Y
hbg5SRqkTX2dkNEe0Y5g6ZXsj77CaZQAllW9ffG+2hmlESUvIBA2LB6yDDNd6Sqx
LuAyYsprEVScD/ZKjftEMkE+ElwGG1j2EeP2VzbMq4kMJqHwR/phCvk6IsdYd8m9
54DW8mqZSazvnK6ce4CWhScODQjxqwkzgpNU3lTXASwjiRt5Wm8/p0VNU4CslJSh
hnrCCES7zk1hJEJ6UvCOM/vQ4mxepYkg38XNyeb/vMnsjpBQV72Kd7yTBrMSVEWH
zvdBwJZCPAvigjc+1eairERb5ZY+8uQ77bPVK4H8NRk3qqTDzqtV4bS6Ho4hUxI6
9RURcLKD4jP09CDitcruGVgbJL4lvlNZDkRE5hEJ9WcP59jDyCh1LpHF6nL99v3y
oFQPMM5G/tqRsxdMzdGIlgamvStKzPN9Kel1PmS8v/yUp48dH8sZYOnZBbbzlhkW
yJMw9IE31gEzB/j3XHOOc5JgRjNgTGpFeLN3oygXW6PH/SQHwpAYAqpNed9qo2Hg
XqHPk9MhDMH+xQrRGEk5Xn/CdiYu9AWGPkG20cLYysLtWTgNYQ3Bk/4rFRcBZXrW
+oTbHGtZ2iTOZcBC2oOL+HoDLVXMbq9GCT19CiVyP7gCLw00QyHaIybiJ1OB4Vfp
KRIKehD4gMFoVvKfnQC3eK59Y3HInez5WES8qfNuWTwgUohr7bgXEnzDMt6fPyCU
zq588uhwIp8CSVk3eKFhIKa7IRTc5LwxbGFNSpKTYniKtVZNNh2ixNk9p4/Dn3S0
/jHxsV5Cku2a7QBZv8qo86F9KdxCAVUKNtx9gpzfCDrJS8TUPiFlzsxW1I2oK8Sm
+QOC7eYcN2Y1CDUm7MVA2WebtcItIZDeInycdIYWKwiJwg5b66X3caDCfqKuc/J5
OZXkyAKnNfXB/P8fei9nAmv03lzE92V8oOoH/Rwg4CuSZekt4dgF0klc4+9/VGA/
KgpuHdC7caYLQoW8r6smP6fyzobGycmm3xKBHVzmLYEBDyQt4T2XuVzfR42Dih0m
yqElImkYjrTYD57ilJSL3Wjr3WeICrbvNbyUnHaJ8fM/3fDKhmTaa0i7+y9xff1f
6ZWxYPOmm5qFXn7RHfbqwgF55ZLvRm1zHbzT23yynl8EpheUWyxadT3jSjRCjtfk
BY5XOMyyMSw1QaZ9hj1XS4eOuKDYDINixXtAt+NEQQFgKIqtI9jwGBNlLjgA4VNy
FyydPS+2ImqDJ9nxov+TYXnOQ3idvfuTKf+DHDpKk8LJk09abnCqCETUMjLQYe/K
P0SwzMgUS6MnZOqLiYmQXSR60TdicBaWBiYX3z0QLfPc5Lcsd15f+rlz2yLx9MC/
Gk18Jsfvl/uoZyaLQNnky8Q0MdoeAuVFzRuOhkACj6n8qGhqYC2/VMe2GaqO0Sve
O36cyY3H4cbP0EYlYdwZbzNjkAxZvEaKW12JagUGtFvGWnozm/Vv0el9oOX5qfHu
QoR4wEO56+PLJe+RSRrf8nZXizsZ00qhW4gLVit/7LKkskhnXVY9ntPTrN8hoLiB
ncsLRcpA3462oMIXOem6UxoXqaVvsYGuYa5GM+olZt2RUgi4b0mo1PmJGl5tWGG3
t1+EfZAUmLjRpdHHy3Gv7eWnp1xiIN4uuw7PkZ9yEZ+jbXHZOIguxlFqfK42MjNa
YoEgIjBXnGlz0HuJOEWtfLFkIRM7gkUDrxwGM6Z6reWcnNq5FISdpCiSILYqucNk
IwELsC5RQ5dNV+KrbP1D92hN19khPWS9zP7bssX0Nx2dLOATa6buiBBljhVJ9efL
uLsngqesoQv0pEEtzPm/grRN0M/Seij2IsIy+Lomg5D9doKl0CdvD+eRJFvDNlJs
Ny33BPZSWkcwmitTE81QTlue6azAXLJX41cmuraopi5djz3+dfqF8A29c0GMtpXH
XPcyhWL3UQK4ZqqQ4qk7oLq61T/WpmCzT4DQugAUFJnJqzXloORjRXbPrD7fCbUg
kJcHAKj5d2V9JLq3EQuqxlUiVIKE6BxrOMAuRHa8w0bnkeYUPSzAxn7tvabL1BIb
FZSLu0zOhJRorBJr0jzGswGaXgVr7+4VWfhj0SL7Hpm04R3BnLnG+lhrh/HhRbh0
/V9qtskoSrFseFV90+dRXqu/Na50WaOMv88LgNETeBWW1uGP29mgWmCGpXPayOS/
mK5sHyFd7aFPHAIYg4A2ci7MC+OPxBboj7oYDfrt4A33NMAUCbs/MES52BEQJsXK
2ySci9dxTyV0QVQP26yDIgRAVuT3h6G4eoNYHgIg3EzYzL/MYzDtcEb0uZKhs+kf
aPT/yTkyIkclJq5Yjj9rwFGh+bzGV/QCMQaZtVTGg+V52inBsQa/lBMdgTyUcaFA
5lMApHECGzezUP68POa3e+myJZjo5t4sBVTuv5QXOJnICDy/I54bSfDqvQIfalkl
4zCFkFEthynxdBYECQCPuL8SOB7WGCWzyYZH+yhMyqdTnNOVSFESEC40cjgqnrzv
BDeDD6TpuQDdtnvFgf/7YSt1vOsfJpwGO4cufHBFV844KGYF9ZSfWyCIuMTVHgRY
zUvqAg4YLsYJfKM5yGGLmsDgxSuUzGqEy6Vkxr6s8GU4D3sIHb9AT99G0aRaes9Q
7q4rfFJ8uCsWAsH3XlncI70EsCjtExnLt5/uKzMsGdce/88/ToXatKC+/y6AHeeK
9XwFISfDf28lp4lWLlGD5rHl6TEE+v9vUBtl0WeWikIHxkqyIV6GEpGXNQ90yOeV
bu3eU+D2UidxLY4cw882+7OUeDFP/82OzFB+eBi9GCerBodVvkfxjD15H2DXWILn
lDtmeV5jJHPyDAIrArbNBsukndBuWNPg2fuhmngQCKYq6oLECTZM/L2+K+/esrpj
03ISMU0Ad28H6Cta4LwsgvXBN3PgKtbN0Cb5sZAc56rcwO9PoAwacPHBTtEvOIvC
qMPH47v2MFuVUhAZTljr5NYaBy6Q/s1l/EhCR7nBa/bC33sJU2Cl3y92icqwlGLM
urXUVA7CXrnELkA9eIHbDgIkK/4LdHfGK0MuycY+TyEjjZJ72dGXVXncR0LTprAE
3mB+ri/hDCmZIWpQrbw+5Du7hjWZaJATT4ZygI1xRABiZ5IMJpgBYa6m1oROqom8
5AinMM1ghNFQrsgXbjrtdOYWzTtefeESq05Xuka9BpNrVKiiaSGMNPUCe1ZbRJdH
eSq6BFPeJgYLjbQMXmCbO6tzXRbbIh0E1N0Vsz6gCUoiV38ANGhqURx+AzmCOfV2
Fi//jAXm8PN5D/agw2c2UfOB4mzv7lpoAEYcR+zpBLfNt5juX7zQPjM3RxOIgpay
8Rn3Zt1BGfbUxL9uCH9bc556Wv4gQNxcPkCi1N3CJPIlCxNG9V50zLSRiE2LDQyr
adxQA3xnfxyqfV22uf5zmenb77wAV91GZX6pnDCnKigKVD0wic7i46h013QigtXj
TaID65qZjp1KmVSUOVhDRk5r4YL9V48ycwHRp9Mb6e3/phyKGzL79jw+gPJX8WXr
7oxQr0l+3zSU8mJdJzyggY7885MPnHNgmIxwVrUV1PJMeLG/nJSGNFQVrTv1RLUU
2wse3gEF4/+Z0JMu3ZZu0o9iKW/NfD/I58rhFmZzr/CaXM7wlG6JiQNKunlw1VFp
IyV2QhvBuxTWdTgYkOrUbc9yaXXk3Dk8gec8eyCRTIB9gG+aR8kCpzTC7r6AQSy4
zncVYLvewAIaEXaRC6r+dr461vzvXx4ijCt0apKIeAiVUg+EoIvEtrfaetMaqkhX
9RhxBiZKMdtL1IH9zVQqtEt7POAT2S6wXhCFoiNi32jPqweVzSRl+2gPdwtp34oB
y+ViTRkEGA8TsqzEqxuRO47kHcXRhvKzFi6q6Qg1e0wR0NRIn7lX+Gdb3JyG6zrp
3Q0JAg+HY+pxX3+tgU2TPeDPLVVIv/uPahRN1YUoNlCH1uOqlazlAdUS0EuuwEk3
e+i3tqR8M5NI0ajtMWzBA6srzacnIxr0s8/pACrf1aLLgSaKIjcIiKVjxDs0v3ce
L1kVQDU2PRxs3PCNKlQ0UgolSLU4itjpN0CwNnVMNX4sEzldbEtbA/6kJVn3bkOs
aH0XlJlqPFxJp9gZ2j9IAg6P7VLqdRz3R8OYa3Zog6mmEICvqgYB2SFLCRh0d2L0
tAT/hlwaWTzNvwWTsLov6J3M7hibRNohc8sAIXwTLCDxG77qUC+MfsXQwJXF5S6O
aPLpw2DolLwdpQLYxQCZaPIx61gDhOOG88SeYhMNmN52ForyAGhaVRrRF2Swsa2L
w/OFOGlt7mIZM6Nbu2t/ff2PrQCTHoOqZh+86MwjROqTu2jiVomEIi0qCnTDKD+A
eRNr0XtxVs56CYXUbU6uZjXO2AP7zCysFb8a19Dqcl9wDxXITvojOioCfKKM0p3N
1yRwgtHlugLnCUysypHSPDY/YwAuaJtjYOFv2plu7WrUaIbGoNllrk8meBxzRjHb
i3Yfiosxah0VYEKoimHAXNgLtzPqxfJa7/ciN9YhWxcZko4dWncc8DXi/vsGcP+a
O/L+JGScnLlGrCJQ3CxeV3TOZ+LGt6iw4HJSfvE+A9huLdtQZLTpnxAYh78GF5a+
lCJPlrr12PcOP5KaLcMvK5GSryD87L0iPMZnl/x+su2gq7CSEhkNjE/M3QMDvZFR
rPPGHaSNIYYT60Wpqfpvej6niv7lIMCd5ElsRR/l9yPixvxRstX383G3mbXndsJe
+1BMWzKUsvBZQx4Qik87z+dlyrmCDQ7JKEzrECUbioiQIBxNdwW7bovUjufJFxaF
Kfu52FlUD2ZbqgJp4N0T4bra1fNVoSIdtYQMmf373KctuHLBnup6PGpaUrjWNE4o
qGhFuYgqqI/N7si6IfRv7nBgpb2b4wwanRb6Gdpd3OsaBLJ0sgQyzx9kQfqdlpus
X1lcpVm15Fq9JvF4p9AU32vfsyfcl2qEGThEpdOlxdnrATWYPk2zlgOFmoezWa8z
5pTJTzytm11bTHRFsBhpe1XAT7SZ7OEXV7Z/2dhkqwkrJC/KI9ku5ct9RvLSyb30
Ke+j07m1+rk2Z0QVuX/nBmlOzrTXDxmsHaFT2i32vKSxPA4A7Ja7QVnsTbYPY/FD
bEUkWHxJP8Na0EpmVGDjkvXTBZwTv31FEeZwgSzDldvcEVcz5eW5YUIKK0mMDVJi
K/PkfsiyM61wmSQP6phyRjZnjkD5VgSb7I72rqNlouy4XFCgPoNYQZUR+mB2ntsQ
KsBxUVhhm+VJNmZBiRa3xZqYgxIQ+BQllMCjbcoHIQ6Kbqq7PMU9QV2sdGTknF49
2pWC/URD2L+ARxQGDU3BU3HzcyGSlUha5hdFAmDfpKPUufl2oaIQVQWYYs27UDuK
p2F10KTocf4kGqGG1kKJTtmAFHG5gX0WSsV4UTemncN02Y1hm47rRxAC6A6CgGNN
5syzihNUBDopwj/1jXJtToDeVciEX1Gk68FgpHMRlHdt7K5T7nBOYTue75CVGwT1
M1tkD+0nbYz73e7kKSu0un58BVlOYtBX7/jOjSqF3riX4TOaLCtJZwrKFPSi0/jB
5TjR+r6PBnzwyDBzUbCe9aOZ3wxPUR0qQ14V980EkC7mnWkDFMYLiWvpiePGTpsd
P9iFPiuwKBsapfo/EBigCes+Yp4qt6SFM01BfQLxCinGsoNs3fx9BcjMLegBnLjf
tQZWUule+JC0bnFXYrwC1g7SHevyuhcXDG3qiSVwmEwh08opb2ukC3EqF6TrsrIe
cOcG1kF4wmDccHKjOdtsUEj9f294JTwELOkeq6UFqf79dXhTj5mxxP4j6UdV6Y2W
9vOIge9+Wyr50Vn2b90gLk22ETFnLlyw3jxB4Lsq5mVxEzNEfj6wvbIaGrdQhujM
IF3R0KPvWWvcpwBigV4Aeycb8f+4Rj2MXMG6zU1jn98rJHgSzk2yPoC/L4n0QX5P
fOBqRWaR1U0DxG6WeLXJUZZTNODo+AURlliH5QnZZPLok25NI5Uv6lq3TrWSeMeM
RPuS9FC8GyBOiAz0mxNDtgjtCYQa/Kl4IPrgI7JMujULDcqBnkHwkENUfkVNZSiV
k1s/Gy62YlkdG+j1KgavHKnppSe3hIqfZ7EHHDqhr91Qe/KXsb5h/l96b6ghIuIs
eQ9k1qq3emCyaLQ79rQdgLuaFOj8uZM8RoGJ5pDjQ3ZU0WfXfeinEW7wN93vP4uF
Q13rVc30Stc48z//Zfx5vC6gzKK/fe1QeyF7XjOMjTcf6P2Wc+1TjbCyq/X8zDOj
H/DPxBkcIlbY0v61gfvB49f3aNqpPj0CC4had+mNIZ3QtPloSBbsefbCtKzzg192
aIrGAf3JFNS7Y7Yv3AUcRO3FlkPPBIhILISVAPKYRXqj9HStlm0P7/vNv4n2vS1p
Tdsd53Yt3In/6/Hcf9T/L8f5hfrHnXaMLtrLOxJtwv7V3AS2diLCjzlA7ipb+MxC
DsZFsu0N88xNcmY3kdnTQ1Ny4xKMYhjUZ3WdRYdiGMkPmLBu8qmCo1ei89B2qu8H
nWIu6nThZAliHKnaW1gNchKBHoaoMbxcmN/tRI9oMZ+cQcO08MPzOL+Y38Ne+gbb
GFs22QdagbeXSIbCV0Wo7LxZD2rPUCB3d5LWuGCH5oxjFo/AIEOEBiygRBR+4egn
0iUmPEdJTYBDPsgRefE36QxgpVgBpMam/WaXg/jc3e77ii4BsLvcOmP7MxllV6Pc
R82w2mHE3xHExX8eVSgdlCW9UpVe7yLSn8rwWnAUiDFdf/MBlHQ3/HYlGNVL2Gev
BRW0TgfWWfultDxLHgA9bH+S86R4RDvW1j0YmwLk0WQDw3yElqlu9oeyEebgEvO1
jqM292eYRmb6g+LBCvGdOWU3g29BmIzF7v/PdhTq3ywR84uNBLWZMU1CZ21a2crh
ofXMsVlZ5XhC4fMtmanuYfTW0vx06iPY59qyaLMi0g0q1QJ3vf4YHbA6Q6UBsN6d
Bm+KXmrOa+6SjpurcaJV63fty7M1p5zZquaChEmPYFFm2PnoFSZcMwtcakT37xpV
e7M9K6D1uQfeQhPD4XYBJ1V/P9C/WdEb7oIc51XoZfcgVFOieuLSQdrmH3JvD+IW
vpQHsv+T3GOhLmhnIfallzZoNLQGcXoT3vjIS5mCX0DxyPj8bztNrorUXi3fjqv4
w7xe2hl1uLb2DvN1OWn/UqdbaTh6/990+YCBtwQfOWMTR4HIwil9yFLoi9ptVWXk
dzhEGApS2wToV7T35QhCcKoIS0QJzMlnp9Fey/O4K6ffh+3EMAyYAXN/eWwlz50/
FO1qOPICasm6yW2rlmTYjAcL0RZ5R+vJNm4jFWNAZ4DOfiL929YY8FUNaS1Szy1x
st6eE15Xi0Iu7LxQo9q2jYXqlPRG331lkeI/eCwNx+o08Ff9x2VH+t63i6rGUCVN
m+LbS8gYwiN16I6TpAMJvRRxwRzD/aJ5kOPF/AbwGecEuRu8E/HgRnuilMkhUTKR
xcMN5Ukj1qhuNeopn2Elv/yLHwGcZaLjdTNK94ybUht1didtSPwvN6Xc9mI/I7XQ
xV4hiB9bnDHEQt/+p7u3d8yBTefvt5pw5YvB9e4M4vIA1BLlcBW+Qfm36UW9FD6f
AnoTqxgBkkpTXtT7PK5d7PPeP4oA4dF3es1Nlq2Q40k+pKB2UoCBUdTmHm5HlOiv
rL3FvikBjbcJyzLQVYmQL6ZcAZC15h9TOP4laDLvXir1dvCXav7yqbGSUlS4LUYX
wA9rnKVI7Bw1Ansu6uBBzeV8AfP1xeKV5j6fNBB6uUjFuVkZUaPv8E4EO/bzXlxt
XOATiDvsztT+Dpcx2hINFu4LiFxLoSd8RVJBgMwy5nPTH/Y1L6ZaIEC7z7QaZxKq
zz5Xzrjy/y9DkuTW4eGOixZMRaFJUHNUVxKf4AaCORnm/IqLzU2Dym0mXNuiEaHT
v0UgUhJAbdFw17wJEFDQXi6VHZaxaxzH+XYnAVYyBPHh6QAR135NaXPsuDC/qjsc
IiH4mXLk15IXtAzHKSGVUdLKsmM6rhDr+KxOeZOQZI0K4PupW98Q5we5xE2qpYOJ
UxbwH2rnODqvnBo3fatp9WM2X7zWd14D/yL0sIVJ06rTlkWBsejJ+9LPQgtCFz6+
SFda8HnxZwahF42yYVgEyS+NlzvrOZFlBtkwUcFE3O7hQ3mr2H2QZf8nYceV27rU
BvPI9LAUYbSrxDDqsQKRfudEDcjiQCOFdI+5fit3p7p3VsRKKzrvhDUPtTN/kttt
jZ0Og22BBwN68hDs52J16ZRAVGtrHujZQ3tXZyoKRyLasos2od/IoSd0IQ1mdtwg
2+rOIxBEeMdk/c8LF6hASYbVi1+tJmoFYbA+kA3xsYeBvN/dlhThmFG5oVT6IFV3
pGN5UniT+0ogFVnSfwWSq3ZWSvHygkIGSFsYKbrWETUoH1G4U6r8yXjDs6blGNHN
T4UH7vzxx/+sch7jh9+YcHcSDiM6Tm2X3xaKghvXVxkJPIRhjgc23wnb8rgipRfD
kNJjJmW2zx4/uwI1LRe+7Ke531IDoNAnh2x40ILEjHRGIVnJy00Kwl3IRFQCZilN
GeJszM3ozGksaFWsqxC7ximTl4xjYmaFdlKq8swfRCYxqZiNmYCbCG6lsdCaqAJk
Z859SpUFgI5ve68TOomD62idw3olNb/RTm3AW4GsvPRn8BA1LEW4DyY+eROYyXLF
5UUf8KCi6p7buteIBjTbgy2eIv4wlwAOe1vKa9xVbV+paacazNQcp4jRqwkO7leT
kcQaq4T+8VH/BSDz8jgk0Zj+U89klDjTgGEBLCLKiHe/+B8af+HwKSVkS5nRuJxw
Cu71nVHeKr7RwHY6B9cdeOgD+ZJWZLmDg3AVTY3kX9M/fnuB0xpkBH+sthc+ocjc
/YyFP8eOxPSF+BOrvFRHEfWWCo8hvWdYS17THpup8dWJDexyFEm3irHe3HsQgGuX
xOS55j/9Iv26jtcVsXwlNlCG7F/zRmCgdwzrdLxOziTYmT/hXeVkkQGuOmiU1dfD
6vtc/NqfLx/ofGrgGLvTpDPZ9cVw4DOi3npnNRhl9e93JPH1K1jmTof+CPfobTLF
yNchLzw0YLGowyrEMF71s2S3en+tJ1htcii9Kxi51eA7wtUCTKvfLTZGuF1WQurP
qf6B+Yu56/xvSlYdi42wqfNS9YpmLx8+Z+UeOb041YF60fPcX1YvuVoUJSA4JbDJ
PPj3f/8tOE7DEmlofHiKSujyoOhyrTm3u0y/ED1i73fqvdEToydCxaZEgNFe0cjK
CbxxNiErwaq1xZCSe7KwQ6SFojan6S2n8/0H91qUkKF81I3EPG+jVfLq+MPYqwB8
VKzwr5RUxmYFMG3+jvvSbyDERylR8SQ/lWSoiIwEUB5ifTo6Cd3Ws+aGhwONHI/t
X6ET892bfRDm4csBBX0kI6kj1YpKRJnbyNUZg48jfWebWGkQNv/1JR4Z0vsNWA/1
2p1/PNfjXTfHj3XrKS852wntGozdfOGdfvbYQq8BIDg6xXT4Ho8MwXIMKgSPWiGw
AVLtfkfMrlIDG005y6J4Z7xUTGCoY+ETEoLERyr2GUsXIWB2xUnBtS8ME2P9Ov8j
jBLtkG2Usg4DSg4+I8IzpFYXfrimEAc2dLgS9eoqMYrthjEfWrO4V2cPPuyPVq8u
jaav9Ca0p9fGdcw/a0BS8MGmxV96HSnhDlYtgPN6ZaFHP951g85bgYiSOn4Z8sNM
8cjaOpYo4TabkpaaKnC1mWBda3iPhGUUN+xBUwfgZo5yOjm4WJstHTTE7zG6p8eK
xXm5IhUFecPG4ORygXR6mgPHm/J91ETzwF3JvulcNDr0hxWUlF5VVXzZmiNsOQXG
7ceflPH2uLPNkftc7UpThS/hO36d/ghhAMdonATZ1gBGT8AcRGR3uZ7lZYXfVdxE
S5l0CWcqEUQwjoSD4Hj827kP0yruNSevUQZfzd4LO+kG3yuM1JWhGMh9GTrExlj3
xASBbWTIUv+OcosMkWOrfoDabt0pTQmU67lJpbKxfXOs0ixvRZwVgru5tnXHnv7l
W1rPElzvpZCTEQOmZIfIM0NHdcw1kdSP+oZBMPRX1Fc3QUEjjMx586n/0kvn0qZ+
R8AWjKz2v/dJzrZHrGwtVvR8q21p80xwVMV92bkdGUrFxIiaQBi1gLQVcyXm75PT
Xo3ePfsQkAzg60v4ZONPInhgXOf3UJNJqKMrVo6kvspO3pREv7qYeKiJYxnYAPNN
GaKVM2ExVLO294TKoneD2TSCpoT/Ji8cOkMaT5an1QSNU7PLwiEvNpe6KIkVi/Ob
dQ9saTFp7GuhZKhZTulTRmFho0LJdilPHqvClUKACiELVdtAKk33BNYXInLuPsw6
jtfqhX2ic3Wd3jNBaLZLryk2MCgLOgYlIAtkBiAeSNwQJtkY0wJ8KAxy6JwXhQjS
WnWi12skXXF5wzDGVHU6X169NxoYAfoYUirE/L5UMD4tEEFq2RTYxXzebuwLx4Fo
hJLlPTvEAybpIeOfjOHdAoa/dwmLPTowB1V2dfirZ4zzQd8O1Q5R7RIN9XI/x6NY
E86e+AHBMzFoO8KNKgFH2TMYCjEZH3wWexMnn+zux3JULZdKNaJ+r0sbvdD0d4WO
8fmQs3Zp6WXXiz+rrTwOKIC2DUHbMaZqbKUHImaOOmDgqUikz7hBYn/QXbCeIGlI
v1qP/TMg+0vGFuJp4tZRxHKn/jiXAu83y//rSjnv6m+XBU0Hpnv8usKf5Loh9ClY
qGgJzXsJnYucvX0CoC7hOisjBOr2odHnORbjdpRETZqENpK2jffENzI2Gpfa3XbY
dvQolqs75xE0ZUvfBysRnZ4WxhKogD0GIZ4NVifuJSzVPnvG0mjg3HrP8K67Gp4K
/9312JkUZFnE7DcDxs2DCBP05UtUdB2h/wkx2yNdUUnJwo7AnEx0Wsr2+G3cUZjV
/ZQ/axBfb9fsBIh3P6DsSOVDQ+4qNlkTw4lsb5QLYZFuOG2vucOs3JYBxVH1vUSa
ZW4UTFldF5ldH1y4F8AWiomROA8C7GNw7YEu1bGcraHcmOGllRm3yVKXMQ/pqfxo
sQfJJH7bbRLf02LX0skpOE4CtQLHtEtJ2NAx7lrwjb9LwRyIgUxseF+k7GeVHE9d
H/xpPia5Wc7OWUCecDd14D3SfP42d2W5SbKyirFqsOrqaOLQBtvkLbn1Fh6FCT3/
ptWSfPO6aAGEuPCqFmu1nbgRX1br/NnDw4+ulxkVPGpLUzyAALUbhAV6nhukil22
hdwukaV5QF8BYFM8S+wImxycZxutS8md61nAG+x+UPjjIlr6bDSdEfhjZ//d7Lz7
o0i465MxKmpdzLCyVONGog6fFGMLG8W3ZrcpIr1uS5IN5uQDVSYwRE+orU3HE7Ai
8unBQtFM40s4DCT7ZMhQJcVqMWCJWesDOWayvfEteAdeBLINGU5D7iAjgexGzy5N
vwTu3Cb8csL7G8w2Onq/KzQXqlzd4SvFe0Wo1xtZTsRguvQRG0s4ZQ0dn7fd5KiQ
2+so5+YyEJnKp9BGrI8xX1bqLhAIPFg/DoFIiqq+PxXRscpykHmB6dbpN01S8Eb7
JiBmNKpH/Zx8/S2BGNcO8yJZv4OloRe8+K24bsbHJ7qxLoiP0hzZFBnNhS+tLelj
m/VjvXO+EdGTA6FIl7OJCXqrKPi4GMyIrrFqm71sUM5BhgY3wRysk4yLyADaQPkj
7b+Qv4haiD6CTPrQPx5Qk6chUIP0quGc3HQrytlUInd1TKq5LX/b20YIOzehl5h2
LBdypA8SbtwR17ycs2HKOOwIwQUhqcPx6Pjaix87E7IAvhXhlaAazH38PUIdFEu8
Td2crw2RN/u3T6bVwpNJ48YrNV/avWNIOtJ0TWHTK0qunYHa6GljTblrHcYNasHy
5H5l2aXsWq+TPkXxb6OXFzyxM9KiNwCG/HDJ2EiTYlKWuzv0zQ/AuHfscn54pIBf
3GWByeTnHzB2/MCeC76BS79AddJojkEhZDkKDzrR3SdzitIiWgX46GpHxR0GRhD0
8o3eWyKj8QLjFS5S0AgjLm2ymBai7V15YLjy/stCfuU5TfwMF1EbONs0eQmOyoLG
+s0wd9wclpHDGxPG/scm/BVb7tfHR7k56quAATKl8LVtUmcDtehi9yGVASK+yEfj
XuKrkJBeD/4pNN21rQA5Wz/W76zjJ/ygHIJrek613TTrBFOYINvx+uq3tjE4b5k2
XYw5qaaOpQJCt0+sK4m2Z+6swunXR38A7aO3Dacc0AUDaqW/zNZLTL05yfE/3RHH
drO9y4L8Cu8qrIbeXblUpmA/6+bUk2XEeSiktWdwtvRgBPgDLnLu88CNmpizhT7I
3xp085wiJkUfyd8PelaX6Cs2shHnKWDFMqEv1LisAHXVSBaKVjLy9rJ0ptcZXAaj
ZxUCmRRMjQckHHyFqWTes/I+uNfv464ds9oACOGa2Uq+gWGHbDCJHy+xwCRD4vM6
kZSneZjR6NcBz5kMC0DdugLM2oJJKlF5IfW3dC+iFHaKcCc7whHSnQK8u7+GuwPe
0gRZvoRrskzVrpb5B3BozdaBMiMa7Z4iZrorPfftMBDBYD2Acx3j4XcaXDY1SKjx
bNsAUf5Ej6zeZrvPyZcYYlqy1e658+Bx6/Ej6t513KHWoXUNt3I7JPJ6DskKzmCd
OatAngyodcaZF4vBS9JnWzkJHK2s8KzTOh4ANVsVntaBkHDFEsD5C13LT/jdaR9A
3iXchMcQUNinJeOYvWGB3wggcHO7xoNAgdnzU5Tr65Hc7q/H5KjgkoMjbOkVGCE/
Yg4JsV1RXCK52yUozw5sN30u29GfeyiQ0ivXMCUK1nD5gP4ZNOnbfX6Cqc/U0tQT
+bJNuKNiP/Mn+xMybghJjFmF1puTmVsaLXTwtMli06YhUpcTeGGsdIeoo2nEhsI/
cydeMn2qItusxGbO8eJCEqk9MtTFLEWrbTPsc/pHATcH/t4/LotOYsrAd9CcZhHC
KQ+iEeC3knFLSRbKy42wR0ILvC/vty16+uWf+WAAMkAfIG03sWvJ3MXKuPPZOBNT
2+FlZP59B7kZ/CVZ9mdUnVngAa6K0qlhyxuiGE5cqwc3Jv8LYq4YxZPtd8soa6+B
3Pj7AW+2PGya6VDMct1Zl6OCX1V+PEacSvd391jm7krPUnNdo+Uof5Ive+bAfIjU
NB+qMao+lSn3X/Q6wehsb87ofo4m1dIIA3QpJzFpbl5KuVjOOmXPL1V+zN/V/Vh8
uFzsqVUDbU9BEyWKOgXo4gnsG2tcFGugimK+K7r35QI7TfCi89RBfEwcC+pu5QeS
F5++/QOSJRhB+9DkbFbJn19SQGP8EqjZ44oiTUk54E5d+W8HjZ3waOzF7sM2/IFo
dh+KvVwRDEv6FZNS9Ey/63Hs83xQtu4TZtLP/akQKr9KZywhYZ9xamzGsDDIrZTX
rpKUbFKjRDyzNKdcivynNsFw335lPnYwxfpNjkA6aIvqzQL5WKbVe8jJrHtZF0hq
t16WkR63kX6vY83jKcdMFh7d7YMqPFnKTu67YMdHdYoomJ7C3xYkWvYBN7zxES0G
mr3GXeCDRDIOfV5nLK4jcXkJHqkAcvKTUybvZpQB6yXlrPxWfhkiMk1X7kBZpkAn
J3ELtJnua718MiX8k6xdJ6XlrPRVOaHnDnzTgP3X09oC6DsW/Xv7zJ5lz1EXrkye
0gar6vGV2CALKuEi9B4jW+3zIUA4SufPTpsb3DyHyiMHG+o/+V/KN3olaD1zhp6i
432+a+/AqsI/vO7DxiAiNDQQiR2RneIKsdggsdsOe07I/2MqhHM6HtnP3bQ64KCP
M2QZ/DYOpqHnHRbjrSiGtc0F2pqzZDMIMvY65wUj/UItRzDxydKeA9rYg7bsvkW+
6atY+fce1gYT5mYVgqUF3YLeICgkb6IyMdfdlflbh4aLWQdzhRdUe1Yh0cXUYahC
FG+99O+9BlzL/cOoXXrY9WgccR6VxVORxn/7hS/kmkUjT+dMVZNpGzBt3BdcZy43
g0li1nUhqJgzhDtWgOazGtwN/qdSSxBxdioxlB0foVtRuWXYPR5TbYNswggYMsYf
uXTNU2/pO1+HmmYGedu3iLeWipqUzYw+sm0EQo4a1k/jObzdLd9rShL3/HPNQUgI
HffNZeuswdrDrC/tEDTYhcjyZ3TrqJwtCOQQMOlZMoMVxjoNrIQTR8aK3QAu6Pt0
oA2nG2xsGXn/POZlXT4ThO9o1ltZLFGjBMj1UyioLePPpHx/v6b7cq3iqUfhadYc
lwM0xJz3UKHubQLwEkgWDYTdCd8NK+bnULta0GtVJZ1Q16+Vb/VZTME+fUtOWZqo
xxn7nfNCokI0OzXGxIosNeNYd0bJOd9d7Uhg3K3mKWJ/irVcDcn9ocYVndXig7tK
yUD1HhgC+kIw3E+RdUVOvAvq+hstTLBeiub/Ej8QOkfgCOb90tTK7fdXZlPFjaUU
8Rmh2UjiFl+JmUxDfZxT5DMmYAwWxgPRfXLEzgF0lQuzzkZ4KLbLU9fDiKsFxYZI
ZCq4MSF68+9LjBFwRpRuXy+k85D2y7edX+21ysvSx7wbmhMxlfmZWKrijWm9uSmH
RdKbMIfh4aoHowvOiswwkP/6eeNGdHetEgzGTf6rETAbnJAgtXBZpGR76+jyqIcz
WK3l0yfIHF9EPVLVh1aywCzh3jhBU/05L+nujdA9+l1piYv/CtSwENe8OI4V9uGC
mp4Lvb2JS6UouJdt+1rDbPaVEA/3q9z5Lgi8etjQqgh1GRPughhRygxiMh+ShNgz
UUS6gDEM4UDPXpI1NXQDLs9CB6dufRcIDYydgXlGtXALw4vhAOCB/YHp+zfopE29
g9pdHPUXCN3K9+pZ/RTeIAIXLXPXVEtpA/2lixlS6kLJk0/GDzfiAUrtcPcMthfm
oeHfszapL+CcF+5RxfRC23lVHdneETB7w2GnAJZbwdk7GddAuEIwSg4haKlasS4s
oqPWmHUPjl7LXxfOGqNkKIrjbQVsokX6kYZsLg+RTF/Nx4wekzjJRYDBIoPx92bT
LFQv9Ovaxb9ubBCIPM6epf7YaYNveuuqqoSkec4XNmDBQ9JZFRDg4/79bRVEgqJo
SvXiqWvfzyXQRuZSRF+DhxrjT1rW1Gbb5fTJ5WDv8szwBr4gyJiyJhziJI97OW84
gsDd1ozDceojXRZIU40BcHFDJMNz1cd1QSywt9yLhBvgmeso/urcoTjyh94crCBT
GNMKVG8AQxWPd/kU3hSsiU7FkIhObvxHGdZr51yRkoniRC1FR0Zo1GhuZGyc7OET
VWv+UWvACaYi6nlxY0ZGJ+9LingTyuO6x24UfMyhD+pojfZVTe5VzF4xlDbr7KCc
UmqssJ+QRc8wdCoOkUt/atrzrDxYGuK/Bfpw/OtfMTln3aIlpXE/B/fufSFF4Xh3
ECtWns1O2EDiMtWLkrJWCkdHJkloRRGpj4wjOZ4yXLloL/Ka9c0HQYLppSyatYy6
ZNw6Qat2JmmLfQ/dvor6R22SS5HKCiusOlAcZb9aPbQgwvdA0ISJr6l6B8BGrKNA
jqRDj6gBMMDmjgdVFSbafZmnmoU+4Titp2ZYVkStW4hlxfSM4jCVPgBejKXbaf+u
kiZvRBn6/Ryg2pAD0DUcTf84dwLWYzMbhHLlbr0kRXx2TcWXpn7qACuowKWBG9KM
PmglPB6DrsWcrKQTfc4WSeNiwEX9DdPSw5rlARPh4RmAPzVGismOqna05Pn+/QCv
KtwPolkPD+jvcsNHtvT+RZLuxMb+DxbEoivBmee3QLO+Df4O5DGVE4hSj+xEdUB3
XefLninlJgoXyXaJacgm8SlQJhq5a15xhMPSU6kXROJRsdjnYyBLz2dXBI87pK8X
pohIjnfEgE7DZ2/nskVQNXJKCDB6XBUQj2U8CNtEpowh57zrPEnB30b4RIGafqum
EtAO96OKR5oTUJ0bdT+nfZh368y8jZrXh2opuiev5Rm1015H26OlQFy0E64TaA69
KFALeVEcBK1+6xCy/pxuh23MVlSW4GaVz9y3f6TmGr05WFRR7KyW8PGkInsOGutU
QDpBpveWr/fANz9CGGZJhbxMuUUXyDAKE0fj36TUH0YJtk38R/6LCTKe3TQwmHqz
yx+EraEJWeLh9g7LxaElA43cTPMmiHb9Ya43Mo7qSn8XKcI9zcMHW251Hsc52958
rKRFoF0sVSdabncqnh/uGREjv2Elv+Mr6lNxTSfzwvvL8he9cvCMru6endz5L5O+
oES2ndr8styglYHaT/3SWBHTdCTc7H1ETavvzvasZupIqR4lPqutro4/vR05rXBj
nK9tx9rj8TUAVonBXiMSLxsFNqChr7lYm683+wIZVD62Ou2P6ezjRX4Dt/Qw4QnC
0EtfNQPXgoOsLhnZWChaCmZO0gb4+fdQyxvW0YuGHCQQ19GIiSIdDM5oFG9SmMgq
IuJzAY5wJILrUNc03RpstpGO0rIi7FfgJZBqEd2xUdDzkwFJ4UUfXzgTdqhweVcx
zlJlXG1ZzORyfBnh6I1v68LuhkTWjLxU7ZZwVkQnUUQ097zSUX4hfFkFWrz3HiWj
iErKdr6QOcKpCFm7Y0onFqlArTZq7bvPNgNLwtXlfapZ0HedfPVlxA25+KKLyB08
3lNpLpVEPJuM4JEJvUwXPLGrSnpT1SyeUIGcrnLgansForXvZNl1YehiMSe5TgnA
rNaOtZaURujuiy+adoRJ3/qPtzNIqDt+T9toiDy06PFMsyHHLgshGGRKNOBKsAXY
GJr/B5cUNixRGEECG4NQRqeZVgffhdv3yDtd6M6csIIj5zn7NiIupi+a1yyfwD+v
owl9hIEmJwoKUKoYGRZ+yBE6/RwttUN2T3/rRh3eACs0o2lJurM9KOFUpuD4B+Bz
ZhM9OnpiCmDYoOSa0PBxEGjp7oowfHHRY5QN6U2GChue3mqzjtQ3WpM3y/STEHak
HvTXWrYZ2NEy5HOuV5pJJ163BXHe7mSe3u2OEC2utiFkOmyEhvADbE0dHgvjZSeA
HTbVL7K0o7B43J7XcLNTx/z0OP7eLYwImTzHiMdx2YhmG0oQ70NuPLTmXQ9JN6fz
D+VqzQ7ylbbbT+12ngq9FEfZdnAOQ4ZFVF8uCK7AwGOCa3WDCuwvumhg/vCIacY5
V6DxY35oGm+YOqlilwH2kJC4eEYZkUD08BI0dkgyI5kXmq8v+DkwaF8iOFLXMfQ9
ABzOKGNikWqx6kyIxd3PDSPHzR2KQ2gZbIzxj8PUUs3R3/R8S+SE8AgPWC/tV64O
4jplL7ZHXUtwpzkKJVHG9UcK81rq1QteFej4BNe8kenqyHJJ05QNyKu1cyvLB9ST
TQBvN/DWqqBGeYocvs5svizPlYXRd8lyGKfw0yfJ12efJezOzCmZwnYGGAE+H5MD
RaSyC2Loc9QhCS7mZCxibyApdc+/+IKye1q+mKcCC8IYPwr+H2SYA+JP583h4bPY
z8JjFvwLih5ZHio8ibFNTunNHxcMnxOE0IgmMz8NnSMUWqp38zALsSDa/Tc12lS/
t58/33G9svT5ZNeXdbuYGt0Aniuvz8vxXcHsmx/ie5kqhCf/BhFkXA1yvTGXSO4X
p8wJmhhosQt0nztnyo+RHuTyv6XbeYjajscVe9XaR1nRspoMRhqW60s6j2+Cj4Pg
XeFFfZjWkEeu65pSA6188QfsSUi+DLr6V/MYpYSpKds/O9bxQ6Yt40O4gqlWjd9O
nhD3bQmiNNZ+AJDHr4vzpsNlNT2ygOfLdizkzQcQtNVHPDpXvxUG29I3SXHlx506
g4pVFKBgI8L2RI9VNmO7RMkd2I/opQm/w84n2ncFISJ39moQLO6ZBy07Fr+iZ5yE
PrCmnqROvrLaTXGDDz0pift0Qq8ff+ffF5UthtLrq3JFs2IvHgmE+RZJymQOB26X
+aPyxo4iuHuhSGHdC50bNk0UJeAklN8SBJJ1fCK3lqiq/GNB/oXKk28DD/WkxH18
MaeqOoDY1ph+iqmo4HxyfQMx/oTgEzrqCHS1U0tcvCsU6z4XXFjU2maN/9C+dDG4
QoIYOS76+53DLYgPh4N0C8G/zdiCYgRtpIoKC/AXYhnUBXpxL4Y4WpNhdtAFFuW4
I5Dxty9D/QV7JHNc8G2k+788Z7uOdsWlEosFpyhax919ou7D1e+aDbS8D8eF+T/k
l5ij79THOIwCiJqZjDSI9nrG2SdoY6SR1k2buEZJQVq2pTIaXS4pspvTpda4gbpq
e+x2rpfLogYfs1cgXClwwp+7Cr4mkRp2vdMATM0C1ULeyXTgMcgxqNKDt7Jqn1/q
q3wlajGvfCXeYaIjS67nalUugiQxBTkSvRxwQMrZO5ncrGuiHlVtXp1cVCYvtPtc
zTmEOxnHRkbdgsuoiSXbU+s3GGDAwbRwjvPKLImuBspXIPYbVQrXJbqeP6FasQX8
hsT/1/ExvHyVOcbvlfXoAGc0s79xnmbItpnAUaGep3PiXf61JH+60dzfXTH32lMH
xOBPOQfHNT4rLq1BjM8Ugc635OtRxF49/B96resSY6/BryE1dMPTpuENVv8IXhrc
jqIIeCoUprYSQtiH2/Z5W5Cqr/ZICrv/wP7qdjwI0i5kPeyG5b5GvEpZWl3eTKO+
/rQhugIrcPH96nZkAqAHcKDqNj7cLrQggmpAqzuVacZ3rIRrkAML2n7YRP8W+lq1
s3mfes/wuMsccE6upek4y96MDdTyF6dmFB2JuhilkRDa+kZiREXflCCORUhNQwmT
ak3aKpguWFiUxUqEmGIbxnDhh8jG+EqdypxQszL8QMmwOyRmpu02GrNN3fSASOBE
KH4bpa8tQrjWg74MPBKM3nFwF6MxdxGWohTRjGOnGoUGqCbeWoP5xdX/ZRTuYAbm
LSQiAivqxM/wD+KBY123XZRGrJlHkTlzAtZA4sWciqWoK2rMpa8oRFRNsvXj7Sms
QVuj9Qbp79GGIZjRfRVL834S7I9uAkij4pn3DZ82ctQRd3bDJ5EhmI+CRRuKyYHV
oHcEuH66rhpA6jY8kiu2YhqOp1xTFXxhK3eLUtxsxDfP0mFTo146E5+7qY9e4Rru
ADNqBbCc5s5aZ++A/gmO0pyPsnucflHrNBkDieS6S650EJDEdoGslJcsx3L+Q9cm
BbcEWyk9jTOnRTGflzdq0Kxe7LHDIKxpSw39/L4W8X1ueE6uS+/hGcLL1pVg47WP
1QtW9+Tp+4hfA6nzssSU1YEm6aENcHfubXEhMdgUoBkjw6leVSf0ogWF5gb6Kr8H
XAMijnsx1ILfnRgcXbgZYwC7gi4Wp2pXAVNoCt2XMXHKuKNFxvHCIr5ztRVxso87
UsIwyDHr7y/T2ipGE07X01/ycZdSCN1NPlq7dxr1wkObpVjOugjBSbRhr1wX22mx
OvPmmoUl8VY3bIBdcuuBi9vYdAGGxkWWPqAq81nnNlC2fMTkc4+FOuFHnYlKyzlG
eOIqr2dsvD6+7fYPyJnf7NwPRyKtXu5YRRRNLypjmEn0bq3bQBVpxto+OlyXTnkZ
4ENtx/iKPDOez/1AmLofsSBa7nxi16z66i84GV97euE7E/OHsPHwTBuMZz9LnHTx
Dsv0Btw86vMpV3K1NkqV0mogcPFHTiRWuZDlknejSrOOKULSez4JmC8R2KNAuERx
ghZZ15TFYxU4Kz0lNFhi54EGzUKEdJivAzsavJ0QMHHCa02nNwgxsvX2fuBITwD5
sRtMH2xI3F25FOEYDkTuH12d3oCljcpJ8oSFa6O5hydSd0bXRXfOCvfcktkoMRgT
C+Ww54NYLyJuQCXa+bb94HAnyEDdkByxzW1Z4ReUPmDJD4dQuDPDi81tHjqPhSFF
ORStM6cV8A9LvPrr9ouSuTKyuuQ4rXsNurOqjUSmOZ8G06BNStL5RabHS02a4rSa
eaieLn+fq6qhd6AthEdfdrW8vhnkLiyQxpgLbAnnbskcxy7e/z4a8Kg7cRolmtnI
YMSkFPDO46hxcDAWmebelx/HL6bcopWo9AH3A/Rtz6Ef1vW+I7S2hYY5yaE7EcAO
3UvRERN3A5dOB+v0K9LfgBqLzsBNd6ERsXPTo0KkgFLnzPBecuitukcXF+iri6hQ
pGv+J0sZGeXMdOI//NRFTD00fdZW6vCwg7uYJXVv9VCTz0o7PMFiRWviUnX/Sw3z
H48sVGBYsLD1o/kOMiqVQOvdeZo5TqsZLN9S8Jv7kUwJ6WgmaHCMHbEZHrdqWyzZ
nhxVo3Ww88BWzuiotkjJVFXnGBih6NdWMcOb6Fqpq9ImWjdlV7RyW1d9UV62vxob
JJ6GBu4hM+jFB3B8MTmrThxV1BfESt9eAXbUZEwEpiczfLvwuurGmaSuvqUCL5Kh
+1gujXfGqHwQeaiEJuIpHlizoq7H9o7vGJ+8ybJi0heYyES9b1Xlh1NBAVZBAAA7
CNomLLK4khZD5kydAg3Ttrxwdvg4w9UIy+XKWy8DY/F/Wp9tYGbUF6zZJDuRPFVS
8fYWIaif2MVe3xajY/6VYOUUhZRuEGXx2V9VH9Ub+ZKqfjajCiRdUvO6FWSyaLOx
fU/y6+XRkaWIuSvnCyEm7DOpN1m4mFo2Zx2i/mjZl3w9w2f1kk0w8VFyUplJaHR8
vBdgeu84onNOG48KHzEA7shtEKqFUUjANhQLMjyp0BAZxqbhYUiMjorFDz+SBdGk
oBTys3QE/R5GCVml2EDfNIVlBVVODsJao5XrQwNPZYTYRTxrNOdKirUnHadljc3N
+KCUorAHVoa0kXQa3JA1IYkwGw6XgnUij94KO729hVJv248xvDTamVs9nl7NUkWv
qtSGPQ0OLEMbbIvLbhKQbaye5T1xxpuqI606Ifln8YZFb5B1nCKFU6zcZaztp+wT
O7p/9zKSBs3Mkhl9kTXnZuBVEXgtCAdNORe1mu27AO/47kH10Qq3T5qk9FWtbIMU
QnGcj2whASDkGgZ+Y8zMLMhkamH6Qoice+vf0xFLNS9cyAq8N009oETgDzcm1L+5
NMWzGwQFuFZZNn9H3Bnk/UrNVciv/cxoMuQ71lEEzBWcYm14e0zwNAOn7O0b8oHx
sBdiWoJ62WAImnHAlHVr8fgDQFcA4RjWUH6CV5RYiqMbUSnDmR7kYCFZ0GY7uG7Q
ETgttZ29MLS7bKGYFK9kY1+2lNQtCqercf20fRkAFbt0+8UJPk/KJuSc7feakJzN
RLtb4CHSUXNWPpQSseU2e6uxFVICg46ZuY1/4p3+oXpuH4gaw1siUIMMwXLCVqLb
1y+o621sGnuRDRDsofGTKFSYkbYx2NTEzE891UljWbo/VW4g7X+F/rjRM1HJz1cK
RUST+RmPzBFE+A9kSH/BPzMjtZRoNvzt6FfBYqo5qZBB9ZcXEtsXPg4uBEezwBTK
E7gMl4CS/aYKIWZk5fiyA7EvEbBkj5pCSBkijrDeMoKCz2qBaknyCoK7aG+9+rrb
xmRUoposmPsL64hiQxZ3Zvd3mPcep7tQrpfXrkiFd7AfCDorK3RKyWn2YJLB//22
porhWn1Oygm/v9UTS4hUrDFsoMsGudx6EYDu4uX2SBhgweU79NeqA73DDkz0Kpp2
MvDlbV3o+Ec8bijEh5+sbOizO2HqZuCKQMpNa1cnnifurQS9MG6dqpMUUHS3vwmY
yt33TTeUZHQ+230ua/hkXlFITQqZVWa4k6bMZqY29JO4XQH0RZwu/TrddHT+TUYH
eDN0O1JjboZkVp1rk8K0pBkKAPWOrWUJN112g/qkngc5incw9qdZzrYFZYHdZurg
vuRjP1kxhR5auO7PAkF6cDDvAPBTt8zon3OuIUr+xfE3+yb3FILFeYRIk3y2ZFNs
g1kM7/uCnlUrEZ6eq1hDQjB2iAjqHjEOYTo9ifrvX7gPRmChgiFvI46tpXR+A4hG
5/HLRj2yoyBCG5MErcmzLHF5mUEeZjC08sznIbZ+4Dd3XWQGXKOCqp/dHawEUECt
vGcf6qDU/wQTXiQU/BcWABW98V6mk20IkcEQD7EVqePd47vlw7zKa8ywBUp6WG2L
o8vdC+ApWCLjU6aqzTZRucTrPg7iJEHMoc291vpe0A7HKmycOayDqqBQcNefO9b1
BYyvGLVahgOl2o0+1h4CMMCmVBuoPi3P3YIQhtGow3Q4fTI0N8nrZkxezyYvi86P
mrBkKu5wjcNp61M9uLEHEi5ZQxvbzEEjM7k9N+KGMzTL3c+xm2K9hb9Jv3gCdpT2
DqDsASiGlCf5TfROJJzmhAISUxGxcaPUG7zauqXzKkSR9/pWddL3/XmAYhAp3U30
nHjeVnXtvmaeTpl4hYphD+/D8RjUT7nK62fhPU/FymqVshelfIvznRQHJkfJdzFe
Tv57LluwHKsfo7LcTEu/JTfJ4qs6AmhlLMZ5AxNOHi990TaaxS3v1vu+ClgXMj9m
OgpIbJin6TPZSsC12l9y7v99QlseGDDLYoIvdel/b3yVJfvDuOZbuKWy/PHDKvM8
AhXG9kaP48n9zQ/8qM+zzJ+j2TBl6A8Td7BeP+BD6WsuJNkLqAkhH0yFHe/q0Vqd
jaR5LxnxrsSYpLLbIY45uQLbg0QbCmt5wDaIoxlPK2KaSXT2X+Si8dlzjwb7QFJH
8D6gpqNY5bw1TDT97P8BQ4lfifPQ7suHlX4nQlZGncwBoWeGeObDC49SE9xE6z+N
448hj1/vaeAC0hJP7hm3Pzs0+s/3zoerxjouYXdRzgCJ5QBJ1Tn8Uc1lhhX+6zgk
AB/XCup5/CkZiw9LDj+m8AoobJhaD9Sn6JbQ0+eWe9vIRsibzDvK40stadoU6ceq
KcNQ1LeOjkFtXJj9EI6g5KyvPB3rXx1WdGY2KnDuQGMXveTagIy5i+50o4ZVVn9l
wThK6GlXXP/WMu/56MhVALfTahLZYuu+Vb6kUnkED6GSjUwVXhFhsGeiiXOh1Fa9
WtPG57gSJDG7s2HsE+lOaNnTIdksWEYvOVIChCNh4U6yZcVN4CCOCkMJuG4nF8QG
Mjprjkg+xurtbHs2hNyQcxlI+j4nWC80egR9HULDmEUqiwQAFfP7mY27KulJO/Jb
XkK3BiJG5eCZnF8EarA73hLnaNKwpQHL/aA9jmPCYP5H3LCm2wVDyspuOXT7a7Sx
oNH0B5P8dWW2NpZBcr+PKXZOroFsaF5NlI5IWdpgPr/6yPwe419gMdZg14p9+mKI
4/PRXSppGP69Le98Ac9AUhIm7iyiIc7Ji+ymGnuCCpqx4cb7X597nLdlWXIQg0zK
+kaNUlUSrQ3JQXDnqWfiodkKQAfZiNGAFYgKlw00599Y8cLDpq3N+3arJ3H1uy1T
ZoooZ59AQNCWIYGjt/QMw/whnTm0jUgCyIJaZh3CE4HNyLhlI+ZbNx5Quh0Myewy
ICdOfaF2XCS99uRGclG9ePHJQP5MjO1mFNtuvJJOOWQRfAA7tM+75CBYdgsuuGoe
4TVPBFV0NHVUXiRL7tjG55d+z5KMVp/vFo6o85awc4P8CEdQZM7gYwIdDzVbt+Bf
Jo+8pd1/zefnizXJh3kBT7UHlP7OyDLaKqZLyoRfbsUDSojvtCiXBiJ1urnT7Ez1
/wLbcGC5qksvYwGX033y3HNN8nDS7f26MXvs5E3ymqp6hJ11joeUY5xx/BAhMLFH
J7bDczd75jhVMgabMsGXFLnkMH9DO1V7kkHHJlfWXb9R9fsUvUHl20jwfL7k2d04
vIFvy6HOv6zUSthOSmqXtNUkV/auZU6SgLfNUVgNk9N83i9dHIjV9NobGY/6l98H
E3O6O/MPOOhHbJGCV5QErWF6GC0/n5fAh2Uin9Tdx84YwZ0x8DN9mxzN5tDs0hj3
R0GiHkngtmlTW9Nxu/YKrX6zkc5YNj5DMBMfLGMwAvyQucnYNG6wqqpyM96qvQ4P
nD2GRNFf1dNecExaYmjb4KL9I02AkCGQQE2xmrAdM8YRz1hRN6VPM9sOjWSxJoWl
Hoeg1bvJ1h84tX31GcyKGgPoL530du6dlsRt/zIoST/0fvBQ4a7izJX5FigODaf+
ntlA/Ydspm66WxcUdVV7RbPPJdpLmQruytX5GifR/9VHqXkgxN8SGC1Yr+cJC8a0
CghrjZTG465GkkQtoXDCKMqsDbJ65t2zGn1sPurXC4XMxIsSVSFrsihzR/eoso2+
HJZjwJh2gu4fTLiJW0oS57s5ADK7mdg5AUjEb41c6EIjC9vNTzre81g1NLQTd6qR
9/X943PHE2mYddPxZVw/Ikatv8cPwAGp1S96j2cPhBr78SaO+gztjz+MAf9UquT5
7gW5U6BWtnX8cqq/7xzvvvi/hYGb78YXhwLyp99SqB/KifZEh8Ti/b34Gy7FtAbc
oDKuZR/PH1ZP7Rha1i9rasyPJHE7QEtft2AAXTrVx6I/mXIwRNbgy1gZNwoezbNK
62pNGYjmfBttetsF251QGjwS6mvTRARlIav8RoGlTyJPZfl3eHpsEILNQeXSfdoV
QV7lY62WcTS5wCLvRRok6VYzaQL4DWCo2AvIS9lrmUYVdXfynIM0oXL1uXiGGdec
FIOWAgE3EzCIYW17CT1QRVWHlQ1hmlhM5JkdD/dcpIZRAoTy7mWCJrbSKqemOG0t
ladeyyohWjWfDfc6c3jhk4D6TplCJqcJs/GGuQHAZ9vOymgwWWF0/uKc0AXxxEmf
ksvwlmYRKLyhF54Lpb3i08FTBMXkOuZxqydd7/gyGYhxhgBo+uAyfQb7iUIpf+vA
3xcdpXEy5sDeCAdYXiGbfHlH2Vd908bflP6FIvBePXYqEYyymVcioBdzlbFbD7sD
z4bk6B3/SLKo6a5C4O3LHSI8PO/9vpKom+tsK+n63e5ha++oOYalkfojriclx/C2
oKIgm6gJ88xj56B8B+zNlaQZmgE+65gBFm7NUTy5wksEcppo9ERqIvnNwujXldfU
oYXPujxSQVXFqHPwqQbX9XnIORfNpp6rxMlkPXSfi77/kbLAdu8ZaimZAcyHtrM8
l5079jb7pcuU7Vr+ejrzaxW6j83WMZ5gykuJ6P+/HUZHzpdqZeuODKYtclq1yUZs
GeYvzQj+ELlZ6I1xisOWpbA8TKE2q7XJQGX07+fukcTPOtQADd6yoEFjQAJhkShj
WTZIcxgyMTmJZLGjonmRBWqLOcDE24uXZyUOuLqqugPWVNhoS5Ukgu3ysm4sdW0r
L4cKBGIAwIhULcAH6PqJIJxokBXxk0eL755yxp59M0H6s8eOp5TAEy99JQkGV0X2
LEpqUQejqXfB8XcCvTsqs+aEDkdEddpqmDEeXVJQKp6fyGdB0Ap62RCl/6UxjXJH
CHutoDJQ3L0d3Hx2dMyH/COAmTA8L3Y0GxNPKNXacliLZKWe1+xlhGPphx8DRFpG
LR+94Df+C+FSvI0M5WSO/w/jsg/kOQJHsUdU6PWs4hupIwp05q3mSgT3Owm88+tP
+6gsOUpxD3uc+/dBAvlkccxpt4PBPT1ZNAFWyNTdrfAq9YFqQl0vFuQH7pf9GosJ
4Kqm5nHCcNDhtIBnCixe0gX6EeiQFu0lg9XAzGR2nrpKHPlbVCluVB+hYtth1gL0
r/tVxrH3Qpq9/FItwsJ3t+Rad86FdEdhDXhKTpA/Xo1bNGKpCA2v3+DjIeD0Iv1N
REMwM8cf7J/A/FO0pe++5U2DnR5/yDG//EfYAVMcgmaG16jnF6laWuOyi18qQL+v
HpJvayf1UgtddpoAw80elFV3hwX0DAPJOPlfDK0PyhunL6rItoU8NwKFhTMpMzE+
3CVqgwZfhDbxbHniGKm0KsWE2f1/oOHmXEvAeAgBWOXrj7r++v+BvscER9CW22tl
rulj9zpziSNZJHY1OfSQwA3t6Vmcswc/FS0yBpP9laYj549kIbRS6Oae+2wAUAQL
Z7C8dDAGS08aKCq1FULeCqZ47Cif7wHSGPfV/IqHcp6oVqIiIHXQQLTUx1vTOKFy
Ciyn8oRi2L2WxQHm5xeI2oVnO2D6wgBHKiIBw1U39ydnhTjiay16k593TG2P9UAd
Tkf6uAwteYy8hRI7lc2xtNsgSdUKMJxtxYgFqSdSqIwhDqv1Ln5mXEdKstZ1Eu96
IQPE4gPSHC8fqVycZZpMLPRPQ13C7DRt0F2dCNvJ8b3ocY8COfnm/zyRGCCxplK4
Ng/j6WM7p7RXXAWBvi3R3D7G8LG4Fi/IrljAeg38/DHbrnBH6Y/7f8oMwwHK/gbu
tq7VRm1WQ2ND5HCs1hr2x5g6Gmj77XojzKQIIV1Jz0agUDYQ7QIC//A9K48yNLAT
NqvOBUDliz/vTYLETi8L1VXAEGiDxsOD2OoNtUFUrH7Ee8JKn8j8ob0KVLDkTbW2
Giahvvt+l01/0lH3XiRgrnsXlGsjsKi51bppEOGSy/k73A+dSMRplr+qG5118lKW
QO2Dj18W8PY+6t/Ncm0iYKTawaEFHsGOGlBpLsB/uPwIN9T0m4cpzALfpgqPzjE0
pxhGqcvGI2jwG3+i3/wBdNX+2ZdnuLm6mYbTwv98uaS5iAo3AD5qGq35JwxD9B39
LMRd6W4ZtjkugdFKBT9DSq+pKz8UVK6UDrBHhfE9aWnMDo2DFF9aUAyJ9OoFrO8s
y1TkhfYgG/x3SDfnYwS+u7B0orjpKZIzEEx9xvNjtGleVJ/9PlH3fCvKwnqSJ+HR
elSzEr/gNu9S92/RsC7pGcHoD8VqOe1qWRRZ0vGcyv3zun+Js5b5bD6bd/frhRc6
AgsUIA18vJOjTQ9GiDIoDQHF1+LhI4JjZrU/k1x5cfB2BfaSlDg7FOQTvWkgwlS8
GnNvKAHKITLIVxR0rVWDAVQj1xySAdQC7pira/hBsWyQp9a3rJaaxMhr5Q3VV+Mw
niQIuk9Betp09B4/c7foKlfGgdtqksfW1hfnK3ZixSj+7C9t31rQws3bFLbwyE7E
a+iEPYhoFlbb2J22ujT/ldFpcn2+xggRtwhxQ4rFyKobXOjtGC3xSREDzUlYApEA
WlaOyP85U9FuUBmVs4wXrZUTG0YhKkmDQyuSKE7cmoRfyG4wxoXe81+xc75DURAi
1MIN1roPx67mhJAQQkbxnY5yb0vgM5CqcvX8m9mhMh0kJs5ZHm9pRquAGuTzMXYk
8/Yv832YkekdkZfkaNxv6mzU4yAViQQQ82EVIqwReJL+fHCOobzYVT1qcDfnsZCV
ThJHevdv94r1uj9/Hx1zvofYN2k4xBoQgLUFrOOe7sYoGByMA8dTPzFb+9tzAl+M
jws3hPUEGrKHGnnDs51u3EqiVsTHSnfelfsfFQTVVnIsrx+rBwxDxg2/sD1z/+fE
yHU6baejn0gxpp/HAvsZuTy5wyRNZ/zEWPLtJiiRGjVeK7FY1ogLMejd56JMUvVB
O8gZH14DN/cOYfrLRvET/fPUMlp1UfCClBrOHN4GMKoPl/1hrM1tmtwPN+Xu/dh5
HFyWev7wVpZ98CZNhI8a6kuH6aGfgtGhBckHb5o1wLgP7YVdQD0cNfTLvL0Qqsb9
aNwwlwaWtIW7hrksbdAtPSsHt1z8TjuW1SzKmm7DcaA7dyW1ZnnpM1xUPdkzeuzZ
zEtMAkcah/zTRDjsj2sVzRxPI/xmThes/pv4M5UrjWLD3WcoPAAnALUfdk/oj7de
qYubTnSJ40S8v1ptDmlrbCXvmfL5MS/hjlfJHIeD4p5oU5FZOz0O63DoENhnbVhd
Ejq7SU5mLe3pVA7f6K4xxKbAts4gbizq5LpQvoualiu3I30+F9vTWsl11Jk/7ldh
zGRAAZHt1RxOJYN0zht8hKPHLxDj89Iqc0mI2KbAfHKe+i2brmTqVrOzGrp7sGHv
jK6fQLeeO3nVMGF5HwnvDaeTvU6GmPFo5XD9dzywir8qkzOYnu5J8vDSNnP4tMsS
w/RvpupMYpWMIC8hEFYlG7T25megMWlgiHL+Njelhhdr0iigO8pP4/4JLEnDJZPP
yz7o0yfy4LLIkmNRzdbrSW+OT8ovcPOe7qS+dnGYsEcz6XBA/9manCYjxoC0CIVH
wmo3hTwnQbdMl9i/mpPKzZNMEdbHTI5bSdyLM3q4xX9O+Xv8OWfw/2USjrVtGN2Q
jKgE5J0pFoawqKF/xPZBKWambtAWT3bN4n3I9rcV8QPDthrdMp5ZQgSn8JpMCBKs
foNndkyXsx26G0zZbHy2exeSyvHAvdoGTtyQVcJV7xMuLJ77exzjzPIqHJE49+YL
nH3M5KBRirZzjETF+NW4O/eN0FN9Hj0oogu3R4vL+N8xrS8JWk9bmxEHYO1AkHgv
1+db0Kk3piyzIc6+2uOJ2duc+LVL9Ui6s/I1cFIM/t7B4mI4/8mkWhRzdFYMgtwn
5BlZMeE8Yj/faKRmOAXXJwDHVfOQubde+zTUmiHdwYVS/1e2BEscAQpxsHuTeVtz
IRmcDeIkloi+TEYiuJpLbOHNb/dj2w+389eVzL9sAzjnweE+hLNVWDS1jqWnPL9i
9zx9yhQAQtxYObA8UoSi14X3p35Y+vD6gYoQ7r9dta9bwYjgue2dSvGSOloSu89Z
2xHozenmCoVOAvuW/cXyDbNG9z6jW76uCDb6uUM67reOnypa9f0X1OjRTucrVmxk
zaDwY/wyBgcvGEJLZb+D4yv3Y/WclMwbpp+YncH1zH+CVX9ZyMR3kqL1gdMG4Bvw
qWPdrvHWkC3fuZ2zF7hB9EcQ8VwGzQOshoIaxLfSiR/wM1AiAHw89tkLGYJaORpd
SFbePXDkyCSgdPBAHobXDL9u7R7hYGsdkj3rOVU/1e8fmuz3yK9pE6qrL/qVb4vy
JCNQPQkhBgyUnVUaaXMKx8/caXQAcHPfgSdQWP5xZRFe98w3nSOsQOM9BdmJ4ZPW
lxPCWlStIuFeQNgOiyinlRHhTFU/BHH1GhGYn4AH6czxrGHdE6LsJWsPE+HqE7Pz
g2PUmtrPX9LDhAqMMgC64MgNbqapZ03q69EXJ1r3W3e55tB6dAeWAJxIUacW/R2f
AjNo2MGZV0wdLmKqEbhU9kQbPN8lXYOIlx06sJtxb6TNR+pjhwZ70XdWQeQkmPMq
JDv+45+3zTbbtNlgn6AjeIkXEVpcwkfgTtGePqqsZ0Nsof1dNXNBlhZiIvP8/iuM
fUXtDBzze52S4yKe71AbHxg3m7Aan+Pk30sNC/4H1jFYDnDMkQKTl5gkVvBODyZO
PNvm7OEimWhCdfvmZNGIiimBnTmAaOOp61VRh4n4A51uJB+ic/ob1FPeQCI3szjB
ONRdoIyDp3r/u4iO9l6NvpSQ2EWpHQXk9Zf5R486LYr+tIyIiM3y9rRxlccjDcoj
OJtOJLmYK5cJ9iSTsg8iElG5gCqd4LTCtVdmcysk5gVGHzetyjQuhBeJwhnXhMVS
5MUxvNOIpRe11S73yUhzy4y/fhTeNU8eJoaU5ITkG3LVIM+jrh5i11pFZVGSI7jf
wbDcv9GHQfXfXi8eLQMJ0eLFt1OAt267DZWTAiR82ljx1H4BxPdjqGspycgYQcfK
hG1V3LEqXIaDnIB7m7l4BO9yPc4lTJJP/yCSF/ppIcSSCdJrZZ0HGZhF7+NMtmRx
zoiN9yvBFWLGnB0hqEwgLusCyokgnN2bPl35Qn8Chz71oUyG2d9n/iPtkn9pq6QH
KuQ4DXhpjvCHVWTEjCgWh9TYyLYjPUc2U6CiHkBVhAzfGlG5tnxQvBtwjVjM5/gj
EiiIW4zAMXk1HeU10ugDkGfADYBImI7/fEhsigQQ3xxh57k4tVPO7H2v2GY6VSSE
/gmdxK2niztc4AssS7daXbs8U893e6P4Bcsezt1wJU3OqFxcfiTFjrYhTX9+5pQC
bpcJrgoP5T8WZOOSUfISEXGFCPn9Z1ry+7uRadiFs5CPqt9xlayOJZsho0daOaXT
Mypll7ACWIsAx9Jn/schNMm2NNgwh36QTf2aRS1aZFMkxWfMEgZjZepisxqDKxqs
GkOZ+r5Af4gxEUoJ52eFJaiMDlH14b/CVmR9Pf+vfXgLCvPu5S4perWEs8Ku1W2w
DHuGlA2rZ/3wPaTDjwZfvEOzNnEaZTMb4mtSes/FKBMAQip9SOj7+ixjVeqVnb4J
DVQMHpgujXG+Tl1oCe7+oQMvOon/pssjl4/G1vKYjH6LSCkBUtIczMteEt/Nw1Uq
mo4I2oSSL7KENZGUR61hRC4wZDXOoPJOGFYkcQ0GO0OsAfhI33coNJqelyq6KLlZ
mzTwHHOUT9Hg9J0bXjFxselJG1GwCiTIkDG8wNcM59zwpP/HXiXWZ98AxhFKQQSq
wb7kAGGg9IsuRqYHQnOlh28DQir0zQFSoj5YWD9NvVl2G8VoEMZDefVF8qGqh9Pb
G0vJM/HSJzy4QJmC3rBylykCV7115j4tDqEH28fYOwm7uKOitQQFWyM6ihrvZXpQ
9jxMPDA+xLomlG/PyBJ7zk4yEIiEsG39bJvqbN+TzEoZw+7sr5go/jZBseeYKoL4
blj+owUF/A1JqB1sianPx5LJIorxcsSSAdrvc0Xee9pHOthdUuyWqxVy08ZHMCx3
XTNkVu8SipE3794kIAxVRJuNbH31vxtWhcrJmFfJpJ8r90xcwZD3hHRKujRFX4Bf
Fzvp+QeMpYoyNAy2KODJpzbVKaS3qGLSVOGFXHsdhf9BSCqNVG1NvHsQ+D6o9RCl
aFsfX08CfWMOW1f1kxTwUGmFEeMwhMuq6Jqo/mMrHl8N0h1vVyH72eb6ytdzWAOW
LUPszdxpxmT0NEh+yopDVSmTSOuKuVMslL+MNeHoTlgLk+PKTI8eN+VYeM+y1YA+
T+AV4qZeThC/o7uh2/1xeZ4En1iI9qPYnI57F0blDVKNPWlzboTj2CQ5bMIl7W60
ist1RHjR4HQIfBbgb6fskMHUV6+dFhfa4+17a5Omn+iDutVh+45Hk/vw4747BtZQ
XZ6xGGi0WCw5E11uUfeGM1UVCBdqmJ1uf13SCE9U6j2tcc20Vb6F4jMmfNs8NMFc
aKuem0hWMosylx12uHg7pL7++b/689fbyTtfqKSgowJQoE27T75ggciKoNACNNJA
+vnHYQnaEO9UTBXe2ZBFqK3PjBRYVrNSLtEiM0jkj3tGQu7YX2/VZXFVmUGInHqX
cKhcc7Z/9YBjjneGptyXCrTULXsotGmIs0nReX2fyO8bn1kjnEPx46micWw+Zumo
xcI14CVOCUXYKGAodk2lqtD2QmwIUOJ3J4jtPZ8bxFrbm8Lprodz0a+jnucJX4xU
xs58ndGd801fi522dXSnRXj/8UMlWqwcaxlZqTu5rmJfmCOV7DIPF9EUlNhBHiks
7lIxAJsV0A1RIlIXxpMWzcqEPSeJkyALP0rmZsEgaQrwfrV0q18KgI+kYCcoQ2iE
OPfGwHUBNN55tiEBs192FQoKwQpoBSMQ+M/yxF4L6zjcasV8lU6jeGq/LDBq/nwF
83Ky83FJYobs1prpOwciQ5RAzxLphkgn3lzibvTLtDM7SzWMhMj99+RtaaL+/Czw
4QkatYjTGQ8hWJeV3+xv4z3v2qfg4tLoBojJjjvhlPAjozOkW1kB4zdpYotNzACt
FzcLA8IsGpRDTvzyun6rIg/ByOEmvMAwNOV6T7u8CN5aMYPVEnZHW/f75opn+pmP
zs7EbpP5pPtucTQwNqgmVENVGGgqYeKdW4K6tfSBetwKKWLDuELIrItsZcYJchZX
HmfAN9C8xRA0kxZs8snc0KkEZcIGRfkxtf4qPSjYevPwJyv9coD0sfqI3jlJb6xY
Qesp1+FIKuyKKBLfK8r/5NRXJz+bF2Ke5wJKOT7a1hbrqcsMdFWpZAAB0xOvLlvE
GNzzRCm6gOvkNsf+wbZHaMFovH4EJCcdoi99j2rFmL0ZndQ8M0LX5xlU5cgG1aJ9
i2UTbR94NToB6OSgQZElTN6E1YhcOAC1j8jlDSDQs8aZVNSW9fkqYxpdGaWZD4vC
JRr8LWaVmZzmP1zv+w3T05Pikyp8YxkDmLHTlKIduIwcFcYLiwn+SJfPgnUpheZM
DbLkc739IqAYcN6IG/lUVfFmQjTeYpeO94aFqre8Jm9ZXnc+p9hn7rryFYl755gH
gxsQPqYlSXvzgXlP28ZsYtvQGtrTcxgASXLDdxMw968cr0kCQzvmn0CYZjBuABzA
UXi3Yr91e6Qa87eHCbIupuVt3MpamS3m4cXFcrmw/HEZKyMeCmHUlnZX6cJLx65Q
5WIKBMiBpUy3QDrrwDTiks4DCsC5K7JYdOflXJV48w9gZTW3mi83BwXxQJ9TjHDO
zlh6s0yVrW6b2KMle2aF7FlmO8PMwttZmlaF0n9y3QNSKsxNwd5kNH9hMhryzYyZ
EmSDNiP4AV/ZQJVIE/A7phygmR3BC7mh5QB+llbLEV/QrLzLGk4nyOW/ySNqOuy7
PTt/Tdp0ORpjd1QTBAydBegA/Ob0zlRSNzTrqeKvaXgQtfUNHY5K6PT/OGS20pNF
AeSfqXty+Oh9LgPGnYlNp75PmEu4Kn7ToUpVGii12Qda/mnfCgtH73wCbzHDwLgr
rSWi25N7BP4LaUmcJW6R+blXIEW/ii7+RZ+Lbbww0YcawUpET7Eddow3PS9PpDAt
HAwu9I5wPV1wR3oGC9T8EcJNJ5hQDNWfldD+CJZCKl+cFxtUU6ZXkgJVgGRgDb72
Ck10ChzzWlcE8Ey8Hc9OnR57T89slol/uLsthG9QJgUotTjbs+1s7yItyllqx2Ay
tg/26AcrEKXDSuHqZO6aVMcJfy+0FQgu2Qn1rOgi27G6D++pzy34uD63xbUFpKgV
YCdv6gXbvog6s5PTZzoYUBSnK+cFLOpSgc0XwQYbTm8KpAiHT7mWGoBTuZkbfoaQ
SVe3BWf1z5tGMtzB6VzA4kH3WWwuvbxuvDMtdYWz256umJwy0htJziHLHxF6EEFS
p2IKOFEIrjQEnl94sUiMpJpUAKzvGN2JCoRJPkEyW9InEl3KxDYU+DqLY64ZAqQN
0zDk60WYAY7M1Xg0l3neQe/Vv2hJMyTwOCFnHApjuW8z2IWlfz5/IVRtCXqRM79v
qVpXttpmjHT2WRvvUPPd+RqABzGPqVVp4+bz/+zNQ6prwUfzqArR/7Ldk5d7kKa1
WjLXFZ3gQRJC6BSW3btnpCMdBW/NBtZtnkFWCk2tOyNvB2l7dBTYe19HVN2iU8tb
5R/dLdrpHqLlnFPjgzdK0JtZAlGt0eqIRDOh3PBRJzVH3wVBFpOz+F6SXxnpufIp
dePvPDYWfUZEhlQJ9iES1o0qgkKFKLslHyyoSTdXU24aPZZv6qZK+JkyvDCQyhqM
sD1216L/0abCBbSwzY0EOMfd1Lo1DL94QnTEduSYQTMWafDwhAvgqFHEJrVrxTHJ
l9oBTT8UDtzQPg29EG1qjGy0K51STRuG+EeVvtcu0YfQJj/lRW6WRZPSh/0t3lRK
a1kz4tfLE40QL/A8RlSHwQyDY2fOiBE9lc2sBPAaxD/mQj4R3d+baYAyrl/58jZ5
tZHaFgQ9cfaB/S40HtquykOQP8/3vhLW+1hwj+cSG/AAOu27Kce1DVn22szQ5Ukb
aEJuBI3XUVgRFFiJeNwjy4sbBKDKANIIhuMRv0Lx3YzO6hyBe5M4zmqV5qh6d7Mf
AZ6lFSr5M0W/F9tp8R88bKxrnVI5MwEFVYVCnCsT++W5XyH6vdmFtv9EthfrXPFF
l3LGCCwO5RmxPGAhV2PWwvhVuVVQUVtUU5+OHlFaDGPg4EutUp8iGyodaTvfPSqU
tJpIvcjua7C/lXaGJYPYYB9CArRuvJdpONVrjdNrch9DmmWcR2dBSCySh5Wo2af0
L0D5DynK7dHLEaG9q7yDkkiXtcIQOnV54PIghKPv3qyjdHr0qxgPBcWtMAQl3S2N
7CnqWEZjJcOEt/yYY6ImeAirilRdSs3bIkWlfh3x1uUNGZ0JR09UTf1dimOoE5hC
1J3R/BqamAEUk0SW1cDo24ETPMBcBTCat6oFUhOTq2lSx3bHURwUUSpZEsh+VHIR
WpmzAfMEwprUQF/dQN3y9vp5aSVVeDmFRKuMiaNRz31DtK5jmPBuBiA6pOAdBAqs
Gv/0bk1/3ITNbTPik61jiLom+wSIs7wtddstqeWSC2J954iYTXOCvzFfoK8vFJV5
HOBLQJ/q2haQstMZXdeEJlmL18PJRR5mZDTSwJntMBP2oxvtHRa1BLUk4a6UhCZj
gyuCXEzOh+Se2WtcFUm7fC8IQzfFt+aev/j70P6HtVeLgrY5bBALdQS+HxhLzCMG
Sm56MlMPgu1YpBoRkFSoExwZiygZEMF/dYsCTFC3PdtBRC/Z0dbsKdr7z4S/lc85
ikFX6/MNncc13k0sU3Bj9u6XE8jlbiJ6zW3P9Ys0v3KqzG8GvLgcBBIyTgdnllTq
VfWAvuoxpRIwYYfvUCBcvfTdJI+O7n8frkSH+v5i55oSaofWkmsNVmAEIc0UatUu
Ydve9Zj2uQM6SYsFl5Vi7WMpebMJz0d37QmjQTvvFvQU7Cpt6Eu5moDHTjiX6NCO
0uuX9mQNd2+NUY88Oc5wgfId/8dIfPGv+3toSWTDljt8FAdSvEu6/LDPxU1i+93O
AURkuMg5Gz0lo7B0aDsKe+L+WN3uldAx3jWiaVz98EfASvzHLsObiYkBBZEiEss8
bgZdWsV/15msobXtKYI+UEO/6xMNwMMxIX9GGUk8e6x2LJEcI2a5sqVSKvHJWmY/
26amLSbGenNrPoqKT+4d9Kz76T05EWt7Exq56Bgsd7TeUbp3IJkVZdHpcGKwuymp
kGyaBrht+9rg8KDEJ1e3JfR7XzV79oibDv5Bsy/K26TzI6hF0v0zzxqEmxTLfdNy
mjU0SNDuveaScRqJZ0hTOoy8UjtjgPrGnTj+I2eRasDgAeKo8ZXKflLg4psXCKV1
lPG7C6QYEiF7EaXwJ679IaZbza1lCgzs4VRK6uLawCnS4p2/ZxDyeEIqNueVIqxU
WfL8o+FByO9PCH+azHlxNiuyDQR4yoLwPXzeR4sILE6P+no+AzRhXStYyldT8v+H
6cJmYjUyOPBIp9jd2/pbUzNucB97TwrKfVBPOs1EAAgalesmjy+0cHdWTBENnAhX
yxhF1sxH2VcSYT9MY1ELCpNgNx0Y5jM6EQw1Xn5w3jvI2uKo8gLvhi0ssQV1cwcG
DpQrKDZhLSUkXQUfzBLTMZTlMdtUa0KLpUxELjQsAuPjcOecOdzSN5+WzlCAH0xG
Jkx3tCqFR4yK+3VZtsbwlJtdVUUsC+UF3R+504H+V4wIJzTXfvigue+9SeJyiXU6
j7xsLawbCbbh+rK9RjNsA3xX3mmn9qzuvSCAJyAd3ICrk3VKCDMbigGRzZF8pFY7
Qv8ycNVibSqELJiQZ5BTeNrXemOlh6MK6TsALJQ9JpDbkPSVVfCKei97KCELOyrz
5oUK++3HHeJgiT1PLDvkKGHneUmrKJyWiz9Z7A3ynQZzZuoh5GrjSs1H9fKVo0Rf
JIYnfUTWbym8gKGi0/udXva9Vmuqj28bLgzkreCCWf4YS8vf3RxB6WC6p6onvQ7C
gq5iJa2KvPJrY2D1rwTpQDQSJrAyTkVPGYoLr8iut7EYZZqoQSy+YqPfPVih6NEz
QpgCGZvhn/6l/F+0pS7GtA/5/K6yQvcmobfUR9XzpkJM0eNZstG3L4P3k9IyV2c+
Ruw/iPD4/i/UxVRUITA4TH272uqmAaiTVAXhkEFtmS6xhdcxrcb9pE+JgVCIGpSe
8QsDTXLxJ2bm5gagQQzEChBpUXxkXvq3jeuN4czW/N5SKcfEfCPsXrIU8Q8ysr8R
GuhAZ3vrWS8kClKOImUcG+4czEta4zWFWU0MmGUW52DyABUdQJ01FzkioVh8YJxo
c5ADPds4VBGJ039b39HdchIrjbxDGZgqR6Mg/jZcq/5uyoIzHaHWxygrhlHPjyEs
sXX6Vz7kGC4AykL8NQ2E0aLLpRL3nNiE4w3LPZNdOprEVMfoGmnQT6mmBGrNM8je
luRT75ONcbE6afd+54NfPpNuSfN0PaMtEpR2UuOffvDbg42IrrvtiOPmONfO0XNH
QErHHS/e83x4YGGHoCQvv6nqHN+iQQScZyaAEAIJUUOQWUL/tlxxyvvxP/t4VN5i
KhVK5I71AevqSytRYilnHSR46OjaDQCK0ARq1rA2hhZFUdOvHJYIn3kmWZkHhKfg
hgnAuODRNtgjEkxd3IS6aJVDtTk9X2qIEpdfOIaDvPnvFJh286Ky3ZwyP8uF6A7M
GoNo/ZfA9xWrP4FFPWphvVxe5orzbHUCD9EPYCf6nYrl+BEmas2nGxI+xc83rY2+
b9ZdSfD6+LGjkEhbb1xdrz03+f6k4WYSA6lQdGoS3HIp2Kf56TuHI/Cx2aTXcwr7
4uqiFC2ICMQWUpSnl9CAXp/erjERXy+GzKq8YxlmJ6yqwc8i7vJdT3cKPBomtVSE
NcmWU04SVzuxztWYI88vkxYiUQwSQKXxqTckAVVr56lEK77c+OxunMd+2VSaIZk3
MuvWmAy40OuvDcXp1QCi42QSYozuNHLezA7lP+fnECWuFl/6uFlkyQ09gjiV0Rfe
17PSYgyif5I7QtEH3Gbn7GzmI+JihgbaAhLeEf32ukAV9vxdK3pvqPdUiR8nT86t
8CwqcqjYaaQXTgl7gBRLkZunDwAqsC1ymnzhN6Qab30boskRUu6uqJPwu0zi6pZt
5dJBS9Cn+wp6jmTZkAEsrg==
`protect END_PROTECTED
