`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ABQhFA/lHDqJDMdMEd2FBpabfuNxgIcc70x6/uOE576xSV3P+91M+k6WnLjYdGiU
DcjcyYROjiwGtFwx2/1Le0bb01EBwQ5QmFoewK6QmifFyEus5InP8td4+pgA4G9n
8o0B1Oeq48u0W5WIBhKE+Un2W2quyqjNZXCn9JxCtL1g5CewFxeDNaNsT7kaFmKw
ZgXMXvG8/As5F9dGuXawHPl/2JizjDGmDChIASAIRnPt8GelUzO97GsvrU3cLgS9
vAguMLWtrpUY3bcL6NNlr1QJVmoBa/f5fPwXxy4r8Ge0kjCAUZcgJJpijUD/Axne
0qyo+2KLk2vJ0ZrAZsb7x8WBA+ouYGIhtID2eBwYUbtCF7M/XnzE5YSC34dgwzRU
dhxbnbt3ne+qZ/E9O/FS6Lj0zFNkjvdrzgXbgMoYvgknJTViG34sMJkSbTTXMrds
i5QrKj2KTVr9wLQM9/Q8hq2irW9P+OQ7rrG+pAl1lt4/pa0+WDUWT1Ep7hiAGnvO
QsbU/4A5+MYVi3E98wuu+GhFoVoHojf3d0tNKMKWg5z1nVwf6ltP+Ha/H7bhPdTK
Zyw42qoTrk3K7v/l2NAYULVBa2CDjBYA1GMektmU6LBRI6Z2nOA1waYoqToHzlG7
7fdbtvnRl70W3uMI6NHUiT1I2WxZPM1WeJfyCetSB7ccZlwPvREDV6ICSOmfEljo
pHV7kqFEBOJYlmor3S1JKy19QyZv+yq20wYLbw2CBYbFh9tmPKpg+omycnPITbBe
D9cii/NjGFJpEQc75WXQOSekYjiUL4Mmf39mj3+7JN5pT9U+dq/sULxkem9Z3LyQ
C8F6lYNralZ0Dengh0HwPkHk1IqKMLFe9u6hGkwMzT0/lQXCBBOsLcG1ET2UgWTg
C9mJCFTzwLvyfN8Dcdt0sCwn4z4fm2QTJ3jyvdZinTo256PyE8aST8nvupmh/MyL
Z/q950YGZdYfCzLirVvigQ==
`protect END_PROTECTED
