`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+VnsspWuv7//CnINc48PLvh77opejy1lPBj6WLW8le8Y9PKI+jhY6na6vKhmY4od
7ava3oIQlntVcGuRcmhpes+iP0SV/xeRm07lfVr4z+jjY0uvfECFXM1cHEEG+xOX
S0v/ENmSyY3betXRcndgAo2eayPHnvWWQzX9J2GSTib8YSviwWdnkKvRfTl/zyMG
vqVCSHbeOUyVlfKkooE/5IIgv92U52vm/lDWgMNwhZ4PkpVDY0tCRBAY27KSzjCr
hBoiY3TqVL+RdJdVSdRyWIyIGTnOUnOuiEaJR2ZVZORNnmN0z0BtqrZ1Zg8NE1mG
OzKjO9uJkNhPH5XAvnY8uKlGgsiKOQr6q+Pm8vao0MBRWe5pju6aJrbnbWvaJC3e
ysRCHCx6PlsKupaAesKgEw==
`protect END_PROTECTED
