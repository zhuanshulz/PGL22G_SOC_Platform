`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AS+CSmygfc5WKupo0PXGScS3jinIOJnEZVXHLVvSiZtfK6o4e8Z2PcKto2RCeXgD
EVT1+pAwH9x2JTdCljcmTYE/3BGBhjoZZOXXaJqrsDb0OErOyCRxCbQytMNxoDfy
URvRvOmFfBBH8xCOFd6kg07XO54/NDpRFRKfHDZJyYKQtOebB42VTT5uDgK7EP9v
kWoSHs8jbckyDIDbUj5TmxtYyH1y9F0VoUiz1PSLYu5+hhmTX/tg6TJp9C8y3N3L
CHbQOZz4XBQGJnRgqitAACSiPITAeiOrF9X3LfHUVzXbg7xXV/9gTODhqlPmj2Wl
N8eBJ2m4rzNLcnWnkx5vinArzqh4U4M0wsJq6Ve8N0/071zqg7IkMBoDVneyXriT
XMU2Vi6tBgRfZPQ2XDiNCzMUQr8TaVZrReiq15wWfu8b/2SqMnj4sHVUVDsuRsNO
JvuLtW0+iuQlnmmb4PAbtmNm8yCy7UoInAy/1s7SskHIoRR8g6a+MviCuT8D1Iza
swZCcCpJ+9Qw3tB48U7CpDc4/3y77O+zojJxmWG20OiBSM1DGl6kGCxio4305Mbk
8yJoOwLnIdPH4cFhAQp+Q1TSuxVWwzVuNUYJGFlNNwtkwHT4GZICOG5v7+AYO49b
FgMwtNLgME/e1opY0ySty8MoDGQqyAGKLUiJiNbxHhNip1hSvehPlFAKGDgaJiuh
zeX0Mfc6/4Z84VuSFhCTHyVP+C/uer6f4oG1xMz9dJ06hvyTDlz0o7xLkDaAEhC6
FFrpDoIhaFDStbjvCJEm/Ov30/uuMnCQo+n4KyLTkAB7RFRyir2JTIt0gG70EKvY
jV0nA9kU4g1y3ydtYEg1hJfhvDIQgFz/16GwmczQBfXQ0o+R8RSgk1BREgnTYlth
/No9pcLO5yIKxLbiE1PJ4H/CVZ8eWdsp3YXUXVb5hn99c7+XRqNhh6bUA4rwReM5
sXJiMhUUC/Mat/tjuZ1m20hihoFuInZAkq4LfEcZ2nh2tuYDY9lrTi7OKIVFpMsA
L11g4xWTwpXOIeZj4LTGYuNWwPINxpjDBMkd+w7aJhMatzLhmucHD7yjaClpO9Zd
UFUKrNPJaoQLUKvflE+ClGCqGtesocVxuXvEQJc62P0Arv09CAsQ+2uh76ok3sd8
lvHS+4nu2x3CajkQ350CujSxU8sA6i6b8jZm44ZAdmV7xgXNZrykLEqlg0yHCTV+
3SRVXdt5Th9WNU+iQXwodefaguzYsSEoRnUee0bIhDEg3+c+06VkXmZKI1QNEWmD
MAQ3hzF5pc05JeVHXySeAMmfJYCAzZ/6kUgymlFJFbI/tICpythR1nGF28bu99FV
QFwSvcRrZ3JrA82oXcQrXYo9la5uJFUWgWoyNfzU/1qWs+UT1O8lMQQf6OkX/XKY
jn7zaU0Xugrf9s+PeD1cq/4P2kmzMvWxx7oFF0uiwb9wl3zPbBksdZ9y/Zhxgsg7
/lLRTOtH1bY+FGHEBvLs53QJmjVgrU7g1I8ZSoKeJdIrDUu39mcpBM+ZvCsZzmlb
XRl/sR2zD+a/9hxd979Xex8QquHsLoFaE8JNgrAIkNZ6RodMg32Sy94y/G/SLXsm
W00wPwu243Vpuv4VFqi32Nj8HaVihJS7q+A2xTKNi1joMv/q22asnhUAPqT/WfuC
vGSIC3TyUZIsBcEi/hfnZWvjzvlc77NLqoQQTaNsWABh+y9eRl7j/lmenxkar+8r
SHAYx1b+Hey+3EE0Tkt5WA+Z+4eGPgV1IhLZjL5NE5BU+TddbQeu3Z1e0mmE+4lY
vfyGs6JT26lTxkTmWVbLy3snYxqlyUPPzhVfrum1EY5du1+1ZZwl4Kt/Nc1YGIgd
2LxT8SYU/lVjI9jV6YrevWAhIogCqRiKd2rKLXGKA45VKpkhEPrL8v5Jox+Qf/h+
Rer5Y2eUtZhgq+cXmyuWOhwGEzOBN2j+HM/eX2xVPWnnDJbj2OcpHcLxXuaFx57G
w7nRPxD22N3TrMUDbx9nuOhIqTe2TJM6kpHAPeZdz6m0pKsQmXV7y34/wUYjt7Nw
+MzSQphk3naJUMaWYyGAVZU8JhBuGtMibAMw5VAAlc+slNluEzK0qUpdwF/1QQQC
EjYSWjvSbkKYoVwI1HhCK1cRyZ8NkmLm5fMU/4jVwJ1sJ90ECI0KXeJIFEA+OH4r
iEFgWC9/pNBhtjvS9+FEyhzFyc0O55mvstdSRZjlFJ2ymGypxj0ITWwKM8YOdpMB
WoI4cog/4jXrwSGn1Plzgw6mWKVLNasI+PUSjOwr1LOudMGHXLaKZfiVLo667ZtL
gLsO6Z1qpNlm1HNLG4IKURRvJwNL8x5Cigovk8d73OVWwRjwBizNarea941md0M9
YAjxTp/7IX5vxHVGkjTJnJaZptiFy5slLXq1JXLyoxcnVAjgT2KjZ9FzdCHyXyv8
DjJD0fFSbuTUlHZZX0l5hr0Nr1Tx2bOH/WcVs8QBZu9GW3NeJWTvMHYKcfdybUMQ
miPPBdyH8E9uYVMEoAWajp4UWmRAW5TnxELQ9ELUWPhwMyItVxMBJwQ481L9cq+r
yYwst11tRLfdczE+UWTj8bgp27X/VOynDhlxma/M9YRedbVEpb1s8sj9YVNZqf1Q
2I3pBXV4YFdthn2pKNU1vA7iX7wrbARG1M8Bbg4+H52YbloFMy/OFr6LE/cK7/gX
1Qt8HY08FdOS1ARmJD8SK0TaZUsVXe7exxCW+ATUmA5OsUzGLavuhGME7m/KBsPr
/v/TIokbKU9bVDLLgU5RyY+nfVJ0OzFzSAT8ccW5QixU+U9kwkJgEDYGlgjiR91Y
OXDrkd+/GK0kosxzLeBbgAgLxvrbUKUnx4ELeHoex1ovHl6vFwqYRNWR4LJIBQk1
F96DhAXdhuVniZF9XDgxMKeQjkfoqFGmFe+ZaJ4XPL5xuuKvB//ACTOqNV8AWhia
TOJymWUpnPaUzo3R+Y5fjXQibpSjFaUqOjYCzzx7wEaOdGLpmcIx0yVsI/JmsiM9
JvhwQEoS1HrZYlNUFpRonUubRnFtwVTQ3k7NmrRcgvcsj2S1FAlvPRAT9wmNWbwM
sCprIr0QgFYscXg3taUXeDjjGgl9l+ts2CTdJsQxeTv55BpGWVgA1wcus0Fyp/MN
myHNQBc1LbboOUgi9+IkdUvVGyPx4uR/rm/INRPnUksvNzQ/ZO+650Ld4wjMiZ2q
TZwFC02BXpLGnGtTNGz9FgVuGRGyToTM+/QKW2uLUh29YVDmxp0Ed2To/6HvVbKP
udA4NgpCjbuPTuZAGgi+xXk+PERBr9jVYxF1fMDMcCtEy1TBGWKaBs8neIxPprEG
Xy4b4Ru7mZo7s2reWcGQ9ex6tac96eyvWFz9UUl4tWBYVQvJg6oyKvT6fd/b4tUu
t2p9ixBj5e141Z7GgaIEaaEHQFdx035sD2WfWU9aFKPRi2PhyfPc81g+5bkrjs7K
2DY/+TeMtS9JUzo4YqDavJSgfFwf8w/BooRLax61Pcdja+2f7nN96bnHeuMtMAk+
SBemQ7qK67HB2jrVW37THG1mSvyYWkphY5NZ5QqAWylzBL+KBSiCh9KiweRJTSQg
qQI6gdRu8/4Gt5oSptLaLkurUb+FQ4TUg/o65+oFolWnp18atHo9K1qDDwUEn8i6
xV3/5MgHBRQ6lVDok2SYkslOuj00418nEEifc/tZHmcOjw3ARs+puLk2KzuNaQAq
moiofWhxbbCsC9XtBOAln9a4ckpgiiw9Tnq/h+euDPAb+WYFD5yJMwRRg6iJsr8l
O9voFWy7kpAobj5Rk0K52tDKF3A97B80mgR20Fb24jjaKU9vFjmX9ImKlyboDX1k
9/cnsNLh7IVS9VZKZWA/+v6QbZ2SeodJzWhzsF8vLNA6YmxwcIdbE/rRwB6/cbFi
2Kb+FNH/E8G9qiOb6ZFhwbSQNW9u/fapi1IfAc7KBdlCCZFN5dZ6dtWplEA+Z3E7
iYj/hxfBdr3SU6FKmjhMcjSblU7A+FtBeWdHa9q8GkLm61celG6xPaVPhiH21pSC
viZ8Y04kz63NWFzprRJ1ankcqIO68m9tH/MuHbwkMTuedlawxyv1ssg9tqbxpoNM
3TPHGmX4YRZuMWl9Or8yl5xk6lYKZoEYnfuLHHi2koNPwjdsrfMmo3WHZcOtV7IE
naI5CLea+MO0PIyWS3hEJ5nr5Xft/Hv7pJAM/cK8rc1SksA6N8Nbp1C7WSL+vz++
h6OHx7EKRJuZqt5jZh2kaiABPhX0kZbbh0YxzjikRjvOW7Jux34f/BMKFWuCQLNR
XGssNDlUJxI19yvD9FtKtltCakextzjgf13CXFviY15OG2r88UhG6WulN6GVnH6Y
h+qwgnmSsMDB3IHOferPDkI5O5ABmjb1l0kDiK8poh5XUGQAKup/E1Xn+xVd5Cny
Yo77yIL72hwozNQ6zbg38DSzcLDbEM52R684695AMGF63abZDRJg3z1Lmi583s1z
xtf5cFo7RZ/6z/E72+kLvsHQQxliL3R54MO3vYStp6HkenJTPwBpwaumdrJXNfds
TBvaiI04a22ZzcDcqLehTE7sDzJPyhpwklfMeQYPv9R8VxqN5879hGZQjGa7I/3j
cjHB1Bw5uysVulempyQW9A/vfDHi+7zmNqbBq+DC7Azq4RYAYHaxcVT7XVqOyYrJ
QP9LNHdkNFPao611ZtmJ2VzSg3j+Ccg8CVRh/o+/C8bBMLvPDj2H03tnSTV5M4n1
PkJJEwwBr1TZxfb9BtzgGTef1tWIvLf3+MS/Hw6UQb1diQ6iYXp9uOtAZze5l2cX
miAWHTGgRWXX8kAbyIrRwk0Pyv4o7lgkGjuEnEyf0bYC1Pgoiz9QXX70bgBV9yj+
nzFo+RAHAtSxBQNP1jJLyirGoWLYJTfqXC2YcXN5qsSjh2+O/mQQcBUQKo0rVZ8z
xriyRwQRcWRld+UV5VrFT3sP1SXcuuOKYVB8YALwsCLk+vBIDCUb73j/Ws+1Ub/3
pZyyZbjXAB3RakMWcEourQReGQxifMaOD/mnFmOLwrh9U2ZfT5x44Vxp2GU2vqsb
0nOUG8wJJLl5kO4SUbZmpE9JWkTCPkchTp1aKywbfWm5DIqCzVaBJu2g0PCg4amy
lOf81Uy2HrMeWXQ47+/1orIV+ifOsY1IiCO/czTlv2mkGWXKovKRObsnXndo+9i3
QWmCqWmNQDvWmIFKV4LTrFPW/8x3CZKNWjAFCv5h6qDtMoVMHJJEkBQ18+N6SFA5
ktlgcN4gj/vuA1yrLRAkOsHcv+jMltsyqZYRHdvcMEvKV1FHniDxiYXpDDw23Boh
/41STUbdIKXlwxcrQlCJx+p8gZ8LlMCMnGd+BLcqzcGC7YB7X++7/awBeLSOXTSc
o+2Fq7yz3Tgvv+6PgYkgc1EwubdCLzvHPY0qeZtcZG9NcV1vAEoh9fmnOT1xPVPU
MHWD2CusDPuTgtGlai/5A84C5y5vjncLx/i041XGZEiAOzC6vE+YFhUK+cdhbRVp
w6fcdQjn/er4HgfLqXFFOz3sIr2EgSqnWOzRQ2zuQs63v8erqPRZguPoqcSVJaF6
gsOhV9urafg9d/Hy6iRss1Xw0Bhq8pnN0DmdUr0BM5L1lnS+qgyIZaptJlw0HL19
gJwB+ucywKE+2u6oJYhYXVQQ5ifL7yt7nrBg3BfLwKHsrqAcmPQAqu7k89UTlipb
PzfxhIGAI9VPSlQUOIPqRBJsYBWe8DtM3599/1GMS8ykplfbzqhrwnqnZCDL+6A+
L88jeL6SO5KGwRGv7b6bBZ6lBwlmRfmjdHRfycD8xoc3O651eZhTP9Tg0VyuzRJi
xTb3UD3tfD3TbMbpvtDb5q5yvWt+RWtmFgCsgphdZvGHhCNtpUC2JxL07Rcai30p
+nOBkzwphf2McFwtTXyzWWvV+kvdf95sHnFvKj9iN670kt7c/cr9dbMt72b//+Uu
h4T46wzrXlQbF3LUAhFK5ds9CAHdZdpAYgDFb92Mdpmd8y5rhCnH3ZFsj5vQyA9F
JkPuJ1skRoyq6y1JlXZxfRKNJGLtRWopKUGK/4vPS4KuwDJGPWVkPZBOEbrzkHfF
Jb0LkYyIDB9LcWzCgKn+h1HJHDxU9MO+sjJeR775t4zql3eBR7jozpNwo7uIBx/i
zOzlcJuJu8kA3DDgaFIFdspmx1NjmIBIvK45OedQBjlB5WjGdTJufGPJK7DyZvKG
yJZLy60jD89hvWCySY9auZWvWBEekpF4cTZk5Wlv8VWKgMAQsGnOWU9Sldd9N633
XiEgH2Gd36iiTC3me/SYI+fpZcVqrXHTwT0a+0QOFnzyt247t76rSH2M7IMFEcQi
3CniwmsvfyP/RHVkfCIXa1+EvdRewxcIEzOZ69jZ85ehOWWKXDtDUAJ9JJpgLnin
Mb+dpD1bb09siZvlOjZmQzQwLvnQsrN8WsxoAaVu6Jah5HOEB85zLMYOxa95hBv2
TksFMdmqAvm551IelcFRSf8fzsStBySGRuMUbMQfmG/1M299MZ6V+aeZLDxOK5sU
JniQKpucrkQqAFP2Ug6KuWHmsnsZNTJLOO3e8TexPnf0E4ejQ2hVZxYqE2TGCIBS
B/wj1zaWqTs1npXjW1i72EQtCAzeULstCCr6rHRX3tLfghWc+1pAIaOGGizGOsQq
5cxkVoCfa4JmXWxgRQN2NnXfMHOl6ql4y5Hpnm+6+AjxjXug76KFIHulZWFDIEQW
gz0J6HebnN8fA1bL02xjGm+cxINqp36tmVQin9LZPb8pWNadassLWcGOPhT7zvNc
9OrPATr1dg4ndORLREU1ag==
`protect END_PROTECTED
