`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EnrfilrLyzZPQIKNTM3XS9zUlGrhjQ2CY1v1WU8yuehRfAL16oflw28YA+/HnOG3
qs3pG3fbEwiNXAukt8zz3r1xCMwUTgegiir7//g8rKhc8bprYK7Sac83ju8CjiPR
juHmOtT16XrBBVN7Dl/xGGwEMAhiLfMEDoopcw69/D/m4a7sgo11JxKJ/cuLlA0I
aQ9NjsrOhviVI5kwZ/DYWSXRuwo2LLNtVpe3QFg6C56XM5X7WFL8RJdgRpeNu6On
WaLn12wE/dzBmiqaX4OyGaVfVvWVY+oH1Ce9IHbeJmJo3qi5UP03uINBRg5WYoiY
fnMpKjLGDa0JmSZUBWew6de77MmG/KG1nK/8AgkE/6D4A5NwXG9mDCIk0dM3D9v2
dj6Sz0nz9ulNUNfrx5bdFGLTP1rb9ckGCyFeilGocfSDtOXqiPP1+A7wdiyS5ocF
K8YXFFyMsSfi3bOnzgY8QuHktfB27MycGsP8R+ZOenybzkwHQty5zOoqZlFPK/Xd
evE5BrOiKHUhE3Md6AnkFERsfYG5tGWvLNeQLSyqn48Py4UPX8ZCJltRM++/a9lF
`protect END_PROTECTED
