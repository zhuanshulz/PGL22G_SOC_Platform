`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gHrpEbWMuVZ8/4dgDgZZ6BeUvHxY8PtaHpdxL21rtmrGIMCJaJFTqhaTIoOIw2nK
eY71RpieKFsy5YoacXUxBR1eUvzd+GDjYABEBzuhgBHooqoHRB01mM0qEiFYXdz6
kMEl9s+lq5oFPDud9k5rj0hI59bnQMTC20iD5w3KlvxUQk9kkIjukFhjWGDTc/yH
gtrMvHbvyIVQKQ2oZtrQK75PFPPuSXasTHr8YCB4K+sUYmmHRCTSCo+ou/c4xj93
tb7iZSKTlOP+mSuoLQcx8x8lq/2PogvyEpzhnjA434ney4UP4daSldn2To7Nds79
7ivQtdI8eYzwqSKEQlGb2EZHEHzk9GvPXpmm5ysJsCjzS3nq/BZEuln9Mg3uH7ha
X9r8w6Zv1VQh9ttwBQMDzyqIOWnd/mxBFcocYMRpuEkvKs8tsjuyIjTjrK1pwIgr
7rspq6swidUv79E58dpqA8kKLTEdiFnNFYE1/5hPu0qvmJR9/8of67RvJ0L1DLEG
/LbLZBAifYC2IZfxI96mBJiU29YFlw9lctch1nh7HaTAn2LygGRpP481KF7TbdlO
psEa/TYyMW4GF7xslNoOzr7xesptidrX9cTCRjE+FbONy7eH3MkQxtfytLul6/iZ
`protect END_PROTECTED
