`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b2Qr06SS+pNt5lJ3GiEgxQqVUrHa4B/DuvegvGIiEQx51rCsFa55l8HKbpC6ZjuL
A2B2D1rqO+oJ+iUu9IP66i3pXaz90Ckb5euhMQ11bdxHNgvSlVnWVQN57ZwSdEA4
2zwSsxqHyU7mX2l7osf4PRNAR5AibTHDx0TIEKmHvlRxQoqOAwk9U3hqxjwM5R25
Ff+PBjQl/y+GGFvIodxHnt0HaE/wNfZnwqaMWyQSEKFHogje/uTnFKreGoX/EYUx
vJvf2q7g634zcPTYgNalxIm+p13N8o+soEsg/byL6Wnm1b73y5tSc6j/fFxsl70u
SXYwlT7OeJB5vLrLkUVeRNLViBsDXA1o/fCugEf4/uAtNglSoQtQbIZQ2HXvfyRT
`protect END_PROTECTED
