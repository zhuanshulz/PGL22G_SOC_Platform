`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aj27W+uGTDahVBxRCicciOHIAro7r/IzfnbXsio5TC1l/BooYzQNN+aV7CwgwQx8
bBJzJSe96B5NzBjYugfTV0tVXo75wwvH6i5x5UmKCb+IoTt1zmk/+iarf1DKby+Q
HHaN4VXhM3A2Za+Axau+kV+jwGQoEkWy5iuxQjvCU0WkuDPutvE28qK8YcsE8qLB
FBK6O6Ph0AyNPc5XaIibHwFjJ1mxfc1Dp4R3y6/+5YUDLfCNgFDWgY4fd9tFPGTd
KkMrbNqkKzCUYc1CU0wa6iRiW8SgO/Gk+YpewWj3WOifh4fgJ+Azy+LO/c/7+y0m
ptSKW/dgelGMoHoAwxbUuxw06ujLU6nVd/Sj5hsCUM7PFhubyOJrkjSR5N4hSPLL
54aACgBRBD5R5/Y1uEYhnyxBM//G4faZsEK8TX3KVrQykLSnboI2IyXErjoO27jJ
qTYnDx5xtOnI4sNb5BYB4NoiOtMwmSiJ1b6jw8J+mrbUBQWyMRsvS0oP3errJIBg
+q65L9UhgeyLagvLUNTV/jrMoK7+dktlXHMnWwVgU3esaXcccLXMQPdrH9YI31OZ
YDaDSynqgRcP74XK1OOWn0N9KQZUnwGtMheYaFg1yjRmyWinHpmkF9lTYrxeUXfp
913sur8MjR0tUxTjA9SDu/eDfpXCmZKu4X1UHhIyKKeY5B87/fcrzL4rGxnWI0l4
bUiu2NS85tzX0DNsxyjC7k2ihNfDVSWC44kPqGz2k8yZ2Cq4DDmNRLJ1N82JPoB/
baldWDTbAZvUfLfEYpwi3/OXmEv0tmHlqntsk1mLHjdLtP8VU2BD2XJRqTYXP/8f
v3nfv7IQ7oHVulC9EqGNdodhFT+zs7vAUmrobewF7zyvgsJbQpMzmztr+4Zm5lpZ
wwvnPoWyB1SUdkjsZDZxSziab9IgBaTe2q19+M1ZQRHv9RwKXTbuphLEVTBBeenr
T4Oq8DWEHAuJ3EOeJzO7rKtwr+v3R7q9AkGSDxt9WOn2BKfX0kSEpAcuaZyKRb4S
R2hlSuPEuxzP6xn4vPhr1Q4gDYIstIIT2uqKw/JLuueoENfbz07rwJIUU7ybfnFj
HsEqWQ+px8LH5FHo+zDNkGUvZ0wO9IJzpnUwvK5v5yXdikWFHAq8yfOGUnEhWBix
YCMLSsegPIS7hskArMGaHxm8j004pYbPaeXQbvbelbDRnDfuthkdeMkIxvs3TwJq
V6IE3f213hV+TyhLVP9ULWzsXtttywkwvsILKtuefezG0+m4DS6U2L7YyGDniXfP
QTb+4rbBk9IrOv9CjhYrwNwx/hcp1n90FrFgvbWlMcIaZk3DlyosER1jOmRhkyk4
OvSS8YaZgGAOY5iA+UKemw4YaCDDxthwYDIPhJv+SrDOJTyEAUPygWeGlwaGVSyP
Vg1GcderujtXhUjJfH+8zfhdTfNaqeG9f4NKcOzDDmtFMWfRnCteNbDycvorJy/X
DosP4MNurYsSNoq1+19q6F2Xj9268FSS83SJcaRfamml5RFPtOaapJ+OhOVWxEcA
6qh5gC2YcBTXugvNnlz02+uBzztdmFCyXiUq1eXCJOU=
`protect END_PROTECTED
