`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GCq4sk2AkLPMI2jmgcped4ccZX9K2XSJZtnEr/8mXy2ABZ080U4NtTCxCOKUCob5
or0QjJ+BvVZUMq59kN3BZSWU6AMeniBqujxs8UbSDM7mQs0Rl+9UIzyoywQACBhU
B+4n9V+1JabE3FJmZbzu4NEF/GffhyA14vR8QsVld8Sqx5aqEVD9Zswi6RuIg2fp
xFeNbbOGOaGvIpkB9zPCn284MC9VyqW24VQIHORJa9ayK707rlOYt1H9DM+CRDiw
H1OaUtKeH4mtKM50iyuHMAzZF9IsYUZSmZNP29/7BpjUWrvI/MEj1SWyTXjKWB6V
GAukWFzxM6D6yRUm+5nLIENJoy8ryWjslWTfJFqtsTsRQzOURPORmpzVUudaw0bm
ISL2hRWaaepDuJ3OcltzKPskreD0n976NJrny3TYbSrKEpHkbTXdMc+4lxEb9B4E
YSo8JMhESjFfPclyEC/PiW/k+cNz3z0j2a12t1BkmjdLBV9j6vbLeVHsJSmQZbMv
7t3zm1dCcu/k0jOGV1fq2A7wS5nIGESOVeWL7RjksVwpk4C0p6Ebi1nNVSytldIR
v7V9zFtgoaAbA6GGahmFCLUaP1Ga+fKUmzm23T7eGlwZi4sRJ1LMcwHytQncqxRV
RFO577IA/JwSwZ/bfsPfO9TmEUO+tQn369fVvCsI+MByD70C8NPYT7lSSPQmYR7l
l7pyuiSRROw4l+FM83RH97xJKbhR2ugvjGHazfsd78WkSjSEwNOG9LZYaBMwpcPS
3bxZjpgaa9bvWIZeEu5/YP6Au5qD/kWha0jz7qi3yl3wAAJdZzbA9krwkPrdq0jT
SU/yVavo60fJ6NC5/CQX10ZV6O0leFKEPC95+lYKH9a9IRk3PWF6vACfql9xuugM
Rb6zf44053pfZT2iyzC4sdWs1VZ4lRbfMmiBHQyu99JOLxuj7Vs3r4QT2LdlY396
LmMl/9APgJtDnvc+GQKcly/XUxaXifnANYQ7gZTdr5PVJpTzwlu2m/gnB9Laz7T+
ECeF6VToCIktJcQo1JrCcQksTTuXLoVuUtGZPlceSj/L6u4RX+lV7DJpXagGhLqK
jc0qydXsvzoVBdNJSVxM9QugTYsXGbfigHjJOyiBvuspLXshH9sjC9XKSSwnimYY
vgod14EWCJhv2L5oQTQdTwWsB/fCxkEOcb+D2AUaOSct0u82zrIvaS8TrO5vzYSL
gpzNicMx21Ys0bMdd+N5rqa+uZiRPXbpGmjOzX0m3+uhsP4006pmimAF580OSUTc
cDUF4qe1K+ks9UssIJeCuqhS45excyVJxHnOOYsrdt/OckNih4ckbmv3GaW2I3ON
e+82NbLA2c+kU25WaFx5BIP/2oXnaEbLHMmmKjZ76NdCV2lHvfGFhXPokWl8T/sx
wAxPEASVemk2NMh/kjzTzByhiuGV1pAGBIYRg0kcKutM9m6eF12Qw6rgEN3AD5lQ
6k2L1/m9/ajWEPlf9EJT3lM4tBQrACvd+7RBr1S7nHXOQGNdU6U8/M9302SEfYk9
XWx9wu20dk63MxJPFPGDpNAbfztNa+lIYoEUnRYBEVP0QpRUxmwiLMwKDGKTOaoq
kxcsqplc8X08ilZNpdsOawz3YyNZnRc9vh2yG5VU7N0oTSjxArSG6lBEw8kwP7Vy
kAtDgSaSgxMMjAwngD5fCuXShCP2PM68df9n8FJMh2LuJaygpe3XSkOInQKNi0+F
9Jc+qOwzOWBun1yH8Jl9rH7Vwe8bcQ3TGlkze9kExOI3gwx4wWSBowmlXe+aAtF6
5EO6jaM5JIvI8U2FM2h3SYzpXtxVqejpVQeloyHw9NaIBjNSwSF83WXLyHbWgQlf
fmYY/Z/mzONto7KwysbJADebtASH1LJrDee2OTEUsjAB873FO4tTwoppWLQBorpA
SWO2r8C47b6kMYdGUnJHtbPpma9oUXIxdaw+aGHEnTJiQK1OePDnltJQKTRTx1F7
5zEBCPNWCFwWVjVggkKbBaQf4khYzCePHHqrwre2iwX2ZGW4uKRZHVUBCrXGSsaD
R6FYWePiWFmgl658FCFgMVrxYJX+ZRUXltNq6VRgtsoW24DU70cfplwumBLsCRCo
Z9tEFsNsCjP0/M9yTR8+ihF1U1hrHr0EGzYfmkjXD8xteiOdK9RUeFJff7bRMQX9
vzNbseBqBBz0dUzPOPUEyWpNusRnw8gTmZocCLWw4i34F6NWIPgNqPFw1wv4PZIG
uH79fSx0qpeIDOPmWVt1NtUhkctbdRFMPi7hUN7R0pLTmbFZCHdJnrEExR5LYjSe
0l6TbTB6vKwhhvX/fieYaArt+VXSGt8wmz/eyA0qZHiLnSLrHMF4pgpyUzRI3Y0x
`protect END_PROTECTED
