`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hxo8FzzTscVKQlcD7dhfZFOeKwKMwp3ZxfSrFFB59ihQguTovGqzoGrwr+pzkjoz
MpoTVNB+fVAA+E2SAER4JJcp/Txb9iE/520bPppaNfQo8IsfqV86YUW9Z7ysTapl
/uxq6QlegIp0iOZoqxrKWvs5+AsoSNxtIyqe/NbJPUtmd0uF8e+Y2+2iZkVAaqh0
tCgLnDJ06z6qo1vFk3nwid0YSYM2Z0LJsfZV9FirQpqTQWWMvDE4Hjzpo7RcE6dx
KEOBeCYcMyLCL/BvjSJdpLY3pgjC00HiFlLG2UmrtjK8phgQMqmcfS3upYMLFPgq
pDz94YpR5q9p3QEScJfbpmvlYTzezv1rE16ezjauWNXxanp8L0k+IvUbhZQab+MA
F63MMGoUbJhMcKX58L/OsjyvI6q5HOOrnG99RqziXxNbJ3jwYhQtB/UcQqx4KHfR
T2RjKuFkXJkzb7cBH5YYbTEBCOX+YvgCCo93BfG7ECS4U36Jqm4zvRo3E5SqmKgN
06hP7htCkwHbyGR6GsjxhotVR/SVqMQpy44YrNpqdgwb4ggJj91IsB0UG4G9TtyU
z9JleCe5Ce47V/c3EcpZjQBIeUvxQLIaSJDWKvKIzimKxqI+xoYmc/I4VTw2LO8/
xaiKPg0JxizNxW8R+SIeLh9DpMxZCQnCQyqo5BtpZjChZO1bSMn8LlMLpyeVdixb
5LwFsWwwkDpyCewSkawWpWP22QfENln4bfnVV23+IQszdN+ubOL2Q/WrAD1bwYEo
HpifZaco10g8pxJy82LeBRpmAWFd/uKev2nFgDMkCeWscHHSXyZ9+LROBu3JdG1a
Qtytr5WCEgKnfpGJxYqfDOAcGr1w9mfHShXPRxasr0dx2tKdtgu4K6g4S4hsaBwN
C371tf7xz4+eOVq0C5l4uBZUdN99eiugewU8fFSx1kUhq0s2/mxf8WQq88adVypa
bw8JkzSywxsBCrni4c9aorZh8GPP0VTn8dYT9XZUrpJUThhBq5JuZsaSlUnUmUvU
SsmBdWH/wWJd0XcRzNZeKPrQ/5HZ5uZKmBeg6zOQo7VoozrDTXADgsyEa0kIyAUk
fsxeKRdd/g3RL1IEj/w42/3U3CE/qXeOd45XmVqSG1KB2A1k5Yxd+GMlpEB/I/Tk
1t6uU20D6hz438LrdwF8G4vRGKJC7oDwOjOKXcU40SQ/BsHUcUR/GFQ6Zn9783Ks
vWyXbD8Hjz+XPb4CHReRjAfrHI0kv7eKeCGnsmtmLMtZtUKrCqf9DyUYzVUHg+wY
VDff3imuCueu5EfsK2YVJAQHeyyFKQhHDs434Tjo8onFXw+qsl50CbaJCSD2u2Hp
TngfPZhAdtx4/+8iIuLapNGeL+rRlHUJGMAatxHpgsnqaTWvHf7nJticWJiV5sx/
s/T7qpRk6jiHtw3nCCjTpAwcTL92IsepdL22jQwWS6QKI6nXkoNZA4sh7wOHyySY
s5xKi8Dw/p1WXIuVyuRU89KPkj96hradyzB5UA0Jzw18SgXCy+BxCl63hI02BnxV
GAGzZeuFG9bYAn8bNy3cT3yg99Qy97pTzCzSWblfz9PEdaqn/TV5DAUZuK6ii++7
8+Lqlcu0hPBTeHPC1k5LKFKaZe1VPnOnp0o5/BIv3FkmtNkK/0rjG8d/EOhOuNmC
Jaf2nKac9yUWkKqWag7qdQ3swGbgE1GtXKET0qkC/smOu80Z9QrsbpXk26TIO9ZX
rJC3LZ5Fy1eXD7I5GP0l2w==
`protect END_PROTECTED
