`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ik9xMi9CohkTu11GRn1kvEDDx01GADmTtRiV6z37SK+jbgsturjHEGCdWFVzHTm8
vxVszx8ebgSUqXu3mX7qXhIZeE8WAGunZ7kc7FpZus0nu4HeBncNMM3VuGUtS9Mt
1GAz8sHHQJxUEMsJRrXm2nnYMk7gZoMHKQDzWfeDd8erK+3z8lWsFc0enLo2s77t
hIAH++ARJx/fMm3FH08rYe+cfwq+3wNtcJ20hQfHGCj8kJKyf9YycjGZKQlXfIiY
V/fYyoP7pmlDRfiZUcnqRyzt07qDMIqQ34o4lMq3Vy4t807xdRo1RaCW0wWp4D1s
9ItcPqSXhDMU++1GcUwL3anRDIdNtfbFPoULTyrHSRJsigbmlduwsG+s8C8lfBFF
xUCtm+wLb0vRZXi7q72qUHNkRMwJ5R2JT7FK0sGBI4+1s7oXqyeVXhUVWbWvLrOl
82WdXXuAk5Q0RbQmlkXFKURmntS8HQ7eUzCS3oa4cVtiLMl90VtwUXoIOPWYRblc
IS8DC6r/XY8O/90clvZ3BJoaWNdVnz85HccFdGiSLG7mPXhHXqWc2AhH3Qp+SuVg
DYQBcswLKOKxLj94ABHlY7nynwPOorcvWRVC6VxPNRr4rdTYZzEJAntMj/PWoaF0
xmnaqpDm+eFulUjXN6Cu2wT72aDnZ0DNGEU+2eN77ao88K9FVXcKwkkNvAWRTeRr
V47RbQUOaZTDBXOfro0CB/JEmiToI3KN1KCwXemUZvYkFWGYoURvEDSsMeTVJGrA
JAaP8tsLfn1478uzgt5iknv79KiBCp37hj7ET04JFYDOkBAMfGKYbvHhPcf3GnMJ
rSfuDQ46o2vpWLb6ammazGSTKf4PqL65oAvXOLYKrfABiJiGKGjE58eLrWsPxBNa
1MKI/YqBTKFCecCM3OAwQERLX0pG9UbPXWcjN9V4tR99XU1rLWGJJuhxvB2jjLBe
Nak6lk66AW3hJBX80oe3cMaSHPVmLDnMcxTygolC5rrM5tXiVPE4gddmgx9q8cU9
LrGayapSuWv49+9j6aADL2gIcwdnpVlgboLugrr4iK8X/vbIawvkJDhwDgsIcHxe
P1qBny+xBu7kSRDjox/kScV3esf/pUW9NkaC6xfYZ9EkBW023QucgmdoN4g16Lwp
7SAwRMHx6HG4neJUruMPTInYjFdytsP2jykj60FMXcp5mubYhsaKrWY6Dz8zbJ1p
qz+NW937v49xTRwky9zSGJCAzVbfU9dwFZ4EYdpiFZ/QG31dy7MOtbvZn/U3H4T/
0fMJ3q/YB+1IvfAuCeVtVFyq8wk/y1OPrYoCotDwmdpF13ZjMn+zXq5P15bcehLx
R4X/nIL1VXL4cb6To5558v+7S1naRpSWf6rqKwXagepl8hPkiWevsI3BztydKX9P
NM7NZqgptdXzuEy3+8CWP8BmyBt+Q5vtZT7vaT6bX7u2zrtNLbtECV762ZKAjM38
ZZskw6xkadnUe64GL+5b74Vj6RYcQv5oKoC9wAbMj1uZ5DkcdmARMxhLraSJ1zi/
eJnKQr8zVlO65My+KMz1nikzrxu0pblMHvRITD3vZ2FckKjkXEtx8YkH2WkgMsua
qeq38HbOuGbtv3iP3qhX6W4ucv/OVqLZKT074twRMm/PKKbSGvRzy8asvJIPeF5A
KCiJFU75ciWtisoEW/h1ExvqjyCdPNZ7EGjVcJ+MVtf47SVY9TSZlmxwmUPlXByT
OENqfJLB/rEGh3d8p9NS9a/hS/j4zE6Yn7UbpPz228XIOtto2Thehvt5enjwck8X
jiobd6Zg9EmZcksINp4kEAVrqZlxdKs5N55r15DzAS2Igy/vSBE7Pr/zXxZ3t9Pz
s4oBTRhfALNfzsaQXYDuZlCgubOmtcJkVxU3SYKUMiuizgL/dv/52j2GNO5stVc/
vwchiql4xBJCK1H71mwcAmcvgaGdCorqXXPZRsInIdL5gd7g+TeDIonGB++5apKn
GKy8BkveKPTwVTdNOdnshljf8Q6k3OBLvSXBnFOYS7kqENXoOpFrzSqhP0yRfE4Z
3JeUDNvBdqBP/QBwjcLO7Iv5te1+OxGhIZ6twjpmadOceV+uvz5ECv14iCEtHarW
jkGlds9S9Dx0xUYOVkuUqcLoBn8lj7ZE4klry/CutdpoBAIfce0kO0KNknkuXfaL
+0nFhUSzE5c5crxodlP7t5ok8WoIfzS/tcIgHh1s2pXSiPZRH3x+F7NNUEQmWpoj
k5u1vsuG+63S7mRq9ZdgFtOykaGPuIg0K5FIacsaplU02Bsi6qddI26DG7PiaUZW
wJqVHm3/mDWKEH3cOHk/thdIWTYvLdXQ6MP6p2UmGa8dtLYSYncRplOgjJG6llHv
BpkmnaUnCFSMTn0nuLW7X4esSRYUFPXlTznYD46M6iuNWP4xKTx7Mupx5ju9Lvjp
3q4mNUIYdptLPBLb7Oj5XxJSeoCQxCuPKs5/PHNjDi14BaSNIpbAN5nIJCTVwsIz
SS4bPX/9jLeLGEqmpv7y4iMousrrqvY6UpCLABbg0kIIaVBA6EkzLNBN8G5t2aaK
W3r4BRRbiYqmc2agiyRGHXbi+VOg/2hDI/G1g/FTRXvuUoCmvj9OlmZ3tvFJJxgs
g2uFTrjYw2fy0IXPXh7QgVVi0F7MGWnWYjO/2mroQikToqvrgK+CmyAn3e2yiUkR
ckJ4YM+krrlJpbRC4FS4xm2FiMRlGKlXMP8AmGAWnlPd70W4qVehCedOhy11BFFY
2BG60ae2hB3UK0z+hJseA7Pco5nL07EbrAYjvhbih/1DhqDCOnEg0mzFQd3lPudz
LPCajSJ/q4io4lL78pLmntb9NI68HtzQXB10N80Yet5GrMgAVRJ2ydGqjY5caONJ
G36AYdbqqzeJy+zfpZHAXARgSNWYefRJCZ2dmdL2+f4D4R/jcP2sI1n2D/fIGv1g
+lgHk1HgBV1w3oJRp7kakPGhmZgphtLxlZAQaxHxhInUNXiq6RbIRpEAHm1ytp+B
xobjF9bIRHvLUKEvazu1XMPMJY9EWvtkjSYATd1JwXczfR0t0QA7T1q6iuU5reLI
PtRDRx5DTV+9I7cuchbXD2bWv11jrbMtUf+IWHK6efffkbXGevdBtsxadfu73a6q
stGdtH0zgcy3/weTLF804jqhSREeQzbIHEtSR5TqrmJW9ae7R7dTRMHhxzBelY84
d34bNitlUEtKH+mUzMqhYxR7UJQzTl75F9OlXcGyOtmnRb92rd/Lwo/VE4iUqNoY
BFgnFN00Haip0UaOOG5EvvQIWLEGsxzGXb8ur/iaXO9KRHbjwPHr1iW/rYjc91zK
wPqcm6bFS8H+Zg1ozqaZ1+MzHB5NoF7AHwmFBClI6NGeqmRykAKQUJw9EPwuN0Wo
3ZWNotbRUKCzsizeGhl+DzQnSK9/azjwM5YECBRaIH0FCSvUAyYdAVx130VFTemW
EcYuPRIV8TnMy3m7QnY3sBgY2CDiTZiD874tfaW6JVourChat1RuKn9XKWjMduiG
TzmRdQqtG8b5d0bJkP99y9P4BZD5Huasv3IRb/fDGTm3A8DLDIy6OfxhmLYddbkg
mJXJJOrjEAT/wLiQn+wnmwGmZfZyZXY4Y+1IDfXEDqOT5ncjx+2+uInGtl9w41zB
bzRhOtETfZECkdf3AAwsE0+BV48iIVAr80Bpxjvd/lNUmBV/NS5H0fh9K8Jbb4Bt
zO41qIy2Ecga43WuEd1VhaDZDIDDEdIe7I0Ff31+JgUc11FSCMKfX9DSlCVvo4Re
ErRdwxESuNyrvYgnm2Y0axh0DByvH5hbEaLDNEdrRbocKILgP2nRadZSyFCTOCHx
qupt7uDPmfGHNlP3vLY4AwP00VbpPr18R9FDNZa2uISk4VaI0LnPSirQJPiWxVbc
WL26Rt67+6Pi7vety6XSU5sNVj6VMmknkF/c3u59REz44+52nmdf1YbH05125FsZ
kefTj8ONtpfBxndhn56acD9xqTE2A2pGCkP0ArYW6PKJd2n4kVQjruegFjUisrD+
y+qLf3Owu6FK06m4Zc7QLyCM8F94/I1IziEp45rVdpCA23lGApAHzf+SqNNok4wz
mzSWnPKkL1m9nM71I4qQYFZdvwp/LPCwMrGOHq2WtiVB0DtyKvblB5wM3070IyQM
uMJxjQRqPyVIWysMTtp92/sRQpPSQqDRDAJQuGwkj9h7kahRGt8E5eDxtdnt/k3V
/7uTkU+MB7wqKHZuaXxi/wPVylaEcvDPx+TRuLHDcLywAXCAUTtuEwGOjj9bYMzQ
/CCxDl/kl8JJYq0f+ridfjjcHqqPwFjG3t+Hb75bGDGAkbSTDPScnWubflyv4yC1
gUpeE95WloDTE2kB0DgZPR3+5HRNchOw/LK3q3No/9bbqT+jMlvYLi7USxjakAcg
UIgqtH5XCPQKzmdnQ5sjctkORVmwzY3PTJofAytnQyd87www5dXK8r/OYcM2TdH9
g9eAMtrXo4bZVXeThWDxZOjk7sS0fY5+aeGboch0PF3nX5BlofgXTIAn4K1Le357
AJuwJl19ROsMiPsCxmn/nas2TcYG+d9Z2xpCW4xL6Jlj6Qx+czHZjQ1UQvrJdgbO
c/wjS+jXkds25LeBt1IF1lsEW4yvZP/++5M6Q5b498SEVFxB3Bc8DX7EZ7fYq+y4
v4kLCFUUi4YUub3XNxhkN4Z3s16ytlVVWrZthKb/+A5Nwih/mjXB6JMuGtWHqymT
r1a4OirbFZaBvbYcFt2fzuVlWac8NYiktdg0YNf7+lKBsWuSX+Pt8VzpB+tWZPqV
0EwdGwqWwvqOiK7maxeJMCN7uUQOzk2JaWIs0E5xq460jWpVjZfOFrHjLWw/0lZS
cFdImzA2/k89X6iKuQNbmBBasxTfReVgF2lVzLCHWj2QvUeLSkSVwOqVLQESx8gm
RdyvdIqDibSZnI0FtTlLn33MzZbox+OKaJcVi4VmLTgDSmFkKgjoTKDs+5+UvL1U
M49Q+b8znsBF6SCPg2dPt0pp2zHzF9DCKmVgB/Rg++5o1SQP0nNNjLwv3JdKZfMs
mm7WLBhmfD1ZVlil8Vx6h9QuGw+/G0o52I2RCnMGl6F4wSrJmrZgjppi1BI4gytV
SnpQgK0d8jLwiNHKmZmw00Jrt6qKM80OUnS2af68Rji/vp91Dp1+EJkvJRk6KVON
Ob16djB1IbpWW9MwDU9NdRCxnbjUoifxNw7HxQQX3ar3oXurDBzRvLUBVxrQfPxN
8SzWD8up7Tkg3Kjsv9nI+Nr+ETQk2Ek6gbL7kU9WZBd+nUVIxdDzbzMh0Q3WXzpG
JPAgFmGYunNBKj+puoguiIJzpZFSCRbF+EvsNHQ1wUwW3V43X+COtDgF4j7HEYSs
8665Ip0ys37bh7Z3ZRvza/s8B/e7skLLkPOfwFDnYiG2AXNfyANCgzQe4gKBa3Qu
1lpW8aU+V4D8tHz8bDvcQz4LyPCj0z0a18q0oZgMFDc=
`protect END_PROTECTED
