`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YBPy2ZMgGh3A/tpFYHe1QALGXMQioCVfw1lsoZCUGSw4ecOQyxQrMs5W3BAlJcFP
WcQpKdr/Pm3HnsV3Bg7lA/z0BNTWLdeaVWAqCUvwWRUS71KRkCgVRCLsGCVNJyyR
LRljDZIyJc8LESIdxwNQOidhnldsmWT3diFOd7uD/is6YjomwD8IyiOSgPbX4RrL
GSck3dTkiuXk+Qzhn9R4P1DbW0aIt5/qTCJKDtd9KmovPSe23UaiAJhSD2xlJKvK
nt/SbSW5mX6B0wt+rH2uoE6MfJ9LqUCALp4C48mS4e0zjwIb0gPZMXkLbNNTsK75
/ZV4jgdTyGdSEMEyYYSL13fTCoq/HHj+L01SuyeXuWWb4m65+XLPG4oSnxY58bMk
h1HnFycNQvzYV0zw0NZkcDVOQNdlDkflmnmpSxypl3lvPmQk//VvgVVT4biqFT/G
3C/ZDj+6HKaHznf9JcvioDPP0nTn04wt1gwI5ETslrXg0NXqqG1DhHvpFnRKABZp
UTa/TjPk4DrARM/OgI0t44XKyMyd7c8cRbGfCp7o6BPw7fBsKfKp8FQicG2OMlyd
cm8LZT/DYFXGK/oc9TYdJMg64nK70GTIibxPyemrOrcmdUhEsLjBgQPyYVFxBeIU
BVGZVTqZwB4awPoXjrrONgA8iG10pMecinCCy/IlrzjWsAdAb5uJgeSNF9fjWY03
cmEnmi62lKaztutRL0M9xjscyhFA9ILYkjyewyfVUU5V6rA+8F64yAeL0kmRYDSn
uXmILrbfQDqX7I5x6OCZ8/1aura4yD76oFGD5DBtURw5S0NyQaDUyMnHZuUMrAWS
Q98OFkz838PfrnEmwYBBiO6/YnJ/SIfBkuaHd8R+s8TbGHOjJx2xPFT0ohzB2O3Q
aMoBSU1RjJBLmdmt7Jvpji6pJeqxUqJCrRTbYqL7LhI=
`protect END_PROTECTED
