`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fMUYyoC5hOFbbTIG+q74eoUk2BqX+3Va4+mvLBdM59sMp6/WyfdJzk73EZthM4kT
9SePI7UCpDkGww1of9503Ymx6vbSjbgfxUl0x89mG2OhU3qfmXMK5s7wYdW0Es/d
Xo1trObiEUCXVtCpn7zUu5yLWjBd4ixnhxpbP2jBr/TtgHofV0tFI368Bfv269wX
6yNt/UiqpeYZiDOrXeFfrul66GDdL6SLHvI3rU0hloLqU0Jl6aCUphONsoXRNwVk
1vaIzPskNNEWDd1+DMkjr4w54RLn8+/EtRJu+SjeUoFYqql0Il4gmJ/YZKiaCwz8
+KJe4EjJ4ymGZNs2BDp74gN/ZmZcEXZhM2yP0vv8wu3xuntDf2vAqWXabZ0sj0yY
sigH8V1WG3fVZxobtLXjiI8SBBkmPpkeQE9lxOyvjuv1uNdyLvWmD2KNdbSBMX5d
jWrX9PNSFL0Ey2HZO6m4R4CdXGU4pImSvOp1KsML/7B3Nu0wSrBzFsFUHQapTmqY
MkFms1sKJd87tQ7LFnk3mIM0pRw2Xp8c11B8KeWFkzdWH9NL379hdrCrFpWht3yb
BuA+6ikWDpWvS8KhUKosq1PSHHdvYk5HrJwjTVEZGyCXeEXB+yIS2MQ803UYrIFT
xaABzcy02CN69HESE3DoY/RFPJ0wTNSzv+KpTVW72Cn3S/mK5fxfZOi1UikIkZEB
uXJYOuKGEB1DjuaxNlcs3zL1Xu5S6WTbJBfXIb3llSYahuTvSkDLrCVZE2gYAUwQ
uwnu/bRr1pmOG+qYxinQ8+RcpjPXCQUOEdhDUfug/SiL3jhdoeWaljYNU/om7k7V
PObrjSo0B8RUazvvTSl+sanpeHwcp9WCIElX+mPTbC4hJw/Aldbr5A1OwAkqMFgf
YRpFOxBquorH72Ux6mG2ocmMuNjXGjmFofVkzLuizPvgh3CvnUAAcNQpLfn6soAe
pPYGSmHADEBZ/DpJxrdY3neOhnv9D+vJYlvmaqZMXMOwDPf88+KaQwwzbeRY2TUY
s2A+LwrFhNAT+GURUsReLg2rpdNuR6JhoKC7pf21Viv7Wfh5RsZ5MHi6e8SPb2uM
wvkalvN51QbwOupZ+FcpvRmOomQ4kWJnSfi/5xhnpMsJYJhwSm3cg81i9Catg0b9
TTsbNdrlsxLhZfZqPQUW7LcXzyH0AKLit2zMdy8UiAYBS+0pfWMf9qr8+oMErQDF
WlzrUdyzLOBYUVp1d7VwWkMEGJBuhntT/ijKO4c8YqsYEcgApqeHVMv7ZigdjaSP
qaVRTBH271W0fdH0LLPkwWtpTTGmwBaYZPFp9ngwW5IhlPSPtOkzLl67jeu+2Fj+
ZKlyJNlLmR1JZKuxbk6KCGGq7+i4OKCh0rwECQtr767cMxqGhqX3X9wpMzMISukL
hA4WX16y7SMNXFbE0WyF02ZBxisYbzQ4lhRhj7U2Pj8nIaAPqViYhQk+MBu3OVQr
gCO4grteLzKmRJce2D3k2obb5k+jCAPCypE2WalLrZS/uzfYZgPmExA4LZd/odr4
zB00QSgH32dw7o0ZSdxtVwlJBq7Ward4bCG2wI3HlO8UN4CT4qj6/nxxpgLAFnQo
4HjjxTfYOClMGYuJdUSE8RV9t+GZSUMffrvMAtbLMWyz0OoMeuT7QwkkaCRljUf9
6behDA7Zr0cJihLuZnjgoi41J0Our1zE125r4aqwkRP3GgxFdxeqCFtO7XyvIkWx
L/+gpPXuj6hPK0UW9UWJFfK11VeXPaZpuJBkGze4YqOdlj/YsfdMB0fvJ/2tstRg
x/eKUrFUGZPMlCkSCrBoZxoVcoB4XLR+OWGOb2ioGH4rxiCSL65Gex8bv1IOS6C4
RB2CeK680Z8sE4aQMmXDa98PbMGJu9Q4YpHZSPvQbVRW6spJb8DakqJ9Vbb3SscY
078cgC9ts0cu/HrEdtfhLUWH6QNrAPo0GzWabvsIa1KCBKEluUQYH1yyXFN6UN0q
M/5ftZWc9mH7mT6ZiOjofH3vxdWli2b+KiDZuUZPUsnYAR2NnJ7jTi7pDg1rdAtw
dzek6cO/UnHzq+3Es51JZ/iKVkuYWG8MeHeSdB5dcaDEmg1Kw13N5hZqYKUoeu+L
MGmHVTmM7j86NQAUQJj9402c7Q036NwyG0XHXjyUuMBjgl+uo94BVD2q59THTYkS
ti2hBmKjKo3NeMvxv4gU9IGpZnYpbkZCCQESiI+O+UsXcZI9bJ6nDBPo0W1OPFuf
65BG7u42lE1l/cYzur6Fc9acxXhtBbb0RQrFBk3lgvNudeljXIj4PJbYiUr0xhey
ElOmsLp4dNRw03vj+/n+3Jd8NgYj72ilQ0oKVhJwiRnZ8CFiQ+C3q4GW71LYp4yV
rMrjklXzDYASShzMo5fNe5ih8VW9X6hHN/1/v5fo38cufg+NQQXNZ4pOPLOFi+yC
ATkyhX96gRw45RtcqI73Iu9YbAXtRkY5FvLqn0kcaRM/p5Rzx5yP94JPDjVEoGNn
RRu7veMSM6Y5IY76c/WLpPaPO0w98sxpgh5rUgzORT1hCVEKwIkG+4RVtYLrOjCb
ss/DHg/fHnby8sijAqDRWNq/gM9vtcA55Bb28XA5bY3Es2akqBWRoD52O3Jxniha
z0Vyx4RTiZJe6obv3jvdMpUssbrcsATeBRHCwy3Oh4ATrrCGj4K4Wy64AlOUlTTZ
nf4cQSzMcUt24vPi307oJrwXQOO1G6Su69FsT+gr+DPV9kPGL8wwZgzK03CxMdmp
2wqYHn6tfSE+2d971fvZ7HeATwW6bAsUV+nPcou2UU5RLSXsZRyfDWorQAwtd1s7
60rO6unzIgtU7EypAK+wDRaSmG7n9OVDnYHyUDSmC/fZ0/Yq50F5O4ahtFc1prna
Yeq6jOpdHybj/lC5dqnaiU6q9m6lIJqLZF6qOy1wDpKfgd+S029EdDQbbIZMq2Jj
TakxIq9tVyq/+NtVojTSkj3uxuqSP8WMIEgdFupZfdKm203hovNvkzk7X1EMF6Qp
0OEDx8ZQXabi917O8ceODJTTpB+LWwH64w/DiZhA7dk+dYyxLAii1hdn49ATBX5i
+sL7Ljo72M6zGpeegTAawYK4Rc1Hrk+15Opbn+ogin3EHwEwPzxjOMP8PqNftsRf
5nUnWpC8jcU/DmRgmS/LkEohC14K5k2FUqD0TYz6xW4avZ4ZfNTOTsFNHIZHFlcA
la/LQ5V2fbHpW6W/WG9ZnySJyyOio9+r9/04QKp1wYh2uyA+Jyb23JiL+aTpunpe
DbuDdYlNbVbRg/diQ2PQz/N3mSo73wb9kzlwu31xl94ZhFycq+GK9zwCB5Ypm4S5
eoSQ96rl48zWf6FMNepaHrSVOgtn8uJgCGfx8K5RUyLZQloq9r4HNnM7449veH6X
+ZVpGpxfSrTQgKAhSr9+FlMnlb883vh9H6u9UnqeKMh28qMMGVbS2QPrQD1rURHh
luAENYDXhZIxAQwFwRtpnE1fxWGvu9E4rPnXG2JNrdgpuOAkGfNGtOoLAK8GxZ8P
JqFyHQW9vkeB+yrL4C5WnHohHjmuE4PLnZcxWJFvzzJ/J/84jZt9MRyvlNermfa9
SZXvyKxi52THW4rh5TZBVukrQ0W5JwRwiTIyCww3Robif/gv98WaZ6WDPTPYaQXO
ozIjHX1nWxEf0tZPr03957AjPsv1KEIXc2syWGKd5ggDqlUJDOt3RG1nm3XY3KIw
VfBYOoowWqwHcjyNM4boxEvnWOoW4nykEOr6NO6wD7i/AhlDSSGenPWvI2ORUtii
fsZeJwZXCRaFI39XL2pGfMMGroTj5aagHFsYwNHfOScGLF9PT6aS5IHa6uvuyFOC
Y1HFoDblzWhxL3EHmFhoxIiSFXop6HfpukMoXWeFV54eM6Aue7qCULHtMO+45Kg7
oumXZw+9ELmLL2PA+5jy10+/DNA7HVVoype7rzRW/eHt7NhYrcYmYwrxFY248q6D
4C18mjuVk7krHSWp8h4UJA2Scj0MqYUQ29K2ILR92zzKzwlIQFAtOE5zsH74CRGp
ldcI4ugsHbWdgevADJJlBIQ4I0yghTjeOKt9J2qfUvGMm1XExVrp1NUV77kVLoqk
C2yVf6zYoib+tWBYuWvKArLqTojzx2yOUrerkLQ7cmKxK/YGz1EREBZI+iydOFKF
gIV/GywkY1/4Y3gwZQLx7yZ9jdwjXRJo95Azm8tsy43NuORgNU6zNnq/pVT3sFfR
HPTwbBBlZZY2vOYlH0Xmg67qHAvkgcAb11K2Vth0yUTx6Keeq1RHTbbuUQMPvfAu
hr+nCU+vG6roxpRXTeGkktzCMLaU8Dl851x/znU0SsXVqVj8lHCUOh+nAv+tCIem
vdPLJuGINF7bskDDMx4FdpEytd6BzzWDn+9/Oc8OgB2xTlzpS9iozJF/Zlv730SL
HYCI2FQR/ttVMw2XodxrbVkHwPIkNs6q3bbIV2OiSQGNwDol9jlaR08Bx1IGzvTN
XbazLzI//bjRJ+u7nj85Y8lCezoeUvXE2SLcGYh7w9Tsq4f4On3eQv3usw9FXGkY
RhRkd8y/xIoBmjGmyaDzimRG17L5Z9D6dO5h3f2jAu67W9SMfI3J2aQfYyxFsOFh
yA5zPHUys93M/o+Hdx3cVx7DNt9fPTdh1eqqaMmkWZOayjO4J6nrhlCysoxsvrzd
OQYCNqcS1AGVu+NSnOh1jpvNuNuEW0+csqLXG6DAoY5qIpvECN9lSCG0xlWRJKnO
VvZMZO2wr6FNJb0UDxKcBIviS+hrbFBw9vhs4/EeT8uDMCfyRhFDkC9Q71mCKgjC
4OZwEb8gnJVXFIcmUKjAlnevoheKW7esQh/Giu/K49R5kRNjrtG+PwRgizV7CcaF
ZOZ3B1sCwz+4eYjAH2TJkHCDoPvLFT2wyFK+ilWy9TYrFS437fbHNaYb5FZpRz5n
MN26EaonIKes+hZslSTaMyz2xl525h/BAlISQ4f5p2zRseVMEJSM1bSGatxpRJak
Xd0+gl9yw8nimquzJefqbiPbyX5dQGB7It3NI20N7/GLGeuiHPaqn4z2zBJ1Qc8H
TMK4vTk8tnQswupuxYpcHCElLRaz7ivflXLLzi7bQWl48UoJP5tICVzF5z9ICvJ6
9LWNwrQl+81KAYXiuLCYJxpwMSXMbqhyJhi5P5bhXRSUvLaCNAWlCNz3xyu77Md/
C78k7dsulkgxsm9TfLbIY1ve9aBtnqcwLH5h9Oqr6FKBC2iueUXhTVxEnJpBdPac
mtrtwJoqWfbam9tdnIWpU/J4XGo5OAr0X5gzN9AHyTwaHQS1KRgtCh9/LY4YHI5G
qBX4KPgdw5H1LYIixYAY6rqV9cqQnQoK2Fgmy1wJ3+XCYYtL6lpi7accIrkOJU2j
j2YWQkXHCSEwYNXNDV89hrgg6TCmtPwPlrqfzAZDuh+1WOLuMdr4UMP6qVCWI1Ia
3keAUUh6l1TqyuI22G+xWkd4XR53rH2uc8E4sUR5rseF+yPVubh3mHjIodQ9ucO1
BC90bPoHCaK0bV1Te6fx2Vxg+HSjvwUrlIQ1vxSWMS4eOTmydC7aLPHG/pzkHdLq
JVzA725S2YGkLKOB4LcPhKmqoIiQn5/+70tSBEYOeRaKi23kdnsjrvv4W3dTE5JM
fCRthlc7hlJZJXnwNfKDKVTJTi7T7NbMNDBnSXTvdNuQhCWCVWtTrtHAloJJCXXu
VWv5P9RnDl1eM0Q3cGCZe5b10SU6JIhj5j/XyTs2G9FFB2Bkl6z9UrcsOXbbQd4g
QTdhRa6NjTsz2WRkw8C/OgE3VuWGbXuBvKYftMP835FhqtauLgDdaxxqIoLf3fyQ
1d8f0q5KI12Po8CpWsgG+xWmD4QtrmL5pZ/iwZCStCxx29rfIDCuMPre7MNAL00p
rG+n5npI8DKkNDmUfXrIDnjBbIPCeY+KbTYesUzlH1N0SoYYB2q3dGYDNvGA1nGo
98VCuu89IOTeZeXiZatIG6VPI7B2POCI1lSA3eXgyyK66OYnB5Ej/Qn7yXcELcwP
HdlEE7PF5jnzQVUUdJrGIGb1Xb6IZD3hBUt/TezRvJSLCmrpVz4yNbvFsAwHXQhA
HslKKWvJSxLDOnjTLXUjhfbgLALjajmbb6MV2dvGRB7+EYA/iyMBVa8w9dulbbXj
inYAKzEghi5r/krnD3G7wgBIrae2S9PVujwh52wK/yAki7Zc/pwgKuFScSeKN2Vh
gXlqXig7bHGmVCzD9L1d6rZuboNbXq77J38tQinrNfGQw0fldfrQoydddoyf65wH
qImGJ4OL6kkCsyZQZe71rSEpx53hPpd0bnF2EgMAWgXaOBw8f9uofmhkGI3IfCga
7sdSibh4jumglDVzrxMKM+4HR0lA9cLB4NjrFLHQBesRvFlUNGhMYT7TQpz+vcZ+
6vqcU5l/ivPJ2fVjU3F37iiHcWZOxKinzcqh9Fe2vOhHfO+A4ZB1NL2tIXs738eI
1uxtq1HmNGEhnHWASSmr+MqwNbYhz/PsJll5nn8s7fFjb3lbAOd9dNvcX11Y5Oc8
cfYTxlT6jXf75iQZqe2svJNf7bk98LQ/BQ5HIqP+b1Z0fE/NQjjMDG4p7hqWbrtW
aIaHtp/LUICqMc8UETSvBada9d0A6Nb2JA7WRxvjIpn1Eq05UAtZORWSlAtRuhjX
rQ/WpY5JaTtpNDvZ9Z/4qZoDuhemqtnncjchFyMvGrICEHCtYLmkmmvADznkNu8e
zRjRN3r0vDCQTVK0JcE9+onfUWatg9KPb4AWGIQ5IzfxUJ48bMKSpmqvMFNQyVcJ
P6UDKo/qOe8Zynq4KEhJ0uNHQpHCFrO2LhxKpyvh52hpDyoeqeXKeIgSVw3+kGjJ
VQp0qr9LPFGFo6tpQbjI7BHkoByMgrQ1iKk6ZvDQa3oGhDKOLvfLDhnrZNL2N5VQ
RYeKiFzzJ+rbyD3/ec9MnBrEqtr0IsnNeWuIRO2qOw6H2FibqAOYbT8oR++uiR9c
GWU6+o1Z+b5Tun9p6JwN0pkwrNvwUf9uxSxnsCb5plgJ6wx3CGyvX2ar2QgHSoQV
HmmuPgIbPwdjracmoHFq359GeB6Gk6jabXRkLr7qm7lSXPeG6H06CvuyMSq6uj0s
DXmZf0II7A6HKmQ6Dt6SWMUuX61uBP5/HjXAuvuMPTsrk+qY8HugqVGY3LolGovf
Vq6zIODEJ88peHZssFdlW+3o0PqmRhjewfbwzJty1rw5MQ2HYPuwBqGbgK5Yqy4O
omDPQTSjOoTPLyWrPRWh1wZj3a2rkeFnCCtKGs45WTU5BAp6PUbCUdACTy9XRUBt
Yxcacw+bIggfcddQExkThORHXKPTX3lwh3lVlomS30je29e1/68PluzMRassw68m
`protect END_PROTECTED
