`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jWVyfZ/ChLPtCiqyldwVVucmwFalYO0ezsCIKAbqmaKGnD2Pw12852QC/Ifb1BWb
BW0HuzbeaQBhctAp5RBPBneBQ5iAjySGeHdOalHxWGXR75NoY02XHSMdQ7993T1m
CvUfXhTpaDOWaFRyUytmwFGOg+RpE6roDO9/RBnYssXDDAAYYy/5DsvaR+HZYZaO
RnXEeB9XWGau19Em6PtOEMTROuA2LtCU6deMQHu4yo6jWHKKa4dzyoBjhgI9s2c7
XTRr8zrCs4ZAFip/RzxF3OsjHtmr/NFP/XaYXWi5MoawC30fjsDJWs82fvMCZwR9
VeHSCH5+BN/BdMV5ta2CykEEnFwNdcS0bgl2fXlbKMNpwjI1OvKmOElsLq4zf/9a
G85fmV3Vs8yqSvoUxYmJRJwWZagNZr5Oj9ODvmXMO57kp8tIz6N/CuJ9Hn9muyta
DAAA4EX2TQVIVRbKbcF6b5HrmarzVnVa6wzqhQ3Q1TqrihZPbbf3BvL6EdcTz+79
B4KJpN0BP2lx+qNGck2jWfdmu1GcQkWBL2lKKp0YQR/RlYwKZF033Ms03VUF+c4v
cWevCJNpjfxztPPw05itx+bu7CsI4Xt/+MfSsiVYqZEFYzrZkN2Jw/Qhpo2opeUT
foRzTbSo+qWRQDfSrE/q1Qc/zxtzTSov29/UZ8ZSOTbmKPZo3eQTiRLNJ8tDgkfY
NezSRIPTNUvrNfgLHPJd8Frt2TibhV/KrUsl1N5C6Jxhem7sPmLjh9wTFoTp5Ou/
veiIuqW9r3Xyh3jJXwVb2sCLdHmjZ1hms8UHNiZh+e6c7TUzZ8mgn0OBIlZpMT44
qK2kF4dIXLHa6B9VCJZQLIz/7/3i+b1a/Pcywpi6Kv9bQRG7YmSmz7GFGG5/xkC+
C2O8LRJeP0Ha/pxkIemIIAdtKHvD9cFgb+D5sk+IIpaiRjRqjdC9bjeXr1p23wtK
YI6lKq6PIj0dgMvj/J7Z6MBbi5nqSzDLsQvpGqo5lkAf/E0xQXHgtdLZeltfM5VX
GgcLVxbnCov4LLLXSxOuPSj6krAc8RMwWXxyFo3XO9hA3BaSZ9DpBRR/HydzXlrj
iGPzDyqf/yFO+0+Hw5vKkVxHiPtat/BIEM3Q1wIgVa2zDBbepkiwmaciOgvf7Nve
iFC+QEtVi9z1FBHAf2btR//gUdkIIqFkoV+nTU8DVnt7htn5XQfS8OiqTT4Y1eCX
uUDlZsCFB3k1yjBN/byoLqiJUN6LWQ4zP9Fa9ViY/+gLyre4TPB7IREsmjILB+pD
8U0E0iXVfyKU7ETaR0Mcuj0ZrvGHwJSFdBKPDV1Jbh5ifCnsbrAG+YBBRkh7prKJ
o6Y7IjRhG2+fo6uV5qyGqz8PuGAsIyHnw58ghsdiUXugpoRRZWyDeO6boaYAP8Pv
xCdDLEbIUCyCe9LZoDeIw6Bt194tzVKxRz2IiUWhNQKO+YX645kd+XVWi6I47OdK
MU5FcryWjxIFG67xRsm4hmNP0gZM/i9irA7aRkon7lUtoz0JYMHTCwwlkPAJ/FYQ
6Pw7vGK0LFq1i4E/7kkCebTabIskyeaftEtxOJNs0pCPumBfFHJgfLyOudP7mwM2
r6rCavNpGByPIGQa8oUzu2ykWu7Rb/XMAl0Q9NzUgHhUg8GcmWBz1V2jYx+ZBBq2
FF+0qSYCtUDRJsKyPdjxGCZC3nFeuM7vWfqNxm8NYuoGUdX0arVbQOad7eiA+Tay
Y3qCm96M4a9pZTxHzXgidVb21UrBALhE4BhundB6S0M3GyN8jVR4ZJqcCEu/uefQ
6VZUchw0r+xVipSW8NjP0f6hyMSe0M2xFw1itdzD9exXECDHxjIIh0uDQ2QniA81
mFd9ebE6EdCIlBShKlDEK5yxanetyIMgHYAUgr8rlCgdYlEGMEoaQuRF+IWGiyLD
Dw8/BfFTxt5YijwhfMrPhgvRndMdlUlAcWo+FtGQ6wK6PzebWEwjaDNr/UahTTdU
5nvhkGiD3szktVC4WB0GthQp0jLHo9Fo9WIdrPmFVIama8lP/m6Nf8ShkXDGsfkw
40fbc3J5qPRQ+Qjbju2PBN9cz8QfvKlVU2owLVLNUHP+fhEU0dVoxzjzC5i49ZXy
T9qL2gRBkRnlqpI4kqia2cD9/32rPVSKFHCzmVQKS9SClQbEdMRkdTPzRjog4TXI
5hdbtPGSJEJY+cS6XmzMKj98rJRVTiwDgAzPshjusQ3Nhb4VXOh5LnygBcI8Zv6s
0WcNYOgxmg9/imnO4a2y4MFfIe8uWj159ESJ5pTBBeS6zMQfQj4hqtBlli+vkJL9
MuOdciImbPdj1Ze6vfUO87nZu3o5oCqqLTQGfbls7F7O9wLNkQ0EsmzlmCs/SE2I
lNQokJA+p6RSDjP/c211rxETdPvgwEqseqvFdynQX1wnMLDiW5rAgFxgBfCkTPRX
rZq/E585n6QlzB4B5buuvLO1IRtFSnXNil0nmPz8VjqrkK0LAZWmCbd9CN7Y5OMW
wNuf3KBVlDt0QbV2V14bqgoCT98fxEFk55YQRq3gBXMnQUw13Xk/WQKvXPFShDUo
320KhQ35ZIH/XjMTIIEtqbm+lWY9DSn5WQhTxCs+zMDM0IHAbOD8gJ6ndYiwM1b+
P4RPDTCYD/y1r+BmsWaYuAh+fJfpPHvdM6TbwMCAOaorTvvI3/ot49yQpCjoe7HL
c1vbA9+aFb/4tqU7I+rIIqnjvnUF5SqLFakQ1+DrHAGE/iu21GWpyr2AhaDi7oEy
nhzDNCiI7rLZBoozjI9XeZ3yNy2d9lhuOpseGFB9j6zkeILiOUnp6DWuU+zY9D7P
MzPMczhTgawyJVImtoDY8ssglJxGn5d6eu4qfX2eYm/RMd8bJmo0BhqtV04yNsDj
KwLyRR7vvljvJt+hc3qTbWmfbwqdbVFKZqR/bfC9dnTkRaWMFk0f2QctWdDpDrdQ
yupt/kKaN87516li//QnCqQokB7p9Mmobiaq+COpLD7EYbCHjStZ1wZMIgbK4fCV
X4UYF3OVnJIuNITezBA3Bmz5OJXXKrp5qhr1hLFsgY9/eDVgCNncEEFquQSRR1j8
LqCVwkhpHcxN2zt+rv1JcxyO+cCr7w0zoZF/9NRJ0wYS9YPMFFZC9k3Shj0LEASb
jHdy2GH03QugBMgqB3UWs7el1qXAm0V35L3I6FaqWAVxmrXYvQQLafZH1eGBTqOg
kODp4u5gD97sx/uxQVRbFMcUhjel46ZyQbhVAjr2g5Jmse3knRExb1LYn3pvqsTC
qL3PFMabSH2sqs8Ai9grUspP8ODjLQ6n2aIJ1TX3ZbOIVq3FQJzBtXw1m2Tce/Oc
MTp+xAgXIoj26tPsIKtmGksXCB315CPntY1Sm6GU2y9GpcpDx4BvSlOAhmT5oW70
nBbsfXjdZRD6kxXeLjqk5BDDoGOv6W8ZutSfP+T9Z2AXqaAZS1LZKq24cxyj0JRD
9XKrl9Dn0t7E8AHgMMHmgTdxidf8stjd4FCHj+vaEU4AJyj2DUV4/qFAhGwS/aE4
v/emYD+aNBuAE+3xHMbxrkqhRXhhFtUFlkAIGOl2ZQD7gxDD6SJi4DpPrqD1pRz4
BleCgNJX7tpZE7I2wKZODg0C8x3kc+82x3gQdfyBkotxH5ImxpqjlT44GwyC2FAm
rIiZa7gca0qDTm3APjVM92Y/LSX47V3s+CtZ01EprCoVMVHZvBDla57sKSdrFK3d
XWroFC3QrqM5L6QmpkYViMzfG4KpSp9zVEtYfWoHl9RVYgzJU3TLYxGZL5n4ARl3
a9dOIl9E0gSKmTqk3Qt8vBJSdwzsZ2OyOc1K9DrGhUQlCmt16oPTXuJLgaK5Jhbn
9oWBGx3wECyghAH855MWRQyrHewM1cilUzoKAXxJqvu5AKmte7krNn8B9+8K7yK9
++zCf58r02mytqOO4tzY6jMoaFOZ7qAkAzQXQEY38TOZCOxv+NGHRUsC6uptHfud
ZPPaY2BbWZl+na+aYatTh2/QhJJ/hhnQrEgF7F3f7mTLWrxHxNqMBiSyZ71vGZW3
xrtylG2BmfDK969Lyrw7jykC6IYJ0Bgm49AL/eIlOmmpy7uZBy8cu9b149DTcxaF
wWsUWHCp1oYGtPTuyMOZAV4VTQGuCCI4umntFDDcBhAziX92Lbcp44nxIKeTPAwX
lwyC7GbZAbWcq5YjaYLCvvUoPph5jkr20t3I0f22fFiKBy8T7/cp7n3mFJEazhAS
rtz9nhTVOvl/t+2OhBsfD+weu7NEp6cdbwLDaEHUp/Q=
`protect END_PROTECTED
