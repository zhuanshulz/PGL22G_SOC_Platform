`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rE3hQCf1itjcYqO3lReg41vIXku0RN+9eyJV6FY3OYQ3ByxHydlOQV8QsyibERWB
yw3qMVUhYpnzzyau00in8WqORA59F4dkYJZV8ZVaZXUn6FVcXwIWpxkEbPDk46he
1pUa7OUJlCwx+9oJv7bhE3eGdCBOj6tmruLwsW2F6gG6v6zJJLdQI9rxEEnorBsQ
WE8s3NAUo6fjsZMN2cuoNuYyTH47bcTHKlLWFQH+XMwWlWtVwH3SNTNbRiEpdHn1
g/8ig7JqWZANDSw21spSARh32pvXEzwh8A1yVRQdheljKai28uujnMkBg+yVWSrH
gU2Cc2gr3NHdUwTKqgZhxHIGutNMfA/PT5sjqcum7X+C0BaGpzTGEtXWFFKEEC/i
rxw+llNkkhbwlb4pyIC5wvRjXxSoJmvJpoVOkBSRJdCfs/jw/B2eC/gKN8pqr2Ta
5WDa8N73TziIBH3QM6Q2omLTRe7+bLqSU3zW7OkkMG8b389/zIrNJC7CpswMNABl
jh3G+VJt75cKPuo2RNXFw6SxLCIrk7gLFgas9apFISnNT0PcnemujUI4tzObfZF5
6+ksYIndC2r1/aow2QlFVI9YtwipKYoPDWrAiVcjKFZt+UnZznjwg0w6kcS9RL8j
MKGDrgW819riRwp9TQkLrwZ2lRkSWJS24GfNCYpH36fcklKdjV3Np6Sp6CvF8oPU
T+/NN1m3hkJUcsD8hfg0eS0A6zPJeQKahHbbLqRm0LfB2KCyNOr2lruE7J+pKXCU
taHfMkRaYjEdtBzq466qrt7xhmyVA0xCpCFv8b2UhHJHQ3vpSzrVGx5SEM/zr4p+
p0D+C3Z0Z5xESXqSazy4fkWLkrXtsu7gCFgrvlA0P3Qx9tcvRmEqE6M8NgLbZQR9
JSCczp7QcT3BDm3SljlcpPOCEF7hhowh9x+MIO3LjTiRXemI6v/HT49LsoQj6vNJ
+e7PhBXOeJIkfoA0rhUgisrrreBSEl1YV9II4yJUbUI2dzTKuXGOCJTC8QPWPqz5
ASl1JGMEFYmZgYs4vpgmHs90X2twg9oeT5xtiuVeZ9cQAKw3TOb1bZkyvM8K7uAs
nraucVi67iEWF2zMaRFCVWf7cWFgcBwcNGZzyMVhvCXq6QUYELXSym12HwcTkGJQ
2pgfGHaXm9lN3F5FS6ZuVzqB09eZOxFY1YkhBfMPNdHfoL08K2UjnDHm7D9HsZAD
MbF9Ojctb+iH1snlYOPmjZ96OFTCEyUo/g/AbDERwak=
`protect END_PROTECTED
