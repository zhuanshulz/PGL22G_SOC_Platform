`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2EJkK2lKdREyngNqG16lWpei3mSI6Qr/9X6Ai7LiC3sX20lfhwsm3RYbF3KZwi96
2EZQQOOwaFeCLpHU1BBdCUdi6lcM+aKmcThzkptRiQezDQtpiCo45OX4F2fNoa/+
QQ/JXiGTR55klFwA3jhGp9iAXrZmtTaIwdYVbP3G3HNuZM1TF0bS00mFqkALN5aT
pyvDDTsQJnIyuNWuNHWhump6c/bPT36+E2lY/0Zi8RP2q5C1Za2EnXE5UMPQa9/r
xTz6pZi2qNj/iuiGOd16qM0Zo/3iC22LJf1e7UK+Z5VzzQYG926/I4AO4g10Nxzr
s8rdbV4j2hY/H6L+ZxLm0qm1Z5iDBagv6/FrP4DkAKvGsY7xo8UW0zkWaRgw60hO
6oOZNV94DU65dF/XVahz9wz26+XfwLFa/BgGGqiBa0ow10wRefcu9DJDKrOl9Hs8
BJ3wAz3L5b47tI+CJJhIF31k6KQ2NbsthoFmfoRvSIQ9RUzs8Dl7UoA3vGwIVHfg
BT+9vZAKMHxmWEMI0+NwcqIxcAQPBqRXlU7pw4UG9MNo0jRQGUzoyBDqs7mInrul
PrmU/yAeA5622XH9mcl1O0qqzAlEorX+V77VR0JPY6E4e1qzWe6FatnXACUSsikD
rktUe0Sh5fh6udwozLFo+7/zfFjep7FFvx3RPEkELWpoXr8tZRdIe+XHHUjrCqAd
WC2FUMBCHvnAOhxC4+NJUQG6/oUReDrJyEBla6T5vfQhnH87KrlVQBrU49lJBR8s
SYTuqh5avIXddt0uTdzp/p83YohjMFHK5UzU+xNG+S+Dhu5OsqW1Scg8Yr1i+igb
eu5c7UD7esPNWPKKZqE6blqrtuRLzS+GSLlntU7KWxLUGh4daNyySPTMOcsiSDop
xc88QS4CffkC1hjP33XL8Tzl7OpZuUAXEvef1l93ZX7m3a/SjZFeOkNDsZKJ8INW
U9y62CmQb3GlxCwLXaHNi/S2Pm/eJ1MfzbBg/MMqny88HOgAchI3jskL6Ski2t91
Vjkqc7pEDph9yW0ejDth31TbSv0UvTGMcXj4zjDnpna03cPeREBDzxyNgwQ7XJCG
IF7l4Q/zqtdMgurzsBGsGo2wp7LGGxJLs2eGTFsySRonbfkgSpQhd5Zt6gzg1K7Z
/FdaHo+m5rc2nc4hBwwFaElnIamokDnUPiA8XCgov65S2oZ7bG+qFwariP2wqUc7
wonN75nC9wgUd5hvvR5QD/1cfrXOiNr3Iwnw304MHHpd3K/jPI4k5d0Bk4dC4XwU
b8qQZ0BS4AXp8vBN2Z7NkRAOEuhi4PYiLCGkvoMP4to1MhrfqEnGfY2ISTUDXpez
e8e3pZbxqGvKnB9BtOql4izCIw9QFUC5vVl8YFuwJo3UJEf3nHkg/O9jXQZj3E2a
ajU6/Aw/7YGWGuUEBZA9cwm9V3yOZwKe1Eh8TNT6L84SVt4RnBhHzI0kjG0h+SSp
/zCUrJ30PM3P7cLy3oktwzDtUSREThVjMxyL3xr1z0ZZ4bUU+9/XH7+3gs3iSSAn
jHSHeH6uRY0LCKKQdviYI6A9PfV+jRbDJqOMgEKcaHuCVjDspZ25yTtwdrbkXqWH
mI3GtagpJBlViYnSBSL63jH0O1Nhwknm+9TEkLathG+1kTi6RaubLTc8f9rqLogV
Ppis7xR4Hr1ud39bdxxoUz5sRTqTPEZdhj3LggqnH/llu9Sz6CqM/xFHx9oFe4ZJ
yuASkQGbv6Bvflaq6F005nPytt4YF3oC5AfjwXEPaK288H6HD8qGy6FTY7ZKcuCt
FSDJ8EhUXA0jEX4tksjZoC5GEyIvGRx+dpjiUa4sIwsVOIpj0jkbzql0ObI3Oyh6
ze+F5WUnPSO3aLLDmZz0uVltGxDVgHao2ae2AQCpvi4fhJwZZyuLpB+H9ky9VOqD
5mjqFJjsWDmAsf9P/mZOQ0k0/R5fw3BWtOZSFgqQfsKJxeiumRaAOvxazyTFBy9/
nXgzrpFfM60JRcGO52Y2mN5pWSrOHpmTWY3sGijBo9UEwusRRXf8MnNC9SCd3SRk
pvnWEYYiLjzk/o6nWaNIjrkkoKxnhpGxPdtYYnF/ct14OYkNMW6u/GA6SHyqFPT6
mb3ZbRbpZKmiTxLr7zhStw6dOUgpTBSd/6dREgXh1NaGWehIi0c9gbROOhhRFPJQ
Ig86iuxA2thqjMdGxG+TkCMrH1xFJ5Ihqu68tQjq/6yEJQXJqrtfyk8YLhfhN9OZ
RRxpmjKx4Agqyx2OvQ8h7PD0d18ev1LCYR7b918awHLiSEIHHb1qUU9xgJUrlzlB
HKCNZQRnYyrU2B77yy6VsCQk/Vlri/J6JcFcR5NW4TSrJWfghjH+5K8Rc/c4kELj
nl4aG1bSCn0ojIyFgjBvYyodTub8z5++GBBuGkk0UXH3/UTMfChcNcF5C7tCsrKx
Yoo+qS6Z9Ki2TyEt+e1C823alKLzM57Ugvi5AFBYR5xr2dKaJfB509TbP3EFFYft
p3xr+Fb3O9/BkndarsX714mAbzJORY73Y4+2Fd6dsDrZQxEZYIPrtY3gpmTXhECE
dFRHWTiULIlrBAr/MjrKabKRWaeJL55zLh6KLkOFcMzBNCkSgOG6cH+8cxoHEUCz
kvX9BcnWLPId1xzL6NG1ygKMfTLc+iZgR/nfNdm6YcPciiIMOyY6UZm0LkJCcTS0
B2Gz7oenQJn3R7SvR2TBE8xXw4P41cV7tvHhdVUabJaut7+ydiU3HkllgcX+fbUF
+n7ZnGBnHSEqoNY7/sF/tSdKaDfbSmWPgu7ZmfXRfA1H/pllqHqqg3GCi6lw7SC5
D2sZpq0NcwFDPgJxo2/oUQ==
`protect END_PROTECTED
