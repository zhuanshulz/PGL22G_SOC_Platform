`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/efcwTn5l+cRTbD5fgfedKYIvYLfTpjU07CN832BrOwHRYTKSQSEvaZOSq6oVbfJ
NT67O0uygz/wwgVMUOncTwpQMU6TnKfOfbnf4cZ0ZzaH9VM2LyXUz9zAwgq1PLN8
WHb8MM9uX0QlLZMXYQwN7Tr3UZZ5VaUwaWtGJmdOr5MeWokXaSX8CY2tUehdVD8h
0SwrLzvMXCxtWegDZFxPV/GGUAMZbfuPlK+Zid+rSPlI58U7fuF+UR7VUbHMzA1x
GXVxYb/fcp/vN7BMj+l0gAb20AflX9kmkUsW98uxg2Z5hgGhD0Jidsnko8YepuqC
dDYO5BhAB0Ua4nfVquyf6TLSSRpkxlESBdD2JIBfOpSQIru0rKmCBcic7kvKiOxu
P5vd2h2DhwEE9AakFqiJzGf2tjh1h+pEwt1t7kFmB3/6b3Pt97XIZoAqhLbjTpOx
pzeivMS80CaOHQdyihcPtpJmm0GyZRYdGBjDR94acdn4D2/icCf8B7N+1f0te86T
z+qV3TfWTV8n5Mve+YXzKAlbX4PhNeru3AseljXzfLA48poi6dmXY/eYzuSXyctQ
+vgSaHlBsDnD/IfzM7D7bhk1dj2qbE58qYycJcS1f3J45Ep+XajcG+bu4ZyqDd2h
CwUO0fiLOQkvsSUXw8kJjwmM6OS7R50nYFwx7knROSvdlBQyCV3+39tLAFCKLh6+
kEllhjdLgo97GTJ8KmAc3H2ndo80aYECc5z8k07zvEUprsp7Ed6NpFzVuHN8la5U
OHPtuXT83LRqEK/dy7p1UXK91aCzeanhpa3V0gUHdxzP4WPXKXPqR2IZ4PClF9UT
ZOsy+OMN+K6USm5uCF2mHzAVgpdQ9iv04KUToo/rzG32BLGvcUQFtSikYr4CLoFl
P7FktASmeChhsG8jHAzOwa3VePOIKj8MTanjcRiVMwnHAkuO/HCM9GwLTb6FFHfc
yvTrJU5XhWOmbyCF+q2IgJCr4mtTEp+GNUuIKNwKnMc=
`protect END_PROTECTED
