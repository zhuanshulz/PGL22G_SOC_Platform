`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4r3/diiFfUZqo0OLQiyK9N8FuYR1vYSoZNPj4JMCbNSszocf0wXcYeM5q6Td4Rvf
MJeUmc+3HPrgyjNihYHzDfq0aB+fngD+lM2/LieKxaKqr2FtDsezq6vpQ1uso5y5
V2l02O+3v2ASYf7DicENBfoS2poDNrDH3CoiqoqBoKapJDEgBYCuy8ltuACYscA+
PI29RtGMwXC6IVqeiQvacQ4jntv9Z9OKDXXIjXH7jV40XdPTyDJE1xc8tWzVp335
Xb+ggtDAS64VRwQrqyMg6Gln45fBjrAuu6ePNGeACeFnaI3siQvZ5N3Mb0l2/8v8
TsSh4ex1C6goE8lnu4F0fBsL6f8FyOrSw25oPU7KWafLqyd8oXUv/NyBIfGHmiO0
OOK+AP2aItCU5lreq0pqC2KHPO2QvdkTlXQHeLN76KGEsMcFhdFEyyGLBnmieZsC
sGgvqsoIOwcMyTDZcNjG67Jnpq30wOl0rHJBjJ+WrRqMPJdhw1sFPPk8rMwPn4gp
4vMhyq5PiN4+NwRvJnvtkzbSyBhpNQhe3MShT2Gow6uzf1cDk7ej0/EQLBvlKxxF
O9yZswNKkoyZsGZ+1KkkvSmznrhieb4UQoxF4d+NKpRZkFeDzIT0zPH++k2gFY1h
rE18qGj1wSTlQjz3NM3c6fOleXkTxBvooh7pyt1BMrWi7Bn/ofp6mzt3lmeXZbVI
b2S/VpZr0UaijRaq5tI/kjcaUths+z/B0Z7KW9rwo78Ke7sdK/sv9TG4SZWfKBtP
GHkl13BjejqReCh29KHxSKVttrddzeTPZ5cUdqsJOEI6P91o59oJCd9H5eFaYH21
dj2teoXxs23CV9A+xh29bl2O0jHqMvF4fPw6LCPaFZt3GMcjLpL78fjkEp3G6FWU
Xa41/rk0S96nAwTeOohTObTxmdLPbwNosemNozHowl/OBkosGGWLzAPUh3oMJYf9
JJTYjQvNoEhZ1PfCAHJTUprhmPH2CQXSu5SoisGbzOy8qxVW8wXRs6PKZXUm5+5j
FXsIDUEE8s25qheDCzSRqe6aXOI6NSRXtjrUqFuOn7unQasj/QFj1c2az72S2DiM
HfgqFSEWpXzu3yp4bFXqibKn3F9DsYPd1hVZCwARDbl3jSZR2y8p2J2yGjpYHMQb
CKODsn2ZTh4Q2ZI7wzxjnqfuO4eiKB/8sTLE58stJ9bQZeivF62omcsqBofW4IBD
BADOcOLs1YB9EBVIw+jR2w8t2kiDTapbgD/q85JEsU8YonT2qKbcK4nev81AZ7Or
2Tcbgl9DF4kCIotTFl9Un2jISjbkrMNU9MAX0fRYFC0oxHyxnu4lEmx12wvrrLvW
FIdvMF9PtAxf0MmcutUUM/TGXOsrqCFMojjyY3NhcXEnUJbWiTabb7Af0LoNtB1E
WHZIymmMaMm6Cv5VBlrjELoTZIyWrMhNC3uqwFOIQ/eODXyWRJahwemVxSdNgwf8
lINnXto8+Fme8WU30SmeePzuXrp6HgtYDKd+qouUfjcjFVA/qnM7JZxFGXU0K7hM
eqtQ/jTbzos3dIcTuOwDikxb7GOmxvA+6lONdqQLo8FyMUtwIOVQX6XNk4ni0Wji
HLfSjpooOdS6Rq4UiYxbtUTvxuWhzd4jndWrGTBR7S9B+WXHC3k61mtrm714nqrR
0qRVQ8tAmR50sG9P6BRQ197CCzPv6+yPggYhOGHpC9D9TvZRjfHeIfaZZZskT/8k
JQmb/hb0N1O7dk34gsAWZfUcf1pRv7vlY6WkR4qkwyedPe4JW2FYU+0SaX8HaJyK
dtddmAeVQZibGMkNJ8ms7/eyMtJb4mecFrd1Rz4Ea7ck4DFKQznf49BaQ5jbhgjC
4nd9NeS0thjsdh0DXHeigVg3uuZbhTK/BJSypB+VQWt8rFJl+2Dyd64wzRRmLOyN
CXxPVPt6r8Oa+UeUAeOA7FBzBNQ0vw1QyvJ4JgPwc0tg5Yk7RlGTtQ7z0q/uv0ZF
Sudaxl6uqwWlBVOeMFsKA6N7y4t6inXWJHarOwls6pYjLwDBkncxGBg6FewE3uZv
3M9txQC42rADyQoCFkyY0M58ocD23LmC/C4Y/5oI5J4ykNPaGSrqLG9DATGHI3bf
+cLY+wb4g2deXxlymKGOCeEXgsyi9SnoM4Tog2rG77bD/YmGn8OyNxBbSdqEMXr5
X2fL5Cbd9lStrRoFdXGABlYkHV+TGJthEtPr+jh4iJ/0foMe5ETRw/k26qXfIOvn
bHjvkoMSjxUgh9XN7dkCQ1+NwpgjvVAhhlNNObpPk/5KYRWgtvJXPy2LCgbI2a96
GKjAbRvoVfMzgUGi3X2v7CTooz6Akid66zwPMid6TRP5NST5nor60UlcY5Cc5gsB
1sPCeT8rZLvPil0P917wbZ5Dk7o+Hh01ZdyLHffJu1gTO0LBaYJY+vPzcB2C2QOm
vngn9jn8XpVX6XamZBIX2OzsN2ltiS5fX3NnVQVgN+17VwRIS92Cvy+YhBjSOT0b
0rem2kXI9nh5dh0MLzkrP0MIpY6PEvqwvImMctqCx+w60RmvdOOhKZd/zeWU/rDR
0d/raOnSVrK6xAAsDelIbvGLwmPQZcRUpYFB60A+tMWdw2iFq1Q3UNssUKOAUpNX
zkSuDwrWWuleSeGRJWIEjEFQP8ibAzZCvs3/nfkI6lWvqCK9b51OISMKkeW6HgzE
7pB1TXUWmpFdPPiNejBT+l4UvbqyQM2sexr5PoYRWhFnyzpHDRQW1joeuufoZAd2
Q7NPKQ3KHF79RQ4kQBfQKJ1UTD1bv8Kvjxo0vEw7LH4yeX97JE2QMbimjv24z82Q
Bcyuj+VbymsiUdjG+TwXYzeTT8vm5C2AgXhwfb5n0TEEc6uAFmtQIg+ZrhnCI+sW
Sw5sDJwbJ/C8ES+07Xrxrir2bb3aukHwdsj/xS+e1Z9GcRetBhBW/NHonJwIoMSU
G3Ctfl6E0JcIWmeFD7zzKqEkEZmqF0ygMJDdukNpCrrwVLoVSuYzW/FtwdEF6dhL
Dq5MJ2cCIWkqNF21dsvWXeSer3sjw0FSz0qHg8Jsy8rgkTF5DeQwsaO07CVH5AjM
9itEtjEGblEWYFmubU5KAHfnHu1ALqFyttJTXsYO01uMSQUSexdvP6Em/WyO4zpl
m7DE7BLn2z7B1YQM6yd8ylDpRg/E1Crng8ooOG4VpscBhI6mbe99iIoPL9A2/fpP
Tbns2HFE+MFj24wTV8wSY8PdQ4EG16GhVwy8wtdfKxviWzGdxFGKWIAlP/2bgu/L
WnzMFUTtSkodiR33lyO5tpaQru8OaZYs7wB9vj8eBHF3mOPA5KrpNhTV5gzQjyzD
g8OaXhPlKeI69C/2FLGh9Za30cSpsKg60I+0FuwzH0yGuf05cNN0sVr/aH8CtKRD
uzucQAg9nF7hDE9Bom+o1oBMYRnHpi2blr949suC2lvtV6s4Ig68V57JYOADqQ9U
LqsImnHJEFV87ErrfBR9LT/HDVUU86k7TjoERbhJxp4bkZLjgmOA/XiuO9G/R5g3
dYTDyBuvdXk4kQDBs0+xt8zXMW57jI4sHeodhsqLar3gifFOBL1ObQ9G195au+4r
UY/zD4mRKN/g+4+KCSBeYkHfA6T1SAtwHDX3BCK5p25pqwEkIptQ53VF6S2naIi3
lstbEX2nbpUfnzLCqMdreymwyUSDOfuUGhFR0oUtdACPW2qkdbNKTbYoT2WHBkIA
ZCJO8tX8xyUJxgqjQkCg+bH2tVP2YDcp+eX/OrYlZN5cU+M6o+mmIfHvwHObgCov
36mbANPNz98IHsMNViUj5ub0A9iQKkKLPrYqpYrNATC9DrnqftsyIsbYjRgkmuJm
pqwyWZkZHn/Cap4eyQCS9bnx4WMBNbqwydnYRIvzXfX2K/jBaSu5AEtgAK+26B6T
24xI75HzA0+Ez0s96ZHs+/stVq1P91x3T3uIgWOU+XeYwS6+lHq8J1jjOTCIE+MJ
PJwtedqgMc7Czg210l8YQ3P+h+1Ku6GjV66Iq4iInutezk5OfsWcHDOKeCLoEeF/
q8cnTvOwHE5SqsbwsRAZwVLWlWixhDWnn3EoWl45IZNAih1nBGl4JOtVhREfOTZ8
qsjlOaPRkaEXroiWezEqD8m9S4Klh+qAIUekVCDtquByrrxTVivrw9Wrp7BGi1jV
dL+nMj+vHjpCh1nkCAd/FoKCzdX3H6X9Zo/eTQk7hKlRVNs3zVGGjuk1LM0QC0cv
ofm3kzu/39qtiL5O2LwpeeO4Lexgx0m7HSfAd2+F7MINc1iY7C9FBc9nBJ/JSo8m
GD70+V2a4s+HN+05Z/SA45a8TKMJL53kD/eZMEvb5CADw034Tef7iF9G4Dogjgky
WrNbcuoKUPb1UKBPVjpQ5bxa11ffQkpTE0als4aSJQcdEXld/DW/PInVTn27eZBJ
d9aX9XkRTVbBsF0U9uMuKGMrIGbe5ySdIYKYbQGI6mm9t7v8zzU6gN8cKGwqFFyx
pmJBmRyq6OCTriz8Bo7oHtj5UgYHcG/gZMRtIORqToj4h3dfRLpZ4eS3nhq5xNUg
kq8/yw4wYyM8etx5foxCmijEJuETsMaJ0tofNzaPXh8gjpII58znC0wlwIjlb7HP
pfZHwYDeUNoPJSUApaylsO4iZa2WNsUie0wXzjMNTqcR6I2lU3hpRWCIbiHnYsr4
ZksalKecLbR5FEsXxCtxAdspUz1n/C0C75lyrYs7GaZSPnxrtoI13J482C+Z1AUG
KVCjzxkCw1wiT0gLOduudFsfZoQtorM+QodlAZrvXAyqS2pUF9iIwvNgIdLCDTUJ
PMZkD67WOlPigSSFbRKzTJh6zw9YBaDMh0+YKQ5S5/QUt+hNBeaDWE5zO/zrPOex
V7bLLZ4slM16GZ812IM4Y9Jq215AHVwSF3YisYokOqF71BO902KeE3vmEeFZbD1x
rICFk9EOprl9ysrnebf4hfG0y4qMXZtt+JvWwgPaR3X853MvgjjTqpLJraUXF1Ea
dPhRS447ydJzJuZBN+u+bhud4edYOCPZdEH5x3Gu+J2YpGr+ODy/+FrbdfUS1+aR
GfCMaHMUomfmTL5HlxdWjOmqCE57nD3mNICixV9ACp9JanFhcFGbe4nK3IxpWsM3
RdJsfWQIWWWV+qvFzycpALsUCclYwMYb8a5Nmaio/xraHwneNwAkr9xPAUskSOjP
IBygAWiqHdPAy+UD3xNpYDUPjgkGo6usdH00fsqMu5yEuCLyqii4oQ/vpOdhiov8
eXRkAhGTbg9jNB5Ao4f2o/jbVvaYC2B+jqGOgjD8da5sExJLrUUaxXBUHQXS41ac
03iR1PqEvd/SHHWtDAuGSw8KLEeca/KveN6ZkJvHTepvkLv1DuJ3A0sMG23bG2dR
6zLwGzrmOv4rXNIdRA+r19gsbJV5DCR8KPR0GfMufTI/XMngZHVUFYhakL+A1TnG
cznwOD5k3ug6+SFVGANnl8X5Fms1kJ5WGB5JhNb4mOHLwQ9yTTTistWWKGJ6Pchk
NI0YkpyYcepxyKnx5EeCWCuXQhtDSegm1iO8d2QIXL1ih6B569eQIPMAyj9CmzQe
+OGpffDEmrvi8BNBZ1ayv4IHWhr3GlM8CWT0vK3VaOuCNpkdysbVcDpJ/be7KQ/+
U5XNyhqrmxbB00wpTv2ch4gnrrrrXL4EXi2R7N+mz29g/D1lYiRxNzxqcbZFEpZ0
U7243KuO0VqaU26wQWHz+NH0FSED/EahrfF/ka3BDb66VDRyYYOV8mmvU+dwMp65
4Zuj+q+Lg+uq+Nl1/hk7lUKG+O2TG1iuiCKAuIOs7ziGUR52A/vs8/TPJOpozTH1
gjklcl8ZZAF1T/WNI+0832JD1xk4u0eH99TrxgRKT4cnf7vXFcZBaXUCuyHLAZDJ
XC7L0ncPOT6vVcDftKQMJmIkb+vmAGv+ygOL6m85F5RgXMmUEEsiNbUPBgOewcOc
dT23i3OzmbIApDDU8M+DFx9gitX7EmfjJwROFJ1v+KcvJdSXvK5HFe+UKFnohQt5
vwb135v1E4uHP4L8JRdsXo1mV32jQ7DbMhgMpVAVhscIcaxhdin0He1q/eHVpCyX
XMUPfj+KWs5oUacqJpswI3ghsE8jssne2/1uQIcJlu0k60wt2wJ5S7CtSkS4Bv15
tBaGvgSmw4bpQcC7azrpXZb9Fc08DglO0jpagLx256282+M+1LF1VUHn/MqD3K4y
l+9BVg2A8TPMhM4CSnV1P+OGfoosQlnYBAZRyqVrH88Y6wNvOGVLmaoiFBNLzWQR
4208edxOrSHU40wkCdoSrxIBZaZtAjB8KE94+vSpmJLpn7z95APA+Y/uig8nut/y
pa159jqdHYbX/Wy1DGMYWyi/FAsZZ1Sr7/k2M4/iG8I+bg4VCXN4ow0v+gVDTBVh
tDyckB6m9X0Wz/+XGhTiR/t9bUabnOyjRDFsSxpjqClz+Y++iFjA6E+YngOXqV5p
862g2fi9rthxlFGxAacUqIcRcqb94P0NsJwzb4eNsJ1n5BdUt03BZSTdYuELvxA6
b4iQqTs9WOTJrpZoqp3EGUoESHS3IKpyzNHcGy3H7E7KiGHOBNASLaeW1lWTIXA0
W6B+qqZDpKgkYRemtP+qtIkyoPt7zU6XCHJ6EKYe0Tz2lcLJJ83qLSk8MuEgYRuN
/1bIt7bE2dnTe8YOU/37zJHM19jDlzh/mVF6DPfj8pajX+HoTeuh6fhZPyH0/eT/
RJydXqRePv5fG9a6wf7UoD+UcLBJw8rHg7S6YZmBIGpi6sOednbYSrkVi6wM7BGt
7G/3VoHjcBZoe3blM1hARxcbbMwNVRVWgTr7scz0KSpV9DBiD1FQDa0VCg4j8BF9
0QaZ8yylOGivmXadZYMfQFlVKIFFTS7WNo19YetWdiwocjoReYvxb0Fx6Avwn0xg
xuVzE9pWGqHV9Pcij9RLzMKHGDF6/YP83m/rtoYqOS1TvnhGb2mOZQQvDRGC4loy
hIbbeMl+SJ5IwEl1FEIqLtYxCzgx74M7qWu5Q99E/n23xQcBuuDYuYZmFt7ZvckG
FiURvRD+rJuIduoZcIko5KUgyD3R3HIUG+3Tc4vNelIxfj/avZ0GbjoxyKwNFWYq
LgNjtjAXleM5aGx5z+bghWo0CCn9bsWvt0KrWk3DV60hcIcP6qY7dF5iZ97G8+IZ
dt/GwZZoxA3CIrrICcCSeLvnUP9LoXpBEVACm1+gyo1O4leGLdyqJrZ6szt8/tUX
VPxe+NS76cMqf/+AhoPuCMkzbvNFJsvTfLTpBcIQRFYnOQZcwwQ+mh4QpEXcRKpx
T1iPnnlsKNqI9vWPKrloM6gCE5UuXaTgcYMTyI9RaGCAlRDWv1J98wHA1mNw978O
0lQC9xwdrjUNL9117Wb+HjhoQBRHbg8Vx6ZVoRcI10Rq1xSr9QEQ5f1r5syoBPjm
5YtPTVk8oAgMW2yPrCSsdGRvjCB/Cqz5HlvLqL6BmAzYuTbj894AVQYZtdAFW7hd
MpZscvXPlM7A802YC5xGBKq4FhL/S3bO7TB7Jvb/xLDfUwC3r4DXSZ9e08UNl1vW
yIymSyekiz5nDqUGSeBHVW5y48On6setn2q633Zo80d81iBqLXPP3oDf3Zl8PpB6
AnIyaTk+MeiNFbzfamNU2EVh0LzFPWMisyeYlNGOQxbueE4zVEdOBnjgB9hAEX7S
meJL8USQOdw1oenO4MZJIWFdclRKS27EW3smWoQwws9BGHeHsYC5pKdpHtn8JGCg
k5oIN7UpQqYFwt/7s7cwZDhcYLrcVDJnq6IIv33d2y/j9RbAl8zXVA1OG0tJ8C2r
JaUsu9bbFH9JFT+l5zamFgLDC6sCU9geprGEx3hDnzfadnglgTjJkx+wM/JBNBAK
og5iaIivCySlOmqMgnwzQA/6sS52+4JJSFnIZh12l2lnsuD1RS/oRBhqDzd9himT
CpqaCcB1KBP4Gbqd2VKYgdZ0SP5olHwg9+bAMqkUDjnS00e8BAhfdXqtFrdHcvVr
eyHtfnGBrYjDvo7VrSVnKqvz6FEY1nCUdsPejbRwb/JAAhIWAjNrZGzG98o4NrOy
RE12fmt3oSsnNoKMFZEA7m95or1kNHRufgY+xFt4J3anISetYxOiXyWZ6lMxsvyg
niGdmu6jxLci3mdsTLr37kCKUiVFly/OxeGVFXPS3+Q+DTqiW1XNag8cBXXFRMc4
aHkGew90kmewr3OPW/nuvy0pPoFgkiP/VKanx3Bd14CT3Q1upNEmngFAVZRTo+2E
JIrhpHSoEZS5WtLfHMrXgnLnKvBTezklo/Lmi1/Wg6p0mawF9IW5WWojQESswWJ8
xUocUx4te/dSzVng6/BZ5rHGufWpKHKwJo/+ECQBID7ZRUdsWe/nb/1+OBNlT9zT
`protect END_PROTECTED
