`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8L/c9f6vj7X/vhcprTZf0Vxqy8oK0eqOuaKXELUwZIS4Z6GWw3J6kAQr4WEwWnSL
5o59DRuaWc+vRNdypISR3duDTtfW+0cfvPCZYIfOHtIgPUPvyNe+6bL77Mjm0HVV
P+KHdzt/jNJUlUjTj4uqTc60Vv4n3zh+jcDJ8vWyekOl1IrX0qldEw7f1rnyY0av
hsiWguXKuWcK9TnG5f+L61vOJ6iHd+4vkv92q0Gd33IDZj4rvDIHEGsu8iWsD+6K
qjvoYfMTnConr3T43jJErJtT30UFhe9LXjQJCQr8Qw0I2+T8L+8ucjDBxhKYsA2a
CDhQ/sWbGlPrg79SkRgZBZdtgWgX+K95DjxGPg0Gwvp0cvPGgZ6zp2aDfV7ZlTL2
WAJ2n4yXPfyuMSkBswJ8EIFT3EAbN7Qh5OPXyneqLkDS1ycdjYdfqFkZxUAcB6PP
tp8+5ndz28ozUmDCFPMALbDDX3E8K/ur67Dc1bSiC3FFH2Im6X9Fqf/9Rp/q7lRh
cxZLpu/zVucJbmTVQom08uUxCiNYzgOO/K0+WI8KNs7zDl5xWSGgsg7U+PEsFFB7
lihR2CIusgHfxDMefDPX+vz8uq/3RbyKhjiOEFVKGsDyOdQBPxSGG5yKMGk5rcpd
8tatKGYhE01Rxl658Z+tNSEQZseji7mcfIAjAZ4U1T3lsOdpdvBZ5z+EGXbqP21s
N9QIne1+ZgNh2pQEbzc/5n9F4z0D3Z5oJ97gayKHTCzNd9uqWw+iiptGOzGrj5YZ
S/p9dMGOgrUQ6Hu8IB351TkZ15uChWvs56bMfEmXRHwT33r0nE3sMfISjLd/RXWF
U20nHULldy+d1pd433dvyzq3Kto1RlhAM1FLnWUKWfu0EB0jAfe8GfHVhD0Gd73z
5P2Xw+tcPbNqxXp5wxqozFr8bqWiz7qtCWwnI7omikhVOu+3icirt2bAEIkt2eFG
ze5tLKpYeXurhQkbs7DgdxwVQu2bhGDG0bR+wD6WI8/CR6cC5Pnk7U/1K4ZJpk+g
big3o2pU/s4KpcTut0fxU/6YWGEkfPxHZuG8AYPMxqM4uxj/LkuLz99JumKJTEEb
vmw3u87riFr13inGPjuhVeqSpcgZmCREO+0Xg/qkRPF1ms7bDM8ntL1xUruidoyD
Q+xI5eF6zrl+ztd+oDNJflO9btNmlwF9ToEz0YY6HUOB/qlgZWyfd+Nfy+7o2W0B
Y4vts+oodjGZoU5l8qfEkG5E+dBF2i23qezdxNCBtJEaAfYW4e4p0UBPPhbb5Cn+
uI6uZhBjqaoXgD6jAlxFgaXbbeaNBUrglihPU1ayH64Cq6OACp21Zjr97fMMPZd3
D56yiEnuKIw3VkivmgpVPI0Pbg0S+OypIUFhXi1xy2MOy2OO92K+MiBEKL8USLy5
`protect END_PROTECTED
