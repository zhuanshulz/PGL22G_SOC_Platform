`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2nSs2HcVwi5jufmKAICQGAk8bKwWqTo0R7Us9Ete5yORMezAoDM8F+y7ahXMwYAi
OrTWLKT0XNzj3ec+lIw8gCxET/slRod2YOTF7auYtQo+3eiCG0UQw2j094nMoUp5
SmTop+F81P6vrjDulzLYEyycsREbq37ZtDock1ivwbqLl01ZeciD3KT8lAIpiD0j
knpsLvYxq6LJVfuRADIA1GqbBMPTpvFuv5qUdQp2rlPJ4eyVVCXPPV82EiComHYQ
S4iOzxF3/vkRklcC41j/nkj0ufaE/8dWvIsLRvd0opZPeG071XETt6PAs1Owvhbw
LUpMmW3PHl2Vx8KMtyHeqTXMIGKEmDdM64vPULwVxvOgVyrix+TCQWxwLGbRtIbC
o7CcQpfBPfcOESmVR5EfqjBKbxtLIMopaptLLlG8jZ7taqi5K09evzfFxEtgtIu8
iFsKnCBESLpQO0sg97m6H+Qv/9SJwGnpV14Nc6uE0Ct/+LiRUXBQ+o26PRT4555Y
blF6Sefj8jxmba9DWybT5b0dLtwzjabdSSyaHUerEU6WAqmwlG8M884Hsb+WCvd0
ePqUWJJlg/WdgsngrXEhDp9WyN1jRvbL0sipojgYek0qJyXsfOKmTdepVKKRthL2
BYmCwbfPGiqbVLoW5mouxxA12ScDkPgrwlLqp2HQe5MLk6nrwteFE+pWvbfDnF3W
qp4e+T4Yawki3Vf5hQjMcRaU8YrcW1sa0jn5FOZFjIsuBv41ISpMv9pCn5IC4zrq
tnMD4c4RAUzbpkiRJHNvSMubMUp+JrE1MwYU9SqH/dSqgzLYH4SN6benqY2Ne9xL
t0vpw0qb90o9+Ukar0EKaNf2JErFuKuX/0NWMWuQls7bZThCwSnE7eipoYdFGg/6
3tZILXRN6bizq3UbGIe2daiIp9r7P0txjD4IcFhsAniLaOppHSuZSHhw49vzgK5l
u1OYEwDWW1Ed7JOHzzFV8vuDo8GpgmTaRUV1l2jS/1cLGX4hVe+YDDp9zqqpXEiU
wxw+yH7K/CD0PH5XLsJDSN8QsCOkqKyFmKJO/eYGadYHHsLrPRmT6FSWjVyzKRx8
Xbx1V+YUdNTonw4XBTA3rDAO6U2zZHYe0wZKsj9P8q4cobDLuvMS4JWmi/RdG+9K
CReZbpuhxiiGqtOf+pIDzrJn5HP2tic/LUjOulUU18Hj7BsWGjfMGhWbiW5p6jxo
s1nYV17EWXQ6btmkWMKABO7YXFzt8khi8H414sEgDq02QTKbzjxRGpP2jHZSXNkn
AAgtFPqpDQWEzAVxmg1bQSeOW61oT5gkrD1SO76CnBL0ck0oZgPMRzZ7amOnV4+E
udUsjgax9Uifxsf9Dnfc85/HRQqJvS8xAyors+rylRk8zRoqypT8DhuDsGF69WMO
E7fm6q1S6brN288TeXIhKQ/JgL1lftdFGjoKt3ZywwjyidZpQSKoZcYr2ZzMIbuz
XzqRzru+AD/0aHkiM56W3MUcNzL7Jkp4Xn10bmlarKh2i5sr0lfzntwtfm8+nFXZ
ILDriuPiydwidpw6Y+rblopNAxF0wFYPFjjE0mgVef5hUSI3nQaRfIeKce5vxeKA
qqcJKUzhRivcQ9VnyrvB1Lq7CQRzEUvBxK69XiOr7xvCPdDBq6YItGCkStb/b5uy
fjeHeR3PkG8RztCpbRuddHbDrjNd/c9g6GZMAjqiQbNScFXZdC78F0I7+AwhT8bM
S7TbbbHxpxFEewvn4GA36fd4eP1SvCVFeFvItf74UsnX1mY7OhYsFKviW1uWh79i
D3WbmlgYJkJOh/5nTloQXCezyyf9dR3CTANHufBp0ycurh2ZjGAbdK7cfrvKN56A
JbAhIhvbQwa/C+GLe0VRnVIUOgzsFLtUlYJRpxUoveqoMNuhSh2zCrbMxxDe9RT8
KJ8Ea76q746/QVMyDThlILVoG89tkvGY/fdgSd9dV3aX86q43a8xAZmvDxO9NyJH
gr06xYQjDwSC29c0YJ1nVOAJQ6lG3V6/fKz+N5kL91gF/wUGsSQnpUzOOc2TfrGw
XQZky7Ndvv+h4U2b25v2naHrJfyu627v/hrbv7ay2M1ShrlFwgIdNuAbjj2epROe
pNJMWjcYFbmO3Q4KC53pHQidlBBqh7rzORTzo2fgVnX7FjIGl2cB4W1wrHVpbj5u
uYZGLwNogShRCbigwJmWUKIh5fpRVuy7YSx1um2oRe4r5eRTYZiQWevnclrT7MqP
2Eq9vF+OqEoHLvwUYHULwyD6Gl2oHRe64PbWQBLpOerXiauGSCzUjsVsizniVJ/R
MWPeIGTGXBPbrjAaLEuA3glq6r04tVQG3E5EmuwnvoJB/Cuw9opzslq0RfmWKOJ/
CfRJiBRh8VfwPvgvMxQGcVoMFxdTjITfLHNRwSfdHjwbYzMoVkTHAyAtMDao4CYB
6W3ZfS29t2WnSHy/MbapJJuYY/Zdlwed2twQq8+jD6XfE4Fh+XI2RyyKUTUTheZg
apKspS0D9VQxWG4PIxOvI71hMFFq11N5IgrlQrQPHFdR/RUin/VYy1WvO6cfb+8F
xPjUcmY4qcE9Rob1VzRuOWfbhmsp94cOMX8YgzytYeV4gCg5hINciIats2E6uL3t
mPVRdRalgxGpZ5hm+IQBUh/W4M4oHs7xQnopqt3e/mYwNezkPmb6PMa1weqFndJg
0asE4Z6YYprAjmJkKENh79BTE3CR24L+RK1qrJ786HmhqHzjHB2FtsE7JbuLrk0C
jkyWv24/F0N3cHym5ai5uZFR9uP4qkzLjWWIlgp9qBlfLbvCNAI0tvw9YVMUMcCG
YxwnUuiLBPNJpgwAIAeoTDhZyhdWaXW2OTIUmQx83RaJTMQ4QN4CAPfLHvaNPPkW
TjYdfXYH69k/XoNKLDZMcxDrAXRIl0unaV4JjzNNe0+ea+TV1YNBecnvsSSw8nqv
9LmBfuczXeG1T8WsEeEsgzyecPGEeSMbBaotJYkBqMBbrK11gTHvH6WGAvjmEoUi
VwdGrah3azRO9zQ7kUa4CJBr9iPsK+qvMZQvnWWvC6pQ0NQwYziQVmrI8dcVkbHb
BB+fgVEoy/e+E7ZYS/iXq1CN0k6vVFIU9NJ72EdRAn+d40Xm1GU7OjnOoNwJyzXU
b3cN0lFdsLr996uKI+WtMuw4D/BCih/UHrE9tg/PyD+T39/ktyIwtR+2q58hxxpP
d5aLqEpU5EYuxHz+d3DI1hIWEtvHJXivZ/TnRDczSnBBV7WMB9rRSrq6NlSB5ejf
C6VuUBZa1+gXk9S8zNEpxODJ31nGGkcdRaYAoaPyOJmAizI3k8vMbE4wLxW6DJ2L
7yGnQAga5JIrha1qSISOAPXcgNef8AVdOvKuE2S2owic7OTXHpaBrVnUEBy8LJhd
+s49F8DVgKBg316pD6LABGg5Ps6ItEHJcEx/3IDOUgPlG7ZkpMFR/meaO5wdRPMQ
BOQ5Wt1R6S+s2tE1uPIauyVfAhkDva4GCvzena3Yatuc3gcebRNzLcx8ys5UhoIW
kWGZ1bnGXPZZ/QmndYMsljR5ClgamL8lpFfj6ZTpZOw6bGN4qKjrlBNagi3VooTb
+tpHLLh9aFmATmrYsnSxeK68ipLrJw0IGiAL84OHL+aocryZ6rpEymeXzHTfsK0s
BcrARQC/tGlWJeIfmhR3ZUS+fKHaPByELGjrMlGF+bC7CyB+K2BqzYWRODL/N8va
JcJR2tDuOHYazlVGlmy+RRSqh7qKAg+v+HXKKBnftptPmK9eyQMYIkL14IhqXDBa
/p5U5S/fLOxSEoyh112g1ST64z1anFBEYKhgxD7uJ30EdTa7z+8RbIWYlkshirgD
0hpmdym5L7AUc9JAmeSGHvkCdGaHfe+4oebxj8icHqwfL6RDEpBQ+Yfg+0UK5kVX
fdiUPrDq66rH3+3pcTbWr4u2J3mZ2HfVePkz1PcDxTjCcQGXMPdz3q6PmYZzxTmG
gMJi8INInqO2kC+Uk2vdMExQZkwXZHAVzLMEKuQjs8vAqr8Ieh1Ss6U1zfKnzPKL
4ClLZvL2UN0G65UPw2hHSQYyEzjMHY2C61gX+Wsxl0lLqw/A2Julk5Yk669138YI
I70sJoXnD3/rwBTl/2qP4igVrUmTJBiHLKxA1jp1EUuT9gCpj/OQQPgOlgDqSmsP
54S1fIxV/gsHoM6iZD8ksn0ShixBxFoKeXmXEJ0UFwqEcZOmUaCceBKsPV883SNs
ss7rTmEUvmWpR+S8A32jbL+XS6kYDEMI8E21ZyV4XoI5SKLROaiERitxOQoeqbjd
dJ5xa4/feJuIn9SifBM+ctIjMvc5wUBayI4benKZeFE4cVtaITuLtmFWzEE2lYG0
iJop+1IKs962XwRSZH4oFIhrCfgsixcbVSfmdUihuQkPcYJV2immlkldc004qfh4
9PEBuA7bKw9lApKebHHlywLp/LCh43/RusYX6cKaBxYuE9gii+Zi3YGUUY/qasUh
am0Shfl8qqwJlM0yN2xrI6egiS7L0sYlmF9BzpNalTjQVoeGDoTGUs3rGkBAPw3Z
Lg9O3kVYzraxZprg6VzLX+VTWfkC1LR1lMIqvnSGoTIVCB2jGodTaMN/CDALujwI
qTCvBk7/TbjVS1l+MBZwXA/IzLkucWwrvLaloGygV+QxgkbMDhTdo2xzJv237eut
9poPIFSWGg6RlGdps0Ql29fKxsn2P29R19q5dCgjSb6LI1VQAMDRWs8UTBhfqb0H
F22yyPnChtVaek8ipJcubI/BA+oQjNRRWGttYE3ydKxB5GrMwNYTixDqkTn5sVkC
+blARvPtZvgfOYOwOrZDZ1DRFDETEWqdAueo4GCJ4gf7MOeddBooHQj4XXXODwGq
D3BBmzIU0mwtwuD4MeXZfqMTAFI0rfgRpwzNGuu+J1uFhcwAENf+PxYdvSksGqpZ
Q+GIXIzwlYIGW2dZqxSzWLfAX3Z27inxAicUC+RENodCbyutEpoI2H8+NVGmFKLp
ws6wkachP5AMGr71F5XilWzC2ocwzoFRvmk5NwU1S8DX05C03w9bFCnxARlpkWaE
Zrise7DE1+kgL4ui4+tAy+b9xsfOR8QwXfZWajWZNzc+4b8jFAcmnVFB5IicVdAA
NPQ3uLEh36/ZsRTN9MHRwy2snU6dODeusjQae6abU6TSwhV9euswqvypt8Q3nDaF
0s18ujtbXLQx2uJhpxW5jMIwjBKAp1Eg4iFR27nNQ4jnCsjH+0l+jVzhantoFyht
q+bvna7y8tksNq8jcYPWFRrvB4IfwhuldS1EKMeQ/WZlRE+Iq/TmLGMY9SEJxj8s
goSOMnR4O9xz0TWjmO4EhW43DRab81RGGJXJWbnbNJOLQNC1dBgUXMElCkNS/7pH
fHIdssXTQ4XF6LEPM1IQeTw5NO3/Whktacsrd+oZSmbZGj2R72s047a0B/3ASJvb
BIHRaCCjXzA6qIqwFDJi1YK+6tOq/IYbvSEnyiZnzlwnQhsLLXqBufrAN1I7oe1T
j9O4CBWZsdZFkWcG5ZQfwfSDt8NbHpH4bqTN0VkqWfaGgOJg0KrzLG1XlROM7sA8
TKvjzb5/j06m7pI1tGNuSIeAveCyCgOiTO3hHkJvYcUOlSGj3Md5VHKYVeljNjYt
2U9Syasfzk9qxeK2R21sbcnfMRXSxixQWjD3ZqVvNsTFszRYdwOEU3oSknF7INu+
htfRoOyvrl+X4/zkHSQRSD2ffp4vxfTMuUVmiRawAiq/tJIqjUDS0SyxDt0K1K5A
QriCDQ3AZValvE+DNrUawG+o63IN3aExMaoWgSflHf1Wj5UOLVeA2oY4+dto4iEw
OHPR6+O1V2evQbOYfEK3PSkYk25LPZgHheWf+7FZNhKt8TKDRXROubmzRSQdG6A/
`protect END_PROTECTED
