`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b2V9ZIwytXtn+pRUdYk0BCMTOFdg3nZ+8uYvLAIZCSCTvLF/6tiNeeAiTbtUWDTD
+FvehXaoFxgEyt3h3W9VTI1Fu43qT/5vIBlzGYw3C4JaZx59r1HkTXkw64uz3Sm/
/GSR20KGP9qECVLvY5IYQSSnpRlhGSuwZtbdaowwUVtMooDGZABO8saovDPwrhRy
1l4D3EfHr6OP2SiTIWG923hsoNMf/eCJEU3g5RNw8svz2ktWEr/YOv1EywCTeih1
s6rQRnN29Jk16RYHi8zCJEbl5BiXCTJch1zBA8MggMTzXGkgjGtYaVfLKpeaWgsM
s2h3bxL0QoF0A63sji1ATANu9difMSeiB9qhwvqJf9CERrBAbDOl6QOSCr2atym2
RDg86rHhWoH89GXTtAIqHYaUZLeEbsef2ilWGzjOTY1Px++A9yB8BRMuRpCnZan6
UUwpAq5b6OYBPc4xBmHV9jPN8HY9yogH0ukLKBB6frLgSI2v24mfIfLMNWWkvzj/
UV+T38XZK4pEIhzSvTwzZCAw6btEuuNgirXqGZvkGduNyhwx5+2sbvwMjoy0QQX9
EcXg3TP4KA80m/7oTlRYYExren902J+SadXoIxJ1eWI8gMnRCGDLydRfQA5L49XV
er+DXmvfFqtskpAMjy+XXMyh8sELK0z349EN3OZO/9nf9I9w0WItu70YHMzry+jM
z1QrWrNPghDnvu1YzU25mvfIYeper+aoonnbYXmMggFAeOvy/zcYzsRM2hFdR/U+
KGRVUn4Q1nJ3BLSZ3En05M6EhOKiypNeHfC9sv1VyDO8NkxP077UJSz9B9zu0jyw
tuyn+iGftrNXJxESVJaLb65AwWBO3oPMIl4RUxbb7VslZtCrkbt4uVrrDrMeB1cF
qQeEl5QEa6HmwWBvFGNZ28Emn+v+fADzvCqfbB4STfjGVnA3xQGed2qxTmbznEeW
iWhVsx+CBThAtIbQl1jGF59tigSZ5noSpIzv2ocaQiv7iXtIHcRaSycG2bpSshaS
BeOv0p6orIncN/fClbcXRjWPbUof/hnW8FZ4hqA3w8QU2cI5BDiEyy6s4n4Tgphe
hd/xES1OREGkwqnbvWl6aAqc2xKBDnKX70iNgzfOTRHSf/8yTFH+NSYyGuZobCJt
fqzcfqP1KDBodb1O03CZ4iiF5MFesv/F1Y+WjgY7FJgD+8NOyVctnS1/8+bCxYx9
8hfJn22Ph93/bKk7P91VNlKOU3BT0DUBGw7aZVHu5XRXbchNIbNtcOxUC9s9zWTx
r8dbv4ifyUTuda2b3l0c6U/DJi0+ULQaJl9PYUgKDEpbAnrXJ6VBpyKHMjoEyCjN
PwqnVum7N8ywKbqAb5YwoAlEPpMB4N5iCm3QXUb11RJFiSJG6wW/qPg15WFva2JP
01Xp2VEuGmOWG+3z8hFA9hzNNBVcUTXDvXJcrAUmyEIHtUOzQvpzOVD+z7AvaUZ1
IdOHMX7WkznpZpLvDS8eqo3DA/sTjrT5agGHjvOH+bnQoqqdCtvqb/Tg0pCN7CUR
CsOOKZVaHirNVAE1TEj7CJaJIMjXKFI9pCZNCpBd5WOaKM8FKkLoGlBJmSyZ8PVJ
9vq06gwTLQTs4UBHfXMv6WBTWpOMqfm6RWUvKHUADl3sjwxFv6t7k9BWEgYmiS71
fTaOgcRGFIY47g5ITpfj/b/xrFfpYPC1aJjX45S06zWFua67QYj1YrxnGhGikl1/
fpv0qN7or4+JL5hZQ353wSj1fYpp+NtkKdrMtdWP0Tlwx4WNooDM2Zv9qNQ6RTwK
ABxpj8QuhuQ7YTYtlGzk48vFH93vJMTix9ojhgj6Oo6WgVep8kJ9qfVjd/cBUx4e
xDVvDsbnFoH6zFDqBjcJotu3yUcx8+TMLtK+iGpOzZmry9itiQjW8zVqojxTO8Uw
7g8pUe1JnQ5thNNzWm2TxgtzuJXDkK/3QofWDrQARGNqz6BQtOG2fw0lypCzTgTJ
jrp0UQ4m3Nmc4mCNSqBS944ahG8Ea+FtGnW4LadOTYPlYgQOLzBPKVOTFV4v879C
v2r3bUWQc/yU1uvw8GioYERxTHR3XGhceB/xn+Gw5fwc/KrX18zcQplIoQ1I4xxk
ZfHV4iQnL3VJY19q6zTPxDZ2W1UdxfwFfcUvxtIvAkJPNBWQOIfm4XMxZeWRMzQ9
9eCfbDeldOmBY02HtV8wW/LpfN+00Qf0ubBEvKAZzl9DVxIlX9zARNBKTtBU4wYi
FvkYkaNCw+dD8lJHG5bGl8fiT3bQtMtvBsuDVvJG45EzeKeTxBnEeEL1lyDJ/dI4
8OR1sn+s0apbapf9CeNWwcto70rCIZhsw4vdBDNd+fo=
`protect END_PROTECTED
