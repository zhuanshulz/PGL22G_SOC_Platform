`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I8HBOzGpFbt46jQJvu56rwtT2yTUJceKPND0ftZU98tTvk1betzT79jtXBgVhHWl
uexd7887Ex4XFN761nRi6ay9tKYE9zFDKMDXExLCebkDHB55NvKIVYqF+NtOI2Cs
/cyhoNv9Fm9EbyycQqG1DU1VCky6mbACXEh+vmiuN/lNe15Q35eNws11zdoSfa48
yqacJ5KJeHLYaxWvpygLboroovYCsDXpSYdry3ACG4YtuyONtWRBWY71foNwPv4a
RZdBLetj5/nBSwSrbBn21vc3MivVxOVOKOu25BGBb2A3TMhba9YM8JieDXZWkMXs
41GromcPn4yPEbEg/Ks7fg==
`protect END_PROTECTED
