`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q6dV7tjeOvqH2we299CNI5qDmnO0j3ieE85AHehNIkqzLvtscVnMppryJsNa4GEa
GWQ5hC2xspaYsu5HRFHD5zf7/17I2G6k7S/ANHdymRjoMlmsE5SK53vWEw0xEQKb
E5xBaUXAP2PPh3Bh1IECEgtvoWNQ2EI+J29LaMW1vxvRVBf9Ex/PkvKqD4rcgqtq
QlJefU+v4GjqrDBKeAGWXz4Sfuz2RnLjAO0FtTjH9NC1bKoFU+WW1FYPdnwGpmLT
qGv1B1vuzsgTYE2PV8sstv1jimIOr0kvhgkCeLcIFkiXjCnhNcYfW8l02JL7i7UU
55U9k47BNFHcSEjRwDj60IkY4F3zDTFmOyezunrjAqscPXthoLrwuLm7OEhDV+wG
IwfnCLzRcjBz5kAz6u4NolDVzHCOeteQfqxpJXzn0qwHrFGFnJxsLl0RCL3qj+DE
ChQ4VVET+VRIVR09gVyFWM8awd8yN94ZTyzHsmQlXXcta16Sf6l74oiIIlOCjoP9
DNvSm+0bqE9L0NAODnKZAMpnGVZN7n5zvXCbCz/NgPZJs9I6hCWcQXxiCJqNpn8y
G2ZGLPwXQUsaIZtfB8haogIjG7Nz0ivRB7sB6nqlsfdfWa9uC390DwQ9gMSEU0Sv
GwsKPO/ArVtWhKy83H9otQETgvoyvWUyYunTO4NgHeLCleoWNGhg5lWC8VkLTiYp
HWdweQo4TsrcgkW66momnZMEZ9ovNxJP0NIl3VuLsErkY1qiD788JRMEP4K6nWCF
GW3d9uq8Ev6wjOrU0s0b2qfAJ/vefaLQ8TJZyK8NFuEU/cGkRLWyy2wjY19uLuXU
B2JJOSofxIuvFGqp+MHg8ak4cjANlAphhn36dO43FcVBiyVBTI+fC/UKOWaIAizd
2///DJ+MkbWCX3CT7cFa5JSUS4+0ZK5tq/Cm1313KFpumtLEYeHA3rK8RnT13kEy
hVFnzcMJ5Hl+PEjsoYq4cUyBDqf4WwOqKhRLfmNBSWhXVLsQyyACqKYaY92fuMJr
o47hFU1F2yiGuF+zWWUomiMApo3ji3SYhreYu2GcxIgr9pqGqdeU4PfeOh94n2b/
RzCaaNarT8j5rhAT0g1x33qmSCQknyQJz0Lf/c6gTnwh//ONGWWPZOdBML5u+ywq
sL27NVQPd4qK6HFHCY/+HjPOv9pYqksoLgTNiEr018UXBSuOFunBluiyHkXxT0be
zQ3TxexDzRqKxJtK1ifr2fakwwe64udgY+3AXTWIuHfncstqKflSAvy6ZJEnfVY6
ZUTTdCZbBAMsG+aXVpyfpatGhBfhPk8FvFObubTVdYWiE87lMgCpbPamVFyWo+LJ
iGrEF1b7dbmSE9CaE6bgUunOVexr84hioVQ2kUGr4tg=
`protect END_PROTECTED
