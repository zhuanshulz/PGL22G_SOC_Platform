`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rKK3sF7Suib82QX78B1U0XPjHra2dhgXtJ+JWst/Xd0UfC9Rt/XlxcSdf1fhk2/e
aA600CnDBD1Ebu+Vqq2TWmj5pNoMEwN7ynIYGBOlkjWIZFpMB+eHGRlF4UvVanWt
HTr5TB/ChO4873FpvrmSFPbosQKdR/h6sa5z8J9/ZAHxey5BV4leThpvcVsFsHXf
qCO5VtQW8pA67fDgyvEqLe3LA+tiXHnQiuLeiGnC+U49gBKBKFEXFYEFKT1A95jB
1al18Bw++TREiCofwypVsOAQyf6CNnbly2K2cywt4aWRbIrKJfPlmYvfn0/MgZt5
PpfV9bFPSb+YtLn1qULOGW1Vmn0IMeWzFFpx4+mELrS5A2VwE2Fufs45nR4xtngw
CK36RJog0EcK/TgMoSoMEGFA+Szp3MdXQjWlyVLVnq3t+2QIR1b+Qax/WxBDSPdx
TvujwIrI01L0557UmuwPqA==
`protect END_PROTECTED
