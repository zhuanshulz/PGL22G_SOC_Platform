`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qhxgN0Xsjb6OVuqg8n7ZXJ+kFUkgKUmIURlFGpB4ua/E1Fou6r2ypNLRSh1orMyD
3XEOqxXDjMi7EedKuk5R99HpIGGiT/UFAwONtp0O9VhDdTvz9kggkkL/j0CMyibV
xAj5UUWgUvqe32eITgKM6nxiY5GcEZicUZnE7cPQ+M6J+HwML8+nGtNfakWkuTXr
enC4aTdqbF62IkXnpXBd5+ePrZCTFsxOkSgYDxHJaphXcoQ8hPllmn+QL4Oyab3j
P9UO/DC4/M3LLrZxG5viYlf6a+GQ/Hp7IOSVDeslsFC1Mjnj2YutMUtXoRhBwMPw
OqUUcPWSDFYt5i9Oiu4vM/anH7ShmpdX9uk+8xv8re9GylFY5qVbblRwSpwGFtb+
czjnIpbnMWK8zKFm0NqOFiCdepD2ngTOFsKfwVDsyomkT59NfOqH8dwEHyPG1846
QsqpszA4I5CY3yDm+YAbv1Sn+iAlJK7NB/Jhb/TRPM/t7L3IDcNyZwCZ86Zp/+TJ
V/aUZdHWc+DSHGXtbg/yRcyFR9kcolvHmmFlMADs0h74VnNumGTngWnGkV9sC0BV
sycUjiiEfzc7gCLRplS9pG5xzq6FENLyX18Ns10m6LcmMEdpGy4dSFxx0E0pFrrn
mJ/zTylDl3Pa6XBDYXsca8k/X4VR1X/jveQbwqQc2nsKpwym3DUJBxwg2i3LLHRM
Hd8qva0CF51Am+aY47DpVMys4PyyU90Mgj/M4URn70ms75oSmiZAxsBhLbA15cF/
gKOu6oPfcwr7a2fYd9DxcYNOvd4+aF57Qb/+FT/2ZTBFFvW7nOE1UkyHcYmKfMQU
6ScY12ruCRw1+zfN/Djzd51xAwv0uRNAttWBwgki0jXN+ajqK8bZjd5L4lAEU+Hz
5V0M313vFPaFWj+n64vSdn58IInKocl2WkkkB/3o8Up4FQNtRHYXI5d/pjQjnsuO
NzZ4Lp3PDoAgvTW/eDDxqy7NoW+WMvvw6brJTU+YpREyTp3IupXoGGDizsQ1u0kR
ETwwv7lRCr4LksQ/+Jgi9rDGAh8RQTbRjuTlQoO4o1FbHg2pUkTazc0/J6ZoFW5t
8MFKa/QtLRUD54nZ/Cu1N9uahL6YWe16oaOftXdRkCJ4pOZ2tI+nNKR5L56fIl83
A3qAyNfOAiFotk54aJZmyeUY3XT5P1Nq6cKqfKasacI1OQK4KZmktXk5TZ+sCFTB
AUA3K4DA2iPzW9hfiII0TWL447zj0/44gf54PVY+5FLUqI9rSymLSi2YqPSqt4Yh
bK5it/IMhQhhVtnTe9f2tM4wEqFNERBd9RGiWyTq4p+b0LbHDHRKS8Shy5kZaH25
hs2CDJn7lpSd2/j/fUgsKkj9FVgr0hWgQGBGb5tNTct99xSIZMTZqhewLzQe6mvG
oIE8EFcfsCZWsScpe3vBlsxwCBpApE9mTqy12w9ouG4wdwWJG0wOh7l0Ei3rXa3J
0JapKEthaWt4+ghYmjwRq1htoILF4Nm6QWFsI6rOhwmww35/sGWMPDhXNNvq9orf
Dpi0eC3xeYjb2RAUpz4ogY566uffRTOLCg45XlaA0XaoToK/yHoGP8ZsKKJHUdLI
elVa6tJb3ah1I7fwKwpkhB3oRYrj5hLKYcNPtX9lly2+saIj5hDYrWV+V7qVvGB/
bBWrhLX3Daz0qtEpbOiHxUcx1h3/E8dJWj5xQ7ppy3u1vgd2TqH6N55H2W4YCp2C
mDPxP4irY+D3b5x/NRUF4B7Jc75tkSum7NT6MdNBZdlaFvYPztfGA7YV5c/8/OBp
VDP1jACpvL9Owi8ErYkZnnBpCgubzKAgUUbZsZN/taBLdQB2TA8qBS8grjGkjat2
9RHNHx5Glv2zaYERudydVb4wQrv87Qv2OdHod5ULb6uq7hswFUSunfRBPn54i/2U
26APgzAdNE54JgvgMpZFKOHocyR7Dczj/K59Z0v4DHNGxbT/qBwOISXD7VhSTUx1
hZF6UViM/xPQJpBBdKwqOtAwHqVUcLyBLPBdNd9gqecK5pe17FEoSQ/bjE2x3S+L
DDlrSEn1ev3SCQ3lBtz4tZeCK+p+lpRu35QwZTfQLxLcxBjIwN7LmFcWIBhJeWt/
ufANbOgm7JX0B9FuJD+kN00rATnVl45BqsZMrL6iE8Mf/8gjhV+1wFCfsrz3fUd1
jLgFux1w3eFElKdsh9YfmexPpANKI8DXc4AzybZV4m8TwUlG8x6wir4VjZ92xOGd
Qp3FCbnFAtpCpLv+l23kpLaE9hTPbTzqLpwflKXYBprETNPrd31HAd+qAN4/ShPD
k1Jlic4Q5bz5tcfmS2cjchGpQHNEEFdL8wJJV3YUFCEIg3CAJhDYq2QubyDCCAab
3V8NHuVZK5aEjC5XxG/98S/RJSqo/bnhktKsVKYgQv5QZQsylPSs63Wg8+vAAGhs
zzQu7Tq/GkQAliyLpG8IlguepKZJFKlDV6itkb16cIG0hyZFI9RLRYzTrwMEMjYq
aXZa8kWFAF76Nj3mlvp5uYfV5q6NSWE/ZIf2AJebOCiMcWXIBpRe3qf5mAaSyn/u
ny77jO7pLQl3GVi2fsXuIdKSs/dvDywjOeJ8uXzPKa6N8z8r7mVyCOEkaB0jUoyA
hyuendPE6X34efrfiddpUDsS/rFm6RgGMgU84slWXYi2YIig15P2ExNdsIJd8FIq
sFgweHYz6NTUzrgXFkx6w3cNDfK5lUmlx8zU7DlYSppDBmrlnO1W6SeNeWi1sIm4
RGop9GkMzM6Yj/SOJMfoQ7CQmjUrUhgZ43zBT2kk4BQ8JgsBguXG1hUxovFkWCUX
gY88CnBLCN0s2rN2TGsrPQJBNaxrCqoDqW+YyvMtgae4DMFMvKzVt51NGQeYyeFT
iWuyQwplf1Nbn223K1kn6OyONB7lB2bojc54dMj/HFiy6PFCAE+1FFlv3GNBHUjY
MYfp/OfNffx3SXk88wMEE0mYBVe8529aS8QaSGQS4pwiWb1ssSsAjVA9bjTB4o2M
B5BoOaQwB8n1wXFTc9g82fWhzLU73sIXcpUPdpuMwh/9NelahAC23xykNAY5ksLU
CFLkEp5DAUsXVdiO6khH1QCdvsqpYfWg36KzHGjzQiAblbzDegmqtjTDJO7uR9M6
Jc1IRIdbzslDE4gbFqe8Ow4vtxCbmPtTL+Xjk1iOqkL95ttvXEOClavz51hRqENz
DtFW1bpuUf6x6/Y5kxxlM7kmK78MRzUdMxx5pU76PwIZ+uba6490qog7iTlrJ1EI
2AWcfgXvhmcKVY33iYpyI8rivBH3jIGcfDKCQJldxikDmCDZcHuAxi9r6NwMaf87
oMT05x1Dh33VDUlMKe73CFTzj2aQj3rYbbXen7U6m8ttBi6zOHjupemnAQZfOhnj
ZrLiyQdSA7UZNVrXac+EKNfum57RrdTXxheJ6IjbCihB3qseObhh6r4l4v43xIWX
0UTLvwcitCsRRYJfBqfqnl1dhHXpYYr+kFQDRIuijswrIiwVZW5NGc9C9/7AT+Lr
4f/TamONvNSCMPfbJg2FTA==
`protect END_PROTECTED
