`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OoLdy6spnAB60P94xPrikZ1M+43oOgpQ05GHsKB47c4ZxL/zgZh47O1Cm0l0OIAI
u1mk5PVYzfnQSjsHqEcXU3rUxQZuGs7P3WdR4JJZn/chfnVmy053RD0BDsnqqWjT
RfyOjHNoU3lGwJSk4Efvix4OmgLBQtKk6LhNri8RCgE6Yi+T8mb1IpXaziTlDo6B
bLRAmWWvDXHsSkRqxmTTEmDIE6Fq6ZgYxTqcBo0ytyA3mJf2sbSKkoEFOrUX7nDU
UHq1SDu3gU1IAhGR345oKS9LliH85eYrqDUbvTcI7dihpv0k+C/GAFGFb4eMDvuw
+k0Ata82hEE9DO2kXr5cGnJqJ+Hbj3tlGO+oo/a+904NfgnkCG2kdx5d9lhVb/BE
ygpdXdp0HIPk5557whH4NEzKqqhnjGj+Rl+ZwGDRD7Q540vOu2DR5h8ld0PNNzGD
nmlSSjmAH060xgXFSd4LPv6tGDo+v9TtMZKPf/W/PaIqw/G5KaWIJVyW/2Ldwwgk
qDtYiY5UrjgkwEHD77XfZW0hSnae2WfslUJCqqkn5grRgkFFUmv8BlatZQ7bq2Wr
CO2djUAIXC3rAMOe4x2fERkYOCloedGXOrkwIxBZz6Phsz9YP7+zUg7mdE4sdG/5
UPlRbRdJixMDenDvl0kxyxSNC3vNa11nlpKi+NHmcuTpyXrubsq9xExaIe2eOxJw
H6GGPByuP6aYV5FggF+TWQ==
`protect END_PROTECTED
