`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GtOVpGRzyYNGhlLcSZlgcmbUC5altnTx1HX0uzHjYePgQU0ggmZ/dbdu6oA3M4jp
NsmcoYnYiWwMsItjvScPEoeHBpaY5tgqt0F4CRVd81ZH3EIUxrlY5hjaAj2755wY
1IRkFeV1MP8hAv9g+2MNOI7D+Zr8prr4H/YG9AVjsb9MxVXWebkez6vJ1/v8ZE2h
xOmwzRkDCYUI4QMPNT2AZruG2C+5nzNOu1vwId7lxgWgNRl7RDGnv4qbn/Kmh/jD
oAq0wMjgNnhXGfj1d6GN7PStfXj++H55r4mbSsn8gdG0tOAVTDfRl88+IEeuLzcG
c+C1vVt1+mcoN2B0cO/yBHNyJw7+lNtNTMyRRQd2k/8fNNE7zKA71IW0vO0h/80E
rmECQq+ATrAUE2tpnptJat4epp49imS5yPoElhncb1ddEbw3j1BWcqHo/XJrFD+p
NkAxUzvDymCeKZB2V0Um/vK7oEXzvhciUXanacodH8YKSue1KhIehwfxProYCEwh
ZMlWmUuX1yPORJHWRFkY7KmqVYaQtxUap5tOnFSou69tKOYC2IkQcZ4XiIaNhZPc
8jPyPhGYFvsWStKrXDqfBaLoSWRlPk6lhLYqIIyfNNC87bKiOV2JbwOxjdeH3omg
JNW0FTLNwNpM4jpOcRgkOMaJuReXdwMQXt7ez7zevBVKFUXlpc/XFLf5mUAJNMHY
sORMW7ALBNXbLvETdbBmCNlwteQGUitNCxjjYNNv2jsicPPEi0QILVS6k6QWi01q
3d/2LVpcxyuMr4hbjLZFYuw3GlmdrNqih3VH2Dbcslft76ARO7R2fde6Egc2UoRJ
4MWGntRUAY7shwdvMQZ7iOv3AIS7l+AeUIGcZ1MZz5jm13tgUWuzAC2DGe8XeDlr
f3d9S3sXcqIHUNIfSj7sYDJjI9da7pyPJqBteCAPAyq+P9rGAHUBihqGhmxxxCc+
jt7rbN1vaH5bB0Q6hJSzAH8kbHFtuZCxkrYeexm/CBJElm6geq5pbNiuT0sXSSXm
pYlYXHJuwgblSEVxR6Aezz+Z4nhD9JscEkgngdDgu9ogrXUVMJCX00UapMbcdV7W
ZxcUiLH9FIDShDi7O9vAyeIeCwt5IB5/JakbkCQxu+3qhxmWipghHwd6rhaClt5f
jMqfcGXoQw+qqNMeIGyv7qR1GuxWF882KvkOwShbB15ddEdmjq4h2gCp1ZHmShnW
`protect END_PROTECTED
