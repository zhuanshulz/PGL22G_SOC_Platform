`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7E7UV/XdIRK2a4e+F2D9HFTQ/sPAoU0biGfzpGAgRTlumAmwtTcHDuUamOW15n9y
lRxkbBovavO3bn2iDQSBeqkzrCxrDlkHicdYCEEH68M/i3Jr0Wca8m2rJoJJq5hi
MHQXiunJlGFtk11cjmV+siUL+TcjxoBFZTVSdVe8LK/JRZGojwz5xUzf0Zcim9Mc
IoXdCSF/Q9/VbhldhKjIqczSwVyrcfjIvl9JlL8mwojktu7V7UamPzZQwJH9izkb
`protect END_PROTECTED
