`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
js4S0Zu+EXyHvXWDB6RyWY9HkS1Ef7lNzltnMyOA+0vD4Jd7Wno/+kfw7/tZ9dE6
E8kTPEC3JP9QplUQ4/O8F8EcM4BOfy/kDqKwigVOlOIBT+VXbV7+mZ5US69i9pPY
tLuF6ScIfDeDZqVGAUxANgTFFfOPOFB7hVN2b+4fzfcbo+s+FzvQHm+clZ/jIq96
DKotYk+UTP7JlQJOpf0gTXqdsjjE/QEgQV6wyBFF3Cbc71ZsBNOp3/gLawsIt6K6
WLgmhYJHQswf0kJGiGfmeLaA4doxRuZRgObzjKZ0KWBkgcnYmPmLdJGMULmh3s+G
4HWh7dWbveAZoFVZmnvJ9R3mjNdSgVVzSeGRUyysYKKHp5ere7+GjlbdRVHBEKL7
lBS9HqFSBr70/UtfQtDYEqW1M36IT26bXDSU3FZMP92hGeHl/Abpw91XUbas74Jp
Azk37Iddo2doAVipY6e2ahyKIQn5X4WGT5gkESuuROFnUkWwBH+igy1A3MueVYb4
egKq8WUyndIlO5k0MR7pradKWPRVqvn2F7udHOeBEW6v+PIm8WoHLbtKYSCkJGiQ
tRYSpj/RNy8aggBfSLy/OnEwn08FDG+pa06NVdF3HI5BooJNmfB3FOIW9ZwhSXPt
BCiPxwzXTGBumSbKenkhb1xSATH/aG9YMI1V6B6djMfVWhFyGEsxRQPr1SVMniZ7
X1f7RCkjHPRhHV3xiwLZ/fJse0a8Zidbwp9w87XkAWn5BvtSNqMMOJQ56YstjClK
KFlcU2QGPqMCPXf+nj5AWGZjY9jTU7RJKUvDRB3TZ0+/LvSHstzsK3nnSFO2KAQm
mascae+N75P5WHGscAs3npg6iWYvkbi7wWL2OLKCLx0fuKRqrTc5H166gITjMBHY
/ufvLnJwmK1dSEELRlwut/SVFvRkHrDyDqttNJrcQ36ht2PNEOzeT+NM3ABIp272
1c6txG3G4+gCLhn8WdNL4r5lA7tIfMPXtKUPsEu0QVaV973eGwKy8ZMnCuOgbX5H
bdipLga8cnjhzHGWQT2t2MkBLMSE9Q4mfRtAsW2I3DDTimgaqdKZhoU63iboJhlW
9jsd+oQJRb5JnLEbNqZo0vkMCva/sA+kBChiH9JW4g83f64CajtQS0bVVqeB1OCt
qyzKPAXZlQMI4Ags2ofYr+Dfr1vjy0H79jSvkWEU3UVTuBEWZ6hDIguUqxy/j4Gz
yrPtS2ePzd52qHYS4iXv1tLQUfvue/pJEYCg265K33AVPMs6Lct5OUeTsfZxGAze
d2LbNWGtVte/nhDmWOc45NrGWmUz+VRtAq8hW+B6Aq1cf2rUQ4SHG8UtH8JdSyRA
DWWpObBX+0K3LuesIHRRhevLive3LyiiGCZAiyTVyKAWcpvqigavkN5JZb7ekLDP
jCLAB9C07H8YgUpGLIiMo3bRFBofE87zKFAFGsYndH3ghyTCA6fuqiN8PNIla8fg
KEIWW9GbsqQggYiBgGenvFg2b7XouQSI9TBcVsru/jePAURj4JZCS3LJc9uMVljG
Ifdm0Uq8zFrUovZFy9VDQJeUkVvGbAa/XislWpyWZlmrbHrTGXd+qhT/4EAND4Iu
b+vHyxiu3HevVmMw4hxYcgElW7l+2aguYrLEabo9HK+kR/nVfanxR0HWIvFaslGP
QfHslxtdimi7yR68X68wfKaxxyrBGBNezY5lWBowIOw+Z8GHOIa8tas03Bn2sHcR
npIra/Npu0RGpbtwPtJH/1JCm9TIAGQ/h3KEXmb/Lcu0aaexJqEkaf+v/BBt1Dz3
NIv4pIzWjTZggtuIQZJpLLv35Mx8btR1aKGHAnU71CTKnJfhK6DSyA6ehO5/gJNp
7NTOwnavD0zhp8GWRDXUlbPy5CUhyJ5z3fBwFvHe4NHPjzMu9uDSibvP5MsX9HFO
PtjW3Juoc68KmHb/GWsm2tKotH/6L2NwQsUJJU9yWUmOCyahn5vID+26v7GzdpuW
ak1NwlfuJg+pHbYUlEudPslOmFDa0UFICW+6DXbO6Jc0eUB6W9+oy0RAzOieMIZi
nuP11B0igwHUA+IuWytgSC0l33BM+XUsuIRzFKGb6UoeDmDARaXVjvMKA+YFXfJW
nc/kX1YdN70jbjq7UJRzHDtaJDw3OsR+GpijoE6wU6lMXtrBGa0xIiEpJ9++ya4e
0TAR9e98YDNEn3vHvdnFMfBmCp9/mMW5CmZmTz5FZsC74LHR6xeErJmtsmwVyRjU
D7N43yyud7HHs5Bq/5Sw+Ogt54D78Sn/tVz8x2ck4U1wSXby2eb88xJeIUwmApM0
GexmCKenVh0KbmpXZjHz32t2nFuaS5Tk7Cw8ZHibk5HtiK6YlweMn7UWNUmXme50
TZ18qEwfOP6fRVpsuxAbW8SegIRISoWLscbwMnq4jRNJZfIl2c5P1GH0gvobN7EV
qwfcWIFv5IT4p886ZU0qKWwDiZbkNVkKKLbcg3MhoY8NCNhzUb70Pt8isUXKE911
sANZkfQkISlY4tNP2ugtIsbmWk0sYTMVyAKOgdLRdXXCLIkesrofBt8Mn0nuKYNx
1nzZi3I8XN/amwYE1mt4XUePIl+7V2Buk8xszXH2XLkjujRVW5ggm+2pgRV1W7lZ
BP8QE2hRVK4VLLwrHqWvEc8Gr8BpAuJIPAF1OsssHFILoHfChtujeRw0Rg26Uild
TMnCqwB0q+3uypRlCxagZh2hVb/HRE7DmDl5rnYGy33UyE+llRf8ChITIqPSa3td
CORYR22OigHmYbMRK/SdeHGM63RWsIo+mt4r5kmaPP4qyY3TYNTkBznVubTZLejH
n8kdzRoVMjArXOQBlfjc1QdC968I+mV83bn59RZvkXYCKklxfsp21e14j6TuSlvO
53HjMSxffukUlaxXhs1P8Np6GDIxl7ePH3POO/MHG21XmPAxofDIaOAfH3IFGYfN
COzggmtrT7jFBND3m/rcFV+3ZW/3XHGhwKi7tlkPVutFWo/zZBIGsaZ3Enbdh0ua
+imzwefbMny8TQRHnarSYT3J6CeMnVdi6//J9J2eqfbKVk14YWhQM1bYrrkjjQ4g
BPqOj1KCKoOHFWi7WPj6GUgBZwyL4eFxstsDG7djWzVeIlTH9fgJprukJYXOow4o
2uJ4WHjzoOXGtB0+Wp9wqhhjzX6rISzaSx3SR/9U9cCDkcJr088ry1PrSwyTRbGh
E7KxI45Mk5csZCN8vVyLFtN/Z/ZsA281HAtP48t6s3dgoDQsOL6y4t3Hsh3yYkTw
pbffwbN0UjT7U4Xv/uxT+2nTbVUsJp6Bga0w+qFFQVIsy1anpQv1p2v7l0BYINz3
SRq+SK1pbgvbnMoXLbu+SjoR+p3bvJm1OD4ObJq3lUCda/2/mDvGDD8cRsFpobdD
gM3fH6yQbOe6ZtMLZnxTnakgI0FGqsJYMae8LinnHABliCo6GHQ8b89mX2caHYym
ivM2LtpfbR9oEyC6OglDcH2AcX6XJfD8LoOKZVeDEq6nX/QHvKSNEySeeiHl9h4i
fqMLvURPUxQfMof4sVM5wlzcPEVoypfVQjTpKGZXhlY7FQeouDxqH/1eZNlrUEwu
EB3nmH7frO97F3/phdihSwMh/UbBrg1pMTllCxdg11JqgftpfCr9448rsw968leQ
I/jT9m+6H90NTz1obpC6Fl+nqDaaE0YUeC2z4u3EQNgGFefONFpBxel9+vZVK4VF
b7Jm2eQjBk/mpGJyu9Hfv4idHASQUV4M4PHN9DDidQutMLUR6o5qIqsoF/9l8+Iu
eiGOw1ljORIsHDQbTlhChP2dqQ0NNbTbfNYKfj70FTvHRwwljt8hxSKACR/L7DKz
f5bHMlDaFAbKgaU+zJrNIYz1TikpcY7Q2C3pDuXeIexmoszsnf80vPDfEjEPFeQd
GMToecwbHnoZv0hZNLhOhwhaFo1NPA7sVe4fP45H51TAiL13mZoJyaIb4dBtgGNg
Z20Dhqd/8S3xIqC1v1+wnHqoegxGVikZUIT7zVNqRRmrdfTvGbH/MEhdSfPYY29i
TjnRiUaFua21YlbYIUtWZwWbM+drjLsx2jgBRQQjmLlKNRdHYnXBq7Hhuorv4M37
yJFTzSpVlrX7l3322v7l4PTKmy3iYZcKhZG/Yv2xIoUVFXrSK67bda4cNIYsheJB
Tvfnwwkrhl2BfCEvrzWdSNCf3DLfK8l2ghG4aq++x71S2FDHL0fRjWyvgZRjAd27
DXTckeQmmyRGN2FTn6MlSpLv5xcQYfZVLpRUTcURUPrvCW7zEdHCeZWTB/Wq6HDD
2T87HYrgaVPk8LmtVasGeId5a75WOCEUpRmhzq42MuBKoD/z9lu4NmKC5P6v/DLf
vfnWiCAFK8T7YF8mN6vaSIOh/cVfDqLfFD9YutcOh0mEZMnkZOnhC2apk+Mh7WSi
gbMdlRCQ9tg8ChQHjDy1IiEWFNyTSdxFy2XoGz20UAyQ3JnE09anbMudyhE+8IDL
lb+ax7AvqYl7SXqDyALUeaq3gALqkPvjczRS4KOSQ8JluvGU2aBsakbqf6J4LyTT
UE+wCRlH6XF5iQrrPtHJY61kRQiUx73t9Fc0bgQmQzH16Zl7c6dMeegVyB+FDQgz
DDYcJ3rhlpLOzo5MH11rGe8CdnfigtPdAWjeiR9RsU5nyu8MQxvnxdvKZAgZyOFn
jS6hRGLp6fD8VGS8kmHijnlGS5rXfLKsmXpTbDI5C2YcK42uG/pj13UZUvRXPRJy
X3uVNg8GTzqO9CZ4Dr3jd1AbcqkRAPw64kSE+tIH4Y/M6nitA7JbuAhgh+MCTnXz
vECUW93tUXuXOB1QVzSgq6u1Aih8SzQa15jfEGt/lzGsHWOKC0ki54rFiQ3FIzXo
yIbkLEVljil3MffYe+8HAokmYNeV8SNZXtwEf32xj8POONVSSX3ms1+I/JlI8XUt
ZZS7LHoqiqdEOIXWoVnBYoF9dBNJZH84eZ0DvvcMTp9EvU+tT1sth5fC6W4/Q9ZB
J/Z7KG4nswwXstpyKQk7Ms6gXeVdWzLj0KFQWtDfsU1mvGh11ZXQp/+lmDCDnpuK
0H5dAjyek1GlcOzVadWlMI0/CYBIzlg4tUBwuyIqegDexkI/tT7eijcTW8wCsfKf
cJvKZIQWoM0OGl7GXqcYXd5Eq0+bBoGso4LgH8of7SRwQRUKxuanMwgC8oOYQPOz
W9dMGkp9vC6SAv0UUzV3t64SGRxJ7F3h+hj3Kzrsf44Llc4TFE7WHHymg5aWilW1
vkWyqbAUtpjXz6S25jcYJ4psLGN2MjDuxlb/Yu+Aow/yHRtkyYGoxSPR0USv/kZj
VoF4sUFzmnt0KYHScGJtrWyxf6j0Npc3pEYjqpEn57YFMOvt89LVb6MGll0iqtvm
7s1NHht+SIMqqE81EQTKAhsPmyK4Ln9PWbbq2s3q64vpjzjLiZByb1yO482uhZZL
Zf+RzAaRgQBJDXaa3KMDI4ymQAxJdTKdm/8k6ZfhtHl0OAydjwfGeK5+4GTRYpEb
6uie6qBziVYblGcElh3w/3/K7NsJmz+FK6m5yVmwnmGpto4ropNR81AYiJzGV651
EFw68m9jOX0u0zPTUtvc3Wb45RlJ+zaZLj9POmO2jCMSesuX8T/9i63Lbem0DvpT
A/5udHEft5e7j280YZAOFCqCZX/za3pXUaZlKvEOLdsX8IFiHESG+H11/ITn/L0u
2VSM8Z7G2bvH6k8z3Knt5dvnoZFcPls7aAu2tugp0wU8+azrMGX9vjjcyR0d5P/b
7i+fgfJr6M2/3RKu0dX3ZGso2dZRzPd1e2e11VUoTDzqLuvI95c4XPCPnsGLGGT+
h14iy+0iXDbaiqt2XDCBkJ7GxUnUmwR8OtzNGPRQU5Eiju28es7GEwGQ62+HBGRY
MpIZOA1GalLZ2e16VfOnDUpmG4vfovlOcIWFO77tIXH0QakWMm0ejkkIMSUO4wK0
Z109P+F6JctxgG6Xb+HSKrNQ1wwnVK3RMXrYziS9q6xGBz9BbK+DYvWKtjrUcpMV
pxPwrq3bPVI4SO36quYNN9wkGRzj0JVn5ixaLr5jo4mJzwOdDqyHINVF8W/JMGqK
f6xNVmdRuemxQF0hi+rMZhluAJRBqfD/CcJmLZF0AQGsbTv79F3oigsUG5k95FTO
3ZYhruvbkt8Zn5LehT38KTe5L+VphIMQYZuyTRY5bnV8tz2XjcBz8RfEfJzTe5ax
niwsnf3pxhqkw7Ydd2kGQpuHVHdO0GVmnkgQ4q8YYMi0cBPuL3LjhCTLMUhe7xEV
Rd4Q7lLpmI9a8WoGf1LxXxC42/EeW1i2s7eYg7e0yaA+Qx0glmvUcArxNEqQmqvL
8muFlk30WGdZ/RNj4EbahZRpcbkQkQiOpLDwW5XLBVP+uTF+DuzN+OYSBtOO6CNx
87KY/T71HfE17U7rjuQIpM7QJsq+JAOfoUGnr/jO9pmnTeZblCt0k82zF7fek3Nx
v5fQOpl+YijL8Uyzh4FbVCBrQkl6bTw0BHldsblOADZ0tQej/mIfYlcKnJYgqXsz
vAnHcrrj7irWDqdstFL41ai3ipl1lpDWexCwO9zWyA1Mcl7WKU/UVHtijbavrYF3
HY+pLt8SJTiVFiU/pTaudHvwx2oGw+Yhed00ahcK8HyE2Wh28qao3iOo7q0XcRf7
MkKxls1NslOx7vdAYpcAxpQ3wsHF9TGd+Gq0JQbl8NRhBciHgosiMqgyHMNor0/v
A8rg/yazjuAXq7sdEg3aQ4tc5BrPtScHThPZmiLqxGZY9ueJg8eCNHsJwkoIZ8zZ
S8U+He27ibDMkG3BOdgQ9X0ZRNncb8jzkn6i6hbsxG3Tl0nUYOgWZff33BbZtFA/
/+DRFojbFZWfacW3/R0AFzL8eopbYwBfjZ89wadmH1rn6640ab9xJltQx9yumr+4
9F81T8VzrZd14gY+hQzyvQwGV+SBahEe+Tq1fLeGIhjA+eXwEy4++eUrXD6GrYcY
WYSWTsi1FpsmjScaDtdfaKe3r49mKPi0h3ZnSN8joC8CP9PMcSo2lJOQ275kjmFi
GEIohEKZIQVZBIwuPvhAh1PgkO0hSyNwFsnUg0nnADsF94EfRa10qsncBTNdv1pt
ojWj/WJzQ95cmE7/AMUQiP04tYvqB0GDdjZ5FxfxBMPmd82H3M03KGbmY8o8ySsU
OTV0Z3e8bQ8kvo5LKE7mSvhqtLo4fPy7yc7EcNNOhkrl2j6eMwXcUOHW+YYQYlPq
BBzcb+kDLIgBDAqlUheZU//tUluIJOKwQ7hQnukTfAO9q/Pdbwe3x6hpiv1pBf/Z
3a53vO0ZXc07o6qVfv/eKNkFT0d7e7iSFlIgKrVk6cSJn/KpWHNBjVDV+aH5H3dj
pV1IfAh1d1jN93mJJg9DFyhBwCCqO9kUeR+uvitTj0vT6aGG1EBfpWeljvvoZc21
igw8m+2E6W6p1JDjrCCtkEg6CuPYoCIgOXfPRV0FS/BzL1dIatAS4TWjBcvdmz0N
2eNICqGuE9r1fx687YqXFICAkt8arKr0J0ZTvTrje65uJiDB2eMe0Hx7vwynW5V/
aNoMspip9tPcG64CUoAEHHBnat6GbpeuVwQi51SecJGkBHBEgCraFLElXHN3IdMI
qKYjBEFx+Sm6lchdqCEHHQqafMnmRZP+T/cJ2Jgy7yaSlEEa0/Gw7W0M59eRbxSo
YoPx/ymNa4vABx6aP1vXhrkgiftLEKDiiE0ypQdHHDGCjooFuv94vZD5L7aruKFw
bsSWS/wd+OshlYFdCs5Sfl/5s9EQEHhD04AyzCk5lvSQavVtCIcskMHQ2VkVXnZU
GwwiQXcKpv4KWZjrEkMZaTadxLszFnhz9kgEBk/eRibzTUTy2xWgQQ2c8iNvGyZe
+Sb8TLLCAfVSXtBtIqXvH0Fdz/A0P0K+t+zNq6mTqp/ymuQyn3G0Mo8jQ79HasBH
wsRVtXA3d2MSZxC0io7V0oMDrVBwvJcfF4AVh9RyeOKZfSoCUpRAYPXAgMTsJN2+
DsARb5GZ4caeqKlQ3lM+KHZP/h11BtdMFZWjoVWp5Dju9yuHmb92O6tpXhB0cFfh
u6Lhm7RBY//7yER2IPSZH6pWEfxIKz25uQjQpif62fzP3PzECj/UnCtnJi4nAc+7
0/fN/4cKxIbbiXBhgtuKbeKsA7fUf5pa47qjrqjpRgjzrTDk03Mh+ZJCDiTD3ejf
skvzAazkSuESLP+2Sz3TkTmYU8lNN/VuaXntTc5tqlfHtQWssP2XsOAKJ5BJUqv7
Drq+OOaLLjx+Pt40J6HKr8WgO9YvIwikS61ISlHwHhZK/iOoflRfsoBhvlMrU6e6
++Xt7reT/cR8WfGhF/dnamHbTzitOUhiTLYVeKRlQhXM1lasgU77Try0056c31fp
Da3cc5Bi+FH+BlW2DROlihqBNimneXPY5sDhRikjoyOgnlxjtTHnpwhs7CMYz5Ll
zEmLkimdzjdR26tjZPcolUzaYQ/1ryrPE0Lk7Zt+JFW69Kd+D8S81s80YSiXFTDS
BHHkKdxgQRCyWivKtjMGZAjGf8nO3bkyFYGPathkwIH/xvCudLvGH9ZqZShdRILt
zidntZeF88ygh3NXIAcVrAb958YsALKOi8lh4utUcWksDPLZL3ZkMGup8Vor4pgd
Ygwl+g/Aw5haTlEtbzSlzeX/1mQuzsCdiQE91EWYBoEEUA4XBp9GzDsYPgYktTl8
LQa+7vVA2TzIAZw5AXO7sM/+T0R1QtXMZAjVWZWU/6XFhRGWwIiguxm+dv2gi/gm
uDswNKSBUDZ2Tfe9mIAf8HcvaET9eQjLPo8toyp/Pj5E2cKJskNCBzuJNAHpLYe9
VZWoiJVkqH5boDlTnrD/A/Ubdqj44tpu29s4ilQcvyjTL5u/0a2sTSgvwxPqgWnB
KJw2/CzzSwa/V+lNFxlAA58NQWrH3327KIydMQTEMtlASh+wP/rQhjDbMPbYm42C
GzmjVa4HFwb54wXlrxsWLdHDQqvK82fj7sZtDhtd//aTFNdj0Ivs6LVu85WDVlbq
TOCvvmZKQWCSppaw1kbeOCsoNGs++2I28nvFPIbVklVIl7GcXkITiD9LpRHhGet/
km5jCn7Np7SU4PubvH7tGYZwo76KvVnO9QdyMNJ1wmm1NHV6aikxKAIs/zV4jE7s
gd8bf4/1Nn3X+RvPHGcS7SNZH3a+j3Ag8f88PQa++fNSYAKUL1QjmFWu67BOCz+e
KCzVmYjUUyufK5SxBdpQGqCxtR3cSbmortPcLlv1X9hbp8CRH+bk47TmKAcc2qBi
dt3NJqIf9/xJAU6pOw73bGzO3wQFAWH7NapkXGHZA9/nteDB2W2Bpoalo8V51Cve
uVv09hzyrdW4mS9Vr0iSAwebcNU2GhLNhWvTapUQnQiIF0UrmfgAJFoUBQ+iMP55
/eVBlXBmIcy3UqtBhKwkdTjVu/cp8Yg8TyMlOYu5z4wjl7lvHgtRsQW8rClPYlzg
2o6baV4QiQqogAuRs7Wpi34U6pIJ9c7+vHIs56X0V/ornN4Jsvdmu5KkuUN0T4Gb
1P2m4+TFme1vg6k0qYzexNGQCpykfApT+yaEcfVtj0+WZFWuLkvw4ZkKTxYIjf1B
ElWjhVYWVWwdiYm1BTR6Lg5ZO5FcFnkBW6sJsTIq/RP9IbwCeiK2CI7ateGjwkXi
U6cZ1by0AuSImTqzt8PNlzWrXfJSH+y4i7X39o6tuU5WaKkmb3wLJ/af6TXayl4w
31Xzss8iWN+oDEKNqvYKk+YXqiuIbCWJPcVhPCIltlx42x5IIhrwuZ9IFpP1l5oV
BvWU4f/ifXhZesnKLJfAf5LxL8GoDNciJFATSeYrTudRll3hLkG2GUU5JmNy6rpw
Ixcq600U2i9iElDc1SZOytQQTUhY6ZrDK8AKJJDj9j0Xmc+ZX2nAW9Fn9FeKy4qU
6xszU3sYh/HDhrnycdtz7vRHeBNVPmNQELPJDMMRSQ0h30fH6Ia1RarcPzdBx87o
VK3qOPASlpMHLopQPq5Wv6AtvTyxiXhw5YrwMYZ+Ww3nGvDLIMGlwWEVFX6HDMnW
2Tzjy/s14gqqOZjKAKSbBfQrSgW1cRR/wQKqluJxnhd06osT0QwPwzdV6k9g8XaR
KKhGgW76PFYrw3fMZw4STs2LkpUd9AQvCeTdp+4sLTonIu5Vh4skXX62866bsJqT
ZnSoVgFvsYuT6fnvunajW7P6iy1bEsbmIoSUhCBdXAr6ggQ36vCGtoXvu2tDKwao
PjhL9AZSLjm8EKUPal3hRlEHRdi4QnrwvA0vEyMJBagCh73IdNP3UYjpM3xbLtQ2
QPqinV9NUowmDvV65NBlg+2ROSU5wdGUj6qe6bWh0S6/ODvWBWt6Ptr/dElFkIj3
6x34PtbFRYTFQt9uqbRdqg27THaEMa/heUuxLLvYLxFpbKStmFdUMY3qy+izT50z
kiEDM7V1YQ5GOPVRjOgwNEscNjeEBJ5ppBDIFuRQcHSgw/5XY9xyhQnE6zLejgpG
n5EAgtPF2T7xih+99Lzebk19dcI7lpmRfZFq+qiBqWm0DLmDjaNOk6c4ZHslLZul
pmBokomaFQiCY9FyVZfD6a/EpmUOLals5uIYRUEkxm89vA+d0gQtymLJ/vno/P7y
1ah6IdBtmBvT5ieBI3Toa51NRpVImNUplicgHl5ITGYVW51RwAPrHDLVlOdBbmMJ
ysak/bMNzLqHINgfa4ifouuUVDKOHoHCOXkpGxi0QWUCxWQLOHQDsMNWwcT3PAv2
zy5zOT79xJ9iWBWlXJ8LVXDuDQHwV1XOB5VukqyC97079H5wUAVhVH/UoB1nDJJy
Wu4iHwJwasc7czou2gf8z/ZYvm6/nOoXOMWdDlE0ia7xi8R+n4pzi/KJBn9jCiVm
V/cRMHxL9G180FInG5e0DgOW6cKRnLr57F1ABLGqiUMt5/aBuyOJ/tzyZjp6L/IF
wzJe4qvcEw1quwuJelr2Gk+W2eOjZK4Hl/NCw2Oh3inZAQBbzIfnt+8AxohUmTmN
roMIbKmM8uvh5H1C0nlZN0hJmXwzaUXIDS06WCv3R2/Vq1ev4UoNIQibzkk4bhjC
hpcJeMd+4BJdUZloc+w5qBLTlG93uGYaTQxkwnwrADfczk7OfaLdr5zbT0ShL486
L3Tmn00itCRz3EKawpzdtKxTBKnjiFAAWVFqJ7V7lYjF6LCj9yQU80faujo+59Rn
kyPkE6/uou3FVLbCbHzHt97qq5afokNyk6EoREQIscE+4k8N4cXvx+fJXgRuKkdJ
rb8xn+RKwKN5yVqJQD9m3E2OZP1zKMHX0XGy74P3u4ElxnjO74OOLWdx7dVBEEjg
WSq+lDG2vGCzP9x/epazxqUg7hYaWNwCElx8dPgoeagCBMy4kuVQ/Os9lxUYDxSp
24W1QfqfM94KAbscER+6zLDPUdIR//l+LCTdhXwtVVntSsll1qktH5RbWqDZdmrg
5eLyTJHwQ2t+14s54eykh7qtN40GkwhR0GT/I5pFRmHhBK0J1Z+3d59eWPCoPuSy
vrMwQZRLcXOSiDxYb6jvnEw2lG0KHMTF4FhQQoZ/I0bY7dCKyn62plx4Q0MJySL+
NlkbWNGQgKew5/nXu0bLttV802+eWAiFwwTGuOuYZ1iq6PIwqAp+DtzvxWlKo3Cp
LjhNEa4i0VfJgLhUFEUr/NMpQy+XV3xmpWLaSy4xgnFxG+EhjbM6QyLkYjA7Ofb8
jD5JS37c1nQY9HHIL/nM0tuMIqaN7E4KLn4psFa5JRiF2ujKLLkuxLW28OdPb4Fx
lu9uGb3ogwSYRYG/94IUYz555zQfKqX7iOfM/Lr9dRkqROFOrDYUcDapI4p815i/
zA6vMh3McZ4yFmRHFiJXJcPy1gbJkz0xqO4R0pSLpm9SIaYFM7NNmYzn8Rsasf07
HFALOONQ2yOX/EW93Joi7qh0JvMLsj1yVPJxSKpMzKtvOS+S6jWv7Wu3FoO7HjoN
thbjKrn2BIg0zVJ6kDsFIVL3hXlN/cuPd5nXWkdR/JAkgD3QQa+iWTi7sjCdlxNv
RPTOIjP7o9D0VOayNYcHfa6kAhgqWiCR5sExXKXo86fC4JrbBpER7wpZu5XVBo4Y
IrNfquQpCVaLeCy5QumRP3ixtFS2HjuqBM5QW+L1oofNnvpCvxi0e0+l9P4G1UP+
uY6YrIPWQp3RsnzFyb2zC/5+oBmKZYfGyRZteWYEI0oPXyY+9e/kIK6azO62qDVg
4vOp93lTx0vLUQDG9XLXQr7gQlm56Cyp4gPi2ZBkKPmtaNS4MkWMYu0QFYqcwE7S
Pe7q4ttimyJbfuTcuXQrMVyK3mO4nag70bfEJufJA6W3Oa1HBVrYvprP3kMIRVTW
ueoIKUYTdrm0uOfdDth5H2WbWkdEofDGz+srH/xCWvdSy6V/4ixfNCYHs++I1VY6
mZt+Gzlprn3LSeoaElbjNHxfXwdImNZVZFlrOKtCBK1Y+2uBf/Lsn1EZTtG0apxl
oOHBjSC9hJUrcHBYq3ahIUJAUTjZczyDb3myMzjNphB0SbvZdfYeK2eDH5TgxVgI
2a/v9wpCFYIMGy1/FvBCUzNAaCc5vkscEFUkRabUbJiJYrIXSEu1G6V/cK434VMj
GraOEsCQyRA3OdQLefB5EvRmFE9jHujZJE4lDz3I+7UFZfP7tziw1dwQknzww69t
+5tfVsYE6innfGRM7xJRPt36mjRm9VeBpPK1jSxNv5VM+s2G/EN3V5CEXbVCHkjt
znZ+xBTLD6Ag7aPjmDMQDXxM+uBoOD0i4BV+9ZjvTwW9MgWKPv9K2LzTG8XOsJmP
g8lKXw+CtaOojAN8GYJ6DsItWvcfVZF9dhU510IWkf4wERTSlCcKoRfl5b6swPWf
xwQHmibr81RTiagso18WCI6pEwhQPaeFBZCtvV4lp6uopoqYGYa9v4AF8V9FkKiD
tEwXFwqgOUJaA4ofOximVlx3JF9aWj2gr3Y30zjgZ04tGpJHx3N55BjJpKuFNrTX
fuQNDXhnDtQFTPYQDPLH/gT8GQaCfoY1wJtlNZVw+a/0uRP1P6XlNWZS+a/yyh6H
lJYg3mb7UGoMVrmI3hC1q7h8IR5bnCIJMm9bVXgKDrtK1wfl4CUcuW3HFKkE7/Oj
yFrhEiha56squLAL7/CFdLIM4fvTrTC4zYDyFWIFZRbM4Gjk8e79qNWAUHyytacX
Dy/E3LdTN2A26N150R/4NnbBVIvOBuAap1rIy/TE7EXKEokYcFhj4kg3JLWirt4V
MqdEx6DWmGL0V9UjIHniJS7NdbtkSWRw3epFT3wjP1tC4aeUuPPC8MmqrU+raWgJ
rYh9WBYgTknPvao7iJERhIi6A30+c9HupRQMJWbkHbKWd+KA/srK+u1BKl/7+Mxc
s8tv7d0I8SEaoDZzEL7PJ7ZK1tZy7Igjd9ivVzAQ2WVq/t5vBEYFGGLa7w9pUtwb
O9T9XhqH23gJL0t4bQl3YgMbgKNCbqfQRqCPld3DTy3K7c26kJTdYec96bFJZTQj
zWpUbf0MwzNvTUZoaGdHS/Fo8GnYn3otcFdWv5QIRGflAmSEtcR/vWBcNC5ofBt5
lx3M7pxrpLbBaSxxUER5oTl2hmFiUo1UR5GXLZTfkwjANTHEMaHcG3Ci9dWrVv3A
3WqkRxzRdoTyQ041vHD1iMIek8DsZBG7NslBAFqEHiXI0XfrcuOwlxj3gvh1DAXx
QkXMAWnQAEV43tr6HlViQ6JXYdN3idHAOP1IXu3XTeLKXwwUB851SzSiIPf0NLs9
NcvbXhGHgWKFKYcg5jE7GxbWcFaArekezgh/1VliFKeEGJDwxy4ngKuXxMCxr1zM
NQ6WJE5kNQmgsSVYs9SbSFqYcY4qaPbyWfla5LRfZBvFkYaHJ6kOzn1XoMuUcbDg
2TjJpJpjARdxybcDId+opPolmQkW6Hpso1/Bi8HnOp1fv4C5Tn95aQUCHg5czVg3
6BfL47RqEXe66qyLHwrD1dYNpRareWs7K2d1jzAv+/gELokZ41ukDVsWvOJ43fy8
WRNCaISE2U5KZir/5338BcyrUmLSF8i08ci0eMr4XY0juu3s0B5SbHE+Wi0sI06h
2zPeZJAe/AqPn1YElBAZAC5bGWBwBMt5Zom5RlC5V56r83mMkVdoM1qDC97yJN/F
MFFkUfWbx49kaQ2CLyLzLchwQly8mKM2L3K+A66m15jBCUEjAFZOvQ5uW5vg30Nb
ZW8r5lTbUcCwgr7QtqVhtbshCMdz39EsdNWEPGWmmTZjKiqTCqN74u9EDD7V1/W0
8TWwXIlA3PL4ezOwCj2v4LELusBuFRPEvdgr0SawBBvNpJTZK9nKzpEuJwQYVTa8
Z1Ok8ZVu2RqRC14aQNuhpU7AzdtKD7ChBcS9k+loGPIg3WErHh4NHzaMgg89zUw7
1daPfPR6mwk+Rqen/VPu06/MKVEUo5zsLPAO6iFIcR6gpKAp/Y3clT5O+K5/1UHL
QwVq+66qW5n8DcyIeAaLz83N5gU/xyMU1b4XYgHtaUeYJPpqV8tKPbDgRHatShrx
aWETSCz9+lwslqcNX+0mFjGxpNMNBejmQSIX92Nmai/s7CdahOr5XCG4p0PDd3Th
lI7yvTfCboCBQTijbcvQLthfsXjmsifj4orEzx8yc7xZo+JNhV8ScQBN7WVmoXQB
6Y13MIPDsxWvxtS7tSomgimcQDJpxmv0PWt89VfqIDNRqwskAuKLKmZbvfISNF2E
fM2PfCboiCQwuJHQHkqOQqZEzZeeg9nm9Yw2TM7NlwpajHQrJGu3Zaar7oJVxaBP
UIQ11GD6l8xqq1VeYOcL5k4LOsVr4KrPZFyCnYrgMIjkLc+GKFuA7CrLvzG729rN
YAyrWe0FNzVx+j2MXw0qtZeHpt7+U5lT/Q/DuDN063yUReRqNTQlKk52eR+99+1T
KTEOROicEk4l/SwGhRTSj2CvP9PYdXfnh/oIBhdlUHUwsKkqibrrL7Sxz589qute
UwNzqAs1a2cPbhDCQNHoApjPlf+rFrRf4Ty5DY8Pi/JRfUlo3j2XTeMc9hiESqI+
CjpvAQMm6ywmxwxNBM4GX6Q+9Jltpv9Vi6SmW4ls3N5qm5E7XcU3o58qLvdpfLsT
AXSctMXTY90nPKVQaw3FE+Ogm9Xlcolb51xeDPtmMdXnvHTzfVdvR0E5u5VwqTDY
CwBbQMBPd/jAXeNxRcOHIuV6H62D3mKGMB0+eeuBupeHYwcmBf/2yWaMQMjuzMKT
QQd+jQSB7K9VntC5Qw6ZcwVnwbS7n/w3LUP9jeENMyMVX9wZtjKlrSH9ecjLfHcl
sGkUtOd1rOqNuVgI6ImaoEbw3FudM238G5+0HwQIAW/FiLOh24UO73u1lwERCeiM
4YPdN4+jWC15lkKQgmoGQg5Jfp5EQLIA4U+sQfr71V7EY8O0L0K+8O5laJITUDme
XVTeN0PcAgqGm/X7zNq+nT+EsN7rPLnwoFFOirXK2DkaQpw4aWRrxS59NfDmGXFh
AB7Rq/u27Yx4g+tTy377Ok/4P7PfXLPAynfwdeH8B584Fzo/2idhRG0WDEPjUOfy
Nk1OvLJnNDavQ3vt7J4K/jHzhjYPMhx+mTGlD1brtO8kDI5JJaf9BjXCDXh0izJ0
3TTcB+SRjVDXkAFkJTos5YD1iWpfa1U9iJgealS1ZULgNlyxEGkIIPll1WtsltvV
lprO6fisWTP7qvcTBwMY23T8EhDPRhCbOkSVEYAIgCJQW5uWT6n4fYNxve0uagWz
PfS12Gexx4MHMbOakZnp3fzJ3HAITZWQdagT+CDkzfYf5P7SxUXA79kEy3uf7irL
PjbXJMClbugH5ZVUGYHlK9S8GPqqb4dTwDWoaFjuRrEQFa9Sxj3P4DX/GE4mP5/o
I3SLAroaTGzHVv++yiPAfo7HczMgXz3IFEBl/ztbmHt/fCGyV2tjzs/tVJ1gtu11
ttU3XjYHTKvY2hwcKeXVD9/L/oDMslua2Doiy6qxvXUUPiWFI2Fj0flGSa+gNicu
A0WjF7+p9UVNqaUgIfZPqs6/M6Gx2xUrY+NlVPCMTfUKa3e9yEdDoAuOLRfZCNl4
9Hxd3GngKDh5d1wY/EDJg58zjLlrdw0gIhk4SP4LiuGBvfXk2vjjWUVYoI8TAV0Q
FwYbXr1UUaPU3UUEhCr83X8ssUYuWxCmTgQbTqapp4sXhVkjHXeG5P2iQIKnyTBP
qDLp37OwF99monHhJA7CTX3u+fzXdT5NRdJBuILHps5odzfSviZ2j4THums/12jj
ovYpr77j/+K8W7edCHMtWuJzZU2po96GxUncE1r3eWUCuuDAxzLr8FW36kkoEanO
UwKYVr5hgj9yl8+v1grWaC7BwMVU6qy7Z824ygAwsOC22wlqwmlgR5olkqy1tNus
TeezpCbKjpRYigLYa2iV1YVsbHrqOdSUICZip/MtdcNne30d7J6qB33jI/zpS1Lz
zYRZYUYH5ALYNjvmu8XNe07wspKv0VgTeTO/3QmIHu9YWbsZLsc0Dm2Of7ZLrmjj
C1fVw3qjH4kdfP5ZgiNsLP5R8fmWfpINYyuSy6rwntWkYh1mceuUtipUdjyaKWBY
ygBwYdaP6naTWNQ53/tJbnxpeD5d6mEdggJ3KuFroHwDKTNMPfjJW1EwxDRU4XGQ
2zQpuJqzwe3uMBOryhTCixi8zuza9yjKQFDCRgjnndutFXMqDz33LYQq4iYvhePZ
mUot8CVUa3gC0y2xzY6mt+F3rr3bJXdIqZYvrWgi4Hy4GcQGZW+2sPLYyndEyZxF
qUjosyG4wr09jMkQERRZWSdrbboMl0FYJKjHe2oooXlwgXBDk8g49aQSbTwvdP6G
vqGwY53kLwiMnWNM71mKu75hO8YLyKv+dTrJpts+7hK8opvUNou/LGez5YHv9giH
k8uyD/UOGFttL/TZXAmBKtm9s6pYN82GOqMjTgZMtJhe9Sv2yG7MAanTmFQHOai3
fQTq/tMVqw+RLMEUTaKRLMrGc3C8L2R5jHgJNYhe+bac1tEnO/jOo09sNUuvgO2l
PPOZICwg2La/NBkgaSTdu8ItHbKoSGR3c0E+oUOYp/JuYDdAM6FgcSY4r3BSngiu
o3vchzbBUW3grje/n8/1NPTiyRx+IMlw6zf9y1AEONbtdihjMhtfidkWkGIgnKBB
owwaDQicDfZSp3G3IvUtw36PFGrgfxQLrOvKyOlmPc1TNlBB5qdvon8BJ0PYCqWz
WcdK5COHmhuigahUinVdCljFoAZ9Js/xEjxK6Dn9LqvYgZMtLrxIii4CjFTNjBW+
cTzvASeG/gRtgPOb+dGDsGDrVkWFYGsmUXGU5dt3FakYsjENa9m+6KZz6h9U1Z+V
aI1b2OlGvzmW2ZFAI/RnjWSR5qQEWYn2fU18W81PVVTZ9Akj8mNwBJg1ytJ7jlcI
1BTULyAaQFIilG81BWFeHDZoDCp5Whbvzy1y8i7GTUXXh835yEGSDDnQf43oBgYc
Qb1IAi2n1kzo0xL8QQoeLxrDTK7mZsJAKN9p06xjWvmaZMgxgHDvHC7Huho1BBHT
I55aXmXnSZ3pU1A0FRZkCUYzN+FurX7M7wWqZHeKztGYzZPqx6aRcvKZwKOJH6Aq
wVNluUfJa84ctQv5/JA07yUUyNLPsBCEgw319q+MSwvRUtCjEKwG1wd6BcvQdlzl
shiGWtAj00kfeY+jdicRgtTvtdaHzc+vzJniUDbtQBLEs3cBJOo+s5S4Oia9z3hf
TzI3WVCNLbEvChzy+3PXUEWz/bLNA1tuxXfgXZe1DtjQugntyF7xmt/gXJng7xJO
haZSjYeP+JlfzZ86hye/FacqOFz7zbhu/y+8t6MFoxllWZ6Wze19BV5TpOcFyIlu
Zw4trhb55ZJmBrqkIBUiESLiKUbVombGo71Z/0ezKQ4KOlTzBHy+yVE5WE9iBXxz
pKf1Tp8TQbUNNbB0Y5qU+Z0BcI2WzgAZtQzE98XbbyfPw9yQCPzDFr1lgvZ7QbzO
Qi8WTPXoXzzuhQBhdQH7DqDWCN7MT3P6xFVzfm78N3LO3qdEGhVrwnZgH6FRF3vq
69O5wB1rQGNUfL3P8mDhFXEano4Ccc88k8AxQd1eP0Dwj69DjK9MBXIl0/8Yzcxc
7eTWNQY75k6V39LmZlcL04VBjYsOidPZ7hs9dRoyVGaiP68lsqhG0cYEuAeNGYzD
/we/1TO4rKSKjeE1JawRBa/DX1W1f0TfAksvCs3MOgJp4161+avBhslB1abX1c+m
R71Zw0dUhd6FTJ46NCKQd45zsXGkvhsvX4DpDi2HvaxQ/fS5GsVIFVWTJU6YvL84
o2iuw060jArPssr7WVzR7TbaSD7cMof2DKF/tvDChK6fRQUIzI6as6sfxGzGnc6a
LETrXYSVH5GxezoHimVoKzbWCZ0uMAxTP98GJ4CMl2f0rT1xdAUHw2hi3afYxch4
DOzX9iw+Zu6/YK4u1Rg5LT/8Nw2NGUkTkhS/JMX7kgt+J+szEUbAL+joLxD3aPhf
7d1IiIOpout7vwHhLDCVViQBp/5nGNLPDcWQAp+43VfrQuOmn5GARFljnp3hmklB
Rj0oKeMI8c1pSSkJ7jMeEwdIaZHwgpfwkwaiaVq4keez76POZDYvFd17WyjCl/75
fS+Nw9/N+ZzxLQ/1CS7FMefNZaDU7hYx+fZ8jb2rTZXwzXfHwBALJC5AGovrxBzE
IlerVTwjQW7H9lxeZi8oPsJcoXpQaPaOAwBd9IT+YTu+D+X5oJ0iO2imeGuQAFmq
LbmaPLMp4fsSDJS8XPOqst3ylFXMc8uuEVdsb/TmKLj/5r5s3NLT9zolO2e4NdPe
9dKjFM1VdbJefMXkwPny+P0G+1Lj36iWv+ULxlS3Rx16H2+cUoyWt2qz7tFBDgvv
kkIDa0z8eSOtips+a40kVl7WKhQ+VgGU3fuNNYf143BJLRiMbI/y7TL3qUkgseXC
N1z+5rgygM3+Rn1JiYAmYB/hKPXmtdoNgfkAUgRQRygD8FMMWoKEuuZjBdzQ76j+
3kl1NYIv+gCyW+RtCvPoK7FXeu/1JU5n9yXwa+dYAEjRA+keqcO6cOg9FBNgKu8F
gT64v2rZQhXhq7OVDTVEL/EPymN9cd6cUsvhOzdxIYQDuJK2RZHlp5aWbbZI41qo
p2nHW5fsQ9LgGLF366/hr3rawMVTPGAYVeGTdUlaG+gSCQlV6kLGlFaN8n1NzQDb
G8arl+OLZYrzF1Ah5/YDjzy+E4Q1IDNU8k8bYEHxjJ8CbLiWjurCmrwuBdYmmwbe
kgX4sFqosgl5Cq4JaqiVax98yPqdMPZfTm9lWPgQVCAD7aAL0f7MwKPCusnDvWi5
yDsLruR+pH9x+C7/jugb3zZwGtbg24/DDz4kfsoBI1SVcltakTSdOdVaPoympsLO
+ex6OUd+StfW712opgWexc4M7gyQjhiYs3EK2ZfzIjHXoWfEZO54hRodksowGM6O
GO7tiz8YnwQbGl+N/hN8OD+pQvUS++UbF+OfueuwhKG4/I6gVyY0MjeOEehS3i9z
9L/Yf0pRY9lhy0h8uJ+cmFGEBV9pGQiJEodFQpfCHeV8AigLBWZK9I2jWdHXs5uQ
ydCkzZxeKIglOQmkPjoAzHIVgkF3Pfpr138SFiUJo1AIuaKjDO912lqS2+WeZvN9
WrqH3YLZGrAwJzqXy7NLyumk1tIEaPMbpd0dWdnsrD24WWNejrrjxGh99V0X+Rop
qb2RfVfV6rXTuqtEgoToJFlCZ1O9WrpJ3YUoNJugTMfNWgQT03HutF0ydwgW+NGw
GfRj8NWl8ZCCpJAOlJYkP9X2CERifuRD+dPhtWObZHYWZZJqWuOdtmzq0jkW7nZo
f3FJiE7teJUBDMYpr0AvzVvw4K4qB9QdOl1ejldCEkYb17Hw7pAeXU3Y9JQmxM8d
13yfW351nyb2xoQ30plF7pZLnMIf88yPjlRdLFfcTm2LcnTPoQIXc7wYbR5hiM94
y2MHJidsFa2KTR1iGtlY31MWC5OZNJ/MJP/fyUJEgsvtImA4s0lDXgqM8OsXUq+a
fEc1iP0WpeXbuWxoxb0UrYEEcQV6yBXMkviU4qDaUQ58NxbevRhK22O26XglRADW
aB4yNq8kAW4iypZA7MXeAXehGOjlkaHh1jpMjDDppRLmbSBsBCi9K/gS2lHDbZsB
hZgXJ7Jyry4IWGMMsKB5crVGqK61oRPDkrSCbLP6Z/NObHdmNN4YBPDV7ktlF92h
ZqPgiUbG67715RwV/Jxsv8hMzO+liCoTdBtYjA8ze7ik/xFCoD6FA6kFH2MF59Ge
9f3YBrfGAG+1alWN9CwpTKndV1C4C5a7P+IANsqCWUwROYERMKqr195NFAKtF7hQ
6gBYRtav/sNi3h174KaVury40YWrCiuDrt6iEIDTL1jbnTdBkeg5phcIDRfnSBss
895dC9nBO4iLARnbdkurGfigas5AnKwfHRWRhSGolcsjfX20mJNkVXEYSfWDTQOE
T+KL9JZxHSffZouUtM+O+cmgRV0mS7xo60yJ66WvqjBT5fZ9E8Vi8UEbhEwgTH5r
GFkRw7HjQBrvwvDqEfPR6A496ZpOTOXPyy2euCO0PYCM2XZJKcHYuGj3Z7I4MGEg
/66dqBQcXjeqmpmfLUWvRtOk0bFCWfwvTMXKupl5cajwWszd4CLT1Xo3EQE8Ql3U
LykKsXfwItXkDZK7YSBnoqGG4w/jPNGGc5VDRYHcLL2Dvhxe/L+TNBpflF2CIOQv
PPYlsFNYgCSxBDR56MOOEPzde4j3tJSwyQl4oXrupVnQ/e8waTGc2RZhKmCEX3Kv
uznJgFGrXL7FGB0W+o3nvkZA0X/0N9aUfg3rqpQQXUnRYUEULyAExYC57hnMeZLa
VCZxk3ui3DISaENdjjFlpEJMVQ4VLWorKiSFqGKrymoUM1ApfCatSotxwoH9b+tA
H6NAK0KHLjNz5lDV+Eyf142r7inJwfUK38QIjU55xBfdSH9PlAl0p8SkDgzvwcYM
9lCp4eIQhRdAZcTEf736SY1/ngZxgZA1IeN+YzHpubizdSrx5+CrzUxJHVGZ3YOK
fr/dhlXZVlY7LYzjnslANCE8Z7KyEma5BQbmo1pgCAal4QPYkoWZoPG8Uw+U1yvB
wElMO6U4A+IWk1mILjdV4Y35kjinshumuTocgPeBO65tZDNt4fezhMVCOb1qswn8
xxzryqswOzryOozBau5LNOAQwkW1/QN4ru4XSWUnpcBrXgyd/PCPtRmnbsC+dU+3
OEFzM66YpkjCnu1CipgHoNjCdyFSdZQL0OF2qakqJUPA70TBXl0zhywvAC60o/yq
otZYZJG+4dAs6vDY1SEZN+59DPlcaC3VcOPfZpL/dWFBgNVXbA2jwF93ZBeTUJTN
NBA+6N+dEPMSnQqHKAtfkEUEjaPTttwHKLztKWQQLP/NMMdtntGA/l3bvOC3u2WQ
WTnms5MTmDfGmEIOon/jh/zaAsIboQu0VLRn1IpsYjoNhWDE4S1CRaKTWcrZeNks
cJwjIIWSHdaKQktlf3fK/Mfe1wrLjLaS8S6LZuHeKt2JTNm0QoMGwohBQ99Vr8VJ
SZZBCrb5nG37NioJXhSf/guiimp4P0i5G6reTJUicgnv4MhKQWOjI9KLXq3RXPt/
XBzX9U95Zj6lLSERxb3yFUzq7HOmbeB+DVED5J90TXeBHC+adA4FfbO5hkVznLOp
E1gXGhUYtJn6t7gLMS2WY+YaWFDv1UYQ73XkD5YTd+vcPXF01hJ5MdD9v6yX+Q6b
0/zBYVpq4mvJZB24X0JLaa/cOu0/ZBbLD6ytn+Hj/UomKGbiJeVEIaEn8HwSD0tb
W0CIk+achdUNcfvRLIyPYRoIk0LnVoKPkyiLUhCaJyupUUffTMk4HQ8y9d2/KD0v
MXthTn2r9Cenahneidv6xcoQts/ehs2ii59LY5YgKbAuKw6/sulZWBvIFyfNhPNw
nJKXUSJKiZZZvG+XkAQynHLNGVEADPkbZtx+2tQjjno2k/S9ydP3yhaylQW3fWdC
HeZWVrz2n0Z2jmu4bExLlKXCxo5AG7Hcl8KuXjBtrLhmAuSVUEA/3G26C3xgPt99
EZA/Q06eYfLrh1EGARfwgIJ63FKuYiLxKwgac8bCsU8ThOUEET/ZoOsrmoG0J6UV
6Zpw5/tSBZh27kFp7SW22ArNcEXKXJ1UeQnlsYlnjC6cB+TfxG5VfAU+I1tYeU+1
PLAwSI/4lm8OQyGMQqslxIUbnZ+mx9OUqx/dv/H49CufXvwnbmHXS6B5dzj0Cky5
/TaoAsPN5jxct3v+OWdjPIO+807xfD4Wyx1KYJDp+JWvbKlPZpt4o4+tJHKqMqi+
CYHCi2J/Ow5fg/ykUcZ/jbUd52htu54Phgci6zf093uaPt5Z1jIXQUp6DSMuVtwq
7qtVmD3twcOemlYG/at2PFem55sHSFAbofGS5P6Rx/rSEdA7MelOQhp4EGGCW+mY
lcf5vr0A0DRPj6U3wtLBF181F2a1RrS/P+W6fnRip1i8mHTPKjQ8/qymeDzCqlJA
J3IzNBo+UKZnjDu+VeUfLq9VfzPwbHgK0whoEFcZznt5TFjX2RdBTjLDDPDZ5q5F
Fo85nDVGiXUzBxSGFhFnXMYo7TiOI+FARag/J8voXQEnaJQQX/Cq0kYs2EWPYDZ4
E6hRkticAws8jwKgmnPvARgOcZNs2IB+xRnpc0g5rCjbaJl/B4aOghihyaAiSa5e
FKcZx59iFzGjuUmTROG8tkVj5AXpTf8WuSWXptvFpH2scAtrDksJsKuw2jUs43G1
8QmMsE06wcZQAXQ9Z6nVZ26wFN0xvB/38LllMi+SKf0PoAw+fnGd8RMhEnEmZro+
72I20jX92++uEWaBGB7ry/gEgZhw4uSePnMTfmoH1VREOPBT4GqMRVIm8oYlQ4Gz
b9NaS6KitZgOj9R1+KnSMYSyxpeTUdgGZvuSJJ/60YzToAEH9MJfA33KYRfRz8C4
Rz6hF5e6MTUD0gERDSMUG1qS2LECYmKWOGux1QB/M00sIDfTqpDBZESe2EQtB/LY
kunLDIofQg39oEIW1gk2K8vxUS951we0os3tZ08RsI7Sm8wCTshi/iwokrjoYz66
q6xe8fzGyHhaKFOwp6QX0mtLofqEvD/8DwyWRuu14c/JuQoioF72mcX8OJ8sBC+c
piVh9RVJAlxrAfmX3xNH1whe7qX0HsZAH2SGlgTxFw7XcBEC5d4327caHj2q3PSK
ofbP6EjxymWZbzKC40plidz4jNvVB44nCDopALdYbtj5S6xCyYgLRKl27lB5/pKu
b6HyuJ52vIYOaRV67fpuigZUqPvKV6Uxs17F53D7YLGWSpUDAXtn56vZ1Z0uyqB7
hz37HGpNrz2bbarDLmuZUp1v1ZqcEjZRZIvDvFRWwXOdz90Q5aI/vgSZpKbhuWJN
latRLRTbIAko8DmBncr6Hr7yxI3H4WkVdfc+DgdCMk7n16fLUYw9u+pipkedQGGb
LeopvvzbFpSjatEVAsASA1591bMyDVJHekHxSjjU2fbtuz+NIYtWX0swEoiTgRQc
RipXvd6GE7wbtVo3VqVGZg2eGI6bq6nLwKvfWtsntJqW1C8CNWcxymToSHknVhi1
/0bL0nmsLoUroM8D9t2DiFeK0M4ZuA6w8XNqww0xc+nxuD7qSUc0/O3oGUtXC1wS
wOX6u/UB7tvrvz3XOquGzYdjFFdTQHb6mX5VAb8TCVbkCWc4vDXeBQStVolMPfx5
nvz5GbZ+bpkiuM2THLW47uxFXC9k92NXyCRTHsrWUAX0aoTMXF1DalRJVca0frdl
HP5jzey95LRz2ximWAWjFDmHIWXFa/zDvUC+qDf6awXWke7VE1CWLHkMk8fzeA6r
3VXPYfPo8mkfQBNVVgH1EB/LhObV8/lCKaRiiutlrt68GawTIoLZMN8fT0au9HZE
cKg45MVoY1jeQUNDyy1Lih4z9YeK/iafRCuIZPnt3rhMlvfIuXc27LvgtjVSJEpN
GiOh1CUNDIuU9bwKwezoYKCqNRFsLRNKVpoYx82FFAEj5opKKXe8cgosYXUhb93n
0YxLchjishnNkoMnWCoJt2/FDQYCj8tXznBQe5Nsqk+T5FMM356uBOS5Z63x4t9o
6RO+WNc/g+IC+6xhuyFnJZcXvnECPDBDo0yN/xCM0ItGIN6SoVa4EHV6j0eIeF81
BY4m7UzRj445OwtakE5xZ6v/5IkxRnCKMzjbio1gs+733+FBHQIZgNCMlSiYpAoJ
aWZcc7Xf0ad2tP9n/ddybog4wqn4HtZJMq5B0GX+BNZd2SxN6FGQ8rFdyG8aIE8W
BMranUlo1V4IUgq3z+pRm4elr/jUQ5YxEq8rcKviVZfkx5PpEahnZvC68/4S5AZJ
+VWjyCvifEFLodOW053lGJy4n3klF3voTT37HHTmCf9PLOmLIX50fR9dgQ28ChhJ
LLID+gAnEgjpB5KTMSEz044j73kdpx9K9ALCL5QdwGrZAPLbtyDRioWSUv3Mx2EF
/eqP6aXgBwiBBrfW7K+B/qm6j7KgI8VUv+QKmh8i2PkfqxTzhGE/LNsmVWrCVSQo
A5BUJZxdnFuqB78MdTa9lnGfRcen97da6cOlkYlB+cV/g8zw6LnC9Y3CaHEZzPAK
raw/gGE4G3F60w/pLkUq3+ExwGZrAm8Gyb8CAanYx7p68kcGrXnV6fBHdz6Tyz7d
zzpAA2uvRdprR3HoqLlch5OKOvXnudxxTr3Qxku6mdkBVak1B3Z5KV0Tsjk0md53
hJGqmbkhZf3w+zoRAGEgr3TITJiD495VBnmzLp82wPJGwfu5jNthjEqVwcVda9fD
fKgbgedcVgweIZAVSk2LWFopTJ3hEGOvlmtm8APwBnfqczQwDpQmVW6N3gJAN05e
Xy49G6qZe70vbNiroEu6Kn206A1869YIpW2fl0mLl42Sv4uPWdCUzNoJZkE5Dw0T
/cZDSc22BzDhYCuE0DpHGg6FBG7xroNa0N7qJrB4sTcwGxblfnWbMDTNpoFnJiXH
Kprbhbrb1GsEJY5uxpEVwBYzrYcyipIgQzrGG/GDqBavlo8Y2ZvOLC9Hzai+zHJK
3fwfat4+TWpcBleg9MI1vm6sPdIKpEX+W1RYBkfYCu8nn8WgRbbhdFRVKywAvfcv
eS0Z6GyQ2r7nyjEULht3FsX8MQHrjX26GRKGzPY7qDK6M6OxDKNuDvUXEZJAVLCx
ZZkF9k5xpz0U5MFPj2+Cde9JZqTaMlq2/FEZZn5fl4L+0dpj+azGnuUMXj9JVbHn
5oroeTSpHhRqy80yPIXtA2vA1eNSNeiIToEfORm+sb7v9+NHjwDej8T0faRcf5GV
BZmUsa2+lYruvje8YE5JSx/PzKnwELs6blhmKVyqI4v5CDgpxyWKamwGp6w8S526
Ax11FP29Ur+rguj1eoOdQafCW8leG2NIcb+t2kRHfZ67okGJEsVEvqO4y/9iOq4W
o7kUdoVNRhiDUdIrqRuGiXhpbcn1pLfA1ZA5YpwcRhQE6BsC+fta8M4K+y24rtQt
pbsMhJ2uNUJ74OrjOPAhlqQuOtr3F0DN4JSvm0KAnk7N1aDYUcL6vNMNbEtVPQvI
QOMdGWuQQLtNSD+W+0vhmQHXP3Fp4ONTCXHG7BMVO4fPIBm8WasOZDJD54SdFPDo
OPs0sYuaMxixp25EeXoKaraVbMauICIdLr7RYgtPGYf6Ut4yTnnKyQOwENNMjh64
QjHHNzqQMyoMYnXKbLis3Em1dzI/ejUP64kEoWh6aq1GdcyFEPImkuoqUBHmX1dD
ZgXGBuyxfDbndASDg/EC41KhCHEL2IMnBIxyOdfNMGkO+FfoNZOMOj0bIkUKDvYb
vg75vErMXniCdCgCcg/xiLOFhX4fy0vWhDwM/SOrxNfDFfDsjRtp6H85Z8gq4c50
n8TmdDYKK1C6ruM4gtB5JiSLDEcT43cL3ISgrhLEYeq0F4kVr79SVSimg7T44JWr
ap0KNtB3Ha+FNZCxY0nGI1EBi9UgxJJ6vZCqXT3urp6nkO5Hr+60ZhspX2vA0ZwF
p4wH9IC89TvaIzbFCR/dCm6tXGsRbRxdPyCL+ehih60MwXgs3LYPDjoIDINFNbRf
GLJTmzv1DzuEqu7DxasyRaoye2kHCeZzWM1wM/mLmZJenbWA+4qHaIg+0aY3Cfas
NanMLKskSswa3QlYC9FtG3xwBu1BufkwgLoIKzUL+68lITvSJzlD+aqyeCmzZXMh
3YZ/PItof5VV68Dr0gAVJwrvFHgO11YW4HpDcJ/qV+q95lbQqrtjMKo/14mwWtzo
P/xCQsiw4Eyct3eah0L+s7w5+7pXsL0+QPj9pAjMpwVyy8aSvsENbdYAQi7ocdQF
u8pLKJB1Fr7dLJ9Cs/msvUp3Pd8PC+6+9JJ3YWSL7X6v+W4aEs7r2fwq+Dw3MXGr
poe2uOZAz8z58dfB3ZCQRj7fUmhW//TveVYHUhEyaPnolcofT5ZsHn1098hHAQkq
d3cjQi2rOH395l1ih/xyWJM4/eWvN4CCXwJdrUjPWphQv/V9l66iBbeNnuZgfg2f
wrZ+0R7K9J5Hn2a4+ILVH9GF3wNLbWvfKIVOGDihBZyqbsM0unZFmBBhI4fdCi05
TFhWmGJe67JCHlZB5c/F+A==
`protect END_PROTECTED
