`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wfiv/4HXg0cJQVtNOcWMD4zILkMBjbic9vxSOsB/M+LF9M+tZqM6e7QLKgbp7u44
ppl8gX0zLK4yDWq5LPERehgAloznL0VEhdhE243Tuf0h6acFJa7nL8dTyQGxrMK2
kRrGdmTxEYIQW+7So/6Lde+sGW2siUu5b8lMC15Y+SiIYWb+sP2h2XlnxZIjW7T1
TRfTMQFG5qoFhzJfSqKlp8/lJhRRkN1ayoCSlruF4Hv+YTjw1YBUrA9RJxIiOoA0
1+1BnOzH6cIUsxzqcjQLEJaVDPxZiQ81yGEDsl4A6rv77feEHE/TJULj0h3i9TpQ
6ntR3xCzXY+CJVQnHafIRBRB7jlP3dHMVXyZllmygKZvubg7p+TXcfeZsmiTr5jf
m+eD3Iqx6miMKQtjPQbK/JRFi5n8Kuye0dPZlV/tu7OGrdegcFpxg80kI71wBobU
kgU2lN6UJ+NX48grkIZ8/tY/OzB2vg34Qv5yxm7MksBYF2lOcUbbaaKr19LJIugM
Xrh6MMBtzH+hYs+hCgPZAmZ6hMEsEBklLxQCtZn3kw/P5ywDFEHtkUvKQvZYrZfD
wZbwtFCEe9mOHh1FEQeCW2nFheDqcfqXHj3u/eFKkgJVZni78l3i+RI9oM53R1a2
gvj2vbfjJzuHzY6lc81YknNh839jJZdIrwqz8xhQjdv6cogN0hJIt5vhpD4Y3KXx
8tVRx2CKcY8jUv2nc3mmi3/wlRMu/WqCmRIR/Hkok7uqSH+OK+IAi5106qwJ/d0f
rgB1Rhq9lQRjfzs+rZjRYtyt7+gw9r4LVclMsJzeo5MSnfSDl6aqhVWIAGhNjc9l
rY4S2907cBzINZ9eEYDuug==
`protect END_PROTECTED
