`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CT8NsPDAtNkjIAQhLQs+mTKvUcov5wRpflwNkLckPnbYxm/YkKQ6Xf6JMqZ2Es/l
Zb4lWFeD65yf5lQlxLxQgvUoWswOJ9+41p5b9K9T91KxMka7c6fITDgYyB1Fx/k8
WsCpBgYmrhghOrD+PJK5TNOGeI7ni/vZJj6z9GZcsIOCMm06ZnPfimxxVTpF8cP4
rlet76BvMwI2T2cAk1lBXapEs4zdyjsOFuDSojlPF1EY6TsF7FPjmz8CTYhW3iJs
mkGNlXEJyarGlcxK6+CGdaXOAPrTOcUF/y81oDrJax74AOlbHt/u5/0HrUwZQ9yS
JW4P5jIkt9xjq+QS8AXUq0afP56GIEUS3enNQFdCS/LaHmZ3Bg+/ek6LOcax2lkT
VWefcKUY/1UuzqlxUio+yzWT5s/G9XoCbjrrSfDLrK014zOAbd/GMRBd8ToGaQDn
KsP0/HG8Oioo6qncsw4O4T9nG5vAPRsoy2TJs2Lz93kngPcYowyQpaqZ9fuFAJ98
Pm1UN4GdLLvsqWXz5LZIWT2XO1WnWjIDpUn6qVjKV4V63sR9x3ZmlCvT6qFM//ZF
lawfzH3TZfmg9krFUOshwtzdkmIgXUj9g5RLQ+Ns72amRcX6QraaUoCegyfxVEDv
B6jHvbv/S24f4WQEt/r8yZ/nzuf4+ZbzVVr68Tgj6H5NCf+Oa1foRjPmhBDgdvXh
n6IdCh30EYrllJ3oSBo2nHJxjpnmemoCUY02VGs5KP4ekT3og1a4Smd5Jmk9aeyJ
k7PFscrEXZgV23vN/hUy1qDDJjjJOADRgmuQV1gqwzrjiNzJgGf/lpmwajzWD1qJ
C9OasWCJcixASmjz2ZNwMPbR6+d+rxiAykVXhjk5at6/Sri763+sEp/q/3e2SXaI
bUQiqrsgAW58XEbYBVBfC/AmwGx2KlOGE7QBu+OA6RRBqFgN7OLL5Znl3S0u2HRQ
vtQJhbukB+vkO6Ddqek648kLBkSt9bltVyfKveDDQwLbGpVTYhQirJ/XpKMo+mPq
YCcS3WAEV0M0dDdhD+E/xjKQv8Y+sRbfp3BoQZVtTPtKdxQOVLjau15Km9mYgBzi
inGjNdeNwrwsq2yzCZS+8kcLibTzUn+aZOwO/dm4E0255aEUyTIMkNK4R5er4obm
G9GAaBPZ+fCWE4jyfhTSIdtqEBud1qUEZTAFGN6BFVMOBJTL9aEtKttmuOMc+byH
+jusCZxA5W+pPu9FkswRFjJKBcIFbl8m/wLg5/am18kRLQYCnkPF+6Bixxgdcdmr
Qr923j+nd+ocm4ZvJy50jMa8nVamGlTyfkH0IIbEQpJVnI10/7KlTbTg2skcykYz
c7oatbJU/C6jIDsvT0jjolg+IX1n2rlWyNj/bMR5rmcN9wZsL2sdFSLJcxQJ93Sv
nCrLhQh8WqzHY10hE9mBlYCKbPukW5focPNXAHH//upTjZn66dcw2/mBaaJTZm9O
8Nqq94/nAkEiJDd1d6ym6epCEIcCBeCcjpjtffZxgg8axzJzwUtNNCn3HdnhVmSd
0EHt7A0CJJg0ZfM/rrH9zeNiuHKa3FztgI20i1SCQqdUrFvlNXzoIA4OdmiomACs
KnjhnBiG3Qy8hPso6/ToJ0e6DUd3XUPAYNXfmHw0ciXMggvQfCNn7a2Chbh4JTPS
QVNuehajDIF6a/6BEvrn+38mKxI5yb3H0cyF+mX+dX3j0jSkHAU2y7J9GiiAGb66
OZr9HEie4yaxmWKXTWYhNKVYbAMcAFPwvwnePQOq8kEULDDIqUZmO4P9dfExXgsN
LoR61rJJil74eY9tYH16z3q1k8zUarQFc1eEG2ZDxJI=
`protect END_PROTECTED
