`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u6530lnFTWuLijXgRS6FwYj9mL2YxeMl5QuGWZup9z3WbPt3TIxhvfNlLeQXVJ/t
wPwUC/xh63pESf9RdVil9mIrruU5KXACaTBK0EPplNMR+0/eBmO+bAQkvsKYCW9A
Chz3YHltaYGAEb0wFv+1IEUWR84Ne4pEqzmrFJSTKPWP2ESqK3hIboljZCsKf/vI
jIM4NDPm3rW1bIpVg3GyVnFVKf+zWSHrM+4tn+3eMos0lPGSXwChM9NfTes4sJmL
cV8s1qwvw+6LUssKyaq4r26Hv6O2QG3EJbRF0MDRZ5ApjmLyLFX4HOsqTGigZ9mm
iaXmA6i2Zm9GanSTG3HztCi/T1DcQaoTHntoUy+XQ7pwJkg8o0tXMMc0xcuq9oN8
uvDNw6YdBXpQJHzv1LmYc1dfvVDNPZTOokIxDLrctk0hTKaSJVBkGTu1y7YWpt7I
SlF5tfmiNv4sICsuyCXxafYCMYEwWvcYLZlJibJBhUVhYUVMwr4a2UOsGPuNoszj
LRLBZ9rEhJNG9VVJDQr31mLKI3SbJi1UWRZNiVVV+gydp23FkXCQ5k8PE29jKtI9
vN0ekCCNjUgPWXHackfCN8wSXY+Kt8YH00AY0lAhmQYZCpPCMKIyXwTrvh0Xo8xT
MwlN9vRpjmZhfVFF1/+8oFYJP3LobRNjC6KXV3OfTo8aYY8FLHdmz9WHhMbEeVb0
bWEY7WYR57Zz946vn3WgI5B2bAOjDAmM/UHJNutoE+of34m9B54AhdKoOmjxgf7M
dR4/qvmdOUU4oDh5EAftNZozZCMZGsZExP3hyeldU2E6blKbb0gTagcbp9KsxXX3
SYeRtinwKzUX6n2B92dcL0yiWoG33o70SnN01f9SrAlCUWK/hNrLs650cwg4otFp
HdM0UE8oHtkVxA5qwx0K37KArOZVgC9EUimOB/5T7dy8I9TofLmMngR5GV9z+/0n
ZKMDG90TS4WEcKcjlX2Lww/t4uRRaqkbEalpbZMzSBV+r8moM7IO3yvSF2H7cKRL
RLwKBo+qwt3XwkGfEIBBia185zSKqMr6baidVqwo8dviLJskKaOCvqEX1jYbqSKK
h9ekAPH7L0WupyCnKtYclyK0HaGYiCq4fmL3IjrVdGxcvtBcpfbo0u/9RqUjm3eB
QtL0LeRkB4MqL6cA5YrR9KNmxTEFVIs42j6q3plbAD2+Vexy6tWvtn6Lgzo5q9bf
t1gaQ284VYtLLyb1M9clo7XH+AEnLSXalSZXjfVZakGIUA2IZN6nV1DZnC77/ZKy
xxNOlaKt/Y0dooyhIAHTtwpPEXSpaJLV3c383g/jKJaHdIk/+w5Klkka+VQx5SJG
MEgtQxKy6iGuImCOLBa1YsHedidWbkAiZS/zFwUN3y3Uf31ezrNxrdEuAFFxCbbA
y+R5ZfQga17VvUJU3hFrcWwsYBojm1SQHG+yhgoxGdpOPXzOIWLgkUutK8n9saon
XqOJU2VXjVk/b+a6+VdQylk679P56esXlr+QYR/+3tR1ajzix36mURrDrsOhlonU
KyTamSVs90XZ2dWLzHzRpkHTEeljpWFEUU5Zi0bJMzZsfcvialtCyOOK1oga2a03
3Ixp77FbQ7jTvrjfY6iAdQlhEjFWWAGreVhcel/ZhhptNC1FtdKcc5K4ysXl/gZF
40UJF8enHy07A5Ao/uSF1KZU79AbCs4jm+U77SDv9fJ2ja384PV26JF9OXtounmD
lH72exFgwru/whW77xR63YD5VnS+6kK6QLg8JceThgOOxGI6owHS98ptefhGPAsd
9sptUB0b5g+adEWD9E24N8R7KsnwXc0dN80PN/dsmIBIk7n12OSgwggTKd1GD1NC
K5MXZWK1H1wArPVF3syWZB7+Jtq8+dl6ezBvWNhGWCQSYtELYNz3oaS8NN6BpPYs
t3aOaCb004CFXUVMKfIW/7mZp16vM81wqg/P6FPpShqZe4IDawiNoIrBugcxlKLO
bULgg3QedGM1Q9kX0pZxOLhnFLMARzPQnrfSwqpS8ICJMiXDEvoAAOnfLJyL8AN0
1Tu0EFMREFFta2Rs+/Xmk+NT5V8Uj8h0hsrjTnmYj+OricXqnSbVAkFLCDTmNE/R
A0OCZ5jNQGSYjvLgKyl1FXregL3UdU2w5G7kPod8c0mfMHKITN0mbyigweFCbneA
+PE0krK9ZpLQOGhqtvfBQTTtbP/GmlTPxi+WPhrZ+LBWk4WpvijJNtgSwIDqGOU4
bGEL9sSr1D8eI9i6+kktH9l3DOALmqgDatrrHtR/Azn8fdKNW6n8D9CHK+htFDBH
gSbZJSL9cr443d87+kL8AH63e9XDDX8LnjkRFHmWA4O+TTxUrjySDg64+EniVVfD
Zr2bQgq90UBkwstDG8h1NkizEJjel2+x6xqYMSG8i9UPmaVFIteMof1nlxH1eOsL
4bhE8t4zlwRLQap69bzLrn4r+I1bAmuCmbILRvqIo+Jr2RB6xXUlq48xqZ4+7PPP
mCySHlpqyjeS3mRb/LFTWNCIix72dqtG61+v8XS0/ouLaJMpOixlM8hibIuDsZqK
CVGrqd/AJHCw9Y0dvuasMt+1vxXswMIvIkGgj2rZrB+V/oiiTKWDuiALGpOjTAmI
1IKldmMeypfsZkpKhVa2lGYHJD1yMS3SjQJK6Uvw7dO0dXCmdub34ik/tnnTtrLa
EMzHFBxRIxaljK1CCQxrmRObrz7sB/JzJ6UOopS1Ozr3ljzBRUx5V4BmEOELQvPq
Jhw81dwGV5LzyZxSbLwSZ1DwTBT2/zfg7j/1R2OQW8lSxp8+v8nMDyYSHvYCPLYM
9XL16SufgGdvPZZZZEWBanm8TKLnmzAN1+IKyNfdYp5BlffzQgny8cAzKLILTpu5
A/RhE25/xKaEttWCVtePkFR0abCw7Ijg085NuTG0+u/YlyaoPKh0165fq8hu5xoD
EQR10nk9V5rP0eCXQOPYuokLYB8DLD96tysofMy3/EyD+u+6qLcoynP933uw9BLJ
kTtSyeivtA/7nFfmNN391ldU8tHINh1o+duUPwzxNGR/fMSVvE/9tD2ftC+pvRdy
L6ftF4jVvHK3ZOLYT8E9bVVUfDV1VdaU6l5dsvmX0Nlw8zhIfDGm0oSIjAdmFvKe
O3PA8//43e0qCJ6nbwSj060/ZATrm6sU67YEziYggQVqiCrx98d9MiK6dx0ubgzs
V/BAvtEfqCUkW6Zg4yim+xYqPUB4A0McSYI845770NyBYLJPOqOUyVeR97xbE57m
vJXNL911tfLJKKpSHaR3OfojEhxt9o1gpq6JibbYsdzZ/EzdSLN1IJktcbIM/zCc
8RCSLq1NNWNvsNy4iya7webGLg2CYJWG5CC9oGWjBTuNZh9AIkIhaduQO3fbSs9X
Pesoe2T76lB9zgEPYTU1bJcSqD5RTIgY7+PC0YAd+YPTHg9y2gaGoB1CPDj+yIlY
JL+j59QgLmbdcJfIq6fr+b+CmSOe8lEUTb4nz3UVmuKjPrHCBW+SIW3CIOilawSV
ZB1TmU2J0COTv67GFR8v7hWHnl/91nQVghO/kjf3433jN5cMvc7ievYTB85AKC7W
XlSdRBW1ODmC558cDSNV2KAV4SG7ebDE/kRRHDIg9baexA8LtITtQc5FM4ILtu+E
5tCcplRaOlVAsJEpmOfzbpKFuybQcMdDoQCcNvOA6xrV0bLwOO/zFuc1mCEffsam
VrAYa6PgtmVlL13DbZ0pOW65QsZUyBkcim2G+iuyQ+VrPgHYD7tTAuViQeF3Q12k
mJ1PWxkE/JxKeb7A3PA5lJbz6qpN7AS0jGZrxt5dmfosHGyNeQkB9gx9ss6vkYuc
llIgcYSkQHwfoV/TNdpDHgNAogP88twkn01LJq1Hz7iudADvMxHI012PPfYPKSDr
gD7PCYsRANvekyQetgAhm2+gds1T8iO/aH2eexCE/slEi59JtmoFqMuMybSrEqAh
LLs1/uVl5QwwP6qAIgnqrQXz8BSA4FbD/U/QKETK1BDj785sDHZ4OAvQth6Fwv0h
An3FB4pxB63sgsMBkbatUs2/N66lAQvteuIG2egC8+0E6eMS/luS8CY/sl5KYBkE
XjyvpqXbVWoRbEmM2jq2hseRorax+S0L23EJe69n1PN76IaEISPuu68kb16CcRZC
+Cur7B80gTZQ2N5f+N/+M0KJ8M+fB2puqF2WLHKIVrsFRmByQGMoMpSQ7bHsjLCA
/VwYXw2oyZ62UBgtcOg4ZkAmUVLXvQIocKwfH8yTsEmNpLXQvNVyoB0ypjiyk00K
/IpZEh6B969AK/s9YzeA0rGrnqruo+OUdJVYMHf62hNLDFTUhQyk/50feKQ6ACXj
2lXlPyi+fh5MB0iBwhd4KecfItpIeeJcjZCQ3ljMTZGMEeQ8c7ZP2aaIr1uAkvVl
/YHppj4M4F+pgxxEHdJqjMjWpeNIhTNKJXGaIFLFtLAN/6jVNysBrcNuxurpgIHt
N0qzxGw+jO6yho+ijqOj9yM/4Rsb1fZEzQMyYOVrXA6Jl7s7GVc1mMkHblyQgBAq
6BHyhr0eJczHz+nGXRSqzTEGvIDcO4NqFLBewN1pbBedM7strPRF7z9EcYeAbmyt
gdm3IhdrbRVIPe5RNzY0b6Yo+IN4aowGb5kqgqirB6ksmaMW7KGnsx0R6pEPf2Ma
tUrgrhgZEA8elGZVAhbUln6kggZFy1zL4pfE/CBxAE9qt2wnjq0BO3MVST8w6KSX
aodY71Cfqe1AXcxTGME/WzKHR77YxxI1nK1hq7MJ6N2j57omlIRoLQ26JmiOV8EC
9jJIxwRxxUKhobtjFoSRj8VHq+cF3gZk46IbtGVTy9JXoGurmDodEuLUNN4mxq2C
J/7ZTXA+Tnthrd+nt/futin65SwhRx/+3fjEShCIYwqGo7bg0jD/i2NOmfR08apE
OUgzF+E5fdltEgA6L0ncVXexOqwbzYm06SB1yPztzYt5HucsiC5QpueIQwlmd59d
r+9hkytpnIhOgSAzuxwFOBY0FkULkZHYTuWC0HOA3xEBLTTKOkSaPp3uog3DO/oF
NQIiZEbIPGnSrGUt+9izZpBOTKPnctJSFxJtXK3nGfLdA3JYGjDVzM9SKbfTwisS
51+PHptc+a0WEcvuj6HTASNadiHwzzSU3vUdxTmPfcCnmhFBdIn5jbW8rv2rWRWN
m96cIySR83JktiNl+jKH3IMgxXFG/U0eRX76hMNiAkvRz+yc116GLGDw4iTibj1e
ZM6IYfbgVKXXWL3dQmYEMs+0sscmkfSd9v+IcV8mDXzfdajqCb18IO0QD5YIXjvz
rBo0EXkUKwpg8HwMGOPqJENqO8SH7FGsIUqu+lL3gWN4xt040mJeJ12HU7ROnyd9
i//dYvhWn+h9Xsj90QkILf5ArTYDRWu/Q0LeHBDmFL51tIu2VC2rWf/16jfQNRXR
FOyPNVE1epgs9L9HyTH1LajA7BToozLVCwMShfVUQw5s5SAiUmH5qx9raTxRCGbS
MF9oGrgvpyzJNJk+z2F1EyjlNr9WNoLBIvBftB3jhG/P8f4l1M6qLGQ3lOiLkJxn
e5426q20fUxMSyg5pEwrqCLvcUJr+JHqOziYSNv/QZDa3FjzJNAfMqgfL0PzOngH
zQKCxqqU9CQz/Ko6aHsMDjicKkavOJC3WOk4kvTkNjMEy8x1IkcDl1VUjam4qQ9b
vkiNUbJ1PZBGl77HiHzxqsJo0QY5E8hx3WoUCd234w3sqy/PvxzgrUiGiDKUbq6V
Dz99yNDNMhRJscw7aCizD6uHLB7NJxnr9/d+XT/7lfUm5p8VjCQaJjYbjDhv9slG
C1eC6icLZ2yhy05VhiZrKiBljbVE7QzeyETE56ctv5xaP7xw4LQGds2wf8FigDJQ
9gQu56XDUoNc1OR80DioykTwAp39j7JU7y9oKSLb75PWxkkiQNVDY2PNmElbQbKT
ZXH1AufPNVgyxGGd4nuyPTIggjPSFedk13df17MyIyBBsHIcHdSI3It7aS6CUfzO
qHhRwtGUvfgIXLbaY0dssZuMO3EBL14De1Wn63JDxTa4y0aqahm/9mzdAIS5PLJk
oxQt8Ndws6PhZzN7Rc0BLlgi0rE0EdVLeR60iBn6HaSqzuJUOPvO5OAatKMar3U3
5n13tHaYIFXHdBhh2SMQAFIUBdhyCy0B3DcCxxf80Q9e6IUDI+BXmkviTHKlH7vi
4arI2QkA9dXy6Uc3rpu4vIQJBx7mvpDzvVfum/NMDQ812Cj2IEal5sN8FqykpA0P
2N8sUwcEbn+FLvSRa6/zQvycQXXbSMvHc7NS2IaMKlRlbkOipkOeph99qEw66i/6
ZN6ylnaNY+hv4j6Zxv+12TamfrQFND1vSVyr5ycVgk3BDKC7G8wH4KzjDEz3X8UY
MdYkgZ0vqwMOjBaUl8N8wAolOK1eDX1UIzviJS3iU/PI8WzZ7AxIYyTmlEITryeL
Zsw2NSGomkoAEEr9hyV+z4kyBg284hcEijMpMUe1q4DGCr/U66XlIDl/Hxl45GP/
raFzOanfsHm0KaktWWxNwYX6ph+/zmcXm1qR78VXmtxMlnw/DdHc4etoci0HiVnO
gRZTvt6v2TRI8oUNxGGIp0uaMDjX6+cFGUr3ivS/4R8xVeCO0igmzlRCq02hJXNf
0kwHEnJpftIfQexUhtTcQ9ztKHek0eb1f7OKyul/RPMU7rjSt+WU865lcAJcX5vW
AoV7AHG2k6DsE8a4dHp9GNqg5k2U1RDlh6RYdeEHp3r8OKQAWAxKXJ5ntDPKubiY
UjWjkBn0ygsEw+tKEzAMszdMROXQZ168sCgPfu3yuhLTMWrI8BYQbSu2z08Gx1+s
bZmw+y3szZcwgHIPoaG+JEqI4BiomMwPiYolT3nw6bLdmvDL1AP9yA4/8VbVedvX
A3wWEs11N9zcdTJkOEfNREaNGpqRZIi7cg9+8bDpsVeYlZS7X3bFK6YXokFTj6bY
uBWIPh+A/jz17XQIbAY8FEYVJwynHcxF5fdzFvdCD5HKRNwwPCGXrZz1EG0QfbcR
ICnSSAQwndW+jMenL91AtRXphzZDBvylq3pt7CA1YsRvAJYhWHf8c6+iEZkth85g
EzNoOOyKNmYgiGZUxdDgUEz2oZ1evT9z+QtW+m4DVPvwboffw/MXpdkwIuImD60Y
nZEdiRy7iI/FDGaAgjNZp6HaJJSHS+OxIUwA4gmuJ07gu/f4vq3qLp0c8N+I0Org
A3LCByZ9h3o+m59SSCdyElrpml9nSsohgYXyp4eEUV+ZdmFLO9VpG8fnZKTkI/Q2
/OccLUHFdb7n240r8b1dpbabKLcb9HZ1mSUekWXlRyKCymjIdeMLmSv+ls7v+WjR
4fQCkhnSY1XQQaBTU2Yz3NOZU76pIvXEuPobr3IK4jejWtOnS8oqZgVmihXr4iDe
VJ8oxVNXXmdo+zH7gQiHQmAJDF/zgd+BESXs4ynMpIYxlsVCDp26qUufQCXQjHc3
iN5pJ22juWivzVnCdS/FK6tpv8iOoeGal1GcXe6O9dP6hhEY4aftuNWYi09+bdBi
S3X/sEto8yv0cWlQi2BDnxY4koWmjW1CLG2cw/Wymt+Stbd7JYSzUM8lUSU7L7vr
lABl3al04B6WrHZauVQ77MoNlOb8jKQ+TszkH44468bdAXpjVKbRGNJKOOKLHhnt
86HO/8e7gm913Bu2a90loQaxDXo9fHUmsKMAlAS0U29drFaq7N+IhWeUnG0eNhIq
LY6Jk78ADr4VN64N4EnpAYVA3XbMrL1Y4XgH4L96UDJBtYxHW2Eh4JxnfK/cmwKQ
0yzci5gBESGpG+3TYoxgnn0lIPp8RjpKyZ6/TYr+GK2/NLgnfd8DrWybDiGM1MXR
nZlxyj0CSGTHAwVDpj+zohfilb6wkDpHDv3jAhzTGePmDcj1q/UDQIo7I4Kr2Mp+
B7CTwhs54Rhi6RM0rQt8mfNMk8+j/Qdj+BNAhoouZlLajHH4Oqq9sas2EV42lxY3
FzfESMgEdkjN5swAplXtYPu/TG/gJJsZk63xl+VAjZeU/P8jmbeUPYucdNLQyVbb
v/balRT+vxBYDLEp04d0DU4tJKofTy7o2gHgH6dH2q7T3PHoUCdoE+EHNfRm8AXJ
4tG/Lwa+fWNyOz9CM9rqRc5seDwjFff0tlAs8jwhRmvF7YmG2skTN42mv0XqHE8u
HV77QBVzmucop1aOE0B1fYmOiFeoRwROid5k86OuW7N2XFGfheTwRiljf/XM4G0F
drPP1I2CuFFRY9HMs/nITx/R9jrAFLqdMPjphny1ctt4J9ETJuprFPAWIVl9bFqs
x6tjFBX1iH8Y1/ifWAMEWAkDVOxlOceyqCRw62wCV49/VH6D1rUSmhNbiGQCu/Jb
+CU4EC3zwzXbk4cxeIWdNRu69bx0eGV7CJQilsTa/AI29BUieE3Zh121w+0+cn+M
843J3td9pFTA2rPnej/hAwCi/MZ+kt2cIWfuKGuXmCZ6azfbaZinXYz8m6tu813c
6qIZ5ciacotvJLZjBTUQmxmyVqjcp+QYHuK8JL+ybsykOJaY/VVEVqefGC4s/pcU
MwzXC6YBKGrkdfNjtHg1wtOfGTrYQuVz13N0bP9RkBp6h+sZK5lXKxtDsNkMO34l
6szlk3ZSrjV00lyOqoeIy2zRjU/KOtI5g6GYRs/ii5n1M1ma2q4rsI7Oph3sVesr
vWjFt2LuscRRYJUC1f2+YXIxVyLUmuL0RL2H5tqvT/jDBSLqnpZDWUUI2II/NbeP
gwcqOg8IWLrmn1vmd0gQRGGqLzRlFR9xPxxrxxBHmdeVwOJMDQ+8Ai24EyPoMRF3
Mffgh/DwV3x+jWGoT+4BdfSOaTxG1oyGcfIkrzHJBcJDavpG1feeNt9liOdLkDT0
CyjTPzpao4CC1fqNtt1J6PezxmHUw3y699hm+EoIhlupHTAME8qRfe1arsxv8/Nx
oj2y3lhSWWG+YIp/9Se8xxNUBDu+TWAX6fFxFcuYqQlV8sINyscpR3sKxbq29nXb
1jpB37oQD3jIysm6wBXN57WYDPXrZ+3EmHE4MzG5d0aas7c836wnOjGZWVbnhtEK
W8S8onu+CI5LjkLyAxhWy5cWw8CokFVV2uPumSyOcp8=
`protect END_PROTECTED
