`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DKAAxBlula8I5inmFhh0+0WmTMr+Y/wieKcaH/vUsdUx45p0xrCpIcDqTF9l73Xv
J5YR8pgjjcwQzY2rf45X2hBBS87+Bi1D9HaY+4NabFNys3kDy7NdKNeACIYY4u83
aJxQl43RDMfwnpppZLiS02wzjhSiiQjy6gE77IFAFNjbcJef6BUQkGeg46R6rrvP
yGJkaodqvVCIAaOrC2CgpgbFTUhnNPElloJzgnZRclC4dXfoSeKPovZXujG1GjVq
GDm3DNBvVt9CpH0joL4DpOEcuyf2E/4fCHXruAgGTSV54NFbJbqNQvrhmwYCSKmR
uYKwCzwqNxMhGJqFNWHVp/zsKfiU/oA2MefRWCeer6KLhUEm5yQslbutvlZnx1uH
ymlsByjll8GTc1ZyRM5mvZC7B8x7SH6TcqU6NmaSyKtJTNv1LiUt48q9p5jaKMvH
fBqJ+IWm/iwbkaOvlb6/J5+g77nLO6gv3dUzxMXMkHTK9VWacAbSOnD1N/dGjO2z
0uiQWZ4oyLEEYiPOmHtKu3qZkhJwHiybeknQCSaioGbXEPCk+X2oAxwZYDhvY5XZ
xXQAs09MJbNce9TUKfaY4Krc91+lF0TAIZEzJ+BdaMiNnLX94xDuvQa9PIZMIpA/
`protect END_PROTECTED
