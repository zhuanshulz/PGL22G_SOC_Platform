`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kmMNgDi3PFJKQpPUIMQQv4ghp2/4xP44LT5Bh1+Av1IEd++zd5VT0XpadMwqRNA7
lqMAZ4BRItggvCWEGfx5Yg8IPH4Sl1GxMt6DCGtKhNCFu39mIdsCyEmiUJL3rTcO
xLVF3Jhl3LnnQFMXaKi4Mfw3PozU/jIwhQMjSAYsjHaE3SIVJJsdZXc9kX+A3z30
+AJb3d8EaMcI8LVozhaVbY4HtXYZNK5E7fw/sR4TbYjbAYlCCr3EDNWT8JMi9WSY
mzDBM6vve5fAVPJ5aIgPpxv+2ZpvqiiUynPX4ssZEiiKmnKkEDl8pPe/bMJvIVVL
tWasAkCipev98NEuEGT+i6qhdTIDADBOKTav8aOH1FIaSRhEXer4SBGuWPRAVoZT
vDCIGOsFy5V2F9oTI4E9OtPE27NnkzLUyPsQIvsZYcpI+ate4XNRwpG0eNmyBblc
TgJNPO3OpYLIGT1HOYrjBZKQHHzuidS6BQugOfMZbFOf1Wm2U3Xitp2BLBVt1QgZ
`protect END_PROTECTED
