`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hy6M/keJF9AFkqymvLhrS9pRLaddtFIQeMUZAVskd3gk1uizOmXQSupi/W8+zkrJ
PHumzBhKQcnKLEnDuWP+KU6eIyOcisiBIpFo3uVfyKHIl9WODeY2asITXS/B2VHv
HZq6I2sk3WtBtIdZBoRURbhK4+uZxAIYL7Q0A6uVe9IvOISAN08B0nlF1LDSIkH4
T6Lt09d3PLo8SN7UHrslbOu5WHcrqPmnOGEoxRKz/BfdjkWF+5gOudx22F6iurMe
9f7d8iXwYtlkHysO37psw5KkrzFNtpMf0wi2/zi9lagH4xc1QqdxpY5FrxVIbqjl
atvngqmFag+nyLpx8vikbfvIabq8cAp364oEme4NFsTx2hI8wCW0eCUOKJEmQ4UQ
Ij9N9zyNg77ju7OIvjg9uD0TJ9XKMjXFP5Od+TDZrtqqOtEN1eLSYICVkCd2Xog9
E3+JN2Oq4WW+I9VB28dIKUYazaX8LOgrN+aPZAvLXT28VF3/tDRuTUCOnsKjvAar
+i+hwbU/CFpDec0IVWEiROUZyL+7NptGFwjTPbzcKisLHMkNZY18NzSJVcu37MEw
DXwcQDYm2mzEhoKWaDT0A07+gzAk19A6GWRoPUqOHH+2xlvTJFxlLsFrTKqHp3/f
ToyHsfhd9XG0uU/r6fBxynX9A7cBzSuUK06Lwe1iVpeCD4uaeDZCCXqxCxT8et/+
00u9MDtGeJe2tZALdAfZbAF6aTStKrSmRSJl07EBW5HOGLTfkHOmN8+7wW09qQS7
HRHHlCFnmrPla2/Ehq+DyP8fHXCIn953c/h0PIx6s1/QisHOy6v09U52QU0v1VoY
2uW7/IuchtiapnV7n8XHFsC2y2UMEhdfZH/i8rftEZXuLPIy5yrfWmd/TjBeMH7L
e+ctibn3EwRbSuGKrPgB6tdxPgF70OlupREKE0gBdtYeB8joIe4jqIn4BnoXthsl
5Tc/GsjLHY9cPeWvZqQE3D0mkj7XgayhUKDWsoNhoz/ZjzdH6Nb0/E3g/ScrXzdF
dzxIjo7tqnsXzOp2BcAl8cc16FidAwqZfbp8jTjE3IuU4Jct8gvmtLbSto1tqbo2
CjYx8fOXXFYV5UikVMr8sGdaBiMyiZKKLt0yDjj3A0Sf+Kl5xghL8+A27t8gyBEA
wctILH2mPlnEaPOb5x3Q3z6GyTk5hkzWBE+u9r2CqNkA+CFlblrkN9aDiJGGWn2Y
4WBqfgL7F3UYdLDafauBspNqj30AuEO9cgsb+5Ao7vVbZSmEcugsqIU+fliM5Clo
`protect END_PROTECTED
