`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3PkMrQBRT95P0G/sAA+eHeU/EqLSUyV2UoOOl/hGUHEKJ7Htp5LWx++f/hHR26pE
WMjrOfJwG3blVMyk5myt32Sd/FejTQTXTX/rklPHokRIrgKCBUBfGmaRTkRjqt19
Iq7vk6t1ZY149x/IWUeClaIxmfpa01nSHcQvFx/nctmvMtELbGIxkLpUKXMX/PQ7
A5RY6nw0GCQ1Rgv+c+jxUKCpZo3SKZzmrevpoWcmWynpfDr1+aw0PmxOE8BZtHX1
oCdhKUNNWl8tcbgm5Tzf9/Oo3DPJYYqRp/3JP07TRq9PEz/lmsAINuPZCeYftDY/
Pi6KWrnJdLGGmiQZEwmSG8V2/ZNJkxA/abS2NQEIWaOoZIjLfWPIYoBYvgXnvz+F
YCFV5HIYEJSvjC4ywha3Bu1QLPjXpgEb4oj+cx4LOOk=
`protect END_PROTECTED
