`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Br5Kq/UbM/52IznEXf3cglvDWwHAf/Pgk1plDcAZtQOiBg1csA4g91eHlrjvPdiW
ugRLZQSP/25qs71Zvt08QAQmBbpJWToIbxzzkv8SOvzOB+JaIK9Y/fw/pQHNGSR4
HO8oyDmi6heLg2Mv3mGpKimcJ8ti7D26jbFSQ6zDX7Xfa01na9i6BPrgbyxQHvVc
yok7KsoMZj+RaWNCw93x1MDg2MvRveVUZXjicRH3IItA+6nMAO/mZFqQB9O1rRBj
BA19+VZ9KkCqrKAMxwrg9vI5+YWuFnYkeK74CvI5os33RYrZP4/xbYm+1wuwGM2O
ee68KG1zJ7p95fSD2tiIHFbBGfUM94dkNOQezNt+d4BprsYrw8Xno6kRYtZIDdRj
E7k2z+sCHPzp4lZiK0XOkc/lfDgqjZyaqoJR1ZTyc0U9yG/M6742PY+sK4XOroAn
HnE/ORepLAgF1yBiL7YxqDiFApfa9P3FqtQdv4y/LLWmKNu8DBTFyGpioAM6emFV
s8HEasPhx4Pn95IEMmLN0A==
`protect END_PROTECTED
