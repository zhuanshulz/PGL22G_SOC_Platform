`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FoWDQV/VF7U/zuE5Qx54KoFkVFuII9whY6FfHDLbCyfOh6P+4EYm2nrUjLS2HL6o
42S7DJ785vAWONus43almhjng4rInGWeq7hOGs4sQqsIe2ai1bejnTgXGcowoN0h
KTLQJKcu5yap6wi6ApWeiaADHunTAY2/QUeYSCP/BVf7sFq0JiZomruPjO9U71Z7
5ijHOf1d819UDm5kmclKvrCHjjyagaLxdESMbvPEhz0WFhgfznRY5Bc1woTcFUPL
S9xrOWjyklk1xZbwVhHjjrx1MFM84kpcPbJqchhTeIaM6EaXDFEQpAIHuOtkPmm6
Rpv8nNzur1NXBIkIQfvn5D0VaqM0Req5A1cuIasMJy6IN121sMp4b+hWkQs/hBDk
HFo3/4kzsH43i8rlWbWsWzdgXgoS/WqwW0xa4kTgosrYzzlPJ3fc34NhDoysUe6I
Xc7kmJ+hcdl0pwK9qDTI3/XnJYSrTlnZB0nbHdRUFlyaIuvtR2RAh6Uwc4V6+rAY
e/bJAx9ZIibZ00w7txMvohPs4uHV8gd76yqqXK2FknFWvvtFyCIxgz29AGP/2xrv
/EyRtXVjFSWdGXeKBM3RvQ==
`protect END_PROTECTED
