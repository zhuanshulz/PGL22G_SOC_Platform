`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MDFNhOZCOjDML/Opmew41No4RWsli2nB8dHZwKMQIhMR0o1AHgh1ijN/DWnvJJvz
FBFNvDjDvUvAbxZknXwSqvCfN7zzpmgbQa1bXKn1QIVtXlLsubJ3LZ1QYle/C+Me
n5uGM7AMPaO9+Py6QpEMhotYEUgKZRJzOHeb7jSPqg6tv3zcDjusvKr7DDSZgQxV
yZG0zRUgvBon/S+3gXlY4/JELGnrGVZL7uktd8SEtFAy69aDOJLHFfP/G6xY9z58
9a7wSV064SRAf2rn+7onR1saxxv6eTxCuu/VqB0ddSqcaMBSQOl5ekfTESPVNS9m
izGaw/5iTzYGmQ4WGKSRvmaO8yIzrwAZWW9lwfjAWhP9/6jqQbpqJqqgWDJdGdxh
Wl1YWonLRZWGzDEKAE3tLA9RMVBZh3i7Kf9OtwpunKe0JzgNr9wauUDRobMN4avw
CeOLkNkExWV+v4niVRGfFg==
`protect END_PROTECTED
