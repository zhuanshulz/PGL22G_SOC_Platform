`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T4Pv1in9+luVWuZVODkqBebL6Nh4cqeRXIahnmprXbJglrrgsai8yviFY1Wj9b+N
Wit6D+NW+Y1XG9X9yC184kY7YqiPOxXWVWM2HolISf1D5FALomxDCniSXXBzzgXN
cPBB45332OiQLijAQ2LzA243UcB3lcuvnwJGvzk5DGUQ8fQU2m0NIOiQm8H6exrn
mEh9QK6/CGHbSe6gZP45IrKThva46Hxn6NaQXX+tSfP2Gcu0G1OGdeKbP5VMl77B
nHTFbz+DGn3JW5+oP/GXpg==
`protect END_PROTECTED
