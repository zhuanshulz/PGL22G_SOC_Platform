`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UnW1m7sEZ+JCPJaN9QOa7lKsCWscPqc/h/eRN2tIiJqvQJlfK6V+Mqi0hiC/kgAu
fXKU4EJh2vuLAq6tWtkZ97Hp7jk/n3gTv201lUYydHOYhMwX/Rczx06tL1dsrciG
gtKVv31os2g08BPy6u1dI+n/d5GnalZEkdmMSzDWWd5qJ6MgZU0kcruguvZnhG9i
NP5T/5cgAgmoRv7MgBCqXxL9TFrdqfpEwtmQxRJaiMQK0cfDKliHWocM/0/pFZEW
kBYFkBFTmPRazqZTUklEJDXraEeCSMuMxJdl4vcBe6cddOt6WH6gksHYcwKci7AF
ZyzXj+EyY8fnuQDwvTazWEl2tLKKsu62tS0ycAmrbu26eh7buM/4/eYL6Iz1FVoP
piILVsLXT53t6gqwRpEVNPfBe02hfmnEfsYDD9Bt8+ih6ITlVNAFgm++NRpTX0TD
dXBd4p1cdsFciBtxEX64XNC+dyr6F3REpZwbT9bDKBMK4S9RvrTrUYNqLTA7D46J
uPchdHTfs4FneIq81PDyQo4JEqlN/27INGgrwdmElTfLZ2CGlm2lkXkTQhsq7z5q
AMEr1R/VN6dE9Dy2ZtcLLRd8mSKtkWv9dZRO0sJzF/uf8nI7vC/3tOFliR9Hv+CE
bf6jt41Nlx2yQCaJGJeUMNA7A8+vp+5qRICGUDP12ZiAXHWmIwKHrs5K0iaxe4al
wUyMRYSXi5Zh8HnP+45tjC6JUzZhRspnwyGypv0HpKdGiKaEH5Ci7DTdWkbLE6cm
0Hac8wMAOjDVLD6Sbvkmh9308ofi4pL1gk7y1JDcLIjSiGrFjXKtrew1jD/cqvtz
ZjgMEcGofhyj5ZJE/0/V12xWlZ79wqdhUruBq4lM9H/kHWFwmLXLYaOypvc+Ojjj
5stYx5YSKcpZ7qahc6txnWpOd04s4XP6DAnwvbTlBM5EcjIw39/SU6TXW5scuLYU
y6iwbIQZzeh75boFoodN0+wU0Z1C8zOUHr48OQDlEbO/bPzfF27pJYuo35Z5Ps3Q
Gx1e/ypoXVsvAgQ5fcpYFFym6jcPF4zkwpIqRxBe4qla9la4KmboAQJIXMZgjLiW
EsnZeCnpRVvqGl+CGWqg8oIX/ealkGG7o66tOcMZhIC1gn+rSuXza2cQQEHILRPZ
jbi8s5eLAPkxa4j5/XVx5aKPreMdjNkH0YmaoilY+2zs+n/4aI6o0nwUjk2K+2XN
5JJk/00hDllsm6uLIN8QAja9fNL0ScBnV1Lf0XaZT3ePEmiQf6Zf+Lzu+nTpj5FO
ShDCDGB+jePpfCgXJNsYmTXBkjWVK/CY/h8Aw3I9b0meKbh+si7weIr1EB7/mxIz
E4xCvCE7WXGjHRWfIM3I9CMf2NNY1QnbpzdNI2cAlCrCl1IcLal3F8EfiRjnIOAS
aq/WnGaArWeSAQheqtOl71nRxXQIN0IfIIjvF74wCRGg1Sa/PGH0GJSmqMvsp9ZF
OUHS7/JQzNG9rcS77xF+yBkfXQosDHQSz5ihWYNP7N/wLRXA8U405L5LzPpl/Hmp
5YnQa3BMdQS1VL7ppz11Hyk/5251KniEpMfyBIOd/WdoogkJHdQXYN79rp9NYb6E
Gh3+DRzNW2fWSsq/b37PTTbm/r6TIgFa6JVRuZk5bo6Ou3d+Il0LiEt6+5mH6LJH
Jef+hm0PmouBlMpIQIJ1OA4IMcSYRmD1KQN+Ynim35ugG+19YQ6n58BkZ1GWIDby
vYrZak+w50btjQPRuOOIj6xZBqtVCC9dXfn4brNOa9qBfYMJiOyC3FK9KiDYzqFu
HnbvOqHTKjqdyzWjaPpBeM2FMPRBnLSKsCIvcexV3JgsUehFqDpyB+kxIBpPwZXk
iqnwRUywXR1d7+vsynOAcm7IRrmdKqxAT4rLKoStMnXmM51+1Cvl1bHgfWpvpu/g
6/ZH+CIYUOXIeUnfn7dIZcGd7Yh+D1+v0xWgRHK7qcSxJiOGpIdcTHliZure7dsP
v8Gla7a2zOEGvbAZiploSM7DJ1IvgZaO3RQpKyeVHOxwUSGzxpfwMROkekn6zFAN
EbUi9AIYeBw/sOMiU9CVqLCgApon9Wnd/uiSK3OsYxXJxzxeiU5T/uEqjoquDta4
G7Rcg+Pe2XJSAusp7oaDPq3IFuYxRr8PxHsYb0vX6E8YZIVkJH5TOVpV/DlKgf/2
YBXbjVX6+XeYC7aXkhUtFlQxjDt7E04FtGn9ygW1AGlpLy9knb2ZLDpBAGEiLRRH
ldOqps45I1WmuOYmzY/9e1vq46kji2VjnLu71X575UDx+l2D2qeOsPVv/aXzA6zy
BYqtbFydBZNgcjeQwly8CQ4YVxjWhysrBa2BZbNf+raIxHRikdwONr3JIV688uPM
8oryeWbBei74ekzq1F9AvpKbPnVPPeilKr4pJUn7z1mVfwIV23CDmTG/QZxGH6aV
SKQmlrZvT1Xv4o6ZzZEbS96oBiPmNGks6lw8zVl3P6KQQVUn5UZBUWlr7+vUeh2s
w9Qjdn7yuYU+/pB/F3qicpRK8AbKkF9us8S4dhFW0iDmtKHLyIPhVVExL6+x/6dJ
hwJhxKISSd2eKZ4S3zeBaX8eDZNrqi/qoJbIZPoITDOaOvWGvUnLDnt5TUMo9r3x
YvMjW4YHRxRltC5TlsIM8OSIdR00yIE9/cpECLaJ/tWh9CBofn0Lpvhh+fZVmt24
92HqxbLgwHwR3qdjIHyfLy+dmXKXZvrXOYBhKIzkAuU9+RBaukiJ9lVJDLd41w0a
DJSTjEa4GERSfMueH1UaXrNClGPE5nkrJCk4oex5GrH0nfiMMHa7uEZTccRL2BGm
xIwhyrnV/ujPM6FeCtyL/0fjtKg0gKiM5JieCZqeo/3ktH+Sx186VEIpoJg6e9zt
zVAmLDVq07c3H6czUid/a+WAHZ5UeNQTGF29mnVo+O1hI0V4NNBhJdnr8YHKv23m
3MKQylqEc5yyUJTgHCN4UnF23EnyxpykZPngt5h5kXYNpoaxH6o7yv9mGkV+ZEzu
JSIBt+q/YlDM75ttwtwncrs81+KVuElzZSEkAJopRP3qNPYhRlrEf2z5OTdY154N
SOH+tRfKvEXSsU0QZU86t74TzNrLasocf9LNqdT3abMEzzmk0uAEUvdKAsNXNn1t
bjLAHs1YahezaDnGcNP6bJ33wvbc0SlbS03/gm4DGRcq6MUxGjR5gBbX59WJ7mqj
0Ha5oW0qRp02Zzi46DxtModn0JRncpN1vNqjg48VHwjc1cSmfbczE94TANzCLp3K
h5MlQCP9CYV/FlZQ5lVwklFTaFxdGd+EvDiHnEFJuVNz/ZGxURRIF/x3Fc9mw3uT
ajKe+DxMznVgEgbLlDbfSlsi9otLbMgEWjuml46GR4JTVN/8cfOK7rvoEP28BQT8
Y15iLRwQZcMZmH+xcN7u92uTvHcAf+B/XpJjeer8PtaZrh/cTaXfW20PFnSG6Oaj
fJoD4S5N+x3NHGFqqE65AiP5HEdFtlrnbI7NJimlhrgaapcVQCMBsBZaZSa0tyoM
2ZBo9uleeffvJmruZrQYqBj9TTMJ9ElN1IrsBnJzKvOqNpTTn1YzjQSYWlr8WVho
wdTAYrukwPmVUSzoCa3raYHDqiVYI7w7vxQmpnH0Qa0x1+O9SBVc9GjuLvH0dP1V
ikvkYr245NnbPqCisJohVUDJuePIWPrMTD+1yu0lGpS4h83jekSy4CW7lQmi6Pal
fq8PSMSlvkejWXiE7YDSw3+rQTHg8kzjdomujF4/gLIIfdsFdM6pr1S+jHNbTEnO
FlmcZXEqizS1SeLnY+y5TZkdNGBYySkInpguyHT1S63XPavTct6dnmnWFP9B9LH6
FcHchAvpBDdM38dTA2yg7ZxXDSqNl9RahfkudwPJhAKJcU/dz/DYw/1Miij7fIBc
UB/X/hoZlO8VJVbSg93nFB+b6l43hdbKNn4VLYwQQB6jF6lAVrDP8Dvr8hapk+TS
z1K0NT+1Bf5lXSvvPyVOlVKYbD2SWW6kJa0UZX6Igo4a3TwrQvjUS/MEPba9GkL7
DcbW2WkdaYq2CXmRpXiZ4nDUwwEsB7CxRW8vl4iZ/GmYQQeDo8TBhDW+W6qdOioC
qn3yla+fBfU5BXOdyo4uqulEzjG5CJInsBCwAPqy6Y01+QeP3G9u9upkGHAF8c5N
RqD0uiViIQ0HHD0apnV2DRbQYCxeCiRmPkz0XMxztkRSvsGUZyxzNKWIr6ypY+En
T5o+VohZ8sFgnKvkLMeo/hrLqIaSPapkxTAnk9xzOB/2YLgwC+m6pQDS5hkxPUDY
GN+uXgrLie8KztPAcEc/HyNYHJDr0nABVrq5AQvc81w8h2eozz5jIU8fC7se8qIQ
lnWqzUP9bR4fTqaAKtC15GLQH3cwb03BONekb56jLDDXglQN5HQyw/eUGhH0r4cd
E3xmsICkqqsukYUeWnTA/Ler1TZ+T8Ym8dY9qH1aZs6SwAybe6R94TetqLzU/o3R
9yqagXTTYGr9aJKbt10J5qsCX45V9ICkr1pJGNu+3ro/FYcxm56P6xnzFAiSfxe5
jRGhcHIm/ltc82cY42mDDmrK5dLRM0cgdPAy6BOPO72YEHslVk1ycHqr22t7H4SP
RxneTKe6IW2303TXWgkALn66Nf3NJ8D3SkA0jdXTryMoJVrNu52n0HO9Haio46y9
hFW/wQWTqq2czx2rNkDx5gzljS/1IBFWshHs4BXWPIfDSVg+e+NKdHfbxrtQONQC
5yfnw6L69WsynzHmsGa9Pak19Q/MaZpOB4EEeQAVKCm3Dh4DLXmlA2715fgyXK4z
Sw5se0mpsStdidzHuMJioLQmg9HBa07dYORn3NeD8o3Y6r6sRnQvRYrs9sRh5bAE
LieiXP/PlxjeU7Vzsnywj6dek+spWHZcoTjIHN+NXCXetjNnT75TpkKuacDhRu0x
ce47V8UvRwWmvczluMLa8CPeTu/Dib6eTHsjP9z5o9EfMZGwUPiTWI53WpXTazaO
S2LwafDq6GhWt0lI8ruCyqyW0AiBJK6EmiTZqRfTDaLxSIf/gDguGt8RvHCurwWf
xU96kNQVw1s23etiWgbs4BEOqn6SBrX6CleTn74yi6KXWyeJytDrC/fHuWHH0LSp
ibqf87u/h16ZTq2LMh7JKjydwTMH0kFJqHl0h6xYKs9vEy1YN7QTcMfLgo/EScdK
AGGxy4tg6i9rXFszzNrdW1iKrM7r2QKCVzqv6KULTsutuIhhRAxQnJ3MNleAeM4J
I3xAT44jAwW/Qa67BZJ+UuT1eJr7ji9SnTbeJGeZnZoOx0ySL5gB06P40dlI8VrJ
IPpevdKivePmAP9B7zctWBJw0b868a17wnu3Plni8nDtKF5aUiym0pj0ySbEsKlV
Owz/MztiTWgePxAxE6gH1z3Mrdovp1GsJibpvzgECmD2O8lqMrDirEfrC1QqGx+4
3l6o7TChVeHHLzca7WgbuKNCNgp55iXGLnRssFLWWtous8FgGv8XjzDh//gFKa9b
Attqz6fUXDRS1wJs4FlYl33/dWVrBIMPLmKGXOItQV1te7iBoPaXIDWO/x5LIVW/
XpiDloPvIk82Mf+RKBUp4Ie3jidDLcGoqILmZAFkRxV3JkFxR/v5QLhNsXbiaDPg
LvDyDhM3RN9OT3oVoagQmAkNBahubnpLHKyuWg3kaKQl+Gnqm72j4A1YJPue1UsE
lQ/Vyxp9mLynPOI/+n0FDhqktovFAhyHEoxTpMkOd00fsjRqDPoDrVGt3MGhHNMe
j86AX6Twp3enQ+q9ldOyYEHQy56rEHyBdtQwc0yUImYC/mfBA2wKMuldCJBguoca
Qt9LLmk+pWrIa6bljYyNEnlijafz7STT5KpjBin/lWt9TYsq5ddt3zQAU+AVHyxK
lQsVP/630l4z3l39Didbuoc0GcW1XrRx0giwZLLKLIlUR0F6vWzqOHc4jJYxEd5y
oEuyTLZmQAYT1rETifcdeQljtaRulJX7W+IbkT9dfjUQn4urO6itYWA2zV5rC6TK
vECEz2GYQsekP3Jijrz6f0AVEZO8krUW3QtcCT/O8Zi2SChaxg1CC18yKgAWxVpI
oOhbBkwPPTLsshxwQGXliin575O5AizT+sVCjXrOS0qhYRE5NYxhV7D/Z2gaLvbW
zT5wJlKuzhj/IgEM5xr3p4P9HapJyMSGbHdPW3NM8cwWaDFpcVhPI9e94sTsRZ2F
Gnhkb1i85Y4wA51qB7ip0HZYcJg1fa5+INUIBeBpk2Grbl1DhabT7LALnqln6lV+
SlTOordkv+JYW39FH1fWNCt9HSNgX2M9x1OLnrqu+nu3m/9SvoEwD5FHpvcCfPTd
mSDEQBYDTaJWLZ/5L5hn0DL/+XIAGwUvXg3V8uWkAxxMFed8NTU+J4Zyv/YvzTbk
mi6KYCaTaPHr875wh/8VjAMwXBPL+FMNBesXpFIrYQKYtkDEq2FrAEWZGCWOIgv9
VbueCAJw5isp/AA/MlIMV4cYo/HHCg0wWQpp7j1jyFdVR1d31vZ6EfM/fk3sYngJ
p54UIUHTRGbgMNrz5GOhUuyPkuLAHTt+x5F+5/Xg8X9dlNH8mEGhhtEk5hbGYfs9
rs2LIOoe5VSZw+KeRIm3kEVtin3PyGK+RubmQXTN5IK1IYsS3KgwnIdKrzzwQXz1
RIIrOrIe9O0nwwLKgMtfB0ng+YB3XkIoqAR7sO+n73UTn2pHIHrQ388f7PlHbbaz
bZsD1Z1IoqSseIHFttwiz7H+maoGKJYFkim123UKf6qxD6lbvgn+7q7zZuhx8nU2
xuD7SNF3aSjwzNcutYE9FW+m8u3pPJ3lIY4ESZLX7SogoYZlj68VZV8YYnCGHZEk
QxUbkSC8onQIgoeLMLqPLFzgyb75hZM727jsF3GIiw/bJj+0rLQqtlJ/KIqqBaMv
3EMw2UxRT2cV3bpiK4qsAoEIqAOFa+Ke9yhJxhFEi0JnGi1c+IoxvgKXLVQ0KSw2
dfKmZYkhaP3lnjjKSxp/QxF9pnMVx44odKUYAUAa40NEHzs93rDKO7chaqZzoQCk
A6+SX4JYjBz5HAZu1H44MOJ4/PLr/Rz8ZgcgIGli3dz9qD46Uef1W5D022MIPES/
hTJ1EIv5TPYSceqYO/mX73CQGeJx0TSJojNh9a2BjDfnixDGIiYS2kA7U6cctEJb
O9wEBWVjPCf0UYXpZ+9hsV4wkch4kx6U+wlcqux2a1XwMqfYJ/A2CVFpnvGlQfw9
oX+maUwRMrbbDpXplWXFeiUQSuct3cu/WUYP+GU3wXTLGpzdqqeTevcg1ehIac06
rkv1If7wd2ryq15qxwHh7UPf7tb2U/Lne8qNGWjaOkHLWgqtdxbT6hmM4o0Unf2T
q1kh5g4UR6OXYYqVoLHGqKXuHZoSpbwPqwUE/xPT9v4cHneHaEZ11LfD/nfUby3D
BnCai0aqmXN8zXegl+EzVflg2diDnNVtmtQaFyllY+r89k9s9fxNxpt0A9K1lwHL
tVa+VbsVin3iVumu1Oxypf9yJFCWOINWNddEChp4yLshccxbJEJoEcjHXX+MGiVm
2yrfLgZPHe0n8ze7op/xGcO160O5olwy7htLmTm61ztWGWvigbbNwrisJ85uaZLT
7vVvzU01bcaz1hqYtXiJ86qjHdGOkYCd03JK/upK+a+iFNQ2t/omc4szZ8z53SjT
L27N56f0wuFAF/2AP5nXjpy/ZnXDgOgc4yoa0kHJfI8hhdpoJ0knuXeMml8khldk
Xj61OCuadqkN0tyD+pF2LKooethRMOQWrNCb5blXpyXXXG7RnNdjducwpnyxiLQO
NxxTkHTrjKGTh+ViM8UbehrdIYMK7aCogGUwPV16oDIf2KumRR3oNCfh71dza13c
YulZxycn0pVn8h1V6uddmOSP6wlTxCDMp9IVD6NfZ4hhHEcEPcjAKKoJLdmwnNuP
R6GeJsEhzP50zGW/UgZoKCgxmwzZJq3GmipW1OcnxcFMfxkX6793YTqhyaRnXNSb
Gds9PBIBpGkBX+F3z7jokQrZftzA6PRte2Sw9DCHpt5STXymcfNR0Kt0BUxC7IeB
s640zNc6qEbkj9weqZaq3tObkjXr1fbZSyPDFOxriMTwOpvfH7U7gxTCiL5inYbJ
WX8QYi5GCY9B7QW8qDxjHycDSH29S2OT+b/Zkgq4aI4h4QPcZBqyEQZQtUzZg3QE
nzUG9g+nM5jJNWVuRD0GKy7nczFce/4SW4nrbtS1fXCVpdrTVX3641o66Z2hdt4u
zV0KRWavabDkWqrbrr78Sn+GLo94CPR5WDSYfPthrhWoskv9f4+6jRXTqfkGrMEY
cR2YwfrKxx1I66i6DFvFGqYQ4XvZa8UNqt9PoVWGupXAjwbe0R5Gaz68mFrjHrjz
IQ8jzLx6nKswd5v7+HnQWSq52rdzEhbShLLAP4YCc/Tejesd8pAOwJrMMfVZl+A8
ymRXam2JPGHQHraZvtFTZb6NinF93TlOpF0T41Ufca9CZttJG/G3peHg4cAmjb9e
PqWvhVou8FYuwgnZZn4a4+xGfB9CpwniGA3ZLZv5G5OAkERl2FgWNW4mZCFcCG96
UopaExeI7bCAKvA1djP1YBptO6n1B5dX8dMUYR3ndCaIWutFjJnPKiMGpQpVA+vf
f79cgsvBEMngwu2wa/aVpBMme3oYUGR8Pu2CSi881CxeGG8/5EySnolVzcYRcM3b
TNi2mPWn5CZWEVxQsz8OtyqL7MrbyfVXhvkhJrxqyVX67XzAgyUOU347yGgYjEsK
MxiG/+HBerYKbBQFjal2ygj4pboXHd4G2Y/uRRXfMH+dAtCnNTF1ksszT8sCH5Wf
q3eKMuMY/qXzp4aJ/tmI01Akf5THVgecs6QU5FyG9PafqEH1MM1b48PjVczFJlVU
GVq6e5vWlVBrGoeXW9799367VGu8zSVPfqgaMHfI+IOE0dv5LFGf/wsDVBdzNXNK
o+wd7OFmpuii+lEhNFE3OXGnu8jmSIbUNeQ927er+cQNRcb39m0mwsT48TD8flv7
JmuaZjC2Av8RHrMduOCH9F0RJflT+mMjkBdLisLgz6CnF6LAZOIbUCqxSSQj0mLZ
bYHDCer6a6GlZrZn1iPuVhptquhpJIEdXpWJoV1E34mDY+orxocbujlMAiBolsFW
Dr0FmKyMn3Sbpii6DFM5O73O/eny2dKv2XoEu3vNecvthN7aUyPgwxRlct9Huhsw
hA5snGEPx8wy8dtjfE8d4Yj5US8leqR6ovMtQMxi0ud0/yUDjstUV4Xqo4B6/9V5
ZBhQA5rDhzgKJcmzsIjUJ4an921A7jL4mBMmKkaNMRGUGDR3tqpaJ+5/xU+QGLNZ
Xt2K4zy0PxAO5cLqYuPseli4OHn79Xm148ZUu0KB6c3ptrtAUL5QEaQZTNSDI9Nr
xbIt6DETISUDOb769zr13GZtt9fN937mLHiYwyEB1MEC7ZmtzRXJ5Ay4xwocZm6n
Ac9yf0gm9PAt6PIafHETbtU5/kRiNNLRe+2KCOAWQoAEU5KmOYCUTOoz5Phf+Tvb
r3qhPA8rerHQXtvN/SvUMaRscGkKJH4yYxLSxLIrXztuj9eL+GMWy9USsPChEDbo
eh55rARRXUbEiUawRwuHuI3cqGlxXoB1jR5pPcPhfFMe69WZeRMZIWyEr2dwO3pL
kJJHRSdX5YxJl7V+H7tpU/vD9B4vFyjJJzH3KCFSKz5x8l6Ys6PSgDWpABvjywoq
M8qcOwngZvmHWTC7YkR47m1hATam35QKqRWr1grtu8VoDGow/wDnwAiVnQx6yKy7
HfpQNGbxHqUHHCCpoXDIMGWwFHt7asQCIhVBDtWaDrxUlPtSp34BAE0uPYPi0x5l
7nwndUr7EvHXX7+GTt3VnnFNaUnL5WN8hNrYX/8wGGVzIJ2sTdCC8i4A8KwuGJMP
wIWvNJQ0jRNKGdUmUa6AgI5cft2a79eC63P/9gO6ij2SN1CITR+2uh8suAOjXrcm
2fU4HtaRhLSH7qhDH4qLNmW22q+O8flmaLtRjJ5ml98o44xjAKAHkGV7N/dXNgbP
ZJDIOxCEyF9fFUY3MIbkjsG8OWwmT+j9vcu145PKHX94uJ1SXrQSzbtFkDfn/n6A
ddDbo2qliKWdassSSSX7M47mJCAKDaNZRe+0xhbns4Z1+VDGvTJrrDj+vTkxbuvd
K7Lgv06ajgmfAZ/lmYChgeINYQcGR0HUCa1Yl80J9IK/f7ewbf58+1Jy0w8Ud+eG
QNX1nlzhByQsoK4BYzQ//uqOwmGjn6CJwsBczFqsb2Cjd9ie2KoaX7Kq1VHimgI0
m9arJFEqyaUyiTZMikl4NVWg5fd6cvQR+Y0JL1dpjMWPty5Cnb9O+fze1HEEWOgA
cubcsYdALHo8RI3Y2eo4Nw==
`protect END_PROTECTED
