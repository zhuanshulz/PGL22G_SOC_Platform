`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6RPmdMxTgpE3vlcw1+7NqBJntCgLwrCBWEFP3YVrlwPndRduPwjjlFO6cdiHXhFs
10MwIAlLF9vguCzllX/toRd5YJEKdqprA8txg8EpdqPOAfnJZe6isSP2krJgytEl
LApKwg8sxTmeT8fXSyn7OanFSYwP+RaZbZGL0PgWq2UfbWZgNaW6jCJtFZF3slRm
9xlQ+6M1dzRgY+O6LZqMKtd/9XzIim0saT8vyjqRRbmP/1AZ4+rbzJ5DFIKm0dG6
ZWWl9GNh6wnUHuKO0fbYpFl0vNk4XGzNsjErhHfqwalDxxB0DtzK3Wkgs7MgnZf2
QJ0PloJxhbEx22ThF79BNjfCKQVM16vALw68Ght0fZV5ypnCOz300LhfLCJXqGKR
gAesnW5+Cz1WsFETyDKieDEM6ErjWNtbA3YmIP1fl94NbSgrNST/IigIWl6XmDsf
h67dJwOJabsWapPwDZqZBBHoEm6M9QxXw99Llgr/9lmimk3DZpNQmBr2v9S0c1ls
EasohvOxEOhpmWbbzanYhGUsNcZDxy3eo8akZZ3GnCbpuacPwlt5qXm/FeFnWW0d
DKQqoVves2wXlQ4T0YAeEz5RN/X/SQnrhsr8YivvoZS/5a3/VaF39uXfeq6XbBnu
jW0ERI8MtuNlej/C5DfYlvtQRBzFGjcoU8tWmTPeKjwzMVSYv7QoF/9LYdVE2RxE
jj8cnxbGI/imfdvz3U3soq/8jQxQ0tyDlpUxW7AleltvA4gGdlknVufhPtzQyK6z
JhQB8webztTXP4ZCea74+PVoIz5MNVswSHd3vhniG15pHAnU7GgKiQr/8FCt1kfP
mNwdvg8M2sgtCcY/y90JxNTaL4s0iVzsnnykK17wrmJ8IgwjYc7TouqbYwjscdk6
SNMxO94fTZIP9hSu1Vt9wJDSTW8+NFQPh+bu+LZFY/DK+lNr1/8aDQWrlKRXgkSP
eNzewrXMvemNfy5+lIKLdK1PpIsSmzA5gzevVXVbs/FB57RtO8RjA6+zQrZJKeUT
Xp9Xrb+D8+7h8QP2DbmfrLsq0NI+I611aMrUOmZDYkygBntq0GnHvfRMgBrXRZCR
9v1JyBXtT1JE0JQ4TsYo0q0AmhkMLMO/XP63/nXOM3k/Z5kFrNJUjmwVSKz4MxqZ
fw+tYRgI7F76W5saQ8zjVJRufnAiAWmSsDG7CDd3emxzg3vdOohxtxZaJmkA0JTd
xNj4xH5CzqCDUsAmhg7opDO0SmQ9THyPR/vMiWBC0VIoIhkBUErfHBlAwfCRP3RY
YUMUL6eQoEIfygE9vt15RH1cHoLia0NhQZOW/OQia+vfBpUJd7xM6ZPGpeDCdjwa
+OxJzX7ZNqPDTnKESr1sAc1h/KhOra7Up160e9Docn1KM+HTotkS7F5sjT7sEYn3
/dgt6ro9vM3ujlzLLhjn8erIx0IRJ34Le7OsI1hfeb5jO/4TuoArSjEc1N2ZJeNC
7dvAAlUqfmkHHlUtVArLw0uoRqDusbscTXX4oBMBv05XtOrLqEKDDOUOvkO5GV9e
wCvKSMypZ+5+2BHTpbvp9B1K2ARYevR8x6UTadH2j2MAD9EXa3QERUcD9e6VYAy6
DGhOefNylggiUOqv/AoTWY63sJsqqPxWyqVf43NRsDWLnMuPfPgMi2zs1bZyHlP4
5pPowtfeTRbt31ocgsJISGsCd3WIAM/Ych2JLugvNtT7nN1SlVsD4xD4DngbXuVK
vFwr7bv3asWdH6Dp7mOhSU6OgfYliBzerTXVoJpAkCIJ+o8PWLn49Dyo1oZYGer+
UReMGSZzeVcpRIn9mweI4Y6vxXB/d4FRmDD5tWqiD4PrTlFIVj4/kafRW60h/dgd
6jT86Jof38X2CCr/5U2eJw==
`protect END_PROTECTED
