`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qkyEmE9JB++lLO79a3qKh+UpncruKMVBrq4c3FrCYxAjnvHJKp/gwUQd1E6tukcN
7ULojL8ltziHLbg2B/So9KA6mOptC2sjh6EZkEKhtqvN5wnDBNkGzI19GhJUYP5P
qK9PmUlj7mCE1pq35TM0mLsNCvUMINfiPGNepyPUOgrwUvuYKbPbJ2VfN6pnen60
zWuke/1MGYLovE1pCYPDH8DSyfdckA3HW6ON0J/lcDLlcgdH3BquScK8m0wqUU3L
bcY9MrAQ7qYHKVVQCZz94YlC2GMBryCvvdVWVaczR6+L8RHQNHPjJdOXnqEu5ho1
vuva5/odgoyMa91pKpGxTnXmj55fHpHnfHTUkZcrUuO1JRF2ZN6QNOcs2SsGgPE8
TFF/GwIY2qQqzlRON7XtEg==
`protect END_PROTECTED
