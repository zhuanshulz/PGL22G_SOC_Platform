`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UzfdQ4o64OPXfjceu62Vqdj7xMY7QJGUwTGDvZWDY6gKLyJsdub+MUiph4OrsFGb
TB6cBXOVz+Q7aftqtGgkR3tdFlFaxEBxqz+zexx4BAGSzchDLQ+Q2NBFDlq1Abvw
t/oLGxlm6+JAnf5RfAUUvFodZwzQaoZf0UTxq/UkrfFclbE8led5d5BLbm4FpujF
DvY+fdjGsH0yuUlFWvgpMlDHduZGYCzHYAxtfIx6OepB93MpJSJa8Vye9lW8JpuP
mxhsbnvF+fTEhRgp5wccLbn/EGGWNyAHvQM5iz1HRwzm3K3myQ22YLKXY2CxyFhN
DP5pqnrNQ6Ce1D0RAvm2KokFPDX/9pK2KmuECwHMxyO92RvkR990g4GeJAEUUWzq
6/u/U0EdX6XbJLso/5jkxBEdlPb2zC4vVbstXKH9XASDX/bLzsiG3chmpExIM/r/
el++M1/cUglAS6krUAZNJw==
`protect END_PROTECTED
