`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CMb+c82QcfISehiwS7lv9qlQVIwXjRdo7jYxhiffd9B0c5JDBlAGDakMG0AzxqMd
+x8UW3K7XmR+LY6RN2xWoEyNoT88Vx6utkJEPbLMOaZcVveKvxAsJmxJzwqoUNlF
vB0Le2pt3zR/PEUqeOZ6Xw29tUMMLgzLTNPyTZLZAF7a7JnVCn2oiVmmz7XGKbKz
A6OK9ccJU/nd+FOW0WDgWZBaJTEWdsbAelVnhd8LuzH2G0/jqmM+ShUoJNGwm6yv
HJ1IXb2ehDBC+fTvTCPf1+GI8g3LcYKUDcw6aKstOiTocElpY3ZxJtK/afx13Dev
51QgOONsaNf5sNZK9JuiurIayCFcUlJcBAzPV4wz8IDhlEe7G4mIdvQOpCNrmHls
HXFsCvyMEpJ0m8jVc2S3LZ4R7KX6wybe28GaOwt/97Yda62MWB6OoQCk0uYlR24i
eKQAAUBA/Wd/rgMBpdbAm9yvnqxnAOO5l6plqJ5wqsq6anE1apF/DhBgJcs7/PQe
U2w0tMBmsSXH+Yw5OexWASJPVxn+zm0QzONSTAI+STusZv34YCYYzypVudUjHgGm
a7D0CTlz4u+kFIvL5QW8hx4jXNkWhzRDQ4dYCX4oARMlYRXaR9qAQe/Ed8N42yo2
CGgnDGz+krMGi92iKJ1yFoWQ+Grxw8bEwaZHY7ez087hZcQ1E3V57m/z/35pq7zz
tzmBBTKYTXpAkh2a1ZNJ+n3P6H+E8tJu59u3PrYLKIYBHo1Kr1I+UMCMWYybyXJ7
KMq6kLVEIHkxhlySapzFE7c7CXHAbl+Gj+liOQBJ8Z0kcY6Vv2Aq8emJflnBztH9
mSRAb4h3grXGlYCGQE0mEAgUb5ebYnvYPFeXhDw3IiSK81kxegvAYYAOdZH27kRJ
aBbCXo45wXXH6UOUN3uSvQ8PBR/FURzy0pwwZt6liT0=
`protect END_PROTECTED
