`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cM9O7wDVK/9u/PVDoeUOw6rZng7pJCcifKNgtmYQJFE2l7H9/KGnyaI6mOrrIQMA
hVfqQByWvhRM48X2f728ljnsa98TTocDFifzVfLV/bL8thnBtGIKwqcr3Y0ZnXpw
gThjM7H/ERj6Rp4FGkmcHIOVLyzAEi+nC0p7v+3ZKtMYEZnRHcOgio6G3QpmcmNK
PzWNi8BOqtuiuQOgY+6P3ay+qGajhZfP2743oo0CGg5MRxDypDR8h5eaUUFEwS76
B4mIVFkRkxDKZA6j+KmmqwyDx/5tJ/shM7ELM5Tj2d2PpglzpD8nylJuQ/AM9H2m
bQ9ydAZ75hRp/gXDVzt0Jwoe+eI5urA3T+0mJXZ1orM8+g0x80CMa9waMXXuLJnR
CvuQNdZ6HmfZR/b4AlSHCwWGohQtJSN5Mn7Pc4ij8Sslhn37IDKKgPutUiXddugD
ycqYpqUoqRs36d2JEBtXojre5gEYr2C/YyKA72d0XW89YbWNIXnUEtVQQa5lZCuj
1O7HsAyPqo9PWzKFShJnJcP8Pm42krIP6fhLYQLEIxhT2pQ68SD9pJG0cUbmvDeA
10PB4guQyirCC583d2UIuA3IpAlGNrzOdwa2ci+GPIzTf99nOpuiCok/9+jqrdGL
UpOFEWTo3LVzBXHZPvUwVw==
`protect END_PROTECTED
