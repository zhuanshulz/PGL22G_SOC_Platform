`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v2d2VzEjSzlr88R5kdbNFn6H65UFTbOSLxOh4o4tRw04h/IsduxiiXI8cgMh7jd2
XgwISYTJBukgCS1d3H1ASat8umXfaoB5EOC+TXkcsXbrUsSaZ8I+EVswyttRj5r7
TtoViqET/0PSDMplHH0W980ox39DybdREaaR6kObGOiNvGCGIYfI4wpbJgraSseX
KTYJC7aXNVtMx/HC7fmMwwWaiekUSExa1TqSQYqom8Muuzu0IWfiWM9pqifBavrM
UAFLzyxJBOsbOBEAQnOPyaI8uxIeMB5LuYNBWP9i85X+Peh3h1xsicQDqE0OB0NN
AT+L2gup0rp3veMVSm5Yiq90mSgoe81grkMx4im6MFTx4dqcaqog48dkZhG5seH/
m9ICsM4teYOfT3z1A4YowyeWZmwEnuDF+7XE79hM3VxhqPSwO1xlYZxFeXNaBAqR
ewIXuEQIbzuzlnBjGyKvODc+vK5ANwvUNKQFbUFsvPtmBgeTTGXI47ovwiVkUBl0
fjkumIP3vSYhcN5r478QtAp7Sxgj6FIlZ0feMw7Cx9PiAB1jb6XdYJVbvaPHAy3e
5WcTlJPVAIW0Pgpo08ZvGohEFazW+FO8/LQ1hLln2T0qE+wPd4G5TcaEkEWofyfq
Zf6rvWnJtDRMWFCvuxLDXQoQtvdH6Iw5jAS/+BUutD664nFWIz8Bu+xDOYNzBVNN
w0Dvn17u1STPSU6Q6zz4EI+8KDNifxWdNAaMmEOgIjWwKGQh/6++SnkqDoXUrpx6
QSfS1AqD/Y5Eg13/WQbChDQOmH87yA74afsmI/x+9z6yyUCNshspRZ/qzyu0tTya
4qNpcTuxYUlmSiIaQ62s9A==
`protect END_PROTECTED
