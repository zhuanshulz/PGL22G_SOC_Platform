`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UGLg2aBSOleoZ3IAbl9OaT4yk0moVdyDTn8/I7lPg8ff9pWAXB55qX3mT6317576
hjOyw+AqUeeCJlheYnVOCThHB41GsgRaUPgRTg9GlyKyFEY3PDUzftAE2Qj3YRQn
CSNIK0ceQddesK/bW8rZ7nG7ORLUT4kqsDjRkOCrMfsjX5HIFtF/KnzDM76LjsK2
lcHEnQSUtyuflAPOOxWy36lcluL2/+zNgQvTlRxUSDA3EF9DYyjSZHpMXwO2CdKh
usA61Mfp3GAaan0nCUFDLEVr73avT9maaRfSDyP7igh7mlvHg2znCAuHE8HgikKU
kuJ5ek7tuB8STsWFtqQPHlFqjkwKmO4haolDyu4A0dOEIExhNrUxMAI0Fa1gAA0R
nGCruM9keyGbmIqWaQfL5ARrpTscSdh2/PYd5TdFnR+/CwzOiVj1PHmKrVqbAy32
fEgiZ6USzRspt19vmAAWv8ov8+CNnjOMpDTnAet1/vR5I8LX6djj5le7Tb+2Xcl4
so3N7zJTHmdjqUURSMo92LgMJ5pVHDSFA8gChaKmRnc2VExXs067H4RB3V4n4zWW
64Sb7xf5qpRVU6bVG6d8uwd7yTC6wef1jS2kREIEd9+DBjJ3yJ26c8UXddssHxwh
nNSaYhi7ikbirE7tgqMi+y+Vewcqd3n5HpxmUkkUv+7iCgwKFX1zA6LGeeBbjeW7
HKKzTTB3ugpA6/lB1z+5taNXv1eBIPeK5KJmCflkSiU9KOf9b2Ni3wDmrc3Y17ZD
Z2qMqN85fuSpAbJRgG2CFfucHP3cU5+ad40XZ/nJS6i7j3LQBwk4Tj38K1od1Q1r
vIC9wRC4dW/9bS9OyEH55VW2E0GQkvpqzM0kDsR4iL4Sl8UEd+nZaXQI52kdbrpC
DYjfGowajexHif1zgbBsuoFhmhF13oElcYahZ3FetmUzzY1H8gJFljlilL2QCUkq
0X0mIanWfWujitO3hHaU9o+ga0rxk7VUpuK3KTo0PU6ODAP0cBbu4927NRkcdzpF
jpMb5kWoYUPFvyU93mP6NIS2SuUxO39Q2I1B1SVBzm/B7Y3WSeXph+tUB4uuI4oI
OfDUPVZCz4HgA4UWNf+2fypFWs/I4Dd5f+MJxYEAWRyuoAbGRppo+6PjnEJ68fgl
SniyGA/HdVm9HEze4GE2ZkgTmkvt3lVbUQgRbeKn4huNp+NOICgRa2j/MCtlR4YH
uOMUrvNMr+0o81DgSHwoGDD7vw8U3+FXAvtBYrtQ/n7YtN9+jixa8Q3z3GDcYn+X
HQBDKoUa2wWAuc7/WzLZnNtYblIAiTDBvwud/9FsfqCg7kep4w6x4szTyDP3L6zy
r/sOc9RQAl3waWfOMCisY+eg1+x5zQLWz0+803keLH5i5ODQ9Bjg7ZsDvuShti62
/OmPagThh/shLcCYU26S0X7eRZ8dKKMSDuHHqghJIsEsW6tDvn22C+cpDLTF9GUo
qE4PIOeIWBO5Sj5k8G/B7guP8LOkRUPicpCUAzPMLYLj6PGhfh6ExSY6TEQS5Krn
sGNyIMohSSNjYvVLejVeL5aYNINAfAX1IILd3DpvTyUa5OSjzLum5v1UsLxi0bzP
gclDj6ZgzRJBwaCLSLBx/akd2fIy4RvD/Ted2jrDOPA=
`protect END_PROTECTED
