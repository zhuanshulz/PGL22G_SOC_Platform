`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
whgz0Zk4DPOCIvMgBe0jxh1LL5nA9NBXIV+cmJUVgHEfo0kBeb0NfyKiugoR9Xpg
H7r0s+8UQ5MUOHgpg5Ckaq1LDNhQL3b9wzTNRoyvdY6zDs3WMi7XGUd+fXLFgUpA
Qsa4g7U649QhU2LelefCrSmaO/9pF4og+5BGqjz1yCsRawsENXQygUeE6VTzOiVL
+YLn0KaCFc1plBc5rNhWomMwDJLw7HGaYjQ6DVBQhL6bXtsuPptcujWXR+1A0hbi
pRntMr9aqrskSQmOu9YTr8J/rJtz9fa22m3JFJX5BF6rYNd35e6vnem026F88IwC
AccT2VnAdDAastx0gdsykLN+CG7ZNU/bqYGTX9kVCJE+3pN4BqoEDuuB7XxHbkMR
yMSZqbjJoHeCjVCClqZ3kj+p1NvOFDZm22EJnLVojvrXzAo5gMfzkOLoV6dpTEx8
TOnY/BgWeGXoCR0q204wobF3BOnGLPIeh0OsltCeJRBFJUPEuL6bBQb/OSoYFrgI
yoYVV2YkEmVoeat7WFV3sVoO2Y/gY5eL1I2u++Z3ykStZaWzy0KyF6kDBAaDHz9M
0uDErZllV3vCL5QLkeOdMK2dbEqZ5+i8OMm0nqzDIeEIMeQWcdeuvzauaGKk1/Gj
RufNJaFuLr0F5O2drKtAti+5BLcpDlPrDZ4XIfjUb4VwxVxLpBISdLCFkq3UTMTc
Lbf3oIeWvbl8kuQxWOykBudhAUw758PL3GcEPUv4Uxyf8YXMos6wkpE9EGrobi0z
SvKQZ72Zu/mqPO8loDIojA==
`protect END_PROTECTED
