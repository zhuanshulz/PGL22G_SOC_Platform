`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SAOfvdaOYakByIUsv60I5+iQJ4osC/KjdcGdSP2Co8f4PgArXr0VW3tGmXykSMZ1
v8nTvDrteAvm93DuoV3x7fvWEKjtTnF4ZYu+SWIavYV03U5iYzX3krulvUuLvUR8
KtURka1NkddeAU5dVsjFFldJa28K521EsUa91ISxXOB5+niQIxyK335Ooiq3vGpU
FAsUW/jWXzSe8KcHKuP5OVp3ucxi/8S7YdY1cHx4MqubpHWCeORGQjIpYZDcT3am
/1lHYX2PS8+zMSzQ/zRCEk58QRNHiJw1mLcr0ZGsdxHZXGqxVSdNA26foLbAQEwe
T97thSnS55kr4hRvq79uvFPxGIXXBWKbf08k4tzOz/b3/AHErQ/YminVKo7rfrK2
rAY5/s++OMmAMwioRKn9Hx5E39e+e9vLWtgPcLNS4FcMLQbRr+x/EkyMkmNjwk4k
o7TdS+nEmxJyLQpZMCEPDD7dSEI4SzBESXYcNbFIz8vuAWSzYCbdTxEY/5Uewott
22bdeZDBPKdQTNqhntO9tp//+A9qgDAKqMARBKWry2StEHKcX0ryz9xMQYpg3ro3
r2eyxOPrH9oW9It4hhBAiuGaow0BNmqZNHs3DvqQMsTV7w/Nb6Isn6K1ARVciytc
kfKNo+nRlTzEkJ8iFnGNvDB79Gm2dQlkcZiPffWsgbpxhnCizszjshYl8bhNCjqe
gbgEmUOEpMQAMhiPmZ61tFlhX3cvwoo6FYPzmLsceiyjgvEBFnBIH9GrT1w7WK2Z
plBA02XNRjlqeTe6fTHmkUG1ffOHu+r96M9Z3v4QLvAowFSzcwfyzwWx9vjhcLg1
3CVOhpuOJ3eQpjtgMbf/Ua5+MTdyYBzPt8ExkrLJEfxFuw6rUHF8H/zP9Zk6uZz0
qntWSUOWRIFFexCyjrlMudRxyhXuweZoPu2xWDuGZQeEY7NiCukf2v/VyF3cAKsF
aOc6ooQGRbVHu+R5HN/7yrIlj1+ZzHQIU5oaiLCrLPcc99Y6slAF+YfGeivrBFvV
7WLoxwzQFxLaKf5y0u0s3ABmmCEqtxnHpfDUyOnl3dT1XueTpoJnOd76k4i2bFys
BK5Q2W83NhM0uj9odjFTO+39f34ncSgcI2+2QjHY8nn4jPgIHqXMq5b/L9nN6ihT
Km28lqUeTo7XvPZU/oiT5/JuG71ERgHHYK51P69X0VXvq2gCcekt+Vf2regUC0m4
Z5az/CAawMeiBFH3Y9SV0YK76r//UQXpgcLu+PHQESLHEoZmdqJy0AqfWBIOg+rz
`protect END_PROTECTED
