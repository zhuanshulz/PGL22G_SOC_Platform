`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2AhI0qETXwRk4aWR+W5hdz+7/lH1o42AEHK0hKmIjW7QVAtk0y2qQ0ik0ggezAJ1
nKgJGth4eKpart5nYfIH/53nm0z8CDugO+S7hgxoGPS4Ols0R5+m3Erhg+L70/E2
ZULV8dqa7quNthpp7S4gw9X6pmwvLxEm80izYz4xPAUMTbsYBvh38sHqm+GNBpOh
/P8o3osxGVnaJI+NF43PNW1ZmiiCnvkV9hoE4/bx+6C/KKarxI+c/b+E1Fv0CWTU
0BlzLdjs3d2ECU5coucheCIYGBjcz8IrChEZBMs+l2cHSyB7bHf4xAlZe1fjg6NV
LCQPzuA1aBMJ+7GvObumwlRol71xIjNVgS6LZVinduNB7HHygvoyhI6BMYH7cB46
3e3iIUYe6o+6Mfr2v+Ob9SgXkMb97q6c0GPJcTl7bzucOULnsqlunw3qsbdih5GU
FcrYhXMoCzQFXLzgWZ0RxqF1KfUR3Cpcehxgh2hQY4n1Rkmr2KdXGEol9MaTKcF0
NTQBDeqpGraP7FjDWFQH1eBaH556m3EUKA5TmLE2cuE6bSnP2rPiaweIfsskEgQd
QM7wm4Q9DoxRjG8C0NmNQzkqxj+tKR/lWrpGR2/qJmFkHphTxgmoWGIgM+aKhz5/
ptkW7+lKpfF+kD088QURthDXYdq6759+LbxE+F3q5RjVdbObvFyKIl1nn4HLY9Ax
s8/6HzDNY0UrkF56fVtW5GKzpM51OBV5M1ULZQ9GI/M3k1ylJOhgJImz3dIL6yUR
96QeErk4qT8zQER+EN2L/P7XYsgG5Vv+pomWoRDlGtu/0ZxgF6W3Ai+BNEkFBG/6
nWcbKLlff/SHSU/AgkGYEv2Y7OlOS7H+Qg1a21C5v4E7k/RStzmPmA8gf9Q6OIes
Yvhr/0vF4JtjptWFZMkdRmF802//2yvNhqLaV9Y5Wy3V9XxgG6JPp/gRzrxfcvpE
5JxqM0Nj75MvaPsx63+j2YsHW08ebMqqjhgZ/n4BaS0O1g3gv22OB23gK9DOE1li
7RuskxkvvdL9ZDGMWM4fKLZzn8NFbiwzKEEgcZHH/YQcPKxkjcbTE8/4SJTRuwYK
hpQCdE1Io5+vetEtNWUwIHU2v37ZPJFsm4/ccWuP2/fKqnqwtidQcQ7nuKwywBbV
HLAYB9MhrvjmizAD5bulREszSxoGRrmv8KplgGaeGNIEejKWdBYaQlj+IB+JdVYN
8ZdRKdb5UaP5Vqb2PlG1q8L+AvTbMR7s8XP0G99NaIvwC+ocshy2BVAvcGw6BRGi
cDk+Nl8Yt3sdaD9VcN0zH8o7gXAiym0/sX8h6yrRfzWcXInnZDr++HsS/Haq9kfs
gQC+cIGgxLbfrpYLG3+qPalNMFcNsmA4drUmFUoA8r0KWGmeVn36ORl4YyfmKk+V
SQ3+8HwgKdkXEFgHqr9Kh1omkhNsOSO0I3zxOY8uUDnGK8UaALUkYkF9sMb5H565
TJy1GsbSrnnl8j0Dh9JjoqeLOUKOtlgcZUxWjs0WCpuHaEfdnKFdWszceBhT9Wqf
lGrTTsRf3GkLp8YC/bTwrX1y9ENVXAMVmraYbtz7X5mv5tKSYrkd6ABp/t4bsm6h
rgce2H3dhjg5yHfHtD/Q1pIwcYNH/UzCscQ0dG6VjL/+7EmqvWiyYFh4bi0ddpxV
PKK8dmqyUja9ILDszdZ8OCR+ucpcs/hdsabBceLP76gPkLQKREfkc3SJZg+4l5nQ
YsVuJCZIJTtHpVq+49C76gkZbxZyPZ1xPDP/IE0Ha1L+ztqV9VP+RNN8zzXKUn3r
M6tLiDkZ1BIZugQEE/2rRKvv8ixuL6bW7EI5Y0kVLldcjEpNdHKm9Hx6JDuLbw3m
Qq5Pmew3RgkmufOuK+ry7nZ+ExiMe9RHX1z5cA7B0Wi0ibDAYI7+qP/Dj5wxTey7
K0NqEtXw4NmgZAY5qLIUmqC/5b58LSup+1bfcE88Q2RusD97QQdOHHoDgxPFZKVG
U7R5+Hm78V8lWC+iH2fdIk71pZ1zNk6C2aqFm3ix5MLsJPyeTc79pmAdhZR8bWSE
q3xzLkHISVwRpjgoqc7YnIMBbKpUIkqaB3rVcGqhYBaxbqFzYkZcGR361ZS9oGL4
l4CbDSk7j1Ufq7AnqkQBbpJH5il5wq89raI+3t7Z+OK3icT4FzWlnFpGPMb3VMkR
rL1/EA5xfPTTphH+/GvIgniN3ILbTFGF/KNS73KroIDfg+CBPK+ZNOO7R7zYBF0p
QB99YD3mEK2RRVe3do3z80QpDgfyZ9DTrrlQGgkiS6esGSp0tQ0d0Q1eKBULzqK1
ym8Mi8ZueoJMhf+zNbIZInXdsJYsePEaDeRw1y3jm0+LCNgI91K+683I1lP3AK+g
7kWb4UBE1riCYnOgNnZKpln6/goXAZYWmQIMlipC+xqET45K4+lFVHtlzOOtByad
govrI71Kw/tgPGniCM5Gr7LyX/10qUX/ApBfWwpMDbnPG1tKeYgi0XYSeEFc1FpD
2ePfBKKTS2JLC/0JNXY+KuLtJu7Q4LdKh9qyeOATYh/N0kheLLchPbA/YcGTKcAy
G8wXcqbnVVtyh8gIiluGBDY2QlutYrYFdNlsyeQ1v1xbmKb//UnQhMQXC16E3zB6
z0yhQe8Onr2V2K4lDOJl5E2yS9R8R94PpGzqeKbchjR69Tdb3fsu9Rd8xzpHOqz0
Bk5YJjks/H3Cp0cZ0bR86I1S2uT82Yb7l5545aAGk1nTVGuSiJ5TPN+3Ga1869Bg
NYm3F1FIN1gyDJaSiAVuS3ybDrhVtXpupM/xBe7KJNe510di0fnux7nwg7Qbx/TZ
IG8sOxRhXTPNL2iALTRg1oIs/klxuGsQ3Ck8m13YajYfA3jg6xV24USWWBdAV1yc
vsw19U3fE3G0YJf7hSFtEqr7mOc9Prbkq/wigl7Cu6NPAt1fdp5QRkHS914Pj4rR
5ewoDh5B0jaJ+yRB2lqqNi6IOCY1UOikq71biThp11RsKrGlg6LOY0RhrvMI8HKG
ZctAFarx749MjOJ11aCLmJmmt114ESSFsX8dgUfwfZyYCPkbOw1GebqAhzgm/+6L
7xEJA8JgtQIRSLNuJoUt89xUVJ6Egat92TvY6s8fZSHM+lWjCTs+tCq7ZHF6Wd+g
CyCgBkLn4YzS/a9F2nb/YMSMkTlCF5eujpWDt5lFV15jxCNaMO2PS3hZen4pnJol
Y12rB2HghoKJ1tPuKNJwZY68Vz0OTtkvamxIIMzQhgecO33NUN5xvv+MvXWeTMB+
cV0K4znUmTt5DBIJTGUZO1tcwklSgh3X2TQmth8paNBOfEmAw3fuZjFYo41oIXf0
Beqla56Ob7+riRDpHoXzqQc+vu1wNMoQRVvtEegRr0Ud0JFeZrGeeP2b1dwir4wS
DWAbhPfUK6i818nNncsrBaSQAgt7hgKww706usehAWSGykwZvtMdhISY9WymCBdD
P3ASFhE27rSyAYnCCo7SsUmBWogV/KLChnxIvwH5PZSJRqG6WlzQhEfQHOxylsh6
ktyfLFw7MvW9wDa6qhNR9J6eNVcUGM4JPkDLh3wIfOwowCDWPbqwjp6zf+7E2tsA
k0dZpJiiGb57Zn5hUd1fK5hBJ4EkqDxwkYjqPaj0tCKN5n7+u6hCrEn/mbd6hjMS
cHaVSQfQzUXD9n2+PhpK+p5fT99nl8hxxy7ITK9SCmQWg/A8x0Jhk3JhAaQSH9Uq
MXrLEO07YhjavdAYpT5FuBB4lINu6IM4nSN10J8ub9o4wxfG+CERVi0wWEoYmJdV
XVGCUBPQv4caB1d1Dlx4dr3IBhdRyslCZ3PWjZ8CrmKuwhKM6FH2Xuf0+NS22CKe
nmcjL2EaH8sjHCzpzoSjjAS3d4NABh1a4RvdmaZLUAkQ9pBQwYHCjLIvI/dM8Sic
D98F5aNviIFWqfn2XzkqIY+yfArVk89Wb19dqPKjjqZbeP6FinwENIZhswb1OhNT
hkYlZ8bbVvmVbuTtBOjRknoSoAeVGYkRi+4jmxpkAAuqu/nep0cRQ4V1hjgOYNyl
54qnFWWG9ZUXaGlzo3Csyo51q2XNtu08dVt4JagU6nxk/kLO5HriOFM43J6WRvgf
j3FprHM86u4HlkVTqxuHXJARuP2wFg5wYTxhGBr5ejBUHoia7BJrSPok4w9BXfpp
+rZhug1t9DjSWjaTmKQ1xbWjwrZCwsIAk0HXL+XFMXVFKomq9fx/A7TEqbu7AxZQ
0OxalfzRHTSQQeYmDmo2CbpHVw56yPBYy6Pmjny/LPaKaWA5h+XvQErmMIuJ1N3N
pBIpygo+Jp2pIUFJFfKYjl08sPQpPVMkb+7iYuZaXHEh0JsGqZkb6A2p6EqK5L/Y
kMhPDSBpMpex3vBpdgmNsHumpgLslo5r6tDmgLgF0bImQGVRjelrIqISxnP9L4aH
ljHXZjmaBarKI31c3oUx12XFsI/nS3+bKU+Rm6Nfk6EL+SbfQxrVOtbfeDGhNAFO
sUKn+nnZmSRKW2MHt2ForHn2jsvSwr/lpu5CFu1yu+A01H2b6GWE97vvRAWap8pl
szaTZ/PuoXoHihrlNJVpIhNoGguI/eOpCEdnJhLXIrPMK01/driMd2sj4cG2cDc7
S/CuAD64Yg0y/ExCPrX1+zsvFWYXs6hgWYYLMVpYA4nIX7YMkG93zYDWT6QB+83c
6LoFaryg+Z5bcgKh0DDgZi43KQglj+X/YL5j1rXa7cCK2FYAw/HE+SZEmmHPRUdG
oxKKoDS5hRiY8E4XfGgJ/HynlsUsg961YWXvO3dAzz/p5gnVs+Cj2uKXyUnrHQyu
VUIfoCnL4jBbEpCQNUkz1Iuo0AeM3EpFCgFMCDIhes4cmIW+gpvOLPRtlLyD+Spa
ykUTdqSAnrXmYGj4CHPaLDuXJqehLBaNYdY//jkyQAg/MHZxAIL/FOQXQfY0VLW4
HdP+xG/18BpW3wmEV1PVwKaLllHOKSBc6ahY6zY9K+S48MCHJPoJTxFZ2JYJj1To
8EVNwzVGj6Gig8SlVPaHJvMpjmjjk7OM50z07y30bJb00q0pisnGxtI8R+LVaeXH
S4VLySbSLK6CwlX75LZ2qSQgmRGTxJA+P5ifL5yYKwToHITUPMuu6y9bVChx8u3N
YxTix1CadnUPKV/iI85KRR5J3XwgSnnNNRwIjdTzH/MdO/+k63kCyhH6U9fj0oqn
l/5imP0AXaUJxTTf3NB0FqsvbwCLqJtQpDTxlgRVyWQ6g7P569ptvrfVMar3icJ6
WKIixkzbFtHZKyGUAdyT5d3IzXBshyTvSNGWs95CWsIStER/chYToOrzGtgHqCr0
xaa9JN4O6Cf/eLZMhceTYkiRnmb1F0g6Mt76TUM2Uvh442E0oP7I8R/X3nlJXMHV
dIAmTA0tJ8yoVQYlM852j9O6iMWCUI5YGRDOaWNV92Q//det5OtGjvJbvTf1ljuq
AdoCBGo8kGQSuzTp75pnTg5XGPMWtLKrPXc1DBEbfGmIFtKADNuZPU/gLOjwkqOE
Us9yoP+5zZTqB1fgoBdiCtR4plLHLR1TzPYHsORScPEsJypo4QN3ZRzco+ju4c0v
vd2yGX5bK0KRRtydQHgPdEF2Oc74XlU0O05MRDHo0BY0M6VE5o4WTAJAqKscywiY
3WzWdgZaerao8BWqpqKdMcRPUMxZRgKWBbh4IGFZ6UuCTRuWHRhs7GJr/pvKgLzC
BvU2/1mz0EY+abRV1zhBrp2DLed7//xscHdwnxesOsG64H1SejiJE35ZSHtxoyQi
oTJo5zmAfRgiaBTpg1jXDj5GzAhDbFamuxZHO74ipK1erIBFPRmtevRYRcbPHwiq
goR37GtvgZBBjfY12RxNcs6zLU7/XEu1QWJvokrVXB/BU/lN0VDdLmQpxh1dy0gp
kTG8M1C3Dkm/kJwLExpVUyaIHCGspeVsSlGUW/PbZTHqJe1LaVdiwrgRTofv0HT0
78K+PhQIGahKZghepsKEexRVgvXgPr5HhnXEBAsHc5G4+4LI2WftHhDQqoM7edcu
h3a9gTeeUxwnhTOojqRv8x1n4PjURs+m614aVQCiRp7Z/+hzcF1O/zW/7tgYA9Z2
iASutUnzj8RN0MVIoniVPTu9T4BjILyuQdxyokx9TEzcBDZtIDFmOiObSo7LTE0B
pZPH65hGrFKO1pDvpM86aPO8WYwJn8uRYWA4oGIfu1jsCpnpEFzHwohZ2tM6vJ3S
fguDu0CyupEyoC2DLnTQOU1gXWsasgzQi2bww4juYAHUkEHCF33ikJNfySr8jVGO
Ga0DL5t3jT2zq222ihgwjJtaKr0/37qWLbCphNy1cAZjjuNVQlVaTRyDQxGCtwjW
HT2huWC9nYNxiRGrulBtWnRUu4AZtOYA3NPHcCELr7KTAH0BZgFlnCeNteRXTC8k
eFUjSqdwXp4fcs+EtMy9DmIolvKyq9v685FdFb+3LOb5fAnuLGPElmrzp7vUWiBw
EHcUwd5cPPvSOAATQpWeKCyxoyFjTlmSUWcEtudsectaNdQP57UvBIqCF7/Vpahs
iYmpxrUlR0FcQtmHbYIbkKpQKVb6Ym3u91ELV0ARHncVLIvMOJr6UsBTmGqT7/6W
fq4IFslTvek+rdmxqIZ9GeN6OqaLh7rR5tpFM8DH069KJ7FWvZC2rr4Xtv0xkrKa
ZcMLnaDP4L+vS9o+tSIOmNHqcmAEhw41jlBtTzKJTxL4Igct93dRrY+ZfRYKEGgF
3GkPt1ZReo5Na7U9xsmlVi8f5irYNCVBnIJFXZpeKFpEv2K2QqWBtSCrOpKoKND1
ImZoCbJsYehZ7Aea82OcREX3+4o5k5Vj6aLNaLe+FhuLpGM2vpLWUoNjbvegAeiC
FrZDXWAUCUV9ebvbpPpN3dGocuFu55n3XcHb8e4YE0b0HSt869wJyd0zOZszpMsd
l79okhecGSm2C2VaqVPJ80vT81IzQtCtJeuutPbFXEdCcLGrd8iQ7eJXjZS6eXgu
lKlxJ4wKtMAihfzP7yrb8mesGVuwQ2pfN05FyNlIp8lydpGxpyPeKz95cqVpMidE
qypqXCUy+VwwrGQ5ZKimKQj4Yhab4GPg9HII0uxfinLJ1CIUfvubV3nJpiDdHqzm
iqd9SvaEGxHmdvVVH/av6r5JvePk613DpzgorVsFYCzNGUAJoSu/Ik79PODxFbGl
bumLPJ0McM47LL/g04mN+pnb5w0tS4cq7JJ6DPi2bnPfDjmiZ8tj+BdPMfwUmUGd
lDbVpiOh7sn8Kl+mhHQlHL6U1h81iWc3bZL0JDlUbkovxbJ80lRXoI34S0yTjMuM
+Iqy4tWBYBmS7VbUMvxbB/fYqn2ggiAmWxOg8xFeCCuo8LsnO6ZL1sxDNFQDT1WP
g35YOhiX+n98Lr/YflJroNfaXq1lZVsdObPXPumkUHXh3qq6usaq5ryGxNtCXVoj
PMvwPzLL+7U8KzsEQ9AQ0utTCdJwGF1nePpqtSPHN2pdeFJOU9MA0wHjX79dVFEh
YfLUZOSI2I1X86+i9uh1ncaRXsVIg+04Rp5SQll/hAcQbd4QiX2qlKWmmeyv1vB1
5ltJqU9+Sg5oWy93+txJcEqJPzK+/b2415XFoiKSj3zwZbMDJFoirT/B1FVMwOWH
+4q7Yi6+PxjRVV1yBb9oaiE7CW6FFa8xpzifjmrF+q3kMY5x9fvDBDcyknM/dFOF
GWGt+n+rVzyd4gXqUs+6JJ03pr61LP0dEvF0uK0xCkZIwr5pbNkgTYAZ7OUBQ1RQ
fi7grdWZ9jb+YmdXfW4e4X2aEuNd/FG5hbuv3XMDCGqn0iADIsil3X3Cwxnu2QHu
jqPj5N3F4rlZBnr2sOXUTF0Oz5U5G9JJ9W6DvLHm/q95xA7wa1bOl8QvsGHKxX5o
730ksE8GcxfcdtmvLnA+NfL0pcsU7ZyuvWstIBSeSfvmPLrDQWSizBIT5FcfiaEq
yvjYn1L6gP9APVbmHc+2ZHHHX2aa0TOV3G77wOY4AYgWkJOB2MPd6ula/xJOXxLo
QdcBMTcz7mgF5YLji0bJMYlMoD5asCYxCBiklfz3fHrrMzFJ9Ag9TyPDPjXbDxrW
8rAcpVQYuVbQD4f38RkJc0seOx95yfuDIGAE7nnWx7n49zDzQSOqiVJErnVlz2gj
kSTY3+QHKVz++s2wEjwHZCbIjUbAyCeAHB60A1CP5pkFDix9GeEAacIzt8RJJ/2l
r3LQrv2F+03vbGXGbJ8wH2XtIDbJvb3Qkc+SGKB4Tymc3f6a9p2p7iUFQsdiS2cY
zCv7scRUGpwLzAX9xS2zg6OAKRgTE8mmG98yfv1vdJSR9bjIBjJrA5aRE3vMiRHU
jw8+guB5rv0mrNXwGdLyOk1FLd++xL685suMbXVZM+Q95quFKaGebVSSKP+HTOZX
bhBa+T6GJThVwjCPSajCkxT4Xv2NsuOkVh6HrcJhvYeAeNC4xro0yAUwMyiBByVd
1L+VUfVW+jcEoxYO6ymQu+2Gl+5SuH+s2Hsgt3aP6rVLDV85kTQMbjFaK7ubJlTP
UZUXfwSpquTPZvtA9/YK03B9zdhzNVzJzsj0peOE8hXQHXkGgoB266lVR32Yh/ZU
1nOBpc9re45plYpC+f60E+qEfNwcWLiiGi7II6V5pQUxI48Jb0yEJ2YqfzjdHNkk
gflAj5KygzaGY6vvr43W28rrW5pblDEkK/K5+kDZJBmC/7gAJFY5FvP2vBVCHkXq
NKXwoj388DMLKKlD/M2iuSa5dcCEAGDvGRRcpbVEm/Q8FsulL/CEVBrfKUG0th/s
nvjH4zj3jCmkCcm6ODluah7OoGo/vuM4EnDjJYlvU5aouqfmFB9s16EupINV/57P
kb0jJinIcfpVnC9GpDACf8Wfz7/ReUmBQrTLR7QK/16J8n0K+IHaGlVjW/cffMh3
CvRXhLpFRC0mQpzPFhnnUQ==
`protect END_PROTECTED
