`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gMQ0f6lRppqkuqtga2/rKJvBEcN1O7xs4D83uZTNfS2WTQTdLNN4M+i+ax99pzlf
rom3B/lKje4oUUqTV2HpKbQgND34z2ZXu/vIpGJ1fnoA3dHs2EmOUaq6+S8F2m6f
ZPkvdypNge44+Rn49jXdouZSYXCqxAlHYgsZdHNF96T5Ls1Zrp0a01qWZo2p5Xpj
+2yCgS/OWG+TyohB1xk6GZ2gzQz0xRTyO0is6H0VCPYJLFfM6ywrbvkkwYMs7ihe
YZKUWCrNSnIYc85dQGdRSANniuC/duD88TwiOJhKDHzYp3ew2opBfZV/9HK+hnvD
RhXkpw44ulgFrYoLEEz92h16zhuF24IDDnXlQwSRVaJgWoKM1vCu5aQ7wbdZbXX0
vlFygIMgostVSkxsfwrUWEmr+zcngq1UtsuoomiUQotnjHWBUO+CtJByl19yBHlY
zwTA5snK0I5vYGs0bqLPYsBwGreb5ouOo7AycSuDK6Xfck7ldv9mOBm5zQ0vRjTl
RzPXYPoHAL5CTuTWMe7YmMPMO1YuVLBogyFPp+p/W1znOsUjIOnA5k1xcHpuNIBS
T2L24LLlunEi53eXpQS9KgpRQm4jkPFwseDigQsAytFi85+bZaSZjP6qej94zro/
6l6Q9wRovuoecsYILAaUaByXZkql78w+BGRN6SvFkA83b+T6uQN0xPG93jdLDq3u
7hDBSZhusmjhbgWgBvxD8UM2oEPNHGrE5TmTm+WZqBgUEuEPvtOAkW6SgkPNwxAx
7hVP8TxBFQARs1/K4m9qz+snygKcFBCl6j6i3OQYpn83Nehy3cnQivycDiY1YMiS
B/dm6UqoyYD7C4xbQmbsYNHUY6rgucCyfeb66E8Sx6FX0MpbloB1LMpdTdIKkOx7
qtoaJhtgXkW0gvTzYyEu4hOn6w3i38MOKk7/naVEuohwRtlyuROT+OWf8L1dqIBN
7wWoEG/cpVfXRYGpcH3uFJvNKYzyLTAV1RJH9OamDtVvcI9XsqjkLwQxMzwT2FTv
m6dMCUP1FQN4Kd4D+tsBLm7QXTCs4lAUcAP74tiF9X8Bb3t8l88Tfc1nuD5NRXcd
Pu3JIgcgiMTcByegbbnUTkyZDksiiquleJzXjgCgN28IxO1RwEq73N8or7U7+Q8E
CzEHaTeoPiM896UOmq/I2XUzunvt+ZjDUFEZ3X2tyPkcnvkwmWUdpP8/62sEyshI
ZMUCI0LMAwtzBVA/ZSVEsT1ZNsqzmlMLD0TarYrhNA1ECdq3cI6PQ8ZIr67S16yM
fM5EGCcK4YH+ohDo9bqND+BLHESdka2VEzUWeplLbBXeAs45TsbqE3zRLhGI69SA
zpopit0sUmzJTiBLbjpp3G6zWBRTFjwSHCJP7bwyp9aGe49LyGSAbFskt1LzXaM6
dRGh9ClNceKT7rRem8LplqvWIU6E+nmZ97VouDOPIPeUaWs/Ct9fsTvmO4AhUkFv
budqr21SXeM3Rqa66Vc+PJESJjh9moOAwZRylTcSxoF02LDwdKP91MTkS+g2bzf4
9VewYaX1jz4+q8Vy6VzUu1YGmA96TwDxcE3qnbejmIeR7QWP2Z82CwR/3OyqJWWI
LBb7537Nfr9WhoF2BKAv1COvVfoRk/fD+isdmHxvV7ZZqIxsx0o+1JuWmOjjWTef
wB7HrfCLyaXkVp8w3gZClxZiUSEWWTenoE9J9g0av5YZuR/+fRD6XXItmW4voj2W
KXm2P+dUUCEZzFUE3s3bE18X0jpy8fdp9KDEckedsMABCeLS5Ep3ltPyceErvZLi
Ft2AWi3ZV038uWxkUrbj+5sqxHeJ9vYPrKzF5KT6khUBD7RUL2Tgn+/7HEc8qdlY
CxtFRik9B4TgA/u44hgWEcpQL8VkkYwduAR13IVKCX9pJK0PWObOyzJyHMlrB0eN
GRj8TrsIRXAirOKmp6WshPp4BJcOlWC1KuUT+YVMn0OaIQGkeuGdYqAPWQpbXDtw
u3GVVbq6w/suvkt5RZC0+BmQXLinOfhIEBc/jNm/G7btQ0Y9qnlfkjigEMMkh/0N
VWzFbQ80Z17cWmAGk5KzaHIB7PApCv+HDbcipEFG/NlP63oFOA5+wx8A/q4acnxZ
CIdTjd120iQqYAV1FsqjM0szEmHhGmmrPYDnEtvOS8OdZQpOeRV9BzrZV/Swy4JJ
lAPtOr3E+dOsc8HBz3LJ8w==
`protect END_PROTECTED
