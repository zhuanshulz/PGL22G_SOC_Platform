`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vTpPVTc+dU7VgMemHKeIf5WmSgd50nif1P1RDuFrnu1nI36U2s0ynDk0h0QSIv56
Dyfgw0mHCtE28K0ChvLbA6Kg5eEbwFSnREe7QcfhVI1tiFngyKi8foW42MYhvwrn
yvJqGLt6eVwG69sjCPkbH+6vcTXyLESpIITvTsbkTLhfiamIq24R5Z+PveaZkvr2
6JK4P5b/ZqhBV3JlFKiwSYQiI3ydaoRytUrhFYiRcuJbh5Lsy66gEulhsGpWEFF1
/T9GXL1mWijyetoK43fdIaU6DhOlfDwfoEarTOpXlv6XOit0A4lK6DwINiZKwhoj
Hxg9x4tZHoxHSDhX8eHM+q6ZJx+d8HSBjo6N3B6cGwTGQ0pjLlzc3CE6KpBJVzWI
C7ExbcUWxhS3OloacIRKiW50iqY65Z25sdX+b06NAyXdWL8Tvq50972wHFsaGjm4
P+fmPIt3rc2W+SUPt7m/+UHZfmiTUp5uuQSXezmHSyLjz/QqA7xmK3BsKALGnd0Y
KKLKJzE4kbHb1rNP8TEqQWuSr5tjKFh8iHcLrzu6OrQ=
`protect END_PROTECTED
