`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ClRcLnEHx8In8RzvVubpvdBHzOwJFMCh5Kg7gZ4/ym74vDVJI2UFYj4neC3bHoSN
Em6XlVKeEl0Rfv+08h+e+KvnE4lCI/5IFr1WO0vYHxSaf9wq1dS3rGbZESeRhJCd
ADsuyPBIFTiGyLTaJ5veG3rdC2PEcIM+Jqv2BkfeP0bWLdnwugQM1rHtmovb9N9Z
hn/NA91akfi8JMkoNUBFK3VwsBev0O6yZh6zispWM71GAvFYK/6wdTbV9JWWqA10
oMlZF5ZsMGeCStCTZfx4E9wKjoiuumrpaih0Lhl/IsKkkrse1qiMcWUpaxN08G1A
gKEmYyeZxBqSbi8CNqoGW5hP/NmDvrk1Sa7JDQgTpwKK5ocovouFODuEjeuMDAPB
Srq6GR5Spcxum1z8E1GuLPpDx6O4UpqgdTlL9pcpsk1duZHVAtIlgzJV+FrjrA2o
N3Hxh863SUYSeHVaAXFEkBRoVpI7BD90t/1JbLPoSYebyc9hsmRNh1DXN68x2Rih
zrs20XFmjl0whkLwaaC5B/yLVKLTwrZVpopohoAvqXsYi6+NfIl2ycyzwSWhW7Gh
MYNIbpxd+GwVkbG5slIjbL0h4d+P0X16MIfIEcM37nyRBV8OLtdfquHD+Ok+TjGY
tuMEPl/gy0Cl7vyMJBAHP2wRlX6KdEUZcg3eFasNH5cLBmFvaGn5HC0wVW2OKSTk
B08aQ/jD3eidl5n4eoBfRQkCJNMCDwLPctnHpTYaUAxopPTxeiYniJhSfHvYjP9O
j4d34hCpk0rtP6z4HZRRzU/3VECmbml2Zxs2nP3St/ToNa+PdFtzy/lh4JNE4ySV
6hOGRXdLfvHObQ5kPkCVLDjMUUm0CB8s0v90HXr418UK9zCybWBWNwg/LWYeCRMF
2m7C8KVn++/l06YJ8GKNWBZBmhr0/JU6Kj0ETt++mXZMASasaLgd7LIJ1B+iNcEH
lQqqBmPAEXNkVqU3jutqntStT8L+8hDfr7zJj8j8wSQ=
`protect END_PROTECTED
