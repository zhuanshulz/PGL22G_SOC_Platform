`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a85vJu+QcUjO4EMRaE/EsyXB0LWPPm5B/R84hyyTkcwjV+Q7REQEOKUySbefic6N
8QhbTIdL+B9q0FufLO2aIF001XNbI9ovgvFjsc5UkQ4a8xWBPURlqjejT5jJIlhz
+PQzV9L2aNNLkhxVVjfKiXBNOt3/GMqzSaVhVSFp/4ioAh8K2rV5h/h6i++Uz1BM
uGRGrQ81FC+bxq0Y94kwHt96YG/PXjqhypetS/D84gqmdqRPHdcMmjqpGrMdNuQa
I82OOHJB0xWeQuOLTYIReOJWNrrRLxPwKb2Xj6sKYEVxjqonYnurZtLvBQshM40X
Zil6QuY4+uJtwzr8e07LFPO2l/hfOLcqnBb5vf/51E2qeHVVeovpqLfLTFBnam8i
zaiTcvbS4pdL/cjNFwGTw9kBFzNgftAWdZd0b+LtMR44lG7WzaTTMkUf3WbAh1wr
Vri3PIR0DNEoYZ7DV18N6uQKM2afQq+6sjmgFFzUjpBJBZ7fqXVRjhP0+pXBohiK
4ZTyj5dnymODN4r9Bcr/QW4MCrMm4F9Ozo/r7CnU9rKX1PqadTs46m3XAVUhWVhE
2E5PDmfue+yr6Q9pq+CLIZdsUVhmeoegmmRbur+OqqLjXt4/vlgltxiW6vRbT4wM
hIJiW9dKWzcya2M25p6Z46pNAq4E3Qzxg/Nv1TWa2Sy+IpWyFZNHggf3La/yJ943
nK0DpnlIhJYrddkXbG4y74rk6ipZEIaZ4dG7FYz9HxHGFS5MVELotO8WSfGBAImH
NNEa4XZC8xXXNf8jW2XN06Z/IoQRGRX8ybkNs5R8cb6FLsVjKS1A1UStqzbLkCfh
43KW7c2xMxxOY18joua9E4q2YXS2w4QHdIxpqNA/UtVBF8nivl+feFzL51oGyEN/
0BwAcP0SMS6x8qYKWUOzY8UqoYVLp51WqkRjUhbZZoAsBEk2ijZt8j1BNThP4tEr
2LsVtAPxQuu0dMKxxOpL1Ucv2XZm+ZigwJDODnrCXGcutrL2rL/0M58lsOoKGpov
jjTTl2y8hZ8D1TbL28GFm2wvPeniYnZsuPeN3CbzNYGirS94KlvsAHibb8uv6lfn
M1MUwEQO5ZDqXTOrMgfdEVTXMcvwLIpfVo8P8L5I6tFQPDCuge4TJ8R9ijbPHPrN
z/QPVo1Dlk5TxqJm79DGzoR75xkYxIeWGrjdF0GaZiYp7bltL4/ScbUAL9HZmxWW
mW9h4FlNL+ugbtNTs93xm1ADti4JATtZv8AbiCu+juHzs380DyuN41V9q8fpvhel
TnTH6oAun0nMq+993YbN3pYOVXyE2C0I4EjCBAQ/Q0qWYPwRprkqQEqws6t4H5RN
CEm0gwCe5UAqtylbqM+l3qqw0hsdhSfbe3BpW0DG+f6oMn92L5Pv1rKsAFROij/J
snKIITKF50aLCMPnmI83Fi6x7NyCCwVlm5Y4oqDXEj7erzMqOspJOmPjN2bxUJIz
iQssxSo9JZBmZ4B/JyCCco8TeGIAVwFGdINcK6wNSygCIfPKrzZbvt+BJNeQ02bS
if/YgXHq9RdI9/GaoGoxyAijoTGUzDAuhO43c7elGKOSbgwSQQs6d7gZ4KnrwAsS
6LY3+9KgpPgAtAeu2emH+2ISZQWDhs3xZ4zeUXBwcj45rH0lkrS+mP1mBPHngbDT
qyk39v0fdwN3DQBZZkYH0YOSkrzEAC3t2MfvoS4JXtLVe05UhnG6+VgBjVw/COq1
l9iIk5eoqPZ/M/IvecEH8XeJTRgEiIEUj7qTsutDsaw+Q1gl7fmzggdLUeO6yt38
XlnWATE6U3wm2pLamaQOoMJ3uYah6JXhHP1+6WtUHSUgfNB1l1xPj/eolpDDB2rq
koeaMo/H6F947e6MzXaAYcxJUgpj4eBaNYXvW81P+avGA1/i+Y/A1XVhU72jApmx
3cNBUkNUlSgsq6EDLJErPw==
`protect END_PROTECTED
