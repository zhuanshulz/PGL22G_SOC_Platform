`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NOjarB/bB8JhDfjOcdzdLrgItCvPqnVkh9mwh/HvsScrlS0BnwwxMUWcXun+xwTM
MDvXoCj6A66ZcrYf+5wnpTGG7dErx+L8mzywOFdsJhFYm+K0U539XVwhg0pRwWZd
ngVE4L9Bp5QS1bJsKvnnAhgOkU3ahZ/oxIfG4165XWshpjZtrhcfhJmG0dV3uSsY
wHXTXP9ZRmr4lAGMdVl4fpA9a9PDMKkcYnLsQ/4BYptn+Fbt70GwnyGIaSQcmkRR
EVcTya02N8qZbbRlyPUnA+Tmdw2InYyTX/gPnuinIfH09DxtXijVXEFg3NVHGXwY
EHldG4NVJfVhELZq1nWODyrXawGXwWWQPI7cQaUpFssuvavbb4kUwj6kkloYkzh1
K7uLvzUifanTeoDcFiMKqhJpWL6fTg/5NbRkXAk70/5aeeby+4JJzLVLNozEhPMZ
hPZY9jWv0QnoI/lu7uUMQzXK27NBRLf2CR9Tq7Tg9NRjoOwhpAWRNK04dH4UzBxh
Ix0MM2Z+TdXkpvu9KjcrnJyMT2pzQngnpO3DpelvVIk7HXI0HCht1LcttnE/XIfs
dK7uUCLOn1AgFw9Rq1L/UE6bEhP1NjXv/rlzBA2Ui9BpYnVRe+z5NimHdfhvaY7s
HMGMd09Q+GNDfN3VhoB9WbaoWEyN8NNRucFwWZA6XLoLa7IC8G6o+zXk8AqajD1D
GnIwJPil/z367ckz5Gado6ReWa9x9586O2M3UA6qd/mlx/y1mX/nrRzvr6U+DelX
KXnrNFmZqAfBc8UBcNrr1mY7sNsepTh0qy9q5uWUi8uuDdaMQnYIIxAnaZ9KqlcA
/eMGxayux8sSwMNsq78KbNYIb1/gx1ECfTrRdN+CSTqXacLSoJAfkM9b4Tu/nVbb
9Z4iIIXZbx4kP5/19Ynqh7NHpln3fRme77L4JPfWJw/fP1uGyutznnHYLNhlar6f
NEE4uiDF/cFktFIOQjkIZPmjIC1mhCprdJjORikIVQNyUEYlybFoq0BotJgvQkI4
q6jsIAPHMnKMoelMDX4mapeUaX4r88u0Qwz82or7dsCE8wdYipISM8EMbPtztHGi
43QW5K/Aepxb3KHqN+gmsDW6/bIobSmHY1uBn4+7Zc0whS8YtHdl7O0YQOxm+o6l
mUWIojhjXRISIzbWfNnDbOsI+ZYkl1powp0MZxlJfGU9PhwQz/iD9VqukZjhq9oa
NwXoa4N433Xq0fDP6hBUwmwWux1gvVB+BFYV5lQ/91uia6f14TfmFVYJEjwSsX5r
njgQWjvYQdbpUM3+pPywhVTryVbdPsLgOwl3Ltw4Q5xGAqgMgLt4KkH+Mx0Ydg7F
pCek24LgPA8baPrYEFz89QF+WD4jIygWFdLmxBrs5OxyGBpTi1G9T30LsPdJB3Qe
CeEBxb8oOncMPjIlXXBnWlAAZ7pV+AQLgU96uVDdAMi+FeWB6e7y8+plLfj/+2TD
OhCJ8KkApPUYTTngHzAEv7Bh1EeJQx9LqKr1zSz+e8+BjK+eI88Sn/8Qlw4pSQge
hYRs/Sv71m5TGKYDxWIThnD3scvaZdQBRR3iubjE86wYZM3d2E6YfemYQwUdK+m2
7X7QpXfpUNWLIHD5nyx8qgkQgOfgzzwE+H06GtRzvgCTRyE+sGTSwwRAhZWxFAn5
ZQ9RS7w9GRFSm6a+drQXMVLpiTUatSZG06T4YwcjZDY9l5R2ZChmpAC5v4qSqSqS
y2XxRbhPvu/ySiERTuRC5gjYAUMAKt5QOmbVD1kUEyr2PDjOYrijVEubCPyVOl78
isqYSZPm0S1g9r1ES5psNys6GxVOw414YrBlwdOAU32tirOfj2ZkIzA646zqDyH/
UAqqhOTBEKVrExei/20eeNzidGUGXpkdAmmgaRwVmksgFmMU+tkZwdIt610bUdSg
L4FiumR9lYFH5URIkCEm2ETCwD3/+VgaluFBRqOo0toH3zerJgI4zFQG3zXRN0EJ
IrpAGl7bQ17FJAOIGx4W4a7VkRZEOjOuELZKqWBFVnjUuHeJwlYKMyP3gbqbzLZH
pBlxHLVB43YUL16GuRoVmcpmElLmRqLsB2eQcSULDmPdWuYQmG9k5yQ+/3TJwWdj
DBZcb+Nbdcr/2YjTl1d8Fm/O8Cj4W9DMcsyAQ5ZbsQXIKElYXV0M8jLpzM6TRz9z
Yy3tgkyajxV9fdinbXwXhvDhMPdFnPWyuB59eaUgXzyYidXA0W9sMljQfOHIzatz
68Gg8heBzK8ea8TMU1npFoEwCRRyXd6L0tBLq+26nrGjwHBk4bH4iQPWsZ9lRTcp
JKYpQrFjzVeCYG0u3AiDnHOf6QW/xjK+H9GDjCZPh7bnJtAfB0L+Et83CSEW/yv3
MDtxvkHcX8xNMQ5JjKQ6g0p531LuVAbv2AUoFj7NrK0JhWMsmNrcEWAKIyL0+qAJ
AvkMqAZmbidU3hFMkoVKsic8JVt3ooMQgXr1M+arF47ZOIWE7tTTnnc3mt1f2pxH
drNH079TU/oZ21hfzhBT2CW8k7dOL23iVO3rCg1b2ii8Ol4nh0uO0MLVRJjRhK2+
CpAraVZ30f/lOEPmjjY8JHN7inbRKQNA+EBca4UW5YrzB27UFwOUS6Uq/+VV9xVv
lNsLY8EnKvFoOnnQXST6rgfylnkhKEMQddXdy0sQnkI=
`protect END_PROTECTED
