`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K6bwr6Q4P28ssAEsOAAU0Ny8rUnp5yXYsmqZ3YYtvdH+w72+THr2DKzWieGKudQK
0XA/BrhDhZVHU+uDXw7R3VQMTF6hl8B2sgn4iOKjK7YowO5mgjYujkTlsXYitxT9
9pn4h087Evs2wPx1GDe/IndzqTuHMzcg+936HlOAFg3kKr9TOz8BWtldsxrKC4NW
cl2y3DnwLR6QulcpWyRWOfnZMvXiV+xVA0IAV+1Z3Hap9+4WtPD3FODnmktG4Mv4
jXyubOmYQev4VpTaswi8NOt88iglSXSOAGawC+Je6PlSepN2aUjR693pzcjAC46V
U730QufxfedfER9ZjyH2FQ==
`protect END_PROTECTED
