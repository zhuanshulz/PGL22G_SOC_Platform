`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ORHzMTaaOAD7mKOgLmrPIcpEYmawVeYp9CXctzQjPao4VCJxGU4jlJfTey0AWaJp
5iqouwq3rkpk5DXJTdFb7K8LG/5hF5zLwbmeioqHbqCZSOmgTvIsjK8LuPnEpCxZ
NwSC+oyha7t9Dv7glHxJ91uqg/6XQDMh8xbfWPdODhKT/7zJDqkxaat/64bikKy6
0f1Qs4MHZeezO41CUfNgZKLjXFYNRoLF2xw3AM8vVZIDjmmAqLaIznTzJEs7I+3H
ld92lEXKniThHsVgf7sjcwqSkbHWGc3m4+yv/o95jrBK5V9RFvWv7eCJdQYqTEt7
OFeEjb+ri+4O8Wma1t1kt5s1fykAXPsUDRE3MPUtshZ8TcF2Leu/W4VPG7Xky6tt
NrxbrgXg0e1Aakj15N+cQNmcjUCIdtuAUr6NrbEy1hXlUHkAKo8EyAB8chUZwnvj
PZrzCh9EMAhlMF2NcsgD2Wxk58JdYw3+8lXTnPe+Et4HWUZl3Jj2QaU494aSlXDu
UTPb7sPps1hb3tN6TsOYqK25Ui5JQLcdeDuOCNi8loWELM3p3HBLHlX8Tx8xHy3s
3uKUosn4+tZM7BU2CLHmsu1uFT1hCOf777imghCViVVsrstZH37F9yZiFq3fQFsn
hNkv9H9VJ6PcpXr3srgg2ZnzTXJUKOaM5ABfcMdGSLUOSB/yM+dOgPehIUdPuK5B
FccWiCX4Ca8LjmqJPqO/h6ftXi5p6c+D+L6w/QV6k+HUMT05M/WTCmZrlOvnrS+u
ik16as4TF4nRgCs4cVGMDvqxC6Ne8U42qHjVgNVbYx1gwqVldmezOgF4xkSpeHrq
AdF8r8q5Nabx/BvuJpteBWJXPz31FMi2ydtWWbmblNpZ9P1Ff+5RaaWBjNtC8MPR
VzXzzxF3SymcyfKqaDAZcJcOUBnqjTG8DzRTnfFczv39u/F5xj4mwQASkD4NIaFk
c1rsnaATBPm2+K4uMQ7SI+ZIaF8/yuChxy/Wl+w86XNRckwTVJGG+gKugwXDYLaT
LPxQynUB5v+Tbk24e4x9L5dlWLQOknWG84R2EauAM4XEQbdWlPTOEDgFqLzkF/2A
j9thAFaMMuBsaKJ8FkIgYIRImWHZWrSorkfYzQZ1pSRls+rYZoqNqrM4vElPXt7Z
PTwveQvqfLoEW38sfS3K1JUks8xDADuT3hIzF3TTZR9lmrb5bUBP5iss7qdkXkzE
ava7ejD+ZJSP0xSfQihydziIulf3trA4UXfrG7wp11VqMdl3vRJs9FXeOvRzEnvA
1AbWP7N/LoAh95eLG4bHXR9QeklPm+PvuIiz+BslmNbykh+bJBDEO7dfQLQwItl6
XrBugkJ6eNKNYSdPmZB+VM2FHU58hYQvquYpx/hSdf5qPPpyaHZj3lPsHEZGb0tb
swWxfdLbFFcKkkYACEhVqqnK/+tSuMcOImltrKZI6SIzZcfu45+uxVqEaND9JMft
cIGpAi7Syr1S9/EL6X6xLCKgS2NNWVttVLQPuDQno2BISkUjqzuzmLe6T3UzBX+o
mYENCD508PS4TuRWeeOPfhqMVR6tGN3Obqo9D0Y+0SEySY8Zv6nEM6q2PZrB8if2
C27pMtPy7/nfI4QegxrAT/5lADzhwDqdJoRJOjBTsRWXwjq67Mh1zzR7Odx/bcfg
GDXfFt+nZNF3/hZh7cqoQ7pGcj7AEEmySQqooZtOIx7wFXUT0NtD7hS4nWhQab02
OtRRWexc4LvLau3hWLd3isC5KXWkkhgw/K6QCTOXQV6kCMyjTyzShaDlcrzAU+Qf
DQTS/sXiKSPnAqsFoWu8XlBkkmdwbe2/y7lMraHhZl5/7WQDk/FGDGQix12Gg2Xr
cpwxhyHJ5ZOc47r35OOv6hAvU1SNG4yO4szEbqAtqX0qjsK/vDUc/yDvNhovWgAR
UaHld8WvsNLOrM7amhHRbSJbIKrtw1mwOxDGXS8WhocPXeXDLmTVQyiptAnKjzl0
UBaHVUsVTgmEGogE/3F8krYIQgvJyloL37p97aBdFAbCQHSFptENEAR2Byoh7SSC
Lq+8djJ4Ar+6+UOKdOvyKwBrnWNfEjYxodxA0IjA1uuqKxIYY7VXi0gqDgDixXDK
ipw+kzeAe/j2mPIZ+tm6AAkUlqgZb+rZGSjAHFTLTkwMC91CYKYxew7ybr8OKfqc
yNk0RsYCS+gIqHLLKY5Pm9I6yR+2TYlf+ZhFJQzVoFt4sCnIRssOFMhFaE+PSDoU
ukAmvEf4EyocxW/r1v/vMH5LTw6hYem1GahomfOzQHHUDSmf6YW1BzMxI+Ft3oKN
DbED6c1+MJ+7EGMXojlRfu8k4KaEiVrFBu5s+KUhGXLcsZ/+3YKDpRE5uFp2SjeN
vgDRl3L0OtHvht6SC+RPY48Rf/5g4ItiZqhF9Vs3sX+pbOXSfiMJhaKOkyaxdtIB
gT58dCZ50uHmVM0rkJDQxij9ZNF2dOehMGUCRoECeInlSWa/VfxXJqt2GVcUpNrB
RGCLrL1nyajE800/7LVMnuTWTYw0cdDXxWBvapukP/gnf+0DScKjtnU900WNp+9S
5ayrS2aX0CFwXO8yw70nZ2JBQxdNt4PSBpzBikwucFGPInVhCx29peuhROm5R19f
oxJfA/htltQNdQZXt9rpFSsVY6hPLh+KdeI762QWqbLe+/VvEBtmFIkZ2vbf1NXu
RBUBTHua4NyXqJvDRXUAoT4R6+0crgYniTSBSDRSpdU+KZdRb7px+FZdn/tt101H
5gYZz93SSEJBpUwyKlhMlqCMdJf1v4ZuEUQYfktyAjhamN4rRsmtxF9rU+9m0pSf
SJ2AvFpLIu6fl6jidAVFhJjwGcIguNKZTlyJr13W7jobnL1+c7fqQOMrlhWWc0b1
KBHo5yIMWQpv7bPh/F8BYihKFqRcayzUSM/j1ONhFJwjX6Qw8g9Ba/MJ2uVxT6Ap
jfXV1fIRlfvPaQAglPNS/X3D8+TLfEtIjc7vZOSJs0ifNQTJU+cj1krW2PdZ618P
EcVyWSmhQpOkI/yTf0lcuu1u9hNNed8hYjI35Yaoeh3tOa9lpjrGZ8hHeq8Qev6F
KRp67EGZuYIx0Kf0Rq7L/KddCyq/igWCKzA+lgzLVXehvzYZHBKMynHEi7bPjxYz
/DT3+EuzqvCB2W6CqnyidkDCPqro1bzjlvEDHlkrE8kAa+LEQXM/L89ELqCCFDmk
5y5R4PXZ/fA/63WZEcMLS6Ewym88LrtC/mKHCJ9lrLFEyBG5m1GgzBfH5gUxX+7z
CqrrdnEnLVNxeSK8LhVrG+C6CBMJzBq8nRRbtj1tzKCp1hbbNQI8rP5AN0hpzMpu
89y/o+HfoVd+CnrRNyD2+iaoLx+emuetvcByPQh9prPmTCQ5jgjjyUhLosYRTLbh
YvaFGcIo9besYEcqylJZTkN0TpRd8b59ZbQx+cMgFNAO2qxVgCoAsdSSD8mWb2Qs
9EAEM2EX1fOBuwYNtA+3OuZEu5uJCpgPdqt362qFdoO+nnQrjDu2ETY3QofWOeE+
958AXHcdgW3ukw+1CA3gPw31tHk1FypMkAo76lgipR74qTbhbpDu4Nn/U0reJdj9
E6yUu71hKfOvGtNmlvFahHZ2I/zyhGYsrGBDBKIYlnWHndTcm3sPaE37YoU4K6qo
S/c6P0qhm3tMhBn/NhJBuRlHIoGJuZ+vrmYftTj31VftgHSLLA35Yg0ncbAjnCMP
c0AtbJSXRWtUy7CoEFp4+tFOx/SNqFPi/8k720Ix8IPIryqqEJ7+jhKyNmMtXrtX
Ud+YQzeIs7v+a6lbCFY/TBzFNKcBgBXleRphfiKknKl7FZ94MTQ53kdLkMlDQ1eb
CzxkruCPZdTRRqChkrqKJTJBD1dLAINtgHKM/9Mpr/f1omMd6E+AFuPzcUazSwBm
wsvJmQtb1kVmxSOCf39JfKv+XTW/DLqmaRNGxqmYnklIqXSUrpwDCmT7CJGtNrsu
yNMfpl2/8i6/sCdEY+h4JP5QS/s0Zg+ofOV8xp+68WoEyMR92ULeyXRXZR5PpRzC
HE2JJJbH/iWtX7aSUI0XG+8asQ7Yrp1CzJpF/m15lGuOUUhXOleAPnL7ifJWenbf
DzClztObHUUwHREKzZAXiNYP5E9JIRnHo61BGu2OoTvIIVr+eLI6b0NrMXedduG4
l1NKsflWZ5HVEPPQ6msbNvEas9SqZTWhG/rF4PFWMJLyDISkncfIdG5ymcpHV4/K
E8vam3k/drHTmKQslPc63pp1SwHudQXYY6Ad33Ce3KS7rn91lmluoHjRUGAOKj+9
SH/8dQPaaU7910LNhAM3+oWDAxzX1Z8+rPMJIm0uVgcthtGsrG568y6dzs/b1QY8
wKeCwNpXmctZ0cvrZY96BjJFAsvkg/KP3OskgZYmZGALmRUYf0CuSydk2D/GjZ4c
R5AQo4cquSNiYs0wIaaIoAvyK5PhJs7Mk7ZXQsG8tOcUJl1kRXLZ59CYgFtikFm/
+/R6axYaA+q1tLCdeS6zbUE9RjxWSEVZ/GwlTSacFdht+a25hgRo85ndCqLKzEJM
rNIPyvSM5ej4vHR3+L2aRcYZEvU7JD+F/9FDxOCsZ1F/EQvPNBagNig6mHesjQte
oxdrbvzKK3MNaWwXONWbjGlhN34c7Am3RL21pP15qiw=
`protect END_PROTECTED
