`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f2VAYy/+oeCWchUDdIPJAnKAB56fdq2L8/oguqVgZqkLznfloGIhGRCu6v7tpA4u
54mLVrz6ReyJ9HhSutAE48HWqK4P9VVrG9sCYhHiZ0Fu7vL/RFKvGsYDZb+CaVth
Rmu7Vn/vt2/C6gbulxgtRwScoZKh8wx/g/eqtfQNe51LGbwF7B98rjVaUd49GDOn
ewHYeCPFFfdi9hD8A0WBoaSuFVZVRV8h6cpW5qiuG333bSJF++7tRl15uNQ27sDw
NfNXu9Lg+Zu47GTHGgVih388Zw8TvrMPqZci0eiDyEc+V5lSo6CTbX4NVfZmu41O
GtPq074pmyxKMLGCvitCn77yS7Mpu2BbEiLFmK2+5Eyuk6DcaeTPQU8HvIHeho/5
9yVsbqBlnCM5z9OV4M413r7TIQ1aFOgeS/lNFS9x1LfsAtYhoYFTIRJYs43elXUs
G25MiZCZruxMxzQHsPSlvf/9XA4r9ES77B4nIPiVW5n20E+MHNKQoXpJGfn4udGo
4ZDFJAPUh5CeR4LEPxDy7w==
`protect END_PROTECTED
