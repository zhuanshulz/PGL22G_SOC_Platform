`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KdIs4udGxWlB1qtZydQOIFmzqDPw9kcmE91be19LD1ojAyzj8u+4CbfKeeUpT3N4
g+0h2s9Uy0uLnk5UdF1o8rpuDBFXfmM9mMrtR7BsIm9DKtZuiPeJBs6JfjvjL1BI
ZnP7TmTpwFoyQBlPi4IJ/RI9C28Asf7HEtMPHKteJd5syTxlQvuui5boYgHGTugX
Ylbg/QRIBxBtGRlmBGdtEEec5riCHSVa5iQVmu1Gn2HsfXMyYpLUcD62aYZtdJm3
CIWp4r2UxApDCk5LO/VEqkc/QDqiejf6VZ2MTC8vA/h8AiTOQCBkQN108EerCaOf
Wd9v+oqvG8ZnWg9i7DO3Ddv/mHJ9pw9qeJ9JiWfOJa+b0NMhNhgGczmIxxo5hDtZ
7Vy6+noaAogPZ4cgSgGK7PZ/O4RlR2PYtOP6LpAcijgqF4emNbXkmSRmVZJ0HA0n
klPR2ONFha2BSl2nQu/2oL0bFdVgk5m6Z/Ixl+KiCC6CKebUgNrm9liOWp/pRmTd
`protect END_PROTECTED
