`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TQMZ7bFreiAIpvCeN+JMXB2Y7Ia8wzsJsfg5Yt7YD6u0SPVWtdeRJOWtjLzkwXbB
1StLDxm4bmu7qBuvcmpRp6/3SCoPeFKCnA9Apdh70Mf33OD5aKLnjeCp9U54hvkS
HNzdRfh1Y/ysmqVrXm3DezvgJENEP8AyCJSQ34YNQ0XpsVDH1hZmvnMZe6fs948h
hV7eGSwBLMBWpvV5zWKKF7Z6/4i0GU496Urs43PI+lwGFvEJB8F4bDuu9bGonFfC
RFp3wtPoIBMaFt1CQsii4Q==
`protect END_PROTECTED
