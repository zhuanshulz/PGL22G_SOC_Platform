`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E9zQdoynkOlVIRLITN2DwUcyimVDEC25JgUAyJ27CNsQa+P4CiadpFIx0LdqIO+I
c0cg0mRGlwLg+FotpoJNFHpliXrHnbAPGV0Ufno+NXmlFOYK8Ti14+XN6xGIck9w
MtzM0ejokRq5uX/jh/uWGARkbq0aFc2DdA4dPTwIJjiSVK5EvhTmvRC2WyAb7V9a
LD9ROWVStP6Av/EmPyiRg6pVFIHNf64Iaexs/41VVYi42wsAm0JGlfG7COlVldD+
qCx/PMrsxqBdLSGYZ6K1OJju/TlMSalX5A5R5syurYg9XvBJZvlz9OTWpdKxIG51
p00mcjeUnpg6UF7URZ0E0Y9ANa4HdwQH3c2RJJ+SvcRq5Wn8IakStc8Bmmt68wIC
I0LlFR4ynn8wt9U1EaLy4gzkCK6MEKJLg1M0uHMWyBqIlqU96TpHM+2yQtN+R+Ye
4Kyy3ROPKmNVqrHWrr/8kyn+a6D4LRf82kvr6NC9ey9xwZIELga9z2koz62jj2Ax
ucU8XNL0tXin4hT8zPpkLHTqVsRmpbZSaixMrs4AP6lRXiyevp4Fq41TFx3ctUmT
JA8SR6niyXrSpRGN1SGFjYvCMo8zwYMTCbUkWNpvoOziXNA6Ghs/5IC700V15PzE
bIZTdeSIKbMndH00SaHw0DbOTAeZFhBx5qUuNXswzEpywBJPHr6Gbh9eULM4SpQk
9TB7e1AJJfaPJdcdJINigFejiJe3h5kz1vQtWIuCKMrvtPt7KBjhsXysFUMATw92
gLqQt8dAa4qxvkiBaqZrE2Le34nQwTNV2ZPYuDv4sEySo9HT8n6+AqhRRH29VwUf
z3X2UL9t9dWZ0QFSN9GOx6g62uoBOTK5kAMjwTNRBDGlcTuGd3q51tE8Av+NmwQq
2pjMd3IH0ILFTnYj9CGcLLkBypAKKfCTXjy3bvoonWUpAyjKyEF2Y3NG+tQMb6iy
wNGwnZvSbJGAKLjC8osKMgLbGW6rSZovPNUzOJa2tOcBDL4xIcryphUuN5UXG1Kt
WON5ojB2tnwYtN4wRLMVnJvgPVCBIdhwJ3sOgxUzKKILRcOUBg9KvfUwPJTkJ+9y
mKNxqlEaeQWKQujUpOhzGhj8Y+30Bh3+m4PWzwR3r4ri6089DTzuupTejSXg+Xl1
GTGGaLbKv52X7buI2Uyv1eMzGTrUe2yr9XDXz2DBIXIsaWdgHHTjMvgjPZzx/tjK
SnJK5xW/xJs1mHVAZrlLhw==
`protect END_PROTECTED
