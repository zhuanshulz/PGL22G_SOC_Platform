`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SY9p/G3odKE68nUEr5+daJCj19TC5KTJgWfjIAVR/R0xfeLlGsu2fYnE9E2CHNmm
xqnXIDsnJuMImV01+VNycPd1JEoA2lD5GpNk+YNq6lS+uXjavqd2Gxpr5dYyEfMA
ZI/cYyD+oQkY9VeOG2QCAvfmwUJAQYIIpSqhWvmGZeGSTLPw1QrDGMY+x2lbLddT
Fh3aokY4+px2ys+A2K/joq+Qnudy0fQv8qvQeAfzZMen5ZOgQcnk62YIsp7ZCw+F
9MnTI8LjxloOmwHwRIQohHMlZVFhroJtGN9VrP44DBTntLnESZr8s2s/lOqyATtS
IIvCmgTVnWJmrnk/S762xodhugS2o+PiqrcUt4Z/fRcc11kFGzVW6wOl8NbsPMKf
HV7DJmVQ7R4vv805KyyPZTCCWHZo2yFLYia0V9dzNVIr60g6qP5ck74YSoGfSLIL
RXBlxOcw5rpzH2VfW3T2eaabVqg+6/AMkO+xH1S05aot/57esy2DqXws7fgVEq09
YR/uu7j3RNIU+txa85iLcw1h2YGdGy1AL723zgGUUhD+uCOYuuwBobyCcvlzkoou
NkQuiseH6fw+IYyly4MN08YPO2b948d+kVWTWAo8x3lLyrWKQAS1NpUs9OfSQ4QO
A8Q+kM7fi5tckkMQfR/oCBcTwLKcqrO9mnR2v4QgRim1LW7DAja2+SAffRwGe3dk
6hHKkHIbl8rrySZKgpJpYA==
`protect END_PROTECTED
