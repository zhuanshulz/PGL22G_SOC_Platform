`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hrY6WhGFjh76ccuYjP5869llMlE263OHVaOAAn/RD/66E7FNUE8rqSeYlCBbqWQ7
xRPqmxrWS+Eows5w91mvbpIU2PsSFDLZ7R/8vL5agM1THhCoRVFBqwPCRr+y+ZuT
Vx/y36qDux5+8nTX0nKZkTxET+6uF+TmFnjXuE8ZgesexXGUTQAPFp7VCH1Xy4zc
ZusywVXjyHQQv+rmWlNB/LCT71FguhOoBwYh62NhLKeZNh+QBLy3tGNrm5FB8lj6
TnOFXllJ6LWXm3TjjsFdvQ1RFHWx2kvDkx91fk1gqS06sPe4r5rMJvgAYtzUZRrj
slg5vIhMfGdPryJQVmzKNZa0pa2Q/b/2Es942fTqpE2Wve19JAngNe3kEjTGy3Bo
HwmMlW5uS0GBxTs83P5YwE0BNKR9fVkp42CwQZqlfIrDVd9RxO4M8W4spok3Vx5C
e4FVImeUt675Equ46qAIPQUCLlms/oe/uWiwJ+hy7PTbwgQcJH9Mz7vhrrd7jfwz
hKQJG0FKQjnt6nGNOvdPY6nKjJuyJkKr3eqR4a2Kk92+TY6UvQiMOKGk0632+S5d
ocVUy75ckWfp8ZRcbpcgEg==
`protect END_PROTECTED
