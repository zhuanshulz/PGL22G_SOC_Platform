`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u1O6XkVjWpW9oL2VEeYakqWlob+AjWlkrNRfjsoVc7tzGvB8L5oRPaLDuJ+QyVgb
ZUTygzT3akfg40U+tMNPbuPMdlIczK48oM6kbbwCl2BRTheBF1iiW24uG6XtYZ3H
tnX7g5yLB5SzVWsEwhW4asF/+qhzBTLmrnACVc1tcBGYg2ZfhScOm5AIv1PD9SGW
Ze5OjqeZ0nuMVg3eYvN4pmT2LY1T7draK1JSryei1As3kN75CS3ucvzkhnNM9GTi
wwA8BA0fEwK1XpF87T8HzO2/LIfDvr9mrX/5i9SGWgvDcLTbN3Zrj5xEclOY/gk5
hwAtMY27HvnV5MfyCqTANT5PQkHDF/QhYZJe17b02Ra+Zf0ON5hUoCPPjNvC4SF+
2HqWUhaO/XRc3AMNf+Ko++B9AXoiVoe/+rT1qvaMzTdRoy9dJ3/pnTWhAb+bY3Lb
`protect END_PROTECTED
