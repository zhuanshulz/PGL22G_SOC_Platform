`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P4dNboJAMWk0hAeb4As+ChVjUw7k2iIwLn5xkbQcffoeG2HrvvS5ZWiRhhmWMA8f
p47w7HTfglpb2ttlfY856OoXv+uqurbuPniKpzL4LRSZMYpyrKrcAtbl/UXa/VC+
I9NDnP+jn0ShokFuMfD1X0UxPzLOBMsqt99lzvJVNFwlYI/5FhtjArP46xp/I4IS
Dfsx79Vu8EbSbymW7R+GCJKcmFxrxKuzUomCngy5EHstelKsH993W7CWZy8Blz5r
nC1NpGzaPx0QIymyz4/p0t37dBWuPPXhlUmQU8+xdEEjYHoL4qtPvvy+gXtMHBrJ
i+HF31LrXJwzmn+IAJBgKDGXbb0nx84F0/BMGlCQItkj5efsOvVOXz7BlF9fwY3U
TaB3pjTc2WYMKw+H/t1dZ9IjASVkyekRlcmQ8XHTIhNWdvNhrDGBzleru5+sqoer
fTPLIEbXa3YjXRAOJORFtzYxPJt/N45sDzo1Ay7Wlr4FTMENM62uIBdnqWtuOpIY
2v/3xG2cVPirOX19aygyYyrMz+HY7eAb+lJHfVOeH1bwvu3iIJQtvMqe1CodZ8K1
izhPuQQ8wNSNLWsnoS2IlR8KhmLKoLMd1c7sS9Wvr4SFVqJrCPTPJqE/R7LlUCA2
lH3tPN2Ps3hejRVdP8HD4YeHxDPSZT6F0A3BVUjJha0hMTYn1WArJoeC2tCU0bd0
U7ZiIMo6vBlSXpI+fYZ188TwCeVc2/WgVkmbPQ3UvKx4qTG4DzU4Jn3ePVYZ4IRR
LJxJfTucAUUegW9BbfulEDLpZxE6tMd8SJOiS08zbYrsyE8wUgAQrJNxEtTRtX2I
FFYNeHFP+Zmfmr9/4aDNIwxKbosw1rdNoYeHDfJj5tDlDHx70iXyED3TNH1Lec7g
vxjRjWVqNfV+20wJch+kZL5Q/RH2L4j2MicaYU6SdhqAU2oFDRzHah39vg5CwjBh
Ld5BRRJ78yJvceizAcXiR04uCnT/XDzje+R+tqGPzWo=
`protect END_PROTECTED
