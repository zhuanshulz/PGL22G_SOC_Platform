`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fyZLIygl8cB8xWiMkXqTuEzaKHExXe73O35bkXpaRmaoxggPeToX0bzuzp5stxeu
wG2Ot19jjC3hAZIzPrpmQycz5930R+Mmxq2D/BeatCOGn3oIkGoGW/Nn1mWkj3At
fZRrbCHjEWxZNUvmksYWA7c397KW/1YjJfn7v3RuG7wf1W+fMmgK8fV9me/eewZF
TJlRFf/EQymXwyOdKKtBDC5Zxwo4nN/Lho+xxsDk029mJ8GkTa2ksZ8Ju58yHDmY
TwQmBm11wiR5CEejLenewKjpAXQckAN3Q52/iVKhtPSmpcFyy7rTsKXFeeOAMtZB
yYk4abrAGoTDSkwQWzDza9XRLdN7lRp2abmn8Jj/z4emWzZZ6hC2TYhEeg7KcGlL
BY6jKN+t3KNgtk0VWSrHTePwZwQ/YLmGxN3tjm1VSUZtPHpDS5bepHwDVBE2M3B/
E1DbiQbhOzMu6jUf9shPWmGOk/bxVTNTfsgocLLe+LBHpAPmWJwRmmPSiU8fJYaN
zctaszfpYf3ujIs3dB5YbnpBEjnkxyR67YkkfWBVtuJ/vP7jFbBXJx0whjfsoavX
Pvn/2vtOcpbkMdo8Ucdis35HE12uOML86xaJUhZcYayPDwJ1R32OLnnfkNbzJSb0
dVUA0FcrhclJn7977XT8CGvdCwQ0Gkep2dard2CpnHg7naYu2w8kjMn56+YtLpv1
qdMzYTzSBqFIfZSq/HCryBLIuaoJpXfrLzfLbls2eJKAM2itHSKxGe/KGVCKapcS
6Cq01RHY3GnMi2jc/V1ylehOoTZsVy7r1uAkX5MfYEN87/NGdScVDkgRD6UzrJpU
e5htb3x9tMKGjInM4kqG851pWwM6sR8CyEKxchKpqP8vSoZwrpJ+Q8/FOxylTNij
rYIbvXrTkXsOGqGl+cpUWFgnnB6FNYY4v5c/zChR51SW5C1reMpuyQO4zaZ6GB5J
+xrO8i4K0mt6qc8XCS6YcWqnddxdlQCJbjZu6iBXncUuffnp5uUsmj4Q7R7gQoBH
VAJcABP6P2ig05Hj1qzrzC6cBTtsuSKoGhEMQYYGeDGd51pwQAJKuGhn1k0vR0eX
tfppx3p3tGfnZUv19SACfxPXVcePPCKgrEmc7YnywvjUAbWJts8rIibsF3H7n8l9
dPSW/YJ6BCN8Q1Jd+LLFXgzH3blbA6S86RvPBfy2LddSapeoqUX2YKSCOlklwS7q
KMNxHKfAPATUzgPcoS2vvuhcpltvRpJKRMr4w0Gpoal74mYWr88Aa5S70uvJ4lDa
JkUfMwa4JPm9FIUdVm74SHFSKYEMTNorcZyP5HoqPnRQbOeB6orOzBgVqMPuLkMs
W5zJ26ShcarzECVDhM+bJkap02e7Gs5udZtWt/OgI7s6c2Od7AOOBJ/fV0nG5K2y
TcrquaI2Nf/1EdW76zNbw5R9NnTWmjhEWLtIU6M2V5hmS6z3UROzgTQ0WL3FGutq
pCBgeWHg6y2IlYpJiKDRwDRdTCrr3zhL1mrVQ76odby5bV3j0dwMU2cdPVFKxHKv
MyvQ85SA0+IT2N0fmJfDU2eaMcSQcaRnmlW3deGw2kcA6x3XpcbWbZGW+Ku/Ejdp
w8WudF0fY9fj0IUOsCej7CoWRN1i9w0eCza5plfof4uAlxFXLdILEheJQT+632F8
/LJnJAQfsPHb8yzrdZoJypBWJ7i9QWV7Bvjo7gjJ0JqvISyABozM5bnhoZgAyEPt
IS9isxs9YZe8b/5Wy2l2pfWIi4Ct9yFQOqPoR870/yyhhu8E68heP9yTu6ar3pDA
vhCpvqMUTjg9vJ2ulSJzrCGyamLdcX8ApEhV+yG7zrfWxGJVuJuCNX6WKUw3YZMX
UtrZwLjO6TXloEGECK7Aoe808PSXGc50af1k5zY4WtqehFTPq/2/lgAC/YzkXnZF
6PBvKkdOP03yYTES2PrEABJIaMvGloFuc34FV2kSRb5UdGhvTwpXP1y86y2Heo74
dM8Hy+o9U9LKQpmBAcItgHuqWXrV9zt23C09eaBYswpEm+fo3XcUxe9ELoOdjk7h
yvOp9Pjkn/hXLagakS756AHeXPl5sOrkLEE2GUei7rOM5ItZWvmtNIji9SH2v5+T
XzaiNFGswJZjmFwByD/YyxVrOYatH3w5lWMuwqvTI6tw2YkPVWPH3HqN5rtREfxV
i7j9aMBQtRBbabO9XT5wtg==
`protect END_PROTECTED
