`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8YqeBNpNga7PNNSxWTreih4+gYYdEoxF3UDCc20TYlK3F4JQMuJtQJ+rmy8JuUBG
2mBT0DXwKcci+wuVi3M9YMfO+jpWN2TXGzpVuCB0Lt1a7mzmtmhXz/bPbjZl95Rl
57ehoJcL5xkZcUal01MTgL8ZyzX3NURYAzZ0ulcWpj6mO16S5UE9aTNR5smoJDj0
PDKG+uSO3V3+Ttigr1zn2TzC0EnG1bORPUr7r+zA3xI1sWLfRCh3AllTkkTAIrjT
Qs84+4Wh9jewIL6M1U/up2MJxxRckn0WnPTU2UVFrrY3OyRLWuKEji3KkSN8WPrE
srQ5URWQkW5ViOT0jX3WSQskMTirJcYlhcydGtTqa6Dx4a3JwfksXcrBEdbN8Glm
KZ9SLDLV/Z6Tyag8mtDvLtQ5rDVKQnYLqQX2pJMW1BhxM+bVYqM5pHnlBoW0N7Cu
Z3ZwKJbre9e1O1Q6indzbqronAGL5ANatEQJaO9aIlpwO68LqPfELspWYCdGtdCz
p+Z46ZugEjTKV1MF9hVtrGZBwlAckmRB40F4kSLhoj5Suw5PfXC+VV5nYfvGbriI
UBLw9LNy/xLv1bmQXVAI/r3Ukk/ufnr1fwXh2Ixjth+iXE2xCDwUUa/J0P/V6waj
CzvCN0tS8zZ9sR3iy63wbxAt7fGfrCj55rbKGha1RRTV8NSPwy2LlrcQaaThrIMF
umErFtL+W/3cZ7tNvh/v8zl/XyLrUrcmXSGNHKnWs5T04z4BX7k8roMCyp4XYDGL
yoTxQmaP/rYRDof+1AiVSFN4igTYzcWJziRK8OEac288ILLHH7X2ugAnwiiK5gDA
cMtejx74jtS6vZjRJW1jS01JU6RrSu7oyqXgRNOQMszYkoM5JaghXmv3nyt3ELMz
vMXCci3UmQLRav8ey+uf+dmVNu5AtdKmegLfF0uP0eQ7gbKp2S9q86BglDJ0uDsn
Z4/A+uoR4Ye54nWO5c1sR3fcULJo786v9unvwfOwx14=
`protect END_PROTECTED
