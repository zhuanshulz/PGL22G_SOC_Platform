`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5SR9MEA0rFHpel1k6wZupOPMos8L2u92oC5PQEQy+iye+dP7aBrWmevkFC5o8pR7
q9+b8XNPqeN2yKQZ85Gn9ZGUL9ami/Fb1Mg4y0V/lx7vudy0cAs+jKbKbhuNLY3I
Tn632VGhmQTY5g60GMFwFRLhEA8aruq6kfd6j12KXHbSfQCD7wGye+TqAdORWxRI
Pokbv5uH6p2glZJ5pZfbWmA+sLSoOHaDp1VsK2Kt/MC1VAYyNNiNPP1zF68tdYNJ
ETnjqhYI++wCvlX9HrdK0UOLrCOkyHJHdB/zyJetgYvD1AsvDvKMeqN9fxmYABHi
IsqqLu0eSR4w62d6qf2FjsFdIsKbQk6CTWEjwP4wAHnCArgMckky7iy0pcrN9kwY
NiaxBoG7JO0ILbFw63yuEY8QMipg8P/CzJikoeRi8jIgOCxtynKUhN9YW0byRHkI
2QqAhBc+pwL6cZoS+PLKOFAZiX0N/7LBAm3fdLJvOHMFnjVKvDEEcDB1e2CI61CZ
+6cAqEnbuSncDq/KLCcYU9sT4lWneZ7iiAw+WbNIyeZPQy4Q5EiCku/cJHaUsB6h
FDodZCndeRhGztktCiz72s3PAY8rF3Tx/JI3qRnW6mVdgNefjkXWNsAlhvocwNIQ
WK6DkJ7QDpwESt7ROn4+PlNsR12ACS11ZO7UXwBa1og/F20NCA7z/0X7vI2qfN7n
GYCj1x3o8cebf2fJRPB87ao2GhzWDcLv+GcnseJEXAm+6OAEv9KCPeEtu97vkydv
Z0cIkvp9hPUIJHFKjgkZfzF8ZivJBAQBXqm+PVtcCgNNF/udByGKn6RQcEX9JuWs
bFIvk7FlnibMZRepNOyymi10tOfRbg282kXGrC/ko6FzTFxoKQbJ7Rngo1q9ObXi
WrVctpkRDqdX/9svT8c8KG+0oYQiRm+8XF7srIwRxv2uHbW1z8UVf0EKw+nWXvRM
6hE1s3qThuvtEEhX5vNLGMUTF0VkiwdodQ0IWnAP0tAj1DiWqneCXlCajKjhTcFc
tZy08TyDWCZo4mBC3hncblGLMO9ANPlCwxh8zUwyeNaRr0lcTLYTYTNL3/GENvkO
lqsibXNsUuEipqRdhxXTHtjOcgrpKgJblWcU0h2X6UXdN66QGgTybTyVr4eXk0Yy
5tZPAj1u9Sm4ob0M467ftRR4BNNzJAe8/nxSfmfNR+/iZKtzJBRu6RiyFyuLUVKh
hLtNF9noKfvs6ysjHWJwm36jpoLrlgAgizNdWdAZraHvP2BH1+RIBZWStv16Xpvv
xFyTLp+VMZgRo+vyzKjQeF1nNkF0oBfvxr5UInwXn3mzQhpt+6iNwyXhNjjahpAg
Z+yFH2aLvHuLe6OEY1i8LV3fpmqAmO70vn6NmXw0DYpd5Jqsj2TVv7W9Mw8UPKPf
yyKqtVhBcifwI29y6P6fNYn7sRY6XuU9KZWKOsOwicIBcVlQlHDN3woGNGGX07e7
43L5HaOf+BZRPWHXoTawHaCp8MntrR2xJzCBDwWl9p4/RHwlQfieyOrjjgGKMhdU
2D5LYfWo1m1PQE2TBm9lQEQ4rtv8p6g6XypqyGC1KocEPHSq9VPyibL2JKOVwzt/
B5ghT028SXO16QXv/FMaTZzm643TESgvGSeTWBs5Lo+8voChMD5tyGr/aCMqAvDi
jEzrSw1UCifWQJEdxToxGl9zHxXHYNzkjscr3UO3KXflSIYln1EzR/k1p9X0t2cu
wm36fVBa3uY8jWo8TbKed51cb+y7pn+4qZJdFdOzu90x9JUZWq9e+iOTjhIdMmzO
5IgplOxzfpPA1uEZrR8G5lg8W29OUdMfmf63Mm8G8zY3zcqOSZkfdyv5OfRvt688
he5bdwS9o9NT1ahiSEk+9kqr5+QQglKBFsdTWjfyetqrrbPCyn+karOHlhh9u3cD
FBhXVLzHekkafX23ME8GtmvpKS+RSajRTa7mY5CcufHSnf7o0qGn7pqtU8ww3L0D
/0LXrqDsxoLF6VRwtOG2fQgDN9bU0APt/z7+x/GW7fUfSsojn/HWwq/9FmAtCuxY
eM4BYdfbijKDO931cQv+Nhj8HMcAcqx6m3YW8jnNM3RgXqEJ187cLH/jMHQ6eN0n
9jbRA16i0XK1qPqWFiMJSjyEzP0XhCb1QVuXV71/A25QFyGdgTCLQ85gbDp5o/qH
XUlj1xZrFaxncsqviBVkVo+B3r/iW3hiLKP51mFpzUT/qdtKI14Ld5LuoZuIeisx
SaE2buVWQKx5cY9qjh0U69a/nHFIC5cC9NuxJOsakJNaygVi/gfV49CklDHTOC2T
hstpllLKQo/okG6f5YyDnmujThXfl3a1r7xryuGZvqbDgwIdEQpx6fO93FiXkpl1
wQwTkB58e8IUgNgul7BeQt5IMB60pcQVT4udTNA1K2sg2xv7klHOrXyO2wNCHbfH
hyQLhkWgwbcNj0a8IsH3vCpYfM2dzh95YXo2HfPhuU/rQ+3az8pM1fBIfS9Qib64
lN0Pbw2OEQ5kzZjqe+QC3/fseZrc4s50pMh3H6h4oqSI9BfQULuchZ2sqX8u1DE9
u2qqwub0FTO4KiqLA0d+DD3SnJeTT7TJdOyMt3ZAmjRHBnlJ0vnjmyKgp3AEeX8F
Ao6EYMPHACKf6V7GT38KEa+ZTdek1moGvKDKFERH37EKPA1v4ZYan5elXfzk1GKG
jQ/+wwT4F+FuL6ISFwnrjoAKTd3lpBI5IRDgH24ueSq0wMlp0iWIyvrzAtRnzGRu
UtZ+r6R5P04mtYjXWQQvFtnaUQbtoHa7toHr/UJVPIeHGh0ptmte1P/2jZF75CZS
1dPov2I9oqn0pABgykZYRiP1yz6Q5cKDq6OkZu47z1jkAW2t0vlWtiAW+mTY/jCU
YOlsSE4oHF/xQH4q5IzLP9+qdIwUnK0xv9p9IpqQgi26B5eGit0eSI+f22sKGm7t
qBH2KoB54M4QN2TJidPun7xZWgI5lMskWgc6sTLQnrBB+6ZAGh9KUkR9E70CoPlq
cBn9zcXG0BNUbGLh8Ou2Yb8jWB5Hl8RJqA9m03024IgdNOikWT+MNUGmjwy+5R7X
izbqB2UzH4XjqMfo5mRy7rDc/6ix1QJUT+cjlA6IIQqeHltL3TgU21ie8NYu8hou
havTwv+eXPgrmkh30hZoxzIVLtqMmYgl4ZrR4xGy/GKq/4JrC8kz2ZXkccjbmgxz
`protect END_PROTECTED
