`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nu/7juLHyAVep8ElPkK0XG24lUYf7hM5xjJsufTbCeGjImppXYFGyo4QpFBXu4ht
e63qSdQBW2Qq9cR+lucXQBXJxZTbeGbDcy6bPwO76A8EP0nhvv3o0i02syNI2C13
QEWYInyxyrX8yfjcYAvJIAChtILpPlUX4aKJofQ9WXkDt/cI02wexT+CeVTUaYY3
5D4SB0eFVSvMFACesgRZxPhFYxhXmLgADPgTwfiFkIWBqIXhNykDfyoy9xLhDlLb
BGGv38ih4YeNuHVtrhlMOOULKgdNQnFQe4pSP9XiBHxirRC8NdykVZJ+3+IYB8kK
+B0/WN1gqJz9A+oh+t3qoxN9KRIZBB7yKeUQ5UCZ1j/YefPwQWf0mln5c9K0GoAN
NjHTMR1uSS1/HLRjkKHbGAz4AeFGsg8JTyv7AVKKItrpuGcoMkRfQNN1afTW64Vs
oEi8BAbUgiF/eB3qHEfck2a8AjGAhDYIYA1eckWqgSHJk7EPcOtlm9F8dlpPmH/X
zgYQjbbYl1/3E0IoclIWOqGq+3VzJOuAJiG7ooaC+Z3xtbiOAR0R84fTOzq5OfEg
KJ18nFgoGMJ2xLXM4moltwxG9cZ/YtoppWZ0mnuhFxYb7c4QsD59Ar6jsDRrnhAI
ZB8NPwOszZfsETMMVtiHVzHXcM/XXfh6MxJ3XrcedqBkeJAZ2Lq8Ac6ZAJCrOEl0
Y6dhY2nJ0UCZv0AyT33K8KlqudJrewt1uxiU1Qm9t8MsXnHIlDrcu7K9e5k2sxQ8
5DGvJhsliG+H6lDeS+fBSwDZk2Y34FuUgIE8NJvfCwVoHYAxeu4pF1lOMSJCDelT
y6Ryz2vgJvvxAqYvWNUQCzhXLgn+xcCtOYXeey1WEHPkMC8V8ks4jgJPNarzAmaR
Cw8Fpo+gtqdfajaq6GBbsBTymrxBN0r+iUceL//3nO6MfDQTX+CeoyVKniWNCZZb
inSv6shtPeuQaMZHd/0IbWEz6L3K3Z2o8JMIn1uE11b8rmzuUoiduZEtCpG4bdsE
tbwktr27nxK3Fl7EaTLmt9M+CQ0GKra+PN55gwl+W3gvMxXcaAot8wHnKoZ/n20P
1569K3IINvkichJ6F/5SGZhNdprK+oGLoH8fysmzJ+ADiz1x0FunNsLyQYdgXbeb
I+j8vlH+Y8YrIa53+ZeH2yOGhIFn2zxEoiCTkxw0oVGfxTchq7hurVDkDrzRb5YZ
aeR45YOulyfUV2NF09iOAErVLYSrj5Nf1SzPcPZF7JqSbSxKngk8pKgzGmrDSsUQ
znhxWhDslGqxFohICfmFnSu+BQL99zIo+E1PHB8L0XvdglAM2akgAvfUbcUuAhcv
voDjXDd6hcg5KAyFSePGNRnDX4OPZY3iWXRNChBsRV0auZMXDLCh0Q+dr+wE8vgv
q/OeTr5FEzKGTQiGhGbs7uYIh2CA6ta2HXK0hG18Y06GCc+uNlzV1b1yGTtoyUWe
J0LiAZjbAICQFTAmmulsiSfkXFyhMx1TBRzIHCChNm//Qn8qCqWPyoKJxOYx5knQ
KxVipJS7JT8tK3VC5fEuWdXnr91K+VPQNlOzY+UqlXjvGiOE4Any/MutVMI7/LGP
vJ9M8GbSRUEg6NQ4zUOeXrZj+u1qIFwRulLEVYS0FY2lLXr0Hpi5zO+jGGR53phO
DgT8rjlknqSMsc4/tTh3cuXIJ7uYWhKa/tqNOEzKl0EFTX0SgKvtDxf50g8mEJgd
xxeg49fCIf/BGK3pMAJV5K0CiOMby09eVhxTDbNV8YoXZiMzJCRS9LWIJKDfU+EK
wjSMwcxmrrpKCx+ZMym/3uEWLrq9L3wgpVWSQYqb7RW0ten+c7GilJbu03XMrylp
Dvv4Op2NluE9f07yIN6kYgpNkjEn2mmOY+itc+7lsb1KeYLv4GRytV7CvZh18rsC
B/RY5Fj68XavvqbctY88Ds6N7ydsROUuKYDDTqLBQBQqeOBGY7lAwa97dbhfevFx
cJJDESlEJgiXuQkrSCL/WDQNAuWtv4rTsKG8M4l8BmimDFFQPOTleLb3weIbsBOW
KW9ggQ5xGnR5ap5YDU7BzToWW62omPncz4NPdWhStjleqaMjDeSuoKzVFz3jQUtr
awh41lclkxDJTaiXolJ42F1swZnb4WOYhkR30hhBxYxEMUnBMHgJA9MPATyXGTCG
U6uq3TxyfCv35oRdM7Fkw8wXUdlyCPZKJgy9oZTh2pYqWBkfOKI3khpirwSiaXN3
WFlzur8c1b/5ccYDV25fG5pnEtJdqQ1dIrX2tjLWbPAweqOVplpu+MWe5hYfL+F0
03235sLc1CzD5qCGZ1bRTv7Mbd+MXuoXZdXOfe0sXad8g3kG1XGcYSsqo5/w+FN5
QoR/zA+TDRRXzAOFgPjQSaEudmvCKC9oqLu+JnnMkt2m9z9Lrux4UVwdbuN5Ll2b
j1+BTJi+Ow6bKGDO9kup6r1OpbZODb3ekM7rSxrcVxqPNnVcP+++3JEImVyCh27U
QD56cikh/7hm9X7xfOOXc9y3RbHr80Djm8C+E4v/3I+2VhAHFUDpT1ueqb+mYvJ2
YdZSicq8TWQKK9ZoIvp4kzReaUN+uZWXyqOiKtam09PYyLMS1T0RDw7xtGJay02a
UHRayY5cBCltoADgdEYIGE3KVJjYp/pSOC9xo6ybNJnMELg9SGZ0xIsux7DMrNes
xXFnhiXMUnEND0JJDSnJGNWktbjS9XtxBXnli6p4kFLU97CjTOxV9eLSgw4WbSOD
QfuNtQqSmzowIeclwS2JrBtFhHqRTDu2Ouk8o7nZzY6WvSASQ5STmUhSb1DhKD3p
ZHUSOa6gsuRU9Sk3XqpH2GveQ14umrzkSU+ciXLz9fMXpXkiRmqS9tgG75jXp18T
uEhnI0Bd4+kp6s0ZJLyuMZ4jc5uJr66dxJvjVTpSYR/SyZZcaM3v+TB+IeDRK6TV
v1ZlBR7fYrSpsTbSLMKILKeH5d2qgEiTaOIcF3MG7Nc3pPojYByhNvg8C3Cjj0+l
CNYY0ht3WvfqfTpmy3MH5/kW3yizCvz4jli0T2+5MUFk4y6+goLwLhP18+olc37N
sFqrk5Wu9DQM2TdCcbCtWD20YoV1x8gMmSOn7ylUGYgwawRd9vQU7qL/eHg3Mgia
eFI4ldXnncqOJDTKVBFb7l4fO3J4RN0cSWQ80V4u4hILko6tVeP5QtxKP7kM95/Q
9Ic+K14aAVO9kPVSwWEhbspET6dIFhWRhD0yrvXZ/aKTBjaFblGegni8wBsPZxns
aD3pUlAcuJ0NstnpKa0pGYtzu4Oo2IAmf7XYiw6XdD4XpSczY86dlgmBtJnNXo+v
9F5vGxiepTSOKpDlgBQadQ80Kb6FepnCIhbFpEt2X6JknVdZFwdKJI0yPV38XK+W
hpJGwo739AAC/ecaEgvOcwj/2GcxhEhcw7oeHLKIq1yk57HcCy37mLvRXEZtiuiE
kOvCUZHG17MZVTdVD/EtTvuZ7QYTJdnzQUUM2zFfxKtEYTvrh1CYYITKjGKI8kYA
supFd8ZNStYkWbt4zhNwJNrNplO9UCdaGrc4sZjvrskSxpGhbOUX+oNtbofMgELK
aiOq3p3B3pTg4qCLAVVHGLfRDnciB1lnSMRbNnBgvPAskfKs0fkhDzldZNZwgsWa
Pb5Bk7q8suvIJNle0X8WJY5KbXgBdkAJ3DonEKN8VeaZwJIUpg4fnu8UwAPbrLSZ
XwNVdaGV6iFwO0yWeq2Gt05ZnGqkPP4VSNbJWKsOFUuyIkwF8f178LD3QlSuJt1b
ZOTQpsCzP9msVIFZMXuqCCpE5sOWOmXf2pgWJAyQNd+KxkTdO7Vuvw0VCSr12+X9
KzgPELacYBvm0HHvpZXIelVHi0ZdI3NW5M+uy18Bo6FxfDASjOy4sJDrSh4MUlF9
ZhkLSYDWrSRyEbcOh1FU9mkaRPNrpxYe57ps7po2xedhsOIjr+wW1LfksjuGkSoO
jBcb63D+wjc/UiAWUQkkrYNVa5FAc4g51HbexFbaV1MelBGLWxo0A5o+5aLnddKI
ayFbzF0CWaJVAb0ZwvbITLlUJ8U+q6ND/+yCVWHbqOunVcSdQIFBmXSrWtxXuhwv
LrdM+jVANns+4ihEQeoSDJ7Ypd2MiARoIf9EHMmqiXiFYG9swVhEQ2XgRQe4jQ73
4rCn/kVITQZ/2dEWS9vpHj15HVxkXiGefIvdXujNfhD1hhI1RRX8iZmM5tj1NZcO
Q1Nru9+0ZlpaLeqbLH3/D3TQ/eErS0zf89bRpOcmX4/quE5ysh/sGnYibaKHegFE
pM/5+Rd8U6XqxA/VrTFoENepL1+DISkr3K2ZOgADD0DBiY8OjqY9phgSVJsPbn49
ixsO6zb+U+0XlLkpPhDvix33VyIJXQro2Y9lSf5Ufplh1xDhcR1NFt6d2ja0TOT7
2bhhJg4wpe8QLe4yLxsUEMhnjECV3zoJgd6R76RImnVVwuL93eK2Difi7vd9Ch9R
sPZc986juLGVxZ31Ga2rFO4B/C8ocvjs11nwL/HwGASV9QLC+aLlXgUiGScMwx7O
WtZtPfGvyXyozwRZPiORLEG6qA4JNkCIB+hFp/hlPePrx4HwOEF40tg0NdPTx4we
K3TduP6Hoksy9OUbkGhjRjdUvz97NHWrTentKIKd5mSuIew3S5z5dJo61XmVemTE
T9QflCVJ8MpUMJa/eXrfvTl+7VkdqmIPDNvA6laRB9YD8tpXZ68WiL1kQY1YH40x
QR8xv2HwhING68VNLnWf/3C1tVHSGAP6id3fkcjfUWTGJzJbmlB5RCKPu6NbscPb
IL1ibHhLw0Eo507OWdN84knZNIrfJqfwOkKdedRhb16BKnBT2TCKHQz97rMjEWea
cNCTgYiN5oEzJqtyqpnsYHwPUhEtkz22qwc0QqxzUdDQV2I4cOee70Dx+axG25hE
EglcitNkRJldaTEkOfQ0T1fQEcsFADEgLBUp7hSQUWVc3ZkMJge/kCvoXFi7lIoQ
vzsbixpC7+vLG5uiKxQxjVb29XBYrUsgEHfzGqpcA14OcVzbCiU7HEjukOHI57O5
44XtSuCdJyF7snGDpc3aYx9Emt68UWf5WKDZs8hiBkHoPwv/lt9/yvy7pNdSpKFu
cS4eD7sNf3tolpZPOTTFyEZKy77we5sOoMeVWY9Jyz8N5x6+4uVQFQjG0hGQRpUl
zl40IcS/7TRJOuTTMj1C1i/EXXf8JwhPf5I5gBrTE6LIDXNkUWRk2ePS4ZbRpTt5
Kew1ySGM/5U59BTVa++p9+3PrMPOpUK91rIQb94le1f9SS+LkDqN0m6NbMu+2e1/
EHXiyMAJtXEsFNbN+dqzisA6pGkxwCdLV7/o8PT4KiiavyL3hBJWn9yBfbSc/IRK
MXvhgg2ww61RKoJAOUV3vlT7uFZWJVZLzyvIncVze38bJakzNKjO8vpc76g4QiVz
V702C3NpQIYpwC0znT873oP8XWv6iCZC7ZCQkJEabd0DdoOVbVg7ddHIIdP8ZOB9
gGOxNt0C66UHBEDEv5h4jeMfDyATz2kvA6+ql/IT4nCEY6q2/LJ7B65GuTg9bx2Z
MEeCWZqU/613RpQa7RHnwIH/XnLrYoWk2GBEBfIt93qI7UboXKnDKWNpDCGb7TKN
FixDLJnkaFb94F0SOI3IVzpLvWw/d1eFiswsV0VTn2lLPYv2vgqcC40KU0tu/xFJ
cILcRNTmW4eCZf0nF5PSLTtg6QCTBceGsvF6hjrdlx3uvKf3EZRkkAgXz3ezhFG4
tvW3iYnPT/Vi53tE/UZ8xyE2YrlkL2jXKvJw7UBX8wTYk3GefORboMrktcGWl/rm
gh0y1yJuIiW/sj5wUL6uutk7ugWkkzjU2palS8nZpJL/UqQ9unMnM0CkyYx3odhe
B8cp4Uh8n7tL2iXYAhx20SZNQs9+TXrpItuKwBkT7vbeBNbCJq7jA4tt5zLfrMdc
NQUG+e6lqQ141eL1gE6pTaBAkyxJY2H7ddQBycfD/B7r+hHOZpDjSrxgenL4TN3e
gGRETFB02tOURDdxpXjmdI2GV/odXG0p0kdodssRUqY7yQEpGNTEzZPgDb+mfTpi
uvnVqJ1SQS+a80zFrIY2Git189lislFt//NQILmtrAdsyadigR0yDPHbP1yacShj
epqZD0RqurC2xDR2hvzvRn7RvQnFdTq4EC+hTvKQzFyj12zMBhMcdsFspCT8QZrV
3Z3CcRJBL18+9qXWoMfEe4LmaQUxn1++C6yjXIl8GeabK29F+Y3WUyxjn5RAzPl9
JAuY2zrQhZGAAjSHYMxfMDSAI/s0yg8uU3KhpmMfVStYg3dARs+JIJK1EkxXy7NX
03Dx7zUUro+JT7UjhBtR67q5s4aDlkAcw21hqLswbf0gMY5Jt7QlywTAgvLnG4Z0
K2f71Xj2UaqCFtkAk/CNvJr4kpDX5wsoQJzmdmRp1KUdg8tWaknvjV95+/9vxph4
vXTB+4qBdqBlpyQr2+WJmpOHNBwPFjDAhRIiQ7DBtfBx785DwlqT7K0MmtVIn1Lo
6Vx2oUYlgjmySN0jQPbfurkSsfB/9AwZs4+274xd7irBUcfWAcbma0/Xu2IW/tEI
dYlyML/OyvRXBmeCMnY1KYzEWlpolKaxwyEc4xHhXX7lNsnRCoGEBffdU+UBMNiW
6prRinRosg5WgugwDWaW+IGMwG2dFE5iUeEr5/xEEKqikBKte+jfJeD33RL3sqID
7CRZEvxKg7BYc7mZJB6jbbK/itvpc/KyCu//mShg49C1i4stn/KdAYPxEnvLysYG
f9ztOm1dm04EpVIbm4cuvHuVcPvBSipfdYka77AOT82LI+EOKVYrRqvyhvw1Xuzn
D2jcmOnmjSB36vGc1CtuJgCmTeMd7izWOQNW5QPwkJd3bjXdphLBFPNLkwBA9Mo5
RdWodGiRn/OPjceCyEAxy2KNE0z53BiNupyUmuWBIHsnaL5cg2eRcaafXUpAfCgw
25CyOG4PtdajLF5/TV5whiMbVTUBdV8FuwrvM8GGOUXvGpydUH9Y/VNCVT/FceOZ
49BgVIHxhS/rDN+SuPtj9CZiAsQGvuiCHQtV0V4L8epUsMCMrg0U+5rcPEzqI+oW
9vbIL4rl1WzwqbQirQyPt4RodHfSsIXDHh+wxheLrOjMBpy/vlBGu4RStNWLAdVO
Qvk7LILrAxgwBtFvVc0UYwKXmicgpOlRFRCaFBlOcgcd4Q8Mc6lp5hsfKNRnxx2t
ZUCdnaNiwkysrZ280eFWUkihu9OScc/+TBXWE29S+O8Bdmd7lKmqgGVGiTY6/vKj
NkB7KvjhAQFMZ8mR9THtTu2yqrWJ3bB+k6HK+03h9EhUJiSJMcTuZPiXPwOs6FfF
kH/9ioByl5/PW/hRwY6ZMMklqNSVV3MJNkBBNvc5hGfmOql1aMA/8haW59gnUTm8
i1PTpDOoh8y/PcPDU+AtZGww5HHq443PjWwXr4vQzFickS2d5QiqJj234Uy9hcaA
Q1jCJEUpVC1UzFFX0bJElVQ4UoZRl59RZUyXj6mWYzXqozPqaCftMNuq4GWkxZ+I
c8aqBBMtSI9L/L5c/4abobKF+yKLsQgS9dOVmXIhx4OQ2Jx3oo6uoAwDdKS2a7ys
dYvUivQubyo8A5a7z6ja9aGMzLfaeQUttwGGACw/LJczZ+v6nzq9MB4Ej0BCenRL
FPVX5ppoJVuxIgg7DS3lsP2LOOVZJo/r6oVQ11AiX+fNI0Ym7T6ZV+XhGCIHH8a4
fTbUxftc9x9nzZEoczEpY3QPM28c2bk2jHu/A2xkIOxQef0G0/5ecjfg1CvM9WhQ
sgm8GcLa3o4qXUj3RZt2NquaUJsmk9jdLFr3dTDKTVl9o86Ekh5MNmILsmF+XeV3
WBel2DUhRTqmVnfPoUZ/l47l0rXKX0b5nkv2NFCmq1oqPZTC07TPIkq03QrYcLqw
daQSWyJ5aYZXchSSjKIYdtm7k6a8AizH9T96DXSz5uLj3yhlkKuSCzydeW6zE/YT
BW10c1FkZ7QybAR2zTUk0LnuSf2BS7KrD1Lv65xYuwd3IgmxJjN7ltqR1/KGTySz
1tJMSdgrIYRc7tfNbzwaX5XfqVY2zzLxCPBuG2SoM8Rzuiu5QdqpXZ+0RaMT/H2T
pvT94N0GdWJKBuIYNhskO5w7KCqmuop2gDGCbG6hSm3uan32b27w7zZSerd73j13
6V1o4YpSRpl3VVqTLUE60KzBHC9gwyEkHowziHCGGrK4Sx4pUZDTK8rHrisWZTTa
+GfoALEL1C3Vi+SyPKeNhgKDSO3ih0J18FDcKN+RcGOazZdgm2NNa/e2ewnADLne
BNKM/Jy5mD1a8+h2WJCOJ07+eRZwC2pgvSK1mSc46wUaCRxtchwJVRazmwvXuCPl
11qZXRnULZZijztZrmLO6wsW6XYq6XFBaIhY6/B3h3eZ2xTWGQiH4/CG9WNLMTgA
vVfOcQvrKe7UsTFNTC+ODMfwWy+MEM56ntsY6rMvk0pQG1GYGmlDgjshn84KBmvt
+aEIZqBY4wN57Ikr9KPbetoy0rZnv7tBRwQVwDgd1CzY8LldJGDjT8O0nWJ27ATV
VzsdQ2xKwlJzGCI+asdu7LzEG41X5kRsfAvoDRNOL72oiUo132ygxwEzCnwMABG0
V019qkhv7f/w3EOuMIcBVEvpgSvje6L9uGuBGcwY4QDcAk6ic6P4MRyYuj7j/29u
Bd29yrNDaHVmQfVuWfEHUGV6AW9k79GpF2TWzGnGkBcO7wfS/FuQw2qIf8k1QHUE
L0X5l6RAn85Ds+43G1wYaZKcKrQD/2kcR/mbih20VEFZuuN5ojqKx/zN32tTRz1d
BxpHye23Mkx50alAbfJ+qLoD2rJKOSUifH6Abf4KsstRIM+95Z1qlvTc68LEv+sq
rmihLpa27I4VIng5zTmpL0gDGGzF5MZxrcZ/Sv41sEES0CIusTsDXDsSVtAuMzLD
BO0pgOPBncGXNLyDeEj75jbsEbf5hY3k39d6PgN2hWV9/MUJCoiMZkmSe6GaEE9G
Nu7h+cykAuq9gtJa1oLJMrRZjNyDf1ppaVzOdHX3V+ilJejOjvyELtTcFLJmTcW0
WhVhx7aZ1N2haQzd+S1Wlhw1ctBG87+fMfBJTvUbe7Y2JItBCqfeTpS6jMNF4Bh5
csA9h8cRl6JQS2HcbebEpgSUJIZJy7hB57apeubpfLwQAuVzfhQnPO/K9a4GFS3m
lvGH3MkN13eNHBiXq0H9XdsRG9lqCZ/MK4BgBOrqTKykSmTqhj/Ns2Wnf8q4Lp6D
d+k3YE5FAUcVymUGKiv1TLiWa1BzHdF3oiureo+Hs4pepgFWElzsV0KEoEB403FY
YMwk41UCWoeY+Elow4+Z3RWqbEE+V5zIPcnqySqllXdA0lGyLJCxsLO31nMusMfL
mdvY9+AH1d96La2/kp/aYiKTCQVt1CLvOP/svqW+4Jw4VontB/Vnba86o4KozY5u
qLXyg96aF8oV4rA/PWXxhyS+e16lIYEekCPIVhrriJZDYtOW1t4gx3zX1mB/8il9
O6nA/AGVlCvCWSX/AMQKmS9P27sCCghyGIRwz1S77OMEhXyUxtyVafmItZR1trZe
kNhomESf2eXA266MH89Vw53QVeENUYLfqJ9198aRBqnFcHbcKBiNZApJ6O5GMAuF
/ELWeNMt2zxxFcwyyiuMsEA2+e1z+RRimJkqvfYm+zvpVsAZOSGPow7D1GIDPGpq
5ToP667aqkmmzqXztErtjmSFNodAhBamcJMLd0Cur78HxyaeSrwoeSoGau2ewJMe
wMsBrvD/GgQa2SBIs3a4W2bt28WKZ8w+mbUlZoJqn7KS/c/JoD9XlFpsSeizAF6H
sGhirSNyHMDY6kCINHCbLxwoqvsKdkzfkVoB7uSlgtwCsZi4HndP8jYwpCIrtpU7
2bQzAwpehMdXNrg4uIi6uGAm8SdoItUcAF1mquH/b9sonCEPTJvsvoy6sLNSaqmf
pRc2LGIcg42hxkDtIz3Bjc3MFCB/4jQYr0masZjr/S8oTQkWs+XNsLTo3XdCF7+C
9oeVrnqq1yE7w4lUBmfY6tvzIHQ/hzJgYBpL1qtFoMccZpBpo1PtsxK/3UvosUE/
VcRVmIJLzGrDr1QieoYloelQHnXPqMNMELPxPmt1mJnfcAhT72gXaHCFqknlWxGo
mpHl90mdMkJAfVinS16K0VQcnp/f9AXGTxVSXSKDuJQOWpJGH0G1byaWX/4RHEvF
luIvPflZZF/Hjb8eK7D8xhriWLa267Vo4HYBN0VzdZ1rH65Rwd88WRQNdH1ctGTA
tMO4Re5H6g1xBg7U8gVmppdBQd6mQNdNrfJTWtzLUfInv6JPDakTBsACx6Z/Krey
bzhcgMRs6pDSaqqSKrB7JoWMjvXmUawkqqclRwILcb7UCdX4wNdMvHGTR3wTfGz6
qBCKu6cvQClI7xS+ivBOTCwwRRRfuvSXnWAtBWyDaqHRMs3HQX4M8MHn3UngBCzS
bLyHo5CIoacw0iuSiu0ia9NKEferbaZU4Ta0Fs53JUXnDA6QvQFK3QRfLTUFhGjf
QlSCugC9/JLnKvS9EpeLjuySiLCASYNeMAOs9KOI1qkNWGqJgSoqAgvCkDXINmuU
oaR1geoc2utnK+FDB8sefBlODPIxbquUCiWBiOKKMqBTZNJCKcIzS73UEfmBYhUv
6pN4YnbuKJcYrmM70vMYJpPtdFo8qn+sQJwgUUPvqZxMaVbtGHPWRXf2JpWLL9Ur
oYgwzU1L96DchFJ0Yp0UYpEG33pX0w/x+n441eHuc/rUIn1CYIJFYmSpjrKtuums
gUs5Y5bak1EcHYqlhXzCeJl3cTljOjJjeZf3aFiHEiN0zGANta0nTfx7axhJ9yjk
vD+/s4gwCsCiLaHoLNZsqlRo/8XXk5Md3S2LWxpXRzwwdveZCLI+ijpg/3X9rLlj
++RFCP3Bl4Itkxy4HTnnTIoFxm2JsOA8McVdSJp0J7Y04brPFCtiT7UP9GB+pmQi
zu7Vth/pxDxZHPXlrPB1Wn9L5Bida4BVjTxhQ4AiyyZGSbCsM/93UJlb4B+ZaaeY
mL65ufwcaAGHTf3szTcsSJdg4VlP0jKDQdRbO31HrOalYjMNGxCy0owEg/UtZdhW
5y+HNWL4g5d0nntxN/83RII+sBDuQsOgAbxNH6cSKWyVNg5R/eg037oQoUma3qaK
XHu3WxaX8OkQiQMIv8kqT/rZ/b8YMK2d3C3ORcl8NBHAICeqHAhpoGKJiGwmYU99
UqVoJQEaUFyf0cBP4jfybXxuibufHqDh9MVjZsOM2wcGy3By2gZmzCmZR3c/QgXv
UwCifF86bClJR+yIlD8ftgJyelHs9NloZCnEyzvRxdMGk/wuHHMl5igsDmIzSLcS
XMkUJwTWWCQJsT9VGwy5m6zmuCg7pDz39/wK6CBGObLIs5braH+muku4mV9AVkTa
MJ9vsln+fzyLc+i3f5Xk7/lqlss6UjgmYfU/DynjAS2MVfcZ8cUPaor3iRTwfemi
iYKL8x8vYvrdRJ0kILv1UoLRWIPlZNYDyX1Cd0uEITMXx+Hc1/aUMuzUaUN3pRfJ
/XvRk7fxRNZIsps5wxrRm/ZxLig1N87BYfjiMAtWLqnrOEp1kIRJD4GzRimmjle3
ZAvvLtYcPXXy9Pm98y+OEvRhBvJr02lcFwyxC7ZzUdmOtZGnQihxmVxQtZiBkoru
Qw/x1ZECx2npzW/VE3gQszMR7A/8vExEz1XBv4VpUIGcdwyc9ywbTFNFD1RYAFFW
0x1KddbsomnAu80R2oMW0A9M1ViKcIwnj8xpALfe2tlEXJLXSytxJUcKeSmgkNiH
nKMqC56diX6UQ6vLPs2Jc5izGNVuOESYh8yaKOmIHTtWn6NBfhDSJfv7zwz8KQOb
9TB6AZ9Uo+i9WgJcR0LwILL1zGuQhp7U2sJAr1LsU28lr9ZEuBl+MrsGmKc72aSO
FsCrvKdpWtrfVnTNVKcGkwZXsrjT+V9+YzDembOaCFNNNn4JPQo85PheKrKlkMuh
K5iIWdf3CWYDTflJHkShgMrdHhlpnjngjzNO2zJOoxz+Aul/yssNAOr7EQ5RTsRz
I0rphb9024Hov9GhGD33PFzdBjDaJ91kbdOvhrFDLTHMssDix6jk597C1T5fcRJP
y8S7Zk8C35VgiLVQnbb0VAQPtKqe69FAJfoIedwBSJoHMhTUHpDmpH/jOdK6fXAx
KMNgArmmFwTOkf5m47+NjH1+YyiXXEkS37Z7Fe0akxfwM+BNAYBiEluFe07vVKAh
cBe6xexvlAHfknuItoGvAHCXuuTq5ZUuoR5H9DGsjxcuyLhw3Y5ZGDoAtanCtLZY
I+oAzs7hEVxMSYyPm3mfBc70NeqyARG7jdyNp3/amwnoXx5qA01UDlmRWG94/p6F
gWJNRnveDuvdn5Mq5gDbUcsd96buU8XSJgDeQleAa7O0iDDY7jb0vpb3ophbhLUz
eleU6jKRTW0C0py906ZziRNVTrJpmXftS6kcmhF50WgRpCyH5o1XkoSHxNvUPwiW
l9kdBTVqfBv3yn3va9CjnpXaPrT/AAo7w/QIp8g+sOzCV6ye7T85MDDTMi8fmpTD
bavQUIyUIgokTocoSqESWaXJ1mp582egUQ5uti9MYDxXSdvldqU/QNR0/BsLNN0V
C/QKtiLCiyUmrNqCPxUdoYzW3NG2gxk9jZCxuA4UV8apRVbiKy4etrBPpmUiLspX
0sV1XVWRww/zDjlSbxmsowg5vqQI/foqhURSDXBBXgIfIT4hVyk1Bu7VOu4+LzP/
YZ5/0t7MAAJeUbhgpBImV0u25uvzNLCXOPxjJ7le3BBrqaCvT7Wa6mQGskmhE7ON
LLjgo4s7aiZSbPGjl4JZ9HcrbgYUSAelkm0CUfQAYcsF575ejK0I2rRcUTb7Juey
2Holl+voEBGOGoF3dMrIstlbWbwoY0zgXt0NU3UcPs3qpjG4VIbFofdGGskmd2I7
9jK6Ru8bn6V481mXBwTDJewftN0Zghb30r6/12wKZRih+sDpB5g56Ihodi0bgjSy
zQyE7oGXLoM5ynsjnoakn99I3oIenKWEtUdiUon/qb2Cy1npXH93HIqSugvqCpuG
Ze7o05PXkmwzPpAtuWVxZUrOeoRBJyphTeFFvXWH6Lu4rfuf4Jg1QC/zDiX/KTpV
E+bRniIOyFgyWf90V9AnOe9XDMcd7qpVwVrfzksnBpdXv3nUnQL2neXu8o3dm893
xi465KBUyxZibt/oPE4X4BdIYSX/s9zyp5sEwU76wPk=
`protect END_PROTECTED
