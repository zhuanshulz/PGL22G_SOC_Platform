`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NYlkKGLRSDa0jaJxzbpmChdCNHYpw1e32Sp//R3ndyTiDfLgD8y+VOwAx/ehZwdv
AWiy5nYFBP9mgl2PCnZ3v8o7FIBReIphHnAWwLDH+l2a0TFfuAtZVmBktYYRlGNr
/ZEfhnz+uxcrtu6dzCLrpAxllcNa+fiZlQfmI6VrdUPs5UQsjH8pz96DBXJcIS6B
yM84LKB2aYdTjdLfhC0ZGlbsNvIUmoWOph4/SvlR1J3zUF4xET0GFZDzq+SHG7LG
TzekW4Bk2paSmWew234o9kcDFI0SJ/u/DNCu4DZy/ecsDBgnXFj7xuf71bTvViks
7qHQ4qFoYHNhT1XLASLFLjQ8D31KoZqFZtQofEall0KGaLsghrXj4J8AygbiY3JI
CbC+7xi40SBf4k0lcNb6dBcL0Z8M+3nfnIQxSpuSbAxAYRGNnUrEXUUns0vD0Zoa
6DzYGky3N4AKQfKfy2R8wws9hUkixOi/H4VQ3/Pdcj7ZjqQ5zEJpWpqm3HJLHBCC
x58WmWh85rMv78l8FXCY1pF6RtwA/IBwKBMTwVLEtx3rf+RV1GLjQcO3uiw55b8q
/Xq/K97o6/qsp3DrvAzIJA8z5STovTz/NvxIkkCdWTILN2YluToMxVT/f2NlNqic
0B86lf4Z6Y52XParsgjHsoB9e4mzb9R6RNjyGZF4f4sugHhpEHJHtO5UHDJF4Y/7
mXwbWe4wCA2w4qTOdGz20jGL9figoz7c47ANJuu/acJvdRXQM/Mg63yXNz3dAx4J
7FldRhZzbiBL15o6Ksj6FcKhB7tHYHaxnL2KQBn76442yViICYDWAyJBlfJEnCf/
EzahcnyCPM7UKxbrBu1ScuLm8Q6FnLMkQSOMSUR/fst2oLsUr3DpBWhh5ug2Wu78
i5pYK0wfHETQD70cdVpIon4y3hrFxz1Tvthe1lWrYS47u2N0/vQYcbbhTT8yQPNl
a6Bfgzlcgn+EUn6ve1SpiG85iZImlih+aN1rJyJBEvmC0g0onjV16LIx4q6wPT6o
n69SLvC+Eq3Q0IBPG+tKEwpDHIaiXSglKB/vduVlRjr3hFIbF349Tr2sSftGXKxh
ezccKDY1Mn4ga7pzSPDsfWUZqNUaw6WHKM29LzAiV+oqDcrC/Uxv7rDJQ4MCWxlw
uzRQkhQDaIj1Fwz2aM28bq7nOVLsNHkiWy/mA0pDA73/4Aq7Eb6r1JBNdO4IQhk8
VT8rL1PKPq+4VoAjR//cNIDuB5ukGdUgzY1yT6KUAbdge7MSNvDcZAjNU1bF7INj
OQ9AslDWaaPvRr4eO+waVvvM4L5HU+UFHf/uOg5EOlSW7/JLHUOxBoWd9+DUO9R7
lsEdaDGW0/BnWfIDdazZE+7DIM3u4I8jsnzG2QKjjPDJvxn9xYdlcNAQ152H+FDv
/epaB3IOoHI8mlPG3hUQ040mKqfaHKNknyXV+sLPWC7Aj8QaTlozieYEhR7T1j3T
3sRH0ry/cLO+/HpDL5ACGFIyHkss5AjPv4qHbyZX/A7fBGS0ZSHF5rlZWyxGh/We
mQ1wCCsM8nK4qGoHHKwkOKte/iBXL9nTD332l4gQ/UTihfbXVvt/nKpDT6WAUAz1
Qoq7ic4ea68MlC2yscqGbBz1cGuL2uL4L71jAeXEddwdZ2dRXDmvsXHiReBS0p1w
e6KrJWgldjhtvYDOsgg0F1MIV2vbdkPwQShXkSVVUzf9GMAiP8zuTgbqS/9jtWjb
/fFrGTL6TLTkLL71dbIOgzX5rcIYoqnyPKipgYNJdLNmlHTZ5iuB4MCDRx7J8LrE
k9+7a5yA2mjp1NRd/i34gMaJT4EHfTxngEDMiccY/MN6W0tFkKoMC1qUnNrWFTza
73SgmIgerjlfwyxZTHQBHD8RG5VH6vAtbaFmetPxhSPPIOzIYUYD4nPaO72kMR55
3jSedKQY7++hftAbKTbRlea2zHJGGiw7vayk13lt5DV1UOkX3nqv7LThmvUYX8l/
7MTu++dbKzSTbFSmKxiTXjajD3ctZ/ax9100pHlKHBX0eA3NNI8ggkX7GKWbGdSG
H5ztjMyuF6oDF4p/HCQIii2A10lxT2qnQ8MWtjvtH7DDZ2vV9d9ji6DUrt0+fzI+
1QinTnD+G+LD+lM7KWLsU8OiX/QNIfHTKJxapxx4M1l+HX1e5o7XIHE3WY4Lu7Sk
JW+lBsPJHcoVbbe+ov9jZA5bic08uK3/5l1Ft41iAHeZna7MTupuZl2JNR5rgo+a
KCVlsUiZtuvdyK5co46yaBDJPfl4LGdEt8MVbI2NQj2/rH5smo/XUY4N5GY0Mb0b
j9wHYhAZ4siW6YklNAxfGMnExoo1LfneZy6TCfZu/MHj1f0Q4Wl1YqRNoYy7qycx
X6DLzNXnVtgXigBiSVGg1kGrTWoqprwJUmqijSAv0E3mdut1ccQbSZ2/m047TafC
3yhS80VAgyfsjU4D796lUMn2n6PwliRiWhHUnlgSIVGMTMBYxKpap/e4tV9LaClH
uZ1OcD3MDq3KLgNJfXT4MqfVtZlwvElr+aQJatyasArnrQablwg4gn/9QUYqhzgZ
WR0Lxp4PjAFkhX70g6CCFKwQFWpaTps9i/e16U6i6g+iQUmI5CLcAcUTSgXM3jdq
flahGWcfgOXSvsGQJaPtj5RBXr7Xq8LFGlvv3VQ/e6FQrjKVRRu6AGMkomPVXtLh
VHPNDO/fZljrvRxbAoKqi5Fa9s/XsR2uVNlmDK5WEPuCmkLvQyFVQ3s3GBVl0C+C
b6lJ7r3O1h6xLg96QpC4K/CWTrp69HU4lI+fbdLCsSaaQI6U78aaWiYV0mdHYOMO
GnlMNBmbvgUQm+Mqg4rN/3SuHiLpEB7B1BA8bS01XLLTOKjzowYer0CGh0TMbYQ4
prSvlE7Vj82LXGztt1d+WxGsH64QQ3/ZzFW+Gkj5ZHPitWyIzLCb30eL/zwoLlBb
oRW6yzTyTyw3LWKN3AkKVcmDdKxa9r5LAoWmSUaB3u/o3CKQgQe+0obTnjqru/T8
cFJnlw+Jy9nBDUyB1cRzT54GEdM7mQLx9mrVoR2BhlYYvFIWj5o9ZKT/5oTYbKJl
gtABN/IFLDbbwQ7STH4shgetzhu4nYdiv+TtMjkC95r5Pp41jZURlOKi4ZqHnyTS
0TNR/CLe7K/3JyCqWs5x9aL0eWH/MQz0LLZymzJcWHLMmGWwhulJRcQJ6chdTqMq
FgOgGaBooLAuRVjqO9593yrxniW7epu/I66gLMRnSiJ+4AX4abfWFq7zHtSqh5xJ
w2ej7HMmbYzrrcHif/bH/9UUYLypsEfk9lz7cpAVlRbMVuwDwfj2JkSUN/Wkar7C
`protect END_PROTECTED
