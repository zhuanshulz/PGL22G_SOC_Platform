`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BpTy1BUniDisicKrgVmTwrtL7JMDGkRiKKgwF4v1l2RrasuZualM1kb5z8EZXMTN
k/UwhJe+SXvghwGFrdG9FJ5m8qMb2jA8L5NrD0A3i+3SeYy/X0XN3NDVs9U0RL1Y
nvvVoxkPI63tWm96MK5XdYr1PlKBDNAij6swXZnFSRCFCGnC5nWeC/VL5tx98rwC
jnLiyHh8aNzoskeYb+rK3/suI26JdamEzJqDqPTeEyO1sFxx0J0dYLCxSb/l4Ivn
nKoLz54aW0DVtiQPPstAESG1OuzUKcPuPXGAqUoAO8AV185ncIJxfObJmJncdiOr
Tj2HACHnH0Nn4152lL1B8a5MHlmST/U0lT7ot/31hobAqXuuxUorndOmLRgNHWEw
DJih0iQ+9bUAXe0TP641oeWk/XGf3ECLtW+4yxIvp351QayUZM0fQeGueWb68I91
8hwNeVnG0Z2UaTk8podPkCl6HPKZmAh0p2FAABcdx615O0GmAz2sm7mO/wW4PhdT
8eWMldtmrwyqXSs6dS8pNZPyoO5+ffdxc+9oV/eO8MSbN6fQnRfbxIbuqqfny/7K
s2LEMrEzOB32Dq/zeWzP4jkCMhkJ7erO1sIhLCM4kaJCPem1YxT7/4Y2b/3rbETb
CSKFDCszP8/UokqozrigQvWzjWS4m3OQrWltXy6ycWqEUIH5cLuRGQw6v9h4RNwM
cLOMWxAoQ7/H6gfbqcQ9NhPw4fV0X7PLeN2jkUGB5jKWxTHVfEYsiaZqNshH60CZ
vRD/qWeNuUdrB+vbKNbXLjiOvJNbKehD+lyTm/8suhvh8a0hZkyvx90vNoG+3VU5
9T900yjdW8SNftaNuqxe0DqL/HQtWbopYpXwCVloaK4dbUnMBALFMJd/I5NGZRNr
xRacOckNroEx8K3CrJx+dXQkrwLcwEH0syQmTP98KeMKLDxPYh+AQv6IMLMvBlG7
wbf6djUm6uEbhicMTuNetSxEUxvmgUxqVw92HcrIQv/xnq6ZctMLx4teOqzFYOqn
29zdSTS+qTZFJ32V/4ntZpuSl5TyLOdpvKxRUSdLM/AT00LHDzMoC9n1unziMaOq
MHdFdWKkfYl9OghdOCejS40CG2VIX6f6NE4ijH8EYpbpDirKMtBd8R03cB4l2TDQ
h5aGhqhI2A3g4r6d9FDAnlDZSFkjRRPx5Agx6Kcy6fWG0Un954x0WZKnctBukWEK
ftY2JC8fNoF4l4AcM3u2DbGposDjnafi4GeDEG88cmLrpyjxH+do0Nbv0TzuFXL9
yY4NrpGu+EmW+J5VgoCqKQYMuCBa0rb0pDgbUN1GxzAQsWcdzrs0i341kmItRAtm
knV877rmtpOl2p9q9Uua1KRra9Hh+ZesoL/oAlc4EuCGsTXbchqfjRsiaZ9M7Rgg
/irU0PfoFf6tvmQuOcQ7kiR179ge/H9JAwYGp3y9o7ttWRV2i/kUbxuxmtGggUU3
StYJvJI+XqraL584RQkM7fhbDwsznfVwDEr56JTJ86kweqfBHLdRrOGYDmABKszo
`protect END_PROTECTED
