`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gqbV3nXmScKCNk8kOOMt0Vld3LRFAOoJPWQ4XubjJG73w/dJjKwcaGNlPt3Bs61H
8VSYXIr2hDPXl7rSWmvhAO/cQQZH3uDcVTrb8kZevYq9ftbMt52+8fuU5bkTrMR8
jASyvE1Ddvf9ssScyf4+wW680t7ebJm2fKYo4+6luxEawO2W4qg39Jgi8HcAwsFB
t7zRu3aRDkto1Nx8Uz4LzuqiNwgFOUp/3QiNw8eZBZNPSg7P8abvuMNG9dTOAJuN
4QYWEYsK7j+VCdoUo4gvoXsSBTAOgQMxR4OkjAOZNqoERYb/4cwd1Qyl2uvbl1Zn
8B1QwcMS5sJL2TDPS8A7LBGTT41iVWLIawSxnntbD71td18G4RSzoktiX0Wz64gD
YHWFZBtGAiyJusv9eEgNU9CrkE7dK+jBeaZgMYTUbqMdOLq5lClxqudRWJlTkO64
dchywoR1cu0pkRgZ1NGvMJaWDsfoYs48VUIA6fQa0t68V1RO5kwMpSOp+ab0Hmb6
A0CiJ2EBwmKJ77pnIbbbj6fKVLzZDAJ8DN84HRQLi/5M3e7bD1r6gQOSnEULZpJY
ThTSxFR7a2+PhfZYiERAHoEc8Dt5V5lQylFHiAok/pBiKWORrYfd0WOX3/wNIfjP
fXWJD4OgRx6TA/aQ8pk3l0yWbq/KjXPNvLIRyjwjiz/dBTqe9tEJOqM/DMqrHDp+
E2SnUtI39VRAVvtJg9Ai9lGsUKHbyIsyHKCCk/PszdmOsKLHh1IHt9NI2UaqZ517
IhZOZ1qITYGa8ceGVyU29TBPLAoVtmKMJtKpQcTbfSeE9Fmo6dkcXTwEXf1C/8lA
`protect END_PROTECTED
