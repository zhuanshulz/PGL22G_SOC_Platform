`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VApDRIVzPc6rHd4IBlQtrqofrHWi4QUoQHA05nhPD/Eq8DfocsuXAKJzpcbabZTz
X0II990PhZmJzrej4eVNYZIf+Y7q0SR791hb4DgNA+rHFRmyj5zICbWSeBcb6mU1
MH8COPODvnoSfupIM0Y+c7POZtjr9ytvNgsB++bkL0R3RgEAp1Q86Bm+CDwrdvik
qAwaxE1aAm3/iFSdv+biX/sff4oddfOUSdU1icReQvRfP9jCAL3XOCXWZwJ6lx2M
RHEn5yoXcWghRQTsBrwEfYbCI7E3mxkpPE061pTv3uIZgwRLsmbe7e6gJWOE0En4
aWealyxNjgKY4RpN1MSwBKmGZm9AGI/nzRxvSzCPBzeRCBfgSm3NOSXmLNL3xPF+
t54Ld0hPulxdysQ1GGM2y+YqeoDYz0Zyb0qNN2LjH19D14HzrxxjmbCIVGttpb9J
bvAKc+/WdVsW9UkgIKIiv7qyyF1jQcygUeY4+6PXASfWN+6Bu3LNmw04d9RUpnD2
GQmBVcCZapyFbM6R1aIqKkJUbv/FXdtGJcaQAtoN6UEZPs0Ky50+2r37TPWN6bLN
zUCH3W5lgdY3uZzl4DS/dnZlBz2Gt+cl0Qj25tVxNc27+bl7zeUzlVXc9q/216J7
oz9q5ZA7/S+dGX0/HjoVBJHadPrxeUe98zidYNcu8wOg10/fGDOslzUx9AJATVGe
souEwQFDGbUlJag3ljZ9gvuAJ58CVsrhb0BkgesvwAZWlyeXQ1Wkr8qYItFVlOkx
nUBHIH0/w1Fm7+fq36A0/cZcROSVCkUJWteJopsA+S1ECzI8rpmaCcJipNXP5UiZ
9ndNQjV49wd+d9DSlImUOEcrJybrd2QHSF2p6gz8iw/mgSzGJcgsk+sPjVzUQKL6
1hpmkapNeKzkPhFWs98XCGjmysX7fYTCBxw6XVQy7XfQr1qBHtwfjyOKiU7z2mlP
8etaxk5ygtxCg9SR8Sx6ONHM1dd8ew8AUPm6+UKC2m5a5uSJL17kgPhY9KFq78pe
A59/k722CSQ/atDfVH4s+wv2Ef8NuGTnWwHKOdaogIDigBDg/Tk79VuxCgHd2+5U
l2LwFibmbj5SVe7bRMtZXiPVgCFC5hfPt+GGciQtSDrxD86cdW0WVNGl0i1BeWNQ
+MgpS1C/AQ6n9FDxb4I6RR4025VFn4ffO61ZDVLtKYUTtvdtEj+WZyTrfPGw/ZLp
18hI/OTAH0+mWzDvpAKI2DzCfiwu2fd52S3XbnItPPgygMVIfx5vKganD8mBOvgF
s9kE+AyBN2GtZsRun3xTWfOUKtcYx9uKzzmO98icOapXiTsRZsJ4SuGGaseOwxyL
Bn2VgpJ8oJr3on8SAJ3G0/YQd+7fnXCTFTDT71DD7wLfoSxHMbATX3klVMkBpXY3
Baptqqf31HzRRa19onK/tYZyoEE3E39rKzRgtOZznEPF6y64HKLBdDrzCD/FKLf6
c6i+kGa676A+QdFCh74izZ73G97209YHMvT3ge6k+Xv1SgSure6gqYrvW1DG8oX6
XRrUtflkjNtLEPxLPVk39TJ++2dCuHkBRrGCPUNoUgkw9OswX13I5P9migsFrKu3
efnf5H1pumYJASKdp99p4kJL6nMuheVG6RdWd5ijbDunWzA2yPOta74dBu17VD3i
EC8depE92OAK9jucD+viJJ65dP3zdGKESY4AepFqTg1eNTylJxGDeYnR51RUdRiB
GYTCn9iyiXuUUErEMZYYGMVzJUBfjttHZbvMmGI5pdQ4wCWmjJwgc1MV1Js6x3P5
Ka6RY4ytOf2g/h30XNYOktvxpKd/pxGRbuRC2xVjJA75IOmLjbT//kmGo8TmFN7M
CYU0XBTdbXHxJUAua6Nn6T0ehNWK3q3A6b6CExaAT7evXlQumAWBKy+YXk/d1v/l
S6dgqB9gxO4ePdmFdt/BYzmHVXb/5eMFqHQDs0e2c9G6PI9nTDaF2LaZweDShdUP
IoZonunxDVcq52lTp/N0J/5AAkr4PrdPI5FlGRQ+d0RvUIowgqWZhEttU0nEhEIu
t6UnZi1T7vVGua82Cv5E3YYk9iH+/vq0YBWEKD13/6BHEsTxuNiYFtQe1bi374bP
6/Un/P8lz/t1Fpc1qy1FaDPQEk3Qj6kJnba0uYGVG0St24L0/TFwCy6lFIfgBfyp
aWUJgum9xNMlgEz/oA6fUivigif76bviPeJyzcfGA/yMWT93OyZA+anen1O2qbCt
hSafDwE/wv+qugBCWeSGblYinXwrBUTT4/JDKD/VAWuPZsXjgdTay5eRnLcXgpPA
7depzba/2p6hD9E1HyMCOrozpqbAASr8ZV2L7oIznyH3qiXDyY8slv6Yz25HswFK
QptN5eYH/bGpnTaDMu+LAe688e/H9MVE2Js4xj/gBUvIhNRjuw8XSUouBHfH/cf2
cyh3l5l+fSXV/QjmEqEew7wrAUKfPte2l2sGPIr9eHM5JKHTeL0/CVRiI6BMl3qu
x4okdcpp6Qcw8fsA5rSRzUQ2+YgW2nOSq6VRopNBbEJFXE36+5ArGPRDqVgvC0Ys
DCa2pO7SYtxt7wgzT4fapEiQjE7Y4FyD9vGYkT/sw7/7xIDD7uh9i7yB940Y5jjU
Kyr5xp3o0Z+tsMf8hWq1gJUN3nWJEYiOR3HB3nfWomPedVRAFLDEUwDbtojBPmmt
BateSWMXUzDQzYbVR7N7HyBvR5Dpw3GOtu7H6TIu5MGaEukhIQMoSTz+VlpZLtdO
hoIY6qYXq1pjIK+ELCDp0w==
`protect END_PROTECTED
