`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S4VZ9pi9X69b4QBq/MeLEUnxxR/2l9X3w390ceLGHAw3gMEJSpAF61MNXcV4Qk7D
hlpB9Ecqe33P2JC7l3pRrX2YZ3tBU76PCwvyBUNd3OTFT74CKP3sg++kyg22gjf8
tkYCpup+zaz9O0YMHVkyccclWJpB5Jl8kMvDipn8FvowFQs2JcCwTtZ3Kxr/3hsO
CI64ulSMSAPBYsJeeaiXTIUYdxpL0Fm/VYe8rUVTWavaXonPnDcpNvd5EvjNXeK8
YUSaRlNUGG7dX+NPKRvmEBQN1Q3sVOCVNbJp0ljLXzgnCle2RYO1we9dDQyt/D5q
yqbokYDy3pjtkY6+pk9FTyMiCfQWmVLdAbH7ZqhNO9k2kqqQKnpXX/UZi5FbJ4h9
4+ScSZTBlkfHPeAz+HovvEpLN8mCZ0SbFm0fZ1oVTrCsID/OuvDOr9CCr4jcffV2
JDOGeBV1S7aM4mWLcmfq7FG7/cIHo9h49U85khpCyS58puollfyWOTiOgG7drpaP
s681Ap0un0vaU+cXEo8oCKTe9IhAyT+a5id0qGC84bekqUpuNqeuwqmiTgBGfIFt
ulerwB4wxijvjwnRxGWPdg==
`protect END_PROTECTED
