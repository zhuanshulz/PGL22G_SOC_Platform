`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jqLj85YH5RX/8M8e7iRnYrE53J46LpdERVzlDTOZRXreXCyJI4EgN8neAp73zviQ
7aCA0klmB1XK+5yh1rdHK8UMVJqVlEZwfHVRBGZpPrNFBbwzlh5EhGmIPmXcyDj9
vBrqiSuv7lsR9X/vx/13fshKJ3Qye1BuqVi6bmIHAt+nHfDg0bMGBJ3ipQFmaakA
vzHbWcuou05d+NoVPK9wTacHAt3eJuGY3r3JO42w7Rb6JpMa1MD7jDF9QJ6HDxwi
7eJu7tpI9KVS3zaAu1iHc+djTKsaI0TGC0hJ7XeAfJYQ/Etg50OBKi+Vdpd7yNq1
PxpdlvEhEOfx4X6KRRfFVr/eHOX9I3I1Ra4VjMBUfV+YGb++FyBLnQ8nmQF8f8kt
EHHkt0IcYSb0fHqlE17/BR7E3HBlbNFGGvHqPUl7GRoPmnZgmO1vsXzsoMFNOutd
TpKz1NfnyiCO4C2tU/TZPFHiqc7JyW4aw4k+IEn5vYVVyqf8xpzsgpea+mZEkoPs
SSoUuyP6u3yhxVcUX633wGjgMeobcuODH1steihAfmCyT0q9xHSEsSF1Bef/Zmsv
7ojklgibCy5wz0mV5BvZseCVLcS8XWRrrWZbOn8yMPM6SN7FcCpQ+5EJY691VVP0
JzT6JJEaMQWJTJie60C+oBoZc6on/1ehS99cgLOhsUQiTaAtVaHp72dpZf1VZJ+W
zrtoXmIO6ChSlAO800tstYpy9gTYYIN5oRoItkPX4ryr0ZbUjiQM6ecgwC1lrFzS
CZ4T2xvbhXb/Zy3jxiRsiIRzbUzRvyvwTru9b57zsN2SkiMH2DGQQctETBqF0rR6
oly1SI0m6zuO1fBZmOaNFDz/zKkGIK39AeD/NipT1iHf5/t3kmLkHdcrQ1J839Qd
0739lE7h6kWCLVEm/+GLekM3fmBl4ripEOEjFs27+f1uSj9qDanUHJt5VYZEl+R/
xRzlR4wSrrojNmFs8B/TMb+VzAvjuJ/36fd9AVKr6p+uVXhNdZ4GCTwv5tqDLf55
Ii12iZ4o0iXDHwWAcYrFOX6P9/8HyBQwAza5QsRF8C9Pb8QevbO/NGxRBXPeLYXu
vjMkVVx17S5Mpy2lj7vWZjMmYmvynhKFBFUIMayutJilGU/pFRy41EcRLkm9xW8q
c0TpAj0ww3lJ0qqR/E8I1g1dnxkKPWIE77iC2URjFI/nHu/XCqOY0OqcIlGmHnAG
WfzSG4TDdEEzyXA7ztmLiS/yWU/mR5EtkT7mS2Yh+UziBgPiVRQ9MSlmGe5hMtZt
6f4rDsDQjCBxXpfUgDiDHypueCERGVcqllXmQ/dOG9tqwcGmzBtOA+SzE4Z9unTW
cStYFT40DkZbnMiXC99C8xXKUd4deCJfDLKcI7aS7yVyLzzgotZRdyumOaZc/cOT
vYvkOPftoD7N2nDoXbqTL4k6Q6og6l4JLQcJP5QOiHKm2n6vWK9P/0umpPtvOtK5
QI4KCAwqGHpP73Z9rwphD2EDnOvZvUxlcpFRIJs7lXTQ6hIzq2PLOXqQIkfFAnjA
ASNrPKyGVJFkn0Q9ARAn6lpDh1yS8JSUEvE82Z9D3GWCapMGsR4XlHTLslItDe3T
7jllIMUtG7ELLOmita5SdwVTemhRSIkpfAiq2+DMBlAl4xfrFRnoWH0DhkiK6YNC
Gz/XR9jAMzqvY1OsS5eB9/d/A/DdJ4fFOFVY8D4+JEbvI+vuQOPHTOqsTrjUWIl0
vekwnu+NDPxL9q/qqhOCMdRN6G3te3KAh8KfFSSPso0=
`protect END_PROTECTED
