`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1YYfFmjZEuCrW+RwLfqhEnoTpKh9zu6lq5hLVCcFB6SZMZhD1kx0dyE8UhboBULJ
BsMIcK8ENIqb79UD7N84ID6J4HcBoV9CyeGNacfniwgKyrGtMM4vvL0BizUNvsTi
Pb3wPV4Jx13kbL0AjMpZ8etW3UhD3HPXEkq9fQQOgRvdlYFwjrRze/oIPF+/PZlX
N8WoyocgAH4d45FP87csHvvlGEjFzm+4wpnVGEKJcztaWT7PVQumzM64HOdnD9m8
6b6yNPDx8Q3JIl++SGQkx0nB48O+GYn0oaAoul17wo0iZGIEXmtqVEt5Y5VZiuLf
kvEIIy0h7iyl5L68ZwmD46T20fm0AB7Z4nQMvM7Lu1E0EqUNv0wl7vxQzKFLdcN0
y6fWCrh60R0qUKlJcgqaMWvIMs7sILj3OWF7AS2Sx9b0zwsIMJBnL4mWLgJKecPY
QDtUCHKWlkEh9T1xJOS5S4XYxpOKlJtL8A6yvQic9P7kOmF0n+vl7bi0PZ8uEiX/
/3+12mtzOkLpCxmMl/i0YDp3iD0+WOXuB5xfhEy95qCfZSNdp7F4ROxBiMXKaYh5
mwENujJ8zaOcE4fXCs9ugZtmT+Cnr9AofIiygz6M/Gp6SS9yAscRt+JQgrvQiWLb
LT+zQl0qYadVVHa71y9SRpsQxf5L1QkYVPGBbdWm7qnlWGjTvvbySztvlxn4fP49
dUiXfNFSjioeVV+h/3yAIe5UObGX2jJECY+bsbRM5IeZN0sr5Q3yd5qXhT/h3xv+
oD9uFl8atE6qUD8GcK5yEPTNAdM/pf7Jn967hEKHTrgSfy6LXrYEpaPghObulA65
GntgDJKpkHdMVEUpoN3L9wKKaGxdBpFQ9ld/xyLikFPOCKlmhJ8xsOSREMXG/2VS
YcQT1mG+9cmZZwY6jo/oGdXUwgSNUIrFS/yf2YqENwdqpsFzFW73r1SkdYBadyTC
CsrXyV3LEs/UXbsCyq+0gbnWW4sSdT0D+ngcdsyiXuG07FE6JnW3nwXXoYQulGX2
3b310L7G+0nEf6J5ldB4vK8tMKCTe4i2zO6JViUEaB3U6An2vt9b61QIxt6K/vyR
Ab8MlP5SuV8hc/KkVEIXDb3C8gGMxo66Oe/rFeDRenJlJHvA+QsROevGBK84D6Fk
qums0IbMAG1DTKN3qjpdJ/YoRjjouCQuKNhRgJa/pfTMtybGnR6cdXgLQfd+R/5c
h3wAXmnT+/ayXFc/8vJTRuW3ZhHWg4SmdjMjpky+M9zH+P0oLZABDqkTvPZBzvCe
weOuan3aatqWHWWRpiKCd7EEmZRqYhsnbyIpCPZ6f4pymcumAe+9s0oV+aAsfMn+
GGUlf0OihwOxn1Bw4XOz8Tj0RXyWXc22L7sMLyItZdr69IwjcDXcO0cY6EgbGCZs
0trmp3qQxURJKn1yZ+P98NeQo15+7et6Av1JgQ69FNTdADHmOnqiavSyRmh4DEEs
+2ZhW4+3VxUTvHrnTrYF026Mb6Aiuzv1V+mN5g4VfFTwprNPe4y2Vc8H+jbYw+XC
2sMQozb+VzwoXRAGB2VNDRxK1IZkn8Gblwntzhmy4I5S8Ah/u5tTg96IzqDvzhgc
7IefEiPntJ1NKfrimH3emQBQHZ9GWK8Kf6wkGjGHxtO07vwdCn9sjM/yOcOf8CM+
wMRS70OAu+9F5Xrn2K9H0+MH5MF7KA4Hw+G6t2CHITg=
`protect END_PROTECTED
