`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xtqE7Enp8aw2gY6BAI0iFrdAeC6EGFMjD+KAQys24v6O95huC+38yeRuw+vWJxvr
ZZBGHfhZsad9u23HPNin9UoiwmC6TWkSa7t3SJYx+/qGESC/QaQc7q4y2buoH8Dv
E1EtQbA7SLvL9Z7WBUxxFwY076mjq4IhlNQbNrS6fn3BT+udxXf25K+2uMuHrMVr
mPQG/97dpjf7s8ZlF8m8L8ChW9AHNLN754nV90WZt3GlHqL/IXg/Se/vRaRse0QP
pAmU9o2F041ZICy2VvLyfhj6ieVm81YMBhz57fAQQ5IqT5Otiyj42k5kV9WGcqO4
BiD5biSOHkD2ZNaHbvl9fQjnb64bejlAxjs2cK3L+bGHt5tUKJwNMO1GNfM50S8u
jBQWi4YmXb3RFJq/ZHljihtW2KynMRXr1dCANQt2cRj5rLNGMpvEXTHdsZ2MNs+Q
vUbKCYmNHoE2pkbgRmSeHP7/3U2QWm+psGBfVXnRr9saI33RFmsXzLRR2lnNAZoL
8wtr1E7ILSNE40U4GLm0GsMZ03ZmsPJzTMbbwPfVu4IxJv8rStH4uo4ZeUfCs4zz
hnWvBC3YCxEa8aH1Eu9yJUW+5I2lenB6uDaXcqRcd2zyUNZJcOeJB1oSNf/bnBsY
+LOMuJZj8R/yPWWC/SfyB3Np06kum9mkPeTINBzFWmMAhoBXB+gzynovWxZ8MFmR
hajwIBixVVd33nNvdJ02LYIEDnWakfhhWeHQp7GfgPvUhwXR/r8e/pT/mTZw7F2Y
9rVSYuxyqLv0WhF3cwpe7Hcv6oHgV4Tq/RWvBPozd8e6i59C8bc0nBQWNItoEYa2
9rL7eoG0zWKX6VL6E9PbyKSN+wTGtop9uRiNYFP/oQCmP5nWBOGdNV73BNvfiZDy
76mOpZKKDRlCZHdaYFsPej1g/MF5akNucjEpx56NL9mYbbtpaej3KYHw+Yr/DwI7
UlfpZZoFoMALFWZLTA44XYPa7mNpu0KYEH8ejOG2i/SESZ4b4G0zUmkU+cJBH/Vd
1jsbmcqsv29reIKqa3kMWcwEzZ7gkXiklwfCUtqaUk4HzIBYdYx2wkCBEcsetfE1
f6RxIZiuKseoWb3WR5HviQ6OnLasCX+m4TtDTwFWl4tE1jLKPcrCMX9fMim/Hg+G
zAEbaVh632J9TufDlRUglyo7t7D9uBXci5qLPI9E3VKlqr6u8Vb/pZ/rp8jawoR4
uDF1xhquNFtzAnpYMyb6BkfhHxnGmmmwBnzzAp0EgKJIR81b5T1EJ74sD0huPJ75
zSpPugwSij29BVDi+mJZJyddbkpdEaQV5qkWvhsjg0pnBjLo/LwtzcN0IjwtpQaN
Fv5COFdSr3bFBl+votjghmpvvP7JQMNMGrqeo/laXpB7LjVqHQg97ZOflmu3fwpi
1gzL/P7RQYFoUF+F4rcpdo9+wcz7URAbWDJEWes7mX5GyCEYaAkzgL8sPWo4u4fo
Dk+A5La97py4Rm4Ayt42c83tNUqJEOuycz8OiNIfI3sAa8dstdjfmVnZpNvTlWCa
4rft1RKlovpqyBy9rGLwlMXeQ9uXG2skZ7pWNhwjwAJQJSN/B0BBRlk9fkDuFDiU
L5Rk882yq3xYlNW7TWEjOy664rS2DaYYmtCqThgWFnI+W1ceRv9qAm68VEZIy2Ns
/nfbvQoqnV2K+Xj8WLFUeKm4XuRIUEAIab6cCsv6M/HqHnomN7SE5vhssL+3YDHO
80P/SmT/EbxQTt45Vmhx0km7rc1SDIq3rzWLRL4MkowO6XtWgZ+WD2EGTb984TWH
e4n4hG+UUthRdlMBoO5nPYMdAyiYLBpE/FuxWjYyAVv+KVpraePq+BmVDjGwdfkU
CK5C0Vwbixt0+5LUOmKluNdNXCspj9qF0XtVtRU5CBcQUJmbZOEFDE70lbmVsAS9
qiI6rROszrqYzfoJSleC8VBZ8SrkfaS2ITthALcx4W+BO4pi2oggw4IyrmsbfwyK
cPaeLrkO1oTuHZ50xpQABw+K3rIZmtJMgKUDcGwy/YNAujy/aGbkKrBGXqcskCJP
p+LpsTf4eXzM/x8gjxmK/K2FfDXV7uFZZ3ydlB5YN7nClyl/rBr8n9EmL4oBTJp2
XjZw/6sPm9ikmUYX4pQVgTGDeq6GZRWX1CP6XqvQ8uS5qjQGU/zNQ/43goWh1yFN
IttZG/A8/eaT76twf8JocuICSkYOY0pSELqcmfGOqvbfNSXWvZtUY7L4xk1fK3Vy
T3EmaapTk/PFuQMO+b+ZoWMZOxB7RyDRtbCnQLW0j1ziQBT3QoiZAZE8K+DVV6+Z
OW8LB7JZBtrGIzjH6Kb8cgXZo+6UpRQ0JpbsUhwuBbELBjXkBQq7jQJTdkllOEIK
NZAESClPckYdZy5vFrp2iBMr0M914xyNAZ6DUomMVl0lX57ZL6LBGX9SH4w3mknX
gtBpTsybD3QzTBGVkw4JFF7NMi94pgyioKRbTD4qwFfPT+1f2k5YrN5bIBsELG54
Zndii18kIBtmIvIosIXfO7QKu69m1Bf5b85DYON3LA1zWK+u5zQ/tlHclMQVB8/z
sFDLb5Z5e+SH42aGkXyJQRBy01nMBO6fyV//XIhiQtXTh2M6mZBMPUsch0cJA4FJ
7ukRjdPP1Sc0VeJ0ZHqzCzksH8m9hr6cnmTU3slX/PZKLozASxLL0l0/L5G2KhRO
D0/DsSmZEHjpPlioZJ7QAa6wPTw5Az1R4jXgw1Od3fjC0xzcD/mlw74gy9PDov38
98P+tsEpGCjPzDdAe42H/OgyUfaPdUhvAV6iyaZ6XLqMtMrG7VSAuyjTNuRu1j0z
X3ny36/VxXw3XOXLra/SptmE/UNcUrkaYLSfe+HeEVIC0XXAxdO5nFVv//MPj6og
lwGOIUu3faUbiBCA4aViJ2K1Q11fssuF2TZyoNx8iYYZX4UgDghqxInGT7lslg4E
oa8THIIYweKM8fX7e19IKwZiAx9jgg4ypOEWcbjByecKdYW4t9vaxWl8UxwMMGxh
thtcDyIaZVf8qE91FgO3IgsoDt1DdysAbEkh9nviUwv+jsrh8WX+fti/rSWrTIkz
yIjAmyh9HSspxjYPM1V2nQDrxmqSQqtCk22Qb8vVM3+rT0vr+ceH/VD9tFRAf+vT
lQztRRRYnC5QmCQ8i6CaSM+e5v1nS+ZAccY9fISIxJIcZKi+A8BWxqrlGUGIHksI
TU/K9kudOB4ZDBV9Te+sPMR9BmNErIE35/w+2xuy0ZycIKbIsG+D43qnJNhicxB0
qdWgJc/tJ9UV4ZdCpdSg94U+6ZasKNrRnjTuaTuL2fXp8VFLe5fIv+V3i4e9BOKz
61piYYidVkqA/HhhOK74IORgkuq8fGI2j5GKe1FmNZvsr6NLXs75R0kMD42Ga0eL
OA3swHgrqmltWSzGA7N4Yb+hLWIoXl9vtwIuglSqoQeuLHK7MLols8BvCnNboUY2
DdVWvMVnUL21i5WHwzgzH/8F0ezdSWZ5FJ03u6IqdPIIMAGRw2+woabkmEKWMwat
djZB39YZmJZ27ZPB85hXun4eS4q4QH0KOsEFF9mL7IkG6oS8TL5nDtLgsInNPlPS
DN4DLbB0laecnS/bPky5o+DJuN88IjYe9y44FAHAB/jGTKIIDtwFM1qgq+ImFJjN
j8qrYr2Q/JCwF4+NG2e4qaefKOH3xB/MuyXEITE9O96e8iLL9tib+Jrtx8lsnrKw
FDX0gVuexj15q3SkXh3MGzGhApeHe+4rpafNR4WqrUKnpeUKF3HySvsKXCWKbNFM
lSWT3EmCIl5hl4TL/xU/3YCkICkx8lCEW4KEtHWw2ErZnETe1yYaSaIEzSHboP/W
W0LqATYISe5s+TodtcxFSawA3kHDNVGV8VzFLIguaE83kXJNfcVtzCbf4H70wt2e
M/qXoY8ElYz3FkmPvGn/jvEm8ZvOQHy5vfJjJ5oKknnucBzCoaGa6OSH4iZJtS6u
pf2eVo+Fqf9P5bGcyiuD8uxKxrEBIHNxqEurTTshUx5tRtKyXI93Dl3MzzbTB0Rh
HUeOh5CGwNYV3Ye37qR6kFeoC4TplYhygNtOLCwSc3U2UAjPa1h5+XUhZmIMOCnJ
76osRWOnEttZctoFZVtX8ssAJH90deeIn8VCLYV92DrA4XuVK93rntWAe5LAxVRd
uc3WhBlIJ207ywf9H1C+LEf87JOmJ60i0H11x9CzEdD0KjXn+/fwAK7c/HelXYyF
WGcECq//r14ImbN4GQAFbROvkpCpGs6VIi3aH/wKIWnUx049yTCI0lJyrw+AXF06
2dYJU3WElI5fmiRF6gT6qLDhW4DTA6yqbnvEqWGAW+9mIvcc7Gmlx6Qtf6Lri33b
map1R1ohZh7CTtzoDLQ/jmQZyXlBAk0sKL0Aigc8pIQjMbRZ/dVV1o01xQOc5QSZ
ZKYQfsAfOcJXlbmcK1RRgUPoPjsnCtRQjGXEu8ZCGqxU9hAe0Toz9Uz6cbQPOUzR
YH+tUB7wT3WqnI6Q1TfWCmnyFgEa6UrDqvLeuESXTdPHH54nd7YamMAl4MSRgsO8
q2T/+/cLm+Pw15JwwQY+XzkagnlzTrjqDaLUqtuE9E64PceVBps92GUG2hpsyivm
d4eA9f7vJcmP0HOG0NFeKGCGwrsQC+cp0g6HxltcOFsmrqQJq0+JQuQnJZQoTN5k
yzHin0jEN5jP7zsZ7MbZE/ZOCylCN0dgkGNT+pW91Kt2X0oFBvqMmlN5OMju2fqD
QoQ0gGWjtLfI3UXgjmtdzafvPdd7d+8hF5wWueEsqSVuh0q2vJ9LhKMVhSG8r95P
TEhR0ieIGa5w6++XSguDc3UlQKd3JDAlmIg9G3mbT70NPPykS/sVhc5XX/1VFT8u
Ylbs9Rv/IZv5grqiV+u8ZW5yPRYEvzxDif5S9YvZeApSFrQWK835zccNVzQasqu6
fVeBZzrvLukoN7QPXYQ1AzT5auXAmtGeGnmKOOz5ZsA1QwXWSQ22lpP3LNwGevt5
sTAPIfiuRuYbJzM6caS/loNC8FJUcv4DbkWFtRU6Fm3KTcpn3/QIN5iVmU1Xig3y
UrgYWjux+R9wXk/AVhjUydrZmqyl/QYshFVwQcKjA33N3Nn00LhmexGhbChBlLu1
elW6g78a3dvmDq6ii2yyuiOGRa51Iz7EF+ZdEcidvqZGd2ZYDeVbBzA4oOokJF6M
IAoYqyM24UB5WXiwm9couHrhcu3OJ2ecbFHkHNbZkv1KPMISjtDJBFfcbe46V4Cl
Rfd2F7gC7vDj5zkYW6xsls+x9B9Vsxnc1K6NsEPLv5fn7PUtJN07xTwkYpp6JQIA
KVD1769S1wLkrhwofUeV3GWWUNbDDOPnmhobJAdS03Nw6Bl/wRlzoDPCUW4i2jcC
I3THYwWZVqVH8R85kieuX/9ivBf9yzWqW6YAOcIMjtZ5j9kMg2lL0vsCT3KZw5C/
iZJ8LPmkfwhx303iarg/yBb2CAWFt0dnP7tzjfCMtysRVnhnO2ClHRRQXkqHyf8e
MQXkEfoUDW55b1IgA7zJ/ohJtsAkex7Uvq8fCnm95JmS3fgNU1Bwwd4hd0QG0LuX
5TfKh1NObqK24qpp2hSiyGcPD+TUci8eO4IniZLKS2DLUcAgr2FpJO1UpHxRqaSu
Q67pL1kHQmuF3iVEp/AHg7gaz3NiFlgn65ClhySTae/JsBYap11AeOGmN28zUldV
/9SLCzq2dgxlVppXc+WWOVcNc3UBy1aRKNScFZdFq1JWNSqJitq3CFu3ebsji19d
l6PrnQMsR2ehMiOhVVutkYceo+DCO/dgnq1v1hPmYK/GL4eykvBXp5NOwaTSO76i
TRFG+iemib2itI4rdv6EZDbbaV+gSaMfP6f+o8B++9dJl5X4OPCL9Ugsx6W9UbhV
W0KlT7/89WS+wBx6K1LVzjEQFo5Db/LXojDWFnOh86uydFoYWcLFTJgPIQftfDId
TZ6SfG7PgXqfaJqZUU5j56XZRSXsy/yHgZ0Vl+tNDO17DkNRf5Z4LwSltt15UfCv
vp7njf7UIroU6eBvvbeJnSMH7fCDIhzPCtaEux1D43bFSTwpsbsVeyO3LRpB6brp
XGePTqQXffj0YaZfBLT7mQPgLGr2/GDBbtJBukBt+KMV1z6SKkI3eURfH+zbKjvj
je/ciZKznqMCqonfo96WxcDsIcAKtyewyGRvvuCROI/+rxaWLJu73Y891yA/6IKL
11NpET9pHx6JkgtPPvk7oazYfZhHEXJE3L1dL63fgtibC+h/3HV5N+NPIJx8GMLV
TEWBLu//GQL1KhPTJFYeKpCaem3CUcZn+moUw41EHgbLdq9kEL7IEPAEXqpYdcOc
AVjZDLSD1v7ZJY8ow3R9/bAgFQ/OKmWsaPxqamEKgWEeK3IyqSo8ooyAnoD2jbJ6
4zv+gKQlinwLmdDeQ+2sWRrJ/il6cO2QyMtNxzGxuGnorROfKymkyI7dezY+nXdw
GE9+8rop3Yu/4lcjX03pEvm/kcXqen2slznfdAcHjXDWSgXF4PbUrQRHiUDerPFW
Bzm30dT5dQuVWS4COUkjE6puYYvRlZTDt4JoX5Xtimj86NTKtpVAMvzAGIzrDxGX
AJqpfjgmbl/X8hfFiEJiYOQB4hqk1LWlOYdL2SmYkyooP3RPdHlBRLsAmJJg1AH2
rMYbYMCwGjsuktXXOQRevuTPg4rEUrK14vTycAHaZXajEr1zrYDDc93NV2I6MSuS
hKlClkW06CoI/UMTPiRlJg6wPzl4LweihT22n/cVnwFirPot8lWJfGxKXctixQnH
uI0x/8F2srY2MtTAPVGc6MaXBqltxpf8A977z1DyOElzU32lSA1ixe05D580D9KV
WfzeOsbrukvur+AfZyXo4Pu5b/gZ3MDdBbt8iIATat5BUcEB8jIN4W+tLI1YVKPV
q57N0SQnjHC7BOEzEE9SmNxN1ToJSX25HZ91pczODa5bxMvFq/fhZUPXIYjBDMUT
W9+Xl05CYV3ARJ4O85XeEXUS/UlnjeFwA758YJEXg689y/RfkqAtzuBW8KKFUGY4
mqtpnBB4SbYu+/oa2Kad3Y30LbjRHN4BXabMx/+qphPIEIEHKOJ0m43gFLNJUorC
mHNdctC6yuxISP2fU3nd/flN/jsAUS2aUV3LUBJE6jA1VwQNbs43QP5W9UYlvjca
afmQ1DsAb66Tejr8S/3s3CKWDBzoKDb3o4knL6qb6Ec/TwfKvNNLhvnnZ0y8/lpv
aKtkpGUYm2tV/0d0PkHtg37HwiUs31M7T5g1P5vlWhXFeTE+cn9ow6Lrid24o8DD
j7IdDtr926JSTn+H7zLw0Sk3RNzmGUiA6A4GzJfQqXi5o8g3zDMaJi1rNQBoTrIu
6/zDmi0kyyWq1RKuIvNvvYN3OU5S0NM+/iJq89pcveLdJQT5Jn/f6pJpMoX/ovsM
YIFKBs1myXIw1epUQe2jOxk2kg4iWn7bvwZufltH5FoIZxJEh6lS7yiTxhVOOntC
e+89Wgjn3t7FPW5z6/E7Pb65KX0tIbN1DzdIlBbRc+1oq0dl53Z0kYuaeX2oFZ7Z
MmhuuP8/8YMA9HQoN/tYERctmBewledZnCop4ZqKEF0Wmk/QySCs5uS4O7UhmOfJ
7EzhwnqJBZiHdBJ8zeyDHJNI+bDCJbRu9vCPa0vmR5Z1uvlw72nBqzZHOpNnVpPa
n0QPUwFiodP6dnuQwtm2vUnbL0lEtc38iDJfMo48F3r9LuX28tffvcdViNZrqSVI
/GV/ZefvXiA2spdo0hNua2oSeJpQ79HIA9150wvzwCCEnb6vP93Is902EFapH1A/
ut557TdyvQmdUTI5rn+KWPiLXmlv7EchYrnmHFucVrkT0L+LOdgmPE+4y08bEYVA
RUIgiO7Y/z9hzZTz7VQYE2suWx+c+LYQcG+4aP51/B1nXu4/Fn+dmUR3Oqixv20G
57r26Yh5gVnN8oB47PpLY/kFnPGonSYJiLEl2UGEiFEMybxM8XXwjCGH5n7T9JXp
0yXaGA9ATA4e9jHD+Z7iBVJWjTPZ66KUQSdJeCFGCIbZ99bGklcwjB2991aKqw2R
TyDy0oqX/S374l2fbWPnPeUxV2i816o6lEzC+Le3PT6i6f/3xFiC0ZHWFMTKqPVS
i8107R4qIiQLSosA/DFau/+z6PO9I73Vufx8vpqLodxXABe7PpN8hIYa90fyF3PI
PUTGtm3SGrhcubrLf7egHBClIph6UnjZ3N4AxEcmSqyWCakrSMBngcx1VnkrxHFW
eBpqgSQay+Sk/NWV1Y78Vmw2Isb9LRZfOBl9G/o6NqsDFo51sL5ZIctaJxvRxoV4
vPHNwUJ946qqcLiaEhU0oSrtb7fddzawEG2X+j0cIyfFT3oyYPiVNCLiCtGrKc5P
AcR+dnjoqCdHic0ieUeu1XJLi7tXyttVor17kCcIWalwqsyji4Yvo7eP2IBzgP/G
dR+Nixmjv4qcGhyEUKZJVNFteW2oAffroJvS7FXmNFKqQTUQOBLKFGzeSI3xtfoJ
ljHG8FPzJ31gggjKvlGEElU0MFGzPIZFIvo3y56vLBtWq1TikqMlgtCCUwn4M9wl
1URkHLlvGgQ+/pkadyboimZPXLbmhsb1US23DzBRyEAshtbJdpAH/RUJgIjXLCRl
WPZa6aBEbv8VOYqZb04KRMUTVlLCUssDzomyqIaRT+AsrizBVvAj47/wZ0XAe+tA
FDJumdEJqMQz26lSuoE2l8YWXWZVIF7CVf7vVfm1J8OmHG//wVRcVnFf5pFx4YnJ
UM1ZNGLosHQ9+HWXLOB/Jr+M1weoJ6yUL7wIYwVop5wshHLgG3CmfjFEbxzi0HMW
rakDKptpOISYimcwD4E9fMrhc1L5wfQ7vyXlHEJ0sfDHSSYpYqDfuqONsoFkRVTU
7hpV9VR2NaAWU4faWo9uM9QK+xqAyCvOdcp02d5NDvoytcnQfsop6q4+BLgCL8it
VqZURjxC1UtaablvoNwReYSnDndso9Icp5N4UVRDsiL0rfPTqWDT7Al5gtUkZvwq
XgK1UsZ+4AY5qZmuhxks49tQypyKBs5y5SWzbtiBude0u6u4xStC9I/64NK0a0mH
7Oii+poLAIutbLwWfUE12M3lDLf2oLjAr6vCZC1IFfL7/a1wgoz81d4yHvH+XYX0
IgZAIue3KhVc22rMJ+arSrYktH5F/i3SkO2XgJILrCfMq9vpBA4R2A0KPdkmygKJ
nieKmWl7E7TmeFcXNlKAFcLpvyXlpc4WFCpSuADMJYaHYUx39iJR8QXAR/gDmqRz
9nVR4BFdS22sa3lZKvnqFWTQCy+K5qj40uyHgnIVj8p55T/n6OUtV0qNwtmZ04Ps
s1yl1uvhaE1+AzY/WEhxFA==
`protect END_PROTECTED
