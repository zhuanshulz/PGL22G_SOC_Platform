`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gup6jiTvHiWURD4igv1c3fownwYDfAj1UFE4k+F7WqCqaMkoVTIHDTV0mghxJVRQ
Btx/YxazGnf6TOyJ6wPtWnjwHmhq6VdHavR60RCCSKafBKKfDVhHYq8102mZU20a
mLOtYbdGenXE2M/+fGGPJurHLH9vTtxjqVuP5jN8v5fAglA4w4Mv0p7gIKPlSCHI
lcn+VoAQiwtjmZuacBpFwhKDqipF8PDAxUJzmerGjZth7rX71zZfa8PYvJvl69nq
6F8KMnLJMLyACEPnk+dzoR1J5F78dW56LiTidh06iL8eRNtH7WxRIt50Ydub1um+
0ZKQ+54+sZ+11R17IXNShBcCIVKZu/NrRD3c+wJ7SNTtV0QEKCRxXux7E3knWycI
ztzeVAKCSRkmxHHevHZ924adSELNpr78C8HWa3tHNw2tkChuUmO6HIgsxx9rlEKt
ppTgpoUOzG3PRk0IFfCfNg==
`protect END_PROTECTED
