`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tS2L/PILX65anfjvBfnc3SVafjMEKIaSi2E21/b6y2fifVJG2Rvqpdsvm1d0vBrN
ZbP1Y6ZpUHf1FlT0VrEaJp0nh+T2VLc6JLKNKqMH+sbJ0sBxQR0u3u9qEn1WSVB7
4NFSKUS6EfhEfeTIJKpVTPvpZE8ZSQOh63bhnnA+tfeNWUU4GSsrho1VCewWXBbj
I9vC6oBQe+fONrxox55AglBRJ5QPlitekfMy6cRZoVokFwshE7eK9qYdjbyIXqU0
8oJXEfvzaJi3xfNiVJJ9q1fMRL5cjNUlwuV7sAECjZV57cr/E56VX4p5Dr943VXO
PLxkHZF9lJW1D+kdiBW0pDQXL/G8xn30T8iyyWXn+t/DOIUW+ItajN11Z+Fap499
WDdpEarl7xtGoi6hOnpQlpsiEiQHAUdj1Z5+jghUOI804BumiPwuy/z/Kkbt8dy7
Xs/JWhldVJTNQ1otr2VZVCuDr6VKQYe9tOkvSlmMaATWVKbPBlB3hjcOEiHCUOKp
EUlcatjzsmboCiNVI0AMYkSvqnMI4raYuDejgOIK7QnRcy9Ckc8FadVJk3UjjSlC
e9H698jQJ2QXBVszWY5yIZwfa4zkAtfBZNxyirdHwYPFEIIpBDnDAhOak23kZzjc
0xJX+yMqlczTB/7No7+W5ovKkeXcawKGqpaEqkq2DSmdgWLVrzZNVgX4q3TlTiqn
gsTKFMML264pzxnb5VzV64WzijgnDPfVlKlTO78NstUUIj8CfscuI52B4I1T2KZO
m5VdhvxRC8zwC7eCMNpPA/Ggx91GVdVJLQNLlpJgflKvPPwpU7FaDFL4bo8DUdSS
vrUoc18T+goMveDOr7OCdsFPyNuO3BHQTKpjJCJlus8e2JGd4B+8lnmcvJV+409k
6zUDrmB56D2bQkWwd/ixoXFQkQjHSWrl5m4v2i7wq6srYwkHUBkf1/+JITpV5svN
a30jgNzEUv7gNQGPmSbMWOdeAxfobzG+xQ5r24ppz0+FY6IO7Dz9tks5Bid+/OU8
CbmkhQFtQSRiThamNvk+4dnudsf8783gyNc+qQe6NrvfkDc0TZPByDvCZfxTfilB
EYvVyoQCM5wexN0tu+nvgDYj0Ltx6/GFGf3sbiOa751FjGFk6H/Q7of/HI4rdlhF
rFxIwjLIBdLnz4Lq7vZqw/A1q7HeelH253h9Ts2xIA578CtdAZExuwOBF23lH9d3
UmirijCY6vtkYu5C0GX5SFJGUqfhGlYl/q7XDTHINr0Fbd4gL8LjfABZs/wfQgHg
ljRobA7wOxVUreqQnakEvNh5N8gJ664stCsCn/h+8CXOqo66thHcA0/ioYE399Eu
0IkL2KH1oG2gXn7SrD4hjSCnOaMOxvTPJsSwUDiAQgFcxGwYNK3QbmpkFhHMCakW
Vu0NwYuBayZgIjwgKjE5aBpDN1P3uBnM0CD64JQKUlu9jLorsjs4ayn9ERhZ7ZFY
dj16SjgZ2dnFumrFnN2D4vDWNRAjp15IT+HdDO5HfNDp8+fFc10/R5IyiJV3TFH1
jXhCln1+fUnx6A9yNfh/GzSpmo18hybTh8hFpveJQdqKdUE9s5io8WYPhwCTYDY/
VRQr+dqYSFD1xJtl8Tjqm4nbIdqgoS2gpqdoOf9feg37tfyIzHrRBOKSr9AFvpjg
OpIBgpjqobOfa9n5SVilHRKrJvq+cDsLBWJgD+yscEBScwuKSTrJJ3ZJMTHtpEmd
HQR0zf5nY4opHg4rarXzZxCYqbYN4JESY/dgKF1stqHPzukZ+//+vZPQguDZFK+N
Q+WQFI/sZw6PLE8R0v7Iy1K0S8cByA5Dk5X5N0QfM/+C0602tLwxwQwBSN9p5eJ4
6OuFjwEDdpibplQsg3oTu0xBFA5OeQHasOuBxHHYIKy9wwyAUGDwsHcoSqR/dXGq
7t+UhR8btdJavQvrtlLKH3FCkOukvYbmGEQ7BmlXZHbe7UaTjtiW5hFdaSySplJy
HdownRz86/0SEZnLtKksadi80LODzhRRw4zK+gEbnP+9q2ZHbNS7bx2jteayG6/a
sK8cM9z+vSp+4jLPfbfks+7GNVrgjORnRUwEzKsK5Fyxl0QAD+vptHjB9ykklTtw
P12u8/dgLj1gKpZax7WJ2byv4IoJ4pGyQoemirK2v9onN0DJw06yTO6aS8+qamMq
dPcU7AV/kznuWMqe1jUYhq6OsRedKR+iB6CkNJQJUzxcQWGTz66xblbB5JG7p0HO
qykUay4GeJBXvIg9INNpFZSPX7ttsebkQQTIvh7AIqXRYjsXtlMV2tjzUzz6x6/1
eY+3EeB8aPtF3AbVqzT77V25vLHWIOUt8ZAtDSmaAwYoQle7KaHfnBZ1kTSkDAlq
Pn4WxqdrNXlTKTE/Z5a3gXuW82geyHkDUSxiqd2dIZELfjuWuCh21mMAi5xJylYW
30GqnqQrAKVYkhV1rqdBb3F6v7sPgf4/n0lR1mkXoPC3mFv2LLbcAynTTmWzzCzz
iUtnTxUkYEL5ndxnGf5r8Qo7Cuy41LowWApzlhZw8gxPupQXbiz5cEcBTzv+cHU7
rh9lqWrcCWGOtMoKypDv94N5jIFtynm4liMhmdJxPKCOBbcU65ot2dbYsLwSjHcx
J24Eueif1drok9jcAQO5fF6BBr+ZNbbfiNZ4oSxzNj/QL/AOBxbT1C+6YKHIjM4f
S0jiSMdbEyEN/bpeM26WD+w5Ol/ag4R10AmCqll7VvJ0x1hHcjAhM2YNSJminfD0
F0qL6jZBGv4oZ+bAadePFvusw1Q4ByMv0iGskda4OQPwDu9jwdVn6CtibghBHoKJ
oadBMIZdruH4A0G2PkNVPxxy9lzUtj74FG3qu1sbpgQW6yRxGkF9mDULduppdYnq
57uV5QLB5Qo+As8sBJtlFaRFmWu4jm9Xj6q+5KX/CPg2gOBXkqHBmPkT45gSB4S7
9087dG/xuQjlvxrXcnbNBUSc4B2Zxckfd4I+tdWjhrBj+1+4wAVUOjbFxHK86WsG
ERCYFgPrXycDOJqlPmJgwvXSwaWDxJ+iy1aJgZ48exc7OPXMQgi65n+OZmHb0YzK
HYOd2LQVJSS9uLcYyhCK5nTxBBYV0hb3BBjxWnOBH94D7wtea1gCsdc1e+mswGN9
VYKS0AAr2xrZx1864kS0bCXsPq11jmheeUi5aVvf8mX39iWt7dPD4cf+1uomkvTn
I5NVeCfsoKOfhzvEoImy5virAKeyuLkmfTYs2Fy288P1tBOX1nBNw68yLrd7RXsn
s3KcbrU9h1iaWm8BeMOcNG3cB84r3OyyPLIjtUiGNcbrz+qI76b0wtgzLiyvDiBa
2T8SuDkldFmd0307YszmxiRPiTbuPtHaNVbJNiKHY0fxeT5HbkXbKN5NGeOJGcpZ
wz6A1mEh73EIT+mmpGGnhR9v2Ox0bxLEufMj+Gw0wMw+lqQFSp71Nn+mHqeuWIbo
xHL2BfBOJsKOpuMGpVXV5j0FL+aRCOfXjAaOpQy2NPSydPFsfl1INoPMVErIr8BW
IG3DsQkIUvmujwBhyt952JZJrg9glM+mC9GN16F/JbXx2F8cyo/ZP3PMH4q0JuTV
8aUbtOoI5H4fXpeTJxRWNQ==
`protect END_PROTECTED
