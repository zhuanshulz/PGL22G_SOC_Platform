`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wjM+v6LA4YElJGWxOuJzpLfwLJsqmNPUAZFSRmo5/xNZzU5UYNQ8KoEL04CBCAtS
NG5Ur/64jaJ4g3wFA6iApp3H4wYGYywvKdhEj9S3f2mqFTndg+UoO/UUkfOd4CBT
e0P7WoJzBUf2us4bTdan12azm0OSl1blNVjxBvJSxBW6RIJHgav8d4wWy1q55Bp+
brNEUH5iuK0ZZyAwJxhijRZ860dv7/1dX6KH7Be8zDPojinJSt8EcTYFlEB2MfOJ
7zZxCpx6a7kOPqXO8GMDC2eObGVJ9vLD8NfeLrdX8UKDRcGyAtCYBnIXrTmRq33q
niI3MoPt7xM93uIIh3t+FkqDLkOjkfLDngWe5VVVuOa0p02DPG98AkqG9plpJpC5
S5JEOV4SCI4zl+DBgpKDfdzxa3eUiyhh8VeFUFMCMosOt+cnnicf6u6uxq6s1hqq
2ZB+JXn42MNv69sMYZ7qaQFYUUqylB5m/Veu9xlvUwmlt3YMjOSty17N7VCMbUo8
ZYa6vP6ixRiqab6qYR53wChoXB15jvcVpzxMLx4Cw47QJ/AE1zPaZePtatnctfKR
5PeXnrjSbAUBlZX/LUc5JeLo/GLhYm2AODQK0JBu3s4Xm7eGU05t4uUkkDoo73mT
Du0lZfNDSy2A+QR+zD54ffD7DCIt1LnQi0HNMROYniJl/V2bNCkcx3O27fTXT7P4
tr3WY9KxZX+3oCZzMagXPdJ7bAkyBJzhHTC88Ex++oZ3IMqF57yVbJwxr5lxWKWl
aknjL585WjP+IzemGXEXaO/lpDLsdm6cZBj7p8UL61XXrDNNfYfDAnBp1xykckI0
jNBJskHaDgHGXLGESKsfX1ApGwg12OnvKP/i58xKC6fKzkgS2ZzP8JwmJYyXMVOU
JV6kFouDJLsmfcs3IGdD7sRGZqrU0953fCn/V6D+ezomOCVKG9ZuIbpVuU6nGR4y
efR7B4Rfa2alMijFxsweNWxOLKXMJ3SxwVGgbAx6JRuml561LN+q9FN1VqYTg+zn
PkVt7vh7Dg0EkWMTvnTbyHlSk0NepQg+6Zd9lKuQL5FVVmB7cwLMUjFohBOUEIF/
bEkk4qHWmJmuYJph/1G2D+m0ZsCFTUDEMAyxVwJxU7QF/szJSt0lVQSvv9Wl+PWn
hdb4tD3jkqRJYmTK1PWazVfw06wPBBF0XYGz/hJrr6YMgFXfD2dRhy3aQALGi9sL
V4HZ5xnx3Ul0ap7IYC/N+/+lZvGrSGUsvoOnEUPgvqJzsB/yOMa8MqWW9M8U/GHe
orJiflG7sgG3DuUt8+nNpd7Spy1qD6jTNugp8sDDpyQjQYb8QEUg85sAXTiOqujd
`protect END_PROTECTED
