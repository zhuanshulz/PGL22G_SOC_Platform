`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T25tDDsOLOPAtiLDizVh9qrY1T1YRIBwh8cXrb6n1lFmyk8oDhNZR02Qam25LWz6
BkIyH71xVD1XJB2PbKahVq7q/dXgYvobslviyE2YWH/yTbBhi6h+SwgBFOFbwK1+
cCQtjykdlWhJEKtUSLsk8ZOq0DVYJHXXH0cX8/NAUIIHzKF+60vV2idQwl5ki+i9
08mF9NsOUhGluH2K/nWhcS/OcglrKCwYf8eSoaH9BqVRzhCiJiaXa56I9Z7hactn
z5kpBBCACWtmRhIc/l7YrDahFBuIzQmnih9PDVdlPeRN6Hfs965hIZmGYAC/xeV5
3CKRTI1lAcPoaOf9bbnSdw==
`protect END_PROTECTED
