`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iGH3ZI9T/HaLqPJcLLunZ3K36Im1uuKhza0UmrMNVq3H2dTYAikCAtjQVHk0gqaN
q9aCQToqoxfvMVlULVsmbEm+6syuA5XIWg9aCQ6go4Wz2kaVaxE5fXl9jXw440mm
iJJms24GZ51oh4l2Uqt84Hp7RcWdVaY48SsKNRqekGG7URet1XXkrVd0wU8lfj7g
OzdhSAHNURUwHIwu0hBeY8h0WqOow5cSs1pz74t9ODZs/SvhePs7lZCgN1RrUMyZ
gMa66eAitiyriOJc27rsuH+XqiZO/M8q/gMVucFUvooTE0jWfX3Q3IQBetj0HnUd
jqrJ415cplEwzazMgQlSkLqu9WM2uKQ/Bg+GbqBcQpGx/4KQFE1SDyPzIlxkB8Gc
Zf0iq/ImhscBZT9Wtv3pnO4s4mA9LBrH2IzsBhXkjbqRTa7cArdC1BGQRaos+30d
XpW5W5y+kInZMzjD0FYyPEbk/QEP5edm2ESKq6nxQTN4J/Ep2CUK7gxgzewsSA/S
xO1tcfkDDz+vifcKyfHGRCzgWolLoYlH7IPFS5kFLDFct+oOK/b+NhJqi4LwNkr1
JqrjJYkPzr0MKa2bkKGr45AcK+2dx/99AbqncQPlT+XEQVT0PpyRMLci7LBn4/E0
95tlk40GnL+ZGygUsSC1qpJLr8ZbWVmDtPS+DkLnmDEXQQglYWFY4iMR9DBPOlSx
icX4QDYKTJsxZE3hQfXQ2ULAvaMqivqPboGyg3RjICY=
`protect END_PROTECTED
