`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5GiTRd6RbQ/uz8Q4aKileFuKogIwaFEdJJR4wB/7xgwIR5TC5RadbbVDHJmVlbRO
h9UUKejY83DE1nVpn5ARs7HEPVCgQEN/Yso6xPlWV8fFtIl1gfseQpHtCKmgVQMm
rUunsHyLMOjtc2mMVoMwU8ymio0+HgVxVAtCbURUwtwKnOxzgwf/DV4s/Kf7pNbn
R6h5ApBGCQwPvFZirrKMF1j+Xq8+YnAeiOYWUR1puIM0R+Necfmcra7lKdH5Hf+E
xGqYZ6jfh7pbmgsQZSMb6kYP2kYASaELUB68oxwNwLkEg6zL8WjvL+sGrqWc2lla
y0+L9K/G/Y61Y59d0oojnG49zUjTsYOAZ9ibE2fQIuxhA14vfrQl7vanxKzP5u46
MGd0yq6TKLOMYj5bd4qaY7Z4nOmrff6R/iVZTQ5CYCk0ucOsw0cnlYsSE+07qZEy
gEGthPYNaQkzHzTO0tf+9u4G6NQBUEl1zgJaT10Sxqqz41OqRjEu3DvnTN3JVIsi
r1vFUTaMlb+nyC1TPiSO/qqHwr3L2Lpp7rUetLhtbv4=
`protect END_PROTECTED
