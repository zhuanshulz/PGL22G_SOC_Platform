`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zs5SemmbPEkBdGZAIsS3xsu9MyHDJl6thaAnX5h7bv/9qdTrgEdP6j8noBgb72lx
OQzXmKrX/kVV/HHIDg+A2PMGOlfPEDshG0eU7af4eSd0J+OPxe+yIt43yc1LQEmL
eGkDsaHqC9YG+9JfesJnpehBGLCvOUIwNgklPgkFpLJ2mblzBhW/3ruXGo8dw5tK
NECgPM0CBmC8xOyxEokJu3F/PhicH6CeeOEioMubscfFEs3kvfhcbTOXEiHZ8LIz
SmxaljGwaljzQpo+qY51QO4lQY38MsmNnE6lMiJt2VVzs672EjtWt/JAhDtI3zba
Pt/kDlZY43VDDlAAi8F6h1Y2Mr030Xak4FX1UUSnVrMMrlYiLfj4F6JJKho74WIx
pH+28OyxS9b627EYzpPNuTBd0vUM98OXP8+L3UjRAtn1p3EjAZ5qqYSF/EuY4kLB
ecwqV3dya2C1xFhBlUP0pbQAZMQLQTdG+Wr4uOpiVflZDmKZBqWWTs0XmzqhLUTN
ES35EK2otjjWQohgoeh4yNKHcHyu/nADe+swI1qvYVhXFT0rx6Y3GyEfQ8S3O1SP
c3QvJ+fCV/a66+6lSahaIvv+8OpS27y2QvEwnbOZxVcVmaOIT4yCzEClXTJkwBeA
WtKiXzfPoM95r0VXUUYZRApgagJtcGzZXcggKj3MrWVea5PlzwpnVIGBkPcblf1e
kMsggNDlOzXYc2Osn9Mge+AtFSYf97Tvpzrmp1u6mOJyyq8SJuICTydgTMOFB5m6
vOY55w7IbAnxagGMloPHWSZuBRlYB1q/1nXz/mMyD7tyTunrh366rAyO88p7ecZW
KoTp/pyERhL7z3IP1C8ltKoFyMh8ExeCeiKYIdnA0PxewTJImejjOLowGWX87lS5
G7Uw8Rtpr3d0eJgPIlI0UyHJlt3Mr1DAg8PNtpvDZl54ijHpJr65PGlLbPQ8sE9u
vV3kjDmp+AyyVLdj9SDOzFBWagDSbv7lHD4d2oWrQJSguI8LVs5PjvhxIizGU+/I
IzyJosw2A0mdpzDkiZ/RcUzFiHPjbzxnNxb+DEg0uzicwZH1LpfN6dmr2DFI/1pa
N2Yi4JLPLfhc1snQI4Pc9puP5QKEWnNCj3TgwEi2XfaZKYQ8Jo/gF0s2jOJ2o142
IQoljyxs54UWk3sc4MBxsdUEmrLekIVd8rIZHR1AnnXq2x5Z6tB+eb14G1ThloZT
NiLFszlrzXwP+hd7QUyOuKnXq6RoOd+oWjPasigxDkfUwjuUR7Ql7L/arQml980M
ZFyiICFrhBbrI/KXUP8e9aT90MuB5e3pbrhY4kAcI9ItegPMCvCUvSk/UJE6GVWV
IsJlAn5IQEoOWgQTWHa/ptp4+aVQYsd44naX2gT87ZAB1PawAqnVmAq6ex2BYSLB
IR/YaDm6/my6onrzVksRlzaZsKmkWGX6pnuRPky+UaUBy8xI7fKjLRZorFrb0NFO
HRfOCDscCvY9gGP8kWbzJXR6vEDpiHRLJ6XIexTeHYRuuuD4rZ4PtB3XJNpZCo7L
N3Kz7+nE0BN5ylsmAEuuD6v42+U+yOVBwD2kVtQFTHsXLYQQTPRdby5KjnUeR5k2
oKYcBLlo0SZ2n9Cf7TOde/M2KAgsVKQGvoKBqknou7luys9ZAdIYV07SMeVy5O/T
jAmeXeoIIK2EKus/oKAAcmv/KQglJ8foyDz9CaY3Fy8p9QSaLlZ92ulO2lBNtmiU
`protect END_PROTECTED
