`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1HRbI1pfuUFPB1SyfT8mcJedgsawI/sgZL7VoRoSE/zvn3L3wCPK3T09aQRRWED6
U3ysNr0r3YYwmMqeUcFExzMq1DAz76ku86Fm/iOzK0BZ3lCWycijgb9dKpo4ZF+B
cZhKKNjI/5p7F6m6cz9mzt/k66Wo8NNzLk+gNSCvkc/c2cHhpAUx0d82TAtvx6NF
8sj2fk3dcCzwrj3D3eZQir55S0jPJDizfubcLziHfPc/ADUVPDjpbNINYZK8IDA9
60oiGN2m33X+0XHpp2QMuSPkYSORO0X+3Ky0OGt+hcmgvu/CrMV735F02pZ6dy7g
m+Jlw2mNeAmugPfjqyeYnl0ig2V56Zh/z6BbnBo0vAW8aYKC4whd1XvpjtyrPPj3
+t/XxFdj1TBFtxwqQmv2V1C7HJkqio/fYiMfk2kGOf1TV8q1Ry2oKHQ4Z16FT5xc
guxhiS4qCcFguLufp4QZ4vjhHu4arpHzq9rd9pGZMZOKmv+nOeKMaZD3LHa6egXb
DFsiEJPQM8wk9Q4auI+43UsIYRpwT1s2v5rEJAhDwzVNZbRtJAJ79paByxuCuATF
0xLu2PiuBlRMyy5DBRg1DNTmchDw83/vJ4hdo5KJv8q3qjSsRZaK/m9CphU43Dn0
UPRUIX0IPs0ij5MdtiDINJFe6CqGOZQzl8nzr/kWoGe5vxhqNoJdKKm5e+CwPYyu
O8X0AOC7p5aPxqcS/9oZnlWsRIc1gD765FqBADzEc93BlLheAAXvKQYagD7oBRSn
RMqmpqCH0/vO12fQE/GYoMNruvco2paHoqYExQp2whxgeUoOwOe1aCazzHLO02yY
noxPw2HekzgpnNaQsxEpHtIXhNLB5ma+lXrFlhDdrMeyOeGFjpziFCsTByedCBOZ
79G2j+XuefsMApL+r0Bp3oF3e0EUdzFS9MZf4sV9JqOJU6f7dNp+54Dx5DU196PB
vONg+Yz7aqUwKzgjbUSOx/YyEX8MFv4gByTVA9RzgW/c/qcVGqgsJwXSHKC2rNhZ
PPAtJA7LZo+YHwAw6o5Pz5BNLUcBprl50hBqKUIXy9fNAm3UUG8zPW18XV7g9lQy
EnQg0Kf35J8KuD3GPLCttZMq1dSyKaj94Sx6cgO461N0V9JzQs7nn1Z+pETjXtgE
p/CSL/g/TONcOjqvXAXYDbXoMID3v0ZvBuDTHl3C6uOolQr+pSMRoGE69CYZftpU
bKaAlKmuFRXhIrpcndMxB6Bvo5OCe/1TlCtJWdxJfCN8JNGO4ojhIfJHDMOm52Rb
Rf6Gx+kyAHCU7yFzSx4gyKuolBezzuigFcNrmb4SKL5djnOHNt8EYd9pcUYOQ6Sq
YzaW7XpGZ11GONhfTJ19AD5RKdySjYTFdJx+IgiXIw5Som0emsouYvPFkS3aS+M7
fcrzUC1lGI7ubjEdeOuaEbBb53Bw4po4et+vSxngkmUdKrh/cva731sTs3ocyqxv
QhPj7F6Yed0y+4z61JBMErVQgWLp1zmQm/bYVis97qfmtBtVznNYzi4SBGCWC7Wu
oUTvYfG5KJ2UIZHvFqwxR8J7QLwSRr6A4wJaSQia43kMONhpqmTbzAfk+w9lzgN4
0gTQLw9YuqHtZ8Jumn29LrRY2oxzXYigHcH4n+HeyiEsOrh0MfKle/deNhq76Y1c
0eEsKC0YT2orc3e7OpKsmmOhn4IxMgDw0StF5qINi4UlyCte3QZy2Z7LevPqmQnb
9QGORWn9srSDSXg0UlLRxsJaoDy1DoTsdwxseI7pM1o/ysuNE5DNIQudR224nbNv
dAB6KLchrtY5/JwBgzgpggWZDeaB1KqmY6krYkdwKOpHOJxmdmYyQfCuvCMx3+wJ
9syqO+FRyzwiGUWg7Ax4LC9c35hdyVSxikujcPM8e0hPXYeM/E7uC3YrcrEQ8SRE
zuI4Z1h8GYjCQKfYraVpALPeEl5YoznOFOD6eFB332EUioE3CWgSjEp4FvYAbIop
v/2LfI0HF8uCXirSe1BMt1gs579mWCDL+MBHsJZyXbsCbPKsXnudua4WfSaBfkdM
pl9G/VKvsIAWZF1vh8znDcvzO3IL/gsUQEG5nTemCImN3B3NZ2FjZal979vhPUib
RcWze5GsDpjov1r6qtcaSnYtPc/G3WqGxFyoGGT+N7Y2PfWkh9p9QHVVQY2UFkdj
1Y2k3mBIztDwE5STdzhSa79PFX4h2gwygnrde4UVDxSNVhChXibavVThysr0jEdf
eGYzr4o/5bOawVv6JyvSjvo1UAtsg6Z6ceoVrzxv6hwzz3cU8H2Ys8+RAEq7wDc2
Koyp9ho02PAyN6qV6LEdRrlVCjB3xueSTkGifWG8j+M7/8HiuhprMsnTHSdSgZPb
xqZEXNwsXsSzplJc+e7GPo/yRCTywn+X6jNNh2vq2TgiFkXyU8WXQUO1hbxoU/Ye
7N4qJiuA7RJKwZIVmrHz/KXhlB+LoOeSgVeZI7zZvdm2PNUeCLdk5V6/9cadZ5fR
N0DZSEHVyPgY9XB83V9h7QYDwjz3i1G86LLGOaE5CRzAjZ1KzFKIctiqZ9bmdUEM
AGf80zpqw/LtX6ePXjeG7y5gucNJUjdeC+q30l4ifKtJKPISw9iF4NcwZvhw4f6Q
6r7U9krVk/N1R85ueh6V/Ow+rSZ79REarf36ukZntvujLPT++gzyrhWVUlbaHjmH
tV4IkaEm4WWH2apXL11hoJT26yICCmjay87XPwBHwXFHC4nYfc68pakmY4XuI57u
gz2y4Cj2t/MLDnVFCmrWLkQk9BMZyGQBZBIji39I9krEbP7aUrtHiKszSIqaSZhx
fZOzHhNemOaxWzpuqCEUV0FDpFCXihUMX1ZJJHtL5+r8jIZyUCkj1v3E4vE346W9
pqHYtfNGjtgdiUeSnNCp7rUVj/nf1bWxnG08NKtCZ5jLCyepimILslQp8GVapske
GC50A1GUdrnAXt6toNIewWKHsjdahTfBTuaMScG+hSpFtfhM9HN3IiIzSXBSOJmq
TL9qjTat8WPqxEOcCBNk3YN1ejvCXaHmR6LwvwLuPJTh5tYuuu7aX+Y1bJKBlu3x
HylmtIhNJ8CWv0KvlT/Vhpc5hg7+EQj+dba5sXBC5IdQZ8T1LIg1IrnBpxfyTuXn
GDq6ry6Kw+CRBMYhSkrrdlcdNXWJUmxE0ft4mMjh0MTSHMbbztM3tW7SWjBgxHc/
JupL5irgF8y89JqwjGEVH70zNf0IIKDYDsx3Lu1m2DRyTNmqjR5Kf0apGHArARn2
SnoGwk5eEVHXoPbeazvCJMbUIWStV5tHZTRscNVT3fnvrCxFqP+hIMd6g5mexuIq
VJtbxKs8NTrac69a3TADOg8q997rl9WXy0zlNssE11Kvmnr9uwy7NliKTU8OPnKn
Z6B+4zTexl+VPj5MLfcoh5zAGRV05RN2QPRa7/Udy03d4sOagXIJ4cXT2cqQGkLO
sr2Toc+5lgHLppAlyXg10w4hYE2CBUdPbwX4iT+wtfh3JpNJ2u7Xir4JXn9RvdqK
YcS4YCaDaajLfrr4ZYN4t8h76kCAzsqeZjgiLBlKXs5AoZqkkoxMXeE3evspI48X
iYH7eUNdh0CWlIQaKca10Tduk/VbDMDKf0rxKewPU0hieRBN6UAoaBOgESuH1ZnG
vOVhHUyFObjQEt4wqUDbMHHzCKVMebSLaMec1QWKWj4mL91ekHHcbBJyMqR/ha37
gmkzDYUmmffwjURopS4+TU6Nb+g/80cPanPRqj/QugsfGBFnS5sNdrCfDnfD7WWP
`protect END_PROTECTED
