`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tse6XcbFcANu8RkHuWj7qpX7wVm+v+iN9M1tlOiXiqDahxE1ZeuUpuNzz6fnb3Ju
/Xz6oJXpXn8Tie3F01lazwo81xSKX9FPA1bl6Ba49ogxsU9WQ5TSxfsdqvhsaq3O
76xf8SJF5+5BFEls1JN/Ig5BjnFis0VTFVLoWaJGw2QqfRLVMzxT1vip2IuOD5cd
Nb8ZnLVTCuJ7F1HD5DjMcpWrlolBA8YIs0Hlr56tNROVDYW9iW6RG00IlMPY8gfL
28ZMZKizmM1M31esEpEZYpX5901kkDtWhnhIUfKYu+a/uQU3wS2r7pPx1Kkl+Lx3
y7emqCVHpxHKTbYq50UsK6QqKcdNMmk3cNQ/pP3R2cw6WGk/TIQ+wtCxO48sCPjk
P1drNdQ2nA7MbnP9+zHgf+bRxECaXsXSc2UD1TdlJtQod5HFyvlMqSwkn8h733eS
J2C4pxg7avCOv8dNhMC1DX0BRh5otY1M4pPamDksD8fAhyK1wphYePkYZ0NOm+fN
3b19FegVW96Ea30CIY2Z2Z0efL7a6cW6mdvfedk6jCetRpSDV6mXz9LguIFalMfS
0pkW6F4fO4Xnx1wj/BqLcrkXQOeXqbWXmeTwx/RclVQtt7dYImISwbOdZ+sGB3lk
fYXCLSMZQJCbZFj2m/Z+3OPnwR7j7GHtUSY16FlZYmr6dLRApttR46PsSsXVlEbA
vRDxjZXjOemXYLBsmXtZ8Lv7njxwpVZUWZ5bOWoDOnB1PV/eySU7CzMNuko4uxuU
1+aGIqeuXPqN7PeZ6qMa7Fr8I3LqDx4QyG9NApp2+iuai17jBYufpp836kzfLUsG
9iXLEk7AT42kF89E83GFzg1HMTy1ZLV+z/UhcHxHNPtuqo2N5gA8dT5+xaDOy8gg
gQ/7Xl/rxuHcLb+hTSNHhMZ92/17tlLgrvPv+G/NuBUMzLEFCHMnK5irtiCkRbw9
bkz4eyqnPGBpDWcB4ktP8zQgVZgdEFgsO4Yh5wcqFI7RkxCDl9ZLu4bVQwtyEWrA
ehioIkmYI6hvOl3xZgmbChkFJ15nS/xt4z8argNStHtzRklO5x1o1VM50X/GWRlB
VZgawE60f4ca3QwoF3Etakfje4MyyTAU934CCd6V+ABFNe4RaiAJWXRvJu94wA1/
7+GwQSdFdNVWQjP2Tld6A++PL0gXpc9hocf0l6zJCj1F/p+ouU+OpD/BNE91OCfu
0eOkBAdwIWjLJG8wo84QR7YZsnqcsRaLkcJ3WkVpMuDX+RSIfe7U0ivliYlO5kSE
TQMr3sJR0FqeJ7ADEgPJz3XDPCq/+0uHEj+2iP7/7V2wc6FCjgTiaDjIi8TWlPzz
HxUabyJXQxK8usV0Lzn9dncZyIGGlp0y0wjElCypYwkI3sxeqgmYFUn7uGrhgij1
/1VouOW4M+Efgrc1ZYp3hqepFzqsgS5HEBzgGxoprjqAVCaBZN0/baS7KxsJBo9A
wYHSt//8XGxsDco01hm5bF7f89BmpGwApZ5ranuNDpodQ4G/vUNk+xryBDfJotT+
mlhXQDCz77GUcTRIwar0gaboQuDqQdrqd18L8fqgc3YprR0GW2EwjzpXUcTcZH9s
51n98Y7tuB2lPd79MgASxWPAA3eFAk8U+fh6FDcyMRJ2jS/gCR5YbVOp0qBaiSGn
`protect END_PROTECTED
