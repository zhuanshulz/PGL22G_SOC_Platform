`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DBSLV6oiM+dJO1oXcgjVuj4rJNNPjnPIPpHBDzUtm75AS+sh/CMKhqaTr7IJ3AIC
Bohu8X9AIw17b7fZQ36LBgFnuhIVg+FPvHsejUACc05P3ZXfXvUYe0iejycW1nmA
IXmL1YqfMUrhZf1EFhtbjiW7l4DmaSr20n0CGsStuTNw0Yut/PM8lnfg/kh+o0HK
InXe6EhckgS7xzE4J4i9SUws+8RUJFWbajU/LL8oWjoAlki3a1RgaFcH944QLRJo
w7SWxirBNGQ5P+Rm7LYNg0KCM6lWLcj9fXXXlGWN3LwpiVrsA5WLAnjsY/XJzCmB
3RFYAu4DyDDW015aeDj2v9Vwh7wzZuffI1c+8X9vKtJNV6WY4e2w7fpuN0tl0e28
pXHYRIhLa0D1zIHhSkfHHsHMoxS1PEKnh5yVujO/BU742CIYBr9oTcLF08xvXTcy
HMxVmTFkCaI9WLh3x9rNmdRUPrmGXvRr0Egs1qWZJeySXtRXvwmbiFIfCEq3Hr8q
+tKiQ50cm/9O9IxTJEmvtYhhLwcRMnb7wy2NjmfEEKcZF9wZWb3Minv/+k3K/y9n
Tiw3F639N9fywcqmJsp1qEcUdYymUqHOXfMDu1lzu/ugDvnsKisZWfFSA4KkG3KA
jMNu0+rY9OIKoqg2TWTKFOsREgLzkTui2EIQyOY3+nBqDsSKXl+9Djt1yL8LH4rQ
SZwOccf3bf+3jAc8kdCJzkzyEGMvX8x1aP+ZVa2b92zcJGosM3WsCPPonVWKX/H3
RkGSM1/u+K/67VEbA4uTx3bkXh034XWJoksh3UIKqJkGSrbekq/LvTiupqmaQ+W8
D1WB/EnBQmeDIq2ST7VhoRRCgmlnXckyK+CvH/G4Qu+5WoeKkBxeGkBxVIxt5+pP
foIizRwsXNY+lxdmoo0amZQ07cXwh62awV87fvLQ0NWDQlGMNp/M9fgwr520Kro9
rOLAWY92dia13imMwXPXYk+TtjX9YnBj8McOm52KAHsHI/8Os8t3ZLt9C0vMXWyo
1xY9OvAAaxCYE+0ZS3tbsGGYzyDIyR/K227/1R8odVNz13oxdHVISF7yoo+V5Q+y
El9QvApChXkCkl4RvQeP2RZOPm2BLtnDwb8Z3p/y6Luah+B6Q7vtXT8ijktOiOKQ
UfJRsnG8KqOzLLRJZHlv8azf0Bnza2y8qRT7AHt10lmu2TcLqO/YlWBnhAsSWNkf
jdq1GEwA43xs1gtrngFxsrJW3WedV4i/IHbOLZy22ji6pAlVbUMmd+wVX5+FDaZ9
wq1WSblGXKyFzTgfeWBqDiRw6PaKTxcs8TIlVN9WwGCGE5ljJQiJfh6UPBuy4AzD
NMreGBIa2YPmAN0VoBMFW9ZpWnnWVvzOI8YSnpPUzijQxaeX2dGGIcWsu/YqZSDH
pbAW6pIQi1fGzr1FaezyOMVU4UpZyRPbeYcQ+v1gDlxxDqwo0d1CXley8NEXB9fO
CB99aOWJtiVjQqT5jfr570QKR99wXv9G5DWRsY8ozUUUtQJH0kGhifpQi0bVcYsM
mNYnqE+YUPVgGzPd8ecmD+hdjI8hmdoyuJ7W2p1usqPBVid17zfZy1AJ2kgmWlrQ
N8BQreAbT3ttntcFaVNi7ilXFLAhNPk5yLwzN/wiP+cr94+ExL20p2+9pv1VGXMV
i0Mt/Q9QXWE//5QH0eUkTR6elYcjytyTOH4F75TmfdHRbB+bAley6w99QnwpYGGV
Y7tPADvEBugftIPi3SEcxU9nXsom2OT10h7bavk7qUFsJlo8CuuOrrgnehuvNoMl
Fe8jbKrdavktjmaa9U3Tv66RufKmriy5cpkFK6+iojAD0Wwrnef1QFsm9oPYK8ko
ubrTqYBA5h8/LEIesHUdjY2dztzbU7ywi5kPyLfQ3MdjhIeHfNlMWxpmr6cMqhmn
v2uP6RLXJfoGHRFvXlbJHMsLrDl2jnHPFwANMrP0eIoyCR9fm0Ubr2vriASf2v1B
FUTHd7TzyiVhHwJGqMWxnJmkzHns7lA7kUdIoFTmMP1fLHRp+GjEIMWvRYbabL2J
V3YXrg26fIiHqzaV99axvM/hWlBwOaITFvjC9fSnnm0oODmR4cp5kTxVQPLD8C5i
R8wO2A1BP8yDnQGH0vktKPbSWu+kSqisTCU3Mh6pHpmoF8dfLErtBtZsc/CciS9e
+5aMl52KiODB6+i8R+wuCv+7jtmbA9jbQgeXrAeJtNEmLXyM5iibbYHdYXWxhUqH
IGli7ryCcehdsZYq+/eitBGat06vBNDWEdwC0lcTBGgw25D8F2uN7LmIBvMryh3k
U2BL6Nt1wpXjeczEZxx0h0yu4/At/tL9BB12Dyu8FEJoDJ+nsVkhcfMneN27KyrB
xNObSwN4qfD740/BinEwylFDT3IJLHgiTclyoRbDze7WViEgjMUZiGU2UtneXiDv
8+Bss4bdiVKoXxnm0p5EiPMmcwIgq5nUzrOR5saHlCB0Xi+0JKdCQ/Cs0hNUIv+C
0ZxvzjRYXuPaL1r3tu5CNTgpktLQqh91J6wvDHRypEJ1zxCnPzDwvYecpCOkcq1Q
Lw2qo6/eYvccnVcI7XFNRrRPKM8Ms7joUYkIzuR5w+2uP1duCxDKrd/HFbUNz2ok
NXLmB2jlBhZCC/YNRQhAVGReTHaLcozds62/tUpywAPFI/9DFwGfh5/bnU9nIQh1
zngpsW4im79CZwYPWPKATZjLr5wUufCcSNl619we8QvtEgEcy/hxsHoI6PiXdSAf
ZjQGihisklWcAuM6hOKQEaG5jrOiSvof5C5Yc4Y/uoBKReM4ULQeQIThfwOqn539
FsBzxCivIMLdHhUTZQwU70343qGvX5OKC/ygEy6TZ8t10nUX0j/w+MdvIdYDEADn
Hyg/DChKUuptlVVr0iWL9VTKOA9oDxa8jrI/NTE6Vw/n9iZYWIn+BrhW4lUlvDSP
S8uGsLYm3eWe6SONQNWWW4ZOA0qPMP61CFyH4DpxGlSTV7uB1KhdgGaDJCOTHOBh
QOG8UMHme7GOg3xuwkrlq31oXywoN2ZN/+91XLov14NHe3aFjNMFN2lCB3wEBT18
3t22XPpkiy0Pb/V+2y7WowVJcImv3bZ6Z1nZikxNScPRiUZPHySWuXpZFxXbD52f
be/KBRjsrcBriqPWEh3yGZuGr/tn1+f9sCH+HO5B4LwRXGbhIVOwyCloDyq7K1TI
oBOkzV0SAKj8wuEuz4zaTilcXTcHeKKZOPDGL4kQb57YfFEfLEnO4PnqIEt1bwNw
/ET196mPYeZb0E6eodKmtkqbSczP0USHXq27RP+lOaMZJsGZLExxJApQ0Nsnjgc8
LWX2zcB6IsPuv9eIsqQV3+JE0R5z2HYcDK7SIW3KdXJLXTOpm50IPNiSsBnIiAPd
Cuz5s+lEnbf2apwlX5GYNnxJRAdSTGkrZjAyihnzLHBUuxZOCyc7/5h+NhUq5KAE
GcTFbVFhLx0B5D5c2B4U29VletSWIkBnkI0fXwuGhr/b4aaZV+fXcxHu0FESWEgm
YD2MGCVnGDhiS7ts0qJksBolbMjnx0zwQi4Pzc5qUOruISgQtu7VJ7wvDb/fHsJq
ZOU6vU96cVc1Zk3tamm4JJDFwPfWCo/By2OEyLKBRaIeC7/KruV40518HaYBxXF1
bOAU5YDsp7ih7m5N0c17lODMymeT9IhlUu6LtzFdUuV4MhuWWckMEyW3qUamMRhd
ZdP0MOnY7ThB/Ehj2NkL/PbAP6+4lBTgVwghEBlcukU81A2E4Q3+gehcbUEs/nlI
SL1eHWYYv8VvyS1YDdVzD/Yc5O+J5DR0gXmz3kCCAna//15ynBRhyzSxjvrDhHvd
dXHh/g0DIDYm4JGXj2jKz3ParNUkawc16xUi4xhuGlRDLsY2l9vuqIvIYq2LdD0G
6G53rcqk7jgC2n3mjQ6c4E7BrLLjGfHiNj87BX7aOIh2Pc8DO7fS6GxhHfQpWvZb
Hgo5hhqo+6cs9FWjrlPJaSAJPcsD04156eOaVzuI+Vvs6nzMfnJ1LtIndZZ8/r7b
zst1JE364ZWR1YgvGjXZJP3MjIW29g85sL+gnNKWcmQ/mJQfu8MqhSzJ/ntbdITL
HHWX7BAIiLlQZ+mUasMCDDGu3r366Uru6O4hfpbBdQ2fFpkBfiG2uN70W8OXW2xo
pnzGTyVZnTnihpN5fFh6f66HMzPEqMgPSg8v8GyQjMM4wKrM0IAZdlraDRxjW17z
kWxUfLrQxSirR/ZPMG7QmErx10SB3K/IbnuwbQBtIrjvIMdUZY9sZSKWND1zIaXz
yfqPSU0RyKY9Tz8D7bSFr6ca6OIKhgy27Qgb3rk08+a42x59LKFlGJ8y3d2VNtiW
68VoSQHDxp9VPUFAnBJZhshbopCf4nErbZ0fu4CRkw+2f4D4+S4brHQYHr9wgnJt
rVVIEKWWOdLRJlaSbd26xItTkrl7gOhyDxJh/6rc7sp7S1nDyBEBsNt5BewA/P+k
EM6TZGHjY4qlhXFqZcuGNW/IupBVlpQGt5LoOeS90P71h0+cOaZPtlqE7ispLxIT
wr3w4z5eB11RxVS/QmYPsWhGYrJyv+TtDewxdl9vqTxiphs+FiVnQ41DJ06bfBML
hsprcT/8326cAM2+A1eJCyVwraQGWloNpVBixQyfnEfAeFNLffenNrchFny+4Sjz
MjKMk5OWFDvvksfPaCw5b4oi3VFZhNGvwM19v1I4rLk=
`protect END_PROTECTED
