`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pdmUlacuTNdTFAfI66MYzotWL2sz9FkEN4wmDEsbkrYOFxIJnSoGc4D7/avic7+k
m2N/yhyFvyW3+Wpn2VcNAvD0mogLOHxLRtlr2Q6pFXlgTIr0Lgt8sQrqIFXQDVOJ
BkvqF/pehV2HbYXAI0hqFhpX9rHEAfcHQrGTOFBxkoPR/6CvtH8Uby2ETNp4L+xg
xR+LKZhyIrjCfFSTvfPr6h5N71EukCKe+7oQxTeN2e9JVmhohAgTPs8aC02AXVRU
ktAF/mTZ3MHVizxzL9fc2YKiCm0Dk7ZbokWgx04BmuVSumLo4yh62FTrPoIXIcZX
dlnBmMs96/64vt3uvKpwLUqeYM73FKwkKK73W0DCf9G8Bx7aVp4o9XNZxGhlfPx7
rXawo5dkKPqjgyLa+btFiZUlr/qGs2iTszWwSoqSIpvLN/73qA+6x2LKBvY9TrtX
OwYLETQvoAIWfAQ9WMaQAR5WpXAgtUX2Ed4LiE54FUuEMsNWDP3Hcu3uqK9N7NeH
JL9hFxPHEVSBMZpWCPF+UYn/BTXh/nUf/ukuO8/KgLCnG25kvJ4e9wfWs+yQ/8E2
cWZhIgp4PMxxbpBxZjf+XR/s1q25CUuywk/1fDcZmIDnmnzaGxSoAu20aucuiDXI
Shr9uJYhM5Bi3R2zkbvPKvPgnZHFPJqJxyQBbXw3Q7O72tZWaBxkPWdK4cP4e2jX
I4G4wXdy/QvGwtMXevJIaXjh1IA6XqUpuS9Sq6kGOJKidBWetL9QC5YSmZPbgVeF
VI0zoycuUdlonvab8gCNpNd3hoerEF8f7Dm4itosWgMWKQ+HWccscan6uWrr0xlN
sU1KhP3ioHYt7bESLFW9c/0rR8R7obf4rKU6shMSBmh+W6GEjfAbSJsx+vQ491Up
3bkLKROws22aCUVvTHRf5fANUmVNA1wDjaNMnk1h0eGx1AGLarJ+5Hh4pk0QVUaG
/H4MjjdIyPnXHhSDIDWGcku2Znu8m1Tg5QXMrhJ63jWe5qAI48SJTu363PZFiLhK
APXQWu5GQgqC/VplCg4SsCVijc6nlu2fjmbXMxag+UtM4i2upjelaNcHRwVKlQPL
GIxZP9fyoTiQ08DNdt1mpcTvtHVzE18uy1Ubc8bNhTtCv7uqlosb9wS4p0mPkEgQ
DrxuS1R2KyA7w4oCm7jLsG7R2QxU/YJN3qed3QhrPdzucK6TYDDGd2PIVPQMq7T6
ETF5MZeqH7C/QhAUwBG62XJHAyyN4r4SW4h09QlgB66A4GO0mhqFHJ/5E8HQVLrz
7opP+XAPFZu1iXCIsXBm4hOHthhlvHrEeStFF06KK0G9VcI1g+zJ+/TqdIIUztvd
4f4ImZKX5gWexB8y68DmhBFBvceUGDq0QE3E+jugPP0kzjXXIOmL/5k3AUTy4Vvu
L/i87yJHuwT1yevBvuZL1nQUn4Z6FDB0gycT+N5zymdXKcTFvrSshMnZ2nDSQaG7
RQvlcjvnQHafFM5kYOSDpUOxgIO+5GFrxJAcIyFuNOTODOF0HVtjHWS3upS2nS0o
bUyTdrYDEGXU/LEQBj9W+FwR/FYj3rYOYKbEMrtEZeSpq4ZiKiix0ZM2F84FNA2I
snjnHVqJRueFX9eGdhD++KC0Sy94HjEHZ0GJFxAYlsKvHyMEVfvZ6Yjx4pzXUMbv
MiWxb8ZGUkro+IlerX0SVuQJju1iq4d71fqj0Lfj3/935FvtWhOb+r1Lsp6EfAKy
46Kxv+rBsh6jiUnWvZ6ioJA6ceOFIL3g+A+ytUEPUOgMcZlmqGyD9/8cqHBetCUH
av87/WYpWJh5ZELR5bNmnWeNPShjsdqdUJ9rZUCZp29WMjOtlx6VrcpxBwsPguwI
0e1FwieMCMAqFxt2qCH++B1er9ked1OHOZE1K6stom2RlFaLcPl4EmBwuVHKp/8J
AYeJ4YPSO31X/To2nLlILpOM4T1eVMVzxjmhqzzbAe6vFY6M+9r/PFbStec1ZavG
3y05HhQxfbFueyOVGlRiEXXAIrAcskhZS+dBLVxJPesc+GdKKO9mM+/zmI4xrmK2
MFusZyhrrdL7RpivngB1L2e22z1fi32lLzES1p2VdBUWCV0RnTlkwqio4D363BKn
xI7zgr1sh526xI+VbhuXLHKpJMMoDZi9hOktImmomfHs5Z6zrCe7SwIVKTyjDh1D
37Zhu1eUCh3HnfsnrY2VBJIQDIYt0z0H1YbvvPvWvpCRSj+asy1kslxOowbeZLUK
xybYCJ5gmvabcC5Ahqguaw4mGIPtViXZzOPv6DUZg6MDReTj1qsIfyQU1ZnnLgal
Pt7NaGE87QkvroeFzGiCpY4ey1re8mHYS6rKsn9NYp7cDKmiixrsdaKsBibo9rgV
8CQmUd9C7jS7eGN965AvmnRtmN8vWxhP119wdBqYtU0zbN90NPjkys3eHCC3g3Re
6/b81ab3wHj9Thm1yoMh8cStVk8kg7d7UGtoPed73Pb+cA7dQPEdDLdzttlaNnTf
`protect END_PROTECTED
