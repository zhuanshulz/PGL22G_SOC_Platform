`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I15VK+JBZ6PmBKTo8j/Urmfc/JmaUQxGKqUFaAiyMFH8Zxj6+mQx6mAzXWCfB3Sr
OGv9godMM4riRRrv281DZxm3oFZYHPcQQA1GZiQuT3E8Bqy13Z8JMsh+F37M5EKo
bPYQwXmj9kVyAmjAYsXacj4fZuYn0xqT8UxiN2YqJAlp/ZPns33AOD1VXH+WYoe6
+o8HUUU6NhM0M4R4dlKazvSRzNxgbTXobNvsTTH+dAE2U2lwiThLCRVQf0M49fku
bRLGlcCAq/BEhZvvsB+pS5+d8ROxxoyHK7AFhKu+qNwBfd+0KGEtrOyE0AsP6kDB
8DxiQmKODkQpMYCOOWxgLVCm622rVF6tBzgUaXMOrfCDr7WHv91t2VygqfBm0zUD
jn7Po5pZdWLHhANsKp/hBKK9iPMcUEaoH5VwNRIgJVnX6dwxR1X02xWEwdsaeZAa
0xBvqlOUM0ktS0ADqZIqm6vAaLXCZdaZr+a6EnsAa+fnFwWNv8kq+eUnbMop3PaL
QXaLZi4v4vqSIQ1nJZMyiQ==
`protect END_PROTECTED
