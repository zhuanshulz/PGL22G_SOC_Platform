`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dYIX6mMStLEi9qxR2ICzEPW1zDzWEhzacDbNd0iENs7PeSvZCc8XH66nx+ij2Sso
GtAFGVpmFtN/BnpUZQN9hicgotz6E3ID0zWMfFKB+AK6ESGN6iNiMAjPgsrLjoRg
RV/KCAdXrxRF1njJmRFDr6xm66itVV5LZtOdPLmpO7x8UQGIIlbe/xxsB6jaurc2
KmV+pOkqnY0kzSFUMr3PH5ClOXv5xkl4XNj+NBkwLwJI0LBxGRlBkK7of9sgcSGC
+PjVmeWgoCkhFBu3FXMIZTtrIFb6cmnr3chko/8f38UgI4NZDOMfXTmgh1ZGKYaQ
PQMpixxmxxfnQp0M/cI48GtVys8/Q92m2D53ey5VP0npqSev2e12uuKIlDqXclyx
79bLHuK+jvTFuC04od52OWo4JD5dGl6AGFBSl+TsIXW9LC+iOHjUJGLZFuWmX///
SonKVmN6xmV+0n/uj9HE6R0QuWTzWqAZCk8rQ6lpU/xeR0IV3HIh/LDkHHzmPe6D
/wJ3rQ2Z2AxFtezCfmN3dwZSemcYtkhtbm+/Vnnszhyd6cApYQ7TIhR3s6X6S7/M
jD1n8hEJ4Gnc2BLsDB36gMHFXMTLQYPQlzK9zFShJgMTXDhpEkR5pA+ZzhEdutaw
`protect END_PROTECTED
