`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L0MoNSvHotz5/EBJYh/p1saj2dAHrb6NviAMSGE36B1dACRxZnROx7lHyYwFbQz7
Xcy4asLxejAlJzslGUf+fFwRm+W437Ckpv8zW6a0Xdr1SD1tfXU+1XyLm2I0lOIO
BnFuaFpENV3xgMzRk5fXtmBBjkKFXfprvWNWs0gR8WyMtDAJUFRjmbQM7PhWgyZQ
80E9F5DWBNaMO44QzrOZtj+/kcSPBcNHmQGzttguqM5AR1WkWFIw/WOt77knvHFH
9boZsjIIDt7+CSrMIQqPz4LxwaHrEeaZzYsU9kDn12x/kyWTFJwekn6u+fKXNMUC
1RtbgQWr+vNDEuo+c/Z6k2yc8RLkDUVzUXEuBA4bjx0h+OjgxZLt4Sc7kSbjt7K3
zdHOa26G6n8dJwWeMd4uTQ==
`protect END_PROTECTED
