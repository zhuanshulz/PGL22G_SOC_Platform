`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TkCltJ5uk1esLIfXucBJctBrCsEp2jA1hwYLFU5kH3XERD0x0b/K4XFRojSBBHhf
HzMeMm7LVfjmMALLTgTBV04ZXbKI9dozWKyURKIOU7IFh6X3sUbkLEPFNc5tnRdg
n3tUKYvVaQtI2UTS+Yc87ufIRLojpvnGMvv6tqOVulvLriuICUGA37pZgUlKWK8X
RDXgQfXjk8TMDjJKx/t/AqjackQ+U/2PikTMLcHj2+MO54J7mOPWwEuF6RrpjvhL
tTjsu9IVUww6h+KQyaUhCuiWbMX4cbzV8EbFfCd1cpfCiQFe4LjyNlO6vyua8CqZ
VF2zBuIpNjCX3FFzZaBn47cjAH8OrEWpoXMf8Yk+TL9YVqkwiDEjlbc32cea3hth
jCfbqedYI3F+pJCFWnsKWdPsrD2jpHgwq0k/QX94vsl4XEpdFHTaAOKOlftrdEyZ
n2fuQR3vDpkgatm40UVH3P+5rCXARezpOX76I2bdmtA=
`protect END_PROTECTED
