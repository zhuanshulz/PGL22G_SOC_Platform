`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nV6Xn76jhq8Yb5zNJkAAzYsnOYWeND7l8EbhyL7RirASY1zVd5Qyx6jImQBg98Wb
2wyik0ySRvvrwXLdhQagjm2mJKnGGisjnYC1kaKaysAghrrPu3dAtFPPT1b5sMBM
lh/WTJvVIJ8uL0kZ+zLpzyviAZWMy+ZtaVckaDJIrx4r/WHpytDo/U7WFNdVyrFv
wZKcM/l11EYfVmBKmCV/86Ip7C9WJT/5mYuZOXG+YLa20XLgIVFgSVlfW0xu2ZMF
HuLNBlVV0BKHna/lUoWIvUXle7BqHP7Mh4iLYRHYS492PeNp4CqkhkO+28mAATec
i0Kjb9D+qgS4ihuuQyL28Y8wjU/mzVpIIuxz7bXOdrH1561fUc8AY6Zjvp+Ieh/d
y8wBkyr21ZpnRsQF2iyZl5psy8v8TYdRYKDJQu93vf1jFuDpvVpX31OHcWESjziU
j5OLXTh+EKTKQoUc2W2rUyuRk/wadIlRHKc8w0ezSP4z4/3iJm15A6Vu0VHBl2XQ
41mFWG1p04COT3WNe09uDg==
`protect END_PROTECTED
