`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K/EjlqVDkZQVayfaIXEudwEfwDO4cqBH9YSupU5NryLrG+yRpHtuhG1eUQFKqNln
Z02SKa6XDfNG114FmDLEJ8ipzTgxmdvgFJzuk8pTcSbWrcXaXBrXxuqaTg5STl9P
bdO4qxkQm7RfGITLpSek5TeleWu8AW6PU0LTv0yc2WRyoRmS6W1eNWGhh1uGqKQV
0mEMhke8Vr76BokTW5GYmhC7jNQbMwm5dNrvmCmp4GghaNj/rOYzpYZeRyT3mYgy
sFKKRYiaforRpL9UafL5j+4JpyRk9aW7gkyh9EHN66b5RG3yHIVAp448JoAzFiGQ
SYKt8Uc7IN0GWHxGPhaRP9qXLVEQhdeeRzGkAb9LCv/S8bi6QG4RSWncArw1SYuS
UAgU5WLzJOFoIc53+y/3tB0u85nIeRG4rSIpCfJo5EjPIaNU8Yqa2Y/vX4/+N/5g
kVAqnNey6qaZ8rxea9c63me7p2/9AuQV+1BIDigZY4v6L+voiCUbt7sBDmEdV8wf
kxd27xIpggmg+Q/iq4pLumHA2e016IakKGhK0Thceqng/b4I/nvo8tk1YEMKuHhh
88ktKbJCxeGIIR9b+aVkNXe/RIFht+EqqYSuHB7Fws1xOtSUExuwe8eTQZb3TuYW
7xCcTl5+1qfA46YVhajZN2hAtQJ+hiGyS98ugTMj7ewD0mLW+e9HB5L9GM4zuJz0
vkVw6uBl33tiYrxxrO8un6ieYGkAZWR86s8nHVrvxW4Y/fNNmJjAgId//dcNrRQx
`protect END_PROTECTED
