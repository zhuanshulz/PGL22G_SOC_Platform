`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FPnN2FR7HHNEgtz41t1Ks9F0GN5giqcHGnvcuYkJMpvGInMU0LFXKgkcvjuamaLT
zLgEAwhcMJQrvE4R+4zYPL0GxnjPupbJCIzUSE1i58veV6rwRQLIbLxJ3hDww3vO
yzeiNqsgpCId1ZLrUrLtj6JEvPFL7tO/S1WYvNln3lPtDNGAENup2lQI4Lp7g2wF
bLJulk9t7S19fIBCtTqMKA0/az1IHo6qXUYuUpZ5d+SA0X1R8Cbwg+aG/YjllGms
Uq9VsilrOozAeC9ZLo2fCN9umj2LQBCLHQOW7AhIqJYlnC/Y0VyUL7KZtoJ/4I57
eztUUmXorvPWod60yG/TXNNVVxzYNIFvDhwWgi0qOdO+MBeJ8qVyzWS3ELpK0bjb
8RusSYj2M6CfpznlvDxTzJKO8cGFZSpfUbG3TqBmbSQViiNWwoxsn4VjlSdYLrd1
wYVsh4kNY03AN7Eimr8X/Cflw9r2gndCAx8eZ4zUv2Hxj9JUoTJggyzDUV09Dn23
HsBwt4VQKaolfvMQVYZ7rKX/Gytj33S/rkIkS4NghCSWUE5Hf3ij01BpHfev43+d
e472jcswUAc+hWfjc9Gbagn09i87Uu5vPM0Gjbc4ZpE8HZkqNVoUsxkQh+9PZiWg
1Rl/MeEcVTb2ZNbazAw1psIVsJ+nfS9AUw4t0jonxzNGp34Vfsz+TlnVCE47vNLt
BMKvlxNVQu3EcNW65WICikRC64hwKtnv7nxgSw/g0cawCzXQwkCGq1XSSXxtKGP7
XmZuGG7efWYvln+dhQ6FuznF1L4jB+fRn/e8l3D9gPS203oFY2YqElAQOvAYVlev
DQdtTuaXnqfK/numTE3eCjWVC0UvbBtRCQ7YvAlEpCknP7Meshr4m3RIJI+cKyef
NrUneKG2aqaplUxbbT983SJ7KI5z3/pomX40rKbw5aetGeEiOMPImX6V9lG7s2p+
ltyG1w7KZ9FMAHrR3ZV9j2TKI9i+hJ/8K5efJWghAHeiF3wMJLh3HX8x9BlCXlg+
Ufv0qnnEPPhLRPBgGr4ZeAOf1OSdT8IhwNspS99AP/c2A3kmOsMYgr5QRcTspNBV
k5vsm4C3lcOR48DS2vnkGrvStwWTYafqk27oXtx8w7xkONbvhiqWihvNoQyrslsS
IRyzjj6otfnsxxF4VLkmmb19115Q+yTfgPwCanYH0eScBnWjQq0rilRS5iGZIWYj
mauWFsQYezj2IkElI/2Xo0K+sxYdoVJFqr8bPK9PDPX9xI4SstFE0dv27av8IcBb
MADuEC70cHUspmJ1ZEjWQaipwc4Pkc+J02G/bT3lCiKOvltC+60cFJcHtSeerzl9
KNhwnv/2xRZE5vgWOGgbNuXfSWeqg6V+7+/smO7MjtjOUWoETej4YlGAS1fj2Q9m
WUJYuSBkUFlXMjpvmCznkt38F20+vY2deVxuppEY4ZECvQC/OBzytWxJGYgOtbPq
KUAVO6MyxcTBWcnHiDFyqfCTUrOycE6ynT1jS2AU6mjazySgGug61dv6FoVm/9z+
i3xKw4aEoZVy4cS0DQdMC5W6wkx0S0te9Oczj9s2XMImHlo6L2qhaY+n1sBchAMO
96bz8vFjaDOhFOm5ytp8ACBgV8bY/YU7lut6ICNd1pqhtBxoo4eI0MyoyoWEvzQf
fQ3DN9jcq/WeUJ0LuEBpFutcV3o3YG2zJwIgu6P2VsuJQKP7XlanJkdPAng6sRZ8
OnZbA/apg4ssZpfdno1ouk3LAVS8Y2QLPL29IN9l5B8wWCqEzJt1l027C6eSnsIe
Q68yYmFQmS9/XyM6i8h6hYyUpuCjoF5ZKRb4eJ94tz5MUNYpuDxjew/U36R603BV
H8VO/5oc4Z5U/soZsG2jUhNs4087VcqOwEOwMOyth1I8yAqe4JJ/X8+WS66auxhM
AxJt5CKEMqYPRb+/2wI18p+btThb6fJ38x/bOMftZK6Avdok4FHe01CxxRiDurSO
5ijX0ayTsb9maMl6YjmmT+b+vfjtTDe2QWDwLDuzTrYyR62mTU1d8h8zxEfXHGpq
9ZFOJumNERp5UYvRt0DVkyjODWmmfaXwuySk86rX9qurGUMVQRHeErTIJVOoz8KF
+/c5XZ78RHOO4Wlnbugbpg==
`protect END_PROTECTED
