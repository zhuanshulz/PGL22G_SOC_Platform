`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5ayT/y2QuhD+aU156uVC6BN6wwYR7Jlv8btcrk00wm0osm1Uv+U+3edeaPEo7hKR
/GYQgElBlcQqPx174e7ZqsSBFiLFSGjO0RXR+6JjyHyY5rhv4aU+hxzEkSBeIt0E
16E9BXH1+mGdJLpFxm9b8NCvAi5O0cxf9O6GzKXyApzNXVoKWA3K9xZy29+MRoQG
FK0F6DQrtJIVt3nwjIzbCIbOXW7zY9pwne00n7xCrmJv/kLYDsNOkwBNZygTVvx7
ePq2c5f/vkJprecYCdkRYO04cT+NxuM+w5c3JFw/UFs8pDLrl+OhgKmX0bfhaiOC
B18eKMhh0aUrLojqY0PtZVX4b6+CYoF+i9DENSXii3Mf5sBR4dttMfCJp2dXeHQQ
Mi+TBT7Frr8bS8aAHCfDWpWIVa7LgDz/DcERSXMHCW2ePW9Al77aQwzQC0J4andK
mPoGcxBS9pjhus+Mv5WlsLBz5bmddL3wb56soL96+j/N7aOBMECSCricVPCx0CVR
yWIRwdPTnnXk7cF5qWwwwcgZ/ZsnYYaUqVB2Bd2rYGLeF6nnIQxjC3uVTRgcZUxP
9SVt+mj80yIgh1A5bMPZcoKlDgRhSIkbPAcTYbggCjKnJqA1iH1EJ/thPHW1q1tl
O819nCpht45FYm9IzC39L1iR+kfh8gbv5P3mvIDQG3yIpf6wlROzCjfnwAvaFqMB
oHgbO0gygbqAH7k0EsA3By4Edo1AN2fCEHbEGCekWJVhWBd6cSpQ8HVgWOp7glzH
UV2WHp8XsF9fYDHlNbLK7KWAUg2reDp/yZMzaW7yiDIDRAwHs/sbSXsDWlx0ok1+
O+P3L2y19be9sq5J7RR5W+Hmnhk7J0FFnxRxfNScUiegzU4cz4W/Q7/Z1nPESRQy
mw3vRayx5Vch1/MMpRDHiekk3ZhXTYqJJY7dTGxogvMq1X08xByo15TbwjO5VNyO
lozfNj3oH5BNYNg4TUJBMk5U19009HQ2wzo0iMdUx5mSjzeMRIusmREt1Rm5lqkO
ENMj93DjorkcAAYrakk8lg46hRQY5OGnhVZ3r+83bUWttS2hl+CpwWJWaCCVTGUm
9aZmvwOboxebcDbiep4ct7FBiJi1sBWX8ob/AE07Ir2B/dq3LdKH5wRpCElqMm66
EDJP55q0xygqJHIrfvqAOV+PEJ0hKWJN0Rq4N86A9fB/FpjNqXdlNTrccpSGM55f
Wpw6p9+HRdRxA10ZOXi4rt0q2qIqhpKSufe7WT6E/+MiyG6muK5YpRyBt/APSw/o
BEL5RPPWN8kbbW+UoEFL9T9Sj5hx7HsvVcIjvboFa0IOS0s9ILFazwS1NaqY+fJE
BQ1eA8rnGfNwo4WM7YDYAfUaTw+y+YuM//hVkSVu9KguwwtW0tpM5KS075aQ9eL4
OIk/q5AANrEtFEIM9Q91kkGDMPtRPhvb1XFixdmoa8QdWTJgIHiKkN333wleoReI
//1oom5qZNF8+SlaC5QZ61fjcTFsochCThuJtF/WYMyrxvfiXP2cbMcULnMUip2W
bm2jq6g4CNawmIa4U7V79zyfY2pLOH4kz88PK1/EtyCM7PG8IjDZEQlNx4df7oHh
3ONGBwuIVijv0t6Kvz8i6qk34NjvORpQAdBSwSruW7mmd3UiI8HZ4PTjUP2XAIKE
hLCC4+vJXs8QTm2mcMgxmORjJUmPuEQyVNZNTKAdI2QaCNIYRXtgrGPXhsOAzThj
Tl6USMqC5RhGPHrMAD47Nu4WJardmh5kHJDPS8qGSr6OR3FdXk7llPwj3SFeVdgy
5mmQodaxKDBQu3OKY458O6Ao0kXb2yIuuEQ3STlkyZk5xd8v9fnyD+DdBYqeL7UW
zj0CzNHi2AZzf4ZaWKl1OK2TSp0Nmg4MyNjsf3fG9n2VpUq/MB8M+M5CqfakCqY8
AaOgarY8KxufgnenaFzP399wlWivUGh4MQtxh4Z9QxT/NMFJht7KITB77TASocwN
F5UgZU96HnieGw+QupAT3dk8YbwRf3e/ANXJ1V+wyVdgYfchASyRLKr8a29kYQ31
91PBDss12KulBgPPpbmb9th0aQ2FgDEIcXQnio6ifcxu6KVrR2tgaecX7dKbjnKS
OAHn5RD7hwpGVJswLYmNKHXqswt947nWzglhlimwPmBvQx6rJSZ8aKP2qrd9l2rP
LKBSdQNiT/5ez6ZstZbJspOOJc1yRwYthWpzIwS5xqodQXRLLOXKvnsKzG5QpJJ7
lc6OdUJDXcNjgKTmqAJTY2zr63sVIc0H1tY1NB6lrkleyl7EflPqmC2n7ajRpx7n
nscxaiVy+CcCBvxLKX4XUJEw7Vl/kPM03jVd+KyVIIDhFNUs4bnnC2Oa1hYWm/O7
0wCjvDlW5Jnjtu/kI9Cp1CQopbt1Cj5wFGDHE0p8DaWLjcPRJcJkalg4lbNAs/pg
EuCQvt+63RxJgtR6Palsv5ZndDeiQCr15mvxvDv1/64IBkuhTtgeLTn5BesbdSjL
eSUU5g5Q6F4kKwk2Mm1+1xYmFOhoEescup2iKRqKghy0F3ltxXK75izLhjLN/IQs
V0RTN9pa0U5T6znTEL+YPA+DIiraes6i6IjUArBUY67SPqUJu2JCFWakrwdceq8o
FvAXJdRkbkB+s7YDa0XR5UQ9JNH7UfMA4d/40scnUVtV7QwYp4BkdODsd8t//EUF
4fHsc3rmuzcS+5EJirA+nZYIsS6tjyFGe3wH4HJo9Q2fVb6laytYD7TPpoYNq2uD
pV2ehot0U/vuPTy3kelkKitSxjVX78hR8t/INT5/2cHgfB9sJFzYh5AtaZtbd77J
Ex+v1l/DDZLZ4BeJBvj2R4/QfMA/DsLBobG+4NwRPTiv80H8d95neXUSrd5V5kNS
5VG7X9ARcp6QXqT1RNrtvQ==
`protect END_PROTECTED
