`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZQT2rZz31jDQCYLXk9vH/2Zxz2wUQfrq/0iA/+eYUv6ug3Ua6QGYqtOoBgl8qQKX
A0uU3/kWT/Oc+Ba+nraclwF0h7+VZRxgoZcY/2f+2o97CFEsNEQ1xL7aspAukUF+
9hjLoNTJXFqZ/ltdDDimdnNvZyZwFktH/5ZtjlH1p2+j+1PtGpXvn3oANaIz7Pb6
oFacNE70jQn908r4XJEcO1VATHyJW/qJjMyca5Of8Qc3zpuZ4omaWDgNGNJLH6En
qWQN7jPTbRnVwr84nEVJ1k1+H+E/gIBQLcjmOotHTT6QrWpZSw4jYQp/cBpONYiT
iMwZh5nLZQgXCQGInKByrCK1pREb2mu5iahsyhAd6WLmulQ4EcmF2OgPxc/C+ngg
FRev8AJ+Rpg5TJh+Q05Acq9VvOhUiCtqkQHSUaIVuSqUv2vgUPu+Ga+cFBGOlGjE
2GwtO8llUS/6xdZN+eGF+BPgtbjuiFjh941bKaeVeKmRo7vh8fkHPtNle9owoDFS
EC+p7tJjOKGrEGjD68CPGUoacPe+SyCnUVjuOOpnRefg6KlDTXNkxPQ0aeb+KYqf
B+dxIT0rB1eCVAP9Dxv66I0J7RBOqT/uMyTV+GfpSDB3CdycfmsbEjpHpbu5QEEV
9I3Q4aZ0D4vxDKCIfJek/1XsKHSrs7gDqQzKwcfykDnEhlP5dwyacwilBmG5sSz/
deLpziRYhiF0jUzR5T/2YCnOdLm9CDXIrj3qmSOhR6Loe9MCQfQ+0jA8cZAXcoaL
F0y2VRcVU4kvWc601K42/HpGeowElyDJLJ6cOiX+K7aXWew0OAgeAveXEkkjk+eN
ACGYm6ItVGX4RDMA8A3PFaVrzTpc+dlNTGmuwtqzwfJeCVRyjhVyxYL6Xfyr1New
bNa52Gk4DvadKpIzxcaNLP6k33yhLk+yj1fbC/7yCV0UMHahj46PD58HOxpr1z14
Ga7OX09f6NloifeYDybUPwG1Grl5dyc+3gs5pE+qoejvurLf5keTfuANHL8egbPg
JUY+jHWJ2nzDMN4mNPcsE7ZSbf7b1j2hTgd0x8P68l/SKnrxEitEzzDY9MBVbgiV
oL5YOk+daw3YT5RBDcE9t7o571RjPHdZOyotf6lrCIk2qL8vc08hizZQLYD9QWFo
wYYUZJ/RpNEz8TLtFSSYsLOw7ojiTLy0zHSnF9hSDaG5YZBlWz2NuEjerLDC3B0r
VS3iHiiXEI21w8rZq61nOFY7pwrlgJneLLOBGZnv3rVZMDv5CcCst5Hk4Zo8EpZN
VazM1xjgPlYsGnCENzCNt3ZV1WBv18hIRVs6JRcpplVfVUoZuzLbx4LSXA5kU2l8
NB5PsaCu1FtTRtRJ14BhwCTyaQE5qUsP9U9/WVr7UC+l7b59plJD6NrDUFqWV8as
/bKfDTlEZgqCGJNPOqBDDC/VgSYrnwx+BqQx4q3EwxVeHfxzRE7EhI+EYw2Kah21
w7N+SJdLPsIMPA1TTS4+odKCYWAnWHMYi8WKF2bwsm5d4p+sgFtFN6BwBvss89Sk
CxdBxSBOpVL49sGYTv7H0H0PoqjddysCD6QsdZpzt/Df2z1BxVQx0nm5cMyYlswt
wQtcIXiKAUBX/ta7J8YwyLsyoalZSFUGazAkiEYDhQpD5WYiO3IAx0ilDpf2U+fU
DDzIo5TFODQ2/Ooxbz8l47NsctG/pEEnvrCfS+pztHne7vNxlfe/XfI33//TSDVb
NgUtkaehFq2rx9pfw/TJ7vh0OjybkNuARQYOkFQtF6qVxPeWixp1RXkarQ606NWq
I8Fxj35DXgz8Z1MaiqiBRKUVO4kVdtMbjLlo/Q4GrkBKGEyyBU7tzYPwdMbXTci0
EWazmehrQ9gqma4hqIQuBs0wuHB6+B0AJMsH+Gw00+viIc25gxwEsEN2F7nqlTID
LIBw5DedXlU0tWgtrNf6jj/vVLBwuzDUvmhtSN5P3lhLtg44Ih2O0RE/EDePqgmU
epFFwh2t+NeV3kgEYBISxzLalIXGXuCvvivp3UaNmcdZP36/aYkw5/3hGqSVElD6
cCkM/oesAu6E3Dd7oPWeuoEvNoiVVboSk3Vkli8MWcIB16IhzGJP/D2i12wFTRk7
gWgsdNL5bnazQ/BDjda5+7PBWUFrj7UZSYCezGYMPKMiqyLNyrcAVni3l+/lZ96G
D6OF62M21IhSLI44Vbp4P+2q3Ox194boT1ZJXdOKhpx8sgB54aZDrbnd2Y33Tiut
5QTUXUkHDj8SKlD0EYNple9tgdVzixIN1OpYmKQ+HFBkdcDs/WzED8J8wT82kL2+
vX2Wr1mfzEHyH2WRHaysGVM+GqtbSihCRsqx+Cgd4z//9sPu0ZlM7iyAC9BsOzf6
DdTsm3mokGD3g4tqhHrL6oPXFAeVYikl/YhOOIKuLgHvZP+AZUj6S1co80rQwepg
Gl32Vy1R9YHmUtO4zsbKHIMi8gDf6W1hQG0niqcjLLEs6tIMUZVYJT1pLwYQBf0B
URDJ8zGtVFitiOaSaBDEwjRA17jYeTxh/l/m++pDKwgCVGaEXmajUilx1DadGRxS
yYANcpAMEkc+bCLF5l1Op41ppWD5Nb4dx6IMQRX4aYXVxNjunqePR7cv9UKmO6LX
P0SlZqNQ7tu5A9QVtDb4hNlFah6SaGPnJaze8L9cQMkRjnOT7+S4sNWQPRAlGeWm
f5UHBci71xm/zf3ld3JorhVFYXgUx/RAaaUILjXspj42twDQgt1AdBHOQFrL4rja
JAX3zvUjbEtW6kDb+Bc74DS/qEP5C8U8UFUybspUC910SyYbxS9N6LUzeR/8tF54
Ge9aRqm6QTQApBLlBI/AucA/tdb1aIzXuKQWveYPR0PsIIr1LM71poTDN9VAZeoH
gKMkZhN/RI2neii+pzXwYs1rYFUWQoFB5tQ1Pv0odNwhWVldZorbGO7ISobYqvQK
1/xTnXtlM298SfiYr4wQFLnRq9ZunLnX0TMfNHuL2RcAn30nJeTYfTip0+8oRKPq
elWsVbMKfg3/EIXZDtP0W2yW8qPkCmM5LZuK/mqj+dhA0WwPzbVX/r/WMurN4tya
P3/1uMXPlDDMe1jpDYhoUtSfJVE/VODZNQwha7s5edpDm7ANAs488VN+5LqdPvmh
fPzvY3too4QiCsZHlTjpEubdyTDWs4mbOn8DPE5LzDYBuOTISeafBjRqDICanLeC
RzPlcWSdaZUBB3y8JMKSBLY+nncN9EoIPyaD+TX5C7aO4xJAXk+PUyAU9mWWNPFt
rEXqBNBxEDNG7d1sAjs/meG73hIfhVzymyOsfO+RzZuAYUQwieD1N3dag9IhptrV
T12Cb/RLAolBal7M5xRork+o1v+7JB6tRvvvhlzfi4MUoG3iprrsXOomVGh0Y9T5
p64jT5RkK/cVZbdyao66yFBkomxxQOcj2DSvMna8WGMJVVSJ98lz2CkzGgwAoyyH
FocnfaTifh2GYLVO1WINBtKyJutJHzB38Cc4ZMRv5rimqVZ9u5SnHxXZerF3HGFZ
wBJdz8g83Dtr7pSYPPjznMNmdilEd2BCvX1Vlczih5UEPbgTxVvFAKeoPGqHamrJ
4HHOXXuZ+zT1SLV9eLxyK1cz6p8jcKhel2Nq3/oM8cUKW9x4n0g0hIUkujxh2jZ3
Yt681jkx03p8Pm8kyzb2FSmD4Kyz1YC+D6OmBuzQ8iX1lpkio5aXM7NWrRyM0EAc
MogOA/e3gy+it8HHb2B+yplQ4RUu98s9kEoD8alGKhSwJFzF2Z41aanPfWOYJLBc
bQEkLJac7hpyHb+mv9yYh+Iyab3Jbb8/GYzrtI5M+z4k6zHYfAN3WKElb2xhyW9X
emMGn2/6AsjRww2eE0/E+BaxSONGiHUw6OdGWG7OrzEYepfpm2jKRefgKI6FMIe+
DT6sADOiUKidv5exdlGU6FpL06JdICwkz94yxS5X03Hj5jSmT2BjnPV9aaLNYrKj
2lU0XwC4fBg6STrnftCkw1tKe8aWT9BGOTLDh6qczo1MpkfufI7Lv1nKkdBstO4K
ds6ZEURzAXSpkkUPNsI8pvlcwyJcFwwka9eT9hKcMiw4xJRD5VTbBEMNVgTsM+X2
Jyy+MKPVQR8bzeu9MVl9QLx6kcciVO38n8nU/CQiq3rYfjj8PYu+licBoBtTMrnE
9rJcbv2mzJeNnyjFHPW3PeZEd9qwigfxsfr2U0T8dzC0e1duCBosXP7bR/rcAipJ
GLRJtU2VJIS71YBBNim0IJf1yBg1dhc+2QC5zFCjNm1l+cpBd7OTYdwjoHsEuplJ
71ufY7bf0JCVnKhRNajzOKJyBtKpIHFNxl0CEUEY4hWeXKgihuRq1MY70UV8x58G
cVonz+b70Z/1hscN3zyIgB9oQQsz6NazUKkcteK4s4eFhcO5G5LgXWye0TVpW9Y+
`protect END_PROTECTED
