`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VEMZXPPMQSGYNX12FOO5yKcMVfsJipg+gVYqZm03b5ja9pa01xLPdVslzcw25kzt
j57BbvvnquubJa9KbPe2cy18CfNpSlsH+QZviHacyHM/yp6vtth58cxpGnNNFVI4
zcO7t8OICMiwBtNihamRL4ER4qR5EKkdpiwQYaQdtzbYAVGMo32wV+DN7TaUGaiu
I4wRvfOS4F0F+IYyZ63OAVMEZh1ospmz9Ae5fb/olMq5hiV6Iy4kjOb/JXfGka1I
gNt4L1awES840xk6wkAOBpVmMaOpW6wxzZYWJ8KqDFhJN6+OnyCTp5y9iDySZqKj
mJ0XnbnAngx2Mjykc/81vmJ4VNNh0z71DuMSmvb8QVU9yATl9OJI4bfmPA4SYgLd
2XVF55uGRp4KQ5va+xn1cCg7N3dpn7BTb76Z+NCZztLuH+KsgYVCRw+CWWW1nO83
SZfumGSLkLqIFgCrgo/vnF3AmutrdPG2VeYVEETOsiUwadBMtjvY17lfVq7jmof8
oJkwUtw3WmgfUejiIEp/7fCwq/GUa4ROc5z/7C9fzyYu8wxzZekwGN39MI4M400O
u6FIhATMWJYkKAuG2lthRzMBSGcWbGRLes33HbX0QL2DHUM9Act+H+2BAS9oBpay
cdw6eaqfZ2xkiHWbTetXldfnrFCIQ15dGCKS+i7z3F8i4sfdfE+gJMj1e0c+BgWl
N3ronqeFAHu59NaubW5goK5kf++wFEO+91XzCwdXyU37KooxtCx8H1fvYoSUua3d
HfmFf8CHHAZxwQL/ltF/hBrvtipHggyvcFMYpD6k0B2zFxwmdFlsmNF42Evxb4MF
hcVc2RbKeANlCMYhh5VsyQPH1gD3666kTJkYwzpcU6m4gQY9rQoKMAxtouvCz8zz
bJUH2tXhAwth0LJPsxB5t+u6EFKiAr/04dRKgcovD1UFYKMJkT1QGsGxJNUON2IA
P2cy5nU+x9LDOWzrquXbfq/wvm2B2ztVwJ7d7dp61GKOZbvF9K2LH7Bbit2ipJVF
AbDAGPrAfA/wRGiZ8A/qO3b+M3mOf8Hr11HAMH+fFTAAppKHB3o4SsUhjwoOBZGz
UzRTzuIesIjgoCfclXDovOSsZVFm5baFJQj5NLsbIIa3+fD0tHJeVOuufc0NPLm1
SRjV/McxTbLOv1mt1mBgfylt4ljeNhIhqXW/05MZwTPBfG6z2BjdkvDtxnZ1JnI8
lYzm5TYlOV6Hf6RcfwGYfNQYAssgQZrSNeuj1QqEj6T/AWyDuO8FY6TsujdaT+Sq
IUWDmacI+K2D/qMdpvTjWu0J6qf1sBdIhMq5Tjs6lgrz9yNlf3B3zj1JxT46/mSY
xyp9POzvAAOYCrT6ScuZlW2+zMoKa6dRK/IK+2PY/sj+ThNso0YxjkWUZaz8gQqC
R4zfV9wV3JesjB/FADUfehm2a0Di3jymya2qS0II+JFsgEU/wKvvhZPPzkGFmz9f
5e++hfngCNqkuGal/+WnQP7MfYvgbN75pzpvQKNbNwCzNOBUIkCbglnsi1esTCcI
OLU18biUyReExmimO1QBcm0jdyZR2+m3wfbN3HmbfWeU5j+szvF4J6/7tuodKxG+
P0siUK0LaCMPxio/ShnyqpfZlmS8RYr1shSb87F9iax0V0vwqewwL7YcmzilfnOa
zsCKEXAdetYaA8RUrq+K+q6ahXFSrsbbbBbLjObun6NZIaec7UwjLSThE/eRwOSu
NITfgP3ZN/eGTSC3HqdJXem0VZdIHR5U4oHTr4+AiPxBiSaySmZg7t+lHE2j/fYL
73YyYGI4Z8qUTjkhX/+44rcGWyM7/Ew6QjQTIPb0r3kA9ZjfLRZNL+1OQk/jOr4f
K/J3Xn+UZe6YILFKOp+6vhvNMeKNzvBkPKjmhpyg7rZod6QpAwbBXJBWi/cL8d8Z
EFJHr6Mv2sXKOsnc1cYg6IYeCtr8BNkNUs0b5vIltFTDR+WW0PP1fAhI5Yp7pR80
//7rjRpSwgOWDNYfdh2EaX5ctZNBs3jHy3oUL+DW1SiotJCar8rrGzsQFMHKnW/j
6mfEkxP0DI1MtJfP5bwSaCR16fG/DDyaTO5P1rtwFquQ6wn8bRURXjkRZpkLC6DN
FoCtH4egDwixx5m2xcKZ5DaCvvCB0apXXJ2UZfZhuT1Z7nMAxqM27fzpuQ/XStsq
ndDvsS6zcWLuDz+dSwx5Cl+b8xb7xA6aO7vkU6HPr3s0mGvrG+x24+kALhV2JweI
rO2HsjBHCETy/IAjoCshBOOX04CoUex4osrsTvbYjnmEtCCLEjZOdOre7YVIrbbd
GGhfjcxgO/D20GOzhqgiiTizY8e77lzrL6qy5wwp4H1PMKBDH+8tVTCevtqrAtnX
2HKPqyC2MiBX9F0sPmnXKCORGXb7KwiQHv8NKqTYLmR7SXxsIJl4VbvI0LarV1rO
817bwVAjfAG3Hk/gFDFKhHTJaPTpvzYpA2zmPoFeKTZsRbnAAkIYXIICzDy5YEis
Lo0f6Ec2RA6hsTS79/NPddrMXfJ4/eGv0okUvUSQBakKZN/YNjvLchfT13f8edkB
sN+vhIJsRJyZ2j7JRjLc5+496qlzalpnQEA78y5YpV6mW9Tze3sGkRLWYVN/K6+v
40kUlhLg5yNZnAlC2JcAbiUGQKxSJZHacRZTkFeXNYoWtQADRhROoCVyFunb7Ba1
yLanQ95k60T5DUcfMe4kxVb8fcezbT1ZLGXroogtkVfBA69V2q5k4Y6F7Mik7mgq
ortSU+eBRAMmHNm5djHBe7baX+QZefq5v/rBLZ1FcGvpYazLzd5IBQ00R+lh53+H
QvjbGBVaZym9KvkNrj8lFTfXF0ocb8vjewQy6x+qdG43Ju9jfQtpwZ/AGbuKEGKi
8IdWmOSWUtyVCNzg9ZMBFuDaJ3vmegwXDKIAU/9MzGv/Ie+3w3YvdIYvWRA1Yx5H
gnLFZ6/1SXgeHz/oU7uc95Zoetd4RSWhGftfd5U9iVYp3qwMbo08yyd1+EncO3N1
jccuriPbj+Aiug84XFPCnWPm3mmi3PM0E7zeUi1JmaH8j0LZponOlyqCWuc8FV3g
olh99u+Nmu6SStclTcBB6i8y0HEQHGaxt7/vME+c7cgwRqNkc6zY9/NcDy2p1k3+
iKmWJNhdCkz+HI3E8JCai1qvQhH9qM/qGIUoPtMvJJy1fcRICFiaKm2bEaopG/mZ
`protect END_PROTECTED
