`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d5LWAXHVtGpqoE9fvzaYw5qEaxf+rDEdxeTlNcWHJMTBP29iNMZcahqb5/7+UNtC
4oSxoKNYezNVsg37Du4uatSY0Qxx0KREIjk316lPChxARGZcpBgcnP1uBHxEiLxL
+j18EyDw22uJBfuxMWveD1M8VqV3NZZHLyy3gUpb8UongqwSw2/Q7oFGUgsbHLuW
Mj3SeJtuvErZ0yEwgmDxGwQoQVDdu1olOWhA2cm94kDbOckxAyl3HNSD2OkntrSi
Zscr1SpVieXZfucBT7srSYTSz3cBjCckIYFNYRJU2kCAlE/9pCwE0jioIK81rhE4
WAaixIh6eFYo8u17lPJJjh7orAIR87uHqDsfWYJUdLwrk0tG2HWSzdKv83NtCxiJ
kA8gRcDQSwSzkDa6aTm4gRYRFRXII0fCWYVRN1UhUf/1uwm0xBfSTDZTdVTBcEDA
xApMnMvAlyji/KSgYMjqMmBsRNz6n6NNIAyC+okd0UKG0MGTjEKEGKsXrIP0injx
Oye05OeZzm/vhr9LuLsfhg==
`protect END_PROTECTED
