`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gpSRFWuXzmLQyB+XbwWFPufVfdYt7a/GKA9L3hxd52H6YvFtD4G/KwOyYzWFi64k
ZT3stHrtq8j+jSXPCSO30SxHbcA32fHyvd1xgYc/VKd/FDL9CrxptoOs9SCMfN3S
Z+9bp9S+REU6kaQJG+UdXUrsi7Ps3PkxQ++X3AI1eZxzn4otd3OcTxypFAx68UJ2
aNSz1RjryEC4beJj4tdkSvpUtP5nUdVn6LGobv9xQhT521fQc7/35q/Ec0VPBvtB
TnE2wJ8EfcE3MFt62rCrn6/2MexhuFyJFIued42TuJ1QG8daLqzy2p/q5F43/Hnt
+LHEO05fFKz3L0VBTWLGVHu1uXdkDEabEpUv5YaGtZLHHnhVVm/Bri8KwPPXQKzN
gZm2GBN+HLZe+pQzmDvZMrLga/AlSt2zTakWv/ptPmR17uZXS+ISXBjHHetKUO+T
9poZDCDFcsKjdtKb3O55hisVLRgW3ET+MWfcppr8itzO5AMyhY3Fv23dO7KnMEfr
s+7/FTHUIG0P7UlteLWpLDkx2Nm5sHlURTAM8HT+7I8Q5BQvjxm/p1xiaBfKUj4Q
j4m6jsMpANjnPqbPEYxaOK2+g+q/SI/c4bymAo9zMFrYG7BVnxzM5D6KZSupIOvj
KtMEC94C/GSUMl/BltefasZxx7wEBf6thDKJpWOy00OexmZy0Q9Qid71yEDH2/V1
72IJ0iVfNZjMiAhsueDIwqSqo6nHrsqVNSOB6ub024VNozx5+Fe3wpGjT7+zkDyM
dId6CzknmqkzFUoNRkPFFfHk+/I57I46a2kieHsM3xOwovR/lqHF9Vl1unnF30xM
U+p8zRVdKTHhA5zYojL3I3KNbAftcwykjXuM2cnrwxdAGSzOdYddlFp4/v9H2HpO
ZkQB285aP2BjXHWIxq7V2KcqZDxH3Pr+ooborKQMldjzjCfqiq6ZPZ9nEQ+P0i3k
MYFVRfIQkKSVDQRGNXL2adCvmgW1kJOlZ5EB4Vl2a5P9VLfprAI6+TgAhdVjEM9o
/yelmreRjHBgbiyq7NcJ0of04sbWTfRQNJqe4Rp1ahQfeH9EbNN7sk2Scvajv5Hv
JAZOFUy9pRUa+D6/FWSZLg==
`protect END_PROTECTED
