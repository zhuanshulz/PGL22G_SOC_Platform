`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4SFEupksxuQap0O206Mhc7hG97pYoW0TO6xphjEgNW5N1jtTpEnFMyalLTBzSK/x
QBAHWoKPBiSSQp7PL4YLzyvAw/EhP0MsH+/1bx2dYUdjc+50pO4wSMxw37ZiI3R2
NjBGoUDUOw3vxdW/lcq3573iWC9Ei5BOfUPCbLprvnNns3g0e37Op5Njb6mLnNfl
B567CF1M1Clp5Ryi4+fDRloACoAR8YAfKl7ut+hzEm6Ia8Pmsjraj7FZYydy6uEl
8L5tzSAcrVBgrIkCBkywq9l/HLc8le00gsMNaD1zpvwb5vgkN+PQnccHmABGx1Ql
kMkVuFQ18s8M60K2NLBVtcUojUjIfP0MwjV1SPJ3cwnx8dgp8dfbEvBoKaq20i6p
qlVM3pgWLEV9HFYd4npy/tScK/MBvKPBK+Baz7pBA2MyNb5PnbsjycPJQ0JWzCa5
ciSiIGRxWXJsVGKbJ4/fFbafia/swaI1+8nqWEBAV2zCi3trfhZMylrVbyJfuBou
CfIHT1HUrCbiPQrz49C1CWs7LGZ/rHSQshyDE4azrXSvpSavhHxk4MfyPq53MW+u
Y279TANwtFKHfsSGqD0XAmSnwLBYZoyKSgT7B6V6a+urqamhlOjJGBnDVpGkE373
CdB/TdVB6GlaLvcw+r57053GMiUW7P9kgEHqQJeNLnrO77GEU1OSvXeitmkxMwjx
grAEjNV2LNY1/eIjQ7sw8vE+CS3PLbZWUSwO1UXqeMNT1fFLtky8aZpV5XYhgA+Y
UCIUjVl8Kwfx6ztOIiS52z5R/VZr1M9wTQluJlO4yeq5aWv9Ixolf7ERnv12V9wW
QIRaLX+r3XfRLHTJLRcdSYivi87CiePv5wtuLzf9oQc=
`protect END_PROTECTED
