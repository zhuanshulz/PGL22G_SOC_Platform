`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ljCHMnOQIt57IQ39Bjv61Psn+/Mgsj8fmSKTIxdo6QD91zxBhI6AvMtrkBVPAhDo
w3PZIsbtco4jSDNxE6jFYc9cDbkwxjJm1am8K7kEuNJkRUyTzrYeniL0siiEYbHE
ev/SIuTKox97elQNeSJta/X+iIigkLya3EEGDV2+AyJ6dS+bKiTb8quYQzbyzPHQ
A+MZhHOGZtpAOcDgnMmGq2r88dlVgWdzKO4sVkMcRolzqVc7LOp+Y79YABrlflPj
UfHlAk8z+h58h32ZyZuNsX0LauhnVkfCvnlGyalCLNK6pccL7BaqdcS2bW2CgDUf
5uI8NUdAi/YsbM1cFxtVNm43XpDflOf4ugtx2yWopWsia1jaCYlDZKq0J8COcRC8
uZG3i6TzWa9QOh3WcLCFSesmS4s7ECVd2x3WCZx2UerFZNN28bzrfFtTq6kvmQNx
sDlkIzbYUmLzK3rweGsTBCa1hREifLHyxr8gnBSoXYLGV2zRRl5A732ZWb+7P3MP
Ep6Sje/uQjbf6k6bO8Key/UZF6vOAnegLey0HfTCv/dQW9uzm+SJamyBGlGK1aF2
ijN1GbhlTcXPuaKK5iGJtTl//uG0WYiqOBCR8lwDdeWqzzIzoCIM7p0oLqcF8cR7
EOBe//o5PFIooAZnSQHh/jrNo4uFYn5DT2ENJkQfDNKhDGaKnhfOqGWP95pnwMRb
Qw7t15ZMirFM02M+k0953259bKIKhJjtt6gzX8/b2064yKhGR8KzlE/MtmS7XNz8
ZRDstR6QqelCCch5qMgF4QvhlX8hqJ+ZisH3WEfGpi2rwoujz7Oy1OxOyAEA8uJN
1BvwAmCguHV72aRMcyzg2GBWZr+mCAyKnJQ0NSu/3Wy0H3lE/ImyCWPxQpZxwxZP
54wL6Lzs3cT+4JSoi9vxUZ4xJXwfvlnFH/yjnAyAV7ckgAazaQPD1PSDtQyq2Mpx
foJ3LgrGbxcsvxVFVF84FhlpfsN0IYNUMai+tTzY9SSGKmHEfG4J1c2zpn/gz4t9
+bIUVC0TX+3PjtIXrApwEEBMn5gahIjp4VqQUQAobNeP4xMB4HDdh+1lPMfgDHC9
te9iyynhHTnwio4kKqk0aoo5x2DcyzrDq/kSZBMN6k1/afZwADGr4vlNmahmfA34
uZara1fpNaSzclfUR1MFayoLHvPh71Ny4JdLbUwpugpcn537u/NH/CG3p2Nn6If5
y2tFR83EMKFKigkeTfCKiQP0AY0Qzafcustg7ROQFsF7gM/DEtdKiWoqKIOHyaKk
t5O3OtDWSJ4Thu/aA2yqZqlrXlyaI3FqHnxuX/Znc1/UndJgO7K5Sb0UjI4xwJHr
a0hXn1mPYH86LZOgu7r36pM5mzqQSCKfXi9DqakiHLrmgr6bU07RwtE9trxuYuFF
p6GTXv+HyK83YQ8zBERkNJJxnBM6y8OSoDiUWdgZmMrAmGvE4iQFcjxU0sfkccpT
6Z5TqMU9kJmAOMYGU0PYrH24oVTmFa7x1RQFD7ThC9UbU8HfjdQcFTwvMOP4c4s0
oM6EF1OBkfCa2hhs9Pr0ngrW3Sun5qFZRSYEQnq2k9DIWo0R0ISdbqETd7umP/dD
GMzmjfGxfJr5RXST+APgZxt2aZTQRoYv37C4fIbUb13bnVMUPi0zqSp2Gvpg6e8s
krSKJ6DNxiUFpD8zntUHbfRfaRtWCY4O3jMQP6K10D9aUPiisfhmgLR3RAWhYBm8
f3zAXy5G7HaxCxj+VV/zrSUX9R9qS83q24MUVXkwqgTAtfwXTPYwxX64CD5LLJ6Z
CQ4fSllLX0KlUXVWBQlhk/SpymO/lQrG5tA2CvsjNNDvG48/FMitPuy7pKpg9Aq0
Cg7wt/ZnMkb1nC1oZISH8UMdMaZLp2qGdcEQLnxFrHWuP112hTyhMy9dXG3LG245
X05kC64eemNGmx7Izc2WVb+WIrJAJapoeEKhj5D2pXO8WCB2P1v19K/OVQ13Ufh1
PQoEB2PEMmrx6FUUMMQkwFGBvDD1zG/4Vg2MS+JM3Cnq5jw4CoY5v3WgBMaLkEk3
2UhCx6Oij3Z/7rfSJu6suofdk7xSlnOpNW7V/vz+1DNVCknxk2xJ9XmJLbNfIUvW
5F7p8S1msIGovzEqsdREort14pnHBQEQEPGk91d+soR9Ugj0/EX9Pb0t9gYDGT8S
vHCUgb5amuNGVNGT3UBegia5TTTq8lPAMMKEphiXKeSMZDxQP1/PaqUwjocTrBL6
dibyqoSeA/sPFt58N1LSgc1qADpdZjwlqXmJI7Te9KB3cQdKXMTNUa/R0az2aJ8k
zw9oHRHy5lbEpTXJ9gVNTU34fOC8xiB12lkjsXk0uXO9MlnfPNnxaSRpkGcKlRTX
mmeBL3ehAcc4/D1Jz5i3Q/VEHFsugYlRrhHZA3DS5grHmYQF+7NfUGvrJe31q8f/
6cCsSxf6MmRxSOKhcBVhHzNV5GA7GbD9zu0r+1PbNddSv89CEd2esd3/nM93X6V3
tgrinkGhpwLY+sw1G9V6I/jIMaZhg9rlQzuMrNBFAOIaONbAW1yyQDTAMsvIgDHB
CNSMdFX3FbetxOmkriuPvePWcxGLqS/8OUQm+3Ed2UoWkRUdJxtrb43Z4J7m3rBH
2C1sON9A1ZO0QdgxpXe6DMf/TZMoxnux3mLhk5yMpIbdbz6yxhzJJgrPMBmmzysr
Pq7g/eTx85X8fJQA/a6AKGmvxlyUEjFg6h/0BcAwnjjWVyQWuAZrlz47+PUNzHE/
mN+uRG3qn3/bko23N4vgbTjZwvBPji1D43T9Anoo/jUGQq3KTsSYktoGmTxXQ4dV
uR20+OhxKbTYjepfASQEbqqnnEmF6vqkKOSG+brX87+srjHRFcNi/visPjS+OW2r
bS3Zwgezi/zptRLar+U02Uw5bjRqjREdHWFKCFhcbqxymg3XTfVSgCUDal9l36W+
x3FcWR+SCbV+EpSsuK2W+7ckYSavHtYR2gb9xOVOqtAFx4A4wwn9G7Bt8HhYo7PM
QIOyHiRBowOjz7kr6BXHESB+7dNZk4kqpxfl0ilOCbZHaw/L07K8xZ9u3xQvq//p
8swK5sJmhiVd19LNv330pTrfW/jmsw+wYZ9td9o56F4oiavSsnEV3dRu/EMNhTWg
Vuj58T6g9zDE0uSoN23stDMFIw17LlvVpo9oWBRcY7TfhvmAaaupIMmBBj/mbbyo
bwOwwAvNaVptvRugg+CBXVJ+9JY/iDgGCYnwV+EUIVuCG3qtgfC6ZxcxdydHXbNc
XH1mfyX3j/1vaiMFQCtWO2QhYwToVQTtnuKjRB4CWm3QBtM4bwoEx5tbUjxR5EHu
5WNDj2hOStAdDtmKwscKiKbQ9Scx+330CvjbciWax7Yxsb/E0ENaRXbIAGBwwXv2
6AeZDT9N1vR9uDNLtZuyYff9Ia3vQ8ys3xeIgJXTJbQAQDLqGzhfw8VUWSGXI4Lo
PLbTPIeRCFLJIf9dDApazVZoG/sGQJuK+bIWCBy8bGoIzNP3gS0HQ8oytZcGKd69
pjbyMWPTPw/7QSZ42yc3cOVGQomLZWRiRLRxxJRTMYznZmtHOVuy04w1GMzgP5rm
DBFSLurqXaZYvjji9IO4upWbVWIvu8NEkxEF5GxeqX0dlSXbGKjpoTxUp3Eq78bC
JoeqqMq6W3KLRU1I6vUKqZk7zbuUenLYHum8JqjeF8LVESGElQ7TkgrE3B39cg8Y
fbABuYe0lZEFa3mWmN1mCli+gu7XXUjP98aI0NENILdq/3njfS2UC+xW1RaREBmi
eSKc7q20tJC+lqvKXEq+zHlMfcN/DIbc+eXujB6clQsiBGL9m1hAv9vkoENbpWQX
p/SUO8xg8W7x+iFbDJV/uICfvtbr3KVI6S+an5AEP/+2N6LqOYv89uNSNp87+6oc
HF/aYiIn85FfRUvdxforLq2rAxuJ39q4ixk1QQh9XEuji2HAk0sJaEbmjSzeK33m
0vDIAujsUf9g1ul7mIfYKblET7rnM3XKoaUAGl1ms3rrD4XL2vvjbmvrGqSFpWxZ
iRKY7fBxUkrX7jWxGip+cHJ1vp0tS41Fi756S/0kzT+OXA1lo7zQ2HTrfxKT+Dbr
9c4l3tw63eB+0lDeQ73d5qZNxwzdTrHB1ev2sn3BI7Ll30me2fXd8JRLYfnCrTOn
s4bCRS0LJgv+V37GbYwcLME9ZlZPUzsyrZf3It4uAtS1kR/QxLl15KZCshZBgEPm
uyWPH79Go7c8Lb+APbMFJ8qfA8KLSq66OXxyDfOC0ApbKEWg/kW7fsRot2QZ4oBb
umoUSK8vA4hpu/vjeVEGFV0fnFeYImRNCYeHNaTmcJhUbeeA2UnANC0ZN2Nm3YQK
RoaYQF1DKmcy604UTho6LhGg7YwCJnsRWUvvUvxO11ZBo78pMnLP38myXV64x5D9
A1AgOOhYMrTdtAtHeGJaOTPbLT2ABLRPVB6vSPfYbd1GxNbm4nbHcbEFrok1k9E6
tE40CobXxW58Z8nmQ+L88lIESs6d6HvtThxAvRrzCWmfBoT3bmDsc9kNB0EOgPMs
ET3fcxZSiDD3EmlTUaezbnl79LvNgVQpnoctzxPtQV2aEvgx/sYGI3aIaUL3eELW
ho88xBa+eUYIa9J/ukC1tzn8SSx8o5DxjEJ8jllBCji/UgBs38MrsMTOdoM7w0n3
+7CzK7f5sJQe98pawAMEe9GxZI3lEH1/yGqDMP5DyvAUqnY9Ao6lpRHDRn0qArC/
N3RjMAExkImpwmgBBh+r83Krgc5o0C9ufp4C8UtAiQ8LrEiSwITNL+0ky8cBwTgd
SnSvJmwCFTVUJ47HoyBMWJ1Xo7pvG+XhAwG0lHmbr7RcmEK6/ZH59LzOx26/VcQ4
cRoZGeu55OAQ9UbH9jD8W5mHAPE+2T59CI4rAuR1Y3VLJ98N7ia/Orh/uorlCDO/
ZNuEKFH5z6h8wsHJQTIEoulZI3L2gSec3CcSHE6DEWZmLT84jGQgdzh9iFhrky33
cbUFhnRzs5bowdEcINYMOakGKsNcW1Us8dISUm77HaslbOhtxA43EJjhFusw+i6Y
E2HKXbwa8ftYXSEtQi8t7QzvjS35+ETA/5QZ/piNi+F/V8PWWoAdrAhUM7LtglqW
bc3EHv5dCyQM7lF+P93G6vIJsGnVFNbTKGuDMpFcaTbEeapXsMUvnDAgB6DX9SN+
g3uDnhKNkY0IKIpw5twlntXaRtVh5Rd0wpPviZ8V5OvpWBRlujIAxPRlzERXB2W8
aIfyp9KfXGgdaxcLhNe+QS2kDawgOj+Kkd6T3ZkoHkd6ULL8Mwb2wKGQNRlYhbhH
TNtQGorANJGuAgCoQ9vJx3ZM69w+Z99FXrxrvTNceSHBWiRiFbtOzdk2jfF6Ji3j
YNMOK+XGDe4xHIfuMONM6p/wdIaH1BIX7NnbMVkmZJEJnsH0C7CDJE4zMD/Jq/Ty
`protect END_PROTECTED
