`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oSDo1agUrGtcpAPpWP4c3nAUeagBqXOWXOM3Q126CokrMFYSlsfHRVLEmzpTax5e
BaUw1GENs0qsrw5HRPficuL0lccxEu+F+BOQW9+hTXonNpEO7e8Ka0YaYiGfnvln
QorV0TEm0Z8u/bScbAm2eQ25uIyNDyPwvpLjFctBiD1JBN/fLqg5PFGKBxpDQpA5
fOfimpYbfM/EZ7j7FcWN0zqk4TIJgB9k1dRZiTHfKoSQiVsswxgBoUmmg/UeMq5V
Ma8NZrEi5AUcwWVKika3KtwfO7xp1rDzdvOCYEhFfysEQJJClGpdG8EfDx9Wb4Wc
WA/elKTw0d3wZ1wDQdHbhgcAs3ZNoSUFI/RTnBzdQkzWM4fNoiL4uxzpffFdGpXy
vFv8om0Gr0W1FsJrGwDeM5SaVn/zhnOK/Z8b16NBrF1uU3gfhwtxzmT4mm6SmZEc
XeYSTNvZ+nEDhWIGGZ5jh9XzMzjwDShQJ4AfWWlUZuDXbUAgEpXfAmrOvLP/2Lg2
DCG+2MsSdmvOtuF+xoBUxntyI0nI4lHalkRQVkL3bZVtkmOnt7IpY8Puwx6/kkyP
ji3pHbQTu+Kj4Cg5wFcKn4lotj9XbZcHenxbcjERiwGWGNDN/q9AwwiLamefHBEp
6ExBah+gaWHZxATZEcgcRMAZ6/MYtIlpVJda8sU05kct5pB1hws3JvDc93cLOLrH
gjcK83dKWk/F5vHUhikIUdbGVqe7qCVuNd2U93NAKGWRjs7LnsKjooRODdiGYnYL
tUuK3KFZlWTXS0audmkj1u8hEOGwZz8OUQNxP9bViwGUFvbD9iav41ExAkYT+yXX
flIXGCGNKtJ1zFMW7OVS027yDqgBahQDaUN9BwIbIa3AArIu/jDHXL8m/e4tj/Cq
gCoikUd39N6Prm/PzY30DW+KPRY1dWarGSs9iwpC6FlDTnKvyMKt76G/zO3tjCqH
QdOIMsd9eyF3IT76cCewoQPkcCyIhy++q3jZI0GITXeX6ZJWQiXepmXovd8vOcN2
WY+8vH8EEWpjqBkcHVV07ioK2PMr/+ZmN1g5aUwBbEE+BJzxPQ0/8aJk1UIBoBov
a1CCZbuSkucUxTh1lNgcN4cf90L/GdK9g+JW+CpZk5pHmsSjrRxNxImQiIjbld4/
R8DUmzGwCLTyen3eCfyK9r1Y0Qo1OQiwFnr2sdvUCNFfU/l/uEWn/hMZ9xC6TKqP
qjmC7IjJMrYIQz1bvXI/QWIE+vAkDajx3jpEFeNVzc1vY7ax5cphtCageB8znTt8
K47G8YZ9NcrQJqE1gcZjMtrVczyER3CFaVbMBSgJCHBMewXQ6a9+k4bo+XGjA3aA
OlibV8PEyN6jrGOIu3tBRPbDTW85VF7LK0RJONTMVKIm58LWvsIf9fxoq+f82miV
9hS3FFLKP5orVthafFJBVcJfKUCD9D72GQL8DKcUXOvcvqCBPbDJ9Aw9yaR8RiM5
XpN/pT1WIijZkrocOZWJ8tnRqTp6Go61Dp9aQuF1HlkZ9HaaAsKQ9NTXMH5Elp0n
8bbsJ2F1sxH06e1q+MXHJyQXa/8y7NMNgDdVX+pAXR8fgY1KwqATBh4cLThhv+ir
gvVDgvvLlYMgw6IQvNL0HsyLo504C2bWTQOp3GVqpvY072fAbQwgIfmXNNmqQN+c
2/y/tuMXnITSbdmjdnxeNa8aLz3gdiNWWiKl9/bLbCVR5Qkq7JNTdzmgdss0Ym8K
7upAewi0GJPfImW63rZDf0gX1ueiHF4tA42hsYrwzFPqSEovMw1EL0wTRrT2qqhf
bdzpovvLmOUItEGDhCfJwP6+Euc38Rx3IJErnzKcbppr70Q31bBEBFc1JVcsNZcN
p54OK426d9b90C/bxN3hHfySG9BebAFXhYtYNjL5jTo30NidTp50H6f6kxegT/ss
Qj3gsAcPZ8iF6hkQOAKZQOGiCzhqLgAOlz+GFHpNw4nHus3nCh/BuaIOAf7NqvO6
nkF47z5JocF74R8n/E0ucRe/PT438oYVd7RFsolosaoyiitwEVcbKLcE1EXPzM5q
bYsfD3vQ94sBcLPsVA7VXQzrwPeWNedJHHdqS9wIKh+Jhks82MB+hDChOU0/4A6f
FyAePRCvFVz1VNL8KQGlzs4lrGl+LmsJ2S67G97Qf88Ay8Qq5+Z7KQmgm90Z545q
nsjOv8Oj+tMWR2qW9ICNGkHMViSQlAMLzADCduNLO1wcHdYzNomfENQSUru0+zyJ
bJG+pSU2OAPrCPiKZ8OZmptLBj0aUwORXBxgQ9QTtmWnPHoIDlTIa58s3gVbQJDQ
0L+sLfKzS9kBpUynHbd+rjqvRl6RbnFRu6qNMAHKR6pZJk8CKD0VIWFYU3B4ljGl
uIHA8I5cGRu6/qIh77XTXI0+vXqlo3v9YqoHkMhoagjY1DS/X+9SCzHqN3Biof7a
/yxDPuVfQclhdnknlcFrGmAkrNrG6ZShbYKHVGKJ9XkjvoF6qMuRPfPO0oK/pUru
nbqcIxBllAB2eiPI6lptUqEd2WO2zF1ZERFX3JEl2nXTcjTeKReW74+Ocw5/Uqfa
i+FtsIRQUtklhPOFuSIefjkGdZTDuNV+EkDl2lZy2F3zhyauLuN/aJvDSzbHrHZ+
3+VF9ssNp4Z+WtEC6UmYYRQqJz5lxbBYiWgPIzm+jdjjgrOoOBOEiFI3NRmkKTTn
oDy5pNs2fDSw5RALHiDvjhK6ZXVlivSUkRAuL30k6rT711CzrTW7JfEcY93JCViR
fbGyV1qHrdc/T03S2J4TKF1ENwPxzfnw8inxQjNkDFfpbEQTwu7iig0NnyUqOp0s
1gn6kx6Su1XVB+Prq6Eqq868XJKq844Fd4Cug41TwCBbKQS01tHK2fzRqO3Ul6gk
IPyPmIxVcK6H/ePZGgXpKU2oJx0tEYYwVZsdzNPuQqztOrSXrXDkQYaTeJlqrfFr
gfa61yFW900l8DCUlREf1RxoSg7N2IbTlVFXDNBTxD33xwpFNmUC0RKQeINnj91x
8uOUm2FoKHYcogcCh1fVopzOY3w2uKPRH3iqi0daRhrpMJyyEAiRVokxQC0wEacj
MQ3Jto6tAQVHogdWniqjzU7GVYGt3wzsMYt/202i9f5Z+CVK7M6a28IyZ6xZiGd/
J2SbtNonLBpdFQLNgn3LbkLMuTzDJmMeby/ycYH0z+suK6QygfnQapxwa2RylOHQ
J0rMPS23Tmyrmlp9+A2r1z5v99uE8oV1mII88bwPGr6zAMo8c2qzqNsVk+X2Y7xt
xO4LO90QmJyPMSEdOqO6R/cyf1yQ2UUiVaK9lmyznw4IY1+WVOMGujspGgjra1T5
uq6ATH5Ew1R+irvC6rFobY+mfeyZXP2UiMffQYy5AWwf5T3gvSw8fWHn7mcUL9ex
7S2g7tFXT+ez6DWXeRli/DAKHlB/bAZXeVtF7kjxIeWIuLuL+M6nI6e3VEEDUs6n
tjvFp74AcbetA8K3mj8ytJL1OYhdnV4mTjf/CX6mObNSKSRzqjvCKVzBM9IIvVWO
kVtEOm7k+tY/v5cxvdujsNVNzbgxu+YBlc4kljS2q4HeuMCCU72S/on0ru2Oen8I
f5UV27E49kfwd00Gnakl1a9ZPNP9K5FlStMKzc6gbtkL8zSivmewCGZ6bMt2KXQe
yZDXezaZG75qAIoJUVppqlNg4gycBZlCmHvQ4AFkk1WPGXxXSTh+itysMvIjKLON
IVTqAO9v4u4RTLQ4UPoogmmJ0OieaENiJGdltgL3KudNeF4YNxsnMlRWg1sUa8ue
WFccHkP6Qkt2WKQIkN+QLeMY9h5zHe3h/J+cp6jUty2Ck4FBz+TlBh4cqt/+bqfD
o7/onA4TaZ4HMVo11+dBo1PY2vq2/YdnBiIMTbHE/1jgrFw5y8qV4xupEG93cvB+
xtzhz1u6db5W52mH9+3cC5CQsXbL60RMwgkLgcaHoTBAFjRzXj46VN+1Tc0ff6WD
2R/7lCjbWah1t5GGiBVK5zkETmyPltgR1tyB2MHxZIkfqf/wIKpn9bq7nBx9+JIR
KdR3nrLksRmiCOYryrYoEyhDPICTBHPVwIUFm73V1wuopzS0lWSVJzw7blDaBI/5
Hk2VTnVzawRh0XFUdlqm+9R5L6uFv4WnQLfaN5i1qr3h6ecpcuYmLQ3jQOi+w1ut
ztN/v2btQuJ0PApN8mp6SfEcEaOX5MnbWzBBbT4eG0Aqw/WwmjlLgkSXlElJEfbe
4snBrDFqTGFqImfrrJ24eYmASv0kpvrDjWKale0Djl/3BmVkgaPaEx1VCFDwewrC
N9QlLxsYnX5hpziuPUhKtyY7cbC0nmqZ3gkyHaasmtYwHSFDeTwHXph+Oytq/xlK
4cwNJPlWvEALZKjymahx8neumlqY4gotQb56x3U0ahLn9DBKWrD7zXA4ELNrd8qC
Uk2oVBP/YP3xkyKyG3wLeC5MsF3tbYrqGWbf3Oe1WnHYBiBaLP4wSAu9VFrK+GGF
gt7jzwJBTpG+ugppQ1ruQvLGY995LSzVXWnjyeRERdBNWVSmsIeMAMVh+U5/EK8f
b8FW6mkEPpZBmTuGc/kWCaOXiBKbGh5a5oP3C6LWgGakyTqemn3igLWI4H6jtVf1
t2+mjR9fYWfj4YTgEalskYtwDIsTre3JUwbvUXj7gp9Ls6ja7+wHKEwfoVQEWxG/
do6/79IhpmHhpPYFpCJ5QxD7UBTqQ/pLlSxbmXIEYBRMFBYbjG6kd61q8fSbzHEk
RZyiunk/B7R9FPkjUsa6XUe38J0OqUXkV9w9BAxN7uM00zDlbTVSE7S7P+gDemcK
pSWLCP/7x3gXiw82xwz326umXp/s+PX4x/J1DiN0nZqFMSkXPBfUvQLmwtb2VGh8
ZiqQ71niMzTJAfx/gVhXXYueJFoJBhi1TyjLNAV2BE+VzCGV9NtaN3Z4hSul/cAh
FQgfnltdaW2E/rLcy183shEz73XQU1krcjQw1bHhnDMbRvY1ycML/enLhwushxMQ
y68onVILc9I5/Hl6BEwNlr0LZIw4Y0LICS0yVPliY28G7WgSK7tGDny5GRwsq55Z
WNuCzj/VYgYLsCJoAXF0AAFP+YELTuNnibmvwHNgZvsv2M5RXF97PrWOUyWelkHF
Rey9Rf1XwjVJjVQiImS4TlK+QsXOj4iM7E+HRzUizzVp0KlAWFXI6qK3lbvRLCEX
Cpb9GaYScX0r2RHpMUtWP+nNQRl1/yLSYInzILVMkpIZU1sKTgxNxQN+3Ng1WNxW
ilTc4F7lsLZkI38ezp8qE25ZCdghV5Y3rzw9e/EjgoWl32odp4ACoyRr+A3y9QIG
ibqn3lRkJFMYpgR6H2gZpBEsHM1MTr5jgDjTUBaQiOfHRqmDxMjP/4j/FaLswJIv
l4MVuMxHf6X4z2MH2Zlqh63b4Uz+R0QlKV9r1KYOSHwZRb9ZdwEdqyYNjcQX6EbM
PMdo3nle5QUqhqA+7124o+eX5e3PsjnjA0nj2/29ZMEOqfbj8ubYeQ115MIGgIOT
JS9dhR+kVuEXl0oHtgkkTtIN9CO+myJ35RjXVIxKsDJRHXZp/2GLhr/T8B1Y7lSC
G6IAHg1f/MNDagcT7RWeygUeYEtM+RYwP/D+77oQ8xPaPgzdlEGizjMROiv1hAWz
SjpLS5PiqjmAoe2WpNLfqRTV4ZX8nL8/zvBrG7vbkGIiDGRCijCzuMraZJTGny2Z
hgzRS2tk4ODO41+EWqMixg==
`protect END_PROTECTED
