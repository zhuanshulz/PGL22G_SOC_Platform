`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d6IPAaVZtyJFlhfT0ly6KW8Yr0Ue9T3iTpGwEBfaxgL5/B7qkKp+1AzXlB4MCNcM
U3OymDU/ovUuR8neQxFgpy9QfIWBovX0aYj0iqsOcO+lQCANmpqO5mPcjT+FCKu6
byfYjR2JO3T9F3MqrbWYtv+JYDlkeOeT93SGAjcBWx9ZhtKArVrtKYJt+gYPovEd
Qb/tqtsHNlBxqBOyx2YDDezAYpIs7CP/uhKB7kG1b7iYhP9MpasvlHWZu5/H+tDa
uEcVK2NL7cM43kTW/udC+cW/eyu2k8mtOmc2a+H6HmZZPL5O0wCBSe0KvU2nDZAA
t5vVcWR+38qTbIr+PJ6DVdOORs6Ty2ljiknQrvqiz1MDU8JfD1+pdzSY547rkLbf
xzIIRg2TIJuYJuqt4CXy6Gy8dOlg/m1fNkkEmBdiu0yZ/tXJuvhjZvNLa72lR56l
2FxnZkqrFbA3Twj31T4q8KIUDD0MqwemABcYUA7Xl1fIy3qa1Boy5RsJ0yJkHj3r
HZ/RpDuK2/DjWpm574+LCAiT90L/x8L8mbASJtBEnft0tl+kgdp/RtZlbJKX+53h
tLwp2ufdp+AAMvc5gdqUXofHEqbL6TPf3VEcdyF7HGTmOeA1Nxi56+LuTpPRvQZv
IijRfT5mTbSecNqk9zWZRWOs4+N9QuKrstSBeh63lD8/pbunTn7SC9yJobyK1jxa
sO2cj+Tkv8rJ1/Jzwu6Mrsq/PX65pinxsiy6+d5ysW0JApevuaN8Kgr9DG4VRL/u
xOgGwQs78QoTKurn+qzyyCVfHZbIkv0VpYklAu1QCz9YkCnUzYobkGXSdNSNKK0a
6WKruXuBwZIyVzbvock/hqXT5fPjL0Xl+bzr2zCdZw3eM3WAkK9sNTnQH7g73lz2
7/5iOdRj25EU523TZIoC7H2sNsPnw5wuzjV48YDIG6/fEeO4JpDUGu1Ih0Tl+1cs
7mOKkPhq9gzSgj2n9nZXdrh0YpIoZQtcXsqbmRvlhRJ9X5bBlxKknPBLuOGYntLk
nsJGUGKaAI2TwJn+/jl4jfYkFRb39Ts6N6Ahk33TsPHZXP4e7epVNDUiEcAyz/Qj
9wU2OaN26jRx/PpMJRkfjILMNlbMQp9PMAesQf/kJ2WknelMdRf5Pc68jNle8W2i
GjMydj7ev+pMrKxCgPZO+7I3FlKEDPE6pn9D9WV6ZYOGwMsJTcAAHkBu6NEG5HMw
rsBhFyRY4zfOKygmuWxb9BVb1FQVg1rce9bJMK+IE0C4jNSoKUzZDo2Fq5e4+TJ8
nylk6h9Tse30DMvKKeYZfIkhQwerIvMbFGbUSv3P9W33oSrX5Y8uL//enifYtdCk
dcYtFLocONm1XpJRQgatUcHGOKcHRkSVk8oWOzzJeYV2L2bU6D3Uew9kHF8ywvHm
VQlatDeJWUuGyG/szR+9V12M4wRNPKOKHsNMQk3TEFp4LmVVQCNa6iutrFjxJy5+
LvCHWIeJguUxtyhGMeFLASdRCouscfZ7QW8S94thLVIalRYoLas0jY+Z6tDkRBrC
zyFGBZyPwUvLdj4je6vK1628gBfU8/NZaGoLhF9wkFHn1LCJyz4DO0K75ENBpxak
raIKBO/QgISDENbXeWod9PS5Od1OwsTo5q/UH7MjlIxHw65h7tn0po9MvaQAIwYS
q/N92By3gAyloPLdqRi9ZopCBgDVtQK6XJiT1sIQErd9YlPTELs4a1urCEk1v3MM
PkhrhRvtyDaVWz+vySLeRnIlvDtf5c0ZyyLAreIhA3IJnAv6oc70Aiq1psYF5EaI
xC9CBrAWJ+1WDeZe5yRnLPzs3niqdBdTDGyHRkFXBZYPQYYVtrMGNFJ2KRNxDIB/
m8Kd6TEpWfaiw2yQ0gMPfw0MIxuBJWGgiVch/Hxoldd0a3gp9DW1Dbmw7RluRO6J
WQDxDpDBexzdEHRSyxf2IJxR9NkfV6WxrCWOmX46BvuixnHOfaRs4gLZ2ibJj1UX
B8t2696SB1I4E387pwnqRDfQbfhfemLULgs4oC9ET5TI41zc9HkKbgqztDp8r+Iy
BFkZZ+YtKm7pRShDHD0+PMZbV5Hqp3JL2drt6TT57EeFYgDUsZH8RylLe/CSo+uh
JVMIZQ350YIk90QpbET2X7gN4+Z7irpATXe1ffRR/CAOo+3HW52VsHg43G5t3FD2
t0awt6JpadrYr1m0rSo1el+F0VyAFi3OUqIvboXj2Ni1FZYTWUNbRSBGpaCzlhGl
Z8jMkENfuRSSNtSw2CQkhSuH+IGzrS3KN0DpY355zFDIux+l4qDxHiFqQOfIQANL
oEuePSF6bnb3qutn/ceEOecycOJ7cQHAXX+QsgkIheYetK8vHYiX0oOyVjtaGpKr
1haXP24i3kKH3Kjl0JQfDX5wmarNk7vpXVOCPoAa6T7k8a9/O3dp6CJuQEyIui3i
FYgMdpQ5LQKYoQZj9sZDiwsfrW71v7UNkXLMW+wS/mm2+SuRc/7IqfThxjMlexUm
zFqtV42VSpZJQSgkkXXVPycVOtgFOkSO2yPWctwQymNChrCccsxJKat6Q4I0QUOB
yxWH/8VxvKhayxUZYg6/+8aqQrAe0WVFhXFQuCluSPLnAR20DZ4zvKdCo3/yctXY
FTHlxskPth4Xz0OFqBnzi8VDkeK5zqD5Psfc33hQuo3rOInLe2LUEiZOAELRLZcZ
ObOWT/tmWvNvfyG+rVNmYWRgLQv+sC+bhVG8Hw53eIOpj2pI5onmfWZ7ECRubOjU
/gcOOJuLjpi3qeEnhkc6MYXXK1OLF3daMWOklFwSoNnSKklUJ4rDh8Cc4RJijayB
fkVrCpxXTYVS6Gp0HpvVIuxd4BvGoc73B6V+gDnibea6f6Xxtf+mEVijug8wj+o3
aTFScqnrQXtOyw/BfI9V3pQfIbOivXgNwKUdCEBHscf2ZvtbIvCxZkY3lf4axNTP
Brfeyff8WH9h7ku41ahFuld0BNSClikTda9PSzYiSKrPYddORty8YFKnWR338eHS
h0uuI5+8ty+vmVAxxt3W4AbfyxtFDr+mdARw5K1v+biUiH/d98DkqqyhvyAgKNxI
lLSYYw/rZKi/NQPJpeefScgIw14r+o8DreAU1CEcHWHoTKGass6SXADBTNomxkYA
uvQr5jXpsvGxhtcigSAb9UnYXuksyxcPakb6jfrhm7CYeKMDIvqMBKlj3lyetsoO
smhTsY8PlLUiOu6UHd7AwQYp13a865LTthsbTq6mmyisLA/QmKEwjdnxKkY4SQQl
HQ9Jh7LvU+Y2RDKuiCk3bfeCEwJBBMgMJr+xCFQeT9z7iINu7z9juBsLUuNtLqyA
T03mdpNejostnvqQKFkqnfO/zbB8gXPk/kAfRC8UF0Pg1H6njGyw/g12FlFc9MxR
S3UbKGdbgtDA5GlM1z0WWykDilM6/7/2KeWQczsia7Uo4STypDiCpCLzCPUGNvcH
AajbKz49d3SZzSB4LOVF1OJYvaBwMMm9Xqj0ZvXb59cicYJPgtwCfAN8/qSq255u
W6+Xg0gcVWjwzB+Vml+dOmQzJ53eD8jVyUDRBUznF4Sg7eQRQP1BdguSLdH34k4F
PPWZywfnYNY2gqRPlRadQzsHF/o6NmYrznNJHQHH9ioP4Ty+SrgcQZKdFZvJEIBK
wyDYbNBK9cCE/Vf7Sv+x/Fqasm2o9BAbZW/tkQFzuCIFXDSF24SXJdjv91/R5Luj
xJkiZd+kjx9nRYEGvg8o6dSsCsRQ7WILNYFu6ToTwg/1NAa7h5sGVGePrq7JchDb
/87Z1syx6FGXEsPooJn4PFs04/exGqwl9aCkV9s+aHqsSz5dslzlkqRenBdydjT0
hlVPjBBVaqa26dGp3M/LQ9hDCQPVGoq3Cc+SV0PbL4lLvO2AXGLeYWFj8SjDNoip
QwaRJ7Q+McT7sWfGblbICLKkJQwfR4kZa8GL/GulPwuYanBWeqCq9hXMDn1KduSe
du0y/hdClJ1SqvWzot/AmvYgg3qar5gCnN0eH0/BhZsEB2KHk9OT2+YrGA33gezW
Oub36FAcWpCOaaD+R9CUxK8pDXgH75K5kbjyIJAjzkGgbvS7SIEmhLNNQDS5SdS1
C3LxH4zcmD17WaP2+M/RKiz/ogBg5YVba+ydT8zLp/jsRad6UJ0mJkMd0OBe83Yd
sLr+jvpNBSNOS3ux3OsQcRrWHRF4QF4cpEwoY2tu4anyWu8HGVUxv37SPR6MBpGz
LHgm4YNIU/dbtFEgLDqii/nbIZQh0hbB7OwJWOVIMgJSXryu5lz2gYqu856mRgd9
4ihPcWLreJEhszjJfmd3mvlfzvkx6F9wFpqrUyu5HRDOnc614tXjz9T99E36Erfg
sUL5hrLmHqqniyxzwnijnf5So75m8U2VQ9C0+g1Qf5tbSqE0J+jdLXdv3JhEOBFn
U1ySKUi/VM74WVtLWA0m8YdmwNM3hz/WSlVHo36r+9tSs8Dem2U8oFScR4yoDrkP
ik/f8OG2kiQw3G8bhku43E0S77+M3OdrGpwyUwMnX3JlyyneXnF/Jf6iwIYoN9Zv
l8XA7YVGmMXybvxGTyeum3dfFlnXwVzYlAo6InHpyj2SyexuP5yX1k3eD4wP8rC+
9KKbC676Yr164OhbjquuKe+i0/nZXFKn1lwid7hdwDdG81m3y0PfJi+M6eG9YaAd
IJ29YtYAzhxYk4/eB/oSiX+Hh+GXFp6j/HI18L4Rq9EaR2WAouLLu8u1Fj/s9Fi0
tU9rNX6a+PHoTVICCO3H9LKSwsi2hx76TLwOW9gZa1XikMCi9JOHG7c+k4ElJ9Ng
jpMXlhtuLdDxS0LPKPzAnQC9ZvgmKco/ZgtnTsa5qGHdjEI9OgaY/kVo0hEzRa+W
6a+XeGRNwF7HoDrN/JSz2GAU6xKHmRYjlEIRZ57pbLk7JxCGpWIJBXPzbM9pIirs
9eXIrqDmEz6/a639VFHi94pXk+JwsuVZo9EI1CA71SmtyLC3bTF1yGm5GD0NfweF
Rc/0ybRUwS+nFqAAFaOwcK7CTLQtj+4PjtcR49waIpuBObK8BCqxFOUFddjGGGeq
VT7xKMkaz1EL81/cpT4D6Bd+nlM+yRMUVKX6dKpzXhYqZNEJmD/+9V61GUnEM8wq
lec4hBgYUpsaEtqTeh+wQVglyUwg9lUoSuWg1SVsJMf19QP+vsUJwjMOscfM6oG2
ApighhtL20VPoUYK7iarwC3q6+21BkKcor/enYKRsZUNyEqcO4uMNaOiM7hPb0Ul
ZvFPRdzNn13rmaJTcd9RP+hAxQVOt1U+mAtuEAdfpsMwo0Hw4Kba0foAZOnWhHUj
B0zq+/KfEeMu4iz43yspVJdaWF0ZJJTp94lnvHk4vlHGhBn2hMXI1O3V1LO7Rgy8
I9ZvFAzYFs78w/aJMbZJjvJ6jzj+ScDD9Z0hJruHywUGMSn1bD4Af9jq+8Cibmbx
qjQLEw+SIpxEWdr+OM2A6n9Z5RqZlzdU8ApMi5F3F9DglNsSDy3qwYmATwSoWjnP
xvDLJQFI3FH4YtvXuIgshw0wlos2m9BCWo3BeoPAIHHMz/GaltFO+7yT8XjBzB6C
WzzDYf6EKqmkwDPoT/r+ZRbKYFX6UrrEcIjmF71MXjdHSGmnEN1it8qpTndWTYsT
KHCeymbuugUoGgd2LccNiH8GKGGTlJ900tJV5a6daXaXn2o+PU4cWaBbf8XaRdsp
VGM24cLq0+geVwWY2d+a5w8EEd/VTOK1ozxNKu1htytEGvF+5TegI3ysTSPX/D+C
c00+5jrDP9SM9BcdfNnQXozHLLvXw/8oKIY1+vRvbRRPljMmZEUjdl+bPVJIDku4
PF4M0W/sG1830KgI0RLxmUudwqdLu+xqv6IYLA4UiWJu0DrHGnHCzpz7RNRO5CqH
wNKHJ51mgZwdlKPR1XLqFBMEb+dicuqoyfnMan9w8nKuiicvm4uhoCWeFvEomgv/
1YOsi0O16HKiOzfprpZ2kQDV6RWbNZ4y35cRgoPkmivP4C2QoHgtKFaOsWTPYXJ0
9FlUcO2nY8NTfho8f/P/wimw3ClTOUsImqQRtR0ovPR7wC6y1whNhQR1akKu0amB
wjY0OkdZfuqaXZRQknywEP9CV/Yj59eWAdi5QJIxj6wPQu1A7WNHN/cPLI8U+MW3
9tMDgGt0NJ3vSVPGS1Dbvwl/W4/lamV6BgtlQMwyrfYQTR0p6nXu6zELzwBEjoIh
pK6O3W69A2jU7cewc1SRmP06i/r+YE60wr6qkLr5vRS650pDDA6HlSk5/XNcxVgY
WGTz28JzKt0fJ2Mkj6pB6LWdUeR6NjrVgtGSKHT2N4X6qMe+MLQyr03dTCgGjSjo
+AhOipc1HcrXgODt6OJg5uZbET4TfBGtuRAio1m/u0O4D+pqUddX9hgX+teR0hXC
VIMr0InTvvnLlJHr3kJ0s6PpQu02LA2BnLYgWYgeuF71ReZ2PamuG9AZrIqW1DJy
aD1ks2TCrR1v+81OqDL7tu0bUg9ctY2OBHyX7mtXf1Z5HaEcP81rl7EYeauhBjf4
eTg3GVJ/6eRxS84jScoYDJOyRLqtlYjHyMhr2T8CihSwnFqHdv+3ZWDovXFY0Wxv
na4/fAOervZ0Wc4R6UOufD/76gMix9s1VodXS7m55yjtC1NfvebGZ4jWZ++4G3zn
bHoQIX0RTBs3iwWaPlf3gJi80XG2BKV1YD8FuZq+fOtYD82NGfhlOx7CJ0UERnp7
srjvPP1/SZNn8kTXFm7lzUaP4YZwXt8DL0/CI9NDINffo+bkUFvz+Jx4f5Dy/rJG
R8uJDgju24UOTS/9jy7NCaS+QTh55RS06hZg4mHyHcoNWb4Ypk5wIUdMne1XcOlI
rbu+ic5jvC99mqlfhbpoJGvlPdAOYkbg6JfCQS7FbVOs2k4QFr+KRDackazJFRuk
9RFq6/3xjiuqGuaJmyEnUrZu1GgK64zIWqBpNxIbxT05ZuS4NVN5XT63Ue1chcv5
xcisEZsvbIRR11/O4qvWRfQj34Xf8dn9SVn6JPdufciX9/8Dw93GNmT2yCZx9aOS
uIz/uGh4MnilnrnV7cTakLan2DnBP8wB1PZETBmYpjPdmnz+VaGvbQYROPmZ67TV
/eIx7Ny0nGoJVEN4r3f7gIX8HeAbfoVzGDeJ1FQiBcdDGXC0LivcjYQJXIyuVTX2
9YR2JU+VAICLJwz0bqJxj6cdaVqhtBlJ2rodaeWDPB+cc0BuKEpiLc2tQCZ5/G+9
aRAiCuclBKISuVUzrLTdxKcn7GfmtoKw7oyk52TT+GtqBlkCDSxaKj/fjTgDQ4I2
69fgBFKIpBra599Z/eHtYz70UT3/k4goeZji1KEEyHiGTJmg53CC9so/eSI82TxD
ChtfEzKo1Tq8LyN7TWHhTlS7JMoN5ND7cEw9wnOyB6ZAJRo4bMI8QFQsLH7voqOn
AZeJjDBOQ9l4kZdlPLslFbwpph1XAflXOvGVzKNwowvNrz0TiT+/QRgefAWaNfQv
6bDlAgkW1x4RdOM9QZqm2I2z6u5yqAmG8JHJbcUd10H2udevVunZTR1x8FOmzCpk
aUQeZZCoYOXZwvh7I36WQphOx5v2OmAmhbq3UdcvyFgSZArvYAikwqZxRmvoEmMX
N5fwBqyzxMri4TbPEz7T7/q29OPirQ0s9cIC/MNeOliRNhLlXXwyH6UbbPzfmqls
VXtO9wIcRvLCA339ejmC6JAyOaI70ukYGVtb+vP4CsKuNtFz/Uqvyzid9SzRuqJk
Ea0tHfT8QTB75VyFVu7DOGaDRNXLRf9kCpciUnWtBardBy76EisepoOKnHdB9heo
dY8lfMWfJ11vFEX8sixK8g8/Le/6v5tH+JBFHytFVP6kBaEC3Oj3eFvCyoqtRsil
6bY/JH9R8/Q0QBeaRlaL6XdmsPzt9nVSo323hg/qwr8OlYFfilaoS2yIAFBQnbsQ
F7kjx7s9FXQOm4cFaxGWqPSyZC7yNofG8eN9ps1v2Nj1Rb7b57A9n26BIOmGAFo7
YH5krvnmBiI//uF1pBiGIZY5nlrIMWgseaVPk+dUOqd6+jGiuXMGpf2cvPViZZvi
s5F6UHV8TF7GfWxSVeEJ4wmDnDFmvOubmogCnZD96+cGODcX8EcKoWtSBrxz0A10
UcH3wWJPPX1qo9y/UbDn8ZVex0ns++pfM8QltCykYZ6OmyTmOwiuAuV4xffleciP
FYw4lTzmDOL2rO0TVB5agcGltLN/Sdk4t5EpLVlkVqGTF3CvE1AJ7IBzXtRmHD20
0VW1CIsmLl80YzZMa00sseu6folINRobJ1uSdRLzzCFZ6JNXzRtwYbzC/qJzr8Ot
8HaoQfAk/5nnBBzE23Lb4bFXaTnsxxa07u7NHpyXYKEtP3UXyqrJmg5NXTb27otf
bN1qE2Mm4Zx8MIj+RQoC44Hlxx8xV0AMJt+F0miV2Mkus4QKggAgjbIT1/Y5jhqW
dFJjGjz0HAGHriuBJX7c51nBC+O/dPPEVtyZRQEptPRmL/fJx8odIMDpGYiB5ws/
7KsviPmF0UvWjCNTNkEu6fuaVDG4HYlbYmP+DqS0PPFYDyOgf1pEt+rZ8U7F1NIp
0+8om8YdZCSweqWfzlNIyfvKmqJuGZrz66Nap8a0vvH98J+rs3/Zl/7bh997QC0o
U8TF+q25lDP1MuPTsFlnNxAAF4DPoNvedoJAJ9NzAoEQFkLN6pcQXjuMjejrDGi9
F7PRYt7vAavim7odZH72bogN/Iej0h8g+S04IG2Y53sTkKSa38Tvpuxl6BdRS+ET
xVXEJdlS/QVVGm4/Cvb7ImsO7fdqhXVWMv+1HUHWqat7gqZOfzQ5mXjs8JbxjcgN
jTMkXy38+Pq8dHOpI20adAZ0gTk1KW0+A075V48I4PEU85rMn83IEqMOuTxnmJHD
9O0quUYw0m5f63oFMnn3+PuBWw01AYNA9KmoLwUdAPz88hcSSZjhMQBVsmroWoPf
68HeJiMPoI6KfZ+PJUURb+Do8AIrG5cP3rpTcFELV3phWPwgQ8GfpgJ1mqQ42Ma6
aBbEYbaPiNq3+ybIAV8OW+Dp1F7W4kpSqWkTtiLpYfN+rtCzEypGCzMky2BRrI4+
gBQOECOttP/0Gj9LUoRhL3z5elMsjcsttylNDI/0VN76zuE4bTmLotApswYAtzVS
gAbbDwAqJ2jGRMszKyk5q6+29k6bEeWRyJujMC4fW3iXu+s5M+6w91ag5KrHYxte
fpDFh4Wdjhy5SIvggJXokyg8p3RzlqorAhHJj359Wwu9uZzdDhly+rJ1DsUCAKkR
YaZ7bhseYctkqk486yGS3wvvmmaiMUm6j7dtZcH3Il0l2H6cYlC6XL0+GUDSqe9C
n1rgjvVCtv9KA/7Fii/bvVDYwnTa1hKbEGTsDAXWCsFd7XlAQiUS3kh9GBoDk/Ol
eW0tsxsAjiB19UUVLs/urDvHaaLAD/ScRpEjFqH48K/gBU7jAUbyBvdFbSjk7+lS
vvYXlZJjmSJh9Xh4XW83sT5blgwZfSuTgxCmDBLeIduExqVKLXakOujKt7vCLwSz
qRFN1bum1XFrKciw21llwxRfvRGijWTIblbjg2xHvSFUX2FEQ1AlLljjmxozhK6U
t8eO87BaChPiy47Wxp/rLyP+dhf9atzDS08UuJ8588574r/KoRG4i+2UOZOgQ5PO
F4K82UaTs6aed51Bt8/HCm+Z/nEMNwC+Ky/ScM7CPmL4NEJtmsLKOxlyvGTC7/zp
bS7sMF0zfqrjIiRpUTKXFsqY6AmK/yC0nTas7VQa/wvuzk/Pc+NoZI7XVirM9JPV
h2BIj0rUmfQvN1OakwSUBr1bmrBRFpG+0Z4oKIFI5K7WzG0wiQKkNX0JRhZZaLzJ
yEm2iU1xjYwQQqLSVJjEq3T/Cu/ARXk+zrocJMLMzuFp6dCC7WkVSnV+jdVjd89g
SpyGhZpeTA1ayOxRGFCtcPafPUtJMC3dakHgoFEk9v5n8nbjKU8xhxupeXTljNdF
O+gagdb5zFP5N/I0PznENoTEukUCMPUNe5e+drxYZcY2Yjt1A0SHh+vkn0PZx6wa
mgVuFKxHS+Vvj75UVztkvs9x7Jka5Foccoe92lwdPp4ZfKNjBlhoDvHl9rL2UQz9
BvCek0aed6FMt/EO7poeO1UPjBg/UHP9/IGYOMq6GCep4UXllxsKgMln+d2vUvdq
dMzJVKyZkXIH7xb5OovJ+EXWpvGMiMfOyuiluSX5HN8oZOVoeDef73XeNanSX1B8
o9zQCxgTEhpVYrpKdue43UAhrZ2NBNQbdamL6DsnkoyUPuLSm285067zzw3u0xap
JA91f+eDs77Kz5hVulmetk5dG8wuqA6AlpwOrPxEFOZAZVh67q/hZs1dQyvzvWNy
yd3hfq2NoSTrm/SJey9Unb9xifYL3E2Qqo1PHlvpTr/6yIEReOgQVWZ0SVZtuUWA
MAtgZ/RUuIrqWmBYaZ1s3dt7UGiViofGTKt9hhlNcU09rOjcs6FX3XUQ20idYY12
aTeLoyrVMBuSgNg7x0OwcSfOHCTsCI4nAgcwkvKnj6RLT3oow5lrMa4zC6jPNv9s
6rb+z7KP0hA/a04EftVb/sbbpsevTc4wJSLHI8MQjG8LZx2mVB6xSSi9EUwU5uz4
iHFJgqBktJXWu/PDaCgf73ITLGRb/Dj8fLng+HWqdY+y2pG/0Wn++O3q8bBXZuQm
2NvGG/Y1YcddexS55QvnL181m78XnTSUa0b/SXxIjnyQ2jimxsr+ghQFIye1GWFb
kmkwLh7Nbh3HT2BUwGta49jS+PKndpE3abafhzQF13s1ycNOYhXhVbjF/b/Ce6L/
NerhqPqUOnAxd03EP2TzOXDz80sLLnVbda05H2qtCa0BEvQsoXfYSDRrnGMby68/
1LhvUgoJm0labavZrL4QNsGB4wq30LuR6LO5wWXW8cKZOw50tZzcxWtO1qgv81mt
hWGGfrB5EtQuEyfCzZ08lK3QRThChggIoOU5rMQuDJkgcg2NHZm6C4HkJDA7HV1V
uppqf0VXGE7N1e2NospgtBTbbj5MahPt5zWtZ+xWw0cvyfZHYA+xvtErtibebLJv
ZOj4dhSGUehQtX/bDrfNix8DONeDZnmKKvkx74YfigWFPjOBlcoarp82uu0rIWjd
jC5ZN+uAlC29I9O0YLRleKgV30kamx4bScDhm8OTNMRKGth9+QrBpB4zusdBZ6Va
T3ZymVsPLaSiFvlMJHWGaoMmEEqoiEOhdFP/pSWAfaoikojZQATxOZFaxL+GzkX/
il0YpP74h+WwRNbXGEOYe9ft6XggyuCR9hLUkCbz2ZhNnUpFewtKXe5heTfuogTN
OkVsyrw2J6X5zmMCvTLENYRQwFu++gjTECOMuN09cEZAIEa7h0K4jNJA6jHeJ7+8
VIaQakbT+jOcXdv0KOVPF8bS3a201hpyoauf4Sj+ep86vYeCljlm2QPzmTAIg3UG
f61DA2ZXv6v42IYB3A+MVr7S7fheBUFwiaKREktW9nuaLZzul5kqEeyV4u4QBvcN
A4vDRKloli4PDPNB2w7E9g3NrTB4uZrT8xotJPimN9TElXfcqAOhUkuIMUnaZfjl
dALk4gxqhxS+jhiQnU4aKbghGVXjTC+iXeLNrIFKEbVaMubsdkygWjfIRtzhDioC
XhzAW3rVGjS/IyEzWP6m7csjjVIG6e76QgjPe+VuE3Mp16xJVuA1JtsZ8V3GQTA2
rgigTc/ydOyXrVlVXUgHoeNcRbr8ONwkijsCkpwx5PCgFEaQfOZBqLb7rpi1KvTP
Io63E0kzas2UCZEmZIXLkr5kMJPw/+k2TAiGvST2mm3fQLMikUZnsLMJg+PDfsrO
Q6Tb/j29oS9VPcO8gmQjWpeFjPmOqTixpJzBGXVuYgPhikGaTRUlAomcnAjf71bI
8958mld2fJGAWe0rgxQU02xqzsNlqEB7iv9yq5YwwpinS8rgBdt/jflFjkXamRwc
IAKNn/KGayQo+3i/oBq5J3r8gYhNFW0QRCYoscWqLED43U3Azq9hzdas4vFZ6wAO
zbjqM4KB7OhymClE5bQjtZWgBLc4i8xBu649mOsCN3TJ19H0vdBRF3uTVo48cEJk
zEpGVZGJTXuNxLcTljPJohza88AjXyx0n8H/uddf//kMEyp52tqSN8n+flJ4IEIE
Jo+D8Vk/dYtloVsNfRcv06f8P2PdmYgy1oZ1fmx/HO2acuY86DMo7H2wbv4rAa+Q
0zK8GQM8OZZG/jggRYtK9anvqT7fEvbFmr0f2I3Sbp+QOrQn3HaqFaDiKQUd2/52
Pr4AxGjfvQvJDQW1KSDF4P45wRqoySzFmhR3qh43Mm4gEgQHm1c2dMCptc/IIpcH
W+g5VIFrBiXu+uk80w9YZQpYsjExGVr6R3nZuUz5Y1ZKbrLn4RVZB8cA4WtGCJ7G
wOOEuvnlyzIt/u+BesvWrzpdvHFtwH0I5leWQN8Lx8bjPPUVh7djd0wV55Gaj4G0
rwCNn9XkHIu0IusnqJugHClvqdCJC3Iu3Eswk0UpKEWksMtipAw/brH8MiKJKK1J
2OQJZ/vZwUL9YvJx2TI4XuTo3vGGM08zTwNXKCN1CH+sxLLYk2gWKMkeP6etB+7O
H8djrJoQcOhzM9Sczcp/k1JoMc/OyqPDEnMLkW6vqbGp2FwtKxloTGCuZCRfwZg2
2BW6pAQC3DdNP4Gx2hNg/RdSpkxEhAG1QAPhus8TSZLC5BpHL8F6h2QDBtZ6LHdY
6ooUI4br3CvdngMm1OW5/jBf3c1CLZGBfTdKGDl2IhoRbiGOdoGizXZwmvzYMoRH
BNNgNmr9H4zR2RVdJelLxvIN7wjxiUGOjmAikZEfAYKgeAXTDRUb5RR4oeFxQIq3
cB9tl9fFJPt4aEDWVJHxNpqz+1S/9G9aqlr+De32Y/LjWZeSEKG5R+J+Lja/Sj0k
Dgo2XD71Cj6wbJ6OkEHeLwwJGVRzwLwNDZS3L/NJZHDWjkWotNjXB/VkejIRxs2E
d0o6Usodb34ZguniLOiE6wEJZ+XIGdSzdx+pBPpdpL4D993WR2spUl5B29fUyLQJ
WL2EafVCwAqsTMhXhUHdcW26ncTnuxRZlrEnXClPd7iP8WFS2QleMmg+esVJhjQM
qSALD58MDiuK+6zhUGklG3oc3oAFSM7uVUvy2MMh8VR5NcytKBkwN+Mq2nHcByvU
0YdvmZzgtYCpkUkjpZvGYTn4ZZpxE/L1O7Y8TiDaAw0pxePg6/V/hcjcqU5wx0FG
4fSP1sIEepw6Tw7pf3+7hBOLA74j1069FOKh6cZoXz5mr7rcKhzkYxGamMSqWZYo
n2EiwK5nzov5u7TZ+QDC9/ijaVUlDvqqslrd6A6XIRHrMKxZcUERmokK2NSl0a1Y
nj+bXsBgvI89d0xetlMze059JbSQlMy4BUIGe/9bwM+p+lEjGRD2xnm9FVJ+Lnfb
PTr5iK5Vqt4CXnmX7qDON6ywz0BxAaqcQTydW8DA3la8BD6CqXvOpHM/EH9gpCaT
QFZKQBlY81Zy0EJZjh8RuKrG30KL6SmitkYKN9nARe0GnR1o9PHtZJ9yBxAOvp2A
8bAly0nx2XTBcGyCmLqHuKffOhKURqrU2FLKuq/VJbRpMhVmSibFm8o4tgYw/Vl7
KFCZlToVWspCZ7seVHLzRdsOa1LT2uBP/uyZNNA/hGO+AEv4Eqp4jyaB1H64V6dE
ltfjAQwUwtiZavLoY6osm6LIm0xUQZeibwc/wgDKJmUF1tzZ1/OXlQ4cepYB3MVM
ABMGwkH6AtAM8Z27kXgi+DKEUW3KQUCOfpiRhrD5Wt121OqNLjGJOUSmd1DppMlq
Q6AWvyuKwOn66WgfjxL0IoNcn3Ew1jw0lmW4ygznY9arQuNQI5zku1j4xdS4G0pm
ZAocnT20zPHrjpekikf7vTubeWhrIEdDK2xJqyOZImFQTOYGPYLkcyHCJ4E+myaT
JhfN6mqqa7hwvMJVoQAcITO++fd14WQyri3NsBQ7323KNC9qUzYzroOaegQrRWv5
3edYhLiPqiPrTwK1iR53BfYKrPlA+8TyS7x1IpckgKm7gVKdyiQp/eeO7cZ1e3oM
xs5AyMNDiMPP/wvwYRQVcQLrzmPS7+znHnHPYyCRRVAhmDmL6Nnq3tad46ymK3zZ
mYQvcr631qk/TVSrlsxJddcpKM5RsHKJZ/h2Lv2r/YjjRmteHNbvkg/1TeMACyId
1Y4R9F+2CAgTGbDk23LVK/KQYfYUGjuRLFlVZDcV69m3cpeVgBoTHW2CrN30/frk
EyB72wkxXMAwzfUTYvs3W/HwSAJDMAP442W0GNnpEEjO7l4cS/zrlBIsnbKV3M6i
ky5wYVBMHR4Ucj80h31uQOVh4R7gSfEyIZY88adB+Kr4Ah1bDttJKXQSw7hFO16v
hAe4o4wlR0s4pFHdEjH79LjcOqLecxXcr62XgGImADtxck9RWE6zmJa4XWXuDA9D
Dc5oJmHRU2Dn6bCcV0u3bDYZgwJce1+RT8Y7vLGA6Cgll6DZiu443U5iqgpApycL
1lk4NYwoNArqDAUSsc/rvc9JXHMMkIKAAFosE3ZvuUuE3O/RIkIzpCdGvmRA9a3U
LNo/hLaLTgfmRudSNeTXAZF1sENn2H3WXzvgKrvj5517NYwEk5T889ADoHEUcN21
FAHzicxp/kQRq7aaed8OvZo057MFRiuSz6Zvrtx1cra0p2pzlVNnk51A2vxsbSes
hwb6rIAbrgVXiDoTTw4wq7IY4LwT7cFtKIWre11tINs4yNOTG8HctPJ92+UO639J
XgCD0m6AlKXOmk7Ue7bNelIXACRwRECtOXUckM52h5Iff7QAaweDd1M5TR2coGGw
J7it9qOeYsm7IGUv8ZKR1RJ8pTwnfKnD/dmm2YIVQPubOkCXdoXVt3y9djskOlxQ
HoKNON3/IeZcT342237hoYxhjUkgdl+NLnAhshIxupLVYoljBGlbbhTEghfa1omv
m4kWUnEGZ7xLjMV6dvK/owb7PHrqPRcv8YlQq86ti4RnplaHZsR3QQECDgPUh2Nd
d61uYjsOjUi2VOaQxl6OufihTuGLKGDWBUoVGwgS28RgreVUWKFC2FZT4JTar0Jd
OWTTKtRcsP2hdBLjOCaBwNArrh9FWOzMh71fBTOZmcaYg+NIm2Imjo7KnlGFPW4e
CwJYFqnLkp1/u3TsKYtZwadVYv34URykcwCG/Enne6uiV042oSQwk7zfQzkb+EfW
8V/JUNwJCzejTF8vkkyRUNtUZhD+g9m930o72lgMqYvd24kKt5c7vR/xm8RiaZ/T
PbY8qBJry1oRIZ39s0x6sEL/jS6exwvRCWUnJaHwYhs73v4kfBA2CYBfI0tyvS63
1BmOqwpH88Caa7F7L3AOlSmBV3q8/6IU4yBJpubH8zQtvk86qfXA3Y0GuzaHBUJd
ymxLaHCAt75T9U9dacQIIi3lj4l80ai86aOaKnzIHgCD0nPVjkK7XZTAiIO8c/a2
rUfePzu26HxirtrN4LxnXIXfnhnTj4viIpZCwd3QBVcmtxLdF8gjnRfUvEpvQboi
zJzbjn1sWeIpkgcvfFmXzbZHDoz0dM6yGL1qxcQjVVifjH4hlf+iXwxpuXGsoTkp
Sc4HD2/dGdxzq9ChgvyVMr1K8PJZsfdQ8sFsY/l7B5BM9QHq2jLg7hIQgwIUuvjl
S/koecympWyIYasuW9MLS6lywlysNr1yO11wVJZvWyAGddsjRiUAsMYiiC1iZhS/
yLBIrIUOUuziNB70y5fc+T0+gG8LD9ykMLyKbKdtIz7cGr5FAFFs9qEhkiLVh7UF
TndBDfAsz9JrBWjplpu6vbX0iLKxHCalqPzmySpQ6LRI+NtcITvaAlnNs3i+KTUQ
5FIH/zcX3yeprdGsP3o5k0Z4htMSlaunHCEsEjDU3GhEO1fbB0uXM7QiAQ9kzPuh
wwnTIUV+9KN4kctlB61B+7ZCefg/oNMKLJuW2vQwLzF0I/wn1VKm90zHnqJcX+Zd
uR72wBKouylHGwM0MyhYWoj5+hWS4ZFvPU62zx6JolSuWggNs6RHRPBmB7ODw2xA
YMgTwChQSi2D4oXH1ibz9ALeiJjYBHlxNl6AdNRVyL+zJGrCgjNuaklROwgDEyNz
SNyNmVBuLYfBxDcdhnAp8g4f0sKFpb9Xvn5HR4lH0HALZlDHWFkIQzC+K77D/08j
BGLCzcsp1Jhl7rMo76eeyDmJFVMMTu6YSuEGAoNocAvS1maMfqRrouDK5y0lzi77
7KEKCoLi6sT7r1w38E/VDiZbBQNmZf3qeYDC3cXejBEFl5KGmvIwIlc6bgZvU1ww
nbpfB4c7bECm222zis6KfWZnMUZU8cq6MtFjfmrjUv0oTw8zeHYavEnLMLJO3GKG
CM6uHdDOAb0SVh0jJB3LHi5Ha6ZbP8G5lzbDOVmXHkat4V/Jf8ez8qXgSeuKLEce
5pBvhIcLJ4i6gDEYzxIeC4uGciMEqS2NTz/sWBGD220XQKDCjzWL4whRk/ijHS0A
suF9TpQp4CuZEeeHvX9DSRgwPrAT6jiQKhSkE/ncd7rt21K6Fh2MrymIPZqC4BzW
7sz51Ejxoxag+ttg+fmTaRlpLQqyx64jvLpLTD+VlAx0ebzcxZTggEJGNaVNmFNv
WECFs0Cr8kRimUwLlXJdEwP/0ia1iCOi8dfG60I//iCELcCimKcJnzmV9BGIwPgC
c71DrA/k/yvFoVZ/XNE1i8Bzfz3X8HeqWlaYKwddPfWM4LRL2eZA4/yQX2VVIjhL
hA2X/n0BJHuRtzXZ6wIj9G31PfuQ+DQkSl5jeXXZfAuJEVw96pbfCBs6g9mnmzzs
d4D47rFUCKCTkjBlKGRTk0owG/6HJMJfQd2Yz42UbgnZ4+qhS9+iYWE4AQI5qpV2
subo8H2CDsWmSVJpACzB90QALF0j3otE6Wt+3MeTCXoSnJLdTpahTwckObLKmnDE
+VptD4gVWBZyJ6gVzHSpi8Yf1QRB+srT6QqVg8bHue0L2zJyshOAUrGSgAkM3hMu
3b1aLRO0av3ThuR4U0g1pqDBJh5JH2Atrnw/A7LQikBu6n8VZbsxIJMvnXJ+w+UD
INDltiugakLAbnIp9+fcMIB9N/i3NnkwYNwoCv263vEFTRxfdLKJbdKeT557N2Uv
DuZl6oHC3BFb1WGdRLGrKLpALD3I/41Q/eRYxW8xKKgPDD1em5FfcTfuH+T2ba7h
rp2Yvm+wBmuQ8VlpEipBY7+XejclepuKu+rve6vEaHzDkmo25MVDWDGYVGVGYTSM
cF3Gsg3kEBEo6IjhOreZB+Aece0w4BReF9u4HIbHGychaRMeB2OfCD8B5zBPYnH0
k7KwmioCVNfe1tqN9zy2gKFzYSfBhrhJrkv/yUc3CphTnzGqiA1VqzP9VGG9M0q/
xMqCW1PRFWwIUEfkklupPvEaJR+ljt6z58b0MgJDtBIHOsg3TD+gMY2rOPlEjt4e
HZ7wzqs3sfLlCmKnKj3y6Qw7slhRaK77ZOR/GDWmciVHpI1V5aSCtRLHte7PMkXp
F/M8i/KS5nUG4KtZnVUFCFj7yX6LK3qwoRrn7z0HmHNK28rl5N68NHLtEmHeGqPc
LkUIkgLORFnatYCaeJDYyoFCZvC2nWngWF4MB/kgT2BCPQCkwKw9fHmrwej9OAL8
ZoRnYHwey4A/MD2/QPSdC+PznE8NZfCPJqjAOMwjE8RAiDjNrQyjs8N1HUQMcPvq
LBsTM/UP45uLiRmTxOPD9UfrhxlH6PQKNK/M2UR9MyVRoZ9PdYGUc3LcotYXz0v2
Tuw6iBJP+GO2BII8hM6a042ZQSun9P2IXO3VV4g19nGs6OTOs1Q13Du58lQMURNZ
b8ByqrmvErELao/SygLwi5FT7C22x2QrOM2IWIAu9FvkjmMSr6ey9AStN1yJxa8f
qcz4K0oWQ1WcClC06xH1dYLip3n/+F0CszsI1JEj+rx3hZe6YTZ+DYAuZ8rieHEb
9cxxHiiy3JkYAsf2UMRZ/tQU670jUjNaWHmpFJxhY7nDS9Egf5ZCkZv1Ql3xtpq5
ZgFE7OMC9rWWmbhSBYx//Q1050V8lgezeJUQFhEwxvISju++T7CB9C+GBPdKRBmE
6xahP80RFwKwcxxhpa4is7vKohIbr9SztXhQNQEZ5UKNaOcHvazveN03mIlGKkgD
403IjOdjVU/zEmBNtGyZy6N4/O0/nSc5iJjcxNBGGwLCTEt6GrMl421fSxyQKlod
FSUOL93ydAAlngKeF9mGc52bBK3MoMT8NrYH0qQC3/VAt3UPW5ugdYe+rM6a0woG
EZvG1eGoZr0ZkVqgz8s0//8d4Ue8T+8XYSgOW28PJWC+a4J8uRHW2RH3j4eVzpwO
eCr+maSwGDCzzUd/OzvxBrnvYcUGbZsYRYSl2t9sOwS6qPBGolgc9zS+yqcRRB8u
o3sE6gFLBke1OTq5Yne4Izj57mo0lA6ukGirbaIuzJRNRU9QoCW/GerhCEYsVqUL
X4MOOY9lFApupuGHLgAzn2K2Utk/CUTFtauuft7zCVMwKGHhYM7cOI/E888EnMkF
boNAvUcIE3qoQtANIsb8Zz6YQJfY4XeD+Fuf16Erf8g3aJ7ALbLfFAtcuwcCP7p7
WiLI39OfWcW0OeCzl1RfFZnNhyfq2KNu0r1S8uC8SP+E1iiyqeBzQQdkDDnL9vUh
xcwg++YwzoJssR9/8uxPzrfr2s0NoaDO7kUiqMczeHTvwlXpVjoC+jARuFm36mjW
Rt3czMWxCtqr0lsJMwQciY00ZVwh3tr/6qw4Efb+Z5NVKVgJ66qzLC4VeKtGnGs+
U+BwamR9BbhcHii8vs8RjCHLR3tdbTeVTws16zO6KEEBbjCdb5Rna6qnsSzUVYRv
/xVBTqQvyA+AmsLOV2mWiBxV6yhLkLCO/d1cMTE0P3/hY+WWRht6S0xznynXOH44
Xzongc0aaZv2HfdSSJdRHx/YYJnlxzcdiQDbgCtWcAx6xpWNXgZqqbCHIAXNnWk1
KCc7KVQY5X0a08StstgRfbJ05G0RZZNjMyQJZgAv/qdkl4EISVhw8rMMhtep1j8F
fIE7MG+R9n3WE0vvNcA+MZwYjzcmdzAvytqHUtXP7cjbZjbg7hZviaambxHxQN2i
kmcyuvAmYnj/5vZ9NyF1k6biNxq65mrFzGCCSdaPvzbmfGxEs7jHRVfUuWlMlL9N
R+o2WKID0PV6c8KEjVJHZ9y7YB2mSL34dv909U/4SK4WlRPmRH4iu3RGeHdKNRc8
F9cXD5NRZyXDX1vvwJhkEcgIqEYuBNq/3cm/XFJ1B/QsyA15Fy0EDz2z5FPv1pGx
TGB/mswnESSIZst5dkxwdl6AGeRIxW9HItLVaNAJfVrUIocCBVXPFhmztJ7Za6v6
IHa2zblMJKicYgdjA+d8SSAW015ze4V4Ff+rJqisdt45bLzrQOmqrCZVsWRG58SA
jopsMdaspg/2jZwuoW8ChdioSDKjKo7zpvUGTe2t9aSYoJgNzkKQ8xuvJUj38CfZ
/4BYdlT+hYT0zt1aZ2QT+fAl8vH/ikgDYftMepMsNLFaEkFIXbH2NBjYtntDbnM6
bAk17jDa3zY8Rt5Z4w8GaMSgKuIx7seKa9Tgb2N/U/39i2mH/Paxfusf+MYmXjYY
MICtNskvK4h9wJdsjoQzsSXp9spwQzWZZJm/aRu+kfr4kKRdNjearWm7uVVnfifC
aPhjzbXxKzsCo/UuqDv4wydnv7YCBotRAqDmIRkJZv8bmu5zi09Up5xdRALP+7dX
RcblyUFSLR7WqcaWWta1KiuCfo8GFtP7sxNIZS0dcHkYZAfreqxylZ3YudAF8cma
O/qWiIa2N8TQT3+N0lczgYXYNlc5/asiX6Lr5hPhOJmA0wvxpg/JyZ82GsGLAj8m
bk0gFvAq0YGfo9xesXTms3DRA5MBk5bMcBWH3vdEhTMqKK0/xoP7yl5Qe+v6qQcl
F8RKqBgEdCgDUgBj0oaNDC0v6zTO5yL1X4XgfDrX+ybj7YleSJaui8KBN2t29yS6
2RRrN+W6AGC+D+MZjzmAAnVaRvZRYspn+0N61kSLxtzLkkvmZ1nC6EGoB/enb6Ck
yCMQJR/L/1TttTd7WsoV7iCWloUNWyC2oplMR/YgJKo5YAbMRNyxhWPnBing6LkS
8UdBaOfAbNwSCQylNjeqDfHZBHwsKYuESZ+labNKhvU074QEyyBrP2okiTo3zU+l
9IIdus3IUNhJjsCIxIBh4dgAo281i837kYwhEbGNLM8zNpHyptPPhq1Mj3mLNc9b
r4tXBx1ndVElIn+a4THNn/YF0MnOnJ2vh3vf+tOdB5YX30ypJyHuVFrY9Jl/9AkY
gHJtLP3MklW2+q51sUi8UeXHO+fUB0NPAD3LgQ2atKcMpQxPE6g5ygj5RTihieQL
riBl9JnD44qdCxjXrhHDUjliq8kHxCHQFYwEf0Px3lfW9T+boIsn16940+6ozWgo
WyTQUIqAKoxkKxrLd8Gt6AGyQlhAxyM45uT4IZ68lPE13LP8w1IhUr5Ye8VINs41
z+mjOfRqDWvdkINoRhGdj5Oovr7D5X4i69/lJnKEnqMMPCtIgumtkcR4gnrVwfky
6s6duWElw/pvvJccnEdTmuy3IeLtJ98f9JZnHLtU8y09qSQX3jXTAjKEzeEeMDAR
FOd39uD08NPceqqaWKYJpIDl5HA/1UBHbDep188p6Y+z2lHETJtMk/ipvudDdA7N
hXl2iBtLWrR7TkCLPFz7tGqnkUccTjewkyFsGVE1WEEEq0BEelbptL9yaie2eQdX
Ph8NF55cCZ080sed8/4/SWn19He7zf79a+BV4euUhdflcIZoOjegSxu2AoGTL8Fi
Mm6Hfw0yux7MR/kAP/W+LmqOHmObdyLMJMzz5LwJEtf+2oDa2L1GWZkpNfP/R/gl
UMcr8rCIRW3kE5qyCPyDeQ/D3PDD0Pppno/ndIHXToilSGJdGM+uVCfcKNTQxxsw
4aL5d2a9/NZzLmCDA5BbnOVhcexPwK3/5mgNKq2Zd4iBwV6C/MUMSZR1/ZX+ioR/
xPfkThQl0S9nH3OaVfl/JTo7wRShPUwzJ2L324rpwqhJMpC0f3D3r0nGzTaFv6po
Yfx3c8269+h8Ne2tq+RbFv2LlO4qGAFwusvPCqgZK9DbtLSi9B7Swa04ys/shl2/
OwBw3vOJSWI9UB6r727jkfG4rpJV+PI8VWO9qCTDP/DZXH+xZbdPRFW/qRhvFW0l
OH+FhcSsmEb+zgaCfHq39vFiDzezzy2pYUoC4uW0a+dJQFJwqRD8iOWto3lU2F8K
qw9fwCiKzv84Ssr9gWuTPCUK/8cna85vWomYN2nmUeo+6ZuHfKuQwc9jkzKW/6Z0
PTvpXkhvBzYt7oZ7qPHoePPE52oBoktdekUpiJXvfIFOCq6pmBwbg7KLNSe8CovM
FL2HwifudV+F46uS0M+9r8joNH6mErsal9G3IL1f+mZ+d3SVSh0bkKXLuT2iPW4M
oo7KIyliYCpDUgL/tWvzq58/Fr/RrS8yqbrtebgdYU+Ojky7GY9YJJ2WbPFX8xnB
IERrM5PXrSMDbblAiDJ0wQ82Hm5ifHsR3PGpRd4IG/JAoEWApk+Tb40LKvddt04Y
3v6XOWaGd3vOtlpGlJZOpAWogfM15IgtpipB5aJJd4/lcQbi3F2jm7JOD6Vbc3iL
RirfBA1RZJDJD28WwnRUZvxu8VaLLjZ0ttO1+QfZ6ESuSS7iZviEn5b1iqv+SIQi
C9skcnU2RxRdNkBRpm2DEjVLVfuhhMTzZklGZvjovPtzodXOdPSFbCrgZqhbnf+W
9xt+ZctwA3VkTA0a+RDwChpfYZ4oHKsYWeW10WZxJboYBYp9AUd7ne5ss2uTe7q8
Y9fqe4mKWqE7DgaH15qSsrgfT9W9WCvOroTbBZSER+cE1GFoKvvlHfF4azaERTzD
ON/S0sPRx9YJbNdLoMmcBPlxDTKsgYePbWy406tdIeIH3CcjAi0gEgT5JSG8RNEn
1u0V/OzrpI/slEGfgoyTX667IGxP8O7gnCzbqb/FKNAlxF1eB3pDRP50kOMA3ICl
sQa5P7rdT6Lha1RATnLQ+KOyMgLPfw7fqjT7zJ5VLnKhK4lGNkIndfW8ZoSrWE0n
ynLGbtBvTnJD1SZs70CQ/9Rf+8hpyOcjAxXGUWvdDWGV8zatduE9S2QedGGErLTl
+xLmr+WqS+ZUlQkITlUa4RIpxsARcbfMogHbNPXDTfaXld+chS11qP+y/36z54qP
S8oCt5cNkV+7LFzlKfmBKA0RrHq3EvUSC4sdXT+cGxpYBIj6sF/1KmrN71D/4Csj
qGxEJKxODQMqBgJRt3A9Zq9dUXQLTMR1fo7bd+2xGoAT3exHGBv+eLve82rKNjOc
TqdbHF3l5CmclTE7bOb81aWHEBlYnvdZrlULPBemqRzlnbfNZ1pPFZzlAn2Yezdn
udmGkAwH4hT2l1otQn4TNFMBcFFg7eDjWp0L7iVddQGpR4cmzm6u1JcV6SxoGLks
DHuLr8uZuXwdPvmWcbK0VFBeOjIsTPaZ8GLam7NEP9NodUnaZlngf/xWrlaQ9Xrp
jd0mDz25OahXq0+GDsnyvlSC9z7lA/I+/DU1adJ93o9zFeiQapPSlTF+1RsXsDWT
iIMQrdtMGA09EFhdJMM6Wc8nI6vMySaut2KIyWkPsHodxyOmM8EzC82rrsArlKpc
83SZDRtmj2hi0f07iw0MRmCj6HZuWf2WruO/omdmGb9gFP89zjyCcqj2KgDrhAp6
YF5XVBV7NYj0YUKTVFeIr105f96easggHyPo/j4m0VN7IMLz42i5zH2lq1xWLDuN
iXLVfy0BN4UOwrdd6JuyBKMpygpFHHsO3Nt43parYa/OxUblCjGFc7fU/6R2NYH2
9hwiXI31iq6qgwUuNqY0iIq+vHJ7NdetAuw27J3oGs3nGzIztVB5gOWSz9rAxVuR
esRosJSEyjrQw4qGCEjq8w1CvKo9PuKDfQN/EcG2oeDUVOp/lUoF5/JuaEd6sw0K
Ux5SAfv/aCZlct/IiNC12zGqajfaZreyFE4Lqr+h+Pat9nkD5Y1zfEVwc+zPTtv3
lYEYdemQV1ffKLypkGSK65Y1oVSSWrEKC07qESyVCv5G3k7/oIHxzOnn8PmLl120
qZHwVs4U4Pc1fqPzJiZpi3T+U3BR5GgF8/pDrBZ54SG1hOX8eicui+RVZzVPQUNP
kSBthIEG7xtgqs8rv45ahq2TXUoRtBIGlB8mtiHO8vFG87cn8v2ACKa4i9gZraVn
lPZFoFE4zYKAZfL3A5VmaN3J+XMM+BXBMhg1f/HaLGZRs4IxAM968f47VYQb2IFm
LgebtXL6GWO2VmNsoBujmK8F71MAJ246je8VOlm4RNDDihsEFK5mF1XTBJrrKMBh
Iq2EbMfwc7uCou+oKTFhW5VPgSa+31RTQ526v6aUTiI7y8Qx+VvUYt/557/GxY9j
et7FTR6M3bQQALTu4sxAg0eVs3fUmr7fi8sPe2jvtCyYx6UchA/iXPM5MNBX5bhg
9asF8smyPgkN/+ew+8LXWxzlliuitFoZo7WD2IM73IeOS7SgMIexzmgKpflTQftn
nV7K0OEjo6Err/NqIYoGWPGl6hGwgNtNUkik9A3yhQlx1RojMDNMmLGcMqR8iDIP
2dOcvs++voBlqJLyZdAc10FDTqKIICXIrxc3J8jDiWAEiSed0wEh7WsQXv/dVW/v
5irg61RKfcNXvgZBqCF1S62mInigWZVuoEhyVVuTYMsLatXmIuk/07ZnTD8M3F2M
v8KhOfuOB13ebECrgKvbEFHdqAsDCuiiZ/+0xO90iNSaXa6R27rE96nABF+x3v4V
AmnCjU/JWZlBBZscwX7XjHfJox87SIzWjSrF7Tqvtpw6ORNDimbcAn3I44qsdEnR
9nVYfHTeo2vkQdT6svNOnu0kCWIDMEZ6hmNv/J0ebawTvCS0H4ltxPZdu67TDSF9
OvdaDIvRp9gxQE6vmGl7VSFq0Z+t0j5/Ru+II9TSt1CprockeN/KY0z8AFj5t6LU
exKhqDU9j7IOBU4oPtYlF2ZINlDUaG/DKGswxudv83JzN417Hbuntb14uzMN3qej
q/HEVhmnCXWtr3O764lMVCzYOhYQ75QOfl9gpFrwCm47wKnHfE5+U/DV/F5A99vg
4EC3WNDuLJTnMc4P0LE5D9HjyFIX0GpXaVV8bv599I4EjL+vwph4YEiDMb2YeJKb
HIfh5dEkWySgOBxjMCa0CYUy94At5vitLNxNyEX8sxmX5fQOPTAIPrSfIcYunRqd
XV+F5WEzxEUN+Mfm/dDO/8LUh2htYp6ES0NWvfhNOej5MQasnIfWtQXmEa+dOab6
pX6zIJlwrdOw+QF3akSlKg2z66GqIY1nEk1pVcGoJ1i/ySYF6bbCD6CcgNt7eeCg
GYSWJR/gMHbYL9jErO4EsJlFQRRlJyfWZ7OJoSWnrH+ogycPO5t7g1prd1jt1SM/
m9RwznkEOa4X2MvVXFaCR7CtQLq+8nl1NR2hx4aLpoGaSS8A3icKXZyLXjIX5KRL
SVZRpQynzRW7YPeisvqvwGexsOmYXP+TzTFLwDsOqlBm2He0yH2NsZ8kVjOMvpn9
O9HF3DI4twv2NHxuaCglaQrayMxr6oa/OR9+ulgA9H051T9EyTwONOjfnS7YqTLD
`protect END_PROTECTED
