`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o4o7yyWUY2EMBppHwdfYoy0iaS0+tClSGCOc6fsQPRm05LEBZ7MEXSveGIRndYk8
4UeVmzMchTXXxaOPWKWKgbsYqn3nkJT1vPbM+P/eVrEYkiWfuyps7QD5Z2xYDvtQ
pnZZu2Afj35YpDXM/eAfyNjOm/WJfpkntf95aSDlxg9v+rjau7nP/EE804q/fwxG
VXKcYG666EGWYxblMlP+4r5R/LIzsd6CoEUwgZ2FjLiEDyl5Lvg/Pf+CfPNGe54+
WPyEXpgGE80fUyBnFHTtNM3uqimTMTqqSX47y0SkXDzQxwwrhExHkA4yAbuxyr/X
R2SpEs/2xRrvz9eWhHdylZ2iPlhCJEH139O3qxVK5nTKSCLQ+UQWM1EvkNlgRDIi
SA+eGA1AsYp43lq2zYySq9R69T/eVBcpQLhn/Hc3Suc=
`protect END_PROTECTED
