`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
myOGuRUDnQJJqP4vHhsiDpYG8tThfFj+hbvaCTbw10JFlaTN5HQguZuTc3gto4oR
WAkuUtWErZKls0Gyf03Wex8KIczxKzXCWek9ZW4GUaCdn7pkPh+70HUaQJofqrwO
wdDKtHLTnnrNeHoQSTVSNmFs9s6JcH/mZWq+RIKAMmIFxHrasG0Q7hCqiy8Mg3ny
a+sRY+7lGvw3gZ+pAuu9thytKUAsTeeJoRwd/OUSeu/hy9DqUz7XNSjqEyogYFyY
05ZYQIysKHuAwrhkof/NykSY+zJFx0kWjTYpsK6emwpWn/7u+OlIqIQAt4Ih2gH7
9XDHfbxb3CQCJsvQ+q7XwaQ4PDjxl8mHa0htqecBEnQIrQNTk2aF1qeJF9v1+PVu
YSQbs8lUqXUv8xSQr9xg8vbDvBmtaZvgdx3rzk3TfEZpiq0GcKTCAYC0dbFl3NHa
WU1pogKu+InsIvo1IDEvxfFjvHXBdjQc5Zar1G1i0jYCdRg+KUdKOi1S42c+Jbp4
`protect END_PROTECTED
