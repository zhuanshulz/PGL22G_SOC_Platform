`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+xv4dswvMV95jHExJ0f620zaxBTtr130E3mqmhsv2ZkJcSTVuuVaOMrw5Yr/KOYR
1NkNuXD1z9K34FS5VZC827LQr0iMcUcgWBbYs+jV5IsW/wOjflApalMqAA/p06vu
qGo03IEcpB63fQWuqGpOV62oEiOyHOq9xT9BLt9wvziYvFKl5/nu+qAqyP4OBeHD
V23bQiOLEMZMiKlzroCzOXKYozqqQ3AKE928vWOqkryIfGwk8ipulicz5fdcio5M
bNNShOulFKbmPge3F1MPA/NLkkS3mD/1yHmQCUggJJJUfE2+Iyqr4zcTZVvWxNY7
soBCDgslY2YaBtvbAXBI+lJdK4zQBmkIknUfMR+JdyNAbASAR2jVVENyplCOaVAp
OKjRBB5LRcRf60nu4vr1gIRYArtHVfogwUAXg6R09/MG1SBMa7NjSe1WXsN36k/h
j98xYyuI5587LEB5cwxdoAFwzzZdaVRSrZwYqRe7XvI5+Hb0hbFer+olJa8+7y0S
rW19OAwn/tfjE4wLB34ZUJc72UiDNEEcPz9kQGBh/4XICq+abwmkds8X3ZKMtYje
9nR4FvaS92OPNFqf8bzepBiANCMcMg9hdShJrqAe6TBY8aow8pZ0KZX6Woy8Umbr
L5APwwhROqd2nDAqCpnvFhw0iZpV4n9VPbTAsrmKWvolaPAAYHaa+QVfe1Id7aCR
Mh4aJcVy7r7dxKxWK0msSVCi2VXUuCfApbpSHJXB7t0THxQotYdrlhwqnwJ9HA5w
kMdGDkbqrcSU91CbTaY5/YJUgXjtVmPDdDMcDNmy8DfJxxC195g/dRvZCsXGLWy2
j6D/YvoOV1ZQpxT0V26nRMLvQN9TQh7oyWiP8kyR/8wgkyQGSOGC45hQMVyqE0fa
t1bfmXnnDiC67euVcm+8Y712OslC2qjmpbIqzYNxjgjJgMnj5+Z+eMti88BK6kYI
H23aWVvw8aSY4j4LICLf9b+KblLiQNzbrbgUmflaawXkv/AScJps1UCYfR2jUPlc
mcTUPkHjTROcAHEKdUg0Phz7jsomtPVtCZPmT8igRyKFQBM/WD3LPE6ezBf8giOM
UJrTcg2CTnEOGqZjeL1/2jbGnc1LLv/p1SmKmn6LRZh9DSX+JsbgZEF75eZn5Z4B
xFj6Cpqoju9v70g1cJ+V2VB+tz2tit/+cp6AwOKxRhDh0Ga6rjVAvLOTPVwy2AV4
yIHGQIb3BvNWP2HZ2n4fibAmzKtH1A0q3e8+tVi+UivR85/cRhO+I3uXX12+dzQ6
XGfDTxVOV0nsgogHbm2JtLjAprU7APGt7Di+lKG5tkmqySNt6IZMKRl5X3SgjCws
b+Tp+B0kRlcyYZJT/Edq0TnwYo4A/h3XHFA7BY2nSH8PN0DLFSqPBoUPMxT8H3SJ
JP6yI3ou9Obke6NLb34RuOwWY69gOaWDu1kq+yNJHIoeF5WiM0/xNRqxCuB+juHd
/kxPXKpZXwJuKx4K+cf257uTuSjuyKT2aK3VbLjvToTkJ6M0o5MJyu2DbmzIxsSY
RS2fq6DCRDp6UYQkHSDmj4upwZu/8b8IKb2X6K6UVeiDQPg08NcuSa9IQDxFZwlK
ZiKvQ/OY4AQxtNusuSufbOyuG2PTJY+OzJNDjoLvow+AsKXxmaAvWZXClCXKuI28
6o9cfcHMrluWGkMOMHFWpyP0yyIydYWT0gQWVlFNbwq0P6ZKARZO/LvDG2R7Zi1q
hW4h+RCSeKXTZKGEMXyWq9FvGIC3IOsgKw/4FvFQRTP9PqkjKZ7bAbi22ZXkOEMw
84DMvR80+PsCxJPC5v1BA2r9vur8lsYvAm0MWSQdpLesUrYLJMI6ZZPR+6u7KFfP
3MBVVvQiTDE2+CuaQYhh5zU6Oe8xn7XW52EMGg+JMAOZYxVHvEDtnxzbAL+fiNZx
QMcreZYiDAyEs3uSp30bEgd42qoxjne/dlfRvMKzax3mw05go5D13S7rg33a0YSR
Hqixsf/CkcFetNY6QPRzh/h6AdabcrINAq/vFCroKlpOJ2garTcO0s7zmEcrqO7b
2Nii9qSTCMNy/1iujogBE6a6b1cXvJwzJSP8bYoC+uyoLlQDMveuxE6a7TfQNM+N
UmbEWnvYOQqEt5CLZNmAC5QXgTaUxDkiuhqbonYvPieznvYPSKzVFzFnvwbBjUSn
t3Br/F0cj0g3q5M6y+uzTzrOIC4rqRizLD3/Rutzjmz7JesDvL8Vx6ES45VQawTx
yndpRrRJN+ia1E2t9QiioVawaqNdhLtGQZgX/TlY9T6wJ1jEvV2troNsTK8OUYKD
pcim4UzaiyHGF9iY0zfJmrbe0qjIe3Kn9xPovR3Pw0dbDjnW/RysU3fnf7COoHW3
koAkWf9zYx2vKjeOaNXsRLNzacr4xTq/OfNa41aw10lef13k278rJ+Z095pweQJd
EnKUMgdNdRnz98ru/64AePVEZfgUsVZKjvxmXmVcJEnYKO8wSkPDCcVNK1DF1vXH
N9tMZfcvjR1PUIxB4JiXxY0FTH7qZKPVvsHhm510drgYe2P6Qw2RqX0ucSSbqE1v
rlXt/+J1wuFgS15Wzitcecdx3W9pLEJ4OEBek9G+YZNJAHHyWgAxWHAOvKQ62NBx
wjH7LRPKR0dy7Af1Hkf62TAtR7V6EuBtyOHAcVyX1Z9K6G3zc2eOTXvXVLZ6LJuR
iiwaQbbu7squUe+X/uyVULipDO9iH12jEx2jqYfEhlvoZRl802TsR4rkHZnckULN
TKPejMsiRNFRm8WAuWAjPo4hzSlmM2UC/f1X0RgYj3C6JPpGkuN8uYpF6NUrmNZX
x++S/BwdHU/ffiKuBYfmgbigLUF9OXUHuZKnYD0qwImWLw0QGFWWT428Q/W/0GQP
v8B4qhnZnOEwAw6pSx59PtTIpOUn9BER/koiClF92fW6usdqkYVNUWSHYfFdFCwt
QSaUDQKW90E1rOG+XoEUUwL0ovZujiTL9VQKaoR8C0/3dXu5nEM9sBJkeA2ERoyF
NumbTaFaqMMSJBlOVrpRXkZIdh8QSOEQ5bE+PsmcwunjlizcCcYoqhuJYiPAs/Nt
AT96jNbo9qKCWzAM4KLzjaaZmy5HDpZx+WubY34yGhPody57eIazNKjR/elVq2EJ
L3Mq/7z/56lE0KgHz7Tj1vkJzc5yORbqj8XjCfnbsWFauWzzPR0On9UuGM5YDRi3
h2zIeSd7eaJncDKvLVcEl40fmwy5BydlaebR6a+sFuQ3xiEllCVPKx0D0itzED1d
OP/c4QGOCROpKKZWi1sjO+pt7bw05GCRGk8U6wIBppkQk/XBncFgnIDp/9DSRuqR
X+g2Nal0VgkQL8aBXMVtBuYOlaqwMHvXNGIFlD66ABWffwJS9EhDKP8aQWQp4aEI
NRHkq6oFcHqiTq/9X+STrtS917ZKF312qrtJtCoafU9KSEJl+q2Y0WLWiuQ/nmSN
WuxvFTqML9tjGHFhKMS/GT+/igZWOPqgk1tRFqgAsv7CjF3NwyH+lOQYB9215kDp
zztRiMpjvpN57wGS2pKVf4wI0/im1Enl6QguLTuOCwu+FeQRS3erNJTrkpHX7S5q
vFFcoUcKm+xfS4VKKz3lr/GR4w2HorUrmj8KauBVOJXwQrl5A5x1SwOwYPN5wM28
QSMH5a/m8glnrsLb5z2oSxZlsHFw9rCoTEvwn690gXG3ryKe+aHzYym94lowzsO3
LdNTHYd7AP0rJHM6osxQwnJt4/VqhfwJyVFNp+690kYn91QGmvRSTsg76NISe99X
s0kR6bXGVlSZGmjhZtqDdJNaKMsAT+yrEGCvpGgTo1eM90QtIk4BhpnNehHP7h4D
M+Q2hV1Wj3r9C7x1xPAVePJXAl/KtGqeKr0K71XzojHS6gKf7eHOHZ60DyVIODxu
8LxlMk4D7C38I5X0cXLy12IR0/n5QiqBoL9k+cIQs+Ty3Ezhu7TakSNSgSMmotRM
kB22vcHNYy+BEBHiylEz75+WA0KjNdOlLWVkCDCQFL05WoHq/WGp3LOQhUwHIg/G
76ThNbEILl8BYKZOQ15aEssd3Tp988Kcxe6wia/E64yph+cZ+2/ol8+6x5ph+EPX
9I82+KrxqaxzAs0P/04iS3903mxlH5UEAO/6lp6IHoSwF94lI259Rc5dIcvDBfRU
xzpfIU4iWDDGWwoZmWq4wQe3EKhNfrieT7yxEV/Y5Ls5Qh9o3yfFQmS2laV0QHiz
U0b1oPBq5IyEaxKx9JHQDmlIT+7lnKPzIOb0QVC/g3oNjqpSep0uvoVOjRpZAycR
czjU+VAiPyqZV0DJ6YMIvp+ahUMolS1sRJbJZ76zBAAwNadXUa78F7SLwmoB4PW8
0kZC1TaOiVnivKkvAIv4vJTuogjouDmqSfOxo1eEYizaDAgUt6xtFsxVkJx5RSjY
CxnR3r22XWi04mHbkiXzLQDHKOnCGphX6pBmbRXNGfdeIVx4EbskfqKvp51V3B1G
dg2ZmV4kROK72Ld83vFqHUGKhpq8GDFHUgZB3LxObOFNZ2ZOwztmoczk/Au/A7Ip
hUjF03XzCwz/XVghENnEd9LotIdV1heG+g3mOLOPfJcpCLBmRyjJHSERXJ98kiY9
fzr5o1k4ZqjG/6B0b5k4sPlhSOVo9UIapVSd1b5v6AFbdoB+A5e2OhjYiaoZ3c3p
9iLmz97zxom/2ddToSSkHNsY0hqIXcwyikuULRQBCwfVcXdrPolPP9KL8WAuYO2H
BG9vaaWtuEYWpuPN4J8lofjlwrC/R0H+PSJJbrqrrU/6fX9gb+ioalU4EvnKMr1h
MLDCmZuTUU7+cHRV/RkEslpXWA/vQJglItXPvo8crvI=
`protect END_PROTECTED
