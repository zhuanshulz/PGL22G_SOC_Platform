`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ggU9Y+b7anBWhIuPr/SrxXmCfv8ok76EFQkfljyZbA45nP9utZ6oPU/WHYMKjq8I
juVj8a5QhCrkvT9iD1W5wQDLMF7INY8da9EzY81V3bFChzSyCzSQBTv4nCHRz0cw
k/Z03Z2WDiK+jE8we3B2ztYxjBNcOtOP0EACdRgFNdGkmUQYF38tf98PlZzScSPz
CE67/945a9U8PQpAoxGZmmq7I5PsXyQ8NwZKNu+XVzsU/FD+5GzsFhgNHtPiTm4v
nAiGY0AJnO03B0clJrvksvDIvE/O2F1b516zUKeNx0B8arDwU67OFE54SpcnLOIb
1Anc9/u+FSxFyVYtC3MKRtJOQSiWGtnt6B90+KUgXDyaPrOgCeD7qYvlrIR6AYbI
bXNNX2iWkAKiD11jxMEoWinuvn2ZOwYSWHg8QsEdnkI=
`protect END_PROTECTED
