`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vJT/gFMRUSVTiKh0ebhbVS5GQw8KgHf7nf2MhVRwnvQ6v/co187BB87NxHgHs1NV
g2l+A8+M+vycw8BEHGNnkZOOiiza4zGMww8ckHAcNmd+mGPY7WYTmhOSd0zfJQGs
1HfBAQW9VZVlUaPa2Ps3YZMM3lV9Em09OG33plzumofDCMk6KYW6OChvlZVGg4jR
k4DGuCNEG5hkmfUD63OQCJanLYbUbyPg19w0QdwU6l9yTU1iLJnJDDHnelfXYkS1
/2MkQUYiIer/HjOuxGC6LG2DxuLN6PgYmNow7lHZacXKIFy0phz87o2Jy7MVvpg5
OLXb0J/VUM3M6NK9rQgQEFFo6IDgFYuVSNn9sVb/MzKXn8OZwq1g0DnqAiZeocHP
hSA/Xke4ZgSRJYPYbHckUAVA8souGGls84qvPeWOqIvH2a/eeHkw4rzxHI2M8Zpt
ANomWiD2Nu8KbQgzkzOv3g==
`protect END_PROTECTED
