`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yK8jm5rET17MvzNbBDRlDj+qNn2JB0HhQ5eXEoS0V8XLZLK7YRsaJTk1a/v5DUOq
dgOWeMJ8JDi2BE6vpimW2UOfl/niExwzInyuj5Bg+hLD550y5zh3FN+OR2Sy5YzF
BdPtUTw0BoibpKiBTJhqAc3bZ3+XgkbFGoPhAvjk23WnqrRFYSDr7I6yy8+Gtm1K
0asDF9IiE6fRa3z46LOocc3ny7AgHO0QeO3JulcxlQgOW05pxBXORPrDcrJAGZxI
ghJPt3RzGatVfqXMoOa0uxfwM5JmersP0W91+ie92eq9+mYzaU+1Bsw8IlKUIVXT
EnKlhcAdErdVAegqrC78WviPAVFH3GFSio1t1S6VE8o/goKbXCS87hWMqP3M70cg
7B+m2rdO3JXcSnx8d9yBi3wQZBebMdbF2cod5CZDxF4=
`protect END_PROTECTED
