`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ol5IXwWJEeofvUOfJsVBaZNi4OeQTn2D7Xdz0itFTnSeVmhSHXcVGc+LsymWEo9D
Y4Zgv4J9EogLrEChDQIR5ItKL1p6VU8aL5nEW9J/gdoPeX/LKfkqylVteRoz2tl0
rKwDX7hzo/6ypJwBW27SjIK6qGGsRD4lhIf3WGtbaj9sfSYC+fLZDpwcvyfyhkUN
faO35OWdQ+OvhAlu1y/RY9wsvngOnTDn1EXbaM1gzTzjsx3nGtdtu41SnSZIzmvH
57qAl6Zcepz1GazYD1f36dxleyTu2A32b+QBkP5eGNocrDq2tAQ9yJqNkG2FQxM7
RiFzcJz3qmNIJvhwY0oXnsIK/vgwtpxe1eSu+E/MW76n24qe1N4bIG7aWqW0yWlp
1fTzvpN1hJTHQNk4CBaHyGsP6XC8o/5sFPUVxXVaGwcdRJR3zZyZ+sJnTXIVpisE
g5AXeHyKrNAqL63MyaJcap59H2MClhCNjgxMEONuJ+rcXVx7yrNQGoIwYxDquQIf
lz+Bp/kA5JD07yYZnG8wTP6eg2xQnPuriJEWF7BM+SRrULEO2xkPl7dUkG6FIJcB
ATDDY6Zeun+hzISxulUsgcWK+URCbAPUu17nKVBch76PusrVDOYAAVb/EmOFOBgx
+s9IZanyYeZbuz3bYQ30yt9Rv0k7BmbPmnW1l32Dq+iu/gGD/wbGpxnZZwrcJ8Rh
6rpyAvkmrt/+iaFaqTm5PTq/ER8h/NFitQWE60EVKfdsr/jCja713CPmZ8qNyz+8
+YjojOo+TFyCzslXW61y1kCRbTgZiAvMTWxq78hToR8MKawy9ZzRn6V6XwSJGNmG
gXSI7dNwjQTzJDcEFXrum8pZ187QjFHXsx9c3BR+VbmkesMHIoxRdygwpyoIZlUE
K3DleWqB3jYMul2UYTvo3SL7lFborXIyUgyRi4w87AgXii9ndl7zTR7d+AtxCJ7T
q4q3seD1VwkXqCLZtEzWLqCoWQezjqTICvs13h/4xye+Xur/umoZdP4fk5B1AZUa
effbfG9kOxeR6n//pFuNEvN4HZ1NpX87MbpMhby3oNSoxPJAgkg98Lg8hj7FYwao
ABLqa1WpLqz9IT9Y5KlJlyddix/nXfEj0noRmv0Z9crAvusIA04w428gfTbqz7cF
4Ifc+E03/BGV818oDn8Z6K5vfTR65bxX6HTKMkrb/t1khn4vgG4H9gKfzBGG39M6
rAwcvhRl4fCLqSNRtjFnK/719fUlRtjkdsvomyekhXK2hRhZLz/gKbRD02aLy4OP
`protect END_PROTECTED
