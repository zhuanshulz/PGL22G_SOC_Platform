`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wE5wGdqOBY7oeC3WMo/M11fC+o0o4/bfjjtSrdkVp2zyCBP08FKoknAwyquBlm5H
wsaaWpQC2aM5Ac6kC9NDMZODORUFHQYnCzyhm/XGwmlbpXbiF9xhutCNszfAIGzS
ao/rEe5jyQeTngD/Veb1+b7TB1ywUYcyni5r1u3by7I1nXzWYRLtAEQJuKJ6vUjO
F+HC2MGhqZebwKa2XSIdZ4VWz7gUaC8mRdMEUi8opt2yl7V8Fy6YpKXuYbdA+t5Y
tN5gYq6SvWu7vXRAcDS+t0lIrXOcDItnyajpnhlGzhsS8ZKGiHt0O2wZHedfJt56
vy/wEU6IuzuPkiCdDRtr09T+TgoEFNDLIznZY2jXDgzWu8H29GmqcURORxT0Cv9L
q/9rrdEjXoaHtbl+83l58sO+81JVGiauyfTs22lp6NH1nT2DjvBZ7F79WNdXChFg
ilzr5jED9IPQpDXu4ulThQ==
`protect END_PROTECTED
