`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L8jKe4vqDgaK5dItnwbJZXNLtFeyF6dC2FF4ZB/wHJ1LBKvNrv6xdo+aNT5A9nPd
2JefAQ4gxuaEQD4rkRFAT4JkISUsRdqTeC9qYPuQG0DWZ76BP5l/jRaP+c3jJcGl
Os6i0QIu8rZeCuwhL8sCAcdT6B2x4cQ+HBqs1zAI9bdWbj10lDAXGB9JNXJWQkSL
17e4BtO9m4Vqa+N121rQW9RoIbGSaFjgr+ReyChBCA9wnUm8Ih2XP4Mb2ickOhrx
9P/ZkKEMGuWhvXW1Rsu/2sXUDkQ10kk5eRO0pgacPgotv/ISjiCfZ7hAG8MhQlwI
Q9q3qltnociEcp90qao/NqdEhX/I0j5urvK77FrkS1/nErUMoZNxEg2HQjM1yV1G
8jtXm4FsAHIn8akdSsLUlYN+yWNfOtqeAQF1dkgd2bqgp5Qz9ODmJSiCOH0f17jj
9g5/eAJYkWutS/pNQBDpMY7FCVIq6AQWlh5zCZ1JlMtWQstTmsqCMiNOMCAQ8vSh
sygcVPAzE82vGDFPenv5jw==
`protect END_PROTECTED
