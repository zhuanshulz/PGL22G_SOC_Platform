`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Nw59KaAAWf/kbXaTJewnh79fE5eMkw1HU7GdWMCx0/EFdkryRYPQcnT20Mor/HXR
Y6kRMEneWpHUlimE5RApU0JFO1EIvxnHbxVGhQyf5SsnlNEY7q3R6qFDH6P/v1Al
e9vL5aNTxXiPeNmNrZ8Q8+evq+PGDAg3eOtTqSRgZCjw/WRjjier0xWoASCLGZMW
YH/ueTbVyGZkGmxZ7zQegXZPkf0sGhLu9n8dVVarUQ5uP5eH+lbJSSMQFqyvAbo+
xStNEGq07HfjVCTYHB5B0w0uBcn1Dw4FqMgoIsScLwNCcXgxpgRBD41iUn4t5dwB
53aZfvoUDdD6p9IXyDDq5W6jPBimHU47gladiZoXJrA840vt/7B+cR5IT7aweBdJ
ivCvMSXaTfvH5eQ/w/cgXnscMHWLO57dy5RQG4IzVPNdIRQevQYSFCMHZwLugPv4
AboT+FUfCiBiDhqa5VEhnvKZtHRcIEHefuYwI4wyoU6ip9rrW+WBEd7N/eK6KqDD
/BCGvXg919YsL9Fj+hU296377uXMsfXsYPoMAYWUhtjToMT3MEr5aw8p3ZeSe8vy
vxXCtQC2sJYPwnwMNA8ipQ==
`protect END_PROTECTED
