`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ArmCQ8kBPIZp0EOSZBO5m33W5/Fo8vCB+KyS6j2GZlQNwVL0pa4jHTxF9nxsb6Qk
/dvfoKVLo9cr+3qw5vR3PwG18BzhzLgXRJ97iZoBfBAukSALmH8aLOthc9PJKbzF
l6HXR+cM68TlH9mAZgP3j0OgfCQYyQ6n+NOvxTYC/hf8CjYgO7Ee7zRlrQmK+tUr
uCHu7mzd7FsQnHJwdaL0hMUra3LqUnTCzinAqThVRqVHFj50ve+k86HBjyzQotHB
f0RUL3/hCiLYzQ9KfT9MXWfdkY/XlsP5sdzaOiaAafS9W+lC52tF/ptSU6Nbfq5+
hIWcZGybivmeqTj/vYOKhAXvypy+qqnzaxAvbLalSyBLi/+NuvOpRx/YkPDKdHxh
9VNst7u/CkHihmMFTKA6cTvM6nspf/f9SuDfIz8VBEj2fLKalXC3JdrZmlo3siSo
JC6mRZOlGqhq+dwz6Q33gNkapZr15YcCqwfJEQ7j7tra604WU/Ev0Xrv/QKVLngh
Y5aYmCnAMV65GBJe4q2omKFX6ma2P/Yn9t+ORqahVlNG3EepLYgUotBudmv+k7ur
94AuLN/C0coLMXha06H2Uw==
`protect END_PROTECTED
