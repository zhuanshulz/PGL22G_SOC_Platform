`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F2G8AeIMyowUq4Kh/DRix35Xl9EnC82wch/aSoB1h40E+3azsqknEFhwAfTIJsd7
CQZGOpBammHgJNfb1fJO2QGYnTg2Kyhy2zErh1GCZrmKG2vdypJZjZYV1O9seou3
p0kgxGB56JGg6u/f2G87lSJMxGfdbEn6Ci75++DVaqCmfnvKalfLTUO5PDDddb4g
cRtUFbu9nrS8+mQ9ZKMxUZMmg5Vo2F3TsENs5Bd7scGRdzHT3b3PLB+cNqKSGn1r
bm2Cw+3CiXeiZ8NERLYEhJceNnLhYV2mfmN+V0u2ArhZ+Cr/CaVFjk2wxPRUdwT6
iWHyNQ6QWx3oDT0T44sieTpMMxuwaQgPC/IgN5qmVFxPntvuS6xExAd20WeawG98
hAR8h1kKyj2GPPoVrlAR8sIs4XiEWshAd9f49hwomjUdh48mTciFjv3qJFHmIxYs
RqXUF7l6kT+Mo7v8mWDr6h1lK+XdKDras37AtGgSHPL+SaZ1XBYH3MNVgGfGFZLZ
xt3+DR07S3dh7ZzBNJg0xMgGr2kZ560LUcFVgiEH4EWIqXvogxs2VP/0uhx1D/Bw
f7EJ3wxLo0t7+szrPSC811r9Rux1DTnGiDcJcHoBqfa9E+1iFxgTqM41QrCT83rm
APc8+bvxJA9Q+dyFEiYz9EAAIbGLLZwdd9R3USrJXl3ZEfDdqfbz45F0+FV0Iu1r
8vtCOexsi6LZdL/quoE+Acl6cj7U5FRDBtWX8J71aiA7/pS3lVcIT+AR0FhDfzq8
yqpSU8NLTWV9EpKx0Is5dbuBMaKksyNgh17WJQF9yFOkHfN62R+dCDYROUtuUfdc
FxsfEWmYDyBIQ5FuLwtP1Lo6Ni0nwxL3E4P4e36GU6FcBMvFVdTt19ob2dnjbVPK
NHVsRttlkqIDC/2pSpB0jnzO13i1ZxDB/iwhM0RS2H/tVlxRKd1IUn4fNJURJBbl
X3jXJ+KdEf+E5lE2VLjB8NRGjCnsTc4kXqtQgKJ0iHTQ8ZAgNHM67CawUaPTXYlH
SJrPNTIHTXGu8KSaDr0wgO4+cgnUV5Lmiqv6wnPBtcxv+wIOEFlAPu72ovgS6lzl
ro86Esda3zBKUoVXYPAadqC7GRHUoDt++fXYRuxpai+jJ5lRedHMSHf+pMeuU5nM
N7gCyHRNZXtvbfYrgiR+xGQq4aoj8ro0Hh5g84ePPrujb6EEkGjLDOtN9pD2rlnf
27xQ8Pee46fpiru19BrlWlWIJAOQpaWz1DbzQlLzBoFWhLs3yPVDRcLFSuXykoBe
UNQtOnGtZdl1Xo5pSX1E9AzKXF9g9rOAaJrJZn7TGqMLIFnwHySMQJQuNINOM2Pn
ffx/+rJ8J/iaptrYA0vAimGln9otGwRBzF1La866xrkANRTmgHflchN7jVz9siMb
GV5q53hA3YVko3SJaIlGoqdipgZlSoEvc3BDacPbdB+7w+XjA85y62qrtCJHy53/
SAlwoaSePYnRjt7aWv/rTJ1X5/sYRNgelSHqKTMtPI3tDaeSffTfxLSwH8RAbciq
SiPs252t3gd0q2iP82VNCGLhXwR6rHb48/b6+irrS1QmejZigiiLzPSZyTW0ngMK
YMWR5FLE6/mscJXH5//IZioVPKYH1r5cqNsCHryYNZv60zy/kdi3QmldNoN9MSlo
2qycmucY8wlwq1NtSiVA6GwC4tZbx6p352va0Gyjt6op2lqPpl3dLxuWuf7CzZtS
S8wGCwVM6IJ353vKe5zdK3ooC0nobzY75GEcU+3RvFsFZ4ZbHMkgempiT/nc3wiq
PaA8DCh/o03KRdq4H7eE9IHCEyhidmD/mYuQLfVBVc5o+54VHoUmKessTYy7M0O9
1ixJqtEdy9ZXXDvcK7E9rB8/fvvdpJw6MDAI/4BXye9p1kjmrxqoRD9xFLxWZc6k
UKFrSp1V67+/Ps+91Xf6T0SFhojJz5VwsPvRqZ/zsskhioKfikINvLE1tkF6kSWr
b/945pZsdBSNRTQPrcYHc9qxVkpdR1qMww89tT4M45qm50eRfqOq2vJFfM04Rvwm
dlw4yb5zJShKBFTKqQqd2vAopqB1uNM8INq0/xcB5Ka23WzQq+W8Eqe5acUA/zrE
ebeJ/eJzSuxE6p9NEkx3mBDREGS5DUx53xcCVBf1xMIR5UCvJ7+8hMD6NR6zuiFZ
NcrNGHPvjmGo+h5kA+Qwg+jDy+gy7P+GfukgnqlQSvi0lrev6e5zShXLWBdWurAp
BkNG1BxwiuibRDSfSwKTXRXVEdsELyrvwgV2ExtPn4WOsTWR0dpba6LRhCsXO2mj
puJp5bErE0K3kMt+9SwYbsJgAqmDSZ4IY7mkH3LT2wzg0PXehuZL02I9nO8ose2L
ppJVbLiPndT4mh8sgMqxg+qNlg7Wh9LqQSiVgkoZpc4pw1O68xOe+mVe1XlE6nCe
MVBfrc4E5aoU4NBcOy4eP7AdbXLqUdNmOJY6UAG8T9TA3Xro8hioWc+SfD7tvpi1
GjKi3tHst+UffYrbQRrsqOtNZAgeExbIg6eUNJlquzh7Emyhkpp7plxJGfj7lL0P
dkN9Aebcy1Fd5YkyXDmbV9YwEYJr7morQ+cu90ex1CQiJZca8RNJLpb0g9EXwjkY
I9W3wK4PD/ex5RM0o3iGkv8sAH47oxKrf/8f+UQdLn5jYS1yWohIF1mfaxc6AjDk
Vz7uMxFkskyJnjzYe40Va/92BjLd9B5EVACdi1AWsnciBfUzbxxi/og4+kQjulRL
BkRF2iVpMIoxHgutB5fB/voNHuyAWeAiiyw1ZeJqaUIBpzuXF6JZGpwu8lzGDRMw
qehRtGcgvAH/usvTzKveulhLQSiraPJ/ZSF8WI+7GhpvmXyCOav545N4xQkZF9VN
j+8n+CbsP63+DP1ij3Q+31mAbY7zkGaNUmVAX+uFi3j5NSh6b0CIgJfYtaeCkivM
TgXKyLKogwX9vfuXgT3WhPbSkgeEqj/82tBAQKOMJedy1dlSftkpvBzTXmBQ6gkn
+b/ElUyFrXE1Uhfs7adhnDzRjTWbY+jiyIbEYpBH/78noHwg59IFJy31zfcxKyAA
QFpxH8/AW6KfDt+Z8X86tGGXC0rw2VhojaRjvhEtoJXcdo6uz47iecBARH9QgVdk
QHncelRMdv2QrZZw+lu1y9oExMsQ/zbob95NXCsiTUGN9jt5o/SekyZGAa1ouL1r
yYQqOZvgyLoRpH0uU6Y8lFVz5xe/ao/WOZvuUCzn0pC9EiiS+w82PDSVliJSCd6J
w/A88JP1pvrz1TxqOSsOe38fkSyHHb14psD30FYObDnHfBCSUWqUGb3HUIbdfu9e
ZrX9t4jw6P6+5hDRBONxTw0/fkSnfS3VWvDpqbYdPwnJ9hZNoBAgznt3vbVezPNr
TQ9qwCVET9/itgTCpKFwvmzssriU3X7MT+YH9m4lsZuYpgZ3pNC82NsRzH7m0gdM
/vZNV2bbMTyv8o4IQIeTmWFb/9+Ayp5raNwlw+tf/Iv64RkC2U88eQ73xnq9o7eI
d+37h5Eru9K3bUpzB8Rr7bS21cdhk4XlseceWr3AVHkCd1U8mTbNklyLCpCYXLUj
74JE9jA5PMO2HQgN7GpxMleHYR0/tAGYxSEfjTkspsDpaPuUxb8TbgQ0kctZGvPl
e+3l5oy3p+n8HyxsTczeuwIt6VuulLms3TVfSlBW0CDksmUmbbUkm293k98sGvPH
aZ76HXyRjCmBkoTAG4NG89Gj1BoD/CvoJI8iszuP2QiCvq0NykmcJ6yCoYaKP2Yb
JtSSb3J0Ptti5rqc2WVxqI/9dEKpoEI0FRhQqYwEMPuwYNXvzfgnbTcMle/fQcAq
k/NOEsYJKrUN0LNLGwANUnGjabi4PSpQT0G4AsN3eXfYxA9F7wzKQV2CxdYJb0cH
fZ51tF4vSPbcc/G2ewMVBzrnZre9+FGg1R5i5ysApdJx6JnVL8p7bybW92a9CjZO
FD/ONMXSl7OZrP4FvNFBgcRKqoomuX+lCS45ErTZ0UMbgUjyr5TwxzVWYQWtkRIk
zfjcnNJgYz5jPhm/A/uE6moGKV2c2oqFc2JcrQwgD5Wb+M4G+46RfBhjP++2mqCi
dStgeAKd0RPGbQtXWm+Dk1jRAK3fKeIiVJ5+SYdSMUJ+D3qu36MNTr7Lht86En9u
0sv3bn7sDY3Merv8E6eBvzgS/GfQm0SuMomICwQ261P6AYp2+IN/hdn5Ip9qseB3
Wic1kX51T1lpRpucMerPpfRp7iwnEIljNuqnvjYBwrks4eO7H5B31I7SvOBaSVXt
6kCRq9FDUaIgoDUhE8yFOxLeXCnS04EHDoEnP2VsEs76znOFbxG9+qFD2WOsVs1e
JhLZUrrVb0YFKk99lleHITUnGymeSRgl+zzW6Ow6VravKJ4JWDT8iGFo914WGyc7
1CyCrd1kRfeiI+O1JuqKZvdAwn0XpJk1jvfAPHFo0eTKYMZl4QZbHQUzM5+NBFB5
57dvU5YvWj888+nCJPneM2Bpx9o4+6D7qRFKm8qDyJ2ptqJOQlG/a7fuqDJph1Hr
XrJkKJh7vxgANsGnxIdIdTvt9ypWi/vzytKvWwQvUGq4Quqa8qW9nGbIFgG+zAQC
O4OzgZXxlhaIWnIcX4/C2stlHXE17HeGAYDcQmn4le2daDieGTtTC0XA4Dl7oRNJ
sIFGM/JM6N1wgFQLNZEltLWSG0vzffuGr+oBDb3njSlel5oU8lGXqIhs4yJ1ogNY
+y8ok8BH6o2V6Be/RzXoS2wjJtrXoz7v/EuMEjZtWU0GpCDlG5SCRGqUKVji3LB9
hBIji1zRtoq2uXNpoytHYO6wTrphtDzMoW499GA7UApHBBzzcg4lOF8UID053AWP
NfkKZpdDy7EUnWT3OaSuDor6+syXRTDLdYND1RcO+s70Sx8gd5X/OXuUICeCIKCO
j/yXV57E/nAC2vkCfgQSNUtc0RgAzFOIocAn0UgB7kA7VqwUKOiTUmGlb97Y+WCe
ktU+/Z8HUMHVb0JurEmFuR45eULuDmBLUvsg/LeIR4kE1trx2JZPEqdafvuDckds
7W6+gEZHyYVIwIyH0HStje7kTWtTgk5+MgJZSAEVBPbnIvE9U7P1IpTLHhD1ACYs
r04VhTCa3/pErm6vngtUpAfDWBofSAG4guPk4ZiRiThP6oN5j9zwPfEF/uD89UNd
4wvvThX/ILLHMuyhajHjaulRFoz8wXCHMkieDCtK6iQnMk9nEnmIPE6X3S6o59NX
E56/ATe9UhLij8kr7zSP3f62ENzCwUXyRz/qcD43K3XG9lIUZjXocV2wj6Gm+L7Z
RDzFDGubODt4WEvtQmrryLrZXqa+R6DZj9lHbZFF7PiEvYuf6TjK4KyiG7qx+VWQ
H5IuqGuUckNjGGlyctXPXhZT3yFCq2sE6lk6DE9oY9e2dmq7/s31N2lx5K5wZFwp
YI0AndkIrk0IJ6NKjtbSleAg5PHFnVyqPP3lZCuQX7lp5Xj5ROJBMnlE3UJm0c2x
XHsvfHRqoKxz8av/ZcQ/oPAvzA5eroIdbZlO5Sv8i1z7RHDvAX3S9KPY8qTP2rTz
VH9tXdg5JgT8D/qPbz/wSrHCy1VkXiu1P3W9IMaHJRSrtuCVdVCtM0YodbM612mS
Vdz4U1FcBBWoMs2GQVrhY/beZumiU/lQZecvIXO3unmKqb6Z9cthz2X0V7e++qLM
bS6LTSEhMJKlGtAaqlSv6IZYHY7YtVX22Qdz1NVbqEb7JX1/BAgTfDfl/iPHL290
VglSy0OoSzdSCGIKWEVogsxCqGcEnZj2g37gAtQVFmB1X3408L1b74MnVDOOdQpf
Po3dGlTJyzz3SfYzF0xEbsyoA1EF3h4Dq7aFoGhGfLb/g+E/X7zGfYInxan5/8bR
S/xNB8sqR2nQ/9cDgBIkB3ihmnnva4ScvlcRWtG0T7DMjUdutbkRX7wuTko3jnLF
y8RsJQbWudt6St+mpMARuK7FYyG6BOITwXpVw2axcye9m5J49nkIwg/kAFbiH8iw
XeD95sNGhRD5bT+5IHfQMvziV0CYKkaR7xFcIUIfudekj/E8ZW0LiL9iZSA/bLeo
SEAj0CIAFdwhlXYTqNPcX1ddiopHuuIwj0YF4VIjH/bz3Yqi3q0zZUW+p5B8qonc
`protect END_PROTECTED
