`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IcRGA5qL2IrI1fF6nLp2I5nDkThwX0DT/zA6vuM8j8+hkkCkHeFn7jtFGQWYoaZ2
rc83jas4fdI3G/mu1x8sOjQ04IB5rozneU/a9r49CRjnwUPx6HR1HNMl7V34Nvo8
yEPwkkr327CrIa1v4FOJycYIFHj1E1jHugNulTFZbUMX+Fh5ZbwMLd45q3q3W4CV
UG1XxWPautDaoeXZZIlzViaJOfezkh4JLvyjfGKvRiypl1Wr8AyT6LnQY4zsApJj
XdsAh4HunqHE1fDRWqAKcA==
`protect END_PROTECTED
