`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
peAGXsJ9kkdkg/V/fU72xE5OhYl4x6ioIH/cn3T+jk86EMcHPOZpl/Nb7Z1HknOs
KTopOCUVz/LvrXtex/U6rTLOxAV/u42LQAlJN29dElA6Uw3EfQFZ20hzrRLtof6+
IVUrVUTn0BO5yM1u5PN8KboeoSuVqmNsV1ods6ZVq540yBLu0lsOfxo00XLocw3g
LMYqI+RzaN750vHKZeIk9AlEDMsetFBUXYavYZXfeJNWRW0++9J1ssxRGMIYYeOa
19fR3ick6KX0JbbF2mRTKB4eKCXivG8fykEqVwTs/s/ToWr4EaTuFK8Wt9U22yYf
KDL5DEwDteCuBENNmX1yjQ87/BXq6sbxSQD6dG7eHnD4cltsVlYLfT2U5/wciP6M
k3q1tlFGLSDpYQ2IhB4Mrv9ym5yCDx73EnBhSrdMKgp7t51yBZiAqAtiUHcULdk3
CANAevj44F/LLrDC+SvBQCu6kbs7lo1yV7wvWRNDKzrNm9khN2ZkF0I0c2XmKPcD
pFpzomFX+VGkAuE50u9U7D0RhHwDq0zHKifZgTkEC7rxykI5N0RS3aen2lJ06v67
Gjug84IGpniDXwKv1PL0mNUsYKyMlioOO2Kc60IXWTfI4QL+NZGvub7V6c67cSNc
fSYeMbGfokPB8Qn5VRPPrqwZd1QvC4vTp+KhJ41f55AXckY2HVjZKtvsrMLNnJH7
uzuPZIU4guJswzXxw1B9gQYJhHl8zVT0F3FOtlo8riWuHmqmlOASBFC9WuXxMQs7
ABL7N6zUhL7kDv2DayPyMo+sqAXREU8g36T99RoGasW4td2xXGZ308k72+VZwvqM
1+tFlVBGiGrVg7cNUAQT2oog7a5p+295faUaAZBPwOtDSLUQN5Jr+vTfCiLjVGWL
thzY2czp0N9NJEO4hLQf3+HeAj+niF5AYI/VIOnPfHMqV0H2A0Az2Afm0mvYtIAw
M/UmS1pPSqLWLjISPGHdMq1tD4wZEo/74NPKGufEtuOeUOfXhhdhxCAC1AcFG9z2
FFNUYXO9qe/XLursQNeI9jARwg+HooTmZM+AjuJaVH1G/Ghf+VjOZlPRzemHTRjr
hGtZ+qIhbYNNeQ+rs8vynGi+tvfyGVWArrRpNNhVRpfvlBjIigDRAc/NHop5oPhr
gSXLPTD+Qz6cBUwSVDoqL239iNYvblCvt4AX8JbpSlfFUc6F4mvMKc3nYL4iI+dk
U7L63CHtFrCS5X07lr3ybjMbjxtqOApos+RJhDmSIpT+s5ckQF69qRI2UddRjmUr
iGUCC6elUQ8Swl/7/HOgTUL4rYkZt6pvhfX1ty7FEJFxG3pBnVM1CghRyBxlNeNJ
oYaNOl6VKslBwad4kngqnt1HFYi0JailxTTN8slNm8+oUJ5k6UPLPzNq9OGhm7H0
SfML3C+bW9N/8oCJxzjoVZYP9UiXMl3jEKFuKcXUtacZmKKyf9wLQwtA12K3NShZ
/9vs920UYAehWvof0+kv/xCj/kWSBcNiSFEOIQgYjhX8HU81g+2D43ncE+1JKrqk
wqhv0e8JB3+c1CmgtyU0C5JeMtf5tH+NsSbswF5RUYm7q0OiEQ3U4ZjUChuu5Tll
fKYomqznkieKBIgG6XC/rJhpIqLWGKPvFW9u51F4KYBfZimjgOroa/JgAdLpRbxI
2956Shq9KU7B8lV6/htHser6mG0NKoRIP6yC2PHktK/jLB3FPf588VQzCriySc/j
IuBQbyaxjwV5KkPeN+dQ/mz+8tKt8VJQsMWgFvHV+oo4Abyev80ncMU2ZfZrzKAu
VlzDUdt3Su+ijWi7d87IJrZEU6nKlB5OzRk0zd2QjkEoU7ywh/EG5tk8Vrkf6alZ
6veLEP45JV0Bb06xEUVOc4NWJlD/rFQK6FzpWMydSdXkwMUXIKKgrDcYaXIVLu2y
aDnkgOpHGB7tTa626kBbNUxrf+IaANlND8zmVVnG57M25EXIXlnIk9YgvstJvBj2
Gvrdt48Etf/4U2ys8XYw7sT2D3cmHbK8eIvu5ESG2uEkOUZV853gb3jlvUQrwAiZ
ju5PwruWNwUhpe1a2QcBY5uB3YOHadjJAQb8niyRoq0t/AyqJP1JSDI07Hm1eCd9
K61ueyMBjAOjfJVtA/cuKoredgYezVXeWhY1dn5UPS76VmsWnw6wSdsOGAJrSyw4
ZdhXHI0bFaNPMLD0zfo6CGd6gU5kkzCW1AyJemZu9df6nPork3BBodLzezIgCvz/
Sub9bcUczRtibJO0hONdvD+r3eT5420BqRHMUe04XrCi8pzos6Ci0fvWgj6Hx4Od
YLFMPf7MTD1UALcjU9Kselfkj8KZe3hgmdUI2OtLwcQ3kCZxTdcQMhqEIplk6YAO
dCGCjhBn0B2oQ1mRVQ12+W7cMUDI1AQ/exVjFncEetc5d1BlblinWPtacBw5fg7I
pqIhFsPG3PdZimwJ391oO7KPM7WJcfWr0dg7v6XGwf5Up/1ZPAycnWlrykNB4Shb
XC8PGO3Pj8isCcnr26tO5fGDp9WJo2TjwiSknAs0u89PWgx5O4QkBf+uo7qkulGW
L8/JuH4F7YyBCC0d98Iq8BsPzaTDDShoq4IpTcvmDw3kfDZzI+691Rd3TDpgRddn
fJopWU705eApPE5umqymvtO3r5Rkps3QKCl6RaajQqAolf70dg4EjQv6ieBZb+AK
FRd/TXeGdlMaQdqHlhzzLthm7dbJsy3l76+AGEsv52zkdAkew9zQnu9bxWQKwJoW
Z38ub1rBjRfRDCEpp2vXJfJzysIAKk7zQX/gvqC905vnI7GUjyKRZdGd4b0OB2e5
+l3extKE0+y2onnClx0g3elfv+ra0Ih4QQG7khunEGwr3As5vU/SwM6Cr8J60b/W
LBJ1BUswqS+C07vSiGQYpDIYgY71PIENpWHaxIn1lrYf4k0tzIohRhzw3lWEPRyJ
3FvwxiqJNKqcwsKdpittrz6gKnpS4C1D1WHXYmpUPCWPHPRJzUOhESVnZmM8JcCH
JbPFl7C/D7bg7kSkSdsSOW56iH9/aQG3ihw1X+4iX1PPLv7xeDo380jBCIk0frSO
gp4tZDL8C3FAYO4oY1Wv6cUMrnxDzfCCEk1GTKlZ+S2xZHgzm0yN6Oyzn+514Fi/
By1w7QKhu9Z4L+Ax9yTDhfbV4zAn/r2FhLSyJv01lGSJ9R4K5hwfNuiOh69XDcXu
QdLWV5nElyDGE4zMHSGgkhBvBjvuIhuS6YAul1aKCPI2oxK9z0ELACeImdd11440
P5UweWQgYzwAqf4P54s5ZB3ETNfJzn0CiOmZMIgoZJeIAkDOP1OyzV5QARiyIGlo
jKVPsbubS7k7//qc31sewIMRVGJm9X0ocGJjH8xRAd0pQ2rVv2KzK3n3l7gy62Rn
4i8//JP3G2uUzkUddldgIc3RetVECrcP8Z54W08Y3TnWnIqtdQfoqwY+DjPoPVFM
ILdusv4q/Cx2OmM9PW/w95jQFdbQU8HBjtV7UjTJCjvUxTV43mhcoxplg52A3cWQ
HLuD9Mj8AvVeYkL68c2lLkXX6JE3AFckBpjSC5pWCwMuo5/PQtSE0oOjsgHfsaOe
Qm+KU+9MCfPODj8vnAXadpFFPtdAZX9iQBGhyhVlCh4a8TEpbpxujb9z0otJZu0T
2yYZ6DGC41MdeW2A/rb+ad1YU9DVpuPCDTc7k/hhTlVCS4V7tAR3SQjQ+p4e5kQH
f6W26KIwJqmBupRxb+CSFJqK7TCLWNjZGA76EVz8F1hc3KYEobLOhFOdeLVFJgUg
Vuhe1Rnk5ZLghVUoIVQQtFexGjadGc1QZzMchddD/Tw0V5Tl4IeWsPHjANC9iYrv
gDw0I7kjAqV5LLJvnRqM1fcusJKPeB/GLdC5Cm2cTd32Facrp5zU6udF2GvQrbXJ
GSZImgH7U6Uf1LZCfcbeQgnNAXCYYIle2rCdaRtL0BeohcGPW1VedGwllvJ4FbRC
ERHUwUgp/GBpOUVHjwKQPOADnazEx87pZXNAmvkIGoCQ0lsQ4qRkeWTm5b77Hc8k
x0iyGm541H2w2cZj2S3yq9r7dR9FOc1AvKvtXP434wQKU4lq9ABgbpeqhehCwf4E
YD6Tz8KE068RXjrHXg0+I3lm5KcUIwKoa/x1f0940/vvRRnVyhyje6JBEUPheGVR
tlGMS2F4omNkeMIr8fO1hNifMTBz2hSdck2bRg7XnDzC/vuRZ0IkaTHFGrtu/lvR
buzJe0wHW716VpS7+lbcVPNaeZUEG5fAm/57u36uHqAcplcU6E1zlUB8fcYYWZta
pGgZKnaFwKb2FZTGJ74aPhdWxIqDFf4by9suPTjd5UjYrg0jxDPhZiUrT0B3D6L3
hnrNozX2JHrvsNWnlzjlkhAMCAl2Dw5fjkA9+G/ClYorH5TQovhjfp11eiLuVUS0
ZWVUnkORtmVAX5qhhQczh2a3Tobud/3CJaFOCTNQT4CgyINKajEfYbhieC4ix+kF
/FNFHzsL7zPgC9+1LR/O5wIb7D71kd9LuYNaCuaxwb1ehPMVizr7KTbMs/ihirGh
bJ6RhKOqY1l3zGtvpR8T9vMJv9hFQRG1m8kZsBkaUlkl9wJoo/nfqx+bByQlNlgX
y74mpZ5B/Q93i80QyfrgpiDE7KuVmc47qWmBA5uAO0AjPiI4XGgS/J26DJuJ4ESl
2TM25tA547+PzlOye8U6DKOQQqJZSZuUKhJ/4ji7Wy6mqNJ1lYafWDmosomxlGwO
Cna8KyDlYeQC/jcE6Wz+FDkb6sgXe79bs/D83aejfXfAWt8/N2Ni+fVfjn24QcjI
cnNusGaCYn5EgCsEe/+tbMbEmiRruvy0yBsHZ33ENrPwFk67yt8NC8NzyIslbTnM
POYhEeYLzvGeVezcbDD1Y6Gijt5IdgZ/5x84Z3oqp4FC6Za61sAgfGbN/8BkSzhq
eRE7oxEQBJSrZGp1ANiygIY+3LCFxAwvacKzlmD+mpzZsAz0CJrhUb7azuSQ5vwR
C3E2oz2Q+GiiayjMra7fHXKOQK+nqC8exBdmwwK2pPTC6a5xVNEoltb+W2B+RIHK
9XAFdlQ8D5Ozo+9K65mfbiSgMghhU4zRYjuTn7PwPCoR1H0AjTIxkOHi+oaGE7Eq
lTe4OE08jTiVYgmFyXZTDaUFvosl+C15Ryqjwhyge8Xr9J8BWSUiRtf1TPm2ciji
GpMl1Hut2dXXoObsaBo0gV5DiU/G4s4yXvVZ4uEE7DT9OWPu85au0j6EWZAbnkxK
98nj7kv4KYC++uSuvDL5gvuQH8v0Mrfa0hTPPdQULXkdpoqf7dGfCrO3vG7PszKt
2nPIuAO6Qart85Tib37CCYYCqi6F1EUuMoX0/lipnGnywSd/KGFSDIJitgSEusC0
FA1HRIhE74lg18JLIenePu0RjRfUqCFakrJczCZ4Yy3fhoyqrbS0RO7VEt1gW6Kx
UbIp5tFOw8kCvcuh7tLn9NSfefcw0nIHSRrYzBpwRlkV/h0OOqf6AIhbnNjyDkoD
voBs4y6HacAbX3DhWUxvt+/TV492+7G095e6yyUrCtRiGywOLQkZlozshT45C0yA
s5JexkNm/4zONDcv2TFC0ndHzIwWCw9loIiQ4m0t+MSSelLHyzU971LUvAni0fC9
OfZmCiJO/D8BpTVCX/2h6rHSN9kWt+70KdDJ+cqsGTiVFS7CLSHRRsbaPCZyXtES
G9IavdyMI1trii8Jg3bXi4aDQx/Xhx4Gp7WwP3EXt/MikIgBNS6DQ7BUDPDqQTM8
daz14s5nrl8ZOixZRKsiszC2dd5gTiRML81X2MiGMK/vUAVjDeL/cECKU8ln+hCQ
ZglZXySXer5pHZvtSD5SUSBP+40sYTxZb0T9ChfMRb8SamHednpDyzX0p/nFRJl0
cdlr2VRXM5VSLCFAgyDJsWW1eVtGFWpHBMZ/KhWgIPU1RLNafMxI72NpQ0NTy+Iq
YXn1x/UAn0uCW7u1Q9Zu9cOljKEs5IIl7aUk3loJCt0A16B7WAXWD1E42c8i4jiB
RPXecS2a57h9/RfKLM7QKNeFjoLXd1WPr+UA7xM0riXujps2n+rJzm7YHWn1/UB2
LsUXqQevw9K2ff/LdNNIv8XCDHrvpTM4wpQNTb4wvkIFuILeZRbTvozjJiJTUYQH
Zv6bb0SBhhHWD5MiNct6mZyLHH4LAkQIvuBk/4nK0jbsQR+cn5AmyvJYRww2nvGL
oSk6hTmu396g3uipPjMYj5/gcI70mPJvOA7HneJ8tX0bJH5Vxn2socCkbHqE89sW
MbZCCj3jIPnWlJOhDDpcmzVTV9sc8XL4nJ3RqGQ5pOVZdOO1duDS2DspZU1xxVY6
CQgXkenwCJ/TjhyySuKw1KiPHt26poSzVQ+cEP1YT9N5YhaNbeZ9c9lmqeE23Z3N
YLszcqgoNOsZoEi6MuLVDh2Skspmz4wWEE8AWJbVwuL+DdX3Y6CqRTnVjJMjXVVO
GAqv2xChW5bMhAug1JMq8/ps7qiq/QSrnLui1d+jDJHH+bCXNtU17OKaK8TuQu7T
Bdwi90dOz/1Pn+k8Nmne2g1tM7ry36F5kEQSdb0gNXYfXBDeBfR/UBfMysavXx8A
xwOTfq2lxrTEcVkwrjoPi1GK5sHmyJ7JtFYcsnec2QMTvWj1n3DSk0Lttb7bLQ6P
PQaqSTVf4lJi52AlQta0XVIq7bTtJPGS41mxSccLKzH7Qo8WpUlY7RhX9KzEReom
ZXkKG77PaeW0ORuihjyApPbCI2t7cqcYkDTwX2pF2qQKKDJdRifcoNyEamuHSnfD
Q1Ezly2CEsaNmOid7sQjLZFAEKm1SftXRxZ8EhSFZj6PZNdT6rJKIwgXkAl/Kf9j
fNUHD/KyBieJ7C9EEbeiR7+LVjTRCIWBWyowJFb0RlslikXeS+cSQ45+MoYC3wnu
9cxIe+uAvXlpnmqVvZCsvOMdHpC5/2vMCw6hwbRjKOHpbjMnRJ32dFSpGTIxZbcc
JW7852sMx4eukOq9Bom+S3lRaCSH6UAmR7Fsjk93HTUwtlv+4eXkk9vPgBn916FN
2oa+vj4l836goW4J/KCk4ScNTDBO+cCrRdz6H8870JqEjJ+9/PQdEzhOmKYswx8G
X4j/UjcSAJGPGQ/ODFGd/Snp0iqS1/NDLvJ3EQrtFj2SZ9k5PcmcQaOou0izwIme
3ZNlgEX0WfBaCzswlIIcmbMifuCJYYTU5QvTJMjtVlwS7rIHQ/XsnNSnApC1Dr3y
ckzJNXuW5AHGgaNH1jM3LlzwNvdgtvTAkSdois2M3dfkiXXcPEJusNS2ubFSam6y
2WA2iAH4uEV7NCd1H2ZsWuBtcxzJVM9JM+Q1J848LJXao1sRF+dAXZ1lTSSdvZij
SU0vGphbhnHcKco36XbsaOgGg0Vcz9X5D0Ux7ymFtjSuCDuNGPfTJH6PfygNJZGO
PWEixxUZMZp5hqlGseTcabi6kCEuOUuugi78BbxJXudQvyJUY5csHc8aoEdrkBFr
+cD2iZ2DdxXkYbTJlf2XiAUKw2LKRO9CAUm5yTyNTNIxWT33L9FBEwZzNhxP+eCx
3tVkFqCm6jQZvQhhNSJ6vBuLVDS3MZU36EXHByeupXSiCjiM4fK5jVishK7xZPjg
BE/uyyBthBNldU8bV+cCMLrX9APIDYSYxSHwpXzLpF7gD83iIxlICaXsK8zB1STp
NQR8zFC6AkdksEiJ6PbNimRTpxYp++O4pFX3wly2PQLjuNshTa0X5d1c4dpnq8FS
0V3H3vRSY/hTuzrppU7Zhi6UQxPddalg9GdHc1Db8b1uZeIkiu4f2Va5PRzJbQc0
oLJEJcHORTJK7OU4DNsjRDa7PVg5pFvwow+IHxPh+Th06c+7sYcYlQGBWG4GkWI/
dDuAw+EE2SRZi4gEXaG6AhbQiQZvUh7QFR6+kjNIEarBRksA7pmzHh4ojAZZeC0Z
xlsqLpKrNEZNaxXw3xG2/S3CHg7cv93BJtogfxLdGPZkFa5q4DilwGGQXv2mCyz5
KuCgGA0ZHIcHX7lVDZ9cGNYOZTwgjavM0BYFSfJR9mu0hEHUDRqEEBqMszmFzVXR
4L+6BhWqm0LElhAs3LZr1wxld3rwaB4acQ2Aon2EygApqnlvcbza/U0Fr0hOvGLY
8mUB4hxwGHPCtrVkrOy56E8yIJRReLwKGrJPdGxxsrvm9Rh/xJQV1UfmBTudbLUV
SSu04k4aZ+WSxpexrJ5S4BHssB5C7czmHdZOdejFcCHFO3ALJMw5ztAAueBJyigP
Sy7mjGhoIyGHvw17AnyvvZEeSO8jUHj5ksaoOdmnjDUdrTo+BCp3C3KlF7MGmiIt
PM4Ez2kk2c7x57ad91Vl+I+DvaSXYApUfk8ybWzQo/N/xYxhCytV3hrJpW9PCe/8
F79FrdVASzLjHbou1Hs4A+ll7wrUb6blfLHP07aJDlJhXsBbPjmoESQ5ipQqGfTB
IigyNhyquQcXeA9oGpDK0qrX6ykiXJYTZp8IPpT3hvC3hVdTyjzSdK76orfqutx3
zyJ1QtCxnqy0bTfwPdcTxV2fpVK8dQEwuP0bTN2nSgKIsykTH9c9kxf+X1uNljDl
mjdan78pMGP7ruZVk2GN/bQ0imaSGNZ6/FVyjAyAFLUh1XkRywbltV31Jok/Dcgs
YyVfnc0p/JKc5lERQipR39Rg5p7c6G+be5dJB5IBZ5Y0E3fGtZcuJVEAos9xJkkW
ld2Oyd3Awkjw8bHXzK0T7ZDV94GACMOmHSFdzj6eYeD68V5xCLcZI4JIZdibhHiA
4hCzj+b/4pkuR2qDu4aRCTl5fK3oTXNUzKqRkpqblviJkRISD0uG4LaosANTptsm
VpOSVfsrM+xB0FjvvPZ+aJN+47dSpbc2eLfEj5sM9LdMUPZpCAq92nqu780MtVJ5
IZIhmiJjR4hmXiUcGJ9lZptidWB1nlNaiOaHdgr0323uGIB2aJWYMFD3sLK3ozBY
suxL6U+cmbRSn6paa7uIrJhEAQz11rFSHYV2H5mW0ueJnRhWCeB/Mr60q7DxKMg1
O32EQl+sTIU2gW8K0CFo+9o8CD3XSbXsb0kZ8Nq4q5TqqEAEoek+NVPwfM32NNdL
GvEjS4XMZyFE7SZj0BXYHlW8HAaijFhhzE/mIXUXJo4=
`protect END_PROTECTED
