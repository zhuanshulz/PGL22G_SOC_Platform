`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6jb/lZrKs6zGiFgE1qNaIdljp7NKxi8znbWW3OwnM/GmwDl5uA2azVelY94Tb2nX
9MRf8s+zSPl64V0qmzdFfheySseP76NGgj1jokqvFfIg4h6LupIJMFm2bwzD5iUu
aSaBYHhE4aIw660z1hTurr3xzZHwXE69iAT1zXquzTeObwGLtjAaD79U9VOuD5G4
9j2sn3QOieIAKw9iikOknu3NPwyxLXLYIsaoItUPMZS3c/FjbQmXvBH08bVsF9GE
jZ1o5DcMCiSRF97BJL4hEztpkXwDc+anAz7NRgMM9AkUSi5XNjL+ELoa0aluyUoZ
8Rwj4wRalLlpIU+DiqiwEhH9rbBKpg3Pd8eHYbO0O+7+zZbEi76FrNYQgaBFfb0j
lPJMz5TS2Gh27rjQcMXrdSpZ/sc+HdkDs4S6UxPsGMHEBCmpbiqNjdb48hLfSAOb
kuQgRoCQ8Jyr78jmHsum9RFJ+pbbp9Si5/TSYarCPV3TY8UGKOHopp7T5fasf+qf
NM54oGI9d5FyjsLrzkcnXayRuwMfSSb9jHASJMT4fs217FRyyTrjXeeAyqnwId/7
6mmDY2VTW+v05bR71Fo9F4+ib/7zCX6XdW5ZP5UMrDGp/JMNyvccRqYYUpGc1xK9
S7A0IPSWjOM4Wm3BroeFOJUSYoOv3bNZzZkABVvyqVYhqi7IWmyfn/qkxn/8TrZh
h/pfCKV/FIZMd3JYCQpN+qiK30ExeJGV9mwYNv7SOWFPI+3wT1XxdAAfXIzAxerP
xIBKKEuf/rL7Fc2OPyCl0rOAnqQ+CvUD/9U3L+HEVvi4iL1oycGwIi9ivZqiFRxl
zphotL6GnQYlohgAxx+rTWOnZKDUNL/GxhKg8bwTKQht1XnUElEmhapvxbn0QUjZ
D/kb/B7c6ePRNzJ9+egxNiOV8nRjLlsCGMj9D207L5ZbJ8OW6de12kdTSozqn+dX
6Wb2H0/R+0dW1kn1eMMhb9rI0quvHlfveExDJpW12428ZfYNhV8Y2zIph7Kf9z56
dEAE0bswKolxOnD12oUosv8JBqG/wrBwT5hqNRZvYNRpPLxIyRRKezddv+Bfq2xK
xH7FSlPfMvaEzOSJ/Hb2uA0p1FYRxNeLPbLSy5wwQqfLl2d6Bhl4BJg9gl/FgOzu
fvKRhpCcCnTK15YWdqO2DIf1imM2OhLZQkEgTwSznnaAYposn6f0h02xO6lyTJZS
0P63j70+bqc8vrladrALuq0IOy7cJBu/nFuMiXfzUUf79AyoddaUMOwuQwvDiWnV
Uo1TJgbkezopAFTJG0S0jnr+5MOGIxj3nsHxJ6Opjuqk3LJD880XE/asgnW7yqvQ
0AiRM30++pYfygCIuRzEQsGUgr1lZG52a46hn5bpbVMT722ZbxdzAVX0U2lN4Ddq
HFbzgjJO+Q1xon+6mRvG1UyyY/SRyUwBx17OgmL9iwciE2oItzpRRsc+5zXZX7J/
l+nQLT1R99BvOUgpE6WGbsOrbkoP69x2TBtewrBfdQskWLA5SwE8EZoysI/rF5e6
sE23DAqVOGFEdOoev0Qkjrlx//x8o0o4CfkECxVhKrkHVQw5tjZS10iqFa/a6LKu
hVMCKxzfhDtIm0SFRWN2vKGPrWBiP3/Udu6UB8WbjVq1N907XfrMa2nWV90Ktm1y
e8/m0clEKG623IVwlXSChnC7R3gL+4KrVK2FWGW/clyErApdJFu5mpOpP3aSG17D
qe96SLJShPhdwrr2GW1d0+5LQHB5dJzIGab4tXBVBOdGRB8o3cHvLAGrpJKpIsJX
jpEAfqdQVnHZSwz8tKAui6DVXHTgdptC8Ps9xhF8g8v16Rt/8xWIHL4Ka8Na+Xub
25vkKGd58eKb6e5AHLhfvLaSw9rtMWTH9aBVK1CmiuobmziyIci2Isi6af0JXaVC
qJst2jYxVIWr732z2XJA3qnktUcWllw8xVw8hucYIL8iOCnqwQWgHLdSZ+AZ54Mp
iQ4tYYEQQJWo4tcJX4OQX6p7TsibhSWH7o3LYOf7mto084acCZ7KpcWYrmcIfuNH
248mJRx8nXTVKzzZzdN0UaZ5z7DpF86/x4abguR1LH8CyV1BUY9OUPie5v3UYiB9
N92p4UyVXAokxKwbXGUaBiybVaDSsUoqPTvt4rmqguQn/2L4a0GCW9/kcQ/0+n8V
ydwtOlXj/9jJO8gpKEEorQWZ/+5VQek/HW7jpXubfuJE420Q6c8qFGFDO4wzp71x
AY1Lj4Ja+bzgwoNMNanD4Zys3hur2rR71bQdQ0rEWdYZ5T/TakSxmzixpARM+6E3
hqqTNTpwqlE3RSrfjJQ4/ewLWTpRyaQF1fZ7fKLyxCCOTbdfX3fNAJJIsyyj5eYl
W4oFmcd1uxpEqP4iLdhEY2GO9oSrk8w8UIjGNvuVXnKD+25IBJd5ld/wcF13bWls
TUR4IP+ZwXXR4XvnvXbMXdHX6nNk9weoYBkncXPSdQZ+Wj5LMnIWQP4B0RJxND9F
Z9OjebXHI5sFt1Gvdp3nkYAEh0NVQ9fFx4RIsZGhOdVfG5qmc7tpDtUDgt/RRnV1
+oFmMnR8jXMbGrjDeqbP5zLdeBL69N5terjbYFfPvf0l6TphKZnkLLMHIEO6SozU
8imQXWCwr3XfdF3b4VFwm2u3R7PpMfX5BnEln9T/+sK9uDVQDulW9yeTXifllVG5
P9Z5aRL2Wqecbht3PBSh4l9fjESba9wtkuiAmR43PmEYncChdDP4Ko0gSblGVcPx
B0XHlEUj9VPAfecT/+9gLwEay1sMts6azBlUAGx3GZ1DlwfEUhR59vo0djD8nREz
Tw6SlgRv9fqIqsd1XAz3geA0yUARJwTEsZUx5S45UX+v6FgZGzNUGw+4kpqaNGgI
UK2zPTahkzMi7OsNfgr+9yaTL/Ik+jnreD/LmE00s4laq31F6TZd0p1DcazQpF/h
zqgdUnrwktOYXjxIifE7K1whqJ87ji8mEzBAfVMDlf9pp3a7F2s8+DVyWRAsNwKP
nKe9zyfXozNz8vYJrFJp3agUYtvDMi/tF65WAYJwYeRenXA3YfLoVK5bF2dHcUIM
RXOpWJwB5Oz3PobbNsnPrkMq4tUsqHSME7oR0r3AXAy80MkkS1dh+rp+draLVLkj
BulcTRkqmxovaxKG6ShmL5uMSWz9GK9NP1UdirmD3yLtbAXEPW3GSALNBwO1xCOK
GrbYeOL8ejNmWa3P5C2U6eNvAOdk8hJbuY3v1WKovySJNj1l+ixZfiY/IcRXFYak
xFDt2518iNJ4H7XckGGkELGcVH4S1NtPbpxrLc7TahWW4adl9sCBF5IxUM7DmJZX
hPM9xDdl+T6TH+cxrJV1nhFSjOaQ104RYYTojGNFUFDczm6kM1SvnLnAmVDn1coK
rESJqv+gA6LHWGbUZ6LZPL+wSmNwnfBcfB3vF470jil9F9lxK6a8OaMApzxkYzgW
iFHSQlbWYzCTgtJXRy2bJmPldJ8bztOAE6UmmJlJZPpW3t4md+eQEOknpKmf3vKG
yWNR/4CTVgB8vNz8MGMouk6cCkBLC3KqLApl5ebfRK9FgbNiuBCg8+OM/uQnskaw
dh6jTR5zmahyApjQJV06UJnA1eBWZcEnHOhhfVlcqw7H/CNZanlm8YTj4djVbluN
Rw28pmLPPAmDnY4KyqQ0TxdFJI+Mcz8UH1p+FGEV558ojczZmA1fGkl2Y0Q423Lm
KM+wyXzgnqOpnC9+qINBOYOYBmwRG+rdYa8m2t29mivi6G4x9JOZc11Aj28lpoiO
fWOU1m0grv7MOVwFcVAHYfyhR0WYVKqV6lhhNcVD3ExZCt009hkwCdVLYChTATAv
iciUWnYionj3Q3j99okXYF2TbCZitcqRw2PJHA3wUxiXzlnnvrGVsIYlGsXKBWaA
StFCgzQ8GE8b1IYvMo4tXkWDlj7Zh0OFHudSEVlJAYiw68P101tMOlXqKqJiOdgI
iFNM+ozH3a26fpeTgEWRUewQazev8fwIbnJCVbQ2kb4rcWTqO+zMGoWDDZydxUln
RHsS1rT/3Utv/RZ+4Mq3JwMcarnUZ9v/y1EKI2SPqgQqrVo4sz/bN+6pD8AlyuXg
t8XcUMtkVr0AtFVnO5RGl6R5Hl7XcYbDgJ/LvmXb5R/AAHzaqRnCrz8dFwUw1HJD
4b4RPODClmp2xTfPz1xe5+3e3wDBlQeh4qF4XEwEPBPya/nJXJcAH7tKYKLiJDJh
5we3RHf1anT3ZQAVZJNsM1KLKkFBWNpZCxW54s5BdY0kaS8aLu/L7yMONSXpHfMK
ecTowfQx9fwT9Sx3sXaW6t2tNHutWdQM0/KCXLfIhQvXUXRJ6VnbXZbsMi+EsTaE
8EbHOxdx0OMc1YKlCxZvAilQfsQ4Yp+fhhAgsvQtGlzYdofrtwHoNXfmbq3cJ+ah
amu3z8dq/7zvlFOkXwIXyO9iWs9tTMUG2fvwxrKbTcncSiJjN7Atbxq6t3FGGw1i
CRzTubTiw/lmhr/tgteVpvPHTr1VsWjXWdAsAPSB4jg98y9AOfWIgRY3FoOK535T
oynSbHIYG9AzinvtKorK7Z/6OvFzk3Ynn6CJd9XaUJfCJbpezMd8gAMNPFROguSk
VTH62eFl2vEkm47KXnBb/SQeXE8tYvz72EwmDRyvs74=
`protect END_PROTECTED
