`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7Dqzi6guc5GdtoSra4tcKp0xx/PVCnWyy30M6oQLcK1Vg3aVgDv0j5sbpByXqWKz
AmeJZKiau+wQofTjRXsINnOTf7m3J3U+gIPKx/hkUAy1Q+6Xm6vATVDzJq+Oxdib
B6bO92RjVSlPjH/+BeMI+/RVFG0ykiLAv6OPOw26QC1kYmYHYaFcjEG6dV4IasEA
rU89pvMNv0oZausqq5U8aiTrkiVXqagb/Bg2gpXDLxROIvtd5KTt+CFkPkDsfqQ9
4Ti0WWZ40S3T7DRrStjEPJJrxxrBFlJW864Y1isYVLtQKqKWPcR/eiEdKEvPzWHC
1H9ciRh3GnqtktZrJi9YZ4Dn54WaxdTmm/TMwpSIzrzrBH756UFQmbZHwcDOsbS7
H2xiYKVU5JbJ2R6L8aRSaL5yX6xkKzBGLW68qnk4E/pb1LE7YaHsICovlOR507Nh
Ypagy6SFEGjoTLcrA3Mdlbjtke4Mf/Ei+VTkafQTvFc5xziQLTXwW8GSLbeSVPIi
aYIJ3IvLMiI7izreanPrYh23qk+vcLsgCv+S+NiH1KEze7Lcl3B85ssrX5ujO3Lj
JbDoBnHYZvlp7XsCj+IWQ6uc+c8YVi6lBf6tLoKsGjfETMYA3BoDz2PtszQxoygx
v8tsNYTJFqYAecQfozQE0htLr4gvOJC/gv3LY1M3tG/te33NqoCd0Ww8D8vWN43s
PgLSoyvjeiTs7p3s0You17GRRr/kpKDcANa5ldHbV6soqtFNrKriZvIQaaHzlNe/
Tjp8GwOj/Dl6qCkB3JrDu0COGs939Dmm3dVhizlerE3DktYbwBNfSjYrNmyC/e8c
SNFtYn4pVvvZALx4sJMAwqaRZyq9mJdJG8XoSCrf2tq1oxqMGIuRvEcy0hBv8MOa
CktdE8uUkc4AIqfzHxetYTdRqR48mrupmwAZsx+1IerTB0e5gXQCnF77cHMGU9tV
4gnHG6OZ6D6ZKOh+oVRgYm8kB1VrvWmRbUAyKl5BO1uiEkyPpZtiPyjESlTpxRFc
`protect END_PROTECTED
