`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2Qe9LMD+8BfJMTxJlnmsM8zk65sarN5wCLJKt1fVNaxPBQW0bb/DewvlDFYhwMux
7Hx9+4VInAKIhmzcaiMeyqgJlNYqVmiuhfG+uBu6CXyzb1ej1RQ/6mAXsRpzM31W
Om2ns20uwDx10T1dVMAy7ryl4xIj0PxEisZagjcy+jW/VnPb2FNfbEEOaALRjLdG
U/8KtVD/D/p7NbVbI+mIORL5+154duraQsyk4TqoCkgAeA+C8RX1Gyc7m8pO16KJ
jk6Wb783/EiId69T9k9hHyCwxhz/ryoy+0zQM3aCTlyAhaxhVIyndHp8G7qvxR4Q
8IfecW2B/sWy20T4zb9dcA==
`protect END_PROTECTED
