`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hMgOlb/G8WfDOj5wqDgho1b9QA7j05mC7J7bX5hT6P/pg3CN7h3AJehtPGqvpEOM
mnZdB9BFMeAnuaXhUoCZNEicBPRNWdwcIJITvrmVqL62gPCeHMCx0B8A6Wc4Dw2x
NUP/9TTLg2hBnUDlNbzkde3PDFDXyCC2iziKcym0XqzcVKoXhxSUXWBQamuuc+g8
LVvk6HSDLC6kCJm8snPVEizG4X1vpiJUFB0WTDDk3od2G7ITkXficq+E5cdGNFy4
hZqrpSIEB0vRCW2V3g9Hu7hlvouImeas6hQblSDfveHj8xWPzF4h0ajfcK/wlLSw
3clSvqXJcotx5iWe1PEMiwiP82SDiMUC9+nVI99P94CG0Zs5CNqcoQSEJ/3eH8Qw
hWM5pUbQE/1nIwFPbkebkY6bbOw2djiobuLPytjqG2iGuCRDqdJv3QnToOEVFvll
yTqxhtIxa3gZb3CyQxmmNU+BMoFelL8XLOOArPSJ8T1wiG140wYwKXlf83bH4jOt
C1LtAXtJ1k3HrY2YfW0nWkF9LAha1j+u9MdcGk78C4ZchmFoJN7kcCdHmY8jhm1/
c4LDdaM4bYK5ZrMxG2M3upahngug3Z3jmy13XGtML2ZMtIhEaS/dqub3PP2T2rpP
jJMVI4Hiqj6NuzBzB9x4ilJbZLOqzwexYeDIl4ZaEcdfEfoN6PJVwYPE2yNWQ1ha
37iecN/amgiXJcQeU+4wojYChwlM856M3BovavN4zuQ=
`protect END_PROTECTED
