`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
08NvaGjeg6RCQre8aKFJv2srx/fKnuENndRoug4dY6JJWZSlxB9sdJozJ8chPeUr
HL+Xg1F8Z3ygrlI6UOzfi8Xv+JT4NOR+WLWZDKiBXK/guFcAdgcA7+fFIgul42Gn
PmFtXB/zUvvEh218h6JBvzX54mxS4esA5hTnEu/6NBiRNBsQfJ+iCzi0sFcKpEIX
aAa/XErZALi3yNOsIju/nYXwPAjuCqj9mre4o5dA84GNHMBHE8ldcICNr/l4mFtk
7jYJxL0d6P97WgnLnDSnqUCZcLiNMMl+GN+xo0HDWdVjONYhAVGhcTUIAmJETIKL
4v3QJAtA543ixBwBo6fOj/eY5V2/PcGCrCMN3WK6M3vdOxcXjqnO6gTqv6ta/+0K
yf71GCLHqBE/bL4DhgQCz4Wks/2Hc18vUtyRYvxLVvv4aYQACJx1u1aDyOVhT9iH
1i3dZLq61QDXocL0ll0O/5aX4ypi2McNaSUQoPXzQa406tfgNcnirCgsdYmHspLw
6cIfusfQ9TkqQ3ya0uTDjQwO/tlB2RNjAZrX0TrrC0CKwSk3v0WUurreNKhLUVtM
/9widGRW/E93OKX8iuzZDoOHeFDohGg+JopXeFW7nE7K/Vok+oXsKPo2LqFWIcnr
r6OmfnMr2UCFnYARbG98NKJ9S39h4+BHisg9IhHyJE+AfvrKBPXda/DN5oln4P/e
h58xhmM9vmNjy4p+C1xARXStpaDXvMle+zm2qPTxyQvaje9afjmDyFSuDc2W9vSi
QVegOW6oIscV6ubyFeQG+g==
`protect END_PROTECTED
