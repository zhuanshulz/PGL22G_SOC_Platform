`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AHGg5vgPEs+XbToXvNkeo0PteZHfBIm1u9ogJPRpSi9dBVaMtI3Zd/ByDfR4eXS1
T1EwwB95f9IvNnxXNN4d3+eQPnQS5KtDjnbMeKTI3WAHpLe/aqHAM6y+ysOSv1B7
sLm1nJh6UPqpkKYfW1vIuVce5OvTQU9U1B/iijqbuoQwEgW/gYP5qBlPNMdejGEn
w51p1T86sLa+AHWHLascTSXVf1xYCXF3QqAQdsc7wYX37drkgPa0PMLxz/bFW2/3
HyvjDCS180nZUUAXeqdmbtJok4x7UY4hAUS/PxArhwlHgrMdkQYAl/rF3e9xzAOY
vVAb/JgVVRTLoPb+4rPDRf/fgsjKB6TBHYNOMThPalQ7n/5NUqll9XKWjnNCJeSi
fqJP/fLH8T3KFvkiwZr6VucLSVBbZNqR1OJZYdEmCIKOC1gqDWffW9CvnKBnFu7I
iLyPdWljG7PVmW6gJbZcMsefBCaGfg+vwMrtsO/JQ9n/dpiaRs6pfzeqx5a2+G8R
6CyjK9ONbhcOfpWymeVfvl5KzwPInsdfDY1NkZ4MmUMnRH2TGLNsRwis7geZdeLp
D+KiV1HzQcAp2GAvXabQSfCKbRI/1+UkU23zR1eKSXavsOYxJX7l2Db2LnNTkXur
5HtcGKdiYctozHG5Yk4+mNKZTTjH/M+BpUQ8OIyAvsPWJ0MmhhGnwWSLOscbXs06
4/ITipvUCHAgaxaF2LMIKNxjTh5ys/r9//utMMJBCHEV1VFAV8dM/+TzT2xm79CR
quls8D/9vjo3SJLxXcsbGidiYVPqP/eG8Q4letpgNoovc6Hi1u0Ngc8xnpkIzRfr
QvkFee8gQfrnj9P7iA7HNQMdXqpupTRCoZJiXbQ15dueESF+kMG5XiBkX/73yWzL
/48sxPnAllIEp2sePzcA3ckqs3C2W1os8b82a8aoEM1TRaKKOmI+zaVBtaYhiMiW
8EitccPK/RjH/wBo8lVTEwFjyIEItC/Kdb9eJ9srL70=
`protect END_PROTECTED
