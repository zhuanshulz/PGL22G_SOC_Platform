`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tMi2Z96u9j8UTvS4UpUWsHLiqDQWiUF0OjWNJygh7X2MEvBrIyu/tC6WVz5rISqk
8+Gi4eQjmFzG6hU9UqNLfikXQEqhIhp1iQz33/c9U+9ctAUqavYmYCaRK2g9r7G9
1DaiDdecQuHQIjW9WoCkUdky+o1kQcj82uLm1mkIbsTup4kucOlW+Mx+eicTuv7L
x2G3CLRe8Teod0CDgrgt39QgsltvXDtMPYc3g6yMqtG+a3xsijjprUDCtC5pG9Km
Ixbru3qpAWLtORwBYvDUhlt++Ii7bMBlmp7X4BUB4nmjj+sUnU8nFPGr1nSPMqYG
JAhv/D+98VJwk7lW5yFHTEGJh8qJ2ZQfitMudqIMUAOd5qQjWdUJlya/cuphzMS6
JY2yJ42K86klvITWUBihCdSkGd6taPJkNbe/oUEXhhUFcDH40qMMgq7ao+StAmHZ
yImsL8ZBqAHuX0Qb+VI2hhh8mr/ha7AZmGamopnVQX9CvxrQN2C7gYqyYDhYYbDc
eGQm/ndkJrlZeceLWsAB+DT9G6ErCYqdDrtCdb2dITfcDlTGt7rg61B4bjGkMmz0
uTw8vg24gTT9n60RfWNYnVYnoPHlrTAL0oNhxSPzek8=
`protect END_PROTECTED
