`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wpcpgi37AOceIW9cL2DcWkN8MugZAV6LpN/o264BKlWxfU1MlWQgSCWEzHoKh/22
YVz5tBnqIqW/ck1+qmlT0JNGtVwhu3unomhoR8hg1cqHnLj1d1pUU4fibqZRZWDO
6XmwMghhrhNo8YGlYUASI5EJ/XjekpVMQ5JhMOPIdc5RtXY3B9SLk8FKe3KkArG9
I3Y6AtgFT43NNOtpUNo5S23Lxw3pRbUKZgVsLS1q2p+aW/Uvaaoy14UMBEpiUvQ/
zkyD4ptgYmPhAfUt2bAl7fuLB/bV3SAFU6HeY00asV1qHOg5ccIqEB8/Wxl95tAV
zMiUuyHvpY8olspVxUdwyrpXJbXL4K4/9d9p3dZqDNaPwjQHB7AJMtuRBP8di0dX
QaCLhtOQ24ooEp2D+LrmMye8qiLvq7/PRcCFUac3aQ9SC05rRCclO+SyeuhPvCNw
8k+sORl+ZDNH9nVFQPxwTX99cvzQL/u7O/zh3WQcLrFFRdfEqhX1iGLf+2K3LvmL
5fKIkk/P1RnFMoY0ifMUIOWtQohqCHNojW4Q6hc5nrDE4qEuaDSQ21+RplIa093t
eoLQGh8r/d3PqauosihxYBZuC4PHWIfKJODbAN/Pe6I3ADHBv39RDn+OVPPwb+WE
GL4m48lKdBpCv/b+CYrMD6MoWr2LRkGrhFkxH3kUAQibk/2mGpo9QIfkcuniQzTF
3bRvnqjxnUS3YgSEY34g09HzTiRJPo4NiHYftgQ8h6rVgIlq77HEcoyDlsn0h1ND
suLWfq4T8MjR3Xcfpp8ktVMQdnSttBDmuIq5X16dGuk=
`protect END_PROTECTED
