`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6OgbYi7gLUqPl/QDe1kMJHXPRUY2laSHWeJ7OKxlXN1cczy+KcCB89vRiZQ3lFTe
e0xT/fI4SaQzvSk2QLYBGpce/uPidKeO77z4XfuZ0sYwUN0k1DJibL3Ai4mzgkoo
7gwuOcwBm2fu8S5Sa5sj8JOiAJwXs8Pze8f2xbw+CYJ+Iq2nFNt1VVLjrjftzxIg
K/WlIHDaw1u6aP83H7OnI3gPTHoG44vwn8OEWBdqtNlYQPI7hazDFwYBd4xqVRmU
WTsn8wCt9KbcQ0/ckqRaiw==
`protect END_PROTECTED
