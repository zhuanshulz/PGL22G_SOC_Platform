`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T5VPtrffkZ8Vz1o6az05+R7BlQPDoyEEacV1zzKfyJ8cxiBapu+z5ryV1Wj/DU1y
XtbNcwJ0ax4r4e354kKGRUhotq9K/1ZGS76jS/k1R/H8M7wbxYoWL0zawr66TK+P
Mvy1fZguf1KavAMXGzba6HgxRnAWAs9yFqv46WpyJu+bX+TVfvHhRx+00Kh+wLl/
jJ+CEfKTLWPaK/T2hJ6+UwB+IsjvhcMJqxRIEwMEwimb2mdsvdp1x4JtK4aanuQu
l9yhWMiXehWVaHC9he+uHCbIgTxH1M9o3+15SS02JkaBzThKl7BjxXVWAJrxdG1s
zPHlVZW/+hy+uM8nKlPSSKE++VIzXPWiSGkawDn2Ekocbg/j3Qxhd3ZAjfN1sxU0
SrISLoAG9BALqRj75NeXt4QHmJz4d7yoM06o1Qrxe9yL+oH5NZSpB+15lqB+yY8S
FJ6xhmZ0XzpDFX7ff5L6pA9VGGCj9dEnRgV5b6RurAzhi9y61uddU4dFSV1SwlcM
MwTB8qeIkl182vMHW5XOfDzlCOJZzZU8ohD7uZ2WNebVgFp6ZAcrO03FmBkg8idK
GHUAwRlZADdKaNqh4RQ240dt+gT0pMqvbHFoUpW4Jj19gBn1RpUCjXCaPohFN1RV
vPqWIqAYd+xyZnNj96ziHUlZtt53MxztRCwVW4Wi/OM=
`protect END_PROTECTED
