`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
waAdpstqEkgzFUM/YdixELbLfVddSFZPLeqviiUWK8eM2/WpeLQT2pHDgvLSyRTs
qBKPYwJ4In4gY3GZAQeIdwdwX9oTC33VKH+5B4Kgc8x16X0XHdBnvr2kIRxitBfu
GBIYdlUJBwZQr4YXEd5IVu/OHBVKPB2P2YXUJNcv5x/5s3/vIdqk1VmXanuqp6h8
ZxqSzqS4r0OsnbTQpIcULzjZiwusivFXQkynh+rU6hp14AbegLAQXnf5Cac1WYCR
RTWK9TCGpgbMHq3p/sa1fPZ++FZZaOv5jPGlJpouVa4/xkZKyLF6yZK/YHIJtuct
4hmfoH+bADIjq2oBmTd5Nn+ex+H/ZWHTpBEdUgMSCh5XPjZcaxs4MWquuhUNU1iR
fsUNLgsr0LFX8fB9cw5nhdguzDzCAzdR0hAWdzpci4vK3N2nZ7GkrDUND5aKrhoX
tI2C8PBnJRipwvSsDvHwP8EgA7mDi/j87ZLVUDJ6wpoUnHnQ8i4CEKVAu0lG9y2R
yBet2xCQ+hwOyaCgpowchYxkZO63IsaBLefEmjy5wpSqtMvys/AMVuVfHbQFVDaL
lOUzqxeBsnzLmAUbVgKyYn2I/3Lq4Q9fiCXd0jdI7wlvUGDJiRZM1woCpiUQdTyR
FKxkG3M3jwAE8dqpetzB83KBOxdpNbNGCATo0t8/1E2IecX0JjcU1bMjsQn3JKcf
CpHi7EuKWWlHCKry0hQzhemR4dCiBGHRTa4NNlfHNY21QQji9PqpLHikyXtuBPB+
PxBYKaaZmxhbndR3X96zT+PdUk4vSkBZ9GTVpEOUQLO4spvPKXncWd8n3wV8RjuK
sCPkcRpJa0hcivClxjBOq8i6RSwBxyh1P7zQIY01fDofB/X09KJtdGoxKfefTlqI
eL3qABVeDFsJgOQIaz9+eyc68Tc59a1AYZUcRhKOvXsnshCbkftDWY5nzbnoxOnd
LMtSlC6lYKQPCkLCuUNcLpgeJy+wLAOu672xVu4JNZe/l+XNHub7fREW5iiCsoJh
j8rEsn1s0yzDDCRhh7w169YnKbLb+I2HXfIbS74C4BwJVGySFxHIpm0pIWfjAglT
kG01wgKWKxDCgfVxaZBhBv3OZBDlV2PjGERzY5EyOdTONy0dNX7FdaK3ESb0vVoY
PrW0eYfw5wn9YlOIQxPru/isKMsONf17uu61pnMwTrJgbWI3bjgUbmEmA9xdxqzB
X6RXIby/3wd9xqBodOscemjtC8gZ+lR/6kcL7dFKyoRH1P3OG4IMRGTilh+zgpxV
d0bMvL7r+pQwtdN1PHvCuMQItrLw6YjfBKyzAgZbOYe9y0UCAqyzq6ePrb87pVVm
lnERA6Ei+aAUlHeE7t8uR8f3had1dP+1NUqHNvgB0/zluVHhbpCCIQj/baadW0U2
YTUEbn2/4zf+YEYvvqZJMI2yUDtiLRPC1G4WVr9dHcUzHKO6Tjj7k7v13eF/va3/
uGpTe95rdx40q28ll9FNHCfUmMgFSpbrBQ44zICE21oL/tHjSKz/0l33JXiBungx
mfuBQmvJwArhW2E58+/FItSS9tM7G2d9b+qv6Q6WkBx1RXBTd7gBDcrOn2yjJ2cu
NYSBuZvRdRZgT8ONtFcFG67xVhzVQR1Qp9oEHWKYNZtnbYR3aqCwn76zY8xH7fFz
vVCFixKgosvk3sHVRzZoVw/0WPZSLopxa7hJ0u8EMpZNdEatN3O+W7sQ8DilrHVP
R2E4qo4SoidU2eJxkxw0UNdS1CoIhzopHddivWgYtluocfINBfFGoOzrnVCuYirc
krtCnjHWfxue8Ort7e3d795VUfLBzanGniUWYPWvJN8EfAwqEHeM+VfVizRDf/hK
NBcff9TjFlm1h08nVhSnTMPNdPTwvKuuHuvRuzSyLZzScntbztYVSzmYr6OngUm2
1m9A3X0JKVEmier9H9+zrYPUufN0ilKqShGgezOauh0JGHcGX6FE6UJhkuGJtvuL
2PBHEZYGtDf9+99ytI556e5te8loaGies0McQyXHNCwnNEOtI8FRBv/wyrB2lrxb
n01/rj58/gBen8RHH/p+OQBdYdWkWjHZGb7ROTa9HH1WOyLXTaJC5RpXiY7MZguo
+60G9tEctRgXMg1ICFjfOVuif3wZGGVGFiRpp41VDmw/SfGdIxaz+sM9v0W493/D
7L9zscR9OnpYohUWdo3KUaYK4z97+9C4GtXZ6z7kcsmeufWURVoI0DZjPvxTV/bp
NovduZ8w7GAiV1RYOETYEp7HLaK9qDQqHwBZrHTdUlzEYjp8m0unElV+Xc3JHt/P
Hc6MA9yyMYm7gp5457vFwhrbx3b29+xHKugBKemTHK0K6mI+AXjmUlNjtnon9m3+
rOCOgnt2Kg8EvWK7evwgOMvaYhjQaj5nZaka/gV5Bi6zWS2aG73hfFVRjW30x8x/
Gp8pM8UtsJVVklb3DSvE5gcGOC0y0Z0mcXFo59GTRES7cFm/FISrWdCrP1AwJUCC
7Pj4BgzBE8+b63TqYQ77FKeLgF27nLmPdyF0uDiqztBUnEr9+gpubfWUkZMvwjRQ
B7PjYfPQIJiYxTNHgnAzXS7oruvEOw4S+bQiqgpe4SdVW2JVi4ElWoMbxcdFaiTN
SWv11jVQ5WYJntRZlSreKPT+Tb7m/6a3T+r6bl8CCAfh1R+9AuG6Y4KqFYNPTxC8
V0fa1BxT/U8/4zpvkQY/cMteF+g2eF+CMLBv3ogrZEvPpj2vXK30trbsRuBSTbsK
m2A/PuHR0dlUTO77uNgcd01Ek0JPzIWqkkwRWY5Oaf9PjMMt4267DP8uNBwgnarG
ZTL4tLFSqPkf8UiTQbBLaZoDSsKa0EFntagfveb0oxc1M/iDLRWjNx6LVtSvNdql
Cy1mgLP/dOtUu/Sp3uz2wKwQxc7VJcGYTcHdJwEFW2bkmk4ZLyWOEzadZ4gRZcvT
+MvLLFgpPQH/0ax19FWP8p9e+8D+ZkP9XAg9USX3QXYW0xEie1qX2zqUGNFGl6Lq
J0oN4Upjx6+hgequXbaqcBtvvxkRCOwambh92YtajNtP7ukbda+yJdAiqhm6QIle
DB68adjLSHh9E6LdDTpOwSGW7zij6F426b/6c03xU7SiY/gw8VivPN3cjHN8Ecfe
sAx9kdneq++i4ItY+mZ+a//yKdQNqQQnkpghhYLgJqcksq5/2D+L/h3SLl43gk/f
OuPkg7y+AsgA9rUC7SSwD7PQfYiLPeTraOWLI0eYV1kfXq8FXDfkeE9DPNnKgxGO
VLRpo59KSajxOGUan4NYcR6KfpXeSv4qc5X10yX7N4aTg6q6Cq6UYZhKT1LOiQu8
J2rDT1Dzqmk2M9AmUbqtRw/UQkv6EMcMKzkIL2G5YlGG7VNS3EddK/UKOLXK/mM5
0tJaGfFysv6ld8SMrBlR96a2XRLNJtH38egqGGzHq6r863Va6dL/etMvW0pLz051
Vv5BH8/5JcE7PqsVLpLZH5IYRcjSopgNNS40VHfR9OsE9+r6DUVnnGAe647u2FmP
8iE3MoWYD2wTul5UVB+IVgZlF3xSLY2LfpuCwuJZT7OQrQxIE2umaHqqG1qbvEi/
tGsyWaySvWvodOOeUPrJcoIUBrNnCTI0EWtXBGHIgpZxuSVB/wW3cii5SSfjTtBi
8UPXqDEdhVxUplB4IBypAoLCfqRCAe6prMgwvfDRJ67XOzyGFz0HYvK+jf0LItOe
bL1YRfoeqWOVizz7b6MNxaSwO+Cc4SMFECaUDFQ7LOfGLBEqMeQudguFDvFJN3ci
rtbO6N/Ya859hSDKf2ldUkrF1mhRpHm3fy+kkcgq8Mw=
`protect END_PROTECTED
