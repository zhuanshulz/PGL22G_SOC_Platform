`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Sda81c7QjBVWwSIDVXaymhBc8ppEYV0N3y4miEZCsoHeNQjN+3jR+J3CAfurka9/
FACh2IfZg8YwUABsz56Q7Km1kkxb9OCl9LeP1Tp1pw9bLYXZYOFTzEpf0I4R47lZ
tHtWMd8AT2sVy3hJfCBBnbbHt9ITOpaXfUx9MAeyTfJVpUYeyA/QxkKhd07ORKX8
1zb48iMb0872IZ27cMylXWbtv+g74kIO5XSk80te18Ds944hUk0gqhMNzCOQhHp2
sNa/lVbmBu0nxdfR9InjG3WkX6FhgOagjJtAQIJ8BiBIE0yAF08E1LFiqodfKZRC
7MfdBLNuZ6Tivjl4pGcjtaGAXzbpCe4NwwW49ZvgMwnZOpBQMD94dT/rFBve7VWc
XrTJPkbdChDXdldCaTmjI1+UCng9DGqxpoADDVIzLkZ8ltJgRFRrHjlSQP4+Iwf4
AO7VdIMZAXNOFxKNNm/qQ7DNPvLLKFi/PzPr5LvQRYig+w97JbMdVDF9uoDcQzQ8
gHE2ZxWnJsaCs84AG8O2gKl5sy5U7PBET9A8s9krsmYe3jU1dDMXrpx6yIGGoqy4
llLI3SqgpI/CDvBwbl1QTXvlkXnCVEZ7lw4ly0HuiqhO4rcXiJOCP42CVqjP3vSw
u+maVAI0GmpqbVccRqOwsIQtF6gXbLgefnSrnO8U2S9+jQlYtcu7aL61e6lLRfAN
gZ7/PLANn7juyE/s8xMj7NXsv0ao8SByYIz1elr2eGHAAXh8mZa5+i3YeYG1apVl
FeSQGtl0fbqqgk1J+cYDgc/CWFW5UMmySFW0/6NxVIlCFVetICKXZTjFnFt9etIY
76FgnnWdpvmqejq8eZ+FeswIKHtK0h2NHdo+gTvawBzdo7RY2Y7E5wHIO1XNuO/c
4CN2BqkUjc8JzdDiyb/+8EaTXNNbemjdS6V4lJ50/ghFWVNDgLiDEOmNu0WI0byr
UjDGIJk2tcnWiKmWBe0v4BdYY9PPdcXxRjcu9NmmuWGlWMo/kHSMsqyE9Tv1Z3Cc
3YpTR8ttbIvyVXLrtBTf8EQWtZio5Sa3XiZrpo5N8B/SJYHxNPvg4FTdgVwE0pls
U88Ullp4Rawictdf6lfbw5h9OSLn1aQ4D96w5MUk9zKx24f1wLCSI2tadWzUBD3t
aZxhnrNVNKhsfKVJxmXkMV3isLO6Bhlq/qIqotjuPFuvQgDbA7gpoaxczggwSodd
4TDevA3oqzCNjRPujYKaDflUjmKJb7iC8Rt5yL0E9CK5FOeNr8Va3nnQl5sleeUu
I7Rs1v2QzunszpTtLa3SbaQxQ1YwYL46kBGBZTOmLyVYadXdsf/Wl9zzIKW1oWg3
rPSUL42JJ/LZAG+WeajNJTmIxkYemHQ3KC9hK12vrSpJ5eFDLyBv7KoDWFvz2X7v
y/+Tg9c1t7EXih7p/4YYocwToZLQXzq+yKAacHeRrl2OuiZFQpQK8XjzNefSzcZU
bnh3mR+KTlGDI4WRB2dUV+3YK2iA6alEeCJ9BVgM8KCjjsyPBS6ebRvXtWGwXyOB
l998sDcToq06vpJKT7CTxSFWQjs11/cAHCLpxduIvPj6xdftIh8Qc7tONtyJynJH
4RdfZVxLq41piMN+AJBmRsD9rBun+aq7ZlTm3CUHai9q4b6h0BZttR2gVmmLS0UL
O1NMm4E1NCmZjrlNTyiagfEtAARhQ3z3vX17Yz6WSEhj8SoyqxBEFu6fC+JgB7zy
UD6+QzfxoXScLGlhHQC/JlmaL4Y+bJ4djXl5ksh61MhU9nXCR3filIfQq9xpJfKF
RB9Sn6BKxvLKMbFxK9/SlESYE+1NkgbN40hjSYohOEOhHPnLHj7GtXVZxojiXQlX
4vRYV1jvjXa9sk9BcfDMbgBXeZqdg9yIHVJLhD8I1+wnHupMZKNSh1VBY8e4sUpc
QZ1OCgpoyfyBYtqiAPeUK6yT6PXidhogYK9nfaFxC9e6bJZf2GXSJgw+9RWIjw/k
XCDe2WZZuQDIJDLKde5HcbT3932ByBCz18hBeyN8z5KRUeMJedq0ZL0ll9Xx7b/Z
RCPcijYMW481rB+5iXgbQCY/ict9gVWST6R8v5L06GUlmlroLhnCfrW+A5OgGtKU
lvrmBCLWpo/jAdJci/IDY5MC3HTxrh3LJBkEe1kTdwgQDQqLkKAP+IpwtsL7/ZNx
7m5DO9JUCc+F7/nQpUDAxxry84WkH5gXfWsgWC075hLbwjUW06QCD+Gk79zU/sNU
ZgQ1V3tmA44n+gNz0QVesT3hLEwd8eqHxYlZ8ezZ38CFCyPoAyF370PEd9hJ1YVm
J7kH2KqixzsxH9avnfkjse/DMnBtB6mWTMRUJrBJps04fNqeJEkFqZW8Xteab3eh
JWUAEx38sp6xnrGpwQ4xTJLbPuep/Ntqdbwyv2XpDt0AwgovHgYndv6LUd2edQGT
lbvdH7vTeFAQepq+3NsMI56C52kAV9034Y1jSAzTLMH3iO0pGwThbVyFJCYj/vgG
ZGLFKTauisLqYT1V1dW4S0qRz2Z3QOpQGn4sfy0PoHbd28RPxJ4yhf4Zx2QadTyv
DqaZjANE0VbaLPYUouroFZDqbxNWiI3jWgvTQQfngaEClo1z5pyuKB3FAi+QBQ7B
cvS2YEvF5jKr6qjLgZ3h64f2Z0QIbyv0o6MzBnveXnvUw15IDiocNWrQPG0j5irx
fJ+J9VOcVsMjBF+Pn/lEzm5doi+2jSNw5OYIhypNW6FBxyXiqPur94XqDwe27klU
uQmtBSAWaGkn+wFPj5yfMJKY4SKcdoyUFUE6b1rxDuWV7iNZVWUwKgon6/ubW0Mk
SUeP+MYRZ4ydWM+JYlOfjE2XJiWKHJJtDUu2kjmzGvlmP3NJvCu/utvIZmoDviYw
qEC0bE7MCwJXmD84QPHhymYP+nNxJbWrWZqkCapeAWW6k5OmSWUNVCjDlRhCS+Nh
KV30vBu+V4cPL0AqK9Dz/hnL/rzTSFovnI5Zw0szo07slPOzbSmT6dDzW8u113E1
pWKc+T5vlKo/qKTe8ayhv1UsGhPNHDMs8ckDvigzg0ipN60PUXrjYlXo9/u775l7
S8S0b4LOfz1GqmGOu9kPcnwoq7vN1w4a3VTBYd4ACcam0eNJypFgdAup1QlM26sS
L9Q+SPfb7i3n2oGCdAhjWWQvzZFTazu2YDcqwEuAwM2zAPSDlX3KVyGfoI6LZGwT
IXfI4WbTOcuTJao7WNXZzfCgs+IrZsktW4aAsAE6jQKAL7KjqdNq7y2AcN9uXMjQ
eowyMI0CBPT7gPAo0Kypf+cFy2gUZ0ouX20qDvW2ZAnz3SPNnz7zSggLDSmZI59w
rfPEXX1HAI4lcnz1v8cbWPZNC6fK3X76WdMaX318cAWlFFMR6DNqsb4W1UNxVtl+
5f2Rc0yDXY5b22GlrQ7rB/vgSioXSf9Dpm9fCn9EoTfpbgXUjvxnS4UyH2Ud1EDS
7ZsrKwn0ngEolCDJhw4hR0vS/51GpN/XmnxWt5Tw+ms/BplQSC7DeIcEduZ7QkHM
q3lwLElJDzgdHk4uXRSkAszZVPZHNVn9MPjvNtQiak/f1uy3YLFlUx/UdvIbJ4SX
m7qqoEGdUqiS+aRjd3bdk8gm9CqWDTFp7XeVFiiCB71NcGvj7AraRsCtrEEa3lr+
xRZ1K4TcGBbTlegh9LCEBG8aiVGeZyXTZLR4ezEeoAnh6m+iSafzxwOudL+nBOtS
NqW9eZ7GeZp6kxqcThvoD63eBc0hFSzFG0YE1CmxGk9tPV0p4m5QueJYpQuLaETx
Njca/8MIF0ia4CFiG0XjhCcJCMjJAx+4TZBiVFTvfsS65+kFC2HiaQRGB7apHzQu
Y6Ky+q/Vsl8WLOyhwYdwTfb+iyuUY1BfE9dDphmyitPdyt+sxS8oH+jG40Zquipv
Nnwpkda7vezS8RBz74BG+S6LduBsCGQo4nB/ah9DHPqW9igJJnmBf67MRLXkG4NN
oOFRPowUc+3VR2jMiVj4zFe06hkV2/z1DUDoYEaEHIqv2Z1Il0RDSyjy8BlK/F0O
zdjtR1cuNw17A08B6kCx2hbm+PGeknOLKwQ00T/OjPNKqrmRYOBpmTB2BpyRFBHu
f2pWPhP5YctjEcAkdd/4OAweEDXEh4IM3+Ce7bZfYdqCTa8hQ3Hh9MoEOrP1PUqE
+xpVBt20gX7aHiAQZDxzJxguIu53jASHCQFRuNV8XGIXUgHKxKlb70jKTgie24uj
e7vrtpwPtQSYz+JD1A9/LOec08xDzB7gIdC7Z3x3Q+rs0zCn88Z7Zkt9OlO9ey6G
5XEj4Crj0K1zhfslhdg22IKARVZqsGeFWm+9MgxSIlvwpd2JmKjpUW3SpxD6rDLC
jVnM988FwDUnBw1/Sys0XnBfZ+Z9PCM81ZtUj7ZLYCJbdKdVhhz1Gi62+uPII75p
sJ4mz4SYoquppDTrr5bQA3O/UA2xQkCHi7ZolotMNyf9QB+9alsqux78c5FCr/aX
7OWptsJ5Ld9Ur1fEAk4o9XgHPBMskPt+zVPPHjR0QueI62IMHfGMjY+1SFK4fJJz
RiwkgS/0Emw4kzg15ZvcIBwQSH4DGG5HuJXmM1nd/49kGoVe3oQH8w8WnRHO2yQ/
FiNSbbDcsibTrjf5LZJwkcQTcz8mkbUkOld1//izjz/tPpypGE9/cxy3ghvw53/b
xMgDa4ZG++1HUFY5Fz18JH4032tDpw/MuqJINgpLuv8TnB/eTniR5VlWukbTkjvK
9HBWnPEwLIPd8+V/FRo2IBQkBSxKbq5LRfB1LxNjbxeH2KRd0Cbib531NVVpKlqn
J0WdofJ1PQl8hW7LhIJKh4xvkYIz4D5leJRp5cjcj2bM71c/W8yq+/Ma5x+Osb9P
WLdd86n9vLva+uQsbRcD4uPagwn1X4kl/SXWevqb1Z6pInvvQ12rZH77Yh2f2qcO
KMmCPoqbQd497O4e1n/FP8sMratpUsAwalMx0ZSOHubCImSRaH/KQ730aBQGOIqY
W+8oC/SjpbNPQgCBRX+cNnSFPzG0QPbzXe+GC5O57qwTpk2wtLnv3xcqnNxkIVaC
UKgH8evImT30PiA4hiqoKhD9B7BqkAwwJ8EyTgNzCmrCICA9svTj9OuM4ppjQ+NI
HsoU+rPEWn2u9pkfhNsgkkcNeCXEnwuRbEvwrKWr9ccOVCSofsos+6lFTr7P3uMh
FEmTGOwka3xrRSB9hzJUnTyIYy3FcMHKjkL3KpBP7CEjO8KylNOJFr8l4hzNWmBv
ZY+npWKhFP+LHJ0hOEsViV4Bwpv+uoxPCKVWjB5O7qsG/8BOedvv3AmVHRAEaXL1
UqMsQnyUVsP0yOpViocL9Lkp40abXgJIMquShzdAFwuWNMcFootYPKgwAInZYB9y
T1x27FLCdo6DUY//CPm3Xsm9eMMarHBPuDg90ub4vu88NmtiAF/qBR9q0eoaUIcc
f7q23Zd5kri028R0CsvYHZYaDZyqJODeJcprlyJjBUbKQwytUjWJUzJO/vLx7Iyj
uYPWt/pkR94AHCibeQHnbTbY0XAgWO12UkXTn2SAeB5cP/noIPiORwymz95QEFbS
dzUaWUImGFrO1oCgZpHaOQZnVd7HB0Q5ly4+gg7czQ7jJuqrkcPoKSXBlueukeBO
P6kyyhrs0wcA2Y5kN05aEL4TDKCDDOiudUNQ1Vmh4302RJPAmpx8ki0o2bLDagCR
wIq1q8cEa7MLV1rcPsZGl/hE/hkMG7eyTH/PzupD0/rr6RSxuDY6+SByntzhLAXC
UAYGEp6wDcg8va900YpwdHO9mPVqTM49Ej1TIUwgY0VJsuy7OPlUP0Upu1UJPEz7
pvXV0RseRCGvBvn5vFRu+QO05lAYRaQdZ6e3RkmdDRaZ16zmmIeKWDHYRygeE/YN
Q5e+3abDBCH9t9FS26OLD7r4Oln/Cg4ZVWVPtU3N7najBs+uLgaErRkQqgjtvAGQ
kko/711SlEEZuMROGGSga2CI+aTJOnnf03IcNBg6ZhPWl/6nuJBYrEe61tVW2wgJ
Zf+LU5auRNbCobvgu3KxZPAqM8fX64rQn6vheO5P/4at3xZu62H1O3/l6pP6M9GV
jjFszt4iPyZJmc83IEO9GQmnBmEVAPK9KGf9HECxqgh0dpvUAESoHXaZP0dz5kb6
p6dxN3K/sSWtkiuvSvPepcsW3yTwmngvc5uSdA7hxEV3XH06NG33+rFcE8ETdlOX
2jYtaPsyEBvL/mW5dpjaohq8v3jE9xj61S/+MeWb9w4Xi3O+wkw4wFMjkKAtU2N3
6+1CdszaFbO0OY3HUfOmPV0jP21HWJikbb68sAj8O5WGFX3bbl0+KPFPqQSFbbCM
S+TMIfLVYil+fSYQAqx2uEhWRp/nwRkkkbx5qwe1xAB4i8ymUcaGkB42VFcuo3On
v7l9sHDxrZ/f/DtksWPOj/LeKNiKusgmymQ6iZ7Wv1rZX0pbd0WxsvytEv+rRkGt
eBAyW8dgiKAq2yIskuWlL/GYXWK7R6Eb278TL1lMGzPL1WTUyNI4PV+hA/Rwi+2q
0W5WYvH2oqo5S8WgY2LTt9+xukY+pEWqgyw9BKZXYBEmKF54s6lbPMIza/hPzq9z
g65dZt68ZJe7y9vTGiTCvke/eNfI2+Xc/fL3bCLLLveqMOHHjCFJRq5bDtYKcGkv
06m+cWpitTz9HetiVTLx/Fvt+TB/ZqLUymMnEI1kOklW3R4Uz6yPL5svNOTkexiG
PD3Pmh8tHvkALAW5DWdioSSJNEU0vsbKLa8zSS0dfO/SMx2IqEufD04zfozUF/ji
43Yn3J53a8+m6UaPm22tF8YamxNQAB9jE+kf9YqyNGUKK948Y5R1rL1GIVmyLqZh
wq5V0ruQ2XR0iw72v7b6eR3om0xlngU3C7pjnCZgT//0/8QW6U+Tg+75ffufErNl
uJz711F1bWw2LfNButKYC9AIhvq/axub4zuyZ9OOH7HD9dRcIubVID6mhUcXZ5mf
X2fZb1ezxXkbm6azxQNhKdpvFoEoc9rPrz4fLWOmhhZIvqik8nSIB/rX9mgWnjMy
ITF682OjZ+NJkfNAe7WdEXhxy6xp+qHmLR0+OMlwLXLS56vu99SHYIbASCFaiNiH
gmc2AsYv6UUOtq5t+D6G0qajffiv+CZaFFLO3zI0fUJGLExPBA515BK9BjmLOypE
jyu1VM+duwrdhzLr8I5mNeBgL0/odmJdg/areuUhBz+rOJAPRQTgeS03JECKkr0Z
1mbfD5UL+jYUlLCr2D5XdkXJuRjdZbYsY55KaJrV7QgRGb86mSmQdRRWt7KpbTax
LVlpp6wMBM/HSZgBAZPXPHfvodLLmjc9dea6YK/buL4VPWVoq2ayYJTnQzGd+oaY
lMNU1ovRsgrdQMZwrs3p3r4RjKD3ZKLTrKkCEWv2j1PIdzemRyZV7uPdgu1enBtZ
KkIEV4LZDbXZL9eVE9CKlUhrj3niHs7suzrnXip8elgWLjGAZ5lSS7ybDJfXXZWn
h3wgglwPBri8BYi7Wtd/wdKVoAnXaI6Rg8wKqJgp1FneBCY3S9leFQkEwopkjHpg
0S31qWYgtwg/kJqSSlKu2qUxQ/cE+XJ0fihGl3q1geamieNKHBdMjJOkrMLBQ0L7
3X5cNf7O+kcUYsEHX5W4Mg+ncLCC9RzWygDJdBAl54xQIL1OHo38Ts58Caxz9Op6
c/n/ivvR2EGkE9+Yk+LOIFXuoinLR+TDglBXNQfqLNUqf9EejX4o7gngSVUHaAcz
3od6KB9IRqbh1FxFf3/3+Ja0CXRhjwUCa5Cc0N/ADQfRNEicTpQSubatGyXhHmTO
P/O4q/eTmWKwxv7d4v0iZwi3/vv2hlHZvWf9m7wFjqe8CIQGoVXkKp6uX6WR2wG7
mouMWKlkPuBwChqzNjp1kc4LOSKSflHc9TVcPvYEi2QxFNJVyniXJcpzNz4MAf20
bwUA/Qv5wRU6Tf/s6huQbh+61HLLrsn1l1jycDpPQms/IfDYdo1dZbRVfQ7QHCkk
zdmsJ7CRwLPL7RfNZUk17fRUW4NzFZqtKLhUh2YmP0j8xdD0eKb43crFGVvVSbRS
MukJlZycy+QNS8FI5jGfHpCDlDk0mu+LQwHiiSL16XlQfBKJf6ioczBclvz+VVEE
T6XKb5Hiul6SkqNulWtKc3Ch6Fyiw8DboFkxOb8Du5rFSt009H2tnevbV1Psj1zW
QeH6W3v17mLeJbj6FhDa2X/LjFwS2FTqG8O+NJ6dktCQnmOhU34KmY7JcSpFEQPq
1+uEik/LTmNmJMI7JBgEjdZz0q378ZyI9EpBMSpnQE1jMRq1LBNIAPRH+Qm5WMAz
QU9ZtJ4+/YmE7hJde/FacU0WAIywqaLiQkyVHIcWTM07xXKjyQIGg93oPAV+yaw5
cQXOvJ6HWKcA6PhZ32NmQThzrgSBsLZPI1OOgcrkLC1sIa4jVgTUYg3W67nl39l5
ww0t1vUS/iq+ar+YgP6j5BB61uHp2AaEQsyUfA+bIjWrIOSlIzlEEOv5wXICNDsY
KWOIW2yPCtSzDb1BfJ9fa4LOnEj3ztD4m1+NPl+5DI/1O9zA9FLdGguUSECbFs0B
V7ivXG7CzPUwee1oFzE7RKdAU3yXajFbYIqKmCA4vQpGEIszM39dUBDKl8+hseer
xPlt6/XZGs+3/17dodAVjlv1hhimn8uJt+ERZSCmkfEx+cCqMUyj92YsqI5qV/pM
g77LY9LVj9UiyyHPKI+B1z7XuQ3WVR8VpvgtHFi7a1A5HohRUZwPjqq1okZGU3vx
ChWeTElUML8Ck2pZw5W5kQrLrzN2ID5wXUUIdLxTD5Y8k009jq1nsQx2YDUPBG/c
cnRI8z4s8VzYPFhMLzzc84Ln3hbuuaJ35qPApnrn0uZEp/KtQbVWCExBqjG5TMpK
2us/xWISPtWEpGok9tVP8SYN0M2qgQ9jN0Xr6ckCUAvmxIgV6o7PSg51ZE6ghJRh
SXooXnSeBYP2VxIMHpHO0tDB9aC5ESaptP7FDdP4InxLkwRxo9fPifqLzP3e8Wzo
9Lhqe5KJbNa0lIaOM7EmwnvNTae4gRbIje/zVu/jdbzTnWCvZC3nAkIYvQjFZxFe
cv+Da7fPynoT4jSlhjyTbZPkMtEokVZuJeQUC3wmqGE8pEqXfDik+N5CnMC9NNp+
ezg3DFQH4i9qEYdQwPyzxNXZKxmqhSSAFQUv5ZabByiXtkzhE6WY+N9POjYrRSSZ
nsIa33CJpIwMZkOm6hXpO0fGA5+lWqlOmUkvRtPwHIDRq9wgdaViy1eaBZV3UuCh
pbq1JxVWLHKtoUKlcbdMDQmbptqgATqr3p8shT7JrhV001ChsSegn1ZsxeFhaWSb
Kjfm1n8WYx7yotgDgFo5M78+4fdWqNYoQ/91NxLPAwGxtnTzj76InTF20LUKLJDP
3PDIsiqtIR6pUlJWcjY9Jt/7g0rU69J9HdD8rzTtofn3IFvsLpSk+zKiyV/ckrAh
9WxZpEOpC2b2qUvaqNiWg1CaPT/+XtJG/saFpyl6+0oCXYACkodSK7aKIUORGQPf
Ha6eyCLLJIIx8LPC5nl+yjW7qhuS5kOpa1jAHdCdLgj8UcbmCsu1pgNwUM1zxUGs
RAyzNBjML3KJmbcg7Sogb5Ttt/7m0yaCIuXalHAEsw6cj6azZBlhvF0jUU4z8I0k
19uWjDPfwXxkz3gfCuRrx6Y2bsy7uZq4pJ49Sy7pGvFHLuMDnfNN5RKFAs2e9lM/
jQYS4SEElRnSqDUKhYPo08ibk5gIjm/4lMYgSa5UBtCdtlfzl37zydfTPtM2azlT
esl/pFFo5TAAig9FWv/wE5CL2RvKyWbadnT85xRri9bqJlEM//UpsyIRh3qGJ9dz
HzxT0R8kRwXyAXlZnZYwUtjLp9puOLcBQki+hiDuLIYiOBVp/6GVq/3pYvAZsZYW
Qp38ZH75sndy2TXVpj4GA4emhH6hb4hWPS8feyby9LkqL70Raj9EQOh6zOqxdT1A
eybEVEWPD0oUf9m2limvzV5IU31rpzHYLBd2QFxMIlNmHrpMwGUqpuO1FoHY/ASx
wg0JM37FCowG2JO7xGkGRLrpM0Z6c1C8bKBPtDJRTZIHThEAMeCqQJdfzmy+IJzY
OMvJd6W++VBB13lJFx9Q2QcQR1tJx1jlDKUFTVCWc63TFf6Z7TJxmuuDty4iCYP0
+J2bshgtJhVZfZStaSIVCQ6csw/tZ2DhRg9MuCLScjClZ1j7+Fjv6GQOTFFUuHai
Y/c/Xb+ex7jwMYb1dt6VXdcZ6jumFf0JcYcJmoOCgpSPbLXw0wJrRR/DHWULLmZ3
qREDGfQ6eR9UPECnP59uJO/XCq1jSBLHg5+fr+/oS68+du2m3G7VPM+qXeWf8hJw
S/l9EMjY9tvLuff2Rnndv7e1FuTA6oi/3oKM8X8AWzZFkgrOCLKa03WDQeZZy7GE
wfV6PtHf4hr7CQnoWGsWfhINEp506bYGtIOktNuuUPqpklyXk8eW/4h1J5M5OChM
wzRC9Ha26PLQAcoKzeNw4B06M+BfoQmHBdaN3FYkOwDrTOp8YclnxWyZUGNGKxhK
3HJl4I0+UHXlc0c/s0t9XOyNwuteUTgXM7XSYuJj7GDb+nTa9TolV/zFQMdyLwG2
pb0fhlP/gehjVVyq9LzALpUGyQHi8w0bsU/P1yl5BtXS3pjvvpYrpjKgWU25n54t
h43O2BnFybM17Eb3KWI1mtvmJW5ddD9Tn5EaaJgLzDmswn9NHAUOrf1yJM/EhcKB
tRU6OcFXjayV2Ir7InP/xiROxnNh3idB3Y1d1vBXIH5G1n167hgEcXPAAR3cZT7Y
CkBL5pTD5LMKXjA/zllxsrSPsF8/WztRL0GtNa0L5mjFdOULkktFdg7MMR6Pvzqg
klVd5dICDxWzHH8VMWTXgIoKc7tQlPnIy5Xosx1A56bzgGSnIrU+ifwCDaKqyZ5U
npP4wZgGzd5wifsJSMSEnRxd3I9i0Q42c363T5bcKnx4P9JJBTkXLYpwNcX+pnv/
E/8/Vt5TN6x2/R9X3/FUBsvxriVkU64myr+eLYCXmEqqWG0Uq8tvKEKmdcy6Ru55
3ZUc+xmoHhtcc2+POx7or/7LwVQyReLfI7M3UrDNJHIT3J2dbN3X/tbrt86ZH20a
UqYnlZX3m4V1FHjgHiun4VIADTuyimVzJAJLu6vPpYGNP1UV2cnThMLxhCLTTHwU
qJ8RF8XoN9LxMT6krDWZDxr9+W+LIXygjJrpcAT9U+qVV1S7aPVGQYrfVP4NdjSp
kOXD/UKkl2gpg9sdB4FwL9/6PMZePLVpe61oPA7bv0+tV0E0a8oJ53a4xtt/ouc3
4Un+cFktvoxZl7xQVmW26LcXGUwH2S7sDCtMMPMmsEkShADF4ek1SXa1AcExKDda
1ayKW1zQW38ynNB/XD24C5oOL8kaKqVuxJuj/wir4Pod6844/28pd4pK5NgikYXf
EH+OzeJBZHgz7Iz//dZrkETQt+fq5W+MTzbyMxDL3ErXP+w1HAqVc0CPVRYA23QY
UiGHZIs2dtqXErEx92HOoutB6V0q1fh1ZFGLU3B0xmluPH5qktF6bEnYRSyliSbj
aJ1LbsNk6air4POZ4Yk3tO+iQTTlI+D6/FUHRJFH05GP0YSsgN0ubz8Y7bJdMCVy
sq0v5+2BVCGpnvDL1N4utyBofMNABQ16Q9177j68ulg2Pcw99ysCLi6DmqY4qR7a
FxGBN3GuESfuExBubyG/z9gehBnRhA/LoIe8TC3PX2kECJ/ix13DH+bO3fL6Bq7G
GBhoBpKlTEc4rq8xBckN3452pmSh41tTEHLTcG0eEhoKbyYfqGMS6XpJLZf/3+A4
jXM6yB1PatiGqoeCZE4wtytqF+bmnB5TfS4YuLtk7sZ4fzWf10HgubPSqVbyPvEF
Gdl56zxDQaYg2TnEBU/OuhV/dch7dwoIAb+2V4yysnvVXuReJoY9jjy/aOlT8UaS
IOfcDc4MeWYjhu3bldv8XHOcj0qBevQna392HxaXaZHlepPTVRT0fIFVqGJ5UUGR
7Is94mFWgk08+1qdZ3wgGcmmr7JOGs7+xW5yzQwm5bpkFbIQATuQbo60SXpuPVlC
N8XnB/V0+XBuKSxipYytLFQGkTGGaLlrYTJ2Nod/XEWtB+/mCYD62pWR8st+BJgL
qkNIG97foRufBwh0UILBeKB4lIYTgY15MnYP7+npYocrFwN5ulyI4BYQKAeVmLuv
ZpGrf3q1/J2nbVDEcQ4Kl8UCT6CgP37FdcaPbVBpvRhGa6UauTgn5y8DF3p0Jqou
1Q4fle9eHjvB2Okbf8ys5w+lypV0b96nOa/qVgV5gCk31UmLRRgdpiKn2zHfam7i
/AWP/PX+del9lj4WiVov+4i8TtMj/7Xj9MgVoAMfyHz55EDOhzCU7n1RyIfmnuQr
HWTKu7zRdJ9O+N70Z2hSNZK0gO41eHp6Cb5eXnhom/AgymeJMW44UdaWXowPF+Iw
aPRmiDOMLYMB2l53fposkMqI0tnWRkwUXqDX4tAIxqPjaQeFVyueMm7qsegx7v9q
z7qfZvHdcOPB/R+NYu7Rl8xaZqzasq21m7qhG9/VMHqlAwGIDtBpjTk5ngoGQ8CU
TnERA/1Alp4y/D57WNlKkM7ERKuCU30MoVphlGYhTxuWerjZQwXklB5Q3PgnEDgH
HxzNrbJM5iP84SqZRnEEvaBUVGN72Tekuyq/XWXlyaMuwq84p7EAWXx12QXkCts8
cxqrEK0YM526+7XeN/PKrLye347NhuxN5HjWIssnNAhdALYU10XWhmUNOLVPo+02
tSSUaG5TTQoqXLV3pAcFxhDZzC5O0vhbtftz3THIVSggcxWqAtAhRE8fSxDtU/n/
lY9GsTxaGo5f6MbFE4/D5dynX0xaLRs7nghFiYpjgDQufEeoS2oy7E0Hj79Zr5vY
TvAlKZFgnVQ9nJfPRWsHN2atCin9LRksLqdgJFlgEKAcEtk79zjFUYPfQkPSLS8T
Lo6I381gqB+Ldcj5q3uib3GlzsbXYYPvFIwhmL5UPr2Iqlk3CtvpeMnqREFk3pI+
N3nRH622Gg+gXTT9CzWPW7udhdclfC8185Xum3Jrx/KE9Ps4RKy5dN8YBW6Q90vi
cE2WXlO/u80M15aYAvBN96ZPfTLiCULLV+A1AAPP0XsFVGnh5txPBTPjUurot8EY
U9OVnqisKvtHmQ9BwRSS5mL5mY/84msDNUILocNX1xNgFSNuW2YdhTXL+CBsCfqP
81Qj5pFUSFD5+46K8d0NVhpOGEIKtzpTy6NfSxC90lB36xv9+nIy4UGKCVN2/qKr
PgGKkdvat7hhIzlL8HRkqAYXiKmQZOtY0+0OSHClAIm3xYfIPsKISssSYot70byV
wE1xsQqZ2vxd+saPzwjfbEMy2he9EzQHkmDlCn+L7RCwYBQIY5Qu2YELmIH/e9KE
EL5vJEBxkMG9QKZi8CWfB3PIb0kGA0p7nU8tls7QjpRETWYVx2P9P/Y4HgILWq79
rEg+bT+M1NpoiwuWw2YBr3e+TD51rXtpsRc9mo74eeHm+O+rQFjNgdqWgiavLIr3
wjT67LlDRQKRjwIBFzc8oCjkv8wSLjg3sB3C88k4juBW4rmFSoibOf0NtJd+NDll
FusLf4o731ilODFqQ2/Jao4Je0d3tDBFdgWJkcPWWF2eixw1AwWcu9DrtwinbX10
udEh1jQDXI0CeJu6EyTT64zB70mhsfwGFyOQtJEQtcsJ9H8xNzSjZzNUTTSUijfA
xqQijabX8HAaiv6rn1C4gGt2zPU+54eRHec/VHHAHmMyeYrtC/6gDvmMSj71ELRq
crROhz+lv06/8f3yLK7AN3E0i2iAdoSN5BfYgvEk0MMJoJmssP1hAR8SyXoZdu8q
t1G/t3LTv36AqDemNekvdTY59qKy8pWzzFGri0PhMlegiwIvYTqdgJrGs4DI9mR0
cEqA4VskuJiDpECUQ7aaA885uDJ6neZTqtm5jdjzyfT8jSVC0FtiMCr0jzPTuH2S
MjVe6Sw3CLwIRNH11GU74RhuSZbmM5gxdVHySqLmo6Zc5NR4kIgJgsYc7N+k4Xac
hyZdjNxhHitrwEOYK5ni+NAtY/9bTqg3KA6TZDO3gXINu0bUkl26GS3f7sMHjjtj
KDy7JASxHovkD+iS58GdfTFrBogQgOjCuOfRiCoLi1MUFuD7smXeQ8itcA6x4wxp
LLXQX1Eh9+S0jpq4YG+R2uG+nOP6zejDqActI+xSAmvtU9RGXV4apYfSYTnv9HyB
bXNC+2XrzwMKDfrteuBFbeF+FBpC1xiANqLXg4klRoz42Tvu6qF+g7pArsur/BlQ
s/0L0zySi3Azx3vdfJNjD8OmJtqH5LPGA2QorX3NwyrmvuZqCIPfs3Lusjn6MMlB
lrH7pV7qOv4sJShTipSZr1QGpHIxQaloqI6hAOPyb4t+jEOdU3f25okA8i/EgAME
huSGZxU5JC1cIWeRItW3dYm+LVAp4LjK7KMaBk77MCzmz4zPOb7yU+w7agpL1a1/
xXBigKE654WYFMtF92QuC4nctorAW8iUYuOxyT5lZtD7UlJLRXfuwgE5fRFxUSjg
OBdfBxE3Ll82OUnNd+7kvEzDmmcexx5FJeYcvCklQYyq+JWlby8J6QXuYCgYRcmg
SojQ6WJCBRjmabNbTYPyH8qw9Uf5ir3PbrCE8u+dlToDOq+rlTR6ZlvCoWJ5mZIa
dHKzylo7NM/BujpmCLDO+GdJE/5vG/Y0QgDm3IsI6ckzkRfvijmpUxjxY1UPNeEM
KU7/YW0hGuoeXuINA4MOvEya4RKFKelb7MDhf7c1981MaZXROnsLhDMebpnhRwKQ
lXqHV5KHl0TR61B4ci0/EXzXwLxuxb3eIBbM9TObEvo4q2LkOtiXHDAh/aslgjbv
v4CkBmoWzx2S4J5HqdkGvyzd18ymcxVfn6joyLTnUnQ2sUeD1ieLCHPqFw/9G8QM
FSpHQd7yjpD3ULWkAe4cW7+DgT8cjv7BIL0Evjnj7GmpiUJD1SboN8kIxw8O/EL5
fs2QoFCvRki45S/+M0hx7OVY0IOGxrwqkz3HXC8r4WuxuptGyp6W6ryXo4uP5DWC
qAZiEQrD9qpNTrLlvpuclE15AiHODIzHl6qgb6sBpXaaTId/wlVjfcqx9prQ+EzB
9B0nt8aE2jw8F/LUnLiEmVpAF7DGy66VkEEHdAMvjsFJq/S6t9hnE+HR58PU9SYM
3cs4jSEUCxxN/z+RqvU4FRkhYaEF72d5Mfrkh+C9hejE8oycylyr4Js4J7YjFahf
xZzv5OMRIZzg6/GWRbAsLrVDln3cFjqMOL14ntKsWrGAWhJa4wVI1EHjUDr2Q5DC
+IoGdjqKlaGwOQVEz61WPk4EAHp7JU5/mPSuyfSl3gy4cX9/QlJ0rbXRcypQfqpY
8jnLpXErN4hc+NyULj2e9dHzL+jXar3IlP7L0pu6VZfdEXVLdtc0E2KBREz0ZBrf
sLTiRxQAMel/PsEOQPTWCO5zoD3DboTwRXfv2VH71qs56EmuzXTqTQ514pEYgqfY
J4OgHBN6MQW3+/LiMlOv/9BvZ4ehCA/6c++OSZh1j+zV3R/8wrWvZuTjBdOo0z3e
MCSQae2cTtZKhO78ss4vpiVmfPHSoSFn57eMx1uExBXR/XucbU7bZ0wy74KhXNdA
lI4UbzyYMX0q73g1JVfY8pF7twwKhF+eAgGtHA+I9L6PNClkoDluml4cxMGbUBrD
NmipXgDcti/ceqwgPhaSJ1IEOTEluARr2/SBShIYPmRyWWjRA44QyenxngQ4C9eZ
8xhF7OwqarDwzOQCh6YekBhK6hhFux28wwJPOyhbURGPO0IEDiVXNQHlkyWnop3w
S2rycESqxjBKff7tn7ShkUjheFiP+oS4ZGy4uYp1RAPqerzMGEF66Qe9/ebpnLXz
b1OSsxWfuSW9UR14wAOXoHSEpGtontzOoQAxka216cvv5CW+LMS4KFZR6L6AQvgY
tCSLyFe0uYuv5AEtTl3aH1HgjAm+qexYahyXk1hrl6YqcrqDZnGtRyBA+8VzxxlQ
GcJxL8Ryby7H0TIUB8YOZdtuuWat+EAoHGTrO6npW058H7eDQMT3xfcl7PZEX/As
jw6+zRcfK1QE7uQkfL6BlGdUPfwFf/MbllZoQRn8fAKDuBcGVSAoUM5IbYdxfRVd
Lx9vPTpdIlJ9E7zu4kvel8Y0D6Skwr0GRiCCh0T3CVp/UcyRn+9/g1kwhx0EGLKz
n227SjL4fMMWaePrkbKSssrWqFMWrZR+/7N9fBlUcUpqU3OzkWkHpWAJmwNbSmfw
eZpI6i14wprtWizSDq7MdXZ3mm3LKtQwyrX5Q9yW7zfTdNbgJKlJjK6CD5X856dd
HNnLGt90+y5ymy8zVCsLqyDp+DQLsDMdm/sy7UzcPt9CBGOdA4i9BHKb2cYWAOBv
dDOwO+YpcrpysENo5CNmQbJ7fRmY7lIlKqPxf6ye7pqRs0gSPbdVw4gvREvJDLvM
bL+f1nrEGwL2w0LO55seh0FIqbXDAuWe+TwpQIyS7mCKU5bah4CdW529qEHcsN+/
WPzYwsXoikTHGjTHhQCJWQT+FKxjUJLtF08F6Qmgazk7rIrtw2r2l8QeAexSrzPs
e0UdjbIBub9hlDuIdlLIoxAx8CaU7vZ9T7TGAwsO0eIrawgfYeOBpar/nhEfOb8W
WBm3EgzRlJtsVqKwZ6ZB6j1MDd8VB2/pe9UyhuzNc6ZcyW1RRSFv0VpPZS7swX+j
ewvkIxz71eey1gIg9JKQqg6UFDC1Acl6fEF5y7AVrySguNnVZK6IA+SD9PcVPzhm
DR1GpXi8PZy4mxh1wSRnSYwk8X4K3izgEWSzZV7drgGW7FRSkWQR4H0qBlxrKaiY
+licUTke+CJ6morSsm5VhQl6rUif8of8ik+8zrEnnQOhW6N+mPHvZW8knPVJxRGU
1Vukqd2PslVU4uLfZBzsldBqsjR0Tvmtrp+QH6q1F1h8+XoHln8qgD5b4d3Nqtzs
p8NW3/7Yzm9d/Yt8gx1QFQgLj2lAo1w0huRlwS6cZ3mtFoYy2poWTDvGTIOt3A15
a3ZibdmXdrCL69cUhP3/dUFw60KkezqV9dV4LrDGURzaP8OUpLTcAs5ar3bExe1Q
6WqYOv6TpxOxUpcdTg5MkAf0wAyDqpBBEZwVey7NVZzEVawVwjn+qPRiZN872XBQ
RCU+FrMphfclNf1kwMKmWEOcHu7jccNIhavdL4pXj/boQp2y7kDIQoP95DQAwNW4
NllgJUmFhsJ+oRB5RdsCP9tGLjQoAyXbVpGgfh+6scsnU4qByb/wwATmOFu9lpqA
8bF/5nXWHIl2vu8571ace4tt/pTVyjVxFnisDh9xItpafm1fV/FkrTGbwSXp8X2v
YZhYTK94/w8RUxDs6QBCfFFFciD1CL5vDsnK0HPoETWt/m56wl5rWSJQ+rrp6+wc
IMr81pT6nvIXO1vUfU9Nl1SwNWEohjaQyxkzyRT4HRIl+dJicXn6SH/1XCnXh/PZ
vlcisodXaeMsv8mt/6ttFedAZFkG+QXPBcolyrYErhID2Ex6+aJc1lw5dMy9cl84
XopxXCKPFimAI+UJEkeN/g6axoACi8Mxe7qAej0J4L8skvVJ6LurUBuwlWnWbJWC
GtnS6GirrUzRkd0TOZuTEuOUWWLEpfKErMtA+5eX8ifwvDcFHfczGlJC6xUE5ztu
gJcSV2DwBD+dmuJaxwg0RBQWZTKd0c5LPmlu1qZg7gZiihxJY8+cZfTnAUi1i6cv
GmpO9fmBPrLdk99CW+8VXiojyRDJvMVH0eTAReiHRSnwU2wyeWWBdUv09xiGDjEt
s6ImvYvQzty2IfM0N8bsdYDHDQ5zVkzPJAPQFwa7C4JkuKj5+5vjUs2cP9T7Th2s
VXTgoJhtDn/6qHDPwSodPv7Pc8YU5455RtdjduJiCGgS0fHhigyKsuGrEk5pBu7O
gUJ0M/pmQMvJshtdN4w1/hmMf3dXkLX2uhH/EAWwZc1Hu5gYwG0oTC29WX06SMGZ
zirdsv2goBxUNMUMFA9v/2VVAGV5b6A53f5LzxMRkSMNBcSJliBDXa/+YKBtmYek
gk/gB6mCDN5p3dK4bLBzR/SjO8MOii8//cjX1dwPD9Qn1yLGUrULBc46qArXnb9k
O0puNOBFZReZiZC44EpPvoTjBoHyp3hrzdcdbiDpGdwCYKlKF7P5vafOAcENIYcL
tiS1SYf69Xs1bTi+XeLwebcgybDpUY/AT807uTH9U25Zgo1kQBsHti6QiW8odAnp
R0r2Vh4yaUDqyzMWRu0JyRKc5RPu4cLa+gWTfDRip+1utMwzFEBWUGaJ38fHQ5R6
UIRS8neUg+YVcu8lCzLuSU6ZxUpoEIwWDdgw3kfbLmdgjJGF3sLyKhc49StZk7d6
JfSeooFceP64xzkE2cny85Q8M61htXR1dIT3P2oO9dnk/wfZYzYusXMpmP6E/Nrv
ar8FS9H5X31y/0POsKKiVpKl2jYGKZVF/YKhya24lonE9UVEyo7CLazsJVMZkdqT
dt5ScDyJJVNykk9NzFvZMiSHh57wAa6FHFcw8tIFOkTChvqhKLEun6pQrSnvo5ot
gfBb1UJ/cxd6oP+LkpSSPdEAsu3KOhgiUlYOiBcEFv2AzSEQj76O7bvdW8TVtB1v
usrIdsKKaG+lRQO2Q/oRkAwr1ZU5+/E3nslqr6FjArKA9bTVqHm0d77huFvbq2us
YT2lJY/zy1SIw/pwPheno0Sr55++TGQKEap04XwwQG52DK/3ztZuX0J7hIPYNCPC
NtZvJlSONXucga9w9RmNFPwYvS5zEiYoAtLDWKmRPjyn6QZzOG8M0lOZRZoNgE5U
UG/d3a+C6PgrBNFB+8LJ1mD0Zqaz6EnEaJd16SGWJerHg+laiLHZ9wvjaZX+b+vW
BNl8LP1l8KRzUCzbJTk/X/tl95AXhupYXV/G2GjagXrhI8gJa+rnr4/NFDGU5u84
vMG16Bzz0nOKmjrypqp58pRi6dEWVrQwEmE0sdrCvXo/W1WQ9sRjX2wTMsER+T8k
XViMN2s9PPciaeRjhu8kSKyLT5V1jmmqTniqBzP9L0CE5mroCfaTaHUI8rXli+mc
C3nZZfVkG41w3LoIx+twEmDkWhQCjGcuCMLouA1H+QjnUqZaKwG6O+82sxWaU1Mz
/DU+wM919CZlKOzLtqZDSCGhIwAjxhu6u+nLUb1d4CVAf+7ZPOAyruQ3D5BtLx/m
BvEXHkXY47E7FbzEOpheQyit5tHMzlQ4XYIlrF6X9ydRk65JPDIrF7I6wclGAHuq
g0R6Yw/dwzixqaTso4gl+XwIVkIEwoT0owNri5hC3BqJf7uGkkhXzLRslhOgW3R3
a8UJ+H+knfCFMX/NXlv5AS8F+SEiGaEn3LWPB8mKRk6xFUgyVrdNiDJqIU+ntJeA
pFB9/hTQaglIzBd0LHKjTaajohYaufx3hdwCgxM5defQW5CJSyngTqtWp6JYW1Mm
P8BdPG/nDIpyqHX+Ssy9ewL6onO5LTvkPyfWr9eoMSJFdrZSsgbyjK8NnLmXLmDm
XOSknHtl+QF0FQj3vyvTb6QEovpXoAUMda5KOh2Y3q3pBxJ/pMeR6haiBH5VX5bX
XCj22DyQCk0IcoJpBqSNLnoF8zLmFkEQP6QtIl471zg5Ug/biswxX3vulAz6Lahi
Lt/vorCD0lacW8UEBdXS6VS12CmT4p+KVAhnFQY9S0t8JhzI68A6neT0ssC1uVRr
QLFg7DO2PCRa7T2aUgyPM2bzWRkx32yvNGEtaC7f0dGkvjWziGfUeLCGR+ku1Pay
ePaBQRP82uhIDjgnNQ3lbOIrg0jqgJW1IFtzNTxesP1cVTaIqRijKuwUuRTmpfpu
NxPpDH5+/pGnAZ/b4DbXRn8Jts7jkhqwpx/NAfx4fJaUUjaP4F8E7iZpx+OtkNs5
gwXcf/eFX47F8ioVjIasl0WnipdbtNGEun3xbtwpGiIno5ddn7jeOXPNvO14r5L2
hfH4xBpuJEmQ+PHJjss+rAFdZ/yAVk5iJWCSi58Id1ETyHd2Sne829JmsEXvu5nk
z/nR1v4s8q49WxCBk1yrGb5SAylfszVpt/8N48GXqroymYD9y0wQZEqjK4g3p1Lq
UYy5kgGcfrRXutEIk33fq2B1PHTKrHvy1U81NrNMQFYfOpYZ5mm19oJnpbSqhMqc
HjeNJIOIpn61jRWoI/vM6513idddjjyJxnj6VDUyR3h62RMQqvtCYBQgk/7bJ/np
NMHyInuy0jK9kV0FcpiUGrFRUJLZkVQldMFenAO+Uxk42LGSyKg5YcmdoW8P+Pta
m30eRBCbylHOCSMCOQYXzjpYE8KbplW9ApDnQ5jeRItP+J51Yx5LYv1qmfalslLp
eG49oidlwHIneq5XuhbBHcwEv0iB/ma1b4raThVBbEz5SnTDsGQWU/hnHI6Fn0lR
Pm9AlyMkimOHRcoZwVRIGxUPk6eikpHUxW4KjDSNb6s3afbj4kK3SFfc21H3Z8a5
GRhQJXd/TrdyOuLvAAT/OqL/kWldsJ4OrGcW5K2bSz8UzC6kA2un/DPYhhSVsVx+
7acsruq9lTpq+Upzem9W5obh8wPsEy7p/uLry14aoZ8LHOadWTekzxD2ZV3e7W8B
Rg8vZbN2SIX5i7aKf7Xt0F2rYd+RKXY+qr082wzaF5/NM9b+V0Rz0++YscjeSaz2
k27WorkxV8uSuCOX/5D6kv363Ejby504GVFGYxaMEv7vjOvkXSTaOIG95azeVsVw
zbwFuwBreNPqJos7dBETfavK3aTkVs//RV7b+VlwFcRvUDZ/XVwRr8SwJPbV4KiH
c9Gm+A445nx7kJHm2jTQPt3L14wYVlS03Qb08ivf8zLmBcL5+AF4Nwz9wxtI3FjE
l4MtohbewBOj5NrAQuSag1kWV1MiSRXRa3ygkff5kcwodicBV/vw7AcspKnLkvIK
TeyubpYtX/QRFFUO6XPhfej9R19K9d7KAKk5lsVVU4tE7+nCBDorZSzXJRN0EBVG
8U57KBfJWxUZlHFPEY7O7+czm6iU9qBcEK2ySpVvbe1NLXYNPeoNTGvU7UiXXFuI
K8tZ83WL3WSZNU8jUtkduAtElF+A/plcboGzyVyVpvuORV0+lEfKF49HI0xltmnR
SNTnV1Lm/OH2WOMjh59uosMwY/LW+uzXN/bzwXKPN9Y7iqrXXLqhRtSfPyf1uCtT
U9mjblsCdIU19JA0cmE2TQupK1tubKtD8vywJCOm6eqvUaG+6rqhWqpon0vPO4so
VM9bKJJfSy1PzZ3Az6MdHtM7zWZE1Y3zNEpcnwL0/dlNOl+BkTyTgtCuy0cNSLXT
Br2SYCkpEDdSB0ugqJcsCVOnWja6fXGBTuCPnuoBPl1ijgHJBfRSJeVRswN/q+1F
Fye37cMNyk52fpwZEg6lKBuw/cHoPpuWPj1N1zasBUs7nwxHmZWA9ceqGIHmFHlC
lnNGcrNSCSXVOsQ71uZTUydS6O4QTPjO1G/w4nzeabT10npi+vJ1839Ys1cC8MDF
dKd1WuyGlvATKQQE4N5PKbK1mGw/c9FqirE4KlAF3urUbSJ7X0ikAYD5let/ELtL
GtxvNSPScDKmla/q49f3auUahuyouMz/hYKuDjRvWZPdal+WrlrkRVfzvNxFJIXR
F+bsBhK26AoFwZOtZCZJYnaouJeXhADsd0aLpLfbOqka2MUZD7i8LMnM4fsxsKT3
9+6FXjpCAky9o9cOQoU5eE2JwlFEECBBkIiRVkpnevPa4KEd+ERxy/8fmCbEe4qy
V/oBAu42r//1B97gVDm7iAqFzXK2yfEmbP2vfgDKhEQQqOamp4NpAMmtlN6dCCiK
Zs1ArYTEBW/XE62zPs49iw7IkVmyyyR97dcCU1E9vsC4RJrLDILZuGnhHiqrY16l
jVT27JZCZ/cjGXZlXO1SfGrkVYFIgDthchIq4bMfrYuhT1+xuhV/ymepHQLgCVsU
V6KpwS1kcz6VuR0bTA/CCzmx1KD+Re7hh97Ge7LnqmvPADflN12ncPpwvmLoJJFn
c5v9breG+staatw+QQunqYbUyaAvIpkQ2swQuIR8M+FN+rukzNUVbCtQR/MyyUAp
RiF63R8FtF4kuzYe5rI9yBy4Y0VPpf2mXgyU5jPc6r1COCsnnCsa6X8s9GO05edd
CEPe3vNpbreIfmNvputVQ6t8Yut5C9qkIqjHRE4svpZ8qSbTQacTGOcsaGWRwnxo
HIxvAkWjb9sq4Cb7So4GRJJAfj/o5sjImdPsiuBQ+j6es+7ZeJa2sbxCdlCjaGZJ
YoQFgDuFhDRei/Kn7Z8LelyvtiZZWZb5cPBg2BXnlAXWgiB+kWjG/xYjp1nk8z0F
dRE7UNhPVtR3SA6m1KMmUciTKX2gaXZEr1gYQxHO5zI=
`protect END_PROTECTED
