`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Peg0yChHErJ5jXkZcyaqct5xqgxQ53FoR0nHS1PSuZhtH5XIWXOx2jW+/sfs5AZC
K6tHe9c+cohHMdC3oQmEDXcFk7h0kMWy8A2GArloRtgvuidJLj7jwk3Fw8lZ8ymv
LahesuVazxZGce0fH6Fot2aeZr+oUhlcFp9cQHK1MXs3OcdS7mKzHaqhxazRLHAl
giDV0VfEmOTGyEjHc060uIAU6yHRSg15ubKUO29OiBnTIQqULze1us0lCkEdb0KW
LXNMu2xwVqePXuNLwJpoP/QqiPBC7oHMLgZL8kRbaWvOpd3thi1biYrBFvq5lLyQ
p3Wa9Mwjx2wWrCECGQdmTwStfyRzDd0E7uEWi6a/JAyjLRQ9/byxslzyaWg8F7I3
TDaRHykeeg6vG4Ay10KdpAA1dxZtaZJ881PW+yK0KDCg9QXf2KAGMIHlIb8LIbUD
7P2p8O1FsflyXipr8AJ6D9oGwOTCJLRKZejZjgh4Hv/3/zCwdyUzaWHvTEnABtgM
8/2fHb06uELFTHA/wktN/qib/zkDnyo9hquiIjuRAOdsExfppYgv3KLCcq45vIAj
cwoDMNYH+1MsXXcDEqJUffBwUtoFihDw1pmUJe02XUal/AT9RQM5ddpTRJKFewfP
ETWgJIUxw3HZYfi7aFQGMWtGoWfHWuDu/yG8NRXrwLcbPuKJS8D7IB4NiSUdDvAE
5wThT/ktq/N3AuFLBnxZKWEU40vcISNRjwBuKenVolTihqYD+eX/DZcgEazTEvac
XQIPWs26gRkDQG3WQu1BPVkzbHw/QcmnlZ90J/xNjTS8K61XtB2wTAyFWkHkrW/R
W0FPpj07H/iGPuw3nqH2naOkWNEXZIm8ICGMDeMBm4Zysa2P5UdlY0O4wV91XY8b
j5LlWuCCejxIatZyzq4wU3/p9y2RHS45Al/qPbFLtqCG3IJMYYJ0e85MUC1LyU0x
TNu0dYO5Q5NUAS6lckbiJFGuv0W9G+5e7nvjI+3t4RYKrCZ7puTjwOvJOMQYtvH1
ICYiIUiHT9kOi5Zm8gY80J31IbnI507bG6gHdbB6Msc=
`protect END_PROTECTED
