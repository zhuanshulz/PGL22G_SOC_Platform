`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2o2/HOyZagcfg43S5eyE4dujyBL/08MN1hZ4tBW9sydYjiOl5MIOrc2PReMZjD4W
OQ3FIiYuE670/rd886RyJzR2v0FGuDLAOsmIJp9ftOzAcI70xATST2CnB8Py+KUJ
MJUtKOIaPQ2ozyagonC5wB11pTYqx8dOJ9C/H2uWJhh5CvbSmcahtRSY5+NvS/JI
LwFIS+CsJ+mNvU2KK6kNa+Anj7gVMvEK4tXVop7fPa0QHiQp010J3+1TYJ+bjCQQ
66SiCQW9LEP5Rt/EDPqpHAwILiv+nPtQdXbTckueEc7pWhkivXaWgWLUtXLGB3sj
sRHQf7Gy8stuL7jAw5JjmOS1UkDGbl1s09yz8hrQlFc5Y7wqUnxZZRtJJbGuAkzZ
OIhhWIZpLbHgaiuCuJHXnQ==
`protect END_PROTECTED
