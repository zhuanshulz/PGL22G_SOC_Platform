`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O/+pfKI5ip3N+OlQr17n2KrkbveGNIO6Y3Ub8l/Q0MSllVb+rvOO+FYSGrdmrbzy
ZEnfP1OdRdmiLh/NfT+ig/fVdNXhwtPVlErxx1bgk06AOeilfdIS7GMUKW07SiMU
BEMhpqf7LzgTSEddrNUQrH0y1WOePgSCQmqVcPoKqSY/rDvoA3CIz+viHCqoqX1k
+AkXtfG97XVQEq4+8xvWnqHKxI5mYRCnb5ANQMEQhnqnysc+nsm7TJ8EfG7cPhqJ
/UyyDF27NUqnx4swe3vCsQ==
`protect END_PROTECTED
