`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hOpFLeBDI0mRBL97+1C/9uZx+gW8oOrQgejkP/kZTTAy38j0wxJzJPhAEF9k5+VI
xmJ+JTW1yfo7yCtUGplguofMHWht31qoVJCXEBaeSu0IJhiDbo0oigBJGwX1ou1O
bWIpr29cj3gioF+u2OGDgGnAkkHwCdHSShEipFoYV0OIrhaJgh+0T9JJr3oWIO0G
wkQ7YQn0suhMSXl1clkWbRRjleTUygQdr05VJiO+iSSMycfgxK/Ym08UkbiWPcWl
2uDhPQRgmqdPBq1CFjWMyV0eGnUxG3spMskN/gjK9KlX/s2a/hsMKReMYgrkLd2v
R47cTe0AhjqBxBQ4Dz3cxg7DWVUN/qgWSLClFg5LTxaaKIKAMjF9/mEdKoOM1s2o
WOWMXYq0MqZygr7QOB9CEdlnOvbFJdr2m8vqFf4xCfi5kOHiVTxUEci/Y25oXcRO
sUKR7fe587/d5lXseDtzQbmp7uujDJod/Wrygdn+sNsJFVRgfGv6M/igounzhqLb
wct9u7EJl08cywwhOAVJiLF17BOGLV+k07dn9z8ARYTGu5GNmC4KxK8/3Afg+HTv
MYnV1JWmd0fGhnUTQQObNoa/iiUimM8TLnC8Z0RW1grkiWudL01AgtUg7QXjP11S
bit17MXH2LGJNqpXt+wbLYAED3KZiZTi3pf4xTbv3i6sp7PoN67a2WziE4axyGEq
`protect END_PROTECTED
