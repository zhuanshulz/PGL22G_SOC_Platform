`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LPN6EqujZe//2AtL1pid7uR1J9cbx+Fx7YKn2TefZPopAJAK66rvVjZocWbOZz10
s90PAIFzArsSrjzbPNMNJoIFoRZYjaA4KfSGXgoyZCZEVRFmp/2AT3AKova0EP5K
u+XrrcsW679kE2d/6PHGeoiTtny32gsei30sNYaPdqigKA6kZ8mC3u5I2iPE3Vhn
PlSAfk+5WRfPCWuwSAKmUgAe6BN1nYkxYr9ZNxG+7L7cjJ4E+Pv9Ni7iXbOe/6cU
zb+wzcB8UDZxDouqOly2RwSbhD0qK30G0NCgBwwJbKeb4C0dsKGD4KrPobLV/aOT
hjgN0Wr7cp4n9Yq4G+XWSeeRKsIGRXOvxg+u7mWH5CVz/40aX2LBjsOVAN6zfKMt
1JPZkdMtuAKe0X2Hs1tCxu0TEC+VeZq5QqZwCTzfC70EaC4B2mTT+Zi3WfKx27kH
fC+HxbJuX07BbyC8ZaaKOScr3EJ7w65uYy4apUK93w2xZDZOZQYe2Ti1LZRYXrQy
OYAxyvgFvDH3J4QpgxONPIKze0pAi4YWGvknWnPNB8rDX1pyO+qRKe5EbejPZPjX
fEqhIs+Ps70IxgoCk3N61Up1smLzk9pKNdVMjUzQnIu0INGCHsarRi35GKOgZGgr
sX64au8C8ujDV0sgyvHd4DMukgO62vtWdgmp8AWiK6sTVqiO/MlKZvTluYmhITGe
8NvxxiJbIdCCn2zbtTB6ZZC9Bj8v3mZe+kgqDxXxFWhMqXwPBoJ9Msgkk12LQZMx
fSM7inL3FT1Sf6xfKRNrdQ==
`protect END_PROTECTED
