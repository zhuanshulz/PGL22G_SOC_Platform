library verilog;
use verilog.vl_types.all;
entity GTP_HSSTLP_PLL is
    generic(
        TX_SYNCK_PD     : integer := 0;
        PMA_PLL_REG_REFCLK_TERM_IMP_CTRL: string  := "TRUE";
        PMA_PLL_REG_BG_TRIM: integer := 2;
        PMA_PLL_REG_IBUP_A1: integer := 262143;
        PMA_PLL_REG_IBUP_A2: integer := 0;
        PMA_PLL_REG_IBUP_PD: integer := 0;
        PMA_PLL_REG_V2I_BIAS_SEL: string  := "FALSE";
        PMA_PLL_REG_V2I_EN: string  := "TRUE";
        PMA_PLL_REG_V2I_TB_SEL: integer := 0;
        PMA_PLL_REG_V2I_RCALTEST_PD: string  := "FALSE";
        PMA_PLL_REG_RES_CAL_TEST: integer := 0;
        PMA_RES_CAL_DIV : integer := 0;
        PMA_RES_CAL_CLK_SEL: string  := "FALSE";
        PMA_PLL_REG_PLL_PFDDELAY_EN: string  := "TRUE";
        PMA_PLL_REG_PFDDELAYSEL: integer := 1;
        PMA_PLL_REG_PLL_VCTRL_SET: integer := 0;
        PMA_PLL_REG_READY_OR_LOCK: string  := "FALSE";
        PMA_PLL_REG_PLL_CP: integer := 31;
        PMA_PLL_REG_PLL_REFDIV: integer := 16;
        PMA_PLL_REG_PLL_LOCKDET_EN: string  := "FALSE";
        PMA_PLL_REG_PLL_READY: string  := "FALSE";
        PMA_PLL_REG_PLL_READY_OW: string  := "FALSE";
        PMA_PLL_REG_PLL_FBDIV: integer := 36;
        PMA_PLL_REG_LPF_RES: integer := 1;
        PMA_PLL_REG_JTAG_OE: string  := "FALSE";
        PMA_PLL_REG_JTAG_VHYSTSEL: integer := 0;
        PMA_PLL_REG_PLL_LOCKDET_EN_OW: string  := "FALSE";
        PMA_PLL_REG_PLL_LOCKDET_FBCT: integer := 7;
        PMA_PLL_REG_PLL_LOCKDET_ITER: integer := 3;
        PMA_PLL_REG_PLL_LOCKDET_MODE: string  := "FALSE";
        PMA_PLL_REG_PLL_LOCKDET_LOCKCT: integer := 4;
        PMA_PLL_REG_PLL_LOCKDET_REFCT: integer := 7;
        PMA_PLL_REG_PLL_LOCKDET_RESET_N: string  := "TRUE";
        PMA_PLL_REG_PLL_LOCKDET_RESET_N_OW: string  := "FALSE";
        PMA_PLL_REG_PLL_LOCKED: string  := "FALSE";
        PMA_PLL_REG_PLL_LOCKED_OW: string  := "FALSE";
        PMA_PLL_REG_PLL_LOCKED_STICKY_CLEAR: string  := "FALSE";
        PMA_PLL_REG_PLL_UNLOCKED: string  := "FALSE";
        PMA_PLL_REG_PLL_UNLOCKDET_ITER: integer := 2;
        PMA_PLL_REG_PLL_UNLOCKED_OW: string  := "FALSE";
        PMA_PLL_REG_PLL_UNLOCKED_STICKY_CLEAR: string  := "FALSE";
        PMA_PLL_REG_I_CTRL_MAX: integer := 63;
        PMA_PLL_REG_REFCLK_TEST_EN: string  := "FALSE";
        PMA_PLL_REG_RESCAL_EN: string  := "FALSE";
        PMA_PLL_REG_I_CTRL_MIN: integer := 0;
        PMA_PLL_REG_RESCAL_DONE_OW: string  := "FALSE";
        PMA_PLL_REG_RESCAL_DONE_VAL: string  := "FALSE";
        PMA_PLL_REG_RESCAL_I_CODE: integer := 46;
        PMA_PLL_REG_RESCAL_I_CODE_OW: string  := "FALSE";
        PMA_PLL_REG_RESCAL_I_CODE_PMA: string  := "FALSE";
        PMA_PLL_REG_RESCAL_I_CODE_VAL: integer := 46;
        PMA_PLL_REG_RESCAL_INT_R_SMALL_OW: string  := "FALSE";
        PMA_PLL_REG_RESCAL_INT_R_SMALL_VAL: string  := "FALSE";
        PMA_PLL_REG_RESCAL_ITER_VALID_SEL: integer := 0;
        PMA_PLL_REG_RESCAL_RESET_N_OW: string  := "FALSE";
        PMA_PLL_REG_RESCAL_RST_N_VAL: string  := "FALSE";
        PMA_PLL_REG_RESCAL_WAIT_SEL: string  := "TRUE";
        PMA_PLL_REFCLK2LANE_PD_L: string  := "FALSE";
        PMA_PLL_REFCLK2LANE_PD_R: string  := "FALSE";
        PMA_PLL_REG_LOCKDET_REPEAT: string  := "FALSE";
        PMA_PLL_REG_NOFBCLK_STICKY_CLEAR: string  := "FALSE";
        PMA_PLL_REG_NOREFCLK_STICKY_CLEAR: string  := "FALSE";
        PMA_PLL_REG_TEST_SEL: integer := 0;
        PMA_PLL_REG_TEST_V_EN: string  := "FALSE";
        PMA_PLL_REG_TEST_SIG_HALF_EN: string  := "FALSE";
        PMA_PLL_REG_REFCLK_PAD_SEL: string  := "FALSE";
        PARM_PLL_POWERUP: string  := "OFF"
    );
    port(
        P_CFG_READY_PLL : out    vl_logic;
        P_CFG_RDATA_PLL : out    vl_logic_vector(7 downto 0);
        P_CFG_INT_PLL   : out    vl_logic;
        P_RESCAL_I_CODE_O: out    vl_logic_vector(5 downto 0);
        P_REFCK2CORE    : out    vl_logic;
        P_PLL_READY     : out    vl_logic;
        PLL_CLK0        : out    vl_logic;
        PLL_CLK90       : out    vl_logic;
        PLL_CLK180      : out    vl_logic;
        PLL_CLK270      : out    vl_logic;
        SYNC_PLL        : out    vl_logic;
        RATE_CHANGE_PLL : out    vl_logic;
        PLL_PD_O        : out    vl_logic;
        PLL_RST_O       : out    vl_logic;
        PMA_PLL_READY_O : out    vl_logic;
        PLL_REFCLK_LANE_L: out    vl_logic;
        P_CFG_RST_PLL   : in     vl_logic;
        P_CFG_CLK_PLL   : in     vl_logic;
        P_CFG_PSEL_PLL  : in     vl_logic;
        P_CFG_ENABLE_PLL: in     vl_logic;
        P_CFG_WRITE_PLL : in     vl_logic;
        P_CFG_ADDR_PLL  : in     vl_logic_vector(11 downto 0);
        P_CFG_WDATA_PLL : in     vl_logic_vector(7 downto 0);
        P_RESCAL_RST_I  : in     vl_logic;
        P_RESCAL_I_CODE_I: in     vl_logic_vector(5 downto 0);
        P_PLL_LOCKDET_RST_I: in     vl_logic;
        P_PLL_REF_CLK   : in     vl_logic;
        P_PLL_RST       : in     vl_logic;
        P_PLLPOWERDOWN  : in     vl_logic;
        P_LANE_SYNC     : in     vl_logic;
        P_RATE_CHANGE_TCLK_ON: in     vl_logic;
        REFCLK_CML_N    : in     vl_logic;
        REFCLK_CML_P    : in     vl_logic;
        TXPCLK_PLL_SELECTED: in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of TX_SYNCK_PD : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL_REG_REFCLK_TERM_IMP_CTRL : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL_REG_BG_TRIM : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL_REG_IBUP_A1 : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL_REG_IBUP_A2 : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL_REG_IBUP_PD : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL_REG_V2I_BIAS_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL_REG_V2I_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL_REG_V2I_TB_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL_REG_V2I_RCALTEST_PD : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL_REG_RES_CAL_TEST : constant is 2;
    attribute mti_svvh_generic_type of PMA_RES_CAL_DIV : constant is 2;
    attribute mti_svvh_generic_type of PMA_RES_CAL_CLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL_REG_PLL_PFDDELAY_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL_REG_PFDDELAYSEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL_REG_PLL_VCTRL_SET : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL_REG_READY_OR_LOCK : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL_REG_PLL_CP : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL_REG_PLL_REFDIV : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL_REG_PLL_LOCKDET_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL_REG_PLL_READY : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL_REG_PLL_READY_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL_REG_PLL_FBDIV : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL_REG_LPF_RES : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL_REG_JTAG_OE : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL_REG_JTAG_VHYSTSEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL_REG_PLL_LOCKDET_EN_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL_REG_PLL_LOCKDET_FBCT : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL_REG_PLL_LOCKDET_ITER : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL_REG_PLL_LOCKDET_MODE : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL_REG_PLL_LOCKDET_LOCKCT : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL_REG_PLL_LOCKDET_REFCT : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL_REG_PLL_LOCKDET_RESET_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL_REG_PLL_LOCKDET_RESET_N_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL_REG_PLL_LOCKED : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL_REG_PLL_LOCKED_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL_REG_PLL_LOCKED_STICKY_CLEAR : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL_REG_PLL_UNLOCKED : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL_REG_PLL_UNLOCKDET_ITER : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL_REG_PLL_UNLOCKED_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL_REG_PLL_UNLOCKED_STICKY_CLEAR : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL_REG_I_CTRL_MAX : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL_REG_REFCLK_TEST_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL_REG_RESCAL_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL_REG_I_CTRL_MIN : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL_REG_RESCAL_DONE_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL_REG_RESCAL_DONE_VAL : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL_REG_RESCAL_I_CODE : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL_REG_RESCAL_I_CODE_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL_REG_RESCAL_I_CODE_PMA : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL_REG_RESCAL_I_CODE_VAL : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL_REG_RESCAL_INT_R_SMALL_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL_REG_RESCAL_INT_R_SMALL_VAL : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL_REG_RESCAL_ITER_VALID_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL_REG_RESCAL_RESET_N_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL_REG_RESCAL_RST_N_VAL : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL_REG_RESCAL_WAIT_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL_REFCLK2LANE_PD_L : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL_REFCLK2LANE_PD_R : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL_REG_LOCKDET_REPEAT : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL_REG_NOFBCLK_STICKY_CLEAR : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL_REG_NOREFCLK_STICKY_CLEAR : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL_REG_TEST_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL_REG_TEST_V_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL_REG_TEST_SIG_HALF_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL_REG_REFCLK_PAD_SEL : constant is 1;
    attribute mti_svvh_generic_type of PARM_PLL_POWERUP : constant is 1;
end GTP_HSSTLP_PLL;
