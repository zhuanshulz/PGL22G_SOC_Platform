`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WhXWtB8ubymTkHm4rIcripdDPLKaBLCakhUcJP1oUszJnhrVRjKt11funW87qdOI
OU1UEyxptG4hzQgf3/HsOjCKgb9p5s38kIHpTgc6It58mb7ROwMJ4oU/Mb/aqekU
yX5Q1lq9+l/m5Pr+L0cN0q9NDgtFmpnIHC+q9BVWXX/MdathPQZ2lUQW1RC/WIcB
IwCcU5RIRYV5HBot6tllzb9aE7HGTuuxZn2YW5LVHQKiywaGrj8P/HXi3NBKUdUY
pn3EM0hzNa6EEfkQMFVL3JMrtE2KAA6GPw85pID7M7H0yZlO49z3TYCs2gPNpW7b
H1VT/wJYNrWfeTNaJQTARlcVpRDBGS7k3DygLMsEZeQrtlBPyPTnmC6eHVdORJWo
oJHTB2HP1CB4kyFxu2p4GzpHMAemVkOd/7/sY1Grp6aQ3q7Bmj6YAppUnZXlkQYw
b0Tu3CujvyHXkDvTtDFdoRzILDD7ITP7lWiHEGnpA2+slndMTZJexEyDdKvgqjFw
f8CIJs62g2L77bR9SRlxzTLBmCcJv3XOBMEg145w31y77YZ629XjOOwo/3rKhZPd
qLBQdZkopCmpQNfD9bOsA9fHNuKIusxA0q3nnF/oVixld0TNyglnhlqzEIRw0IkP
TgCo/VFbNAXKJws2x7POGS2/yuXQ2fKKG2lpKrpglGs5wJDS6GT55TpI99yA1G3n
uXkXdW6P+Ts38DNewqpm8MrjSQvtpQFJn1JdN/Q+jk0e51OCtqJJUmDiKNYPwbV7
rcUDXIKTlZUCbsHji8tb9ZqZr4YtL3M6R26r1uaLgR6K3gm7oB4lcCx9YEPfcG0J
lYGDRspj4ZaLsYsAipaAFqGrU7TZfYCr7idzNJkjsVTbYkC0lOLt3VG0au+eXFCR
NQlcYire8ry2DGbROtNuZXvQAwY2GhVzja9hfEqFg4zKIJH7EDHxwjjw4qkVwQ+2
hdBe5hhtyx42w9zIzlL9y1bv3NrVgeinoiIwMPXlYPxg8wNwQL/61s4axdvmrObW
Dm1ZbhGeHD9AbzBHeOqQsm7VcSXps5NBMInsWlSkxTtAvaG+ic9DpW4orvI7x/a0
oAdIZ8ace1leugUMxJ9RyoHhZ2TIFPi0FaPJsdKHhSlhhfdsfJ53kRv7zY+QjVij
4q2HE2cCRvyTLJ6anpk/RFluI6O0Lypc4RyPmZmNla7wDfE7Z7Lin7dkwFXsoTEd
S8xhJNXAIJRahl7Z1IdQsg==
`protect END_PROTECTED
