`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fabQd83TkbfhzdaQKBAy68Usk0O9xhEkCgih/jia7Rp1EWSEw1KJp82VadFt0C+H
uyPxWbCR/rrfE5oxFu4GpdjffF7BZYHWAOij9JiCgUOydybVzGOMaiZK7duFpA+i
/QHjEWVQv6Vn7D6B7mX5+5dnd/wm++pJvOn93EP9G2LrDOjOZiVuMF/BOYYhYuXd
rXTDtjRI/D3XMOvII1/76EXiOXLqh23JsNUqMX05dsHb6p/fP6VLuipNEyJaKZbz
yyiUB7qeEqOoaZLXoD8i4soXX/Y7kWLgu5Hp++p5L/SE/QZ2YNwozur7ciajawMX
JRVF3ofeL0dtlbxoZvIuRsIw2BQdD6QoGkdcgLQsxW+SZ1v44CEKaWR5GfYLmUBT
79eRN+iW7fonBgENFopMwAjXsGI34Y1/n63Ldj7Mhjf/4/StMSG8u5MjtIiinCaY
u9ocST03jZIDb5P+kEEW85iYw7pxnaJIrTyoOpi7Y4VJZPtRNfHUi4yP5qH7/h4V
0nfPcOrlc1Us9cBqL7KZWeWpNuFv25Mtg0VU1k8vreGdL7HyLuoTiB5xJDq+huUs
uQ1W4Lr6qxS8PZlnbCjy4p3n79HrUFUBoAOfsXwUysBhdaWz6T7TYUSIA18P4qBj
OAtfHE4gt9sVx4sYOIBOUn4klAx1aDps6Vdo6u8wpFZBApz+asPTDx6ayXyNR8WS
kO9B+WzwiPcK10K/PB9dh8leg2q5YuauG7d1IpnXukGAkwNOJVYs771WqIrqEAzH
A6UcnMAve5To1VA5x7H43iPUDqYAq2HaANjtbmr+hGu+jv+B63c9YMnJ4FDDzSto
H8w1z41ATNZPnGXkiTADsbpIy3gPNjAMq+B2X1ZsOwZ1BZ7X47VXe/gOemFP491q
/csT3feAstjoDy13HFZHEChED++u/0X5X7CHx3GIAg2BgEmWNZlIpK34nI2tczLI
gpqS+QTxk9jtPVU176O3ZAs8nbpHXo0VMQ2AC6jcrG9RvkCWcNe7cqMZdwqjrF7D
50Km1DBzR0G0N59DMWmII7USU9b+tUUWDLeBKLtmJi5NmRSqpwEq0QxpGlNHwKjC
MF/rrWaBbbMd0s8p5QexCTGuzzlU76PCBgoLoUT11aac7aPHZSP3kt5a1Vo3ybnl
g8TaYKLpCWqDeCBsc2ktT7DFJ15s1/fLQAQCQ9mTKpnHVHiLdbPM8vcisJm6qimG
gGEphatl6SsZIBNl9qvsQKP2CzPitGdPhM9OYtVq0bi6PIE2Wpg7Y2sJRTRpBNxK
PCd/F2Xjn2pDrIwrWlIujGJnRyN/gb9Y3ryjkwMKeQWonVu9Nmhj8bLqPq/hWYMa
VTY122acJfPc8iNE3sFsM23hQWpzwlJrqJ3nynLKnOpX2JR+2AI4CsshhN3it0+t
y83QytT00NyGqCXiAtM861949PcXKnLcf2BgHcNaSoDlBKFyTzWWULqgOgqe+Q6j
R2AMJZB8EoEQuLjU/7tgvhKuN441sqDLhKDxvQxZdetUGsjmp87QLHWwwp60LXYG
iFIN8iCDKavrUL8AJKvLGQ0rnBKLCy2DSyMgbTz1KKPXD5DeGAL7n02+8ywQBAV5
ZnY4Bz0qk3gm2orGCSXIdFfdTwZY9qhJ07JBuCI8EpZgeTc8Rp9l+kOgpZsULpeT
oD5ALD1sbzv1cE61tGcSijdBMfFIsuD6lRAopWm1TyE7fn1BKKhs8DxUt08t4khs
RdlYJxvhQBC6d4/IkF12RwjKhpC5QZBxqYvSwrxLT6PDJAeyFMYW4JkAGk2mAEol
mJN52P8F2njb7SiUmIHzrTz5RLbA1s30ORNJFR9YmD/KTCCUQNDo0ruY0fze8ULu
Kbe1JPPezjqNkab0yErtRWcqIXZhkHWBrOWHl5c/yvXRXNMutIG3uG5oT5AIDrqO
pJhJCN5ZaPVJJIHAjFmbqCR/brZXbT0uamwljb2ToYTU8ETfMofKaonwY/yXRN6E
HPVIuWiRzcNpoVKNjM7tsbBK5jEgSjArL2m/FEuslCOVSr9D0XncAZH1dQyC94W4
DCBMV6pEb0HdCklFvWVbSCGzUn6uTjjC4yZreWHokl2YCWzA+Knxh3QKXTOSVfpI
JK4IpGRzDmW/+YmQAwN8BBsIJ+hz+HhkWYeneX/9fv842PCc4OuC/NcS/eGDmDzW
UMoqAglDUO3hNqz0wn/9H4HMnu0NrDGWM51LQkXL+IBQZlqhQqDVAdy94PywyAJo
YjWb7iGSUALXF/P8SJ14+y1Z9+PqxPg9f7XqvOUqfAFGYFwE9IUc0aDquammUSsr
oXC3JtEfOaNEa92vhwbNbp5Q8qtCJLDe2Bca2sFt4nMN1i0SWyYs1ofYR2nEgmch
1vM5ViYr6674ZdOL70nn3jA7a+pdiDB0/AqLrQycaGwvxC9ZzjP6kruRjAkaFWbZ
e6FBPRTKRbRrwAJ6Pa8nNp0q+vM5Nad2pufecYWR8ksrxlW3Sl/CuVidtMSZW4SZ
L6mOMFRtvoMrwxp8+mOsZ53S5AA6SAbQuVEYh9mAn8Kt9zXDpQeAymeTy0GTOJDB
0VzBXNaosIm/Igtk253t2+b/AOBnm5eiQo6QPixLGMZU20v/R2GSs/TcIZSCu7lK
JhC9tMzhEHczD74GWvWqmxwLR2o9iehCE0o5WxO/KRJ4AouexT+CftOHZmVRYBv3
VgbITY1w9JNq9Ee1v4U1mTja7aP4dLMy7guKjjzKbhbuLafHY0k9wywEgc1N6FVI
ciW/2iFseilj5KiazRd3MEtr1d9nIdrY6MKYZqCAEqWloSLCrVI10vXbQmaXxbMH
raa75jnWipcXkJnIbUhRt2PnGT4BXQGs+Sk0anODYCbH/fLD1WrFN/zXrUfC1eU8
fWJw9jWW8YyC6dnHM19gpH2HyPv1yyaHAGJTfwYlu0k07m+YWdaDaPBTJFMKNzMb
aIKBe3R+vNFWgnfnfOKeZ7brEFXYNWRYpcWElqNqLf8RnJkQsjat/n1OlODl1H0g
MfGq2BlClR0+bCvzSWjrxIG2Ugi+lY7VLhkZUs6/x+Y6/B85ZUTo+TE8y+sqp0Bx
OOWgwt/0F0/frfWsQ/Hsgzb8UUWnS7n56IGsyqCICEaq3PbEHPJYynDvip/vUZBA
XV/0bvsV3pCYAgEB25cC7m0Ux0at+XaamdbjfGn7jyKjqIcdMVv6whaYkl0FmRft
qJzA0s2SezCmM9DJmDvj+SNFo3AIej/IEUEPbie30QTPjm/GXJ5MsloCDmRzjLr6
F0ah/pq7AVzPwXPx1O3wp2quYlHK5YH9UABvpDbi8kpKaRkuppu3E0hNR/zR407Z
yY22q0/57OvQTNicnIDmaLu8X0LIwD/xP+WOPLl6MVT+Ml45nLYsY3Yiwv1yhHSd
itQ/tKRdsW/mifU4Metaj+H4ptkg2+sCOkL0zH4W1rySXlf+gvMA0xxTg1q2O9k2
YT2wVUaQTyKzpUZrglR7gYQrdlE7nNJM0w9CQSWgo0ELxeNuhymdfvPcKluXNZig
dODKcAEEP+keQbGYF+vI9i7fUmxvqn+/yxdgpH/Etxw9ieYfbLagxNIFieOnV2VU
HP1ioRU5n+tI+PkbKeI3iwHLm8i6eLJF7Vh0rHugQt3SOJomZ4arp4+ZyHZu9NoG
WLn7f8YiDMZQfpqvQsHz+vh2FjPYqoiVFZJiaP9d0Ba0Cl4o/jS1pJO3+5UO0U4N
86nSnzdwwbo6smauwbYahUQTGEQpHd9XT8THP7w4WUeAXmdzWJNiChuna+28j+xK
+jbETePNhmsEOARyvK+OVbl7kSuUgh4oUADE/U88XmgNa65pBqlzJyIRRwUBWZxI
+doJQRqqTn9agG2VysrLj0F2+v7irqfxXfD0B+zJxapc7nX7sE2Bgrh06k2QmbaN
YAA44DRVR4XFZJbhgB61h7ldzf38uZPyQ4qq7N1lWBpkZuoaJdvoPR59JY1VwCMy
HIcmxfhzEJbvA6V17qMWnvE60E/H/GZnHQkWDdCy1rLPEZ8lr/N0I5rp4x9WXwBq
rsmJ1xelCgpogtXbMsfbBMBQtRu/DLHefctGNFt3RZnbUE3tNam8xvf4Ok5r3iYN
KCBbYHKdlV+BwVeR7ckbSoZ980J4I0QPGMQlJgcKI6VKo0gipJU/WLLUlyRZCQxu
Axzyp7/kd+d0zZlPrwi/HZbFDZtavYA4TH3V1aLhNYTGZQTOk3j5AwU0Sx08OE1I
uyOdLGRKE/kMTgJlae+21XRKjnMhm84gRQxv04s4EZKE8btIcLMxfhtU/DBHL0sH
Isv/ZBFrqvQjm97BzmZTwRK9NYn10smijGZya4fptCRpovrW8dPAf9lcitoJy/SN
25NVzxhSddrC4ItuNxuWfaX7wx+KcpoyGHx6CwaYP1Ly+YTzhu6do3a5yxBLMsff
5ROLKX1A5375SurDYJ0+al98Ms4SDf7BM1ut9aDJJWMw1cyICZbMxXt9l1T93qGr
MkdU+/tyn2cKBUck5hW2swdfafcovq6+oa3T8+6GsHdV1rYiugqataz33RBVwFXk
C4KeWmRGEEul2ybTpmAOSyQttQIN2Lks7GsidYDhlSQZV1uF3zZcafq69SIsQFAo
ZKlTxVU7iKPNRzYT/xjPeqRKlDnuDYyE4Y/3fOIec1Y9c0HP8es6oArd/MtIRynk
WSh/ObH7grJA36q/Aw7kn960GSNpUjBNKIwFsXG7iY1uIBuO1AYMYr1gB4ybnsTz
fLZljyF9PTiVmxW+GxGUQ0s23+mrcGuRNZHPlk98RfHzEXg/Rkg9V+nI/A2SS6bt
Xf6wmc7qvibLPAzYO5rNGobTkRhmbmFItGtlJiFmgioNA++RMSCQ/lJE9EKcpILW
dXL1tqw1FFamanwpVzb1rn4RaizS2lrPYLG3z+6h2Uj5JisWBut2OsZww75VVZya
rGHNpWFSs7OMHPBMI+fyDYYxYpn+utIepk+oZYVddhexURKFgzvSLEwYKRlxl0Gr
qxrqnHP//kHiQsKm5DW5piolZR6NaUoevz3p3zFkf8POWWmb34Wq/3U8Crot1ZG6
yox8lNaVPvkRerGSjaqqZK/fi6a5WgfkAyneXWbMyQFLmV0UeEiPzbgejH4ZZhej
LZBKA596ZiZodEFDZK0xr3tTAKAkaE/mXgSP1g1VoMJgBVcY0jY1s8yDtzYhFSzs
VzrbsDujne0T8BxIMC/TBbBbcm75bA4mfS4c1LIwlOjoFTfJoxZYm4vhW2BIw0hr
A8stTLJFrzTxZR7oZlhkH+7DKHAMhdj5J7d2K2eN3oU7vAsJzjABvJNYA2F4ZLUG
XBWUY5Im2qozl4xUk9kptTh17x/ufkPxw3h9fiE8L3/olRU0mp5PNY0VZ+nT5YKy
vdYEm9/QFJUltebVH4fEAIHGIs8GFmi50a648RlOQaM5VZcuX4clQ7/sKtrMlARi
CEUJFEjr3zDd1XYS1UfiQNw2VKBTi/04pesW4VomQX1SaKocnDniYd3y19dgkp6R
O3GCp0j2k2qr5ASNjYNDk9OSICod1Rxq3xCZwNZYHuDIfxY2JEHv1My6Yx9ff2Ob
I/oQBkIi95JHPjtmTk9YuSFh0ro1qvBuzMce+/du6ededgvRFOKjWzbXhscVl0AK
xaGycjp0DH12r3UBlPD842NLU0iviPBehYp5L5o3jp/GYsX9jX7rfBwMKvMIQXfZ
nMcEya5EJydd/9wwvNe6Vrcc9QuXMFrzrgDhtxXyeR7fXsTh3Fr6jGsJseXojh1o
zuAvtQn+btnVBeXrkOsy72kM7fosfOlju4Wigc6NC4qCUjO25lcexRof6dPLOzWd
RsAKO/AyvW3BFrwdmJlyZdKEto8rlWQUlt70oRCihDNVVhHvlyHK0iVBYUeGrLsx
llihdFtKO7xOcXbW1VDuT0jOERS9QAvOX+PHDIU35DZFth8PxnsNBhhG4GsQuQtM
pw31wxyPToWIn6cXJ61G5CEhVl3BOwBS8OGadZqxFfDk1AxfBidKtJ1MPuB0ewki
olaEgG9oFvOlcbsvJlY8eVI58FjSm/2VPM9yoMZyHuE+aPw2ruEws4gMBLEto+/j
I9jPBLqWaCWJz5GV5b7/sfRMQ+9Bs60z8afsIhpy1PJwQ84vUncHrAXqqCEli5+M
apGIQS9NaFfUxYAifh0yz5vKgFTNFbeoyth0JuicKDh3HM/aQTA8JLWznlzsHIQb
sIXJrrGVAaSr3XVEJeAHo1kqgN140a/gvh8ql4cLISfky4B8usMY2HcTSELMWOo7
qS7XRmnY+tPCoz+qtmbkOou++P/aeMO8xDazs38zdddjyrgEhBA0AdlGuZFa0PJE
BtD8A5itcmyml/JWRxd53nVmuH2Jk2iK0lVlNvzaBa/d9BT7wzIV/YTJaJVCzwsW
JWh52yKhuaPXGTXhubTa4f1oVULS6ixZUPbpL+V+mjcpUxgdJMQcI7n3JN5ewTSs
a4EqVp0aMxmwOfZWyiMYn+/x+AIyckVMgC8fEJa5wgCXfnsfoVOzGJBHyOoHyuOh
kphUvKf41rbmaXFPRJpwo/yUNQ2xVxlMKCsTmtJI/gppy91sBAec1qHfwR5sPdvk
tX8tlHsjYguzsFYEA9poTyzUs22wfYO7DIxVF3xis6+Mfx0iorccDcbj+VnoY+E7
Pf7ON+dxQUzbcV6Jr6NN2pnkYKa15WrEKkYvOyDtkY7O9gxM406OC2CnLx2nn1ch
6TNL0swk/hKH6PnIJOHDEVdqT5tM7E6bXIvYC/tlq2fTysEZv0hIyfwTm6z76iV/
mpnSroRadFtSmjuHd4c01tADK35eG2WgCjHjIOI+OvzjcfERY/8P32DjN8o03Z3i
2bFFBSg33T7iddLpVB4WfImb3reMbNvkkDXXDE9Pqz5CJuxnx0k1xlKsB7K5d48V
W7sShPyYl56puST0Q54tENiSDC46EPweOvTnbn0yfkGv2GyMKgRHVe1KAnKTwjSs
l9J3z49NLJImM+1MYRxEf2LszrOBGzdd7wUZ+1nj4sMojnTAMFEII1HSoTCjlhJa
g7Hn1le4+/BnQnfTwhguAV+LqxS5ce/KbS/yfbffutqhhdAJ7qIoRrcK4tLVDGQ9
I1UWD43ZH7QXktFOnw8KYnlFuXshU3cnCcKNHZm5NiadRkPybe/ELseQggCCnwMR
mp8LIXZSSKOoK72S/pLTDsvw+M6/3sGVEoOH41eAdSIFuBqYNCGJC6hsf6qA7fgq
DPnAAAIwifYtmZxK1No/3hy9LGkBMafdyG/9WiXI1PY=
`protect END_PROTECTED
