`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X0JtRQ9TyIUJruqN1f/tkoaU2jnR93i55SjIm2UXIeSmTXMbJkxSrdcNkNUIJ6+L
Grw/tUmkV1iAoacKBTbVYCTaQAaDzgIHKJL+/dGWj5xQ+z8GihRHsDI+StNcvRQv
tMrT/UNExi4VUplIIEtKVQYQPHJB2kiw1fDl1WG6onCQ2V6WTs9DgyII6r4/MAbM
ymDSP1aXwNhAdVeglr787nQs/9YMhK4uNX2K0A8+1D9clEY6JuNVpgcwH3r+Ijz5
4cAi87fcdydqeNrTxYQW7FWm/NLSAtL+fljbHCSo0q4w/AkWkKIdZ81UGqKeUKFd
1S7NhEwheBOaVNh2YtugAMWdCM7zejejquta0Y6IWrHu4XdmQOwOx0TjWZOqgp0L
7MLZmMB+jE7817Vlq7QT6V7yU6kO1DcAzZ5Hcn0kLZgBJHa2PI0lJ+i2faoI2sIj
38n1lKol5jkZpWph66VLZgPFnB3YF02XN3FqiftlV1GG070viSLY2p9wavqlGWrN
PSWvXSE/0BAX9AJ6cXlrFuGd0D14B+9+E79PrGYKdgLV7nFs/+yj/1nuBrHMF3Iv
565BVsYLQ+RAA1TTct4fyBHRnwJLWz+YANtPF0T5joSuMF6A2uzU9Is7AlSFJ+9n
g+i3TfQt2L9WrOOnBrtiky7LDnfj5RKvUyKhwItdgaE=
`protect END_PROTECTED
