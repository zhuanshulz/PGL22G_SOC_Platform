`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6x7u/WwdHMiI/N/rpW1jbym3ump31Mrt9fBHff3AT+So1mqv6qrtogbLQ6A0Uydu
/vgYyyO8EqYVO+tFqOLo1zAX6rOHYEvfqDy28HJ/7kmIwMHNGQmzVM0bKfBKps7O
m14+80GecNncfvg8TYym2KvW93xD6PzL+FZaUybxlJrgfSucPFTVnmdFCLG+lqq+
ZN5vLFAmwKQwNNlZ4kNUH3NholzzpPOjbjSaiPDmWvtP2tYLJHenRaF1W6uWlYxP
ceRuVzXhOomUhR66h4vOXQ==
`protect END_PROTECTED
