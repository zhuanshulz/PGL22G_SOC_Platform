`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g4l8uo/tT8zronZaCRZ9EAAxkxEXxBnFZd16/++w11TEvfbIz++q+t1LonEXpEZ1
+KqaYUdRUsaWBSKVK6ybydseUNrPBm9QbcPqDvrF8hJYQ0PUtFceHQg3SSUe5UZQ
C0zc/qEa/dhBaQ5epPhtNkKXl4wRZ1qvMsiwFTxJaA6eZe1ldqNO0TF0idkZzk3g
1DsOLpso/3JYEhvVb/BZl9pLCWN7bTln0bUR4MgoV2GfIthCR/XiCSw0+Tdws4vj
J1P7NN+wy/ux7L33/bqrVXamcNQ3DhLmcZIlHdC/bc8TeiMWITaoDLTnItK79xe+
PVNl3PJ2b6FYjhXknmF9WvBc4CIoUhnWTW6adxTii/DvdtZIQDoxLNAE8q5b9Bwb
4j/FT0yP96k4OhKnKjDtHAaQyZYuXdpfivIXNJNCf3Ts3OK7Lk02wtL8v9a9tKaI
o8+sQEtfgW1xN5THIwcrmUQHr5V9q5Bfjv+fcQqFTEoR9hacyoT4/jFGJ3mDus8j
PvB7FSkMNrSqWeZ9Lw2S8laCkpKVje+USKjkiIqvx1wQr68x8fpt+aUx+HlnDhVm
SUevv62Xt/73D0NvxNfnTmBmqke/GBiYbqTkTpB7LzEbMMz2urjxpR0MgfX6QYew
MpVyd5MkJHnjBtH+WVzA+/GExOIsUcyTB5liDkCTj8DlUYlKmWukV+hYdwDusEJS
SzKpil8aBFrYDdGvPJhaxSUL7laYOytca0hgPD9lwWx6cjH98aNUZ5FmffIMPipK
CH7kv1YfELMkQ9fHE8E5THRH9kp51uY0vnEvNjt6v298yJhP88o9YulybzGvoQe1
`protect END_PROTECTED
