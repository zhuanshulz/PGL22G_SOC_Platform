`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w3+PlhACIAmFjTg+Mep3tY1SOXKuiAcODo9KTjkMxw4r3WnxKeT5PzRcWgz7dv+i
Zfmij85eXVMliTuPd+dotUsa7IHwm9TAME8PXfpXFvGowJHaCa5C6XawDV+Yey4K
czkhHLz+paeQGG07qvmSC5+vtHGGyXOQGQTUr83OhW7gjbwwOLRdk+ejXMvbS8o3
O3EczOzTFCQRsmbvundDdrKHGbacF/6RNq9bhi2XJJndw1ayaNH6F0yinxpELn+T
t8toKNW6lUaoukRzafGSqyJoaaDfAszi1/WrtxIvxvdGovAlkCa4WpXwgpOohBr9
05Qjy+snsiiix/rUdVl9f4sR3wblzGfqJKymxRYIag4cxkz9LG2ZeQTnnkQbrOOO
6/1dSoA96ntnGMCME8bwmNGJIJ19ZqZeN2hHaUo/Kuh5kIEwJeaM0+s/ZThitnU9
9JgMj+z1gZEKkTYg4UtpfTzVi45Pi2XZ0s3/IALMC0R6S82pi3NRZ3VqW5c/SlPc
oB7l11hOU2QM9f69CTC2QCTfhhWfF+eJpawC0ES+HS7CPExIsf2CVRfDxq/Q54eH
kAkgOG55HGWgpS2iMN8lnPp92UaPqcbA4A5UCyOg9xdZCMFkXA+fr9iBCldbf8M8
56PRkPoxxqeG86hPeOMwDDKnSTTH7P3QW+ZSdwY2zzXc4cp4bEBxh+Ie158/G0UD
wNgT3X3Cr1PQizjeOkSfHR+vDAJPeUDdyx19uvXarg3ZnoflSMFeRO926qI0IKiY
gmArqlTSy/7pQY8PFpbNbT+rQ6U0D6hbpWcxpZ2B+7NrhFrKcnMePHEJrm0d7TmR
Xdk7A7bDIMrYp+ay6jgMd+d161Op0QgWB5ITQbvB4JF8D/7pkmvPsf7z7lem3cAL
8Fj2JlcqWOxTE0uXmKZIipAQdxd/sNlFqGzvo64mB8tkTgkPQRHomWZ8fN66sEQr
URIoNiRL8SCUrzaI2gJ0M7qrsJ9rx18IAFYIcTfhZiloV3DYJntUCbMoNx7ry8pv
6gWLfnValZYF7rSgjLBxP15b3JYARWAjKi43ALqvNzpOjav3hEsz57WNJyJjcoUP
7Pp9rCClSckdWCL8MzZQQBKdUfvWTqCWdV4oyC7pKEKmw+CqClPX/z17ijyD+pWd
ieAGaV20TtVHY3JNH9VzTKXuoVlGFbqYBV6OsHBLgKAUId/Bm+9ksjhx5X598L0x
UjLL/64owXQ1f64roMHnuv1ou8Ut2buNn7Iqchx7md3ebQ9TxVUrgs9DWHSu+4Q9
CbEvGnm3zdUNRvKhgwwoxYQBIo5C5Aw6N0Cp5MyMXQbwJ32dg52ZlrW/hPpXDr0K
FVlvzBRDJ6gP+jYbO2QgWnKrmPE7UdIJdu9UTe4mpSuntknED33jThRBehJkVWWN
ayrncrenM/kpYJcYAKl7tfxmZhgq2tSYY/3bp9fyAyvETaobe25RGDrOIm4VXwGB
axClZuIrg+5QfcyPy17smJ/DOXm9oLSSK9Xhw47zfilKu2XreLbYCPjZye6O7Pfa
w1LDH9tJnOTzpdQWOT4OLuHgyZLdeBZqhQDdzqBp40UKXwhZ9Te8TemD3tAAboYM
2vYl9ZEFb+Mkq+RA/abz0WFLHYuk6qIqqUBU+aoK0Xk=
`protect END_PROTECTED
