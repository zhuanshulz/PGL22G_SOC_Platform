`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/zNSsNHNlmYRjfpidSEEpwgyvMm3WEneUvIBIEIuWA+4nofRy5Mlu2rRQhliOy1z
6OdUbid8PVHOh03IJ47k5N7rc0QzH3zw5anQ0OrefwnBGomTuHxNLDN4x5jbzRLn
PuVg0nQmtudy2h/X2u7Z9NyHr4MSLzLFcWcLiWtJxeVoro5HEwnpbuuOerBAYEAZ
OtoqCVG1XQhG80FcGXIBuKpWt5rpxpX9YML7pqL1qm4Xe0Q5RoocUQX0BjeHwCKd
icYQUvUuVkhZxTqsiX3jxqDsyZJirkokJystj5RhSqIQILhEzvMLX0zcQX04PhdN
pn8YCB3HCiMPXfY1TMIDrUwa9XTHcQuawf+aj8B5cc86sapCkbU3IEhUnQSFI2VO
9u0GBYwk5K8qSRhkhL5or6HStdOpVaJQNo3z57FB9wUuhhexgvP47Afik7MVhEQz
CuUpSCNBnYe9ZaPUtVX8T+uhPqm5v4sb+V3ROL80b1n2405xEPqeTfH/mMkYIjKa
Ih7uv7TLVsxEu+YG1BvEoXpfSuHxO9Bfkf4B8ltmoy+EgvgEKCvGNCvIfvPgMwh1
lc6cs8geDnIKCl/1TK1mIw==
`protect END_PROTECTED
