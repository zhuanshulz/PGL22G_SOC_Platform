`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/SkfD8RYXsvrwaJHYAKXJ3Zej/i/Rz8oXixnpqEeeGVnDw+zTCbriFbkIUQ+lg3Q
myn/Cwf1nN7dK5PcSoBLYNvxTnx8DVBDhQA3OEYPkj8lwS7U0dlRkFP+FWUyHs0c
wBSh2AyAej1HH0erxxfE+yHZ4JGNaQe4dycObzbY9xLTZRI0jImTa7aDOKaj538h
2cAnxDuQamg7fSldHNM6ams2RV6lzau2LOcDw5SfQdhYC3pscPImo0M55khEkFl5
VP0rwGhld7QTOnOsPXJ0uCs9+0MqPYGqnU7VyWkjnCsEGUKAedkyynn3YHeXIpf4
Wb7DZX4RidOpZT0HbgvEcpw2r491O9vOx3Oa4PbOroYmOHzXHqLOzJSPbpROsZdK
MVoNtA2lsOCAfS0OhBm83+dZU5rbRj4/o+VuTYtej0WKDv+lNYrm2nyoRbkTpFuS
1OU2xNJN97PxIirKfvVoX3Qe6F2g1iCXIGDYpHUNq9bHZs5Akbr+8OcB4opXmmTV
pUiCwRBloqXxxGrOnF02srZHPvLupjy45ePidUeIniP97LE2+stcyGsrcfdJYX/S
pe4l1i4pwN9pOFxgglNzoft+4n7r18mvPbueX5RS0THRK4rVgmRDa5xTmWX+zxrH
abskT9bb3tvZHzbFHhRUR9cww5M6Mo7KiMuTNhxmZPGC/t8lVp8vHukkDd3XEFs9
UCbG3R01vEp3xpUHKAiOSsjHttwLyo3DZnjOrSP4BAbfuR9KBf6Eb91duoTSRuGJ
HbvPCsgPPHUyOsIBJOqQul6PXdnQyOXb0Xwdel/6ewOVDMCUO5ffJu0yvCI5KnCS
uiXu1Fo9OqjFGDaNzLQ/sS6VyKCCiXqoFJ/4XpvL0oBN7MH555xmosevOqvyhCny
DLiSUENfObbuPk8AgiXVuvUAU1K5LmYbEVcsmyL9wdPBkmHVynkim07O2TLVlJsO
9ZvlJ/qk4/UUWuxbQB3YjVK+klDQBp3gEeImo7d2VxH8oJvUy8yb/FvJqnO8ECXc
cf2jhsjLIPo5bVyWRcxDdYyZA5ZhjqQA0WftZrAhyIx565Jk1Aw0qujxy+Fs7InB
GvgaA+sFV8Fa0fILuYq6pCdhC5o7Xu8gWsqulBkM39H9xkLrr5C3uomgu6FISVUX
4+NdU6OpFp68vbZXgWOj842h8leWnQomLME1H7hNK9Af7mQ517la3MXRq9BpC4pc
0ESQ0uDGjl8DYUnOYfaPe11KHd2eOvw+v0AlQIgAjJBO+efypd/6oot37xSwh8iR
DiazE4jib4HheHfXqY+XD5SmBtIwsQXxbee4RO1j3C+MeqdlfZm+UlvUE5Jh8UYE
vlWNGfRx6ncSkSqmVMWO0LNUNDehqq8ye7XN+uIe8vpwaXh9F8q/Nte7YqIPfyiH
8r/M1edUwFdREGWRtV/CNFchl60+bBLLx1X+TcR/BoHiVzUDgLW+s2Z3yZg1MVjk
7dN9yNQgv3DG+HjQBSAks+Ewr/d6FW17bHZO5MbsdrATMKCIz/+bcCNQFj/uQX98
LdokXX5Uidhvila/THczJo1LLOlQLqpU446k9MPK20ZFqb30KmX15YHj14CpfqZn
5cC2GJI8j8GIxalG0ugcoshD8t+TgTSkxJ16mkZhLXo8FT8xQS0V+3uHcn9iHI1m
Jab8N7H10AOfUzWEYxJN8QjUZnoRor5TJz2fzA15e/7tbW4OIyqzyEQks1n/bAlR
ebK5/WAFMWWGTD1rzhovlGSTfsK0WOZ+xYs4CHcaOOCSz4gj/ntdiIuvwi7WULG/
WG5tss+Q3PVZfkVpp2A3kk93uri6o7U+mwZ/QKz6lnwWaXXhh226MIBgoUMfGVwz
I2EAJxUwIovLeBKndM1oMevxq1PSfekAHhnrrbTpv22LL/duofParSgg99ggXXUP
F9VMo1ulwAJEDwHdDHc0hTxMqfAlXra+f/6tDjqtsEJBrR0mg0Gyg0W7vWPoyYHA
jkew1h2HrR8xN26A2QkFtbfFrn7Efps+eCvavG8bn5sAvEoZyN5++72DTj5TUNjP
AwFm/fVc71im+yg9QXOSpad7X6g20MDprEaFYZ7EQndZAas9PmXc0MqovWsY1Fe4
Z1et9//HHA+aCSnCivwbG/4pEUR0Vwij/Ml5WCU5aB3rqJRuMvUNx1Mh27xHScWk
bY0CL8zybk2SbFe/3X6jfnSQKdqCKY2daXl3eOeG+l5z3L2MSDvfC2YV2OuKh1BA
ClvH8Qjhb9rjX0xM6jX3K5VOnzzepQy0nHrHfxGtqL1ZKlnMF+g5ad4XU4ABwct3
UBKH1rVZeiS5JAA8IowoAuys5nhlzU2O2aI+sJExsmSMuZsBh4p1wI/wzFAeCv5B
vDfiCfxV1zy6h+o1XhUKHuFY+hnHyfFP//VM9ChXu5V9HHMHwDmHeEbl8IvF2tkK
vHFx9vtZ4VqOX3GcPODy95+HnkWP6xkpKQNvuguY5c0E1WVA/IgRwA4mratmE4Zi
2ychr8YHFJJTxKKt56dLqqwvL3StAwzseyjh/GZ3QfTzdlaTDjwjfGMLt3OHmq9x
FtKezHSxa6dyqxAMyUZjzYV871MbnBXodZQPmrQnauB8z/vEpSjIhHqS6sKvBKS7
D/zQMgRpcyn24OZ5jbQ9CYPgJKsjq90Xfxl1SkIP4YBBwx4CIdfWC0Sm2ixWpqeb
n/2j7zdVBjFKH7gpwpwmy0C6WRKBNJuQ2DMhh3lFSLUqezK0ym9LGEWYm3cN+Lei
Cch3o4DT2aVn8QUB1ZD/yshYnTI0g2GjAQHBQn+/sb6qzQVCpSMO88WDp2BBKSSQ
8Q5p0K0I5KHy+SgJSvjXC9UBcXB0NMH5zB8lpd/m64yaulwq4ti70uQSm5UJm8Ha
ExnqxlzRBK6Od9igUVvDnd17BK3Z9Q676dU2foz3lHzLmm+7Iq9uv+Ln1ys95Nxk
WAuTVX7eruuP6I5VSCZo1i722Hzfs0Rs9r1fgInTQ8AjXuZB/2pc7sZPZTYkdaAP
hk/Viny1yGjD7M2Q4ID1w4ZEC7wUnZhLWC+lg5GsugeFF17OZPH1NX0iKb5/UaM+
Ac7FH85NLwvnxX7B4QQH1upk7Qx73KHePJ5HHIsqtZRzgj1odtf9G7saTpL/f0C/
q/LjgOp766eLVJJtskZy9g8bxaE4oEiTozLZRdQWJ8cYYBgGx6HIMqvwML4/FIbi
if/8TNP+DI/ldQuXikIX//V86JpQt1LxOHUtRd6UHeWO/aLbgESDZzqsCROxLPE7
1U/YhfmoDymrNpxrKZozU1AxUv59FgrQD8FJBRwpDcPys+k8CXp0xqY4kUgOBQyZ
5BZLPygUEsHM39wWol/tqHLYIw/DQY8oSHsrAlsb+v0E3fKCg8rB+XClr2z7pgq3
2j7BgjLL6zzMFT2lGx7xlR+6tqRewjpyzODCbPTEa/QTZjHM/90nz9gMWnEe9kik
tOWHHnFMzAxPnuEVi8VFpHo6wES9C6Q+vs3WSiPhy6WC+cYNuV/N5w+L+sP5h1YC
Xtq24EWE2ed2lp2TmsMyXSQx/meAEJXvTr40et7abgc4yE4LBUqbPh8QOz8EV/K7
RMbW3OeNDFXB0VFpwkjQ1Y1NePzSKqdOgXGKxSo039o/cmLVt3Y06aT7lxZ9TeAc
Y0Co/tqqdp/Gyl0/WU/UFVJGY5p+6tgf+IQBHrMuqqjfhQGVgyEcEWSrI2IDca1V
+6YX2qmrSvHRRBkAXrXYbveBPlhaITGE5lPkv55PelP1VYuOQUAbznF6YtGW5m5W
dD6V26yUPg4eQiPeVvO40olioBPedjl6d25UoTXevP1fIsvosm+UuaVAkB6VZpY0
zVICI0DYQsLMNYxug9O3vr7zXWF9bfKgZYSq2hFOVuBrQ+teaYCg/r5sYDB/5Zs9
1WuyBARdgKacTcLzRMxoZviOwIbvRmkJpy0wtI8RkMTtKIY4QXbU6OuFbCxKnbto
foxa3iIBmUAguH55lYrjj67Axu3kjn7aI11lSlDam+Vt8aoBjF5YN3jb5f7zXvcU
tuvv21C4HcDcpwW6UrjsPoOO72fapwzBh4pCf3qaHORCTtLAGtDk4zBTB9pXeaKL
vbDYKBgtWYrOexqgGXErBlXdBE+rJPsyEyIMVJokqWQKRxXCbNAf0tu9LesBWn+9
7sE3+khVSkzCINfDrTfgVrwgQYBMOK8IVsPg/bn+03hFUH/l5TLP4AHPzGB1uMKB
FQpbLWb5tgBVXeKhN6KByiVtqOlyKN8L8DiI4ooAofe2uUdAjy68+qVHTfjYhQKx
86/YKVtz4VpxlW4rhIFbugJQnMNYTHqsLFTTcF53AbGHPDX25W/SzgylbYz4SCb+
LE5YV03M3j2lzP6Ckc0pBr2wGRmCD+fL8QcafPA7VLi4H0esKuU/EfqxwA7ZfeNd
srTLEajLsEMbpuyNoh1loITCHIJ9tvE1zktjTFH02XrkZsYB11izY/3t1eEePbGq
syeBkOJ/CRSAZbV3TY8rEG5bW0y7tOJnZqb+5TigYsBl0gFYaS3ZfCv5lFzHESGU
66YXW2e0Dmr14IYDq8FENMjQWL+9NOYRn8ddyp75EBwlLzEjgeIQIX/la9ViiRwf
6kKgvT0uXNMSg9rAjUvj4lY/NFrmjWliaE3KgyNOPoUKD481WUNLWNIk5/SmnmaE
sPg/V0INrAxUiWMxMMah7zvwzgYobVfoDFwHvGOXxqFAP0G0+jJ9mirSqOp7LGFE
vliFQsa//gsh47sycK4TJu8DrFDCMf091lrpHX2hmrCO4xTzqoglvUBTJ+OR2MA6
Mmw97bdv4I+aYQ4zZoMSuwCjF60i+rsRhtBz9XCzCaPnpTWSrXtMwucndyMTxxnu
z6unjiWAu3U+E78I9IOoFzuBsTYWlCRAVKPFvpvhrchUq3iUdhGJ+u2q97sGwZ34
LGhLajaoT/sY9Oes/KSu6wgvdUzU9rn/HTnO3hya2iKMR8w4TuzZOVFHOsPWM24r
eSW05k/NoxkiuHHG1r8z/P1i7pwcd3pcT9bwDO+QEFaQJZUR+k4WV7QMzX2EbaFR
KwB0oCZiBTHrDVOJ/uv4EdZcFamQiiU8W6KVjop6L2kgfTzsZJZQGeLkvdR20JCY
GIKt/gCrz5UKmJywVJc4uRWgogg8OkNwz736Mbd6I87jZie0AgTO00VZdVNIstE+
8m9oZccPUlAxw+qTi8Vw0Z7nqv6IDPtkGmHPHHa0YxjYB5+LS0DeEDyMpS9bbi3g
c61UbRyJ1KgdHiPFSQYqum8d1yVzqB2P3aH8/4nSHHbuQT737x4Vmv8RYRQVpyka
FsZQxwpiVgFSL5qc0OyH+/BzpBQFVfLS7w1VPddRH1WWcQHffV5HyUO7AGcxp7mC
Ty9i5HCWpMleUDkJ0SPfeE9zLCQ1+LaUbw9TIhb+DBZlJpLqTROou9uk2tOgvCr1
RjSnndJbhAMd4LvaZQRaiPKn6cpfuv8+tmF0eilKSiY3G/OdwJEeMckXgWTVTazP
IZ4AR6LJ3fhcTxbDA3oTA3TIQJo1d+vocf//Ju+yDI9LhhGAXrd1WWOzD4tiN2mw
M4OZqIo7AOpnL/TpAnuzvRSm20vNmfsN4K9QcF9v5biRzO4YTQiCR8ZO26qpaUoZ
pFna2zshy6G4aRRbcMkWjMhnelOVOMrTszX5CssR6chus5vD/k7Ou+H4l3JOFOW/
wSV/I82Nm19YHqpsmcQWsu5/Woucy0pEp+lSHnEeOwKL3vBOC+KaXBc9Oi/DdiJ4
wfTvbL2lczKPfOiVJSlKt7CU4kzTJjMetS8RB2UaMVfYdL/teoI0frR1po6/s1NM
7BpZWeOCMpBJgKWAm8hKIX3DvdOM+4Hbo8CHc11MBKYseFyM/vGTv/qQdrDefnQY
5nl826ArNKPAGLBTQo5GdiMYvc60iweUJp7qm1VIKR5cJY/L78+nF5Pljh5oPPZO
hHraqkUcd/ao/wIOvyUAHoeWZQTuD9fyUkClFZQ+hUaK62iWaLek9siSSDEsJdg1
ZZSJkLXomSx0YvMZTJ9y8iyr9/3mOAfu7wkceMFWl75v3zfNi60oiqSureJttXDq
Bd0Bin4ns5hgE0oXSO3ZLQ8zABD4+zslKZfb+hDvut6rl/gnQp5Cflvy7ObUoMJv
Lr1fGXV6C0BZlRWXWOK59mMNAPy51KHPf0E+cICW0wd60oukPUiMIGSopKVwAqcn
DHujpR+BcTVsf/oCKCaiIz743u2w9TJhYN6ISFL+Zct3nbg0Yh2X0MXPX7xWf6sw
EodumdULS+tKGHgon2jWiXslOzezSRMtdfibbZu/37cSI97j8x1d9wRpdm9FLBp+
tagIgbM+9zUHcxfFT8IqjciCJ4ULuR453Q7Cj9RY7gc8U6/qL9qvUMRHaFr/e3/L
6Wp3pL4JlQNm4eHGi4Klc0vSm4vZ5RSzoY9pqpRvZ0XalBUroRAco1VrIM7LhaTf
dy/D1D3Xq2mxq6wJiZ6w8rJnnyQOJpZBXNCFP3dhMy7FV1aZgAKSgbwxg0J06MW/
jbcRhZfoXuee/249gCHVocJI0An4xpEE+LQWCgUm7Z9Rrf1gbJSNSPx+3xREx8wk
rWZKY80IZgR5eGicVgTQPFiNrbaP3JzyKOFzyehx5c6YzOiQTANJBGEYmpoHEwdh
JHTGAqTewx6PP1tva1lS3Nx2JLxVlxfmMxtVsCcDyU8+ghAAePtiV+UlfYt6bKBV
5xo/QXEOox47qvNozdn0N6k7bAxXOJy2psAIAqFWdI9eYYqc9nYeIaBKEM0nAiV7
lv1QUsW+Npm9Hh27boQCJgJzkgXMwf6pmBrUtdRdDP8mi3JMFBjXIHcyQnIxGbZr
4DOqvT7O3z2AiH/f5QBLyrKN2IBnxEVDnxyKFemlHQ36KOaeZHlEwhmIS5ZONbnO
xjHUP2TF+e6YvZhrZDlNQdzw2mqoKkd3MURHo0nJ3SziUhviOXaxCFjomzsmcYnz
oeKUnzMcKk4H1N2Be899NiNWtdZeYPi+VKdqOE5eWcs2JvZ0DFy57u10TB8+ntCw
hgN5SnayB3YV7XQnMwqcv5pSQ9N46wclNGvUn6iDw+JOcN2Cmkq4dKjk7N1ZUmkf
52+1+GHgcoJ6sK2QiHxCGoJZ+6p8zcuQ6afuKzCy3u0zOep44kYm1iYKl/O2mCDa
Nj2xkbrdE0qpHtGkEZA0UZjVxXW+mb2Hd9vPm2dJDzSxgS697Jpg6egnBpCZ9awh
LKxp9tA1O5+NJ+JNyHjXsJjgsU0nD+/l+stcTzVcayaqpG9TNLPFjddrI0V7oNwi
JdFLrwD+KXJsUJy7Rdlxcbquh7NQlq/PpOqMizA5SUREQ89jBuxZkSmeUhSk7z9q
0kZKHFCj/xPt6QRE2kthZGbLMvbVQ4kwmh++3bh/DuO9Rmo+8E/qxOEqK7dsGxPF
We4GSIXqhtz2uPsP0WASu6wgtt1qZnt2sXWx4n6vAFstk8jXmR+yVrLfE278l7Ua
DVT4J3N+jpbPx60up01pn6/W8rRmeG48VbIJoRZR/zjaDDftqd896upP0wooDXCE
Vlto6U2KTJDGGhUwi5Yy5Jlx13SZd0V54IeACEmM7JNgWi1PwazReWQZaUvOrd2G
TkP+le99ufQJpphQgP71bvD/im0PeGd3aYPTAOPpDgl9Mf58v72sPKNhOqfkJKZr
4j2F9uhNarHZ+6h/R3FjdQJa17rDu30i82jU77jvAY+n/PHRCqXloAKZs/jfjW+K
mNR/QvyaP+0Rrnm2jZ1rVraYn7PClwG/xgWL5dZg6OfeLNFQIzNgSzqoQfTPRdHF
4w3ZpgSmRRZZimGuBwN+9mz/Mc0NSV+n7VDh1o5soDaJL08yvopcuBaN4L5m7EsX
vEoq+BGPO067HrP7fGGqdN1W7RfOJZYmRKaFdp0igzveQFPEU4WM1V4pPjlzyMTf
SuiGyzAt5zUKv93B5TuaZ8zt51G8qT61JZcaoRfVa6Pks19//AhDgwH8XQZFXIDS
d4SmEsyqekNbGmrKV6nq5COm7YfSpelL2saD9tn3q11LLwotCoilhM3+a4NohdoX
Fa7w1AcKJ8b5Mc5ikbK1pS++JzEtTKIz6/7JMb7DAXh+WmkGNQqhUhC0bGAmB/jM
RLVUidy5lpx8uCvMnM3fXYWXOyH/2JKplQ5e7YijYxjsPfOhzD8h9lki7rdpWqN9
zYGyEr0nS2lJgrpZJFFZ4/Soz3nQVbx0SITwG9k6kbZ8SnZ9ZAC0HgtCrmYYwi/d
V40PeJRaHXrmUEYfFL8DDT/7SpjpCNihuYzpSoY6+Qrg06uOluCOKc9aWeBIBW1y
kTiyQiF/1wRqqPptN6Z7LfqabfCYgNLPOQh4ygGivpdb4iDSEScvoaLcXywHwNMo
w//imw8QQe13nBQZupXG8diGVaYYx50SEcvnYZpdDWYg/BsQB+zhJF3WRb/UMGUu
LcX/VUJeTN0+08I49U2EKUDls6xHMo/vubalYzcPq1JeNRSMHEUR+g+hiJAuPXJO
oEFqvnP40lw575CgqrXRMyEuTP7tBMJE+MmR/Du50GYlxXt4qeVxqtJp7gPYbV8k
xeRKcB1Vk/J/JywvnWnLOqN0+bgkoqmFAvfaWSuCSG0mhDgevofQP2CjTr11VsbK
Pb4gRRGVa4CA8Qy62mEM6SlLqyzXkYvILEF1td6LfCJEmPBsZ2p9qyQNWRaO2koP
W3pgdhglMTFblH4QzQIDkrjZW8p1YSDqG25qCudmKk7Fm8R7WlO3Vt5UgaIWkmeb
vKR2qZDyxzxffIvcJ3zj+HJBkEEpvfhhE6UleGoGiDJMhmlY3GuyEyPG8Zv4x6fY
Ry9/UOqRLAT1HL5AJE0thkrHnL7LwClKl7euwh5qhj7WbXoFdt6tx6Lx40kUqeGv
kgogTGJE7dv2voH11Z50t4tSwGT6Mal7vX5f7pDbSg51KrfBhkupd/ZorKNwmr3Q
0gzNJPTHMYfwE7Ab9Ibru+LODSLeiHlCMKg77ZMqpXT0wK46YZUZu3j1TJGeshua
FxX5Ie0+TMahdS4+osw/9nOz/hrUr13PNmYDgiuexOayJGkRPC6g4nmQ3O5dUODk
AKDNM4oaiY9ePSvhdKha6j7d/CV7fYxAk0W67+yzvl0tmr/b+5923OovSGM2T2ss
f8ikTaf8MHKKKcrVQMDhkahN97lQqUO3VcJbt82AaLSMfW8WadDCzkQZ6E2NTzKz
FmV6adN8B0jMHPFRjKpppfZw/bvz4JoqYuQ0Tj8HsKBnnu67sahzvK7xOgzOerDP
XgtZvGp/5tfTtXRczfcCNNL4q1JfkyRlNxdY7LZPhlfIgENP1q3VQcnhYBf1wVKl
8HmVESZMRBTIkdoLGmdFCgpZBxkf1CcHwkOhOFAoJLhokAbodbrY/lMQp3jZVpbd
2zGL5z/yJiYK8lPZNkvNOpbNrgNRnHBFQdIGKQeOxR1n41uh9eH1f0rY0RCgOwbD
l8lC7PcTpWiVqDl4dwQD24FO58fim066wboA/lRFNgVPSYyNHXvH+HagZEoTQESB
my5ay7INQkEPfpdJnxy1h2ffu0TvvawfB2rc1xkNohcNs7mK5ma7CUm8fAb0JQbE
Yz1f7Qg22yUa45EMkhXg3URCZmTJAfvMZShEzXX+mdbmpVuy7AYgy8d8LpARzIh/
tMWUvEjaG7xL1z2CCwMrIrzAOxtjF/892pniz8pVlPhNJAnNBBSuWhXw0oUYnbSi
MkjLF3y382uT9BuIb8u/NfwxIa0emuCgeV7h/T3UmM6uIRH0YLO/Axm1L1NYEHSk
jR6pY0IfUZCiA8FJHRv3Xvs8sDZw41omkx15tW2PH+4P//TTbx5gRXgMoCMQTq3H
1bU+p8OdcakMhSDt8Wr3AQ74ec2Eyabz2+BGrcq5Ey3zW3ipUrKaJ4VtwXHg7Rw8
qySov+G4I6XXKJFEN3Dni3ZRwQri1dC8VainCpgOK6mhRVrEGhWUEdnQ60W+mFLO
lg9bl23qo8EKuNqQRwatjoXd7hTRCWa9ydmmD+QKNpRtpQibcA8bwgH1VIPGjvZ7
5KmwwypIULD6tCyCKZu0o9fUAvmbULuoPO5lcqQmSNk1n40WDZ4QayQOOJfSvPfc
cMJEFxoNR4vt8WVG3+o2PgCIhsU+hLEFA+z08Uomq8P7b6HSQmc9MDeTzG4i0u4Y
y+yQXJqx33pjwY6PsZaXQjMhiMt0TAgS2nKjpw8A9tCXaDil3duvI+gYt+wDLv4c
64xN6Gl3Y0BrcVBWNgoMyvlL6yoljtXfgyh3GbsIlz+b7mTRtbzcVc6JXfBuz/Ln
jUSenwaINaQd47nohFsl+ttiwA99DcogxgMSHwhIm5S4KnLreKJ5zOLsVXKDv+0c
Ggaaf7ghJ5K9LjO/IldFlYuprN+6rgbaYnZDVXLNRez4UNhPLXu9hT40a/2JDiV9
GvWNIrTC/yYsBsvHkknPk1jnlJriqKEV+Ndi46431aivRyWh8Z++hIOXBdD2K6uH
pWQt5q8SNQWiVymDqz19eEId24FoMCMtT60ZlUQcGiO6KJtp1LkxSogHyo1gW/9Z
`protect END_PROTECTED
