`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EH7/Bwoj2NrZLn+Kx/X0DZAoV/wkpRciCaqgs1f/0Yju6rfK9wXg+iMGWkQZo0tM
lc4kxZe81SDzxd1dBbFYWvvqetgx/IXqP2RxHaJ8kSVjmNZHG1SsdR2PsbmBOnq+
9HH7gAwePm4tful40gw3K1m5z2ZpBLmljqo5SAuO8oiY9IL04aRqtxAhqbUPXaJz
djf9XbtEDHiKVLwCO6s6XrpC3+C3nQG85Xo0dVSwOJKyNrp0jK8jX4ynSUqFYzEu
X6uh9xb/F/3/J46zlQjpyBCB/Bhi6tMRE1UlHfbz9BMw/J4Vzh1Euzy24UAx1Fkz
bcQuYmcjzgxTJolK+qvl8piEzGku3lQMwbp5M99ZDHehrfFbRx1uIz4WkdODz9uf
neLKr58H9FkA0+0jOcPZmsoxezeVYEP/IC61Uq8+loaWKIy1W5haoHyPjENJu4zl
`protect END_PROTECTED
