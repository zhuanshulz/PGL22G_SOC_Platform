`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o0SmNp1i/qRE8tJIVK9ojb4nsAcRjMP7Yehab4gkHbJ07FXjG+oq+sE9YxY1qi35
Y8J+pAN7tPyJLQAgLgOC2+aPeoRq6J+Z1N/Y/BgAzbzA13d5Gd8vTFDFnbUDJhRW
oiQzMMT+6n03VXV7u3ub/F7hinF2PiEEeTCUq/nPsgXPrl28WtFuoUUufpES/3lw
1I96hjKUrWJCNTxeZKtiBHMRslItmDRecUO8SYCwa9XU5Qz5vn2ykVhd+DmBPgwB
hhIuanD1FS7fyAVbvfdTMMFnNVSz8MfHMWOrB/SudbanPUBUHg7Pvj+p+dMTxtqJ
jDmW94EPnXysoTN533M9BWehlqS8C8IAZT5yP2HH8t2nlQSIQ7/w3oUkhXOWbqxz
KwgpWclPrO2rh6kiFoIlUcje5iszlWAs1k5pbgtva3ueoZyI/+cTj2kAGEI32k/g
SVt6DaTqr/NlrljMTbFY9/mUs5WvyoBdUbjGOQZPnXSqqgcTKNUQ+FDnIZHAHSzm
poFpZZyRnLc42IBXz8IkVtrmQMdw6a813bB6HKFcG3hyVybmqqfMYvqlh5jc9ha+
A2PEpFXYgz0NFB8hvdJqDLGTvEadbnJfqKcbNbZ9/BowjQx5ev+ZUE9nuxESthWi
/qV5/MGAWw4JdPFPrHddNZg2/C+MSI3ZPXsrIpbhih+N8Q7AgS6cYWa7JII+f1Sl
JTauxZOwBp7z3tOyvVglTXkvByAxFr21Y+LoYfeXubJYegoN6W5hX89LgXzgi/Bu
XEspheQs7UpJ2Neq+Jh3VO8QbChoWk14jWFCovkQf0E1l4wVrC9Q5Kd/lc96dFRq
lchdoG9Do9xZgloWxA8zz7ziXdyfyM63qW5R07Fh6yxg18ObHKocp5N2TFiNulcL
LG6EcvxgvV+6zgkPPoOMmGzzg7bMQir5GqVFSYBBtxM=
`protect END_PROTECTED
