`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qnVxTgQppBErLH36QvIdeDSplhjp1o90I8YlwRFW9076GMB0wc5663Rw3absjp0q
XvrfqCgfiekrHK6MiyVeZ8E13qIg1tXeIdluetqPgV/45o2f3p0fIScqtV0FWhrq
i9Od7z6Cea70bKQOEj5RhhcEQrZpRTn8Ys3W4DO2H8ACjn7bHH91agxR6IwMIhIa
4Vqdrlas+7R9RpRtyTXqL1Ecp2VRow3rw++EYFv2RkCfKybhiXs7bpS3oty9lWgI
`protect END_PROTECTED
