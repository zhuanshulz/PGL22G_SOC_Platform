`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zBjDjhoTFbPVpmVcmZxCiCHZfK+J3U1/vDOXu2QLDiDadPjpbiTIUPclzW8lqAGa
b2FaATQ6864Pst4rV1fU8WwyyWXoFu57y84pSkLMpnvynAfifT8lC7xLSGDR9hRJ
36NHuAUxqguFwajX7zGUd9eVJn83soXPUGjQOW5iXClvC53FcveebDe7nvn6vLi2
0r6fJrGKTxueB3zEaMNcJ6vzyBGVFQXdLYng+yGhJs+lsL3x7TaQw90NEYOybMyP
IAZMGAJi0gTY++Poawd1Mu6hj+DtLrizFGNbCgn2xTFALIUlOioUD0vxbtoQAXvF
+NkznXILZw8XTxmM3Tky5/j2RbMdekuYKcXEdgxT21IZC8TdMvfF32MV1bVzfd1u
5RtbOvqbthltqf2qEqr/VwZy/Y3+Q8YB7LpPSYobZmvAPt1M4zUuQ5ATZLEKicgi
AE9L5L/YExX8BtyHAVSizECEzcMmlBqY4f3ncHDgYf5Ek5x/Bs+iK7ZfqrLKDwyt
JdxRijfX3PN+Lbuq+vBIJdlkIdLG4Qy0d3vA1SVUtMbz/X0qE1+/SjxycJ+fbF5L
bwGlVG963K0ZHKfJ+qQMptmZwe+KfO2szFgXTSBD4zB9DPzP4dKOShkSLIuKzdtJ
zaMr/hve9O8ml8wXpPewkbwS+PAdghGgL6Mjjbpb68z1NTE3hEctB6lRRau21e5H
CbdK2PVyHhZdHDXpBUxXSUJLUSy+gAvMTaXFmlArAVToOMR1ugdShJ+a6QikG5QF
+r+CnQN7dZbnD+piUFULrVjUYXPNmDzWYWVMef47VsOLWRG88ZNey52zsgQqdYIa
LDC2/t5PFlm9R/uKCQejWF+9W42OdRzrbwoqcRJjSBxGHJHv08PRQYNC0NPQOJRZ
90uA9kYXPcEa74MNRaRd6RM2CAIGM/LtFTedG06vFlhOc0O+F554oP2IaJCN94Ri
lNGXFfmL5dBcbB4a8HV64jxPy5u9/fHtJIOfikpp9npsYCophk0Vb3KmO3MoONNX
Mgmfh/GuyMFcl+jLgYXENvTlgbF9fNxzMx8G6cpn1TrCXW6322BMOd8zW6y2fSbq
Dj8zc2McySa+u0ITmLHGugp3L0sP59p+TCextwuEWoXO0q+t6ECgUr/Ppa2W1rbU
qfxvbvekhalL+Esb4G6HZwhBZcMW7YaK/W5WUG0R21yxmVX4SmT58arvYemMUOTf
XTL3eFG2Udcfn2Y7FCNuhoHinoFSgK+rNJdnj7a8nbCIvkqX1ngO33LxXISrNKvN
h5IthkiPNpM6bSk3dAscK1D8mG+/9DXm8HzcM/K81wnU3Zb36NhF21Zd114dQ8Of
259jtEplMhlKju7mJvA7/keVNE9vpN93M12uxGAU0WB8CLfvW25t33rFqC2XkJ6k
vKdgOqrqIwBeRoeejpb9U9rxaeZNGxhHJUKMuOM6b1t84fgu0CUem78UdqiRLI0r
ii72Zra/XxbfZeFuKUBtvOq1Uxv7X4AFPAqg88sDM25hcwLDfp5b1M5wRLqYxGz7
bOoIZw/i6Rmk58zCDExSLLwCWO1MOiZ36NaZPdrWcIzvMIh0EMO0fUOmD+HjpOdS
7rTD5w9Tw2TjotA8cRoBtSQeuQHSRCKiiBXZxzavq+kDQVeR4dxhjvaCLLHg39xs
yBzT9naeTBl6LcovDdStByVEZQL8kE/iIgftQXicfeP6qa/bUva2+OaxHtFOK9o9
xTrMTpVj2D0xnORT48j2jz51JRXHK8RUzoA1wkI1dzzE6SnL1kpTQBWJdjua9gMR
UAYXBiyCwPVB54/4rw1wvwDU8HgsAoJAKMoNMrX1Fehsj62kKxtdZmDuWoehc7Jd
/EhrBQVnkyoX+YDxLvjBPf2JFD/4V+IaH+csD5m805zaXYkihdcL54DveFxFpo9j
lmAWvkJ+D2e178bg/pIAA/R/nPxAtqQ17xW6jsiv4iYp5hbun/YCZSNBXZHmfTfK
nBNdAWxpSawk86ysRr4JHs/jTYK2xtmQRgL7P+h9mJ17zuh6sxx1UlXJbbbnNYS3
5bzM2rzKc9KbI2CbJQjSFm/klwXEe5xREc6l8S7ZaENj3nVA1M6a4QPKaPxPeGAC
LM6RlXuBJmVL90ldCPmLboc3JXi9U51Hn+hfA2D4iveWOaboeixEbQEXsgfkIj+A
zBHzMUyJJ8rwALujk8x6qpkhyA/2wvDBPlNqI1sBNOmU5T62jurY9Q9wGcJQT9hj
dn4uoeh7FlcvdGINXqlp822m3/de9MtWf2XzrYuwhz1o4Eg/TSP5z49BiMT2Y2o/
ACUyI7V9JABZqwKjECyIslYMg+91RRiUFfB4TSd/tW0gjEmoDyegN96gl1yUnf4s
HgYIr6nJPyp5/axKKwTzxNUSJRCSH6yHDwinjIORsKC6h3O5cvCxaAixt5NSIvQ2
2LXRYSaXIVZAeaTmh3/NxB4MW/GRbinAYUo6SKpTfzG9R8F0Id0t0szp0Z1r7BDV
FluhKEQab1JEPg/NkcvoFuZDXYRs1lSu2m1iZ3W2RpZCmzBese+WBcS5hv/dJzw8
WDygSUQJFAVHwDF2C4UmUA==
`protect END_PROTECTED
