`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UDiglfguS79+SzdiL9WMEcaPtq+5ZhYEkBROtvH6K+pVibtTqGAyQ7ZjmiuUpj0k
+SlrxdAKjoFMAGU1HJSg2+kguhRmOKdWrpQac/ZdiZoPeoHi2sBSc++2E3Bs4VhV
sbe/p5P7UsbfUxi8BaQRhbVux7h4toBQ00cJfgDfLfm1l+Gb3pkkA+kbBUIPUG4l
wRIcqmf0EnL3srteAddx30JKWc2uLtfOuk16se35L9UBTR7aFbbjAQI4GutrqAFq
xVH+T8Eqkv8jzM5N4jCWZbmZmVqzO+pmOlRTtV0KzQm6YOkg+5XYObCMNfLJ6naZ
OsrPm+wd114b+Dvh9f48WEWwyWwi4mDU2kT1D4I/15qw1HMwJx3WGHZUTl7CfN5/
n+u1ntyKCZNFFiZ7W4RuOsNp2Gf5fisDi6KzLbqPuZFnHl7hMXJJsByd7E7EKtrZ
19dQC8RZiZ3t22womoqw1/aXkcoYem8ByUS7V4YjdB4WyPPeIyOJvQqrBxzvKDGe
XcbGcX/hQWJ0UcLZf8xs0A==
`protect END_PROTECTED
