`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M6djipVAywtr4fmNkyc69Rou4nMXtJH/e6f8kLwDu6Fi2tJ8RWJYEC5mOqN3eXDG
NDxHyWi9p/UW342RZ6CEtl7pb2tLKUkpmCGGiJM7e6Ea72e1uwTUCK3ZNuZzjlkC
uldyP+bXmxk4YObtwxiaPQHhaiQ3PC9pSq3LnpdoV657EqUdySMTHG5855dR1opu
xU9obZfVvYwNvud3IIu74P++Nwe9qOnxKgR/XBOBzB8BK0180oNCDETyWBdoV9AG
lxfmDzDnQxStmGhsGtswXLdakqcFRR+XblNiRSeW3vMG+j6Mr+JIEPg7xeAF9t2i
DXJ6Q6MW6gjkORiq5IfBMeCWN0+FO4zaGZgniQSGSF4hT39/HYihR0WVbq0SEKmN
LV0zE9+Lj3m8bOFLrwCXrg42Fyglh4HUEc/dcYF1r8CqdsaTX00iTL27Q6w6+pB5
AFHPUIIyUCgX/Sk/zKcUwizhZPVqwwI5Rzf2FYVtPPcmA9vN25OnvmKkBdQLCIg2
dX1m010JtO/8dHBk7vRyq40lJ2NSyaCX7g8C190dpl/V2oIkWv44IauRCyqHEoax
1eobtqQNnWLoPZNWIEMpzH1e/kHo2TIKRobjtlFerwGUUKr9TP8DEhLbjUEzqPzk
hRsTKnJ3z+KpudGjEcDWCp5/yGa4gUi/xkezVI0LPOqZJHoZ5r+TqJGOeZERqeFQ
JW3gsuW1nIorc8tik3yvY598Zcqdr6PBHYp1lXbiYEJSck/K2RF2jKUWyOcqv9On
Pn9ll2w6lduyRAiRr0LcFJjgDpwqU/M1m/9Nvb3EIx/LlU2/azIxGFVJLBVyFt0U
yrToaSQ7nWfZJESbUxqNjjvcscdyGxmnFWgqzR2jNDf+vsgKCIPo9ZDFlMQN8YMJ
JvKG1Nc1zD+mNfaxE82ZjXyFN1cyHiL1bglteCK9hEojq4vI7prEx4XIFGDp8VFa
StglzOCKrRvk7PfqhuzYRxsBXu0V95kO6d6s+rnpCmFYYwo+Pz9XeLHr5uhsBb8s
nZe4B0BhngbnW+uAuTY5k0cuJf1kAy3cUTDUCRf39RZhnDkOigy+wTiaQZAdrqfi
HeamEI5ymf+eHIr4p56P631Pd+5ZCC1D3pO6bebs//ruexg4dDld9esZUqI4nY4j
qcq44L8/I/wDKukr0ak2De6spjfSGCp2IhAue79OiRTMNzSBFLQ38cUwHZKveL0w
z+GCJMQ7opII80n1/jbWcxgcSORCFMWrlVL5HoxDabYT5B6MN6UXQ9fSxw/O68na
OfJ5S30ncwt6ivBuDJ1ChXh8o/olAePfrLD/5MsXJ/m9Lm9dQWjylWY2cc83B/Ej
waeHeW+5IXTx95TMt7Fw0tfJO3XDJyDht8+zNmWZpJQ6FJLD9vtdElgptMfM80T5
yj1i88K2/9oBs7fpIFHcX/n+LJnvkcnhcI2UapnoKER+V5B0q4hk6dkJ1YlhQ0D0
B4S/3hg4zrQoctNE+5LkbhxQrplJJsH9gqroCxVmNzF6oDdmJlbmR/KB9LN96dAV
uoxLC9ZHh+hJqvRxDgsBeeqaqDS8ZplK7fGTuaMryN9Bo405rTlzNMkLYGJarEih
oBQLy2UtQFNEKR0C9MyxaI467GT2xjDO4a8lE36bymHdZQyjKEbEvlupO8Kbl3xc
as6Daw5d27A0ozBpLJTA1t+Rz1omfh884C1qM0hd9OG+rn7Ka8oBPRLZ6p4AGG8E
Jrj76v+RaE/Ty+PIQPn+vPdBs2JXw5kCIfim7xcTBnx4yy6z9fILqTj1IJcSSF4Y
w0oEKND8rcwP5/lg6fbXVm208SqZSr3TOs6JFpCkxOtTBrh/LBBsaUaW41kGVfGf
zbRKOTAK3z2krrdt8TrJM7EQ14eldJ0OIhZkbeIXr2lKk9AwCpdcyl7h9nKJ2BDI
5dWb8vC0PCSq+9rYeEmm6gJgmM63XMozx1GB/frkdednbldc3q+u7Ye3VLFyd8fr
t5EoCTFWRNkdkRZd6NaDwRSDGiOrrq/KmUi9ZHjN36J15/a7lYMkZ6C0oQlf7wFn
hS26p6wDNDZGPvykbYZOB+4dsJCPOzm2SHgcGOZUeeXon4jGbkqthxDdrm6X+47e
/JUkryt79W8BYA1xK1BVZmlfHWRDvUprqSGGw6Wi1V9qOZchS8NR6qXTChF0vWa4
Eg0ipHu/Rah8tLG+M6LbcxkrLuR/f06MGbuYQYPb+vwzZFNbupRYud73ZiKbiR8A
66omHhXs2vz/Jrt6rMkC7ZjAUY5nDpBMaK59Hq0ugHVEd32omPO40p8ZP5L7hdIQ
WWrdbrfZKHuZ2Rc3jFSN51PpbVY0Lz0FN40Pm8J6caDhF7KyBhl+N0sdl7GNX745
gqg+laTUYWans6mwD5tk6L1jT3IwVF1zeP+6tJD1oJkT0gXO9pGmtfp6V4POU7/y
qBa8UEAaM5cX1H0jz5fTLj0I6FoUCq+FCv4FthYXvhvJXfIh9hgjYzPOh8jL1WQe
KD1bW3sZK8MzTYfsekTQdQ6luKVwkY3c+mwBDIliCND/o4TZFRE6xx1v99bBsQgA
sk9h2z86iZeyEW9QoVowf0sMVobf7R4FL73v5Qjrz3l1UawDCPYdYM47c/V/Lfrh
DIg29k6XE5BQtaCyKDf8vubHdzLJiN2k88JZf3pSPPvHvyinjQAMkuEmGYUi8vIu
eOGtgN7TH6zQ/EAW2R43qDHLpAk+D/YqXEGtMaaZpmLrqAXHMSu2ZlABg/Ikkug9
dDwC5yPE/igJ62MI9cqy8nZSJs4w/adnR/LPqeSKc8p2bsfGKZs5hy7a7skGD1yr
`protect END_PROTECTED
