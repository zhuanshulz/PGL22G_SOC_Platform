`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uSrgiyGWr7txcMvcymvLIYn+2gjMInUjch8cbTC1qoq7mVEpM3I2oto3vtwujb/D
n9oPvuIyacJ8y+OpgToZV1xngyMPzynel93bkyatny6YaRxW87hBw1F36jVtygT8
UvHu5RQMIvPeWxOb3NjbRz4df5n4Q8Pcj6mkTX79lG5IiK9aqzUJFjLB+BjSNVui
9sJG1jnJLr2OnICII/IMT43z4X1FUKV8UOM6SBW9P9ykwMxWARNlm3tGw3AjwOOy
eeR3FjFBtr7hxXiWubAM8h6dpdhC+q03Hp5Mwbd3vzbFdsyvh5Bztnm8CY6L8Sr2
3F1rqhTCwkmLejscuO7ZBrG5nyWOs891KmmY9aN58wvwXZRh2kFjVZ/244aS0Cxy
RzuW7ucAvm//0TGLP56M4bjpP/ww4GUdy4PkZJGo0e0=
`protect END_PROTECTED
