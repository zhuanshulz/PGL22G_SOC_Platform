`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hTT0ouLGCsgKFP3SC8U0PZzqxJJ0Hfh8+k2/+Rro58F+pbF3oDykw42llfEypu4g
UGIwzKtUhERDYg6YJbIWFCHib8zGt0Q5ZkT6AQywFupXP37waa/pvqemgBEztWXf
R9m8TRKYhV0Vbks4egduk6jh0VS4G7bYs3oyRg3Qh+HBel+ZVA3TNxGjt0Tpx2hB
vmjQCCEZve+3bR+2ToAweQuwJuiPOtvZ71kSDPfi5ldXKBjiPXmpI8Oz3vMYfx4y
Id1a0HXygVhsS5w6kS3l4tWjQ+DbGzhFkk8eYMzJTNOSLxk4WYZp5gy0u+I1stO9
g7P5AwLyBqpFM5UEY93nXZHAwV/ZFSOmQj4mLBQAtRk=
`protect END_PROTECTED
