`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wgsmddW76xm1O9KHIyE0xp0uIBjIhJHJojjWhv2HWcNEMoFFDK+DflpPn/WVmUxn
+oT2gGJM2tBz/aVwTbDWn9Y8dgmRjkXFvft3SjirYYMJXYxST30wx1Sd2Lcr9n1I
sT3cam1Gqlq8arYHK6cjMqvc77LjfksySgHWf68DCBK8tw0bgz8PxGOIg0LnSsod
udEiGJOfUPMQB/cncWZ43Ys0zLtMXOi2KkUa7yv3edz3wzkWZKoVr4mmIxsg6mJk
GLScKXbCpmvib6RHW6bzf74GnvsrjXAjUbr5+afb3dHxuB67ySp5QrKReBYnfy/X
vK1p7aPH9I8riK94I6urc7/bk5uNWZpSJlO2OhBthHFqDyNLZzO73kHbMw6HenZt
fZUojSZp/JoyJXZv//BJK2EI9IgJDaCkZeEyIKfi/me/Y0LiGwqqiI3EmpF2Gi35
NORo+xhTWzeTkjEiVzLEMg==
`protect END_PROTECTED
