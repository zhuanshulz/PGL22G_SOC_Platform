`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zwQ68ncqPrJ7EGHO/dD8tmKY2UhAbm4INAgXehnP56LfdxcDIPGD3pu2hiDXnk/+
neDO2S+cR+4eSwUfYHzrO0EHH1cKzh3F7h2j1Tt1fxRUU4vVlUE4GdxWokQKzmvk
AKXYuSLQ4VmXEzS5DlTWu8RCdsZgUxF5NwdX3SpbmmJbbsRbbJmQWOCyIyKRLL9P
jjwei1HYcuJPxxnuUZBPcxYjmu9dgzqPalimzeQtYwvumjAN7d2SfDmzYxcF3VnC
asVxlddVcpkwTy5qCjJzvAoajO1cAHsA7WBZgK5U1ixylyPM9wqP98Epe6/6GJcT
pmSDpmwSwW/kDfgUrbiPm8bE+WtKFGlcOzNHexrPn+RRBB/HIWuNwmxWLNBurVQo
BEVrMENXLcKHU7fzHnw+O19CGvW6jzuL1SiDKHYzo1UNcHqPHXex2MXPhSQXcXNP
+cyGErKtYnVoqghKvAR2ObV6NpHkZeJe5kyYM4eEhLytjSTT0Dx1Llc7jP/GH6/O
aqlNG3meGo83qQM/0WZyD1CbjZkEh29s2a9eq0HMm1njIA6JvNJB4R3zWx8EyWoO
`protect END_PROTECTED
