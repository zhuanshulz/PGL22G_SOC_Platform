`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4aBia/srGMbBb4IrQVwLZ1XtjXQCgK4/jLO3xUZ3NFEz8NbmhenXlc6rlbETXljm
ZIcy1Xc6CekoUUT6+xV58bpMUXZx+womrptzVBSZt/3X5pA97CFeno1K6j6URDlT
oFQW1fxeBrBd4ysoAiaZmZ8nXvVuKJI6KoX60Iau5f6OiTTSk7JPKPFnxSt3Itbl
dIov7fH186Tc9ielVKhzZzWPDaE+XIBBWDQl/wB2a++H9nINpQ/YSCTR2+bcf49D
psJyfaZgM2B19EwCFZn6CPhBAxnmaU2YezxvjKC5T5Pp73jggJWz3nJYU2GNoxfK
bGGCxqFPFg3lkJQabXkNNyQiO40Io6iU7nuW4817BzY19crMFG9Lju2qUmn7+XAC
DGkVr5RpIoK8oyLq7i56mZ4hJ3kOEz/M8ADSWNMvDs9N7jmvLlT8AMJPzSwhyVMa
jkWM5VMuOo09sYB8ft0MV/QAtzuwIxkBZxj/Mhy8RAA+N/Ec/+Sflm1IFUu4fqIX
8cnkVJfhl1hgDwp5lw+Ribcgl2OLCcST6+FQKq8Zq7Ih8uHwPYf5/o31ooMdBTkY
Y82B9UQVMAcH9u/bhq+aNThugN18KQcjeymFBiiIKudCurhMdzDpSsjd1KxzY2wW
1m8Gs9u9kgHtDJEvzJsVXQglvSdbxj5qtFYBd2v+dlYNnemGEazbSNIa7jfQe+ci
ocwXL9sLs0smyrQWh8PE9H1YJ01N/zSV514GKTii0r/6TdwSop25rIxHVnlcB/s5
uoa0AFov1T7bKphe615t6t3xS9b+mABS+Gis/s4KvPbcI/8O5J42IuZ6dTVQoPWz
1Hg6qCS2CIauGtHvUKtnmJ2lZYHmo4SH7yYQp3RKMxsZIhZ3zGQsn6qTgXjXpVeA
KrP2u9KnyleGrh6onMQu4rI8S6ehdqWOA1g6MDixdwqr3PvMeNk9X6txbXS/b/TM
NKaxbOUiw9BCp6fptmmRIf98BxMcmB+a6GdAqPJZmTR7CUcqTYoHpCWpTWpsR8Bb
x71EJ8sYvVF31x8l++mJigJmU1IJKTkaTlwDGC4vdjNUVVkAK2sx7gbfF5nEbwRp
hsNDHp53kGfYUKypsWzUJoKCkcb9THUiSFfQK77IRHap0gUTgL7hqYrxHsN5iiHJ
`protect END_PROTECTED
