`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QFMTnHsEBe6fEnT/e5BcDORmjRQQkyVSgw7cxJ4Fx6nN/Z0/BmMq4+uDsT7COQA4
RYMKYEHgQCmlbNGWBv2qSk1UcPB1LZLNvwJae2zQCJWjogk+H9QprEgAMY0fBJj+
PNLNcYWLJBVJA8rHkrDv9TikDTDBB/r2y8a1QywiQIhTb5sPJLvWDzuJ/YcLL+rR
4NSP//21jdaB77vD/FTu9xqsjii5inngcVLI5EK3ajDOQQPdRZFwL+XMRb4dPK3Z
YurF8dTgXjPOEV7hBAby9Gx04sJ95EmwM/hlda2ocl2QepQI9Hpi3ZzkjuLMbni3
ItcWRdFLmLt3QmGBCd+TNJLJouRtXGXIt4hIFxSpm7vQ/foP//k7RWocfn4orUwl
oUo+d1qumUj4sGoEdeKOCN2OMELEQvUgovnd0t434eAAG5Bv3ttCavvO1Z19xoV/
NVZaoLot0mDw6oEQkX2ybmFi4AVtE/uWNWdF0yx71ioXkDYumqjshGlnl1xIhu63
hN8vuctDK3XKnMLT4BTXwT7HDSQ2H0ibRRf7gmwr9tIAEaeZUiQoHqT1G9bKMPdV
R945XVEFCsy9ed5IiNNRzsCZJLp4ugrUEj34DDF9OrCsWOqWMdhBxxxXWVwNb4Cy
UN1yk7LColZGa1GUUgU9sYX+cEDhtM4/VrHvS45zzB+n7TtObiSjrQG5IoxISuZE
L72kcKdEFjp4J/jxh+KkbmnbQFwz7LmkJE71W3aBKRR7cVHNbKbLTTvrpcQLKnJJ
3RRq45A7LoDp7s95bKUmCLO4Z0J2GoPlYCJ6AEb9CqXm3FnnSWSfi7wrcKZVzkJ8
KC6fEZjrkKf0SjYg9d86OcS8NHl74nqSZ8QVtl5YYdpjJU4kyCVqq6Sc+Pq5laqS
bCJ4Mlr/z07L/Vsw2RFCf1gxIx8aL4OW7SAyG0Ef6IhNroEEiR57j3rCoq9vUDbh
rxcV+HMXsrWHQSN+WzhZ6LcV5qv8nLeuQKRmcO5kJCnmpeGvrW7Uebu1iInYC1fJ
60nYd8PxGNsxrp6z4Sc3aAf4+dL0kW8MnY14HlZ65JA/4svke2l2u0HpyACC7/uM
FBbfqrMA0mfUhcRHKdx5gukmgiSbr3W2JDUJbXH2GCbzzMJjp7OZu/yP+FdPIbJx
RUgOfGrR4Y2vI9XM60ArVcvZJLJ3M8ZYESrzbnV88LLfgtewTyaohGlFCqbw0oUJ
POMSdrMVRBE7TdmyznGyElEFRRJEQQVxx+KrTTOBkE1jLsjMj6Awm63CPdDByH2d
BB0IhKToBopR0lmq19S6zV5cjR9FOwEcElzrqwWPagib7ICmsz+VK5LOk4/Aj/Wd
z9HQ0/ev4i8xAn9syg+NTOKvAxmsq0rsOrzcvDK4RPnUPQxUzEARIhS16QDyzwNR
ijvRtYhF98k5DqIC8dwvMiLIUzxs7w6uSdqaBRZwRrzJeNxER8kec0kUWStinR4V
pzQ3YFjD0AIWazhAYeZiWye8behurDzrvWa6mUGacwl7XvQwypLYCejMdpEmV7c0
8rOeaEyVp4HhuAv8Sl3VsM1r7eaM+sKYpnCA/a/fMXiUp9tkqXJSjqSJYVtuC0mT
1I8IaOq+vrc+eH/Np07Ho3bdy8Boy8qpz/KnH8jFDz3ST1tDMgWitf7yjUrhk5uf
6D0waMuUyCGPHEu3lNCqo3POQdWNJUqC930/S5k58WzGibxE1T1583QQ7D2UPRxQ
grv7rP/xCPNWRdDwLVsLtsX3VXbDRAm5SX2VGMAJa8FWlr+I9qU0gUrrLMbwWZXn
rhHzcX/Vim4KFkIRElACFXy/nI3aJ9eYoHrhCdXJo68df/EzfuVao2Tu3AhcD/3A
br1+H9isbh4B3j6T8YZ6ICnJuEfvnStenfvuUyD75vi9iw20Ei/IIyd3ZMHHDGeF
DSGlfYdRQgYT5yUUcPZ4KLx+YSS4HDfn4u+vAJs98D18T8vSEknRnMfP2bc+Xs5D
v0Xh/euPsZQddVMNlFLADFtRLtKL0WmEI2ekER70aLljg1PImnvuSo8Dwmk/fEM4
uT45WjzGMk0Gk6/AUAmPuPX4+ju8X6wBSGDYDsC4zbpzrET05geKU0vTTG7zh0y0
bVv2Tt+QAB6nxP4IZ8Qd7J6X9ZwYl5UM6nQibRMlR2GwTkTIWAAbmSBnAybkwY8w
PMod8aRCLYaPkTXuZQB9YhmX42Q/re7wKpZlENcHbjH2pK6NFkiB8bTzBMQgFxUM
b+zuznNAzCV+IBOr1q6mX3rnFC4HZvesbLytepZQFp5CUXkTdA8aEm11YofwC58M
dAJ4F7OGwNuRQVDNTCeiG6TQjqO0qM/5oH+Ie5xlW3SitVJeH0X6jMma7a6+FXgW
J1GDPzvwfDkL7qL3GZppRUb51NbEl1vNs7L4Lg2o0dU3sGt0HDOR42Qg9CT2LKBM
LxPSKLTiCoPmQ3ZfS5js2uwqXksQ5D7Uhqea9FYi/Ec3XW/HVyGqOShnCwsQ91Xz
CzTpVrb+uQCJOW1uymkW30Dj3CsUB3Ksi4rZBH9FNloY4ITbtz2wItuk0SgWtAA3
Xqj98T1R6IcLgmW1UKAL9Zpcrx8VxFJB2XRvpo33bGe4pBhaCchogGgV1VFVont7
x5ITrwHDc+wLWwLNw5LfDRs3q+2cg8RPltKuG0991SDavrQSsdqbJHRmfjuTlNRF
9nkY/lHCs3tE0XcEE9soA6rlOryA8lnMwTCAYdLuwiQuuyWYUL0I570TMh/Sxkk9
opfM7jpDn32Tr8mIxKp7e6Y7Kf8DvdJOuEiTDq9uOPMZqoMPjYmL4teq4EKXn+Pv
mZP+R5Y8SdLV5W1Sw4pjLt2g8+ISf4ycL9zNcB+z5t308NoX9BHWbaOr3J9BCCfg
+9I+yj4JNNugU8nmWk+JWj55sRTgV5Du9bYErJtkdem13mcgulvI0AWz8yz7qVnd
WrqT0PK8DRpT8yPXGj04684MVoQEhlJ/wa++l+RPZfmjNAYV1gk+wFLVD1eujezs
KD0f6zLmcddeCn47YUv6LOAncUO51ZRVR1Cs25pwFKcSCzooefYeXXMOn+JwGx9j
n+N8zLD6H+YQqgvXwvRZieWB0EWR17mcb0FphqM+ebzIzYZrswf45qJ2NrYG2jjY
sz+7xi8XFkE8w+g9/KgUWQM9lVhfEa4g3xWiOackAg6s74hKKABAO4GklRviZiA6
W9IWtX2FcMLnnlWzc+dMpESWivUH71eE3dG/tEv6yaj3r9TLSKVDQo1OEua676Oi
mVOZLtYTVaMCu6kkwgxC2iAVdqsnefHBG1DGRAReB7L7jh/hRHX/lgIMMmgNMkiY
bbVPElvlTimW1LscfxFixNrtrMI1iWi7tUsKRuvlQ0ecwzwYvC9aNcYMTfPTSAoJ
jnkNWpw4+BYFTjIdLoDDPGAd6dUZOaSIpHRDfLGjBxSpw3Eo2kg4y92nxvwGJ3Ut
a9MEsTsTcTUzCqISaO2J0JkNPwzl/kSzfio+calhLFMhbbK5VcE9vng7TWDzPWFt
kPim6+Cm1Fzzhfnb1VVDX7RKRV6Qxk6nPjTR7UdFe8QCbaHd3Di4n1aXDKj1h75T
jasQlcPbpJIIZRRHkuleQi5zLFBCL7SytiA7weS3mb7XpRl64VbB5Vs5598suOGc
Rd8q/gVZcdQL1G82M3VZ7ii2vOyFdr+jRM+FWNpX6245FK9Jz3DEqT8eeY5ycFah
+Cy2aXVXDbY8J+mM8/siZUaWfjHViTB5yd8KjLD0uLTbCBWMqUoHd9uAlcAjhAf1
FnnlKwaDviQNBgP4qIAfKzPGh+Y8pGB2bQ1nVIKGqLFrFmJQpSkDsIWpyg9wFGan
mFdHwI6PAlyxrUPsRKHj5duRGJaGlKYTB0Osues2p59+WnMDYDgP3aB2a0KZRMT/
ylLwiAokIXlGFC8sCOQ6GfHk6EKx6OtYHbFuxfKwBbKbhOhZViy3Fs2RiYTBq6F3
w+OwqOKYyoZrqvgEO1fgQ78fq9C7Hs6THQiWuAemgi3X547EnU7W3XbM+wXHOPGy
4BwjNE/hPT8rDdEVjPUvI3V/yAyiGtv1HH2jUONXYkQb1kyI/p9wGGuQ25wIPBs2
UljDfsCDCIbrAOq8s8KUM9t9eOfk2QKAhbLwau2KF21RZfKmjGDgotNSe0lWx/PK
9k05JxC5Gnw+GKr3ZrB7Nj7P90ueGyOz7tqeeYQXdKs+/OvT1OfS0xFovokdi4XF
vJE6VuHYZCUCqzKV2it7jkxJiZT+tEIkCDXpYQN313f9bMtu+05akt2auVGq0/gm
MBO1IhVl8oaYWcn4fXIwxBn7Vx3+nB2HvM147QuP6N3+e1dcPfjXS/Uf2YziyDLc
v5qZYUMC+QkntQOHPvfAfnJDhbvJ5JEWAVCdZ7aG6S+eoaUPo7U2TYy/ntJel536
xTQbfymPMUj5otD0U1YFtuLrSLxJ01U0GmfJ2SB7QGmZ+KeHMpJaVQZPEw1JZYGG
wKPSwHEoMyjewIG1a7BqKYdzFpb7/3sMNuMkEiK3kH/QbfTXsXmFn3cyVSpzOo+k
I+Mh9dRggR7brIMdpjQqhnYJ1rKlMdtv1oPsbd7xKyr6XAgB4SJ9MDh/o23pblDt
9+N4y6jx8HLX9sAuc5KorCQIKXQ/5wq1DEPZ7Nemd9zSHiYHHO7C2tagGFraOhN9
Zc8fyio1iBra4TbtHrHJfCkoS25XqzDj8b9Y8sJrsjfY2AiOiCHS1Ho3QABsZPxT
BekVoy0Iv20slaKFnSP+8pWcf6/MRVG08feZNoe9D2MDfwue0XNlutxkWLV9hiDN
foDCkgRvF/JKV4c0tN7GY1Nbz/97c9qGNzabEDCL+T0ryKGXN5rzxJkjwsTCfEYB
bsLvCIfR6Z0WsqW/gF9z4gitnVFNOEOp4KjMwdnVZwWzXT2CUpg+JK3xCSe35Jfo
vszzcLfyIoD4IrdPeF4PtU0ytGQ+jOBallAYTfsXMcaufkRzta9DXa9Fi7TiHNdl
Crp0qHH1lD+mPoErNJSuvWtCYvWC0ssajc5MFX0LvP5xv3GRT9ViLSA7xyzLiG2A
EEXgJlNLVCTv0iAucfuZDIuvbpSz7XqB0zVmIA5v4TVS0P78ZXZpKtiP0GsMdD4l
Z5XERl6GYqH13GdUmUPRKUB4x7XIUD6FaOcdd80oZgB9TH8Hg/Skr5fxz67xKEwc
DARD+145XNBcbHWnQbVrRWXqh0m1yswIr2j9ELiOqhM+y9Xkw6Xr2ulf9hEWBrqd
7+7RB7N4h3Jifz54AFInmJqIcdvKYmp1AjmWmaHpIrB6Cnkn/UjZCb24Pk/mxUrh
sRepxmqEcv8g7BN+eAzLJuKVyXBaZ9dsH0+nCTFCFeGMzv1EMgVREKa+8uJw+bdm
7BeW3EtWGMgR7eIIxYCXMpv2Fp2Q36RjEwDjum+Gt2xXuxW3gXOA6aFl6zhB5FUw
sFUjzCmkYHeBPFP+UsZid3V+DSR8ZVpKvalTsT4BFhvPTSUiLHz5o6y2RMV9k5Ja
cexX2z4ufr1vfqLZr6r4+v4ah50Cmvr0E6vO1puxfsNHLVunmJK99yqxdaGz7yJL
Cz5XTbsvb2/X7pMmnzvRNrB0qUy/WsNRgVmSj+wwhdgxsgt2mdEik12la+9NW2Ks
5WGZ4KegmIAjamjYWYekdHioq5hLwMknvh5cZyR1BzUefW30Vpv5a/8Q1P6qNv5X
RdEEhMKCrvAsJG+IEhD1itRNBujlrWIVZI0SDuVDygC15fowAXHSvSAWSaGtWMfI
yqsdacUrjLdtCzL4SlWlZXvBBOrdRlm6MdCTFR9nRrXdSH7q1Pzv2P4RTrOcz+gK
oBPRpoGX+NdA0FBXiqrPVVUeakDGZuNO/F6AIBmbJy7ULZM//auyadVsWhe/q+DW
YQDuRlozp1NpF/yprTM5+22/FMfGtXZ5pSAGg/KcpYAXF63AMN2iOCsXE1T4d2fF
Hzk+NQeyZrw/Fs9k4BjfRSM2OxN/oC+GFraD+GC2N2iYPK1GNS1OpkGmQ6JN/vOU
EbKdcD4ISFfiP3i5+KSMRzWDdqcvRbFzi1vnIKQltwFAMESu04ux8XMlX0OK/L+Z
EcNA20iizWoGE+I3XzJh8cJmzY0+ThovImr014DwgU61Pa0AOc2zkuxT/CIfr11j
JdB7rCatKsCWNCai4nAsjDOo37QbZqSjOfiN3Dl7xwyv+cIN1yPzjtMMM9TixE8q
uYmme4W4a0LXtCy9VtaTdPL+Hdn4zsdyBKzUGzUotlfLbJFrUAbas4IOLQ4gQAmU
TjMFjO3H+TekqUyaVOCE/UmIGQtTjIO7RA8pYZ6UfokSuhX9i+6MXX6Q5r06/X+4
lXpJDBeebkZmIMJy7JFzKC5vQn+9g1Se/6nA2xXJ4f35h09jrdjl3iJu6/2FurWQ
1GV+cA2T44OrsQIujC0MTij7Z1STQTujjapbb2ouPE435VQeacpcaKjsWo7+hpK9
mtTtzNm19gqdeD+ZF957jz9HRnOwfGZgO8qPG+ThltTD4jyFlzM3dAHuIBFSHyye
fBsYmPnLlfP8HZ7jWPkwHevtCxQDAGH6InNfgg7qKX0GINMcAtyT4RwylVirj/sT
IWEltUX1eoZ4wQbfwkhAtI2kMmnDqfFfvOp1OiDxBxT4Z09HDB9u5JMf38w5zb2X
SG3inUoSQjHAi7BGhJP5cymUSs9tFW5iZcYsPHN+9bOE8ZDKoqw6SsrKGQMX0bIE
PMj6F7SLuCTnPJtjJsVMoBD1OBBQdAFaCU6GtRmYib6c+dM9j0lOxpvaGnFytmZB
K4uGaAV5SGuO5rGnJDC1LbT3oWgtioIV+g3hq/f0X1GrTRWv5dHa7/TW8qGM9QmU
dfiH7sb8DnpXzODrOrZLb/xF+fcDA044ofxhP+0JmbFLP5big/pUkGA7+EhsqZiI
u/VKExoRlV31s0PKAR/uDa8h6a1lo5FSh0ZxX8wZC52+p5KOFkvttdT7iHbLcm3R
6sv+QMFGDfBKVMTm7h+Hk2Xh1zZcpx+akiOiYYAcgwP9L8g8jZUnZ8L0Jf+rhDsV
NqhnxiHVf1kvB+Tuu4nQCPc4ytvKajj8nGACnfNe2iUkHeDcBJG01zTKt5C83szF
Dm+Yh1KYInQhRFb422Jnqco6aoCRC3VhvHmA4OELdb0Nr+Y739M+v7Eql/vmcXiT
UO7pcRaFrRKRmopdgWE0yql9qxl3vEZRQ/Z5zKiO7qCAOyF4do62g3f83ty3qqeT
nE2HhfJERin+takopy3WE939LyEYmvwcIBGUqmazSN5OLswXkawkNN4T6VjjL5tt
1jtHFITBDHUNf1nsDjrF/M0DQNYkQRZrFKY8foWSkt7haVwSdOeZgForl4yA7B2R
QYZliE5OqsF0n3WVrU8KCyWdGKldGory9JJtm0UG2tYno+QKQtBSynw4AW9ttKo4
Jj9I7jnFRrQ3qCN0D+fJpIv5uO6/yDiAYk770cG2KfWMbHa8lRsTawI42e656ie0
w2c8CiKBhIRUjk9nTv3r39g9ZyT47lfs21fhFcqoMxnQCRXOC6zLvwUFP3K9PPKV
cL8b9brmUzEsgtWU1gFWqHfgmMTBaR0Xwp/2IZtLRaLvY38uNp6HTj880j32zI5n
/Q0WyykhvcQMTWAUQMuUEKMa28xMGP3e98g7t5wud23/YMbuup7KS8AX6UQivzsu
59M4MT0bZbBPDjw95U+CEqtEsgvbleAftLYr9KBhV0Yn3DfplgFVOKU8TudZkTNY
mPNHjjFspCz801+XhUZPMfrrdwQfAd3qq9RcwHr6Iu7IM5Wq+9I8rK5+Z12vrdwL
viNXDkoIuTjXPFEsQKqH2E5riOklgdNi5UW3lEDHkCdcp9ce3+6PU6ZvNlC1OnOY
HjhSW8FFCBqcicAriiVDlBhk7kYn195dO4jI2/LLNeQdzJGIWu4hr3falPYUvO4R
5zSDFtf7csYc464Xy5PA4I1HUr6NIp/A2IoTSE7BEp4IgFo8NCVs5h27rYkJNP5D
UJ0fEUoVLOjCTLor51MotiH96xGHLGilW33SBUY9GrxJ9LNIi3g6J+2L2vW6vdus
r4qstKw20EUelYLsB6JW7Ac/Kcf8sm1LDColIdEm+VMg/FqSKIRUpx2H8Wvr1Em4
5yM6VIR/4vYzpijZnQ3wGPz/HI3MTBj5Q/7ma81fraibMATTqbdvZPlJEUnkLzv1
az8YK0DMD5UlsRJJhfNFE006Xujq0zm3ws2mcXZ4JL92Ou2xLSyus5qejTIAesLH
uVG49N1zIBGUOnwLveXGR1/YaMphLx+/yNjcM2XMVyavRdCLq7w95VnELBnE4EVd
q7sDe5opl0WyXRBSb4v4MJAuh6TKbNZjhi9zaP40mJcuzI90Gles+QS19KlSEowS
Sztpru+f55G2ijx42Qjg6qFIj+zcugr4hmwTsU7/S+UZQD4/Z5jZ5RcqMzQ6HXw4
jLjJwK37zk2M+ko/YUdpyWd2Xjvao+EuloNlDuwAmkp1bV9a/ig/oFoqGKgCkr3b
3G1YRNl4RttLpnyuZnxljotFVB/QEoiZVfGlJnMFkftaUFFxB///7xIrrW8aiAD/
ljFnN9X5HDG/PcD4hA7QjnX3F3mR9JLTO9ea3gdK7vq7S9ki+grymXMC2yY6fdOr
P5C9mIqiEXL4J7C7gS/1e6WW9PPsFuC+N2kugtZcPK6fYJjRRbeeyyO77HCABQVi
mdm0Is76eH7MqP1AK+8ERrQz2DlpTYHtcyWEzQt8aClqpuLJbzu5CHYoX2TvLtJu
wKIW0HdxjTQfiYpprtF66lGFSHgUlDffxw+h/T+m9QLdTddENtJUFcDizVxhy4zt
cnWrZcuR4ti8RtLb6KCcY3/gm4xaZbWpnai7su/quc0eMfjB6gdi0W6/KjlMr5md
imZ4ewDRiM7toVx4EwK1k52rnShN+QKG2FKvpApcD9EglU+Vkzh9Eq9ISAbvhqxo
0HztOYaHPVObTH89PqE6nT9MrX8DIPeciwcjaO0ai4du9IXFPq7r84PsNknNSUne
48fiq6iOym3OQmktr3zEFMEIdbm9+OWo/+Z6lIs9pB/gqqxkyUYFzjtrt8h7K2On
ygqluJdCVrXuWOuBxXibr9DtByen3O3/avGCN0Q6S2zu8dxzrwpx6yTOgjzCsphR
79sYfllNsdUIxO48rk0jsJKjTjYjtWGhaW6fMQvH5XWqspDHCXooiPM2toJIxu37
zrClW2Az+eV/86fd0q2/UONNQ4Dz5sXbPOID4gHl3S5g+BM5z3FsJcAICatgJoW0
UhdqZRxDD+UDul4uvpgDdoErgesTKEUCj194yCYT7y7WzPiAvVTJoUF3OQI65DTp
FmBD6fgQap02ltzSSKzbad7toPbxU28D7agqCKK/vcVQZE30IJ/5aWnVN3FAtXKS
dxJB5XFFvy/OGu7iMZCC5BEIgOu7oZzhqgGkmRT5Yqntm1tnIetbNCe9cDFqVsu8
Kv/qiGOFTtmFUiPYN9y2dolBVA6uzLLKwrus/Khylfq2ndsb5rS7utM0G2Y/Izgh
Q4ticJeD3hDTDqON7Pj6y7cTvsC/XOSvLFiBozkRgSJ8sZN4OCC2xyp1yQtL8Tmu
JQ5Py0Z0geJ62Iu65ZT1cF+I9E3dZCjoALDjLONuOG5hXNwVFFvt5E77tV5x/Tjb
VJJ/cQoLZr+eqpl1aKGQmelK+PXQ2at5MM8cKcTzJ/IIq0hu7D0dfkGwYVxz2ily
yRB6fhbNhcF2O8MF/Nj/gdhSR3NcoGINLbkY24XdAO+DSTQX+MQEid++p/V8CXz7
UtGcJz1GIC66hr4zZo0WwGk+jFJWkyIojMgFyZx6LGiNzUPQLy5ooIalG1bmtFx6
YYtRVoeflqKt0RybRnztcwO8ANYlZvpTwjXvOGCAQft0EdjRmLD4KLMn6sJFKU2y
oNWRXIQHlsb08bIxjBGPnnrDISLCZbtMW7n3ReQ8cqSD4WELs4wIGTYoliDOjgzZ
JNabV3nqSNOYY6X3R4qBdTAp/CJ8CJz0XbEqIR6q/4x0AeOwEy3B0VsVZvDv7xmJ
IY1OiTK7oJS3Yo87AJyyhEu3q/E88sMtkqsv/mThTRGy4uuVB/gMR3q4a8ghvm5u
o/sItyC1ueff6Pnpz/TUSMxaW3k+616Rq8J6Hz9vxt6XnDS+xzpfHNHKGloqsRj3
hz5bwoKe6JipzLHYwWXdHsden/KeElPu8V0EqgdRnvQPGMB9/+xHAvcq9w6INrqA
RvX/Y8AgrtCRbWeeh+/v38RlsgxLLVVpVk67y2aduO/PP+fRldPbGLmusg4tWtai
DM7yare/f1v4BkCQhzEp5Gz/ztJJmE//d86Fw8k+fCYjvAzQslqqtSx3FqN0CBGS
lzUNuYcfYtRUGkNY77vtsPlaF8XMcCyxhE1qagT5Y6XMoDWXgBBCkkrM6LRTqR+f
HOrlc87Xdlzf75/8d80LNfyXC0rblxmWyng/kdPwx9nBTTAfsS1xK/MH7M1tAfte
yaKYJtFplOTdc1m4oaU5BSiaO3Ks+XzV87eyzdJWrSMiHpACVkFc/YXvoxwKik74
C6ZDkvMjWhAmvJLehOfjjGI/hLHJGHP0b6l5aDvOJeyjIna+nz30fbxsrKQLtLH5
4xkbqas/unbTbSiPPfmRFf69h82KAgw0OvLRd+eATumwpY7E22EwmIr1J5vnZATs
VlecgwKQ6ChbQHRNSiqIgmNf5HcAgBBI3YcFK2GMJOYaBYlHd+lnVvv14uFGkgd+
fqedtRGGAUzLS4QTsGXeSJo+yv1CB3/k7NZsO2/1mXYMyUik2/sUn+fZCYij3AVW
eDgbW7HT3pDsy/tSJNRvjmw2ocbZ1tkLUiJeUql91YW0zU3YXY2VnpaaygBsjIRd
GAJu1WxGKEo2crTmMiztNdJc/DiaAqfrg438moeVuYpAKX2QHFGexzVZ0TTqRz5A
ltOAz3KU+t7SZ4p+ss/hsN4IyVCAPwIJw/OyWsTOo2r+ySQleiDwjBvZdUtUIAES
KJomfYiGZmBVwUt9Ln2nqQ5D2xaCQEQF58Ai7vVGIlb+WZKHfhOz4qL62R0U3WlL
0v4aLs4ntD40u5VypQyYvNcIM8Ni/Slo1L9cs7b1Hay5rtk7X8QXOBfd72S47fuM
AJ6e3++8rpVBMgc/xUgmIBXZ1u3wc3/SFks+TFXIIRfjhuvmBkNvmkFtFk7WrxDx
SQuLP3ftwKo3ugE65TvBb0Q+WJIIEnBuGZB2yhSUMf0ffyXZJDhj6E0WCW1y4v/w
2chpyO8riCvYH0w7PR7LRALtGLUqRcwb0koxQrr4OQwWZSo6mqkucNd1BaoqtwjV
3LAGJDW6ElF4lPJzAkCRTeGKmAdrbu7nD4yfFY9lIow+spKQnZ8hudij64VuCEw4
KOhCxgHEQJyuf3Ude+86G5ce+xUJYbpiGoWhQ/H6nBXyigTF+IB1O9sXveGoFYs6
+ovrV1ZS+97fdOK4Zz64YHBp52KyNS+xQ4imu3yn2Naym1kpxeSQokqHe7vaQ7w9
hgZBo88UnYQCh7o36I7k0Gl56kownWFTdWJoZIm4Ma+5Q4dOJ9vFKHiKtPoPeLfg
S8FNOA4hg0NWaTKP+Dq/ONedhP+5ZfSLCpv+CPqx8ph6wmFujugREDbbUZ4y7Jqt
WNpnM8SLjkiHpIrIIOZJW3Sl+iW+0zXKmXnURV+W/nJU72+3LpWHK8SKSB52NFlO
Q0hdA59Ijqwhm9+NRH0Er48Egina8l7sj48oHIFrQQX/cCJ0EhhjIErVnp+uG7n2
MxyJ65lZtMtLIGEX83tgpf9i9bjw0G7x6qaWS/vkeBz0A8sdnUkH+3nV1Luj28i9
VT7jBUJWcCduVpDz2GzCmMswz0DoUGwUUbT+bfPKW24JvvB+0Fzvzmu51XSX7FKb
xw9o21hQDAZOf65mAsdsIoAbma/Wsj73t7LH8bUox9KEMXBcyN6MY6S+uOn0jsGL
CQu3bAh0oe4uqniKc/twmRyTGZ2Yool+m6+VAznHryewhxh20aDPtFsaX4eGSyVL
ECUWqQ0lrIiMBrKDBog12XoTE4NPge++4YeZ0feR6aghXl2F5XREBaxvEV/FNmrv
y1km2WBWJFLQyftY85fxESG/PZ2z5AsAHBvAdPZLMdGXB9bvxd75Ytj8hQs2i4MQ
b15i+/KW6EKlgYwU00/lZxuws+9YJkPoqT7vT1ixZREIUB1vmH9kWf85OeNMTycb
bFGlfzvbtm0pRXqt4dGQAjl9X7Cc+fWSWiNNpnU8Ke5xbIFB8EaVcDN6pWSeeCyn
fHaLLjFNHZJyuxlcgM23xQHYPPfxYzY03z4EC+27RgPOwKqZ25IDe/2T+ZX1rLDG
u/zmp/csFwr72sD0y2HwwDfhfDeLIyUCwriXuHwwTEOEIAnTRz3blaLif31O4trg
6xLAFANTNGbLXe/tQrTSUbylv4qcmwTEN1gckFJ+cBAf7NkXof8Zrh5umV2e+pVR
NEnkqaPLFMV/LiQ5qLsPPrQgBsVYinXGqi7iKhcl3KeDOq3pv43gh+yFsM8WWGtW
qCF4N4NsPXLZHdsvIBRHs8xC80vU8ccpLqQ4FySMkgvyKUlOXue7glLbKw5JdmLK
0boEdKvQrScLgsjzhXIyT5lHNs8YDTZd0bltmhpu+nPx2nnbxtlXVhdZKVLuRYXm
aQDD3TFYSBmrWSfuLqvaojTKeiNoYpfO6QAoh6SqH22w03L/qK166B5gGEQ1vfam
rg6hnnyjIqTUtbW5YAY0+11xySL1xLvvhlI7f0BIAiH8mU50QiROeWBdsSQdrMsK
Z6v8SXAVGiCECp0Q5QBr16odaH0Cdb/pxcImRHLYQ/a+OqIIMqsJIPMStekuzx41
PSUVZLj4uJr9tLk4DHrbbdk5c9nUHvKoGZVjoqh1VYeqiTAmz4rLw1rzbxkrsASI
X6ACOevHjl4v3jdC6VG9FGdtpqmAmO7cdlzo1ocnmZUjpRZ5hHOYG0iAx1ScUFSN
rqrm7U/KeNwediyBrdY9RK4fgJ1kDRUtHM6wfXWalXaqcfo7IbVaOIug3Zp8cM/B
V+YN5OB0EYOJdmDL42DOFCYeacfKaS6mkiCMA5lVX7ROjCiFExw6s3my/Aq1jywj
lyjEeqOoT83rLfFwmL6J8TWrJUc0woCjTsuUbLZdoJaEusMO0fzg8qPgTK30zbk5
/Zl/Kbd/O0XcmBicKGJOmVmxQd5Kz2BZ8cmDvfkX5Va2Y6D/cKCMGaPe0sPYdytq
0zXNR/ljm3KDnYUb9YV6MoJQz7NAksAq/4xBhJxunTeEM5hLzjat8Zuok4Lu/SND
KuiZz51cxCljca+iY/HEX5CwP08DxtCVh7VN/VDW5ODTmFziASfL6G7OadgAxAs9
VPOmfqpXZvyZ8zbHnRpuy0lNrL/ps5pv4CiR9tfPJPA=
`protect END_PROTECTED
