`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
97UtspWxdW987Tn1vpVp44/ngPCiLNE9KCUjjMFy6UBtcPCPERKhKKSbSRp9TxT4
ewNI8vHShS8vucQMTIVdRwrCOsEswKcYnO7vrZJwFdatFzJlA++eeFT+Dy1ZeZcj
tgUzQ84TCYgKHmXfPUNGhJGJ6VDYS74NSuVJEXSfrHxnSQ1c8TEKO1n/w2jkc8aL
HPNip8tfarXZWpjI9CPGJ9evwF0V9zHazxIM/wvbpC8kv14Fd6KKrA8glHB3KuU0
hRdphCOtcPNkSXtEyfHatmodwpuKuLJD9818DHSzr63j0GqCooW2x9jdUF8odt1E
mwP7z88bCylgtKJtQSDQFaG/h7Bvi4jS2vhuSWDZLlaW0usuPGH5u26BTEhJqR3l
sCnuoXt+7rr0jLceir4+SA==
`protect END_PROTECTED
