`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KJk5bYxyiEsowFuVF9Y+emiVzu91oHNplBjYbFFWDLZ6DC14jh6WkkqhEWsIw63i
h7uoOEHcP/wrelxG4IYA1vz5HhDYEv8JFgj03qic9IG7h9Zy5fO8bAM7JKKH9BrA
lIGtMpfaoVRTrWSzwprBR6mxRw5GgOuVh0WWep++YnCI6mQ0s8kvxS3cnyFU6o9/
4+xSoEJI9K/GJtMnbexVqV0GrLcXcjtH72mB2fPYaMnSV385bY55OAPKMof/cC7p
Mb3+NsvvrtKhnCBTJB/vcVvwSLLdkJeWqwGldKUiBZdoWPe53UPGV6c9pBUYRs0P
EyAeTubo1oFLUFEtVS04hJNJSTfhLrE8aaVYoAQXMSb7BQryvOuWzy4nQTBBUB+/
`protect END_PROTECTED
