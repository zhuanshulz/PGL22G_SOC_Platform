`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
awCUMd71L2UMI/OayMwZMRguNYA+L74EpiQK6U7nNNqZgigp0iQqz2bp1OhuG/hv
ZK6qIcXVs02kzUyD3h9w9u8Z0WCyMV5A5/oNr1NsmLX2wj1Arpzw4A0gtplVQfU+
uF6JEqi1SEBsVImGAqtcQiD/32LCZIejcUDhBUL3iA9zrDP7vueXU/5FsdAjM5Ai
i3R6yd0UWpxj6BGjxOtSXvh373FdBiddqbpi0LFwLZE6nXALogIEserie75khdt9
n7bbS+9QikpnBBLVcGTd9nRhQ4r7y0GMcUKrXEJjahGVJ30g2FSgTYILoOMPMeb+
vvcUFEbWXR0syZFnTqKGRoFWj2/G+BJXM5HPJisLh9qsfIQiuM9yLPMIydvAvYKw
ZO+5B30yOKDosOWzB/2/FDOvmh/lQaWz0Avz6LMZxOqed0yovDUtnUrz6KGiv58G
hm84fC+P8olClqi7bEJVsp0oYuWe/aQUl+EPbdYpA12jszjiU7MgxxabzzXKvvtD
WAImxZTmaI4HXCi3ZvZTok6m3tkXQrwiIz1OnGoh3aiiB0TeqeduUbAxmMtD7MHV
GxCjTrFKAHogGvjmbA+yvugOdprs1gQDnBx/XMGOhY5qFTn7FnLF+x+wn1vfbtu/
SLFr1whlNs9btatdoSyo4EdN14W6D5pNW44oAcSHFcZvjOaq1d50okeggbCc29ez
Wv1MfTLV1ZnJviX/FDq3qYBrGw4NZZ73z1PzVaChfzuJiN//lWOVWUuM011SCXQF
yjWs18N3Ctszexe0XtDmO0cEZYRss6BK+Nza+sLS8Tj2A6P1KNPYbZ+iYhFjUiRr
PJtcLuXCBnsrGodQLcZNs8RD8uephJ4bDn7wtOZmSYlhLboczmwdIWGAlG81/HYq
suTYAx6b/mA1DhlB4lLrd3mbnOzK13wA/JWLX3sWPHDoW5tLYiOoLL1aXY/U38Ck
HMX/g4VtlsAHBVU9s/oeXAiSz4Y/o/c9lvoULjQngteDDP+PMdH4Nx/AcqQxpyO8
P5mDSl6O5BaN87ICwTknwQ==
`protect END_PROTECTED
