`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sGLOn3uKgn7Ik8SLTVrI7dY/YZKZhptSjy/Ray98gz53lrp3t6rzl14Ey/R4WCEQ
h4lelBqPwj1FPV3+0fNW39Bx3NtYj0+dhiTjgnDgGs8ElMLLqYKszbJGNJ6n4SqL
w52pAxuUXvzoNlVARdlZH4K225Ykqt0AaAih4IFMh/NWTPCkaKF+1C5bmpQ4O31y
vgshqNrGoUrekq8JxI6HyMm0crX6mcyFrhzjG5P1y7DVQmscIq7qLsZOTMXSgYu5
pa2BhTqTHksMugAYZD0xftYBxDRXHySAikuDCHPTz/q5SpavryY5tWKO8UiTsV3h
HB1qx6VOy4/Iq0PeicGCbSxngqgcaoRIAoD7hnnhTy9m6ylafhbMnk/cDtJH+V9x
0eq351/34rpZFphRLVY+MRuQgpx41khLbiycFTyXpj3npyEJ6KmKaiFtc7yW+hOO
hg90Xav07JoLZGn6XPIAhD9b+ntudpmWE5yCEf5jMKRe16CGicCvwE1T/F/1W/aN
dUjg/NFJmAfZ/4OQI94btg==
`protect END_PROTECTED
