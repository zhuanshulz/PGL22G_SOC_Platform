`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hTRWWnULruB391+tOQdd7uiq4/ou4QERBoc5SykbZHcVy6B5uZnqwpcFZmFFeeZG
t7BD+w/pPQ8XkJeQiLsbaEjGdfsbATmT7jY1ZMzD51eff6isg70uwgGxdwiGctFd
xQB17EFiEKsYGPhvK0WnlFUjNNdFtVAv2zgMhEAEpLkKay2a4NgqffxHPZCcktIe
W0XfZec3Jc0XOiUwEy2p71sto5eCqTpcCGm8mzD2aAysnUwhVsoeGOZCyShbxLhj
hoZqiZrj+rabfGKRvZFUHGzF+2o2Xca1rQeLSN84uuFHFr9fG7jqLKSqw12qRkkx
M1/ZtlFE083CImKvECiB+Ky26ewQHUHm7/ZuUmE0RD2SKsGaxsy9sNDGTH37Icn9
ECXxnio42WDrYRNZA86Bgho2gDS/2x3q2ttLCzHeHsJFqa7KpqHUKa3gEzLZ3uxP
Njs4CvWgBcIZgWpopIVJPDcuEzmiSapz7z43hviyVrfsJuf/GWIMnpblH11gBbjr
Itk1Lea6fYISUBVH2UIN/F6oidFm6amWsYHMd9DGMUJOKmgxGlhdRcqxnK9nsDel
o66DU0YWwm4GefEsKzwNeiK9yrgiyDFpi6MGpXGZ/cRKIT4woRJ1uQhPPWwEJEb3
8KGY10T2gbnUuGAzTfNBYEAQ7iwDi+EuNNnhbx6ctjEID88OdH7x3/XrmBdwTdGU
eTFZKaxFOyI+cxIZMe68DuLHp9FXrcgOmivdCoiysr7oge4wWrnYYrbFbYkd5Hjk
4KUkvwzR6cdC9ta0dX3khJ56SB6LHuHFBqDeQaOr8d7zeHesN4Eq9wsG797tPnab
ZRxsyO+V/Bs3FuOQFkR2D845Fw+f37izqcXjc6y66FXujUWAcyHSgLW4mdZ9bfbt
Zx3uigPV8GiuQEGxyGYXhrfARdvg2jAImTSXGcJwZI6XrN/ivDm7SIp/298jQhG3
R+whDpf7ldj8n02jSsi/4TiIV3Jo3qYjmES8Krtc5VBKP044I4dv3Uhoz084uqvH
LZ0TzpzWNeoKIrmBGgE9OInOBSTjyZS23xSjQvHuwOhGvTmuaxc/lJaWbQ63o42z
KJk9yIJnphDhWPga8bQvV80d7sPVm5o2GGaZEqbMqLW2S2vbeq8ArrEQLHmyV/gI
j6xbm2T86kiDohMqm6t6Q+dTGYfCEZb2T3xVC1MZ3bBrAZKR6fjrmxg9l6MchQ8N
p9A2fneMV8KaWk85uGAMOeYgTkqRFlhINKpKta89FFB/rVTkTXdNei/YAvBIMHiy
XnXtUSIE7do17lCGq4QCyx/0HouBZ4CnjqTi+1olBkK6N3aClrtPWCqA4CMJB1AS
kK7HhnVQhlX+NyGIZ+0hjEySL6mWYYwciitHuptci6XbpgTn6wCLQ7WcIdr+a69n
P4dP0gLloXeajV8eueCBysmCJYbfcEzMyFc4mL6LYs5UP0iRGdWvZD+Z8ECqdMCv
3zjkYBWLSfLg8ZwykOh+m+WOuFQDp/HiF6gQmx+9GiLxQ1zBTtVReqo15I5BajVx
opeBZ1qwxShKvROaBY74VgoKCJO3bV7y4pc/fZ4C2lc7kwtDNfEp64EWYJrAeg3A
r8f3EmDvGdk4E0ckqvvZxctUE7rGaJWKcJk6yb5mmhf7yw4czli1V4SrG8aBx2B/
ONTAmjWsJ7WrWuodZ+FT8pk0pHtnybJVAfe91sBXnoNKUcl4Iw4pfriy6kaInZnT
P3xk4NNRBAsM2RiPinHSndkqxfDGnQYWOAU0Fc9v2thJTJ1U0jso37574TSVBiIU
7lvn6NAgWxwYUS7j8fKk3af3161xkjUNEZTgZxhQKLeFxD3xr9cfY+T5LvLSwoyy
2gLh9kQva5WbP6oXATBswlUfi3+9YTcOKfWk/i4v6pFmR5avhA1zDUrsnQprHOy/
QoHD2dEjxqjiy+fUnALA2OLIhZM5UTr+DgAV7s/vUtu+uMaxQbHsu0ofb76GvZI6
gp+ALFRe0+/Fkh5azI5NR9upNNvucd4g8i6fJpJBLlQl8P3hbnpsFYq1mYurRLLT
IfBYwZwYCC/Ys1m10D6DPlrrI5ZFlugtUYhAFTDOSmGeXATcrTAkljavW01oLrWi
78vOMHzxToHAnET1gHLp0Dre9nzucYWac70/mr6hTzzW9abxy3891ESdF0qNT+7e
na9GLYn8SweQfPCLWneRL0j3ADKhgCZmhAF1vL9mi0dUuyoXcXKQjDCb7xklg8BE
ceoTrV/rAXDIpMr3SqOENQsDVhLKafVLnx70toLkUAUX5MV5bbluGfUPiEkWbEzl
B+LQW6CoH1mnUcbWOxOUI5VwBv+rNAJjf99UQe565Ra5o5HFMOdxv89BX7HJlWkK
srpLIluHEEZp87IKZlgqcLGIv0mPuQ4THSvlYAcIxq/TYZt2u6te90EJhzxtbSil
d9ZoNPQqL5jhYXyPcgNxnPfE4kuW233z4I139NvKQOifSQYlymnTZKiKWyMrjb3v
A33pPGUE7TyXjeHpSDvzOfhmQynqAaNy8ebm7MF3+PaxfSfF6f1SuudlJaguS+Py
b4wiPFWQnXK+lP9+mhMDJMmZ9SZdJYBoTso9HuXm81NGW99F4OMY6MuTIbSFjua6
qPZzMvhRx6ToBCWcFmhu9sxtWBkYqGn/qzIwkNjt9PBDP2DwtAMExgkjwn2C4bY+
Ykmbu6eoGaGGAAZezphotFYx5+f6Jfum1b+cPHXoCiA1ZmDYlj8kay4EQ4xR2aOP
a3sEm3jXAtZoBfhe+unFvbGlF2Bi6bjgZ/MsHVuzXTqA6Ew8ngU5Jhz6EEuFn5nd
W5B9LIbV79b2gOlpmozi2rQZXtZF37INysuzmnT2ghRORb84yuXGfVwiCEZwMgxB
x5Rzi+KBhAmkI12qxo19f5Sipm6VmVKsT3UjfTPRsV1K3jbrbtNb81sDA3bTf3wd
+irh9N02OTBbgOngxlL2+UyR5N1DInKabcV5XinO9uG2NlIX58gSUHlWaefuGtaj
mL6SMVaHZacF/WCpM2RGWc9Ic2cTGpHNc4D+S83GmLK6q27gaku2j+mNseRygOrI
LE0/m8cGU3nQqD5ykAFUvS+m8ATUE+P9DoKNU6zAI8GkA3ganLpR0yrR1pCdl8PS
xzv5gO/+IoyhY5T3OO/luFvxfsjwYsbLh9Fum68abV4ni1oeudSWD2dM7VMZoVac
sV9NhmLqw1y53l8Xz/qTkZW67wWV7mNnKxsuMuE/pAk3CIrQdIG86FVNOxciLb1b
O87Qodl12gInlNhEPs/HhOYVXvxDVjrVcAtzZ6rgJA9kUzGMJt2APo+utDos+L7v
+0c+ujfLvWgxym0LIQTepL0xovQr9DVuVNzWebi3vo2Og1aXFOI/lpvu6AwzeX8w
vzZERczZltMlVsPmP5erPov87LlvSTPC2mpScpr/2n6BlEH7tNxpO8ydS//9m7gK
TgfwZPpBglB45aeLyAJL6ZsliMOpua5N414UlRzJSSV/aLDpF5RPMes0aG9MoieK
Y7GISw/WxLg6ltv13ZnZeKKm+a4XSkGHARFR6OTfGlNQgV+Qy57gYenxNJHUQqdk
PfOh72Yng7ZjWZf2BpNlkvUHuoo7efTa3axLsydu9SBQBS/dhEtFVYqKraz3KbKH
xJ1Eldi+tOhiACvixPK4lRhFa/PCN0MMPRNoW0rwjSKdOWvycbPnxELTeCT7VIAs
ieG9ywFuscWXwSaqNca/ZgUla+wT2WzUYG4hBR6cbt767m5ZNNqbRkj1cIFjcfTK
iTDd0kFn52EHWAiytQClNxMHer8oRD6mq+A8cNPYD0KBtoaZ1E/OlQ2TngY78VuJ
RJfhveDhi1bTP/L+cpmv5cbmdVP4ehTdjmQ6V7gDwGu6plg4dBJNv1RazM2El9Co
VS4sD0+Ad5tfJUtR25aa0uycAMdOh1QUBMN5ZNUOHnZT6qjxz8rHACsyHfw+4toc
gnXCvkyToa+18/gbL3K1S83UeMnNnEB/NjbeJmFOdMXv91k/oyPS3eisPr6LJvFa
72whalMZjA2t1Tgu06QlRtBmlO1Fer2uvAO9Fx3cH5NR2pOAZBoafXLtkTKgowB6
RTmyNfGeI4v9o/FoqYc6KqZtHmMD0f7Uh1qrJYL3XQ5mAl6TX+SCUJge8/hd92Hp
GG4uR5/0LvCYRvXmxMVen3QxC+9Ou1x8LBsvXyuL6YFN3vvdoJPyoGO7k0pueDNN
8bJgKTPhcL6GJ72PZxiHy6yVlLQEO7jbLpR2/pERTHbV7nH+BRUiZJMWHcituWVV
q8rG0q0MepgJAlN8L2ebYILSO3MOfZ0FBChcvwbP+s+c5y1L/dotWQvrQZNOY35L
F4kJ8aMVQIf3UOF1Y/55jLqq9442asUEAOBCldOTCHGuivOLcq2fI7b7SGMLNAXN
/cDNlEzXnKAoUCpviG6+yGAyvxIG6Iy6Jm5CRoMxb6MnGug3xBPmOHLf7lSaKrSW
qyU3Eh/LDvlp0MeMxEakQjDDHz43sS7NfCoeXh2cKJqfA4JvAqMBODdV8VJ+cQDZ
tDVRZXJqz5G19ur8I4PxcgubLtj7ZYetExK0iFZJGKpSzUaDnwgR8gyW/0NTGRbn
yBnH0O1yxLzCbXdn7QcPWk0t+D7GiMa8q1BD7QC5Du9XDJx1PSJXGb/lkyAcs4pl
lXu+IVXQD0TrqPX8zJCmO9qZerrYE4gwL+pchcRgQU1E7NrKL7yPAdB+e39YXnV9
BkTUB4jI6r1dFhwDwKmdJueNt0gnkB78X/eH3Tx17OJcRJkEQDJntyBCvkoiUl5Z
KRJvW3VomAvWlyCSkfYuizD83Gks6SdDEBAW6XazWf/yOCDuHAv0I7uOymMB1/C+
m7G6P+KEYoBO2Rc8k12hvq0EfJGOvVG1TrUp8zkaAiMu3/SaBTCwhQdiwStnuSg2
WHGwzwHPtyhnpHwgNvm1EjvfQsv4p9QbmC2BMbmIET/x00BjB8B/aeVJ+CWr1rqS
LMoHAwI+i23VjkJcbWbMM9wnHYpKJDFK7z8dLHTwPU/P+Gq6q35Y7IEAlpQYP5gJ
a0dbVRoZhPZgGiBeSkRo784njqXSiNBKQ6x8mMj4ndzA7gD2yO3kAD01zQejCYu1
KIGMU8I0myJ/pJuSMLDzWL2QNvxDmCXS+qPTLAnnYnP+Pbiu9I0/kSbnvQq9IBLQ
8g5xnrykKvIx+ot5+VVwgsRYjh0uuy46pJ76WZGad1Wfx7xV/eMmZXuDISykU7OD
IfH6zE26SLgM0MzXB/FLE6yIuk5/cSvefuTvmLkRPmHQf3+1YIU0y6TKbvN2uABY
Hi7w+3DLf/PJvVlZkayx9Sc2BAsLcmlRDYQeE0FDozEWskv+dts2H4xfyUhmxsCD
S1niQXZJvYbpk0EUVZ7CMPiZ3TAY5WRifEIjoKtj32uwXEpHsHndT8P1rIivpRDA
6/eGTfQCkaexmlKBUP3h1T+KE6AVHDDcDN31wgJWRmbCGXsB9++Z5OPo+oW+Fe+O
FAgMY8od4MsbIybv54Y/l6vSIXJjGlQ0G52pAET5OGq7PzNMGQs5WPDELIGiclVy
1SheRKP5z2qC+KXdJRWgVSFi5BlBFtrekq95lPDe0sLGLyfDDvE60fK1wECWVAeQ
S82qtr2JnnvB6fNQF8Ev/OC9+qylPj49rTP+sn12g2M3IvLFx4dmU7AUODCGtVaJ
pdV/gdi4RaY8i5O4Jkn+J4rb51sJaRkNSeksokIjaErt9m5TNvMGx4YJ2Kp8bzaA
uqzkIBBcmDedrLV3CZsAnn7v9DWT2k+5vVnFykmrpmCSA+pp9BXOnz4KAoKq7apM
L9IqGg6j/lpsItKC3kETtGYSW8JoxioSEA8HzEPQ065frUPAOA6gi/kYOkEofr6A
ijT6ALYVgOkFd1lgTyLghGXDg8XA6lDbUhnes72LpFik0dI++RxptLI7TXWsUq3e
v2rwECrVLtCWpoYh6tfm1M5hezFIuhtlOhP1i8aRw1Pt4d9wWcJ1g0ovrtEx0pf8
I1zeiv4v7nYTkn/eMFFAv3qAb4fliN4LVbdd5qFDrumSuit5rVLSFqg9nFcIAuX1
8S3g55Cm7QPE/ERGobL1Cv+Eu1Dyl/9iMyA4w7n2kulfONLZRsTOmQ9z1fb0Ymz4
MEai9A0fcWnlQMJfj+ws5F2ei+yIYfa0yRgbXLDF3qvO/ViXwVcREytnguiH5qBu
aHvNvNSmWwTf9tNUYurda72shS33YjY8yHSadX+JYstfw6WocgcA91kG18SvTSHm
7lACVkuHZ48zU65WX0S8hMs9Uwa5f7OqcbsX2mQ4DHqT7MSr2Xoh1c0r1LjE+GO6
3h1AHVNUftBwjWkHPcK1jUlP2Ey4EeRq2JQnWnmIlA49W6mvlYY0Q0HC0yqyueUT
reEFDzP+b+60GmdLvYdRqn+y2ycho/KTWyqGCWdjCJ9GzUidhuQjfaUtYxKJGev1
bBomj48azNHOaEYdDzhPXx9AukCECXTRdPT9czj4wZ2+ZJAnRdJ4kjJfujM6x/Wk
ZmlbKeqP+sWymV0cmM7l60cjYl6z10WEdOcZrYxyuuDofzyruwGGnC0oVc7MWSC0
K1ZBR134ZhBQCAlnSDAEDiMLszQb4DLf2h8E2eSHDvqr/hXQ2+hu5ZpmDIu6NFUk
YGnKgdv/twg5+Mxv3p7kpTCWu2psSFP6kSMWT0kpWn4dHL4/1b4l3fhxSyP5uIVb
TD8EtoW70eTohAaZsEPrSE/274ClCcTmhDQbcbXGKtT62wbLteFoxHB/Y1rRPWEA
l1c1KwZnXusV73JvRO1dkZbuynWFnXmFjcYm1/C3bJg1xzsfAFQC96DkzVlaodG7
m8Md+x6Ky/kGib3lRbJI69LmsmJ26FFETZDy4cfnuecndmLBiTs3zATanc8pp5Jx
fSWqsMR/sMrPYyqBBRRwF7W8fPIUQmwxX0PE5IX7GFspEwenISX83TQXprY8pIeR
xLeqOaSgWwAK0TmW4JoBgYUdeFHpVY3H46bX2DK6sGnMZC468mBM3xwJaL5GtzEQ
P/V12cY99s5YMWckMvjtlCQdTtXMe9Cpz2WShC0OqWbdEUpI6d4e6elUpwRZi7xG
bNLtDoi+Fsrc6iYCCJezb6ephNpFA/9FSsUR+ZJrjQ5qrr1MWjOClaDN5h0Rw4Cn
yrdqKIJW84QTYwXAHFaiiHCJK7crZRe3pLW1VenHjx6WQargySJ2KkHdF8tp15fC
WVSDgHyLQM2RoE2Xlza9kKSc1L0I/kbteVk9XCwc7wmULo7ThXvO38B3NfIP/4fx
ALmL1LX9qUr0ZdhRkZqlsxjEhRjNNvx5oY7dGPGG24FHhrFYXN0o1FqoF6Qw3GRd
dJ2gU6knYygtNQkTFBr1bYIt8Eu9Kb6Yo5Mn5AVdeH0v6tcfG9aC5bYChRMihJoy
zO3gk5TIJxv4Rsi+hruFPtuQKBMsmIHHinjvALhaBqGbJ2Y3bTLNJ+64yopXbpci
n+HxdYsG+4NbvJvRtlc+1O5EQNsgvjejwwrq4DgT19EUHsWtfArBTFAYfqopMKSl
I88O4Bh45AJhKmfDFJEYiKYB1A0P+drTAtPxue3015sYjTxnSTFDitUsFAPmXZ9t
untHYZoE9eV5iLm8ohiaYECBmUut+UlI+l5/LRwJOtU=
`protect END_PROTECTED
