`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UK/rRGaIQe70c40zSELjjrk+xStT7H/NLlrbvnF6M9fNADxlCHKgMRpqQTFfVFA7
7c2gfKTaCGbjzn4ZOUTuVPuJUd6RKDbsV6/z8rOPwrPA1dJ1Y5Atvu3YNgaLGEkm
b6D0dVsiUtzDrQVElN0HJHsgJ4AjY0fWWXXZiJ6gcrzotfDsEbIgrH+uInuoTyp7
82NiD2ZjBv8ICxHJ4HAqkuhaY+y70f7wWTBu8fTSDaoyXRDTMHtSaQK9hVfLFtT1
eUyiWbNL3R884EbWxl8Id55VH0apx7fh75Hy5MRBnvg8XtL6BKD7gBm2J6Se3iwO
1dA99rx7lWawLmq04+yfJa4xukKFXikZLPqXdmSGP/hE588Pcd1xs4P29BzNJs++
BizlfrYVPDwEse/42niMtU6culo63mmpZVFaJEn0J4vbKatUkxc0wrOz1HTHAAjG
7zdyjrczYVO7uIuAC+xF6r575TC+7SucMdoS3rKhy30+NmiZG7aBNX5ivVwhNm5J
MpCeFJlbVMAAKHaq4BVNYCLyL7Nup8UUMnUIE8uxQmiQxFWvjnvjvrTmjrOxto9y
5LleTrGmGuqxTaa9q2+5nHfeF5jH9RY30UrnEcjuJTAP8VG5XfxEOgWraTQ3sUD2
XZTozlYFuFXPtyWD88L6ar44QddAWrcYcat2bozcTQlt+khHboJJjEcfNoD/bNfy
GXtBkNRlUFKY77UC2bazWADjT/IUUHuRuVmnYd9XSBG9zInU+NKEptOxorVUkAzr
hg8irZilY+c/VF3Q4+4cTe2gd+qSrVQrXUX+MpI5myr/u8blb3K5Zcly6J9sAnR2
2+8ATWdHnEPhGecCnnkLNrkPHCLouV5sFO1murQo49VXpqA30F0twi/uPNlkJRBs
L3WnBV1XSGVtfj+v7CPlZ+ewlISIVRruilZC8D84KF9Wko6xMh+ujqLPvncwReYj
t6HSp3ychcL5n/64JxSsp8As/HuOVecpOnYj+8L6y3J8gHcZG4YPo3FdVadyEnAW
ysmdkpe9ZQhgIStNTycyrEnDDcgus8zhaL9Qpj5lM3DL2ux9XMgKG01HrvwVglD9
nAy+STscGBvULSB3PaGC4ez3hogk1GcyK21aHdMzputzaWlDI9qPJd5IARQR9BMw
x9avRkhD/S7JWb6H+3SwRZVSTgTB+rAmAi32y9fSN+d3LFy3ZNwtrzgS4luPVixY
GqqyOJ/r/GMfRiLVp7sM64EQmLNInJWgUsJus6qGpD05HS0oExJuOdfKORRln9tz
khBuRAWtWatZnbJ2HMUXsm3e95quMK3ovOaVwrzpprQ2GvlGYDYJFw0BKSoS6Rp1
syBbIQuoyP4cLp6MF9Sca7A63hBM0XTucQnQC4oKjlNFNwuP4zfVDahAD2t/WpP1
ifJwfMkDO24OtZpJ5a0xFla6BfRE/Ef+Esf+fY+kZ9+7wq2MrdOiuXEFfbQxYJwU
KBrEY4QeZDG7fPxvqvC8jEMAeFlX+74vZGPGDcPNdpEpK15/kdFwSkR+InzUI0eb
iH8bCj62AaDeUAOfJrdYep9UMlEZQc+sLtSxbf6huYM3gKmLSqJjr+B2cmckBQV9
cLEAeQ3lJESF+L+1KW19wHOjgUiL80gpnUnKHO22h8oQ7S0PShhllSepgD/N6Hqt
IUHlvbOh3FV2T8AoIE9JnqP3uFlswU/rymMD2Kmp4uneKNq8Lbtm8E936XzhcDK3
L85ekcU01zHh8/RghIhMe99l7l1jF6FmOFhubhyQcYjPgQwdyp94tM+fmapJoti4
Oci22e1EoeXjVraZkLvfeJCsODjbsEsURlTf6vInnmkOG4YvzZKPRigoqXIcoKa0
njE8LEPje454z1tAXs4KoBaRjRbiDQBGyQ6CZ1e2OeuHln9prOyVSsIEgRkMSaoX
T0xvfkD7wr+Z/JWDbdWbJETaqxJGNAWqNJL2w9dyDuVxkTzZIjMpKmJWRDkC9m0b
aygpnOyD+JQD2sU2BfAV6MTouFISWJwbfE+SA5fZDJT+OjEh9bY6pP/xKJaeZipy
TV8Ee07M50OnDD8GEBoZD/s8/+i2a9Y5dZ+PyL0NX7dnIEAvBo1gqe9qvxL/3bQT
7mcfdbiK9u3ErTkwkGwmhwNUL9o/C3foZRHTDgMe0Fp/yR1vfB4WHxNBdZt3oODd
O981XO1Fd/RtW1uLE89veiakaDJfw7HClhkKAdjtUc59UjW9SSt5/EQNPt9Y6EWC
ZIar7393YwICKLOgzZ2+AwcqrAAAYwN+IY1noJtZr635Wm7dPUSUV4Rbr9dPW6rQ
jkPF/xymxGEx9TANMlyoX+evdoNQ29aMWZi3/A8gCsZA0q1ksUIWUO8vb/knVMmy
Ks9nYB1TAoq8cAyx0Ter+rQZ2+dMz6tyNzKVCbnffHdsmxiugqr9cVZ9CWKQRmu6
OpLh2bSRCvqauirDxphbMW3ot/+BmODLUL7C0S5/62488IoZKL46nRLu/nQClJJb
ZLU02CtzzJzOg3ccFnlbGIF/tU8AnVFFICqQc4LOv/2HSqxtQJHEXuUcAtBHGqw2
X1qtHd7TBD1+hZlKANy5oyUZlQnwtR+nmWWY5dmq36vnrssbKr+Ub86DGP9XYrch
IAGug7lYClg4CpBadZtIuau26KrCRnKBQOM7z3aY7twqoQUrGsE6m07FqIXsb7/O
tE1mdRwW3hclDcMSNifvo3Qf+/5311X3mtDMiAzG0DE0rxcx0Kh87lmWXvN+9j+t
3brL6opN2zfVKANcdAEeQPG0jAE0cKwzRvErenB6QTI4ymMqT0ZNo8IBzUcpHzM1
3QOOxZk9oCetjSe3veKopiwyhPAqDlVFdqtThWsQgMQeZCQ66YeOLfIVOhJgBHzL
IbYaJMYCj4vCnGuSpcjZMBDEUf+wu1E6MjS0YtUDRiN5GYFHjNf7zqrYW7jWwGzT
FsR5lmv/o5Gf9z3auYPTbEZaOlCi/FZZ+0U4O1Cyva34ilpg9FtbYZAhxwnGB19E
j8mXJbX2M2kG1pwEKr+pss6IbWyuFfo0WpSYWHVunm3+vTOv/g0dL7nSv83IoA6y
KWC/5kBrMEFz8uHLdAZIKx4dIWVI5jb5ACZ7hjxgmFJQDvK82A9whmqZzsZZeh7n
eKoz9ob8kONV5Fhp+SaBR40GdSqWK8mzduREb3IyND0qCACe8e8T0xERN3CANW+n
e9UFyhoZmm+NtNjRHEOeSrbJdrW97SAGJum8F1+8GfoLTO7LZ4MhaP21/FoFouaP
9tNgJkzLZKKWA4qeYLY/7EI6HgsLFNeZCvLgAhFdMtPmB04RyBpui1bjA8bLG73N
DBWLxYRzdGdMRrCv/xGoYFbouj7O6XD+obEFQ74HSWWLA8h404dYMjWts/jUj2fZ
JFU6yYiMVRGV/9catpvkFj9zoDNJfQiyG1p6UW9+aQ0ege8mrXirVmNGd/LN/4aV
qyZ0PTiczxAu07MbyeKUXQ9hGbOeG7EIUNC+GgmyJ7md3YRHcqq36CYQRd20vm3F
gvt76vkkfGAO4q2AXdjIxYH+YDQF43E49klBrNrOVqEBfJoLlHqnHTMDS+cd18Eq
JmStFwg2UvuLH435+QSlLiBvyYdLlcNzcbn+Cri1xkQiWmN+Ffk8R+eut0+Jtlio
dFLXp/CSyEV2i2EYRL2RM/OeKDp6jyxqBP2RjTmv9tjYwFMzZCE6VSjpBNsww884
6bwIOZIoKr1ODQ+DfUB/rPVKMZI9Jvru2A+SHsF6CEHo9IkLD5FwTywHw/QTrmQJ
aEwvhLsAVyLzpY4CFGJLqGW8ADwu6kr01xTQGPTkstTlmjOdq6nMZagOUS/O+l1P
R4Xa+pzZ5wy1NjjLD8Na+3wR7/dpVUaqe7h3jbFSrG2i7JLzYhFk06VdUrlIGQNM
OCYTCUOtZzJiS0aBTT5S0tgsdqQ9ZGkZ/lKW9pMtNh30aRybM5euV3QmdMWF/TPf
7C2A6cKgrkJjYrEWiBNRly6hoFD/qpltmjKnbRnrV/bo8oEW1fPkTQ1tWpn+7/US
7DixKrNXy9/tWMkZT+vndVNpiDVyht2e/kd1pnDESE4pariqcQ+Yaw6873xRVoeB
gM11oKtyVZODNvoYkf2BossxQmGvPJJza7iILe0sIk2UXsg+m4iu/YBR4/920w0h
2cVkFeg1UYUUcsyWlD8KbeAu7qVdPGg3KP9SHdHrRQOiBczu4O07A4j9HzDhP6Wf
3B8HpTapIDeGvCM5g8FAyGZyZNPpOAv5MwcFfe3ikwK766p2qhRCfgQ8zQsdln5Q
VOWE7Pv2x4u+Gcd53379XtckUkAzKooAh1hiyDbNevd6CD9WjPs2LnU+I6sKyeTF
KggPQ6JlmaNmNaFmBkDmPvEWJgXDFWZwqz+jwJ8JWxluzutaw9ygSrNGHq+M612T
0feCzyFZg+/X8XCZENyuwNN0mEpBSTmyL+lyuIEpOxgMy4B2+cv+NyHy2karq13Z
MaSVOMGfapqVhduNgwUvoNQMwjIokxmIe9iS0dpfl7PJcU0s0eoY6IqPWvHUet5u
LwzCPztrIm2ne19WN4mcvwbfiku4K5w9mOam3Gkc5jb0+hcpNEj1sCkRn2CYb6xb
`protect END_PROTECTED
