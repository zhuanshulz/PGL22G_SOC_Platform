`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CcQdHIdCKNOKLHrcO6lFUdEiXirgTez6TRK8840kvYas5ZooKjE6ZXdQoY5dz7x4
ZhSEn55wp1pMy5Omp0C732FOlWhJiTIv2fZ3h5wIVhBxUnociqQyAgxy7yt41r08
JKUebjlOVbtzgj/s03XYICbe9RPNWFviBTztSS9nowLWCFw+NEf/KXJ+BD78O4Y8
01RnVLL/Rm5LQGG+jHwMMRN0a4rcn2YH9ZRj1+BmjdKjrGEHya/2w9LSwi+IckL7
po4n573T4FfreIBxGz5WoZPwtQA1XHGyNPeu7QU1PGUlD2hjli0Dd7Xqu/MYa8zP
VMiSx6JbGEcvAbDxhzdZzR08PV1B34kvA4+oA+TKZw0HCkeiq7secUtSjINq3e0B
2jb/bpUjpokBklxz+C9bxsz4pX990cLzFdnC5LWqJA4/YPXazM7PB3+akQBnRNZ9
p10+4Nc7IrSyk+qtXSklmBYVFUJmfKuN84iUpcyDqAZNq10ShH5o8sSgG/7NysS1
2l5ZXdaUIqLyMKU+Q2VsOcwgQSpWN4TUwA520A/wVy0DX2wtjOCN6MsK6yQH/XPA
Kj03+b1PwiBwjgir9vGYUg==
`protect END_PROTECTED
