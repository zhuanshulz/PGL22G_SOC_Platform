`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rymcUq3UjSIEkdrg1cl1O3ZAu3oEOqSOeswhVPiTh1CXlbmlcTzVIVzBv8YJBHSx
a+noCtlHboQuod7b505Qr7RYP4piNByDxSe7E+EiC9GzJxQtXB1XVklpM6JWDB7O
v62OTVu8hvAtEby9AOj7CtSSWaFclayozqE+cPOQK1qELR1s0HMYIC5nNXVscgnb
nV9VrcL4TwaoWYBaWhjPGtAroRbJnc0tYt7pfArj2qdYN5yRySzLdYvWa+Xp6NS3
HKhhaYSYmFXxuPO7j1yCAUIpyy8CGLbvl7Ve+rS9Si/7WzMQL8++/4XqWpgDSoPO
zclcb1IFjy2c7NoPUvWO+H3qpZLo1Eu2HswrLgcC5OAGnIRvWEkEDznxlucHBx7P
9vcXcfC//Nzg1jitxQVvxr7ZchQ/vDnEm0bvNxq/4GqF0vPTBbWNIUYIqR0F7HCb
3/GyYDOW6S2nORmNNkH3CStK4y+0jfxqrOyE+GoCLXwzZLFM3+C7reHnvo+Pu37s
BSN0WJT9/Wfxm3GY+CEIhS9BHqjc9es363bol8oFtCq98g1KGL02QBcI4lFBG/vK
F4/8hKztm/hCZotB/uibKdnOxG0ZA9kibSrHeZV1h6DOq8KxhJiYklCqoBfxFOmp
4sSjCIN9ijd+/arGrNYMmEUYonmrdCPkQ4O+IhqkoXHdlaVDUTsNLj/KD1KwxjxM
Q7CBzHP5f9s0+Jq/834GsBKpTYWt5BJMjpa3H8Ilp90=
`protect END_PROTECTED
