`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yf2NvFZYtmZloQ8z6R7kLGr9XxEqDmUtZrO5Ak8V34rJooEyiet3dXjBO+rrVZOC
/8rsO+5nyQ11yTJmHiTf3IMi9wTBMc8GppGY2M36SVehla8tfYlww5HaDr7Z7ek/
IxLYW5UbuQjxsE18cUPeKHXfNYc1+BVODCxypaKNyM6Z9pYRiDUbnI12oU/qMcsi
Xry6ianyzmelnwP6U481Ir2FPOxw6NMa74EPCFxRltYBJroom/dFItPX3YmlAQ0P
8vw5wxrsUsAfgoLsKL+Il+fam9ykOUwLiBy2IX9ALb4SD3v3vl/+KJHj8HgfdNLU
NrmuJCFUgDyPTPTQ9Rnzxd0AKUVjXPsR+VJRyJ0ZmzZySr2MP6Ny15XuLouo2qh9
YKDxffWS/GDQx4KAM2mYlIR0hMaNUhqJZ+7vWW1tIce6dv270sR/zQbkPC8AhrXN
BmR6loGLaya7GwfU154n/ktALn568QirxWcojbLeTfknwty29RfDFTYcV2/gWouk
ajyxWwE3JqwpsF5QVxXo0oMUVFsUfa21U9fgD17KdtvF8M7YP1DyhMmN7zLmaMfX
0hpkiZLVIWR5bi12vaOPSMBH0rQqalAcul2OBjW7zN8cKTwmMozjIWlJXhRZqT6Y
qWLF0ZYFSPSvOQ+AvHGRyjRUk9aLWNGq/zqBYEc8h+22tm7VSMmYrnwqxIzTW8bi
iQ71pz75DhYL9FOZhx2fzUuJqAnlWDIO4eTHSo6p0NaGQFjczDt9fO6AsqGOx4dq
Abe03MSSx9YUD0dDl469qg==
`protect END_PROTECTED
