`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HF/x+P8PX7FAwJ+r/qlmRWEmRfpFIJvFF1X4J1+5HmoJRwl/ffySOmCdSTWTosNn
1VAtSgUsP272/+eSgsSLQmukndM5HEv+5LFKPF5uK5SZx1bJmx5CQTo5HCe811F9
MQej4KQqOkP1LcQ6BMNMHejpIvDe554GlJjtm175xt825kDGF41rPK4aLINPdPsz
jcCyi7nvW0kjcCzVsuWaUtedxQqeLZ3/SEE4IBwh/PhOYSlnNsg3Vb79PSqA5J6A
IUGZJXV/vtrQ9Wck7rwI8vOMC1MAyA3JUrPtVAUMg60BwWHSIZb8sm2pzRTnuPIV
MS2OoyCFv+7E0FKcno1+sokyAP6dLj5053bWXe129U0bP7LXaipVS1dXwll+Osq0
Z0XNqbl2iY7F6vRJyqz+95Sk6Zd6RpO3jLryLuM3EMkvvxg5OLEbCQpmgOHniDAi
JTYyWi1Icb/KNplY0/7ZhxhKCqQCqR9E2pBlit7bhZrBhIx1+Oo+sDFIFpgbp1u8
C0JX8aihiXhBsPKBZUcwB7tfqlr5/VnmbGqA02x4fdXJPGjLVaDxKi8H3h6yn3ln
PTjxApWdbRuRXKoWTDKFeCeSIajDXH1v8IdB+uBXl8wkxvUdCgh6rRy+rTFISzlV
Kmg8dXNiA8O5yIeY8bTBIjgSz5XLK5t2iUnvY5gpPYY8Gfwvo4z4mj3AWzEhXIBv
WM59hq/zUOOROe6IrEcdIp0qjM6mxOWgnj1RBFo8YEb2svIpJZRkV7Xzm3gcWPJ9
de0c2qHqhGOKk2oOs7Rf3UqcVdG3jqaLD2xWVKD6FEftuZjLbBowfCSh+IedcAX4
s+MnGi1v7xwWRD+fq6UpkQ00DvgfNK+AT3akfSOdwOjZnakRLkxb5LVDiz2IHPdt
MGItjMcb7G4I9fDDUVwcleF5sIs6YUBITUqDI99zmtMAK9jKSi4+mgWSdUy3xm5n
qAtAsjrV9mOPubvrVuXzUlJeNIXQ1uzwuekzUOgSK6QcGLU5HI2SnYdJJjyXviVE
jz1yRO42j9OKODsl/Mk+QGWGqLJDq3Nl7WByh76PiVH8nGiFYcfteMD8lF31UA2J
KnXyjOuCzRpHpZdlf3PYWHKEhFCbllyQlBCeJehPsTiOYZd2ZFDXyv6NtoaOJkSE
U5gnxdxLjaga1sc6C3JwmrQ43WGjMVJYucZNgSf6hRprfkr5wJsv7HJsRd+4ev1B
1qGwEGogxeO1TFRy3OzudrPGQn40dlogfJ+9xWbdCBNHbwq2zvWJkjxiGXdosg4m
d/99M3v+M0ZLpVmrIjjjo9mVl6juCxvty2uO+lNzX3XpcaHT+OW7Z8fgEoQbWdke
JYvylvkx1YC6QszQzMeLxhfUyTpygRdSxn2hnMgQRs6g3as/DYJ59sa17FezYGx5
jj1vrGrDBD2e9rSLvmC03wxnRMbqzdEVR3nw1SXAGPkt1Apo3NSnohBXsclIoEXP
ZUYm+imJ2NcDsMGpH1XbsHfr5mf2mp37IDwLDw1B+d5BnLRs9PnbiQLyHDZvlZq5
vOqRjzQjNMetxC2s2hi4mVAlWgjq+soN4CdmRpRSj+diS2bQ8wXKxYoyF9nWxH6l
6RhQHOFFdS8/H7du2JFc/QC2LRPUYeiwlbGVYmE1F9YWekiKHWBPfINkZTWOiW69
qLgjqDQhQzqH1xslxjJ31LGQWRwtrXaxVgmjjlvOCo7maoKKVgZTo+gg4JquN6Ti
Lj1g5vaRhmR+7X+m9Po+S7E2y8iodfYzG/krpFuNf6VTBLovHku0DfjOz0YdCk5r
dFtWaNTMlkk4FHQ77gGXoR8i9XwIZ/tP49sh9cWBlR+gElwbYP+ba43weCpav8Ud
d6uwOhBp3BMkugChV4oFIyk+i3q4qblytJi3s31RCo08UX2mNiLW0BUfGgLQLY7j
9U0oqUMK5RZTVwUvgBPJfk1SvYsQ6QXyyOVgMzpHhqXPoDmuqcG1bP6XUnPQRwaR
vdOjEPehiu6ZHMrTN9W1rXNJip0DDqa/QcOKX57m3t+aBnqZOBlDTWPeWYOul54m
DW6/J9emgxHHpwf+ziyIO313fZRyXBZW5teXVNCCmwM1Ki2EK44e2zLN/ieRexub
JpORhwwafdAFnmbt/pfxrFdVkLkDIkj5lIfJi49gaghNv33irHUJPmQReWd592ea
lm+YYnHgWjlaALsBhJBypjdJIj35iz+Z64tS0B4BXaaBHjkAZPqqosBaNZ3RF/1L
/TAChcHFxvfYby+8E1uyoCY5t+4Z6n3jKV9KtbFIghPuPN2euf0vKvh1Tf4snGNi
E2K7vReU371A8/4outF+Ucje3NaKwBIPqXY4K4di0OxlxrFZqajFaYstsAYH0v5R
y0o1QzAi/mbT20LNNiGoONnZlFJ9o6Z5Dm77hPESN+QPjWTOmc3a+mP+OmbfWhoG
4mHxpBoho/okRrzZuB9xGpdsoJGZJwspoWtQNFigFYtlBu3L+S8gY1TkHjZxfDyB
yieXjogzCngrjuCyJA77q4Nc8VZnnhHDUza3KYv47EOPN89R9CfRbGhppf8asc5h
0BMNp8sb955kp6/XdzupuKl/g3CbePESbYL7MTCixKma3OUd9ymyLsYu3hUsRGVV
rOKp2f0rW4kpcgo9HXMnIQeqmInn1ifg/4klDGowrZ0twTDvr16yeIFOOh5vsCKT
S1sVvyI+0MaAmsIEcGznGG7k9VKkGVAy9xURPfrV1lQ79xHBNyQcMDfJ9sLB6IMq
DvDmYi3cPHV4U1cEVYwjLXiboqFzc9eGtcgihRkGjE112WWrFaCCBJKm/0bzvjqP
z8uIRliH/H5J6Lb7u+AUFbgqwRsROxt4CivIp9nGLToGJtplsNOD/hqdyhFch4xo
MvpmFhsr6xVqM779koYx64wrfCwIdyHoHPgW9NozoMPVIcmllk7qhL8kyyvAbA9M
CPO7gU3m41jLdaPo4JTrn7uie6V9OkjlrBiHp1b2cQc97eA6iLYKFqlFGkgqLK4j
gpa1IyBEb7vMV7znqEZkviydzE5OAJwycz8gwGRTiYFu2jdIjGjFII0uZZ5ArHa+
HymreZCYxrhVWrCcXQMSoep2SqdRfxr26bVtda05yqXzOxkEjnH1a0bOqJ2PiOlz
VhX/tqBRQm4xpRlX1kURYtTkG6ZhnwgFvYA+pfum9UEZqbwcspuDAbgzd7/dO3wx
vNIq6hyS3Ie9Syy7I5yszlGzoySWE5BklrrorefFRghYYVQcGRZRjZmx2/DFf5Fx
+9ijJJvnWk7wu2KinMMNYvroqwsUTTlWgri6+uE7Vf3C1vlZlSf2k6rDqlUil4Tj
uwpwvvbSkmwSwGzUUej5YoUfsipx1xACqkQoxWV+9rrMsRvSsfKS3TNNCbHD4vzV
Vao4m2Z7SAbAiZh0US//m4zvDI6iqXSAu4g81Cpz4FMAvOD0ZufZMOunbQeyLkfU
9U+4cN5+67LgrwCssdyjKR+l1CGlA5fWQlcvaWoiXxJ2gwTcxQ52hDv+j4nAv2Cz
M6kYohort9wMKmUKbKCQpowqPL9I+hBteVHIpMou22rDClIHAOMBi4L2HDt0orMh
PHDgYB9QijDwEFsfNbYa+0+NDO29s026Swjrhn75L2vHYfWmaiB5oIqDqSBA3asp
Lffkw1booTnoJypUVQ+E/Db/d9AcooOTIH0v3CyayLj0LySulC8X2zRvLhR+KQH3
6kiOtRbRRLnmedet4/gvVA==
`protect END_PROTECTED
