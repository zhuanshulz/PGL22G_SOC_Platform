`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GglwzCB5uP+8Ktpx75+gwZpPL8a3BHd50XFRRHibOP2dQBCnS8bY/Y6lhhr3Em0r
OmVIFBhUBzG65L/c80Qof4SBp5IZ7gjLSpEmhJIB4Py5PRrqrA9yYXD7xS30fm5v
UfVGF3mTiXbcrQHtiL8W2pJT1Y4PswBwqTj4AYMLDMNTwr4Kpy04eH+Z3SmT9HwW
qwU8OdQqc/W5WIblbihIwF8EWArv+veadAQjTGmZoTMdghNUOhJ37fofSYIVuIsN
FKKoSE4Cp1wHJouAofAqBWehzM5PhQMH9pZU/qXzFKC6CT1suOjc4wo8B/oKymxp
x6mk981OD9A/bX7DC853vtNleamlyr3SOISSDGDmtR31K4ptw25TjoanSnFeRHQt
eO8egnZGNjm5qpQX+PuuFxD2nPqHGr/9/WqG7SO4qrlXXOfvvJmHGtNsr9WmI79t
8Vb1RtvZMRrIWS8KAdIpuXcP08PNX9f78OllQ3aBCsJ5kLmV9NcqyGWbmL9oAor8
C9HkRPg7vng/9a2r922d4UILBkuzEFg8EYBxe9gDztxADWeSERdnwqpYc/cDVToG
E1g0+67MmA3Y+N4roVcelXT9ll/J7U7MUS5y6/Mx9CCyrOEu5Rv6/zq78OyehBTK
ZH1gNPkKI/F7hhjEFQRQSQMjnr1jBgwEobzUkd+OsXi5EjCKK2GwikaEfpkBOex1
0ESU8y6Jf74kHqtnPANkc8rKoPeW+1V8QOuy2m75u4Cwx7UALt0legDWpM0AJnIU
TLoK9XTvAvVVbcvlrAQEtX/krPoKAuFuq4UbzPi4UPI=
`protect END_PROTECTED
