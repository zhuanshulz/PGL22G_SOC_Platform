`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7v5rELd8LwbP4c+RzkJICUlhhcie6r1corMdV9tEi5SFc1gcCDEma0zwlSlRK/92
C97WEBPvO1U7/MtzX2c0fQ+hIrhQAvw7uEy22uxnBf+vDU2g2ceCCBdrW5E3RaO1
G4CaN+8On/KhqjFlHmu0LTtXM73DHp/L6a09+vGewzm5H6t3/jKMgdQ08tju8XWu
Xcg5Bwb+VAwTLY/D6Rv3yGeHGGCcC9bwBhoisaP23tSk2PNFfFFNrcgmpGqX8hsW
ATJXW8eSlTEfJYX/NHsAx5Zw3L9siWfYoSblU+dj50g+5wTMdaH/ACyFtzm0xVta
smBaOwHu13dq8n5J8VlJwAtrihQyzkdtyl4g8zxuGbKU/rA8H/Hg6UG2uOUvLhzR
Bp65qzAqxd3p/jEbCr2sBVdqxs/XZFHfZS/HbaysjcYECGpgXbmrHEWbzOnhMtFr
x7UGcDy04Obbu8vV6XOT7WQGpGPfTPBClQH8OGHkpiTDddm6pXf6UnMLbrDYSXqz
PBfhl1MMSHvGVKCq29AaqSbrDjMHnILaG4W/qr/yoF3Bw0fzzIOToRN2Xyrl4gE1
D8EIorKtPWzTX/lJNUhaKjXPWx+TVG5G1B5h99t7gUaSSS7ja64ZF+5pZId0deX/
S0KAZ0Wj9Szgu4+y7476/bSxStjSkHfUdvMORiBaIxiEgdC3U4Qy6/siQMcbgYsV
ileBTATbqJNRx+OPJAUqhj5/FSLv5EknJJTdY6rK2xcdVOywFhTI5d1rZ/cxMiId
j2XXzy018GUHnjyZr3GtpOr5HsUtkT1abalgC7ICj5z811lzR2d5s90VRg+1EDFP
um/J5kQwuxxekT1gwlGN5AIOrmsO8j2Gb1W0AGonqBmOtUD1zVlCOTJip4Dj3kaB
loZCjBKa0fn6CmmACyqBOUuAilzQpuriaa55Z3AQOQFr0NFSBbcrmzH9R0np9pZq
mXTXJq8+0/Ahsliz1Obmis43qNIcW7+VolBvd20OH61QG+fyk3PwnhPSxbyOq8Wq
Orr5D5mQjqeKSL9qNv8FHdfgJdNePJXkeyhsPzO4abxRWRFUUiWOa7/b61TlarA5
kBfgFksEERhWx+1ckEz1EsC46YM1G5gJjadx0Nar+OqcTGtU1XsUT+RBbMZzVilA
WMNwQ+pUkhKid3as5PuP9VEnnILjQG/pyVBiadJ+dtunyJRIrnRg/2DnQ6+E7Vfc
+0WYjDiwJzuadpTIWPQCFssfdkDAvxehlP3fxJqabC8z05SDNPzxLqsD6ldzlS1m
qWYtAb5FnD7ZHs3Xles7OqP2GcOGf0Ig2MWiO9+OsgM=
`protect END_PROTECTED
