`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mKaMwL6Q881QQWn+FEcFVla7XHQ9xz2ReSRlJzJ+YtKhWJ628gbNApMPIAftWtLL
fTeVwSPkynB6M/4HTBgtaOcodHjIbgEqTQLh9/ZycvlLhmYMZhfbk3ymio/H/J/A
ZWnLkWi8UwK6ULXGoGautqeZzBzrzv1TgpQI3B+mVeuLhB2h8mY5qW903l7bwefD
qqMLk7OhMiMeEk55119r+oE2FVhvQUEmZPMs0aqlfCpIXvFp/T0WlOQGptP8Pqgx
/xzVOwFRUMhYBbOYkrdz5cU1eTWBqrP0VJkhY8nZDLvnAvRvdQirXI4nvYDa+55X
swLLPzlS2QYGea5GQHs40dGOjmhiiwIWe+NkUwDDlWtFltFPeNwwyO2V6doIiP82
p3/RrZ0ozRUuJqVGNL+SWrt6b66S1uGAwui4U3mk4grtNBN+4voeyGfifuvo8K8Z
TY053Ef3Auv+o5v6awxeuyu0IH3RCALiXrvNxwwA1AQ0MddgonG2eoXEkSMdDS4z
eJvS0Zkesxa3v7M7t9by1G8zS4Z5FuLYOk6+WzV1xCm1betGh9cln3OF+b/0qYYq
9E1Q/moUkehVDurR53lWCg==
`protect END_PROTECTED
