`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aZC/eSWGxAbPiC49OhAB8GcS7nMdUzlat8S6xQtbUhZwvoon+fQsHQkZr9ahw0Qc
0qFGBh5h2lN2tMTh5eItTEqOJZ+MwfDaRgMgvczvZOb/BuigXZwq39TibD/7MYiI
WMfmh4Gmp1mReLrZinSeQMN7GwvHK6/ZvOJ7F7Qc70WHwQMSGtMXHwdw5DhNz+YT
La7rlGlXg/m+sWb78TnnY6hJ7/boeaxLTbaSLlNnmag/K/jk7y79g0E8x+xRWEou
IChJXwvJCQYznwxWaK+BZBCqNlZZIJgNuY7HBNgvGYRj9Hrv7Bd5Vr7PAjDX3nui
jhO2nTR5YZPIvjK1lwPl4Aw6PuyYON+DqQS99dzhYvUrIdVDyRb+niX4YrYGlO9S
4IEs1Th0dcLJHF+fCcTL01IXxkHipFUUeI5bRv1J4M2qwlIKnkDvjpkkXPvELKFR
yBk7VSymkMDIX/BKiavjDKw6yaXfh02mT8lBS/xAjhQKZQn1vlYZBwhi+wDW569M
zx2nccP6vlv7fjpDeCEJnl6IMVNgzOxqfRlkJCu2BnNugrhjWE3mhjKSKrBGj/2B
`protect END_PROTECTED
