`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bnSNA6rgLtP6xfy0f6iXKzRmnmB57BaIxYr4IjlHf0SWy11qZu+28pLM7Ltycb9K
xlFEABas+Z6DKjSqKJi+XiXTfxL0Oa2/tK4nFUcBLpPrbn4FobtvoHkJMPFPPmTG
P/V6cNgNzieSmhamTMZb/sKfvMpn7WNgdA3KUKu4o7laJymcOc+k4XDhI6bC5CAJ
pShnCpFMGiIjNIPJX9fNIejwbRho+4g8Mwj5wFIuSmC9GVzhIAYOSPUNqH8jegCS
oFlhF+54OZCHAD4wwLO6Y9U3ZGw7hCqFQpvESHNa40FVNbsJTL5JjEVDwJz6xqaB
8jjZyf5f5o5NAJ66sidZdpAJDksg448ZpwW8t9wqoI96zhUAzwwbyx21z7srp81J
JHUfZA1fZXOozLVgixoCe7BCKjXnkRKXWf2ctHQEf8sXejVV0Bp75kgcD+PrB/WJ
hq6eLxLaYJOA+DqxFzOdqfqx7/W17PdQW7vVmwNlDJ40IwTst6jDXLhretRpMIvw
EyFZMz5l4C8Yeq5LwcaAuoRj82pVnwPTlggN9ZNij5NlembiG2h0dmxRuzQ8l8aM
zAjrri/hQM9aPFx7t3JhJxkAGsLctak+mmI2LG0kdno80ObgCEJLKXRp/bm94+k1
V3ZRiQS0ZEvRK50Q0aIhpTu/6fqHBStwfZmadmkuSK/hhGYEPyLmNSPEYFKCMQjl
ZqPaXA5lcqeyIbr6fNTahsPf+XT7uHy2kqeXpCChXyUXLc6WxgnGVD86gL2Je5GQ
hh0gWdhN0U6OCXQDJkkPaqwK/SdU2ozNpnR6csyZ6pFAzVSaL7rLg8JuiclOhOLN
DAk1ae41ty/Bw+MF/vPzt7n77vyrn2yx+lRGdB+mJV5I5cbLmW9HhQfl0DhNhg/I
8X5R9Nv3PmA5bQZBbnLqInCxav7680dnbE3aWwyZI9l40j5QnAfDsJRJZpzmPJOg
fJiwkByTgfWGfUj5vfGe+j92SdPDM41/LwaBDolWPih+Hy7RoHew0yk4fjQgHoq2
FYep5nPpXv1WsKhfUWLWa83qbk9IMlQ3YtQeCXHa28HoRw1VCh4Cua4qV9S6NERf
WaV+nqfqk53gNYhrY9IkJnffNDsfKDCTA9z+Uceed2tsJ+kWrEJB0+nwct39lz19
Bs4T8Jd0/3apSjJOLTdrS6zHLf9SOhidBfAN9WiwxBkpUwUEDe9zXnDmJUD5Akwm
yWSO82B2DFCTIxQ4DQNUiaN243boZFPPwNJI5NSIwQfIXb/7RPP20dSSHunvGk9b
1onalosdeUMyYt8sO4w1kO+2Pu7wfEyrnjA2OJeS0EmeqaZ2dfhaI2rqUoMTyYlt
Hva5JuJ2Lnn0kTWaO/FEjX+AgxisnhdOWPCf5AKJVY81EG2a7kZuPyyD5Nb4L2sM
tMEyVmqdMwlRqtUiiY35lrd91wvephka5Sw4MyJh3ug8HC4yjRGbIUcP9dmBQ2pP
PwRFs37xlezcrcobnAsyumByulucyzXy7xuiyTbh9MX8TWskYbfsT9eIOB0PGXfk
N8uo5bOteJ7Y2wfj2vKBf68jlAHvc/kmStMGuGsvO2OpNItr7fcZ/ExX1Ax7lh+C
sRUEUO56K24GWe349SrIAnKBz5tBWCaAal+G1h8yv7Rcw+P0zmM73GXRHGvtUR9F
CylMUCdRyaxhwFNHZX69nuA0tMd8mHw/BOfSycX2a36u9VggP7SrrRqfgWUr/7Qr
b7gQH+1253xu7mgyU5eE5xjG95XKcDTVo7unoeXJwSAPucsbi4EVw1ZkOcIMWRV5
6qsF1UYygX5CBMWAmcebNp/MtGjRRGT/iphrhpIKTKct2cDNHYx/Ht+XVJhtNq1R
L0LeHl0ceHnXGqE7Zp56JC0NQENIBP1TiYin9Qz+nMdbM0u3jx5r80PtQn6NDKbA
vKcVVoeSSOtx0KMujQq0qNzR/wrhLaKC7qJGpPn9Tch9QgYHqNGRfT3K2wkM9RfX
vrAzhWL/SeyfIq2oPPW5t7S5A35pm5ym2UMaMlxJH0U3oBKBQ88xNqEhYQyizpfP
AY3ZasYcgx3RCc8tyMV6tMjCTUYwW95PyZR1Z8pYG0FDAZQArailOGlwUmJ1pA/R
JcMX0BXx7sStwDYcshIYJ+k8GDd9kCGHP1XglpmH81wRhHeGCx3CxjcFObdn60vh
cDnMlSJ9/4ueKavmtABiuWhFq8oLRNaNaFz41eLxRK+uOCuzMZ8oawwJtLiYGxfT
W53XZSVZxl88xrGhODsBMpzyzjByFl0klCsPWRnjjzfRbq9v5G6mpJkqdVYL0K6g
RUyOlCDHeSO23JCemw8D3TYX3I9DWP08BLKiJmyuRdoeEAI6Rnq4vxOLhQWeerKc
qMmwvINQ57Up3pb6WNEc1px8tUBQXKGhQX+nh6IfeDhILBvafwz8NfDA8H4sOiTg
pMtsax2UFEAwsz1BJFrAs8/WlCsAMV2HV8aEuNFY90BSv/wNovAk/jmS4eHaoYle
otdcSAVkD/NYTKQGUAVgapC+glYJ9v94Ed0J0fOHwyV0LwL9XeykfY5RG/ex/SG8
efslX4OvU3OVULpyK2XPhJZNSoW/Yzo9Ulv5Mg62UNeksu3CVJRTscLi39o65gPY
rvT90R6m8+gkntDHc05syumMfLD6Ksb4GLLFGzAnChNi2bVZzrlGa12oOflgGXdd
V/k8j21E6xlFrt2EnAY1hI3KTZ7auBvodqCkqp5Z7+pWX7AP1pVrRwV+QqvWBqpy
Yn941/3LjJrfFqU3Ns/TGVx8JwipyAozl1BuIr/ZGKkUokiExXWyay1BSiPfzsZR
oFQ0iapgkpYFlKF4QU0EV9QeofHX9QIfSm8XuldK2Y4uVigmn4tt6TGYGAr0kn+g
Bn9KYI7PQRLnPx2rvIeeoLz1Abjv5KU5vISAJLJFQkFMf8T7Jos/gfRN/Xvqg9+F
Ffi6SZIyKOS5iBkhZSmeHTBFHv0+ew6AmyY/ab57trxro4cVrg+Ggi9Xxb1vQSaU
HAOL1fm9ZLDNtQB1OQyJVEEEmu9O7jXig1etMP17A91lAilvPyObLVTLxljeccpP
u6vghO9bX98Z3+9I4O/mOp21Fb2D6uCnmtLYSOBUX9eMzF5Tq9BDLUxvJ9j1DQf+
X8R+vQ5aEZVYWsivJGJWfSROeN8C85kp9RR6sNGgniPUbIeb37r023r30+09p6nk
46hgIQYCknwXpaglvdMFzEXFp7RY/vVXXp3VaI9vMsfch/wwaA3hYIn1uAcm8wyj
LVc2Pg6llRfPULtiWBSsMHEvBW0Utw0Rjhi+JBq9jgTp07jz2O669poG7aV4zLYB
hZxxYKTSj+yX3Mzs1v7Df/qYwOpz3g/SQrY5yA6kshfGK/LvYS4XTM8Jp5KKSvMX
s9+xsrVx9Z7cT1mMDU1Z/ZhBIXHRqFf0TGF9laU2DCGLZmsTlQY7rmn0FsvfMQbj
DdrZm5PGXKGBA/ilsACc6C9s+yrxOHIL9RZcGlSrrHT4ftu4cHLJenU7nel58Um2
4DTL5aP7Ue373qRJ2FquEYjKnsLGuN8LR9CP7bzpHubdrstluzB917vBkUAtqEMd
kbUIvNuG26GDzZWdlcpsNr+euGrcKMWpZ2ySKtqlZyopSC+p33rdis26NExlrED2
1HKIoBAGJ/VVQTePZN/s14ytWDWyWY6+DmhyVt16AvgK9xLEKFTau9Eh/w6e5TPJ
A2dQcr78lhjfsKGSf8pqNYp757RS4MtXKD3mn4n0zTn0wx3RDmMJURZk9MByRw4l
oyggKQadX/g01/9SYt1GJLl0J9Ls6Htdp1JUoGumsam6j7kTrc15wnZFEJQup4Gp
RsT4OKoBPdNdB24Dt4LenLEd2rRCV1YBS3SKHEnvJGzeXEoiaQuA6VH5lzB2Y10r
XDg48i244nGZK3nRVauGqel/iG5cFTZZ9+UtQIKf7o6+vDRAFy/Hl061Gig34n8d
Uh5qclLn5EnuUR/4MqJx3b2b4UFGX63g0dJMdTzzzY8PB7ttxs3f/yUBoQEIGw+A
1dGNQ/gFiX8BU5wbPuii7MW3hNMXSDRJlUZvfyN4GCK2evabnPCe9kHJWiQqSHyg
OyC4st2rHa56nzuR73ph/s1MGuAbSy4sHMibVLpTgbOK6dG4R82fZCQl5dd4wluz
Yw24qUNEgcg2aZet8laoC8lbwHN7k+4maUgr9k2ma3IaPNQmhLuCNpCgOQbfsdVZ
i5EFh35pucxe7UU/44VHRBxCEZQBesLDms6J+/eCorkHUD7p9Jg7fih1NVhnysts
fVTPiFw6XAKNYd/0XWwW7RyhepqeAAtZ8QtiW+RrcNCQzw37OwRKWlIDxF5HL2OQ
zueb0+j+28CbE2BSyEFXgZ1Gdt3W0LBTpKh8jORfXwt1bbhVDOW1iJCIh/xMo4YL
vK5c9mrWpnNYCNls0D8C/r7vFthmFfXcWVWuU+x8hIA/ZvG2JByYnNawT1rvfTvb
GsyRr63caDI7RInaY5X7iRT5ENDTsQ0EuhJRYG/8FtwbTMTefOoq7fPsKKNG+O+g
FtyMGxabQa+hpj0vw/g3ry+6Wh1ZkXcdX8fSMNu0t7+CJUUgHP/LzUVWUEwsu659
7DHfy/ISMqr5D/Uurf/sZY7gLGdGo2iGz/eXwIyeg+ibogaIwkDj6J8MqnUgKM+O
No/NsS4deuLfvNnTsDcLXB59FAvcy62qJWt6MExsvMBmKKBs3MWmA7f6VihHjtRD
31VZxX+Q6rWfpsmMpe2NAOhg3jCpJ6fYVEFp5DK8ZzpOTeANQea2x68Dm/6iGrvE
W0a1B2xxwj24b8iOXN2XQx1bCbL58esycTvdMDYvvpRMQea34u76vS2FHAhS4peZ
nIrXUZng499EygnCMT2+wXTXWyVrhLrrg08R80K+z/mUvHJuoJ8rVAtbI/glnxXh
W04Lbq6R/97p3VIpwWnRaNvXVfBgjm6Pn+3mbETXtr3MtwgNxbJ+dhYqF1CdITbv
/kDysUxzVMwANF5c5u7I/EnwR+tNxeKCzp1KjED0Ho2TZd5XGvAe7WYut0tiNbB9
/E0Tjjn43Vfl78ClbjzpwJaqVttJIMa5Ta4VITHw/Oz81pt4hbW5AFycJ278E8U5
8+q0075DEgb2AaRXHHUKxL61J4zVW2ELMhS2ZJzgYvszZm9sHHdhT2RTjo/XY/Y5
5YDYzIoQmBqaovlRIQqE4OBl78rVoxNUFClbmmsb+kJMDOVFnZ6/71xCZB1unUQV
+qYffuq0KJqyB+Rqg9Q4Ob2IFpGvRqdwNWz3lVhn0+XznBJkS2FIupjUl9Pu4dst
G0urq295lMXYlQzodL2EqPgvRUNP1y3WWFnMpdhmhEzlj/a6Zh2ukU2Xurgq1oV3
EiBCyUwpVXaXxfvss+1RhxlIlQlXbV9YdkOc7vgbNZaaK6+FVg6MWF6Q4993jZ2q
htyeRRI+oiQWdTiSCYY/8QV9aoywo6K8MWloCi+6XVUQu9p8FzhZg2dovBjkgxKu
9OHEy/JvA9GMBpHhKhQQ2Rp+nZdX9XZFcErfWsf2bk7AKZiQzfyHJPRK/yV1eSYk
bMdqNkr+wVw9eNarNDasoff6n97XCiLRztcGjBnMDwRfIhxwHwnTEuqdLc+LHWPM
+oPXuUpIwKW+cFfl5pSlghVjlEh5QCTlOBDEurwxZpr9uPuqm1YLJh4k5zGEqJuE
Vk/vacMeJhS6NaPdFIMvzPYinvbrzn/vKsqgeYg3jUMG6YEjhDpDBjRE7YWeBxwN
U4C/8TH5fGZ04Jygcrcs45RBls3jI9MNajtRy4lqKBj/0z2TXfPQfQ9iP9hi83yf
a5AyosAPANzfk5DQkP+OneFdmQv9lcaZ0pTBJ0JrBc629KFMYPjmyQQ3rV/Njquj
MgeSDOZFE/8CfuMlP9+/cAJPYfVdMwnIfCFfwWUIVPiBP1Bg2/AI+mGdbFUZ0RzU
Q/Dr7y6ii7niaTq83DXHSWr8G0UiPxvm1bA2uYCdnxLCiurHUGT37hEG7RUJjq7Y
67SLj3mMvS3PM0ZrTgvms0FZlmcruHqcCh4RkHr2ye72yBG4UzzVl5OsCctTt3TP
7xcU2MauEsQodrEDrm3u8gzl9uOuG8TfyApN8faI3qbijMwEcp1+hJLIbmU07qJI
EbcyVSTTBhiTAsDCUv8TgpqxcJhO+XbBOVMWx8IxQ4NgbJUaHO5ccUReZX6aGcX8
BibNe2+y0Zh4XXN2NM6daGrTiVEZnOGYIvngDFpq5+9UyDQaVMtiXcFA5Dn86eC/
7his88+k5oszI2HyAJF5G+DARnXs7n4aP0hkZjgTX/0/clyUhoL0/ahcYpUaTLyg
VrFgHebvzngFvjP/CN6qCa6bYzlskpptW2gR3e9UBR8MAtVZMLRYBboo/jKU+9n6
G0+JAwVeRokPV6vQNXZRoDTzONe0+tYEifmj8O9k2i7c+SdpwSjhYPvDt40COkPR
lW0TzGg/ACL3vlsmPLYVhgMc29ujQmr0FCbn6eCdRogT5sr9tNnjWWQMf9eNeHFa
+xxD34UprN6z1/H1H4jVXtf2yxeKRGtXdzMCysm0l2qhCx0VfZbbq8hFOWixUOYm
`protect END_PROTECTED
