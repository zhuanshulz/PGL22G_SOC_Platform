`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QolTsB4P8k0RiCVwCVza8erz0uWU9mdcgLup9f+wVEhnEwRynqEITB4FrNm5Kym3
KcujjXlSTC2DG5NGvbvJ5Er4JIO7+LP+h/gvpGY2nrLSpUDTsMvEV9bSW4uqd0XA
cel2zKvoQ67dJAjTjlq3BsmLJSnG+s8kfA6TGYf89oTCJjCiDPNI1ncpiJoSp3HX
k688qc8bzwxX2+HL763HAnKDPAlF0tMPWTym7y9MFYitJnBQxs8ZK1OFfHKbjORO
pGzY+uXb5jrSjmMvqfljRgRzOwztDGfJAfiyYBW+j3PPKqOUMSDNkq/45DJqBhii
u2MrC3hNBtuKYWF9P/72EInSblRPIyi6AaQR/QtQLoW7o6MV3ix+472Vt/zDMtJj
2sNMFT+9a4HAddpT8maB8CPeBcb3bXTWcIR856qE28cWc/geguUp+eRNxMWLtOjl
eFM7D3yDcYnQwA6j0EKN8KwLYFhnhgs3Blh6XQ43x1y/LbyiH2yDSFOWhKZkldTL
49knnT3F+jTZkjpDkCrZ6xjFKHXxe9zpYGcjMWESxzCdHz6KGrFGuHDwOpKzPtBv
kDn7+4cACUlvmc7qoD8X8V50RQBheyXZmzFSnSIZQxc=
`protect END_PROTECTED
