`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PovfNKg6VPqeNLBJ81uW+CPB2nOtBrN3zyIh99hhvZVys8vqMDCjCAD3Iw4yZDfQ
nFfhc99cLOgXiU0ihpsOkziVo/R9DmGIVATOLm4KkTmvZjcvDk+SJdOCMlDWRVw4
N0M3WoFziGyeGK1qVPgqYOMT1/XGqrz3D9LyXRUQ50lsPtrx+F4LUK0bVjIoO1yP
L+kzlavxUaZ8PnouP9avidBFHvlFPesJy43rIcyTV+9u13bVObeM9E+zFk9hDafw
TSQ39QQmgvREiizgAwMYM+UABpUzuB7iOIR5yzlVU6G9KSj7bo8iSfFGdNLaHt8U
UpZ2T0buRx31gXta6oYgBGoZ5mdDorkVECV0bAjwHxF0Aw6W+nVyhV7WZmGGPC2N
USDNpXNv80nAqgl7hz+adK6z2zGY/wfecDeyAaeplS4FvvXKPc+0bhjY0GqzfOh5
mkOL6j7Hsq4NFqr/JBFw3vQxXUlbAQ2MyHVpHwed8mnO9231CWs0WXvAH758eZCF
OrFf1H9HZU0z1QgFeQs/moM8TVMdgdf5JNmD09l/sJ+aUTT0jJl8bPf4i1rcXYIb
jVHrUNa+X9GGtwRRjy9adz9eCsghDDUguGnpP86ilOxLcM9qWmpOrwNshVFw+LUb
OeydFi4F2jMFKrByvERVPtC0Yhtx2LZX0l8hAaXit2AaOaltMPGhvReYjVB4Dek2
i06zfmcq5tHQUo2AnEgsK14ZTl+NiwciWo0JIvTBf/1Phl1vCs/vm/9uipiYxUci
FzcvTKzsbVW7V1qsfnXwC/gQ73kM87PqZjfhWzprI/fJASwxVu8O8CmNHVY2VnEf
ooQAvJNyLqhiQ6Ho7+FvZWK1WUlsEiRZC8W4BHsfsrFTTQuAWLKEB2pMI9TVaLGH
czM34R+PFeUrK9mTy6gL67fuBEAugyw6t5pEgZBnclvbIoLwzb4CjMnBLhTNgH61
z1GE6LFH7sO1dOXtiGx2QaLljMbT2aQnzg77bnRAD6VfEfJzC//bqHRKtNI6y7Bq
hMZqFpTxB2bTAgnT2YIr1Zj55kC7WzKT7tzGJEcKllsjgFobicAjgmGcscWKtBnK
5+wSQjukFKhAiAQKbXn7XiK80cO+LXCDSamE85CE1l3VM1vg9ThYmsSV+HnaGDn+
UWuIRfdCyrl6d74wDyf1X6x9C7vwsqZMTDFr5UvAJ12JQX6eu48a/EpB/FxwoR1B
/7ZFD9w/M3e8STgxdowqRmyz3dYaN3tBbnokBjs/M7LVjHsZaPlIDmw/y8bZkY5f
JX2f7arB1VwVTRtPqT3arE2jhHdKEVIXWAAGHZZkcdnafZJ44X0iUF1UIWTr7Sb+
m6zWYEhcRXE4yFhmE3LOhgrkTmmGe10Uzy8IgVq0yvttq3uRk254ENjsIE0ybaag
NobC8EuHj+2QGicgGmYPOgS1jm8LZCWGG0bhca/TXu3kzODvlWw2doC7RhLl3cKM
5HO7F5yh6qbpRN+dQOMO/0kvBxpdlAL9wHJ3duvkx47WLPh9/TZc/q6r8CakUmE3
ik1XUptkXs3foFUSQLHsFlyFB52Wznxmmv/ymtU4bDgbJp/CXPk8wreZFnfiSo0T
fPEIsXQePBngcT720pvsnKymrTUoWPVe9SUASUYDY/nLmQRlgPvoZR6eu3ZZWDqU
+OxJmOwALBu5KyvVriz/IAc+unL7ILY+wPuUAb7aVDIPeYzaTWszLNmCYlnUepy+
HB/UCe58DXKQ94hrZj/99ocBFzKkkDMIdYFoWJplC72Ksb9aTz/FKocIQUefxOFq
MEJUzeciCKsV/mk0lY+2JZqBwN11veFBK6sFn0dENUIvU4qKpF8qIFGG/Kb+ujt/
mqXTlAHXbUaEk3d/cxVkuvZIG6q1ZUBPeT4AX5vzfcjRzu1kMzYoQm2yGArcSNy7
v1jZqf3bvGhtgDY9P5AbSGGrkQAm1NEMNN9xTGqAMflfJ813cYti8Ef/3vo26kxC
qpVYRXh7pSdSYMb9fnCIgIn7ZpRjSoOIW7ksvd+2fscTw9ng0a+0nQOXY3EDc7t2
6jw/Mxqwo7SUctMFZRd5fJYIymgX7hrH3uiXEYxuwJgN2lyEMFDpb16p0AyFEdla
5WAyaxN2u+pBa1s1ON/VRnbyyLxbrdjO6Py4xPwIaI+Shto+ZIPcI7a2Rcdur5f7
AAUZvVkQ4r2zxE+Df+1xUs9vu0cuhQ/EHlwRcKmqR4NGRJG8F0Q8Q+m57nHk9UFe
IzEtTzSMEs4U1QBGrNp+LXH5ZrxlvzHTJ5Y8bBaXU6RuTCZZGeclzbGJDoU78JQy
7xHDaNhIwwVgvWR3hdRpiuQQ7HZEW7OhmxrgS/Q7g+ZfyUsAiT1uPhdImAHfwlSM
2CzB7Mh9CmqFc78hD3NqT9rl9W+7JG6uczubTt7PYn5mOO/4jbZZbAok5dnLfU0O
JKPsjm3A/a+fRet5RnQR6yCfmreRmSJKiTJFpyFeR/cNtJdfo8qTKySjy5E28DU9
ywswx53Z1G+Xt90OO4h2uEQugByv9wetxmXqRR5pLPeXbT1JNmRqaiv/4OWMQZN7
eHLusarJmAV258tQfrS/Ksp8m3HLxNXC+CNCDWtCyS/XgF4jot1erODEv0uNK9Ag
GnhO+XMY+S680GJ9uIYp1I9Q7xyyp4t4JaoMcTKz3+X7A2dhVu+YGKybWwKppxXu
W6z5AGGZ92wwDpKPSYSp7PU8Dvvj0MeoLqpoPi2MZeDA2wMTnSkQGZ1O2V906QCH
bcM77zk2uf8iMf7ZcvjB5FFKsbc9pSvIzbmP0wybiKO0p8vN+PEGM1/mrspwTr+y
K4jH3vxPWu6nqEoOXACgDg==
`protect END_PROTECTED
