`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5PwxLcQKUPZrfEXmO2PJeNyTdqamm7VWsfPFDqbYOLLrauqFjDhkpe68kwJpFOUk
wlaZyIEtaSnx7W/b1smBUHaBdfCyG4BaolBPfQzBtSoya+Hwdp1IWMR5Cy844Tdx
30fzTac9pAH3X5rXZSGnp8e0FHvTBEDenHAell5CqkPc3s8IsFsmAJ2jO4mMnboI
VHlMpeevdX5NcVprlG1PmTUOFuljzjM/c+d3hrr5AJeHg41SpFsgtyN8ZiuzcrLs
2lKVSw6nteMdEdwnCVpLoMTIiTaKyQk1vLpzhOpjuXIYGOE3rf6vgneZ+9KtW/iY
DByd4gvKnuFS6TGCWoICZD55XBLH6YyD1NprbKPZVgcDIGUwvWnZOo3LBt2eUwBg
RV/+nBiirjpfAm4jdE61ZOxw2nu345Kh4ad++C4s1kV5YQU4KdqXqXhusNXTe5qC
QO089Ze181XMXDvkqzYkYtcgk5bd0nzugTLPLyImzvnmy+m08W+gXys1fP/on41B
A+EPAuX8Syt3yfjAIHjFfF00z+SGDd1NqhBQSzBwXTdcuoBotcVWB0rjd7iu1AhL
g+trT/un3k8vdo1os8+zR/dkptyduoR9sPtWPHBNm4UVl6K5uySNVtJ6nwnKYlWL
i5AEaeuaEAduzJ8pEgeH7ayDScr3EPEnE2kdf4UqzdQLwFMNO3EVYoqUaNi3wQTz
dQf9imPx2kWwUsRck+YyxKRLdSj9QXb8KgOFG0BkfsAPYTR/QyuRKq37wJTIh0P9
GOnhsc1dMEQouc0gaMvrxNQX7qQAVBWPprtOHsifjLFvJlDFCoQB5K3TY7vGv4ed
GVqX5JEEe99zqt0GR3DJqgs0wIUG78YPzj5qbzd0+aXfdRFWQc+DCF8x0UvIIR1E
sJDGQYNrGtev3O8XLEUCSjE6xy/uuEGBRsCyin9lMkRrVEVeOz76Bievp7VtGnpm
XFmm6SJycujm6VW3GM2mYeJQCtER8tfJFFJovW5oHMyyBKM8ENJ1+RDtw9IyhZjk
NYtmuAYOBplLguC7eJpl6aFYQDNtnGfuezoLuxHIOo39vgcmwgqnvkiUBUL9YEiT
SO6ps2RJ0r/L+bbiYi2z7xWcRiqUSK7K7h0XHyEGK/j7IYHLISAUZ/CfrGyVc07Q
sGaP9ICu6Gv2IUjm2lZ8jOCERz2Xh02BiKJVubMXdyfI61D+pB9V56puigZM3urN
7BJCDAqylc5BrPJck+UlpXBrmalSaUf7mYsBAJkRDjOAWAyjzypVkk13GKepoMGl
EppkV9QQxJrfKcdeOhsVwY97i3NjcEe5R8TPRzTF09b+wuyVUP8tYIa3+rXkS7Fk
h89aRq0PaVBtzNilmjRmXTLynCVae5+jKHt56c2Yeb8/KBlHsZh13H4PGmqr8/17
E2M4isz+pey2OPRvYW3DZM6h5g9g7u3zIVE4zy66y7sUlItLFUaKmPvl/1dARiad
hizlSgBqpeOeg8umH4DcmoSBiKKgCAZcMTXwohO8K5R7XUt7ngWCSrwKmBQ5dGnm
14k44QgmVrwikjywzfbAP/hNZ0PjzeE0ljDVsm5O297oLamGSNjFZqVdzySPZnR7
3K9kxFYejVj77k66uv+1OtjL3Q1wMSb5nRRYBplrYDd1PZQxniEoWk9j2vZ+20VU
UKr/D0JHqEJdxPBFDVKE7pwYhxLDbwv4s9BTXy/l8Y9Rn/agauBNuGxsuAJd99Zm
+vqRZh65r5nkYPgv5pe8fX3wUAh9E1SfhbQzdQ1wykgj2W4WPOtP6z0+/eJZg6bk
EAlUnr5BOi3/Jv7uGc1kkLC6AsCw6SZnNPWbyEtOx8BqR1Pr8gdohgGfEfkubf6c
B3jBE5e0+QTD1KsaTnxTcoAAkTf/8FiA+4kiIIiXLwEUN/5D+JA3o7tvFBPb3ikI
ljtIXXiza3hMkvHuvUgXKb5GsN5/alNhj9G7JhmHeFRbDwubRZ7M5iZ2/59mtxsI
UqMd4CljOC9M/BZmo+x/mmlY5cG/fxltBhhyk1QYMbhO2I9w7RSCSCeTxXI7u0ka
mCGSthrfMSunozwdrZ8FcCtvFfQwwrWduWbkWL0dgMxkQ8ZjtyPU83Y4R0oAEca7
QwwRak2SJAXvK+YXDmx70cWv8Ps7p1WsbCBHa1O6lNCZlQ7FsOGXbtwjeTblw0AK
ZY0VqPuzMNNxmhuD68hgdDl24CsjJG+qnmsRMQYdp9F4LAP/MRBExDhzCIReyx8e
VHrx/FidPkWtZzRUaYgiQVCPZGObPo94xiAuFhknPSq4B8wdywlXRlHUqdjVBi0P
GI0GujjUSx2smMmasyakc355SaborX/mbErUmOgZQYMmVkjryMhRL90yPSrAKKce
pCT89rm4mrPvbFsm0e5KeqmjiZyv7SfjqEHjhNjOfLyuCXOWnOq1Zf2lZfGLIxB/
VqocvQWd8OeSwGjBKCqbdqY+7x3gKoahXwUOYh7U/cTFz8Th16eC4jeqwsASQu8i
UbrtjumpAMTh0ELhf+46X9D5l1dNWAc4RUgSj1IAd1iEwePrD2J08BSYJgqyhfhv
coBbjlYIILOIZtuBIXOSr6xNeRN8AP+DlvKp5cqqMUv4TelnTYYCbUo2VBsy+byA
x09AXAJNLnb+Zke3chs45ZQGTfb0BLMz82qXO6XfuDATuCsH2H4IlKh5uver5C/E
T2jdxRHtnW5xvqVEnciWzz6QzfmTuC1X3MV8KC8nq8VG5syhE+UiDMV9BPrHdNZD
JCyFklkQNurlUEZNFPMSOSyYRMZM009ABtdJM+S7UI0sxul99QALpx8NlzEiFY0O
i1zJX5jKwCyhdMOVgyC3VXo29OXshzpI0jmL9pZuQhNMWkMBCKnijt4ld94em+7/
MoiojOauQXreN3prXl0MTZnq4jE8K01j3dTlBCNy1XskWP9wIS9x3rzGG646vCMB
zXMQE/lURR9Akrnk0hebRg9NGjimJ94OepcQXm4dRQ4W1HjBt7O163fwMFlBe5K3
ATNuNatj4kxrABLuwfzIQRvn3//Vd/aINlDn1+HtEngN3wDOTZqe1yHrsdqEKBGA
RGhrT8Q2rCzMGstGFyXnF8c/7/etD6MInVYYNBOkXNnr1E+OpeeqbAfOYYZMUzMA
bcAb1twdwDHxfJAML1uts271vOZwUxJfHpLM0bzUX9s7OnO73yD5axqk+L3yLY5z
7ZOgSLNyjW1zhnPfV3zhI/YvHNMoZi1KTpAYI76h6F6EgfemxGdL9uGV2FRN2LLU
y5fHlp7SCCWx7UhjcEe5XwncZzP8LdBKyAOTC0KrExjWvJ6ja7hS3DMhahe3PXNt
JO3ZLNQuhjCocPlZMhx69f41Le1ek4UE7Max1xwU0RVDvRjSX8lCqQtVk2ComlVP
wMtJr71X4rz8WKuxO6I62E+QXC+gO1uqprfVlGUxwcVqkzuoY49ydWG5uRLB+joC
lzslcfRJsyedztVe92Jfs0XvZUmixTn/NtcUPW5e0AOy2gL+xam88S9XgNs89pUd
TSDPtIud+/Fv4M8L++Bm+5jf0Ndpic4+XC2IyiBkTqr5grEPMojlJCVmaBAkBeqR
NQv4VuagBESxmvsIUKyJQCJsxNMAiCjXXdPAucJPASWGZeP3f0ruiBQZDvs0KUBw
BDUEkqFBSQFY+DAA3mqpV/jrA7pg+1Yj+JSHqUjWH50tK/nFlK6V4+M/MdjHxVTB
IZt+9sJ1r3JrGnbTrT4EqWVGZLe/7oveyG8whLUsS0jtHbP5TQ+g3w5/NOSWqbjj
qCvJlpLTVzOli/UTd/QxzhuUkP8a+0qIZPn3AL6/jC42dOkfdmzBYPuJqTGR2hUv
LFNcGqIVB8AQMH7peVz8mnk0dSsTlGwQJx+Mf0S6uetoXNJjEbsw1739RC/m5h9R
QxJQPkz8mg+Deyij/BKWcFBR9F7vJudwgVFLjWBmZfcjSxrWYzpJmNi7TnibjlBG
QMPwyVq19FKO2D7O1t7tYVDlPR3ackJEuuMp+wiwXw2ABMTphkgexYjUAUKQSV4Z
d2MqDg5JYcLrTY2yTPgw6OAiX60wLz2xkoEz6lXlumcW9X1qVhmK+WdhHusL3ShM
f0DbeNE6GbBS9xKZ1mo43+zMOOCuU5nP+GpKGp7xC1vbURMpCEcY9FJxPHhg/oBO
7STJ52ysSocnq2udgvPUe1F26hwAvJNo8eCs7YpOOjnx79Z5mHYLH08W7s6GYmOY
mqhzZj5vIbmpaU/Af6XJdBwXZvsHGOLqCTCDO5UIKaGDJc32YgswuTdXJvuEc9CO
lz3jP9hjFFeYZW6LuqKf9Zl2lbFe8kwXvnuqJVgMEccD1OWKF+UYuoQROVQ1rA4N
t79LR7LCZxssnC9DqXAjtGVvluCf3SJe2GpV75+7RBxC3/HG2wwsQzEUc/IPfFKU
sWVFPP9l6ZyrnprdWi6DMn5ksTRGzFQOLffg1Pl/jIzCkhfMhRnzjZldyIG7Sj4W
Cargy+if6/lnBemPCeM9MSOkvHmbI5ZLOjoA0XxhOqGiaNT4ic/j3ouBGXXJtQzF
T8EjF/tgXp5PwOndejqvssiFcpummk3eX8QRcdyGpPmjfpxsxDaLPdJgMXrvOlBz
z/Q46mYIko5VBUJiOgcXMuht6qCWT6wdNpO24imMTMv3QMpTi2s+aXCArhUvZCnQ
ZIYRhxPXC6aWEhyy8e1kNPOUKxIh42KZlo4EhxVyba1H36tvVgiHK9ueSRZswkpG
BQOdVXdMHhz5z+vZyGpgyckgaRd+kVsnaBaZ/pDFFtW9mHkDQeu2BCBRsoxNMkCv
KMwAfIiUezqfqkcCvTykUUKYjnmF/3fh/Q39UpERFfEV4tPEqyeobaCSzUlqTs2i
CzWRXMswgA3sk+mPEBrEDVcAm/df061hFUo17uPlUElDKPKsdsUBYnQ84Z3dkYrQ
6+pCBSjdQIofTziV/FxgW1dyxyinowFIJEe0lJ3Pk+jezBu3+8F0F3BdYRevMJ/O
oYftZ7aMJ8q8qzV2sfxRlXdSFpVYDV181R5AjA4zX01b3wji/GFdMVJ07UK0MwHo
+0tan9vokDkKwvEpt4Ap4U8z7bE7fPmnBH0s8OwccFHxISLOtgJfeGVzYq7Av4FH
j/eKvnMCxsJ4vlC5qbBZO3cfK8+tL2BHGePCozo36GmnpzK7Svjd4WmMinxqirz5
9OkvLlVJzfmrhY2P3sVo5wLOzJuesM74jmxIUQmkXB2BCrGLT/7lVNYBvhALWiHu
v75RyNP1tsb4HFvgovR46D3hcPZbcWJjVE0S3/A7NfO0zvyA/Yoazlz/rn/CXipu
j4NogK1ROW58UkaBJ5UJ24edOmxCpwb9L0C2le5pS4d1qAmvOkoLaZ4cdoaCNRO+
SOajrr4Jwq0rNXSzHpJ1BTW3CwsdWr/UhY+uaGqOfBQLVflYJPVuhMWj8s8Zfsv/
pGDKrB6DZL+ChQRklRv65AyATQTqccVuaQlPBKpmQ2xkoqsfgLQJp7M3I/6X7yAu
fnXJdc86YlJqDrHP6yTwbtJwA02Z4X7+Dgs7rNPjK9Pzmdg2+ZPjYv+htKejVWt9
E+xnly3kfpJq7PsXFStyjd9awxIplzTQ44H8kkc4Nnefolq9s1oc0K/8SEjutuAn
d24aQmNp/OS2Wu17R1z5GUzV0j2I+4GwoxTh0e0xgzf9CRyAYPLgHEdzIJOGkQTA
b03wz2PVw7Yi2KgZAr4z484D6OlPxresFGJaTUpYpgKsFfPAeaKeE3zd2XV8FGTC
fSmaEutGEJEf9Qc8M6471vttnqA2TWW8z8oDNZi6+b83dw1dI5D7+NMiDqneiS6q
E2DOu5NWUmWS1bk4s1p5VxgFdOqa+8J88hephnvMb1x2ZWl8Ud8Je55c+yf6z+5Q
VcAnEQocWJ553iDvMUwB4rR5ZugrSSNylPh8m6cX+2+uMNPa5c2SLZPElc8PuwuS
hMqBmFBhMSBiA9S9bidTQ05eZplgNA1v1zVnhCXLmLNOeQERYHGZLlfkamZoGHkp
IHYfO0NMOg3MXlAuurme7qE9e0xUWUNn2MLAqoTXYghEI4kekjW88j7RO5uHa0Lp
VGJhQ7E3Rf3+tDmCPU4Zur1g7ZOB/2lXifdu+nYPqEH+ak4VlvXZLN5jzOnBPeIq
tbr8PCCXWm5cdNMzwocLGo+6FAQys/OCD8FXN62YAeqMEzqImIim64/gd9eTGHS8
xTDstJFz/hwADOn5ng8+chXXL97N6i7NrTFzfyg2Kk9G7WKEJOVQHkqGIN0E5rsc
Wm8nwn4Yenb2FuWUrPr6Z3PA6g3w5dHCRLcoXsD7fY7suoO1hV/xtSx4Xq5d1PGj
a6Sg1vHVMADnAA9L0Ktl3ggrY2Y5b+Qq2pYC8JXZCoyZVgOfx+LB5qoLvvVGztk/
Wz0ePeB2EXgrvW8r3MUSpuXq61eDk+s15MXsRcgLgfIcarzOtDzzCeTTD4xYA7mg
vYLS/j64K20ajzcomhJtxAaWFupfc02ToLJYI369z7qgVT0FGg5GSyV14tVmGqjg
5xxQN3t9ZgSBpPl/TFsCnklhqFBj7USERBMWadKekOvbdtNrYyfmp43cyc1yfl97
yjhO4pXI/2kEBJsXIqZQV9ZwXcjBNyV3BDKVGD9E2hmRtg7g7jQBIbHDk4enio1P
WN2fyjMk/ujLY3CQa0W3gDEuQR0MlEkpGtFOzoO/8Clougfy6WSGz0WW4zsXABh5
Amwfn2PLfMjY76xnveI+Qkk0Tx/ln6okMAK7J5tShroonQr4GDOBDXq2QzjrEBsz
tOvwWGbJYJmHAXjjTj/g3JdWYV5a6r9aZ11MlHezLyotpH6FKtUoQl7VeXwRkcfh
et5BAqfTWJs2DH87rLLTk1WHqpRrdDJxNja//m4pFZD3/aA16I2xgNjXlp4A6cwd
Ew5Lh2K9UFBGeLvvKE+/bM+6OvnUhRw/Y6Xg/KmnJCCu0s3VlGUuY9gHK1ZrXJwM
kwFiRTxmrW7C8UrwdZBaqrQFTdmNUMU5jWAkoNX8DDRyViFE162V6JMN+VWE/JcJ
X2JOXas+iWzy7z0GlWeWjZJZ1yjMVGVJTpSU8l75rTK3z+FyIhXEnRXkoYI+66Zd
GLGRktQbSNAkfsmCVa1rA78W9QnTCRV9k2EQ74EZB8kpTM2nSuZeCQWAvc5yrwEg
8IfvaoFSJaj9l527A3loACxH80DpL7Vgc4+GYI6mNHlAWytfmHgdAtOPjpagAON0
fA23erTMv0evhMeCTeg0X7MnD4K94zW/eZz54TP1J1TqS2OfvpunlPHksGCZk+LO
rdN06Y+KXjLh9TBBZRLesiBbpTKjWlWLM0jT9Y4ym38F82eiWpA3nKtGF+podtYD
na2VzIiDdkIr5Pb9ZRFhTe5+zQ8gO70cl2VeMKZCR25a/3IML3BlFH4NaP4XI3IP
f9P30BDxxVxdFrT4Jxc5KtTY4n/ZAL9PPdWffg7vKJF1tAhOIbuOY0mHINXYNPYw
KU/KC82HRkuv+Ut54bd6ZH/Lt9v4HbqObFhduyaZZ6Xh5XIUMetvvPtW0X1LMuNT
JXZbzHwdsBDRnUDE0sCYHTwF+u6ZI5EkS+DMgY544bxp1b9MryWIUc4H+pm+oeUI
aoXU9nO1o96gaBXYURMPJM1XOPq1QGBA+2OnsHhR3oK08iGq7/DmwzJSLPxT75sy
HwjT24Z7g1rdP0I+RfShbQR8atm5OmTMNGtU/qOgRGSrWfRhjp5yZEMl/UPwWf++
jV0AzQVlhbaFTQMB772oGoDZkXWW15CLfc/ZhGleMq0vsbAdppC6LnbWhBS8U2de
HOf6JNL2AWRF9fffZKLCEjFKLJ0QasCjTL7wEjhhrM61lNtxOYTDmkcXT+q3m71O
f1l1SH5wBxR7dWj4XPSzrl5W/pLvOJYaE4Idrt04MeFpVkipKG4+AXaOOmn/TsFl
6UhChdcu03MV3dZVlmnEWCCi6Y1iUdcqRe1SHTAJKkKo9O7DxpjsNJw4bWMBW6k0
sFnbU4/sgA/7CaGlOA1lHYES4IjRWqmo/wOiSmdhLKfqL+/Sr4uw33NCW0DN013j
Yy4bD0u1Bv7N1ysJ+DejcPeJkrPpwyzt8iiB2EKrcBdZmRV35kVW/3Kk5bExIcSi
EP0XCd4cyd5WA1jq3c4o5cbG7pFLWallN16GpROIi6QbL4jBMbDpDXezQIhhwxHj
+zkJcI0PPgxYy5Q+scgel2p6rQSfcJEh4tvS3qu79ZR5ehhSMM1Yt2o0tHrVUbDd
VaGZNkwZiQFwEiNwTIZxswVGtAkwTrpngWKn8FJvhak+ob0eGnn+KVOImkKO45YO
fsLtw1rd6MEbc5OiblRyeq1oCWNX1m0mmslnVy91yxdKDuojW4taK1+D0vy6mNeV
mkbP0I+ubGp5ZUZwqLFY2AXLcOl+GU0oRErNcFhltUTiNFzeeYPKwxrLfGNfDRlp
PWk2zvndscsPJalzB3wv873UfiaZp4q2ecZRTyJEWWFRUil3CGp2WvxGuR1+12X1
+y/tdZ+B78j2kyDhJNZ1+TPqff4p3BnVFTTGTEiGZwHqEvgE0Zx2PxfKDyF/tuOp
wZCICojPNlykPKfas1KXQ/2OJRrofZr1dGYVrAoMsC8GtaoT+SNtUw3vOAVkn0JF
`protect END_PROTECTED
