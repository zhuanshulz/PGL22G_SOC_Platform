`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s71JliBC2Ym4opwCVu8AR4UFEc8/+s9SbHA7ZdHHFf09lfjVWtXXWJBZyXHCI5GK
2hysaQuqoa4RNjufxEoqIBg5HYGSb+Lvgzjht626tr3lPnyZWCTNUb9v1MHWYmzA
lMPt7N5/+KMIoNij1nqCMd1C5Mufo0Z4DBEINxEQuqIZGkSFTtgQTfbQNwUswbrd
WQxrtyiSOgKoUlmkpzcCnYWy8wH7eUi3PzV071OsbFGcHE1XhywOMPRm0bKKJ1Xp
5p99RzCb7U/hnz8KeYlUEFhAhioGp3IHMK3RGcGNTo42CXUs3WD0JjAinHTcYV2v
6YTywwVjQzLFy18VfDavyp2IWP43/jIqy2NVLA26fuByP9Z4/WNp9Sx/ANro7H1P
MJA7k40Qf3Hg6EfQTCWp0HBq55AgGkiThqN8HuzHdkoo03cjIxRU06utz2AnTbaz
tDXxbUz5RbbnZcy3wzNMUgU9ReN9wNVmnzsOcNHUNzoq/AWbNeTOL7q13jyl2dgY
p+4HdlUTSGAI9reXgYoSi6TyuXb5c57fuQI4C8ypnhCnSRqBVxfBe3+kTLvyt1Z8
tq2tFqakwYHAqQccrPwb4j6QWSMqd51NkHwmsRhg5//Vd/Apgoh8xEG59IGLKcpC
ddY8gk1Zr1cm5KzwjhG3806ngwWGRDBX3ZUv2/YJ2Y5acjMh+TQ2LJ3bIuv8rhfV
CVUyAIiP2RIRsdeR5jGADFECzCfFm1TQB3GgnO8MIP7WpQWxDpnElb1boSpXVerX
+6UcBcERyMd40VJeDzlwb6Vv9+lUdOkiRdsnCuzwORymfHgk3wRBFJQVPjdwIXi1
Mv8q/TKSI6yOexRLlsnCnZiHR36yuYuHbDVWLfh55IeqbQmGnd1tXfft5T94WTsP
rbZonJR2aPnymMcwZ4WJXS1b3s/p+OdSqtSl1xddtGL0OHopPtbv01ZrcIJ0hMce
6IYgmQBv5cHRQFWce/LN7ClT9d4TjWLxXIDLLmlF9HikqdOrnL7BnaOTIq9tIxuB
vBNP5NDVlmUVYGBml1LeylFQtvkla27MAGgue2uCiVVZu1p499tuhhwrx/1c8uRd
L3wZ5sW7qOIbOchTXqcbkuaeo5lChfCFwGf97Xhi8+ni18gi3+xLK6OwA8/CX+M9
3KsF8BDQarFbXu1wRJc1iwNut0J3eDviCzRTympoYTajOveGHSCdSFEo4AFxKy+i
4wCwsHCT65uETpc8eQLaRWV5wAnCEL27g0hBbNZ4KVCWCvjeuBhykaMleH0ipJaK
1Yj/aRhC+FGWBb+abz9T5pj+JR9/CQEXcxmm/ECvL/QNU/3qH10sxqVAO1FHKV6R
SrdSlrJIUUBz3KZHS2wMpl60DpQzLIBc2pnuHmvEuXK38vM5hL+ivv2WI2WeEcl1
yvFxMog9j9Zb2gRSMJCJkk13a4lnSsTQtv0z7Pcg4PDBZzKdgKW/biEE8X271z3m
mMYDgD/3AtXO2Q73zcKChsc6UdsFnUlCMDKKTjpA8O0lRU9DWNMCuN7nNe+nSZ9Z
KsMCDjfogxIa4dmS7u5PqYSLH1avJG2Dc6RBz8ORMCdv7HMptt2C8gwCnOwecxZ/
9E2DW/w4JeF3ImYDLiBpjNaQYz6W/RDxbyPYk5Kp132OUGFbW/PPNrhfL/+qNGEn
DTLYXgSIrv6FvHhPm5DleNniGwRHVd4bOxedt2giBHRHnqGyJZnIXeOxQjKt5eUK
MktRVhIRdq7N2nmdAoqtSd72XkNX77JlnkCsWgsfcuuPfND83c/QpR5MjjjsUevv
iGhRYFuI8AnnNRaUrcxUvUEN1wj3kyk0r8qgv323zv4vASnBNLLFFYhIe4qQqRb3
u22Qx2awuC1SnKK+huXm+pDcsBgbifnD6kxS4TmXamlJwbry7PG9OtYasX4j+B61
DETtnAZVhN+b9AXGh0bIWgaGhc+7FV+NReIJpHJWckQFxxGvfjsi39NdMAAIFQTJ
OvrrxUb1e60z7ZtT1jyWtrV4FIarObxkFsyxHmMPagpU4LWWc3fA5/tkCjFBLOcX
chm44tW0kfx++fwaPdRLqrWkx2bc7aS8M9a1XGL5Sz+lOJ8TKYHu2Dy1vdojSpws
nzdXQR9ohe+uNhI3fpWX91+HSkfKy250dTkOxbnwdiaoRxHbvr91q9a5y8qFP2WD
O4LFNmoqWEctAhZOaD/aeyM39G1STjaNe+2DOozUXqvYKFGkDCNOXkTfiDbA4PHc
3YFRbIq7TDI0c2Mbaid7Klt9viy6x2Qb9d/+SA2z8uz2YE4k6Xy/hB3UQPTGNqNv
A0PCbY5AacCD38P3tP6/PA21BlJKx5uBTH/6Jql+J88Vy9qKavLwRE1eHU2nhefG
Lfjw1UNx6hHqeQ/QelC+NkQ49ZpxEEV7VAiWgRYZuvthhfzQmTaLssc6TXWz5fPw
s6T5q1Df8M5u+j2CAlySsU1NTGilaBvUfP+HsVLfm+TLUJOm0Ym1aeXekXo48GFc
AaCSDIVtHf14uzxhawV7bpnPPhjPeFaImYwM4jQX/POvo0SuWvELnhVMlblSb8EF
o1Yi5MIYZx8mdirOUl4YYAytimMwGs4u0vf1HELuPvxYPm+9KZKAGGmmN5bLKxOt
paHXApJBPQMesIrvIYYJEM3zSyxHdFPpPUwu+ePoQOuaTuBsLkpxnfNjZ0qQpNK9
gJLRL5r1+SW/N9AZpFgSnQeLtbuh7v+p7JmIfvcJUBDRqm+VeVFJOzEeyDlmD+7D
5u2t+KFtl7NPCqRueRjeJdSoIYzAOpkBGsrejkPdeSfiAAbJ/5ETd68/6lZSWjbi
8erHm2GAGZ6R5KnWysdvP1k49F739ekx29gHC3tSAzwopL1c9Y93ZieGadY8uZwP
5XcuQiDpNchh96YJH+QMVifXVxB+LcDuneonQsF6yeZy5d0QVTHAVcrPntxMNWj7
2NPahkbUrqnc4cf62w2n9uuJ6U53vdO9yYBh45YGdU7m2uujvRtGy2tNDK5Il2dW
A5+l/4dx4uLMR2j72di/hEy3Nzip1l8RpLldXxUsqPuN1B33pZOyNG7bBlSJovlY
fsb+KM72oUI4CH6+PqIg2vnHGaDnGqFxi931YEUtqWhs4gbSbsQbdNKn+ni4yeu+
VVFh5vOkAJPRC6jZFuNe/llcgVZE9ycAlxlyEfSni14xwSPUBFAKKsT0h8cS7pao
Wso2QdZzYCTIoqzSdKf2McMDv6u8kw/BrOW3yVrogwzT9Su+t3VxZZWJ71YBLiqR
hHXeu2goCj2RUf3yw6osdaJ6cVf9YVMwN5qk/H0FLrLLXQm/oi6qXGQuezlmienp
bPlzO71OSgMv3+n721D6K6QZB1mUI4slG3KPVNtk4rRLUEvqmDENojb+7wHfF+58
h9NfR39clV5uPIg2BwB+K6cos33f43kNuE2RGmLeVxMb5ToEPVBXVkBmRg5256oO
OfNN0HNtOjvNGkBVSfg+2rnZ9KMmDKiFtKQAa65N3BTJVg5nhr1HbvQVdkaF++V0
xMB12ii/fJkP+HtLIQAzLzH639I4OwdK4JG0SlG2STgIZaB7rsQhqiCTEM2mZbTY
oNrnS/VlDqZbWbK8MV8x+96GU5x3Jl5rDlTf2fwjpdUShtg/Fex4G7M8Yit4Duo2
lcCE9okYSb/vyC05JasyXw9y15ogS3AwzCMWtSEHzEYnQ6st3FPwvw8LPbt7kn3J
dVQIjOgIToV7W8UtRbJ/xG8w2RMRQ+YHI6GeWuWi6DvykQKLdxJ6N9Fof8B/UHK7
E467yglj4hAqn0+8RDsgMz6G2pLATt6BtCqs/TnX8ezYu9uDdNKoCBaGrR63TQOR
TewWEg7LTC2RvmS2FlPeFFbpn/JDLRcTn9j3comtN5c=
`protect END_PROTECTED
