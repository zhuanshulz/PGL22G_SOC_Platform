`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ga0KCNUFS3besLRRMiEvUqBdQZ4udwLM0af7L18Zpmq48CbDau1HQfS663rsEe4+
mEmmghgY/a65V00MZUPsIAft/LWuxmT/kINlWCx1VdFB2ZnLfxjtpWsBiKSol3le
XGH6YHxymmmQHMeuC80mZzM1g5Xh/OUdLsR2eTfKJ3cS4Nl3AeCI6ZI9k2itQNrw
HmhUIIhzXJDfgxJbs53/KrqRo2386pTBxCMQPJohHdJjoE2UWdvB9R7tnbhE0+vn
yLNn/9zKZiyBDwyXImXqA+EAzVPoA6nJ62Y48HNsPsdqYkhdIGQ8G5UNnbSAKGZ7
kQeUsLTU78g0MW/bHSfZ7F8P7RdCcmXnpfv8yX85668tvTd0Mqffud15JznqWOLI
z2aiY2/5ECcdICfZ2xzRuW4c3/WWAGqIWDv1Z332q+R+sp4z9SN4fmJaVNo7YW+E
08sNNWaylSSUNEIMU1IFRkzWCe/uaV1ABgpwfJwCMnODE9KMDR0UM+R6GPslKRd9
bYo7hzq/vluL5W3/MkebvQ8rcex6Rqi6vmRb4ItA2S9B+VvtJzmORk8alQigIqwQ
FCt/ur4BLCJgGFxYIQwDa7J2m1lxSm4OaLxQpIDCh+Kgqt9yAbHQQvnfC3rrPezf
9r0JEU7wpzn0WpsAJCars5KxVE/dbfomX4Lj8Ra6e6c7ROUkVUDjVPuU5sXtZ0G0
7fVmeqpX1HeykZiB6O5LKyGuPii4itb9vIkW9ZPSAdauWvfL8uZqx1elRoD5mntr
0JnSnbaxOMKm+g03L3YrQ9dZUD9ucDc+2kUmYeUkCHSUsWaNmqrLR0YMpc6RYvrR
+J/YP8BO3z49AvhvNY+WdNUUWFlQhKaCWuSGGmyOzEMXLzeIxe9VXmgjFLyGhxcE
MVcSn1mffmiBmuAJ8p486EuuiGtle9wYgkKizFTr+MbQrKbT9Ex25PJLONG9Hf/R
HGaDaJ4v+7NC9R/Xnd/fTfbayEnkfLqXojGXIQICwg5pE0VHT0ynBPEkArdsPFjJ
EkvdGerAp4AoTbi0vXhRhpOi/Y0t9ywkbgebpk/x75b7gEAWAM+dHdvMPGvUz+p0
y+AoX0+Hp3Tl9/CBlPjsxg0/UY/ND/t0Zt/XTPQahI8m4vmNlP/pEKnXiSxvex8n
Dktx6yiRNUy0EwpN5zwqeIKaP4qae1mOG7/Pu23OM0FpFpoNZiY0Eqg/wIep8rgl
YNhoVDy9GgWuVKHa/u3oYlHudp+QRKMQgWuPkamf/a4pj4TmBwfhDSfbgJ/Gy62g
DQngSnnXPYdYQcbpbmZZmhLO4RCdHjxuoQMTA9o0B6nMkwmg8XoYb7HEL3wX5P+r
uHFDUeGTChFLJzmOcSqxngi2j5F9yUNBYKlhFucwGnYqoPe+ojwNbEj/gqIfTLyX
f6YbRePicGEUPgt3LSQ3b84l0W9dihGrs5sm1mfxR4vj4Z5KxjZ/fZRiJ8Zsp8Tw
nG7lqUGri0nRh8aElAxKGU2V2TXLuJWrUEUBIopAgTkD4UpWtYtY3rMzAM4xCfro
+tzVYwcYFFHTl2lJsjxE71yjKf9O9WhOQCbNx4P2VgSAmPdTTt9Crlw8S3iJXX/v
RtHqbItz7dO4kpofi9V10VLv2riBsbCY8jVGcDkI6GIWaU6fy5LgNah7GvoTJsJa
ElkA7M6YDV6mRj71LJ/J9rcNCJMjD1BE3oYWDDhBYmshQLmAiZWcCaiWxa0HMke5
2UpHobZxYslMTpLVD0qqa+m3PwbhJtaBBoR5q50XQUnwBci6HD1uodU6XVY5hMGl
G2VcH8uZ2mm9KRPk/WIy2xRIpEzKKtMRpMItYs0jhqa6Hq+EFLEGjyVyGmlbqWWc
Xvhq9SjUa8ffzgf7oJkclKt6oiZuOgC4Bo6bksZ0iLPs1cZYzIsjBTCyhNXps3TY
7RaMK/gGlHw280dvELQe/MJ4NgYdn/ANAe+aYJdpACouLQJFYPqUeBPmvG9lKLwy
rLSIelGwp7SB7nB0LfWPO6EdPUSvhtf4sGWyktlHIi7nU1Yi537SKawRip55N0FF
hMBMrWdjqFuxxAYzla8aE3PrKs5e8mgszuNUcXQsHNAovJYy0owRAhm0oNUMzFCG
n6hq/rWC6xCyx1/uSzP83mZJ2O6i3Lu9lajZZay6BnCTV6z+RldtSBHYQWsHtznK
jzbvN7Sc+nh0BV/eH/bB697eJTfYlysMyFMGUxBadh/v7tGq9NQmIJNbspBdtuCJ
iMOwHmuswfEEuDx5TpPeNRg2I5Eh8+EYZWXr1kCKd0NS++LixV6V57xuRVkFXA6Z
`protect END_PROTECTED
