`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zyzy6I3eiTjeRZ733//kwfkBmv/k2hRLIFk9hCMbZYQDmQMiLNdA9Ujvq2Nq6Zh7
MqGejzw3ZZXqbSNBI9zw14Nr+4o3mhVW0TMtTrPKoq4mG5L8HuSfmdlMlIVC/Avm
RFt/P92+xFBALxl6G5vJEeJNAngc+991EMZNUiXGgx05pkqSCWzpR9HIhGnRxMQi
ZzvpVIb7IJ5JAJ0XBMP544YDPjkG35xTU+kZ62Y0jYI3ejFviedDTrnqHWHfHdrt
KC/+/M2/1fIoGH4136OMB6FfasfXY9DqhntBO92GQ4RhwzjVu7F5qpnfZW7BLCfZ
4eO270wzxp3kbguLZrNkXO9emcDBOWhMES52g/bdqd3MeihobD3RjPYBdLGkr78M
yWp3x05pCQGk789JDp8KTfgltKhBUCtcArgGZAy0GUO0H4HERvWZH6ILI0gw44n+
oOxE7Bo6y9s+Y4Yo6YeM0ALXQ9wM4nGN3dKWEyNJzgATumwiFVOsLnMtUeuzXt2n
eNIWd0Xt05wHNc0Ney2Df6oWBP9ACBv7bFyr77BoTm3SseUlKutwZdmiWacZAzC9
haZR7Av+CK3G12PLA6lWv+GwAv+xYQ/mi/FGcuRHmbtg1Xacx49MK4iGE0he662X
8FuOQ25fNNOrMdu9lPN2ib2te9uEPm5gefNm4BRjuSuvXjnwmi9orWXkN4eub3qK
5Du3l/1Zl+7ICoD8efROPxXPKFrPv6tuvnUZbvPbYm4UGxivhZTxaV79VrVT/7w3
Kd8nw02HQ6YvJZBvwsrBoUrcZw72+vrMhQediQzLmjJKeSOfod40Qp4ImDdfBP2i
Hb8ikxzaTY6tM+RovafPpctCY+6iXNPo4DyONdm+hfjvhwTulBtVTjtlHaJ0xr0e
kwZuiH1PT3d8uLKTwpnpV5T74Yied+UYsP8I7c7ZZxjMAp9ZBGCBrdY4eC+8EigW
NSmNFcPy8cyhgQ5/U0gfjTkliwVAIhzKl/8xwc/EUho/iCVsheaqnDXMQERsF7+6
6k8pdcPiTW9u1nr7OpsIk+QH/pHezdzrZxXT3U872GS5CilJLibytTracQ7J8h/M
/haProE1FMAXJRA2MvP2Enk1lu1Cq2Ylw8ZKZK6aRogswyjoAG4fIk3wJmkIbB8Z
1rZP5fHeeeQRikbBpgMeGg==
`protect END_PROTECTED
