`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lDlsjiFvWlqPZW353GuH2k6nee8FSk123zwUcWLE5bhbK4bqumbO8WuaXncI/RU3
CbBXJF56gBAZnYZ5eEF8ozmzeMXaYCNspqzIxcT7/JIkpnRqh79EifiY+RG1gmC/
omqyLXAWqL0rQ92V6BwTD0E1Cgg+BVqQv220a9UgtWBzRUqp6VC30w3WibMJJArZ
MrPMyoW7yRjieuuLYMJwbL1Vx8zENBmcNCMrWZGsPItWE1my19f9UU1evM+hWPKy
c5ayrBMMi+d9qWXtQ+QUG/wP0KE/49iCzeNb/whW+LPTU++DQbEtJltcBiU0ruaW
v5gnw/+OpvQnGwwRdW2+kJNKQcceWkMECGiNo/dpSSl/01UU7hh+mIBc/OsmmOKJ
PyETExS1gRQqI56l/Fjn7yPn7NQEXjI8Ac8JnQElALIVnbEo1xh4pDoCRt1gcFPT
72W4yjoVtPxRM4ZpejL4IbKjo10OpWqIsT28dn2zsiwuZGpVF3F5lDTMtoDXa8BN
aNefKpvyRzVKzEglQ44p1Uw9LfIVl4JVw4I/rcgR0srH8c8OGuWJZCzwYIbb3zka
fLf+jCtdRRS/i6KjMjWV35XeMOGHdotq+xZa49Xpcnc+3KDmuv0J51WxiBOKAk8C
ujRhGwUlmxb/Vxk8RnwvxgwaypIy1SCW6yEb+3625xyjyJpPkuwHpOODbJ/xEhDJ
kL3lcUnQptEYrzTmM5Io4rNcz99DCY8xgXDOrwlZqVA=
`protect END_PROTECTED
