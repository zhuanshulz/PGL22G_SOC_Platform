`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
569joKQrqd4Eyzit1dPw3TkwCKXsISiMbbxzvLuuviNjflnKQGBFj1EjP7xLe+Eb
OcQ9W3sk+pfBmaHQMPpmHYD9P3OGl2q5W2wj8xg8I0qtnLRkNVFgg41rtJ54SAfR
3f3MzSi0A0ZXgQcR1V+8GRLzu76KdjJAaaWzRAAKxHO1Ij/eQSw//7ttW0GSGFrw
o63q6wI016NyF4ob9GQuqay/PJcF3/0A13JLPaoXCJZx0oShXX5JRQZfAqqJQHjY
FDjBeJgQ2t8LbpLfgN4uMLuGWoEL1kNqCe3RbtDaOKqsBwxOiDOaqNU/mJ/pwsbl
Ab3F72hXs4NxeCJ57sWUdgFaBohFeJsdthx22FFnaFNH66mU/6yQZML/OIJrzkhi
ZueNYXXVlQ4vQ1j/5zUUhg==
`protect END_PROTECTED
