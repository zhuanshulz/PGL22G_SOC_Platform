`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qnv9tXxQpsiORctM4CL9I5mSkkjjQ63t/lbqM+TzCwYvLltxDuIVfg2rC4gQoFAd
YEker/Bo2TsRx0QItkzWoB0+wVVIVSTyr+GGldOpLx7TftYc16tH5s9Zx+D0FGcD
f0/aKGhzGy+isY6neuGvzMkCgE6BBhpdlZD//x9ii1juQW2yh2kSA0Ua6leDvv8D
bS0v9lEi5WseUt64IbatNFA45ASyrPNMbI1W5uVea/gjAhJzjoNLju4gBo7Tge3K
RXgRcJzyWuIE+E+6Yg4SaUs/gQ9RHZR2iLDZXpjkeMPX5S9UPdly4vho5JpgUlur
jZkuU/ySQ8k0yHoe9tiTh+MUZj/NralUNrLhOS5iCTPQCiL7+S+WP3ZOVLOXOgFr
vXv+cLZanL1OmbsBE2HhfK14OA0A7Whmwc1neA4p6kwC7tupd8KqLxc86q85qJ5U
wHvihyAD8cY36GAFpd1zEP15FhGM148Cv6F569beY3ifedhHpQrEorj7eHAI4IUU
96hTybIA63y6QMhW+3WDhaFhIrTEkAm03ZqZoXFEaUlg/B0m2vVzYYSnUuHq1q0K
QP8TEXh/gtgCqZ/pyZSPsWgKIl/FxlnqybQDDKyHN4WTel8QEIMWjVS1ui141rCk
gKhHUhIQf2CcelALrI95qcqcU5zCdowyIwDxRr8p5q5KfnPxZGo7wE2DTA40PfhI
BWyKLEkSC6dlEa1DohQIXiSGN2B1Z3nzbWaC2oHZhGOIa2sdd1Lm/kbg4tzg5cqB
H9QolDiI7veMQC9ukahl+K1iXSLOlnQP0LDUQmTteDdZS9BH6HO20u+A1RTqO68Q
FKQLhNd51VW71IYEJjOJTXBmFt4imhdf+G4pVP2tAajHZ7rVEvOU7AphedvkeZ9j
s5I1E1SfywCTb+2KICPBbRXMJOv0tTDjzlHE4aY4BIpmrE8W7eTyqN31qShTRTgb
Zf2pGLxqh8wUvOez9HeFS7Zy6IQB95qcr/VEk7Tik/5ft9/oKi7Nkcbi0bMFJGVw
MQkb5JGffFlkN2ahBjarCTPww3t14g0H4HHTIloCp/EPsVpHM6B8JagWtOOWkRqO
aGgEBdWjcMPVCMI6biy4ekKGJq4JODqorT/VbG5erjhTeVzH5bq4YlDqPxCziQu4
c94b3VvPD02tK2h3hIvXhyewqiLU9j4Zu02hYjUpqACT+KtaJOoBYhPEvCv1kyBF
ka4gshbHpAFgn57PGi0zkJ215NJQrgXmpiNXf7apWbdSW8j011Lp3JoFsHJI25dp
V+pyRkO6z6Hefm1ovYv8Kj70bKnfeg/oJp3AShh7c1yRvyRp0S89YBA15ouKh3vy
IFhNRWfmlhpgwg2CXIoTyg88Qe95u0cmKeOBzYU6039fghHQDZdQXvgH18TygvFc
6lsUDe2ZQa6ja2tIPIbbUFcMc7YocHkiBmOGFEIY/hC4gBXWZTMH0AvT54OVZ/WC
UCabIl77l9M6G2GO4uKp/U6/9CLNaELknwh87x98u1pGNwr+m2Tmu2af+vhe1dOv
fN+LpSqTjmFF2DtKCw/GQlpqwAZ/8GSEGeHQXDIxTYvbTnJLdIafOKz857QYGxe5
6RcmbRdqbvYVFs7w3+VPBfbi+tQ3WGLMzoygva0jOATxIYGSqA22duUJLZ8x45bn
Aw99+ejBWGcTq56Drb9BboKrj3E8FS7zajz4sNebO99Qbycv7s6oLKjr8Ch0Olbs
z5Aa7dWumxzoAIuMulETXmIx31mtNkf/WIj6wqjx06Yz7APi4zm3QX55CUIICpu7
MTSdqJLX1j68/kXlUW0SUMlIPdviVNTbtIijz20a3aVSU/pUXcj9bGPWB9T2ryEh
koIbb3o3zvfnm4IZ03FuVBwI3qiwtqin9S0Bm7yaReyQug8PzzVU+QZn23lCr3LJ
LJScU6ZBG5/YkyrNnZw335YCU3xsxpSuecgVI/afHF/g+B0OX2TsWqmhjiMqnLg9
Vnr+/GiRgUqyLD+G7w3lZOkb3+RMsj4a0Xw+FXVaqEfUl64R8Hfmd63EfGfEo6oy
5yiHRMfcZXk7reJTIEtkjEFOI1OBMmTGZLwT1Wo9l6vLY7Uab9NftMaEJKhEePRc
79Z+lc95fZWijZ4gH5xys97E65bONzafqgl4o+AtRFQbK9cq4ssCzBAOAumreu8i
sLc8kJfIAP1PFIoSddMDQY64lKdzuEo2ayrJ6e9bmb+FDgKIl6wdZhEUxFkSIOak
PJLl2oINvX6zxLm6RFinFRnLuEqe0sLxL7pgD4BX1o4QkuZBcbjLxHC3gzd2sLtj
hg7ym1VwcSj0iDLJ0Kf/bBjNtdykX0dMpXg15RBq9W1QLZlOEELPsXLnUj/DlfgR
BALuVM5uCn6RKboBfqotWL1W8T/XSAOEVjsOUAREXNEnKMUJDEii4G0ya+Ogm1Ed
1Iuv8Hs2E9oJF1UW6Mlf2anT1h6ydcrnUCKFgiWSpposhUKC6EgXB6iM7IN557+9
rEal+lQUgxiQSitQOkWEZGURK4IQcUG5JvsUchERqYFqVfrZQN0v9h+Izt7AfNxZ
0AnpZkD9Y5wPO2B4lyyfAzrAykCq81TOZ0QC+Cnf8KzwksTW+sNus3z+uIy00re8
7qWBMw9CqhgTt6c66JUUbpU50ZuL1G+iN7tlHEufagSLLr11m9x6wnUuWuvevQP8
rksSEkml/6EMfl/lWXZ6oxzIRy3jrewk8GQ0Xn0RACf8MuSNGD9db+pwebo6wx0q
YhQdoSPlDxtNFZlCw8UD3SkB4gVSz1Xc6mZT+fyXvzGo7duzs9B0Hh/X6LfEj/Eu
VogyTgpEx+A2yecCNcSGHZowZnBTK0BD3MHMKoAXSWpPUy6hJNkPD2ixSZ2b0sSj
VN2Isa8lhr7VtlOHeb4sDSkKdNfFza0G7mAiMFUPZFlRYnim68FLRk3RsiuL7f4p
WX3KjiRwMiZrwwGXPBI6jt/dc1QmtfMtAuX8YgNGFuJc/fPR2R4nT499O0DBHJCP
iYe33y1t/cCEMFISXoyjxdBzR9Qiu55Ssm0uCMRll3I4BYGVdGIGsekVDnMOKKR/
P85LmAZ52gU2G9toPfJ/meyI9hVKs6Pi3CApx3WlmuxsKsrDHoiBn8QaRR7xxO70
aqaHk5s9XL9iz6tylNK19I5HGbdJXL4y7I5iEpRZsPdnJPvnNTCnt/8YRtL816Se
bfB0H4XnWm05GMbTbSHBWiRH/N9GbnsmRhcNpYGIPGH0X10PiG4Laq54Ak4FVuvn
8GyTBdo+rKmeY+EKnZHWF899Tdm+CI5WfKP4FzyEZzpfWVyMpsRokEJqSMjSr9Rr
iAXav5GvS4q14jrsTt+1w+cbWZhi5wkw8p2WSN5Q7cFtj7FwyN+e2yRrF75OHVNH
niIaQm3JDwLshJuFHIWcQw7SBdTJ6sHMRAvdD8N/FcGjq6hkzGNPzKVJFDFnwf6K
OkJlkrcI71x1NBdIyk3AqsQQp/NUSSUhWIN4lsBc/e0g6/Rq9/Kl5pWgYH7lNFFH
tJ4vJ2eG+IlIxr7OWzO2ak0MSLopgN+do7TxjZL9vZKyoeLicFQK3oEQXcw9xcG6
jH5FwfC8v4V3EcFdPKTJo9bfbNgUW5omXcFBiPQiqItgzmJWVX1t8LEfw4BYE1LK
tfWlGWpFYyvvDyQTUE5Gg4U+l5a9v3np0pjP23NcNb1vDpmhdGfI4ti9pzwI+aMr
`protect END_PROTECTED
