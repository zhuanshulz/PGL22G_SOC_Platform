`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
daU8fUK7aIL9W55ROSV5C4o6AyVTjR9YYMrNM3C1MUDEcBgjov+49/+o0HNyRIzz
lFwpOgxVOajBWce7edMsRBEA5BvJMiQ/hx+VvtIdivv4Kr1A0fQecHK5ix76cRgY
nUHwdsLyuKZQYDVOEl4eabws9IaD+h4dTI17pJXPyFFL2jI5uDkaMrS2tsZnDHS/
Elc5iYEWMsoRKDOWW14M0O1xzvsflLx0fkoqh8xOmYlEBktqsCQsfqXyqNLFFU+o
xbVqZRKylwzYe+3dfaeUFcxiQ5oik9JGA7cPRk54LgjpFgasUcC9v6jN96vphjZv
f1GQERZ6RUru2R/LXCzIeBJIgoVD5UxGLEYsygxaDC22oqsPevmsvXHBcq1eB1gA
lW61USzZpGgeUY79i7C9O4mUgb6FTMDlfLTshQi+iXXr2tKPPFf6RjvpSAGHcEt5
yXJUGe1zNApVoyWjRnXPR11wNpWy8BlMgKwb7koxFeESBTMdFZZ2MC7Yvsn0TTuC
IcA0WGaSQcUSmO74MgrfoM0Ys2qPlXbBvBsDRIK10nGEHk3bPoeZu4gkT+SVpvK0
xRIaErd+l1SJx/0vF/5d8OIJ5zp+srxwV2ZC8qbUfo3+HRYYzOmj4t6BBjpaA5Ll
itiD6QZso11c51gbZMXVwvHsszAK6X1ZObZ1Fs9pQEiX8SJZIZNoo09IeaTqYPzO
IfXx0qLlCUE0FnPktO+KMlkLPU/Hn2rB4aFYa/kl9KB4CH36jLs5AOn92bnxDgO+
hUCAxUQZKRkdHkH17QsNcmP/yvhuoLgZjPW9j3bLGO3NBuJJR4BI7B2jMSv2pduQ
e697YBy1XwbEZYTpEyjiCMcITc+yKtk8fimrE4Zq1y0IIWc+7nayu3VSjBzCLKON
xtGThuSxPukbVE4y9aYlaTn7mdbwBb+xzd5A0KFeoPp76DQYj+4AkOXZ2oJRyerM
ZQkwsjCOqgVZdmy5n0JassovAPSwhbY7zOydg/AVOl7NokNeykoRjyHSgzoUotqD
tKB43UF8KLNv0QoO/foiAdj6BYF7+6wKrKfb2qs5sCSNt4+EA4C3ErnXVuDyS3tx
soEduVDd4mDDNI9qRUHU0UtnNhvyHCuU6p769f8EXWBawYhJu0CuJO8yJoSGFpiG
AedUuYdG3F1i5nFM8TgQbNjKq7IyBtwHmFAgdL9RNwokHMqW4iGT1OT4PFln4T7o
gBqua1hFyND8jTJ4it4zbKrTb2517wh9Pd5EkPIwwoWGL/pbKFd9yD1IFBvMc5sF
vIVJ+rzffFS4fliu5JAw7qyxoej1JcE8nDrqjOviDW+W9J8HHT2R1xn0Oisb/ZyP
08BZ2STfyFCYfJQhchTzvoe3pope01h9I+2uMtxS/lEN2hJ4S8oAV+wbHBgIES3d
3Zs8GjZZlviBOr52QBGOA/yw1I4Cxwo9e0OY/jylsQQZqPaVehLWtsvuocRjXJ5+
qbjJjzK4b2VWB38PWSmu0UKu9AyWTvV3hqxpxNPFDqm1n9mirjH+fWlmJmo2AQzu
YruWjqW48NbrISHywLAVX4kBGZQeKdJ+g+9htGxbyzoapuJbFidWro942Yvg92B/
Uam7TgbYzDl4w1l3KXgG9EIjgBCor4V8ucVZiDsJR9DSD5NV8c41USUfA65STkSp
wCGePrQO8zbPmUzASjdawwW1OjYxai2nhFKy83UiZhnsRWsHTd8cjH3ZmCoz/zLx
6lvEdSIOZE6RetPP5sQObVzN9Tz0HjrVq3fb5sXhvxcBG6HUXiFKkS9b2U6VRjSY
ukdnpIx3Fw6tloTwiUGPyx1GOqbCSo4BaKy2ym/exALTQ8KPvQsso8+hyyaLQE/j
TKljzb3cYyqgw+bmzCE7QAbG1Qp4E4mHP7p2BpPFOhjs/KLeeFvz7fr+ULNuRxC2
0pwJs3Yq+kZuC3uQL2EvndJ55cK+dWG4QK73YBT1d/zDCmGj+3qjZ2dkRWwJ7BNV
imb6FhVaUM6ueoGZiCNUaZbkwz49Uh/Ty4SkWpO/+rqaZsQEIiBw+k5VXigBTrbt
csYyYKuiVCb8zEf5kEPdaFzjljd2cAgnnKFM3a9HWRlVML6CfOp+mEeMRFyFP6aq
VIdJaWIbcUU9XPUlgqcvRIPZUqae1U67hy+RyRa0TALi0eN6YRUgI7zzDyUl1tA2
woMsIfsWQOLYbhm1uTS1WKFPcHhyg444TcjSTQkG+y4BD/YsnlP+uDiJnC1KIpfl
3wCFUW19VnDSIAcHTRG6zqa9dP8kYIH29CnT5POHFIDaweDGcq/9LGw99MxC2L1a
hQePFoVr/YEv3UKH40YR1oWpFwbcJmPhnIadCuk7WqS/Hp616Nrekab/1u63rnDn
422XCKt24dz+Rvn+BhCq58sU6rLcXPZ45gk0OzQk/XzknEp/VM5O5FOKK2YV+1Ah
WXw3WOCNhgMhKhP+MjR2/S9Fqb6cgVSmDPEQWjhAZEAoArWpuDc1LTSlxCaTX91U
iZdXWkRlAfh8aC7lo0Ym5978w1H7OmCekOujrM5AT2oTWWfsRJJG0yWVH7L5cu2w
gn4tKyiAc8klWwVjofwvgq0hwT3QTkOWhNTxnpPUnCbhavwW2s82dDgvIXhhojRO
+JwnfecLOFFJz7brlQpswwhlTjXPSeGUB8qgjVXW4nsDB7YWUwnZIqfFQFRXRnnk
P2L2yTqisMZNiw6IN3tzWYG9of9O9PkwmRh0ACslo8Pt//mRHm70tPoDsA+GOvEz
JoU94Z6CJG88ZcQLQyLD7W14qz+2KCO4BEV2mmc9IgPtxhnFzeTGBo/jWyg715BA
RvccotNred72LzbWKxSe90S7A2+F0Mc8F0G2GA6ylAcB1kg4mtW/sr2e3LprvG4K
x2LPpUOgL6rqNGqr73F6WQpPWS9rS4wxFKqmsC/3UrTJ0ZzPGgAC5++weoLK35cf
ylCCitFXP2W+zwj5bWBMlKZUFaCoiggQ1pDVKTBHYPItd2ZwrDGfaHa2N1mQ15vT
IvYWCJVuj2bi5HwCU8VtGz2uOOLreS0WCk19K87N13RneNaHU1fYUeK5xFJhg6FU
B65BjgxCy8kjwlytKukHRIvxjAVaQHNaTxjOzVDAY/ZeUL4J+W8HntI0uHuZW0Ks
DYgiPk9qylQ09LgSXv2OUs49ZOOIYwm/gCY+NUX0jdho+Olp4k5oOG/3o7RtprRC
xsQv58A5E0fFPImhLUrxYZMfz8dcrDbez0c7Q1BcVGXVE9X0up35It1BHoRtO5nh
7q9IG0he09nU7FefN5n7osWmUpFYVYEV/qg8AERQE6rQUVR7oDFvpFCYOiUgZ/C6
ALkx4KecZ6vI8fBPrQKB4Cn2ilKKcdKy9rVyM+aM1ESl327bDwZbBkNqmseLB6Uk
yHEi6II3RgP4HHhqzyeG8vcs39kitBUnyzZMt7fF/Mkmk+wkGZyi+q6ON1tdwpmK
tYwNt7ZxQICuNPBlcE01Vg9zcKOFdLSSGHNIYJyerWLFtj09VqFSkvFXGiZUUPmM
0qetVcYcItsZoX/ZVM9Od/6z8j+Fh/11hFVhQ+UAriqdVExBvAzTWgSVl2U5VRv3
/lM8ng3WKwLom4HooxiLY6mKoxU5l+XYdtEl8CL6HJ8koC+nSJS/wUmFJ5U4277H
GLhuGVMNSqqiCNj7LFjgVn+l5AadhmGeQyHlREdnbzMhDUHXggBUTTVeM9akf/fk
ptvGdF5RktH5NBx9mhzv95LM3AsBgFBc8S8RACVjTEgAhQMZ5Pn9rLcQKoawDzG9
O1TvvcWnfV3v4Rk5sma5bClHekJ9eMnF2uQkGTiT3PZQRwFXetrsreuKLw5SDANo
dnn2KrgJxzl1icI5yC7YnbI+sKC2rXE4XG728vMiwKKUlIEkRwqLu3ct0LqNs7lx
bqli4y/mBgN142N24pSHkqrsKCjuqR1RnVDZoVussDBvM9qeg8qMX616RgzCILI0
qjvs/zN83mOABVoRoLKsfr/MeN1jrCnMEcYhScTLymVJwzTComfRY4Wur5MNxXQZ
MfRATMi8FCqpgHNHSpKEjH447IaL+XnuLtAi2K94dsLhR6oswWPlFN2HkbzhkzQn
ss8SlNtU1oQ/B9ccFx/G7v6X7QnLPtcwctXXfIFTaSejssekoN6tPAwGfJh/mfI5
tyJEiJaHtCg0CTdRSLyPC6s3wDfkmwmBhE2RQ8BGudKMhdw82r4P81oTFdFZc2+n
tuUS4xUMWwm/tXIqON8T+vQymrvg3t80jHGlTniQDx6x87+0iaqBkUJ/isuZzpSv
O94VBb8uoyArXvTtOQT+C3fEpvJeVJtbIXk1Aj0e8nnD0EThoHHtCZjA2MA27Uw6
mT29yb5xdSkIs3kX1/9PdjIDOBg+nmLRnR23dp5GXfmRl7N1O/H3Uj9unVn+yMgN
RVvktfR5afwkJK/qdsNbzehiyJ6KujNoodkCPHsTYRoeZaLQ8teQr5zq4m4JvGpP
0lqQvX/LlmkbXd26zqNuDMXwtnNquN3U106GgoTER+GM55QViNlrS2ORdKkCJYlJ
uFxP3Sd30zUuANUZMWpYuuGlrxeAE2cgceBFYzd9ye9om1lN0rw12nvnq9vlJMk1
SbAegPqr5exRnLInF5vnoHtpm7jDcLqYtFB0gPDaYh2YTljPIIvX+wGJ+Mwak8oz
01P3MammPGxpEITVF2PxBU8/hu4S6lhtEb0/SizAFnng5jLv/l747paj6rWptpOz
9BWd1kn4keDOATtvR5mwt1eUpj8jAluRtqvzFN+gKxfr7dmccxM78huB3hrv7b3t
h6F4j7TWJt16kOS1tpdrY3NWME33mRMgS2X5Oa1+W3IOAONRecoDpgUaWv40DySu
khzMAcdMW4kIRIIDTjAtFT26ZRnBbLao9f7SjoAwvUesVr61ixsKmaGyT2dhRf2Y
Vk8fTV6L2/weoRI5W2V4gQjKM4if8yO2aB501a36Q4Uyojsu0SeRjjPzUOh6kvwD
yRvOw3tAIA8h8MIsC9Ok5QNJgsabUOo5w/5UUbmk7tt9huA2sPL1bJc20wei2zOL
IlAinsq77GyRf5w7ZXQoWYMTdUkKTvb1KY1fVg68x4gPozjNpwsaRfs2URw6wk9n
ETrvzwFfWnvzKYBHjqOiLyrDNPQ9UvAspq79+elkjLKtsB/Jc+4bWkg/1z9q/Iid
vzPq+VOBpDOOuipL1kKnj3wvUYZsC29i/+AmZF+my7fTwpLnabu/X293D0LlWeZp
O/F9BD/rjAF+2X6F1iuVNuXdPMw0eYoeOvC5Kd3M2g5ztLMBDgGbM+xM2LNwf3Hz
dHtUzLzSPWRg8xCef40lKLT2axciPKutcwmEieUcsFAz3zJjLN1KdvmpG9Cnlk0I
WZHvCo60kOOrmshnGDj1xOyx0OF4Wf/Gv2NRQW5ky48mCQFU+9kDSAUziMWs4K7j
JBtXNC3JgfwSxr6vjhWGN6J75p65gPr1Ih5WvXd4p+ZaJCLQ5OH3u5BR96reel1z
b5Ff7ivT5EKpWVZFVIzmFoIQbo0mmgMJkx6BI8p5PNXnWE7xcT/b12GtcAHOiqIP
XBN54YTbClbgIaQqoDC7/uINKpura2bAg3dM1yJJh9kEg+nzNoMtS8HkrMcQeBh5
8p0xjxHvRnfQfJloob36JjSUBHGnkcfWkf69MyW3EG4Nhfk32n4jHxp8U6WFuOft
cddcU09K/kcG4EtAR/WYHfDAiHMQmck+LwX3D1rcPzJ/U3uH5jI/Wpasz/bvJBty
R2wL7aAXjBRGq6QipvzZQLbPwY/XPPKyaMABvwBIpidp07Wa8x0LvdEKOvhF9w6H
NqR++sTaR31Q3AbaQDI+/jssiiIg1c+q4MI934z7GeEgNaFKBfCS6o9O5XfwvvhW
tApwsYp0ICPRc6t4/A1tH+ka3wfNeL5OXOiNUjF9rLVuhMzMyoK+Qhkq/qRdjQhe
l1zlhFiF1OQiWYoVNLGfz4lhA8SworQJN5lTqGnJ6UqY+JXuWwXUs383KGTpWfAl
iR0YdH19rMC0WuVSnSXef8ecovy/+VJQPU69q8uEVuqaeFtO1j2Pp8ND/BLROli8
+S6kRJ4SpyWL00qm5dij8dwQRneI9eCroDFi4S86RQj0ERMuHzuc7xKC7wnD35U4
JG6dAZroGUHkmyFfYwyNnp1mJ3qGEF/MY//7het6XCd+PSYePDRju8DLgvIfwCvo
Igpl+xjRyTEwRgFk0TAMiqMrjzxnWz+m5K2n6vWt7wdV5iOH5yG9MaB92wPvPVxk
CBR6i40BlwP4s7IYapki+VenC5bVri0espzSi+ZeqCMQsLAaBbxrV5N6WcLs1ZwU
8Qg5FWUQewep0AViTCucl6AoN2W/v/sUzJgp/E1FOuB049lzQA2Sur0qKi9BUZeo
IZ1e38FCRjxMG475o1JakagIKQLPoZihILfLtBuj+YulopNEFtX0LCdSy5qWNnuh
x1rXtFB1CxvRfFKuAIgA2bzPzTjmAw82WEDZTUUBuRvvtwU9KI6HKarcxRWr2kLP
btxfvkZlspldWMd3fCs7daJmRjx0ML/5WOeBu8cwc9N1coAiylO0z7K+eTu9lirt
HH4+LtUaPVHooWfL/9a/WVdBJ0VHymDa+GpRJqV2ykFtejwpm/GuqwwJC+LgAWcs
1EMvPz7zIf8vdJkyZ/hmgQM8D+tAaz1JPPOTPJZlh6algSxJYCad/KHK3vpJmHfq
egyLdGMw5mNWVT1S1byx/fMkiucBBRWsxhWDfhhOy9AXHLlwHYuLDnC7f9exR2r3
KRmDUf2T3WaDR+U/EqooAneH01DBuAFdDv4fLwtWA2KoLl8WSSX1ZFz1O42IvZ4P
wdavyR2MwQFPwRB2xVJDnYYNfcSPtCTQ+5JN7kEIsKsTrVwty2ibxfAvbqL6g63/
yQFeJMMPrbmJexNeI0k8PJX+fwk2pyCq+jC9tu84fRbI1IxCn+1ffTQL/kO7BZw2
91j7gGUeFlAM8l91w75WO7spxJRJjRrezkjYjq0IEd0yIf+L8FGX1FKxFgFZDXjx
3nDDkdwKiMjXzKl1nx7iVAIyDk2CPlwgqraVtav+34v1UyC2w+theYOEboSAolkE
PVoO+UkKkJDgukk9UBHRLr64azpmriKBhn0+Eldm5FSISsLPwIMZIYUbVBDxtJ8O
2af5YJdWsU/tvjHpafZ+YnwlPS5z+EdOFL/99pxUCz8Djh1q2t5RgMriRUe8sCa3
8y1NQRa/18KuABpaegdbCbBC1RFqZ1tABLZX80s3ZTF+xf935k0fMVUbGlK/BJJ1
LnfLSR+MrtILn5ERH1nXFt9PmTfmQ5eDdSok/GJtNKqYmprncvV2J3Bm2pR4aDps
iM4GYRHq6oUW9lBxDi16DbUcStXYNS7bsz4lXmIgP0qrTDpHksGafmVYrMTcReRb
yGb6hlcYk3QbQNVIZX3trTbVJIM0bjKaP9nGmkLHzUkU08vkiP4/HEEDS0GrBo/M
aIrdcHmezHv7PpSgM4Xa+8ouqMPQd/eyNjQimAHcz8Scd5+yFkzbFt9+LWxFyVa2
eYfeha12WwdkZLeHfvG1h4NAcuClCsFS6DvOiYYPRidgwwwoQuSLswNbAivgxYnD
RV0x+zQKSK+HpH4L5DKwrW08+0bGPXyRYgqk2ZEBajPFlcM09mFKOYMciUunJYgD
Cv0Xj2WgW7MyjVCMIOlzfAUeA014V5OxjAk4jW99nTGUa6wmFIy7n/1KJeHa+sOL
H8mrfk2DxY7e88dsxiAczQ==
`protect END_PROTECTED
