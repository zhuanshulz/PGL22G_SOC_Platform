`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MKuoR3VWgSXDWliSW2YEOOt21Q5TqNRPvX9TEpqfrXiaiO/6r2hHOCA5sho30Nb/
jZHWZ6DuM9NQDduZClZBjFXrce3GnnF2f9NXK+Z9lDJjFf0XyJ2nwiM3+4AHq4uU
15TEsr+F8SuZPExJRUdULdZOXIdUmP5AAnEaZrkQRHYnikAnkuLF3J8pfA+LtWXN
dSXAO4fJL5hek3ask6yW77heCK6kZCxYpNQuY4EmbzG9FHGX4zT0AC/AQrRfo4+w
xa4Y3i6iJXEGZys6vD+5k1XXBDMXsIaQYQIGRkF6svQwtaq/T6EGDNW3GO/JcJZJ
Kt0V9cpFl0NI/jsru4rZMXimtZAUeBbmmKtYp99hubOqtdFk+vdYp0fEvKD9yALE
BCCr25h/CoYGolslOAUkYQKZchyhJv4L0SsJ9lTWzMSx0EhOnNqYaJvJie76T7e5
SIor+zoA8cq3U3OWRZGM3zWVSQzC2cbVec6JhPkMDGe3n2WNkz+Dn29yzLYb4ilL
0D0pHUO7S5Q9iW9msqaPZgMfiEocUfIb/z/AW1VOcSlZ7MH5YrNvhBZX/DwhXwpD
Px5qoAN9hX1Z68Y/NGG06JaW5+pnvHuJ71rb5T9usju7Irj3uH2gbJlMgeoom4Nq
+K8RXsOoDvPyJq4yI+v3yw==
`protect END_PROTECTED
