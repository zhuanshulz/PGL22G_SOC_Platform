`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wyps7tbW+einwtBgay8BCyKj2indn8XkedFjlXIUTbVkCX52jFQcvlQrsG4H7twS
AaiSBNuYWwkf433Ir5kOTB0oncTpOhveg5ZqNl0RtkUtSUOwQQo4LD5DP0vvtU0a
oRFFetDHH5G4hUE7JhEVen/MXhkJBpTmalPDHZ4dBAyDR1lnxigWZDI3EN3kqUJa
Ppd+1qsTKslTYHd5RPsq3IZrgDSGkSmdAwIdqUKai8IHop+xms/YER17WIADFfvp
kJByfT7eFWNkCN1Fy6AiotUw9qgWGMTATSg4xbpBZP5dN93lKF/dNFPLBRaGTYAT
DJN5UjxFQGbRW5F0BK8pkOD8zjcMIItSZFGwVNjXhj/4TwTer5c8JCH3cnIPCZ/Y
HLGEgzOuVYXcPgL5fCGz8XGRvJjY6srbG09lBtLsnBsjxXtazgMMPl1SReF9313E
l1z4uXzIlnqeMOj28d3LOz8bBuLCK70PHoKhzIRubldfFC4XY/Bjmh3KGhjh0XJK
SPeIJu5yC4gm40n5BJa7KSfWM+mVb8J/HDIhaKscVU0El0wmM4w7apcHaIOAs/OT
qAg8ND+0vUmMVi0+D+c7c7D+MvAGkVqAq4gOYo31GpG/4X7o8+tdgcopwTV9yLzz
Xh+EIUM6yDEQUQMEFXT781OVSb//1OyE1gjE8/gbdEywKd5tle4G3cnx2Au2zmJg
xn4IHpDnrhVqMrmnHvCcuyxUN7LbyUmzPz29xPLKnbnDounDQedM6qVVNrXqd15I
gg4kCi9FT5rDPYmHGCzck4Xr6c/J7TIP7MljJx12V7pLQjKt/ADfj+hcC0zTVv+r
u7PsBPjilyey8SSmiq0LQhXDCqPs2Rf1GeHpcq7CZFA7F4CM1+1oIQjKU2gnqy9u
bATvMJx/ekSznt9TaDTZFb0FqSdpjvGWpQA9FM8rP5YSgpWYO4U1u7L//L+mYSnY
WmopdLmLe2qj3yZi8nEBIzNacDMLUmSzkLVuHrDU5a2jzhXOQIySAXEEJtBSNJLW
eneJVku05CB9j29kqu2v1+U085dcZkmlXK3z8+loUFVJbSg6ns0/MwTx2jbXNW7C
ZndKo0GZMrLweceFngNxvVppqJUNTg6Us0TRTBk1whHP1LgcCNsTyiv9x51z7/5W
8tucjl5W24G7zKQszF3uIexV3hO1rI6JfRgS23zu9GaxYj1XO+P5bsSGLwUuKEBf
kSnEXekRcHX47aHHcaSC4/AKB6PbQC4abXlSUCH/quZwTPEUNOV/tCH8kSNGCxTn
`protect END_PROTECTED
