`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mhzc8FRt2MZl/iNU/SM86PmKk1Z+7wjkDRJ+susGwbQjcrJyYxAt9mbQ5cpP4gOQ
dodouyzbKv4tbYZb3otYncwB1s6GN0SIp/xbT0ghzZut7VS23mzvLNZo5BSLQele
Fq48HF/nveK0gvdrfSJyrcF79MdiCV0WuB5L/lpTIK6zSgRTW9QcXRmnPal+aLEM
obEQbVDOoLafF2hk0/VoyEJLgPln0wQ1vi7q0CLi+lYuwEv70Y1ubUn21Mp7i98m
1UcE0nIurZ3KCQc3cscz/wKorFyUsQV9z+7kt2Y95xlV87D9YGBeLYy2uUkGZEOL
GOHfzEoDgtiQFKFeZDP3Z+8S/qzqTFzn8MhFTK3PImZavbV1V8guRWbMZ+yDI9eu
rDqFL4HQYoeNVTLxlfpfvAm59u+9xlprR83LJCCti2e4785dlAkVYXaIiCL5LhVi
sqyBUpPDKxU9W+ZpBs/5sMwbLai04h0SsclAorTB6UUvWhM2BpjsL7AhX8+w1sIA
deTSQAJ1NP9DWsEiDhjRwia1sYID0dfMw4LU5gXiUMI=
`protect END_PROTECTED
