`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w+RnNDipNR/ovjqVLe+5UkFWKINNi2pQYuUf/0S6xafRRojT341pKkYgnek8Mug5
elpfLOOMhzUobaxEAnGy5UH/p/FagO2aOg2L8OP6k9sdi8ybsyYfgevHSJx/XVZ5
Rp9zgFRuF431Rkv1wozlpYfpQ91fNzmKAd08eSN/68jvzCf4BG+I1vInxja9sFRC
Az+oFQHwjRge1Y2nK9vqU+lSAfJnk4r0dVOeuQCCKa5wUnuql2DfFl0Kscu0n+fp
IsDPP3FPfNqYZ2rr8rUsIoxMtFmoRoog/PNX+9T2qrmkRUb8Md+4Tzt13M2cq3fG
o6oTWKH1gVB0/PYrzPyiL/tQaGr5qsyyYZBqrjthuQr9MB0tR5rvMyR8Xq+SkO3Z
owWZFUWOPAdrgctds2wLyyyZDnXEL/optwEBZBtLBDj9VC7TptnAtcO5iqcAqXTY
dyoXrAEe/C4FBZ8oFOUxwy/e22KfNSrCZgOW7IO4cr/QWbIIgVqH9ubTeJ0IFY7H
qN0397LDOJGAljrhB/BV1UbCAI/NqYW2ax2+lmkDIPI8+1M6rOG/l8kWt6FYV6bo
Wkw/go+p1irUrgWE3Ff3Kg==
`protect END_PROTECTED
