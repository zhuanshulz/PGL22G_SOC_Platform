`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hnberDQ3Ak8WcO2Ldq76zJDYWNsn2RH+68g9upTfa6JE7daqPvnEB8xPc/Gy0jP6
Sr2YswKMN63+XMzKkMJHkLCnTYr1V454j1PsLpKB0byIOWCL8iCbnCM1uazgR5BO
oF8OvHRFMf8BMdB+A1dTNUqIs7RBpZuCtISBeBL0iBMsCgQY52Vwr4BQAjHd8xYe
8NqPZ7drfT3qjv4B1x1ogXfAhEPEEJgQtWfzZMVxdp2C/lXlW448UfG30eHaHVtl
R2ISXavanbUDZOXPSPrFEz8m/cXiObFQAcN89be6w6/mnD76fdnItywwAjVO1j7M
HRooKaK3sStsUqhzyjkNewdJh4VN3hDFIMoB6N7pq8HeMXywMcasCN1IyhC7Xzwh
1xqoIbkhHX8lU2XZdw/Edl4K1PXgxQlvGECcmiVMCGbZKaNRxTF1chx+1w+NtVLM
fFGlKhKVLre9VKvIHmSyTAoG1VdsQCmnjkscCZxzmSrEmcyY6knlAXn4Ev938l0q
DYDzegHwOKWnMVOoIU2ch/mwO1ZaZZ+w4MSQTBZdAmtsQSKYx0ezNbA7LhQKogL+
Oko0azQK2VM2/H7eV3xpHnw+d/jnhyNAaGTjF181mVY0TyA3hAZgTlaQpnS29R8R
DWiaBgbAtiwV6nFS9zbE5PBLAYm1XBolR5D2n8RfjtN/DFyL3DU94L9pFML7HNMf
qOcRTI4xf+B2Wpt8Lk/rrAPGdXWT2DqRiTpCkxMpFm8JSWQ82vbbjxN2+Eogd6Q9
rC0w1A4fbXjmDtAUxdeuIW1PlvT/ruMnv0P1Adwsolk=
`protect END_PROTECTED
