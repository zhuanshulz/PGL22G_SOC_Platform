`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7twCmxqKKpU8wFn3OtClnMcvv9Oi1scZWc9Ek3xpPfEf3Pp/x6awOmyE8LTJjAtM
IMISPS6ya+CiOq1Rm9gLbMmVOcck5y+q36JUTsWTXBJfo13hyzTM7wlMdf+QFrGd
Z4UOdqBRWT0ZWxv8OJ4WqG/YynDUeQz73jzEM8QE31dZTMXXfMjZCZ7sMoSqBJvK
A/+zQAPBUWVS15moPrRwQ6xllVgJ0ygiCCb0vqBxGoY01IIfXKBq/X02pEz51R+z
mCeEaRUpDO5bdV7sbZQ6AdlsS8u9dbz0DIwHi3FPDcpEszJKmKthmLqw+nwT8Efw
FSX02+44Nqff7rY05h2jrPl/rGq7rv4KV+jdAMcHYrjETuX7XnLS9HWz3LVFHYeX
xyah6bJuXNCTgnIkjwqNWNrnzNNrtXXi5p/hKvaIdMvWDBoAp7sXUbWN9hgOnEsl
vvBcqnP04ZSKyibidFvLVODxLyO5p7x5MR9kWs9UNUCrNLGBqNUa5p0zejHxlxcy
4qOkStFRJ5lxhG4+MYWfCuJOohRJY54PKYvrjolkzdZVa0DsAzZFcX1Qafb302af
7pj8brJa7qrt3TRvuu3WEg==
`protect END_PROTECTED
