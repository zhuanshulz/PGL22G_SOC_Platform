`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rsIWI9f5rfW8x71CoIvK9wLTlPg8eGTzorlox3unOwXrpK6xqWfAyNUkOBLMTTHM
RB3raQF7P2lDmhmwMnjIqGiyInM2aftr+ORPF53Xubt14w+FnPoUULopN7tgql1b
wDtQlr3+mvgbXUsra4qiB7n16EcfRVxmbt/kx6pDEqls184gUKZiMORQiY6nzjHu
qdSslKkfEFZoOxiSnUvoRxGQ7sV11t/c193qbi+dml/n1OCZ6N16xepyQJwO4Ocm
YNTpuXgT4h0UzBIdtRkJN9/b8i4/2AfoA0W5xbyypyJHXMifPo13t6homj5QQ/zt
FSJw4ft2VUwALbFZZ4IvzaJvxex7tB8WlOLEaJHq76wA3klliIg8gL1LTEZblLkU
2jttBW5Lhedr16VuUJWA7BvEKCCZ9lickQaICM/yk5RiNCS40IuwSKeqTzfuvTZi
lZzhVm6wLXq/Iy/1PP8AJaMy6P/U3gGo0+qwpYP+8YMJWXwyg+TpbqYkmXP4mbYa
A77Ump+f7/3LCCC/EyI3b6bdyAYPlfNjVtOEgKNaXitAKiL90c83pynS3Pijv6av
BU0uGbnyhZE92zRultctFod4yTM142XRV2QqB6HB3nWC1oN5KwYw0WQ3mgXHNOO1
G6l+oZdxGmyyUtC/sKK2vWd3bZYaZjyTq9G0LF9KzO86WtaTY4hUJH2LbYYGavPT
QHOl/GQdvbwlE8bIUsKVoWU6o27qzgUPzvUm++eoPWf/pGH2IOiX0plT5lKsxFwH
9xBVoTmU7nSXssJghbKuqjCbw0c7TH5u8Qd1Ir4NN7gPPIypJan9NWW+R38F8UOK
HN3oLemfUbDjmyAzH14rlPJ0ckyBLLWt2/+SEMy0snCojEYRKOjWsdafHYzCPKzl
2enBcou/EmDoIJtWpTkDLtK/HIqaE2AJ5WDx0cJEUsUbPt5vjV61SBHAk72kHlHq
vDwQCV0HyOJezQa8tWEH3PnlU4qr1HrfigLEcZuWi4cdA26zNdigF6yuAmOSF9LK
zO3KJZO19VsMUYvViYkTT7zUC+80d5qCs3lmdsm0bDhCFlY7AHFw1DsjEVlRuTba
v8Wvvynp6iDYN+EBmxTbuf+xrV+TYUPyrp5B5UTNzr9feUvetEVMkibC/yLF/R+R
94xsdSQuCINsabILW65g7OMeUXi2M1jlh4XoHDmiWjzT7eldei+QrAlzGkhLaSXm
T/rBei5KnuJ5U4IyDWddXn31me6o3RlGOT1dF898+ak=
`protect END_PROTECTED
