`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ebNU7hxrJ30fLQT6IVBZgf/+oe2sp1C1vcjG0QwDSNxepnDDCakSOqVTyb849+Eu
WxWKGtmyzj3PRaKmiz8qW19EhwJk8+CbM1gI2+h+tpKeEzyuq7cYvaEzp0Z9SrCJ
TQH5hhpIhIliGj1O8EKRKQb/Yld8ncqysQcmVvP0fVPHWh9JQao2d0uRIeWgWuzZ
TxPt8FsHcyEkEe69iO1/+7xg5EBzAcOD1b6HSH8+stiAosNj23bd4d4y6b34vb1a
ttQ+WMkP6u0bnS+d3mK49Q==
`protect END_PROTECTED
