`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QmJDTLmS0/OrGcT3kNeL+/LW4QOSDdSeqxeFi7nc+gqtXZBlYZmwdBuMfC3egXRY
yzfDZ62ONDJDMPCh64qTiurLsWMF7Jn8r1ha2lhkrvjdE7L0VLK06JzuAHDzHBUF
2HNLnotzLLWfYYR3AztyBWXrmFJw4USZYrxDyzO6ckZ2dkdDHk0nHJXgvRPDfO2J
tyr70UBF4dtM0d0sz8VC1aEBx34wQXQFk5Cx8uC6J6Vu9+nCi5vG63A4G31qLHvZ
AEwfUDUKrYt8lQTFLyIa3ooOf37il01ZdTUTON2+ZrPZS2wUogEf4K4GciX04WPB
gFI1MeS54cCe9uJU14Gfl+n26Z4NpOLUcGGldRr0uK0nxib8UW764rwStI/ebmyy
lWyY+HLnemzzWhDl4luqiT+KG32u+WOAPUN0NTz/QpkXw6EZEDmdE5EbuQ0ReTmc
I8X4nqn08RrVqerHdZpRBqPZHTJONETbir19H7rMRHR5M+8T8PSoZQb36oKSNdmy
s9Rxu7Ogltpw9mCP+m4ZtW+lSleZoIRjnyzDwvKiPYeoCzGeHAp2vfQoP2tEuj7+
bKJgIQSifHCRAo21YfCgTP4nds1yPDQlbgaIEEEMw2mW6lD8FfHh8kciOhjG6RKy
z5nPist7xtL8t3iDHeT/fMpc1tthzaYKAvkfz5BjssVZAkYPvWvBZjYssYGiqG+Q
Xl2PbNUgZKL58H1ey9zlLa/lvM9xgJCxH9/PxF/spBUv0sQG4z/0+oEullkhWDKv
lOhSH4NF7kmouvhfPKN7DssZlS+/5yFr1cGR61G+eTCl4QSGy7uSxcJYPIehOHQK
sKy8vzAR9dBhoT2yGST9PPB+yBmehwqcOV33x913lD3Mmajmj93NlDZs6T2Dv1yh
pnYaJciknZmkS3KchkENXJND6GetnedESBIIgpM1GckK9FpR/I83KuZx5ZfPjv7g
6Sa2J+TjOsSso8ltppFVKHRSAotturLlANkmCBJ8pSpcibJFVCj+vtedspsXUj95
uLdraViUyNqrgAdeZaq80Z1x5V9XM+BaxbCUb7/pRLrc/YTmh1wuQFoa5xTdOGK0
uZVBnhsHmQplhk167+2u9SwCTAXZ2GRe0vBzKepLuUnyywShnmNmKEVsKMEyfiYZ
IYq1m0iF+KwVBXMO0ozuE6legdlxHihrVVfvrrB7R14sA3wKplfI1cKDrzwWpqbu
sbCQ6t03ai7DXlwr5i4qqTV7XYILwxSCGgWwkWEDjqGSaHLYWDsYN21v/YWSSZ9H
MizCaFceYsxzXrSUjIkcbfnXEsoBn53UHkY7jaz0Xb4kfH8ydaQtTRxxUr5BiJiz
v5zZpL7qCU5+44EnjNegS3fwDBxrCFOWTkpETYYYQNltFCHBanmywVjVJ9HgniDG
+5UH11kid25mtRdjSgQ5Axb2kxgaEKbRJJLA8th8mKGs7K0ttLsP5RkmiBS0UDrU
mu7pBF1VpPJDLGLlpsvOgHochrN4+OwsJDMarzBZ/FBvTUIQA3ceaysCHiikNcKD
O2sLLQAVQSQkBMOAirrNOF+jLzPWHuAVOLtX3uE1d6CeVCCMDPM02ZK+fNhP2KnO
M1in72UwPcvMOfm64rPpiX4FmFeMPfJjTlikDCYlbOP6yRXzkQLm2Gvqv3jTIOyV
C6S8hLqWCL3Gu5Dn2eBWnFSist9ZViFS2X+P+/QZbbLSdoJe+eF5gW/2uQsYlb0u
Qei5GReN1LO/Bs46zrfSQxrIzHVlm1CJaKRLloK8UnbWc2VWfiCBm41AIFBz1xVn
Fchc62CiQm1DxYy4JI5+KqAWL+Dyx7Ldu991VRddkA77if3SsT/Y9kMdsiBzSzSr
HTiX3wd+QYkzY8k+Ypkf19Kcg4w/cO8I6Q4UexOB9kD6fFMHJ63rNFSbkvKer5ba
qyH55F1TqLt4Dmn9y1e6k5SkjYnT64DsAAdeiWWwcCRk5nOwvUBX0m9xquAlQ43Q
YJbkhghtJ5wKLmKoay1tZ7bRydmgFnF+pAQQVEqt2H2sEQ+tpQjK2poSPAZLhrRr
`protect END_PROTECTED
