`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B1iJ2v7fx/SJkaCYc09E6zunPNtnTkA/9KrwO5M4KfQ/gyX+Tb/ADRJD8mRPdRWq
2htQGf34WFCIXOFVxcKYHnhgNeHYpeGF6hwgdEZA9JpKbFf2mvZ6UxM7pkXsB7pg
kh3VYsp9WyvdBD2s2KwMt7ssyuqB0vs0TubflTy54A5JRwEYwg5A0J4jZSPTLi4x
mn3hZ/iBNz8SvZccdfD0GadMQvA2M/ywthINiYHTLbznpr7BRysy+glu4PkochzN
mzsu8a/2I7vYipT4hmUq7QcW1zFXshaUyJRDynNy9UpuSlAlXpylTNx8dzhaSoHE
aIAfcwKG4MI60Z3exbYkmjAH4XFCqW6rNVLwdGnDtUsjJn96EsdzwYZZ4BBq7kx4
bvVTNamxjjC7Ev8uQClHElz+RDTkOai9sQT6y6cD0YX0uuQN3ITtjTsG+ThDqu0O
Mwp6cuob08OBmCaGx0/4l0vc1yA3UqVnsDjMUyH2O0MkmE3UwMgx4tFXFbpm1/nE
4I0z2KJR+mHsbW1wgDZu5SENxZFby07tWEBQ02oeiDCWOInsmkvZOjsMTxU1yOJJ
JEYwwl6OZONDhFAXY8HXuPV1Mj4bDoxhLIlRIK4ipsWpRG5sFPblQkfNeoYFOwYD
`protect END_PROTECTED
