`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hbIrjEbM/6jqktQl3k6wP6FvDWdBodLknUn8mzA5+rbXH0/00wXKEpvTEBlJ0U4P
rvfhbQ34Yad7JrklLR8jvR9OOVpfjCs/G+HBGbUEnsBL2jUaL50emUtUImg3aKNW
DPIe2yexLIcbNKs5hW1LXiZuaNsF0x4isFDqovSlNWokgxcg+RIjCX8cXkPR+Tvt
1uw3qOF8BHpGHpfKSVBHu7RdZOQpFyCMJGK1ckSMJmHYH0CZNSyAoen5j3O9FPbU
svw6jxBsxeeIGlhKcz4MeldRY2/+WiDwsI15xovhXvPZGVHckBrTdqxT+37hKwPO
pgZDC0cuJ7aVMutjLhCnpddwIsf12PVfa7s6pEiv49YEtz0ejWboOiaMF4FHCwlw
5/VV5EyzL9usvxVAMeEpr0fAqm067URKBYrQGqN+3xXbj5CeFtPZ5B5CwUBCOlOe
fLKQ5xLTObhxZX9gwZvmeXjbqRkXocMQtlUudT0+l3qYGjbQ4ibHrb/BOmZXsthb
+g5YaEFh8dll7XHYFh4rmkaLIowJ+99uW1782UXXaBMmSRfkqDTHDxEt0mXjRQYf
IUB1NpkOiEEf4lXyyTwoG4o0SUhwBihGWPLOdOmSA3X4XOdtVqMnPnluVDTI9nK4
QjMA+6Mvi/dVy9aSwrwOJlm3EdB2UILK/5H3Jt+FJU4mYDa9z9S75poeLLkfWDwU
zleXjtjGHyL87Rrx8rOSv0BWw10yJ8px9hMr6Y+FCcHgEDUlT77k31QKyFFCMReO
M04GaFAxqs9u0cuvJxKSmAWWt/tkOwc7wa5rBEV7mlPCua78znLD2bk1NpmM8R2g
OTnFb2Y8oyMXdMwLK8Zr3ZFRZLoDTj5ILqP5qg1FTEJNTT6FeUZ0HoY8lnUmvr0P
esJuM42gTelOoC7BkBOIr31WPTplE7xWwZi2xw9x30ognbMLpZoIn3/qyzA7tzJY
8u1LGwy0B/MHkgG5wwOCYdkmId2daWdie/DK426GPHfOl+Fh7wvBr/JwjEkkCpI3
LcAX8S5juXq7lIc8Sf5O8NTLT1woa1+lBgzVyXdyquZFx3xCeaujxaHJT0bXUrQU
8Fwm6e1QrJrXmm3jUuC827bW3ck3Hr4KTstBYq6gZLFFvTDImCLBVXyzHyzVe6AY
LU8ZN/41F6+t0MFb7Ud7oTFzNBvaNsKpXpneEuEVG5y4wG3JwxbBtO/4OevrFdzV
3V0EdbUA1GqiwnDt+kxYVcC1MvbtiTlZ8d+U2gh9HS7wzOETad54+L98Vwubq4L4
RJqU14E9zCnW9vb8Rf6AS89x2ELg4N69IjwAOkPCSkByMiKeQtRJcDRehvNC6Feu
WASQFrHKpICTu6c3kaRID+eWShq2qXzfOFLMdahxxb18nkKj7CCpAHiVor9dl/So
QqSGakKvzPWiuZWfyJsgy/PPUtEt0O5yMbEFrvRIB5uOPZaDaesOxQ6Ktpp7Y/IZ
QuuEjVlIiMLxAvHdEaa0CGAMUFOAazHt6aU/sU1eeWdqQtmTmBf6MPSo3hW+OpBU
el8/U1JjOezDUflya+dtAAEf43hV/0hEmaSYn3kpaHK7VCIfzVtg1xZLx3B0JxR5
CcOaNlonbA7ov9vWwPUi3JdW76ZPOOqrSbgOrtPj/zl0g/si/F+ujOqW4hRbOx9A
QJwIoZyXSGgj+oUJDySOykGY3kKszt3uWG32MgqXyo5kSdEhZwiFZCAmDvatIPgD
73gcXiN3GU6hLAx6x/KYMeMwcFuqQd2rz1WuroZ77WEraN4NYyDvC2gfRmHM7YWi
u8us0LSR74SvMIsMMAZdHitrk8yLiCebphw/8M3Ph+uzge7J6rR3K+xMzAPyg4wV
nKLI0jxMLK98/VUQzXhy2soZRbsSBKMJ3u+f1x71e6OO6BxJ9umBadQ9VjV6vSSa
vLZX3gQQ4YG1Y866UimCOugh+xJztpF/e0/zc9pWXSX5mayuXf2Y0GWWQkXESf/d
O5ihPkmayyIOEAnTyABQbue0O0jnpP4EW2UfREFz7EWxyf/zzcibz6ubdxd1rKIb
+B4J159bCTLDMHh6Dn/MDq8IuN0vEeD/Po6uIx8VQ7A=
`protect END_PROTECTED
