`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F9e/vZDsWK4GdfZNmnjA5XrXzmjSOp1rOdLNkuDU2eaFp/la6TOsf8SlJ+x98kGZ
4QWazq8NPOmxQU+O8l4Qliaq4Ty4Om/nlWzq7Bmv6EbMy0B6YIQqAqnstPXE+cQo
IkhBq2tq/j4YMyYK9zm3kI22B7Y+y6yq5dNJlAiyetmEYqacwqFMwV/7af+KMFrK
UjllO2+RfNimWMBFOQN6VgR1FdHdF/CwB73pazUphQRFAhuX9h1aP0vu9DUNnfwr
bgp8RHnX6vK9YIqT1HeISp41W0ut3TtikRvZv71djCjuGASmxYKBTsXX506zx18J
+rIT+iQGs4gcrG7SPVOpivB/aOFy0aRiW5TmGAiwCo3Gib1a3z2nRjihb+SyItNF
Emlw8LIkjmDCpMAVeUVSXgU8RsnECpJ5nr+vMjxK7RK2vkrGmxn69LgFB7JdtiXN
bVB45K1P6VWrr+bmqVhjcA==
`protect END_PROTECTED
