`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WT1suXeHMBWKSg0qor17bqjXRdikWfTK96+bpNYqkw+3G16GhKX513KAm6+Az1i4
fN0s+ajOJaDm//gPDSwNMeTdGluEJX248rxp+CmvXLInT8wgHgrhv83eFWMlVTB2
TrBF9QVejsCBjLLRDelP4OTm27a5JvUNrqTJTlupA22ex4t9JTK9uVu6CeXy+Z5k
Si5oNdF09CvlczgfpKWw+JdMEyVDG5tXzSba5KZTRUCKf71PMhnUtWfZypl0l2r+
+PDWXRQTHgC8IEuvJZUD8QOzL00CNQpamHIftaDX2IvgX3hXPwFSJvqwm3zEvAkU
uJkz6lzzYkcIYvcB0PNPUbt1pLDJgPIfrdesmNM4DyGvz0X5JAq581gvfAGXPsIF
dXozWXA1lBKvp5oCFIRFr5nO+XYaR/+WJ65M2DNdsQZgV4qO3ol4UpdZ4xrgqubR
GgbobIfgFINy8rSYHGj4EHfonC6LIG4er97pV9RyQehYcLe4OLfBxpY46J8B0h/d
Pr3J876bL/nNkjJEF9pcBo8vhpoJjqSK9YiROp1spj+UYrbo2/RL1J2BCUsUA985
DJuHMbIae9kqnsVRxSV1tr7+M7tp+2sildpmjD2MX/KDMygnuUFjret+7bmWreZ8
u1+74k3jLZOBs84giOVltIltR5RQC21exwZGE+ldAknYjzj60KBtHzDmaGtKNPg3
75SiXTCVx6H9oyzqWIIVsm0kqinYkqtopOop3bWCStPhUfLCP1iAV7bBa7T54pZH
UTLVFRXVqJb1LizvonFcIuz6Su2W25li/LSr40Y37/6nyQKkfnPOM9CFVF8buBQ+
5log7bMtiYTLEn5cCsZdzd82p+zDtTHoiGqrRDNbX79nDJ+kpIR8f/3kLk1wGiZh
VHp00vmqygs7g3ch1JQXy3RduOHr67zW4ecLLJrrT/jtpLSXyHBGiWWjM+D50xkb
nXJUMI6NTokKRveuBAhPDiTkiQY3uXOnCK0qU5enr6ANgrkVFwBCz9czrjw7pQgM
DwUjJu+lluD7pnPuId3Fi6YtRJHFO9sWvI5EcuYPvtCZiE+NhadfJceks/bwje1A
w03abHVj98NXf23+17u2r+VQwq2F1Y5VRKcYRXiF+o+/Y9LtKAvcd2ZeIKxFaRiv
ZDXKD4Zaj49T1T/HN85CcZ6i9rBPHjWXpdGCm2Ls6T9YKUYGxm41xIxmtOleAI4Y
/qSaWlDgDIndlkBEklkwVrkerNT+3mh7lJp4ZhgW/BhabEPVveO+lN9NtOH4hIz8
vGUF/FJP8dyTJmemNfLXHPTfygETasYWZHh2L8WvNm7xTs0rZQautEX8IeOn7U7M
aMpLi/G7mKFJDrdxjK/goeSdLu3Vgs9NPhdBw45JZPPWBLycx0wHCLQYm3rjRMeK
73dGWVJrLT1XscywC2dPBKa6FWmafZyqAIBdigROkgV6nKj75U1gd2G7Jk9X9oyT
iXMaP+mOqpng3V7Ky1B+wyh1DM5F6jMrmVKEoiS2txkSepjG8fAm9ecymm2sD80y
m+uDJU0jRnZ2VUUrSsDIWr1KJXba3uBHqcYKN+vUUkL8w0Dkf9TaaljAiY3dc54y
TICMrMQm0TxWWQVoGbJlsJ049Ys+RxRHdn4z93z6f4I7wK+QB5YfPWo+OqVdGNvl
DJfDsygNUlBKUU5ySq1l0Wuln2188NywjOmpXWDmhv5OT/m8Lz4AyH5XbCBGTzvD
VJQFNnSYsVmLS0ktAXv5TrsTp1DrLjcOWwA4qfL7LLmTwjZJejN2l/FIZ/RX6haE
5+P0HCDMFGXY4+MemzE65w==
`protect END_PROTECTED
