`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VDWuqIU42oAgo43lKLCK4k5V2jk5LoT2tRphEBNxCQw+WUjFqCQ5QNf+2lhFOF6U
CExNhsc3SYlRdF0dvGZnMyKZL/+Wtrk0GXHEUhsuqPWi5JgYXEGm6gNlGIvd+gIu
vI3qdEG85K5EVvv3O/hinRcwW2yQ13yBbPwI6tDordCYydCmNB0JYH9oThZH8WVn
hRYavYXbwrInyPrHJYQmCxRUP3YBwk5bG2pt50kEnnRcxrhTWiCuxGa3SDWbJmGE
mde7++0Mai1bYz+dsRRD5GHfajuBR//djfS5EZRzo9XKgTSs/g1TeETVYpPiaHhg
mJRBqincN8aPWIDAEK9ZBlOelDYLUHU4dExXzF/k5HsqJrzJySnnaKvzmg5q5+4Q
nheeC/e8A9xrbEBK0rAgrNeC/36O/9qlTon3nNzkfUYXHdiLkSmpfZZgKQNG+v5+
dSs9PmdCbKWgh/yoHBog3kXzwPYQwVOsooCWUw/47eVxshQw7WDJ4NH/Qax3CzEo
kLO1mPHkBpYqRZ50PDHZAcNikriYQVqqOPEe1UDm/x/zaAIonLfJiplfxwY9HzuJ
I2KWPFX9i4ZwDRKJHx1KlgHEUQAP1PzXdhNwIUo8zcUophtrCC460IPrzDQVdMld
xKxF6syhONDzPTnvbao/q6k+CPvbT5bUhLlDZFg3AE+SQb11bHc+BXoefaR9Ajza
dXz8j2YnorHicSh2tkzxKWB3yoCPyRPIEg42iAtRNX7rYV12jI5Iln8oDa0Fgxgn
VKICE5bpn4p8qxH6LLPP6B0vGoYJ741WB8s8+pNroNDHhFipyUxJuMFIrKd32yo1
Fo7sG0Ku9tKotaBGidYYWkb2yU3ucvX+IRkZy8YjHnHImeJZnscS+CA4wS1zvUjs
z0xB1Sq7bmqGiHdGDDn73oTJnB8EwE5QX79RRe+IXt1Wqe9ZAdgPnQAIO9VhVffL
Ak87ykHx151mxrfYExQoAUL5MsvzWVmM43rgBI8a4OJ+Xt3IueJ2umS1z/C380X3
hIpN7IriHk0vB1ASoZbGycRpjbL6jidiXSDDjc4/hJgka09ZRXj9diWeLiUVNayW
m91aQbf+QEeRmakvFJ5Bqrbg68bjBSt7D1T3WkSHjohY4O+TrC3RjHUjo4mkA9tN
v8p09vUj1mvpuKefzlxzxYE1/kwAB8XLr0By11V/DVDAjb9D9JPRjPvw5baXrFJa
ln7iUnPOfLIpcMbBeZE99fgescoM0fLTJfAOB/cyQvFx5rZFMmdv5DiiyDzlRTht
YbbeMs5fbp4QlygfV7U2q3gKuMp7TmSOdqG2sdO2N/sPKVMtoJpIABtwZP7r1cLq
f1uMinPr5Cc9uBNg5JtQxkUU2qjMCzwq92XQD9n4cRPEJ7EZfA3jaHoplSaJtjzU
98QnU65+2DoydmZHVGy+fgsQriexmCsn5XwCqpHbMwMBpfeKUNw+bkLXo899HnZZ
tHQmzsjveuyXF8/ARqiPNZ6/dihaHQb6QXRHiFHmWUMZ6B1CA/TnilAagUj97Zci
JNYUPFjgNxPri+mEE4bT4OsztFNAtdnkEtdt5Khsi35kRxKgPX4/hL3uepf1XFXJ
A8Xp0PSxpuVm6qFytH1cVfbIQGXdc4oS7VrX60BqBnVm7rbdbmsd0uq97ZPBCU9B
O97RT9u4kPhPpbQB4sntqlaEiUYEIJwIpXGr7dRUmzQP/ALnZbUYFgJPd5HE0sZH
aogXZeYeKUpPHlHRUF9hlnB48Os7hZjZ0R/IO0Ga+NS3aSNduRSRZ7XXm4d2lNJF
URjml5b04tiVwWOpFjBYygu894x7C/DR/0vvWpeeEb3OfwbBKeoWjaUqvGk2UvNE
a2bBgIcIC87L6ig38hNJ8udy6ZAQ2sOHN5+5NrIpvyJ7A5Mb85LF9JaNUIc0zMbe
R5QJy5luZrO3kCihATiq1c/cMnoAegVjTexFLcz6Ryjkd3FSHq0F6Tye6/2Bof3A
GqMS/MxTrfbwQ1tt9vmBwqdVVxoXb5uZzZqiqpnn6yYSwkqi1mCQWnQL8haNY+f8
ye0zpOqEiy2gs7E5Ay2oC1LVv666pxpp4p+X9VO1/S1IExHZx1SYc0x5UrAqu3Bq
tRW7tQKVZ4J74aP61Dq1qsOuQ7gTEBIYwwOSbbXmXwnvL+ElfXoKyafnIVpXW91m
E2AhModwSLh1jkDg3voKC+dweeLPDC8Ur+sArAvxLmbHrPwIRrwDiFgKaRZWTGF5
gLhcchaSszt3Dd+q40HxkGeSuH1A+vBmIPmaoQOXCTE6yO3gMARSKH+0BAhXf0eA
zi2l+lsUIphLHrZ9neKjBFwps98hXZx09Oj5aywZs7jr1GZ70zibItNfFBO8YXZC
Tncjmb0EBVhgm2AHCQYEJbdLJ/v20lgTklRZg2prKlT3yFnIYtG+rgw+/dKE9x+7
grUat0rK14woKR3/N8t5lpun/pv3uiRsmgQiboZrB7mlGUsY33x1qJKls0GGQcvB
scmzT3VibEbxgJgpmdbywx9FS1Ebq3qe2zA2wd2CNoWbOTfSukbdkm7JjFt5mLf5
CfI10Skz5BzFzR2NASEBcxrvIgS1mdiij2vHYwiLDxrP6302XT5PEGd9htNtKJR7
AIFCaHhHF33ZzTT2wR1jUAcgK5zr8SLXO0/tIN7Pd9TzyPEr5tBWWhcXvF5QeRqc
i15o/sw9x3seFe7NKITKutlFt9csagnCqq86CDPYxEzO304JEp0/Yt1BGyyFzDnA
c+cWMhhIkcwYJc/OVVNU3jwgUrQ40svV6uYnA0FEYlnT7tBMFIq4mdNWa/eqx5qQ
Et1abLI6XLBm2j3FlfTDZNLRhCSzhWbr2VMLJ41zrYRbRsnD6Fn6EOwXhqpzp9Yq
h4bYK28qbXZpRIljSvXuARTA4NuUy5DoJ+T014cG5ezdqqDtKYgRTTRZEPjepAs8
KLNCQSZGlrbd0svaT5xg+cM1JkiXxt/euZfj2tjZn7z+SOeuGlMQa6UUfXJw8Oo9
Yejvh7CzM1eIrz8Z1foEorReoXl8ZkEbX5wtawvlj0DNTp5Ku7qAcTQT6LeFq/Kt
VhmHj9hdHBoR2ZuGCGINJkQXonqeyUCA5Twgy1DbNZONo9uk5vksGPggQ/NILrut
w4Erjqs64Prm47M9DQH7iJ1LzIOa8oPaYHHpQvFFWJf6Vs8pqf2wmlktdeFSisE8
CSa2sGu63OIhm/SEMXZkLAY76ksLrZ5P803BXZYfv9EH2LrslQlIvQPWlq+hXnVo
Zkr9zMdro0hsNFHM8sbeMf5LEDqzH92/diKDo196Qv3u+bcKPq38h2+awnytI6p3
CTn42/uEr8AC+ed0zBRv3bjrTwhxuIIovR0rxPRhV/CRyJT5OFhAi+VYJ6SmyAep
VuiFMyzAuEvU8VyaNWBZEaBpLlCaAM7gryq7iiE4wd0DSp6KsDq2uE+nQPLFuawk
6vpdQ1ZHJCYJ3XrRHHG1FUw4YpVt+VQiBeKIb4UDS332Z7xuu3lcNKPnkCXP09H6
xtJtzJN7AdcjOWJEBAp1/T8dQY1JujA0zAeIeJQabxDcrE9t2SdNlLprc3FfkWSj
B2EAIZZ/LLioYPBDhWw87cuD89glbOMVeYHzw1njSLvBnBvyrO83s/NKYp98LhuC
0R2Gnjz3BXKW2DplyeYaHRuyZPalau2dNwC5O7xNon5b/ur8VlCLUa+olEG7v7IX
RcjpXUk/WfbVZ0yboqLIgOFc87AANC0ACnUBULEMFrS61Ucbf+hGEUgeX+nPD1j6
juCC7dfwPjjvGMKIDrXR2RWYLGkHWIc0GqAOfgi2B9FMsn6rWyWxekAAfyp/ecR2
Ny+Q0IQkkNMUXWPhjxPRpyIScQ/vFMiEKH+O8aYge+uTHUxnMvw9A7JqRiXS5GUy
nJICbGTKrN5tebWOOBMLNTjqjvnlph5hlQ8Epl4q6csxIWfltOjSNJSXw/msvoEr
Yh1uavk/XODbsYi2W8AQ9U793Q78URTZDKaTgPpp6xkMyE05qrDBUvX2tct4/zTH
PXccEYxXHYrxV5nzf7Sm6cvMKI3hXWUjNlSroiy798UXlLtPe4Nr3ZbQzYpRZSVX
LzuUf0JLfIQhIpaEorWzPj0d38qrgEqPNTaefOOY5vaHnJIoZTfL0vsjC4X3JilV
23QchVpl/NAo9awlL+kKhVDi2B8pMeO5kSdvhWX5mIedjVhxBUbuLkC2JQE6xmrT
pmx1zxCrSS51NCSjm5DlCGtflhLbNg0rAeOOEyp671TfVjbQG+7g5B8SrIN0cvAB
EPnkreoVSkVNRN/leLUXEqduZZHeS2PZJ1tV+vP0Io7oKyA4jM+WxjJDAfw9XgrD
YL0wWYZ367b/5SZDFKz9ggEVpY1J5aXmQLZURHymUs/ePKaVKlu90IMUOkoW+VEz
7vwBs+BseEFZ1MHJEWeEw5Hh7aPjHVnPsQ8eABlUAwVn9VJeO7m6dau9sgBtkzvu
cnoBplPyACI9GUMVm2PhFVYLDyljsM7NPqazhoa9OCA8eDAujCsfR2g0VRPuDf0I
GBalGDZz5egOxjEkwRtknPzbVr4GjRhMLqMkgC1OPdRhzBJUcLUznDDGFRIOqUyg
EB4bhxVDuSJU6mr6ROGfzvtXYaMQ0WsRtVePpRjeB8j2M7Yu4iNK95/SvmjkjHF7
8ePEGmXPEmvXTiEyPuYf/vwfRuW/47vUUafDB8khG0q+QKXrORh3chNGbQlpYHqX
9y7Dk++XzqxmQVAES8yFzzG6HMeaazzzr7T3OP+N7xiQ1/tcGwd+rpjuvNS1aJkY
T3w/IczLFImLK+9zND1SyijMVgv57nbOyfOGdwx3a1lJCb+bBlXwHH1qWVsYvzSk
ny/l7WcRiC9WVxlNDClUsHSG098KFl8umveEnQJe3AhTb6UmfhjYpSU4v1JRG+QR
W4nax9dedYrFUYS+9wU7SCHVaaVUXyj6vgNU5nSLRIpKm1yNefgPgkdwI8QDVpmm
yB24qxemlrqy1o2E5YyqPVRYrnzHggCVaNDmusxhMh4ucKTXsuWKIkDaFc/aE0Vu
OpTVQO+NXBOR3rVRGt7vWghHEGDloZytoQaY3eVSaxuM7MyZWAC68NFrrzMgNW34
o0q9FDO1QmbWp2khR/7kJQtRb0mlJnEhxlUoh260T/fVFyHA9B+zBwsdKfhxF9oS
zoLOnu8xMVARkKeKzvWES5l2DoeIltzbRhYHGHIAwXsXvPgJkfVFerU52sV+tG/w
m5PFDSIv/cldsENWaNkifveZXOblgbb42LHOC2QRR5ca9ezWKoD+5vbT/SPcpeeo
EXsGl2USLqwZRhVLPVV/cM8Y+LoIWNrLsDawbto2adl3303lojT+8t+1FTk2bSE6
HHx3/+fqE5XB1OuleBAUCeAO2+GHsKEESRV97XtpcLyhYC6J7sWpaDjvDb3HfOa5
GdAzW1X9Cvk2UpU1S2h4kgV3igGNseXPIty9IanEXVNK1lwWq2hJrIIFjSb0h2k4
0jrpgKBacGY9r2kcInZZ9iDFTnulmUNEZv3nqV0UDhK43vTxoZYnUOJfyuNE0sCw
c2+eVWksA/NlJKQg4SzZSsYSMUwgyPxfWgxy5axi4HjYiX6MsrGC8oaN2lTZwB9D
aUx9VU8E8zcoVLgAEDguWrWEFFYrSCmykORqZOY6Q4gsxb7ej67zIASwDTiNxQtR
9wwQLt5wE4m1WoNSV+4pF0HuA9R/jPO/pR0F1RB06XmVqTSokZ6mf7C/5e9DG1dr
JDPVW3gE696PkkW6qy/ULwsO93juYkV8r1Uqm6NZU68v3VPcZH/clSKw2wDcqfkw
iTKh9HRWFQIOLpjy9idPgE0UvmS7BuMGnnAQqfYJhGp6GdQ5VHZr3Ze6jkEd0sa2
yvta8YfH+rNwAz7LrdjBptpjkeIIEH1LhZmsDCnOEn0x4q3CGJos22bD7pMBPJOw
ORIx0WJnkOpYzewpym1OcCBa3jkEvdY0ip9aLEtWtNF1a8aqg6X+7qeJ8B0LpFQI
6ZcdTobjN9fi6QzbbAMuj2ySZvR4KWWWkpxmIJyv+DT3RfUCNBYd4SGDIfa8q0f0
P1CyfwwYLxpF9hnxs8eMfeizQ/6nV+Q/yYcxI+RToPBkek/oZLs9VIibFRBviFow
REZLKBb1ryXGFlFQIwvzNmJRxjPHj9KRCYoKaaSX4PBrMqZ1dTAXPx7/1/naF597
RpjA/G07dFD6890xt1TywebBYF26WxhfjMx9g/TiT5khpFVTfkbNtTbMO8mNz6Oz
nXEgw2t9xAn8nReDHlheCUuiRasndUSV4xvh7RuCvSe5LOT0oPT2qmAt1jfeifTF
exW89SXg4hE/eTJqOby7IPgpGRadRl/Gcx5rBvqUfcq1mqNtVCnZbUIadexavNwP
1I4YDysSIBPeorQVyxZqo8XgTPSOCDm5/Hl/JdffxH/nr3XLboDfQE/SCfS/0H4o
RASLeYMz5WuHQ7OQ0Hc3ktsqk9yESB9Zz7xXpc432teUfB+oxb9wCUM81RVHh41/
2ip9ojlF3cisDF07QfCANuELA/0k1MvFcnoMUHkeAjI9H/EBGKy0k1cbDajtFnRc
Wku9WMJLojiHU+0VOIdxFJzXYBgpJpl9kyofntewpBHRXdWuuEfIjohjQt9HATSK
0hGsp4blPiFd1NtOem/5b0f5vocQZab4ocz/wncPCfpwGfVJ76b+293nwYBO7grv
Y0UOEBtZRlNriHkHW5DKJsbNgKXhbrHOM5o1/N1/NXId3xdywXR0pWIps/fL5bKO
urswxslV67odFtD9k1OLIoxIYnHuI/Icuuqyz7lCk8ZO3ZQBUvQSkIjrEf4mj26v
R8AGVpLjXpzQaHyQ6F3XaCrC39UTiL10MjE796ccAVw433dEsW+4yIpHs5+m77FC
UPaNOW2bdfBjeMgu8gOsTRisYaJqKCP+oE2klzI3umHYI4sS70hLmLXGvYpJHj8U
JMWR6XKHO6gKF3KaCSQuzvLUEFgzgU8Al6F4f1AeHLW4yMYKzOt9lgYFsDx1dZkS
C8J3Hh+VDvUWcL+FdPshkid3wCjR+TXKlzC+3KTNvJvVUrSqAJcFAa/SVpwlYW+r
sJfi8byHwt58GsN9hABOq7gjSzQo2Xl9sJ0Au36sm5Tkv+LRaRdQ89u62iDEvfNd
Py9qFfZSB0X3CfI+CvHit0YHR5Av3onhEWPRUVnpz4J0nr94mlKtNNzgHDD+wHbQ
yKkRP5TFGH1INw40ZcQ8sz6I5qzWyXAKkZxW0JrgKYo777YKptr7AjoYxkgqHrc4
n4khkhFNDgHdR28WpaDS23SKYqgYYdUESgsYszZWnJ64CjBY/CUkfrZeo+BZnvom
Ta6iKxgg+h/T1AsOwheVftzWoduPlM9JOow5yCZfd12NrddXVl/oeQLA2FdW6Mmo
S1GJJNGI9rBmzQdmiZ1r6JeFxckmwupfyM84ZXttZJDe6LB/6K2hqJlHpgcXIcee
3JLJ3OZS5oLkA4EUppscYfPbdl2z+U6IPm7o5oi9OcSOZUaaj8X+RvdvcVL2X15W
+BASHKmZuD7P9AV4jlMGCzeCYWKfZL7Ggk7HZtatAu7I63KPM/tefNQPhdmQUgjS
MIGaQRztU3xJuj/+ql65E8f58EvlYSHy9v59lqHh6GPhOajIY8GznD10STd69AZb
Pdrk8eUdjvwsJ/BOCkTAvSU/eFzDtTJnUeWgwWvyE/MoRN83JXHe7/LHRDjnsveN
moFgwjZrgcsDibmLC3QTcWLZIR6k9zc5Kl1tBilpT1BhaffyLFf5+arDanzm9TnQ
r+yyPANIu7TD7vxFzes0vzaewQa2rCVQvcJbAzSE0Dd4GgB6XywLF87Mma1DmueI
bM0ftePgZR5rLCPj10Zs1FS2Eni8Iso7S9cLaGr5MWWAH6f/DNRqaEWazWhLLDA1
hT+pyZsAeYP8upmI3MOs0qWjXPM1AZJZWfb/UFKKPl2AW6LU/zenHOhPcTKM/x6b
LyBqRbDTTeWf3DdZm4b27Hp4PMoHmT19f6/k/1oyozoYORo88NNFhkkTiQYrlRI3
0yRuTD0ABUlNQoERaA5KGI62lqKXmLBeXwfSqfbVDFBdifJOsMPYodN5h4g6pao9
OA2GAikU6pYXrTu+AR3XbR9HQ200qKvHUAMmXiRzcoyB3Of6X537qplAW+VWGnsM
s8IGmzNpNK8gBnjZI8v1s/1jrO8cccaeBYJcclrHk73T22mz40c0C2dNCJT2GrVE
kJLhuThtKGMh5tNGJERtAPVn6EYinulo7NVHFLw0goANxMy3PqtX9xT+3/LTZVo0
qn9N5ok1k2zLbmsZC3XfcjRt0bfGqad9AaDMF1tQ0c/MUlIhLAcbDZt9xSP+dzIP
lySHWUJjk4wh1XSvdpjvKbGaQy1z+t1y6vL5+3ej+VRJnBYpUf2Dwd77Jb2CfR6w
DmvxdYFPwc2L2QfHkdyU4cROa4/OvG+VmeLZiMxkyRfAXwIwvEa6W+l84GawlK7A
EeKDQPrAMYWZOCtxaUYc1HDaaDbj+KV4VC65AXrDRRUpsogZvk1ahsJjPEkhO9l9
3MvaxhJQdgkkzxRZ+Oq4DR0GHNB0kHxvCPorPHeWA2qa6MDp8+bwthk41jQCzS88
HCQyfN8WYedISoHWvgh+XgMURySCYm3I0A6V1OSxSdjNPJV4B/+TNspCzLJj9S6i
ZjDbAy/SkaeLYnJWvB3XowQwEsILYZkk5u6V8iPHbPnQl702VZh8B5LiBPhmW95K
4721ysoW1o6yHMJoWas6TUevtdyAEwqbxUItjRk2vpY=
`protect END_PROTECTED
