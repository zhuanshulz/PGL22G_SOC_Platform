`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9dPvv89LedYnmaPHtsw8gb9d7zrLjQdHLcUIe2PGYTPgEyzz3uOy07GbVoDAWRZb
+SzcHZXSRSa3ULj2K0TZFoBB1AR1+cC4XFK5RMZ17GUSXxk8oHvNJFHAy2AyseSG
J0hD6DCtWL7yXZevq/nmOZ4YgyPWQuUepq4dgtCWgcUQLxalpzDIaUkjIBP8a7HH
uaRBd0xvT9247Cr08JnryOMDTNeloRATzVt+p+PuakUfJZA28B7desvsNb/M0pRY
+mMGgcXUkSd1huW/gYddqWtnpdBuc+0oAsmkZS74bS2W20HVUj66+BmQUgfvamAJ
DH6xCYZV5QD6vBuk/0boAOUwDMYiMgvov3QC7Pndx5szCY9k6E7zeacq72v53FAM
SXHPU5+heSGtGnTsYOsB2VOicUmELP3sUj4oyHVXz19ZmG7mH6GGavLqpXYJ6RvV
fQ7+pSCIlmYea435eWxMWLURP4yrnUcAFFOe9RtPnR97aDXnQT62EWOsVuigjsmr
P4NHtm2luQOQX/diPiRHaDNxTPEaOUxKzwzNlbddUN1Cg0gf++K+KkKzMb7P21Zr
4jnszVP9w6f0qVVWgXEdFWR/p25bZo4Ekv6q+ae/DQTde0QciLeQYwlVSSqPGIYU
O02IVT418kY5Il79q1jrHYkGiLnkRb9PtQyvfuQXjonQ5xc19ab+bF5kaT/Fy4Oh
MNLZci6tYuSBnbJRHXCJgiZ9421Ca0peXV2aTWnYDHFNt6Re3lB5zzfcvAJ/bv9n
RGk83DJTCvIRbOpSxVKJSN+3MjGbvZ/92HEX9ev60P4EQPlbPOcZ1o4jSOzL1fw3
41QYX9mivERtho6sUbwS7RfRi0XBe4hwmOMyMvgPeKDtGdCgygS8lqI47OKcte2l
FJdFYanes+LNIjJkXtpgN4GmN2goS2VGNcxag1rlBXMyGmfy64QUkxp5v4EJGUlY
BKu9mApKj2+22NQB0hos49Q7rosdSotaRFWJ1F9nzdyKqezbwb46mL6lwedK7yjm
TUrcNNelfZwSdWhI74d6ItN9FffJ0IDSDxMhX2oZBZbu1F9wbB5wlSf4BmVNUaZq
pSdX0vD4pXdAC+Gg+l/eRsVD5/WbjpAF7/dEk4iugzuu1THgKHPb868NH+NZAanM
vOPDY/nfEEdELi9FjzpKEQzpuQp0QupsWowdklcCo7CBCsJB1nPjfYdkGXgoXMsd
sfHN4B8f69NnYE0OBNsXeG49kCHY2TBbbCwwjP9f8fLoV25qqnrxrVHG+owKkY7t
1aJjE/WkulLFfQxuNjBynmkydcbk8jqQZrmtNYQF6c6guVEWRp+hruB0sNhXshsw
/+WUbyLLblnw32UUmKH1GR3wgVPffMdagYBtDtYnARY/XD7edaGfvj2HkZJN4i0x
HzWK91p7vetAuLr3lDQFwhfPUWWvDkbhfjaKP/g3VBSjOHpqJBiG5pgy6eBARlTR
vR2NMMMFYm0LWg6gyiplExIBOmXjWN9ZebmVg1rWN71zaVXjhc+SLmzg9ZPSkDl2
`protect END_PROTECTED
