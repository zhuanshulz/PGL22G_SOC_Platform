`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cT2gvLUBdRFwn30BzcmPFtMd/Jm/W0M6NsU2NSYhLbxI5DyMjPFj4Cd3NdUS+gTf
0vols7ATwbcoTP8XTDdgj3kiD5OlpWbgAcpL1H6k7ZTtGqLNrngM7vF55JDRC4R9
++Z4b9PqH3a6o2UP5fkrseu9yDfPNCKtvCKKjxWX9z/iDNd24N/SZrLL1pClBnDN
28VG9KKzf2riukE6f8aashhYtGeEjXODmn5Sd1lfYah7nqMojgOavIODvYWE2ezI
LC8erzCnNLsWFgCtY3pMYzyR13N6LngmYWVMQvvTrNjJoev/dblaG5Fj5y2ukC0b
MF94GjIxb8s0QrnagZdHY4spZPoNC8z0jM/st0ySm0uwXWkmjWQFbEfFkQice4dF
PoCAqWtcpTqPU8mzqsjgmn3swkgZDNBIXOtNkqzi4AOIvLwdRwVSuDttu/d7RPj0
EWAo97cWqqhd4tJzA+JgvyXMQAWgy6HykUYKahwtZruWebOReKyEMhPpAlbO0VwU
aTzXDqZ5YcmQ8wJK9get/HsOd8d3GeXUF6CMufTPKjdakvMNcyIVi202XELNJPih
TUEbJmduwZ1uBVmWaAYX871iqkiXL8kLMkqYtfxfbi+EB1Z3FbGqSUECV67JNNJ+
bg6ddNfBOBBs1GEnrW8AFXsl4fQYXzF+VcPY93I1ROzvkl/uxtqbXiCYLPCkk51t
nEYU8ILwcUg643OtrhDIgwYJjaisFudPuASTXvEpwGSRGzokwf4KG7RHRNyRl9Sk
aYTGcto1fv3kOgAKcnwk8PsYA/8IDuADS7tY2lcixXPzm5/BYCCCRiDsGgBBDP5M
YCUUW7d3wiaWuiRLfO8Wv8hceHot0NXknmkYZFhMuh/lGO/A0LfDyveufiUBDTBk
lSHrTRdQa3w7lalULPlIzjMuz0DwcsERfTwgZZZfUmG13jGq9DVOyQfXyC9qsd9K
Bty9dPU6cIT+OgXvY+IRVSP+vyd5jXtg+EwcnJ5DCWc3QL0JJ4gYiWSXHZjGZPs6
KQ0EQUaGzTmm0+6vxkN3qi/Ou3nW2wlM4Hrz32jH82maqdWsrKPhP1jhONS8hOc6
LS27bXvsAMUB7D2xlhsx1xdTqVLwgtzln1gLFT7gUMgkq2rcj8JPYk9pPDoxEt22
bmTBX7pEsYteGg8/w8Wn04gcfHcUFuzoysjEA7032qXGiZiUHPFmwR0hikVo184N
8DEpd1zoWCOueW0ZqiZADrAnweuIt84B4UmwQ7O7pcFIj6fBhtivxZCKUHLZE96D
wSmblBV7LZFliSnbexnJFxHz0m6rkFdNqnDEJQK8WNA98QXymnmp8mkU/5kWS34L
JtI03hdaGA9Z1uXyZYh1/A==
`protect END_PROTECTED
