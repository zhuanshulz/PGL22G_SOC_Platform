`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MYa+M9Frb2lv0ipgQpgpava8Uy7F6qqPJf/YKB9xAKu5jZKhMdEdyDHjkrUHa3JS
A8DN2naXe485euxEqDPHfhPFVENCZ+4QZvsdz/twZyTUstBJqKarLtHzOu9zlfrE
926tC47LGAjEAut36Ucy1s5BqJ8jDddG7PdFECJwAqjjWlltWDdUVYRSP/xWsELk
5ZIAYy5iK4XnTxNbzQ6ILyScxHuYN4OY+pQYdR6jlqaI3JbIN9IgYXtShw5eh7Dp
oTgqi9HVwm5+8tRG0/us7Yun2yVpXWar+DmfpuDKbTt9qBu+U0vkHlTZpu2RgRng
cR6bD5lGnAK/FrmKKMMkefvvb1gI5ac3J+DCr/UUvT41UIb3aA/OzVDymyP6WH0U
cH/YkgeqS4Q2GdeZsE44L380P7WUUdF46iADezlEeLtIBk6FcI0IG/o0K/GH0P/r
zPENv63OR4oetc/2SUwt+3ce9hptfTc+UoAK3yyfEOP3NCI0WoR4cd31LqaArsyL
CGeOUxvi8M7D+hmbQxg0qe3Awlrv7lgkGOFmdLkLGhivdo36MZaPYV+buBPPvwNM
huDO8snDBrM6ydzKHLfrt2A2quJAKQPMp7xAaHduZ5OB4ewwc0LZil+7FLK1MafK
8o7cJ6ErMBFcNSINB0BHGCrVwwlmk/Uw+Y+lVtfO38jf/nNPOnt4R5i74GvfRuCR
oEPTsbqgzj3HxNeYX0eAJy97+mBRO+J4lSwT6G6AHBs=
`protect END_PROTECTED
