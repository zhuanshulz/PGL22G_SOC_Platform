`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xW/abzXaRw5n1s43AurNPRyIyhpToPFCjhr9hTj67Ve6Pnv+agGtR4o4Jg2406Kc
UGJ0EWpJsL/pJAn3RXNLgCsbZatdL0CwPQBh3IlPEhqwf36bY3fAYVOkCGv9yoKS
EshqIr/K9NZN13XfaCHZFy4QmHqSCqYnPvLQQPPYXtoVrpuoo4xzK1thUzMBUKor
RNxJmzaHDdrFUuiZ9miEycM/mDw19cbs651frP3qSZFWAmyeqxOl9TyYHTrhaiM7
2w1d84FEMKnp/uzMXMsO690GDi0M7Ex6pMKlGJEYc5wBMjaOeCbPd1RiEQ271tmI
FkgW12LHZjlZ80Tytbm69p3iFy3QY8VXGESUhb0kHs2Rk6Qmo3IB6qAzqj6EsETz
+8letf6S8RAR0au7/P4RvEaEDVIMNR7KNpMUzNZFw4n713adWnjEIRBecXcNWvQa
+vcUZL1t9aGOvEPuxwVYlcdsC9rvtT43d5iI5ucIJhf2+bEuelj5igmBvj8mK3lM
iGTqQ6Bxc6ADbQrlMxiogCaLd3FDaVYYfm+CzeDpH2PdFv2aEieoStTBw9+dKhFa
zC3S8ePe7/BFfGSy5fEZFy4nz8QlyZfwFiRWCr1zvBkYEjQAdguP2mF0f5wcwnCn
rEqvuhcWY6cNRVWwr75wp7VO0AQwpXQQNFZQd4XRJBEIZhBD3taeJF5NZ13jcpij
RHO+zQfhVKDzYoxGVw6jnT2k+he4WY0tBFcJlFs7AYA=
`protect END_PROTECTED
