`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zVjiiwpUh65F8yiydFEYpbJHS9rbB2rJw+CmS1DaNG904Y9R/XOyGmaTENxm1Sx6
SBvXnZ7OeD94TFXpmFmzCiRcKemyR/SM7dcVI7KOc+3MPr9svXCHJOF2qoWsmrVF
y6JOCBAtE4tkJtfJEBiKXFKDMiuE9RlOnN8Moevh2ny9P4Nd5cwfB4z4c5Sb4KGG
MAoO6oLUI6/sDpAC33agGfJByhgq3X1CPKefkZ+C/6gbx+xwN++YmMYs/XS/MQL3
oOK9osGWp6qDEsXl0/d+mePgUMYEEdY3n0mfHDEpElY7qXr96Dpkb7Gn0WWbhf0+
uz3HC/lZwZYUaY1e8XGeEGeRQXt1dlN2Ggq7cDayKtXXFqPqZOpODQ++A+vEYe88
IOWe3QFCGPKoqJVa5NH5ePrQIKwVRWRXq2JpPZjM4ipucW4dt1vdeDrODe97i/zR
0Y9FDXv53Xp+Psa1TDOIxHghqCOkozheJWg9sqTQYEtRcrZblXhRqtUwLBysCKGN
RC2mm0MWIw6qt6BK3r2NZeW2ArS7mXbFyHerM2eXCxf4QaoK7u7Bi/IaGlmpAOeL
WYhVMsDrANYm6GxMxsfZDzgWchZttgH+YE04riA764D5YGOYFtJv/xJGDvJtElYg
MvSIyzwMetp+/yIxY+rS36M9YkLlXqqmiD9CMxHM6sLp1acZzzreEHZsyL+3dpqk
8n2QkkRIWMxUTNDOWmmgC94vjKUh/BeatXZSz8K6f+kG0QAwQUsaYEMC6EwNm7SY
zBgwN5wPeuYyUgtamtIqhYO9Yu5B4B14B9CCwxFZKxSG0GAM0WOakw3cOSkiSgYB
HdMIyeEECoqMf7S1vwJEYKDhL/sMp5rV55r3lql1F81HmIkb+loW4vKdZlev1gi0
PdHEZ1iqs5F0MO4nWClvx73UCp53LoMwBZOwRGfHDu19xPUNytz5X0uwRBtcPfFw
HrZEU+gq8m0fOtZDX3OKt13w+m/4khbGP5AvjVD01yldW8q+Ktl2OPFxZvPmCnan
75hM6ZrqmF5G7wwlHRV8dg5bDTXOTUwCJaaeGIPmKPk2qWNtYWsWkkgqsuHvffkT
QwF0eitzS/M5BZRxk/HZJakGhaKnlYzt8BoTWVBvK+V7Sn9b5qTWDIQpF2kBkGuv
WTdrUhIypAuE7fzvnwrH+LcP9trg2NycRv8diAFdYe0OE2Fl9po4QicWNjUQfjte
bXttpDSpLrny9ePsborATuUuxXvQhDxBWXbZbX2D4HZ9apEaZNk+WIiZFpeMKcEd
dP3Lp6Qlebl7mUhs3lVBXfmfOm1Aho4A/aGQxOWslYq28TlQ1sd6ouzSaFh0ANEZ
uqfbvEjXYpovYT06kSADlGFzQDKBA06YBgO/ftu12rYE6uKZZtc1CiVygljLP6JX
af/ECb3S/HoSTIZjY5Nb+ORSmAEJOeWS8kPILOgCWgbpMarwE4/H4ePEBGC9YDP7
RTEyZpCRpfDA8xJB8zFOc2nm9uVyTlLCECyKCb9cZBuLJzvHkXzcGRqhKA9zrPoN
kS+hsiLgU7GlxvFZ+omYkVDid3EfIj5ciUNQMfC0A+rXz7ByOfGkgS4AhL9kXYUg
o3mFg2e0kNYLRhzHl3U3zlFkvDDyVMfb5GYeC7vksgMt4y3fbfzdlysfY9E8jF6Y
V1Qc5/Zd3K2rDPRZWUBHiWo0voupEjJ40lbvwDPAWOQl4mhyMYUMz1N3/Jlzr9cw
a/Yv3jxKWKoVRkw20NBwo3e5mCGTOj69UmAxKtPYdhdxQaOT+paga/Oa1jTFubFK
oqHdzJjHXGvpOOQZe2CizFKRLW2HWoCVXrLVvDgbtP02cTUFEILa9yvco0FGFVZD
U4Nf8HguD6mcywhdUSmtGhEJjU5y7K2KerL0fqws192nGlYO0qfPBaWavvFlaeCg
Y48VW0ufJMlPB77cY8CVOIH62yQIHpGwNUjPJr0Z4ys628T56H0yCTl/+vGrY5BZ
WzfEhPFWUz2e+YlHfAwGqdq6P8i74refkQRRNJ54qFgSBvEZf2M5YcL6XxZtsQBq
EDlWzzEzh8aqfaVK5Tpw5xTnDo1nALwG8DnT4Zpe2npz6D2g+C5ubykNkr5WW7pj
ESn0GYoWRBV/g97fLZ/BETvCZghh7V4s5kxlWfZ3yltoad2dKDaDmyecff8QZRMx
hOeaePFvlsgUAFquXkxBqyH7emdLh/uup7B85vMlwcE6WUgffkNeP9u3A3EWL4dd
QnKaZQ5Oq8OsJfjjyI9YCnmWFOewnNFEOWydqc5q8/gn1LbkLfgMWG44l8eDsGMM
6Eq4i9LVDNDfUFFdbTT1jX369pf7qtnHaZGc0WL6R7P1ruDsUJI1JpeoH/4azbz8
btSmlzxHusOMmEIUKm1vsvA31jsQnhxfVOL82qDJoKa0PBwkiV9SVHmdyrOc8eKZ
pKqjqjbzkcVxBw9utY2ItJdtwS5OWjQF4R5LFl2CjnC7X2jI9uUTZ8JIZbkuQNUB
a0t0GWLFExS5u0knYUzwLy4nE3EFVMSqcf8iYhPO5h+pt+jNVDE5eTxnxdxBjEuG
W5y+DQ3VG4a/h57wsgk/TtipWOidp9Tu4tXpIkUsdEN2kA/pe6d+j5PXl/FIxWaS
s2+g4gnesktGJksNKcVkHdlZJWgrxH0O87Cm5KJUeEOv6lWu/vhSk0NXlm2t5iDp
BadN1IQhbcyNeo1uD1ipvH7SxlpEP2k8zS8IielpCM/SSlbyVpAAJwRMnkjqgHts
+oHTPItutMnHutUU9vqsrYGGkm5rNI+SXicro9wk5bdSqHQnSSxkBT0zVKHUiJ5a
szKlHkPRyJcC6GHbuMQrKxifbfaMyu165XV9JXi0JmSBNGa8LufO0VgXxPKlvnCN
8wNY4PO03EI2FrL4AMSKkjW3bLsrYAmE18CAGbt/4RWrvkUW9dmlNAUSRjTEyRDH
nc9lieONtl56Gl8us3DIleMSyVbWpnS3BXyKDBZcxIW+W2fbzqMLcq6YckkLpECc
PxUjBSQ/XLMJrMLJup/XmaX9WefG5RcsN71GC49pVNYKPkTOh7OfR2AoUdc66avy
uik47qOv4elvUzxjBPVfi0tj2OVzEHcc0hM5uUl4eHfwgRMEioaExls9aeiQigFS
Rg24Mj0yxc1j1Pw4+GwRbWDyk1Z49KA7l2Z0IVoltJ+nd0WU2G7xqiC3ZcFmStGA
ptU7eZbHmm3Ec3Wyw3HgE7sSXx9fGBMfRtQzLkUpsvWIi8VIm6IyLhZn/oEH9mFI
LJESjwBiZCHrNrh2RqSr0eDtzbsVlb3cxVLqg6xKrHQkPzbM4A2Ec2PHW+RwiY8b
pi89Hy++AL1FgnWchYFVnxiS7ZLxD1HT4nf0Bb0MwzZxoydoSvu2uRQg1cOEKlWL
2TjltPaTgh7swiLii8Xv4NB3JN1p+QaFBMO6o30cQydj+wFPuiVbcTq+InxP/hlH
PQgooQyftrRgqTaypvdsddZMi9AD7ZlpT/JoW4YR0hJuP25Wmj1s0lFMtv3AjAEJ
DSFmTCc4RTPbAfv03AXjRsp//FG1tUGUdlFDmL8B+ntDG6Ip80KAPRBYwH5MobPh
2xau7HzkGB3TdDJ1ukMHOXowN/3xYTL3RjSwZ63+5cCkyuijK2YFjwKu2UEryhcU
O380miu/Q3YHQuS/fM3Kbmh68rGvQ1D8by04gCITVC6rrW88iOAiizBnTGDk1c7Q
mcAt93mrWAgfV6sP6kDn9C1vOp2aPoBTwno+O3jBYqSkYjxrI0C0PYJXPgTT5q/A
mzL1QjqVmP0WegIW4mi4vUgO34Ambsz0/vCMqtg4gu0FqQdT65ADO/TxwgT0k4e0
i3Nk4DEwwhtC5l3z1IuWJBbo6daZ0wmJJH9Nonpnjdq78UJ75hmWBoAv7pJdPEYl
uQGXxcogDbua2gRm9T/Gd8/Wcmn7MTA+/eTp3xNsBOSx4GkKjTaxa0b52gmlC1wj
yjcyOjla+tEPFazFio4MgGh6T12iChjCf1k7QHAat1hHjpSaHWGezYx86clc3qgr
GlEsi5i0f0eq+YxaH2+o4DPeq0U3djAInJqtwZFHX0vQwQgknYunlCFzoZ/wUGHC
ONWKze3cGTbmKEVOA/RlfU9eYHHThSLr1hgZHkFrLbTzbDuJ2VZtK5t+8OLEGAKB
qOOsiAwhtS32aFUllMdprGhSI3iy7n7Gl5g5hi1npRMLu+zZdVWXhoXHa/UTNE98
71aT1EORVFsX/+H8UxBBDU2sanwJQs9om7ZSC+wXTLYS1nNdFUXvFn18nb+Codyg
Df8U7CfE+ayWRSYN+gMZmQDSeGg66ReQYVcxW5BZj9gwnoOp1blpGSzwgNhqoGRu
MNWZAL5PRgl7LcC9Tn8vGGA20YffO78PUBmUJJ3qVs5sCY7zSNeuP8wqY0Rtl1ml
8sYJfZ75SYVO8p9ifFXZDBvSD/L5coyCGKEIpqCKwlUL0xHSAXhLZrADEs3aMKXn
LWi2sSsx62OE7L5rwUPQ5msuvZUrMdVzM5GnWEfssnGK32QgAeS6waZwWLXF2d+j
5ZsmflCG8p4NurERl0qrZJNvqO2T6XLxt+jT+gr2p/mniJQ8omaHyMsNPHmJuSNa
wGomp04/jyS5RqKSvKkXcsvhNcdWSNzA2OWQ9VgKqNo8sTa9RtbBCHBinGSorHCh
YopiqOyt0lv5LiogyyTy7CZl6XNz3AOJQl6IcM7KFL3Pz6le/K680WkMWbVvqphE
6tSr44NutqZh76pWkb5N1WagBIJ2finR6ShHspgZzV4VhVwGWPrm6XKo2G/2uYEI
1nrJtU6I2/oeGvVCwVs6gy0mISXTc71xfBjPtiC7Zrkw4Dm3sMVC55QcOqsnKeI0
JBpkowhcB0oRrU2xmdp1HA8MXJx2LipWpBIryLuJKb5jq2OXnsKTgmfLR/pO1v9q
beCgA1WsPaYKHaPeyiebsPGCVR6p45mWHbGD5f/d131d+JUtwtV7iHv3f0q1+xf2
DMr4I8yHiNxO0UOf4Bi9nXC2hJ908VMA9KuFqZDoF4mCwsadxSvQhfLufb4x9s4a
C77E2Cp8+etsvkrI3jW7Ug==
`protect END_PROTECTED
