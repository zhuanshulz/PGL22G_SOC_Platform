`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Po6qlg0F3pYH2PpHhac3VYf0P8fdni2Tp3Ng1uPhV8aA8X4mnjuUSJZbExs5buRy
OSdH67e8p0o9yD/tWkNzVvXyX1RdecYJYHPzR1WANWmXWwoCcBjSuEYWZ5JHAoBp
ejygErlxFt4w+9N3ANqoFW3e0ihfkUwH+NlRnR5wC7EcOkxfcv6nGx5dL6QLn38J
RjNricXZccpfvPg3RjJuwUMq4p+zgQ7LyI9lTD0R/g5Zh2dzlf3dhNZO64khasBK
iCH4MAqX8jADoHxs4RbOnW8XStr3NDGwCwCoNuanXS4ZXDshU5MgxBFvne3GetsD
deC0BYWljHs6hc94EnYU3KQYB9hYsNrjEwLXUfb5oFSYQ0P16ccEY+3uUACwvJ4M
HjI6zPlYsWxB9AN/5oUaBg==
`protect END_PROTECTED
