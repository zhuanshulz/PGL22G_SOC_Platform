`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TGVaN74NnMYAttja+KwbG+FFcuaE/nTw6dnPTI+69CbUXv+vBsvdqgB8dSkkju+t
cZgLh2NnSOeuQ8PVRmDieqbzaDxJTVKHXvVR5kQlnfOg7xnmnMjw4zjv50eo/g4+
cAdiDJhoUYORM5tbblsDwFEmi/KG01EGk9rY0/xTd/X8+b+k80jmxFhaPKzyEJJv
0RtM4Da7cMyaroCWJNH3vosgVZDS1xhHqwk2ekfUb+7QbtZYozdzDz41NUCKHGIb
J9JuB8xZaYUYIDl8dMczb4KoswF88sErE/WvriXgN5MoaHunCaXPWkrof3FSUj3D
GiOJnBrDLGHO6321FQn4SYeGguoDee3bbl3eYmJXyv14ZMsXyO65aSp8dHY3+te7
KcvGnkvzpTZSHPyoVebJ0OPzgKFxEOj4uMdpZBgsahDgCcQZgteFmH2qdjXdfGfr
vgP7ISzx5TIZW+/Q8nsOeuA2OVVYBmnbYHZJwTxrH3O2GfJk+dgGVfO0Ee6eW1sl
Y1gxVdA+tDqwZIobXCrBdV0McYR8rSgc+UV0SC7ClyHVhGo3PiPE5kVf393Cqz1A
ixqPW6mTtYv2RJaP7VmL8N9NHvCAZXWLBoqxyrYgYWpGnh+XTeaCrYO8YXuZSdU5
OdGZiT/IXa9bMXojL3KxSP0PqhEEanCh4YL4vIh5jzsuoDz1CV9hIQ+aCwcOjntc
TEl+Z7OsTu+shAy/YLXlFTOwen8qs0uOzdUG/ySXczSgwXScqFTAM6SOyqY0OVds
Le4qxEf/wwRXO64ty9A5suSKtgnNQlGwx0hc02xFhwRGtH7sEBlVLxIUC5f9dSTP
pLS7RflKEHGxIfb96uUPN/Tl7JqwsoEt0AIbBlx4buqiY7GKK+Qz6nJQcgwdnfw1
cVIQ4o6dsNIoNeCByvnqi2DDhhXCxV9Y8pyVeozknLp1H9jYs7r02dN/2+I33BPS
2BzxesAZj+OIfPnpKKpExhIb/Ze++TBUpN3egy3zT3TPzt+EK1ZdUoT5lmKFJj7a
fc9WzcUkuuOs2G055pVtVx32QfecQKzXq5D9uTdmU6LOAzyW7o1CYzgd34XG3Ufu
WjxJvfbTuc0ko8RDudwnIAuiCbxL4iMrT52usjpQRP0gfVBVgFplfz8OyC62X17G
SjumFaKFzDmOeDvZFw4+gvVO0JyttpMFGkZ7QrQSWTJjWOZ3VqlSeTcc4rGEgQWY
mfu3e2KXefW5aueAKWitd1rb+lCDuqReRyLGE5/5UcZpNGpktguzqeXsAICe2uED
6l/cj+UxaELAc5j+PE/OZqe/PwQ5swk/lfpIk4oEDef85lb4zhFQBAiHP2d3QF8u
/INp2rOM/CYEBaGhgK+lJQ8oN0tGmXDoXIeBzayZv4gQ0ZD1aRxoXvgEGO8Ab+bN
w+bqyhxZCmxw62ptoehH9KwKb3+hAk+stoSTyZtS7/V8wZ2nnXDpOdrqfaVFYuPi
mwhs6s7ShEbZ6SKlMFxZEUL52m23fsiqLKGKIbKKAGBivNZI8LwXaJ+nPbZhNi6x
+ek6PfU/NuJbMFInL4tEOOCaVPp6I2GKq7QVrjqdv/ledLm5U+V5+7gnA5ry7DfY
bBSp+IvdKFsdLJIr2qsUXUvN86RApLgru5I7ReLegHmeriuAvWLqbqdqyVah0OqB
BY6nQ39oTnrtUPp/2lnTzTW0wMI+WVT8Thac/nfihLXFiJPr/XKk9J7BUKz4RjMH
4kL0PY03I1OzcGNvTQqCfw5bjYZ2OC+QAC+5cExc8T2UElZnZ2T9OQHhKkaIaMTd
1bGvg9vMdWCZWKVwggL5ZytkTZ0M8Th4c+S++zGlinrWNUrOk4g2w4H41VYc3bk3
uiVXlL7jn5yhhNtue4tmISwHdwnzuJofxHcj4MttktXjH3O21cLkmHtZcG2SLaPF
s5/cDpf8A1Cx0VY5TSO5EuTghyyySVUEeX3q7ODeqLlK98iiEaL71ApJshDggxk9
Bt0I9bNJDQeA4MVyel0Svny4fozVGy8OFP5EB/AOYmb7J7pH7gwCavu86Gim2PM9
`protect END_PROTECTED
