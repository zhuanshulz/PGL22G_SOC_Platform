`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BHqlWFjVQ0AMU6kCCdwzDH0LYI0hEf3T/Yl67Xy5hkXfC3JGOuwaaj1MGluoswt/
BKQqCI+iK+sflocNxV3zMamsOFm9dlBEce8y1VrLouE070ADU69MeYb6rK5ERs4N
MmkGoOuoB0obT/mUB1Bnz2XhVS3wf9ExoDLIqTz210H3Y40dOaOuUFvrcfpZJv5K
oKNwHmn7grViJM/SW53ffE15WITsEU0NX3g8WnpsHMFL5Cc2QxYcV1jgyRX0ON0r
rKZbvNIZdxMsLDCyXnleM4BYJUrbUTZ5B7BROqwtcX7+kIIQ4rSA3UIFzu+cYsAs
hMW8FrMcPx7I+vihDjqVPZV9OXB/hmHmlRIaGIrU7+3Mw8i4kAXxAGXRZ2shxvmP
7chgmafFzTpql3F4lJnf9DdJR+vpiQEFOpWjRiNPWl2tetbwIyes7ljM7IBT8hWj
6F1cISEqH2h1dULEtShYsBhyYO0ATspCDLcmW0uIXluBDHETsE1fJRihWjXub9rr
DXf8bpdDucq9ubiu1QgPuatNqiYXWbQxnVAkDxbaJk/De9bJUPFSBvEkqKA2NSak
cz6zp3M1loNE5m68gZTWmv9Fmqunkkn7mNN8BnIFxawNS6dbKMUfXfU423KTsaPL
rmkAT78F7iRGmgDBQ6oE/c5+wGncCqqr1x4PXJBGyT+0FQcA1NUjnW0seWgqOWlT
lu9Wz0w1CoX4gSoXBIorERApQ6MINS9MgF9DFJ3id74reogZCWLPXsmfKcD15hYu
jrcUx9HhS/kjnjrJSLkjBujknb4sUxpcp6QllJYtSahyQOx7sLLXu9pANaWTUzso
NsZDW95RQfpQU70MbFl/j416DfX3qDjiEFtZnVn7TW8teSlorv4FYN3x28G3LdJA
0YviQxlcCOLJKeOUAXm52+9+QAHyBx2zTrBRpkGumU343IOwmVFWqtmPhYZ1er0S
d90r2Xd+yIinSEgoDDUTUbLYvpeeKBDWz2cT7hIfCd/vbF7WCzm0QJtaiqMgLKZI
/AUNy/FZhitDVWQuoTquelCixN0nZFMhSD5Vy/aAZrO+6SQ9SaqL8RkGo7U/1hu2
WWBe3Dq/kiGP34K4PXFYSSfVvcx0G0mH+nqRVaFj1st5gu/NaHpylXgBlxrVEN8B
tMWV5Uw3rZoNSeok4RaKLapTHsi9NvhahE6daMD24IqO9/hutRvsmt6PyZJjgV5o
5TEWh+xtQ7qx7WKxunxRbpSBFQOOsOHr8iV/mIAUk7Smj81Pj8qQnnIH4bqhku39
GBuoTutkwZ6F7lbEyZuoT+a0aVbmk0Xzs/c47fnLPIcHuAyzPFepO29yiral82dY
L239mVn2TULAYWmrJYEPJgAZ5c4fgZJwM5KwcuowsX6C8FBE7HWl/CC9LCQ68cVv
wntBCX+rXDLIIwXm4T4nwaPnGTFne+QlTg6+4DvQ7WdFUx4Px8y43VPRztomYlIr
hlS8+l6GET/nJGT4MTpqtvvHPq2TJ6TFTIGyTy4Cjqr5of4tZM4wWQssl/hlrRCQ
q+HzIQnDmfvqmV44m/x+EqXFTL9sIO+zwzdgBupwz6yDXdXKM02+jxSmWqN7uauG
YuqkfxQIYJB3gz2jQmgHEvvYl6NxzcVK0L8V0RmjvmfIfD0pFFl8v0UDNyIuS3hb
jnbWplPQ2n1iuU/RrsOpg++/06cpdsAlaoBPzV4nuLnaUQreZuQctfCf21mW7wNT
FF2SeqNceSWfk6TDnCjzGCZQk1iIO9qOuo0YfdcbcKFTAUV1GAzKhWalt7meAasS
XyjokFrLNmCTbjn9vA/iDeYP3qtO3SnWjN9c/C+UP0x+0XNYps2mjWDMZsvjHDiY
QXNb3RRe9PLvKWTLWIcxp7WY+A+pQNfq7xNlIQl127WsCIPYxB8zuEWKYJkejt6e
VKTxfjT863DeT3W5r/MaercW1cDi0RJcSpPkMKNDm+CK8dtgnrchbyrhVtQ8q7BN
knYTLYC0LcN0sW8TCO4kfXGG+ZswN1OsxhOdmtylxL2SQEVMReUEe61OEXX8dP7s
utRl0S6QAOyJgWNrN9cf5a5SuQge5obypD0Sc3xo5nzK1lrmQWOijqvylFEVKthT
Aw+MqpaGLrER/cMjlulPFlZqky9gWx6rUC2h+teavXDNJlHoiixq8JVrOvF1soMl
d2Uaz0/RTwqOJP/v70ylQQ==
`protect END_PROTECTED
