`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hha0znCS3uwmhT0w0E0rJzW3LlTuJfSIQb3SsIY/s8VNSkG4X83Si9Xa5jbNQEjh
cJ6taXP4r0Gcqprw+BvtDz8HkOJwpaSu5W7kC+65BJwUzic6o+F1varhwFqpB5N4
XiOHbxbBlwQfxfakPdhvo7C5hhJkMbpgsJyVA/pLIedBUG9YvR6NmIBcSOxI4OSr
txV6BXVoOkXfqBtPCG7hTBaQG9pUoLbqBnvXhBmrDQRn/axLo83mq25J5ah6ByXK
peOegQLYF6pGTfefcX58Alj+ZdrmIkXkrSSU6m5wbeoR3DVJO7vx+OBET30Y81iU
2BXQFbWMszkXr+dFyOSLQSLp3alTyxTV+1gVnA6nvdEvT8rjqufRww77LoMKuSbo
rUBraN9nP4++M9GLPMSA4JLtYxPTt0WZatCIsPsyaUY8hZSRcTpt+lR61qDBVPlg
p5Fr+E6WnVE8tknhapddenKYJ6NTpVfjncK9vjbx2kIxcVdj80HFhOT1+V2Op08F
WFLLc2si/yTqhhmUlBIBp6fK1mthqOZGXrbhbjk/h3J4l6nkmk4qK981PXGq3s64
OmM+OCtNOOQ89MWHwZcJ8YBKjMenIiBYBHBDhM6SJFNwAOZv5ZyAP2oJkIOb4m0u
t6tcFvcs6qEUXAIWEdbuIfwVw8FU8JRXQ5bMp2cdRfeC4rdbYrlusHcyux81+EB4
O4WLJHR0ShF07dpRPRZsMOQnCCkm+09BdV31gTm5JVJjezHwskfmgsXjA1QAZXpD
2m4Ult30z79SyMbUQljN9jlM2A2h/zk0BlZuVenK3B03ZpizuKMbYTA9zSCPkwX0
6OuFlpSN9BOSgtQQHK4Gg/aLkwY2Neab7PfPdnHcB2naWEud2W+AVzrs71405FUG
rO3B0KofKz6kNW3Ue5s43thJUUX5a5qPni57fi+3h7Cnn8rcFfikm49ni/os3tVI
LTJQXX2fVqU1cBJbsRkAGf+TJbuQNW5TsE/Xhbak9J+VZXxYFALAV4xWB9bCkJZR
Nvn46I7ke6duJI5th/MszC8+p39trdm+BjQHkKKm50DKFYjp+0PnIx+L4OyzSSCl
B6ezqaGvVpnWe0DolxmA8x+UwW4p3NXDYWkHoNI3zYr0YQvN7Xjp1+EH+XGop9KV
LCq1SEA7mXiHGfsQI/YPuR24033FWEqDl/CxRdU1COmySrkP0/I7R4w0Nw3lwobJ
Xq+9f0GVQy3fr6GxOx5Tz6QCtZUtgfdJEFSMJnHa5vspPWSwIiPfB/ktLww6WIwg
Av88Hn7r+DW92V2B4KSIVA==
`protect END_PROTECTED
