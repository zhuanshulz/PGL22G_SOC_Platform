`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8hsJ2Guwz7LHHNr6h3PmXEVv04OqAoqmJnphhtrORFSeLXWUVHEKeAj6WnDpri34
xdCt40/U8YBD2LkRD9bsz7sM2j8hSXwbgM0J8c6ZK/JoPNHI9BSKULrGAgvmSocz
usFiKhkVpX/pDj+eaGcsgLm4KGr/xopGb6R/C5nkEex1PANfzbzkIWEHNcu5Aaly
elsx5oJEiQx+kLxBxOBYu2dT47xjfe7a6j6rapur+9tYsi93jWUQ8xrsoAQVmGoh
j1IfZos9hqLDYNybdfJV6w+KMQlDZVe1KW3+aVBA2SbXEuQm/fFkCNSGPu+wSL+K
e0fOd02LrzoRJxc8s9Yu8xDMq8O+PC5VFEGdv3f3ITH6hbytEy9ZeVoywxzgcPoF
hmjlcr9zciY9ZlV+lllUNodhwPE+ONgd/XGWZXMHEqMGju7d+L8Up6NrPrdCyS7a
6ftBhYOX1f+xVfnA5g2KWE8gtC+8zq7YYIlrdDY3jbVF+0f3XocIhXyGoN00Mqu8
/4ou7jjddtSsj9sWmE7BEFg+QDeHKN+3kTxOfkiLQWEVdCu0c3AJO1a11oDJTO3J
p8SCwnzyJBofguggEZO3kNt4OKsUFAToyQIqHEeUQDGx4w/xI2PPFI3oN+S5c7EF
+J7rMKGZ5dWzACslH+YL7zl7MI2ZnFexD11OCCEF2uoNPoZm/YS941G1+Jajly+R
OtXWTf7WJ4WCNvn+oL9n/4XW9I7Yal+4+mOaXg+IxpudWKvG2qK2MTdALQVPd7XE
h6fnaabni01aDbXE8t5gRZwYC7WH7Oc9qXCRik/+evYTyM/FBPW1PjzVqFHW44dk
`protect END_PROTECTED
