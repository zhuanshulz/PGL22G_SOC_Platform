`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nOUgwguotK6GRJoElNhfusfmANCd0wmVJFvA7ZrS0FrZEBp2IcilqlziaBJc4IMr
rBVe2NOOAD9R60zHkDGaxdK9dhCWhT5Ds+8GpVcToOujBGZd8LmJW3vAsnkedIVL
3RnM3NupNZZmv6mEpbBRR6qtcjXkmfIHFsorXkp1xPoDuIllpXtdx5WmxXNRojDA
enH/TOD1mSsxpFlNrVAXp7ATDudSGM6VqZ+7KHaH1EFE5axqc0UKnpEXUKhWq6r4
fxo0mM9bM85zOovrrtW0zQDXQ9F1J0hXQrbnWRSfeZeZhoMdE9sv4elDo3n7+eaE
sj89xODMy20o0ZQwmr3UE4wxGaMU91ZjQYz98Hqg4lr2URPhd2irNaOWHn318mMY
5VpXexAhbehqLt/SZuzOzRKXuOdEmmvKwtLXg6EpmJegrS1fwdRfTJv+S5hvBL38
NJH3obFxeERJAfMMJmfq/22HuVUQZ+iI9y9AjAJT64gvz6pQPmE5SiK8cnwSOArI
YjPXbzdWy62GnkwOyLr5ZoHuZCgYeJLbBZrI5b3/qb6YnfLXpgq/K8PlMDQN0cOb
EyPzA2wztkbBrHzanEdAOLclYSP6xp3GmY8a++DsAu4YQGNzp0rCUFrdwjq+hn53
J95uSvSwp7YsD/j/Ry5Nx3R0kTJEvvIIMOn77Ea/UsoNqGBC0pakc511mv1q3WGt
lgYBS1Jbpe9Hy6OuPA4s0ynHpkuSrv7Ol5Z2QDI0wkDfYBlQy5SS0YY/GfyD3/OD
ILIAiuAAwew5cL6S41rQnDqa2D6DpYmigl7/zDWJQkvnvIl2VaDvorE5ZPh9ZH+d
Scs5pzIGiXUtIvRK1kS7bUl5SoZBxcfaruzF+2EwHOMG1aed+MeCH96oGtd+Lq+6
AUheWY2DIG/pq4N9MsUOQcDt3T7pze243/LKwr74WOvTEcYWNpivyHPpWqQv8Uu5
gLfd6wQ50PmR2UryclJMveHGfHdwgsI77EzkMIvtJJnxtamNGdshL//SXS+i3GIB
JH47BSxOU8H7YUCejLCRAesBIlD/vB3hFjsSnv+bK+BFi+4nk0gH6/ZjqqU9uPQz
vbYToE5/HNrpKIMZxg+44ZN0O6qzRAVpYxzLp75VH+w=
`protect END_PROTECTED
