`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F+5qZaZW1RWki3duoJhBR+In+9tfBMg6enfyTF+OX3GzmdaG0PAaaRptBX9DuASf
csFKLj2x/p5CCNc6cZ9RtAdn3EsgWJTVlUsWzmttRiWVtiekQdKYoD4/wucKsaaJ
O5D0mVJwzdo7FPAKcZthgjWvX0lKBJsUH434BY8u1MPlErIy78ouJGHvTrBmKdu2
mLn9DWs6GemTGhQHlyu1TKXI8+DcWK7xlGk4lyCRmuMPuo2a0DLdewXhu64pLQS4
XHFE+pIin7dtZo6N0z/zN6AeAv8tmtHKRondQbes7+oFHsuGuSf8oX2WGaOzn41y
nlUdbYemsX9eqoVEiPETeQCK0i3o/9ssNEl8YQpZxuVLrqhbBBUe1JnmafuHcyTX
iiRU4dBWZ612Hvo4Vu831XtNK+7azyttT8U15Xpmg9/Ea+qyKSORXnkOaqYBmVt/
LU22+T1xzDlboTkZwcgj1EpQPSJOOLKzvy2XObiZJMcELNt8nPoLo7/pjxUYQh8v
hBE6ksg6KoJ7MCxsV3jzzyyqyiNNRNUc6odPY0VE7mSmZWDr9/85sF+30HeJqIvF
7oolMeu2B4ADimqak2FIDi6Hjk18RNedqXmLXN6L1I9eHi8MFtdKzKc5vzr8zKza
kMZTlIS/3NC+L8uEntSEqseJ/nLxO42MA6X9ab9GqbZ8vNb+8UNy6DSDiwbh5UOB
OLuOtEFqmnpxCo07g1NbN041wF16PLRKR0ojxX0OEN/7p520G7ErNirRHYxPe6wf
NPdGv52spIqz7SaGxikAQHMWdd4JxRBRki8hOunzcR1T0lQSzOOej6Rer78pM3cH
58zF3U0Sgura4MaI+/3/wHc+wBOvfZnq3a9fjB56FSQ=
`protect END_PROTECTED
