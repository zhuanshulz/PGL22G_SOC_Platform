`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4Sslo3bFIJ65Q+P8P1miUcIbAC8sCmEouVqSiAc2dTVqHYZH0HDvS4oAv6HW1yaw
hXjLUcasJ1MpCFpj29yQLzb4P4V/IthfOGv8DAEOKMYmdp2XuJD5EABR0vrqH+0c
SEyJVrlLObFhvq8JbOZ++qr8FkRPRJuiR9+wFmTFUShdnPyoW1DTaCHPZTxP2JlS
eg7c3hotBqmF+wd7lXmnZarFYnvnucMvlqdCx8Y+KC0OlBFTGYGFHrc0zPlRP181
9UxXxvT4X/gZ+E2ITn4+3TsUSgbAzJsU/w6DWJX3ljjbAzk6E27EVg45SncCJS8f
srLww0G2cgsbflFw0Pct6BAU0V1XCygaAQk2H/MlRRqIRomFJvvsPSFdpTK14Sy1
AQmgZQkdg3D357ia3CQ0GCJJsj7lvd6XxL1pCXX1IK9helVmZkfobkowCS8CfG6m
knCO3JTsffUE4OfCnth3jLtHFg0yMKGmaRJtPBxCnC+9L8UMmnlUZkXGWA8JuOkA
zRojOtNWS+H/+b+3tQDn5nPyseg8nWfy1Jf4a4qThJjnbCVDuFrUjylUoBBqhNRR
hYyOaHRJWRyNaOIzR5vtTjjJiNwYcUlS1A5+u9a22deiXnBEm+UNyRrOjDSwJvCD
ObQuIXtJOGp1EudrxGLzF6VpHIY2gGe4yZrENWrNPIsnYrGmAHHtR+VoMBjKc3Qr
BFPTimHz4As4rum5y9L+hJiJsyV6pCGDIMbA579mOJqgRCNNkBAA3pbAYJrSq2dT
tyeayeKZ0fZkUCG/FslxO9L29NZ/I6qHHg013f5POaWkLj2i4emmsf8vginCgres
sWlzZkCdTXLruA88swIDc53kGAMd5X15oehE2lwN7x+1K2/poFs3rweCvjNMZpFz
`protect END_PROTECTED
