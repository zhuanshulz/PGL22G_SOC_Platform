`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1y9MrYkx5+/cyreGB5yW5Lij9NmBdQdvhkSuWfQP5ZJOQlUXxEOvMc+YSmTDx8po
5MYdh9TOjsNb5mSTmtp2xqAZDmLcOsdlS1rwRj/h627XZlRslaP6BVdS+MWmP8DC
nf9T7buDKbxpADBNPoHXOObCUq12A21bm27E4WXUn4gZg5R52iE3bjqiAXuUCBpJ
zpuHIfmRZubkxaAMkkK3ouW3lQ1wRwmiR0vRSQLwYRjB205Dy2awQbvkw3d40C93
REk9QYLIsWZMMPeBrrjzSzjkTOkV4zYoeiF3fSibbMsh4SOjUb2flIpzS44fSGVt
Hv5g9tJeN+IwfPdKzkYtqOu10OP2oOP+PwByUXLPOEK7kj2+TiefVX+m62yKTi7P
9/RapiCxobt0/b9WaECK1NPQbdKgNvOzRkio0+39UyQhuhMq97/iR7Vyd6IekyXM
WTgP1CApOvYHzErbM7pAUn44Cp3O5tTuBXjjYFgPg+mf/grS7HIMPBQDMswlWGDo
RvVQDcg1fDP8xZaRs+n61YDwur42+PjPSShqbWjf0cgrKG4zzsvexSpffNkaAx7O
`protect END_PROTECTED
