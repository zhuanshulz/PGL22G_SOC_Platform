`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EbLhmmNRAJ32vZplUW1ggDaQKaKBpGFHUDIoA/7fGKLIhsiYwWEqucUz1/x+Fbrc
bhNbux8uKxB9Fx98F6bdcJNtHI99injjuzPpCqh8sqY0tuL7dhxgIJ2l0jVFUVBn
kcWVPFfgEGDdt1qUmAMEz1EQMZjpwikgGfmixrBOBlIhwLlEDG/ld+5SqDZJ0Gyu
COdlv4exywWdFaiZJfq7HVVOoa06pCL2j4WG5nBKv9oxcDe0Y08iLcPkjbnymFPM
e3OOUKFgbVUuWLnM1LsOfg9mjhz0KHoeg+uCqi7R+GyqcbOJgfHoKPCp0bn0KgWK
l/GuKaZox1CsDuOgljNe8j9Lx9YsL05F1jdIBLpEo61WGrNH1jP1oIo5XO/FYMH4
FtXUVc2clHSIh3BRaB6v0Q==
`protect END_PROTECTED
