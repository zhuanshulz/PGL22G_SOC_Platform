`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bizCAUrWvSAFr2o4EFnO/zYQh9shwX9DbYMgrmDZtXfFtNSt+bcpdejAhuUq8PeS
2hAj/vkrFF1pRg9eX1qP8UgsJGuapnDbEBzhxUQWmuullgtb1jle3jum1lq5ApOc
aZlKBUzZZ22nEXnf7AnPZw7zA5cROrkFvtzUStFgt+JOr/ssWiv//0vcit90D5nv
CkxvbFLlkquEQMs656YVG8y12eW7O/Vnwxwjeb/9uF5XKczDgavrqEF5jo6i6GtY
iyYLsA0Y+Nllk6t4Ygb3nEz4aUQiWwdWOwWuoX3VbKpG7il8vmTmmLpPtw2EP0B+
uQwJj8yMh3gbq7AHatWDofwYwTCq8dLD2rcyn19/N+jZA0yfCJOdMpDDPYID2cLW
BB4t7iMf0oiaOLAk/Epivmqhj3ZW6+meunPYW7nF05oKC4xSOSqse3TlPHDQKOUS
X0FQ1w/daQ9hM0197rOrUI6GUkM+CFP7HATHo6YWOIalVfg7WYWFEHV1ncM4U0f9
OabfPn4nh5xG6kwWeFE+VvVvPjT7xiDvFOTc4z5dzmIINepuuFh7U6O99/bd8so/
TMzCD7XyGZLm9gNfapr9KWITi1H3aKospZ5YFeLNBY5ss5MnoeSZ4aqmoSfCcSkR
6i2IfR7uUxifCFYPRKbszaw7uOM7bPNSmlXhqarvl3XlFHfU6Xccbhq4pPCrEcE0
WTdF3CK3Q4JKjtMQPSX2HCUCjod+ZL5GZCDfDIECgdeyEPkd+LG+IypxFsGQa465
A6fWzWzroMnmZxxpP/eJopVbhwKHCc+e0B5qesOH6Myi6ALUOUx2wXqE6yzraROW
mvpBwOl1LdjPVIvPIurUajqXiq3GuztAvPAcI4QMOLzzZgzFKpFEBMhHHqiAHo5d
sollRYcAv7YIYTuklUTCqBbD6Upr3AY7fGrQCRIrK8cNDILJ6Y/UXWYJvurVPgUn
YyFzQBFQSnPP7jkQRS2jgDCVZQ0txwLsy8S3DyWTl8LMgMKxx4/YvlzyEkG3iHj/
EBq60Wnl9NqS4MDg3IcI2Q==
`protect END_PROTECTED
