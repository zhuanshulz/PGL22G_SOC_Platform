`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hhMlXOepIaNo0X4EKcP6B/rtiG3W0plifdHZgdkjBHlDL9X5wWIZBSOO8x8lwqM/
+EWZF/1og7YXPDYT1aC6fP27/EJiV+t14HAqJfAi4HVFz851XyHfKSMweBXY+3qP
jhjQ/0AftyAMLMXz6RcW6850OnF1o4T3JSC5nrRImQ2PRWsb10nmXF2IoxM+Ouxz
C/XjveCmA1yVX1mSop6nbfnCytnFXx+Rnkt97cn/D20JzGeJP1DRgF/KkzPK86r5
eI6DoZejIkZDgAczWUTm0GJ9Z5Qur5LDR8Ca8xUXk5cFA50CG8XP/5gqSj69LXGu
lQxZd/mWuwuGbgDWZinFTMXhNtA1l4zegTxbKF72IYFm0qTMbdroTGAY6G77qL3X
Apk5eGziSkD5bkWrcCyG6jrPLJmI4AktL0SZVtmky5cGHpYIibAxhkj+nfIuKA4e
VYbmBwiNDHRW6MSzdAJ6+Q0o8jg+Ak64vxgJqAksclMc11iLg4NDh4V0CK3vWUgP
6bfDp/lQpUId1yj9iLxtd6tdXgKpkEPZr825do9Mph7Ml00tTDLNjMX5lKuRJVOR
JDfTxAZ3mHRMlX8Img3jCuuAGFuuZQ5+7gu9USjCj6sAyMZs9WsX7if9je0Qnn9D
trYy740YogZJJKT5QFGFQaxAG1FWXY9sdnI5kCCHSk0rfzPKdfSi6sWzRlq+CHe/
HpLFdgsE4zZcSvmVZx1UH/6kBVvxL3akvvJVKXFqNiUmAa8QvAOudJq5TkI1kfoO
tEnIk9yLo5poCwJwQli+5IV6WWC2b41w0m3k8rMwledoTXxaRra000hPebLr6TNU
0aa15uXDihe4i/dDhJiq3wxrKgVj4Ho04Bb6WrDs9a31R0KRqJXVyK1O97cFTaaA
VJcvilgZlZAlJKIRn38u1fupbujlBLcuk125KUo4m1l3cRtcd1p/HWjZwrkRsH5c
VU1R32PALWrxOAy5qQV/C04tXPc7Qk8RuLMIUSDiqIXnTxu2pADRjUWFZdb9jk1U
SjNZvowBaKF1ELxzYYyQ03GXA3jTdxHktQV6gr9uphqLDgk4TI/sIZ3ytZQ1Esbr
wPpKaOVR3K5uyGkR/DP8QMB/JtZTOAHWplYgpM1PfLdx3CaAaJ9yZSkTeEGE5m1t
/oTXb+PLmKHK/JTV8DNnCpUuhhKZChI1S6fR+Mt/Q9DrU4+OLR9hgxc1qH08cFCn
nMZ5KQV0wPRt8eARBsHpRmWX8wAz5OYgH9F6hTO0fGZV0SL2GcHEMeFCfREGH02e
z3AQcsIZy4u5znQicgf3UhVDCa5DFa4qZKu/YYsIRvgtcIc6Km2inQB8o4TqlyYm
KNCd9JYMd0P9dkjQ/gumkiiAr22aeLkKRwuFZB9pGaUEH/IBdCb5HWQPE3liss+D
UCRLtttOabGQDx/9sWHUuyE9w6XiJG5agi9x1ovzLs4mHuPp6C0kG1SnaOfELCm6
VwMrSp4RTMOcWmBik0ArOecRtYWONsddGrlU8GUn5j0aprdx2YNyVcprcVu7pDsP
aUJFmTHMeob9eeMBE2kytCKROPMD3XyUwlGJrvRS9R6QMEg5zPS7kphCL4V6uMpr
5hhPM7+X6qFJ4L4EEbV66czS9NJ9bLgEatPLkrQDXeXofwGfmhnaial6KH9rJOtc
RavzoReBgpmoNQmpMPCd+cnaJaK0hVemLEHPVA/H/Z3JMQ8q3QGZwtTVMv52zNVV
9MauJIFRzWpqcXTNsYZo0CRj+A9i7PgXVfcZZTTO0NDnWr2VZBL8WBbgDFeP2t38
l2e78mPnPTUOfNh5LghBHMZz5Bm4xVExhWZxiV+h6OJlzfbLHjwknw/Gk6PYfP2+
j/DaDBqloraGexX7Ey3ARwCtrLhS82wmumFpRvidnfisXH/kdXIejlsieEnbOFK2
fyCfoYO17k7Tivzn+QyqhD5Srdh/SWKAFl9zau7sVCUUIM+J3b7UdOmqqlMBBQYW
Pv7pO1sOf/EzH0JgVanabtTqncUcrWBjsdZtHKuHI8po5oxmEN3KOG3XJsYrzC80
fsrlYXqRKcVVsLe9h7C33XCtdwgIzzYP6t79q0DhvqHeCtCa0tzCPCmy9l/kM08a
IkuzotNFIhp/rw0JiScbZyOUYGK4uo28duqLEX0u00JID8syr24iFMmb8mWvbIaN
6jrMtyVCbVdIdE8XGi6q2SpDuYKPh4NJV6pM37PJ2LSL310WrlIsdIeq7yPIkzaY
BPsDW5oXb0yqstR5zAgYLMcuYFmBQAfpJ7UzrNTOqI+CzForK6bVKFvgKAG+8ZN4
b32J50ypucUT+DI23YKA9ua1EgGH42696Jh2/2h38eutiw4jXBYASygb0OSfBscy
nD9WvzvCfpY45ckkpiCNp21/cfeLtLQ6D2M0SoIxd6gN2F1s8GYUy2r8tun2hiXV
O6txSMZ0PhjCIdzCnqMUehOP1s3uwZfrMPORSwpk4zGPIOVHLL3cfvVzCvcZaiz4
Zl+wsJ2Ds8KNKKTRRsCP21wPexlMVFuD9uKdczDiX6EdsrGIfaxGIrLylA7w3+Rp
khsstenxI0s7r9f2175/3rF+m/n4NyYtg1vq8TaYJwUOog1b9dPyeXVuea+vBC0I
gZKfANIkYXfscSmQM0Flx+N5mJPOIHsYywspwFKekQ0npPVkC7QwXm3kU1k0bCne
N+B595LBYk8cdYNV73HaMSDbz7spvGWQF/cqKc78gymsoZyiph9n20zLuml3zPcL
Mb9hxAvQKHE8RurtIvLigjsU4uGCy1Z0kHoh8f/rYJtgs0wB6iu+RhfpEp7w+/R2
WmzN5aSFg+/OShi9izgFlNhCnmp59HtNlAqofq9woF3+TPzXlGifpMgyCwAvUhhH
k0ceoPu58WsWPWtYk7EXtya37ywJKVqIL3bsJIuwoBKDIRfKqA2MCpK4hZGtiMWS
1y6p9goALhASEnKpqzPZMphUDpsjpxIl8KRLe+xLT46B3jHskV02uXoLvLQDIPAa
3/KYL41chzSxQvYoj2ENwZg3fStfShIHspO5A8hKAG9Wc2fhVZoHrueHeTVH8Y8G
gwlb5UZwV1aKOtSGdvvKWWUclaTqaN0ICGZjMTUX7RoOJBOKJ1/v7k8yrMjiCarZ
gheeE3F5pU8NxiA5OQZQHPu1LSSbhy66Nu439JchzmR1f1iD66dU9MCF3g9Q4Spj
MKJZk1AZQOpc3agjDqvpeQF5FlB6NAwandR+BWc+7gE6GtJgNG+gJFmEZU1YGKeL
1+jQpc2d9TryGLVii50HyE79dWgHYcVAzwISUVZpi0sNZXocLCMIiyNNJtpIWsxD
MPLCdntJUUUW6FVamFDJzoyyaCdjtNZsNaa5FNR+vRfdU7nWI4E0Q7m60/8m+hUk
KiT+ff9IPX0EbI74ya9Epd2GSFy58fbwHyrvmcScGbk2wGnaMv+zqZDZHIDA02Ws
iEW7W3Ezs45/LUoyZ40qldQMqAg6zVHWdo9+Hn9DrH6seYhkx7bIpphAP1p1nTTE
UYHGeLDqjy6inkLPBb3xnslMOreCqvpbqV+JhOyWRBAvfIemOKf5IYe8tNi/8nlI
mjI//NDdYDBKOwDf7NVBPbGbwFTjdo6T3nKRpUPZEI/jOWS4Umrp5Op1tk8WRquT
h4bfl05zylQkaTDq1O1uVLJRU2JzNQlU7yjxRmDIk1MHu6iF7xZ33i6Oz1QnoSvn
uL6OL6EtjYX3GrJM17mLG31st9m/RMEzZBMWMfn4Gu4qPw1eGmpf62kiyFBqC+9Z
48m3Y0oDosViPDmcjsrRM1bdFH/xh8uaEYw81+SZA8qqYqCUH8EqQ/NXJLCNGPZ+
CalBejDWcjf1ycJCRIH4f2cjDAy0nDnpPGsxvAvD41SiDRj59HQZ+OqigCB1xaTd
lLbn2TDbk7FAuwvnMt9yl6Pcq4+REz7phJKnYuzYJM2HVeIencfr6wwhQcGaNCx8
xxET6l0gVDoSCRgxHSifl1/SpgviFptegDIPDbDGPI18f/zJOnSwH6FZvuxPS8Jk
DfU/GLbKSYnsTOVhj/NMzepz6jPomYHVP1ZdwEQUhc4IiCgHz3lecTewRUAW416v
QlLB927F2Zx8M4PsT9oavWbiAowoFqx/9hpkSU0U8tfXd/NOFnRcd2meDDi6HROn
0rzuwWP9oBLxTj5I7qY1QBgrzWj0ZVH1iid3vPEOeCIeifyDNS3mfY9G9+jOPjhp
vXJy1M4khxgL09scan43vP8XsfUBENRHx7w9K8oODFgpo08HF90IO33Qj2j9+dxa
WBjZq7E3MjduhrlmDU1QrdW9IYBkBZBTrfigx27S/CwxHmktLwk4r8GIAiCc2/N3
juIx5Ab4X1YETaYElMosj74TzoBmWOFaSNq6I816evowjnaieskaIXzgsylBNJyd
QfYP6jzew09tG+aOJBHDxxZIeyz+hT+QCjHz210azWVg/bfBJPpZvQ/CPX6x+uLu
hwIypeWyx15yj73GX81sIDnxGkl3T2wgwWibvi3cacczJKO++dokz3nkQ67Sb6w3
UQoYL70DrGUOH4SDIIBPVYnjjlcr3Eei1uh4L0/69XPFvXfQ533dyjySkXjDR+nB
nNXIfuVrLob2ciPdvKuXc84lCng+tn9JfhKn5Wj0ecM2Foc6nEFClY8/URvVah21
VloA7yQcUQfq5O6PVhsyCDUz+4x9uPDWIiodtYRPno5LXC/7U3QBvj7YucoPtja7
snGGBT5zBy84+3RqxMVsXnkpDmTMym5O78+W/3zxNgvkZ8vKtXL6xjzRaG1R7jSc
dcyWVOpLdjSlIP07gldElW4oHQqKWgynY8A3kCwFNemEvo7PAIyp0yE+ojOtAjMm
7/2B39pqvYlPdHpGO9iR52xLCZOZV917jB3MCl7U2b/1JH9Yh1xSIT3eMOdatjvt
lN/vfiHqhBF0lQ2w/KFdBivYW3TOMDk6MzmR1gy3F9aiTBqsJx6VqJP3O7PUVkJO
28RKUsWS/hplQTol/BHhUukLizsTVL0O0UL4dv1J/qdBHo67WrwbMkgl+eL4hlES
04tf2uE02bukBSgd8XXISVL+Vm4nrdqG095fkWxw4TRALPhqEGtmfUMO3NEVvz3/
XSJoXZA4fNrDnENYFwEZJCuM+ScRI/1KlZzOg57dmhN/Eo1bneGXEWXhIoFIiFr2
eS4P5dUy8420oHKLfQB+8selRd5E0OBjNaqNUZON4D462p2hS8TQgCI+nTRojJgd
VX6YHam+LCBwX4RwbBACsapxicTRL9FsOeRyaHhLjo+3rGfnlqB4k5gKvh8dxAH4
UK7DSJYOjxmFe3+Ckc1M5xb23GrkAD9H2LIcyg39gvMNE9ZpNYDRmLjpn1K0J4Yo
v6SKbsb5Uv2rrRAKNW2Jb9dRc10iHu8P1OrnqiObvJHGj3k3UaUTvb1dQ8cbwsAW
FUquqmdltULz23FKm6WQVp8W8CLB8lh9SfOSRtXmRxOK/mMZ46S/I85Ly84bdH1y
zjofTelAgKMELRssxOTfkZRuDf9CHDOqhRKL3INjDRKFTlZ1eD5UmFWJYEj3hqi2
iy4V3k2/0vwy+3ycRZolKjDxo6zghQ4xCRwPsGo/+ODmAXMtqdngN1T5cYNEt3Vh
rvarPa+Iaak8FfRXUO17eyu3W0oAB8S6dy+EVBlTjrtQRH8utkUUidGcjGkQqIFj
cYCtg2ADzuKR9K1/G7zhPqJaUs/Tem/2vYqrXXNUkhxRziSFNo8y4/XQmyofgLuh
Y3WgyVUAbHf9DjjscTmFOrbGrquZaBENVbBARYodSVSCnSPr3Tdu7ryRr/SUj+Mk
1RzdtdYEYhyAe6wsvFh0NaCxEAmfllxpAQdRviZg7+0F1ZyG3Ol7VfHrMfBMzkA2
zzIhba4Evjb/jZGACkVIERKZUnlAQGNbAi4TMfLr+AP6HTGiZy0avJ4Xq2ODXauW
H/xDYa5iL6P/NbrUkcFzO7w0598yS7+C+g2rBvzrSFWxfn/Oiqyuvx0vN7iT5pRW
KPhrzsFVUdcCFqe3dYs5yQ==
`protect END_PROTECTED
