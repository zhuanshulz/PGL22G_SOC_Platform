`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mw+1NKjNd881l0S3KQVhB1QSibTp3P+eVkTtrg4vJ40LQ3wa8nTj8KnLsCpXyAG5
VL+NbInoUrIzfk8UKckmylCaO/azWm7/IZiJRYBtNcdQAz93C1APm0OvS/xq43v9
ZC+i3ZDpHqMl7CnkKoie2uKkgmIK6CHy5x4LdAlzSM+ToljLgl3OBBYO97kSDFhn
dwfUTqOBLVXUzYTdQXEE63oyySVuEtkXS8P7oNlsYoIm4L7H+nC/USXznTAiUxcX
hNQkQXP5hqJwE05S8G4r+WPAfIqfGHF1YXdU6kJiWy5IAp6Oe7jgjJDnJV7qGWry
/ZoZe2XOYm62QuGZ4J/0a2YR+4iEv0B2Y2A3v1pZLaOsCu2YOBKQJbIK77C87k+V
HEFCMiUmVhz/EEsthjgADO67VEj/SW529BKQzjC5hMEzLs2kgyEzVJtx7HUMxpzO
AGrdNWM9A9tbu0efx1s6UNNVYaRbL1IX0We1449/bkNaj5+VVoS3S38xQwjSL+Eu
JYGsMsIUsbYLGGr78R4c3wyLzamUdU47SXaKiovz4XI1uRNcMjoitSZtltICSlxD
sxah0LlPEsPsLBFrytcDKXoo9iKLRblzwLBKCvLP2njAUlAjHSHWtkxJBKmODdGi
8dYjlu8tk0M8jGeJpUvpc2UZKtx10tFcIwjKEbUDVPvbPJEDqWmadbnCQVAtq0gE
Y7buQtRzmd2Ln36RcYZNS6XNGkokiTDTFRNzNzhX9OpvXdUyYwuu9YQUIImk9cCy
MYUG0RfEReNb48q3tZ1DM6IYB5CUMlVcexGy82l7UE6g4VWNFUqLMWOLwhUdZ1J8
xJ95WjakGDdWk5fsPbKV8zlD4klazCzY2YLHwSdUkMb5oK1a4HpcTIA+B3hzye3T
XrtFgH4MIq+eDFf9BXAaG9uiGnjlE1pFrFcfm3XhmHN987bia8ZSKY2sW0k0+3NU
KCe8KOjcOFVTBnhpeFbk7SYB6TTGypRrXpiQkSRs2KJspjYM385TkUrqCm+/26as
ADtkrt2ykov1kDHbrI8sDUxFQ/Swsfyn8O0N+Mhkte5INV/bQvnKrPq56Y9Zo17w
tBIvSuf30vITuOySH7DDNbfZZxaB0hxChE/e+366SpQU+Leh7UC8vaqvV8XfPVpu
B6HGdKDfxwK1Kuwk7XWERqBrcGhjIQmWObjFKcOSfaC4sJB2Y/sgTKZudXYqORvE
lGi4r2wSE54NKmlv+pP6QTSTwbku4IWDRvluqNGNMIFN30yTf5Sqb9JV8hFi0ulW
QeWioIJLD9I7KUDAZaqiT6Sbc3QTt4UvkUXb/MOtMKvTS8UERSGIOGNYmdM7vAXk
PbTYNd2g6ZJJSRzIvlNX5/751kRXZrerLpEzGJRoEnmQYHlN8IYBZ4dxfaQIqX0v
cevov2ZAP1TgWMpT1CwPUyIz6VzUBw0bcBxHaILeTM7I9h5Kw0N0jXQLwagLi8fG
U2YgehZ5Ubfvt8IULc4Clt0ZqF1pPJRCocwXq1rSvT6C7/pYYJgUuDcuB7PC+jyZ
pCY3nUu55SXVWUPzTUNIkp7N+36eKuXZN6O/KXM8TbkyYvj9pE9q/fAVlnUe2N6M
+awpTeBuSifTN7XF5Iny7tI0MkamR4oQcig/S/DB0Q4r4C5dzE66VFLatQWdZSRC
/S6GM6XOm88KX8SKR8nwheIzUNe6CXjvi/RcVF2U/OxdVUNN7UFj4tMIOie1Lck3
YcKHpc6oaR9NddiRZp9JEjEPOxKKg6pYl5FhTP59RhMWDvbpQks4i5vOS8VqCtcW
oeBNzebtRHWoAvXQE4Y1AHCUjWIm6sgRuHdZ+2vFm6hGGGICx2vDeGBqy0zgs7p2
Yy2dh41RgVcGXxVuQBu6mPLubk7evQLaa+L5G9/hItpPMZZGbvEgV6SnwYSLF7c2
FLtyCE2Mfy+Y1nnxwkZ1Sp3T8i8S7Zr7sjhsihqQBJ7vDJIdUycCH8RxfYa7e+xv
w8W7qBvIGukatsfGKiLmE3FI/tad3V8gwKoW/BIilIVvxXvpnjcu4JyMR6pPgiRX
MknyxP5+5P+YD/52y3HyCkfSkLPTDPN8yEWi6jC288+hnEDIsJ73uRGiI8HjTFvs
+dZK+7SIZzDE4JD76SUU6aXr8LgNu/qx5fPN7uMVbhIA8iJhysrWfe2sr5/pcRuL
kv9A/Nxz1RqKp5adozdTjYsyNTO/IB/MX3cs2fs71tIOAwYAYB/gV4hpke5PQ4+d
Gz5/neTS9VML93SHJ8OLFKzYXVyMde6jXq1GxD3mqpl6CkXHCJlUKtKpdmEmA3sP
Dbjl0lz5/1sGtJS/C+X9b+Edu0OwS4X3k+3W6YYwIjb/mHe3Zi0WO9C48k8rlH7Z
XLeq3m1jIx0+N/TRGjxcG5Qx5Hjov1wGcGGncYnG23GqOKKBQjyoUk9ZcWz/mpkX
EFDrcFEQXUMxSaf3gjkeUwNrFp3hDwfgtDXTVryT0ozaI3RNRaWXh8/4y6jK1FQ8
5n7nqF7e9eyJB3DiiFBJ6E2ntp7nrQ6H7e0tIuWmWmyc1GJ86ixxq02XrJ6z1vok
r9EL8GayzvS0j5K6AWwvgfYejRDzpGBCbmLZUFhZC3p1V5BTfEMQ86IppIaoMelw
DKkE7fl2f0SBUrOLGUa0Q2G2MLGe9//4ZZHjwdVv/Nf/OQ1bHlo2vBPcOonRdeXX
vXnxFwefuuQMac5M5RJSHyo2ipw7VYiczMs+EliioSoP/Ufhp+4AG/vTcfwNtYIp
caOZ3Tweq7rUaH1Wh5cb6r2bV8zJ5XwN5zAO6lFj/nT7rpSAfCQAXZsWoYpmPawG
U+hHS6HPFQVceF+VHqQoD+Qcz18PzHGulxsnQt2twQz2jfPQdKmlACcSkRCtNsUr
B0ndTYz/QNCn8zssXURbYQrnrJlCVmdK8+SFZ2r2Z9ctBfreu77cQE40I8Q47NSg
Enh7Jwp/m1v1w+DDVtPO/pMCmwtwZ3YmSNpfec7wRVGFxODMzgWKaFNYuVNGd9oB
okjhqvhBkD3Aj0M/QOBJbajPiaWC66Y8DB6SSKvmV5g/NCpRB+CE8/07qeU6WU14
La6FaAVrzfCthg5oVzBjoiWNzL1rkwy/uUNeBR7Mz5YkucbVht+GAgvvF0qnGJpD
1MUKuznPuuMS0GFroHwJL4H+hm8IEFr9kGxm7q3r/RxYAETPZCucz0cv+yFUGcMz
zOwBWCvM/6XK4SKQjV1XSvEEdh0rf/z2qVbX1vt3DIPkhtAEmRGikBE0zEhwke8C
gSGnn318hv1+AUXBPYMVoymfFoSryi7RjXeWtGE1hhKZNFERNefDn4MQN6TKaR8P
hCnW1b4SecguPwE8ersVpSbK50U32jPFj1hw61w2OtnXYClP3Umg03HFWLLwl54s
+oEAhebdRNIbtEAwLFdoifWofEWRrLPYT7opVxAHNLmAh92XXmv4WZz4NqLaII7+
d0NuRmCKbKSQLht68cWGWiSvbLlTaO4VmTY5G58JaxGJw/vPgl5k/bnrAgAHF0jN
R32L5i4sJ1Yew55g5GiWMEHYeYek1UFDCj8QRkORn9K9gTV1TKpBZwhetbp8L+Wb
PTmSJBIhGMBK1XtyW0HW0C4mHJXC/wu6XW5X6msK+3ZvblFS0Vfh9vrVWNM429mn
Idtx55bS9cbI32ZKYR2zg/RghiYODOw/Fo58hJEHUSDbt0m4LemVEc08SjIPV0Gb
h8vgSqmXxr7rH8D2kRgkiyjnHH8iHFoWrQn1MRArAYx5mbX5xVTJEdwnyVTWxcHA
d03QWWAei111Ck0LwuWa9RV+2zZuyDoBUq0Vh7fVUNj6qJkWWYdx6U/9+u9a1yjJ
md0OGN9t6W8tt92KJAtqcCFNoEi7oSxP3iuJe9wz9UaIInL2Pkzmaz9bFT0ScIzR
esHWewSPB/PiXaGEcmBreJ6tUedmIFH5GIExapprq0iAeFKdbscAeogq5nJVoosr
wZBBr+1FW5FVYQdCgoZ7nWUkhnfkIERaY9VIOZco2QF+o68Q7r3R/rurZRyDoyrq
bztTZ/w+3AU8dshpgiQ6VA==
`protect END_PROTECTED
