`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0sFPlpnvxQtn/op0pw2cX709A0p9/F+TCGhfaGb7nH4B3ZF/LYn1/eMQJERsAU3N
/CcchB/vYJAn81dlTt7wPjTdMIT6EgVz/M8UXAOHsjIhhFlPPykkmKxr24TpePcA
mJiv/GjrNc+pMfnMBiIfum5CKcUixi+Mel0MVnkM9fNIzs6yOzEl/0I4R5ufoPLa
KKOZY+ke0jmsDdlTMyaXZMw1JaP/Ozbb0Jwzk3bk+aB4/nTChpEYJRKeXfb5OHOI
ywvlpYJugPburs/hRkRGV1rpwP8Ghp002CtxgPdhlh59TXwNKgLDVC71+Zypj390
00wZo3ZnTRVzmw63ZqUq5WzU2bZC4DaThHs9GZDEqCFdLEP3huLe5vYtiPzt+wwJ
bghmfV+pCkjMDTQlmR2lrA6NBMHPW7z+ty490MuLshMGSpXafXd4rpgUla/6cNwv
TcrK44RlpXfjcdPampqeppGtZbjFmyhRbDK6SNaIl0vYBHFPN+GhCYbUzaRHo/Bg
P57DcdFBxciagda2oawXkPuGPatCBm0tjiObQsEj7fzz0wHYoMBNUmw2k0yeuX6R
oCSCq88pkmGtuOsEhyYwsWmvDV25ACyZdrjdaGwWxuh91/9P5cOv0aZGNK68Ejm9
cgHKZHGTR1wfI20LeBMDBEEdG726CfGyvQ+XW9cFHply8XPeGcV/Ox7jD4Jps6Ud
IFWqVKXUNTq7p3C8WzICHDHSVO6hBE+5F6D87CKCefWrHEJoe34kFb9hEs5ycJfu
S2DvwJhHWwL/m3vxUZJvobv9IDlbZrh3qmtRwh8j3h3cSUpLZXeLjLNlrpOTWViU
ro5A5Fdz3g5lrFflJWyjhfJbrvlKnosCXAWqjgyJ6QJpDPNqa8Dh7WDVHN9DYO0Z
3G4a3TvK2x2tX9wFvCe8ei6JLgbh531PDeZelyAk1+1C+RHciDtBIhDppaZrVeMP
`protect END_PROTECTED
