`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QICABuedA/RlmcgCv0HczZtpTjV46E4p5RbmsFGapAAdCnFTJFJbLsAiIsQ9TM3V
Mt9l4219W3Mhd5uS5psNOiKVQelCLcZsaVtpNfHy20+80r/gossaufoW0qFCCbgL
2P5dxOeLJcx56SxgNfHIv7yNcPCiQkSQ5DfFbfvxgRgKCNZAYWz9TcsrAV7Zn5mp
tHEts3vlkC+u8YAPpLsQRwse9VRYpsny+t9EK2czf2FI6hdA0lrUIgyi3qlLaYZy
Rcm26dr1YXHrAWb2eD2pMVY/oQVPWce9yP+TU9TMnbIppa0NfQWUZNYjB7EL5r6P
GcyNZ02+TIS8aJIQagG8ospTi/MtIwQynNvVuGmo+mf+Hfholtb5zwGpMj4tDRuy
YX33sBdLxKVQ67ia2m+3R41xuWMKYC6BTd14MuH4sHyFWyDr5y/desoudIR0SbGY
/0FYzJ+mC6rrebqXu/nWwlG/7VeTWB2QnXsJK48SCSH3PjiUmfHEFMMB/abhnLD2
Imm+/SZI1pD6UT/gctMsob/VRH5Z5N2gjyBxMFjxfkscd7lzBN4kYDKHivQKZXc8
utHiwSWeuwkIUAWQmQ9J5g==
`protect END_PROTECTED
