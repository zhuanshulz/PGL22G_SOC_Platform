`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FjnGKEq6oj6wXrf74q9MM4MJuqn9/Icrxoi3ZoyKnbCq0El7UZXnimsGP77EloOB
345xPJvYQOj/fu1fjSHDkbaltsh7VJq2qUMM6oVkFJTy9qVr/jmwQfFxoxcQ5Lc5
zMIF4dHzyqzswzjptX53PlQb/D2Gd9G8FrZNfzbaitBGLA/lGOJEIvrcLwI5i4WA
7HwnlO5aFGPRxjPKcV513gu0Si11B+dWDUqydRjQgQ3NnZCY8eAdoQ7rGt7QYm+5
u25jTlFqop/FpYwalRE+tww7U78w4eRpYmkIBl/yfrGgm+T1ISdVhbRq4gNRt+iy
C27iiYtQx1T+gZn0yEtSYSEsMnQ+u+9dR+HcA9QFNNkUcVos7iEO2xSaN1LvXnmx
HitmL+iPAetRAwGmLNEpKK41h1j+mmA0SfJRfJ1jg4t/yu7WQAqrzlKlVWn0OESQ
ToXWmvuhzsQSW/xUlwMVJocyanH1IheWuFjon+M/+s1cRfnwYNq7/uQAwBbUqGWA
Ys0jHxZKH29OYczJX+gY6fqqHFLebhuAlmiEkEJdwGVK7Hr44VN5c8UWcf6xq7LY
wkn2dln6WAk2TS1NptwJLw==
`protect END_PROTECTED
