`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lLzr0Qi9MfSkMOoxQIx9zs4ZxSViQdmyR3Z4ycYsXRMkupUg6+2/nNIMNP5iU1jP
uAX6B/au/0EP4OI+h1rcIAgkD+30VBgnGrxl4mFyTD/kyjRSd9fUYWYA3I7QavKg
/m/0MBFkT4vqZ8QNNaO/oTnmfaD++QEIxJsSehlOwb8NgbVXbwu+KHtSb7oB686g
loxg2lT/V+i+dbBjgd6z/h7ucoGWWQiMW4x8SBlpCQfSJP27jPOQNM7Iz4vHYnzh
wRt7sMbEuDgB2s/WdBq8i4OIWyiRmhWtyf6gtPYe++OUlOaIeOgen0KZLFN9syig
PF/L7TGQ4Oifg1og29HqDH+hinqG5QTwq+tPU6BB/rspv7qVGTEUbovgLfvI0T+d
88LMTpDKlAAFo0HTBwcjA0yu7Vt8DnnYhVWAH1Ska29Le/PohaHGXFLkdnjLg869
/ZI6JgwyLsm1c0kWsC9Crzphjzv9Rwe9qThYyRq6UKuVx7neVKF9rh28P7kl/eSI
I89m+htt+90EVgnWaIL3kyC99Tqkp3PVbAtmijpjrNo43oD2G3rm46FWiSU2unjt
FS/rL13xgJXP2kldwplw/8woG7w+c6OUkrpQ+mgDUYjfEa5qUwT3rTNxjGv99CFM
vaWX0lZdOcvLyD1AQhU92HEwnDj1nkArKD+Zu22zB8smrzmTeE6EqeKChYSHFaUE
yChW5OY/Q5nWi/tRVTiftL9+xopKvXGpsupljOarVMgHStKURPhu1TQfaEA35wgP
zO6oyeUWU/QHJfhUslCbozXYfE9XSG5HcGQl08CjV7NFzyqLm0lrMHT4ivARj3ju
1yes+F/lts5AhsbfuAMoHsbrd841mWaSTi9sgnn6W8SfOE3TZqhRIlS0SID/R/tO
Z7j/8IM0D/Z2GhAiJ+oxoNLztzxlbQKb2JmnJH3x0Bo62lRG+YEG3PZ4Py8Y4Zxq
xiME5bd3wxARJ2kJt5bSqnP96Ecz19GfcHsTb5K5Xtm+DCK/IdDJCzECdY2g+8pN
PNkGFOerOaR0N5H6/peqZoSJ1IGktSXaUFHJDiIPQRSLZX2AM+g0HtBR2VzjWwnX
jwGZA/aGcKi9jSl5zHwb4cF7uRcF4T8btoASFheO4Gp6wl+6D0cbxKTAPed23qEa
ADf8OJeFAG+vPtg76OAyIHK3e5GgQ8cQnbEFIxfbOmju/dhotqXBW+gsNH209/dz
IsxvYAaj0CEMpJSoWU6/okgdoVi4rwpZGJAB7nU6Yd0f2s70shAlYsOzfKbxRNIR
m8Kbl5ZCTK3Yt5ug9QaR/z3KLdp/Y18RotSeeK7CM5IwFYaTT5UFXizHRxNR2a2W
bHQnv4ALhTq/uRSlbWkY/m0jcc9nWnnBNxSuUfY1Rxbmzd+dBD6aYu5rep6pXmIg
eRAblXrs47bbmck94LGYKNxMPFfq1D1vsrSkNtr5xXgdONTGqSI93M3nZKE58aF5
ku1tJXrs8iJXN0gPIlM7B1IeifOIzPK/Om9lL0miiPLpfMFMSBf9DCQVantN48o3
tC7Jaq60sd7YO0VVpqu3nnN5ce+UKl7B7K43t03zo7k9gxBT59FWGfbF1ytE216g
C5rnq3VXp2Z5++RsrBx0hghmRPLAHqbd/5yamngNuUHjAkx/sjMnCg9ML8cryO5y
XLTKuD/ssD1e7bQmCzpoQI2TvkUTQL663a60Xrah+MMWe+8GqOhai2IgOdtPunKU
4Wfkw4+eYo68/k+l5BhSHKUwztyrLJ92acAV50HK/2ZGQaCM2rMqYBuf6VMtJF65
tBddezrSWlWCbdp6VqIk4nv3kuP4z6F0EDbULNQ9tB9w42YQ9lcAS3mT2GU5o2ID
PsbUkYPaIlAu1qI+zkBrefUY8UNJ6mUABdJqTiW34l7GnUigCHA69evuAXOcxS1p
Sr3u9REP7AVtOT1hhysY/yrJ5vQOrdB79mQtGb1mKJegVO+7mokIs+ml79+cS/mE
7D5fFiqroyW/jyJtnM/NMx9EAOOCFUBP4BLYGmHwYozeDRlu6oyYTm2uiP1BWExJ
El46d/b863j0NpGazPjdENHQzOIQrMZFVUTjQILzByxIDl69y5N9SuHvHniuWxAv
i8zK+HLQ41J503p4s3yrg2J5j4tm9WmkEDchj9JgoP+wx0UcYN7SHPX+gVtVlsL8
wLV4HkMBALDQtQwCcfxXfDm/88Odh2LXPaw5xt/9KBFQ6pFQwPakGmGsB2i+XKS4
DYfyzDtq/o41MVSeY5rog4ToLfDGXeH/J/duUISG7i4Drk0D1aZyKcKyvFjiliMw
Adi5BBi7YP2vBvc7B/7ecPrriWDd9Khz1FCCUI8oz4Aw2boP91YBU6WB5DD+RLQS
ZsnjLFWH2jfILkRESamvxR5FL5Zhn5L57X0uejdT4vEPobhTFoAI8t9PHYyHkFhN
uXL3g/LiV/lcJ/zHSxmYVaDdFbTMzNZm09P4drq5oxZFXLCkXpXDsXzyq26/VOz4
KqIty0iRmxcMvhiQwP2CK1TPBpq55XeLrqwuKGVAMPf6bwSgC1YN/EZnxPWzqEq1
oBrtSyFwxJ44yaw9c9saX/VWBIzkaJMUFCA1lLYTkEuelQm7kpPEN7x8bXQXDLWc
8BMmNOhgKrYz9Bf8KoO5EaaRRAbN+3Epvp4EfF6Yl8hBUUCT1ao2CJFRM6NU2wsd
wvpjZeSC8c9wbbI7wTCw5t+J7KCEVXxnYIDoUJQfytjjacgtVAi7qnTwJK7uOFip
teSIZ5XNjS7v2dfd4+d7F7/HUELS5W5h3Is38E16upMCN4IXNDkiHa+m5cWPelqY
E2UOlLlYVR8+MQQngnU1FEOA0Jn+ikN6q6CBxkJs3cNEeqz+Mw8JT4ARYdK6HDVE
DG3skEFNnoicX886ZbK/YR1+MVfG67aO0lggnJScIIqqtZlSjdILJIZnxa/BpVb3
Jmy3Q5Fzf/hYfIsuv/0a6SXpJkuOxNyAC6Cof7j3f4wcOdxlKbMFcnXpM0FXELMz
ak9H9TmE7ZAR74l71kd6z1hx7RotnXY93GSHv5+sRfqu/iOEhmV9MAkoAPxKiSOK
fGo/XBdcrGkCAkSfU5o0po6KjnX+Ak3qz6eVsmpOZBVbN8rxcl1SNoaEKchKySfZ
ysmDOuyIL11w2dfXTO7mHxAXpym/OsZR+dZXvK6hPSJC8fRP9MMN2dHvTQ8ysLkB
2FuDR/Bsbj52AQ2Q0anoQCmPFJ8fvHxY0vAiZqk5Exh4gPGH5W8KMC3Ddt0B9B70
BZ9xiLouAKoaug5WLx8gsjxx/BRK+1to0wEBpkFE66DLnGvEEgZLGEPnkIkJiusR
6wPI6QBoS98SmGmu3Lq/0KH2KLK5fGe+90EDXiyuw/rGXqElIjuqcubGdg2OgdZ+
NNXI65RiQMgI9UDEgl3YX1u013CxqjjXLbYxdk42lr11e4WBJN4u/NvRlyTyVmOX
6lXyE1rees0q0VimBEk2kwinZVGpH4NzVtSwtRIIcILTgaZ7dbUQThFfLbekCUsF
PEC2DoE8LNRkyX7ZE8E2eEghnE0MNdTUtekL2BYbyto61Dr2pPE/HeM5ndLnobIV
ssFshI9igevwFDIU/mT+GRd1jewjt+bYujvYpqIKmr94+XQAKW389Kf32gEnJk5a
35DCnVqmRsyal8awiRz4zkKrFgwbVhKCGiZCX4j3QPW6EeQS/uygR3uU59FT8lS1
/A+opmOeTIQozQ756mUGarGXagbKjRCzfu3sqH1UmmMvLET+xxe3ZsSkMbbXE6N5
huFDVQqqBTlQ68xC0QuobZo7kPlhdPxOkO9u0W9Resj3H5j7Pc8iEYh7zcPw8Ddw
Io3QzR+IhIYwp2pqbaCSm7g2tCuzi2NOvAyqp6tJ1mbz06yeWQyF1dpfdVCHGCbB
OBYQsp8gGKPAR7ZSvdJIDcweThUgw+JRpz+hn2gXspfPosMMvUPNlnyS7KBfObjv
sg5eoZaC43eOhCi1Ks4T4g==
`protect END_PROTECTED
