`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mZCS+4BNFimVmXEZ5F4CbLn68ThLF8yGXtEBdflWHlj9vO2fwpzU8Yf+Bash2yyC
991QVLhFeA4P6Vg5oA0i1/GEMG/zadMXoQYRlvawz32ugTf59SFj3QrbIp1ki30n
akOneWLYYch6+T+DvsyLSuWNx8u231GwiDeLis4kWOeIpHhfnB71mcOADjallSof
Kr8kC1uN68/pJkBVlQpLvDcjFOsQVaBNu1jTZ/mlyZbWlCsoBOKhLTMjkQMvRqj2
2nt3Hu4vhLQ8d2iZu3wlF4xE/1e8FHGOSRwNzlpzZCAWY+DA+SPDnDLhLKAXVX30
rfkl442UKw1iEc7skQP9Exko8Wfvc047ZgQjHslU46hibyrB73vkrYv7edI1+hMn
1O7m6WIvhGSZTU2rV/2xKr2M4pF3l9U0bD5H1ry98d7GnSi1oMBgGYY6aIo6I4dZ
S/ElwQXu8QmfngHVlsOIxiT42enxstTGFMZ1HwEaYZ0/mCJATPFULSu8tvJhJ4wt
IxIuc4EjJohRZFob9UKq+x6Nja0a3Y4Zi0rQjTxbsQi/zvJdTt+0JE7vU6b3JJnb
SJEOAUUPHBYm3216fSyp67+GM5Kxk9T8AgfX66EETrp/nArunRxnc9Q41dHWicbu
6qAr9rPvTZMeG/ROakxZK3wBOzj9IdFhahLomJJkO/Amqjize8i/KX4Gc9uceLOk
KE/lnHcydJgt4vBXsKmNe09GNvMf0c1BiKM/GJL/xg/GWhaNtUlmhiQinUIGPz8t
uDv6movn5+d6WZs/ab0pZrusHekIt6DSk7mwIVtLCAIfGSVm8qXUYm0vShVOZZfN
UTOprIkCgK64+om6AWc1Zg9r6+kCQHetAXdq8nYO+TnYEyvKKfu/lgjy/XcPZf/s
NCU/qOVVud+2rWJF6pJCWQF0ZdRRi187kB+vTli1gwWHAAytS6+HpYQOyEPWxGew
l7fWni5IQqM0bxbGLAbH4jU0bZq2TOtazV43DQQsqVc/AVrWZkSzIxRig0Sda86h
dBMfhbeURoLJSIe07zWmKgg2wrl9sg+Qo9ohJuIZvXyAOlAsayQcYLFZQwe5slcR
tTEvGqisQfm2vyP7S3wWeJGKB9ivPH4noKXv+H/w6Jp/FNho1aezJmZ8VVrT0Cvv
e81mSwjXlzWaWiVLsDNpEBIA06oqYaTnLBh06Y8sIYMKF2gKUHuivG380mpF6qIl
NPh4UN/d+h11288ORljh07ZwG6Wj5RoYYRHy6TwqFz6Y6QZ5p/diGordd3MjAwaP
GbqBvo4hY4WZmBXaO5WDAsEiCPHKgfCPydLt768mbYK7WmPc6tMUCV12wIq+gNCz
f+vJyoJHcp7DlNKd+tbvPlt5G0ckPMPhGEd9gL3zX7e1VHC1S4mtiX6KiRPPnu1V
4gf4ToK33DRevU9VTaqnn8/q0L21GnVvRuiXo+mpG3iN3jBMBwi+vw7rHMAJ/Lbq
tjdVQ4DW6Nb8khQ3x0opGK9k9wAaODRivAad5tta7qdseXH12NFxrLw8rmy2DHeB
7O54IoDPzviDa7MA06n9+AypvjNeJUaHdnrFx1b3vuYwb477MJ+VbOZXPHnG/kl8
3JHWSLPaA4LWH09am5G9XaHD+nxGUnjbB3kgK9AvcXkzSxbA5OFdA7rZsU6cVTbc
RtNut1ShdSWb48tR+I0cUHCFpvAtAc/XhNSMLaskQJgeZI7sdiSqLwHkc079JlDw
i2zLSVfiFf41kqAl/haHAjD8kNDD/XuXRMMuMsUvHxzeRUvq7B+EFfWaExus2LBq
hHpn/FL4DyWox5aG2W8W/UJFgXl37g3WmrxinElL+r7Lt2+wrK688JOvB2MBapPz
IQPu3fwK+wW8n3RVPwMCPZJNNq7Eq9cGeR2gLqrUF/lI3LjfjuqH3x9wDqbYIudz
rMkhFFKKdnu9u8I8iy0vyQOdBs900klrI1wruA9xKsUtowdW6kA8wV5RHVOWCl2o
NNeKSStaoQdfCSUQB4K4U9bJQ5p2Ti/auM3IgR6ZzEizI62hD67ehg4yFm99dv1D
3CYmug0WRk2mxuCw+ylv+b1gU4JDEgJzU7y9gpw+TOi0TEHy+553xWft1laUR5jj
PKmwfyAPXn+iCMGtGXwTddvl8IwD/WpmBt6/nyRT6EsdvypgGqt6ZzFZeWPveG4T
ddOwQSVvU/nj0gcb3iGQLnoVXUvpxmoEyiWWMWctYHqwuDQc0wGsKX+g41N4EgoV
`protect END_PROTECTED
