`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eWscfhKb50Umc7pU95dKrH6pwmrcIwMtf0GBg22wqmTUI5CiumOBj5FyhfGMSx37
v81qMxs6EEV1czfxa87mHVj73odSSCQfi9PBAJIuPI1vZ/sFSMjw3nFLpdjytfqN
UhHnLOTP8Q+PkloqiavaIIdkeqUmhKNbR1uQUgbzKEUcsDNVxUsgM/XN7N1WDqi6
kQY69Bci+KkeaH9W5L5ZE5t81Dlmuq0Z79wz/yvHgaM+DrQOCTTxSn0Irw9NADgB
OA2sg6IRKLAJ7VW03NUU3DrNV6Ie15D5CrD6XYCvGZTmzLaNSfcmXI2rZ1bkeWAn
AB2r6kDR55oW+k1yp9hyktx+qrNfZqLkopXtgTVHGFLRMwtLzEtl18wWecYco6cM
lXPF0PPjXZuJGHOD4WnSbV3H54CwpUEmxi3OTi7+fy5md3nOodgCjejDnGNYZuXb
LiyXmXVr8ZKYSh+4bhd+zlRCdgBKAzRlxuUw3QuWqoIx565ImDm+k5HSsXvzwrWK
4AYO3h1n9zahGWmF3NGPmq/ulZV8OOAwncwPRqm3v/J9FXJKuISzEtSEQq9ZEltP
NbU5ndD0ubNNoQqNOSmKSIouluia1oo6MDT3UcBRqrd/dZkXQv7x/oq8EEGOdKbg
A9S8XbWnmd9cVOSGSWX3TRH00Vf8lWoNqZRVMaJcJc5bEUS8hL3GYNYvZjXnMzx8
X1sPwRBf6CTlzpfdiuLA3Et+bRQKAL3Med/L9Iw+rRl6JngLVyZfKQGVyBu7rJT7
JsOW/CwGK+60J2al1tJjQYcTtQAqzd2x2vfXSbIjwtdMDbKSa8xpjQDiIq9AdItB
18Tb1t+FnTjtL3ebbr0pIjGRtnzM51ThSjFhcghyDggOjd3bO1OR8mD8qE8TaRCn
BVe/q57soN2KfDwKae3IIJoIobeqWAPBuQ6r/6dLMNyK5bQjcKi4Ph/Gk9SHhCqy
AyBR3LH4UtI6aZWopj/z7co1JixWQV3Zz+BoHAYwYkIj+Ftjk+RR7SQKoh+njLY6
JQZhwvEh5UqrHw0IPEoPXI+rzAln3mioLqNOt1i5v7zK2B5Nv/kxQRGuU1zR0AcK
oCqxdsfhUCR2mJ6c/OBVUZcP9g1tgw3OZfROZG42281BUozhs4Fi9TVNaabF33u8
/jJS9zeQOk+Hxho5mHUTod8jKYRFmydRICi+43vizr9EK0ugNAAx9/xzCzobMsgv
AwFJyRHAIa7fU6Kzf2KvK2ScU+Y4fXfJn1dncWkilfLFaiMD7eZ/6Ajlix1aAJL+
iXuWidfs1fz2XEbXC+iz3LM8t6Lfh3LMJtGcqqnw9zo=
`protect END_PROTECTED
