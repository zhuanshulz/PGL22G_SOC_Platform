`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kjhnGQEYOlDmu2t72WwGh0UWT7YSsEu046inVa5wtIj9ZeZB/no8v5S6t7rahc2N
ZyCLczGJlY2GMLmDtlEouuWQs5OsPb/qLSRTG7DIGptiMowYoCwXP1tvuJMbA7jv
BUyI7N2dWpanej9pjVMSCxC6KCbOa//JoZHJOotiUsE+0AUiZZLs0qcZdd88ElEm
bH4xPbtFSCjubJPJ0QJaVTadfrAKAemIrpFX+ZSjHi/7b+7zSNq6Kb/zbHWSA83c
PUONwQ4alqQnCwLxwqy7e10RBwI2kyOHoXak3U9y58HDabrTI7xJJQ5bACkml483
pZ5bU+PDWITViBgfF8c/+oMH1qjU8m9M/sGWcJtiLwBg/T0zyBgyUbHpRqIfEpjQ
gF9n/4V1DS5xjiJ2Vb1Ka718ad0X+XFlHwfyst0pJD9+6DClUBfEdjVowaX7ZOam
Lgv3f/EECGQQ0zrBytFJj5y8dACrvrWYsOIJAlIkw0rS5PWLrsBNV22BKp8L0FAd
OVi2EHlBGmSx9xjX0eNBIzDhSJgewfo688wMtMRYedQ4ZDWnXcAqML2xz2rJToFr
tWHdNmRX7DHEsIpQQ8NZAxdac6KG01EDPH3ti4F/Ub1MTaOkaT+giZTySJkpxfO3
jmSJgP1FojokzWD+qKWZJlmmfoskj0TgXQzDz9moHREsDr+7TA1bdOW8wUm5JCoj
FtX8xjAZ+GQkngclZsJuK1SHAi6Nql6QH1dQdC8qI19OkDG+PkJr6vKMGjFUPuZe
Yyu41v9338s6ciEkNPPX+I1TKMErP9XELqZEfz9i07xpPwWlhhuruXKv3b3eAN5t
+X5Yp299xaR8vi389l1DGZDEPGK2+5IXcFgrsNyVTxq5E+gRVMim0FlssfbSMjpi
OCdTi5Z5EID0hVzjaM9wRmmrkbip/eagCNyASSFdTqqoWxDablzkGkkYwxBUQqXX
DuXIven/UVBR+uhsHhkgnOVzqOvgYGOCByDEONwuKGuUBh0vkC8bxNBBF/JH9npw
Jer0jq5HjqnUEtMYWtbeZP5BsOqlue3Q/3L6hXVsnvT/HU4v4IeBtQHMWlrIlpkT
l7EKmRxac/Q6QNrk6lL7Q3YHr2li/28EnlE2x7kX8NmQyxuxlhsvaik6yHcocblN
OhzBHr/be6HCUzQW8zI9v/Wc0IHxBMSGYU0cP32BvY2q2LJ9/h3dFTlnVZTRclmL
goE14y5Q2X55zDc47uhEF/uV8JzjbGRRlg82+y5SiCguW71gCQtWrX5w+e0QQ1Ap
z6tIxwLbiqGcbmpQzr3fYPj4HL4DtE7Ak6utbTFb6awPTu2Nd40KranrQJDHpsLk
n0mq7+XH2FredhosgQTzPW8c2yTfvWOfxZR6eJRkHAmElxi75nACFU1Lsl8KGIYV
xChnlFcjh7nw/eznJA6XLHazFplywPbMtV9qGy0Oz2hIdZidNeTepFo9cSiL7Agc
+0S0UcUmbRemv/ldDjtAoM1rVBjk03h2q7PK1qaU4YEJ+JCa3Rpyw2YmX2uDcLNn
JS66dUfuc6W2s/YYFN3kA5sNbPTSkO337J5eF1mjbCMHW8MRDWyn2PVR0y/gISOI
6SKDgEjCTFO14oLf7xJn/eEby09klOiPuPjgOe2dXKKU3M0Voutdlvjtq3+3ByEr
ssBmyt0T4IiWoYXSi5Ar6hhzjt4TVItgRC0X6YS9enzaObljVmk3NqbUPMJZyiWo
4Xh5GHHTbQITX9k39iKsUFhmhDSub0EzAtpGECfASzvokObEvYapSaHZW/FRLot1
XliTxbDpwv3xViBxoeKfzqib1hnHDokQQk8MSbLGDSQlLRGbhgTNkJDpUuX4v4xR
Ft1nNVpcvTYiLuOB/L9M/ONwvSZv8jQhOwASFPFUOE9POiYKIMbsqC/bxt66d29V
44yRzgC7IZNOnqm12umLYQE4BDABdVpExAQqahrC/POZD4B2g1eAkDlFrDThzM+J
F/lP1L8hkDhU4Avme1i2R2skKmc8fxqsZV6xDr/4i7rZ2U/yg6nK6s2MaXmM2BMS
BMB92T5EX7N9LTS1+c8n+FiN02jQdC10JQhl0lkYXiEFX/WtgZshCCnHWwS+B2N7
h17zWhp31iZWzV6975yPiamLh1buo3mms1ZVFCEPz9NvoxKvN4W62lCsQyNVpV+r
TYSEaOV+xisgYtXnWDKln5VLQtEdupbBJrwyqFSUUwRzDZpNEQE84CSxo1X1znaK
Kk4vQwULqRDohjRN+DdfKPzCblbxswv3KEGcagKAAUDppgznRvxD7u42T1fzSDoF
5AKWDdjMJo8RJuNzad/iOu5T6MsgKGtH1cHk1cHDiJ3Cl9rDgbsE7abUIhg1QLS8
xY5slWMQsRBzUFdmhSsbcqKnWX7R0r/7g5LIUiZ9oIR99tL+joVh4ZxgUcGyvB21
oLVfdoEFkKiEgXDHA7VZqkTqms43j/ZzXSQpUg3+1Z/CHMGkYyw3/M8gzLtlmnez
e/jwE+SkCKcV37bvfQ9imdQBlNjGHrDQbx9KkXOd/NWxgnWx1F9WNCIIrmShA604
4URQbT0ghKxFfUKBimTlPbh1KXzfHmgQSSkh19TjFHgsl4dch8iCWu+I1vH+N6kK
+N47jugqUjjTAM27shI6HDbdakkRHexTT6va6qekyvhxDzhiLpk1IlJ3lJrfa9h7
cuaqbERGKiTnrvBGDqma1pAVGUbY8/Do3D/SzLUg62t+84h1OFXLnl68GHyFAEsn
12OpCtZt5e0PmEXXGgsOfW24IJhbQmd2XwcEvGuF/RU1xhi1fkIzPGWd1lG2eb2Y
8OzUqpeNBc7R0d1s835UNgGYhpKq8VQ4IXTgBnvh9iN6ErfiFVuWtTaSvruQvCnY
2e+x8ssFybD7y7xGlc9ADOvGc5193neuNSopOGozUsYwnl5oxj+ritMs/Z1xAnxs
pD7SE6mTkqU3TRV132DuJXsPqsCxMIlj9eCcG31hIRtBD6eegPFxA/bsluWAeNFG
M4KndinhpRI5n/mx4mQY5veTTkDEi4BnC7r4kH1VItBLw3zPlW8K6pPgVSQrr9v6
ClAUOyAjitRVsFjxKlLlDh/7FMWOiMx6rrOM+beaREnOOVRSHbLHdzpRjmg/l2Hz
2IClRYpJMsWHoJBiel3MVfh75JT8p16U9vjRUCholrnwZuvAYOFm5yw3R5MAJOao
AoWRBWk/IrV/GR+PlKbmCeh2YvBliYOoF+7CMXAWcKFNcZv391seqjkHCk0JNNCn
mzgu8IXf6IaKKwheV8FN3h0s9aXer9ZFNYNuoTVGbYcuJ3TFky8OObeXUm6kHJ96
FDcwQ/518tMhlEIxJbwmvrFOdNn4PHf+JeAIMbvXCsS38Wz04vCT5DofTv6KUa3b
iG0hYgggnbL3Wa/SY0u1U9cJ1u+ZtYzcb2KE/sdDCTSJGt9ysOavRzZX79PnAoNC
e9Y0h5G3R56l3oOaW3TsSxLSIZDLH40xat6M4lj9TQ7VvLTSUVXpw7Ty2VC2lNqM
RxvYhyE/Og6g8ZUqvzUVZMGwfToxDFCk+JjVuqev5OXWL8jzcJs9yHhmN7xBDtYO
VHUdgB3EY02W4C/UFR158dU39MTT7JQCWh6Rv9J0cug661dVZM1QpahBAEWAIbki
EiuqtJqkGZioh5NtdrRWs7pS70UoxymDhHJ9kD34NX9nzHXu3NSJh9cV0VcUk1mD
Vq8OrbVuxwjgD0qXEpV2pbY8cLRNSlkKH22GVi78rLGLk2WmNCgldHs29P2G9Hkh
yR+kHK2Th0Qgw8ziLia/oMtb0bdPoCo7IYKgZW+Fqtbk82M3p8uWpFzxwXYgKE7F
zcp7Evt8ccRdP/wQCMbIJUO4imKwjAC/GPBbiR1x00+RKt6gQ9iI1Ksdm8U88RNw
+YotNN2y+3Yh6ItDmXgFfzLQjKefZYlr/302b99Eivn29AaJUVcGB1USHRad6anG
qFD6RYkNY9EWjbhbdGgPkrTXIBufB5reo6N4dfaFu9ipPcB7SCL8w1BFfFXTRxuO
X3vehaed2VpE3i0ZUzlRw4sRNRy/DaVQiLR0HzXsNDOAWE+KMZiJkeqp1wq7kwHQ
+ttOuBFQtq3mt7UiHgduzNBHdQPXw4HhJO8+6JwPvbUngbYQ1aJ1bn8w2gRxfH2F
sv2AFQypsJdGrmKRn6daroWlfOEFzUgiu+a2gSvENJfXdqzNkcP2Wc8rdTmCSg0P
y7qd71R4INy7iLnCi1PT74DdHFg+Wpc5Xq60ZJebIP0a3Ad+rMvlgBCLHy9cph2G
rUeWN9IUXYJJb8MIvjP9c9k4RNLCWg2erQpHbdyvu/UND/H5EuVIxn3aFzW2c8vB
j2fIjY0WnvlghQrCR2CqtwnfwoTxjqWg0/t6m8UaYH+WWba1vUELXpZYSvG1ZGXa
taNsmCstwvWv7nfukUzx6MGW6k3owJE+yYArG6tjNbMUawNvKj2mAxe1H9Jzty/O
gubrjScrupi5S44pGbo4Dj4bV6qBwCmoFBYtWKpDoLlUpdq2oZOiE5PAt3Z8/W7h
5/fRhBKwrUNmqsgW0pWSrOkKhDjwqvJ/sH0RC/MR6A5tYIkrpDal2zcN5amRaJ4W
u8b2J9r+ou7OScc+6zPSwLNB8YBI8QZyzFjIlgSQsy/XB/gnSZEoHpZ4p6NgcNax
hQhuuymDy7zP1YzesX38tmPPg8NosOmzB0V0+Rv+FhRfJNxG776ZjF6qHb+/f3yX
pNalpufyswVzUdNfbg0UHWHsLOzTrksfw+VZowCk/ddr60WxzMOeOXgQ2vBvup6d
DJ5Z95pIpDHTRIppTEJnuqqGKWrikWQ4CB3vr6HS8wg1m7wgLH3lzygtAn9HkkPv
uWU1ZfLctHUvmKAJBQY3MqZ+vRzF/DxJXqHABv+u8vZ6TxtkVoQaPctDJFcmybfk
DeMefmgnd+e/ntdBFnWUtSt6hI1Si9MG4ZSTX9Xc2kjuGKGUVt2dACaDK9zVy7jY
r87YwTotJbtNvcZJVUmwtnwPI1GnwRZxwrwn8HkwfNg10LD8lEKbgM+cN2w18T+f
mopME81N/MLMbFETBb1yWtvAup4X4JWyVpV86TzqolRrSnqHFIvyZe26rWoRvDUY
OPl3qLVoQeC82Yv1XNyc5Bo0o7sodQBOB3nE3EbTSHIdClmBxhHPSM+hI8NHOsGJ
+/Ow+ucwl7fOmnGZm3t66tm65fdxxrtwyCkjW0Ujsvp1iQGTqz6mx95megzGWFvf
CFsPCBHN98kcWdTLB2hB42yVhgstkLv63VpYGyap5qSDeCgIohxsJ8JcMYMMGv8Y
nd1HxAUuRE/ImG3dl2Az+kJfwQqC0i/RtY0baySPjXuDUrqcEMXIFuTPrH6dDSZz
3TcChqbTUa89d1hnLkQN7bUWzlwAT+VWsVgEEIc8SxIBAVUJN6Atfriwoz5cMASh
bqLA37vzZJTmW8ata4qW0jP2RQg384WNjuGHrLMZo7lESKq1/C/z+ysPzaqX/FTw
BzGlTn6ZcoWj/zHfc534jZxZsnt8Dp4NmCwRPYQtbn3EU9zK0K87zy9p4HjqC+9k
PsH20DnlYw0g0KHpj04dIuVj7imUCv65Ewvx+RldIC6/z1sOP69rozlbcCNwu8Gq
clCz+v1VkRlM0NfE4j6OV/RmwV2WHsQWw1DhsMc3Gh9SkCv4tBtCvsFyxA+QNXbQ
LCIfjl654avPwGeI4YDnNMTGNXsJh87bckpNjvkaAAdM5ib1NgH9hIZ7Q2DxLRHu
5PfDTHCHS8kgHnjj7gPvSnNcFQlSTRpid6ZrKgmui7gVif2c+KWpPcf8PNeXXsln
zQppUJ5SGt3amiBYy2s1IX7ARWj5WPdHTGGg8wQ2XLmo1JCRp6CaslRDhO68PN3f
JmEcP24GDVpmYQRir/QyEoPbCNsW54b0KRn0fAUpYxxQWNyhvXcCDBrDbOW43OcM
sEvhUvcjGgD2ckHTpx4RINHUxBMrvWakpPRv0uMLrDjt/+cffWcEHFcQ6n/kxnJ+
8/VD2vKKp4P/cL3F/nISBmHeCDyq1k/oL2t3rH/yqJVN3pfZIk3yqdRX6kSj7oiS
2IJnAaY7e+su2YCXkhrEMc/XyMcb0YKLiYCw3FFM3U3YJaZxfT8rJPsR558yI4T7
KdxiXWGy0S1qlZj9Zm6rjT09gJ1xwJUZzZgjk2g9mkGxWyOtNRNYOpQwBb4AfGxe
dZOKocoe2DaO06UIZWiPE3VhrhwroJgEJRiWaSpWWZ4CMhGquQuvlIzADF2RDGEy
V9P83qIsQ40qeGNvi3GY7Z46vzYkM5MJZFCsIXCTcZ3GQv0/Kg8FNoD69sxRcZWy
2RsHPJWC1jLEWbavfjg61CguZDc6VuISOMw1YcDcoqRM8PmPgC2WEKp9e5gP2s1R
Flj6dUYYUCxAguU0ntxx7Gx8NXqyxPwDbvXBIPYNZ+1vp2N+vzMHFcfwLxW55YQg
CCKYG/a8UHOh3k+f3m1P2RpNl7qLbXExa2hPHe6pKwUNtkVvqSHiqukLxi+GNVQK
SMyRKj1PVwFQEJOsBLtzmXfe+JU8p/3UWpM6jTTh9Tn1aEsNYnh29jUOR6KUe4CJ
Au1CBo8skXH4K7r3L1NS39hpV4feb8Q7YwwCYIOYltHdHalZKf/sdtbjeakRLCoo
xnS2zUzessNcMTio05wa3mauoXTpVh/7PedvB559wtXGpTkOn0XR7pzOjcyEymT5
7tuzGlv/RDYb1nJdt0YCuPBDKVWv1QDMVjmneubhPzDPKlFjo1WEUKe7mnEiK4d+
MRXF2D2Oz2N0F4Ci0RqTo/ZDi4KMb8dPe+7/+hhluM6kgafrQ2uuoiWOnj3kJlxb
j/VRNTQ/Zrd5vZQ5LihqHMGKbq9w0iUwR/powm/Vyt8ZGeo4V/sFd9RirmZqiFDq
fmRWwJiOHJkkE9perVEoycmOP9rV5xm/6anFuStIAFCd2jTBOnaSh/Wy6t6mofS8
FUTEGcgc8piW/5jV16l1TYqKBcdfitnNFFv3T+circtMAnczuB5uxYKsdH3VVtkF
LBnQHMieG1sK0+wmy1mF2diQG2me3+56LCNiWETvcyZBCEA+KFtOEcV0PjB0fnc0
OcCuL7ElQMENh6hcMi9r+8fQ7et4xbn9uq0aVs5fQT5roIzOSjcf3QSCdCI7V0Vr
7EvYf9clxzPbRYix8pKhQ7vOsnfCmKoi3sCP9euPh7MMDPPPP0j5BFbC2xnW6crk
Yc6KFNF87ib/ymj0SePaB2MTQO/STZJwWTKGoM4HzHSZF0c+VmSM4vz4H5vtixLm
7YMAawihsnT/wUOzEKBYUn/wVkmmNRwc6CXVByIvipSu9ci81IotBRh1Sh3k3by3
suWRpsoT29ZXjfAKZWIO9Hhex8HDucp5BAtD5kYThVwQSno2ehUcHiKUtlQwZrSw
T7ZSxDxKaaO82a9RfZdZ+Obxk+6SRTmnPpw3PDwKNEDZnl2XA4ewonV7oHT7GLpN
s8AUkhqimp1VxerN2Qn0X/pVfgd8gPl00QVkbamKV+M0I2f/7Bm/n9LpRvGxnnGO
QBmFwGoPAmh9Gc/+2Zbqquwo4tZQ4apcqJnATFV0TKhs50Sei006FzQv0Svi8Otd
RPtaYCPu9OG681lKYLl8oMthI3KkU/ieGRi9+jg/wcbkJpqUirZOR+vAHCK5Bz02
xAy9vWwfv1G8jGx6QaGoykeFdtGQK4/jGxTXebJRKjuG3WSa74g98KUx1SQ0puQt
W6kQo0kH+ab7vOexSj7Gcs1hbLOr5kzIVoK+7AJGZnXSWNidHK58jvH6VGkDuCMS
G1qN+VLyghoeb5FSWPzNTSevCpn4aZuwjJ3tChveFu9OtAf3p96+YfXNfPoRQOQK
KKzlSFfuqgYixUAGezWaO7OCIUtP8Zb8DG6R+dw8diQvMtdQtymDfAicFn/YvQ1l
iIlRnJBDCqaClm0TosrGM1FrudAkVdQA1Vv+xkZMnS+rZTzlnO+sajnChi+xnJso
BmE4LpD8RdgTAggHFLIqyb4lVuo4Vyim1YBVRtqbSMVR40GBZ3h/29bVhnK9qWY0
c4qQCd+WreaqUlJuaMVnajEdxLMBlmpbrPhTeGlTtvjKZpzqkjIw4Lv6N8QWRjIu
6y+tzrHYX5Hzgp59aTHQASBWAiwjWzzFlc1reID6+tgWOX/MC3OjOtlPz1Q0NvWj
swZd5HkEnEI+FGfCgObOM54hI8FoTZbfHopcmL/+/dbWNL0CJr8uHd1RnJi791i0
gEuPmQ58HLDRH8YHjP6EDeRd+ysEgwi9EfgowwJM7oB4Eo4ktzXiwnC0KuN9C3xf
DD3g3sr67fOFJmVR5vnTFkhBMABlMOrVAtUicIRGboRYAH5DxIa/kikobT3cDj6W
hxKbgl6q3B/6kjtFr2tIFEyViJrHqviysrXHNf5e06nge0LJaB6nSYRRrzt1UCm9
pMPLDhEGLf1uO6H7AkpJZGyONgvhnYad99RLtE1PL0nla9Ps4OgrKm4mgaKvTMV2
N3xzekNNYl21FDFJGe8VHkB7lPvhsRdfxZRwJY8tK1v1oX1cir9l4G0bJI1i3V3Y
ll7Ub+w82JxrWaPVwIeuTxAWG5Wevx27Z/en7hn2Q+goNehlZcdMCHwRAVNZVNpj
LyXY3+I2Mtanv1vacGu03Rexq4wWal9egYTomNcyJI/xdcX+u2Q4PYR0wHr0HGtH
JcbiGbEc+W8v1rdGXYHdGlnYUfNKSmetWTQ7+AhYW58xVjpUhAGu5Vv+1C6/ahOo
etM0XrF9GIyFiDlQTRE512WynUuE0YbBc0eHpGHMlAYUUqgOcRp6D6pcgBkX5ktR
V3EhoSMIgEP4xYhmF1zjAg7bYqTUyFxhm4Hd6McGYCXalAtdjEm8mpsuAxxaKaWS
+Q8COsH3yJsGMLcBmZie98O2kF7+9NtTyeYCakjNIMvQiwS1tZ35ei5H6NxU6Yqg
7rX3psJAZcjf//9aNmZM56TU+AvbmbpZqlfwB1Qcbf5/86M3tvSb6RB3xJP/MKLF
xQuhw0G6oG/dsU9yX7HWh7F3TEqtOUaGETz3hAs2UL93oWt2QliUJeemNM5uR0TR
Df4VeD8ntTiQapTzxW5+9x3S4HXVHpSlZUXHelDEwv9eF4Bcdjgs6NAf/RCPdTgk
Ku1TuhzBe1fB2w7yd6Zp35n+bRZFPtxQ0Uol9fcqQ4/olQcmrAuQqWaN7kDg1qNM
CFhm3QylqrEG8Mv2Jh+MoVuZIZ/HY7ftzUkSkGUdichGoOkaUEOjGGPJTHRbK46d
vAxfQGGQwCSurYqruzsGMZf5/vmFGilhio7LPcjQKNUIpqfQvhQEyFvtACaRyT6T
HyJ6mTq0nhzNbIMvbFx4hiExr0k/QW0pdjpR1gU4M8mh5nnars33hTD80j8h0A2I
2/6xFIlWGbI8Ce003syfVZ+p79mxdfWVCRA/I2x2zmR49xuqptn/lhaCQcWgqeh1
hDGI5cdGXGQKSK1ZQdZygHtfDHRSE7faeWCMlZqYJxfgJ3AMUDuwy2VO335kpaCT
dZ53R4+n7G3PO+nbTZ0Inxj4EMxZ03UkGTEjO9qsKdLY88DnYYgybZCukFmXhBe3
KPh6BZL4IER+fL7yjIpEyuigVm+n+NSgOgfgmBWq9moEETkN5pNSqfTO2HgS7kar
JaFIxp2gdNAr+CQnvIDmNyQJCyPacPufl9e305YF6bq/uiUgbgt1YSViQ1bb/wtQ
2zTVYekcdModqaT4zbjEA70pX2K9JXiztHBcWVJRyX5ya0T2KQI75LRbLD9amxOP
luExlYsOemTjFboARGuT7KdR421hhmuabfFVeADO2sTkkbxHyPo6CvvAEtWHH0F2
ZQWO/0bd0/hHi7D0WnjpMBpoK4A2PMKhNc2N1GLp9QeF4IAdAa5xy/6PvRuN/PUX
et7pWSe/AQ9lv69WhRgLTm3ZVXGnDdr06iSXNTTvzVNQrETM3dyM9IH+E0g3HJNv
3A9NbLkbhqaZ6xBAVKkDg/y1Ia0UdWg8kQ7MOSI+1FNBfpLBIldYkjRrUysSFp7s
LHMTLKiICURUOlF8t2Bd+z407Jr7j6hVVx8AHkXKV7TI7JAqcxCre5fLpEKrmVT+
h5jhaLXXKxC+eb2BNu60MT7oX5jtU4pktLcfBZb8XsF8YEu77wFdD60nxbHSrswh
cjMsYQ3CLQd+KkgUh7jZMPSUQsvdakIYzsPKr6K2coRrqxSd5dIgY9QUUU+7LpID
UkMJGKj5a73em7jBIwvfR7mRrRzmEG2VIxE7OAqXs3fV6tJ9hcqEMx0cDONvV1wM
Xs6t4Hc1N7Zv98zHFJyLSClr6Q4IynYj8JvmKHDAj6X43ka9HXcKTuWiH2cJNbFV
zRcM8GuiRCmNNhkLxnxJoAni++hTEmiXDLgTeMupDL4LUSD5jgmpBOoOQdG+rdDl
E7QDyIhXiLMnK7gUFuQIwpBNYE9swpiSWw0UkX+1gLW39zu0dYgDeSYbEJ3pfS5L
3CVprln4HJ7bBZ27+snx9DaAndBtPiotMmPEsrkV2jaTmYjYiV0jIpb5rcNoqnfQ
0D51jUIo3pkw9SC0mX5WPF2Iwv+ma+tRF6+8D+gRUlgGTgrFzRPN7Q/CypiM8+Dj
1gtJcyd2b44n9TGtiBT0xj85rRq6IawvVX9NhtQqUCci4n+rCJIL/2jZr+CNhFqL
3DIZLxF845athWWFkmel7rPF7sTx7Fpq1Rf7BM+9jrBGVao7NuQ762qgEZLbsvzW
gdobSEN2/hTRvsPFLMbp6u6Z9qy5SbQzZa1sb0QotMQ4JENQIq2CPJr3aVI2Azqe
jsfTKLCUKIgsZZ+vJiiCS0RfWvNLJBKUoq2WRwATNp+/l113WcY/zaYMM0JYds/I
dATQ05QHVjVqd6DjOuecknRAuPSQXbTrVBuUEibcqyntfNlDSjjXl3SkC9vHwPuh
QRuAWvTThpCvVdEoKBXIhANStvQaSug7K3MQ8sLfkPC6PegLAq60R/bnwbB11teN
MG0DzHf+ByQ4jX+Desq6w4hoqWUXcEfEfZocvYXUvWlOUFc3Q9jkCQIusqLuqcWo
z5xMknPzCU9BCx6QQx6X1676Ki8uRveu1NZt4PPrwzbECkM6B7/+sNyZALiEskzY
h4Q6370ou0e95GhbVolLPWniKiirTq7EemnbaklbvRoynUGSPf1Wqr8luuWErH0O
4/XEQz4IRXYS+hSP4D4BQx4FKTAS7V4u1qBZFQEYSVIfCPYThobfPlq/LxSgrHfb
5cdmWHf78vVFDq2T3DIE/7E3CrgzabiRYbJLwkEedc4KNMV7dPhjgVhHmSeEtZfF
nbNkrMXFnQTszARTF50fT7a5AV5KKczxpboSXxMkfFNqf9cUCsH3g5YiwhwZRveo
t8su7ljdI4Dl3CuoRd7BY6W0UFKTlIQdqY7E7tcxG+Cul7HNY5XjDIKoeM/0y0I0
f+rpXiuTYZdFYcI/4g0VNX7Cj9qjzn9taHMq8bdkKmjQZJ5OSsvrO9ULywoa/cPr
+Y5k0ehgUNfb93JMmv3QZsuvIO1WsRNuqRvYokwYTAbp0rrqUElgZlXaA6DW0KpP
xx38+h0QL2KvpXJ21YxoR/51EZ4NDtNCZZUPAkydw+YPYwIE/WNWTEB2T605yBM2
NjQTf2TNQytpPXpw5BkblOTIrgG7sgizmvbFHQ2cQlIbFdMQ74l54aPXHBGbA0xH
SPx2WMszvs2bMJzCIa404gbMvFQbTbohsUsYUF62vDvORGGNhjrmBNIyj1PlIRxg
cR+tdnqS2KrxMwwVCXDjnpe3REBD0Xc6hcMLaaRmUK7stHjmEioalVWtZkuMZ9GJ
E/MOkh2LbDYwzZY1wN8Y6TkZF/7mmaSw9SycPF+rxntbeeiMasMkmHUOQyir/JjM
npc95v3dJlOPFckxnU2lNgP37KwdWWddXH+sP6X1quOPIqvSrtspFqEhHA4MGIYA
7ZAVTFFVUcU/ArxPfeeeOu1s+0xeKadhEfsrZfBo6XUHwpGQ9/myqOWMsXPK6ONy
9sNHOBtqxM7866DNQxrwL5d2pLR1E5kUs3L5eVkFZo4sczc+rDOkuojZ0knJLSA0
sCstQ7gfehs/ftA/qBIl1BvCD8PRCPyMfW0eaxTS2veJU4pXcceUJRazzoIAFjX2
SmfgKIUO+DWVnXLVAMkMhclhM+rcG4vFgYp6Rz83sGiI8bnvY24AGa7ohRCxifm9
HU6F+xaHH039jUYrXU+lxzFlHhAFC+Eq7HmsZCUNDPRDS187B8KtF/nUP8+Mu0W7
EsTLqjQh4lY8oHvo/84iAK1ptUYMA3mlRoAUjnk9fZ3SE/aHGxloI/m55dkcRdtN
7Uiz+DsDR/fN1OClqW6AOW1mpxgZeh9c2nAw6LvAuwcFAx5vSLAgeSvQ4P5Dybkw
/KA78iL1NAQG2ax6M23m9eJLcN8CEigtBckFj92rTJJyD/+BsDgPAE/YWrFNTvyg
qOkrnHXfl855PdDujJijinsjV/mDjMud8UEbUJDzN3/aElzL7V4UfpUrmZ040Oy1
unTkB6M7UFHanbMa/22TVBalBwYgCPSvS57gU+jioOAMcn0c+x7AK5OnJGSScddp
l6wWxutO4/0Yv1F7O/3tJq7/YMMvrfbeYH2WJfY7VM7KasxOllhMIEB4a/bOieQY
M0lLbfhFWS8MQc8U3MXnZFtFrXU3RRVhJR+/jtif6DYYnDbOFbapBQ9vQNBofZHt
QxUSGFEhjUM8UFW116drww==
`protect END_PROTECTED
