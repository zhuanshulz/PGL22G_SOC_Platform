`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yAfu8NSdRv4Cma82uN7/+uAkvwAh5mCQd+LtAM0ov5bATjtZuQZ9zpwQeD0k3TZU
pBPBhCwX7pCVZiybFI2RTos17JE3VFuD9SO85NfFlsPzp0TyjXfL6hjb/FnOZwWG
iigB1+FJWeFv700qYDU1OhIrB4OwOMFFOw4qcTc08MY2uPYrjcZ6xqn/mXE7uJ9r
PWU+GuJb6+fH0bAMVRqyyuw/gODnDoRdP/eq/xcBxlRq+e+SC2nk82hXXNoeTZSX
/Zijxm3E2h+vo5hZV55NqpGRit7DxykvtvMoMxr6gTqMyR3zYmATdbWuxrhsvGiN
KcUYptvU+PvXZ9MDYm7Q+9OhhsCFmRWOjagBM+447rtxZOH310HiCrr2dZ6KgUJL
wMnQa1OC0C0lTsbbWcnLmDZQRnNP1JyHyOaWL+KryB763yt1nIwPEbN75MmNGL0Q
NArEFyymvr82278qO9K53Tx71vAGPlKwVD9B7K00gEIZ6ABycakgCbD6f2P0oHNg
pv/37nHknJU7uJz7262VnuaNvHhXKJsSFMgGf4XI+pgC5puXH893c4atvwbjmDOl
iFvn0mAEaw1KhVBOYutsSMlSiN+hle/tYW903JP75S/ShjugNmWgU1F3kEcQhd02
9RrqHoKuEAQJqP6/kYkfJIh2spcGt1TD4qnSywtw0Gt42pZBKMpCZQ+jiw46ZFb1
YEjJD1gMKmDDLTLIAeM8gA==
`protect END_PROTECTED
