`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uXZy+RC+9Q/ZB/KP/iY3+MDRuN33Fi/mA8/UHdY/glo+hBTPK30E5SQJoxIrUUN5
TmdfBnQ4Aw2owRXGYMVa6GQ6ZFZs6reJcKQlExnkkNmgnNIL12OEIwEK8ICh0ekf
mhwubVgDl2F5tH8wzJwVQEXM1wNMJo2W7hZgsrtv2UweLePsDzlSfHeMgi+dnzRq
rQvASki2LK+Cjb78VstXPbGJrBUWd39MTBQoQUiO5fhLCQ9Y4kDikK+I/C9vzq+z
RO/xrnJF1TdVZgi1H+34ZPmDoGa1xpW+9HmXTlt25KDJDCw6Nki9dyst3WS+cOuO
MESjU7lt0/+FnNLjqRt1XmqnGf3CfBisOV7mB+IaueaH1Lpg3Bo6R3EBgr3hXC6m
cpGaCgGrDtNwGpft2FO+EDQV9Dq7+rZl54lrrU1mrPdRqdxx2qibox4tghI7XuAQ
6Km/APWsYRC2YrB7GkSRhi4AJgDaS9BX+OA+/xv0OPgCIb9wXihnrpriZwZ1ojIz
L8ChbzQgf3RB4kVySd/BuqOP0aUjxtpIXwTT399gM0KPS8IMldXC2L7WS5EsM4AU
dqlBb/Tzm5xt1ClqYGHEjl1WVIR14S/P1DK/VnQb0xg4cmVjtt7rijEBe1S2IexH
MZt9Ww9uxbuyuq/22oEdWoU+tHG66ChQjzZZRQyGdWmoKxhmppVBhcrXH3/eezDR
ezy7TOGTdUUw+RgeRgOdghRXn7kmI+WM4r7cqJn7xrthuu4O2BKucdq9wcVzsput
I3KPeSZiu5LD0NuURXcpJ+uDyFaEKQzUBDFCO8VK8eF0seoBW7slwOqDsINkIVwN
808np1v7vbPo+zoHtYaeopDWfdRuX1iCh12C7LDCURO8Yx11rkSrEsc3HXIIZXov
z1uWD3V78sulsnTNH9+DJWuMnGL9kqLAUwcASuN7TQbKocfBa3YqjhYbzfGeHYO1
fwrj1DDv5BBSNziAYVTD3yjhbUXiNHtE6fxrVFUEEgjaXBVgrzB2n0nEHggan/X6
deUVocmRuk7s74XXHd1FG7SHlcLS1GuSE5UrnpJnCplKjCRdbAEArhTnPpIzk3UU
hW2cfLAhhPCTjC7IK3rEYPdByC/4mnHlu8bz/ONqxssc1bas04Dhgsd2RH75pFSy
ID0rv+QpnVqea1z6cG6bng==
`protect END_PROTECTED
