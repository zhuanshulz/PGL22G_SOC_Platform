`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WrJZQiCRgNT03UEnoLmU9xHBqI3ValHiRwuGJksg7NHlAyJdQXSZhQxg8LB7gQ9w
NUNGTQINU8ChqJ/8GVv0tbcboMB8QG+4x/B9DoeW1NWANTp0NpsJ9tBwmC7IOZoK
+1w187de1xsySWQUhiHQXVJFO8kRq8xdcWB9hGS3jSDXmB5J8RvC2RXeNozp4PIl
cUCfYFxYoX90GZ9LAk06XzV6KRLrCq7ZztFlEUTCF46DtY8v4XBNT7577CH4AH+U
Z6iLI/94CcTyiYj3k3gwjvHk1JqnSGGpno0sqZmeeaD5zR/EpzjkwBfskQqqks5v
CFS+CYsU3CXlMHL8AmZTkkn3VPdZv/9hiPkPjeWab5JhDT9USVrCvch9lWEfpTe/
IUSMSNsf6LydRjI1/L6LwdJdHpk4BgoRt4RV3VOZOrj8xNKGDGijOtmLAVNs4qQ8
b+vhlGF/RgGd41YtYBMgDb2jvm27eETVkiL2t9Ixv8b+dMIsTPTObGCzSX9mPleO
QkIWf5zUcQ5pUENH1F99ox7mKlI43P/ljLS+l8XRtqLU5/epPVpLia5t0IV8TL2k
xpVW5sgATywz+fVimQYQkjDgsOLuF4Qd/J6dHEH9O+78ISb/D5ThhwgLH/sAW64r
+TgKiWyEQ26e4d2PRee+6WZG9Ua50V08Ae39sg6fT5IPoR8U9Jp8uVhz6p0Q5Vuf
Q5fd78TdAb/ZzShHiic6ji3/LU3KwUw+E70fwnK9euRGYkQOHJEbjQ2oPntENSOZ
1WqaVtfKc4NaHMOw7KH6oq8M+0eXBwTCW29dcUE4o4gS4sRpZJjjqoBBR7f+Vqv+
XhkjtUaQEsxzIe9twiF6F/MFgwvZ77hl1BdUJ7tHVhobX46OWmkMw0P1yBZQUIVs
aGd9hi7J+L/uXT+XUgn4+fSc4hFkbdv40t1B0n/R0ZztD7NbyyYB4QtN9VH9FW7C
369LSiNPf9pgszDHTTueAlXAz5S5OUC82doEmMCIQLrFHRruYjdAJgnqyCNVWkLw
nz/LK64tFekFT/BGOtzp9eUvlhAsHAg5PbBab/yJHQfpO1RDsycws5Ov8hpIO6j3
rpF2b49l14uahRG8w4TbnOJ00eicj5MJLxmT0CYI82YxEYjdXUcWzXFdaIJMfaMT
4hjivihGmI76HL3aB4ANCpRjpJv/HzfC/H47uMRtmhl+dWoqDVluQuD05W07Db/Y
3nrSEVlrHBxVrkqovXFxHv2S3EqezaxcQGsEqVkWdU/yatsOkowDGHFeZSRvIx8q
ybVFOhnNz4NUQpdsY1OlrCQX1T7rO9Eh3nNbjCr0Qu4oSTihxMEdJkZ/DvAYTO4Q
AddZmukrOZJtGFrKyFZZbwSq8wOT72rduwdiMt9EcQHBIibIAxHgwEf4LI/Uy3ii
2CrgX1N4BKBo9s2ixus8Pl1gVha4VYNJttb2BnaQrjfx3MDxwKDCajYOzj8PrlNl
+VzYOWvl/pg/2Xl12L8tko86JTzJuUuKfdtgUTQryUYKzltUFNM5XQ7DzD5ArCsE
XsPHtm3U7wQXkgCss9W5H5ptXdBGxnm+FDV8+e57etM4DXomVhNdUo4WnjP3lZTj
8M3wcd2L0SHrIu9p9M18U2e/pS5o0OgHGjwPmW2aX0U//ybbmskxetZ+s7kIULxq
ejzPp4D1W+KVcIiIs/zGJbRkFy8gvRhLfl1pLL63yWvppnedNLDyDfc5z1SZkxLh
acRsQeHQ3XsewMIOqq5CIgeC2ZKwyoaxu8lu0lbq3gno+dhNvu6yfu994MbEuDP8
0eK1iCeK/4VCmKk1YFnIqKGmDHx5n4e1gSQT2X7L0TTUUZQI2a7NdM6BVFXz4fp0
dHp5rwRtJFm7GoPb1Pq419SeAFG7hw/pZkNICGu1O/XU6fXwrayzpxfS/3PWhUYQ
VBy32gh9Fk6/Ai774C5uB9EhKhCfrW2GFBg51+eJgR/wLfX6uKwGZZ+Pj0RTs1vF
iX69MI/04QgtyGmvnljeRYQEsVDM5BpURGXZO7TUuDoTj/ctZJW+Yxs4Xp1u80ar
dygfVPGo9+U6Q7CVXxqmwpWKNWLyiPsFLq/JiUBK4pgfhdcrnhIjDyyLWvF59K9m
ikvuqyGn+2pg4BBiwJ6m9Oy3RIfoGF35wPbz02GpzEEY4Dcwp/otYhibut86H8Fd
bSvudG/A9zUSg6WLLGdJqWpJ+IQ5Fp0K4tVZXTGvbNs8JLgM4B9cq9p3RcCYvucN
Ux9SHAIU8QHtPXB5LXXZIT7WcC78R8UciyTe3a34OnKYKKre5M/YdG4JSOKqwoYa
KtHAs2SJ2XSbwVwYYd43LcZYy2ifBpJxPvPGi71ZZfDmGLah1C2Bbyiln85VSdHS
8lmZwwr1Hzr9o9WaY822hzArvNy0qC/Hx5bgBoecwsRDQp9SIYTdGkRr5sMTQtTu
JPqXizPGtzT3CgpmrsQogxpZj57E3qd8EYOgAC3JOE8ARKmBaQKI7i/LFqnybu8a
8qkx0xMH9nwah1jZxUhE3TfB6V0AbcrbSXdsCwWPDY15igBg261GCXDLccDVnaHY
CUBnA4nKpJF7vL5QYdlpazgM2aSyGqdGPPiLAQgjKJxtAlGe4Pa9MNWppEj9KzDm
3Ba/aQr96cPgTfG8HdwtIwP1tW3DC1MKiF+oC39ZUTT9hratskDxsJLuDsQtwQCn
5rmeNS60PHdUXK8JnqJetto+ugerBocqDp/8AJDSPNaygC9HUDwJdmWmw7VxtIrC
jaVKyH5THGbEt0NTjZGC3X/RARUgDY+UcpkbwPb4qyBnMgrIP8xAkJ5UVRUbcp+i
QxiS60YXQYTbDtggNrBUSziFvdCC+FGU8hV3nuNSxheyyawP31yY92xIlvibIXcH
ZvyAil5WV8Qo7o/uGA6yLYBjtZmuheztuGVOmEQpdJr0GWoR0MJn9bmSL1ILaJsu
Eo7AMiBGfHAKoYhTMYprpOCnEC4LlqThjDTcInOyMB8/CVVK7Lc1tyMVCNz5ImA9
9Bbcw2UiNrmoFnD9b9kq2h/BmS36Xozvm5Ts7OoRRL858TPyxSrnQYSDtILidOG+
3vi+YQMjVO/Y4ZMUwdiTQELJciCOCMxCrwf4tuM21jyhdWne+1GwMumdD9AJkT3f
uNAgNEydMNV4UsXIVscB9BLB/YjkzUA1tIFl4jj2KXnI06+Xu/35aZDiqEMqsjfk
n/4GaEjkbChXZjrrAUBxUJTFP66DI3E2dIa+wVYyHCmjipGkLDuVwPD4V8L4G0FZ
3ZGferbTW2GDqiRKV4Ne5wSif6+zpEa7XFj0XCJPDQ8WV+aT8I7ILThzuqqUr8hP
j3OyRXUHQrgmFOVbYvXMb+NS3538GlWBtrMEr3rP4aQlp8w/itTn7oQ9Ap8te5tK
BgzvMmNKTNMyCBMBL84B/5s295OpMbqTKYOwsD8g4gc3CgdmZ6MqVF78RdMhsOGz
l1lilqMG3YJMaD3MSV01/0FrXJBI5n+p+a+X0LnPvVaVK3douIrylMnelltgAoPm
c2jFb+X23bRsGAmbmYA/bCyBTw4BYswSc0l6kL4kJCfv6Dgg/jeGsTN1V9HDd55a
IDgDqpR8/Sa5Q8SuD1tq0u0ADj0xKmi9VweMk8GBXxvmghwSpzNB15QOmuWc+Uab
lDWD9l1K65i8ndXS8lQmTmFYIcY4iwUXKEHmCh6InUJws+V639xOlRhkxeMLUDwN
KymvP7474X7/pkAxGR9Ijeqs7Ny8UBrGA06GixMJ/X527IPgJPTnVozxNceDaTFU
weA38qJbDp3OFw/JQy6Xr/ujU7afZKn95EIZM63CdH8dedxLbDCjqpWlmoQGKfa2
IS75FogRBt/onIyx/PSOtq3rdvGfpFVTLAzoYy42fEwbRxvOdaOpqXoLAiXQGOfM
bR1rIDuF3lsphlvFqoJd/YR3t20YL5iYWTJ5RYSZo6bBZQeDijMcokcQdN73JMYL
VmrfPX15m/bAO0n5lWoBZ63v/0wkOhLA3rYVM5cmq171sfDF+bhLKrXBTa925OXL
yJ1k44Qub7ALzBdbX/c6k1KRIMxduPiqdv+I8Kj4uJZss3KiER5WL0EdFMuogvdL
cwyYOesTq6X71tJg9ZNUKAe/hAcPM24Ph6/ibCCxMaJMW5Uj8Upyi0uSA///d+WW
fXYfprkIjEGQkdcUNDo9qvBSkQVg4XupoJn6WEHXCvPNe47rPL8Uw59XBlfztQx7
rk5UyJ1lNXaOE4yqgzS3X1zNgBMqUbanDFpX9He1D4sszGX6KnBNxO5QRjRxFM5f
iNb/YhxUCQxkdN0Am95RfyN3Z5Z57W1RILcUrqTRkQb/BKYi3RXQrrToGiMt0sL+
k2KY9mvB0f6x0YSjCQcNhuA4OZwwl0ZFNTUIWMa5A/Xla7+BlPtfetq6t5bNXidQ
fSxLZF1v4p7FRH5GWdsfZY9LmliyEiyOBdntzLRhS/oPNI1uBqKZ0RE1Exd7EDnK
LOnigg9x1l6j2MphrU2HLxWc3JM1yzATzu892b5qPpyuG6k74CaYO5WCfNk9Q+SE
+ck4hishdKbSnVsU/UgGlfMaSQ9T3Gj5P0ObateOLZw=
`protect END_PROTECTED
