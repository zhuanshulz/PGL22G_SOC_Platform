`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U11tQqv+yN9ogNXCnfPmgNTo3uBsDXOkxAy3V9fjXi5ddtTKYOrjayPTF0dfeq3Z
a0sP/hG8AmQLvHSS7pZo3TGE3vUu0z2z5OO4cQ7GhM2L6626av9AdClySInCVvH+
iW4XA+L11ZkpxCdQ9qeHn9HvsTfWlEwqqdpKYbo0Q8ZheWIxadrgjhU2w8adqRKN
58a55vl0k1dbsSl3tb/r+mWpQd4Lwn/CCxIQK6DwKvdOFkFr0G2+H9dyyB++ZHhZ
OQcFBpkIhgLtJ/CBbcPExn+81r0EhmHHlcYFNirylN2Gy8xaE9u8Zd3mVkWqSN4i
lE4L0ePvycCJZdQLtR9BeMXJGldFfY9RlKCyRdTOQs8vk67fXbldLV6BJG24wyVk
EHptAwXShCsFihM+xpdA+DZKQ9e+AiuZ/2UdhAbM6FgYLT6Uq1KwHMCMKafycCCQ
oZzDfysoZW0GKxMFRcXrMgQ2xkCFcVbRLwJo29yZxnPC/+ax3qWx31LMrqILm6Y5
OKebff4u1Noq5mJb2aDtvvFfCur5j/mqRtelw8rqPWc9azlPvLGH1Vfz0OJo59Sc
k1cqL+Rlk+CcpQfNhx0x16LAgQ3qvIeB1UzzzBDeX5bw2sLRa71L1qRoMIrPtzFZ
kTgEu1o9NUORbxGrz2Eb0bjSBI0H6J+g0KaCzwJba7oX64cd4mUiePjPgTA3CSGY
6SwtKg+0kL5+Xz2APWr4uQQVnK59Z5wWwncXi9RtUzcOhELVvLHQ+W//1lki0P/i
5IloAUvaY7rv7rmlTiq2iCuEhMSYC2JiU1ZwQbCx4fdKY2lFKlN313/6oFKNqqMe
wJY9VsO+J5Hnpe8fu2KrCUDRFb037CCJzl+HLfTh2UgyM4HJI7C2baScXlQu20pH
`protect END_PROTECTED
