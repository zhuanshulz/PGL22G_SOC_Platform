`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2SDE2oOJAN6SqVUWq6L9Julfjj/ENfUsCcuHuKnLcX/xb5vqqQtd1OVZnrbLkesV
48fe9uqxSoXuEsgXUfY619rDBwzDz/uaQ5nhSo5cGt1NJJNYTEvc5AnDdX6poFCS
EEQvQ17cW2CE35mIOdAvEN6n0D3Zg3fC0JNK8rMhTUcObfrGxwq3pZL19D8F+Now
3jiuSHYLI49YeDBKvNdipZI9O6+phPsp5fk6vYkY03I7zWo7GfbxOV5H/ng4ikJN
hnxjKbb1mrm5RL3DqduYVQUs+cNWka90mjcSdYBG9+3DNEXVbeRzvcg8otyuNKWY
BAj/ePSrKlpCWfnzf2J1VytmkgnDZZAJ64VHQvpqLvN5E0Lcz5hpm6vxWwC6UhPB
CmOeru0GOw+eqvwsqNmdUH5hkNT7n4+dv/kEMu8DvULA6CQvMvRmsIU7yGTE0DFV
YIsH+eAxcPAljtcsqe0YHLB9Vn17IHIe5DX3RYVvXwGplyv3SsLPcx1yFdKgPbL0
BM8MuRT4PRIggFF2U7s7CE3fgymjrtZEEk8B9F9hAL5bFW847A2eMLiK4FsHvCAf
58YNaz8qTW5+Aoe0o7FEZrPOLGdBrQPEumyowzR6cl6hDz9QUazGTpzkok0kgdZ/
yarufs7rCJTDpNVcdNJauR8LNv9dMuT94bsFroeYPF7/ZkYmVtYWZY1i9zURsgkt
5LUl42DO8f6hg9tGTZfzUFa2K8vU4rN5lq8YYTOfu//lFjSmYt9zu6AiFKxFZb0N
+3IW8Tg7lwqfw4MDdCGJnxQqay6eNjMukOfbAaG2qurwzMW6S+8oe6z7RLeK4fRs
KcWJxYcyTzB1f9QXo823W2nf4ahejqlpl5bE0jyj0iBck0jwtijchG3/cuixtFZS
kuP3XGesMkpVVLY/ikiZ8EfhH+nFlrFcrawjLJEBRo62fyItSR3WY6WdbCP2oBK1
wRMKTxcOS2fHcJLoA0maX1f1Fr12z/PjpsiY1bLZpSp1wUqM++PE6Gdwu0tVieZi
dbReUuHmCU+IzvhAzSyUt7h1W/0LBVGaf1e8tBIfOUYz6fdBTK0K7dCD8nfIkvwU
j+9EyeRhaTHl1JG89Cj3qvqDME5+wG45Mm8mBMKinA1uk23ClVH9Xag9V8cuDLAu
MPK30HqkUyASgMW0eQSXLE2fdwnzVSjzQFTxJUHOvwzRxXIoYANb6zidGh0UI9xX
qIcKLhSz/o7BBzcF4SVdDPNVWnVMY0m5ETKFgboR/x6RtfbLKuIHwQNf3SH3C+4M
FSiUOyU+axCGNoJe+nMesRWou2ejvIl0TppG0OTKPvabgSkGo/BaWOBz92IBxvej
Th3CYY0kaZGoRLtJ0q9zjzNQf8tTvq6EudbRe2kg0ZIuB3Zmw8KnPQAb0p8DZcGJ
Zo3pIBvamZXpEHBxEzNBnXGOHi/RgS84cF7QvVRecILh74i1ODA82WGtvRC0DgPk
VortTjpAD8wHGy6wIWeOqyTbU1XvsVLj+GsD9n33N3H4RvzX2fl2r1DxdBVGdjgB
5dEXJ6twavN8GN/56WPeo3E1i6ez/DFtiwkEOwB5c9so6Vvy331rtj0yAX8pDFdi
raglko2O42WW7QmFAbUK/QI8357TTCdxImwUdYP8YaARhNLraieLUr/LO87+XLRq
4iLwKYSleDZ/0osQXzHS1WDoEUUR2P0r4CSOQE27OLsAjTz58u1p1bfg8e+MPk4F
e6x1uplrwgXIVp/RleVYXV6am6yEJ+NHXsEHYid1UyHuAR8X6vzhpWgR2hb6GTfM
jIsygw8mvhBtCPQ/r/c1ogKUaBu8SfQXycEsTNdc1nQ1RugalUl9B5Vo7bJh6joX
Tte1PYm0p0OTrSHZ89CIh+SLwZhxaMhM8SsSoESlzW4K91FtXd76twMMGO5TmfzQ
xlL5wjzQCju9lMQpMuMqpKURNGKOh7jdqgWD9G8v9ulbLViQkaQwqMYunTQXsjxf
zb8OjmV4VSayRGVi79K61KORpFk/nPLfvfTyNdlTqvxigOLZ6g7Bno5NeRkYm2IS
r5uC46AnDPyM4oeecoFare5jTpvV8x6IsWT8V1qfNbJ41Nd06QEWuiGV6kPbbOpo
70dVj0a+sri8guWYhMLRAb/TIseU2ovcSafCoZyG/0GH1glOzcsNlmWgr4X733M/
ADlC1hnbXIer0ASGPJsyBa3+D8fu7xAqWvLB/PskTJKwuN8C+56VOCVYNcAFzh0C
NiQHwMPnv9RBOVjHP1+lhfEgaHovUkF8poqQUf6Oh0Up9zaLIfx1uuDtPpdKpERV
57UAHBmGZ/AgVGgd28HNH5SMVqYnf+kiEUwEq3Hi6EdWYrDeNEYznJwRPPwbzhAd
e+Y2X3++Ho6RGwK8JcXtWej3gCrTyuoWHmukViOsXvXEUADIrG1zJik4FEEcT5XD
OcGKQ4GDXRuAcAKa9eQIQ2HcnS8zju00TV2n8sKK31cAWtd+ykQxZpHuk34qbkYm
hwdFntPjdfk1RQFShx0E1fARtiTKgIHUiUJVTlb6vDU9sx40sarib5StY6lvIG42
VqEmpVKWiAw5/4kGEIW7exMnjiJZkCzaCMgYPdEhL5aFp37GOwEZf0d1FFGQEXs/
8dNGHUMA5x+4ZS7dxczAj68WMMagXWCbrte/6JePbNmB4mw110otkmkcJRVKIS23
sErlYoLFHuC3XyqXk0hWtNBkClLENajQGk1eI02cX5OFE2PguGQuGc7Gpfdiuj2q
ib76Odc5OXcjytmKqRfqe6eNPThwpdGcZM6/yoJxFPhfFTGnNLho+0iA3F1o0wLU
s7YEVIhacybw0kRMLbkRbHlpC42YcJrVw0WfA3+pORu+Pf63pFH8rRjei/uuxtno
CnHElR/T2SYdMsSq02k6isGzHzBrD+LgzlRZseyIm4ysqRHKW1kd/FEXYMR7j0bM
r38T+JDV0qT5Y9C3750i4vUOMfplcSsVE5lsYDOi0QLKpHfOxcEkhDoUm/hre2X1
RD42und5jKKiDknV9/Jc2SkwQ9HbcSOWI8qzfkp9dpcMmyshq2/BIjwpHNQeMZXn
gTTvkgH1jHhXdao1FCcnGwKqwEyA463tY1zOPQr7cmS/m760cupNw2l8NMHyFRr1
bqQRbVo810wlU0DZZwXeBtPMpi1JwfbOM+6+Ht8mXBti6dzzLCawgeRI5Fk3wcgh
uZvNWwe5ptfenGXikNw/x56Fxyr7efOb5Lz0TiMNMC2P1AnqdahHQkxI1SWCsFUQ
HhgzZ5YwAulZLvUvPK9XszhcEATiUj7Xdh305qH3gXN2TakwGJsih7v0CDlUfzEx
sMjBe1AsgLoPeK9IdwxKzYDlvbU1ASDjZhEq0BzldeY2Z6w9FPDjpzwM8OmVfzGF
jE++UKB0EZiLsv3OgkRnn60TwnE8rgZcXUrbp3SD6BsWG5zp42uUpEecG9OjoICP
tlCc0qirHuhoCm6WUiVixQuDFfeB//D1dKXfbYhYpNfGPj4FcsjXtVIGvyg/nsTP
HhqoGsUzaaSg+7ZCstTlTVtl8PWYHqnHmTfpG5omnEI1eQVQ1RCCwxFMSdzbCiK2
BzrSn8/B6nmoo4bSWL0Cry3D+I6OhYDbDY+FvP/xKRZDecah9nW/+cP4YEXXkpAv
GgRFa+R4dpdXLMyStrBeDw941+29mdD/P5AqoAQoxz/GV6aK0GQ7F0qI2Oi4/5Hn
VZwucXlWyusk1eJkd3vK7EmUygtpYJkwUJ7bdzMhVL/5MsaXoUJRBkNnpNYR5AdX
Zw/yFmJ7BD4UbzxPzv+3KZVQcKnOTb43zi2Oc7yrBTWmD/THt8yXTeISTHKal3wO
OvwlKmEPUAZD2uO3BV0fztZT4wtldL6F1c+bWB8GXsJtZewBk/ZvML12kt+ddtx9
2o5QcszpTta2VsFcf47yhP8HnNN5ISGLTHwStCxEDqWUTv33Wlud5wCVrY74WmL/
f01oqPeBOokm4xj7+B2O1VTRrX5j/YkZTu2DoqCP+OKhUQi/bTjxzplxr5LA1Jbb
Z3hhBWnQKMRfnfap42i3drFHtlC/UO23GNT55nZbNE4nsCu++qGgjk5AlmjOvhVd
fxGK5rKqJR97+hS1BuDuQARwnU0WvsEcylyLmx2mT52LkJuxSniJxbGe8aTBg9Fe
FfTZ6siuIj3AArDa0QH1javL+6WqfebTYHBwHVE88VOLdwVMQzhyWqqXkmV3FIhi
A7RxlIruvwmokF4DMS/Xuqmr7e5LeiCzEh+7n2LZZwa9Vkq3USCLvvCWtBo4c+/c
ImDALalf4ezy3elPYfV233crnu7FWIt76++weEpKcMvXX6WZDkwC+lC788g49oYK
mrCB8rzFmbzdAqYFvLCksJjDi4/GCardpOhpxuo8K0YJsiJhG8xAO3Fvtc63UBa9
ba+7lCcz1NY5/IMe32NbVRFGGKS+AII+m3LJPPsigSJAPJzUU3O7oQzlqTGqCN6A
AWTZsdDvqGXBCxxhD5PkgO8r5CED9Wumf45ANywqSb7r2ofdR93WCkE+MkdxAPbh
nfbdD30EL2gufAA5pwDvrd+Xp7ZnrAvEBYASmNsgHAH/h/4OE4IRUC0zhV+9zAGX
hW2BhZ5+DaYcxrBtFS8I5/krTrQxD1SOHYCxwGn7lzIV3WjV/8YNUf86iv1ZFSES
IsDvHHyFgvIavQUMA3ObNKviZqVkgpAEHw2hfcyjLNsKCDgD8uCNa6Na9cz9pIuP
yaiHBq2bUn2rkR72oJDEyLh9xYpHr1lKQoliazQyPkFrvJU8ymj2QrPQWc98tTDN
A7K6xJBcysFdlg0MQp0KiiR8sQo8BFZy0n2AvJThr3zpXnhrEVy6Wa24kfcfwKbA
X4u9QROTA/aridGBKmY4CdNXqHYLnzWqqXbqCVYLHjLS33+4pFRMxf1LijSsueWK
Paf8R9JEMm0SWrnglJC6bSheXtQfXpsUgsoTbcqmslmqXoeGciGNKRjS7JbOMWU4
XYrnxp8VP7LUYHa56pUVQzdgFCgtMoqib8UyyciRFJnK7DNmP238w8eYLAvkDY/3
i9rnQUx+Va9efjXyDOS6nWOAvHaawesGgJore8nrHrB+63Lu9165LUii6g+rTJQj
BU9Gas4MK/gosku+1HbiaB3je+frjVg/eocVDCu7CyCrBTai26hnqKugZl+kbIpC
CPTKT6/jTn6iOlKT60bPEtwTzeBvhhXWytb/gR0orcjM7RA1G+qwfU5ZGqjaqMlf
W/XSa3X0U2uyvk6b9tEnmc2lvUoy3NHZ8Ll3R9OMQTLUYf4d9ncxLjJ8fgaRCdql
UBlmj9/0sfC8hQFe4in8bqMD5gRR2Ar0hhX5kVRVinlSI18p4JwYuj30YsnKVnB/
9UOb8q7Vh+CYjDC0f45Tzt7brQ32T3D3uftZ4Iha0gnsXrgECHZmuqvpQzAZbBbb
qqiSeu9pMHOMZWudZXylUFESQ1skt2gqeMBIU0rJMTBVJ3a64s5ybWtzvy5wytUc
Qz05pnrWVyRfm2Rj/VUSzDuTNUTqnogStc1aBoD9ct5RFMTYgQzq/ULehQTGaL78
jF3k53rG3iG908zdNxKO0YqflmDMUvXIS3I95yHF24qF7FDvAWaTwrA5YYE2pEYp
75JV7iUD4ubvd2kBXkXazrXwg31699pZSqJv1XQK9nSaizXWCCttmCRLyMzTUjgu
ZblaGJwW+fW4wihlI+TqcIiaPi6WXz9GJY3Kk8SlqTaF1V+kyJkJ3BW2F1z7s8Ib
Y1AoYzJUJdwTD9UK811aRAi+DgLS25rjoXZA0PjH84lD2UIfmGSNtJeZS1oSlTHJ
mFDmFYKlILx85httlGgnzGbtbzRKkQRh4bKKBB8drxcFsvIWwR4yKjaqK3mpW6XI
VGEu+7hdVO3WZjA6C5plI9HXyKLCldnN+0GeQF++4ARHV9OD6/mxudbuQ1RVi38W
GcSn+dDru2D8jDHEG3KOPgBFPjzS00ppECCjDZGrGVSoLFuu0nc2kG51wYxhIBSM
hasG8K2GVVztUo+kegkvWeZVb28OcvsivCNr4EKucM0yA4XH0kHF04BSwfoG3ljX
Ysiqq6e/cxjkAhv5pil5zqB/r4ezLaC+sBKen19PztOIFSTekqk39Ps+RRK66DE7
SYQ70IKW7OKJ3Tdz/HusJhE+hsF0PiC9rjn1OB7Mq3uF7VjXH7HT3dvOfIFI7t+V
qeVuYm4QuOGwGOuEoe14RRKDoF/3sHOIWebDWOb4WFvRNx50v/g+hbcFtvmUFdKU
01x5ZFINu7zbYqRluKz3ExqHIHUP3FIMDxZaHVSQSFxbdtoVIWFzq65opZe0C4bP
YUnzTZlb6K19Kn4I9dd+ranNK6M6qNoL7co7KyVoBLguzdnGK/yT+wrkJFSsQa09
O8U53TUJ3xjcDdX8EGtfO+Xigxq3tDIthH0vxbqVg1GxbZeGjIUKuykTHH5igOoR
4Bfo6CZcbSGd7pbTDMvthGP1w7/6ipbCbhftUoLrJawiNkWRpnvNz34n5srsLhJ+
Dx0fpaq/KXTy0HnQGXUnwyP6o4eg4PXw4bH4JazMHDuQ5Hxr/kld2+wI/mOa5WtM
T9nBPCdSXSnui9wltzolKYYKQej1DRQpZJQ6wVDhaW53roj1y98oFlbY2vkY0NmZ
aTn9FrQ8zpvBAOU7iWCQ3lQ0f2BJKRUV+8GPKu8cwAjYCmcym+fTY/ZSFYjLeLCJ
f+365fRNn/l24PCNajsxcI6tE4Y6LYdVAiZ+PQ/rv2V3BDKXaAl2EBem+3jlbfmT
JioPUuC36Xoas/WE1mjShyrae/TBgCYKMsmVla4UdAgKWAgoi9HZqHGjiORtr1sJ
Df9Bi2i+Fq+jtd+YfIMItLToTALbUDCcU0uoJY7R++mjMtrFkfI8vzRNff/fcqA3
XXS6jCylcCE1M0PbvXIBwDozmWs33zS6LpXGrblt0SDJyd8w+Ko/wUL4EFZGdkaD
7UztTrN0frc+DhWumlKtwSu2oWrK4GupdqyLWO+IuoJ+cmuM3FBJgECwaDcCCGF3
8TePQdTL2UShiJjRklOkSK7tB026ujaJ2JxcPrYgyIhQRV0eBk1HtDBMkTaSrI2v
CoSQ2zoS39/nAVg99uccFIRaWaz2sriGO55wS3Grof5xAZv1ehR5PqbujPLWUT7l
wWJguNWpHXU9rOUg10Krj/GFzbpCorb/WzO/R0zgmf+q9ykYdKUHjBGUuAf4OS6E
cIIyE4KyNLTjKC6tM0JEV7dNXPjYWWL5p59RhbmU3QXcaui0FHqMxSUlMUNCtuJS
o/GVd/mL5J53PwA4ENjKvQePoXdnlQewidxFGes7Z7XVT7aYMyoXKsODt4T+IyKk
PqSPGJ6IK0PXkU+XBJuoc5zWoizRL1GOCyTy5AQNHvV/abpwtwAJZNM+73o+J8r/
cMxjMqufpAINbcemuR2zT5++ZOXREbmwET8J+0v4voAyIoUqByQ4PicmsxWlkztK
dCeKewMUnc482JY6uxriR235ySRPpDWM/ox6O6Ys8CdPB9gkM03uac+TZi3o6Vi+
8b710wyqsxxqjzlX97u9mLmPEG/C/hpaeCTXFc2LJnEOebqE3PM95/fn2YI03dWA
Ps6Rw67d6KVj8412N60ZQEbr7PGmB8KLDZ5/AZEnPR8qC+oasnYeuPqwZj4PrhkO
qGnFaGrL7nnLwt3V5VCCsfWuIKLL7GTIdIDSUrTIiPMC6U5crS/0oC5bi1wbCck2
6GixpXCwJaC5QfJNbn2hMKqWkDYk+BSbEzDmDmogeyU=
`protect END_PROTECTED
