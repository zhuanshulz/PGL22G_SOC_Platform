`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EQwQjHBGY8wKN0C8jDSIteng+NU+y9Mmsv3WuMBO7SKYsMmJDYAlC2aFarKNklQu
/2VvmGTcwquUrdWFMN70+oIGvzeev3FyLVkXAVxixlZJOG+EdAhg1xEPndf+Rxah
/7i51xG8U8HIyd0wTMyvOcLf3C+gZuNaAaZ0ucL/APo19iwSCEWsT+pLgzycf8fG
AlkzjzNYNFd5adThmK+OSk5MEhDem1QFIsX04xXtx31ayKslpsmbqcHOxN0nFRAI
cGYc/81pkONPQBPcFS7myChBGCq6n1qMqXeAuqZx/FQgbHyXosng78VFiFzsHoKG
rDnzHaZMcwJo91Wqwf+7f8t7oMM4a6RrRpCR+WFQHuCkl40lXpzOVsGuBF6eLa5T
4mG0cgp+zKgmNe6YeH6H7AbaDxRrp8tsezgUldZ9KDSGEWFaMUdO4863yFvXL/yc
LhyL3yEENCHtU3yjixa5uWzj++ByLJgQhc0mFqfQk8/ta89yppFT7BOSZjl1MkTf
gqMq7oMxOOysIurNee4Jrfg3kAPtVmfH7fFfPSvV2Z63SQ4G74+09aIqXd82jzTF
zm/QEoe0zDgLeNwy9coiHxJSJhJXWgUalNp+XSUvhnhXsz8SUZjQo4ui5gpzzROo
`protect END_PROTECTED
