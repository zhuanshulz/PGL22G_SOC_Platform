library verilog;
use verilog.vl_types.all;
entity GTP_ONE is
    port(
        Z               : out    vl_logic
    );
end GTP_ONE;
