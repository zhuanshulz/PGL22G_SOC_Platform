`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DzUFwM1ytlvvd8TOz2X7yVImJDZvbWVHRGk4bmfVAtQKLG/Kn6efb/+jYXwc9lCA
1oLrrUgDtOP0CHuoUGHYcPTahcJEu8/QE2eU0JA5tHKegVoxttPjcqSsAkBsJ871
pvsgC5yl8qTOdInS5ZFa+Y3pnx5I4Mdo/f/GY/YW2Y9WduuWXTYHxnHMq49YUVbH
JlsKkBFjKnvjr7uBrcwUBVwvfHijd9oZxLgc6RYbfLcQ7tRaSC13XuozpGJdn2FW
oYx404DDv0hnj78xNYh8R1DOST7D11AR0Ta1OA2Br5gZz5ebsTR84loeRdKDWsjI
Ge16yN5pJQpzdhDE3WxL8SuUN/rrAgp9H9FvDeCMxx68eU4/+SUCWyshU+uMs0ta
wUmxyVrweX/+Vj199p4vABXlXuA6opRox998ayHgDCklNFSAukRrqMuSKuVWuDcz
ffcsFHytp5X0OLK/ZXg/8wDdGshdPGKV7JokILR0D1uyV/QgqlRfBiDlW7m8Silc
SO9trUUdcIm1/gee3ffh/VDTf8zsOFA2Z6qe9Dm1dFCa6Gx58AyKdwfWsw9j+ozJ
pO3ST6UxJVHFSVMnvYhqiQgMbSD+8cV8ve9sNNqDUQWz0EScl1Yo7H63dlJjwUCg
WFafIRcWRJxY6oqBV46uMd/ILwnASr3+TWkB2kqGJb3nVZA0+6fNf3pHAhg2Qm/E
x6T2KqkbM57D5OZaPxMRqAGEYgAAzqvk4ox8HLBbQ8hkugGbpg090YWSPI7ifKaJ
VXDOjRVGxOXMiSUvTPmwCpXyk/Iq8uNgml58ZF3ZGNM5pDnkZCf1Dn1uIUFgc4aM
IFFc0B8qvQOHZNX4vIzHWiCINDj39SIRJvMwIYe7KsFqs09jq/jgpSIwO4cB+ZFx
iU824FPUKVc7iV1qdPwRO+01/LLSmVrkVHlMunihiy2baO9C+2OhoaBkd/c2z02/
0prEIWCFTPkx4EZ3O51k2gKl6CvDe2e3udza4y+6Cg1tTz+l5Gt05iZW6xuzwD7z
WISjO64PDe55E6hEDVSZI66N/RlMjuo33aFP0dZnvPTvMgC4ioXoWEHMfJTV2k2Q
zs/RBZfdyFtlVOcJthY4uS3q/3Aw6g6MOG+KOWjffMKK2oyeETe0iWGM3AmtMQLr
8BENCog/joxJlS+GJoxo5FKbfFEcnI7QSxK67Nq77v19R44gUlZPTUeNTwn0Ouv9
TaThw08+G9xKEQxmQnG3n4BI19DvgFNWPYFWx2FWMHshLgkevyE48D1P8D+JPB9o
Tuw5ulqwCY1WnTEOWnFCMzFE5c3wluNzDvRMUcmeIKFUK/NYU1S76TXSv7PbEDjT
EjRqCb63tnHln2brYYX3Wq4B0akUsUkVOw2coE59ipLq+wRDCaAnjNq2FGYWTYSi
ePpTLltUTpSu3ApU8g5RJpCORmXpdrz1EHv5eO8S4A4dYWnxJf/xLSt9PGuV7FcH
1Ye1ApCBmSQB4GMQBGdzmKW1lx647yjgjpqSp9AQ+M02DHVPtx7rWyVMsN7B4Dy5
zOxJNnXe6GH6cW5BDtoYTOxyjbxYAbJyH01CS9AOgbvRAPKwtonbSAawmElv81Gq
+p2CcyQac4T2DX2553HJW8g1zI50apBpxrkBv5HkBpkFJSUVazzar/hJTtoDtSSn
B2sFYgWu5QyCbEWnYlvzOrBl/GjQaJpw9VGUJrYVMxyv9L59zRXjkywEUIdLoZLe
tkAt1jtgdyUfP98f7K/1NjBCilaTZc4O/IA9Z1GrcKUBEcflekNMRIBzNjgWglyU
3IuiUTVuti4ccxMQMLymRqe7Jf8pt47AN4YkgMFHrnSMNjl8w8nYrX82OYJtDldt
289OgySPfaIBnzTl82Wp5+AvUSflQs4y7RgDGT+uPIufYeQxw3eEO9ZHWrMUoZEm
rsSfPdFksJ+AIalPoiZREcT4BotB5jyQozCUKy5gc8jg+ZOSwxkdwQAYtUwyQ6P8
x63ToRGx+2qsjaCb7NRqFRa5SZuWfiMNVZvqvzdhgBBfiMylaPQHcVQFeU2rsbKy
EolTVZ4cCS0X7n5i7gU5th0IjJF+5RE7qMw9ciI55NkBoeRtcuuqz9L27ryiySkB
wGDnPyFnItDgLopi/I03iHUH7ROHbL6/QgYE3KeCLkbG70vSUw7Bt27h8aAAVr6Q
L0R+uAoJCMyx7d/XEiIj+PPRlGa3gtJlfDG5CqCfsl5h97mHbCKBF3XZL5bdXCkh
RURs205hz1Aky6hym4MJlwYe5ylhzIhCrZ06v8rnKBX6wQVHHIoaj/WYGH5L1LiC
f1bhIBtOeCVORLOY1ossUHbpCYDhT2IPujKvVy9Qfqylzm5voBqbK8lKSiJwJmZL
8NoZl9aieVXhsT4QLfPjy0FgzKJoPmG1NUyCOmn/KfrRdjQlYsHdIlhshdbhSMjx
lXW3KUMrW15TDPnFj59MRYVrR3e/Ndo8f4DLYYA+qeeQxKlL3DP9PZ2KmvL2CrT8
U/t6xLt7mowcrELWCXRZm/vMiVCOIwQZZN6RAm6xzUCKJxtM8w1qsEWRC0ZmxJej
Tw8bN2t2pv5GMx3jjOJG88lnPgLgdbGSwImXNadYEEW9LH3X+ibAUZSG/3eSqxRg
K/OH2tc7PLLB/LaFCTCVt1T4GRH5HZv6MQaV+LDSD1ayhAWmpUXsisid/0dgGRPj
6Ld5pDO432m2Cd6uIGuawUgvlJ7fQC+7daem2jWKUcCjQboEBSF6Nt3GbjUgtxjI
dP5n8LAggwQeIE3z22DxeuONbtOwKAV2nm4njNWITk/MDDb3thmxptNsECwI+yo0
ShJddaIMJ6IeJYnu+11sCh7FXSbzmhz0T5gNQDsHTrbF/2rhrF60nG+Y37NAwnYW
xK4olJR/RinRFdzdlV0KSYnX6JGRH+q/fC7pgDIajLRBvG5Ex/AiXNiCvDCmfX86
ird31fvRPCVfI5uepHPkMJ71V6sZrzBiEzc59v8PMS4ettpoGfD/bqELPDtwMMcR
xXsvBE2SY/6EiHtgI/Hu0ykE28NKg/WOe58sKat8xRPGtkH74QR/2Ho25oUUjfhG
d2PrAVZoelVCs+l851/9v9cHU1NcxKdoBWqNkAQPfvfxsLkQlS/dFtFk4v+ZV7Fy
eDScpp7RndkfLC2eufOnnJ6AVBzi4nft+QZr0f3xTj2C2xWNjdA1JF2RuawWn+UZ
/Ot9dSJrF1BvvNjHG9VXH7smcJH77DVmrzVZ4V53MGs182XQx4WJs1H/NU3ikUor
fLDh74ZekZzVxZRryVHl0JJr+TULIeVUtZDssDer0IC2X8n3yYAcudVdl9pgOxhe
k0xVFSmf6Y5bEHcrYqhD2Bq1HPUxDB3WJlHCqL6JtvrSF1+dTppbMua+wcTy3jne
E2hzctv/1AIF0LjRmjpdzn0dZCJtBf1w1ynHpPOMIKwnaBzyd/qaN4TC7Ol3Ni8b
26p+2ePOVtoXBD7jYlH3/Tnn0NbFVvq9pCGlMBfyaFVenXgJQBDeUrff3mu7p6Ma
4AylSf9OgaDT0pw8I2U4H/Qud/Ou7/PP4tDdmo1HPiJ64hVthEwxiLGp9LU5Hefc
pIiiAWZbr2vjZqGabEDlAIgJNN/dMS5nZx9bIqqocTfkoPQSWNT67E9oUNnGHzNV
BwL+il1ptbOU53FBGx+3Fq8cdwQfF1KuZoBhrbO3C6PahBV4eBsyABi5LIsnGtnL
FDNFRuXLEpKv+yR8FS/SJpsftGwb+yGQ2vHWhF/Rn9y/shqMkKYwDu/WEOg5zDW1
hyNVrry8p1b6sexYbH10I4BKb4QkeDx/DJ9JRULtjIHdigXgPiwW/6BKzlELJa/G
Q0uFdlzfxv0ieJ2ZcWjuFRenPK4+FVLPTnfO48NWfyLVvj/hDXUgMT3aujsXexem
aEYuHqTTxsD5K1PuK/QKGMiUEE+sr/P/GHeE83bveQu4z5VByZtN37CAJQByENmt
0kQDEtOa/KP9ASeXgXJjZS8HRD2RA9/30yVECIUgkPiYaDazvR9/Xklz/MyNhFYq
F1mqq+7xYm+vB8Z+L+w0X63fLMtyUSy3rUxrWCmBn9I=
`protect END_PROTECTED
