`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3yGiaV3F4KKg3aIVTgki8mzmae/VCn8jop/vlWLb8HZxfAR9KzgoQqclpTYS6Idf
OUGi8hFDCMEq/39KZXIWGgS6Au3KgNOJe+SYzu2syMay4Zj4wbxWgPlz4ZH3iI2E
SRF8IIVGrL3ur7ZelPWpSw8GqZc9bg8dZAY5HqhbDmo85zfImvaxZfWiXbtius+h
k4k/8Xib8sRKZ0qOmDNSqM4uOL0el81G4t7YuLqfhBrgnV5DsLev7phfRtISUjsn
MELYH2leTwCWMIOCCdcqU8BZxgjWO20hqILI/uaLZZk8p9l8HvOtCIkGIm+8RqBx
9SB10Ark36Lqs0AojeL+ltH7+RlQRgVKULqUMHnv0k/CoK5p4nQ8azIBxaHtVI0E
R+pWTcbiOVdJ9zDd//qhq2JvLj9tEbyezwExRJgBdqUKk0DauwnytmKo2ryPught
N7G7lqJDxmVWi7GeZ0K4VVmsqMqZm/W+oq/yt0AN7l1K3NwaEihEGOI7p/SoRfpv
6CZKtl6tRr1I1JoqeejQBmrqqb63T/brLFXoKyZ+GUUxqvxft1J2DzxpIfXvx6ko
HokuqDWHtfmf+rX1BCpCNBlIMYFZm0I3x24EqxToKxOrwFDy7Au6T7YIdfdY1zzV
4cJAy31RWvp0oadMtXpBC93QR48YwK3miEa5+bS9rtcZS0Omn6F8ZGk5DDbWZ/kM
z5KWUaTlbrPHwPleKiio7ASCtvOtL7gF2zIj44JzcS1elY5kmwh/daCypgIr//Jl
BKiazLbsrJ6PpRPjBfSPfsPHaxsmgCoxpKtGrED9Bt47VXqSPZfH4/1rCwKGvCDw
fVXo6vBQLP2SkjlgxzZ0Jn7fsZ430/YDoFMOILI4qOlIJnkHUNQMWgSizmofZTyQ
G8fp6DmAR/jnODC1NuSHVSocP+Eh4htwAqL8Auxiui+QU6Tkil/JyMMp7u5bzSYK
mvU/RfVWjdVQI64aSqjv/xXu3kansrYzUTJFUngGYBjsPBLlVNtOimDf9U7sxZFR
731ALCWhEOhqSnEE1cNN7pYP3HfWDWWU/zY1yoK0aonK9vzNnHqwsPmTjjMezbAT
AjKmvbihTzF8qaj1o6L6PDvB2bpzXRrGWSRijBynLsFjrEWYwyYoaO7lydXsZq9z
objI7J8rpudtgVVMnCIktPHZwn1zWclFWSdM8XCy3porpNOwTvZCuBsPW6w89SOT
r8QKu67BI0om33ln9hObJBeA/wUNkv/J1Km/lv2b/s+hM1jBPuLMmyJuS3r4DqTi
7C237OnaQyZwdCuyzfOQJK966RX9ujOBB620I4MDY/1raEAanfBukf5Ab+T4736V
ICLrWjMbPXcuc4qD9BaohGNGp41Fkg1umdWkaOhv6LQoPkDVXnR6FmzzBfjzIfL6
13iP8McKfI+sbLt9K0ljOWm6q08Xglx+H8oyTWyInpq21MRUHuxnZg56Lu2EttDT
hej7/vYe7U/J0rDIdlrVnNMQ2Wm+6GXnWo+qi+Z7AfHu1KVrI9LbKL3O2syQ1gaH
JL/uhhQ9sCjbVy/jlit8uhRM1X3Q0aHKCW7j7PCwkvWXYzMejhaqDVLI6zrvnrKD
9R8gJEzhm/Ef6Wpo16pjg74RVHyxGXMVshXKlX3xYcudkLuAjYf9IU+sNv/IxLBP
FTVeide5A1xCXjHpWkOpeY0nkrVfrFbRZYD7e71hxpM=
`protect END_PROTECTED
