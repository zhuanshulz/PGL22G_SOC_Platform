`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4jenoMBOFkzQGDJP/rDRr/xHpaQn48WpnGHzXjR+KPGRcrZEq2s7h+Mvhw6nH+VX
phK7q+xOBpsqHCiw6xLl6moPxkgMOHKNo98EfhC6l5Yz0U/wWgBY6OJwVpEC6Yrj
JoSxyrhgLTjxfGrAu0VTRThnALQnFgW1eaVm9fTx+4TGGg7VxYpXaTGUiekSIwXZ
QwJLaLzb3uYd76vedaLFMjIOtm07t/z893GPNf38wDLP4PVh+hzN8Y9pCsPUUBg9
2UvQGchEH5ZIFpM9TQdP1WcZHMfYsgpaAG+IlbJsvx8mCu5l9tael7NaGTViQmv+
R36iW+FqiKTYm1+G4MOHh9pqJ381NqLZHWqBl/By9NsPC5kElRC26f40OB7I1yzT
s5yrrfavgl4Ba+ti3kHPggGxq05J11AJ4CBvToQ91sKOH3M8uJLN6ggWtRIrD9vq
84js2ETvRku6emOCmaBH8e5YV/mTXL/M9GzmMgatBmuiDt/5Mo1+P9ENm6Y2ayff
Ed9XZtk+71FWmTRt2teH2ie2yBAgm0lFJVctpXXWf8GsDUUyZ1lTkf8mnRHKs7bD
J/4HCJALw5a+l4uEr9cuYcuRIj5vuecUZVQfFt1puUpXOf+ATsxp5nFBSGIr9kNW
Szyh5vL+F1f+3gWMxaLowfaTk1Nh+kiTLmZZubwkhi2DAqwj3CmKqXo+S+LFAfU2
bD1pZFxhVORrbiwRUpZ31PJSe/koFa7WwQFWNhulavl7FW5djAMQX7QSdHtC0aSn
VX1miPGEBVfAkty1ST6Dt5O58vs5TqZd7vFHrV+B3xMwGXv8/D1IftLsCatcs+Zg
`protect END_PROTECTED
