`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IB0YlDiv5xjFeiup+G7LPYe4g3av7R0+//8ECqtG625YfIW/eaGkdjwGyIzZeZYC
u+HZ2DZiDmABZggkNGsQwDOOdBRlFFyKbfZDm55N6Xpp16/3hzHgEarnMxmLfhZA
hQ4VXhmE9lIkUZjjyIZiGe0Apc3Be4+cg8XsEjViRqtibO8BVA0oAdheGFeAT572
0SVlzzwy6EyZn1aOZKJ/eF+B/CPP72YyCyHMEe/rKpjA4ERzzjGPsOTHAUZDm8Wq
doNU4j2OTbcILmL0jVk1KsZBge9LPYsgbYBSH3tKa0Lb7s8L+qGXKbS+gkWOWHGT
a4JqNdzaISWMNJ7kDcNKm2T2WzXSPEHuS+4gWEUO3wx1SxY/xS9Q3ABOVmljdfEB
m7VJ1m8th5siMKMkzymJekD3OpnLOoiAqL2J/T4LUCN0pXJ2P7Prvq+fUCTC0e+K
uAHZqgoiae+jMrke0bAzNBKUPxUPJaITm6dV1FNNcygOXPtMCYJyY/YrJx0s2cyW
Dp9KAdL12Vrx4DKxDOYdcgbG3kDCbaH9jJFw+SR2xP7TZs2ACTM4ZviZQ6waPMBs
DLlB1s6wT/Qhnw3rRhCRsQ==
`protect END_PROTECTED
