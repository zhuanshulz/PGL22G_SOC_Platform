`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8yky8UxbHillrLc0Y3BOgWZK7zyJm5RJpeU5tizdNUAjhJ4tJ6/OKnsULp846Sg5
kg2Q6JdMjVBxcuFdaWKe0cgXSRNKP3z1Ruv8C8h/f4udTJNBxatoNFdS8PUBADaE
OU+frx+b8D3zZ8+xl1eyx7U24Z0AF/EbH83ND8NFesc2/hYmzgJ1EW3NLsK5InON
MFSNthvYslbjfcBlHKoD7he/AkVyA2qoc4snB5yTef8nYl1wq6sbQqpDVCs2zqcS
BIXalL1Tx+1JzZXuCHCfx1Fj8Bnum9i5TyeBf7nkWY6lyLan7ZAePSB9qA7vH8sV
wbgvftqxVfd7x0RshFtk+VBNq+0M5J04gkXdwEMk6zVuxfhB2AmDFIg+3q9sAd+e
cuOMy56pL6+mpERxmpzzsRgtwdOLk4crqCUBnTJto03bHZD0Vuh3sGpPAJKJ/FPq
NpZi87FruzmUd6+DadL8T8/E+lSzohLn04fgzf+38EdwkCPkxaf+PuIPZlkTvVaM
3HOe5pBPtPluD9Z9mgPHmk6SOakY0lmKjxYT1dTb1hbrsugI0/ZBFon+MB/6/+RJ
qy/ak0ouDW8ShsRUNS97ch2/1/8fyP8Fzvp0z274yRYM/zJAkq2x4vru++KHgjjP
bCyZOT00HNeQfGIPEfKxmzuRQhtGP0ioy+wiJ+rE7ZHdlU7pPYyET3ITIZEtep6C
f/RSipRrILrrS1an2vTqo3q56dejwD68Ht8u0qsoOVOWNMxWDujRwmE8VIVXw6XC
CULO2y7pgJ6ctx4+tXmNAz4yADobxb3IkvTgQ0w2+qynfiwOiPzEeN5TcIEh00lR
fK613suf4mnCHtvJCmCi6QibrSm/1hmhEJvaTvKNZZcAZcVBsN2J2KFeszSNYs6e
3vW/qw0b7XVlzjm2uHTQklnVsK1i3ip5RlPcYRwRF88Y1dryqiZPUTga/oqE7oQ2
Fs0LNZ7WdJcThsX1dTNqDVTMK+at+V6HnYdEXRIP/ORyfRmdTDz7uvqpuEjlYuG8
bGAmvYNxagJo8s1HcTKXWhrav6U6/t6V84SBLMPsh8bfsQ1KFE+zutICubgeSWZc
a76XC/OvcGTJvDNZIgYj7AJMz3qpiFa/xAVbrE1rwWconqcyUCdsNfHyeoC9q8Gq
6d7WchD2foPsgNL09e6BxGJx4xDQlmMG/qcgX/FPawu65qmxc8I0wEHrj4PWpC7Z
M1mc8AaalBXzb2lB72UpMa8OlV1hWG95Z40ObPA0ntdjVSC1IavX8HFAFe63oCw4
CYlWeiQuV5wUGPuh6Rb1tNB9mgK3sODz/yVNbxc7SYIJN0Ietq2d082m1j2/Isuj
g1F2yXin7bBMZa9PltlBk1p16Sg35WIq6Wj6D9VeO6wGQAjSpBan10kJSW7WEvvs
EZr5Ej0UeRF/OpuslS4zbN97dyLfKEW7IosYUay5bSJb/l0M/npCyaFy0uV/eu8I
IW4tR2TlcBzGQacuYJLRepfIiipIf1UQ/lTM+D1GH3nP0G/9SdXwjmpGyuILn3vA
1v0QRGfBR68Q/TmmkPC4nC54o0UUeBX5UCQJEMzktUB2WWZ+9fHTnqK27pvhMt7B
3sYBfoiF13MvN7fgrcqH3f6vzvok4O6MKGolFeWeImDcTTDV2KGCGqxIVrA9Nw/6
11QRAr2upIj8/vwYBTf/fn1lfHXCtxbRR2lCRZDOGJ+YveBAnC2P8I+ANLZoD5bA
Ny90J1ht5su9b6MucqxJzv9WNE9oKz07mRZRmWmFqPlOZfDuHyINXZlnSMn4/8oi
NFmY7Nt2GRO1MdBlXSutSxuWPtjA/aKUMqLTSZRvMb6c0EBLjUCgrMXYz3d/7Hl4
3xTTBs8v03ixks6ot45XUXfHwAVS/QVReV8uFRhrU06nebxp/XD0u4bEjm77lukP
nDQjKVXOMnOtFtM8sUsvKftT7lhgD+8wQQm92gRp4uTJVQnzpWAS8rhDdXB4wcw5
YDjqr8ziakiGMN/mIo2QvlRE/gY5TREuonlJjHeMxIs5LUdI05VeZ9Uu19Yw7/s1
6hfPKOKJq1khYuc+pXvyM2giHRgjxYl25dX9XlI8SAQTQzquh3cibWyVh3lqW3YD
zzmftvXtIJ1HLp05WINW19rBkUUp+8YOzvsXZ3njQ2HmJTCMQ+H8X7miF5WAZBfU
RPBuGdqnCF1jWl79c13BMYwG5PNiBabkd1XydsiztYKYOMEsETGLFlhQbHpVPN/r
1NQzzVM4JEn41aKXVdfs3QeG+0B/40fq4kjfAZ0Y9v//uBgXQu8F2DUC+kIsMzH6
+xfWRNBeSxNZgekOhOT2gysTztCZuFtaNQRKmv8BwYsBtFBdLOzjMe0TglGZQyqm
HpTZ+z/SIsw1p8tm7zhKOd/VpzQJbTJxr9nNTjSI2CJh/x4kiqc6LwrNIbl3NCrM
cocSdoqerVxjuftlWeXyb03hI38VNK7BOCdSBZ5iv3JredOLHmfR4Lu5afH7uyZO
9hkrwqF9Rt6TNXekZjvVofvmMt9zqjVGlxqwel0puwa2PCse61J3TQ786WUmc7Iz
YERcGKgaeOzA/6kRKze0wvifij+Dffum0tPnRvQS6snVInwK/rLSdrqmlLHeEZH8
Y6ycgCG/fvf19pJ/l08Z7g9HSb/ZVWj9n9/luiT/uIHZQTfrJcEmqny2pscqcvnu
HTA9DrSJnMxlQKgGgfJjVKYPV15itnTiblkRmvR+VWCFpnrnSkh4SrmmZBD2tq0M
ozUcJbJyWoIIs06OfMSl91Ivw75+q3glDZAn1F3NBu3AqKeWrsw+bn3sUUz98bA+
jnpAdA8D1sZXEqMjrAdqM4SKkTJ4eOrb9S5invEjIf5CElGdlAtMYvkNUFv54fne
LgmkiYfEJeEPS43XFylh00lIV2/dia9kJnAiv4gx06Vq/pwF7DNew4kW2Z3pSulF
BwkDpvT5Cnm0+BDqwaeePn0i2jcr41t4CdK2TUyleoRxQkvIz25vwNCiYYxXuWB1
rTzlIabkUU0/4HgcGznl3Rr1eW2++JyVhzq1jU3z8gH170G935UpQzVkVs/v9LVt
0lMAiQ1U5BC0uoajGAwi9sKqXHrnwhwMAwaiIRxeB/nyLGr0NJzXDX4l17dNm9zz
Eo3Vc7NhaMJPT8yDo1BHalPN9+/Qe3rQwqu8455wwJPnFFZtcJrXGcwjuAPQuJkv
tW0Royo3BM4rKTzzWBcqNVtweUnE3ndyZectOfq2s49liyPhi3aK7kYNQIBwhxFu
4mvqz1biLgaiMIcBBy872ZwjbZ/OEE0FFCtV12uRpItj4bJCqlxjpab8A//txIO3
9on2MHgrKNQxnPMcMrSmt0k/ilG+xUHfaBrRrIUwY15WrdzgjEEjjow8XHe3YaNw
5eRHayo9OL4GC41sIM8eTMPZ7djc96VBlui9mP0PG+ryVlkGn39UhJRZ0h1laLz4
ZUj93WRhwYwFSZebqUfuSaJ8HldKkXaJPyPm1T77eJJ/AdrtTwe3cF3IW7XqGDk2
05pZTaGhFc3+3iCFSt3Y0sTuPYD3OaVzl4IygHOEhPZxYum/4CvpQPjnI8Ve7VGE
SP2mrEMBFoQRkSo9sSTmkR3AU3xFmIm9BZ0G/I9+A7+C/nDwD+qnZ7e14yw+bY/T
BjDn9ITOrBX10M36ul7u7WEne/Iyxu7hxRa8/fmWNWur+5Ld+1fLYP558DKsHfi9
XjMSN7uEK+uIpmgU4OJAlCyMMaLtt2V7ldePIhXrQajmG4gYoKS3gSqnVYNxFjkt
zWfrF1czlWJaEPh2wC9Js9UoNyXa6hKGFt+oiz637hHRcw3MzWIpMdtTdIaCcBw1
Pl81WBlyk8U91Nvx+XPVFG18+zaFOBle8tq6svl7sZ1qFy3GdKF11sOES5GQzLJJ
zJnrc7tQ2NSiIysRE67o+2UYtoWDIzfart7hXCJpura0usxwiuNcVFYZiVk4XGm3
CvGYKJmECwrc3NphrxbMXeLVYqJQuCtGDUPLjC6rL01obPxTA3NNCwfwxefmpyUB
tL236nHoKycevh7yiVzWvXJoCvlD2aNabJlSbxTWHeVk3giTyDxiILfzpDgtEW/E
q62NCzjTtTGOyVx/+JNEa+mrxvLHCnGu4qN9uhnEA9aLH73BTIfD4ftkEgnipgg7
wlKmVLyi+CseAYZxh2Ig25/I0zUCmwAjjXxjgc66vcgA+qixIadLUAXlAi8BtxnM
v+zmelvoyJpMU3W/x8btdPbsKPnEyNAdRpQOXHpHkvlY6KjC42YA3wEJY3DB2dPH
ZrtLy1ydTp1IOrkxtZRE7zppm3BbF7wpOnPZWLT0AtgBLxeOYrurfunEWYED0Yid
MnrO56hbh8wFBe5q5qID86xwwD3PWU+6MN7WzbczT44UOVs/Iq5/D7lU4BKFyxiI
VsXK2vXWshVy8Zn92mbcwkmzHN7JBOY1MRb6/xpSQZPlYg9VmRQaRbxOIXJxWbxz
KFk0uAMZ16c9/w/nunKK4TskzI1bpcnFUOtM9fiZGYXKa/6xLyfXjr4ld/E19lGB
R1IKXTZ9/E2jlUDvSHU8v03LmR4gQwDyczO+ln49WuveWIK/0zpgWkiuASfT/y0B
sJkUCKfKjtNlImh+1S2uVreadnuejWIU9ulGeMvSNc4MiDIe27ceUqj7yqLzacVL
xJOjXQHP5mFL+BbkA0iOpS9t0bJ+vLNXjqH1v8o5RpLNyWi5vHvqIh54hX/jrn42
HMyfQ7lSULkvklaCi5TbiKzF3vpfxKCTuKz+ZSA6SeUbyAOnAq4Tcql9sqVe/T16
a+jIKXe5XuWtEwmmGPJmepqIqXwVLPzCjif/wsalqwsR3XdeGQJzXqKUgorhHZyl
als9aryEsXv3U7KhfqfRTaAevvLiSH+tmjO430nGiGLMEJ/apV80d5IC2KtLvo8d
`protect END_PROTECTED
