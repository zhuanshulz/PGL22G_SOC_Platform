`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GjlIt2WjyXr+ox8mOeJGr34w7YI//CsdQ1SotPdtUFn/owS6E1PJXLYR9zJkj/ml
YHbz9zLFEoJqa0e5aXstKX6LLU9Q31XM4bId/1M+iV5XePR+Gi/OQMPdKYcECvPS
MmjNyqKaNZC6MLacPQyGutT/C7UlnbssR7BW6bsDLQTHggKiHcSU2S8m2TZroV0+
LCapNE9I/YEe1Tec51UaCyvTZtKPLzk6uGCocHLmBeirnUGcNUXIVqSVeYRcYQ6u
YAd+YoEC0o2EMuZwK8mvqkNrbWNxU70PuojxU2g2MxlmaH8Wi3goRs1XIXOMG1+u
cnhIYOj62JWPxs7wLGnEdbXSPkD/KMy+3PSw5iq8yDi1LbFri3QaoqUmcLcSj9Ft
rKMQXl584aqhBr4vA3mSxRl24vKJJHcD4/+r8n/ijKDXCFzunZg30qorM/nskBoa
hJ0yHGkSWE3n+yhLFfaWwbO39rZp7120EvuZyYUWbneLaGygLRb65bm73iuEAKk8
KbwTM4DaJ62CM1pm5/a4j87eOq6nwYhfa2Vw2qiX8S0nFeAsCKoEX5zkGJ74wwUG
XQnU+qedqzelrwA5ueZeyoKNz4WNkWHlUg6obBBqBbXvP9F/YPCWeduXt2kwUT1t
`protect END_PROTECTED
