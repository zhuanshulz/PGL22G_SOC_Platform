`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H8NvDUaWZg0TRXY3tNygP6ZIdD3svPy+VtDfiwdQ9zKm7OUedDPfn8qW+sTiPgoq
Iz0AHd3JlqVrlZA+XbXWUyoqXWnqPFJWLt07+A9l6T/bE+18pZ595Gma4vQYeIzs
hpDe1OaA/n3zZGF+h51Vwp6g15IxgBcbuINJ9bEDYs5kkqMElgCdnaov3EE2/nEE
d2VGRpfuKS1fK3E2CidMkd6UlzvItKFtQeysUfGeyosmNC93dSvPN2/diGzm3nuj
5MhB1rwWvsBe5fJH4rBMJvZbMkf7QigkhGcMHtMQst/+TwCt+u1j3nBWUriETde6
9BFkqA5os+w+CviUrzR1ExIYCUsk0FIN/gE8hOOuMrdim5teOr+seLNz5/nDEnYe
eqD799xTKV8wiUQWbxMEXy5BZtZl+unebCrPGB4BDXTy26/4DCJTLmOd8AoYWKYF
Nfhqsj8zxw7y92Rs59oBNe91HD+xTup48GHyH0daqtjatJKVnRAtihDfiPbnhZyd
N7Vb9s4fRgAaCUey+SS3A2x4tONAGvZqlNC7T6o0bSY6uXZp/NPeIpEEVF3pyt9C
MGj/5AGVLykrMDhTebOXVWIvr+86zILc94BCG8IgKlwR0ohSldI8NStsDPQKRRsx
ohwqBNNYzCaHvKNkFdIxXm9lQ6GsAyOrv/kOUgjADBMx6Q9DBv7pSMwjKlwX8r+Q
htmgO0cvYPA2NupX3V3cqZgavLdPavtqCzPnoO1bI2/8RvNjg7TIi78yH0EhOgM2
yse/TP/fzn7SG0TVWtVMHp+e8M+MRbTITV+/nrVyuENJ9TPfaH+awzldRHm3C3Iu
5BZE853P6EIz7GgZl+z9AwfyZMhLK3ap/+qH4HRQS92VCEtgEj1D59Qu8sc7wRsb
CI4xlJHPEXtEZFZj5YWV0P+WFuMviFqac/ePYNolcypnNZF/A4dHFYqpP4ECQ+9T
zMgWwagg4cTNx4CcRXyQyNRU9Xi0bFZ06Kel3T6PshUrdGdXiDNjdtdTbnLEoMVS
hxHLFJq0fr77pKJ0kI1/HV/zUIi6/+L1ifyLYsGuUIMTnKxS/DArKVQa7F8GxpNW
jYrSobrP5Z8uIXjuyrZeIsJ0LcS+hLD/j6lng55bTGcZD3oXWoMYfWo4+SnFJZ2J
jd6bdAQrXWKJYbEI4UDoVcWnZFQyataZhy8b37SovOkCtoq+24fyH3QtQJQqWP2/
pRrrrrZMBbntOaQAqcl2VGZ0+ZxGMz2BGuCBVEJ3pNJ23eWzRUPoHBv5Y2k3gB36
O2+53vn3bXGY4ypUW+QzNKjOqvEJUIR6Xw49GB41FprWi0x0LegeVttb/ZnT+xQB
3HWLC/MRXEJYrSFbfLfJh2+qdkRE79d/9qmlWDKGrN9vmnpfuJXdYsVpxXxjQfih
ARiSV4NqTAIM1Vu7KqRJhIB0nhth3sqUVVhuqvpKs1Gk8ZdAOGS1oSSsmJ/dRlAz
SjDRm+TQKYrMBgOb0R8b7dPZdGZX2o5nlP0c8zrb9jt+oeT+3JyE/nUGgEMM8Kp6
1yPz7mHXos1oQ6mGr5GoeubF/yJbX+qgliLq89OwqZhv/7h+rG1TOfKEIeItpHzf
IQQlDFMnATx9LtYbjNgchl68tYpR2cq+KWdOpCPN79P4BzDZtnoggc8AWzTwFZsf
LNWLA5kYoZBzyXOOyTD7ohKmYfS+vCh8oL8wW+N+/cGmTxD5KAZGUHPr5BCSHB5P
XzxEs1Y8zLv5CDGRRetN7tIoMKJh1BgFV/+yPTNHkNPVU8vuKIybYu9qTuZqXMs7
/CPFqaqkrxu49R3R9Dc5QU6WpCVz6UHEm+3JLbyPpHwHDFitDHv+59+5cHGgslDk
TmsqVFBID356wi66jbtOUHJLZOI5iwz26voEQ63L7UvqMsshSQJke0CgvbD0AaDY
uDq+WZSJOgLvpIJ08kAHXFQYJo2/9+1Xe0hsOcbIaxdKvNPtKD+1qbOc/zNT2g7W
UXN2iKTeK8XDMSuj6bMII2YttB8Ngb91eu5B1yWpNlCky1TzzSZbToPIQy5fP7vs
nUwJRsrDWI457oMvvbzJYFPFvuuU1GYz3WhDtKNznippAJSvxiUBy8jsh7KIl/vC
/+kSk275D6g3bcrX2VDkgSL83pZA8Idml6ZTqIkcWqvsF/dWOrd+sHJpTlyIRnGc
Z69ao50cO7s5nrDiEhNmJh9Gl/oN5v9Oe55PrhZ4YjF3FB//jr36KXlnqvp7Fsls
eepQ+L+PXZrUJjYHbLn5Q97wCAM1+BveqyxHVI0m4mIOcOA31X4zSL+Ps4Txxssb
PnGJvm+6kIyjwmrKjd8zE+8qbcniJL2h4iJ+yq1BAFEDJAwksyVnFvA6ko/Trs+X
VQee8ycp0pCF0MkwZ7G2HU5Heiaieh/wj4t7qMpeLJYF4fsHz+ym5h3FL+De8hnA
Zpf2qoJ+MAX6lE9hBr04Z4WlC7byjUJ85hZGurYA1R8fBhAWG2pViww1ZFHcdmyf
4DY+T0MENwIXjqmsItXh4d+if38YJ20bGz4WeUKFp/PaeHEeeDhKGrKZftutFrfe
Hfs7NTdlspIvAFNUJpX3lxW+2Pl0wY+Gdq+/Efz7Gyp78iGl/l2lq2/nKy0Ix+Tb
2gLuw/0O8xKMkWBHAMLuDZ2kRjNRq0asLJqdf488kg80CiWg/AvC0SutSwPiVXol
KNHbwJNZG75jR6DDmttQV6AlN1cW0S5docPWeUQLUr3oCGlrckRUUJMRoWm7mm6A
fSKNENWB+vqQA16NQvOyTJDaP5a0Oa1EDGVMWv8E5NJjR4S7pY3tzlAVix7VWTL0
KYadaiZRtasb/3PPfb6DdYcF/1TfSd1wS7AQvqtbApIady/ICg7JT7i8Zadbsymx
IiMBLNhCTE/ByeOBrvFNnTPPw+2BNVyudhIfGFFsshesZJJxjPB+dF2ldKqSd2tJ
EnKlGlxsy8Wi2haQB9V4/8t+PeIqsj1BNPtWxVo+G8wx3n/p6AviTXCK/G0qPXTZ
7LNcyQeOS7evEwFai1I0DBUumy7IRQqkBQiHiPpyxSjU018mknTZ0uvi2EhQDVAA
Kj6WgulTUpbuOo/vI5cOHis81VmiwBAwawX5LFh02hvlIoRnRBWmEy9ZH1fmkoj1
t2s9EYP0rcs8Cu9xLaFKaX+ImNR2c2c0cb5rJOygsFk5qgo/bcL7eCYcHgPwA1En
NRDmxHhnuCRp9cdfxE2TyyF9Oc8m8pgBqNx/SrEypd3yUj3+4NzMP2gey7u5gXEQ
G3LZDCBI69SJp6JOGCd67cI7NZl0jlBcNFey1WNj5SrWXAMuYrKOhoA1pG8ldVVk
14vo6KAj/U1o+9HmBW3g31gskmH/R5XjnJ2znmbpWVYJvRMkjE3fPZ0u+6yR3ITK
OxOm/8sVUnCnnykeu6LHZbeQVqGRMn+dp5u02bYT9JUcW3ZzD8sQPX4ysLtj6t8b
jVkc4mjcrGIumhyAyjA0fkvWZxME2PO1PChaJYnQdiqBqmq8cB39uBLu+3fOUR10
oFZ9xxMxpQFZVujWdgIOErh8wemh6Wb1t+4hpuGNkP/jXllOmCRsxLygGB1pnhnD
ivF4A0gmN7IGMiPe1/8HQMtE6POcVxC1bTBzPhKR9kfkjHrQuKEM4/TFbkXNI/UB
5nulDNeujCsxJCwXTEPcMmxvpdebT4F82f4EVJAKseou1hPYp2qYdneo3hXGW030
CItsph+g5Qwb36qqGA/lPOiKHTajyKD6eCYZ8xfjtWboOCXF+VX8B8JhyWF54da/
oedCMoWbsPiA+/LeFkNiDbaKoojqAqqF4Iz1idiId9vILuB747+t9dAzJWiUfSFK
zVjAC+tAIb7d1WYHua80z3Qtm0upfxdZSDopOFs2l3LFJU1y/nUHg9keJCj5XoGZ
8c1vXxid+YsVGqXYkL+hUDx6ju/7bnfBzm17LdTbxHFM2e4/jE9GCA0UKxWn2QgV
7eHG5susTejIJ1RTV9Z1+dw/vhp8w+N4xuNcP5b7pDQBqpNw7TM3PMlWg933zmlU
2qUwrtACPKDPIcJGAbg+F32khPkKREnhcZrnKdNZoiYxJBf6Q1JrjtiTP8IWNuca
UlbjLctexd2b1i6Pv8wrF3yb6MzjbBoKMKM+rk7byE0Ga8NWHpzZTKKQ0LzbE9Lu
24lOQv4vXhVFSSAgFMmInQGH+i54E6miSWLkhnfL5SUxvOR+0jkvBL+/Ktz/Vt/q
5w9RqrdR7+hNledYDSZ/Q4O9RSa6s97o2e2X4krj8FRLr5KbUgAlecUvbdeqJ06/
UfIclyABNiuPtwWHJLjIWZpboHpTVasXearnna1lgSNNceyzNCi77ynJnQH9Zyhl
pMExzDRA8kvV/On0VJ48nhXs9fwmul9qCZndXtgFhq4ytTEntEKeTT9bueGJkMrz
ECoBeQPyg19+QGKciffmnknKBeKsWGihWcdzRfZLGbKeUh9+YqWz+EMqd3PtO2qR
95+LQ1i3ih5mPQDOIx+J2fpRJ627wDkc72He6MeecN79JCU+Fd09MGk1MVCJrSRr
NfWEz5Oi0+gDDTkw/3ktYNH46hAcD1fy20jkhjHMhHvFf/vEgMmKNUryOXBanJ4Z
J+WIAXZ04rsgO2jBln2do02sPvLpkYO3IIWRJQqkVnMdESv4jBDIKQcUZYiEzOqV
G3xoLFzSlWJ+2fYR/m7KPZoW1vuzHv/DkPLFzTqvdixROxh6FtbaPnVu0T5OzSTV
DKOFgSF8LvNlLDEkZeg202v72HDtzdUgK5pLjRSBwL+tVPnaFcpvqgRcN0X2u7LQ
Py72OJhl3Jo9fszfVMylOjiNj9SIFBnKQa5e78kZVTXrj1n0JFTueyMZToyI9tv+
SQxmUINatUPo6oiwfTtNbTwdbp1ieYh/Tw/zA3XTN8Aj5A2ypdGXsrFMjpYQ0HKJ
Re9h4P0IUPF5F24WfhZUyX2mMycQ0rZx9QtR7tbZeP2laqwcw4w+cQqzyPUwL4x3
+wvw+5bZWp+CCTUYVEVwXiGvV3Nh5MBDadmLg9S0QB8HvjbpoibcMQRH7d4xx96j
NyDW12T9IC806sU83qaPdVKFTPZwKvQlq8E5P/xTyEKdHjluNQI1nEhthaJyxZPX
MGVo9DNYgJlPYf63mnxik/iuIIckJ9TJu1sxAvER+Fjc8oUDPt5+/crLsfTutseK
YT7vYSdbEv6JUchmewIN5deimFld/TxOGuE+dNUwCBlxHW7U1MNcsM0A/bO1vDn2
Y0Wyffjz9KvXqeTKP4jDkw5unsqyhgtbAsSnThMrPkhBZTUaySjw5E91Q5gX1ROP
Zktgv6aHTdYhtwLMqkQNZ6MQHTisBC7hyQxiy+jucwdiNs+VHxpEcgmL7g9f68ww
daUjMMevsTxM98isTSfJsG3oiYj+m0lNgql72J8YI4RyjiDMqd5g2axhUOXCoyVv
UldIwyTnYf+WNBo+TA2m7eATjkFgW70Hc/5+Gtpceqs=
`protect END_PROTECTED
