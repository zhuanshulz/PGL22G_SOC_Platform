`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vLg9R+x6ydPrG2kg3aYTS9roslldtHv9SwFbsLg0eVbRnjM1W+uaeQC+9wq83VbZ
FDNamXeY4w/r5npvN9WgYcQj8kDS8eQJVjpf8r2t5PDho6ciJ96V4DEgObmQcV9b
izxtuzusInqk/CM6KvQf5R6BL+EeDRZudv5oFk04h+8Pm76DcRDpK47TATwV4Z5Z
Jw7dXZSSprvHNqKNkaV/aTNQKHdBOPvRoUtpLqfqpLNZnyU++KAEr6Yg7YJm5NNH
WsXkUH73CZwtYEACl8xvc9zpQIqvUipEWMTrlcW5Z0V5Enl1Qr1F5pomITo23jde
qXks/gC9JdTT9T0yG3QnOjbPfcSdDCPGk3ZRnDV0iX5nXY05X7W2G+rAmwy/cxmE
`protect END_PROTECTED
