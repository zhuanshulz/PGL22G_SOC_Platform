`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SVsxo8PRxZC0gRGqGYYoA7dKq2HqEZ/jOVU1vF9ANu9gVlX1+09x0hhVk0KPLOir
fwi/fp/pnlmxHZK2QIHkeCoh0DyRbCtLp+cy4hxqwn8zHARj3WaD9R5NbU+mQ2wH
eqqtNDy7AwQft37Lak7kM0Ar2Cdqiw7RAL1cJ2GR8CdWI7rhFuNiQOJN7TYNKCwp
pkjLnMOtIRU6fBMu48IsVYdlrZUwg10003CvTL3gQJqgFP6KDH/YaFsQ/MF00wX7
Pliq7SAWZNK2ismkt4tXEIh0ulbeoxWNOKGafoEkrjbjq4kpOzeiQtzSGt+vlSlc
Hq/ufWMoCY+IhzNUsyNLAMebUMIHsRV2OaSlEi+bGKPzr1zkdtHtWWgLvnCIANcn
wMCsvWsQC/z+nf3JJZ4mue+x9VP+rWLmYlRil1EpbaJfsaHKRV4Zqty+lLgxezpi
eKSBZQ19rZTZH/cJF/23OvMrjwne5WJV7OosC/1lX6RDXyLZtMS4uap37X5bv+kl
56Kj32DlRxe8D/aN9NjbljmcbC3DkCHLSo9KkbqcFyfAnBPSZeICTFdIMa0W/l+0
o7f5Q7v92MwXkk+dmDXbsYiFdNbvwjeCpH/sFoKQaQrrC3avDsEF1guxo41IvLbw
kgDiHzN6QswYWmbBTpj6qrG1cLWG3U6kQFddJmOszMqWNozE6HfMY05UUIzxC2UR
rwbAxNzSa2slIOCDpVwbi0IC8+o5pJFV/qLjOzDjQZtzLohKeCADzMWofLxpIZwy
ur/kJj9dS0VvrjBSa0RSrOaTxtdvc3DgvVFicmf63+WdkWC74dVTxyt19GPA9IDr
3uz+qYl7xpxkrPiWyukUIpp8z+iBgo7VF8iJBx2rZTPS1suDk9/eQdl3avI3zrr1
dHfj5hYGK03kJJcLk4FL4ZPNRrEXm7Tzx/ghLn5aOjQhxlJV/4ckgSI+cyXkUtzl
6KgI+9az0VWfhKC/eSowGtZLlNaBaTZd+4475DhAvsrjjGlGpycjJEYANvH5JSSn
ToQWSNcU6p9uJwyKC0+WHQ2bKYCI2tqgmJ+l6NMVKRpqYtiLzT3n5kSlne47MODa
enyYZURDYXEHRWBguxQjFfGU3iYDEzrEXsR/4deCl0oGHIw3jgBVKBmN16NJl6pi
aDONmVHfw7CfeQRZ5fcp3cnDE5IjN1ugkVTt2ajibtsZ3xYaf8lPVBdUa17ArQnU
fTini+J5C5um36h0useirAzA7xlnlQs4kQEBEO3N92OnC9uu3ZDbK4PWcHIGhYFM
hGNvSA+EKW2zn1H3E4jD8Yak35VPbBXdXER/Ui2UEsZV8POvGaKls2LdfNeZqVJd
9wL+mcgDMxoQcohKKepfIMZXmCZkncNAoOI/ohW0Ly+tJJAlnnjCHBmRISlLw9Ox
kdXlAjjpyuMGUt99Chze1+guSgm8KHS6zGwi8bVEUEmp6+G/qBJtRsyvQ6VZqM9y
ZWL9pP7gKCbdGuhql8v6wqnIvxDFfLf19q8cpteEprNnJr7uOMbnBJbyG6agbqbF
2NZ1fw4niQbr/zROwH4bY50zYy8Ov4CbWIA07IksLV/SLpjZQC0uZjicDF+JKefq
Ex5hvhRy+0nKxCR3CHcaR4KWxGeZthn0H6HVXD8DeUjdoOCDmbOAbHX4fDaE/s21
1jJF7RT2ow10QxbckQd/cjsfHtqhhbE2SM/I5N+eI4TLF/LOwDs2v+ZUvP8B7nn9
Lw2mKMtNnzrmJg3UN7hmC65uvsDO611Kd0l/uVgATUSXQg5/pV3DQ3lTCeV9K8zw
JA3AAgRBhv5J48FIkU9yt+mvARi/U99oWYbWnmTUaxfbbo1CcZty9VdHGSf6eyQn
1Z9p1zkw5RQ0ZUSPUhEd1jngSb4tqaxM1rTIXqtu3YnV3hYquX86J8K1OtUZbFdj
2W7cgI9KFEUP/gPe5Ix0MCQo0qZmiBgPgZJ6gndtSnSUwxI8QYYDOLMh8x5gQTS1
18mwDghLj25Rffl50LSGNR5dDtuWh8n7h0p7Y6w15+yvVxUSXdMQ0vm+h3nNN8oe
nzBB2qR5OYebcLfKWI3xc04rKO8SA+7XwC7FySzXzyFKBlqwz4IPmC11Rr8+9R80
lspgedlBFmFonJ/EaJNC/6sxN6N5vZu+yZJCHA+lGkFXlWxRAvgrfAs7+Iunoq/O
8qQf755WUKcMk2Hg2ywGZxxg0mOjokKasgYXsc7XXgqKUmuxkb3i6VI92mwHoXBY
QLwvzxJauzY55nIEsxu9YzllVG3R3YYe1yHDHD4qTE8AcmzkgFwlYYyjgbYLBjCs
89XvGv9BbsxwD+4f59EEtwGhs12yBwJaht2sKVbkjDHa1+uBueWIURuYv7VFsaL9
UWnuDAshldaIBCgZgTE24R6y/FedKcfy8aWQfjlXDuiKEEur07kmCYUx08lzfcC9
++orNhlrVy2n2w1KQPFb5sMZOjClt6WWoLk2edxfqQOBWIFCdbldq0jcyj3UXk/w
cHYqd9QlrgeqYvYTfOlnEmGM4y4uCJcVeJjfY81RpcqGlhCr4DZ+BCtlvIRj/6tl
u0EZHBzKj9ZVP/YP5MiHczR+XK/4i7LccTD9eeWWat8533uavhQwac6ihuIHLDH3
vfJAWdpAWPzHIFm8obeDoUPctgEijCtfYlZL+8llhMbAThX3JeLFaxX9b4hFZYxA
smGj2O7NHUnuN6OJsZolV1WEqI5nmUpt8QDE5ktVQ/TtTBc9cBYp33zBzMv+Z3++
mtDJi14UEIsUVCaqd6O4Yh6biJ7qzwv9pzCgGmgcQuKE8mcpY6+nVmoth3g1C2+m
aIZzfE4VP2cHYwbS+4eSg4y4Dh2l6A4WowtyTVAjO+arvsh+D1QqaOanRqgkvwUM
tX+izWeoCuebAHbxEiRIi4un1XmDrJbudChHZDH5LhIznRy5fkgxi0D2CNHlaMpV
5+hVwTVIgYB57lWK9IanMezPSpODU0btS6rVXc74JwEX79bT1v427JwjF5lqMWLE
GzRPTLpmlftsP+qp1NKtI9fkg++2Swptqt5VpVLtr53Pbj0KFklDNNPNcW6yGgMa
Ug+CKD85ClR93nqDQY0QbtXPZJJMOHSz+JNCzmfXsYelewt5dxAzULWC9/rOzk3Z
qZQ2Md+YMm4GOj8+NtduVXzS3/Y5zrH/THDRFys5bAxLoq5Fql5VxG322MXCSHG4
ialQnknR8/7IXcGN9q51fTizWPNGogyjnhK2vsUr3daI7X5NoEYlSEql+cT1Hial
eSADbrVSNJfhdD6c/2bN2Yf8NM7Me4pkmizNNv/nZaUGaeySNLWpuSbZUPy5/Imj
bltHF4F/NAyT13CgIZtDND0J251wLXx9SKxGbLSwtJVembfgWMO9fPpJNyMXRu5N
NGNMkr7ArnyX8GLIykRxVEF9Ftdod82SE4MORoi7IACjcvXKcBsSnLj6JDmzStoe
FbnRFh8S98DU8fK5YkZn32fsUnc0EdgK17PICrZAAxQnvvOqkCpWCR+uTwSS9zzU
Kdl2ElK/DheyCOvhbld1iQ18If16cmN13viZNXjLrLvjPPivyJmms/tONMXmbYwv
T2wFsHr2csxrP3+WSH3kqCGESJTbpjza/zFBM5EdwMAmDAcc1OJ/700aLNHQwpKh
T5RMefB1BhW1WrWquPGPvsT0p6kdAuggmfOmf7Sa7ZCxSiOhWul+P508uifptrHO
fvzpFUVCiULLX8/RgwAlzxbjMVkPsDQLeUwatTYadZjULpIzpaSEbkR/enga14eE
mwf0U25mStWW8e1ilg5nSV/+GO6TntR754JG0ldrQYr2lY+KWSh9c/1IVZqPQZkR
vs2/83BDz6yLrxb5YQGkNjFdEMeycu5AXz4smzSfnn6e7+vCkXie8khVZS0xD0tB
hQ5Acqn3izFsUvpxLEAqx7tyllQ72/9YEkNn5dVPvqyeIXKt51u1iKJiLrCAWbQQ
8hjZJGvuG0BjWbpi5Miyg/4tIECjPc46Z0WFgW60RNYmDeGlVWZ8QAW7FGiJSH6J
1O2D9aTkzvbwh4575PgMNKUXCgNnKbqpbxMS6yitxBRoByD1r/i6joGWI0JCqpf3
mCvKsSsWyHc1qbggVja+dCeVWSBdqsMTlztwr6IvM1b1SLGyTuEFv65yS1QIaF4G
jgN8i4LOKkfE9TlerEnEHKC5eXYHHvgrp/PuPzJMwt0+xx3e5g4z7n6Ij0kzKg8S
mkx4nfwVsNoAoqfThyfZkAtbsLKq8ndm/80R5aYmvGz7w4DR7K0nupwgBuk2OjNI
pLXK1nWpwZSSnmGM6dJRLboBz5eJLCSRe5hP+vKfuZc1gETV0/CtQedeTyStGvv/
sptEKVhA0WdgUd3aQmL+t/mKqeS8Xp45e0dWyobtT4DanYQ7rgrbviGSvqx91fhS
lKZwChPUbwvT9OpDyr8seEa9tP7CaZWWTIJHywuYS2XUatR2KY5Gmpow8lWpL03N
bwhwxxAfzcXSGKeHHOeWbCEBGelNMnNrRha40x+0l8u3jQXpNvvUu/vdgXDupQiQ
pgFfKc4R+isYSZtEiIqjeuzybQddKQnK+4FiCggG1ZRaxyRd74CAwbYzS+e0ZwmN
Lar61uMXo9Dl8W+UGMtNaQ==
`protect END_PROTECTED
