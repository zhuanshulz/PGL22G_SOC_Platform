`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pSLfgPNSm2/zYcof4dePIONh2DAL+L9kBXJOtxW0QuYL/HYeWLJj1PBze/aaVjDZ
QNTIWSoWF3H8PvlGn7yGeE+h+MORBxVCPLIUAcaRy3SF1F13O4Feu4DFjnh5Ol/q
g5izgXKwILLuiIZUD+I/8pfVVFX9Oa7sPnT+kyY9vTESRXv74sY9DkttYrGXdZ+k
QNSjSSQ1P9WYezG/fj7vplknn6TbSgUBFo4ZOqtHrjRNYWSR1YCZre0Es/8/NrTO
B4q1Sqml+Cg/hQriUINn1F5X4l3iqPco1A/4v5YxIPpJetftDIvYh1p0/wUnV+9h
JilkKQbjWQCzruL6KPT1GN4xy2q5CQSxqiQKZ4m8tT2lAVghD1btZWNEdFjgD0O1
i7kn1+N37Nt3+rL5idRmjT2UgWKpvDbM1pjbXtogqDZKpmDG9O2BvQLM1yzMMPpt
8xVv5Py3GF/bqDUTxxY3z9vNvjqoME0dU6bFCusyEzQwxBi8Zcd36kXQxLmFLuJI
idIR11BcB1j0LiByaa2o/T4zYlLo7kaEqYr60zoTuRViZ80GPBYrPLsayvjKAxhB
YI8FYeQ3JWk/Qyr3BQtkU503pOwYztbpf2r5HbfmMJOay33df5M+KVFGjb7BTiR+
+P+/pJYNDVdS7JG19Gfj2nR8ZFJ9m/9+64AwNYVh0ttlVUF8b02fexE5MkOkb6JS
uQUequPPqHKU5eTGt1IHHyXtk4ZvSiR/nHIaQ6Y3bQvk7EUxniRKlF9Jf0HdzXOL
ZSeVLA/kOTXVHv0yugvtfmTUmvGh/tjRubLvBVaC2tJ6ngNUQgYXXNzakwUWAHmb
FniKZIvZ7ffIa/ZQMZm8r1jj1I6aXUE0o/VTEHA9v/DMKtrdqDMRRw4N5Dbb5VVe
ld4YJpKruq7y5gtvm2fP/loTULjZVg5js/lOQSSemw/PNYGW9oLaYZGc0j8cTYXD
tZ0RKafcg5a02cvPUm3Y4aaN0V1xfAFlHUmC1j87cnyK8S2BBP5aSnJuyRUFIlFY
W1VgAPgZVGsHOXlzXtoQjHv0cvCixfXFvLP91+X8r2hIJ1PIWqWywyrIzMbTjJQZ
heV1YxqeNd2Gl88M4Pjlh4AZkxuvuqHNsxlSihHg/ktnjqambI5CLt5gDTgimQEU
a+Uk2n5M0AOEw6gYEqD9MXAuziJNjeOyqqRzhB8D19E8PWNy2FQiana6WUWbfGal
MYNRSjKDApKU5fS9fmCMkYSjJgPWKBI6HQSKpg505uatxh8SxvJ5pUGsLmY986NA
E29SbCjB7qMCmyFIr5C+41Mwfe3y//zAF1fTUndHBA5SfQquHilCv3EQrmpsmM15
yly0jLrbSJrGFt7ZYZ3ziGwEshtejLYFFPCb5O+MAmBtUtQ+gLvqqdofO6N2nY8Z
NE6qZ9bn1cvO515DmToW97M5WmJr39kjHT1RgUmQyAkdBTLlrLbathxUOH2CjDdc
rj+JddbBB42hoKEgJWBIwq26+wMmHQH992ThMVu8WqXYhlx9MUVjZd9GqLhlVmR5
A0ZwpUIQLxVN1TJwtZUFn1zSIcVSgm1tizP1Qxy/zuGz5cp/F8YhnqXRs7RfQ94x
kDi4UYebGiVngDuleYViGOK2px7CawJJ208azncVeojA/gXCaGs3LkIrBcYN7q4k
i80Ew+wJW7usN2tenOXL09GLwF1yng0Bh6omIXuu13I2fsRogaxRS/e0Ib78BQDO
oD37NPvIPzuv/DdwXsNfaC0tWYV/2qdSeRu/xIplAOldb2SZbiILSH37EEmxkho7
vbpH7tKmre/EPvq/b+WEm9typwFOa/PbKz7uiouW9cegkkG7YcrKdQOKG39HqzKr
fhFQG6S3HWR1FqhZdIk3sA==
`protect END_PROTECTED
