`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uTydzn/K26M4vJrZ3I2c+4FDow8Xf7WWVUd7wtCrMh0ZUKp4b/k5fhFVlRgjCkSX
3J/riofiVH1tll6gtrPEkRU9t6qQP574NCSz3XV/pMOFxlhTCDYnlNV2VRtpAAyc
hZjRsbRB3gg0ugjzTfzMi2lFSKNOMHOw7I6677vWfFTAgoe3I631PvX8iesvjWGk
X3/lfSTaYpqqg2nt1hBlkpa7HUwE2pyHohWIni+Tj1ngzBx3Yy7H5DtaKOhkzzkP
rkbXnopfAxHLaVPGLX3k3PvMDlZm9ttq8p8zLIQuXqOQHjsJbg2exXKiN/qHEqeX
BKQfnr6UJhbn5YkytZhF5EZVBiz6qEFroYXxcdzjRx4rY3LbHATgVq9dfjgUDlqE
1iOLAuIxMD5IWY5pUMbkLwvow0vEMmpXmFxRAZcIuxHJWYftyWfVRrpqPv+i+EHC
gXlxu1+hFQuREkdjiQ9jGekWd98JXwBav3gd8ABaQeMYfN6QrwatJbi1javjzzZD
8LElP+A7RxQghtLP41ElFZD91o1Q0NKdUptbALQSNR0Ormv1aaT4ATbfNVIkYZzs
mcR/30aaHSkgxMDTRp+8DK2Lwl5Qdrne0UEvSzNFnfowqgw03gvH6ThESIbOZEmM
ZbeqgeK4jYS++nU3EWXU78CLgc2r0EyvtIH3ns+PI29gf/2hZHro8S5D16o0/r7w
RNvz9CsUkkUe4/emXi+/1pTxyBl3LWHnj5SsvT6l/k1xGieIBmIR3U9HgFl8ObvC
iPUf0S+YxCVqcZhiZJgxUf5kGGznXfRkxUMmuKSuyO392VM1yoRLKM07yMp8liIj
ya7HWgM/Qagn+G3+qRZUmtelIuuiL9qs4un4Dmr2vKCHgPB1z4HopWkUmIQX2rhk
TReqOd1LhAn/rij/jIQf/7jiNJRsbiCBmw1yJ1EhOpiME+OMuAJmpkISJzfA8yFY
4WFt2yPyUu/51gXLZfc2oe8d9lLaY0jsMcd5hWrED5D47mxMG7MFowkK/elOMav7
+luMuOUCPIhNmYj1wudYaDJpIpE7/DSDi4tGVy0KOipGnwjZJkL3Lc5dAEIMNsYm
3EszEX/cqMI/8ayBrNDf5NoicZ6b5bZQJDhRUi8orrekWyLsQJzuZHrN32fx7Fm+
0GCODrcf8Q2I8aCqLB7mGPRvnDrmdvcaYTk0KHGlOLb1oI3EU05FlxdNS8ZqG0r/
hAyJN6wbPJuO6V1NpntNbiojhqz0Us0yp5mF2w20c/v7TTWfNrrB1k3LbJ1DBQc2
sm00yRnew+E5EXEcrzgcsrnB1oG31rCJgLWsgUi9utb/Pa7kRe+HFFRo6NjfRzJ+
bxbAAx21hi0oLpgeLjKnQ8qDgjti7Rd87EM6y9HADSyWGCg/gdkx50nVFqCYPgqM
HSvnE1x39iBniztq7ez288Df+cuRSvINsREP6FnIjOdRKMyZ+EN6l+J+yDHYfjYF
9A6QZyOE7xGve216rVQZgiYEtfQSJ3XUb86WHBzGr+ttxwhkrZYLLuL4xxOBCEys
Idxl6xepmBUEy3y06df4DaEA6HyKW6Qhmx7VojWH/kmCJOzL0oCXiLD1mww2yLoE
n4nRkH7D3UrN5X5+EBoTveHrBx8bm7bWReAySpkN+nhfKTQDERcLHG4Y5pu9lp8r
w9Gcpu30sPAFrKTV7A3WxYGgBgrJZTnqw50uBlSlKgcxy2Vnb+WEdYsZ5k1AN8Mr
OL0SCaSnVBMEVbd2U/f5wAyzcxfiNjo8UOmJL0D1W+mCa43LOsar3Ybz3EwSrl35
EJ10wKphGeFz+9m2T0AoED3IOlHGfqcqEq6QnthDcWojV7oX3kgbr2849LCQau9E
HDqTC+pQm9mSvm7cY9l6rBCW4pOxP/wVl6oYD0jDAVv0QCmLdExyIRAST2P19Jo5
/pkEIdPenpQx2j8K+6qk68KXUEiIUERtkMpsmY+zUkSzVJRfGItGdy8Kgp3mm5Vf
dy0awt5okE9HIwYaxdN/LhAWOI/kHgPS/JVqMEvIIu5WXxEpJoLoFlavBEk4hfd+
Hw5ZPD0UGRzmli1Rbk2g7OC0G1m36F8n6T8QOuKhSd6hJIxUydkTzx7f1oKHg6sg
sQP8ksb6FiacV6FToGGgECIgZ5djI8yqoL1TGnPJbrCZjbKShIOKPmUbptWHBybK
7MDLYADSHYANEnxiAJhqW3qkVEv6nvWYhhxqKet6DeuTP0M7ILtdwlFYTpkdPUS1
XUTIdGc0mzOx6xyl4kyK5Fw/0NunhkzbxwR/N14F/NEBxagZb/lmIavbC4Vp0Vjv
fFLUej72upvnLtSfEU2cbXmuF+BuWzuOBEZbD9BGYkoTpH5/OEbhN6zckl+BWivx
YkBeKunAFfmG/MCP/E4J6k32pIisETvmpQic4ITmQKvqehRCyZot9XU/wEznjmF3
aDVwRqdOsXftEyjbnRAibS/RTqhlLjwhfeVRXJaiddb+PtZT0EC445Vls4wJurwb
elJIBCK+M5FnJYAGq/+DdzZ78a7LaZFmmHR2davbgj/TCcEfhc1ltgnQdiGVcU0c
+7kDyoNUaPlk7HubX6TScmBFAJG4hnGN3mhQ4LOwsfCRyMjNiG3GTcCDvh2q/Hvq
0HUEIw6a3WPEx5BmnI/x44NOjKNG9werfS4luU4lsdNL2VfKi69hCvbCXTiJtYJL
A9Ezm+noGezabpIxagPm8IKhENn2Wpv+bZ+ayZwPP3uR91NzzPnWrDvG8gm9dcAY
zZiBRGxJis8WWofxg0VGTbYrNEgSpzxlDrH/0p5pjID8YkCn1CgEn/sK77NqlpbL
d4e89sPU+ucl4+Nb0C+5tlL4RQzU+HK2QIvGxQsItZjmLdB97y3CG2TKzu3/WrlJ
dtVzb0mqsEosXcsW/jc0suKPk2NLn8JK95P1vO+y9kOnbssKF0m1lNHHKMj5apMp
+tPp0UDF2BsV02lyAlG4IQ7gmbV+JJO5Y4+4EwTCq/ko6ImCeaCPDWTpZs2Do4p/
UL93yeHin1P4NoMdzgQZFkbBg5RzAeN+4oB7i9lnTZrGeXjnb3YqwtHUR3ZquC4X
sE83wUDDr1Z342DxaYgci5jOmT/tzjPBK6FbFBvwobjyM8zRua+EUW18K3/HI+BT
SQRE3QlaJw6PPptBVfY1Ueq+Td/+ysRMnz4psN7WciTG/PRYhn4uasj/nPqXDruG
UDY4PeSpvLlOpBVSh8WN3mMsB/7nmizQlbhUx91q4F/a4CJrHXWFaYk+uD1/sJ9w
WElsbi/G5EvM6UBd3WHtwP/Gcn5WSmPY0O5gxRvyI9fP3CjHDCWfQ8mahhHB9EuB
XX69uGuN6S1mWK0MdU15FyPipN9PQYG5uV0kRcJfwrdjmJCzq6KTRcNlUGcFaWHX
NeWU3wPBxLXYmoYpUKsi0p2lBEXsizFcBO0XQzQW87DC5i/TZSy5IQzwUv/i9cHK
M1O0rNY8UWpU0H7hiCatmvl/8SrFmXqG4Cs0qh/iYrTeb32I3RS7lUqOWXKOmEXn
u6qgBU3SHWivD14wnQ9sSqNS70BRr633+czZGG0rioUXMmt7Z85oclyUAvzrTjOh
DC0HyfdUDiq+/x7TXjT4MBCuIzkd8KGaWisRwK+zVuad5RCQS5C7KgQxmPjsUSE+
siFHdKtPaSA9bPaa1UK5ha8+uiyNZjy2J6d9W+/EFiPfIGtfzT9vfpAmVAI7pn/k
0Ka94V1iOdrZqm8pIoIJZG1haH8kkgvsULH+izZch9KpohYlPehj4t8LKkOuAMCh
Mk241qazLZvWtFvmhTzz7NpK29Lx87HfGEPnvMXQ4OlPmIQOeKqrnZQxAdB1Gd8b
JGiZtXLyRJaboe0GQTa/SfgeCzkPAIPrarrV1AK3XoVNPs58tzvcfoClXJ6vpEH+
biiBdgTsVyElRwYAIWVd8UrQGxA7p44GzHJgWPZtUwNLlv5zkspYpA05QvfxELQ7
`protect END_PROTECTED
