`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OKz25SPBEhQB99i2ezMtgHPEfahFBH9auVfzJN3wOT7CFN7ZXV/JN0cpOKrHhM6D
EUVOwuyDO68v8casXET4Xd1iqytVRXsiIPLbeiiNqbLrTOPIgDDBSQAIFvooxz8Q
jv7iEyF/RDR4Vm95wnclYQEbmUxW9T77Aza8ScrYyzF6UQC8QuX67zfIPWFF/PtV
hdzryZID0V2SufTA4s1ADRs2IUUZPLKQFj5b33cgmayrGqSlYwj1k7B7SIuFPEa9
bVshrrsFuqsZObbABMafjiG+GLAAtsMjSPZSS0FvfSlwVMo+ON3NDVmmeqp1hXGY
sJoDzUuRfDB36o2dti90e4x9DvS9KcGET8fOTV6OzEbwvSj+LAAAL7YQWAOdCRjo
PZEtcXzhPyGLvrThEz6elvrwaWuaGoj/qMC+8e7dg4aMmlz6eRIFGA9N8xCARKlY
X4D1yINMDedarJqq00IZDkYDMQEnPe4zgqieZD7x6Z2GWIT6kKhN9xKvB/utVQin
k/gxZJoqOBZ/EEJRzTRxpQ9c6JbQ+ynubaBj80bY/FwZORyk5xRQaxUIn1mgNFeE
QYQZoMQlH4OMIWRzJbX1Heud+I4AbJGdO1PEdTE5Wuo6eAEJmkwl/kER+2EnL979
NetQcTblWLRmJmFOGsf2HYXwSXYJ7w8qiH5s67p/M3tT2RC7mTVYxpNBsSwNIL9M
tWPG4u+rz9cqrKEz0ebNREQk/YMGvQ/dODRi2NwlZYj9qpKI7JMfUPbfb/UHm8Eq
BkOu2vdCJnE3yGXrqAYKuzIy3OK12bqnZo7zH1LCI9oJrhfCWxDW0yWaBRue/lC9
BHPQPvCjSvc4Q2Ezh/zNj2CNPVuVDqmteuYLIJlooT4vkZOOiAVyjNvaDdmDfAPK
hb2Zl02eUmsltcrxadAmfEh9DAz9tQmVYfSU/LiBmOtiuRD3Z2oOPaB5CLxJPMVA
Zgxv28K2E3r6xR9yd4Vza8mqSQtoas0hjiEk2f4LUxsumfE7AIuG/4trG2JXQq1t
Bw5BYyFwV4bWrKuS3SqqskQ2p37TEDkM6CG/5mH+cMInLZNr6kAapJ25pBqglEcP
8NHNd+hKUGZih62+bDy6PbGVkdaPomGlab/ph5Z9MK4a7rV45rBg23532LKsga0C
9RoOXN42oVy/eFVHMWPWkLt/nf/2nD/f+eFbZYBVodcPUX4JXdiDxHaBj7+rz/P0
+Z0iWPYZiaTN2pRZLPSBhtFIMPts8QTUB3owywg5z9WpD+lpH8/1EeGdK0gXjzDw
lB1X8DMlpfBpYYUFzObrSF7c9tds0OoqlZJYu0B0jzYGX+owMp3SRo0UFEQYrNwy
H7/w5GZ8qMgiL6jzxUgxs7lnOIsISsW2rsbDR46Nh+vFEoZ4yJKXL/AMmpDXJM4h
4FAlggsfrWh105DH1DvikJxJIbxMxG0l/2NcOEqlBP0xmb6G0SWoabUyvza8Ebgs
f/6twXTIgzJnwC/sgtCzmd3IsbTViTepeGGsGLZb/3VRBV46lVVlNLD5uobhkkcE
M+BvfnXMW85gWHmtdXShssqatznchiIrrybzWveEHUJJPFwN4Lx247NLiH0n7N7N
a/2HWuCzss0fVzpGc3Lw56U/szat3WtlAcWJtOPgAZwY22gi0McLD5dRT3f8o79y
GD8rtrM+lXtfNPlt/yG0MY56KQygvAHjEu8Y5KiDAaqCnnn1Rh76wFhTlIHGKvDE
6G7PeDBRNrYIhOLt5HYG2hVdojoFMY+19HsTQx7ddtK5TSCD/9hOC6QyhuHmBTnE
H3793cV1xiyJjdChFtD3uBiCq7o49bn7p0a06RYLBVq1mGg8bJZK+/pc+8CcmMUY
J5LppP+OB+tiqQFw9Kv1eFJ4MHT/BXXWQBhkuCmwPeoXBf6hX0Cyt0PXZLgfvQKC
4U/qqZCze/2h8wzhspYu9dqWZ/GX1LwdOR7OKjAGi/yjDSsbFpYQnVhxb+aXOrH8
zdXq4Do6fwtgkisMu/v5EhOssKb/eBZn4jyNxqC3F4X9mO3mf1W5mamPBSdP/bAG
dpZl8tcGZMDDEltCgTDJKDTCdT2YJR1G9H5+qEE3tukVHEAMBOhmYk2T2QFh5TI/
YlBcD6NK2zIjxoZP+pfwonj6cYoqn0wkPPgzkyeFp631CEeCQNoUQzZIvoDuibQH
WYf0O8Qok7M897q6DOr2KxEpPuDI90i74hQsZBkGulNhRrTgX24nxZingzumVhVh
2Uo8U+TrET5v7XCGIW0oyq6Kh2ctZFppNaNa6g+TcCHmwv/Xr7l7SyfP/96bTvUB
wA8Vd8zKDMB84Xp5yv8aRhMcpfbVRgssCktW37q/VZczuQZOdXjYhk55vQ88qWFz
+mSnXrujThjt+xuvCpip+ZqyetZEDR4rKE40af1AlIrNi2ZFmiGtEMv3gpZXSpug
KF0kDxJAxfLfCgNYOOwnhVoaTVwfV/ofUKIuj8IqDAWE3iH/cxurqV5vqN2GfbXB
UMgPuMpZPdg9vXMK5fz8rRpUDFUqpD3x4onpgdCN5v5/VSvArgpo8XKmYHRTr3rM
9n3JVU5s2d/Jvm/ph1EisvbNDncet5XD0dC9KZRsFRWb6BnZUNasXpEe5pIAmnGZ
SjWl6zuyaGZtgNljHrFVjirppjpL7dtiaqxNYvfGjjkIRAZX00zbN3Z9b4cwxKCX
lQ0v6Hbsa5Ex+c9dwEvJEFhTXs70QV2GMYgJMD66VOqRsw2PScBeB9ZY3kB0IESw
LjBiwR/aA7gQUacIxCWQ0T8Nys+l3m5kDLVx3IwsTt3olr4Qza3D1ZOoNH7y6S43
iX6EavLXgt3++LGHxqvqkvHsZwPoRmgtMDhag5xrYQQk+hQggd4C4Ma6CJt7fsrO
UWMA/U636TjtzrwJTijdDFQELSrgkgaKEUibR1Y2oUXPidVszoH+Fiknf8PHYVdW
zz3tIzeP0kBR97Zg+YF+oGSt6o5JB459VeWUPQlOHe1sOwLcHYpAmor/pYCNJEsb
NT30w80RPfod2MFYYluy7amaeL2ylyuvFG4ufP70flyXET4jjj9CinuP9rX5tD1d
oG0fUSIqN0eN5BVSWvmGhyNPrevx80qTyMaSdyaGwJOyJOuV6B4cBeIc6iGAHtFJ
RVP5l2Zg42NzPbSNhGrS71UmpLt+pZE4Ef2Gqy8R/j5LyAUy4lZE4TdzGAM7/tCJ
hO5FqnZCKBGClwPGwThrRMYalu3qcMh2pD6AHXuRNpLZRmbZb4VqoaJ/nwSE6K9i
WVERCW2tJsDkWMbVpPQgC4Pe6z56XQTwks2eJgaYzYqZJy9hhyaAuPCWAJIFCs5K
zTu6/kssR6sS+NTKZAC3dq2Jjgp8MCw3SxdgHV5gPzWWs9I4fEY43o87zZDcSIov
RSuqJBwleNuTYNENfX3qjhgmcSHYGxboveK06dSV2R2GhhuMXv8iQuQTRSL/pkOP
PpO113HJPr1RZUWmetp9zgvftQ6aT/eaipUa/E/jCIqBDVMVo9xbdLfZQnzDyEaM
sYOvAcQ4Soi0GkEWWP3R454qd9X6an/dDWcB75TjB7n8zYxWOQSNHs3S6BHPJY+s
tEDittuPqw7gbyYqElZwEJ/KAdnSg6szV7KiJlI7DMdkKn+3KFSYQuyLCxHHvAAM
vtdngKcksCposgwTWtLvFHTnTESOj0E3092se/0hFY6rdBZE+ErhWgx/b+a5QvA9
O4JZa5gi2xhSvo2eRTYliyg/2syVIiQk25c+EHFyOJmVLC+RCj40ZVbVl2zaYqN1
ISGYpDNU+AbAgW9pUuJJ3FvxNcLMj4bZPjaoKy6XSLetzTO/wR+kecTSKHUnEYJC
auZq3SlTbbkqBAeWuvSxHG53QJMlC94O6vANc7R7eVy7yW49/vdpK/VNFPczgxW1
hhZ4/7HI1j5/Qy5K7jtJNJDMVdLIJvJLCckTOpCmcMGocEUL68r69oVnQ+C9u1Ej
oIHFfpdFDk31kmSsXiJIspeN7CtQQ7Sre7+qRzKTyAjWT4fcq5AsmhKhcnnZHYCH
dd4x/SO2Qzdk8LSHQevkuxuS35syHhCOOGoP6SlFButBvI+qoZz+rWQn+NDzRTog
B9CVORW5eexLHnalOt18bGJWnebrqoK+yEW4a3Q9hcrT6/bywA6NgJ1YKqUEKAgJ
bb4KKndbTj8gUec8gdCIyKI2WQ9wbC9/YSDXyXnjVwQJRC9/LaYY2kaWRrYTPJow
0ESau8iRJw6tPAuZAgwbq6ukqmecTPclFXgm3S3LN5JRD5xuqAy5RA1BbUPQ70A8
zOEC0PPuXVAmFLOG8CBdiScl3NDOO8D+av2sUUjPupzHzWQ3XFHiSKI5fH10DFHq
FKeFu+BV8iPyG6rbLbxrzq0nfCW5urgdoSi9gk/DJzW8SMxVxPsm70WOZFYo4B97
eIgccN+xxNiQGEQjy8qs7JCEbxhQ20SIbnD6b3yfZznIp5BJ+WZU7lBqbZ/p5z58
fzOgYx1Gc/C6Kp7wYXK7g0XyNfCVbmyiyXnAOHm7IyBcIn0IHe1fVhxrjJi29hCL
3I49diRMf2NBDcFUafepfVnt0l4vCAAAETXANdQ45br3FLDD5X30XqVBa0fgD66X
GJ33KsNEnWtU13PKLIr1TmtHftK0v0o5GqpvQRKxR/fKPg2Vf+FpmMoxDdMgZQOn
G2E+0LsNhffAgQnWkjJTZHATv2dflNTSE7Z9xE/RVsSNUTZ48PGVSjaXjsEmMe/L
0W+hDVwgxhBFriToyE2MHC8tagNI2dyVtRi0gu+fH9Lknghx8bfAy2iMLAG5A1jt
GDwDcY0pWLmfLhDPZ1kPLyA+hUKlvYxXwTkobpd4TuY08jcXfCIY1b4JiGPn99Wm
tNVJjZXLQt+pgAz366tdG3G4rKvJ55Uz/HMKto9aClj1p0Ca7nj1KEcllvvwHF0K
cVSNu8NjZ/TOBoUXzy+DDyS4ttc24irUnGV16vkxQcRTu81+PiaTcax+Co1VdNte
fDl+EjSOMiVfWoy3sx90Jfp3YEPSk0VRctJf3k04S54ghkGCwR6rvPZ1iSsD2DE/
dLiS48xYVHb6lZREQMrs88kuCyHiao79dVmuxMnStohmn58pOWJd/B796MVgChW7
NgYsN/9xygHNbisKR8T9PHjxzXvqB7Fk3GsgWI3cEe+1+uOvsw/JqenwEZftMbKz
BzeOorAE1Bjn3AgUUcu77+h4hu+FXgbKFaB31iGi21tD8auOf3z08rUh65GbWKqi
+aKqSy0LkZzLciS2fko704wn9/8KZiuyu/KxfSs3QOpsBuUP1lqSIwLMpqpIAWbs
84b/O+zJzXt7WfCzh8y1B/V2Ld5nHbHCJCrkFNmBrSTOYLIezEoy3K9lqTDBpQYr
x5kBw34ZHx3U9+dP5mqIwgGqT9hq70RFYBex7peYfomyl5WCZ82MgMux1dSk7Iax
Umjv/iZLYARLKMGia3Q2fdxjbSZ00/mM/tqWIt9OeBE7OFFVlj5Ox9NiU+439amg
qs7T7PBdvURVSEUWx2fpJTpUWjw/Nmw7Y1ijOtIP1+pLWUA90jahIcGIhORTlaDT
ccckMaY6EVIaWoYbp/BV6EqDyNJlvlApKCugP7UaMlkuV7seDHhqzk5S9Q0jEDKZ
K7qpLzunkDiUCtGHfyNWoQ5FNWKDgHV/f3Xje2dpXz7K6Mg9SBmHmrZ7Uz+Jb1wo
vgOTaZ6SRty9UUwOBV7LOp/JzrEeExnZ6WUd5c1cfChcuSR4swEjetgxCtcASvfE
JJDPKgI7T4FNStdJn5hlYFwII9pQqCwIpSCEPaB0vbr76ULxAerY5uXu0juJwzly
niNmLK7zXu/dYZ0JtS7O5Umre/TNycyCYNfVPcKAvPSINIAhYZ9+waNVivr4XajE
hqakmRYNgADrd4NjXIJgZQWeWQ/eCwU40+qV9M+TcV8Cpk3xVUBIo8VN7ItifW1m
77KEsXrq1PlbW5o/ytjpv6po/bLt+AFBYUXLhfSU7rTYgXiPP++6NhSu9W1ISXei
jtsEwiRXT4WY8a2toHaeXbyWFhpdBDjxoq7iF6HNJOKiIwa0y/dHHAW3t7g5bKVm
efSKsYj1Mqgd/2f32MeucU2smqsYnUgnuLRddxoYYQ/RKNA+8YetptOYeg8woN65
JXXTGINdRhL7gDb/COzxSx9y7/o6ZkTSBAA2Dil6FRNQHqi7mR1ntOg8KCL7gHO9
BZ4BHqSPX6XoitOwiJRAVwoThWDYEps9v76On4kd8bLYqQhgJsuUR49qhhRhTjyY
EChN69kY5UGTk12s7wN5WwdNM22USBi4E2Tz0r4LMcW9T9DPwxcpZXY3nFRIDMqx
ezjFVccWW40uSOlW2CsnrOUI6UmYlMLTwdtpQMuFoCb3yPOGrK6gXn8S8fO3tyKL
+C+7/moQrpyStjG9y+PAZJJVjNA1kbgM4q/mXhsrsfQNd4ri5DH9ESszdY9AvCw8
iwNd1ylhrxNNGT4CN5QnCLxMp0WGYZ6EoEpwCj5PoYQrwSxv6jcrz9ngJjb54qx1
mVGPXW/bbiWsxdzcQkuqFPwyQdmnybQhh3EpFdYtOmRH/vWtleSZhXD10SGhKQ3N
XoM67oPmf5oF6pZLGCxWB2k/UQTjujwi8leUaD4XFiHM4NllCY121K6dP2QYtfTV
fS5QodeV8brDEZFwp5KazZ+nLQeddkper4WaSb6BKVqFuVihxz4IMuTeXjLdKj9L
be3enw3k0oZ4AtxIelxEPCkhOoIyR33+FUU3JQVHZoYvbxcBP8xqsrUfm9m83jj7
J5AbVncrT/ctfKD4RVy954VyNlqrAJATz0h9In2VSp5y8QagOwOHCxkB9FLIDivN
xzzQx+vwsnu28UE6Ynvd9vZ9jLGF/b8dE+c96TIqKSAIq79hcaqIV0/wuun+uzVY
lYdFe0shESsRxvcbpgGLj0+OZXx913QqjmQ6qxspvKph+WNRT++nfhMnoV0CAJt6
S+kM9M7GVwJtqPKuFtxYjd09CYZioYBfRRge/sspaR5SGuMF5R+1RXhFdwlgp6vE
Mu/guEo5YXpb0kznU5DphKBrd2aPpwdmop0ZOLNDfOQYw5wtyme9d375z+4byxFJ
rcQo4+5lvoiNFOENJWzR4oW/UZyPaPs+C//fKmpIeh/qU28GMF4VMnojwEQ/Mr7v
rMXzfY38XAxXruOX1K73OJM+9IpW09MyPrSSNVuMQDa5UHxomE5DKsNc97WqEu52
n6wvQIoU+7Odwo7wHZ7aKytFXlGucBdVH75qB7f8xVrX49vLCw8ynuVjrFMrec5O
4ehle7XgNluBBBCJFUnjHiNCrGxtUaM+GdVEnwfrCnVOrpY04dyuQ0OIwbLdmbg/
Vm4v/2YWOXMB7m3rsy9RzP1rHSsj6xmxH6a2BwYW4xBbdfJ1wRRB9rUH14PNF7ha
wo4AL7RIKK07jKQtplXy7HyKZWQfeWu0019zE58u4DA5XKvSMP61ALspmOK0Rd/X
Fl41Z2iIzMDf06+SCTYqyKBrI6T+Ox8aPV95z2p7wL3x93Vr5yRCB63iRELHhHJe
Ij/8xUWk3YwVxSVVOAtRkxb4YbsNqMXKQg8FlfFCcKZTaujWN1vU1YY3mAp/EdCc
5PfcB630gjUla3YzZeTC19M9G6Z8aKVkx1xak56agtemZdwYj0e4FqsDamx/Yh4v
aOrGE4rOOWS0HlQo+nYT8N3pLN8BzJuRNUJnsf3SS27CAeeEpfUk8jREcbVWWWkV
XUjf6/NftQoQzkD9Kqd/ZlO2u6KcIx2mR0VgxZKPByChLJXbAzdrBVPqu4sThDtM
RyTrH6tB9MYoBz1Y7vatu84XGo9ow/sig0iKsozXqCN4wNw71lwUMGuVfO+lodys
rICs1VANO+S8Wm2R2kd6RnovYIrdjMMGac33NDeR+REXSdexA+pe5rF5aT+rpcM6
TyF+Wymyt3ZAvPoAh/TuSWw13lbZMwDQsr5ogkHaeuM/HtiXOA/v+dBVMvlM/Qma
tqYjTG1pfhaJSwFVBVhkdoQJizELt3gwVOeMw5AJ2Vq58jI0BAEbKUF0/tz1nn6J
zz8aOALyZVHBAVow/HNkfisCN4SGgBwPhRGpAGTeH/Xkf4+ES3mlD1MkMW5gwEHo
X4Ey3Ow+fAYWI5ugYLcVknh/aC0RgIttuYJ6T9V6aspFu4qflGUaFr0moADn5KYq
cDzJhHdQhsuALsAMExQ4je9neVc+kdyoceSQ3Fr0/f0=
`protect END_PROTECTED
