`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SUW51IiS+Y0Ecxwmb7L6LjvCz9EfJBPWdcS4gM68S3C7UxCQJd7ryPTGkXcETXiv
phY19jBnOlQfuqfABTwNih7E6RbvbmtgXmZb6+4APhB4xS7TQ2zH0kOfV40qwpxL
dqL7d55BHCjugpBHUQzP8vMKQO08sRMMCd3AQJUp1oq03A1x3QYfQfMNQAzx5ND1
chHWMj9KGnmjf6lzCGTe7hLPT48AdniD5diX7s2Q+Qj4+jcg3LyaxAIn/8OygGZ9
MKDmfuTQQcVjYZ6qahofk7dVIzbnk28V9D0Cm4m8KXajHMcVfGqcZYdeT6+TYXcs
oEaTWF+ehc5Z6gLh5ljaKrGEeeWhmddmw7O428KNXxHSXY5mI7R+fd8ABlYhJ7m1
mQlxHFzvmzYuesIC/xJYOtNZFBfXG4o11PUoB6LcE+gClLLMZ7Rm242Mw/PDLReY
DyzooZ83Cz0YhlZBDEj2dreXYbXVrAmA/EiR63RUU5wOPMhTvFYJFVLcXMwSUia+
gClCIB0LsO08/s4hLKIvKjsmMJxYo6azj5+mWdLlsbpMsGPvSZwbJbY/572mANIf
lLRHxBvh59RXhZkQlxwzEL+wGQ6matvU6M40tnCxvyf6QePwgA56Pg+r5mre6Mbj
MoCjZql32B/cPrJXyLLaEQ5Vjh1UMMrKlmPeS072HxSzHOrwRkYQ14sHw+72L0BE
sWPWFtpsJc7jnWRDiR/qP0m7fS8ZC8hX4q8UJALRgiVN69iw8ESr1+RMLUbsBFM2
YbSldZzenu4qZoZN7K3jBpcpAOgDLJ1gCygRMM2GS9FbyLoLyd6581xROj+u4UKi
yo3iKv+wF9c4aM95jRioiW4bx6xNHDXdas2Cs/n2a59ZaTA+UigRc1YVLffY2/0M
di2LKnWUCc4kqCJ8+hbMT+L3w+b1ImDqaaTKeJuP7Z78MQ3S+O2hxx4ipsDRMzBg
AQBbo8hngcSuWDnDcE9ojY+adXau0EB1nny4GpKPj09S980nJp75VnuXRkaor7Ei
FhjrNn1o5f43Lx2cArXG3Lo1oZzFGaiWccle4BBdu2L7+Tys9eo2zPrYXAf4gXWC
piK6tWb46RC3y81RpJyzIQyBYlPNpgbcz2yvG6l0ImtMPftbUrhuV41oOQBZ80PI
EIyUR2mvT4S62AR5X+O9BuQtBUenwPTlRpeD0aokS2uuNYWqcB/3yazqZiJl/gcI
aF1ZV0zoHLoQ9wdWjIZjSx5hPPnKJAUeQ+D7fH4Kh8JB129oy380oZsMdPC0tOsC
YX4hzpGi6KrmInDIdZxY+4UzWESzwJURCFwYk0S43/NSTdA+4YRroHHXvhKgSKgr
knS951RhVcehaUUS63DcptiSnlZDAl9bEdORj6IQoADyen3Bzyqaqp0yryaGMZgW
g1pC//AF5Jsrr37hbcjulE/QAH6TYsS1ob+vR7tIuTXKDpbL1+KmaHbVdVIrqPYe
PTDdBdvsZIQGe4llpgFjCM+wvGOzd0HTERsSMYYkQsKVqTfhTsaJMazNfkybKs+P
m0XH3DKgfue2P0qNLNzpGHgiENXOnS8V+SIXvFlUSemsIR08sQTroveKPhX2ojps
ol0VcL9D2BC5lY2CyGVAS+BWFbfyArVIlSP9a+jNuLc7Dje2yJhY/kobAbEm1PP6
FYFH+ndABDujtNj4EY+W+Gp8yA4a1TZiGTaVbSL6vM0GJcBnJfkSjlUJ0bJYLnh8
uLn+nFTkRzk4+s/NDmd3CTQeXC1197FlMTeOa56nqMkKcY3n9BJ2aXa72IHpgtsq
gtM5ymrNK7NEngDQ94dZ/tdSbWn6YvX3RA3ZnTlsxWQOd6oZulHeZZ2Rf7T/F2kH
h6Ej2jHJtP1hgrUuHBBbWLe7X9uo5CDKjdmpag3zcCNpUH3cfWd734yTh/ISgqeC
BkVKeM0iBIwJ4E7No7+RHzxYmibekGmAAP38ziL3xfd8U8o8i0+9euGPjvRKdCQl
fMhIqTlOtEMg0VluIBTGWTNm6m8K0vwGEZWMNlqJ8YeOjUvqeY0MO6DVTRgUO0ea
UDZTzEKTdlEd9s8cWkTw73t2/gdTHOvo1/S0qSbNX9/4j8QoOcbIqOOQi7UhgN6N
oJKfOa0vQ1NDNjXjsL8VAWAW/UexBWAN2LiKLYPO+r1ba0fmG5friVTpZ1YSE66/
BhKMdtitRXN1CdDEs6OQqrjKX3AGhsZb6+KlyN4JI6Hvqz7eivo6BiwZHUa0ss1G
sMXFbkyaYYmjSikVshbV4O+Esz5o1iTEYM63abBHRdRBT38weciYF0G/33wA8auD
GVgmVRgh3CIYLSN9ggyHxkxUyT9po4gKRc59gY2El8gVAvkntcksmgAgayI2noXA
VF0+dpS71TQ5lnsR+l0ivDXBrbmn5J6zhOnnpfsqbPwkevRYrCRRZ198SdmYYxAI
93+XCVG30SB7jLt/xawy2nqNFyZ9Eoz+RPNNCO2f9BhP4Z3V+OoGZetyBixCnfgz
QLA+5lU0vMlDs6LheJA9Tmwrp79EHD8a6oJFEEZe89FkSvFSrBYg/9ObqvI7h8a2
IfiSH6+B/CehiJrLhLMxjft9dhrsiBk+xkLCAzPTMnePmX8qwi1ITBGxc1Ehe/di
wbHtO8Ta1OQmdZ6QbJjKEwdJVVWiH9a0cdhNyVhQNc+NEFdazrV4cbf+/fs2ovJz
5bbTvTyh/uR4l9HHsm7RHIxtjZF2jaC9sfDRX/uBUdbxb+TKForm/ka3Z1W68G8R
YF2gV6ZcT98L9OAFbeKaSrQYu8U5OmPi9OwrkLtRQ7ZRNHdIDZLJD9nnoAn0FCYR
Bjf3ssjmmohz8n06y31I5D6kEQK1nRup6mj/ADXjdoRDbSR/tH+p7BNP7hAtS3Jg
l18wTfPXL8aN98U04yd6OgA9QXy8LQraUHvU/8hf2Ih0vG7xRfFHa4NZUXnzl6QL
HaTeQSCkzwLgqIlGbOMi1SA6yeHwFlyb2Wbxd5mNTYGnwCK/SzNV6AK5G+YTSzNy
uvpbbuzuZ3k06yD+6Zo0PhIjphs9UWc/AI8r4uWfsmkD6QeUUMj1fahHC/E4lURx
/0UzQ6KEA1jnnMuvhp8a4xEjr6PwNgp5y9dqQsdrs//UKt393lPJ3FXVW0RY49vJ
Zs8cb0nmyRZYp+6AzT4rfKLk3ZUgi8RSC2WEarpM3MhLy9EFl0dVvorwTrGt/yvL
TV7T9OLcdf9bU4f8NeUqMaPsDqzYURJvA4fkgI3k2I2thoU0AazvP2XJRd8Ulwb9
ybSQnMNjGCGIBlgqcadEY874AWnnJ3hNJlHoN4Szr9R+j7sd0EfV7D4/R+rRdRfp
aaMQQcXk9L3i8heshvfGJ7cNDguKP6E6AwhS4Bu18EH2J9tQciAM0jwrnXoYfsa5
zMEtJwk3GN8lVxkNvYPsMLzgxEwsUMTxb7fykaOc7EFpanDZVXeRY0vTKY+UzX6a
mIEevu+50zQAXWhtUUgpT1M6LHKKKMjF8eYK7cYUngpnVN76nHkKvzOf2CT2oE2d
uHyWtT7dksoo2vMIjNbIW0A0DPQQQu/zT+BR+x+LL33yWb5T/JAI6gcNBWWQ7f2k
WvvfFtl03dHkr6idX4Dz296LuOW27mLHdT9Xlf2fZbHQ1CFGRXgqhM8F6syXZBnL
K1ePw1Pi/VBFWKq8MXXcG64rRiOUFMnCY/GZ5+qbmZy2fLXgZq/u52PSapXFlwAe
ZJxXJ1hxI8Ry5kOhUhhUB5QO/P8Ucx9eYM5y2dQ1IRcC53czqmKecr8CeAuD3LM8
xiXoDmxoSDa8kv46308NPL9gZ7P09htHAmoQlRO0QRhQBpbCpNBAolzNTc0O+qsH
soJe+GHo8vYiR3x5bGf3ZHAZ0Dr3O5GL94U84BVcfh7OO62G7TmChq631Nivn1GM
NNtALFox+MGLCepge6fboCernaodoUGol3pYL10cF6RyU/J+PA9sIXlb6XkAtoH0
moVpqUgStyneBkcLushhzWEqD3jibzsQzVj39/ZDjF2L0+LqZlZEFwtylEtqW59u
zteA1SyokYe6HzLyD0lEixEtFKH631/zWGR2qV3p/l5Gajtcj8wTj+bVTQeX6ac6
FOTTGyZOnGYKgSFEQ6J3DLNDN94zKwZxUrAegWiPO1IMwTuag7Tyo39BW24mHEZ4
9As2L5W4OvD3q79y1KaDQ45lT6FMB/5tGK+ByPdwRCujbbiwdbEAumwLQyY2voB6
QtgPWomXbAsmkZTHXP2MlqMBCROo3srrYxo6LFFkPitnwkixX5reE8gv8yKejGTf
LdJYf/C+hN0cJrE0slYeo7Rjpanl4vz55CGe+oZTg+WbjWCgJGSEaaLrXbW09WX4
w1zL/mH4yMoGaFeIWPMKLpX50Ejpm0PO7+GCtdm3ApF3ydzRokvFWX/FJvSqt0hK
LhAvEXqstNuB7yt0tji26/APFyz/Eew7vz3OXWYO07gMGmgRcUJGKx7UOhGpluD6
2nXo4KkWqeW8JCi36of9M2XmzTYvC9SbnviGaUb8bfDP1EK20kT1pNtVttu9/7pJ
KSYt1jSQRCpI0wtkeBCGSUZqmiSL15nkoRtKcBbhoOw2fqWPv4Jpq1F8+OrGnRQJ
ZEScC1ILxSH86tghCcdZoxThOZejYzBOGIy5lgX5SCBgBjBeTpfZrvG2PH8DMx08
hrNKY0oWCl7QLVH340/l96g8AlxSoOmI4ZlTVeRCALbzFz7QbjaiE24gkxmHnZDT
7gqcqzoka9UGQUonxqudDE8eSIIIathhjach1bqHgXiemyFD+hxIx9uQ/sEpnAQX
BpGIgnktqXpwtAthP0rFh/rYKIvw/1stYDnJT9qcaCD7/oH9YvaGbT9Sr2nju0Hl
hFpTx4Og/N5ahNf3MWi93GhpqPb2GRvP0JmYupJMiCPhgZsphYfVqWEx+lg9IEY+
AfX451qc2VbM+3zgu4ktIErPOmd2TaKKrmLVfEq8i2lBFtH2mTaBmqGuUXBVGls8
E9OJx1cHYN6YBqJGJk2x4bbymPa0LIYtkAtQnQGIIyb9Xz2b5OmeUmpuUuEwvnbU
uZg3hDUklXVhnFxIuyYY3D9IG10Xwwa8bWAoP5vGOWt93cGFzVbOiRhqjOIYQ5Am
XrqK6mTxC1lvvQBuEhubf7M0IS6UkMgqoMqnu63gXmlIVK6v4ZSm6UYGD14kac56
s4Ga7cyFYPK4kS2lBGx33y4AlldjY9bg7nR1JxxQh0dcb2Pn8m0F0NgHFKRzxyMA
PSj+oU40i2mwheoYTMCbG3ZqlhYyV4K5Y8818jikJgUm3SLM1c6En4CDNxIQ8g2f
25LhrXLBa8nV3WMP6Ud1r4GM7k4yoMri2BnyZpjjORxtu5OncFxBWdN8loqHAY0m
BYDgrdPjBrddwRHo9ETudI/XRfLDHF0JqPC3P4aTbBGzYi7ORd8mSke7jRl6PmoV
F2EaD9M7NRKR+TWE6DVbAAEgjPRUJcTAkaaOxNe9YV8R0tTW2QmR/wxmI8z9NRTJ
OcVCxO2o+YdUiBY2QRl9RDnSHMRyeQwkTBZnISfY6EqbOW/8cMFpujYqkCIbeV/S
4c6Qbhs1vsqS3/w1rR/wAOsBZi/tzXNp1wbh4UEQ7FWD/u7TYiTq649P9HgqdCl2
jjwAQbljbdQ7RV1HzRLiZgTcVeFsM1L80tT6xlMRvphRSAbvWzeTuy+TCCVIPXKI
LIHFam0VtZMeM+trZrGxmQDvkmbJzHyint6k/f+KcvKLax4qdVLKTQJuwt0Tx1/7
ksv0aDoZaFRNgUe+MxFZ/ovf+zyXwuU3lEEao1QFMR7CNchGdbmqWrMIAr/+LKaI
RsSUhAsgI01/hK0qb33z2qUgg26iY9eQPqYrx4cfe5rxVBCeL/EtvSsQ3xmyb7rY
JIU2c+kQ93oYzPxxH/uOyy5LYZUK8tUj8iL1+FDXPVI2JGR2WjyYRnmWA4gSxjlK
9QP2KlnymNbIp/PvpPwrRVxckNcylkk9/Tzo05SorEUOR5GfKJ1I395gC5A1U+za
TAG+6/XRt0BcMMJFg6Z67oxe04ZIhkJ7gOiWbJxffaf/ueEs3aj4k1Ja8IIeEfAO
Kq4Bd7CKbQ6qIaEu3LrwDMjgSyzD8hrDlxRTj9Lk5I88EvyxYHYo1ftWrvLdVyot
zTEP6D0aRRH8+y1G53W5j/qGR2AbtiOhd5vLvI1Is6V4IdX+GtWC3KwtVZ4XnnTj
JTHM1is8i55QXuiHz0/VuLYDvEaeSIMQWCBbEeYfj8vrZ3bXkkSvMlKHXoZBRAyk
h3BlOYTmVyonxBxXoUvIGzkqFulbv0aLi51BYZzGNx0rMa8EP3K/h9XW0PXW9jPU
c1q3GWrInlyyI4QGRoZDX9SKt893cXFD/9zUA3NLaj4XDp6s9nNBaCqzKDQ04lvh
4lKgHChIsq0vo4JATwI1yZV6wiC45A5MlhxGU5opE5o=
`protect END_PROTECTED
