`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6XOMO+cbyjLa3WCSLedcFe3mJba1virtHQKluoPvjAbdV5p0RviCR9NBHilWwa83
zABfMi+PiKEW66k/vg3PWu5SisLEpzJ7CUph+eYUfjp44xFZBpGGEx1yX0I2ntMT
GqbuFOA7gH7YC1lsdsO2CtpjjU/IIjz38AGJH6nSmI0/qUbXPeXlO3mWTVGwkx3+
F0FRjxB4+HLEabUrSzmXgWhECCPJEsoYPIZRdE7F6azothqvHaZMIHmuciSCR2yH
ELOglvM73ZqMwLQIRhFIkNKCV4zIz0WaWASEGDaMdekvI4h/h7q3fT5lAlWf5q9+
ohYMKYKFowz6bWMt2MziYc7S3l+GgM/AR3sDAQa8tH8RR1KnW7Cnhd6fin2txExr
6u47SEu9TKRuPlm+u3fncPIUO3wCBQ0495w4fW8qSCUFJRIC4Wh93y2MCumvwFrd
mLt3iMnCWhHz2cEC/GA6cjMUeyuMR8TbEDbTkjpW1pFLtGn4g83SvRvQQPgy3n7b
K8POw31DbY5pkRNSNpHfqCMoRQ47wHusU6XjtYTzzO7FynHjXd0d1Rq7VA4dGGKs
gg2OdRejeCCAt/lxw4LiSIq4uSvEE+uIFpaSQQGz0YFrgo9+FhP06hBNItbwblWT
doR1N6wrN60zuRxnWm1oXZyBUiLEpmcnMjKh/fGhH9LJQKIrhCjoWvAVhvJfArEd
4jk3Is51grolNoBsP4OgvVwf6rvwIVw7TOuPGfDpJSu1kh7YRMvKGCph25OFz4U4
od39i7HirkAovO3xb2tCk1SsQrI0leAsFglKPev6+x2w9Nl5pMoGE57Mm3ojqaJe
OwwtM6Ni4YCKhtCINF4mceo630gpz/slopEinPyYvvAC82bOYSui2hrhHjhq8Kt1
S7rQOedKi9MtnKpkn1QiAzPe2Mp7q7a2b/lMUoEMjhsZdFq6kLwrCbiOGsxlX6Ju
RSvYiobdP1uzAeBTunmTmV6tYMt/E8b1flE843GcNFalodJfSUOnqlmc01RuyTBs
y5POD+tSdMPDuD6Zha2tdMvgOvvAOri6LAqhBm/eYg3L7sRfLhE8YtKUJE3YPYCE
bODIBu5CKnt7Cg7xT5I1DwrTSi0rYG/7B1V8ou/0neyl1O45godeDSm37254Osr1
gAqYOsMWhCpjRPifPzOmb2p8/xhw/XAbyldNOZZ8QZSqEoJJetx/jtcErFNnplrC
PuawmMhPmfTiTEi++/ImrePom83aAYVBvCz7OfuAduCGsnqBj42TiZNvgtBAQOnc
1t30n6CPTQPEOtuj/ApNDyKgPCliMMu4y/Iinj+m7++HJT/OMcAol3Nb0BveB59R
yD1vQuxdKJWmnFT4LG9R57J6kR0q8vSCs/waj+7C+sPUyl0rA0Ye8jm+o07PzkYw
svjAbt08AYzMGW3ro6F5Z6PfDitqqW3dJE6Kd1c+BIgq/+wLvKd896FaxRWut1Ll
Mt7x4DEKsNt2Y8NmdHtBuw5xAHGIpOkSow+a7NbmdpQ3I/pr60rTkvLF9bUWAR81
bAyCaoKEzCs6sL/marYJruTz1IOHWuwEsFyFYHLxSjWmy4+LvmCCX064XzEfImwe
1pZ5Lzad/3V6iE/+0LykA2AuOBZQFoWjoZj3vKvP+HhBtanED9tYiyIc8TOD2Wcr
AAVn/uKUIjLuPKe5V9xaq7iathRVjgYfHdBtiZya8k4MTmbtxk7DXUrREwufGnXY
0/jjcSMDu5sRZgoAFo4VbwcH4wBxLc8maholzDQh6zmDk5nG5RQ6sVLqyTHZe/Bf
Gqwv2ccjxuAiq9/h7D66cqk25MiP6pOgZMq2o5kPeVAN4QwoqK2YpZeK60ZqGaCX
vUUM0OPVEsioA6V5KiDBYJA3JffmgSogvBc+79UCru5gsa5UdINYp3hdSheREP7f
OXfCzD2z1IGapLmM9LebvCvaNu5L/xl3dRwnGxlx4yxo6h4uOJViqmrgrTYx1e97
BdTFV+Vsa21LRI1YMPcdJdzG/o7gzYCwZ6bglZHfV9EMjNdAyh+JNn+zh+4SDWFF
aGQSwn9/tvNkFVSGlBTRI2Z1vTJuUayqBv+QqQL5bRY66vHxhZwglkvRza60x1mT
4XLAr8LUyt7N3Z3ClzMlsusbOckYKfjRB1w3UPAlYEbx9gvUgl+Tiwc1McxH1i1/
P/9bzd0LkMMCzl1xTcGOZMmhuf/HrLqAOZc0TuUyOnPMve+jkxJVs9XwLMOy+Dpv
zs0erupw2TDMKCxIoT7VHnBXhDPyRQ7vaZbwm2uFvJRrA+tSDi7VRJcVpPIXNT/I
8Kttd2rECs3mFqEyFZwLgvjHf63kBT7Xwta5tnbij0EtcY3sb+8w6JWpfR+vBMSx
XLOdxc/rhFPZwX11h6q07xrHKPZGt5tKI+CBgZ/AT+c8YlCIlqVi6/YW3RNXdPuf
VNQ+dwc3w412/hL7E9rSgC62o7YAp9Vv1IB623VDMNM=
`protect END_PROTECTED
