`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A34hcSNSom5NNI40fDZB0gFPrpSDkmXjrbIt3AstnUWH03gLAPpoG7wTp2/5vvF8
nyo+zEfpWF5BuTVUUXNtyen1q9BK+2Qsvs9fjHE7CqcDPsh7xN9Yo/h1bgtOaTGj
kPY0tKTR+D5PsT3091tIRuMFYnWANT4GSwmGLSKcWIBune97VvCTpVDz1Pv6lRSP
QWHuo/2pn+7IG/54/BRmS/KbTBLHlmCuMhSpnDhtTWVuWSjWks1LoRrEM04fwlSX
nygGMxJ6Pcx81wO7lDx9Hm02Y+vyyfhI3y7uzg0lwwCMm+lTYWOWoXmtHFn0p/TM
q9NAzm1k73676AybX/z67zCJKV/WJDL6MTEJMtZcSP4u9qVAAtu0kkI0Z23NMMBq
ntNVcIKfBYv/9NcksgtQaxlCVpGdQejcgkgmj8rQrp7EbHrI0pDzEV//sDubHDN5
SzOjEQa4wxXDlH7E9Ht8k8k0r+ZZruq3TiSG27hwESpMm2RfDK/mJIFBWdhDxvg9
i5pWVP2S1Fa9KxRtRe36UIJV4Legi/5B8wnrz3xZO8RBW9+t9CzVpy3cjJe3C1eP
wkB0x/2NxOUm3RnVVw4Hi3ozFkENLCjCAdsbp9ZxcxYbff2kUGf5N+VJv8L+eEaD
42seU6jjiYpTlc5xuD9D17Av74dLmC5Gm2ws7Av1pFb91GJUF/WCBGKYa7P5QBN5
+B3MOAqjdagA+r0IxbJE+0rH221Z2/ICGFi50rWWUcg07vCBCCa814HhtU4qjJTe
iqO9Tq3zy3vq67J7TKizf+mZvwTYlN/FZxPbVufewGw9rAiLLyQO9PghwLcaAlew
5b18ghQzjzSqNMu87i966W1f5hgUzx3b0GJHF19b74FzOqi+8ZA4f4D3XA79Rj7i
OCdaJBn6gM6YVzWHqQVrBZAcfx0IwJLpSu0oI5FrDrn4meBvl1RkStOGUBLLJGPO
QddSYYfF4ky5C29IMuNtQ0fEgkfWEAwCEmW1v3r3iLemJ5cykwjGpaPTHJOBvP3q
Q07mG40U+fhIm6cWu0H3VwK+DJ9g03IvWMamKioCbfXtCJ19O1yqkyCCKo6Ln4Ls
kihcHmbwXIU56IHKa2OujR53mltpDHIQcPDJsDZZeeg2L3tX/z26sbdw0pH7y+rc
T7h47nwhzoiNsap86v+GOJMSmEWb8eMmhozwEfUyxeErskgoN7BM70vv1lHrkPku
kpLeRjF1Uhkd9qIWKNdefYiEycm7B3FUlxFypzqTOySQ5MHMGsHj4EB/Dy4a1JV0
ziWjZB7PHoLNulfSAsY49UHjV0SsTyFdF0acdCDk6P7iQ1dKBDY2EezDlDyimXNI
0kd4R+w65dnzfGNeEMZ7i47DSQYwn6J5jDTmcb7ZHGMVjKdLDBRWYVAPUWHTRUzj
yIJkeo640IJYtexmrevlbrISV1xHe6iabc0M+RK8ZpOaWxlEXBl0tgVvLJyvRiiE
T2A/t3Hcyn/qXQlVpcZl+ZwweEIa4msL9ET6ZyErLP45VIdV/fLhCUhvV/d/bNhA
g37EK8/eVtlldQlNWmNK10kdb/yMY/KyYjknqFLphAnA+eJjTGBtSJg9kz5l9atj
naQZ7DnKWvCwNRSZxm7KK5pM/8I2SNkwohl4jy8DcIiKI7jAA8tbfceq4F20wOWA
/UaAeZFjlgFTlTvfSZa2U95vY31WXP44SmMTnycq4rG8zfeJz0IRDYxHBw2VEm8a
nk0AXGZuiyLlhR1hwEUN3funI7//Zfwt/+WNYJWZ2Z1+nWSWm9ApWHmEDp6vm8WH
Qx0tRuR9Fb6d/5yhwcRPwZGO1t8iokdrcMHYqiN/rJ9hjpZNKAKj9ZkhP+gE37Xx
e4EPBxcy+1txui/mKa+p0DJScMq9Nj40LKmE9jzUMlYvhk/BNdLMvBD3Bk/bo9Y9
zIVeL1pj97XRhAblv3vAtrf0aqIV7fdZECaT+9ORnUthjChI6inpejGrt3i2WkFU
8ZrnctUiGIVbo1VHGXKWb78tEFSpZHQhC9UkyRE6L2+IgpJxOcpheYobZ8WUoJDN
Qhg5G7w52BKmUKbgcI65TMsemvwHLcLLIbTjcYj5ABI7d0tMO4CHqq5NM8kAk3UR
O/bmFuCH2/L54fuR/SqFxyhhDStcC1BWZvgdJeX42OZFyD/o3pESSuWGz5D7EZJk
PPdyjTRG70QoneWGt0bfT22+MTpUvHnL/GNZBVYUj+ZE8eLwmsWO7s6SORa4UP9X
o8oAytbWhd4n2wJuHXCXBh4MPEiNrsDiHgz6Xk09vVyrLLjTLKLWLWH9384p864V
CIGbgxd4AbSP7WHU+uP+owbPe3PaUZLJ4uMsjmp0XcrtSHbys9wW0/EEMxA2lAPV
Aso2vCkhcMxXaIoyFqiaVfyo/fztVqODzYtoNtuKMP9EtXj9S7nbHfuc9UY0rv2G
l7Kke29dTR0U18+YVio51xt+XmP8xbRY4PLZnQ4gbuxN5LrQNKuPqiCWM794/p5Z
CrUTpYvlH2c115ojWtTWoN+uM4c4Lsp34+u1EnmKChgSbfLpOozNSS9DZpTue1qc
NfR9PFrfA7alSRlLIbeipmawhNkEFH1U2O98yAzIsqZaoswma228cscQ7sEcuEdB
T8JACkDD4lG4+agbiTPeceKoP6KXJnW1n0PvmQgrOxJ6th0EHSvuWAA5/W+8sSbS
BLOGjKmd16B3P9Y1wa3da0ob5FRje4lN4d5RHsKbNRPVKE+px1qTJu7a6peX87ph
TlHdmsdPoLRJS+xsXRpPhZam4MhayCjW4IsHb3I8IuFcbT3mrcenTFcOLfhtkxgD
Pmyh4EviizDHyuQMNLaPz0mJWHREXVdKc25JLhsoP4jYCpM+NEwIMAh7AMxkKedy
s551/ochtrEaI6W+YzMwG8FKxbyapEzyT0yOGDOJjJEB2qPaLa8wKrwGkwadapG+
+F/feQCcM7eCqgbmjqragY53xvPaGxKAeZmIVJGplBclYCpcZ6D1KxN7eTb0otXV
haW2fY+rWtHGgkD9Gd6/9atu0AnqhSyUwY5j1IjbfkITBOaqEQO6Ps6aPqp17L99
5kzvsUImBaFDhL8Gk+lgbaa/4D+wopx2PjEHIJ8idMhFQ7I0YUzNDnp+xLO89bL6
FKevAnxcoGJhN+zcice+8heE7F6C5Y/j2hHWpX6juPODd6ZFYbNaCLOnxwTpJAH0
Z82/0nbDwkW/SiZ3MEKGropOo5YnA7mJ4MSYSH0nqDNvyKAdIje7uPGPtG2HjJgz
CZC4hAPeMTU0LYBxyi7cmey/sGk6L3l8fg2Exl9XkxUjBVeI/TIoQbmJbpvDy95C
148atCGRdXlTWSw7QVRngKInl8yOe/zTESTZNdUU7cLqvqO4dAJfU37p94OsIXVy
PYcptF+yWuDA/qxohyBBGzvWNUtwspmdBYWr+Obndhwik5h6gpHusLcIXr4futF4
WwmKEVCRDxsxfABMDhUhmO52aFf3tr3ULgo3nzGpiKwjvjhVJVgD2qWJMWNyI9/3
K5QgUes+UySLF1Unt74XGZVxrJCp3NTN0nsSoh09ZVR4r4z6evB5ijJN+pzFmH8V
txLKKuvi2jc7KL9JaXKF+pD6+W9zP2ZlcUZ9uaiNg1sG3nUG7+QTsZGSY1DbiGou
CbRqhqXVPPJpZ1frL+vRSFx/WFDQSwxyA6Wx1in/Zu1zzE/mx1TC+VSSScV5xqO6
v6DyF6iTH18fSAhD0I4uqX49qhM1Pexc3l8LLKctUAEVhpcW6RCmYWgmAX8GS7hj
DUaGxTGjmYO9SarTnLG694GhMgSDyj/MkLU2jEPYePBUozf9z7Ze9gN7Z6hJaEEs
iIAn29KK7Fb7I7akrYUtrgBidiSYGycEo/NZu9zD/WsWMPk0CYC1ERNEoazYzuVU
izc9JAeBZ6cHO3Gp8uLoC3lvkW79EINn+sszW0FNCO+jXXEjlL+emsmChnQWAwrY
VGXqMHW3NuCdKTPwMe06gBT9CXKrbQbKyvrKgcYapKXrsDh0NnhoFWnjcRVsC31N
buU4WJ6e3BkK7v6uz1UTz917W8+E8IHPnxY+Vw42Ab3M/srMyu1XDi1MvVCnfmuM
0/93V1rqHdyjNlGGkSxkcd9SnE4QGdDMrLOEO5ooiW4yJbaKJCveNydtZntbAH+d
i7lg5RDd0WGnSvwhYvBlfZI1onAWY5m4dQBeyqU8dPPhWApEmMZytqDBPMfbrZsR
6kV6nhYzVCZk2ele7TzxdwSg11zboZgdjGgDmcQUmUFmVIsnqcTv5X0AnjmMM5Id
1c0qZXoGczhlUySmTptaQ447vM8ZPrTcvvjMqHkjQc66ly2watsz+bwKY2pUs/OQ
uR4sP20z4dF6MkYaEwznCOS38qEeDKcGYXqoaBcl+W8RHSWycxF2eoTFzjTg/z4Q
PULBQd/eeydsPcUzpYHEG01HEoonY8dTYyUECLDmqivY/v4eldBKUSBFIZwNLBhD
PR02WGaBI7zcM2WMHwnzqm57FASuQ47qkJXHebPdro4BdRJGgpcU9ajnVOAOcJ9u
WD73O/Kq3PDuMrXCvydwksR6fS7g4WH/vShm/QKk8BYP2shSgNLB/Mr8ypIsuOE9
zFzYojEykh+nTfiVWiPiauVEDFzCzdAyUimKRATOvDjilAhDrDkbIXJ4OFkrUI3n
eqyNsOdYybMuYs2UmDkcYR+sVdo3UK+v44J5W8mH+4UNeWHsdUEfiADMcLNX/iJM
i4QgB4IUaltoFFeyuGSpmOAIIZn26EKKj9BHOUBTRSoUK34Lp1aRCy3xH+xrITO3
lapovFfd/0sn8Pk1fOjCNNJ09R+7kKDPDeIskDJMdm4fM5tPSs/f0G10AjxSRAje
1K6GsWrNnFEw8Rglj4EYzbS9Fp1hCO0n4hpqdtW9TN8QJffkIKl/2HQziaCb8aYX
w8oR2ReX8pgnPmRmD0FkA5NBPHPg4Tu49lJTL4Cn0EqzhLh9sNqpiGvhhO8yeeU8
Q1FTmYqW54C3iWCFgjQZ9RIuCcD/3bo6rwPgeFcc+yoCNdtIMeG2MFhXTPXRSV4A
2AiQ1w7RWbSUt2yV080/ju2/Tt7OIQftkefbkFelb556g89pXRP7MZJgxDyVsCQc
wvjuU1JUScX+dmlIr3TJbRPOhvnhKf4rO2ZBjT9SXFPK27SChzCpDquyfUdRjZh0
+JKngn2k8VW5IC5HnaOANu9DYS1Dn4qolz4tFqotbjQ2Zs2aZj0cC4uEk7R2YOdR
kJaStdlPnGEYXX7J3nJPREorFUxRsXH8IKtB5vMpMBrowb0YwPi4sBf9UxLdIstV
YwB/Lm2lSaw7/KxwNPoaGjHCOv31VGDhQKAju6MG4YaXTVnl/Eu0/ztcy6S6+9pu
ZTSGbN+HgmEJDSixP2ovSKn2XgrwcINkxZ6Uo3GTnUdCpUMK8+scBylArxE9hJxv
S+t/f7CwAkN709b07mT0h75zIbEDNXlD2e4+v0ruR8CQ9C7VUzS/QJBLLfzjM2KQ
yMDRipgtWofK8o5etvkhEajbAJ3wf09uTjFw0gTDbloUBzRvqAuFGf3KcYIfMyH+
Fi1FgjGsTdrkMczuOWymqoQAs1RcjCtfhuHxUNxFJhZhMHW7tZj6Nk1iLylkiRaP
bGw5uNGy1bT50lCxLdt3h/69PmfFm3MVkl0w4sd3b/NkNVoEM4TiciUh3jRnvnUj
0dhVawRkLlDvu0X2bmE8IskdhnCY63Pbi+FJzjNUuw7iDKl3G9dwM42JQnk3m/L3
VcXSBJlhZHirbtDP2AMYeG4DZnAkWNsnkgVb/iNQXXxUBt6JxfuUfDN15tnrxscc
t4aQUhBpMmVVbulkfnKJgECFnmmESqvmW/WT/pEcWhHJS8HpiaC4Uk8ZxqgsEJj/
8s77WJU183mS9d+BClctDdUo6wxpmPNCMvaYa9cn0qvMjGPdRRU/bNnjdPw47F6C
MgSssPgViDbaerZFNXHPnCBIxqSB+nUBOCVHQjxcBqfq71lUhYmKOlfr0cwKvouw
/WRE5kOntsVdNpFJHf5I6JWA7q/DOjulfp9uRxQAtDFPT3AY2hEePFd62TxMNSbs
`protect END_PROTECTED
