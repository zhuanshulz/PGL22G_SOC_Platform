`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n40B1OMmSJqOP4SzWhWcIpe7+3i7V8lNcVpqYKY7KBAuitGr1FWLuzgIWf3tPkWk
Xh/XdARuZyn9L0q/3iJZqr98MfGjOoNTtmy4Kp92i0wbaFrNp4LlRW0ND3WADhFg
4+i0PAA7mdYWP/QtO/Xpp31aC7SocepcauZyY+h1skwOCxJwMFUqnrx5ClLS/fd+
kWLOJ6rdF5QNhA/LUZytwKiG2P1nhOAzAjGPpjsb6/gIdITkR83vbS3mDJ5oBusF
OA3Fr6gZv9NV/PAuk3KVeeBT/y+TibiL/ptv4B1CgjduM/edU4SDzzSjpXd+8YHn
Mm6IRJWosUyudfeIlXiKdAzAiW86zPy9fxy5mQ0HvRkvdXvLCHmGsfDiOqYYqRTd
4bGT6to786PXZk+IhpVhNoxUezeljS3gr+aJCk9Awfqvb1rKcFhkzxQUrhBsDXbv
nUHmyQen5UuUEy0b7sb4o/iAJdiBRpOWQlEBf5aIKOEqBlFHZfEc5SIxmjeEXI+u
Niuj7a7/Wz2QDIhYrqSdktAVBcYjVHeMRP2qaKsHt7ZR7GDPDKnBQdlF2EMLTbk/
3uujKBTmslTZ+R9ldXG4KK8x5T6BqDDRHDOCfpYMUPB51zBJoc1ShximHwAIrGfR
i03C1oNhLVO6OZZrARX1Kc5FPxfBLupctVFiehrMwVIKNFoilqwATlIDHGasmXX3
58J7P8IPM+jfyCqKcdD34QjuOlAkP2Tp6tG1nKTijMBB+VtcJcw5cwFL2eALL1dG
ShjxRgKiU4JbuZX8iKB0ObNnsMXccLXTxUr+izl4gfl7k3av5wLakvFFseskyq4c
WAwubDcBGzAWQHoT2hquzXyri57ksuqna4qPern0FyS3YpmrkeQ40pas32dUFAic
8JQIb9Yl6OMCsdaybinySh8y97SfuUDgQqIiENiANBls/alBNFemFq0BXMbDniar
p49FEfOby/BGpPckWD1vswYqwqWljTH3IfbPRp5dyeDBhrADGnOcV+uU2sYo6RGF
Z9d0nf418R082OcKvfWP6+t0406WmPVxx0znh+XgBsFGej/Ch9sTW9riv/H2RVMC
ddjut+P0O2NfLkMbcmKpGUE27LtaKqQgVLkV8yb56W7PTrvDxIJQpW9L64ZIGdfv
iyLtWRbJ1VSJbzCjdhlgdFwAXrFAO9KbHlHp3ZuWWFgcEDx1cuiHSdyUxadqZusK
DpAW85PzAE6gT79HJCR4T32sqcqu1gTusl7LBdpwT2+YFhWZNV2muhym6MDcwQGP
VDvL0+4Juu/5lsUxhX69uie9Uh6yWZWt6XL6VD1YYhXkfm2E58eeQiFBB/88q73Q
LlxpOf9/JFgSDTeHEYhv3gGjq3gliBJyofJQ+wdM7Q/tZRnEzxQcfE7qAt9ftmrk
JmVOjMG6EksEVz0nU/pD72Z8b/nMfvrmtOvM+I5VYrpbfLoApouuKuKlknH0x5Dx
oqvJQW2xkftKK2Vk7GKmLoPQg9fjWldDVMuF0DAVnTMgffuf4wq/Vz7CLaJRcQHb
q+eetPfCu/The7TcTdA5ng6+dFdKNJFLcndDhYwtJMQaWf04GfT0oOwAUE2ml2cC
EObQAHJF8+PGds+C9V1yl3BHPEao9wdTZ/7MrINLGC8zO/bTGvU4QEyuczrUxvOt
GEvLsKU8twZeXc5LwKLAcCLkc5CRE8poNF9nioXNG4XwaijRIwg2Xs1VqvrxuCeA
/5Xn4tjxXlddUpnFej1dy7ah/vnQtz4k3GnS5JaRI0VL2Zs2UMKCFUjpNNxm+KTj
GmcaGyWVUa7cLllWLZ9ryYecGv0PrSVPP8qRbxOiXebmlKVKFomDqnHdT7kooMPK
0pxJHinUTlP7QTIwD8Rtar38cQvOt/MaReEnTEldZ/PfDK4f2ZxSg4fYAJRQJPcX
RAJ0eNpKcjbpml2c1smdnEfeUNQxHLJFKvC2Gme6gzaT4PurcAxRD7nK3KSW1k9/
Kp3+NZ/Pm5IzaMWUvNG8Cm3mCF3pPxKJsaViksEmUlx9d/Ruuyt/Kw6gyWNFeTeL
fbZpweZ2660z2FmDIv3XzPulWnNWkidXIqzLvP42u/qUWS6f2YvqgomL3jYrblmz
wevAf/clLqeNuzhdRLkNdPeG14qdN+ACVQmXipDZjeQJ1q/F9TPQ/On7OWOZM5ek
fJ8YofJtwK25nOwiwA7uMR5ZCN1ZhkBgz4JxllBB7Ut3vY1anZq7jGSyNrP46sRt
icALIkOGckTv1BI9rKW4lHqHFTkCKoD4mia4KouNV76SfnXNhHbvWd7kJ+6ef1f+
X7zc1ctHEDzPMJ0GLJvhTOmQc95qzNNWWLb9CPweKWSkvggGyL56M7rutPO6zIaG
DYp5wdM/UbzDTvH8Z8e2QTGBfzS9PIHV9VIUeFiVutkX6k8MyPNYmPQj0uupsugF
6++2UVzHf3Ry5oxBJhAwK55n8muMS+79gAS7SqcZLxG+hxuNlPttKwcQY9eSs3ce
R6KFuFWs6MyWnNGwQ5bb/IRMZyBkbADhLpKrwgxY2ICIro9kcu6hsJy8976H5R4r
He0n3fAHZ8Ni+1HT9uFgHefMprEWekuqyq8zM0vfdwRbWYMn7EkkDLQGg9pO6x8O
wt+SEIMY6UDLnKYCUl61LofHVomkS9E+3+molITp/DyKnZfAIZLD9VTdAW0o8btC
b7nxRelIYvCGusCWDrzkuCqv2DB6r+UczFo2sTBqO3YrYkWDxuj4XohNs4G23CaQ
pLykzOSesSSsWuB0lNttwGca7LDDwvjk0nboKUz3d5oU/Zos40BpRr3EG9W1uOn9
ZuNzab8pqFJq2A4RBxcLnBIQWotERqI/dh/XeyVenE8hYvEPqB3VssC/VrGtZa7y
Pgp4rLHMEPp0f+2pLSaTmQEe4Y1XWimJx8YUDnr1i10ofF10HCbJO2B/uGHXoRKL
9IY49FaOKikdvq2hCiiaBjJmBlcwxvc7AlrvQcKPllGpWameoEbsXKlW3qnY6oky
HxbaWa7Hpqjf+l4gbymTPhESJpVOQM3AYU6kdwp78wRkomRQXJlbcodm2jxZvlbE
IiWOkaJXQMhMH6Ff7rlPvqdJ35dcnCYg+O+10r7ZanShgCen5dNDsQcTxmmjK2yH
nniBeDyWk1Nl830lqkvBkvJHWPdaxDAnwABjsX5BEGOO/ostuXrmU9AVpmWZusdf
5fZiNOnYsE6YZND4sksQUCnRiJ7e/NNtuJd+sLNrFlGgKMtYvEf0+EGCcCFKXg0x
Wxhvto2yShvzWLDtP3Xqd58BCl7NKLZO5zjiZ4QAvzdLaMvRCi7bNQG5PnDDQlFj
PR1M9MRtry0oEh9gVhbpBBbTT3E4an0HlhytS+YRV6n47ophfccLbuVCrqXxfWFR
+JIojTyM5KwHceMBbLCuXF4UNpjtkuG6Ehe3jmeb9P2Ns6pubxG9YnpW/be8Wsf/
ZGHF7Re2mwL3eBCvZD2dAFa2a6icJoa9Z6eNMVQ7Px2duMTJ/p6keXcWf7pvHHCe
Ytq6Ro9wrvM6mhNywCZFUPk9hlu8eZzMti/XPRFy4uPHApyOPDFIser1Wei0n4up
AzxkZb6Hr0MuvJ5q4po8VBDWLfawRaYykLBwb2AgILkaOS0FmorLcfGuvmBoY7v6
XG+2XI9Wld59Hzy9xTd6JjaoSY50GMO5UbOzVnpkIbEu0OL7UeygXNjKapk8N3NQ
qUjCFaYVq6ULD2TztqSBWLUBu6X3fAzhjXnkrbrCBdKXVR6kWCWpCt1Gy9N1klek
aZsw1Ypsnnz4tvnIAkcNy++7wJeZAWqMvvd1vRVCWxPzxPt5l25MMpQiBPfP19Z5
8A+gq/jnb/YKFFST5QvzZwNiAmkz7iGSpL/qqs1d6v8Uue5kO64H428dIvNyDpfJ
N7qtw0le36DziY6VmYCaVlO4gEfzRqGnGRDIy2HLg/OkMeLZaRnXLB1x52cxhl3u
Waasc1LcIb7nnXQ6nwO7XlVFO2o2nuHfsi2z/93bU0O8AJoQIgahjiNsQtHu7QBl
VOTOtPT/Jyh9D8v1ZZdq2v6g7YNfNPVL79ohQHhrXNTqJps0TpJxy8boJd3EjLML
02j/Th1vQtlW9RtRLk5gBn52iPIGMv5Y6jCHUT21B2qHXcFeQDcrsXegxBY71VSb
6hIZqP8SG4cf2JEKiTybH/oknAAv7qUZkVri2qPfZiWjfbMefdyriS70d8L19vqc
ixR5xUIxjF+eV/Nu0Aq/aqAQoN3bXFn4a7tqU3LtJstJH6ky0OngqYUJXsdZa4Me
LX14UGqITiIucS2U/fRz2bmKlz5OCKM29ISk85DrfxPxLn/wgRF2m1ElDiAHxbAL
4kTOTgTo6vM3rKvpKSlI0lO22SxMmtykjZF8J4Ulit3gdNNEIqIVJyIdsqjsPyVM
9MbIyzN88P8SlLFh5Lo58t3wmijVg9qB96n77SqK5/ogqRmPTlRUkLzsYVSBy2ob
vwuLc4ky/Rsx5s6CmhEVu6OevNYehgcm4p+UxAMeVMAmaQzSpFWwQRkWZU/NYYEZ
YErWOBu6BXLRSq7ziwtmD2zmYw+CvZPz7PiPNMLxjBeIDFxynC3mSfjncvBUOojB
Acm9eyC85cNfuDTVcZKME3tUIcNxyycpq0LuNhKZ9IxPr8OS3FjfPTEKRTqGWzFl
6X+1HAsW6i85sAK5M/EQYTVKT9EFZ6uJhfmgkj/mEWv5lnUHDOVf3SYwOK/0dJDF
ttlE1UbwN3AdNaLq+T1MJHSwv7P82NSJmOODwM53Zt9PudhQQyG9UEQz02RVeTb3
enAUjeUk+H5c5VJucVgBwlq/lMl6V/gN7IlC3VX/7R6C0qhQ15ifET16seipWbTD
Axgvv4D0y5x4FX7ZA5Dnik9AtWlsiedVTRtGkCZe7ouTNyHdn7xGxfkBgF7e2rib
1rZLC484Gt/xXGFCEBXkxUmmDz0GdxwlLFaLvEHuYTfINBIxC8+LAaiBkoQpwKPo
xrEXK2ebhxbdWZgKAvYRhw0FhCa9/qO0mbGKG5Jt/TosZmBMpkuByRtEatrRXwG8
oSKoddWCF21FkGYQZmDRwaavh+rJXsKLT58pQOd0hC8ZtZHHYDh7nFZ00yqV5/ZC
+jAJSOGkwDtIaEIJYOkH0QYG5ar+FdaHfwCqia3K883vOF4U5NmSsc2Ukzko0sYi
91bMSq8PP3/ZYRrdfFbyQbLbMB2Xzw513woEdZZgPNQ4tJLFo7LM10/9esnSHa3i
dou3EAPbe2iCh/fZkQCCL3cCtmy/daJDpXF7BTMVd0OtrhkCSbq/OtQ4ndB113MY
ChTC2l8oo0DaZvjK588yMUcx/8XEyLHQlVMMF8Sua1AgE+0pFCl/VL3RLuGrDS9L
yxRvxUBtSSBYlETBnBg16L/TDLSIFzNR1Agvz1u+g/lU4BDv9ug6fku0FpwXjRql
8XNG/1s7aXXWU2FyZCzD3rdqeL4jctgrYC3JXEU6paxbzTixLJ4rrLvxi4qkjk+/
8BjfZr36erQM11kx4oxYIxi0InsaFfYfS7Mxq2cbDiXYcc/UjolEBNU6iYG1aNCn
EGo6PsNZEk1rpiSzRKqYVSTBQW4xSRNK0JZMUjhuEnjKWc+eE7uLKVunhXxWCK7t
7kKC+uSOxkotuzDTmSQay9Bm4dNj6RK19VkA9JoIbk/nLRfu+M6xWLAWcqN3Ve45
3JOxsV9QEBiimj+KznGlphNn4ILA3GQVGOkKfO1BARg0BToBjGerFYhYSd3OvOkG
4Fs4wkxgX7IGrjiXTFBV9Ce8YLfKdTlKgxcChOIX+BMRdDcYKmok33oL27zOhXdt
csnOi63keow4qKNYJdSAVTUtJRjfQRoDkWiUvBpuaX75P4KDx7Jn0EzWyl9fqsb5
EE+Zosz6CWbG+ICx28U4aB4DYpzcR9dJ1PCSD039jHl4ARus6e2DGfgRarBHOun4
e+GiKJAAYvArn4Kjvf8qqlkaDCBmXNHHAUeSx3ZJcUgKbwSooQzCBDHpJkbNrk4q
Arr/dpDf/SRd2m6SySWeBaDAZMLqnJzjWJJWjDNGWvMRik+rY13XQl3OF/1y4yWJ
Amh+Dl5IR1OJNEKZofHopRYnIZ7sHZl3L1D/kkq8VmroOAqRHYOmX3bEE+swXE7S
`protect END_PROTECTED
