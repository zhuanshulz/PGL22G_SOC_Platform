`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tkzkx2KzUStMhey4sKytRuPt92UQAoZFnZdSqiBvNexP0yoKuttERVt8ueL4mbXW
Phof7E+Q8y7ZKEgIvukhKMGPIjMh7A9E+BUNoBF0xSZtE0F6C+c5iiHAu0upC+4M
f4fqP822USgpnahJRdz90rzvSjXeAKB8pgZSl9ztb0ioxmcPRmH7saOR4f0xeeWy
jc5bglnPTqldRjghB5a1YMZ6L98+UkGpzuy8CKkNlDlknJ1a4G7+VRpQRK3AYjsH
2i1F9hiLQrc66qkpeCw0iPHZSodezfWgAWdb5ojj773HamKEZ/u04nn3T8WNALMm
vD4HEVN6rQHQuREYjI3b7g==
`protect END_PROTECTED
