`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p/izcLV28ERRQXjgLPNuoCGcQJsY+x1yYJBNnSfYjG+W8E44H7slSVV5GAMc5GNH
laz5+uy/f2pEcwQI4Ek4IbQ69afhsQHS4KWGt0o6NoGTBgUsmULUDo8FJssGhNAP
GQPzQnwhQh8bfbeeuVqDz+0v78QoJm9oklbX9PNDFur2+wSgYjTo6vYfRbpOaF/6
9wBZE0W3zIGTUd3ln/c40Jvx0H9uChObboK8sUR6FHistDz8/69th1LDqioO2ORH
gz+cXzkNFU3o6i8d6iIX6mEthcNHyQAH79Am4vKT7iL089Q7mGWsuVnn3cZZ861q
TWtTuTUniGJZ91LBoJngshQNBja2Sru5Xzy4kFhnoSFYunP7F9OVMnN05qkp26Wv
cmnpczCLVoMl6CtbFAZ2NyByUVvrj0h+y+MIpf2xaHEDxoxtoxrw6k+JRSUN8Lc7
XpYwMLPWBurkIuD1vuiDRWQjbALeBbJyItTj5amZX+JnIG36CO/60uQ4JuWIt2AJ
ets6Mx9+j4JHu53VYtOetTO5tfWvqI61gnyuy7dsR4h/6gBPVU054lbN+Dl0bRnE
nAg3j6e+34pkR1TZZZCVf666QtWe4wQs6qMNR7UF5dXDkcNXSeMvpUHSJnFwb4uV
Z0hthbfNXYi5SB4A6qd3q+r/xn/18dOv9CNODRKd8lrRf5giIqprdu/RMFVM0S4M
3f4kI3+3uzmpmjSc7BFcLC5b0EfLg3bF1a3mFErON7nRaTdQcmgils1YeXhDmXAh
Z6gFkyO+FOTTMr3eSWPp1vY3AnFN3Rb0uwfp67XDSzQv+wVj5YIDxmiT1ARivfYe
vbY5BAw+83wdOefo/gGhk9sd1hBgVzF/7SROrW9WvubWUssyzNQnMpM7lRe5Fqra
/DdLnj9pChsPQq20S4rGlEwANdr7oRbHncOPm/2DUtMsdW8U9DBiIYQWFVHDw8Xs
I80oOAkHbkSz0aoIkR/VabC9q/KAJ8w5Q6jJCWXxf0R1Uyr42+nwRmt2HKGs1pMu
4xvU65B9ArHAnA2pzr/FVbkr9vh2yqf1u6vFterF6oPG43TAj2rM6OInp+rc/xvk
WTz6t8NPEOthR1kHlXXdkQIRv8OHXyBl3WhpJAat9oTNADkWibBGKNbFiSuEjDkB
/3nb9hUbFezT0ZMgfTdTuGJrYxY21nizSs8P6toSca4tYLXlfncUy0E0wEjCKTYU
bLB922g9AUXoTN3siJSw/1aY9FvGS8UNdqUlF+YwuRPeJS2ntOmojJKScsr1fjUP
USuci5/mlf/zm6k9MJFhyqG1fGSIJtMBOqEdRnHRjx7SQq00zaN0PI7VI+8yYEDo
TwlpgIrXiTRWZAa8QAeFQR04HXqHBaMGODxHjw7WofIjxWy5vP4S0CrWYjNV0jI0
o+L0TuGx8fIVMDYEwnob4KAq7/GNtheLXcQWT2qoAl1T9+0bv7WIQexPN+mQBJaW
XSYmaWlb01D40JkEqaAz0qfZXlCYe66l2BeWOybDAvRVkXxJSiUP1B4UluKn1BW2
TrzdkDghFVaIhjm5OgF8WvCmEgJzhR1xa7m9Fw50UP77aYn1ANmI4b78a24rBDLU
SfgBpTVsYBfkh9VSLDLI2FPMPYdNOGO9MJp/E6cM3aCGbzmAqVAGgeCk4cU2E2hb
wVoQHjsRARyzUesaRyGDCtLCjHCkeGzqPuOMcNQgHHAt75PsUBryYui9hLpeiLnt
vKjkh8bC/YtNNW35kbwv23UkxEMpiQpivgvtdtHpMGckmmmPUvCbyC7slKi33EvA
MTHzS1okYZTOQiYVXZy/XmLnbk2NoIofsX1J2L86jLJr5DcjX3bchFBv/PPiSH9D
wE/KeAf95+73Hl9/S8e+88sOaCWejyY9QRd4/ct7qPcLs4Es8UOrF1X8uQ08OXVg
gdRXnE6bE5nETZOGCEC4yjxEws2c5ANMiZ5jttwfdT63J34rihmtnr8bqaaarRFH
RtqwnudOkaAY7I+gOyCCqlL6yVnme4j/LThogTxFqjUQa33ZpR+mOaqj+FvxjsUD
K2C9Zh/BGzPFWTkIXDTLu/fa4RcWBNDv11Z4rb5rzqFj1mBBlmz1uPMJ20QuPHtp
CJCP9tHZdPIiEOOv8EPo+/nP0ktRW6ZxPMUUQIGK+gL1N/7T2Oxl/5+01b2Y9KyC
lbPjBzkSX5lfOdDvtNNFslFwFFkbecqKE33Fo+ITEtfZ/2JZvCYryj5zjthVS5H8
h6WeHmLkr2FBdk9890/BkwJiedYk5DmkpdWLh+DdatxVfFnZpH86jUpGibnCDphN
m6aswi/k92v808dpGNASutsg8XzkrZC5DiaPdrH2FQzIBmZ0sJ5ZM2cawVjQC8Zj
0NUlECKeIhHz/kpRyj1AnO30xc+WS6n+Q6RLntdAUDL25lGu9I2h8ZvNNfWCU8D/
`protect END_PROTECTED
