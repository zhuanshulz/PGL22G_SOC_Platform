`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pziD9MxyRvaxD6ssLHMMD+92I1mo8/y8uGgdsezpbYw6j4Pd+AgOTrcn70+Nc/Ng
goLBf7sV7yDQr7gW75foPEcL/Yq09BQpBLHF/MjDapKskVHdcCJQ0jNc6BCrTesT
dMehWOabQtv0SoQIG4sIAvmSRpgJxIE+wotvylw3I5WgRQ50I7yE9Mf+2SLovVDV
uhWBbAFW8nWmS+BvfXBVn4YZWKXdpZURFaDl8MYIUfRFrlL4N1aePUbSSqN3WAjR
Y/kLQqDqpVJxHcEL1y+LKl+CCurtAA1/9DwioUZ5/s55gG+Xur6QJ3rmWs65h2gE
AZzL9tWkSBalB7nnDN6t/YrQt8Jyg0nhmJGCxFPBc+gFEWts0ugyMdMrUJd6f2OL
7O07N/EWHTVx+raIj+VOIHdUDjU2gyfLEcwORIYxr83U7C72hZL1Qe0EJ8itb9oT
VYehhX+aPGGtw9jhyu0F6DJ3I2ycYtgRQqnVH7q3DdKF/Fu+oH/X0jL+dDYduKQQ
hd9DTLBQxgzlEv0vci/R6XA7o6K2JMyR509cgTwK3e8/O+tuwIiulpwEqjTMC/vR
DAqnlR3YYjatrnIL9HKGTzNUZmfOzydZqo0iapXLTLgLGnjAyXGt8VQgLfLsGOUp
E775WbIWhL/GP+M83P8S47pvqCpW8cJphtMF2JmC7RHeF7OAc2OIw22rSBHkFrLz
KWYkqD1TIFmoG4KieWQv0I52oz9klKDidsDn4fEI+ihW40RU+nq5JtTjpigLDxB7
cuI8weuZCUArnczBTE+cI+munFe4scJqVam3m7IchpmJva4Yw8Hha8L1eHGjNvex
Yb7wxHl2zRrQBgAp6cMq0rOq2TRk5J2RBsTNfJDlUm+OC0wu0mwd8xXsXYkieWI1
9RJw4NvgtvNmLt75oemlyd33RiN/9jyRR3KfPeRFqBHJvTl0J1CzasAgXzTNAUpK
xEQgx2or9zhMelJZ2sHQLef1z2qm1qNZhsDI+HvlMfe5xRLlmPN/OwIiGbdTJ5Kq
TnlcIizsK3tJFeA8eGitAo34Q8Iq/2hBZ1Ugl3YOkeHWF89peAy/qNHHdsQkgxbd
tq+CRz3toNoeOtMKaFamoL28pqQdjavtFescimsgZlO0LLRpO0kGopVnAxaKjxse
lyfuV+lOG63FqF/NaCLOaSLBcYwyBIJ4yFIgZnIKWs/JB7zSXMNW8DFNExuN2pz4
sgf/MlNEia0qR71OsSD6UgtiLF4pFYM8MbjHXAFotmlZNTG0TBQ//fdGoSWdqDj6
O29p/JPXBx6eQ1KGFXkPYEAZhcppFVoQeiXzZNUZcyHqQggDssAYQRdOHNaSw2Bk
DsRrfaeNrsKw6aN8AdB/DB75yaTBlJmrqTqThRo8BjeiALna1Z66gQj4lwYSanRp
g1oncd0TdM5E1FHN7s0VlTsACrh/8PM1nHXIlMojja+q6eztFscjBw875W28OJce
6nZITkxytG1rsHNRaQIockgYQbq3XjrFQopmIFgC8mBed8lSMLadrSVVnbc1+Jwr
87YHZ8wc9cjomHCntWaOOqZfCPDtCfzqAD0SJusG84Mvj0ue/nxyhssTlz+rLzwT
OlTdKQ6SQtvVtV0gzpyZHsShdBHbFsHx2mxQuoesWGJ1JP8vYxShjDLXbWk+PDK2
n1JY+3+ZCeqArD/TeXjWVc6PkSi5IjzKVt8VzvUVGaYtUcnzbnN93OJUPYMOTL1W
2cwqOi7zMCXW0lGqrR5GHkTA8atoCQr7pHC2koz89mQ=
`protect END_PROTECTED
