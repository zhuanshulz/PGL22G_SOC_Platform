`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+sKGf+hS82oY+WYgYN1O2UImjxUAG6j+DZnvsnOMfTpLYHgTp9mRq5gsKqWH30IT
wXkecBUijdtIbVn6XXGtJ8H0iS65Ci6QJG7Or5q7nuhxTZCBDwQU6jR2jktiO5hi
MaRCfSCuH+4kz8ZVR7gMrtzj/k5+lQq0PJ5z/NRMpRYSRgWGhEKw3fBqfnfkIbfn
01fCCjz+idWjQrKMLHmATvORJUXGJ+RpFy0w7mn4HqOumAZiIpO6P7XQ/+uxsAf4
kGXsRW9x1v9owNaQI8GAoJULEagblE4UWMMN1VUB9K3TlRPYsnvVhVeXHsnhbCX4
prDf5ZmdKp9ogWJbys5lQfDPNFcBse91HQgDMjZofEL8ENpRqlx12TO8AoezElZt
vbWz8dOWA7OlBn1J35+2bxlTzSuyHNWXjY2HJECjqomQxiAauAQMQHaAUzYk+R4/
ECNKzpb16VMMuzDTfAv2HwpFTKv6tR7aYHU/p8aOfVfbBSmct6mEH+71QrSgJQ2l
mPmXmJbLNEgEifoR6p/+f8TglLjiZtZiAfHQ2Tld1z15dDtfxUKXkdZAivczy1VJ
OgjrUqbgxnA6ZTqbF/jztYKkgpWWiOTyDJ0M4Y/p/wlq95gunIHnp1oflFwTL0Xo
IHFb8CoEu6fzCkSeVdz8+r81Ze6gb0xFApMvjQHfOOYZC9jCYQ57ujWMQUJOogJI
Sw/ljP8vG3SNtDanRqCxYa8ttNjn8xt81KHb9f0+zp1wb041tEjGRBQkePVtXnsj
eodA4BvEy3LLHjXVHX+4WN89H7v/jaEt4zOI3F94xVnkeuz2o2TmBJDemGUwqZyF
t35hZT/cwhJmrufRHbsoajUBuImOUUMJUQtDr4xqLSJgN21bHpKR8Sxq/yzO75zY
6vWFAbNIxxbna4kHf+yj9A==
`protect END_PROTECTED
