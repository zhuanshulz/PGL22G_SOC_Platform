`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eeQhnZI7yzVRTWhijs+9PairLgSg0Z8bnm9LZHs7owlmbTiDUqZga7mK03UgDsLj
WyU+S0ZI7hnm2gVSVm7pGdbyL6QJLtJfz6k4LgRfH43euPT64PVYA755gX4xbNF/
GkmE9z4gfncfHXrWRsawPRGgMAGeUoovzXoSgiLYsfV+Ni6SEzLBOpECOmJXbCBd
Su6+XBh8aUL7woQ4Dkn1Bp3GhIamnVocBEh4LBh9OAny6NnL/D7EyMLHbPxgE8WJ
3JgNLbfXkVe71g6WymRAJOgpOAUvjcb/TMA2z8Uo5PJ7J+2Xmihlrac/dsNdXq6P
ofP0/fbxpaCUS1/V0/zmpKIE+HuZJ23Haz2x3roGvZqfHTTC6xw6WsGWIUpSRGRT
wobKB8UNydthtTafamh2awicjXzviODjGY2F094d4//xSY79imHXR8Jdd2WihKIS
LbvU+29mn5OVo3KcwqUukG5wZvGe8QSM6/us7M+Qc4aPUahtTl1k4WCILm3K1yAE
FFYHJJtxLyOR4phCMxJkRwXwwOUWw0ujHvKXG7Bt6YA3HtaZ6Kto1k6T3FdP2Cx2
sBnEj+lmnJQwLxaTPDSO86Kyp+lWxHUd0ev2ngxz2cs1nw9eJrDI+uue2mJa3AHf
0BJ5mgCk6ekSj+jBFZVyh1MFUzI9EJNHjTrtPyukHdVr5k7nl9SZXbxnPdKiztXx
AYlJO+YsdXwcaks2Hk3KADLIUZe0ReNNqAER71Xa/AtVkxzKHTsi0HHAH45j9Vwq
IPKrd0WL5cdR7epfWD/ROtEcVQ/V3QQpBzzFFFVEp2Cn9U4ITu2AOEnndtZK7SaR
lS2CbxVOiIA5n8W2CFAV2F5uBIrT4t4ZAQANWTsdoLeFLNpxmXLbcjTzsio4Sgnp
UrvuEjOiSwXdLxZsQPDOjEWl2wtUei1Uud6N1yjxKj4cFFIP/DdeYL5awjOjS6D6
HTmwwOcbMqyvJj0hGmMrFDXGbrKkBoHLZ1UmibvvjotNbQV85XK0BQGoWTzQFwei
QcrhG67iVQJnpTs13tM8N4pIyQhfpwrvyep4Owhc7KA=
`protect END_PROTECTED
