`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i41JC8a42b3KkXUgxa1fWKRNZP+CB33TQ9V9ijUwxGk5QCu9y1w1FvE+oyhxmqOq
BXws0j9dvPgqGYmcPK2rzzuoloW4Q9TrtWC+eUr9Alzstv1pm/ey4Ujt5DpfJLYl
OtviWBolSfa6HmqO8tPEhq/ILxtkOtqug+1Zg4878qPLovZvfpsoO1D2zQyWKXIW
oKIPIU3hUn/exGmUgOLaGJKXX3Hw1l2lyIMxuNvjHSdyhHfB9t/0ylsd9o3VgEFU
QMpZwL5bHw41GrId5B9i1IWg1H/5srBVJY750jMUJDZJKXXorzyFZnfgzPxphUak
vLwAEsgH3F9XVO5N/1OFS+9sCDWxH6MDijNdPv4gJTFRd7/MTEqwBJ2OCdb3mJh8
hEijjkrQa5Iy2d25Mh3dxY8bubg0FCGXDCRZ1gVA+ZSaDi3qGqix/ljJFcZ/nAb6
YlTfFiARX15mQm4TvBPak9YOflzRQIosPAFaB8aGaKZImqLC++T9fVrsMbwQBu0R
X5UbqLmDSspNupL46qBp/r0YT0iNTpxkTpMxgXQikhwWrfUYIZAKK6WLxAToLFgQ
7AuQHP88y1RI8OXRbXMVRygLKT2RrZ1DLyaE9iZaiVH7q404HHqp0uiwED5Q74b+
B57vdvFYnwWnDlwRLybc0DySTNl5K2S1l8saRFRhNxapEtjaauCcB7gsgygp9CE2
`protect END_PROTECTED
