`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JSGxMW2NBBEaysWMRqB6dTvzH3DJIgcloiG/5dcU89y3tPjHPmGI2DjehC7aDrkT
o5/IicYrAYxa49+u90SYSRmdXJdNA8bPgSrZCxrKp3H7i8cavDDDP9jDuS2ZH+Pc
chm9pqj6Vd/U4TtlTZz9pjJZnYyPHjQxU3u62exRcnhvffqwHl5prjhoPamRsnSa
KZkY8zahGq1uf05wPeEd2HIBR2fIoJArQIUd0TXsaV9AKXca0g7+BeIoMj+Og6SJ
f7Imk9p9MQZSkPVhwoWNAn+UV3OzSla3h/UpmQ47SgaJd7YXpG90O3xpOPZmOIl6
VrTQtpFkFU9xq4KU9Ll4P037yZQ4Mf5kMZyO4lHAR625ieFlQDn+9RJGp2q8QqSW
ErlllMOiTYKMjS/tPsrJmUBROC7PjK8zzeqVqDaPx01jcmzmUtEzJ+xX7uDKdrOD
nZdem5rwszMMr/jeClvciJcQENraMKNaM1oRwSk+VYIpg5ejr6CtCfNFIyGj26uW
BwZAdtmvrKlQgh351AtuwWsGiVq31i2Xyj7Cc7RUt2p7MBKCAcEYlueiaUzHjYhY
WLqnqVWRkar9On9zgO99knCaC+7biWRqsazLDuqB7shCPnTEwBds3xOR8n5ENfGw
OIrBUOgraJpfxRvqQKjWHyhSfI4IDf5TFltjT0a7Nv+N+LG5Eq4zWGP7WMn1fyx5
B+3p2YTKlbPMFjgUZrRN3rPLpAlscczZVoBgsDyUhJQXpNnhyOP9sBioIsB29I9Q
J9ExlzZabhIwueyA5hucZbJCd8dxTA2mmj+oDMrkPeN4OSenRe1g1pFVrdHoir1d
RfllowxaFsBYLnku7UnSptlxYzDN0sOkC4IVRpMqZJ1s3W0BMZjcAALBv3FTi+FW
bt1I9nP/e7wit0NPTYgeJZYqDEC1F+0zgfWqlLoT/J0=
`protect END_PROTECTED
