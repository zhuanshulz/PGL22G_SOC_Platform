`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XFQDLv/hcN/680lqSWeL/6vrkMg6it6cPQXvl7fSZrnILiKDtJI3eHXClbFSI+dn
cIG8zBwIdFgmbgKW3+GAMlRzGh4rMwaBbGR4j5iEB2ldokZb6cdZyERjZTwtWaFl
V94+eTaDeKKV0rVmbQtppGIk3rTkAAJps63uW2EJGUHJFv4crgjoTKRIx0zOSniK
oaUPxPrOWazBI4j+ngl8znTDf6Q5s61LeWAUffHjgN6G0vmR8T8jvJUJn/r9K3rW
U/RtH672wg7eHL6XE/j5uXdpE0h21WJEFlqbdWuijNu2mC1epCM1/FfUVUO8A9Gr
P8KnZeRHLbPTCRmiu88ZfMOi3otPHLSJLwwImJRwqhRvUGPPzoUhJQ7Uebh27XK8
M6b+zDEAx8eN2Py4TJb4m4ijy6jUH2/zfdMxrZlycbh3rJDPnc9xDPhIdLhJg7eb
sLjUsRfj72B5TD0zITw/GU7FEMWPw9VtnawEvSoAkFmluLp3bP8lV2gScErHyYuJ
Y0QbNV9H9VLl0eimqFYFHwCtWFLs0v6Reru/0B6CsV+O/DctvAmxtHSWRWCgbweC
5saWABtB+r8niCkWH4UdWDQpjTwExBNk3Oouz9XUC1vbIRj7cn18IoR1iYXr7Tu9
u7SwQ4g9DyF1S2wb3FnRGrGUEtWwMKFpaavf4JOJlHlDp+VMQDdlu7wG6s1x+KmJ
Ro3NL+hoXz+dguf1YSZZ+Lny2YrBXPTkuRe1WdGBaUs4Ztlz/lcGp1fpBnWuW1f4
U449v2Cf6kZR7sbEBHw3oHuhH4iyqX72bZftu4HbHsr5B6fZA2gerg56ThQZVHc3
YfBkbw2CTQQDC7aVinv9cbT80friQf0CcdDlEhcJ0UQnyIS+6wIOv1YzFwtTmgKo
7zjTThSLnAAuMvhAcCuo38jjxnUk7V+O70cR/xDFF74hATf9tNY/DFu9icIX5ebq
lew4NxR3xqEDtvgoZy3KkwwwNZ30n5u2siGkoZNB+1gptsYmP3PyjIPNChbzthua
4EWlPhp87iKTixvtRIoJCesFZdPRTwyD7MnL9tAeygUZRRJeANF5jtVFFuGIIxlD
n+sTwQYydeuGtY169nz8uokkzdRK9lhoeLJHIJsYrRUyVsY7DWCwZdhzjr7/DtdD
Q0ojXNPi0HzOHzVAaqfTyodNaK+3yhr4P9CwG1Kfru3WfLC/TFpkn0XYWeMDIjBu
52h7ECmKhqD/HL50w+NCBqjV8T2Ka04jRlkIeSG2lxPdnDjhRvo+z7+jAM3pTn5J
8rij1hLl0zT5e6jU4qblfMoz3zGk4TIlEreJPTJajToZ8tGINLYCZi9C06k3qXg4
f4qzUcEV1bNJtNHy0ZjlpyLtfnWB7oSHckRvd3My5js472Sd8yAsFE51yNhFrCt0
r2qRozEAPzz4Mat14yyR4OiRBK3tOdEZwfUtoodon7w8t4aQD2Q/8uLJarCBE5t0
CRH9X6FgKMp+Phw2hgz/M/3cCNMo8YtO44FepcPoS592SmurU7a+G4ltmPoxwium
HVjyBE7nDWxjNsR+Qn0eo8/o9GvfR/YqEFreLR9LFUfOBYxVKZZQtO8ZWSo7B8v8
mYOgvJh37GG0YyIfc1w9GM/n9GaQE90T6XleyREU1zA1oXL1e7u+HTfXUBl3Ngd0
QslRSz5Tj5GVgPOsQkzjG3dT0DKwe8ANI02QlMKtMVkHyn/FVXKRjX7xKx+JjX2U
nLnB/Ygw3zeBR0i/JcSulGV5f6ge5iyXlG+E1HuI5FD2+OekDGlauk8c3uP0j4tT
5A+b91nB2vpoMp0ClqJ9F4A7zEPv1CtqAedUpyTbRdYqdTp6ATbttVhwRJKTnLDs
+vRNUD3D0gp12DbB8+lYs25Ylz2m8jN6VrqYGx7jXmMfFmTC2T5130BlZxNL/HgI
+Crxdjrv1n1UbVIuebfBOg==
`protect END_PROTECTED
