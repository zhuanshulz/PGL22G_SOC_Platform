`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f6NKdjEZYaCImOUg04jYaYUiHsPd6aJ6MtGFsRfi77oYD4acqjvRxLZEXNZGacA3
xZg9AmFXMuSvVVyn5Hk0ssRnenzeeltDeQ1UGs55irnF48zvO/PJLI/A82IVeOxg
e/10bINEWl4QH0JfH+lwXKl/Rm4ML9NIE93SJluDD0XqkB3FMzJwmYRg4fOMlU+q
6EqqIz5H69ghyN2g8bHnqPNpvB9ZEwt2MEqR6TpRmNk6ZfprUUZ5dDvTbm5FwOaW
y92iCZiVcrgW69UobCROErdsyzYmhz3Sp4b2+QOA8PbY7jLMUiB7MXQ8ZIDuLk07
p+oYzIuWlt46shFIgAfildVDRM8ex2XQko+StvozgT6txcNEf4k7Rc4YPg8FDYek
6K7qD0D45EudKuldPX5Qcbsg27LYJHCVJ7PeavRsOlgWKOYZWFa9Nfw6GciNXHKw
2966DspRsVvBezazGqEztfm4bXSEtcvLyQZ9lolg0EowfOXej5qGVhi789Ii/YAO
AUDBL1pGOdOYDidmzfrv7ELa2bBn9PJ0QN9JIeKgRHZqpoCKwUaBgKk/KMpnY/jJ
zD6nZP3XwsKdU8nNX1fkaB9iKAa5U/69z9uxkSCMhyAwpkmpPPdCv1f8pSQLb2OA
HNyy8Bu6fFzHla4EmT27e3Vn89ZvznkdW89Z+4RPosiF7zReZ+IzzyI0LIg15U8o
C9w95vhOQCQfB2KAWSGj5CWpm1iW6TF/fini6s89FiZA3JeSfyks5RDIsbb/JJAT
6ju1jg4x4LINCY/g/LIQsO6Co8DTM4NKTH2jz/5/7NOUyW4iWkuBmDaj/W3fmmTC
BtJooV9oLh7p2w0o2A1pHWBoQImwkacKChK3+MoendpssylN123P/OU1NnTQ1XD4
jGSbsyil4F166z5nPw+LLJ8I2PT5AoqXsZ/pI99MEKsMHOAnsvcsNEoUQPF7bdff
OkGq0KBjMF1AbZLDe5504vzFp4RvoAA6k/LzJOYU/kNEYOUNiGlIBfCHMbGEgg9b
d30q9Vnxml1Ftq1EAxleXsFI421xJhhsHWQ4tP2aOsI47R4C4e9y52Ce5rM5L/cd
ePnc1UDxFFpIzUKUR7GJcXNLqLaTkFJ7UreZv4UN/bWd3X0Ydkni8AGQjIjn64F7
`protect END_PROTECTED
