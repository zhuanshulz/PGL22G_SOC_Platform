`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Pg8s1Ene26oP5aT+1GPzP72fRpDjzEOFKDXpRpnHANY0Z4Ab1N7S6qD2E2nB9G7R
DGacWeEZ1Ws+kR/aX4Bar2adiuMVJ12tQEW1yjTjrsJdUbL+SePRqQUnPPVvfbDC
kjJQBMm2+aZISKdQCHV21mGyR7O7RIXV8DkgyV/g1Zd/8tKHqbGGrdJ01A3Cu52X
cb/BDG6l1Ez2t2y4S/Uj56RQS31nOqmvFRX+slbXbbiSz2hlzY51xLdpOSEhBXHX
pA09wlUU0G/MgGInPhHFTsiYvdHkXXRGFPNt8PnZIHfGKD094NeGFP4km87f1O6f
JjNs5uS2GDrlUFzeWeGMV2ecIp7Wp9oavz0/Wz8CrAAv9bxBTUjfKBefbrXCS5ac
/E03OxuP/03DU4yaF0z6Ui3NE4yC5xucW2uK2GMWOGCvBt/NL7L+d0RKucTivjDh
RoVOjGeaPQeIZeNPCNAheqDO0+1CP+0jMWy2GLsZC/8JF8TLMC9VBMOsNd1l6Res
D6DwI+Heb3ETUlGUUd3P2VhxLsNQx2uAVf26qdS1fl0BMaaihJDxZJyckF4FWxi7
thKcU5MlqyiU1TzjoaQ5Ro5LeuYanr5kKD6j8I8P10j9iZ+4rWpuIaeiqTMLItkv
m7MHtHL+tsgTo1q4wk9JqROzB4GTfX2YYvdc64WrBVrbjXUEk+yn0KA6uzDybXMI
IwI5FKMlqalfyTcnQHWVuD7zFtAweGnvw9O1JcViFab/LMayk3YiuJ2KExVuNBO/
s2FR2VJQFbDcUciXKwm3erIgmXiDiUppV9cSVcOdZ3XP7/YT0QxnG+qRc6bTniv9
pPShAaa/4C5+4H3FHmLD5lcAsPqdFIJ8O8OjBbgR/uwAHvdlaF21+mCXq2vEgONS
L94mFvwd5WbzNZcYoSgMVw5nMJlztJyvSKz3Mw4JSv0uVxVdBAJOzMhGdpLkHWBy
bEuuR9/1RtjU1WlTtL6Ei1PcQP69IHFX+5k6Nj/WDU4k/s+iLGujT55+kbN1XEe6
D+dgF1gLePblmRmgbcZ+vMuj2zlNRKpwpVsYYWOJxK33fyzmEdM3JW3uIJUniXTS
3J/yQzVqPK2xpUfe3joMqoTzQcnvb0+yqFl49DkyVLO9/M6Be+wvH0QiFP9Zfwwm
3a8/WIswq8u+Zf19n03HcfnXI0fH/sLtkxOgLgG+F6TN/3Iie46QjsURAUupSQga
af8o6ehOBzSG4j7GKFu6wtAPGEysAYJ0+2RZxDZsLcVKWzmwD0g4GW81Y8Hg1gOg
l3lkgIchsdWeCzR9vYPpdtLWhjxJKSw+Kzmd79QHvsBu1NG01qBOBWK79zSZOIE1
PVxm1478qf99utuXo7/ejP8w+R8Are6FguWKLpxQYX/+H+2eFZ4ybmJ4eaMS6Tw2
PjV7WYX/o84g+aW/y52T/gNC3nncd59+icL6r/ZncBTOeCWgO9hNtMb7odWYcuzu
c2e4upvDO5yboayAf4TgtSiIRLRep+8nyW6iWUBceywbSAIVF2/F+w4xMjxUuGqp
S0SdWxuJpEBnpwhuBaHov+5YwrWjEct+vvKhpM6nO4Fgq74UFd4zwzsX+cbZHl/2
/JmzgFXg/4BtkryI7fa5oOycG/Pa0gYXOrbJKrLJ7W4pWiPhG+JbGMzOzuR8bGdd
B6QzbiE0molgMv/AoasiJR9E50JVHaKUTG/9+nYNbH29UpBll6zOHFksnMsZIBtH
16821qrCZD+TnouzZ8c42PA/pFmSJyo066Rbd+x2qNCuQadbb2wIWL4eiw1O+kwW
TorGZKgtvnJjK/W7atR5WroXgcetIBu6yQYWkTT7Pv7oabPnl4tfvVng564PTnCE
mNAfeMUmqSfXWQc0tgukX727iYoKte+dkehIMvsc/O0l3gt66v6ddPmiZgItsv16
k2fR00KMmrAra5nV49hrYw7xaE1/AtUz422jxoPesTYCJyHSR4j7hSLSKhQex6vi
Dd9KBI6jwhvOyTFwMPzx4qbOrcloGqlvmNB6CFBXb88O88SAu6KF7GCbewe8Dphe
7cdZy/dFXpDMssT9bt8yn6JwKnJS7DKljZoEK6Tzbl1wQq6uWxyC6cIZ09QJ/81H
hdr7+nkOrDlkBGN0Bjgji+3WU6CoddeQAbORHiNiywB2BdqGlzBAcZ4IFsFlQ8Fg
dv8jbr3oVMW7WNZjIovWzONxlRHFfXqfYp12HyhcfcGOwdyjXJTU8rVxugFxwsI5
Yd5onYMFfxIVZhthQWPVLA==
`protect END_PROTECTED
