`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nCBqAFu7iH4CJ4UyCeCzUGaZDL6k03gAvoQx0qiusKV1gq3jqKZLwNwynfp4bOTT
IkjAtLIG+1lbLeIf966mhaaRuvz+OheHQlkK/Yl/+JMSrySXhT4/611IppAdwhuR
fNtKA9KfXpMglH7d5jvCFyJcev2DXoX4GMcSArqZmm2lp+OSndUUg27Ga9wdrS//
+TfKjgkCZDX4rJ7poXwCnB58jq4LkvO+9xqhaFq3k/8Ln5e2AztWSZ6bOWAZmOG5
JkrTADtNe++jw8uOcwODcGQZv3awfnZ28G7mr4036gOTK1ENmG5LX4BOaqsSARhZ
SxOezFzLshcQFN3Q0HTl5qGrbDcZH1YGx14dX6xu6rIw+DlU4sclKU3xCgoRaf3K
LBG+XS3l/5Ppp9QcotDjfcPaH+uEa/sHy9RovU581Ll9yTTU4t0j60BfpQ5EOqkD
xg9NqNKxZjxFe4MDW4vsCF4yH5ypnvLW7QwT0yiB/Rzg2uainMsUgd8Nx4L4Z9sL
VbgN60gjNOvjcy1xPSBe91uQS+1mrmRsVvmAXhLDgHqtwqewmM9tVPRRJYkCoMlW
qSgzKl4ZSTXKMhKDyEvytyjHWdEbGT57Do5A8L3IRMTXY89vQe3AJzWZBVsaqNDy
xLZJIy48TlO5BN/scc7/eRAbQC3O1tpyN08Kk6sYOSAtPX27v/Sb2JeRM29XKOBm
x327H5KHy2G5vhEYjMgnUA5P02iOYg3vOPQ3J4fiS6psSDNihYbhEZk1iugEpJ0I
y1YRvLNgDZ+lou3gvdtLUA5UvB5wZLpHvJptoiYUen1xjo+A3wHWa9xFeF+Mvq4r
8YxcC6hqS1KplSn45TjKltH8clQYeJKptSvJPeD1Mt3TD/bVuDZVin6W2ocCHIel
XPz/0rT8GZwsm4oncBt3N0ZqNBwEWtY5JyR5thTj4Ftl64OEfq0lcq6NAG5tJtjM
aYMu0K7L2FNxtBM49Ul0EeACYTrMvQS/WYMZ65YW/Bd2M0NgFJADyUSjNzjtzQhd
4aSaZLjgSSpxI4juXt48q3KBPPkFPq06yz79EyisnvO42ZtMgPkoMvseUM+JuvDZ
RrdxaXiieXBToqwKDbmuhkttfFm71ET9RDAoKeSyHmcnE3mYB0OCwcgT/GAVJjMX
/QvKk/247rUh2bHhwinaf81262s6KBU8otII3EgM232LyUyCUOcXjrIUhTcllx/f
4IniUHZUuiCQzoTqIkbyBPmzXbnMoTeZyIHuV41q1a3/hPd/nYNacVdaU4zpXwX+
pFx91pU1QikbU45nnUs0SbqP7Dr63tDtjNtWQO3rSpy8+ZyyAf+dYnPZ2kAZgCfQ
2E7p0drTLOt5DAAypZEl54zkZltchuFNDM9Uval7+ZMyrMpG0uXSrmwFYiweiaRA
wlniHolLTLrm2xcfkyWFcRvcGPfHVMnrbaSYTk85oW1AMPuiKxv4smDDW6oKjZD9
HjgjM21kHQGGXZ/fA/RQBbmXjb1Ms4elqgL08KZrw2v4L0iu+CqkzLugaLRqeIMH
C2h+36DFGhvlIsYWMe5BeabSzRib/z0m2RmaN8LDxhKYO/lQO2BSEfsp+f3Of40x
le3gRW7aqOXNuro8rDTzPF5yquZySGSysy8N+fF67UC0ZsSJ9EbUtJG6/Ir3JyiI
tDoBfoRiWTLaWAnklX4WGWNdbTVv07eRQUhFEcycDpBwi7vY3gqcYlhSBrslfbv2
b1iQ6PNRMTjJl4gpvgsGIzSnGdUFSw3j3tb3rK7uc7Wjg/8rZQo8F83Lmhz8shcH
GWowtn+m/YrfOiTBwqlA4d+DPVVYw5u8rXsDxTs4CAzkvUkG2PQDCytebYbpHrqu
bmmcCHRkqYmh8+KllwFTOf955C6+ZgUe0NuKxXxkWQJcVYh+N9p/Ije5HRiN3xH4
raVE2zsl8IPvmyZ8i90Bf+DlS915AKupybHF2ArC2Bb/fiLEEE114e8RcAopyZ2r
pI6LMAqAJyfMlrS4MKXOpu+04AkxaorBNAAv24ufVALHYylwchZEw21J7srlx7z9
gg3gwQXllE/WFj0caioLfAXFceYxbs0GOTqSEUHGgaDZiYMvChzL6OJIUki3EAN7
lpg3TMZl7cdszLQtv6/Sv5SQ9jjb/TVCXWN6aGhBSO3rtM6Js0ZSGgT3A+AwI8yX
h8Q6iHG/5sKR4G0nS3mnWyK8Ew6wLDc9XdNoeOkndP10xLj8ASDAniCqFgsz1MeI
ZmK9saRP1/w5e6kjDTYWxa2zVwAliGUS1A9e/SUt2NDLV+ERUVCNsggQqqKdDk8D
uFdlr6BZleXFa9x56mdbkc/FpHbcJ5vLCRFedKqITvGERMawDrDM1FJ+2vxZ/0mb
16JSMMAcmsgKpS8H4drM1zyf+2e0rdrhVzW/mSs0B/Jf9rME/zoszWfR8jIRoWEG
1kNxTI9iVEkN2gcv8MwL6z3tuLG/Q40w8DgdarSZWYQ29z5/MokqNxYOjs5CNpaw
uJuU3wu4i/7z509mC1c9ep8WnnzUi5m/+hKbZTyLwUsB5Sxa7WINEXLbciCsIkNS
nTEcTwaAKgJ5t3nIl/KbExA2giX65AJUAYRbfbov9XafSE5xMPxCbBvJhvRAdqRq
vJndryvbh2LNbK1bUfYaWv6X0sg5ph65OsY4VN2CQvSF5J7rIpF0alZDExYev4MU
HiNteJWTAW2vUz2BN4xQ6cDhAkbZSLyhJx1LYHk2ODjZrcWoLLvjBCou9RIY0T9g
PwH2VGruJc+7IqjtNYc4IU4KrjBY+w/bjGo3xRapRAhMxhZBJXqI4VuSC7jom+Nb
ScP+L+VlJSl6bXnlDXbeiXUXqEofEwoGU11ApZpmJvUfC2LQl10mRNRhdD70u0aT
BoFxhlgXDPmkABQesSoedhlUWkaM4lpYLkSqTN5endmlFAsWHypb3XJZV/vlefn6
M7SsaCml8IuI9WhKkL4Pub7nkZlFrTKBpunhiqUArQ2D37WVccZRwOB+XS2pHhtA
swTU2D9C0/4t5ns4x5BJOGOlV2hYiK7jNRWAwWisbQLFQTwVs0esjhbC0bsIN3i9
0dM8VztdigWHcRJqSBSpmZH/tYVOnYDC9B5gXsx9vqo/tHWTsMU2xztBsJmWQnfv
gnUxYYg+Kju6OQUJEYfxWY1wGof19sWIF6Ivs3EPTEciFhNQx5o4VLbDUKI0Rdlq
hiIqSt/Q3Pa1rBICrayCJpr0xJRvyk98bG2qz3SKe7kZzSAlwqkfEak+sGwoTFqA
5vHYm85Q0FLE3vmSuMiYcvvOD9egB6Tw1uejCtkIQsv/xbNyEjLQ+TJaZfgjWobL
cW/7NR5TqxB0qgXJL/JtiViHVUu0c9dhyCv1cHxtIPUYRLgDYpx5+Lpi0yxAHmBL
HwDQESawPbVU2Ov0+tu0iaxx7YKKYg4RjuUzWLzoSXOJqx6Tb+N+L03zU8SCdvzh
NBuJX17owdQSoX1y2dYmKcXULSM5uN4Z0L5BHLXWuCTX68mL7ZIEgpzIpWH4GrbQ
d5wiErEsnMsS2P+iwgLYwCq1hDKWLfmZKZJ1G30dIGh3upQxvXzV5L72MlUX7TH+
gqX2OYCAjYR0eXQAhvWzK5bSS4FNdmONktkmD/QH3AaNOU5H0FfvGBHdVSQM8ZBY
6FLvPKj8uz/Iz7V+GnGxFjxWP/nZ6P5zniSIEBYmSlyFCP+HUbIlggOcksSk4wHC
nk6zmrvQVgMxWqBHiCRT61zXW1selIkLKh4H/YUTEW05QV+npI51tqLII/cHtDlb
MG/CNiJoUifj7ovto22Ul5az6tWOHWDT+Rw2PAwr5iYrbB3RJK3+zLTFq4m1w09q
DHcvPpZIC2PC+SOqQzaS1aRf3YCV56PBRNG+Wf6YLYZXikSDcvuXclQ+3Ce26upp
M6CtD2sRYDJcFfHHrjcixljtLh/lSyoe8yz/hk5ntlsdPBefw2pNFB7XdZdhqUCp
zdwDfcG6N5zIYNBvkCQck9Qk1LgOWHr0ghldrFFJmJ1RpFtS3yQb+1khxmWtMByM
duJJWUqupwaulLSb9U3+BT13s319IVEHBhBh0o2OIfzNujmtiBl6j1st0WHPggLi
KcB5QvEEN1SE3uNdxsSBqCtmZv1wZkeZ7wmftpUYBbn2eIwTKVu+TzaXnFU0KtXl
O/hrNtsbtoRu54GroyaEQUCVv9wTlLRQNr6E2NvBy0Gqq0fZ1sEq8TmYNcgc3kGS
gmeufX+srGvIzihO3ykic1AMTN4e/m7w82jUMbtZqUsy1LzLZRFb/7fLgP5i9o8B
gvJ4uK94cuDukEPn/B52zIqkeIp44fpdkScnJwVy/faMlQqIlXlPToQvsEDosjBo
ithN2/BT/JhF0GCbCAYqw43vCKL79ynKduFSS5FnfZSAKvgPIeWQCdbzPTjDrXF6
0tRyrgleaGd2sDz9bZtRYZ2iHXMMvsHMNGSIuYGH284FGri2IiAVL8SybLkdS8Gx
ALv3Zi5vNtGnEvfuUyrEJSoPU5xcB9lf0zEvt2ydNkeZ9CJ4uA4hoIAagnGFIsax
rvzB9odFxi7NBoBcAdxXe1TQQQvsLTk6a08rqUT9sF9N2f3r03MKIW5b45BvbEXl
zyoaOS727f3U/lu4rP9i130F2J7OcxETNF60+6DR+sl2jdr2ZwnNvagkDMltMogG
KAE4OI4wyECjjid2p/2gg1JdZtUzak4hVMy1ziTsRkMJx9e9KgVInAtfWMF3j2rK
DPCfcQBdo1RfUHU4u4aJuvNzKOnsa8lQqnT9OxGeK/d4xr0Q5hMuEJSdzv01QuTg
T2gHCx9K/8cJmgfRcdwATaotDhbM7ttMzZgCGDBYI3RqscaKRFdM7A0uoIr/7TCa
kxWbJtPg/g2ewtjLZbfQrQXdH3fazLhnqLdK5oBYp8etsao1hbzxBw+50/NmXW0E
QiZgYPdF5N6dy4WufXAtee5KQVcsTk8jVgaH3ngySLMFPHHQbD3CAvm7sm1X8D9s
J39/w17MIp9Ug2+93XgzokEWh5UubsOog9AIY2kjIg/uPK0AX47hygqwVg07Ca0d
DQZxhU1IYxh593o4WfhUaI+0tM95rclUTu/DUq+qj5TdpBtbSuKl1jI9Ps081Xrx
7RgIPVDsWkHn849205h0rknihjbofof1lic0EfDuawP3cAmgSod8G89gG7HAWfnm
PEe5rzbl+u4R9BnakW9udTqh7LUBqAJEr63T3+w6WvgsyLimwcP73exRzD5mW2aK
4ORUiajJGo3ZKirieATMevcjIb4o7tLbmrZaQReF/BMnI3hm0GU2ZtlF3mAleT7v
sxiPHEQQzdgN5ESqk2pB+ZMjjyQ37jRjBPNx4DyF+Vn3QXsxuN/kf3VSuyutizho
bCZGH+V5dMWKexeHV+cf+vxi0OZ9HCavNchxQUHTcs5xT4EnzhFr/EWH6M3zNqda
YrUxaXA5tgOAKkK468pN5lDNAFmVvpZN+dOodIen4BOXr4/dTQto2fPrc8QBDQNd
MmJsJ3IDg3zmGOqil0Bk/4kUraqwpL9PJfYQJ2+sJysf/+EgnRsfRtqeeFRAaM8B
2y8h7YtC6JdwlMAET8foKkKbfHmXsjUD7C3fGhm+0Pr4UcjYj7C+oApk101SEFvt
RiG43P2jQ32OEDI8f92TcfenspQjFY3ZeoxyWmPX0oFZHfIuJs4VCgvn0AFIDIZY
tZ0nl6YsKprZAvAQM975IDYG8MnzIPebzz/l/wPyfP5qbaEtcXyYeTWsAllGaoZe
7b5gFRI/A/v68IHTMf9zlqxJuvnN31zZ+OxBEg3CihEsQzrFrpu2vFGpSgoqNcGm
PFpoQ5c8fJ2zvmPvoh40uzyz99SVC2SI0ihPlcH9f0956wcuqLgZHeTusZdni3Fl
7eJmVGtwX+iXWzK1fgfVxBmWcZ9K+JLKWI4rD+a00P7G8gyouVjdkyBmXHLHZUzH
12jlhPFpf/DwXHCZqka5copegeE46Tm1GwVZXvSDE4cGwcY3DJFGhbNPG/E7Zvoo
2SIAt2jhsiSsN+watQphRNtBnlDPsJW4A1dnaNlKvDOLNsIHfbJwDSU4Nt9bwxZl
1ZMsG4yH5x1vI5OXQXY/LxhuVqc1R8oYpCQyfAwxR+4b/78wdjS1BMBbonHCCd5y
vuj33+oSy1pkUFqPjawmBT7Ch7UiRoBst9pVWdoAkBXi48IXlS0WcvAoZSEpYanr
DuFyvMk5g0cOrPcqCRSty/DPmDlzO9nt3MXuDLZplEbzhz/dLYRp8+xN8CVuOFpa
2QNb+Fqs5HBJP4A5a2HKk9hzbx74NNpplWPFFaXY7fpCNmamQd7gX8N3VA57xRXX
6SEhGJnv3YWA6FFxHbIBUXGZ750k4QJk+fzxroZZ7PMGESG6i741B//1RZY6cEYg
iqPUBd3bvMHr5fDA85J18LTfGejy/EUG3De/HIUKaNwBSS+F3Oedqhni7c1wfamg
aR5fM2J/8qBDaYCi/aT2UbnwXtJAAupA/X03KsYKkKwmGsROAw4OUWnM57qNFoZj
1qiRzN7Iv+fpTQtHYX/QXvG8b+J+k0a+KUIxHzqcA1uLxDlCSh08dMWyDmHnW+M1
ubW+SMkbr1kAEXbeVfB6p0AO/Oa8wfOS5HBp5Ay6sX7bc4MZ69VI+ZC/hFgud5Bb
6NFDX+QSjMP15hdQAmiT8TSIXGWpxyv5hFyTIqsiRPqJV6JC2UeqD7rutOOnXIJO
L9GNom9VuwN5CDQZ7cN7jYGmzmOzWemHoOIEjosF5SNWj4MHphYtAlrjH++lohIq
kpbQUaUrLfDaynZnQdgvA+tktkQO7FM28oFuW2ag9XOEjv3nuEUGhx5wc+QkezVu
dYxYYbhBN5RspCvs3uvVOtLQH0sW/t+eVclNrr7LnPwihbQAmMBe+aQBjIw/awPZ
AzgPRo4rBJW+XYohdK3b4XpvsW1mgqF9BnYkuPpH0Iv7Gb1DdZldDHEg9gmo8S7k
7K6h8Swm3k4AokcPf0Tjaz5/8TnvCdPpg7ExOnHchvaP/X+ozK9ArbH0oVjwj/gY
rETh7mfERzF0IJn2+JQXK5Rzt7SpB2BRSORVSw5/RMBF6qz1KtfEHlN6MSLawob6
wo+uuoy38mk6uiIRsqhiyPc7tw0XdKRs3U1FXEbxRSzh1p+F546BxD8I/WjKYypV
IvZ5b56QT8beJl8fewi2Od4bkyqrqhgca3DJp6zaP89L8EAjDe85i8cLNgP3b4pN
Hkp3TACpyhwBRmcAGPEePJYnb5Z6mBL0vspX1UeTgPTuTC4TVXKFS2nWJmTSWcry
8nRLv+ByMGmMfI96v0BMvu5P8VLNiITYVRElzynjjacfPwFoTZlrnhEeQ6a2X4Io
h+ezq3qRbjS2loGM1XqyuHrmiXSgkbafJUnNhmbYe3zoXayhjy1LrKjOZowMghY7
hIk3FWu6ORmVjfXZKB5Lpah1aAdKw7mkqXtdX+EzVOTBn4K92KJeiE1Ek0ipjHsE
hdZ0sRhC76n3VJCMfzpWhoobl+TD8qPjQ2/HTgE/IfsTRAMRYnRNFp5sZCAeESHQ
GAq4TmFW84atoHnhKfOYh7PPUqiDJkBtfG+9KMyaeIcIZRTQdgOnP+0PCyA8PSsB
juZFEGRykEVkXyEK4mCpbyGR0immcH+lMu16DFdBgNM1AZXhZh5nPtpbgWLJMidH
rVC3Kcb9OP7eVGplPBMV7IYI1oDg6YLCAnfLPUAjLUZOZQwoHgw+TXDKNhdagbYH
YAxWVIlVNncj1ue4S/O6cDYuB6k3zEFiNDML65TB3pZIBtfufx9IU/s56mw8YlRL
5K6u7owgBI0PNWG4w18be0TuWFW/SDDsjiTJxkoBSUpFpHeKq5kCc+/EBw3CN2KZ
/0CIuaeHevsxAyMCL+wOAdZY634OXqPZShF0hY7pskK6Tig8HswxuvLZj7RIH7RW
HFh2PZ+e6lfWLB5XoBva2X9gmHFRhneLsCr6IQ3Akx89oDNH8XdWaIaEhb903bdx
65wzF3678BLoeY+LBhtnjfXLwf1um+JXjIW9NN8jcmA9mSvSyyqsXZ6WeH4AKlHB
uvrc6lfwtavKjly1rqF+IpPW9hRqeIDIeLDsLIFABAcYQaUEzdGbZ8Rl9A4PP1zP
Lri4GYo+WCEMwQAAkvsqBplvOOHFpS8LFL4QlNCAiSrGbJ9WF0RQ9nPMIF6JiM/C
fS7z6syg39EUdHyw3ikLh/JnQ5nVL/udvV5RVEI6I86t+pC0nyjeA2oN0iVTI8CY
UZpmdDK+xvShJLMG858d02Wf9dAw7qGpMM1AdRNHMAsRc6WmWgC8qEr6mAOuScDc
ejo+8NQVRlP0ceiFtH+OdMfTM/oN9m4yKoZSQQFmpoU0lVw8LRxTlNsNOcAlDW2m
HOZtiDNAHiGdCqhKA0+Rs7RMfmFiNV4jaeuM83vZRsCT7UbLm3aRWIz0pSix+Nni
j21YPbykEU+Cr+kWkdfNIy7KXR/LthXRdhEG75hEWHlf74umnMkye74m1wzx7kZr
AwYNMMjrkOT386zStZeC0CDjh3l/YDhHTeGGqHEO856xkRHSJZlz1uiAFjMUjOsB
/hsP3lqK8RqD0uroYSnQ0Pr/mQQpUm/B019T7ALh90L550GB0GMOOzry91WZV403
bqBFMKvmFVFnGAzvYea/nxrOefzpewjwlrEnG1cekg/iyiTuGZpZveJ1S9l8nKEe
NuZ9goiIBYtm/hAmCnI+Avp7rRdr9Evp0TzHDz7mumd9bg2zCYkUXyYRM0sSKKtG
7MOupGOQsY5N6uUicCCrbF0NBIt8nK2ekjzyfs5rF1+lFxtFv0mBFAVSdfMnyjZG
EPmTulW5XzElbQgLfM7/Uomb8nRbQbPEOc/Z+SF8GLrgKW+itGfF1CjF2+g3siN1
SPzxgqkp917+X5/2GnRo8TvQm1DWpInZXOKL0M/JnQBlW1ou1Y6++QPRg8n/HjS0
bn6AS1sfXTNjNjXRpjFABzygJZr/dXN/V19glQE/1XA9a4AYsKPh7vvEV5hfexD9
4T41SeaGX1T/t6ThrcYalzoj62Bncrnk/3wQwnmLSi2uGWuQvJWfASqdME2M3W/i
gPH4KUlCWfatYpvZkKm1+7ArqnUosaqTsPzbFTGiwgl0Qh05WBb9L7HkEBlcfsVL
MKHWSmhZxV2RpkGtEgi667F3akwQy+okVNpm6hArbh+d7zqFlb6j+bxQyfp/1/SW
SW0mL34SdMeWj509j6MDhFUg1CPi7IxC0VG+q6PeGS+hFGY4BA29YHBQxZF98UbY
z8WguhzqCGkvLfBe+FBRJ5ZBp72ESDpRrizzHoFNPA+X5zr7Wjk5qKlM4B2nPXxd
7a/fy30wypBup3OllllJrOBZLF7Hagx3ntknE4IP/c+IZnOYYRhKVlVMwS1OS/nI
KV3YZrUbtKn4nY46n0fdc0GHTMaVSGPBURxNcCayQD/d3Fz6XzgzYNoFPZAlnoar
2gMm6RgDiAZnB/fsWSZaP3zQYQbbomji5IbM9YFJEzxp8NRRo49ZRim3eV7DG5OH
Xqkf7CyBaJ6EsI/WYUCRaekuo3bTz574aLN803civ3DJLS1LPPIMSnwHab1ekev4
4S8Wg1bvCJxoyuKLGQpjsibQ1NsWUWmNuahtNbhUjkJyD+lQdrvdw0kxb53ymDV7
DOsR1d9zd+I4aL53zXugKeX2x6Ygfv8BH81fe9MfNsGjLlo3/J3rOapKtlJAKM8D
kUSRf2Rg82uGL7puRTkSBZdr53COMaJ3xKqlM9zIGMWC+lzSSoQhRUCAQKbe/5SJ
keTtOwd76x/SA6fEDhKifsj0RaCr+XD6+W7YLFVYbVNfWZAhUKhD4NKKO+/MHGYl
o9cCc35dVP8T33hvGWZRQMHXrW+IU07zZDCI24WhIbQqJ2N7YhoMCG8ft/DVk23B
mtH8GZyAmNeB8awApP/rlq7TNf579n116JjvD6cTrxrOZLio8qixO3Q/8jX9xN+Y
iAehVxjg9WI8Pi/mLYEIBES4Wlw+a3Bl/2q4ZMc1W2/EBmp3jtDHXeF4anfPMCOX
7wT0ySq3eYJLolDsBMy6nYlEchNehQpxjhyy3tgmor7mkuZzUB5H+uitH7558mVZ
s/tlLAWmyRBj0Eujsnetu3brZ4kMqy+McnzctnhB5AKHALqy9y7/sftuIJToWgVn
Ib6g5zO8EgfvgxiOFyW2b9wOvz6HqcAUsC0ncAlwUOVZ09UFvUDTOtcbAOjpkfMp
QPBKYONqnrFLyLsjqGTTvVRfNJyJhDDcf4uKdtToleuN+3Vn4IRl+tGbesTdMBhP
8bqASTPHcfpty1YwDaQSeB4kJfwSTbCZ14VPEAkhAu9x5JGyKRydAsv2bQG5mgoT
I672z7b7cp40MrnMhsu3PpMG376AS31GlLo73JtmGS4qz46rtG24G8f4KHSWomX9
SjERf8Ycm2tlWDKNCvraaHFuU1FTL8Ad4WQL7P4Sk/CYjR5wYMLDCVmCF/+ZiCUE
ce8AaoV2QoGmkH8olK6fdZzd5OnpzCnRvPoZS/CH2x2pXRRwZD2WYAwKwSfN9VRA
wggYdUDEOQvngQpJxyUuwfEtLQ0sxBQrsEok+rthbvkEZ4VTyHzb2tC497N8gMfa
ihBkaN7LsA44tgY/yF5FdcZt0eh3k1pI8lQKdcHGSn7YPLzEu0cb8jbw2xicaQHC
XdDShJdl7AQHlawQgQDUGCP9CuK6ygXzcPEzgnE0VR7j5aIjVCq5SGMPSS1P/q4I
lSMMnuB4i1oPWm7lspx04QO5pgalLDqIcBmi7Hhl9graVD+H5k7SGhzMoKQ2k/Kk
ByBCuDURCEtHEuu7Wc/jA4eKfeQUzKLM0L5gYHQa0JL+XBWeGSNRjv7gtwh6LIqZ
kzrSZsu/XnytCFUVx66TAJZ4UzLbS856ATOOQA2L7/AHBkARvMyIZLMe/F9Mc8GZ
hLcGrduPEnDAP2v7rHTY/4Y5ZeOIAC1+hdXlU5mFGVT5czUY//SDB+ItMM7wzaWE
dDyxVifUVl2iTVpOKTYmBw5MFpAW/KZiZzjUptG4N3vQ+O8DaaiCtqL9LBOu0NkK
g0T8ebnV1hm9I/NKjgL+eBYk3VDC7frNOk8YRS8Ny60Jvr7aHsBwIREsTlYtbB5Y
9AHaXGTRGoucpy0111o3XnvsjFzvHy0p8BJ2N2JHm6HBwA0FM1LET8bujY7ow9g7
pZwY3szFVxHt+C3PaOOzBN+mg2i2hvX/q+L3sJyQs+alAmOZs6go3aL3p53/RU95
DlYsSoRQX9oTGIaOo4cgYBkIb5Q21xFS1zgcvFPhmIx7XTKwoas2VihGH2sWWyWn
TZhdpSYhH9AvnKBhRIBOkrZsAJIpa6MI+nUsCy6lXNaeqAwwFRH9QlqCvSrGdwXa
E7ZjogyXNIB3IG50T71I1ynbrCWi/Bq2I/X6vREMSusuVjhOg6KFwA2lDSbkAV69
v7f1JFi20aOfVf73yh4hdvuwTSQ6QAefhACIoIQEHX63mJIR3BhIuiW0MCsLC1SE
mOc+sZuY8RqGOGk3L2GyneOhPD8iPrvXUMOSB73KZd2BA6Ue32UUge5yj7YhyNET
vlzvQ0Po5AhuuZHVozEgckWpSAjz/gOFCzPAs+bbn+k22VT71HrpDrFuX/mu7QKJ
+Pzfp6BocxKJBLehuChMq8BFkzVeMIc7V1YcmI7LlY12Fxcbfp3npLotkHNila/e
mr00idGQmYaxbkq7LpHutKDbCB8/pWMYkXsrrU3Ca7NaQrYCNt8quc4xUtiJnn00
Zn1LI/lb7YYcP0CrVmXBn6J7MKc/3cZcePCDtGVo8y2NY1WX3N+PeRynftEKPhfZ
+aM3QOi/eo5pAvL7yrp1awYMohLXpnzFAaZNSlbQ4uPKTHp3sCuZBpBquPm8B9hU
WZ83Gc/wk46AL+AqGt91Nrqfb3AZOp8lZ/iCv0tbMDBBHwjWzJpsKGjY3SjDV+7d
F14ltsLta6TPj/GEQ5ylPvAdDXsCGbiAPYgSNuzWdyBmE5V2GIUp69tuk1Dzvh7Y
mCkiyyJWtI2HqsC/gQ0XDJv9SO+d5yIP4v2ANZoBwgmTK50kuq//sd9zzv9qGI6Z
bJZjZU0V4iA+wj/t2FByj+Xv3vYPxUHiaasvznP06Eiia597uedTfOuLCCyaazKW
Wevsfc5371u5URJYkA6cp7cUa+5fkZcDBE3NFR4Zxn7iJoSB77UXy2WswLiaA1Po
+t2aVcuf9JDpJ0lh4j0AxXaOAicBfdd1qyUPrIDv4eUIoPCpytioJPQbbri9h9VE
C/SdkZu3v9lm3c3jnTh6diYMcPIr3Mn+C+dNEElnwtFLlKhsjuRCmdsc5RRWwwNR
YKSPvdBQuXrZ59xVEMenwhFiMtuV7lT+urRJvYCNT5SzT2GAne80YU6TKq2Wgfxg
wtMx18xLrrEdJbS42MkW6UVv7/twO7xUtqWqhvXoc+IQPFRB+yhciWIkUAG1GGqo
GxK9KRE4btppZCsQx1UAUJYleOqgy6EWSnd3udwvMCZblFALMjohy82WOv4CWKJH
50MUIGy6ICyKytpzvi8C4Z52VT6NeUg0btNu7tdXnmIyH2Sz2eDn3auza0ha3yPr
cdVNC+ILJMSAbcFDKHaDoNmxRg2LSE0cT6/ibEFiRrMANNm4l6SP4vW6+wWhhREV
jDceO3bxcyTi6jeeUdvBB8NbvOhHXYTS4REfNILtRWQooolst5nhr/sfKlLvseEf
ht+kzRyV8HfB4beYY811/0uIWhPxgVyaWcL0skbJmLZ5x3T0m7Dl/bJAqN69Tluo
yUl3VG6D1DlIBD/sywK/een0qkVW3m8I8B8+aKYKql+wgiPZwzUAN6NKG19mnAjt
oi/UR4hjCJ2LxHscvgO5f649kV7+elKqFCV2gzQEe3uiQ7kwpv4KcryWcw5jc0qE
rQitO+wRmve0Bw4FqnuCYTqeHg4t3xh3CY3OGDHAN7ut3N1lnAvX2gBMY2OHmupP
TZVZOrF6ZaWsuyf/bDHYGNIM3G4vONRS29O48DHGygV8hzyNlEhOOFPP00+7rtZN
xlvVwrCg8D3ZkCXPwRqcOC5Ubqv8k8qb+n/fALChFWl5QD3RufKixFTzrkrlYtVI
jS6nE8YeXpHbHK2PJMQiuqxqlb7W13Ot8GOR/sivdMR7rMIEWGSHQWUfmXgTiLsg
wuS1RRd0UyZeud7MMiCxcYFG3kmqyCJgTC0VsJxQuXZEcTxJrbg6elNZLIgI8JH5
oteQOpkCAvMJIRx/ANnMtp+HlQT/BrNLdzL6UbaFAhZYneGXmnKgZfXfcljWmopJ
TZlUbxpDjNmsFOsLE+oSqthey7fUbnHqwpWo50dMlovA7Hv5WMg0H1ysIrw57YIh
CHjZTxypxVShxXATXDfWhttAbmAKvIIt89MYP4XFYZ4rnC7xtNJq+1OdYpD8YrLc
dBTzqxlJ6WpPTJzcUlhi8Y77ACo4WyK3GI6nn4JdS4Efez6+aPJCyyG7AcVQhk5z
CKFijvYS6PhiNhlhyr9wX/dxT7uIg9zpB4S/MFFrVjb1ke3M7YchAocpptq6b12X
kgAoWSuLa5qRI1aadfzqo8v0Jwb6BScI1rmZ9thjFCoLfbwOCWzn1x7yCO7fJIn9
zPgk7D2lvRXfNyRaxVCHbRz/+9TREwLRc4NyMIUDmDPRlkloymoGf2mWAWaF9cVc
AHNrCx6YczVBNL6DVLANeW8PbjuAYzxgpBE1op0AZJZipI/s7mP5bKN/lLqXXhxg
yQAlJ9MFqMx8pAhrdq6romPavLmWqBjgnDuaUrTw9TJsiOOKuU38+PsnnoiZhrn2
Kry3h/Jj5HANXAVFA9erdFJvlEwdVyt0P6dMZc7nhfY4HGsYpNmq8Od6zoPHUKR5
dfp3vWDYFQnvXZnaj7CsXA6tve+wKHiLUXq73sHLyh/WrhxXvhu5wNBIRGxP09vA
5BOpvZWsvVuXldfnx5VClQHCFZWe9ZR8FUQFrU7jcK6WbsQWU9Px+9amtZ92ZPux
ZBG9dGEy+oE1fgqRkpgfNwttNQYKYn3A9FmtQlfyIn7h8hW4dQX3peUPKhDU0qdw
NLVHdm2JFcBhlmiAmE/oZdQSAUwsxWRiKVTUnUGuY6LhSuaZb1jjW7nSUxmvTB0o
8YnXFYo4Qm5PXnl1lJ2/l5/V1FRv7EtrnFaBNUZXWVWiAmXTm6/JF75VN9MpgRYZ
8pYnn1LUiFuvElxmnz6ARAsAAaquAU+QQ3no2rZTT/QXBUZpXTa7AboyJ8g8bzP8
KoeUDmqT2aEkfVeacqe4IFDhkDBrSm3ZDVXqQ5kM8wjdz0IBBagYVt0rGO60ssig
oP3COm5Njp/D49Zwra72oIiRirAcHPGO9kQVfhB9nFOI8np4O88YXOTnYboJwi/J
GI3DFoXaltiBKX6dPC5NjUEn8fFbZtYFLPGl3D3owA7gFE7caW7Vu0bZcdYHR5zM
q5x0ChnD9HXV7cfN0NNrJCyonFjPTp+TOWpYSgC7irXLxDEOIszFVcWHJpZtfM52
tmX10iuxw1mox0JsFGOR9ZcIvixY8CIK1eF8vwlfp1JMxoydZ6JlksTrVcNLbpki
1+atGBKWIDjE4K3B4j//NbmV7ngmZAeouOZxn5b2ySu/f2TYxaFkv9myteksxToI
OOhvzq1qxRRA4fHKNEb/F+JjUuCNEzjIdhZW/4Y1R2HpZaBDM5/CA0SXymZBgr4W
vdz/fbgAe7TGv5pvgU+iCJyrSHbNhE+dWlqsVLcstTzWpWA7Je8MJho+0VM/5zFa
Xhza88u9u3o+19Y9ljolxxyS/1rRwB6SpJBcLRDdIFvTfOJOXKSkasZeYR6OHGMA
OQcjhkzLObHr9psTAatwlqdyZJeeryp9bwkTeS0mT8uryiTYmfRhb/T3PTNZe5JH
OloZvC23DoHoxPFZEDXYepwcBD/5bMmPsvUsnBBiBnvrDa2RwG1K3cgs8sTPakfT
8ETy5KWR3o4BjE9M+LrYtZIIfk6DyP0+7jrmBUFjyM5HoTNVZ8yWp4gUqXc2n1Fc
leb+R8AyOV3w41fX5G2Hqu3rU3u/nsqy3PUuzkE30eZvBflSyXDdKk1R/T9N1Q5D
OeGBTWsPtbF2mfEHhLxBCo/9J29enmrreLbO9fuA97nyC0RA6GgJdC0/Iwd329as
AknotcHHTFlL2x4+0kwPZzsFj7pa6bjp7I2LSrsWeqWqRTx/XoAWwBwgewAQI2mv
+zSv3mk8VBBj+iEDMUgPjZJNxWMQRxREOawMP8DN/GseDdNQ67Hu62BlMx/yqtIe
/Rc3GG8d2vd8xAwNYYKfx/24IxD/vz5HTl6tt777e6qfyNsoSaFMgO6P/JmcdYR7
KcllvoIStIVxymeLC7xXEysq9gcnIGeGAeycWI+H1YaE+EFYCsiEKgG8kecIO/Px
2k1Kx5UIuys/Fk3vmAO62zKqfy7JL8OBcULbJizOkp7/WUHJWXbvxJn2/GbekR6V
geYGpsZBPwlIsGhzN1iU4OKzYhvO2gz8RLNjUYOTYyucDThvpYN9yn0WByw7r7Th
Vug9hZdYjoezhhAvpHCYPY0oCXHN4LViStqbJJ67Y7nov1rKuNZuBJnFiw+Tso/S
AwYYSy28JDAPnRoQ+goPchjOQaALt+kihzPpTzsz/OBSmLQQhItzzDWECAig6G6e
yKM5JG/OAKeZeGlS2EK1MHvI40dB+aOjATAotrSOcHkJ4g+qRE2u1hHGY1J1QHBW
Y+SYN8w6GaaVNioKnD2BsR8E1El3YMhOf8gshOfMINoRowRUbxSMcUokBn+QCij5
t0C1HwpGFLoYUYlvg+4JOo2Sr8hNN9wVMXViNVMV0gb2Z2hJEIUxFLa6lWezx0U5
G0UohCdRsjp4kzbbMQfAXKpCiAVygZ0W5kQzC/QifuEf/oB0DgiR8htJzRmTf+pj
oyXq95tZdedsXdLsEYYHHXcxEC11gez2xfuQYubtMNst1rUYuSOA6V7XPVKOT7Iv
vJAekqWyAIL99ml/F52wGdPQpDcF6nxEKIiLktrdkYQACAxyGH9fOHL+KWxBmpGW
qJZKCnhOcxVJDWNjLYOlyrGcrOtZ52xq8zR50++yXSVhTrNKYzVBiTIEmQYnm7b4
onAyVGK3oej5xg9/2gyGF2aSQURKtTv+37QOi80t0B0RyhircMCLq5DtQWxyKexG
YKWAPIrUOEDMkhLaR/X5ucFwx/Zo+bvuJruMe3iJ5LG/SsTHkJdBlbN1bKVeJKa/
18cuU3os6QtW5XNHd5+BtJq2jwVDoiywqhAZ2gwJPH6TZ5sFQam5DZO/ZpddEGfs
9XLYwTXO1wpU/ogHwHHNna0mFA7188h0JGdIR6+8+byAi/qdwKeRrH9LD8SG++uz
DNVKvMXEXFDm5lCnRj+xFFzw2LtJVtQpOD7VTH3S5fVLbZwkkoH7yZFvKwRw5w2L
xH5Og0KSvTW6HMCvPDz9wXkl5TAPMbmUphwQ5WIPcw1mKft7t97xbJtsTmBafoIm
kqFpWZQr1LBh1Ldhhq0US5J62AANxFK9+Pn/3p9oOj3olAMjlhmyEsvh1ls8GnBA
dOx224FHg/q8hBwVp8WEv3c29eml0RuJScRU0SWi90oRgIIeQBC3cftmnwF9Wfgd
VXGqNLBdtwWS0SVF9Tw9Y+zqzF3Fy2MM38s4a2uSCczqvwiueuFWTHR1VxJsV3f+
IJRPHXlK+B+chBV4Li0FX4mHjkEZ7sUXHBvHbL0i4piCVE6e+u8TVDAhG6jt+dGx
2zKvPQhh200GLjd6Om1qtERzihMkQKU5Plo9VBekjuT/jEKjJ23dhR7r/1lS6Bes
OFfS9FKm0JmZWJCqQ7Bn+zsoFfljDWabytx5DcoS/SvQXmSRcz9VO1iCvxKIkxe6
gf/GK1h7P2BZM/gdlH7xjOga8Y+KwQSn+A9uTslJFylaAE/+ejQSCG+2KmfxOgCy
iuycC+H3Y3RqieaAPrmbTb+AfGSLJaCSBBkEjQZGvF0nj82Kp+M4/z7y7CqhUxWD
FBoMIeMw7CwgHOvedimxafKDNdhlSABatGoNGuLzuFndoKRjB1ajbbaIK8pcetdI
c2fCQjruVwWts16J/DPEnTEVvws1GUCIoO2fM322TLc81xdFapLwhUATROiOg7fW
Bg4gQGsYdV0dp8lEqutO25oppEMRQ9rBSL9HeMPi332pBXs3UFX7xg3/CiQNwtWx
+eRe0tezMdfvkH7mTEleD2HRECAAXq+CON1817bgqOmbAWdf9/DbEqNTPc1Bv70w
ruWTsbDgrqNKSRL63cBJhzQLZ+Bu6HFGWHucSWaxFJqO2SjtPfgV3B0Yk6EdX0i6
vxxpopMdRsXl7XvKbhEeZu2mhgZroBZqiiMWs1IhslR/ST+xHclH/M8rik7sIO0M
vGiL160F59aVnfQTAcfy5Tx/1CWSJKC22m6YIzPKIkgycOjYPNzQMo02466hUKmQ
0Fv47IlRdrPMhzkkJSvPI+UELQUsEvD/9stFh9hDP3ph+9wEKYrHd0Rcw9zr5Rwn
UO+knqFt9lxfLPmlYQPWQiEAkqtoJc9+1kiYhSL7HF3XZd9AkxWtozPaS1dw+sEB
amujB41z02AoUc+IuMs9i/4GL6GUa6WfWSAToDbiL1fEQUEwb5rn9wnAWIUXwgWN
M9qe2MhfcPEaYt3VB2UcgsuNXJKCvifkq0UyoXAgfrSe4tsr28UtdHsz4S6WK/5Q
CSEhtuRxRw2V3YvQ9V0mcr3qD4zV0zto5u2NXicZ/J/ZGjL6sZgrFaCWZq+M3R/q
5nnkjgrEkQPLffRBLyBHF4BdFSqSDam3JZu4Ak0BxXD+Fnvt9vs6GtTKl9Gjygtj
zr2vc8Po2mvknukpKbxKCe3jqx1sQbN9ccPvJRiIEq6Bp7Q0M8i3KcqMkydsiiJm
5Edq6H4qIUFWnELmO4ukVnkPVjcyMXEBBcw3GFKQCxQjjIZrrtjbHg0qKvdpHuJX
JohADo322pwKz+aE615LqBHX68I6LXc+Lg3Ui1fK6LhMUmIid7UM3M9SI5AqiIa5
mC3hih2qC8h+kNiPi2DnbLohJFyQ51E8Lqhiw/yOSDKnacUl/Qc+sr/0tD28qjuV
IGVeCxoIxWjUs1sgiHB/WfUdn5SEocalTvoJorihy5NAazaJO9FUTV9lmGZvhnuh
KVUhUsVLF5FzslY8gQb+faHsQd3d1hR43azsyzTucavE5W+0zXEXaKJb6kYlF5YI
FGF5dktCO+X7q93SIFOFdVVVJ+KtLK1SPv4zZUB6eRiymVm2OAOKoEqrN+4znwu5
4Ab+IqHTKm8ogg3ie2wKXw3/0Wd/cYZwmBYqBeiIpwpIply2SLdrXtZt+TPMN37X
w/DsFCJ4Z5U7YS7xpn5svjsN/00YNX4MAinsWOtu4RrhwZsLX0NfhGAkjwMLTglk
XkAg7zZcev34A6AGxPIjeGy5GgdMM0TD+TM8NloRF+o5Aq28GzA8nYGTYv1oZwlq
uYMsK8GxGXcTiJ7KMmU/BDFL1wa5yk3M7sW7z13rkMFNYQa7gKgbu4eTdr6ptIVL
KhDg0AH1/FKHdmqYso59kMddl7eIGGDuitM/z5yUuOAX9gJumZYRkvfyAqBIpFP0
LoQ9ljg1n4EK8yrjinlXenveoNvx9UqVO5B2erHNsmB7mZMFpgLUC8LjNrSMk346
Mm7gmRMpEY4Vg6S7Jj0TY+wl9kose7S+/2hyv/fb+Z94M6xqgzsK0JUumwolDhJh
JO/RPKl6Eb+53Z5m3/t/tsdOB5zVWWl3uXlv2ewmKPNQZlZp6X5Ia/JXTvNbZfWg
VdkiHDuFZ4nltjgqAhCZCcO6dxGPV0Und4cDgZOjqbWBQFxOcMY54vnN99gpcUga
nscjRYEz+OhNVdtlgaJVOa5XhWZEiVZ53iTJGZ1i8WOho1w6/+mnG+2Avj5iffo2
987xVctLx5OZnQekKh+pIevaZwhNn7Z9zkF/XE9USRCAgfWbcFlJfr3odfl9r3DO
gQ2sATau7Ss6m0n9JH8ZXzKANJrl+97PxiT8OAT/dWxkf7kZ4Qa7w8z43/F8XGbK
yjtsT052onXHkdQ4KwW/d8HiCac6XdztpGNOTcm0oN6OVzUVLXLXjFopyuzeYmK4
2XU2DpSwoBqFZomTlA3kyNBd8zhd+yweRniyd+Mkqvp/NoP3CtVSUShsO908j+Sm
teY5c3nTlkiDzvgd+Ea1dIO9s8x/ZFpQ4o38wvLQPb+HF6b3N4pDtUCCTj+wF9jf
87+rfOcre9qWxBuHmwMWLlTTHj5Ayc+0Oa7PHpSlqrhB1trjw0m2AkcJmGrBSMxy
NMv0MXJvBPOUWaEs+zo0Kohwf33r9I0kPsQ8SUyLjpAeyx2LB7o5xxucPUxQ5rvY
uKhDruYgirOzunwRShsA0hL6NmyoVfTw3psVg8mTvffqL33fSa7MEAcMoBYt4T+R
3Xl0wSW4bXf76AG0iLBquSIuWyGIwfZ7/MeGZbnjW/7tz8FXtJ+XbCVndVpu9TV0
KHvGmOnSQP7OWGCOq/eExqWp1I5XW9FxHrIeWctQcBVAQkNmvtYc5Y51XGfM0X4t
dUepucRLORPKSjwYggBK8EitDTuC+bbT1PPpNzCkvRbLVUZSIJGM67rwrge8LVyL
wfBhp/hZbLUkfIBHAAD0CnWnJWBZtgh2+1KruiV0u6S6VqFIdwiEGevA7kFOgnqN
yGrqiZBaiwN8MSaKU5i5IQ4cj/FyBlyR0WkHONSLK3s5+aIuT2aZXclsavhyfOJX
BkCm8TXLGYJwRcKuA8vS1Dpv1mFVj4Lp9nh4eKCOTFzgTV9sLZvP8jhGn6BeYEff
wS9fbMawrg4wXp9H/c/TPM0zeD45KAq60apei2C88WjuXduixoK0hFG20NOGFaFh
sZpbb/I7Oj4ZW1ZWtbqKCSsxfSi4hm5FjBXuqNREKtvOE+vXHAIDalmcSU4OT1/p
Y1g/zOBmSQ4EkJHYLovvVfMZfxCXlT0qhPXEO2aa8g1NUxynOAWEsPs5noloAUEz
o48wceC63bMl1K1f6H63Q3MtH2nqydYfyds+403Txx2nIs9i+yVU9NztDWphy0nG
pLJ1XWCATLSshjW7P25fWz/mR8Iv+8QpE2TposB0OvzUqFmQVdutw5YPqGM/zWZT
ZphHr9U2n8RZ3iucIRYj3qmiRNIt9T/uBJ4x1I9UTM58Z4XZ5edOoR+AjnoYUsuh
lIqnAUI6OGfIwpwAu8d9tqPMdTwHvzskqRqm+1ZIYOjkFMWbrqVFc6n+UIuALWfl
ZdjD4H2cvQ5DrUyE95VmitKwJouvtGmSAkPE166tbogV11cDH7dB0+fcff8WO/nv
tjY7SPmnUYaU4tYOEhabhsAXeU/1cY4Y5zfOXqDONcG/qcPcq5JFlMv2k04ACzpD
8LCj6jS+xR+Xu+2M5Ero1tYoeAu2DDPZmWxkPRLtCwO+8OiqLn17DlxHIhQ2tN3h
1gzoJfOGTad2CdbCbQ6A1GUWF7vDejp6RfWuk7CZMb1BLsAQ83qpWdJCwccrOL3D
1OuNONMA/D7fNy2EbAWmhxO6Awwfl+/W8j8yKqPQtaF6mwjucNd+WfgdPgrwzwsR
/uBCnsr/SmVWpPwA1wGL1SxifFWaT0PpJT2Ccquch7qNM4X3xl+7aENog6KmtIaE
5yaxdRbwrahMAkiVZMEj7rpP5Lz8XefC6/VuQUMqKBCKqp2rUB2jLHQmLz4oA22p
Q0/sbwHXhxlTTeanHcETPoFT758m8J7akep0wmLz2MUqIIs3YM8hP0pDRCOC9KmC
EWD6wKTPTi5MO5vOHiYOB/UbJl6Z2VrMH3A68j0KzyDEPf866lT8R+422fcWfHSC
xfhpmmLstdJCK9kpgXKHXbVV831HVxbgU+SmoTb2wCXn0pcOjn+xilcBqb1i8nrt
DMtybEhs+PkDIwuR9TOYwBs9Hoctd1TDo3ed7hv6ObGdh+Y9QdorgM0IuVUXHNio
QNH6PxqwtYspE31gc9p1TJdV3etkIp4SWJRROPhvAe3KZbA2BdL9wUPp3/4STy6P
V82wcFrBAnXfXt/aoI7kbexQf6E5py9gNDiQnBJoNKMOKYzPVjwBQZnSqp3VKPjL
L6s18DX2+208h2GzqMJjx5qoAxeRD2L9Mc78MEgyO/1w8RSeT6gGE3j/J8KF8Kd2
cfLe59HVAom0PN2E3wghuMUmcSjGUy34iCmVbzCXZ+weWezaNZb/Ef2Vmz3Q5Gyb
m/z71Nd3HREL+2mi8J3NPJ5GiSSA9U8+4c3ojnoi1d2KACEW0uZ+/1pUaNm3qLJV
ZGYEdXwH0TzEgFDRNgme3EF/UPV8Py22LpMzyRGtmKFFCLeOtu4oUJmqea/BcdIU
gP5TTtAUmi33iwoPmWZWusziLVoeNK5vDaPbRBXZml49y3UoiJ4LaQqUM7jjBeNF
x/E5zSNe65/SEF4P9Xxi3ag7rBuedmrwszPTzcU9IpFHFr2sEtN336bGJ1g5w2yF
rznNDwbdzGDsm844pyWo+JElU+Jewam2OOnlFTj8j3nrjDQFKX6tUkX/dKcYs0pZ
b/IBYZKu6bK2dbHZAgfcqtTUMrcx+FScYMFYqLH+aAFx45YPDWt0GZQpB/8xISJL
OzgsVEkz6PxVv04IFazT39ARDXjKG5r1+PhJoGPay/X4VLbokKKaLCTN+bZCgjLT
Rx9foPnjrgVodmH5BsOK+YLLhoY2cK1L6clHr3nYrXHiEvxy3/6jNKzvczbqEO24
P3rNpBk70FaaMdmlVdcrX68ynfhgvlfExRTx9XObusuIhUJuZGKz9gB6SSH5sWv9
woWllOa7j0fLAfnIg0eC4apKDQEA7c+onhZ+4UMJyjRmlj+SlwMQmipLpxvq+9h8
zhD4P6YX1jdrKb7IEnUfjYcU7CPUuJ+f73iX3PzKVqNjVYjy5Pga/j+zNW5xmq7W
iY39LqHBn1Mi0KtQewhVa7H/odKH+9oGlJ2zg1XzWUXSMvz3c7/C7ezy/nHKCBCK
J0h+3042byPpjn84ohGf/7022n7QvQzM6Zdq+Aynz/bzDx4p3hQj2iH+XGI9T1M2
1sxhGtTE1SHID4/ZUgZF9ybHsNYDy/Tar08gkK3JBer/gFwoiMs/6AhlVTG3qvrp
54TV3KaGUgGJbbjuLt6/19DBLkCf53nSnVqsH5aM9lNCt0VIsA6N0A5kZ9P675aj
4zyFf5/zcF9hx879oRSEc9pvrBPUKDUfHeBUlco2GmnF+3SWnrsRgJeI6K+4W4GT
6X1Wp/oiMH3luQrqDjSGea37PGC6cE3JmuwIzy3ZnSK/eN2zh21wRfQA1FWPW5XZ
hBFoS/WBdH4J9IIwZwTL+g3seUupOB2Ffbm/Oy28i7kDy6u/UADmfAPBv5v2BpFS
6PTcavMqZ/EC0dBQISRLq6cUEOH3uSBOlixPxkrFkAE/CUDBUYd5JbINOwURVRLO
vRMOWaLm6wQd9NhLGq17HwBpWWKgBduaLMJ10d+25colVZanc5KMWH2qFBi7oBAt
ZydCxBdIvJ9XrItPDMpWGz9i1YknY0IN8/fCLpZfcpIJR+8tHWMZTENNgtnlqM4q
rKelzDi3qpr1w8nCMsdhZ54T8lWpqyYLjimBlOZHi70cnJZSBuT8MvonT6WFk16a
faRtOSvBBVKdQdl4Nsxi51tvZRXu8wUt5ExTFpao4ZYPUF4IsubBlqyaTv+hMP0r
kjmPdVkXrnFnn99q1wo8jWyXCQ36gADJImPoUqNhK2ksFTgH6zEV91WQZjhcbo8I
159RpHAOQbOXUsEMGvr/OEVjo8vM9Mp05QVjkrM6Ha7jdFmC5sYopYLlcKMX9FKd
YJO2SrjiX9ZjcLFOg5rwSxN5pepTyJQ2TlwSbtU2KH66vRfna5GGgE8xbGjAwN5+
fnss2blrCKlMd0DuBX7pjAbnnu3o2dUlFw8/TdiDCh18qoCuaJZLy4TVXyI4hMuP
ffyfD3guqGYz9ZLnvph/+AJ+SzXx/RtWcQGc3jY703O+MapJYoEZsZTG3/cvGPaA
Za9RLkQwcjxrvUXleOjm2RYzAXJg1r+P4zh9ahtHQ3BVYFUXmOQU6+Wfh1r/o81J
UWTBkS9PYOnQ6FddUCI8StMsP7NHUY+viYqFdMQA4oAGtX4WLG8E20PbkzBwZ3JC
wl4dX3miv3dKnc7yupMHd4M8P6mQKf2n1+5wkWIhNXCp8lHUNauMrzBnnTnr6Dz8
Qsp7Y+YFWsXlYjnX0JTns0bVbGsgTeLvLt1zDq6/oBZ27eShz8yyikklpPbOqF55
GwOY6VVFtprmFEwMTH3zmjPkUvEy/uXJzZkmq2holw3LczV7LOO8wDrKrsCmydzh
5BKXTIeJdJi1QnHv699mgFKMNK0McaMGbPI9ALlEIu35MGBm0f4WLiZvjPIm0xgo
gdXGedU3rBzjlI8KIl08qPGMbrYDC9tM4PsCfJC8a+iK0AFTtYpTONyt5ProbT1P
wFb5fzg/hRvzgqXhYTRPmTWpTZi9lTZ20Uia3efbo407bUJAAiv2UvkARh8hWvwD
YjRD/s05BgG/kHtIXgtEHdVCCnaQi6cLWUcyfTENxVff4z5jn8tXcEuJsvbZYQw8
LB1k5y78xG4DiDk2kBQkG8pwIssuXLXCpxyzwbPIeonRmV5c2IJfNH2hzcPqGm0i
H+7fJVUrRY8+WOL/HTgZA2dYP62lUzhLYH8RwZdVGV4fDH4Kn5mm3njVI901x0S4
ySczOLGLC/kVNb0HrV93cJWO/X4JWVje/Tt39G5bI3LXN9jXefOxfh3hcyNEeukh
HRhvTqq4uhBLVYTxSVfj1S3rqd2UWplJaZIc7HdDsiLhcIjeKGP7G8I9aedSe+Xv
d3Pcrzwq4PDwkag3rTQ2sMlSO4xiS5CuN09RpMOGoilFjRJ3zSvwQzqFSGfgsfP0
Pwsnau3PYg4UVsyrh6xpQfEkrRm+XPQ24W0m5Y4ZTcLmM/xhxuyzOZ63kduJjSCr
+KjqSsB0kazmGiDMDHQoD/uQ9C3RLyg6mroVb0n3C/sFFRpo/z6Ri/iFkrXHsN0f
pmbyYKdITIXtHGpWIERvOubJk8Dc5fSDSJYcxQLme/6clONZhvbMmbkaxorGTLyq
0FByEEXPqPYS6SmaqcR9fO/4J50pOF+hwp2EZbVMA5RncpkT9pWztUywKe0w6uXR
McX80s7CP3INTGUoc8INTsnwoB/yKsDhrzBnpOX2NgWFjDFZnN6SGie9fegoxmJ9
RvrLlrSY6s0U5ENtlKAotmbDlKON8oNmRdvyb4UBy++950HEU/LtDIX6oo5G9elm
4diHsjQq2isxuRJwISFhpNuwH69dtUyCIlrFFTq7fNBZALirquab4Nq8UKGk0CdI
clO6nkDgcv1zRutmyKoryAIGnk+wxhE7CJGnNIixVu/h06ER0BDIdgNKGxLpEe1a
tTYatrcdvjzokacmbl8Ao2znM8YOpLhKKT3g+nZFhWzxe/J2a8AiH4v/2454S1MA
n6pRGVZJ0gRD0HzkwQQWT/vXU5ZWMUIVn0qWxYhCd1Mhi+M9/4tOigA75xAOgP2u
cCSqhnV+9sCu6Br3TN9MAtVzizH1OLsKJ40OTTt+wMOGwqaGmrT6xPYk5YlA+M3L
Eo/W/JlqadM3+daXtoQr3wfZYAHnpgvCcpNLYi2Qq6FXtHuXboysTSHYURqeH8Le
/NRdXZZmLlkjHTNVQC11Nn1PPGf3Ad/ksFa6diZSoDFqUFdRbDI019kjp+PPIdC8
i9Dj5R2j6AvPXC2h3SN8vfeXF5s7wY1wMWn4z1DlPtrrhzfqHRmdfbNni3pmnUGR
/lzN3BscIcmPZ4kp0VDmGhvlDi+zdzlZx6TYoU1f9kdry4epicDaJCyI84BpC56S
ErmWU+P7al1dQCSOXqqc9I94ltOxaq/4ickkWjT/+CQs2Rol0JYcVKA3ZsctWA2b
/0iOTd0On6ew2eSYxFCbyzLG7bEVUFJriFZO+hbSSPAFZSITQ7VZIQDDxhnpbXpt
ON1l6YvVRoTZF66dCB/36mJ4txDbI96qSnHaS0RytqFAUZQPCUTM6tr8P/KRRrQs
d1ihaWhcQr4BWJpIUr8is7/oijdSFRC0Sw1IyCBsOiakDCSyIIlJx3ku8XZlT6ou
yQQ41kWRxnCiLg1IGOi/9PRojKPW8QWwYKhvPa/OcWKtmNdD2bGTUEkXCN5MXsqg
y0KgIupT4HNPWxGnG1LKBOpkOcNbrgezQRAdZyl9Elpqprhlb3p98jH3s3dueDWj
xNqgZmV+YLfIrz9UOwr8KqRlK8te6lYnvA/mmsMIcahkd4MMTHUMkT2mKBHqLX5J
jOGEboYyzYEtwD/jqjmfcfwElpi6zbXdPNX7dwlVJV6UPAMUqDCDeR2Ey9NCNPf4
/j3dbP42bGNqdJLdSJBszAwkoN7qhKIWk3oUjUgfsnNgV+TDaTEV+afFrlAfHpkO
8MunJlwvQ7UtQ4coM2Yl1mGQ8eiAFm4jppo0mML9J1G2fy5lnMxBvsIopQfISnq8
U8eQRp1332L7be7F599RqzA+RbsF2Gom3qdwtZS9fkMMVTne8eTpC/SERHcoFGg9
EcGiqqAgi3X43LPkVoc0uehoSiURuSEV0WqXyN7f6nXFUfCxK1ERqdEm0c6SCiPx
UR31YmdK6/glfgkBSLRYnsv41pgUJGiNaC6sDEVEfTAxZRIAxF3+R/aRtMNc6Hpd
SSV0VrRP/fKXI02MbzPSDxWR6SnbRpblDV8s78dXWmXrlot+vf9ewVMboNzNxx4K
uoycyVGU0TTm9U1GBgzmZ3jbRxlcFvcDFwOTEFc95vLr39ewxX7h5ABvdfvrij1O
bSjIojTU9uCpoq/sCE9e2FTqbEz7k9vBS8Xml/Ioy/4AHVInIpNMOCZFMKPnp+V9
bMiGBFBf+gkvrjX069FndDJdgiyZMzbhHuojSdMf9JnCFYvzMYnPWABjZxGcu8y+
jZA910xYp386mmgKTUUsiZiDSzUq6hPvfNzURiK0vRAPuRqhc4QFbwwTnJVx3fdz
qs1YjC7BTIQbLGtrjrovt4DrNo4r9fqlWIq2eaA5PDrsyv9BWHQXsGYKatTqyfyt
LuMpq2qKqsnuFyF+ux+hHm54iTKV6z9GirWr2TlF/+7NW9/8fJ8okhLjsNjnRMAn
tn1hkIqBpkJnQ6NMwPgleo+zBJIeTnAKxCiQTkYGQTo/5NfzBJ8UipfvLQHulssN
93W/GZg2nUZe53nwHN23JJgdrUMXasY1JyhOoFTGJJ9L01iYugqy/NvIy4M70qS4
q8qNgOBnD0ZYbvb9Am1qSJc/iMVoIJsxfp74rmgh2lucguUDnPn+a1nv5WtnjS2q
pyThMjCXX2aUJP9gjJZU0PcRsGnq2BzN/6BI7jbbEcP79YlvF//x733vt+205uYh
0MlO1mHGS39VLXW+FRZV09l0VvYnyoBFW1YMpGdfngMHPC4JlA/UH61x0/zHaYdZ
/99bv++Xz8g09RJmrVSqyRiYBOwS0Hu2YX8qlOYzvOCnxXwjtNgkHfmwq0xGI7VE
QPVuC5egLbg6q8GbjMhrxpHGFUsPViGwxPjy2vBR2akB6Y5pnAIczGRnxeXzfzEE
2GdGWp3O7o7C9XBWggYdgXcmFQq8/2sK8D3DW5b1/Qu/d5kmmWEe9BYutT1x4h5J
+QgIVtMRryErs5mkdH3ljfPEfmUvRKR2bCZjz1ByYS4NRegRB01mjWBQjB7EwmLw
kfBr0YED/8ogrEPorjzreIcrR4/48QAOUE1zZzQjXhI2xHqaV1yaaR9YKnLQcdO8
5D1Mi6dOhom/cqmNAt5pRCN1nLwFUiZLOOXkIPz7EY3BxSUVZb0gE7K79CyMAMLS
m6bM+CFnwMlr1fJBrvnpeDDtvOd4/GG+HPnkuvznFAoi5aDIwHaewt5MAC1AzpVH
w8fGMrPkHPF6FUw6M4Rj+YaTWAJujzEykT2i4UHhmF0Kbcdom7JLFtC7qNfp+yke
VddnePyo8WyWkeusDpiAmcvD1ctqnuuWMIJuu+fsXn69F/uBAQpSv5Lti6e9ZubZ
Gup/YzLjKCjPuNPUztUMTtq7BiSLhGHRuMGzN50ieYxXVcTSZD8f/uxZxqF18ip+
OnJzQaPsHzpJLKU11ejrb+CxPe5lE03gREdM4NbI1shvQ+rbveK3NxLF0BuNUvBG
0zWrXHPe3lFnQzbJbSOY3mpZdczX4q0TPKXFJW1hUA7kv95l8W8har9jXycY8rZ3
C3Vvzk3CcH+aq8Bfsy0Dis/vCPw9UwjVOPF8b2HC527vgOti3ImttAzZKPKqGQl3
xzDFRtCDJWbVhhRXJqniFh+R7aajTVU8NAl8P4JUVkJKFg24bdM0pdEDiPEdyIPa
ijDUBUohsE+z9yIUDSSi1O7Jw0yz4tE4MFxbdjv1yRTlqi8Pc0THEUg2xkr00SWM
zBOEx95YUsgc+8Tcq/R5EUgWl838RC2Gscv4vLGo4lI1tdYxhe1Nu6+kvgVyqQ8Y
QBjVcK7BNA4wwufK+qck+7L+bVYv0UAFlDMYTTm7bOIMtsu9OlsOEUT1C/Yuk834
6qxsLXJrh87TymH2IgPr5voA7UQVPFvKYiQHNJcUB/AijaGsgZMMnAsAlrTOzm+p
tn+yIncjktOLvCXUi3Q0rg39hYJzV39/QI6EFCtVUNY7fEDR7pfD4KT1Zj52f6RI
/t1lu/Ol1/lDvmtQ425bjbpL9uMFdrTCwnsZOKzzsd9p1JqyiPx3Eo12bVMLE7Wf
Od7Ks2Y0C9C8brvOEBmnSW0+aKFoiiHUIl5a5xjvpQq1DPhSq9EvHaeIDG6fpVAT
Mt6d8NfNw7wT/tUkj5jXaEqhwMcftVPm2NHZ0KNjAAbfQU9Gl+Mmpj04PvCXF6pU
DiIfUdAAyPw0oaqNnRaWMRwkuk+oKlKIiTfAbmOeqJ3QQGyqSFre59naLJptrICn
azXLazmGggtEPJO+pj1DZZdU6C/LMVxJDkrQ5F/L3BLkwZIBL+aMQqZP1b+TGah1
4JoNrra6bfmeHDjCyaWhQs0xsCNA1x7xWPSIqKMnH51DPgtGfHHQEDQ7GcP0na9t
Ah5iWs9tkG4EYW9EqxA0Zv1C14FZynxxxn134hssvY8Y7cHL1/UGttH7Zxr7MJ2o
lA6QBhBVPXpJzweu6tSixL/9W7zuSmLXQK7HTDCvl77IF+IeLYIZ1uVXlz2Wy16P
7073efq952jRKwKcD95iK5L7ouNugN1J482Uqp3nWftUIVGlLbAULSUzXC/KleXa
rue+CqkBOK8Bb5mbNGU6yPkBxq/bdR4Bsl41g2CYIb78w1ap5PcocjFfMeRUBxkw
GONp0EcPu8tqvhV9kQQIuetmxU3TBpfxX3mBFGA/ma8PMYYiMGrKNF1kBADbnsp/
a5+vIciS81cbpXU0d2f9vZ0r5+q/1y5MyMryz7tgxGtjR7HrzpcLbsn07Q+f1oWj
H8+2jKTilKHsoXX9yrX3Aqt2Yh/wTlhDf82utL4tu/WrgAcb3YQM6bfh4LhB49s1
1igd+CLJ/7fpdj1qOqu/rcwRKWnwC0iEhd1o+OKlk1EYOOsZW+1gkyzd43scjog0
oki5Kd4wopHzmC4lqwTSIfExYLIZXmilTFRaLpiGrJOsTIf1ONNb/O84Ty5Ciskj
mYQh0+pTWCvldAVPhyxOCLIl8bH5GBU13/ymaPWTkopVWsqY8D4e/5SuAmW6yqYq
Tug9yVBvSIfdhPHeohftxerIWkXTh4rPl+fkDShGKwzSRvG6M2AROBxmFKGCMfFV
zm1rU3kqSWUdwtNsiH1rrltGVQmVqjQKEv0u4qCWhCJReZ7Zl5B4JW3F1eWh6mhX
U2l94DG70kDktlyxIWNudBi9GgPh6hAoSDZQC2IGIwFE0eM1p5tlrkwskFr3nMZe
204JYGLlwGXMr6n8OX8Hf7qXc/XTCw83ZLFarC2uahrlzal8khyYR4GfxSu8oZui
g1P4xIgCKp7xuBCMmOkzUeO0wdoqvWJzGQ+Ea7ipbGx1HOIuYL4A1gjcRfyVinq6
BWKh/e9xe09ktkYRwttEyuKYxFVSBomv/+m9I9JmEBOzABensXlpSUDx5fy5pI8Q
q1L8P6TSLcTKlZKq6WSCLZu3F1UN8iGsQfn+GNdcCGpe2qfKqcxgTtsYLSFbOg7c
UrDSdkrK/8ar+yPOwHw+hWVFy7P/pE9Fmh/t3khRfxgCkyi/xVCt8uxVSbiTGThN
27jEcSEh1yoWLEjy4O4FOkxCAw+/7m43OA8ZIQa8c0Sw+MpjHr9lZGfM/6JhMcKl
txYdzHTeqb0W8kXNi0dvTPUPF8iB/tnRkHkDP+6OiX2sLhS/DNlFEE0Z+jTjOzRh
CZUivSe1MCWWIifMguLOKQgfpNHPLJ42kO/WJYb7H+hZcnYMNrFTNGi1FTZFgnur
fVg/neaYdcHKrAyvmD3ipbXyPD3NSHHO4ASN0kOKyc0eSpPYIPNCF2PSiSr/ditO
t+jhpoHS4uuj6UCCFira/HgxMOdGGjzZ46r08v1EzQRbMlOkhh6fSk9D3Djb3bg0
G4cCn4GAH5gly6p/zdx/R1yEzFM3McuE/AQ0ll8c8XGkeTRSCV82vcGEu+71lr4U
1cir9kBmP0LOL1RA4SGyX4Va/AfEtqaPs5DTLlzJ6ihsY+X09stUsbrlVwV0na3F
ExDNidNaG0Obe3tUIBrRnEu9O4PjxwZKkZi7dOOkwgza3A9Jxf1hsiGWNcDhatsN
np4OCTFqJzfRW36JVlQxc+nPx2vFZtSO+y0cz3W7BPJLsgqMnfTlL5vStFiOy9Ta
KkHAOPznnIcQnoCCtijrSjf/qdVKAvGI1PtoWKuE5N73W5Xw3z4M9v7T3/YYYsCj
ExPy8A+yxnArLES1XChd5ML44ImTgGsMIyHH/M0y4kueJYjhQgtoIR9Z/Pggh3kS
qtX3N3EDxUhlrUrSwPSYTyN2TJ3GarRlYRhrQcMw0aN7oT4tp9FWDchm8Du6l1wV
iOPBPNXcPEWgYMNH1GcigFnfuaHG0ioEckDFLNqnmK9pvbOBtzpfdzstHcUC3FY6
yiL0VaMaRVdFYqhlob/AJHgEujAOJj/twJzmejATLMXYAU0rXG0mjuVr9mIi8MNw
bmHYZ9tZK1b1jezPCEbHeCNssIy5nivd7r5SxlzUdEHKAxqeyeXW3nuGQFsdJ6qd
JjyZ0F1PD+uC8pgQ23rf/iksbD+pfl96lQ07FT7fwCSeVCe0JCim72euxYq/w4Fw
WLl7Yiy2gtbbmb6i4Ec4TP/OQf+uhArMdPnzhRzD9+qC64ZE3XCG2/ozq2kU2Rnq
gm25Od7xWp03L/+50XkNQR3bWbt4leGN3xkX4c+V3aGwdwt4GtlM3ICDwHrpU+Fb
24nJXdatAl5Ak4LrIhrSI4n4JsrA63xqc8f6oJJ+v9U51246Uwvmm+U0jRz77pGo
5BVXS4unJHWnx3Xao3HP4S85/y/lNypGhio79Qd1OpbsP9x3gpkHIpeMdh379g68
2jTazRQZaGnWztffAWzdU1Lo509fOBrEnk5570NiXsksnaUm0VeZd7PrQ8D8FuOT
jQ8633Bz/kBwePZIn039P7b+hP/xSFefzLCkjivdZ+w6F2UnPXruBQstawu2Hxno
d8MAu69v0pdNe/vyeNAm3V8uxTmueV58DA6A2o/lDjDipZvPWI5M23beruGAG5rt
QrxVqlfzqaZ12RSKtWXigIq4gbNhSilrA0NlnxIFTyj7fKXOoOOPj/30MFQjGptL
muEvH+PdjREz7MK7gu9SVeDCLJ+4BBKXdJRvVPYA61bdh+CXcaFGS0cUiRb2cDyE
Sf/nBZLkuIGd6iAnWqfzukU5VlooYd7D6jsBKxjsLgICdS6w3+9dYs8YkCc+sc1V
5ETwF7hFo0ubSmqEMMP9kWxMkSxfvraimte5nXQr2j4R4y2cfBCGCk0FTujJu3cV
Aba+w1/8lUYW3cQgi2WzKyMe4Teu8RqIKKIQeKjajYrDaCveMyIc5Xqm3Dr35xdk
A3jvbHf98347CGjssuxuh8j3aT0XGnq3rr05X45fM5iBq2KQhPK1gG91lccXPdvD
ON0nIitmbCSx9suC4kCyCsbui2YjxhE4gMTm+ArH0QaWFFgcixV4JK78DNc/J9Ee
8K21cuqDL8HU1/TIG/KSJznp+AK+xTSZyPzxK8K/R8ZA4TxWI+/fL3Dh9gXESVVT
zA3kln7UVja5DV120YhmdsWvyxy7YzinYtD3uPVtrylDP8aZuyw6hilmU0mA00ie
RS+AdmNbOBjIIaDTK+FSN+2PIjSnq/FZJnDbNMhEExaZqny//Tjmnt52biC7Zxyz
VZldZamqcPxJWYU6b1Ljl+Mpu/Oqs383lQgjN0cVD7x/N99uvFNWdenZw/XE+XWF
rObWpc4efb33hBAVP7yeWIo/ERFQfVCHkMkEa+/gELcQHmqm1Oq0Cfu+FFkGTynF
BPvKwwInnnGSDNu62DiXTKxAkKzToiyOckCjVlgmUJXi9S9EuHVd8yvAj325ic7G
w6XoMgZsfEz5JZYXJl6QRhsxulU+LWM+B5RhNX+9bYG9jQIkO+/7aKQgEgFga9/6
1K/tr6UN7g6UR2StjRDfBm455nhUAw2OeTnuwWzb4d7w5dasiXMBkjEmgYsEj8FE
Y7ad8mizFgvSiaLpriVM4X6q/iqSceL+GdwE+66Datx6FPLyF4MaW7nuCkjTH2o7
rKHC7PVJdECLlnCqSaQX2pXCVlDY+8qa7BYbL8Q/JTpU1OpljymioeHQB7PZiYlc
35X207fEu2TbV8rKY3jDgkfJOpbbYOb9FUbxsDu3hMGQs2sDbWv/LXAhcsVbepn4
yErkM5Mk7QaHLllQEQIAUJ46Ru+Tv5AnFlRojdiSt/OD+mWdltFWAu3XEAYk2M11
0k6zbPmhtNKIn/hX8TZCdNCueiMVmSbz1j+IUtWkYODYlZhFUYU3PLGElzkrnlgp
lmhenRu9QNvxF6ueEUZl1h6JmCroDlbD2g/HlFFKjjJOSaZwdQVZqUO1ITAP4Xwg
MifvTTRx/hPqHNe3TRfyCa8iRlLn5jgMwCkYsUUmzfosXHTIIo8mFxBMakLhwTXi
dlk3Bqo3canmF1AjS/HU6ybkbF5uR2z6eZIqacPa8EYqKbHYnep/ChfqmM4JMzUC
srD7QF0fZ5J3cQbjlrrOf6nRHMOxEI4JzxhNfu88EER2JlrlUx4aUq9zIs/Diok7
YDQkZAQqoG0NemPibG/jcr5jgXRX3ICkGiwyEwfgjxKmiNr5K2Ifc8NFyYLFfPN6
kBbt111NfKK/J6MucoKEBi8UVYCGz/cp2cCx4MlH0K8YLE4uTn4n7aUVf0HKzPKT
X1wTstLlIYV29y133UTZUcCSt2nIuHS2sOQ34LLfpacR2WcqdznnNvgeTc5xtc/1
U8G7BM7ZNKQKGfNLjXkY3HMR/iuecQ95ulJ74vVli5U+/mVXK5ZCdzfyVWKJIj4Q
10rdbMczU6yXUlsT9o0I49BfbM+lZRVYhI/nNJnS/o/YkkE+Lv2Ujv5Ly95Yr7GK
NZJ1/3wYg6F/y3KJQSDpceeRA+TO/fw7M53Wbauj1dMMx5nhVLXQ0HaQu6CXoFcI
eW3Z5UYNMUZNtpAfefiQ2WQ89yhtQvusBdjiLxK5P2BF4pmVAs2jA1UH1EbabhXU
gczRpkvqVV/3G7QRtaJlriypJl28Le9uIQW9BUCeqx/E4XTRfPM4p57xgraN99Ma
DbWR+QgQurcjv4vG9nP1kbfZMQc3JyFGouC6cK8hyned710xHg6Xq2M9xITlUekt
noPSCFBiFaeiVjjzWiWv28hUkK03e09BblAxJVoc9dzvxTHPtQhjYWtcl+V7qmWD
cTb/ucEVNQ+98mc0M5ILG5kJP04D8uTnGPfanwQWnHJO/qlId84zOaHUxE+PO96K
QGWCqPQu3DhJz4JrGOc96Gq0UxyRgi3D12+PGP9tU+/gtJbjqbyCaQcty6I2c/40
UOsZ18WWxZjmHNgFOIkqw3xeX4Nro+pGFFeGmFDxSHgjSiBHW9mfoCOlO/EJ4/vN
YRUf79GXEdA2Ur3g7Eu5fZjcKOp3HRlQl2W16cWAvaYGevW4wPFkrLykFb0+JvBi
ZDQkeUSEqV/oJUNMTEM8ADOOvGtuEIQmWds2EnGbqlyy4dU+mjO57ABK+gK7C5+x
ZI80kn6yizuW4pJlckwBRUKlNcOWDCOmMZh6IcqFBc0hY6rJsQlPc5qA49i7AlBU
6eGoq5YRVnzh0gh+SsTtMm90ttOUBlU3pHp93ODVokLRIYHfRneocejd9WenL0Q9
14olJ/1bV56XYWQN0kUxRguNZtehSb8ce/LveEPaT3HUyW05z7poGm23NIqy7Per
cH7NklOjuUiNSbRGsPQoUdv3+h8DHeTDf69jkf2Wi35HOUWdjzBRXfwYK9gWAWAb
z7Ki4eKy1F4hnSYzYWBBddHOUgZxswyLT3i8KVisFlC5HS134CTkZn4/9ySArUds
1ajaFsYZfbx3+vwCFrtVftahY7R3WHqbhLer3lJPj6wdTSS2xVPJ6JKzg47g584z
4uqH6H7WA0CHvAeDO8aJYKWi/Bmher+oGqInIB1DivFjxxWZ9CPAp8NfQa4TEqtz
FVdSwaS0icFuObAye5Y5AcYuUEHH9kXolsT8TyeTA59IZohImhCxYfmSO8jR4iI+
z/oCtfjssecZRwel+NyHE/8Up/m6Y/U7Xj3Tjycyi2AmSgAVEMxMokpxHIbfOsDM
3h9ozS3TWupl2vox1QP5+o3MG+iS42DbN2DCNE1zQVpKGjKucOlHLz7IZ7cWTIEW
qWVavFmr8Pqca8DNkcGi3j+DND3bIb00Yer0Uo6sJIy77ULtDXVMwZ/4lJI9Hx6t
kgoe136a/guczS80TxhtHBuF8sJr+hTTwX+K9V+m60sehfL7oSGqlRaNef/axlZT
mGFD2hgeM0JFaaz/O3ODAKaHeO76qF7fglLFmIBbikkt3RA3dcGNZcHNjVw5Kolq
T+cLtQtThzBoW4taFtuVaWD0Rw++UM/Rxj/k3K28S62X2MAEGiFqxJRQKIdZfl36
AQQxzkooHtubia5HsbgzOc5DyGmh326aeysS8Ji/mqQnXQWpe7hDH3yZP3yHjmvU
PVrnuUSVLg8alHNb7TZnJbnHW08xYF7gjskAdN1Qq7zchJte70ojyKKxuqanj226
MIYFhL8hcX2qJOskuQfvyhbgVNFpuDc6bJun7f8tOc3OdooWf2wvRchxtBT22W7E
d7RRXsO95Bc1VRg5X//RXiYucctyJp/TarH0+R1AFrToq/q2p9FLhA69V35d+v8Z
MiRp891bU+lwQg7mHPLH6S9bLcAAPi/73wioc7rgzczBUBcqY9I6g74POkq+mjHZ
uXqVyQjnmFIkql59YTEEKCFnRlBY6iVjAIYz/dzhRe/0TojaiQq2XMKvaJLFeEsA
nt6qcVK6cNw+Rxh263FsLFqb+pqU1aOQQyCx5oLFTigL02iIn0BEZ2JYMQYVs0rm
OK06D6YiO/FmkxAODf7DrfDPh4FFXqDWI2J4oOHgITyJRQn24FDI5d1YtZsS3V25
pUU4dY3oMC8lD+tK6j3VPU7LZviQdT0+Y794/6RhcHb/FMyfwNo7/zebHkwAHC/G
pUZp+uY3krpYYA5m2SZpNImFcdlHtvLZOCmrzdvS94O/QDAaw6NZb9OY9q5mdc4S
d4K28muSHXesciuY0veIifhE123vlJdCSFce8VpaNWAVaETYNsByN8g+JLxgmiR9
hzGHAgajMdAbvZFw91Lf4u2MEc2XDGmxUKNbiHrAX5k5VE+oT3wTfatUOkffubuF
Mb8tGCfMkA1+4tfUr8JkFyXe7fibgx7oPPTNlkUc14MfAteBPmyFKAj7Z+eRpB7d
CH833xG/ojkJ2hXoV47IDD3VHDfNGf04pNPDtW2IonyoUiVipVi9tZziETTHkMrw
66ma2lU2mR7GNSnmv+wojq9LXzpBuFPb+iTL8TFjEEmuUiji1i6Igs60VfJ0VLVw
JnUdrA484eIvI7fbQpQ+Z3IinLNMJwQA2JVK7bTZVu6KzFp24VPm7fDTpSzRa64O
QciyuFSPFalPebV/IoUcfDk7/pXtTXDtOfM2wVXYUfswxz/MLZgas5LnqHaGIGBx
aBoQvNDXJUGHR5ryFSlAeEESIbbgTb9kAXuPaL2LkgAIRId5YnMPIFPISWmr62Ic
QyEsyJKYw4MgSRzkvrfoBk1oRyr6cooy6pgG/e1PUy9t7UZy9w1LhPbhW65y5xe+
WwhZ1bENzcoUgpyoBEwYwHyPG5isBRUI17DFgLhcmuef455i0iooqygzI8WlLMhO
rpOUlkJ7JNBJcMMIwTB3xib59qrLJKXD1n1sUHTtIN+9oXsqFj5icr3HiiyiUu0A
037KgOIoedF1Qhkfec/tNhXddldnbBIa53pAxVVAlngOY5c9evqsqH6ENu3JoGV1
vZbuO/WziHnaZDW7Q64XxV/AqNPvUFQypwruiSybcDSQBJlTByzRUqW+eGT/0MfT
Vutf1smIHP12KowCyXP6RrsGHafg3Czm1QBX7NJxlOAy3w+KvxWA63Q15+7mSFBu
NMGz3LcUCCP76oOalHhB/axMZYD0ot4IQtfL4dOI4/yKoePdOaLwz1UfdHKx7mHD
mZFNCjUl6FdeNUU5fMCEt9xI5xjOm5XFc0EfgTzufTBp0tAjTb3HRtc8VMQSxOOa
3Y9gJ/jEU+KfhcoOrDQaq34GigH67m5f+Tn3KzMbcS496klGQkwJfqePr4wtaWUY
DxXwUdPq18YECPoPfOLjBKCiEhpop+GrICdZUFw+6TvO8gWUif6cB0VSp7vBJzVw
G/QQ/XY2Cs8wkvLqEAgJ2KgiUQWsVV4LqC6x1ab2ZEXD8fjpn0y/2OLiVyxokDHI
clWHKM8iJnrokKcASBaL3Hfptp2hJ5PRKS4DqVm/g7UUkeH7ajaI9EGd8BUq4ckY
KuhZTLr0fuRLQuS2xYtonzpFzvMoUNZ9qGy6+iugMePCXFglir2AFbzG5ag6TyK1
wDfX1XeSZzgYMhRx9c0lnknsdBPR5jyJHynOgDtMGfAaZpjVHgyNazaZsAUg1bqy
z9odybI8f62dlJkntSxI8vlceYlfCNsiUnWqLcK9I43htWZQzKq3g2nK5coefB4m
sb8TM4t/Hn2exrbe0Pb8kyhUkvpSEhRNPXHr5nlY3kE1H+apqSvjeEkbRqdHjxSM
CWHU3UIiwVh6u+ASkSW1WexsauaWeWy55KmjN0f4HZN5YNsF64+30wVjvkcTm9kb
3zoWj2rxuMgyH3iRYffrbPUHNS9QMQbagVKVNYdZ/eDDOdXpsZS3OQkSbTNbyo+w
T5BIvoUn5zTmj2UP3PjC+e8/0dKLvStvxOt+XmdCGCLulAlLb4yfRYKnkPVR/Alj
G44gF4eL1dkpm2w/lK+ZNFxgVbQJTg2TAPHR6s4zm1+fGeFne8PDHNo41PXCJVKP
cUKv+eJ/2ZL68v1x6nfc0GEcQqrLsthnOxTO2c0Zbmkzf74hf4cMs+wTLbXDRSCg
1XPXCcCaV5Db0b2dVcG2bZ+7NG3Z4xzEDbM+82TCxdubEsf3/4zWthHsBKfwrKH9
8K8ho301a21utEETuHvgUjQisz8oRF0qleyimWy0WEiI/6Ox8wwvaoxauA+7ujnf
6YmR77aIjqrANDhJd60vG83wM3oO2pAuwImwKW7tuFsDiM0TuVcUDSRduoffyFRs
9G9fLHzgJinYZl/T9QquBQd1Lqdv5q5+fETWfg/jrvUwH3cSbKIaGHWk3rAtMmma
BvTuposP6shYX12z3VDXQhaz8gLN3xsMeg7IEaCXvFd5XJj9xOBOcJTqP3ofPPIC
QJv/41CiejRcc/ozTK0v9R6MkfzdsTGp21NBJLrSFc1cygRvlocK2lWGtksu7EKj
L86Sj1UU7uhojJmr9LRbmy2jcNjoMQi4G63nD79wisCVFW1YZPROdfINYjyq6o4V
cc+qw9Fn2VdOBfLk8G/jSsFl876L/rfGejEK0EKnD+2a1gV26yzh4uH8ivQlGQTW
VhG6C7/Y72swcaAOq+9wNhxrneugwSzhBtsQJvzBTtRMMCwFIh4HhoGZBO8X6Be4
iukMOlKsck0t5ibPmy+LK3xUt0VYXPyIEzuGhlmwo5Pzg8kAsP3PZpGYf+WkhleQ
WWnXXFXuKtfKhexzlmRYRYapK9gvoiMkARAS9X+7ORYnNQPE+c2OSF2EU+FoBdiz
3LaOGN3jbJHaBqtTzlPONEmkC3WF9cHytyrhInsyC595y935aJBJLBS4e8P8Z31o
wk7AHO2XoT6FN2dr6x/QXqWPGq5I7LfxREIgMxGFiCZq/ipkysWmj8DuUeSYkoen
zEccoK/ZdtvHDBzXRMaTxmfsW5KnLD8crKsV6oYArDXjANF4zigjVoswyosnPo+p
nRt45V9nNf+JWDrV4fjtSTZrLyihUdahqgh1KzND8Qo0j1aM0W0rrTRoLgQzuEue
rOVP9xwGHaYxdxjAw2qfcB+y+8acwY9j6fD6/pMbKupxBDrkXrOUUKGezbi6y7IZ
oSwWHvhVgrOUmNsrpLDuBW6cZW92iUixlUuuK+tNWJ06CKX/0f37E9fEgba4LfWZ
I25NgZTfTBuSvkyaJtRQ9owdb7pMgsUPe6iIOlVBpWHU5pWJsKY6uKASK8dBMREH
2vXQ42MS6iHU7sKnHWSq6S66Fm/bhmFg3sGp0Z8tSibgHi1WqY3PU4cpluY091Aw
mDE3fTaJH6f8Yu7Q3UXTIYYXLTrH24zU7xsvMlK52KtzYzWOgt3zsHlUxTYhfMD0
vEcRp3H5MGUx0J76cl6F8zOUO68kNeqvVuxLhrAsyLvMVFYyHIs24w0xJ2TiZGCR
rj2EpK8kw6+gOG1V2NyBSSRh+XH9UIIHauO2PL/ezPSad+1zJeDlnZ/f755zNsom
Jn70YoFrjS2+Kzg7Y2zKSeRtdM1Gp8c2+88qlZw1CrW2OpvpA47UgiELETXHBgX6
nzHcGhyJnyDVkyojkDATKZWRbf7mRCgnncr7f24eOkwpjBIQHdBU/dMsWpUDWuVb
NpkyF0mhzzsqxheVix0lBg9kop4EwbQ0xIQzqzcyLfOcOwSng54jJ78ySEf7244x
EbrVwrH/JvkV0YOPIbhFRFjIbOO6j3Go9nRdvHJCS/jv76jMU9/Hp1N8oZi0ofsY
ChPr4SGz8abl+1H1LjUMwqOMoVQzcv0P2TxHxg1CWcKnZKoMgddf/Ibg/794wO87
MIbM2MOySksLl26zyXZ796z8mK9v4pGQB3TeGAvdxOpsCmjolm/7jRivjLDmWxsF
lA0bV//YSu5BB8dVFEtLZpOBC9WUaFqumCsx7/ItM3nlXq0zilE+MjqRYEoy3B/p
B24vysW6kT4db+6DgvLD4rHvGOrU0d2m4mD+427ExfECY/FY/X6PoaCksX8khMae
q77riCSzmTvOS5f2Tfdie8aHhixce4RnGAF+Fgurxvqi16rTwdBuuIWVRytUjN8u
Ux0u1R4bPS9EdmUqNgO2bKNuQpSDmFMu6dyD+AG5gsgrPGTQLOsjn9qYf0Liog7G
1LvB1D4B0MLJB30QYUmPFVV6aqLMQmoG+4vOhyJZE72jsewdNQkWIeRimcOfJM/2
/2b0CeI6rKiusNuA/RcnmX677z1jIMHXBek3ss5/DkzxEFzpYomVTxyu1tP6Lr6/
/wKckmSGhwQ/z5bJ5Im2Bj7rXYY6y3ilvnuyp671MjJHrcl35xo86qQoQdXIHdZ4
QB4gwm0NgSXZRFXVeJu7cRGqTj2S89U0jvqit9zgeGY0RFdOcnJmcTtD7i1O/gGW
t+jXM93j7hzi30EfBOoq7g0VvzOQEqKxqOz8jNYWQZ/qdCcCxRCKqdzIpK6fi54w
QIP3Y1iMI+d1g7sQNUO7DEJfs9rGIfXrq77cD0CgP72uQOwOXwoODnlmDiF8IK8d
yIch7yzZGWAg/+V+wUZvH3STKlbvKCaxqy7o+FjGzpv7qa1ITf5RIKU8xJdIXw63
1Nmks0VCrv+127kNGM/ugiLjjXPWaedttcy51zHyGKOoH/ANe/2DTvhz3wbUJ3yl
/y7RXYAZqQSHUgRxdmEy/52nVh9gqoJgqvcSwis8zbJl7JFedABUyIMh7HhrCBmD
z4kI1c4ebk5z24/WTLgGbUcZoWUxGz7DHkKmyugN2LDESZghLsvPKAVI3d4yi2oS
/OGNSN5K13ynJ6SrmHW3uAax3iPN9/+jON6Yypq3IR+pGI8RrI7aZzBgNAfBnFvx
J4RPXNJ9jVDf+ysfU2KiTP7ricwdLxKmqG/9yLBLSBxUBTI8jOeQXqlNK8eHWYTT
Yxq3dihoZvr5c/Z/Htfe6crX7ZpaKG9XYMuJVh/fEVa40eDdG9UcWRR88e/YTiks
G7kSZWzS6qjWNEfjksxRY/uEEVV8TpH8QYJjRFUIlobps1UhS2+mD6IcWRMiAZG/
7p7bF6VFOqff1E6yK4pYIMPqjWwthP8FIk/L29mv0O17modlgliWgmmL994qJDSb
ZwkjYluBwmwUVmuJjbPkJMjV1CDTQgrm0fELZpj5BTIqP9d/MZ1oUCCYbIgHuft0
UFXOSupnIm8vQ28Lz4uBdjNJKAKlIgOQHikFLX4sLn+o6mAVcEuJB9qsnyhJ/raG
ykoqJTAtif9e2kkkNegSbMUCk28/sFAjIo8ijrgLF06yIjXOkgNaiO7WqVD8y9hW
VuV4j/sjMOkwz92UOAapywTDobNblHB/QdRs+XKovZB/Hxr3/KVTtwaaVR1MYfsU
HiXNsY/9fqY0QqNll5cK1S8etir9VVRaYOq3+GKq56gY/2iQtKXKVU9DqOGTlTkb
vJrc/Qzk4SjCCFFJaUvoFUruoVrCNoCPhCPg6jXYCcd9NDq/N9EQwPF6DFnTJcHy
cXG6aOJEhYbr7qcl6NveuLLxJ4PjIMUdxFZBSrqsgOuPSAr7dSLsmV32CDaCo5me
24ohHgLn5fhrTHmFMTpIb+U6d0AgRNTbvTISp8EQKRPEB2zGYhCTm/5gU8rC2HXG
VkimXO/YQeEZZXqRCZd9hVh1105VqMdYKfqtdJUqQekCsdSOCKJFfDRrCn47oNRw
O+hCN6o0IzwzGznjjepJ+NApYueGCrY/uMnxpm9h9leh+Vb33u7quJa3znqj9DDw
m5l5EumiXU1IAUBS5pHe0k6C8cSDnvZKll+r06Kgb4CO8hgjAOZQd0Xn6Otw47Pc
3svCE3bgrA88BZ2aU8ldHPAe0SU+VAMELsuH1DI+fytvWWhMZUfDMpm0rQLaEM/d
DnJOnMHcbbzbwC5yEevrBHTLn8RbRSoC+g8CUgWoJKZC63Af7isB6EQM7NKgutCG
FZCUkIF3CPk/MJCOZdijGWGwmTE5BBcp7NHBdsAniwrVqDBvZFO2drS6M9ndEkG6
Tb6FaKfBSn2LGBjr0iu8/GDbrmrHiqiLPUN3hjIf0UEBclH7mAtBCX3fdMOkKcFW
pnmJXn2HwW8nIQMJ6HgS3B7tZpfKHnrgumT8UG2oZzZ3VeIRJUNh+mKWWh5YpqXQ
UTThG9LFLXaTqClHHmx/M/tNeXWzx6OH5Wz7KXietz9XQRiIlj/4vDJ4J/WLmlvy
puiphsHvRF756pkydPR5pVNuNo3TnD9V5HmepleGPCCCqunf60zomSW/1YtCMiUF
FKdxQ6SvPEcwOuOosU5hsiKYhFHbPyDxPeb7rZ3sq5QR6XOKlAicOwfnRAnSULi+
2rlhubi8F/ZOpM+Hp2NrbMfcCTcZBPzkeLtrGsgHOAf1I1SGziq8opDFQggczRnY
+mKPAEpbWrCop8CDcAGT968cvZj5r57LqckhQS63oKIL8Wgifs5VVM5XiCGfMwRw
NbfzAjjPPZZHwMX83YAO1u7sjRCL2Lb02GFcn4DCbsEq9Riiw7KVSkACqlANFeAt
D+Ms5WIxNQI3ld2uHYNpD77onHQLp4NqKmauPiioFmXMS8ErPNB1AaMe7IaP4200
potIqx0bKUdVP03mRwn3Rwverhw549xnBwhLFrvWBLc0bZX62rjHxAO48Hj7Agj5
JtbT41S8sKFbb8Pngd9x7XQmNy0cVBewA711cCV25YyWDOjSwhJt20WMhEzGT/P1
pB8B+aWHT0it1UJdV3Rjhivwe9v/bL7aYDH1FLItGBuI50AiCGHSi4u98AwdlosN
jFEL+LFmzuWdXt8pb+NBRUdIeoThvtKfNUoR+hJh9bl4SZF3hMBETprkTn39m7Z/
b8cmRqJugj0QSd9Iun2UpFIxuPbi4dNmL4zXetwzwyvn1G492XMYmy7EzeRMIR1y
xmAfD9MwSKifnpkcEgIwJGqaDGl0FByQLZRwOv6TgRegNE8cgpvnvlutKcfTqJEd
METRomQbF37pbA1I7UBYsgdb7WqvhEALjQwW1f+0VFD4/ymDI/Ot2EmLFShxQ2Lo
78lJk4RPnPV/eOPkKBC0K03bYuAubwA03lxbrC49yAD2ykXFU74t7RH1Keyt4vdB
Ujg2BPBRVjP+UtWMc7C1wScF+9umOAW64bSFNnfSP5nCYeIjkfypljrR1ccTnwYs
eHh9vkrBrEwCsJKQVTjHRcrBKot8fcc/TKFaSEeRskq8KS1DotcMdwM14iZ9HX9g
FUBBljg2d8ow/oq6tGAI2t8hZQ4AmR7Ld+7TiMouhSUMACM7xW6bf2JFMOOHu3e/
pMB+UJCqr+hCqhv+Quj2WpP97UKm9cHHuaNRTZh+HW261xjHak6LZBcRgV6mQKau
oysobYjsFNFR/lreiCs9SSD+a3pmzoJ16n0R+QszG5jQpWJUXLEELaPOej+i/Zsu
xtN97HxSYYNX8Bqv13FQ7NfJxkoe07w4ilYoGSWn1eltx2l7WdbFD9usd06/dl5X
SVHr2mL5UCaAAitw7MOvItpl/daAyMSv8aZ61UmcQDmXGC13aT78XFtE31iQ/znO
ny0VB+/HVzWEgniyOi8X2/IbgkMnn/WFfFQHgnu8g/xFMSU6q2sjK+GkwQP3Py46
MIWBd0aZZcc+7fXjY+x8cPVya0ExUXKC4dR4C/jF1oZHR76cMoo+U+CvZFPj8NLA
yhBLECRQi3vh/s52sGzL8PTkErSTvId89TTkklPxKK5Abd9QLckZtE8nCY16glUY
PIvaSDCO08qJFt3NZJHDuHVbAQellx8K6RHsAo+2KBv9miiRqu44al5xv1VAywrQ
UCW0LnCGWN5KaKNFsecLitVckdDHUNxrhECar40qBL0B+aL3L1AIouVhyD7J8j9q
v8AqmHiNAlkCg0nHj8eVoj9gZQE0HnasXrC4KleGDtlOvsu9VUYClC1TKdyl4YnY
aeZBprmNIwGOlmUVUYSd7167JnypDH78pwThOsEpv81tQFNR23GmfFTFD9Qjs8Yp
7emoEzVBlhrL5GH4t1ZhJSEalbO5U0IO1y+dtk7bYmeN0Wl0tAgtFO1wq184lGxy
Nv+n0QjfVMNM1XSpuX5RJIOQHm9kEfoTCRN0EfOwbSLlG8H0wJFhwFVoqIeHmdrO
6ZB+SplXa2IoQ1n1EA8MXZKZGi6BdmDQq3DLE16J9G+/u5z02OVn500yyPMa9chq
VFfoiwPEeNd2xFkblxfX4xBHVPdAomD0fV5us/URJjBnE0RIYX7QttAP7DVWm+UZ
p7+dOtfLhzdjtr0D5ymBM9PUiJ4B/geWTStWz4krLpK865MdpqMRSkOKDBjl0TVn
U8BpjFeuPeqiLzOMMU4bfh6dIWqAuYBZPk/plsy1S6QNHvDVMpu0A0eh6qHgS92U
QgYrrx6+nTseIntrdmLpCXU0B4rFjb+fcruTpHvV/uHP4vxCGBPdQG9d861mWxH7
feaPte/ClBgDomokG8ymncXXgnYJoqeDNFlynKioxsyxdrBoAgeW9uYfIe3r/bJ9
ed5JnGgxv0qprE/CeUCmPHaFQf5NGHkNtZsviSzBSG/FDDbhU8aqufIsJgueSQxl
QIn35INGmGq/Fe3b8q7kGt6imdMBF90zYLk/jvVvVmVScyUkaBPpnyllpWfj21t7
Js+Uy2SB+9Y98KfLfx8unIZSTvshw7cWn/7mDQqmv9Yn+ls6YB0Tr9iOSijH191b
wSzOYKjJKm0yHZmcst4+GX6pj06Z6nBOK6wXKnI+1ahIL8xOKpUOfJziU3Rc9Olf
wGT3xcY5QVn9LiUU9snz5QVLYWG5Qichb38rx9ETfoUACT3+5rQr/7UIhW7gwQJM
Pk+FHl3mu7ZgL2KwZd0jdeomMwl7MgIbsRUhwM0AzSVIucav3SrD4AWOF+hts1zp
kpe4ndQ+6yrPqfo6OONvHOfsK8fb3HNgsY2Xwit1cjayMz6ZhXj5YKer8xuP6RxS
/i4+CoB+WP5JMlo/EKhLIZvq1Wyrd2OwIa8YD7JCr+YkZO7W6nGjokI+DLtnviiH
H4QvLZ1UqHIPxv/OaQRTkJf0+VlJL4toH9+uZosVCj6dm9RoSOeDt1P5BstWzskH
wZIRtIDMhaNqSKGISa5YkQVRNxaV6NjxFzBB1PCPQ/t9k1dbpJFxCTIG4OqMgkIO
yjzecKpoZOBf111mfulhDG1ojTwKGO7vcudsa2gC7eYVySyp8Q9im9KLkB+xdmdl
hpk9VIQ+HbriU8WaG1/pyOJP/9OBgQ/R2yFVNOy0Ll4U16Fj56e89HqMQl16HJ2f
QVUXW+u43KsvVkpgELpciIVBae377BtDSp+JpGvBp09XpZTYJ8QyU/Lw/fX52apd
Wg/j2gTISuOEviv+iHIdSUdA12+Vcu9vJXEJH34NT4Ofl4w8vvJsi/T8zvt4yngi
3hJuyKVPqiiqmbTjtUN8CU4FCQfTX89EIIcoI6H4lWUmpxSPRiExNbjICzUVWb17
hDORQaXoZgxXttavhT5wHlBOvL784n6RNIANBgt2NdhHwz2WiCLWX0RY3La1A8Wv
tNfgVMMDk/b7KGPSodGdSi3xe89ZtrqBJJ8mxyEoL5Namp5FSCl6U0h1Il9SUCEQ
0j/IjoeWLRvohqfCDO1caTLS7rOu0LPeax4C0L1Otw7wvWpLRN+sl5b3NuuiBeVf
V8njTTT6X+Yk2yY/tcTHEzN9QdY4au8Gwf4UK1PHoZ4/NZb1PBiC2IQiwG01EHv5
TbPqF+QsBYpr/TI+3SYHh9AmQCbpsZkoFSiEFf1uGgiLAsW1PioBG7UW5uWNvNBV
3esHKioZod19BFbjl9Gz10/N0p0W6meudqyLwSDbkBLtuQU6anZZtxL+R91oYQCh
IAQFJz+RqNP1TMXsgUMxRcdtKnFQGVAoZVgXkdrUZU3o5SVulzLR0C4/h1JeYSSy
YANHFXbpIrTegpt8UOQGdcO2kF6HUnltkGMeRVVAC1c9Fv+/oIx59fAXmuJ5ZGZF
por2COjlHHot1rAKc5lps1YLvoIiFU4QkPD7yA635JmKSXhC5nXvsvuOiaCq8for
Z5n4rPfndVDgTK8+hGZ31h2CZrnM5ZtXcGwObN8qQqKbvh/Uj5kG+kzgEQkcyWrO
APrXUeVqD03H7rbTGjZK3VOBwi6YsqQFkjTssBubZwR8ro05ni0JsSCTNjWSMbEj
yg1NOOIwGkQzQuGTdwZjVjTQeekhihFRAiuopciJ/ncLp6KgFB8IuB/+Ze08cIQ7
UKXiImHvPzd1ZDReGxV12/gajbRj6qEWSg7uYvjGXpOVQdF8CmVaho3n5oIOQJec
s0MFHwfRyas91kqB26UjB7IE6rTIAPz2rS5p3c8AMG4334YDbqiw0/3HrkGE2vem
nSYkt0uUGVbC+3qZ9YJDG6IN+ZeYj2NPAwsp/dfPsCu0M2sabvr9ByqGYqU6n+ot
MAlfdM7eROHcxogJnU9jBHBLcGM1Aw/RukJfhdVuaYNLpEUZEISw654AyvqCHCPy
zRCmASctfdrwaAKYRujP/geriIxYF5lkIOwFAJt1PXbu141tDwlhM64NdLdWs/zp
CG+DKdCDZ8zQUzhL3eKpTYiKw5n2XfSCMf73o1HrZ7EErV6FcyyJc4oTVs2rSGB1
OGigCL4U730bjRNbagJK/1eticIyjEM8So7tN+6wJHIwrc30ZnvqDnNuGvbTT5lQ
u+aQawr9SV9mWS2hIhJMU8W2zzhCx4QRHlPQFFD6uQ6D/70jXzbMTipCzL2vUT4C
fGXwbANv5ulRzOWRwx1IFZ165qehE/AXS7dpxtEIvTxinuOFkQm8JphcV8oyvQeJ
cOtXTh4LHcTir8yNJ7xsJvhqHk/06Z2ITyuQH6RmZL4FNhlu+7QnzSlKPVZZ/no/
UErIQvwdUTnZfgrTH7s/93aM7Dq9fmFmFId3230kQQoXrq5NSuPITpkUFJkgr84i
p78h9vLX03Ku13a4anJSj+LkrragukLHUpYUC4qYinmDjWB5LM4JC9BEQTUz8U0Z
8Yhc279Tce3d/YgbzNTYyb6TEmGDpwcbC8dR5TiUZH721WDwixzBnT4eFt3Ltagg
7awlFfoKNmUiEdvXfpR/p2HfythMSBc6iDpHPJvv1QGv5U5TsgAmPNG954EirXRu
kae+xeUxZP/Ia4csnhXjjwKuK79f2d8wweem8j7ic1CvLKzpKt1AMU7SJhdiYfpq
JZg3PkRzxcivquHPm7OQWR66mq3x892/H0rUKMKKIzaRP39Eohf1f+0r4HggiDBm
bKUhaq/QnaDbbL4aOj5d5NqPCJynafl0V5MRHFpSlMA0oHp6Vi1hcF/mAZrUEW01
9tBYFETM/bo32MkK5T5LDpKUFud9eSpknD/XFGJuDT8kQK6QpECBsII98OjY9Oyg
40yJ3jlcoiQUhPno+sPSeVt6tcRkS5IfucX8x00ulQIX1MWZnJgdrUArM9jq3y5t
16a3wmcfM88VEi+XHxejZ5bnYmv8hDblCJp6nNswHY3qzXjJTWa7x5fQ2bUlR4Md
juP9cFTZtWR5Jx5nClkmxcjDBbpL0ZyzKijyt8M/YAVXw1iRpljwNLoOGO3zTThL
UMIgvGAetDvZ16mGb4jIigq9AjKzCXI7U24gt7cwVsJyEKpYhA/iyS7SfV53kadP
Hvb/zBZXSQadUgOg4K1ITa6M5nnb3YPPubxrXf0E7FbBXo0sMRaCoeVPn/PZEx71
dXojFVkg6bjsQwPwh80vLGvKFEBm0jafPyli6USLTUrGxPlfHGAcFOi6frZvUdc0
M5aWDW215m9BU4RkwytOvdFjqnsN3wCA5/UbUt5AxCyddYPNUqkvpdaZDD/ZSnu4
XcH/pMJv2Yq806gVLH9vwhQ9wMP+3wCfXJFjDGdmJfQNwRkW0WDlig8gsawTj42C
ajzSRxL+YPeEDKBQSjR9Ed4AhhhgiaJRo1GyHtQ8hZcTIvIWBWbxvfBR5IJSkpMU
dvqMDOHG/ij2Rg4qgfvZy+Ez98AGHfRvhh95W5M+jd+NJ13HVZ2RVd6ni+8WBeAt
kMxRvvDbXJ2ZHf/bZhFhXv73jusiFUDSSbsY74MGiRZe7Et1vmIPX+mCaD28F1ZI
/wUdwxULhfL2sx1wP6gjAue3jsfgzKK3uez/AKFFSjn7BcN+WyOpQ5+1A6g+Gm1r
Zo5gqpLuDsp2VK1m1T6C6OC2rO2bO/s4BR3FyR3LHbRAEPtZm4+qobVBV87SRCst
PjI5kqN4bAfhayV4++5yghkaAky5J2Xs2gqvD3Nl+ywDVHpYvX59im6Ls5GSy9bZ
MLwHf1I1dNcugJ7PEgHIhjMZbfnFGA0763/+zwzmJUVRJYu0cCCD0t9vMd5uGpOn
KyRnj5cw+RvfgECbCuqS6RDp/RWK4jAcb+nSJBYQJ8YiOba08CXNFxFjHKQCN7Qg
VrvLPpBAWyziZrMharTL68apr6wM5AL/jhSLfpEqV/V8yixgfTdbLVIGArWnOBJ1
5wsiGnqPSL6GiF4pvozF9Zw4TV7Cpv4aVxzg+yXZvbSK7uXgtkV5E8Td53/tmWrq
z51Uhy4KJ4pA+eLsWX08sNufQMa9CGDrPLLqYq2NULVMJRIYc+De2c9ExwnRLiHp
/redYOTBuVKS1wgV+d/1i7yKMpg0tNNFUl+BdS+ziGPD5/DkhtFSCO4uRuxdooNH
rGZDnovZVFDnvyb+c5fF6dSFjIxmU1MForurXMOj0+zDsAvS8wZMHDaAmsRHGIRf
rrOXVLFFvZtNeZ8NdsFI4mXdk+vhZQ6rU1lsdNef1y1P/l+/hhqyz2pZ07ZHpK4/
2p2cAcJrl+dkE+i4WSJ5QW7baZ3ihT5PgfjgkdJ47tJYMKt5rIAZYHjL4K9qcLi5
QP75knd+n5CryRO/1al7FHIG1Lm8lHy+wDd7IuFmLFfdBMiV8WfX9oagcfH8VXef
1lbTT8WTQHjyDoFBNjCkIncBSoGh0NQUIsLi+RDkb7wHFCXCmBpxDoNlrZlEWbS4
FtmrrfT2G1zlwE8Ak3shkU0lgvRJnIoYcGax+6vPoVG5uHPmaVOtKPxiZyreGqyJ
Iqw3cSdrx3EjrGIrlVmttrBPyCz5kA8FqQpSkQs4mOYDjHfbJsmNR+kKmwEXlp2j
fIc/Witf70yCeM8kW4zurPeq7wZLOn4zWEYE5QgUOIPDmw4PmhRiF77Waak8H9T6
1Lx5f7V5PAUG6tCBjPcm5qIpn24yMj83LNhz16ClMY4iTWgH+z/KRghcIb5uwCKD
HjgfbHMpoRkQ//kewvzCAP86wUyQ0H7JKqSgAZsi02ZIfc5aiBrZ/C8yZpIWDkSm
CfNWXeKYzwHr7AW6iDoLDpR91uEvXnTxowvKNauoVUDEpeYXQzqzTkd94V5uNK6d
wFwt1ZaNr0u5Vy8tPX4ucvDfcoBCGOxuPGIcHKyn4WMX0iwR9b+eXhPe5uL5I/6F
n/B4jgJUAl8RuWk7tlD3e+VxIBlGVzDkTM0EXHASNkcAE7MyAtQZGlGAY5Jfaxq2
Ypu0LMOkq6zToPnF7KxZDi8YP+/q4aiFRXbYFnha4SJAMnVlQa1KWyVwBQfkx8Ij
c0OpXM3Tq0J2UgK7Hny2g0IzytcbhIY1MwALLytk/mCkVT/3aqfbC0gBRDgO53DX
nj9WNa3gqASKPvlGOM3yVMqEgog6JOwz9tOXMLF8zFa3wJzaPyt/K2dyCJHQnKGp
VQg/7/axyz/m9yxlX5EYyA47N6oBt51zX/datrT2+YWpDuvToHnWMR0VVPA72oRu
lq+Zglv4eHMh5CUKmmgVMy8XNiJwB7oRT+nHz6+pxkt8JN8BeXlo81AzOSNy8WsU
FiXTIgOAJ0RdP5FZHx42bPiFGhJAvbyLMgadX9rC7KHEET8DWfHrMgq1m+JHcXqG
bvS5pC78WwbIIgFet14enyNBW7aGDBLbJ/Duzp/Tan3CwOEzQZzB/O1NObYYOshH
ADO4PvqGCOyQ14WXXivqL39un2NpIabYQPZylLEFulLut6h77UWzYYAi5O8y9M7z
E2v0JN+/rCoGgRLCyhvVoGUvbBJU8DB9eWpRuTbKnB4kjpVGiolL514udLCozmdU
3mOkiOrhjDoftLvnUhMq+xhQPa4rI/A1jSdt3lYgH0K94I3/4OXvk+ndEB4B4BU6
c4+V6HMbOj2f5Nn88DcGyrvohWqbBFqEiIvuErAkwIH+GkxYtJHxadVTZSv1DHzR
iiDYBHfHyGhRdEdojNW0jpqHBtFG+O9w1Boyp9Npa9G2Fyk/50RYG8MKdx/0hiQo
Zb1lsDpXbn/3MnG9lr7uVFcKsaUqjuNVVxeauhyw4NGZqI2XfQ5vy/sLwDtNjUxq
Rlb0WJodNz88Zni80GmqCv3FrXkUALQ/oHCmPqmFPcVSnEelFB0Sa0LJJMNXsuWZ
teDyxC0dEexVxu9icTv3yBGMrTv8Q1559tJTfZY7i8nluGO/o93dHXllA7ND4j3c
mmpqXkBqoI0zCHTjonj3BDDqk8x2V3stUR39W/Vo/7o1yWOR8eUZlkSnN2iHvEuk
VCdX6D59DxI8PmfkCXOXwQT0NXPszYZNOf5+qUUBrPW2WO635+VUw7nPgoc5pcEv
urdn2aOow+TR3LJ6i9x3mEKVcDVhrkCRcUiBbW4Ji5vQqLyISe+4/Y1UsiqsfylA
eSq2fRErFIzJIYRY+7ILUhy6bzvRNhLj+T35h+hkCwuUxUxCi1l+NckD9llkY5O8
K0HNRCuBiBMs7zgUyJ0dS/xXWApz32wfrq5tR2eHiZxUV2bf2vcjNS/rmLIT5cJX
ctaAgEdDh9YaaZJAMJQJIqzvAaDcDCHXHPW+cxoENd+KvWZfng7XPRViY/OyFDix
fB6mx5Q2QIVYRqkPeJ6a9ix5Cvgc72ts6fd9BkBx+J2G5Eylp2YJCWd31+gMRLsS
jzlevycHjGJOnM0bjHd6cMMWROlKFHXSoNXeoGDgTlcFx0vzUd/ugxd/DXenSlFt
owBfEkxC9kC3R3N4nGAP1UpNxiEw3aM97N6oq/C84/yuCT4JDHokjRk98XJqxYp6
RIBpMzCuQbax18Cr7NnR522R1QyKot04aFjwadSOUkJ9+KgThC5Iv+hUAU7HBQDj
2wrFIiw64nR6XXBzuPhsMSCsYHJjZuPdwGiu4RrlbNYNDm1KfMR8I3qPeblWZwxH
+SeyMGWwideSMAiAPwi+7GDqOKBWUZ+wg8WJ1RaM3WaM++BzI3+sW5POkNvpyU3n
BKxUk5hI0D0qzFdeoLiEaUIY15mnw7iErkryBLzFqb8NJjfSIQrkbzcG4bgot3df
9A6BHfzC/a4minYPaMGodY4+ziBZeyHEIOOC/jxcnV0Xc0pye6z1jYJ5jFXRtq+7
mHk8MI9+RGDSFcXuSCLKgHGAnJWeXOwujHw+lrSzAIFdgwKn5Ppxe5v/VI8+BvdA
IhUaF8Sz4uVUBnrnwYJrtJut04mXQ7FW+biuwWcnG2w0rV1gzDXpgUyxdrJgT9J4
oK18FpTrKkjz0Rp0KlbWluXMD0+KXN2nFmcP3OHiH09gXL+1q2FVZwxKfPke219x
ck6gWVeiB+/3n5GvLHtFhiTdrnPGatW/cV1NDAlirXy0JmxyFl2q306+jm4zaG2T
6BgQQscO3+hd2Neux9TplM1mMY6g9wQohuSk+KPylqHu0RVu2UcjeL54WqRnMX5K
gNGrzZxxemSBwsmg8UcEjXWnFoZ3vYrh9nhMbmD2lxoIF4oxs3VlN7Vjy2lMkZX8
VZCZPu4HqkYM2mcDbsWZdDfWR0K0RMiEnRk8PNraVOtD7Jd70V+e0VlhPUwlCEuR
ot9gk2oatL9EqMoBdeUKED6deE/H0TBbUIR5eYvxBXcghoNxOxN5vOxye7b4gXIj
dgl44RPPmIX9lS3vohu6d5lYExz/AuceSx6jXqE//OlFAdGEFoh5GtGm9OTKT7IG
lWO0S1XbGTeHBrsCGBNN9LxqM3CXN1bTKv+QlDbpVLw1uQaUH1SYGPzG/ZbdiG2z
kAwuA2rxLW7j5Y0uZlgT7RheuuGNTwsy7459597mhfACk9otZE/dJXBAGTkkNNJO
dT8v9Vg4SDXzwgREA5cvFClRKS587c/QBcLtp3QE/oa61dSVihueIDYF5AtYs3ry
Ghx477r5KgD8d5q29k2jEFZRVxeaRzqk/qzhL04qtt6yNBIt6oXbEFXIpgPl3PuQ
DwLoE+NpzopW3huhR87cwgRYAxWm4mN3x6iLt5NqNu8d7pOBWnSwdbnIrt6azi+F
bAS/psWJP3eJl342ul8whexfh+z5S/BPbfAVs6IZ+JjDdxZQPpA3Una4rMC+80Jm
hmSBNxWRxXxQi/8JZ+6eDjAk0EHz2n48zJCcSG5bDiMvxdXCZh3KdvD3q5HmTb1V
wy2hNWqjsJN8vB97aC8xEvPdNIOTZC75bmqa1jcdmrnfoTGlbqRo0Q0mk39i8h1z
7/aND0TEIh2ol1AvitunzsLYGIRmy3FTONTWSpeCzxkwiCS7EbSOmHsemaf7PPRY
uZHfyRb+D+7gs1unzWSH5ACVCsT6uDrm6eWT97Equb9MteByxZmKyHoldUkEecX7
CHIZ3UjP1S/b58q7rXwazJXqaRYmBxHaRdRbB34CGWp8iJFFbarA80u3iUR4JXAZ
UHeKHxi/1e02H/pNRfB5txSRr/8oWJ0EuaMWFk/P8nxjbJmOdsWt9UssrrkG1FAG
RQ9KlIqjuwMTWr5R5rOzm5YfCM/cFq4DL/XId0wam3jIe01LV3Zsn8zq3wmTbMuh
N+8B/YpM5zYXRRZc+oeUbCJAkwG/+sMEWEOuTXiKWrxCB0VTz0CEFlRjIY+NiaFE
lK7QISHGeHOhpopmTnjUaRxAboTACfe8RKzT4JAuh38iFaq9rcHLYA7wdAdr0CjI
7dyWWU/ygroV+c+FkP8qi5o2d32Lc9Fc5mrsKfbX5BmkRDd5YuQr618MPb4sGoH7
09pPO/HMYCM2OOtmbCGgfivrHFmuJy6xhYn2UqFBrYkgzCN2vjmw/npUncX5wACg
I6a9pI7FXdpdRx2CCoyitZjoaz58NX7wKVzoVFgZ/EVA6nWyBR6YYmdjGegbU7L5
iV1iINd7V0pgoFlYOMc08U+MU34G6p21R9D8SSw+UcY+L5EUdHCI3epdNQvEDb0/
jIusCkQzVNTccn1i+5ThtrOfCmoabLe+OO2HULQsvjuOv44aNqAiebntdzEa+6zM
NmxN4lnd+JXYxhIIdW0VEJz0Gc6Tc9nFNFH16f5t2qyaSARGMDTUINk/qHKM6fD1
IUQBuDUAf7HmXWLptvVLsdgggY5VW7dp8Sh94izmEjgwVhaWonxaJhsX6cPDFuqv
vGP58BBpsdp4QHavVKkDHK+uwS14PJXPopgw/qYoOudgQ8ELy17IVUlLn2dEHQDX
tYJZr9hdqaXxDS7cdGYhTGWZy5WDgKZCBZ0y1Pcsq1waMSvEc9eHQbizcfIII56l
iQvJ1uzfooTng9lL58Ru++P7kDwKg/NiBj9qT9DPHA6mWNMct6z1AFazbq/tJtWT
lJangzq7KyvPF6l+vG3c98q8038IK2tN7Ib4prqrozT0gAkXtUnmmVgV2H8ewr/E
Av1cXV8omsagIrO+8O2UqDBckm6cV5ZV7Tj78yR/o6YJ4HIMum1gyyCawwtYhEuT
EElF6KiXBArOx4ayLajmXeskZT/nOCh5LPfbVBrgJTlAT++34gPsm1TzSLa218eC
Kf6GiWLKdx2H4yZwb0PrmPOHlWJCrhPkjMCTVL+O/ZcW+smREC3s/ux9pGDW+XSE
VUsGh6uLldJC1j7LmrAboOjGD91F3NgVDOPeOCaDnTmhI4UcODryz0FQ6LBSKxBe
ONlRRTocWTz6QPIRDX18M4x2eUlbqBwrTRMyge2Wqkyi2szcweT8MhxSF7bfK6/I
i5iS05rbgfLzpRtkeLSzm7H8jtOzhH27vVrz+VmO1zokwMVmt1UdE9PyK++XsF2V
+Q21lAE2+cXBsQmrW0ce/MJOE+zel9McFldpY2e//zp3QfVOVTDtC551xCcoJq/P
a7MMYQyB7ZvKr07RmbggK9xaGkikqOiSl+CldI2sMOmeW94dwZ4aTjp/k1dxODlO
PxbFetqVozunljeXJUaOJqCE8wU4I5PlDhb2NaYolhdcQi9CgnnYvxkeZch2Y1ab
n66BDOvQT0nMi/3x0c6DfMNYxHQeE+cNwmnre1Vz6ZTSfKw/M300dxV9z7HWWSRN
DOKm45TQYLa/InYC3+IrtCa+CwQjNjZFExg2A/wskTDGIQnUgQlpux4YoNmu3TGH
we1TLrOQ0xxXq0CZL8nhHX4ronvt+9SXuJZFJXFvHX/KuiiaONb91AVxIJgvyV7s
bJJGoz+Ff3E0jK8JYbxdqNhDyuE11U/FwWGWsCCEYBxZJD79SHLoNs+0yfL5Cvl4
TzK3yOHy37/kF45VrTnuFDjK61cFRW0WLAvK81ValjElaS5nTFV+L+xNk74WShGg
i9XaNC8uyERmvXkDepm0AoJoSwek+poJqs25HeUiE9+tnjKG8F0Z2l7m4D0fPDOo
MXr/3R9URlzVwplR/q5sB3GZ9GUpnC25b5+DIAC0kluYfvthLBl1VFpfXk1ovAzK
jCbPQyYYcoGuYxq2qQfQ4bard03DJj6tFvFmwrk0PrGvOnVRefFn7YNpZx7dKKEX
RMBtohbHoTJQn/OKm2NICEBlK4uulsbMKagB/gTXtx8Ni3otYMXkoay/1PtYZkoY
zeDoGW03BxtqYtfdb2+iNKNAcoecyZIYmibxW2TOL7nus3fFK/Qz1Lu+DObBsxAA
RGHMLXoBItOOOrJEUCPXudTNFD0sTBDzb2AnGq1mLlGWoLMl5oCthvjq+oBt46VX
xOT6c1JJAjER1NkiudFhsXG/RU1Y6XEZKDShoHMMHxAAWgpU/k96Cn4Bs9/vOwOI
N2mqp5RymTxC1Ys/69BgH7J1rYo0SDCm8zHjdy0tnUGSLTG0sD0RJpurYOMK39Hq
1oHBuibbI3dN97KayZkanucoXmNUcc3tr91G/gDp/myudRAvvvklHSqhxba3GCRS
rgLsOPyxzA7qfif3wsVQF9vU/PkyvESg+o+0ldnAaBGh/2kqZAFrkS1RVOxyC+pp
pgHGNtSnhy+n3kcaXrs22p0omyU4bqnkaX3rvQ5/hfvy2QOAWwkaFjaXbgEQIuEo
dWyC3ucOMR7QAWjE1sjrnlHgY26DzfJqdN8acid2EmCFxvgra3Y/W71+TYfL2y9k
n+6SoeCJOfXXNMdInqJgTXlBVXq28eBi4/KhKiObOdH6MRzXgj63/FWK27ffQshO
KYVEOjDntApMRYkh/Y1fmmEb2qGps3Nk6xgRo/1TpZgeToMsmVGCEqZqBBZ3MO46
eCL/Hf3N1rbnUasVi+ARU0HyAeMTDORuk4NAwEVb18is24DGx0KC4vt5aKkeOENV
PumNbmNjqM60Vt5tQpfsAtTAJb+bVSzkmF3gdYlq4RWk9qlaDODFNdnCMxowrtUa
wHn0aV8ptpUwiUjB5SSImOrrHKfCvTGSU5Y/URk5NRmiq8SLj1jOjzdGtw1Wq1dE
O/7cwRPX1ICzOI4sAVvOv6VyRM7MXC4HIIK58WVKV0qoCppmCFyQEIO/YHnCe/68
T5XcVFLykp9AWdZnap7uY46GhYdNUNg42XCJsHkIBv5eiwaPIVqj4w/kiA0vgIVJ
XuzoUTpOeEeGXJsFCxVoKhKCnDYnycOROul1jCT+bezPGwWax/S21RnQpyQfnhMJ
+GTv6siTVCzhUrzccJ9Gg9NX9RZ13GxSbIFbQjLxo9TmG8iHax4LJihQ8WbR1IO5
cEyqNO9O5jjsHYz0YzG9oGsQjdmVVMFMGYiB2W5ANywQP9zLPyEQNzqigvJlV84m
4hnM1gscQw7pUMYepLSJxgsEjgD/g2+SPfvQlMDxId3asiAHfwHXzxKVnroRBw9J
6UKVinUGXQGBMxmhYKebTfhQU6tlpI0i0ueqxcXTtUZp+kfzpYQnIq8WuXAszUAr
hn4NGaRAZrEF4Uv68w4ZqmFWHZhC7+bWgCeB48ijPzVM8WcnynFVQnvmQu9JCwnq
IHYaX1P24qW+zt70I/ExmCFqSCYDX91C/Bowuw01jSRBv2MgJZmX2L2H4ZaEY7om
JqEhkVUurpCkc7G8wpzkCiG7rinZaHuDXkmHgCH2vm/zfgTddGecjMOJtPPYdA3m
2PRsiD3oXKw6mV1BlbW46OIVl9vDE9XhfdCJDKGDRjMtaQe19jfgbxeF0J5ROfow
kPdJr1SUMJWBr9aIOUxMDANoWUVllPitWvA4yvUMcQZpCX89f7Ks4QePckcsIPiL
RglTfjkgZWbtfexDzKUeakRqFlCkLb+KJgQSpIVN8ZUK2a8MJUkkxzxqVsfz7EFS
X4/u4qZH+tTj99vKElFjop0IzofLJBqLMK2A//p+mmxtVQoA359+khGLE5Glxg6z
KuADsYAY1WwfIcSA8wYV2drh8Lo76NFmh/oNO4LsSEkAVjnImIve03GOBuTOQy4U
WQDLvYXIZYEoj6rVF6Pt6OrOLHEzX5dMFabcWl0RAj5yVxVWtppwlfteUOvF4Izt
UBw/BvjLhSRCdSmpBhAQQu10cqnuteZSrU7zuhyk3YoeUSIzC7mrbn0pg8uUSyqi
rvr0GBXHLR8rGfkIgmfuYqzoWeI3AP8dWdzFnCqFBYzQRmDW3xCsPcGB9zDUcHaC
fjNb7AsS/+jByuNGU6tbgOZO8TfCaF3e56QyJ8wM5ZtDU6mO7EpYt7kY984J6IA9
HDx4p4mCUZC/Bjit8swAUc7N+grPlcos3bVj6E0CnfoFQev8zTz0FqEmlAtmqajS
yQaAnK0+XLMeB09qfKUoN2X5AxyQHCQse9YnW7JGxMqMtBOA4JeyeceqFc7K6pcQ
Tgy5EEE3Xfpsi8KfSxa+7o7PhuHUFzp93cA0Cg1VuzPfz5Xg8sxpqydXenE3uvzt
9uo08qxjk6MorTd65T0adjXgWF50Ofp2Tm3qcR656t47Gr2OKXj2/ukj0RV3SOoK
PtCFbv6G7BQJwSIPh1u20e27/yNjmhW4ElN7l04zsWyeVvHIWyQUSetwC0AsXj6L
ZnE2izSwT85bOC8ibEAS+6le4MGKj13yMB4LjLAvW5rsvrbC6Oh8keBDvYzbIqih
Kvco80NJTyD13LBQXDewzSJHD/6vJLp0Xujgh6gfYc/YodizH2MgRE/L7pzqy7ED
W+/KKCss7vo125TpwcgA3AtZQFVdaI+ejFT7kzsSp8ZghirJ2KYg6OfpX44aadpM
XcY6gHRRQP5cyDNTo29/W2fyAkUKSl8RXg9nV6o0/IUfTlz/rOUuvf9L8KiLYki7
xjsbMnm2YFFK2Hzjt2OvIZZllL4X8r7D9NkV6Nym/Yqtro/iKWLbZk/FxBeoXUnS
DTFHwxCn0MqhFSSWdWbeuSzzMnqGalNUly3sFFPpg2qksTfv1hwumQGESgD2rsYy
Sf8CHHpv0OpgNkgkg9zN5sFbvqMaGquoVn/CCLim37j5COvrQaywXbrPhgPENO5F
S70SHbwWTTH/avxgNNm6UH5L6hieBLsa4XXbyhw70vJXAiV5ANn4kA4vqZudmK3A
jqH0UhcYG3j7DzvRRzJQq7g3M7zXA2eg/Ud6r8EGgWoKrEDJIU4KRMVN2Y3hLeAz
RsVMLhD0L1lp5IeHb+3sFW5QH6V35gx20iX0CNcqn7dM+pyBcGNr2E+7eyVuvqWx
DGmzfK6KhAnzEtbMqueJhgJt1GUp4PLliZnS9MbMwCjp5O6uOV0PMdLvuP5kPwYl
3IC+xAKVe6bPDvCscnLA/VArxrn+cZbuvjhibmN0s5E5dk8eZQcmMqS1uNCwKvVq
uRjAnXy1x3Bp0ASsrqnbrhQUe0HAajFTnAV/Fbj3jndStPkpR4mWdkVxYuXeNHr9
PUrVMJs3a1CGeDRkKYF3PxpYYzHj/XEvBcZJRcvSV9REtjnF2loYDugBc2zK1l4a
3erpBZWnjaCEfntRy5uWSHcKnPg4UBtfXwNaXSsF/YD3lY+MLzbNsYqdrAehcMtJ
CsqrRACvKWpNsMvGFxPnUyZzLMuZrrJ39wwEnpTjcXoWnAzOrJRQKZdmEhLfkyQj
gf5p3SHg+RS8MtaCk9VROEBvf2Rqdb8uMvAjbNgyv9R9alkxdT63ORcLweBwMyIE
95QZW2NVgyoOsClttaF4g3TB4o5du1UJJoDfpJsGN7nqD/oNMRdDcvjghiLhZw/h
D9cVW9qs2LIkivnOBRzAm+v47nWMnY1HsLQvlx3N9xAdFD5t0K3XYwodKyc8XmGm
Pal0/JETZ93OoFQqOCHNd4QLJC5R2GUw35rNnzZOmBJaJIWw+CFUHg3A9cMas8v2
d5wr77ApT8bHDEf0AvTvQVuzZAhNnA49ttsTxjeU50n0aDM3uAOWN6Y36ICuabTE
8a6K+MZTuUXaMImGXpkm6CJlGser8bVxrPiVaokp4CVYzopT7ubw2GAl+/A6B8Xw
yrlidv8LwP21gMGfY2uWj7fdJUs/L8/cgCx+ign8DzcfrkX8Kc+A+qJOz6Pjod40
fbx3FEpEaUHtS//k4aY493M4dX/UuowtVkFsraMkN69b6jqx3Nqko6dBsF/nF7Ix
rdB1Fn8kJ1Xai0PoTEkbcIYV4IOZwtaVkK9sCe+g9IKmEQvTbV0/XeymHxmsvHf1
zxeBPObjR22+6i+35wHAnjyAbucttTSGAVTXZkQlukma5uiahLBHidPJZbOwVAnH
sNZEPkaTfA71gfOOSJnLlX4l8I8Aa4ZMeeMtgJJmgKwoLkOlGAXApunqx+usPyI3
VidrSXO//MguquOWIqTwGH+loe1YYuPRuACnAiGvJ99OObBWJkUZ6UnPRi5hExEE
cpdjW8vArFfRVea3Mor7vY1NoOw1saL8rqWjQopIYgjz+rXt8ZCjxPldDDa2ifHZ
gE8odKtu7hEiyV/jRoLsMxeZWS+WDy6vnTgUpLmcjDe/kQmSiKqAv5MmLnL+COSU
/4tWkh/UfuwLekXT/cPqZzHvPIXrFz0XUoGpabAe6wDUg06tPsJ3JP4/EzFB2Yoa
eEoOaPFtNkJF3TdHfsejHSzh3XMMmmzPYfi02qbgDDYO0mcx3ZM/w20QqoiaMzhV
M16CrvefqU4I1HYc90RTLDGeg7iB7w2FauOUZiVzdafyhInMb/mgaip7IWev5L35
PcBrTnEhhbBWsdXlufZ9VQjCOSaQubu9H0/8S9wKdt/VzbPU9hkAkAdoU3MqiWmS
/aNZ3Kf2YjQZQnus0EXKFXWXXzM2Z4zrzeE265E8m8x+NSAS5RRfO/a+Qnq72ZMo
+enAvqdunN1iqQV3HtDXgMn8yc1CSlf36qJ+IhT2HmpDghAXbuPdRdHWQEEOrQmN
fT05HbZ7J9YnNi022ynRLRJ9BRBC5xUNxPD/2jXWJxBM2qssk5vua6ULLRluR78M
fL5BiE1PdV1cOTu1NcpA6VHJo0C6mTtPWISvoaz/0SWCvjxw8DYNoemH3OQ2QZTD
yBLifobdcIZW7Pd+bW5Cf1BzwNr7nJMUzADGI+95ue3a0+BZDRPlJsZYN5KMqMpo
OCq3T1BsMuaFjzEtD2DQYeVy5ysu3twVd31Z9mTfTUna2LyNxXpic+AVAkMESc9L
YX8DOdHwPJNst7kM49wdzAWuQcztU6RTKMAZOwLoPqwIWfLyhZ7hDPdH3S3ytfSO
h/JeCpzLNGLfCAHez/82r5FqIe4kuvzp27Jss6/wzP+YS1UwrE8020jZqBEhu9h9
m02M8SvGW7PTganBPY7ZyuTKt2MKFRaEudYFztGBL33xU+6oJCX7Dr8HxxbbZFk4
RhIWEFaHm5ej37BFzp21MDVqNZWvpBnvmIUCguJ4dPzf9LvfmJoibcSxtQM5l54z
iGtNTHhh/VJdZpy3cuy/bA9cu+GbHAGwAs7VfnM+jF6nxbgXORtOceR+cc9ct7tX
chCW03k40W96vz7VmW7NuLmAQOi//PLGKX2+EEs/bLIlZfBtJGE1UgJ9mmxa7yFF
6zkKdMjSqEqLKDF2KTCDAxxSvqG3dvKeN4z8P0P5twPR2V5iOlR8NfF7R7mPLJTV
mjbnsVa1icYmzdDj8J62s0DfCq0ChKj6wTKMP77aoIe76kpBbVfXclQt96i4eMd6
xI+jr/xnFY2sZSS0IQbR25S9zbQOcP/nkj8p+zw0SGQKQbHj50WZ+0j5s/fr1KUw
1cqo8UF8+khJiWD4wBtXGCUe5x3jAnGZXCMLIvhoZ0fvXL+j3LH3z/q6edfakibw
yJNMAIPLtmDxGCsybminypC6dIRjokIvFEKyQEirT1KHmNLlpb4r+PrqhEh6tOSt
9kbtnQojNj6si9b919WUelzlcbOYfsvMS/bYHXCsX6FZoIpx+o5RSLGgViXSlVOa
BgEMTlc+W12WI7pBelGqph8ZnxRCbcOv4xQnUNybU4NUJH8hG4G6hgPVTqfhkSsM
Z5w0YdmIS4l1goWganlNHGiFpL7l/6+6gerdC/ka4kpc5tWHjbzSgpn4IruOQSE0
gP2NytaDR3wptX3bp7n6WAcoXsve7VsJkHcRywWNHb2q2JZB2OT8o67CY/uUVPXq
yXevGcd6ZmJTl9ZlizDpTU/mhJEwAB+T/ra4JfIIfMaxEj0v6YrXQS8NkNNq+ir3
03GWyALA/vZ1zvxPkGtxGt/xyv8moWzI/Q5RYKXeD3hL1DhbM3485UHjnrLCTWvG
VQgLwHPiplrpGJsNdch3PJJvpBN5irI0rjJ4N3PR1vbdVbs9ZTlrp8O8l/rpnDaJ
EtmNUUNQeSLz2m10Iyi6ICh1Ib48x4BnMDoH6QHBL6f7TwszoSR0N02jQMxNQo55
SG2QM6t0Wm88ygpykYbcZEcnGYzXbWgJWdIoykwylR1wIP8oa2sXULgpz8BpK8m+
fnBvtx1Q26XHBuu122giR6UtkXYXAGFF/H4ZkzSWEPfUMTi3QjXjZ95b5h0GXUp3
hAmQ3+GdidWqWOKogzJuYQYAcDUahCURBBLjriLgVaCYLhhxJaunUmDSozU0lGG2
/pqoIJzNHLzNHRm81ziRDzN8GinSKs1kkwvLo4i/5lpRRg05wy/bxfkd1IedqjYI
0+B9A7i30DLEvB5xaan0pnyjDGe8oXwQVSZl2NC5zhJFjGP/C25YtwyArWAnPZwc
4Mlasp73uKNvQfbmf8aUR1k1puYt15P2m1QEepuEOf/7ZUH8tkCsP1N49DRQdys1
hQVbIsAKjpkOEr7vLxLOmEOMOVTV85J746VEWmCprEV/YqxUVd9rnZWUYkSoCmYs
H1uZzSYYzhevKcSuR8xhyPwvmtsGdALGP90j2rDxFhdCUj14lJvPO3l4kb+0HQOO
qTuC0bzaMovQ+lC+UCelnUX4DdKMq47ZdR+d8xPi185XMlrdpitoTBSs9Y9VZffV
pP5I82DVmtFnInMXuA3myFNOD44g8t0l8UFll5Uq+8EPp3mrCuMWRsAJjEH8nu3I
x3j4uBcdMbJ/VDjV65/lgckeHY5RrrUrKkAFjo2rWDPORcbziZD2Yu8quGb7qH84
Meh1uXEmFt2ApusdZB39k+eMeCP5TqFJ2DqcV+H+JS3ErIfq3/I1zVqi11QY77nV
4KR+TCzM0Tj2OghLQHRfJcbLozMUDcGndveeSawETwq/MowwBO04HvjNfktMnHZb
7H56GXdkFIJWBn5MLwJfYj1Oz1NX55JCdSdhKXa6UZZVUgmEp5qM928do6iROQF1
DdnxZKjB+arNh93s7a4XBfvMfRf+igGoJzoAcuBckXwZrDEHS2edTPIbQATH16jt
GwwDvH23nCg63nfx/pnNqzPLfycOwIJjNMhFaGhWEPGTHbDRfm7iSF19uEPGHwlG
lqIKzrhlfqy2qlfYKkBzVYecG3ddp2VGBwMVkQr60AEVbnV5LC84GrsWIsMMsWG0
ofEE+0OEaP54mWv1Jvj+ktLRopwKbGZCwP99SmXbIQrdGbnR8GbDbSly9Se/szh+
xtb+Fx1AwQMBnmIZOTVrs++JNm8b6csMaT8lk2V9Au8HUYJfCxnQfSv1tUUyufxL
XxCKn56D9lAwELGaFYj+IRAEjJAsf9Hfm0bVAETB68oQBp4cpuWaVTUdJado7V44
Plem1jJMqjmp8O5mTTQVWuaac1HdSMytymI0XLp9DuqrPpbFTC4FIqav8F9xLnQF
isWQbjsrNlfb+/6SN+gjk4VI4UyVWWR74mHD5zNlZKvmRXn4anuurSIV2DEXBfJV
qaDfweFQMVbYGN8S8uqaksse5D+INI74y6u2LbI8GjYEt7OC46xxlR6Ihf2UMmUs
OOydpeqTGr5cdcE0LUF83i7OidQFZpJmQrCUh8AO6zjFbmd6bedEbbBo6kXchPUn
2VI4im41ms5FeRSPwwSn7gRrsItENVtUtWnlWvKjL15pZd218p5+TcnOJu+KYFKh
VlLzY4oe28+IyMyKKGe1COYroCb9+W6WYe2v8C1ec6JPjJ+BzIrhpc6KW074BbKH
Be4OKyecKBAeZjyNRqhP4VSa1I+kverdlV4S0TjP2HP9+eRhgapaSUTJCX5SpJc9
tqFusHlmnYPf222hw5TrmCdLfZ7jxV/uo4dKq04KhPBjJEGDA4840g3maI8QI/2J
ey8N+iNQ9y5HzJHAF7Lq93BKHLeobMd93mzWnyvfGXwn26dZAikwWdzcUG8hLOXT
9E+kIZkuZpsI5K1EHJHZk5oAcTubAhG2Obj0bQSwYha55ypdWxGSfE8FMUjLw/ZI
xoLRsvlUd6aYApJ+ncRsH3XixfQo6XtpAujkTXpcHans/HY57uuLD16CyyBpQ9Ow
R00gk5iq9nf1SPTBzvtSTo9T4duaMvXXvn1ogX1G5+qP5MVEqKIXX8OotRHAdCIF
h53vr3Fibduq3wfu5ufDz2AUe3N8bxJPoUOuLgBOnh1Pv2LBHM8SD2RCJhZhpvgm
cFQf6zpRhBK7dw39QzcDF9XlUV3PiGH27B0v7nnxiX1JTLT6uVPPQBzOJj0VFNAP
hS/aWdX9dxzPzCjCnbuEik6WcjBMRxBfXNep6g5eA1ooA23vTJeH/uDFgdea/crL
pdAObD2Pn8dzOKE5WIagoHmSrU1j73qOSBsfyh7dltHugmTlwXJhG4Jv39A8+q6W
qq3BHMb1yfv9GGroTyApwC+uf8GugknQ9GFtEnTpRY14Tp7oc29BM6x5J/h6INJM
KqLJP56kITMvXNo8XI6kG1nL9FXJxIbxltZotD1beqZ5Qbo6G6PYAiFMIR0NvhbZ
XwpLjks96HFcQZUZnvMVC8ZCXkbx1R1pfzsyLxbuj4od8D65W0elk43k0e2RvB50
Uslhl7ZYdu09I6b2J9+yPGb0jjdKxzIM3zuJDX4ff6OQgjjzKKFYfA6Jb/3RXy7z
0kOQNlK5fVLHD37WXTernC2Ml48gDsFgSQWykxpbwQO7Xo9s5Cjunbsf6KhptJyY
2SyCtO55pGh52D6DOtA6eL14luNtXt/nkk+Sve81iBkmqOmL54LCPCWMsi47ywu+
isgkBc1SJtgpbUD/XNVld6b/N7ktBm/IAoySxtZZsC04KarVU1C4VXSQ7CWQav6s
CaSJH+G88k/v4+PEzMqQVJhBshmfMERbUCE+KHLkhNxEFCdAeOhihQaSEDsaFP8B
BHwZt+Is23EYhSXI/jFlT18HCewF/C24f/LMTVqz+GdEeEmMhm55ORLWjUw0zQGh
3pEyWO3QF/wDKYOhj34bqrBpz2NbmSOycVYwUqOMMdTAf/g+LhKR6FD5E2xYe5+H
scheqWVCA5Z0wi87EgAX3kcOXRrgcC+IQuVxk9qdRakOR7burN3aKmifdxuDcgOl
wacmYbp6MKAFiHUms8TxYIWp4On3XQSrcKIL3n+/j7kQJSmrNTXOvFAn63QloKy/
SykXybv/aAdQhHEH7DuJbR3JL6Kl1Z121MqhR6pleHENNU7jpd59HwdtSPhmfCAn
495he1Ki4/xjK8KG6NPu5EwFULomFPI4y6EPBGlpu0aTkfarrpB31b3SeEKq3Wk6
0FiI9SrRZxdpvgCnFFa4tVF633JO8izr4x0BQUbLgNzIauZMWgC2dr7hrh8qV1uR
bZv9nB3wTvHWBpX2uk1pfQal8CRdDH2RcDO7PSLXyClz8vzlQsh45swfETTOLMMD
ysXSyN/Ubrb4ZiWX5k5LWcpnMjFk3c2MrHtziyVi6zHbXe8Vg/Vy77BtlIKLwlT3
odyInSB/EXuNpYj8NF+pU6HBzsylytu/AOTsGMfCDpiKJSibPSDBXKDT7Wlm6hJu
XROAJJJNWE/TbdQjWuJMEpxKVpFLREcOjhvRUzXo9EdsSaqwNaFxu4Thkc0PdlqI
LWg8EwkG2sATHYIYwIruarTeM4UW8FUyxaHLJFah8qIxy/zQbrGqLwWDfc9UnYQP
q7x107p2IOITHKR+6LPHTBAeJyXP8xAXE657vloWwHa38XJp44G1FDgcYZRM4oK/
1tzsivi2WD8ZzrVcEtuSHj/7sZ/MBBQuj2z9oj/1oayVMvxNH0LheeVSRZn+HGM1
ObqqZ14YVI5UNIz5kg/LiLdWheeedasfS1457OEVXXICiH65va3E4AOunsmxytt7
R3V2hU+KCCuKYCJxpZtkaS9qRRuT/lQ8oGg61CCe2+Sd4rR4yaW1jP9eFYTGu7kF
thhJGp9yOsQn1NjB7G/pPSv0oZiTvfSFFpC0xKMQwkE+dHMtCsIU+flEX0IP3yiJ
f4Bh8dZvuykkRMrs+7qetjA4zWlzvo6DsWnUZPs/OySx/BjYgDfu9MgpajPfzKXG
sfVCnip7yz0BPivtDt6viZEL8UJKnnUZoUC+qmaIJVDlj0OzZhUaM5iIhq6+96PV
0qSxo3MjTQLmvo1FKEuTCDQcf5GEFDkiMmuN9zJSL/55/cygU0CBStV+jHB4uUJy
0nfSImJpMXN33mD9MOTbxEBXODap3BY4IgMEuMEs4l6lMJjxJSL4TCy64smpXUfw
BfzkzwGL+dGcC6Sd1bhIEyLMzqrpy+Z7ARtJuRh5SPns/X8PauAB1x6fN/Q0i5Fl
u9t0OCeb7FpbCdDWEtk239wVwJTUHS6fL9sPD6aby0fOfWI/aBdelWN0w6LtLO11
GDvUZt1/qRDAeXQga4GHfbVf/d4CesJ4RKeXQgXtaLDpJnDDjuhTMH1feZrsnzxT
ARhrHMXUQJwbjYeSbQHHCYcCHieVYFIwkG0slnGn/Ba8flTEScjVjbGTnwlz3BVe
m1kHxYO7nRWMYnUqrn90bTxiSqj7lwj4INkGWVcfmljoce9pIJN6+GSmH8iQkgiY
sks6xRYMNB8bH/NpYFRJV7jdl+89wbQVHqt6yg/GhyyaBIRxyKEy5S4QjZ3TxpXj
54xzbcWfAuptkAq6gSA57Q6Lu6GuN/p+NNIlYxk33laMPDWfEljyM/cdS8k1qLZk
LNMCSRXTgrOv3Ov1kXn70DkbjN+gFU2dIRtxl+5uqHkb6zyPaVB8R5wgsXaVxphI
q2/3qtjnS+JaVh6wUZOoesc3wPgwkMdzCdqlLd9DhKdW40BLs8OyB2FsOxYhDdJW
f8clrNCdadw8kZOoOlyT3Th+MHpEDlei9WZQLKXiWKk8Sc2perbAgRrXYt3LkKvG
nTPERMkuHI6jP2tuSz4RNa+3zKVXqjGutkjCeXez8asCQmowV+1rruT+q5Csdbve
KApPg+HvBa5lN760uET9EOQCQDkxbeLhaeKq4pnjHD/RMUMRgRuiurhXbHHnq3lv
HQRyBlElYTOzLROpqv9Uvvbt1D02134gP6DXxc/mhr0FJTTtwzJ3nvRk3UuABcR5
FtBNIKoeEwqBwcIojGEdKLdvB+InRuKFGAYrEp3ltj0HDjO7GL2USo9Bob9sLUij
+mKh/SsGofgS/QQnX9XDLqrglbg7iBiJ5L/MNkMJzC/pvrCJ76ZfnmmIXNUIOu73
ubB633nwaEsE7q5FjiPJBuWi6vidTYg6Rvb0dbFrJijYjdnxhZZ1VTgchcmyr/Je
rTPZS5rm9qbh7P9raIylEHe0RjooW/LxvVxi81jL6B8eeWmRJYNMvG1jW9uqieD5
LhcBUIz1+3pdm6nHuZ4lycIKYsOK/HYaW6q2h+5afzIBWm4i2ALxwTbTQrSh9LQX
SkrXwMVX0rFTVkaSeAymRXGFEfJ6XdxuUXIkdE6MlqlWuPZfWvSqVGMq7LeWOydQ
+v8F9NMSqTrMOIw89DGxKKlbtyHjGmKCe7oz578aoPK5M+idPE3Ji6Cu1g/1ucE/
G1WyLcU8Q3lawNmkOSTU/vWcZO3elAeGFls6eKA4BrZ7RP8qO9HP6z64TZNRIU93
36apAS/1uRtGCFA5Uj3UfDvlxYq51g4LY1xdRUb9htnI3dvt593BpYTC59zlxCnj
OvjFLJnATKIDazvsqSJmWQ1MyXt3/0iPHrCvetTOqQqx9NBn3wdN+ACLgenCCg/u
81oSHQu2xudrU/d/nhhVVkbN7M2P61vs/SDrZ+nnbrhe3KIG8NVn0V121MYrghR0
h6flDq924nox3p+jFfk8VfXdjVoxTpnArg8rnPDUpjUzyWUL0I2vut7cD2Hm/2te
3NmQ+8gUYAdUM1faDc/I+iuc25+3fKY5gAr6o824IuMcH2N9B6SC35Xf72K4Yh80
R7nuyP3g6ccSMgpO0ZLhBcF4m9BWmTXecalryFGVnJ8ASxb0JJgkbZBBQeuojEPt
bMWJjoS2BNct4ohtPSbetblwWaVFWBM+vecD6Ca3I6aXyUurMajlLUoyPIWT/jb1
3nFMrq9rCAhEFhD0VqVMkhsrNseOzxDNqI9kftL8xOBWZDpMe3IOMk25KpEwT28F
n1EDpxHyI+x3USjGmm8E3UMPnt/hCgVYlC9IkeqBVEgwdQVECl3Blz7dFjBefyLv
Wpd78zEAUtQF6zBkLMyVbOTXcTbvFA5eV4NQ9YCpX0jhrTH4C+Ty6OvVBBLpGeRl
ox+ZgoI9uzeNm0cmN0rDrv7j9z3q8ZNgSzahC+R9Llzz5+1uEiOLYV7hk83rOF1i
ZF2VwGyvVofqC//RCyYL1Chek/tfDR+Loi09iv/nOxCCleZ+H9t0/oUqlAO1AU+Q
kY1q2Vxl/GPQckqnohfrsqYfjAd3VtdlrB/PTDgDREWa7n4/Qq4CvFngctRDmU8U
BsafjyaMckeC3IDQWtl8/5srqO9nxzvW1kY0ueQzrwwtgAWCkVXW4f6R1ZuRYB7c
vTwYk0o2Yv3+VgJnTD3w0IjQ/CWuTrHS6R8EmsVVUpgGtGubkci0aqLMNyvdPdUc
hATwa4o263qIGZElNWbiuM4NDs9z3/YOrrWnkBGVlIMx8EcDUsTA5pmTVXfxNWZo
PyOen/hoAYjsIQpuw3o5Us9GSFPPkVohzSwsXaXwRzdTZPmwZZGeLFs22sQvcbV5
u/Bb6IxxFN9YGJQ3LdUkAWAjqeW35PFbPfAf8iJhPuxHaYeTACEgWlobPh+PRdQm
QZcj0up9rCBFdULvPXDYiG4OEkovitcIxm2TqOf6J747ukV9P3s32pJn2fb4/KJ+
47y0ZDI7j2c+iwSoGAMSQI+JjqBzyxznDufnFfnQUkUvzbkVKaj8Utng1n2lANBq
dqA73+DoWqiyJOitpfjO2F73D72XSoKOS61aRqnCi0/fPg5tz3hVsZw/WUVx7odv
6uP+r39/iWw6J/N0tUluDjUtA1QmAfN/IixDlrtXjGbSqGrMAbSWrKTOQTVXsuGW
jWs3sGpGWHZTKxOgmlH1a7EfAsYUrPszFWso8riD+2Nlz7sPb6yAlIUxVR0ISDHV
wNJv2c73NpUleESxo5s2Bx8+2fzjMT8Mh3H4hANdacgA/wb86wM2Nn+HFPpTZPHF
vbw8rhYT5yOW2nJetBBvV9aBrPdti2NUp5zpzt/PlsOGRVdoCY/1TbnI8yEPEO7X
EhjIm1njzSdvMALJHltiub7pQ88tQoPzScu3WwkgxI0oSPDtaWcMuNi8dK7Uxt78
zyfpJ5QyUaTff0F/BfCAhNrdScWH+VdKP9lXyPonumm6uC7t6HQskQcB5Whw6Xsl
eQ0UZt/O7n00LHOKPE1zaXs5DNQcajMX0u9eH1p2KpjxRicjTfiwtoj0gCHcpBKf
SE1WEu0J/Vu92oeVHe+/qT2uM/iDzHYsNa3udMg0qWDzDKAMaNLW8OlOEyU7ZKd4
MtMLSLpv9peo0htfbs1oXG77RgD4JL0mlA1MXRwziD49LORnj/ZON4XIOoQC8+UV
D9dfQQkO/sM9sIBnGUm6iY2FffJ+Oef+56q7yZXUKyLpDtTdbZ3inijEJNslpCKH
4u6Zp+/E1I1A3ieN3Wahxp/FDP8YK75Le+e9mNWs0Vl+MftT3BY4UBGyXdBy84el
QB8VbDcLyWff4pBBRueRx0+o9BWsLRX22dwHyH7vnaCzaKmJ/UtDdUS8sf34IYSn
eoigRgk4FPNJUQUnkg7Ok0TXcekGRB2lmj0kfJKbocgY/ZY06J6r66+zF8P7017y
GlNn6Q889IutXGweqLGOeSCHfH7QTLOWardvd/6IStftRRYKj8NSDN6MMB+W2pg7
ZWYtA/EwR6AjAVPc0B4M4feV0vD8pa6PSj+ceKqSA9dIaBi2FlTY8X2aesAoEcFX
9RdEqjT05MME/I1WHOZ0n/W7JZC7F4efO9zcWAqPADc65+5YXCSTWWT3Pz3RR9Lv
nMdI0xDcYOaNzY0HjkJz42tni6yZTwyv1WQjz8JIuuZ2KoDRZJ78VUNL7fYOEzxT
jUFlDHXhojz4fa9g34COJQB7vhXmmMev3qvlq2NlugO3dEMYT9lbBd1YhgIt4wWy
o5fpiWAS2ilKgL72ubg7jbmFPi3UxNi6l3Sc4cetlOWOuliN4dHHMvalCTmGPUku
7hMDlHFLWLPtwLIcU6U85h7L5e0p6dfZVBPiQr/tMWn/tc68FxTbQTMQnzfNsHja
t/g96IHmigNpFdbrgZfsInpUd5sDL1P4J7sDL6QzVg1kz4EVxE1e0O8nVXHoUl+2
05ZBLHi45We4ck5Z75IdJE6WqhCJAW+F8HOL8q2H3NF6y6ZJKnPc6jSt1haNrwiE
3aY5JLJNAAUJ12Ef0zc+4eyI2VHRTff8h2VOdVDUUQJ9it/fS7jW2Nq9UKynEvxt
X82z7roEp680dF9atPtMXYjWotEJOOKQikvFOHkmJ2/SiWe4qAms6R9VzWYncXD+
YXUhoT4kg5JOwwmAdnmrcKMgbXAl70ToePyDI4unFj/0fE4xSldAE5HhTVWjU46I
EWxzjDWBKJO95sbUuFwWFdxx+i1Wxo9YLurzUE1LiheoSpC8FyHjM8EL2i9cMhjy
96kCoZ/UM8uu4r08cghOA8FKZBHG9xbZq+OAt6IDF7r4/2/8DE+mm6id9xTMzV6T
xy9aw/ApCNQud2YNijZ7Uy9Av4eSr62jmncjwidnnsKyuj5qdPg/hTnm7FPmdUjU
xw0OfviI28zJJ+w1YApudPlaNrqxEEQKhpZtU6CUPjfGimnTdOU3WPejt424AGBx
7L2AGz6TExL+g8oggo2Y8jOs1xbGskP650J92338HP6JLPm73S6QqsNA1MTcqkw1
1n4Y9UJWwFtyITYhCCunibn/bp5a73xbNKx5BmHw6W3iw3fELPo15t1p5n0Ex2KB
bq46Ge/pyMg3PfxLoMiFdVc9FgX5okudhu+i74ijhqQag7czgEnQsdY9jzlffgfv
QvY4PKN7ZYTdbjaiiQac/7ujWPUI7rvxfP6a8E7/WkP2p5W/NL6ej7ZN+cddye1K
M1SVXkaNvvKc2BUMmhEbr9Dnmp69HLZ/dOlk5ioQtKIgv7Jumeg8RSLiH25LA+Tb
ACO6l882/CiUL8UQ69B9+vISoFaMYBM9QZ5S83vEd/4swGDjHnDpAdDFyc0wvHiq
H3DlCQWz/gCU6UYuamMgAj9G44KWb9k9atCbOYMCOG0vcPVhmmFDEk6DMuVAXmaE
2thzdaGbWo/Q1SOyZhut5Lk7jB3kemX2eP3euZiIWrUqnGzZ1NLb+0LdgUx54go1
V6Yalc0/fPYQeQtkKD8cErrOKeApPlEnhV0YoQysW2mCxreEtNlqe4YYmfCgt9mP
PRhO4BZ/a+HWWWcCAz+RO8fQSnp8VuaKfqbZpCQkL8f8j1uI3A5n8qhDb5FUyT11
yvg3WPKnQGqCsUWie7+rvLU0sfCiOSOE4CqdM40VjFNHoJmaniRNRj2b2BGVNBqc
RnpNZEF8ek8I3VPU01yl0G78mWq2kfka2Nh3jGgMLEm/CBxjl7ILyDOImS+OWQeE
uiyLneT3N4M+JvDmUoBxsw42bGEV8/zRtYVqoPsioViFLVNAyuAqcudemh+pYgPE
BVzDkO0UXc2tToClDyJee7CnF3eFRXyNhWxN1iY7aOnyzNMxLZiTBMEnZasKXWgP
K4Cre7HwD1FbSxENfYPOJjB4Kv8XsOuOm5iaPN+0v/nkzQKQix8yL7586Tu16lVF
pTULDLr+gtFWAjtVcTGgTVaAqehrfym0SlZQuOGhQbSE0Opiev7HIigN1ebCCxDq
hgOgYr8mzbHtEsqMuUNoC0rrM0Yv8C+acqRHYKqIlCIqfFI8F40DKgke/DyykrJF
ZbIvI2eKT/pmO582y5A8kt3Gic4v5cuml3xo2q/zDsfeW+c4cSVka08mDE3DYTob
q3ExkydckOnxfmmAc5OSbNayDQna13heK8VIBl2six7M3UxF94h7TFiuMHAqlD4I
kfH9bEbtGH0Mh9IZJXNubY3IfMnJLnfPpMnXr5+MI2Wz6a69bviZctQL0zaj/t1p
H+RKahqoIcLWHaH9YeK03gBv9A+UkYTfOFMN2CTzdiUKU/zKCfn/cAjiGfKGjZph
mZmM5f+wsDkdHaub29VSWYPA4uoqfwwk+2UYmSEK4lFhTVtIb5FNgc1fb8bVycwY
h1p/OH98C0n2X3fY/MzeQInk7BmI8L+3/ryoHnL3woewf8mqEkNx9DKqBIy8Iqk+
5KXfns/16Pt0QGrsR5d9DvCE8yLJwSf2fovCJRF14+McYBU4+mohuvyHnmLQz0NP
vyavuVqLQK5pQewHAg6nyPALz2JonkER/dNIO+eYGxbk7odfc+edUHcpKxSPhp/c
qfW8nGOMvdbsr0uCg6or/Uw0ziQsD50680Dymw50wQtiJmkO6pqNt8T1mDQVZPlO
Q8nI0aet0BHfBMOtoYLdsWFOhDqVn5v25+RXAN3WvVOGpkiuPnlQfApWb4z3ehPh
xmruGZAiE6DZ6EswxfG5gvPsliMuApaf97OTFK1h39lAlbuxJeCTSDzcj4QPEtAq
9eVDU0ujyQH/YzVpUR8FNKjRt7K8MDx1NZzAh7Aulg8aXf0yzNkMSwqdJH6zAhOg
LU6ez7JE1/j9AO6vnpY3tW2k5ALNRwh4ojQD4UN8HhXvIIUGhgBqPZRWHwch9+y9
5t2brB42hwMmps56Eesu56rWR4NQmUijP1T7nuKHSGdI0jI4ceB4XwFCIHzMeODI
fQW6NgdYVHxxsYM/9g6qXzrqSm6ZWGOePf2Ece4ric+ILkN59BE/EZnqrc6bGNIj
8heuzK3xnZVhrkM58cskJS8af06e0ZedVog6AC0trtgjgbN6FeI/S/ap55LomNON
++EJXeDMCPPf1V35EMsSl3EwaTNHZrZcmTQ7iRHJr56hM6rLX0h/iMwtPsfDxaaw
xyUsmkHNgcYcnnVYvDx7ayPsYRQVbX0tCw6pm13SkOh+75NwqdWstCUYsl5cpYW5
3oQuJDaRtQg9k97ihhoOZlHzm5ecJACpZ8H4Ak70aJrkq8R5R2+u7+d21xYi95+W
qTHUg+bROMABa76vm7MJq37dBbK4+adDYWjzUNQG/RFvwEqmADP8Djr/HpPZSFLh
6Hajw8EKjtfjEIU3USM4uJAgYrLWoA+d99MZGGU8eS44QdgcFAYp983t8CKll6nq
Ys8u3nzoQuQWlhpCJ5c92y7bJw6RMOgUPSc0IHSi6tv1oL1v/7O/ErUzKEJqtSTQ
7JDoaPNICnDJG4n7gfnhUHBIWQ0zyQBoCy/6zh4KKRF2dZOZREdgZb4SvhvIF/30
xQ0OcN5MvVkcUqnn+Zt8YiSUMPG7t1qMXNFb6TzS0QvGR8f+mRrRqmu+Thd69/oV
nGqAbitoEkpertPXGBJDYzOZDFDkBpJ5spcSDsHr4KP8pVZOOgKK+czv0wRA1K1j
IkS60vfcWy2zvvEOwwTnJRvI46/m3YX5AN2i1f32tOp0HU/Zz82Zvpyv1LCkkoRP
x98FGWbL3KS6R8tZUXVUpA+BSXfuU/YFpj7wW5vPgRJXFR3V0ZzspikyAjIB2Dl+
gol1wtITZlMHp6ufnSD85eqJXVm/x2T3qlS2jZ4VcFv1TqgIzQTiWCcY0yP2VSkR
g5Si7sfuKPFJ3wVn0LUfAoDuldKAEwlVNZOixqJekwEl27CPZHPlbOYyJtu3L6aG
H1CoCy15fQ5WLOoXJ8uFhuzV9LZZGt1/ZWL0tgqxujTpZb7Ob3s/8p4botwS1lmN
79yNQcz6GvFSxqX1fSUiox9f+HxHHseLbuspTeT2MRF40qo0WbiE78z7yIzy/cjB
b16mDYpLWUbPLFdzUIVbuIdz/zvvcYNFkQtxvAY81J0H3/ZSa7T0899fTVmBWf9m
G71LzzBpJdB78Qh7y7WffIFfB5Z6SQpy80vKqnKko+FwqbfIHAMoRwlD6n0BpIFi
gtPx5ZGHsycDnT6ALZPqjeBIok/KK86CeChR2BUbgy6j+cvDWESLtneGaCXCgJ0A
UfEw0gln8a8FQFvtJ95L07WHPjRpWhKb1GTtUKGXpEgkpieJx3v/TNoDl+05DRMU
3lRpWPAN0oW07o1cxVSfnY+Ps4LFQ2899BAed/+YRPXP328sTfIFA2130GakH3+w
eBRwlJJA8AMrFSuzCox+sHOShblmZBWEx1+S4urHkGKJsLUTuT9KZ4QkeyJbEbvw
pNe/AENPQa6n1Y7ltCEAXSHYp6lWk+q+LZr2+kpPjx7Y+s4a+PYZUYJNgs10dqje
5HTPA3lx1Dx2POkFvJTLTr2fj/qOUkEp/kNZ83iURbtpJhOVME2uZqt10WpDc1Y/
mEd8EEuXp4pKegpAWPUt8uJalVcAuaDuKwUo4odXwIMNjrYsT7viO8AsnqH7FKYc
DhiHbmDlwT9bMqo1mDYF+FmUFMv8Kd0FgSeDug+oXU9akbzfUS6/RiwCxdU4MVb1
QplKZ4ieLhJmz9vEdt1z4OFOUhvzge85n27cG/LoCZBAOKWXaS69AGdqax5UFyPc
xo7huUtokSkKlAoDyhHuXbYt/e6Y0Ts8UhwQV+GQC5SJuMcrtFpbA8PMoWji/2EB
DwHrBJq8mwi0vi1+lTZOgYE7H7VpLFkTHplxL8Pj3MkvnSrPvWhQ6bGaMrnO+CNZ
2h7YdptS8U9li3lz+qaHm0GvqgP28GYgHB9JBsOCVEXe3iP3YKa2vXrxfDVA05sF
ThepXKS79P4GNN3Qh1k9FLIdcz256x1q6h/HMsKVDftyyLqMtPJyNx8MjklRtHHh
/2rBPqmaQHvajscFXKZd5Z10NvFCQfstiTz9R/nQR/x6C94UqV0Hx3tJuZp+r+Fl
iSfdr3ZE4sK1O1uJ5hYQehBfG3NOXId3qZi3ftAQ9oHexjzy0jpGjP3o/pOHPvVb
vehh1SeG0wHZfw7CR0dLf8SCld+Utt5F5mcupqBRBcpPSUD58Vr06JaZse9R8e2G
0hnAZD1mLKPUZqiOFwpOuUH5dNKzx7PsGoekSk9CNKOjG3X88A6WM30QFAGSOiu1
pUgFkPwM1ph8gLzFEGxtuoif9F46fgk0uMwJY1fcC+iMYZbH9OctcMyIT8EBb71H
sHJSxu88BlzQMjyEH4iIslG/o/n8xmFtH0fI+Sqy+jh9GP5Bm8KY/xdHqtyoqGDJ
WsdHpqVuR2h/G6s8nBTBCJ6JWWZYwDPUY/TLM3GRMhsavsj7dPNg12a1cRnQCbKC
jWQ9zNbPo3QP41q0EOl5Mt9z4fzk7cg0RvKNkVecrBYO7om6E79MFIZsfqyYvzYl
7kvGAVKe9CiPN3uCuKeja8By5C+gc5YcLelsac70KAqExJpcB3Dc0hqCpH8WaREz
x/LWP37+uHzg30P6/7ektzosTnjkJBwTYFjaBFQxRDZJR+aBfTGShTuUEO/JSKrO
CusGXf3mW6CI56UhcLhnRd6cAQYM5hr5ARAoLzLYJhwuTqVi3mo10zwlKDAN0ji5
Tl0hpmZPnptpgoGZn8hopSBHGoSu6Je5AlNNH8WFIIQWC0HWrk04RPlEmW5XWAKC
Kl7bV5e8s7wUf2llgqsyZBTBhBp5G9iGzsvglEKsLpB7oq5i7owj+Q4owltthTy+
IYdvC+2tax6MTvTs2zTSjUb9olNRVLk3frbTp1AC/RxoAdyLpmmtWeK2wrQQo8dU
uzAPEvkUuEYWsJ/vBCHLhZvcGhGJyN9AZWJ6XTli6Z3IcpGEu7fqYivBSumlyrty
TsdxEJrq4MqFwkI63g0gGaKdUy+sZf4FpKsVi+IYiUr/X1KEDbJFxR7UdRKrU1gg
kYXYUaBbjvekCoHlaSr8Em3jYbaD3Ws5pFQ2AHwIShDIZ+XUk7cXJ4Ihg7UmT+2a
6OSVf4T+YSH6Cuip3qpPMPdrR+58IJ5DV05F6GBap5C5HqpcU6dzwvtHUCpx15l+
3RpFRzatWCWzZrJjEkj/jGChfz2WbohM4lnZEFksMCZCndmlO+uhOjgQAbfOnWK9
TcTuZD7//tY/MZ5Xj69GdA5iwXkLeJpMyi2+8FOawZffv2T5xiTQFaaKuErn+7bQ
njXQ7PYC5B6PJ6BW/EGcds9QCt1NLaeSR6hNScbYsQokrGUo9yLXQTe6IBUgCXzN
dT8zLnan2oJGvEo/m4b/0MMR0OS8imruMSk/XEZizl7bqHpXTTC0Zd2J+wK/j3Ib
WY1GNSDivZXuzO8COAzS3Xd7wPqC4q2gXKO02QZSw9I6luXtbnZP0yHsTOG4xsVW
37JJiHOAtm+U/vg+3+ZxTwmKGOZ4rxkX3zjkFNRjKoBoWZfhczI9zc0zrtWAWK6+
5FUePa+y3t0PPz36ZBpsy065OPfOahVfHzStDqZ+kIFQL6aAYjCScUNYV+I0vYP+
hJGL+MbbsWp4/PaPRDUokTJVHMbi43ZSixErVfqwXWYsMQ2Q965rt1NldbYJVNY4
y+GfGBexSJLP+KZ4aNNY9m9axa3FPMw1JApa3gE1micA2WUo03/0wr6st4JvpPp+
q8TZk/LpmAgio/SYDX8vvQZsuvxMawcsDSrOw9DK4rm0o/9U+r3u6CkucVZJdPh2
vyNXrG2MegDNDRI1FXyQYagsz2BFn8g6jrRvSnBbQOqqGSGGPXrGvfyeRV/DO0wT
g8gR1/SfL1YkX0g7Ko2zlJPdyPn13IxiUNx4e5MlCoCU+S+fh0mVEL8utGmMLbsi
MWIx/jeFZ2qJrNRhmOMHW6lDCgXqLl8scFpAeu8PkzAGmMn7gKT7eYIw7oURWNMF
i4yJ7viIT3u2ULXXoXxrv+iyi0xImIfqtXSfpONjgveag/X6rKjCQ2PgBidi3dTS
AT7XNd1T2rFgIq06WIY4Ng5IUiZxNS6ZBdiyIc/hMRfE5hR+u9vli2cjpYAO8UQo
TZasdFG5+KP7vHdYMDmyatNiqzicQr/an8CXDAhxZMW3N0A1O6hiK69fhHLEiACW
W+KMVf5QU4icvFcYDXxY9kDFFY7op5qPuHf0UPtarE7tFR7qF7ZMadNwATsgeaZh
GWNC0n8qQDd25kXgD3BB8pzOR6I65ceJNxHtGDbJLuHP6cEhWODIsIL49nQQgEb1
uPizHVK7RVXQ0deLf+gmC58CWnqu+VRZMPMIGbQEDCmkt7eAcrFsjMepe415pjrs
xlza90S8YGACKR+qNFKVTYher/dIkdgbY6ZgcgRpJTnXtoyOu2YwTrMGzImhafzt
dKx+6HLSSJQniKtdZ5ZJjwPjHwrtMQMubQNlguciHMoBn+p4gdEzxUfYzyP9VDte
8yuEqa+9aYxppj5VE6fWPthNpRs5pXblz2Ak0wNkI8KePNCkTV0f0GPnjIQhgHj1
N7AJbuMG1PvN1G+OI4n696EtYkhnMpEyu969Hmk+JFTSWUETal/qZeIOqnZZfguc
qxu0m6H/G2JnD6GUYluVca2PGrpjfyRrZE6mJZIJXCazTJaZCkSN741dxA7vcNiS
OUg6FncBuu3cRPcXe2InhxO4r27h4q90ckqPLWxP8SgXUGHPbSv+VhJFOgUqBU6x
N3ZMcFtoG+8jw608Ow6F07oeuYbZQW5isdtLGifmsWZEJncZdNma9leCGyw88BtJ
LNVyW7TJDQVJh7efMr1em00l6FDCIu0F9jD8D8Lxot2qYU7+LxmMXf+wMK1pAI+B
RCBHaeFfUla3BJKk25FvBa87hyHOhomIWCep7jcRejreBKSkG4Sg1lPmdcPgYO65
OO2ltrJJctlsGqzl77rS+PXl8KWD4RhDv7ef+AbM95hm5ehrx8pP6L5Pwyq2xaDk
mCTV11C9E0n/iEI88kkeFcAMBPrP4YFTqs0bhfOu0wXiBXcD5G2YfjwRy4vHDlyl
aiPVcKkCEFVbEbhjYqO4gJBs19WBzChMyCP0OqEfTIPI2JlRzeCL2JBX5KQ3U82C
gKoL3bdbB19rFM7WtSsR6//YFN9dkq1WECB28+mpZ9NRoUCmYs50GLrS/Xpu6kls
8vtZqvFnWuBqOLjJnaOWyKPNU/mPI8U6vbgHYjNIYOluC/lex/8nvn3efd7eIFcL
mWYj21AEJ61teVCkV0tW0mnDLs8IBhq8kH/H4sBFYxxB5lVrbpO2XrBJZAtQ12Ln
2zlgaY4y2vtU9fxLyKxfWqWerii7oIm8Z6zCbwaD6LyjTysgG2UQIO3M6zy87Eu4
/Lq3UGwoeM/nTyx+4CyE4zWIpN/KMgbfruDDtb3TFwFyqNg1SWLFq/QADGYp5RMG
+Lf3wZueAMPFeQARUyZxVgEs5hG9gksgguPeDEOjgRtvbE3qZ/HWHEwmNDktTvHg
V4o3B3z0aMHNPlzqMJ0hJEY8ocDtK1bQ4AE4Wgem4t0t2dTd/P/asQzLYl+LMre9
f4Y1ymm5hNOZg9ovM+9lAsEEABB/rPQx9Uol+EAQSEkcvU3i9wgamgnHfK2UVR+q
SOmsdcL5P6YgvYAecY8eLa390fFkIgAtzFc7pIhpIsGHV38MK4kiZrubu+5w2UMA
PxjugyEZqJ/feHaq2MSD263ZU0K3f8JJojhAXSPyM8Zc5gmTcNNcjtYiqjL/b+dh
Z7xFSTXTjRy+G/ZGdDiry/ufa0OU2Ras5irnsPdgXh+2sZbVICoK7QT8nxOIxEA7
CRQGkXeyNejAuVKqQjvopWwNrG3gIHYJmfnu+7W4ePz0B13rmwtE45zgWQ5mUygJ
0GD1up1Igy5Vvi79FDNISrU+yGY6GY4t/xJHvWxRGyw6xsSYG0Q6zL4RAGbd4u7w
HmXwAXavfI4xvl0FbeB3VrLIQ1n3rBNLSZpHu/XMYUts2H/FpWKxmOGmInKl2rzY
ysFF/26WJebzCeHvFaxwTju6ZQRVUCOlQ/nZvEO/aV/Q85N8UQoETRAC1Fija6eh
SYTIViPs+lTtV5g5orlWbH44ij93f1wEZcedeRHOSQ7X/wgrrVficvXypkGs58cG
oOOlhGWOn5v3PAt++pDKjeWM4C2V89pBIZIv/+rvJrlU32HaS0ZOlu0jYyVhwRpK
1xQy4IFT2lB1pmNgLW0eDqrLG++19nioNwrq5rQHvqcvAuB8Hqi+yCdb4tfo3hsL
M1CDHQfGdNSn3udxgOll2Ms/v0VAB9+0et6IDNrOrWHAadmtvm5rinYvWRB3kUmA
cq78N17z806I+sd3SIWAVxR+SkLYZNCI+LJz2GQUOwZcA3FHUH/ZK+icphHmMVAL
OD1SsVY6hcp3IHzEE9+3GvfuP1lGHbs3Mc/wqOiShLeE2q0ZKUMgu8Acgg2zahUF
B0/o+z3l4wmzskE9GLGeM7s+FtWvrXEEB7sstbXw+Bh0S2VqxAW3AVaal6wX4x4g
+wkzulv1gx3GtKY0+FLMucTpBlRndgXqY4rwT7GnFxPEr044uHS9ub+VqwkerKEc
N/lhZiNosgL4xPumjXNaciN4JuutDakNSjMjeIfeKgUmJLZ6KopBzm2ov8Z61H+u
I0/kuFIep0j5WHeZRVNPv2WK1WPYF+VEo0UmfPzTAqvvMQPit10q11JpKkG1KESk
8Qk5PeNa/NOxe3H1WkpKjgVOk28n/h7ysXr/Lc6cThCu2f06LHuWg1DbGtjnjgO/
Z8mZt0Nf5vd3+aGk+Mm5aAme0Cz2EcQGHV6a8sPm6QgJC71zcSpk0buf3V5v2H1Y
NQci+FH1xfTs52CwBsH9AY9McmFRC5YmKLYmylBVg6m0kerUv81zfE/QAiCKuGo5
MR/AE6OIMiivcz/qGx0LvFOgnkCP1I/XjOvuOgPscXORO9cA7OqkocNaBqteUgnc
s2nKR4gF3ZTxwovQTn/PK7lGGh2sLyzmG3knPvTsn4XdrKL6ee5DXv/40XTYC589
S0UEB72H3ELbm560bDGn6l+eMEtKWpO2BLPNaJ47DeWkLNfW2y5Nl0D7vLXDU6C0
myUJJCqNMQQawrTGgJ/pSoYxQwTUjpnLsELRqNemitLj+RHEkGc+RBKs1ViUf37U
gphgQgOs/qB24Qd4EG+G18uJs5Wv+Z78dN1Qc9Btuuf0wbmZgy41HWa6NM3zY5Jo
yxCsH4d9cC9CCdn5OkCz3UyEqYlDNeoWCkuqvmIV1L8T6vLIo2zbENYA1kM++vba
xse360ScDAdXDmNy/OMnvvAZt98ZZdAM4QcPcxnGgt0yr3XhPeQD5G2cjz8XmxXm
tPrRuQZbIDH73h1lOBi1tqJdZY+aa+yhlqesQ6T6dVXDaeSvJvgvAOWQuz8BcWq5
yo7Spjh3cgmnIbW+v3jtpHkYfmOFZRKCo+dCH5SVBqo1IxG+f3vpeTJDHh/0oKg5
3sixzoSUDeKH70yO2TjoROvQknMT7LAQ+clOtuwcUy/NJ6MCXUWfpceR4IWYksZ/
ZoRrW0zjBCc6OIMAkRd/VG58t+npJlDPl7GuATsA05K4IhOlkkDW2MzmOWorRuqr
AujgRKukXWt7GKZSKTM/gIhVzz9mSpieGeo23pEVPIB8aMBrVdHgFnUt6LJJLbvQ
a68U7WMh1+V01WJaeSJsTw+v0cZ7sdFy3C+QSdzt0MctbaHSag244FYki+5VVOdJ
r3MNFn+XxAP422s+2VnRYasWFmi91sCXWbYWqXHv+bLaizrq+n/GWBJuna0pC8ke
lqLt70WPYp7WQogpfCgsmCFrZBZqz6scasw2QH1Iil2eNlrpQ4wa0EOGCBJg3ZKw
8upVgDNfwfPIHlUKjx8gHq5et4bdD81IbnjerYlFQ7SugRmTFxbg76/SU0Ev+whB
ZDqr/Sw6C0QVhptU9BOsCb/edilBua78DhXMlNqgvXp8W9HJ/gQlbpIlZ+68+5qA
aGgIEvBTweEBdqQNZkwZLzVFuAPHDbTSFoCbUUtMS+ZKyaLMuJ1BscTgGovDbdna
gf0G8YtC6m7+sHJLK3kwG9ED2eyP4fYmRdwICmIwWL+7GM8bGJ5LUTpTKkPyDgji
nZ3+lpvmdRfAwHFfN6EBTeDCg12JjQJdAgG6RVLS4OMcHKe6Gk1cx+9oVJPL3cY1
+LbmWNmPpk9fsTBLnwpMQup48zNDucWbywMoeWtlz6GChWi5M7wji7xGhz0EV11i
rNhatfJQH+nabE4poO9RLiM88NyQvgRej+fmQlu2UrYZ79yuD+TTZwqNtT27H4Db
ZWYak/f1j6CM6ZFln81tTqOfHgpE/jLQjyLYffK0NrH0J/YTkQ4cjJYyERzDEYCv
gxVlWuu6E1mBlW0oxALkITyfOf3EtzgZpVTtx4RuLs2OfvmSnuz+ETmbUvzbC5y3
qdYGAe8K7tErc94mRUvqTkF7n5lL/JNO6d3eUp7sA5D9QEOmA+JxNrpWrvXyRTFT
221ZccRS/sQeoLNkDTXOmXuGVGKSdZ/t+pYoyEsrZuSP63GSVLYhY25usg2arkjE
HZI/ptBFILmtkYK4Ex7Lo9AUpYVUZp2SlEH02UZwQBH0Iwf96yXpuHXoym4KAs07
MlhxL/UOqbJVsQfx+r/osTX4z1zNj/wk6TVPNSW0IWQ7IM3sAAFegii8z1NzzxwT
rlGftCmxwgvBrnp8hIC6lV0fsSxDbuFb1y6Z8+DLvrdKWzKSFBWq4sFnBrYnuWAc
83EdtcIhY1EECg7KbmDaBN13PZ3reckvR1q5cW9Bn/92/4sl3Ysjtu7dxsDh8l7s
SQsos74ntRk2nIiC5h/QmnwoKJs+ctiCHrCLEaViJlOqnXto4gE93esduZVi3Qdt
oA5crGc3YrAIl1we9jJjqHw8qYegODkXAn6I0ZczuIBIzlE1DRLHsiJNbCb8VCwA
wf0fWv0Xf+DBwHcBEgasLComJOxeRAPtakOoRqsKGsq+XdF9wiSZeuvUpsJp2gti
OEUGFWGBm3/6Zv+6e8XD1OaRoLle/eU7rNCeU2k2g6AEZfqyZrKkuWWtsEXNPew1
V3YVbWsG6ywY/Bj0TCmmg6BHCTUWTIMQSh/V1siG61uQHJNGr24RhPTFyz9z+5Kj
5zx+MC+d+u5DR7wgXI1x3T39B+WdsB0cXkpEFvCoHb+HhT+Oavlq5q75i/3HRIth
3V9fX+ptEOMGcEjB61MuzwkJTLabzsV6sX3XJao3oTeeJ9DSYIXfth1WSGWD5gyy
9zBCxN/AfkpIovBIVmVgGIEGhCfnGwiLucYVG1/cTx4KrBPkmXCxlNeR2IW2pXjz
2Sju3SSaNWE1fKZ6s/+CEYSmedH2GyzrJSz3NxDYmHulOGGKktzqOXSH5MUsb9jM
ocOPdUKlFdVNKxpJcXm9I0q+tp0pAGcKNYIadUrNh9BTRl7xEgOOQPEba4qnFmG8
0luDo/6zof9W2qJMw+qz5q6ikwBYwsYezYE0JIsURmTO+DSNWCetHIROD+KBgg8/
Fl/4SX/dxKVTBXuaZt6HABbzHmC9jNo224rWdsZAAk2sR0VHKHgvzsEFf+spmUFt
jJuZAUB28fwEuHzdzYcWvRwJ9/f+8peXxhO+Ri+rDGjLfBBhb4wkwnQeakIaAsAN
JES0S7kdakCDl1xxTAnqiPWwG4LhA+iHxWR1ruUn9oTUg1EMv+RvCFVoMmo4hRso
B5alit9O+GOjvbcimEvdHLqVzKlSR9KtvYeNMAxSlr6JRCg1ZoQHs4i9aLCZb+UL
zUuNnGUQZM8EyUPEp+Gt1JdPjxRvljAPBrtVU+GzFTVazeZmSTIB9/7yGRyjNUKH
kt0+l/xPHPj8ucYmGm2TEhptkNGDzZVwWBExIn9Guve5O5lDO64E/nRq0IxZN+Z8
1wIpt4vwLoDuqr1D+srmKp/JTIQd7Djvjsc70WNEQ3FE8OeLZZNRV/fXOJq3uRv/
5gZhz+ivKgBYih+DxvnrtYFJnp3W0snVdya+nT2dwfd36YHahPClZ9WnKz9HsJTg
dI7iRBJ7/0XJz5lvgAourjmRK4xUDL9oMggO+bla0lSmFZm4cuJ2mfZYdqOXG4kC
eH8glcWdWyJ4jIwvN6Sz8Q8CtIlHRtg1ULsBcRzZV4qOHHLOusHaQW/v7kAgRKx9
S36/F1hc1/SCh4VUnrNM14DDLlNF0ItJ2kSlWSNmIaLPxfFcrS6iwYth4Dc3FXIn
NybzEH/Y4RUypS893XpXhB+DoBOocDATcT0A4pKvQxF0SZDKvLl27oysZUd/4shs
4nVkxYp6Q9yVnFZPHfD9e+Im3cOH1gatoIJfJwIjske8RhE8KljddnhI/hTlKIFj
uyaHWyAgJsrKa36jM9fIkRC0ZeK6G34GonGolK3lX8l/mhkMZz0oDGValMDnMIFZ
hlHBC9NM/iq3H7+ZLnspxXM2gVppeZoLdTIkeTVKfY2MIf4r0CwAylUHfipZGvn/
REN6b5gtP7La0wF9CMv8Bol1n4FY9EdCPi2fs1+CmGTOo7/sog6HGNsNnSFl6Qd6
FTL4kS2wAmOPg3ItA2sM5EO/TIAwAzEwXeh7iDQDcteyg3Fj39vWwFd6M7OE6fIK
zHa0z8QOlA91skud8RtU7mIWv4J8F4+U5hfURv/1BNtZDxUNI+z3dUNlOmo9VK7l
yMARZ5vkV+tOKeVeRPVYSW/YvE57zekpKE+m59w5PE06MxX44FoSsWv5bPEduncB
5V/pcYaQBM6nPGTcGK9c8M4d01Xl2ubSpSf8/KB79Rn07LX0EkYUC6BvujGpLytK
ehiDH14hNVouRP0pCgBSZ3Q/D/MZm38RpmBI/kzXnzmmdfBXjwDrPENmXhCgv8h6
8JR2Hjp6TrglgF9Hk60LOUQ2LOqWcwW5Bx6BKo2jnZW6mdy4nJlSN5gnIsjpJz7J
MM+bQW43bLLzVi78kHVbYw70pp6a/2oery2bx2Zz7lGwPoTn8oh4RLFU7FgVojlF
VzFikZxMKwjsEuXRss46PF1Q10jqg3xoc0Mc7Jyap+NoaVprfebGg21vNaO7Z9o8
KPPWYNmFAedb4BVndV3JGrd4BJpHpXoR/GnewdqH/zVRDFBFpHCvOp+xJrlWNwoT
/mqITY+V8+BRKtbxqct3ppOWo/OusgYCX5ZaNcCVncT9WOcQLc7zAtrTa3GT6vk2
MfIfk2UE9khNBkY1LbFp0K0+Pgv9PkEicftPOC+ZDvpI7ivwSwVJKhFalcS9of78
0ZO8IvEFVqC2qtoFU9XCr+JUsJI6fV1wagB28bx6wMYORRybuV25fJMv9/Da68BN
akKN6Sf3DHiTvTz7kwi7N1l1jIATN2HarvlJYURkF6b+1T/m45xDa4yhXJuau/Cf
uFpZIkYyg3W2tUAgvCbiosVnU5snvJ9yADYkp51x93Sxdq9Pcd3nZVZsWh/QSHGl
ESbh89BXLh6UZ6WT4fxUSEvOx+qbh+wBajrXto1SbONz2bUTAY22BX55czCZ6U6e
UJy5jPK/+RAbGbsh2k8siRgU3VeXa2lxCggEBxRJthYPEVy5RUX0Lrkc8dZAYjsk
P1atiynl+FLrOjJVXV6t8f0NFH7Tqmrpbjv3y14fzVdyjlk/zc1nF03jwnk8t1sx
PuHCgUgxjOjkJw1XuW2pYCDg8o2ZGfdaDi5y6UqpjC574QL2Djc+9Q9ayhMcm8p0
nPU0qwtMPbBSqLQB4IhlXtGV6gKVEIxKV4ZUPzLXE2oaTpj8Xt/ny726ILC0yI1B
kGMXTrvgyYRYArL0DbdCryj7C2HZFgIKvVwoMtsG8fQwglBFO+2b9GILNcONXAyU
pcieGUkl1yO8zO+PbGgvTL5VOLli0Y3IH7LLgWlJs+inJffdCQQ/1h96suVXJJ8H
SDyo3jpTZAd0fJ6dkuwIoQrpsdKqRAPc14EXfyofZVUiquM6f9T4eV2vEsJa4DDy
1dFEOEV3upV6T03jU1jTlg2OQZdPI8ghBrYnvYkzXbFuvIi/vVU5iAaVH2nsYbJ7
JmBRsa41bMMZ/CTNmOjUEgJzhki6JRZ4KTDrYeh6Ygf+F8yP804MBKYae0WRvP4C
6PKGyuR7JEYLn3h2JGpkrUDrFo3qOBqgx533YGXI4G3Z2dg5CACNmAJlXRpae2Db
ZY7GfUChupPLYCk+4eTrYqOXhLZ0XMvUlFYoDa1P4f2ALmEOq68aC5UF/HGp17Ce
MUoC3+KkQSjNMMdcoSc4WwL5m2z6U6uwmwasdcdz6xFQ8gCamycPTy4/33JDzQ7h
w1DTGMlJsI3j+0z7ySHqwPuJiuFBclreXuFnc50GWJDsPNocB9zgMo+2foqYqsO4
8LV6S7Z8RGrzmcFGTx+nVrALzV6lyDYSGVqKL5xPJEwL376miR5eojzAlp/5vmYT
+/pJInRbfBsTqcWxnut9T2mCup8Ou47g0SW6uhqiyLEOTDInu5B2QFoux2ew01+Y
l7djEsl9unZo/iAvsJUDa01QMMaOMTQGnnL2vs3lOy6hUT2E/hPxf60t17EgYXdE
4f3kdZt9i7X8RLjTmNW5kF2thtICjyt22eKYNrACi6PjGHQWGjTuD11ndMTV20Ef
7/FbkSwjqMay/Iu+sgxJshvs8sDe+UytDhPb3AGKV7M8CIYUE3wq5T91JmBGJAHi
Ssypq6jbxv8uF0BFlS6N8BSCzzFSm/0GPanWpMSYi1xgD93Dcb+N1iRO/t3GvXBO
ZxrxhZlt8LSXOVP6fC6JJptiZLbhmLcKOetCUdBIhHw3ixyyB5Mf5cKujUGTzN5/
wexppX0zvCFbTup0st1innyYbQvJlxQpqdgSZ+11d3G6sUO1bdRIy/IBus3+6dde
KzIvdsO4uqqWY7axU7ljq7s2KcYZKYMtUToXD8ac5bJCt8WAC2OhuAl+l94tlmfb
OlOEr2yD/xnToDbSSu/Ec7eHjEoyW+w3OEsCc2DtbnSTZ67EeG22UGqRW28URTFR
2yzQTVO5zXWGxV+MECO/+jItiAE4DAih3bQzn1CgqdnOjzsOtLMUJ/zKtqVj2J75
dMABWhx7+o2dT56FludEJi6AOWy8AezKS/HXFa4hkYewaXSIgR3GfQYSgVggob3l
wG9rLdfspBM585YP5e0CCDu3upyTloOu3vkRNVrG65eeVnBZ8De5+YUctlNYMmN/
YBtRU8Pm9g+Ugwb8h2qzYztTJcNXI/sf0yMWSie9liyK0gHFQSVzOMj9lGhXgbPm
/jpToRa1rfSuIAo/fuTqdFO+ydo13eKUCEHhXioFIzhizBSpgJ9Hu8GLHDwPRhcZ
zZpJXa/RRwa1rZynP1i6NNOuiFFmVhuTNoi5eu03kklxeRz0OUk8XMa4QDY0ROYV
1Xoy0NEdGxHuPneUvINzRe4PpOFJ17n8bY89B9qpWZdud4KHMozMdU6lB2gQZTqw
6qrb9QwJwXOIcRgOckI4sWw438y3c+PBjnsUYT+aBEaAP46AlaZKiCRc+ii/MSsZ
ARY1jWXjKQhrdwaTssW01mcfZPw0RATMW7iRs6uIaKpDXMaFbZQGPrFWypeiMzWt
KJXlbh+AbNYv7wTXfCoH6ef4CrjsORnS83dk9Xt6NI+aGWgFywvDo+q30VnmkO8y
Vcq655htjAh9uG3hrr1e0HFRFmD3TbJLPtUIjKpIak0GziEFlQOVbQiKhcHTaVLk
xnvJO8ihBOB6mQ3NlMVjC/xL3IaC03rW5M9lIkYo7H4EFTnb65HWPAO/uEytyr7t
IYlnmJd3wuNvK6VjHJYWryixByNl2w3i5Kf88UB61k5mx6IzpvqTTXqET8fs12lO
ug1edOP6TPImjyLVjMR9XRuS2zdamfyL6JLKw2iCyhSVrO9yt/YAzcqrW3oTTAVY
WUSSAOlQDVZvafBumnoaE8vetMyBqdmD2Gs7UPmfCADRxC+nn28HNNGNaVxZ6HC5
O+tc4KCcR3OOoptW+rds95l5YBhaO4ZPtkmpJtAGv4NbSNAnPsEB7Tg0pUZJWyk8
ggj7PCWhWebSMWS3QEwJq3x9kqCsb7+48GbnTAd5r5vW+/SBPsD4FSRH9TQVn9IX
rSjokPjCd2sqcKBpKPYgG4T5iiue4R5Vz4g4wzaow/CsQ1pQCXTahMBp2TXIA32e
e8u0fN2fR6LsGaeIvSzaNzyLxalR/RUJmfaVOdjBjYmU1Lh0wY8YsDbo0piKlwiX
aPJ/Z8HTuK61rFgRVswfyfoCel5rvfva27Xe+kgFhZ5S+iLBwrbScRdXiTqhKx/T
KCBeh7fpm/fCNGhIs5FPnu+v+JpnRfxuoM/8wQwGmWGErVxEqR4kVvOJTWRIZVdS
Tl1aWD0xFcegFzInop0XfMrl3mZA1ISY7byrVP0BgkvWwN35G494X/zNURUkraPF
2fZmMxyg5PGojO5cU0Xr9ilIbyZH8FP+JLfuq2bJ6bfl9yTskGJyT6W8dyufmpls
95djV1xZqt5ar7UBwmZYLKLha9SENcUuFqLWd5evibuJydfpSJ0ywVV9p2YyKAqz
PYC0r/4reOeHbiA4gM8rVnNMev2bP1dTh3+4UB3I8Cm+7RdWnejiEoz5jw8rEzmj
WB8HLZyedIG1VoapvGD4GkJ/oy7uMSbXxFlFQ7kRJhiLkd1Tj6YtuSdkdhLH6r8G
pvQQR1lLxYO8/IItSj9uktOLhfdxIBqdK0jRvzYWPn2GaazpeOqGCAyXKd1AvJkM
KyDIYwBLVIWoaSKhcdTX0L9koZQVVee785ZeeR8X7xjJgmCCIx/gdkZNldHXnSjZ
hG9rAHPgA3xb9yaDmoVGdyb/mBt5Rhs5x+KgBcYsH+QvZk3afqwlMFCXvvbPBTLT
C68w9a67mdxjXlQm39we7M33ylb9DGMjJWN6wNDjARgjcrnjm/oLq4zKDtkeUk5T
ZLX0rFyol19hOMJ0/7hDxBte9ojVtqY1w7oBS8u94/5SMGpjQ1yy8aHaxtrH3ieJ
J2Oe+FJigkTqthxSfgSTn8lISaTx8BzCpp6kxCyRe/MtkYUyqhG/eY7GUKzD6uWJ
JeluYtfM3En4tQQweWeYFGlwRZiR7epjhbID0vsB+Jw+6g16wfScxZDIjaglvzHi
EfK8yfslqHCCYovTptmRt15XJv4rRSVFdO8UK+wNaOPynUFhWhNWdBR/m+P+lcsV
DdUXbQs89ejpiz/GyJoYbt2amKHm8NFYD3qnGoubYG4NYL/H302UFyl/rGb0upZV
JuWLmD3g7CnMvfox9ZU1ETKghP6wkhKFGfac4mOlu/VYTR0K/kYLcudePdCsqphe
5muPRV5YRP8dXyTxU92tUXdpgfIDXqZUZE51vauQrAK6MeABFwICFrTuaPLTIyeI
cOvwm+QaQ7e8GJq1apaaRo/Mv/5kroBikHRM1EvvDGllAwirc7IOir6MFdMwA4xm
znUp0BOkzs6dhw113kmWyagKSeL+x4STG7xLs/itKDKxVQbVG8iivwllP3/UFEGY
84D5zXLfwSuRREg+jR/NnKBlscAZhrT36AjUX/dpAhta2ZVZh4+A7guUlGeLP7WQ
IxPXj1XfHrQhn4Gm8xzuWHbpQicOr0+7oGbtoRN4Ic9KC+dk97GcoH4Mrs3m4vIt
nVzvFNhMxIbaBYd034N9kYxY/6iKDIcNpnXhYIauPTBSbkWXteONrKeUqxY4Y6sj
RaHF/VWXSn+BHvDiHXULFtNGEahiJKCjEBG3vZvPCknviLlueCmKII8IrbV7fQhW
Ws59rv7OPCKrTOy+hp9Q5l+CIyrBzWFvtiE3HHhopQjpB+vGaNSBSXO7QOPn39EF
Ns0Y11o3Dtayw8jsuAh9PyrEY/NUk7vGbNWWwm8DSOew8wcBj9NLmBsXNkV/qCsN
29GFLz2ZXsiiSI/+TcvnFakb3Mwj2TeOOnhiz7PBLDS4FTk2vxrMmWPFmzNKuQX8
LYaw1/qhz5jFbc+uztCkWeXtoSxMUktIUHYwa5zcTDCJjDCUD8x4h5pajQA5x5mR
dPTGBONs4rTN+LK13R1Omt7JNAe0W+zIdQsHJ7MEOGM3KwJiATqgjlsuy2Vq2DZT
N/RXo1hL/K74gAZFZerdPBxBpgSWNU6SXtDbpUfymdymYMANS7nqu/9IKwkV7IvV
zYPjrb1STyypHNGglvhJXddnOIyWKp+E+8PNva/63QqeoTDsuA/OLalMgq44Rxr/
775ac+aeX5HqyzNfX6diR0H3z8aCIMPr0TSK8+v1uWO17HwSIrmxFkwQ2qKIzAWN
NbTk2IS1zPxV49JozUeqUcMlPb+Kx5VgfWgPs/QXm6FJ8866UdyqbAE5zE7DpbTh
eMROgKvX/Ztsz/oNIvshzqV3hv9K6nofwAGHfZhHYe0zMO39r4Z4CllADIarbOPq
p4Dqz7pRiyXmZNpnnMfWCuIvJoRM1BI8JBryLMEe/Kzh4OY9InRlUJNqgzDUAbGU
O7Zk3Ni5eaf/mRZEndqLOSiCiwAl8yHmhjXvW4hRY/Ayu+ptgwLTCL6KamhCOhNH
NsQY9Yob2Y1hY866YtaUwvouPcQTXqgZN8jNEmHsqumozJPbqkSXF6Z+dy6NNtot
RPUXQmgYbf+LR1pVxGW0/vC9/96iQ8sAEaHSxvLsTkdZedVgSfYd7mGXvNqoa9Bo
1X0OfNtYEZlfMs50mO1qvq4kqjiVGG1BM9K6qQX/10SNo+ZAFgPSHG7oWwusE5UE
Kp+zvXPGSyttPuuEsMAdDwYPh20dq/BsSD6J6pWD8T4GoEcWEu8rzFOzbuP9wFgT
zF1/h5N6VF/bHR6TdWY8H/o+Y6TofmZSSW6XD95+CEcAQHDdvGcPk0AoOXWsFa9j
fvBuA4gYWAoT1jGonEBONt0l4NACZhH/0o7g6ZYVzCWIkGCxtbPkv5OXyU6XR8iq
8NPO1pe4Pm7x8ChBXS8UivnT9RbjyyMcERZJC+2DXOj0DhTSMl+VFOut1VIECbRm
RqhZYH6CkDuh2ZOik5cRYw09QtcBmRDenUstYSellrD9UdtOicovIYN4yS8eEe9d
P5180XMEIynww6ybybfeLakUq64GRwSYf+YlS183dHC7PlFI3ylkOJ/qk+rBc/PW
aV9AviUJeKll50nxqTfBCMz2ph1kjJlSrOYLMmDvFRQBr3ZAugEwIvIYGzDocgCk
Zb748xwGbQRCCAWd5oVAb7v2osJTdlCpgMEEtBjJmbEMLBF98WajJOsjvj8Gci1J
2ru41A7+ISOz0qxX5IaLTiDpIpVeIty6DIAh3C/pNZv6jQjoZK907KcxYE6XfEEc
amd011bKTUO0KVr9nP/9m+6LVx2iSNyy2IYjVCtuFjgFCRGFlD3iHEuLddC6S6Bj
9272NIJGVKXp6dbFn3b22e12fP5TA/oTcawtzb3MQM2g9wlB571zJqO+GJmCtGNA
kz2+K07X/mLssn2AIgNSYR86BNfBun+bbiRLeNCBOImNIEMYCwsz7WHDxjBu2f86
w5FNrj4n8FXDtXcCJu7rEnKYrQuei4jtlxLCgkEuKQlQby8bykNjb7D7I0OaA+hM
JW1TOVEgqPRzFlUyRNUv056DhfKesQZjVIwdVpBi/6q8dpJQzewnoj77EdpMZJiE
/kzKug5cKesskH+6egKnBiPFfVbaoyZ0/U8Gtv/zN/z3krOM5PzkEGNLLiIgls2a
OlH4AjP8XZJDi6DrUiFKSRJ0ey/h2JeqntihnvQWANvIl7SYpw8g6xGDDreMoevr
pNFruQ2Nxpb3KcSnXaniM5jfuQOKRuxNaDSqHH4+8ORwW6c5cLvhuJwGkKoEOuwz
+4hOnXNkks5kpd4rHfj9AHmHzcdsDQV63k1w9AGqyy7h2X4w9ruzogL8xnnzQTK2
AjnQgSOVEGdaMjnxdPLR7cbsb7UM4jiwAZMDUf2vbjdG7YFbNgFYsRO+4OrBVEW0
BhzbBzWVeNkQLoD4MPxNnTYzGSw1piYmOEbyTlvfge7RB+YYJYV5VzsdzR7Vwllj
Xhe5P4x33flQxcJRgQKOXsXsNZvdUJlf0dmbaPJ6zOxfMMF1oGJ3XIk9WU3gA1/V
R4cI5ULwRQ91shqkVt6BtvuhoQQ7awKBX9FLj9LnG/F4m9qENK7qyQhik8Oo06Zp
1CduH1YuqfmV2Whj0FcVREGfWBnT5VCpd5xY7oo6AePmKj6+G6VuUqbXzHNebREU
+3tcic82yfr8AjYINKPep4Uxz9fwKHSJ9/z0ycGLnlexSfciRQJuSL3EIJEVxRjS
gT9lzaI+7BxuALflf5dwi0cmCpAV4e3zzQd8Ealf74iIvdlGS+/L51Y2LonRn1F9
iiUHiXTTC7Gi/HFryfcwUapleMdyhlOxQBMq9uhRHQDVLgcDMW0QxP6fb5rbpRDG
UZoP1nRdMzCIIhSQpFT/mj0MozqR+CZc86JJ9SzguSvJilVdUpfdOhbdpBEcgW3U
rCYe7gxArJKSmz0iRS/8slbv61dXFJNtRsKtFXxpiANFEquNRBOI9cVd4s04C7mx
E2D2zntkUPQg/HahFOY1nOIWo/rEkz7q8M6lb9qTLATzaSqEMSFDYy2Vkw/oXC+W
zeC9O0JfEVgKxtYKZ+azJroyDZriAezK8f3HaMDcZ5URGxS+h++6S+J+loWP61YU
w4KPCXoONMsgm5h/pqJHNi1SeWeNvMYT+wbk4itK0+TKFNMkAYNBJo9J1aA1xE8j
BXVb8yWMWoLtKhDJXCEDMLsdedex2IY5Rh8FcZGP6020qJhVToL9lYtlADIRFPkl
F8u7kuISN9/fgFk9VyOA8KO0euaS6iK0m/Y4LCwDeGavwPo2uHk+izV68ChTkhmq
ljAez/A9/oyb2LhyXc/Wj5ojErHUMLDIoGgyh0RDBEWIPpfuEIc/Y+c87dkJpofG
22Ts52im+IaMkHbP1K7jfa17elM1vLbsmT9i1k1wzSg91i/49TYZGViAoBRDWRdx
aEgjRUukY+HWYoeMw7N17xojwanhRBCfYzFfHKZkaAvLwrEhlvQLeg+PtujSBP9N
azH+sgCI94BP3Nmliy/Jf8BChnTcSvBmKXCvWMAo6929j47nqHQVnVNf+JOj8To/
RIwo9t4ZwCX6TqdHqaKh1npwA4CTRlKY2U3JuSdLJAL1Qj4tMfAPHg+bqZ27/b4l
JVbUt0cCvFuPfmv67130ryy6v5S7reY40HgTfI1wottuR5Snwzb6Sbyc0j6Wq2nq
uqwBpkJcyKSxduAZ8PjgbF9DQr+fdm39Pqm3MJAHnrBGr4sj3d2SMJqLHsSryNtl
DIi5dksbfQdpvDWSCR9VpyQ9QUqQN/D4skYtZIsqhcxIu2ykpz+dnghXjAu55B72
ptvZU9V9HmxZwmdFGOEBNGW6GSBHBJb+wyRRy5HRi0sXRDsguCKqqFS5kA8XqAtg
RHFSaEYZGyW7geaSrTHJtbrxp3/lamaueFtzqmpYIwkwsMD4S6VaxDrjvVzR7rL6
tv/7xmWeZDsdq7WNUWDqahe3VbppggsNf1RF6ADbQlgsAO1e80fIzIEixPdEgCd6
m7clms40XNHjg0yqrfJ9xiv3Dhk1mm+m7KrdjV32IopSXuzCPSnr7n/Ot25KBbxC
kAvoKZeVKGlb/Q4AKL8RVwv0R1SHRElsUDET1hLjqO4VkLZv1GR8V7+SUpPVONQs
MNY+BVz3PUIvhu2UppzwvjqzMyJHglnepKSbNMrpKGgvG5sLmSaS757O0YV6jOy0
vhLlSflqiYaVBaX2jWnc8L9RjCO85fjh7AMWCwYvny0uboLDJ6X/swghoEyBpyRR
rW4o70/MUMhNKpEjYi6v2xAkvFbUk9UDNhduAozzNDwN5s+ZVCf0/pi5+QhyOOxS
ES3fW8pJi6llWUWQYe6ESBMkAhfqxsjMNQ12PX67Q6QKSEweyTvBgc6zD8eLEfqt
q3Z+vaUmfDwNgbgqJyJLJls8Z5NJGWlai/E9LfnzyxDiESjY+FfqINTpwjU8+1Dk
iD7uN39PFeqi1MUwc+dbXP2uh7FEaTRy0t2Zjj0MVrVnlLfDX35Byau88tcNRoCm
UpISUdZoYgn/vYBigDzfmflr/LqNCinDUE/2T0VafhM0W7ud7uEdr3Q7maEfsa8Z
qtNFfX453pDFCIz5FUOFywZx2XS6EGBbZTnQYfq8cU4D2kHTXdblrd3ngM2X4lk/
LETRd3ylOJH60ZS6Tlzg4no+IoiaATFJKOApE9B/LTyxPhe6NKMLiMIIMZuViRDQ
2NlB8wA0mkujOuHjon8QlhesgWbdKLbxzUblVX4DGWDqW/1McjGUoQ9BG7BwfoQz
0lTezHoY2PjDw5fel0lXAgfJXe10TW0XUPLsRh0Nisq8ekIOiCnepO1D8AGfcwfc
UeFswfedbTwXjXU4UDDUChs1zIm/wuC/rYF0u4pgIFYsoqjx3kQMUypUC+imUzsa
N7aMJJSLX2qTBR44MKkVCFt09fYg1tXFbp6+M4IbVGk7y7hgqSnZovlc6+yHhTMt
M2fuWtVOyDYoqY3/NcwL8iz8gtK1cE4gh6gPMzJQqPnXfY/IaaDWwQfvyKqruA0M
3rReAFe2h58FPeG84H6XYCaCSfUF3NtNWdng+PN0gCVZ0uoLdS/bSAN/Hsxc9sIY
2iThp+BP9CZYroFEOMLAUUooE5Xs5B9QEbHejdsVsfsReSj/F1nxbb+xS/RpADr5
/iT7P0S5YIxIyI5nlkrmrvkO947cwWYK3XabWtJVaGKyu1pH48JOMLunFuCEncud
bv9jDah/U73IOV2YVYNzdiDCy0P2oBz89gUJoe3G3q1LEZGkR+/QhZgGA+TEIDt3
//QHmNV7fduD49IDycto2+4UbLBA4uZzQGYAHNwKj+PZeMhl0eqdUXDi2z7EX9lb
PVis/uud897HBq2UQmQ7gDcOp1MECxMkalywt9xtr+TUKC6uJtWsXvdcWz7L2ZtZ
z29natK1JGfars+R28CaGQUhSEEblOY7l3OBxYELhO8YP+rdvJMg/Clm/mbUHwX6
lktt2YlPgXcymx/YTZR7LDq58qJd9fAgeqCATozn8OIWF5OLOK47xGNyy2A+7GFS
c1L03e+6kFMugZpP43EBpZQsPeB9iDRizvT8adNn9fofqtdgMWIyQb+m0GXG+mDg
XZdv7bpB30QrNRiuBXz96isqNWdn0+J8X1dNXDGOt+UmEyRgBbmAIm9CzE13gH+o
18xDCZv+ILHj/kAtC0wJrF/zoOSoRKl559nb5rBo301rqW4Cx8nqZ2nzAyX4zIF/
cvX7i1ku9/I3DomjP+gmDVPysOcEIGBse8pwZEh4Hbwj/2WRb9OYzMLs9lQZ1urE
O+1dRW8EG+MD4ghTso/51sgY6OBVPsVa/GZlSJqcxRO6WXUdaJxj6evIhqVcTw5B
7xFDWFfUHyfzPg84rCRYJp9GJVTnQpgr7Z8Hkw3EFgAYSNC668R6ajpDOI6VWPwM
5rHAwQzG7iU9NS4tC/ZIses+igdDpqyhsXMnADyKLnISAGGnYMCk9PXz/P3p0Nqh
TMsGfSGwjQ9Od6LJIdh0TsWvfYz1MsBCY5ju1KN2tDH8mCYXVJH3c60JVF3dLiTF
BgMjOqxCFdukL9oLYnlaAIuiSPxZ6SJgGqi2nBL2hZUknfsyZBAwXIOyDMe6Xk0R
8Xvlb9C9yZvlV6T71b0F2UrduTXPPxI8IBPH1Q/TwS3NAq7Q/QQtbM5Luud0tRE8
ITPljCbjnXfgJYBn4nBEZ9XYRvJJ5/ZbPJMUeEsgqtyfoAOM7JvkJP4n6GRWQmj1
/g+LycA9yOki0BctWzj/OPvv4DGxqrXVWfkiSwWnMHDW/gG/9TtvaqADgyoxedgT
kMdpfCMiM8VIoITBBnXwyN7IRqK02ZZBoadv8waHE5KnEgGPNhPjV6IuIHbmVpRk
MVZ+fx4dTO+P5wRDt7ee7yUIo6Ml+V0mmijdtDCLWaMYZyd98OvzE+XLzMMayJp3
ArPUzI+oxEGg0c0v8DXd2dyVhF8ndRXwGqjl8uS6FtATJBXS/1xPo01drW4UqKDh
5VBlyZW+tON/ivnAsmHozKOq0w4uDtelPhh+aZdvf6CfiAY8iF+hEsXRRaAzrqZG
XOhoevGKUrnG3qXhFBIsdAF5K31jCVnu3XLI/VZ9TE3zjuzx9x15d5X5SgEQo1Up
osOmkmwgvwFDDWGE2tAMrttdAe0F8/pDYXxdFaJh4zdZBdHd6LLyJWhx8N5AQHoo
v5+NE+a8ZP5Y4TCJ2gNymEsaFhnpQE5sTo7ly+8LwAduQIWgw00w1ab/na8/+xnt
vUi4eIQmaClEsv7HmlwXdbfgxjmvZ9Fn0/kUSgyoPNYr9XmiLFkEKrApUtONlFtm
WgTP0puP2nCvqi9cQLCjxAoxTUYcbPF9A07+A9/zcR9QymXv6umt/GS45LHJFVi7
ykmSa8xMZP7Up9wMPxAyWy93TMjQurlcGiS6+3PptEHjbs8rmVHc4oilG+gP4ZMK
6FpKTB0LpOTo7efcbELJM2YlJ9NfeWvxYruKAdnJ4g9iOnSVqjA0qZx/vUXbZtDF
X/9VYx9A33F4X/D5mbz+lqfNY80RQboHHsvd0jKH2vM44SocMlf6TVPRTpZqz3a5
HGirE8zNAXy2ZPhg/75ebXsSoZW8rvGERgIT31X0jLaQuw21wyEpWX9GGK9Ybv+i
V7eJN3gt8EXdFo7RozS2ztYuMN7+0eoPivgzC3OsR0uYCQI0yr5+gcYo/8QG7Xfy
SBD8T0Za/OatOfGABqrL4Ti7g0NgatpAmjMOgvAcTVbOJUcAsoVxpzmefwsbvgPr
rL8QXHAE1Nn1IO1IQwIjaO+XUmG4zVlKzquRQ06AhMqjMqNl6ZV0bZF8bO5/u4W8
Go6bV7MpKetHjKO/Pl2NrHZFpa8jeHuaHMe8DJ9z/JJbxYUySb04N7yNdD4U0FcI
NjnxAantsCI0CrKyIWJDeQ56bb9POAgggdxXsJR1nGepynLFrr0Ac3iRy5kd+VW3
sACQFyTfy+ud4kXPbMAHE10F6Xql/u8qQS4+9ECN+AjFoh3M+4GRe9a+eOPMDI16
eXkxAw9M8hm3EJbPGV6f/bFx34SBr1cJgN18x0LPcEX3ZB0SxRZxQylObcIfZp8R
gjjHK7SVdjv2daelEJnV43SEp3sWQQuo45rHcmy7DWEv/xY8+20LzN3N1Ge5F64a
WjYxQz0ac25Dy4mI6eos+EjmCt1aw/GuxgoJ9lO/3NlNvZg4NPjmyytZ9PW0MTKo
9tJJy8m5YLCSy2U/WDeQmvcj+ZvfShwWmnthC4C0LTLrqbFRGoHW/BTn2lE5qFIp
0k8U6VwGv+O38ff9EUYuVgXT9oup9+uS2bqQWl+6oOt0tEv6h31N1TjckHol6oB4
tlid2mraM7NHF37kFo4vfzNhBQTXM2Ws6LiFmEGio7u1ulsLJF3lNUHPDjiT9jFV
3SARiOAP/1B74HGH6S/pW2nPRIMkUYZ4Ev9uU4XoSfqgX8ZyVEzHmsPfl8I9y76y
AhwWzWXH7v3RB75+Qz5jdLzzJRB0BEBOgaJWy6JmeYJhGLWBhfkS28Dj/GLiteAx
BGRSboAuEGksX0xDLyUjKj7BWof+wKJ5YGqIDt38l7gS23CLCKwIaymLN5YOLKP+
wJ4eeIf24tjiMMMfd7NfyzwTzquutGiLvm76mHd7Dr3UHedhRbkExJZryREOoTg1
WJEC73MZ1R4Jaa0IplixrcHkvpUwuFiI5nGAiRLp4fNUzzYaNjuQTK6kLrDYNepH
O0K8452FPgVXxkvNc8C5CxVb7QnxvScO/zBM7++tmRmY6trX4IGjExjwZbHRojjb
+K9xRb6Spu0VNbIVS+u9AnRkcO9n97flgBHNX3euRAlglUjvInqBVKUQGjHeSmoj
lgFRiCdY/FzBdfKah8NT3bKJMvKV8xhIrJ3j+qlhDGdkk49xX+KKq6gN2x4EJjRp
xNGbH1F6xUNbHTNRch2zfgLHtBEYskW9aW7NELIFR0ZDAWRdEDvaUyPRBCgsqTjE
fglJfnvZTu6/TW693/Q1vfTsr/xjTXb9dwRZqltTFXZLOnhblEiMIgbQyqz/EO/q
WZFn7nBFAB+4u0OCyB8JqTdq00kUp0Hc5L3gDLjbhrC2iZXogAzxKsl3TAo+bk68
9oqxw3MazP1qWtNWnvIQwDTOWOxAFwRcLmkSYbPvxSlSj7Y/bnd+0Dr5irtcqp0s
yEask2Swcm9cC2hSNMbKrrbtCOwLNsx3X4pWmfrOL7OWqaxTaDFu1ON+nxwkq5Np
5j1hdJZY6/a4uCkhxAhh3IFIxUXv+cpGi8giNfn1Ixei4UvdWN4xYwZDHdlb0XCa
fJyWEKKIe9Dhugjg9wKwnGkPOeEMmukIbcmJJWbfa5+4pcPaWkxXqItfZk9uFfsb
7AvfHq7zHQdPPn+2bsVmbmhjp5dxUgL9JEEzHnDom1Ion+kQ0ya/VACfqpe280Bi
i0DIFdzM5fPt4E4qPrSkvlPtwhExElyIWjfIAt/kc3pOYsnPtSl5mxKbhP0WM0f/
W4snzchp6/d6DDJFkaauGpt+NEykaiMbdT/tOdiAixh1gpY+Hpz4oljEgLQw375r
iDv7fUDGz9WFZ4Lx8Bxm8WBeEdPBcw9m9SA6e2k05lQO8xcNbbHK9rHXK6j2Rujb
11Ha6LKip9OC96yKgJ6zNDWJWo8x9f25Je6x+wwHTmOWYvFYk9gyxrTYOsqkqgEW
A4HbfDySMJ5Cu+KHFFcOzlUXfhoHUB8sek72r0BI4hNy3001nSPg77CTB0+J8mXO
aG17Onqx5+ymj0Ht68FmLlVlAw8EL+c8yJxjtynAVtOk/dDw7upJ5zsakQNuqYUa
GRUJ/OiJ1cRoxX7AD6dEJga99MNZZVd/cpbOe1WL8aBiHJaF1yC7qGFu62uuE1Rm
TvJTm9QbchnIZBQeMSEi756WTu7FJwyqNslSA9pOnDxGycq2DOCqQM8uPkiRF6rP
CFEKN6FRE4sMpPNgZl5qeXEalXXjm/+A160cix7JQSjSvONiei4srvSCKnoy5zaA
wGzkGndBwx5HgmFENFhzS/P10oDa/sYq57mgGSed18+kQjdoMrD8WqhUretO4Szy
WrdYCCCXbHnmNNZuYRkwXDBfw0cUgtDVpuw0R+h1+PYj8Zoa4yTk+TFZ8uAgSjYa
L6FYiNKACwyiof0/Lnja0C6B2OX6tVuyOe2SQtJ6W8wLRJoC1hpuPpLqF+8iljEN
6ZOdvyCxvrD5jgh82e41e6Xh8XxUCNX7CKGilQCBzSp1kDvn+bAscRFPxeKibpJ+
a43KPKqFc3wngTFKd6aX/Q6WbIWOMYtdRtpJtTRBaxkCwavrFb+SqbGDmIyPxCRq
T3Bt9OVjd5VYel1lXKdTwD8ItWdxEfyyF9sqizAnTbMA+/YR94gwx6Oie5iUTE3O
lGn7SOAcsu4pL0lYw6tndm6Mggazx/p5r6AG6njF9+zbzFn0U9yAFBt38rvjbmrC
DzyqO6tknyC43BAbXDIWOlCNxmPs4CiTWp6YcZCybSjxCssXiNRgG2pgb36d0Jfm
49weER6+dQmiMqHvuIKROfLYDtMhHqBIwC3Wv2NlJ7P3mOZaqpCppg6myv6gFzUL
RLNPa1E3yBrrGU50EL7lgZHeSfmEiNviKuivKXKYnyGYE9Gyt4owoKDu7BqfKAmG
4hH5ED20wYI8O6YKOi91rup0wruphT8s5oSxljEDPLptfwMvA7PUWwXCTK5034up
gqXNzf5gsJH0VpHCyhj3Y1Bfkt0HPEmhMptCs7JRylzvMzoaJsghoRKrOOByWE4i
kFyqbxW5vF+jwyY1mL2izbjN90v+EqrnrziW6hW1EOkz68V4+8RV5jLJATDHiN3o
qF6ry4k3ZvaMkIjRy4lvrtdRb1c7kgq92MjYTqOOGMoZQO8q1FU9vKojGX7xA2su
kE8CnEaF5XzEo0yvIK5U0qq+XCtbPGQaCx3cQwKtWtixxMtFKk3OTbSpkToWFDK/
S+SREaUhyOc0LeiYARbIp3p0pZaRRUtLXjGVM6dtINRW+7CH7SwNDCiOYbI/IDb9
ZF8E7DbVQEwbzRPpjO0wb25581SUKzKaawnvsX4FQVI0H1lMmG/0yXFHETvUkfjD
qbqN0ty9CTEWIZ1kWdokyiA6B2Gn1eINrGAkt5Ey92V5MOhuMOe9Z6trCgkb/dsk
VZO4VxYXwUC4X1mCV+xqDwU5EPdIrt1c0QYeMTOV/d926XlCuw870ji1Yzs51/d+
0SGGQT81eZxznBDjzhlEF7l+NW08nBvvApXteMPNufe0108ftl0UJvD5IgTYjiix
bz2K7T0Az3MvFyECb2HbLAAclDTmNB8rqHc5WzrnB78OosrXYXWRLEvNL8m8r/IL
4BZ4h0HXkLGNqR3MzNtH6C/FBZ6geLE/3VP/CldlUmUMuN0LA2agLDb+n3K9QZPt
4rOY6lo67/27wJDagFFzIAYuqzJPqSuLyCrNTRhMEWPA6BkvVDsMQVW4hJBQHYVi
jFuYJozRz3u5Hze2NSIQ3R1zLgS/zkDaWu5hmpqedKJzHCvco9oqgVHGPpRcy7hv
RKylDQ2y44M9cstryhQt7e35YcbW2IFmgug5y8+Zz9EgQZjJ+FocBBq1uPPc4EsK
qQO4U00vnRZbrCeODy45J6X5Q/0uhe4Hsutq1geHLdS9YAgUhdetTSAa3H31qUIu
dxHaJ7YQI0FXWX9IhTphlmtOuXSabVdbI0grppi876kxksMPbrhwAvh7CiBDDemE
FgPzhDlXIgt2o/mQvqSki7TF7yyq5hyQZyhECbrRueOeAkeWZu0SLqyERaASiS+U
Jks9AnMX33EM9pFrTOR6MCWZc6geVuMCDq+7FBeNoJTAMQuxitsrLtNlVcbdVxq3
k0d8tKfvvjzujx5M/IneN1EZqwXsmPmeh8XXe8G+V24EeOxfkUHYnSejsQNqzxuV
GyvEWeyP+E7qp4zKddKEgpmnZDKEA2EUtVGQ4FJZp/4OeZQ+UPxEX0hS2Wl2n+AJ
oH+Wyc7XJnoCnqStpEl3TrBIpLsfO+LMeUWGn9mSllELPaAzbO6pbGBbtQSUiAdi
vc6rn5nNaa19BXuKYfKOD5ftNC+6eyaQf4LetXmMGzGQz5DLIlnAEhBzwJs86m2i
fo+bwlKbkrmFocyf+7WMjUDuX/eP9HmcuO9SlDnXEy2sQPR48djqcph29VGJGh1u
oy/Nwrjber7eKD/tHTFOXztY6XuBfmY4kHnU1+s7bk+vvt03XGF46r+gaVwaC92S
hoodxuO+ZVoTGhGmax6BJcApIpfNKCUTmrgtz90IjDBP1TP4C7F6X1Jya0LBOqiX
hbxNI4BxXNk5S3rnOGmD38dPiCaqn5WyhmN8Kt+6O1Sn4ldEyTJwyUdFrG5QCXWR
D2wdmiVeXwlz9R4rOuKGoC4X9Vma1HQBVx9OAtAkkAcBzTM4CeDVkWfc5WnJXzjh
uS4U/QIlcvkWA8eCM03bQmhLN0g/lyM73KheLiyIVDJR7Py2mHadT0hR37hMbft9
ekuuqlsqUcpOj9XfLme0OOysuLVuBe1c56yaeiPye2HaBDWBHDuojnjbKMmISi4g
QOFXdi9sMfsWtmcwwcSPTsyCoHK49Qf5YLiM9URi4sDqsQam/jIYTNzi8gOe7aKR
pRuSkgiS3j0pKoq74VHzt574T7g+LqOrJFQJ9uLywUAoy893IJI+d5Y7R3Br3ASi
2qUmAnqgNkEr3D2KYinQRDJnTAmTOnqPTnttR3UgE8B/gU/8DyiinvcAYnFdMmck
G5g0AZOa5rE7BKmbs5/d4AIlRmoWrfu6FgbgGsIHX/QQdR7In8IgnrCTmxLxFFn2
6qC1agiSt7d7qKLGw1M+OTY0DQpQRrIqXNDa3zzheEsYZsXEjkLkYZp8vzPQAeZb
FUZoFamhZ5HKyGWWYEzAWTgtZFxWky64FLQ1ufrLm//aK+q6Rbve8Nv3R6tIiHdA
E97uBP2gElEfSIFlXzWJN7kn/7s66WjwQsSTVpe48wpIEI1gh+NcM5sgOYA+Z3uk
zAPmTC3Vcm1WLJRbyoDScs/7ZdYDXLGRJn3ZrOPS8qwGdxBGDYSpa6pu4I+jOUTU
EhafvaroOOnZhcr7Pj0ZL5tW8miJTaTQL/oBrqjhQnC7bXojzK0bmtFaZZhtIapC
J2yjmIJvX+xJt/7kYvxFOvAHK0j4ZWlykfqqPL6+mxWdmUFQUcIYMVzHPWpJxooB
dk8URNLy76rDXK+k7LHh/wt+Dcou13LP1X0cNS78KLxvbXcU7XcX6xqGluWreFda
AXDol1oNq6azv1cm2yfkhXAoM7p6zd/uLxa828x3+fHd6tQ71Paw5Y6h0BmwYj2R
rELV5ghEn4wKl/s45pFrkaNyqi3oToPb5G2P+0G8Noxqfm1uGgFZlZAwTUUDKNhN
GK9rDhqENbUeDANf+CgyOSrgqOl+AG1TWLbxB+uc5DsaemjarFIlGH7CTIMgyJXw
HflJiVHvSPr7KeXwlM1d+U6W7AyhryDsRXQLej19IyyGjQxU1WN32RsRTRTOsywr
qJ2QyTylzNE3nB5fCNG3zPvcw3cBG4Ym/G7VOPkwgzvrffHkS45JbENY03k8KCvR
M2xiiYH7YyMkLHpbINR12zFWpz0TFvTuEpXhXMG3FjhmKOEI4elj+4cXJyV+8ju5
bQJjpkTBPQCW8bOCEkabBQ7Aop9H1yw2ZSPBpE3FQsFX7cukiTFWlrBZa3AqkYSF
uwSS1qtJjk84uOkGDkP3EYRx45HmljU+eXlOJ31LHSCFOdU9KCPkCnRMtDV1ppeb
hVFbgcySIwHGwIHoNBbsQOF+okz/REzymsUwnnu3gjCzo9+Auz+Uy1maK0HvJep6
QmqVnEmFLZQ5MyyB5yDADy/tB4kTOeuqMm9Ji6DKpeirFJhrFo4AXiEc00FLdte9
fA2I41MZXlYc1ukT5zuUeLepoNY2VqLd4ZQ6AlZ0dvwVD+mogixVtj4/yleIYPSu
MP2/H+TiYE0cV2A0IbVe64HRsxZ/XrU+5wdnWMkzRon0qY4MQmfFEEYGjO6I+b/i
pF77vrChzaGTiWXghajn7HMvPcpLnqTVNpzINgyvBbjO0V00e/rreJFQkdaNEJCG
Mzw0KuMB57R5HLDuyma8XF6EJB+cyPQJAMGTHsLHHPXZz1DXaLzUIAHGTrn4XHlh
CVDoNOPpODhIb29UsRJv08OXDUbNlL7azk60rQhE3G8ZOATzdnYBRZToeRy3jgW6
gMo13AZmk9kF71mfteYLm2JUEwj8QFLobzmmwRbEc1lo4N47AxSmgZZLTLxZoIfs
OtZKl1uJ1mYDSSuHTRyWILwb5yMBYULM/FEVMLpX0PRRAcTkNsdxa14aZyI9Qth4
mq4L8XyLhMuWJMfsPzbT/CHXiccWjmBObSrhnk+Dy3pIHctRtRB+CJpcoJEafrP8
Yp9+Pm5+Vl4IpYrUHkAwI0ozNCecvyvl2EuVARIJULghSWZwDS32xrK3fpfz+IFM
uKUW6ssaRy25ksCWT3aXClkPF7SC6Mfs6Txmj4TGPWDAqyHf2sspFlh1L8lIOqFC
CXUVM083DwWSDxpOe3vr8a4wbqV3v4HmicgXITGeQBnVbMNqZlcXnvHgwyC2Lqd8
EtOiB4FmtR+9v4U6S6XBBcHFybhU/UCayAo+pTWpHrbqoUSCqa8ArzRbF/NrxdU2
48NzPiIuUV/63+WqchJt0HTi35aOtYFU03WoNI/Idfb9IwTkejB50Q4LVlftagNB
1cR38DIyoesG6dDxQGraQakILDESi7ANoWIVMBiF4yEc89K+kww6aiAQZNC79han
EF7XHt01eQAJvkPW3minUTaDCDYX1NRrXG0LPTCE7eEsH1LrPzOq7FmKmwR2vv0O
Z5D2jcBWwa6tj50c8YU6vKYpW/P01iBThzgcrL6gT4OQjYwdIeR+KpvuT2l+3LlQ
JrVm6h4NdGMMNGMNTgk2N/qg00AHL/5E5nGx/t/0jmFLVc4PHEguVTuoP8uP8lty
m+yUMvjTKyvA2rXUGiRBSgFYbNGcn00Xj5ttfmws5vOzIfXgTXxUDlWaCVl7xFeS
4UQ3hP/iq0Nr2NGig01cpAt0NBCl2sYBEeMQZW4ORcrroJoe9FtsPeN7B6PYHmWp
s/UttM9GfyzTRdHnaVjtpv/L5KQwQ6NTAmeNzYU+cxGpCfcwExGtHVEfet0nitaV
B8XSEPSfk2kXcEkVf+xrEMmLWnvrxE9UmCOSMciB6Ygkfv1wbQ1ZmHwHzmVwiu8m
lPmEsaN9anmQ7E/F8idsCC9j72FvPMFcBVpJS/dIuyBDXKiz+S9wI0OMDH4Y5Fos
dFDQneuRJiqGocyGBokZHu3BDlAD36eISGQ2B8KILjQFXUXESNTZXBLK0T3EYHd2
j94z8aRSy3sK+yN6z8QmL/w6Gq5fKLlTSsIaZnozbvhJgVNy9ZcupcZqjJ6YlAqT
DeHK0QJok4E8dAK/dCQPcRDJ62T6OkH1Vzchg1XRWTs55VnuO5TFaAxej9pKddiz
hPsr/4nBjLI4Z6J4bkRgzyYpaO9z2hImd40e/zASs9kVSl9/T+kxHe6eVhN2ONp1
Hc1bsJEItxlVRREpL3aC0hY8u28CbgzF/3b/UpP7d42WvRQLKU45OXpr8Jm5CQrY
aP0rfRD89vyFvAdJf2IOfrbzQLE0AxzJgIFhk2ddBBXMcU5xOTPTuLE1eUJrmMlx
pc2O7RGNSIodFMVPsc0i7o5+rdWUn4ofuBF9W3X3e0npALiwEyMPT1YsAIP3j21M
42fgLr8GNSLEj/7EvzvRA4xb9F0cuT5xHdcwnnYEu3TahaNCONMrlz1OzjE5ssNf
OAsBK38W0q3Wl2+kVxOoZKvYT659TI94Vtjd5Kr8zzQYd3mp66ufdQk0kizYGXEw
Z5kklPPK0Jq8m7OEFSvATtSkUnf6DAv0QyhkhzG1Om1aVBsxzZyLupUbwaFE5Lxh
P0c1cADowre0oAsayOEESfmpEbXe9NhZNvM/G1oGsMN8gaYsJnanSCHsOrFs8BqS
mLBxVktp/c8pds1dBaXZ1kY+Tm4O8C06JU1bwKMGponFrt9qwUKJY3T80id7XbtM
MNUqvVsRxhzQMuEfF6OB3fER7goVcLzkxYHQ80E0gioRFxoajQqFd0nZ1S0CrKKS
4wz10iWc5RXDsR9OM2Yu877xsqIPfla4Gq7Oc2/aolv+XNEgbdqng0H0uWAeha9v
dyKpVnrSaScEanDboWZKGRmRwCmqmXuGnahvXJcs2tOUEP08y8FerH9JwdZMF6Jt
RZaKHLblYWaG8XBer0LVf+275DMx8u7RVOpIfqzef0PZmH+5LB/SEu6fgM5a/OHb
bbfNf0RhgRF5s5WibOHiKfxXrso8IiJj/H7FhXzJw6u/fGzs2TxIPljomvVjFVjl
W+iFdXm7kezFJVP3UrEF7K8Xe3iWjzu69SvPvcEKNLp7brIwkjAJr0Rd6fGxEl+E
Vfx7LzKaJRHWBG/5vPs1ZeRf0dmh5G7SxzAumTs7QtIVR7oQCk+ZPuXXroCOFUO7
VvO3xm66WUrej3pvZNlhF7WdhUHv/ifxu7Ip0hIB1bQjXin3cL/6S1cLKjtDRnyi
Oca5DL8hG7VKHVHcPlgVEgE42tmOEkcbvHab4L4xPh4De9seYnKnNvMg3zzNhzHp
2llGreGDVD6UbiGuPa8pcWJ+xpEudB0l48Qt5Z1Gfyq+Vs5NxGHVRbEXz17rR03X
X8lHgEsa1o3+1XmpI8/uz17LUysC63Ws8HqcMBnLNbnEhdvvAetV5RVPFH8jHkFE
lb7EEc0FkQx5Hp/VkL8/RBfsfsdMpbwP9CzXGyUojzMw0yC8vivW3G8jmmArMOen
+Uh56/yBUxLESe+sF2r/j7rwcb9CHclX6aeNQUSSla0n7VazhGEft7Gj/BXa4xOP
7OmgVR4xpplFDOK0GZmCxC5PVg2SyngKF9OJmHjsAvowHmw7CI4SgF8g0Wspv3f+
IbW7x6r1soyT9E5vISoFotcnOoEn5RBi6+nIYnlMRdeG+Ck/UF7VYCgxXfeQ7CSU
YpCvf1HvHgoJpMGwMo3XKR01zMYVRlwtCqg0p30HCrN2T3LhDved/dYtKAp+EsBl
bGLfGpoCE/i8FOfTt8kivF+R8kvOVUFxOqvz2c4K0vumYx8AqVzrd4Q5eUv7nSuX
iP1X63MC6yooioZZRZggJ5vvcjH6PS81RUWarj+QbBDQyRL7MIpPK6Zn+JLzYnSL
roRonhDXY37K8zXrKzwAQc8pFqPSlzxbmAPc0ajsGHwWrANZ4CNcnnqIP1q6d+jt
BR79z+NYIfQwWSAyWeBkC86ga8k+Z62sA1XZlp4JBM/SXRbqQrh6FjbSnSk8p9cx
/yW+1Ik7cY/RZfmAXyDfF2LhUcNuoaF6jTrR2FLSWt3ZWUoPpXRF8pC8ooBIOPl6
mEcieKzWkYuzqg1Snn37GyajMgn3lpr5iJ6Qprsq+gr/WISh96EzdXB/SRaXSC3i
0rdwHyYgbp6WijnqSggYH8fAnu9LKfNyjAO6sk8KSXqmU4NfFrnkqSpSlLSmwGPb
TpG8m1gNIbtDGn72GeU2BVp9OyuT+hkL0mpRM+qOKrLG5aipUKUrbTBqiZaz7yOH
Kq1KODDJcgc9tIa69CxJEIbLdyrFO38mmH3gWDG9Vz3bD1R22B44Qla4PhfBUxNk
DVQw+AYsq/JK7woqjv9PNlTXQIzzi8+slsNeirFewLiBXFb4ff7xUh4bVID64UYD
QP5fT69Tule6O9jg7pbZpLzE+Qb7Jyyx0KWBLW4D8ucydYBiBPbU4CMQukMVMj3p
zvmLMor4cFyf6+KXeUEwuBT3sD7GVMAlC7Erqse4OElzOHGrpKC4Wfj4oSZSvQk9
eEEfD5xkr3ShZ1+8LEN+Y9y8zNqmzV1SUKMU4zdQzlIGURZUPk5UStP4L8zTs4NK
u+R/YdUnv17ohMznfUqxvpTgKnSBh6MaHxlVMx4mmkHbOc4V5wc+pY1vBPz6Zrf0
3jGDyiui63mWf1nDAw3KPosMP0ADaZPSyLjGAxg9fARQwVmy5+T1727o7wD6VLlg
yKl3vVnP41jIAOZqG+0jhZ5sJH2G/tR1epMabt0iPQ7PtEWd+amGM31Jlf1yDq2G
sYei3flkMXVEEDj15UaCXYZ+/yCzpXc2UR6uLSnp+vtFftbZxjISvULyLRgnxWJq
7Ci5tdbqLy5ndyDhVipiVCFb/NwEmeQqegr5dBBoyzK3MkG72KgufpHB14vDGlCx
d40CMzp6pAD2DD4E8VUivj4E7Ezh6Vojj6npXRlxT8z9iNC9PYEvnLquER2fCuag
gmc5Qjuu+8pLZXpsNGHHiVt6W4exD+ghNRA341KrC3oXCocJCAjzJxsq5XHUSfKz
/wW7XZiTAwwXB2T5JTDzZTAmsheS6myzgkrJ/nDmPi4GP/ocu6981injo6MUHZHH
+3Me3e1VaBIbQixge55g8A5n+1DGg9YVWksEtf+eO5T8+yPKOfKu+HuwqpR5CSlU
UfYesVOMhgkgpAe6M06WOmnOA3zPwnq9rcgdPijXzWMbjIvcoaIrG7EDXB1SyQZR
Zi7AnKQu2FcYplXcPzVaNp4z82G6lFCTtz+rDZQCtT7fUseO1bJSyQ/BwC7QBBPM
zgAF6KuW2r8lX2UhliEGqfyQCqyonLPPAWGqRo090DrMKPqZe2uJkVJ5B+rBtJ6P
nPhifxeSrKQzP9yFgpWTl7BXDO5IHLPrLvWk4gO0qf1t2iSw2k7TXgr1PQ9vEcsR
95s28jxT+mJ1zC/gd7cleGXjVQGsrMS+gWft2MJMbsdWeUn2SCh/yEJT89kH4Gq4
O1why2u3g5jYuWhas0g4loGdQTy3/DtNEpJqOhInzHMCg/tmKJi6N0ltUxkoalZf
z2YF865yPM3ZLf4F3YOGSEEUBGKq+74SR9Fgsyy04BtZfQC42B9X0AK3LwzLpyGI
bb6MSg43Gac4IkwfYS1Z0kqRd6mvZwA6QcmAotIvF/GvkDUSaW41UMg2I72bfksA
FQ5J/fiN4gAkL1xFZfigTNCqhcZ2/R1t9Wssr6MyLZdoWJJnyA8V5YCxNg7S2XvS
lSrNn4lZQkoNynim5uIIv4EatwQRFmBRjZc8BHUmdYLNf5MEvn3Mf16OFa4eM1Ep
wjoQmOq3aWuVuMDeRXg14A8LpA51HI1CB2PqOpBOg1imLMUnWySJDAd+bzsgBUnY
hSgXg3g1nRwfsTbfRwhqxCzcTlIdjTmv12jNiAJ+hkySCEBUPLJ1ZOEE/tfbetIe
4TmMu3b+cI06JF+lQIVAHxDQfMKxdpb6sJ5z3DQLeDc/MdxPFsgJhl2yOdvsFGF/
lvYYQ6QkM2UkniiS+Rhcp/IG+L1ZV81/3rTpnjods0L5PmkWJM19/hq+JhL6UDyf
aPsQDUAe+R2kxVp2136/uzAcQ0jPa02TNkpdzsHneKRITA0zgnM4qa5w8dh8Rg0t
MOojbtjBkwpgAL8ioyT4NcOm+WH00czgeWDrJ4MKILDufjlhRV+bkJzjPkivtKdX
o1pD87eTaIMfzFRCPepTe4rvYICE24KhsQhpmx65rJsJx9/IgSuqEw4QD0gQdJmN
hMkeRD5lsGugNj7PKVAKD9ig+8ET9RhqMxhZbu3NG198gQas78pKxKtqnLT7fwY7
1LLuKPuicliXRVSU/qWGI2k0Vzk04irKeSdtOHVLaVA0zlF2Umu1g34224/hYf8a
Hp4r0vNZ54anFrbsd435kfmjvQdJfxa/onMSbP3pxZ9caKhFXCwdS4ACq8YUdimL
TGlFaLE7jfwyfralIeDYbqYQk2ytV3lETmPheMyuOE2Q29HHB3nObhfStAFzsC6b
RPHnMUEmqX2/NnthBmbvoz9RtNUFgwmPN/cXQOvacivC6Ch6QfPCvJxkJSU6HkrW
f9EDfRsL6xsiw/0ZlXmMuVdEr1JXlCk8jWYX3oN9IdP8yqNAmZozVkUbviWkf+R0
LsG478i2JmWrdmcxiSzPE2m+49PVrP2avv9tkPa8cNXp06G1u4FRWzy0wOryEKRB
qScQC5qBiqOrFHliDTyh7vBsRnCOLGjQXbjpqxoYm63lPJ9aZbDGkFdaVZncvXys
SpP3ZXfbiF5yosz1//Ei2GmamVLn4tGqa4D6MjOkzSoCcAl+azzgn/4TPanMSsM5
jnFL6P2Nkzqy5jSdE5qHmBB3J4R5j6J3yw7Z0ERMKQoxcsD3PD825JX4qq0PmLfN
KobM3zEMrLb/48tJlWwqs1RgSMuQHqwNDXR4098zMrCBE5nZLVUuvstnRHFKkSZv
efFG+9Bg55YDdrvPju9HOnKaTGj1uvB1rVDuHfVMp/I+IAS0TGskVKMbveQxqYcc
C6+o5vqi+GOqIguiW4/aySb8Qwto8BnbxLhfklAvfXTD8DmRXvmp9AT3TeUVUktB
rn7dCWbrAyYEWmw31LZJY/Av5R6Ax9owivPDqQZ7ZQJAi/yGz5cpdveMPsv435Oj
B1aXh3UuSRe62gwZFP4DVLDhrB5PhPPywbq4hohpEWimED1LCZ93JopcdQpoDqhK
1v6S7NbHKz0wte0CjmJkRIyxzh35YENYH225SwcQOELVYNNg8GhhMVpHAAEVEjED
eUtxe8q9KWqvG58T2Bl6J594ChCRMgvbTuX4lMms3X34G7X2X1RVDu5/v0M1PnKa
epqBO/YkSZJ6Shzk83Qn5KGvGjo6ZVfHp2/MA6Epd1BIhrO4GnX/h91ttGaeEz6r
iGXXdBDPgmSVLQIgWsc7SrqI8BMXeaFl7tWFFXviqcQTR/Dsj6NQzTteZ7V4F88Y
TAoEoUpEubnSiGLwsfYqY5ahrmN8nrKYQXGVEM0Ux4SkxyceeXRyD930nLh80mCE
2sgzrAfPnAWEXyhnD2ccdHtv9INiNOye3XIPj3Ut4yJqqI+muzDxHvrhc/NX2YYq
0tEW0E41r/sPXEaJEocQOkSFEdo63UFJ0ZW9qXo9i3Ic9E0QQzeiWR5zm/9K88ni
WsIKeRrTwep9LzBC5xemRpfPHbUJEjsLjld9NgWMgrJZgjN0CDPtTSFgaEhD6ojC
dcL+w/kk2at3peDahsLcv3lQGSetx+4HxwdTXQUahWjvU3pX6Cw1V35P/khHsHgH
0RTxNvYJ24pQIQFVvTrVga3CbnNo1iMdzM/LHBP4JylgkOu4+4X/TqVMycDO/Gv5
/gfjcl93tqm/LJByLpez4RhGDOKZrcUoEr6IIio5ljn+ka6nJVLvB38gltmTk798
Q8nM1sVIiIk7Zj8YL7BmvuvICDSu6LpXlCAwBtKxIZEI3Hdc7KVpc6nfE2hZMc19
cRQYR4rJWqu+MpaIiSKBihQJxMFkmkS7e19zWtLzNTfpZHmcv7ElLvGXK8BiDTnv
WKascJL/HdgFUdaxPYPObeKTYwNVMJwTvgXZ8v2WoL5xEk9i1mGnxu7T7iQ1UKOZ
C1CybQbfe7Ews2UDloudXy2lkxM81FCgBlejc7++me/JzBup7zNhFyv6WNBMTulq
PZBEvUe7ksxc/NaRUFQb00oVsmB/0A8wbDJvHVbzujtE+R4WpX2Y1IDhfIqMBgp+
n+VBf851xyz7Jbmu++C9tq5+LpqXpT5OXWBkAzkC13d4SLgd0UU0wCGSvEb0OaL3
Jc47BI95ZJ0758YbrJGzJVeRf5T7pGTP+y7aBFho2whaau4GPt5Iw/IRFVATC3gK
KdddLuNWFT2A2liKCYPIc+GLepzNyENy+WdCiKc88v92Io8ifxma6VxQzcbFqMaL
cNr3DO1UD/BBrertZdbJXK6F6646P8kdF0rGnBoJchrNrDVNHcOpKFk6nuj90lap
AimBCLxy6KgtpCPoNJ/gAJRENcgPljkKawdKWhTAOzxZnynZ4gVbqJ/FDdnnGd2A
ScgDORUMTEMw9oSTCHyzfSZUnSpRVaEFHtlEQsRU4QQGaILwugWnWBH5A9jbsgqc
EbkK3j5kReU2tDdnEGTwk3J5UvnRlG7TMPdek+iLm+bqtlgPmOCIKjwpIA934MJf
aAHUkPleuiCPb8MpEguggdMJRKds59o8+XLeLKUPJMUejURgTTXb6IhQrAz354NU
65LUGkr9XhpKpbzQFpDsScUaHEXGlELnLcJ5OpAdk44Gor+xUUtAEYziKkid7B6C
87oHgD6unjPJOyZG8jLDjMRZWjR/zq3FWHHIJCs0qxZG2EdplbGMku7aQOewpTTl
UNtWdNces+TzDD4FGnhChRYUSTCZGSbLuCmP706c1UiU/yLXT7ykarLPVm8o+Zn/
DdF3ogxrPty2wIPK8EUt1qQpRUlIpk4DFbF5nrRAmA+6cTx2wTJX8QYze/dDSv2D
wovFxYK4L3srB0Idp7k/NcEQrxx7JjpPZTzPGXPRc1uh0F1vo4Da+9ZKYszbg3rA
pS8CBoubK0rQYINLp7ZfeP66zbJWiLYNQauHjUR9zDmkD/UQedjciSb8Gsp9WY6U
ojaetpu8DmbSennONX/OL98zaWBzVyRuVWrJYcGLdoGMGXoGoMmLj6t+nYmD9WNK
IV0oZGItJ+TlxAvrvBF0aLkKVUCS+IHxLpv1rMLRFNHfwQctB0MGUmbv8A1NVG/B
3lQrND86hd2NT9LUaNPqzLkqWezxkOZKcvvjE5K19h/h8IW3LA3d1Bx8rSbJ3RLV
iTNxfJuj3ybP02LVvPk+FC1Up/D7zX2VhAXXbz1RZgegJbo1Gu6/If+CMJtCCixS
wSDOTPq6PHvB6WX3BhZGa7zBBEzdfphlc2HYQagYAAzRMmDY181Em4mJuleyIHMx
RcExfIH1Nuzqo/Hg8cMNMFTy9z++KXzyM7lEa5Zvj+CfK990HYsoivIPbMeMe5eO
Ci3C5/ttsALYkJZ29cFBDfdCahJ05FddgnrKkAl3opqe/Ls70IXUTJ0c3JTuhs21
AzVEEdzvKdJcoC4kE/gtmAR2l1b35Z+3Xxb/fJTm5SaZF1DmMT/SK5wGqoryQHzp
buPHL6YTSXMSQA9r2wegcmJKA4VArCMCM/lHEGSs0UT4cZourJd7mRh4h9a8xTuE
2+0R2aCBQQN3guq9o0cSV+wgG/tyzrYvHXcv0OwgjV/DKHYc714EXW8zkOHweDmP
IIl3N3XV2FeBSvh+UFK8q7vDLLIMIIWCWrdzbXHbe8TFM87trAUD7L86fO0vdxDc
2dTvvz6sfXzjXt92Zxm5DTlbARrjykFZIeTJj9f9Z+dw/q55wIU07Ap+djdJIA2C
Q7aVZ5Y5HxEExjHpBsX6cWvYmYRf+6GxTgj0WO+Hhctg7I470sdsw/t3nyCZB/W7
YuISEVqqiXmOk4oBpBygDWkGbkIvN7cEduXeuHS7sb/gI4TwEAE2iA6l4iBHkM2K
qAd5SNJZlszzNKL1oNdvgsEW/PQ2uR8rxzipgz6bEQ6hM4wZPs+chCm+QThvcXpC
qlwWJ04cVIpN3NQtQhjAgyfxos7xjCnKP5PCJnHTc3o3lbrhybPXjsgYSB09bKMU
JEojIuMWZm3rPrcMSQl9K+dBq1+KONopuse4f1JGKfdECDNzrf2+Ffr9URh4VFWs
hXHxi1uXrSjb1HbmkfFqfvYSNtROn7lm/fuZ3bBCeLC6cocpKUELlLBLEmeIVIt0
cxOcBn+b1OXVh2tahxPSSCOTCMvkAkAFMy9N3vCHv6+JPq8vTR5CP5tfPXWqG+vK
N3Ss7vhA6Dir+WRSzrQUNGmHLDfBU749c47flZAcrvANjI2UqTvRJFH6qeE5g2a/
2AoTldkvi9JynY7Ezne029K3Xth8CCg5L2vDeX3r/EFf/+4QcOxObKCLD+9FpknG
YxihRuoctfMc3imARPrudKIVWkNbms+X7MuakriH9ZVm0/TmdniEdV7OTmjrXohd
DqC2wzYdNLpFjT062IXYPLWU3tjWvjY/ZOi9sKewXQoa29z04UVuvAr4oEvdRt88
Rpm7JlazKzKmByFsHOWa5PKQ4g3yADaTIAxhBtUpjnIqI6xCdqLEasd/r1WT+ZNr
xP3HtGy5EUJVjQv1Mdd+sWn9iFHAJ9SDNzShhAk9v3ui8X+LDgZ3NTcyIDCKg4SC
3RjjdDRwSxznIh/mZvdvBLIcZHRhCWJD2ze70zMehLZnyJo6CnHmJqE5ShvnL7DM
MQgu+KVsMSqzkdXerEo7XhhK2nkUir5TzLdlqww/YrZQVNzfvz0CEZmvMkXtc9Ik
gfE6D/miJrsmF1mSlqqZKQaYZB1H9U+ZExvGdnkxrJuDqGIanQMkkYr7FeB8SLpo
U0NOoZN9SVUT0shBRUdibi31up8mAgxWvggM0Vhfvxkb3D86NqXv55RE0tkk3ZHe
+8SxG6awjS6gDV3+7nO53fbaIReWkyezwFAy4MhCRG7WT17I9Ql2l0KODQDufCUb
gDHRq8ngZc0+gqTnpSo1cYouFK73ct3YuQ0h4h20GK98OddfD0f1VG0Pg8svwaDm
uLTFFQ1x/9/c+L55SUvrWkobO0mgLebjW+4v2LQ7XZCGockX8B2pZoo7A0nORkQX
JR2qG3GwkGV4X3VCXVUxudAutk/1sVteRK7cK3wa2ijsbuS8Z0PXQk3Q3MkmuNAw
bD3/rMdeobNhFLQQRjHAH09zktBZ1thgwm1hErtsv8ID440Rt2Rb/Wup3RmcWpRb
w0V5ilnb+ZvoE0IyEYtmFgRUZRwglbEni69Dl5YZMC4OLXUo4johcF9YJkqnm//J
9z0Wc2fEtD23z9wgLdfsPeUtslD5PUrO+YbAUcIKVV+8JSIytlCr/P7bZGx69Smm
IFnZcKJyeQXQ0Mj1NS2bYxpL8DhwPhKdqc0oDgW5js3ddRYcJQ/dQ4DPRWi4YuIF
ikqVpAfG4PpWKIKxBvpT3d0X0T3P+QqdQm1XcuEM+T+stYTG3Knkw8uP4vPnOYiF
12J8bazuenoWe6qPFow9V8YQn5iNh3UgCT+gX4KS1XKIYYKe9q8eP9S4jb7M+Ue8
uN3I4Uo3VoYBkf5Ij1+3EVxvCWkeXqtKNuSJ2CYQ1Nf8dZke85nf5/gBh+JqV/JT
6Gebh9I1tX/JmSbkKfjp42LTCT9tZDQBHvafPZcJuFXBGgm0hZRL9zzRfp20u6sv
o13HkTsJPxk4e+UeK5AJav+Zw0Q0bNeLT3DGC61C/8NbMWc6fChqGk6uLkZekqfo
5Y4c0hDnLATlh+Aa5BKM25b+pndoij1qdFs822anL4tWYhXexyXX6+HWVkk4SprG
7S9W8f6fAnpTLfD5kvnaSxmprSena8S0O5ga8RTnAFOtpVpTR103lLdYHuUsP3KO
JTwG0P+nydt8m8bVfuzYE9O0UKrpklRiJLnvU06qulstMTfkojIMRl5LV6O4yXWo
aP8eEpNjDot+U0XNwObnsJAY3mSCntXhvcDqwp8C/3IzE2KLvJj5kQvYOVpd17Og
kQIGgQSjpwa2r15Rwi+Xm7CmOKr+K4IXXz/5J1XvMsScRW8ODpXiRsqVvdUrlo0H
t2RCC4V1Fzr0pzbeey1/3mOZMbk/v2M9TtnC5KcL+ss2mZ3+74jMmyjhqMkWurPB
O8MNVpdy8kyqhFgI4GuNI3WbHVLl6Xc1QlJ+BfY9ms711uOtgIGnO25O07b1OyMf
jycMhoFVCkYL6oEpVB3+94pKYM7ynKr68WP9ezB9ZGClLGqXTRPXqLpH+9/0Mvey
1DIE9tL3QnRuQClCzExY3DR/dno5z8TOt7nxKZtWWi2RDi9hFkpYMtQP5u8+Z1L2
X8nH37HZNV8j3cvuDcPZ2Ln8t+3GA+3sJS0VcbXnmtCw/GCbF4rCyO5yU03mBL7M
o/jJq066pabaEFp1qpoJg90Z7iFboH/HHR3QzLjspqMy4GnEGYdP3IKcQQHhU2zn
HiwXkz0l/Fvx+P3l2+X04N5qrWjmK6xkLdak8RreeA4GGi6H1lUzshlPx1A9gKqD
vjGSn7nuLSt5+dDBM3bg4ArxD6gh8yc3B4h+nYgQVd6HSDy7JGcVLS0CgE2s4Vuo
M+NH52MWi4Vaon3B3VjGcaaFABLekXqJV7Lp55qWdNzK6UJgJaNu1QXcqRYBVjxZ
uj6jCuTSeGIYv/W9WqYpJ70xyjYVAmSHQ1Ybg1J3c/f7ubw0ZHiBDmOYdpKQXxHr
YK+2lewYdtdHw1BTM5yhzIHuFUvC4hIuf6tF+ol4TWrEDCNzjBCHgkemudCJINJG
i20JQ8xtHa5bgptBgNc3rdg9ecs4CESF9b/WURMQaNiU8p9LbbCodAH0UeMqckRT
NuHHVHGlLjTxLQS1y44tdZkt55mXMt4iUf/OyobzvGksNjLUWgTY1kre23MgsV0X
Z27N6Ds+FgUyrcJGJQ1x8s4O0aj2sb5rMvZOJfxkMhx1YL2O4+T0/H6R6PMKKk13
xHNhr9OLirh9rbksKvwUTMl788kma9bC9hPAsOH4kmEVBAseA06DBu/sbveKM4Ze
enEGD6z5VF3SUOB1q/phkEnvXXergqT3xUYD5bMEhBTd4IqUkQf8MJgRyIu24e90
EwmoOhi/b7pAaDhxu8L1KTO8YIDTu6fP7NVGu0COAfXabbwaO36ExvePGnvn9Dis
jUhwhc2Zce/nFQbBJ3zq5zMe1Dq71ri7Wc+GbMbZQ/mFM9sQ2EP8BPrdIUUFBDg0
UIl/cDSnwa+2hNUSFp2ebRrprf8kZM6RD04g+MlJPauv2w23wjQ77Jwc5AmVUqiF
S620lPgq1FGDXvsvfu3H4FPvp0L39m9QCAahV1X/GZgGx28oZo3l9elziE/1ZQVj
03XIkNYb8qKOVdyyf93vfgxJBswnizXj4kSTfW8uxwhdKpyecyKaBjiLZ9V5WIV6
9o31DHVMdo/NvWIQ1/z0k83G+b1HKw+3AOBLZmNAFjkrrGtgEEdecwCKMvnGLzjM
AZb7P+er7Q/dbL0V0Ya8R4StWRqlUUNdD5BxL553NV6hHZ4f9obE3NttMhUePAqn
0xLNJcUyWIhg9xh1y7PUCx0V0KBqf/t4sHjwU+74GXkdid+Q579LdogRNmqhHpl5
k4ehzbba6b3SAZgvn9mFLI9f1BqSVd/Pz8MTe6Hvjqo39ixa3QQnM/mjSg0pPCGL
T62nwB3+9VKbyOqTevS3RnMnmjVkuZpx7num4UC/gXESrhapoY5hX6Qclx+Lr6bD
UGODG6GIKo8Q2JOtTSWdVj9LSlJ2OTnPOngH6of/Ik7YgS4WHLXnPhnnxO4pWVo4
GKIveU/x7iXdmKdSbvILaOzd5jnVudaB38mzs1qLwNw4AbG78wCsgPrNpu/1yniH
E+lCr7O9Ksz8Ts6lwtyFMnY6k3VWKnH7Y6mYmlyb75N3ddl7OVM+aOa+BXCuGydI
dLu9mS9ohJ517ZfTuH+0cm+uEIaolinzwKw1b6NzdPXiIySXamYn2Hb+jWM5LQ2x
qgIuWA8ry4FdIqVnheQrV/9YKkniyvN/WAujOQgqHMa3QKI5e3B+iHNWZX79Zb/j
lIgHAjkszW78rClYbUOiSJlrLDO+Si62Xr7dzBPMJSEUQ5THJFiZQkREC9nWpOk6
zorDRN5XTL+l3f5LvE6pHtEDuy8tkBE+pEs+TM68m3R3+dJafWC3INFea5F+a4kQ
V+Qj+l2WpovsHCF37bwpkoCm5lEbSPYBtyVvh/nlEOBS4zaUicQdFTrNiKJu5dF+
SPunn9mhilzmn03FstFnu5anWM/tTyINQBS5OopS23KDdDhwugpoMENpcDRqalYJ
/b9pdgVmy3QMi3fr3FPo/EH2vAmDIehnnfKbSzzeQCaYJtgB4GD2PkITpqfJq+3B
AT3J7ZhG31LhJKTpu9HGK+AJAdk5cSylutdZxX1/27i6a48wjC5IOMOtzH40MwtJ
hL0owE1RQMjtOVY5vBNc17ii+qkPXpYrArswqEhudajIsoOfIn3A6Lq0A4iqvBMI
gaWvYWwCQUEBD3pkGDOOeFAexO8NdeQnJV+vB+7R0gbvPrhCmAbVU+lr0oC2idmO
FpAA8HLKnl8epqULVtfJO4jPM+h1h4y35Jho6lyvy/PTtAPjMBmwil2tAzuNEKTy
tSUxxGpDs834fK+AUS6pXf8dyBUwQiPDHh0oIaqyr15oD4bLpd4WGkgP8lKId7Al
/tsrXEo0K6QHz9Qu/zWdCkCg27pK9/j9ztulQ15Pro1Mn/d0y5HUXBZprIWjHPNX
4QLkM4Z7QNlF+S7VDM7aquGPIpcLE6WXsVHtvixxsNGRhToN8+6b5e62AQi14lNJ
4J/h7dFAkzQvA54z9zZb3bbGO2Yj4L7TqHZrjULZWY8JLcdGr9WhuVWqv5E7GT/W
578+9aUSQseAON9JUFlpieqoLG+XL8VV7VL0gMyysBISFH8M820o6fAzC9h4ZDbs
0EYYtrjh3zP/gw7rJd5LlvRIyHhmU+nUf9VoFY1v3tJBkjDz8T9VOs2ORuizHrDo
h4LkM9OiE4aWGDlJ8cht2gSdZ2wSyfSmnPdTVJGa16HGbrjLt8JiYF64rHYSUabX
JItA0DA9BsuhIODGVjhqy3KAZhKzbXlbCkBAO1/7jhXhCr76ghv6k+Hp9/7AwcL2
COsX6yprezOjKEg/7vI7agWMyLrlj48GV4KKec3opHoqYEA1RXzIC/KRp4QkQcEb
5b1CuunRhligbRx5pJeJxghoDLNfXRYYZ6QcKeE/NCIQvV6aWBJbzIW3U7C/Uunp
P54DUDnk+qrZ+q59qQRy0Z4YQXcBd21ZAmrozUbLkca5duHb0amMtD2f6TtHoEn/
tFQK4OJ3XMvI7Vh6rILQy6nEBeCRN05mU/2oZ+/h8U1yld7hb3Im/ZTOyUIymhbO
dkkvPyaGkOm2k+vkDSzYAkbtG2bLXaxAJhaAJHOLEuBDTLJq+MvTYqPMCeCgmHYP
lItJ0eJ4optCrIWxLlfzrE64yjm+Dmn4u/2BWfbum3xL8DSHwxItDKLMucWc4HK1
a1FdRsqqWjFByDgau3U//xYBBBC0Fcl5lCf8//GpbpfhfU17JrIbDDV0kBgLPhWW
k27V/E2ilwhxl41FPhdbmbNx2CO4UY9b7VXlhUbkBo1yZWbTYYu1WUbJ8Uiuzi56
Ut4PgK7FKKSyUvu5zNkxOKsVyyokQVzc797HZ1MgbaDSM/uzOXUCqAWlBQWz3fYx
uIiazPIiO8Vtw2NrcznOQ9bzZgDP1PUNrEk5fuG5b3DvpK2hB4W87bk928YlwhOn
gBcmXNRC1ZAg3upCgLyyge+oTaW/K6TNVLnNi3FrALrXLFYeHRvgF/JV6lcQo0er
g7/DDe/P161hBUwTRYtYCuHbufGuF4T6ueWcKdSJnb+bckkd11r7QPAyTKk2jE2A
geWBTeLffxMOae8m+QL62aXH6lr0bxd3zDiJul1MGFKXOZFSzwQk5gg4cpHFtbxk
GC3Zz34jL+cUqVyyN5og07CRtGwQtS6ozCDFMw6Aer6EEjG24H2gE7cQBFgMR2H3
8tnB72zeP0Pkoob5T5GaddOQ+667I4a/wOsllCnLVWuMuCre2pgffGytiouIjmsD
Cfp82w7cK6ENM3ClWMry8C3OgEpcVwY2x1JvF7IsL4SWHuxi3Yr4ODGQZN2lnM+H
mI33oCbSujdArvKT+o6YYNvg4V4UaNpSbUmAlAQzuOz+1vCr4UIzUWnthl43IFrK
+9D3ncMUoqfvk9UGyA/j5fYp3VL9AjIoKpVB+RFwAk27+Os/LPGyHxEdNWSyeN9K
10FVSqwnif6oK0UKEeAJtuj89N3Yls2Wcdyppc0MGUEtrd5UhmzAi0A2kowceXoU
L0o6NjdA8d1k8Ti++1vmDyVLOBKPAGyMbltK1v9tn0WSdvMvOtXMDvfcmafT3Cmf
oSAvXrAVyjbf5M398WgQZtwN3lM9ffSmQx2hYUANAvuDw6HQhBUmLsqILTVQMJTO
2l7cnmap+nDot4FwIAt8ijK0/+XAucojsOj8KIA2rbTVPkYyzPK65TtTsT8JZLWy
3agr04UgX5jIcV2hpCUFAEuGMZlwYzqb940QXEVOuAKQs4SNrPjhOYgkCOxO6y9d
bM9sLcbKWsy6g98/rEConIT2ggcrCJi91MiUol5vMX0AYk3w0r/XFQpzp00FtGKB
cDstoS2r9gQiVtDSajefmjtxaRanSsIhYG+hB3c47IdLGOZOVzwVpavmi5wlLro3
BUjRPM9jPH4V11WZWk2ZM+BiFEogUbM5hDS2HO+KgLADg4CqGqAq6lCNu2lQNpgE
LeCgaZZUj5lJbIvC2d3tzz3FFIsJgjM7jXehurVpQ0ojHJDAYYZBxHxpMIXfoobM
PsnYco9cSZ4inTNKLAfuWHFeMKlWabPITzK6dQSNKs4p4gJujTwEvd7VgVbyWFkf
fTPXIt6k2Q/9p+GqT4W99maacj+/SIEdr1cfRHz3lTxbI9MA1uB4Y+/+ENJhNUCQ
bGpxrmjfL4qBX2sUX4d0KqJfYQRrPUWsx4SlrDVHsYTdTMiawU/FGUgK9spKDSAh
Pocno5QntR9fjBPWP5H/zTqjPtxCapL+eFK+71ryOUwn3MLuI4e0H+oeCWdDEqKI
9dBCADowNuAQ6FzRa/16JExx2dEc3ww2MVK04nhAp950E/kSEbM613O3n9OEmBuP
cJzObSoSUipsH66DAyXnIPy+P/yQJyXqI+DeHUWmWEKh31JKgmTGcRAVVmE9wy+M
CXdFLzn0Y1cie8L80ZgPm7RqyFDd3gQEm0whYBYNvv0lcziUmqm2grHoNe2BnGZy
7r90x9UziawUhLaecaARkv8beEPm3lSjpePk9pN6yVv1QUuMBaiZ8tefPXJ1JPW1
gFgfv+gANeKNfLAIuLLXKRhOtQk+UtSnPSTrQKruo+tgL5iTYdhHVnvUanPZTSXv
YgsSLEZ/WQUs6RhvtUcngjpkOdKN2pmdOEkbbwl7idlU9PyKV7HmbV4WsqdgStDe
0emBomT6Sbz/4YKbIJnbvTFw9JLhubneezJvXak3x/BKQm3RUPfN3MAPOwkZ247Q
0sS1IXdIO6yyEYUOmeDGTRTsq7VNujpswnP9BARGkpnsoUijj1ZghyHrJp3pXs44
c+TYpuOvaLORkCfKRpuoTL4qC+KlmWg+i+QjWxjvhafIknpNqSzT7/KaSfLC4Klj
ttsycEvzpvCOfPNmgGu8/Y6u/nq/3r6vAm3O/FYGtDZVzpmHUA1SSSFMTuGeiSQ8
g05j5QUWRGdsz0qQpY5Su6srFfmvq+nQNasxzgmUqbADexHgtlj7E/8DE4g2LJRM
q8T6+qVuHkPvkPVkVVbqPnIoX4hyJYFGIATVD9EDEzB4/W0V03006ahDdaEOeDJn
iIMBEmWc8wUA9DHVnWiuRIsAB97opoTxkTg7bECNPSdF2/NxeUnJdHRRMQLomvEM
QsgnvPO1ldj86Elv2PhLrvILacSx5Mx0eAO8Z9hZGpdACnAVYP1dqmohvMxWij46
co5iMFWPpSpv+uvWgyggSKlHEvG8Y2Z6WO0MqBdHue6bAJsWF2MxekXnyKdIXc8j
A4zs5ji4NwOHKLDo6W+N5IUt6FBLoTnL6sYvU5RoF1JfMyFPhWzlkS7RYhBtxDVx
8EPhGxMdPYW9f8hiDuUAMEERgQ5k/6Q2FoZqZazGc3RCR9fm8SawYXIwwNFQIzbM
zBNA/zuIp1dvGxHASxMauEdY6tgSkbMQ/pfSsyQi3Y4P/yPEer2Cc024XDRrm9ud
5i25Df0CH8hZ43Cn/MrfM79XXq4Nrm6gs3DKEBsSCu/4hvrI6Oq90uz2hrXlTI/X
Sar0s2omM++Lt12iWJajQxmO6StPLk7OMuEZdkBPRvqmTCB1zKVXHdStS2VijSAx
ax+Ltmh1b3R/dzaqMh2GkCxoDbadyoEoIyOMODUpYvFlzB4MK+3GlsxnHpoC63Nb
ChuB1OHQzrCecgDpWUSd7eEuRiPawOBNlSvdluRqNHWezXeahZFJ878fVxLeFY/b
/R2zsAbj3kdeAwT99lqBgfeK9KirZLpDCXSVJV4teLHo7jRiTP4xOlK0Ke3fTeeM
PYw2Gii2eRUpgG4JT9IBVZpmIe64gWZUg3rTObPeIo6bRCQ42MHiY6kJ7YB65BbU
LSbqdxjkyknjavsleL4Vk/e4LgGHar0IOAuvy8MvZBmpmUVfrhiP92KBilNrG8Fu
fP+0gIK9HULQMMcNjv2WGZxpiNm+tpF77eXovwmNmFWrN/Jy2ndGApLqPRyMG/Ot
mzGi2wiZHNJGhy7IHcJlnllBBxhQaZnaWxTpcvXY5N3vSMxb4MLO/exgGfXAVGQ4
P+1DecSYe7wVP/9cOzsOI5Mevvn3qVaQ+RcT+6vJcK94G8/JEsQyS2QYMVTZyosJ
0oMEpHYY1ed+p8u+6ecEz4qbJgH4eR5uf4yYR3xcCtY/y15e5CyQTaNiT4PB/A4X
ncSRlF4dmQiTImfLH2LSsAXbiamN4LrzYqDeZUoDxVIDdQbC51BqFYUlC+UfdM7g
O3dvgkBBYFZa0t35agUeNufAal3sltBkA6hqhK2HAaPV0IN9Z5W5bsoZBfyTWp3I
vuxz+/2EeKL4svkFtMS5f3Ie9b6XorIm88rHgd4wiClr7tcVnOmiosn7UCx+RoKm
tdx/G2Zag/aSjpw5p8P42mK7ER/7g1Dfp2CITkWCNzPEhbCn8IYykmaJmR0VsZTy
bxyYUzvkwmO6fTMGnDO0nRgkyXje26ZoH8qK/jOfByMSPz8TDQiRyq3OjJaiG19y
CmOlfh05s93yPmFoY9HRz+FZ4zC4585MIuOAIHuX20bU7oem0L9LOkte9RP994WS
B3DAq6CugDMWuGBCFySaibJR0W3TJpafqyv/GF+grUkTqHpzPnHDGhRUbUaAwMk2
vF3kIr2F/HFl1ybKcKfVRKoJ3VLdWhC0yo6024dRzuUByCEVYwSq0GOP79h/muGM
BqIhPoDFiriLIOQnpp2iwUmXoo3nu1DhN8CKWAR6GeV/YhwbVfM5FxJbwWZcubqv
Q70HnRtOTHXqqCkGjZuaDzThTqqXuf00NsuadZPcmD1HdghoY2l12NAdlEkU1aL9
9lw2mIiiu//PXX3zwUUQ6NZk1Amqk/db540+uuwl+qN0gyE+1bzq7lkLOlMMOBa6
NrsKBCSJ4+HRQL6gT+KHaTQL2kJuNE+1EQ0S/i0ZdGsB0F6WZhh2sGoo/xbUWT9E
EKqGlB7K0QyDw+Fn5IiwUZADYXDmVcCn/qfrIk+BqHvhoo8ODfWlLMyQA3FZkYcf
fdt6z4EkKN6jJfrqdkNOF/y98aJ5jlm50Bu4vcbdoISw7SVvebJ+tP1GTmaO/6rW
v0Q5S4XN+4QINLfO1lVws3dckrmdNPBAaro/JQVt89RClckkgTjSnAduZ1hOlqwY
KnE5p052viBUBwW9vrntentK06Lg0HcXyZymunuN1Cg4kUygHH8Ao/+Ye2m2ThL/
0IS3OIP5eGMhL7t3fTXsF0cVDmFw04as4fHgrUtAc4Fp4UORpFzS9hlk5Dnrtm9v
2XecnoH3KdwhXtvc4DGwfX51CEcvjlsxpUunTbl/0ZV/giFAH4s6zoCowX9++2fK
yKQnu0CU3Is/COfc44QJUkDl+76EAt8fGBXST/AhiA1/z/W3DiFcHK4RXHU5nOWr
M18HGf6ZcXy303dthVN8c+GJU4tJKD4cnPXJzCVSf4kgKlVLQFMT9x7+gU4Ix467
Vz/jNYIOEZL/wRInUI1vfqqTVuzPgBFvm+umxhcLPnZcfLW1XS+LCuXYUKcdKx9t
Dc7nOaXPnVIw2W7HBFbO/DMGYhNwySlycVYdgq1aahCsS5hTL8KHfBO5E5rFMJir
BRDwWjwZP3H9gjP01+FKqcSMLk1IRf2LH0wovKo5fwiJ3/9CJ4dN8ibG2rh+mhZo
Y2uom1Wky/I2HFLaPrHe2m0iH6oZSXdJ0iaQ2xHchvDMoxGpBZ31SoyrYPsUJdGj
BEuP25AdSjhybC0/2UIZ7VDpmGBKvJRo2ICuN8KN7jVZvkMkM3h0IhrcKN80nadd
dhYS+N8M8Uz71t1N5mP4cvIVvZ2O4oCjQzo0U5cM+b2DdtKpmTD3c+eOyFhUvPUZ
idlEmcp0FTpLHnfBumQn3ejqB+Uwg3S3R5tYWeD8C+p8tZXBXf08VL8HoVMfC3eh
HSocVG+50AuxtF3p9hJIIvrILma0eAK4ss4lGt5Pqp4f8yyCerQUo4zGayRmZaIf
uSDpnCr4KUVdP84Ze91UKaVj9uMNxb0GVcXoHtSeDLqXoSjxiHUiKq8GiEv6kWyJ
KJ6CjvXGweIUCD6Jn4JTAmEDrz19Jz6fuS4Dl4ztN0NTNuiWJw3Y2B/4Hj66OIjL
G3hHLkvgsEVuTWy6dsPwG1KlHgYisLxKNFm+1VCSpugI/5d+lVHnL+LV57QXo4Es
4w9iro0WFR+pE6F3RsNA5lZIa7UC8cCNhxvIb917AoOoK8MyJrKRdpqrhhPED59l
Z4+zUBmV2QUvKgIUq2bKwwXAB1WouvMZ0R8O60Vjfrjs027ZglewZgfGkPIbyihW
VBLEp6UEF7Ivqz1K1X2rf1iKln8mpEKoDuNkVM896dv9+MA+t1U44A8YK188WJsH
3QkhG2WdzcugkNVoF52qZlXXTb7MOzsJhzvJVOhFKtxDtXiK84acu/Qkt7MvcLa9
d9an3kj4IPI9fUAMRnpQbe7TjQ3AJgPCLex7rbPaKbV5W/+bX7tvJyCZkAxeoikl
wEVftSFFvd2PON3/4gR7NB2ZK8sNqsSze5qLg+k3djsQsDPQ5XWaAtoEKbkF4P43
NyTggX/RcgKS4AQ7Pcw+QX5TNvCzdcRtecbm1Qgo1OTrAhEhygkoBH++N+AWIs+j
/5dCjHunFxWYIyUZv4qhhrzBficlOSBjTsJyY3F/HKsxtuls57N7OLb8ZygSB9d+
DkRt4+0rK6kaXGXfIf13dazhH/lYvAOZzp6O6Hk/yLxyp7co6o4wQRTet4QsLnMR
6UcZ5f3G9o2BkoXevlaNTiHt+J/dvxlwCcfwQRw27iUj1hlFQBYfICHijXDd+2QF
kVT8QKR8vLYt6mg1JN7ZcYyj1pmKCv5fOQZjPNc4eLrB9oS/6VpcLHBWE2PVjMBn
E3oHhRjE/6bOQVWa/sxg49HyIUeuaxsATAkg1CxyT85mt7rhZ9gGpQ9yCpCSRU/z
r4V0cSKxajMhAoB7bUDWlygOMkbU/xzkdTr0aigxtECVqqcUcJaWe44/yzukb5a7
KPhsVSWh0z24glxjbTDdxd8aq9siIWDbXc4FG+TIC1kE9Xt8baHE1UchxdTMdN77
Uq9jR3jSLiqYRnQqmboP0RYNU6eI8c8ZcXnu6w3PkwvhXHGsCVpqWaSDT6Z4SjHs
Nic48gAgbiGGCG9YviE/6SN7UXaUqQX0SIOrjINkaNeoHYRK5KxcJDjOPp62siMX
kiRtNak9yj352V1X8zx8XHI4rc8r3V8DaLlEYHbzzPQjJoI0Ct2qsBBMakXyNAqQ
pDOQkqta0ZGUP/M10Pd6SeI7e8AGt9+1GBqodZg1119en1mG/2cLPwfNL5nVuYEs
zW+3gPWvGtR6VRR0DW4cmX70FsR1sO5TrYc9jC+I+70DMrxnClf81dwyB3ZWesuq
pu9eDdFU/1sDmoCXGmRXpyLol/2Xzl5n+YHfP5sCL+29JjaDf3RagaN60vLUASbQ
UxSr0eUUT3lLP0o8PKnHSsxQD/kE3q/gW3U/cfW7qu52/FJgvPynG6KHKjmuhhbI
6/qNZR56X55evaSibIESGsZPJjk2gyxAoajk/gvGApllNUY+t58Xs9NzQys4L2UD
1ei2HsjKsx+Aq8y85sIaS7AjLq4TvkbdvPU1uXj4oS3+5mKLqaahzY91rEYzuUU2
IZiQ1GRy8owprMyheBg7Rvjyhu1BQ3zuhsYi0JrSbOYE+tiqFlHi+uJIIE3CwnOp
fJv+sAPFda++/YKlTlwRLa8J99vSfsCJaN8yoM2EttbBUU6GlymSMqMYJxIa7YXr
Vh80L1yOYZbN4nq8UfDI764u0tIkX9EY3FZvcFpOa2xX1eSeuJUGsFmbSxN6g+kJ
Owp/iFg9GQbjkTw9+SICethpfeAJhtGyJlB4VhaHZ/9jTIltrISnc/NBckaLAunq
j/P2Ck2lHnrrMj7uKwlRl5neZ/XRxn70bzA+zhpZVsqJXL/I0vH18mF4nWyH8lml
GfAfnbmRBFbOwHsOhvtrlk3RvosTjoer6WbUJzXDnw7n9Ss0BDWMnt0K+Yy2EIn3
rebdFjEQEyYlm+A7fTtS1PEMD48NLUAekznmlmva24TVANr2SfdPUKlt6o+H48zf
R7KATaKlHh28ESbjSnmlYxvbVJQgYzilaXcjltRLAWfqkV3c14x0EEbPQ0P4+lno
Xfx8DatpqGBcjJJcDBOYobBbUxyt4n7mk/7Th2Uy/Kf3WEgqFWEPc1VGmtxbBxoN
u5gCOwfn0mOmxcOJwS+YtHukxk7HozTaReDfvIO/9qkm+Jvu0ENWNSkVxkTqP1Im
u85b5YMTdWRc5nmH2cYM6f/KzX6V8sWG4wwTPlrCFHeKAum3ZJHuMC8oaFwt4Vls
irBT/kxGCz194NQSc3t7tC3S3fpdn+oTAfC8eyCIYkm+4CXkINzY1TPYj8W8mTE5
i/ZzCsdVyVeq9yTUZ0vXgEWmS7HtXXtX9licrfkh2KqXZxIjUdGagR2OxHO5I+w5
i5GDWP2+b8QNIshqDq+Tk3XdpZBSVFuoEU1E4lMNfXOYnimQ0UB8Saob+N5MCcXY
vYw2A9VhfY9A9u5l197g0agfgzOsX1zVgxdkNZYEz1F1ynzKZ6g4hOTtD7JHeDPk
EWnt3fieC+rzo9wY3Eqclet4xhJFK0FKb2Ae9X1oi00ZpabqWn6LmGFiEmSBXupx
WpWD/mp41EoQXVwEiIbJGP1MNqF6PbUVAQLhwRWnE99bGP9uXK6ueVyzTLs+IywZ
486WYQ6RRjig9mAJ6T3e8KKd5DHEAd+bm5kAd0UBH7wBOVBeNTGmycAiOTO887Wa
zn1Mfz0yWazBryN3Hx1iohVjtpNLBj3yRPQVi6zY1HH+AQEFH9gQskxg68AsKGvI
VAnOCGHmusv7mPDR+7sdfpeXs8zyW1dbs7iz4ZugomEygHj6IleOoEUC4NjLvcK4
+8UZukOpZeFGZVdO8EcPnbBVUeJ/mA0NerlJ974Ihy4qBgkW9gKpi67nyerXdp4z
w807U6O6GsDRgLJuob8mzFp7xms7Xq43T/ygQQXcfbPuj7SbURG+ZbTcRftMZHNr
bTsxrXt/qhjRY2jdLR6fQkgf4a769mcmNzKXYPaXX53Qg9wNcDWPzYNbSXihSut7
hMKto1Qnr/Rd2DL6uaV/ZM0WSjV+p9dSwztmm5HMjl1Ar2UgwrkVjIq2jC9SFJlg
pinhsQu5aecSWT/InQeGS9PDsquu6SMTQKlfeo/elMA4K/vzKgh970V7QgjrGtku
+Ut2bQwH+Rx7oRv8JGMgbdt2vOx7y/Lr7xehd9SIVOcjIOC8CMJk6D5yqxGevN3a
ZdKiFXa9POc3dhOGXHdeNhhqcO7VxFlpBHfHx/EvrlC7irRmrPMUqW7azpdXgCGH
kjf0iuvT2DGb7ei7jqfVr+oDB3dDvuRdRXKN4IptSn59sy0isDMOs/8PUXk1t7jr
6avyxsnbaGdPm6HnDzEKMGf9S9BD3cFreVkd/DpBHoRGsDRsLTkiM3izHNHOA7Kc
IMOrw1Xd+TfVlz15ZCmFtgKXEUeU4eS7mAPZ9qGtvhpBsmo6g6QqiYfI8KwPKUE6
187MhtDbx8qGJe5kkumQLQ7fwp3F/zI7Y5brYtkICIN49KZRoQkHk72Lc2vIsEdb
m55+Bh0irimBnUp7E6/Bn/hduzvEid6DzthgtD6vD0rFoz666THxSp5PZJXWYQrq
QkHtqHFNSLq9cFvIc8QWAXVfqw46+VfDtUTAOI5HzOt8/p4l2BGIDQJ2fK03jx0i
aPknYre8WfyCWHlFzE6mq1aUPO1ov3zFAzFp0qE0t4593d6h68z5FN7RW+V3Xwm6
BfwggLN//VppzF6ycD2hFw8fKnvKQFhh2mdj7QaLWEds2kI4y4mBVVMYLnd68eH+
AF+AVbv/Bqu8mLYj3qF67RZ7XpfWwAUyeotEgFCPdXYzMigve8FacnRkL2BVSJ3Q
QVEaf+BpzkRZ9GtrjB6Du25KNePf6+cAnuXd8LPgc83Egc2yYMiUmmDa6TnKDGLQ
tvDG3kT4+0ZR1TEU3WNGttojqwhli+Q5mjI3rkaqN+OZXfnLFzEY93hhFZgz9Bnb
2ox//sb6nyu6T/S176TfTk4hxpkPN6fa3d0gbP1F70oF6VwF0eXz4mezX49UIi1a
G30re4ySsvkuCD2weniMZR0p8cKvTluoMPZrc0o3e+LlOwYU8OIIWEJzrmkef2Az
BQ+MYmxXfwA5NXstWvmsUjxKQQsKWgiKE6MId1r+2X3muF3kSSRSmZTVje0otrEd
tiQ9d6ItbLb8+JVAark8wuhpSR1z0PcVrGLQtdqnq6oUn7xbFQ71gvtCshPJb1oA
q0PHbXdGe61ATiIM0+j3yiSr0MkYDE354WJiWrdzVf++oanGYrI3omytqpdyhx0W
8uf6AfCmckPHIHf9mv85iL1jtocjBq4nTEwau+gbG3AidRMRQ1TUFXsHL1cnAqBV
SzxbtyBlGf0M4EMSytN1Gqig9d/aKM52pZ+Et//CO1uwFePLvYsH66Qlc834kZC0
RrMTlyuOkE0kxQ0SddEgblyiAnXLP3U57LEnwPN++MqBKtjqJp4C0KCzG1jcH5n2
LIlBTHubVw4s9jfSNkPXjud+dpjfOTTtlMUdYJmyq9yWLTmhcb5SoPKbuF24/HDM
DOUPIuoeJK72Xa4iB19hu9DQuLH+kLJBjPnhe9VSk25LICLU75cgNPKnyg8MDlhu
KZ0D30rUhTzFDHTCbTTF6ydAYjsfR8MH02haORAAdn/sZwEKbvpNpUHTlqYh+cdB
kbDsWpxjdQ8P8K2vPTi/vnB37Pk3EJsr/G8671uZQE6FNaMpOpYSx/zv69tDTpOM
8hLwLGS7P9RUVZsZaqfBKuAYGtK9GEkU5lXbG5ygCgAORTm/jMcPFbVkhX1pcSye
5KpOBR+lKSCnFHseuzWdzQhEOhugzugM1kZO7yZg43lJa832ciAYLpnBvZZ7tGp+
z/6q55WWhJaWSUpZvC1sYRsY9CPpFpW31yhEbuj46MggdEFoTZQQVb1LpGm9u2LT
/B/8jgUjycNW3PdRBjzVd520QF0QxlAA5hPHQZwHg0gyTXId5+f5iElPgv7oJY5R
5Dj5/soV1SzhKoRie6uWl3AmmVoA2fcyFhygACRWWCHuZBO+adz8NQ6YSOyqabi9
6q6HsNw4hmBQbM1rZ9LxwCoQiKSGbLUi7a2iDgISUcD9ndX/9tzromm30a9Tux3q
xu3xVL7Pim0uGgp4R+dk2yTH/SRMQId6Mw0hThYpw620QIJtR1h7/J/6uOrJsD7Y
wIoYllh/nC/MdI8Bj1HOHwsLD3oujeRE91onNEbyoxj0Hrk33IkWYulBUPkh4Rka
rmcu/3TaObMUHONoe8po+0zyGbnt5jC0kZSJN+IUXXGzPYHkB8HZH7FM+lmZTWIW
m/d8rkrKFZ0nsu+7U72torBxvHyNFsqTfyIZKZDHe5M1EIxp8swK+9vnGIB5z8vC
jl6ySxREbCElQl8h3f4N8CMEd3bvEDBZjCsFb9ydiD9RTglcraQ7dZtR9nwZDbBK
Zjfz+qvXEewkN1bEkZ1YC80c1ArahHdqRu06UYqwGjyMkyOE7unz0NUagEZD95Z5
qMr6bJsW+Akts+KX78O9j77z0ft7LqjxcxGGK76KX3SSfYgytHKAT9d5MQfwTSGa
o3OIhoxETucnbtZyZgJh+4LjbL5d8tRNiZzmVaS6NXOn4VUUNWuosIfJb+mgwWvU
1sEEcejBbDJxAuKM9feoltRSB6WD7E3uhTCfaSo4dg0u0YLQDHQsgwI0eqqvDRQA
jyICAmFHfpKSr3A+qyRACvHg088vt8jfusosMVhZQrub94dhgVmH+8OPrhjQDFIQ
HH4Y+vM2AEILw6fGbxMAWrVWK2nc/8MCI6TRjU0h6Sgug8Wubt8Z6NPmy+z+HaJP
/Cj6Fr/I9tV+x2b1NGcohnwWl+bwT4bA+/GyGVhVjrqr83fH7cb19eQRz/ihLtxi
rst9YdfrJowWxeNbMn9qdepWzjeuPdnWFmuNzclnENkcmAbqeHwfnsTyHBl4C136
LcuzXywyp9qWxBJkqOGrK98xhDDEe21rMRwdQ8KNi3itRQpgVAvrldHSIUAiFC1Q
/mslEOywtb+nnKQZYn1/i5adn7bL//1V4B3A9AWSsIgRXlvaLbRbMi0lTBsQTvoG
GpHZhmlH/6EOGrBW+ZjJiAVYY6WASOdOU6Yq842BUXocD6CpUyW83tiPn2tDygHN
bygJk2PELMNSjAovsrF1ZeADku09K/vpO4gljl4vdXkMIJ9UaEuSvoO5tgNTO8JS
rVtQLsT6vLAJ7syvg7PXAolSf1Q4D4IZi/uf4m8l7frwPLAWXH9ZpkHvs0XXt577
srJkthtK9jZJaWEaPzLhR3UGArFgtxgrqipPNGUnEwA7wX5v1W0PRcoH4+XnUyRh
EWt1Sw6XsvADowf1U6V1pHzr4FUImI4qecrGyJ8jEK5JfDjQtixcWVBDrjhNlxjo
Bqyx1Z+ukr8kBFSEpM1v4eolJogU6Pnm0MzIwo96g+G/0lToPQkNgRnePHWVkQXQ
Den3sa+Q1UCnhP5WC7UG50ITf7+JsMMwvZJkpy3wamh6V2tcvRYsyx9zHFPEtXSM
ekthyqu4DR4ea9ODEH0arCvVRqZoiqQR/ECo6IWV2eJUBShE7LmW4l5xyOWLMZor
yGB/G9Mn1uMqCfZksDfKhBw95M/AN0cREli+ZApkI3dUbODSmG4wxoWShTlNU5f6
ubQ3/rkzsZTQmFisPhLBPBR85+cRGxtB6hN0KJe8U/sBx5JjhxMaTucgk/tlKlhm
biCAiRgKu3L4dlr+Jm6yqccMnm2SYvEB0bhsN5ER1AGng+5E3XCMNWTXIFl8tvE8
D1VdW5+LPOdUvBS18ICaYt2z+wlOFZJDD2X/RlVJ12mjOju2RxU7Eu6Pk+fRmCEN
jkQxVheX4YULj+PHrkrvVB/kX3YiY5X/wZmtIWl02+XLO3OLNwS0Rlifd8v8AN3y
86Jl2J9bEpkjGJNDvPfcXPVTr33GDHVrH9NH1ygoGeSBvYBdgEMmWeIe5csHeLwu
caXfRNcZw2EdqkO2i31ATmIH1ZbWmPiixtvsXltSr9PYl1ex5RZVFf7ZbvrmERq3
dSvfJEcRy3Cb1VeA8rZMUwzKNVFSZuDQiavg4d08wW7CNxP+wmQKkDDsNeNX9OEI
aPd/fP3MFbd4FQ6aoSV8evOssdYydrhcpcAcfmzkB/dRMmXRrhn203csFrRNHnkT
+bHFut1SoPw+piLrb3hDf2ebRqq0sUqnbOww6jl9hE2CQGKeepDmt6OFn07xUF5O
VEd/GSw4kjRJv3pJzL3Dc0lZQRZY15TqfvEWMG0JJQ7b+KVTCjy+CkynEu8IO2CP
gTNT+KdPkwSvVlLB4KY5kanAXH2oteoqOrua+j/IztW6tqDiWqWIliWXaFHFcxTN
E4kjx0S+tcn7bszovnIGS8kmn+x1ike3zm7IKe76CTmal3e+z9hAjWJSiSnWN8Do
0FjDDIKg6LQhTj/JbfH4seJxI+LtzxQDznJzdaR7rGscB9fZ5CUByhedxAqSfyAk
NR8+kro75UVxMQJvXpY3vCJb5EOCwCh/0ogwppz8uB0oOxmmoHpsy4PlnHTtJ8OW
4OPTHIi7N2CsX8XuMITuvu6wquYM/LGzHYC0sbmYa+hyWGbadIE5PRpjukuLFbpB
VN0BZ+4kLBdGSAMW4RZ1iV+Ov+cWqvBshbW2AZxnLrMAL47lOL6COSTqzePsPTKO
O+t9j8hrwWR3lKbzSfpNfSOEgO1UL1d0W8dVqWDbqq70hxmICJVmpMKkNt9nfob6
PCUUsmkFAbwkh9x05hr3jjwThVbuwa0rV1hNyibkuIjnngyP8FMeSHJPy4IIrWSS
ilLjB4Xq4n2y9WrZzxoXINXeqzG+e5XzaGKmCQBA7Zs19tFTlqo/eRe7CaSESDWH
Sw7ecUmZKiKrcs/FUzpmaDN+dNeC5vtKQ8ZwFLttlN71juwa1pfxnSRUPD9Jzktb
D8tEF3e+nJ3EYW/DeLYOZxyUXFMrI9CxDwV/G6cSm+ssFFkIW9B/tvU4Ud+4NL1A
QQqhh3sDhG96P7vutyq/PRdkE2a8N4Dw+Bz5K18VGTsM61wuiJtazvvx8oKA6W6L
JlrQ59sZZqtDzCmYeKoPyna8NZ8pF2uf2Y9wa03umegH3uyF+GGaoIPft1ZVm6Du
pSFESieBFaDNWJtN0vp/4LZKbq377CCXB9Q/wr7c2NAGHQtdcH39k6I2WJ1b3Poz
EkrXNxE/zvQl1ykfpRE7LKZDD0x9VE0wU0O1vTFW6oUp9PUZrDQCzIU4KO9O/HP5
kZ8aADwJQo8kE01YtIr/i3TgzdrpColIsKa7AQeEbiu99ZodEOgC64BPOYvzACq6
GiMAryUcS6L37OA+1HAKSnXU0lWyzgmLYWhIe16BwUCDT/GNk9oRhvWOTWsSU+ow
WkVm44anwhSV34Y5MmyQdeKPqT0MoCRbSYFglwnIm0cwa7OE0KC100xScyqJu5nQ
i58krhVAw8JIKleW3dBiz7Tm/pps2Gwugxk5RzJBZnSJe3Lp8K6THKcoAmDrdAoP
vyr8mkzdg82ttncOK++YPn4e81pu6ZRG/MIi+etOoT0B2AhNkbYPrwd7EbRT+5yI
coUkvMxzpsaBR4ULrvZAU5n/aaJxk/1bc1zleAJNGzMWXhw7Y/PSnYNVeHLk0sKZ
1s3+aUOADjXdTM22z6jwjkyfL9MCaqlwUtfGV1eg0PLFPiOMPKiOVYuVFSlRk43r
X6wAeSJimPySGDu++98M1pfkigqAnHRE3lGRgQsrmUDeKTc3+JRAxrhl8f/IjHbZ
a/a64CZvfaFnmwgt+f+rc8sg48AUNp8Is/BQw3sWysdoSaaaUZoXJ9l78TIXY/rI
3ATn8in2hnIkoTeldjmtUl2MGOBHYIo29yR4xFtX8OqMT6JX5nhbmb7ZjZPb7hRi
EKq1aJZIRQxsuROHCW7RJBH9WH6iV6k44dkGfF3fMdOpZJgwuWV5l1POnOiIqQZg
KOQdX8gkq8a/1+ep/wRmCch21Ol/Q7yfQtAiwnh3tsmXR+jrcK5CcMHJ4BphADVO
MP6+PICaeIXCw0olEuMVxAw+WqjODQKnONdt2+UrJ8xn89jdEL1OOYiN67LKaDy1
4cudK6snDi1zCW3495RFkvEo6nKt7+zyXVbFflCFTzHnI+jhX4fFItxFAy/pN/wh
Olvez7A8uscjxYLXCTBeCbA5/eNucvy1MN0qPucUIniLNR7obe6Yd9NDSiC+it/t
x0+aaL7nF6USn5+nB/Rd/RBDD29L6vnOAVqp4aMovTuF7CeaRv51y/+hEP4rQDh9
MZlhQqQZBsmcixmbkBumCNkPRSyjA355euCsHNvaOhw54CJ0EePwgD9kvIZDCNJi
bnMhfF+j5btgWwv1riRU/qD1+cCgMtJl0pASA1mvekhcdNkc0uMMWWyoMDyyIEBv
hJ3ppxPtdwNmqzZv+kUo6ilcmCwiVSHQxP9izjBziB0+keYuZnAVRMhiwRXTQGDr
Y6jFbBNWaCHa4SnrEqpMUD72ZGjdMW1L1O7KKBtjjNU9R3KMhX69kyTzq5sE45Xw
MtgaTmCHNhoh3XhFXDopkK1hHmbdqB3cyZDynEfk/Qh6SiyUnDwm71VC9+rbBCWK
LEwSumvDm3NruD71SUzbEQ3hmVEuYh0mYRXm0kt4IuQSAb1IjJ56nblrnl2EdOCr
drG2Dc7F0Z6R9xElhbCuXY8fMiXFd8SxcIPFoeoqAfmPTkZn3hqG+wdjDeyvZ4Yz
PDM4c5tHa0S02GU5C/V/GfoqhNjlIAjtwmSXo1wv0ntQUTKfdNAXJZ1yPDcL+Lq6
CIZDYbMVzi0VLO/HUdtI3j7OncpkNGW/0O9b6q4QFIc/zGHz2+41Qqireh4YG5/A
cqC5p/qi3xgHi5TDR0dwjhC0J9Pt09lqTn1+/sNh2SI4Svm/t6s3eNy0BiyCij3v
kkMtQjfuvQBSzJx22Bucu/WLaxy3rVixdlInNne07HpiAQsOTmYDZxR848GkUJ2V
PRpln5cbArK8jcyGMTkfiyqCcANcAcsohc5px0a8CmyR9OSme782/ywLOlr9VKRm
tL3IpuVF6I2NYkjXJ33qMxh0eJE1qoi93GrdbbuDRUeDTAbKiScL8smO/tB2/H/N
F+/zB1AgYCbqix2H3nDAKhJAxkhYWj5WawRKcAwHU0qbYbVQWV/fizptyGlaNNqL
U6dsW4cMjkdkKClxIYkYZOjkYPBMbwXtXah4bQkwJOHF/diMw1lt0OH5+Ay70OI1
OhKfQamdPOIeq4PRYr+Rr6MaXITDizIFDhE5RzcEeauIChzK880/evQ6rIFPjqvH
3fIxRJRFY6ubOJilNbbjeqdSUE3NB7m3SSJ5tsCBTJuvAYokXUNj8Vx3+nB43esf
ExyKjRsCdfwO/j/QpSen8b0cTF34qu1vyZYkATGB5wgjshg7oMqEd3gGPk5ien3S
8s3iH6gRcCKo1R5J/YTp2Y6r6xW8gu3DCzqASh4hcbJhOFJfZfhyB5d/YDw9bFc/
e9H367XDa+4ir6i4tVNzb+l28+Eq4vH3XRM5feXZQGWNFzHGdtaUJUkvM9Ni6TQj
a2sNQLZAUrnw301IfGtFpOsiphmhlLgDQo51s1IA/M8jnv6Iwg7iO5XkwCg1y1BY
LoqD6YjltoFx14rTFoLLEECwPhMh0nIWu0gMQp2on0BKHZf1XQTJ2B35eHg4/9o5
Yn3CuHXb6M6DbNPAQvoV6AntbHqdNf5M/ZB1sgHCiMAVhH0I8QjVnUrJxJwwnQY+
6xLBLXCCEqZBKNWEqPclqYoYOXAkKKfHgSvHepkXqmDpFPlGFJbJb50K+rn7x96k
fjC6lJZ+h/aNZVsbcpX14ecT9Hd0zQkTur7W5iSfce1grSAEJk3T9bG+1ZZiZxVI
2Tb1FlxkwmANPTmO6CaTCCdkGNPNJC+f53wiNbPst84Uu8Q+N/tPredJ3VJUXXnL
Hbkz+ik0h33evPYFuGaFit/n7rCqQjgEqmwOti9fW1T0HihkjFUlcAd4Cptg/Ulr
kzJrlnED2Ka117sOhQO8Qm8AHWddn0CmKxeI0FMkTvnNjJfm49zy3/c9A4xUr1rR
2EP0e6B1fMArQ0/XxkOTD77sZSxM9aq4pYlIDmH2eMc5M1VtxfvVusTpj0bfCTaR
zBT7x2HFk3P1Upruhkf59FpvgwgOB3FVEmnDbO97K45mxczUqNLw7tVhie+snc+9
+RbBH/kZ6UwU7QMnI04NUTku3RU6cSbHNNHpv7NZWe0EVv7mA8rCHmDpAjM57BoU
juhzmelu0uI9cKsadV0dxvqLZEYSMfUAEPWjrteJsTO3fICllIJIrHAu4Ywap20t
zwMPYVNDe4m5YKBd8qgbK9LtHXliqeCgyMtnOd61DhjUfi4RjqAFYNQvuRp980tp
hWg+WmXxdN8RRiggHcBBy6cJjmQBQRO/dqfIIM6mzRajuRLqPBEkmEIVRvQOf1Vb
7qXFvdqO4JqVQfLmEv9/UknZgvCqetfzTgmHqRgz0RiIQ7n9+vT5mhB584ToG5Pc
iKycaZyVt4/aPs4hB6/LZAPI+vCqQKKaRCA3xTrgUDE0x+GWTagGT/qHJU3J4dW5
YOz5qbkK7us0399dc6W41ICqPehdpSszwtyjh2D1jClZa5OODSZgdmw8ko3ffsJn
8RDdi5cRV0ni00Wb+O5pwpuPQNukNGAixPos9I6cigGfum7MVLVIh4FzAzj97xqX
fbZ5l9WZmryjvjOi6XXc/t3hOsWUIPDgZkf3VMkwjwIlm4HcDwEGXBWVgSDcSLDU
yfM0y5PmwqwWaVUw4lEwbsaVX8N1aRvtvtJEouqDbyIQnNvP4pXlxLZt9qUtWsmU
urXSvGg4HtUaGunffd1ygje2mupp7w2KcrTchoQEU7MiiTBb8+eb/8ObWtGAKHTs
C8sdUubU5F2IayTWvNugrzt8RvA54+ZX0Q2fyg6yhVPtF4TWKBOoEAD3Vdt3FE+V
hiSsbzOrVzs4mCOitVMERU6JtBlrikbMkGB01gwrRK2DZjVpaq6Dj7Hsw7nlLekl
zCKZKqIq1ev7iWa97wWsghdwEH6lFQiuy772I5w8EQ83YGMWMULFviMtqLoxSYhV
FrwqGASwV6O1XliOAAFmFZbFCBg0ETsnN475kbPDeJZZ2faBJAiBg039aekDrvQ5
Aowg65QSzGdt9QO7fAX2dTnf2Y3S0LQ+/TyHRKYcwIsX5u7qGMxVx4toZvKp6ZLU
4dKj2aVms2P49cc0ygsxf+ScQecbKRJSD4Da9FFHPmiSWXBEYQyAFj7jjfztqChe
5MSH2dcmJJ3QLHgEUs/LtmjuDr32LjFvyM61Cd+26WbyVe+FNl58hcJ/TBjuI8br
jbNKgKY6BkTD/v7l4vzStUsRMDhYD12DUicxZ0jxkc/y5G1HFnXanLMWkLSf6dw7
NfYJ7PhnZCCmEC2HMfPwAPtdvO2td6kXtkCCAyvxNR3RKbeFPwZsJ8IL31w3GAT5
oNmR/QehGwVB1jyW2wdbegL4GjobwCznkKNQIGubxkzVR2AHoOvZFabmjXQgXlad
qfbZS0n1rtr3dqtFXcjy4l4LCTr+d+J/4u+hg39UOPePdNDwF9jVSiTsUWDb2TxC
+A36/+yjMu9NvcunjCTGpOeTKJ0VlF5dhJ07mqMmcPxOJtjfc9CxYTknhtx2y8qQ
sIpVWriX8XQEPHm/WunWxEOf7l4ST87Ev2WvSKf1eaqVHpPv8z3oOo1Rymju/66d
8UyZ+vr/tm/DFX4wvNKT1l0VzSq2CSyYd07nK+oeAnbVbseW/IZtUHK+0iL6ru7x
gCwlIpKtRth4fXGBCl5vHu6SHIz/KgdS/I0TDND5LiuiyvJ96zzpbXYCiknaf3lQ
ENCYjuTs2PggcZPGKUhfWqPQ22OHElNmlDHDRM4BTtRWLtKMmZzX6gX0DT0s+CtL
70bkr34LH/IcsGDVSf9pfHo5njju8GYNm0KtpUyOynST6hA7NwOkGWQrMxrUIXSB
7dw/OjEjCCYvRy9KIFGSxNWvxUnizV4CtmtCqRyMUo8So/AtHg1+H9XjCSlPrC2A
0JD+ZtOIZ7RVTwussVgRe7ltGsNn3rLZXVitGUpj8zDhv0STqWCd5xxkhRRDZVZo
k0u0JxmtLOl03tVHE3vbDobpN9MjItqgq+l/QSOQ2DHPz+CIZpF3kH8n70ZWl5jv
S7QMV/NJmrKkFJPMMnJoj8p2g2De/qoR05rOPY4FRRrZo3J+KHpjbwhdipMBKtvF
D0Qdb1BqBYzPM10Ylw2auo+hr22RVjWtwEnfmFr7e2dq3HJxPmu8TnbenLW6Cslq
zVWks/o+ILXWgm9sCoqkp8EsoUrezM6WlOIOfKQThOf5M8vzJdGD0LYFpxnZB4B2
NpJijSRwTYuB0zgCDdCRXi6l/iVzvwAtQcluS/p7SMTK6GqYiA7orHG8J7bWWLup
SK8IheP3QDjLfh3Pa6DCawNmvnmsASB53nsygrdwZSgqzwXCr64283rWPEFqRHYl
BeOmIOtRKPRVZP0Eqczw+/02pWDeLlvFyMIoZtuwomwItFW/uEssvP5fYhsJaCAv
9C1zJXtiAbLwnjSEl4+fqaqzkoA/gplSd/745Pxjb9uqqDeaSymAvX9qTr4rsMtf
BnFLXo/fGHsv/MHQqqf5RoEBwKA5DZcZsHJR1l16iVOq3wsNOj936j9Lg75caMN/
gDPWDw2haYMbBjCF93hGTIH3nSWU6wyF/qmXN2DHlGYuHdPxXKtM0EKTQQcCjWL6
CfgiBrf0qyvXGXGa6z8968ryB/mXU2OaDroAaIHf/KMQCFvIM7V2xF7FkgzYAzHx
4FCX+NqYipRrxfwqQHpRNhP0I68g5fVeRdnRegllRcpV7aG6X4/0ny5gemYof4E5
QkJHtpX/h+j+3+6vT6nPE3pFuJfNn24JVdFinIm7YDqhWQvQj+Bj7H3fyy6HFVFO
6dU+91f3yX0+Fbse1bZPywjF26zhBmGvlYiiMTlcz8pwykRQG27daQT+kE96wzeJ
AKiyFxwmFwGYnDLZzotV/JUWupUMPhK4NqsURaHKlNipheu7JWwFtEWGGLoesqxI
gtj5giEH5LHhKLcuimW3L9Rn4xF9vb96eS29F4oFN6BO22tOsLAiO+IjQxHK7+k+
cSXQl+QxxDvJTgPRAHjQyiv5wgmslw9FQJeGk8wqDUO19hHmbSFnTnN59GukFWqH
V+bIoXjtFvM45rkF3ngAs/y0KIp48FdB43wJIQRaOcsLrfYNQzUdezP2N/mbuLZQ
McbaijmVrr8BsGd9zhm6iHoE5Ms5YHR8EunYk4dCMBCaLkORM73xqnzUtmRyCsP4
MDfdZRfSqhF+8LNsAPlA/GvjBtLblKYLSQOmHOLgZnayKjhj987FqtRnYojTZSgd
yGpzm8rcmqVUdX4VPu72JRS6zGKkvWX4eLffrzChqwKdOmFObidPcYY21+eR2NcN
3pLuKghM/yKlZdumjad2EAAPpP5Wwq5c7Hb3mUAqx3nSbL8KjUf8BUUMz4EieUYU
u15QZTTLgs7yjVxVlg6WtR7ttOKnby3U7YYXd4NLmlaLpXo1ziYKMoK6/MK9EmVS
p+ijZinY06djT+q4hJdpV5Ewc8dkz0wB1Dw10EIH1Y5gpE/FtQJUgDGl4KViBrTB
1NkASlJ7lFiJk6f5thMGnZOzJTvSQgPKkYy9bzziMqSftivTMyVs8j8b+nnD5Wc5
Va/lip57w5aIdUuq2YaB7/hINYzuGWcpD22KtDH1v6nUcQoUyuPJFrWP1hJFwj5F
WKrEOih5eIImZA76mEM88uh4imbkIPOn+d5I5NKtXCn5D5h3WVyTTuzaTI89nF8x
ADHveyP4qjSfSeyQ3Y9gyGenZSCHGcKdAQ1jdVYWtbbR4JvtPm2KT1RcitaqcT5x
UJ3fRGpQ65QFJIFoEWa9tJM+lA449x8pIs049a50m4cvPEgSaOWmic6oYu7vF6TW
INXvKCAsIP8t1n47UKw+VIv6bq+GaIRisGuwRD9h8Ub44wFanyuHPaGoFDQEYhVA
DghqfSENu9yVp0sxeBujGQtTX4jw66w5Zq8AJet7WT5vwpYm5mVUp74MmNca5rtg
5Z/gsWbwTjMn/sSQbiRuIC3B8GhraoxXadLY5chICDfSNOj/pVsX/5djrYGm8jFP
Le3l/STm02V2MacisZCrUuF4xyAf1Nkx+Qu0LcielrKI9yd35ixbwpACVplagdWO
Fzb40ku3MCJ6lisSDc886Fmxwz0uWE1Yj201zvU+ODNmMoQQD4JXmUlqAdr/gx18
lPrY1ZLwQGQkj9idNguyY76GXaRz8R6KNFj2D2BKa/javyqui5Ttl0mRII3vH6Xw
TisQHs0YOHTNamlicXnhAArShGX8H39OywgpS+6e2g/aRzQU0Va+6P+tlKbU1Hoq
C+2cJmIU02HT98+Bp27zgsifrsCoV/fTyBAvkxDTOLst9uti5YJMJH+JcwuK+pi/
gue5Cb1w58bIhzN57zGk4tsXFt3Cr0vzreBIDIX9zVQ+i4pAxL+znhPBVX+nx9wl
sty2koXO/f4KtjLEgYFufaP0JTIUCJCzZ8d0M0G9QdQXa4O+oPIQAo6f8LtwMXS/
QSKf+nDlmC5AHR+JBoomYbbFkU/g4IJQT2TW/I4i6n9/s/IriAAdM8XDrNGbLWIf
43PrgDpOU/sluDvfNtv39ZW+hyy+Yur6BKrkFkR3r1ZE22PXvEoHgkO+xzNGBJGE
msFyK/HS9T1mbgmllPmsc9wheUZlqodTdnZT5aMoEg9ZDDNiW0TEsEhEMajznSb2
NtvgPjTn4+IxC0gnCMazEGAsmSWJCMldZjy/8huk2bowJNI/Zltmsez0uZdxrOoe
UaayoHvjnCYLHwe2GkHsdkvzeC57vFtXk4hzk2m+X+Svra087mUjuF1mHz3RHL4g
ytMq3oaFOChqxSrTUvx+9CoMYXvjrnbIBEUcHMx03+za4Q8gBpTzVQEA+B3IXBLf
ul5KrsOVLm9mX1x6B9mL3KW6kPG3RtJhBVUNT/9LpGZd9t05LhIX/m9anWHEeJIJ
dapoHnJ5TCNrMM8TysbBRMoEHtiZL7AIx1AKJxhcxWuevTAkyOiyIgPXKpLQIfJN
0xbvh1VlGQoHrivASIwpPtX8f+hdPumsbHJywkx8wZs8fxe8LYXw5gW8c7/wNnyZ
S76jLhzMV9SkLMRzdNJqc7LnVTk0VI1AHNJztCqM2+4tA2jCf5x27LKqdYXNpXvU
a9d32Lzr0Y9Cb06KsA+08msCZRV1wDGad9sjMS+hldccfcomQ0hnE/UQJXkjBBEt
/zg0NI3rEWiaJ8oN35/Uprybx+LuZaBeX6tKH7mTg0fbiH9Y0ZBBCUIDzeNbl17/
+4nVMLArbXKPl9zi+2GEtfHuav7/FgGQPLJ5T2zQmklUYOTTaUKdx0a1z8Pn1lTh
ZNH8OYmhbbYFVCcnTqTdT1vLixs6scYjXmsYFEBFZG2stm5dUqnJsCzIIWYD6tlV
e5rKR8wo6vLBO+u3skaECgj/J3NdfpAdSPnXYV30719kKi2vFTFpW4vMtvg2wRVI
JTuIgwdhQBQbf82dHLSEnvLY+RI4lxBTufCuicf9xpTm4p/5SAxe9LOzqwtsfQtR
4IwtiZ7AjH+dFyiBBjQ8r6StatyI1C0v2OwZryCMaxLj1J3WndurVcmfuv92nvYP
StScHNfph0mZqarzX4ED5/fmK5jM3Y2r4zvkKKhHMI/u9cLAUXpHMOp2DMUOe6Uz
98gH3MOJdKnun0XxtByMQ2T/dbUYrOKbI/ZthfB1h57/i0DMNA3FsUdhS/QxmJ+K
kgUcna3ibNBQx4eI0j9zBj8/2sTRgXdp5bsxo8j2YWwCOgGpu7Ii5NVtAxExnYEW
VhyTDT+nQ9PXjSs6P6UOmL2IsX2MC5RAS+1c+ZAIE2BG6DlBnBr2ntZPhFIi2zlE
77TNzLwGPAout6wQGqSa4wOiAkjm37IGlch9O0nDukVDnbKqZ8LLryBLq/ay2RwP
qd4Cg+avQsqNepWbMgEMzLsF+80FGQchTmz5vlxkM1fY/uTe8oiE4fLpTv+gOHwV
tJ3BANlW2ckr+/q0yqLpM2tppEHUUK556fI2LwO5Hv7sVjrjFQPeNvUD/gE95eC0
eX0SCraslQDNDiu8kxHG2VtBB6nL8VGwEdYdw/VQrGcnrOAnZZT3AdMDh+6xEETp
qN8aaq3HaeSPFdUK8TdaYgLV3aupdNpR/kqdI4hMtUExKZuF1m8fZUkCWAQ0hYS6
aPb4doKKTeTMapQ7arpB/TL+kATTNVUJOpyroAtrHjPW/PcEbfYh1CbQEmFUCoNv
CjIrpVNFIS1Nz1KYtu8JGbH1Eh51XyiKBoHyC5/CgspAQS9farXEVWE3RYLGV3AR
zlufwiLd0gtRCFTRlplzLsoMMVN58TVNfZlDLCxkx631QNCIV4O51ZMNcxLO3J+k
pU3KaWvlMdl2GiPRBxyJldoteu4IkSe5k+eEtb/CsHHfjcthB+Dbku3HIMvEetUZ
8EWVYESPD0upLLGz6VHZjb3VwXK4v1ayp2vLJmIdhxQaxrok0Lwsf6z+qd6ZfOjb
E9caTd7fxW3zRJiTDH5qYYvgQWMI+uMOqETnyxOaH5IzgiFWGnhyBZKjbThhq4XA
Tp/TjeRna6Qrq0HPpd9yE3ne4dykY5ErESUe/qUopxZezYDVSIldybAwt5+ckd1I
yjxKyqztmw5Uzexk7k1183iTrpMerj/xVslsxQJP6fd5She2s1bj3TxC6gNteHqp
rR+7HkAT15qu2gYKJrNlE/KNNvCltgwGK3StJx9R8W5yV4fysS0EhvElZ2oMPcaz
7oPmJhXXW4C/pexcRHusxRElhh/i6u6J/mkumKpT/Kg30ceESCgAS1Ixfkc5gpQP
ycsFsOzofz1tESS9AKRkg/8arGZ2FmBXvtxaZabFrzbETgva3QBaV+v1yiqMXvyl
wVr887ohYQMnbSwWX4Mex2MGIbhAi/GcsC4MHvmMrUDZyMrLBaaKN7asgg8f9i0o
oG+rMokWA8J++d3yx/qSpp08MAMtcX/LIjhnJVyJ5xXAC/A5q73aVmwGInT0CDvO
O6JVvqq0XjiwQM4kkkharhuvZN6H0OCTSDBbQISQgPWIo5AZLg9aCfHKwHkqRsm3
ReKp3bJuEyTElr/wQBGTHCmIMkwyWREJDOBK6CQtMz3cvQSK/p2MvhKytHF1Eoqp
unqJmyoinmuz5gmPvGbYwl+ElOpXHyr3cqMdOf4bq2yVsr9VpZSf9vgsjyqKlAXA
ysz9eUT8lrav1yX4mC3suJ5u3/7MXOobKhLCQNj3eDIgD7PX/MfnOs0TCsZBLuPx
nyazR9BTEz5KgT5MTCk243sN07Eakq0AwjD1zzO7tDRXWAgsz2o2AWjVMWRL/plG
8NmSYtyF+hu/GGOcorCfUJZ3Riz4mAUHGc6SooJor7FYAvbz3xZ9ZmNqwxP61BYU
0iH0qeCeKqTqEqZJGM5hnx+MkUourJsOowZh7IKRKLa9OkymnXE/TPeEC0r0NZ1/
7pedEjV8r2D7iRZg+/9WNLvLUGrdpPGD7tJhrtEXCV01lTZkqVqX/gp/b0vUMh2y
elf9NqX4fc+h2SlbGUVi9eTh/JOGwWqluK8EVuRJZaig+Zyqmd5BtbUZDwgdyP04
RZnJ2Ws7UIs3kyzcLsv95+pKt9B30eYCTfqmFidcdp+a+MRBKsjiSiQ+StH3RLGr
fyMP4bqsUzHo/uyW6x4bJ1H7ZfGTziI+nt2g0PnB+pZjwCEJ4Us9egiYk4qmeOTy
yh83YA6YEcNO6R7pJhtV7lu0pYwFetLcwYsye5owGS8CV4vgzDarMssJqlRx2m99
IfK8pgQPXjiW12duUTx4wzO9CQOme5t8NLgKQ1hzs3Ez77yZC7Edl0bC08bqnumN
UTqRuqo8isUfFYxz7Ir4HEeEV6YwjEKHNz9mbnaZNiKeRiyPqbbkjcLNSSzZ0Fua
9UEhpBHD1H6htO6uf4K1Njv9x8uHfbhiyfnTnWHGdHbRcuquob+3x2KxgcUH5XUB
y0AOQmqN+3Uj75s6AOl/HQ2mrZpCyNtK3P366OH7IidkuTX3oibjfHVJmf1qRqEQ
YEjb7Q4LA4VLyhFPsvyC6W46OENrjXDRlpGrXES6SSMBMVVvwcxw3eHfsjFTvlJ9
CyXz7LpUFH+V5Eu8Iio8gUutb9FRS8l1vRhoCtv/Ka3V8t9Ptx1vGL52wKnJBN51
8GPJVP3WFkWbuCmCsya1r9qoG3fJc2romdliuvQ844NSTtewchqmSURioynQH2Hi
sQpFq09BMXqRQnxN9FW9sQW2O502ZQnEArixlT0gK19Qorh0XtlvKFORpFsmkDqf
7qL8T3V2K9n0XUKKuQQUvy3GdJZcTsna9yjpYNyAN2oOSFoNG8yQ1VqnS26fdizC
+szzx2IyJGH84FioWxlzVihH+1jxJ9SvwE75s/4w76AKWVVzfn/tVQLeOJRrByP3
m1kuaWNWs1WEXEtwaxGA7i4xVFWtMvPZhAMLGKrri+qVtYFlbYu0qQdOLEFM+7oB
09yJ905ub6880pqP7N49aYec9pkOObNq0fzYeyd/dqJwF8LnvZCSv/Q9Rr1u17Oe
ikZsRbzGPd2cUFQ+fUKOQMHLSeAsOj7XWEU+FuK9aDdlsVn4gS8XhHPUXxkBmsJa
ykGiCP0hM0avGzKriHYI97t4kv27ruE9ozymCh2P9E3SbOpHb8A917nVLzuzNbLS
zxLd/iWBHbg2kRTtdeQ/uGQQHCtMIU1lWmxOXe/GgkzNSq+Hg4nGUEGYmfCrIHO4
ZAs+nJzMdR0WRmeOxNa5Xb7fTixkqkt4skY3rFoVlqsbWdv8dkYLlpOjRIvG2lmY
Du3bbpKzjUAF3yJXO00IvJkI6a0fB4Ut6QT9fz84mh07mXztmwqj/5DmNvMdy5lM
0L+9aqFhPiNcRmrr0uH2GjP5NASHAzYQkjOlVKvCfuuXQuMAk4SqTM3F667CgWiB
ZI+U5vOjZ6KOvZwmcw2T8X67PIL6lT7drPAiqhh00nLyyt9fn0RW0UxelSdAsNEK
VmianHWoWU6h0Cv6kJmBU/Y1j2c6Rxx6GN48dRDKXtqMMjO0GL9stHWjPcLT/Qva
Z8BF4IUU8omNg5azHawW3wT5y6tuFaZnWGnXO2CDSy7Ztu+617wJv6zMKd4jIGhY
cBxBOQLEDNUjMjK2Wqo1hGvxA7mj85CjQznnQ54e+ZpgR3fz2UDBDjarqxX1hdzR
gEZOBHbX2HqORpqRVf1ht/sY6gWL7fz9l02vdBVwG3/O82A/vdghA+FZtpUcE8x+
PLfxkXysmzOs4RkShrrU9oZomawZnHLxcJ3+0uXyPB/46irv+DlV894MRrK032pp
7fwYc0mUT+nSryr6MxF2xWJHM624qOmmWmLo95aw458izEEzEnvcAVp8T+Wi2CEP
PuQRIHCZCYEFjFYDI3o7nAeuC0oAD+HnMdat1QhKnjPEhi6uT6iSbimfCQo9/hq0
dkZ5KzKne54HbU4wWINCh3z9egRyJn1THjSgbkodngU4IerEGEEsZ7T+unAGuVoC
eXm54E6hQXtRQgH6eLjOfya6ALm6+hJKpkUQXOUL+8sWfRZkGRjeaqq3T1VqMbdr
RroTR4+c22LFObJwib+gS2ej2tsYoZIjTTu/eK6wsO969AZkZREejcOjrhl3M7LQ
RjBs9BZskTzhHEIJflnBuVRHoH2pRe/hB4qTsqhDt7s628H5dPu/exqMnm/AZLFC
z6gbLZ18BL5oE4024qGEa90GBOkT++vEtAdgax13uDhuT2TBd63h86gyUFEZbqzz
f+sA2L9i190uzMZ1rIzU/VYl12Om4A4dFx+ZMvtXzTQdURxz1gLIzFlELiP5AAEF
E8zXlkKUkFToElFfN5X5SockUtnzgYNHLetMR6f5BeGBhce5woLmtpeeRRndTOEJ
PUxfYRj7RE077JvCMaNLoiAMydJrdK3dCLolRmNfKPE0wil8ZPw14h9XUUYlRifV
mABntfMTn+84uaomS/9JU7uaM2ILvbBpLmaioX54chyHSYnjWtnoVUu1L4zAMCpM
IJ8Bvjf6CbyXoDAxtPRuul2fwMcDw4euaOYND8PJW+xkh7ou9Xd8lhX7HW00GloL
uUe2RvizLRCDctvjqne3qEIVcX+mLPqQMbP14pPJPT+mdVvI9RBJXQS6iPIBiE1q
HmblccKNzjPp6MqQBhKd5fDLqpnAIRJ4aKOnIxdN+ScPlXHDA7zIqJIS39Q8+a3T
yCPbAF/GFvqa6eh+JCw3zDMnkvTAC76GzDUsSR6w6OYGQDL401UG6vg2Jv/KhaAR
gFqLIKvceOc1B/TH46rHTB23QJ5R/66utAhJ7GGRXEtfYg0I+I1EjeoEFMwtIaw4
d9274ExtGTfJu4dJEot2noomOlrYlFlRP3pPP+GQBwpdxyUN/LL92Y3JF3k0X5iY
q82xdRj91fQBr2O+PPMVCcwvvP1a9VuCw2XxTVqNTMhOWOcloLAuaxSunLAs+mOQ
SivUUP9jDtWzBCL0WmBYWClkbWsOI0eut30wh88apUTC1fNqBzX7HXrP8q33T+4D
yZc5gtp3omL0LE62y+sj7J0IvHVFQaPlv5jmySL68xMjBB7aELA7jy+kD/T+K684
0O/zLJgsSdk8o3GJpFPjMRlwqA6QN4B4/S+Ev5ZSEmXN86ULj7fAVK+d51Aw9ZQs
Fj/OdJroeue/TpRRHzEcyctdPyXFQ+KdxZIkayhmokEiti2IQfD4N1e4Xs3/BA4R
yyu3rQcdvhaFZ4HFIMVuYeNZfJhd6QES/zCvepXjLdCE+x/uKFuMHq/sp7XMnIiI
bzndf0SHC6FtMk10FLYDlWpVCAyeHDVBSE44zyzmZHBPtw6pbGSdgmu0RLpxJNW5
obTImC6rSEHbGu3vOYN8VGKZTh0MrdPHSdWB+JbtZGmWHtru1DYxIZeahzojgkdP
ngJlv282Z4VwGMEq9Vv/bUoOCz6mg8QhsznCH06KkKRTPc6zdQDod7SybzHWoOo/
InewrbqghgP5KjDpu0V1qQQ0iFEJmkbRc8d5CIGH5RZ6nqKBuG+rKl8nrc/nOR0y
8cwFqDrwzwzT8tVlSiWo0xzyJT4BcFyTrnP6QCezPkl2br8W4PxlGin/limh9lYw
Ttlvv9xoOO8tK91T2lVePiCFNPOM4flvVbpGoUDYtvGRAfAX6ZraL7sQB9DM68Eo
lKE4HV4JSXrQbVXgqaJwlWz2iL9Ig5v9TyHJUBzyqahag2ckSMAdYzsd6owAU9Km
5kf+2AkoS1y1kIMEI+Qq6LWz0O/aXRLbJiR+t95LKox5Jq3gu3WAfYf+AhVQ1Ndl
/2/TXvWxVqPGB7pTMdVpeWSCCMLd/x9ShBg8hycOvJok2Sp7rw0B1MNgMVzpdwWR
sx9K88LPQpHROTDVc3kHROVJdI05qpTO+3hJpk8USH/E91JOAZcr758TyLHbMB5x
rJZxnY7fES7XjiI5HeCL8zYFGjE11b1mqzlTqEYRROSHy3jsCuqd5YZ6icP/Cbfe
CaGmTYU55gPtkY2pVpY3P1oa4Tno3FGHR/GS/Txjxo0uJwlF3EhljznBbLyxwqYj
+RAV0JfWGpPuQYLeTQZGkn+f6IVwL+5jjEnBH6n34C/FHOMeRSMrQbCCS9M8y54L
lZJmCNvG+FsYAyP30plek857QOI8lG1of0DK5s0cViK23YK8vVN6DguibJ6t3gwi
GKx4ImGER9YPFb/bFLkmH8UWmKc6tfvoGqpxVcB0eKMWlJWDcqXPpm+XdmH7kMJA
si9vCjlS9i6p6auFtolnrwWzIoCRb7E0v0mkcDXLR5Zj5gJHRFb9iUzKsgggSP9k
oAhJCgr/s5fFpcDyOvldtEhDZKKhLcvFgJHBlA7xrhdR/m/wFngEXGqy9N20F/HB
Tdtd1pNkEOmM27FHDTW6EsrpJbitk+o9nrdxL0H0lz54NyjmXAuxjYwGQyR3sRrn
tidTtq1tspDgSh3Rv5ZfagK82r25cpCJYnETKRfwZxSUm0NHKSGBnePGZzbpEF3E
+105MdkY1t5A9+3+VXApx4npaWt7EA5fMDApiBnoC7DHNX7fIS2Mqcyct4TIxMjY
M4nUEuSFYy7zjj07HPt09ObHRloyVXxl6XHpvKqH4sMCpZBdIZyp3BDr+qPRVrD4
finWDfZcfRISClHe32PIuFPvbJ04elVYa0cDxZxdM6n3dj4BUZKnxJLpvYeRjVYN
FCkOs3dSNBs7qwFyAzTPmvarxbgr0xLE8lGOAXgTk1W51HeOJfiaeD9fhV0RxDcm
tsGXcwPfTYbGsZpChI2dBDnqailpbFCpaZQgcK+j4gXew0rZj6eO8dNN4d7OugXy
tDmZ4EgBpsbpDaclQZxQb+rZA7MN+0gRl3B0zAsi4i5M3EzVnw7KOY2WVsGNyM/L
aTHL3BXVx20rnLjOLYX6JYSJkpUMYuGrLRQmyuEAvVUBb7fcz5poASctnaY4tOuc
LDd30oDiTQ3pbb7mRNPXbDRe6wv5mgSB9WsOFFmY+zHkNKIwUMMZ3lv+sSWHc2pr
qBM3YaC3S1RFcDLR6bIXM5Tk9iR1a/78LgTRYpJAelIphb2NM4lmNcJxkCdVmN6C
3UdNu4E3P3WR40X4TTw5O1xZx11sMYDYli8sZZcoAlnbOWIlBB7Ud/iWEfxSAcLz
mphCyTzEARsNXGGNor1GTGaZEGDha2y1JqFhCOcm5FzPqMe0S9M3fzj085IvQrzR
wjgGIcuJmg0aOO534JOKSHQgmMFiyEVZlpsUxdy/yZnulML4rDDDb8YdajlZO3Q+
YPunh+XA/SId5/YnSLP3jilP9Eveno2FNqOQmjbj5GueWiRGkc551egQcvCvAiPy
uU73pQ72DGdwF8jaFPigr7IHg5mqP+Ny11SqeonOzTNnODQKeaVlp9v8SO+WaeDV
7B+f8xOnQzcKnJJYXnAGuvb8rjk9ui1zWPHfJZmH5GK7Rk3Pc+N9FC8PY1Uel2ww
6YdOkSjB1ro2s/qtrDRC8FbwjCwdVvrnNCbSZAoUW2jGKzpVNgwL9TSGlVrap8X2
S1TVovyE/81gr2c4AE8kAt/XgS6A2gvkN5mxRSDDl1sUzREi3j9iK6za4elQbLJ/
1QjLWjpF66kGwJczM1RLuIPIUsB1GaVXRIqJT6ZQaBMM9FiQNaGrL1S4PdHKgqL4
yN1oMB9/SeQWCtxglNd/qHd4mtnXcC5/uusVMN+upbcrNhAm69loLYaP+2dM4ojj
mwkhLeTZ5MQz4+BOhpSs0icZp3B1R/QwLBigBZVys1h4OJWzVUk7Odjrk2tUUyWk
CGmyhYOTU8lGYyKAnA6gSzebzpImZYnk1GcVAoZBY3KT1un7PQeHFVWKIpUF0Hye
TltZ2lFn4XcAahMTNtJaoyl4Y9xqptFjEgeIh1r8iVssao51E/34SnRyxCgQRMTD
yq69wD1DwoG7A3db/rySL5hWYZHlxBjXZwGxSGXHkJQYy77N/iWx3DFODcb3H6lK
4zoEpgbDhAQi3uz7MvW/UOK7AuH0g2MSFNll5P35NmW7NdgT3ysjVmTOoqYHxoBe
x2vOxMRsb7VS85eitMjLwxMss1HEqJjp7Hx3RiXZbtOn2VC17881r5I1as7sffM3
QNb21rJSd92rMjGm0a0cRcybNm5MOo/6U+Pwe/LGH/6gWwVEKvI7wkoEZXPI6MT9
67kAPiiTVW8wXYGog+4Ikk6sCa4DMEUJDd031zlM/l6+UgKg8ZuMq/X3HAEf2hJA
azfG5b1p4fc+Rw6nTzeqojTyBAfG28rp9wRoZx7GJEFTruN+HfcCoOIEvHttxF02
aaD+Tr7C6C763ij/RukfaALzrTO3iecu+KFIxg/4WFoHyc6siAdy4d+S/iKioqG4
sfwi4BGFh/z395tZi1btz756opM+nUDkd+cEgURN/hA4N9bnUlQNGM8NDnJ9ieM5
SNEkkO1ugAl/LGuBykM7/U92Ndg1FXuAv6asPirqTzTSpHElmGnw/lyYw3rMIrGK
QMwJBpRQl+U4s1tvEksD5ayxdU8T6loS7tvnZ+BU0rJlRdxAKYixHgsesrgSXxly
dlcZoE2h9ivBOy7LTjc8uslHujxyekxukcmmuAqfQpeOPxnOqALeB504O+jGi0Qg
dweGzNqGbeokqT0+RrNjnGvyAu+NJRx9aUIBceswkAo4T60Cj/ThXHHKkKjX7ueu
kZGTzrkSxMlc3xWjNz17FXk3r3WvP7aPq5qFAS2+GqrxkzvuwNy+/oPcnbECZn6w
QyU8IvwyLItcL3aCESU2+vfoaFfJtFr0Q1F37oxZH/tlsJNuYF9ZytoT2VGADa/Y
MX2E+Un/gVOXOYc586uDgxtaXM+oHqX+ZFbhUUGXwCR7g4wQuu0BwvSisnXIKD5d
VAfpiKotcRpL7kjGTARtgD13NlMEUNC/XDvuNJZ3pO3m+CN7T3MSbvICnT3ganK4
aX55EwNmEcqc5CQvwCNhCT0FjnOxHLtc2ftiDANGWXfjY7lFmxGRJ+1pxZ3poGw8
FoiTaRJBEvnQ3M+tPOq5DMuEItfrB1xUnSBcLBOHDTd4FqK4wVyb6adCilxDw0ia
SJdjr6PtkcFMiZ9GqbdqLm3vawXmKdjn6XQ083JnuC97FQarsDIRbYJAdC4DGsoM
jDvRxTH2TJkzbbJY1iR+n3THiIRlesVk5JC2LPuy1eeYw9xr2rgMDzmhvAfU7cco
gnngqk8clA+cdxkioj7pqY9egS8znp9yxI1zOYwzH7bTNnQl7ClsqInCZqVS/uoE
xRaQFgijwWjwxspL+3jtUmpEx/i3IduGJ31eO5VZBy92GZLOP0fi2u1t5IukANsE
eVZqDq7EcX15eQ5yMDqlbpZeJADVzcbQ2YellwI/Krq6gt+egRx4oFoBgnPEZyxy
GSU93T80W04GGFhsuIBYnd2nACuA3c8HZXfOSEW2ird4ULOJGJanTjVLBYVxpqAq
OqNInHp6LMc6D4RZb0+Vo8XhsBnav6ExVX8HypLyyLM5rRFPgzdg4N/X/MKyykoy
5JBqvCQuib2bQjM4M7FF+HoJwsmunwUKwOIJmpTCPYcYhfbp4KRBHHAIB8TIBQhF
bxYXedJohpllYSUe0n/ttjkxaQFFg54GQAxi1kXD5lGQ9ijD59vZzSFZdWG+5D07
j637jCl3+TlEZKKGBrr1RjtDGl/TZ03pEGhc1OYGCZeh7lb+TOKXmXKkiGFfU2xS
Y2mjTxaeLX0IW9NyXwyiHEaQEIcnPfkzh8EjjI1cqENOWzxpSlUO2yriZye39ENt
nFVqQoPuSOsly2FqvPhwWHSktIttp2XOdI/TboU66l0+K4iPeE27KdrtgFNERkfT
2GiyagMf6/QUNKlMJujrE2LO3SjU/0xnTplfKcHaxcaFN9Pn+aBSM6mgv4YzrEN0
HIkItRtT2QdJO0ilQTU8ZXB2MZRuNaRi+ytfk/A90dosXCpJfTPIofed5a2f4xwy
W5ZVY7MgGOmVS0RgvZB9GAqnXMNadzRWM9j4lNLn6e9WP8cfeBZnAyS/qhKJ2hG7
uDirM8EL3yzKM70eu1TLRdKaBN7mhrUOYwx9R/Tnj03klUXh4gi+1DwpFEIbDgdP
rcZCA78qXeizopzlEFeMXBDuwlg/2v7IbFH9kBks3T2AjPdr/S2DYq84QiWzmOg6
EBaFgS1G1KHtyI1PcSpfWM7TQ351rv7YY2feUsqiurD62WZmsT+ynsFfeiQ6Lteg
mHf1KeA3z5tyOCCbdAUeMdygpVTeqAYMSHhVR03HnWP1G7TK6BbT7o8eFnO/mL8Y
Pe4XoYFNBi5zGALGQ61ygQxjaKCYlquqYp2LEv77+80b42aJN5b7OEOmVUETOzkt
+2pWCwEnythMZ311tcNn4o/QpgmHZg5scfg4c2zRPhhCLG01z14quy3fXHqfIKvx
kH8psTEu4FkR0H4rFHkZDT6aZk6SxMJc0/S0TUx0xArFhn7FgNQEntAmEKKKd2Zt
Mfgxgr0UuRcKpyNjZmy5yDuoQPSr9bbIHsTAqSayYzYgSlu19s3O1boebpcfJ9/w
xmQ1Sqr6ROj+ybN9T2mlgrVunHlIZcDyyuNlbvbzISlMkFjRNbJGdJOArcZv2hYY
bF2TcrTsA8xq55mGv59RfAcd6S8tB+sBhdW1IVPQYGNaQBku1N8k4vO/IvlVcjvy
VIzOiQywOAUpL/snuqVYafcJADoiCiKPxxN0UNFmcXYvLceohQj/Z8SfDp7Mw6EE
k30iYpiIFzXTr4c9xHdyrwlX70ZuFStXWMLaKC5/1H2MxLIa37pF2s4KIjtZUKPw
uOUWm8kWuk9ExiSxyBZKUQQcZDEraAeTDLKccGwCwNLByestvrQx7+4jCyvx5ObS
qGXHL9D4BrERGe95yLlNoZqN5wuLwo4Hr4RsrR48rCg98DURo8D7L0JfI7gFsBlj
ONpnrdntO6sfGj1bpNP/2cdm8lubi87Vqluo/RrDijawGpeIRe6pEqh0Bkg9waGj
lqQ82fjOxFI+TkFxchZmkYI2tPBze/mB+qfKy/Ifv9aU63Idzs8iCxRgkWWzLABt
kRZNLNA7H407p8l/qyHpjWdmsrBKtpHGjS2VvatWBhFW+KXzBOEJew12i2coxG4b
/IYqr8/9m4aXyEbSsLFj/CrG/m2QfMIDjwRKAUXdYHn5cmWPfFsEVKvw7LCAeKG8
IifXpDt9/7C12M2hF+omlosD3m0jPTb0Wj3pB9FfOejg6WDC5PyhExrdokeMBbLC
hLdV+bxDmwcOZiKhTzVkuk9lS9PetdAP/UagFYn1oxteyUdLLm2UW9sMalkvTrvV
slSunTMK4TbUut8CaioU40nK0Jd66IO9gcG/w+XVbAfh/34Rpke5aHPmhISGZg7q
7T/jt3aBT7hYhTFxJYW8vIDVx6SmAB+CBTTfq1KB89+vhqoOgnX90dSV1EYaXlIP
6pWopP+sNi404ZiVoo11Bv7rN3i4Vs/tPNM+OqmhrOsSUZTgQKIUMhQoMGHN/E4S
ZtOP414t92OFm/JldVH88U4OhMjDoZoQNrI/0meOp8iu/dhAWY5xbNu8M3L/c6lD
1KzjSTTTfowQYxIbgdZhfHzyLC9IawdjBw77McI1goWsMU4imEgTUMWNbU0XxsLT
73UqHPheh/crg0YNTuzrKaQRdabTZ5/5ZQdfzS2mAbf7ogfTpqWWH/vsbg7ez58N
CzSEHjwtj3rl4ApAbPmUw7+8jvZ3ZrwYYxdhcypmSDPhrMVIAINsslUkq3/yqY5B
aefuJCsFtJuBepGtBrsLJydFlVlMdc9MSoJ3Rl6E5EXUjjOVvdzQG5VItQO2ffAV
eX0b1GPKwuaP/DovtxA8ZQgfhXFb6PjsG+E4VTR8HDVqB4W8bjtfSbQnNvygB3wQ
6otEgiNm9I+ptuTvVoe4snvL+MvFs44yS6trvCGBEfyV3BzIOXmxt+4AEgW9bCSa
4poRHlV1vELr2b8wcX9OX7vdkEV2yv5cGNUVygS0nUr9EWnZd3ufBeRFr49rMoYy
sAT5P21nme3rM8+ZO0FHDcQBdcMu46FC5P0Y7PoWOBN48ivoK7y3jVpFqTG9NsIi
pzpC/8jeECNGzrpYaj4Gge8E22z0R7PfE8Uu5Y1XuUN1v1uJ1Oyp79+BU4+AaO/r
gko1oabZ8asCRllN+HGz6nb2+ZKw1tb8txwN5jiJ5IZNaT6vP5PncsGObsc8uySY
uAIjY/E/7NwglJcKZJNCrEkaTxqfNVKaUkEVrTS3JYK+hltqBBNN4toReuBnTDb0
XlXXp8qi8JBiiWrc3QsV0Xmm0OOBG5t4gciq7DwStDMZ2ck2PgrzG1jjjurEgJac
XunLZsGkG1DJsIxnNmCWEhOWWXGe4T6KpisCbWIYt4aQOXiYYbQ3brebRRW65NLu
bntiFptzPXdHJUx2F1n/eNllAE/7shHp3ryCFYlRRrXCEzlx+JyIwgJSui2UPFxB
BPnVr716ooaWAAQpy8eZbcYygqCnKEyokJBoblNjBJWjpj7ktLlmDXX/SjY7hhqz
C+PRUFK6xN6APjw0RskkkiUbm1gPzP796k2tmKk28WJ5whT8IapNFf/2JxyATfEQ
Ql1O2g3v61fpLEnVW7wstRbbcI1QTQY+HNyhn+L/1sX4VWxmTGm+YSRQFx0lRREL
qqYAFBNrccAUMQiQG7ZOH5+fbmrY+jKBZKGx2gZL/b7sRHRf75FAucHVAknGhzU/
u+f9GZ4bLqD567ZZxcJV7k2PZZTIDiS2Tb6wb2TZWlOw84fyCwlEe7EAnPMYYYhR
T6QGfzVG/XwSxHzrkjk6d3+2Z/NAz5lg0CMD11Meakjzpv7HsZSMDIERpoZNYatg
YzVq3ePVC53meiVns903TxVGgcQr1/YePnDaC28mCRMGiNhTS6bjsgT3DfH0gXbo
3QbAmgMEAwxKBlJeWUASbNdQSE3/Km0TcG0z24tgOD6Nch9vJ5B5Dbrvwp7V/l9C
DgmacDx1FTXpaZMKBep0w3DO2/vNx/1yNZ1STktPvcd0QI00HNwVltcmWC51r3IG
pN9IzobAq/LiHg7ZlGq+pV+NC0JZqZOt9Kcus5TQwBdu8sW0eQ/gUMyy306Wmcij
5JtKHyzcw/kx34oNUF6pmk1X9YPLpVcdo7xzziUalrR7eMF9oHD+oBb1AAcIUnN9
Y74ln5CzVPyJ8a0u1fjB3NdsKqyZHFWVv0I6hFyxKdFbzsw78RevGBF6VBtgRoiF
1hC2k4K6SaaNfZNlD2WSsW1fRFNk1XqzAkhWPUYX2TQJCQEPcpkor8/7r4ITV3PF
GijOhHJhspcwYVOaWmD/gTRpti7IKgNm7YExh+vCjo/cUywe5jecM2GLZaoPIeJM
JQL23vOxvqKl8RoS+EVlJgwq38Bf4/3Tduo0b2twOGmCc2G0+QOdqMBA+QqH6/au
HI0WOF7JIIMl5g2vnKATrPC/+D2uH/zQjjbPy8WVcJr2q4DkcKuH3TGMR2JtAveR
nxcsJZVgC7PIwxoNUxLpG9VrSgb8xokCjPdKVPG7BuaZ2xuZJca5pfofPWeKOxHF
5NCMTc9sWr2n3iUf6+krsM7ABgd29rljMCPqPHnLN83JXa0A9T+9/Ze3IC01T8Et
LOi3oC2n3YLwthS3GR7BEi5XaBBebl4UChFfG5sQKbMbP7mD2UPj/66hM0NElwg2
0vi8NAHJ0Eq5nG0EQUmNgAJKG4tXZgZlSim8kTUc9Jrn0tYXSUNpRraf2Uu+6Vbo
3+ENjD+S2dpksj0PuiH+mB5cJ5pgH2/JyVNt9OxPWXXAuSZPd0jbOFwAUJK8amZ3
bi6tSX08c4gfmFS4unyZZaHPNqtLj8KC44C1kCbgawrPlF9OxHpGCiNBzcvMLXsM
IW/9Ci8kEm83lNRuu02hLuuV5k/0q+IqHXtD9r5CcjmCaivE8PNqOHubi3mZWvVs
wqccnZCkCpctji2L/4z8Y0m05v8AZGgcQkj6AKBmBdn17GI6dlnMdqu68A9hAmCf
fbmUQ6i3Mk3k67WgEdHJ30AgHcwjeTz0tpvBjsjEKxtWrvzQg1QbYzlaO9Y7IwEX
RshSlGZgxp7EEcNSnz2ooU46L0QCywsxtwhNwQ7yht23aAlQAJZeEhX2OoTSvzbA
EA5XD/870NZicV0U+7VmCDeeH2O0FHbF0PYuH73n8XBxL4aRsZ8T6Upqd0IJJwCo
oTxDrER6CC+UV3wTuu/AfMiCOMLEp1V24O58ok9SVhR2PTM1PCVPBTgQpYwXqCQM
quvAqHj+oIz6wyUQdiEF7UZ47lX30gdVEuEMBkfq5YsGCephke9hO9lbViVYZFj4
8ShojV6UeENw4WSAXkO034cdc4wV2BgL4T4/q6P5qx2C6zp+0G7fUa6/o8FLwiWp
9ffz2o8TNwJYoRUEy8oMeg1xdguWf8oDqDLL7DA10GMb0ea4ZHz3jQRUbtiuedFH
GMitf/q7PMqgKSlR0TJZoKOgG5F4u9spbA3CzLy+X4pGJP0FD3eSDqFhMy0rl8e5
dhe+JPotmE7SdEtHUzN/4LZMJG5+DEWZf1h5k01tS50l+MM+bFIAHF48u8venw6A
5HkEPw4m8bbCeCsWvN1cxBg5OTJQHOjVvrSetKNLuGNmC6jZtjgjGD5dzlgjrDW1
SjNTntSLUb+oAPZSWDPoV0+S0cwAM2fj7umSD5miJVgNUd2pqwaMxloQQYgWzNKd
vCbZR9HZ1YRUbgwQj7cwK0HqrH3Jw1lSbjnfkt1zxAj5Hz71JFQPqeW6Z0tbm12N
l1pegj+VaIKWxuOkinY04B0nAkQkIaJaKAMvdvWjrFy3qkJr++nwFzQ6xz9Ao+W+
FYJ8NM3E01/X8z7wTi7QiDBf8U8Dcb+J+D2YeGA5klWV33aNJkxWh/FynHlMsevF
CnFJpAedppRlBE2K2kAUj+7JoxCdcu/USKoU1uT3d8L5y0OIy+dje7gfytDMYqNs
iBraHplaMZxtjx5SbxQjo4fZBqCv8uZjLd30kr0J8+I+dNHTdQEtafGNW1OHMsPG
jpbgurQaYvNQRqPdZ0Hc3N+p2ZdFK/LBIW7EwuMQ4BC9KXbK5V2W+BRkNg10ydsl
t+KlQ3Jjnm+Bwc16ykvNMGLTrHRFMbfHx08Gosrz0dpo4ce6SxfMoR36NWEZjul0
uEiAAx6daXDh4nOQWg3E6WKEbzZrh/oyTy7eMaMDwyhxoS9oMtFKe8oerpU2iSbK
Ky2mnlwW34gsJGqoGwP3tjo10PZM2yynNftDx98ZY5AoFfCa3dym2Qs+iwzjeUx1
QH6t7SXd6stCjWKyiWibVpjR81vSEUzLIK3joogpzB3t5qziv94EPWa6LupMAm70
f+6QE9eTShKv7Aom82gL3ZL2iH3Rn8qUYFjlTtEV5puS44G1jwONImwrIU5i0UNp
66WJ4VK15l9JQ45A9vPmdxl9npIxGlUQUgT8VAZgjJ4RxROWgQCQ9N1kopuRYTIE
9pe23k5HiW+uJI7FYuvE4TCee5BaNn8u/w+ce4AZPEyJSRQ0nDRwR13lUQHPWV/A
+2K4SfT/td5GUoafOi9R75D9s3zWEvyU32on0t6BMmVQxFeJZTGvEZGM+8vWA5kH
7e3ZR58pWl2LhTnTjYghlJqYPzJgvh+j1217HLzX9vMlEQOFuBtoPcsNr3lkNF+C
wckNIFaOIRzYXGi4/asr/TpIvTWLrpp40ggOzsS9SwNo9whoKYXxvUFzf5pWLbVr
Yq2YTUyft64es2BrQ1v3mSpjsQaFzCuJ98JxP0NdbuG/F2dx+e55f36WsszieoxT
pti2wD9nphNS08o2lHjueryT+nzbGhiouCbtXPcSlNI1QsupbpimHNtZkJTqFXwx
hn1LGmwvXB9a9lLkxXbobMaRM4vBxwR3LWzN5eQjXA57RpK2QgBLARvi48hGDMtr
vcfuor+gXbOVd7adN6J9lzZVHmJY4Yzgl1JQSHbogx8obI0g0OJFxqrGqlcCqGDC
bDB45ZvlvYyf2zGyuiWaXqJlPzSHTIdJIQm4bVprUN4ep6zy3mmGVyBQaRg6VJ0M
5Lww7XHGm29AZsXvG2DnbA2/43ytOEb+eEpd1cgXJ1p0HNaWn7/s0S+8lStpECZF
eV66n65ebY/KqXCmy8oeyTo8lTxEyaOxOYwjVGHnMZolS7i3j9x/VPhXyz+RLjUZ
jjaYLpYgnFqd6IdSlPhIZAbSRUyolDjqU4zif8aZcf7FhzJ2Izp/kqoEfGZjDv2x
DXueqFpmF9GbNFWAJAU22bKQdAouFxx0KDF/kBqy/DBv2W4rsAnsJgZJFVYlqirA
s0364L5jA2O2TBu5AECfAFbk9RBUWh2vsmT4uo9SrNNmWlqSSc8eL/cYsihMXfga
WwL/DafTtaCsA8Tdg0dZWpjqXcEDbXa4b68ZsncsGR8yffrapadFAlW1Fz79PpS0
2tkSpgg0LE01kvdGAVqG3hKgV+QNxGtCjTYHfTJiiIrdsgQMAhvQgUbBD/fl4Hr7
d0GlOP92dd8g37wJsKpXcCHvUkuQN/0MfZycnrv7vB/5khWE3NSWXAKis2GBw/kj
WPmjzFTNFJxephQBfPlxZJSoJUJ9QoVS4zJNKdK6j51rvQFKsYZRac04qMUtBfcJ
aJioSuNnbR0kzSBDeArZYdm+bUfORZaIyC5BLJlaDVP74xrT6hjyFFN+0AhT8soy
YVeIQ05cfT11Owxr5rkRq5LPfPeTotElM14BWxUGPrc+bXD9cyYmwsgZjw5AoiRa
8axBawqL6HNg/Ydj8GOb39E64KBE9mtHD9f4yTThVVr9MnNke6r8bR5+wtRJaldI
b+JT1lYQICpCZ3ttlJADoHMgEMdHUUGYE3tJPSQwZzd+JeWwj0tAbP6UC9OWSfyg
N82rOFWSSpwi99+05Bs2MDBRVXMqvJ+pEHemZdMVfe6PfCrYqRa6puWTWXMQmSjd
JrBhAeM77l/OVcntBkDoSOaUqlzSDI+fBnSudR6R49Qa16AhtbQtx3/inMkZevoq
Iz+QaeWktqYIMeTrTRCGJp1zqT6tH/lJSplCh0uuHqPv6Sfdkc4yr+BdZVS/pbqy
x0h5RD2q+lcMY+OnT7agFruKasu5NApnna3MQVlRGYw7NPZbO21ONguGaYKfR1Y7
kABxf5+yW2quvWAJHOh9aZTwWnmP8ecP2YIwE8thQtX5rOzmZAus9rMnV/ZOs5yP
DdpIGSXsQh0gwmVZXoroEMbRH3vCvbBiBDJGTUmqVWWHZeGbjrVe2ehkEFAOQJiP
yy/b4BnHnWNsEEppyXuc4LJQc8cee0HLP4+JLBlFkt2QUMcZ66Z69dWTMkjGu2rW
nKIOOcKkwuXiO+kw8/gad85fBV32SVXP6sYvMxMfJF+5FDo6emUGcEbqoEAU6nn2
I9l3K+mgpYpb1YCnIh3Zzm4KqC1cw3v0SrNgP2KLjRbmcbNICqWXbz0UN1c2S/Js
Yhkby0DkRb7Ytv/QTOg1EWxijwgPGSxXypqPXzcAUwrUu6A/qeQHxBHlp4S2lCD2
iu4kwY318FFKskRKrGxnm0s1Gs/wgcyNlqYb8cCTOtumuzBHvJDzXItjQfCkExNZ
0EXyCn2QAZ+2Cihj3OtfEQlrMUczd0TIPphjh271g60W6uVW7O5Uzfvyf0bYlICW
S8v7/Q5zWV3Jvg/XZNggH+zcqbO/sxVYguZuqMApfFn1OmHS4J4fskhEGdL2KTGB
RfsbimvVDwrNuP/0vK5Nzdyfpfl4DHm1Qfs0q5bahkTikr/sJWANhxpEzDs3bcpz
AhjNwDv2sk1fPmn3zUlVMeOUlsaIHQmcX2srQB4UOgnfKBaHPVeNydXR9aQf94a6
cQr1OgXrgiCGjtCZf4C//hgkGbsPVVU/pNhiMTCChYOjV1b0o9Yt5Zt9XDWpj9Hz
9oN6eW1tgm+LhDHKwtaP9L6hPJ8WK52IRZH2kBnlpepJNKYCqwiRTP1ZUgbs1zVl
4u7hBoikonGSvPwKNJSLTX0V+iyfYObx2FZ15wssiyS56k8y2i/3Yrm6yA472nps
tDU262EDxS9j11kiv2yftbXEExL3BvIoF8CvjFlrRQZDm88KEppghDAv4+hWckOE
ZZzoIL+vmDreNxs5aEL/Uphr9PCdXcOCyn4RPN2SaUGry26oZgU8Gioy7m93WNUd
NJZGO0w73GtY4brAc4NewglCh8tCu/YaTrHschiR3IQjBuFt7QqbQEVCzMZ4eij0
ER2U01dobhpo5PHapZ/o5x8H1uELGfBjHFn/rOAdai624V1l78sjZ6327DlaLlLa
6VHh8z7531CpB5AWsMfExG5D+vLwVzj6yztaANuVk6UJ+I18nODIIzvT9KxVJIgj
P68FTkmkzZLfM1nNYl37dZFe0fysTg4RyEtzhQvIpNQuDGQSuovqc0z9fvgGwSav
Z85USowKeu3XEz9knwzU3AohaPA54OJY/kElvyLuN98M35d/LHXgDs1BwdN0L9rD
JdYauiEu4nrF1Bp9eJ9KRu6NAl7QsetV+xRepeo8y6T5ZyVuHFn5uyE7VA40N0rg
6t0qcJkokqk9m+th1bB+6giMHdmhs+iVsoOIeR6snfh4W72rvdtLwYY/DO6bia4S
PePWh7pZlyfsQKABX6WBVay0XNtl7QEP1bODyH6vuTmp2Ko0E35xKbp/uZl2tHc6
JHhrtG7Z3gRUzrsFqMN6Bpp27noNEwppKH8Resaxu9do745BJKY6ZH89FtHyCY5v
qGKsfOOhIRdCswUc4t5lcZO3sB6E4flzW6cvj0btWh3lR++bAIKxjdy+BADwleB9
liI+DSfruVlz186RBYPpIicQNMa0DPw1wc+jAAIAZFwdPnE86zbJ1KPbhC2/oHx2
NW8ZhvHAVcnx3oFjbVyO0URLG6fxU5fjYaWh6Z3qftOSPfochRMeLhlEUvXzatpp
Zb8vzKHDJbBm1EQ7zIhHXoeHPuXyz7FSeCtfr3PJXlT3gmhT0DJTitd9ZrXznO8g
kCDIJWX3+PxXiFamRa1y7gj0/E8W8EQHdNAUUOSKCf9j+MYSEquIxcKJfJeBxzpy
6CO2O7/xbcXEKyA8AHSMUfzemHRE7upiJ6lxrqtuAWoEUOJisoeeEUO1LbPOnW/E
OwVCM4PuWW8f4FqcR1NYjmHm+bQ3Xqu1uj/p5In9mG2HKeCIRrR9O38Mh1ypYpbs
K2ijc8ABvtIzukhTs3U8Poy5X2jc9oi9ctvCB31iASRcAA5hsD+GZPJAIifOmWbr
bZt8kBiUxUrfrPgD1O+rcR5lD98xNJzIdudBw8T8PtVatnQCwbMaE/tq1LZzShD8
1YXnw5rjJwUVdwce7gRx4/vut0Gco4w4u6k1FEpauu9C6NCdtbYk468kQFSG09B3
tri0pF9WmwqzxHZskeTQ74ARS9zFD0zqjvfBTU7NHqjGBsDf2gPqlHw6hGo7xgkp
/bUZZFkzAz9BUMZcuwu00MAVGHS9e41bw4lHakvY3lPTFbZ9l7ftp4pXNLI34iaZ
u4BcMZyhTB2rrfi/8buE7QFtWti3cwlOeKXO3Zf9A/9BYIxdwQli2UnFUYE8yrll
XpHI8lq+Uz3viOg+3PAFfhXFQ5SqIwT378SQ+Lev8LhaaWLr/guADx9O/qm2gA4+
hKFdn6gCPrThiaerIFaFrBO5kjd362VnA4R+FLdWiYieaHM6vD5fyPRLXuuRIlU7
ZZgQxLGtMHslbcqkbt+gHmR2t/heIQ0NZPTKW9HRiSQL6c5HFkbPAbkCIbmBJ1hT
j/vRbkMpCPi60lUc1aHTzM7bBFqpinhz4Q1bo0NpT2apYxlVxCcf3j+xV6/bfCdi
lS4HMtBYBeeOo9NSMTYg9qCOporvobIJ1ETn5VT3wM2OwQeNCHNIUfuLiwTrh4dZ
xOphuNmnFW1wJwUKeNmlFaML+fPJ4OMN+BLo7o8F+lb3oCbsMgcgOYM5ETZdT/WC
sjnsu0HmR1/awVQAgWYdGxe5PptTT16bPDt495SQo2G2M/hjHRzblsnho5Tzln+E
Aum82qVQksmcF9sw9Cqg+1o5BGBRLC7nOi0eUXf9SsqLQZoIUC9/8tgecEEywU/T
IO7xcM+Mxcyc1lnoIIFv8KKY1YB23QMH9RYkljhOSfD9xhRelAM0DS/Q5wsb/WFW
og1EenP5i3ol3y2NESkrhCsGumGIelGtmbzY4WMa6O9aMLvJzteq/2UmmiIo92tD
0rM2LV/93/jPGUE2KIe6axE0/8X+UtGMzUB6NYeZfVUnqVWCvMBi8VuzYTsJOfVd
XZLE9Y2tNb/XPjYZBVO20vRiIxU5AKOacg259nafWjnMLOX0TREifRrQw/9LwOsh
Mttn8dlalulGkR6MRlybDsIGVyTN/H24WrMKh4qLlCYhKAUiEVtDPtXl0sKKJ/UR
fJEyaMakc9aAnUjBG7HEOwEJSCBXfeFyw2O22G7hu+27UV6HrAk/Kz1/DamtsVRy
Mdlz++FfubOLZbLfqkYEaxgwCCHQgzoTFFUJrsja9A5WUtIS5OyZGRasAYdka4e9
NDlAmuQLr8yhf+o16AkHWJ/qHpuqz7CcX7CsNByNvtAXsuBCZOUJ1e7FgF8Vnqy+
QcgziKx4t9c1ycjWEI4eqgRAsmTtQhCw9BT3i0HsWtixPPFiXf2gGeb5WcRzxLzC
13Bdhw67JLfUNkJhIKh2JV/6552hdJ50pElytNTyKM4yD/IGr8YjXTkv6iV9eIYD
GMJxIJ3B+qYMiuX7gEX5yT7ND272KFfrudesyJX180IvW2VKa8wpV3fyX8NqPkIe
2lw0gWzVqYww+UXrhMaFQLTZcNdPg5CiwgFTvmgDqWSCZXhkn2NRB8re2HorMkSJ
eddUsyaQSjW9Rhe5FOJH1BQ7JWZnodCSTf1n126dgGioUc3P19fyTy5/8xyN84wG
QycM6ITaqNu1A0xrKoGtQdXOgm9+cmsnSFjan0kmznen408XC2LcB97hLvtrE59s
Lg3KsgwF0PiLE/VVbLcO7omRNIazPhRK2f6/dgIlZoKGWAv1h/DLhycNU1Nkgmoy
pC8qlGg3rb4Xi9GpXKANKiHWj8BPrAWRv3x7fST0aasFVkrhVWMxwKEHuh9lCOXE
VlxigrBw8+ViGydQyDMnoC7zIOGBZbmGmhzjVuKzzxfPLNYL7Z746+nY9srSlYtz
WPlVQRpqjgnyjutzYbs3v0xPKMFB1YCGbBeZKt+VhBq1G2r/7/jdRxBCn6kpcs+0
L769JaKQNj/H6YYJtly+VsMR9f5W7HDYmBFrs7hYrp3OxGTkuYoKhQRLcVOt24L5
XPFSD1OsIwvcJ6OpY/qf/L9N9IJ3c2GXygu9fpoYBrZ7VcnCAxXnRmkQygyH3B35
9c1unJM9n4aly8yDnU0dysbQoFFfKcU3BysgHh2W3UsKElLIuK88GMpS59UXQoCk
sySRXgRX1M0p3IH7DCmMA6ePDZ7vL4PVN4QMiRo6wboe+IF0lU7nkgBN2I537YL4
YJHE2d66Zko3JzWgHoKHfs6pigp9jYjGiNqga43vM7l4tABhNlj6MVeiBRtr3d+S
4mW39cQgaxFro8Y8kydgs9WFIHeBy569DkLuT/shLyzyjHUSQbV1Z0zAHmP+e8Ic
Y6iHch13zp9HIaWJrfef2SIZyRQUFFkV5hCiGxCiaxI2H59bZc33ILGqLZtsN9Vp
3rooTasJ0cp13GPAwDW/L+fentffyLWgJDA7a1rMXhIxj+WSE+Dj8byi6kvfnXMF
YasMfOdy8UehPww29nsp/Pq2CsBbi6rHB4pm6QMpjl4d4VbdZ9dL8o5Lqhne6A72
wi45B5OZWVGq/aRdmG4WMSONURJmAN4K06Rz3dvgpyJNpYWTcTMjTdpm4wT2rYAg
kgvYJfq400mrhRTqy0XwQVf/IoGkv8knI5cJizS5nCz1gwKi4zQSotGKEgLZve5Y
oLcvYnJgp9/A20fpiYMVQCT3U987tQXWurYmcXL0qjDpqeU2jw7fSQ+aEDFyko2T
DmgT3L2NVuaq0fDNceCDOxSRYkvmsRJGEQFwUpWlMTOMCYVO9H8zVghoebQULQ1R
Iw0vlVds0WqjUZcBjxnwBwn/6ngsZDeOMCnYa5H6hf5uJKAIFPhXXlWOWrvYHkER
5JaN5BF/4myBUFsHuo5XIuPjjiIcV9taxnGaxQRMcVh/G6nkETuejNC6gsm1GMnk
5ZoGQtwShIQRn80idsQgK78xZ6CUoQNRzTVdSz6FE+ebjE45AvMtOZTpgwqTxGja
NUaC1H0IKfgFYYBygZ+AFNsszaBmrkWHPrendaqNXTV8/hDsCjo52J65LZHDKaNd
cqHIs0I3YyFZUeCV+Ia/B7OPGpAfcE++HZbcGkZtSZ659t5zYrM5NheBJg6uUtbf
ZrQp2nlGFkZujOvcqdYZDpWFFvy2i88pkYL4C149AWqg0zusdDkdoty9hZ13PxaR
Qd7iJUKeNL7/Eu8LXIVzYLmiOG0kVRaIFCj8vnpeElSvL6M387WIG8ch4/s/Mo4V
8/vajqppCg30iK2Wkih2fh60CQ7UqgMCz8rMZQhfHDyN4mqhyAAvhHG0u2sOyL7Q
rxLdNgi1zOJ6jfhVGp9FUFbUHAuOYhi7eF61ppMhHOw14Vcf5X5v9EmbFhEvVLRz
z9d/+GOpRgBpTGTQfdWkbxuDQTOJ5kIt6s4JlxwvjagapDSTHbXuu+HCuVMWB1tS
7spTW1KrJVPCFHhPmC7Ai+ma4tkrKepim9uzS4QPO75fwbjqE67mqaAu5z2qf6Lb
Y+jjqDCgFgGhOK6aQ5wN/0JXNkCShCm4yCwjCXCKGpP14Qc/1mLYq4no4LkDdk+n
aSNu7wWP1rRd2n/MY/B7nZg0mbGz06vVgwX28s9Qddgg2wuWl/xA4un/U6Gas50L
j5qhwMk37isnWEt8hcmFXCsyBfArely6X03Btu1wm9u3WcO1l1pGTh8myXRS0gER
4/hEwFwBc6mL6de/2soudkdQB6yrvsOXhrMPBkDSHsSzOPDTAF/sNPjklHUAGHQS
b6JfWPcOxL5nHnnfmctiXkPJYpIFXP/eRwmiSEWv++HyOIjZ01Cg6YPAXJ8DX4Z2
2pvlNZh5oznfcuRttyGbEkf5mkTEfusQjKcKW42ivo6ZxBHtHhRt+ldtUBix+30f
PWkcboHrXUE4Nz3uiD1cSOOxl8CRTGiiPsaoDNuemLjeHkMgyLjFPy3IeTfBxjKm
gw9qdHBpJRG93o7+4sojG+sahid++6SfE/YPI8S7GsGITkBTKP1MdhOuYMC9nKkD
/EC7/gzjXUSNutBX40aAZ1EOahPlmVjUyTsJxZc4/ZcqolDWNlO64fuRf5/83BOm
krpDn2Z36fjHQmTQEQiQTendVlNO0+7lKXaMKK9uQats/iS49D6VnQyO5NuSB8m0
Y4lprb0Gkb3sB+Hu/aGQdmzvGKHLt3fkn1Bq7tmHHVwvsoNVmWyFrrZTb8Kaissj
bqM41VDk4bS7kxV4LoRCIOzJmeoAkhMg1IKnYEucAxvElqDwpHt3eqtqRuM6Jlfk
H6cQdOEN2BQPNz26qG7F6BNLF7noBF++hhi2AQUApqE+1+R4De9r1AMuf9wNXpn5
WCkoOAIebkTwSBmR8A7Lmt0YUI0F1cbtBV8Kr8VHRYajQ6bqslLXtpZEqdf3hpDO
nPfhuPeYo4N7DKUxxsCK8K0siSLS5cvqkPBoUnyEMeFTts8q2Qd+UhSooGr20t8I
P9uK0JXY53l5nk6D6KS6gxJDd8o/JqsqjCggvnWTiSDmSlvW4EDX3T4+1SW9RRlE
KWfUVHIA+TRvx4duchdf1OIpO4ul/wfcLiO9W5h3YBv2m9whffBqaA0WXxlpstA9
8m5c+Xy368Gv5XLPbI9wyKcNXicAkymq0KTAP5XlFz6V6+Q4yQCZNZB1mhEhImEs
kS+e8nHk0vVVeKGqQWcbzh/qKJDSeKsFTnJ3X37+jWk8JEH+pDSOBP+jRnC4kxeJ
1xO0aisvmWRUljf80YpTmByPnmo4676Xl9O+N1N2/FYX2dfNbnRXNAcYVq7Xik3v
RCW8o+ha3HJuktr+K6V1UzixFN2KxF4mMHVtoQWATBqfIcIj13wcoDPy/0N3nhv6
8q4/oa/ysmIzRRTFhXtKHwy6dlZEM0K6KtfvTGg7P7TCFJOm6lyWrBN07k7QtAUD
Pt7mccEkq/Rc4TWrtknPamtZ/cjJHkmtdrwXQq310pGw4lyy6QhIHbSWcgga+8FH
WqBUKwjw8SFpfHuZ+nRXYIC0A4kb/L2UWmhQONl02Pifz6Ee5J8LPGmyHyUpMTom
MIvc7BdaVQ/0NcS+ocBaFQTgSyCgXtM8b5GLqqLfdY+VcfhmBjIXK75uNgiGNuzo
BQMxlJxQY/Nks1ThdtgqErl3/sCjxOCuC8bc/6zSpS8lXpmV7foWnIKIiyqffQ5z
mw4nj090GqypQSbJBlSFCOcYGhH05TGgWJuraGiHZMGQ3hbGKbHBY9ObSOzHyAEk
lefXZ2GiqXOfPhBroR4A9NG5LeF6UEVPSPx+ip6LkocSK0Bq55zQGh90BAV07FtC
5Ml4LHuRSB1e4rwMiACToilAc8WrEy7ceWkhqn7DeYEpT+XrqrIzlmZeOAHOAX8z
j5Pkx+kn37IKRR9l70ihE7GsvzyM1Ndm19My8rwacicDOffVy+bVb+v3CMme+DKl
r8s/9TxoLk70ycSUVRoM6zcMmkIQ12xUPZQbNcbyWE2sHz/EDoSAtpVsudWa1EnZ
RVnJgaz9vVUE4QqOfpWXxAfrUTmPcrp1nKkHTIpnzOHd0Xi98+9sZm9bHfdVILRY
q7vY4l+Zl1ezynBjeOtp9sjwYIEmR2YrkTX2+7vbtXsuVx7AA7vRxmGkAp5OY7gf
bQM8OABggnSCnZ9del3Lx2rO1UMiiSxz0YGOjii2GcflYW/3RC4vf/zIPaIUZgUQ
eHD16m/Gzlrhe9NiSn7lpSm/UN3243aq+sfIS3mrlPRfjtqTGB6yBKt9xnFSgIu4
X0F2cbqMpKTvql+wszotSR5lV0+KFdmqz/xMDtX3+caB54vowwW9bPuuO8Gb8kmw
yG3nWqWUFRnW719koq8vOMmKPBxYp4Y+MGwLodtgS/9sPyYhVebc3HxFazexXrM2
8Pof42FSrQxpWHTYdxpYAnTyG8uo1noWvgm8KkG9v0Rr4RtTZJpvBnJSUWV6z5XK
6IjdTjvRK/oo4txT8JJQsMOoveyGNhGlJscJkNfB3kPPAB4lng6wFfVltl2yIs5V
VyVj1Mtr57M5V+2fdlm7lcSaYJPlEcxUbOcz5xIAjCkifvGcEjmwNPqJ/FRK3y8x
RysvH2wlQ4UlCJ0IFW8hRoRz6tKsaFq3wzzPwrkGVj465a02L991pQa7/f3SGnFH
qHqQQfK3dlHOrH3VcZ7gKTFGEzpqLyEoFJVIVgfnvm61iFVzv17tz8h8gBQ09sS0
5sMF8u1QPcRtZH+0/2c4+OeYbsBYBll1fh/tfW1480ayimDwqjLfHyxMN2FM73Et
N+AzSyjt6ht2Ni+VRqNF6aBXkuWRAoKl46LfNoQVuEL/6VVnT0Gf4y8zDpag7x7+
INqVJoiwxTjY3Uib6oy4m9TfT/GaV9xNmryeAufZ2ngBa/xghIy1fuYVYCZ8ON9/
OlMqsXPKctljJNVJiPkOxPMgEadYT5yNGqK/ls5hyBzHEvnzV2dQ4jGO5IJxFIKv
JksK3kIOU0cz++LmtBIMZ3hAHtYtbprXtVKOPETxZWqQv1ALO2VsFZdEg0gRTvhQ
S2Lp6pG6TUaOUzUXUne50JzWfiKAp/c0qXGQ0ywL1L9hP774y+zbkmkWM2FAzxUh
Qb/TbmwtQ+7IF0Up/AB0ReQiaDDl5CoZHQHLiHOhG7WOFy9j+SVJkqDN7UWgqDoN
wfvIqN/gVfZ4qcFxKusxjsEcQv+5z2W/ldXVM1AF1LyPDyDOnXCKRbpygUnv1HQC
PqQYxuRZrnf76NjsYnE22PSGLq6RIGcRBv6BEb8Z3LMP+eyWK2Z7NfWnWmNAnGLI
MOYDWO3YeqgxxjYCyb8SGaJMuzqEZQ+/N4Y8mFqE+x+lixFnYmUiF+6Q4VWGcD2t
JTJnreBlLc1RnzzRUgndhhG4y/qholpJBuolZVJx3rTITYlrNBE3QDQ1rgoVMqB/
u9mAawjsFk2Tl5auefCN2VCY35ClyU/KXDUovBQaDhfTltBwJdKSXDpHur9922Ym
LO1vcHussi6bib1409J6WglGxromyXGlDjqgLXfxzmyDwrzU8RIc0xTGD/0NDn8G
I24h3Guhph3I4YUsCYSKzU24p1l+fSiwhWRTRmG+Vd3yOmgWM6HxOKbudSlplPf6
YL9DHW425rkLL33wDSHSPg6Vt+19jTiA39OxVCiaudiSvMiaA38QwcvfrIKP0Le1
Yb15yIpQuiNlrXp3KAj+ZXOyAHpjRD7sNNjGQZfYJhHx/FSfWRU9EOWGIY2DmPuc
MpXrj5ay+44lj8+RJ0seqenIacbb3W+1Slh34c63zVLs5ZY6qyvsbHibt/LAd4hN
AhI8zZICuSV70EZq491aGJZqST2ApM5kgbuq/fEq7WMKKob1vQfub/zLL2QkQqW5
QtPDGF0ZlsQnq+aBJZ0y/1nn5hMzGWdxaXeOXJpFKLmlrChtyCkDScMb/MnoccpM
wKOeRrqKzeqzzZkTzPret2nc1t2HR8vRdRCC+mFn+oUO1+0iUCuUPgPbQFZWcAMB
4PI8qYx3aXqQdH2l7ObQBSi8aqd/wjbeY8Ay/EKEzXx6i43fxCfV+T93OFAE2/uo
WeIBlF9CuXdJZZV1hd4miR8eFeGKuLNGuDrtTSUsgqwfZGAhNlXSarwEQm2GhYAx
d4R4CCYtjF0vGiVCAeIVMnI3PGVtrPo/UiHc1s4nLd1eTu4k9q47STKXU/4xkUY5
wzgfVxRah1Oma81neGaogupBRAPAk4NbgCq+djTzSl9tMKHPeW+NJssHy9WLiuOD
N6TP9IXh8rrMQt1hTDl2VJ5MguDVeJAg+RsEOTswGF/Fu+/4RG5bXzHl8TC2AkeV
bU9lPLkmRum/sObZZpwNU+CKPjRZDXeCzw6Zup9I43psmMk9dgBcWpvImH8aPOhY
KvPFQ+DJRE9PL6DASE+YT5A62qnHWyijNrSUoURDtKVkLcFr8q54qERPbHZMqfGn
2FWy4fpPQOQkODuzXPedVvLHcLMLUepQCT3aF4liWsYDr88H0yoRJA5P+MPA6H6R
QkU/JenXgXbKG4mCrSY6ZwBaVfxKODOeDo/SwdrUT01dhf4tAdTKWBkWSCnxYOxk
MO/WhyW4BLxGyL0xBakeQmajC+6DZ41arCRdBimyurVLOvecDUFJCIkgU1AhFFHS
ZjYIfsRaNvfKCpE54soPEoQwlsWf/36hRcgUIygii2AQc8nRFaHpTku5Hx+cFjDQ
HB2m4S0imh9WAlMN9O+J2wa0v4VVqOrNrVhVFNa4B0+oh2mod70GogH6oFFv+09W
9AydRaqe2U7H7SXRI5owDVjvVxrRJB7e4G1eGhXxMqgoS+bXnXPQI3q3T8sA+dkq
FMuOa7aeppBAhMuMMSiRfFlxZ+sRM6hcZQyfaI+1tlFXkAekbyr/2nY7KjXVoV4i
9AOdElCgetbXBBZiggfrci9O8d8OWuSRBObLUa2vzhOpPlZLttUzGBAYQ3Z57+UI
IacElYGGjMOnx/h51bmPzScvms7tNikFOOlP28s3JyaaZniB5eti0F6P0by80ef/
eUkj/viCSy2mjzwXeKiq+VrgUdJ6gc2EqHi9uNuk+cMUN2+Dm4BzAPoTp2swIOHs
9EG9+Skr0vknBdN/Qm4ODAmFh3MeXWpT6nsbo68xyvCFbf2LSLOrbicM4AI1p6Xv
XElAgi9SuceuLPbn+/BKWR9ya+q2pLxNwkoKYqrl/M2wmviBot9C0dN8KmCsH6/k
qWYLm28D5ySk9FIhrqM5x0JXmbzm6bnh+YwOkd5+rsVjEXgp4rgM0+tAiXCz97LB
vMJSUfF0PkOHGu0l2Cr3/FIaXS++hJoEOJ0FVp94559Zzlp0G4AK9qFEnYNwdDoq
6sqvpptvibU237tPQh0JpVRFUzB24lA7qlzjA6d87X02S8Woru3LsG+aHPom1AAA
N9AO56Rel5BiNx2NL5OVRzNdMfVFjJu272bKtxvfK3IfgNkl1CYM5cwQBhWE81kJ
v+x4avD1YZOVTdst3pXmECQlhjX2mkLDLLwg9+ATFZa0LOcNMwlSB3Ktf0iqnr8Z
pjAGEBOqh5FsNvL5HTNbo18utTPX1Lw7H1xb3EC+JhkCYbVWzD2v+f3+1M1qe6J2
XCIor/X7kzHbCczhPQRAFC8fQnVuO2r/PsiyY1CaouNUxmIX39Mzms4hTklPeKxJ
2BVXVkhYOL3fCEO+KPNZLoDLhRm7TCHOWi1j8kjzP1d0FKsZLOXvDUw9Q5l8AFK5
YqpySRYkfoxVLHIa9o23/Pfto3map9ilQHl0WxT75/XeeeCpEiMMnGjD4UUFd9Mc
xyi+FbBEzhCbyW5Yi9GlgKU7K+/jdGt/ABoNQBr7MBoWEabFtpprgY5fCCEVgVBC
W54f5+S+E/ybsJUk68h8OGRH5Fyte0yUibBlwUk7YPWrJvTOCkq+zAcGUv6huRZG
CpcDhS7SzILPLh3GRounVeC8icpS+5xs3/y0AVYDcT0RN3/eNsDeXIeOEz4qLz/2
KSI5H5X3I8Ub9DunWFDrx7lN0p8RbXeqdwNLWC2QkHlgyEv5+5a8dhCeH9fRnfYa
/dzzbUdszDDG5TDdt7WiGbC8h1IsRWuSkiHPha/JDviRVLXw+MWG3Qq+nA01sUlq
9dNw66ie5OBtbt34YIDYQSRqMfwBtMUML0c9drf2mA88GSzyVLnc4490IVhzBHi6
VAJzsLkgVoAyHsMthcipXuWA3TXIq4S6U3s1mxpyqxNmMDexT8UNZNtFHv863kt1
kXTPRfSOo8Ja9uPKoXtjHXvP2AMtLFD4GraxRz4sL5kFKH5RC5H8IDfpdji7dpoM
LM+mR6v6RowoALDrQ31+vfKLsni+nlzyTpsenNnm6O2k/zZIgQMOVYCSzecja7G+
j0OgZbz7BdqfYAR5AuqRafhW773YTazJMTrdwLyodhKFyramLBuzsW+Ojo8TsODU
jTEmvDfBhkGRVkBQS2YtpdbbIAC/FQ/Iy3G4hsHgYF8l7bZI6nJtFswMvCmXpWUp
V5NomRDZ5ypqXu5rdPMm7hdFv4Ew5lAT3b6lxS41nCSKgH+7W+BWO3P+Yip/NBjL
KexeALgzOcTayY5MOpFPlhRPutfAjrCh+Oq57mmeeTOwYlOYK6X2Na+psMzl4M7J
1R9bACcbIS/yGWFXd504Hn2VVkidsCYkFfv6dQpQZZcREjLRdHCE2cIzAO768GMV
dJJvqJYflEAc9dWWANQCvlOGtSuU3wx5wk9pq7psJn/dHUbr5/Txrgx186ztmjm0
1m15ryeTJR2a+oGp+KOBN0r/0cLVU+WWKj8pZ1VVI+vJoVTbve098WzLncyw+bAe
1a7WUrudSvLjgQsWFDBX6+jf3H7wrDLAZ23mhbG+0TdEGPHmE72NdujYvgDEwGc6
Vk7lCTkPw31hhCPZEhjXEU0Z+onlitnnijySzrqCpdiJ7cPTUPA/3qCW8UEcdcj+
bJ1/JkK20DQ+LQv7An4VHfPUn0W1j5HGBndR4X372v3hKZGU46KbXBrtTSFAavCU
d0aoosMCUxOhYk90EeGStQmcfHOmfMxQqx5+jULwx9v8fLmK/4QJilbmBgSERwXx
8vKMeDfZRYXNIqB5e8NGlZrFB+4uuIiglgU0zMm/CeByf8CXIla9NDZfK0Bl8/uy
l4QoYMX9ysS6PvM7eh4Vr0j4RpBj6hO6hAH7CKYRqtC0lE5VeB0LMa8WY0kyQS74
Bwb4QOJylKLUI1SdeXQ2g2VAsgwdtWeGNe5X8z84HnybYOfK/z+QWfNCS342jRUG
3YlPhUKUvHZWoJQgD26Lez3fDprL7mPt9xb9rNIlhUCuw8iAb3KoFmhQ8Y6igIs8
5wNfkYIT9Bjlcb229U1SCPhmtC4NQVOZ2rQ3QeC2Nvt9/BFkBGsGJfW1pzrMigMm
+QnnxUvdU2HyB8CsofeMPQ7tOhtRt9E15W+tQCLs5a1SvwMs2MrbFkXknnp6+HGu
8C2XUq4r/u35HS0tH2cTdfp9eGA0DSmNNDyBjHTDunSyl8xbkHS9mWLy73Y6OV4+
QgWVJLxJN4HUMKeTa/1ljmGS81Y3EIm9Lj/j0Rj5ocPh98w+bBG9Csu8XdFbAsOs
XoilWDE+Gn7rnhDV3CaUk23tgMUaM+0xcIqDZvTusoptrF6nZ/lBJdjG/du1aU5p
jJmDe1NgR4e421KUWbZpQLb8SyTxhzctW61BngithngArn7wElWAZUsT5DGxP+jk
0v1TtPLuStokksi9unqGHWeoo0aZbWgqvZTmXvhkSIEg0ivq8NPu6lMk5OUplhOE
lCi3d99jcoH//xb+jtOtBKr/v9NDkEA2/thZUJ+FachD0PDo3fqDV8b35Z3RZGCf
V5I57MTahlllTYwYzzsY6yuoba22EPoH386bvKP9KLrrc3vY6iFfgs/HsfNlAGlb
h+S7kS639L3njwNN2l4oNxMHYQ8gprNV8Yh3DzQyHjq0q5EohnOe8099u/NDqFnq
OzlWUF1olnbY/2jFHY2dpt9eNO3R1KtMJG2/SV6xvFj8n61i0FBaO4fwrAUdiylX
U8/liqvSGaNdLSxP8dev2gPEjif3DHSLmRW1NKDocRZTY7eOD70U6Du3VP6jJpkg
BQ0UpwvZZ5JmoKRlKASCGwatboFQb+ToxTqnogoDibRiSXfe9VUeBAY1APQbdq0x
xXrPm3FACCJzHfhkmV/5MkmFkPDiNim3FwLGGQrtT2AWxE9uVkmpdRqIrF//Wawm
L0hSnS1j4CLHwIrS8kGjudOjHF1Mrq00aERQDt9fDGkicsT/b1duHWijnhkDaB/3
BChlvFZhcsslB2r6C/ODX7Rv1gWvyKBbK2kt3MTNBFMUFOFzGHyUBHxS+FElsqaT
wjwCCORnqk4kMgxlWJoQ/NrCsmFUe57DfaURpyvPyxRnVSLD9XpC7GLHqhpJ1+GS
VYu7RA0ZbRaM2FhqdRdVnKlLm+VxUzMlLFEgm9cohkmrLj4/gAhVIwdk1M3cj+II
CX1r8mA38qPAoqc6QryGwUNbe0tLYDkOVgtI9LDrjYYShLCC3uKQa78QEnGjGVsR
Qq6xflxzrg8vgdBK6kbtyMUf518a+/FSRLaGExlSg561Z2zECCTQLdeMvTIAU6Mg
tYc1OeCr31YXrc9HHgg+so99TyeohI39Wr8sty1J9rJte/eFtnKPeAyLZMD8bqJl
bv0BJvmfk8P1Pq46sg8pxuBtsC8BzbVCMYR/Sa7ATLGObPrXtFSshqVs9UtyKioe
8Om68A1Tgn4MzK3tD+J06vfgQGpFvLSCk+2PbFC30flSNP+2fEzJc+XNYlSMTdg0
rZsRsYwIbO75kjtFtCF3KiquaqrAjIn0JID8KYKyJ8MctHoL7iCOaWEvHXvKENfk
1JdYQyFT1x2nFeCgUdjblSVtRqVuF3+FQdXhVdSZzBdfu1fznypkhoFVQ0wxWlEY
ajAdI/ullLRLCoI+DGjAHU9RLFOxZULW/sI2XYhFN6K1DEd4OK0OpLpjs+1Ty8IU
kWo1pBg5HOVYJJl82A8GzbcQwfGRfKw1tuIIJC5Ko2DRU6Id7CLAOscc0eCZXOcn
3PFolq+J4FrzNO3KHPL5YXyK8nhDwmI0ee13zwRMqqBWkjRCDgFs6Qg++AiI2Og/
iJKIia1Sb+Fpe0YN+Pg6qDQArL+ipfGKGb99sWMa1HeKXCR70Jpeo7Cy862c5BT4
OK48jaEOzuwNnRXd8vCKLZqWMzQeOH46AFH+LofRxpkauYhj4MVSxnWt+3dE2sbi
y1Ik8kD2DuDkhOIFT68NMJxI94/2qhfj7FmB9XS/dZPCcYrJ7tuHe/MrQYRoU3rs
EN+2//8JB9XYgSJVODb6bXYfeMlEVumdBPVsOtrqdINibJzn6zAjBMLSn5IoydWh
Em4Re8Dq0XqaI2I4wpDVDpEpE2AsdDE0j5HiQmNwxQOliMXHlhEOiNyIKb29JdAB
BNvxBCShS6HUlHo9ms37zGvpdUQxZ16QfMoWADN2THgGf3K/g40HagGwtFSILDCm
UY6OQGMX6w9UDv7OeexCgsTltuzqhyXuklt1X9oif5RDUoSijgdCzXrJHCxz313R
ybWfIlhBZj/230j5U8PvrEEZ3jsYOOlYqPUMUmKv1CGH77smQ3tguE6IMNSnB8Fc
t59zl4N131+fJXvjsR9fSMeIor9jEfminko3sjdWRzio4fRH2cbHWf1yUR0nDvdV
mvKWrRDFp26YtyeMZCR4gNaOX6mbMSqY9cmJWS4Xq/0R6aG/kOftfY1rrofGLttx
MrzxbRGfbsiL7ssi50eYM8GbD1DnXARvrm6daCiZHnqvdqLVG55ZKHhwSTVf7wkP
6Woj39CDlkfY/bdQm2MpM+fA6xwdLrL+usyesAFbNR7IDwG/cmXlLnXOcZ5wYYHc
tYW5LSbMCRFq1Pf4qfhUmX6QxC3C1gEc/1O8l4ZfCkgr1sCWI0hV+He2H/201W6y
Z8kD+t9HncITgeCkDLNnwaKlTPeoQ6Ww/7IUGv8m0Xvz++xy9+8bUlLUFY/frs/E
B+8hBN22pNjskTEtnkztQ9FtKG4LxUYyQx07En7+KjkphvhDv7mVk/ZIZOkzzrFS
WviMuyHdN+SsZWYH6D2b+briJP3p/A6Fjgz1MjRgzJL7M4hHeZ1AGh5S7UEZUMX9
OaYHtY3Dc8H9J/JE6UfuN85ggVf+5SCO7OSvmi84yIUxI6VLhbaQNfzcpLkP6G2a
6VZCj+R15qgzBXkl12nNWjJNjPodVQP5wJBBkuX8jHz/4Hf1fm0r/SFmUNbS5jSn
Kz64Ezx5VSvEiOReOpgS/ivYmcFyLrRWGn3AmimA+dQWcopFQvS5jYtegggvypgB
Da4NkshfuEuX2J57u8IZe4VsMFbcGfdHC0F87bfuaVi2P/2QLxLJJaEh2WNOzAaf
JpyVBpliXqV3X0ZoXahlNFb5jfUE0WtSv2KG1bHGoLGlCKXJz4VhLlFYyZgmbS4G
wJSYBNWsijP/MvVT8ev9XSInqkqmGjA+UioGoVLTR8NrXuIxs4iwz1aq0644ClGG
hZ9SR16JvBiGl/5KoZNwrCeykbPpOdzOpYYRNXM9ufb6ZIyTB59xJ4WYzKa2D/PD
0E7wGIAfaMZScSM1P5q0c8KBLTncwEiE+szAWFEDx0xulBPIbyJ1DM5UANDQbG09
0Uy3j6c3hHWddweDFMY/tKjln4NFA/U8mAG/pB1PjQKHzl7XWtw+Blg3Qo6RCTWq
Fost0q2f2sxDD+U9Z+qOYQnQgzDZx+J9fE02kA++UBkTZ0SzQSuUKB+oh/48o3jW
o+HFOO0L39ZlRXyjZpCNkrP53keeqgoKoOKxQ2c9keVcZ/mFhLR/Q/7ijmK4ECp9
aTkZypVsF8Qq22lcJRYLCuWRr3MogMnGYlxSrecyIdiatk0i0faanfZKLm6DHcgL
TtOyTQB8Z78AfrrhTEELngi2hcXch+lE6/dFaHXmEPW21uNU3nNS9tOdXwATSioX
BNDz/U7IXbl8ogEMHYwYobj2kGhAyTbiQ8NN7ldE7lQUlLg2O618cTWGTR08czY/
UFhbefsJOfyl4a8oC45vWclehoq2nNeHmupzfD4ELLyQhIhO+kYytBMUNGX8iQ5i
hUvOd8K3x/zoCEGV69t0pTcTbXR1e2+bJHeiZqb/I0Psy07ZV01STNxZ431urAZg
Dq3WFcV/f9t3eE0ZNRD5UxVex/bVnB/aFtji0tdi7ZkfyzakU0kAi/OLeHqzvOGV
7UkhbemPQbuojJn1uKClxlx8PK7vM7qcC7YEzR/RqDAZVuK1oeDvBxikfY2CYjw+
olTSOV4bh1isJXfEYkEOuLBEhKZ9QXXJTYWwvvppRcaInsX1zwEINus4En2inH9k
glfp6z+p+a+RRXGEoz+PTtc0z51TpF3pDuEBuHXgn5AoOQNw3Kj/jj0STVw3tLid
ioQM3oT9LLGQOKVdQFu2v2BOQ+iBcR7w+lXfM/ZqWBQlns/5NWLKd+wnCxHYcEdi
JFYTHAgNaWXp9GVQntzMxCoispx3gZs5KkQMwHkB7UE2Ki82HGkw9SxEePHDFvil
/FVCYwSPY+cNlVyB+6PdlnmQBkZSXYG0VXZ+Wm6LCPGc85wsrLcLav4wsOHmFpe1
n45Lhua6j6YMpwepACu8dLZCR01Bx3rB9VgpPVQJOuFsaSTANpNq73FjHAbG1cS9
oefQKosm7g3DOKM3UaF4GSQFE6/wxdsOjyM/nGpGBqeRwicu+adR0lb4YHVVSLX6
CtyO2AH76J1QzEqG6wwhizcEAYrqSCgdt7wsXUXXtY9tdkm7R4v3DVVdYY/l1ZJ5
TarwfH7+sN+5IvYWYqMAuyzv9ZGJ0Ip3uE000J6D3c5v1dvgOmGxBlPDot34RQYX
dHBJWO8LHdzfxOjS/2FVRtuYzJMp8kwCe6bCXFo2wC/DkmjPbxNRyGU+/uoaQy09
yW7JAw4UoqrRz2c29q1n86afYlhb+hEMdCd1c6F1u7rEghY7EJfxAfRTIzwbgAcO
TTj0vltumSj6km+A0TTx9IkIRTo5RCOAIJnIjS82VG1RrPGiwfWr052+2Vaoxpm4
nST9cUHtI+srsg2QvHT0Kifn6UHGkG3744jX3A1/ovwJy/YO13qokMUHEAYLggiw
1r1wm9UxBr3OwoGwyqMGn6BP4ftDm0nF9XM8/pIv/T2tcRHo7tL0GzM8vSxFr0pT
4kqH6AystFgERN5PqN4sILPvbrfIv0pk2DfHvlMHjPgRKkT3aCefbDKser7UnxmT
Ru1arkcU0etNMEruMgLvel7EqDetxSJAiyFAgRHNyZVski3nZY7V4Wn/mE1Xe3rV
k8iWUndPcKdvXcCFCXjZvRx8c2q36Cem2czrocD4/IjqjZAOJDMu35ojMoXG0G3U
6JZ8CXNEpJNHwGiUB+VbHEzeRnMDsVNwrXhvHOXTxz0Z9K9B/aEjTaZdEIEU92f6
GwUK6UBXoBXuluqoGpCqZg4ZP6FA8o/fFTaZUbW6HWo7nSBHjIEqkd+PhBg+fhm4
+5RQflV3pgIRkqohqRixkWVN/smpsoTd6KPSs3bekEd9uy6sCq+MhfAGZpTe5Dvn
FtB5aziZBCf/zkAC6GD2V7Ptf6iQq5dQGJXiRX4OHo7bFvJN/foz/fOg8NIaIMiP
X2gzwuVpW4WoEbDBgyp4/vvq5PrN2wM4LdvNV+Jj4FsycOci84RjcJ3MHf3wwUAt
vQklR+natzO2TIEJiJDcp86A4xGK69Zr7WAd1I2YKiZudWhqUi4SjzUqfIsckvym
aypO8hrJM9yCyXhiLoP5+5UWqQImc7Ov++CkM23tdPVbXRVyySnn9xzY9bOipHK2
1CdK9O3VTuNAEFsvy3phztwRkxaPPCN8uE/6SO7vfwHcooh9aDLXiBsPK6r4Kl2I
qI6IgXyjY06otSLIpqlhgQzlzm+UbmhrnPlGx3gB8oj6N0eO26p9vScK1Uwk7dWk
xKTlV0sHDLGfdW7CFk0oPnA74sbkhGQxyt6ZfMf0+C7y5LXku7C120OB+nTfM37M
V1OSMk8g1U7mXQdJjMQZN9fvp2K0TcwaeVK97soLpdi4w6vaAhiarkhl5lqLnosR
Y/BiE+T4pF4+t39RU7WqIsiEXrh+mep79m/G09j1snU+5zRgTqRVRyxFTH1YscOG
CLnsT9OkEeeLzLQDi3dX0Q78PNGFOgbxkjge5UtKDlnurmkYUyeVz09+f9470Mw5
XThgmXMkwWslBu6R2K2kvePIrdWGqyC+AJDvBQ13+nofJsWnJDW2GVBntH46ts71
CJZKJqzNFSbB4NrKyyOsmm7krj/+Zv6622ApFoFh1RwMQXDQ7rvXUIc/OjkgQWya
3oZx6lKY7gFhlmu6oqie/Ag1C72/UPVfQsP/HXe1k+GC/xcvE0g2ZrkJJT+YJoJe
RNLxRfZwQRvvvuTMjxb/SRk78bABvtf2uwsLgguajbUpYK8xa3oXeHorhOHae60H
9anWCFb4gOdJCvN47DbJjmKeVyuQtVkGYQ5AL6r/QVHOs29NFGHs8CGdelNZuoxL
JkJZT1To4qTC4lBvUnzFf6hL5jWI22c7OVm7Vg3vXiaUpNDakqHg7daWII16vw69
50kBfvah+CbYukdr3dIeRHoURbyRuhKqMd+SLPvBVjlIVkol85JvF9y665erxg8p
s905j8MxW1B7BQZmFD7WDebb5/fhvIZv55+5xnWIPq0uCnYKUSoFPm3P5bBQtdRc
sVYK95tZm0h0qcEElqvR/Cw4e0zdrneMkTCOwa6TKzuY3BBzVYNPoxoJVSFSc4oc
8eC0dxu5KBNw6C7h9bc56pJkdJRoICr4GKCCQjXSHDWNjp9JdC48U+n2YthM7Q6R
4PvG7K+COAJMOXVr4eCDNOQQ3+nGwNuOVZU0NQ+DS6S0T87bttWrGCiBwWwle1oN
ElwVj6mvEdUS/fWTsjFyQv2me0sm/h2aNgAg8jqhHDf+3zzVJp5QyMpFE46cVGco
8jvdPqV461++Uz/L/lnx2KYbIg1dq9uL7wldH1Fpkr+Y6Ub84HN3C3VOjplqPQ8R
zH0qubquksya0S6Pp2F9aCCXSIhFMQWOIu0kt2DGRtSkTzBcNASavx+tE21swdnj
YBPTY7sxN3zYcsN6NBF0/qSY0L+MBTfU2Bv5F2ZoF2xvM2wy52tWPbEuG4Myhr1C
eAu+HuGftXzMrqbk8l79cUZ/KkD0NHsHLZbuYPctm/6e6D+kc0ZSgxreKDcybPxR
RugkATsd9/YQ9S02iAGo5cMZm2Jiy6ckRihUWi/1++JJtgFPtpW7tY/i8nFZJWNt
Kk3hU3SPtkntd2zsVs1RQQv3/ETf5mUmUSO1cHx7JC+TW2xpxSkl6O3wFYXl+45l
dDgBV0gCBQ9MqnheQQXezvU9IQA6Hdpx4R57ViMGLjw0FUarhAoixOu7w4fhtiKd
9YOh7UAbykhNhJ0Mu8tw1HYCqfFdd86r/BiEVwkvgljTQTMM0I51yvUYD/H3kX50
mK4fjB/VfaC050QseaMlmP+dQRTIWQAQn7vE/1eH91tVxUnoR1joGLiNOciNVfj7
cwyra+qHlG5pRJqcoWEWVU1ZdZLSFUlyYacCLHBV+weVTh9KXWbVqCNlcn5gYp7j
J4h71v0TUefC7gT147p+kvBkTiR+5e8fMKMTHQqqYUaID+e1ubnDMr3IZLP/RhoI
M/MQpm8d+Yw078Z12+G4bNeZdJtDxJGSy3VQt1Oqn/GBc2S2B6cOX1kesS5ltYHY
4WNrCWXSYwh0tkSA9LAJuRzeNxHosA7lWYAyqCnK8gLLoWO+RxAx0mFKc3AXBOl5
q36bZ05bUiG4ZTz+KGdEA6qJpZca3rhjvVYs/ZcqmSRrVhhBWSGlrxmbpxkcK7lZ
4wutnvqjDTrNzKMi3IgrC5MfMvq2HgtfLBh8kB6tB3lNGVH/s+aL46s7TPQCvEqc
ymFwviYX/dbJ6F0L0xqDQ63qKRZsxLEOwGS0ZGl+ait0i3XZofzkV3QcsYzhevrx
gJ8d319dyPurKIKtXPOZoGO8TOpDtzfIDn/RsLN6CUev1jYjN7NAa94bEJAhW7ZU
BBwaDeVpS46WLYwFtC8HEtUlxYhvLIE9Qx+LJTevdgRCA8ZfJ9zK+GDd03oxins0
y/Y0aE5hNJiMqJyGBpkOC71tg6eoMsFakQL3GoWXxD528tGSWvM6VW4jY5+N8hSb
SIHHV8YcFKGCKRhcBRbPcg/zh4Mx/XjJzFrQaNQAY6dEUm6Eth2JPEPU9G3xLJ6k
eSASRJLp056n8woXbr9am6AVFyYdIHjzpAUg+t+eHzN94D9E5zlgFM0lLxFiP2O9
r4zEhWz2grfLzpY7/y0rcU9z4TbwePWw6eliIRe/FA8ETYBlwoHfzpU69o3xFrLH
a7WPZ8O4XuE1cbcDuba6c6USWAtWqtKraQa4W7vvcFt/vH4a1R1/eyGcosKEfLR+
/wYXEGy3dXqJ00pC618/X9+AwyfUK4AZ6P1IRZBVPorkBKs9kEbSgJTsy4EK8otc
zmiXjGXmY/EfKJ6+UPzXH165atwRV2MaTtFB+5LCHHtahrQnD0yuMuxQv+ZYMt8S
UYgstTdXeCXZdOUbUu4+N0oxgDD38qQfsveK9FxDojBvc39s+xCu5o/h6Arfo9bR
0DOMuhdXZDpbm4R0+URWp7XJwtIOhd6BzWyZgx75DLEX1vnAKN2JaVZd2AMV17QJ
liXdsWjYJY9Xh59Mx551aBtxsDwMO6nJdFrhiCKP6EdVHd+0DFsVJf+LbF3iP/fD
O4N1aJN2/Y5wLz3QJW0etHQKFYSurGZWmL1s38cw3Irrxb6O0Y0s0Wv0Vt4ySM20
6XUlOfZZbNEaPXoW598jN7yonUNd2OKNKYulg2+GhD5pwBG5QiosuVc/4BHvTrAQ
Q1kx/3h5Lkn/A/VYFXr1eVBu8YObUrwhuKetTXX433hqqDEtWwhL3iibs/JNkpGx
kR6fuY70/gAdd4QiO7njpGLQrQbMWy/kzmV/Qf/PuymTpffpx2/+xoWrnQ+sU5jq
nVlR+xE1OUh+x5R70TM4+Q3slrk2KacPkal/yesp8MPBNufmxHiecIU96gs2sZ7e
QmRtG62iu901kDfbXtzHFt6wAwDRqJBc7OgB3+ySX6CP1iO0zL0rLBYNvm9vNbJj
2CHeIHYvk8f5XAqun1siuX9sFGYd+qAotfsG4d/b7RVx5G/ZvAtM5crzlpP0tDd2
A8qRZcsmC6VEINIS58sC3F1bPO141STAxhi0Q8UimtbqUyyycwsbhEoNBCzyVRFo
ODS65pPeBgHebqZmqxt6V5lFXqI1dhjIj5rlcHZ0zhXL3WmoLVJvGtRHco8OYoLe
oQyvSjlL9/hiSuUA4wgK+iKRms+WhvekAcGL4BHL21q5mzrfC5RdUps9l2gKVKXp
e6bGa/OE97xmLWj+fvNOUNgUXZChM4A37dRuA1igk5/m0VUa6f1Uks2J2W5eVgTb
ka6RpEE/NN/I9G7tx0314hCbXJJhTW+A9/1fS6hcqkSBkggtp/61TtbBdCyhoRSx
mFQNj00pb8j6OQcxYqlCrITVB9RKKX8nG37FddOHrgTrP02T36HLWlCLMie2ibhR
PrD8kUUcs0LYaobAkF3ij1q+FP2hzAd3xcfEO0Qze9RiSAd1u4goUSoXIC0Cjrcu
QC4z6UHWuwW70i7JDYBwA2mqK88ONCM6D9uVEBb2SrpkWenAdxukrqrrpxbZIQG0
d46P2A0Z+S11S6Oug0+WtFTtBF3w9jAgMQqQU6b4zkl8mxRKrNJrOTH7ApeIj+zZ
+Kk0MJPfnToOmvFzP/YiFpyHb+RNY9iwFuKX5EN9phTZPNiO3i67Dk9uqV4QbGRm
4eMwcTiCfByOZzWmfj1uq8Rovjv8jAJf4R+xJrN7L1QhlPRTGIUxU8WBG67NfA2H
0OEV//M//fvSBds8YN2kaTlh9/t2Uli9axuBDG3EVu33IFM1itkJwFdpmd0QiywW
IHzj6RMMQ7WuCRtsJ4jl8Lm68yslJzpTZSruULaOLhBS/hyLBKmTcHa8kEqsnD7l
iFCiOveHdPFuUfyfSTHZfuTCiLy4m0tVNzjvwyYQHmr1bqXdnA1HAC1qiraQ2a2l
roACk2IKh4EiSb2el/j23K+ttexp068283lJvW6GEt66oVkXapuIE2rh9vtwEx7Q
5BwWDCnKQw/GKsQqiKXTz5HJMWUyYVklczpT6PIpzkUsw4xRJ9TjQprHIHeYOslb
5xSYRFw8kfU3S25pHalmMccD8maDT/xa4J5VGeXE6T7EUWRjwMn4kB+i285N6XP4
FqJju6XrrnsuhQAbhJf2G6E6slPs3wTB7JjyOD0opRHx1VFeoNQpojOi06SfbCJ8
ZdTirWXuQCJn6d/3g/aMfPE+L+Ubhe+ZkAWmyiVPPk1yzCOvHv7+fxdgNYkBBEQa
G7V7ZgdvdJ7qL/LxCj1O6+gPCe/UKrIXWL5cGheGCd4u2u9JCHUL2bwqvnZVHG18
bybvdw59x1RlJQN4qZt4Bzt/2Zy+8CKegrfFB337CGTrsZqxAKBCjynMZvWggO5c
ZzfKTlD+yyZ9+7W2JLKuoZ2X6U1MaMFbw3mq2X5k9JlXHQJYhpSrKogP7GloDZQl
BeGJWY2Ovk1XNDouE2zrQGHZpr66xevpkXhLYPiuPl4PV9JkQGn3GBHeThy6Ml5C
Ro87TmMDkr2frYC6/ydMSrg4b8ZS4eVoCpqlA1Oi48BFCrdlGap2P6Qq0rDzdJBf
15YCOn+MFuC1nigNHaxmQ7I4lAb/59qBWJj9gN0R0sVNVj/skJZeqRtMBjFq7RH2
kJvHQUZ8/p/G9qCe257VN0/xvBmqTEDSTRJl7TDL/+APRHMf8THprvdFE/SHAJ75
bxaGIxjKnZw5pOEbK3yXlAf7qWRyscKbl6rptcZnxzXSxqev0OGzYP+EzaJzNEe4
T2Q8IrB95r+zYv9XEHgbHfxRVC/jp1zcGROdYkrUbg+DrAhsX47GLpPBMBHDhpBA
InEu9sqgwn8WVljB0/rXsFPjtk6LKrC6sSudgoFeyTWnEwz3N4Q3OGniHRHpLmc6
NHMo13uk5KPsEtVB9y3dx5/nh/tlIygjD1ovmW7YduZov7UnRKYLEM/PN7ivQdTI
LqXfeX2GVojb43XXO+RchcNpCFP/nE+vBdmlVL61rynEEsKXmn+2ARFhLg1Szf8b
TXKmQjyIr/puVtY/jSvRQvSeZtSsuNHkJUsSYyhNRjNX5pe3JBdI6bqvjVB+msIb
8hzCQIDE2r8P58o8+Xm3PiXedZ7L5rDnVWMy7/6/mWUzlqkzVB6pQ+Cao2R2SkGp
L1qQGDNicI+d+JSX9hFwtxJZPCuACi+OfDrLe3fmPo7gL4V+7Fnr5HgGMRafUqSs
Y5en8+g2RrPMXZOwD8zmkEq8rc7WfoS9Iih2W47L6wftIMPMPyLAD3zHH9PrzldB
QLfIrvn7cR0QPgd85o7brL3X7IHJRG91la60dN1Nu+abo/zQ6VCXw0hqh7o8KfBD
UXdTmFR/hQ0TqDy15oKjCdTj2Rjqq9/1hSFaR6vG0otxrZn5QuILnUB6Y3/KeCAE
RfrHXhWeZit7oX1FGM8S4BQ3BylSh29yRCYjEG2xne+0HNfpanzkdjNu0P5Umnm2
HCF2CGT1ubQ1qLG7OIg3aSMM3DYxX5s2hMbpP+XCB87UYsJ5xbXpp2+xjlxUKTM/
eN7WQKT4E3LtiAr4Fhyv6wiDuXeiAbIyBOMt7B3n+kLi2GRn+Cc5GIbmbZfMtP86
363OCETVcwZYdoIdKF25jauvgRqii7dTMt6g9Ck6DbUPAYvV92KvQQgnAE8LZqMf
Zl+ISKozuzm4LtTMsQyA5oyBBEXmx6u8X5Dey2HO6gj7OPjNw9/MBQB06SVYMYdj
7oiF7yYz70EuwRujYcdmVjy/Lp9SDs3WzfB2ruPpc9NSMvSHR6H8XazVybuTJm7p
8X+f4VjezDHEK5/fIq2KE1tPTxpXhzL8tCJjToF6frrjGFMa6MX4FXBkA3ch39fh
RSMAsc0uxqdvwn8QVlzUSxCw7rNRq1Zgh6TvnCAiPFc9XiPCsAYKbiHqTh4m2v+f
Lx5tNKGdwWHJp8OHRhQEPFOxgIloIHbuAIEGUY3eoYmIl5NGovAE6R+iMwAyMXd9
YsiDna6lIavLgVlAYJm1Dmkqg2/ituDke929rJ4p5U3Lh4kHiUCi8P9MrpeGCNIO
ZDeNfyf26zMo/Ao3Y0+4FJoCanMBVtyqbeJlkZmhd6+rDtcUvQdu96Xh60tdO3xe
VYJh6kcF0idjhfxzo3yCfdImFjLc6CmNT+DocHSvNTt4pVNi7UXDioYMrNKV1HRo
8gdYaGwU2Q3+D6XfWJdbyIOQtUgexyflY9U1biB7zcYEa0fgNM88/kWW7bKHK0l5
OzAtPWZ9ROKXlymzVauIle40rGL87GYAvWy0il3VZ57R0+vDENmImdm64uJo0ozX
V1kyxTZKZ2qsyyJFZIYSjxYfzx5eNxS7tgsKEfezR25DPF8jzGkxPOv0w8OaShRr
6VoocQZiIX6DzrHctoZJcU5ZQPAzz8IaLN6ucITSVsvHgW0o7yYmrBWBKaBU9ieM
WXyS6M7R11ru1p/d65F4CsHTa3PISW5Y2GzBQ/coMuZLOuuQT0FgUr/qHU+Q5fu0
owUD2uG6hou5DZHP5C9bUmRP+qLEiDU1aPFLYIKCPwRyfvE++hlfn30XsUNS4bFv
Sem+fVtpzr9UD4h2AxaqwEoPGtIy/4kyfe+vqA6X4kt4kND9cajrPrXh/IVXgAeg
EPlZPGV563CryhUe5GWzGXLB/WaahWW9pXPfJR+ij1HThLnblc3ANSZmvsG8aeUF
BfimikWD42vhwbD1Njs7z+BqJb0Fmv7fWa2p0ELNhaa2QBO6t3PgxQJIhl7QmPDN
rIJFJ/N90uWmsjh6nDAsobaq7Tiae0j0dzcxMTCjeCT6T/48W8AgmQgH6KGvcx0O
DN/Hqz/lOwShy3b3Tvx5XavU5oEBkNmHFKCoEZw9D8JDV05zn3Lw5YKr1z8ClltZ
1flAw++OvV9ilCvvNF6UCGB1Hfscn86PrgxHRbYo2e4PlVMgMNukU3wUyFQzpN5R
m78me3B6N8BOVOgAUlvLg13YU+H1R+qDq2wAD8tJaDrF0U9iA2usRPI8EuvH5PrT
Y6b2o+NBhk8sMeGGbf9krXBxIxwar0boICV83kE9/vOhbekZZOVjzjOvNgb4onGf
FiYvMtcdAntOA7HSFyyZtF1DU0Ys4jTIs9fVh7ucKvVY0YFuDYVyNvCGZLTOOGGT
PzFahGOZbgCifkhM6NkXP94arE7Lm39n3fyLRXTLjHHLDySMtVMC5612/7EuEJYN
o81oELv/SNqLyL9a+QGOvkR5SUQaRM51x0oGcwRJyHB5bkBTk1cEjDz0BtygNIvl
Zx0WW8/va8oy0xpBZPoX5MUYMGPK4ONEfuwrfADkKybk4U8tucxDZV6CVVCHaner
JGYMVpNMK1+VI9fnqeHl+5OlllwzizWrsFEbP6WsOZv9OVb4oKyguAmJ5+xAVnuS
rM0lwvbg3PLStSQNIzGBzRn5AOQwBDfWdj0cSaTv4qGO7lE0PkIL3E4y+FNmP9bf
vIRnCGDGel6/o1l/LSIKwKaoaezaKX7ZNtkwS/mNbHa8Ns/Dei1lw8BDVB5LdBMi
gnRdijk5SjND0kK4iU+J0pDqavOdsPQSv8BhZv9wTIecHqR5PJAAjsW57nNLEuQ5
CBJYIcJTc9CUtOTff6hHMdZ+VQgCvUbXdCJxrs2ovI2SAVgPs2JyvcjJxxrKRgUR
CHkZ+O9QyLMvDYerW+sk4tU0CjApWB6VvJUEcXKDyQ1fiy6i5Krwa0m5IbBAD8ct
w5ePExd5NMMiHgiU8XxA2WGgdA0F3H2tDTPHIb+AKIk6IbYDhbW/Qk0y3M8jj5jZ
DFwzjEHfKfdV5Wv1u1T8xdXVlDomODtmeihhu5prVa+HZirDCkBKY1ncGjOsA2sb
/sfAkUNIJgmC1uxwPRAffRqKXMXSJuwYSZL1SNkR+CbwcIKUnanHjsNWtEnrlKHT
Tm54k6nQ2eQ4U8URUE7yruBSN1oAybRNrQ6mMQjnEZfLJDR+a809ls7xhgCpdEZS
jPKiC8jDrOrJ7+STP5xjgccEG8O/0rmc/tNzqc2JcHXhpV+K7KvX2fsV0GH7tVof
5wbW+n5JudLRyfAz3MGzA0MHeB6/UQMFzUWRYRW9gdBNkOEW/tHmAzUvoIUs9LiI
/1vRXN8EzCp2FxLwRfk6GJRw2MY4yS70Yl13AD30p3IpWzzNhL4aAUw2IBmsYx0F
ljerJy2QLve4jbqJogXpuX7lbHlrXKKq0HymlqUhPzGstBkcyrJG/NsJ7fDUNsBq
eIygfu9wliLvdZPlphf9nYErryUWz2BDfKTcmd84cNErQ+6mm0G2RRCjaratMKCh
l09G/Tke6ji1K5UoMEC0ApRVoM4OPV3LhSSgNNxPG+RhQmc7Y7Gac6xNExOOv/8a
IeO1EANMfEwdbSAp3uLwFSbmDV7v5BjWzoP5/YvhMHLEtG1pbO8qecRzT4c42WUa
4BTmGC0yJevradlCM3xrwOIIapjQ+f4YxRAEaf1qKAxQSfq50PPR2sjjSeuQg+1l
nSvl1hDk1bRIzyb84X1dcFPv/Qy8+wjIDbUiig/xTqih++7UrpkPDHojivYRwJOX
Ke6jnqA9rAFOTvK4QQ0dCAJAoay7TN3HHxOnBIJ3FIRxQj1YFYHBh4vgqZuSmD3U
0YGt5isShjFwNytCtaKztmYzWUrGvTQhIha3o6GdQhbwLDhlU35REnMf+9m60i+N
9zYBCuH24+IfgF0Xc1ciRFgvjiSZyRnlSOEMEKz/2Riw6UVaNXjd3n8c+6w0P9p6
PdshsrtNdByle5wFs2XHqnZJVVHzRLkRIdfk+IYgEaAq0ntayorSSJTU1JnL11ZV
0nvjS6x9wFceQ8lQzGc5jWa+GV+QmREbKyVKQ0D6Vc6hBgFs8k07GRMIe/fCbohe
UcotlRlPhCLGsap+26MXvoSQ/55YD7kO48ZHylwKOBeMD0TOgIPmtVX5q+ex2M23
LZjrDWrawm921C2kXUpNASeAY1uQkn0WMK04wIh7wHbVYSiJDI2fC8nG6jmKy5mT
J34Bwa6N1MUd+/FfwgTbqo4b/aGfiHCVdSgRejhW2F3rvbg1/BYnbYOgvwsVhMY2
p2WcKfqTo+KCNk3K4vZuRDDjk83/zlFPh9HKgqch6HnPZpddFG91bd2Kpp8IeGKJ
N40JV1Ky7CHb0OskCQdBZWBEvSncFaNM0/dft6M9ULLXFqRrfWXf+lYg83fExCYi
1jQO0ERQdBJAhOw4vLdv62nCOecTmdB1VFpQzajLqiiXRbScxq6EYyB4FfMxRyvL
WslB0Z458pwOteBvzc6+dqUc0zQsnMz95dz0U3dVXjI0gdhklcUk5fXZeG8egHNO
3CVDNZlMmSsyC/G/KLyQ6T1ZqHMc9RfR4b3F7FT0550pERCJ17rE5rFvkvycWeu4
rTTWZDJCdbYEijKpJ/esFu3zZqqff2runEzP9L0ghFPHuDuJrng+GL1WnVqL3TT1
XidK9PI5rkSIiG0sc+7zzS87L2j1XxwRAPuUCZiOnpiBU/oq13Ug7tnrC+YtimP7
Of1MAKTbUf07PbahUsMWkcKLz2Kj9RaWcxoIk8gIctdtf0hBybtleFLlEAA8TMN/
vU2UpaWWHFFsvAdc4wCsuglgCIR91p3DstAh6v8RtOcUvu+jwQMkx1Pt5/0WhDG8
zlDrXtEsx7nIHqoUnGqK5GfwuOaqvQPqZc7SDV+y4N+G1oKkXNibh605SA7lrqbS
cO2yqbPZKp+/+I/agT0ZZMkM4stbQ57Asi32KZyrrQab8W07PXlRsbA9Yy5VGFe9
ONwzaoCHkQgChtOVQPzB1N529Gsh8sAiTjdphq8UWG5bH1UqXIP9N1OVq7AMWqGB
mpvTulmtxH99LDGRsl2kZjudDLoUK2VpXP9tPqezMp7XbT5P2GD99KbQOzOKguif
G6WCoFiZfSjtQjE89aehYhT5mynaedBq+IY23FeIm3A3wO2apLsq+OWbi1PFE/WG
TZOSVpJlWh2BX0hH/cFO111CEWT4Nk9BvjyqDobkDXhFwDS/FuzQtdGHz8JG1lf2
Y3L8BV77JtIuDGRSaD7A8hBnTpRZVv8sqFPbXCXcpg8aa662e+NByIr2N8BqkKWA
r7Si7+dORfZfZ2530IQ8pa8jQSbkP4w6ZMxr1dlqaspas68X0bnSbAJH3ZpUEdyj
neJuQhRx1OxG2Y8ft3dIx5r2+xBpbk+8fw6m6duQK8j/tOnGhXSucHiZi1rnN/Vz
9CCeS8Wn+up9ARn0eHt8M5atOT/mDiyEkGuCDrHCkxZX99NowVMjVZ88+957U7KL
ZUbOlPRvuYeUrPPVphCduBblqTb+1/2PE1PLNzdDYL83pGlojvtN6Ah8ccHNZOn1
3oTeaVWOjay4F/OVT6ysYuBIvcK3ZHtytC59ujZNdN19+c5nxAEsO5Jh4sh8wiac
TDne7LDE6I/SyNurH2yGacZFfEaZNAdq5gPmsIN1ywDQXus/JSwEoZhIOWIFNvdm
bxP/eCPaMldNqI+8CWa5F0WDsGKt08PMgdJ4Jsh/F+hxW/TST/nr660uot2hw+Y4
8B3eg6Q8PI/fPVzABXX1SHlUdE0vu05IcsSZlGWUPlEzVCq7m41so3lAdZ5jVLqM
EGFUol19VUGEx2MhrhnIHqIpwoM9Q4Ov7M2G6GUky7GveNjNVGctf8MwsIM/IqmI
5Mv6a3/gYpB2gJaMgLkGiS0Z/uKs+Uk92ywuLMIevJUg3C1TEp4ztDdQaTmExEkW
sGoI1rQBVuJ5I3BpBDHErP+tVlRj1iCGAoCZGLxr1pCmNBtr8CiEj48Xdnu6lSNl
UEsRCWqVaaBTSiGdT14RYx1Td9VGCyXHo45rapfN3CAKQyStIB5dmS+JnwGCpdM2
XKmOxlYzV1tBe6MNG7dcdLjwrEXxbw+CZLImhbD+YNNks7otadica7NUzjK2vlrb
sNHYNyN/ue/d7FfTloQucq6WFF0r2sv0I/k5QoXGq5XprxYEdifExSUNpa3AL3QW
bEjyBqZLIcDt+J3GwGBARB07F+iK3LE7gEwULZjOAg/dIwPtVJ0W8vwQy/isMa9D
9+HYcdNEnJVXDFfJiSxpqJxhOB58kOiPyyTFEIxvHxC0dIJvFWU+YnwOV6dAOnLW
z24m6D4ms5M66Z56Uc7+gqgu/BCXyr2hqeh+k9ZAzWxDOZslywL2Q0h4I+FhzHAx
i48wVNAnsMxMh0z9dnZ2a5WYBtkkcS5zdciTCP7XmP2MBonwuR6K813TaoA54sOT
3/AejcvIuBPlg0Q0VP41Zx9g5oRXPK0gU8VBhtmQA0O/2yABN0rzD4Tz4/e4RN81
WLEn/ZHFjOajOkEMitDlQx71/MGdHqS6Z+McMVYh8EzBJSyrE+hp3Jwcy/KHnAaW
WQJ20jpmCVmAwz6XVNCvFONAACLy4tcs38IjHWAMjbINCACEp+eYPaAkoqYK7o+k
gH/Mzd1aios0br6OD+2yFr4sgKwRFm8NAniXv+r5x7OZpKfZWCNC5qtg96dT/eel
wLG7QXPdk1710IlLCDk9a163vrsPCn1zNd4uy12b3HFBWwtz6QH3Rnx0bWyL4tGN
ov1QzCXIoFD9UTb/HHnI/kC5629qwHrQW+b7utluAFnSLqqPvjKgrfD6cmeB9XL2
5B3co7OPIGUcQo5SBU53jpu4vi41uUC28aO8iuOjnuzVegFZ+tT8uUUI3NMpk7hx
JKpPFpLX3uHaSCU5XQ+pXycUd25HKlTk1FBSO+XLftYOKrXhH+r7/5H2peU5d64U
/Tw4J1VzXc5l66JeonMzYZt3tZCthOxhtbYZ4mfPtEZ2TGWS3oyZ/4pDcbBgNxCR
1nqadjoM1YCGrny8Gqxyn2UNRdN5TaaQKvAg0Av1dtZ/00dQAeaQX3aKIVnGdGTY
ummzGux9gpgks2gtWXPmuyOobS2Lv1isBJTibsBdKUdoyRIqWMQAbGTdkTQ1Wrdf
aHmvuirpN0YqwdiLPwXzOoZKslJK9pL+5FH1jZ0vK4+7+1X5xKmih172GXNwczIk
GJObZS1grTEMg59oWcHD6p4PdjabDzFY9Z2cHE4R2gstwKCDu9eBjXP4evyS1Naz
vprB5bt8NOd7ceFwN5mAuAAPtgGhviQjMC5VucJ7eF9xeLXrX9fHpBMw2A6vY0tg
tkOPeYJ/g02JWqMwXeEktKS8OP4hs/eM9yT2kMmeLcQrT+5W9Z8/BMRujkZjWIBd
EaTzaKkktgcvjy2f2NO9sSovyMOfXqXserftShw9RCkv5YeAQBB89OqCWHLHcHpb
1/SF4JKwhF6A5p83HliQeuE0WW2iE9wprSCS9ZvWiPvsfYZB3gbcDYVcKrNWXajz
Ebohoy5MsS20hMW/DOiSFcOSoNCH5gJKYi/KgvTv4mWRIpN6NDy6mnneO3ej0Y+Z
h94estHntXgIuhwf2P1QNIuPYsZn7R/M7csgni/lXOpD94n1CSDGMxyojI7witCi
Wey4iNjrHY1wVKSM5JQTV6TNTf48xZt0cDtOEFq/30tH3lryEsx6T5MYm72MCYh7
3oxC/xbmaOsuryZQuYmZQ0wy6xInJLaWuV4zYO2FyPJPmit9M7h6JVxm9wmT3Ozv
41i5wpgpJGeX1XFNWFNLZwuH0UtibmqeB5t8sqBj45LFIm4IESsHrsyyCI6zT5vo
T5A483hTfEV7g6Ge5F3TRtqU1IfdV/qLhzLm6E/7qfjgEejMWDNBUkisC21IoFiO
D7iZFdue1+Wq8jCg5rZ2LC1XbAPBjwxgdsCnS8tcF610KydfCq2XojLnGUqjeAaS
XjDZb/f+yQAZox7bgajXgXc3uAec16Hl5a/+lpC7sUtQGqqwXKb0lYXC8UA1WMX0
mbVgNCjGNaoA8kicocjuy03K9skp6n5RuRUJpxo8i2Qtt0/glwPRGYDMTr6c80Gk
h/xwBiYweK9SwD2tnpCG6JywrsqOKnlCIQBZG8Xae0W/o5Fv/xg3+qps8t1Pumtw
1TmqKmQwtxvXwVDK5uSAmidu0PFxy0yeUCQdEvEKVN+YBByf4Tug783Uh5uRpgOM
pFnKojhBr7WQ7QhYX+Uf+uWLFQa8+nb2sDEzaxDihiKQM9c0enCLC6LUmH0m4paK
JAIuXbLMmn+21RxkRQOJ8HZbDknsUjEmwrjbyxOQ+FJ3PSFkBD48+C/FLBIEccRn
UcvtUgQxAfq5SUSgLit1DSiOensCAOwqoBD8iFEsOBK282KY+N6P0lKM9N8uOP7r
WK5rScZRallibewjcfmEjAh9uQAOFhRVy++bchcuJcajZ8pYoFdb4gOaS5WeG8g+
HyXmleZB02fzU0sFu4wqGv267jGVGXdAmbeHVZ2QIjpKTuflM9a5CnuL62SPXlgl
DqzESASVTxOVImZT33Oe97ItovdA80iCct3LxYcpDBjRqnqWXzUJWJT9Q6dI7jyB
FQ3yWyYKL0NuDW7MFUW6vTd4HpIhMZEVacnWi0tdfwS60qtCC77L2olbt+TEsQWv
udRaPfUdvHHkmptzc7KGo4q431X0vDL0e5jvRVS4cehoWE+oDl+gLGDv7w6A/5vo
4PToZqihfy0/PvFXYmMtbue5a8LOfF0IsCLLhCemeU2h0Uf6JGwwbkkyKBLifgNP
Pn2Gm+derhbABuLBISdLuQOyzB4gk6rU88DXWbm6IL/ZlLfsFtk0vKzuBn5U501V
FvhDdNbaM/q8YsRJF+7qvA2+DVdFvr2KIQCobk8c+G6EfpR61Qa+g2qL/VaWBI2m
FEMjOrqa22+R+KG8f4LLQ2nARDIoHPDehhaIXmMoSFtLULQPTl6JXg4BmUqhx/QW
Jp1DGcaq1NN+wrozggqjDq388mvyl7pAFw4jVO+x4BccsdFqcTwNiGYtHzP8uThS
E/flmaV2mc6+sTUJ3ZwKVvfAD6Z394QK9hxtAxRa4Fz0R2UTs/LU8ux2qkYW5+7Q
UmjTflR3upwW+beT09s2Y0mVklnRB5fFuteqcZ3+joneu+7S4WHso8gZIkQZx7Gg
gvK2Obft882AmqSSoxJwQUWdqfliYOPvhYgqH7xnWdZxDWNdd8U9AkaBKP1GPiaM
ksgSylgBgRUvkjrpuzPO7oNpw2MGWIE8J54okB72JiOA0CDXNHU5UQ5/TEaE902A
LXLC7sv6VRlIQXvBHnYDE7+izdLr2Qmbjfx6iZAioi55PZc8zVPexyBQPhuE96k5
tcpCcaI4oApIy77KyD1WtDvYTc5QSpb0Ju91tfA5xtP0WJPQ7fczXS7hIJZisbr6
tUTbYLitlxOje20muQa/FPnW5Q9/yVIam/l535vV914BFW0+wh1fEFO0PxnooNl2
fvqo/GtxJ6p9BEnkrCnG0XuOBS72/eQ45v74RvR0Zw1cL08uwlhzncDYGt7LmlVm
D6Y18ryGf/c/RjNCphaebyHswTUke+qMZhIeUGi0Jxe+ujmxQGyL79prnqWh7pje
T8i72S8+L76c1yOvC/2RsFbnZgwjz9K/wIw/R5FtZxUSjIqlV+SBj3fmkzpcPeai
8xKXMICAYmTX9GgpJOtnfv7etU12P8oSwGjFDnzlToupNNho28k7C/1ReM1Xrwky
zvcXosrRPLY8RfNTrhp9ErYochGf/5LPCm9RNmOY9lbqNFBuvraPei/dZUQuSdtv
FcfkOJ3h2i4a6fu4S+y2vWkNaSI0E0/B7FbE7zgrinyBtuWEsOYTm7TuSEv21OP6
8+9EIsD0sbPlLMViuFm1rzIIvLFFlwFVH9YNuo/lRIyvcTvQOtIdXjC3CyvWvCGA
jKwDaWgGZ/7iTDWkSonopRmecFpaEsW4JHDQkbod68FgCQHMjZsbXMZsTuPdJURB
wKPkbpza8F6ShDS5SOBz4hFOPXvjKSdaq8mKSKuVy+f3yiveSfE/uMveq+U6M/55
SR1thwKZyLE9eHouAlLELSP7jucBeYEdKcdevitQAm5yKYMHJp2um6Km3JyuIwqB
opAPDvqWo7y2oenHxJWWAFZq0cw/HPVboK/XDhENhan6OOUU+Y23Kqx3BXphCMNc
CfIbkTpGjD6SopcL9dqr4U+XGaPIDo7uLANuUi0oqEoHx2NYO1WLLhiUosZzUUnL
1Wd/1JsKKe5F1AUVCPqOTVqNkrA92kRyW1Gb1Dc6BhYMdAzE7wwOy+S34TXFrUvB
m3ONYZODUk4IYAtIAMM7l25tY4eTsUdLqXb7rRPnHj1G0pjujZRR63BVRe6oIQFm
adolqKYPynxukH1EIejpoxqKEA3qxCNymqpGvIywpPoeYTPlXaWJz4N8Iz1yfrEI
x43O6NiabSdep5mLLzDwuVvsfzFNaEp64zAQdJzKFrkd7yi230Nodg56TEdUstw7
FdAXD90nIgeNkXn2Z+PdPb09QsSa2n4B7VF6rcPLuU/ahtG8sjOvvU3lp7oAVVsD
cUo5l8wSWvKGkTvb+kystxR+ToPg1TsbAQf47bXSLOZz7ckmc2pFxLYAmcpluFZ7
6cy4UaRxEttUHnQE+xN847zyXcY1ymAT91IaYQPLOld75buzHVO44xmNQaeIRQCk
DEUyXTP9+67SuFY3RgHM34JgaojHFo/pnnJ1tbDEW/RjKiRjDGhiSsjl/4lSvKeI
1cwFbgs8PoQ3SE2WDFg9lxelgFAYFlqgBBcnfAQeD1Lv5OZ/PsodZJPj9CvwoUaF
AMxLAQanJOfsLhFny77N85CfsUrQK3xQ+X42e/Ql773EmmsW2uttg/EljidVg/s1
xqAaqIehOkUlcdhWs6DKV75PtikTkWS2scGNKXAU63IU5nLI6ice8aQ56voCNcUE
vhIJG+xlzwg4WbLkZ8juatNDWMjSbj86Y0/rPurgPanUTbszeMK2SFHQX+GJLlH+
rqv2iUm1NelmV+pd0vIOsGVJoMUffSbUsKw1uz1KMvrZpOH8oSG0Ow1/VHzmm129
OxCQvyaQSt2jyLlLnuL/CDkU8yfC8jC1bZK1TkDUnp0TQueRT4pgrhWdTSu719as
36MhUZBaThird5D/5kuVBryxdJRW7T20YWD0sB6zcLcpXiMppaQyHzIvW1zHyOVE
d6p6K5fSq/igoLFLHABWUQtIY4fNumfVNHL5zc9Yx+OavR6wF1G5derNn5a2QThZ
jG/BIAOn2f5RS6cTvHEbt+dpi4bfh/xJYz4dbv08OaO8v93rllqNQVzxrhuFaPyt
fBnGdc2AcHikJ3fhUkZtCRLiOsLCZONj+IWCcqu4K8k37mzxl2/0DbX1Xlf057PN
9OAcJ2lnAr0cABJFiWT58OqvdKEWg9/JpFm4BH2kMvp/ihUGiqab70utTZANzjGF
ATMzxdI4NykYSFLdTVYid/MQW6mij4CQ+daphVZ1pOERwTT5Mjc3lZKxFSAaYgLT
nE7oaezT5mNNFI3VTP2C8tiyGuVKahSCRG81Xj51eNXVBsoZjFoDj7UW2dkT2vXz
Db4My+30oI3NVuYKNM/0ifr5odGWGZndEZWKAMr1B+E2v2hFoRJRYE8yZD0ECT3W
SJ4Br8UWe0xHVtvb1Xy3R82idrY1BYTH2F4Nah4mWaqGKg1iCA9dzL+u3RzdtNjB
vokCj2HfFtOnWBluiusb3324OyaG3rqsic1aSaoYDMyOML+GqZnkhZV0pIqcBa3F
9UmmSX2UAz+R7Szx17ZHD/F0Fk4atyTAAO9cNt/R5glBWiinI9OnZLGg+web2tK6
0x28/Ju8SpiXlRiWiklfKG37cBFmOB5kZQhvNs+rufDmJ6KPSrvK8qhENflWu44c
hsUqu4y1rE7oP4NBZSDb9ZcrSGblHk7r6calEVW5UngN531kL+ZpcuOB6LTGV5mX
mPOQCYozX56ixcQeRJ3dZFxqTWnVIWXOQCrsrm4SJQEeMDi+bso/MoiuzCy/Dx0/
ym6xiB/+axmO/obJTIFb1ofhYzNCcs5Z4k4mP0IAdX2V9qihRN2FZRV0ZBb0B11t
W/uzqA0Nxtz2d0ZiXZaJs4yzjzrRF9nyR3r2W5if9g+JSsnN+2funWCIooLyAK3Z
xhRX7ZkwBI4XONCnXqqoFHZA0M0U2CJSzb10TQR0BsyCOUUmuPsu0wocLqaQP47O
TvacxyGbphL0ep/etHKGFPbN5r+TLYr6Wlaq7nuG2eFxg23/pQ/uTmz8wV286djz
gdyb80P53Z3zIYCVxsSWyXrEF7M4tauoQmWFEkE6sDvda9c33S6N5/Tm3G5lnx3L
BoKaDtvjZO2coo6YcLLJuCdUfD/hKY/uDRqietjkVYqYcAsmYVdLRAHy9TK1yfTz
09+6wGWjVwGzdEwffS2V194Udfw8+LHt+kmwcmWFtR2VjOOP87e6c9CuHp4VNjc5
EEbyyrMPNVllMxLgTe+JTo/I1bJloT2R7SGsVAj1iWyY1fh1aitsBGH0gATbuzwA
99WPxxFwswKD99KCmPTX/Pn5x5gayDHqxCCfZxmHabipgr5aOVBr99pFFA5NS0TZ
OZyZJ67fuNWwQjNfDQioW3bMJCblS8PXFoquhsaGacSv16yjf3XJTGFNrxL4uYo9
OEOgY3m4IcYfRpSosoAajgKiauPQgLolcRt++2yPkrVUosvbMIu3GpKfLCq2qgM+
wj2yg51rooRfvwizKYaHYVxaDpGU8KzoeA6Os74M5zDDg6OFdvu1s1fWBlQYJELh
uaYzFM3uQA+cQDjU/rfaOqFIRf9OncKfUujvkz0mxpzBH27+4pxx9wuVb2JAShE6
ROBjItytfChbDQ8op6YPCsRRguY+S2rraY7vz1wnbqEfl57dXM4US3B7dep2QpIT
j35IKx4wjfMH6UAQ7VrnRD0Y1kKbPWl05/397WQQiyeik8CvSbJhA7USe7OmuurH
6ei2iuvlh6jFxj4VqstKiGjd5bVf8xxwIF7g0/M6UJjoh+UqNkCxQIm3Hliuh5il
qZy15DE6CDbcgEvORp4xQh+ujkeUxl5MiQDAoCfd+/bnu6zWwaaCCZaCV6kttcM6
N9a0H8+udDNXUCjalIq1FdjYwQT1gZ3QDXvx0SFqvSkH3vQqs1zArSlf7Q6mSjt6
PoFxP+51YaJOscwfC1d8Jt0ApjD28MLI2k1nEun5DAg2uE9l8T86r4nPpi6ARcEc
WojNt/fsK0tGG/dXLyZn3OlvK9hVjsRXJ0Cb9ylf5LGREdmlRK+3/W/r1OeDKP0W
HQ2bRtuAE3AEGQ9+yzRFn5QDz9ccj6OFU8R7I6KQB2aYx03GQ/qbAxLG9AJ52wL4
T0mQ5h16+aH3AbIuHIk3X2HEwNU2qAQPccAjZH4Pcc8FFypZa9MSgBs5W0T76zKy
wWVnS4GwZ5/6ctQT9E6iLe5imZfopLZsTkPq7s2WtZpXB8yeOlmqGt3QV95Xamag
fnaDF8kdjOPBg+IGjKaUARXsGS9NHdvuyh2A/OO5B6WBfEU7fCZAYJO8fL60JoMl
5LTAKyF3YgsB4XkBHmBPIQpiPoOczXyEohIj1avbdhHj9NSW35bTkSgKaCW+QKr9
cj55oyXd5KsFJQt+aaFskblznlDI74ro8PniWv+bEtNbxjEbXYTm8pLh9lD1iAj9
rvJ2749qd7SnhI9hOjIjz6TRRSOecIxeYvzTvtNjZSNW4/xzY6lFpEsV2CMIo2v5
QTQhqKwYiXO6DA13FqqnASJ+JtV7s34ddX+qOSLbC4a11kJUgAEbeSxNWiXuNlEQ
580mrz4AkjNYclhN/XdYmHRwOQuXF8IYHtCAmEpM2awnqW0t31YwL3LD0nf/sic6
2rTC+aMKfSPDPBQQVV+7gqmqR9dRklZUSOz+o+cvxkTLMZu3BXoCiphl0scgU4YO
X1CjcIsbCzYLsLPQcGJQKT9rxoRIP+5T2tzo0AR8d+xPvvZxzN2h1doNmDbT8wvS
sHawOz2bnG2Kj3Gt32bMOuHWWlkTu12ZQDpckS3rxmo6KZ3+R8ekrWRdUZiTkRV7
SjDZo2gkxhjLnPKKDMhf71x5n9A7+GEXuJgpvcLZSxL5JD2hb5eQCGN8iLYz+1gy
R/0p3syhTW4M0k494apc6Tf/5VfAdC36Vs3embZDjz6RM2Ch9kG26+tEsXo+cmMf
KoFmmi0EyEwdfcGLZDJCIo0WLXjRQpLRB4BMjXtDagKmhcwXJFI39txFKtcMp5NJ
lFwUxI/jPHJ4XE9cLEhj6FLmejc7iXGc5mWOps62Vv0kTi7+2c/2I4ya1oN7nd6D
xdvpzmOyVE1P8/K6DSta3JlLb07UUKeTupvM7hluXK1aTLkdM0pYflZ/dSIiX39h
aP9u2nCZW75YQnv5MFxWAL7dpjvpVM5zOXtjY9Kx6XY1Bfgh/l7jVW+D6+Cp9CO0
WQYwgzihgMdJ2q9ZQvkvXo9GtU/IoEikC4OPlxQaAWoZqyLtJumxm0xsToocaClG
GRzn9XPE6ivfV32oQUg38p8fsLAKQ0SlwdARzJ/WaV+cex8pvU/XbFLqnOQv52/Z
KuTVjPy3eb7Ls3Bk7fj1MOoY1zBNoA7ym7ZZNrmp7WExBXS3JqsBlOHWhqA3vMeN
xxg1Uh+ZfddiYPOb2dk0lUJAfINTNykHNBtHSRW7UjM4x9BnAiGLo18JI3JN7SWL
XUhZckuaXHb3xhWnqh4foSjisZqvWtffU3QEbifIQBIshZ7r1K9Pk9SDun+yYGCN
i3jlJsH50yM10N78g/6g10dmVo8ikdFwE67inR2WCfJlXQmuYLnv0PSqh/m4WiXE
uY5evfrMyVMUOzJSsNwe868EyRXqEC9Pf4lMGblwqVM7ZTQVWea4P2jTI58IYE9X
7sCC0ohORePqp/Ypxkx3CbjsdgGRSMBOWZuz5zBRH/ed3jxmovC5RgK9P+5t3YI8
XRqJmdvr2/v53X2NkEtJEzEaYmYBsGHu6AbR49OfQt3lPF6wvojqFuexrElzc+4G
ziXZIzRuPaWJTKZfvTu9yhKG9z9RrnPgFaafw9jY600QDuEZGAkgVhotLLhvoxLo
gSvgjeMf7aftOkXpOYsStf28CgZJ9fVrk68SyXS98025wGwrfsrmrEumuvhYIJlG
EnPQDuHwaiKxsBCSl3qc4mlpbbC673zoSP3TerraoIF7bJaBUcrrTUkcnsBgf7EX
44ckr/TSO/xZBSSHZWTeBHd5tP1nyuLVIyjGOuAWdGIS0lldkHp8Y6L+ho7N7JLN
iSRRPaGDaxoGbXE+Fh2rKn5TOI0UELbHzBmw3d787dpr23lPwUA421rfAW22ob3R
cqYAgvHJjtkdhV7yjoVZrtP95aKLPeBmnbExHZt/I9X3m7jHKq7UgJ8VxHsgnzfM
vA7df5rDu/PHpx3mEZToepxl7l8HQCZt6+oy8Z/bsZ30SP3u+8JItxGe9q1MJNDR
iH+MEYW91OgY63scDZ0x978ysbGsPgdKQJyOUciOPM8ilpkTZrI/jRR1+yUsFtKk
2J1aUctMi/+OoDaNg4NhwJOFprAwK3W8Ywg4lGmPFt7b0Wic98l1udAAHmNndvhh
4kiop0ktdJfF3Lvzf4j4QwytrjjBNe6NXypSG5G5C15LYcjMKZi7ULe3i+RgYMaE
R1u+OprY8QmIWV0+HmjA5AoxH6heoRIVc34q/uzrKReLTGsrjM2aRM66OLhIgXwj
gGdixMSJXUnf9WrOJcXjqbcLTvdyKXBBXuiw+L1buMtbr2l/suqUmvoFZ1egdMGx
h1q8x9XV+ATdQkcT1vdxqGr04rQ3CtKVY0c4qDqHSkpTZZPf2NhAU2lWPnl9kIUN
4fsGuQgTtXVDPmTnk1LaxrAuiOMahaUTXuUgg8PloAWZHh3GXcmD7emlIsoriEMm
iA8m5xkNJm85FTighU8F23pi0cKJrD7ZNu1lb0poHxvQ8P3+N60BPx7GTuFAzXfK
74OQAFvuxPVJQuV8+S5L2JZkT8spDOXjl70uZF4nP9dGT68nLykDAINS0sui3kJY
3pqsDdzus6d5/+Sl9hEqtF/1T4kILj69nMvuRkPNEodnRPQmE6mpMqaWOKv8fMes
8Gexpyn5ncCpVwhh3RiHLCDW/PtsBDxm9s0uUiasLHiZqQ/TL9u+M5K1FMp3xlUD
8ycoVyUpVt5g7CSZ5rIFPFFrR4iNwH8n9ifQp5V9I2UflBDKtV0OMzcFtqoifsr5
8ArYN5Kbubw3B9TMETED3uJ/9PUgLaSKuEDDz2YuZetlRgAdcscSzhdh6cCh98K7
USykjA+64LoJhq9ufv8xHnfsxXbmb7BVOneSBIIofvJK4F6BPpSZ5+yet/FYtRZ/
t7kypOVoAPq8/ztCuN+WlRL3Y9OtAFJ0vOxmacTs4NeaLa40aMjPYk5T9/HCUpjZ
XQ+ofUTava9xwyEYXqgAZ8eG4FnqFDT63F+LCeMkJ8TqYgMw7TkbtnWAwbtT9iOj
Q5FZU9Mt1Qsk7rGlPA/hepaPwmRP0Q+0xp05sZJ20UZTE4k17kEjTK4tF1N1mIG0
rUg0VHIX79sfXl4/IaKNrU/zUP1T50VHEQNyj6VZV/JU+sIdE7HTDd6Wwc+o8y9r
FGk8QODFgzon2oe4pGTmj/4RSHw9pTqbOQulMaAXYDYET08eGJOax+30QiS9cmK3
g8U7HFBLEsJHsvCA8tImBT16ff2dBlB1z5gx0fZzSuByh8KIxIxWqjZVhoFVxl+b
ctpI2NN12miNKw+h5cUzGJwDTsL5W5GU1MEx+We+8CYVEyY1LLAITbd3FQ663fl1
Rt9cjd1hcPCxEJ52bwI1UkH1DQ8gskSfbL6xdatDX2a4/0DrPifP3mlIEY4pRYlP
rrfGCJnJms3QFhUMDp19da1PMu4lG6qpoWQCmZXv+bRQJQN7IAOqe4jCcr22zIic
s+2xsvYZFnP1ggsTtpCMdBWmkKPGHDw1TKqI92em6jKZ4frrglHX+CQCFMyWGsts
UKoe21ah0B4t5FS+j+ykf9UfTVeXLXfuTfttAs1nsInHD6pMSRz9WYQkMA+6cQWz
BXQUeRrdEgJ7SVLXt0wUJyzwX7r+bXQdxY1nBAQgQOpmTTnM7JJ+y1lpAcOitHIF
V+cU8lBlfWGmZ26wmO4G8FRBHq8ZvmIKLhCLGH35WZyZuq4NGmtKaItq8VhKl4VZ
dqYgJQwMAvNA891zY9eefsDP/5E6pLE+N4L2wiQU44FOlgQit9KAna5of4OMCtdo
zYpIA9fe0k1QAFxAMitffezhdy6Y5FXVS28ISsxJwOPK/L+26OOqV5SkJjT85NiU
BeUpOmoygq7wtpSYdxC9fGXtD81wBCLX3gA7WzzLvVifFrEBYs2jW4/bS4Ufj2Ff
aZTnoY8q1LTHSK58uWULW3i4c1sRJZ7ggFMJpMi80jc99lv8JmaYvW4c/Vd/2F78
FLjNCXxJ5kIKVGXSFMstBPyh4HDNnth/BIW0yciGe4KvJgKQiP4YlPDceb2QL/Wb
N7L2PpnDI2GH8JpoB4K3Vzes/sEr6PQrZm3nBwAY9a/oKDmrylkAg5DWaBXFAhBR
HOEdA2Jl1rBWL3W4vyQ+kdmgc8XW+ZubzheaD1Z0HV5mnlp3dH88JvAx6zO9dXm3
vrd4hYWLYGD7q9pRHNh4vnPufRJbB/29/w8Eg9JVxejCMXMz2dooXpEegNX8IQPL
VLK1fwfdxOHYGEStuj5hWKIOwRlbtbGwNKKHcSutYn1N+Rs+EvF1qpFhB5NpyQRv
gEY/T38W+WlJQYrEN1Z8SUVa2KzbwZkLmEAPBx7TAVHJ3qUY68MasOcSBvTAHGUB
s0Q9/M/Hpny64uvjWtrUcbtt7FPEy0E/fnhxfYK35Vx2P2CBUUoAmXb28OcDlPiP
0aC/FnJg9CxSk8tDEjokqGBb3zJouRdYmP0YV67mIEuHVldTGLKJposXwPf5V3oI
3bTNMMCyA/aoQmciQ/lHCHK/6arVdAvAHevrBGSB1qvw2vWJYJa92SxdDElM213m
G7yHKzlz3PNT+Uy2miwaVqqTV+Gra8X2trYNMllDmYbb2gpxYBZooV1q5TZ8sgz/
tfM1j5kJqwdixrIe9yA0JEISEm/9qFG6/0UI94EZ7d/FtkU2nhj2IlGwPR6S5qsR
VYKXxDN1Gd4HdWfofEptNeW8N6Sfy9QFn4VUFvLfTfHBUiPIenf700Bhq3yuoABJ
YZRB6KIqGtagdi30O0yNr/wGxr7jk9hawc0snnWT7sEICI7P0lB4xKC/XhBXZIpO
WeW6SC+71GGNQVpIeDC0p4m0dj2gr8HIfwzo+UHIhnl9AcMB1mf1RKBdVRr7sCDq
Oq7mznEFQucFsPgv3cFmJT/TjNj6moaTqm1d2qUTuIAUNQ8e2jejePaKhPihJjH3
yF3dHZdkHQ9sBi4Gl25i98QEX3mhyurnrccHfDEUHel6lQvK40SIw4XyZJgmYQKO
H7n50XmA46NULZY+FlHwR/DrY9lj7KWEVOeZGR4+Kup8JJHnQGvVE21sktBdtd0b
ofUcMmJ1iHn3mhQQi4mByTn0VndOadMrk4Z+V0stCZ0TZP/kfX4ToxGJqN2TXHYL
QWlvAh+6W+i6Ijt+GJKixmv6bv6GUQW39CMMI0yNxNxrhd95ZAhB0Sz708vzACZF
6NkSJdLVJG40nq5rnun/51kcD3pxeUJgGco0VdtaS8Aqal9ESjXrEqvJXcdOwYok
DfAdCG62OZomsGiaFHLl+x/7kfR23cIbclb3heqg8VrhYBbScOBrDqfCtKoODgUZ
rWVIjaFOl2yrWZxBkuc3DMHxwzMsFCHc/G6ty19yeG2daodod+h7JbR7KvqIBRAg
lsx812qN5MRXtBSMFMgqdDM4Kwfa9T/t8CsKsJv3k9zvYJ7S4j3atQ8kozZvsu7i
IO3eHu2LTfgvz3knt7uVkDvTP8TM16/ErVKQtmf1J9shkayTYaaHSt9/4JSzrD05
i/immGHT7nLYy1C8AZ94wcBn7w3dYt5uIRkPbyQkihtbPNqa5vvkpKKHdc7t4PWV
b2wwW1feuVlseZ5KMG2+cK26tAf6oUDpi+r9bMngFXj/tLffzRxloN4Ak5xjnCeR
pKLAQ5/CovYfIz2r8K/4atzDVzXUuXNGMWhj4+czBS6elece/t+KxCxGtM2j4pwQ
ws5znCIYrWYl8nm8x5pUpaf19PH7rDZTDZIEEB9iVlFhsDZwJ6JK7brTPPuwg7JK
LdxY12DB2NHqpYmJSRsKHl7AtyjyPghqieFutAPFRZoYby0WQVQD2XGzc3DTftcj
m+jXcJWK/icbKH1PJ7HMFZBQ29aY51teW4y0vXjVrjFMIdzXonqIya0IhcZb+ETs
dKMyC2FfgnBdBbz29CWTqAMoG39bLnse0nMDOw5FLbs/rj0KMnv9Trr3IAc2bZir
+EaJ/cnOmuuIKM1gOxnmUYIu2QRpzOufy0lR5fRjD0IGRLFA66js+cqSzc9k9r8J
tEdxB1AY5XQ3YAGYIajeiTzIbwvL2L+xcoseYB2qJW1l4NC3/addY0BuxjivcoEj
EjnlTF0dwfofnvYjt72EXPRWehy0VYIoGUuDASAtCFH4IhFvSkeTXEeQJlFPNOo4
jqgA2mMQwX87wriWkmvWNnRdigEuNOjPyoJUUbtuOGzIpLKzqUeJqhvCm1Ygocnm
LUW+Ios6xv5VJ066VrdMItI8NHKHsiQI1NZeOqb2d4xo6LcpLzMuBimjCeRTFjhQ
siDyUyNZL3f56Z6voKnaRNeTL1anNAWVVBdaIaItY3XiB/aaVuVCWoEV3AdaAKav
ITUyPXklZIW3wcgUJFspU94rpMNfxhgD7onp3cW43tKe8h6YYhq5xI8ZjG4AnpxM
3wdqfgngVY7WK2y7YGdlU+w1sSly9g7+zMqUC8kgZD1xT33hitLFERSwQsGrqZ8e
ebfDm1j6YUw4qkQ5v8j7hETMjsgpOu2ImEVWhYuuZRmo2CaL0L/kUhzYGiVbvPff
Tb8sAUUcQTSwbkpipCgf+qNfIQDTAUITOhBKetcBtp7fv4hNpVpjlyM01HjoAmWw
gjtg6gqsHkRPVGRHLiRIvScrgijxRx1zG5LfwqoUtW46g7RrhVERmuAOfK/xLxu9
jCEbX4MSv+ntyyWehf0fn3K50xJU4ew/633uYPUpXs2NVTRguHEC1ZQuoi8ao/gK
Tbv4yvC3LFAMAkmlIOqPn120AWVawFVnpoFB5zx+Zab7bfnHKNp4U/IHB5Wuik9V
cAKtzBIYKKwyVU7ewC5IDbOcWc9Ta+xen1c8NhOJ7+C5ZqI+pjae7H7o0BV+jrZs
6e9xFMxtt+CIWPEw8CVMEEccl4ll72lGfY8OQvRBY5niCAhJgnNb5mI2TS65k71c
xXcERgMD00faQSCxIGa2yChFtJDF7d1hzTiCCoOjsSQvOyhnSAORvQUTitZoAesm
FVJ4l2oIx0J6ykmQVOzgp5f/X6q4jSB+8/sVGdYHDBvW7to0nGiRapyWg7L6vuPq
8xUDDTeEA/tH02jvs9uuUbXhEbHUqZTK8EXGAjiNDpC8IgwxqfoUHCeOzUR2GRIo
qQyxDh4ASQQVqrlyRRMGxCdi5kvdAL0+KOQAJ9iYQk7JuRugPRv05ZQm5sh2Oqmx
Yf2VAvrwKrGsd49VUfyJCF0Aua6GdHZdZFAOEdfnj5QBx90hPrDiV66tFBSoLdMS
/XBMFPalpX8Hiy0b8iWdOF7ox+1UqiV+GmDKNZaFTVZgdf5GNokQkKh6MNPvQxRg
tYvxYkY55cFx0sAqoOHPHiTIwNZ/r9ulma4YeIyqCxpwyU0zeHCV6geq7OVbEPHI
zN4/mJgz51s+mSo01Z8/rq4v/W+4BorufFzk/MXDkVVfyeKcFhxYNIZz5uvy22VR
Ibtfh49qEFv5ftBLYo7Mw6yicggTn8Uugt/gcKUApsDWLh/vzn5WezE3T2xEFn9B
JynqZx9jwxCREuI35dNhaWos2OoXR3ayeMt1kJGCYSue1pzw+GfWh+9Cq9Q/4SBb
rNGT3X0RJfmTaaRCZQrECfRTNlqiXOJeQlEmsrUWuv99kPhb4vTzt+mV6rAS3r6K
lUIDKJW2h+2v5imN0UfYpKEF1lg1+3sIkIGVTipDY8Zuoi3UhMMFGiC7zRYtcTQE
OwOnbl0csiA2zmbbh5jsUPWM44aSEvfla3zT6TXYY4J/35yTBeAnlvQKd0N9V0Go
3jsnzZdoj1S6Bq0k+BJkjqlBi/JwYgphtw9AhUMV6P5MAF12NmgZ9NmxHwGPJhb3
O3+cu8kv/lE1sD+a4Wfj5H/BWVdODlow8G7DFGaZiAzG9k5jNOmJHvSI0sk5Ipe3
ePrCkOVzfMQJv2f7oRsscoPkrTsE1ykibDNbUksUmKsgx2lyfVdsrofMNNGfyiR2
jNYLdsqTytH97BDe/gOEivWKdKzNhrbq82P6rAWxiVIZFwmC1dKokuEwwGQE5uwA
v59pqFb7c9Q7sz+OcvSK2HNbatlCnSVIf3rVIzTsNX3bjBRsyT26wXnHPOdZEOY8
EmSW2sp63KpW6Gvv5hmisyxscXeBAUgHr9bcrEwGeIaLHGAFphCycwclHRQBBMlD
Z8ZZv/7369D7n8zFXzPRuSW4uqNUt72xwCUmwKwiC3Cun9MtxtyVzqGGEAPG0lod
AeixI42BZ4SpY8Ey9TkLfA7KnVvYYOCU3NJXSAa9YWJtlHJax+gZ/IbhLkzZ6+mg
QYOKvzog3+o0Jz1hwD0Bg2s68A5IaKzr6FvGkNf7Fsoda2JQs5fbVa21UmyyyqtW
JnlEDXuRSqHHkCsHXku4Z4No53huXyNThhNG5kBaibA+8TMVh2D2l8M0Y3MuI5d7
MrzaYTDPWHVUSiOQI9ig9tP8UI0kuZA/E03YK8H2a0dxhpklfbABhnItN5c5/vsy
nG201tUh/TQozZyX1M3n1yBXmk31Qe+O3W5eDpBnCQL1fmmPusuMSiAaftwKAo1D
o+Sbdna+NqiMbXGiu6fuwkIFmQFMwNcc0oYLziohLBpClJUSk2JYzzfltyOYOOUk
Y+4QGICsmVmyYhHsDDLmpm6rx1fL+tr/G1tARva9DGCrWQTLkSYFPtbCnrjvUuDm
MUB7DL0HUAjtBAQbJfjzy0uzbr+c67p5rI7xNxJk1RyYxO2X+1vESvBkLGzPSQ8n
GKzfD1UV0vP3GG1RW37/OuftMamh4d9tydWU7llPfl+a8yFAgfXQ8V7QQfZbHLP5
dCeNh1rRBW9imHvazw5qz/xWNfmNYtG6ieRAFTsxfInWBTtUvMzP9/AM/HrWBokc
4jwsJOv7FZovbMFR5UowaU7htx+WCphJBnmBArOlPuFgJFcWdKJY+Selp/OOSCB4
T1wmowTcJ2GL2PZ0Ph9GyOOugQf/A9gVcVFRwbxO3tx6wFE4q/JvhwzrxLiYcveQ
c5Tddrn4BCrM0oJzwor3CqMneP3kalEF5oqPJlGKraTab58Sbj3wPIGYnVwhK2q+
PzWrcw+pq7UUbG3XLo9wpwtqn0iyGuf5EBC3V+RXb0nVu/WoT8XoG1F8hcF47/I9
YQkg9i6fxj5hWjk4yU64WO6ScNiHYdUp8ibSxjGccwfKpyMsPGYgJOfLcEvKf5o1
nGgVnV6IWBoXu5V/ShKZMEiz9hkLJwzk6vpKnsZBlZV0qAmZyPhb3dHxPkRjUxwx
uQUF47aUq9XcmNz3vQszBx1SbLW+CPELDGylj6eyPpjSIELzSy78Qey6r255DXht
1au21m6PDTKLIdLccXjOWS+F19N0o2xqvS3j3VKNYYBihfN0Cdcz+UmW/VcW/5KQ
qF0s07Q0qtWvtuumcGfy9ATeQN2SCvD79FMImrhjorDl2p2zmCGDb0NXfguXwoPY
Dq9EuoyQsg2E0cPlfm9aWE7bggBX9szBWl5HY+myCX01tvu/Cq8ukt4tDsWbtBP9
GF0Uu8ioxGfSFIF+JZJ3/iRSi5DIm1dajYY7xwyKlOtjKhdkEveimXwby92qevih
ZDzFNL7qsVeNZ9i54AJnar6h3R8ri6MEDotDnhDyw5S9LXplf76d9thHWFldmKM+
pwsA008mtw+LYvdhcDABaTsFKKtzab8/VWzOdRcxOHTDEiMCvLem1vGp07jFyvIz
eWt/Ma3foPBzpySsHfzEAR7bfCLzWZwWt0h6ujUtGat9MtYz0aYdAfHDD/ti6q62
e7xXR8u3X0JqmRvCRx6o4TDek6QhwfB1CheQnHiLZB3y+UcUdrfCMWVAPo3pFABh
picAD0DBgTKQsq2FiG7LZyMO7jX18cQH7TmTyfJGZbQUPmA7PSkZO8Udr++0iNOj
PIwx0k8u417HmA4dfFnrBfec9YDa/LcSDoF+8P0B41lvAIByheG2Mu7eQOepfJTe
fSlsuWi5bNgZ4ju2Vgoqn0J/ALLcx41/YMs4+jZ7+UAhzJ4Fo9RFUmLa5l6JMZy6
xVXEU7CS8Xv5t9Hp/QStq/iACwv49qU2PVHR031H4WWcqP/uivNKIFw1W8HY9D8/
lvLiXe4FBsU4cRGgzRZXm7rRNWm7Xcuw31RvaFxDq/IhcZlQez3ly+3RwZVz2sxp
pXnIfoVDX1W7M94H4gg0BWxgjPP2ha2+x4kUMIsxy9h4lETSPvaORmqVZ/FagyCq
IzW03ZGokJ3jfQlp+xzp6RrumcEjSlnXy2WblwMfp1jU3ycidYYsJeFOYFkUZFwl
7sJqxSGYVI3cHwUy6BxMGDrZvO0uyPIqzG1MHAtU0gq+hx6T4LSvfykpkNyPmsTq
+Haefa+RTK73sfJr0kAX1NmccMa0dJEAc8n8oTOBWdQ3SRu5uzFoylxfl6rOXFuF
VTH+H9QRjOFoD0prk3pvHp27g0Yl64HeTF4OwXRUHdQtwp9zbf0efI+yf6KF/GXp
/lmrlp9+iOOKxFHCPZoNGU6E3sa/vPVCZvIYyi9OhgH9NvzWPk62KSDze7hZqTk3
8N5RIuuP6bYcNWBNfhC5uDg+IyyY0hJZVbHmvfNFa5xj6UYiwddLgCzk41DYA/pG
mum/vaOJiEx1VhBB757+yR6+82sAu7hNKDEWtQVQ84aA0eMhnM8zOyzCXhyf/t0Y
5FgUo6lBmgfBok034Fj6Gy4UjB0ZC/e3GE+bjY2K9l0v7hLm5BNtPcXHuAKTNXq2
yzuZxJ6VqJ4QBT5ekwZUsTFE/8B5LrwANBYq0SVRWJ3VjtluC23dZLjIqmRo5B+3
XCZ5Sg+fY/15DaJMer3iqjoaeBesaT25JFi5kRHlmLypPtk3mSJn6yYPOagA3HA7
x0djaCap9MK3mHQCTQtZ0t24eZdxC9Ob2JXmu01HQae6L8w3C4eV2ULJKulO72ZU
epX1yXJP2FVnVio3g+ABrD/cVk5UgwUU70TyA3dE2LDcss2TjwJc9loByElzdNsP
JVZA70AOy8js/goyEMnqQV2zGlQkWq2PUlv8BDOveuCdbwjJAkBTDkZydOSaR8EU
fUqRC3WTiZspGUzeMNm9/poKZGe1SoLpr4BPnQ4SCASXplqFum5zm/ThcmjUzEH/
WJuDhoFTIuvpFIUR6jcaVKIWGStKz8EWvoLnmfoYBVAvdo08cJ1EztBU0ztmXgY8
TEhECSG4wCfypL6MM8vbEodXM5QZCx5n9bHw/gES5H+HkM35fBvEmFwIflmbZ6xl
3NSKhiEZidJikNJkYnXYa5N8t6tr5oAIugOTgAgt76WLo0z9affZcwKDuYLLClqG
mzWbLduPDgmOQiKFXGAJFfFJ9RVEv0BYP6cHOOD08ShAHMbVIwBa9QfzWQE2Ik/I
z1yZkQeMFadxSMeZOav3i67QghtKT8cy5YAPaXSiibo75G+DgtjzsEjtX+yAIOGe
0Tghpt1y0/KPavVUsUbVU+g9Nnxr4LQlx5qkYQrggEoJNo33C8HtQaxBXvOD8tQi
wpnPGcAydum06dwcT8+vbfWIexAlj4cwHkJKX4Ziod1t9NfE9J3JFNY2PdRwuYJ8
T6NZ84W40mVMX/eM/YGSEgJWRQMtRVWazjYj5/Oh1vfZTsAz49+8vFdPcTMqKZxQ
PPz/OmbdkSa61L8XEDdsFrJaQEgYYco/o/lDClKuy8MHfelXTlxKIUPSSFv9VUth
aanzl7c106eUci7hAvvk+K8+mJSC/KI7q7glL90IBMfg8FljhGvJf+dURdQNz/Y/
AFez8aS0LWAZpqdqd1BMojhwELxUiUbIxIUOtl04pA27J7WMvEe/f2Y1YGsRWdGk
1I1B1oP2OWKgkTba06PSoUBhzX5rzZcGMFg3VPKnWU7500F/yr97y+O5I7+YRZsc
X6IwmRe5RqlRbD1oF0cQjycPmsR2CuyHACQLh9lr8/4CgqBx29gWYX/IhAsFpD9y
7scrX6BBUa7bfiBwB8KYtAS+hLpBukK31Gcekpqv83nN+cYCTGoRQtZgsNqHUqTL
Y9LpVSXNqZ5cujYAWshqlVYBEjZ7tNGowYohK07vlWCrMerQsoqGERN+bKGhJ5GO
pphaIPbDZacIDHy+nnk1vI3KhQmdv5Tne2bVb5zqw6XzKh34YxqkvgF7MzofZb+3
/4lLO7SNwoy+BFrUawu/xQKzshgzq3G9SMPpmsQPWpvT67PLhYreQ0z4ZQ21GP4h
E+sd7Doj+n/4y6XReTVW400D/CAzwSJHqZI1Cj7W56Mzw15Fjn21dOicPyK+QttY
lY/XB6iupnRj1sDzRBkHg4S5gvwsqzlmxM487RrSZEpxlHXrJj6PxgSJA9r0o4dG
ferHw8n+0tKh3WjL/8oZ8yUPO9lbCu2oz6M0I7H8j8kiMQL6ttxgPHidyCYhKg3H
kU9jpK2IIARLwOWf87KeEZX/w2HVLj8irws04ZDz+ECTAGWqs644kLBAI/XcOjGt
0JxmRK3Dorz9UOEbsTnXV1v/V9uY3JL8xqP75RJ1YS2OOP1DpdtyRfJ2qnTpAq/F
mOHDbZc4Uxyv7GRXHsxS1KvypbUU/dEukKkeqiNRglFIL8FNr8pWX5ceGvA9mMBw
8mb/VSvVNkWQKW0/jAFofUXd2cYI+AnAL/dGr1EieO8jtyXF9Fv8CdfpcEBDdFaB
yIIYeg+ZY9yqDe5OR6OQ0DGxqTDV32D2yuDXIU+Sx7dRxi5+PkQyHFxo/ecnOp+9
TOMi+GF01K0CpPzqUZ+wj/SoljfXLYwFqLGUm9NNLjzkOn5ES57mYDsSHPn1j6qk
AYsrJ9qBZzBdUXSWwX8Aqg0j2OJd9FgtGXLZSyJM0wyQiCj51JKaemqilemQJNy6
CW/m02s6p8UAu5uTRY0dgljddD4vBEe6+8pIZRiCEbcMDdnLCITgVb5Bvo8oQLLx
Jd0TJ8nZVeKvGqesiY7UU352xMZfD44Ibg1Z3tePVGxiE3gl8yCus898TLbhHpK3
cjnPCkk6JaubLfmIx42n9pB+uToPFCcB4oi5ydfbzyw7XdasVUYJQ6rQVAu3Xm8a
D+bm2MHWUaxpYRCiaLatjhg2M2as57DkpRFp8SnwRdLgV26fIoKx9RypCtMqEfcn
waSFK4I9gS9WkQDaSt7Qi2uoV2HV/WtbGMtcVW+/xHR0wEGlP+0XRsOPPChwphcE
6tSxfRsHQBF35CUsp8UUaFdKAzzRaHKYyalSjqnHV8HGlWM+a9LQuKB9ke6xFx2R
j8PQy1xTwwJWud3WgMkSyRWJcDxVXE00hVtjEqV9GZjTK5BlDc81QEX1U9KgesEQ
cvV7+BVO8Rp02wbSfqUYHNbrYwAd+KFDRgrhOwk8HxawRL8opBCTGhADj/D9UF9J
X7/jpVfeWrKOoMzFrWwWUrf00DY4fTQdVl6ipiYgYEoH4tb55LE6yh4Idgg0zDqu
C28849Eh5S1QDAooLikEg/ttn5Nqt4564E7cFbbzT7YIrq2JAbWVcq18DnGBTQjf
Thktw+VCmbrCtyoH7FnKRrLw+9cgzHZHtQ8ARTVLAo+YGzby8X4XGh5YJaUFJFCQ
lzFGKFdnyI/53z1NloSj342azVgEFJkprvZUXiB7mScR/bgW3DyxJkZ4AqwZ12D1
OInZ2EtpupGhF8UqHZ17vFaBqIhWPhTo95gnp5pmNDCTt5+V41BCoG5qea/733wN
7kNgCfkqo3vwXJNiIkduMwWJa6BYYcsxknt+A70oAbB92n0BBlkoerKz9gCXgXQW
13Djs2rCUNYoGrz4D6mSr8Zf/sXsd9oc1hCCrwpBHn0qN5kQ3ZXXwIGePcGGSXBa
8dQsKhQ/1QxOnhBw1aX4LrZy5OTAY7c6UvCmpAsQzQpjN/XA5PSsl3gASvdUW5/o
JCMJcYP3nikojbLKYmy1xtH77NXjaE3NjoEzUR0ywRirz9MYfm0fzANhEJ7D5vb8
h/eU/lCUznwevbchG61VklktYUj1sOoBjOIZq4b1U0jGOnicjAr7Ved6G3iAMvmS
nVVGJGAUrBwDL0uP8ubUfl++KWY4t0+yudTwRLgLiNWULJR6aw2shiJkbKcH68kt
gGUIehnosFhwgcjnGPjLuJFcOHbgEOliX6BnuBZih/NJBEFt7JMOSn39Ub4LQPUt
NXT6nFXCx35tW91KfDMgIkBZHkuERiFC/uaswQdmfM5XUS7bMUsFzLq4eftJm1T6
vfPHYMMaWKuEqvPkMS597y75ty4w5SFmkGYsmn6Fb8fvdXZPg5aPcIGW4NPZ6gZT
HwygU7vNX8AWWFK9ORHMcV2gNIm/wj6CaGULVSmmaflQkfV9ePClo2FrnAtrdhTr
ZrnAD7c/3z4Jyv8Lo6sUMQPauqP/S+MT/cQmZjh1MEru+ZSEpgzLdVZJFn5X1sCW
hgneSwf9kjcdvhjUd/LFDp2NE2BOd/4ryYoExUQN6vbytg00aQ1du7fIH/16oos/
kXUL4gRx2zz9R8ynxqoJaA+fx5q5/wV2vaQ+x+9M+u+7PjQsTbguLODYac4iVqc5
yUeRhPpUX9TXFDM6GmR3SpSe0o1jgFIXxpEW1yVwPOV2DlS66YcXt3UQ2ujonHbS
a4mjxS+Ms/anWAkfLCP5ZOjwfTo49CxBkeOrVcIE4Kr8a1Zlva1Rs1VSENVAyn6q
/++NGsPmSUPQnMJOHTv2iA6UcLJeyzpGA3xFcBJtyjy/0B8DCZ0QpY9Rn1QXDDwU
dpD88Au91XPm3eJ0eCTBT35AjJiKxu+LnOkW5B4ruRS6wSp9LvNTjZkV/F6uTSng
2Zv1EbCqSGBP8V1e1RfFXrtBxcyUouIuN1fGPq6RriIsS3P/akZkWC+OHGrZ4hkp
xsVLc7bHUqYrOsXCLwAnOxVEs80m9ga0N4Yy1MEag09ToLaGOI4twDTs2jS/ieoz
N5493EAkaNvzZQZ8GLpoyHpWOIT9im9KMCw8XL2Ekhgp+Hjw8qjFNUA0ulIv381r
USmwTY51Xm4tDE3iJuGZ2y5UxwtDfvO0ec8wpNXWoW2SbGXQlSQXazxhqHFRfu09
M85j9QTlmwh4JqbZ7O0N7fgLf41B0HQ5NI42e/ayVHmJEr1M5niG4C+JtiM/cq0N
juEhGGnBtLeoubHpCdNeOYN/31cE1BWaII5PFLh/XXpivnBBUVKGEB45CgiD8NpM
lRz2ofjNUI8ekMAprEmhqRFLIbo93WzGMO+JjE9qFbgpIMonXesG50OE33FyQGuU
fBpMnxjknx+PeaIAU12OwTBIQ4HIZR9AUlOZo0SOTsImrB3vwPJsLo77+O/NRVdS
ytkA57/1MyvrhmfVXahjzmeBdiKXKLH8vcdCmF/HOU/NFUt9AndS5m3rGjsGi98R
TeLRE4o6bz1s4qg5NYB7RY1EkLPBneIJToyXfASb3YupyOmN0uZCfK3PboPRks3x
3mZPCd0kzMb6X/MubZ6Sdgwe7fZrBhBsmgsSQAz4TKHea7mhqBTQVYQHScKduN5k
snStLIsDKyQVN/ib3GaVs+S7hktKyILr1eJpr/zoU94gcr6W6FMPK0m9+goyJkAn
cfruEnwptarXBUPnx2zuntp7ammzwwWcN75in9+Z9k5VXhjIvdvRGfR7bioH9Osi
6PGG/QFWf19fN+VQyqyuNzF+Ymrz7TCO1gJ6Bz+3XgWHpLq+TkyLtLlrQzWnt3wN
p3hyJMdZNySesXW0GfN5ackcUEQ5q7mXLnGp+xIqQn2IijzqKYnDLUijw7j9IBUv
sIR8ltzCITZG/fH9ESTXEHKy8Lh6TcJ6mx3K7BAJKaJHHMUsnbFinTnNMdzo0cvn
DLomrIY2H0QZORABCFO3LMLE5bsZojlrJG6qvPx+YC9AMi7cFe+gcXbyDQJ5DSfi
hLVwY4ELTCzUTICLr4pKJM0sD3F+bsY9v5b7aU/W8PW+KBT47jzw05g7cJKuphkD
5ZkzZa8IRDvUNEGr4BK1oF9VRbisBXkjkb6tmZVPvpOW8hWe29URKy+OXlOpA5Ak
T4RO/HMR0TC57CwIfo+zDKMrlwo5s2WHXVCJJISq7cLqTL+w4bYYjeOXKIigWdy+
lcwnQRcrdFc4wxAZM8mHboVvTitZmlObz3hZGua8RdJ/v737YRr/MJFhNdiF6aIq
PzJns9sVb4xo7UoMUSmUEWdD7E5rHZzWO/aDfbMGsjt7IJaBWbBpDi+8y5MZnvpO
2G/4JPJETgVJ4xknMnwDw8A/RYc7NgVovCdQKr1TKKL+agI8uLtgaCo+5Mj7UB8Q
N9kP80KBg7sfVrsfy1KzCzq+xHX5MDxlVSPNnGibWZJVWKBj0BIeeHUbKB/czxrD
OKMoaGRd5WZMBwJk+lEHCt14J5BM6LXZxu+JrAAaxgJBM9mZs190cpNTMq5J4Y95
DMWk6aM/w2HDHxhn6u/gfR6QAHwhM5MU2L56WEVzzQtrfnTOCMmRlFyVULH0Dn1P
x2YcLGMZy2mxSvO/SOazuW5akM8mOMO/32I+EOEYO2w8oAwscFrpLIQzGn1/Xk7b
qcgba9bXHVW/b3oBZVxZFFehRLQ8zHSpHNQWj6qXNWZLMbAyR6lXUQlzWGXLAxb5
HZHbGfN1AWEwU6zVrQv4JT6LBaTUoK2g8PtE7yQSE+ZMEFhSWCGWgMhBgQazkRh/
C2JOZAqt9tQCTACUUcgigAmcEJWhKrQIPS/Fv6c8Mp2gy8gwWArpmBtpT7ZorWxG
uLLxWK3OLtHq2HTDzeUf0zRmnL6qARa6pHC3EYtLvjsRH86WcVsCO+8zP+rx4/jd
NuG9dQUzCf/nqDl2/kng25VgsVmTlfntZ7HQZMeMiM4ecWHMgM4QuGi+1AzZHh9B
xs/gjEh+aaWhwkDQUAX3bAcGuNb0ZTuurBEFrIrus/25gRIjaKfHAtHJI23wZo+v
WOobq8YoID3OZ2WQfVv+FzCli8AXnWT+SoLL0V4QhpbP4Jao5TG04M4CHGT+XRYK
6z8XUynLNI6D+4c58HhYIATM9+2bjIHSjXnBaOxMTfyhFNsi466KqJv9h1iT2vcz
4V3BQ3jGGqciq9T6VeORvqXLmpbmY6fzrHlT3NbwyG8/KZgLDNBlhxsRhULabQHh
bG5D0Fj1Ft5CPln1KotEmkUQDhdjrlHOLq3GdaY8XafBlYrHpZsoWjeZIs3TaIUk
9AVNbfyKv9o2OSvxfV6dQWVsu8PQAJyBAFSnRm3cqlrcCI1j1UYc45aUbEBCbIK2
quP/PqQckeoNgVxkb2XOSp0tj4IH0CnNSqKleeWcj7jLeiOFLl2hXvslI8265nE5
B4tqf9zwjzTp2TdCaW+oKLC0Eiub1smhuyhf3ZySANbWYPcVqEdxnuE2sv1D/mmj
p2JA5bvwHlocmVFJPhGN19CONRTJC9YQJWwQ3GVRE5fEjg/3h0n0/aXtu1+uMY9w
uvT1Y5ItvkFnAJyQAx4EuUM+SLhnmlV0prNhXbBDE6m1wSpLLEwNw/D0dRvXp5M1
CUGwZnMIUF+x5TnKxV+p4qmlnFv/AVGQ53U0ancPciQ54Jo4fLh0eem2ifqinUqS
4R/IcztFSdazC2JjtXjPtLiUiSPAHtDAwGiiU0GRMwffnfME+HQnsvxSf3b40B72
DtdpJNcWiSeBxabgzACmpX7acLQ5JoV4cvd1wyBVT2tBEUJtVzNlhsWTUlVMlH6M
uoWdT4GS5+zrsyckYsq/tqBS/IO3HQZA/cY3KKyheWaPGgjqU7K32pL/EIWVttTL
K9Mcr6d/2SQ+waoGSRQJ0kzqDrpGnN09Lrx0be/uPoziyMiCTFmURyKWX1SPT4mt
a7BL8yiI2s0xesP6hpkuyQQS6lM0a8kDW+rrKrdrv5hY+ZclgbllKWsESqrz3RBq
ZiphAmWZwT92RSJorMWA/3RZXAD2PQiZAVoWH73PHVG0xkv8cleOW8wIuCuu4Ikf
2QTpPQUtmqcAe92Qc0Gu9SWjqF4pc5MTcFkGpnQohsvbrMxxr8wsKXcGSlLGmipy
Bj9zENOs3AFECYGrqQEIUowL+CQyIP/1y+O4VDECiMzZp3jGJRhoCBkENjP0luVg
XAvivZHR3Rv6r59wMnDcnQFBkOZf3sFzKHbXBd9IEiY/kHL0trQjcYLL330lvn65
r+q0L24HX8TnY5+/JxNHQUK/oHev6fRJl7Ac3tXWHdwDrr+V+aZ7A9Po4KK92CpY
6xCVmN8mK0za07XPGeAAiOpFSRIcTYgi+se1Ge6Vfyxpdy1qB1Uztc1akJ31s5z+
ldsJr3L1oRroiUfBTZ+BCcbLH8q1q1Mkpw0ImTKw8SgloUadLyLsCslZiCXf1Liy
r1Upfr1rZDhbxBQD7guLhcJaGbsl3p2VjZjTOEcame1vtMzDx/4Vaz465NRbQhoJ
ZSFatPmxOHN2dKAWu72qpxwBwPBtbqY0zWBGPPoJzBYUpQS1kscmWEoiSNiIyeCE
0tFGKLOl8iPbMvb4YeOXPisADxzagMlOgjY3g0VvounGZ9pTuerKzvCLALOfh/9t
NJhV72yqUY9d5J/ENRYOS1VLetZSz7FbYXxjP+ig625R9lbj6ap0gGZCZhq5TbvO
cZtGU1+ggpUqIpyaWa+rVcKXUwj31pZOuVQTXgCe7Db4QJUbX0pmcDmdRYEHL+RA
Zu7SZ2eaWNR8v7i+dsMn2xrCDG3lGOj+1zK62rBRYPcLSlIeWQGr9QEIJ5Q8DzVC
puJhAFY2pcHrFdNM4mUWz8EVF0tnsqqTUGjnHBcQzL5y5uvMiTCi7FfHwg82X9S+
P+n8UB/c5efK1Ztt7MW6A3YwM070aX1QSws7rL4vjHj8KPa4M8ZivqK11bykp7Io
7l2Q2c1rOFPRR9Sb44ZAOEDKaN9fhe653rh9vZbbR8wJaRNnTgYcTyeXoDPWP+Yc
ZshlKDPkY5zMpEzP/qfIdYSydmzEiTCy4gufD2pKVxRZqM1aPArbnw0yixlPGwJr
hrNySA2Z0/lI0brE0xlbKxr53e3BPHpNVEPoUDioDa7J2qhudpjU6KFAf/a6vJP2
7ixW+SPFPHvVBn2k+fPV9IXO4gWSXQAc9h4vQsbDZILO0P3hS74B6SbxdONQ7oLt
tBA4zYWof6mvM4W6wUx8/HRx1J1IklcXKDGd5fb5VOAoaVXnZhlTqXz8+j2x6jZo
n17NUT8GAJYDLHPGi6WFq8g4UNbrqkW6ysQ+XhxfHGXg9GmHUWv1tt6SR0xnQAwt
LUZ7FNFCcFnagIKT7q/hZBtpEwea4T2sk4/Ja+lzg6Lav0chwFkikk5li/fIi3sf
gno4M5nopBVwTJaLh7F3R9DwDjuUUhhuA3651Arx9dnUvmdViKEGvC16qeCIq52b
wHLFbl2EHsIw8+KTXuaq1DHkGi2v/2fnx5t4/3ezzb2JxvIkdo0eEfEBkXxhjPVF
6B0pnCkU6qvelWA5tSB8arKvq8pSglKzYBsy7wjqWIexkHNuKXotBaeujHUDIzxP
nfTZTV4gVmNHVXh94f8pZZ2ktMCzUejSmqCAyda2RwbsRX/LTxzUcuSsxC4H1Fx+
K5Zni3JYoJWJrB+nUyVmmj5eL/m0mqfX5Oc9zAIfjpBzHa5rQD4ZMBoMw9IGVtkt
MIPvU5+p8Z2s/SngYy4/0pHTFbY9VieE9vDwhILfC9ZlgNp41bgMQxF2pGHPH5ZU
nDVkX93MiVt4pPegA0ew9KFGpO7mrBz4juE/cPvWODuPc9j1VuUo3/MhwuuVYOLJ
fT3gITWNrkss0fBOo04sBD3KHQqNCnA28vpiQUaluVGUCH2r9QU8kxrfGUR1OwHh
4AOSwAW7YU72T6ICFpbaRA7/5ruU/b5z93o6iDKz8j3BQg1jYCnXCITykTO76+ww
uoMWTsjeaMmudOM8D97pGR+W77ZejinmUaKI2eYBkPqrt8SyzszpYpcJa39w57NH
MxYX6thB4KblRT76peSzDgqBoFXEf8OOFkeYfIiIjwPUdcMFF85+GRTRNjyyWA9I
E90hAh0RkeSVsfBhCnHgXoCyGJRuFUe/dZWRy3/CX2r736rw8QtTiOQfASLUPX86
gcWbi1sPPhDm2isZ+SgSsreXhYBfWLD8H9lyzCyhpJ1pnqEhsearRG4eDCNVNbPq
+Too9DHx4Kyb+xtBzILwWuAtC/VsegP9CMIao71p6xYEDAnKuxPEzfGOEg2ZrIFb
Gnxm1AfTiuxMnIi8Tr2/6IGSYF0+BQKuml2IkfxQhjf4C7WYIY/+XDzxTR+67eXN
BHnOEC7bsgT/x253usfNVBJeHhrUxSNRA74I6oHuIQthTnsYwuDQGAWnNstE+9MY
7bM2YHKYdaUYZSec5o6+2fIhQshlimfHQ8a1RNqDR4JGx1FTUspvXg9WwCXhm8RM
6bqHvkigtFpTJPq5wgXyNIlXYUUoW/SSR5l6QPlL87UWVF2isgtni9qLCFV92hYN
qri0Z5xiidr69qn/smSk7DK/klVM62v9pLa8HzNzHGyB8fLueimt61hwlbxW1UPO
nyTE3nRjyndeg6LpqK5edW6NwN2dDeGhxXqWJ4xE1TY/6IaCsSal57Ohh6jZ2QVo
lp6YpAVTxsVwuhns3/U5vX4G0zkakXA8vcn+UirK1ExBivbXlySypqdfbqt1yFbr
NogDlJddiSYGWU1roH20yGpQuyfPt9zN+J0ey7tClt4rD4iAjTg1oPpfjvJrLC1R
6+2OtC0Scsf671crt29uFyNz7Z4ZsVIXBnnvHOEZ947KdA2j8vq8BkBctidAG/a5
R9NN2cCSQZs+pQUfpkX3DU8lx0KFaQ8hpxZeX0w3IFW+RqMuBVcRgVb+sToAqogT
7QonJkA+hJCt7gLrBadB2w4z82IM2FIXhyaBnJ/hPMXb2uNgiYnMqgVuw/OzbY15
LXka8jHkMW0rjphgpkDbxY3nwInpv8GTE4CbeDGn+//XRRmckuFgfH3rMdN/bh9x
5pVaI948FXmey2uM6gieu1QURpBtzJt7zLqjKbHZqMWJZbkUA9TSSgpE6kd249Z2
fngcCaj58LDNrwDLbWWJ7IeJx7hxq8h9fPMZpznvNkS6HddVaHbAa6NymIjcE7U9
r4jQpucipooPusG/7u5JC+9KuJDeV7nwUU6LY56JkXENt2SUzfHF414tqMIwFKSI
VybzyQ8Smk5WrLv+sRPcfvFjL0VEZMWGDw9HevIVAlO8CNtCx6BMBNY2OiyqhGOl
oqEAA/teXxnBoEkEYIzM0EJMaPAUG8+EVGqBH1VxIZbwbS2OLWDGVaLcmUILypw4
ZOQnVOD5gOhBLWFAe5ittI8UAIO8NOOQeIV+gPIEUW/4uvgu4cUMJoypL0asJjW/
gA20fEM59lK1SyX3qd1Z0n/TqdpMtq7HDFkIpZBJogazj+ZNY8A83aYNZ4t6xqmc
dbhHaoSRt+nHSL5q9XqlbsdBSBRwLRJleemwS7+7uJTpyZXsHrh1B8l7tXvqTnsZ
7bTYzc77J0dJLvRuN8o/io4t6U5l7eGx3ftVlP4ZIztAnqF9mhk4HsTUUvGmd4zK
q8iKwCPVJu0FGhAGFdCGIwqglMjmGD8ht+7Mf5KKd5Ne/9WGgWYmMhyreN/9gymN
AQf7yi9TxIMqwRZ278LAXoFt4OoeM+aahudzmeDKCCmKntgsMzIG7NMjU8KS5VSU
II0Sllt44T6McXvx5SKRXddO+tJdtJ+Fwa86zFIUnMyQkmxFt6hbdA7rZ3DxyzVI
CAIv44/gWgkWa/1O1E/tyER7hKpiu5T62mOvZNaFIw5tJc1Sq0Qs8sboaLaBKAuJ
daSSqAeKtyd2XV6rPKBbHSohR6jE5mMtWqF095/aYNhDg/XnNRditWt2Kh7ihaUm
8SXldlFmq76F2DbWbuTxcW7get0EyQ7at7iJOfLWTXOZmE6UR/Dwa2ZKBBCb9AQ+
SbyUfjPrIGBF0uXNdrCxRl7ZMs0xJmJp1krD1q35Jxr3YI5zdAUJ5Kc+/At/Gw5b
WzPz2ZeQC22fSR8WJ+6IyXPQTcsI/zlendL0l+nd1N5QmCKjecco63fZtAK0RRHp
JqrwtHq5ymRr8EEF/HzPlRpiCyWUhOxu2DT6aXkitByV7zeFPrVp62fya/+DVgff
SE9fyCIs2CJFXZ3O5j/O1CY2QebgNWTuTZwNZs0gws2imqxX4QZcp73DEh7fX6ov
dhrOTooG9aRLy6miu8ullgUc1EGehhV5t2RSpmSgs5ZgzGE/kqy1wxAUwGbN/FkG
aO5C3vOSzKUzladNtOUs+QBp/Gfou2yA3B+pGGER1S9+IH+JB0GiPNE4CfYzDqXX
1XLNEUzuBJbEFSqgfneZftWCwAXr4B9HRQ01VEFrc9mTFYJoRbelES6K2zFw6sVQ
BmL8hJKkOrIWkABlkpAKw381kWc545lBIrn8pnJA8Wq95cCuD2OK1I7JoXkoTTXy
8xHDn6VqLElMQ2xd2/83spn6+k4a5sVHb17tF6x08qFidK27LZKNVs/MY0VgcNsi
LJjvSAai+A5WSnh8IKvWBn8O2RG5IvDCaZYWszWwq6IZTTkRLgROsQGTBZJN6zW4
fGnzvrVbspNgYCoLE90j9KFFb1Xtm/sowEFLR0SUqbOiezmoQ8w/3StGEgc8r5Tj
IbbTlzyItc6AqW23Ec0tj0f38WuX4NH0oTvlK8hem5J0PpioM4zO945X3MgYQl9l
mryWuPThqFSsvekQ4s/8QNHoXrmNCLkLvlPxrL0aCeVl8Ppuf2Mn2OFoIyD0nXwH
iibACbn+NpbHsp054gmXo29R04sGJMFi5+mHzgX5B0kTIps5QqhDR0+aqzVXVLHh
pHkaV/TmKbEFFYtXsCw7FQLAk6Ng4tPZTuX/F9Knm0wacRp/bsVq7WfZGa3JzJ4S
wusNUbMzdvIjVEl71ZLSv3S5+7DGdyYIzkLCQx/meeGPFIwvvf3s9IZNZ1SUdRkC
HAF3TuIOcIS2GiuMHNixlVpNJXs/dI7kcpKAm5CpLNsLz/wntUwXm6EFPu6Bhu24
V2VSqtX7yUCb4nQGDm9ZvrqiXbondB7Zjs3a+BCrCAj4fzr1EsUoC5KNNp+B2TQi
owEqWMKoRNNOIQ4FQoYSsWVL7daUl+658iXQoiVaX4nj3oe84izKk1lBccxcqoqh
7FdRRypaSIGAjLu1Ppbi4H9G5839EokrO6rLtzt36diH4aIiMPZY+DRIkfXE9D3W
SOS8g3z1iUEgJb9E7pORfH3OU6yh4CiEGcJ0DUZaDXYjGwIwSyeO7PEKny8vsVFF
/9Ooa4ooREZbNrUjbwY37Pn80BZ4JUjIHaejRLDPJjFJyCgYgj3cvxkfidzRYNl+
RmZdKzxht4nJm9hmRT2F29uhpIGaQQLPewDNr6HVL5mH2v8e8+L99h62qDyJBgTi
BVFn86ZpdvP3qd1fdKmZioO2E2pwGI7hT5odTfiIy3+P82oHHcLwn1p/sRuOm7yk
iZtKpFgxxE/lB24d/84/UoAO2pXM+UtwraYZrOX+HfuDPhFNkFB23oq8spPIXhH+
PRhmouBXi3o0lh4g3TFlVE0XDUEQLdaCelorUmak74adG/97/aKHJPlsFQyAL/u+
vtD3KBFDTe4+QWYkFsC8bstdG82ojIxuaxVh+lTzVpEcqBKeSPNMHoCURhLbeSKH
ScfBYwG0Tk+2+0f5yYP7nU6rwpR/0AW4J6Q5tmEt4oB7NUoCQdnGOrGWeEqRhFGO
zBPhw0smzX3vlbVV44N41Wx2XfQCdDeiwvcGja30u0xJBQLx8+qzmmthv+DYCQ5g
pW0Hn/cH+fW0K3Vvw473NWqSru7xkiaNLrO4Aon70SOpxdmRWCLA/f0SpxyCOrLF
T/NkfEEKsruUxoMfl+Cm/IticL3JCkhHSgUMjRcFzP9iSLu7q4c7168ToFiD7nGQ
OX2rqPsoOlMNbfvACNvX82FWfQ1WXeLbTU87lGhzX6UBGNrKOWqFKHULv/YuYFzo
rkSYlgP8np2jMVHstQlR5YESyrQWaM3TrR2Gp6eikqOmJGGYH0aaFBs0AOZmgm4L
U7j3bCEo647r14U1csoqvlSm2SY0qSp/uCOGQlLjl1y7gXZUNiSfVKerm/kDl11t
NmALeUCQnD38d7gVxVX4biiSy2D79rFqUYkO0n/roNzTQYCkcartF1ZcjgeJ4HUx
mSGyvDJzt+yOTn4f1huO+boY0QGWvdXjtmvEhb4Y/fSSQ/FVlGkpm6GzHUEIpPHm
BbhEeSsgI0CO91aqypKqt5DAnstvoQ7xc39IY8AmVx71CQlGbvpu0lLF7tIwpE0L
jqufr9zCIfgMZmeD4TcxTNe1vKUNQKL3b5Oou03u+7PgLtBFZA2qvznGfW8K3aGs
UWxzMiFvgxw0+7KqZXb4uda3GXGrO2Jr4wqmvewEqq0WP/OJmpnYBmSJkk2qPHcc
0KVbq+6A5HLU3esRsUCQe0E23z1UL5GQG4rl6NW/ieFbL0Da7CTzWxhxVxCfDIcu
FYYhtlFr4f9Jx/BW5gW6WdkfRLNbZYa5BAOhGy08KlS9ZlyROTypG1O/1kaoC61G
kHL7Ext98eKvUd/F2fJDpCAg6AtOZV+Hj7bt3VOC17DD05gJSsYApFBwNCIsh+hX
fifpKfJWNu97EL9u8rE6+9ID1Avlv+RrYW0/ncgQbKeYvc+G7LmTlG2qyGr6M/bB
7KDQ8o4KiHOXaqCa/tZwjEz1flZbKRXGNUAW9pvdiZ7ST4duY/uH/GDHOTPiBrNY
DJKk2F8eEIg3WkAEvT+Ub8/s0IbbTxVjKm/5extfPS3sjaIXe0ywmGImA1PwQ83g
/AP16XqKVXI1KNB+0hplG44EQPNPkPaQTzfsJxP+T23mQslY/VNnekqKbbJVuo+f
ZZXra+bOvt8PyYrtjWAsIM7M95mJVU8DbfWzBzds/wCV5JTdhASOFdGIutS5xX8B
zzlji3m2ol38ahL2u5Fqol1wE/RsRzwH/PKwzuSKy0/gKPEp0wkAuff7ul01J1Yt
FK5uz3+bcpAaaNLJpUx6ea+Dg7pmQKA79xMP7/08f0T/H+xs7QelyUqWLJz+DdkQ
9iAK1JbVGQ1xnVj7QNgwzgc7X0RnsQ/ZEh6tblHPu7ZhcIsJoEMdu9FQh0TqGH3f
98biLhaSwff+z5TaKFxErwW7uSJBT6mXgjAElwQmI7LmpAojwIwBkNa5nbC3bKJM
CaoA9oeCfDBKBGOOzOencvDEU5jyUIqzseeNi3cXRFuPdMkeyKBggwTJVvbOhk8/
ErsOI9R/WyUWbh4p0V9bZpUf0Kq+Gyi2an3q4Kxaf56eREtnpf013e9lYLt9wN5M
ML6HbPOYARbf6OZTtTOSHZ+0D1QJIlJYsKn2adwmNU/3O0VvIy1y5M2NZLkK8Wuz
acV8SSQ2LK80rzWUCmmHxSzPzWRFLM2B4FI4dznn4BXFkP9jjSQpnfwpJHAaMQM1
rnIz73EkQ93TPHVhaeMPNoyAmIV8lPzABWT5oit+hbK1LChWdoEP8rstZLhAT2gS
RTjRxcRww349/FfTfQBoGrirRZL2E9CQib4zG2NrA4IUsfCduIDFQ344D9Jbt1sd
g3582CIxuroFfiej15ord3aQ4NnSDWs6HS1RZci+14S5kqn1d0+U/EujbX1SyWBa
rYrYW3p+IpYIxIp+Kmp5Yo4gCF3FkAvSgv6ag7Ky4LmlCWG/LjrMxLMl+pgI7rAX
JLTyc8Ff8Zg/q3mUs5lt4l9ubapia+CDLFNZK+yD035vbK85jH6WEmQ1aJUO074C
V30yqpvfEemkXbOb4ZaLV73l/jWHLuZtcB7RPHoFGqSqDTwhxlbJXoT0B6nebGeg
m8pm8EzaRqMzu2/9q9buLHmqlW38SKCnaA6+YsQuzO8t4kcBSqs/CmAhCdw3kOvW
MFchkLMav9qeR91KlLQk4EMBalpzGLYGtZFtbfBB5M/sYb60bGS6J2I5yyaSl6zK
gpfJbub8li55UI+I9Y9DTkB8MISOG1pRwatFaB/iUOd5WDJoAarlmftsW/HlsqVg
AGgbZ9tk8g6Bpw27ukrOanA2f5H9ITb/MvGsUi3XQslxruSp+gtXuynM6LlSjJB2
crONunp46bLuYrjBTV5Bc1ypOtg0Qc+KpbPBVHG/4x0q+U8KbXAgYHmmrrdDGKxJ
yrr+V+fhiKBhngWX3ygQYhAVkI+jM9WAo4SjWNCicQQnFAcyzA96VwBCV06Qq+hi
SqjJW2Kjk6uJJX+CDzzORrInI5mIESsxPBkzNaH8X8ml3yM7+OOEONmtpsVrIB+9
qclRChwwZTlyhBvvQtm2cVcFApanRfDVFm3a4za8ST88gz7fwtlMEwQCuFBwGe/w
R137f/ulB6IEcC/isfpeIJq5eGVg9wLYUKNW59VzQNu1qKtS1VxzdUGMEOcKZEeK
rjYl59jrGzydFHTiSWPUc9Uc/VNxAGBotfwB4ovuRdUQsVMqxu8brdaYb4sYjUiX
EBfne91RwB/VYfy98BHBhrmm74DTYbFFpthMU9Pj/JH4ILgw22PpeVfAK08L8c1L
xRVvTrclOzyRSnplOTltve3S0AZiqGN7pVRjN9mOFtXdQLEhE1EMustPoPmuAk6w
Mj/wVOZLGSbz9DkTYRqHazlhSnFGig5Br63kbRFdCM8ZRHix4wz5l7+SvtP15bBn
B7P1nlJQQEv+L6J0AP9u04osv9I1e06IY4ndzNVV/4mYsUjk5xabt8vXLpyJhtk/
Z4hJfdvWfQVMwTbGhh1dlOt32MLZTcTOw1ge6GhGVYIKwOV4nF3BL4IfvMlA2EwG
uVonpW0SE2vqwC/7K56a4kDuIGwO9sx+TsjQ2KmbLcwcMvvg7RQn43PWOR0C9m+a
vtyP2gmt69QX18rmuQ1p4KPXflD5ElWSAMuZtOnrXR9Cfuvdh/C+Fs5BFybcbVkM
+5kDiAQ8e1tTfmzBa7C4CFjYoW3L8AtTztUujuWIwHUmUqMvleLY08J888LC7lcq
8Ps5srH1gQ4jeXzE2clEz/8uBvEfZidLPbw0WwFlOdRcrtoCi6mU5IJDZFvYeC29
90mK5va5wTq4NdCYbGturu1+1alicmW1WxPURkZXggt/oCEKONOuh+Q7q0NKUz3s
RlmtGbbQ8PMk7m+KqGz0T+Ms1xoklHyHVGi1AmnkDVKiOCWIppZ+D4hb/Nht+8tH
5n1t3N7DwXxDHMg3B+/zI3N7T6DVrWmPHM/tcvOb2BRcnSvGnzIzX0/Ks/xJWjON
e8QitaePua6ujgEoBQFk70SNowcEARvY8hG9PEj4ryiDU7pIH3P7ZYLeQ3DYrC20
KoadYTMd25CA7m0vjbuYjSPHmgkXhe7RB085inBxMCNKuvCpnUVe+AodxIQ7hzC2
LZ2gTGj86bj1PYePpXoa522RUBFE7HDj/+8KoTirZ82GRibvYphVVJro6L4aCaDR
wdgAHktoBxCN25DAZESXCKiX3O/Rf0CmOa1ZL5XdSIt9ZudduWZ+X5tXsmUJz+iS
izkJnuOK2e3QU8/BFqhCR8asXXpY2Li/5Haltc7Ze8XZtrw1w2gge5beThzaWEQc
erEDjL0O9XR2NOZxpnadjoCaskiKBn9tWEBPqTd94qoEEt5TNofqsmQMbgpBdYEb
sCuP7hzmR8hWObz31i0wnRhCjf2DnrmdSKiKxAVU0uzcRyNop6u0QUznc4+Xbs8i
FjvWYDEi5h9f+zXY7jp72tS7b7kBW9mZC/JAZeU+lrq52yAdRaJmm1i7tPxoVqu0
1xuj7gNvBi82N31HsANXHSCsdQ4qccfXLu12pqGM+j3r9qh3Zt1H6tHxDAEqqNC8
UmzG4qJZNibUh/L2Xvge+W9+Hb+dM/IXT+8dlE+w/M5bCNZu9adx2Kto/jCya5r/
r4OaCi5n8vziwZGYXMmfrmOWwGucK7bU+VVdtK8zwWii01k0yYtMMtUtQ1EWcqrO
9OlTTM8iIGGioQVjx2CnH+2AOed49uamGsBgEoVpNFPdRSiG61xLKEhm7MwP25SR
GBug6qgSl75Fs3KPhBsQXGD//UJPpZCdXdZkWGP5tirDy4IyUTbLSpjQwHK6sHYQ
ARTiY8NOzZI31RSoiXYwq3ST6SQzlhzgrwxrLUa2r8feyNBDGI5vByVHpbs0g+Qp
yxGXFzjRNt46hvHY50NU487JQ7LtO0jOJx3CVzDPlLFEx2Qb5KDnvfS5/xGynX/2
6sqRmqxqSvxoxUdkf9I0rOePyibL1V8VY5Eaz90w5ygBf+boBYeU+Y51OQenydYN
YxBXLCYqm2YRX8nIDjepF2pzQ7V4DZURiNg5AAGig4KmxCXN0WjFoQ5byVF7ypKo
G0KXCggrPe9Mg3Q83QOyl1ivjHSdJ8+hla9MZOVgs27VnBxxrLIVrOMVYOif43I3
ukJhBPD5PQsIVbAktiiQ71noxzOKYX7tiK6HVLEht7K0LWvlLXz1S1glHnQFMyhs
WT0w7+uZ1sidDZ2BHZOuy14pWbVv4iXtVyVfNK0tQ5SEvZEKbe0oG+fEM/Exdzf7
6uYXFC4Q321XnVEuZc76ySvC7p5p1qk38BGeppGJ0PbztiAEjRTPSG/4fptQyHFq
1IUNVOGo9Mi1y4oY4X64UW73gfEdeUvtHcx+DfmjCjS5I+lj66RH7n+NyctDlAro
fskYFYRtL5f+Ylu0torYM5qdrOM0nsjHJiaj2Dg/6yoQnTM9pmBt5Lb5pJ2OWUYv
sGK5eytcaV7PkLSpdEPgN+JF6SQ1/xxuA/AZM1Y0qf/Jo15pdcGLgDYCEHi01zi8
ylERoPfOgi6ThTooNN2+9zqR7+ZhzIqpjaXJ9Soer1BgYEL3Kc4vP2T5tz2X+YvW
iyaLtouGO9e9Dq8Zeavvyyrrn+WtfuTSRKoggw6O34fHBB0zO7kFvlAriJvPM2dD
8FW2XWwseLAV3N67s4fDJ0gNMP3UFjHcDxJ3BPwOZzYp2hA9QUzABSrQqzHsODs6
5EQPVOjXVHTojUq9pyc7g4MjXXJ83mPkL31IsYoSXUzKR7LzQXPQPTixbTDvMU3+
C43LFdVSnbIMwnAKZscmgN5m6HKFOERg104+WC7DADJubk5d8hRljKVAVTiX9T6A
IAjFt73ShekxW4kt12JXvD2KdfLGjNiWmINXCx/eGypo1WXwTDZxrP5+NqeczuXh
k86lAQRr0ZtFdXfhW+4BJtevNsTeUyVuR9mm5GZXpOly08zJzVRj5wbSaJHvHsz6
0fJGqda8QkdDhYEE8/YAcrK0n4VB/+kMFzju7UlvraPDBKgWDM2esy284hOh9Eqg
pTkQi5NxqG+K9vZ7YcXhD4NMQxpGH+j8NLFyHxAOile2ubg/oCi05QvR8XodbHPA
BotSVmJCc0lXZ1XCLk1Q/Wz75qHROtsgLwvujk6+0lVbfKsmczYExaWB0L5K/SEG
8l4JE1Q6wsS+/PaMT0Z78+33H2r9xco4u4sCtEsuSCBkfvtz80YM/OJLppEfm7hb
n3nKIkEqBy4IEUBx3BgiKAKL/0tLO8z9qM9XMl+leMi/n5xdCJ7VAnp4FW7DShPY
fmzjT/paXodppZzwdNjoEtDfsmagctOiPzlPSznVBOBcvsPT7GAJwZb8gZxFnu42
zPBgSPMjHVRKUZ7dkThztOe/c3mj4dNUAx9IttDPZFXI2Hc8s1I5Zsq94zABaSFG
8ODSdnetHQbTBjnna14Fw7dOMEAJ6vALOquxbAK6caftXM5M37FtLgonOtUUrVqo
2I3HJL7jzgP7IF2fuPaehc16RNjUb4I8nQhLfGpMLjpqnCQP8Ht/5yQRgNk3EVZa
At4uRov0K3cty1WDTy7vVr8qkc1ovPqpHQ3s7A+1FLFSMiDERW6znKRg3ZQepoCK
woib5PHxIx3NHomW1LTl8d4qEkGy3PXKcZyh2dHmli8HyKvrgCG0sdUxr/l2d5Ei
qJh3bycWE/7Q8BphEg+OCHlJLxk1gjtf21EH7eo89uWGtJdPfWJ/pSdvEmwpEJXd
6Ct408QdZ6tjk/B8LrmSQF1Oj7RxS+mHh6QaUYI3gKwDeQ9SHu9321X9Iw7fsF2h
n/3mGFK9xG5CD+9Qv468kov7Q/ftld4xDQwl5kgnl16kfs+TsPXTSq6//2rIxb0E
mf77QZ9dgmBozBmUccs0jNOimzfMU0sI08e0H56Re0umGGIXMO244tVlI8CrDEGz
w1YQ3BogY+gw/IdJMNW1MDmKGp/YSbFZwkO39fcQfcUTPFSzS7qDh4ZZHgX2hboy
/CnYCRVjeFdnvA8V7vPHf2LEMLQQvzI06032FxGKe/Xn34jqINENfXEUkpwI/WlZ
x5JW3NAW1yS7jmtGDqgkSU2z39WQ/9vS3kVwG/S8eCjnoDq868hfsGYH3HXl1g2k
lVkfyhB6Btly1pIp2S//7D3skV4XQelvJZl3ZZbyatquZ0HACs5u7iMNepQWRqe4
sK9DADeZ1i9ZfpOrbfW53o+kzyfGgnhJDZh/u4Vj118V0Gs4utBsvwVgUIPp11QM
Az9CeHNQKEhTUbiiYDlTUxIDT8NBUdjStHRqjzFykLQfrzyXM5cZ7Pr8U+uVU/c1
P3WDlCyA8GXRSakgvC3PBNPu+ii43ExkgMD+gnAKxm+UyBIdlrFtC7I1Okd1gcPR
P4Hy/BFOrXuxmyD9Sop6W7DcJUNkseViBGY67TCuEB0U1wBN2m02cWahT6fPwLBF
xk27yzwj1auHWVztDq1lpdVcG6v9Drsgy727f0lZufmZlxi4qRDs3NBEH2zbK+Vf
clFFJmi4m/u5T4PIhzAf1aj9bEJtOX/m9E37crOGoLDsArX+D1RS+qcweo9+E5Rt
enNVUKO8MGFyVONORYFUImJ2f5XwXdnXhVUYtFK4NVcXHeGSS0rSSC8IvJVFmwNp
xv2gS1ll6k1DLI8GflaAt0hqiVjDZEvTLoq7SBWk+spVP9cwt3fwvCMvCRc5RzaD
dbAejb9wQzNKFjeMS17R2XUNP+FRqhUHGR8DAvHn2dRfa0i8v6lu8w+Q1lFpgXxM
0PJ6uCOBBRS+Y2GWe8XDVdWBr1tOiT3l710E/TdGThjXen4wkc5DNThbWiVS3ap3
XssuUTOfV3AHHyin2bulJFeG2x6M+MVSqxcsW6uzr4lF8xs+Q1yuxLhI4hNmXIB1
jSjbaqurQgzxV6qlkNj/1SbLmnRB+/tagwLMXnV3QfhB0D5CUK4KTHsvvzSh6Uol
iD0TEVvRY8bWkx/swAV0Tgs+Iqx1mLQeTAdWayD2RNjDq00iO0B0IYbDNCd7Xi9/
0hQg82c+bFMr/r81cPvuG32otBa3Mlcbi1FmB62NAJrTLdjM5FJeicv7zYBSYfsr
fbsjmLbxDyL1WFrH46t6Klyn2Wl/Kr0mD5OaoQcvOtTAIB3mgec7VjOjnYwMdZB1
+KHjzYGjqXw+wNEPTDAQmiwf5ia5L4JLHahTRHxj0TChXBYOHe4LplEM2grjlt0w
3ljhiiezCeHjDGzvd4mS6HFeMuHwZFAe6MzZl18zaEUUDGq6JEqlhvhB1xH1Bv/+
3v+ai5gaG0HJQHvKZ0wxLkOvps5h+yF6c+jvaR6utf12qbLLMZGBpK0lt0EMdaM2
Je/jVZGYXPIYTZwcJtBMUKhbIDdMBXitEaX4Zc+CN2t8HGZaZi1GNV06c9llwrLt
UVXrYwA/p/ljUNIEAM6qusnatk4ITCnq6wJSMPFE3cdvC3LvSmaOEj4il0lGZy/g
T5a8+rNnLHUJupIdL6zEBCXSOCEIl48YJTHLMiO8u/uCQwrqDreael1TB87U6bLN
/XfL7HhLABPC7KONh6Js86s2x+Gn7LjHnKFN3z3iUJMgB9oJ/MDLaVj/8TAchGUE
Lc3xzNFxgjkVEeEc7yI6fKPhFeNMxLqzquMhov9eZRIkyVm8AYZgPBmxIzoJKf8b
W+dHsAbP4/3k0gCBgYiXPKuXOsOFvocCmVleulQ6tBCJnNpVTrisYEIs0quKlzex
dk53fnGAJA1R0l1UFk564tHa4q/6k3IBIT1v5kWIPnHLf7xTKUPIk5adA0E+ObOn
mcqSPI3d7nPUENq8ag64BdS9SXvwD19V+0Eo/U8u+PE2TiypiTuBNfKMGB7Q9OKQ
WxNpJo6ezEBh8bQEC2kPtUIOBScp8f+pcIumD6l3+n7mNnH1QcqXIh3fYJn7D9Wo
zVHHyQ+aq1ZEL+HYe4LOQdBgb2fuIcavkfWlfhjP+N6kNtmdtML5X13298BAPcO4
walOcCp5iTRU7mBjihULApxC4pDQk+zPuRSSKSZhxWtK16ZOrZZIOEiOmgVl5jNQ
oe0GT9nqifFAHA16vV4cibejbMIenB9idR0UfMf5m6fFrJeAMsPh1LJbjzxJoGXW
h7GKbdUb4edo7tb2OADPVoghtuTaIRuS0brW9SGHY8xQ+cM++y0PhaD7wnj7Yb60
4m04D2nZL3BzeLooFojB2BDX6wi/rwtoRoTEzI1ihG2EvVp1i1NZ/CMibw2JFWH/
XjD+vNtthd4+Qs7a62t5E6IbOnv/DNaV/1qf6DS+nhFWAYpxkmbwmDdbJHfT8U2g
bNOKsNtCmriQRAz+VGcrEVntckUhSHlSAOC9twcYPV8cE3E1pUBPlNZZyJkhdryS
Hg9bO647JaIgIuBiGEJSm57ehxEt78yVWhj5xFNduieNvuPBMLU9KX8ErZenWgvw
7GCc/OlxA/EH5KU+bBw1tEyzUPS0ErjXnkhax8jqzlKin2+AhOx5mHn1xHHorIvu
rmBaJJtr4P8vQhd3oMzv366Flhgce1okOLFe8eBL+7PgP0zCzvajraWX8FA0BROn
A+9gaK6jDtayU3jiTVwC5ctkfPOHFrqWRzQ2qDc+mHek7XtgE6bYWvWqWAma6m8S
xud5I4yo15bWDNZ1x6R4YnwASC6YMfrP+POyobsC6vZZz6B2Zm0g9Zd58sWDi9u3
FGNbqENU623EfLRgpVuHrncLNaqscz8Q7pYkUsXivxnYl0l0KlhQbaeQ3bdt3kOu
JyjqoMs+NwaDyZWp6AQ8wvav1CfLjlRRoZwBkVyiu495xzwTPJRDXeiKBQGe+UAR
d5UEuAK/wXpfG/dcNlXiIcusJk44gzwPPOkGhQ9hj6fVZw/Sj2zpyCp1J156f6HJ
uBMsLskEJaXAo5zusiaX689UDk7oJxkhvWioE+Na56IjJpLNuzw8QGBZ9tz+jcLr
qPJEqLVRqVqQFB2VsJAfKA6uBEMpu+gZ4BrusviUyBo8YGDXRrk5PXswPe9EwMXI
cLIhWo903xzgN0iRzFi9H9BptgcKJeU33Mj0GOPuy4IIU9N1wZy30ImEvFK+Sqmv
ZFY3YjcZEoyc8LlH3RPWjaji+wcV5v/NzUly3h1Jk+B325ebbGNbCLbRJVppUx3H
GGaGWrK287j/C4BKSTCFia9/aJuNeuxmxCdH5XhPTAbkV8OFMHSapPOyo/S9GoXw
u3gv/2B+c9FitwqDCk20Gw+WoMoanQkAyf6q+NfuMGKpRi9m8Ky/CSt5aVYry2ti
PpEqMEG9WsWEhbvorcd8yOqjgAnSY2CoEKLUIVUUvUSksdAvk3narOZj/wqPnoRU
41vYgIiW4aDzTJW3Wng1J0U4/lzA8EBBP8ucVrf5so3tkt1YV2LX2AnVzOSfpxhF
9dJBHj51Rzg3QXPSEvuRuGUod27Owb1rQxbI6UGHTpOfo3QMbrsRWUGzPLK4Cu2T
IpCS6H5GSB9eWEMDVbAIbC2KiaLpzofEN3OIiT9O67qjHtTF/b/KxAF2qSNZCdeD
Rolnr9Nrfip/9iEkWSilP+LJtrzvmKGG9ZWy1EFLldHSqQQTL7zGLhz9DBmbckkX
cGlILG5Jo23OoA14C7mgUEpE+iY0wd/BWn4NGsgPnZBcHUV+DLBoAST2tnqSbqge
h/WWV0aqadgb7EOeN3SjnwMGfSzpcQ6gYS29DCF2IeeL9CEyny45cMUSj3kNqi59
kvyf9rpTIPERQ+Q2Ot3KMkdnW5ERh2vUqgtkVrYK/pXctcW0gx3tQ7iDffhj1/E3
2lieyP5kbFufbBUy2A1PviRW+rgqWcwW9WAFD2ZOksA9PccNAXJS7hxADy4WhkQJ
6TSa0Ypkkdt2V3w+0zmyBOFM51XqCjZBkefrXMlQNyRDS1Fg9iqPHYUUBZwmTmEh
EvzjHGR7OM+3Uvu8tgtLsE7ULaFCoq1tQGspLCoIWP/p6FKGPpTIVajNEccugS8w
rqQVN8tny0MaHpAgzhbOZETfoR47oylzuTMP64mzouBUl2kDxnJLgqcbvAC/58XP
vh8OYWzY45FkD39A5CrMEXG9DUBiK/H/iPA1wLmF68aypNPAFq70PomcrX7yIsrN
VqkUhjMJ/Xy1GXRc5HLos9qrh1hrs3YdErNyltGEQgMxiseJws3Ztj6f46MV9svB
6O3Kj13J58t3O6r6N41zTiNYN9r8KQLpBF7KCdRqxHpXucJNInOB+9aIumAuzqYF
E9D1oSiAmY6HOMGFbvd910BzzHbftzcxYmg4FOzq+wWDVBvXg7SU5dTRdSF8/8gK
ObNesj3VNEvmdm13dhdiIQkTyX7AjC1aLVmLeNpqiyCiJBoslct1d+0waJLdAsUu
yHSPEcFcdopawAcE9VUOuLxe48VQjyBJi8I+2B8EVLpr4hlbd1kqIsc5AjI0oja7
d9DMuGthI18HGSu+O3AFWjE8i81VHIoVEOTcsvH9VsGkzPNKblxYvgUbh9ZqUkMo
yaYYrbI361PN2CjtMgjym2d05CGA2LxMNJfH4GiUfaqAwETjwHXxys3SVjJKDkV2
7cOb6zte0+7bX6u8HSaCU90LLiE/WqJeMCC62VQ8MW8O277uHLx35M9lNmfCrkUK
9xvo4F6QaxJkHlTDD711XNyP54yK41rdXbL5FiSPL5MnqrCklT8jRcs/iakOGT4S
0XlzWVkgmesBfZ5kX4V7WyAjXiz5RHJ66fl+vxxLuNjQ6LCfCSUmhUIvN88jRFTq
ldZwZB+05tC/RcXOZBO8wbhVayxNpWjVOX+CuJns+uEGpa9sr45C0q9mAu0XZdLK
DyKV6QxMeSDLCYDEKClKGTn69hWl+Qh9pqhWMcq5lkibsNkC9c4xDVhz6j1P6MiQ
M966NFDybZeSxkDBKQMBS3TYjrS0ys7yJZvYmIh09zF6vlhAbHHewlbXOLAKFTFX
ZdCOjETi3W0mvsmbi5AKYpM+8s/G4xcaTw218hfI+6PdMfX4dq44/LMj60spjXq/
5N04ivPiIQQNvZkRLaOHo+haebBp8hY6FrnU7n2GEJAPRxMq4G0nyMm43Q/CnGyM
GL+bg/fyUG5GcMcfxBgTzU59CClgoH/V4b45skHBgw8V+KnMY+d/TrL3stOPJz8j
e8g+lifcilc4Y39G56InfcYngQ4X3xFkV/GAsFdiHkhDKTl9qHq/qTFH444ENQ20
f27c/WbjZ70MXD4szw2sAqRUt2iqFCWATTKL2S5PDLRA88HS2pUNpM6jONGem9pH
I9Uoa6fNmKX/u4RGb1adqO7bYzcNM2Nt7wa94jZWLlSV3I6FG9VquIO7QVRVoW7I
r/UUEpxP6lRY/TLr464PxXGD15xhjJZSBGISBaW8qOovauUFoxHJGSzi1RKmfcEO
pYgN0PvkgJZ6T389DzOhyi1fpusNe2+gDzjnu/zy397j/g3GiIwAhMUFKRl+nACP
27AQu5PULhGeerQCwqlvOFFyvXQ27ey1+IUZOBuDYtLShPXtrI4/2eu5CN2b5vZ6
bLBFBTfKP9Z7rombf2k8fEisVcdk47eZ/mIiYAbqUiLg772PbT/9hRH/esWtO/pX
wPum3dDfdhicTR/TDXXGu0JYBnqDzrfX+3AVKf7wjzbXa6q11FVBj7rdai/Q6w9i
Cm7BgPJZ4BXmhQWK3IPpw8d1USFBKNe0m6V5D6Fy5EVCikS6iTwREAVVaf7M7qmm
YI022g/vtRr6dkYPazYPv7UbTvwg7AbFyrXCPabmctWZ5d7dWopCO6JSCZZ1d4KN
JHNUZM0dHEWNxGQWbZl0cgF4Mq4Y6djSJ7cD2VqyRPeAnn2175s7r3LpWQQN5Bot
5H6ZPzsq+V6fA5tYj8Biz4RVlqOpr3jxNA5gZvmUlbNAWrgc/oJlteJlfcRGQCeb
fVjcOsxrEbPicynDBeJttlFiY0OVJhVsn/XeQLxg8oWstS6+yVVFo/CCY1h1Xdpz
JV4kU/Ev9QRrxmpaaVYcZTJDPzrKtzBKItCAo2Yvlixwnd1PXlBPnrnHIQBp3l+Z
HnoFF9t0dBACWbgyMJoligi+xtF2g81fLSIwYezy6xo8JXNMgUSJ2O1EkZsWZiiV
TDPVHEP1ZNjouEnb/YkAdUeQ5GvzoWqASEOL7rzdWAAabMW0hdaBWsv48lVbf+CL
+mxt1AqF8FGmFyN4PVhcVB2dy8Ww09huphp4PNVaI7mhRTNWvGhvhSGyaRZLmE4M
RBMYxNPz3hobiAhzIa4FYHoaMxtJGNUCzOnwqiGpaG8/8aHkJdDdXtKvERo03Ai7
9NBZG1hbOwZd0QPaS8R4sO9rGEnmaFP501EIEfl66+i4ndz26tzKK9PIp7+PrB85
Oj1KFXiVXIntvZEZjXD2a/DSfWA4/oBtWXxvpw3q90DyLnH5Y76g9zusUxN8eA2v
cqleD1CUH4tQhryoMpxoLkGpBjfohuYWBi2Iseof4sLf0a4K12VuSEwcnn6av0pH
neSFIpaT1N4KILDtGlzN+oddwOOYKOKmAvAxVRl/1qQ1+4RxT9Zbzy0aRj2ZbeUm
V4/DvlLploFV92vX7EmgydjDckrdnJNrazNOaXKhrkwJpTZ99RLpfq/7NAou92z0
2VuUNsKolZMkgG8npFDuaWj1sGXBsyndksNt0x9U7t4mtV6OyQCFlNEm0Wi++VBb
r9YUwiNCX68iOJ2kBJWtiV3yxvn8qrgFPawA3w9EYvY70k24++W+b0wGQvsOj3VM
8+gkS53L9wLdhyaPfwSyGOeQFvScF8DNT3STlwCbcvOLjuDXvIiSYaUB/svSWxaa
M8eOpoP4i9fn+rY9/fxuMhl4UsryZ/15in7i4SqdMzrNM026aLgYEXZecHqE1RFV
hkYda8kj4UEAK/LU/LKkAjQ6ZVLR0WCwtpOiDJc4h8Suu45/K1HN3uf2b0N5ooS7
/oJByensJ3nI/zmiTmSGq+d/CpnbnNAvxVkK0AynDhdcDAXarOjXR/bogRcCMe70
ixDK6g6LVeLpzU1uKTBzjRd8yzf/3hr2V+mlo2wtdPC1F4Ek3+Iwcg1QzAU/lK/y
nH7ozTDGk6djpu0WuQhDScyuVXgND1UHOAL6XDEZsbp6f7Gby2ITsU+b85RLKBva
buUlpHgLIYhmcfPDTrz91Ig8f0o1x0qk8usJRJEt3LVvN4UTQgoaQu2TmNADwetq
5xm6nCEgLucXvfa+8HVDdqaV7nF3VPaZFzJRZghucvVzJvLsFLXV1jNrJuXFujdu
DcAZxtIX1tiJ8se1OumiFSXtCTkxEFT9MA5V4hpddDPjzxDnE1+0fX0wZFiQoWfZ
Xsow0u4jWtrUrNXT2mU1wab4CFZKDyuBuSJRfxO2zKU+qhQPUq/w09Yap5DGtNhj
1DicRFUZMw91vsmBi1cgiod8mZGzT/MaDOo7PD6eAuSZELtigzjkYMoePu0dlwV2
ZftzzPC2vpQ8XytzG6ZJYgUn9SEf6sMSDqcZtC4Sz7M3jm0SD30g+RP/6D1qF2Nw
kOnOnlaRkdYyZscwUiy0TxMSOaKRQUAYpI+XofoepzcDWo78tp305iteJR4JYtq9
QbKPryj+8Xd7UCL51s0t0H303Ud7n8vClESuG6ELr76ARDLMwihBtQ+lGetxoVfW
R2VYEcwGh2J3fjeb5HAyWUhHbQdVn8YjpGGiZFLQtnu1m/AuCrps4yNSNVHmPnU4
UL1zGurk5EwhA1OGFEM3utGa8V0kIu9l4rMaHPwBqI1LYwxh/yFteqehZVsA9A3Y
SHG3ISfUMGrigZITERWuN/GQkCM98KW4f3MDA7Plmjy//WhR2/2pOizKLqJHg+4C
ZzI5dpdLcQg6IdkuLU2C++Rjvs3FR33z9eB4Zt6vFMDM0kLk5lcBBUrLfrR/XuvZ
s1gKTlRn0NiugTnYlBi3rOQzr8ul2eCgF2EZVW9K0+mOY0kHSNiQoOuX7fn87Qts
MPKoodikUHWHyOD5WJdxg20IQjlV/2EHvb6i1Ucm2MBtSxIh/kZNREokImiYNCGJ
/mIW+/dBZO84gyl8y70cS9T0QLnqpcDn30k85yrA/myBnFdKo+hh3SpQKTU11BjX
MKqWJOuXc1wPTTb0qq/oke+P0ejFppIjnW5qnJjAl3LMq2psOXOgXd4j9W/N3t2U
AT9kvNsws1WrJqNodmvytbJ2/LlhkRFkz0w2/x3YHloK52MfWwRWcC7ZgOOPncyn
u4l200K+v4I3v4ae99DrHruXLG1LmDiZPzldfvqAhR5bsK4kn5s9NobPpIh62V4M
V9fCdaNEeOrlMQj3TMKlZxG6ezu8lKcsELP9pEkHI/E2ENkPGJPscHl3950EKobs
qDz70LLJ2wYl99h1aiunSo/wEVmfD4jiYbWmG6CoPi1AdIFGRHx2iVK+K7aKDk2q
3eqNpKSiNgyrcqLe2mxPTiD2IVM8jsS1xXpnqyMyfVW+GvhIaF/m4XDEwdbUAWOc
P65GWhj9UXZbl6sFylXT/kxgDWhx/91qcH8DWy6jyjMnacIGZPwHiBVkQ1He99y+
SyYodM8DveeVbYpqsX4NwRsChP/3lJD9JAAP+er2wj1Os3fqDidD2lh/DWRQ3B3+
N0XO2LsaZE+Y9Xepg/094P5RDcdbkWeDMNklBqWUiJRgBjf5R0l/zKiFpJT06Jdl
4tSf2wk41bVtnV2QYToGPmXSzRy6vB9cZeIVBL4OgJhTSKPhQaCTbXc2mwnycwJg
xeDCCP/uSHIxt3UC30/1Ki1nDtvBOJNL6YALLnVtMrt8oJ84HA4ZTW9TJd0mvkZ+
2DuHCbHghBTXfBkvzfwG5zbqKgleYKHdOBLhrOTN/NnOLwGgnqRwY1i+gWPD+wuQ
fv1ghcm8Q87ERKFqyQGtMVrjTAgoWZIIRRUDO8PaCVC3KR0qWk6Y8a8x3NKt985/
J6kc2ArY4rJdLXg1CtiXsf2C3ChtYE78ng1LlLZxAmlGeTaVBaMOXrOAd31edc9p
R4O0usvBkM2wfkew9rm1erml0ojEj6JFO40ZRldRwjWfbLJlFWI3DVGUXoBWyARf
I4DqVuTrVq4vCG6MQFdjJJ46A0agf9W+1q8j6v7XxlPtgCwUOEdA6HSNUoS3xMbq
THEJ37JyRIn2Z0A1td0OwaKN2M1KxXMe/wPL3MyLvZ3ruDL7QBnWPdlREBYM2MlG
lzb5AnrE7urEbUWOU9KGwaq84hLK3O9Byh1yZaU3S2nBb4WitABpqGOlzzyyj9O3
sdLTG4lY2AnVxR80VylnHWqQTqyWIbHuIQtGyZnJxtSanrdvhBBqPzG9K8Yx0Ywg
BU6dqDH5YBDCPvYh5MxnxWRW0UdJbAQIRaoqiOT3W9umk5+qxwXJL6M7+uCGoKdI
/ABS6wKQ4rxghxnwq86P4Tx9TFvYfvRaYwpKw2eyv/30hXVnvkdehENwFZVCfXFx
RipzrI7eZfw/LJpvFPFZJ+RWi1l7kh1iDuGXV/86NEkZBL68TAepVW5ymv9sp/rL
FqhnyfkjhzOi/dZGXqRQMCF2SJVAR7N2HvmkKIVoQCLq4QSgLkT8Vs/lh8/Mxkhg
M0E02qSHKvG3km+Sw6NWZyjNWStzkA5+NwivzHZpsbmaPuYzk1C3q8Khpi2rUdA2
V+1vlENBdgtwtHCkwU6aWei8CWEii6QH4cVfC5mthmm+Ufm3cgMm8jNfo5D8VjZ+
W8Bf+ppxW14RMxU9TXabEh7LWq2Vnl7MsDi69/RBOPWtQksm8aNGVMqBq209h5Km
kO7s0lCwd5dTcq8Esofaxl+iTGn5XU6seTPGPWEOwVSKyYK7Y0TUSoQ1OpriTOVs
JewLw559xspwzcOyBo5nmrZOcf5/NaBlXtuFF1bRIcMQ04yyyg8GyRKtM2Kmv4Tu
yfEFgxhbMVUryuEMNtjo7aXWGU5u394mHNlUwJmfx/j15oiYwvIBFR3hdDKjJK0x
IYYga2iJty5Q68zQJ2TkGeuKnPs+/KCSu5OuQMT0iIn507FFu595rtmFBa5MOzqw
yQHS1P5PrYEQOh2oV4mmdfSX1M16hLx+5IKRXxBuZy3yr2MNcnzZGgPrXvOrgW72
mqQsx8yGHUKsisQ1RRBXvjVAeRksHYYdHnz0FFmh1jBr0fFgCMrBpBeBUh0Eye0y
iKmB9Hhp9XUP/45a3Pj3C1zMuQBce2c4h9UEp26qSnxQRKct9k3vqNmERBcbfVkt
w7ActLtdG52SpRz08Z26GVxcmeGYPOGJk5Xi9zx0jwMMtk9BNLi1fvwDg/uy796r
sUtsRFXlcug78AOUeCZieVymlphsqmbS9aXAnHymBszg6NIYCS7jGcOOe4PKlM9p
3Voe/CHQjbAGUG/R0WGkGg2AzWW4N15mTsT9cgvaaxQsQJGBjxm0oj+y3SjZ67UP
AqQL7xrqb7R37Gb/25KGlIhoN+seYz5yZOFEWl0Cf0JymoLO5aHGk6G0cohz6IUX
8eKvW51XiS0t2+KMln2cunwR4KrehGla+fKBi8y/VqlOaMsZLCnlPPt71fG7qWLA
+YOSz33Q7cM5FBLQeVp9eGfMwIxLjfgYktv70d/Sl53oXiy/fOpelV543tkcISV6
Djf76fa2OcD55LdCYYu43A2C0UNfFM24sn+SExsGcCaQE5MsPjZuF6uekgL6zlVr
sPx2mQ966wcWvixFCKBrZlO23bp8AFDm4gTNJuQRgGMPw3L7YRIODAvUum8tZD37
VeuiQOUotPdn6mKuCIeQeskQdrNQVJ3ySg57Xyb4XsLQ8J4ghhn64Exh/RDD9va6
OkjYgz3ei0Mg3g4+ndYo/WbXEC1dN2mB5TlTUuGXzVrzd+8XWXU6UaycqceRp/jQ
LZNfbwCUZForabISq9HMlqs+nQ+VDrFi0I9uhpj3MHleYa/+5TEbbxp1ClNcthLo
3cF7HK0eTc9cquKT8PW9VdJl6K6Y5UxBOmXvTpZfHGy4zke1+BS7VujCTygRdTtg
VE9Olf9Ak61pheCyC6p9G2aAhYoiweelnOOL/vxiC/nIshwShN9T1PCOunR/ZrDX
abreavLy8LZPkGUk2OTqkQOMr1xYXQ+aowgmT74+QvLHoAHYml+Z3WZ+og7Zc/BO
RHnN/PiF3ZmPZ329Z18vKvMhtJbpUYadacxKu4+aDuRg57MwhjD4xPQ0DUgaA2PA
k4AaUvJaTNAmkQgNS4R2nZhi4qmnHWb24l35NkVLyqK9oFdishggxLnczN5SXwRm
m/Ab01CmnjahFmCrFpwU8krAKOGr8J6/yWdTd51zQPgqeMXsJuHAHlZz4TKM4zWa
123jykjP8ZUwK9OcOUrn6CsRKADG3IuLY+vRbr8EK5n2P3xABW6T/YRMsxzxKvob
TgJcvJtrfIYcvDI8dcTSE4oLq/J0j6iy554y2N/C7AAxPdHMIe9xH8Kke8LtqI1F
2sHadM7nPXk9bORJvX4EiDc59o4wQ365qz8X5iNKtaeEGZS1TeaBUZUjp/0CXYDH
rJ0r6uQpGAyDlKC1+9DZM9NcbIfaGH9YK9bOB8tUgvnTv4cSW75N1lh76LEn/VgA
zhTE1MOWx0iozk88upfbUnhvATXmgkGdRnTY9UDYK2VfDjCexBRTUWLKDWEy6a9d
b8/1TKkaVNQYlbsXL0gP6B62cJUPzbo4VDXcDpvnce3nWwpPsWMAyVUB1dKbFGiK
2T2MUoxGIjv8gFzPb0Y9FXU9IhMNNTqzc1YLaAMilx417AeeROz9qWEBaRe426oa
rMHy0PQ9QNrykzwHIyjP95tGxbCqvtNUnRro6UcUlI3U77qgfExjg16n6nDc+MBj
DrXG3YPhhOZtomeb330ODBhmy9LkzsrahQyoadav2yCYglDcytZZQGpQAPrVxtEm
kf1a9NExjdk0WQEUFig8ukOnDZzJIRQxCLx6FVKwA3i08QMUcu/OPN+lUjfXBhgn
4VyGskAXmqIKR/WdQO41sNmi2Kc03PfTjS/d77vMV/fBzlWR6qrj1Bv3ilx3uqkC
lkq8VsHAG+eKA9HmyqZkouQW0fQ8qs+9v3ENSNjZSkr3obQVZ25So2ljnlUtKN3x
QJU9TJOVJQCF2Wz3daTcW/FOg02SEmXB3oq0s31IeYaxioVWVMQh+rKiLcxNOwtk
2LaSt7wo6vjGAs0MOgOlgPZeqCwjVLz9EUOdry7U24iOyOFOz6KBFGKC0tev/tOZ
4/yHD+Vvyhs8kpiayNEbDMFv9nO5rNGw+O664KRs4UlM3Pl8kxgG6WYRm7/NCPyh
cyWBPmyB39+l+8hAwh9IMYOGOlHcRqKOl+8zunZwAQffT+okC2TKORJMG4q6KeAr
UCOQEaoyYRa5SVq6FM4o/VfOFUPOwJuQRQLIIOO98sc4X6a8JLQ2zLKDEWKNb+0y
DhZ2A1oaaMvz1nPkP519nqjCD8U96HaEd3L3oDYBxmExpOyzkT8tzElz759j8rEZ
NqL93HN8CB3tnnPTFFyKfhbXgEsfdGE09/ztOzzGrznRzCC8fzOkKIz7pOYsTrIb
J1/p7WaUEbFdCheQHPNGb6Vv4g4PoJLUtk14k0IRgAgdxBQdhAz6CUdCkfoUYMyf
aeiYFG/9mJFskVLStoBHwapKeg1uYg47rOd5zMZtEz0sSEvnOwyQ352zKeYEpCgN
9VY3DqJNm3Y+8JYTjCzSg7eFnIG24LIwJXm5Luv0EvEHPfyZNNRW2mZl+YfRJ2iY
G+5rh5bC4w5Fn6pcI1b2wf5Tdk1gQxnYKR5vVyyjoRtR0EnpPIqyMHv07Hd7FRCb
Ldh+fkg2lrROlaYLbRQbAdnS0NoHPcDotu2fEJ9jdwp3nzRtNynoW25LjY2wtdH3
cfRn4AR/b1ZKWqMruCUjovZvq0KHHzTRgC2jnwMQIt8+tDJrs5in7ml6n0LJIr5L
evewkHDa9yyjXZUqEr1bixwdpYB7F+fJoJxSqcBokD2OybR7ZGXLkKI6rwukw4qO
kW3XtRZ7eS3HFTyMv3k9ru6pF3Ovy2cDVaT5fjDuaTO5+LdcExIWo+ZJL1ejdzmN
a3nrs1g1nwsKhmqkTQ1QWH9npTytlBd21fiYGdx+7NkV++4PoVRCQ2HcamTVXXx2
mv1RwpcjSKfqbW70u7WYHssTctO6P9QNcGJVlHpNRDBEoQiN94ehtZuuHKpZdLix
pwf2dmOT1MKo2t4iNuAoBYpyT69PinGuGBmuN7RhF4Dm1TW8tE7p14vP2AsXQTAv
kTh4VIOaBWbQAFOn3O3rWKWAvEGg5vO8AqdlvBipoGc4hRg593dDWbyRXo6Bl6eR
V0AokAQ8Wrum32vSS1orBHpjm2Pq/xzEcrGHEWZFDRcsYUF9wefcDTaAdXr9fpmg
uU3dlH21AuSPw1TYfGovr24OQP+KhDkLzFNk8KnAhlAyhXuIVEHzmHwPbZJ7VVrW
K4Pvawt2thHllQN/XHPBzZhxAIo3UJendOjr+WO7WM2v+Dx9UMIOz78cOlQNGDCv
Cd9blFGalAefVunTiPOxTGeJbpLN6/EHnXJh9bn7xvOSc2IaeQUGkTOP4KrkJE7r
CZyWKVJ10+RayJD+he0luZ2f7s+u1jUQNRZm8v79TH967D6nsga2qP2uXocfRv44
WWeCmLt5OXF2prmbFpGVgp2h3PIlvQEUwCsw9hlsRtdYUyXCwZCZJD8oUyJoi1nw
8IEsnZ5CuWrqA+ROeogjlM+27oom8H2FBFcij8kmIh5cHhtDYkiHlPgXvSKcgOIZ
8qJ0cTU9JJYF66UY6S95RRn1AOLa12ojPoKlN3q6cdRl5C6SfPrLpZX0SRm8dZ6m
8eHQ7KS9jtIKIHdVNQnvad4ZwpiV5Je1Q9r2eDOMBDFV6O23Hrht1RFX2aN7XAOC
L3W82Y/+Yt1rLzisSRfqC8wimoLB2MQ8PCDHODN4HJZm4o7ZncZp71BzaQd6jyfJ
Q4SB6aJnoY8Kmu/y9Ig5ziHGHIs458Q7y250ZFHi8KZkxY0Np7ejWcNWRu8iv80W
flQ9DaHAVTa40e7Rudad0Gjq//Nimr7WP98i4q6caOv1wcbOW2TD6zm4Ecsast+Q
pXruabcEKbGsQI+aWoA5NAcmrFThLm3MBUVZaHx+CmDmEBb8mz32rs7B4BKabkb/
IA0XIPDwclWmHeO7C0CRuIoB9gcbPAu9z99nX41kwbsfOuBebh4TL3LvPZsue7VB
gAlL7xlgnfzNDxpUUVjIpyMg4TdNgIhpQg7heloPNUrwzNtzBX9JFH9n0neHu69U
k28cdKVAN7YXogEBHLtQ48ueXghDaY2Lc67nX6+qgRhQbCADt9ekU/9mvmJEg7o8
L2taYdWYv/nK/AxS5aPiudZM3eEgCWsMYrjngntTyyr0zch5kyiHAKgP5gysc4Ds
ZqITNFdz6lqzOPiT1d4o40UYXZaDvYgcdfWrb3K01kM3Ww5cse4ZqQ564Xzb2Uha
3wTNUsVkvcDnAD5hKaOb7psI0bRoOb4LAQiFbrR18/5iN93TyHh/sKUNRnBvOAzW
bkzN00Ywd92EUnUrZSO78BHExtup141StNgIXkylOGMyYHZAdcECY4+FyWH+HTWc
QSFaPgYxAzEhsedh/bpvIdpL1W2bbjYCzm9zIwv4R5QGe/NBHVya/XGSVyQ7ovh8
9D7pECRQF9JstXdI3t+9+xEEi6D5sluzhhmNwUSezHHqQVvCsl+BtesHAZ/0KH8u
ZU2KjnP/G1l7+FSWLIASWyPcyJhjR8ljTQNfKNFTcoeACnR4RnLZT4Vu2XE5abEr
gh3sstXIbAxnjoGFSvTcBdB7UgeMtja85ERNpmogXAQZYXXThculHqwDIMajGqZV
tvkPrXjLsrWc3zZLnrzFV+kYORJFfvMtqEQ7WSpPppVplQYGFVYTPewcDfK8Pw1F
FNLJVcgFwZLRVsXU8ZzzI27hawciVvaqh2snWbNaMBbNAdhTbkCd8STO41h7Oz+w
IDNQ+PuQoGH7X9762shJaXHBskCp1K7+Xti3eI55lOOZC8c6HQWxIYR9UbaH3xs5
RmktWUp/pnZqp/3/BJthHGmMI7T2fzx6xtpbSnMnu2vB69C26fDHaY8eQkbxig5h
MADqPSu7k5ZF567k95sREXODte1bw4SSvyMB4QQ97poWfNvvoYhhw9Wg7c4L6BNI
rdUiexi2uQ8lwH/RaSi4lcL9x/uxCN1NDTQTqGKc/TIgIrpn30+g+SUuO7FynHvq
cSXdM/aPlbuIYuWyDRLa3Gkee5vNFGTM21yFdg8+KRNb8vP7Q7/+eIfKM3XZarS6
nk9hxnKSnuwq6XjNuuz7yWzwWSawvlciaxextbL237VzDkOXiY6N3uvwndUJLyng
bIXGtt7JSSZzjL2qxYVOVyZkxMaiOGlEafnwdbTExf/urCPHklxm/f6xbqMLddld
tqw2EFKyhNJReidvrCUygNbZC2HYYwk/MLaKiZ6bM23QIzYgZI/KurkJ0wXSPv8c
v3pgaJs7FptsVp+9e0uqhtz0q8L9PZtqFwrH99m4LSS4lHPJU5vlMwlxVsDXekj9
XrwsIL9p35X+CPcT75nBnsevqcJ8p7zTYl0fbMhSQEqzk0t1gSZdO8LUVZ25Otpr
b6jaeRfbdF6KKP5qxg7eopDN4W7M85ot1JDR1pmZHPkvXLk8ThipDD2DXsKAlfrQ
Ra/sx2fX5mZp7e/mZXYbs3j38Sx/TiJPq4XRnC+0mrvp9sit08LyLNnf8qdu6mb/
IcfcZGTUhmEDnBdDcYvvQ2VpG6j7FW0viYClD/gzz+qn/MebmMF/X0njTDBiDVLN
6Qk7LeDnBw/mLdH3qoR2HBlq3eZNjQftOkyy1UaQ2wCwW6aNgmL0wLQ1A5m7kJre
ImfKR8r3ahTLAz2x6JFebHcvJigyKceoPyytCI93SJyXTnfgiT8ITw+x5EPvA/6U
iraAviHfmrrjQ8E/GlR0XO+gEvUGkMU0+TV9mqubQk/YPrjZ0zmLaJwwPcOrS/3S
QCMRAFBiXiNSh3xE0R6lgakoDCyw7Ce2oFSu/Ii/7Nd1eWt948rqfY3+aBTGXnHo
X/SDdCccr3vq5belNhPfdcujNamENmejsJPbzTMxzLLREojXTLZD5PSKUvLMGkef
KlRPN+DeP4lHvWn4XZS/Fsr91HzLHGBWWjgDERZFQhUCFXyu3vGeEGNwj/xLxx+U
CZtjpJnzpCa2Jj6ebO6Ys9CLknT9ITSSMn9UKpPgUf4KGFf5hM1fyG7skcZgD7wK
SfirBendeu5gtDTyo+cmR0BSYpNB+TvaTrl0+9bU8p8U4vlP00HKQbtCg8+9j6lp
q3BPkemch9E2jBxm9E++gar/GI6zzxU0lbS1PP+JtN+Yq6FGLmQRvng81O2aay8A
NsrVUy8VneFvnEnDHW9jw2/JtLbMEj1Ua7qP8NYzayCcp0s2zgbMRl7vm0Z+mx2I
K4CbU5C47yof+4sbFsfCawIQxiJvhs3fP+qamKMg5tQwS3Qv3taGsrqgBERrlC8u
TjKIaaQVFxlt5c94uiZgJAR+65SCMHjsa/LaBeKjvA54ZX6+NM1UYBrYE4RcrGPo
ckayHAWeGDrT6oab4lIRrchZhb2AqCB7ipM1I3mA2TRuTW2mYHJCIUq6Sp+LCEy6
9ZuGzzeExeSUktNDadQo/OTtxDALxqPiIiPs8VJ0JAFgeerkqooJr10G9z4MfUl9
VFd9CJuaNE5oHZZVACeMzSwlKVtE+TUbmYS3YUQ483IUhdcFMEaCCFzvJYxxcOvO
gFWArQ1GM0ixOQPlsNNXom8VZy/nbLqgctQhXioHN4tR0Xl5IB5zDnQtyueazU2B
5q76i6v37yc/2JeV3JUGCflWsHTTVA4knN/wxKJ/nFNsbNcQgcTeJDpJKNSum77s
PImKIdi+3fi1/4dhWYlWoS2Bk86Jaz0DtiTXoMZLNekKKj2jXn94swUQXaI+QV9Y
r21lt7lgjmwUXautllq9ALAhKR2sT2BELdKafLz6WyYAN+xFrX761YS1sGXECAl+
5HYvOroVVmYHaJxr/8lXxK4PpDbH2QeuGsUB1dUO95OmZWY1ldgGP67aNdEjZBSS
6CU6P3tV/x1Yq4mWX9r7WFN6WSrY3p+vK/Ox0KZj6dLkO6gndX5MFPY4tdj9UEPv
COIQg1eJPQTlSTC1/Iz4lJ3RWLXju8cLkY9FChIKUX4Uraf08G21c+GaTNdJT0sB
g/ryYaSwtCXgsG2m1IrbNFDfBiA3oCCutFC8z2PfJCpBCI86ylI4PdhnV1KVl15f
svwBUIjkfxKJb4hevpAkA6LM7QK+b9hUic+xw41QhITGSEve2X2JC0MbYwDv7Wgg
gcCFFZ8ZwbTVMTZ5ijW3KeBt//nHEuyjgYMVDZ2DZVDm2BGjwZY/2DZ+6eXwau+7
ajBNLLAbUXmbH2gAAsO97XyNsECYIKarhNxnSpAbIxEHyZG34KJct/Si0LpvDuvp
iQAk8cFdgyckJFCwHiNdOBrZPeZ+zGxVCmZT1Tk/3aZZ1NVwmoi1prq1gJVLeC2+
PIpX6vqUb4U0K0+Qe79aL8F0KFxPhIrGlSdmNWIJAWiRc52fmSMO8u5rVuXYSPdx
7yGCEz9EmA0d75WubqQlMXwRpDFIfMRgsZTl25ll6eA1bVGqKSqXuiQNq0DMUw0F
T6mlfTVgjbrfs/L42okKQUoX6a3Y/sveqaJLkoXTxBY/l1tWh5JODreYsUTiJB0n
E31tJjxFhEuYzODDO87tVUU0huuM4tYapxPSrRvRMCvcxUArb6RzoMfBe/WmRvdw
X34/DDtVuQlRXY0mDTg4206MQZ/FjoH0yyWnWM37WD8mFg1eJsY25Scdc4R9Pj7K
MAUPpxclZM2MR2LxQ2tAeGG6aSKnRbi7CT8WLEXuckvf53E1Ie8ZgGHEbLmu1u5k
WVBidLnsbmo/b+mJB6tnQ+1kDpMHNJpitY/aodaMXm7dmH3wlIUKT1TjJEl5KeUO
cIBBN+oj35JUYjeFuo4wHf4FmkGlTAdErfO+9ZJjaYrbM6JgDBrgiza2oVI/mEEr
fn5GqDC7SFIHSdDAYto9pq8u0f1YRAFPIRs28chvP0yOSJ38EVHsYGE/07oDLkaB
zgf1oXbis1XFdZqnCh6Cqj8pOMOPk9UIf2Qs5qxkLD+bPp6skriXunWz4jc1RB5A
PMqimm2h716uuoAqn5xCzSAkkAi8eDgbVmqNaJZKiyo8LdcRKXbvjdTEHA1R2bV6
F0D+UAIW4iMSDisw48BaGr/KYstetatKqapGYGF7T6AHRYQbcNf2sUdnC25uguZU
9RgMuMrvm07Tbi8qdgRfkMCG2LAZOqoZpcyPNZylgqDiZiRUi+yb+1H3OeW3hRCR
6jpbpypS5HlU3cow9GR+U5syNY7obFBcqyShkhoBn4oQ/wUgt4tyaG74V0VdZoiR
AGPh1mvoAD2zMHmuPoMrHzyskHWXndlwRkMp708Lg4G6/l995ejWwtTBIPxKCnDz
JI+MyZWM2VjElydBt9yOqxELYeR6K3n+Bo4rupLOSAfbC+eMIUP9W08BuzRM9GcJ
fazbgpGwjo+6sAm5DRmXypssOurH5PiyfbkEOhkPiz0izkDZRfQeyWaIVEFjOBzg
26/cXHsMYX9HIOYu1CUobdXWRV890l/ET5dWo9qwY8VJRANVnaVlBJ8MbJOGQfUA
vnWh4cMRucqU7E36lJWgzG45u60hqF3ZFJCZDHURmZEJhM8kdKCYy4OnfrZXz+8E
uqtt+tGll7OWB5ghWFhXu3gNgebMq+L2LRGV+dKgfY+rLZ3HUoGb+pqv8TayRLyD
L5GMjVhT2gw92Y8WOtsGwGR6tAeZ6CSgJt8qDMOAPEzikO9vpP0bVMCGqCi9ejA3
IYrgNlSDR6QD3KyfBImScA7TpSFb1EoQXmqfdT1j/GzaK+Hz3waE5qGXDgy1oG3n
bXFI7p/WPMZyrC7dUkpa6Tw04pKjqsJtr43kwt/cSKn6ofSZXuYi9ICvw9ZUGl1S
xxOZNEwdl+QQ+axTMdMEKQfP3iR9Vf0Ip+XggyEjwRUHW1raNo4ZMBNtAV4xZ7+I
4SYIjdJB8UhrcXhMjGGawshaIOwx8i7ducV8Pj/AV4Wc2lK61lP3G5jRT6s6gB3B
3koGuAPMIzpr0ijhOyzvYSp3mnY66U544jvwELfr5AYymuH/CBHFc2j83PZ7dOq1
8Jv2gZxBtLY3pqaM2Zv4ZQEy+wArAcvdtH5Htv29i96Wb0rXQFzcGOW1i6z+ZAtB
KVE8tNXOxN1BkdtoyVb5yg0pAaIXfG87et8tqxd+1lDJfraD02NYs179VzmtY7tP
fNFiB3ZNBVSn7R9iwYVqyE1pBvlCVoJHCLtqwd176wF5wcZzrFcR819rbWJ8y51L
t7rXBBMII7+sSnAxHbI+79ycvhnjnbXkeqsfX7UpiTVUrnqxFHZAXi5trCRel1g/
lPDSdo3MGO5rV8a2EcghZVE2P4cZZsFehkyQwCiJqTWVB/DUxSgZ1pn3x49HEl8t
IdIdfioDJpcFBxb+/Tnfjh55+JRGhwZMAL9cgUDmQJauoLSRu//0aWAdcRhHW9jf
Kwj/pP0QUKK1dNndhwWF32m+4RufOIKuBaCp6iz93RBkj8zJUs7a3q2hCf8AgKj+
Fyrdt5eLMAYVIlJQ4d1uc+86/0RpXyRinS7LLatNxa6CbN2Yq1Dyj8Sn7nuxfOKq
y+in+YuBMOXHkiAaUggkJtbsAw2+B6ixz5lEEdwt4WDWoMfCDUHDOrzLrB59gMTd
8mERuC0ea+q6jVq6Bm6XLh6q1Mw4OLIM0Tr2f9gMa8sGwfCH792DIbiZEJh9OOuq
73IkbXjBiT5ZJFrA7+kSM7z13ehBshprXGGgXY7TwGs8cSls0UrGzxNQzlrsNuwV
UYSbwKSMbUz149DbmDS08MgPGgfM0G+mlc20dPDL2HncdL1rVMgl7zSwII2a4pHC
sFuL+m/sky1rr+CTvVav6KKanDlh2YayYIVrcquRo2HGaU9LouvbUi9n4JaR0+2K
hxsksady4MIu13ZcJdoQDpkbso5EmwJ6u1YRPX7G78JmGFR/xgzGYNyc27iP9Ijm
kpcW3blOhl7kGEdgiJApZJc9jeF4Or5Vgu759YvHQxRb62q4ynd2QNAWZiMd55tN
h83BpFHuZBag8XZDL6s7rLxP+Z6w9oKAFWe+WN8BxoOgYvPjoCcp9eOpHQraBp8/
eoJ1DIbkSbiD+wZE1HN6DMsAex7VdbG+ochF4VLlckCFDam/yAJiUB41vAGJX2Bb
Qtcxa2rX9jTfX3vrW060eZa0DddHsIRO2WTfC5lHN2Yenh/3n9IMcwO0wIb2ItfZ
dz9mACxoQOXf7n59JyyO12PCdhCrTVmDqzLTSk9RrfgELRkxs/xVJCXiCt6sYb/1
kzKFj87bPCPt8SzPuic9gWneK8/ZwDX9MJd+Qp2I3YwqwV2aEkzG9Kys8Xt4M0e+
uNjxMij1HH0etvjBMZ5YIe8DGqS9NlHpB/pUv6kbESFuutqZyqwvYmsTdkafRkcG
Ko2XHFYhxsODQgxH5Y04r3Kg3vUg2TcEKqFmXXP3JxDi0RkAfEs9M5RxCEsvqDDs
qzAyc+P7Fnm9asbC4IBlOEHo1/M5fXnY1LOI+3W5EBl3Qdm1E11Bw3/Zjki0YZjl
kyrjBf/nvgoLRDimJUqycHrOGed1PjdFXhP22dYP2+7QmzBMMMEI5DsdHE08AaNb
N7iAGf0K5q7FLIKdoHjT33l5Wxk+vQBW8rQXA3pQnmGOH6ryGIETM3fRtXz3U198
lPrPz+uS2owfUhYc1J8rvEhfo1KPmMvVDbKi25GtH2q5cXSPvXd0LD9QYmEQ968o
lQXRMoGihYNP7i3/N404qJQuQzElttMaqWv30IsrrcCEpibZFXg3iv3d+zdfD8GC
rklA/umMS+wle3m/Q+0oGvGdTyQjbzOxDjKC1i4f+9QDDQtolzQCmpsaFEgc+ijw
Tg+6KvXaB59nQoWCGdkGMKCh/j6R/XRlk3K114ayBx7zM5lTvN39fUBgzwJnGnRH
wiOhcHWgqgpn7Wvw6hfspMK1QY1KzcafLs1kaY6kFDIIorPeKLSEfh7+yg0wyWDQ
LujBW8bPsRbu6vZ0RdI6nXnQee10zLD4gEISDSy5f92hlQ3rryMFL2Erko+vjaqC
13TK2RSPAemDqWt9sHR/I29j7UxyzzAhNY2dyJPhKnAAe48PUcTt1+Tumev7hk8U
Fw3a5uGjb//KUQOBVucd6eCJMap9QV+6TVxls9o9Oo/MeuIC8ILauYzrSF9fkKkL
BZO+EAYToXVzYMrfLIt4+vqGt0Y2MQdsauQ3C2PZv1/1bDMPMy45BowBckQls5yp
9WvogQRv3SD2F8N9PcrBmTJgyKXHCh7x8LM8X3sf/mbyBKujApEeqbCOvhbZkEja
TKU+tY5QqyhKGrBEDqgWHqIcfZZ2zbwYeAOA6EbeVcT2c1Ke68KhdL5vmxI2hJhx
2P0v+OYfm5oGR7pzfIE2iEj/q2macCMGAMQB7X5lYsnlnaUxM1IoTmOrYz1KE+Kx
OxZBy10EyC5i5s21m+9D+5nDU5kAlal2jqTG8IpWbMFtvWjX3SgVRBJjlLjM4jxR
FLh8V4PBrihLXsdQqsBW4lYlHeBF9mBEXnwUvEy2dh6rhJvMYqrC6pc3cmBHGaSf
Ddi1EBnIVVXG3o/UMEZ2oN1+92e/Oz7aSGhW7Fizy28UahVaup6T1a6itYfCHOVJ
dsSvF5aDhHwYnQWd/eQutUYq+GfoOuqRFg1qH8IZqyDHMoeEFSdJMZGa9+ZpP6I9
8ooKgb4Pp8cxDlheg/PL/hx94B6/SyL0Rcsxa0xuvLlz+r2ezAl7KBxTyQzGJoNL
JBJ3RusiPYPAM6XXbhfNiZsyS/A8oMiFa+QHSl1syeC5qj8lGCFdM9/y2bf9dCVD
qsPAN9ZvyLQZNbu9xzbiu7NT+KamdjiE9Mkvua561tifDanOcgxclrsOUDzqGu2e
h3g5BDjJxJZbnxM4U79OVgzeoxT9BeHOQdk0Z+rtG30cEdSgvj+mj1+Jz3jgQtf5
l0fB8vl4fHY1jZA1+8PVUmFDgecYDVToZWNMtKGVb7mHbIpTNi52f6wbwRHbFpXY
B6uiP8dU6BkcEVhHMbSZUWmKfnzcK3IQFWji7YjpDLopqTP0yDwEVPDO2cosLfiR
NgAMKbLKKFjT/6QnPflDQd3w9N/mcSt+2IAMvMpo2oe4EgWufMJjYT9SPTwilsib
WlxfPWdQ0ow+S7WKSOD8htRUrX/4XI4CZetwyaTKYQK2dRdac6qPj/idxEKWVTiA
A2XfJ0kEREmO/ERxBBQYh6CfYM4pttPJ6WFrWVLkUHlHSQOY9EmmUGAB5WC0YIOa
jPKbCW25weBom+zQOp5Po9S6GTknDZRcCv+fkYGLB/a76vNXF6yNisvqo4RA0X7O
q47ciuFE30MjHEQtFCrDt/s8USBGkwY1pAS5kCqWbY0X9DNi+wHaL23f5AM5HHkO
v7Uab+YTBx9XWYOnZI1z3EdVlk/zCLJJr1x6yWu3LtN4z9CszGe0POq/5OTek0Wv
TKLrX9WIcRlZDoh/UL8F92I4XcQ4SYSHWpaW5lb4dY0IWY215ZUb1CJ3GZ7a7sfu
BbhJjioRMNO2BruIRKLF3WcsSttHhhTQkG9tvdIZ9t6nzXKaBFrmN9kMp1ZUCctV
AqxlL2/7GyR9ema78PrRMw1EO994JvZMuxitlGePYRbVwArD8uKVeurPM72L9NIr
xP/phqpWhEK/S/o6DSlyJ2J/G9/m9Wc17w+rfJufT8SaCpPcUZkXulPIBCo3laVL
1bUy5jr0IElVzAJdvIcdIZEVO9tBpPY+Kkh0DPv5g/dbioiMEQZaWnUEXH4eHwRH
4DwrbUU85+0K4tj6SQo3m7+7tukrwQs86WeaYrdDhYhpbzKk3lwevppeQJtVZTRj
Vj6/uAmms4zw4GOVxGt/RdyYfatwrFz7ks1kkDkFd+PIVCFtuIQkGm4yNZgGYtug
JER4TDlp93D/EUpvev3sIwk+DCdfL0L2Jj/GUgyvbIxLvq5J+yN1TOg8wMFeBEra
CQrx5/3GcgXzyIHQGqa1aniyt2hYdfq2cdfz0mshPjD7mi1sohbCyP8ImNVORbjg
zctbcVI3f2otFIBYZYl9Q0gfFNTgZ3TAvzmTRUwQier3HLMXC2K9C5EmLtuU3enJ
Qi3HKQ5YSAShWd73r1NAFLyrlJLD/LpIAULrFipcmV6J6Bx1wmeLfXeUcsV8IA2+
h/3TFcCP0BiS62vCEca598+aVmh4WckWpWvENSoIiJ8hhzawhrRXUI8J6y9Zv2Wt
26I2OIGwFHjPbu8+gNhKwvmq4tXmuCMev9WrWMzkR1U2QJE9ntFQpD+YMnvgPKy7
LcqyDrGL7oRxFt4ZFwb4vh1EzbECq+CB3Fjpb5eBerlj2efUT/pNjAUtjeXuNrpg
DIqk3jU92rDFyqNU75gh7/PnavJzByG/iFsCrCqMzMsfod9S6qd/lHIQ4rR9WIjj
Jra3Z3wHfQYf4+LFAfp2u928v7inwWhnUyR+DxBKd3dN4AJ2TUeKVRQN+DWE5T8k
wUv0DQfaqOS1TDHcdmMfxfy6VCDocwb2oUAVSD1MpISDAyNiKGAlvme9r3coCT3x
O+NxuOr06DVl/TyuFokio+zmUOLKugtfQIZBl8oPZHniNcoum04oGe9qtEJTihsr
R8erSKjwyDdjukroNfxOIW4v7+vpHvvKhpex02+RCL/tDYZ4Yd3K5XzSa9a+SZ57
8MLHLKt8z2EDgKMALeFnIK9ImK2Ujzlx/13BM0hRnMx2iqNawZBYKji+Brmcabpu
D5/bxNHZU0T3LYssvpTZ1yOhQ722jo2B/z/hngFEspin0aSjlUInShYATNFEhBz2
/Y93LNzxCtqGrb5I+AkwdFx6vM01y3yySyri8wPqpY2/UPPNrC5XwVY3B8Pno6js
of2D5msRlKmgR0NIzCC3bB9RMEimJpjEAMSMkZDA4G5a2wEOxw2uOZ+D83mCTfJB
xEGu7n7JDeHWRPjTFueUmQZM726LSa0ntg5+I4XyxtONJ+GaUsZ/p8iYENenbhuh
EEyq4c17UwHY8PuSLj5K7qLm4Vw2RGvs80ZGDwuilmBRM6JeeRCASxTQueipofNt
v56jwuAPR8nRJ2IRE2BvfqQjljAKJeJwaXyRWlchlsFaruas3x2kvFAjQ5HDod69
xE62sdd1j6PsAcrMcuFuSw1ucM4lxTuRuyfGjVJY/yYjpJiJIm+rF5s28117SFOm
qe6SupN66cVSKJdMYs+qgrm4WaDPZli6g4igghLKm3sjm4/oANgDvViaH+ObLD5M
R7figyOEd/TyziDCfUXBbYiAdZaH5b4Cu/+FNKQ4DkL7fxnpz/nVIcC/iObd7wGi
fmNaX7AJ1EQP7Tc+gl9/1PDCX7MwPSm5sDJVvquj82e6QuTiPXMVx/PRNlazlHsV
CulMBvZWOBlhAK/GULzQ3gYLlzn2LBkzBNZne9F3JnVL4eHdrHa1Kb+ZScU2v1UK
AX3pU5L265eQlp5sZVKaV0XSN13SJqrh0oWrugRjjR04ddxfUR6jM0Ysr/FA5Uq+
hEl5DVDEjr72yckEKNAfVjFdUWeM2zIZY5VaVYcYAsvmUJOUX9iFDkH9VCH5IgRv
mOSLPl1YJt7hBspazqCZwjx4wAs41UfCVuxLf2o+abs9TzM33gB2GpKePf4DIwkN
q3cJRhp35Wgzxwk9bEC8LeS7xFo8ATZ6rueXwOrnXZdxPc+aZolYOKCKSsgLONgD
b/dPikHIVDgNM6Qq6WBpQBi4oqZ+BK3Qr2s2eoFLtnJHlR5EKdgPAC8lMNwCndOz
Vhzuc2DP+moPmmSPMX4AKJDsC1gVsfjFz9GGTibinO398rzxAAeRK6bcWwasl51j
lwioojtb5eyAmb4jSGELZs69PW26AwCDoOtryRSUcqGMJZsfiJ5lOgL/o522PD/P
t8nWhEC3LPsZZOBanbsw0OK8IpxIWUMq6i1eCK/kVoB9yH8TvONLDXZ2kn0JX4MG
/xXUMBiBWeS+R1EgUGsGA5Y16frsWs36miGuGjrFgSG3udLoyAMgVKGn28B088d/
gjtV0aA1bVhalvFAf0sPxgGbsALUo4fdPl4a2iuhYWgBc9o8yRQr7BNAY5uBDb3O
SKemN44ykMNKoMQGoy9U5KZJy3yhM5SbVCVIY3yJF8JkqL+4aIcGAo5V/bUCOcmh
n1Bbs04gG33dNteA73RTmqTJWxSrThj8H4aM0Gd1ncUzgIOB8EuAU/Kz3H60YXQO
SyHUwZsaYO5gPgLgK6AF2DstepQSm52QoW+VMMcqb8CH2IgGI6/G4Ma8ZVS04isH
V3Z6VZNHrF5Kgs6PMWj2OmKP886Xf8qsM1R5eLHIt6wyJMNJ5UvpFYiMwTOyZTba
hyQKmhEntJPhcentk3PLdeLGV5aU+3MC9mHhfe1fxinWSp9htXSY97YjxV9Tssk9
dWYH6KiVO27yY0ZTC9iRGl1bDlOrqrHU1FZE75LJya7zupaxISBcRUYaPb2q1Z/3
TYvkX1j7VSkzewz7bSQCHNrD1zeFD5cPWun9rkM8OcrH7FkRnF2QOuqYVC+iliND
uCLtjcaRreiZkCw8U2z154V5Bn7lZOTd0BPoxZyZrxYwvrbbqI5UL7xp4xlfHPNP
eHrA/GlFfc87VfPj1enKFjagBb01lT3VfVJfrJmQjlOy2JyAcoTt0GKVBh/elz/E
b/SK/nu+djap8gomjSFucs2HC90g6kaFFQ45bE3I9Qgp9eVqVdeaTE0r0ps+3Jki
Cu3No9nl1pEpyTNL6JDzQ6sRF+bKLs6j9ALuJXW7QzNMfvNf6VNFRhnak7IJmpvN
2zoGyqlEgxZ3PJv9mJxE28r8pkPB8eDRVhMU7Qu5amZiXTp/cHKzGDprqB8bTNIP
jyhvkOaQoy67wCbuJZ8yHZh0NFlaMT1K2gaM/Avm6Hj8deZ+UDuUh68MZMUD/b9A
bzEIaSOx6fvUO+WwKt25YgY5xfOslRIblPZ5YSdAgmnSA9KFB94xMszRi6wMvaNh
K4elNqC3CF0MOM4qiKfN+ZSYN1kxUuaFJtFW9OvRT/tzrASaJb4yh3kgTgYcJK7r
vp22GqjVl+kvNp1bLzan+6jK6+u/nyawom/pOkalqhall35iHKcXBFaZ29kiMe1V
Oamdxdhxl5Ve8utv1aJ2n269CxPbDELUV6wUpnLndBA+I24IJOMa3+pqpxiaRt6r
qy6osw7kHG0ZAafIHB4TIs6dgw1AgxLpBDNarRxDJPkflDaNae8NarKwHM3AjVnc
ZBGZyh6IRXUkogHoNXgADT8RaoomYfOdIP5Q8l3ch4smZBqoCjqyJ5qUo5foRYFA
1gv9YaMT2RC9zT2AsT8aX+SfYgr5l01rMGSz4NUNHgmdEWYfg+5oqtw7kP+9QRq6
WtSTYseFcKzQngH2p4DGL1fIAjDfE6zY9JMRUYri8sI68cvfhvKfpxWrZDtwUV8p
V7JyEMaCj2usuoBvWKAYR4D1a/arCEisj/kmdHBNALuxtARZHYBWntRJh4dR8QGj
IZasQrnwJPd387R3UPAZq2XX3TUQL2L/NFX0Mahq8HZ1u28Ec2aCITco273/dUw2
V3f9Dpjm7QVwH2fKR8DLmTCYVphdIrw48GGV+YWnaY/eU9UR4DaouzUGma+fElQ1
6qvCOPbtSURX/IOFQZjiVHvBXcmZRPN6AS9+Gank+d7fkLIyZAy0W8Pe6MsOfVQQ
fwNV9EFyOUzzgNYe24gACZi7r5Juya6bcHCJNGCEE/GIF+1Lh1+onqYFHaRSgRSr
ix/d4ZpKVA9XDCbXV7Jb7Hy16fX2SKaPL6iPLPx3HdFsNclaXJlltgJ4oOx5y3LL
L6E87V23c6uGV34HUR/N+JV9bR/R8khiB0rujGHzOjDWujn37XFcg9YpkGLb4KyQ
ovP5x2r4FATEZzuyNcTY5RIELX9wKz2TwsbZRuKwiarA1e0niqeWxgC6q82WAQr4
qxnfhHAE2UyYZnj58AJsOJ1YRBwborKgANiAQR29bym/Txczsf8Dcfc/Nj7FygYw
q2StnrPDO68stT4iF62J/uamLNJGK3UCQzobO6fO5BQCHK9H3R8QdEkkefwvyHQ4
TmazqbZePcQcnrsJkTQySTlXxuN7tTgkdp8XmhogiXMFPAJPVqcO+dMyk02rsqAP
OjXYUdcp1Pe7fAN6cvCroJ1tVrkGqlstxt2nxBO+1Mq/0CnI23XfTaWSKneKeKb6
PSWuRhDwvhiU1bvWjonyGClIj0mdu6y128kCcwOq0VSANUdwXQg+3x8xJZvP5N8t
1KqwwSvl+SkX4lEHyX9GVrIqQX0uZmyriOwSEOt/Jv7orcc4O3lW8DQaaDOcRAUh
e3qPlioSqpaZ2F+/Nu0GqZv4d3IGg5+E4TdoRGNB3irU5mZ8bVEQHOngKbQY2/WC
JlKAnQygwXNEJLFzi2PxGtE3JdQyMpPHxlQ+Z5CQLmN/XUHtIeSiYrsIom7NW2Ea
W3WjBj3uJCMhrM5nSv4DFCGCTv7pFT9K7NeOS/0x8OqwB8jdraD0qtUc+dzg1zYu
olHQqUt38re1+hDxsJqR1Bcai8xIP+OKS6GDtnfWgPgOOUvKSp743zPCNUrPGLQE
uV6gfDeudTURAiOiO1b35CbdQdaCQvoBtnZvB/Ihxle0Z6W00J4rN+59Nd0rPkH7
b433lP264o5L1WHOzfmC65JFBnOOs4kRbHT5rvOJcMnmomSjsYvfqIyEcdTdoyXm
lPwSFk+XZQDgvAuPajlzD4s1iB2pmWR8yaXA9GbfElr0eIrLWCnE24PQ67bp02W9
xXZFzx/HTBvlNnTgVlc8cOcmNL9TEghZg1oVaoiv/gRbHe7v23hZ6TuR2BPLo76L
F8jzrHccUvU6saKeqKwa1saCDX/ITX0EMdF3dv4qipBsqd/E7rgeBp82dey+rLdt
BZOS8wfCnH4fL2s+Bu2XNtWY3xLCbky1Dkp7jKegwKthxfI/etTbPiClrW+0jWwP
2Ig3LxzUo7i421e3k7WMkdxTPU0Cm/3MbK2YVTU/e0Xh9TaSIuiLOdjuNduipa1s
1Y0+a1mh17ls7cU4IkmJnqHdpZ92AM332hNoGbg4lxtdqxtiHWAPgcpZWE7jsbQu
VcsgCfPUrwCuZknQWfHhUL+ZUJlZPO+KQJhleI0bOZBZGRbIKmHSvekXccjjrfFw
FXIKfGezTcDl8BowE1qIW0zEEoFv92QYMjoykVOXYEQVi1IPj9OsXDh8rsMVclPv
fXF+MHtTU+VztsjRm3krB31Tqs6C5ov6zCbRuWLch5zaVQObTMfNjx2Z80DZxVsl
X1MkosG5Bt687E/0NF8DDFvU3Ov6sf+0d5g8fHUz7ON37EagiXpKGE170wvzV8k3
y+367m8h4WWpzo9Gk3XMr0T3a2gvDJCp22n0XuX9gOwrC9HW7QsLOLMjPv7P4p9t
SeIRSZu+WXSbuSoqPMCow/WlH6ZiX/gQYxnym0yi3a+IxVjqAtEtuQwt94sQagI2
N8PuUDNcSxklqtIgOiT0CZPXPMvcDn93FV42wTDeAE0aP2ebnfrI8GWe86tM23yW
6WoXCyPzqmWGT+mF7apsJw5fFYgt//rvOr3WoAJ6X2LD89j4ZJxHhd65DMWmrdxt
MOWEQdvqNHEfj7JnIqlfuyc6lGe50JQufirhXOEP0F2xWtmHm/Dd69x0svJA8yQm
uiESoLHyVwKVpIc6J7/M59zcrzkDDL+xL8jJ8cUIcMoSuYuj9aUTbBgWgKJriVye
yUyzzL9F/W3bvrVa1BZyhiANT5i2lZDE/iSmCHq3Gl+5HjmKtHIMIMXwtmsubflp
7trlms3AkRdoTg53UGcjonHEAqm4UW7fqZeywd5a7kaCgFxRVrF6OzfeyqOKoq3e
GEtHrh+fUpdtWNLibHfB66lbVggzE+8e6ZhRNFF1ZFQqrExv8rMNW0YeogxvaMXi
0Me2loDZRgj7X+DycUKBvqA0zkFFXw4k7IwXi4HA6CWJHABX3RpDhsl16OAiQl4R
AA2YEa1BvAae3O2iypx95GMIY+sfphH96z3ACWqRrry324gmqNvAmMGXuewBoeHJ
oE5WXphIWcGN5sHBrNnf8y2LVncLbEuCdqkt3I962NnO+vsPLfLGB/TlMeeAvT7M
Hw542/UWVwuSnQa1dh8HSsXxqd5Bxh6E78IM9penmk6NCHRbnFQipK8miW7vaVFR
6VjHMAC17967oly7mjhtIi+YpMKqx1LjoofuvJtjqaIB863szcASLkprxSPzTx+M
yQBbSo/ZmrXdatoxnDqkXvZSTweY8BklkjEAbRdTSvhCP6cRCto26xfu6zZ8QOaL
cobWSM7VaPAS0xPcsZ6xZnbEPBoxqkG0oDl4MAgZu2ZicvZC057PET8wvmLyu6k5
8qQxxNvjxYxELx2DterRroRzXJZ1tbvXXzmaadvDB9zFmDOf2XWj8YKd/SwlZ1OI
i7q33j1fOMU/ex7vjg1P6w1yL8EP1+IX1MAnV9SO+BL+/p3a2dxDDMeonzLTHz22
EUERQ2g73xNlLIpMOtUa+Kn1HAfk1IHr7RtociihTMwJRcRfhJV4mgbNPbqGnyFS
d+Iiqg0OoPEe6eA+n9jg3la55d9W+9e8Sucuq8BHtYXAwt56l1+5fQD8x10zPv/T
ozJT8v5yciahPYU9HP80iJ9no/JhgzlX042t2kmVh86Ls9YnYnqK5iNEM/Dn/Zlb
cEXI79enw8kLzL0icf+pXbwLooHNgQmoAMvu14cPd3hG3HV146lgtFF+BVdnTo8P
3mkHBbI7VFM6Dr23yORhvPrjC07FFFsH0xtwehoCgz1DIBhBHjkvFpE9RP9NdYoR
wMEclAQqQAKsBE37yJ1EHTZqxPuVqobltoon994qD1V833pRNCpuWB2dJEoPldxf
tvopelmgmR2DnsWlQvvekC8BeE+EEatRitBaIZUSR3XPlhx0n0fu+hhYhizF1Rmi
YUoqSk5uJeSLS5tl1TgsLsdYNK1mvkNdgBoJ0lDyrS0T5lnTuRbPVKroRf4fwqOj
Lhug8rltW/7OfRsZHY0RCZhI88NOPT78J6PEjWLEJ3rNaa623nA5/CX0LdS+VArK
83TrYRp1bQFU9XabTh20+h7QB8b9bNTYR1IPjf95chvFsEPu7tXx4QJoH3072llT
zayX2CwR87QdUlPwCA0Gi0/WaWLylGWlIw+zVUAd7TcAr/iDhoH0dPdJEy4VBPbM
pnBYG92GJv8HiA/xm4ASbu0g16aUx+Fxzp6IxUgCJynDLNnQvPxRtf84aOwXcty4
B0fP0+6pVbt2WOh6XOklAMvKvh5mZrj9lFBZhuKHjBV82tt7KTZQmL9GyLu/DSuk
wavEUz2W14jNIUgOLc1b0SSw2f0qekn07JhjpdrEQT0ZDnvvd4dv/ipHCIvFFcLq
pa2lFhhsO7QRfz8HPDz/XUhW6uzE4f3MmxOI5J9VAbCspW3AeKvWwiLCEhnfKe82
+4jLNZ1OjS2gv0qP9E01oorU9ztTk7BcyI4XpP5oCYZyNg1BDq/IowrojI91VhhF
SwN54nMvlR6zUx6A6j69wk4DcZ5t+HDWnh4vrJ0tX1GAh7mrlYeR5zzBL/LOT6Hd
CVEJu4GeusgtqE5qlu7BHHEuwnhcRma+awMQg0eq+uG4K8RgGZY3+gyM0OqVPQgI
ulAwVTCXvf91GMtFvMFsE/7vOP7FXlE32Pg5IThfUMAmzegA6GuEW2Fm4fdLHoYh
BfVa0T8Cit/x1oupmGZiCEpcvEGvB4ZrKEF+xZ7TsIjwS84rv+3gahL1Cq8aTIMa
yAl/xvJ8BdyQQJwq3+ap+TXUrLvlVj6O3djY+hUCgVv176meU14bzM+HIv8hcDxt
bP29tAml9Meocp7L4CsS9v2O0a40JYEi8AdJl828kPsIMKfVF2fpQ2j7kWjI6ywJ
6edebSz128s4AHbcMEpY9ZzCkWPxXg17NN69MyMtZHmyVN1UxISi4a7vkQAmGn//
bYAG8rE/qSZNtzqREtkLr9MMUIA2Ub+LCeLrLP8cvrIkaOQWy51UJFIVrYpfMKKs
XJBTmz5fyTamISEqCvwoqtZGaU/5IHsNsmehZ+aKCOIbrpyNQveSTg2l8Yc82V5d
C30rLFwBoK/x5uuc3Uzay04siknY57GoiIyYQS23Z4lvdwVVIOqwHrqIkv32ki7R
fgabFbpylQNx1NnsWDGauCL1Aji1e5rRgDFd2JZsIVwJjkUsEqrzbihPtGjfXRx4
JrfYOpVbDf5h4j3AKCF4o1qYiT8SDrMRj95oXwtSsGI0vu9ZQSXCPE0l4XjwKWcT
hg6WM8X2KJVg7Xp7w3CfGCWDSTpbe5mZzvn7wQ9R7i7wc4EBt/KJ02jWX49VsXG+
wP8G7MTXom1MxMTeOpbOw1Q4QAAT6PwUlathiGWH+BDorKBlSWiIdy3VW0dbxapb
QYnyulxSeoY3FAAznEHqdXIlQdolmM227s+hlKixkQWzs7VPkY1EHt3xpLX5XfM3
GlGJING/2GywQT47jp9bEMmLeggUBCfEsUIbZ8z1mOAlOZTpvVr9/5V9k8l09cjZ
4H2GOnuEQJUyCGi6Zl9PrTDC82bHWeRHzhrxHf2JSKOsqpF8WuO0JeIQ1msK7yHy
yhcM1ebo+RgqXo132Do29OFYwazdn8v0y/WfmHNB5MRcA/bvjfLTB25dEtL22gK5
CKtzjEzZmzMjFiAPVpSizd8h+3Rv887sCpYj8xBma1f1r/nPtaBh3bzRjacY7CdN
f8FXkeFTKOGRaZMcQ7q9zy6wwAtp125icPHzvO3aPtHfIESIbygZZ4QzD0y+HF9y
IRAXiJiUmoApWnGJ+KW8gsDWtm5ITU+ukjRoNtByWmgAhKrJ1LoFZAt6ZhhsrU04
Ob2MTHwzRjPFvBjrPB29Su9ksQyoqI4u6ToQO3qntqvH0kygOqUb9gki2Fm3RmBV
i3psUELbxvyDezOF2SXvfyh8A7ak8HFcGaXCdApNl5cLvqaZeY1Rx9OOHbEAELT0
1WYTtZZ4/bmlIPX0F/yoAz02LR6DpTiqdYInXO/E/nFpy8nFcaWi7YDVqkU4xaVO
ArhrpW8OwierYQrA09DnK9TSl77viUtI8PTZtLEEADKJIHPeY7mwIBf4hM2O0Cfq
o7XbB2olHChxGGaxlirR2Hf2Owt+j2FKTmKM8YQ4+vAvuCkucGGfVrr830ByytlN
+fS0cL4tqcH8WMpgrHU6pwxzXf0tonEqorM5+OPKFFwdYB1ppUW6XkvNJrI75Q+l
T92lZL/bJ1/ETII/i7jN0FMkP/fL4jZ9efbR1ZaIpvkIA4OZy9HInKV2DOTuilEX
EjcnttqyKuYTFtBaxvCx09EdppAVuGysFv5rqDspr/rvrxRoDAst9L06M0jNRTU2
OjwSXEYKfgdNjU1/f5DnNoBZDthUc8UiBKmnvkpBSoVtuQmK4/hE9iKgSw7Rg98S
3Us/mR5hMm/7cggLo/69KssRBzoAb8Zu7fUNZEfqYqjILKNwiDmfS7CR6NhLJSN/
ooGBPmCsWUKEqofx8ejgvsrv0NT20fkeHtNMN4KdlYanIZu0i68Mxc7tMoD3Uxt9
dAb0lohC8l+/aqASw2bQB95fgH+L7rIdZsfr1fY9T5mCWvH+YfRYQ9NzbDQLR5II
e+93NnKCwmSR03TgD/UDNU4ae4GFfXnWQtd7CVGedeFtFK8vD3wMJEbZvLc6OlOa
YIfL6curDP1tHa5Nr2LCnQwQBzYz1lZrvEpQUw1B/ZKtLLEpuG+yOnShvhMMWVcI
0PIrDZzoksV1gEtqNsX+sKlQWi2P8jS2F4BNqtdzSJ+qkTb6gp2dV6YNvqiW384w
XFllvsbGCbrSHQerG4396YSTosdi/6OaFuc9VEPvJRw7oMi3Ee6HqRvXSlh1e2jf
qZ68LCdDzSWrGWRR07dME9NGOY14bOTuwmJUm4PtJ/jMaoca7SGyXdazNoyhrjSZ
yyO5I89cbOlRYYUtmppwsV5/llOdmwMaDe4My6DkL9OlkD/vDUYJeZxHwuNQm1S2
epi8heUufCo3cU1asNwEd4a2qqK8VkjxcC/Tr2pjyKhjwheIoDcMMVWGAS7VAODg
RQdvUNV2fN7ASSVzt5WpugCxRrh/+TdR1vwk8eCmpG5m6RHRZXoYoxVYbOpQgN+m
b4+7Js8YbHSi+DqYPeJfGjv2ynA/Wd+B2soxI/ITO4+drajxjboTgGoigvPpX7F0
fxpRlKG7iDZl0EKl7C77qPQpQzLv7zR3ePQYVXdiKSN6sR4TGMFZfa7uHlEAtwhZ
ZuihQHGUq3sJbqt8uzdphG7uY901ZK7jrXnFzhwqZaG2UPNUGqMzfUYVpy+B4Tl5
7ZS21E5eLAN4RpsznfkOYCnps/a+iVhkKBiKXaNkNf3dczWPLev/0kQiMV04GuWj
9LZxgW4KwehHirkmLtMAwgIZw9dq/VC0OL+maFmAVXocJH3c7e4vZlVvRoAanH3v
Hb/HWmSJdQQNRNcAeBwukcd5mTNhd0k2sjR79ceyqBbrfnkcgzVDjLfSHlg44+xd
al7EcZOxYC+HdJcl6SAd1WhPnPPOf5ebuvPOdBeyXHPl/Js4Jes43FQR/ESyP3cu
uIWv4Qk7f4p0OIY5IRr8qG/3IYmldc8X3XjRRrSKZt/vBxZSRel8K/MPIrBj+cNP
18tXmK4wxTl/H3cWjl9d5srlf9ZWJ+aAAsqtGqCJseR40+eD6O0ybginRF43CQP6
P2bARWqMI2d+sKUWea9LQ1AeIOHRly/sB4fHrHZlvKzj2JVzsu4LeouyEo8/gH6N
GTgcF1nKrg0R5+Qj01SxqkzsDoutQySI4FqiIQcYaj3eDm3JLuimCovrkXgRz/+h
Vv92P/NhzaUx+T4F+L2jdr0DbQsrF8m+kAnY1n8DsGndvsJGS9O3THpv/pxi9xBT
hiPfqd0CHiVOtGGNwi6OqAR/BMvAVNBG12Ah/p0QWSWglFn+/WwJHWvRSA57Uudq
RUdbIHBg+jtE2TSf8zSCFGYbrZjpl4PVntoKG9bGXjvabntar+x8N2c8shKH5ajc
yVod7vt3QAECfDX77m+7iTyDlysS2nLVKppMynG1sVGf8TLOAS62UJDMevOMSN5c
HVtxMm6iv74j8eRnq2EWr28GLZXpcT7wOa2HQV9mTFPpdUlkPKPqDzGC38bALj8G
OBfHvoTDSnnf4SdqeNC9HrwLA7t8+1bVQLg8VRtkR0DjgHwS0JbobOjoGswkqpJZ
iHpZb9JzHth2pJCe45Jm7UxWJkWizJvswzNbLQQR2ARZ2Te4i45IipKY6NkYvQYz
yxuFhU7fuavwrUWZJVWYeRVT6quWEmunZxOjDPwbsZ6r5pnMczls6roYEGhHorR+
qFeh4vgcdn2ZLT7dyza/NnAjs54TaK75TCE/2Qnf+NOUASpThUl6MnL1QyGr0awK
tULt+jn24oDFR8wLJpDAB1x8cF0xZvyAiuF9J56Cs1R21PAqs/3EEBV+N0LN7tCL
ECXdu78UgFmbiUkBeVfkrdZj3mRHk+9eYEO4ZHIEslo7jWR9aLxzCMRbaBHXNGfM
2zOTtiWPgKmnFBkb9QW3RbTrgKHcm8bTlRf8dCMYkyHzlqEoytDYwzQcZs7lxwuP
hx3lE/pftc5dQFIwEyKLObQbzE/9BuaKqHHEmiOItRr1g8P9XIgKIRIwxkXuWhPK
rolc1C9NYxVXhx7H2pURX4F9QVeH/o4L1KtmNfv/n2qX6P1nqUjYGo8Qwto4TwNg
NGzF1eo253gW10t8rQcfgNHeiR7DNp7nJArUOte31OB/v9qNu8Fnj1RUwqHLwfjJ
F1S/O6eVcJV5GHTveroPMAMjLKDFXZr35XyZiphSMVH5Pi7W/WHDX6C5U0yzSZvO
q2drVWElBjIeSL7HZDrHtgrOWPMSHVEN0hOz+wbnyIQzeN2T5wZiWam3dNL02RlZ
lCw6EbcHiBT/4IK/aV9iCV6GKLu8JdUszDjx5DhUY34/dWkuUUo84T/r5AbN1xnZ
gvZLFMCd5vBSQWD1z8AqpHZAKv/WZIR7qJwtXtWOGtdbE8mRtOSAP0RfdjU0zBdS
D9QRY6I/Wdf4zj2gyQGOTYYQr8ms7SSAFZ8dRGcaXA/CRldPyg2xN4mP+S+1TwV/
gh7OBpkvwY5dg696Id3SzKEyGFB49WQyc524nRtf4NWZnjfEi+rWXAFBdoiIlx7W
r0ODx1LSiHwlkzkjbYN3ImnmdP/8vQkq7hgvP2zVkhbga+5DdcfYHA4XZEVjwlzw
qtXAVJ7rDtuutnhYBU89m1x1r4bKJRE9ecFcoN8hcoL1I9MRCjZzL8A4RWW3737p
i6cGijaCmZQPzXUzcKWwCZxMv5U6OU124f4PkCDg+zrOyI/sLNhjjm7egT3xq2SA
pI2YEMsrr4lk1Fj1k+Vjz/vXadijN89LyTgXpwW34cDFzSh+cIKSZQfDmV0wARqv
dyFiB7RyD7qmLlf8VO/zlHsbmNaFq4aQHf9yH0JbcocDCiBKmXf0Sll78kZeAIBh
sqgXFOoBB9EGBs2m3XN1cPW2ObftqIwsKv9F7fXXmTevzBkI9/8yQw2J6pYh76kD
wY2SiLE/BNjp6PG/pWj5W45i4p0kbGLid2w1M5J5YyoSSwZOLbfgYoXHTmDhrfLo
flq57KCVFov0OE7SlrtY3gQLtaD9CGwKLvtGqLwS8DdbEwq6RuGaaWulThL6sT5N
QzhD8gXGb4nX9JH1zLouO4R753sE3B7bZ5NWGqKGy5Tu4KkPI9wBJU/9W2kjYegT
V/O9g18sx8P1X/HGGewOaIdHaHN8eSS/Yl3R/7GzHE08RGCQyZCRIa/3dd0dzAo2
ZHzvFdi3OrKy3qFyMSMfgHODZb+3/xrx9XmWzo0PizsVfNbx30BrQZf2YHyNtmr1
Ix+yVDONA0v/zbV/Qhm3TD9/8+Ub6raUlK/knhND2rtEglZItmsMygTEsWQJ/YXo
/w5/TH4QcC8Y2X9Ykejqxabd3e6ed91zJn1XZZHEDlSRZa81EYfZOFQCodCxIYKi
fEfiqeW0msQo55nNqhND5g51CHtxRFkIAxM3uZ8gY8Tf+PSbSW4DxRu62rNDlj9i
52ogerd1siW5+OdQAtthwjOja8T49rY9Pr8QuX6+hLEj2O4sPpx1+hLDq1m6USdK
ggImBQnw7zVKM3l/vL1zn3aeOVkWfcJ/1YWBa9jYFBu/azPNLy+GMxH4to5hNIP6
OmjeZkc0eB7F3ibdslXoVwsIbv1WmxlSjasy7uOJlZ8POJK9wwMIZwsrfYHtCaCf
LtTwnzIy5QVSkz6euU75yl6hvT09cVLT1W9H7OOEdT3X7CeGMlej/aroJ/XclCys
7RVREgSbaI45uEBJ+GPb7oJVejtJcEu9W7Xpc5O5/fROaS6fJeB3NuzxUn7BRd1+
JCJ5dQtTBHW3LFKb3dWsm9CG01uTU5X2NFrZd6fuxP44uA9VZ9rPxORrpNjwyAft
JOPmpYaD0xnclFjrnhfcXi5z+8cht0cwbuW3zCTgoeIa5ORbMFOpiL5o7z/yOhhA
4ayhC8nwQKzUKd99I/3FUeUNxWyNyR3oCZgHOS0qghCGXx1xU2svo0HOAvSrudHo
VG7/T227IcOdHLKRHm7ZgSHusbc0BknLjPr4IVRXnzbko3AiHb8X5RZnVK++4s1L
ejZiBkA1bZRXkaKn0yLL8C/1kIGKXssdk8ZslPT+eCblGgZRJnaPOlNq/efEomHQ
UecnYqEcqg3kRFfhgHAp2T8Xktyu+2hZUkrmmX3/VGKQTBeZ0R4g1R4UI0VFuzgy
hi4KlpFFKTTwajvI8NGv0R21VUxBX5Dp9V+4um+BoP5n6xAnLwl8ui6HHtnRIb9C
T5/KosICZkClPhYtJJdVPDjnW9atmNGZwNuN9Zy/HkMHkRzfl9LHhbYvhAmfahF5
sAX6MWVe6akUyXOBuDxAA+VcGGXMaHKGQgAT/iYrv8wFXQn1KJE9e2lUQa5sdaZq
l7qKolBuJkwD4PSvWA/VVXS71HfIM6kfJpxXuJOwNws9Aq9C/68G1ksuMiIgv8vI
2hDRQbbN6QdVIKLUfFZ3HB5Ai69kW8b05h8F12HBO9zjm/YUXg48nGHClmJBOJ7y
dHnXQjvpFibqS8r48Ky7vC81lIolDMkbO8pRSE37NHf3qzIKF5z5OUXQ7msojoQw
fBV/1pBvqxENiYa+eRX2YVJL/UhgTf4lvjWoXRUhsAAYzMMh/cS21AplKO0tJASE
afXFfxbn+b3fpPtW58RBEQnOJxOQ+QvjNerqumeOlNglCUknYx9yR818c6//LWDW
5PxV1DJe1TwZWMQ/2BsYoU3lcySkGdHkUxVK+u5np1Hblf0VvKJsgMjAa6YLZ/1k
FgNvHAl3HLmDAJSHDsZB4gdpaF69FZUwW5IiyYGH5uj/yVQMlrwQTYstiWhEfxj4
jACVjx9vOFYK28Yh3tevgmKbALaqonCJSPQjR1NnMUTG2YAbxIIZiC2csRu9VTUp
Eu5A48Ji4ehmpIp/iyF/eCJnmvdlS66Zl2xDwgpJTGuDHpobCL7VaiRDA6P2gGP/
qA0vNodRXvpEGYO6eRk3CjfrDzmdo2aHyJZ2fM9uERg9ZsNGUm8YgxfUlsIgkqzA
dnWQ6jzDiNX3TDZBkHxkHxe90T7RcxxOKUzvNUSUE9RApSxGFzQzV8yG2CxCkK1T
IUkW9zHUFbLigx6O6GHiOpl2UfArEcMS2GfpRtsfa6/17m8NYpnHBuzMF9/1yggH
FweAyQ0wUplBV1RrBbU3l1iaVL168j14k5jZqKJRgspzAOVha+CgxHqJK+irZsH5
NDR01hfMUukVqlwlIrSRli+6v2zh7+JSnDwLLz32vUolNXIrNN0eR+cHxbCFOP9T
pddIWYdLEBEGJfG4taa01ArKdOZdJGIrnWIDXGNRyYVM6mJJyZOieByxW4lLezRf
qDvlI6j/llrsN7jZz2KGBdGsW/Oa2ep9KhkxEcPZKzPbORmitfBL0Ynwu5MgvG3M
d5UrL8uUV1IiNldUkg8taqWqtbDCo1w7P4NDhWrLVQD3033FBQDiwS2C+ZiH4wQj
YNnQxVKw7LdJ+p+j7edm+1TDuBPSIfxRWljZSQatxvXj8G2qpN2l+aAfZ9wd91jM
Gego67rk0uQj5PY5XdfW0VJ4agh8FdcmOvP5Kq+2ZXjntzVU8zc4yVaJ0TbYz7hc
4j6fOLnY6ZXcHKVxf7n2b4RGW6DmIGt3dNSXsu0w9djlJyI8ZBWLOfzA2M/5j4CG
lputq2F9yUvPT9r2gGCNJoAafia2KfeGu/ARcvyobKboz+fPJW2ofB5VtOzvzVwL
2DxRZ7oL7qxIoEXvYYmyDHCxXPVjaTRNeMPgd+/+V+Bq1q5M1FwU3Dc+Kin0hRFy
AU4UrYPXguwOQLkIyj80pEb1k8bQ2Pp7zW/DawQW4EOh9y5Fwkj9EfzE0Fq9iSmk
1iEVQaVMuDyxeB6VQeeLQ879NNBEe1/y343b6VQDOn3UgpnFTt84GTfSJH/DxZ+/
+E64wHKvFKZSOjNUs2q20TZq91NwuO4CYvCHNocUTK79n9Hhl20Y5uUuRAFSP8rq
B1K6Q4XlWhQVWzaC7TnTK5SBdZ0m1C98f8ynpUoZhVvegFdbDNQjELzj8mCaPj8/
VlMPOKFNTiRt5WjRkH8Ri+BftgxeXgbqP6Frv+5bt4JCzllxH0Khut29MWQlgQmr
lyyYG3aYvDT6URyan7jWoy47yakUSKLtGz68OjatzMOG2bHK42HnMCOEgSw/wujU
k03itdAlbtsy/71m265TiCfVvu8nVb7G9eIM1rp+7kTLfvLSY66e38GPvfQ5m4fl
syA7J/V2no/YTLWgy+/UIo7vHvYC/YP/VxabkVjdyhgI+i079LPLJwQA1FS/sbvi
So00U4mKM+tMHck/LWy0Oqoe59kKjphXxsqCRmuQCaZbsjHdPpqEKkRIQxhK3mkh
wvVZ26Z++a3MIKtEF2ONaCl69xrYqd90UlW0PQ1jUypMZ4UVZQwmPQObLhVY9sh1
0N5ZCkt+xK1WQO+RyojTrblTfwVGn3GQRbcQD9bwmMbiyC/dAxh87AYjVD25D2MX
RBoYqa/V+9WwFQrPWGqHbDrhXW1WqR4kz+zaHiyBW83JiWG8futcBMxs18UuGXIj
96yua1lSUlMT8ayA7Wd/4Tjcz4LVJA7BPYXa3lsIzwxRh++dDO0qtqL0ah3FX+uk
GVFaojfFPQA7cAMyXfoIp1686m8d1hsKLkkCn3U93cUAb+5Wh1YFsnGKtgucQw/8
FNDTo0ierl4pBAQqb7CWdURZPZWpdLQXfDZ+oKmHoALoaYkifH9Iq+kCI1/U/Wzv
AJ/fW5O+kWQ3YepLBwRDuliRul2QZBzn0izf4Ij7b+JoATI/G6YLUvN45MJvjUG8
5p1kh5GQZEmOhYF2Lk4MAnXk6hRUCZKuV1ZDsQhDObttsgfeq2kIJG/u5mrh4RS4
B/u1w/3RN3bTsYwTIAPLCRi5/ILt0PbxUXjAyVKirup9snkdhk7jpi+QRfymHzTY
+yD80BPbHIwUSqVwe8UUkWQ3yRQHislfm9ugqkPUyVqPlFn15TKqPD4Ba5jp4oJq
FeVIhtIrnoZEbVk+7q8w79MHSvojrejdCwJbtM70xcBzxkY9gh2ntfCsnga3e3o0
lPa9ITsyVQv8dhOf5sMH8OBDvC55B6c82GYmKTJIs99SVgjvQ069PVrRe8cY1dSW
A2js4T6kdvw06KZqHEC51c/cJHFLx6qoSS95HORZMo6QVVtLkGjRHx4W+it+YZXE
8GCsIK4phBWcy+I28hs0lq0Z+ccPyOutgzUmqORQ+dbtAqOkWBzsLVGpBvwKYH2U
ha1JBq6tqhimVOThT9njI1lY8u7jZsru87C6AJjxQxX8XYkglw2ZrsKm9TyO6/6p
XCTw1GCCZmLQkf0rcsik1xkXPAo+haHCNpj9O+SCtN05+RhSQgDXbhjr1Rv27Ar4
/62TebjB5GtySjZTFZ2m7GYFCR5I+JyMawgePA76G254t8VzW57SWK9IDzAO8tWV
9JKoNFINrAtBzxlUxZeF4y5FTYEMMDYmx/3ugtHk2RunCOWecdPHn51jhn2tiX33
12EAFMweiXtVn0a3SSEUa39MaPqLFtMQ9x1AYYwsRlN6Wo4ETJIuhm98tLpxwYuW
xVvqXvreNfo3RopfWY74W89qPTOVmFps3M4J4QMRgUDUKZeQvFcmdU3mGDpFyBZA
eB7bzCQRQmvlsWaseYFAPvyt9QhvcvkKapJJJHYR47EvBTkWdQN0y1DV+rauqmE7
29gIkyOPqaoFKctN59nbvjSduXWcvxUlDkhB++Bcf1Z3OHXpVeHE+9A84MgV7LI3
3g5LCjdgro/2x+iTs5FgMvrtI9dAek2pVQq8Ch1AB5vRYBxPkSp417FHAAE6jS12
LYQ8LL9T76Ef0kFs4H2PubH+BKbZpsMzJKGA4g/senBdL9lsHvOlBfT/I/OI3KzO
c60ztCakcwvXofIlH147uT+11Son8GJhz0tMTsb+9lqoRDNJgFZ91qDhzC4trZE2
MBRB5YxZRhqM49dwCXRc/ueVj8XLCGCRwIlrG3WQkOr3js69N1zXv7jC4Bh75Jkf
so2cirzABlaXzi4RNOSxooRyYQo75gR8y10VTLDlIXCfCN5QTdMCq3BZYwdgi0TE
Ry0bdzN5vL13xnReTTA+PKHdanIkWbRZTGZ7n3OFtWoZgvkxfy85Gbx7zRaojMPt
D/7BIiMKexBHCm8Hvgum1fC/EDma751SXiMpGlVsYDgdPDb6A6LNK5B1+yfsPg2+
nPMPxh9ub6Kd/13NcFZdEqsTdJD8qwQ1nPa41MeG49MPxii6yoAPjYJLOspwbnAT
HWPX20wE0blj+jIlzbPK5/CydjyjiC3vB2ZUaiq4GBTyI2k7fhksXtlWPFjgetru
+1bvH2ZHtK8PBrOkcN17hbcHNykIvBvJcJxWiLRobjJJa1fzwwG5in1YwbLwrtNU
BqtMpwhslP35dXB1QY7MoRGJspyI5bXxNzRnMO5ZJIXhyTIreRBhSur/ofo+op6P
ajV6LQhIQN3cGGR5fSCvwg7MdyJclF9ZOWvvCD/oQJkn6ZZR1j2qgS3y4a+8jc2t
Tu2r98kJPtrr0qoKlJD2te4vVGr3GciF3mbwBoGqtTXHE0AlOXEAEZFiAke6Vh8D
eaTmgqpOsoq4J2K9vXjG9/YnEt8/VYBa+VjOpUDlky8RQiiZ41+Wma9+pnHdbnw4
igTAltcP0MUJY4SUzyDjnMImryccw1gUjotuJ1me3EaqQkSw86EuocB+TtnACQ6/
461BBjB5MW5BR74hl7/2/3w4039t6aqEex0RySSHpkyby/5zGc8gbRDMWEI2R8un
GYlcHRtT2z3StgKFbptFMnyLyWdN/bAstVPt6anHyNZHKswZ+zp+27eVnp+h3nP5
DfKeVLfsLcnMdPxOCl2wN/EKx64x80uapYQf5EyRsdozJRwpPcHO6LnTe5E7A8hB
ilg+OZLySFbNvPk5G+K4RrOv7tCN3FCrcgHSYsCD4UrovTdh7AMlaZaFUcijpIXH
Hc3C2OGH1QTVwl7ts8oZOOYNjp5D5WeFxDi+p7dt92vpFb77VS3xH+mGdtsWJPF2
hb1roX3LzF+fDLs0d1hMJ+z0KprgmuI7Q47pMI7sawIWIzBNzuWseHXuFd0erdHd
94vAQoIYUDHNXZDND+/nEZWp0uut4P9sBW6K6SgVFw7PkP+IzLtfBR8Hka4FLRd3
seoS1r9CTSPhsDZyaxv1WpwwIkFgZWDuw30YKZVkPUh0XV62L/z7XicMr092WsH2
XPofno6J4y4BbKOXCIRGxyD6kgQlntfwzJQU0zykb4IGakz1I04skErhVaDGJQbI
uaBJjyJYp1Dfcg137m8sE8spr2UoaadZ0BjIv8ZXfRw0+CaCMVDyZe02zrqhlRx/
m21z96Q4gb7pNqamcEpC3hAHm/rFIub9fgYDuBA4uN6ctpQyMcSBxOXJn3lx6bGy
Eug5Plz0hWKNGVtI8xnudex0vjQSaJOmgZrsvJ03cpAyYiQnoPQjW3m2klFViUfH
t7fi/xnEsxaQkWBvfTKEG82zb+jnnPoI0hMrvDt2afy9nBccgsRf7TADgWsgdVNQ
iEVBD9kdLs5tANblPZo19zLlx8e59tGeE4E8hfk8qtkaQttXJ/pbc/7H0c5XwszU
yqn+c4B3w0W46LIvSMnwe9laqebeEz5BCllXEFtuOZaQz85rtw0JZVzidxKmFf6H
g3XxosHPsMApawfnbVoBBgJ6MTbs9TcMObMZmf7QiEUkIRK0e3O1Mc44iHFSw0GF
HEaM9BABk4cvjqYZmofk9R0mapIt2+mNssKezhnx1yTXy1tVWfUGy95vrEKhqMki
LEgqPYb7jjrWvA4xjNubIU6T6oXJVoHnA6sgQbBxpq6JtphHDOHHPTSCxdH71kUo
vJEVevZWB3XulWYZNTab1eeqTGha1F5KbbJVdBsQR23Q25zH1bmrT51/EpmuW9Kg
THPlsBOmoUI6kFFNjY00Qq/fIAA7iOLsIb4q9aEgWYAbc3sWvBwBN2yr+GfyH06Q
PjBVXBsQ7yvr4VicQIbfGJtLNjoLhvZENhDLcXjZ98LOl7m5M1Pf6ZQojgVbNfzv
4VFU04pxoiiuRWyNB9FQldLCZawlkpxCc+LOiqqqbyVwSqqAnPyVUKALRGpMdaD2
/ZkFc4numUeJJxrzjOe9spPo1RguZ95+rUaqMds206VdpcLvjq5UjIuTRQlrQHFq
FGELu/19LvIe4hILeZU/0uZsmk0Ab21FabAQlViSU/TJ9q2goKtjTaK4rAFYSDH+
zLz+siM9DstqHU/PyJ9gf6f6W06B1Gosm64dkqXMBjnE5xRyOtZ6edDZaZsHsz1n
Kh/NArstpWa6P4zj+4m9XIBNbRHqMuMSviF0IkvquvMSxnmuLfdr6i3tHoIzEA+I
sgncnE8UrhyVoLWofW3q5err0/yxDYdk3gWiuMrf/bpIAeuRW0rgmU36jjL8Jpdp
CFjZri7xISECbR+u/DF71+UTEQm9cnSVLHD4UaTTPqcC+d87FmVRNfvc1Qqzb8dB
zzKtAUWw+jcE7R8ucafVlvJNVSqphOenhTzlUM885VYp8sousZSBvMcFl0IJxZYJ
cEDAn0XgMPIg/oCY79pkoeVa1wiW9LCylbW+awn1O08n2e8H0N8j0PXmSk8uNHjx
51S7Ku/KTDgFI+pohhpy+BN8cjv0O/TDHHG8kaQmlx+ZiPZi6PwOMtzNmgIkzmWp
iZiHtBTvk5Evm6bvcLe7aJ/8GAj2GlrWJEAQbzMN+T0D5Cl8nX2ntBH8HScpe6fK
SjsQtn0iGKTIo1tq+OQeilC2eciDy39BAdL2w1yokV2EmOmm3Psz1Ato+g5pFkgy
jQQxp8IV3MsxdcEwlfWBxHwTR7wO86QeHaqjaT7efAhDyddi+00dOWWMFEQKkUrH
OEdPt4Xy6lcoIAbIT0X3kFUKpkGXbh7rBnLfHJBEd/7kM+TpHTGMPoUE6tXOE9p/
A7cH8LjQpkHPPAMZuPBpsa67T8mfcp+CGOvquFK9WlM5n1jSn/ByxHvdhQRtiWay
6rv/PqKF00GtDJujFaBg3tAOTtENMGP9SzEZhR5c6D5OdekY/1zm3dg0hCuPnNO/
58Unxi+aw3WkAQ+RmKt0QC77bMgFSDnXMY9xUPh4bt9NxMqe/7j0D0ryL7yPGmRp
ZCcK4U/XmT/HjiesUZDAb9XEfMAa6QGD3FgP4a/cUzNd59byacEzmwCUi+lo1sHS
DzBp6tuKPAtIHhxPE4E+iaYqKGBJhI513ryEcxNcrT2r5dtP5zgA4ZEq9PibvtMR
COHUtX9iD181UkDC+3agvnrrdLGCHpCas6U0sxaVjvKzeQQw8Jd1579ajAscYI0v
7bXOPHCnh1RxE0kfmG6WEz6LLdK6ZOwSDdEfq4eUS4he/YbkF7MsW3IQxRzR9PBs
nFetlZGGYpGA+FiuaOB33MOCV57HdQGrugdYylUufqOL0RZYgIG9KRNiHumzA+jP
68BEYTVPiGk76iNd/CfkuTDPWjb18nOWOFcuzoMJqOuwIJzKS56vMGjRsajMgoBm
mf0VB0drqC282YbC64Qhl9K/1nM9CQGVtvhhnP2sBGPE8XrrVCyNPmGSRfNMrdSj
WEDFwAcXdXOT9VCczQu2ih0ifX8vEObvSFIuU//zCzAFzFfUpga8JiTgXx4b9i8x
sVqkL7PV7EzMhLgEwmY0a/zVRxBliPK6XbaS7qyRf4CdNnSxUym4kwBHEuR1ok0F
4Dc4XL9DGmxoa+xJkQ6Z0WRw7u9HyZoOZNnOAugRcZJDdvAT2v4HuuiUR43mo3Ll
nhkNFsUFRrhW3iNL18kVNf/H2v3sh9sypwJOOfMc/FhTaJEMr/G2MoV0uL8VBtd+
T1PBYMebC2KJFHQ+3di9X3LihGgbUrajhdKAvzcjAfH5+eH+WkMxNo0F4RBLz1jM
Mg+93vjpdRX8ltiNiTlObNblgqdrmA+pwSPUmiXe3rQGfV3gSyhIgop62bd8sLoK
ksH/1RbfVOHW2hk/selWgIM/FaPCpitEjRT8i2ZDjm3Qh3p3tzSY8TsevY3kunf1
HWYzEBba1qCgn23YiWRG2Ti0NP80xJ2AmpTm7WMP3/A8/wXuwwp/rKcSDRQrRrMe
mNI4AtoQxXaOZmwAUFUeEHJpva8tU3J46LDK8dYN/t+Vlj5SZR+EkNXBeEBZj7d+
TZV4zrT5OF8OVzfNQXawbEQKBDUk4kWTfSkoNpHxU1UMvZB2HSCDIyzHNRCsbL7E
7hg8xG9iYY/256As3L50MbTjdMN+HpOOliHzqNWj6mR54E1icH3yGpmzJ/6QBZPk
vzypzGy3uNRtM73SS4CuwjJ9CQ/38U9H4h5UWeiQRIP8F5pLSstc1zSU1dIdLDz/
KNtlLF/dNxVPl5mGnmLN2GcJ9SEsNmBBtfzgKADe90mYMJn6VRq7kPzfU+27hD6B
SZf78hpKbJGeifqT5KPjKY2w85LeXRBaeepyFnMgYxbQiY74qPSHQaJAR1BbByQ+
6uHdeOvBFm5Wnm+Yk2wrrgZyMwoER3k2qr6x2k6/BgQBg/HgtQWPH0ZJ/txcD3h+
+/9OYSS8FYSqZCjJ52NoMQKUOB9AB6HC0759fPur9IZnrlWg/z/whDNcotzfbXlg
ppecSULEDrOHaMPI4cTejbUGpyakW5qKsHCR/6Eugt0GRH/CvlEAgmAioTUxWyIR
q9XckacVO+dV7tJmGtOs7wwZjWYlCQSXBqETqIpgHZz/C9YFATNK5BtLmES5icW4
hYb6AduiS2l0P7c/cg0kSNG8OARrEGopjPWAJse5VwV6VDGmBt2/jfHOfZX491j3
63OOYovk8VESZkjhXsCd+dUZv7uRvVydqX+5NtbbMAQCjEnj3ZjZJxPnaqw7vlWN
7gD19RJ/RBZQfUTdlmQOWI2Lwk5KNnESa1EiK75MwHWZL8+8Vonc1NT98YRcJVbR
3Ab8yVe+8OT1YhmHn1NCWLrvLbmruBQb6eXZhLgDJVLO0gcvxQyr3e0pZqElU22O
2fA0Do8lH/IoaF3lpgXG+zd8cuDNN31Vn3efMU7RGAgjNNFGV4lpa6Ll1Nl/XZYq
zxGur6m0WUjj35K7AjGTJFKsI3cNDDtEgUFNfdafjJRoWsfXZhNUMsP9eNp8b6kI
ojgVnWlRxsLZ65UA7ygiyqD/1Efccqdvnuvnq1HZxtKtc9kMX20aF/BqidqH1Rtx
6j4iWDQDs+134WqczZXp7k6hSEJNJS43d6TToaBETuuSmcP84W1U1kuW+VAuJ++K
kaTKd+v2L3k+PYB5WvCgMFEp+l5g07+4Xi6WaA3KVaYeynSVArPldj2LMFGXIRfl
6ENcOPUM/z7L63wkPSUVpreHY/fdbpbix3HOrupIJp09BNxG56qG8iSYd9qr3fKn
F+VR7Afx+DRZhB6IXz2sXll8uNWbGlW8pbIWkE+RRDynLv/XFyPKgiqBO3BID3c3
EoZ4OcYwUhRTd9pWwzDqT+Q+VQN6/S+WHxOexxLLP8exegwqnSbiRR64/lKipmGN
ZaK44rDPUWsWplZsK/uukxLxs9qJ9nr2uy9OdJFGMZZs5LYddg3kPVeVMyQ5ocao
QW98UekARFuT6+qaJFioejk8GQz3V85RBhc2EbMSzeL3/cPK9lxksAoSyuR/REy/
0SndWFcTiVKV3qMIT8SwReqxjZOgRu+E08yTF7TuDFMN3JCOpagfEN870nebOkK/
FiJSGIK7oI3FKiw9D3cktZa0qxZtpWpjuo1pzl0quBCI3LpWX8Yc0D25j1CHrP0W
+4Fo2PPqBjlYrvb1isX0d/zm5dasUDhORrVZ0aRCoj1JBD5rPp4nZdD/da+hw1UB
eZFOlt04uO4f/Au0kNMVEE7rXO9RM0ilQmC785p/Ox3L4T8yzF4kNdTv7xW9Gw6O
4YDZKVWdZF+kfB2tEYldJuktm6UtBRrq439mWcaj9co+bZ8Zb8aIUEPMgoQmnyuc
FMGZb4TqNvdd2rjXkzLOuGLY+F2AYNFRu0FfEo/tzBZS/9e+GJeKdkVz/Iq8JRDE
g07dPmwCbyD/exNNzs409V9OvZj8eg53pbdboejKGqpEXyGK5ydFepthmXsAzWZ6
hVxcqMUdQYp4Ittg3X9r21Q9EC5tzD1jnc0rKgBZ7jxgW0eKnV8Zs/1SY3b5Muxk
xQRn1jW+yI1+WZBBv+iPn+1CEMkzuBrAd0qAHdBXhATfe+/lCGoezeR7BWUCneP7
KohM9KQcFQqNKdj8kSRRo3d8lUrQ9gxqg2y7HC9gDOcosWI/M1QpxNooTRbcLvqX
XYDAVjuyJ9Cp3X2I4JstuouRwoo3og0HzgYfy6/RukJ/YKJidmc9BzVPEwxCnRlP
p+M41tbLtYGqs8a5KSGHlganD98UkJuQANBagbfHx1kdcYpjLQ10vLtqx8TZfkgr
9z55G1wKSGgmcLgXyR79QtuzGXUCQnldMXEgEChvpnn0OPbrygnxycMLFEm9Lfc0
Sv0D9ZvOqq0BnHr8z9fb2ZyrRJqI8KgI9vxGbzNAFsTUmkCfihrLwnSXTuvhTCsa
TDgJR3RgGphY4JeT6AWHGYQ+vQq3/F+55ywGPIhb9PaKg2o9FFr+IG1/5n2hw/Ok
d5eoQ5K6PVZhaz7bTAedYofHF3vBK7Ze5S1+xf1on9MSYN7kn4Zdm5RKJWBoTCkj
0UVJym2JdU5uxhpo8ORG8E+S4GLVJHB3VjUd3Dh2wBUmJwIjlkCZPlkWz+KmdGkX
HZhkxVO2CV3dcY4fl3gqcJ7it3NEEwDPWXLd8ddLLxY5EBI+UyDjunkB+DHjQ8O1
DEWH8H30b9x/whw78fOxJ8Of/aEEPhMjBxZcCXFtACmoacz+iIdXQTKwt8SUMPDi
GlN3ps9xpluKe1YFgxA+E5EN0TvDv2j0ea0o0RjsWWsBqQWrnK5Jcv4LDpXREHT1
w6B0fcAPxr07jUH3qM+B2MlsjXZGaW4Ai5HyrNtO3t1ILmWdTjqN1oG+39TwG5mR
n8JRHGjvEg28G73pjFJnMiPmzQPL07Unwz5O0Ip7e0Sn4LCHFJH/CkF/bEeuOk/0
fYegXkJlI+so0z2qgl5UiSVx8YSijAIRFzAvfYtNeY6kpN2MTAmsU0aqFw+WwXsE
NOT8KttVyzTgUNxqVlNVKbYQdSeiLiWqu4RVnGt5IRWZ+Rt8RPJH0CRNTyAb79D5
kdluqEQw6jYXZ+NqfrEXgzfnIzchyUTUNeDoTnZsdDW+fLJTTGrPQDF3zszCtaOP
xrx1OZVv4ioYNrGVOua7YeqZLMYTagdKwtUF2JO0eoZRbjNmNRDR+527nl3Z1RSe
ZBKEZrOMtmCeuw/I+M7kx/oHzj4PVg8Li6uhiZC+CvswXBu2g9x6aYvW+lrR7+bM
Zo6ZNqdg2MPnToUV95h/QgBniyPxXET3Kw+hAcT89sd/KkZPkxqwxGegTLPz3lNx
CBWlN1ZzOeVXWn752+XjjDmMacUJjUr1WlrOvoqEZ2p6HjfJV9/IGeQ5GSWafTjY
/N93VT4ESOx9iRGLOjmLYBsP0kCEc1zadJTHcRSKBll4kG1m8g68KKQ5xXPV+vQF
D+oT/4Vv80AdA9wfjGW7CqMtRwnuGlRx15Nq2qWED/F+AWckNoG76RPtYMGSn89x
lZfWgQQVh4LhSHI1uWmzPBcl2QRAXwS2RekwxBVZM1JyGRQVXdGqcfMqG+U97a9H
UcsM17y9tN0xavaIlrW05R85QUhUewuYvP0ueh+3Ks31Z5m7jSlNJZ3i+nZdIDkN
0GF8IfsTUT/QW/rHAk9iVmNgMiaekIlnLbTe0umkN0pOqqOwHtC9MgZ2pVMqae1W
xhSE6BZkK+MPT9VaUkK9sK/LlQ/F3kQzk35WAzdtbmiEUYC/QFwnz545tMvI6+bX
XrZZDV2qiD3TKHOOKJoHE7l6aWnJgFvcPgYxklol78PkL+6vAfRBlc6GETkiproF
iwv6+Ym8AsPqFtXaNexayPipae+ZxlowoS5CGt6jd8cMBq8CqauABMZEn6yzc5cu
yKGQ1BvdnxLUZ8H8piA6SzHqyQ7mQItiRHjFhhllvl6xRzWDJpvt954GDjYNeiXw
EndENzEnAuKg6Q23Jt+udhInYGzk7YR9W1sMIc8fEN5mUaBHPuFofMmmIhTuGpwT
LIigR/fNFgji+1d6KzFI4EHgOjBK1WrKo23ieu/6mGBCzGwdVYfiyRxnyUxFWGNp
reX0A6Im6JTEHEv3ROfQyrNmQ82SQCKTT4q8Rj1+sDiDQo5m9DDO2t/JIR2MDfsi
1cT0vXEHzGS/cs0TuVoRQymYV8W8sXjibHI+HlFJT6nmhsMqW9d8X+uGCjW9irxl
BM3kx+VFHyw3oy5GBnnDDykU8EcqHPVzSU6z67UVO176jB7abp6eDJgmF5wu2Ml7
kBnSEMQKbOVcJDyVJbpteTGoBBiOCAEMOXGzVvU7z6pNTSQbJoflS/yiNGir5PbR
0HjXJ49Xkptpb79DWZ0AIEB7RyoeUzn6lYtzCPQ8CAqqDZ+Lxtl8gVyM5mo8+1eQ
QeXmDQh38+IIZNSf3dhoLVBbCN2e6XCLTew/23/rVTZ7wC2nBY8OS0taDbyDsllv
zPKfSrcmMihTRtpe7trc6/uB2IBr0DdJlX7xwqOqR+Mgab+g8xLTfyniPgQjyiCg
HaOiOShM71ntgCViUjCbya63LqsgqJ74R0wT5F8F1QL84s5dAnEsnwr3xw8cebqF
vaVsPI9VG4ivGtKTtDCkR6k7MgO2XlEsC3yVTgbnlH6Yxby37Sf4MZqSDfKRmqms
O0Sb3n1deLHUr3V4Nf0/cVCj0zrNKxU4oE6a8U3X6e1rYxogb/HXaPhd4yfZVbnE
B2k0DFHmgRN4I/qDbwQEYFWDdh3jDOHB8FU+GxunRooMmKiPIV4GdqH6kNnGfcP4
OePJo/+olwJw1za2d0GFFcnwgKOAx/1Mp9l2L2K1DYnMD4NvrdXQH1L3wjJ5ZoK+
DU6X0vsGiyE0mO6xZPHJ2crCkhE0iljGCP8Dgbd40VE+sP+uOHs7QkAebtpDk8Qv
mKpOV7NnxKnUTZxbVpfjFibdyeHZuJG2kx9Xeuv61aQqe78tfT75gAfZR8R2RAE1
HazX1T/QKUasA1IrGaJCKvVsn0mKf2s5hVMbglu26Us5LYwvLjE/cVo1VOuwYzKk
O03NY8MNq0heW7ubz+YE5qidSlA4hNWS8sAOPq8I6k/BDE3ZAODq2vVPCiHEQ+HS
ff3NAj5gvXHFFdeYLVUdhQ9bg5skyUgrdPq4Vlb+qvtcl7CCH8zgpFjJrD/nU5a+
pqkQX5hA7YYli+ZvzGnxXjaRdlUDYREhrDFK24Id1cwHIvLhe0u3x5ULhurXDDqU
k/eHM5jS7MhYkf0d9BO3XfYpil4ftdFQVbwpllvTODDgm6uIvpWLF9jIxMHjMns7
0MGW/PsLpzjCT3wvL4URHK2b1DadER9eIXZRpX2Irx0sd5pad9ukrY+Ezt03rmrF
8t35ZbDmaBMzTive++5Uorbg/ftzIxyECUeYkf4sDiPRcCP8xdIce7RmfKjJHm77
Mr7T8I/q+ot0Hqnj6zovggAPnF1HFAjoz3pm+Osatmx6YN0oYtXpS6XchFVL4EK3
CyY/SzABwE8HOwqpkpaD6pLLk6U4FPsSUf0ZF8FijHfkFxJb+07X1hFwGT521j6+
bofzGL3oKIAEyX2HlfMETZELG1hEnjJ7FqYceTZ/SCO/GQtlh5WeR2e459oItsmU
XwfwbvCzWtg9XLnSl/zd7Z3oI2JoN2cgMR9QKfeaCMeGAPuMJ6hCMe2R7CbC0iYX
kgGunC6CQCLHCeVQfertjAdQGOOpUf5Do1VTJRWFvKGw7MC8beY7rAE9Oul1H+86
lNGRyUiSuDvzT29SIE5XTM0VCh5adF+ziTANrsy4iyZSQd7HszjSBaP4ffTdTPYO
1fU3XPS9WEEhMW0DMyP+O3tC5YQKL+vJL3IxTlCz6xUccimhdj4aHGQVNMc6RP6M
gVc9oWLwmz493++0svJ8fwvXykHa1ofawF71wcjL0JDuSJUalKuibfHWGtfsJgKX
YVUqFQcyCsLguJQoRvHoa8cJHgJRlbGduVMJk5JnpNrgoiKC8rRZ1xmvSPxS+YBO
g+9B2t5lsmp65K5v/KP4zNtf6vNcxA86VKuPSc98ozeefShdF1Mua0Nas8dN623h
xPDlRiZPUrlV6L1uvCJkh/rP216MbYt/AMnPXfYae3ck3G7UcX3KfkKijsyUqWNQ
eA94V9jpBB3lhRbFvqCWcGsBItNWQLCA79QpfFe/05ZETNQ87SnSUpo5KjaGHCFj
rkfdYcRl+Er1wOZqzrYW/Dd3W3Z189BLzFD11jAIO1IHokH5eC0AyODPfFWYxFtf
pwLW3afNxCLI+ZKfIj799VaWuCiywqY/Fbi9SYaDLb6R8G4zu7ZUwOLWBTIG/opR
MleeYvA5PQ86DZZfk3dFhl6QyDPW5kI/N41jFdoQU3p1eCkrb1CXCqTGzN7TorqY
CS+RtSKG6FlygsDWk3dFJb/PuHhOQXHWdrJNoM3cWW/4NAt2LOSQq6u10dfgaM7f
P2YLbzW3nQ+7oon93ggEra6aoa3Ksqr4Ta89BGSSpKL7ISlOM/0g+B/xOx9FDaDU
u8xY8Mvvi83PLTC5DtbEm3fB/2PhcK0bSgdeIivTtQJ+3e/jDEPUo750dK43e/v7
9MXwGqnF+3S02TJOK/lCLQlKEb0cD9iywpAiPD5ggwk1030XmubgcjZ9ftxnCCC+
urL2V2yz10D0OL1MasaCQwAjjW5ISJDGqDsGo+RWJHjL0DbP7KXXFv6KbfAQ1hxM
InsNr9qMsmhXCuf2L2TSuyB+iLaQz0Wldujk/0JRHVvXcyLXI6B2kDXVSNv5aGHU
cyDf3AuVwIf26VDOK/ER+LzIDCpYYWOSTYd3kgIyNRp3f1FxAhDTXmvMir7M0f97
dVTH4ibIoAuuis6jn0Mi8U+1kiTZ5oyvsxqiYfX23hcd0R5GBmt6cvQMXYN+1iHb
mj3HJC9OyGXBjOvNoPWVwJlP58sRtb0cPNPdW1hZi2bJJIiCECUpXXt+CCpxR6eW
haYMygUZAPXOUxyFU4dQ5JugV3uzjOGayb4MfB956K/nMsIpaHy+fDXcdskXS4dh
LwtwxWamxe481gXHgzP4i/CDVRieazOb5CUEmEsJM3NCg/dGTu3HzFBn39eXtjVa
/oSgR6bKjkjfPBOt1uKv2jDYO12Sfau/UbMqk/OAiuGcK9EikedNJrgQ6rtdUEu8
WtXmCTh1TKZnK+q54rwFUuNUBMVuZ4aci4/SjTTJyqae1A8RSgPOnr6sheuzy1+f
ZPJmP9y7BkGE5WWKAE8PaO55Zpjj6TgDnvyh59e7XcykM43GNlhD1TMM34jETgvs
5vz8OB1kSrVtz7V8XRWyvnok8SEtrk6wUu4dS9Xvr0RrqPcpuQaTYr/G/rsPavdq
olt9Z7Ccj1JciKIHznhjkKTOovN3KgIwCOa2Xcc6eQdqh8bE8E9lDk4Sc4x79CpD
Glt26qC2gASXaV3piGVXB6pfWbAYmSG+3cgme1CjV4zutkJiRdAZQIE/ExlxhG/P
SaGaDfi82uschRJIMHrDFac/eqwYHgSqEEHBBAADgqUT2at8kwdwGVnun+Ioy6fQ
B48bG1CDiBdc/4PuWVfY5cnJOA7fyc6WoRWCi8HVkAp9et2PqwgqYUyaZVaueUAr
CMSTOG0Ce8TcXZpCx8eKE8EDrCVn6boPMuxCXGuE85AgWJOHsZ28Qxt/ZbUA0gGf
sc00xTMJINuxn+a9v3mKP07xYYUi6XrfPT2wmY+q0MFpan07kL6dKf3ra6DI2f+f
qt9FO1t78g1hUTD6kHBvxK6Ib34+mlYA6ghlwgwuYsMw0QonOl//OgUfHcXy8Ny5
CZ+LpIGj/fcxI5c56n9FjmKD1ksEoTtb2ylEaIPYeZs9vQnFnjn6eUGTQWw6ZzGd
NbJVRj4htONuw+jGJ5rIC3YZ+XcdO7D59bQgbtEI9unrxc/T5mHh48yU7XfYVWay
5+RKq5rw29QseBy2Nw4XZvGO3wKL2q5H3QjQ1LdRzBlWG4JI/LSwvQldn3b63qdd
QmKbhRX7mhPP7luoP7TlsIZEWxnqQBoQAUzg8OL1kfucRTgUqW3ppMGrc5OfstZr
znOShC6HPRT5kAudkR4zweHeJ2rDxxBAFAf3a1RuNLqWS+Mdk63EnAh465AS35ll
GbwDGUoYQ2I4/thoarGIN3L2KAxwGQctPNMjLWu1qRqvHqneCYo/24LTw/V99xXy
atjkWOrTao307Om9PHyFDWTZ6FuofZ50eO2EU8655yDjpHXXKH+MDeLTZa8mRr2K
AEUEG/hhw0yn50hcKQYayfMSeGXgApWial/EQY2mUV8aeVEXae3N8xI+Q8clN51I
iEIr/bW/PJ1e7BqOu0K69fsJ1P1FEbh22yBubit7mMa7PqKzzJ+2gr85L1rhBm2T
m83tJ84yjjkJ3o7Zh9siu433qXBwaS6FTPtSR/ia2CT3u8s5DdZDuiWk3K2XkydY
FtNDZRslNtoTYY8PyKwu3QQ+e2iWDfzeOqqQRNqoNbJqvcUhzI5eA9IBJQ+UXJCc
0brwjXpY3bDVHWwSwlRYQOnYZ5EqwJW2gu+J+H5ihYxre67dRH8jYk5uuSqi+kNj
AzjiqwPP7LpW53SRCT8/Ea7naTyzgBsKQfdGMTahs2syn/zHgMT+hp9Lpzhvaw4Z
Loh4oXpb111Gdouvjh6oMAaHerk1xUh+TZDJRP/Rpj7k7g1J2/ummwOQ3wulvXDV
/auPDL/Y/VDsG/LuwOG3a7glz5Ynb0vhlKqrRGosPWEYIXWreh2hl0gJJ11SbbRt
PHuDkQKTrbV3Tm+kpjLcS1CWvvJYeTvBk5z4QMXUglDPxU8dEU2Rp6CWZuFzEvge
aOPQOeTJFPChhzZ+jN/lxcW+3IA/EgiZzv65/CPX6b+8RT7XfePdLziF20Kr+EPX
MyFbNbaB314jWJhQUzQ6WU5LhWiPA4SZOryYuBLGB6GTv+d/XpOEkr3lQsYUZ7t1
s9YrA2ziB5VvMIGE6A2daKPPs1dZOkIpt63edmlK4jSf6juQvDvLI5cSBfGn+8NT
yVSO9bOXl1VxFhPanryhJMnr0BQUA+DdmtgB1wEdeh1/j40owLgAbYC72HoDW4zo
Oh5z2IGVxZX2CCRggxyXV2LY4kPd3IIOORq+jQfRtLP7ex5E1O4ghg9C/SNeCPMQ
AxPXALF0L843KV9OvdP5DIjnH0gm/euRlYZQhfzIVNLtW7h3f67XyJFuUq2zIJ97
L0Jv7X6p/2VkW6v7n81bdc24Z7TVfbpsj33mwAQya4KKllQoy+vWMO9W55E3ZhW2
3eCATpDw3iB3PVpsuiHaoEnL3nkp3Drk2xt1g1Lq2AnakXP5MEFO67wrAonTROKo
LAfDmohafzscwN6zULPyzmhdUAuUdB6BYO2eSewI4JG+CsNYdVfXvaYZxeL8K5M0
boeyIES8ktRkXQw1asuKxh+4v/tEcXzEneSNM+YXgnOcR28tI1i5hBxFMgJrwoD2
sePomFMjxT3rACK8eJvaUmhVWwfZJuUqE8a7U42GBWKd9i8ESlhKLnd/PYxQwT/0
ToSXofu22MNIQHQcX4Su0t9jmWEgwt9j6H++foMADBXkjWMpi0RQF3XoUYclUGKg
CoJs89n2mmUAPVB1vvb+HL32jmGDijd00nAAD66H6/EctF6hzAnjhAwqf3UCNhZv
3Zkv5sj+jogURrRiU+iKcbQlvbMW9El1esOSbGF+y7x+QtGUQgyP79jCbfb7EId1
Kmsbx8wtb+jF4H/KG1ZSomA66jXz5pSXU9XugYLy16cGvvTqtJEoOrDC1mD86iYs
0Io3lvVhYdYg8sLKVn6lIofneUxsgboIuoEFfcUSFYbMyDJrM/aXP1XzOuqbE2Aq
aKnCuFhbmfBAlQXP+UUr2nUEuVrJLWA+5PM961ZfcpZALwmLK+rSvMQ2113zac4u
m1qF0EBSUuUWzuNoplCcfB3OgHjcisCsrqqEM5GTUtyGgcl2xsjSMoMQyWExtp9t
4LOOZ1QB01qQCHqLTGI7RDfZBcLhAhlU+I3iAjtTg25rDzyheqWNotbUMZGZc284
hNABLgLGfAy1aYLA70wTLWl3VTIYVy4LFERYUHAtspWPCNBtJTClBq7ctVDBKCP/
Yhd4PWphte1YxniPBF5P3SmziKAtqTNB/a7QLVEiN6A4EOzJ+GRi/LrJn1TRs3Wv
HuMk8GQ9U7huXaSDjVIquXR1z5grBez9rzXdAIIDj7eBDZInYY6fsQ3q7YrONm66
5ViD+o3tP5WTXwqWV+BuIWbCJqyjtaZ+eFANES255K8zyQCO+YIIxw4E4JESEDNA
9Wt5EojY9QQnzxJdatojQ8lJ61+oFuJw+src6yk/JX2rzswYZ+T/qrPnflEPC867
MLSC5/6PGKl01TNqBI1aV0hoe037cKJ9T9qv+i4xrJGYlv7QKu3qjKC5PBj5hnnd
9g33g2RTqcLcCE+IoT83DmVU/7Ij/Mjd2pCrEiOaob7tRFyiDj9EHHsUNMj6cIMB
/nkT+Ht1ZE4mFnrAkhmTlJFUqLDabPewLNgPJ8fsA+JpMMbABbJomT9qeQk77KGX
F/VSGPOWG+xTTx7TyXKBwTqCFkkTeVT53jqVboBk/Kz5BO/msaJNweR2KM89kTej
4bsXOADadX8ENu+P7seBM7uoXD+Qp3OoO3U5GekZeptaLt15NYWjD0SiyHTao7kX
i69jGOy1Zvg3jtWdEso9Rj6T9KNKOwLa5CR3BnithbHsnd0x/tpdpYiY2cGX4ave
LnqGyeDK5urflJryYVhCFLp9LpmQ240ulv4Yf7bbjkMfUK2OvT970A/IIttnvf9K
kUKlj1VO7skNm2rdctN6RLi4fq9B9HZKqOjuy52oHtD32G+lQx71xUwrtET25XAS
B0tR90p3A5vyju3/0y101V+4+L8oZ92T+f8euc/SJ1C/LniSYisDahkEjIzWZr5K
B7qO9eQujavPdUaIezSvFTv89aESmS9tFqSZW2RaWdKFk8ImW7Ea0kL4ld2DW2Li
mCdte60bFni4YEJkbjCYf1eY1opAHQUuSpNICXjIudq6MWpUlU1FGLEuUfSOfQKn
kiRsdQTqy5wWJS4aRvZejfaOgq5199UPdFxaxarZ7ywzk91MJiggeU4Br+KfMi3D
uROzTP9Gj3akeqrQs/ybKFFOCYOgQvv7hZCtji7suAwlPBH35ReMywqtwfCroWDL
lDsDlqiaQgG0yGI9VRl3hDnCIa2hXucI2XrTZOJff1RxVdSV6Jn8YxFB88YGf3RD
pT5kZfg8bveXixG7n2PztcUD2ZsScety7GiPlpSREi6D5vAWRiH5CcA0xLhGTJZT
RR07Rc/TUTXr6D4M7dt3kH7WF7xEH/S2dNnJRB4d9R8AZ4ZniKs4vcZERvi3WVVu
ZqoL5drZrEbHVsFqh8GTkL1v3ol0lyaRgvUOxm8Y4zJPWSv0lKP7AEphsQrjJ1uv
vb7LonRNlEvhsWBNkET8wSKssVKp14TYQ7igS/iMtgoHT6D6i8dgP+PvApn3Lgfx
RR+FgrEzOmkUrq5hyLktLySgGvRKj9gqGTy2A/vngkbCsdSfIneB2yjYMbbgXQ50
BRFh8J+eYE8bzPeSyAQJJlOORuGXrzKo42PH7Qo5u3NjBbGr3g4GRNWu+XGTdzBn
q1vuYXWfmDujljwYWp35zQPUSNEdgvkQPh/gMurh6oySrh/ze9QyCoY2eCGM3ssN
uOfyuCFgMYihD+F6PX8ec+4QolySsWcby9K3hGS/KhVnp4Ht7MR6vUh7TS85Z5zc
VBtTlwqkxX3sAAfRPF4eaTHam4LhVLR/R/IqQn2I1mHFLiby3HMlMC8wdZYku6zY
9wxhMj8IkvG377ddzWZKdYfkwbIDSdNb7HWtga8Le+mf0x1jHI/wdPWZZslQqR7C
seOSgpIkldpEy4QfZV4FgBGcLzRSbinYWzBnU9aT4Ayfv3S9QxDYt4dO0U3oxjEc
KdQcQ/gytw1Y9uVCgOBFXVXp++hIyC4V+diaL2cxY13SqMrVENEmGPPemkQEpyt9
Jla0nBrH9tVB1onFOT27gBt5lATU5QMkl0taNZa+pXxLcuCrplq14aZrwBNjf+vr
NLNa6Y1f9WtIuW9CVqrlsZRPucwaElAioX7qBRXVRkOMjuM7EAX4YYDVJ8nlAi+K
HdojyJWFj1rNqq3twFTuWhf3hjKTX63QYNu9/Y8H3DH+kOsxL/f4iCgBnExZOjJy
5hMJPPl3eY6lNjZ7Cc15Ak1s/RhkNfi3Cmo6gBzpmwMkpWu4fH2tJ+XzAlAycxQD
O5uYw0NeTI+jl1jwekxqtCKL3oGs0AnGhiPxaoWz//WBavvqpfk8lJfFQn7dRVXm
PCcyr/neezFGGWQX69uG75zrxEhjuUL4BKlPQfRiYBgtjqHYFBl2jaPkNvh16+eF
3YiE3RIs/XSRygYRitiPUSl7lLiTxiyrBEZBs2yYZxSui+eZmIb7+OBcBupmkO3g
UrpQQ80acJW7N143RRJ2Xr3sRHn0fE+JvI7tPYPmmElrcgKBESl2D9IVv70zPxyX
ByWzxlZoBq7RVudxAdEgUgEMT5ySouBfwUmfG82fd2J8vzYDhegWy831EQLf8mK4
yQhmveplcucf3pKTjPrb4kVxsuW9ClhATZk7vZmHo58Wvoo0JaFopphV16TZiXXH
zkADWJ8y9qUGQ4UCiOw1UzofZZL4rxhCGU0uPfeRwPmYySaW9+tk5x9RtE4as1go
kQ4uVtwHxYeg7wzCyFpVwU+dqp3zX8tpsAyMwjPxm+11eIiEKM2vpRBuMiY/HViL
C5N6IP1SmYqmRp9nGl+84Mq1iC7b7zs5MOEJYYos6hnzUGUvdhZdH5XYOqNOHGzR
TmZD6GoJkEij79uzSTDJmSmiJqaSAVNjS4RPgFCCRhcesfIAy/vUO4yoeaw880Ns
EeqjG2FnCojwVPkPlRjGkJoIWBQVBHlruvydSiB4ACFW6qB9698Z46Vxo0Z8zE5k
u5AMdyghSVLBWN5Tga29x0xvYgt1c8s8ATFrm0c2nSPn7XaLf5trxXf3y8mJPKqI
ZAJPSREbsxoojN3ymdXl5ik//N86MqZ78ntMbo9BBnksoxbHuUraG9miHAkZeq4d
tnWy2Bi6a0q5wJTFzbn57OjJyUOiy1cB/KumMxR0ICAVf75xVZzILqpo7FkMgJkK
lYYGNVtpbRQNLbPnrH6Smo+Z1x6YfMcKv0YyDbq0iqtgnmgtWykLgBQgXsoltc8/
/3tSj8yf0G4T7uXAEYJIXYRbDB9Pm3RCnWsqd2eO2gO/2aC0hNxknFmmUH80sefO
QMf9ttCQhtSBGSDh7wIlRgQlFcE2UlT6RtK2tDvAaus316szyV5Fa3TtNZYLLmx8
AtCceNWSK7EAKWpBxCOdItZQyCJkX+Pet73oIU2C52BMoI9tLIdMcpuApvUJ8nJy
HdEY1HmwrgiBXM5tXAOZ3LhZoGqOamP1wEmyoTyL+VN3s2Em4rSUB8QFdkIGA/07
kyKplliWi/wzRuGxoVmqcWDzm9pMepzBTuMFIAPw0NSaNHRnDJYkiPdanW+TsilZ
03fGKw4br2m7ayPOtIpEJ1Xl2prZv9fqHA/8a1L7Bl4q9XyILaioXRE0oPANbNUR
VatJut2c/DaQJnwE4GLijuLApTI4i1H+596cLffPJ9DZ/d456CPKe4P95CZrNfWY
b01yN5CCEVJwQO9oNQRnr1I5ZrgC7ddggcTb9TgWRdarGcyiSFRtcXb9f99XEiCX
5AyDQbmunlD0FfH8k4OJuJV7NTIChBtJEcJcgfTZ/NWVsk4WpKF/Si8IDO6qo0dh
5SfdiwT6HX05veUn9fOfME5TMpPga0UGG+1L59tolfBeE4/e3m1ZFcU4877pXpOD
nNM+LOj/4jEzJSu/bFT5ObvyabDCYSJgxrStFsVAuyaJ7o2PDta1bZKTbb6aJHrg
yqdyOI0JPmqd3LUKnAllY/U54OV2R5Jq+v+AnSw2NvsxStub9I8mohI7kDSf9wNd
Y+H72ZzW2njzJ8o7t5v+ZOvwETOeWEnHs9xy20JgxsqRYYjaGwQyzfRiBuEHTZ//
ZmVvP2j42kAdiys1ngXxlLsT+hHibcsBCW7SGdAbZojixrmyMORxQO2PCxyE9kfp
TqropsSpAUh795R58QiFGcQ8VnCYT4i4NZx2INt2rluAEK34rS3KM1vQR9KviyZO
tOPJ3HeewYl13pEmrLssLYS+0pg626ee+0UUUt60AJc5NkqvU4U2c3xL7Ld8NX1S
FLhUjMjGlY5U1cOkRgRMprQR1+EM4OXLAc2TJlAxi3FxplyFxg962GDIYeKVfGEg
QfZXz/P28na2o77YpNz3/LuYe2gRcEmAIoCpBSSGA2lst/nNZyqIFS85rPCN7zYD
pKoEnLAFUdIPfcXvw2BXHUe8AePBijBi0t7Z80ynBsNE+pmJyp5i9pbXIufkmL8l
oT8eyqp90J+yIavLPEy7sjNJQsktzhOe4s92tdzgOyEB2/lLnU/91CPGXvpWin3I
KduNMcK0u1hHycBON+p0t9H1SV4M78YR5dTI2teqjGoPCYm/F43GdIVNhWK02U01
1+Iyim5tQdlxjdqvqTKB7rt1jPWww8Cfz+xoOmQBpynpeschh447XxV0ajAWGIFf
XBtEZGDxTCaUoKdrxLZq0WBew3/4iLw/2DWfP9JuNSqiGOzQUtU7iQZ3As41OWX9
cuw9We4bVxBXRBGxrZnVJ59v92OsiBMOiuIQSKVMEc7gNOa2yTJcIR1GCGL4ivoC
iGZZtjwy9tktwsy5CFaSzzklf9olZoM8YOgKk4e3E78nkFvAW+lE5WKTv/DEGZqU
S/PT3D4KxXA8p4RJ096Gm1WBD+DcK58172c/skBMJkTzKufZYdFng24VKiTB1OyX
SzlEbHpsfGBWxjhOGEuFEK86fSxbLjb2jKL+Z5DhxTNiR6azDA5/x0yjygeHitYC
Q0qyR1nXJQTCLhg/hpoY5Bcmcunl42IgcSdNRU0iQpY21j06q5pT/NXcMAvQDiC5
+AG7U8qnNl98K1qFIeB5xlYrqK58OB7NcZAk2ZLeMu1hVt0DoEjRtfS2B40U04we
rmYHFNQRg0wZnMLIgBE0U2ASyDhAcO44zompk6k9D/aK+sXn4FSH5pOzA2tU06qb
4iJ2lA6gh1c7e85wAt/uS7EvnvFMz7tQpWJPgZlzuazGwQrUFji83ZnBF6druixF
dia7E8SERe9fsA2trkV5J52pygWGtGeGZXbnfm8KHgpvxhxphkQYp+g3wHC14suU
mMbV/zfDws81c43ikW7JAEjIBufarMNkLbBhjKdPUpM97g/BisgAh44ElvQcLAqy
uzUvdk6Up/7BhDddp2NagDeHpI+GvChNRqPImHH0hp2NEfT3pimoa9qeBWyuxXi7
4NtuElVje49n8lHzMkKGNcDRIXExI8UlKWlyr0EGCwEoGpH2R3m4R3ZKrmVS89sp
o6REdkyWZ3sX226oZ7qZqMsDkCXStVa0j/QTSoiZRBbVyhm0ENv0saQ4OGnaEe7n
AFJfSMr4Nf1XmFURiKiKnvgK1+R+BXHT49Z9naR/Nk7OFkxiSLd9NJL+TZqXCcgN
/USA6wD7ocQMeCtFzQxaOn81RbbLTWaloyrCmf5e8SDOjdPW27PaRF98BDnruz1z
Sl48mGPI1+uCZvpkXxR25qqOtozXWW3+vqCgJ3wOeGnE9MYbjYujDn6sTnB+gRav
x9ydBBwoDLO5VLPBHtd4LhxbfhAKKExyULO/kIiDDNBl8lecb/+vBWc08BNF9uTe
ObDLzAl/vUWrF16T8r514RlhOoRLF343jITd6u6yScSRl/pf8lyeG/H6O2054ql2
RUn6/CU/x0at7JZCs1uiVBRfgubEmX3YeBjc8cKk36rwsjtil1wSAmVRa2BVpIpN
/U9+y4viR1g8NeLiQXPbxKVVBsyKUOo+19BupLhpGwoFUSkRDx0AXTnukzIxRGmJ
4kOdpEB7h0CsXeGQaQ7BCfMPWCLLwnjNybuMMZaQAVIUqJTjc+AijecaJc1pi+Nm
3GKavF4oJwOumWGNw/FYtLfejXf+5B/nkWS4sCvykxv1eihcXFmKdTA0YVwOH1wN
QV87TIbOdSMXCRuisYqbnyvi4BEiPl+U7zuLTz0P+stAimEc3T6vNrDqB1FHikBW
Rn3KF3RBETOSkCyJ73bg3rhqYaDX5Fj/zZairOHcjrq2cd/tY6+JNEz50H747xUu
xIRxGbgRpJ6KkXb0d1cB3bbYsvN/5Q01N0Ew7VuPeGdVHH8KXbQA43+uVgI/8ElF
tZjDBmLCffPJOTsskHwNItc2DemUYloS4A3JzkHvi/OemOgFBoZDZrpWVtLjVozT
yiXtXjxjbb4SYajFKtNFtNya0C1xaW5y11mqJYNsterC0No6qe6YRuxcVGirFf94
JdIcwkZzAPXvEyzze8gMtI2HXS0XG0rZcaOdTsXVORknRh7oaPTXPeQ355UU1utm
R20ZItUINeBxNF1oC9iGJD6RYp3BAqvd/GmoVuQcVTsgVHNuIYJHUxAzElYMoggp
Mfro3BlS7t1m/573aFjC68nNkdHfPuAQ4qVXS4Fbv47+PxTpMuBHMnMg41c5RmfH
wD80Y8BJFPzL/jIXdA21BgP+7yGFIgIpqWqTdkerdXtboQ8EWc882o7+wdLRkR59
nrR56NWL5ecmHSH8GwpiDuqL8Hg3D9o8PWJSxjoV1dT01oCLBv1IoAp+6TFKbtMF
5DbqZ+B1CPmC0Q51vlU9em7Be/hewtY24d5Crd6BKz4HbXfVF2cjavGWljBsKBQb
C/DbmHHql+NllMhjnXK3gqi77oiB8q+oqPNGu1mPaJnPr1UaHbrFs4pdY8SwTXKW
FWGpHvG4gpcDtu0nYexnxeOqCW4HFMq7PghXEmyvLWRlFp6wJaYw34HnphnT2q6j
JB6lJ2LpgpK0DiRVK3oowKGMcafQRPW/AYjZ8jBwBiURA2QIvWhDF3Qd9Go8l/Fj
hWR7c/+cpYn2DiQG9lRbWl492PSEBCn3KVgp/EX/Ucj8bVS2Ef0eUXqHWY5gGebK
2BH3Z5JBpbluZ/vm6At50zrjVENGgh08l11RO6Zu5GUpIz7zuUnKuFxUeAlt9t/Y
kMBTtYzL1iCmgmFSfpelL7Epqx3wxudarukn8DyPZajY6TS6wap8H2hndjGgygb9
1N1035cYMKeL1meKYybQFVkgrU5sg7iRT7aP5d3RfN1alzCSRcDQx0dvYiEbT7mw
3mqv7oWmqEYkoG8RcIvHzW0BqYZeUohGY+6s2++VddO9kOFgdfkcB6H0eLepQlUO
y58nPWu35C5xa3psb9ypiMeay9BLcYOtvXP44NWuLnTxuEUOUB4Y6q9tJ46Mto06
OuixP86bqY4Dp9NpldiWWmr5gINDJB85ad+6QsXUmeqmn23UTcjDVoLRNTme8fPM
lwhNljebX5wHKo5nooVNvfMjLNgbWo10b2Hn8mODappx+fBviPwcyhj6WjEtTf8P
nKeciWbsbEU2ZB0xlMHLbU4vGxz5saKdkQN/+a3d/XTLZvpvi4ifWi5FT9nh7xdb
KhsL76ZTmLH85/w0I8sTRP913uaOEqiyQ+WUvwZFvWvk7QKuthQRlTZCxDuBeQSL
mTT11xBAWZZ8YRjVHF+3q6Bj7koQWPK4IVBL8RJCvMSpg3HgGcx8iSQgTOU62ycb
uMGfNPrdtxdKINfLHwQtrhXZRmFlOW8/0jVj/rthBhtKkEHOo+RhamxgYhscJF+/
5nlvgbMM6cbzUpoVfTezx4fIJQkER5aWCmNqDcTXoH1FexjR4Bj5ejim0vnphaVJ
zc8xF7qHmFtynV7TJEm97uWDqZxPmiZNx9r37BSR/NDOJkPufhxfgGNxbsfZVVKd
b/neJ7Sp7O7CnJ8FFmbXXslF7iBj4bo8IEJTg2eC6IqpldZ1PhZAzCUHNKm7gRGh
y22iu1LaweGyNGKx0QhnXha/tzSbq7bfKKU6bvwVetkwI+wPsgavBeUB53KC9ONJ
9eaWyp30q5QxiBiC3TRGM3V5UUQaeE+bZgRsy2sIZe9zKrJGAhfaTW3i6omLQ4R+
JyOKTnpbzWcjXwIDy+if58NJvwcufBKIlqWe6Bt7Azz8VPQdHGbSwsgAsA7YqjtW
rsp+vrrq96jxBHTN61FKzaTuDvyfaxeV/a1HmrxT3JAlL/1g8Ye9iQMCtKesTLag
TIp6Ht6njTYS2NOg66CpcRUIdRWP9mSim6+L9fLuWAw75RP3gE1p/HEvp6zmk4l+
S0+Qhqt8S/d8ahnfJlxvcUansDphEWg8kTQAiwlSfEDyjG1fsNagqVzV1YkGqdpG
i+7w+K7xFvE5kTIuibo2o5xmGTCwM8uGicixj7nZH7LAlGAjAtin5JltPXX0jtTt
fU7pN/M6lhNoJXrQYvu6Bc0I8DOVd+hDaxvEhfkxiDfMdz6qkcRVlek+FMWDcYFT
D0gaKRq+BtNqwEl7cWVZuNPcfPKsAPv4uf8/J3MSe97FGeIIwaGv+Sdw48HuMiPV
sjMwlkOIRckXUBasy7oH8DPfwn9rwLlP2e7632QkGgtjgfwqJV5UH8hBq4cR/3vQ
1QrCVH/EebbKJH0KnYkheHvJu2bWxZxbQNeDefiQQx9Au9BcBWYhfXt6K5YSH+Ue
GeVmnOi8gKUlUl5j2c9qFXORSeMQuqEqBdKcr4HOMdCNeRuyHnbn+J8iAyvqH8dq
AIpem7DRkvWKkEsizmhkpH22g5w5/Y7RM89nZ5BSKtpoJMMebM52TFYsugweS8og
EsX/lGAhuGKyNP05NVCH/bGvG+6xdn/ymckrC3VS7mNbsG+VMYkd9hu388GB06sM
EQVIldwv/A3nm9V4oR6JeciVoKLQyWODb8En0kdDEbe/P+OgyJSTd9IhEmJQdCaS
NOSSpggzh0ZsW0jFskJXbJZNEu/aDy9BTbHMvh5CwOSd9zfx1nv9yTMPnJev5/pu
qLTnWH4gIg3tmZXE0JWmSXedRCG30rDLN7ckOvjhwxjiQ5bM3YUcUTscmhpmT2sW
US4U4QGe41W2eX0YKKXJlUIR+XI+AfTrRf8zftewo1j0qwLIXdhtEL5oYE58K2jT
k+x7hPvd12GibIbLNbJtiLZBHhuP3kLDFZh4oIsgpQJTFebQI7gMNq5UEr+mfooh
ka/j+S6h2L1tlwd/F3+P+2tA+bsMzLfH95dyUD/5nRdLAlCd9INMU9wOnXvRQGJN
C8zasqqulu1L/EPaoPZYEuAoDBoTbOtUJLXR+ACiCVdsLmEi9799QxRs2kSvJm0C
cGUHnfBiSSpYLz3Z4CYtEaV0g0bfG3gIwuQXXS1vc3TMSJkknjfRBJaZG79Vms7d
oOIDQhlsFelOuIAYSFjoL0tmNVi4A4vjPqC7T9WZZ8ICobVhxuabPObsk+vkSinr
DOTbf+fneCayA5D0iRxX0rHt+CDs26s17DjWXy/zuHCBGxwpTFz7Ay9o17fXs6et
E75IWOq60I9NWDoyBHewsO9h98Yaj9vT40VKzM+0QZDOtWluewketmXdCX3L2F01
l2ArFGjywNb1UzE1q06/VEKINpoEP5BI8TI6Y92oiwUt8U1Z2u5Aa9NbqzTBPHEF
83s7DxLovBEI0aj+LbRQ5zL5KBdhcl7Gqftxv8Ta8zSDiHZLeasJT2kljnpjCOQ6
1qUwbBkZLznKnSlTkbWMxCeQh3ljnYGcRYQIKuipclh6kJqVP+m002DWsL0rKmgj
SUE6EvUppMfeLP6KjBzQX2Se+9t27NNLDvnPrPJNbIPk3+N+Kwup69YGLKm1Wa+Q
cR62eZPrA2aiqWPoaaXvLwGH2vm1LasniZ6QnPUyDD7YuzkobyeEpxhjdCVnnFQp
PIF+dn3OGeORQx8Cd+3R6ogrSdDurlUMCx4qFAz3rp+KAACjG4xH2LLxAlDI0Jm3
f5JsjAOIDodued0BWQwW2wdoX9RJTGnqHhy/sAuRTmM/Zmpb4Q3e7+5wkhFzP74I
+wLwfm8phw1D5Yw3dwy1mwZ8219xekTED26M5vXgsQ3UDpFxU+RN+qyezMuGzCST
7IlJDDBzD7qy1e5yf5ljc77TbnYXYGqUJZuqYihwngfJHDOXMjOtQdSVf3cD5F+n
wDZOuuA3MQeexeSWp2hVwkyPCR5RskQcV14lua/ojU/6lA5RD4ZJd0/WmTFHvPa2
+eQslPNWDiMIylm9GbTe1X2joipBN7ieNlEwimhgSAsfz4rR132dQ5sJBzinP5ST
la6ziNa97gBVaklHcq37k6bB+PugfnIBrp6zP6DI7nLqnnoJYFOIzDRqDm7T/eFA
kVusGsrPqwldrhZMSRVfYvVJDhstGMaXPQo284i45XZnP1260vg4m11tV9l4WcaH
oV/c3NOCqnoDbgYXT5q3eQ/Vb/YtL6V/qyRcJ5YurV9gEnqzfKpAK5IgLIROunHC
PoVxH1eV7hRZsI9Lh8jyhvWjArHuotvtDCkx0ZVjvLfAibnvknXxaGshX31Hiy9Q
p9uP3mSF5pbqA9IvHUeA5elsr1HudbhLeuNm5KVib1YN71EHmaurbHnUiUVnm+P6
awx7v4+vNKjV2GNKSSQ6vYR7Icj1cpWJqH2hurhfSTUg2mcTGmgXCZ07Sx21nPEf
shTk1jeMmzTmGvKxHa4+JeOjCdNEivV74cLgqCK7nUkrxaZwcp6du1i5wcq9ucwO
/sfDVR4TzVyul7Sr494IYQ1NjIyBvH6K7wpKsAgd02WQRb2ib1H9w+Lmm2m1z/JS
b3J1zEBXRkSWVMFppa+7m2B0GQejESbqtci0u4P3rD/CHxAVmf0nLRXti03yEKQo
o0pZ2i/nL9LnfpCMagFILOmCw+0vGw0IawQMbhY2McyJL65ZbXS5P9kHB8GUnJYW
vqgaQ5//b1l+MOeGboLaB20XRG+9Sb8j6aXcdNC+Hpg5ncIw/b6ejAErBUZ6qNb3
zA1vl6wNUtQ/PTSzvtN3P3yqa0zoaFFirMTLJBUBKVYtihoo4ywJTb38QZpfDgs7
x5QmbckUZQeKujLjVbveoRBnaftwQZjvT2XgAGqgxu8K0vAO+62PAz0cj/5YWlEH
m0l+7RiRq8F0vb8KUwjGTgwTvWc7ZqfQ/hGbxqnDOYFLZ3Mz22jhTOX2hAUIsqlX
4PKJYwXE4rcTYLtRYaU5lt4tw2tUAP4M68BriZwjlOW2cheCiX48sCMBrSC5g1fc
/L+ww5OFhj+jUGrGbuHn8F2h/rdASAS5SHlq5ge63lexn+TTQyjp1zPjXV75+5iy
u2Epls3lCuLMC/5yI8QGAwYKVGBkjpDuXbckWWAfLVe92uAyjSseJkIoLSrzypnG
8ZrrTfmBI9AdNRGwgvrYheM5aXfrkG9JH649vhyCFYPTIxsS9rzOBolJlcOyMlhD
u684nV0LK5KcX3EnEMz/yYyL7Q5nkTfLMLyPL2TJ+xP1WTtuSWiPsH3pb8OtS/la
+f7R6hLpjHZTbWUxjTovwJZI/oE2P4b1A30MkFxlgGH7FEDTMDJFF9YQF7fAHN7V
QPVfP93pI8aQN2QE2ZStkadm0T3LQ5+adOE+NMenrluele6T2GcRRaIclnSunN74
je7hR139PY/tGUaUdzQh13CheiWQPtcDDr5UQXxhuVExNeGJn0hx5vLrm085T/l7
8Wu5MTlSrNNw76/RxZjmtiZJKEsglIm1BmeO8WRmsjaGLUfoGZszxFnNZpjMoWW9
QO3j8Cu++pDbpyiNVQkMHVyMagb7JdM5emw2k7sVpLyMYPesivQneGjb3G9/w7hR
qXpAQV3nMGdmXsiKz2pZuxHhmJzBYDch8vtZAPPDArLb/10YzQgQd//KQC1JM1pG
NVtp+DBjDGPbXzMBXMjzAnbmr07DMzKrWGC9tNnAULJzbuPIK3gN7x2Sdg9janAk
W326i6ICBE+m7Q4v8InnQr2q6dE3sgjDJEBn+CX/mCiTnXJBvsqcvemMLxcQvXnG
L42CLP3O1egHN10TL4JDk5zS04agDrKZTO1nrHYo378s8mPNobgq28KA/SwS6fuP
irgmtYyi1Rw+bI+akW4rjjMgZGj3p09Djt8Dcid6XtItCBYaTWGjGzgRzei5XWfu
BjiItnLDZC3LPslNk/AAcERJ1y7eoy76KpGCAW+zOfsoOU/PWCD1GtEiBDXZwzWz
2teIOdFkWAuHqNZVyz5XAy5oN5bfjO4ieCUNzSpvhIA4LnzeSTScwBosK6LV+8pc
Smw/kKww+TzftDliUVEO3Ypnjnh0uKtZALhs00sEsNdwulW/lb/5FMUOVjeI1SDn
xeUTBfpC8TOseBDx1YgeaKGlDQFHx7MbS0srZD2EFl0FpEo2t9JtI8+Te77USfar
u4ymxX/hPYoZU6jKJKBiqFeT94shXweSq4u2bIBkTnb1Hg/PMgso7AarsbypUzK7
nFwLeNG9VmqZ27u0d9Jx0VWHw2Uoz8EKfCjZaQOfLHJ2cx+uRN/7v3tLC8MkzNJJ
bdExLAUwYcIhFKr2Gj70TxCZWQV4jQGpqIkT7ondc973+X9jvrWO8u68qyDA/Tqa
4rjuBFvk2hZKo/as04V57p8gHW87wZqHoWmsqWfuTsbsTLVNXw4wc44WQtQirFPi
6yz+w2ltsD/BUiMDszJU5IxwtAEiMCTucxFu+YqN3YUz88O6czkyVUr6zgRkUQrb
w7HLkso4C4PxA/FGPMOX9hJm350b1V6H6KUhTzK3G+1xXZNeTvMrktjUIJtncMCg
mlPJ5ursvntUccvoiJLhisoZVTY66/RAUqkCFi3mf+quA1qQHvFLVvS4I4Rh6jQs
dJaEvFFxX+ViHGfX5U6La6nZrqkfPx88sDcRypDG2SWAknGMTTyYL6xsQPMvX/br
PP9LBNe2WWYXKOKoAU9YSFgLIVz+7NCcxLzzy4hwB7pnd7hA/eHnj8lSfsvF39r/
JGvAvoiZW7HcTZ5c5Cucus3+wqnZS3t3U9FKTB3S9udeXqIGNE6Q2zx/GTCfdiWN
j9CyLvsyrFbetObST3JJKlU8S2/AyQm1waOmgd6EiQuapLCTEeQ15ZRHqtLOZ1/w
MYSyd3SyLc35xUIRtHzmMygL+0UPCHJgxYXvsZmB8rtDodMUvLxI+wpWyZnThZsa
TTf9p2n8UYT/it/RkdQxiTqylI1AyFE75kGijmlpCwLBURdh9fojHJBFxt2Erlbq
hSjf3IGKLmZ/K5H9rawYUehvMAxwxLasEGA5ljJ+SYd8867fPANY0u3rhohhlg89
iQfsZe7WQURyicHRXAK+nPbq7rol1CHevPv1VO6HDWt+IPhKXOkNldfwpB7gzsDB
r/G+KWhsBBVX/nWdAVfPchWscsU435aMkmI6rpKfBVaZO0reZAXU5JCUwnU6gwW+
KaUJggOhL+tvrb2IAQqxdr3f0EkjM3e7FpfkTBQSTqb3knI+Tfhn9ArlQTu8JaN1
de94GNAvIt9xyYOrCZ8tgoFeoRzjGI/z4nLzjT2B3GGHRO0IojGjPFnIa6usYD0d
NYSM6e1HE64tymeuWpinXq8ANTW5VRFoCGfv6cM9cndVCJByx/6nK40HQDlSlAiy
jmM4VtXIA+1syO0n/8cvOD4ZM+tgsBbM2zA6kQuB2fZtLhER8Lfzqa6XxsGfqnZB
MX4t/7h0tkhl8jyAbu/mCpNR/PDgBbInovsC3WksKAPza35nPHwaz3qYqYyAF99M
Yw+YZojGLVH0b154MLoHUnbrMRVhZHvCTaoaFk+ckJ4ScWcOhqe9paQVjO6qc4u8
wT2ikAq3RbupWjXCRQBbqg8cuMiaTaSiQWrhP5oIhas25PYzEDJNrz4DunloW/XJ
ch4meHPPzKyvSQqX8EU5mHRunjlDnmBBGQ83t7MocKRxvhlVk3CoShpJMmieSz1C
aOjadjxqnhqJakL6a32k8U0efMXARQc+yKkDN5Bglb3/X2UZwWk4gCxs8yEgP12h
3x1ybw2s42aSLd3jb9k6RKqWxgW2JKiC4iH3JpirpIgzBP5ALjvnQ/1RRAJiFmsA
YzmJ38/A41uirVZ0gzwEq30Heg2SoY0E9VY6df5kWsDozHRgN83GKRrWX8/4JmnU
D3j9FXnVltfGzAA2RFwOblWrTIx7b0agxUVvAfazN9VVf7sOPeFxkdvUi+4cLChz
5VkvR29wR3dI0Ki5c6YzEM8UugJzQS5Ss0/MhSHSmgv6GALuuhwSJa2/vy1UG5cv
1dZApsNO9Ph3W2fPlUfkzaMFSGdXWZolM2NmODkRrK0USIe+AR+ToV/1pY69l33s
BE0eZpBU7BgQ+QNCpPTUoCB+leGCzqCK6bDBxTUstDiM8bPQYTUc02q8ssBSn0rI
GObCyeYCVABLcPCDQcpqlr2zz1JgOOXCdPifKsB6RAHKfCE/NMp0veYwYbAcQRDO
5w2oAGiKmrKkW6QBHBaWf66YHt+rT3xFVLQ8HQheOjTDuGnq3bbzW/JH/QMjTR6M
cQSFgKSdHXoqA+gBqU2Y2N1yjvNXfqKA1iaCsarytmaONstFoi7CVzXBI2gNtX3D
IDTF1r8cJbf4wQsqrK58YY/Ic0/ptkc++/fKeQu41TcUwDfiS4QWCvVPGGTpW5XZ
OPZueXX/OTpHUew77nJ938+iDZ97y/JZuXOHEfPRnPjOluPIVMd0Tv3keFZuGlSp
dKrGuJk9JG9EJmGbHbGI49hN6wotdMvrNWsioM2z6DJvwSP3Cc6uYErPYSQKGDiU
BhPRRl8u0Cam5eE9D+KZHsY0PKEB2lg/N78UofR/k1+QjN6rRd+Cw8lSpXVqZAfT
W8IqTjKqhZIRhacZDStCieFvWvq5C+XT3AK4fzH6fI6gC1DdhCW+O7jMa8mPgsvU
BXz+BVpRMqA6H/qJo/idRgJ/ASOFe9SY34FnoIBv6LlGU+3ERzFbTWTQFrtHkfW7
+X5WdPBo27WNZ3p5+hmWlID/JJYCU1yQRpftsSQ3uhd9bbtvTmpT7pIHtSHixizk
LG3iUsAqweJCr1QyaMbr63Xx4WT97u2L0IL3uAfM0YsOVt5Sv5hwcbH9JGnV39dp
04WCSb8m6rV8ZQky7eKwNT4OQPrgM9wMgHD6rDdIh8h2nJQmT0nMj4EkCv90rBR8
6rq66T41gvx4NVFhncIoakhoy+JbR6emKZYXx+YK+gMM6pChcWd9OtXNB3xWfRZs
qJLJhloN/R7DqH+2kh+31ROyDrhuJ1hBEoGhrppe0S0nEpeP52aYLNQ7qT7ec0CL
VHqAVYIyjOoCN0TewZxmE/ebXGcI+z5I2VdvfXuet7ijuE8rlgxpHtg2nHrHbasq
QaRwhY61m/c51FMqkChnHIhSGwNPn0j8ncbQYOJ0dIMXzkSrK1p74fCZT1j0/zQU
3vW6VmwxVTBQnx5uqnPcfbI8mlaf4TW7HEohnhsP4c1ocGdTeAH80hAyomb/imtz
ztdaDCJwKzHt/YwS4SaWaNXatFybfZ0xXoxFW8+WvIQKcFHkaixGzwqweaJ5NNx8
zWS0cyKS+NgCPtJNv61HQ3/b83+Xv2XDFjacZloOe+mc2T/lxYoIzfJONv2iioJv
Y97hi4yrYcX1JW6t4X6un3li/p797/48PJL6z3lVoIvmyzAEpoQWR0yd+6QJF0um
mK+/GxEuCKasYXmISMgYRNO28Lr1xPGusklScpffTptIBPQLuLuBSye5yCyzkHxm
mxy51S5aITD5hS9V8epOZJURoNO8Tto8j72iM+2eGiI0JhxrrvOTq0yowm8b1BNi
MRUBTLbEHeJ3PDcgZF9ehOFvUZI+XCnh5fnOHdGtAi+TyWhPKTTZDMlxhhJgGddR
WPabzG4O3EIAgGVzNrLwXu9sEn3iD4VEMOinaQayuLBu+n3NiTbh9/AoD57FT1kd
WJ2Z0O74wIp1etwnfjT/fzfGqN4XM4+Vs3yXWNl63dVKWvtTcdI31ogiIfAEXRsK
DSd9vCFdvmC1BMx0tRXz5Wx+5ezw78TBFzX1GE/P4UwE/Q8L9wJlH7RFCRXyk2IF
Xjo7ugGXG3zEHz/krhWSq6OjfQJsggvnFHh9ohynLR8+rK9foUjddNVxKH5kzX2Z
RfM5DaQphcY6jsaNSs8/cHinSJq7JQ74TF6SA4KWQByH+6eFwxUuZYg9miFupvn8
E8e8RlrEHtxXein50Vn5Iq31Xdf4PO/mWKdD2XszjVCCz3OagIYjis3CqbWtWcbS
vXpFKcyBgJvjcPZeOUhvEyPoaiep3IUaCTE8A7YTDfYe41k2rl5MUcH7gdIv4Um/
SWZ0YBksVAZ9mkffhQUsYRuzZPY8B2qxv4lGiKWmIZTSeFqlb0YmlU1thwcKBB0+
a64uo4aK77xUWV8hrqvqvyMb/WT+9b816dSO2dOFj75p9LEQPyZrlH5S1J/8ZAMA
BM0ShsXtPdgcoO45DbqvQ5E+rmDzT80UMx7jYWEf9sfKrPX0flJzLlDY/g36S6iJ
x4kil07C6F6qTgFTT5Zgkh1PalcqG+uKgM70LPGet28nLI528QygSv/IfiL3sBn1
AuifAAjJbpSAixLMKF7Il+Jd+OyQkShd2Se9P5sc1t0teZk6FfB7oIzXkWBni4w3
SXTwDWSKtxFJ8FXIEU09a2POaIIgDlGBkqaIUTpShRLmdraWRX/WO6wMxuAiGMjR
izajyARbOX/BtQzSuxms0YUo2CN8haByhFUewEaBhwWzt1MTaxjiDAmyouNzcbOe
AlvDEm231ijuz6yOUdY9/lHu5Cz4dPok0zujsOfYZUtd3TqJg7h1x0RbGGGIzniO
6eK8JLV7Kmb8HFt0Ag09G9P3YJWb26668nZZ1knNa0Kcs3XN5JmPvvkvtLz0ywT3
/E5/r1JC0GfVIXeKcxUI1a3r1UmOWdyqQYKreExAjp2UwnB/SCbvFwfULbPKTt4X
uSp0RK1wJNtSrFPKGN5Rl2XXZvEegSG9wx/v7wUvFbPWJ5jUoTVlYB4fHZm5pCan
e4yTJ86GvoW7AfuBYhYF4aOWG9seKzA3pB65z5PTVppGxtVwPEvAjGX9/8M7AQAp
LaAqhsv1VXcT84XZDRTXovs3+rXNeE6HTHruR01Dce1MIJkfx5V4tOYzfZESI2d3
+k3NwOFe00hyfk2r0Hru3FCgphgP9ErY2XDLLvWpeRwZVR6sBYK++3Yy5heye0vk
1KeC5Y+tLtlbCbReVL97aU4BlgUS9hUaJI/LfYGMZD671RA6NVPdETZo0iObDkqU
YsQUgSCzH1/fqzAIBBC3wZr/X6AJVqLt300FfwTvv+tOdmkLsK2VHOAyOiutuzn8
9vtJoHb6tmP7TGi9DHPbnJdXFAGBprz7mRMFNbvGpep4mjBXpfeJ7c7bqbuabeCG
s9CRQVxr79WnMReSpXK6gOw1A4mEyOZbdMYldrtItxMbeu3VW4Dgi452bgT4xL9P
o244QY5a8gaN+6v5yZsrbQTfCUg1qGvLsQujGSoF+XH/QEx60vpYeBJa1hZhyorM
jlcxB0v2e4hwBoSKzPSN/k/NhO/wljEuRFDGB9cwDsq/iJrzaHZaPGK26eNmbUHc
bGHDAmVUcBv5rBDC18nYrIYxz90ykZ3dCtiYXGTetORgNFZfaGDfuNhPRDec0ouI
HpUy2OCAszY+lofZ2QVt/PzxiKf6in+ADvaOxa4zwxiabKI5GGKChPZWnkXK3urq
/qKsZl4UYmAep2O4j0w5F+aBEJO+JI6wuxI5JsC+AL2AODRlY7Ex4wbJThnnxAWu
CdxKUSH11ULFJT66JFYdpprgTBIbngC8zz9x1JJ6JvWK3ev7FA9x9elE7kk9bl2s
Eps9f1tSV0CWMEIGV0Zmc5vMVpU8OmCk8aAOwc+WrNtwWCK/Ik/fKf5NHajO3xd9
xKryM/xi45YOLO1/5uO5tLkJFPW9T0ycVDBFQyjPRgo0pwInhTRUo1U6wy5WrtWK
ILcRe4xkpMPTCsyXDvyo5MqZ1iW8uI31vqS5XdqSeuSPKYUNkM5BlPcMOSC8bYlZ
ITI3LizzWvKg2ykz4qe4xvIsldC18GUNfKGVdOAPAS8cSOjnKz42It8zvGrda1vR
E5J4uRuZNnTlDyYKj1HuPfOIGk5Vabf15A5Y7/jzg0M2nD5DpyIHT1d1uewzdSCE
KB3gZxmmabVHxzwK6UgM95/eRxHIrcQxZVLsdEskkpwpZQ5jP8MDUNxWJStqejja
7OReRmkqyegk3vh2sEM1E3NAMBt6UChX67yH5rOBUlo62xD13aJ6ODIgR5Ku9I1j
QJYwbxGW0UMIbsSFrXGszV9oyKE0bBdTZ/4D5xxXSpvQeVJj8CL5pIIyY6k2NPw5
XxfyQEZ3JXzasB9ihyF7Sdsy+1/pzC7NyxRvsGFF7hloNkZ1X6Wz9SSUalOi7ztx
bqRvbhhFEIWtcRWK0mPgHBPXzeVDhwooz91UYqWvR6VD5m+TEc8tJsCxDZmv9GbQ
TKolygW3TTTnXUsmhGatU0UVflFJ0ikM9p7scdwnYoWUEHLBnNkGPYBTQRkksO3h
QhIpmNDN0B6Rqe1eYOH8bxCJSx3wCj2wkaj47rsi06j7dPYcQNVHuVNoIa88PfQY
P0i7LYMyqY6ocsxITiP2qIvI/gTNcQvxkwzI0To8MU/PA/xEUnXJDTcabKY1qyXI
YTat5WAsuJNf0DDcm9VMeIbGc7Am+rX/1JFyGxdPxtMvlgrrJMBuBs4vCE4x4T3C
yBG3gY3VOtPeIIQ3A9YX3C0kuOUfGw0gioqFl9R6f3BCPt2jOu5hDEKM1G2uPZhG
2dpCEDQp3Q61+MRhPzrk+qGACYODt6TIQOiU2i6CRGWnyVfoha56CuZmkfEkKcJ4
7JGS5pE3ZzyGwQWkgy2ANFoJV5pfoodYT9Sa2TO/MEg9fXkgAYWzWtyEVqNVjsmT
Lz8ZSSkEAYELsQHC9HVDoR1duLD0gi/8OwymLv9/lHYsZqceEVnXIrwCjycyDQ5K
jmmPBeKXZUVRouVCmh20WO6soUNJQ61Ha1H3V0Yn8yLFaMTITEPdBE+8W/80sOWg
gaDKehPm3tLSPQvPsiWbD6N5VXRLsTErDDJ8l1B0tDpMcifAK4XxcanC9CisuTDp
R/vwinMABxQkKitavJ+yrfn/mglzQrUqU/KmVGrJjbi/zcAqqQPnXhcDpfzY2Ulp
XcPknxs72gpmauFNdTfxSLI19b7SvKuZDIW8Sd2gGSlYI8td4MKZm3omnSW/4t8L
WnFQc0HqDHTgK0m04sjbJRTurxMmsbWLpmp9SNBDscT9Z/5zoH4OcY0JX9wKoko0
ycu94wkMtCmUbgwSeGwX0i068jqnyxrEDWOstdD/aCPeO/UjEzDCryXjzZNy+v+N
UzXBnUK4onSoiii3f0NQaFohUJdMkII+RJQ59zRVWSzgRP84FIQ8LyZ7k2RTDzDY
Np+iBJRrmlH7fs2mYWTtxqrS19VhPEfrQo3HPykH9h2ZRdgrvJsi8/p9NjEuuWoC
s3U81luvg/asVBjl6woVNntdgeUoETIHVyztf9T+zDVQNVxm9t5rwSt0TlULGnYm
YzvU3kk7Y1Ac0qgucOCWWOjS6CBboqgr3HCPAIvdzP6nJKqVh75MrYHjfWm4J5JH
nP/iJPBYECBPVMTX54CN/TKSXFqq057lye25C1P05IJCYAqL5LM9UfAMM60psDsl
NV8l7g4LZc3/cTyOxm3yeqvS8SHO8VOqtqwVFAWiLay14Rx9SvPtDDZPnbpFovlW
H0Bjf0ojwOQ+p6ihYUn7lLcDhVYp6s9ODa0mLxFkIKOIeKWZ0bw597Vqm0v69yDx
V7gVRS9RBh35xRDobAB9C+kNfRv81AN0HH+hzM7g3RYqvDZj1ZzduZ5zs2lSopLh
qJPsmCXYwIBg0jVW1RA4uR5Bn/MnzoMwekDPYA6QWZ3+MCBj7QdO9ZBxjH/nA7O3
upzD33szYV9ma60RBToLBGt61kHkyPdwBA04GPI01VWHubWrz+LGxrHhwvLdI0R/
pyYN8IylvAka1BqFZlSTf2xMrGbQpxRuY2FWnX7ey2qJNLDXhItFAOwHmufV6m5d
MT7LsOwOEj4ZMROWLK7i1kMh1+tLFzCZGwSDWyqbPR+9acClDaNAH1jkNW/wemc9
uuoqscfkRrvfp5/deoa5Ny0vK6R/jM29+pP88loxbumh17eI4ofK+DZ71B8zT+ie
7jQSnERugOazKYd8Jb/geu9ltI525rFf35Tk60JDhiADHzYYNXvJ08JsHlEcEuWJ
7ydkistjZXrM24yq5jTbyi9+IVi8LteRSKWu8Q9XO2CDTlj3VKFxGJ4KRTU22Vtn
DKI0QB3sjW6xJOLgNXpJ3PllJtX9Ar/cbQOUz3XNvcJvgsxO1xZDpUMGEpTKD3n4
rWp2xej7yIbLOrZSoygooWnN65PM8HHxZyWglPr22dd1fJOkXmhMM6z1GqRy1Mqd
RFfbYw7K1FAjrQCsK3cj/tXdh8o0GP6IJ5c3+htSOqyqWR2LdIeR8u+UNWOp5K0Y
VYqPQ6xzbquzZHWD8ynq+TNqCdR7GrjGwcNhfEogQ/3IOdwTaMkJzqsIPcBnE5b6
/l4BRZOZuxaI9LSx+lrBnxsl/WAmVRKJn/coLTUi8eZCV/K6QGoN8cwMNrph2qav
i7VgGYWiQfF7DoGrA3F2IKeFR1RpjML7fSlQz7wIstXA+QQ2uVyoc41zOQhqsWBh
AdUcVuM+hQfTHnzh5Cub3rT0LvP24J5J0SYEPuLBgL90ZlQo4u33exVhQnsOEe31
nrPA5PrNGG5evwXC4kX6YXUx/pIxJR/6IYfXlhnMkNRKr+rSJD0J1FHD/SbmFm36
wPSICbAstuAn7inl+prWXbyLucIZxwR6Tdg2ph9KluaFmjr6+u85EewbtTCrXuhm
OBTl2wfUrxt7QGlnx4AgNFR9bAWit4wEBnI5P5vdg7GFY4rzYJRaA9Y6q3nlvhiX
DlHVDg7H+fKLNO3k3GY3TYTWNrFiLJFfr/Fdw4DxJvRztUSA98XxYKS7T0NFArTy
LyWCBp3HrSaS3+WtxEQ5We9LFnqLXq46zazY+ZMIy0sTlm+Dmyd3V/EicCmkcXGX
TzRkSGpMyNNFMqm9veKFart04cudGjEzAphPsZkhMQQXuTyE8Sar58STiYBZ3Kv2
dHIoxtSz5iK8zaTnibBhLrrQY+ZSmjg2p+Nb0rFHlkTIaTkRbsoj22J58JT7G1Vr
qD6rUoGY6l5w2GcwxOa2Ap9a/G6u4NVxD79QeN3twVI2JsLwd/xVUsGlx/5No5e+
9o0O34QDixLjAyaL4pFerLDBlWHHQWcIGyjvVCC3U1+hEw9kTaFJOT4zG+pW34fL
WS5EPPNqDgur7RfppWaDeav0/afdZgrpOjpxwqw3SpfeXiCIxj8bWevIdIc19pdS
vXgLwEObxd4ZH8ChYsRXy7yOtYzvXlb5lEgD9WT2lpNAOQxY+095aiPi4r1xGAPU
iXCeovRKZOWzU7yZt4axUPrtY45tPa3OygRG/jChyE4sj79QfhmnqfBO/dGMAO7b
RRwJS5TOULqbMZeijGJpBF9l4WYZYnuBiQQH8A0+9qynlpOdasVPDjGqCQgULf3g
u3Au9lHnDPBVxpMDK+/qzkMg5YUs1u+DIy0eNU1f7/btH33pXmFyrccg66O4IIiX
WE0exrNUJCqftuzsZoXdw302kN46lmSJp2hlL+aRzJnBGXeYCcD38+6GWCSrl/TD
kM2KAt510MnFOyG4H09Se6lv3PYOm/cRK+JHnyge3y/faEPdLew2ErDfOKBA43xt
WDw8k3k0O1W3wNuHuq/NFKBmKPw32RIccOVLglu6XD8Wt3ZNHwNR4OSU9Wrr1Eb+
RctKcl+kLklxSoDq7g7L/SfSAn6KcEGAa8tIYffP+UV4wq6UKczxwR9//PjIi/DN
Mcx30+cRXwCGeoca+3fciaRJ9dfV94vtvWGb8eGhVmxjXQvtZSY9WG2u4iMzsCPp
F+g8iHBSsoqPNx2PSDwzgiTrKQJYo5yBjj0g4CPBMQzK6QhRr5rKXVefpt+C+Xhr
iAQWvwZjd68I8qHLkvBH6nafqsEKLcMAcJ0dw5xDL41J7RhwC1wNyCpG9byb7bZn
mK5vGe8BlcUDVLURv9BmWELJ2zEH6+RZOQxZQri2kHPrnNiwnfJKUUS8pRdN4Gfc
3HEChNO0pkq08eY/jaEZYi7BB4vZnnlWZz5UUAFxEH78NfFc7QrRqMNVGdyZs+mL
nCKJJLddhyuIPqustU7Fbq9505dbvm1upQhioCQaFRwgLNj/c6YyWcHKOgEje9Y+
4ZYhLF1QhXNMjAKj+dVpbf4fjvmfko2q7o8sE0NsudoJbBr712wPXW+VdrtFGUSO
aR7ZLQbYOYyciIWRqk0eihiHnL0g0+ItAn0x4lDSKRbnWFB5eHE5WMbQesnlgMDu
OapcJxglJjYpBhoIb7iPdM7BZ+pM9WAWq5mF7y9VosrQf60xfzJPcXMBnY19v7IZ
hDC82SzP+PiICo4OLq8caESP2AQP24k6Me+BMS/pORWM+20btc5elmTgDDVAVqIi
wewacDoG6bG3F29eEdrBUHex9Ig6BmOaIuona+RukWpf0lrfzdZ0bxXRkaCM8xGX
GVjAXE00oDzCR0o63tJZGNoNOVxHDPtNyc+7qyfPdWc8XQSrd9ZFvp2eLqFLf0Lg
jY2vQGge6v/XdncL7WmMdnqFXgAgpmR6lwdp5oZI1xtIFXJZHdu6t3xsEr17M2SZ
dBocXouA6DqCLiPTXHW+MBSVGEYIEzvbJ2Q1kY1Y+/cIke/kM7XmC9x9W+lDGS20
eyy/rz+25yBDbTvgoikEj4oQtGmEDnaYIRZriAGK7/pOEwc3EEk4GE862S+C7NF+
G4dP2/9nn9D2bfdQpQi3Dc1OIKx/lM35Xm24kKkOOekeneooDs9d+9vI2OTCIR0+
dxmvvHD2mergmjC8F54sAtW54zkbQSRFBrltuvjWBcDZOo8EBMLX2tBk00PbYOF+
UHz735r5Q5fo2ChZvBUy/8INxim/vncvPnia+2BdTAYfvkCG6QoZyI3SNHc0SJlJ
pfZVPac1CqDla0N7ruoC4P5o9iZdCLLqJ18gCuPNWlFs4nkUyo/rfYlkqWHVKQZq
isSZsHWjXKcvsticMtICsVY5nmMzdnmv9Q9ux83/NpCNFTHFP50LE75tNXOuWsTv
HA5Z0yxyCSkU2DiUdYnB4gX+h6t5zCdXHoplXDjovSoc3X0wp6bm95Z1t9DbqDEa
tHnnm6jwYYYlqO1g7GKNULGNi0r624mA8amFMhZniqjceK9dKLqOs9gYjHy2liRq
pxbrHdIfZaQcf48AtUgmbP3xBejat1CW8JKHfw6l+YFWyQGTMDWY+BUPhpI0pp5L
qBkw6UKYp3pUawrt1YTJ3+qYDDO0/u/D5Fq9iJPcx48E/ofb+vAnIRRK+0tXeB1T
xgRCeP7BTPctfoEmHppVBiMsU4CePm/8TTjWKYul/nhIIo2jYuuHqWz2Ae3ig8R4
lTBnJnpOOIDf8rSZw5TjFWc56/QIRF/ol1zse4cOsdJQQBcI0R/mTU2s4nnOCQuP
qN3hw5YEtYi9xLP/CKk5oDEC1Z2mtR+qLwaRxsI2fFmxbF3T6k/US3miw+L/rLyj
UlT0nnmazxu/yeTKqtmIj5DWKgbwHgwTCmxg0gU0tLFAVxq20N2vucSftQ4Ovs+S
rqzrOjxYUTgnypMEJ7ydlx5ifT0Ue2FrSAUXK9CNUERAD2WCKaEe+CgeUfvcBXfp
wNkQDOwmMlPh/29F8/NL1GNsyGgZQQps85EJURzBfJXhSatngTPa/EwQv2ixeBud
cZkfBqZ4IKd6saZRh3OAOLKcJznYdHYf2TMmVYIcvtbmKNIsZcQCsgw/nHFqEke4
rbo57EXHSAFILhs69Lhb5dVWtEwFS8hNY9E1mo23vLP5UgLrNA/JKiXlcNj/OjS2
AND1oX1Mckl5SUaOXwPp/KKYAa6YclNB//nxuDdj/W0Glj1CqJzV9St/74NL5s18
/Z9HsoJ5W6fpYrBGMk/oYZmNfWYBY1hDIo+Utb/m9Ex5BTZa9HseELbXLcYcGD3G
aZdXdB4ZNs4kaSgKlcsEFg4Ojn1uelpw2YszxaK1kJV2YcwjUVsInnnpOjd1W9lm
P2SRS3fPUsFph37qRl0oPuqwgY/yNESjI//iruigqUTV/JBiubJp6I/zoxaSUg7D
55JTwqgKxyLwaNllS/4sQdARbWj3XOcNyPycWgStHx2CufpO+4V+d5m1nri7OzXp
3w/eHR4yButgg/jWlYcnET9rc3Up7neh072X1XLQJ3JdLi96UUSpyS1CdT2Ha45v
Zd5j9D1jWZLo3YgjTho7tYiYHORF5gLeSF0m9ZteNU4kbUtqLgG0ZeK7VHzCk/bv
+8tMaNkw/UKZAyBPNRT6obu8YtywjPI+R5OvJf2jijamtubtVJepkO0IQS9dmXRN
MVNPzNN94rMWutn3bQh3CbUkfysUF5j2G0GKPej3t9XF+C3fuXS82/qfOAd93j2a
VvhQd9G47/mPAV+rbrSLlMVlRC/4Nxr9odN9UY/++LPXPmToomqG29fKQm/JwGYh
uHGuVppIuiHrB4IudgT2PTK/sAux69vcIXQv/g/1KNOPZjopTU6V8URZ9/wUY7aO
pVRg63XJOCkscXcsOg9UAqA2WZo9HW48EWMIABsdT9K3Oz9EYrLreSJJhJOp5OHH
OJ+Mk9Ot/qwOyNs+e4HSl2LsUdeQ5rH6OCB80QbwsahvuhNMrJMghLLYCpQhwbAZ
MrKhlLJKAcZAiX1DOnpUyUCgj7iHO+rCk6KsDBTORvO7X3MhwPEpZkaUr1kRGq7z
b0VN3koLp+g19UAICmO9dkJxPhBQ5vH69enasIY0CrqfHXgLUrRGCnUbzK8Yjbpo
/GRanNEkhqqoRY7fhswuG3K/b7+qUJf1AHvnBedr8BBDy8764n7QKhT/CXRva8QE
VEwzqqaQOmafymXzBxAlfDL4URHBJFeFQCaqtTxAnUzb1V1J5uSnrzvsY53V5r7c
9oLf3LcOkAcruA8vQsArFvXcUIHnm7KHX7lsTda3ODh03w0o1NYSXHALQHaPuRmW
qXnmgdkqSZ18WkIsnLRaVaipO91vSU0CSLFMPHN5S8VctbcaOwuzMUVXx/7PoOjj
KLl9Va7lqh9l4HTmX5BTQKjs+aPSQWMPX0+dDVuKxEnIfj3rkkYoK5hUt3oTp4Hw
O0Z1aVJXiQRqEzCe0eoHRZ2ejv5WBhJweMyRy5rttKStIF+t5t5x+UbPzfRyaVy4
MxWrvsQgPUBG19J48o3XjXhQlMJ2P7L2J5RMgysnhhGHZ3ZOn+IkqqxvM1dGo1a3
RnAsab0QLnjCN1lKsoDM3G2c9Kl5SUl27OHNWY0SyOtrtNkTrIP7avbamA2VkCbC
BfZYR7aZewmfnnHyB2lm0SOd6pSP3mGbGruwBnE9zPt61QHZu59MDhNifVEXFmbB
MZKsYV9JUwg4w5joirCE+IQqZYsnHeF6e3F1k0g+6uo7AKiJYo5ajQ/pi30VFrAy
JCgFWgaF3Okw9Is662WigG1RMJ0zuvxi2vQGrcUPY6ATXRLtYRLjvlgEJ/d5JNL7
OGRMWge3+xoAg9wQ3BCBSetm7X4JvYvIt8kuJAyicBZUQfi688Jx2odO0Xqykfc7
gXOgeLcyr92tTb0PXeo9JdovEuYVIOhHIfCqV1zmO6k7zGFeWgyckiZmIgG2EaFN
hJv/wfKvU0gaMn3KQkebk/SQjEHqcoWVND3BlMDsSLq7c+iQHDkDRAHhwRzEjc45
R6CsBN2sy3thhrgqkGv3HazU+/rkqSQZHPqVTnKZkFWVimTPzzJf1DZ27T4XHTi5
7Wo0+6RKWyfDCL61H2uyO1jS0cP38EMkT0y6rp06tWskdiNucWZcLhetfekpg1PO
qckS63XRU+UwZGpDnpYezF8BcuAJ77XVn6Zs9i2ElQmxVdZcewN04eEA+Nwd2tpP
jNQHIKg4Cr6jTc9WdEsr2y8X93nyLPqLs+J0CAvjQ/guRpIfuOrTqILuwFII/Brm
sjDGcTzMr3TgNL/ri1rAWZiuk6eqY91a5vAa1kCxYn30Gx0VXrPQsGzrdiIusFwd
fROuIlQl1oWXBHvpaJgl6ft6XAqdTJLTmtY89+p4apLRjXmj3ARS3d9HUYyRaVMe
HKsPoC6Xue/CGwnEElB/IdTbwFuBW4aIJMVHBFjjvVGtI+uzEdrcuzi0S4LTzYpn
3dTW0oLByUk5ARPWXQv0chHLlkzTmtUUl4CanG98hQRgKHQ6Ue2BFKpB6hDBerc9
B3Qo4IdUASxq0fSTIOOu6LV0ySJW5odVv0lfFEkHjn84BGUc2xGzLnpC59HZe/Lt
mVRieBAc4EanKTd4h3a4U78U1PRJaW7p+A53Z0MuomSFi2unkeRcGAXZv/o5o31s
Myj1GtTCMM0YcExzQdtz7TpQgHGKAI1J21M4QhlODChutXSDE6t4WfnwmQZxOJT9
xKS2LVQwP006LQ2g0YxYrMeNWIL7a5Ky6X1DbXp24qrxzd6kSXNTEBx5tmY2Ugia
viGsOzM0XTBNigWOnF619kek8aHyhWrYl6E3Ok/HM/WFSWxu7D4V0wSbmcmi3+HW
E0pCB7dNVFHG70zl8FcI7tFtnT8GA+AUajgrtvicmLIwU3z0e1kWY7pxbGKJj9fQ
YdOAy1Tu8jsVvacnKgWhWKqomQNkM8u5nIuqQIWNvSHcJo4l3sWHczPnFkYQu6c1
E39md7V8/h5YZUfKPWTcXnN0VnfcvIiewRdPR10S+gSTgIT6njVyMK7YCt3Owv9x
XP39A1wxe2CynNZCVxBtWKOGRw0QbZwZ7vLqlCuvuTd6o00liRpMD1gqgY50rhdY
hfLHMgAdCYgPt2/uCX+HV8OWzyrAgfk8piVZyh2zFYRexnPVpqORc4J29pXB0cEB
yoZd5cWDBJ07FbExfsDbIfWhfexZlyUJ8CaRQ7p0HhnwsRcUqoLNB6WaFtZt3nrt
6qxOyePkrtWshuJrXeRxcvdHDwZ2qlmbIMpmktwMETq1Z1ELaKHkbk83IkJkiYDA
2FJ1O/uom0Qq74P/fxIg0G7YkpZySvM5/5x1/ZetMWJNv15uJEmtVq/2sNC32WJ9
LkHNyozA04lkX0O2OFN8DVbG/bHNnZoEBDvl2H2r6pNwoVM2hvf+bkrFMcBIDKzB
NwT+/hl5t3JD8HEXHam5Q6WuZ+Y1AdkipG/Ri3I5a+sA3qlj4wpPJRbAyMnet840
CF6kfDDziw45uWAmtaMLqvMMBeuzVgqgj4qEWzTCLmZ/AV9Ln5GL8eUpjb9/A45A
hK9ROp4bHMFKpSjnIZ1Hgt/Wqx2rJlcdyawytwmURnoCOWmNqkhcEfV8e8PhWEsn
lpkM78VBXWUPPTW0l+h8NUzvL7TFMjfCpJWwqCEGJ4j+G1EzbIwmL04UgIaivj31
YBk/w4W+EPaolpxaBeMmWdzRcpwIW1KxKo7OytWZD0H/z4v7od4uZlHZwkeA04TZ
8efUS0a2W6vEdsVPYCGGsrmj4YEKrZQXL/nwVgVgU7Du7c8Gcn01Wrih6igR0L+a
lWJPJtqE30C2u8BNkvQksszr94/5YeuhOFDaeJLF8j2qgLgvPUAdRZ0D810x6cdC
7jEvCKZnjoNdkjlFndNGaLG1SOm3Ss58O8NUPVc17cYB+ONRFYOOGuwGsVavRbf6
NN0PGA4CPs+TnxxBcS8X8dt72I7tZeOMTVzB+eVte5BLcknkyfGb7V4MKlEZdkw2
BErKmmI+3Zfdz0YnBJcdItWzMStDrG0KqRV+VmrrBGmAW2CEIaWUGtTW0eznyTUx
+CnINPTkfjdpmWxEs2wxdxQjVZb9c+gsiyjlPvHxNKyg2nKUV+oyqDuA4NytHJn4
WbQecn+JiBLgH/RZc9Bqhc8sJUDbI9+XflScEL0tag5jN78BAF8N2V7POZPpKJzG
KpVztGRcpJKAvJ+LBXzsPrWLcW4bwpCFjKEENahOwF+h8V4wXkZhpvd7ZDtCFajF
eqtkdJWQfFJEcPnmrbOqfO6jhUIP9a52cgSP0FDLwOMRbpnB++ogckaXuupGDhoG
ketFjzH9p1MMrleHBTm5v6tEPwi6fdYsPuxs/41JIl0Ku24C36njaJAKm/AzrzZg
zHeEvUAW3v5TR9E46Qdvyyz3boKaxUHidRhX7m5kiNd/Dovu3i0WCRdhKlKPtE66
gmlRFVDLY+uAUkFViHVv/ZGQmLjCt1/4fy6hVgKphdssR1jo4JIA6cybYvc7LnYD
vm5Bwm36crr1W+GEu0URTQcygcB4KGAy+XARtcP78gCh7ieuHA982Y8rZB7NrG5e
wGd3Wh2HSoUzUUif3b8McaT7+tCYNexdvqcMf0vPzR+xwnbUMzMGsIdPvCIUrXfC
1sEIC3IW+85rpQJ1IXsClF1hQM3vOJTDq7qqX4eGBVddipW9W8KFcsLkQRkRB3Ko
D1yI6nYHYrOnZqojcWFafx1xeh7PAGHovkyIBsU3DsCVCklevVR0yBg5O5p3GsWk
4wCCeam7TQZ4mgIRz8gVoY/a7/O5CCytihjiBr6ntpPW04l1Qo+Y8AqWiFpkVeqm
UlbH2teYTHUKJO+T5P5NccxqeJaepZ+eVlknkTQharkNDUgrPMb45hDo3e5GonYK
tGAXcPDayDb7ICHu79qOoOSUMF3hu1jCFoFY9lqAYtNi8bFlZt2+CryiTEmYG+fR
5yGah71F9Gpns9nJKwGnp+7bD+ZsdWaTl0J8n4nEwWtTWIlvsNL4N4+zkvbsLtm3
Ra/v4eHN9x05S81qhji2qjSo4MiUO2t8EXXs74p6E8OwvLCuMSi0VkCKoxVHxnQb
GVv4cAh+TTjngKUhifBKWrgY03myGavvgULKVAdxAhm4niY+jHStU5elAJwYo5Y+
PTx42TLXM64kL2G0JIluSGPLfFw0KK42LG4krL4ZNOm781+J2DkXsjaYhAGTorq4
6hEuMznVJERiLkfb+7M52AOoSk193jfuDUeCQGgHNFoceYkD8YBYJPFYjdNVUgwb
ctQeCJ+TBMYbixaLX6aofXzrSe0xPDhx7kffuIjjCyrFAf8haz4ASrS5nzcdHrk9
qGUAxLVRZmoBekgFjCbe4ENXi6Wof+bBPpO6F3PRY6+GhDUO77msvGhbc2oziefD
mIWAMWXci01J3akG/aLtaZiI7OX5KZ6ziNcGSEOjcm29B3kJT5kzqhqxzxrQT7TO
SrADBMyWO3/AKV+LBTMVHSHjVRpT/M7s0pTqtJLzYfbWQyIuYQkoo811YvcvA8sj
DYCOxp9OD5Udt38biZYupFTQmh+a6OR6jfZHoCDBzQfpLfLlofXamkE0n/M57Dzc
mZryjtGmyJGyU22OI72mEjJFapSgorNrndVBIxnMKUe2KGjuxYp+SK23jqiqGrmK
CmchdC65RY8xWwBohiHT3Mkc3ZCmkin127LOzi5lcNioQDmduQEDDbH/3J7SOlWN
ijBgCvqSvDjZ4Ho/Jiu8RUf5NZxQxvgL+yak3IlnxRHLMfUFoC8OzJktpFjxg38J
pcaV2PJ9RXexnR43vQsRXFtWUC7nWkbO0w3wiroHETlqX1738eqy4HPa1aZSE18l
d+MTPkETxwaxX7oSRbf6qafx3GfPo+pnCas2ELIqXiz9saqbhd3h6GQoIRbla83D
lMxVEwcHPUiwKcM/ZkU8y/Zwe35zZD0AmsT0CebbL5i8Ym0Sd9lT9M81tWjk3mKn
HJ5fGF67GrmQslEbgegX92Unzdyw5KCaVOv6Sxb4jsS4sqcjOZF9gO/2eYROuBvx
00HhRMgjcLbl1RBPhxqrQfmbEKKQNGDUKxLZKmu8gvK5vsHsjTvVckY24Wuk4n3u
IwN3TdT/Luq+3DOZ/U+9QjivaJNFaA/FSHaESZPirC/C6uVSVn5n1xsM7ZO+cuTK
Cne7HrsVh2s7E/7czzB1+yCTsOW7w8zyFQPIsxTsgthvQoidBmIrqPRlW9JRZd2n
6SxWccTg/IYpNavqYx1Gob2Z8HUh1N2V+nl9TT1WDXKq0w//y4256yncLU2rXcHV
xLmbEXrcjgbS3VKhy2ZyP199qWLgw5l3VN+AachzqLkrOEtqkrpfBVAOYwuGazdC
0V7NbE/CQ97+mzn4/e2M+U0IpN0s8/YiW69fx3WLF9fkg10m6HlCPEzGOChyAuqM
xOuVylZ/V2ptxR0D5sIdRas6vgsU7Nq36bYAp6FMCHEZJ8ER7fXPDQKVHkelbWfA
g+b04SUoHmTYzczc8QMDzXHDWRuRZ9I3fgK/AeDzFFtegfO+qn5rX+L9+fXJZvbE
3tlUSt3mOo2H0dMGghBUsi80MJkxYsHBE/VS1LdBihu5eLa9JGjeqQbUV1L1uYJt
E2DezDRM4MyFL0kHi+rInP2XZgCSp4WInrMmQvSTTiYxhdhvI3ji8hqVKrO4I64m
sjdpSaS+bq1lv7GwEzCabWixicLobiba4uYsLKzAtutVdFEfJY44EIrjW7nHJoM8
H8CNulNqzJuHL92QSGpwlu9K5fZiS7SpWeI/AFYaTARiJoFeh3z1+xshnKSTA9I5
p/sRNyElratwm5LcLFquaIOcBKitH0bjYVHK/kza/dcEOmpVyLZUAUOK+7xhyio8
dRrQcOUo1KOgn+eoU2ovmASiv/BhR8Dv7knQ5ch4RbB7+QF9Q5xcJK6Zml2m0Blq
oyt+17RSbtPJKNlpI+RXABC9DCe/J1TXGKProXkoztZ+lZWMAc4fFYnQOG7egqan
Zh/3EZKVmtOrvFVURdF9FF8hnn9oALCj+1/4f5n/QvlIg0rjYkF/AZK2ZZa/Z0Sq
yYUeWDxAFpCRDzJIDdsMtDo64Wk+ZvidhnNN6vqXYNRWFkF6nHcBiOcp8vv3m1rH
t1nZ+zeHA8QcgfgZ5R2Ym+hneolzggigwAAnZ8BG6psikXsWdAsC7PtsyzdI1wcC
+78fbEo8iRBBdGFbQsLpDSj9V1ZrpAoYSWDYCkcggCwebc+ybNahKdBviArnHQDg
42UVHlnslyFKUx8QU/EI5RGPVL7Ze5CaKz5dsAxVvrj8PCcq9vnqzIJ0Z8NgfAZL
0L3BiXoPENK/Z2Q6vjVtNBgvwQN0Juxxr3GA9eY/I0mhi6lu4jWrqYmmtwbudmyS
pXveJkRa2sa+JG77yafM4dt9YigM4nOGj00XVWdNQFM4uKnANtsWqI9l36AiMQXa
KhNmtkRQf1yCJOSYwF36IqgMz/3vOVWfZaPSTnwA5kFi+ccFAi6+tGp3COAFeT+4
QcYDsl91MroKMYIZLAeeh5ziH+ywdsgJdQanv1vEJ4/gF8NJH7SGW4jePv8GXon8
ahsx1J/W1g7WWPJCr6v81ODvrHqm1gBXVdSXd2E1FYlQ+1mjAHN+j2ui8Pm0iLXu
WdACcwaoWSszy4QUflLItaZpEeCv0k+5EaZ6kJhSSGM17ho7raf/ToTvOQJjsNPP
VL6u9RErBODl5+offJrfPxuriBRDC1Yld7/c9esb+Z32Ei59TUnrqS4lzL7DM0Fi
/ecEa6S+RftJa82rORsa9GoKx6+S6AOdp9WkgeRK/pzT16j3YzzjW0SyrK/LVbFA
EK0NgybAp7McwyVRbNgFSfig3FNY5fCLTG87f/bEnJnkeSjjQ80A15GWkOS3+4f3
jAUSgEcwKDrvInzeWY/rYgn7o5GCdbfpD8NmTnPor2UOB0f0QE/0O9RA0zCtZxCN
jmq3BEVpSWvLYuMVOYk+QfBaQuNu+OW+0Awyz6VELfL/ZwLAjVy/zceiIsFVFqUu
JMGlxE/ET7o05OMu85dJhs5RkXwbWxGkWCm+lOdpLbl72Ks92oXXENCmZ9sxifay
IlssxkoaMIWVg8yUKovy8wkrWFLRJ3pwFeEVi8NC5vO/guIp3WGkt1h7l+e9uVV1
W4fcGOutesiCqG7fOqn9MbYMwxzN2bv20OUTyjGeR61/4UXeReFSZ3yIrMymBDWX
xu7KxNHeRgjAdJxAFogmYUvSh2Moa88y6Yy0VL+wTmaOsgkK5w/nTAqkFEZrvmHj
9y9ERQ9PkcCVoEjCacYLW788nDP3BijvRX5eqxXl3SNg1gOQuvM7potYGcp77DhP
zqRWN9Zw9KZxQx3U9h0wDDp/uR34lIt7/RsF7PIGF+M5NBTtAHooYRar0QMl1VEu
ym9NLag03M6cNSeSnBMf4wEuyIk75Oa9UmdEsAjse9D3yBIY0UYjReQ8bq1U4v3a
ui1s6F8XKP2BLS96KSitxnj+CiTUoxybHIeicYw6IFwnMopu7+9dR3/tKVCEOXPc
wMlgA61gJRRXkEZVkQPyO1VzYYUScGjjOsoc+skIoHX52czQ2LWGoO1LZfHve5B/
PgXtRLX8e3aY/IGZaLRItmkKDbskew1FEnU7QmMtMLOGsboKeBnOCxfHcBEXFywe
o6D0U50dVZ9VsUs2cQYh8I6d1sNAw8x5utE7XFqI0BmR/RvSILjD+wMsNcId2RiQ
gj2z1BhVeKgZsZCIz1LCYmaAofeIAgINRFn3GV4IEyEdK7tLenBl4Sj8ZmlCrruJ
w5bvuwGtoXCdkYQzeqe3ZsU6Xdye/BexyeWmTkwqL0vXb0WEJS6K8wZ9dtSdhc0E
Kti20qQIFyEZgJdD02NQP4nQx8yHXe1XmEBeP42N7FR+Tr5Jey5oLXEfx2G8qzak
EdvUhUnuQjSVLLDE7MU7bNwd4dBJRijyWTU3QNw325fEtB2PGKCQZrJaYgNSs1mu
poDNCdh6lr6/nh8f8mbEl2Sqp8JRsl2XwwnXmnT6ALjpkjNpY8zB8sa33D50Ougo
VQmjLAxaL29ybmUA10jG3m3yT3A8uW2ZkloTMq+Hsss7zptaPcwzJX8Hjua7F35b
1Vh/eqfqeGjwTR8eCRP+UuFu9aMgBjx2lzamPlCcHYhxk3KDiFO1UGvu0geBK+Fz
243wwHDXoF4NJnOdEtNSJQoBjZMi+n7Rk7MS6PaHRRMl6XbohPtrZSCKFhA8BMPP
EBDpFH3EUKjKxkEEOC0T0/df2OOxC51otHq6kkFFQSFGycnt7E7ARDWWBt7sCp/W
ojI2PkI0Rr7EWyf3xB/aHzFraCP5gNoXytZwcmOaRoZERyZKb6cdDm+oHJbLhPeY
UYsRdAgyiEdAPoKTf50jklB7H1YXj0YpCCv+cLvBNk8Z7+XEXmLtaopO/HfjcmEG
dT8us5SvyCdRiQm6Jx75A2jXslLWUJoMjOl4166aeGy26ZwCkfrvet4VQSTvc/2x
nEtxUToEdhTf1GLq/UMLk24DAEN8qCGPgZg4vLBN8+68vWi6XWJAmUT/fpRKbzSD
ubGMZvsJhrGJWJ/UimwD8skHVzlgj18XhhbHEy9TkfvSsJOQSFl2myhGrdWv/IXw
OkpKU/Est84QN1cRAGtxlL6GNVhDo5ko07jKabeQuxqdDrYIgvn4pxdlDHje2Gk8
y61a3F1J41nu8qlyn25/TduWZ0B1M6S+JNzDtJ/UUKah3DHMUM5ufuBlb8JWUnAJ
A5UOIrJSVlNmZShwqXjJsmU+PfVP3kEtYWYeTwXi5P0vWDcsn6gK6RKK50NkwwT/
ELmAOp0mUuqk++gqaz8uozxPrKe+KCK3xfu3AhHyjeR2asj83rWu8+9f2akmdsEC
eB3pUv30ndiUy2Wi9BS73LnZfbCAJIz8lhmj9b/Hh/WcqZwSUlXPmaXkWD+5wyFE
uFQ3VzlX/IAt5GhvyCNowjgVoHQdaPDQrUH/PIy+pxykcYRMOFM/xO6JZZ46D+nu
JN3NXnOgAkXAOA0Edj19Bfi4XjaoNu7RF5763yaGfqQa2HiU0A5vt6Mgz5uguHh4
f/GPPAKkj1Ri/Xi6x/XaJqGUJB0nsu14kkEBvqooM3T3pfbjfChyfO/d4RQM0eE1
alKvtuzB0jl16c+Q9E4NJAZCvD42Q6An8czoLRWXJArNY+hohmNd4SHuP0DTzkmC
2vsIM/9Xf6+3DhkQGyRBTr864wn3Ff5VAgXcfshd/z8HKA67fxh7AQ7vFzVB/S88
2muC0n4EH++DjY5OHQZzZT8S/np7QidF+h0GTHHw5sHFz2rIeRxlp7p4ay4O8b2K
ytIjNcd8K0sh0OML0vUJjAmzygJ+H8Pt/lGYXYGWyynC7yO/k+tRhKF6pu12S+qm
mRZcOEG+tng4hkgAyi0qLbDjjfb4bJp4SiOWqzx+H3KDKrn+kr0RpWpsAvvc+oKS
hSXovDB8RnB2oumVmEC69O82p6/z1SxZmCNQr5oEettmchWHjto+pyRPIh3cUEyf
+cIqwVEPlQCgxBS5UdJRHu5BAxSDgwD3517RMkTh8Z7pcosV2hK9fHX6aAZ1YapR
mXQ951/xAw0X4Fc6mTJGs+4M2k4sVjR3BlGud9NTcRfX6OdmUo+1z6JOwxuvhBqk
8z3ez++wO8MxnMWh1Fu2I7ouUGoI55Lhh++ifTgKYBu6kqvspbaARfr+1V7XxviU
4tj74Beiz7+HAP6fkS2RhQVeBOEl7S+OhEbJDcFgz/exvupzlY4jO9+OuNw1iKEk
wPvqIzbmFZuTWSrdbtEiRWomBIPcwPotHf/sB1QOQVUCwJ9SG1yGLtMo8CS6miop
RgVnaUYy5WqkLu447pnB+XZtiEdP0HVFQ1hjWwRlXuWx5fFM2FAfbs4TVDh8MY27
5Mzg7ZzBG5nQqzfNh259Q8Tmo7KnrTZkXIE405Mj7uDJ3Ac1B8Hp+ECQbj6Dluki
KPviURwHVPzPaoRVHBFi+0qBn2yvQnOoi+D+Z395DxoX/c7JnSqiHoHyRAMQIJR4
3/olZiIIb7AzdViasCjI6Kopa2vdroWGtm+b6QBwFBuKuakhMRlqGUX6NXkgkQVM
eBI1C/7+br6VJoiVJKAlMOw5dUD/8ub+yKUu1XN9GqhW3e0DcxqaP68/5vW2ykbN
ErlVaJ1UYpxN6ulwmHIDxLajpDLkCZ6Oir/m/RU04AnZTzU8Iqb6Lpvvfo9nODT9
BAkTiYC8ZKguo8eKn8H1SxnLslHDbGGuJXWpOZEE6PknwhbonRMCg8K8RLfiqkhY
+lF6BnapMmPKja9F3CujEHvkzHjkreXnvo/Za9oUkv966tZe0GNRxW8i5KyqOhEz
ywZvDAVUg6lWE0NqfZi7bgluspSQbCbIhKGASRQEixmzTGz1C7e0AO9aDurtVPf/
GRyrzjWc3tFRliVkwe7lGnvvfXb3JjmDqXtbZgphU0LLZL5oRa83iN7YOuB8JHb0
1i/0V4bBOKAsTtq6QSbuYYarvlP/O3tluJemqu66YCkcC47M2MczoQUJOKtiGfTi
mZz68Xn8SiacFBWaIXn/Fy/kO9mQTHm9ze5USzFTZS2WSyJhxb77QJe9xVBx3Wjq
SpSvKlaxlk/rNuc0VwZmDLr2QxlH7251QXed9iB2sd/TT4uYLlXlCMSleby16SPa
u7n4fOImVc8gjJmgH/tissdh/sCl49WfEcI1aQs50S+5gDOZxDx3ijWCNWQ54KbD
UMLX47xg5PZ6/K/TOaT4CLUJy0mDZ3tWk967uY4sn2aD+Y1Fb+uSQ5pQZA8NHZJ0
g/eeuG69uObhVIEQBADteQUpl7kkxFtybncNQmpSa+I2R5344GFZxOL49/2zrl5b
nT7wI8Ey3VzKKzAxNl/a4VSK7kF9Ifc1d3j5SHXBB6qF1AfpWdW+cN9zjXUa2ccB
jrYsCURNuQXq9b306YOd38ofgQc1snCdJ2eF4KaV8oWlRP1cIXeauXTrw5LOTSjB
sfJaos1GtkmdbzFDOvNte7suwWLdpBPY0ifahIO0BoYik4tYWdayz2LpMlQahJ6U
o2cEPYxpYAZw9t8Rrr+NokWlfFWj8L1FcAgSsYsyn0XwoYbMIe1evN7SMwzfJTen
az+qC4FxelsF/kWghTe4swUobXUEV+ZNQYuMZfNnPAHG1oatGxRvYHvS+fIsnKAd
o8D4ek/83IM8UsKYMCfwai8eQ8P/3y4ZWmtEGEFTdV6OB9Q5IRrdEY0ChTljUOL2
pWWPqBf3N4Vw4RVPnScJid1lrzWGMiEvwkkqqVAfQBp7d2wm4UNcJLrf4vBDZbtv
tz/LjCvhITmOAx5eesg46lGmlYsDg1bx6DXowIchjfOFFpDhMj+8elj3YluBkmt+
lML1R+N9Yld0WyD2i+4OphmkzLvCuOqcbwkTex33EsyLYrbKJS+rP3K6X5isDmlX
ZVAYs0nOx6PPBqF1oewd9bKp4YbonJ88dSrqSmgT3HvFSaS52Rw2ex+lmykJb0W7
L8kMpoyA2ZUi8FJqjxu15jW29qTAhbBreKZgtN1mmZi0KQf/eXVrMN/ZCa48JpB8
Yhnz0/EN0pkJ0a7RpNV9SHfTtWwiBhau1JsE8pQZ87TEe6+2oxKhXWL63MsaVzxg
+ZkTQ5d3hKFfDjYBTQQ8AMMLCUo99VlILsgvbi4Opx0Nk2PhwHBOCf+X0fcj/01Z
LtKaxl9TegB8PJw6YSujpJhFxcSyn7kPX2en9Q5l1hXaDfjwYlT95hcmJI1kYK9F
UsB4+6jCJo/z0YSKMKG6CagQ0uvZZ/dOizllnDG+AvASxRTnmVEq+o2wYH8v9jsO
pj+BBSSfGnGemjVep5v3UEeQHV0yzNyWLmTgYJ5q/tufLE8zZCZcklsevHbkl46n
QpBVhRScVwh9CrzFybn7a5pYat0Q7XmuUwui4+9fkIGUNbQLX7QvS8UDxh3kaZsM
Pcw9E2g6rwHY/r/i5Hh+eMeF9Q+2Vsv8lQ4zMGVNDobARHc1BnxMXfJ3z1vd/CFt
4KkuUGOyELMkwOvKVliGAK470+owuxLUc6qimYAJ77cSKucmrOdWaPgCz4pdx/Sd
EBNOFE80E28YfsCjtZvvcyVUg3CM44eH5zy4ggrN3JEHuKRTSGuC8YiXcKlQNph+
7ibp8hSQH6DZBHOZi2KUGWpVKGFyI4tLDCRwyM/BSZit0gXO3HWVAmUGgWhXg1XZ
TAQv9eKrJbJI2CNzpAne6II/8huszXpY9XzZguBGfKXDKkS94VueK8xHdOmnyqcY
sXhMJ7aoz6eCz2ZVQCcltpdFj9VaWxvVPeEtbyiD2Q6aeJHoCuSO4sk4HBIXsTgu
QIU9xZq/rZdiJeJv2hvOj2rULkTvvEEi6ss4trHFf5R3DHAgRfcHU3DXNXTdcF2B
+poMkG6f7yQvJKu6qoLkpkAG9LHF+uQwytaCITTgmDmieiqM2qeR4IUiRtBgrzr0
mo9Y00W2QoG7OQau37Wn6XnkJk3TGITT86q6ptUdRwaIaruKoGAL7llKHrN7Y1cu
KCaQNhWNwxKAd6hTCG3TmYdKm9RjvHNF9fIfqNMIPvtoj3oF5D+ftB4EuZI5ROrs
WmMCq2DyVbEwbCdpzCWREro+idELg7jrj5vaVT4dXPkjIyapxpFoqMe0PZJU6Imv
DRBbA7tvjLbxlUv5lI2exhxHL1ZobpdHPfKfNN8mbt+pyeUUzJ6GdCZXIfYZKpXs
eE8oZg8bpQ/V6EWwm5ZFCD9PiwHufqPGy6NUz8UXMO6EWBopa0dCWTxznOMpha73
3IVHUFLKH5HGg7zeyeY6JPxiclyk21Ei9OY2dUl08xgfANvi09d94+gpC8MsqjBA
rUZZkcxivlftWshXr4cwk4RgVYEDIWoMBv36Ee4wAlVyRoK0VsZz+i14rLXIpik4
VA9Kpv0LksZZde3GipuEvnuwHLF+BjC+6EhBWywNzJieScOsCqn0dSDyCk7AJyc/
1vEOhazhlrxF1ueRcPB5e8bQQLYG9QNLfmFQxPZXH0YNuOj26Xe2ySnqtt2uvwX2
jzbC5xP+7Ur4RkTPs4dmbC/pOPGa7lULaA2KPaRgnLpniD8Cfp7skFiq7FXv3n62
ppEcYgCRi2dtHnSrQlMK4E3HRi9HiZCk8BO6ChLgDMcn6CKlc2yBdVjD2W+jToCJ
xcd7iOWbCRtyIHB6ue5CvB0zT4DvQ/z/HU+uQ3eFAS6Hx4SHaEEeDshTZwdZJXH/
6pqFn8iKOuE+4r/rHUZbKubNH8lug+Gfvv02zIAPSY3/bizGbJb2w9JRzoRLG1G1
TJ/u/cZOF4p8t7mXZDr8ribmzW0xQ7fmhK8YmderHDk0ajAZu3tulNZOZN4WdGlS
/oUWHOClqg8CL9/zudD7WCOZDn5oegVjtL81h4f8ipljw0weaTK80bbx4IhB/bNK
sr43ZYYbD+KWClj+ewiuMoqb+C2nb4ozNSHHqV+wP6pUBfuta7nYfOiQJDBz02td
GIy1eAG981pkYTAnr9IM64JoNP92aS6/6Udjoj4xBZKrG00hhBjfQeJg4dD2dW+t
vCkt7CdzpLCwQnO7BRua88CF25IK+nBTV3tElPvb6W66A8xOMWSXTRL922530sTH
Zv9xF7i6o/TGQw+PqpJX2Kl+wLZDKD7PYllIoJOP0y9mi3SK21mi6AzQSKmT7XJA
a69TXypv0WIsUnhc4nVz4xqtQNAyMtqoDrw4bkrI7LJjeeeUScHDCRmyg+HzZUMf
emI1/JrakeZYByuiXdOsIpmjOJuDEwe2b0e/vi0vUHrbPw5BO2O0deyCgu7V7UTg
NaINdqP4i8WinZ1O+0Rx5BI+seGtqmdgyTSX3eh5pb/4B2NNfpNv2qdwv1igeKsi
Wqb34Hqlg93/Kj4uDX0viaYKUYiZyH/P8csh+DHDhKbyfUUVPWXwBmeJN7AYo2il
0fXFjnrm5GYyGI7t3GVcPx5ojyQEOhIO47fR3GIDDO4fL7pgmxT6ij8GI48f+BlY
5QAE3aP76Weu7BkI17kzk2x59SqxHo+G+yrBdkWShMGz4Pl1eumbi0gyVlwQQLeP
ESAUHULtZTAe+bQ+hngAFEX9ZjGI/lihln4CLt+7h0qA2UNv+8cnvK6n3IK0xIEd
1wEDhJ3IJm7u5o4ElNPVE1SA466VtduChP694Tr50gHEsOIa421bhdIAxAXiS8xO
c8sbYtTDZ6d/Ic+l/HofOW0RL6ZAyU+cNZmiGVYScgLOk796JysjnM9kigjuy9uT
R7KNKR0Tun2M9T4n4ViYBgdZcIzeDGWSqyBb+jX4se4Tm+E1iAR0bYGFmX+m0Wgk
8K/qTVj7aoZlmGF7hbEL77gx7ceCENwUyLhKAi3xAXECZI481et01dJNcrvnvloA
/yezmnpJO8hoZLEwm2VowidrCBpyyM/0FMPNmxtqiY+FppOz91B/u/YkjJ/vdE70
X6mVchCeMbydkw3bMzetzuvUcIRfTe2WZmzP01IDXS/f5IGHZO/EJzIRKi5Hkl+f
2fbjxnYb9ZltLPWSTjycqtIsLZrl7IE23ixS+jCWU/6LhbF4Ru9S3sjk4FY5EXQ/
3PwToWL54rFj3imAnNrsQw/pV8KumV+zBKT+Pimy+1T4D5KPagnrQpHJhZpRf6Zl
GCc+wgWx7AkUHOJcHAC+IbKsPXpBLsQsMneVdpkazyR+xdZ/pDy9McRRZiZY95FR
cQjogvxzCUCWiZ5hk3wp0lgUiqVvV8vCRwBSv6BVLwNeroH+uu0ILHE0ttGJdmFf
zt/VqOPNh9CrmqzMLXpXNZ1gLIesNWCIkQtZsxw7ZmLM0YpvwH4EbAfMaHUalmRZ
vL7P1e+B42760yDRxpYj6/1b+lSkOzkbC3LVwLyAwdINcHA4nPWmooK/OJcuP81P
9GvZBpYpCrv3B76HxIzddS5iq6g7cGrwk6+sfyo6FnaD50w0F9j1sZJ32CJLKkJ4
Bnkl+kG1B6bL7Wpyt3POE/7j/U2my65fhqfZxKYlxxVF6ClVjEjlcsjMoGvCikUq
RmU7Y5TckGJli2b7ajX0b5OHE5Qn6FcjIvh+UYEZXDyXzFPlRhFA4vJSWLKU+NI7
eTe1MI7LHJTpeF9Dh0YsNGF1LfMsjQSe64BfJtob3nY39V4ImuP9hS8AJ2ZJ+JG4
8IfRY5Hy725n1TP+oSFvyIuUr/qWIusWaZhEBf6Ly2xQ28cCLKdo7ahuJqXfG/aw
Dc3MgtBgD1QnwaD+/1CrbXgH9J/02Trcudj/g2Wfu15labRSY7kz+5J12n23W3rD
GfHWabFzt3lKlRp3n1aY8AEsKW5mE/LmitqCB9dukALIZblNpXZAVp+fwScBka5m
e6qXQHLfwYyKMDjb31mtUeYkKEhX26BdRQk1EV8kt1KYauRBzWzZCvPHvMvkEyYy
kKpGXWJAk7SJr6/DI9sekTXd3Yq18sGtHm6KFQiezsVoaMJCircTaYh7Hx1TJ3jz
aTZzuNT4QXSZ1XZlozcdqqBR2Szd0dSjM7DOWUKxt1RITuJLW4+oAx24Bk+kFHgl
R/sUPBIlKrUKJ58v+2r+9EU949NWdTge24iZetiKxdG3XRwEQnOrWfvf2WKGykOQ
ltdkFvBSu+uhMy1REETcz7p3GET+pf9XSq6ZWhv75NHMQDmUenjO8/BvKT7JPSCf
ED1fN2JAgQGrI2UbBv8kOFkQB8MynWCHr3iUMYsO87YUEZtGeJjo5tOixAkCKrdh
yKjBJktsBZxwMAv+eV1OnqNxWWs6/gWA3rENSevS/z7pDJ6PuO/sC3Hi6h0ffoLz
p+Kxe4q5n6CS4sAT7dzck6DNjYiMzSTJ1xVP0kqjQoAOL6h+N29OYT1ROtvW2qFe
m6JU+J67h2rjiKkjhftjHsGZOcuB24trKv+93184OIFcNLLUJEewwFcCEZit6Tl2
NEvnj+feAwbx7tDzclqnhFRLrAD2boq8zMaBDjlabToZNCdgu5yWRNdSMQJaaQFi
RuSOGah16CsDHIFz8rjgkiIW2Uk6kFPllsIgH6P8UuYAhDk/OqwrNVzp30LcH55j
6+v9+RY/EZ2YWqpGUCsZmkE+BGxqP/xGOKBreS8EpTJmnBSyysgi/J8SWlwf24/+
LBhi67e9XLKR8E4Z89aRDYkEV55qdBKmE6qrw3Sb2StAAitrO7jx9qYTiaGKorID
h/smRtY5fTuygF2H1d2XP36Ph8xDFdRVV3JA/8R/P/NEUZRYdoB9+rdpN4ZkFJEt
3bUNsb08P2h3LFpYIBeq+KjcLTiWBbjv0p4bRK7dKr1lO7JlXrufxmMliaPjkeU5
oH1B1CfTDVU2ZpWsGqrU6raPP1v4khL+GIq+E9yQdxtuzEOC+X1+Ml8tUKDomEB7
sgXRLO3IKbFh2989+DtBqImH0l03t6GGCwzowsubieXpR5nurPNoEDUeRH47E7rX
hMygFvX6QrWXn9gHQBXbUHd+dxjIUMcwgyKBM1bnJFEAK9kI1CxpFT5MU1ofMinw
h/mBIQsDH2MIwug/uvBaFecVVLwd+3Hn5GSJWq4iMW88rdarkigRH5g56mM28CL8
BjTBD4/KQDUA5yXlj1AV4ilyWoPgyJbE/8HFhnPQt3W/U1Z17/lcQlLvD0TDW/oL
+Xz9JaAYXuJRFSXFI82K9qbzAkGtA6XERQh+h+gg5rH76qpj2dBp1K0zHJkG/wR9
Z698LZUKF3WCc/1h4657z737mrvjukOHlyPJNZjYpJn5DM9uIOLboz44z4qAhYz1
62ltYlh6j+TetYC7Ik0C6QReY71cdPErs27sPgZSdAKgXwu3ELnmhOXXGw9mNT47
wX9o4Zw1lWU8i7j2xy0G8lR/qkrtIkKQZVSKt/ief0KIJ0w9OupDELliVC6HAEc4
JI16X52yHNtQTtHPBLd/jemxgu7NpmOT5/Dy1qR8Z6pDT8h750DKrC21r34DfNYW
VuoktLchT+PKmvfwRExv43ePQGuDwCMZ2y7V/Gv6jWN/UxedgCAYXpabP3p4gugz
5yCaJZEg4bPj+GLjCfiwujtwke/eFc4VhLF5jaOYDyBM4lwHK6SV8BcJJ48GrEE1
FXoJZbd4IDdjvjXGL3tLHejZDegCZxSPAW53irZ5Yr+6vLef1Lip0lhYncByQQc1
8quwZKhdo0uh2YtK3R+IjsxmN5rK/l+ce7kCJhCAh10ulAnVmbV0/myYtZIfRsMF
toJ3BdYHmuUXbNwR3CmJZmjd4G/xW08ixx9oEg625o7h0tvQUtkB8i12VaIHnBKs
lW5+30pFdpZ5GCPH55FAe6U2jAF+cGvBl8GFzg9tAGJ4CdZNrTt0VBZP6CbU6fr6
CSX1hWr0lYSEWPZyBweu7e5rYJh+YpjNFXB8YZlOPb9GV2D/Z7OZEZSGBIeCN6Uj
AKHhVwncpUOkax0z59gTAjh3fSZGbTePNdMmhrJZeKt8mwARBi5WEHYy+oX6tzEY
m+oPZyM4EfN/tu/rxysWJKIh2dw8ZFeLgcY9zO2C7JcwuYyA0WQFJPLptrjsO4aP
G1SGWhV+9HsSm753CcsQFed4S5UiiQpYI6RSHhorywpV6VpWTaINIaB3pRKmVLVa
po3cCN1kKFkIaJao/+8675zkPn4ION0aFe4yWhI6EqmhenH/aGy9Jlqx3Xp6l8iQ
yyiHa3UUhjGZ6/Dve7tOcezcN36GKsF9+UVeS6tFzUnCrZyWsuVKY+FNfugop6Na
H12HnCNP4+mXGYeXsi6U4f8QIwcB0YhqXLPzZTVufESOE4555FgiZG26Q8t98nPO
ZjuNjfC0AxM7vS65sd2wkxrEFepxSFcDAN7RRGoDm5S8M2OCD4SLRGZKlKdrIxYS
VRNNKcFI9Ij6319RXDks44oYgljF6+2WWK9zoLhTeO1JpT7diKt4s7LVFIU3hy2M
aCIKQjEAs7GYqDUDiCtFi02QkI6w4sKDWWtMf9VIAoKUDBRjEQr/9HBQUC2+Auxp
RNMdCvNPeJMbHQMxYnOivkn2sZQ1FEfdaSCYrs6wIZ2b5TP8sSHJK4PfzenX2dJy
dVTWWRom430up8ypnuVg/zXpNUHCyLS90OE3/9e2Pq9EYqcOty5fRjSWhPrjAzAM
p1GDiSP2tAxGkuR23zqdPTeYbOuOc6UFGXHAgTTdOh8rK7VwIoqhdwf//tyxbMG7
HtYmnyEZM4rYFXOOvgflDC11qfAC1fx9MdGg5vaUPniMxize3MKGNnxy+CMAHvuI
WSOOGeN/x3N+B9gsWte3RDD11fL+NR5y5KGgc08CYWp2klVehW9+mynOkCjMbI6l
mgvEIoSr6YhKG/vTTDnVzzZHn7y8i5Ujf5UzRLBHycXnVeU7hIliNt2oBnFesfnU
d6vgawg+SZB4Z0HHR0jxeCMfvV6Y8KCW5TP+0IYDCKvhudWJfNU0aikbiRSN0CnR
s2mYZSyS5U1t9GmT3Fn2s9X1NxxnbQgo4ZLdzXeTTf87bP+qOigTxlBOF//uHtmh
08IPJVlxkXcAbzTmaicETqhd4/SM7pBoftMXm7tgxIuyusqJpXaKCHa7qqp2wD2y
LiOWrc6hEQtZ66q3PmYOp1iQApNFYi0LX86etizFO3UfBP5cB/g1ofjxtPQBdQJF
8S4q0RERfPiVwTZ/QDbFmsq+BlOEh8M697M/6dTuYYsdV1bbiISpyyF09tmiOlyq
a11zPmZPGbiu4g90neyY7Lk8KkdectIduNskND3KR4MHQOqum6StmJjIAoSqOw5Y
9SsnYyzVM1Mep8PUltlgPea47cxZNOUystDS52tu6DLiKcwAhJP4zmrEO2hrcS5s
5LC2V/cm+5YJbzLd/q2Kf6/yZIQ25emhmSmLfV5SuahYoqwUprBcJ9mqKj9zcNEd
o4n1eBGjH0k3doshb3p6NXfvdvjqYlozVkTg1R2W68KDn3eVPIRvJnaIZ/eihwP5
nlKnl9fdnn4WALQHob+pSSR8tf69oi9+VEdiZK9M1ul68eKuzzA/RKnAtBTxwJ/b
f8baaVtq0+ugWQL0xgNewoRh/dDgbfz9HQcTfi7ZUdNDAKxEw3aEF9Vwig5ctFWb
R9Y7mBlT96S8IDAvuUCVuxVsbpOrSERZFe6KbLfN0WgunW1eG9wi4lvGhSG9zvUm
ZOeG/WlExAP9fpt9QdlrZSE5hjm//MJOAxS303W9TPwIMQ3wXLtDKAOlJmDMyZFL
HMuhDapE2UMMPlhr/dFG/hVzE6YtSD2EYrbkYh1ooQ64gz5Hya1LSwCCzD50WaNi
T+86xtHQxdZodI+vhiha9ZLi4IjqcZI3XLSZYHXkC5LY974El4c93XZiTf7FdUUr
cgMWM+NKA8ymNF83L6xQjX9iFyp4KFdPC8dTBtb/Ufo3foqkFGzvD5Z3o/QzmMiN
g38gsouESPBpHMiqPCoS2iLP/Iwpkrz7cchqVQv5LCcovSKutm4o9dRbnNmRjF+G
O5X9zDmbSRnNBnDGoQlTQRiNSImBIONc/7yejLCOj6OhnZ+CIdC5iQ24/McT8ay0
8hktZDk4fs0syyc0gljeXeVPjm5Ecbf+m2LH0WyaDhl2t/6+j71nhgXSfn9F66kr
5wo6juL762MFqqFbyJr5oTP4lI88A8Xu7BjwHCOXGFcAC+axdeuQWhxkC/bK+xKj
RONDowe5OMioRntVzSlquyw3WTuCBufcug+nW9Ps0gjnYLDMyIG30nY/Rk17DoFy
2b7bUndess6J3nk0uDKEYZ3P/4sVGTnkC1rZPUs92vR+6gkgnXpLp1ckcnef3XEu
fNxrrgVqwbxBUlkJ64SOHpZ1ZUGZSQucKxvNIJ55rMbTzpBWqxauEEdQuBI0sTS0
VSduE3NgyB0Q1tgYRXKtBAWuYbir9g8tRcviRXCMoCdDtbgPJJ+1bX9DKdrklWcF
dwgEwP6UTgUk8Th22zvIm5FG0tflVI9rXSXWUduj1PuxpUPmDBp6Hkdqn3e6u77i
3/4Wf9n76qQSFAtUxT191kUbIWsaLzfA8tX/kWAVQTHZHvbFOt9oFGm1lmN5XbCh
5imBIatgtZlrYa9qQpCtc2PfbUp7z+N4bJHMpdT7I0vRKoTqOpARuRZbRSbA8wam
caTvJxYL12px37vYgtj1rZEvFEGkqTA9urjrMluQhBaIe1p46Q6XF1Iam8RhYUCs
F0bDA9zpISXofEFH5INv4o0QBJKyE1VfZrjYK5pFmH0tOH1tr5BOgxCiPfcN7wJR
Krf6SHeDQJiFKtj9v4tWEa7Jkg8ZEx9iwnTRq5ZUIMxsTspVe/rhTo9fTs/DY7RQ
udWg0HbkrQDutZ6SHF3arFoa7WehU9c9QUpkLkpQU2G07g62bg7Ga4JWwr8MSbal
DLxneGwnY8qY7iFWhV2tLPi1CwhUuaqWmzwHctQ2xpKmf9YMQDb2OOfZsaamGsP+
xUbNnq2mDD9kGwJ2qBwLygjxSpKZYf5F3cWrbBRblGndGSdkKyJ5ZmBcxPHb6o6K
AMWlCGxabC9fpYySsoJHh6CdUTYSUiszR8Kj7/sPEcVJdWyg5jajOaQoIamnrPl/
2kmClibp+aWmOVrP1X4AqWZeux0sjCUXYD/8rNMAn1xnQIGAXU3xn/mbeh0KgvyD
8PXA5oN7K9H+rniszxBa47RxeYmTXko3TA2eTS8wzsmxkhWtI8tv3jn9GBhBtkgC
912E5DoqToUYpzE9Ay7dd3eWjwfLr8JktpXBXZbnf0E0AF48yKcDN3lOFcRnD5TW
cUVo++HhtxmbapQhUz/StqzksJyiwpfgpYrWWpuMWmcv7Mf+AKq3z2pmBcA+VUqg
cT5duIFlbG/7QWOsUh7Q7BvDAxEdraPNxShMQbo3yDle0un4+EDyi/uKKjcJUwxT
oaVsoVLhy4y7gcUxVQWc/kbTqIStmOq2GhVu+dJm6K3hPuD+5KNsSF92YPketsJ/
WqVrciyOmNHC2SK1plJrcjBQ2mIojxyuJCaj4B4kpMvenckgD2rlZZush+Xbp2JY
QxSs1HfEVbnmRyt433mxtwVcW2nrFlAeg76DyQ9Gb60eLT/kpXvO6Kagy7CZ33WS
CFuOMzDx0wI9PO9Ig834xj1TFC5WfhQpQgvbv4Di30BKqatLwRMBue7AQSo24BdE
3uPOUfHZYMyiDnE0OAYD5dul6pGnLVjpTJeE8axCN2ENgwBSU9VXwpCgwlqNZrg/
jU/GE3c1JoHB7+RH1LNg78n0M9M/o/2zgmY+CkMErQOGWFcz+sm4104OP1djPCqb
Fx9ciJW0TiOPXqDKadSMMdIu/suUkoY5lNL/beT/KZgu2FxvMqwC66YzUQLN/Vqn
a3s+K4hAjYf5QfBNpTALtbXjGwk3vmiyUCkJn3vEcD8lnOdUSoUa2tUQ18voPodx
kclhCZcfywt/o++hDtRwPS3E0dcWAvNdWmNPZSbTf5RvQ7Ck8z7WU9JYZH83Gb6K
Ug2nR2UMuGoptCKUFeA/eqVLLlNLNnV4Nd7xbKIQoJiHyarMeubYsIYLa0P78ap8
kqI1jHnZenbPL5ZYz0cPs4O348YthRUQVpENAI7h6CZ/upgkIfPUn6iMjRstSWjb
4jKFRUggZjov4IxsdJKDCeO8i/ph1EXzGnsFeRwlcmpmiZAhYid6KCnOlKSinBks
ZGq7pzAUHT71KBl5jqaNQ8FCXvSHdKsol0jvSQvwUj5s+SlN/yIu+tQjFyLIClEH
/oDbC8E7Shc1WlASwjSgjPDne4RRc8heE+pTFmX6yXwaXUXQhBqrUhfqG82bvJgo
Q4F4o1SPhxvG3XRIuQQRUUK7ptALT6S5gtrs1GlBsWMhKx+P6mY8aj/wT9Vgbw9e
hevVvfs483QDqUqNYjYzbqwMqqH74fdm52vg2aRL1vHA4XhL6ScZtzE9fact9Xqi
jY4CQsJcOOYnjDCpGKr7Lc/AnZBTv+OmFqkW+D12YGc96K+7h96thBaKdHq17Kn1
lLF2JNkVQteFDnqThDsjkRbwbWUt7cY/Qx0u9GkMfqNSb4Ds9nJw49tf2JT/iD+/
mv7H87SS9/grFdNuyxx8V1fyOwtpdypmwwIlS5gEoJ1u+HKEjCuuaiFIaWnBLAyY
iMJelP0dvrc/1v/JFTGtzQe3KDMwf9X/uZ2zJ/7ggxbyYXAohCfh06hlK32FCO+K
CqN5i0S5MMenyFONFyRuKRBO4Ej/G1F8m2/61/Nkeg3B0k1XwfQO/+TXw8cEMIL8
ObAk+TPAekanHLgaoWRQ+Z+CHBd336X64jKTiSXXCxtpz/pIH/9YR2Aljo+cyzM6
jtUZhprgLvNRYzdSdLY0ov2h3T0T7j+QHjvQq6eV14vgJ/t3zzOLhTa/GKUT4Gbe
xtXFpwsME4MRNtohJbI1eh7sKHTtyhnoaWzMj3BjmrW+NDG44e4RkIx2XWLxkezu
aBXWrlN5oSj/f8b7OudFrZExlIrmacR95viz6+z+BM00lHpJUPNcujDLbZ8pm95u
Z4Ijt9YK0FmRVetpMZLKEqkwbh/T4gH5eXpYjuBeI/NYrKn2hNOROFzDeMiIu39U
PPCqOUke/2zQ5A9tixmU8xHUM+x4IdX1GoUslAKEf6Abagi+vcop0xOgXq18+iIG
rwvKnEvleDHaLR8LNKyNFw3yu4WiFTxUuvyn040FAsOGUx8ED8cmOYrd5pRhBfjS
r6t4Kt743mwCw/gYn5AnX8Ng6y8OgwN7Viw0h13dhMl5rqem3W2XHz2IYTtfvB3L
5CBB2BTGfJt0oNCecj2tpgl0MFa0LM1ju5mzfIwB4HIska2i+9HNnj3XXr4rzmhR
6c977UFs08gSKJMZCOK3gZGNfU8v0QYyBrZ4C53zVcopqY0JbM0id0AOU7dQgB91
sExA6+ra7EDPqOszS3nrkwxA9PYwZI/leyaXjlSs37QzsKj4omzplQ9lfYTdhuRB
mux3DKNM66P7NncrXdsecHz8HEFRt5a2C4w+UhrOp4V3sRScR0f+/RafNJ56gblO
YEuKd8HWPwJomthRrkCAJ+wgMl4k+B62CQEQ9ehKC7eSMfmggmLBHfvEgGntY8+j
V/MspnhaZfJ+lLnYXuOLpXT6naWLqlFnkHET/qoP/JJVAg+blu6kvcFnXyt96Kvb
vdUNATAKwjywg3XFih/4AfpjKBaGd68QV1c96gApWU8rI6HpyeaeZrQ9Dwchqi+2
2VnPHqvJBe9ZSFoC3u7BCZNDQf34rZgf1MF4sw/OmZEn9e4EjSZ8a/lkoO+f2Y+n
FGCAVYg/dQxqdDLMHphhGB8HDPh/xqScFvGPNRaiW7oLP6JmkI16J4soNdvvGSPI
+EQDrx64+ILZiNUvpE5jrC5KmPmYHp0XkQEumHf0sqXR4cj1iV8aa8dGCOKwov4e
dGM7e8JwM+MdEMFxQk3ezDRywSAmnagwcHQvsylMcMORKjsDAsdO65rajuVpemJE
2Avo6ZkGrncqR0dRLgCNXrOx1O6bto5vLlR73r1cts9hYFQU9TEXymw6P0KYVxpj
XBwIi9oEwe4yGxTiSDHi/erMwWVfgm9ttG/UZmnMc34+RWRGhbX0iXW8gZk1+76o
XNElZxMYHGR+7c5VZTmZnkvrke4viPdtMVr8uw5zxSJgXXHy1HUMZSYmQRtuyktE
sfEHDdjKxI4Wf2D58I2dZuLHv+QFxILKhBy5jXcy3qrrBSHnarODIg4QWBOhT0j3
vTzTedXqbYS6C5JyfENCozNuBZcIOMBmjtAesGeWUqhyHV68NGAHePflTYsxw3VE
gsjT3feQie8gb+N+EwMBufz7i4BwHoIW1n1fbdbNFubaTXo9VPPt9n2lU3+47BbX
+HTXg9LroiCwcDehziT59QulISBnuAQ6RIEOzsBEOxx2K8DbKy4uIoIM7jpi0plS
9BqJVCXnRlXL9LuBKmtlviXyr+eOz0wGSI0f0h1yovUHndoCsRcGIhg8DW6Xxs4p
QKos7HcLDFduTjcAgTbyT5YudY0SyoH0pjPRJn8yZpdm1UPLjZtFbuGCXmzNimbE
x24Xv1BGW5dBfMmnQNtULrfiKk2cKcWY/zfbn3go0ZLjDPKPoOGkJKhqUvtspD4u
/L00ujSmpij4Pdw0i4mDny8zD/OS7ftHDxGr/GhqtaFs7ScwNI7uKojMQBSyF1cB
Hr63yLdM9NT0OSe631WJ6+ojUb4DRJSWAgNEN9tGQWAslVO8Db0td7Jw8uR6hIFV
6s9rSG0yINQiK+B6stdhN7FpEhX9pevX9pM/xy40pgD3xBzHivwOafbwtIOn3FQo
LPBJ1/nMWqLArs/zkrsR/FJ9bZpV1JfqtJ65AGNyntGZgq4VOFdb+wIcrOuuVUmk
cCERT1fXSFvlCWAtleVqMIzFBmmVTwkFoTz0r7DwQlfGdXZnhcoVwoO3G6SGkQW/
460Hc3eJyp5t4wHAn26LUa5Kph0GAKHdIM4HJV7a7Nn7pRqgD7h0YJC+CipF/gxR
CFYvH9Jy4OHwI2jNp+Bm+mCULMfo+NgkZ558Q0PImL2HiqkMBkcTcSenE5Mpupdk
LkfO/6zT8E1z1l4elfUDulbeDepSHe7xO8Dl3Bw+GLtQcwnsye53syYSN4IWpDM9
/q/CN5gXDiCVn3k8Srmwwm+Ai1Sd2sHANV0hk3ZszCiNHUsksD2xZ4aKJw5frjWN
5JipM6fyAOFkrTPaYeKUjblMA2O3j17zJU8IuXmGa6Tv8X5frQZAIfuYe2A0RG68
ejdghAz1oDaHJs052XtvwnZ9vbI/ClM01mGU9avEp5dRV13H3StUyB7u3tttIvlJ
0SX0opGTZ0yo2pUZ0r8d5rsYJL9Y/hfSe8SK7t71F6kvP2CUlaxyF2HfN0IqCpWL
nAoFCuleUaiLbGAhsP5VncyMk+eUWreSmb3oA5t30U6LNaGd1l/EM7eNPcM0ITX5
NC1mZGa3sLsoHgG9TuwAiEPQHAziZDradJnoTUziZiBZNlTAnUfIeMsDFFRfh3U3
pIE3ptEhaBvKMAAb4+IuhqBKKgRQb4yFCk/e9mNqyFtT8HDaaSMx8r9kXIncJDJX
kmPzSnoC5UYkTGpZr1EtetUsAgj4s6EY4iI2itsONMeYxZtHdOtwVnrnEMGCWCVf
mNuYDmn8H27Nd95RLQ71ebqteLQYIajj6esN1FyAi4cJSwoR8JN9lmr1P+oXJUsV
+8s/v8CM58z4SgvCqF+Mdufsr6w4RK/5zSNR7hYJhEHn6NTUnvwqGgTc3qD5Z6oh
VhMEjIo3g68oOct37ov3Ah0AVT7a9GrRlQ89fN2fAVmDa7vCPdfLNKadYMGZxH8b
dtfIG5O+9NqDPoRY+kUDRGag7OAUkdoTCkbctxJcZTgHpCOKNWYa77gnpyrXfQNv
rlpSVfamvMRRszUN3IXjxOAMA8J8zoLI9OQQnRcAqbsqvvKGHCiT0mG0UVESWj4c
mGkhva6MjAXXhw4PCT1zzMpTHEDiwp+Hs7xbxmGbansZYanhcvsJSy8U7eC8Q5MS
XZS+JMg9tRZvlokO2Fe45Bw/aU9jDDTM5dA1p0j6SzBwyEIcEuwhQUIdooNOd1fj
aQ9OhzfDs8lX9BNO8QBO9SMwAzJ95X3ERqVqpO4Ek2ykiNKd8LdZjieFU4237S71
o5n+1KJ9eju58jBr2XXctyV0+abG72o7EZWAowBUTWp9JccXRCShDyrdq0+b9d5W
A5BynwOg6XAlVA65J1uEFgg6JitxkKcz96zDf7MHxZSmzDUZyuRI6apOE4jkrai5
LMZl6EN1SplIMtxn6SD5jpvfPQqmVdy1LGctmlXNMqYjbalLNKiqEqYLR3TdO+/6
/dizJ0iwZVM12V56vzHwYrjuqjZIqs1w5VafS7sDtPtMdFGFjpIr8fpEjVQDz7qg
yVzhv8jjtxuCnxGvacC5SEhpi/5s3Arba44k6mEG3S4qHNA1nGtjf4Dc/RWX80jo
ofnNsz89kSPNRLulSbzyKTWW57+ZTjh6SoUp/HzaPaOL3vcbO/+wm/RgzbX9Bii4
QJwAXndaES/7MCRkzlaThESx5nQXl+2BWa1yhSe2a3QfAhXM6U1Mw1TTeZE/SHre
dn7FWJtglmTsz1jf/TAnxhy9cEVDniRc5jd7gzOjZVQLKfrAClAmwZmaF6IfiiTV
DDhEXwExOe16ZymIpwlYGSG6QgkPwfBll4ONxarvM5rKr/vl4mBqSlcmxB8H3sBO
Jfs/FYKLnp0SLK2vUZxeyhTtLfq4CxW2hS6KIF+CUcqnIdKsdxQbhK6RTCMzST5f
KiiAgDQZFpgCg9xXOiwpcaDdCh8NhyKXAsUfDIRjXDAupZLP7qaUegm4WHfgztT+
mh5tQldgKJD2elCjsGeSEpqQBAjNtcvInswCKyE3LLFS0cYYTJ0C0BHgf4Iqxw21
VcTZQnQfcFY7Dc9detUOFQgsGEZZlt3Uz6E6sE+cAqrzncZiCwtethc3CUv35zCL
vVkrllUPiB4aZiQ1iLMAK74RLnlh3sHBmfnWPNdTxtYwlU6CuHs3LsufNAaA4HC7
zzHvwI5kK9beQiW8fzwTYGLAUbhOCmPbKA8AoRF8j3opjRVQwcs+sfgTs/q5uLnP
X5cSEWjEqcQcmXu8c4pjY5wljHkg9pAaWxDHpPcWjMaZq8PxXa6/qwsLSLXp3SIx
Larv5kwrTOM7dFQRYETk2Mp8ZWsEGi1UfoNl6GKSeqq0p7Cwbs1paBMhA/5r9XvO
KZizF+nHWX/SndGuTEY7uLYCy+d1nSUEMdFd+dDEE00aBGp0OJ+3YqMjCj9mz7Jv
C77bAfOz22UNhlN8HfeU+TWOv4qW0qg5RVU7VoHNV61oCQBlgzA0LQx3qPijdo1p
Estbg59e8U0VAOttinm/zi2U00LYa/siisI8dFbiEFXi8cYis1CSR99eRaL2N2V/
n0mmpZ+hPXAt8t33LfikLxfH7aaeQdyog2gq0USXAp5u3qyFCLRfOpy6Skm6qegX
/iysK3OZymM3QnX1wRxqC7SPOMV/VBDUnVaW+O9GvPpl+LvM6dllnl34Q4qESkhJ
8WWE8HQKNWkyp2XtgQSyeY9HxaRdDJ5xU6+Eh3ST+TcbC1buTEj2oLaDl9DY4Uoa
euX/aF066a6o2PWtBLBG3pKEtx49jKxiqWj9lU6B64HQ9LL3Gz6fcDRz5y1pxxVY
T/AXlFi7XOe+y9OFgBLGqhfdc7TqfrH6n38CEmNBH/v69ujc8zrLBsCwY17LmqcX
7s/rVWq8NRPVen5T8FQetaKFZ7jkdSC2s9lxJJ3h+ehqlADIoQYbuthk9outkDzF
vebk21aVgrpIzghLxwSZfLlfXA/XoDfWbIw+jmT9jj//MR0c5dvYy2Vt/KCj+BGm
A/bNKn9bfvTeUMf+T4NpgPtGmO9xA7Fp9ux42B4NhHNvMY6quWOesm12MbNiAjvB
/B1Qx4JPHv9EaW689MDJbhcgFK7qprVpuGWghixp6E1EroA/dkAHRwXHC48I0Hqv
zGAfPc+uw/KqnyEHdXxARLOJUwfqDEtK8WApTa7f88kupgeTxfk5LDbIJwECuVsh
FW+Tl0dbf5MVJJrgVl0dOnVFXYcpXsgQCM0Oe2zBhUDk9/tmnwgwIgpkOJ+UqxZb
ookCPmf+U6QXc5G57Tqymybo8hLM3PVXhLb1PK3vK/xi1zCy5Vxm1VEazHHHGIIT
8OWKdZ8E7XvjXCJfMJMpbdVBkLikb976i3IIsz7PEKF9JBDbtJGcTnW76eoR/7c6
RiScmukfPHw+tob4NB7iljYXzV0+cZNa36xf9Ercbtmdt6LldfhUIPVtKmi4d8JC
7QNKKpxVp9mQotvCLTmXO+U2rsmbXQ/DJ942Esl4xgLmPKC8Cu77n4kPB7zvL29L
klJ6t9JnYc8+KwAq56kt1HFJZQYPH/ALKzsHcp2eUCEr33j5HEyMrti0bsBv3cRa
IFRhz7t8FfS7NZRuI6XKoFcvXptXkcXkhGEMh6asLrJZKnW9ZxWH8R31F22Lb4S1
F4cOyxz5JVdJR7p4R72OLnbPmV3RC83RhE1FHmumMx5HDbwsvpZRqEb2Ahn2l5pU
DuBYnHbaw6CWO9hWu8nabtuVr3Y9AoKGYerKpj24qPo/otSIxoVjJiiYc1Vz5xLZ
gujkuz0pEnn8JaJjzgX7sS6OxiZ19TtNJbHKgZW5+N6AnolMFKrVQKPtwx/U/cIc
nchLqIH4+sQoXIzZ8uYOeXTpUpBbSNcZrddyy63rJEDyHfsPtPQUArt0Ii7NiXwq
v1mxyAPeRt1seigKfGcZhaxgsMJRn6O/QfsGiRDM/f5N/ZOy20QBF2azhmrk0Zpj
32l+vymRHgzS7GQbJe3vr/o4y8HVay9KzrXyAD5SbpoRuw4tHU0lujZ7lFwPPqyh
88WUzNXKIgohbQ2bbXeSS3OKNunkmxwtYASgDfpRoXVl28lN9SpYR8qS40JL44y1
yoeXoZB/bnoC39IXzjvPu7xp6JnaP7pzofpRggXRkFnVAetJ8mUsd3m+6UYFt63s
w1ZDmU4YpUEcGhnpa+BOPzKyiJVSqMDVLMWdwH+zl20ORiOxFlohjZo+KQVM+cuj
HOmHWry4euwr7VAOdENdgpwzq201jm1tN022bj4Tb5M/BFPYd6G0zx1stGaOPY3b
eFbXwLlidgw26crj+MxiGyPFxYztQqETeV2QIlLEr+GBfszV7USleybMfspBGcHk
ssMfLkuXaUKQDlqr5NFaJHZsSwz3cPRDxLw2G5nMRImMuO5K8uBQ0eos59D0gJ8u
EHpkMUKps6O7L/yH/t+d8/C8xK/N/o2xTXaAVNtBQzM0y4JPnxVREPDni1PN9xGQ
kdKCKQJ/hlzlp44Ioh449QFgVwhDNDnkQYSEw0ls8owb94s5io2W2NP+fI6UApQG
F52Dh5t/Cwu7So5R+QstfQgBCKPiXbyojpr/ZCVyI3VhFrE9Lvzo+wFSlXB8G+uH
HaD2FukXKz5lKDe61CnJNQTFq86W7Oyb+6HRrI+yGcIypM80kFT7UYXAem1WiYwU
xmzJ6ylNKRAPMS04GiJskJqwM40RP/2QcrtrQ3cQx7vAv2h7aFusALkPlzwbTT0J
JV/puJAfy/9xnvMDtgWqyiUnp1t0j7zvXeMjjDJHHSVXEWdkVNDpENdYUf/eR6ky
r+TV2L17aPCBXOfpyVfGWmwNNj+6rcZW43wwLu/njeM+tfAi2Ao4IzR3OwM0uKwQ
HFBSbAwRfwY914aq/DDV/iYg7HJTsl+vmjgaDXD1FWwbZm8+903OdOIehQiireDA
1WVXowYO3kBCwhW/bu4wzfLyYHq95+zveZl8k04ljsfdFiGeGqUgfFgrNcPPdkGq
we7n4jyd4UQg9ul1+pqaPtnh4/4/R5mZshrei+IUIuYuVmaN8kCSMMuvH4/tBrGB
Cjf9yzLDyOhZ7SvGB/XGGPqgMj+Z3ZP9RqjXrdZEG9Ml93iKL0PAWG8hZzG6Kofs
zEWfo8byCeNlJeHR/nMpMnAcCq8ttOuOkgAGe5deie6+58sX5vjzSztpuBfbCgCr
5PRRXR/jhD71vty56sGwOV2nSAMC8bWeVlhiOUL3lPUKjm3vOSRwuyJVL3qe2e8m
T66TdSoTPkZeZnON0ZmjnKPXS2T2UtHV6XFaci0Vk6nDPAwFtGzjBN/g08eYylex
X/qFIYjJcY3HYp9XXAyVQxPI8ks7fTIYual37KHpnWNc1NInsRm1MbnYTtIzBhsT
2rAjjBvIhNWQzBcV8s+KMNuERiOnZkOTVwupt6D26TYanvW9TV6rDmaDXu6ask6i
O8Kvp9ciTy71VmekDNFjBFPuuTzyg6Xvlc2cIeq8y+MvDniewmB7GJwUFy2BRPln
G8LhcRc7LoMOzCL8sx6NoGne9P+mP4e7cqkdfzsGBVIz/Vg55ygZyOa8nWR+6eYl
it9h/y3H+o9NwF145O/ZvhQR7dh2eSrVlftRV+8oL2vlf3iY0fRvwchFr3dYjTCs
9c8TULc24OAQT6Ek8SaPxwV+P+rlAxnVc48yUTfF6/v+2DhoyvHKSxfWdU0NDzPL
Ln8GJtmZGb1hg8tVz+MWyTXKotIukysXMqDsFdGSzYcMccqxbCBRJIKRt1HjsofB
IrvH9KfczkMFm5qx259NBIbFptmHbCPZCJhdoGnGcvbRSwplAKTIb/YBwa9hB0Ed
+iqcJG2PdROWEznoV/tU/IYXNYz6zpA8HJA/k2cr++j/ad3PoPpANzTd3Ti6RT8T
edvH2/jsWJlrfCAfUnCIzYUg+jGbBS6QTmWVSSRgOSXyepKN/8BT1t9L2KI8D9ep
r+rdu86qSGF5+BWWQpXsENYhPYCyXnh/PwghnnL07IJTQkDCE8UWQsZxKYTzmdcF
w1BfWR2uBgz2s8HmiJqYlNNbrhirxTmHM9/PMHawkuIOMHH30s3pQw4ENAwJmUZ/
Kp0fp0p72S/qlbbgDUO1E80ICKtxY9LSRP47LQD24hqGho/dwlst9luNGZET9VEd
SZGjOmTUB4IYaS/bapHROyCoRZoqB3Tej4BFVAgIdK3jtTZbZJIgg8MPPPoyeEaJ
IdlTxXVoCxyfkNEyOjLF2j6LPxRXFqejMN3iXK7lF+8gtioc8GUlnkbQBVwB1n37
hh+NXL4esuf+nPc63lkny7yzNtmgo81YtKrF0ekXyN0JCn29MyjZJ29s7uQ/7r1E
BNsNXpA136ojavgvGaAQB8iN5QCOyvRVhxcp24fWYCoUeKYz/V6ae3yX6mqIZvaB
8Tz+FHIsFHrnV3jU4FQT4vWc80UjkxDIeM7I/knH5Pc9trkTTuasVUjXGafLUu3R
YJgFJrhRTOpGbLvlqraTdpR+wS784OevhsUw/1NHEnn0Fo2RQfpgMbU2fgdrd2Yt
nuzxqYexdcd0zjI0k+iFpTkbMAnyMLDiCUi4W/xo3XPNzbtxm6dhR10E9KUW7XAw
d4g/KGyyim7wXB1ZHm1YeZ6niTgLXUyKi2jDDptUJvCLoS+Qg9B1MMaYTvKCxyzf
fuFaZZ93y5JF6WQR7FfpGal1hja6jOyyPJ5zFiEh9MW5BN7aBZj0wJ3sDkVu5qEp
afmLgoy5eMF54ufGSInt9qQkBLD8ux8X+ShzDiJJ7ozxY4qAaaVgL9O7vy95y6Dn
3TOOmo5YG9FyQp870bNzWOe78QCmaJnpsVxjVlO2u/9vW5GOi2+RosO0I1AFCaxe
6AxWac8NfbcAWzEHQQ0C5PmlN/3IhfexCkJzkbyM3sL8Oj30xKhSJao/hvMwarKF
ts5f3b8Z+zXdyyRKvJvLJsLaRru71o3IIPpi0xMaulQ+qupBCKWCrtXgawO7BJMx
9CeeeZySR0jttXWhri/I2M4Z9KO4nAjXXz5XhyruZHR3Hl6EZlvatD+71+I4k9Yt
OdAjaZZ20rcltcErGICzkflR8L82Xo6Lb/he1fGHHnOwUBQNvqn8tEF3yQHS/YV6
pHqplsbyVgwumVifeB4zlsSgdDUWv1/PSHcfB6Lu9llkCo8JSUxyvb4PJkJ/0o+U
gMEWUl3n5FnpfVAWnLRb+ziJ+J3jPqx2Tmhl7Iti0Vn+m6ikJL9NlrueFgV0lpZu
83HIqdkzmJYzi9wPpfKAIj3B4H5+EpUi2zLa848cFhmbPDBWCLvLrih7EVnfmP3A
iTGdoi1XPPYSUk8t1sHQTjED0yQQeEOTbMlnpV/C9zkD0RS52fZXRYJmc4CZo1GP
Rz06sX81bMsnfwlGJliAMY8qVs9Q1+cbT7OHwGaXebajxktd9S0mSos8wxATALeu
4au2nG+JI4XbOjFNcZgDnAq+TUqDFMT8oN48LPQTdmgXz8Ckq3tdSsNUreBSh4t+
+adojpSR81hz7+o+S5DMowSVGt9uQPzr/JIJrwX4MAYxsOjwfVAUuGRFzHb4HtSF
5lzzTv9Ht8Wa8rD6yDRJS0A0LqixNYBt7pGDbzorEKoAyufGivFrImRlY+Nj9NCC
Y+X+1ERwDSMKvpx5tEJUzjRx2aF8pCS9+9eWI+cFkEp1/io1M7zdxGqBQSJ+8mLx
Z7IPR9FL9sjEIHovSVAW6XtrOKMgkdFR+x+V8hbJfrZ0ViXCcupUxKYi7qu1YioG
WlbpEtnd1cpQb9ZDwwYD6LtFtSPGEvCucrWLxj0IpyMgexBe27BowDGa8kJOFhDl
vESEeAn5vq+WBKXGDT3KyWMqui+ZHvfdkU1viP4sHXu/aSGjyvgwmE8Wx5uN8nUL
nui1euv0Ra+NwdsFaiXIqEUqQ3AReVw9Y5+RF4wt0+VHV1q75blhkAqdvqpALc4z
VI0Lc7reCx2RuWoo9Hu7o8CZq1zfITPf3T5GXccoaXxbqklm83EmFp8lphwB+pqN
N8U/4q7I5F62LqgF0GJnB+GrUpMeZowyTTX4he3+vjAjEycdVn2yaWpOE8DQh6s4
AtnlgOcDLxiJXV5rrZu36kn1cIop7HpYzRTliJkfNnagq+ahVPyyo5cxBGS1X/Gh
FZOsbW1xjB96ui8T2GvondDrKQuqreiwBQIBjCt9d6C9DDJdyhQIp4M4ThZmCZSs
8SZdN/6yo3VKsBnXli2G9mCVCWYgfT9qmVHdmPRQKKOsYTay+XUl6PAgk2T9U+LL
opOIxFuKSWzgrc2gKuHdwq3wy94uP7c0uJDO0LX1Pev2RTz5TGFqWyi7WryUDxe7
p3i1cUJO7tB8qenzDwegmY1RkhteGrA8196gy9toA50oZxm1MwoUcnQ3yc+YNqzx
QsS7Q3hXit25FwFH2p/CQWYRHsBfRmf3SzXRRY69CqZ2ASmR7ihG0YP+dF25hXzv
3LAOXmLFMaD4reO1EbBc2IEJkWihnq5UbpPrvU6ZdMgVzMoTv8oN1HIWD8EUUEGn
17NsAvCKHfTJjeiEAqRqp7SMqff8bZlCysfSJwtyiQLN4B8D+AGFpPfStZkLLWgE
KMkVpDW+AUpmp56f8QYXyujufzKaSdU/m4bEcIMonSzwt4xRP/lZZiQDj3zpdDLu
slB29xptV5yM/rR7A7fv2BrzdOJ0Oo8t8N3M0u3fr++AIfVPuWLNXwlHnwfByAVH
BX+DrvT2B6v40Xc8PrxpgHyLAlHn8mxZhkNWlhk3SzHSIAPRhEce5Cgusn+aEjrE
HRCZRit//bYqCwO+Vwk6g9OZeeLx6t8hzMAg1eksbTBjpLWFJKfrdAba88VuPpX/
urqnWMeYyu3xc+R9K9WI7ym+c1k1fTkTxAsAjjcpxto2Wbh+YTLt+KA4NiQHwB4j
HYPh7sT9qUguUirWgdDqRkb0SBN2VBmnn9gef4N/5BPhQSAXqzNkbBDWYN+IZNMP
0cgzrXIDFKGceFQvBjwtct0d0B9QsT06YZhbWPxDBx+PQDfhR2pDmYoBiQxqVGMs
wL2FWephOn0OeDXCEB2yxJouJ/fL4cxM4MtX98tDbSBV3VJ2JK1XqfVSEiVO/8QQ
bq3lWO9UxWR3h4OjblT0lpBdJWeBIiSnAEhFcLBsxl9/gwjQfV0gMp0lnOnDiYZ4
K0WEFNFawmGGjmInJN2JNkoxC2TAOnorpGS6uRCeBZ1FqLMLdv709LeAQW4zfBPp
l+tN+R2VGvj3aFJFButohHACdc6wKGylNDriffzJR/hqybWUqv7Z7aWwxBJaCj9y
6Zzxi6/1B7/yODwsbXQQr5QdPabKSyIqHuvjpWSPw8cy8/g/4d2SLwC3gzW++K9u
yl9wrubBynmiPkKcKsK3KNjvFwynvTv5oOebXYkJMWT9RKSAQxJNNYrdmywRvx70
hpXTZEm2jAh/5lj5ifVg3aZhSttSbRucEu5h5YKjzUran20AQOEuoklQJZAjfMVx
Wgwi16yupXMG4S/99A8CllUjUO5wP4bwn1QleSOJNUx7ZoO6a80SUCfkyauicUML
sSh2Gx7LTELUP848/OV8SqGLGLE/8NIcGNKSBxy7HUEGH0nX7VdqZ37l8cN1Wd3y
fiYAFS3y/fZUTFMQnffcG6a6WmroMTd7f4RINAKA0/42s+HCo0Ek21BYC+dJ/kQl
6v130ALsUI1H4iVEPWx0+1yeb3sVOn+mWu9fbAdE6lJ8Rfj6xPgdJrrMBaIQ85MC
ZojD8axANB9+06nSvCIYm0FtfqwPje7xTkdMtKBQsZWX2z6hROUf6VYZDxdn8fzk
CWd9tmt0gQfi7gWNNtx0SnvdD9q5XtclsOzuxpCtB8cOL5zC/L0U4NXNYJ3ZTE9j
dJbfQwYgUdS3MHDvNzKVw5zDGKUnItLUp7kI3Fw37/r0lXptpIboBSKsD4KtNixc
7CTUQXPyWDcgdxvRvm2mAAFNQn7Te1MRFulZVNavIU7XRHnEaN7/RApztW7E7f52
UzilNRXxaA6Jfv83al6frp8aTgjwM2bWKRyHalTJRBFjL5XIb4mQ1UF1nub7hHVq
xukBtvph0NB5xeTvGTiD+9lLKL3BojOm1dNMDtPhbwSwPS7JhWUO+ECPMNXTGwiK
kRcajoL2cA6NXWTfMarKijp9X8QhrDB8Rna3O8gotiAw8ijEPT2Wvj9jdepneR+B
G4xOlVUMx4EFi/ink0K31G03cbJxHazM1TlspFd96cABwW2b7cm3gqR0viaJ4uNy
mMM+snWe1U+doXZizkIPVi2e9RyCiG15xmhaW9W7c0wRpR54EKElOR0o+Alep7E2
pxf8V4RWAjwIG6QQ4efoH21Eqq0IAlVt+AXSdk/GENvu4sfvhzOaif15o4G6zovh
Wfe1kj/b/MVavArrzlKGFt6U+7vyc1PW1h6R7JWrDJxn74Xsys943rSoNU0eDoei
qgFmNppiS/bq4ugdjifQ1chz28odNeEuJy72ZhuB8Y3Crfs0Nmr0l5Q0fn+jD/iO
9GFOroXbfyPxlkMqXfkpjfabJal/r0O6EOZZoIISa30dvjGQ3fLf4uRw3Et8Miao
OLDUKNkwbrJeOzi3bivzNItjCo3r8XTzclZmF5ShcrBILQA1owwvdWXo02rPWTy/
UnJWF5c3eViTNkOn3CLBeLW1bjVeZTW5KTmgJVI1V+C2UR85mSPnMOiY0hZHA7CB
Z/d12ppr56Ll6ToTTNSz1p9e4DcX13pW/bhFVOXi0y56CHIoeJ+pBazj91KuTKIg
PKJ8w9fGRGHC9uOBfuLDeQE7/wgmR37TJ08abtMgKkUs1J74obeic9QgX6F0iSkX
BVaJiHDhDZPG2F3eIZkUhgNxk7nWe8r8cuoYyAly5w3BytwdRONULPoeEmvJKZ77
et7zAlmUFqgdqhXZZsVSqdXNj9aCs8Sh/IMTWtwbooBO2UfppF9Pgqyt0QsC26pC
kGs585BCeG9FKHHnwwfmnELz5eMl13sOJ8zL+qHZP4OimEjyK11GU+Yr3hMnN4B0
sfONRV+EFnQIqVr4bagHPKukVlS4dVt55lnEwoes/3CzZtyQh5XiDBIJyvoXf5z7
fOLyBUZjMlybV5LjXbwExT4l/abMNsi3TeeCs4zK+PP6je8bclL8I47PW9OMMCPX
4mChFyV2ahdwW3h/09q0y5VyPv9rX/l7C0Sfiz7hnpS+YeI/9MrdRbYB1NJFM/0s
dzaDH+NYE4SmfusQstyIrF04WXba1TXsyXjvSmoVI0uixwoiaNQP/mNF2k0gB6Nf
8+FmWZa5SEy57K9C9fiuhMFcg3mggQQce4RlTse/vBV4atmmxuzBDBUHm0tRWgKm
D0mXhjhD8fJ/ntzr8K8mYAIbLjYd+ClWoztDeskZctsdLlB7cQYlxKzNwlEWeUIt
Bw74zc6HuCuL+zLzD4A/dDtcHJum1dnDq/Zaqj9gqHPXtxrd76gSp1iyQ/9nZ3CY
oEWytdu4n1bj6aogR7aN2+gcjU4wFXb0pcKZFafJmTjJqo4ke9A0AgnJjGC79uT2
knq/yLISU6b/VcHA6EvL8SUtqdN1c5g+CYufiT6HwLxwHczXV0cFMxCaS36aPa+J
Kert75RleJ+4IBo9ChMVHP4LSKXKItVhnJaRw8XGI1A76XfRgkwXc3kec5XoBs2U
LXceECnPyIJl3QYg2fdmzhc8Gg8eD1LldmsFm9CJZSVIyu1rJHH8UHdNq5GuEZK2
RhU/zcQcZOe/9BGQhudkUGJFkO2hfHtpB/8vtP1UThkP+tfJBwUzNo8518YZBy5Q
MRZdviXRGuO5oji76IWTwDQLf7RBsNiHD9o/CdSvT8ZMiCK+g49eqP1/Bmq1x1IC
BAfLkuaNBktwTH8JpIL3IOMYIEk7QtwR5n207kFqtr43xBiRdnzlUhiu6FDZDJuH
w9Ajz7GFYMJDt/0H8cwKs7r+SQB2HUiR01FNhE5R+pFiHlPzJkFmRZCXT+QWgCeX
kOUA04p1t59l6gkuF9n1GhBcY9aWtfLCW887OE+dCy6cOJjlKRKYVB3tDkIuuneZ
88x3aWH+o7BZGCuCmM6WkgRjSu66JTRB5mLEJbAOmT/mW/rsFjW6KYMJmzu//o1z
q8JSA6qNdNd6us2G8wM8FAX0BhEnTFoKRaVcOnR9y7zQzufgpdOXXeCXv953PmQ/
4NIx51VYmvBMrurDxZIyNlRLFo4st03KYL0CtBAxg33oLQl01ydsTrFhH7Zo2jNs
qFFRrC3i03jOpnVdKarNauedSF5tcxWDAaV5a7UJPhuphf2Q+iMHIZSo4Oml1K0e
2NEln+yyvjtXhI8gK73Kc5bOOXSwkM5U3fxs+qWUgPx8AwK4rGKVash6ofRCYdm8
Z51J+wf6SaW6WsdkndqRIGuWzhIz2eklJ+w/es4alJ7CEQ3rVvctwNMcATz5IimB
pVMf0Keqd5rLtFnh6yPOIcBKbtVETmnCFBgiLr0NNwWIzI2s+jV1u4h685Z2rjrs
ZL30CyPy+OI91WtbyjirW3+FSyhSzG3hUbDUtXUqQ2iNJXRTdRkO2yv8hkQAsWZp
PnZQm70TETJqDa7W4hUsq3gXblTVxLeiTnudD84wfXgq56KDCha0WRdFXlzisRNw
Lr7BH892PxPSTKBUvi+WxeOmw25N2rXp61PbwapsYR0hMsqO88eIvIMgHyLQ5SFm
My5z77nx/IcFTd+S9x+MC1FT9u9OW3wTJDdYKYRt1I7n2vD9tWrb0wRfOczF3CLx
IEGWuYrG/DSWkob2fb4zVi29MZVsOU8FmU5u4sSrJY2lcGz/VFHAvPV21uq/1nhX
44wrG3ZMZKwUoTKeuXQlAFkbKeP9eQRq/+YVW/4+QJIGmZaTBDmU4FJbygMflAfp
P34ACDzo7KXElZS1M+kl70LuxrhhpF1AbyHSi1uelKeNVImjCnzDV2g0MpFD4IQw
LiiP2XZMsrY8nCvGrEnHFjWj0mxf0pMJWTuCBFU4y0HYJWoXCVDCEj0K9keiKro1
Ox5K11ZXFQG+8qe1+sEMwGa1XLEkSqvVyQNsJ/RlrwdZXmvxrqVCNffaXWgz4mc5
IpsiJWFZ+Ju4OTmi0sjC2pdCL5TuNrSFlooYnDN8U9QOa4vnMU2He460S1OUgWlq
5scIrA8DOq7J2E3+icO8xrwhjdwxEYZDN3+BEERJuTIrR4FzTzc/FNW6VgPkLrcC
JyTPeHjgJHGby0/KQzPqs6TVyrWy6CUJG7dajLJJdn19PYmP9I7SKMJMevm8VmvU
MPiEL0P3XWbdgWcJHUlC529HS6n+OLQkzegtv0Osl5eEP/xrNg4KpJJEMoxQOBAv
2t18T03ijEFyVMXvrfkEQMH/9Lt3Ql0wY19ZV3uAMShAOch/uLdxZg5EiPYQZ3Wf
vuJf0FH03wRBH5THKreZ9JlNT1G+ZrrLt7xV8BsU2LrMtdXQ+HM24AT0BVsEVzV+
jQVbymFIOpi1jcW+wP3PQpwfqRZYkygFVmx6IpE/y7Ee9mabFrdSLuWvLCChsmK+
jJWLEDrTSK2wt6o8+unj4BNhDKsax43Ig3PMHYcSLS9dFg0gJqlf4wjLfDNdFOUJ
39FqjV+d47B+g2DuRnLqOIDJlhRvparQeTJL8u5tPz/IdFlmfZ8WA9wKR2939n+S
Q1jFL+QHWur8PEs/al6gB0FVGswHpI7ncc+vC5VttTnkEEbU9ofB8rtsiClYR71r
mB+PyvwaRBSrr9IHbjlxvzPb4qFMmAPB/IqrcrPCeBhV2V8deitozE+sMgR9LJPy
g3QMMFMUxzk2AFxkpi8cEeS4Hqx2je3ekakbpqUtLteo2JWXa1427bRUjI2OHYD6
rlv8PQpjg/OUmuHN8Xw/xOEQCqAgoQWUIKVEwEiJsE8BUP8YHTHZP+Vsgv+4iU9D
HNAgizJSIKWhsxqj3GB6okUGfKyZQKf4rvI4gkAid6RQWW3aleRhsdCKkNry5EgI
aoUoVV22bf3GV/cT2MNBcUxtmSwVUQCj7KG8PXsRUsH93tKVjZPYeMIQJqGlklVK
llPbeWMCdc4LDkRSajTxZuTYlimxnqBdAzJmys3RSzoD/3++lPytIs2W7egerLGv
peRs96RIgJ7CJdMQDZkTgFzRv2/qutukJsnKceed7c4lok08Nu2hCuocDz2kX9wt
l1BRcHAzfwpJo7/EYnWv0xQ4FhhCTubDrsYURNxF16qh88L4ctFUNh1Nc6PFnr7U
KkrTwFplUheVp4gu1C1yOKBvsuGbHfFckd6FsWC7t6WMcIHDxKoKtonEZfj+cOMl
XhMjaz8uU/8YTBK0wfy8CBg/nVOPff8ZyeTncvpqxeitq/aXCaMUwxmLTgFaIKdf
0hDF+/c5xS2FG+g5LTA13KMddGOylnCOUOBKxl9yOfmhbxGRtHG5UD+NgXVoMydg
GW75cTeH7LUBvJjpOdVuWSTX/IoOuz+wx7B8Udk1n434pSLz+b1ANXcrV7YRd8rj
708s8uMv/vYRyy/1P1Eqmd8MgR3lMJH3Y/25hVFDLabEP07H2wDd0PQJAaaClTpm
4/hjBHLVAU3QeH4hsFQSBzY7PfAXjSh68iDrQFBgmwzLS7YaXm7/TIKk/Q9ubFtk
h8IbtOpaJAVM3Zk5IaOvfI2paeTlgJm9+JBvCeJuMZaYztl6MPAmR3KQ4yfj9ZYW
Al04zI/KWl+MdIxlHCZ86PtUvAUL/gn2LNIpvojiyFnrOGWqWJzq3g5x0F72TdAx
MIQJ74dxdk2li6zqkE0NoK+JJG5fNhpO/jJd1Y9T/qBlIGAdudLv44zoQzJf4Cu6
Dqwdx8HXOjobxgNa27wWnFvmuF/JnMntzZltf/Dma9QX0aBUtc1g+8ymnjh0Jqqn
7rYsUT7VW2jpGi99rf4lY6PoFLWNTPH2KqHfzlRaCXWTuhYFHza1Ob3RPFUeiYVu
BxufPnCWUu/Vz9TXlwZiJkC4O4AsLHnsMcA1QD3f5ARhM600Pd44IeBekd94UMcZ
zvszeW8bnFLuYe1Clm1N3BxPG9zvW+8mYvs3zY37d1IYErn2r+wzlmjqJ7wwA5jB
nAgmfqYzQ/Mh4Aq3CQat6ayiR6SsMqnqo4t4FEJV1EQZnklYN4H1GbvFajJotGxl
JzvQ10saBCJBWwsUjVQODzHuTjOeXGljTuukBU+/J2eQIdyC5kbTVtsozVO4fQ2d
mvnfpOnvRPL3ytsq/uQcRh/Glu5bhcKRgMO9N4rzlD1eU7wjgdcduFvf7JTr6N22
FetBQVPHpKRKB+NhJl+7wLtJ9ejynn++b+Z/vEvl5nBRGgdgMFI1lppfCpOaCG47
2+JQDu5/VYlz0wLKOGAjx46CHTPEPREcPtViDy6qQ4nYMhTUmiMKW8QrbbQ13Ge5
SLpvy81y51RX0Ee4WH5ySTN405qUpYA93XMmlUtB8V+nhdep6ZanTwmiiCWRynFa
HZVfDuTyUfvwuGRenBxAmBhKLdyP5XvOxY9cXci/DXftf529uNvG0nMR4rCTghop
/QnR1oPq+UxwmWbVUXStp1Ru2q0dRhBuI1T1JSrn45WIZ64cgqEhWMgZcjykUVnH
4n+dPQzICNlx/CMUCSDjPONaLeQ5IqDz9ecrge14SciyX8/+f96IHETfEkmHgX5u
oTzjmcsX2WEoeuysYyk6LneQmlo7AhpBWDIhNIOTSHzy1SlveJ7mnOyir6ciB6nZ
PERUuYti28Y7QpYm24ppE3M+pS1dFwVet+uZTfF9eLaHugKA+ryPT2hRvjwEGT2y
LCuB1ZhkmUsrOkXIeQbPOpapMjwjjpcJrMYp8Fq8Qzp9Rqgw5hxIQOSTOpBwpj0N
iQd1Q0kRpQfCIwAutdDRoU9sRt8qr6B/r8ezYHxIVCTPuxbkZkqQqtLnWu2aPrv6
sh6dlXyztQi1MycXYN6A8X7vF3JFYk8LTze7LEtH/8FjHpJgG+mmQC4DRIzckUAg
pGjgEPee13X5lUDnSYn0O5fq+hQ9ZhnwcYt2dxb8rDcPR1fVF8V3eHGD8cKcYQ3a
DygeitFfpesOpezAmNepAWyhp+TvumBQJHsCFoufdFZPjPr2r4mRmi71q/AxDHDm
Z8qYhMwNgg5t0WGamTasNIpU5b4o+rSZC7/UV09DaiqNSobHCkZk/4aU4Z/5TOWg
qxAGRx2eOjeYHMIIDbBxbXfT1zRDyalHrMXaI+c8J6YHwtLWjmrxtsDqObEbmBNu
QMviwubMRxKmQnR6B0xQjvkM220+84fLR4p/mLRIYnknDxApe2Lr4CnQqaugPePY
wQrKZ7nlgOwa4sZiVjM7GHryYUrvU6USSFK6S9T/PhaecLjxLsQH4m5PUabsFhp9
gE9YYK+0glWmB66Oht1716Xc4x97m0W6FOKou3TMfuRflWICghEFVbF8KEge0yTr
QSdW3OJ9uI8J7Lifp7yX2W6fa4SrZCPl3KS1IFoza4i3x0914rtN/Z2voc62PC9c
YVx4mdIsTWSghCIlDrnGRjQyWlg+h1qVbnmnUgNKxZZDmdZ5JAsIboJFymI1buc5
VNyjK6aibVzMslQ/UGp6BgCcJ2soAzTVV3MkmSM4qQ5xGI12Dc5UBPrTPfAF1hkG
jP+/6UnHPPXPZMagrCEqJSuODNnGGBFGE9fHAj8H/EXU2I2LkykLppmzGESRM+bB
2L6Apea4bXl/6CTKCHxw984dQ245f3goC1Yr4iQ5GUSZA8fc4c6oihFmeV6b4Uu3
L6lodCunWWOyhDchlOJzrQtvc+J4+MaKPKaevR20XlP/1yDgc8ZtAubOZajDes6E
5jzA8IwXQLtpboxlJKaJDdNopK+6vuoN/TqkZ1aeiLNz4WnoT7zgMRv8bNstmr+4
ReqxNFFyEyXkOfaRF0O3Q5vK0FkavKy1/IaqUh8qwnMXaSQc2r/hG7u884IYoTco
RmVQsVHkXM3uCohPbjDAT+p3qjQ6Zb+T4kKHdZHhqfYFCkAPlQ2z/LQNuctKhm34
iwgeR/Xp5TZGV6MRedK28pUN1RGTSEmOHitRw+6RO4QXZhk/iHP88AT9Q6KOtO0f
xXrtM0VP8hLFOTp2/zMAW+lLGneNiYuY6WbSE6aMBlqUvbhJpsnqBwtEAQy3Bocp
Id33JNyScoSlJlfYM/SIcp7FvrC8gk6XvLJWj0G5YJdYR3qQ0DeTH3OJ7aFQcH24
k3AFFfwXE1jFkV7P+ygMQU5t5KNzamCnToVnI2fuA6PemrSj6tzInK07dKKPUBI8
dggR2IF1H1gz4bg9Tl3rypD3EnmaEU7Is/0FsA8/r1/tUmBqJU7OFWk1WbF6fy+L
2fSzmWZMiPP4XSlskh6Fuf36eVeAYAhtQ1H0iKwucbAtmYPolEFJa6GKvEehcOEy
sJMzptn5TnSOHJkTLFzJdni6h1LuFX8A1aNzQazK3piQN+akGtxX5UHBblFuxr4Y
nqVVpOjnlE1AR+1YGbsiezrkm+VISAZvLcJEVbTyqSHhQhA4uc+YHKRCxBH557G1
1cnejbRwet4if3Mizai43R3wiDRTmYjI4jV6/PjNDjO8Du9O0162SkF1ALXctWKK
Y3DLyZbiBNyUTUbDKKthvv9DNQxnCsie/+EyTN/81HYLD6zAj41R3G1qxiv3TzjQ
+Wv1yHoJcRAoyGgpzOoDtzvBTLT0Z6cGJIoStt17NSAnzH8waJfii9B4cQN3ZvQ7
z4mfEogMxl8WgVfe6U9kdH/ksR2eSW9eU1W97aWd/eWjqYiG8BygIiv6aQrs9FDx
Bh+KrFizCI2qjju7TgVJaR41mrUYYs1SzW0MiqkrGNCy05cy41RIf/OecDHShZ+w
Mi4EU3nchIeSl2LeX0qdorj7QEjEk28pYk8kGJencuJGnYDsKlVUcbXgEo37bM3Z
DCRcBy2LIZwUj4GVQ7L+LVYRkTIPE0fqyjBfxpoXjONAbMVVmlVDh7yok3IWoy/c
PfPhppDrLGmsEXlTksMH2Rjas4iLGAYQnzIO2+A7FHdZDesghyybsFzbshByI95p
iU82f8gJBVxhwpwMw/x6J/CcXOznXPZYdc3XdrZuR0GEahCf+3mktHg4AOHddHMI
s2FWdbW8LLXpQ34S0PR2CTOFyAKuHBa5xqcQLybzk57CYFmZfZgYoUZwS/LyN6oz
FSThE8AQBgj24XUNkp1vsrJjH0kVwwlsKmoiw1Kw+hxsQYFSsYuTqXaloz6Z58sQ
1CkrYnbB5xdmIHD4q28SiI5EBtRsF1azzxHFtrRQk0vJH6fCMZftc/+gxOyDhPCI
Gt8GBf12T4YCY6RnFdvsq7wzurOumGZ+OhnXtDgjoj/2pwzX8DZMyfmf/cVesZ3O
ZtFsHpDsJ8GdWmU8urGyYzNB2xp95/B/w87nkodLf3cKI7Ar3tSIY0O1kJfoGuUN
awy2L1QBo+kY2GNXlfc325hv4UiAmd8IEh87+pA9ZDjJys0sKguLNSMjfd+PUn94
r+oNrifJvftka1xHnhGpBo4pE3gPG3y1ZwSRVMGT63hUgHSSPSpM+ccaJY2aoYIa
RmUDMCW4/Lj5iN8adlhH+lFmTFQFZ6cfhxV446cIMuIa0zt3igNX+pkxJbINvblK
JbRWcmfQFD5bR0pN67LRHxjovNgIXgsljjwcludSuEeIoshdUzTeFjETyxauSNRs
6eHyxHCGt2jpprmxKDFu2tOwQ7fqNV6KT4Nw9CfmCAxRw6vMEJkEsxS3nZOABTmF
TG0qzpDbApuou/fsUd/dcvOIfo8Puz8udGeLynY8w21NFAtWoAGqwRp1uLxlV8Bh
/4aeKh0F2WalwIrfhUiruE7Aq9hhXqY9IfTAZ/SY7EpeQ/ui50IKQKgxJy31wcPy
MHqDm9OmAFT8plM8mkDJGrgufo7N5myKN6mZ5ZFrXArkrgiFDfGu0fDssSkBN7eN
FS+DU4di0n4LtbmmLGTFir4bohymLT+DMrJUbrMyRe89FMH10lLa3CdPLdCO5LHj
lbpROLXwzZfHlTuUjDXFkB60EqV2eYxJolXgbPyeUaRNVc3Psnj5P35ytMC4kgNL
LKSl6s5Zh6mrGWLkhQEajSBXbQU+r6uZBMsiqHxUBq8BdeyWCdhqp8UhBYdD+fGI
mZBu9A3q5P2m5GgPeXtOX1h+3KDz4TDz1Is0+CpALNLKvuDe/wCXcCKvHmsK+E81
szj6BFe/FxsjoX3JkQodrF9MhMtNurVRfNKUmy3D5F3ufrgCDKYNI5kf5KsmaH3s
AODRnehwJuUQuomVXvTZYubnQX8inrwNiIsEiL26+xt5KAwS/pq68qOPB+mbP/ez
pLO9CvJ0WOu9g8sczT4P6e/2JAVNiQ/QSfEsQoYYc94bk2Qqcuz04+7jS4XgaF5X
p0eQA0bUGq4UYiTFSr2UGCZGoSpSmAA1OqoVwQZxh1jvsh1ykuRfIUx3RGR0cFdi
3l0fi9P1tMD/UiLLdhSLTjWHUIzRdkkW34Ss9yV8MvQQ8uXntjgvDne9PnfL8ZoN
rt5dD7PIq0V2dzwTdoLe4U22yfsCi8Q/SopOzVLI2yTWpBVGofxcWExk0sBnAt/k
/6kZH36YaXbOPFC92Tr4i/LfGofTELKD4zP+1m1HUH/VhWlmk7M62/gbHyWZfPg9
tGEmGdF82vcItNcib6kAIyWqWnI/+NKfKGj0L7/aarMD+Q/b2aQfaklY7mN51ZPv
e0x3ZFgrNF1pNCCnUZJzYRFERHWL/B8JyOpeyxBAgdhDN0Og1C+p4lPoLG7qsBXE
VUYu/AVFDgEhEFSsF2wn+RxRLykpAyDRHy1hc742pyx4bh+RojqG41GPiXnbNKzh
9lRuiyk/L4GHpjkz9JJkJlMlPdLWEFFlFo6QblcdwMZG0hSq7oeMbBpU0acs9NxN
gduAWr5DG9QmW72LWi1rzpvQfAjTvVReryoSgGiuRWzWag9oIS5YNVnE/7PyZWPc
JeazfX6cI5y0FiW/+7zl1zdpQ26rdeQEw1mkJK6U/zNc/sJiGX5PuHqFlFHa8RBH
GCZrSdwBZaoJcBAy12ZwNqvWKNQlDT6MJQRAjnOYZwozBl/NS6npwM9fykYy5oEH
9bJdiAD4kbjkXrMJaXbE0LnR8lrh6PDv847oLMmyY3t0cnoLUF3AGa5f4E1Wen4M
6cN19denoFHKQyrUiJ4vldheKsf4G1sMzFUbBLZKQVpCeRJCu5saIURpr7NHQ714
n312PLGDG+yGE1/PxZhdvGtbEM+3UEZB3+RGJ8OK0adXxeQChDElo6UYOqqSCE4i
7FlQXXIFmWD259qKtQJxzfVsFffdGvEesfSywpfG2ku1wNNjT7sA6KQr3wUr3Fxq
hB3BhxiSeS6vbtnyirMJqooPl/wfNgAYxYQ2GeKNtmRFrGhsOfACW3HiQTxyW4NV
9TWef0+YEtbeWod/O/LBiwfzrtkYuUxSHrRqckQWDgEJySp+JZOJHH5FQ+OlwgVg
5i37zRM+vJYv6qXOSMFR+YYgDeitZcRLdAxXh76tNXsI+rVtzwU2ieRU+O5KYC4C
HKkbEKft8W8hrQc3FSqQNd7fxiCEZoezpX7Lrl7PEk80nh+HkblTLsPnqAewQwUw
1aP8l6YERe1UOAU9hUBUVIdPuQs4J1aDj2+nQ59am1r6rtYYdcawni3HmBbPiPlD
o63MdmgAjBQdfdzyw9MKD9W8gWs5x+u9M1BsmBoAtgA5aZpPD4ZxNicS3ajlb39A
73YMmQeJ/8viGTHzuU6WLWc2HBGIzoBuwtZbKFsOq+82iC3E8+8gCUn9E+uttY2L
8HDmyh3K/wjQJ9ZAlFOenWoPhJiwOMZdpU/IfDf6ISpjQSxTESicUNQnlMBb2Lpb
VG9Y7NbNHPHDfSTV7kd2xs+pwA/bdY54dWQNk8sWe/PR3Qpzz/b5W4pXhjnNBk7h
Fb+NjTFryjPaA1FUtyfZjTLoh+iQYtXI4XLrH+OnL+aMiUcxR0xNSebkndrbYCu+
wg4pEnXK1j4yopPxXiNob7CKIcVapT2v5rcjPNp6/dc5OH0Qi05CpgEJ6JPpZeTf
+503YD5FZu+AViuuszFKP3nVfbtP+AoCzojEwVXF+dH53HiwMSvKzULPmK4TsnWn
hbwWXJFQeSStR4MT+u8W300KOv9XJHxCtDex2OufSITJ7Zt1NP2pdiaxt5D+4Phv
19jR30mnn3l6PQ9XHA4r8LouT2kwlCMx7G5aRmG1Mud2+5v5z6dYXbHpHy0OyQDE
Wuf+HGG/FSbg0AyMAEbSZMJ/wbIkJJ5CTJEKUf3gWnQMhHB20U08c7916AVKXoJi
/j3HDqNHU9B85zlMUaaRgcua35vlG1uEH0UMpPFJIN4mZyD5cBixra1mijjxevvu
vz96V8c+quUkuobC+xcz++DnZ7x7nasdd8xDDrCn+xRakPfLqS/RHTtDxfxKSOnr
ZwKtnHrTNxhNhxQ9UfaZyt83SFh/LDPGozFWPElkokHSDEgJ0Ki+0ueg6QoSrdui
/vW3QjyYKJB7gcaUeRJJCJ9iH0MqjxsusikFAWmxaeqZa57nYRBJcWxtsDi43F/M
k+l4kEmN22YnzAXNEeDgtnbworqaeipBk7JkdFew+LKl5F/Plh9q2tdnz2exOKWU
0+CUvDDVwkajiAGb1ms7n6VhpskEWg/iFRbbd45jbPq3SOT9p9xkwgO0AHfEsl8n
atK1ci45HLrzCmVZHzYdlVZWgoAn7gCHHZHFemHb2/wFdFnGK9KGy3EHQCKnVyeF
R4oeuE24r/LBc6mTf0T2y04krBGGCahIJee/N+8mSsAbIzcY4HEIIL2lNQvgjnWG
ziLfgo1rac7fkjyw4y/epcgHOJQKkhftLx57ely6P8wTfsuDphYXVtOYi4o9UdpT
UtpcH/n4jOtrAeY0pKqCA54yrjnpRcs7QNro2E4zkbP9S5ApNE/BHPCoMtZREmj4
H71RNmzKS2UjBSuasDtd0riJMN+cITX07vADcGXR8EWBhCurkUijYKNRvRUM8SKQ
9F7muU3Ud4nmhU43hXbxalGRnmxOeJP/Y6Ws3kfGOl2yFahIj6PtlX5xp+uPTGgZ
8dh7Puc5+7HfXjZIP//o8EeU5sZ4Le60LGEk6J3yi0pAw2q1N57tGjOnwpuQtQVp
X92IKeIPcNGTfZ5U4qu07SCQpiGmFuEC2O8gm2H4FLHExZmPvqnBn4H7Ph/TlzxX
nNB5MZFtCkxQiBcUDJ7GooDcs+l4PRjAeRnVQjCBhtPAjUdnKl+n4crXih07enq0
8g55zCWEKpdMFNfI8Qb+AqR+jr40Cc2r3/4C3vnvWA11hgRaBJb6JuErzzCT53qa
xai+sc4gStf5NiXnszx0JDWafMkMGWpr0VGET+nq1uVkqdo4dHDAgs9JSbIZvh+5
t96D8d9fNVrr3dhA4zUnqx3krzCz4fklAD3JWc6UHwZv4oSRL8GnXuqyoezUh7XF
/75zc5KeDlkJOb2KPj5yA8JEzPdFLn/V1UYs7F3TahumnnOUzHXzxeR9S4t0IaIl
vyp+xTvhy6xLUVAXLrie/CqTcYXxL8GvjBmTz2/a4FCa7lYD6oHhFhmKoWdgMSiX
xS8y7Z9YhNKzkct6zqImAXAYNZO5dDbxKWM0tZVy0ulIIh6jFVBojUACTbg63B2K
pCNi34YPOFVY58rP499uTaGzIuzyXTVHuYJlfrlLiu8PqgY7t39JqHeoTjNiFfOH
9mJh3YvjVz8Y7l9Xc+fLRGgTDukoasTqsmRQgs4UfzvqOc28zOr4g9OSonSKiq/6
z/3weFQoB918kSPwAWBr2IsfZ73HA4e32d5ILCS2lfXiCnrHMzsHSh3Z9gxW7Y9o
/qJVwiRF2Sl646lWIc9/xGYVDwKgTs2TKMuBnapLsQuSEA/zo4C/339aaUMKhBLF
6x8Rybs9IZiykZzcIYMVh6kSMdxfeLKXg8B1IB9pe8oVWV1jCTPWo8gB7V8Dqt8D
nLYX36Hki/VTEP2oXcvW0cf7NDPQa3EdeOYNs9cbu5zbTyrpz/AsqMfxiTMWuEs0
ZNl2WU+pOe56gmKkRStYRc/JiJYe2bVNDMSv8q0EP22RmaXd58ESdSR+jRPAOd/f
i6ouAPHBZ3ImvVoYPRt2oxpESM8LZGawDdBrMYhc4GYoZowKnRjx3LONKIdCfQxv
yqbpS+DAN4qQvqm/Y5jK+9jzR5n+S06znoIYZostBWU6biYOxVZrJ2XYy56m1+VN
VuU8Dm4Q9pm6TL9X0I6HuyOKg9rVoIlb6GLiCo5cFXRu3gIsCXG7pNpe6Oc/rxSi
bogPQFAKQiANiiomSSbLb7E8oiwAFmFLgaJMUAjPJQvyTbgCedhBZHanWNBO9Y92
vir0f17oky7iRI8InRPIv70q89V5/Fi5XikX5YzMxEKlMwrkufnpAERwoOcsi6wt
LlF0qAapuu5yKVfNsUujMDHtg8HRnzSUZT3rBb2QGwPVzxMadZDV81SvOWLlmHfI
tkvYPN/tUK2e8fH8n4gTSfx5Ljp0o5w6hq4g6t1uD0nKQOgdZrzUxjjKB388jRhC
PEqWkDrpw/S057zSTgxvrrk1PW8NtkPmALZ/njVAxm3nxZUw1A46dCTaidjxC8ph
Lh+nPc9zXWqJheTqgC5ObmUA6iuRwtxeh2uRQqk0634zvTJYqFhS2/0P+s8iAKRO
QqeSRJIougFH/PJk0VtF/9GmvkT1Zw4JX5EmSz+WRcRpELdIvlyFrBEhYiV8QCbA
tfFeJPVXlfpuzYJdB1jnTCMQf4j0W7v8KrOaiwxbfdklAlK8U3/OU1PxYRfmS5xC
b4+bp1Slnn9PuXyLbNEw3QOcWFp9kpr/Dc/sNUkDAXOrNarN0dxJRQa3ARk3d3ki
802Lm7COdQ1Pe+l+LMveP+pUSfOK/1Vz18m0Oks/NuCZOHvBPwhYJxw6O/mwSJ6L
F4sOtuXe7wn/ONQnJXzECNbxHDk94Yhufqm8u7rLX50LcHjw5hJy8nJydwPaAfvf
iHVWtFPnqpNTUhEM6iIkg+EGE0JQIStGm/BLFfz6NCCmE8RiZHLyb//XxVePk5Ak
V9uPzqhbZJzv+dba/Pmv0IWx+Hau7OnWtlgNT0RIX8lQ0gxeHcq+Nv3aAZkYmcuG
PNfBIIXV/7vvtr08RwIaxRCA6UG5516YpWhcZX3mH3lMuZcSiSgfWAFnXPFvhKXF
x30nI9pfnWCaXmKyE230ByBYmeQMK5zaQoEDk5gJPqveccjgx5425nRZ6OGoOLqg
7zU+nTaVsRGoJX5oCnQMi8OU2V95RAXtIPbVabVfpToiJqFL+gRwERfpdQbaMMXe
RezFHERV8yJ4bhXhsb1dVGCv27pHt/Xz1hVsrWtTWep7TfD8NX1+c5a32V5a7Yd9
E6twoF3xgIRbpMkkUPhTEGM3UVigxHnJ1Pr8J9zqFGBXnSJ1FU/zWdXRZwwCaDga
ynX2hkeHhNHZKKFegrL9koZ343yCv+k0gfftbsyBLgFNiXHE7hSEcIP2uEb7ns3e
ekcX3JoB+qlQ6LvsYE/Urx1DS79TGLl3mwLcGXFoUfYvuILuovJSINavZiOd3IA0
Dg7nf41iimPfnStLXKbGquxiyInwCt+iWIdGdLyZdtf/8WAXH7NQz1C/17XvA8wG
Zenx4rleYjvqrDN2rURGiaoYSSggxEU9/1nDHln6BpodkZCLNQRipG5zNQJrFIJj
jS+G4GH1C0cfvVDQuSYJ0k08wDKY56zlKXeFaVKkzcWZAtFKQps0jmNn9hJ7Mnyl
7iACqRk+T6UJxA9P+1Av9TCRUWzLzAsGRE2UkZT8llCh6cm2GPfZebZ3V4zIYzkU
slILwrd9jxa3qV6MOVLjVRps50OT9RCgtbZeOhQZEJJZWYLFI5zUjEOn1yRBCaFn
cXzSF3+UlxTgN3009p+w3j3SR/ilVybaITCvE9qvi1/RpBLXLP7ksIQxfQ9v2tFX
NmZHNdko0ETHIFJ9aRYrloRbRsZy4kxN+uAX4C5hSQ+IDK663UGtcR9kNDU8drIe
eKc9wONseESbO92eFOtFM0IVuqDcZGc8Uv1GnAEFXJTuOHsecAzvSQcrV/cisHGb
Buo3gPWYJsfnpvBxyf8WBQTwUS90gRXoTYvVdDqHNsCVE4Ybwmhv62BLBvEP6Ajo
iCRkzX7Iwhxo29mZOUeokh3glto8pxreOXBW8t67QTfeJbTaAW+xzCDtZLC4yrAt
DUjg1OUiqYH7BcjMvchArNFOPSWeM2vRZlMoCt9v5ddtmmMaIvQ6aG/hIjRqosYX
qNxjn/0gpnCs8uH3GTmrFYUgZH4oYWZp4rNjCq9c3FcFcwQsyCLMP2VxAT3FOqhH
8PPJ5EkCdKor3RBFCGh+lTfF5cN4jjKfbSwgNxUWkxtW0cyvHpiH/Jq5BPK83F7g
q8xPwWqKFL7NIcuQNOrCU9yFNwayBxSYzYer7Zrw8ppeRzwnD0yksn3Uhd0jCzRT
Wk/7iIEQAByu3jJ+A5tdfxShjeKDm1+Ms7ngrJY1d3dqo1UNxg6/LleFTiKSigYi
zXUKhQouqf/WYoZMjvgFJHSHv8Z9Ss3DlT2dsYx8f8DWkncdbk3ODVvl1qi/5fza
LaIAVm+eZ4Xp+ZS456gvxT3bekNCuvrhkoiFzYzFBX/v1G2GkaY8AjHnBos038jH
ikqm59YfXiMVpFSJ6Y9aohuU2zBDgpE8c8y5RU3VNvnOljQTSarleUCXoR5Aqvz/
f2aZT2/hP8cgnVeZqjgztk6sIxprkp7zzorK79kzWXzABgNRKm7kDXQS1iuu+Ihb
ecnc59Fp/KGEracPsbARWdT9Jc9Y7ovEpCVdRVt8lrYja7ev5fY1xLVcT5iQNaqC
2+AISowb8FSwqE2c5Dj9f7YKvBLkVH+vPnZ0KJRUlcpptl5xq2zNU2tP3Ss6qHOG
wQOtVymu0jkufzc5mp+xZAQOiK/JiyM1gUV28UBwiovzVE+YEN6P69VMzbbGppi/
mwfxgcw6ss+YGXuf4heTkBGsSHpEL5zvxhDzZJAxkDLLvj+bCQ27OBrEm4fPV/4t
Rb0XMw05B+kEBCLu4VLzGvWLQdMdUk32jwoXmOQjJ1VNabrqtNqxUtMU+u9F02oR
qbO64y0PuKBtDQxwlTiTFNKAFeZ/zh+rWbiZou40Q5X4NGSIAeGO2elTrcH0Qavg
oLB26hEPlkSIH5t0U/QGU6NNJkqWE94d/oIp5nbilCe2IhWWEZ7F8fwTKfGfVWPP
LtJZACMMwITn+pqagETdcJj+uBiX0elusz8rF2jJGemii/Uyraaa2oX+zoEpgIUG
75Pi9hkehqKKU8dpwl/8K960/I4dUrC2Olgs7z0JElPpKDNYi8aQR6edFfERP8Yd
t4F2KhIoVg+9zHv5zh3SVduJqrQtD3XP5o6RCpWzrTlhYqxCrXCrT3Ac3o5r8oec
EwzydOo2GlA8f0OlLD4pvTktuwS+2ZXefP9ulXUz6Qksxrq6vLpin9kUIT6hby4P
YBeuN6HB3dBMLSDDEV7JLz8/jDZBeL/qBxyN3y6zZYiBRAoLlBCwd6ntT5O5+M5n
VBMZgnU9cKnyNU9dBHZJWI6qblS+228922wWGcP1hdYsVbrp4KnjTb2z6vMrByAj
qsiqK77XT4dC5LtN0z9S8iE7eDdflXf91qde1/ep4EgGsGBJ50uQRyTwL22edk/l
k5vsf25RgEpqYKHK848cCvRZIRK7eDmF+k6PLytU4kDudeGND+LNyD3FvNN/9hxw
mlOGyvEIyXcZulUiinlkqhMYQyx20hz2IvKAOkTTixVql9IUM47RBJzEDnGnCN8N
h9ba48McvYV7bDwFB8XHRo9yg8s6qOJVUXdaC+ZrgHX/GuUSEgdYPdtG8v9zkTya
L1seXYyyxJnKPKfCZXSy4iNAmWevj4JfEE6Q1b2TzrCWjG+CS1DeY4DS5vq7jz/A
fa/+bxdPQSzgXIneLeAbGl57TV9J8ZzY1qJwpeoEKORQK7V4uRD68C9VkFaulspE
kpPZhz6Mhw4zC70Hr17RLQnXS/Gjqme7V87/iktLH2ifrpM5EQogHhpLr65jfHP/
1sm1EsNhUQh6sn05sTcjKRBqJHEueFr8nlPWoi4EWCCaEn+Y104gMEtLqyKa8IZd
q91kUgGiHbOQ2rvu9g6KbrKHtL5qU88r/weyFmRA642EXEbdBpe+5GDX556UuHNb
QrqHaNc7D6/rqpoFEiihfzrzAAe4IyptEBAHopD8x+Q9H4EXut60hTbMT/kPLNAC
P7qrG0uBYxc6leUGChHdwIbNw6j741aomgPrYS4mTlzRbhkP4n8xM2rqObcPrtMj
n6aigEgCTyEtVHn8nPug2dekEydUhp1wRKpKYYqGu4VJVqh9KRRca8cjqXWXZN7z
l5X2rSnbz0igZ4llcWygdoooVamZXtQWBNxFoo7kjWRYF/HrP9NRw78OZN/IBWt6
iG3v16DMx107WHDe1I1BItdJHruOZ5hGlymUetYJUc2TWifJuQRfaTxtxRTN2U5z
iZH13gS45CGnCGWbmMnLruwThGoyUHwaFguj6MCLI1gxUB5N9BNSkSoZseS5cAp6
PbVsnKbEgt+f4l2GvaOfhbR4Z3mp1/e7GmXIDy64hBZ3SyN/u0o/aUm8ZZ43fhgn
h+YnI4CF3MZVCQa9rcwoq6czAdRQEKuJL5W/6Ki1kUsd/sV3Z1fhkNLrb9tp1Y6q
kLVck5aykMi73IbzWxEA+FGK6uCTTqdCgtSQszqbFvOMqPlSC9TKaWOWrnZV+e6z
RhhCx5siOKE98OEqP+64A68JLssgZ4QCxk6b7iPoagtuCNy6mqJpQmDhfeyPNgkF
OYmTJs/DAe8rzXAM9ZxE7pjRYNYHLyHQuZ1JvebAkASkZA89J1sUgglaeyHlB3QN
2xr+MC+//GT5RCp+688cvhJ3/J1czxsKXZeorlD1bLL875JjJq5HuceJy9ITveZd
rotk3CxSnAM1OKDFq6tftEszV9vJO6A7iHGPmXmgMfEQcf7arMf4QwZ244NSdldC
543Ij+AiULfIIXhz0g1WoiafdxYkqwHFQ1AS37dM9cDk5E+kSMH1Uxh9Cv3AkQgd
477MNm+YrONXFNhOePyVme6dRSnWl7i14CZO7YU9/MX60wo/QMwjNVYVBBu/aJBy
UnRRNEFdlBDgTy9w7NKAYRIh9571DHQoq0m4+/j++0WENxoJMDIketx8Kuo2Uy/D
vJdBVY56LmsMWCa84QSPKNx5Ofjff8t/nvTMjk7T98KFF8OLnCcjtkhVOG7jRlJB
Dt3YxoYn/gyJQtAnLBKgv3PQOD3avAxUVkDw2rzU6hWB1sSMdKNov9qwxbGv4xse
zewqoVi8JwQBAznQncGT/+6DxUtz6D7s9vvnoVOrTqrxBsAU69AqtvAohoTAVVUT
8CY2/46zrBXq3Y6s6osK70S5w8sIaVlhB7CbZyMA4R+xoh5xUIn/ZF9Ufx/Kkpjz
tdpYZDqkZTWyS8JvXkOEmuvks1VRIUKenLEnAA3GSWi6SPKQYFIZ6k/rcDck5tg1
TVasw9xolmC+tpxXWat1lkxbVGxPlcFaFx0O45grj4CJr6uQrq8/cczeBW/2Sk5Z
h4zJFzKeQLc25QUHB6TtbhLY0Fg+CbBkukrY4HsRP2Ho3FH72Mp6lkdiL6LswpYW
PGfMqFCfXueezeNaRh4L5zw/1C+XskYKuDgjwBKjfHiEQ6Ttegve7I9ZU4KjAO8k
/nJQZxp98YQCSp5DK+mT3vWV4zSgcLDhAfLcjqFQkuvYQd+PPEA7AwjUelovyivT
kDng1ApzCPYS1H398y/Q/hmf+hnpAU4RvbopvBqXBFYDOXhqBNoYZZgsy65l8BCA
mVIsNynnbyFC87yeHRItQEw35yg+Av8E84X4xMNQLeAqd75rBONziycsXKyTkcRb
7UutrImloHIjVockfKSl93MHyx80Zh4nPMZMGT1C+OgLkNatkPKcHTcGHv1P5azh
WJyBbLOSv+cYvtjnGAL0JGwvkfMywmHfHrEL+3zVgzj21l5kJl0+U7KuyYgVcXsV
bd0VwwG7ulFCut+dY79P9Tba7RBCC4EjKqD4PgG9u4qLbto7Lmw+oS1dJKzV/On3
COvJwaAP+yCN1EeO1ixqiKoM9SY2fmBqNFRZxVJpjp0tpxY9IbUpCDNmMK7yPOuh
jVAbzDA3HzWg2Rrp0wiDVUCutBwCMwXEW+tvyZXUESLc0Ylo21KTXXenbEOYTZ3N
F4j5aZszoR6B9RF6AgYs3cGM7OdP+KZGnPN0gGNIKaf6kCCpA9huBOOE1YAQe20Y
WyEVo/wzRsciS8BGTZV8B32QlIbB8gQ9r57uUkxXZzYf5m/HqguY/Oi+TYKLqr7z
6cQba6k3gFp4JMrojMhJClKMoRwGFbRSYRdZmNKgRbgr5sGWrxSEIRbih7cubJbq
WcWz05OzHgJ5nUk2NlKJ0fCYZ5A0G7BRIg0iSiwbcLtHgQZ0PdSoMIDSOCPX95WT
jYHsb8Fp6+taWtpdwcDec9QnVedlgHLgW9fIoDSDGhov21agm9prdfSARBQLdWps
c+4rPR2j/uBAHKTNiSYB4Vh3TOGrXd6znIO5R+iu5N19nwvC2xGQQaJG7OePcyEO
j8BA8GInjLtxa33s5aCsY4pmmHLgyEZradZO17UaHIk/FEYZgvnYMuXa1kPOFwBJ
/Yl4M9zW0IKSMg6IeucIZxuo6qBf+hiVBF30c+FL2bOESTLSCTOSnGvZKBjyaTJf
6Cktt5xuqmYyA+0u3sfFnzgu03UIsg3sGwxqBsu4uxLW/Bz0HqQ707bBTuMu9LgH
CNoGSIP333chHrUHEiDdEq8eff7/QdIQTcPrGPmTO+ruajSk05vwF/O8sSkzhfba
lmtrDwqfjyF3Odg+Y5hZ+09tPsdMtz/7DXw1o6ddJelqYfSSIHy2ekv36wBM3XsQ
Q7Dn6v/9fJzZKzdK7sRV2BqJhRjEcag5xlSEcvhy/2iDIf+aifT3UIg1K3Op8B7x
GFDZvUS7uNDU5V0ziE39dvz+KFNsjJXJNjlrz8F+F/DHKSk7CnPT7LBjvARycUBH
/qSe8lCKaYiBpfR4fPz+Z1tPfHKVCYZ5Z8zvXph9U/hJIxiQRDOahNIc6URL5/HA
jfbu1VzORxUI5gmciQFeKK1IblLY9hK7blC7F2xWVPgguh+L5CrMD1EdXb2Hfd5R
7y7+p0Y51RTA6SAvilmr2Bmukc9zEadxZZ7RHek4lLtlybQXMeW25IJEPyGdDeNh
NjnOG1Lr1sbf5yMcTbg+ewUROxcl/woeQN6UqaA/ijGUmEwHR2WgZk8uF/lKxSQq
6SLDe18BveQXxXBaCoEydKSzMfaSigqFbumiTTSah0aRO3ZPIoY3mXA4l5GhQzc0
afARuY6PIKF5AtQrj2TOtK8DiRIEkUFsZAyVJ0biHcX23EbJs21GREzP1/qYwA+i
o3Fm+/tGNru/jjYi4+B3kWQiwhC2ab08AJt4eMlkApsOA1QqItKjHXT/qdmQNwAD
NF5lBjhUablKPXKDbJiYlHRb0jNoI6OvZ65WMNpKO+ZMHG4stq4b7b/h/Eu0fSsP
JtlgGYAt6ft1GEK3Fej+TMkGwNqmPFvoc+QQhJwi7ayUcFyR/UMtG8rRaEpM4yqE
pG0/oO4XXNexQYuoUnVnWLkkUfR7eQn04GWBj66E48+vdXsPYyXxLuxt4LvfJX/2
wDw7pGrB9mloo+Xf7jBwdJpZdg8KRA6JPknqVaCdoewhEbn0DdKMHYJtnkhKVLdD
HVRLOElurFfnDkOnBP89AOCPDmAAZ8CdcsaGzxgHs9AVVIPpxpG3DGlop7S+pCTT
1yCv7lVWW6MI9JKdNZjag2Vp5O1Ggg/Fyx1FcYTzJg3R6jOiLZt3/M37ohcU6lCJ
F8zLxcB/lVJXNKOgb2tpZXW3OBWISMb/gJ/ikhTw7IurHnp+pA6pTfjESSuEdKBX
umD+mXnXii31hl/tTAAavfUEhFa45XanFCSHyfNqQ47xCoUjXlGnF2wCmzwc+JUv
voUhmCqRFWIQmcXk4zXLuzY+PKlF+uagbWVDz4TTJI637JPjon7kDgJpzd2OJVuG
AIsjS5obp0R/RFxRXpkP0LlH9gKZKTIOwkNwiw77nROuRaX5gAisO6aBwuY2/2WL
WxEBtDhuG5W+80qetQaQGA+sJBhhEIB5FSpXckgpz+hnsqQglt7XSwUUwZZwmOdM
mpzBw9RF8doI/LLUsHiFhTQ4iliA3wFzzGB9OIimz4GzXX8a/kuxlk+tR39LZMYe
0WmMQuOWiUHCuyJDaxPIZ/OQJiAq9EjVUkpyURmynnD7kTLPCByNSLKxbUyn/6Dq
XCPsHG2wY+ny3AQo7nqXzu1dvqjh+TpzTCbuAIWzxLiySK61XFhKxjL/I4y49/1V
fxHBtUjAmQG7e+vf18aFsi/V+5Y3X9KqLyjk4n7A8oJ74zQUySRJUZ/4yDquQwpj
XWIiHtInF2GQU17VPlh391fNIMF5IJcpIuXOcFPHjndCPWQxfDK6dOwqeNgH6sP5
9EukA+5p7EYr7FSxh5iURfDTilRzKX77VObe2aMzdSKCKvrhCUTAA6ShllBC6p5e
FBot/FXfkqX537GSge79ecZEZLm/QZsLsI3Qld0c/A9nG+lawlaT8sgx4MbGXQ8b
kDAj+3gzlMqQd0A2WXfPSaf4U8t3QgDWi+IJQKIdc60dkaEI8c1KFrlvMm1PmKw1
vyU6HqsbnFAdwtikqRwB07KjokweAWX0ky7aa9gu7FCMtBGnBlxY19HPxy4i3V/0
9RqVY4BTVnYUah/XKCwFj1Ap9yYXgAhrr9jD+w2VW23kLFfvdCSz2kRpv8BpEFTx
gM72q802rnvrRPWlvkqoMJBGGauGnXwEzrdKre0BMVs3EK++5UofoyGK6UbUVeSR
F/viqCSG6cYLERsnV6RI2aWRGQFzY5TN6K6mXmmfMwv/zFelg21wZ+ksI8ZjoTX8
Do8Phh7Lg5ii+Q8CXNJo4YAZT/HfBI3uH4fdPEVZxrL+6oI7Hl3H/4IqhtjrPNum
eJJaetsRlrQPENT+6gwOfE6910EYIw793Q05p9uLmfJsaraX+fsjgtUZuqHnvI9v
9EN6AOdab+YizrZMFfF7di1wyWL0cuHCcS2LBj4eUqcUovVTy2oo843N1TdGJTNS
e2JVmxtqZE+WYZcXq3fpIwK9QKe3OdhK72oFfcaUfVPk3BakdF3/4fPonuSQVs1E
AU55EokalblpgSaQ2plYQEE8uepEnvfJwSejkp7yHrkT8lOHutZAcR+6Wlxe2Avx
nbrwaz4NnJ1NgcHv2tegq5CenH7/FhRukrMizIKS+H3ltsDotjZfoyFj7Ve94L+d
uvyA0qJZX303qKIlkFKgqjocWPfPZIq2kNzWm/CDu4aMIa9bTcJxo/S6kjiAwnJg
xzT4XUz35AbKobvlsgT3cQMMEggdKCU4yal81dLUEHbusm7q7MmKjDn/Sj8VeUnX
QQ0TYeNV9vJWidP9Z1yjIbNjPx18/2z7Qqut4DYuGKK4sMC9x9QxSrjjz5K3PiDF
yUu0WjTXOvWAsDARKpC1R7sGljBO/JvypHl4ZfKJsLTYhOSd1/dIc2vXR5NFbGsj
YciSR9PQrVUNfPuThsUad4OqT4jKifXc4sRyw8FCfE/T/nnqkjej1uu6/UzX1kvv
sU/hlp/ablkis43lJ1/wi0ACUBqXFc619jOQbmJfhqVpCLRFkmX1xc+OodO9o5K6
FAgxN4dCwojL/Meo7QXpdQKWg6Ho1aqX9qWpFbBOI9DO7OkzfBwXfNfbvp8LnB+/
0pyeWgPOuML7042Ajn/NlBgsGr1pZxt58YbRH0JHU4iBPzeyjYVS0nHt4JK9QJeA
BkbDSIunU3kuJlcAB2nh5XKAaF8x9lpulevw0/6U9hlLDWi2tZorhHgiEPI7YAWy
kCsvsZPKEdaYUWavhQaIn+a3pfjwPQXdgEl2FI+XPLcLmU3jpCI0Bo7wQjAFVLaK
icQfALQZWMg7N0kGbPcEO7OkqRJW6GRyf5Wt7P85mkXXIgvP3JPqV6HzqboCx7Oa
je1NrWup8hRZpdfFRsO1TCmfNSZ7VnZEq5khc581DqyRPiok8nFO02GRhTBjGJcY
oFuhgTN/b+WUlTSBqG/oNWc8/yDDXRdveq9taWLu6trc/NSG1R+mC98rinKbShub
VlfgdTHpuYeRf4vN8YkgoEB1CUGa1jsfKPT+DVdE8ta0TsAcsQD23xfWlPGnb5cQ
sz038zyZvKnMaEwac3TQKnTkWb5Bv1orb6rlNcPPB1rq4/6WvL5O5hzFDUFt8sV/
z2zURIi3FrjZ0guGxab/DwXuufRHxZ8nrecrY1h9cBi20s42ebBALoiGsOZtsA1z
UxiJxvSaaKWQwCyFHkpGgEtR2i2HFqBgYW/Is5J5eWdYpDPO7b+Aa6FihncaYFDc
Q8+9tWvp3BQH5f+Akn48shvSlSnZRkScEsw5o+IlCCS9qWmITVUfF5vFPuLXdDkt
Zlj/0BkcDkvPMvhC0qLQ1tPd8GxSMrpw8YLrM2EWnOM+5tGElJdGz06RJYtZNUPS
J06YMaD2CZPFEQ48zqu5zQlWYbWEJtmoKEuu+KOJQc6JDbnjwUPh64RLFjQ3WE7b
93q7D/HQA/ViI8bY/SWI99VpcsJLkFmPVPHIEjzw5BRyLTNqh1QlIK3w8fxYisin
0HllY16ZCWKkbVPStWqg+zyVFWWUYSxpIYPXCHF1JPSuNYAo+dqVT0ILU0Lm+JMY
oL3diA4LkuwaLjhcw28aCVp9fr2sH5TvItrRr9M+CB6ZTWMAugLkgYQGxmPZBzUf
soETARWblymAD9gcEC8/Pl+S0T1AI3Xnt5U63OrYnOxz63LtUToVqFdJ6JL+ft+c
u47p4MfX4NcqDeT7768cQ5v65GLveMunGwVbRJ8g2B57TNEfa0WVzL6loESvxDv2
yLSZoS+F1LtIjk851+9Teb1JQMTsTHZwYp7DUvTpUcK5lyYfzb87SaCoaODrPepw
s+Z/c+As1ZlGYtuImON+sczHhXTaoavajyMJlxd/tBQpzzKKor51pQjIC5Zoe5D8
XL3PK8zKgGZZtaA+GYm8++d8Nda8qU2W2wYPTSpgHQmWAP/eijN2swRGDQl9pQuI
oeqoRFAJYEWFh23FDpNC5/IhF3cWNko5mBz0BL98u+E94aVMomBdBgmJlmNXnRQd
FP2PeH1yyhDPkTzayQ/bMc6O9+0zd/9GgvofgrDOjcsypp32wdixKfTJYT6pg4b7
2pjyvR5hZBiKl8KFqbNtKBMKCeTNIyalqcxCDL/Wu/ByZG8UKaaPahNICY/ZfqDD
nKAq70WDjX9ufTD4aGqH35Y8/Oodx7+/pZcpPC6zr0l+4hFfBS/iKLopZfFDWqZ4
6nAtQp3EtQNwAZXOiC1ylfxlT7iwSP4MCU4ZMV+4mbVeYZmzwfOsc1plZdEnAdwg
j+uL2Gil/c6PPGkdwOjY10B2Z6Wdx8zZDFmCLZl6Ohwj4Kpwp3uh2/n74+Piz9Nl
+NHTlDXgXDlN6QU7UkjxSr7TH3Frkx2+hQ+AfXvFzzpI+bOSpP2ePaURpORRjUxd
lPu4PWUOhZgDRpTTQAC4dfjETkTGKhhJKAOZ7LnXz4IKl7WLgDNW1NUa7iwzNMV0
K9utQ9kwZIy60S+gEBMGRaicqGnSp5QK8UggL/4y8CHzr+7JKSlFgusyTVjgjCH4
wc84/1F7um5X2WdkG05vV1Lkvsia800liSJikWOL+Squ0J9S/w0J+ax754e/TpnI
6Yvd/XitJ3MbPLTKA29RNq0HoET28yotRpA5jpacmmbmeUHdVEaTlDTtaWHHYQfU
olmmZjtb+rEpOLntbRaaB5c09QA1IZ2jI3AGB13BN51Lj1JQ7bfYXnHfcx08ZvJe
Q/MWBI5cdQUjI69Hi6N75eN81/wjaHyg7upNLMjH1T3DbtSYLyrDNMq/ENjuTglZ
8oE9LY7c/q+TKqnXvAXcOQKs+DqW1EKCFdp52Afbs0++iD52MAiVLZUPiY+ovlwI
texc4UCvsflZdEYIrPgYNfjNb0TeSuM+aY7l1LglN9MqrRA0IC22ul39WEym8f29
`protect END_PROTECTED
