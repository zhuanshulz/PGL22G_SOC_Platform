`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
la0vqjc8WerGyRtAPiuwrzEK9Zd1qp3SU0rFaub/Haxo1BBoSlCAAfjgSGPtWR9D
vAhLth5DmLucCr6usgogoYNj0Ii7fhDFgTTxe0mYT1y/p+93dpqK0QrcE5wW10p2
/DO5vltxpzsNO3eysesl0h3LFR/wHyc7pBZFeZBxgnHq2cj3go2N2mL8kfBID54s
AuTbwxSFXlnLv3KmQM/ZHjVClja/zUkbxFU1T2SSRaCqhhRIFndx8WXeLc4rdrM8
lzlhoxZgiqZcc9Isdfp0B6R9vZs9JW8/uoBPO/sAjAeUS2SjWS/8SSEzGSpd447h
/rK9A1znZ3rrrKD7tSWxFslTtvKmxvveRe7SgV/w+3DkFyOmOLAJ6+VaBFo7s6Ne
5kusdZbDoE1ukdFnVch1HjoyCAETLp96UmeWirmFbGVFsGrUg32SoC7Z8+fYb7cH
knk6PaMMocC+qhljf2hKnL1CxivPVVEJ3Ym1t03+lnjw4MXhlDypUrZOTZB1cZsP
uCjs14fjDDx1AsaCMcqjvISLEONvUlp98MzYYeLq3pF6Dcut4XvHAixxODdNW+Mu
RcshHqdWXsuOucPY/mVssRF3Jp997uLb/gYIbik9MzvBa2t4VpmJDucac3LED8Lh
Ty2JKxaEJMjmQsnn1uqFP5BcadjOo/xQcRn8x7lNy5asT+IqS+tui0g4pCi7op9V
gnt+meYFVC1w9K5ztYmVSJnsFzUQKOJ33GWdtXHFL6Tt/OBUVuJsw3X/6MzYy0Mn
ipq6MS4rNTS2BOEl9rR/raMnfQyQ/pAULAdTDTXnhXPVtkK67X4k4LTY00AFmI+W
sPdJWD+XQQM5KYC4mgFBZSAyclyHx5Rftv95wZ04ITylHEKwMBJDCH83yVNcE/WO
OgF1j85/uzG2/8TLuOZf/vAkVXUZDqsqa2se+qr770B4EODqKx8c8ATb/xfKqbwu
QXh7V1CYOcMi7Ci4l183hGrK4UAe5xm/+vc4N/Zk92+FKlWGArkqBVq47v3Y2bhX
WT3FJIMkL4PWytVChSGhCnWF1TJtvzMPBxW/cmd4Y4Le0Gadfn1z+3gYb/UHaeTF
B/yNtpY+QZVQZJC+Qe1pyAhDPifthgEnxZRfciY7STRnXMEval0LbkE4Lzi/7/Bd
vyqYqtc0CsAZpEj8pLYruxO4+HyYMMKzqYBWoRzh35lX3K1ifNCDhAlue74LWfiA
EMTJzHB2VS37erBIi0D2OXaOOqANacNixef4dJkwf+rz8eNT79ZkxPUohgM5s4dy
hhLP+QiP0F/iwJPFWVdNiESu+w70j0aAEE8dnVJs81opnK1JWSN9MKBG0fCSPhv2
Juxnvi8wCvpQeWOG+RTzM5HWbpIhy5LaZ+Lkfm3BWJH28VWz7fvyYFVGlEIF0nbb
NjXh4Eqhro/RWGmtAAMA1z37Lcbxv8kNQSO6qz/PpMxNaYAH+TwzJspRbuaaJgcK
4aM2DCSk7LeNmxXHNKG9Jzw7sFe0bgOi1G+PRCGm+V2vAdnSPykXd61ITKYOTrLa
miaNM8ruOqxuW2vt7bPS6XRHCh2hmDC88WKNC85lhbRDD4Y5pVEhKsR2m+E/AlVT
UQu2mZHfDqvHUSBUcmrIxlkdhUeL6WIRaCkOXvHhlbkmFQRBtZjf3483knwfwKxs
mFWkniPXi9UMLr9r1kQoq/HxeEnNA2x82duXCe53uSjxD8Uqrq1jlz3E+BW8NkuP
XOp5+Zm7ErT1wg9sNtnGx/N+thuHEYT60/TNBFfuCnG39b/etxaTWktH4Iw29qhZ
2Oy29U+Cl+ipjGjKfbAzBqlytIuaZ+1ruairdKlqmZidLhCFaedBMoNuNH+My9qQ
A0ogrX4vYBE9+L8+K5vBV9txIpganvOw+YmyZTTaSE1DaDDwMaCw+OGgnWbSJDOs
/qhK+eiRX8RL2owgACJMBw+/3Gmk6YcWibTfM9vuLAQFi15P1k8E1ekVu8nWll+I
luZrtZxfUrS77GBezKhsJdyUaxaSqgsAFcbOYBcGiGLVDycAGYRvbd4nJWcEOi9F
RVs6ZmtvbekR3z0qHcKgHo0TCaz883cgI+pWtaPkMSnmLgm1O2bpq2NyfG1oFYYR
i/K+8umscYDvzSf8zx4r1y/3ACk42f8Gl8OCjgAUq6J5pGeZkrSdJ2QVI0OKSLLa
PvkQmEHj3PWk2haR0iYtcDoUl1SnrvuDH7dYiacaK7qYBK8bMKpi2/7iaUCTcOoN
fCenLJiMURA6Ci8tK2Ghag==
`protect END_PROTECTED
