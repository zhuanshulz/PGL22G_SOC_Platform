`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jemd3QszIWSm7XhL94o/ZgCQmQQ8X0CXazeDpdgubbZTzXSMmwYnLRSOGV9RGh/D
TLTLgkn3o06zujWgGzTPrVIgeyU04UaglmFKLHHFSEgNKBGQto1W/7Qj+412X3k/
9vng24ZbXX1UvBw8/bBBezV5GaBIo+100neuhaGoCC7s7SIhHAX+dxLOw6EOofFG
VW1td5Mij1yUA9T7sykRJ41TNFBolCSJmCj2WaRQb9YehnlT3LT4fXISLMtoLTO/
FxyP1Oz+8nqLd/N4LoK5bM6THI9YCeXPQOmfL8lQFmWfcHvvQXAv6+R/OZliasmB
UerOuxyaA9RTGqZv9zj48Jko4oru7eX8Dnz+o32OXVE2nE9/JmuTaE2rj076nxyk
NMxEapJlhnhc0G8AAXxvqtVfcddHmSedHfs4sobJsrF/pLV5MOKbOmm4TzfecYDK
/bMLEyZZ92E0cNmk4gZFgHhlA0le07L3Cz1XySvIUM5Y+q5QpfDIW538YgPfh9vp
bkfBqBYAIW2OxEZsskSFhA==
`protect END_PROTECTED
