`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vVwLEaYoY3w6RJ1DRi/SZ+sB5nfwryE5kJUc1foC/k0srRzdTzD6dEGsJ6APjmMg
nmMUbZFBsajIYK10lZM3OhYZ4xOaaNcXAH/iHW4Gkmvr1OCeJfNVQ8Qc71e4ehHO
5xvyb4jpp9OcEGxiXZ26o96kYa12a21t8x4HAiFK1L61AvB/yWwKwXIe8NhW+U4C
gnT4rUxVj7JlGnt/hpNuZ1dNORmMRMBNFGGMSR+0J28UnUYL25q8QerMO1UGiTdo
2WpnUPnaJhxNH4zwk8hO1bE8RrJXPAkAiwGCIs2ufXs07/ApvgGWwulwTb4s+Lwu
rvPyUFLQG7l9cgHk7xeV3oxjIF/y9n9hQ0V8FbtGUA37gjZx9Ru/bKt7OorhplLI
OCUsB8VMkgWlkS3XJ6GyFTPh9L51oov3vhti8XexHdISgy4huoOKd/vbCqHTApyu
IqSoZZhBNijl4jvISiBSKBLwY0V9VQwQik3PEX1XEokFiL77whC7plFQkG+GxyST
RqNO/0gNBXEQk/GrowoctmJwfYE8y4HZBbHpu24ogWsZ5YFTqN+vLSkwmHt3Co0r
P9z1H0u8+rJ1rabFx7DiutCha9HTkz0O7/Rx/e3WfZUP1JGBvMB+OwkBBrMZndzD
giNkpPZ9Kj392IvHwW7Y7D7LxAt2dxNb5qxI9ux9Bqfqld5jsZ3vCIg0ZlJxX8BH
MiP4vryflgvCGD74pqF08nrQod+JUkpeZdXdM3d8R3xk+nf0AWRdNsVwnGH0AxYi
tdM1Nbyv2YgIGMy78ENaZYKTyg+ygEo7/3ZYSpcOFlvoxs9qlAoiNkun41a64ni3
sy/XPfsiQspCrqLiJbe64Um+YarTyuQkcHi7m2TfrxF9j1KNGaZiteyx1oa2vEn5
gla7mYE4pmEX5LlxgykZGfyhn74dikhwM5ZKb9OwZkwxgwk8KcBXW2h7ds81hDo6
1IzFFF2bARQjO6VTC/BjrUz3ap1b9xe1ZZ2745AYgDuEGgBY4ZKbmUij+hzdXXah
A+cQBFPL6zfipdA2UZhVSv/DkAbTnOH40FzC1Gq//Gs6wG31Sg8dZ5/Mk7KrBcAR
keZRZE78x5G5nR5ssWikE+X0SMEQgicp4M81PBN0Y25/Ny4RiYEIZlsAsWd6bSCJ
+nzAoozCvW5fIK+1aaMaA1uqWa0L+k89wpX7jQVxxD1hUX+VdBkqIJle/GsnulKT
wtUfbKVGdblYiGTKJrFcOMIhQ5cILdMWZ9JJeMAR2rEy6XEjJ55UdFS7y2Lz6GxV
0/7Ft00K3/DEdOOxzYpgX72+jBPevGg6mveZMKyWI89ZA/N3gFbmJPSSkiRDzg4t
u6PRfIM+34tF7H62mjKsIH7Gx1OQNoHiKlJqOYe3G2w9TKyuWKuCGoT7iR0RCnE1
doDFmlXE5lucwQOxncpX2QrU3UaiKXvkSAR10st2TJiaCEID3bl0MDJWHNrQ4+q+
hk03s88AzLxvjk5mYsfWc68QLKn0d16PGt7IAc1nJ3sW/JqVzgcL2OFwEXhlHU8d
azU1Fi6s9TBkjngkVH9wIEz15HvDMWmzGf1lLcqQw6SNrNvvrxv+2N7WfWNjXL+G
4corEJntR2O75LhmtGP0PXayvrZOjAuwQP1GOcd/3ywfN96wCJdMNhbSYcGCUxll
qnG64meK8w4PQ7xOCIrhtcx2VVEIQO1Dv0dyHIuNHsfDYs3Gl7C/8XSl6jojBOpM
P4wsRu+3p+rXeU/FnV+txyuwG4ApONQp9KT1GXoj/gA4iFYQaXBXKxNpvmuZcjC/
jCd1ATORxYsD9bzOOMb1X0YlMZ5pBGG3ByFTwv1koj/RTMPGbl+8/IYEGonug8oq
Xkr6720gJ8bxPQFhXWxYybTu2naMJ3FYeZOMMeSvzmjQN5sC3pSFzlPyMXK6MQ6m
LAypSP3zUG1TrWLI42DaFF2WAzI9ozDl1z1YsXv5ADLfejbe9sk5fa5kY/3fO4Gl
gstJwqCyMxPZXD9gZlTvXMCIoylfc+BY5TY9pEv46dr0mhrwk2PZxSgt6+XDySrr
0k8zS5YID2aMd5Emen6jKj37nHlpVo5gWwKlu66FkFJeWTOKMXAmpNlsvHcbPHwP
1KSrp30H6r9Lr5GL1C6Re5alg/mtcgxkqwijPiODPLwdZTGccIuNnGhhymczOJjf
66hvBFx8+rUELAiJv8POIsPbPl1vFm2Wrzb1EI+HYCI4T9DmxGbWXyj6i/oxJsL9
bPQsaLokRQBrTQpOUdAxjZyJu8FdOMZzt2mGbhUTrhaSj60Tqyn13kNH3vgv47t4
EQswy59eLydso4HvRsYF7ZWdRO3EKN3RX3SZ1OBHC926enjqeaiJe31slxazfqj8
3OKH1PD1nMtERjoNSypDGdQj2MH9dpe/pBurGmizXuW9GU3QoSjzwYQZgevr6+7Q
OIF/1GqNq7ZJ6v3OwjkEjnWLUc8n8tddM1Qu4WotIMiOb79m08xB8lY/XqRREJox
fvxS2QfvmIXa39YdVoAf5nZWUGaxSuAeWLUqHq5ulVNkE23s4w12wYaNK+WFeTNg
kEwNeIzlCCJxZFtq3EzgDnL+HnK7jj3mFxVtd5twvSFaDJMOqdHJkkUF2PaNRdFo
FwwMcPhtjnuxqMu2NnTvdZMi3XFF+9lJ/pzL5k9zJAALksE5TAt/i73dznO7GT33
NQc7PkGCItFV9iY7mdYfBUGCqrNAl9GWg4LwlNszqAMu00+rENwiBzqPRZB8RSuE
L9GkEy5PNvENWSwop5313P4+CJ/lLdQgrC7u6D8Rbgth0JaF6jQpnk/iPe5+Hln5
GkEr6Hxtvd+20/oyTUamtPn/YVYJ5gy04RFag13PRfWUlry1l11B/JBJw96/DauT
3mVSEe8AVDk18LT7Ez2NDTQKsfG80qJEQkQBKcYr1F7/+b1VtgxIOFtFhTjtGxkD
0pcRBLPWYIfujl0+MCtk6F8+CnaTHR5lrSAKL6p+ul8/KOqGn/a12SuFZAL8cqPM
381FG00r6WkFDQNV0N+NffM8i9kJvO3xlOmV1p+4OuDRwNVU8yYRSe23pjDK86WP
Ai6chk9SCNkdWjr9dIrr44FgxQ6qhEY4pvLWZJvdRjEFRAF0jcYRtSsq0YAAEZ7N
QsiwN+LTLFiC3kukEP7NRorKYrpRJrRhkEnMxQsTfOxiL/sbn6IdzvqNnWiE/qNT
PlVjqF0Ooq7KJtBM4SgyQTo5Vj9xD7bn630IRXaazQ07dChw0NFJgPZpJx6dpmqH
2dUQaiAvsUVPkyNZEZahmTr4u3e8aND5v7+wPdmVuTGtigGcb2BEV8NU1rcZYIb3
s2sh2Iwg4m8eyVF+VSiMYJgf2XtqAItkwooUFDr0gR9s2DLRJFvjlk8O6PHZMfE0
48MLL/wGKIXJCE3Xtz6hR98ra7AIAFW9OdvcyBgmEBcZFhZ25FArOi65T9ZaNwDn
vBtrNwCQ5nJW98ASqzUnpVLQlhDICsAFc6ZwyClTTj3WePyGWpMuFWw+lsHkAVVn
vhOvwha147cHpIkhz46VxHoww1T2pGArNf0L7Z5mog3FlD6bMp3aZecnQ9GjRWOT
01cjPiyninotdOlrRNz0oircsD3xuASUvup1VQvAHtWuFToHR0N95UZ50+FUo6OP
Gf5fTvcFTOiHK3zSt8H9si2/8AoU7o4xw/yt7ScpyPW4fkmMYeLn3toOyDgyeStF
QHMnCTKAemlRpvEWJc1GlaD9kTjHWTsb7M+DsYDKtIqH9r+j7A8+5a/N9fZaqG1B
UHI9F4J2VYfiJBwgVMEK0GgzuhPWJjrzVNTx/jlg2c9umCsSYVG8R9iEu5wc+VFo
EPWSeiuryXWB0uUo/0y9NJ+NQvyX9o0fHifdAAPNQiBuTkP4qWCfemuaHeEwnAUr
gffnch6Jyt0xWb/fYMwAbNn83p/JK6ieKu3D2wbrMfTxDBxtIWjcVVnFDaG/OAem
VrbmQKVHbpgR/+h2cnbcGsclxmjcq8Q2k2hrkaC1uMwXosB59TK43RFpb2wb3iit
Hcf9/ygxVDD2uZboZcb6MXDYi8wipcNrcPEquG2lvu8C/iSyUuFgH3hjXS9m1nUQ
yI7gaoz2KahpWrlCnDbtnhBYrOW93nVY3Zj0d2kSlxnQyOEMq8SYsjJvx6krjlt+
kQsOrkF19qCaxlEC89cIN03/rZ2hNbT6tC5gDv67ehpdjTBPlxb4LyEzAfR3Q64g
5xfQgYkzaXutXaSa/VjzIvINTRFOPbIkJEPgUVlPE9vyffCCRjjiy1SJJTp+kn+m
q+JHDjZxB3TVI0gFWlOgpPcXbBT7eAuauxijtJi2g3dhQiKJZB7O/m/Fq5PVkPyV
6BxSz+gmAKWuHm+Tg5Bq5G0GpTu8RDBm0F5/T+dAgROyzD/Awwj2+MCvnvD0Jb3X
dgGpHZFd4IqlipPFfX6i2DY4kQTtrGYM4xOyfk1qsfuwM6cK+cDeT6NN0he3bx7z
RenFqbbJm0jkOKPdOBaY7r/HlV1lKJHnrxrgaJDYkseEIhqsFjk/4EZSA3Cpik7s
N5/vlBxEu8NhaKjDOTuvDCgqZk0U4Otj4qg/Bw+x6+1+S2/B7sM2knxPJe1AEfc0
OEY9ZeBfx7Wri7kTkQPACCs6phSMQQeGGZ7y+fkoYDQ/z4nKIXzgCbZodwlJhqgl
qr0gFTxnqRVjp9Cju/nAdmzcmURVIyaffb5uwrwZiB7013Gfr7H/fOmZXP+amFhM
hCEaoPjLLy8BgE7spQnZLy+Hvvr1DSWeCjMNDsL7k37+5CChIjBffUtDN5wRNDY9
V4dXfrCDCCuAKmZgt4RXvgFmFy5WxX8phy6mH3xCa+EbzwcIwCNCnTQlX1qdoYXA
m/VpLyrkVROOq8+8WpNkPyEGuPjXTFRSZwLKKaF16GmXwX5XdfDLxOVvbRiKv1aA
NO+uzvgaBcJ3DOeczO+o0XtWOGOundMvCBZWI7oPspj9ch2tgKtvG28/OfkgWOmt
idpdKlu4l36fsPeV2tE3T7A9rVpr3buLegyUMNRaS955Zps6fEFk5s2cdmDbaRAC
84J8H1T+A6gWwQeiFZncOXdIdvBzRTXZZhT/H42pFk+tj4IwkcK/yKD+89/YOrPp
+ZRH/rj2bOmGZ/eX6LxBeODNbXcelY9jXg7LWDj85iT932jMnhcJei/6n6Y768wQ
4T+rKF1XUhPYHYAR5Yiz5jxb9hBrQiHbZSbT2LNv79thb3618CigAWw4r55dz4Sm
KM7eMeetQmS5MvemgtrdNciZ0jXE5E+xIPmASU8T8eu3uCme4vxNnY4V4M7NrZs3
VJUtIL5OAO3EGAX7e3DN992Y7wRHA0JuwOVpEdEK56bli9uT5LziIGKoptndYi9F
wSEGqa47NL/a/I5W+fvhK+aafNi6RNTdId09I4MXcrz2nDBLCgbdJI1qdtH6NkHU
JkcVEYQoC6sFacq+HSLazVGJlH5hWTJx/EmrAVTi7cOPzUCWHZ60u6VIt6hzRzXE
pjmSLz2fLoLUksmdLQWZ48aoNCSfpqMjpMik7pPuH4kRLqh1MbotttjsamMVK7sL
B0HzZw//yWxULHyf3ZnUurItnGHGF752ZNLeCFocQKshIZzf/lLIYEhXCtNhyArd
uY1NYAUBGvO9kZaYEBvBnGOgPC4ou9J3HSTeFIhxGqENtk2mCqqp8kodduDU343O
1/BXnhsr4EcDhAcHH4kxXMUJGo4SBG1pJKxdbD3sAXpcbDi8mTPmh29lt9JQ+AGZ
K6STuAZgmD0a0zm/RSBKsS5aBKMMfTxUs8Bhsk9ypMcsFAibczyx9Pbm+H6br4Zs
TH7vZYdu3fwaKhPDPT1Z9tTqT7L7XeazYCb6nNtZeLirNew/9gncpyMHcmU4j0pT
g/yMkryLbQELObr2Bb316Ede2Tf7vX5rVWMlvGFII+KgXa0azx48MNLHtE+L8QsZ
Emd7Za0mlXBb3IzUGv0PwQ/S0aYBeEVIEoui5eSoX4hIqbDbljQijGjKzxIAi0LI
8gIudCtW5foz6E2cpEhAw+kUECNezNYJvoRFl7ndZoZYHzA43zFt0/UH+yS5JCqN
F9aaeSxE3EFy/Sh6vmltTz5u0ATAWORILbvlK9mKGNHWsBLtXv63KgwC8I8eA0g+
HK065eZWyqPm3rDfViZPheySA1IJqM5wXugxQjI8LTtpsKItqgP8e0Uo/2G0zEFc
yVkhlun3YLoia9suu4j/WZdm+TaUInNxCkWB05U20Z0WCQtE5JgJX12A/hQO0cCR
rfw6haQs9uYr3xI5IdCAcJC4fhhE1eoKXXImOOLQoSLex2jfCN4eWRzdF+0jbamO
RafZ5NSQGfNnIo2v1mP0R2CoYVZAg4qKy96Mhr6ytHcASJRH9WiZGDua7j39k0zy
iNaILH4qWiInB9K+YEaYbi/0MnmS0hoIeCK7INY+XStPsGQVoP00NGUe/DiQ0R49
He2grLYcfxUqwoaAMbSEbIuxoA2ER2Mu6TA10GOxt7TrvQN+enIsL6an3SYybdzI
bJGdBohawn5ZCDNXc4pYJ0Vqhy9m2bmxi3r8toaLedm9kgmCzZ68Cyscr/91lneP
H0Q+IaFCPTsQeRsMw10vNgvPk7BO/F0AW6uA7jgetwQQS9nFXI6018K/IrDWj0pL
qEGEHrl1VTqrhrw1xa77M7VyYkYSIpLBt1slBkxS/VRukAynoL6Gb7OYi9YLZsjs
tRBvzkzL/QA7XlLxKSJ4OZ3P8o7FmZpl8g0iKpK88eUVilg8DKaVhqGw7fQTmcku
VhOhKCz7yBBIqbXPSsNcGppb0vEhIjhD4YnOOPkk88q9Mxa7dKlFkhPuMvBwRZMK
AEmomnVAe0ocWFKMOsPPebJFr5/X87GVczctlQZkVap5qsGqNyaQBeAyO7Qe2AjK
kHAyh1NaY6GoWH2T6RpkiGxy1DGompagyANrTd+ADAMYkUPdmtR69YXAMPdxl63w
jCF87vQzpkJWG1KBcnteNxT0gXuxsDTaPUfhxH2dI/WR6er555il7EZiMyyy/k+S
2QAHurSXYB3wScsW6Bok4we3cYY6TMMqp82GX7ZhGV8bmoobK4Ah6pFIf1NHBaRq
03+/Hybp6rtCfXPX4F3HU7f3wUCz73P6Zm01ItW26ACagjbzdSod8XCOM4z6cfdY
va7jWWFaYFroGsNBmFveQwLRiAzNLPKisXtM/7Fzpqs3g2FOYnjinMFvE4exlHIW
3OqudQKPx2ury6fYE7IPctyQPlwQtIMjzvcJdru8PJMg3cvgwdKzBXwH5LaKfqBr
oyltWpuKqWWSeRDZbh/JaMcNxF+GlsEImWcLeGusHw5mLljdEiCPLCv/x1ALB+Js
LfpxOK//tksJ5/7F6NCMRhp7YN8J1MIP6MWQgwok86APNLP4nWoUDl/AF20FKkyo
D5G+P/mtQcjWjZjYWJKytW5OH2HioNiHP3d7zVlIc/TC+7Psf4jetz8a/qBpL7QZ
K5Lz343OYcM3MCohQYGn5j7USsBIE6e9KWqjzBVWZT9eqUJhQtdfPMskJDjAjdXg
7mEJGmMcUkD0/dM4gYrNFEKktXpgthmEtxjaYr6DDb91Rywp58ovvDR16JP1VzwB
zw+8VigXbJQc8bfU7FwrVjt+btMIlgo4c3raf4H1WW0sbikSTuLTxZT5oLy0e8+O
gTiixrDQg+wX1Y2qXveNZ3HC9aOyH7+IbS6xIJV38I7VkPWUFDYkIEfLbt/90Xqc
LVMoQ0EEDfL92zY8wHevYiRU5FQ+uDPdL5Jp4+rSKSHv2NYm5FQer9CXFV5GGrPK
WMn2kpC2VSGoxIa0TOwEHiyuWHSBv8jcWmLzM+N2fhQ6ACGLr8lVlVfz0ERMbTO9
hXp8/Cf4kICNvaSgr+XlSv6mBAZgnKoI5FDJZEvFOLwSNpnHSw9AlNABbSgfRJkf
dKg31A9y79ElBGzzNpToYTGrSKYLMgmPC1E2sNpOYxOUQ/DBHDZYDhGGHoiJAKgj
xbpuVp5UYT3IS6kGTSIfu76jsI+JgM1aLmvNkV7tqRiSA5E1Rogxk71iB1BaYmCt
2zUVJGG/D4xdlpnojkEjU9ygRa3PTT2NysW9DckV8neplIMO6oyLUPHjZ+9372no
olw02RLqWuTd7GdVlaCtIPf+f5UXTKtRoMz16usa/k1uP8VeVCFI8qT3nccJkIv0
tLuzr5or3OPOpO7RiZsNauERDQa8lJql5LKh5ndSRr7tHXyuVcY/5kYFJdAhnwr/
MfDKqx2ztjlAdMWkxMKz9J6FSwgRCCPqECUZ8Vpq5OtJJ1nznxNRQ/Rf61mbHxPa
TGHT94dzkXMJ3qhekKFj3Btal+UF0K422mi5OfIlgcB3cDR2Kn54/+nrx6K3fcsI
UB5YW114Lh9+cFdAz4R8+5AODf1v20vLDyBnyPMYcfZFEnVJBL6ZTCgdbBNPy5kO
OOBTvWhr96l6w4Sk4el43Whbih+3bW40ZkeWxAxFslzVX/ufzU4mKI5h2zjSxXRi
RIIqT8HbSn02mjEQMMqFVza1Q47WRt/1cyHRYw3A+V7orc1G5Buz6TvgiBPcVyGx
XZKczr4lwxenl1jkJiRJWkjd/AmvHVZvAUjIq0mZX1fIPOZla0UvxKpJCTDPPTyD
FAyF/8jQFrKyT0eK62Z7cGJY7MA8qnfdq4eg3nTMeD9s4CclNHJg6F4Sl9FSZjT4
0uxR0Z7AD5QZBDe/S0IZcU70yjnvnBS9lAueR+QKOYL7F/cC9uGnpe2n7+e0Hnx3
QK+OUxdC8DCyODijGQ3vrphbbrhxfbj9gVpb8nbRMsR9NbRs2SIPnz3tQ6LDrCDT
ts41nTuSBen19qJ7oCDgLNjyz9nhy7GbjF8WbBXXbhGDsbtDrXkMjxcsqwqxYBcX
hOVG3aQ0AzvF+zKE9HclFbF3iZ2gykSlcAkMmklpEpHGnpFu/kNCi2BI9elebSto
wodS6NGP5Uv0JhIZBgtkWW+OKSACMb6gyESLetmERv1l97a/bK1IOLC64mghFvL4
zIDiXGV4tZIerKBkWZcXnoFbPXgZnfCA5MO99t0a+icttOxsoTIbY5cfsWfRFi2/
Df/pmhGpzr4U0NqoG0ljclO2FBroSUG1xkkmkAoYbMR4kB8TMPd0Jr4MZQj14+g+
PpmIXgHVMR0CmuaBTeOuFWryU3NOLdp02t3omVNpDFyitEkgiVYEzsXDJbEcw6Z7
KodoAXUlwOUFaqspsg56PKjhcMYnr0aH7D4FL5O9BAvr0CkanxMCqO754liAPlWH
tQhfYScB8fDIjTYicnHCVxqPMru7qlEzjH76FQLCBIBTrh4D0eBPSmPOBd9j42Rs
ik0EFRnfvqKBMZKX4SSsBEnkRCFHg6gBoegldPOhSFtOVh8/HLqASQo/uAkXIEdx
WZb5qBs0bDDWnP8CidhqAAiEwxkQDgE+SePoA6uAXKJHnelU0ParuymMoeoY++/7
fHRn8BYCXdezKfZeZZDAOejezkHgGFKLs3Wb2zeCVeu/wzbcsDfANNxvwff95HEn
LveVvwSkmV/cnH0KXrr7IlofrgziQa9WrxzMizuHkg4SE5LbwOGG2/l+8x7oHRgk
f7XKe0T8RF3n6dGepUrEfiLHxXRJTV3+Q9VYV51ki7KLr6V073zho3vSJ1ZjciAl
m1VeXEWYSRmKovnI3cW1aWs141K+bI7Zh/7fqoylYxS3413cOhF+0LRseOX+/H71
pfhcSg8aRbb6pGtO4CNeRne3I8OFMn6ts9t5pRB7Mm0OtOsQxX0GbKD63SNu7ryb
R2NzpbTI3cQ5V4DE+s1bj8gDb88cDAevhYK6/OrFiou3fdT5zfXja6+E8hp+ceg/
SooKA5rYbri0lF5HZOx4Ppw0N+4hG74FA6Okx5KUij0ELGrWWj1DJswYQmAlBrso
+ODTCXXz3xc+4LtevbR3j5h2wiIbHzLGVwfT6EyErmAcCXoBSUFFEh95oZn2e9Ht
8RFB+Ecu0RfrFx3SLzR0AM9nsczlzL2K4r+la2s6wamOCI3opoLrNyGGcnX3PnHI
yVQOEAPVXswQpMsZgYbefWKZoZBn6cVh3Iw0xjEzxeUwAsOlXcvP4onlo7DMk/Nk
n+NWuhyueJCjSHsgYvNbSpUktXpe8+Nv40c4HPjp9DbywIGH0nCQvxbUF8LEvr/T
XYUWXd3dMWN7ULgxtiduTD0C1CwiY0D/gU0tY5rSL2spFeZaM1sM9N5MQ/dpJUOc
PPa04FQVLWVhPVuwIza3NTEAnxZTg8oY77QEqnX5psA59cMOZc0AodmjKmsK7KZz
K/P7GgviGW+Yn9jo3KzyFYZ/ZGaythjFP818go0a/Oh6T45p+6y8SnqTllJEbi+5
7caHZyhMuy0m4pYLkwm1AK6iqdETm1yfNBEQ/SkMif4Tj2nYJ1ftM8cfcd00adsO
Ko5DOIBwrtiJ1I4l7ZOd+OO1CAQULTqCxMRGoKRvKfrJ4MjYvkiyhowWpkcpxHpG
kvwE80oPm4RGcCRicH/PJ0mD0pfqtBa5U0b1u7ny3/xAmtFUT/cdDzQHJ4677iI9
o839dOZ7MBA65JpYM5B2RVldQ8S+uJp0WbZLH2XgBYwSQiuB5VizEp3RFnzRhr3J
2RsIhvOoeJSI4myZOaHeif5Dp9Vxbug84gaSOiBuZpSwWjoxQz/vfsk+VJrKxlrt
R6b7M+hzCP8J8QGR8iY95oxWp31p3WhmVDGofbpvN1Mrwm2Segqw4JqNwRpwYqZN
woGdKbWLgMJnRjTrQCii4JgxkCADaX1SE+QSvcJ+m8rcyhkfUQ6G0HPkFzdNirOE
vQdQmXQvEM2OBa4NbrW9PtLr60AcZO/XqZE7Qp1cEyc5Yn6U/c/ApbibT6JbOIRC
ENvbsQkOTgm6KRbUfJaR0/0O0IRo0BE+w6eVCFrE+S2KTB7IiYxkXilNSf/8vhsi
ESZgN6ljeg5sucP/RYtJr9ruPSXu/b9UFiO+Gke8z6ZNJq0d1B66Rrt2LGTjRdbm
G2SKSYmCv/5txczBwVdb1kP63R32xfL4N6FnO3g+swxvVf4iV/Q+pHkmjXk5rA2u
rVAoICl73h59TN0xlGyXyJQrzD4rE+LAM+3DRuJYhvxuKNty7cefLXPNkzLpVuq4
kmVl6LXfwToPkTU/JFHYPYv2G1B5jwG7eut1uSUs9uGk2MTFSxt91egxLJsh/fmn
XmPnzUJhR9cG0Q0J5ompZgP8Vp0ml8veUE8/w/pADm7bVFVZpfaNmqlaJMNX3fXN
P6gcmn8DsYkviiyP3MjZCkG0sDR4jcFlzyt3LgUGCv59GPJgF/yCIXRg9qIAj5Vf
8c6eY6XvtZPxm0dstc5W1QhVaq+9RQvV3hBbOBDqEpPe4oeTmF/k/USpTcCx1cWo
kOayHYUE/etRX1Jakt2CFc42wbmkPmXwxwc899rjHhBFR6teJj0jZagRLrA0bey8
6X9HDYQ7hGLYEqJoSsr4olIeVUM4UPFhXnOORkgVcTeVczOmQN9p+hk1XM3gT0NW
wZBoeLxoafzgt4nLUYsaWpRxRlJBAywNZK1GO+PmnthzQvg8VOSIuqvPD5S8AcTH
pXOoiymlzQhcz90RvmsNYwgR12Tm3qg0hjCGe9seyAkg51W/5QnP40kq/ZAMZxp0
+6Nn+MXiJdmlA57S1+C6dUYjWXS15ee/xavIAHMfjsRKcmXGaCG8Qb6QqufkVjGS
KzK9pZZwOncW8LwYneIMlG4qAuUZoRt7LIoH3O66v+gYjqcoX46fJyE1JS3fAKtk
BdRfRK+zaPxVZyfGnr8uRUy8T4hdDINfRBJDAUhX4ebENUhvmcaF8D0dFPAKLBPu
lrr1I05RvpmhbyzCr4GWYfbSWleAJywzfFoX3wNUThRw5ElC+5AapYN5cM6TJlrZ
`protect END_PROTECTED
