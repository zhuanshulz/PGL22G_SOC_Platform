`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kfh+zAE9FyWriX8CcujXYOTQEv5kzhWGW7xnOdtd74eEdUTL9FSLKDtvYZJh9b4Z
gpVjH5WU5UiMb0iZdym8005QU2OZfbTwSuewYcF6rDN8ty8FtdAGxE2n4Sj2t3yA
Ev0ugcIX+WfxW5QQn8dy4TOKR3vedrDWF8sBdjDji33r1XKcD2o68lwE6zgt+j0k
qt0Xdo42ahGTgzXrpsj/RKOoWtgxErboJ8yBOT7dbLrZAddHSsnr14QAWPWYx2F3
q73Ca6Flp4E2+vixKhwhxOGW30ZLkhSfcCnt+FHk831tKDPVCrq5ML8mrcKdGMQi
+8280F8rY3iAAYD37LGCCrf+uh+4Hl2EGGP2lzEvEuLOruZG7AdokHNrdFVmWf+2
9K2NblAhvfgU8fF21NRB1M+OTfWVJjwvY3Ruv0SnddzEmv7Vedg73r3jLx68yN8T
rYcC/ne8YXS62eNVGIxghB2gFDEZmxWRPZ6gDdWPHF4hIJWTFLGcE6wpIgaYShv9
H2r8gLTX2uBi57TVcatK2nS5+pZ3DLMXNKsWHuiofjVNaBcoWQD2p8GhuGim7lnG
KtHwoBB0kxO4dUjpItOqVPGybXr7qVwnAA1HwdmdM7KDj5LwM9o7IN9k/FHYWCuG
Hyz8ElTpNuwOcBOovWURU1v0iGVDRZz9jgvNW1EI25jQzl+YY0a6k6FSsYrjIUsf
28oxXkLMZq5gjz+z+6jAB4iVsismr5EJeCDwl2rSgsrm9d9Ta0q00tZKScRLNfyn
X6mt0Uo7L9JwjAIyxqsmm7XDAlYOTT3uWcokPhbvuE/4VV0AUi5gEqKfvaJRC2ya
IOZcMr1qAfx39kIpmEoDzA==
`protect END_PROTECTED
