`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HNQk/XyJxLCiQBNkXtscTEjFwh2An5hpmv8xZY3QPR7VHNfzhLm7aPpxyfzXjhXZ
rZJ/cDp6QZtaYcnLOZvViT+ftsY7pdqwceDUxMcv7kGgcEXBV++ERkuyyK5CXioJ
sIdM5URoeYEUR+8oR4tKe5OaA4A4tARAfykDaGhR4UjLPRqXsR8yDaFYpL5Q6pO9
A269sPWJlF501+8Tfh2Aa1q40h0EJ3LA6kPHZvombJrt2+4MlFCh1cngQ9syizpv
Cc0WWwtMwrVTXtDtnZGnIN75PYtqfiOAHbrF4mMkYSbERvHlO1tmcosdV5A1ZMp4
wljv6yf5XIFTkkxqc5EbdX7FWPAkttJKiYYh7QudVJhZEzy1TTEe1GDJUkyHn/uy
Psb3gl/Z378oyflE8iYIWz57of/FlKCKaDVzSDtxnrXkXos/IyIA/BvMn4q2bchq
P7Eexe4axNkIlS/tJEzlzmOUsqG0GdDQdEwcXPZWelu/HTVEExp+EaBRD6TDnoI7
LqoWRkcPdU+eTzKkMQQ86+TGP5JlbYYZCbDxvHPFf1HPBb278UFcDa+nEZKUx52g
c3k2ziGEwCFX0CAmsfHr/pgp3+6FoLVQ0ElhJV/blbx9bu5HMFV+uL49K1R77IbY
lFTaitpqZvEcolxMd5tNEx6B69P4RfxzP1CkVSG0D4cgZ4weUHIQSvYV1+QRe/F0
SahVAPhuD0Icjn7zb/f/wQpOJEUqwH+TsXT/Cv4q4CtQdWaylPN0V7qS12eSn7kH
+ifPm6/0W0FeVnBsxpZmmq25M+EgV27smmbELQ5F5ZvnLNa/C5U4EGbxPPX+tmtQ
oUqDQKsaxIMIwxN/9HwUryftPfQv+gEprIIcOImghW4=
`protect END_PROTECTED
