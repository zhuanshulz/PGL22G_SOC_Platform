`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rvRdRNOVhJdQp7oKLnNGw/5wdYZX+et17V2Ot+oWphRDH4IQ52W8IDaYSgQA+JKO
8pzp+6b1EJfRBUdHK6QvyOEeTNXNkzqCYOWWPBzztmiXwcmn29LwFhVFmvGkWzfw
y4xvewRqW4aF1gk4cILzfMpbYH0SmRDYYYiGoNH0UVmhM4foBi6p5XYMjarxhX9l
XVEcx2jsW0cUaW1a32FsJWPpfZNBErwYVXhbxnYouHVv27LWwHGD7XYfOXa5WtAc
/h/DA43VkIk5xpvp4jbRRQhOm1/ilF7+oKnHamDV9vUEeT/7pLLRU/VMbPFSQuR6
dgpNOeryY5LkTGe8zAksG6/D0mwWemE4DIGHtbanEmHKu19ZE4Qsa1BSSCwlZgdi
xr2yYsF8OQPi1WFCluC3Xz6Q6OflBXk4GJLnmRYBAFk0GEzrTzE+en/C12NIFVuE
2FtaOtE9/CdZAbBX0XJNASdpZrqNH5sA5TPbk1w4oRS810ASvLuPc9r2lhFPLPkt
7VDw0AkQFHN9UpjPWldrY7mxeH6oWfV0BgLVcXRDf+c7770GYebKQz+0EtLGJubg
XxD0fGzJz5FCwlXOLVqKVB+iR3G7EvwSaFRDtSyOwaqXjgfDF7wn4XkcnLhRHIEw
LkyGEcC2RedlhAGo+CkiutdI7CYDjNRejWNNzhl3p79sYT6Y4w4kvAwmKhzqei5o
kditHKcLRB2v86XpWbFj1Gr1DOsfb5PEsANULHFCTu9guz3J+5SG/LwhCPQ3AM9Y
gP+mkNa47vAq+G0XA/kU6n09TsO0DTYDaFZIT/T5RTo=
`protect END_PROTECTED
