`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GWfHnHUs53knUepRyv8KYA04sUNyvZgLk70VUDkx/oK6C0J/YGLUwjIFHHMFowbw
F7aK+INMRsCG6kBekPztnk+7LMeJv8ndq+DxuGIySOxokmmpYHZIOuyRTSwSr8li
91jKrQh0kqQOSgV6GRjS5oJmOuyH2HEDiG4k4Fjzsz/FnTj+bKslNTJ5LHpCZpAZ
B3zqY5C4zLTWQo/BudCUL6xbQorTkjW8JeKAkpXyPrUXPFqwQY2WzsHZJcLvXw5l
kLsSQez2Q3clisBKmnf7LnUf8y6ZIxRx0GfP9eBH00mzvb1XE5vKDuBRZQThnMMW
G8oNkcT0St9G0R2M1CNmfWUzqzekmJSmOOh5OPJeETC3YnDhtoTDxXxZsnfVxlv7
+H/LUhF1yZW00jBv1RYoCea1061RFTwxOAQeBnVoqFRogFPfZzOdLhb1KbK/JJqo
XAeFuTvFCaJdoC25HFtljCyVveO2cZr4Pa5w80JBVJlIRNY86GssBjOmfKd4IbN1
2txIGyhgmLm4rpLJ3QgHIYSL2cxnyfTSPrjJrQDqCLdsytACo0f2dPirDEpLk20x
9AoAi1Nb9GrBNhfk0vQGwCyfTt52PaTffB/4trQbjihlboQSnVthwnJR9d/73lFg
BCc6vBwgirMqMVoyeslFEy/HfR0u5yOqxtC5H8ThIZFD9y3+uZvWu2T0qP+wBYdb
DALYUvuwpmMnIAvqFSA15A0o1OzcBXuXIdisaifDDBVII3vW0HgBgDtMktvxvoTG
9pYVnT1aAako6ZlL1forV+iVYTSkwGkYWL2UWkEq45UquWguGEJo4oqK2fK93LVs
ltyIKy2XZETcmLPPmJtuJ0g5ZhXXq9n+QCTEIc2Wfu8ww5pRBW57kDnzvNfsFKb+
VkvAtb9rNo9as9BT1GObk22qVtCbhZHam9V+JhPu/20UZqpc13d1iFRQpQMXrrfg
jvAISGnQU4a9YmnmSoTPdbeEJZtEkpdJWzCCUivaxFZ5+j5Z8I9SATNhlkuDwWhj
F50x8xFVkJU3MCi21cxAS76Zc6nbQPjTlE4snD46IxmaYWaBI6OJ2uNy5JJAqU1o
+JYIcvywMDPIVJMVy7/2ic18VztEydFJxbmGrqO9vFHVaM9Y1Wdi6HPdfoYvbrpZ
vMu4v6uucxMHl3u8NF5TQkHKCotZHTJ9Ud8GdkzVk5+pHdmNMWwiZS+Tuiu3matK
Hgp/ptJ6qM+XMNCRT/1ofzSS04m5atqj27wQKUO3aLUesFHog3HJP7hYY35XJwG0
Hh9cgfuYdYr5b4bVY/8BGOfmkUZwzzt7tS0k77RHspVguP24jmtuU0HifbuP5McT
Hu5kBdx3V5nzgrYA0ubSLp6LGolql8N0buFH3vpQD9P4XCZj2R5TSkfMTqAfdqJx
sqkddFLRliGsO66WM9qSV3BQ+Na1/quIgc0k17obmUHNuhkllKU4LLeHY0AgRyAt
7yVAwePytkLDInLAmoe0ipb88oM/ypCdkx9EhTaM+EfeOyHMhl4T27SHXbekIQPa
hv2S8yqiPuCSe3PanP5PDXgsOoEiTor1Or24gdaFpTBSQkP8Pcf4VeHPrFDzlzmS
9Ort921ulzlIm9xHYhRekiPainjlnMb8DO2/4Ji4c/jrTMKt3uTQK/lWHb1/55SX
ERIcjO+ixo55SezGVw4jj0VCnkZWLd1IXMYKl1W3U0VwIBWZWnvxwomvxBeatWb7
0WwFpZ9DReShyzyQD0gLyhVRxejBc0CJ8oS6nvB1CZFtt6PWX6uJx4hznhEhmDrm
ayP7iAZUqlELorSSaebr5dZJo7H9KKOI8zs/sdHaGa9ZQ1VClHGxjZG2qVYT0pKz
3CAqereuB2uiMYEYBYltH1zAC1d4/apwtRcq0Y2zl7MkVTcwmypJCwqEEYntEqdR
6H/uLGwuMA/qiyGv+UlE2png535Dn55NwEUOQWUVIGJ2ADz85jbM4qltNp25hTPl
IqimDvQbyIdZqfHfDKW0/brCO2NvDAvWov4rCgKqHPJ1iY6cHgR6vG9aYmgfH++2
ZobDdIOermUf7mWybkf9OozBmmGgFaocs6jWv/ghVH9VU6gW0BK9vCMcw2eGuFRV
/xxMH3BxFrAwMZ1qB6tocEpDFeFKe5qsSB7RfVn1Zutm6cZd4GVGRyAx9lCLnzA7
H6Qti7RBOzKLY0/vHAyABwE8z3TDmo9fmaj01l6UYwF+AfGlt/Idi9w+8hy8/oyE
zAuT78KFxzHAWd4vxai+12DHbZ414hfdy6K8ZPP5JNGUwRZlqolUj7k08n9MI1xC
9HxD58LmItCFmF5MGePgi9F8Thg53LpCn7vEFt8syuniuJ3VZ/0rgwHn5owhqrgs
pZ96izBva1DYuUxCk3Z6GKvqfB6pdtFePZTEIwSeurQ1WyoVpQi2JqnbmIOJEL8g
cO+judpTDHf3yaYxZilaewrWCvfNaYs4fpT5T0KmUhCDjRvpHEWiZxTdf7VPnSUt
8YrDMvPZgTSik0UcQrjM8b1ZpLg0fi6v0q36Nsx1tIBRXEDI4uHi5mU0EPMCco57
gZi6knYuXqubeh23dlwLKz35nSThpuG70BYgv2cFUrkJIc4eRdybRp4/StKw9I69
IyDIYLdOP0TvrzftSsfhewgYfI4qzk/H9K+MlFgQLl8eelpnSXJO8rYhLoM2pbES
Qq+1rSKaoCRiMklk3BDq95aCl15ZotdXBij0yZlZ/XMSy+b4chpeyJ6cJZu0K0ev
giTiswgt1xyIwjdadC+wpoZ5tvFDlYOZNdcfOATGtQuIEAqE9m3dXa/M3WpXktza
S0j4BpVATALO93R+z4v1Ds4mhi1ZQqWJDftQsIhRVOZbVCbbV/dVymVaukxuXNU1
mu59x9BRijIXHQW+VlAUeb7u03jbWHGE8I7eOPXtSUdNkKe30v69lsw4bwHwCDXP
31Z+rncqSihARAekWkZtw0cAj1/uN+IrgUTFrjGb4J5K/StnPf+ddEbEwvbtqskK
IP7vjzj10ubiN7h1sDHnZpkMt09X88ljqGn9y0fYOrQqiB0YHWRGZ4AwfB79r9d0
uzpeP6RQO0ltHWAlvwxxbiJfgnMfblS208f583XyXygNAxE5g98eujjznL+3OCjs
rxhH5thtZTyydj0dgDxEXU+pDk/3R3vZ5+A7NrO8RPDKyr4/e5Zve7J9Kdc83BRu
UrSWze3vk9JH+XxBeW3W+1ntt008cJ2/2rh9a9V/fvcBbAj/v3eW+x/4Qpp7V1i4
MtxL7rQu93KdiNTofrtEZiXhg3M+tz6MsDpctuAawQqH37dXV0KvGsU7+ZJBVGWD
MJm8zwpt/93JVKk2bEe/CeqQADQhPVxRn7pKGSesj8hF5THwdxDvECPD21qijuzH
X1eT1X32VEWUCbAVBi7kJHNMGy6rtioae+lQBiqGleuW0xV4uyFO5EueHYbtQg8e
WLXxCN2sZmm/LWUeVW0ZQOvjDxXDyvhuuWrNgu1DIiCBde8Q/uCk4kOkB51vmCBR
mWnL9hS+/SE67dxzaADxgiGID24taQcYRTJhXTP3ana33AP+EoBIAFyJftf0GqpC
RvpPd8l21dJkN5IqUD50IahIZMbFVqmXWSPpqI+03w2ClQn1uc3USkgPjhKFjuZX
SPKkZLIvvEPvCaOLmQdgiKFAOHkKL7yYCu9L+sDuWib2ymC66Q+ffV8ih/QasFoU
2PBnq3imIUZhuocnR5md2ozKru7d/ZkR2lYw2CGEYqJfmJKJXfkEjMCz+7UtD6Jx
weawAYQWHICSNRnIihL5/+RPJrnW0YEPDkffEac4Ck5pCMftAWgIopLhDm18vE61
pw9A2ikN6rB7kUAEQ/wxVoC86U1TpABwmKsZcYYbAKK/z57su9An8/Fj+hhWwyvT
h+TrQ5MuAEzwOrZIIX04gs0vK6iIO1c50f7y8XInse0RAkSnvKtGzPtiHuG+IZTA
7pCAXJkuv3LD8cYYLVuVL+MPgQ/FWgGRIT0cgAfuy94N4wgTF2kB2QwXeXOD53Ou
Db3qt6uiF+JMWssz9L5K2t+rAkoZ4AzgXvSWInwFmuNKEhqLO/z5IW3n5UfvkpIw
bU5Ryx0TWPh/o38q9ux2DNJiT8MPoJtv2GgdeWVWqW4fm4se31AByfeNl6FIHUGE
KLr29cm8UMZvRql5PXHFkaqEpVwijRWzo63WnHqPk4Rvs90MyDIswFKuVI+W6WzZ
LW2aQ1oX+w6VWfQKcHJrtxjgCb55BfLb+fblUhyvvw/jzo6eBdg6vJwMzQK4IFXz
dy58Aui1my7XdbvN+0yAcjf5815gYchs6dBoUnrQwXDJxcMZxBNgCTO0mSFlHWWp
fKNEZIjCzyX5woygmNLPKtrnf5aFE6ByNkWrqG4oYzb1U8HBJfd8YOMDCPNjpL0D
/jGoEi08vEJXRx7pd9BZDwPNNK4EAK/UNcQeOyCRQ3CH3UOLHyYO13slxz606rOB
akQ3Wm/i6J/XEMhVRApcOob6eJ3maxUKB57GI7SNnDeLUx5BKKkorXrmL+wtUs+n
noSdWwpVOMmLFE5xbv/fEftPyEHVezZ+1N1ggfhIRzKsiA3uwWRxdN0rLYO0FWyf
cER3ptfqqLQhoZJrk7YnYxQniOAdWAXZ7/2gvcdoemxL9wmfDXgO9s4GIXkL1Qmd
w3NHC26P43fZgLnf4i0m/qv/qNL7MgrL/EHs/FhxH5eD9koBAQebxIHbtGcxSScI
IBi/U5xvcZK1paORLwkwWQBLNs/O054SsX0sWK1+nGzJwYjSyZ38mvAzAW26y9fp
uDjfL1w6XfNA8TG8/y01X6AGyn5BRTf7j2/Sohp9iqIbpMMg0pOGeKY3H4NQjPyE
OhpU8J3WyVIwfSS1Z3Xg+34LZ5ZxGXBn6T3zheeUTMuAZWjtxemX144YJExfBIHW
476ourTyCX4ZcE8fZGAtlFlNOcrYnzEPzLxErYGPcJSRDwUh6QU5l/tHyOd5jKIH
`protect END_PROTECTED
