`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZsEXVgRZccN9dL4X05CJvCpO8YSuh0mLzbr2vCrNap8Ha/7M+f5AHixPNpsyj3tW
o93gGuUC2hs5JscVp2MLo51nHUSDlEq39i8XmKm6klTOdNt1McdTfN/bWGg4GBZj
XZ1nG/eAs6jb0UvoaPSxDdRGLpNei/B+zsfpacQzGNxV+iT+8f/xMBgaV52chuFi
a8DF73AEczqM8H6t9fgAJ7ggr7VXOLKnpfwyKjtyY6gVNHHSyyJGuLCBPkJKREEn
nDAtUFZ+007QJl0aQVXcePBpy6htSk6TUN17ptQumM7klA9K+NZ75qxZgfrkqPE6
8HFkHhvmOU2ZJRI5caFM+j44gnEgQ5QKh/ibl1z19L4DEFMtm+CvCQC8kb/ISDQ7
b/eq+g+3ycOR82GlZ5APnMDn6BHH5Nz1PtjRQn316F4=
`protect END_PROTECTED
