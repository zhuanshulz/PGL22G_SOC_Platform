`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3I2IuEtE405lXFfjUJRqLSePpvGlKMSpg+Tf09bAHEe2zx7bwjLP7M8X8yQj0aCI
RV5s3IvhPfcJpyjxmlLxuYj1R1CCk2GrvldwX0qyVG1OAC7DhA4yGreewwsTPoVh
CYa/dZLd7iRPSQ9X0Ys4+FKx37B3N07vO/OTXCTnMjYjNVahfCKi3Y6+mILLeloP
w+k3fLg6sdhApLQ5vCJP5uHWCeFXLHz64KzJJb4eYP3RQ9mA9bxMpO2P3NTrraMR
fqOM4Fhb8FTl3epkglugb2ArUAxk/GQaZS3nScPEw1nmUzADFrSZTFo+tua2nmaO
B2O4uX/1pQ/uTD6qgr/G4v9vxZxs4/E+R50rwVttmA7Xt7VHnaaB3dBky4pcPpUV
Iw+TWBKFzLLSUtMPVJ4IGQWt0f68tSnHsU7q3vfcwGjVWxPdXw79hMGYY9VvpFwV
FR58xkYcto67jy1ZtD1xzuuUymsV/3RlvWY4Ud30Zchpl47ttETK4BSAJxCSj81i
RcA3HvXpJXoYyDIiHNE1atwmgLv1ZuaDie4vIFUu7gtJHnGSPoCxnH40PKV0ruyr
so/MT0uesRlsxRa1snsaxuipRa92jkjMWF1sK/hx0WL597Caly42j5Fh7NlldgSb
SQuzCGaF3hWwU5QoZ/dA23iko/9y0XhmprYSa7pvqUBaQLSlLDussh6DkYfpYyt8
w9vaD4TGu38FtvSC0OWFwwQH7sGIaywqqJy6qcMOUHA=
`protect END_PROTECTED
