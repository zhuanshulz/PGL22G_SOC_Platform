`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VaCu7YJaaQGvtGDbYdIUc87KSCNBVsBoyekCbtMACjxnVw6iV9pTU0DaIBtu7tcz
qFT77JysHPAkO+oHZomWcRWwsVXyTQdfgudQd4MomuN+85btqvaPwig1SlWxJ+qa
JGyn6SzVEP2wxBMbVjUNSzydy5GetIFFcR/kctzE+Yq1OtrBcYagSNl3DKKrMp7q
k+3gFOJVel5Zglq6ZjyEhge8hzIXirBD6hXrgoKhEPZ437EMq09oiowmU+YWqjES
W4tP39RxGIVD1WCscTUUXJCw5spJPpWF89846rIKv1MURkUd/Yc9WBLQutJS+wvS
EHmeX5CXjpTKSovK1nGT1ClmLOv1GpRGI1NEt/46qQaff6BsmDHbPKbiPR7/thHu
FiEF6H4pXxH7VkaBdvxX9nNO9Beiawx3vtZltT2yzLUVblJqOSJK3HmUdfbLIOCk
D6ofjVtCkURcCdjeUHLTJQyrSCO28QPKveuGpi37cdysV4kibXjjJxEZTbPFZSpo
wsGopqerPPu+63+ui2FtPDczcSJwwUfMayR6FCp0U2tuNR2PT3Q0b6Htj3p0NzQu
Nfao2auqZDSxdYxAKEU9m5oIN3ZnwfY/2H+6z0WttrQ=
`protect END_PROTECTED
