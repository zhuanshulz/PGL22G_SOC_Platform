`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
76XBiGg5nvrLEQlPJqLUySOS9pxT5E5Gb8kMHLD4obXRJCjXuDXuDny+AtHe3I51
NRBccCt1TCpVFzOci7sElM2XwjRlegCNDhtzNpOgELfZ3UN/Q3O2ku8BMJz5M/uQ
hT+V1VbHaR2KOLo1HaXzzC37hEE2hKXdrwDRu9Mje77lMsOdwJtaVc+qrruKRJKj
yq9GEmViKxJaFOf4zNl7n9cFlWUSZxlZshQi0//8FYc8bJdrXZkYMs2BcDp30X8L
GylqxsS7pbvDfzaX3zXeYqEAuamEiUTdMfr2XS7K/tkyu7OjFQAysJpduo9/OiD2
Pe9FwFOpMd6FkCJdNFT5DDDF24yq9fCA1ghIXgvj5yM7h7NJQvPdjrbU1MgmB0Np
iNziDMnqmzlbD1ZrhuBP1Q/rFjCAaYsKD9QPzvmyhtyimxoIoeHRfJ5lJoISPU0h
hW5F9QwbwU2q7B6W65+qrgAADWbRH9iVAzKKl84jS7SQjv8CjQLWe+c+VV4u+nVd
7OALqOEdcipKfKTgpU/HmUvrDpA71lkABKxR8VjhW1ahHMcvSHmbtlhmpYoZnNpF
FlfXTNKP0eh9MiClQIunaLzP18HsBGVo7qVD3feGaR7Ax3kZ77yDea7/wE1779GN
4zuh6nh6KYQSSskev2YpiAKIgmWrhuRqQRPcEKEcLbTM82AW0qiYKZj/VbfEFUqj
4vuJ1mYTawrUimdHcmx20LzMvB7jyF+Zv6qIemNQs7PaJGam+PKYuHh04m5MenP9
BolBKFRrgv7MZyxouL+Wm6zq61wEqbFketr1G1hwlFI=
`protect END_PROTECTED
