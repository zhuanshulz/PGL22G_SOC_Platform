`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
an2pYace00aBbPPJuSO6AyZGF8RqynKYBH0ye4Dh8hb7+HHzRxeg3jvGSGXJxg4C
zuJ3rMPyyE3xv2n3ggVRQztiOnGnn/uD/dCCm/ddPZm2ZIEU70DOfdhFK6lLi4kC
oIYFJSjghpAIgts90lfqBoUj+sJFKLwl4HqBRG7EK+Bz8okyGEdKB2+cxIZDsLuG
4yWw0aYtmYR0X6tpyQArjehEjjQShgHH1EoxMfBRu7dj6QjDf5r6uDSMAOzDs/k4
bD5Bc+c8cCDM7mH77D+AT+8hChkY3cAUw4BWBXLjw1Ca7ZiOXN00Xe1u2u9aLSXi
sKOPXrzF0ZkjQOMisUH+bjA604637Xx6kPdp7mghleyqfFxn8KIKdr5SP0U8yAff
EIIyrS8SQC7GZBh0qlYdEmeYpk3jSW/1nclxPoZlRWkd1azpCvTcojhI0Ep9o2tJ
P3FhHpx5bhSPTyIMPusLytGpZyJS7cnx0cgiRC2YYVEqGMOnlTIJCY8b/IsQ6Kmv
tX+wDSJYMZ+9vKlzo++PUSyMFWZY1mK7VwbLtGtk3Vg=
`protect END_PROTECTED
