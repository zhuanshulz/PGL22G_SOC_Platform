`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M46QkQtRF6vssFNd5pHY4mFQ9b9bkwqvEXmCGk06KH0VHnymFjkYsjQgJyhVf02q
rTwsb0I9nrqqb4/7KygWI7V6/wWynQ6RgwHzgbIdanWlO9XhJsq8pM7wNzc3RD1Q
TvqWdzIZb5JV9TPfU3lXV2q5o9OQhckllqtc4FFjBDQeXqLHk/9PYTYMjTKyMQx5
BiZLJPXmzy4cpDmj4ZA/aINSiDmTf5o5Le3RaSN4q2PIhNN9WizJ946vj2Fb85Z5
/83UNDzWbUbGK80ILU+Z9afCZJGuOqkIaTPZ28tG/xNjAYctdgWX3v4hZ8zfZVZe
gCVaKcuvjVjEAVF3tRmdTjRY8yogF8FdU8Ln9jD00aYlL7+gw097M3AAhcVmTshi
2oMQO9kn0R56awaGQ3j2YoZ1S4Nnjs08Y65oFM4AxReUgFOqwYu2wDRhUoj8Ucb3
66UTLaVrgE/XE82nRQcyENezxjdP8O8/pM6cFSFR5xNs/mhlK1tC1xaV4Y0PmxYf
LspG2/b/8GCMsqX3mRVN5X5w6TY4YGg+T84x/9ZY52CWjfmoe3OtvU+wBSV1HMIX
lUzvmX/44nGB1RQbdrUztrQ11Tex3GdKcpBzx2VyfUIC0vF0Js1xpFkQRkPLPHtl
ddU77lGiT2NCRC7qRL7qSvSpuLWlzyjFzdD/cA1HRO56hP7JZQJB8GYtAgbOWsb4
RpKLc21E74bLvj6FlkDzqxjLEhC5H3WshZokKD6xbvcxjj0NQk94cfJK/8V7BwFr
jDMTuIHhIIuMkzQmsE58EwvHFSq6M4C96DDdLOKtdZGS+VVkJzSvmedJ3hVM2guD
LqjsKaZaFS0/5JcZ6ng1/iBU/IFnamtdQrz7VvoA7o//pgaHYe8PAA1u9FRBfO7w
2pGfTJamra73XzqsAPPqmVLcMgC6pSYZNyAy58nDl80VgJood4MMsYBuNC/nVd07
lGHvl25aImDJ4hSpLPANSvA6x/3uZ27tFfXEd4Twbo4cVpJcEB1VFx0McJvjj/4E
z09OBwzOa4XufhMs5JbpablzvyIJfooE2YcERhuD0Zc/SABPEZUeVYdtC9xDrxQ0
FOEESlp8IWbb0WcprQMFlBQaLUO1yQG2WyGc3wfhw4oMSnJdCk0vH+4HkDYAX8Is
YhCX87LqEVmR7n0krRXKIx9t/NN07lqcRoe7cSMkIgTuvJ224DbmDeluN2kGXD5n
DsulgU0z7Yi7lic3S+oCDuqmmEbFoNUhXsSN4CTbjWCx2L9NEJAgd1uj7ZGjcRag
sOJJy9iAX4JHKfVqxQUJ9YoRH5zGoWfz/6tPyjUcGT1ervksuRc7+bvQWZ50BK5c
ezmZaYxlOf9/SjqSDeMo9GDcoPQTNcXqVdx1GgbrcnHmZeYVkz58WHnCkZsF+K86
g/wSPWGhGWLWFUbXXC2OHWZDPw4zfjkBHqmeVf92uNpo7bkyujeB1DYeu25ZKV5n
XMjvPgP2Vqv8liv6mtlgOpsC73n96M4P8uByKnVeUzvytBe7JKgXY14lfagj4Lj2
8McB5zd4GS9QMmzn1fINISxHIbJaFKGQIGaS0DGNmMD4tlLm8g8B6wSzahMIi1KB
+xZ/xqgmOJxU709sxpswk53ci7wnfyYLfipTaCT3H6cbeLGk44Qxmqgjhk6J5wVq
EvCKD/BfwYGZ+d3SZ5bGba/G/muvhTWd/en0MaE4Mxka7zF62mx5M4lf/H7SB+Pj
8+pO44RDb5BXUHVgL9De3KaQh3NNLhTyg09LGumMFoTYzv1TGUwI9rtcAWyw9gsy
egS/d2QBOf4TxiQ/EDcfTQ+bHVFHcc2I6VqOETcOCSKYgQRERP2MWzS6sc5TSAls
fzvku6CnMb3IXcqR64hd5TMRRwNiGqDHSljsMKWmSjlTz21NGMjpt/I0rTk5TiB1
smw/NEqM9mUZ/k9berbeGkVQZ4ZtG/E1wSgGxgQY7NruTNNVxBbD8BSd6X3Y3bFX
W2j6GvbVQWKb0QDYIpVs/eoQSruVLeP561CUACODtnU3PaWXUnQJeVeuQ9N7qT6x
PFpfef5HDx+qRu2aTgIxq4al/jBF77k9mIXtwRt5agnxOdhTWo5E8pKlP58OSe0V
sN4c/iF5vQBv7sJ1Hw6cB7CCZ3+nJe3M+reW+VFksgKes/4joqrldufu2csy4aIo
L9TlHsQsZwdrM9IlUPWuf5BDF+HrFkxiHhSJilhkwtl0eqLPABjGxDPfeLBWOr0J
kCR39DGs5iXM3zUuNLE1AM1TphvGgk6tdRShCm2KJBGWvE58+oyzKHGrir4Kh+eY
ceU4nd3VjBeS+/77hSOqC31SU1V0qmKX27A5+Pm56MM=
`protect END_PROTECTED
