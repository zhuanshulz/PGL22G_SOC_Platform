`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z7LlWqjyhrwiMZ7pKPiaLNoIMNO0JMQwRFM79WEhM9eu4Tik7+mQ5E2ezQ4VNtAy
MVfTEmwV0vbsVVTVxyV6hJCBuJMrH2VzWY2kyBjppYPmuOEwDHNDmQ1VjDJpSWfF
tV6NVhuVBrcY2+IR+RBflTSHfilDwzFrMrAlNcTeWyOdTr07bBnnBq2VJ+lUJjq0
29FMZS0eeWFBaNTNCQUCnGH44ZYphiCQvKbR6LZLfVemKVYBoOPSDHridTDdkVm/
bvKlewOzXYMs4BfA5dhjcEVWoUBdtHEmtQg3FhId8LjTskyVkhjTw2XJiwnsczL/
BUWKirNMN/58iHrGRk8mAjriIIegWu6ANb1t9LhgA15cpZqIFZQGNwgN6/xXTeOy
3vROArQBJ5QBJGUj6xf4OfYbZp/Cn7jXw34wKoVk13SLixEd0FOA7DyX7AuIcX4y
4Wa4rE2dnnKHYFqD0hIi/r2xqb3XC42P0D8vvlxG6vl2CAfQPWmv5T36cAC5apW7
ROshQO6a3+jbj1524m5Nc0Jt4hBYPipw5pDmcZ1e31QYpnI8F4a8lUnpHFY+aG4j
o4tAGNs2fkLO4nQdO2sJi6pqxRFkJACSfgHjpklMTxaxIrRK1KWUEV4yRVWrdxsm
cbW/4qrXaavoyK4jFBHEm6de6+lLvqS8YnBUsucbyEavfp7U352D6Ml4pT3bcx2E
oe0YwmwFetWS4rsyVcJja8MprgrZWSlbaG1AX1kK9CErSygD7BFPZ4uLJnmA9KSX
`protect END_PROTECTED
