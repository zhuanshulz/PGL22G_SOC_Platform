`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Dw10BRThSEyQqnSn1dY5RpsKNbc7H4m0lero1YU9nww7bOw+prIA82xeC0YT5pr1
YtE+SIwLNE8+ho/cEJ0lzJ8cZaDwkIyOWrCnV4tvW0vfsNmYZdjQ5VtRXz4jIbDh
IXDOldiPzF9K0FoU8xjNOboo3TqpJNaO37E5fGKPsByGsjD4J1elUHSa8JBMV6rm
WMb/VczrS8BK3T7p2V3kn4dnliIRpsywyC0ua0pBZW3avZiIWTe34rNHc2SuZs6t
ttQ9CkpCGlmxJgDnO09ZugvbKtmwcSH1AgVyE7imAnxidEY4opI7OYg5P6QrakvN
uG1ik3JxH/D2OVLf1G1WV4ASbnaWNokCUPzOo98eobQYzJIVHzJL45e4Nb5RxfJZ
2QoM7ac9+zKG8HytjqmZo1aAWP6aGGEShLEZYCkCicSgPMLsP3acfQLXQ0KQqboG
HP4Ul1I/KiNaQGfw2z8Fkno2dVNaFOZ2qgMqMIqu2nuKOsS894IaQd0AuYWbV4z8
y38aLzdACGBHwhneu0EG2LO+2mPvjyX2vedFZNJIrKfDHwHXCQAFGul7c4jA/Ikg
/A6RvPgzgEe1QhWakZig0YJNy0VYZs5T3Kbo8qbxswwxmPcda5UY4LzWoDmuFGJy
P3XS2rEQmWIS0s+5Ymn5y2dUAKTIW2bcfcidyRqBM0kuQNao1WDikqjEsanTRovb
WxM5Vq1eq5zkbQ/7C4B5r7zvOlXjaWCNOz6mmVwcSmTUVlrREf38oXq+F8sodQop
n9nFPXc4dWbH6xLR7CfMP74SXhQ0963gw5W/fFAX+Q18W+afGtXbK6NlwYynZdIo
HMVYnWN+13mMyhkUiIJwkdQIxz43daS5Ybol5D0Yd+Rwaz8GbNJL0Ret8+Qpfjct
1uMqCq7aL9SyIh/BZiwvKxoRM3qzsXW83Qm1WL1tV1GkBxxvj+TekTl0Yx8QP0Iz
LH5hFl5iUuEa9s160qjHn625MtMYEgfU1l62ZgtaKotGVLDlffRN8mlGsKDiRCkS
vJQlYkfQW9bCQZOB9FBdGuQR7Z8ES3LeezW3o5Sp114dqQfdvCYK84znVuDxXFll
tLt6mfeCCFArP7RTc8bBf6L3sT5mgoQGytPWcNfcfe2ImSyxu4NGQfg7V2/7C8Sx
P3aR6B/6FGpsc3xYDDWaMSsVr7F61x0g+676OjRg8wh8TdlPkJiCPU0ESVOgSmu3
HJp9/7CxdWo6JHWWx+fKRD0+A+cZo9m9n+7APiDGIcALaqQbPHa0Y2UXSTbEpTGt
YlbTrzqpeQUFBbR5GaKwDBy4i8RdkaSDlf/iLqSvV8rcVOfRk0NX+MTkmQgIkMN5
qmtlsX+SGBVRqL8RHHfrI7jKK+2ZwOjfFhgAfcMScVGJy0FCNg5cTvweuUMj1gQE
eVz12jwC8reywAWvbJlK0C2Ms9DogD+Uv5kpODkf8Y7s7zmIlszxrAnEny7phM+m
+PVjf8cwR5AWYggHmtrfE5ZhZU1cli65B1CaKO3i1aP1ZAIgjF6TPYOc5t0wrUhL
YT7AoYg2Ric5Lltr1DTuVo5NGsAvYiytzKSqOuzKzlQClkkxp7WpXDtiq7PWRZ1w
J1ZV3u3TOiafTLIVq20ia1q/V9IBl2LxnW+jGWHKh8ak2BQLCag87I9P4ibs2x2g
KbN4kZtJX8jkFsJzN3bdyrHfn+aGhTwr5Pr8ylRziKhxUJxN/dATuflga+gMlbQ3
JThwGigtGYbf9CqetBhFrCgcuUlu/XU1V9kVZc47XyQWGJPLaHyJJswropPzkotL
5UZtPCcRLaDUUSueDZwK1pYG9rDI+049yWoD3DPdVUOYSS0s2Y5WNx35PnazTJbl
sBGcCxM35m+TQD7Z0fPvQ9mAeLzTV0qaUDU+h/mz0HPUbkAVpRTpxk7No9ZtanpM
j5agViy+G3U3hbfppUqWV6CsC9YW+ThAP8+RXiSJcBqVgSuKz7urSaGXCEMCmRWM
CHVsWnNwPcU0cMAoktvg1OFbsC/qimzpP1Zu3wkQjCXaa2LQkLd/U0Z5wRsptiQ9
8w9ouJIF6eKp6Q1U15hZjvqKZgvsXYNAoxX3Nrve/mR0Owe+W5ETuDfA6j/xhbfA
t+rk/3ASyyCb+5bRaGyfnek1mCB07fy3HX0Uk+UvrCcR0u4R9aX0HU0cL/hBRrp/
XoZauO9gpGq1stbQBi8Jsivd9g9lVUKqPrUSnWO54krbJoHh01mjFcD+IJJbs7zz
RodI5RJO6dbkQxroQpo4qSM0zlNORh7nRcRQAO1xH+bMXE2psCmS/3Gjxv1icvUJ
BKdKoQQpGuuv/2+jjcBws43TknF5+c4TV5ULIBCuI2Fl381cFkSkO1w0HkoJPfer
dueJ25sN6iBLoTA2YIWFkAb4omRFkpjpQ3xPq4ZBS+HvVPzvQBOQ8gbi+zCM4var
bQeGTEtjGOdbqTEDanlO8U9Nr6fR6YkEUfDvfp6hV5XxXBuKbvMqvh1lPAqew0YK
Mjo8Aur4EUN9Urj2qmef/dsbK2Seke8O8hne1DqprB71uZva/JO/ppBF1QV6NtNA
bVF9rmgFZnb2dkYo8xOL5OQfnc7+A+1h+1+fOLjJhOEhG0nLZ7sHA3GQ87qsTBKs
z2odP3uSkZNrQzInp1D/bQ==
`protect END_PROTECTED
