`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
87ylG5Bkr/nvxUGvPNDdkcwLX2OFOmTIedktvdiG1xEBJTPsafA2kifwuvoYqCtu
qaFxNHLxNE68qj2MS4npLeXkEGc8uRBF9J7uG9e/yGgW0SJf317fPsW4Qj8l3u0O
cx2/he3sCDcJkYB0DWZ4Xrda9LHY1bpIXpH4c8+EV32P5Lfwvau0fsASkiXkeYfy
lxCtaMXsHHZcVpGCoI6gyNvTohks/BcOxQyY7V3ksISDZljxETJCiQgk2XN9Qcy6
a0x5/kEx3vh8RcimBhKzh1jlIknnVvotnN/KU7RiOJphtmAgXMB6v2HorE4vMaNS
w/cdYiP6O3deSUmFEKw8nwN1xWERBpWblCeo2WpHspZtq3XRAeiAojSgVSBDv5vS
flUbmPSDtJk7WXgTBQSDL7P0jtcfVumRCGtKgKCcOXDd4of4AzX/pVz7OamfyAe9
EwZfB0TEikCMKxE+VPiGhtiz1IR5X0k9VD84XWe4wwA=
`protect END_PROTECTED
