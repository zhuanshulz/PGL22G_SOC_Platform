`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4TdBxj57puDeOCf8oR12F5VXUuQ41krZGtSfSg+dbJG8pUyO8kzJnqmhoci4N6Id
2tyPJzxgZWQdOsIRXb2zIynv3JjdAXErPQ0DnCKlVrOIMvntE9MwI01aMEMDSbMy
y++Qp3E+Z1A/tpWJQf6tPf8Qr3h/9wuhrGcGjOq2O64dMU6rmDpKzAXa/7/SHJ76
Kj+ZUKzCQNfC2BvaS3LJxgpxyDKTPpTd8//iso30rHalgEmoHEI2ljlAZ49Xn05x
mI4mIBJu2hizgRMMuKBGPKGsjZ/vKip54P1JcjVx7mst6jIhHrsRIQCzkaksZmKs
OHr2e0vjcBqRa7XyDlZkQJXcxYjdrCcfSHrPTYwSYFprcMFon5l7opcC6OUYgi6R
TCqgdl1s7vhZLwPJY5glP6hsHR6nupI1jXlLQI1YUqUuYPqKLuwADGoIIACW+eRU
Q4GJQ1JhRCICAUWR37GMDw==
`protect END_PROTECTED
