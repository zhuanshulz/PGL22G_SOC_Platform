`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FyevwZ4x4a+dTuVmumRATffePl8zHBlRHmmvis/yFw7vPN9OgqsFboTnOjF1ObPW
HGTUDLGi/47xOIk7SfDe3PjaX6WKDrROAOlC92WcRPirkHrL/rsHm8vQVwJkLfsD
kBF3/soeP6A6vN3Xbp0vtQ4qm+48CFiCCb7ThlQLctzlXNKBIqSTvA4JBm7BXkXs
JBuFOS3EBAElO+4lDyLhtqNLsk0ORPXtaZBRP1HB5vg9gFZ/iaLZq1hqbqE1o257
HcD2qr0PeIjVNpcny91Hax30tSiBLnb+00az1TvUEduKlQsmuCfZm57aR9CXWhnu
GRDXTzIySbySxZ1EmYqx3CBr+Mrj3LkzNn7WivAH9M0YYxczalSXqkV+bsC2cV/m
GYfTB8RawnwwP5ZhqFvVmNmrJ/UlKlvkzmesAyTDNcXB4UgUfIvC/fT4tBf1ryk9
f/EDt3Mk63hdH1K4FU/Vo4qoeae9a1dscpKpT+4qKKoomiG2rSX8wkTp+gYRk6Ia
JOwXbj9Mrz0Q1ze+QFwIPxeGSxh/Pxz3HRG0SHv9xF0y8wn1FtzwoiO76OmDwQHK
uihRwj5JCGdZ1rRRNQxkaZa2rcdUNwnZGujz15/QIwF2g2Qdb8EtL21u8bTj337Q
zsZ3HQ4ZxTTFsoUXxEI9LO/PBdQEUwJK6tRfxiLkHu5huJD5DfccvyQeN8VNVTW/
IGAawLc+QHoQMFcRbsWqfhfmyehKf/xLLl0qsb6mzr3gx9yLUZwVFtvZ+opiw5vp
qGM4v6AnCLvH+vwcSm13f2ykXlBbMbpw+uNATkgHhnuRXoYpQqDvzr/uXLnOKRew
VIkzWEdQ2f1LMZ/NPT6OSVOamqu1Ik9EL4WqyncqoCbTRSCtX8ZHA6ZTA9Q6Ab3d
UBNr7uvvgShSglI3qVDoeMMXg8tfLvkHg66Lk+NELhIwdA8H4O21vZdwT1fbKytn
j5hkxMWtJfO8FcQNFlPrrT2aecHC7cZ6rtwnXZN6xE+cd9sQ4etYSxsI1LA92s2b
1z9VGkW+9UMxcnb0roD9HQlsJ+kuL+9pQLs63xBo7ZbX6ZJOWaITD7MitNepi78m
fx/o+46IypvblO91S9VTpAWc9VzUhGPTEMF1k9g/6slLSvdxsvPou1WX0Dqtk4lX
mlDkCuC1KnmBJD2MEYR7P30Y0YHk/+SaUASenWZpslfOZY85A0s5VxPYJvDph1TM
1v3E5LevHrESzVFimp7+p/OggkHb8l5kLzriixZlw//XHmWhl7Zqm/U+6bDnsS7r
2H4ViTlzyAjYFBbp60Rebm79lidI//+vSSoU3Xa/4IhYC0ISYOjmzsRxVHGSUxRe
md3tQixQZydIsL+QmRWQoQnFx66haW0Af9mS/Wa10eDC245PwFS05zcosY7BwmwY
yNncWJWmg4XGnj1u9thVR3mS4YuIMzD2ayio0pz/fW0DOayLalezhD0wFSOlUo4+
JbYYVlwz5j3V2+HApxndmvPn2WBflrD4vLyb3awn5svFvgs1u6SmSYkOq3I/ollv
84nAI225ybNnSTvBgSPnA5M1P5zlioRg6iioUu6evnDv8LMpp0Nsvhwhg1aioLDS
yluvy4Jvf4FYLcxUVe8V040CWV/CyoqvfPOtYgd1LWxD9AZxlFfaes4+rrNZ7kff
1o4/HKPA3M+E84LQnzsLlbdRygjyU0FvgQqd3nag1TYqv2OVarLb4HZCLGq9vSlB
0aJjHz++9WaEjZC8jwHZYfAlo6LRTFpSOk8v8gqOCPOerDGPcwJrsrnrQkW5vH8G
W7gTSOW7iNiD+GSsO2aOioz0sK83MR3xBsKvPQYWlUhGxEHRY4IuSbsVN99BQtpM
1H+A1MtR3KxnvcqaHkrevcVhlfsbaHUsWuJk3epWbAXlNgNSOI54nwumjFDeDm4x
v/r7rTWD/3n3UN7SKJEoQO1DsyoM1vOsTFJqQTrs5VoKghONnq8dogiPI43sMYIH
+gwLaCPqG0XGr1OkKdFDZoB88L+Adif+MZpSYn6RObPmrJ6tSJd4cC7YDTFnhRYb
c0kAqbIr6gq87eGCR7lv18oQpc7l873I7rDxzysUDZdB93PpNkiNn33lfZ3lNvBF
8sZR+uNGDVVdbcHvF4jkFijhGuh/GXQ/MMZ/iUXuCIaEGFPMCMsXCgxag8iC06/4
yUu4bDEDY0uO7YMcUDXH6zxMRzZi70wV49Q0fuYRrWPLFK+IuscfwpNAV+16osc2
9tcVN4WJ5Alf7KEyVpBgBw6x6iKE2KLpk0kGdFoXxmSLvFmhl4NLaHzeth1ivfCo
jfrI3If0oo2479dDif9498ZGqd9dpa/OyXTOdiLBq74JwaCqZdH71DW6iz/I0n/r
xCwS9NNnp2YtJ3gJZGW51Yld3TmgCc7ATh7LAylC6I0C+lLO4NIY5TNtGpZdCUvq
vQXw2FxxL/nZD1P1sxfFzrPtmVcAocsWUn+V8ACSM95c3uxMl90m4/Xj1vssZblx
KguMIf00+jOV7HSscrpHezLD1pmVzj7seKrgduyqGHBG7seDd72aIv9zkLoB6w5h
BXkD5ZWRVWLPeoetof9WHHCc/WBU6P+t/8+kBWsck+syYg2F82Gk/iOzqfk9DHbc
MU7YgRstbds97Dj13vk3oMe3E3hxS24xDW8idt6cUmODQ2wSrIRvdB1HTOiVBrJq
KaAKQ3jW9/2yQB5RKtGhVaUvrxdnxL7/Oubq0iBuKeBf8JutMPkxvlVjrrzxBfXl
DT65egyfqzg43QzI2+WPA9KY9ZiI1KAp1DSnEvT2iPKhzQo7op45K8L2zZxeKis9
WPpvYnZM4HHnk0sPFOYjrk6F8Ap4goWtXN3eDr6rQrHqLQW7w2BuFZPsCHDV0Y/j
OVZrUiJuemvJO86PDiZ2svHjyXpk403pfX8a5lBjL9IhEJCTOFMZv6l+3lYkmRB0
aLNP9npE/HAm/LsmhlvtAH0/fgsJSqCOxMxCP/SCxczMpB1+fp1u3M7j2qfsI88d
z2dAiN/lVj3scH2TOUuid+g0TPikL+lAtB2FGXX5MVYyaRNQlRxJNOi4WROsaxcH
vlvnq2lm6OR2kpPtmlRC+rl2a7mX/f/09+x0oXu5vPOSBggAnZ5z95Wh8i4VZvsE
LR8W4U65IhNbP7X1y6WrQ7QgaAvmoSoN+dJV9ZWnZjJW7GK00rG+w8NdLd1gzmit
uMnciCrovLoCjp/+Gc0UWr1eUZBJmZ0pR8p0yvidP2v8wtqQZXQsZXgHNHszM6S8
w91FmBRG9PvoF5CEIZdVapGtvXC/muVec6PWlyvpZjeV4r+ZCjsFr/D9GPMvFHmM
q21Py41ps2lD+nuMvBdpcVHRChdM0qBuKAZxtYKw8Q65RknFkbLhfa62b411aPN3
ZUIdLjMDHcRs7GJwAsRtHKJAhdzPOMcu0o/hD6BF4umuIb/FnkIFsDsjiVXQx4Px
YpIovABX+Ttqv3JISu6xOvz3B0xvU/sWvBpaiNVcRWvaekF6DUx97eCd4XI+ATKX
LjUCYFi8US7Yz3YYMYF+3byFZPYx0jiHwH3EG4smDKcbxmsPzL3/g6/ksf0ZjEnm
mUbYY8zEB12oEIHjMgVxDNOg8M5WawujLhMga8tTnRxF2Y9KYsy7bEMqHE0krzxQ
AbJYg+Ysvmaa7L00mqwt1IyzRbK3S2eTiDTv9Ui9Ip9RYTrWVWU/4zL1SQMp4LG6
bE6BREbMm4bqC3LLMLF0E57FkNfxjP4YpbeTqT8lFVuAbrh1GjKBDq7PZC+D5Y6j
hN2tc6i1LLdVXtvBsQ2vweJdPUE6lLNTqmwcx7ywnU8UfLa8fDSAsSIIpzwDsR7t
vi/TVOcDaTaDrUSv8+6w5l6ZL9gBG+51Wg3+5ch7ar0q9ivMAiwJAauT1hP2y+tO
q58zUt9RRq0WiwP/W+0GZ6KJip25oBPfO4AeCB01UzGujpjihJaCGvin9syuX+a0
9BgphNM3nxMMmt+sqVyOr52bfao0ecjUSn1Mw7nIfKBiH1AeEuLHi4y/CSejIYi1
2hlyjc9mlH7ab1PUlZz3lUxGpK2nilGyVHK+oxA+oNcVkrYUnxDgsBlSOY9jSc71
dODkJUMZjYMjdEOHupdXWA5q3GStwxLR0x0zGjUORGp/kOK1Wza0XPu9TxuR6Eha
BdpZhC9YGb++6dQLU5JOzOE/M93h1ok6s2u9eHgdBoVmE/icG3HDWA/nPEcfeBv5
hSW/9w6aH6IT2IKWbDAKBKj8nXGDKs9HzzD1O2ykChQbIgLeyYgxut2+vWtJctqv
4nLYAKdVc+Zq5RboJgPjFbIvq/hFv3XVaNYx5MAKQH4VF7D5U6I95LQC1le6gF0q
bc6YdTcTQJpJRuHuc8oBwIiwUNt6CzGw7kGWcyFg6ZedhiuGnjUrVqKZvet8rZRl
iL3CUnlSUVxhrc7IHHyXo4dvHnRg3vntWWo9p2OJemjYBPOnMCYLagp8ziF8ntcz
+Nq24NLdjaq9s79Fky7a+ugSDCWdUuwFs8r+y36sHjumSZL6N33ij7Yl9CAd4Sa8
zMjQRBbu88vtxcx3SSsf3XJ8hAVTRd96h4Ki34lqX4LRHe0F+QEdEdz0y7f/nvAQ
Nj4qxjGRO4eDLpKa6QmfhR3f2EiIdbNp8F1JE5F4gMRmvUO5SudKhtO+PI3C3G1R
ap7+wY4ntuBiWCKf8GbcyjADC4TmLCMHSH0dqz30yP0camT+uJMM7BDYu5+0GtoD
PYg+34PuY7FAa5O0/n04fKnNYU6vTlBPqNkFCuR3zUDHbj0YcdPHJIMwJRR9CetR
JXD1pXWvDKo8FYQFuDmDGUkBzQ56CBKlteWlalWrJClmsXhau5Qu5W0QWH1R3vGR
cgmBh2Ed4d4WiNLvtDjPG4kPbvRTNuKmfZvkEKsZ383+q8z9af7Bp6QfuuXDqCT6
l/sWoWXo/WAyFqfcgc5gb8nfz+UUtTDc7yC3wL2vf7xR3yPuQw/IvPz1lwx3MnXs
U1RkXgRElTH+/TcuH+r0VIMMLB2SbTB2QN8VuUBNMWBUd/XEo/kgIUsNb7TeVG6D
Wm0Jienyfzsk3D6RrxmyPAsRZhk9x7pu0g4Tiw/St2bholCRUu2vchhYKcDW+V4j
TRI1uNcEuuCL5NBSkPLFjlxfaHl91RpIYdWdk+qUkK768S+Uh0Z4shJbdGCdAsGY
sHfNkfWJsKRuKaR3jV+MtfxQaxa9fLsnQQM733u/s5QDP7rtvJITren55k/1WztE
OHaSmQrdWNCOzlyYTod7UfNWMnGWPQ3YHIBbu62DMElSHKpWEu8bMkhWHUFJAGn6
1Z+pyjtP4kvVXpf1NhcycWjPfwoC2/dW0fjRYtnYUGQY4WQb2Oy19/JUTB0YPLwb
QCkuEJnBVECBhl6FJvXORjF5ZqnzjhzKdth+3Yao/V5SBlVz+CnlMl2AqoEj2Sl+
wqIi76fDdQLCXOl6w6eKIA26nZp7KxhN4j4MEOJ2rkh7iMWJMHyI7M870pNX9kpV
VMzQnJDez0ePFbin4ym9eUUWnsIURiLfzCiBny+F9yrRK7G7uBryTg5ITmWVG00c
U8xTDs+c2XW28S3buzduJGfFgmjA2iE51cCdAYM6J9tM2nYDDVKiBN/pMuPhX4N/
zNm8URkdbvY8nJmFR22OA+BJAeV4LXEppGFakXERLBptTxmtke+i921fnz5sDe+R
sq5hbFuOpcrNRSA6EBAG5ycIZpoeYm5hi7phv/Ygfwn2mfvL+5/aytYNvSx/nCoX
zgGr1yp44SQY8j0nDC8TcRrVw0JXvcPqgEpzclQ/9Tobhsq8Bsg7G0TauSnVu4c9
r25o3tuovEsyySGObOvWc5srphCBdu48ZqK4o8XGEYGhmLu9ZmVYNQdprhAlcdDt
0krg8YIpsYJyf08IXFcTg8QiaMMVNe7gDoEXs+zTmx0BLDVoQRdhWpGvjgxzMPPJ
RHBXYcX5OsosAF0FeiAzmB8aW/zLtpr07PCY6V6CkZGkgOQ/BlGt3TPNd+kwQXIs
moHwiqmVCDm1pUheMHVBsWvhqxVzNLha37ua/sbVBX6tKM+Msez7CqK6PGu4196Q
yivIlD1WjXBN6DXYTxI8VHvt3VoawSceLg7Qjja6OB+QgVCqVF0YLc0RyFEaaHZ7
`protect END_PROTECTED
