`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ol+ezto4b4c/2HxPqpVrahlABvXgOFoQR/8bgEoJtexBMy3hrFdoLyTsjn50yvab
YXEYUaPf6WLIeDMAA3gHQXkPbe9E1k6+QlJVztmxaCacuAMAUORwTQXh89ayIVaU
mcP036hkEdKmtpGTM+LBlNV6Lj4/+eq/gs+WLyYuoeQUbRfRpnrWJNPgCTj1BU02
49lxptykao7hrKs4gXMmaRm6N9lL3LZ/QffZQSDTK/P8zz4SoKhPqR6GQPN/06Lk
OaR7Pc71JdtuWmuG/U7C1rtbqqhO0WrAUqwXKJP972+1bccgugOcno5istfQCgHD
7vkiIHL2TO73YlkOGDw8SN7P2qkLyKkiKhq4Q15heUZOEVbqKOokTTk5o8tdL2m3
RNk7r4pjAmwkgE51/BS2SzZvhXX/IZoMHplViBPFSbNkoyHkw2zuJPvXPnOrCrR4
8djn6JWtd+ZoSjfKJaGHcqYSTDm5809PzYYiNcsNCKQxqV+ufZ3KoYtibI4v3VQh
dpbGRmAQHsXSagDMvMGvMw9sDKNEmtJxCXuXA/W/XwftmEVMtf0AJE7ouOeJ2r76
GhIrA0SBILO9zIp/q1aybM117/H5iXCYOOHcWrJyrbvUEVvaxVxPH8Lz4R4SWvtU
3ErykGclRxgxXLNTw+8KYOrXfSi91ObKJDOMC7x9U/R/RYy7rVpsJTDrZidq4ip4
sbBykLMgpwzOXkgJy+Qj/C8lowJixbJv5OsVyebd+ns3FTcK2a3hLEs1ap3JkhBE
Zc5iH+A67xd+sOg5SWxeuC+ViFuCrNM7GXdHNTrwGHvEr6/uVWCq6n5H5viPSNHm
F+6c+2DKl8ivQLz+W/WJex/aNqb45eyLtb4ltPDlZAjTYEArCeD+sR63KlhiRCvJ
RirOrybZ9K3XowsXhlH45gXzHM9grTbBQd+Sc8O/+cAp15YuZTHKLLidNALgWLmf
+FSluJ8viRK/MQ2wNv6/1zxDboWdgdCT4qtjr3Du+MI/SXt30sE+68BQMY0V2pzl
HkMWKwhJK6KjVlGQEbTovMZPJHYvBsoxqwPSu89jSdhnnPSzu/6vuWyFGGiWLv1j
4ic2QcHnFrRjBq8P5PhVpiiD8HcVYq/ZIVLn7u8Mfs527cw6S0QUietZgOeBw9Ik
5nmhv1UOINrCDc+wwEn8E2Zdb2WGYrdTW5RtoDiNf6yhMEBxlpShLTLws+LoeEZm
sPNp/O6RCSh2iz91JSlTNgtQEUZp5r2fZaJkohu7xm4BJ+KOpP+g4kJfFr1GadYm
lxM6JuLm1ReMFUADNbPLKOpIwo+zaQpNjBYyV5IQZDJaxXsMjk3McII/FYjNafPp
uuf4yryb2LAuthaqxoPiieK/Q6U+/Tv3iAsKfWAH1Y+dr8dqJSNRYVieg8SZF/Ep
U22INH3DcKj5CPIGF++h0U/bpQ5W5DMA6YxggbgWG++sWh6ii+a+n23jSxlPNK8z
x2r0V6q4AhXmOLoBVtvW1g==
`protect END_PROTECTED
