`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fDYLTp3yKVwCRD6/QjUZSEKDNHlVpYQ2udKQ68uDU0T8ypBoNWD8Q7cqECKa3Nku
MEkf4tZkyyMCIU1Mg6c4nxm7OdMN3YAV3NS7/s79D/o4GJbu5F4O0uDbeSSeABCb
DB8ZFI/cKPtyZSKLVOegTpFV9EOrZclz1wGX1jAuaVeyGuggWng8Vv1SL2G4ifGp
iLBOr4oP2bim2/wD/RVDYIjOHU4lilUJ9LvHlGKeH4p2v5tWCTBMTKq/rNfacmQM
AHvNEu81Jc0YXPnYfczym5ZF8IiJiewO1RxTL0e9Vu/Z/An71GswWNuMza6mNPYS
6hHQzoh7UN/4T5sMDVM9B8NlOXMy1K8PiSZJOuxPGNT9PcGks357racbKvTGQykq
HKltddfqFZdg5jcT4vmH9VPU8nb7VfYLMG9u8nHr6yNif3xEzNxOZseR/dWewBDc
ok+ZTLsWJdjl2b8k6ni8LgRNHLDHtW/Pjm6luZCXrbuyEWI9gwaTZ5qwE6JzahFu
ulm07KZeJtpublJrLWZOXOD9Nrd5aGY1j6I76y5bv/E=
`protect END_PROTECTED
