`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
353c+HgKslsZ+Qo+05Q35YsJpj5fmj1bQZoQWgt6WIfGgRZ6mzmvbHzhBE1ur5JC
9EX6g43oLoaGRLDYUmr2D2qU0Ctz45iOcL25S8jNLRIqj1HqgPvvo5Nz84TZ1DL1
zkdgzGbawTzkT7wEwdgvZjua78885aV5BhNzKojFsTTfoZgztKeitvae6IX1e5zv
nP4diCmAUdkuCnVVZV6RsqgPi0bMKFMfrio8Kwe5fAudju08fUb87reKI9pB8jVV
Nhh82WETgwGOcvBwMi5UKKtWpDFxRqqxu6oTIhDe8huvg8/N5SPvlOf4kKtHOMqq
vNdb/jXR2nKQ5socCNJIHl0TRKkNuQB1dkQPlnsFJzsulCKq4YSctfKrNEADt0Zs
a1Tcgv9ir88OYEkMcLIV8bNQ2dXrhvrPLr5u616KDy4gn0NLG0A5xE+RrD++ryje
tXh6uunkCAyKKOKCMczovshJeSy3EVBrnD9dlidF0hV6w20I6YBNToOOURL4BrIe
JjqCFghNDxhacgdscQTX3w==
`protect END_PROTECTED
