`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Fy7Xky8xbBVLo033DI2YQVYhcdYy2zGSG+XY+lmtSjp683flia3DmWG8OkTFDXOT
9SJ1tpn8F5hykMS5FMl2o0Q+53+jkmZEt9Pg+dkZsOPj9RIfH4ZTRZDhlKRvSBth
CjFmdRoldiLZ8KAxk3j6CO8T5h4eol0HTVEaEZfiF0M2eMA44vPVHDKaa52D6uKO
Eo7+2gw7Nh/ARRIDbVkGpnotDh73gAMGZcu8SG3ERMGhovIV+5rENjuNGLNrtGHU
JbP2nkK3W4d/in2h/y1CorHptOglgpKPnDFHEjCadoWT3iEtFEnBBrzXzMVXyMOU
p7n4JtCAHpB/itBrRXO05QPUX1gLdtggcB5n3lX2rRuVXhImJmfCYN5kk33pN1qR
AE6iKVJgPD9a72hcuus4BPENKFTfYRgFqwV1SRonFEH2XB/g8Jl1eN+cng2nN6Bz
UBQ5662kuqhB+5xWp3ICD+0TN0WE/P4idQgOSJ8uDWB53zwjxci7jsv5YhVCh49x
g2UrhtSy6FipLunqxDf5QnKPR25e7CmYS/AmumG+VuCfyZaKe1909hHWMn/eq9F7
IvPPbHoY0sFWAkzr7ry8OxCPmuPMdpQDybJYJpTVX3niTHigyJiwGZbLA49mdiYK
ah+ZU3EGu1wg0M4xsedwUY9CLtuKpNX907Jk1l2eCNtqiJmSjaOe2tPzvb/b7ChP
p2S7f2Yoc6ryObMIPbfP6JzHaaxCIpGxHrn+ZwKDBpMnHzM5d3dkt2qHCFtKkMow
22nagTnbnEaCaZ9RRa0GRhKaTSHRPkGfVF+m1Wxnyuaw2TXZ/Vcmf2Jr2ra1+hcD
twMZG4WfEqu86uSz0TTCTaT2U6vBDGJvH/UxGc7lMg5CcPgT917krUwABAAyJfRD
XloCmO7LjByQdgfRZ1/VdDHdgEaeYUdy+2imKyyTAgcD+b/5ff6b4NQeOZa8JpUu
vvsueu23BbZCrS9408zczR+U0UXMa1SQvO/r3RXT1gN38tB67q8Hl6bmAEjGxB5U
1Cv/xs/NkdHS3LfEH0CfUBllMfG7tF5tOZ60dvgY2ZrUfOZu7SllgceHn8OVKMMW
DxNC6kUfuSlsvLJKmG3u8FSwK1vYWQbZ2R4vg1OvewxkpLxUO2CElVeACzeqpjHA
hrnjkuRweGgBOpG2z3dhY38645I5yLtwvCrv07a/Hh5xZ3zPGzblrWV61U8PpfBe
+vTPxg/ebJuBfzCe774srhS83SE5gARMsrwdqn+EM1C5mRn3sKytyoJ9Pr5oQ6AN
bDkxJGbRlJ4M06LMXCd3iN+5NPHamDT/aqXdD0kPzYVkTUW59HoJQqQn0JpW34em
jKus0UnhkJsxFxjWVf1on4nvAILPpNevZvfXCvi8QlYAMfL923PnsHQ2SHLJgo0s
8ATutIGKcIIM9k6UPzH1UQgY4WLq2evK5z/n9xcOJBoVnoyHupXsQ2dUgkW1Qs4x
P+3EM/S1A1vk/GQmcw8Nqt6h069akPiQfGu9RgH6xYaV8niDGyriWwdZA+s8SQv2
PXByuJ9PjQGWIc9vpEPUgpKNosHDajMA/m3SVouaxWN05xOKkfu0rgru0UnJ/yBC
w+rHZ+PyCXhBCf80PAPHXtBaxb66cdMPMYU3r3kDQe9kSieJ2JV4RE4YWMle7/0c
r54yboMEOvryiFQP0OWHDNpqcLf7rzj8kqjNbOoQ0yhTIY9FFwWxEcOm/xKqXx3P
y7pJTLS2HJ79x4S/rLtRl/j0zrcTpG5LRuOdYwv0s419oTFHlR6Ha1PK2p/1S/fn
6ihboUgRugQUHAlY1U8HH/7Kb9g2vcO7m/hzHk5es4ddiirhgpBi+bT3cM7tvna+
Q95NSFPRiYhq34U6oqQYREPNdX9n2nzIh5G/zJ17fQDdkCcvswc0XdGcVBFUT2I5
vbSwY2h7fjE/4VQQQpQb8/F7I8JX8+SWhjJTig/3yLLGNN+5Oxb2rCxHTf7+FNyh
aCRMJEU97/KDtbL7+c4ehjzEnJ8J3DG+DJWjtiUvIQhswJACCYgnzZqYK8gNuMFd
55dVff4JmdwQolG0FrW90WqEmTe2SjY4fEQBMTh6JIskGKI2EN9J3ExDZ7Bne1c2
we2LqZCczRx8GpG+Sx9HoOrWd4aH+XFwbegiF3sWiGZm8EOL72EwRvvC1aaVymGU
`protect END_PROTECTED
