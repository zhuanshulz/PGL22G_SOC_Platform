`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ti6z8pychiSGW9d9bXzCIfNpaPKltvSMwKg44dgUaDv1ZfInCCk+bJRv89dX7+8V
50t38bg9E4tE/9M3kJwBIyABDh3IUzflLN0ktiDE7akn3ajZrqlKb4LmotFmwzoG
AKpXVEE3NqoBXVdrC0kbNzJirqi3MS8AGknJo/LoEKXUYbiNcEVf+JQJW2kwzF32
/w+yVtE64/QVv99q/SJf0b6uSGBWGi9G5zqkdNIzpZUfARyauFFfrBTG57NUo+Pd
P3fCYCfPuWcbMQ3fLKKRBe0MFMsWab0euABvLSP+WUxXdJg3LqBfsnho31OKAbhO
96kWdmsoJPrSw1H+UzSmL+W7sYIMLNSZYv/n8KsDMcPiCJWa/KLPE/i4Yi1tMq0N
/yvfikIBcCj5BmETTMn8ByVyJCOTGSMyYluy0/B10y+UhGa+/eMDFPhGRmNERC/0
AFbNLePkamMTn0xsoKwr0EfOMHPgcvVABkLzPS3h2/ucFWXBPPQExOt5NKthXUYF
oLvyA09D1c39iNxYObUgz+sZEOknKrEqlCXkBLuh6GmxA2jvnqeZ/c3BKtBpKoyA
LW2x4ppV5oGHKBLh10KFLIRvozHlOL5bENARaqovriEq71/C2hgxXH1eE9DySSCh
Z6thMLlJEXzmmZb+q34aoF3QEfciC7eQDc6R6q6nRP269VVKhf5IL+M8qZHdUekz
I318K8xj1gW+4j0z1+1CB8tIUy8byZ7+ZEN2tKvkbFvw0AB6oQWWc2TCozbV5pQd
obpGhzTiPu2Us6Z7bn97RxhGOx66fVyqzvYsx6VGaraUpPaEG+CUwsJElQvpx+Bb
CJ1zLhDLeTWFIQzfKmEHaTjtAPmOfADj5/+UTvV+S7g=
`protect END_PROTECTED
