`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0hoVG7mlBGVpQOJDBn5TIHgQKdOIaXfQYBek4ORh8hGpxEshoglNOkZGKFggMc2k
hfSeqNPpU7Q6yFXlw8KaB3hseTlBgP/zDQZzdRSslqQnsizfVYNU5yvYQ9OWlZW4
AGFdm4rmIiR4QgR02EiD3TtUYYhpJhEEehezzkRyT8Qfn63ANv1DE5YwERgh6Ntt
KSUJj4A+0DOUuhBOHWCnWW401IYXHj6R/WRhCXrk9NLJyMAj8WFcciCh282GWLkU
d1uOPA5/0y229plqKsUBg2xjSB4GMfMDn+KzKsqtr4fQlOmQQQcG8NORsp8IX13q
Coi4qvqWsD8sBCSpb5mYMaDzmrW4tJSCNw/7KUhuRso5OPHJbjNCPPy1J+sKgheb
Sxn/YseQAgRSJN2/PL4CuAiqhH5fMAWqgKGboTY7T4MODBqOVWstJ0X6gCCag2SS
lat+EGIp/9aqgmqeh6gqNR2ETmYB3EeyLk24kE6uRKheutANCneiDBAM8Cf2Upjo
3zbWoNVBj/a1DhgGIi4+e51nw9LZqjWeFuT7v/XUS5qdCSif+Hz0kHpht/QlcJOx
L6O5dUOJtQPI9hE0INKOiUH/dU9YcSHhPjVXSY25Is6dmHmLZdKZBCKvlvnuZJ2T
nKFbrTNiQFLequaSQQ3x9AxhvJ7jGN7h+rpJR8TZgZMv+RgWLDeICh4zRzXvaJrb
OskH15zkoEsaaPsICAC+tBUv4gWuxqPBvjyo82i503j9zgOsx8u8lDKZr7s/C7ec
63vTWV6tDpX04XKAnBUaIUcvuYQ/tV/kq7id0bl3J8sxvvkQRptRxm8f08WZDKT2
t/iYG/xAEMNfRVyjMRa3ukGE46yDsTfY3mHSY1D+eubSIeLn/+Uq+snzW48WSS9O
hqXRvaACoHLJgDEJiwNWyJc/KpmrbagzfQa1yNPLo4IBogOT2hcyY3jMoichCY3N
DhmRL6tSHsPbYOFUw03gWB7Zb6ICPDrCFHhuGbjm9trzve1E+8XQZ3SeN8eAP7vb
AR+1HBMZtiz8GjbLOq7udZyrev2TO2pVLblhOORsMzo5NBjo+86kPwcMYJMqJhL4
e18PLe1bI85Bb9kLLOjG0lTNZpcLUw2N97MlJkR5bGVNVZUma4A4bOjCbP5Btfm8
vFIE9xgjE4Twhso8wpzMmnXiMe8+OMEm6K408UwWgzNhpJaZW1evsV6LTjEnLLqs
JpyvHC3Ty8CV3TS2uUEaMtyyID/Qq9FgeFhEwx9ZkXzXHbFT+cO2/R0IJsYInkSj
ec/mLsDNB9g06zIctLyRdkeCW8ZrjI96RPfo+AX26IM=
`protect END_PROTECTED
