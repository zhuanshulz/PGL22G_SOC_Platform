`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9fIX+vfs2m4HS+xCSmJNKuUeD/zggGRnpF9AWl7C42JAU9X4RmyUy25EhIYGgi9+
JASX/Soy9A437gUc7fTQ6Aj2/BPZe9rU97jif3TbyVoLt/syqzOL5TskJa04jLXz
EHaWA+DTd4GgjmDIEr88nYUasAPm6tDdtrti8JCDmBvJV46RZLpcY39JiDoYY6Ic
W0lUOs+YW18aTlpwA3lxRGesMPBqr3GVN5LIYGouLSWH4HCvXdGEQxn1qhYxzcxU
Wo4r3QZtHVkJC89on9uJz3LQEJ48C63bTwemvgRJJkxJRzVvzlXAFl4OzUW/3Ap3
Gx18MqKJwke5Rmh68MUsDn0SxR628/Tenm0w3Xu6UzlrQBQsAzoIoGfqfbt+KkVS
`protect END_PROTECTED
