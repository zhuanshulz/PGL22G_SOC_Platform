`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sa8Kzin7uTXbVG8LOMhldL+Dk3u7JpV4i2JA3LkleeTyDcuHK5RAfJ/+Utju1q8N
E+D3oYaaPOkjtDw6w757WEvLEg2izmzcKAoKIJo9HKkUmWWLu/7WRjt4rNMD1eKf
M7tu4WBPjSHrJ2vtd/KNW2/xiqjwct3CH1BMduYcxdh+byRyfrSLQ63V+1KhPy0B
lSKvP18w3s1jWtG+xeO3NVQK7Xl53MFW0buSEqmz9S7mT9mQYO6yUxjWkOWmN9Jd
LTJrjshHwQSJnR/o8GC4ZA==
`protect END_PROTECTED
