`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LbD8SjuUFgFiUPimP2PnSdWxxevUFpbGaUne7c3JdhJ2uV82Lyyud+dMvhS43YGa
EXOG8bZ5RkTVQfxf275i47Tfh2jRt4UJ9EieBypRreziArANzwTozb58zuKiULdZ
R3UnZO4PrpQA9DLBLZwVVXPowsXEzamnXjxFoU2GUEsNyvlWqtZWAaX/q/H7AQPP
ZOJkaTjzRJQyLGkE31AzyZCzwMsikAfkGZomr5dobQypJFRAinliwFe6YiZfd9EY
FfotdkmyxD6Z10YvsWJmr5dR3G0RsBv5YGTuajruggDHPlz53V5ImqK479/Nu1Ec
4HnAqsCnt4Ih1E6hTnuDbMJxwYa9ZWVija5Bzag5+FanNKNN6Co8u8D2ibTnw5ny
HznYs2I5FeSJuicnChyOXQ==
`protect END_PROTECTED
