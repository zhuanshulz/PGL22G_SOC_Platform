`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nWqxiMPxQE8NU7dNCC3fjNw3TpdSS/vgl/ESsJCgGJHkBYhBIsGbmq8BJvg6KZqy
8XdTi7iSKWgLlpOCVv+Qk9Oo/1Wgo+nR+6FvAB71sbIIQ6xrrq6DIZgARZn4+KUa
7SWelEUUXMWwEU5r/5SVs9XR11z/Oz1BMLUH3S6WJaAToYCNNSfJOPcNERJIzkJz
CzYiKtaxQUA0jpRn38Z1thLrUNP257RNATtHsSEJgGyM8AqVZuJyyrKfuKIZTlus
qw1rln7ci7WRQZah5OWDPun0+i52xeQjsX4gXRK4QHCxSyCxqP82smfrT/q6w35V
zF8P/SNGpYNXnHNOdeOXCA==
`protect END_PROTECTED
