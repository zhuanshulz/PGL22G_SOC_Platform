`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5hw4HwACsAWTITm8Xhsh0OFmCcDpAkVMUCIGWQ2iXV1YLCZHmfubY7P/o0/h+XWu
RX9z4AV8FPSVcLG0S2MV1LBevb89Qo9pxjEsJk1+VECH0p+73YKvAtjwS3OCVLLQ
6bWQXq1HK9xW794NQuAqDog3Gb+kKW7LRdRG5nEtuCbD1maSlr03ZlKzoxnHmEPt
aMX1TsHb7WUX0Arakl4GvEr3JAGMdu1EOyzWjOFvTSun9KC752qqNk2M4eWBBQkX
K5ejTUqPXUBq//VjHfcAbwSni50wKTKamKxAAhOMlTuKMM/03lN09OoVHCvTpWJ7
CvZERHcAPuKVPCxz/IQJZRpij0VYX1oz6dVxvpXZk97yLh+V2wJpuRX+s7pHO37y
b764o36StGGk5Gg4XL88y7V0S7zYUoDSHmFSYXQ6ceauRdlrCNr7lU08n1RFLGhI
SWw6nT/U7pKi3fAIsBhazdCB9xWSzeRVh3eS8vVNTPa4FyO3cC879qF85qGDPfbj
g5vbMV1GoB2gYdWMNbuBlZ/umq588tJ5kHMvXSrS6cRIUxINqz/yjKKwaHzi2Tuf
4BVUYPJTBUVTGrrI24G5sxFo2zlgkaFZ5oeK67Zfe4iZ9HfrA0wBiXNjMt6s9VmB
SszzpCw4e9H/1jh4jeKZrw/m52Dy3PKdNWNkfKHVwXanLR8aleHX5w/mhK5mNYrl
Ofx4VFwhHZ+oDSsi6s5p0y/K18mfNPsX+6coasA9WlSMO1SN9i/uNhRvUKTZW5HV
O/sDqjKWIv29UzKNYxknZnFCH086TjYAiTwYLnw9YdU8ngl1NupSkDY2kK/oagDo
wfpMo5yXzRU+/2k33QmhU0QbI40wa7Z6SuwJxB+ddTeEaAP4cXwfRwd3QCGVZUwQ
wUoJ8TNgXhl1M/vs5rGqW8Zs4yMk0bq/CTj9Zj52aPFr//8MOkbl8AgrTyfXbA9q
hFMTK+hWDr75dDmDxEOSiYN8XMxXqfk/A+th5mOlZUOv04pLNuLbuBN1ScH4N0p+
4umK790+BIE8kfCSfyqpACi8Y8JdrRK4NSIytijbRa7DSYKZMVCl9HJJPTiljYt3
kZM+h8M9rd9J1oOqIq6drYGWWLP6iXg/HEcS5ObN9RYZUphSx6uABkDsykcGLGUV
bk5MU+4mhBFefNhIUpC6YONZUtQE8ACfV4GivCkycoRHfp/bY/2o3EYCPeveJBTy
92xz5tZNm7+pdLuQ56s8PiX+HelnPbrEoBVwO0+jiA5X5s/A1+NgOMfTw7wb8uoq
kto23Olm+/wizvsc0TaK9fvSOOBFUy5ay8H5uMIUXmzDTHqJC21pLk1lqLio45pj
NL8H/afHXsc8sk0aqI4iTHB88CrmbCRz6iElg+Fs4vyFfzqG+iOrQnr6nnaQgfc1
UErWqPHMt2rtYJCXRRWtTQIyzddKICGlXfrxGyIekVdRZ53f8BD2/H68dbSkwVEe
50AKC5n0vmt7ZJ1NK1bEIKaNyPVBsBUgSWTIY0UgzrOD03TzBJDOCQwhMqDm/p2p
X084D97W/TqbQBgLA28yi59aKVaObu6mT9NBdzIx07AJtsFT28QbemXkmeVzr3rm
jrKU4oFEerImkvu4HBVfObqZYeOPdbaF3+uGZFQW9kyAm93jOlQqK1SkJq6wzR2t
x4rUhNRi2RghnVpAlMZRlZMoMqtnzNtKUXMwpyqjoualQ3h6G9Xa89wf644mGrkJ
L4AaGrVfCh8KHS3CWcnOBRAZcbk/oRUJIMs4Tsg7mc6dPD/8GqB1RjM0cZuha1iQ
`protect END_PROTECTED
