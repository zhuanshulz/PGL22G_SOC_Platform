`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TjIdSm3WfbVdhGdlhTYFWa3Og+M8O2qhjaXlJcc/9z5xPVEwQpmCGBzVLcX/uHDs
mr3iwxoq7/hI4Lytf+7Mp4ZuaaljkZ24nA0Gbuw/EmUU0APH4KIsOtxkjFwshhSG
OdUdCuoUJ1OsARhUQCK4ysWc83Vld6QjZQaTjWKmlsyAKuRmH3trKhOipnZkF/BV
PflQJDXZB2l8d0JxT+TrvQ7/8gRIwdV6y+hyCN0JG3Q0ZqJ1PuX5cHrpO2X22bKj
zBIK+PBvuESr2sRI8iqidemw5rheXWRVuxlcRjNTmw2q2/FXkyEK/PxGAy0AK1nm
NoK0l5f0eSNOjEx/+b0W2GXw5jrYpGFMO2fRYl9Jy9bbKNtFGLqfXxVc6ErcX0Tf
+jh3hjwxRuSachOAJBQOccSbUB/ZundPGHR0izEVSxP//ttE5t2F97teIB7qNqJk
Q7ostiNYwwkhh5263/Y8GQwh3gKGeQo565v8wkIFstVUsQwba8SQ0BxAwuwu/n8v
pltTaVS2EhxYlrI6j9XqJVjaVtXAquAspVRWTekCM1aqulycLObuS2UhXOiWAiYw
HtaJLDyW+55HpEp8B7CUojcj32NbQl+HCTuti24hoiWmYDY2DWlz/CzgfJAcDj/m
k6k+xxWA0LRMHvJpC0rN01d7bf5VVclCDtck0rchg7ZVdKvEfE9bSA5Z6i/I+XAH
JlZTzmpie1EChstyXPbm7ZqFU6B4M0wlPBlJK1ZfVZiHwaXFRNJWN9TJpTQPRhBg
vGCLrZeIKUVfIXAoRCtbCSTb3EHETXqGqu+7Szzuf7stZInQlLlV+UEZCwPhBdDz
r9wN5tvbBM1CcpeR+9aegSI2wXOoEUnzk0i5axmzRxdTCoAAVM0NibLBMPgzoM2V
Rs+6/Rj2juGbxhD7sxIqwg==
`protect END_PROTECTED
