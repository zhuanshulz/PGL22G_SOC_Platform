`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MC+J+FgkRTNJirtLgomQbYSBE93L/iNlVLJTijcKSOBaIGc9XBxZTacxeSkR3Evo
PqHttN9OeGni4MJtpG5C7z4P4kx5/eDs6sz5CQQ/jLfOdHFCsZDO82qS+V9HOT/L
8do9t+c5aiGxAd974P3Ws/vH7MXmc2JN/NQGf2FLRA3S06jnw/RgkyHtjSrbiIlT
JNZLuyqCKRnhCw7SDNkdWeMQWK18ZqSIgxh7muipCk8q3G8yYh+efWJERDfxAWzD
Q2ZOhKKGd1tiyWijhViEycPigCbXHCbW0BNVtnsffd5XVcoS8Ij3AGSBaK3nVdmu
ZnS3L6LfUMgqqhmhSPxZtwivzIGhbqz+3EjngYV0DzlYscFJbeYVE0dTZ5G4s7Xl
PNTSLxzUW5kn2M8U+BXrlD8SbM/jp6OZuN3KMkagd5C3B/a9nFHZl6N0zZzgvAfB
PBjLkiYbzuxQZudqBRaWTUglzkhksC6kvhaGhYxrBqlzUqF+E5jryAvF9wrFSmx5
EB/95ietNolkIqXv23Apn8hVsCuJc0MOiQQb7f4hr3E9tgeBamU6P29Rq58Dt+Sh
/jKS+o6Pmmia8ds103Lqg7rMkwwS6BFxm/sboHn3wRnN5Odc9hH0SQPGIxaufQN2
mTvcFyXEIAeJQRQ4PFB+5Tnb/N3ePQzyUzvl7+L7SEE5aDPB7zBZiJw6x1o03Qns
Jtulpz9Sr02Zmz/DAJE4ctQF+/m//AjY1X8FgrxlRJQQ00/ZA0871mjJilwD5MaW
qiDFL+gtZ6MBcXAQ0rRxBYTDSXl7OpXLp6DpZBZ+QlOHC70NdXGRLTlv8dmyGlmG
0dVqVMW1Wv0yAqKE70xRdcEn8NC9+qauFDq9qoAroZDObpb/LYwW2LZ/oeCThQkX
NPc2oR8hiDaobmccF7IBfGr1JyU6JB9J2U0gsdpXW16RzKcDEoP5697XHIgXQ3cr
KYS7UpERz664PCDe9sbE3IeBSROs0JkaDqEosQxiOpuCfwnrQsC9De/2RelNIY4z
xk/pD7Ej6LfcKnPUbGRDZr/w+TuZSQ9LvaOFiHNO6fO4z/gjfh5mCIE/g5kuAoBJ
0f122Xt33D25v/fEvSza0Ul7OKn6y75kOyVvigoufZK/Qj+tFIv9TRzaBuAiKGKD
acg6P2ZLhfHyUAWnfm+9ucL//jIt8Cqvj0O5ysmYb59rH7MYESAa5RdTXkYNGr4t
pDzExSZNbjormr4+lY8j8So95KbxFKSnYHdjufiW3iY4zH0ljjUnNEVb4s4tDtH8
tS0/qCGV8H/ZYAhfX5g/zgi2vmxtEtorMPCzn4v04T8Qtr/tKFq2iOqLFATRcAeZ
kKMoG87m+iQu3DQ3jRyRT8PNC4vNJoeMg6RuiluJJFvA3WpHtMqRR79EOHpu7efc
qcj3fAKPsegN0KmLvs4A2omq6kxrA126eUg3SP+IudAg6Az2VMwnYZiqz7u5J+cH
YrpmOiJ1IMtweuC/U19U1Kp2iRtMjM3uFQjhmAv9gOVXsvtGxKiKpq2v5MLfIg6g
XXWbWkiEOKaYYc2F4+xdKDC25OnGV+tiNCqTKmuxEcUkaxf9rALjIyi68CrpCj5O
nholtKKFFYRjN7N8WyyhrvFB0PQVBnSm9k0SNGFTwUGXqfR6Aa+sCCIRt3oigzXC
wX1ey/cMePEKpmSVpMac0/rle7yti6aJlcuzwKy2MGEn32SBg9AGWBqbAbnhlgHv
G58X7VawU1LhE2irWugch+5ZgR+nWA8eaNZ0jIXF28m3RPDDVbNe7GyYqthOZ0LV
A3DY/LQKbYvv+xtO71wuZ5RTGFnxRvNiZaVbXFbmpeyyT/Qtv4guKsCF2eaqm7TI
rAwMJgl2A825hWetayhEtcPcIhUEbup336rk4MGRpNObgRZmBN9bVEUeDAKSs0NF
TyYBQqRaqtLdcwRXGpsuY0qgdKo9tjJA0JD2JnyS6GXarE95oi2+EoTpy33fTiWr
kaNcDr0eLoB0yrehH3W3KLMUGyVwRKEEstI1WXCFbFRvRxJwrSsZexKtaNzDGAP1
Wny8gI+boD72ahLbyvCLmouMUnX3T+epFQl50PfJME65tRy5KP0Wq56UE62Ocaui
lThSTa/M+jl4n0W6Ohzu16Tv2O35tyJYOrjjbmtvrZePapQzgvWDUetxKtol+WRk
Vm2DNDoT4J8ahcKhmpLbDgGWPcZLPANd6eI2D4gu9R1dKwG/aV6KtrgqISdUmtZp
j6bQZHYu0gPGzXUhmMdk1ehwq/zJuy7ntXIxX8ilZb7554Sob+xpSE2gryQUTxiP
LjGFozBmCMdx4/HYUpgAhlW2M0CayLD3uvGYmEwen5JZFC0KwDWhl+ACoy96Id4g
qD90j9ubp+WFtM6CsWRVnQe7+ceR64PeprV2bwPNxfr0dEHj5qdFXo2LHoN2M9ps
Tw6QAYRH7Tt7LodlG6V9hMNlg1Vkh9wd+4fkpoqaltLJt9pAsb/MvCQbLJ6g2UfX
m9Tsostrh02g9I9wgLQPZNz1bp6lmWG+d8hhPkH7+5v2LzH2IaLAYDUQaMnV6VRe
zUxC5xsWCdFj1JbjJTLR0UkscLvxpoPphbxXHAD+joIZDuSnrW6OIvrw2jidEqUq
3h2E2p667ZvcQyl/GEAGg4q6Y46LlrzAvUHbf17NIM1kZfrHNs4vOir2VGIFRVCf
qbifMHdQVTX9oAdmlXTn6Chk5mOAGE9sn2XU4Ls82prYxwFX6plimGafJFl29s4t
j7amK8ppmVx5Cddp4tPg/SZRxWL2dgHEnSrcrwPisLdvuAK0HDHGzCZiiHYAtsip
DJmby5q42bDvYOpxFd+DqREQG/GaHJgdWkC98GtbXiFMUn9zMCDLkgSWWy4eUlgb
12BGrywUdK6gRv+MXPKsLjuXjhcXjvTa2MZKBp+w0zZaoDobi6wmyW6IglX1MIq2
AmHSvQ6Vmq4sxgOCdq787ACNrewUmzFurPTvxE5VJO+JJbg5MjO51XlRLLAV6IVf
xsNKmwskj8mUZexKu2sjNvA1MsGiN4oBSM05nFmIFyGZ6brN0rSpCc5cRXCgymom
gp32M/lq+sKzQtf9SITG2qXC6gdrCd4yaY5zTbQuGLxVbgoex3zQMmqQkHEmzbbd
kOtFuivp9dyaba/vo9XVkoSCe33A1HxAzpOzGMwvKzJXmNH7mbTevXQaKuRmoPAo
TX0Bv6vUnt5Cx956AgrqMZGCmyGQ/7TyeOrwadR7DgfZRc9jWSPHgxD3cDyR0emR
4X5SRa3Xjc3jD22uoqmDcuhIOJJhQSp0IAXh53WKUEDPm8BKcxs5wXSE9Pke2Q63
bKhL4ThhEOMoCdUeqdAgJn4WuyJUMxdbdGxLadOVO0oEn9NzQWLM9Q5i2lcLAt8V
7kl3FO1P53R2RrUKNWwY4IzC6TZ+ZPQRTxXBZmYdwbcLaU7Di4Fvg+44n7GJ4f8z
bPNfAN24IeyWffreLyMmLV4XEBSRabUALyFgFU2GB17kSk5RkGPvjZRQ7OS3zbaz
hdueCrjEHUhjwYq88X9EDAxYxSy9N47OXIqmH56YZ4nIdtzPA1RKbHI/VB+C2heC
c+jDMRVFWK9lf3+s11gRLNf5TV4Z8gFnbjrZkG7Mk8l7uNGZaGoKAKTbRxIBHp3E
XNzgLP9t0dX8CD74o958l68KTjBTtFjpsDC3sO8pJucAKgsbGEPISxazdV56n1UJ
MgqpLiW8lQiUWpqRCJkn8lvxrmpSvDT04i0ZkxSdhIGdoyOhHuHfSBiZv6mUI8Pr
y/MuVOMDizh2s9ucxxdx9HuC0Fl5b4yaaAROWewhrgYeIYuODNSeKCZqtQAUg3tO
rO5lH2dREFpy8yvwQZhoIDyOSBlcxcAFr1tDFFv9WraBWpFaQxDzeQwzK2bRXkze
AXeC2bxZOKQgCdyvTKY+fExjxKUQTWSyckxyTHb4OsLh+sg0wrl37rhSvD5DEov2
I7uXeznv/zxNfsMkGfaSzHn33t3ol4OJ+wDO0pTpFpBA14upPhd0nucyV60JsRcL
mp0RS2EBC4HporyUHd1v2SU1wcQIDyuRbzvwfdNCdbNlpgU5QgF14x0eLNLZyYzG
DwR1bWLjyQ1ydMpT4/hwe2XSephZ17OVU1jYydGxW1JxdYNzRwRtuPbftK+3T1qQ
Cac5ggczloD1EfOcJgqfvE+5uF9DtpLEODdSpcXWHhhcMsr+Ys1zuItzLv9UYBnp
WZEbgQgavIlNyNyXpTDnvitGiUkXZlbuTNmmNFH05AtBrk5C/bnPJ+In3a20GY19
KuzBdZEY4o6KY2pABPVY2Gpzse0JoyD+/TVxvaAUkVQAIGzGYc1muStdS8HwZ3mO
1yb816Do0YruFZK2YBXBYxvK0x0r1xa75ufKbTT4+GBKh2pZgsAhC8wK0UPtFJrZ
V/O7ViihewHYXz9xmd4MTN91MHZGcUNY4yIJZWMO3ghTBnYdbXeCD50VMXGQBLkg
ldHc0vg3DMtzKmKcZDD0H3aHb/9PoDpjU8fbDjYEUG4jLCNFFkyw1v8uS6n0VTUI
GUYmCCra3fQ3zxgkarH07uNY1pxYA+x/ou1SYi80SQnh654BPi6S5ihOIdZqAS0S
yy1DxZh09eF+iR8YypidlexkTyuMPjYM0RbkLMKRyR1V2lgIcB20NH451rjGcZF8
eFQa2OdhbFPWgpfvgr/3ZGlXAnt0VyvTQd51Vux2C0SkO91xXqGhoqAOkBbCWTE6
rD/cZ6KOWg9S1Z+aiupEuv/HphF7VkvX5k18t8HvLWG7EkzeoRRAgs7MxCR87/aH
vCgtOvh+1i2XVLrSqFT0yFL6ARyUAvdcF8sVQfE+zlmAPECIg+wJGLe2X98JeMEn
Oyz3kOUHP6uMMR7Gf7cG88VJc33J8pv40e03FH8LAWCDPYFf9ViuFtRbUmvz2nCE
0EFH0IBgI7ql5PwTPZZTZm/oVddnHrpHkZGOUmvP212vfZn+Pw7TfZe2SmsbyIic
zuLtrylTBdTsnO+OI2O9iC1CpSpk7gvIlIkFfLkYKMMW6bPNSZLAzhltPnr1sEn4
JxJ9SjVevAq3CskfNtHpHyeD70HR9sEd35DhiuVVDJePwSTxUGwTWm4CM9CE/kBM
vjW0nz8qUAQc0AtSLAMLGjTIKQ9P0HAgtZs/lfOa4MmwC86SFeV42eOQY+jgxUp/
iEvidzmrkTCxxThe3B/aNv/y5yddhBpfAnRIUbkdCrzolUT0EAb5ltxwnYIXKKEm
VTF3KP5lT+xGYHXUsS+nACB6xcCF5JMyMAooQmrZq01fEAvHaWGnQn4AznkOfqdu
VfBihib9LL400CiSIH+EoIWiS0TPQTeVp7k6YUrrytMEgtnG56hg/rWLfaFTaW0D
pn7sZI9N3fwdiSiVffyAzTVgPuPY65dd+j/S2yHw8mV7jSGgbBVqivtfVxjQj45a
flYJYgy3E+T7jW3/U+T1X4aDkpx4Y8Om+Txo4g5Qx+E=
`protect END_PROTECTED
