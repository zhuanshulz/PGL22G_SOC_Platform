`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YPVtZEEx0/2+Hj6keop+w207MnDKot4dVHb7xL2BWpdY/NxYGXRrNTQPpqNfLSMM
SikrwpKZ075ReIqZHIpR8FGZOzK4QvB9Xz2HNdJBcqzDRkcMNGsI7sanK1nuIxX3
Pp+AF44rXcwyZfzFHtfZOM01CkHn7j5sCxHTOMb4XL/ME6Yyu/pZ1zAShC9CNhcT
/YL5OAzDVEbq23xcY55DaxKIY0DpzGvxtjKcKVYYDjQccEEjJRYVP/0IGwd73WA7
F/ReQooC00/rPpYZtSnbTE7TvNLvxFl761uE/dyAB3i7CMc/LttNZ6BuNEYgOThY
ftPzHu3BwG3ijike2eoqcSYEPgCk1LXnjVt3G8jrVogxpO0btBERXzlztqhs6wTM
4zEIo43F+w6EnCV5I28XOGQel+BBpM/G6aMentQYSTMJT9Rjp1WwvH20W9bHI4gn
ePirftSRAeOyPzCuZqBLr/02j6bGBuM3esiSOj/4FF2Ox3NyWcqxZ9WT5318D/p5
XJpbKXF1LoG7D/SajK2KFF0LSjvvu9jrO/hEZPE7rgDmDWn6rHIHfJTZzWxAsCx/
tWZR8nm2quegRu2A+WKEPTSBvkDu/TYshvaKXwrugopmpMhbNfKmZl3tBQQFwfs6
k8UMB973OW3no5vw+PoEQWfEEiS2UCeqECMbVl72DFnFUPV9QfHVLl0DR7lBbUCu
YnE240QZ3IySR16oK7deycGOW5rpLuulvGTtuuI7l+kCu9nWnFTLW+816fZtsLrs
wNjKn9eG++EY3/JQGUdkvY+CcAplHYChLGKr3rYezvQtyLwASwOQN2Si2k7POMh4
H3FXScTdhUeDnURHHCKi6Oox/kO/oMKrkPlayKsNJpPVhAdAgqC8YVyDIjHybfG5
k5CUQn0dlgP/8ujrR+NDXAYVzXIPvmqJ43dO5FVyCEPp5rHP72vo8FDCB/hIltbb
dkWCypCvQOVG1SIpnTna9zFZ2nN8rRB4Z20qCq3sbD7KFWPGGjK2kw8pEbFTCB7X
vedyH6z5GkDFtK1/ah8A4ohPVpOqP5L+6glDNY2OTTG2IjIFlV94FWAEgOPuCXm+
HncpugmnPn7+Y91nwCv5n1bi1gvNnHBM1h4t0cV7NT0a1Eb0+tSAw6liQ7o5wws5
CnvBYdsjzqZIbWnv4M1hPi4THex9mwBIcGQbmzU1Lm7oNtvIYFvSqF90pwC0GV54
18RPPG4DG2tttCc9tp3dRBfdBQUwzwB+XIn71mMMwDcBT+0ZZ5ApnivJ5qeRm36+
Soq/j3fU1lhpBjxGpbYzYjAVFeFM7BT5NwStfcyQEss5JROtyAPlX/t+Y6+Xssk9
BOFqSjZMxWY9/uGBrOvke7+kXniGFbPEMpClJuTJW9EgA1awngHPbgDqVbXBp/jj
2A7Gm070IuQxSObUAKojN+nkYcgDJ2eg7qTwKHgKTf8XhCs8+FrXWJGr4YnGpEcI
V+LIrVVrRHcA34uVsnyvFtVKpoXR2fkSRN1gjnAVwK8LsnAMJRy/QpDdGl/zKgrt
oiixBP7+j2hf712rxAPjwQItqkpd9mWkN5vhhFHmX5ZgLjqKIHIBLiwBvcYyU134
1bbYyd/wEFff+c0utylUCTc4akzg6xf7ctYqSoWBnpA//Vxfn0c8q+cY4qZUg7Gn
DnuHHQwQ5h+WfE34XrLnFtB01BljOzYpjma4XDUTlqltfiPPohZRm1fmR7fOeZ0g
HNlWmfDlp7OzvZwa3NGCtJFtkJshxwNFKSNj/2Q0R+zr839h572NzDKK6r3mzMEG
IEpDLKMfnpJGuJKDM9bHwBor6e6Ft95tWSqvOhXcc0hcE8ppAirpnaZX/UkAIAzW
L9rZB1H0vVZZ2R76t8x00kuLba5zXwHBAU5LrlBYkx/DrNXaXApGvIqOXKvn1GD4
6zVgxcW7Qn96Rn/+L900RxanefZRvqkEJPFUiZ/fDOgVoNI1NuXqZJmtVCrirO0M
hqsT8mC8F6U46epiZTIEe1dYFRdvTcDiuKrcK5rY0BkKboQuf9VVEuygMHS8pSRV
hu2C2qJ9MqP4/OJXGE1tTQccVUw0xYWBv9RXkaKyLz9AQERQHLlFgETeVMsEEn02
OfY44Vn5wiFPdyljuyEugEI7dGA4aLVXBTmrTXMrkCERCWcaMK0Kc1mWDoc19yo3
d4aRceGrUjTuxHqCt49M2DeoTCT37S7cb+2k67kWyni4ekCvZ0bAQqDTwPZXP+Wg
7yI12h/AEPKpnDIs8LorjjFFEejd83oRNatte1DjfEqDU91PEAz72O5M3XyN9D2y
e07nGfhfQ+1nHqtBogv68erfpK04rCr2j1a4EqAeErltSFuHGCLHYyqXV/wHSv1t
qub5tiRF3ENhePa3czJqfEpIsDuX13L5Tbnt/htOYbC9jdtFU6UaxAQW1TLyxP1L
hicNZtljXIlyJoYjw3lw6NiLNWvM4kgNI+hAPu6+O7+cTp107r2Llj+fjxpU+fAB
ltYKZrfmytXz+Rnu5+YcyAUJVmnpFEAY4E/6mUGkjyxLjwYBJ5fUOdCDUPibAiD9
EFBPtJnFrCa9TuiBiRyXcKHNz7OoWSsYe+TNipghucw6kiLoRfGMjX1J6ABJxioL
NvMqeHwrFWd8PI/B0WLSUHnuJ01qRoaTBrBGHifD6pA=
`protect END_PROTECTED
