`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZSzFzCUgpQVCn1Ei/AZaIHauLNclLFXp4fWHrhlbdK1J/SyQOYGe5xw6oQjBR+a8
yveHaLGx/HPaSrNSnlSh4ECZZwV74YFKfLSutEdbe10m2ocm/wdXu/6ykyWvIzyk
6Vz38LKnmPpOUCYp/Vqe2EzkdkiD5GQa1xgNo6EtVjIr0lzNA9HEKnuAxcpHUuOJ
H9o42WBvYwK9OK/3i6bMp9UopeiYDKxNQeoCek3/13T1uCyW8C13K6jCkgbZwiTS
yxzx/BXK9G/5r5UrbSfnpCC//a56CVGiZZYC+rxCggFmwnPryWrSV2KGciY4K4Un
2WNdFUq2ZhdUtzYB0NSUt/W4yv4TESxuBYK/aIAzEgZ4vvddKeIUOhCROAvZdwaz
0G2rIbgswQiuIPe6hNbE/Rp0+BWzJrK+nq1pWH+BAsx5kFOB7LL3YE8dFDDHhhIF
arJck3faEKNwGnsJRktcSJNO8zG7sbLsspCQClq1txD+xRh8waAMhcfO642sgIdD
IoJq6+AZTFX+uxHhdlQ2e5VZWTk0HMeUHjwTHnZ3UgkzTOaeiJmveu1WzUNA6WhO
Q7pO8C+Yip4Twa7DXjkkvlpX2bxLD+TiKMj/t7iETDoMJG2PhXNGJcoz6yGe0VXs
ISw3c8AcFxecLJIjmmqVdd92dn95EHQ9WWdV2bvLwgCj0o42JZ+S8PAmjuqBFZrM
tnaarjfTVBfnJuG3FFs7lw==
`protect END_PROTECTED
