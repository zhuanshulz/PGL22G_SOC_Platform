`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2rhNXUgy/6lFxv6quBCcsm+0+14LSv0muvR9BeK2XLK0RKGncxRz/dWCid/3ujdw
s10fJRWXESEeNdsW1rSDKRjlBZrzr0/Wp3M7hJjOYnjn61CKo0gONHqRsghqbJrU
Q/jvMZgBVilNOISR1oLH6t/kxFi6OCR7x7i9tueCI8RkcbiuCeJB65aZZMyE9HFd
kYDTIM36R6yfLZ4sc32SlM9bp0FHl+44KShL0jx+jVxsbqkRpTlH07BkYTtMwlpD
uhAgmI+1zvVt7D9MONs05gryN0vqaHKAVO/m8d7ZYjLYKS9c6F2USHlalO6D+pFS
Il4B2nYHgmqT/Z5s+eNhoese8jtykSWJsoECdh/TTagtJDwr4bUo1ksLCw9yj6oG
r90bJ1drxidH2zHDboHRT+W6RspD70P8WEHecO6O5pSFFtg2PedNhYz8kevenViz
4avgknzOiJ9XjbdryzZLl1RsX8TqW5lxG/2slxRP5+e86uqlGgrxB+lmn8x8Rubs
gUFFFOEXfQCXGRiayHLD402fYMZrwkTSngbx4NODI4GUfDUEdmt95rtCrV86pBXh
+Pak9TrMn+ATe4XKb7D17A==
`protect END_PROTECTED
