`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0yXHAm8me1hE45o23TxQ209n0qHYIrU5iriEHsfx2ecYOFaInP8GM7nBrDiZTrpE
N3WaofIwdF8JOUDwOho8ZsG4lOvU3jnFKyJAKFI0qM4ntQhjbf9wXGVcXw/DJRuW
nI2majMZigfvkhoNVqKCw+pmsfSAbZylmTxCjneEp5aJpvAGQsrv3uiiws4DQB2U
rGL8Av0o6nnOldD4cvOKhGPSZHP7mcAfumrbi+MuNQrIT1STn1PxF4kS9On+qwRQ
7sdR1pdgp+bwcnPAjNoS1UCvpff+J6c0XlP0od0FfihdbPg8EpMT8x2svUYLSL06
w2DKAWYk/9UslQDe9U9WNiem2ZyQtLzFoETMyxVzHIrEfcPRgXtCl3iPHOW/16Zn
HN7hfkp9E1gofMmoINqfLCG9U88UwyN4+jxJFkNcJZvcZ0gmMd5H71UdZyHUc0Ap
JaNl0vS7VXz14Bepw61BIrb1ARAbVhMbL8M67RdARvTaLNAU4Q8bMUc96eB4QW5W
xFg2aW50URCCRAV8g50btCbLtmyrtOM7WzU7xlmH0oNk2b9Gxi1cD4EJRKAhBNnQ
v/MtHe6wrzyRuTMC3itPkg==
`protect END_PROTECTED
