`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jcLCbaqvAlx2P1/w6tZwAKmF2WreYplpFzAqbiSXLRTptLU4JeYP10oPX4NuE1AD
w9lsBO9oGr0sd3ve8pRCRA7CwHQrUG2sqi79Y5htaR5+nUlL3xdU1uH+eENs5VEG
6Y47SZqwsgMmf0Q8NU3PmZcDTHMiG9qQCcCm1fX3aeiB/WN3HqpMubNou0l1RwBs
NicbiNd0Xm62Jdn74AgTv5/HSjGe4KaOJEQbeNNK0d6+zYdGMpr0nyF5QRBfOzND
vUOl98NfcpzIwNQy5aS7f3NWJlUhoKbor6poU2UA4amArtTPpGlijQ43u4qEUXhN
VkbmaD9yJ50fGWGW4/pSZfkGv6QWVt+QkZGeUeP+KeH+v6NL+aknXPrSwdtg3rVs
sZJDSKEHDY8vaJZIFlrl1/68TPHol6aVs5IST5U64vceUOfyW2Tob/00NZ0Jx+St
u9ffQqGP42DtD6+0MbyQxA==
`protect END_PROTECTED
