`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G8wzZanKcmSvf+86cbebq0WTsCx/ZpNV7e1+S6mkoHqAIlKVjhYr5BWhac6EwKLi
FEuUVDpw3rd6gEVmHVxpLkY08co7qwz7ZwFnvjd0dq66FZIJgGnyltNMR0c5rv8f
kJ7NLK93+BG/2aOin6IVPtDrswAYfE28RoikPiFs9kiAyGpwm02naLY8MbnQnZQd
wgKrAwXOYrWRUsLawDdIxtka4tqWhqGhuKKvLKCmCsiwTeUBI1Lbn0Y3/q33CMNX
rmuol2J8izxLatepPvGUB7CjJuLZ7s4gvhntJHQt3JHzLpBTacMeD39pJU0jviHC
UBu25XLs8tHmGZuQhJYjS0i6fjZyCp8XX+50Nm+1gS+KtTUhgqssYsLlit6TXJdG
iBtb0zVzgjDDBmDqRiLtcN7Mka/7uFIIehu8Zy6u6CCguuUaz4OLN0OlH7QhLaIc
IlK0jktlv6X1OQlfIqAr0x9/Ue4eVpPUTYm+Cp9mlYjoeXyHL6XTvrT+uI1ZlXR+
2kpI7vPo+lG0sSdSDsBLyOReNAcI1/W4rao1DB0Db6Y7awE98w4KA+dKgaKCK6Mg
vbTCSJa5Rj+mpPxOICGyEoi0LHNYc9LWjbnN7O7miKalGdui2+gnzllW27/w1umW
muavL+d5xUlToPs/2MU4cYO/GFaa2AwvL99TJ+d7xs0GP/ZYDBJJj4glYIJn+RHI
HfGUrE+q4Wb9gj9FsV6CVuZ7WStQ6pgN3FlBL0mXRabTw9L5sy1Uu/8dB1v4iQs4
xFBKCYskcx/ntLMb6QyL63ACedwBEEMpMSIO4N02OQSIknli+QQwxegE6qowDq8s
U9OnNaLY02rat4NqZvVTZ44qpdvdnTTnQ8zvjbSmmnIHGRzg17U8goUwd/NPN8UO
Ljso38m1AAo20qAmQpVDo6JAD1FYN/ybPI8GFlRqL+09dK8w6Sbw5u7310ovO67v
wpNX0xZoveDdOunCdmpk1E+rl/B4o5lGaeE+YYR8BN9Hpt2xkAP/EHgGk8Q/81TC
B1tigKllB8zmNaj4Xd8Z2OJzT2/48jxYbDu7xa6LE9umXssbLeGOQa1I9TmlemS8
OVpNW+IsITocerEyGzXMh8t/F20v1jfLOJW8DUZF4xJK4nAa4dFbDFroVVC4GBcb
cGGr35Yliz8W1l2ITdTAh1PnIwtGdWAQM9aD1aYiVWt+Ipnul0bWNsfNKGl5PhhI
jbbpFL9uQ34C6idWGXVo+Mo6kucZHuN/48ihbEa0QT/w8u4lutAdrHSfoHaBxn5k
os5selNARzGs5kXFyal0dFQDdHqOdbYEQ7hWRDZYl6f0PYUlNeBx0tfm5QI2xmDU
w3Uj8HVeN8RXI/yj0gmYtZtjmRbJzZh2PBy420ilmisCRe5S9qlo4LfRnQmFMTit
G7CAY8dbIlOppfVmAacRBX18djL1sT7WQChLVbLir8rdg+b83UFmRloGTh5DgMHt
IhEnun5UIubW6zgqdAmaa57pP6WWFsRlP4gYNMzNGOrCSmspI8PZRZnCbhDath0J
qY7+UgX03XaZdLzDh9RQNYAivw1BdSFpBuQNNyL2j6Sxy396OEnG8lKXf8cwVsZf
bXjnPyUQKV07XDPVEJIrIWH8RSnTRY0Ovt39qbG3pWetkgT3eNr1YDGOAs/mfTfe
MuvaBnpZSTJLJZx+RPjvVdQ+guJaCjAK02y1kkoMnHFpUT1KmzerblY2AkHtRVwK
1bjpEhgDmN929o+tbnmFHtFiQNYwWXOMKJaFKnOTTTKwUGaxS67l9WQ9BdeCcbj7
tYzAHAv+bEjKGe2S/5sOt75wA4lQ77VU0rAqzPwhb4xtUTh6hJ5whrChu3DRU/Gt
tZltzjnt3p6JtEK5lzgn7txOeXhgGdC5gQDbNIh/y2N27DU3BrOBy8FueZ2kSNEA
FoZCFk9jglMf4/lDv830r9FFzosYgTs98q7bRzh+0+74ZntZ1NHsPNkvXSt75A1a
8Z2gcVPir+s4t3gwmH14dqxUZQJeMAm2FtL1qt6BzQinWP0tW/mjbVio5pemdwAk
yGyx/y/pM3tOWNiidZ2LAu/jNuMOGXEhvm8kBwRTxi/5pBQxae3SIhbX7SFyEOiT
Rmnzw6fACVccXEqmi1hFZfjRaXjfJmlFr2lDKOZoQb73NRENs6lcNfrUF+hw9J6t
bYZtfhdbKtza0njDhsRmceOucoE5XxtltKMhLDhnW6r7CrkwdbSYUJvep2XRw8Co
S0vNT88I5j8I888np2WAij15T3X9ryFaHPh0TqDR+TNGtWlIqJgIAsozJc550FQD
+YsUwrzUmlR95MIpoLJLuDzgoOTjbg3sqc32sond6q0r9Qin0nGCy9lSxiKOZy/N
qFQ49IyP+diG8AQdPho/B9Px13xZMhHMG5X2LXPO9knRu/5O2LP2GaJHkT2+p2Mt
buiY+EDcu0t3sYlMwaH7JISIrXt/ubao9S/g3/+u64Jtw9L0gumjBc+lfoUrm0ic
FO6dYSy9rp9TIEYxaXBJ59dhe4d8z05JW+0/akUvUTVYjODJxMfqYvK+Ardx+ADz
SvelfjplH8vba/Bds2axl1ZKWYU4Z9n2ThbJfRKVjmXskhuL8/FKTsdB6EGjIJim
F81XInGWGpviLFIv46e4kPN7mr60L3IvEUI0KkgH6d6x8+gfPmFIxOEh8ve/PTNC
jugiv2Tvp8fxb8RWxJN9PyFnGrjLASeibiUpKL3JH/FCZm+ISlaLtlc9sfKA9r1E
PQrQgY4vb2lLMieCUjkDhv+mkRMZHIZQ+nOCLKt1dlV1Fd9pWejvRk/KHkLdKZIR
5NG6Kc8Cnk2ogdXXEP1pt5CNTDtooFrNVQVe36WPqlpU4IZ0UtfN3Vjt0hyCqUSH
L1BFS6ugA4uZTLRZdSSMDQePZanl8+dJnb6XqITtYswmni/S/w8r49dC9ASsfIkF
rmFE1PhD5lzGnOWcVfWetJiUJJdO6f2Ih1Qv5WT00ScxiHAdkoWQIY66WCG2lilS
MLKyVJsDHJFk62TrEfyguhAyMRg6zXAa9Qiy4wGzv556fcBGFXCaxu0z+jdGvp4H
nW0I0VJHvQrvZR2kaDbsNXPqFLlHD6idd8V9htOizO1IWWpOywPgtftFY/CE/V7+
3VMIHq+y6uLgdvWTg7NJCiEHBPqJ4CPefbgRtfbransm4fUY2EZ1819sqJarlGVD
Nd/gfVV7yOIGMeZav8Ozgq9MnAsDKonU0qi5n6TOmJ9nLcWimHhcfoHGdI3Dux2p
5eSmrkIWg9DOEVICiKl25V+XWxnE4k0A4wd45nwoIIlfLQ9KFGl2qYjlN+PTwG5j
jIMKVaVBdzUBQv1UVWK88NSbzsUjr8jZ9N3D1kRsgw365OyewOyhSRHuLDy2oQzz
eOISFl5xCptPhYvQ1ojK61P259zyDMLPIjdXFm/ou3ZF69+eDose5fSUMU4HBBw4
Gl120bpP+m+KGtsIriLeKLxOThHBKsnDpvxvQYkBZ8DuZ0D/X7LMM0lZrWzFEJ+1
RKO8cNMtcFaJuO0mNh3UKg/DX502yC7Z7Xl9vxFXOC+JtxESqVdQcQP2Cy7Ktr0h
fw+95dpAZlweVlnUMpip0cyadZ4OSz6ZRQ6ts6bOZkKLbTzi6aesnQUEDDqwYn1v
nYbl28dzjbuXc14sEWhupDVZNpVbsMf2vZIC6O4lP4hlFWHLVN+Yea4uebkzMQE2
vJS4Dethp3ePXcSWw2NoYYcJgWQ0PV12v0NpaWl7zToNk/xtIRcB9THRDJe6hkS+
zK6kGWwhbauPAfIQowgGS3VnmiNFvl15Cr0Pt5byG9/p3Dj3WNhIVWTHGOy+vUJM
3u2//xQHAuEwk/k7vmhukKOK0GgAcrvjeDcNQnk5ojRGexTpx/Aj0OMPHbYR2jmE
NcPjjLG+hgmAMG70qqAMlT6rRUzI5xi76c9hpLGz8xA6rxj7W/speMwPNkNjm/bE
nVxTdi00Kv51jil08PELrH0cWf/WtFauyN2SXb0MVhM+6zSx5ecaZv8fLQ99nsNR
gCoeizVtfTxZ9Z7rKyu457fuuPsQj0tXOUllOohc66ao/SS68RFAqu6cN6tS05V4
dl2Ha0Vq9wTTlmnn0j1TVyYj2kzvS0LzYEhtr2UpIOAqs0ZxzBnmEPg9oFK/zcNr
QY7nLxEXBYvD9dWPfuar0LnlxG5HKUrvjWUr5Kbc/CvnZpeOLPOT9LB0m2Cd/AAC
YotFdRPUfZODZIpLxyVQ9eM9dAf0QM8RCN71wGhjz5mFD4u++2g2csYJuhPW/pau
GM0PWl46o2XIyYDRMCEPcOFSzzCtfk96DpYmhhdAjCmP+CPCFigIN5vRdvAb3iz/
QkbrPrPjYrbTcTOeZ4WnZfnLS12d79eAkkH6cUKoBkuh1VteyAI+fKFBWluXpfSw
7bDfdZ8XhUix/zMFZgYGVHACzUkshE/3PQ3tg0It6A4PJn0dkZz99XxBNBx73AVP
H443kZSOZVAKot/MxIzTkkOnnvw6X0QiavC4S5z/6HADLa7EVLNgtw7t0MSuS4KO
e4qKcmWEuAruPb8XkMGp0Wgqrz4oLR4WfhaPS/GxRZGGuva+atoq8rOZ/42oNHbl
QxkqPuM8veHnMwS9M+m0WKBCHH4DqHrltx11BEGkxY9IpzscAeeEAOVmV05Qa6YZ
0QznsnspQShDuYUzoyo/faU1z31XKU/obeCHmAdAc7kJsj4Su1hidK/OODb//rSG
k88K/FON+2LasvtVcek26jwBN6ck0ODj786yN+Qbrg0EIa3tLtkEaG1TL45wpVm3
lD5jHoRG2a5wGA9g6IIx4Al7VtHdvSExlXnHcVlo20yrPsrNFWsBvhR5e0fLTtzL
ounPmhS5l4j4/SuYroBa9tQ1Ckt4afmfKFj4Z/kr9diw5vIrx+odz3ZlsFjwMzOV
K9T0t+ElpffveZkTyFma4u6SZwmBJtUbYheGcRBKoX8cINtmBotNw9NMrcb+GXBd
AQCvcsFj9WtDO+VOwQ+hoivISxB3Za30qk97dt3gcBO+NniyBxL9qR/w8tTp6b2r
E9uGqR9LqcnduGAxD/GUgQRiyUFzF5u8SREQ+J8Q9bUDk5O2dJz6tfgyvUDQ/Cte
AMDBuafSgqbzaQiYT1fQJRhRgcPK/AJIzPkhuK8Ajk6LstoX7M0xBG+mkU+LCOfh
Vqqh9h6zWHbyTDM0NcYDSBGurRMIblU9gapFUJqhmq7XliMbpUYtiZ1AYujNvQRr
GLwfhp8K5ugQ0X3ntogNVadYni8JH/QACbFVgy87z+nkxaFV4FL54W2OYGm5Wr34
lJ0APiq9/DLqnBCEhZM4zRPe9AFGtJ3KQJIQesr54ErRN/RfRSR3WI8pyRTdiK0f
4LbVMMc8wglJICiw4LJINQJrutY3H9DMrKAhtqhLs5tnTCJ+Nbe7mmNGlX7pqFj1
/wylGsRiUihD0oH/1ix9gG+AJ3owTneh9lesfquGogz4U7X92ykvVnf22Lsj5aus
m6s1Og6Zs2QbrvMSJwG6mqKllGNo4qQjXenkHDYlZKWfZ9/wClUYlyOGEDtLmNZ4
Di/dm1HTyzEK6c4KLnmLbykWKRlIV3PtG+UrZzmmrzTIdHwNJ6MaBregqlOHqqyM
50L94fLdB2uANlghuAq89ZQh29czWJw1HeL5vxeXj2kvQFo64YFNoPzoC6K0jVSM
G1J0BPk3+HQWBSp8/OqiX475XmRwQZ2mcAkl8EmYj543jkMasUisKWisnW4rDQWO
w9aSdCCquT39dKu2L7BFCOY+L/v+65eASNf75sXbBo7kwhbBxjCQK9JDEVDpIdNZ
05iyUM8C8709okWbiIAKzy/CAdtxNC3btyoyVIaQ7DtQe0F8L+CKLssZuBKBlL3y
0KCg9o068ijsutVm1Y/Ej7SFhr+cmxqNWnKobBFcLHCrnCLW0TmJDQxlrvOpZ/So
Ip8mYvKFhk/rOuZqF/+JQVfFeFsc/oP0ERWs2jXEgM/5969N8JORixVdK4OMfYQP
W6neqkJDE/yDbGLg4zacK9K3oHr49UfFnR5H37tzA/sDCjItduzcY17PYFnhdyeg
Nzo4t4xk/1CXJv1a0J8fVVWGQlE/n38MyJP+n9m1v8jdgayNt25lgZlhyJSfuzAo
d6xDIXMonJXjy2ei8YJKwzUxSRxfCa25cfhJn/kDDDx8VJq2Zh8IT4aCxwAIhgEP
hsEwpjyL9ulBvlBWMXZGsqflujNwum1YR5e0Cy5h86AFCtxeMBgs5fiHk1CxFJOC
V6OqdYS1VhN0XtO+bsl+eYgALfukv+FT41a43uzW7U7JPdh3IlM8RCK0L8OA2MTz
eTiLs4Tb3LB2c3lC5sTcnOooZ4ofxiZ8DHcO9Y7euX/BGvLSO4oOkdEmGzg6gxV4
rNtdvpJZGY7I/3IwmU10sz0qUM7Jdt3iG+UZOJEboAv6tEC9yUKKZvlEsAfFlyJd
tXEuEVv3Au9th7Q3CJ4HaICRQH7MyFtYQi4uRKN3GiSfFFwOftdbnLSUAmGEmtQu
Quhyk8bgY+8+eP6FKsdi2FSp+LHoa3amKkNCVH/HKLVHejmLfsGtMU88E4NIe5qP
BpSN3oyYld2IDybdzHfvDIUA9Heem9Xw7bSLNr9EGRCOIzsbGQb9FMhQqc5T2ast
z7wWQMeUKHrqkauCPj7Nt/09xlI81HJIcTjEdLdZwPbfhuwYDmv0GsA9BGX+dLXg
y+dU4Y5ACCvrN2nCALDrLQYD5/I9to9Ze0M/LXBZDYyoOoaEwC03Xj8xqLUoJWbK
9tugwjTa3OtSd49AdyRvadrMKNXKgCpltTpRXPRQ8Ms8TYX+JSjO8JhEKb5X2wnq
KGeBTADG772HOxEhfeXkp/Oo8ag9jGPtTdIb25kkd06Dg4657/bVa+1Rev6Th43U
8dZXApWyed9nUK9vco9MNrlxOMusQ9kmsv0Mp1skgL+ZGfl5w/8agitTc47pNHXE
VnBvKLFNuzmzcJRWrQAs5zaj9pyA9Ami0OYD7U60wnUEtRKhIiIz1ydtbr1UsyGd
RrGX/jqm1TbnXyVEvtbzkj1dLB0lUvy5DBtYt11dLXOTXqOqKmlMX6m6Uo6P0Fzt
uLDPLZqlDrwH3WDPbu4uEi7pROn55XKrEiqola7SQ5xqIaeUGTi08h/iqhtvm7bi
XD8bs5tRDT8n51y2FmP3gCnp9ECz5p/LILzhngVjHkNbuRf3BaVxui6uq2Ryu1GX
LDnps5iftNkqOoXn/nOyeZ+Yb7/hXFf9LDKWmN1vpV5Hi3H6+DXqmw2coao9vSa7
3Z8ZERvknKJDRsltPgUWnZ2WrkCFgLsqqj70HWwJFgLbkYyqKbBF9QfS6eTkYmpa
PELF/uvslcG72qtXmZUfzNFxNbsgkIwVsjhQPcnGRAxjLIL+QmiiizgafxB6eqs/
k2HSjtu0zJ/BBfnYLJVEqUkjmQZS4SiEXVYBLJD7cg2mRkPWh4AI21fCsBi952qA
o6R+fDYLqOvnYPTPBn/VEIbJWfac4qJqD5IDHVzs5aMIesUoAdt6T/92c7qMU2tR
5KCEe7LANUGGeLhKFtJ9Tq59U6Vkh/T1RoVM4dQkvckxIy+qk0ddqIYVdW/gIVsx
KBzrECdN6uQz8OPouUy1KdswhPD0mK4DoQvPwyhv5JFi4d7JkkG0RhU+AlixH9CW
ETSKiRbLgVRV0/QcRURjLZlf1F6Ii+/AhnXhLU0cy3WqV36L+jnPBY2wOc9237xR
3XC064h82k3SvUlwj3N85BQYO9W3go3vcYFNzGo49jesyH8ofhtlyW28ddNYVW2n
wvQIePtToHh0ChuRh+A3vHod1A8cCuO2q3pCUZeVRdI/Q55qRwXqy+staulWBuAH
5M4iZvYHIc3M39fzjWwKX1gcr9Q+pvMuWdKKfKZfDFq39fYcqgv5emO/pJjzmDmh
q4UX6OWyuwU5guGOIJIDL1Lue85u7moEKnCGhs/aYe8Jzcq9yIdFNQuAsJ+TnFWZ
TkqWsFdxr+0KJrLIkXmb6LeQrj1/1tlV5Iuub/qwYIEwCKUXg7tRmnBwd0p3l75M
671gYSfhXdayZogpPOeP1G2Z5mHyjUBDRF8M1M2oe8ojozrNmTbfAWtzLd75WoFQ
5KqHs0qdMn59HBWGIzoOsSxnKuFduSwHvllTcW3eYJM4yT8qyF2OXOoh6R0/dapA
mbvqHLgy5/WDMENh6ceBSO5U9625ftMaOUYKZj7miQK6vj5ZeTXMI7gpTVsGJmDv
ZEY/PkBIt15NFYhinI+JyHJ99WiP5XWvkfAK9sa30aAUmJs9lYvY89PhMtQNwxh5
SLmJQ7Z8J3O8IW+F3fNtFujVoORei7sEGt7vzEXHv5Vu68vjjFB+vyd6lHf9SwQR
rvrzXWeW8W4umGk4VJZPmdAeiiLdYmEmhHo3p5MYz5uJtlr7VRwBSfKzWVKqGrnx
BpV3ScF3qRcq5TP1CTUT8b6HBPfSzuisO5FJrs23IL2Hapjx8KscKsR2FKHaIHX0
XLbmAoETyL3QrBELeeQKnz15DB+OFMA1e3gH5wqBsQ/+4zusrRc183gu+u3Fj7wF
6q6/78P/ywZW7yr3L5kGuaMKsS8TT2NDLMbP3xUN6lFEGEIERuohBmyc+lKb2pBb
pI/YVErWlj2POtXkkU3wsj8etNxoC2UoUGyWtD4gtWN8dr4AEp2uH5WI6cNquaPW
w1gQfCUdl2bOMA/Z/sxPPceoUB30K9nVOfVl8m9ekdQXuvJCUdD5mmFiXyWnV1Mn
J1SayCgwn9zl5tPShnA5vj0Rq6RtBwqYrPkRZBUrhFA/SHoVIzBSDzR7UM9RVlef
7JNxs39Yhe4OV1y+E6/MtsMmG63Hv+eZnUS6XS5WKeyjCwjdi7Sd1WWDTuEUGD1l
8xuWAET+dDvItft2FGVaS/mkb2Ij+xXyq4kGXAiK0Tyu8HgWQ3PTe62oI7rwTfXw
GrumaekZF/MLAcERaVoWnLCJZD8mAbHb+tR3bt1SbA+DA9YTFaPpBnMA55odQJqG
4TO4gHETPXKquBOlD1ksoORa0TeQdNIwH5FZ8rtSWFSSzXGDyVgqpkbLwEheS8jk
50Kdivc/l6xX0wt71ybmoy/IAim4hHyurao5KpSpF10Fv/YIY3JE3N/UE5ahsJxi
nOIN0j3WpWVCHJjqEo3REazDoJsXdOiU09p0BAIZJQC3oJKBLEM1GNUha+1tWoKI
lVRy05n0u0o4wGtv2gie0E3JAjem8Yt+FRU90wdlqPbbbhLQz3UcvvMuueueTa9C
3WNDHU8WXNNnRiCTmQI680y/dafFs88GPzoVCXQ8Sxqv8RZUIHHX9hTZ3+pcCAPH
lb6+kWR3rv3jaFcJPbdbsSdQiF70CGBGSNvXZyScw4gXuE+mOu8uqr1K9R2li5fk
tsDJ2RL4Opyf9eizhPoYS44XUQgdKrbcDnYH0/PlVIxQCg7ZWs+gGQaXdAnBcriy
9CJVeyWtjRKMQ7OReGKpsYYodWC24CbOXl7u48hWlKb977CtJ32UTBV/9BX0WILf
FTRucmgQqdgoNKNxtf9KSMbAm8WzVmsaATHjL69nRR7wOXyEtN92B306fmB8O+/+
WdamnoOinQjKVIRBy0at/ZmCB6ac54F1nlJuN+/xPDojIUhkYor3KU7otLSmj/Jy
6WOw3nE+fhsWeswEn+wTMpPAdHpCQ3Hm27Yo6SvJkLFEfCq1GCIzR5OApsZgtAqr
DmJmq/rNjTS96VTh6xcBrqJ4Ab4Dk8Pif3m+WroEtRN5MFP509CfFfUbvOtDIzkC
XtU/nJzHXQGvCIKuVT5AQTlMqeb/O4SJaoKcXHJ9srlsTtEfPVFQwPQqCTH2jvT2
ZN5809CVQn1gfrDpRhVrvXvql57RnwjwuhAINsPUDM1iHckEWsMghwn9fzXDLVT9
Cin9M4/Ls0Y8lBludownx2rDMEGdz2UDtIDF0SIfgwOzrYAoE3XB81jKf65YkPgU
CeIQkcR4oW+8jSWxXztuDtDjnsmqjvABseKU7/yxkk8ypK7vJZgvSIwxMoKNhJo7
+7fpA5TjMnxgOrU774Y3vkz4pTFpwJizZgx+hEnbYkgqjfPFSJHirepI998Wzmau
bpXIkWpzKulE5cggsh8x9Q0PKBIL2hLducLTNlZAu4UaA9X7B0Tu2ayQ2OGJD6jD
DqQp9eQYK6dIO9x84FjBv2JbHFKP1Irst649WewPg8dfdHScZXo+BUUkt1dipolQ
dU+dFacHmMsBOoJAxr2QaS+cTpoPCRvvtGJaLuhyIVWvuW8YCl+ilusA2Aw9aRBK
ZGc3tTrNHVY1L/AxiDrCvQKM4rSizuNSUizPmgegdmsdf3hhb7c9npQ1Lc/P/0Fv
4eHnX8zRUu2eEpzt8S/MZiwPzvLPb/fB2EjeKE9nrujvLNv1gca2hNyTz01Mw6a4
IVKbH9TblXXsLo+xbNiF6t9zleJ13nGD9+6IeVpCT/+R7t+HaG4FC5AUDCbPzo7g
pFfeE8D8gMGDdtYkK+G1ZVLFRz0s6hobzuxb9DQIX3RkHiJxOD51UCAB1fFWdrv+
jytLXjscRqY2gSV0sMIvK4WO0utIr7ye9FMphv32F8OzAm6Ny0QrGKtsjx19088m
7YG5BD2sBBdB518WNHndzHDLwJP7JIk5ArQPqfoboNXUZM3nYJCCcwewixcEA/ap
ObH7PIZyqdgEUPVn7BqHsgIru3+lDjoXgp5RAwNa6JNo2S99LksWwWV/eoswWnHm
y+r3Uy8YTnLPG0LTb1KnLLROYNzsP/h1hEH4fg3nRXEia3FiVIJ2zTElagFGEJrn
TUB/sMcoXLCvO1aXAiYQwch8kdz7I00FLgf8GN6crmKXvg0Cj+w2wPVhD4z/lhqG
3IpEHac07L7GXlg1rUjtLlSeN7BgpX5znec1VDqE8JTctv2BM5iqyB70IZEUwIfw
9DZggxzxc1sY4wbVD7qmzrtgEFLO4froeJSIXK0pevflBVJXswFFLggY5QN0f89j
NjSOcSQgo5rip38gYQ0NzchOgD/JdpEryxRPpji+Vz/RBhBdh9Hbzxxkn59RnheF
AaWpHMUDnsncyo739I9uCbs5p4NGX/8SoAtvg5WrpKZdeb3M2dmgoYgNoF07nCRu
TQGz4me4lAms7T0xxmfObahEByDWQwpp9TxKA0Ua7EbhjP4CWAyNCYr2vBADFvS9
aQjG3qZh++EmQGZmIiV+5sAKG6tAMzA1ZosLIOUgx98GZOLSikjFdt5Y7pLnQZ29
MQSB5jsQIauI9KetB/oi2WYcDCcZ694qYlHyhQezBrU9dcuqyyn8K+21gA8um7mt
kWXP+HEocMI0pM/QPNZ52HAH8JOsSMJONnpMdZa4/7y8LaZ7xElg7hQZCZMIqLHr
pkbr1gQN2jhoDxyTKWRrvjbRILw7wvWzY+yHZiJ2dA7zjqv80nnjKD4l3NuY/Qur
dNTdup8rXhKB2skWIGHA+M6x7gHxEMwvLR4UeBPngVmXI4boNoD79lANpUTBKOoF
DE4izjTVNMJY7MRXKZk9zs+Izt+qbR3/XfpUMnyIuG/SZFC1xH6Ae4YlEBvp5dUQ
7yUOfnyg++t28vIH5Dfo9DDOFsPwGIYP4lUrn8zdrTD5v7o0CrZLX1Up2nQ7kO05
OoPbjXHvf/Gm3qDpdi45fgRWSYqSt9ydjMwpXV4f4NXLv5cjgG2V9x3lV4D+zH5+
1U8kO6UL0zdU3t2xx7VX+ReY9QMCbR4xM27ZI5nLWGT7FMmItECRQASV6ho5Ss/T
KMsyS91kfHXKj89rwMZBLz0Nr2Vbvb0Y1J0veNafQF+Wi4ESecnZMJDmW1yXOPv1
fXvdFIN8LOMn763leSi54HPGoakqMdMlaYDOZipW5Yo8hfFsAyLR/bCPd0iCw45b
n716n34n6d/zzwzVRJ/yBGYHwRQlesMv5nEO9Oa1yhTfvWBNXXAT05oIskjDmypD
+s7e53Gf81l9brd5IyTaKkfphhY+OuGuswC5+YM3wRL8uNeY1VS2uoob49l7hRZa
RYy0KJy4zKKcFJTbgAK2kDVzIpkwHpX9qX7O68q/Uet4Oucv/BDPbGOrVbOZfa04
wzGm+36s/9SQT3tOp7qoOGgp+r+FRlyhMjg3oU0sDyZ8yZt6u1Gkn3easQPhO3Sl
kfqOl5FHBM2QfmwQX01ZAq7RrHrU6alUeP3g38C5+SIYzSiTNdluE+aUKby36mPy
LXUF3cR4/5hIf8f2Qb6dsXQZzyhSpZvP9Jr/x8ObZJ1qt+aunKOWtHnvKG3Ub8Pp
tTbAE+s81Sa2yFvWPtDCQnrK0zgIH36h1JxOy9pNS04EvVzTam2b7b5j1aNjTlFc
kj7/XI3/LrSxPHpQrOGO7Y3RnvC5UwJv0YnLoipCN1EISkFP3PTFNXpqY0j5Bo8n
+QfmtVZOyCWPM3fvapBbb3EK1eTBatx5Mojzs2zLgHwLdifueHqwcV5YKR67SCJR
07oA+i0YH1g17+yImlLK7XvffKb3lM5hFs78s7H4I5gINXY14AKaUnMe5oLbBYRo
f4V7nTWUIHRre/h0gu9BBfwbkskh9l8ISaCAK3ltnW4Sg4Sbn1KnIAnQh9f5E9JK
i+vXxAt/rBDzVdmJgD0a0dh2gf7Ghf6YrUiKB6xWX2rsoxyP4Lt+AHspoZLfAs+F
NHbnwZBaWe/U6AdrkRCJWmKHKv7w23y/RqULrqx4SuCfkohS5kiqxFM/a7ZS3De2
49rJQrVhJOdDe59u9tasYNlNS270uW/AJ3EdMUzoSATNMapifIFlOzhX5MMIc+YI
C/4n4jiiiBmO3INqz3zOQsJX231n5ZT0HUCFPw2k44WkEhMS7g7YpFczb5AK65mq
1oAMTd4ZN04ou7Ub6gu7sJ3HpmPeElIEsmJ21xXo/w1BG7lugYbvI2NCZo6aSXSL
A+Bgu870tGAPhTyAKzsxIFGJlyGRL6vbmQr4WXgOdBthFqC1LTdUKe2CUT/DrUc5
rfsAobx+H5JkzN66W6f+wXcWTDNchseyplwT6TxO1N8GhOH1c5gpszkD+YZt3Y+D
pFNegkL2hq6rV6d8xKc/LyZzKJe/up5Kz9jkmOXOR6peWxuHPJRsGDy1APeIQQOz
Y9ccMh4WF71h2KC0dAhva7Y+qkczJzMI/Wlx9FDd3kQ7dx7G8AEgAZ85+qa+H1jj
XT7bHJYqqTuYS+DB57EtyraJtdJZMkBYNmI0Qlyb3INbrx9Z9+X/do2j3ZUkuRd8
UmCDMgI6k2TbcXrng5Es70Rau36zkpnv9JRl1fOnh8z43j9csNoiASWT6QOBwq86
xSjOy0U86E4IqgJI/3DX73atfmArRhsba4htP8wj/vl7MQkxkc/FfzIKg/V6J4sN
bcsEvRQPClb1PIKroHG4VlIgYnOVdyc7MsFHRedSwEU=
`protect END_PROTECTED
