`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ery5OQaeFZOwHIEoQuG7yvzJ78EOoJppgs6QlE/rRWjuGrKgkqabNvZG7niliXdm
jVwgjmDLqjDp033EILcrsp/4Bf8JJySiHOFHQZf113noN0NK9vWy+VsckOZF2BSn
Qxj0Rkyj4YlazPa8l1A1K9YoTy0ZVEwK/f/kAmMJoGOfaM96Jl8xmDNeqMp4WCb7
+roBQ2imKmWuCLs8OFI3myTAmKUNfuaHuFfPMZP7Cwu8QWc4SIfk4cMdhFinckrd
Uebs37oSTt8VSdc18tYgduyrWRrxIEP3XYi4YAs4Mlk5B4PSXLhW9fsSrHorbBug
`protect END_PROTECTED
