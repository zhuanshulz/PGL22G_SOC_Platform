`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fBQTAAkyEUxeILfLZveFmM0MxV8Q2kkUY0bDM2q95fXOo3vbDlj9XeU9SsefgYXs
KGAPV06oB+vMUaW5HvFeY0Tt+IC9zw4PMkwW9uCsdRK6Q4E4l2Lp76MQSNFv9zhN
C0EdQoxRFJqilsjWJHS9H3cHgyY4VnGLka5hklqXEdyZLQMWgsqTK2SSAYRzRdxw
02gknQMexvK86mJw2l8+UnR1xFMsF+q5yvtPShuR9eA9AIfQ6g5WNRhmOiGy96v5
Yo0RruiG9eVkqPdZ909vsFlhf7Z0YM5JkjmzJJK1vG0X5UvmYvUw5AiC/BiQrd4I
j5bmvRXJJ3A/rDUylOpw1A0S9Igs7QTY4Ng9KZe2ZEdj1CvAtFQTsW//fPg8vbTn
2r5/SRBFzL0Y0pGHTRmWDwwmb+tAeR8/WlHLyHOlmly+iVeh6+Z9RAIF+UcFFXmD
9ZHXBKO5eLoBI7ltvE0yiLkjfQpDInRC/EwcP9SwM5Z+2VbeH7Q3XmRgHw19Vsj8
3EADksNnivV2hsteWu4s/n+Vx9O/VV9gygeTVhPW5YNQQIedG9R9aQ1vkzaD2d3P
/d50Xw6HpRXPRXBKZst0HfcdJ24lzIS9qs7iD0buH7c+Ra/sc67qH4tNM9X1drm1
cSXkq4x9VF4rhX7tHfOUrAOsLd0MTSzP5UJCrjJiB2C+ERhleXpLNu+DmSG9Jt0e
jWt9+3n7pddupCgwxRRxXQ==
`protect END_PROTECTED
