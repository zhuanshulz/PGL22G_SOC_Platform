`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TXjkDZum6McP91II6i5gLwpb1PDbep2O4+3wmdmcO9jQfEN0t6NSWqACRBcOPCPg
gkhnJDzK5kMhjgr4sNG1cW8XAvHErbBlHh+b+GExUrrSwa/2q8YBxMV2XyNi9pvw
3CQK+wlPLsQmXV14W9yM6WuwwuF89V0nwOOVZfTWxP75vHp1IvIXy2BQCCyW2e9w
wjkrtos5IFadQEPjWuktR85BogyjK/vakHjvi6aYNrC+dPwz6AC+6ATCm0V9ksYm
HEzcM4p09GrBrltpuifwQ8759JoMMjvnSUFtgVmxBD1m4rxcFY0P/pXS6pfJGT0b
0YIvlcKDzKxI/aKEjL7K1/KVyR9ZEgo6A//f+El9PmSuadSkTPUs5s0RmqW82LgW
+4I6alLtWIiPq9L1WtgedRjQr/j6U9WvTwZuLYP/GKfkMXORQEgWMycZeLoxmm5f
ncolnrnvz1izsmS/A7euqutrO2dZdLEvrMGmbhFwuRpFZTDYgNNdhhOWneAUisFU
bSPJaiwyic3jqAAI3Ekhf8i9Fv1Y97o9rY0PgBzKJfvhii8qX9AxUl1NwGi3n5H1
VPPQKyaqELh8/MLLZhsrjcyDfwt9N71/pI77V4Kctyk=
`protect END_PROTECTED
