`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/Pb787z+QG1LjvcwU98TLtacaEjCuR/dHAiLbrsIq1OovYvtm4tjDQZeXyeeqdgd
6NgZs9StaQ6hyjKHukfQ1CqcQD9WgZGEIJNp+DRkXl8pBiWg7IuK6Dyok8WH7o1C
dJcRhScyTwv64M88OnJM4rXQj8XXKuknOnAb3QQnm2YcbEIFsj+knD/5TZ5ERyJ2
skhUOJuhB9DqGC8U2oqZ6o+iJXlSCK1UhoGb5LrwuYVc9+RSNk9YSj/heb01VDt1
zC+mq1oBs1kQkLDa2XschnjCjUnGmrYFE+WDJ5dQUKpAkQXPRTdQ2HoUFD9A39NP
HuL3/GGSxAdPV4OJ+TiBblkitMBivj9u8f7e2RuwE0MvprQcyETrCpLYm10gfB/v
/oIMaPi+9kk6VQJN1MrzO8zzjjishU+LZkW5F3na/1fYJTKQErizS8Par2l1eOCH
fT4Mlik9cn/l1j1fxBHcPBY6n8kEfC5ZA3fxof6nd1kQ8LXM2wlHcrcRnK/kgDTI
jhNIg3oXQ1/pwKn6Uguo+D2bsK69MuaLot3OPE5qSCginQvvlYv/r1+aKRODCSDo
DmdS0Y5d5IdDwo1LpoDBxzw+5CuF0YODh8YWvmoUF3zTcoPD3qiJl5nIBkfcPXDb
WTjyiJ+1dUzlN4ak9MtjfCCdJudxMUKFslOhVcOGDanBRIJ6HR9GVPMrrEfsa+le
z765NZFOQqa9/CFn8vpZsxuFMmw+ql0QV5m8aEtHqYm33PnlBrrVh7PaGD2yM3Q/
lFsva1a+Tj+2VMwX3MfVBY3WjhpGCudvS9E0NpB7eab6ikbVvzbL89oFvvNuOX8g
tvRxs8bDEVH3RtfItFSdZc65Zg5YrPZSLR/juxhMly/ym1YKB6VGY9aMoJaBwbHJ
no2fln2xfgc2s1qDtcCIOaJ8KMv/Z7dHHaNGApt84N1sPGAMBN6JLNAcJM0eVHo8
YASyXlARDclG8d0dSLCaCt9mVPIrwuN9lrKCg298iRs=
`protect END_PROTECTED
