`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BdI8uQ+uSABp6oU2aaVPC4C4kK8+s2DcV78dvS9x8HQ5etqFG+vFqo3lbcsYvgGw
UpCLBms+1+4M016PdjUmxeIjjON6b34RZkscEIb0JXHzykMseLk6Y6hStYSReJJO
1w5QYzwv8BO9uDPZ1sBgnPmwCQEa+i4gJtrCFeTYnp9THQdvm4IqHvATlU66jOei
RlPC+8VEUQrnnSOmzecsgFx6aMmTFOPIgX0ELt1JoVqZTLWjo8fg44CetI4Y8AQd
TmsoZK2as1XiLJii4tbY+FvLeSgSqClXcTiXXRgUxCK7/wvD1qsPQ11Xv4WoiRSL
A1TJYqHpmIn/uUhTPXzd07TM2MUBzY2CYd1CyABFVRMJFEhUAYENTajXjgdzThsP
/BKPVIqZJfYMvCBY+hR+ANBf3+drmvkGpQNwFaYULodTvBo6A/j5vHMxPVPn8t2+
xXvG4GAWrMPEtsfkXvzxxQlxgIeqho0LfW62Auz0fL03JclXuPMNTyZUZ62/15+G
BPxdCzxOVKlG/c8V7kqsutYDKYl95zT7uND8d4O1GvaOGm/U5EWaRoKaR7OqbkhZ
ygF3aK+LBBeso/f/b84Dr6s8eV3Qm9PeX6qTtMRyJSea27pYaZssm2lqv4PnGjLt
PDkVK55CM1g3XvMQT6EemPU18jeQ+9BpFIfwQ9hz+IAc8/x47dcMRT5AwUi6voDG
dYu+T/GDIr22pj7iAOOUx1bs8ItPC4cF2PAG5fefoEYZBFC4/rRBP+BX0CkxTH/n
vN0ilzyVD0US21J3i3j+l8d5cVpZZfM+VtNbnIsSTVNWzUSZB9YEhcvl1a3Z3Dyo
`protect END_PROTECTED
