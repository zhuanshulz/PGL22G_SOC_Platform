`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u/Yfm4nYf/Oytv1G1+eB02TmFyLq1zeySCnbbqXMtpbTbnlXx6ETifexi/WydmS1
8WVPpobSKCpZ/E+zZCt8dsPznXXjl1cbWtGp8rdAbOFCv8lijPy42OlD9MpiA9OW
YceB8Z0rEilgClJjmQvCvYm9bGd+v0rxW1iFkWbg4I/WzITT6fXxl1afpK8O3lMP
iu3lY1p2TTfymwBzXinxw+rDUYpUYUN0KdIkwwF2cYFTK61Vd20xT8PX4lLp9YLT
aQN+qNVlxx/7Uvn/BLmDvqjbH92M8EZDqTkhwZfI4xoQ2L0sTArGyhmbqPIHx1MI
Qt0ZufxNQhkaf2rd8gh0UzEist/Yyu86hQRToFBADd13jEd7cp/yhMDsoB7+DdB9
fZ0aTtQ0jvUFbtOgnnMsQzMNPcZRO7iV15/z+djL2MYRYm4GdQuX5OvvfbfnoK+n
wYkJDg1HCxjl3bk3caFCeeZxThoMNV4D272ZZZB+cbcfK/FgN+PXCla2HdSWKgDZ
NxaHdXgxepWmim2ZEAye++Fl++3tYqHnAXpY8qqbGSxd+XaCWGlhddt7OfTqRUmL
DmziaoIhKKS8iZglq8i/7ZjqqZ2xp4cT6RocpmphDuLrgfCWGibIskXb+LAdGOTB
z2iFz6m/nKObptLJmXULfSpa1Vb3zM1e+iP779um5PTMP1ZcvxfZIeYLnO6s5ASr
2S2opa2JQgHkORiRuC+8AekJAOLE16H6TDdMlAKg5eiUvh0S1AyoMtcauClIN0QL
efWd4NO3iDf8xJ3d/2TXfv1UbvmWsX+Akbj/WrbdrRkilfGgTpmiQJfEyFIxlOWw
lR/qZ32VV4IXxuG+yWKQwp3YqS+qqAxxXOXBQ4DTWTXTdJNWm+LNxpUc+F3+AleS
boztOqGbQ/gDAhvdS63uxW5UmBcinXevHcH+9e10OJakwKBo1lbuxMgnE7MFjIRh
IlEJgj8NuqccIALKILEAXiRLkLoaVSpRgkTbVgXo7NcmxstiM3L6pef6jetc/CBe
HuTx5Li8SDUYulaJjL3odzq82fKA7fkjpxFHuZxMSCG8MEMN1UqVNeq/2T8htRJA
nZm7gG2x5uCP0ipz1Q4PyBqdbVwTr9A36lCtNsWwXmOxAsKM1wO+lrMSFks0meRz
qUpfTZnzxZHJV/bQAEYXTA8QED+IYXuZL0/3l93+FaNsgVsd5LQRtPbmtz9jxtPu
euTL+PlhB9AUGgquPSheee5wc85zD8zZtwlXbgzlTNCf1992HkUrHOUVInFxmm8n
BOn9D+RNddtinKfjjw+V526hlt8Ow44SX2LhzuLrjsjU0wtH59wtZbpfgmEVoEQQ
V4zkkbFby/CSZWPRU9Ug8T7BndzFOty/D5SEeBz3z7Q9DbVK2eQQEoFCY8UlREff
ZxHQsR5LXtZ01YlF5GbBG8/Qj0d0qoDMFziiO80WlON5oxIeljgPRkI2Q0SakZWq
UkCz0Hfxk3XwnE/ZeYrGo/4SiWkthi39g1Dp7i0c63czedjdcQKesQwuyBdvBW4Q
4L3pJe4dqTqXBO2k7m/vQSPeL9NE2TK3wWYO8XjWUs/uZ7nNA0awYL9MJsWMd22e
UE4PcMi9ByjbqSBPCFsFyWIW/nZ+Qi1ZzTcVRoZ6XrficOkHja79bVoP6udj7VJp
XTAAefFaEsjpzy54H+vQZhh7q+uDKl82fibmEO+hxulmxltpeOdIftTB2QX/DPz9
xd2T9EMeV20N2MnczJCQhNggpCngkhfRDmwwUwcXwdxKNLrifGwiF35+9LtxHfw5
/A2dtxnVfLo6NQwcQE+9dLah61SfEI8uvAHW0RQHgaMnuhMbuKSu8qkZyLGB8qps
hpw6sSI/KsuM1qK/3Ndklx4zCsu5vVYqAtwhMpcLBZ1xV6KWB8UbcYHHW1RJKyfE
V+nq4USs9ky93NLLLewJVSQRRUaB/dwQbTl9XpIoEmHg6EqZCU7HG5OYk+7Gp+Iw
4/vA4Yv5iBJdqEGAvoOb7TM32+i1QWqe3sFyytl3jHpZEFvIj5NnRC1VuMHAdrfW
daCupT3ZItyVj3yXw8IsD9p+hANxwPWQ+E+ISsyz8uzSMN09P6Umx5aMZgBON420
fdfAl/FTQkiAu4iMpSiuCwLQSnUyMmm6C4lhLUPygIsrAgaI16kcw4rHZFULDjfJ
ZLyH91PNZaHNdjfIpAhTiyDTMS3zCrJPz4PlNO1HznJ9tnB2kxU71Ris9DoI2+do
+J1dvju9Vy9/J1+0MtmygkDxfJR12oVFpiazIFYbssRqqvfpz59E3wcVzoUlnwQ3
Ehl/QqQbU3fMPrW3VtPeMqkn5O3cYukRECwckndYce9j+n2u/x9p163JcidPj+yh
5xROVYoM3hlEtSCcH9j5v6Xo58SCwJkgj8U7QKMZnDEZADBDCz/K5pveyDsxWBUb
6U3hymrvLQq+fGL5SqJm+NTIa4NImXDCTWiX/OUqTdNJ4KdjaMFbcta1BkwdD6kz
7M6p8OERdBV5WcSddRvUgd7vhuVF/EHV69qyUnSwKs1GRawGA+dtOFzdxLLRTVzO
MwikmHaBH6jMVrPDpUBNog44IYvw6VGdZqm270FmY1tWN69tcrw+5zdjXqCxoLoN
2emW2OiNB998ffTxGnu6fjbVjviO0vIMUmwqnKg5rV2fu9VumEjFRs4k9P1SUYpU
XqPBZazm6nxkl6O+uu7jH4UZp+NkrYxg+TChbM8CY80xT3JHml7HTIv64cmnpxMN
TI+kEGqNSGclQMf7BLAvRg==
`protect END_PROTECTED
