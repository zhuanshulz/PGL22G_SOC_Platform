`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EVyJ9Aio0cnnHdfmCuyNsMblOViWJEUmwpzhb28sryD6ibX/qe/eLVJDiCIaDqug
/lSiqkKna6iU1oI/d8cghIaV+9EMBZaWV0hlUzpHsuV2nBsfuNCIh411V5THaGLu
p4/BrsPCJLFyfxEROPfwistwI5Bqx4EfLGe9fp/vDJaocydGBoPhvNcGwLV52W9N
IqcXoJpaG59RhDjirSUDBDrUBrrErhAuRHG1fBXe5IgHp7UyrKtR05RB5xnbtgYO
d5auhMgNY+VTtXID2MeUTT1mjClHKGpIgs5mvWZVJ6VKJ+UsGwQJDqjotMdCPT9a
JRB+YMUN1vw2B3wukQy8xXt0Qh73Y3SLahFTjqZ1XoVlQDskz4YWGtqLOm4IqFmT
BMGgz6KmdVCIdeKAEy6fmm9EPj31h1WvT1aJbBjO6kjw9KSlNAAWx6n2RdOebMaH
38EKxrmpiQfaGOqrS+l96DlgQcYMzX7fvku9Ovpi1z80sG4PGJzTusnWx/jwla79
6gR8cXgtHbvw+YrGC6ipidPkYYn77Z/lutcp9zMn60r9fBNAIHiLDNehrICAWTr6
YZoVrwYTLQ1G8iszAmMYEM7tCLgvn8ctNsnR2vmHk58=
`protect END_PROTECTED
