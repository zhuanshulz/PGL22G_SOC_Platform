`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5+aLdaPNxT+PklQKr2bsedVJkHGJYoRIaKBxEsz2qktlfLvektGownJLuTPMG2jJ
zCV+7NT4XTPLYjqdlKCCf/awPlGLihC9nByB8da6U4DPF9LC7kU9IlSMF3RpgQf0
Jzuk41h/wFK39tlwHCxSaXkm+ORJPstbDM1LeIJ/PXJ1XtWFFvWIGxu3nNqkBred
/Bc8SWTXKmqlHSAcWu6/vDW/R+xLnjjvhK40POgi/4UBDWXA+82Xgjp2qNlHVmCd
Ju8ZkJjv5Qoqyh63UEdLLyapRC3sPHAnzMKmH4hd0M5kpAf3FIDjvzDVtNH8+WRP
GN/h6jdmJ8bzaof5VIaYGFVEBPeI5G8gD6N7Mp/fHnyeR+TV4Mt2A7fJWsUI4cSC
bY2H9fZ0YCkJqiK+8YHLLEfolEA+GAqPiYGTE9qNTMDKRXoSQIex3OKE+URSZqaf
GzLWPekmHTMVgt+NrRtYnwFS+U7amJV4KYQaG4s5EkuwiU85dFmhnu3Wpri0m22C
OSB9X9Bc59GyED1QcDQO0H1U6aTqoQ97V2K+ag3VTU6yNGo+N+BC9YHAntPT2tpB
jCePu2E4yPrCnC0F5Pjvs91tovkThmvYv4a6bNAVx5DsVePLSNeByWQ2TsDGpOkg
tJG3Wq8TpyX8pT92ACa08S1prXOqZefuui7os18L7O50eDmxWc0ToC5bqoujMIjr
KZNTRELhU6gvgv+RprlNyk9k05tb7MpEHRhcO/pYPLJWEa4Vb1+0/M9LheVUOuoP
UX5cpLykEPcuc7DHmwraBj1reKmp2TfYj8nFKV7Z9QzvrtDe2i7+u+Z6Ff7yozOw
KOAaSvk45/IiaQfGWUEXNjA6UE5VKeXKNZqWcflve4FI0P60MLDnf5nECwug7QnP
nzVpUtNhSum55+cuw7oTAkEQk5buAL3xdfRQBgRThuECwZY2G4A4qSEl4xyLet62
ogIhXE8CceRfRhXNPB9sWfoch5jT0BgEFVKuhUCmRpU4OL7uw+KKLCB7sjeJLlmx
sZ1DGbd9Lp+hJx+bTd1XtABetChC/kcsixGPrP2HLwO/riv345/Etv5PuaoADcio
Br8HCDzkHyfXUm0UCGzkQAy80/f09eGo4tpOi5GVyqQYG8g86RvLI7oSP4AY1nKX
4j4AOAqbd468eHl43W0reZgfV/VHpN1pspHVhi9Js07DbQVc1JX1q0Exi1n5JgRB
+7s7SldlcgHofVvuxMIyeE5GUIRK0rFDQW/OVGT68bVwvtqA1OAlkGGn+g71RBvQ
IhjPfmBWogGwa/KkE5gm/uh6Pcdh3n5e/ihoEO02z6nlMsG8sGC9d0T3AeYErP89
CaV2hOVy3/wxatGwjLXgEVpWjVhCo+kiaS/O4XxvSEnANwhg5RFGK3vvoHX6Ze2F
bKc5aoHOJWCPou1k8et9hDM54iHK4odPfXhzprc3L3ZO32RrtgKcaY6hIc97FOs1
/wvq3xrrKWqVNYu0JP/QF2Hr602/cfOvMTA2xSYL54n1cXj0Wk2K4+O/6V/46LQF
JIXWObmE5StAydBcI0nl0tEpCJF2P9pKzQ8i6Wqst7o1PIPaghNzbUxQQOzzXKDo
TPCzJ2u5CxhKLqO+eA0VVieWanyqytPIzA2adTqfpTP1hw3DepouyDljii+JaUIo
JXZP+mNqlwXIT8JsHzvQkIHSoVS40soLHi4oRr7k295KJBVcXQbdO/oJ3RxmQ6Su
oqcuhZgluIBiNCRVBFY30+PFpe61aUDony5NQnyMBlCtD0uU3y5j+CpVUpWN0A34
sSbwbX5xW4mM3VZUyC8HrT3VF202xUSpWXsEBFjRDT6aopT5ncdYhFZOqfkGPI2a
y/Rtk5GzvRWKZmW8HV8+vs+W/xWXx8tpjgB1Z91npDexbrSHdZ/bxp3h5OKeUVD9
Yqwoi9gs32v4LEO6fPrKget1rmL3iUQwlHYmKJL65k6uydRjZNb8xy38njVvYG+x
kdqD8GGOB1krOTPiovfQ/CVuGAWx5+XY5K0OSyGVDpl80VdPV7J0Mdasx+dpkw6h
w5R0PEtZXnB+XJ9JmfG/l1SghpXI2aWSkpFhEZGO7Wx+EB0puNO3JsF+xsOFXRnO
XeX4k1gsVieCFDD9XSoJS7z4jrtRxTi6SB7YHZ2XePTTVq0bl4U6Qs/7PTs2K0lK
vRStDg3O+yK2SJSGhr/JONJCmZkWxRUDPFHZL7v6XaJXKn84abI7lpCCrwhj/DBQ
9Tbb78e1fPi1gu7idGy3Ys2ELGZj6pDqwlKvDq2UyeCb0RXd7z2eJ4GEI3nBX+SG
bVsfq7vLbNUAV2+eWzy5AaE1+LjxXRDwIRJhmkZJF1ZkgeEMxMfNAXSnyMq0MkZR
`protect END_PROTECTED
