`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JM6HVTGDLJOvAsrD56DImh0a3MwxYJuoND9MCb1KQujh3s88/R54wLCIVY7uCSjR
/pdAPj3G64j6Dsq4+mWbPY9RTUEbicyPLoT09b4w4+eQwbJAE1SnIKioX2nAnjw1
qtPc8wtad0Tug9/h/PrhPXWQGdI8AHMGyusN+oPuWPmc8UlCIIIR6F0bzjmKh81g
Gsnhyu2hR3d0tfNbYSLo7pu25dIbdSVj1qzvJUwEpm5kuZO5ZEh3S1RaRHVDL9xy
ICRp3cNTRdZ1X2WBaxbz3qa21JYJZkovqJovl7zHER9NxlK35Fqk7ClbPLKnNQNd
uSTG/e/PS/q/+HLO5qLQLGCzA1+It1cNmx3xLv4Sj2s=
`protect END_PROTECTED
