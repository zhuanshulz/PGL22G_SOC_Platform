`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rI0XZ61IUdjASkoeMxJwbMe3fF6N+kDYz425FEMHqoISJShIi4PbUR0/KOzg9DUn
uDtmvg8hlk6aMGgK3NUgJ0b/pucygU0S4dGxYqSanKlfm1WU4gqfWSQb086Z59SW
hHBWw6ogxBLGJ6M/MAmgFH/FglZwiUbsyn3xgK4EQGdACRDLjWCjjjOxcWHFEvpn
LNiAS1ACHF/wYmA2w/r/6lrr43lybGQvC/W+5/v0azmcKHjbeBnVeBlKSLHgiXp5
3UfQVtcM5AeleUMvGWV3+hR2I0fEX+AlE+H56jx/yOO6LyUEwGV53mwTGDqqzJed
c9FP0RD5CDwiwoThIRahQnqXUrWoZrq+z+X/YXdBytL8E3rmR/0tBA3xBHYHR7Ds
oqh/SlDNmrJgEKZJwJlgtj6guBv2n/KZ/Jso0RlSJ/CvOhYdX6LWmIKOEuC3I01H
bzn7hk9r+wzXrbiHXytmRhKZGcI7GET1sewHpnpFoNWobZF8wM8mjPdrlBgmt5JF
5YwDlZ8I6O+KtIu4mJAb7b5mX8DUxichNoTfPOWUMI4=
`protect END_PROTECTED
