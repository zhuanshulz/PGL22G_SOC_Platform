`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rSCYXvgOgxQ0+w1ZehZcajuWC5e5EtV9lRBHuUB1XGhhdZ0vAFY68S0ePZ3o4k1H
5Jv9HC1pH20Jd6dI6dV49uvk2yH97lRbf89dYP1Svq580g5wLhIvttYVPECbiDXi
YnyzHDnv/a33ZEAurl1GYW5jhCwzbKtVJIL2HZ/D9SpQDJNMdUsZTEldhmGviKHi
xuU4l/6875tXwFLQzPy59YoyaG1p+QI3S8rKw8lbpqJcu/E4rfdDpzsFac4Q/lz+
7QXXww0b2AbUDFz8jqWablbifP5LQwfmfGOBywdo/mLpxXlrISDAKYJhKKyZTIXk
l5pSqdokKdViAcQsZxGYmqnnXtXuCoYCF3GdKD4ZlGKOYUtPJzw7iXactHq0jo3N
YtFA0P69SnMCjJMVKm9E0hDfFmW5Y/nLnfz2n0M+T58dtB8FMWZQzJB4K7sTs1Of
0g1dvoHdm2EatFt6nt2PPlN/B4FbeRTsfZxc8M0Bu93JXqvCRfYBcI3viaY49uox
LaEjyM27uqkHO/R/eh8rzrphstnP811EdqOHVq4oLKeIPBdaxFt7kMUOeXVkO2Vj
MnUCFDjLIqQ6hVN3QV7PsYZUw049czqoPn1Hp1GysSZKECI3IRbryx8kT5QF+SqG
uAMYI8ZYksNiKd6dz9T9NRPpmCAzxxgaH9M0KKbA3sQJZTJ70JRnzJbw2i9WbCei
HvbAQlloBMae4mF+wI5envqdiIbAIpu8AX0fIUZXgLTMNDzPY+AbvMwGqvWrDe1B
+vqESc6uIsizJ6LBUHCQgrNz7rZjxXa4LEbaOqwbb5e8qbxKbxSW1zNQb9flhuee
+Qh7oOfpkHWkg2aPAK5zfhGfoxWSKUMRfHEQ5I76p1iRgQ+ITolDJhdCilzJt3cR
FUbrVnb1pqS06Dki6BITMU7oQtItCDxFK+T2s9tmISpDE+9XhDXzJZk8eO4rbeAJ
FG+QXAuDbWeQwejHzxwFxaf4MS/3kyrY4pAHxCDhWGRzcu7ty5KASGPQyZ86D2Ex
lrnbZ3+dflNBDLaLCHLN1g/a5JuvWqDrKB8x+R7WoGBz6PimQ7m2UiX/mZxHP9wi
U0bodV0Lq8SlCFuaE9FkdkTwsA5QiYAJFxJy3/38CZ8UV9HSoIvoL5h9pU1Egn05
7SkuxmngvbeiaVRgQ1ysTDsSeph+JFkUEWbUUVVW09QsD652BMqsv5j4rVdmK6vn
pr8C3fx8WM71VIOuJ6XfrB2ENsHiiDptwf2ucZQVJX1pD6wEArcY31jI9lLzAxCY
7pMzrghNhTZ3cbkC3ErGz9QEvr6uZjup8MPAr7nm3pjWSWxkErrOjwO/78wTwLsZ
1woECoR8ytztET23cz03KLeKaOgcdWyeJMAgdc8d6sa16SZAxGovJIWAmbkJnP0w
WeDHL7TBCW2ItYFbWMLvS4AKhYoO3ZVDMA36SEJA3jJw67nZm2S4M9kx1rTJv3Sd
a5kkKr0ErCo5cUzvxNSZm7APxHVo83vFt6iPuYuKEsjQY7OvHXBsfoiXs5EN8heh
`protect END_PROTECTED
