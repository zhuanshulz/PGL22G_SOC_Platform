`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SrIDCta248Db9bz0AkTdGrH+1eC/aW5VXj329n4nyvU7jDAL06EkJmrfzlq/ZH64
ySJUEkdo10rguYmZ35vWeXdJxPHuljDI7VIXLltEeMVsEzzDHiUtOHta0DvpNxDX
o+Ki2oiM3tm0K407mXvzBfHLhnSaqflILVXf9v2vCvDUErrOrbNXUsoq0KDf3Ugp
mylgGafvkyf0eZziHODzhtwuYpbEC5WVwIniwgGuD04z0sfNjJUrUzMDER+ILBcr
x7vKyF9u1OEW7WGBSjB+xo7wLepL7vUNOv4Ff6y8WIO0jSC/wVlRaY7WCzdfNZT2
7k3hVfE6IBQxQS4mfObPdt3GJMyBf6xvV2mp2gcgjKW1gqprbKW1BAY50kHWmRov
d3NTo98Vx/Swprcgs0/8i9pqFTdoqfax7QQgTPWMsY8DLHp7AvCSdOfN+fuRObbo
/dVrbYW3nBiBIR4Wt7iqt1UBE77JC8HxJQshDvlHd3nsPg7U4DDj2Gx8kIUZVtg1
ptrUhvsA6QdByjZJkAZxKA==
`protect END_PROTECTED
