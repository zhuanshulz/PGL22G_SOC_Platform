`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/hDZvWtFBsPaNECIj0TXzkqGCKH4I3FhzAM0dhNM3DgU+nYupjK4YiFOAoe1Q5TJ
a7eoR7dPKybBEdk5fbM+hHU0WdEps4Q1yKWldYqyQCAZz/7ghghV+0Brv0WGcX7p
S8cFj6uIThjNuww+vW9wNLMnLEhz2/DzupToCkzo0L+akglu1+Suym5R4uItIgg9
CX432RVMYFCvbuVt0Q3m9QlV3jkIsot+ng/C8GJy8TmepS5RxaqbyQxThsZfpyvX
kM+/et+6Kh0f3d1v8p9Zyccbmyr9NanIPTwoHoWFYdefFZJqIzuOamrwfk0LARTy
Xk6OBl9VjQIYncwMwUupjgGEOWCrvHNWkDzGbgC1XkKGoj/ENvOpwTRWdXPBqz7Z
81r3aVSyK2RW8/Vv3zOvsojnFtxlEHUsI23e64OSNGjIijin3LaQjlB7pV4MXsnW
TVljDqhjB4HZ5HP/Oh/MBLNYrABB/9b41hOLQ6/Xh1aIXmJBh9byYf3b2SDXNewb
TXBVePvZgzIjRA33B/PZfA==
`protect END_PROTECTED
