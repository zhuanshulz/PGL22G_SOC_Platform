`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EV42f1ZnL11cC6uiMbOYurpOiwqb5RJ7YFDkLIMxC0ODEYNRSC58/QxhdQd7Kwgk
26LB+VZxwrpD3tpex/ZpCntYeYL80iZeyQXT1utq9LlTxul9vA+oq2LhkMKE4jEG
0FRv+gFLn/FXtFroGmevYske3MC2dlsfMrQh5tGWq2Hx2qrhE5LmwhhOsX4elG3o
LyVWLAou4KC+wrhRheTNZtLakVM0z5zimewJ4hOAp8KoDsYmJWprywbCsG8kbJxw
EKZ3fgDRBbJiyfTFx/epdm8ICmbM9uGAkysR2rqGn6v/Xl84S1DGnC8ixkW3lEQj
Oiz5Iv+hG9RC6wfQb+CcAw==
`protect END_PROTECTED
