`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2F47QZnUnTFNHjIGraC1hJ/54pE2VokMHDwfOCGljSq5OKrRKvpnptJEvWkzm6+n
Almsx2KsY6XctxLXibEz1U6H6LOt3iGxtxmG09TauJ/ztnyH/kU6g09R+Ohh5Kou
xA28KjYlp1UBi9XcuPyBN+CV39zURZLB8QvvEgkqKoBAhpKCUUgRFx2+hCp3IWop
LEzwDDgjD4pQT9CWj3GOXPAKKsPtUOIBJ5jgLlKd1HUVmBe5GY5g/Ofx+eRbefoE
Fp3RnHF52MBchTWRqTogcDYeGa0Y48BWcnOYtgef9xtMHtxGM8581dr3PINW6YUm
xGZOMkAN4oxICanuipTDqg==
`protect END_PROTECTED
