`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4F2G/jn5enoke/bCMfYiVz3v9Mkms0XT9ZDJb/tEfmwFoz8b92yWrskMZ399MRF5
/WiACuvyc1JgFbmx4+ULZ9cDpdXXqBPM7vKkgX6X27wENbGYjWqQs1JjIMrHeQ7g
Y/ZxRlj3u3tE+SNDLbdXZpzAbeVvAhCCr9vjHyywfxXS9U5R7XGfcjQCEQVzgo7P
vS2JHx+Sp4mDbKoIma26ZGQZlc4PN3TyYuInFKl78rXp2nfGDXq8FoTjEpHWZEtP
rq7XxhHUh3l3oFdcxw0aNDfKi2Avy6hmS9anzfJAgKjW4XSV9bESx34Gc0hb0LG7
2PK8rtxiZKfqxc/yS01jM+UWZ1FsYmyt9CFXmVJFx5LXftbqEE9S1CLiQVsCNdpp
vVpk/qkDwuhOMagcVxAXhqDANC3xtETPr/YMiOc9zDNZ51sxeZ3rIQiZodGgQmQT
TcF/CLzgyT0vZFAYqSbs+6Oc0u1lojn0GU1Dnu9l6jLH1D1x1APxmIBHQfCYE13J
m184RcYx4IYL6j53ngLrnDomQLJV0BHU8xSf3/NkWRofW0HU7PdH5ktu1GjCdG3C
wEVpgNmukXNJNDDWy+aPoHG8YsqOaDlwvCMDF1RKLLaUIqdaB5NOLmfJ0u6iEYY8
Wg1AsnVHGdub9JojYuJ6x5TievYHcheueZ+z/A9qMN0V5k/WCq/tfIMOglf0QSde
xP7bRgOWIWSOkIvgv9NLzIs6flJhOXPNAY8xDHNLxik/PHdIEBHoTGl0sZv50J+f
Qp0mK5q3OccmUffbbsMGLhCTguV50NXeIDEsKjrZjvVuUrQ1x5rXCJrXp2vEk2tL
RpCQIH2O3EQuga/Ohs6O0XFLhilXiHpHjum/av8DmlXyNe78gFo1U3rJGu00734J
RF6qoi6e8jVyHYPmhpuATsEbJfkszPanP/59Rxd+7SYd0V51hE9h4q029ombBCZz
PFFksFUec1OGvaiLeNoOL2u8A0VUcjb1Lx/BQB5oGVUrmH+v7Ixvv8PNeNc1yMb8
8y9WzsKbJSrgzko3y/th6VeKERP2aGFtuEnvQgkMGXyfzEXeKFDfPHP2mqVZoP4p
wZZIHuBfTlpwp7YBEUsRa7nf9ldy//UcUp+LUo4uYM/t8mDVamPTorIlYwUlZwST
mSOe3c878R+jxlWDYVQc1HZ27DP6De4N1ZGsOgacpfy6InbH+2fEgKLh12OvK2lD
jcl8SQVsVq9fgPdd/C7VP4naqXDLZxozHdgRJuifv4o00dxF9EEY+yK5mUoEbDRt
/XYAxFMoQsNzXiBXlqlqh0kdWBWwHncpD9a6z/TpPQjDHU1GdJtqfDyQOPR5QHRf
HJYcxRKsCSUBXo24oYUbo+Yawz8nnD7pBbVP4jDA0CVDyJEdWx/UXm6wy1hzUiET
mb57KK7C0/UrATHKfurW0bX6DZopY/KofqbvhsTxG4sXxsFboJUiMT3yi57auv1O
ZUdIYjxQz7yosPw6qcVktPv+FShnxgwdwiI7xY/8p7O7REwx+0fAiCiNMopHAURS
WHjM68xjVbXNwngSmsG2a4f4CnNyU+YbfFGJOcoLLy3naPAdpR1dIGlrdQ7n/2tv
1qHk/D/VfbN5/+5cMkSgLuiigyG/4Xo2+DqpRIt8yJLsM+jIzlqbwEfl0D7jRG+k
A4JPaf+/Tn+dbHrEBeGUO/iAYX8tsbaQ6fgibL83w6WZx8qoJAZApWK+zj+CuExu
9rW0jDX0NJwKjuD6lEIo9NHX8w4KzxumX7GfbgCoE+FEoiE+DlPt6UnMCcuCRXIj
BNW+3QsH8rjEWD0SxVJOJljS4mEpfYDeh7cVoVXhSfReDm37g4lO8U37iGoP3UGb
3m0zL+WUVqVDFfG1psns+kFlaL+r3xvWO4X9NuYLTNFUW6BArMXviNIJLJb66ZfP
EXROYjCD3tfjdLaY2GTtWQ==
`protect END_PROTECTED
