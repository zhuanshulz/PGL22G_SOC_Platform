`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qtTJ0ukPqtc93iGbQz7M1K7hXxnebooLSGKRQjhiDdoRKW51SVt3H773lA7HheXX
Xz7imhNwdgNeWSfM5aqpVRZoHb8ruGsKMlE0kZRYlcfMlARJGR87g08nB+Cs6xHI
rC97Uab1IA7CMKqdtxCvtW/ipRRXFDZ/zPtqtAfdrn84VP09UH3KMNUKqG2u4WnM
It86hWC1M1mmyxWba05od1WeTUn3iRH7cJFx7CM5QPOKra+1J0xhyLM8WpS5tR0S
JidU5SMfLhQa4sZipXtxmoYRNJg8/qG3ri2Uy/L8uSaIhYNe41kL6HSoKX77e3oB
hx7yXLAfMYYoYj3Xv9AMDeahhAhcJ6GmxVR0UQIj9UPCwDhVjJSdKf2J5VKQPCIt
MHBfi/NV/gJ1C3Mihb8tkjttIZk30j05F3xJsz22J5b1KsXELSF7o41peq+2vdTn
dRLLzIRvgMBBonyrjWh4UalfeZqOegFcNJ1GwssHERm/gfyQsrfktAWb4er9/qpj
tZkZy5kdN8mnRt0fwbYvPvqK0hOEKps8Oop4/QFBdT9+NdKItYrySsgtG4OqNA/9
GpaqNyyuC3XCswJTAWG30FS5wu9KQS5FIHvA4YoWSuQq7MCGQCBXu7DiZbpyjTLn
OBlHByVDdwRWCfO+0s2/SD2hQV0YjQVRzjHY9kOBUar4QyNrfSnxCRbsLTSRphfn
qovuc71AE6TIL+II+OfN9wbQRM1Xii+rIZ40KvDY/3quoDBbouBWUJfukJ3QGiEb
5uQKnRpAy4x+M2TIEgoUaHqxFBtLp7enyTWQ71owf0Vg0DAC2bkIUFASWA3SMqhF
V634GWIRIvnSQHWTAwLenwBUbKcpUWqRsRNVmNzdKV2vcXL72knI/Ti0fGXNiYVr
lgo5AIwZ75uMKNz4IBsR30QCev8K22/tPMhGK7CBCLnThkhg1tLtAfW0mrUIwBX8
9GaLbdQ3zt0pmyq1MExQLkEMhmeofn56ZjhZ+G7zUCBWYpAXS5zpan0zbxh36PSd
+ggOd638d8VQolWVZeQK0nhYNoXT+A9hhp3DznqVGZNjUNEMQPWlEGzaoJVllBgH
8ht/yor2tGH7Y7hvJlcCFrs8zOFj5a7yjVzoVlVMr88vMQVwFEW4ZA8tY0jYBRH1
lSN2mgJhTY7i7a7LcXOVO1UPZ/Z4xNPIalucj3pzvNKLNIL+5Lfm33Vm1CmnDW35
+DCQbMDItSKnfHA6sjLTJrET2afwPIoGn4DS+1wR0HyMkylYd5VTilkjDFEWU8tR
rDCZwYhCwq7ZlIZCjGt37gc5aQoAZ2S31V0m5EpTJ8lYv5sXGiQbmjTPsWOw91Ka
YxBvjtWVnKcGw/Jo/V93AxT2e4a1HtSzVNDIuBPS+RJzhI7+HkKLy7LrSJZHWxYG
w+Q6eCGpBMUOUuBsc3TgVw==
`protect END_PROTECTED
