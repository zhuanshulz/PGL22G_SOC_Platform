`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QhiNOii3msNuPuWN17XchlWWg/OwHVW3NhD7L8oOR6u/6eK6BafSgHz3R+Ruc/5B
l80CGCeaRNPwvnuBTFb+9dDan9pR+IhmBjSjElNqBN4kXKj6T+liEmJ/XHfrE83c
aFkFXhl16y/5bdQey3IAP3Ugz3e9wgS/sj9mBQ50O3HfpcuwOQLzFlDWTDuFOLUl
KwG0bs5pt0VFB0VPsrTR/61hZiv9yTMFs8iui4pWBoiD8los5DvL1m1B5Wq+aBOA
odC2fEO3l9KpF1x7coq5RoosNmQO+v5o9+BvrOW3/5Wi+vbqZiLtlzAKTUAkitWC
VE8gFK0sKS9wTbVzFB8BLdrs8zX7mqkFo7n9peDcQq77YCH0L7FU/BgEDBm7Gsiq
MlFsyRkzuVDAXEID10iyoQhMDX6xAOd5YqHWsXebFnLJTnrpAOkdNFVrRZsejDzb
VrBM9wnHHuzEeCnhUjfStRuVtg2wEL2Jg+BwO8X5Rrtla987QdK9HbXYCKXwJSS5
Pp/ZZxV6P+w/PhjEFd5EvT5pz5Z5UF52LFHoNmeRDi9Xg62VzvRm8RkkbAHygQz8
zZ12ajSA2QOHCHV5qzruFitDDkNw1Ln1WO5JhmaqVH82dL84HPfJ/A5SC52ZEGFo
lVhL6vTRNzmHNa8UYdUccw==
`protect END_PROTECTED
