`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0v5IAsuzT0bIwAlrIm7KN4/n0zWy1gp8Wq8+NAluC0p27BXbjPU3MmRYOtiXOVHL
Bh3rPqaqpEv8mdhIBkGTx6KLhzEi7rjQOgWvxAq9uj55Doyf1QHt2C2mY855lIir
wxS27/AuLaNUqhmcni8C5ZoGUFG2YqvrhLbBAbjTqrcVla902ZfUuslyE22Ny70N
Q79EIr0hNXIG7r+EIpgbPfnObOh2xwD3MS2DhhEOwQvrovRZPMDT57VnTO3KoIMR
rIOypHn4fCF7UqftSjrAZOH2Am6tLlg6X+iiqIuyKFv2rTsS1iMNs4R8pY41rsqi
cy/O3TEoftYa7cOVNTvdTmJ0nX8oWSvxtOQQfyu2LT2kPH+nDGi076LrmzyNZeN+
6QFW9TPZ/ESudhj7yqX2w1owWwHINpTYTARmj4i+kk4IBHqCkQykaoDwbeiiXBIx
zDg36IkQNn6Rqf4KKcqhPffOraqS2jX/riVeGxkRUEdVhFnvQAKzNyyWqiCHidY2
jyxBEebp9l9w4Ojvi4v5DYnR8wIWxJh05ZBNiiNhhrIvESiMoTT3mIwFVo6AmsEM
KSpP3ARl3umr9mG26ndG1zvF6zk8dQX0qykuidj6R2G+DkMdEPES6eF1hquqsVjh
dz9UG0ZOuSWVlebnDK0R3inO8B7v8m9FYYgj5cA1wq5Sk/AblV+U99Oui1wWDSOg
hgc3WChYRvUYqJxzD1ylBYGwbJ/jZg2/snBLJgOdrxtF61hgmEcHpPJSlJFhgIoB
rkdT77Q79a1OE7yjlkpS8H8LlPo3WeFql4QqcMZv5HI+6/w5J+XlWE+LRoX6Xv7m
ePw1CNS1Zoh7GPMtGwMPLdqrHZlHN/4UeEN9NHElBA07cUHPKYaxCQ80Q0TLiOhI
ImtqaN2Zn7N5Vk9TfglfFH4/oQSwllCj3oDxCI8kwaCr2nXY+FdnkbURqMR2mHat
q+7iqMD9uhFAP3zcI0AsrX6vzj0fSFP9gXlmKfzlVWM+EsH+IKNhkI0J0/ruhy6Y
EpN9cCARSaxYmCPnIDiICbn1iOOdU4VlfTtrpLTQzBJ2ZDsppNxV4XqUnMmIkRwC
CSgQHuD4DIo+uOeidgww31zosls2qBUHm6tHpGiIu8dUPIAgaLHG0e9JiSzBBUcl
bkTzOd5kBmFtk2cwi5gsqlvwnTpX3iI5rpOJuLfyLuo4E5tgCHZT3z5IXEaUTG8X
ie+whdm+wUE10bbLEQa3Ag3t/zfkbxNuz9lCXTs1LTh3M4v2Fjk71P+HepO/F4wC
FuBsM6uXdf2ggILRSadt3VJQ+UYq3OjabWmaAeBMmCP2109wUpw5MIZK4rFsNy1Z
YbL3WPKlrvKvb4hIxBEpblzwZBJvFirEsVcTuMdgsZo3j11801sCM3N/I255a5Yy
WBBLp7enfv6zMss7jKEyYE9CCuhdBdT/hxN21Ntn/p4LOWdwJeiYtgtlLVScGA/0
7GLck1TmNTmQ/oXLgL4xKc+Az/yQ74ZcdpSQxjnFTLoyEmAwWfq14p9p3yUV+OgR
FtubEBEQNQv+tH1uWal8/XU2rNlIc1gaBB9OrTDWhcF+SouceY+6crzvKLAc7njK
ptb+6isypDIUFBACSP5MyY3/CTedeFRa4t7Y9Bb2tQI=
`protect END_PROTECTED
