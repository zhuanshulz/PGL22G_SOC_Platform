`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X5LoWPbiUQ+oNynZ0hoKEYZwtKLnOv0+kdbm8eR9Km/frx4c8SiYgC7dJEagGeIm
vN1d/FmlrvgmOLshx/rW+S4KGH//sbbnYSeO4S1riC7yHc0WA8F4hzVl6snqpjV4
FAWlIBlAP/t9Ui3yJlf830b0YD/Kazl75eCLKT3c8Yyu/U/qDPpBuMMGJSBw4iE4
B9xJpwqEmTLw9OsLQIIe3SpZhT4bcYax5fuuk6XOQ2GJRRIsPWibr6N14az8mWMj
aajb5XMNhS2i0EGkq/CtGgNt8xhWEDG/ZTD2kmTJhviLMt3MqAM0ROtYU0RZs6RI
RLUxg/VkvDYHuYmpNJeWBuO1wp59XUDEWWfV/Ag+yyErV3hsjpCCgC/GQXMZjx7q
smviLlZNzMmR4V3BeO/M26UsWL5li/x9om+K8XYox0S4G+PU2o7xsa8cLLG43oSo
CRl5tMPbUU7GfeDwDafcMXKv2qICPo+YCR6213NtWyqlYPT0cVQnwNfApOpVsQqW
gWtpSBBaUOPKdhBLUkBkH5e1a/T9ieh3/AC+RT72meI=
`protect END_PROTECTED
