`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u4QWFUT7Vzrex00AmvleNaUzVaC3OWCgHsDMBOytnJoOET9CxXTVi7TdajggbP4F
/tTJjK1TWS9yhg2ejGiu4cZjhpgrtgqC4R6CHvpQ53o3dX66cuzGtP4KpTsssYaa
oWjNBhwD/LciTERDSjfx5vYrHIZJXgXjrOJxPHyP93F0qaAM8XRExxR9Qdq/y4rw
UmVStccilqT5PnjdIB+GPNbdRM4wO1jU/WUptk3GF6s+oKL6Gn++hFnwDjFZRJQB
Swp8Ph5EZgn9mw7ztbJH4CQRNpt4uyLNevM7mow3E1XeI6cQ16AnOFsYFnFx4b/Z
8mpZ8VcxBnYAzNfT0QPjwoEpWNHmH52d1hLSm8CGeLG0/IXMoz46ABuaZ40ojixl
NmOmGm/GlC0HiCoEHbU5MelnC0S4ibcwCObcQnYPWuaPi+T7FWfCYVBe1HSpe8IY
yPIEaikLGHy/SG44ko3OwyVwReIbFChhMqhsz9zW8z/mP1l6c3khHAaZeiUCMlle
QNs+FXu4Mjrin8E08zOKWXwE9R7/PZ0+SPHJMDHzU3BHFDXIQLkbKzM7fX1f4j3O
g5QfiWjMXlqsbow+OtTJHTsobBIG3gfFNDis/bj2jRin+EWRKFuTdrhr9Q1Vm1DL
06SZsMdYokDckHSYyYq3Q3tDn4q4CF6pWRlVPJ4SpWHC5wt4QHw2opKKewLHbIsa
C/Y1nq93jXQhCJn8i5TR2nVtjlBGDxKZvj0uIpKq8lqM2sHs3fe9+Vey8Nwt+RqB
V33BmS+kZoye0aEZBrus0DFjh3KUxup7wo+lh1qRAR9ibDd0BMZcEfaJqcdU/6M4
15dLR6Mowx+GoXWu38f0Fb5TP9YJ/7vMDS9yW177IL0jUeLjmsIfokZ/eGsTnVDd
hRtbPCrTBjoGfpnujGyLk5hiYasoOHbs9pKyjPYmkVMl7IJckAl8JqBAElhXXJnz
0+atrbjz5ybo9ceSARR+jIGggpovinti/MZERLRf8ytOSpkaMloYz13fmR/Bb3V8
8HD0/8QfxuoCJV0PFWWae4Qye9kTZbv8/TArzcp2/q8BWqREuzYkxBk34Sl1M8IF
G++kUV5d0wFGRZPCyRldIbr3vXys41T0Fl9HjwTTfGWccTOv3Ch2SYR880Q5Gvop
ddkn9m6y4QqJZb2Q6QQF2d3BOIs4qrxuMWCbXb+ky7Z2fBYOGejPoUul5CwMu6T1
yuLzaDblZ7dCRqop95NqKnhNoOe83fOkNYUHhFPDUu1Xk5TMl1u0bJZBXAEYNCNe
5gEOlIrHrBYf8MR/M7QmVMQKmdRb0HFXVpBDpNS+l+O15jfbPn/B/GHPkqkk8MhV
1fabIFwvwH95RfXKQktqKwzJfw3XNFXU238cQrRtWUp4Um3Q7djJwsXQCiv+XwhW
okXirIovC34c/tsOXhP/rD7AGTAliJ9OGtrsRqX42I/o2wL0g3nKtXNYpzGFrVsv
+touK6ah2WWmP+Y/XLJ8YWnw1d8lHp4Fmj4DOjHHiEoZkF8dVGsLKuq7aqdUJTr0
glKbfTCjBO2eBZCXpSl/JrQ9xfEFqKiGCjUYBV3QWCOpuNbk82upRWOz/Xncqvyo
kn27D2kYwjtHg6yD1E7bD9kcyjnQIbvZHjnGVzd0FnpmONduhVLHhGkZYkZe8iSE
2D4ff2e/NvU0jghb2EH4O+KEr2/dfmmBJFSUhUPDGWtwCBw1fnf6faL4xKI8P3Hu
nmYz1NLkC1avnxgGKpblOmpw4BQ2YXFooD6ppp6JppSQtmZHz9iWK+NXl4/EOxrt
Ed2SwWx/N6DhJqVOyRi86RPnBNF9UdQ2cPsEgoT68lYiD5+b3jsAB0NwVZQqrty5
90kwmnUWzNC+r8hJbihSnIaGEfSeNiE17trs9uoIN59DvwLyHyXEGco1gbHpXfeB
wWPXlMzSp30pZNE3dpDLW9bypcFxBLHmYkQs69yhqj3jECzdjtpEOhoK2K0CbHWo
SQ9neFvRA4dTLZKrxSGbNS+rbgVYwH/CQwDYEZAEEE2ZBh7BsPt/t4LaUgDpBUuV
qDs+hzxOH5gs6Fk6esgXt/OcBYqHxPkV79wL+HZHXfKSagQtnYu0MRw8KodfJJxD
+2dogSpJdWw1AsVmgyvS76Mr2JRAyxFrjeMZ/UgTTQUVY7jb3h1fmwa9JLqsuJuB
x1G5NBZnj1jPPQEs1D6AuWaGwH5q0wyiahTlyWS6dNH64M2/AegS0OrRVPFam0t1
LYqiKZj1E8eEYQf74PE1asN33dnr/7QR8T2Agk7bQRSFju8Cn8nuGepgM8j5kcxV
9NiwRTC2l2X/WjA1qbTuYEWk64rE4dkh1UbcTjJ2fjx01QVM/bTJE8fhhlXGbSI7
IGdoOr2Mx4M/kLAnaa2atTKwDO+SGrYyChh/hUrCNwNFeBvBSYrSsjxqsyeTEQ0R
V7ZvoUzwi3/f/BPPpRZZ5LFxG9uCIdjf3b81t2xcNFFnm3mPVz//wh/vT1j3cxlF
ej5fHGrueqM/c5gPF++tc19lWnOWvrMMeE0pp5q6SOj7iz4i/RZK7ARNLibxxj9B
gn8QV3Q+tX5pJDlegnb2q9cV2xxSxPOPo3cf6PRlaXKcRzP2k2zSdryC+JKFXM1F
m8D4mC73C8rpwtJjD4q1+qvOa3UwEOm+8yGQWhss1mAkbkcuEzlwQlwBgKQuRyVz
pNH5DyWTQyZ5i4P8OpZUjU3SuuHid0ohVKMZUbRJN9J0HUnJ6ZXlGVxFmvxN6KT+
PLMYi/MerMjnkG+aoDgcrsZvEuEc2qwbt2FtThvTWvo/2NJIW4GoPWyej20bJBqQ
/8i42aiEIAMtIsFD1etCAHOop/Y6JQpP5vr1zU13NN4YLwCmwz+OHrIgyFs4C+Pb
BYBFEqNxk13126gxDEfkuQA7tDd5yQ5zXEaELZsNA4alCgolX8GZxgJgoHlEJspS
RCtClQlTpYJCAtRMuCiByQS6mPvfzf9100QvP66JSNRAnJx9LUSnoMWJK5WPkTVl
3y6iUwV+7uE94num9ZrkYrIUT+FJWnz0PzMhUfOV+VIrnQxq4W5L+OKnqmO2Ipcm
oPhA/WWYq/IgNQh2B3Afjl+je+ntuxqP0XvCfRFCQrNBmp0p/CDCFUPRr3ZAvLqz
kvqMoErOABo//Mk4Ysmw2Sv/m7TLJhcCQwys5Opa1lx5Hb31kswjwSUAh/JWFdFU
FQi0or+TZMV8/dhcKDMn+9XooPt0L4IC2PurikSKN3bBSro4vb//onzKvg8wVGcw
0Dl3cPzTmgUdqBmkidSH/LPMj0q0YaRg9vOgA4TQxkURlwj33wEcUQYbIwon2EM6
GnPgLxypKR2X5n5ik6r/7zRqlz28Bc4Ui056H8W4YI9b+eHxkr6mXDEwCAm39jsL
O0ZTeVMuIBcwvP6YrX+kzxyiNfoJoJ5HpRvXDhi7izff/PHHD5+B5miXfZmcaYwo
xjrz9cebGJR4uuwWhYh+kuFUv25SjQq5c61TPIfwwOKKF5Ee2y81fH3Cb/ZlEyhF
19wI6oZhfNQdcDiuOmWNcBKEY8HuUBaDfEFaF6CF52PhcfI28YZiCkx5tzcK/EGY
IxteDEMIg9Gq6TVQ09fAVa+2KHM2IneuZGhxpiXF64np5iC0E99N3T3tWON+mIQc
4K5yqQgI0v29EXzTAWODOVCEbE1sdk0H94d7wsvIGP0DyuZclk40bsRKXUPE85dc
/nnMfmVkr3sJsCKfUZaG01cLRN2yHL3WUJvTTXiAz0kxE0lQz6DzfDGWZ5ZGh8lD
H65GoCeYmte1RtEngVrTxrSSzEfSUsyU9aMSu8AArc3Hw4SnngjaZTpHHstYfZBt
+SRBfuzcolIlwpxyMUyRo7jxa/xu2ffyY2CIaM+y0D3lGwgJBunJ2bITE1LEi2jr
mxde/96zLmYGuXvq3RiHw05sbfknvRnL1e21aVrUmQjrz285Xj2Ky9ZjVFfygMNy
ph3nX6buiboMEVecsjP5CWtbPME+GOXqmM9scsd2jl0OKBP1Bh+cujKq6l+akT4k
IrauIw+IPkpeI7VBtS/oRKzQ0Xpry2SrsXhruFkSXL0eQW1QbJeceUZO9QmFDXMP
6/e5b+IEhiPQErL8N0AAsS7HnTb0ngIJuHCwxnv4xlGfg5Top4YIg/BoqDCfOwwC
H5opS09Q+Tm7Ec6yWGHFd45Tv2e+VU6JN+KaRNQeQ8KSBYigCw6tgzYRWVjOxY31
fJU2aO40Ce5WfMI9tAIlaf5zfFoaDrQ8fWNXb4Gxa0/wdVOvZ+PkcbAMrlg+ogxS
rH10ykITxiZliybamR8fcpJFNHb1+LpYGJgUQ4jum+ozP9xDH3OEZuiLgsvRl2f5
hOzwDbq7dvjiT3pau4AUSH9N6TG9NjSTwGJN/uPGLj+dN422sd4uPrAmx7UaggM+
TNYQIQ9+pfTWefQW8U0ylibmitlKRQuGoFagkCT/uJCGNVtVOexGAJDagP/jeoZ1
Xz5IS5cYFXvUaq7haB0ZbNtjn/Z/jP2Vrc5V/Fx3gM9/ZHRj9y+5ocYPx6jjOlFm
BsttvHCjVg4ackQrUVChzrRghKojtBykR9ZCjHP38EeP4yjxNg1e42THNzAa5Fqb
Xsa15/w8JHcUvC+y5FuKuF5xy3oY0z74/gqoJiHy4N/ccnGULpulNpZmiRor4dQX
qv0f+5rqjpArP2P4iwD8s5/SmIuC8ZPK2BK90pStWCbL7afLWiXtUPkBL0KCbdHI
QggKcMxRuPSKBJf5fEtYWm3UITCAW+fK9e0j7az91t5EJHj/WD1rAtjnAzbBm+or
49qxb2WJ0r0CcnA0Mmr7mw/axfD6BnqgK2rNFVxvewR+xPYW2U9qApDqTCzLTUuC
nQKJnFnTl3ifppL5/T9TbBJSRf3qoACz7jDIvzPY8RSfMiZXDLxnbVvXvwrAwRXT
v9MXdZXK54KEbEqM0oktNtzvbPwVouSORxdJ1tkYDYmwZ58wAxtZnYDCOtOhkokE
xF3nAiToClNGVj7fjlSXEN3721xZivW3bfzZCq7Y8YCmovTvJgx1Bfg3LBNce7je
pk/dlQdgPMvEjRNq0Ep0ZRl3EICGyyxAtMxLUyuVvDzxrBlX7XfNC+x70aX/xTAg
pGXK4onagZmawhlrPVuEHDV5JdTxDX0BvnkD0itqDkLHs8cEvAWSzMLhaa7jiYnc
1nAw0KrThm59R2bTKbJqfjBw0njtuuKF+Bj9W2EzeQcTbk6ZpGZRt/Uqc+RM5vFa
Tc2kppQ2fgMzVv6cLVo38enDM2nUK/hal8wclReH4hNBoYPk65LHDg6yXx+CWgMS
4CAGnB2Y1Zw6bf/WedIumN9faxhmsnHBpkVPn/rzofw6OEkO3OCTSPOZiGSAhDm7
Ec6m8n/aKvpE5mrPkrG/9pDcgvFXjdIpfaCJa4U+KWlb9eBtF/ZB90kOFEbQdFRG
VqwEc6RBwnHugd4fY34E/eb2PvHE+FQB64+uylb029cFBrVhmkmF0j+ykl4m8XsQ
PE3QTShox0JSRr/7UpS7m5AyVCCoiP0s6JlzD/qOe8wRu3peO0lrgtCHxGAqXv+7
oyrDICOSWqRD8rxHtS39Jupf1vxT6XBbi3oQDuuXtU3T+EnwnHd3RpyjBeja65E8
n2oP2ItKFONaJXxXudnl7k4f4agbVvNF6FCjDnstMRT0Apv59qoJeVB6V1hWj5SP
GeFGWg3YMCd8JCM3+kmUTMQA/QhgNbvOEGx/iqWudZfXsvgthlDdvvk40rYxcH8g
YbQI0fukVTVuOqqaP1srekQlH2lEmdZO/lFVo4iZwhaHDX4b7TPaxP6Q/Fo0O3Lc
zynt98y7RnJhkTzx1ZRgywdhoiA8l9Kn/36e7YHrhmAHqyPVRQvNpzCC+q7iTXjB
Jh8mn3O9T10wf0orqBVEe6uRQJYXrHyLKNLoJFVD6bH2bl6QoMZkX8VLlaYNBeKY
8V8eslyEQu6A00Gd35uQR5vl2qu7gHXKa5AbuQwHjfKiZtpwNKDrcSQuOQqSY6rT
NbUV0ECDQQ6twvBvAKvkfK7IJGdibbhbcrKEdMLmLDtDVhHVQCxacvq6WosZcViW
y6O4GJ4+qZ4A7IJEI+e1y1wFN8PlrgdU7D8CvGE2C4HMpwYEMxs2Z7UAf8GLeSKQ
JEMDHqlFey/KWx6Ge7QtXchr4lICWQJS6Ktqvst81A0a/qNfVaB9T/NhvnON5gvE
DOj51EKJLT3DHjnXjh/jdcbVx02cBolJAu3DVPOzc6O8wKynN1dO8heEfE0B4M3t
yWAsa6TCO/rCICeP8gBaYqixI/6rL7fydRwqV7imfVfY+k0IzGG+TD4ySHu0p1mq
6EFuqvpmzoTA0Rg+YVhELvJimkgz/5PL+tHQeGcwZAVLvxqTI0VkTN11CtTSBexL
iyGy/DOE0BrEXzbgJnXLKkc7D6UunLiRyZOHyXKwwPC5RLJNr39F50bCc2131WEL
QEXtFJGddflRldDVIhO56Knnyb19ghxzIXr1VIxdWgUVwGqLizCo0KS3Tg/GodqF
ZlKqUbvbRZt/O14ggMpTr2/BdZllEW806udQYWBHd9w1dBjOR6cR3omvXLVBSPVF
rKZJ0uHUQ+GOR5675IGvWu1QHjIaelsVgh1hS+M9hh6+U+9WTQ+vWG0ClTwXLuMu
5bsVL7KAiCA38e0de4qGm54x7wRqAH9CsqhrykjIdQmxH2zRlsu2j8z40HEHO/hZ
lVqZ6zGr/3+aRRK15+Fp45n7Y3TiuzCYjC3adEuCL+IHVldlpfIcRHwWg1cNMIte
JnNvFnvr15hfhZq4UrbhOLxS+3OtizvpyT8NYY969jVqaOlL92emoFQ/otYizYE0
TdwAHWlPPALgV21WQGy7SkOu314W5+lFuAjESt7j68MCr2WyrP9oTOM7/zLXXwig
NXFvimHy7it260Krw2HmX5EGF1thYyk2jzEA7Z/JhgOX4xA5sCXJZ4TsWcGYzXXC
raJESbdQQfkySEnVHMLyiszZAiWrVV7TaIb7gpvwBl/c31cWjiBeGsGKQOXFO/2I
iOAF3Wkg1xebhDLYL8CuB6n6imikJtM/hOwhCiHQlBWENPL0J4bFKnv07LqEWdjk
3nMxKah4dPtqRACcRUpQZZK0l65GqaF3Zq2B2m8gY5hOI9utKNkheUQhan55Be0O
3JriVAIk7SAd3wfyq9NmR5wPexMHX7Hsg59x74fq5D7GvQrLNLDwMwJX9pS9Xqnm
BecSA+KMW5p1EPZmjy5T5ftOPM0tyc+FN13SoV9qOKOiqYrimcGAhwlhok2//fpg
fbH/pt40GirNvwmijVVMQckmFrC6W5lAQKd88jcsqxhG3y6ds0Db9UiTccRN2wFU
V/QHFkWAoljmuVyZ/DbT/N1lPxxcMk+/DXBzSj/NZ5B+nASGLIwKWSIv8qc2IH62
9yRtUBVajUnNwYMWCjX04slf2PWaS7n/9eZouYVi3VFaiLU2J8SN+75A2j2FsW/O
V+SpTgCnYZZZYXqB6NphoBmDjoD6rfx79Xq15BHWAlk04QeWSQ83vvU9nO9LdE/U
toOKQRygp9RX6sS+B5HsZ74TngVipwWC5/pVoy8/4kEEADC9h4QEkPKYP7nDVjbY
xkc2Nfh4FJE9Sal42FecLbx30U3WWvJO5gazfHvA/FqyQCa0SBO9wO1gemMhgEk+
gchWMPA5F+QJNrynPm5Dgms8AaOIyTiCI68CdG43SrggZIrmusXtXq9KtTxka3bk
mHD5X14mf5Esb8xLLrVXwOERfPLne/GA6a+a/LHufCiEL6znRambtpqRbJBukO08
qr2TOae8anysoXSqCA77amLVgQJpE7AcQC05FlbN0tYm2KtKPOft7cX8FDjv6wEC
kFf8wUp9o1TrYkFkRi6fiSiFNew/YI/KmFhVPf+fSi3XbvMx3mIkeXqtXzo9PcaL
yTT+LtVvQTcRjKNgJAQ6s6UXUmi/SriMz6PE3Aj3vGffJWSY2se+cYWttjRTDI9K
0JeUqy47nLG5NUXQxYLJY/pkzt3xoCwacIiWfWbNcWWZF+dqNss+oZLjLn3PFUVY
hYVzKZ6Ev1N/xNQ42g7PzUGqdcvqFAuQ4BgliTdKtRYh9QHkp7Bf8jGb23ZP8JuS
IyJ64xw7xu4J5ihYNRkMetJehtvavUP7Lxohy9bCnwVFIUWyztvJGt4mSCTa1Hx0
zgIHUNKEoKT/CUgHK0pHDyLK98x2b+wWO9tNvVOxVdyFQFrYqCFHSueKLxZ/ABPc
bzL66TWBTWuJmQp9MJCDtBvdSjQU7CLQAW/RX2BNx/2SCBCMY/G9UBdYN3fg9u6K
7lzQ5lv8jRH8HrFS/Im3M3l4o++Tf0Q159so6ZNiKADMex7QLkzmMbP55ScXXe6T
u90X07mITAzcfidvi25gGwLhPZqvtvICy+p8gcnQARzwlrxgmk6SxhwgFIOIib9K
bNq9NaNxHb+W91HJNUaasg==
`protect END_PROTECTED
