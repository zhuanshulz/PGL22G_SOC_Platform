`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lcUi/HAcvTF+O6tDlFnmzAgpxujM/L3IwsEXb60UlgZcIHsH83JfmdUYfelIkWYu
BbqyWH+tOSZ4vxKRVa77OJikVuqBrL/MEKZioKh3vVJ3e2uPUNe2BpN2dXVf4RgF
UkNHE4DoMu8m4q9ykBvkZnVFJSpftZidmPrXHRKFcM6N5KRNA5POV2Zqpe6S2Eig
q1jwxYnHTiJp5HptmEaBLQeHolNQRC8NM/kud5Gz1a5gdLh9rt6TZsBdFKUAzuNo
lnAjhOIEFu1CDaNe/P47v4sfR6VCMyjq4xA2xp3aoLLWeMD07wgsld5rhhMb1nsy
v5pXVIPbiXRIQALtLk5FNrK0mleuGHVI5uwJfZ4pW/S63irZ/6VLM/s5XmHzJgre
kSfFck67P5Pji5DZUr4BUIzyTOhRcPUtLcfTjagXKsodeYR1IZrpCNVNIcfF5VDO
`protect END_PROTECTED
