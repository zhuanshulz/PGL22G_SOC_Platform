`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
edSXHhHTAOlYn8b+FSkvDrAsj4wSJxtxJytSDTdiPgUg+8AkdlSKzspJagK0ea5D
VAYotjvFbU8wU5sVr5Z01Xn6h60c/3ztbFdqECfpSysM+X1d0VpNhY8OIgP/7Y6r
flgDe4j8uZRvucqdRsLmFrSEJBIOoKY2G+wLg5DPK88ErAMsw00La1vC3eFmMqm+
iFrgtXp5i9t5T55KUiQ2ekcY5uYMUzOuxizBD2B71xAMNSZObEaWcSHUzAaba3cq
KxSjREaLNn0fyKvNxzhlm5XV6pK77gzWHVx3+rtW1BsP/yYIKw7djme+KO5dkMIL
TXuGcDjdGKq+A4n1MJ/gDtxiws1GDZNSRLe/oxpY8d4I0dDqOMCICWV9T6XiMPEo
QXl6nUyHjMTekxMMOskEiqigGxr8dUjWqSxaot+Uk9A6KcowlC5LcE/6ilIXpx4b
yXaP18cAaoal9vwmYLefSWhFQWQOXmOb05MFumqZuMs2w7V9BszKZjinmmtK55YQ
eAgzVk1i7bDmlX3Hillqwh2pVeXbqTHTV+zh5pW+VQDyfn1WYmPi4xWXGwL2DbK5
5jRmTRBgqQzv30fzoLtm2u6KUWGAnri5Li2v86MRGs9MJUq5quaEs2jVg6yxqoLo
JfvyADbgQUAruXe+JdWdYwa5p0DVmRewsBxP2GHZ6t9Br8GBLCcUy8EeLSTE+7Lp
oZTGY/1Zgj4K8A6v5oU/uT9ipM0H4Qrmm8/PQhYILfw5nLV3hKXLesDw74Tbea0H
0cgvROHP6uiKP/hlm1IukH8Z8F0X7vc7JuQqrSNV8RabpfW5CqxX0wh82nJEDI07
dLaXK+bVnPvXu3LmUo8SGGj1pSc5en9yarejJG3PDfAUrG7RDKfm5QfBDpK/DiS7
SnzAYuNh2EoG6mPCdj51bap0cTnsLz17dbW7yfn51TLgRco4h4TJTBVo91+3aFtL
13kfpfBF9HOKUieD+stEpYMkvKwFxOOlFMbUrzoZ5PA=
`protect END_PROTECTED
