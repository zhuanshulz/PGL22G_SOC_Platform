`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+nyvokiiYt8ON6c9zsiAcgnVig4PfDXZXaL3pMrXX6sxhPNZLsIxT5o4k+eB/GYV
FW5N+cbfk8Y+SQwjMywPZVnLNUXL7evGN0SxOqinkI8D2K9UwqgXjJVlWV5c+2JN
Nx5jnPVuxf5zPFUfph39EPrAtQhjTpUFY/HTEtpVZ1f/8SrlrP7QVcIPgN8hvpxU
9eMorp+nZjPby6Hr4mzJn0CEttDVUKuugzO7HS5Wa98K6qRae8RviU8yv5R9xN8d
fxPLH8bmCAC8+3VgdFwfxJ4hv59n1RpENYR+/p+n5jLmnp9rbc2grUcyll/oomO0
r4OVxiRyKtVSGGqdfrpCVeIwUYSrnW4LavdFF/3laOuj5PKLB0vbtDzDPUPnbdxh
xgQYndAgOe36B3GJo8KazWpglRt98o3owVB1/Cz55zNxkbATG6+3pzBQoVOgbRFR
BP9dKX50ZgW19A8LvzHXpw5HAyYNTtV3kaAyIg+lavS6poognZ9yotK5U2sRVaKO
1Xm955gC3Z7cnRQGmdu3hLaRqZFywXSFf83aEQc5mMu4397mdegSfR7txTWNdSFN
TyqWNRi62K9PZ3P0hlpO1dHePsUQJCqf9GkHznAOQXGAqSJF3yObZVzcGd8Fxbml
H8aUy1HYp4U4sBbvxuqzJLItExWsPQ/VzkpW/jDfII5XmJnc4gvkP2ZbuTB5i6Tf
kf2i0+SBwhoVGqmyWgHZSM5WSRRQLs/cta8yKp6cKZfe5HrxcafnGpSzDt+f/nhj
rY0HrmP/6oyFpNTlmoPWEF59ytrC9h9ldqoGr6bMi0PONy1lAp03kK74pTCaOaC3
o3tsHxEHKBwCKzBiW/jwsHmRy5+HWfdYl82wSYTQvhS28w55Ly6RM/wfxJixFLsd
bMXFgoKsZqU6VB7r3rlayRt/DWmOcA/6JEjvRVmm/b6N+PgZLwX+uHaRA0pJuBM8
FvC+rZTVAjbmdOMErCOWB9WdGGBvciqziDMWQUJlhVDqswAB53LcS4O5Nv53XXjI
65FwLAzcPtOWMpOGEYiP7vBbnAHPBg79POaL43uFMGzdEu5qNnwXn7qJx5p4PdpV
2YO7+Ks4yKfaTDmF6Imlt9UmPXyQb++okzl2FN7fM4okRf64cgcQZB5OX2BwaYyd
GnBJxtiNMGgTYFp1ma0mZJ1hO04J5gjFEJjEJarnnDouohuLNvB2DgfAydgXqZNo
zS5U3CuVSgEfzH3Rw4lNyQpLUpBhRAbJ0PvF9ZrKlcHogNoU5yMj+kStfNu0Xkt3
t+mxPJylms5abZ+nyDm7sWvYIi3K4i6mvgS6AZ54kw0JKkpRbAWcIMd1EfWwOMPk
c7BSJ6TbwhlIoyS3FcOsjkfVzo8DcWyItYNqWQAmV9hpleKcaVev+vY7iDFAxhZ6
VKJa/CU+vEO37pTXSBtA7/J2Dsozpw4/lzCoRlu8eHvy+EHsa8oNSzxGBlXspSdl
YJk+pjXtDi5DaFAAZH9+q6ccpfZbFjJaX0/YNwIPJhBY6NlNGmB51amdcYIlEl00
YnqAlMh52PQPJei53u7RA9/0gSbsu94XdJnhaL+TYmI0mWWyrjNnGBIk9kfkNmRK
s0NYrHLWs2n/7SOpnZ52+NDwpo0QVSDWfcjOTTO14Z9dbIx3HbDyWZJTvaMHGUuU
FahvKXCskBZOeg8xu5U5jU48YPs2NDbdJt78OEox7XOPkTg86FY4Db7wvBGOMENR
YXG2MP/QhaEAb+uxkAlRrLJvuMQF5QkNDoc8eIs5TqWHKS70Q9fl6kNU/KMCuL8X
XNnuuf7qT7ODKydvVFiFeldqGFELLUXWqtlieWdlw1cmqtqufUs59Kdr3BC4HejO
2GI5dHgp7VvYtYK+WZ34F52f9I86da+NVOiO04ITATYmBIsLHS1wa+94RzSqz9PX
VHe1VwopDhe+GtCydTMF6S6JRtxhG4D1QULbbBzkAOyKKzDNcg3gsD8DcdYzqpmW
YrkeTUDx2soZTeCUk2id9Of/r5HPDK06EQQ2oyVP9eXVn/5S29TuDNfkW4gzPXI0
jzqo/irp4Cdjw9+f0bQ880F5xCkilCe1CfbxmSM+9GXxWCzuyGdM7qx45NmbHDph
wvNjw8yPtdM+ByY3qFBlvei4Xv86jUVZlOkQ56GZxJd70zEMdM9CbylQbFWVDtbQ
6ziEPVOe30XyMSZbtZmQnkP3hSVLOhhE88I5xCMGsNY+gFbOaAKaM/6LhPKUoTBN
cqolAIg/tdcgiRbfrKjVd5Phk3lodBHWiekvB+uGHuqJ7hx521Z+oTFhOroCzJVY
dCKFV4btab3VCO6krbhaE5yviW/IT3A6FHccT5veW8rTHolLAZcXqQRtzkSzpaLB
tJJu3SBztfL/QtzcyJPKMJPoyZx745/UG2h4D2eAJmmJVQNF+e7yfDLwJw/DInT2
QTE+NyyKnyj7MtzP0dwjZ/gp5N+nsMHBeMlDWuCljeXTuE4IvjdGoxnenXhPNKTE
JmOOrYlGMRtFF4uo+cL5DMujAfyHYFP0TEmsdda3ZXlaxUneXUJGWZJgCvVDA4+1
4B3RQh7fxxOWk3EUxmKW3bRpQ826BSJ8MQR3DgU4xnxJy3vMqoG4hIJ+RcvohVvq
JwvWXPaUzmr9po8KXDeRK0mL7AW4K7FOPor+5udt0zqIktKie5yTphxKXhmWz+ls
ur+ragVrtmOe1TvLVsMX2i0xz/f856Vc28zL1txfQmhgLZnan+6ImRAYaBHaLI20
1HeAPMfuYdjPDoQRlOxTukcNAQWr2emmGA0qJXppMB+D4vYjDoxMvmaNYo7hOUdi
zFNJ9tA1sxZU8AIn04e/6UIcTKBtpDwxO4H1rcfeIOfD9Vf5tKZ6rKF5SJ49hQl4
2B2eynWn0M8jdzDeln5sKLJGXvUvdhWofMYmPgGdRnYOqNlPmJ9zvux+Ch3XeHu1
xJ7MNLMciN2nhBwrKc+irP67eEbILrZCR6UoMkc71H+J/O6cg1RzUgCw4QY6C5pV
anbo5O5awnvhK2NjYTKTQVSFpkFoFtR4KVMC+NGAc18PjGIMlfsv2u6J5KX7tK8a
kf8+RQX4AjoUiIUpge+wiLMcuSiNa25H1MFVKdnqbDWieTJ28Nqh8FV0CrGv19Kt
gFTWS/lLML8te8Oz2M8w1B4KSO1EXe8P0rea7mvPZOrlf9WV2Zf6v8h3c1AXVMzg
Nfz0vBzfpldUV2DuQNsiimjcb+X39uBeooQ4+OBQtQeVXlBU3dWpNQrUIRNuvNi+
uw7yRwaP/kFdr4MCKD8tUoo3CZYJKPR0GnrjsEKIsLJUYBLnWeU/LbGv1ExseoYS
6bDn/lZ4084eW5jxWEtjrcwMi97fsowKP1bnuVr1VS1/FIr7NiAV/atPfY6udEOT
kXc4hN4Z7BZTl5EwDh5bKLCTz4W58+Y0aDcp2DTpPiyX9aNTSoxRQ13+HVB9gs7R
4PDRhtHLexUzbB5qg2vKkYYgdDBGssvwBJxJpBcD++UlwIMe1AEbtnw87dVwr0hX
qLAnHiR4mw5sWKEmnfdJncDGiZ8XICD5B03af75K2LuYNyEHTEmL93ViblmGp2Dc
/wYNakQDecznyXi6auEsc6N9e5lUz9xxplbhI1Ks3Yp4PUX8kgSiwKzUfyxedS3b
S8cbrzUwmkzGiGJhkdyamECWPoIMj6xcebKf3fmUQBbeoOt6jFP0fS6BPXnV8vPh
uRNqJ4XxhedJvaTAFMD+qVltr/jwf+Roum+rbI78y05/+vF2Kdb5c/+kJsiuHzq3
NRbY2MCj+Jty1QePshzZLu4FnElD2gPi69tIbXDxVS4aJ2QT3MFUb92gR0EFhyG4
AV588sp1Szoi1zXLGtZ2OB0YpMwSWu3OJdYlSrSfHPM6a07zpefmySvyhbpaVbFl
dHTqgPiDLM12EcpZz+QWUxUI3RPTzq+MMF469dOuRDTyWbtNtjCytp4ljWyHGj2v
LEfLh+FqdOq8O/nlYuG+aOclIQ+S99mgKqH5k7ASwShtXH6gvYV+P73Exr8srBZs
U73YV0MfR259sfgRjodyjGxJd1uXY3amhpStjYpFknwHnayFkMtOeoV1hVIuQwzz
ybZpa3XOzKarPJRJEaDvnT4tPTeIeOx7AWdL/N0f3/2dM9eHATSaI6hhGEO2JLpE
Kt2LUeJvs67w2ZLVTn7iFy4KW4qrbG8665I9Z5vz0uh6AKgnRTRKMQV5GwkI4/5z
FwE+vsRhMeclRwem3j7UMSq8cwBlhlK7g+DmQqJiyNjvOhaurKXyyMMwVYo5eiEz
laZQ5kAgocZ8fxtnySmC62hkzwBQrecejfLxWSz6PRjRB+U6iyXWrXAoxeLcQQEv
QkDNufQg+ZpjOFFISSR5K6l1jPLSHRNZFhHlY+7tLqjUBl297HM2ey3EQPtUZ65d
ORSfxZoh+ynCVke6F+4LKuXfdiebL9uHbUKpsmDivQQFXauwTdaPR/GtUquV4kG9
ww0iKPkR1ijgf9HO9TWUS7tr2FZNXGfRjusBONW2qnTCliqvRmCYPDiaXldAiv4K
JsEsA7HzdiPLahT5MaETQqH9KvqNoLjOqy0dxskLIwu/eTEOpDxwEqwnwHfxHKYE
DsAsZ9WyFbH9de8VH4PxYtS5PtR5EU+c9yKPeFDSUxfuYHXTqr/38kTSZvoS3ETY
rISxoZAXJhekYJHnSmDaGUvlZ0WFhCeGDjbihjaH/OJDW0djs1KG2jF6jUELYvqv
wpq4oPe5SDNSZtxhfjxpE2u3R1fvqbguRE7qe/q7E0DZSgsn5vks1m06lHV+02vq
1CErM5p58eKCjsMNkiFwqFjjwJENMNVxhHdLPdk/pzUBatY3cNNxdW8fUq/ukSIm
QMSvoGMaYEecexgAeEXMFjCVp/VJ3RRU8aQxHZQJgk1tJ78484r9CSRMjIbBcH2Q
jfl0PnBcvEzoMciT5OlxzwqRV/3NLsjIeOdV3yx3jfzo3wjVTb9r3pJEAvTvedoU
P0N4L5Oy7BHY3g8G7wd5h8b7ZwpjqCRa1p+2kGda1s4xO2Dj/+8U92jAaHfxkt89
TZm6TanvYUGh7WIvfd5kRSfJzmoVPOkewWrZMjW5BtDfhQbWmL6xaGvnJIaxideB
SwpXhz9Te+cQLZgjtJ95I99WpmUvRsZupx8qnaZQ/1HZZAzLNkM5VFFo7xgA8vkx
zXvNO2n+r14my9m6+StIF/dcH7SOeeziJIVwdESDJZk6Q7npLh87GDegXaUzZubm
t525eVVXs+gJXNC/ishgs6a+7WHnbTkvdnao+J7BxKb1NqlA3wvmP4cjMBPzIfRR
4JoPga4x8jG2afjQ436S6s2bCC1gm5MbQzlXIlQQbTXn5AHiwqyRksg4TZNb3s8Y
dBoP/xHVWGeNcCNn1O1Ic6aMvhOTDINX7W0+yRnDnnHk+jFBwjU/jbx58CDXOD2/
IE9fX1Q0IaISeb/g76YfGrlPiAFlxPDFEUJnsmBeLjMN2ep1I1W8D6bnFvQ87e33
cgJD+DmFufIvd7Ob+weh63oKiPDDD+iPVbptATh+deqg3wXJYOUQdW0PRU3M+/T0
sL2X7S4HRz+A8feW3yB0ZWobm3PTT8GkQMdZT/Ri9gmNPYNg8BX2iqD6rosB7Br2
v6nQzBb1nraDQsBvsR9CrbzxoC0T0mn8M5HnOklUBDZRCYwTAqW7IZBNlkCHiy2x
p2GqOpJ5xEfLtAWwHC7JBzOcRFFl2m4UlElQEwfw7GIovFFXd6QtYU4tKDzJ1Ib2
bGVUGi+ZmSJccRSh/cfcH3jso7NF7KSzR6N4ZGtlAsZ6+78XXOEqkVK5a/qa9lxt
+YwuvwelVUuwypbhSYBVb0Q6wfveAQ/YQ2K+A1CBTqzYpBOv9ZGy3IdMwXiZvhHd
OrvsgjGGHhL5T2rC6/dyVeaghtxZhI58jVNlTWs7LcPGIFDOr4gaetK87R4Ubif1
h+HyQQDam1O+viGLsxbGQk8kC3bB/zrd8YfWF69P1opX72SrOcD7lejEV/NbZafs
f4iqP637EvLkDjJLq6K9E8Avm2tuGS7lKoD/AIUwYtAdrcB78zm8mB+3Qdvr1Kmi
gDJUMJ2tnVVs3ZFZboyxi3CYeXxQGYYD7Uw4NHP2MZ/CgSSWj9RR9a1zJtM6iLEV
69v76HqTFl7sv4bOeCOjlSmWB584kXWX2BaffAdP8XJSWRZcoxwJZd+VLmOlRGZ3
1GkM2P8Bbiv55mTvcuRrfiGlTX9613GAeFX1lL83s+E=
`protect END_PROTECTED
