`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oyezhJWEyoMM4qcvBJJNyemRNuZ+wVATuNZxALuLW99sJF41i8I2tFeVrVXm+Hmd
+hnMGRk+XtpyPOPs2xuBUxFJKoyMZLV/wMSS9CKtHhXfEGYD8L3IGuWbUKG1UCoV
EBtqkEGmN/xH3XHsbiszivahH4VGPPE6+NUCMAnRQrW/h/EfgO1ktu6XH4FNWnJy
8lbUpdnjJn6yMwmiLepvRhH9XVX5AF+zcDCSvxSinhIHtJ/57WySRa2pSa5OQmqQ
dN3Js/2mAQkZZqzOXcA7ppOd8Micuyo2EZSsL/fxH4tTh/W9o9t5TIeG3vv5u/pw
aaXDa8Dh7N2PTEZH4wXSYu4G+gdpjLtqeEl8RQEYBE5ZMkNyQv6nYudD61Hf+a6+
SWmRkmSadEVEPiv5yThj2CiHbJtxTZj0NMIo8xaVYF0hnqFKhh/rKOUFoqbZ/JOn
lACo5tyGKAG4rUnb3190HFlB8kGtygk5NIpPzIaSS22+4e+DdBDrdQWmsXdvsxFJ
g+IhlWUx9YDowM2ycYubbOQP4U3g8bh3JjhJSPAsy5KkYKPtZHm3a8gRPMgZ/JRw
BKuFV8NR0YztZeGZCPaR7A==
`protect END_PROTECTED
