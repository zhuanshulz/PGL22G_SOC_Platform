`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/K7Mo7SYtTEslv3O+vmLFWWYvfHX120xZsmI0JKfVuC3FgM7cwq4d7YQmSYhegix
gciSNASLvJXdjGwbaDoCEo9sxyHKBDOfk8OrVI9BdHUDhcHXwUhiJs3ilN+IA5K0
oLCRvTVXp9zAELWyxuRrOXki0CX02N1Etqnq9VEqky+gVI3eA5yyHk59tkCMswqu
RkDEo/U6LjHa1yIEVH3YeX2xohyQZF5+bt6Wi4TVgb//Zzqk3va46GvYLNEZQF34
APU5ifLZ4kP8TByKcNULCg==
`protect END_PROTECTED
