`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
31ImA9wbhkfjy/Agi4dsQP5ZcQhKL4qTzdqBYJ5T15RQ54BJsYwVSY5YtLfON7/q
ieUKX5zqmVN7ouMd2yrjAUwm6KVbdTt3KAn3xfas1wzDalmWGpyRdYzJ2SSatPj0
CNDBR4Xd4m4zBY+DhehLDqjy+AFJmhiazZtBsyyCByOaATjCJFMnpxqCCIvZ2cl6
HBiWy0ItGmqTfDs3t+5+lEbOdRjmbcffawDI9orORrJnR8omGarhKkU5lI5RUq/z
9loA09jQeY7cCdl4e71pYbbR5zkNzJjEwbiUjpaKuNbTlKkAVPQtASRFbgY0uIAC
CGe2bKnfdm38j9bAYwqE8YW0zUaXt3QabUXKjH06RCxeMPMXDAHl/fo4qRUZGhp8
KrEthc9/SNXUGsHkUYPeho3Fsr97hBA+VnmSlV++uNFtKLphokKaYAssqXeENmq8
8C1vc0XaZXDo8joKGtV9VJaPrwAcRSJoFcIpKQ8OIkJpVO6YBgkZjrivvS/OfVNH
`protect END_PROTECTED
