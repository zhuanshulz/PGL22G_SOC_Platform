`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zAf27Ib5XZOFoFCOCnCQlZeQANseW426n3sYb8izJCl1QAgT3oXqug44YZNlAach
ajopLzJ3laEskHLjRiV7qNxWjrKu1gHVVC7FuR+fepYnvJDA/xQ5HelZ2nV4rCRW
U0sbk+vRsEpvkORqrtiZVYQCkr8MHe7y9vdqFHAZemuQp6WveTybJ98zJRtMq68F
7lVD9bw6TtEwHNcsoihFJaSGM0MREZqEzuDmcn8snYIvzZaM8pMWlFj0CAQP+n9X
JP9dxt5PFM/Mg56Z75myIQ==
`protect END_PROTECTED
