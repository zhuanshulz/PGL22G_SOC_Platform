`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UmWrXMHSqoTUgyr+8ilBm3GoGKdsC/h4hgmI2tWYGG0flUjWA326pBn4uGS5YOqO
zZJv67DVFw5P/exYlsZ6h5UfYsuZ8h4THe1/XGV6wjAfhQZ23totLXlUSf346V8x
GO9guxCaUGEbXbCEEYve8b6hyy3ogIUBy5PiWWqYQZSePoiHWZm4xmBZnaoPDBll
YY7PUxefTdopEJTbBF6tG4ItHqtQry176V6QYo1q131fS4QCG95miHUyX07N1BGu
4/aE79YJ+XSH0OJfwpUQESvQyzAgKs2pDTfjGjYVujSDpq/L2fnFW9iykjlRQGx2
+r3fnZDCNEjugwveC83yfK/zooeerx2TMop6pK/juv8BjR0WENmVPn6qjhO4RLx3
bG+GtgdWMC7gIX09KBWSoG05I/vUmJqE9n4/IfvpSFomUm/L1HS8JWCEQdHMboDG
+Vr1K2DFW5GziMg6C0dJvjlBexPXMmJW19s7S+5lro8AURNumW/IB343EE7w6heI
h0xt7jdsXV+CobN+ZfHC9IL4LHA/zUpljWcoQDwTvl4BWbsbWRB+6Ob5x0KlyQ16
H23RAiMmVXxu4Sm6/fXITly7rncM7Ul9vldIppnlaUHnxq7cxwFaH7lZM/bKTlvE
tPtQtiVBwdL5FtEBU5ha7w==
`protect END_PROTECTED
