`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S6yXmZyC29i4qB47WCzus5TGjMhOGnFLfiQYfOHtkydxy33fqbQeE4kUzdjWGNPe
yPyr1nBqMegBEFYdfoRCwBM8ZUQr8QhMxwf4aDtXIvk3oz2qrEFd0vto7x2lsBtd
9jt19j2ZVY58nuyj7qimFpeGR5z8bBWYX+g3vE4RJz/k3YxruoQ0qdDlQ69n365D
ta8mJc2RIGt7Ytw9CUz9fZi+KknkQVsOQija2hipybJePnOan6vro0dN3hUNjXz6
cFUHjqiK3u8HD36HtXkCUwmOsGw3mMBGx15nEhDCrRcXaZFd1uPsxp8y2LfBHH6P
3p/gCmEJOueo7ymMCvGHFg==
`protect END_PROTECTED
