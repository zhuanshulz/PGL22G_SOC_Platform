`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JyOJDCATsKO0UMlenn5sph5YxdIRanTAa0srlTjRvfyhPF+VwoiC5YQm/9l9tPrR
snyPuEDllS1HaETcs02eqFmHgIBSx10j18yQP5QR1gZDBGH1HViEQeZq9XZsz5RH
UZDJa7ywb7+R4xL5aiDjKuL1HF/B/hkLrrQzsW9b6DewJ9KAnd3EoSyir2stUsnJ
jK00EeTX4l6QLNy1wZn8u4Ax/3MnB1PzFYUJkp8lV8V3x6IxgjlSWTm9Baw5mOpG
0qvpOz/TMk6nq7gJtS6IRPchdNir2ZTwiV8N7EdwNBz1RpTDlw9B/mqHvuxAUuOe
acpcgKykQPQi6T1BCZNa6OqXX8JXnTsZtAzNDmM1UtWJODzmW4wpqEhXyFOqPVK/
NfHRlYjkJB+2L6LXBAKEASvl4d72AkT0tSKmYSwqxnI=
`protect END_PROTECTED
