`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aBw4AdTas4Zx/HfFgDwuQWwB3a1Ct2OYjHBf2rBfPzwwaLhEeFVteivLu3cDVIm9
nfRjOZxyeSbDO/ouJh8o2/vmpnUtMhdk2dM42oEqVxFrWWdweyc7cjZ1RHBV76FC
dadIw/7GDbxBV0f2QhjuNrt16OfAo+hjsdcwW3rggfvvYR1S6liD/g5wRqCmRe8K
pgqdT7iz+cTfoEFpGZqPI+vgcbh1tzkhvEyLCVQNHPFVwskIUOdg3g5jcTZ3saEC
JwuxOrbAvav8UzZ6W51ZFE+2yNO4h61tnGQ8qyYjXp2uVBNkCuhnUYOyjtZneJsQ
pJZ+m2jn8Vn3xXiaLI9DaVkg1fYeDumMVSGNmvEe4dDz5Ht3RiP5UiRMMnG/VVGW
paay5cjSu5H9KQqHmwBFMCXt0CnTcIoSYDs/t7mnHIJkVVnAan2syxvryBYYwASS
3MutA6vJQpyGClx8lGOrdZHl6PFnxMPkGTFhIY71Wj8fmd9exxmAgv9b4NLee8l7
5ermUtJu3L6ztZDfYs/8WEaCam+5cI7nDu0xBPWVFZ51ow3dPDPDEZNzTbcdtHH/
y26kY2TAlWvTxI3VUFsmYRlPrV/mBRB5+5WmWsv1FZICX7Yr0wtbeCJxwAK5U0+D
IYSXdo853oTfwEG5LnjCBuqOq6Rd2KY0a68d6vBpsNdVNZOFq0/XcjNWCTjuTUC/
H5a+kpZ6WgsVIy3hXY/DI8o57E6tcgCUFRU39T40SpLx2zwzY+mxWqRerBUPoNK7
NsTuKcgPRVNtRbZ28JDSOAcWjD1+ewVaNNA4E35u3EFkEke0r+/SQleHJgDafSHV
8Ns+qzXDMvdgWllU5GxAzwns9bQvxqA31g7pep1duzG0FfNcz6TIcF2ktZ6tYnm6
cCDmEkMCp7iIv5ceUKUIJ+9+/k6hlfrPlVXiiT8F2CLqromVSyGrRf4lnSqn905v
nEweDlh3OSxC38MX/C7MhFOeIB8NprFaxCfFtuL2sYrxxrB5OYGTyYPUCc9CMBCQ
HJLaGHcd53vfoeiZk8270NmVEV7+dljHZwNIdAHUx0Qu3lVq+JDz1EptENOxyzCh
pQE8nXs8AqKQwTZlms1b5mux95WEoSGL40XVWUvACQzaTuuanvTQoOensBk6Wx2X
KEuE0G+k30NlTx7hKISHwg==
`protect END_PROTECTED
