`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YztrFdQqZt37Om+HJBXe6d0EntoORM5K/aI9jUm3YEb4luoB5A03E7JtN9WZj5y6
3qyJC92ysmvcNOYfzqcA1L1wOItk0bsnD+IDs4d9ybgO52jiaFQZ4QiLR2ChJXUE
Te4b0r2CHI7UT9t7jZpn92fIDpFlNHwLw/qVnFvATT5SEfYYWch79ykCHhVasAxd
8jmluwTgPjQKrLnO6arSUX52MIcFHjbMXZHpSe9wyOsx8TaYbl/KRk+jAkR4IFPF
kIAnPg/GLSH+1p9o8lROrNRNEgAJ/9UX+nrqX+feUh26RBOtxWyPQRF07RztQ2na
dDhcSQtRLWpfN1R9beuEWDDAtGxdmzpnULC3A95BNE8NeQRAJa/eKOa+I63Xk1Ny
34McT4y7EHyRmOBxH0IPzVJlTdeOumAqbJZ1KdDZ3APVr5kMvWYI5BFWGo4FBNsu
GkwizCMBmmtCJNl4Tq6IReSOJDkNMy2EZh9sMUncvWXicSUa5lRfwC7KlZKNkgtI
jmNXPsmfO9FbLfHjP9Fn+/lBv21CjIdUE/2pCmKBIaZdyzwomefkJQh35xx4sNKg
xMlYTqWJl4MVGyx4A6ZQqlQlk0Jz6PFLyVpbMTa4oycAdJ9CE2I/DE/ixdXcSj8b
/LN3OUsVV/xI84C96caIRacQAmlkLLyga5Y5Rgei8Mg=
`protect END_PROTECTED
