`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q9wnClkqL2IQv1nbxMVhzX5n3pzv3gaKuyFRH23j3SzgGzm602o6JnEKKUkEq3CL
z+du/yVuWaRgaCHXY1ab6LdAZKqet/Hs1Z1Nujveb468aVURMqyv1Ww8sMmD9Coq
Ta0rfgsLO0VJCYan2QD7b4dklStoRDsYsAKD+rd9fPFNHXGtThW2t4DjPzq9jY/t
0CHgnmxcNHxDKvzqwY1CkXmicbzv207wRbg2DDkWwdYjNz1KX2LPjSa1ZaADnl98
NgMmd1zEFAw0A1y+x/QhiOZljopzjvqIKvETt4fybkE/W4GzB3N3gc2cpfib+MIj
PKOkonBt+1tvdRAeW3OlIZwIG2VU6l9+THajAZGVKrXcTgsPGJQt2lY/f2yuXzCQ
D0+lR3+4UQ5cikUvmaHoSkuC76a/CZYG21cTBmz/sOOsoNKOOy/IGmrKqGRg4XJN
Fh6K6K/G/84XayZIr/9PCFH0NQDHUyZY+3b7Y14O2WPTmZl9ld1xDDmgFJkcQGPg
Pekrm6Rzfo4TmltT4JikVa5lvoYCmUuD/5mJKvymz39Bf/LZOwqReMNoz5QCMqeW
9w5mg6kc3sci94Cz9Cl6/RQArr8PTKiWnIrq4BrTVIw=
`protect END_PROTECTED
