`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RZIXaUN5QZl5JuSF10LpMe5xWllIICKWhcKq36FSOs8D8u8ltCtyC8v2mUtt1Van
ytJvfFM5TUiTK/g7DlfNKnFgxjpVPyMZy+reAj1C/TUcKxlDyZ0sJ1tRTAI2rpG6
Diptl+w/4Nd1/8wt6oeMyu/tr5lWlzJ4MOlbK+u7zW6maCm6D/iOYi6uYJxOurO3
I+pdU3qaZaWPxqTsSrSKT0L44arSz16PmpeulwxSlFMPEfUedNNmI7GobI3GQb/5
VJ7IR52ifmZsAlPmC9/y9Sc71eloiQsEwXT9m4HGVqxYYffQuhqAloKb8fSWxW2M
C4iCGT5aLT7f5RmnKRi/4rWFnpFfWWv85/+fornDwB/80IXFV52mkqqoYfKuVHi4
o9msvqmNWRx0XYBSwWHPxzuqQ+3dfCljJQpckLhNvMdWjcV977mXzEbycxZE3lwy
GnjFFLeItv8sQ+0oLeuPiqqt74oQ+3iOpzPWvhRTO49qTRYP/2eU08Fn5oJT6kmJ
aK/1/Z8hWeDhfhWRfdFsivFGBl/E6QDPf+x5hAqfsoiGwvkMyuE9q2PQAETX//Wc
CBaMa7Giji27G4yulfWQOqJTaSKP4yaXieKrIIb3SEFMtfdeyJQTt3kDsPQG4dWn
PYOyUftxCj786Por6gC2RvGBOoxxsi63bbRZ79JrUmFi1fCJq0shRdrIGKlKx4dz
ruaqGpGM4dYdmhVBz0k6pm5GCtiDpQvVWuHt6802NOBzlowssHqRwSK976ZL6u3B
sLXq4Oh7M058G7RBc39KzjEUZT7T5v4MIfAE2cCu6hlcr9nI+RDJ/fXoBXgohbxn
OtmBrhWp+W1hm5XU+xcqVJR4BPV4Ch1BuPiVp1tKJWe+VrJtjOiIbIMGNSm+KIq5
DfvaJ+bRNAg9UCO/AF0Ol4fbIRlUoBih/LrsAYXlwG6raZ3LSx/B8sSYnrc11g0o
qwyim9edqzewIngvzVb8qvQzYuIeFlmfJkTCuWT3AwEGCUB775OotjFfmNg/I10A
cFSQcyR6bKEf55CPIC2vSEvkeQpWMwULST2v3fjW7lfenMxTrM6kSSt5I7VlrgZn
3sdk50REl4PTw4w/11fmONUx+bpQmzjVbdue7DpmMPdY/NURvSCnUHKRUc5Z9HsI
Cu7ymTCwdxGNVjHA6ZtApA68zLagkZOyEMkkiYTWhyfqURaEXzQXLAvkqja+tvV1
1fNhb+pfCZgDgPW7h1ePplZZAlPJSwM+sBZ5RkpFaR9vofEuBN94o81ZAjyJujwa
lbSXCfVKUE8GchPdQVnxwpac9LAubAuALka4buzcvQU=
`protect END_PROTECTED
