`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y2ZIOMPMogQz9gj+E5Ul1u+wBvP//s7LjwygPhvp83TxNZQw0V5tc3TEmaeapwY7
/6KFCvHdgZAaOL2thySVLlSAOiREquLd7+GTTESG3bcMv5sENxDzUDU80XesEc7B
WhnXB1jli+5Mrp2r5GVMTl8UGnQ9/yLFqvoZi/wjaXB2tUNxXQfM+4sK1hSXxpfl
yaxdU+tm5HrFHX3+b+9n8Q7jfJX5m6UyVHoNdJTZEaGLfmL4VTjcNfPtkTwEPmZ5
CXe6V1F8yhgBzzvLh6y5RfpYc6u9XTipX5Zhn1Umz8TubfnDDIKgr+NCz4huuDuV
gbvYA9GSXqL4d+4D6a06gyGaNfX4o9GCpkoC7cq78Utm15Omvm4wg4WcaCe+sKrp
jzvHDYu2GAlLFnJZy4VSjw==
`protect END_PROTECTED
