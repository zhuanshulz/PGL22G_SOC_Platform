`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iKgEeZYuJgzDMG+HjJyV9rRBeLKtv+DxiwFREuKRO3rIXwfFr9Lhvm0t2j1DCt+G
Hua+7W14H/qDEd1r5VZnSoI9Y7LsEvPZZggKhZDVDyKMu8S4uWr6TGtzkpupH5ck
cR7VRgGGz3PN/cWvfVPVrIbqkhtRQI3V0cTk8BxfNjHxxBZeQxUn0RhyQ6BfVH79
rqT6e393d46huaenCMlAROgcoxe0JejV0Ja5Ea9Ymox0Fod+9Kl3B7gfnr38Dvfk
UVqzHADp42lgqGxruBd3ue6d9Lzw9DxGEmte068sAS3KCTQSM8LX72Gj+I1bqZUs
79nPK4lRO0wTWTFPkJcCkPwr5ABMs/qcVBnUtz2DG5ZfrIpgybbSs7pcd12M6fJw
YBnM0o61tj5yWPpTVSsGEkgZ3PxMxndjWiynrShMW6b6JksOokoesE/vu0+ig5oc
bkQ7K6IGc/lOqbXqz8COxR/BNekL6FWyhnvdSjrr/ZAUzM5WZ+yr7YREx/acN4SQ
shamQQOrOvvC6ZYDzVcYlPQ1oAHpDbswrBdNYNaX+3i0bnzXoQoiNhP9Ehv6zAGb
rvHgA/s3xSeEqw8iUfG02RsTHyHlYMRGT3B1m1l/gi5s0alUnGnkaFgXHSImpOoc
XXjZ2p4MnkHCj8rMieG06FShtbcpKO1jgybSFyOV+jGBjqI0/umEI6GaoDrYjLqQ
9nsVt3jtAj1gfQ10iRT/Gbd6Dp487G7+5xcflvGSMo6MeTGcUDafhaVEu963P/6i
EQE2ouotn9xJBvzjcUkmhkj4UIid/qTU9M2QXRpTtALBIbHTZnqxZWVB2f1Lb42Y
2ee3nSoUmJF93DYh8odLD4oXqc5Fi5JR8fj+9aQqDptwVBRgLmJTr0o1lTPKcB0Z
Mi0FDtso8sl6W42oEMF/U1PGb4XsxRXE6DKJRy3PTjok12q0wAi3Jg3x8wkG4/I6
Q7zHJFJdKIs2jh1PdjXggkjAjVEsrKP4Xud5CNTzENX8s2+1jou7feN5MNdwl89w
qMJIWkGe8OO6MHP400OIHx7AY1PluvE2unLhzjxDQ4UcCZhrpgutAO+tQ15rcdIJ
HcTplUKvwEr4uuwqS7iIEHLvJRa4QSKtd9bhAUpQSmHcbNOmfU28iAhzAXRkPwi2
Ah94qe76d/wSgUtQeUdxxVM7OeDdagPBZ5Ab3Y1I9yqwmKLGnvIs1Lyow47zyamE
fW9u4AZ1GOlidSr+2HsYUp0w2lw6XOgOFRfenJdcuQx6/SeRoiQyXK0jd/m5CzKz
skkfDDuKAlPeth0xKiGDkisum+nnh4j2CeQfuy46BtJCiWxchXr8z3b1PvAPhZiM
iCg6xq0djbHeiyrp5Vk3pLsI3nKj/P8tRJ+lkIIbLlxvqNQ8/GA6MQ6uIblMbDc/
P1oqHPi4lQXj1Ms8o9d94wKe0vWRh2iGNe5YONn4/PQkHootQo/oLKB4s6KWGGC0
kq4ZBeS3lxni4SVQTcJDZcnxwreTzbsiqHqXU2OZyUZ7P0qZLYpTD8gh7lRT1lLQ
mUOA9UkTeAdC1G/+qq0o5I9SEa0RViM73BrBlZ8WHuKccZfRgUMoxqYq6CjxZJRF
JN6mtVF5lspvzYGHj6VhcOBx9ZRQU+CEqz1PFNVA6aYrqFClCqRHQ6KsqkZNX2BO
0nj6xCJ/YCZHInxiXMrnyZfC2xU/Z2EDI4lskWGwPCTz2hXrpOfi6dxv5x3BlWX+
bnuKoeukVUH0VT1ZpzC5f9yCgUb9HAZ1dSbjSF079DdZdqu/ielqxsygr2h+w/n1
xrCXsy9JkR7NMOQbAhJgqBXlevFwytmfM8/4zApbNiE=
`protect END_PROTECTED
