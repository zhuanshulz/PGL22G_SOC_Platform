`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eXC1q43ZFBFQ6gyKix6bMpeCDcnACRbE3N4q109DCT2YcJtj9GwOngQa5AqFwomK
dt2xkDYDx7nehtuGGu7ECHE7M9VL755zLHaUNUUc/94uhJzZ1LjLbXSAB8m+fU1r
14uWKNDD3zz5Eg/VKZZgQt69VWXviaXmKu0Zy7wgsC6+J7j9rKwSopHOaMmVnJU+
oxG3MAxtYulic48qMMmmctUAFoZ5RfzrpR07WDwg35E4qkuVRmNd61C5XOHaSCpk
uZ5tIvN7tIzqr+6OzttH3r+4UYwrVlTCQNdekEOC6H8EnendFXdy59dnHXG2rulO
ip66WB8Cai1Qoq5Jn5tfn3Nv3xWdb0RlWpl1h044BHmeG9MaEYJBWht3J7Hasw+C
pRYk7WpiAqVUapCFnRzmLyRH6oaLr98YRO4XgoVRencDo4jDyhthY71BFPIv0Lhg
2EIP8Sdytu3Sq7LzP8X93uTM9hCBVQf0WqaJWfWDR/mBe59NRevr/pSMWoL5Thlo
hr071UTVpiiT4mP0lop3M3M2gHPiUYDE7kLlroo8AdocnrlUF5cfMURvBz6gtbRf
8qj5nLmnmv1L49UJBT2j9POWA0RIenIRMK1/5Jcd/vJ21obvEmf0+X66Y3ljWdsP
NKl7+RUVWErMvAJ1IxcS9vB3qOeEEoqhfFbxVFQbuaoVKawF3WsimCOywWggUwgZ
+pB7iffB1e6/knse1s4UbUHlcWg2k3yjlmxT1O3w8+fAiQRanoPkzrcyOhTvIjzH
`protect END_PROTECTED
