`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Usgi84NO383sv4ku2QohmbWIMEVj8KrrZ1wg0137jQrTgaR3xJdL7ccTum51PDWF
FuACJgY3yhye/vm4hEGgPPeAJjHfCuZ++7UXmwhCzsiJ4zhqDsouaVhpxDppA106
nbDV898xaDHlS977MHmBOefd/z94j8ou7P//V3+ulZop1eK3ibnNc3noAc3kZez/
B8MQRrmPi7WZlSlP1YqY/Y9C4RM4scW5bMmePO+RN1PMaDrMZesndm8TScTE1z7v
s1y6ulNu/qHYvG+aqHA9yC2UkcGyteqrSEPZd8VCPQZX6VuQ7zMiYoD3jPICGTfK
kwvOCd4smxR7T5K7EDL8HKKlkfq0NE18402KmYRK0BE3A3hx2at+C3izDSLFWUHd
s+KFq/knIsbYZgHBkuLl2BkDXUBRvSzC8E0tNVbiIRCAIAcFdEclTSIWaOv5LaA1
4bNFkogj3fgJIUyBtiTzGC0fGpaqtz2Mt++uFTetxpEIPHDg3P4P2BtTzCJ49m/Q
F7bqPDYRHaKYI79gIQlaV/Dj7uRcjcKnFSzRaWKeEhzXa/C2OHwR0dPaR/q69yGt
EocKrleOhHNoHR7n9fbuwWRCi8wEBQI9iOihfc55GPKUJhXa53pycamXtGqj17U5
sQ7bQajTQB4a2dRHMuhce8bSZgOWPkxzBo8WuvtAs/VsHYtr+XWzD9EDERBmBnaQ
Ngqj2eFxG6E5jwQK+eZYVdLOHay2wIBzWOwBFhVytR8Vd+QzpK9xWZgtH901OFbl
DoceKNxl3lz8NjJG4YaEXFJlJCtz3UIPFmQmxoXRCvuYMYoWfdoAN/M4UMuAu1MT
VMlpwyKSuOLl8ve95SnLltAKBIvCnxB5DXnvnEp6Ysq0Gm0yU+TiHK91o6/uEPgq
pab2KhazNPO97LzI225Jrij6kTgORbckwsifDmnPJ0S87APH/G7IbyQHVJIqDtwq
hxe5pUzRZ18Onhu+TDj50w4EwCsUIW3MesBdqrh91RMbc+xzrYA6ajZngCZNTzxq
BGHN7AXYmVMc12+99pdFsLhuCXwjmVa2hc4gNdxrkn0AK4qwEP/JreA/HraakA/l
EMvFnWiqapA5Vc++3LYmdhYY8GNzelwEewsP2dYeO6/Gw5WKRKEKgv4ElFUtQzS1
WFM2T0GnoZJp5gTw8682DEPepsCDccS44+/ln1XnnF6Vh8x9gXf84uiw20FUxgef
to9X6PrpQJOdtBmVh6tRFhgWYSn9MJLVu7KA7NKDk+qyb0p8n/opFFUVkguDyq3r
6EjqvFSH1HJL8FxumvsIj/oLK4ZrtUoYnjjckbBgxSvZzPU47GyT/VP2G6+VQsKE
dDFDmJNvk4oP3GNwI3LVYj8eVsJMhvRpUSRP+acLE8RQs90vomu96cXFdDFM/4wj
QHRXYyiayA2Q68IcTNDh7ewOxm8oknFgx8bmp4mIsDNc1fjgqzxkXdiyOJ32opj2
+IrZrLCgl/WQvNF33x0ok6dwNui1rqGbx1D4n3l2Thi1AjU92gozqpITk5bVx1PG
3oP7btuzOx/4FUI+A6jTRRIv86MnXc7HWJiLz64B250iopIdPQ3xVmsrWVKnBr0p
ncJE2MxHaM1bTpn/oa/JVE2tbvRZ1ahnVV3TRBepHFjo45yMqVntb06T8VKbRTqR
NqH9d97qOXJykTE5hqs5QT35n4LfyEQPSsRtUjHTNieGGRUtBgVtjveDNFhQrSEz
Xn7w4Us91UHJ2E8npp/MmYNMqeQDIAKt7zb9Hwz6MRCUxZPPNlO9TxWQSkpb3wKe
l+ECZFxKR5kExZWriUVXnBUZdsk7QA6EowsS5TA081+ZqzvddNY1YMv9MJW22i9h
5jnJbnNnaC0SJ9yHHSj1Jxe5+jDW4Dm5if3l/fkS4PrOtPUe7XTNey4fFDhwvgz/
tzg4g9T5wPYJwfJq1iHMqOOBMRXV3bPRDFbFcZt7O7x8p9EBz8IbwJ7KMq7xnIWi
K5E+aYqfZIXFjMqAsvI8SQfFTYpABE3HKouKc/ebvOEJVreLSOU4TDTvWQqJ/gsX
MiIrs+rlhenOsu1ybXMw1Vf6xUXfCwF6g6s4P2CNFzZxm0EYHmYy5GXG3Q0iLnEk
2X1nuBJzqaafdsMntCknBQNJsmsgCuof/Zp/HNQTbRVgreI5FCKJmeiI9IVWc9MR
YWX0bTgQLRHXzlZoZfrhxMga6HpfMcHmCS2gnWnz0IAhnh9LZd/+kBYDyS2Qx+Aa
FAwVNuMPYF+Md06f2gkUFO/C5T32N+SFh76mlWYQVou2hrWMYYYkAoR9KsTTMOT8
LiN8o0HN6qof6HBjeZwUTE3nmGVPUYk2BVauesOqLhBXgv7v9laLiHWFOZZjjMq6
guMB/HRPpu55nEsO3+drOYFsT1p4xOwGlsOlVLvOYl4B2Q8PDhrMI1kIYkBQ++Np
DtR4fY/WekVfvP0RRGiW/jKgsrLbA4wlP06thuOvmcGX4tfViz33jm22tZ3V1Btm
B4AWOZgCJXwC+dH96FHcFLQunNsN9qd3nKRIULdnt7sVWC5EQ4XanPGSbYX++4su
6prnveHKqvTukiGbTj71smED/HnnJVEmyyEe6STT12HIWwbWu6g0FMcWEtJM8ZYw
i+7OVQMoFCLfgy1B1jh3Bneq+/sGLcUgQh0NiQFxzEk=
`protect END_PROTECTED
