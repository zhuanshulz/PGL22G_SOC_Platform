`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WpxU60G7cEqun08Z4MFbEGZZPRZOwzpKaTLLa3SuUeOijK0mFaA3ctqhaMgae8+c
Ilw0wUQZPam6BfxpCcKoSaKFmwBzp4zZ4GmlgkXe+9RoS3QAlk5qB66dL7R4oRrP
UqB5QDMOcFhkIxk466n+Ouro0GqsrEFbZ2325iGrIj+70t3zW4r1mgHP62o9UNew
+h5S3An/DgDhvTkKCtphRkydUNDrnyvuocQXNtPbjvR5EPHnP5Tu0G1roiPCxGhi
kTk1tkEfjCIoSOSIo3SnYAukvfVNVQIrjBbj6tQg9ntVjA3qzT3dckTQ1/24dfho
NdqCKTz+8AaMGfEa/w4aAxmYidI6o5FBsWdv+ptvZDfU3zwmIomb/Um0WOZ7nDZ2
zDoY85BYsFxh9tXhlybJs+QGu5tOElswO5x4fXZfylQcY0e+/a/JbmCJCJvdlbgn
pv9rdXfvNF8j6RqmeREdCCCw5i/OPlY9wMPKf1sLXFgPyBBCIzZUSWoLhFZUJ/Cf
FAbyIVsY+ENV9OD/Z1MTPES/pxODGzHmzsuiobArACLkIGq8HI4lIh5VXyG3fKlt
P/uuLfy7f3r9q6NzGWluFmObTOyaix6u2liPlAIkTxplHoX3yGyq5E7MXA5SQssf
5iGO4+fi1B8m3pSsQ1yDxWJzzelIcI42l6KyQglpBPNiRDGeynEZjiqKGrVCr232
zHb3r2LG/TKL+Wazzv8qAqARTXvgs79BzML5IUNYLDbkFZPdkjmAdvLdeM7CxsEx
VY1GXv7CNSFvHbqmdzMOHskiybRtUfpBiMBoeH5QuJPzszzIoIdd6CDQaGWps+x3
gSEXTJDBPkN5yLvZy0yHt1hBJeCWJly96arq5IQ+GSFvYEyxmONaB+BofQBQFRrT
tdENAVbmD26vDvWKvSEj80/EGL23nyiG02G8JAchLKQwkdMJjyZpj2NbRgK/sR5K
LBwiSGJJVc3MZzZPX9W5iMrFGlWJ7M2YBclIOu+R3qmO0X5ObYZCBiFQTCCf3Ho8
fxbR7lsJ1lqxvoVpA2LJfVC6xlX9ggjAg19VpsCUVTye2duS+3S5pZ3XZlmF7ohR
mjnwvN/ShyRKBkVhUvLTiQVFMyns9MBXVJMQvI7+rFW05pSE5TZFPeg8k5I4qb1C
3D8iSxBjAxsKaVTFeUbMdDhhaThs9FyWBgdb2UGYJoSptyzZZG/qzjcDAtI/EwRI
`protect END_PROTECTED
