`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2ce6JmoIh9YdiB9WmjzMDJNUK+JfdpvL2z6p7axQQZd704/aFuCvl4hppYNqXdib
Pv3WMWU9tgD5+p/OFo9ZvvOjZdlxqTberO9o03mY6BeuydlxX9OypNHEUoysWBSB
F45LN40ralL6tNpBfNw36RQGKMiTVBSsrXmsFJzK6P0TndwXH1nbK3Zz0Ym3ptPh
czP3a2iXBhBiw0F5nH/lPZTI6nVk5lOuo9hosk1g00ldfw01ivR7YKUYdtc7e8ch
ky4A1pcGQgHTUqybidVwWn8QwTcbPqUTLyZE49uWzLcQ4xqSaEafpcdkne3so7Bu
wAFpVW03V2pgUpEssLGcWaL4GJeutMTFZH8HEtTnfdkeBPpjMGO3L+FtiBicVNzw
BC+q3m2A2A4e0c2jrSmXqikKU3LhJy6sLY5N9cj9wDALxwc18lPkfyskCnVsOEW6
MFYz8NcvO2mVoYMtklSl1ZdIQH/4NAt/VZ8TTrY9HQvSB0pRvD4hzLsHVaFZz8Sk
L1MC/waQwf/uiYLFMHrpcUaOB8l4PRpmiEeOlb5NRj8YEMrSOrwvR2ldimr09CLE
q0vJEM9t7hAGihxh4QeQi1AY8L7JIJ0ukY4o4CuAnfgmPLnL8Lt0J7tYZLbJG29t
zY3vQBVSXaEDSh7242WirQ==
`protect END_PROTECTED
