`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oKHhBRrYCCTqo6ocZZ0xnMcqYDJD24zSgWkJxMFFX2aypNUd/01W+ZcW4m+JuRQ+
j1yib9Sakyet02LtdMDKicLNQ8KiYzfWGg6lPq8NfwqX5uGClDGeqJTipZRsj4s0
o4WEF8Is/bujKpmoc1CH4x+cEtSO7jC9VsLb8TbYDlUo66tNijC2p41RaDaWvc5U
o3oLsFK1jhXmXVb9WngNtC7ptwBrx5Wnfe00MgvYixxG+BXY2BLgGvKdW95vNpQP
lPbsOpfL8j1dGsKsqjcAjHtyymYdg1rB5BVMkkiULiiRXiBjbm2Wo5kFlWh32JaM
x5oYUq5lVps45eBvHvBJuYJUCGYcbAIA9A0W/02X8SQKFS2eYR2gsTbuolJBTtzn
gQSFjM+/40dRB6ROeSaWbna6BgGmrUyswSGj7dW88IXHznJA/i4btpLAF298DS1j
T1yQv3dv+6tmNH7pXiih84M8AqGrbmlE3EGiH4E/UIg=
`protect END_PROTECTED
