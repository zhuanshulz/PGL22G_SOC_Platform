`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
czXDMkIEm2fSIcE7j3CeV52ODvh4TKBLJ1lRBw4WtSfvirmrHzQL6EAIZGjDfamy
KaPAiOlnzCzYhHqQ470B6EeiWNfRD/Rrg2auHFylHqa18rUW1ciqmjLLA+WSpOng
MVidGQj+yyb+x4xUDtf8NH9J8h48zoXOeExiMsLTuXBQ29cnZJ5+VwI87tVM3vgj
0hgKzqnKPc0zBqpKdPHJGrhl0UZMLqJJ+iFy4mzjWDQ1/nL4AYdWiczl7/L8qVug
5oEeCDCo+pGoHRouI6o31NGwmg4z7/WlbBNPsxkzuWO21zrkSLyr04tsajbmnxq6
pG1arYHJolSzHZr+BHSMqU8Bsrc13GyY+dmtzcRypVMrcH86lJbGVQtIDxJTLMEj
I7Q8+voPqHYM9Gdf3X1chKIFJdeHxfgIt8n+sbYIpxoqdpo6ORfyN6Z1z7RWXQx0
I5Vzfre7O+CZeZfU8bu8ZViTM7hSmgrxWl6QAXKNVD37KfYlYYpKuHVOo6YG3Xl0
P3AlHX+Ow7dqtfV2v3/EsQb5wN7GGGiRnRL+Gxq9qEXrDQI9X2Uo2C9j99zIPwyy
5VV5hOocnFIJixZhWI0LG32yXZ40b3uKu8s6z80P8wMU0344Xd4/b/re20OBGMYt
yDAcMVTYpl1blapLtLktb6LUetwyzLqdtkCweaCYUP/QstdGyrMAlaReleSWpKxo
vf/XPd+h5PORt5BfEoV7mweP4w3YM4YaNKwpR250CDB6YXXVT1rbOEAhkWzK7bui
2qFSeW43wpL1DwKbJY0PUQgJ9hAoiRymtUZgXhoDCYn1ZGmx+6divN39Yp0VmdDw
c1KBsCfhQq5loYaQS6T1W3bbmxYl8wfka7KghGuQ2dwEsRK+ffDD2ymOKBo4D5H9
hktkh8z2EjMU5xqcCiEPl13+T718LO6kAO5ZDB+0Oswrc/Mp6pFbNr0qw46noCHD
0LuCDJBRO03L4HNJYk7WiHwILGmPfYMkeNJvTuDUM9hFWM9ac14SDRiWoDAEDNeW
nKGSK7SVq+PyhBpY0D+ImEZiRKh77efSoORZUCDHUHTaw3UM5e0cML03/YwjxUaO
rPeCOaVVYYtkmpa4EtK5Ltes3jAtkRHkN4OAwWg4ByoZSBoW5Af6qgEZVQueerM0
cwhY/MGKfnpcwAbFttPYN3zQiVPRcBZQL9HIHiiSGNTRTiNz/30exg5GMGYXtadM
9IMdAHXM36ioS+vFqk43aG1Hd0CL6TpcVrtNrr+EwrBf9hrasOHO/G5JvkYzccqX
5zh9rzAI8v1g42L1wY0pa4rW0BDAp0x0Z+R/yH2p/Yj5eeEQ4g+pxdj4EMSQ3jYY
tb+ndQYetH8ZJKW/Ybf5LzaT0il6DlcEEEKETwsvqxjcfN3salNlfT5Zl+0OguBe
+ub7xw5XFgZaNCv8TH8ab8zIbM3Ja7v78OS1b7fhSG8opYFuadUHZqKD93LJPPNa
6RJPT/2bt6APo252lWQfdA==
`protect END_PROTECTED
