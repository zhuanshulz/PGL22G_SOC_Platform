`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tE5XR78QRkipuGjIqWGiKwQb8YfJmaUHmHCJeBEQ7FTOpmFN60o/KeyDjxMDKYCe
rodAG+3PjlfsmknIMvF/+e6ytF15KGOiKPJBzAEGbAYoIAqTDw6A5xYCoOF/n4zP
PcnYy2xGeSZi/YEFli70Cv+MRKi7kTIxBXmR6J3IBAeKCVIJQkAxBxDgeTFZ1UML
LTQjjhvoFUX4B0j+vH9r31mybhoKKLlieda8IhPZBYalQNUknftFnoSGdWkx5TwN
f3ycEdqyYutYtdhKJtuFCeUh69dY3Q5Fb71SqBY2I0GaXoAQZeyNosKqayOqTIAP
IIaK1b9TfP0wyz/CwGgRs1LNiyTT4Eu2waxfN9YGFDOsNV30o98YF/etOnIjM56O
P9OOcmX7XygrVJTbUVjWlD6e0qhJDTe+wwBc7QKXeIusffxQ0kKotiAE/W3mLpsC
5sFv+eZ0gYG3XUq0BuzifS/dG5tFT6FD1fnxwiQczN2CwTmpdN4Nxm16bJFuHVFL
M9QbqFHRHJWpaVJLE15wnrFKCGtVUj8h6pyKVWLbyNK2ymWwZZnerXqfo+AJ2To6
tZbEuOsSn2BeJ6+y8Nwdmu0EDoYcJrCFYaARm2h+GeQY1Q8gdz6lc8nc7TkcBdAw
GFgNQaCKkkr9XWYkYhEJJMtSITOjkymyJvqQskqzBsCyKM7bUV5ffFxSWfng6whd
/Ch8vDA7+FB07GPCxp95Ap6Dn0RGNwVgG+hq4DSyRKgBSbkmbZ93JR1Sj/Xv6+mW
awrzaGEfFuNq4lvMwns55H3CfATM56gbZarYwDWdS1TWzReLiLZ2QSwDsvloZe82
L6Hk2OSpvbasIWtB8NYxZ+A8IrRWR/eMnneFvSw/kVO9CPaJX8xnngqzgW0hp06y
LXlmzMWIvuDso/oQk1w8o73k7RPfMep582dOia/rz5tO1q8fo7fmfAErivdB3J7J
yChDzRdH4g7ZW2XATUcAA0Om0IJ9ZodMPFXxOUOsYTlz/DZc4AoreqxZFQ7ZLPw4
CBa6dFm4AknJXJ4L3gEhFJ+I7GLXNYhB/Q9XDiYRGSsqRA0KIrTKnWW2IVk6lTpT
0pDavKLW+wIwYvrMM2fbJ2+OkrPdCiezcpc3J/8yMnFcvG1fclGll5uogBUIGhKu
ej5IvJYSuCMV2/m0dDfvgF2pOifOoxv5gOr0FIRuBL9o23g5P3359F/yGcc9/4I2
uyJF4KzCMAYXsFg81FvVwoc4ck1qx3qrS9w5j7tXdKnzj7U0jRjA7eBCrWLF4HPp
bRV5U9S3ZEpBCwpjmnad2lWPwpKXo99zF47m41Nbt+amGbh9UiunQ09xSQMw5epH
gyPfSmuNx2GYEVAAb+LcJrMkSqqdI9SVVKOQbRB6kGU=
`protect END_PROTECTED
