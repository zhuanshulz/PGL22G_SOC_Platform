`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6IyeTu6r30IZc8mKbMXyVX3z6SvQFzDfW+1XWrrXGsfo58iibezwrteuXLRL/5MF
Mw7b9BxlxZHjQJW5KUI7QU3KFDmvLbwVrtytXpCVZx6fQoW/U5pZWCGesyNWStOU
SDwKoBOUBJcXilWz0D4U/MP1OowvMeokLUcSnfVA4YJOzVI3b9Npty2CLIRd+Vlv
qEq0ykhfaZOs25iargrAJYnEQYCAKI075uUtFEbNkk0BQbWYsU2OTNSfJmGnRbHl
G/Tu5LXrjrFvizeaYMsQRZstbo/Cps6a9PciblwS00MpPUk/2lW84zt20zrsytW3
hf7F0zKY3r/IwA9VzgoZOjEl4uLMhgPgrchpCHcD+0Rj//Uh33PPjAYd8Q4rkV8F
RhHqdfVwYnrk+NJY0VJFLcTla+Ez5POVZ4Fe4ntv57OC3fHd7HUMjsCxc2v2R4uq
5Mx+GWpiRwGmZr5xA9X5NfsxWaumU1urVGs51xsT+5U=
`protect END_PROTECTED
