`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A9p69HJTKGsCqYwG/7DG6pAloxLtIZtpZ9STdodVjYCfRH9/N3e4F5hb3GWN5WFF
OEAjmGd2yVGJC2r5pW08Y+FnPLRiD2hWPbOQZc9c11CH10WwQy1Tmr6aHxCo3JBw
JISNmFizsH15YwTGWYrqXkjSpaU8/Yi024UrObL8+P7acKehv0euvViDY2Wb17sm
hHK1PhKUlVxkC5/w3rvE7KEpx21I5X/zk3cmZETEotA++6xgJAZAzqi6Aab7jWYP
IrMZT7TQ9T/04ww5HCTdMdgWEQaJUCyE5yRADUeAYiqEhD/3eTcloJxTlheIkMYh
cS6PjiW+Ga4s8R5GL9i9LY7/rREpmnoi5ce6SWwKGkfcSBhrVS0A8iPU7URDR8R4
Mkkt69oxmxX8jCboadi31t/m5sYg8d7d6lFiJRtpVDAVzA5rrbrMg6eapluGRRDq
oUkfQ3ZyINhdeheEzicx0gS/k+tbqmvDSottwwNGHWIa+gefXCmbrpsCe64RhGjh
pQGst6gu8d2SkwU306XFEN958YuoogzvSzgrjy4b68ZWYEeudpci3feCZzv3M40f
8Xy9pfltt7r1NplsrVUfqlHiiQtGtVbjIAAAVpmP5wXu7TWOY1zj2fH2nD8juQYD
yPxuarGQ5QmKzKlrauW/6NInrVX1wzWhHK/UMI++yRrQ55N7aj0kN0DIffLsjuSv
kzyyPhNZHhNRiqtt/2/IPTAXj1PeKTdrS6WZ9WrMHBFUMiyZTYZY6kvzg2XyW+5J
x7uvD+HMe2rmP1UbCT92yD8UgqA2FJUJYCriwfOldfMxnJyWYX+Eqljg+pqhjkWE
JdomLebW3F+vFWQQs3dsWpqd/nHRwYo40Z7sCmiJb4rXFh+x6yY1s0rNzV84XeZg
HJjQTIpI7ut2boxx4nEDNBE9qF4tXvWQq0pc2V55MGWNSfUe1UQRdnVf3IIYk5AO
8V4Smxp5sB/VunCb3HlavKwpeiwgREjbX+myR2lr1gKWpxV6ma2uCDaaYSAbeXrD
gjtX+F6L4dgPm5zNhYMvYyP2SyM6wiHkHVEkt5YV+Uo4P6pCG3CaD1KWBAk3WsLT
mwhhc33Iw7Z6yiwwn7qhh63LAF4z0Z8TDh/3GQytFAKtDDvQ4/AkFeSDmJNGRPpE
6I8QAOGATHwgifd6TmU1DZzOqItiYZNSwIMOJRNyUJz4AMRgmskgMdBa4wpf6ULr
IoyYUoE+J1Jfm0czGNLho1rVP9lyoKilv1RJT2RveM0TYNe+rS5rFPAKLBnKiRjy
A/gCtzqLZv71t0BGkRT3vw==
`protect END_PROTECTED
