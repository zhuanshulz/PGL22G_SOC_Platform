`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7PccbAGEJRs2vUvhhN7gDQpAwIvEN5xq1h7Qx+qyKk3DT5r7fchpvIGD/QmF2iWU
GrjSyqVoofAWlg6Ds69g+KQJeyfheJZDva1J06eOEqaDqUoM3hKGUztjcQ9dmCMA
Dg1iidLoweWVghTPEFIql+OwnqW6eVkkdh7sXzrDNgRGHQVb2k0Fih6P5SnDllI6
WS36AKAr6lLui0ybLOy3OHaobNd9wlQPYN/SyBG60x6Js/w1qrlR4LRqhCOj89NP
9ZNSxNPwskqVUgTUGSCiwawT+Xdv5l7h0ERDgn/gxnKTpVhRu6vjloyKYKHNhA/P
1wMPDw3LrKJvXRIQi45/IQ==
`protect END_PROTECTED
