`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hVTy8wI/wGAQeE+5vzmknYfp53ps6TWA4MhG3o7HHzNGqx53pNhHpJcHicldU68s
hJgUWmkTIyvE+pR0OzhZ/c5OZwuAI7PPQvTX4LsLh70a/uZ4bSLzjg8PbWXp+xx1
GdVwPKCejEo0XaHf9ql9JC2sWzqG3pXzEfdiLhPLslMl4vw+Tjd3UVKA1ibuSfXy
bFO+Sc1b+wSu0NoHJMXuPmtazqHeTRGpH4YHDJ59fnboIgi+X7mTF2dykfjCfuM1
8vM9DWB0D+tVp0MrG7PruLoIyLNhU4FtfT1kFEVqsNchIRduKJpBxT2WwT3LC5hl
6ESpHx+6sakAgIGmTO2fziEl7bmHlk6N8Q+DD4NDHgQI6kTsm9Uu/U3500skklkI
2QgmJxVEPMJhM6dYetnL5g1yaAGfaMAnJiTbEDuBMW33VkmJFQtyf/M8oZCwyYen
gBxTiYhTvUjM4J+GkFALKzw1lpYq/CvNBaR7P06CxnHIMrpEyrAblKqfoqwcZPN2
fz4LRko0W1gMuqqcTOCX11R0t+fCJsNjsLTsNRvG9lJ4GNgefxJo8zWdLSq7A0fo
ZBLa+PaCppgBYCx7qywvQB0d1W+JphN2R962DeNj6bdPUWiP/y0Q5msJ81eOkgH0
xfaLerrmhkV9BPejc8xNzlOy5pSuPXTuLR2c0bBy0Mxb743kmiid2Z2lDQ8+5hpG
NDW0ik23ZXrZUfXRxsjG4mq9C+z3VMX38L3uiRYUY3oca8e3L5nXePzXcZcstiEI
fEAw/ZgpWDLPNdA9Iw+cZSES3QyxxpiGYAfSXS26gZPiiq2LECc+zU3r1QlhQGRn
c9DuVOaOBaAtR99hfeW51eKRxkL2Pt0Zptn2HhXwwd8JbgEnj4OZITViZUHSowjT
w8vE9OJ6orYVLwi1R4aJqhg06Yon6+KvZlM3ZU3/5aZtZEdal/QnDtP0ZsLz1mMX
AnvDGVY3amEW8RNWmiDAvg66KQdqK5qb2EFOne/H2DKKXntjfQkwf6DoyEXOwN+J
SYthMk5l5DXBfi2rbBfD1z5kTLj5CfR+gO4iVU8iK3cJN6i/qoz0aSQ7ZeIqy/I2
PoUJfNlwjxxnFLPvhq3nvRnG2LwR9Sf2MRB3oDkNBwD3stHrsWaiY4vtMuOvStsn
mj5qqVLYvhxFrdG5zAsgTHJ4pazH9xwoeP7TJ5pkB8QW/jEkgrkt9nyYNNiuVHPM
wP5DZUF8WfN8PC94v8REbUCuJrRD+oe8L4esULMQIFbRAQKyVafsVi3eRbp7CY2d
zYQiiBPRRbZkjt8l844m9MGR+uP5EfW3T6/dQEZes70HVj7L71ZNUFIb8uHl3O42
+gshTua/Ak/g4AAhNdWTKa6GlqJP3Woz7QXaTXuzKpU0qsoarpj/SYfkLWmUv1WW
IaULmTqyv4ZcvV2tN93o8ViybdKRG4Q+rAcYcS95s/mYtyQn/LFeHRdLapGxWr0g
NJs09h6L2dVE/e+HJ0aRJHKGPy4BKKEmEOH+8nAIvIU9mHrQQn4bYAvOSwPYlRDC
En+XJCDt4FsmYw2GUibsVCfAazCiUpUcO8v55I/yhoxQEJQcAmRQ056g7yIuhxgk
qsGzVlC1MoOm+1b+DpFH9mc/pyE/+G3/iZ0wn/PmjCZ8440tSSo2dSpsm+GpNdu0
zVdLTWPfB99ntQ3t6m1cJOGGaespSAegiQ5zeQ+4nvZlYUHsYP4AkRDSWUhhaD+D
koJpEz6yWbdh6y1+/sP1x9lu7oLk83WhsfSzn4/HZUiEmf9zeFhKg8xQV+CqY39s
Y5suEV8E1suIEDJsUkZWu6X8oXT/33nyyuHHW+8HjGbAJViMUR6E1BRS/Z/5E/P3
1RuhHWVdJt2bw2bsq93rauhrHrPHSxniQlZdhQUheEHR6BzIAo7gUEUf4a3p8grz
MC5gvrkv9xvnCQ5orkmd211JNNvz9DDC9DckaqWZyxJXl3hv65EY6VX4Tjtqf6RI
LsY2c/DY9P2/gBKW2YE/kX5h8UuzAnODxUYlw6DDI2DbHqBaDayIK14/Qs+LZISv
OELtz3EfeJ4NqdK/APPSsz9W+Rt07mefnAIxmseNt99oWf+oEVme5NkXDS3uk7KA
VpYVPJXKgd6uFi0OK8SxygQLzxAnTqQ4PVob9VM1zu0L35DthhNGjg5vlp/EcJFl
DbIChqgNm/FgoWTeqAF96OZmvADSV8v4722/KN9YetAgRQM9umIkh0WaGUnO4aGR
jmIFakOxM3TAOA0QsXo5U0sOUzbjqFbVtutCFXsgkyt8id4iBf/JMmttJ/TDG+3d
b1XCe4ry3dVPF4K8Nw1aWJo3+TEHh9w9sxDgqwSF6x8AjhsizjrWXQwN7jCd22Ab
tHi4VvlAkXtwcc7EaW9CUhOF/AmC0Jh2GsQBBuXXr9inBjl5t/y56KYK0GcrvWh/
IPnIl2WIJbtCsJwj6pmS59vlWielFixh4hzJXrP15+s+tnapqExUikD6YineiCIn
Yygy3k0LgT5uAMsp9klB/wE87SoQ6Jz2HspNtXea25UFTHmep37OZifOBDbxW0aF
VbCayKCZzcLXAH9hPVaAHt+jcKJjR0AQOBCZ0m3ezMmcc8irUm4lRKZPjs0FlCd7
efGJn4BwuLucM+ts+ROgDBQvc9NL+DlXVZLkaanPdA4W8fvwdgLva5Vm2XybbAzj
GJMWX+9tzZuxLqMRnZv2M9bVMptuh9MqJnKa1zI8lhyxKTVd257RHHW/sR1mUwak
Bey38SK6Xw1ki4wmt43X/BHAeI183L8tzhBLFvrgOkGeeerjzypxNRcAkkhtiMa1
s10UebVuK7TLEzHDUzJv9hDK78Pm4HXvpXyhu4lRvRkjBmus9blrRnKZGMqEQJaD
u9vqCR7hzt1EIVT1agL1YFps/UVOMFgEeqXucfV9A+5FTNcwzJMKgfCzKE8FpgU2
Ul6LYzRVgt9irxUvjEKdP5Lg8CGBC+nnJIeuzmhgfl50zF2sSFQWImfe5c4gEhnC
sndS67tTnn62RbRMwWiykvWtPyQAx0/XEG8Hm4eskwkw3Ky16+s+dLnQInePe7ot
gxfERr+6LV+1XVzbAvSL7LNBDI+WnX7Olgh6ya0ovi7Nlfr081ZxdO4/A8XE5oNK
vxmbsAUhHmUQHMIXjMEwjJnl2wursg0UJZDtTuavH4eIzcFK49T+tUvcUMpnIZvZ
+kvQM1jFrUzYa0xzmFcfjG8S+u5PVBjPSqHLVxDVA8wLTXU5XxW3jx7YU3gkd9Nc
jlvy5W3dFP+sBli9etHghbopEvk2Bw08yHv/QyUfs+RbcmGER8nQfHHyDszS+18F
`protect END_PROTECTED
