`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vl3il3yj1n8ZAUZl4tqCLR97qXy4fimx7B6wrV18+IJnbrYo83CV2RqMpoHJbQqu
jNy1R3l0u1yq01v2TqIdJijmm7pCHYShWFPsb/L1uvJJCOC8Oqbgge6WKBAsgb7c
s6vzfaTif4nOCPcbsG73POBB91vMdxytYMJ+i36DYWeghl0UXy3MUOSaopoJId97
0X8PQ62GUNOoQECe7tfJiGSpArBEDYi8rqmr78aeehYgqXd/5zUHVRc+020TjN5p
R9OQ9k994sakwGBG2sSRLm1dJrifPzs5K3F/0HHIQyAvTqxrHyeKHzVNFsw+iqZ3
NbL800g/ZwGW83jIh2OLf3bteyOlS/cPlWspOD03llabMw8+oL9DZdGRqrExCEZf
7aYpMSIgQzy2IBTdpSzxqDsAcGLVOeeSa9i3jtldj8vGHQDL1YV/yPYwRUgKhbQz
RtyQqDy4yOfceIHpSE9cnFtP+JSMUb9nDFWMqJT7grlO3aBltWc+wFon8xD6QtUi
yq1NxQ8FWAvLyqiwF2MvyQ07wD8mP78rkdCY+3GGC3xTYNrnA9ewvW6r5XbleEN7
73m4ZT3J9Q6uxq0KfXGguXZA646LGZw9vUbYHL8W7PjPK9i4YPMInvWKb4VKW0Jq
EoUsfYlIomMuWw33/uzpkefcdB55LZKWfIGrd6AVo45kI2yIYXVLG1T+T8hld6hs
lCJFApqu4u2RhSfDWPeKhRmCUswFMg4X6FdeQRp8G55lb+KJrfnPexCGzjwUS4YV
Kuz2Nsc8k6iIdBg9iAPjIwmRAgsnLKNSFO9msGf6e+4hlcWNL+8Z4HY/zW0u4Um+
b732wRa6uMxdT2IJ1ae5tgQVvAEsGXIPgQDrow29WmgzZU5WV/C3XbUct4fWqd9e
oqDk9TYiUQ95jqt4p1lLmHayC+825VBQxddyLLYRC5E=
`protect END_PROTECTED
