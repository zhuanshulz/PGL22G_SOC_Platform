`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GqBc/Ii6nEgcFH143cKn+RFgEI1XXVDaO9uHXoM/M1acKLUQC/ed0BvtJ++Tyjb+
LtDisX4ajxt/+VAagIR2O/Eai8Vt8s+ZhTxxIVlXWnl4QFBjSIBMV0OOz4+Ava+5
Ps1vGo4wBLqR96yYevJtl+OVrUXmKezVmztitsVv9sR/ljEYr42kVg4UPRDCQ6tb
8Rs/4cOtE5Pdn1+EHL3GHTEVLXLdvKKF9DDcGiplDycu0utlyMFrgJph+Zsux+x/
BjfD+iDn4DCvQ6Cywyde4PGlOiPnY6I/QCuh2h/vGufTMw1u/fuCga2r94zMuS4c
QUOGSH8+wQC/gU/zfBx9hwQGX3iDMKfZe30THcUViVZBv6PpV3UG5fztd8AhGYml
pOxmFU4EQ8K8VOpMfZN947QuiFNBN7o2jFDFLSxGmiyMKlHc0aVUvJtWfunSH+BG
LUiY+SytVaE8i4esXJwWBn3hQFmliwgwvkkFevr7aGiDYKWx/+L+E+p8GU4AywGP
j1VRlcPLihys2wgxBl2ecrCaf5rhkuiTb1+0QDKp840nhv7BrsjdDc9iMtmORz/h
cFe7VLtBRMi+zbLN80bu4XRV73a/UE/eWusPpkeXjuriY1tH6cBaZYJOWmueHWFl
lBExmaXZx1Hq2wZj1Q15oA==
`protect END_PROTECTED
