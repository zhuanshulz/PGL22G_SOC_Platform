`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VbUf8prfaubjJRqXKp/yE2UIBZY4MiGZhutPSmvvROUa3uTJuEz+6DFWwV2Tag4F
mmfUo/UdBJo85YnDoUh0W6Yzylno1JkRJqoAIsVLywD8UxqFlyxGsXeofa7xqNN7
en8JAoS/OMuBJ0CqfZBMNsVFVSe/c6MFkED+NGfxRd+YUUCup5D+Gm+5AFX7DGMI
AlKQMTKmZOPLyY3JJ4oxddKHne/uO2TXX7T6fQ0q3ICN0fcqk+r+/kmZRnMoyWAW
30tbUK7g2vjEO85PkTusPfQKL1tSKBP3wx2h39OeWONksWNQeWS5HnocDOCV6Mda
3LfC7IB0c0xeWe9RJF+rMlfe77db1lTAAySi1hG6eQQaRD2GNtWNTwY8ndL5kclX
pMnDhs1qckOezqW24/nS++YsJ4NgesMLPUGChtHoTvUA2bYhcr8KE2YXBhZLyAUi
XuZUahUdfbNYp/rJwereNAUWGyr53zy3/sxscjrZoh1oZQk4Eb0IB0vBR8cTCWMS
p5gMvhpJmyTy3QDDG8haKtvaSbX8Qh5io2O2wk26p4ncVW1aOMiLUoXLf/bVIELa
Z0UcOm2ML9YW4vdbwoWsFGv7UNpkCXNKzHYNMaRPoVE+DEQ8m5rN8v5l/18HtymC
irSz5yHqHZEXGsyhg/8Y0nKDdgaBOEER9HSC3aow9wKlyLNOUcJXOAUfadMu7vln
bPU101aYtQwVQX+ICmaNuXK7kDdmScfAWSdFM+Tx7iHs2Ezd6pc3xz6UxMD2c3/Q
o4GgAMbTznxSbx4W+ZljbJKqw++MEAnMtMupKTRsIj1DG9j9SGxJHF+UsARTYJie
BWikJhJbuTEvuNkdxi8olajkTCqVG/lfefzd+1UDUKK68ODVFVr+YEcRWOPAK7dk
IJhmRPGq14nEKw9lvay/j0EsDVCdtilnrfNDFmaD14E=
`protect END_PROTECTED
