`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cxvIzUm2f/YPEnh1SgBE7IfKhpHlEVUpEJ4HCHML4EA1RTsZBVhDMeGdz8idMgZR
5lVsI0W97OGxf/RJ9tc3Z9mFk7Gm60xpEfW8VSbLpO3oAFwKdv5z9SfseQGdV4SF
Qs9HbLtBv7CCzl5UfOaVqqyjUX9NyztwUtWLZ9bcxBT14CxnaL9xNUVErnQHpI7+
cUMSNfJUN1HMrVQiJ6zq/QCaFTR/8UcCA0aIg1rPusNb4UM7kL7H9DosfwOeQDb3
nm5Z0Khz146wNM2nNAh+Trzaz9HlR/0lQhUGC02UfzirC6X+9/+SH9uJs5CKC3uL
t0Log90xv24zqtDvvQpCj8hErFxfc5riDyBTEpd5nwgc9FXh9y08pgQOMGnDbR0Z
HE9acCJS8A+Ccq5fqbH2cDgO7vXbkvg5iYrxn9qMfZgv6U6WXKZUTpmNMATb95Jw
vHx/i1o6md7sZlsGGh0GrXsIBxImIND8r1XYhbtdL8BC98aVoSWZGwb3OO8Hkclm
09I3hQWPNwkhKQUiWar7fpFpxVNa58esw1qGz4LBnGeOFDH2nXEAZwg4NB70KdZE
F7W+f3yUMToWwBhClNA2qzOYkZ8lFSitwg6XZGRjUWLBk0QMpWg5vV4tICKIuV7Z
YYSTyyBA+Hu+dEOeQSbSYNDftDjiFt11l89UTZDag8bU6ZsqYoLc99d9bRXOaKHy
zUC89KlK2JhBp0XGOs+ZOI3o2zszc5s5bPx8oOmgZ2QdZiLK80hAxv5tskNGGyUh
`protect END_PROTECTED
