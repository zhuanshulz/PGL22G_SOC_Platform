`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vqfpjRS1PWXmwMZSGlWDbtXJkgJ8kgHSalAumdsSm5Y6d575F/6U+iBYDQbeP17E
nCZ4A7XLOaoEBwi99uehPM9CLdnhaUU9jBhpRoMQowXSGUtFYv8Mp2Kmc6Qz8iPQ
gSweXKpmNq8WnR+KmY9DK11jnY6zexOLc0kDkBRmE0LBpdF/g3/5QpOWVPe4ZTRu
d2tSDNupZHNGDvW+U2dgjCdxQZx5KmDrR0vcXS4iHMSh6JeF+DVV41mYg2R39ImB
cgoL0NyK8Dz4NsGivtxOzPZ8d7u1TuxFs2wbZM9WFpwE+0nqzHQl3TDCagkem/mc
NIH0oRaUHXnmlNS7nqr1hFhb7kwZY+huCRssbiZMUL8al+YhUtILTE3OGYB/0wJW
PmIzVF3wM5I7eV2/t3Slx2LGKvGmFBdBB3VwT+nnZENQ3ObjAvwAwB1MbZr/3hOw
nYTHUOi4Yo55+ARlz/kdASEgVuh2kA0RydbM5ozDf8dJkEUbKsKvcIIYj8HtOMM7
Bd2Sw+anVboe/AQSMJzbCEHYpueDl2lzK6UmSmByRR9LHyfdfrPaqilOy0nix2yf
hqIEIpDU7yU02Sazoho7W65KCmu8UjMoJESlCdlM3MWbzq0WrgGPE6e3ldu73kfL
EKZCNmu3mNo+eNtaDHoeEpMeSnNYdZC5zdaFLZJODOfikISaaMqtFJKCbePJ8beb
GRW6FXuvAWbG3XEupqFUtDG07vIyMOeDI7qO2cHWAFFbdHW2IFPctNTUJsa8G8tS
YAlrvHO/nOOOMtvV0v8pRhup9/WPIjHL1v4G7vR1ujccQqgV3cqNV2lXZIRCKb8D
/FEeYODSGX9JKkJjr4Y3FXDD59+z8uULHxekoRLrFTuQeCG0SkzFYUgujADehUVQ
FBWpoktr4f/MxPUBDpckWudNXTc4pyleH3jmnUOLTfsX21ZIfP71Vrs84Z2BT7Os
+f8+hxUfRsDoBkwxZ9nnwXsrFp1HDxv2NzphRXum9+EW7tRdsfhfUZGEC0bOsBVe
glroz6J2wpjmwCd4gqSlboy50Xqdj4t0lhg0LeKilnZjSXpGtVvgHp0iP4nmNVzQ
g6IwTVAzNNeV7N1Oly0KIY8nDtwiUsUNzAM0OL8RKNLGmEhto2W0xVG0w3s60YIb
Xo9cCSOvoUfh7QTls10gdrcDlTOAfY88Gkye0wPEBe/oAXkYNeyCvAOurLsiW2Px
adQ7HQmxpSlPazECD1YJ5H5g7/Fr5nzyHH7jTCyPLthGweVDYODIwzdoZVHrb1Ca
EvIKDCbTUEFA81ASXIzVMuLY7jXVgDvgenumMzM9FWVQ2k39BLtKfrzcdOFxGaQs
6zT6R+mmaV97GVxCKx0+QRCwCnp5cEFfWsIXM7kyolT3Qb8fB6Hq4xTLIvLVk1BO
STRiwGiWtuA4E4l25SPOd0NlZAtc6F/Xr2tPvgIOvZ8EdRaQHMPpOGFqhKCg5OXp
7/rwABCvuKZwNeeKFI1uigk0/SIQJa8GJX3Y+kaje/Wmuo+3LoyVVMv/hCCStKpr
qFbKttaUxzz4sBNyFQXm4/C3SyUrcz8bXpl/iEuMLeY/UqFD1prOpY8B2g8DkwQk
7JVb4Zp7+GHlJvErsU0nv3UBIZ+SiiZ2pXkXs1RHk8BNilE/XksWo/JwAYKZtoyI
90kM+/F/y43pU4NAHDKvl62VCpZVYHCzHoNyl3IYClyB8i7DP+9RDz0Lqov02Aj/
47OO1w1+a8J+xabGMXYejM06hxgfQVoCb70wKoHY3UrDkb3uoUa0kuKlaVLg0Xsi
mgIWawX48WOyafLpbU6w5d+mx+Df9pSoUgqp/u7E5Zi64/8fnAU8p2o12VQqBX26
Tv8Lq+2sFhiMb5l7AeFrjKXP1fwhpQ2t+npalGAdd4/wnmu72CyGveXsHQn/3d79
4kHxm2eRJrS4bv6CxskOODIYRbrxP+MDtKHAL0HvhVVm7WTCCYnGih2GBfM0ujPQ
Zxu7qxtgbGEUsLoC0fMSP1IdqmG9ScQsfVwBV2Yb0By5z+XruAINRff/Drl4iTl+
0xFNWCy/RgQUMm4L+Ck9A6DP6ebhwcedEI7+bOyC/IVkBiOEovbgvES4gfadKWTN
/LUNduV5MdIeFwMLlHd2cILp6CdudaWVm+7aHJZLab5k6Ltw3FruayiDXhpZXJA7
UanHnlss0Qds6YVLRy/YP2FahZA/qPLiuE+aOfeEaPOv1Sx4wzMJmA6sg2a/68jI
ANklIqKqCMpWSEAWcoRQJ9z/a8G3iijcXg8c9zkAZTkoSffZzbndi7GxaKIKRBEc
+g6H/4cs+XFJjNzMsVSoqSKjePLMwIcrZEi1VhmLAhB3BoUIvajrByiz/cyQWtTk
/uJD44cufQXfwiuypki8jVlZ/XMGtxzICgS55Vq2WZiE50TChDwBxA2JxjlCMAgR
/iVw+5a6+m5YosIxvelFC93lFQ4b+2xi9I58DEW6wr9TmHzeQBkC3SzArIh0g7WD
4B6/godveJ00Wm8AodjyLZL0ElJrcrZPHY6hQNvUkjnbcW77fDOQyQ4xG55EobHc
iEmQjFr8MzwEot+SmgfiQfxXJfDkifSEisIj3nJ33thM0dYAcTCRyomLkqGray9Q
qxvccmm75etYFCGEfhRYgguQ/3y7qr2fnKmK/ER6COsCxBUqDcYXs6HNvvVws88Y
E9VsKOvB5HxLAuPy5mbMIvtZpOqegxRWpiVGjOAF/8WGgzXaZF3v9Qrkae8wG6WW
BnaAaoD4iHelzBu+OAqv/fRZGiLSMBF58vvAa8q1fdAYOXW6qU6g+BHccZZXfKzM
Yi3vEmi6OAly4ue1VS8tn3q2dppNLZVXS1HuKJZ3e02YZwZsVLAG3gmest33eZYC
HpNH7OO3os6DqOCdV402liEVosxnbXQs1bWbmexxujWMSBT9cMIVKkEQY0baXzXi
9XwZPGZ7ac7V5BeMVKhuWTxL47Ig/gTVqAIyNqHnwLZIF+Xmi4dKurQ7AOxq/B3r
7Laa8Hocvf+F0KMRsxKZba9zUJ/aKxHxrMlEfz98IHjn35UT0t5H4LxpGLpyaTJ6
irHziDUJlm3TKP+/WmeaewxR+sm2y27HCWVth9N+/qIhG2/+4bWJPpQJCOKz/XXy
4D6/w11ooMUevCuEJPJnSCMMVlooJJ/sClIUL2H6TRQt7xGyIS3HKEtq/9XDGMdu
qeFwkYvbGK/slPm8N/ILY75g0Xpisy5aJQ7FoNPOk+PuervgXkrr2ssfOQagItU/
NMWqn7sPi6QbZ1UTdFEdV+nwGyTy4Leyxj/IitGseTSVpaXjXxTaLKbgMlKhxN1m
xZH3FukqAcIcLvXYCgemYZI/cgFl7SnDfeLtKMolcUc41pC2QqZndMkMH+NAKb0c
6z6evft50v/GMO4NtLuVUuymrYJLRqXm9f+MTGLud3HWISmMd0HDnMzeoeK70K/a
NqR6ZPB2lhbSo1oU7kMNDqVv+NlDONkJiceX60cBnUEBEWgYtKQq7Xlxq2DO+nVb
XvSVb+/fXQXTvppMDDlOQYuB1CkLTSHo2Qnyj0LnHFXi245PzpHVogN1XnN/gR3+
ggpM2okANxDOIVlS3f01Jd5zCwKtJyYL2aqCkuscWrGcKk0StjlsJBvLFTxgOHO/
JrHzpN+2MKAN5gsFobsIIyb5LILyrUIaeuVWarPl3yRpcHusyUm4/giTO/sr0I3w
aq87UlRXJA8Ej1sbEBA7u/lqhpVBC7pcSj6430CCiZgXsgqSPEPJQOgpv+Vlkc2G
86cF1c4nufspjtPBKYHLCk+OdnRIDz7fXs3MUQtoSmK4KqPAM4yJlpvhOT679T9s
lFcq1DLDPTio4J/IMR9T80iA83YgHrxxP3PH7/fBRuelR3z6EKNabGYNSG5cLusa
0UtsYJlnrOId4oujGIZ3gVoLcsmWO76Ac+l1ogMzlneKFlc62c89ibdnRJ19dOwN
zW2wM/iJGTBYYmawedQunWci3a9oXsChxfvjK89cQIU3VsdaJU4oiMn9rHySnSGr
y1CI5MGyH0+2xLgpDXz4av4B57IvzNQLzGqYXyTeuIW5pCMvQcE20s4Cec3pBOF0
LezGacM6KKCpt/T8+fzv5V/Oeuory/I7M534moh+EjCSQ8Wj9/tOatSW8xrO+yo0
HHAnTtmGCPWXWAvA/yt9Fk5HZe2/LJwEdy2d2DkY6cclNbTvZWArDDa3VBq4C/FW
oXTnXVXPpEE+e04naPh/52cFEIeA9y3PqgJAlInqXyz0i9qT8UVl39qvn7E3iFTY
jX8jfk3rrOEdmoAOiYEssW3s2VSFsz5s5l3iEfj8C0mi634iZxnamfznakUCjtx/
bi57Nqc+EqUhGwWC7Z86YCPbZwEfpJF2LZoiOOj+Ric1dpvsJVh0GS9zBjvd1RWN
AaC6K5rA6c9j4wJ8CHald2nfP/0r/zLs4z4DfY75ubShyHRlakN2ps1TGBI1imun
Hh7OIq6l7/aeaqIJ0Qd69dkHygDAVEqRFGxihHy3AqdDYYNmTaebfWUYqlrgg6Wo
zMtWv8JT/MzsRie8X3/AyWdWMK8GR6BrfX8sOXZqt7SHTWOjeDTOqazeU0lznbl8
DdMyKFIVYHltNYpftntp7o365xfjzMC84SudX2haDhC4TDJgIdJDdjOtE1mZRncO
Lo7F46irt2c9f7cET3di4y3M3RUzlXYJVKlbbxX9gOwysibMsrG0g/6rC6ScKFCt
y6Jcjgb7MCzdQadn3nnM5sXTacZjLfkQEkE+w/xu7x0ym4gExtrxYRzlEo4jOUdc
QgwbcGPAqyZ40oIDtdLf5+DPzZI9Jq9Q3n4+Q13XFlAZZJ+hsO4tbFl93aWrp9MD
lgrwrYQPmKtl0YvQk6wX5dR6zwO66nkyPJFbQGGs3qq5TD/5JN9Fi8GuRnyaEq6z
ByA6CxpyZuuQnwuxGIPiZHqfooBea40Ru7BdfNfGSHhkByxWwqTKAWx1SLic9OQ9
mnDsaH5m/eCjxtPMV9sqjNny8Auor93BR13OUCFmT1X94MRffTnyQdRofdDNtmkg
4JnTA2BIeHHpVLCrtY7MsCXDeOMbwvC43VD/z+hH0N2NELBjqCM1euBpS8TNqJAZ
QVQrOovJsA/ABBnrPdp/AVWg6A8T4STPP0Ln9xSfISvk9zBoGT4f4ci2QCSSw9In
UIB8wIRMl9Ie19RDIPeyIKkFpKiz803mLwOuzRlbRJ/FcIhVxAhfOfXuU2z0uDSp
sogQIaQhEsymx3+N2Kq2aYV3SwRKKSUprYwNpfrJ8AvlDZfIUr3K/+H7gWIEurpP
YC2Vg6suzuW01uuGsqMQgcrb33TBNmqGLXSre/NKpDasHwJDAG0wQzSlfhXCtTDD
WvB7IhYM3QIgM5A/L1G16W/URRJxjBVEwz2KLxVZxdjSscpaHE4tyRFChOPElZRk
KgFpDKX/Cn8BYo6Ao4a6TNTKBrW/o/mxKHVAGYxMG3NOKRUf1ASRjvwDoWj3tJcK
V5y9fKbdMYrxiuwkqcN6HgaZRkH0EId1AP5zn1RLaYRAIOlq4MEJlg/eMCkOXhDP
1oQqxN/f8zweGNXDtsgT8cD6UU8X2t1skTdi5Q3r/23XnrDAvGwNUlz2k/J6Jd5v
ICDvceG/9+UX2uYS0Ay39giGBhoMutlgvwvHaCfaYoFu5XiUa1M7TmAhwXvLtgVx
27u1dXbI935bqF4jaaUCZSeiUa8Lf+L2jJmv735yvZgH/v2xJUFl57ybMtMBagCe
gvL8qMq+HvDsOQ7rJ9QP4wC/zpD9tjEyHxxb3SyD037NgohaIy/diYo5I9YbntsS
bLboVNiWju+2dOCUlJ0/ISSKdsfLijulkFmZnP2DkDyT1OkinZA2l0qA7gsOwUuT
wMeugtBFjCt22awoMuQ/7ehj4TLI7fZ0Z2Rc+PxluholElOk9emcQEZA/XXgRevN
xoSgTPVnmXtFEAKdgUjvJkbaob6MLT06a7H3PbmlxJ9mpUH/gfdUmd3rWCUXNFWI
Qd4BMpEyI51lSDMwZW2XoV2r5pTkQqZlky/CM5k7t7RuQA3tjyH4KVuV99DC6yB0
7w6WdJvxJqLopufLBZ0MQV8BG/rrblZgS2JnZkK9c+MxroH9+0ke2Tb1bLG5Sy/Z
09U2/fOl1KTqK0C9VX8CjMISxYmxud26iTP/2b0JfdIvnF8SCXyG9lb5Yn08UAyt
aL28xQXh2eoK6vmtdkmyoU7LapdW+ymzIHII5/4OA1ZjQQcVAPssCMxkWn9bhjqF
gmFqkH5g/CXAjGOWRfmdxznLZTnSkWKfCL4X7FexHW7V79XRWlBUJiCLHmEh/BRW
RyxKmnsHq+7HXGsjIHAaNSZODBVSDFhkclyM1rOnGxSON1wwGl4GG/grX1VJgbYD
aIuOIcnbtMgQaoNBVNwxSXjKC+d5r3Vj36LuAzTpyVS1WB07dEIaBg5wLIDyJ2PU
2MvvsPGsgEYSvj06PzEwgKjPdN7kDlkzhraJO1ixUcM+YHQltke8ZzmWKX5NZIZY
wo2p/XkJ2TXMARiWGk98mn0/qZp/WBx7Lu98qXgEEh/L/hHtSvxLCZ4BqyULcmJb
YHX06EnfTSBi2SOuYCQeVaH3GDFZI9hLLG4RdSljHRBV1Bh6io+LoevaZIKZ8gYY
Vp3zy+auzVXM1gaEcMca1ut/hehO95i31k9RTGCbT+DY8Mjeu2NXPkxRNRxVtXD+
i5vHavr86ZUWFelu4naro5K3TaBxVtKrUFvJpMFMQZLC8Nf+zGaZ0mwlJC1N5Qdo
GzPCOw27zoC4U7Nvo9/eC2GMbJLYu5TU+oGDgYIzbhpHC+5gTgc8AOqEyg4d4DVV
5+YCqkBusEnQyKN8qFC1J3/cWBYNFif//k1kq2CNCeKkcpF3P6ZCA0uPdZPy7fjf
lOjZ7QGdK6+AYpcV2XFFiyNHZ+bIxzwLbbQkgDJ8CvkviZ/sR804BgARu98xTUi3
D0diLTToBNtdbJXDUqKkz277edQWfhmD8/fw6QkRdOY/oUiFKkdGDzTRCIWV+ghR
XjpBlz9aabj5IPiULK8KGgTCgOr/mh+Wpw5gfnnSZW7ovHUnCXdDMj3zE7xgSFz+
HFCU1LrHbz13H8+sy++RgQ2sHwLQZaUjq56HBo9gOhlwD2ssVzbZwinm5Iyd9p9Y
aDUpLqbB65qOAFFPYS5wPENT/d11a3BBkfPSE/HVAB1KhvxuR3jwUCokO3o8xZ8P
Vr6A46fUE2wb7IFzsxb5im6PTXXhCSaGlfLBrPUUo0LGHrSV2BLhAu3AT4T0nT+s
jZ9Bvk64pgEe09RUvWQFNDeL/TzXWAcIZAocUv4KSt4x/5Ery66n+gXAWL/2scDq
YPGihfTYvxLKZw0XJbMsZLSZ2vOOHxB0y7r2HPbHtHwn2U5CpNXHMzeicZ/M5jle
YPn4IfgO02NQH/+AtBFkMWADXOEfOONz+fAQdJKYVzeJoovc1LtKqjGTUF+p7agc
bkDqK3kNYx3iwcZT5UBqYPJgCL2VsM6FWt9c2P/dOQaYTF96Kq7mBRkx7SkDYBUF
sTElEmmS3MWZxnXw8oosO6JlGDJ76HdG+6okYxLCxtuuRpBFJe8DQ4nE/bxTgY+A
nopHT0T6DtnZ+7xXFVki4d+x+DOupfEqvmDPRPz/6xWe4FmQBaBbvLG1CIEyrydr
Mdn8/hA29KUzSW8qtMCZPDFd3slexTpK8cjw4mDmyhyKRaEszaT3jHiCr/ZvSIr3
Y7OvpwIY58imY1FDomO43SL0tjHywzJmtD5FnuGr6JOg4RR4ADaXGLweubGr4qH6
x8FuYAwWCB9ALPSNz/1Z9N0AgniWE/eqQlaGnGkYXnxvVB7vJBGQDW0IcOPx1Drv
GfLsO6AnMVbQXhrSzC3Xg1axnozOgIZNRrQ9DfiNd0SVcIpsM+g/WxqXaGLfLDqn
nPKPToBJwcn5Sewgkjn8fIMDy2tvyPcsKoeW7Jcetmu/CkX97UXKkSOF0weCf79/
79ZO/btVJOV9/CMW/QEOSIKelAyacDk7H4tDaxbjUX/MUWFEGGHXpuIjSR09P7Du
+dg4o4Aqjzx/TZJ0xHPPXDW3VHcRBtOwPgaLEqTGuwWBY3HdCMn8Ui7ODkyIYhrL
UrjhLa+UBkGlRlPmnNEZMjqJTz0A89QPk2yof1mQYK4lGurHCo/hfJsPG0xUkzeC
Rc+fai2iH+eev6GSr7hVdM9FfXyfkFi56zWPy0mErpJbTwf3EaPNvUac51EalFlI
UoLqj7NK25C/Z/QYWnwcDFJqHz5SyBgnAXTigkRcNf9Lo2rC8yy5kxtXYYo9DzHQ
i9FZwwlCLcX6MqTqFg4IBYFNFY17RpZRrt7s/9V637vlVx+Q98xSGXEfUCqfbGFD
8gxBXftpZWVrgMba3J8kEhOUoEzG1aEirsLRsj94jur17FDxugt/tRwRDVVfqy2h
UwD8BODYES3vElLwp9aNXBtkZkm881g+Xs28tuxaZQ3LV5OGFepmxPDd9UMcj2su
G9xmPJ8GkuYUMcesPY0G8LhPGHheoqwkqHr1mRNu2WM=
`protect END_PROTECTED
