`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g/qaxSLJ/jXTttLsex56bGrhGfHLkpJKd/FwAWr6VmJ312ip96SPSAkIoRG3jWb5
yEsQ8UpOqq8EgI8Xb8rktpUMlmQejuUQbHljL/K/19BrhXEmahLXwLSAOnVMYb7f
c2ljsywzrN2cu8yZ+K0Kg/1+91jtGHIKb3EWBZOpSa6mo5cCaYx3ZbADwc1f3TvY
PSvV+vOrtf97Bc/d00mFp25E9m33mkBV5gKRcM94khVdOir/kyK8wuOxNyLJAWQe
Uyop6Pc0Y6EaO5iw14btOrE7HDzPtSqZMM6+oB45j5nl3JpslZryjxxNzDCYzGG0
2qEVTKdDt+FEGE/aNs7WmDI1ASsUwOnQso6WeuLvm54d/jnFCkV1qZxDHaQNgrug
ULGICInJFEacc4Wx5eC4JT5JJVCXbMinRdvlnpsEtUB6s5AY3b/v+ByQpd2fnGhq
1NvYPknTMPMrzwaaXw5112cPehPq5c2Bcm8dQ7eWGkBXDa4cSgJB7aRs4Ug0kqHt
x18DYqV9LUiz/CcbWg72COqHHR4uESJ7AHLucOEZyUwqXtvkyG+oqP3q362+Ajj0
/ISuTTyrMrlUfnIFMLITuKCldPcnMmRVw3n99K/zVR6S7nl6JykTfDTuX5752gcT
7ahcbPFcdyjy40pB25DBN2eg6+Xp79aRsF8IbkX9nowyZVYuFcKnUYBbevUkBsFX
TUoxfonOFwS7I6PYVp4GE7n8Ai+mM8x8VIwSsGNLhFZ/6NjbLTYnEc6aVU/iQa8n
2UheN0csPzwp7aDGNXHT0bBMOigeMaEGjjAEctAmPPf+oUr+M9CPtnKgCy+Ouccw
XdsbXkSQkLzUU/e14dOxZakV4mNKZcMyjxjHbIJqyorAvzykskDmxlooP4PDYo8s
fZ+YVgVuw3duQkAP40QSTTdAn8gcjT0o9EMumjF/udL/QzvTLd44JqBk3RGNpURE
49Rznf0vHYandhyKpMbW5PjujFE2GKV4bzU7Hn918Wz/SQg9PFm8P9yWKQrcIDWP
aHMNOXNTL5B91ATerQDPgcO3+dBVrBiyVva5LvTQJKY=
`protect END_PROTECTED
