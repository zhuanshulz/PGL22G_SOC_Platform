`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2XVU9FeMsuqnWYdZ81xlA1UN1gX+WGxAyS6GT5FQa1CHhVYEQ/OBoMGKSlpxR3uj
ibcdBOq92RlYF95GUh6tl0dz/tsEqxeqkiktWBSHZhK3d7bPyqDb5pmRbGz5FudY
PQtdFDEjEuCMmLU6yT/i4HPB+OxnJgZvMlke+P2KWnbvUZ8dgjm883u5V9de4VBQ
Q4ekJCG09LSmN5rxPuqNI1iE0X8LjA2+4Fwm5KIvr3793qV79u6jMjg+UDjREzQl
bMi6FrgOJ79DzDczq4gwQx3X3X0kiFtf9EoMRn/6IKB3ncN20gH0qvILQf+JEOTu
nFZ3zaspFRVENUpiXD1ToqYfa27V09zsRe5VJD9/QIeC2DFSDPO/vLh90wJ14yIu
jWM2IwqkSR+w2qNsr8gyoyJkrwpdDUtq549fFxye7J6N6mWdFn6NDmxRojuZchMR
x1CqgRDxna0kMT9qeQW3ondb1Gk+y93cEH29it6f6+ysSJjZ57OVGpZwTVOZbrkS
LXPtrVoWl757BVzp8yMkNdeLvTv1HZ2eky1XyM4IqWVJrnqifivBo8d035ndq1Zc
Hm4eu30UvT0IiiFBVUX0yA5Y9JEpe2fkT1DvVjz4yWx0SBz1tRVUJRbfj1eugY5s
XUwZ1E/GtfuGURuStVmA6QLkiUddBh15K0Lo34F7rL3pOPlBDkP5Sy/eNu047g+Y
p65fbx262rSnHt5k4xqs1e5LXaGCa/ujaG0TVVKTotRRtJANfMA0ykF3i/a+k/74
FR+kueaaampNfTiypoc+cBWyaK/CVfstJJyQxnXqcYCKMdRLM/Y64uPOC7hmeaKe
vrFoyF3nWroUVwjSHj22yVtw9FQ6rcx9vPvTZnbL7owSdLI/tolQTqJ9hK8V3184
hh9TT/rQjnDoE21fHaTXssZbT3qtlPA1BTEHJBFAxcl91d+P/Mk0BETeTz9SCPVA
BnNWscSgqWEbx1NVcigqyqAaqcrJWLQC5xWWx+YATwc=
`protect END_PROTECTED
