`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dSx+DBmKqxL8HXGkdIUpLlKFh1y3zcV1vWoz9Sc/x+3mMp1SoijgILr3T1w+QmRL
xd9TGlpeP3bbni/Ifsr86g5GiRtchYw+RHKkBKreV1JuBFn4emvoQt+Gt6UNEXxJ
oaLXfHUnGV+QmH2ra4jibB14k8ds2r04RlB3OWNMaFLloXBUnhlkcVnQUNVJv3cw
z1dhZHD5UiMj4ibrCIzfzB4La+kFGK//sv4iTWk3u+7YZCDSma66PVqIYQT3w+HU
3HRq8kDBt3arvCjcJk7s6g9ShRveEXFPHKDxCJXXLJD+tDrcSYDuMZTWJhWxJTtF
nkagDLh26+2PdaebWJYf//xYeW/Tawib4SW5FT6WtXXjGszWxRkTPhcMUkziy5TZ
z+A3DwV2uE5z9L6xNjZNw7c7UC9JNFT33wMP+yrakwdGrUedqJ44UmOR6pk7AXU/
7qfPMR4hzOO2UvFaOMqeVtZeN/ZC74JA3qByGB/GjaNzmuOu02nBenlsitHSiVe5
YTUewOQPrn9DUd4qdbLwEUESVGIoCfzpBNnBvZtQE8DtPafbpmO25uCK2/JeeKC6
JRtfyD3k5tvfwdUdhkOFkNCmWwDBr9YBnF84Z0PAaRpWXqmEI2eGMEsLPiRtQdk0
1r3/r7KPkXr9LWMnUrs/ut7ZmIPaAhJwyuwKLDQRq0rAOJcPEXmKW0JEK1ar/qE9
Z2kSJWRTI3Ssa0tVXN7HcwrSjC0AU+dX0I0jj1AKyNU1v18GtzBVC2EQTbfxKie/
sMvl9ScZyt19xWgz+e31eL2qQ0GpK1vUOKA6y8ChylfkK5IBm6M23cZL33g1o0Vz
AUw0M/JVuVDATy/z28doCwHaUnjrYqx1z0ONZfoZEixjSsHUtRw7vwLPTZUbbdKy
kL1tSx+zhoSd3bZEPyc2pjjUvLvYZXTN0IBe10ES98wtJGGwDoivFQVtlKLCAClc
v3pfk+ciTtKIyJlkd0IvCQOT2LqZ3MQbK8/uGRQHFcEdlc60NMMp9ysQhfiggmwO
TGSlpvq+JBhjiqWKAqsyOEw0O3oUE6JXZ1JReAfDdWUN99iPFlp/kIerrS5wcnx+
nsgNWqr0VeGNBgUm4m8OKrnyFv7t+PVYuNU5EXb6yk9Umn+1GEoueOQDcSI5z/FB
e9uluYcw4c9Rk8Si1GkI1myjBoMw9wlhHa5Pqrdn4oJgDR63OQwavE/PDmRpT39A
Dnil7lWK4ZjPt5yRhRGshpbLKs4ta7Gw2jUrcXmzc7oMt6jXe18avwfZbbFotP0a
SIr7THw9JBnEcEYPz0GLhUSpUJ85Yaoen127W4cEGuVroJxSuKE3CNSscKGaWxSe
0SGA7d/RAS69CMU90r0eI9gopCMNsehXDSbdYaNPFchwBVHSpTJsjrw0kOqqK1Tm
kE8aUY15FE8HeonCYW+btb76IZfl4EoBUVRNCQw3CsX8Ikcfy2mic3zxgAfIKHWT
pXod6iKCFFuN7Wfe7ZlzbPScNvwiw+AlSJceTaP8806ww3C4fU1q1swXeTvxl85r
F8ExgvZSyT5mmhqw5fMIu5GA7YmGor7x0vdH0poFRDSjje8fpMqUiusE5t5S/otl
ZIqAdLSK85udgBQxSiwZkanAdQYLN+evpytvBOFYkAFpq2yhZD83N6v/iXt6kqYm
It18xUsqVrYtyRpkg3Yz5wP0RZcQ+s+QgJsvSN/VPrqV1768cO/+4ox825/EVvCF
c1ST8l33DG49ElQmQcOgBfOs++FWcYymB8t+AZm09WToJ4VeQwds8Y61sqg+Lg0n
HiHQqP7EhHhD1zjU/ZwEnBJ6h1ypKWhig7bf5/aCaNehdZz2ES8R2ujkFBJTirFN
PQRV7xVr3q6peu29uWtBkZAVTX6Vr24p891bFYYuwIlC7PNyh5BJ+sdaVgrzrJK9
ZN7KFk99Uhp00vIlTYsTInQwtkoOG0zfDjemilH6E2OJmIz1Lqy2ZdBIrXbBdIUH
AYAEeK+6MVexcDUHSMvRH/la5AJQo8KX10NFpKxzdZu5+HhA+3tfyhWZCBE1IEMM
l6FcHuxZWGE9zu1J0hAelpVDKkNkJ3Ug01IB3jMsC/WmtMgQcfNDGiEPjLBkbysV
Eue25dWz4f0Rqx0mE+ygBNvntF6gWsySEuwBwMwxjI+JK42/OQ/lyO0NagladnaQ
8iPajI9AsR/bXYqJpszvEmk0vKSKV/lpV4AI9FHOJR77OmhLozKpCTUtucYQ+0x/
9p12m+KXQgCpeJP0p9k1n//itvg302aQ0LC0luhUOxaWjILOg14psgkw7x4L6hBm
W7kPnRpL/X5Yt7IwyBQH4FB1Se0BR8L2f+BBuFD2YXXOXocnrluw6Ca5JHcdCu0n
8FzU4rZdOlD7OV/ZQX5e43/poZ0OLckJpQST1q5yQ3fx3C8zkxrVh5ry5gjViLhd
1Wm9fwq2B011gRO7dJyEaslHQZsmf5P0ZeF2R8Yd9QsoYYg3hd0u8yiZBep4T7nT
0hkhK6Jg+GQWV3GwGKkCJFZ9WAgFlznRIoPm7Y0V/2slvHUpxlMtcPokvreBagJx
a+dNgMeNMwAJKmayD6Pi+ZYGLGtcRfcoUl8UYHJRBbH5EiF5dhVSQWsZri+yT7s7
uqwcRQZB8vUKQN1D8OnLAoq0C9/3VKzBsjR6ot2qiPRepxV+ilvitTMH97PD20l3
QF+M6aCBc7jX/PMiLfmxLIFQZAMOFz514sr2JlnNc4LcngvBZjDWPq37DfOs4bFZ
o+g4thr2KPWyFiUDTzsShEyxl+bJ6/RpJfe6M7IdeB0+0p9/VyyV2uMVOa8hOjpJ
JtHkqijfa2K6Q7TMq+wgqAJCd0K2at/yMxqHVVr3gKudl0uj7lfpyTcOeCURJH3p
We0jduF2WVj76mvwGIgxPNkj7WM7JKQpp65xhLlotYpRJ81okPoaLD/yWt3KOx3u
b3m4GwMyWMFqizl9ZeSWkB60qmfvg12xwJTmHLcM3EdE6O+GebnWJ4W2+D8hPQMP
4YISbFxH94rp9ed6TLHqlNS7b18yvBsQ6bDEVF6Kivjhl0jpy9BH6DcPNGQ5mJwh
jOTpBLx93MVGRu+DpZTZ7Y1Lg/EEOw/YWw9tsigH9cJXWUw8my7JScGigHavO9iP
ulwF2dZVe7Sj+SY2omUVaXY++0KlqCMq5rqkMAyxLMBwPBmWBWAXB1V9M1xqsD0l
7HrApTKSmHWTeeVwzvuM3cJNOi3HGKGpm6uFd2yg40+MiomxWt74v1FPmjP6amz9
Oy8rZ1pjFqhWGQLD6hTKwE1Oe6U8mdrImcdhPGikN0GBfqgNgCGTtczs0+GM/th8
bw70K0F4ljuoVX4J8K1niKXTrnbV/bo8adAPkPvhWlgRIILh87V686AjPs0GfoT3
8LuVC07u1EA//Z56g9KzoGwX2aIJhulx8EhEcM9oAzxfztyPJWO4ux+727fNVU77
TzmFADWagGHyFhx+165pk8sCWgsFOEBR3twPJBYbVedUGjcfkfMlZnTpgycfy2fq
gW3EVF+oqCNJLZld5kHtcAw5FICMLg0rC4RN17y7UV/o7c8WeR4PEXk0wCObpGHw
YAQ3bkPkLZgsfMxg4NjHWupW1ZQb8AJKGTUHzDylJBTfBiJc+M0QzYNDrEgX0KUe
yZ640qzkyO9mmiWhkuSauDRxJXIITjVDmClTAjnqg3bUUo8cQ3gEoXiKfnFBgE5Z
n3UTmbLkp9vwFkMSkOV73YK1w9cXNt04DS7BpoJSL4nyVTb7YV9aHPxoDKOiirpS
P3bsI3tjUMA3Vo1AgD8ECaD+6bWfQzOT+HoVab6UqsoPB7GYVKTh1PMJiwEpL8DP
2jjl6PmcbNMctYb+KGI2zg==
`protect END_PROTECTED
