`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CUeUMj2TB4nhj8e9irKxs7Lr9gZ3E9ntjz1RCZT3fkNiZkAYdKvb/z9JR/jvaYo5
1C1/N4CNLbfrVmBfjkLK2UgPevMP1hQMMDYrSaCgA12xUVPbLIalJxhR2okEAONV
qXVaQZ7H8ymdffpxaDCQ/TD1MnN+CaSWrdt5mdkqSb7U+lW2io5XDKdXp9Tl8yez
OybBILvzcHeeP7fYhgKZOxDXk1mOIk3EyQQ/gQRBLxP43JpdLjymwduwAuclxCU3
/g9l5FJA/0bUMFhRVyYMcwnh22Fs1eRS/ApuSmRt6fWclL5qJNdjMWE9uC5kDrLh
YU+TLqyKerKQvBkmu6PuCbNA0/OPGBuuW9JhtNh/mesIr9ggzM8d6UpvgeD1IFqZ
DIHD0s/zn17s12DP4Tc1FkFisO8+BrpkxmgCpnf5Je0+V4a8FgBjXbnJIHsqVqeD
9mGeGdE24aPifM25Ca9qZ/T+FZto/SnwhUc1uiVFOMSfGGeaLmjGeA2EARJHiAUY
bdGFYR/+IvliAJ4zunlxXMtpZRc8dk+5jjapHkmSw7DDePHxqdkFw59+WJOeo2NK
OePr/mrGdoSEQyHZ3tZt+uSwLTqooblzC0D7+EflyPQP5cmT56wtdicLFdEDICDs
ECC6+f3WAGb1ZW4nSXDB4X2QRW6tejsbFqqigoK2/vYPPrUSdtRgkh6qKqLW43Hd
r8sW4+/DWSIzGRMAId6AmVLx19ZAkYTdRLPHkP1tb3LzQGJqvfGTbTMYqPe45Ger
MlR4Lm5ylN6jde0m5BUeLVa2cnQTvRz9JCpd6LH8uMpH1sy1676LoGwpjzx3adj6
b4pnrKB48FkodZSQrKbv158zCS4nRSjWfVc+F65Ux+44/TszpOgQQPn3AlvR4WKz
9KLpOB0eAIUn6aZPpyv8uIucJOUP67Z/3I8XqCsN71uM+wELYgf6lhyNYNH1AXPS
BnCAI+CkcviL+8e1Oeg1KYhgRrOHHRfUKqNL5lX/YS7vHm8/Y9X/ioGgluK6jSlV
/g3e84e3W7J6RnnZsltho5hdA1+c3H+emTtqsHDElMAdywc+sdAVO2fhv1hYfaLg
0FLcfs6ckTCzydaIT4wZp6LAlvfdTFQGLdOA52pzwBjcUQB2u5sUnWBfV/Zb4MSA
5sJ1oXsbIw1Q80CMYCaBS5zzoo5zBY90GQixCVjg7SuT7rH+R5IQgI1VSHppFzXA
H87I4yZUZ9uocBm6enmUcbV4uqs5lFZ7pn0BdlXpRMOHcfWsacy5dXv3w7hqMUGU
5re7jm+S3cEpMJFRdz2NMFqTMcxg/jYUhC/JhegIIzFsvSnEkJhkrmtcwAsNb4Is
TRt0G8l2Fo0Kpo+V9X4TtK1TUwwr3ebHhyfthjYEpky8nb4LKlB/gKMoiY3JxJ3W
e4D6xfjC/T1GaoX+1yIABdwW16W5e/psCjcRiQitpO4thL7D+A3R67mPGBK/BhWo
er0/PMvuvQVqVV9GL+j/4Ro/pNXTnI/ImWOrfsznEiff14N2YC7EBSy3NxoyccUy
B5YpP8XtRqZNUH2QxJbGDVdipcFXMtpxbtbLTzpeGRac4V4/TwOWznpRAuYPFCuS
eotIu+K4vBrMPBibW8CowpYorIiQ3D4nSFDeNTInUqLOcDWNs6kFHYiEgoQ92LH6
vs3AELD50fKP4rehKU84OAVoJuqgT65DMpcy/aII9g4iUYExaWGDB/bQQYrglvEI
Pqcq1f6HM53MTaXKbBVPO967H1wa4aOTgpSMyT/VjawL7C+ViBTbWpDYgGBOWjfU
erVEx63lI3yZ6R+mbQbiUc2WrpD6SeQfaVGBOT6tgAQ9ix8lttAE2Lo9oEkCY/Cm
V3X4gbHu7nShY4B8JLhHTcVruxPt8hni7heWCb2l11cKXOM+H95QNxlxpmGO+EdX
cvTqDDDOv//8gw+WQmukOsYxpbst2xtVYwERrZZny7eibJrhX+I+cXuR+WqXENBP
lT5/sIGCi6s3Mo6PvmzeBw8uaxhnFmSq15xh5nrHcp2DOsRHtfC7fgBzfy9dcdYf
CnaHgzV2KInf0Vk3fjpRU49chBrxGU6QgoX5SYgyZvT4taMaT1Yw+omhkOKJd7mL
bk2GdGf/zX3LHfkDPJosF2dESto/DZyoF3SiTmYsfHHoFbnBwKvBn+mBhMeYIOEt
iE0U446CIpe6peCQ2miduvwgXiH23cMtp1tGY8Oqkbxyr7Wqcy/dBCQ6HA1BZRoW
Q8po4al1qcyMNu1AmN0mzmugGa+aKDV/LBUgP/wIzMbevFK2gYua5fSMnqK3rsHc
NsX5IopWtnbCz5LYEnsDppmsejOKwNx0nqA7QbbF5luuVJ3XIIY2+CvGYa7VslFX
8p/ZxtVT//DPZlipaHKKQk+EcydwRfnREg/dWXfRTC6QZonEgOw0hUDR+64OZYIg
LtX6alMBSxD6zOe3KK1JTW4T0QvWrult/VCdBwBqI6b1k0vl2jg0E0p1WxfjrUEY
ps7d33NJxbJ5qEExZhYagWHulsVWufaiZkTCc8yu0ElQ+Lruca1lnxyhxQa8cW4b
oeRuSWZhniC+juwha9I9idEae+WxtmYdnBENSRwsd3ntBfmN6gYWPK+WZ9Y4iIaD
g/e55YkH6330r0K5NZahgwlzcQanW1hFPsiBzfVB0FvSNDFB5fddNwRdwiBnV28l
Bqdo7ZPO4oZBVb8hOTttMdvi40wRWevLgoWgWiEZbJitOj2Th/sEUZtj3tG1Ga3n
bVPl22IFjesY1lGWqaw2j0oV2pX78GIezNUMluqArMQIdMd44FgoLJjDixw706Xv
ibVAtcE/OU0UZKC2NAOzOjgM11nQtloFEMWKc2gpkYqpdHOkl7nz8yAGoShRymkQ
5kzJMPSo3qa17X4krM3jH3j/k8sFf4BkHd+Q1+QVLvTuhllPblZrTm2Uo6lZDL/J
K8ZZSdANLoUyBjNcoTXT+IcjJg2bGpLOpBAU6uEnPoqvxz8J7ifXUcK012vbMNHA
vsy7izU8gxBcOLEDanocFQ==
`protect END_PROTECTED
