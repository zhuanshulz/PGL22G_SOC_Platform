`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/I3r/RMfmck5T1EOYstNrVh6I5aKM6BCG0RKzyJ2P9tyDJvubIevKYvoMDwG85qS
adOplzqiWJh5LrcCT4A4NG9bFLg6vUlJuY3EG53PAED5RwMYM47bfxGMARpkpICd
rFuQJgFtPpTsbm3j6pPoIvkRD9Cn4eQccwc720Z8XsoBo9OZeeNUhaGUlTPthp3t
B2X0eHkjgGRM8m1VzSH5lVPlkB8E0i7h9hw9+MbHPMLRMAKWhqwyqcX7VtCmLHoH
rTCPuryoP2Hma2DCA5TKdzSgmyTGzx0FfnNpQ2cqeXbmPwRT856obdPQlwdyBn3E
e6tIqsFNUJ8/HT3V0NOpEelMh+KxJlqIQsyhsp8g3IlluMKoeSxVatNzztI9lgU0
gBH4VfeieD6abiL/xpq5ebLDrrF0D7ATlGUkKfQdlETcbrrMgz9G1F+3breSvpWg
q/zTo9zl/tzPciktQeD0cj4im8xsvGKbqlVahzvPns0=
`protect END_PROTECTED
