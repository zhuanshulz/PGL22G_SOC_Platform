`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4NSWR5Gdr84ra11jiQQizRyFkOg8+JNKIjk0veyY34msQXaoNO3jWLKScEQr+r+x
5dCYQF3FrNPIrjjY7U5Wjf1klcqEc2voZgdKTe9F/gTztd9u6bGc4QF7xHujhzgO
TzbEOVXBdAPcrb7PmD0RuVl21jRXaKVajdFcRDzYiMxTXChAe0clAMslM0SW6BAV
wmLn5TLgcg/fbE+ujPuMfViRyB5qlentGricT9xRAK8af6Snq5tXB25fl5SJ3JYB
8xdvYHfvwDPBvEl5QfV0jZo4K/Ao7bHAfOpNttQHIkR9Pp9sTbhOtIXHhUg74Fdg
30qasDt73Ywb9UWvadYFCHqJAwu0qtlXxArqRk/wlgbNxcQUYCFK46Ib0xPYYPW1
1dRiLWA96YTtdSvY5E0eLkRkubhkJw6b2FAKLuUTu/YAL7yrbR4wtScq08KeB/+F
JcUGhEqfrZW5mzGZYWJ61qQ8It6SP/sERfWTXhkyLur1a0dX8+DNvcox87jhIbsd
XlOiuTajy8rNNswJD0vOxBbZ1CuiIXFLtuI9w0d0UF5X3oPz1l4NlV1QY/iAsoAd
NxDdmy0xoGpytMp58R2lue/IL024sySE4lviHacXf9ZL6dXZewU5b1QM6Tw7n2WW
UxdJu0AtOlYewFestnG1iukv9z/POcwA16fXJfXcDxbiBgVt31jZGi3kB0wDw9CV
m9kbfNATbZMYrolCxmkRzf9Vu1FLNj6vYbhCmLKyGFj52Nadc/7fikTx/PxSZ8WF
kVL8AeOh4bVrfhPvbpCqlQ==
`protect END_PROTECTED
