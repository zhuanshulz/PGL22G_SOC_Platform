`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MlCEWb8uogdMVInWaZjIjWGvevHqZbW6U8JHU2asyhJxH7iEEHIvMn6MCvfb/Go/
yg1O7OKcoPKLf8f/i87ZGRZy3p5KEYO3cKduz4dSYQ5UTZpsGkSExoE1X4SauY3Z
xuQAXfylOUiFrbTXJSzDp0Hw0LD+pq/qkQXvku328zrv0lowoeJo8m+Zvh/5q+yu
IFOLpg5+z/NV5jTKDnfRA+PzaNmMZyzln15rc7TfMnZsOjMbeSFj/bb6RIhcovVL
XF5Cuo8Xh+MGKsWJ/VWu73yrbQvvi64+9y3U6zy/TY5y8zC4E89syYdfM3CZ153K
UwL4V0I7J3tPznNNhi9oqCokb5t25P3of7aaxtlKHjW/QbWZH2fDkHeeXeaBpi5c
zD1pGLHxsO2EaxgPfVA/XUICJ97ElB5D9669lGoeaLRaiLeU4+AoE7MA0Mxa++Nv
9Ya8K1SCHs6VOHKsBvJKPH+QeqxhjSVzwkP+/5gXDj9/c9Ar7NOTpzFm9tK+hzkK
9ZtmC+5clwAdcgSC2K/FdR1p7yIYjlCBNvVZPKb9Ovrg5yTdPWXeTlPBLhaW9cHj
EpaDTkBC5irvd+DbmgIKLcVT+WqPBuYEFgtmfcRyD8Tjr2ftQD4JScNcuG7G1aJv
`protect END_PROTECTED
