`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3+l+cowq9OGSomjkK6J6NMgObfNNDNfOIHXDIYwmM8Oc0FCntOyMubYOM61d3DLQ
+VUuFWBL1vVmKOvXLdNBuBcYFymC77hnt3xytvc1EcNXHqefOlNHIVdYO4gNj3sk
KmYE+4pPMtGGwV/uNuLaqGvElWudh1sV1dS5Ol7yenm/6819+6Ez/YYDCISOYii6
v75QJb9Pfk91j6rTaopxBqE3pKNB7mjggiTr0XAUL4NlROsCbHOT65KE/dHNVGlC
Vzkm+Fh9GxZUI6gU94FnpxPf5OGWvoV/OUn0etp0Ii8/iRQUo56RvQ5FarF5uVoW
MAZaFgw7+FiSlX+NiOCdBqsOqjM4KOEy+xPqRi2k8d8=
`protect END_PROTECTED
