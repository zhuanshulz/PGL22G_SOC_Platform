`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dVQQ0LnCoBLehLeSpcynl65Tb7H9EXGEbUlHPvg8tSaNCiXoC66y0H2L2ulwSeNk
9VsNldXyefcBwXwWrKHVVU9VixudPDD8glqR0K4QkFlbsiiBfI87nIi4bjHrtEzo
02UodtnV+hI1kBlmtyXor7d2/5vEPFZiowE0JSOq1qU51t7tPXFE+vlIcIv/GqSc
vcacDqloGFANuKBERZ64vWgLtDAsUlsI+Yzin0bZTaX6hPBXhRnjDgG9hmmolHeg
KR/l81O+eSfwTakfb07TN3bnk7nvwJ2URHJ9xfBAJAw0+yuLU7n1FVarebKiUG80
9FF7Pm2dZ5UuRiMh+G9+cyh21ZwJwGy9278mZb70lSCV019a3aL2O5lpkHXsdRWL
VJyWFtLkQn+U1vFe+FqyGx3D++oePItjUoHoKT/swwmR3SYUIYU1g0DklmuFUdGo
nnec+i4wtlE7DoWAtzjIZJtgAZ3yZt74qV7baKl/t3mmedcyZ3CoZmmrGevHq7It
pb2SRJyf1F7O2hRqsA/9nLUz063d9673/tgcrqpv/KL1m/jQtlXvdM190XpnKUHK
iecr2E+OAtBH9Vk11JagqWUIedZVsdVW4mopMCr0021MPv6PC3iYM26HOOU21z6z
6OMN4PyaZlQ4EI/WRiSDeskaHfTeXhD+f7xFVcNfN9vOZFIXIWUgUULxdvdXihs8
Imcq259vXNNFhKzuDohTNF002EgLuwAf0sRe0mNpBJbHbcHbn35Y4IVs3YK15Shx
k9i9GZRSs+eG2hcuXSUlF/fYPd1Gi45OeuznYLQO9NuLMkf44KmUkhhYwh0gUC9x
HdMmCBu179197VlFW4lWsaWuryy70TFJkhttr/Z5h2AokArpjhHBTbJEYC+VSdJQ
dVwtq+6KXTOIZagMZm3P0AQDy9CQsRWAY00bJRs5Vd6Mmp5uQ9cERfbGYfX5Mcas
s2/9GJS9+pirtNEPanI2KF9EEnuEB/3kB16thrjMvNs=
`protect END_PROTECTED
