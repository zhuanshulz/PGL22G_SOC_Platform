`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U3hLKWUOCa3LMiGlVoeFIRvPJVFzLCvf0dH5C39IoRmpvikZJpL6Bd5nHfMiTNM6
14no4xs2EQ45EGUuj9zbcXMpiy1R/qLYAJ/tgoZbCq6b5IdgFy2ZLFCaAPWZmOVR
lDc7nF1tndvRZWb7+xUJ+iz+Cv8LAGnEOFinefUyC5YP0b07SpkFNvSXIlKfpiM+
jqI5B//IBqYqYncsvCwA7TtXU9Ir9qOfYJMXh6kbOya4/f7jqKdtdJFBwmdx07lv
Nl2ZPi7zb+/McfAX31EbDvwbgfWvHvRZH/3vlmQNstfqtbXgH3FXQjDmAPpJXdvE
ACUjSDlPp/mfb617HhXEpivq0/Cwf+8GKY4bTWM9lvY84WCf3uU9YOOoUV3veYo/
ub3skA7sFhf94eAfyCmzdWFLjVTwYR2raxG92iA4ZqV7AKvUpGVrUEcrmAFgRRgu
DePVI1b9mQqx+2ppTsCv6MCT2+TuMZ/y4YRLMEnw1tET4ieEeL3GoqSaDpTt4Gxw
HYhqMCLD6sRjWH20AbwCggx9kyuKsOlMCBCiDlZ+qBtVJP6X93tpmEPfxcFhQXGA
ZuC78LZLBt3NTGVdF6LVEBtIE8RvCWKhTe8OU9carYOVkDARZ3lHXZFG7cJO9kDP
CRj2uI6PbV/G1DLujp0oZ5gxv791HTWKulG1CCiXC4UfEJqjQUaKlQiShZfz/6le
kai24d2BU+Maa9KcGYvszZb8qLJ9HJTxJFGDWeH33zOOv7wEY7QrZms9zUZFqiDa
IEwcQCpK1mF2mZqUjQn0oHLjGt9i5WKQi2l37hx+xIchvBUm35DICBdF/Y0NcPoQ
r6v+uaXcbPo+JCOhHoIqKh+Sz0cdhtwojejj4oigmiWFl2Ol/ttLkGjVkP8ucVaa
Ke7AFOkpIg8w570186IH/GCJh8fXyD8jkk7y6+71Db0Fi8y7GrxF757qotzx/1KW
IojDPDUM7hMw7IMssscErCpagdNO0RfU1ECds/Hc/pKC0EuSkh0Le0Ln6N3doV0N
2NJvE6YSBzTTfLQQ5H1JJE1G9HUrCbI9LjDcyYgH8bDYkr/TqN8Owjv07lCjbNUP
6PrqZmoaxzyJiM6gqMrEcNnPzJJnPecfJNc45Osd1WvPRs95iAJ2+BLsFpXObrAb
YbeclHDvS6sh0l3yDWMDZoYukFQK7rBk9uzoTLpER7aKf87+eJR1ywQ+Wyy7BihG
9wqwvJCDpRqs+nEWjfp6ktXhe1/nNisoy/Kb4uAX+N/cSeimKiV5rpMHoi+P8fA5
eNQwXBn/P9oegUBf/lkMrnFSP3knfzbDs0E9cms2yYZ7mu9YIZhoD+o4OFhO4ae2
ilbutAe+KTJbCsGVG+H9W7aii9CPpKza+J6EKnJm83Io6O/pVe1TXF0h/cHRYj7m
Jf6Zbr4pkS3W1u0osW+QYi7g+IobI3WrwybMS3ZT0pSlNF8aslgY5jfx0X9pUGBv
sVxlZG71/YLB+OBSv5P9hANLRRQmRq40abf8aIjgoEYRntPvOBjFSLUwD+q5+RSj
E7aOMc9vQWXWsPi4caTsYYW0WkrqfsXrrjmp/NivDgUiHaBpMuTLlLAFNkTWvSE2
6sEKv3UNDltRBuZRuszd2YuVbU6Ksyj6zh9xO6xrtFOf1NZojVYyztxfpg1XRv1+
NDjSEQl4MMxhUVGYqcviwvPtKLEnvwaf+p+MCiiGQlLFqanyrT4M/597Oy0WI7pr
etDB61MQk9MJSi5dojppsrWJUVw7DCFaHpX6oSdmfhElN4JkEoq/d48XDgLNWjX9
vlrHBoxgN7JKQsD1pqNvcGDtFkQw08J3LWBRFGM33Gcaor/yruSWvHKfoNu/vbrp
urBs9Dy+gYu7flHursBNsQ0C59RVVdBB0KzFlNjvpX2oyt4WaNFaf1kDNkm8ulAW
SE0RtVqod8bgmi7s5E9N2yYDPKexLC/HHusGYLnZXBjHuggFpRnSWAicju8YacDf
SKhYjHEiHzDArZf2ko2lOFy3TgnC1RO2tpy6hwwQ4NZDG0hPJ/bnHxaQm+vEq5+i
PIWBpgYUWRjQZI3HWLuygzZHXJZAg+yXYzqsVX+D4y7t/NrEn3qQH9MmbMgdJ1TN
Qs7wzmQdAb3xQevVJDtbU63VwbiwuROzRXCWRixwgKHXGpAenyoqXxV7LpDteAbQ
BQVGXvIBSA36SoGhV3oUnhmRwAv4algAvrWKD5PHKnjelw9lgixTWY/x0eSUfgLF
89aN9HP6nFAcPV9Hve9/iJ/5j6hwOAqJSYsdwctRx+yHpMAXPMnBStpQu+RWHM8j
L+jO8pMoTkty911/bNMSVtc8oxAubSL6g/IhKKagvBEgN7nqNVt1CZ1hEYab1FZ0
RjTl3ume9ZhxCe1s52jrGIT4YVv+DizPInr2j+gm3TpfXtUPf3jqAVzLK/IVax10
rzEj4w7s3FpdSRaeCwylR+X86A1Za+DGuIxrqz8oUJ0n10hJEnACt0iJmvpsFkBu
4NY2AeJoqk6ARsbu96PLZ8NKH8pQLWCQ8hJyK4Oxl7ssciGykM9mM+gwnUcxII2U
2bVvPdjUGD0EOIf7qUCOdCjfk0kvQlnweVVVEzbHjDivhnWiUAVJF7FboUsGzJZ3
hQx8rQhXlNW2RYI4Hwlx7plqvUu2dXPwDSyZO2FdWmz1I696zxXhDhcrjwwnjlhd
yzTO2MaBc1GKBcO1jQHib79l8fv9Wz2hZ/62VpNERCZ5EBOmLvyuqBwSIkviyhjD
SKgkU17FZiJRk/vooaepnqMbpNBbg6qpie8Q/RFLvndDiPYzdNR/QyhXwVhYkEw6
teho36w0pd2pN+/yUS9XnZBxIGDD0TckL7uvhu5J9YhZ4+x+pRsNBP8Vmm4WV20z
s7fOLbl1FoOhx5aZ/opwwwuicrG5O3Yynj/70LvaPpvPsn+TFFgfmOXt1lIE1Klk
UStEZfm3jPdX9dC0WBXNAUdWWAO8xYDm7Ziw/RDfD9nEZh/mde3Ik36RE2XcoMO1
sihME0e0NzPQ0oVZQClzzb5ccE+7nv8ujKi+AY9JQE7mJlcRMKasmZKuRRsF/yDI
gmLIoApGhQGLkj9Vf4e9+cFjv49ySIqXISk6qGGqiJGJmd55oyiojJ1HvzGfxCi6
KkgjvGCxFD5gYNvBs9/ZjkBQPtRVjT5dorldeS8AXAF2yE+VYD4S4pWY9Z9MGJnt
hOfSO/xC/3w5+JYOJEPj0OS1W13pLUTaBUR5rAriCiPjJD6jtJ3r3WJcyxJ6wzAs
ErAwrjYwdxii8FSG9OD20TSLI4aN4y+V9SyDmD1fed6ThVwO1TMSbQLFinx1MrWh
aep8pSqYGA/9LlCZfJ2Q1IdLgftepqwT5Ev51oRWrfq/ZlYH8EItGwqAI2HGBGKe
25vgyNaXeze/fM0fVmEyWNBp+KkJYlzTtfWOKcq4pRflRbvQkx5mQg2WY9S/F6kn
BekUT0maaKBtscBgJEpe/yXvA0TzJmsgSRBLbeF4nPSZbITfab/FVDrTO2iG65PG
+/NDPQtbBEOOdi61bB/nuZ/fCqh9SLnxgtqdTMtHJSofpdZZ0w67qG7B3SQgQhAR
PT2tde4cHjiuu5a+XRY974gGQzRYUq6gerWzucGGmjV348XILeFfXq9pSE4gLfH3
2DZAFZsNd0mv/hTzGa83ybXEDw7tp5kDt5uZSoK63zwVLTn4Di38d8OfuOd7BDSD
YwnNvobv85JYxAclL7GsOmNgL3Yoqf1Gner8FGmORcVwboO0Sm0rVwg6rvToBwAT
eZEKOC7ruzgMCinGtjva5l3Uy9mt3RUwHvqEjj/xs7AwKGwASSzS0wer6DqnsVAP
m+BFsnONbJEyIjSZTLMMuNepcLY9ojektfRfNCpqjeil4BFaEJm1fjxf00RO3ao4
dqPc5K9hXKhmH5VSViqHHKZPW+74FABAWzTcqa8HNCGSoiI+SGtuSzGeFZFyKUE8
irT+aAy1datacPyi3YYbdWqO4xT7RaV/CF8JXKc8+wsqMzP4HOFz0g/WwmMEF6OQ
5xehy1EcSCCqX7L1S19itRgALsecb2+6zfLYYI7Gbr2RU8adAB70RfEe2dQvqIUU
afgNGpd98+3SXZlOICUdSGM5Pwja6FNxtCLpmF56rL7YQrB00KvLcSfpPoqf8kbo
ENDxILvom691OVhobkGBT86vblqZdtJCohL/ibMK5279ym4vHGHZXnNiON8N8ys7
jTaTztSdAtS2bSdt5awOcaZv41cgx0urzW390dpSRbsBeihV9EzzUI6MQ/mBFK8j
IhQeBjABjUEvG90G4tFMLpy1df+XEA5KE1GKPit2YR3x8t2uQwgqPks8gZN5mTfc
GB2DjMhva5rhccOxDbM6kzQ82awvc75FPddtoXJdFulBveTQ96ZUx+Bdd/NlZMJR
itSEs7trJedKJ6M3Rlv2GT0HXDjtwdYB0RvvFpdzj7UUPSUwiCpx8B10tqfbdhyZ
fsz7SETOkv9InfaEmkpDomzKnvVpC/CKXM4piMOwnCUPdodfVMTH19Z7PMNhKrf1
1jXlQgF7nujQY7pB3BszVHIn4lzlNoT13JlwG59zvn+SatG7hrYq1orjXLaZBQi5
oN0RDN8aSXxu7+smUarFin90fpFdgUqw+VfkKAVeiiVMsX3ylLHW9gDVzUefkG5m
xgz2chSbDblBBp/zSRoGR4C9iea7+goFm6Pj40ibrGXVg1m6OwYZ97iUCDmkKEh1
Eai3AVvqg7o5MDcn08zVLtexpHT0x82if+9GfUmFIsRS0L20zyrh3UXxVJoE+oqD
d2/n750kUlkKWmarRFFv2W98wwX8IQ7srWhtwitYNxWPcINvlp3YWijOkzaQMR36
TnRHQxizx4MNIfzBLkfZnqkqWYxJoyEljnmsPwPlXcx3dEjRTNwx7HIR/wpS/zgP
9fPsGSR1QJ7cst5HlBIJgFGdDfvk3/NEf11Z5mTj8FH6buE6amSiZth+rb4lEpbR
qe+0eYBeBxUnO6h3CqCBSL2GcqVgJ2H3iOSWzxKSB4DnTdJALMh2x5Wu5VvWGWy1
w6vj5h6DmeiGN4JXXENhwKRHaEqwV0tQIUjzWtN9F+MklFk/tSaka5DpNhF16UJL
A4bl8hbS2DSiRXzBihvghJJlE1Bh4RwwsJ2H5E+FAaOHe8+JCNl4+7MfKfMqqFah
OJHhzL/trNwgf1tUpB3+wZ8VHauoXRa5lULZT4Ze++jhnidy38QXD1huBAlCU6GF
iGKuholdf8VEZu5s+aNYrjlFqoRG0PUqLvbZiMYuuQy8FBzlBlMkqx5aPc8Y62QT
NHuztPqhX2kv+/IEy3fXMBfiNopBdWbHDsIVNStlj2tGj+SGATmT3OTC1xxcroK3
bVxxdJ+BxrJ57AaF38vSo2aXcmyGCvtBQX3ur5E2NXoLew21eFtZXMiyrTk4ZVE5
J0Mlnpvs1ZQk85N/FtjPFUC66cXTTUKceC5jhVYAyujEkRszj3aEPGbAjnEh+5lN
kIt/G/AAskn8FE9g35Bk8BcgT6XcILBLUiErkx5vlUYunHJF3bVsuW34REEIIVM9
XAYaVZVPhFDI1kkbpr67gBwbfxWs3/HyD/jB+8M6K7s4SREr0Np3ebM9BejSFbqn
vMa67TtrzPo7UY9LEILWucuxclpHBZrSFNhaul7sEW8GUt5hdm75VPyQax0y7wbE
oDl0h82ewbMnv7TGvdErGiZZ/Rh0xeSKbkqOheBDhdch0Gs3nQy8kcgJunooLNji
iLw7P22TOUp2WjU13fZuEeCE9HzfMczy8UdtHl8dkKLrrJZerv4k/yEODxjSqOxr
PX5DeF8s7eqUFoMmQHY90ijJtVuuiFAvvpW/5qz0ImY9BfcV9pj8EZyfbuz1u/gL
sUBaopB3/9p7AH/sjpHIT4NTUNRPV1/EvuIu6r/UrPVVpDCKOdbbfr/KhXTkNWqz
6YYrkeu6jdUndalpK5Boxjo7zJfYZmjrUV+p4aKuF9j7Gas7aDaYwJlhXQOGMxsX
d3Fu9ProuFUUGUxophzXM7+nxo/20ArYUgaim09vGmDrBM1gdq6fa3RBhSimXXDk
0Se5RTpOHVbG9X73mIal/8UxllYHOdZIW7lQLQQngtl3uttbIZHJff07ZC9tRkBV
LVxTiexhVIPayxCL2Tvppb5Sgl64gafTeCPmCSUylUqGtP76yrspJYJj3tOWSTwE
djmjpb3UbWXg74A0d4bUZqXccmLYBnM2NIX5UEUvn0gKN3jPuWjFW3RzXkmzsHUb
VOiH/didcIsLRMuJuBA+RSHIUQwT3tSatr7k/vRi/FUXnDXOT5pQhuteqkmZKcKp
bYtdoM7SYZcw48SJh1R7rbjmsMXDJFqOgck8xKsKvMm/STjJ/Rskbcp3KMWbqzzH
IYtmhkizhz8MwO8PvcAWZ8VGF4AJYYBXIlsZOS8XS8h4zfyUqOkwaPjugHB3VnBm
E5+xWmXm6tHv4jN8Umwyz/JKqcuAigpTFcVTZQZ94oIwAJoHoNLZdte1rTsfg1pm
ClYrtz/2Uo8ZyDq8Y0BpXqRJ4ntq5IDzvaT2iDlJWBJAHycToCA8y/Lv7oHiiLvW
9U2tbp7pCIu13rJM/sxN8wt6YhJa4+7g9vNytzhwnTwcVt9GtTr9yOTcA73AYI/S
OScEblQ6T/cryFw0Xc/Yxie/mywdermsFJVXotnTbfv8zPg8qmNjdUHxcedlYovm
dpZo7cfhomvzFGBG5vLgRsYozZr0vORMocVy/x9YbriDFPeBl6bvWurHajeny8nd
1nD3Ygh5X2nBadtsH821m+tc/6PSAURPCFW8zxnnsTWZPkZ9KXwtGbL7LugpASdu
blcGIrFB43L2cic9Tq7/u3AKYqUmMoRvIWG+K8kiIxXqIj38AeJncuoQijSP6ER/
gpAxQf/5TRyHQtJWg6r17NMyCfPbQvIpBDcog4QXM81kvhmbGRmcEsIgGB9V846u
Ex3ZdSWb8EIj+bKFEfgEdUEoS38H/j8ZMG6z8EN1A6IxbBm6VASiespFr1vdPhj+
N9gpnW18H+/KXMN47ZBf8OWlN6vuAq7a2DQrqI+pMOiatOcKIDcrkIyu26Hneh4y
a4DqIbbyl9YCI9vPRayG8HaHg0NyN2ye2rA9m8AI+TKsQ06U8LKebEdi32XbZqf4
bvIIwPNDrK6V3njxsBwkTks3JPjehch2gy8chza99IPd0o4ioOz8NNcoMbnqoxwK
y8+DCjbn5HDNObfNUnvC0gWjgIMJLq/faUJQxXzH26SymvJxhSFEP7nuiMzBwvww
P2LAZbhpOHswI8JW+HzZLcqKsTpEb6P2OMpCQZWYjlLOR67imuq0j2hWa5vojY3D
1EFuKdz3x2nRskKcGY39k9RJXDHSokGT/W9CZF55lYCtEs5sQwEjY/qHjXYmuwqy
MYkhUyxG9ewr5Mac76MmynXsJohnZ+xJaRQ9RLG3QRzHulReQVe6aM5VzeOr9Jmq
4o3wK+J77yALxukKQeyIxAtCJvpOh5sYxERHD8p64pad5K0H8KgUUWt1cMfuHqjP
eYPoF0A4esBe8l7JQSjzB4qYi4R7+4r25TZoqyDn0yVaINe3TMJPphr8j0QGwbV4
p9eOrg+C8miJfK3BMziMRw==
`protect END_PROTECTED
