`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4wve6Woa+BmWVse6l7qnxxgq+ZKxFFjVUxgrXhIzqhSH3X+5W0vtMMIekVeSeBzH
NnntZHOV6zWOGy0xbw2IsX+6MRxBFH4QE8o6ikQWK4xp5p14J9rX9/vG7N8TefQS
MgZN/obOQCxIumSQEnpD4AotJcnrIYod9hGoHzg4T2p//VrwDQC6XIqXjQAXhlRW
kxuriKKqAB5nbKZkiao6Yzs9NItDfgmVqJTq27fipnfJTrp/pp3OpEuzDcwRqVID
aGjl9D9ZNgshhlo5HRTBuQ==
`protect END_PROTECTED
