`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
chG1reiW8S6/5ZCJ5O17uYpNNo7/KGMiJSh32B81CHevj4mio9cvSfFQ6cVGA/Ut
DaFzLsdxgqUpy5ssVUjQQvh7sz13Je81jLoDi9PDvbjhq83waDhLlyRO7Md7OKF3
ZNpLR/NDhLtkQFNmYmo1X3G8Cr/EGpQMIqMvjRE42FLLu7B+ahdmOLuAUIklzYem
ZNFxzD/scPHs+VFI3HH51yTxKQyxEqjUlHqSZsj48Uo1w0KRM/5qOV7XoPxgeS6I
a6Ovje9pBRc+/YeCF67dKDXH1Y4EGK+Mt3Q+hAFDMMAe75SAMZgEMDRojcTJhO0W
`protect END_PROTECTED
