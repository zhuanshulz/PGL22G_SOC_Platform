`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8cOeTonBa3jqLDi4OQR/rCztqfl0xcPNEGz47V7Js8/jpXQ+dYDwHr6rupAB6sQK
3mNXEY/Q5X6VKrUafZepRRslRXTNhN0GN4D2SJAevHIkAqr1D7QlSkGCvbMQ91ol
KKhwZjM2yj9frlcWdlIXv+ZNsJwXINBV6vpu4pTxu0gAvmaZXWWywCiXUGULW0k0
bVCTcugYPfz7umFhdo9gfy1pqbtHYq+x8HbLxQToxAS1njVqIZjUqiJWvoQ1NS/W
AZPGPmEDYGccCz8V7UmprZZ1ng7b3GGtFrkyyxNdlmd+004Kh2VPJeePB5F90Uih
Lsp/mjW6h8T5uhNajakGaw==
`protect END_PROTECTED
