`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AKizdK+wNqaT85Lh5p2VQt9OReYIN3PK5HsEcrA2UgE/qn0W2RDJdwre2tcHQP6X
h1FWTYPi+C8haXKgy9gYPHDib66ihzXjMjzhKUyFxmcrqwgsUFKauz62uSGj3i+9
GMKoS8KgidEKMHqq5r0oVkTGNGveyPM0JCnIwPfgrxrE+uc783VD2usrnJUtqHYu
FIcz+V2ZCvXsJzDuOep0j4aZx0Z32SoY0XOR2hsjhi71L2GJZXZBsiLWKLQ+bvsr
lBJaXXIuWLe/evgUlG5x67aGZAMBdjYHoqLnI3Ef8lDBlp9FSk8lSy1e6ahYmupn
pNUhfxL9RP2NSrPf1vyY75w+yliKjjhrUMqsZJ4xyQoljC+jQqTgJ1SvdIWUXQx1
RU76j4aYynATYV10RZ2IP7LxdiOx0oqoNuFm/xB8CBIA8jNy9biDdt9FEXUM9XBj
99syJ5ccrNmGH/eMofYfyx3HzWEL86OTKLNCPiE64CM4YroYEdEi/kUKwwr1+gr2
NDLu/NseJKyB7gp4bv6pfm+SRlcYNeiHwRvK+ThJuIqGhPd9K+rKrO886JOk12Mh
RJN+8BF7+54XlS5axp8XOMMYtls8va/t2o9PActV2ygjXMPVgBe4Xf2Fb0edhhGe
+CS/oN4wqVWKkvU6+509bN5rusTzsONEO7GyI+9NZyyl1HExfWrQJtrdU5u+OgCM
SqsXaCLMXjl8ogYtsgG1m7ze7nqwsD67rKqqmOk/SrsapAXxuAHWrfvKpc0hxnLC
DLrwUr3e4uiHn6WpVNbvZ1VMqtxdeIxwaonAzJVhVi0hx6rL7Y7lD+KG749SMu6Q
Pzyck+aOfD3/xLlD/u8PqrGl4a/qUnKjvL7mmED0pNuYp56OD3tiuwzVxgn2tnb1
T30Z+FgV9NbDfg92lXVCswCgcGeA2r+fKLTM//1djFqRzcjCjIeoeLUvI879jXxO
NChNvUZzvzhAcwVywSGkmc47Z/IVAcLE0kqHntgPcBGhHEy9TBIuGtJ9DTmw67Jb
lgihmHwq1TBSNlLYe6P9MsXzunyOlxKXOHRVQ9Qi7Cztq9F/+MLz82MOtO98DNIH
HGfsuomb6Ield7QgRZRMEiFIbA6t2Tp7eoHvHIRe0JC3tCTz3uTpLwfaosgYFkqp
sctOWVG8UlGmleg5pmTz+7vFtPNomk/hMwCAV+5bJEv6li90rR50zaa2PKcXcQ2I
3ge0k0KM3XEFAa8CmfSnoplatMwYN9hrG8n+UE5RPQX0ddUEPBKNmO1AR5i2vfFr
UAHDBsHEkGdODXjjDeaH0Bbci/M37xHJ26ssHr4WEZju+p+5bGQMoRvhkG6gjAn4
R6lonQatXoBnQSV45/1gqUIEZsI0KQ7ycCuMqqFHV4IqzCd+dAmpplpwH1LdXRYC
bL5f9kMevVNkAYMQmb8St0AUq3zi1aqlFjAdzRW0URle7BaBEu/HLnGi9vdB4ejL
3Ca9dKfaaxUEUouxKVRCQzcABR/yYS65c9tX3BliA4mtkagzTkZzs4ovAO7nNkCe
dHAO4+UbTZJAlR+8GpZ/Z25hggA4g/GJm9jZyo/f2M/ppUqGGxOCHAK4CPIojBFl
FINDqEj4caR5CtU+EKhSRYGK5R2jrqE+JnsfIAPZD/zLDcZGj91wmhDR2o2veMxm
Xt7ckDXXnUUStZQEpBX5bV3U73h0wyrVx5bTPXS6L8RJ2LAr5Rk28Jd/xuz0N/l3
0WyD1IxBt7BP+gdWCFOuiwg1GSA+xloGOoyNVEN05F54edKijoPOkwewJlnun3Kk
zWKCxc4T65gxDeRwxymAC1OluQsTkZXrYveXj1olodFisffsF3fUpUP8pGlFmGLo
lJ21yjK/LwHZpc+XppqRC1AzaCRm9Q+VUr8F46mNOJNtkjnjna9tw9OWCE9+nfbf
ZbPcr+ARAcyspZM7AVHIR1JOoIm/aRDg46Z0T7Nar/TM+WpyecQYyWBC4zWrokJ5
BVs1yINKVAUV3HG++B39ydkXVY0QG5MLRG/9KGZkekWST2l9OU85T2LFnOAONlia
z6WTpRW2PCGfLBACshUtKzkx26scuXwN7+JKL+mfU9seA/UDxrnYzC1znkQTS/n4
qCOulX3mJP5pzj56QTRhslHisHhi9eAdqjHq5Zs69xkWIbD9/unDsQngCnxVhpg6
4+p096ZDlvYbD/2tLk2ANvQZ0qCmyep8WOleKT1fcR/AM8RShRJuKfnlkYdtiO+Y
sInXuzTr5IoVAAAVk8C1dH7zNIFr7UUw0ZCl6oqrfIqMG1XZl3rDPQY7oPF7aXEn
xM6p2nfE9R/NV+k/xsDx5Rn/TjTEkKXAYjiRRUbHecCG2wg0GylvhRIyMeGrqGQq
937yfDgh2Glw67u8XgzNXLTXOQwE0jGWSKBTomjLabLQfeiecyf77X9nbOwGp2qw
h5nwPQpgu4wmVKRwsi+IFsW2Stnx8hM8OFyynva8RyRQZ0j+U2J+zLkii/t4x6xT
xtwigbQ/kmZ7JnK69v8z6okszCApOY5EfU4i/4aGkVUgfd5LFzBP3KCu6yiFN/+E
rRjdRcAe5H0AeY6wuNpzopMMDFdq0ZkqQ6VDLz9BNQ4biUh/AruVyIoYyb8D6eI4
JRxBFrBAGopLnD+KZNM/JFRk471zMKGZGc03U9/zlxYMEAPaFm7Y4sfBDf0qCu9B
G8NyDRI3DQd9YVuwOfFYNwlYURa9QAoI36j6W+NaqFMDakyBLE0s/nWQlRUwtI7v
Y0qm8OAs2QLoslvhYW4vLCzP9MMZVA5FiAXaUmVJCdIsZUpYGE36k2lhkEtt57JL
Pqaye+9q9czrbvu8hMpoJqoD8moG4cosTNgzEnPodvBgmuMYETTd4BwTB3h+RBIP
jtLuxBtPvZyP0zWugiBBemWX1JWT9U+mTAgCVodGpKT2sl7jzsKnbE9PZawfkbSy
2CXrdzUq/gJoei/040EFrFEqmhU7AAImtA03dzoa14U1KR1UQ02Ioyrz9SiT2ZgC
RVn/WIr6leGvCayQtLvHQ7Qi9Mj/+A9nRHyxZnRWEnmgwD8uYopRVceReHHI9MGw
6xYYti3nxWjOtEaofMXCGK3EUfBL7nuIrun1gln943+owFCmvm+NNgPlTDrBK2df
O924wdJ4Xb1ZLjDWqs/89MFybCO0lVIs4Kb5as7Cx9rOlQrr+1MXBn7G63mDq2oQ
7iFeIhVpB+qXIfwNQx4eDktxCeXfBZXUK1DXbanf2khAwZy5tT7JY1VXHwJ/kJVr
BuuUCbHiWXMYLsfIAPJOPoc1+exA9foIUl5eHM6BlRGtbDkMv71QsfBEyFyHfXPt
Uv9ykb3gNt02v9j8KUKDH996c7u63Os3rn2SlvoCdgaoWtSGYzLhRSKhz+cbHlWC
qXPyc1Jf7iO46wbFjjZqi3gV4IpWE1PFmhWqlb/LfLOnyvM8nOpef1zFYcEGYv1k
2ybLIptmwjhsqreJwFstdVpKDNFVGUx5O9VMEEgti14vvSvskVhWlf3IdJbAV2lH
jRcLrwh1czBRKcSMH0UCYDjpPTym8cMRCS3flD46bWy53ovulpkO3JcsY1Tja+v6
OviX1rhaBTSyFR5Zp4091XV03kPOEO32kehyI6krikZSCnHWZSO2AP9wD0opmE2S
0zqRtO78ZtMzL6qvCPJp1fbBzXIAAHQpaQqLUT8ZQJKkmcg66CtEZOwcqYbE7JPr
3Du9JdfD8X0KbZYR6bi7MEEPgeJrW1NZzIoWriZ4JbB+ALCtVNGaPirIHIIqg5Cb
p6aDsvV1Ysm6hybEDehpNE4KVjjyenC0XnT31dDTAjW5yDI96j+utkXW6oe8hR6I
pobnex6NigDgW4A19Hh4L8bd1cNRJs7+wdaVJIkDGB25DtiGIoi5+CVDb2hQ71HZ
PStZ7B5kr4vqUh2eQlMUxrZhajbnNv4T+yxdNo2EKNjlp98QYytsU6cyWUlp7iTV
Dc8CAh5qVuG7FV1mhN7owdyO/tJRJuoJG85TGyFk4R6lcjCx7Ee48M6uEw9nnBU5
X0EGpkRqKWa2jaaSQX36nfLBnWwOMJlhoJqT5suT1iGKnDNHyUSrOOT3IY18r1jB
CLpNYxmt8zLG8vj5XrT9ZOVXaAsO0yCLsyRbeebecDnSBicHvnbFTjS02wh7ZDZ0
CFJzLuT8fBbdpQB60M4DgtuGHSlQluxrI/E/NA/KztCyV3ZBHnv8MzPHOwEK5x5c
CVGMdDK7T/jeRmGhkzq19rpLOv83ZCHILsEi2U64xEtjzF2R+dMyraw+fzHqsWOi
RXMreHgTXRmRaq0n9QPmtfoRKlNIcUtuzYObyH553WkiEi0t/VEBdqPW6D+nvwEA
+a5h6VhqGb6kQs8aoZNB576kM4odpMPY1xaWAtL3X/rj0B/eMsQnI5j1ql3ANxh4
dp+7ifaVR/s0VQy9xoXntqAwcT7N+7OhCabyR72nWwYDgRE+mvsBLz0hDW2yVcPZ
UChc0YA0bV/5MQ75Dbuc/Mw9X1sz6teuOOk35k1SMn5vLQF9GgZm/FjW/N0aDDVp
NfULzRsitfF0iRQRfoSWa0GvOZwxRO45Qi29gnlDoDcGH86XBqY2N5gpeU59egCv
UsDw643nUXdBWQeniVAksLhMgH6jUDnkrPNwIOFFvvO+8MRuoxr5Don5XoVTZ887
vWuwFofRek9WMEiQtUVdikRJiKU6HgW5mzqyYFwWZVJXZkFY02mfCT9O8KHLDW0+
zufwqjRTLof3J7Kw0sQ18a/LZn6S+3WY+HLuBXF4JaTiK8sdTp6Y86tlBIBjmy1R
AONg+2Ta32Emeyg0rFzxds77Q0fSO7DWoBDjgj48vuLCDjhg8Yok9Qs1//cj2B3S
eeNfpEFe1KkIab0uPhMX5rROC8gdIsXpfBRUYrBod0ZjC0+jzo3Lft3nZLCnR1sR
4XROav3QDt1Tc7YY40CsjGqpsgwFEvPPvnAdfvgW10FDo0rat42Wlgm4LZ71cbVo
Cy2Xw0cUikzqo/0zcuOQ0jp7NjcDW7Q+NQjiKumafkHozQ3BpSLV8cPA0siK7sqD
JW2KyW+9VJDg59/pu9Q8qYWhE68libNawEAOSirXWAG9lrzeWrBtzQuM1YzGXX9E
sjnxSx18GMt7RVTuaozuxZcot6QwKcRuUi2Tw6UlmCPdG2OgraG70i4d9Zqd0Rgo
8CFEhAm0kvg8CNJmTkBFbk83dwI2h4POIBd0/OulvtrR6kFHq290GnLE9rZMKXwX
mjhczStYi+9CQgQS8We5u6hFMLh4a0QWlO8hWXjlKUNL6k7OdUs0kbQlf7U2wDmp
J/jeXsC1pl+M91gSMb2Qo2CM6QPwNDIlS/bSHrgkW+UiPyhiLLTbi/1Vr8lxLTzl
puMLc1AhLhpf5fMG7BMmE0/51J2hq0kZ29EhQDx8zB5nBTKE4j7hfyQAP5tKyLHv
8JenR+enQRVBmLvZPXRGjhARNsd3oOSC+dVowvRQg227/Q79pjkIjRUo++c6qCP9
OBhOzw0ONOOZJWcB5+xGYLQpw5lKug5OlnmRZxeOicT4K+NsGL7EEaZFgmDmSK7U
28F+6B5iKpOELmL4C/Py4frwX1DKlvdgWBkTQaNvtVwaJEwMdWKA/64dYUzIKGIe
48NMa7ke9EymoMQhIqLI2Zev2UVJChiR0XvbnJlKiD1T2SNM31rRwvos390JeUUR
u2VqLxQOPZ4O8I4W19gpUvv6E1HfILTmS6EC29o1MM3BoUSBYOwNxGB8+sjp3xiX
EZcLFCHLyOZd3V+/45MYlWnz8/jRWTUWyVIn0dTmu/K5fgpA57RJRWWHfV0b+q6e
gZf1KJKQQ4H1z+aGusdhqj0YDcFqNbVIvux+gSJqO0TDqfxPdDNkZksJdxboBjWH
MRCc+8iPSZVrt5CxeTl/mLOkQbUpfIyEnPOB0ZWcoOS7rq0Ub4ThANvaSF85MScD
J4GHSovTMfyF0673dCN3y545KGd411oThGk1Ex5TRJ2I9aWeqnsAFXxnuebleLoJ
5ltCLQzvDzelFPFGHZpjanl4Yp2kAbjWf5iauF9nxQzOf2l8GtdXxfgFNjpRQvvf
qDqH/ZqucYdkx8H+o32K/ScZ8PMmU7D8UtHvworrjpx1ZiNhSaLbknrXdpYHI8yn
P6ZvGc9vCSRwDtwmQhgRv7sSup1C3LoB/mBu6z2mf2+ichBeiHYDQQuuNkm4q/It
kNW8vhytAWx23rPIg2l71yfCQZnx8nmCA0IposfZzC94QjljKWrL8OfcpDWYHpbW
6vG71ceoV8mCQoxhEymOcddsgCW6bi4AYTjVxseDYf/zyMQYwoHMYDRSkZRktOZg
r3BqHT/SwDEkV0VxXcUUCR4/1lvD42dP7zVuy04Z/blEQ7gCP6SykGQ50GW6u4yh
Tc3vDx20uKT+sngiuKOWbwktrKJry2XTQ6/08iuXO729mlAmo9YYdNQpHa+PRb//
55Ah0H02eraKTNWXTPyMZsm+pyAitpiArMMFbttfHPVZfagTmYTdAqtx3cRx3ThP
/n7EM5WA619ONFs6kKwXRbKDxdfeX7Jixr6Z3blajtEOGNCv9TaulcREKMs1s5lX
OmpHbPL3Y970m6v3lIFSm0ijPsygmnTxH9vtle3Lmzh/QdRP1uuE/EZ1bOXja2fe
wh0Cf2KtTXaPnLnc2PxbbmgyIq1SuDCgve9SKGY9GZELXN6AmJGKq1864iJcpPHr
88b/AztqJbXAssPIOaG8AyaquVjMz13yPzMSsEQoan+UuqMmC77ISqmgDrIfBIkM
6+mPyGx0wP4LjuXKGJS4O7m4EwHiUgFTFdaWsnfo8/Ypvbm690nm/d2Xsj/p1anu
zWNfCFm3uqPW/476/uiAeuh6ZZnmdeoaRnjztR0/qUINEbjKzVCHa/CpqW3w8tKg
V0kQPnllWgEGP4oME2A7nJn2CzPBwYu+fctCxqRpCbCDAfXtDeZm1hDvWSwjKaGo
SRtaBqZRUMUFAc+bfdFHescr3V4v9G36hWDI3X2cvH+IJtISiRptbXOCgWnoR1MO
WTcPkpcH1qAYNq8Oktx7t9ttArcP+UAFCQNeB9uPGJluYm4a4VfCyBsticA5LB2v
0NrdnFAPa74ah4sTe889JFPbBx0PhEgJ+bQTuOQu/xrsCrhNm1YUTOkrcGBluSwD
GdDKziR9vG2SxjYFB2uu8ULzkAwIbPXyfm+e+IoDuxI=
`protect END_PROTECTED
