`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YAMYYvI5w2JBb2zIOhQKjrNYLPkHsr4kYupaWS4KHZ7Iyc/gIJbi4oG0uLTWVouO
8x1G9/zn+T5Y8h5xXyP7ICzuTjiL6ecf7uNcda6j8X0P7ry4S9Gv5UnCYjxdemJM
8yIZlK3kDNO6yP7L7jEC9qiY7IaGtmWMrVDH9GMDBLKvrv0aFlny5TtiB8hwe7+m
Xg42aUqjGRAtL9k8+Wva3NLWAQygJojRN9D+sv89yEvSU3C59xb27S7z3wdrg24/
kyxQrrwws7ukcXQGURpTR5ID02yOoGUuhc8KM3tl/zF8YddUIrEJtOmXiNO+yYUp
lXX19Dro+0CSstNV3KZkkxmnPu+HTZCcn0paMH+48rJUT6H07LNXG92Na3YwZiJc
7EgkI5uusl5hQERjje1D1BNVWLvokunZZKatyKGMe5tqRSGuC8RNrMGETACXef3s
Za017G8lwK8fe+4svIkFx+aHC7gfpOdzQ2hbTUzDSwJ6bOhmCHZC8KkoHc2ujPk3
+cEN/Ezp+M2T19OFoNLoS/T9s8QwOjJylCaaNU0fevlRRUY9fO4hoYYJ82npcqIJ
6oyiIZKV5+kE1RAI8Q7uIxMZ/FygNPlsGDvZOffN3ofbdDjjTFBA5FMn3sQ/Vxie
RvHyKVg40pd7XSbCn8XPfZvLEMjOl3gOHUHYGZtEpUj4JIxPsIoEF4x0JnHfq8+a
c5pLvTFnNbKvKR9H0Hlj/hhFbnZZbKpPkQii+pSmJMaSFw4yRTwQVeevkKxqo3jb
yzoQNKqPOWPdkoiPCoxYKaDprUP7ZbRE8rTXRfZLLvH/Alhfk8Mzo3EWkjQMwn56
iXwclnoWWyUPSHPoiZjE3GZNnM6hVKbRAFNVlohp7co9m+hqWwJv+B9mlm3HWz9s
d2jUMbT+3e9sj/dFmISwn+R9WAa67NXsYn+0C4GdQih4TVnX9CRW1bo8LcYXSdlf
eODi1edeDgSiQLwOEBTb22Jisj6JuwQptRmiDnp53IVEI0lwe0Z1qFmZX5ydzy8K
YbkzFpdW+s4Y+pnbA4akRmFPoDmUDD4puPJyp0fuYdG4m/yfYQTjGtliBit+O7lc
7Ro02WA2RQWgy+U4lcnk8DefcuihH6uxcUSiJXE1KJFypL64KzbSITPdaoZoNYN2
RdhfKNy5+uHE5txuyW7MSdo6kn/7+bo3IgM9bkzglv38ebVnr5WzopAqI3+kL+Rm
h9f2Fz7y5xXFehRgUN/kNFZFQ9/SIJ2PNEGEVnMPqcvZZIfY1rmlkur0KvKSS6x2
3ULN26PFQNga5i1sVIqeiEnzUjyaSM0WSl5QAjQUK9LT699uXwWebo12KGGNa4sW
UbJMsso7FwyxK8O2gj9Zfm6DpIKQbBfigbmwgxqpI8MwRMlld4G+ScaNr8G0G1rb
HCd0P82xXSlFMNhW/etL6utyr+lev/J8KaApydkxL9sALeOiQYuEZJka4J7bvcze
vNot5fP63IWXxw6WN2zfyBXfnsXfLbCKJyKrtcYqQxXR+XdOm2aFsq6fHVKg6Xr5
mq//3uU3wLiahH0iIGfo7vTCKXQfb3ZnVLA1vlBLwZ3gs1DD7UO+Zvn6U+Nem4F4
/0+JUBA1xWlMcLNBGAYSauXuCOKU7SW0+24+iLuAuOaTDjJMwox65bGsWbg1ISXj
7X4VG3QAkuP/6nSr3qOgJSTmc8unMh9dmWChwDLm7x56U5xrOsvTfhMq2ji5zFpd
ek8dAd7TVqX9GUxWe/QOqBQ8rlqHwUCj31TzMuBh6XM0F/K0V/dL6LjblYfvFaj+
A0vMpVAqHFKStaqAtYrPES/cCztvgdXckGjx8sZY3rpwDBJt+zeJ3HVob70Li7CM
YNYd91b4TvUgUD1DlLIk5WP54djdsNB+LC3qkpCKotizw56Bo5LaNHCtO6wXwXkz
sqh07IJ1a1XVqOK7en4DkiRkoyo6yltt+ZdCcc8oLdB9A2emkQ65VUwqPPVPq5nH
VZZT8nLTmx6hCTAOiLbInwRECIIoGrtsUMKdUArzL3amUSl8ek+xokqK+EAYEu84
tyuD3AGnpM3/nRvdyrqGsfqUaL+qVpiBqWGqvxvYIrhhguJyKFBkHbPqCdOF3w+Y
mhVXyfSW+kmJ31I6tKQqinsKxspksFxuBYn2PW9v5UY5RVUkbLOVg1FccqCTEPmt
3Pz9DVcsGL8IDgreuTU3UK8SBMsebhiCyMdZV5NSu6snvmtwqh3notZFlBcVYk/O
KI2zpFBoUY+xOqvi64D/LhXSZFBJ8u8OS57uosyphCRiMeuDg7mZ7Z3glDdKQ7hY
pQxpXdoJdr58ISYFjYmT3diKDtTb8wDfus6Vo9i+FtLxR362c+JD+y2Xmg9toeKI
Ux90LZNasmDqOnqytEnZm5XvUgMChCOHOzMbV3/kbKCF6fjj1qLK/Mu3hj7h8lX3
ax835o4kQbB8r8z9+LHym+DAcCo37QDJhRm2Ob+xF9HR6UndMCBbIBH8M+6flYoG
fnNFtw/dTPSBJp8gF4d1snQl44NRgOZS32PLQdal3j+x4K+1lKriVuMm8rdUNNtR
YtfTHqFl0ne6IXKO+C3Vup6A1uh0p1hdwve+mZNbhG7ok4elvuAXnsOgjx+cFYyZ
jozZpmg78j0t+EF30Tued/1/C8J4gRiCNKDWU81pyjCsrTOTIPg+6Ftr33CKYNnW
4H3a6Srujm/EoxziH/jFDsSvfDoiCAjcCx87WDeRGusqRcvUCbaXGMGA/GCuyfgA
+Ujg+Rfqb1aHY1TkF3nyB3Gb4q0rmk6d/jtbg5hRjtRXeylWMiOPQ9t1sN5a1Itf
fuHryJmhIbrDKXqO0Ujlm+TONtC3R/YeK1S1It7RF06wGxI9HwGDWI7Wh/n/fRbi
JChc+7dQs943H7Tgry+hJDVRZR/Tl8AkTrtDUtDAUsxdIBGniJhpfrKgQxo+aDlc
sVMdC+5ZY7LdGcVPTFmYEtGR+FjedvTXwmn1+sBB2FoZlly8+/4VOWmfCKGN9vNL
hlLMM5lpFsKosKHs7ivywY6BkBEm3lDI+3VxGnmzv/4NcNvggifP810zD0r0wjxx
GFV+0AhrcoWQvU3D/gw77gm9WdKV9q8tJJC0gxEOe9dx7wrbBvtiTSNN0GewJ7pz
exVtEyy5muYLjPoscH5kIi2TX5EhLQIHWc/AS1Fmc/L3t5o8ymUGOD177omHdhlm
P1+xi1MlVhrtXiZfisfw8N1z5KmBFbB8Z6XhCoukvSptR4RPzwFjXim5XsoLprHy
b9D3gZH3Tc2/OlICfls6RttkH7IWuNrkGdwfIkfNw8CA0nkqj/qm9X3lXqoOimg7
fuVh/g70c2qL5ngNzlyyyzoL/vivrTCAYd9M6M/cBLl7ZOVwsWfIUGe33bbZQbSV
Zi/p2wiEWYzs9PmYSfeAkUEW/cpkM2j+Pq33dKETPRHOOM3d1kylvnUnZ4BS8Fss
3+Mq1tfhDAfoac/cYKecf/YIbKleymEx9Ut2CaWk8zxVsMHrN7n7QkysE83Uov+C
hy6B5Dfsu0EwRTK5RKbrq/hK10sqtSCryoHv4o7fOXYQuJO/GhB5kgQ90/GQQQSN
HSTW9qofT2+KpyW6VrD9rQLUl/77K5OWlIYwnEUDVj6mgZea2XZm/lvix8jAlEoX
rDsgGDddHxHAtg2JxCQzIJS8e/ZnIFlqcZ6u7yVnDJxhF8Eiscc/H01nJxJsw+N3
xMRtiqZbN63pAwFcedye+eDA2soACxxyDVcgObOsj7uOvCsN+1QXrUapi9pn0zKH
wOiApV3KY7Hi/j8b8/rPfbUQnwSjb+siCKih+lfMH+71PfyfkbTS963w4WQ6hBlr
DIIq5zT5V4Q+MuowQzTC65A4UMJp3W8T3WXMEhQ7raXUdNuh9GpQKQjly+AxhYMW
gzxLrkFPCKH9MPF4Zfe+NbGYosKRL0Ji8QG0Jn0KYxFV7Z3Fu5mEyo8DPH2Ntjib
YJaSawyPe1A7FBxYIucgk45sl7vS6YvvsmJ0oyjIBNjXIqCbIn5O2Q26RVlxN7sQ
e0Tn46nH8FblGeWXhwq/FE9awYx2rmSFQkuTLgjmpfG+8403te2lGmwEjU1G1NHa
CvsNwfejM6wMR9ZNBIRqn0NbLrbNRXhwQVdWnp5Ncxfy9O3Sh5DquJ6O8/2V5tWh
aaMrEocaiTJNXPMr6nlL2QJcRN1INRSUUGLFzf2uumuBPYJ10924dSQcrBad12Nc
IsGAWiAXbQmNW8z2M5gNLedrGDET++q2oKl+CjDhaALbc+viOqGlrE3/LTiqQRfk
gJXVYqLSESzjHIVVesq2kgSwY8ngo+7syIjlti39Quh/hiehmaogHX/+b/iFaeDo
OqxLfn7gBaJD8bFojiIuXoDWxE5gvXUT3WA+anS3HBQuxpnI+XyItgKhttpBebqO
KJq2GwQjn8KqqWD4Idbl6AK277dmv8J9H2iEZU4bV4GAVi3IRgvnY+4LVkID1TLt
bibrJ3iFieiQRDf1qgda0Sj7hFkXL9LDo5pC60p37OoBH2jeT2e5idnyXOLp3maV
ZJjQ2hTLg4I4308d+VGUWdNw6P3xe0g+deRVGR3bm4d8zLew464BbUa0ndSCyp5c
tcs+cdOPFtfjdJb49H3w5fanAEcbwRtFhg1CBlETZtY=
`protect END_PROTECTED
