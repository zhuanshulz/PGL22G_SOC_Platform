`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uU9ih6n3pDTVwuih7vYv9jcKvSTJk8sj7IYzqkazbiD0glA7ZaHgw/eh2pYAlHab
xFrRvX6EHHCluQtZYcc0S4277ymtXsh1ZekgauFf48gf6FL5n2QUcB5C4HgQT3x1
ZcxXRY9tAp/JaQygap04e/+6iA7A6w5wwuZHiKYzpXarHLJHSxv5iIXhljKxKb3a
XYSkBRHRx3R8VeheRrAY1xUcGh1B3Zza3GuR9yce/AiYIJqZ0vut01oT0SPGl1Jl
jqHX+t/AZSaJN9CX7EduRnIpd4lc3pHQVngkxWEmmK1gogeUgf9zZ/N8McOsulFA
BuhTNONWeu4674i/af7tPKOQKSpZSYP/45rAgcETYkI9HjXUQSjj6x/YYqLW7jnp
/eT2QaSLnbxOCnJHJ6BjpVTpJXWWfSd+yVaGO+dmUTvXgfEKMVCLfdcNOVMfatJM
7AtwDsSa/wDOE0Qc/P95Qm960g2EZNl15LN9MfkhadoST1SviaRhrpBaSYTaua8f
Eb541jxmsA4Z2xfjWBml1bv9nRwTNEnHMThB6o2C6qVD8AMHD0g/CjgfeKpSLDcH
ZPjy+D59R3+kEqUXhv7vzMxEk3jGjBtg9q7xGpk7Ydh8otyi2MiFbill1JYKtLvR
hWnddUFJ5kVncUuSwMzoGoroOjMpTDlnNZuyNbr5n+dvOcr5ov89sWXG6cmJg+z0
TV6M/alp+w9fIwOjejB1aTdOFjt/Vw6Y1VaYg/Y5duQNfuaVLmcN87wWe5/XuSbF
5HJKx4WP6t3Jt7ZRop7bx9t+j2/+6nJKjgUO9G7mynYdNQogDFSdfgzuPXN9mQog
vGP7j4GzP0n1SC0uqMqs1IkJWT0MYaVFecAYteYxYEYYq8ERm5GRD8E2Ujec34/V
1nEiMTqq8HMt/27gXOCNYrBvOGE8t5iX9x66QI2kdfytkX+IRwkRjYyeWbGzQhuC
HOZNk1AxCjiQl7ubyYpqLgqF9SeH9LsMK+gEd278gsSm1cxdzWoztyDnNZGWJSo/
WoRnMVwEwDOrQ9SXBX6rkjDaFDf48x9GxN8AzxgdKju/Kd1o2DwcJkA+J9d1fIVl
1u5ck0l35IWTPR+J0SDrynGr6w/DwdWFl0WLNx0MXQc7OFSP0QfwVAuW1TZ++dRU
YGfi/D1KNeJHs+hZNvXNLNkEjDKp3yRxiA5qnyjpA/z46lcJpj4haLA2fCU7fz2Y
6SvSdmKjKLwAKDa/4Bohl9V/Tb0axjH15Iz/64/nO8CSicjEv+Oj6nHTm9WO5Oho
99QE7v4G44NJlVC6reLwyp1c+YvSsSbRxFn02Ex3l7qRdDfuty2sAFo+w3ocPI+J
thmdw37xwVnRkrn3GfKCxFpMTJHfBGQQ4aVxY4+wJ95VSDl3GlEdhCPLp9jL81mR
x/qJ95UjZxQ2ePlVguqC3GGNoe7KrLp3IwjVGrmnEdJwCrG0zjPHdGvnARDGmcgK
rMp+HPNSe0r18CzJSBtDbfo+7nDfl8ENDkGaaCvXaOn3UtI3/R1zZPOQIfg7rTxe
/AngUdXC1JLoUXhL29u3FZHxmaDJLLPh2dEaSjlWcnP/yzaj5504tGLOh7atp61Z
t99ox4qom5PIJcUkOWby7yODZJb87jADKtuWwmyhk9WEOhGfhoTwTtHRg+tmYi45
0Nx9C/u5KdDLVvSGvD4O9sXNe1M7BbhFQjxebrMXQbFXAY7+LULg87uFikjsodmd
J/bAJqvFf8lazANUdhrp6Brbxxmcx7po4ijABvCHPzWSLz8F8/gy9i3O37iFT4qr
Rp51Eii0E4Aay13pe3awtQjHlAMBB8zCN6P2o/m5QKczO2/C851/4dxjOpdjPz9f
XFL8XNKC5nyFB3//hoS3VyDb/rOmXHQlOGRYlWA5GPr1tX6LtqhKV4wy09FzQp/F
4Mp6R/4hUQE50AfN+7X1WibGBqPW6hbsbx00Gdw67q9VCc6y4gdKEhCD3wHTpqja
LjYhvQXT14p8qT2z9CGXPelfCRhaunxwg9k3augV/gqBshWXoYA9I0msm5RL8UIl
AsTF0HGExam5SYzDnJfkGPS/JwtcQMWGE1Uq86My6LHULZ3mM0fJ+ch9YilbG5kW
asYeJIqmlv75OIvFaD9wSykYcXoQ8w7wKCnACEGey+kJSlaG8FK0yg1h/L6S0JC8
1kU3kUN9ZseZDR5/yle3D0RSgTJnOn4CL3e7ZfY3wxtOPx35m6tV6c1oHcqa5RuX
73GRl+tLfA2A5+4uEZBaTkelwPqcs5i/Jxtwpu4/fZufniop1baEduoc/X9VkSSf
+ADxWAiWQlfOkyOc8MgvFARafmVCDvC/3bVOiJ/mpvmGvLoJPc9bfRCvixWU3jmc
rBPIz/XY1sQ75F3pb9cqE+ucKpJ8hou3xSZHnkNmoy8dUgOdNdisdYtsYeqABYLy
oKTS9ut93v1IMJHk341Tf87AcQvVWY9b9L2iMZeUs7a4TkpZJYFOnyUzgT0S/858
5OCB4I1BFUhglzmaGy0mWoMfmDVkNApyhzObXGLVxR2ShAuX7w5U9HByCWMmcBU4
6amXZz5f7GXT41c0Q8ZuF4v5RO/h34z+6Bsj5bm0b6+Pt5mZA7scj5otbK0nwBKE
JuGzuipsfx+rky3UC0A2k+rFXAMZjBTcNI5gdAd3F4glQA3QZvb/AG/JrLMVkvLP
6XpI2cZSDsqhCArtLztJMjr8YFwC9/7OayWPFuK2T+0wfRKboT/cNm54ged5AdLx
wC/joAn3BzwvBLq6ESYpmwBXcNEhB6r7bzrBTlr2JfIy6DUyDyfFtCpb+Bw+auwg
yRqH8NHpunGSq+JAa3zi59ncEdgStKrPjEADuvLHAimRApFJ9mpkQnVFIBHTMXeS
aF2iwODC3g2uCqx1FH9+rtbB93GdRPnBuFToqvpEGttDjCsiaZNrdOP9NIkotTIt
dJ4gLYV7ToTlw02InNRXSPzCcU55NSzB2utRGoQcR9HyvNy9/hOxD6sN+QQ8DORG
qJ/Qix5qvOJ1R2DWg9hNdgM8pTlCa+KSFWS9xs1GHd1eThRpT4epXofnMYyYJoiV
63ktFa7Xi8tcTpHXy1AsHv4uz4peAu8HMCXhulRWeYbuA7l6cJgdZWrI5atEV48H
IO5vHNEKhCh8oTOOQ0Sd/amifLwM+udwtB3/CEAPoYlFjqZypzdk0O2k7J6Xjs0Z
2tNjnT6BfpFcb1kl+lhpXUiWEHE/kRTGjrEYsrm3JUWmWWwJLGU9hKnfdMWj82pO
N6HpiVvVN1nGHqNLm6JlvLbbY4wbvJrxzkBX1qFI/zaetR/sJen9n3Jk3fvVCAY2
vY44Gmwtuq56WOwhP1COC5rkcJK4TszDIisCjn30bLMONx6rSyF1AsvY92LPIRnE
2r35wb/LtUQFwz7GTKgVJL1kujjlu2MjoXdvN00VDL2PbiKDApi5L906Ik50hC3R
XQP8Bz4Lp2XySIKu4FgyKHzxNxxTyeoN5fr2domHpCqWhu93YrnnIWFgJcyhNJQD
nHwqYTfNzOx8uXwS4G4nD3OHq7GK8l8qqhbh0QI8nN0bPt6I1Jooj3CxMxh0S8AG
BxxIwa2nfzEOQVzM1FP0gkJ9DywcpQqsnPC2cEBFoq9wSZP2VNdQVqBUpb/EEM7z
3vb44YNBWluHew7buhg12Qm+Eee5YgLorBV5nRf5ydxeIQMMSKGJ4uxxZFnH7n90
DceFlrA3qyH59RN2BupMyl00J49YqkJuPv/176nnMLj6eAqX4nCX+eiySDcnEJVA
X7xC22Y6V2t+6WmxK0FJ/pZ3LMvKgjh5RA7vv6rkXCYlAS0S3SXX5D8Oto4kx2s6
aQjc3laSSI7u6YQvtiTHqVj3CZBsPhc5Q+NbLvF6jooxTJ1kmwXGVFIrlq1DQFSA
d9pFJT8A8A5ZH8ujuv/2eqLYqAjIWp6r43+UD9B5MY13rfiRhj4ohCwMhshRkqkU
HSMFF3MMGsl0bdCWPo6ta4YAqr7H1V6K0krEfsooxYU2hBt52+FDApNjGF34ma2e
S5j8eAi0WAzi0xtS6DDrWTQpfeb4X9OWCGyIVyEZ+oBlfwZxQRYUN3lxhX2dvqb0
hXljbABGe58EsLmbjJSBZ9mRGH+SjVWfc4elSLd8iNTrVE7GRg0f7bKKK23oJ8dN
y9YfDwgBlQVozuvjtMjhsQTP2ZdgStrW5wYkkDClfBwxiTtf0Ve/TaYARZm3i8Uj
5k3nqZ0rIUBxaq6b6RRtKP/8xpbvhFjeMpuAD8vx9SstiM3NUoxkKhFafxGHOcGI
x61IvS/aTf1cDGrYfNfO5nUgOOUvj8kLQHJJJRs0ncxAaY8F2n+qUhVyXqhmhlGl
xj3b11fdkem5ZS/mP+k4H7wvfFi+ohPuQ5ZLuWWqgKx+YR8q3LuZ0U3n+dWE43pd
5cFv9pIjwtk8CZ48/lIUO+XRxQvzHT9hDgsauQG6mrQHeT3OSLLzMaf3jDYLkKxD
FZBbnXEL0PqU71wvbTQtQvNboBPo0nyC+mSA73oK0DWlerHDE2vxQic0CHSwKdFA
93chXkFaN5/9ZNYGHxHMXZcKv9+lTT9Fpi/g0u6VeEbebiCRij4nWqosoTh9O/w8
TDu668DxQUPiebdh6X+aH35rrBMegrNB3I5Ak87h521INOKSB+4aO5UaJMghxyZ1
M6Y+iwqAzR+z+V7Yd8YSzyz2WIjS5bsd6hJjdVYSk8n8207BU/snGNk83oae+CpO
ErIxK2mawhyOzul1hr/C8svHZPDk06XmXiRpqmgTZ2DI//WZxrrNIJOxzgFUCpVU
WXHW+hEO+i3xXu1QD1D0a2EHsyVxHgHB2iS+/2Cm/VkXdHhR2pg7M7Y+4P3NtxCa
pEwYll1IMzzYywS+ur08LLEYPGvWgOVIYQD+jE17hGxrHsCfunEo+VmmnGjAVZkc
OyTZS6Xh9fLgK0Go88gibwHjIeTvN2qK91RhY56DdGtUo3BPPD6N7DVDe0rYbH0j
/3ZqTdfkAZeTzjT8wtQ5P0qmJxVU7o69p5H21kaWSspSFh8/hiVEkMlPzuPAdzYm
IloUpYSLfyUFUyEYb/MfAv8D8OMvvbW1QmGrnfibJiAl6s+1w9Mx69W7UDAcQOJR
Uhdf6xWcuMZPNB/Ckc7dcVoPZovbcJLMrDkFjGW3bWPswePmNuFYEHb0/lJZKP2b
DB/7lYZVhpwUd8+gYwvlgDBf6BmWdZq+kzAOUuDbT7ASJinorBfLXKE9Mh2WJN9+
boGTPp6JNXFA50G39MkIWMAzKn/ixLlzsT8KtqrSm6lko5Q7w3kqtxY/6p1Rn73P
jJTpsnVZU6yAqPYEaEp4kLZClIA7q+K3WJzA4plnN0EbHIeOFSOvSN9x16F+25CH
T2XWtJhAWPBaGT3IWeItqW1Kh22DksVHY6S4zLT45PUUEAmW7y2FVZC0lN9+gP1c
pMqu5GQPhMYTDCrkVzkONEgMV0OVj8/ur3jSaLNh0wWmAbHojXhhKkusMVO1ywBz
c3NRsBHgC3ufPa307eds8mSIpR4aycrNpIu+iguj1FARF4aPPV36lYoW3Y0Cih7w
g9aH2TUXLMAwNt/n4CkTmrmm7K4oEzLXZGuRC7ndpUfN3JfSC9nBzwNuudpcn/AZ
ZsEYIvphaYKaOaaYcgp7gtiITlNfxdfUIDJ7P+2LSXgksmvWz2E2aGCAswovdapc
GQMHZ70BUOAhsKfM4Jub+55iRCf38zUh7kH1S0/4OkBXXuuxHrS3xpEggJKBZQU8
vX5GcHAij6YtyXyx7q5UAc6SJJ0o7JTlSwvTLaagzTPza5oiw42B3AagVqWXzIxT
9d+1/wUSblArMlNNFrxY1rAACxZeg+1Hpl6+kiB5zc48YxCJoQcTR43GRu6WJf0k
qplZV54n8ckQj3jcu5ujdS6fYjAxlz+B/oDe5XRmJLIxMt27405jywWyvr1oI3vk
D3wbitP7qEqiOmD+OA4sAUD19R9+nfVc8f+OF2eiUJpqCSUkQTcqulTTSN9SMvYr
Z1GbCxnbWd3k/J5vY2J6OZLtKieL5S+mgyV/z3SSeeMOzU0ntImOmUx9hDFX2r6A
lOlqX7lez7cT9KMSBFmi45a1cUsnqJ+SMu1kF/JAQmCxoPsM9J8i+znkiYb/1tlf
`protect END_PROTECTED
