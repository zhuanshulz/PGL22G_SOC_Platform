`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vA/MLJTVY3cyEixgfE9AIKYl5BFcYgOkjmOkPQCMPcGeq1F2huI9fxWkhIyXuWIS
wiaUdPxex2NhpR06VshNAyhonTtV285Xft/hEHcUMbL1WDpf1tGe/DCCuI9ebhaG
qpc/pBzTqRopXxqvbuGFMPU0Z9elgQ5EhhjG4bHr2SJ/8D43f/5jibbzs3eMJFOz
RNaNgjWg3iIurFVm+lHUKeiKDr/Gje9G2sblG4Z1KLxIKxL1ZaXtxyJacnBuinXH
skLagmEEWQTvOkh5+Q+yWnIGm1BFuKlXlf4BPbp0H46Xk37z7X9Mrk4raH6Uo7Fn
6VeMSgoOQqbFCIFA9pgVvkm+xBYFfJIg9dAs/2lNgcT4v5LVc0qxt0wvgd9QlXNw
4vgA9xI7kpok6Pw6F2Dozkf8SHARsA8h08RrOb89MAAYJsZ/DOsYXAUR0fXGA/Zo
BP6EQj81/u56LpPFWO8rM/hS6pK1MBWZP2/8W7m7JHtQr7DkVv1vnV6DnxLvaOyz
4BWG7HGMIImocQZEQEoDHkOpaoU/SSakNI45EFmgAxI6dKyqVD9q7Muylz08DDeg
BdPbUtsG92zA1XJYq7s7hv1mh4jNbXbVAoIrzdgeMR2yHDmdKTEdu7zKRCPzS0vi
DChPTMPYG6QjJ3ZllzRHN4Af1hJDo7A7/TeR+bzGGuS8IJDXEJ6L15YJg8im1WF5
JF1OEHX4kcE8mOIrIOUWTYwpDswrVo87dSFJzFgerRAreD+ZM3+INZCX0/SRTran
3CgI5OXqpqWlP1/H/gJZOlKM/3kRqSGIb3OzEACQYaYWbqJ5SvTMtOHpmyAFX8r9
T6ixdV99YYHxaUucfV0HK2Tlm2v8Mcxy3GtWDfT2T8+rr+HPzou+FXGb6Ii9rVgh
pocRuajdf7KUod8ZVFUZRbLQz+9w8KPMPMt4VOYLQx/gdbjWuu4ts+9gE2DBUYn7
GyraYs4lZSE/jg1gqJi7htp796BQXFvN7JaMAKYDeDfv2dSJUZVXBsx6g0BzgBr6
qUN7zRpZX4f5PmXKbMPFm5CNlxv9Jh+IkfBk8XSECaeBwS4T59SAnXGVZNszhB+5
kEd1hNNJVETXe8bdsXqxjOThzXVeAhtwWV3i86hF3z7/R+Nfwv5ZNo13pDKJ9k5E
oIpUmUhfyxZKaCuS8FuXiRYJsnbeLtFKNcAIdgT8wnC/qY5Q8DuDdg2I345g48aU
vgDlQ4fQFuYpO6/yw2d61M1jjdocwriWV4Jc0nsHKaLEO3nnnhNJEhCAC4IDc+bY
H+mpns1b/wxdMFvpi4yj+wqSfCY6Pk+rkQKphMexulr4nFML98STM0M8QjUrMgHW
Gx4eqg4W9RB6y172xK9M0K+eXPshJKXy3ySS6+n+LcPf0RkZx7TI+LArdWNVdD+5
NTzvJhM5HevJlRb3n9foTQK7Is3mVVrwPsKojJ2Py8Q=
`protect END_PROTECTED
