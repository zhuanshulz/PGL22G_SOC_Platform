`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n29IQbgoyI2obS/ufwkPArbiZiz27CoAVeeT3QdGvzZbGZJdzQ5262LevGFaWGwJ
PITWBeOPx/p5K4nRr4zpoyZ1VnCbjiR66KfJseAQPJDqBTdqdUsf9juiZTyEl98e
jHxwnJLDCNf2RL48LsVeH6+azCC6/XwapVjJWNPiK2Qh5EqnYKQEp0cPoyVNSS//
9ApWgCdp4/xnxTO/6K40cQ661DJID/EHGnUjPG7K4Ye3VouswaiA9Du9K+pD4iOO
Dfj7lfSSOpPiI2U2y4Wq6YSKLB8wD0L7u7tsd3uz4iOcv7sx0pluwaoWEgmvmhNc
rMIuF1bBdgHX1RHOyy5TlYzZDsOIikvLU82OZI7C1DmAiZx71Y/rEsFUEsFsIdR8
gsAOj8WuopVeL0OO7MggnFMRJTcrqNv9f+bRbbWl395m/NnvTOW8jlZGBsYNbBte
QVGOAdnlBMAINg5oS+x03A3vzaHH0dPhtZoABJrD8qWcQnrNpsMOTs90djyMFji1
R7knI9+UlU4EZp6I4LEdTrXdaH4YKK239kA1f2PLSMJrZffplnqpLUVaCrYIZLqf
T1TMzwT6YYJhe5q7GfktbZc1p1or7+zQRGjNcoqEswXy4Tt8O4NB+IXwMYYCcZt6
b+u30SsEa5eeH0wKXgZ3qOHi6fnKEBKTZsiM/ZFXpsQ3nr0uCWkYmRhGwlUDDKqC
uOCgAsmNLSPHAQcnRSG0wrCCOy9Pe2lo/sDGa9SeMZ2thFnJFSEi5bf5dOqt0la4
6SorxJ0V3V/hBqzWUS9TmEQuLheUoA4Gv3G1e95JDtlz2YFMvXR0EoMti6c9xQMk
ohXJ1nkBvpyoXVTRqzdxuoO89qpIVpI2qrSyyK8M4ONNBVM5vIU8nyqhXXxca1Tg
buhOvKyRcjvLmIx4W2D8Xqdyrh78EOkqAOG3JGpSrPn2/2NSNz5aiECLlv0pURpg
NkPPR1YWo5j7kb2l25FG1MN17IusQf0ko0bhph1EfrI3gv/xZQutLAEifSy0+mxG
EmixXTkrDJKz58y9+Je/9wT/4efhKsCOCVkoShm9HNhdqh8C+IgpvaGG96Qvhl1F
FtbXu/pWD65xM71S9C9MNT/7UDtLu7u0ArGnehV1riAF11oCW8Z2ZVG+HLbnF9x/
BtXn0UYEj2NxoRm6UGn9+AfTXmE1DyrYwQ5VdaFKk6BkWoPW+P3WqcUyW6+akABN
hecRj7vPJcXbTRrA+JB7cT1/IG6mtbJzJuhrdOtnAMmiscIJi+SgHgUu1uzCtauk
7X+/NV5Upl9iYc6X9rZipXFMzTy1qABV6dRk68hur4zVGHVKzqpJf6ekE/PfTWav
r0zY5DHVLgsVe5wBESc7rrGyIbj8gZpdfjPxKkhzxnpoQ0U6cq9QFzUgz7OokyIg
AM/tHLsY+fMvqXs4J4qMexpWHqXHwwNe0vZlbLxYvE4IbXONQo5SlchKPBzSpA5v
ES0SVukeUPsWesG5kCzFIdHj0ahl25VWaJoY5kg3xxv44LUM0ghuaIfxPkfQN2IB
3TmATv1kJ5p2TLtY88MAP1564edtpWckhykj/4dIVmAN/GhuZy4wry8bJAfOUsN/
38L1QdThbMrsvYP8SWnZsXm33bJ031/wBHzPVJL1TnumxIvTQDxL+Ah5jN5Nj1eK
qT9Gin9QbgMjFycGZamFLLdxRiCG87JY7k2Gt7e9xW18XweTKhoPCeqnMokdDKgM
TEbmNT1gViUC19OYKLNIbXqXux8dfxZjmn/llh+X94l4AbOm8ihF12YZHJ3h8drr
`protect END_PROTECTED
