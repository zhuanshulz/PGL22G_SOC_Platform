`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9t5Irxf6orZMaQdH1HTbdLjf4g/Fs+7nspq0FfSz3YkINAJ0KIyOMKmzqu9PXKgA
mQCt6WBEqfaS4lDUjl4wddLSnXlnrDWfinQfvlrPswx8SLY23XxEcV1saStUN5nn
34+y7kyC6Vzro5JIwO5v28zf3ShlL5xOAewsrhI3m3U3+UqYSZsqtE2u5Dv1h2CK
IzFRHKur9xV/E81swxnXkvLTrD83MJH63XecZ2QdxyTP3+0SqdwyBFWBw5kIy1vM
G2VRtU/EWF5w8XKNvpVFGzfqliuYwQ2TRDNkcOQ5CLnB4NxG00K1l4U2XyPoMUn9
XtLomuEPlFEYdZF0LX3uAW1lh7y5vEjD6sqoPb25HcSK1FcT9Ej8FqeePuCXCWiw
UsfYJBaGB32QnDPbtVkmM5ZkPGTsyGh80zGFY/FFsihM6gzoDmtYa+OQr9Z2yHjX
2e005oEH8ySWBaF3yPdkV0r1ieSNS+sqsOUu0DZIX7IDieDLT3ACRUvqb+6HKMwH
pcgBTDOVslELa1hjmvwh/d9oWkNo/bCR9oK8jNqGC79J2wmi/emztoJD3pyfJqCq
1lorD0SknJN0DYyk1eg9+YYK6JZEmZQxsGzzuZK2wfe/OWZaGSAgqdg0jD5HNWe+
cpNIy5GHyN6p2kl2UhB17zYhpf00ATu1ijCJM2MrDCSytmWoyRSUlWV1sgdKLzz2
8Xm7pFTw4KTNG4zuRmKu/cV9GdKnuqg29wQTNMR3jzuzsSvZ8bGjeSyDkzBagcz6
RHaZ04yKPy1rzAZsHMLTcbXlBk0uo16ZSbjesoIu/B4rcNb9YFSuyJFMiAomC5e4
kvKxJ/pLB5VDixnr/pAKq1DG+LO9dkTuxTYj0q8WOnLAKO0hukHoc9iu2Cv5BoHp
6qiy1lGrqXwZWaYXBIJ13T+qxkYwtVE4RLt5h4xaovFwCWaNruUka8j3GlPgekhC
VjDwLm/2KqboQ7ege00FvqT7wEm6NG/RGpv7KNu02Zrxk9WuY/DQ6jKk2xTTN4YE
ZBdyMVFL2/rnAEikP7Wu9to0tpFfjr478S7B85bPO+7HHFuZ9FYJamUvwiQOtuQE
AHbVs7Remr5BMAzGpyH8Bm1GDiZKsUjJ2kr10KQmBrYQx5WKwKxVBK01HHD5qWvc
5bPXfwPrxYNRxOFBmiwtW+kH9VJNOkxVEq+puVJM9As8uZO+fJpo0ur9Vac2Kkq5
8ikXOYH1QyidVeD1r6dhtQWPVqGD+4BRP4b6STL0kK+/nZ4Vg+JZ3s7bx2SgFp6B
32q1C6+4KairS0kxtcJ5eECNHghXJrU24O3B3kAtu4Hsxihc170NlJ5QSVOHvvL6
GW4WfzSxRBqfRPTWPXnI1J/ehfZr1swRN1/oRRyk8nA=
`protect END_PROTECTED
