`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zv7XGWG+UHUiDpAnpILE0ipOOP8l6do4ElaJiF2RgZzEhZeb8Ea7OEI3QbRTxu/n
M17Kzy1LAM2HYJpvwu1OzMkjTom10sYUwbu477vukjICQmCKi5m2ZurouBCfaNVv
ibt9H4f955KWO4iHF69gjUQyDtxXRKn/rZbdw021nj+pCsog2sS9DFal0otY2buK
on0eui1vS7nNzmX6Nbj84ll78vtRqugQAqI7RcS22ZPSkGOv4i66zh75wjzmNNyJ
fVaQNEVInLEWYRuRMJPnrgGC8CMWhR8tuGUcSMcRZCmt2h4kd040ziC5y31UDujb
KaHNc9T61lzxyetMIMQMpBb5Xts0YZoTgCDWqp9JSj4unQGh40cFvlNo6AK+mq+q
lr1Jq1hcpV/2JbtdB62aMQjL88u3EWVR2GDHcWsWIZ78j79ecqNmLfDfchpvmFQ8
sUMra6l+PWUwbNt6QOB4mRcwxCJBvMPQZ4uCarrmd2cNedQH/mVepkkaGmWkaGC8
GYNcm96M5AXnz96CT8cjQSu5K1j/nG7EM2SiCw9L25xrMQB4Bi1JlRCzVx7DsnxV
7Msjm6JJCaGnBKUncXr9/g==
`protect END_PROTECTED
