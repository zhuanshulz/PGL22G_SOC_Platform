`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/mfVSMHkewCwdlNPfcMfNMIp9OCxABP6eR5VyqrVKa+HyTyuIVtPCm/+1gsRYt+l
WX9HT40FKXwgM1Hmy4kPyqDPTnwCZ9dCtsBAsUozmVlSnieYifv5pXAcJATWBViq
fxDOfcwMsVc0DjjiTtN3PhAtz5QMM5iDszG8bA58p3AZCrArN9oZFN86ts/MuI6s
X2ysnOKhb//a1sINDooJwd5IY4RKES4ghGisY1gsjN8vQynzLudQHGMTtKRaA2Bw
Crs02UXzOCLFmbkH5czScRqGDj7VElrQAjEbNkJuRxXLNXmPvwYyTz+hF79NotOL
qnQIQkACSAauZdyCW2Th03hPwMN3n2v+XFnnBSauDn7ENpHbYxKurwoh+glm8dYT
VvKfrCOuxuS7gvTBqFvqYe5EHOAXsW89/y+/zmTLiJbKiiX0vknKSNC+ca9cOk1R
t1L+m1mjNaocW+zPFrdlUsJxxwvj23AYH5F7e7iiN6dCdTfjz+Kjd6hSxkO24EP7
sGHYl6Dko+zuaWwEvnxobuF1MSAlz+si5Gq0GInJN6eejOOxaDNELUVqUH/TXqLg
pQsRwVAfn7GD4B59evlfWgguk1jKAlkiTLJMrzuEzSHdQqC5FMCoxe7+H8Q7GbXQ
TZEnNf91kHk29ZlNeChSb2PBGX1hCI1GQkUCdmXBErmWed40upGZIPtVenW8dHdb
6v2f7lAxcYQBfvB7EV0DXpSuPsSfVcHFjZZjaqGYRr7REfItrOM+GOJSuxzUAY3Q
rDtH1AWv5QZsOxtqGPDuDIRvPcRPOvUHx9CbWLmlmma4qT9IhSWr0omgTQ6Fb+M2
ueseu4YCtR+P2oGMc6PLOcnXj33ltpxhOGfNhjawEBmgQRYFu9BVKQ2WQXbkjK1X
qHLr2rohatmZXs8PgwWqBb/r7ogdsBLv2EY/Pw6pyGdYi7yxyYJN3gHICyCdwbLT
qgWg7i/Jmh1Suzm3t6SRxKOB/8ugXdnzDH0S8YCcJPcM/4gbCS1yEHadx3cq8WN9
omeEi9EBqyURHEaUSHlNRQ3z+RMFVlUhD2C5nF0yDsLHVeY2nxaUop+W5smnfAXt
GVwJf6aHSDXDz+LwA+1FSoq/VOeD5b0yx+C7zg5STjOGIteiHMeacZLMErAV/spR
m5DgPq9KFicODJGrJHHkoB5OEbjjofrVANh1gsr3G0pIzyRGTt8Nh46ML1UweI3X
tRCCJ/npZzYCxW37YdSF0mbesgBGmZVLijvippxG7MpcrbVIJYbZunOViv697X+E
g9qykccZsrt5ckw9ccM1rNSAb5+9iXrvONzh3hFRcG1ZnKL6/aILBxvIL4Nnx3EH
ZVbJqeLvwMKYLUjIsCrjBZXa5LlwuMusbG440ABGplFTvIrrdoLB8o93OWjx8ZOn
9G/EW5tQxzWmPwbghbQPc3JcmjBbpNsDdN1Ph1zH1BpCW/oDYaKBL1xtCXJmCCbk
ovqRoS76bFW0ou4FGBrUzNlTGiBRYWzeox0eEYUtJlQHBqMGh1YkAqDj6YOZJEXB
IoezmHgVRn3siy0kunsI2VfpNge7JLRbpFmR4p6xvOcKEBZUdppVVphUmountXJF
RieTaOcy5cfPhdiZmIxXHDkhyX4D4nz/KPeBfyccUFbI/9ed1fdYMpjQ+wgdDBZU
qPl38vTZkzmAncVSC9FNzZPntMzQSzf+ELtE6O2yUy3uPxnxyWn3KalJgHEAJ6pB
6rvqkfqCpTtml8dw1gXYy0BgPcREk3JqbOrcZlHaaLNue731Ed5WnqnJx4vnyTmP
jnxQGmp3OEaDp7EbopivHladJ7gSF6ZB4Hgt8Jlj6/fPiCk14IubT0JQnYCQvFBO
/zX2KIvqr91ddhplHN3NWS1h/3Ma5y6+9zlYhdP/mp0/afDGywQaaPh44c23CtIi
Kuqg/VKB8zhrKSYq08tjXDn2UcVg/SwNsKfzw7R6kA8GD72nRn35JPwGXdPlMwcY
wq1LBtRRQShapZ5l1XEultagXaAYPd37YHWJRfcnRNiN/ofWeTpSKJ9ukxiAivZn
Yh/4vbrUpN3bGnXMKjEdY5zXgLVKEznSWAIamolztnG4Br2CbnmzgJVtMy0uqOGf
rw2wMcrbFYw0hX1g2LrZxQ9MQQxxkS9M2HPT7DoT+VVdmnR+fQh0K/r9TRg3ba7A
D02umaVWlRNx91ujbH+yYdAHZfvI0BQk9Y7VK4PoeQCiRJ6VPZm/KdO5zze/bVSi
mFECWzlvTdlbzH2lk0+Ghrw6+FZ0sRwQOQw3nKNFXFeo8tekWrWMhUYkyAE3YI/j
e3A+v4vk52fCBY8pWesrFbwO7mSFyd5EEPoCS+CshY222oxcqBx7ozRprn+xUEh9
SeNl0yn/BBBoK0fe718ggIvyX83F7LOB6mOaNEyFUDUPyxEkSPurgh6EOlPLtMEq
YJZjTHKCtg1Oftw4yymYk2cwsG5KI5VbxTqfCJcShlHwBVTCQOFCNd5ePU3dUxTK
GF2VjszRO4hCYl0+mDygTYIYY5k7T3tmKWZFLQ5i1ZZfdOewgcp033k1Q2HzH6EY
+STDUbou0koFntmR+yR/g5krhAlB8rnY7hJ6sRKiOV4lHAJViJC+xZClpNZ50OJ7
OkqD5C816LaRL8xxchtuspZfUzd4syN3XteSlVqJ5TUrjQCOkjPGPdAiQHunmwFO
cAf0ghl7f/ANmzCcw9+b7gyB9yofASlvmVmuoaawYIduZZchIsZEiNNJKhIgoIvL
7TMJLK1uMnYPfGzwfwvxwCI327sOFShslXFxm+LlV4kVPxTCWJdfFlcoppagNyiP
2BcpM2bIDT9GxbMWZKwAaJ+yIVO3ff1ARvVYBfZ1RK37vIFg6mfdXt7I9A4qbJWM
efOOZJGQg5v1uy9Zo7CATd+kTk7yO0A8FlHxGANq1xuifBX+g5Y40g99TOYfaM0E
vPtihO4+BLGzG3vmpydOGoiWZi3AqQKxm2RP0tD8ZaA4wmqdzkk/sW1ph6YuXlST
HwZHNfh0Daxq2pjo3+b8Fn2LqFPh0e2X4LgEMt+iD23CszDt5yeLGc5Zk0zTPWiW
rist9OWtyq9ZVz6JgYKTL2i0s/ly4VUbKCxmst0XxKd490Adlk1JhxMRiCEXwK7T
1n8RXPwpCovqDVzTqDMmCfrZpzhCUdmk9JELk5+9qYeUETrphvzxQpBOBNIk7AX5
C+ADfuAOa5H3wmre4bCcXw0GmxLSc5Vh3Azp5zhvsh7/oc78N2PdR0cHNhm/QK5b
mH8OZpAvhckQqjlrkj43qukIeADq1dLqZ9o6a92m47MtnTxxlUvmPoj4pG+Z+fdB
ZHDTa7JfVDszZ2PRViqa7TMrfeJPdU+Rbtz3ajEA7FQnEOc1qtIg+YmRrBcBEgpS
pa6v6RuYI96MUe7WDqm+tjb8o7XhPBKi+IM7nXwRPbit+vzkWn0UX8gRzNpABwvy
eVDXZ29vmGqLVQQiyOZG7yNwh/PB3A6L+S0edPnh5Jy0LRqWo9mvCJBTv5sn+Z58
j+dHRE3x42AfC1pUP0QOTclCVLiX/nErtA/mtSrakscO4HWrTRtTw6mv3DUBYTIQ
RN0uVy0SuVHJh+aGsXAnE2kor6HRSv0lCSuMN7I5S6VWNqz4iBy5NEnSGxAwCJWb
c06wN9xdHzGqugfKm9NwY+WqIaGOSOYdpfkDuuuzvFRlwpM5IBKS2fWKt6TwonvP
cpIINqebxQQ4QPvUBvZqt6IUn/4ahsUV//X76GXTd/q3gtkhkat6XXhEGDNGEpFG
jftLDKOuF339l1iMOV1ntr6aXwpHEhAotn63WeRKP/3m5VZCZcmL/Y1qs3/77q5s
sKwNbZdRTDR1y97kEgR/CELBv0oghxEM9dovtfJj3SjIb4q+o2eKKzM3CDQRRHdI
5rCWH4aKYIyxWzSFbtaSMPvMutFmmPiIimYzmDGeAaT4J3GT9AMSvfGWisymoorc
AnXInYKda+yKjCBhHm+Noox+XJBDc9VYbME72oJcZPjJzMAnJ8pg/gvL8BoefjGO
3MhX9oJJ57jfrZQRQTZWcvtHkM8pltUudHiPg561D32IesNQG4HAeRZTnlCRKQfe
8/xFJtvMwNJlTa1P9G6eooJihX2ZOjm+OeT+u3qKp4op0fYaZSqiIZX62sEqBg9y
8WR+HjNpE7b72dbzOr8n1dg3iRvp4TJ2fJzDqIM5Gj5iweD8/DD/g/LHdTDWA2T4
ABdTJs98Re7EKoqdoC7bFislfFFQ707j16ZF1zxTkAHP7QgrQE9Qz1KHabt3L+v9
uIPBItSsu2+uuKfV3XgoB/aTTTDXJ2gtlsuEdGVaJAq1S1vo++tIfv1/zt/NqpLf
2sxC0N8/abAySOrWYtgVixnRzIQY5r+GCmGSJkT4adGFjduCHpkIP6Qh+Uuu9G2P
TshFgjCdp2r3x6+VIs7npjhbS0E5oFUJtSZGWOv7tEYB7yWRexU70/K4YxCyosPK
SBNojFxZSBo3RW3OJTrv+8hr62mS+aRkn3hjgdYHz58zjOS7jpKs90CUWOOIY6p2
OTLCSFDIp5gDVr0SZA7LkfqstvBeyKxyltxFGDf+iCyvZL0N2OCX8MWKWEZ+fcRe
tSvb+4FD6SxK2rcwBfSM9JOLomfKIF/VAKd7oPlCfonO9258gwOzAPe/w/KxTzyA
9ajJLT0Ivcg0LYL4ca49lwrQS97jrBQMyXoy16oYTHD7v/+YdsdUiCFv4+Z5h6mn
cngleS6ZUAfyaEz1zD5cGDYByyVZOzMaD7l3r4V1Zh8xSatalQAi9RApu0Efb+ZQ
79/tpjgzRxUNXbAqksa7oia1Kp+UP9Ma4SResggNYBRabDpmJiQqjpJmhidhLihf
RR5eqNP+LymfKKRhtX99cp/xQAQzsq5g7scWR7xHXBm2QWsWQXUGIrI4pCKPqz9B
jXj9owhUHpkBhdF7zAaMuEIvJAqwDBYy/Q4s6jLggxsY9T2PmZDhaPGuxCAlrkV5
ARbrFqVgBgpIz9C8EeOdkcMhjM+sd3G6VFIYlaE3anW8fqZb/BoJiCBe5QD/VdkD
vIJRFM/YdgMNAnypyh9ghyQIge20HYzZUS6jn2V83rMKw5UzZ+ogZjSVQAwt1oEF
qcEW0MPyrPijf55nLbZsDxIY4HaO+TcCyQwa0pCUtQxgIrPKlvBF88W2Kr64GT0Z
TA0z245IlvQQb7u61ix8/3l2FW/Ju6WntoYibnJoYKeVR/n8gQLCxZs6iTs55Ooh
na3WHTiUbOgn3VvaxEsWrfXBfDBknhPB1DDU+5GbRafIuW23dCm64kZbcAW7dOXF
YXoWBJi07t/LPIeZZvwG6MAvdwZMmwsJXhujALwEp3dh1lnnEHfGvOF8JJUEK54u
LMIjY9Vg4RrKydFJ//NIWyCkJZZ2EDdgnlJAX2OpiI8f9vow/CPoIShm9jPkwjln
PCRBnS6OBsQ+vi654K87ToHDP38MF1Op4smSICzNEdNwAfktLWXXIfDJq4JA9K8u
x0WmYglzDgImJ72E8ErxNUaO++oj/TsCgSUs4Li/FRtanq47JxFw72hZWxOIINfc
U48SPcPSTVBDtLAWTlH+Jtj0UkcUWJOesV63A1eWv8Oj7HtW9IhwfyaIY9r4pRn2
YkHXT48r6EzZdNw6MH9+o8ZCX9HeXADmjjN2bt4weLuBHXLUz8OYvQcQZhScObJR
nv7/JKtaHCIywcKWC7DTFF33HGyRkLVHoLB0z5meYXEBZzFsS9HUUlXXQaJ7kFLT
AvaC8OtVyeqY4YUOvI0Ds9CzvjBoC5SUxk8v3SjWQKMSToTYEnrc2ss4fxC1TBTR
6MnPYW6R2bImtVdWBLvNYnvlIdibiYBTgv+ZiuuYcSODbgpd/wQAS2D6eHzs039m
+i9h9hHmo9qwNKCepMgHTWkOT+4oaE5jxb5/ZXEgdSF7DV6z0tcpgAHd3qI0GGAK
B0w0gyBYCw5kNV5hjPlzE9F2ig6jBPQ3NPPIevRxJBq0KnJtt+WD7al6anBd2X5X
r3T9OBrSg/8d0TKIBzLy+oFubwegveFzaER280rp9AfM7SQ8N6t4iBvzfnkmkKkw
5jvVb/ENAvazFH83g6P2rFtck2at4GWRjdcY3rkcxE+con3DyH6eYVZozDfytuWY
4F5tHZRKdXptPwwCu3D2fWPukKYhyNMZL8BUut5uEoPJ37TPpq18Bg4aaYi5oH4R
hKe7owjX36N3INFqiaPks59XGOmbFHlx8HhkpqBXrz71Dy34AvBbMU9CbJyKs4L2
Miedv1Ty+TmxCTTmLUnrUDmcrL8LgPIpRAOD2fieIXsQDtYNrRnYsyrS2EDbBoOp
cCQuSdK1mHZy8aOXeqLmd0S+JbxHPBOye3i4YNG+rDFyj8YtYSZqVfpf8gJgOet6
aScSsB/i7htGqSFRyzZk8FkyORNEEe00yp1oUwufEtRz3vrWujWgjIqY9bwkSDy/
PMbbkm8hhGGSt04tTvILtYXXRVImxtIfV3r+tZp8zWSRimeT3ZM6wHAYbyM64Zmh
ymdSUuAmB9JAch9PTS0Bxz7JWN3WdeolvYab4J0vixySZZVVvBJKlTzuKeDfgmbw
9VrR1YGrvNT+I/FOZQpLPd7XwmMfZvkRjkqLQF8Q4mWYSfRONAZ2B/OYhAOSvjle
e0VetZqLFm5yzA5ZwmeQzODdXvvfsdQpFeNxoXWgNH21yMe1YBPMu7hqqiKn7I7d
BUssRpK56j5hyOuMG6cDvcbh5QqKH1sPfmvr7vzGRsEDGtYVILKfRWNwUvWgsEeK
5GP9zyo1FnKn/dNb5rR0vBwXiH7lpdS4oiozVW4HyPwkSvtvZ7dfoMdfTEIuGe9g
h62/zsi4Vdb5YpcxNqp1Oi597hxCwYGVnplu9aoO22aglO/OspJByhFlA12hL/Bw
vRFH5R+eWipIsXOMccMiqUVq8Jh30/0WTaQhPvOXOp9xAgfGxK1ck1mRIOSooirb
7QHFUB4VpUKFCYkzMZ0pVa7E/hf+afgH+G0XeZ6ngw3fm2gZeG0QYXvBRjfNe7B6
2e0b+5/2n2pXBAMiUk+mW6W08PETIZzfchd9OXs3XM6KglVXA0x4zawXNPOTod2K
rc7V+OW01HdbFCHL7moDcY5iMjMKD1mj8IdOxJfJ7YUkwCC2+x+cbyT4ibfWTjWM
OfhJUN6ki6lhOJV3081BMQkxqEna3/WqFDF3ilISREAl0GqAb0uw3MjtAczP1bhl
gN2XRSUo+glgFt3V9Sw80ICjqVhzr4OVk0rW2aXugAb6H20jyjw1r/cW/a19Sc01
e+YHXnO3hdmR+nYWbEQNsumLwhnZddCsAj6sZuM6fi8F1Q5lptmqZm+EaHDCtZjB
I5E1uN8Bt4CqxKxkKoajd/DejEIfRGcny7sv5r+DLJgaBBUdxRzMK2cvqb0d57dg
3Iq78WP1ZHPluvno52rFZBc3d7HHNJDgBIC2uNZP7iYM3OwVwp8rqGEoa9vh8UIM
drvMqH9yhApQWmMpY/PyYb1QtKfmAqMRRZMFv4gPgM5vzs633lQ/dvSUy0OWcvEM
VAa/eFIqS6t9s+c6mSsJvEovhXb7Z2k/+ZFbHuOHVK46t+0nR/IzwltgkwMQ/6GX
RrxygyAN4rfNl2cobhursmUINhjtvccQ0lsO0vMmi+MczboS709GyUHNDSp3DYTv
K+qJo7fFNd+zIHBDB+wvkFSkBpFzHbz9akQGEnWoNMat3LquLqFwp/ej9HAAn+Ud
bnnvrkcME9xqMypmz+iGFShgcr1Gxv72brRgFIDB/6xAwdvwl/YsoPGgvPNNmBcn
kFO/HLnKSAMGZENx/YmHXyGTGDH5GTyP3pHNulcgP2tNcffyaEOnQqmLgbtr/+/f
ptLh8pXqBNaBG7/RN4bYa+ZbuoT4NwUNfKkNDZhjIFRv8hKaJranIxPn8jIvH95C
nJpZnhI7Vh0Tjkgs26AxgU8lvbpM3sA76Dn126tYI+Rcjx+D+SmhUgPlkh4XNVve
WXEV3mMhYnZeKxCvtfgDbgiQ09j+km/1j27hEiP10HcTg06rJyT4Z5IA7lPUeCTG
zK6lf5kxrqT4tDSNnZ3+GnbtGmn5Md3/8juynWfcK1mMosZipp4MkLEXT2NX//lR
HGd8Q21Zfy2OWB4QSq1VB62pF6CiI/+4odSJhZ2VkG/KG2wOdyS/vh8w8jNv4dKv
qltLU9ofpdFhmCOT7wDGSdytpy2Jldd2ChCWcJoPWrVeFZRhqH0jEw9TzoU80Im9
JoYPGIwiY44eiIyDl3APvSOHOz8a3ou33UWiGZGfb4ZwYZV29eqCKMrrLA+51kUS
taHWAFxzMsyxJk/3fslgsKl0GoS0uJcJEr5yEFG/KiOnt2XX65tm6HYx9/kMeRzG
wd1Tff19Vk2YNIte3C61YOIEgKJ0XF0S5d8G2HrnvSMOrgmOCOFHpGudyMkPtIp0
dlxwcQzCRHdi/OPXjf4RREFmFnCu5JPAgBTXdLhWa5iRmw9CifFzE8EnNGCW6foA
SP1V9cNtYCj/7UMp1+4FLHDq+1SwJOpak0gm4dSEKoicbFda/lAlho0YNtvLSNI1
R5LmoqKtHtRWzbD7e57gpnv288XDTbDU+t+dexFbUShUQiQaHnld+6mRfPcrOwfz
4MmHjpYZnZcWO2SqDD++1EfcVZgTnJHI3x3VuVeqVHvP0vDBdW4kL1wrS/jvzdFS
GCwFB5arayRJwIP6I3iSA0eMxJunWA8jX5htl+1m/vPkqH7YmGlZsb8PhQ5X3u9k
sqhtGFQrp2LaJTaq5WaShKcn2io1M1a2VyYzFrHSZqw=
`protect END_PROTECTED
