`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TlFLgKUiTSANwNUpMY5Gu01l3PN1dJdvTTRR6LCnnEUKqSno1m9gamuozGTu4Rv+
mpMte5ynVTuzEyQ7UsEbQxfz/15pXNsDmaOXayvYDypXcIva1r4AkzvtxNy+Dk+N
DSjv3nYCiDcSHi2/+HmlEWYZ70dvCuWQOQ9lA1dib8klCGf1jM28zdzuSLahGP1Q
VSWkxLuOL/KwAeQ42asJGJ3GlxMmrwPEonh/Ghe+iVAcTn/h+2Pv4LWhy21sEgUf
`protect END_PROTECTED
