`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
te4k1O5IGpj6A8UGH8B2DLlJH9LV88zXrpn6EqE6jrNc4w9tMlrqVMH2HxsR7Qhb
uju/mG7CvFp72OlJf4veAq7Rnpdc7F+WkIByodpc5hzhb2M2lvfRKJXYixQzJHKz
w7kBhgFTLOLqSbBE8Ss143nHBeoXtu8y0Uyf01SU6a67kcVKYWWnwFBQAaD83Z+F
W48z1KxAsx5qh6y5e9hS5qh+fNpFFFLzC9ejfkv7Wn/7q9hU5uUSwGjI4DwVCxeJ
iN4bl4RDstJKILHfB9+pbaSU+qMqE/XE9i/kWcU2hRJ4Kxr7R36JsvPaJdX2DRL/
0+/Up3W51P7Q9/+dwZXHZJYVCewZU7gi3A3q9SQg/PZ83mFReBLMc/B7R2ERo6G2
gkfOetOWY+jwLbcyhHjHxcpeb0+vD0s8j/ph+a8Ayv8cyaTboB+PNR0aFsHji6/t
Ed+qwioCZ8c5Zltdpok20bYIhceH3nMbUzJxHQmK6HwxVylg7F2zPq+WvL7FfHKG
GL8fqbyXazWHGNlbUIHkBvuT9LbO7zU93eCbyH45/3M6Z7UgrYkr+/1icez+J+EP
edurMCJ8Jtvboqz3LUQM55NDnjcwur3d9WAoFmcn5gG/E0w+HYOF2YRRPdstGnKf
vxJ9mVP18yAyTavywLAhtvs/u/0W25lSkN60k2P8YNnczOpp6zuRHbxr6Plk6cmM
TopRCW4NOQsFAeMlelk2f5nb6n8yFE7t7WRt2PdRDhtC6L6cpdkMHTZXka75hGfa
MD5WGIpW/PZn93JG6En8LQ==
`protect END_PROTECTED
