`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CJM+j+dhGwDKK0IQ0DVnJgTLM7x/ZHrO9s4o6uTGPFDI/aIObL86hi01zhkE4Cn1
PQ23pOJGoC1w8eg+8NJ5hUH8X6NOOd0KI4aRZS/GNfQE3iKfU7btolesxEqwwoYP
9Edw3/mwSYJGDg+pDqMRHQ/x3AEHdk3H39DFwdx/ZOlrjd20hMLUuFRiEzK3kex+
eCX6cWAvQBEiwJMzbnYWoNBKLvyncwu2AiOfYTMcGlTHX09Tof4Rq164CU95YdL3
7/cCjG6KfxMg+4B4DxC1KXRiowRDR+8UjXtrrtJTxdWkBGxvESZdOspmeaAob3Pq
lAyS5yXtIwMRVbC/M7HqRtukS8920bDp7IxxNAyFxkNqM6DCrGnzcHkWN6a+sO3f
LG+rxNJ9OFqwHktYfAItU64kCJsD37d+iKZRnW/cXuCc4YO8gfUP/RctuX58wHbK
ZXkL9AVCOOadD/husc9glt0HIWJboBsLHyM05205+/Brpga/CcQc+gpLuNQs7+NM
KDvyV99ROjpja6Z3ZuCELtfCpSfUNtYSfsNvUKgNIuV/ndfPfhbQllQXM2vnneLl
2vAtvazYWimtiTA4/fZDRse/j/L6dCTxQ7tdh+tWveu8gzLG9AzdkiEJolL/8Kii
FJ2zJXgS3ucbGymMLK86TV0QbzXPehrcOusD1sih+dAdBurGjQn0favhNYr3fZw+
rZ+Flyp9qQ26S9h+3SPtXx4TNZcxFU1Coy93nidMXhjNCIpKuGPo19SJuP4m/G+4
dL6axaMJicUda84Cedzyod42roJGpm9rqa/bySpSeDZU0z8fLekU61EYCnWhVyHi
xI4U6gd9FjXkNYuEFXg50sY5056lPvSs9OCO5dmw9E3Jsj1Ddn+5jArZ3zYe4Tz4
24qalcFinRHG/BUfAvVCivLIe5E3Rqrdysai+0S9P4OrUeH7QC2coaQ7v4fE+UkL
3lLQkVjnaojjTXJnHXOisIgDSrl+HTVS3fIljqs1as/bBwncztwPfg7/czE4yZKw
TH4MxinpxFsC2yEOYKvJO7osjK+DETamxUtk8i73VuqHxs7c8H6TRpX+Se1Wg5OO
79s+wJNNPCXOVW1cN4tSAGYKKXOvNyboX6tTV6FxGeyoy2EHVuGvNDF8/2mST9c1
ietZsmIxs6GJsAon3VcDpx1X8whZSA8lj4L7Sw+QZcSFsy0ipWCAuHD0EdFp7wka
YaUH9tiHgp2kgHFesuzuaIgLSgpwQ2cWhBPu05GXBULwpPxbPEhl+44N0TWzgeb7
uGYcCR1BYxRFgOxIv+uS75TQh+jQxf/A5vA3K4vHg9jcIskB7m2X5GMCwJCyv85W
/dzeqXxjvagaLeP94/bdWFF9GvJgXoIRUvpiHATG7UmzhyVOwAV8ktmZPkkVwTF7
VaKcKplYy8WHXut14+JXJJX/oOdHzjPQRch9f4hpdk91Hl8F7uqDT/XThS8FmJLV
qdGfqPgQ9GPm9iDmCZIHUZeArqT4JOMvLYaCLqEe+R+q6tCQ7w+IjXgXUxd9BJLf
pJuz53S3qSTqWfqjVvFmCCCj1eum65wb+VoXkRezybQ3Sooq/boDna4yn7jSp6zL
6uKcRByBJOIt++I31OHaWdFvMpAI4I/EE7l2UUgVrk0=
`protect END_PROTECTED
