`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tVHg2S1xMMid9N9JMqvLFE7x+s/vlVFvFC44FoVzRZmO1PpNbH+na+sJdq0QZPEa
DNC8P2XqNo4K+cnvE3B7Ld7PkGak45+4HewIPwZLJVw8RayFqlNMACUOrnyEpvJy
/4gf8KRDRFGlKxfVu9ia2Rf8txNqvBYucl8b/vk98oa8zQqIx8SMGL+KPaEYCeOG
14dis23pYSZnP3NFLtkEik0O7CMjrDzQi1BLwf4B585rhcbnWq5XV3gwP4B8gsqP
2+yQj2rfxU92EA/HEOH8ORIM2EM9FM4DS1S+Lz9dsV9L7OJMmV0MwtGgZzSumq0J
oydruNLhr4K+ZIJQIefelF7D5OjZYuAWqUWfOjbjCHLO4/30UbUzd/Jcuux2xkOG
MAr4wR+yifL/QgZxrifSVYnmH6uI+fkRVE5jozhl3YwlFj2Eji/wye4rNbWnwG6a
i/R7iJUIu8mVRCFdpLtSvFzDHRpi78gTJCttwqqtvlJyZai7dG0MavYvcIkmDKYw
CGbRsMhFrJypeln/ijaOSjiCVWKhdsQAgnnRPik3rFa5/V8XCugDev6cM24fIZjN
sO2rLdXs18I2Dr6crlAP1m/j9RXB6gU2Ko4hWSvXH+O/c+j8T2AeX/ZiNHxVmsDi
lqdGwUbKHDRdwWJDU8BDBPPTdvFVY7PxA1AjlgA5jlJbXMfa1HtbzZUrsRsmT3B5
0sdcXxkwlT+5mosck/TZiIe8yXKwH/oLveCVQuEujq2ovZNehDoeB1gi8aHZFm8f
poaVmP1cLU8ilhmH+yE598t3+ceAhz6iedT+BCM+X0hzoiK8Io5CBvUDMwDad0ta
552ClOOkIb8sfAe4OMqgQ4hPDn02oRYviKZCq6lhlSrlMQQXdKX70/TVTBaa27ve
Ju01jLCnUx1cONek8nRjhhDJQ8z5XpCi6LZ2j0fy1Gw96RQrh6Jgw2tJ9/6739NT
kld9NmLhx0mhyKuhvhqdCCHC8CvnGtUskqBCJniARukYSiZ1f0hXqLo5e1jqoOXe
`protect END_PROTECTED
