`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mD0LuZT/Ao9aIcpgamVIOQnYsUuOTnQ1SS2h56h4BCWHvp4gXiH6/9M2gMRn72y+
Z7ahR3QbsPG1sHBdA91wtSflF17s1kzGriC0sgcjt/wCuvyLdY1doZacBuj8SOdI
roa4GpMq5zv6GziWiDpwnTq5OqRd1JibtfSjy73qz+cHWB1Bic6qet1RrMaNQTbS
nU2XG7B1bqWU6AqZG/WR6kGvEHvihNvVOp7Go/hiIH5nbKVfXQ4K6FVqDLIWQwTH
EKfx1zke8g51fkvCAb32srGLTu+QK0WHIC7c/6g9TWGBMj7K7ZwR7ouLur0jkKtf
k8F2rd/Yc2wukF4O47T11oC4EzClDUt/EOMpCAHQ4FVXxEOw6EY5ktl1OiX7rovb
QyJJvF32vjWKF4uZIAnvzwhovnafVNIdUugP7GGKubglFvIOQj1ah4i02huhN+ho
aJFanarxWCDgjPyejnJbUAA5yj3ERlcJrq3Z2leIUxBPGYdLrryIVX1RFbJZ+bvW
t+WNQ1l18heEAXXj2w696rzjdbFfDfjQirDj/T1Z5oIT7ymn6hin1cotvsoB07NG
643H7kRXxBY19VBp0wuo/axFUYqLEK+eZRwF2Zn2RtB4Ln+Nh9BdEEHqCDpDpkku
Yt1oIJEijVXTcfXtMn2zN959xFYMdUgzF7U8bSNhMlVFyfrXyyDCcqEA07l4hmwe
Nyt1KMmcCLanbYzDEdWhiVDzC9GSd2bM3FOnagX1taduxY35LQiY9ClX0EJ9bgoY
arf+VnpY8QwY1R7XKaYypKaCrU094YqNsC5W6uPFhNsC6UZ69VgAanAEmkuF1h8o
JYFuS020Ynwz2r/6G/L6zVYQjqrRk4iOydgK7PPxKJ2LWegDw5Je0ig6dyAH/PWu
ff1AwgX5LY0jsB1GOOxuFWM52HwyXpQeXqExIIdQg8iKhcSY4Z/p7108NqpYCk7a
EC7gyWijlkmoVB44KUAY3tJCBuzdY4lVjYjsAgxClAxfTEfWSmF8xanb4PHm2xcn
9gULNr/bUNIOMKS6RoiOeeBlKzKrGOIyazrunixTTULLZSfOPrTNQKhjGf65vGMT
9Vtp1ZBOpH1mA/eGGp4xpa0MFIlrPi2FmzjbZ0ZEB51TE+nnVYxH0E2p9g5DJ8s7
vXugzVjzZMiBJponFkdHBqZo6K53lnUNq0nPP6mO64XF+6++cev2a/OfGbno/nRd
6BL5tPb7WYIDqOrdSCZ+pzSAi9sNGvBGCDwD1VcjXFlIg4jY9XQz8cPbXmenlOvA
rFermC6rW5t6PwjxvjPpTve1SA78h/7JY2Msk9vSj/X9+MQJeI3l0AIqMEwVFzVL
NqWqCpHFi+AEcI/EcEegnNdJW3hs/h0faWCsQ9vt0kwMxqFxXdyjpByD1zyVY6+k
0LNr5nXOqYDrR4MugrohOi7xgr7NBsT7IDll3fUGfjJWVQWdFq/0wjK0kgNmMlSs
7bPB1cPbT4AuKmhn7Nl3aNt/V2bcKmH6NGfcb+SHcakTm2/HwEnC5R6a0Fu5oZVt
RejRK2ZwtKI9eb8HNBzTXqEx7e2Vfe0s19u9BXHVc/ORXC7BmUiKtiIoOBMfNlmO
jd5NALXJ5bgQ8OkhUHoBYnBgrj3WJZ0IIhs22f9TnB5POmyvxxIQGcne4F5l0qQq
DTmOHN5ldKylHIw3aRJBV9r1q5ObulhgLGX8ie6pVkEai3YBZ836gSz711LshvsO
jK0YsNt2M1m9DsEjkvmIBuj1jvtzqEfzVlLjZe4XupRVbTkgPG5Vr2yruKM7XfgH
TPRLAFx+n5vsWU4jw48jiFfw/8Oa07IqvaNa/U9D6JzCpKJ9+p/OR+4ZFDnK/su2
6td/O9hZXYRqeev6EdHs3Q==
`protect END_PROTECTED
