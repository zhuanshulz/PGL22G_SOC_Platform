`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hb1H4Zw8uU3PXbkLQrGleCDLW9DRcofKWeB6d+6bmGXmqcClzUeI9UjmO4TkGkAC
OH+R9np4vmwabyMyDClc/wLOIEGYUKHNlGrreEwcmd+rfEDwVcrNuh2LpXqa1ivD
QsNlnL3Z4Yn36Ngus4T/6/OhI9GDx2+c4lDth1emEATGqfjjNAy4B8m7tHCrvrsv
ws7gxGMa3S7RWd2CMIM54Vog421WBVShVjTDoKIT5XvPbp40aBJFvZ6HDfqI1RkO
YkQhz+Kjc+CXGsMGrz1OmW1FOMyrLA5S2dkWESJrfrcw4g6Abu1xvIQ5qY0GySvb
2QB7Q0mss7QRdt/0b4y0vt9XoN5Rr6BrhG0W7HyJNPJT4L73jc4pw4xz3SQRC+Oh
BYDk7IzTFMl5SefemFvQOdAC8pEdqOyNj3TfrzuOUguaXBI7PtOH8sFFCXFrzcsM
8OjhMQlRESXwrQWsgdgGyJGX9M/rVv2QGNG28pJ8csHkHWsahVCTfPF3xRFYX0tj
bMjnz8w5UT8Kdb53SO+RIE88GfSvHJdMVXoWvTq5xtGc3Hc2qinB09MZTqNVqJS+
xnGdxeJAinVQ6T8Gi4pVkJjJZYMlARUC7/6RyFH8g2wS5VjVidK0WvsduFOfUZgt
9vxV6B1QBy5EZFYP+krM0Yvn3dMMB8TeKowJUU4rAgx2yv5h+D0/XDvro0oWF0U3
742CSKhU4SKrZtNI4lt0bGCYXimU5oCMCWq2Lbh0N5J2ypQSOlhN/uj+wg3mn+9P
nm+OH2rAqMYexKYDXdyW+6OoAtcW8TdZ00BDSzqavZhRp9v0AFoCPX7AXvHFsX7B
nLPAmjZDQpUyTwONkY4x5QXilQGQpx+O7ap8yiH8uMEYQ+Zz2Z3lbLZA+MaFGuNG
iYEVKG+WsCLMwD3PH1yaEXo/+ZOSz/mbiSc134d36CO2FHatiowz0P3IIN/PwWmt
2Pm3XqCHBb+OUWDt1zqQAKU0MRq6k2WNivLTdVUkpOZ6HI2M+fmUT9kiYaYm/1wf
pVak92SLhU43sFdnihJDsv30D/LUDZCTQLWZLEHfi1r+whTBZf7aZ3P8tAWzyQIA
6dTqwUzfPyEhcMOfzYcm22z8alTnfT/6GwROHuuaUhZjVTK5uKuFgsq8bToeKpAN
cpJwWb4VkFzbpXAPQMYGTSuuLUTJvtlbCV8muAL7XLOwh21MP5Smu5crACWElTRO
MQgOHpvsruZDTIn8f89NXHNOCNRbww+V5pfud/+ITuSDPi9go4/QLDt0OLVXMI9P
n6NZwmGQK8VahTkgdbCCaRdMwtVCqJNiNTI1fCLLJSDXGYs/u7eGtqRH1j6Y5ATB
2UkVg10MESRPrjY2axMAc5IDmhErT3l5i1C7wYEVm4AgRcY/g2Qlen6UcYFvDLHt
ZDy6K/U3F90cosRP05jGlTG6xP6XeM74damfNJXYqnSuk31u19R/pFvDPEZ4ymHx
X/unst/lMqw0R5pN7Ap0NVH5waDUyKtaISi0jzab23QAojcrbDNNVTv7E5C+0f/f
pus0l0Sj5w5144KpM88+fIjMrwDgAO3WU+3JLSBSoAEd99ChlVlzvrmq0MQFpo7e
dnbZuIUx6nyj5SAk1MRXh/Qky8KeJgnvWOWi1gEoxRWIIDdfznkOcFGLbIdo5jHe
x3lPafjdzJuNQ8G1GEl7zP0PLs+Dw5moqbIFgLePPu9lsXkSmJS+7Rg6TJHCKfgm
XnsakeO7Fj6fGBJh/J6aBPF+7062bhB2YFtArUu+hI9DtWjGPKi/+/g0eu+PBIPM
2b+FfkpFWcuFDmhQAe4S55SOJ7J1dd7+fa+R7ofnCnozlQOW42G+cFUr4ZCSF13b
zfBW5zBLyBmj7kWGk5lh2yJuLBLoenwf5gtOVOpl7Z8FjhDmNCQEJt6WlQN1+YsZ
zs7bxVsYlfRVSy7uG2djelxX2Yge8sNd7e5DcMHipoGaOz/HJQdxWuL/ef8OtltC
MsP39kgFEbFv3aN5+w6aQHeKBjn9e2EtmGr+p57GnOBljpc5B9Sa0bK5QC93FeNf
5ealuxeTCg+xyZhEfoOT+ClIYvGtQ9/jJRuwvZ96xS7uo/1lTDu35mlsX5TCxuaS
93f1BiEY4A4z2zrr2bGiJmCTB8HFuG/1CyJTVAIH69CPPtKHDuY8VfIWjq7ixWn4
3tKvhYvp33HHtVOcTUUoxI6vTeP+O4LluCdDHfXT0wduvEP+xy8qxeG6to5zjSda
BSWm55fXD407PF+r6aN9eejwlD2bQPXobNTpmL52e5+U1mRWMMT5TomHvsJ2AoRS
hqGhC+vvczwFAqhQjEtHmU+FKGIlnBMh4wqkVzzZ32HnVWhr85RhYiE+8Ejna8Z2
c9Fy9qr+IilZ3XEyFrzp9ZlrveuwEJ7eUT1AbGAm6zdPhkaSjAyTtRw2PvBbs2hM
JLaZNWyoQ76lIKkAN5UBdjbChuONaeKGOij+dpU6PfLNd7yImjSkGxwsOfQ1W/4B
QUtsWuYelSVf13Z9E26VI5MZfr/ImKfuGnUDZjzU+0RQ4icNwKYi67xMvAbqKCEe
1Lnfsx9sA+BuwlcGJKgTyxY16JOl7qB33KghPXq/1rgvIfSoipT2cFrqZ56OD58O
rFdRGSjWAnDXSAry3/Pk3EL48UzWI/zwWTQg3MzH+AOT9kxbiFzOVPF7LI4srH94
4zLz1XW+jhdLs+kc6PuaCdfr3AEH1upHlOJ9M1n9oiSp9ifRoHPnYCnOw0GP4lID
g5RPYh6O4+RKBp/p5etJ8MIBe9KfeGDqQBFtUqVIPmQ5lEXeRYRIX86l4KLDBoUF
J4LJLD0tzIl86VZsB72taVjior7Hww55vH4GyefyX69zKhmoKEKr6jULCYSc4/oR
eCq/IW631KZFicDIyitb7ASYC+s1iiIE280URp2XIMDCE7Z/xWlMZNWX0beaOoQM
Hi6zkuXrYg1yIMhKROjkpmQCRCxU8ifV3bh/ZeJUsBY61kLVN6PPG2PUTrLXsisF
7hZaSvwETx/n6m5Yu1AaAoa7rk6b0MRp0uxwTi29jE1smV9yT9OcsT5zDkW1Krtv
IlLug4vPO+iLhZadchs4zByvc1ZwmkNlDmDG4DqxNXcqqQODbP48BjmhSbN6erQt
DJvc7YBHWaYaEx/zKA6HLdAS4eKJEaZ4VhzduqkRW6E8hTo+0K5toFJOrGFZRPFJ
qdLDZwHJZWfaVpyjhMw8gCzNFo1tNh6ciOi8rREuE7i5G0g4tiWbo+em0sFUbGE/
MWPFrmb1BBi986eVxMzgxg==
`protect END_PROTECTED
