`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IV2sXdqUPGvKc7nvwnAJej0m6VdHES2BlJdUZoXEJysrb8kYu2NiplDZTkg2hsFS
o7WwPRuc8uSEg+ZaIHpsWsVWxSbJZLNWAGJJSmVx+Zy4t0MO2+yWpAvRQ8Td5YHi
aIUqHvVMyelTE1p82ksXSNEy/dIgjnDOsNV3laZ5cRjszCN/yvGTiQEp53Q6Z3ih
PO1N5HeYE/nyamq0BXe7nsgw52s8UAt9erOTdKGSloRdSKXeGaMKHZF5A8U8pXNG
C+H8C+5LktV8/rfFeu1vF6CY8R+q+cGs155BOe2A+Xcy9hLGzrYhFXF1ifyKn0Ow
TyhGMbN7AY+KP8S1BYA6r2rWGSt6RhYRx6ZrnG3EqzJdl63a3JOnP8lHte7IvF8Y
lrm0oHfFSstMevleQGy7sdxVaD+Px3oxSeTJBwgqfZXv3fImgye1jKH/5jOC+jKM
B21ZYbKLXmUl+eXOUCGEBEX57Pmy9JxFZeMn26OOCTLALzkpHPd2aJBNtTOlKZB7
axHHvMEbQ1vKTEcQiN2V3BmXWNYVlxYQENyauFLmoQYTWxmcpzJCm1dK2R5BtD4W
VvlL7dt5LF6GscJ3zJzo6+PtDA96LpgUXdK5ERJniMsguymVuwx+lQamhdA+1k9q
L4HflRaUwc4rD6621GnVb5PwVy7vj3RQqOM9gHs0ERzVxSgAAERlU5Hr506UOrSq
oOWQfMa8r39uCrakFeJMPhD6XJRpvbSNyb10aWgcbzSU8Vgv3CbVpIVxtB1Udt6x
`protect END_PROTECTED
