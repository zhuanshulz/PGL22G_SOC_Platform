`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B368lBSm25XndKuyWb52uVTMn7U4NVGpg8kgG5OnZbosIjZimJiv4ZKqnNiDR2M2
ObIdvJ06fjd3vuGKCcAo4nfot8A9cZS2F7CK9GBbeYHVAaIB+iiM1yavJnh1U6pl
VkiwfSc0bed8b9VhR5OBFiJ46VOfa55PxndF6ZLaHATjZ0bxAtEO9A3Seass2ITR
Mol8U6iHrdTBaWxgTdUW1bgkmwp2N4FVEvzvgmg1XfzKvKyBNZ0WT7jTavpLx42n
wqTt9y9MhaQx4xhWqnED63uU4c0wj14imQgZtZaoWlZIEKo1eLzCyEKX5qiIX1R/
qM7esomsMs3Y05R6JlPgpHMLTiwNlZcrmxwx50v2Dm11DD7iH1Rjqgx78S6gVW3G
is1y64BbEydZpdE2bF+IFvdtE7FBkW3M+IIYGhHmaJXq07udhhXJxsEi4TjwtRrQ
0SdgudZeFZOof/UwmfcLj3MgRyb7mMcPkLmfYNz+W3rVmhYr9kVpoGrpeebEIrVN
FHfSCUwNG0GTuYEZGjiZaWcfRNXlAKyNmZrAJmpueRMZcXGj6ORU6Ivt46o5n+9J
C/X8B3C4SUVigcFxc/v8w7+4fbapbxaWeLzwyVgcyMrEWTXjEuNwkzqXCWeNSJjJ
8VsMThxhoIbVtrEfBRB45xq9qTPgUQr7tk1BLAtdFRpnWoFnLNE9b/3m9dly0KO1
WWiGxAyAwzpp35VLhlo0SplieHhml6NpVCPpY9KW2+mt0VVaFV5MpN0I+qH6hqxD
SRSwpZjwHOnKr7OepxmZhFBaJRNoO5B5hAH1h8yYQIgI8LunOAkvvbCT+y49pJyy
cIkvhUlsMcB0oRUROkRz4CbmJ8n4PilI3LAQ4OlMpTFcKxi0UDJQt7ZzDJ8QsTyA
5sETYgVqLMeUhoOaaFrKLjsOkVvrhDkwFUA7oEPYk/H+E5NxBlj15mAX/Oiha5i3
PuWQN01qAhI4vQOZRrKtuTGWrt+6Fgj+mJb6DOynavnn+kni0U3CjQ/fxRxW/ZkE
xT/VqCrD3xu2VxSnSuWfPencn/lDs5xl+N/jrq1oDJTUTM938jwdDjBWQ942iVUZ
Ka3f8KppPgYfGQc2BCK1OPpJ/8KkIDSOO6HUoctO3qUkUMxG/fnIEE75U/Ud7fPA
BJn8rcYMe3E2tDB3w20I/Q==
`protect END_PROTECTED
