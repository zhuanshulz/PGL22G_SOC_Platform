`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yt+u7jgXRmGtN3KCe1beo8kB8nvZMqwzWB3KSoMHWMA77dKPbpS4obUACq7LFrJR
2VYxB06fQ+1vASSjJVqwSRDn5k6lXFUpVhrHrIrHOIPm50KMEp7nTx5ylC9YPzCJ
TJKaMrX1ihYtplDgRBycNk8l3oUJYzADDVf7FLZ7HOouuXOc+c1z6FPcP+N+HiEA
IueW4gQiC0zndo1lbWyxvFGLoLsvE15sbaj5YGRAxZh26HZ6nFSEa9V/s9m4wUMN
HycUjl8aNhJC0Rt2LiqywBT3PlT/8F6U0S0BxoP5UEzqm9t1FQaF0z1GiSyzK6s2
jb2hykNJ0oDNXZzPD7NyrLKtT9djzmaith1mm0fVgPGQ4PojewqmnWJStOijX2vH
e3xroQtqc6xNYj5ikG8ayIjNpj+bvBdtrHnSK7jAMYX+sQBXQGIbbahHdVpL+tio
EZvKUccn/JAtbzlbvW2EbWdEX9c43AFVUe5qstzbY+cO9V5XswCNTnz5BprbtBMq
1tH1Yr5IlBaylBHfyQvjnxekHutH1nZEbwjTroGo5UsfafgX6ORdyAWlgfCbX42G
NZehqyRMlpK1rS4RPoDj3uXfo8U2asFo6U+TevnT8lkushBD1XH3yMXZ1pzrUpVN
ho5PC5Bf/BtyInyXWWF0pXn4yUZWwGq+ilqDIoMr4jg2BYlOc6I3v5Jv1HA4LgNS
W9cYaQVUpjZzsferr0zej2cEfX2/9eQfz1+emcDQK7o+KYMDHCVDIgQHwWuY7wpC
Rc8/ZGdf8YoZxEGywn5qVz1yNLlx7NZZO9zR9ol0REKpTQX9IXqgnXcEa5trTe0e
DCBPO+Bh00+gDab/9nFoce7Gbe2+Dz8NufYqRsp98zwzP8nduTkwgob/WCWcnVZt
Z6kenoLreSZIGN7SdOhIrbiDaOau4ART1V4irT09n2Ta9pKC1rlSxujbK0gXNI3o
Xj+xA11TvQyo0YyOLEmEi3RofAPCNqSUDACVxFIEHhNMq9bKkWnxfXVNFgpgqIy4
gLElbo7eOlC3ajVkfT1VwjDwq+OTm7DTdsHKtwY60pfg5CSYhU015PqJMlyz5Tze
/gDkBAM7ajwV8mIu2tM5Kjr8qVEew0K2Ii6IAdaH83PdSojfUPOzJ88rHrrzKB2t
JgATSKEB1m96Jf+iG6FAswCSW53tlMRLgkS3DZA41t+J9yFDRa28jMEsbXJPD1ap
tA3+VqliIRbws1/adtgN4jmeP5bzaJpi6vIy5rTV6Ymh6yT/evjGb7jKp1qxHoUd
rcpbek2fSGDhW59Bvv8CNKJLhPVAkaJ07zYoVvBfADsxWDqIkU39G7YgMPtxBkOg
626ZDVIoztbjE70BYf0pmpDNJk/OcCWi64As80V0/JktdlVTwk2F68QKeaeTPeqX
Q0R4gmliBp+WbBfLPK6Fpp8ASR1cKuJQT9vhSgfb9e+bSh7HEGL2tnFaVeewrz+6
CMwMhdDkocqlnHzQ4BMR0kBUvTWiu5SVIjE68YPq387pP73Ee8AND9RNIxrO50Tt
K7MmoBONaM39qFjLl6MLMAuq3tT26DLYR/BeE81+T1Ll5WCuZuBuVD9jp5GDPcgr
N5h3MZ9tbe4ZvonmrsUCafnsBCpvQt8ghe9AF+NtMvGXwWLu0d3zzSgil9r9Evr9
ink4zLmZ5hksxVbou2X27YCwFHQg4mt/YxTZZU2mDp3XNbmt2Cwmp6jIC+FWDfuV
uQvekRJpDMG2JPah5hmOYNLbeEpkN2/pXjeHOYX3vFQ79KXvggxfZRoU1mE8MMh7
+H4q86cN9bW4uggWUSJo5pDDLhupep4Ae0Dbgd5M4gNYVqwSYoD8LSYs5EibZXMu
YYUpg+1UB4fJ5UHL7L0JDX+CJKfwfxPfqREC12hVPOz9F7cAxXO49uRYrkNMSCNV
BL1MZkSL4SnB/fLyp81FNa0Jj0q+osAROFxTVcNWzNreusOMqinybqqg4M/sNXUC
4Q6G7HEFwn66QybCPDoSyTiuub1nA5PFKzeIRWrO2R+GQhTz1z36sk8dGzVlhadY
iX4Y5atNUUoynTowmyhM2OF5faxNTf++vbXDUbVqwgIMT9vXY+aeEMwO7DnwqQHo
mDyksrdwCYhWT54mtBucpK+/rWM6bpxN2Q9Srkrf+mc8OoHZLLZcrw4IG3Sevlb5
rDLm1RzHXgKsENkDJKFMhiToziNMF7qA+8rSgHL6gdODfRKHXZEljSOXF3IXkxXA
gRvuRC0xlODM6dg0MPc4/WUVX+mYjMTZ5/YGpdvMA8ZcaIFRtOtUg57ecUP/gMy4
z4C8fQRjJv0vepQKpMP9i6GWtxavIWDv718++FctJa0ghT7L39mJQ2ehQq4tc0S0
qUJCSpJH6F/gFltY0fA5RwLqLbk7QSH3GPm+RJVUhu17fJkLB0Q1nYGSK4kPVpdn
pUTjoKs1TXT1kx4qmpLomQbRJiFLLvuekL7scIaukBjmnhMkYCF5ujeLDuSDJtXt
bMQwnnmaAjCLPK18U1iqmIXt+HBvFzmlRPOxYMUEw45Kh0qJNcKZwQ4gVjEsEIuM
7OEgY3sh/XZkyU/2ZUmaN+fxC3NDZgTnwG7+PP3BvnXa0W+Dwtgkcg+0ytbDhk4e
JzqIhoEajvxGfksxDy276xgqkV0GtNUkvvxqNbSPaoUwFDDCyzHklKpbXuuU68xq
daoze0MRthEGtkf0Jd7EVgKeT1iSevimg4GAHoDoj9AQJIc78Mju/hpriwbPD1XT
1Jg7/3kzHGPwEqHtvaGm8UUng3+2REUaRQqdvt2uLjc6W0LGilSVJUCWd/2xSpOV
0wk1LZJae20o7Uv/w5ELiOOXqjUeshlqbX0SRcasvaJd82i/GEVE4NVzhHVPy0vG
TtjZvoe4L2i2nsuEo1HLZM2x5b0nrRvPlursAXwPI6ld7LT6KjXlu5sJLLcf+2Eg
W1DWkOWnKefI30NDHn15QuKCwLqvbUYV9djOCLDOtH/XIeqv9eXKypb3ybdXCuvx
kfa/s8Mtf1qp8ZDNUcgLy8QXdyoXYazzjVE7fW4+sWFRgZdpKqP2Rs9vwdcFlJFh
EsxocdkF1Y49D1yZHdAtOxhk+76ej1WkEoqqLbMsxbJ9xKR5zh3obsXC70dQakkp
+0f1f+tiIX61u3eBP3Dy5o95ppHsgJQDEY0fymCM6SwYJmvY3b8cpg5ntlK/iZy/
zioERqu07BW+wYAUNQyKlKlmivmZHnIpTll7Kg/9GPI/Zcz2g1xTlRP3VGNeHhuI
1T+T7sc1X0kyUGp+C/USOHQ8Co9yW6p5joSC6xpzrSGG63SMHv7lCEUxa1THlISW
t6kAx3lV21L0bOr/E6JvPDdJZ58gex+6Ux6+m2bW9eOL2lvPmDwZD/5xXadEPrun
vR4JPUlae45sOKa/SAy5V4E9yE7Q172efVYBARadVY5R3elVtnL3hdYry2xwOdqf
UWk0vWRAnTcTza6nRGFX3K94qIped1bs5EluvowprlYxj8Lz41zyFgAAEqiNIMQ5
8Ep6YLMNZt1WZTT6SeVfpwqtygi++hO1IKo5LDBTB2wH914Ay1YeR4WnrQUQlZaY
StX1wn8lyBp7JkmdYAdni0BK2eKS5Vs1NTGgAIfaFiVvBsq4h3Mz2c/GBJL8w2+Z
THWYSiUrSFw0zMU4fqsWv8+Plx8pwRhnfrYSJBBRUdNI2B2wZLZs1N9URCOxArJ9
509WBO640UtZaVAxgsOAi9LWHNYGX6ml0ckCxFj46F0Xve1jc+pQ6v7eJ7Sbs+DV
on52zeoUnKfqmF7F1Ostgt0Zbld+Dt6D1f9zTzowYQYZbiRhzy21jxj91g7Aape/
MpowQHuGCDNo14cYVz+fs4FqXaz4wESwm42pxYB4Va/edaVLqACyslaD0PzxJhfd
EK09E8hMu/8Dllt3Ez/BFZjlEBp10pBFAmg4K91AvuXgSTUimqQpj8VrzJEVjVnv
R0DptNQfCw5kczYC6bd+SmqpAqqGxt8xLO6JnII0Y63NQOv6K+S5sCx7DfrE5UmK
rg8lDAomama4J8xZPTNONzmzjeMApfdQ2GQXPV/R0BYumPCd4X1uhFUB6ndL5e02
qPHYnwNjRMrMkiA/4O30SoJNLEEwipU+qVawhG15Fd0LB/YauxI5qHzARqyVWTSC
joHomU6cZDsspZupDlDUUKc2I8onuN3AGMX+yP9++iAubB6iiLnRF8QD4pfJp2ux
YnQxpvvQ168niS91ifxHTFuvEVInt/gEB5bxcc6hoG3eU9t5Dyw8oJRbi05lQCaS
RpblkqSBDqcVmBgDK7NihqnPTskfIsSn9QsMNzw3Ae8PM4UJeuXR8T5Iaq8Yn3JK
5BdD2i8tg4+WX9TzdZUIY+94CBgnQffSMjK922oJWbSNsUUDzmhS77Lm/Bd+387H
W5yHsHZmxyaAMAxC67JPFlO+sAQUFXm7kZo9hi9AFR80IkJ8m2vKHcB/lgw9dYhl
ewkmizSbgrLadNsscgmXAaQULnvYrh6pk0YfCSltMkiqGry0pEdsg49pH4IuMRJ1
00dE13W7vBKAPDBjKLqbxZwRE0K3OVsZuFkUtbuXy8Upqp10QNALOAzHsg03DMhK
xSXb+epPC/pUoeQTDrjP+2uoId4ULPd6/bWzX9+VHsjFzee4qqxfE17sS148okX5
MCzXRgQq3tAuhQ/eYLCARtgU++IGdH6cY8f6J2m+i8Ub7Rr8efB8x3jqOzCZqXYD
7ybrM7KhT4jPrPz8T1FRSZQJ48WjsnXhtQOGukP7QMNySh9LFiAhXP1cd6438OSP
T3ePM4XRG2Dim4arzJVIZ3xxxsMlUo3w7IWGhwkSqSy1G/WQKZSdauTw+7ocHSBf
k7FZkrqq+brEXcEsX3jTRumfmJUieeorusftk2ohaf9vQcv50hpaazxH3QGcuzRW
6ZnSlM5/i+Ycwuj+yITO7OLmwYdNVQgDl6gPcr8U1fGVD/0yF8igPOoJ80e8fUco
IqRf9fQBGniXhf4+11sZZ4BOdCTIdVZBS2MorBZYtp3Uvt8AtjRF9f1xRXJtaGHt
UVBVAUJO4BOGDOLYYDmyAe9zRrkREAmx+CssLRimkjlkuKEpQ5iT4SMHr+wT8Bhj
UNcw9e0qro3uHU4PL5ON+eXONrfyz1Q3rHtl8toQnnevRsNQtfUH6MYVqBGRlH0v
JMN9HgqBFCVKpWDlEMJY+Tzj8p9s985Udhg7fp1AjRGJ+yKu89G8U0K1qhO6AqHf
q/Q8tl121FHPLiwXE4+4kPj8LM8cECB3OfwG5RNW+nfB6MwYFEay3OMCsgKqP5G8
321u+OyX20QA1rjyQKDzbV2Yi6/1rpUL4B6uSp5/Id26LwDARNSq5tIzQWt5ePiH
0wG8/E1bhKvUq6iTH09XXBOJ3nQqzS34HgXqtDAwpACA4nwT5i2yhhO/4pEeCrX/
DPyjCHQF0DzK5eNraEj3c0IgMkoR+fyocycf8IgZ6CR5dBwrKg3gzjrB9UUUwpAK
4zvF+I6OhU60TYW/GgIr7+M51veDYe5m9AH7qWQ4NA9rHjgiODizYa+OeOBA7LeY
gqwYVmVHu0suWzqg8uIbPiRCBkHCvw3fJfWaWivD+BUeGY0/oa8eDXrcrcziCZ0N
Y86xc9x/e02XTIimL+kDJzKZ9P+sUH2s2rAduwjrZlrQ/YDhCDXDw7Rcl2kEbRCL
kz9dlg5bhhoIbElD2GI8ZfLGmP9wlYmLVEbc2/oQlzvHq64qBA48UwgvBCofnHMO
dDKSVRcN2eSMWHb1bYwv8Gmpv97Gj1z9HwedlesnY4fD5a4xTYjA5ogU4d5aCrcG
BYL1+DFnbK9MtKsJGxE3hrq168lUi9ulH86SZo6NfVQ7vis5B4dtllsXoAcf3Y6b
3zwTzGGvFGCep/Mo3bHswo/tghzf7b+Hcce9Dp45+I5HD82/nkrIAqaGA2zCpdhn
GA6pkdDrtbnJVM9YAPIPOx2xHHoBYwzhPX+MEBjXiKR3+jjG/1EwbERTNzDJDQ9p
3aNmUq+vM4aLo/TO8gHE0aUdPBQWbDGBCgeZ+oTA79dw/QKkMZm4iSQrsnYjmnF8
R374/3RsMFl/jL+q3KiM3ojpcZn9giSmO0sQ2roVUVS17M7zSqzkgkvVzv/dFhps
`protect END_PROTECTED
