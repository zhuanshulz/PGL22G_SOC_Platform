`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+i+a/NuT0ll58dG32En5vqv/f/QIqtlrjZ1F2TE7tKCo61Bohjc2wB63xPh7XUW9
Wv/NIjmbmR2vxkxG5QXfqypaRddjnUScWok0FEXFIuKi8xq29aHhV+Vp00l/i8Wg
wOBur2t4wYupJTakA34IA35GQZTQfhiJbheODH7i4IOsnna4oSm0/ld9gaoQBOZd
z6APbrAzmYunThDlxXOOlndp4QMATfPa3+zoYp0NfzLhCa5+G5OwSvrJ/1thkMIY
o+iaBva59jCcf3c6U59EdECMBTKX4TbiIIGMrFmstSeH3qGMjxyuIrNlkGYXp9Ko
IVXIbIR+oLpuixom0scwR42cfYFJxuoiSJccv80ME6snznQd/zMRkIWatEHdmg6n
H45Qd8GflG+EMnOA55lngojF1zcO6+XzsIqhUR/Y7gNUFE9TqswH/wFap2O8aKpS
tbUCmPT48M91X2ycQlSRyyUDES4SL3qsomhWay3KdAu+8Ky9z+HKhJSZdxP96jgd
pHjp4m/RnxZE3lPb7kh4t5+vya9XnQi6MVS4E0cY18OyVIUx9l00CFJW6CCPNCb2
1C6EVO59j/CCARzBp55r8e9Eii0b/oYNUf8XjPENCdat91qpL73vSvKKeT+u9kli
CCRrEXNE9jfIrEF1luwjzr7U3mUaJfj6k3kYBfSs+w6qqCiDtxhgsQ5E9MyIBGN0
XEjGA1anlEUoJYEScKeY46OclU4rJf46QR63CWLMn1QBrIbOAFRJvaKYD90+TScQ
`protect END_PROTECTED
