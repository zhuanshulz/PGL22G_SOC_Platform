`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UiGYuRVsBUCOttaG5J8K3nFouGcOP5laz4QJxgD5lk8jxuNlnio7Pu4pzlBBXMEC
rT1lcB+6zf5J+CoiHyYGQ453XIuCegr7VZM//unFgXtXN2wK52lg9lUQUwagKanh
bVHIK9bqMmO5boBuD5DmXhaT7TmpBUIGUOftl95qRL307QyNSokkPTTeEktX1YzG
DNL1AfRoQWyazZLopSEkalUbs0ZYWKdZLTY/JUygteA7tMazV6zHF8XN9UHmyum+
Aq4pzkwcesbQNkmovYK+2GnURjNm2v63yqgKQgyKuoEAMpg3eEOlqSgLaPlc0kB4
3GaVVeexmyyBUl8z4IkP4qdtP29SsSg8PihBSYFrOv2kqlEdcoxrUwWsbn3T46j0
yB8d54q1IXwsibxErsLlqaohuPeGldi47XKrdV0P87DqPsEMCaQDqjeZM4SYG719
k8fs/wDQo45MjSzqiLubl6agVipAyb3OoTXa80x72P0qjqRTnbz5ExCv/wCm/K/l
D+BuZwLBYKndRw4AsvoSmA==
`protect END_PROTECTED
