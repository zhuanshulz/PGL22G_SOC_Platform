`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OZKyAlZgqFMZku+jkzHD+P6bh0rFoeiu+gTljqRVebfqZTE2zXoCStoW8SlNPuSP
HhykONss+oTk+92TwoYbTCgZTdL1PihS3NyzH6PcQozhszGYlpAJ/kPJQMm4zTAH
3SmW4MY5AlAPP5RX4wc9PN5scdLoyxAzBQgIE15XeWm1aDDtEm+kvd4kxim0krfx
hbmic1JJ6vxkP1/RLIvhi03fQFf5JUOAh0tppBcS6wFU/0V5GSDjAg3Jp4RAn1wY
qdSPCoF6RqnpRURR4gxDe5FYvFGmMfcseSvpn98oJzvcCUv0EGGXRu4wJc6hItex
x6f0piwF4HFNOcFzbcc9egH0tniOmOCgM6UTXJ9cntDiWYd3LwbsmP4DerummGHa
nZOPdhzS7VtRjYsNmzzQ9TiUUFeTTj5kb8UMRxu9Y4F7Vvwq2gwUFFGm+Bi/V5XB
cBOTfV8/mD0UJlF8L8VJB+GbmOvg43OazZXmOOYOkrNhqZkLQS4fhq6wQnqMd8tk
Ix4fLGt1pW37w4gSVNQsggHpcFmp57MPlxddvb3fJtiOv2VJkibT4aLTBVw7TGid
bSjzpWEvziZpnJxkxue2yTBUUH6o3s+y1L541At7P3jWl49tNqSTpsXD4SP4uIfC
x/rDWwtn427e4uUd745TQ6io/n0ytmH7Z/w4hCSbUIBDMW1TzzcGAgopDyVNbl2m
eMDCIQr9X4PaXqn1GfXCHVijb9UWRvK4ja//qSoHjr5lUAxakhaJ060g8kqzhtJY
MGEQLFVyMkAXp/4Mn+YgGNiepYChUfEoneW6KweFMzblaJ8ThGvlRk1JCATaoB1m
jswUxFchzyv+LJM3uWFTZ3gsPHr4wswrc8wxcumXvK8xhyqqfFiFDEyze5yWLwrm
dDNyHB9ycI8KGbapgPzNQ0UlRzg2+MTKtxs6wmPYaF8s2ZLzaHkLzxnaETf0mytb
g1DTr6kccmEFafwjs8d6gGFAwHcZa2aKUq0LlmRNd3Uoh0ateu2uqj8+f+TxnqYm
joWDsoSYkuyA/aFYl8qyPGJruuMF97bGjTA+uNsptzf6Zdqpoir6jAHXLPCj2A2u
FBxYOk8ELODv74cAhPe1rqEAs4yZ8dDjVUBLN4Wwsk8=
`protect END_PROTECTED
