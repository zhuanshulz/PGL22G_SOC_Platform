`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
InK9/zTRfOHcEPy+KZPURzcCZnKKhnAyLMNNnzXjKmAFR7zwPMCXQOtJcWXvfjkS
j1DGO949Ddq2+KTIA9pedt8ScoJGJrM74VbngS2gpNc56gCxg8yHPDtc1cdWkM8i
UOwOkVV5tYUt2rzolBrUBI1wPh195ikyMFcwkgLsFdG4I8naJ4vp1+x52F7nLqlr
n65/uQVhSCP3bLYNIejwHAlYFbOZJpvLMN9Ub5T9+xwVyq9xM4D84kdD+YtQO8sG
c65Ct7a83qf3KMRlbDnHSrJROVThVXkYkbQMxP+ltDzM+snI8EVYxLM53pLlDHra
iM4uQA/Q15dZ4wYEhMZU+H6QzQMqkl7UjEDyNS7mASljRmd6C4MMJLWHgNY1ZioK
8RwWkA4c+1LCV6cG71ujVg==
`protect END_PROTECTED
