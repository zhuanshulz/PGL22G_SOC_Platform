`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/YoO/xnQZMnkBr69mvPSEs9advLbc6K77KM7lF8sFj0cGAds8/yOotL9Lvdgy5S1
6Evtc3X0LAzRCFlB83Uw1IjaD/MbIh2KL1LaNhZqmXgpZi4U6f8giIgWuHPDCaD7
geN1PJQCd1PWpS3glXjhVDGxy35xZAp+SZo67IegPu/E4DnvPMlT9aWy4OW+9dMp
LGfYEGqypMTquowJIQ+fu0eWjMdYUz/jPu2OoAhbp7zFJwMvdmOK2vZi5Zo+MxCx
bOqHfVcz4sT9OTunPdLh5NqCYVADG5qAmahJIwQE0gAs3sJGrk7psSEFfpmNjh2x
PoG0OAyZeti6pmaZLWoJU5sOPCXEbVOFUuaIbPMm6Tv8gawasVfG4N+RnR8LNkcL
5NbYKHlq/+n2foYsOPC0Nfs6/oMX/qk2nlmM+lGflThEcJASgXZAcexzOQCY7BhX
2+EtSbECvcNccjbhlpaZqdIKKoF1vEoajbkL9QbXzpl7dlfYc63cQv54o+vN4Vyj
heDglj1BtHx4IK8XE9SIDPT1g4gV57/npVp7q8cArA1R8WeX9NXEoyDCAPvWHvGJ
OzA0A6EHRHzLu66D153rybSesfKqNTqMvTg3WuGmhmdw/R+4bITAZA2cbTxS59DW
iqiBcCjk3TFqRZaeN9O7qyrsWVzkeJ5QNdD9tpMSvnlA3seG4dKpJ/zlJKhTgHVU
epkj1wf4cf2RnczZOzEaXXftaPK2Ai9rnPYgFl6vLuWoNdxN33R1JbWE/D2toCl4
v9lgty2ad/Ot57tD5JJ/rGfUBfAFqFov3qd1IYJ1EfU9nBLLTsvMFPjHCyvKoKOF
onAaJmmQafszO7LU9+/VvANEeIJLE+UZgvW1Oql6Mzv+XylMDyh0avt0Pm1quyv9
qEM9rsUn1Du4u4cejZgfK1lNUM0GswXmmkS/jgqYugA5lO0uhbcHjpy1DGcDkgkh
R45aBVgYVQ4F+BNvvO/FOcC1a/1tLkkuFrfzOc0mVHxUAAdoYaUk/2sTEnZClCd1
intIO5hFFDoajfGErhlrg6aiqG0S/0TtNOC6kiR1V5ZxgVLROQ0EVv7unh9C1kfA
gJoczJEmRlGsafBrkP5EI9WeIypIcvBzlJtN8wHvgOIxOnNnAh3FX0/mev911FcK
Agj0OYJezFi5RiVqfaIhm2EZjI8+ihe+53gTyjIBv7XZjyQZaXoJrExOcvFt2KZn
KJpj+70QbVuu9YNY/eC2CjsvWivM4BSR2ANipDUJbmI5MvqSQNNF/zPunzbO2Fuk
HB46ovptUt5bXnd26aqzYcquHvO+mmAXqNUijTF16o3AI0YSjqpYIfDZeDDnFpnv
9uw6YqkdTiDyfcH11aZ9hAem+sVFG64bM+940yKybc91k6cCDExHHi78+nGsr8B1
Lrh0GvrrsQp3lq6YXZpMkbgwwnMdGq+d5WaRh51IOgACXTfIYrRmFv7VX3/7/wRu
MLUIBxQZcVxPIz9Ekj3X40HJM3kWfy5y+uBTSWu7nEJgCg6mYNjNJi/zTXCes/bo
Nxsh/iuxjAQFe5FHwR2kN5c/HoNvnIHR2vqOnk05YWWoQQx4WVS9ZZlfU+KDkJQB
gXXvVj+dMIGzd08kLgkxJWhfHfXwBj0X1PPmEbXTnUSHsJMaG2JMCr57r276iJtg
A22RGRZpF/jI8F5FAYiFnZW7bdfO7WcNNH8FUjLl6qQENgoktQMMKu75EFxSYoZU
xFbuexII2qIdn2nhzGNJbwYGJbNOLzGb4Agn7bFInB+uGO9GiRINQypTDtLCRzwV
I7va/RuQHlY2LlmMHNK+zXKVC76YpIZqsMzkhdFh/YKKBNOMvBDddu9ujIlfJLXR
JFiplpyrcwLjH3J4ZFDpzMCE3J/zRaMO6HJUoPCcGePvxGe7ifvzobus5m7TKLlE
ABWPaEQsblSIJ/jW1h12/jAwKTwip0saWlVZMvexp8OGJLF+664zxJ4Xv6X1N2kM
f676fZlvnSPBaMHZEeUXQjP8clXpplsymCmbPvkviXVF9gsd1iesnt0DLE/UhsC3
JsFaIrB76yqFe+Ob42tb69aZ4FR5B2tVQalh1byUBMX9sLFXLzbqsUst7a4ws2oh
WfF7DEX+ktuILxMbQxUIaYCwqbVYWibmZlBuSxBeZ9UQPdKY4l+WJcR4TD3gLEQZ
i42Qd0HA7q/j1oNjdtUt0feJPScFNt/6Z72YjTjx6/GHq2zd5Y2Uwr5wPik/ewL3
ae7O3Bwu58+yN75UaVSDWWjqWoj6PR4u1XoKfv131hXEn4kXuUMZYRD+onQaFHG9
DHNibvN1Rh66ZHhW25cxs/BYPzxHcp3w4uNGU720wFy1uyAiglINvpkDGqdDbbXh
7gDELhTd1CTX1N4ATm61hCnkw9F4fekhPc1OrI+XwpxzBgWtrMbCWlFOMsI0y9wa
NVfJaD3sbVRerCW30wi4vvCXOm/2xxZZwwJzA6L10FOJr+sQZt3Lq5d69/tEZZwM
I1uLtygVR2zMcqpGz/k3tlehrSjCXGXmQA7Zdl2mG4EHhetI+yjD4bLm6aA56Qk9
31xFgs8NBJmDAPrC3ZXHl/wUp0sMLHt0dUmyyVid3FDGp4PQiJshUmTaYPl9uRnn
s0JKgP1GqASld5kW58+hBC+mcagSI9GowHE9XjHRgGCefsmEWmBlPQcbStuMvBEq
tWCw/UJBPC38NHzT4c870hYW+D5F3+WuCBKABtPZwwGLaNHNj1CN9IXI1KImmcRY
PsKsvuH2/IJ01rUqQy0YmAMjWbtNxIWqTBkyUzrcU9tR8cd+g10sJv81u9kDd49F
Zhui6gkwievEJ494cl9DfornYe8VljcH6X6lvMhNmm6brfbpGfHEFQjNjztawoFy
Dv0q0c6wKJSol1td3XymkB9uvZSL8YKrhJWVvyfPAIxvKEuACDSnX8RRnkkjofRb
6WyY+Fc5Rq97lSG5KjZd7l+wwdIleHkNwmlboNCjr3rddKPkpkq/Lvavip9rxte5
1tMylohoeJc7RVjfGOlR/MUijPgCudvZffqfjNlIlww=
`protect END_PROTECTED
