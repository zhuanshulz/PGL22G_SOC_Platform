`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ml1BoSVr6/UZJinPCr+kbGIrF3obuigh1fReB/mQ9FEcy21qxTwa+1RlXhgtercH
JhS6O7VZbOnjKQTBWOiCM4p3UfUvBB37t9Ib4vZ7+RP0y32tttuqA14+xYn9AZBK
EROh6sMwyCTxVkdQh/JuXgQfODsb1h4mWV2t6T0/Sw1fg+kPyzn8WMOO9qHO0PO8
nF5c5EgnjggmbM91ih7zkq2mBKe9FJj9oloe3SWEJQ2lbcIRmYCQzRSTckiXF3uh
qlJF/nZmm6GQdQ9+ZeNzFR1aABtdb2r6QlzpOWC39lw=
`protect END_PROTECTED
