`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FJjTiy+aQkKPKSj2VriBPHtTOd2olAWPvRgtn8sYdRW7o0gNet7iCV3j21ONDUvV
titn+qMLdnzG2iha5Pw6R5UBNe8l09eXsC2MRNzXPelx9dKnjZpyGft9lmO7AjfY
SlnsRv7k41uT6ZuexQlOXqmH/VV8bg8hBGdbkA8U2OzzhW6oDRGYt1H8u/hTo23t
DPUbruQAneDL8ARrtfgNQxVkT5f/+Xx+/Wq49ugj6pCSv/C9RGD6nO5Ckpz9qfui
IadyhgfLxt0Y6Opy/GsWAjQN5hSCqwe2xgt5k4+IGhBav+/nKIkxtoWfFn6Yntt0
/w2Qb2C7jFxAgVPI6FlEyp4FRrma6zJpondYQkHqEB0/aQSu45MzqyulT+qHdqLC
RF0ee+UVvqzEqv5rH1MfnqrGmsCAG4x0pylM06690lSVFQOsRwM12St44x1TG6r5
JmBSDegnQLW7aFQ7xNz+PPI8WhkUbIXV8jh1ISC9v1WULlUMO2hLhCHU4yNXhvwH
EIfRc8gROf/AyNwTlo1CQp+/j4jRiuDWAr4vkr/9jHPikny2oMQLqjdX8HjLJxXe
3UakTG8itJ0kCDMcv+4OWb17asQ2htfM9G297nFSCIB0+QSlhUhC9DzqxclSzXmz
lh1bLGuhaO4Q0+L4o8kT0vknQc/cdoQOWrTn66O1BJKIkRkkvpWeu9+gDFnk6xtk
hjqPe9cfVq1Xb04QdPj+DJSJvrX8nWZU2PYddwdVkEpqNAmHW+al7AJkrrrh7b7l
Ee//dEz4mIsg9asusWiUALLNtPDiLU6VfN0IHWcjSuTh9KT4xruFpt1luHZaHkzA
fVh/Ufm4a/3Kgf9x5v26i1dpDYXOFc+L2csmaL8DIiVrnKOfiyQEM1J8uFOcGXD8
shDHf+xqnqfuMwpW3/doie7EwVgVOCtDSROBdoMQDiYDu+KzY07GnVu2MAhfi/Z0
Nh/G7Z3KGye1QjrWD/2l3vC/xgIknQ/kHk7ISkjThTf+a/3sltdV6w2/L9YXxk10
vDMTcW45Q52eqP5b7IRNV4eQZOclY6r2Tri7m4UW2kqgNBm9eovwuqpgD1B2pQ0m
cAYGWd6NUZrxKpxv+E9DF6w6+Qv4YRr1socAji7kAf6pxhDZJ+1H5mPt6xy91kda
3lM+9E61TI7pfhXc3jSIn3kR460lJ/uXjq0A5fJOJjd/2C4oEt7sf5lUhJCvluAo
626HbQa9YrNgviCCvAzsCZCGKdIy7YQZOl/nGk2glVdjch6OabgQRasJEGlTj6VF
yjJaBfkYXyXiWtXQ8BwASm4a6HaiGvU4+4dMniUh3Sx/s0/z3eNWZdQoumNXNLAE
fXqKqzZKFNFq5dKHWNJhZ2N9hbJL7/qY0OLRCK2SQEXYSKsOppA9ac12GSHiDjmh
dho4XKfSNwTHRgDouUGNAXDDmP0fgMC6wWCYnM1fsrl48/2tzbjO9/DwmfCpkkqk
13arLs4/GXLrc0vIHKiJZ9cPfZQ1CkBVSBzQbEXwWO3bLBYABQBG91dmQcucVcBT
1+JStJCX/Gi05LGS6QxMYN+C3pFtIFMHUXtTWo/sWbwxTfo3RTYG18Bg0omts4W2
uZlSa/lBBdQBJNNOCfTCfeHxFJ8p+zW1x+Mw0URITyq3vC/xRC50lOZx+onlQHfl
F6/ZNz/jgbcpwDcOI706aZFFTz3qRD2CJtYi7ka76KWbnMeSSL2Sw0Q/kL20LGm8
tSssOLBxzHw8MZAG+Lf6ltC67JTFWh5at24lT5e5YeGkvhpW/GM5qYRt9Xq8zlxz
+NTsWnmkzhzqTibPw9yCFUbBxdOumlb93F9+E4p4NQXfDoMrkNC9Wf09mGH8SCEt
Gaq62ZSbjdSI/ODAhaEan1ThP8amSFPTP3krM62cBPr8IMp+0HTXg7eMbfMQYWlB
Rrs/n2n5eObbgkIUHBFDbUhqgoCjDX8QXy/2JKt5M/flSmUgfVLPk83n+1oBqWxW
BxVOXwxtKUJTv1Q4Qr0Ey5tGylQr5+zTMKaQKI7JTHQ7CkzTX1iIUrHBNrRNgumk
YYN3K1SvTwLTKkAJLq3eHoIx1zBn5pXNWnPVa4DuzQPM01TS5EuoY5mVc4q1jP6T
/61J4wJfnbPSvuZZJd3J4/y+3XFY2fbXaKgwxQoQFyg6tE4GgeRYgYdq7fu/GWna
LtDwJVBO4RKrxPA9KoM1a+3qhhaDGq84LX1TCfh7BOo0OP+L03pohIXnB8ehBy/A
eTclI7n3YK3asUGsJK5DQGx/vY4h0SXMGHwzOpU3w1cjHmC5QALlS1BDJsGk7ceV
bgY8EDyZIx907/HiCN1qA7wJG8hzOaXW7zQI6/yflWOaniE9AYdNLZtEuPpNHo/b
v93qL/KY41t6V38sPy5Z4gn8ZKBpdLVWzKt/2N09p9NptQjI2iZxf6FgKufepbUv
RRfTZo/hW2DEUl70kSZoQIVjEOer34xIdNj62znwKr9N6js+25iwsRZCoVs9B8lH
9UdrkupXaCFwGvdcMlGMaFlDYct0YkKKauSsBjG8ojkAJhtCwcL2RrFsNpCmU/th
eVyA56QkiMyDo3EyZIPakgRpY9axDXwb1eCTg8P/pb8anzPMbn+qiVueCafqyh4u
eUtK/fqsT6W5rhtpflJ4AxsQTC8B+KnRapwIiLn3Vsi7+LZgnjEpo2LioCaSEJOD
QlLJjkrStOcYeUPR9VmU7/TjSRmCtIs+VTq/OQ86qvkS/7ieqylYv/mruYM1mB2n
ij+MZCF8E2HY+2VLNhVIMTC04uICjV2vZsIhgH1E4u+6XAiDy0lp49+tNaeHBtMs
MeN2ANsVs1Hyc+elIwfBjDCvKYKIuBT/8nmcCrWe7VyWtsuO6xkrgdB8Gva4XlgB
CS7Fpc9fcri4ow/2BogUtiZu6dWsRMKlyUwmgVVraLDw3tOeKAJCI2iC+FVZoePn
V2RQGWTyq0bzxrDr392T6baMoSEkX06yLcoSBoS/k9dEXNz8TFSJMKMkoUf2ymH/
Q3UHEeNGCdxRLhrjIIiYA3SbkL1xq4z0pR1yZGlz/k5cTXplvE5AKR53c1iDeSCJ
4Cka4VwFRadp0HR0m2quOxhOHLF4wN9kd4y13IMHuiL0Dg44D+IDDHBvHX7V8opg
iO5CTz8RCPwzPQdSz6SzQ78qF9HJVE2ZqHYM/QgM18jZX+6e6hUi1JnPMnaFxcpZ
kYXO6LlBIYu3QX9CLgw/qylsPIILERH03ToNCfF67kmMnoExqx6NacBHIfut6255
VQChnQnnoT+SOJZraUhxTZDtE27LiP9c/h9jEnB+I/bg7s+1aQfisNW420LQeqaw
5HSpP8oN+nVr6f5/8qEk0M39N+NyoXmzKm6EkZKn00ZJeVN0xMQcnmeb+IHrLfJ+
/OSiNyCkgQXuTOI2rFxy6UaVPVg925auME2Og2uuztC4gASNRzo8CIhjR34RVOT/
ALfosXULXFju/1+8NYVH3EzdxIXpPA1dHSDEpLoDni0MH5apAniwJc6PhvPWKGhj
rjTyTxmlbZ0HL5/+jbhQT+SLMc2mam/8yAwoZXLyLns=
`protect END_PROTECTED
