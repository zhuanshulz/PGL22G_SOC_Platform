`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
05Xjc8Cg++VaKgvmhchoe4yJTkw9eJSVCLOtgurTnGJoiczVGUye0IGtRR0DkyXR
0N+tMlnhAZ/dt0ygeTMfgyCvVo6Eha+9YSHFW4ZCXkhTLxagDBt4wUqCA4Wn9UUl
KgTTLFmWi7UkQochbqX/pHDo1SGePp8XgmDH8HNQazm/hj+BeS2ElUpvRWbo7ZD6
va3m18gFSXT2EQxtIHcWTJHTN3qqYya8MlJ+IxScaPDBbSMzXumqE7+8qwT//cSp
0XbNtwDqspWPI7/1+OQCmzj3HvFySz+0RdNRp/KbCPp8corBGZCWo9bIsnzWnY26
WBkBy8YXhbhLqtsXDsdxbQ==
`protect END_PROTECTED
