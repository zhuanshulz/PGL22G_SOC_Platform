`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
purI+9FneORKAQ+n9MfISeizstWkQ4faxUP1D0OMOdTmmXMYnvHWosXu0oZchK3X
sU6ZYX1uH7/gaFL/9QEiy490wjqJ7g7FmPPWyqbNHDPaSorqXQPq0DdU2o69inrC
UdWUmkwwPrdIpHhOJ2fiDpEi8pmNXcQyRbLTexdxAqGfJ1YaIc5dAc6XmCdWPzva
ceEI3CnUUx0LkW1Ge/5Uw/Ta08KgGhdRGEN4qOsoit6wxG4JNHo675xy/BX6NDJw
tzRZh7LKUM28//zADCiNSEU53MpAMMswMtjbGWY7MRvAKBlaqEjkhVCjZMcW/UAC
cCyeGb2sRDDu08YjNkFHx97RvNsEeZM8rV8762/XFPxELpVKGEZtY0xFqV56oFOs
VTmrpTNCL5oSJoAthaUuXxaCBT6Mf4K5BFel8kA91QvrMS0XqBCYuEi95KsifIyD
EC10wSmxXCYV6IJ5Af6LAB5OmEalvj+W9m/TTynh+xVHtHfRcAVt07MFXoGX5VvC
+ynjy26qXhrUWyQaiTEdSpTq+T1Zqr2NtcHmdV6AZjT57ZQyxo7hYF1y8rbfTabR
PT2FxDNAVHdbBcw+GUf6NMllZmQvVYcMXv8w59O99XNLaY4+c/+YjbQlQ4huMWWx
fHWedeZjGK6BFHuMKuy7Dkun6JQgKfMuckLYveYCJD0njG68zMMfYViL1zYK9Yi/
/YexjOGeoVK47wiOMgsyaB11fIZluN3nbkKZPgrCvEEZ9OL/YCZKjWTLb7scZKxY
n7Vqkw7e4XtpyiwZfXggGsN8ayAfdUSKfhx/YTft3+/7nC9eOi2LFMTjHUX44NCq
5P5Q8YO959X0Tum9tSL3zBUAxop4V7twXSNnTZFJoRonS7sxChWkGoAZZ2geAbJh
FrHQ3II5KJHwh0VksuVYk5QE+44KwEWDWEUnMgWhP5fwStcBqI+msZ0HlOjQe6Dq
2mAisPWzdgoGB921hawN+PdqGl7U8ysc2AJZHe7/SNt45E/dzxoZAj/JkxDTzarN
8vTEJ4pEEdw+BVLEJI0V/+fUC1Pffr2ZntLYpUXvgDUAgJXY/h8eT/zAZVdiDfRA
1X01BtBYMdyaVUUh3/pSinfOGDQanS3vAhRNxfySkXvtUhL/V5AanH0e5BDfQD+k
aNUvUGBiySwVaMcpqyiJOFuVuP2DnRRhyZ6mCGN4It6NDdpOQTuqAKiicBojdOGe
zHMpQ7yw2HgA698Bv20BFRvdn/vEgkhWg1pUqWTcyNrMrdnDR4O+uob5SZDGbEkj
bahbp04XPc3heteRnUFBWqB1d7YG49DbPCZG5+rqjS54A7S+TSzcxSrReXq6hOhc
fA1JAb8RztEKJzIfEEiv7iAMycb6H/6JmJ663g0wZWr9xORKIx/1viWTgmDW/ko1
521P0QEWe977SS8P94LFwwYnC8M1poDlgp9eeCGgMoM8xBFAxogzopPWfeMHw4bU
THancazQTUwbpHi6vYTCJJP0bg3pqHyYpvC6HeMJAdXpQ17Xrg/GXz2vOQxDIBeW
RxZ8t83fH1O2rliTTyju7u+IQD5Z6Livf3NZ8BjHX1AAU5PjnMyODe53/GvZd+tK
CvW280ehaje7dulsOWcIuB9GQaDaOuoKDR5Qq5UP+KjksdLBsZMiaXnLEbwy2He9
wofjfD+R3YRb+2mWvTlxarBt0k8/ivKlKkY0EPDK0WlSCx6fYkm1FvIY5d9CMGy9
NliCHQGWm62XDDtb+rlyOsRgRXJJ3qGSP1rfCHAZL3LQ3KsifHt6Hnh8furK0tGz
mq54JkK3TBz/jXddK7Auv87DaEsm2bFmPIv6YeRWtdNW3m0ftbDOi933s1TSZ6wR
R1gTOK6+TGuk2H8wTeFDXLL6ZIjAAfp2jFUdUIaXAPGfZWTAM8eP8zU/rNZ5kueU
YMfGA7Xg9L92G3Uluh0iNG7mBUbYCUPzVvaB5fpV/zWROEw60QboSL52S8dv8ZG0
KhWQ4tp/ay/KlPe0ZDsgCPZYkzU0+s9si2OyArZKtw0Z+ZJMmmMpXmXv+BCPZ29N
HsqmDexc/bCdS+JlIcUzQwqTQY2y9lPZHU44AIxdCzjLx0/5gIwDWaCAHNL5QPI7
rTx5Q6cba9BBsuJayjMSm0JMBtTcRr/F6SeZur5RoWZCW3a17vYAjR0Cfz4+DNeZ
sLzdiXPoAHPULCEA9IQ6uMAp3kHufqD4JcXA9pOvbKPm1BhwO4DVKJxlHgBbEOCc
0uzoRxnigB6Vlscnym1QeS7nxx611GEAAIB1jxd49Nk+xDu5eOySwgeWZ5tSV1pf
gQzY6SvvIGNfxTA81s4cUUEmWnq7PNlHuQ63+r70hBSeZKBUakDe0TPzvRZpGkMX
xdRP1pyGXpuUFCA5zc7CGTY5fVtGx9GDtb0E4oQSJ4rRUK4puIw0i/w98nnR7nxn
SCaED9GxGrxwjGN761JDoOVvnJzVebVs7MGC2DhPcelhyyW1IFaRziFjAOpSHXAm
A6qq1mFBXCvYUSQ5LhEKd0H8sKrqXkfvkvZnMxL2rRRnAtUPr20NG/qmY+y90VsU
J7zWYz7Q6s2jRss8anPGRLoxCcGsyAkPwAMwRg9tenDUUNVT1L9gmXR3zWniu2Lm
nmUkXaBxbs3bpoOuNjsGHKmiShx7ag5S8U+/Bx2y6AfoQeFGexPXzDh8dfgi7JIH
GIff53q4vXZbN5KQFpROqOyGzP+xrIIwPY3+5R4b7FCmv91RtIsSsv0dbXdrrjeG
hIPML8TAf75HBSd3HvYlwaxgMwrsA2WFaq4/ox5E9AvpPd3/VwV/somd0OpE90es
E+twHizAu+lY/GQFn8XR3AW0UM2adovpH0hQ9CzWIu6gjBbkoElPUlWqhbaEM7Wx
hWShZp7/b2ppwpHc3QlVF6GiEuBUQJ6C/PU1vSQ2r30k2cnPbyK329SujVWXPtJZ
hVhxZteUpz69kDj6mYpCD11+pY1IFZ8zNB3oXSHA64cKDciRrA7gU1YnYEFzV2Ns
jV3wrGcNMzxpQK5Z57YhIrU7LcA3+YU/xEI+uw/bVGYag0yHU6zyxpoFlyTMsgJB
aqCFtdV5sT/XHF6r5Ez5NdyasLpj+h77fk6SuUUiNOg/z9j4c9C/RA9195Lomrr8
3GKLI9Zb7MDigWl87rcMnI/wAGPKv+Y/YU/ZhRYWt6YWSLJePt0tpp/DTKXtCyYl
ACeYn6BTB+F7oXKHWyH6gXEnEq3NcL9C5Xk+C57axWgboobs6mPddipCY8yhyFfs
fwDPubjrjEQr373xuiv892Ys4u8OP1k8UgxhRpbKV89fby2T8DXewCEH+kNwHsHs
0YVWVmXXvYX5whrDjvtmY4QktMUd+7JCKq4DNXBAWv0pFf5i/zGxveWWI02FRJjx
OR7/JIhsBTygMiMEsbQz/nUpJuZUHPD3TWyuxOtFNPNazZgFAar5GkWzNAb3+nLG
vHXxQGYSIgCBsqkJY18m1KA8N7gPJXP/RhVg+mHkyTxxojLJW/QDAOTO0IoZGjhO
81Ap7ca5+CCOZirvGHJdF/swrdWMccGwVmczVyV+ZAQCTHrG3lrtdGo6gVSe7LRS
pa2O4FfN16tbu9ivGTzpjZ3T4npHI/VVVKqG063/en55WU37ALTKFlv7huRGeoNu
MUMxth54LzL4142f1wOPkPkxNKXMuo3QsOetV98EjOyEEqvt+QgFyvxy9RdYB+hP
uBHXliJH+DFZIY4NQ327lwd29M2RZjajDAeNL7HQTBM0+6iiaZaH7zq3REoh66iW
AfwscSho03ueyPwKWDhP8u3OjFI5UObADQgJv847Dr4RSV1oOlFjFFeVg+jxcZrn
Hgr4Hu9ob+WKZEy12bsRabHV+pdc5jJNxeUMY/ySYMs1r08+tVT3dlPM5hswRxYI
TEJ26u0WPZu5GyNHjs0JGqtFWhVDH48Uif3/iPKl6I/aPLSq6gYEZs/2crTuf7Ve
2q84bdS9JAFgr8C3Qge/hr5g9M7tPza63efHQlGvPgZg25eU15oZg61I53sbyz2r
9sgYRG0WcCrGfI9xJzp5/CO/fq6JePiG0McJgPOA2mn+wMHHfNQGG4PnCys4Zlol
piXDhPXdO7myXqxbRM7umkwzEwAjvTDZIpD/PlXAHRJI7pTuvmegnbOkzrlcUmP7
SpKoouHOZOa6yuYK8FGqY1yTPhE1yv0OHy6aAd5EOeb4v1d7E591/mjLhCbTh38q
quAu28OO8eQGMfyPDEP3/FlneO38UkUe6jmGy5Ydpxaob6eBw4Ly2Jv0/0Ak1Koy
ObmKMuvpMJrMmEGCUSKR79bPpbqTCSj53hLQwjjsl21q0vHClCorbmJDs9r5FtFp
JnZHaBfKVo9K/l0dMQ7VT3ISz8+Wa4x0tYb0nrfZmpM661LpS33LNYqi9nJosLfn
gZn1AEpyLFaYn66ONV78M5RUwAPFiYc3JUilUG4GPu/P54WJ/uKV6NYlha8ZKifw
p0oPqJ2aDe/W5E32SBkXmhgEMsa/ZQ0YxhRbz9jya0wdIxSV5hd2AR0rfHWbIqSs
4DCaELr0Wg57MOiff3OxhCj6JVxE76uLpnbQGqEU/xMvwt4z0ObRdupqR7018mYC
JliFlA8veRR5opiCAJr/ikpKTvREfhK/8lWpZ6rByMZCZrfqEcR4E/C7PnnuSpvF
vKssDFYSuGqXUwb48kK0q8D5w/G46p7QkwLAZCknl4qNwu+VFzyIjdhpwp+OZihv
SvuJzVBfwpeBhbcI0nH+2uPbzxzIkhHYAlH9JF8bUeIW36BXzXLxEAu0C5WwaIyC
a9EK+gOLrO7+/n+hsM270ZjryCpwT78c5XNjyfUp10rZgqmBKwxxT8vTkcHNksQ2
VudIjyjX2QcPtC4Ki3K3lgWpSO6ol/FoZrDW8LYeC6D/qlr5s6hREEnVFdhT5sAk
eANHcCTOY5FDmh4j6iYbo7RfFo/FhAaPdZsNk6mOisZLUL4VmNQwv4vkZR+z1x/p
xT6hA1MXWCRpuNIpkaqA4m0mxZUA3cWru1J0c2olOn+I21C7ZDlV+0OT2j6y6Rya
j9r3EK75uMJAVSccXglDqnj196pXIz5oOoeAl8QwfpA3HFBn1IgWOVjakjv3YZSn
Oodjpfqf2nC2LrIzxgzeFpfArMpmVdUlApI/hBiymKJyz7JI3fHlha7GVuCm2zJS
0qOOkpa9vTBzS7EUVeQbSRIJaUpU0045JYqGMGGGqineMuMebNGs0amKEQ8USdBT
DPw9LmDxmN9wzh+Xer66o0K+jhvYKDl7ueU9EZGMDi5FIWqF6wgQn+KV3CLmoiur
ISYe/wlXptNuPJTRn3brgWhD5uaRnEW7C7Q3lOs9dprBiXJA2NJr/bFTJyYngigq
e7GdGDMPCEqUuJz2SQIWnGu8TG4pDKuIhDQosg2SvECfpWXfevuApOAQiWSnoGzw
o0DAjLwZtTBGrIMFMbIPk7b82W8G+spz+OOiX69l8iQQOo4s3bWoIvc1fa+s8117
ivTtgbQgN8wgoRIGLVAP47jmAlDVPzlIZLWRROwwM6Du2ofS3Chl/86J213vlLPe
C0zUA4/9vIy6vcVvXL8P2rFjgoosr73WYIT0ZE6Zbgc0F0ArXF/nLF+Gv1/P1k/9
qG5Zqp5YpDRxgVL/5uAXycXJe1helxzz7GEhLcvJx2dwrS4h1a00Jy96NAJ4sB9x
wD7+IqMK7oQZJqqEIM5leOJnN6qVEJ8CACFschyM1n8guOrLqc0WJWq8ZSizTMD2
ppFrGurRr7i8e5vDZ5z0wnNyEADdxrl7XfcLKMm8LtYmhAkshIEC4r9B/B2bnFe1
hafzfZ3Jrh5zPF4IOl7ArvBblCdKYUoi6PmC7UgTs8DNbkVzTNUnSxzqHy9vnVOa
AUyGErHw6x/o4rvRDa6R7tMzXgHncouvFGxzXMC7hSzLtgAIq7MAAmQLMewOGgJA
7VhqsU/PT4o/o9Hdn8j7GFIs+sVYDPlDx3LmAXWdufWIEks+TZlsgWgOKlwWXQ4d
tiPxWsowWily2O3F89vTW2DESTIznMsoig55E5iPYj9jHeJwc4H45bLNs9VVSi9P
Agr90biuhTkd+m4f5A7wNDw9hGn8psVSvSjiCvJ+pj7dpXxs8pIWhWO96ZNuk8jj
2UR42/9x9G/Hd0kp7Bm5D3qaja1TupwivG71XuA9cUEBHWE3YHRpaeEGdfhdOSot
pKGSIbB++Zs26i4dR0eRggqnZmMQfesZX+Fi3oU3opd4N3SMidsDIIT7v5XnwjAM
ysozj8ZRmWLj4fLFAXjByWnpBVN+OsTkqCwdTyvOkc2zcr/0201mFpj+VfP6c4CI
EsmPUQZ5Eu0FhkU10oHzoU1qG4h1tl0UbKSAJ/jqDdnAMFHTIdfwB4INMOrOGrgz
eS7aeWtP/t2wqEoQ2xADtwndaMaSZjk4QQqG5+qasfCker7fED6XvyotRc13qyHN
bdZJfIyF9Zr9DNOIBQ75l23G/nqKgA2zByVACMM//IASkliRcZ6dhQWjKiJdLa2t
PrXqFyuJY7iVz1qYOexG3q4n/ACCQMb2K9cdDgbBP24e4j4oIP/AUniK3oOV2kqB
EG0NX1jXjT2/5s7arLR9sk15yHnyfbGk6ucdlCDqkRUKWl2NT3i4e5Tmfn0vfyas
GMJVVQTt0ieIOAFtuFmhEA0Iytw45t6SQgWLUy+NJCWIJi9ykId5f8J/7E7Jz4Mp
x/IBIUR1soCSTbmJROJFfXRtIQHKHBMapkHgcQXh9MyuDLUiOwAdx5Frba6AsW8q
v4Kcej4UFUvQ6KETn6CNyhimRYAmFMfEwtU/lVFxCO/60mnpkO1cV0x2mUWt3ZKp
Wu2GAiET+dgnLPybaszijmIfB6k7AyBOlUxua2/l89UeKxVscj23JUc6O42g1Zm/
yk9rFKjGDY3ZXycsHKoUooCSRURnUBo3v9sKvBfC0wCllv1oK7NFZsLYzCxU4OeF
q5IwfBl4h/g43rsYB37hLVHIWzOJbMzLMk2V5itj1fr5TBXdmOvW1UxqVMZqc2V6
bAPqc+BFHfjXnCAIFHI7R+/91xUt3HLSIqd/HpxtkUPYuG2L6d6PaaH2hXfZBLfx
jLgSeI0GsjRYsGp1HaEijXAisy16ZtaGFCe5Z/3aJvz6nmq2633Dqw0EiogYgBCg
UzxSu3Ule9rQnNuztSRJ8LirCPSrzsRj2gQ+Y63cZpV/uLlH6+zh9b/7ZfD2ysCh
H+VLUrzNXf5AEBTmCgCNYY+VbdF8I05F1hPmc4Dwo7aheG+vxuGwhO3XW0gmsd6d
Q0PqsUe8rF1PA58ys5GjIgyGrbfGFNUyUd7aHmvPb/wh5FyYsHaBPq+teSaeSESH
YF4mkLWDWOidkTlt1thjyQBydsrF1pTSrCztwCpI3MlpHDGGeLci1VhtojK7x0ss
DLCdUItZ+YLcvicmIq9nF0NFQL0lSAcHNsaGOHcf1bErwwVdDKRfijEHup3utqK3
z7ekj3xF4Dci2KmR73OYKLn9TbI7hSrhOO+tYEtLYSavj45oFNPMnrdPdZ0Wt15/
rtqL6vicwPVzc9/f7gOGNNRptEUNYZyD1nifBkWl1l9bqrhk8CxEUFfDVD9N4whN
uUVrKKPAciPf2qhPh1TLoSLF2AZpQRaSkCph7r2ai5HQHBucDEXsjX1Hwn+XOxCM
7Sa7Co30Y3AgOx/E/fhfMMGzCKC7pwOcCiTWiRAgAh8R1EIPYYqPEdn1g/aqFp0p
zkiCZXfJAnAmlF7cnjsbAgTs/YVuNhCk548rxfjHiUuGJF16HfAGDSAMzPYuvnfU
krOYGHzGck82olTzMPb+h00nYgWXFKs56IjtJbPuOPRRgkhtOrEXtYtiKimT8Wo1
2cAoY6U28LxUjwb/LNesu2aB6bnz5Buy6Ug0zQOutr3AeXuKhSXqcXtmJ9cnzm5j
QoIPPB53moxObx8f33nHj0DtwvaRdCmlrEtk3rrO56qoGSlcPmMadriAXlNV4Il5
Mgz8vpda1kp3vFzkEwPX7XVblhfKnGvHJ9VVHAMTNMpq6mrVccb8ledoAOSLWvRd
uLSJLhr/PpNaLghphWYtuBx/mDnOd9qOi6la4FY+Qv2YZM4NgZaBhBV7Q2OPSPfB
s5VcYCWduavfD2zL07Hp8K90HFwouaVX9DuEGFan3L4MR0Jfa/egzykESRLWO1KK
Gh9wJyed5dbz/+5G3x7uwy/oyHVyWNUpsRkLYT0mVIJS+ggtt6iLTdgaGuIid0M4
xKo+x1fotqyfhn5uE3+UG1wV2Jj67iC9A7AWOUyCoa50uhigF8SOqnOjahSruIES
24lao3MNADBJje37FZh3/en720tz9WFRAiGZVhltn4UMpw+4plmo1pYyU0KEcOCF
r0kEhsUr4sFfqzad4It9sOumho016J5qRFiJce7orSWhU598kC1BMBuVhUFABREI
BQmQnO4HO7kUaW6U0DGwjHR4olkOWbA+8prWnPGsKueH+w3aFZo89zDeyrCzxmi4
o+vPL3CXN8VRKuqsnFj4PGvTZQIqtX+Wpcsw80sVoBRvsXQ5zBTj77fATRulVLBO
duKOGV8M3R5cSEEei9xi7cpE/0UWc1OX6UljbbSl05YklT+QP9nvIPv9Hsq9SElX
6fF2f3Gb+PmlKWAlKl44efmfoFfXFapfBAj8s1W+TQ6UfUwaSS6NvaTIWAZMfuEd
iA+/qvbVoXOMmgj634UXLTvgTf3kYaVUmJkde6Fwoomm5LPlWQJMINHqxG7YtgrI
KWSmeZFMwa+BB27TkAjZrSChBwPa/KVBT0StFSL3nLRoYR08QLZDm/VBWkE2wy87
i5IJMSAKMNhiGpsrbIilJLLmn1P4esI33t86XuAX2qp5nQon21J5gaSLXMxj5fyK
TLcIWJEGOjBiv9PaXHqN2IblHd7iowKAMybxr0ADsvLqKLKrV3uwduJjIBbyUJsG
fsLMENICcJtjjHSysrR1rK/eHUz9P7Crjw7srJhsBbGZZmFkCTqeoFFWwIAgmMFW
oqKs+Jg8+ESGSj5EcCIuskwzOD5Sj6C7VewsooJmoLfZQIxR3Xfgq4tysM78L2A6
LW25Ioy8EGTuv+XxIcOyd9zmem4l8/8Bvv9VMKX9QtLaPx5Dy5DLZW+j1I0Zfxlc
SJgvkW6bBjptru/CuevnPhdB8oYbLGQ7CFZcYHEhXDMag8ThMn6CbtH1EiWzvreB
J4HI57Ftp8F/yUJGhsR1LDhKNJzNWzkG6qmQ7hC10HETeyDQSxkTKNW0/c2dZZlF
nFUAuORR6dQPqlZVQ/mxm5Oz14GF444yvyHL84YJKhQk1kmZpG4rUsppeernqeNE
5zpu5WI/vedLCHbu+IUs+o6X4GMvZHAV/gbfpiNPFaYwXnVcEEhe+rBTNW/MSTPy
S+RKpuQ0NB41KsoR3evBohj3AuZcmFtOMqstsxpMWccq9DHzZL6q+vQwbTldewwz
aDnrpFe8kXPuYfYqzrdDODgpHByamjtGiaWZX9Ju5ynpydtEryUCbPT+IqpFJy9a
tuOIXZfmmKRtcJW+F3G4fM8i58FP5NLgr0uTfimqve4JlNFSXMIcP8pyBbbCTv+/
kI9Ge5GQJH0if1HRLAW/1X6y0fGT/nIkEsQhfgXDOEPPf8GNq39zI89mohqGHog2
XnD5KTlUnsYHxEOSFPAw9ttsh2ZnPzZY4Ewn/SgySrj90Sf9OUDRXl9xCqD2sCj5
Lk6/C29M/TTB335hOyQKfeKt0SeApIo652O2n+ONG7AP3MCj863fOeCNFI3nhglp
Iu3roGyKqn+CAhJZ1mYBEMIbtPJqYZncz88B54H1qcc/C+ht7erF0RilQ30rlVEQ
iXkJ6ud30lnYPjzXqGobgaIv9HgMcyhorYBbF+lwaqp0oV8xC0Gto+Iu8WlczRmG
X5LTXnVdx/p9Zut8kpKjYXSodNJTjyrf7tsm+qNVkqLOPb+YBuDUQc8eFjIKpZfY
xqbDaMietkLtdjAyRzC8Ffq/E5Pt9NLyANvi1k0l7qtFL6+N3fFhkPzmwEmwtIyR
jNESmd7jlYUj1q2mHahFUj2OnHqWgQUu6DBkOWSMRUJ8mnl0xE8SSTgDb0kIU6E7
Lq1ftfYhTGnWMxqfS8sefsmPD8syrCCptDiXdT+wMxgfOTU72aRS8u3JxuSTGn6v
a0iERRqveyGONX6MV3Ju/+TtxhoKvoAoaTvwVoV6/QU/OYF6QXxizY2SXPO9Vfux
zKTW2DxctNZmTuGzHVF7zw5pIOO5uqB4SSeJUNsVbVH1cpxaIGfJ5dk4eiU7iXbx
C8zEaIeFcieUW+NGcTORffZ+tjgNLrw1H1iTXjuhMdsAnw+MmuAf20HZZP0ecCuE
dYu5D6uusdhaHBKVDU4ESVdot9TQQriaNKzUJe2FvaWEDLthgZYtmXjpE1/4pNOg
QMAnWIsrA9DX9YTr1p4q6XQXlsbGgv6eI9QRplRGUfF0b1MiXzhAGw5W/Y0NHClS
fJv8701oR28Qh17oB4yutEkHxzFbeCwYrUF58T3dTnRtbqpMCtiSpL5u9b/471EU
8lUVD6oW4qHYQajgZXJcLhIiyqNS13fgRO+RPezbNhq3bwkjD3NUqzOpZ58AsjaD
Vu8P4+1q81G+1wmiw1nF3HFnJ8P6NXn7iapDV4+74mhd1x2WxIYFUjeH+RdSoEZR
vgkEqYvnrb77o02JZD3EFhERKztjlhZpkd2MoNeAJIOKs+Kh2nwfLx/krKvGVQOt
F1Hjd3OWeYcTJjtXof5nmcitRHdncwakt/kM3Lz2quemHjhKCWP3qnhGmiGroEwU
Z9AFdlSQCBARy9gHB508XqBBImIc83TSoicUBm5nV2c0N6BmtnsRxia9QnyTB89+
zu7GxQ3QSPPAc/Pzd6ge3U4zDZ4g0Nf6ZCUzKZnqj6bQQDUxM+2yCa7xupWT95MY
EMKsgYor3xVPtd54iITYsmOUMYx0ZA1335PEo3617p3LI1p6lXsxxyXwSWo3s0bo
zpNnnU/hlogD7FECTNF70LoJ7wSnG2g+4ENgSVz/6wurNVCPdxb2qTYrzgCbWPcO
EPNHwvMopsjSGDP7hKsEz+qsyqvpeN5tNIicsYai/Lc58UGahc6k4Naeoct7qDeE
claG3zY/VvqcONMufH2mEdWzzbnSifXClWF1iRAeYleV+GRIb+SOZeeraJ9Kg0Wa
bfBAYjwFzRKKC2g2CxV/rJkrWNDYNkTDKYkJZXLiETiRgZr52eIQgRXe7AX42XPw
B0tI6yUmbvJpOlZuzoiyQStV4SlJ1bqNIkFcJJ0sHmfAnr63aNVChqpgJUOBgejA
WALdiIJflDLmhFZtYOIrNDz2shCDLODfreuTsTpo5aB6WK9/N/GcD0Qox5pp0Qyz
fNHYsABjJzVjdf+0HXFa7iUdiTl1TYJHspqn5P0Ig5nCLYuypc69s7u00nhI+hH8
Pr04DY9mG8V3LtwzJQV3ar+jxUVx9k1yTQZsLM3JTp34WXMQgpALKNcbCJQqei7R
WvYQvbnToNoL5xmrr8b+KK3sqJB9nXEjEd0A1ueJMVCwRFZ0gFnBCdP+TILnZV09
jHZ5Md1Lfc2OEspJHmEoFGoYmb8QvXRtlkFubgx+h3d4o7AwodcFkjDEs3eFpWHL
R/eoknLs8kihHxm4EDHGUbamp4FqcXFSrV2wSkP6pShE/HpiVgwcV7PjO1Dyow+4
YTQzyBQ5Q7vidimh22LCe1m8clX3+ZSjaY6ygicCt0XwYHUzktxc5T0e+C6g1utY
a20768vcd1SuMXcfrnXJFIZNcdTnKnAkOhTR1D4EXvlYYv/S+zbu+OU7kpX1RfYE
Z4FYCFqVoYkqBT2WIM2hw64Ut64vwuhlRelXODXvYhyFqO9QXqnOOX43fDEiB8VU
rkQ3VY0E4OVi8neZi4aQbLllfksUCOxcYX/p+luLwvJRRkpI9HODpFZF4jo1rB8H
iGbhUoBvDCnit7zcAw5X6qyBcb1LAmV8uiMjmZlMao7V8TtaAPqQD4ragE6wDhCE
n507g4MdaUTMV007Rh5Vghiv+gA/8c4Q58ikU1ddv7g=
`protect END_PROTECTED
