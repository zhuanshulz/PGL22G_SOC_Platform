`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T8NJMCtSvrnCYyqePgL+RJZB6iNGAhh/hakA+yxB7oYUOI7hutBCI2n//eQSphES
aHmtsWcq4QnqhjuYOjVQbe7SHRzTi1Hu4Tnn9rndpvoZThj36AIs74hDlNKs8uo9
5gNx1Sjpf8kQEMsx65tVtOmZlf2JfdIJeHs7P2zwOUFxafsCzXl7ES8OZyJWy3hW
/Dng1k4SQL1QmOuLdBpdzr+6UB0xkHkWE5b4Aq/SsVWqzWu3uP5FGakPVXuXZgUm
OzV+ox+NdzEgmm9jB6Q6AyRkFuEZosXNbt30vxo2ZomsISqecGrkHc3yljuN/xwz
yL9nF5Yn1CRzktYQOz23zXKDeCoDXpdSbMYgfYSaY7PxBN9H+dLvCUAPAgZoQXgW
YkgTze70W48QzsuYCF5qbeh61WrSP+3ILIXqf8+PEyA=
`protect END_PROTECTED
