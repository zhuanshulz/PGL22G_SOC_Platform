`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+SQutedZXIIxLSMrxtUwFrTWb/7ibB/nhIY4OUHlvJc0zvblTD5E0w6XXKsAIEm1
FMOtnnWBOJdNFzNLQIq5sHaA9Rlcmg+NLWlQ8kkleIUpaEKoiTTGqqkMfNJS73Zh
Q6l7PaeQtTYwiQfJctQJt4UhHVwvCnxQVz09zT6rLd/5jF10uJw36gDEaX4QosUj
6HcBD2mbK/VN2T1vL9LMn6i9emIPvik2osdqUT33pwRgPuIz9zTQOLvpwe8ZQU4j
6jMerzHzwLl1ZGvmt7QkD/8hTRoyvpELvbY+k1qMo9mrdiVKrzaPmbtux1J9NmCS
UVLDjtfwdhBU4GWE5TvxDiJh5fo4OCoeWYs2o6/ow0evJj3P6vXBavtF9IDXnyzI
vL8zWu0CJKnzoYmB6Mc2ov5GzE0jEmGTj273j9Zy5XUlHiAmi5+GxGwS6PvA66D6
wUldd3PScbLTzG4i8/wEVxkbZ/XmJAFgX6ONwiW1XCfLKVu6t4l0ZVzdib6Pm3Tw
AQ06scjIHhodou8x6rVaZmJ/iuqblmEqXVpRh8q+k9qvtpgGfy02l9MejlwUN68X
diddTzGQi8SVZTp9FyPmEnmfR9folvgNRxXYzk3s3yTx204OU5j5whXn1zsI1zPq
0WCwBhUorTNZuIlQ7TW+guVuzXCHe8QWH7MmmFRfCvthi0buMbL/KgJjcE4dpKkW
XDs9Ct2ShSfy7WuoyjGWw3N2ROrFsOTiHn6UUCs8D678z8LnTBHBVr5wr2v00nh6
WcHtPbFj4jFZ2UsdSIu2HAiTREsVkZk39thre1vLtEGlK9mFcz1NxF5+FdGx+jwi
otDFhxUS1ZvZVBsHfkmPBJXGt67K/SggjqJbId/z8D7SSXk5oZG2hk//Oio/+iQz
4lC0a/3HZ6XvJ/mnVZMsTmW+4uXx8RvkEXBC0d1hKGItY7z418rMLu06684xh1+U
lAEG7op4yb4a23dge17Iuun/v4UigB7vki/t8m5pCn0UUYo7S3wTKrIPmppg693/
TJiknPGpeWG3BEyOF0PRApdlhz/cX0e2sjVaYNlyIpldtv/zuMfylRKYO+WpITlu
Hrl49tRz8HlSpNd8fdcj8jstAhbIc7F7puuCqmoRSF+wfuUn7fVBghW2nQ2SzYr7
urQhXtWEuDjOlWOzJZL647jhV7wta0pee/am2196zzcAHFmaFkPz1NMYEa9j0EAL
P/1EO7WPr6k9RxTSmxH+0P5Jy7OMyCVvqy24w3y/rkL++pTjSO1u00p3GV6/iDJB
tOQ5YJZgTRWDOeNx+IuxId5rD1vOq2qRrEC80npHh5TEVZYe3CHx6Ur8/BrodJSV
qyakofuUuT9EFdErXizGhiWaHkUh8F5Dmnvf8X8rTXub99R+BbqHCmYKFHwTn4ez
P/dMs9Wlf+haZBLJWFd6/Sa1VtUFhEctAv2rfTMNbEbzAvookY/wGRFhnblEtJim
1O2sk3q9Icd+3Xx2Afqfr/gC/GmAJfXzXBm1sAcMwnJopDkKZGb0rCIWeAkgtWJq
aAk1USNHPZfH7CMe05z50yL38y34dio+64trgGVDqLztHkRzkhxsgB9cgcb6Xpw5
dwI5PRUv/jqXYR2XJPOA3XwrUtiBBKPH1xbNHZ5BW+cOsTJfBhpeihcvGeS/AxXz
c1o8+0OaA7v0DFBJNFkXN8tWJ2wfEMan/4R8sBkyywUD3wVnsPrVLB8xNjsXT+ve
2sG9ZUEHH++wRJbhO6Hy/8Iz7LpvMDvh8a+qVLFP+uhXubWBfumv6qxp3u89sArW
4AnPJMbCkUCZuwXcDiKatYNUW6ufdLXUrKgi75SvpNFRLsbYqEZCGkwh32v3mmG/
Wt/ht0e99nd/W/n6033QI2etONIza1CZDa6KdCkeftrLsm3SsV17BL+VybZKMyi6
YqFlpn7reC81o1I96OlxGZ25U0wsh+zKZPdPhqiqKLhe3FKX3bx9vK5O9rIzsa1T
xe+y1zoHu5VTl8LiJH2VMv+WamSuvrkEED4BkUTQeuSPjhYds6MvfuWgwOIF8MsI
aBXvO7mfvxr/5vfDpl1N/YKQ59UlPw0ISclmYIAbZEgcsAhdSkYZKY2NR1Ih838E
vYtzQj8FhLBPlfF2CHRQbYwZiE62cpq+99G3jNMgbCNzHIEP9IUuadybCaw+JXqR
/fktfcPxnY22cYgoX6YfZVTb+9SaIoXmO09jHEbJNbcoXp0sgX4TYGDZXjSEI4QM
mS+k8Wmf2FDhhfw3/QYxg91K6NP+/maW8x/G+QwcOFe0N+1Vk7lS3iA3GLx1BC+y
ev/Dgc9cEYP8T++ZhCYF3PtkKc1/4zC73HL6oO9TAmlLHOEMepB0wBcJNB8hReNF
tjsODOVLwC09QUAskdwjR6JF91kAZes7U72uJls2PR404ZYv8srZbxh085axwgRN
snelWY23buBIPU2jp6YrIIhCuNf2lCOaHXJJ9j8/GcPI6Wji+lEI95F3SKLhavlT
UL8OwVNL4v5OJNnQIaVS+DKXUyxu0vvBDK4ghv4jF3S7dq7NiYBjLQmynufMGkCh
g+93DmUePymnmGvGHwCOiFprWRJ+lAuKOICZoQgwiu8P/He1Rnt5RdS3qQ+kd0dq
ym5v6hivzmuHtNx5067AqHfKO3/UGEE+3DAoeqnzJTc0iaoYMBEnNd4j/5FUu97F
w7fVylQjdhDkN7Hwh3iALPtBBhA/yJNMI7XOS+VuNZqh6hI3iyhttO2yrYmcoIPN
4lygmw4CbKSxLyQkPMRhJfW3a5ZwX8lnfvsUIeSWFDf1ks2jPxI5FvAMrVQ05dhH
l6/I18ETFb7uV0IkYqCDug/e6tF47uFsCzpNrubqAst4SjslTROCD9zIqqtATDqS
jPTzr59y10WB0LvLZoNf7e4gtCdAxhPArly9L6Qrb+7rZ7aJqMisyv2a5nQWJufa
6zgw4yUM/yr3KHabCfLOPX/+2bnjuGx3baTQfclm7WA3x7bBye8gKO7neGhXjhEv
P6KIHvY+CrwxVEA3ZaLppr8A+cb2mD8Qz1EtT2VXfIv+oFY6XkiUG0+5llko8TJE
WgXQ6/xu81EkiD3wlbZyBXJDxmgdzc6eHhwXYYy3V4gjv2u8orziNHHbYPvqEgKY
5jb7nNCVLV81LBe/FIbo3LHPRn97PFZM7+S2JOme/WDvJNw9vNYSkNkLTbiJ2QJF
3WvMpMvpWwTh50kOAvNHyKWLFejGumhgDfKxZVjTCXEXfYXx9e5Aq5WiS+HhrThg
pXbv2hEeRIWScwjWmqqM6a88JvS1uq9a61664yECqz0UrzilwBPOV4m/KnkDmC3J
Ie4yDHWBJXSnd6mZ9/RPpr6ku+rhl72hDgQzRBC3K5SGtnKysInD++M31BZgoEds
S5J/YBLVlo5EexUyUzHMM96jPBCl7Q04oMEta7EzBKC7xHrDgHoasLE0Qr1mJ3pA
fMpAcrWkSbmCBZZhE7oN7fC0zhHDJGnkYjKSQAmlJbC9L5zFV2CUDmTlZOKdHvH0
QHFqNRLs0gleOqsnL+vNE7twLOGex2olEV54Ivd4/zid0sCHgtO3yRzzC09Na7e7
dHCYHUoSgRO66TcKqTu2HJIcsHJmnGkOSve9ubNv8Hn6u2PE3ThOTzW2XmyhaTQD
01rnw5QCZGYUQf2A6gLHMZvZtDa5mCKYMf6/uNLUc3pvNP8ITnph/8Ydox6JTU81
Y9QEbwgVpn2ODHP8ppX1rSpILms/O1N9GgM7321Nnb3pSA6q8cnT03VBg1i9ILyH
7UUpAxQL7EtXJLqzZL3/fTwOVEIcvn0qgW/0TWJDUPsnXq0uGyCzkMzvsQ6ReU15
urPCr3V/G+UM5QdkOQezUbYg3OqLNzVVhPj1wUVSMEZ6QrnDW/heXbitbefy2kle
bBN4kNCYDaqMZ2IA9Uz+u1wrQrkKgOfkakbYnl5SoKGIOrH17aPrFFrOI1F9MWW2
DS+RKkJYKec/hl4d55HsUTg/mcLMz9Wc1XLTq1OtQnAdOoZxKWZE4PUodciLe15Q
7oxws9u9IYB4HpWltunhgbgAP1AovJr1oI0EJNXo3OFeuYbm8eKKuaSOUdjFEtml
daunGhiYSrQOiZwRL1OU2ofe31FDTfT8NVsLkbRM9VCyRhc0uIvVQuRJHg9oSISr
J+vq60Cvhf7dsJM297k/aZtF8MSObbf3VNgfzPdKulAfTh0UjxABWinLAJ9g/bJx
9kJbpc7rNJyVZja84/NkVK+kpLct17ptTzrqqf6RS/m2Ovgt4RSFh3znI0OxISTD
WzPfnHWLdaj9G5ds+8kHgSb4uu1aEhFR/x7N8yfxmFjXh8/jhSZXcU9BeN9XtD/E
8wOSUVMQ7qI9TB8holpFH6v/+QytPRpYD+9IxZx7M5pde36JNA+bLiw/yrVQcOad
iJGaIwjr5V4TpiXBGjt6N9bggWYQGvusiGPIpL3hjdQDeQwx62avOU0E7K4ydqYv
PzFRlErom8Wz+ZpNN7usXHntg/leqe74mzBtF95atDazsx0pUGErQkZfG419KrZO
vQmkBrx7ZW4ohUoh5dHu5ihykx0GfnlyO8lPxDUeTaPoK26orbjZkjFlmLo8scpY
Uzumr0Yhzbdle9AMyXxQgAenfrjp30NJC3qJSyuxuIHTWE40RJpD594Xxw2E13ZK
HdkftIwlpJ1QN+I8bXU5Z0EFci1pciShW7d3gYflGwpBRC87e7x5kkOCfILFqCdH
+2Os/0w4bYHuFBycd9+qWNN6txY+HTmsWKmyerItx3dgrC+HHtjRWq7VbzLP59jP
MwbCF5JFuoTJWMCmlXCmkuxBUiQgl/oV2QtNmx0I+JTn19O49e2cI1kXGVZX4I78
3gLxMuhDAanfdNZ+NccuTzfd+CE/E+NmHeU9uda2W+kkEU4qEuowDZOAZOk7THMW
HcQvOG1aqJCkKZkmBbvObWMDqvUzY1AxSi8T9e/jnxep11lDl7m1zUOq4xSPSsLH
um//FP0R+s4oqSolAQstDFClw7+3mLF7OlTGEYGQ3DDBY3B6rTOtEu5rrp/ZaOGY
nPcqnuv3ekSMmful/AZi8KFDyctRA/3UYnQpj7y9UJBoo76pxRL2zSYseWqCxl6m
ytH/ZcILcnbFDbyTvlWm8/2VQ3nGoZlWRVYQ3SS4gUR8LmP+68zlraqso0apZOFY
7Fi8p1chBhPvXhPOtcIPG9K3kuQSFAAEGVf8D12SOBr1KZaetrQxkNoqwhYnebpP
IeG82XWa4xTsXSGv9YpjygiPhQ3odxbc7gZypjuly4C/yZE7VXexJELiJ/yX8HBd
vCFVsor7HG2xS+z/kqYdCmtyCQyeQulwsWQTHRdPsbm5lb/zRs/CNGnqnOW+r5bV
w2nRoH4kPX+/09zQwXBg5x0U84IxnKJR4SksU3ROCW3LCL5+W8X0am/ZV828xwjA
dsN9jU/rZx8/2r6C6RStzUrenpMDsfYEnbT+A/tzWjnn2921k5Z00CokVSor8A97
zUEoOj+BQ1YASl4FOQXEOOLomMvRonZIHKT+P+fuSmMF7CI+W0ccxQUqavFV7LiQ
X5CBUQROlSvOmwzdecJPQEMp/6yiDq0DdZyVRLTwaDPCs8vqyEinFoeEJojVaPPW
L1Ujp0lYp8s1fciUfnMvtyRSK9/fD9fXBjyzgAGjgVPl6WBEHVfKVrT5ltF39GsM
n4m4JXusmyTn6yG2bRp48Mn4ptEZroQJOFLv38J8OUglXDiP+8bxC3zdrMJa26cF
gib5XsXe2QlISG7IMtOJ3iy+L3Sdhwm7tVEgSx/ccJGvwW+/fHLvLVR+BMr5L7Vw
Iu+Tc78W8l4iAZARslrPdxhQ71Ithev2JrufLmrdcCcJTtzK3WvId740CPMeG97U
qu6/GVoWNSdZUfG4exRFsFTTdmFRTWm5z6BXUs9jqil7p9Hbk1DnHrY9W6fYVDGn
nomZ3g8YI9XjI6gvR3uHF/x5o8Dr4Txhkc9qFBVZYbI85ePXHinrTIGS6bYPrke5
pTb7+7FEPamP4UehMyfiMlysuiCoC2FBP0uJm/ENSP7OtMa3e6CRBdvLvhUb/qgf
73gdwyf+sBK2EQe7rhwPUA==
`protect END_PROTECTED
