`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rta0iJETNjfF5rEk3PGS3rvIUCAOTAz16WDRxFRBF8QfhLJZq4wzauXgveISmHM4
BnSfU0fGsehZj6H++yZZXXMEeMfWuQkv2jQhgHjlKwPZ9FcGKmugz5TEx5PCD0ZV
dN8843pbu6kfGvNXChtbod030ZW7Rm25o5aabECfijst4rXBdCQTyDUo1oI7vgNN
jYSBwlcwtD3QHCuYlKy3uJHMdCM0cNuq7ew2WILrvTpadrYGUFAl7F+jBatAZEuH
BJpr5lcAs0mysIopXODmB04qqJkZyeI4D8LTkCGfimq6BuUQZj0E9lyoCMRJp6/o
+VCm+duY3iHEUlOtR9c97NgdsME7bsWnLk5GpqsIZNH/6XyX68JOy3T3hD8+aZby
6wgG2B6x8zeCy6Nl91DpEVoUgafJ6XPi7vOCuRkzryQx+jWabVpsxgLlQIPIquSq
iI4/hRfJ/W8uOLEANjNveJVuS+ZzF480TpCmLhBniqS7jJPIfRZxoBQ2aPbprZUg
6qR0zvx86Y66cnksL/PtfeBVUjt2aGfirH9z/r1DUMg+rrrZ5wOilyTQuX/vUsvq
gxmBRW6ddsqIIcVUYwgqU7BbgaX+XTAGedqwDsjc31+ho2YPcRe4neYwu8su4M/t
2dm9PH9j60mdTjlYfeorWGZjgpvFsxn5meXKqkPaIEEMApnhQ43Pz0QvcoDXX3Oh
d+x8EEQjcOQPRwrZVVAYHGOJqeJJPd7jtJTI1wJ6mpK7MFTKRDzAootkA9K6+yKw
`protect END_PROTECTED
