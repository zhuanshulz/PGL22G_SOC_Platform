`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vJ1Ao1M7rjtd+1MRcAg5P+0LbpfrIqSe5fv0TzHH0CFjUZNhhn9IW2VixAskTL+p
H66jsf5VYekS9Fg2yEukAsZq+DOtOCAC3Hkepm8okLzZtmpYB6v86mXkeA2Y7Eld
Fk+y/C8uqLIG2CplIx3vTANOSmgjklw/5V3uYcoTGjExf+x96psbz0Wpa07a7iA2
eCq3KCzJYdaBHUiEzj3yr64XJIz3ZMug+/xla9VOkQ78jZwfzZrXgr0m39S67KNI
D9d0k5hMHUBTkJSKLKg5iO0kA5XXjiuCORWaWRVPxyoyX6eEm12g0rk9H50BS4oi
NoVg9at0y2WTTCjEYKqcOIfnZkKPHTjzQSEFq+hWTfLQx4buCZ13L6ggeURJswFU
lmumeT8nq+Z7tBdk0UN1RXOPtsb4p0KYl+wbmukeFi6T0Rre+AzhVj3x0Qzb+oy5
jmC3o/EaHeLFb+/m0y3wZzmOzg9ioWTKFR8YbApKBASelL86VEpah36NC6zJtIQt
gLukQuhCBa7H8x0yHiuOiDYUtJ7apzhbuoQDKKSO9km+iqdmo67qjTSi75iAKbMt
EXZso7X/dOi6T+3kUTowQR2VxsS8jmNgATqBiX4EGNbuugroU6FXHdVQUxqInSl6
MHx6uO0KoZVvT0craHrg5gwUXywSy1091H+bqngD6cr8oAa5ONmwYGXwBCoWsv7S
qD+yKB6qoQGiioHFU22WkrPLxolQXrw1JGSGl/jgzS17HQsXrSX7/UpZH7rcf3jz
EDl81+NQ1Gfpc7nvwk6MZXUAcWmv4R+SbGpzbrZNvsMcoa+9AJwPVbnaf4628o7I
+759NCEKTnDyZsGmVxO1vfAmQ/trnEQMMEWoUeP6aLd9SQ3Owpaum/IcdLrAOlL5
s4p+Pi/2hIt3wH6xh82rgtvly4H24nWe4dFZyITOe0NpTR1I28Qj3bCEhfQgqA0j
s6qpeW6adktvXL63nmUU/4StQa9fvVxkO3AdQz1Ds61n5PpuCP5yZZEnff4+6i23
u5GQ4QjyIZQF4dsoej9ygyneJN4jEa8isNpIxIhGJnRR3PmWVKeWIGXvG415sbpv
2tDcGH0DNnmf9xuc7D/6cUseu71HMxJWJi9M7tGCHrEMBWdFHV8SLvBuDWgGaQBD
rxNQXxyGWCGIREEzKVG/rb/iuy0IpRNDoXRi8bxKfkIu+1XplsKxzXlOB4WOa4qM
J70KKN1pwEJdI+uH3tcu/s+vAhJv9Yzqt9G3js3g4yhrphrtvg9itaidk+7ewws0
WPPwipD7OBsYky6J2M/DhjlkPhk8UtyDvqbEgj7p5QXq0g2udFbnUBlu9okz/iuT
fjpI5bZ1ZUgo+2InhCVfZE8ZMijNyjG8ZjLhcUP6VIe0J+xTwTNvEFCJ3L/w17rk
6rKeR3Ix8BKuYg1/JZ/VDdyMppy3Zhq5R6QsgNFDvSdN9sr5yZvl3gBMTMICk+if
SlHK436oLc6Vfsi5kQtfnc2WMB45i94O5PNqAxqnTG8zshHLq6W2X9purEF/kil3
4Bl0/3nHuB6IZpBZEtOedfP0sgVguzKTImcs3eBcNIE0Ar9MrBEQ9Uy9YV7I1l5U
SYHzsaZSZcrvgnJ40EAS4XpPyQ4m11l2l6NGNj/h6cvm4uDfvGnno+gTm/o6Tuha
wD0t5tZJqeIzGL73KQsnFp4SIn9Sx5V7O3PwJKDbtRAhqW+eX4f3231giDW1xBbp
YIIItDQ6/MoYUy7TFVvKCWNRhnNoXMDQEeKd+awIZn7oggtm2agmEkUsg9akqUW6
Ig974rJAWz/GJuJQEktrhl5c+H9RHj0WM5Wn+WWtQrSqo0ZeLERffF7GXcoA6oQI
QtkM0R4evFO6CmMprbgTZnFuKLKM/Soa8/xhVX+qTlNGyJMsrlyJjtfkobE8LFPe
T6k6Bg1UVnGOh0zafXGnJ16lS9u+g3AaF6UHsQb9uIIQ61ePgQ6sstKzjlGpzgBw
DTwZFltETvPaH29x1ZMZCbMnJrfzEhilYgLCvs8uj43dXX4cuMHG0VRIrQC19xQz
4ca5ttwkZHFTcWn6x0L0WYPwABOehgo6X9PGDv8zPoGC7FdDm05QuHNpDKmcg3RW
jPdC0ZpRsESJB8tI1f8fz7mkmbINHGOMWpVpHsHUMCWjJFTDIlmTXmgbDu0Gr4mb
Liod1zHkmc9O7pbQ1naCZ0m5j2S8A+NMcRSmf6TA6QtIIN6SPzzY2QXG9DROsJ45
vleq8WUd/xASvNJPrrx0nyt5DT50sWjY5opN/TyNH0bb0PR98TVuc2dBU2wCA/Sn
Xo7JdISjElktEH3tZNf92oqgyoJJdkEgUgTbK13YTAmGaJH70JweA4BgdjLhDY6w
+ZBSb5gJtDmu4H5N3Q9W0wFWEgFFf5LTbDeJOk9yJirlEtejotPcrJk/0MEEjw77
rc5CwvsnYvnMjcDc+hX7UNuUOgCziZgKf+ysUc2Q+KGn8N49P18daucClUnRQvEj
KvnZIK1nsqG48sYyOAEyUNZ+qP7kAE9nh43aCMQ7oo2VUO2lYmuubmSuXJrZ2qJJ
FqONEHiJW/Vqhxz3kHkDdCAoSlYm9V5GeFX+slVNU3nmULRaMkNHUl3e6J2ZSjhh
2++/54wGj+nhcc6cuKsS4prnMnibDHLY4Gw/t1BePAlDc95XhsWGqz1zHmmCRk0L
s7PimNqHRGFgy8ryQoSFZDueI0KtJXMp/8ceKeb6uj5dTgb63J8kRs0m0sWCMQxy
8kUarozHrznlocEJDQs1IfXuVBtXtvBCbyINDEUffzs=
`protect END_PROTECTED
