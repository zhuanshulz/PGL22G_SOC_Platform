`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W/t8IIReSR2ZBRtG75nhWZOv7Sbz34tNN3PVeOODn4pFdADrQP2H7m71NKmgQrBA
oqG3pvICfXb5qW2lH3LMqYL3xO5LfgTtT2NSX372OS0IHz4T1JpAttNj22/q1oOE
ow9TrIZBMYcLoYdhjniUGIGZyFr2ixuYnlbOv/nSOz/X+VHMxE/Bsm4wOaDyFviv
31pXMjpBhza1ZulqWJ+7HSAkE6NPIk669s87l7C7mdNMzGpzVMLXhlx12sIsJtC0
Nz4on4Co9X84TBAtzlhJ3Xx4MV78sSkF+6BnuFS38jXRt5Y5mun7OEjz7sUy4WIx
k58gRZZRuPMEFmKVSrHCD7iP+nlWcMPpChX8tNmMKzlBMAZrPlkfSnWnOYon2gkc
3vOpVhnVRPks+Kcoba1QiTp+w7PxFL+SBTm4gGZQ3UsdwLWkTLc/CZWjVA8Kqu1y
rdddZTv8+VDOKeS6n3WEilSFL0ZfPUKS2Xx7mnGAbnPEJ23DTNaEVhjiZUchXBAl
+mL2OERbiRUoxKAdbd5rfQaXvjaXK/YmunAQ02r5tF8eDrb6zaYH2xmbD2mU+Env
s0XTVpee9eQ6+3tSJRz8AePp5Fp3/1wh+/pc0nydQQ37PwssCZXjj3IBjWS8vu+v
hJB+r9WIVPGt95eg5HHcUvcS6VELcDQlvph8/+/LXRylEf8Gxx/r41WxiOXqrPZx
qyP1yyIKiJU1LEFE0WHq5aEjrDdKv8tj+1ZV3Ao1IhqswAEgaMjyk7zBblNi8AUn
ijGvmAzXy/NIl4YtiQkFxPVncXuS2N8ZORQWJtRqN81Pzp7ZEylo7kYcA590gyS7
adjNxD9MSbIEzzjk88DbR69jM0dtlIDlJDG0XO0cpoL02QWIJsRRry4Pp9i5ZxbR
7/YrO7vhXvvfP8DlghSpj/k22MqZg4IsBz28A3Pk+ax6BVGvUE0NYq4fo0gh941w
`protect END_PROTECTED
