`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7vJnQq0rdWmyxbBU3xkoy9c+aiDh4zo3QG80zIfVzMVrgvWVYB1qSrFC1ke/hP2V
giY+ItP+enTfLpKZeOvAg1Q0+Q+3PVXFI7amjBp5kHBQSW6OWwnc/D4gJGxLC0ja
V5f0CE62+fxZ54Bd5kUZK6lbKxF5tfzoHOyno+5wMKL5CclKlMfUId8N9ggZ1JL5
Thuoq7k09b62xaKth/+SdvsIkHisQjVByxl8Ttdpil+y2/l/h/U5VKR/zw5xhd5W
aDPCnpmqPcx2ZsBGKWZgDDCr6Uj6B2Vls1WGYe5FceGQu4iOdsX2yr1NOylBhUUQ
qiXsCjdEC/MmNMromUAWXeT7xRzyd0RVunrLukEaEOdV3lmXNmzdtJv6met7BpSh
6lEKG8Wbqd8kEyFIK/yLiz3OXeah/1NOZuxOLHGHZnkatOOza3JI/Ibb5EsfGmYN
tvbIYpHsHKcK9hGkay3qtvne73K4m0pqc/A3pcJWPeTZjJCLP4p4CGRNiwtkl9UE
iK+6R91W2ajnhKRtn9tyYiGssVMAfSmG0jLL98m/DVcZNIrJ4nYf7cT4TtadHqrb
WdLLoZbRSA9s1223tbqu0A==
`protect END_PROTECTED
