`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1LypFzXtrAWQt3rFX+3XDIrObMYDzMZtdEen/tGntl+uDlZOZqIRY1E7RID32Fom
19GDcuL3qsV+oioFns73sVoFZE7uFx/dkH21RrXEnyByLb0tPcrubAjKkt4XkLXW
kvfrVv0sU6B0F8DRdeSqrW6gw3FP1b1bkUOxAfsZCbQwqC36jPcLqxsSGcBc05/q
Tpm7w5APj0992YiFx1xmJkZUacrwdiZMuMIWmOL4lY1JhQxKtb5t+eWJUKLw5P8b
RfWuMZdGeTTnDtyFAGLBMziVFJdj746rbBkRH1iacImwWOOS2UZBbg9DvYopSu7O
GqgM9YgZM6ALOd526l3giWsGZtjBGEGiecO/rRQrBAvmtHOIxqpq5Om68BV2MnWC
3B9Wj0tz93UMl+aXUb4eQ1ozsZbZdAm0HzEDVD8qOJqcRxoj4G2PS7UPl2wHnQSo
KFJ/sc8aaKytBSQ52n9L8ZbdtW+5XmfsSkN5d8wA2mzaZZHjknDcSLNkSUyukb+i
i5p0Mi0wqTppfNfWWVGTxxInpRMm7BGBeY1EZ+PELrRkgFdhtFJq9wiDclrPfai5
`protect END_PROTECTED
