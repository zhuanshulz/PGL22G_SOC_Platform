`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DUiNrcN/FkiCx/5i3hkpXWUerP2aH4zkWPCi3ZjFUdOPnrwLmYAYm3k6263IY7qx
EkulYn4DYL1Ede5J+Pi+nSeN94PYsu0+n0kq+mTSMTP+MV4oc5n1cQWqmUq8SDZ6
IyopmX6IxxcQ9W9sLypS4uHYDlaPnTsyneU9HzEgaibiKbnpFg58wA915ZFR0fmZ
QD/tm1Bqez7cn2QwCgjNlLFmg3Ezq0fafWU8cbqDlyNrjTVZpmd+QtMwGZ7GZMAM
4HlxqAv443zxS49rn83yFOpxv6Qis2pmtKnG5UNcSHK8O+IS2dV9PnIz8roDTTgm
Gkajvp0ybG8MD1gAOLnmRJGPH2umW0PfKseNelI0JjfBM8d2FLz7KHI++U/yGsJl
s5I8yBppkQ+5DbE+RkLwruEcWQTED8TO8WAAH3WH507GRKULoDkwA35AENRE7MHq
9P9SaTV2zVObCBwWG1ezEys0yLQREVTC07YrPBZXk4a9pW6Bpf3v4hIQrjZg/oY2
EVf9X0+sI8opb7kbRd7Eui2exWsGSKkjjRL1+zJrSaEMD9ZxvIfklMuJgA0GS5Ow
UkTlenetMA8qzS6qYg6k9WqvJ17TezJIm3U8562MZJdyNY1UTHnP70aaOhXzpZGz
OChcMrgQfvPU2DD0to8/Jm+w5jKJvEur4XRIt3Q+pf6j25kk81EVv5u2fScTqeLx
cPJnqZiPADd1FwZyvH7nHPsd77PVK550TSNH3qlegXVoI9VnMeKKp7xILkb6y9ti
rMDE5/TZsUBvmJcni+vONpnKhKHFFaYfsqo3m7jCpgSxAQU5Q3EgeMm63Mf7IGXO
Wz1dztEMBZnu/HfIZkZGiFZmYpHy5mYT69zYa9YxT/mIF+bTBPRGTyNb3IEIkb7U
Jaa9Ttc4hpV54Cq5/f3HTBCGR6DL87dzdU4SAF+3Rk6hepNWpj40ks0PsuP4nseN
rrE2ENJPwkY2WbB97E68+uW36TAjQPGZton3IjWEDPww7KXVHNQQ1JOrTUuVNYym
IV6/hFXZEHedQ6bOeR0zZCW0df5gDwJrimQf3QboaOGYcItK1SiaUydOqMSXD7Kl
Yok9VWgAW8M9d73YGKv3o5iapnEZEcwGHMGG7MYgxUAu94IoCG1lkpL5LS7/kDZx
/ZJcz/jdLpTgrVJgvMpxn0K7ydeYbWBkL95jlPnovpNHGvIh+M/lc2sq9IBnClCi
KbuQ9QNpHtL/AbFiIsYr2zQcjOXv/xfag6hE1UCApWkkBUVpfV0c3S787ZIE9Rb8
xC00Mh2nzVVw/FmV1UZyo2h21eiZqWGqSucRjU4PwTbXoMnsStHefSI6aInDm4Kq
tRwG3g2A3bmsd0ZsMQ1km11ImB0wvwBuecX2BooEf8zHiNYzyjpPwUfKRBGi6xhz
`protect END_PROTECTED
