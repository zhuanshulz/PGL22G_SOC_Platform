`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZviCoSyvzmt8dYHZw4DZhGVUgHUy9Ai7CwLJePLLXAoTJH5rPi4uiWnPWz/iSRtG
S2GapAtLTSQNAxnWln/DEigv9VlRKDS20cxF9l40/Jzz9665Moi2VNQY4PmlZ2FC
5v7LXfRcGIT4UYHFRgKJa2n+KbDsTHI8qWLsJ6jVcKHuSnYz+mtEF0z30mxPjw4D
aJ0B5E4gg+jOG3R2NxCyxUK9CkxT5GAIxWAIG4Qhl14rnAWtbdtyf1e82daG2OQs
wQKyLtoQmqI7B2jKxQrL4LVYkOLpWmQxZLHFHAEGCGdYf45wlaxVUCPuemtJ714Z
xpcBmqxsct4V96wqJFLJHh4ds/eAjXB5SrUyRDtU7vhrtVRy8Rw9qdCxW94vhaRO
gTHqL4MKiV7Ss5NOu123slljqvYF+Bh9bpgzSgJ86LLIHp+2fz9YSi3TT1pQT/uz
6dfxnSId7AQ4OcSJFl1gWV6O4DDJsFEEsN3xxc++olI6kip4cNWNgodz1t8LScfX
iSJRH7ZNT3nHyyUTAuOaelv7eXWDv89IEf93frnGpi6dpZh8+Na8bY01jFmi7IUH
McsF1WrT9gDEQFxpR1EcyC8yNVHumHFEC90bAvdpf2Ooj4WMWIGQIGTPY+a0hcVz
jePuGCyXH4eHfKhzbOP6goLTSKMGNzyKHI1gWlsD+8jSkd8EVVc58afGAXMCdAk7
Yssw8koK3B6d+znpYS48HuJFdfyK3pK57HMVZwJbmPNzsYNKbiUDzbYEhTPJzTMs
xJD1a8GD5nGgdffYl4V3yFbfDFacYN8jA/vv8LgvKLk=
`protect END_PROTECTED
