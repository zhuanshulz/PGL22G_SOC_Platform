`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
twMmYKZrvwaPEiBAaIvHXj5v4EbTd7xEd/kmNExqk8CGWq8zSnM9hmsZqzmyK/9J
jQybz5Emg0lA17KOMbi99Jl0MT1EnYZ7gbaZ/iwDnFlnjftM6/9Eag/8L6TFiwou
uo5KogepBysFnlR1szFGJdEb9nxknvmFIxZ9SIbLDzNYms3bSrf5SXBQ/hqT00s5
tDsLPVPgdIKjCER/i0bs+jhCyD28etucIgZrdTsMoOj1+zK6BKAHjmTTTVLawy3z
6A+Zy3RsDLhn9GrKFQhenEi+/hItvhYGvy0OBoCFB1AczCmiNegBn0OF8Ll/m1hT
rudYYmeC5wEVc4PX7/KyPxcprb7X6MHjpb1XfO2SzfZ6sVhEN7Nv3pi/uQ5NL8LC
OCo3lHeHtQnLZu7O9uuYnCRiYBZD0aVa0plpO/bDWPDA1WDAV9kXdXVR7T/Q65Qb
gbcYBynilBXocT4/IvTUyzxaTr8HtOfftAJESY9t+wpZOmvgbyj/LdUIYFwg+upG
Q50mNyab80pxXhsLi1jpGOjD4MQfHGV6ZkoXL57II217AjGZvdUOIaaXJMVnPPhY
yJxwkKdx9RAGtkYxpyCHVg==
`protect END_PROTECTED
