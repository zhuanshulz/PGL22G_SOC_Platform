`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p1YAKM9GjmlhNDNZSMI0vjPePRUsALWSL5f4spvt7lm8sb35MRvy61xBrLhWRffn
JIMZhfDgL4igjG+qtotMR/Z1o1hKyJR2oj8Qf0Nhjhnc/dxCUPxqACDUGx95dR7o
hIvBJobLYXbYfFtCWy5ZKitwmUZOPeWYwQvWorKYxL1BjCkrB2AAi8htrdbW7vAP
SMArwFE0ZwZ/5psws6ZETXfVcIP6KJ/3y4G37S5fDlyZRy059L6VvtVwuxTzqSHM
FL+F+r11130lY//S+nJ8lxktC26Tf9aP1Im+TUBjhnAUPITJJWsv7x2QgKvDZHU2
HDpumtP/J/HD1aLmk+gaQe38eob+eBnADx2ycxRorQtRRtOTfmADgKNnGs6zBnt0
2sFxcd4euRTpU8t/z8kTF3Ks3doLCMmdFMgnA6e0Xv+cAY8lEu/TM9gu09xgPxyw
gvCd6wW50/V+cD+EQNUxMlo3CghFEKoPfwg+SZAiWmYzuWV7v7YvHZYb6Wis6QX+
WiYalbRSSADcF+tIL3JniM4CxIFZWDIvF631zb83GeCzkOVmnDZRFPtUTtOLPcKJ
cIB3JHjwoX/0Wa4b3YhkQdp+Di6p5AE283+XKudqScM=
`protect END_PROTECTED
