`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1iGgtvJDkOTb6420d40n4bcKcZAU37hpZaGceBCEH0Zqf9LbcnSMmLEAnydB1D4U
nr/7YX31EIWMV80gW/XsW7+Yxo+5lfUSbHv5tYFNernXJgZPtiV5R9Fe1kzpHNY5
dtkebt1vE7hNGOLLCzU35CTDMau/D66jnMzuj5PjwkE1LXjUv5iLcrg53km50thd
Vo7WUL7SMMpMlisega26oaTXpBwnjJmnbjZARGWEIvRo7utxg/Z0ZOs3ltoJ4X+U
m34OVxSDXlXcOSHacCY1msi1AAuscgHBBOlMxB2tq0zCHqxKlIxoR46YAwVFz5ef
uNPc7lxkE7RXQ6dEP7hpEubprl+gPz7kl7vLHNyDhBs6bDe0T+dOMJ8+v6n92x24
WIJUh08U+QJI6pMtX5+KyxJEgJ0foEdh5Q2eVD3yLejFXr4PuKBcE8vxc+pDUOvy
zkOwhHXlNUngtAJnavP5zj30hN+a0LdyExDBQHyNljoCKchtXO49Fv4mENkoEdeB
ER3BIV4cbBcxGCk+dHcsDCuUTchLUTtEu3WqH15GRuAP08+QwdG3OFRdT7eyNHy9
qJ3yyS1iKIcqtjK41+I/Lw==
`protect END_PROTECTED
