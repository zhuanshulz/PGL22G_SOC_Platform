`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2ge7i+Q2P89L0kU1vjxCLYEq6pJWCei12DnSG+YWnv6vr3oKdf+Mi+F4jupsR7q8
sG89tet8FYKX0ZT5d0SJx0fACfxco9yB1lXSkAjIGkk5XbYs4NvzujR8AGwmAsbQ
wQvzVtKQXmEdvtkpcVY5NzvJLNbXR3guAY21jxc6HSLA9UqeLwJQqdNHS31yT8qE
/OSTm8KXQhB5oqoWBPMNPguKUFqVR4wkJDGRD5LVcCrLvWKOe6M3lYsw9h2ODtN3
0JG+JK5quqysG5ZHnKsMZc/BRJH95BPuP0zRtD5PY0p3quVn85IK2Tap+kggPu2D
Tl9r8/tYPH8uZ2ywZKQSv88GQ6Kty+Ppvmux/iaecxL3Y9ECdrI3B0DeVRJoEgdM
BB8JL/NIvTAO5Hq1hDOXzeAjh15vaSG80E36uuGifcKspeYfNMy+AqMLPXMR+Cgy
i5FkwRFefzP53SimJEb2r8jx4wH6x/TKYRTSnfr+Ef0J2FfKwqaNsDRR79VQR1Ds
i9KazXf5LiKCG5F81q+oHzJse04r2y8yORGRup0rZiF2Cg/ftK4382jG6KuesFTg
Yb5LdVwzFsgv21dboESHX5+W0scBTrN4nEbOW5zFF9aOEMPVFjTbt9qBcoKrpfqu
OsjVYqlV45RuiLGHeDoFK17ycOTipFR7C7pqvghZnYUvD/w+cTxVtRJU5cOmBXr1
F+JoSc6NOQ6sqLBhiXpoTqMbLVdowzWkmEFqSxSoQzi5Muo9SdnuO7Ubk9XGOcjF
ckxSbLQm9pZBTWzw2VLpRe3sBpbXBgZeLOEZISgHhbGh6ejXhrjpFc5BjNd0Mt+d
XUDjT/xl/68p4L5zw9yUoJd9D+wWPQAFXyfas0DMUhQQf5U4XKSdF68X2BMQbW2o
TfpbqEJowegoOFfZF4SSHIEwvicJBSVcpTRGrvjA4KmH0Mz8sAvHVbx+QtduX/vS
tzmbQwyWVq7J3swJ6qNYAUn18SNuUkEu6JXs+ze2MIsSDMgwljJeQTfI2rxq7KrY
yBfvpqxric2GC83ZD04Ihpc7qusX8YTkvapZGDm6NOVhwbzEFBcmekaInYTI+1Vm
bCo22JTbeZi5RDYgYq6MWzfYBgws0O6JrnoGUkg66aCOWlemPLZI7lpKmnlh8twk
HI8Vi/gNGszXKnsdu/xuVnWBH0E0KouYdKP0F/4LvucyfVOJbmFcVhtUtOloqvxA
Yd/BMPwHVpT1S20SwLpDo4p7I62LzTN17Awb7fwHnqrDP/6l9LFkRGK8gukbe9es
bdDiuwZ86UP+29z5/O4uDfFnOiOzOlQxtFdrqI0XwEiGfHH2AvzoKjp8TqDxw8uH
`protect END_PROTECTED
