`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L09VcnCIl/iG6ZXY1CLzmlcqxQa4jWU0udgjQ0YiZ14D/wtnluHCAlRkWSHVrH7G
BPE1DFra26mS4h3yeEJMUNni2b+FxrbvFpGHTX1ksh7JKMRe0j+kBVTORK1YjyEu
MFcif9HQjm2+0+Hpx2TDmTxCeUsJ0rg4v7Kq+7HJKboCBRJNE03Tcw8x+VWHWT45
R8FKAmu8224wR4jlQEcPrB+LmQV4YM1W1nYBubZYiEgAM1gd0MnAFavN/LNqXW23
L46gZ+7eCUqEUu/aqX4ulogVlA63/s237999DG4C+PNVRnIsfl+J6ALCk4DmdMg5
3g1b3UYj4aAvXIam6eqaCdXybcNI6K75WXO5VWiEPPFS2qCAf0OEAU0WpxkgiWAV
6UslQQf2KEa0HpFBBfFxIB8EsiL864f9t+5/gSmnR4PWoQhKKCPZyRktM8/YHnnx
0UR6zI0lASzNIKIE9o4khFxGTki8Vuk4jLeefAk0GiAG7h+RKoYGfzxa4M0h8f8s
x+NHReOBGTAVCnbkLc60/UvRWxWM3IOjoTXfJXF3GodpQbuBKsjCh+YvSKZY+itU
SoMyF42DeK67QQJV2jl6GJjGo0prAA0f7pHQU/YjKfEYUa+GY/iew57eJXsbmh0K
XozLLQLCf2/NBuGQZSRXy4saGHYqX6/UeMqksu9fAd9M2LDdVtIqwRIC8BLLO8tX
O6HkK2pTrm1Ii1nzCT3RekV+gZblOu1HfmQWQ4y8Vwm5UfIFODNaeASc6E2CHrZy
ZOnDr+bJClzXyA+6A7xw7LS9kjdBBVt0aMezmpAOBeYPOiA1jdZM1D8dOIZ8Z3PL
KeEZl581ZKGIHwhzfTbCxRvRIbuxiGdjbQg680HjrCNmE/QidbjlDTcfkhqWRmld
6vuoGfZ4jXvGO+GwjyGJzUykRg23YXg3RY3POoPaUZy/wrE4Fe8mXf3x8rNuIbal
ienas04+QPwLKlIe/4SpwD5UqRYQXwlqPSuQCyrkK12sWJ+8u5DG464GciIwFnPQ
9sKrJub9l0HeHVzpLPHtVw/3rD9BN72pF5sW+zHN+poJY8eIxdau9bLfs58CvS/Y
aZDyAXykVbyiXw2YeTg44rawPr8wwle/rsB9cy0sYzLaF1gBrwmx4h/3AE7Y/7Cl
g0Qnd1dJ2XTXjgrBKdOoDpuwKK/h0U8BESDr7kzhs1+U3i+DpRFLzv25AQuC36jc
ntVneFBMBUCRCInEAzHuDzvRJngny9xe/FKpBfBDr2C8ESxbb80WvIygG81M2OxJ
wjPQnQiyJZwF+g/rZWhKmgZKJlsnI0PDO7YLV8ObGE1i3DRGufw46qXUyRDGfjPg
iSO09qYbLp8Vd48O2EzYEqvmdfcSQgAeJguVt0yPHy17wH2GPpfpEC+taC2EwE1i
BMET7xZs0hr8HMWofzyRuKCpyLQ9X0ziWn9XJBs5N6dzBHcTGcbtRGIvfyOYNfay
HDAMmzG7QDS7qWwqKOOr5/rMq84jVlwEI64DtsMaJqxg9OW1KHunyFu43UUNaS2y
3y+KsHl5Ha05xb33+z7/SXdGgCNUGVJW77A1zYYilwi7ndWouZlr552o/YMy7TOp
vUQnNIIjsnjhS8Xb7U1xDtLo8zHnmI7qte1jJRJmGKnkePNs0HrvoRordYvf/xm/
zSPkABQAf7vJkLtdoM3h0bji1OC25J+ARERqdtzZ6OQdMDmIVTHZ1dVhPnMTVoav
n/UcdafHADJ87a/zFgsF9kdjg/3NUxETOrkNMHMuHuqvEFxF8wrbKyy5TTW8b+ZN
reAp9xO+iYNd1Ym90u06sCJ/kNvUFeK46Jwiqr5cE/sG8X1TX4rZ1ZiQQjpVzjWG
zvZMlswkUCieo1/ShXF634xVxD9cnla2Ihhq7c7FJkFuv5NLrYG8ZfIqWbijRRkN
N/7NimKJXZsR5Qly1GqBuqR+L5QTPAPhWbzRosZESU2ebwoqTKpbBuqXNlRc/Ez0
9XagYO7klGs6rjE6Xspp7awNTQc6ag1SpKLFqmR1kQ+dAHbPAhOcvruCNArbEBBF
KWkX48/m3l9sv7k8pD9DKh7il8QhXpU1zHCD9J5Jefqu/XI83iIO+m9hfhauAw2H
ZsdFFyUMSzlsd+fpsKomOtqKDGS7B1Ow+pAml0i3ygiVdYNQMH8T964dQHyrdBzU
5bshNEMmoEUUn64HdOH8dpq+mrVZNfrV/vJzlmP1qZp5jI5zoYJc7XXxGok7YijM
KOzfjL6ZahLqYqnbVFHcRV6ghZX70LHF2rowmqBLZ5Vff5FlJMSEbxgufs9qgSvt
BKlWYY/tb91KuSWldvRxrtqLERQyFkxzn67F8xdMMhSzEdr2XQR0BBk6AHkrmcDf
9SZQX+mp1p/yX6zzrKrKFsuZw8AIGtPrtOzbn4Lp49fR0MjYL/XRiHJedsb2VtZX
HaamUtxJ9BTQ1FwmpysyZ61p0ZNFMfdNuuNAguiXrbPeiBtjjwpHp7QCGqle3Wsv
Kdw59OSch4SKOsDU/XyvULbo+yuR3BN8aBcqcVaNtSHbQRMLhiBpNWAoGuLjstZP
KvVJx6SxMiw5AOAWLHIJaPq2uS56wcoP2n4JwtVgHvlnbrGFbXp9nb3If0IusX/S
qhrd4GdvLWYYK8QP3W+QLXOvUAtKZL+qWWo6lIPlikAfnQ72S3rHa1yaT77sBcIf
4Apdm2OGh1zosxfeoANs47f+MW7aqYSgJ0Q+qAFW7Y+RdULySPq7mTHAsybz4ps5
HuBjEPPEqt7eu1kYYA55Vx0fOMZ/Y/KYt8aRFR+BFeq6NTxLMCoDZFBPX47XPVFV
rcJ47bZ8qz9yL3HUHyD64ghhVvJjO5ZXinZVF+30hJ+9PgrRdNY5DjWoDzsrcPok
2ZRrp1NWmxEmzvjnjNIM7A==
`protect END_PROTECTED
