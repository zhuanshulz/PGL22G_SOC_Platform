`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n3S9zAGgIq6dkzwBtakbCulTNbm3KDTo+HWWI6CYB95K7Nn0rZxZLlCSrfbhKazZ
SpN16Z3UG29V4F88PLQF0dcuQv6XW5a7hzkNczKERwkCcUNuEhWGbyEoNw6CoDtr
7Gg0DXQSOhChnbYgu/7JP1rkp/ZxqbH0UXAyPRBbhzi9kHHwOB9Sl731uM3RdSHV
cADWI2dpcBDKWBzJP0x1+zDQfOY+37e48xlG1TGaSYoVBecdD/7811n2+eRLXnP4
R32q1mCN9yuQtNbsjAh5CQ==
`protect END_PROTECTED
