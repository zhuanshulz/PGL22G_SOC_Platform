`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FGl57UtdH+plRDcJAapdwDQf67KmbfDLgwCaNkoZ4kx6ImbOuenKtlyRbVq3NgV3
HFk6nR9rLdSlg79psxytyeZwVdoLSmAW8IsLIGNH+DnnzTS1lxETKpQ3IpiT1/H4
4KnB2kEtMt2gD7hPCRDp6FBOIU3rZFEjoajWah6vpP82c9NZpGZ1Ryieo9//JQaZ
QrF1Rl6ze5I7HgGcbsVUZZDesxCg7/RAVFYH7iALmS3RxhR6VwoySvyEffxA3t3x
mizqwbbflTnzIF2AaOjBU+iOb4gfz3hCzE4zX5quLrCjkkUffdzsDD0yF229iPbg
zUeATSNxnM/sq+BokIJ0bxFWVBS7YS6UYdkA3QaWNdGxzbVLyw9+hvMXZOXz+5LD
35DJT/Abo7iwEBTLQn/uvDewExRC48pN8JYnogS/6VohBgOjaJW4ebgXHsXns117
SETCNnJGADKpdxHATUXom/4aM8+IXIszQD6dRg5XQlP7n4ohTPeJ2qrSGpJOKnRm
G9LEupAaRMdRi3w/n9hscsLibJZWC2ucpxeRAliMa4/zPOoZpC7SXhi2tf0uAVAK
`protect END_PROTECTED
