`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+5p1gUatpjmTjKEebH+9gywgyX6z+3UQsPhMpo+yDuIAgrWrQpOopYlR946mWl3A
mpV9dq7BfXNZ2SdCik+ODrgMG2dUoHcLJcC5gQgttv19IwZMI63FRnqv1/SRVo8A
isuGMl4Jge4CglmSGaVYG+b3vLs0HjmSainIhOncUOcT0k84o15LAxcJlhwpq3qc
99mZVMl80d7VZB6Va74FLVRB7Hu7l9o3aU+WbpB68dl7kOjSip16qDsH4mDNB18D
AoiVqU57gj5aZJVnvvV+U1Vy08pKTld4KvcACeWkvgp/s4HcOk9wIoflx/Z7Xck7
rVfnjP0iMObZAlUUKBnyD/DrkwOAR6fCPLlyf7x45f8KtxKHiwia+PIANIiPO32M
36FLosdZAda/+6vB05Rs9GlXhtL/2DJk7b+PYEEWa28ydhTfOXu8Y/kwf6nwFHvZ
4tomGEKjBGPHPz9M+UbJrShgpQRIdycDWBFUkC+q7ITQ2krV/v9EXaWaE+uDz3Mp
4tQOQSn4JvhPPeK4eJQYDQ==
`protect END_PROTECTED
