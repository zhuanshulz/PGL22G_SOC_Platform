`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HGBh5cgKw4NF4Vmb9Gm5Ew4axHEVmJtZb2GdZLfDtP9qU59T+9gMyP0Lt6oiKWDP
2yCI5pPbLSWfhRfrLrrUfhNPHLYgOTrg7JG+S69SfQz7dCQyd4feP6BDcclry1Es
5C2uhLsAlfzHrVquj2YWnsAUqn3Qxzp3BnLFmVo47LOFj+AnHQLZ9+J0apmYhCmW
Uf8I5w2OHy0pS0orlOa6I4cUSklBqiGv3AbOh6TDERsCGZvrg6r5pNVePx+PMTPE
BOXhSgktd7Y6PJyVkvtLNhQo3vSumOmgMzZbnJ3eI3LwET8pLS2O9eD7LYn0iC8L
iytDoqlBL9AN5WHpOjFjoi7T1lUw8R43A1eGmOsuZUfJ/f3bv9n+lcoFYrlVXOSO
blDiJSByT6UjcCOdh7+s5Jn4VHGFAR8TNsIafevJ8oeDzzsuZ7W+rXX2qZnf+9AG
`protect END_PROTECTED
