`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zOLuCg8QTKKxN4qEnKPmE5ANW/eV/7Rz91+W9apeMVBNuYBeVo1fizMvbbMABBV+
Da1Upafh/e167RRrsylPe35S8IZN5PftT19+pGRvX0MimdvgA+UR+GEgyJx69Xfb
r0++fI6KoXIsIGpS/lzUlnN7EKBFY6MoYpX56JO6pf4mqLo2HTZcRq/XfmBbuYcf
+BZmIMWOQD5/ujuJjytFsWYUUELdK6jfqOWfRbOSBo3ZUgQww/B7vqektdGyNgIQ
nw6caf9E46ZXkwyYEjTY0srxQi/KhWjBnuS8e/r0XCil2u8d8JIMBhKQvn3v1yc1
7vE8uMvUlZ8bowsYdm5VyiEyykgSfYOPTb8jTsw7ao55sRGLFsNW7wTqGYIYfs8t
O6gWDJ59ooO0QISNggNH9pQFEp0IeiLqx7yABgcmEqb5frwVS6S3eFhm3443vpAQ
KOtExyjsJnNNWjW2qzheSjEHUCeH7LqGYHsAsnRIeq65kAMTKHjMQShG45paXUEY
kuOavSAoiYHGVJawO0Yo7FsxdMfqxpnkx0KJ6H2kHvunAewCP6FTS/+NfkBVVZzM
MO+SsO4ATRLUONX9Jk0JoQ==
`protect END_PROTECTED
