`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jYxuEWwIgcknBz3/raZutuxvPEDnioqwuX8NPq4Vrj4o28//v11jpVsqhqHpOA7e
16WelSsGuHsOs8JFOmgPZH5G1J5lR2hXParPflzon4SCCjzPnHqmsYB3afTA2CAW
kSlbjH4Ue4VGUX5muR8FZcQ/giJWlw3JuPvbDRRHnsl9GW/Y2gZBrFG/DFuJKVA7
IDNcaghG3Q6BSHTF070RmoK606sPBQ69xU/3u5zdLY4paAx+ka7XlCudMX7W0eYB
sCQTawdfe8jpIDI7HBoZ+NwQib+kF0+RW1C7h4WjGOjvyqyt1mLJozfhQMAPrIpI
0dBncQw3PuTjVVLbSN5ttLvVJ5AetVWPxw4Ae3G8anNa72GHjcYhBEzKSfUj/LIB
H8U1BHmu/zKQC8PTTKn+xw==
`protect END_PROTECTED
