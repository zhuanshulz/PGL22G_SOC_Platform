`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zmNUNUaIHxl58feLpEH30ntsog6mzJbHHQybsFdMzmo31bR7bDs8XzwGkIHlNUmh
pEcwzTvjMYDnG/K3uiC0Ht88Gc/kf3Cd3mOIpgaQUo65OjxRnc2zFUBNIaZPAPXk
KNsRCKpvafc4MKgkaOyfhfxDe46Xa2Yep9h4aS5rM5LeKp1cXwhj388yqjPpxIZ7
5YJUZ9MHj1evWUtcVADThRc9Heght73WNYKdVJdUEWcHFsUq7bpV0Y7fvDueUgjB
zP0uIlio/o2LOJZatOi6ICZHZvGvfU6lCYxENKaqgsSVjr8APye6Y1r9iwoOcJmT
nFKnjwN/jBPU9W92F2pY963EgA3wye5bSHJmEDmDyu6hiIO9+fax7we41RSlR2lj
eCRWvZ0oUjfr2COaWu09Ag6D0g1MfLw+8QlVflFAkJoPFn1MbZN/dPvSI1/jjo1z
jTl/2NAZTxeHAVtkZ4RNiLhS9FbpliJXF+6+uaGlbwl5LgoIP51CEjMirEAgHowu
dCU3clIiCdZG0iJqmeaE8nCUjtgYVAARS7e49SRwlQ72zE8tw77+jd8A39Pafi3b
kvCXQltb/5usy63dBgC+8g==
`protect END_PROTECTED
