library verilog;
use verilog.vl_types.all;
entity V_APM_MULT_TEMPLATE is
    generic(
        GRS_EN          : string  := "TRUE";
        SYNC_RST        : string  := "FALSE";
        INREG_EN        : string  := "FALSE";
        PREREG_EN       : string  := "FALSE";
        MULTREG_EN      : string  := "FALSE";
        POSTREG_EN      : string  := "FALSE";
        USED_PREADD     : string  := "FALSE";
        USED_POSTADD    : string  := "FALSE";
        USED_ACC        : string  := "FALSE";
        POSTADD_INPUT_ORDER: string  := "CPI_MULT";
        A_SIZE          : integer := 9;
        B_SIZE          : integer := 9;
        C_SIZE          : integer := 8;
        P_SIZE          : integer := 32;
        DYN_INIT_EN     : string  := "FALSE";
        SINIT_VALUE     : vl_logic_vector;
        OVERFLOW_MASK   : vl_logic_vector;
        PATTERN         : vl_logic_vector;
        MASKPAT         : vl_logic_vector
    );
    port(
        CLK             : in     vl_logic;
        CE              : in     vl_logic;
        RST             : in     vl_logic;
        A_SIGNED        : in     vl_logic;
        B_SIGNED        : in     vl_logic;
        C_SIGNED        : in     vl_logic;
        A               : in     vl_logic_vector;
        B               : in     vl_logic_vector;
        C               : in     vl_logic_vector;
        P               : out    vl_logic_vector;
        PRE_ADDSUB      : in     vl_logic;
        POST_ADDSUB     : in     vl_logic;
        CPI_SIGNED      : in     vl_logic;
        CPO_SIGNED      : out    vl_logic;
        CPI             : in     vl_logic_vector;
        CPO             : out    vl_logic_vector;
        RELOAD          : in     vl_logic;
        ACC_ADDSUB      : in     vl_logic;
        DINIT_VALUE     : in     vl_logic_vector;
        OVER            : out    vl_logic;
        UNDER           : out    vl_logic;
        EQZ             : out    vl_logic;
        EQZM            : out    vl_logic;
        EQOM            : out    vl_logic;
        EQPAT           : out    vl_logic;
        EQPATN          : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of GRS_EN : constant is 1;
    attribute mti_svvh_generic_type of SYNC_RST : constant is 1;
    attribute mti_svvh_generic_type of INREG_EN : constant is 1;
    attribute mti_svvh_generic_type of PREREG_EN : constant is 1;
    attribute mti_svvh_generic_type of MULTREG_EN : constant is 1;
    attribute mti_svvh_generic_type of POSTREG_EN : constant is 1;
    attribute mti_svvh_generic_type of USED_PREADD : constant is 1;
    attribute mti_svvh_generic_type of USED_POSTADD : constant is 1;
    attribute mti_svvh_generic_type of USED_ACC : constant is 1;
    attribute mti_svvh_generic_type of POSTADD_INPUT_ORDER : constant is 1;
    attribute mti_svvh_generic_type of A_SIZE : constant is 2;
    attribute mti_svvh_generic_type of B_SIZE : constant is 2;
    attribute mti_svvh_generic_type of C_SIZE : constant is 2;
    attribute mti_svvh_generic_type of P_SIZE : constant is 2;
    attribute mti_svvh_generic_type of DYN_INIT_EN : constant is 1;
    attribute mti_svvh_generic_type of SINIT_VALUE : constant is 4;
    attribute mti_svvh_generic_type of OVERFLOW_MASK : constant is 4;
    attribute mti_svvh_generic_type of PATTERN : constant is 4;
    attribute mti_svvh_generic_type of MASKPAT : constant is 4;
end V_APM_MULT_TEMPLATE;
