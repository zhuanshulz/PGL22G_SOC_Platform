`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2DRI6kLyqHOCaUa07KcwQ0wBAEHhgNvjMFu+3IXaYgxsOvpuQxtOXJy9E7H5RcTQ
FJUmN34O0Od0t3dcpb+HnxT60Q+LU5WHs9mIOGPqR8z0I2CPS7UhziuEsX4HUoJe
xZTWTGyYLptVEiipRy7oAS1B8iQqNtpBniqBmKIU7+IxcH0gCYbc5TS2KIja4xAl
5i+qogHomeCFuN/JD7BZ4elrCGWJgp3GH54v1Ca3cuDZR1B4Gd4jgBzeWgqHzBat
fS2bmmk485w0Z5DpX5DVQ6n8+nbP8oWrIL5uH/RNvu3NrfuMdULHGYvnumbB78fm
/j059LLrmEwRQeyw+b4WrRH2GmxvMMfSpGYDrNXQ8QJSYk4vS5DkIp0FldPP3Cqo
tnXljUjsO1EpYDb04JNv+YBWmlSTgk29Bbd7SdYwwxK60Ydw0JLV9nP2mwSl+Y8s
M1zy64z5HjnS+VHzQBBFH384mOxrdEFGc7d8yIXa7wi4SHFxLi6R7izBXhiz5+ml
hfRNi7fmJU4gr028KdMQkPTml1HNM66RzeYq/tzMlECHMVta35gOIADQx0mSUHMi
JI3rt1z5NfWd3jEgRmbbDaTreNCa97qNPsHtGWS4NQ27j1ae8MyJ/aeOjMsVZqze
5swkOZd6pMO03+BJYmYcV5X1Xcpm2syVb9+Gx/aMAX4ich6LVvOurXEnDIukprUa
34qWxPZcruGBY9d5inMijAgj+fDbXk5LmjcGJMoO6sIvFQfcNCCpUh7YeWmXVGeK
KX48SMN7Y8DrClNUOs97WFlEP4pQGpdi/igSFI1WaQ4LwVxmje78byqHBIt3ErRh
FNigk1LwBdRxlur7f7h2GWK/EoiShOBaszsUvvQVhBIW+GEsuQCCUtULW7ZJYR+O
yibs5QMP/VhiauZXjSPwjr+A/08UgMSD2ZfmTsr2+jKkrEeZHjqKdt8enRGQo9/J
f3WP7yWJH2YAOiRgjQpI5xlQ3Qbl3JzpN3V7QigWKIIypDQz10LnvABf6CrgnDPS
ELTZEZoEILhVC+dGPWOPerxF4USDt4zlPgX56fwWOGJnFjrFfjJV2YN/W+ODQcAR
uO4weEAdhjW/ZDoWgmBvApQS3UQOlaGXfcN5Zx50SCMpJYoSc6aCAS5KI6eU2FZj
fIkHbv4rNzJqTsE+bWsHNWJUq5JTMBs7xTJnIbKY5qEKJ/3y3q8WKDSheMl9TYXr
BVJZq0GrzP7XL4qmdVsmtAr8dyFaSL7zEZfy9YWl7MBFy8jOmh+Z+xvk8KFTuG1q
9ekvOxj1jpCpELDX8z4G4RUHWa8ysNbduUioxdLjemRzAfuMhC7ByjELz51jWC9v
E9T8LXZx6IrkWwdM+4MSpsuHFoPpPXD3vDfgE7j4H89q8iXPG2Eb+tTeaWP7geln
ywZI1HmYu53ZaI1LeWH/9qSYGld6Qp6+0AAptMftASo2KCK440TcnBFfo9rasn/l
HKxGPc9GuOKuMHVN+1PxSkuPbGKtffJPlp7aiCxcLBAFURJFWu71y7uv6f02G59L
x+wXO7Q9uznVUMRCchE2iF64eNvD13qNTNU9AdUGAOjVpz36GT7A1NmW3cFxHa2s
6Czo2szUJhte31wD6xRUryfSUEeGZDaI1v8hWEM/RpTc8Hf4hjkA6pnTTPkX/RM7
8TOjjQr6UP9lncrXhTkGeuFGsJigsst9bAsqBbjwDGv4Hfk5QShlYts79xybR944
+9UboxI3CVD6X78wNRbpHRz8f5TlXtwlr4EQrdarpKGb3n35MNZIflEoSIde+ZHL
UAaWFjSaWZg0lzSff0zqYtSlYLA5hkYRRhCYylNcDqnODlpme9QWw/81f1U6Nuck
OmENBsi/abiVlQSqNcZAtP6dYEyi7BAkptLK9WoJzlspNWsQ1okyW8usIDSQHXwO
uVGPvA8mHqzTep/3ZPDMwOUMJ14AuzSPn3RRFE2OcHtJ6UKdRj7YrGl060x4V2EI
CT2mp4e0lByOmIYDSiMdB1/arIt7pdAhmHeBGWFWCM3zJMibG7qa7QT7Og+ER8je
NaHpYdgxz2m1HyCnQ/k+dc88sXAz3v3g7F5Jj+UwS1OLZ5aNqLFV7pfI/U/U3G0l
xpOUM0NCIbZx76M5SnQOyKfVLSlLfrbY2UD14PHdHEnHpG2HdaXoKzz/GaVZZhzQ
0rQjHNXZKW/A2mZkxIWasTAK3VWwztcxis0V0nMIac22BkNaDfD2vmd7M4Jm+Buw
Z6lR0lDoeWxVz93s/8wvSFedBYshpvFrv54/iFbcamJ2OPDp1MyvRRq/e7J/8EUY
WU4MU4heG91m8Fd9xEcI5B3JRMYSYO6TqJw7A4KaPMYBrR+/3UudE1w/9htkrJzt
px1OHQdngOEr0WzK6cI4t6xfX8S6NhSHA3VdGBKUf29JP/p9LYSl+1z2Wh+RAFWP
6BMLWKBV0PD9Z9Yv1gGtxiv+1xzpYOnj4vaA9vb0wH0IB4Ef+rPok4aR4gj1E1dv
leEYF5GL670UMI2ztFHAa4jAEt4gWfff/SwMZBH9cZ8zI0JfSsBQL8Cnyt+7FGlz
dyDRDKdXVGViRJFUewr60EHQ5KzBO3edamfZd6cNnFjvcnL4VIj9GjA+Yf90HHqf
9f+/caeHJhgXDtn+9IhPefePcvaPwWV/X0SGwMbKAz4LlczIUZPhVcyRgaZIPG3O
Bi59LylZhcGbv+KzSecS7ZHH29T7mZjCdeWksqDQ+knmcZNxPLIsynPJyAlQGYQy
KNVJXE8sODj0zTwp2ysVD/mEG+zwHOYYVIDXoYOrEkc=
`protect END_PROTECTED
