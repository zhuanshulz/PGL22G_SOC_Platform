`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4tdfainqJYgf9qnioJGXTTPCcLRLUPKh2J7jkUsbtVXuhjGbkCPmbTlzCnekHttp
9m3zydw1SbOsLwe5myweOgRxpAZ5OuBurtWXu7hUNYY5TLNHt+e+H3fc78hRWL6z
IBzdSrhKP1bUIkKdPRduYiOyQJw38HdbbqfNwKiMlnADq6JqYnj+o7H913gihPvw
0Utn8MDd8zrIA59tGHwLPUriRNF4ZvTxQaks4GfaGlIrRlEbqhKW4zW2aWwK7K/n
hTXaYBEucgJN38tZsKYRdRUlh/uAKltceu24AENBSrsDVCPCtzwYLcKS5eRvBaVV
STykOGOa8/25qO+w86tI/5mQrkO6+7wpJcif+KE3IQcOTlv6KQ5/CNz++8Uy4FDB
EmursKTJHadcncyFcipXE0xsmBXD7kc5D1apm+0IIen52NKeckNQgKshUQ2mqS8U
J1lIE9LKhNgtfwoYF6ukc5d6kX6eh0JuH1ztegv32VW73zIUkgvam6ZNqLimlZur
RehzkTr+fECT7cr8UKXz8LBN9EU0W0RbQt5IfnxAG5VsZBUdCmNY2Hgt2HYdsK/M
cnVPcIDFu4nKKdmNZvlNcoGXRWbQTNfe9VofhLK8NXof/zgKFGxQ3vGagT1NNq9X
uymacfacn8w/e+oERxeZhnc3Yebkm3QbGaor5cJCNG26t5NQxNNFi2TlP3dTLit+
LhljP5fgs2PD9TZzcxanHzlbtKUtnG3o47mTCyLyxzh+tGLBriVz0rTniddjypQ9
sdRjQe993Hqw+AYkaZGIZxi5HigblReAz8Lc1q5+5nSu6QccMPMN97IJBHWjHGmj
NSR8Au/pta+Fz5SLrHfEEpcLeWcETNUcDaI2EudHLRr6LUXFTZ4yJEgIWaQ63Q3o
i01fsjN2c3wKfKsCQvIJNFnM+QjXCoPHucMsX4xCcSkYckgxwtxRkkDMXUqqAvRa
HnRASA8JH4yc0t9pcIlyxmSkZCMd8acqKCO2AjmISZzFgVaH5duXR3I5HbVymvyr
/0LwqHkYypyGAHE+HEaDnPKqiBALoTWa010S1pOqL/dhWp12qwegGj494MFSL1wt
bqAKNIBNzWYk0IGkfgeiEzznwLf0BhOCgaelkxhSJe7ol7GoucEdEQ68AF1P9mFU
HW1DbYmbq1rQyC9d3mnbVdZhxOQ11wJnC2imYH2OGRcYScytJIMm73cFBkr38tz3
Q7CJix7kwhg1jTQgNAstL/wLHFPkRyILpbRRZ527jABBXOvpnVNjGJ6odACvdLj3
8RO68etY0C5+lQK0oiVAG9wbbnirmCl7NFYZnnahje+nPu90vsvFe7H1NBcGLH/j
1I5scmb9MXN+aR3TDUA8EO+Eh/NsD3JhaP0uQ28lwK99JH18qNlupvbYqnjXrlAY
04fGReRl0AwA6SBk7G7OdQxNx+W/oXi2iBjq7PztMGdRP5EyPTO6dsthdXpVnutO
46fqfXEyUUriX6ybJ+d4IgA6k9iArbJtUehFlnrXIhtrjUWd2uFVvEub9DrqQd3I
AthdKzfJf6c1N9OLb8GuVbPZh/ruWw8+LL5nG7JogdjnzpsKIbYIy20sHQ94vGXc
aTk/vH0a2vtGmdMx973de/6NPGO9LZfKqF7LPucVp64aEg0NITOamFGbeUx6Mixc
bjaBhKDseFO+56gJ4xVGUtdeKQDDBJrzu9FL3dlc4Ei7WDw7WOs7IHh7lRNmv6mL
0pxwM1eN2QqkRF3E+btE7Db7Du7S8hU+x5DMV9YbtgXJEokTKSTqrZbw5IygGi4L
X3sLMpzSP/ghRnqHyXe1d7NnCGhnqOfJd1WUKoTk8rE+0kUxb4AQ8cYbl9hHoNEu
ikSd60eDyhqZqcSLUwOpG7zC5RGg27mqHowMgt4t/kbnrd7YwgAJ6o51/BvFkazD
B5Yivx+OD/9+52SokS/zCfGvygQ6FmZtvkPrmG7GUbdgJsn2xuWY7yjYMUN3p8Aj
rB357/rO/HYrMJOmS/Jb9yEKijxMu7ubrKSdHk7VeJz2fP4Yi/+m44e+cClk9/pk
H3u4WK5txecPHFoslUYwYNZAcVi0K0ow12rPSZ9c/YHFiQBWKiu6sUqs0sogQyX7
SQMxHiu1LT2rPkb1lxoxaUxa7G+JchQp8cR/ME6i4lekqVPdWm+YbaY+aRPgjrGJ
vgV9Nju4nwctDu7Io84esEpZwLg21xOVsuuRQ0igJiekEp3+7ZU8HQCOgZkGBZ55
m0Hz6VepjdD+mCI1sv33FE1Z4uVEiGLnI9FF4dPuOYqrLzf3RX43e/VX/qZcrMIN
W4HeGVKu3XRnqzu8xtMkiQ==
`protect END_PROTECTED
