`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0iioBZLIEjUr+8lSlvmhNnumGHLJq8NCedyvZsM2j7jhbHY4IzBNZrEC4RJT7Rij
TUbu6DbGLPOOwhapxKXFnwfHL+47DAwiUdQyEBvnupqn/N6RpbdCkfAamSAoGZ1Y
ChVaK2YarCpUdNWqIrZ+jgthZrlMZA3y8Wfjth339zmnXb4dBn4YI3IBNZ/Nm7zu
hsVbe9mMa3jFij7VcfpQ1I5Ce4co34qBPxysa9gFFn3b/PMopiC63CrETLzRun3Z
/LeQMc1f8ZDgMcOIqIjuu3ws3hzriLpJOGP2XT8i2ZhwNzqQSJrjx/jOfcIHqYPM
8g9pL+23mRf0aKXs3JqLg1B2AfQqeAp8IVSYjrqF7N1ClIwu2tiN1x97j5lLQeEU
bSNUNaFgLsisre+hL0ScLyc0kjEyi3CH/brI0LqYe4eohN6T/dajxE1bDkVCRmIX
WBj5PNVCZEOKUP6nAo0Jbc1lmF18vA2abR898X3BWnVSLlRSEu/scsIQj5JkyhcF
whyo9wj5FPZrgqXN4ZhbyeV18I7IYVyNzfl0L8mGQIy+M6Mr2bTAUrv/kDHACw19
/5LSK68qj9wzxKvMnasC54F4UqO84jR4nrsKgLulWfrVsYvZGDd7QSMmd3OvkMpe
`protect END_PROTECTED
