`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bYo3YOciVMAUMTa/wbatzwIKUiyMlyfCfwazd+XZIgEAdyRv5YTP1WLAiiAmn9w/
H2lSFK1RuQJyBKJL46v/oRFh+yaXsOM7NrKe6UNkBYgw5VfKUMHYbcGBgy+G5xJY
J7AomxtjQ03GcMhfGmZT/tApQcTlICo/ZIZhnGGIDXwgOwB7k4occYHhPiYT79Fw
wu/K0sFAI6dZUJuCSXoIDg/LFV6Lc/9E1hIwZuKri/kcMbZ9d2EWaqG9R/lUNMpn
AZjn9Bc1ia0a9pkcWnYmWofRa+p196afSg+asE1LR2Zasb/Yp39II31CYYC7xMWB
HHdMBesWukIhvr1le0hf8RrSb9IM4uPB+/Fu38dnkFSWHIrAJUe0dkOBx/q0uyG+
Moy3dWxUym6OieIXUsUx+6nAp2SSeA2bJ6Z2Ri+/bNMnzdaKVPn8gt3f0qoyC6CZ
MZiG+egoVMBSzReLEZ3Jf353VtIgjcAZFPl+f44Sr4oUrOF0detcqfr9w/Vmkd3r
hAWS+jprjAUGjnPl0qDg5NvzcXTWhoxysRCmRDPec9P4tXNjJ+vINIgr/p7qfXuB
rjkyfDa6Y38oDjHSg76k+7ZVp5DqW8DDKVjEbqCXHJ5FJAQ5WHxYmmQ5eIQk0fS7
glqxbtJFmSI4nxfxRYy5COPYs2j1B6WXspiFhNikB6X/0GF6LJULTuIfjrfhJHLu
ujFUX8BNlB5o1n2chh8fK8lKubctmcNoLmqEFwPtNIuaMDjzKqywKy3m0N0dYET+
hpDtGDaZYlE9n/Gad1AZHT5FH2e0ZIjxPs//KUweZxIne6z/vFYFLfOO6sh27gMq
0gSODX3kYBNDpnyIY7oIrMstlqY1M0V/fXW6hGXBVv6/p2f6paC4iPMeuqwH4BKr
NkorKMD6Y/AmFWKRP7VnNkvhfvwEljClywGhrS91oEXbNFprA1CkcqGlQ5C3weah
`protect END_PROTECTED
