`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5EFgzgKcUKcPCpLECx0r67caGamoqZT7nhrl9Fg59hniKb5OM0hgmlHDyIvfts4K
1Mwr5pzApTwhw1aXxoedMFZfcD882F6mB9aX+/I6+U7RjsFu7ZO/b0aSCcWE01Po
g/Q7T3tIPHsupYRsofrwKCt2Wxs3iEHO84Lk/90gGmSDtsAhNamRjTP7YtTEqdVt
9G18d1OyTm5zjvGX9qdv/nvyCZgJs3ICfxibwKENRoiz7qd+XpyvJ5HXA+6nE1KX
O+knqN+gU0X3MW6Fu4WsHRIXPxrWZa7InL/ce0hfWcmYCl6QuEFg/TDWJoSnbsES
lZhWr2VQ0NVCOMSsFO/rHtDMfupmqT7WfO0CmDEva0VMlrIBUSnP87aGVnwcSqpk
amyw98o0EulObdBeC9myAJGY8ArcHadZMSQ5INP1Z30Zq+D2f8OLjSBAMaLZkAJd
nVp7pd579g7MLko83Trwp/aRhxXq1Lj0ey7YInrJVCGBSZqx1Zfc/iyOAEva2MBe
NyRFL7MJ6RpoxLEIEb9f7g/S1GFPQstS3KAhq1sVdAADnoD15SETRXZ/LiBFUVkO
LJ06GypJ463LdEkfmtsr8H4HDGNef2lZ7oZ2nbRXxT4gx7Wu1DeV8xd5pZziLkW9
H4W3IH5Vg2AWRNTWgUKe9Fk066F7dlPdTg/uVP2S2YV909gBnWKVW22DS570DRtX
kLNBu7lLEkyw+mR9Y21TNc2QS8SfVSAF6OeEieVXGNVLql1TA1LN19/Vbrepfjp7
Mz6HMefFShx6bvZr26iBVZoJP0+764GJZuxR7s9moFXuYJo9PMPP3kbJvQX/+Cpv
`protect END_PROTECTED
