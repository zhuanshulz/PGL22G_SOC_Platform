`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pA0wW3EbRejJ9MjutpQ2ff/dill7a6SxI0jFKc0b75dgRXEwI5Yj6575ptWGB1FZ
qGjhtWMLFAD9ELbKu7mhZix0xF+QbvcwJsV4XY5mSR69kB/q3kifo3lnr/sZ1+j7
HjdcPZQALo9NnWEYQbqLLuyOcti6TMgTjGVG+BYNaBmed/VRGcWCKBwHUhDqunPH
9qHXZ+UhT/O/cqE4ZeFJqDeUyrfZKkcZmkjaEJBUd5WS03qTzRcKl5K/381jgKHj
VyPeuVb7yZ0NoHp30MC9haCE8Qye3TEYC7g2yaN0EL53msWlzeRsycuzeT6V9sqg
ZmlPojl4FTp3Z6wp0wJCEYaw+ZRtHHqIA5zXZkX0+Z7iGmbuP4RnKBuK6TPEVBK7
Xdo9/zFpJHU+dnXcVwvb0EfvoOlNL6AfsFInZvs7QdE=
`protect END_PROTECTED
