`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UPyhS+bYJermpL7VLosCRGN8qCbkRK3+aqHtDO23sp/4DqVeBU+c5WXh2sha8K61
TjQBANq5KwM+1IE9Z3A3RJZ4AxgGIYbrs0dS56yGJjFIYbB2IoIQ0YDgQ324bCYH
soks7hHvOEiNmi91njGuBkCmMugsyIs1yzvobd0BKwFshJMPtUaJo+gIQPk9jiXm
1eV0iaF+wdlQnznsPv3hNyzsifzWFuSs6g9SB/syOjnqUOTH/bQmahXxbhucTfom
07HBWZ9JCRiwVHkRQbyBMatLR08l+YoZjn1BsPoClZuBBi5+qdpOONaEw9X+ojBT
8Nfaz+8yvzAOIfBaqctGn+W9qFfOSE9Lyck1+FGloVW1ozQcAEV0V71f6B1CjN7/
crSiGPXH9yV1zbXOSxvzvsw8Nz40j/QC+l2WH2PNwoJp/QMmbGiuY2llXDvhXZPg
GBU8mYP8BUXMadjr0B+9URJqmdLoFzaxuKb1W2RB+04tBlzJfmMIkbkoQpRsDCfo
if12sJWUfkwh/nsnA6Pm7Fa0t9tpAxAh/STualj6rdiu3tVpkp2icUMo7aGIJjEP
7td5sk5egCwcg2RMPI+kFrQXNMYX7hI+Cp8XcDFOrAUix4l101KVydZY4bTufqc3
O5sT22jFxwJnTF3Y4UW8eiXJQj0I2m8OZ9JTapwrYAQksCilM5MWnIc6ZFqmjgGy
5r2of3do3YRf0zqPluxCM8rNdVY39efpaKeZoDRlzfB9mMdtQN/rM1RgF9D1PPmI
UZW2I+WVVErDq9wr/OJpYPkl/9tQrjCKZpSeYpcFkFbHF4FuGJzZD865R3q6AQE5
zjF91l6Pid+/t/2KpPpNgh1Z5xCAJpArB9GNhea26qyJkaiwhPyrBWHdAwR6GHbt
N27GEPqbS8Qabq4l5/3oRWwOwqolpHxPNcBZ685Dx+Aj2BX137B2QbnKXV0wTWPY
v6LzU4lrUawS9nd62bCIqyT35qSwzjPz5XJVx8CXfnRxKCfH7S9p7L75SASYVLL4
`protect END_PROTECTED
