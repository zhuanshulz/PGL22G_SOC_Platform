`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rEpnq+8wdf7jU3Rxfq8kPlXLMMp9t1t2hDoVJK5X8Ut2WNkAfbu45Bbbi+UFOXDF
b7Omw6FoHJ3hSSzM/ZtnPeY3yMjOlX2rKQR+HSRtTPW5Tr4PHtTevbJQ+v9m5icD
XbrTTPtbBqB+hMgAern1PXqBQaRsU0VHsqD2EDgp3o7bMw/WgPAZcEF21DhxywDW
YDjgN09DsM89Ckzyc7BTQYNqyUlNd4TJXMeIpWVt3wEZHrXFYXnEDv13aLZijdk5
zXUkAQG+0DaJjoA2rSiFhaJ03/oE8qXyDOuJesYtSJS4qkDirGGgia9m3k2ZOf2Z
QtyxXKrM6RyPCCqeu2ldmc5ugik32WqJmmUq37MjGciM4VesdNEL7T/uRq8pHT77
CEZJHm6bqfST6Ozn719+2Fjxjqzn1o28GQrxbm3LynNvXEYF3fvnDvvsGulI/fdp
ji+GXhZ7k0OKvRdugEWhmmCMzKv/9CjfmLy/48xx+iUgGpWtqFgM+8cvaYcPdf3o
OxZfjkw3epqwqOc+D7oMPFty5sjM6INCIjOOUgNWk3Lwa8EuSks9QS4yiO+xtNk3
1XSoIJxRwJ6cvNojWY5p2sMiGXDhuvGBLx49CEEFDyIYQYzEWp1gLUpJs1Hp/XF9
dQd7yHxcHUeG+Tdn59s1y7YLJzyhy/m6ulh6O4LwgDgNbH38heZQwXEBs1pmykl2
dKF45ywE2YuRZ81BNAXQwBkDSNMgGDZ27yLK04gPInlkUgvN6mePekZtEsFdIN76
Q9nh6m5i+5VIH1JeuuZON1ufP3XRfvk3iK6WEBAzOwbsI5FrPMkM0HPYQCW9NRnd
mtBweNLHFeuvhnRDTlX28sTy+2zxobIxaTGEq2Lncdxv9bQlntcxdr1qmdlfB6BN
+YUjR/+/OFz6tNEFHtZWY3Ip4v2Ro8y2lsE4EJzuCznR3R6K3YjmmRP/jUMV/B/j
XuUBcuQr821W5FHSEvpqa2Q8Azf2csXkSXU097yOufrQh6e3eCUayxDr43N/HzT9
m9A2WwxCDm0flkgFjfW7V+xjiR2LJXE+/p+snFtfBncvcQrE1XlVZl7JFZ6FuYh0
uh9wDjGxbLfFGF52+Oa41Ng8vz1FCojehPkznThTg5tZv3RU/qm7ghtNSgXRYw+j
HOkIyH5Is7wpUvgWUFXV5czY6nY3IsRq3qFLei+TRw8DJswoTWc208/Ky6yE/jKx
frQsQ5Hz1moNFaFdSF+cwGu9vOmmYujYrt5s91WBbXpp4VIsSbWeEZ+F1+ccqV8u
0gyC47mYJZZksWR1onUOvd/9TANrC59syHjUFdDA7n6S+05vOZyOXEBA2QSqknDQ
P8MUQizWgOfupizKrC3lV4Mmjq6aUFAsC27NDYb8fsKkttMBLWe+Apv70FHUG+Uu
Q0fOqgfRtDP017w9DmFHlG+KaabxW8aWEttc092dE9V8NUnexsYFkf0HN9g6mfDe
IqrJ7R3ActDVDtkb2+UMdJjQshcu3o7UW5CYmXoXB3PUCEs3E2BaqMTkhdumK1gr
nn+ITAsQnQNcWhjL+ysd2pWAp1qvSUCSCXdww/vj+GOvie9NeVUMWi1+Mf9sE7Uq
FMKKapxhFhSDJ6xWYAmcM54UnYmuTO2uSwqOyqMAit95h/Fy+p6OovCagw/bEWz2
W6HIT2hVDvVBxJMXSKJL1dcINZDKFPJlLIlvuPwzOmsPDuoRzTTlI9pASbBXMbF6
q8y6aDCONuQ6mUvOdS2pJsq78Yb/nfZwADjWVpcjliwjKH/s9vKkx1wkly6M3z+e
3wymzxu5KE45jy0LWy/j6gfD49O3wzbarL+sCbPabSfizlwo+bkrIdxP5zlmzoCE
4uHH0itC5KVg1+58fdWRuZuGlp/rn53/Tf2vBC3WsrPP+ttNSPtjVEyN9gAl5WVo
GAKKoq1JVbR4Gau03dOzfLhBuoux25lEyUUXbpADOGWR3Hx4Fkb6/cdiJ53gDYD2
GM0//FsDnzMwTKi5clr9qMilP5QmtZlex/FNt75qZqK9yW8OYD4GN4CtEOXD8udB
hpVcl8NEKe+IDb6ueszAf2WWpBCbd79UQCgbMhaTxw03yYf6Szq6dqaxS2f8H5Gv
gHUkUt/D01GZgjjYI8GGjvQ6Qafu052/Ovs177P6l1IAxIJbaCx1nMZxadeq6UP3
W2i5vxCRZcL11sRvCq3q6Jz8ugdmEFkzkLOQ3eBef/9RpbOuoWEI5WDsCXMpJDIe
yR91Z83uFOo8MgM1e8T9dXgHLx7Fqv8Dis8DW5tqfL25JtXQ/qdmIgTkhzCCF8TT
Q01qON+aVmBUcTdVmlEO41s1XXYcFDShK0a0cDxjaZGknelLLsoMFcpO57T2wPhd
eyDZImfhpL+1IOmSFaLnDhlIw4KF511USd9vt65NI7ZSY/+qOuGK8PoR88l7tkQp
vt8xnQVaWxC896Pq1eDih3OqSdX8jnszy6xNS3RjmUg9TLV6uPvBLEYKQ90U0I3N
7kXJmkFBJVn1haGyQl6Ud0iNXWsChg2ZtMXOOWgn+yY1Kbx7X3SSMpGRbrjSrH4Z
AsO7YvNkmayDAwoJCHCe0Wc23ziZfEZ4VYfU1+UIj6Hkm+kCMdSNGUVSHWOIGk5w
cqBZRkzRDwAZtuJCcM3z4/W323l0DtI/8Ht2+ytfI0tfeNn29lJK3C6UJucaRi+D
ebtkbTiUYaoo3LX51fYuoqKwLsE9S3L5XedwT6bhnU3eU1hISpW4aGf9V7/bnM1+
BkrPKjggdK9aXYC82H6YF0z4IP0WKw1gF3hxKOzTzmnO6/PAunHYk1r7zWUWCEln
np9GTRFussZseYrchyC2Zxd48Otjki+0LWAmHkdbZtfLeoBMILZ8yhr0EMRfGj/P
4HKOqIiavYRyndFkoPEPx9sCzACeg9QtmEQydluq6D5OzzE89LyA/rFo3GQQek3f
11o6FCGvh9CxGizSiYnrwB0kJin3Bo3eKNxfpFwh0QPOuFz6j8btNLeXIVdMNqgi
At/c0SwMg45so8b0QAk59YSTAwWqr7ODIRmyrSxLfM/9VjNgnfNQaMMTzNhj1knQ
4CBB3llCPmTboWo4X2h0JNyqX/tCMhODGvXny7VuPztR1Hs2/ZvnwkAZR2IXdVSD
/1ENeyE309oXUmoNhiTEs/7k2ptNS1N+zFcd0oRGUC14Yhbkvs2oTmii+yXB65sl
4YdCd9fwrSKRoUB0mQGyEkN+wTxSZ3rPcZ8GwxGhiZbuoBkimHrWnoubJtXM/nSn
Z8xrcgmpWeoCcjFRPuRZOL4xxny9yomYfmEhATh/MbIcxdRjvU28BptArJlbnGNZ
SJ08sNZqBuXnOZcC24ZrMaarjtOYiks1hSO4uvA/G+IJVj0qUc0oM0ZRHK3UF/NC
SZACn7Hk+s5Z4WZ6X0m36g==
`protect END_PROTECTED
