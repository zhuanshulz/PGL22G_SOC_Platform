`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zTo+rWaoVA65JFkrp5iI6ul6Ei2/X7YFx+jpINijcmif+JH4XV/i3KDcC8N6pkmd
YKa0NBCCTrGbBxkyXPfT09I/jarMFZ3qmz2u2Mxi2YK2O9zsL8DcTGHfW9An0F5W
a+3JVy733H5/8KGBIAPgbFOmzPY8PfmQlwtzfBkA0OfhF6N7g1T0IDm0osi7W47N
aeTBUmCfcazNluGwZMR2EKmKbRqgIlYKbTx6j/iqQV/DiDaR0/zeZJqaOS+BcvWz
daw1fTG0Znf1TpFHlaTuy8lzqPt6abCz6FKEZulRQa652OGWHrTRdHi918aDWG1K
p3dOf3cBy7zq7YvV30JOiqfQHPT8ghqDHUXKJIRz8VRYv2oZA22DEt6wP6ATN2Ly
M6+28q7a6wECidwNDuKCKm9ZdRvX6ZPEtvXv+e7zeZl8QM1uJ7a/UsYg9lt50i6l
53mKY9Sam8XV1tohiCTm9wVieiMQ9gtOHseSjAOqitUGDbRewi0xCYPOgIPL9+lY
OOyFxYSm9OTBamGgeUT13rqFXsCxGbG2u1h2jbUkflG3Pcyf+BBDPfOz6r4cFFwI
aVtmXgYz8izIOiFcURO9au01LKP64klzB8sN53F5T6g=
`protect END_PROTECTED
