`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UH5qpsTDY7nl7kheGDqluocMHg2xBcu6XbXwMsqcpV5mGHirCPP4nALMODINZIBc
gHKEoagxkrWluNCqNIsRMg+1w+zxsx1JIv/uUpSZxh9OJ426GiMkKK0E4EyOdfuR
PS6l3E9BDRwEMmv7obeTdcoPJKyzlfie9sA/HvSokRF6eVG1z9MHZp4r7+jmKyMt
wCys8TKep1CUI+HRpgWCYaas6NpY3/50gqaWAjqqu+fDmLWNB0y7zyJbFiziFzXT
SmgSOGSPy49q4M+loZpI0Xk0999E1uPhlpZpgiXrLr3XGNPadpOF3S3rDStUSVSO
Uq6S/UvVnp2cCgG4YQ8QNwkGDwZ08Ojg6HhiZBgmMFpmiwdQ6XZlLHDJQPQGFTPV
v6dc7BVkvGu120L/ftuUqhR+a7F81oQoSFAZF+6K0EHIikkIOuFMPOhNO25TGDay
vXlDwYiFVOqlvvw8kX+R+Dlb1AzeS0HXiErZWD3s8tsLtxE+tCo4wEvOyNBHmzH4
Q3mzhmXcZWIQuJ0meM4hgljZt6VzsPWb2qaborbm51IFCTi6poQa475tOht2jle4
uzNBUdG0DidCcCkbsT9ACv5lu1S3m610FhI9lu9F9/E0PdjyitTCx5BoQzYfbjTb
IXtmHpMoes96QNmL6qtreuLsY0DVSqRErWXlsMTmEJvWILsrkjXU4bJHxDAzcYWT
JNqv8zsSW6PDT8NmbXrhFmTSLS7Xj7n9QtbydiKRxGla/xgtVbMDxuwPmIJAsyQ2
G7kGntxPiJ3dWmcEX++clD8OJet/sEpYETqUULnzcHKi7U79I47RogGN6ETvijjX
RFe4CaZfXWmruvw3bOwq2+bmUb2hhx6hvb7chdLZ7qd1hvBYU5s+KhI766mHCuPS
2hPuQ1mFT2RA8CdE6kkHMRLneKORKP+feMkHrxmppUdgJD8J5OJvYZvf0g+x+HNP
vprmM4OlGe6SUPZoyintNzY0pk8rfFni5wS1ZAXHn9rRrz/qy8hyFrTS5p5ZDFgh
hVw6j4wSKj8vxPhcrshPswtF9wskoXSaIjyqki7Xt4UOO1kNQQK1LeNxyhyhQQ1T
JFHM6CQ/QUkDw7iVcz6ePGaz/G5YpZSMIkfr9J7l4Fn3gDzIMInKU8y1S+G/3Jh3
B2nT9pb0/HqAdMUePUiU1s03hcPrZC9iiVZdqLvIspMsx8IGfmsf0A6yny3rGsZv
AzbwBiI0DWLigRdp5h65osztYNTxXPF7hrQYkt5PFJ9ZjeMCALOolkASy0m8XLd+
Q0GKYwhjMbZrQRuGeI7VgKvWbG7bG4ujOKhdAzLrGEab+xA7XUPYPDJ1nDY8/7Hf
`protect END_PROTECTED
