`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gk6EYe0g+YizBzbH+rDAQDJz38yhrX9n0HmKranBOCFwPf3LYBYx9XVdkDE4U7gv
s6nbzUpZSd14slKswdj6op0GJSMvxtcc1Q/lA/lYYtLWEmSKZlsvMhuRGePgNagL
v/HzDkbUk66sGW/LAOhbOHCIgEZWuB3WbebGOjWcrA/tQseoL+5NJikAWCUeWOoK
5cZzyv2M6CtO168270Yzg6LDJjVv5+fFBvJz1iYA+PCrritKM2k7Zz8kIG/hcVRF
lo7UuyRIAcyx/YdSmM14TKw15Da9nWIlpGIQADq55Ja1zXUGVH3HkOmEMYCzE2Ix
/feLK3Dx7wRy7z4lvTTp/XjHdkwDQs0DpFFIGh8BabJLJmCBrSBZjxssuyS+fq+S
DzLYy+D11ZyCcox618UfMLcGzvtu9MFbxlzLewwqpUd4NDNBqAIXfIyNgsqrESvd
xEqPyOW27wHhT8Tj2TZXpsX6HOlLCrp1UgAcAnsjDreK0Ggd9Wu9MthDsmC31K0S
ninKuH2Q9KJ26OJj7fnOaZOhLZ+1gyJ3REb2C8QnE48Zbq+gpTHn2s61oD97we/x
/rud7VX/8o9cSQQZJJiCP53JbhFj9hqtLLqx3xYAD2a2SvoF3Atd5JQGg76oRiUW
actRBQ8JwXmaXZFW58jGvB1KqDeCtIsBN9qcp9ZJ0YK9oaxmIl3j+8STf/Ajxf2L
xDmJp3sd/pM6PUf+87l4W5oYEhxTMmvkA6L/NjaFi1cQ6LpUNzg+qGawx175lLkP
5EBjokTCLrdvpII2Se/+7JRroM+Bmx31XOcixoaed60gVVJYlThCZWw545lUi8bf
WRVAcM4Ee62NEMoyADMwpoAg9TjbfJUGoreEij6sI8kl4WCgC5rgbi6ohOPXxllb
CuFIObC9bHpLu7aoMWOgihzVTwj86959/zwUuuE6IHg0WoH1OorS53gAvWJrXVO3
drCZCcaeKFrIflkq7pps3UIBFMOJpczn0/I5t2pwTO9hdQkFtmq7FFPHaj64ijgf
Mll/QD09OeMaA7DK+dpnEG91DyrQlw2E1DWO5Ebp0U7ir7hxCELU9aoyqxmiQosp
rRkBSHb6A3igTg7/VlciQtt7sgJmr1Hd/dz/RV1h2J+Y+EYS9o4fjKCRslroBEF1
sxdYy4jDjKbCPf5YoPHazyO3KoH2lUD2rcVDuXmZmTszx1zf26836kLOGrDsqd4X
/g+RQxi9PzvJUNSauGkL7sECnAfx7giOtDrV+mqb0TNK7x5zHishvCOvVVqvUXwp
ZE7/KuqAqAjwy++malQuY2Vkzb52K5UHABGJ/R4STOWpXuOiL8PlV51ZAMWc6xOh
DeUUpHkQOoXjsRZjQVx2Vs8fhiAWaiLO3Z1PnPvpG5mDU/wdNkQkLpV3ZA6Dlyry
QO2fEEa7sLR+1FaIhNhIJUEeSS/0PmTofHLLYNvUiaXHsTSRoECGh4IefY3U77hd
bzJ8AonMhhbh5sihI8Z39H75M4NKV9jzd7VgvNYydoNOuwFkHQRx6FV7kPTmoTJl
qq2QgAPaxiesNIFOWbAeKsbqSfRQL8dq/FlZWxYWK/t+YeQntXpTE3S64M37zxbZ
0UNVOg5oqjUxg5ge60ZZK+Wz9Zij42gbH4vjNvufRWpbCY+3CKBJffMsXj9HHBoA
0pjynR5viMNJV55oMcs6rnEiNJu/cw920pLH4AQLsCyxK2hA7XYyrzn7ytCT0SvZ
Q1WG2c4Lk0moj8mu6ziOZnc1BUBpcEzGdkWL2/vFTCEaK6lNeFeUPaDNcjwHb3qW
talng7HM+dUQvUAFrCJnEsFMPxMAuw1V3gSpjCzD7O1M55tNdYQr2tMIv2PXZoiH
CQ0uf2PiIQphfUn4v9kwh1NNStzb4On5vU8/8mPdO/hc8dwS6VKbeLYzaGVo8ixU
L8tAVYxFf2jqoOp761B39vU9tZ3zVIs7TuhBc4GqNyEXSb9olXfkqzRqrHiOiP/D
Q1M/PXlYs4YHBXy1J4ncvvNiQQH3Uas1GYEqKy3sWKy4rwdW3wEC1u16Xv7KvdWA
3IRHKDcCGky5oEWGwt+Z16ei86Ycm04IE/1LL6VbAX5EkezdLQZNjiNrXzpHU5mQ
mS2sWJlfK8IAfQnJJfT8eqojBVkVHK3UpnJEswzc/8CSwcpzDH63KVKgLzYHZHCd
KpkKy/fdQ7+Prt6oB0lLyPNJP0c0ZDWkxcVycZnO6u5vwwexqG3iuyeCOJugNH4S
ezgAQNVziEpkYY92Sl7v7A==
`protect END_PROTECTED
