`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5F/RBB5R1nSnEZkcQd8hmHBAPmVnPTed4HX5Htq9xyT/nj4VjPX2X18/ZK6Ny9Da
PWEqAZos3nhLdcmQJHQLIqYu8pxP1avmd0G6jEhCsoBlbB2n0r+hxG+ktkhKn8wr
0WIyacqTpVu4DGPuzKFZCguQBay5LPQoMq+rO1gVUL71pFkgXYrwcGmwiYyrRlRn
z+n9J52SCT3ylPePREBMxQ/z0L2lf4SWJjGc2I0TZGHwpambjU52xv31qqpfJtno
A1BV4kjOFWFEV9bi62YOOT6bUte256dB541y3GtpkCYBQhJqUnXwe/Or9vRBBrKX
D6ObHFq8uzYwRjJmzMDWCOvgpkqjrck0vGM617FX+vI/2nvGiuWMQsOlqiYnJXXU
opzwXIwlkAwbkq4IaAomPQIkvpZJIDKztFSgLA4zszg=
`protect END_PROTECTED
