`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6pPxZH4jGnkk02+LRcm4Nl0Pj9spaBUprlUnzf1SHYDMmgtOWzGLsj2M0I02Pin5
LYz0TviDKnNc+UsVLnwl0+jmtk/3Yo8C/RU2KFA5Jtsn6GNT+jVxBJ2AXpyUruYk
jTa/EJWi+JyIaPiJ0AjxZTwR1Cmlf0pdhKjmSI/IKlvtkpOHFCecrk2U9oExqGnO
M+y0b2zrztPs4Aa9Gjj8EeKx9DkJjKZ0AgOFcDWdVuaN0kQfgvB9++48SsoKHT8m
knvuJ9yEnOmmPpDDje5X9aMlXVTOS91P0Ef6u73DMDG01Pu28PV+gquO/9ZhJDdP
pFhtamf7/11/QMBeKYpMHwm7vtxrx32pCmo8vw76mFBCjRlDm+e/zVSueL8vGmRs
qtN7ntRuMCS8uFiEiAKhK1kto9eEdf+0Duah9TLQi5dIqfbJVm5rtf+DboEUpTYQ
Sx1469ND+h946+WetKJZZvq+9pFA2IOBpNjjHSOfzjZr3XvBpKxo1QArE8oG6lZ+
8H5DzDk63c1uSPH5nrdyeHnTYqIb8w+P0Lkf8ItUUsCjFZJa2MHJQPuzGVnkKIWi
Dgn6MZIkWAM6QP7bG9psGx1ZCpDAgh2cjADYBWwbP4xSNVuP0QJTFOuVTu9v6SsS
vqsmzIy71IZ9LGj7KFHhAshlUHCyBzRTwEaiUP0YFoGP3kCtkI8j7OMpE6Cx+8gB
3O58g+mH2jkXd06GLXJlVuu91S9tC69axRdWWZMcyo02JsJ/N6P58OhjqmAnn+Qn
bYaHaaz7zGB8XF+OkAbmhlzDLk1qyNVRlU0bPSCc5aj0R6+3WKsYyewhH8614pZ+
OFMKHsniWQ11Ht//Ddxc+aILHHCiyHhSBCplvpRIqs9EgqPYdvNSsbmzVIUsP3jr
baqz3pl/tZGwRMUkiewEFJO2IkzGd9EmAD3WLTZ8kmrjE0ljnXLpmko6/xyNKIT8
Ip2MWytagejEMd+Kc9R+pIf7pL3asAUZtpFguS+zDCcpUHUlbbc/Ps5OinOB16kE
Y/jDSd++tzrFK/JhIDldCKRqedLDgmwqSU42yt2Ll1PzgBSVi1Z1wdjRc1Od2mm0
cCrjYTwxUy8GDb4pf1ZW/706V4rtXHRCsaNHjQQIje919HRWg4UIHfIIA+aL1a4e
7XkvEOb4Ek1P7QflHv4Snt9svpD/y0TN8u63XUWCHzzYZt7TqSc8zeLh+wY8IP05
46ZCgSd+v1kw6EUZaxGZiba5iyWQW0vY//SmSbr5zYzBaVvxozHdvtZTMm2xsR9t
`protect END_PROTECTED
