`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H+tyEP+TQGmByEgpKxSBKrESJkS4y7xfe1D9s8XWwzarRfpn+VxcimPE6HLcFy3G
LzwxM21wXWmJcvU1DIo9Hv0q/lhXfLKSGDjzTe4i4+3ST7F9Um+ysN7KRnowHbWt
xVJ19a4IZ3TfGJdkCjhTLCTb3+F/ky5zaE5tuNYzygZtrXCdLfISSzL/dcWUZC1e
Wt//mjXDPnYwjZRyCLMkEZTrJv1+evmt0X5BI7eAZsAc4GRHVLzFdmzKYUPXeiMf
QdOOWb57V6Tymz7afFPZrW6Z0jmL2oNiPZQLVJfMmhrvIpu9k6eMdKnQKXiqfWVy
/Kp3//vwZSZ9uyBur2rvqYymepEe9jUWqyqBhVEWl9rLMntpM+IO7+C8XeMtf1hB
x1HAPn4ZIoNPhobO1esM7rnWVRTixNsTzjwjJi8h8X6jxlzK+CH2sigBAh9Fg2HK
pUBsWmas3mSnBNS4L1LQXfLv/J1w98HEEN411SoWjQeUIa2lVlnL3mxzoL6kRGCT
lfgqOtDuytAH+bqFj5TKh8xhx1Sj9CBl3NDGwluyH6WYyUle2m6KbnXu7tuj0SaC
kb3e9efRHHg289htisZRmBnjR4EGevg/esPrWcRLEHcSAO/PkC1bU0tHAilW7WQw
8d5ZxrlZce5Rj6BH14Yy0vLAtYG6n+WVGG4p0I6BUN3M5ZHgdiCQZEsYsmBcsvPY
1nqqhH7C/lGL19H2HYvBNU2ZUfMwMVDNsOIZif67DZmgRfAWJkJr+ERcGGFTPxpW
ZaQw79dbNq7Zg9mQklua6DpY8zdHeLXqnYprc5Odoky6oBbQDT998YboEQTyfjRm
cRQWVWi1/dhc/+QHItlYc1h5esacRhYEuhtFK8JvEIwAge9rfceG67M4n86ow0eW
9lPoxbOWuzdffKGtDGEymOr5X6keTFvzvK9LSUa+5wc=
`protect END_PROTECTED
