`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZkgMTpJ1ZihX4PXAbzxBGNIlLPphC6bkKMlJ7ELOiOkQIngUQzkUfYJSo150FgKt
F/4pjhbttqFSPU8S+Y0Gmrjs2mxiD9fpKDZt7OEUIXEneke+qYv9O2OON6IEjaNw
uAmP6g2XCqiNdD+QrZzNrkwSSCKWlp41Zvcgh5XXvbfHkLkiLcr63z2zemQIlpDE
1K+dCw1Fk/5AJik3EoLrZz8itgAEJax3nOERcJEgX8a9SNTYQa6KXCMasBa8AZd+
+Me4GX9UeA03WvZIg4vcgnEkpFLyaGn1RX3ZN6wX+oGuLC/Zn43dzjSDADneEl9y
V4TAGdx5+cVXBWaUkS+h2oX8dAaWgOjlKp0RsEU7SV/xeQOzj5DMS4hRrWapYZWF
i0v79JCTKutAKBFoOPsqXEsBznYqMOU9eYnnFiuXDNhCxx8J88yKuX6fSesmJE6I
bngqvRnr3CYvF047F3m4mjKTX8TKFfe75MtMxZzEVretBCuDT/xydEYY0CPgbVs7
4MawpjlmFg7pHa/Wkj51Xf1oC6aTe2MIE0AA8tLtL/cuVzJh8QMR600aOsaCfmJ2
uQIdp0gNZ0gEGec/8ZEJYPmuJminlh2FAen0fwERl0S2aMobW8VgnlqzsYp2HUDe
7HRB8fhR5IeVDMgkF0O6BzK9njx6N/kwmYGLB5Vg4z5fcUbGuYzQw7ucBlufBMtx
oGz8S95L0R2W+K0uzyAmnfsvo7xV4OR5uoRUGq/VHzmUMzF0YTmduwplcVus7885
chPoNVRDzhj4th4QtANO1eo5sZIl8E3pSRqQRBLx+m5fQNGDFiy5GoWiWMAIGNGa
RxIBD9NdlHz3HBxYqQqn5ZBLXz0z478d7Cm1hQGX9oF/MyyTMQPVxiEHXaKYVVoY
v4PNrECQPGCORYkeOCXKrVTpNB+q4+wlS6bsLlPyOzeFuV9tGFZM3Q2T5IG2tjIN
o8+Qp1xqBD+GDe/YSheGfCJYhCGw6GIAJFLDSdv37fXcrcd4POYGV5c2FJmv/E15
1mkJrYvcjtX2TPDQOx/IQLM4kxf0nOEiL7PeCHBUZ/XBCl+TmwFt1tXDMLXfehQ9
h1gzk5yBOeiHcSYDbDgI1YkmfwE8EBCYc/zdewFS1SKWYR1UFoEhXZH0Uq7c5ivA
psgJkmVUwbcpn71ljNYLMgzfyw8uMEVlp/oEI5zLXsdG1f3mw3WPNxfFJFKP+3+f
LT67G1w/MmdRjG1ZbILYSjR4cgLNZiWv/mYGXbQr+BTecnrMUvkT5OaDWhpemV3A
W2hcSjBZctIHRIPV/nd6Floy0lftgmxr83nX19/JzZs=
`protect END_PROTECTED
