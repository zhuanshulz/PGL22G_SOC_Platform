`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SeJ9NtU753+J5pX13mqsDTZZkNJkK75oXxrz6YWyKgnwEmwcdpIGhol85D6xtAnq
Lpes19tUErXWI19dMhysHccRQMjmAb+SJmjo/7btHkXizY7vjs8dWoex+VS/PVdl
Hk9OHzhPVqqTtZS80UhKRW3cWSG6NRxVv/hRFPJ97/knoHDG/s2QR0LVQhRRJsYC
b81H3xmFNk0RJIJDLiVMcqo1Hi8JX1Af3heXbGqF/FawfaOke2ARbvnfw1OQKSin
I31jFnYquaoxNoW+ETlU14dKv+U+O0BuDqyAQLtR2mTVhbHpJK5KOJ0AWbXTiicV
vUal2sK5VWrK8tBsAMALfzyhZ/qIC5v4KPcX95/PI024TJROL/E0gOzhaZlGru6Y
nCi2Z3fJnRJ8omRXt3wjsthkhnO6Uao2u9v3GpsgrxL5wkBfGe1IccTf4NK4D5Ey
WgcDC0FXVWX9kaQGllc6srbtpeTQKX/tRyxGL6AJJfERvlIt0QySwpMLp6igMPOU
F/mjnQEcfXKZlunDqmuobDDdbI+RkrkBo/t0L3m9ujWwQeBr5FzFqhgf1MzXS2an
XyC+k+nM+1+a3GFnZqb0JN3IIHOaYuInlQ+CQlv7bpxu2Myw1oTHqOWP1LobdgKB
CBkxIXV24joYoj/6pe/0x68PAnkoXuMYCrkBYUmrlzhfuf6hPIPlS0dyzp1Fy0zX
qbRgUSMMFXJZakgUkQJ4FZuxLr4WAdJSXp1hv77foCdDNhvDmhbb6rF7MvaqQaSN
Q8RDaMfCoDDp/fpjiaNdpjQpteGMC+cgSA9itfnlobYFubnIct8FBsOw7VKzDKtx
P3VGHlSbY/2w05LizdV+d1p0UkXzgmAXbxfTvE7ZBt5oIsISzXEYzp+hCxzC50wl
FW5mbUW7dAKtg/gEjmmS2r9hqeflM6+p7DA6rcXITRs9dXQdHcNHDlZ53jZJNDT6
vyUgE/U11F2Iejo/qWomj89+D+PF0qnEN3cP/YbNU1Kj2ydDk2pRvjsY6FZuaxVp
VhAf95K5R46ym2dWnZyYKOjxUXMYYl8qpI+sG8tbA9hxTuG3EbXJ4kJ3a3klg8F+
mkmU6mhbexDibklmjibbi2kwcDgFVHO3d48o2D3D/u1u31Q9Cc3k8+OceZ4P15Gf
`protect END_PROTECTED
