`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hWb/hYqjORZODF6K65CIhwvw6r/mVBfo1FsrY37a82NKJWcOtaz3E8qcgpdYasZg
z2G3K6paLPh+TvQnUPpevY+UP3vVzW4vHz4fgpQ+VDZPdVhWi9olgcS6L4G8dtdP
n1taU64wDhI0G9cjsjXc7H58X0Bplf85mewv56bGMQdN4nZxHAEKL3bsMOPnqFfT
5ZIdM1km9fbpXDTpa+bY2zhp5c8/BBjJPMJ+Ft0lLr8OhV1ykCQX4mCCJFN32OSp
jf0OJ6BPmOeyaHkIY98K3JudFmPasq3UM/KayKdr/1Vhxv1XCYKpoTDIyHFv4mtt
9a6YZhaL/8H7uyE8SQ5ZV/Rg7gSfs5Ti6hIzgOkvavsqu4kqpDozdS509paDUjN0
nVXkqM8Bkf0dHHZJHGvgIic1wu0GDh0WIBfzEKavESZEKkn6ktaTCBZmbDfRWI3B
/3hAM08Y0OzRm4XdUayNmKMA0TattMuawvVFWAcpdZWtf1tHBRlO9pRXtJ0Xfx53
a7Yi5Za8Sf5rBMOQr1KwssrxbdyfFAIGpdigUYfXIhi/k7MDmjy9i1PmWE8VYnfU
SA9fZdnJGd3xT9aBndwUsQ751GjqHzci3NobwEPzg84wXzgXpJmaIEWtfcsQNG7q
rliNfSlm9TbIXRDn/wyTJbweHDR5nFEA2IGEi04QtT3VxIkrYJMrMCQIWltr3vpL
j7jafcUpfsAyZAk8HXGIV3TUQ90seksCK3N+IURM1rWufTeetSbJM5rQ/+VC+Cvu
RwKxY5RtiPPoI7ffY7uePIwOuBmhosT3gvJd2D1aQxU9Zv4bZh0b9fU7EYmr+Op8
povR4L5d0LeqOsBXclFxK+i7LibMTJaqJBQLFyr43u4=
`protect END_PROTECTED
