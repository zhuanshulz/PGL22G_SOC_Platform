`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kFEnJA3b2onHKTv5UTH25601d0tp4Fwv5E5bjXmIuKaRwoBMWcni7HNroSalbv4f
4A2oToM7x7deNOBNTA5hh+p1Oe+o7Vrb9Hn488yL077at5aMzDXVBzhI4DVmYgQL
iNecC7fump4r80MEEodVRswtq104/15sq8+2dK56WxzNVMsItoD4zq4Flb2m4rUp
0U0a+EguAnjS4HhzQPHLRJpGLe9g8/NB9hW3QQqHTrwcFNUbyEpXwF9QUzCBOV+Y
4fqguQR4jrc9DDmZDS+yEdWh9/jikT1HOerhGq4Py0DBcy4pnjMd7cSUsLo9ghD2
DouhGzby+7/92EYfATjfJQN095FI+k4poEFNu7lbibOGDs+/qFmXK41PzsqSjQ2r
I8UTY+DTv8TV2HV5hD3xuvXlGVDbEbXES8GkYMYi/vTHYqxMqe6X90jDWaG8LjCD
Xuequ8drD5jJlOV55E02iAMcWbKnckh5b9G3E0akALSMKSiTR0Qd1kr7YhDSDMp8
IrTuZTelPp4LPwAn6L6GaXTGGvKGR25dTgyBtmYSSLy6f177bHQLlhTsHRrvas15
XYUXR0jksJ0yzmjJqZRJqTjOp83aWpLFk+pcK3hBz1rNpW7vH7Q2UXzUgTRkt9Wz
s8fYPt2uBgGmq5l5v50ZVLlzb/nFl14BPE+m7KYJhgc0/EwCOi0xGF+mm+hhnNpm
fOsCbbSetyzls80n5uQn31MG9vM6MwHO/L1MMs9+b18HjfmxjOa3r3KAZSM6rca2
jlPFiPNq957FQzxPHvUD1tvWkvIs71Lp3MpWU1FRSiRwTzWk73aCETWuM+5oL+4M
ZNbVsNpRGuJQte+yYyCWHJD5NsvFsmm5xgtn+PruWsfM9Kn2TpFsWUfkqVnG2QRf
9M0g6aoTOBDZZnuXWrwu9RgXmPXwntGjNqjrWmPYmYlbjNW46+Aw+jnEYkXjnEgn
kxAk5dGVPem0C5Hg7de2jbgZodlTyhJnx+cIdGyAR1Cu/ZHX5TVvrZRvQdiI5xp9
+5wu/0p/2nCJu8belNyjzr/CIReaNqcZUdB7XjgNpCBQxRjztmj/XVFTI2YRhVKc
n0fAJ15UsjB0doIFs6/J4vAh7xnsBJbTGABeCpXI/Q1H9KkwxpEcOQ+nLzyjWKy2
WxLgUC4cI7xkKC03opzEvROw5rXCVNzJY94U1p9pHZN7A8aw7U3M38CChPxX0By5
dcRtMpXNigOveYySDL1Ii9I/XzBAP6FkmU+inWP3H5m2JEIDyAfCWTi4UAp+HGLS
49rDHDshLjAHtWvfft+sashmV/q0Fd41BO/ZbLsKHOweio9k/9mpUtCBo8kulHBU
n0nhSMnwWpXaT7+5nMfIpQPei8gZKw+VodVi/pXLMl9pRngyRtM258/pcunlJHFT
PWCBzxdb2B2YYLmJCYC9FDAnOij7XaPHcXY7iW4rqPue+Jq9WF6zBrKXg1CCB+mA
T1X/Mv2R6rC75RCFFwJ87pPThB2VrYfGPMIGD3AKVqP4r7gOAaibtrCZKiqx7+M4
xAe06vhDFmQIK8o4zSGL5kwX2BJJMuZyESkmB+x04g6Zxvg8mnkCj6Jh2jZ44CB9
AE6WqdXjMdxrT1R9Vi1xEgHYFjYLqmtlUzPrKrjYEfXGkMURPUXS+FWIuCTzhANY
6ck7J1VCM2prfZ6OqB6uiBFTKC1MqLOi7gf9rrNT9GnU3C8tkqx1J4AKAn5TaK6O
DVDf1gt0Ggcw5zB2U98GoKXK7KfkfQLM8pdjT7Pe1zh2GNX+LpEg6POOA438oxEr
W8w02fjBOlBsvOnZC8Mcd0v0Wl1V4F+DqDpY5W5ekkEuIvOGVgsScLM2ZbZdB+oD
O093Ul7amYVzMT5sh7T6E8VOuCba6VZokdpDlxu8yudmD5IVgOC2hS+HgfD3rQdF
ta1kE1JkDqbHYJ+eho8SGINU1oEYPaU/SX2qvr1FSpV2ob+O3mw4Ua93JMOFPhrE
vR0RFwo/SSf2cGeiA9JMyjtKTOT9HxP0DHrgSBiRjtoxL9FWq5h2phftvLeNq/Bv
TK2NhP/b2grymzUL/eZGZbaM11OXpUkYPGaTU3iIITyNtl2KiQPvMEdbO7C/sQce
X9zX0svMPDR5MoXOafF/4IXRx81rtYYFCOEwSfUQ90/6H9DHiHN+Pb24cdeFCN4q
4vmTWj/09G+xomytMqcIPdtts8PiQPkB+zIBjdCbXQbIqTaiiJuiHTF9HdGuK1xl
T95OSk3p38yPa53TKCjQ8YHm0vM1Ui4PG1hKANYQngo5nUMPbKtQ76PuXr5Hrn1h
eevZhO39XHGmnuUsrwOnMkoQJHbGgFE4WbWDeZhlc2bPuJYEigstagIEmLfmbh12
t4tofCAShFljaCYA1GKr57QSA6ntRu1/34cwXr/6fkJrXQaz91fDMhvDMpw7Gtb1
bJinoFNbVYC0xQYC+MSGZ2vdVH+00MNrdFRUfMB+nO51t63M3E/jWl6pGPpk6gor
tRsnEcrwoc9O5rA9F4Ve+JFSbJAh/GaEKAYRxGZSDnT5F+/4tOSlxx/yNiBwD/Pk
MbTCloXV6GPjUwmT5Ih4Ozb/2LXlRQjsG+pYMICMCHbhRH22CNXw/J9YZUcVnJwk
o9o/ELt9Vio5afAY6n0pXesabakLb5sF5W2dzJLHHezuD1zt5IJth8TMB2YJFfBl
6FcAbR3duXJVa+DDbo9Nz8n/K50dR7s2Meo842eLmNQjnkFBh8QITh+9OjZ/JVd5
hjS91j0N+lLniDwKL+A0/A6j9kEyimBf65+bjeAbDL7tqFjSLQ2HMf2xai7tRxxw
6Ka8esD2VkDiaHKveRunkc6KJ13eqKXuKWgC0Y2nMP/3uLlS/HSe6aZASFX349fB
cxDxWD+BnjUiKvtCHnMsM2B7gR4Lm2UdozQIk/Rzn1wd4Tmo9sChhFB8bqMo57Dw
bl3ot4pI3gqGxb8548gweSrQ67TWE1Nqh/nBfh2KwS3tWMSKDceTQts5YSJLfFpC
MwNz0MuG3o/d93Qe+zCf68i3+ZzmRJxB36EhePO8vU2NI2ukNytOeHPxpp/HWTos
HZHy3aargJdSNJ1C3qtrBeBZ1mq7AiW5C2oieUZmg28LQHBbkDHtVGQu+3jRQ/XI
MRukfZuGbUEmDvSNWXReD7dq7OWoOR/TlEJzeB4vKkVbCbQx22cT5gmug9RLLKIE
VXmJVtv1rTrqPAmpefYcRKrgIlvSdxhnBL80+cj8t1T1V89kE0bTokr+2tC796Pz
8C4OyOxbDXuJaxbKvcicrL3TaLEjwdMqAM+0OaClBYlogMdCZrnpMbFMkzRG6tPH
hDLkil7rgZeE2P8vXPDJ6Vemb8eqCRM5Rmz+jE+VcnXcLkh5MdxF3BglzaXyu6Er
RSKmqe2iefgrRbrqTUCohLviTvZJBPruDxyY+hORr+btn0MFVk32/97ZqYFymTvP
IPGhwKYkxVkz37Tji5tYmDL3/hT9FcueawiPrXOnPQk+UU9ahdQGUR3Czhw5ABmE
ap1Q9qRrd4nCOLjEUY+GaH5ijV79CBKm7u3ubgy7+r2PUUBi74lstSoQzMn7VI5r
kSvfRTpRkO+grdKlKfcbz2Bs7WK8F6QVbYM/v+NiLv7h7E6kF5yBxMRziVPZX/oc
SKdfrJ7R6tpf6oOmVFC6kunYdNlPLYyU/r+ALNsRE61RZBbyX+Vy4xvq8/PBRzJY
XB2HR/HJwAHaXnclfdxB0cDYBwX663x1ES0YZrerNyGp8nABfRorJD6oFjjl7+Et
m98lCgyhll8NZIoOJzJhEW7v1Qtu5e2vG4ZKWZMEtE8nXYx/EC0LY/LXXINfNZ/t
0dhzQfhPxuyPU7eytrIsqxUHny4fzFpyhrcUwSWeYHUz/oKi7LIkAYHO6d6aFtUU
wFL33zzrYxexmv1jXnjIHo3xJC6zGmzhxUjaV+NRbUjoe2sWSzFe9eLHqdz6b0EG
w3aJ+qDh8s5RxsxpcCJ5O0qUMmTQGExbBfruL+a2l3+NJ8AyYciTEq0auiQlRJ/n
6Kmj8CXvPwvVTYI9rMRXoisztJpE6rCvOzmIXQlHmyRk5f/ftWV4rSEhVxWsMAkR
MX202sw3eGoXIgmDSHvOqVVTsL5SkU8mp/PgWoUKTPlX8owrMHLrMEZoov/Zt396
ZbJI4nmbw/ridDaxso223eJM5lBfyEuUiBYWRcLrqFJHDuKk/qs8npHsfsG4Ymwn
o2Oi8ni9FCT8X5FwjbbszErTlVb97OUV5N8pmHSOu0QbiVQ4D4u3j1qvBqQJY5cV
VmIs0Tn8YEw+l/YucKkfQ3h4JnWnFoYEd4g9IZ2BrdqVg6GAPEqbwcY3gYqQmXpg
//cwf79XGhm4cQSik4GB6xMd2Hbj59mz6LIb7tJM3SYY4k7m4DNtQFape+ZQuoMc
doCbCtK/DsjKSAUtO6mBKBBAfeDACx0n0ez5mMAHqyUgLPrSPETnCmssvViT4Fs2
uPxAUe0NV6g7c+QKYDBdeRFaXuPCLlTG12zDuvsj2AHQmQQGXG8XRZG99RBRCtpH
atca5GL/GIWVhATN24owHuqr5xHFyZLcuocEaVBUUt27dbQRXFX8+xD0oprU/axi
2TXzQcB8dOpi97GKHSD5o6AbxW0g1lRBw543TX9WJUIglGb7Rv17S4Ki2UE2kirk
WSk9A4tsgblrl/0ooK6qkBIRi9nJ/vTTqzpR0kZQXldjKLAhnjYjZFa9JYBk78yU
OsFE6mvvf/B0f0dxuwVQlo/g+gALj1j2FYF87au2xeuFxNNGzRx3CcskpAXliS77
IU8eUnfQYCLgaOW+0bIstSGlxqnuYNzPkrk8dwZ1bw27R8n/k42chm0shGYjK2hj
L7Mb4XzYj11kNK5FKHZLPHBk3oSx6Jhq+udEb15FMJmgMhMJ7UH796vwhlqaXtym
pGuzPwXYRYgh2yUHDyLgygnM3/VTZFEBjcS0DvwacyM2cVZjrgKrmvzAPBl/McRX
iETAJl5UdwKV8A568EkoAk8TsKK2Uqd5AdavInbiM6Um5tGJVVxvB4gbVZOC5MrO
0YUrrLAO6xngAjWi/7ruZYyh2qJJ1XaJqhWjP6c+zj2jmfg7KGpmpsdGjP+RDd4j
yK57oHL3HeuYzKaY5aROeaow65qzvNNwZuxIQ+3SviMG4w3Keu9Kg3mOPgmsQfPo
PYmCEyZD6sZf8dev1dznNwsYU8BI/37Wrmn6BkExTsaNDUkObIddguKkxk/xL2UR
ASvv2HRxf6ZZWLkEb6Nky7JKrCONDCbqMe2xjH2GEb/PtCjzoTiSf3uWFCJr22Kr
XcqSaX5oiHLJc+QGiZ1L0L4Gn2ZxCt0gcodpxnOi/IhaY9EoZe5tEMCEzYMzrFTT
rmAk9ekabktdwGS/TA0VYZgD7F09JTv5xNypvRiKLQ+XlWc5UHu+eXzUxzBoO6th
b1s+p6pj3WEd7K4elIJHg/dGkLk81KAMGvqslu5q+63w8A5ks66eE0W3a1bljfkB
a+woYDfIE7EdlQS9rRGJtrRE1Wyf2ZL6yBMgT1Iqbeh/9VuWB4k47nksG8j78avK
OyltYSk2bVOLcB+TRhVRsA==
`protect END_PROTECTED
