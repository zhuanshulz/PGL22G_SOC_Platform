`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Af86CJ5xAoOJevzZ33P+ncqCWySLjkg0ydyzafamMlCIlhVXmXiVeFBo7/2CAKQI
EHg657WtZ4gv3pofXa7wpZ4dhiHpW+I6WQWaSepGFDAIyW+u84g00e5+SDqzbGgO
D34/yhPE009uNs4I+Nfr7GHnmXxQzNyjk0txN5TouDn+AUX+/ANh5QvqNjtQeZER
KpuV8S2cdd58zShbRxS95hpbpCo+yPn1jK1shxARr7EGp7qQzHMtOlkGxd3bszS8
8X2gRU2yXnTZ5XvAXEACVKmawdqyM6tkdOerVYCeOWLj+G/WsD8g/p+oikMRXFKl
Kc8WnikoYaZIleWn2shAMLiJm7jBMLFpLykEG6/2oiMOpaDnAhPpk/vklmqvLxlM
clrXQgWT1+UDvaRYLyq+rhLiXNAG/dq9y+8WBQqiWtiyeatWKdquyY6S4rR6mjJh
aRMe/PDJxCcFtRpjTXetzS/EAqpinu4Ux7y9QvVFp+gbPvIQavue3z0dHHP6qqMl
LbtymOs2BwKdso01IxtRURJsb/RmK87wEG839W/ViBIU21XMJWu+1P0yozC0WUQT
vF5QeTyrgHmogEeSJScs/bgC82SbqkB51mRXymmxYMpzVT9cpX/nTAwiIFUDqfHB
kZVELq/AGAq8iOyRmV0fZKk+BHdhsJLz7QyX0WhFxRq1QCyyzZLbJ56B8nnDxNp0
Jl34IHnY9fXMPq30y5rGn9Ofq+Al0B+Ko7W4zf4ul4vqB6cmZnBpXSV3MWG65xDq
tMjYDMpAB7+w5rk7kPmYHsiIsAx5mtHKKaQ/9etNgKHboYMGrfmrw9thKCtcTOAe
yiQKc5DaBHinZjckgDKHwnZzV8nXUoMY9G2x7RXhrrseq7eSOiAbIKWaAsMcFz1j
1J6WntTeBFCDl0Q9BRqniupdMJrQXK0hDDQFgLQQQKkMBdjqsjhMh2BW+GFqQwt4
SSMwFQD8ydtRuCPn5HAGKWY366mK9sGbzDgC+A34CTdJHVChE62sdgH4apGqGWHG
1tt5ser3S4ey+Cpx1OifwTO/E+P/SaSIi90qoarYqaWeebDvCquyYeUWf/veaf6w
T3mSQr5Je2/CJr/RNjSwxzvCo9ZZmpqoosmmeXHwQf08fj8CI4LQYgZ1TfuVBtSZ
QBDOBYp4PTzwMla/iielNHl0+r19caU0vWpSbuHMfix69uG+P8sJVu67JRtjMuAb
Ja6SbyGYC/0Ff7uzSh/mQLbDjTa1ZwfC6o4ibPlEVkfOTvX0xtCIzYtHmRSDzuVB
37H+MU96Yovq0sPIvWFjuNThOJbVPmjQHaBvmyGObe14KAyGdli6w/vGF7GgSzfa
RKMrBLehaUZQ17vGfTOV3Sjr6kZJM2QC2TyhNSdFZCfChV2RucGSx2zDzJz4j6wO
N0m1mQY142uIJ/yz/QcerRtNeTK3zncJaRPe4yj4MY3aUrA/84RqCcQfaHOptCEb
Ofm/exuFGWOtsVHBaXR/o6W/MdwlvBmy/xApxqMCsR+iOhTNbq5enHGMlqTriMm9
0Bss2SjBETmgV4GfK7xHsqZbOyhNuQu4yaOsaxHK1mXaUSmWgal+LCXQ02QIY1GT
jzEqFgnuwkW9s69UM10N2v9XAmEmrjpzBjXnjOCnDy6s2RlED7LopbiDEKG1haDi
ESxeLSAOr5gdGUxosNWFBKjwSXi2nL2opw6kvXNrWlRNSLp0a9Fo8W2ZUuKhdWKm
n6H5DWQwf7q4VjZaaIWYmE0pDtg4DWz7Uk9ez1/eiGeLiqgcwBki8Z97VGH/Bmha
gQt/UQcyE/OYzsUvmQwRx9lsUel5wNohFn8Ek8gC8/C12K5/c/4qGEse12qezqxZ
/XyUsQrEENoo+7o9jwGJaq6oCpRNgOsA4klmZnYv9/AeflNHkaVPxMs2B0XBz5yE
HZ3q80gXnzn0lkmFQNGA9huaQZtYVkjpDQM7XuDd2BAHUNzbQmYNKT7F/JRw5ffw
sFmj9qjFYoTMU9DK1goW7WHHmZtA43Q5vDsvGOr+r4DLDVtzVezLFl/xb+6bO7x5
lsZ1N9vEA2tF6bhNqzwAF547jBwPNxnauLYiQFrtLdjIDZ5tVdle+cG8C1BGiCkU
`protect END_PROTECTED
