`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SCfbz2PayLVJiW7GsyrtCJezodrzDdi45PcJyDFw/eQvXw8NPLLCkKJSO2CitLM6
S9J8uSoLYcuSHizObMTjvugBMHK8i8M2LG1XaZYEvoItF9qbF7Ugm28ECi/hwDgt
UE2hjC+L44ezXV2pUjSjDV05ZMrqs82bDceqNVB+qQqYlfAfvDQabySjA9jsW6Pd
rGhL3SAuiC4OtBXwtC1qZSOfDmG/AvAum77v7OpcDT4Zfj4QujdzXWa15/4hNZaw
78Gl/9mgIDvkzM7qg1ghEL5aDeJv8S1L6EEb6t1dNRRC0cFovwVwiiOXXXK3vLAE
3IQK/rtEpVYexUoa9LEyBUg0PPig4Jp9/IBS1f8fkRNe8JrRCHWsh4rzY51cW5Jf
LqjmP2GR7aY+GqUVBaB35Bt7QBM22WxQ58jScWo7PMUO0hldP4cCNS/z9NfBjJqM
7myUO9Bg85jDn12o/9f+Xlj0cjKAy2oLTsBeRvLFn2hzKcNL9E+6W5nV3GCzWsEp
/DGysFeLCYntCnvge2JjLqB1yGSY8zkP358AfMIu+DvkyTVK9cbusA7Hlfn6GVRW
HBhiO3f9Kw74znuLgvERi04fBtFCnR/f33q2WOdbDGII4D4z/bWS9plOkP7AXJ4Y
WVFoOB12fqtTw6nBOzR4/bLfSgBg6IgI5IT7HYvcJHkXEGxnu4bbWAMeTIBKII12
4qlaX+14KGvDOd09WE51HOIq1IcsEkBVfi1KAIDbOIVW3Blvqi+4NQXKi816hc/S
tCZaa+hT/T+9Dkviwp/ccJZQ7vmmvxfeIgC7lmicxDiIs62mNOlzsH2JAqs+9joU
7O5mFQuYqFq7tdmjPRzI2CalyO0qkAuS+TSgQf7mw163pCFu2WRk10ri9+l/Je3W
VY4Sxud+PZm9LOd+0nfaMIP41tj27wXJeeqtfbsJ0AFmqAYyu8Z/haBCKYFSut+u
ZkQdXXghhsl//nYQhBBknXXsblowtWtkz/AjbUcJ1mXCZYDoQFixse8B2vlT9y3A
BDBm/5e0AM+Kk3Az+xeL84rOwS1C+e1ZieSMelSQjmg0Lp7cNmBmOxe/3uHXu5El
Dgi1SyRauq8NzQYlFOL7NDHkxz8lnfpQytsSeeZ0yjnDRLostdULv9NesdmK1NBo
PAaBFLR3JDFOZPG3FIH6i3UvQSQdsZvskmPh2+JmmHGPtHBmZn8w5e8Zz2iwEk4a
tkjjU81BGoTiMNlO18oSuWno/yPAqri61GGedwGEKNGYkJDrYnfFxOa+MMW/Qax+
HgJ00ex/UZPqFa83dIzyTcAiPQdMRZG/zvdBpuFCT191+QhP1phdKKhWG7CqBHNg
qxvytkk+bb325mHt3ybK98OQ+yB7c7JTEXxyofrgb7tp+nJiOozPsMbZL/vzfvs8
HuM7ZlYJKu/AiAL5NeexklbFUWQX+81mrxKam42H3cmflb3ZkCRcm+sb9ildMRJl
9BGCjwciVAEtaLUs3hkz+rstuxJZowjPzFFShPzD5TeyBdtqEfjsDiUokiF3r+zB
humAokFKkBc+6CwLF73W/r7cofK7+1cApcT/9z+BvqPbk0u0Gt9XcEg7IbUraIJd
HZSZGQJIpAGEO+/LxYaUSNOShXYEsnikfm2hwyyTDVigNigCGrCqL6G8lALtSABH
vWHYtMSKVcmxAj9YFzAlPqMDvc81IUcrt4pgHM59D0c=
`protect END_PROTECTED
