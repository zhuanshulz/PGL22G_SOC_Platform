`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6aNm8Uuik4obxI3++IOToEq1si5D+hRnH/j6ylkz0U1goMSmdZts3ZQk1Rfe8Mcy
oR5NJvOdAsXid2xp8ieEhn0apvLyBc7Myn0EofvUNxQ1PSHxGI+8CQsJD3XEn31Y
e3EiIiC++2G28xVlGf8daRUoRkTlEKuUL/EcUFA+b3Mqif+8fHXesjZihgef5FlR
iDDGpJfxpG68oCaCCXH66CpV2zAt4y/nR6qwFT5RWWHpA5gN1kDovC/efkdAP4Mk
YpfRTkbkwMKBhdf2Q4uFyGD8ICK70DyIfC4zS9owt0DFaUGgTpWZE1M5mIDXw9CJ
iUgrxJQIsxXo72NBO8DSgM9uWQqaT+c5eHWgmEZ1WzvMZAH0HG0UYaATllER4iMP
HhizjEoRBs1PVEh2Xee0S0HAEIRRp4upMljmKdgkfA3ZUkrxLSSscOmfHtNjUAlI
SqdDg/jxmSepzU95JLfVBU25dqpkbXCxtLfb+0gu38392baYxYzZwE75Pz4ZEmqZ
06+Vapz4y2IHZRbduswE07xHZ94FwPFtiEVGHLvXXWxinAi9qG9qQI2tDtDNOsqr
WPnQK4TdGfPOXPibtC6K79KdfLoTXbY94qJ3GbmGLhy/6syBZT+0z4DjUoHKWRCh
8EIDaeoOiLp1uOOeGfXjR1m6VV3K0TF5Z5UdXf8QWpsxCTlPNv5obea6bM/JCxTT
hV0h/wPE4bzvVkw9BHS0/aBEq97Ohhl7ByZVImDvCAnOo4g5F90iWaLTmanSXATq
HvIgLex3DoNH/ZPPqCyu4Nh2vY7zapvFDagQAJHe4BOy7w6X/RcnmVOXTKFWUlDE
8asD6ylQElQdOc2ZB5VRriIda/YZVrOmziQy47JzQcmZBOIVFyHiTvx9puUMJlOu
00qoIBs7kvkw4ZCvOidnbqXD1HgwLJel1EmjX3jmb72CC4uX6fVEGBv6j4T7MsL0
IEFqj7iUv7qqvfD+7hyNseMz6c4UybjFaikDiW4kgdOmMFHLrm3oVjeLGWTKRLs6
6jwgjSOCn4YF4SKLhUeTu+LLqPmYgd7cbS5AsCVH7VnEE1mIiBl9P4iJYvq3mMBa
S2t36QOW3302/75z3Yz7Vx5nSnSYQFkfaIB1OtXv5317lkamLfAiRnqtaDax/fPQ
glQG5YHnAGhlUzIqkVanMRMYSftUhTtpTTInAs5ODS7KdqYgewObjFqU6s8PbOdc
5AcSnqpMvtR6tjzmTgEB8vSGkQC/wF7rpsGcVmFtQmFf5AE9wRMzFIZdwimaWYHU
SNmf+tLhWkGXfmxFAectXGV1pZytdCsaKM23MQP0JgKduPS3Sv8asusBdfWRQA1Z
nm+pSQ2VkTW3gI/KNItJhq6ODzxsq6z86pxZMnq3ll4fVxCSA1AaZi52o1cIryTd
Ntj0tR29nUmAQVTX6Ch+CEPTeLMSKfJK7uDtLiNrK5F3wfrEBSx8DbO1XKcpplu3
CXW9q3MVZt4tGz6XUpiBsOiF46ZnvYH08TrMIbGhiTPEzCcdDoSIwBfL/BObCrbq
lXBOpKz/KtgN3vbJHMdHfeyn5/cJ07nuEVjnYMNOnGGOJKN3bb8pip62Z1y3ZB6Z
MtndB3W+LJsSh64XA1IKJgQwWv9YhH06b5cJNxsb836YWX61j+6BASPGJkG+WVQk
IpkHKfL8hDJkHmz2ANz0+5t6V5ryWuMR6gTJ0z0htg89HrF+G8Gay9y9x0qCuKBk
a5LN8Z6EZA/rgiAPrAsyxJx9/pbc4TVAWV0Gn7yaIhJRrEAUvkgsYCeu89aD7R8q
+qLHENieKmIJ3qfwxFfZzgd3Oybig+fQr964P8T3PnZFh3+9fj8xRemBa+GZB7Qv
fKebyTJH2TxCps7DeL7FqJAX6GxLLr17/7eOWmwQIoKyBj7QUh9ceKO8uT53/NZR
y7+srJDPCdL4ItWPoXGrdM2U2KyupZAscFe+nLMbrqcbYElvvkbKUkRfKhQLPmNP
Cm/yLHziA7ld8krRhJQSiXKUevQb/sMhxhIg0cuzx2cYnYAI4mrpZ5MaYRnKPFWz
nEU+lldw1MJ3uWNP2lpPmsoC1KamKiMRU9oNpaLzFb8qNH8nRo+h0AhUdRbF72KD
auXcKz5AWwWwkBkBpqNZJIPWJJX78gSwt/kNhf8a/dzg83SAsrzl4W60/CGQGztG
9L7HxpiYfKkO/p9+oMbvloE/OMYmx7OJ9ieAKgXaNZxQjZAG21qoHZ5maevKqO7W
rUVWEkpiEudgUB55CESM/+K/vQbRfIjpfi4VEk7/ODcHQP3J0Ux1NcAj51wHdnzP
yiEIh4bnVdlT9ILJ9BSs7+owvGPU1A8BcCkV71t/aD0SR/LL6GHCnBLnOOVghp5M
`protect END_PROTECTED
