`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2Z/79/QH7F/amc3pGLpsVnBPun1SRFYIxguGCorix5J0v/DuhMYffUDtiafBgzeS
Muv1Fh5iwXvl6w56xQDNT8bV9Kguoaygp02wt15pAYx5uV6xfw7EEhk5rNaCfepA
o0+xdkLdfjM0/hXWcgjMZuqqBRuih1E3febLRneoOe2+mXKAMupdpYsWZqRIUxqh
5t8vqA3oFJrlCE219YDjPbo3cCFmj9XlkfUeFEVNh6KQFST10jIArMJDURDtJiBj
t0H5zrjqWJ9WBb2axDkRZALnl68S5zDUDs2k72XiNjqDXyp7YeUobFejVzrjMuSN
iK+vciYW5aQmh7bEIt6+7DrXpvWkRiP296sqAX7KAFnMRy6Ut6Pn7fpYx8Xl+xlm
WjJKjHy2VtuoWd5IhKZ23o9G13onigT6yNz2gJr8P5p65W0oxw0oFE/+yJ7lmpTZ
WrGwUQWoLQA7Z1H6KDkGbIaJUHHt4ZIXQYxsjDAtPzL6SsTI03o87lFPEFRV4Jsi
j5gv4/4pZW6cGDSdvrcS5yhqR0Q5Wz0vMruTeVPksu0cz32cCQKerPquokIGUVvI
oqSu29g3z9RCAbHB9uebNBPLFt24pLiwsWHCUCL3YZM8r9ZeatigE8FUIy8N3lLT
W/TCII1sTc/ElsmYVYvNjBuFZVQXY6U01xCPRXzGfcngByVHQ4jcU5hil+96AOYQ
quu4R3CjPTUpOmzwk/hD5SbVyG9xYv4tP5KeaI7yu8A2RLY7fKyf24F26rLZQtYi
nj9QE+VwKBpu0MhsQL40OogsFPKwyHk4zqekWiCStmoKszzE/E+PMQDZ+aBEkP5Y
kVWOPXtfa2ie2S05ymFhDBtik0aV6S40a/DFxCFYQdgcRhkJ2GnnmOXVVpo/5JY4
dnhixeiKPPJ17V4i1o5BSNJ8fxOIQN1gsObGeInKKrTYUDfMhph9GlJ0FsYwbr4+
GtEO6fhkZ9j70v1Ltuk06ZvMhJMC+Hs+8Z4hYoiUV17PAORs2G6K5YhqJwx0DPd8
fB8fScF0puLOvvVkLA41IuvMpBNCs7Mf+PS4kzk6L/mNOkCUnujRNTlhZBWemuOV
zLq4mcpoU5cmPQ/Q9zHahLKHzazfnKSjrd++8PIpYkonQsYMLwtc92DxJuV2006g
vN12SJqR/szQ0RWSZK8720dxoCMEOOfEnfZvRbKEKvmCPowSWKpc98xgxH26lOAC
SQW/7oSFnI4qac/Vu0coDEIWJuZat9X273KkVELG0baIRcz5m08WNwEbwrRTO8R+
KCqMjG9aikl3GZZRzFp12rZUPXGhgA9QkibHk7jsj+8Z514P2ab7S2Ft+Lg7+3/P
sV3D8Ms10yT2F6Me5qWZjfjuCL7kz9Dyv7CaNdZVj6kK5E5kaJUEJqhGfCkhXFAY
okaiw9Tl9JIb3nScP9dE+YMsbr3MAJea6gXT0u6uxRIE39QCGm06wsJvwDCQKDLW
my6b52kRD1sWlXQKuArP00BhSJbxbNdxVNfOvdP6+kzf5FPADgAfWUkkXlcKbMZX
OAxHz+ve2qB7vMLEgkRkJLY2yONuBIaWBlnwudPXSxztBB6kVQAtTs7gXpLkb9PR
AUyheP1HGSv/gpmYC87H8VexX40jJB0Vo8/vGpnByloawwBFYOngw4AidIzq6qqI
dzcM4a4f2YJJ+NaDv564AL3g+4i5MAK+NS/Xnv3uWD7XvtdE1hZ6OfayxWH/FVyF
LiCyT4ZYKgyveaajsKW7eQHsLx6rP7afgedcXMsmnqxB4B17sOS1abeh66Kv3t4M
Kjv6i0LvgH4RB9rreByuhzmHJZWq5eAJvmXuEXNB/jVijid5Q9CLn/rFTDRwS/cR
5GPOfs0WEugO9EM419DlnWPU9xamugneCY9m2LQIQXEwHEk5OZ5yItD7icNBMVZz
WRxYZeuu/5gsBa21q4sRF6oFvnHCl2QGuBMlgDOfiwLYnapZQTYHEVyF0+a5cHyw
7lzl7oS//828RIfUnr8FXgLHkwLvqscGXd/VX36GkvPWhDulPOSEy97O0Abn/Z7a
8Z7hmYefzd2E3RlyIlfi0u8/BPpnvi2ma2yEi+7O6DX6dKjJOLSn9YS1b6l7wD6l
28zv780v6s+vQHaZtSEXIt/LJ2xj/TZzKKJ0iJHEVrUOFHKtBEBivAj0DIdXqN4r
9x4wvxQfmvRYdKcP6owJQSZUVc0ZePffYQKKcGg1PzlwCFY7nJ84ctI/Y6SsB/t3
6YvlbLllQCOfF1JtkgeRPdvrHh5v+w2zfAWynRm8m/UHr1I5tW/YBICoFdbhI+zs
F702fh0VHxesWuSdXw/BZQ4IlZ5cWVRReuRUe6je2rNA86a+4FOPWOtnahnmK9Aq
yE61SkcDJnzGH5E6fhNEa1DhEWOsN0aTdUDTLLicdTIZExj6UqJWKv9YId/GZwQ0
1GuASM1OjCLU+4F3cbFjd0nocOzAxkPjMXfhIQKgLR0zXCIy5bUZevPGcM4RUBey
Ub5mnqZYfOEM8PH2RobakCzVRa68+Nswv5YudswgOcCPdXD2SyQpl57ja1aNgZr8
GXXczHngteiJ1BZnD9YEsh8W1YI1IM/hXvkoW+RmN1whXEm0GjtDg3klFD15EKvC
RPz1Jn+yVnChuyGriUtmpaffTHnuIX15hMRYqr5kEFiGXhHS9ZtGMH89jxUxEx3O
vFxeFu6DVk5VIsLgO4KwxZbWusP9nxZ0S5D4eYhDOI18nCI/uAhI0AMB82n+v8dc
1BJJcAlGIMdt5PP3+wrtUJT/d2mz7d8+6nowP5w76YKtj7Eto+CEEfXJI6+vt/F5
y8+wUosPwuwRonggziC6gUSwqiLHyRCMzZKcImJ25n2DCN87HJUBKCniZ8BjQ4ns
abH2eCfMxCbBlwZdViRxdEkvuPte46TNUNdnuULnPrNNbKtkSH3tx9Oqe2vwlX5W
qZy64U02fDL8BQ5x6AA+Pwlw4Dahm/WpJiYe+mnVUaNf0rYUCio0WMjJOpfnBXck
MlT1VVrk7lH5uxR75iCFoqLQKMOM/ld6wCtoLsmXroL8e0jc3x0DNxz8nZMsudxr
selI2iGSaDr3PV4N1sweTJn24NWlVlnzE1SDa3NpZKXKeutEFEehEDM4XhR53y4T
YopoTqnneXnOfUax6R7aWVNcbzhCYxreIrBETehyAOac9gEz6GnlmaBOKmCWUe4M
13llh3C4ppnrElilQjgIf0b77dAmDqjOMDR2etJ/Kr6vc+Wes7oY36+L1NSeC9ES
/4/1mnsxRrTaNdRqr7UgRQxaa3hWJA+9utzuDEZw5ZdM7DjdwjyUBZlgp0hYkqI8
WF1mP7yuGhKF+UkCEMaIh66lCVhuNjmdy5bg9PHHqOWVNUlQzpLQKz5UjqJUIAc8
NImid2h1dc1znwBoI6Qkp1veHwxh+RlnCgJjittAoteuFLmisTRHgoFlDHcxnytB
GLZzKq7slDEWPgltVNRt26cdE56/XQrBXOFix0HxP1gKaGzG1j8iaRiWD+i7MQRo
UuqDfIB2M+qypivWqKgrSjg97/saUTq/TI/ECpsGdGz03bOul60M+pmLoqXWNbrj
Bu3UmPWKD1BcDpRJeHYj5Vr3oupqTSceXSzRfRNKu1jrRntARmvg2Qe1Hzph0Pki
FKhzdEYI1zhc3iov7Nlvu/xYIQMMrwmbFR7W2NJxLEOVYpZwxM80Zrze6Se3AVgZ
Glvp96vk8bOWKEu8GJbqfx4V8Etw9l2B6z008Zis7/msuDBXE6Jm0LWFfp5tbdB0
p8RTbjgB3updIRpE2ZhfJmLRtteuQs/uyz7XHWsJwYtwmVdRdmYde3lzf9AWcMRZ
eaLByvRxMC1BdP4oZJLGPfVOdtRblEcW0/kMEgHRpyUeHE3dofTSu4yYqixQb6LF
NZFzRylKjicEHSino1VmMw+mrx22uL2YNvB5FH+Jo2UyuFp8MmvYej2OIvdkGYko
1C9U32nhu/P9GWo74Po+P4o6f9ydR61lTmatkw7LR7ulhQemt9xbAvylQMdaxHs3
IQd4iwKbuG88/P8oC0AkRk8ZUkiScBOpx9WJNlDotBeZMUx9p493uvsoH3elcWJU
csMa7qMcw3pJvM2Ljt6aBDF83ejys+GIZv2QkX21fRWigCNOg0c4HsVaNsQ86IpG
ViV2Q1hnukWlcm0Zr8JZU0wuscxBGF0KpHWTnl7KesxTg+w9MloIu5svTQOAjOZc
C0K4xwKcysiALYCHo4tKbbA6tw3mUysMxPZESOiJIMA73wZW5kVuzZ7Z0bedSZN5
oonsMEIIdNExgMB8OkgW2nRJhxodQExYMhugh5kkxNaesdUBO/+SuLF/nKdTbr31
iEt9ETEVPiT2PvwM4RF2iWqLx+gKLZUjRzklZSA8Gagrm2kHH/S7JQEUwKkian/F
VQv/azYZ3QlxkAyotZyY5xYLedPEMFXwT1sSgc+Zokor+tm36vz6MPCrK6gEjPwh
XMLZaO/9sMzbi5ysQ8MMFjDgNDmkyAnpVdGbq0kkiepNwpovLh9qOuyIc5x5m7L8
UkwecO04d1WFG2ZYUHFA/URYipFHNDgiCBWbedfMcznp7qE9xLZhD1SCKQyg04Yl
DgHZHII4E1LV3WqLwcf8hEu6NlfD5M3+0ucD03zUknKHYzUlwK3tt41JJ3GgGZyv
sjK6ADRKHI5bBaF/Mq+4v8EOBUMXGynS77weNZacQFapi30tieDLnlXYB6FD4j6b
2c4AiicMU3kdhUpZW18VW/kIDFAV93fwXTS6GmUS0VoAU2q97P3OXLk2OMBIvVMt
bQ8fiwwPWvh7pzPj1rfRA4amZAbCCSGEFo8iA2SpqGBi/S5bUwOYGspsecEAQLbB
0I9zXiFciwErHNV9OUuw/Kezbo9nOeaNb0Z8AQhuPHZStkd4LxSnSXaxwWH3L+4j
ztZT5Q4/oMEgpDoK/WpZgbqO6uV2nCiO3w+yiXmiDDkm1eSxqMgJFCgY+ACqzTCw
OqCpHFtbfRQSx9Z18QWAuviDGJwJWG9YxmZQoto1CEntrxhBcHADV7KV568m5CM2
/EjN26F2tbetrNRzU/Oe7PaC7FWLHwkZAK+8fNYoQdxHLcad3N3DsfQ8ZKLi/sTk
CCCkSzo7z5Q1SMR6hCQLG7pPoOnqaCOCHahmabqmZwmNq8HB+Opi+e1fwkbgmws9
xc7V6lHxikHp7thEPWOfNgLsch7Q6YueMQRD1OYCbvTso8eShZQiSWP2H6l1SCwp
ZIZXVT6fCVsQBL4xls0ngtTfAZISo45Yaai44lv1djcIDlG+ZM7YokH/V6s72flO
egkdnxmUSaVtt1rXND56FgdVvaZKZ1LXSQkpfFWv47Ug4D00y0lcfbpdYkndwjKA
EpjpjBbRNph9ZuiPyifMsp42cPHeXhgbf97x+1TYUpj5UQOmB2k0lYsGwv9LmGR9
`protect END_PROTECTED
