`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SkXzPeb7RIU2AUEiWBi4EXlUFAiX9YWi9ucwXHCAE4QUmFnkWvNmb15bdjDK15zC
sa3jQhkaEK/M8IiP2N/c0PTrh25rjZoh4PQAky1mIZDu3XCc+E6aw3IrTo7JdgQA
tEwkoAqdOROGrYEHX33MNorbIrSFmPdEmT5RY/wCzDIJZ3u1o3UzbwjE/Eai0rJA
+WtALdLNrdahZxDbiqV8+OBcgy+UmAKjRyChHfMKOw2P6efxsN3w51InWMH8Ib2w
4qNbccOL+ZbYTjsZbq3bRxpXzTz2/L8Y29kv8j0B2v0ja1rlOQG4KGtgsg696sMQ
4QF/YbM+cZoHGWPMuHPsFrFVWAjEO/CeVQbgsAJHUHryuoRLh6zvFvvCEu3HzSfm
iR/Qqv7u4hUEIvigV5jtsoCJ+QaXtREwRJ5uAwk86a2VddamMNed5cerZWBV9Hlb
YVwJc7meZF/pco2vm6NMtzEOMxxYX/jS6dAQgzGXgqDS56lREoJUXs+67STC0I/Y
ZTG+tdEYaSw2MfqxwMSANKIW0HCeta1KuyjtUYu0oYD5EfBcoE09KpzRcMuoHZ3J
yhYK4REwK791j6MAwPi5YiTjJ4CwvvCZ6VMct6D/u4R0S3fj0geYtgEYjm6aRqqU
`protect END_PROTECTED
