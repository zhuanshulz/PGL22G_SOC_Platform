`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9PNSxqmckSQEY5xMd9a0Y604cHV+l324Mspa45l1lvOT5fSLm/6KPVY58xen9mlm
9P2tG0t5P/9Mz6N24EA0rlVPO1jSTG3oRIy1eogUBVcPTEb2LDkjdgjb27RsxqH9
NBv9MSjlQYzLCCuOpBg7WOXilYefGAto0g1kqyn0nYiCxWMJDUIhXWy/sBJI1AYj
BuqdGlqO5y0Y+YNUBTM2AIrvNvrHaRfLfTjEWWZw0LDTsT8HHSgg1JbQJuVLIKHO
dvJuiEHmWxiGVh4I1lacI+Uci/t/+W0RAhFn60KUGvbusKayTW/sl+H15uF+Voh5
7jimH9E4uw+barpMMT3PAesMWbXCXbHYJcz5/EIMJ3RoFxLxEJQkbaWacrIS5YM6
vqf8bMGORV66752NJ6QTRzAJU/YIJJ2+WhX1fMj6M5F9LvG4lbOW4v9zWdBPzhcD
qDpznx2XzwTl701DBBj9+RZ+DaZkKJdY3aH6DYRag+N9peTkAnLmaXfHQzhZE1Ng
083KYnqx8s/jxMaSToRAqkXBDedjnPvN4JpajCNrpgnmYnKQ9TA5bMukq3lauOVi
iNWLFNzkaUo0aHVfFttbx11wxgevJ5oM5jvMbz2ilP275xZy61mkKoaNATtuMGmK
EdwuwtTaTRvc2WDqBWFTs15bMk8orIcYQA5GrBfWDdabehBGob/lyiTTmRsfKuJr
TNJQ3UuDWlzsh+OC5TMdJ2Y0uyiXB5u16K7WpgcUMVA=
`protect END_PROTECTED
