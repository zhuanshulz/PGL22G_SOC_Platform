`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
42I9dHxYBAfFmmDH55aM+4BiwIX7RwJNo9bIArN6a6f/5i3id2JqwinCatvHKblx
vyayRhHSz3/UqwtVR8GKDFyeavrdNEBRS1Wt0zN27lUz5a8Ll9LJ0PM7vsez1YS0
lEG+D6Eo9ftMkW9U6Lk0NPqQoqqzOripLcO1oRWzyH0C1UFdBtCnRxY7kh8FIony
St29+l0ZU3yqWO58iVMBkOchGSBjjuSYOhG540X3Mo7wwMVNDD4hzJSc6xjiQJ72
bgLdoMfNt0+MD4B1w4PLsWNtQjs61DRI4NwO12Fe60Js1GzFDEN1bPwk/oFHrMky
V3E4P0R9dANiuliYgAWqkneAXeHDwDRBC81Da2QK/rvAvBDFM4lEGSZBLD3dv5AR
hyZAcUbIyKKoDKJP4w99AJixtbtjzrZpAcPF40Kh3FkcjW08hfS+LUlRMWYlmK0Z
TuBo1UdJ44YAmVDXJfzt3rDj+Q1aB5sWU/fjxaTuVluIhLFw1x0R5ah0ILEY8GYe
MBZtn2+cigYkRvGE9bk1/WdrjYWjGQjPsVdOZVr3OphQbh1yXwY2UnxFswYx4zBZ
7Sk5C+T1Cag28OZ+1lvWmzux7eZf2ijIP/SU2NfPtL3p/ZWPG/d/WxOT+7inGi55
RMQI3oUqeqJclaWVePjvl5GMVXedrj3tJ4+QIHz81Zsn3DUUdGNzrdtTUdk8rjad
ycwPsasIGNxu7O7ThT5vcymc7tsGRJtMd6dAxthfjzCdXrM+arR2ZIM7i46917cc
NYCGmij7/zUUU3O7529rgA==
`protect END_PROTECTED
