`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e0rDMswDAdCnar60SLc+SKz1hljNFuTHg0Orp24XQgMZQjD95FfGTqUFYflJEMRj
DfQYOrMxKugvuPsFkONDyjrxviA+FdfP+6QMHIVOeL4//gmxZSzoclNmub6grwZW
rLBGtrZhX2hgfNsBt6Af7h5bscU24kmuQ5i0eLpLy15gr0054rXOqsQFOCPFvc9T
L8EPILyNDdBb/KmRq20UGOdPQrPzOyyGt6PcKJsr+GlDHoXebHnXxDPn/U93c6jI
6EDtI3X46OazHLn3XKN6ml0fzOrGhTLoJmkDnRKoIlf3XAUjg7hWn//5+CRhMpjZ
hbbez/+zQ6Xs/BKaEjsLQ1wzVKF3RJLlX3sD1kO5I4/rfwbbxEyXn1zxiMtVIBZe
j/yhMKY0jXbpp6gpjgdyY/mV8u0NzfFbWl7MSxOnMD0L6Q1oED6L1GM26WQduo3s
P6frKZst520pyGbhSXGZ8NkdUyqe2GjMWl5JtPtG1PTqXXf+J7nv6lYzigExN63D
7qnu3xHkvTAGaSm/qs5DUJPlxC3Qt4Lm5gwT9Hsn1WJ+Mwv5hCcVzBL2hbFYI77r
Q1QvqBRgvJLwqCld5k+nqL9bIECLpPuTpAIDiGDdx1e1gUcCMU7qb2AUL2RLTuHe
9Q5Woesqy8ROllsPO7stkAAHg352FI3RsgPfsNemiNMPmnJNBLTnRBEqPyIbT1Dn
PPmp7tXvA2s/E3Ypw91SUx144pBmz9+BGvVFdHhEpuiWs6HEHYYbQ7mp7vFsbCjG
NHbst84P+FvTy138FIqaQm+imqUQVrfKQp4MG8VlaJVNustxIynxT9o76pGV2YAd
IH2PgWfDEW7tcSclLYa/Y4UshUCAE/pcYgUah1A7/pIMvfzVH22IFuVdn6UonL+O
2MJzHybGLidJby+BO7PC3eY3X4nJtiReScno3huCPN3ABHriSQ4vf2sc57yzIhAM
B3fG2swl13w56AGmvOiR3wRZSF1pmg0sSw/2iPMq8JtifwWPN0Plo5CsdAmVGhLO
NOhAJvBKEc+FfrmWbd5zrTjgCNy/sPhYsUrAucJDHOLdB5xFddmTk27Rz8m1PfwX
+rsO1fDZ4I/hOte/6/7pMQvBIO9LbADJ/wLATf3qCN+5ORT/K1gFUEH99eoSUqcB
S2akrZdWseEp4gMUK+awqbYhDLG94qZYTkYRVoAJs2NXcIJnxnZEvQ7Iuo5VO9Dz
F2c3jQtQaF/5PG2MsisoWAd3I8YLm8EejmVLutSEf1Tr3W+Xvoa628drvGtE40TY
LumVOI58XJ2NiKL1NYCGhvrQ34jBChl1TJaCJ3NhcmY=
`protect END_PROTECTED
