`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BNcrviJDNjjiGVo/yRLtsjuLYvxxbWHJrGjREBvcwbOBfPotZddCBmmd4L1ZJ4oB
W8leKAKTEjan+9iUdkoKpMCheHQ8MEFhLEf2hhc+45T/Rz+lHDEP3s7/aZ/+byf4
MazOzi3F9FnxVaX0/ER/YMlilQ+TUCBPC4lzUesdr005MxJ7m/cA1OT9wuRI80Ka
Xl80c2dwjqkt4NqCZ184rBx7GKs+OUMYJAaFgbpEPlfEsVM8sWHioqzhz89y/pY7
jzAcTgwfeKa1pY5AYR/OmQ==
`protect END_PROTECTED
