`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mY3IsdbSSqSK/nXmcdvFG4gNHRHIydQES7mDga+by8G4w2ngACSp1YReDuplGGF1
j/N0cRCepTu/5ICDpgdl89AFAstXntkYwOHTixM8AnOnJ8i9RJTv/iBT6peaaFOJ
4JY4kxCB91xUL1yoec6iazVgmdukiDLh9lEVp6QgduIqDSoFEnVCsJ32uFZJbLkN
kqB+J8Eov/8lF94qybJtWxduc9Dqzym+YfrX1nUqcx8NhZJvNpl68LZdhUmeVYHX
SmMuYVb6POZ4W/HDJUeSUhjJeny6aM045YEQR6w0UqzfZUm0AI30rbCBrl1owLPF
B6E0nahBqzcKmQa7IHaEEiFsVI8N1zChMimG5vrH7N8jhwyGFYwnWEWLGYZfNACB
1AoX1j/8QsP0vkkBTrmS7nBFOJTgqA4XJEqLywvn63vN3vYTxLmqNt+pBdOP2OIi
wPP6q2zNkhTENRWEPH28JwOlaU0Os2nKXGb2sJS7ciKqxEd0m382+9Q1zc9qsKr1
vToGzQW7FDOVJQqrNcufxcYdTy1Sl48KQfjePvUlES/WJpdBNpM/eJssd/FbzOdt
7Ywhshr2NHRtR5eUvpsch98AJS5ngELJ9FDVaGZaYsZbG8cemZsODsFcqKJox4Qn
C8oRtmMHbZW2R5ls+vSrGgFXO5ZXFEddWE2mV+lXk3jzpr7jj5VohKUIGe4Pv3d7
4ZA3CP9aJv3/LiSmAi6hN3umfpz8zLWk2znB4tzipXbgaDQ/x0Rsn8l8itJPEOoN
LBJTa96BSItKBoeoqoia1wVzkaFV3HYD64M9Jp0wOV2SqBH24T9LQNivx5ila7Ru
zsgw2r+10OvCftnoIYvJS+uGvr3Sc7rwbfEpwTXhtKZp5GNfkgGhjq5A4cyGCPQu
Dge5WIHg0s8vubaRBsnZQtsoGIn6wL1+5OGhkDORW392lKwN+1GJuY5mHFtx6ZXJ
QCLJPmrdK3gBx1zAF+ZhSYvYs4xn/de7hNYpdmjTeS6FR/TQjycTpPGtOVHM8DzU
1NEdq9/6ur+Yn10x/I5ZK4+1xOMerUnq+9sqXlyRoFWGLPjYgqoddBfg/nvJDV44
tqhJws1dANzva8fgtQm9ufDso2QgvLyavACKb73YSX+ev4BykvAZ7LCceyFDXqAk
biESruY8JkvTEsAhB5koYr4HiDVk6GN+cosAmc49k1ZVnCowuuDHrTXbBv2agvEm
KC6NGFcmggEbKXDf1AGjszcGmnl1RbW2S0DfBF7Hj1Oe94NQcjmO3NixvruAr+6y
GudLyaDi9jxmPhvHD57ZJOjtGvFQMyavAZ/34Kgf7j4dStq/A9e97otr+9zn9kP3
eZc66Zo2Fu401x3ML2fpnLL0zKbIVDuuz2G8d2Gyto9TT12gPTdBwB06DdiE77KT
Q2XX9MIHZ6At0DJS+8TnM5zgdh0uYX+TYiFEu7/fLEWl933nFmyXybpVZaNIEsPj
LYcJSCAPXDdaioUpcdI0lkaLcnUkED5hzWVXoGpZLWU0FI7Gp85nFiCg6MYDK5rB
B6GknfSJJsPxjosf59xvPM0QgLDyiPkLqoHGUOs38jbTsxjnidW2Bkg7o/6d0m82
ktFk7LMnMDycwy2R0lMDQhHpMeU82pohIzlsw9/+K11L7lkxg0B8HxEZuAnmCU05
`protect END_PROTECTED
