`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lwwIt9vZNO8UXx8BXcO7PVr80Rpzr5nutUAPVdUw/oWrNpvDsz6B4C8yjY1Ew+pi
oNLAAmEn9XnwR9Jz7Ls3u1qNXflseINW9nb/F/3NuBXjaOZlk2B1EiQw4JRY3Wj+
zwsqxmaVwKvGsHFZS1tzQQi51suLpGNrJXDb7oWZ0vc8JYGTNX6zh92Wa3/DOMqf
r+ePJl2De7V4MyVr4tOTWYX+46799E/YYJ4IV8z3ubYzXbGcjMyIziocdKTV8cmn
Pt62ea9zWqDQI7JEdaXJrMXJCtaaEIOkYA47qbpRlP+6kb/dDs7gcSNZTrS9AAV6
gQi7Zd4E1vl+lbKv1r2Ugvp970DEXwwPxIGU4FuEj2GrnFagxlRLOy6plbrDpHU7
mOep+O4l1OvUhUHXPjBnDzwQUdg961F52EUmLOaUvjjk40eNHiT97Xd5C3RCQnaI
qCVjJ77NsTQgwJGv3a5kQun1bjCnaJH05pePuVyY9wTPsd1iNfAEj92va+jaTapl
sadsMO5G6WpZTLYKn0TJQMIo2fxIJcwBtPkbyKQ81budLNQQ8kzFcUsyI4PPNPR3
rDD2ZW1Rlg5WWl9AVT0Q0QmDlGZZbYFnfBCTZU3pBNTRIeboXQumuPa46sDy3Rab
tMuKFxu03wZBAVqi1IOXBJp0vUOzPCagxsUZhhwChYx7dA208lqxHTOTLvgv/G5N
dZG+l3hcxTfiuhQrNYyc4xw+Dy2rcbnBostwQoaQHandE2lOX7+rDfCtKZXxjUYE
MzFfgsV4KfqlDyLSPwDvaJONl6RgpBfyDVi2HVL7j9+l++PfOpI0jNh2ytktZZ0M
XE4AojeLxDkp5rqt3ahLUhln0qW74bAu4P9Tsw7AqJZh/c+QCkd++aOLob0/zItn
9DWTkDpfqWv0lB4Y6h+V98xzt0Zg+vYRJgRCYUjSM1AevM0+1UThseofSQ3yWSBN
YRBwq+p5592CXj51L/O1yYvZlPSXyLX8fqJ2p9CgUqo6PNobWstzwHiAz89Fy+aW
JwQJJjoXzRx1FnIqktiBHAH3UjwhyAH+xOuaD5SxOY7vhkdNIFePoz+Q8ZxdneI6
GU56jmkMFXhi3KY0ZwgY7gN99cLXS9eRIgdg1CUtlu9LCzsFicCDiKpVqa1GR11a
V58X+73E9AXiDaIMM0w/idT6xKuZaUTPKUPOuICYVodVB0ZtCTv/AJyeGSg28h2A
SCS2vKJLUJfnE1DjMDl8XDybpQLZv7OHLGAAkCb27UsXojO2mA2QeZu56vOEZzzt
5AeGdvA/x4ouA0USdqC4yAxPJrBdOHMBGxPb4+nbTL/IFps6QmuFuQAOFgZRVoS+
db5dZ5COm38rjsuGZqP1t49brPWcymN+zhRXi1wVEDZ02ehPNMjSVzlKvC/kZ69m
L1AAxMiD1L3VBI3ZrCTOQrq1lErjld1LvpqNnrz0a2UpQceJzaCdg8ziwX6m38co
AitTSgZQ/GTnEnH3BT4aOhgQU2RwLBuNltQyYAEbadA7RAy3atQGN05ZVBFGrcBR
nCuu/qSKq6IhzYoeAw64ays4sYk59BWqgJeYjilzH0KGUCTCyn3J/828oaGkybDL
in1/tEy2Puecc4HEmHY7hcmJCxNtVAMOeLv0YBKIW+2Ef2YLYdEgE4Cv/MEgHIHr
AP/98n6PbhjOXnioaB5S9gbaz1hT+RLZZYQeeYeMW3Utz/yUlqFGlFlAKPx0HnIG
AR1uUNiNnkBrzlTXTXNzualbCH/9jt4vD+wL66EOHNCJA3IESScAyg7X4hDm6R6k
QRexQR8/0gHNp8Mrl8E5VLXvLVYlylWW09azTXo1nQOOD2ci+vX/H+3M/RIRozE5
Hc5IgYo0dhs+6ieZtcN8y7n/M4sHvKbm6FeF+Mcglw6ZCUKNmfgS6OAz3chMM6/M
bQY5gADMWlJ4SqJV+OkgOhdO19UJN2oGBxxlcgozS50eDLYh0OKGMUQLEEsfAaHg
DfHEsyprglWi+KVKzW/OpCd6Zmb4/1NH3ueQgZPfyYMZ2JwqtxEnMlCg9eP7WkB+
TIeTYIxdxhvdpC85/KKc9moGZn4n4spXq46fYqJ+MT5vWb4Hsaehh+3v07BoPro2
U7B9a/08F3bwPm9n808qPbonxcsPU49dzx02zLVg3b2JvI+COUM7ddw1iizhyGbJ
uVsD7T+aYsqD1XcLo9+XsjulqsieeXMMnYzJA+m0r6XgJNZWOYb4VA13ESZLry1p
33GaJDj+nJb8LE9rUxI/ufk2CyFRL50IIfP4TSOsbP6TwL2WvbYizcRzPcd0ET3F
oXCSN/k5Op7fZwr+9/RQt5ZKDHyqD6ZIIzjsESGY5gUcgVomRtLk8SL/CI1cXQeJ
N/XTYjh3G2FSscZl+DzhImYtFNPGQcadbBkdp0gR8oZ7SGNWuGhafkSK2LBF3Ot6
0YazKAYPdbVPGRbiqOeHhrVMWi8cZAxrBYIVce4Sh8YRCqK2G47txG/P/fBpZSdf
DndeCAOqhAK18Ar7tp6eRKuYQOTog+w8pPj/t8IXSP3AsnFdajruz/mQejTp4Hqt
E7J+iZYix9hYpucW7jIl2KaPSNDjEOfFTZLXMM/3CktOeySPOv71opivsW0jg/8n
RGWJfqCmHvFankYF8f3gkus0Bkx7aM9OuAeuvcNG9pNogd1NTN3MVcz4NJIw+faL
umiTXOBpZ86tr09PxKWP9VdPku0PYrtT1Wfyo26cVWVM/V5A9+AlyUwh8sn39uWb
DY+xP/kH+M2Y0axeY8u3eIxB3HNYtn4j/RDt5octfHI7SLcBxgGdNEqfpBN7wBOW
edKkBCarDadEi/SlHPr3SCKTTDAt0n2XUC0BFIPa4XggTbHj+NONrz8zTDdGg74x
xg9npk5SUcCsNlVRq9arPOG66rKxDgfwaV7Dyi4L6R+zAi21hUEvMhEia1+l/LLZ
8V8QEd4+hJAqTkHbyN1PqmZFE9LpG6EEDxYvk4SRx5oSdLuLv8YZ5iWxEL6+p1kO
EOR+2kel7BYqGR+Zccq8KnBxCD71kdeBQ/mQXj5xyTjpcxH9uQKk/n/kpX2oSWnT
bV9UrzG+NqlYEb7w00YcGlygoitlBkTVkoM2T7hS+5Dngvkc22QJrihnQL99qotB
1EOWULXB2pohg+oJiUJmWzy8kBXHQPIAFAzdkpKK8xNjDUDN/vgWe4LOCNV3slo1
0dRRo3hSgih5ksQpQ3tGmQ//nGB1mAt5vop2nJpEhgpQ7P7YtpB74N1tcbWm33TM
jy8e8UJdYbeGca5FUHVWG5o9LrerSvEMG9znWH054sX7Akge5VnmrCJW7yyHa9zo
PZPWR+zgkynu5d0GP3GXwH2r3jVncksSckaCoduYacy0X9n4l8mCdoiFr8ovOAMG
AayyNaZjFmvrA6SO/b5Fk7KdFysgGNz9EHchlcxj9eXDiTong+tashot8K0fMJ/m
kRsUrb8GV/WeVqsQ4YPrL/LWOF5EJ17KMu4n2Q76ZiU5oFzIuNtPQGW9MTWAy0EN
RCZIMRR9bYamg6JHVsjQOVvmvzh6Pz79uxZKQTG65lKW2oyVtVUGRmCI5pPVjc33
MBmXkzfd8ywKxh3Qvz8LjGTeLSKq0O4m6dLVVezRfwXXO8wXm5sl6IvL6nOxEUmz
c5txay+ZiErOm2egkAaVzLM2vJ4gKDwK/OuP+NcapCzG5mfw5e6t4U1K2G5neCLv
+b4E7yKW27ZuR8ZfTomk9A6ZJs7ktXcYvnp+b6wJNrRlDOt0XOkyoUs/l/x6sFCi
36UfXZp/XFtUHFLNSHgNdYNkHjNdzWaNHs1lMlD6Bba35XFZooWI235vVQfzF+y1
OZQcb6kZNP5R6xExfcPxlNLgnCMcLy1zIQQ/lfHo7jYJ8MLjrfhGc0TxBiRcQWel
XFdKCFE5WdU+4BFU6YDZkPi21RCo5o1hjBJfht0WvefQUt6jAbmqMVU2ntAns26z
hMhxt+zTJJNIEHnF8IsdC4TTFjvH0au1h9aEalAlSg4JVWtk+fgXLHn7ElOo08Jo
0UQ+wBnrCUH22b7qdS/m8+qh/9dk2gaVcIsNpV768dphg3t7hwxm2f9Xx1+aekWB
j6iF7Ej1XBgipSw6z0yTFr6cxOhn1e3KcseKpsjmuhru2Ryg49DtUVwimAbBo7yc
KfeCIBHQ+OOEG8T1IJZSdaij7lahBEBVD5FqYPgtGEQH6qUWgcnv5jHVwNde36t4
B2NneAVGszHlAZA8LbC56m/s+oDWf+fEzDKRqRLswnYHh3l3+5dGexhRosZuld5S
qa3sYAAnlMsTk36SxKeh2pA501bVvYb2iLFC7pv3a7S05qcHyEl79iIfj0mbKRV8
rfuY552cEWMIYPwDyvDYsn4IGzBqfHESZzW5xu0GsJmlfuKHLHhF8ZDbYb3ceUVW
uNpWvJBigoFifIJ9xu8JgbjuX5E9lNt+lZ0FGqGMXQZAbqF6G04810bZsDr85Faq
7nloZBgEcQV3uGlpCQGJRk14kCyvKfpR96ISGFzVkN5uMNqz9BXt5W6v5Ue8SGn7
hcR+0z0M98t7ih77RAvs9oGodF1IH9br3xuAp0TMMpc9ECYgfDHFiplRivTWZZdB
jBNn3z+1zChCiI74OUEZzDCVYRmo23/2BpoG7J1nN7RyJhEo1w2bpcZ3c4aU9hVw
F/wTGfMQWgHE1gPEOjdboaeiPlyzseqFZaSAu2SXd7hkkg4Ynslc6oLWxpuIvvRo
lKOqyTccvwOYBO4M18az0LUIiqSztm3qVZkpMUt7jYVlYO5D0QYsv8SqfTOLqGOW
zhd7zQgpaXH5zSTVdHBRjVpTuEEqPpgjrHM2p3x7BPX5EtXtl0Bw3RsIT7Y0z6WJ
pNiYpZ5tmMnvadKECdr/gjOjzVm55tHZYEx3HeTsEbrxuei0/AQtz0/6sIx9GJ7K
USG27PH5nGP6j1owoL9Lww7AJFpFmaG7A5fYl3z3a4rSCQA5ioffICEgUyr+QIyM
dpegsyZXdJRnchrnKFWqHnKoLB+nsY1AQi+xyYFVE6cAtm9zXdlFVSfF6puQFEOL
o+PSh6gcbQopL2DbQOWwtEuF1QTwddaqenb1r/mBNFf0Vqc/FLcnooeSIQV9fCOR
Dhrt4BPnJj7Q6O5FLFkmD5SVf5rFY8QfxqrsObijdmckWAp5RgKnCmAzYUF/in2j
9FNYA7EhC+rMmjfjSA5Oj94EBQilSB/CVzqh/Qc8tuh1QT19n9I/WHF1FWu7LrbV
LVWJeb1EBvGufeNw7btgX8jsGCFx43Yc4ojjt17Nm+nvMmUifsKkDgwSOc7s+5gQ
dGT1kRDIcJK/1DLttUH9Us4EH7QwP+k+C5i14dEYPp8HQ5cCBXbxlSbrmyCsgdl9
uESpE2YlzFb47NzxrW10e7s52iIWfNP9XjWMx/HFCEBPvmqUMVIEF2c1e/PR6FGl
qMqfRHQ5F2fbhDHAzlrsy4vcL0Q6kKlU5vjAIZkMiOHj9DoG24vqIlt+gpaOvQdP
0DtC+e+QOvxgVnvryk50Oql8mXQf1usxu77IL82xL8iwQuw3OA6qEZVSmLXfBSoq
QM6OMXohZNF+PsuOK8To6wtk9qtgLG9Rmh00Z5G8pz5JD8c76lKchhix5YyN+tmc
BKkvPwYey17YLW8OksNZFj2th8tkSh+BOpny6tjChSVkfkQciEe/tYUjI+yV4ghU
meWjteQP9P0GrYJCJP/Ih+pRN18MXkuyzu1FKRl3N1OszHcDJw82769yDSfubxPd
8xqgai6XzXlZxPj9g22GhHwd59XPfG2VlmQQoQhCJemRSrJLx79LEO8/t6lH4OrI
Ii2OSVM5EMcWrqf+syd81KclNI4cK5y9BMxobH7+vRUeCitR+044jrjCh/fjTJgc
YflqJ7S4iYv2C1LiLgs8tRZYJy/t2FkTLByKV0w0mqA2EDT7tH6w0KY3fgXVvLdt
upXvBj7tn/BBlATdr/sa0Txw2/JaPYAios+gYRKLlBXjzvjG1RUk5+8eu+pc9mn7
L7evvaHpK9Fl4Go1Hooi23JH8QUFPmcU27XXYZky04lJl+OlYLetwHMM1/QrE2xB
Ns7hhSK4k/Xdcu9C5uonfVo4hVEEZykWiEEKj6N/0PRsj8XDx15b+5zgH1nPxfrX
cl/IF+ylPsC+yaD1+oZTXsDX/6518aE2CaoUmtVrRjMHxJ4wYP7cgxASOS1h8S04
6NPfC5oVYJ9r4iP/5ONUeX958QeMBVouSbbfjWYnqrwPb9DcV0rA9g9zGfCp8MXR
8K1oian5okZNXvlQG2Tr0pXEOlsUt8f3NZ7Gp0m4w0x/g8AUEVT9rp73Pj1fDOho
c0A1vg7IOG1lKrQMrNujYajk9YnidcWUdgATzDhF+3KsrA3GaMCtl0pm3v8GYZhd
hpfZXMdrGRmWiJMmTONp63rHDb2hHTTkvhIboH4fdWz2df0ehJNhhRxEssJQdYjg
BT4LfsdETJGZbSAazIcz5osiAJHh+a+OTjcujGTy6P8wCQdlUOub1a8ONyCjrnyE
dNFBnqpWT3dUCObWVEhRkfvcXt75xlWQpczDnZlK0S3eVkViUnIfRqcj3dwXypvp
cYt2t9fYU3TsP3k68z4IG1w22OMGb4id+StV+b9uufhO9cZ43zWsIX8NyjDZ8n26
4mJpJ0wyRsNS/O9L2WyWN35svo2KGitS5NgwHCTXJ2cBV+sumQpEtcF9N2SkVbRX
ZvJb6x+jeNXyvykh5remH6rKBAYWcPn+lANEHNbDObsGxQnfjWw6n3XVAc5lkDZn
DHSraxr2gNO0mWXP+CpS//sP2V6OXR4XNGP1niD5+QWCZTOSLts/0+6J8N2jJc9U
GZ9fnjwFK3g/Fbxv3JM4q8AEVH/GxHr+WsMaAc5mavzHpjl+8dC1ZN3Ymb8w5Rr7
DasYTTNkRwApq6l4UCRgttcpsB7JBQ5GX8hUDGWs6k+o5Qc+NFLfn9zC+pVUvmCF
W4qlNu/szlFJmYqqtf+PVO0jp/iKP54dt1YxcuoFDZ0WDrdedalv/NvDqVdRGB6u
NKsQFoeAfY39SJuX9d603WMOT2wSkfqNaIBUAlVOkctQAlHaj39+Ftr6mUXushBM
EK2Shv6IbPKbeI/7VOeVHP4D+DqGFZqSrvGA4EJ9bRrM2IP88Q+yFxy1i+wRVRwz
YM7AnFHufEuZStbbl7iJO6PMCpy5VdZ1BvVqK7F539e0rvxPSxTmv0ZFnPEphDdk
9MCJRxdiLAchO94dxn5GjW+eT2DhNMw9EMZq3RKVQO+IPIRbb2Quwml8Bk+rssbz
/2d+YSpoyO+f8lnokRk40BuzK4x7UHYSB5fjM4AiGS/PnCQQVPqUT3gWZxhYi0oB
nQCwFQZRXOwtOOx06arrWEl1+FWe4L1pb9CJNFiV/V2/e4GNm4pD7it0H7JMykzS
zPIky7Tt6l1tKixW+hUFKXlMk7o2ZL9M6TL7kRCAtOyZJ0HSTDyzuXN+5accD0Kx
QIoAogpBoJslbSGnyCglmlnK4MFQW3bLj8LUVInykvNRHLIfdB8hhUazjVrrBHQq
sOmfzUnllg6ejdrEw2851hCcePX4VHtS1Fa7ZYTDUn3dXmEHj0SSDdM4WPUebzgw
34pN3LXtsG1Z3qUHO2EZY4wt0sNqcQ5UkOmObVHn4GkuAimmXq6ch1XSb17OZgu3
l+5C+Nwbk+Aik+q5SQhQQZHXpU+nJ/dsqjx/CeFUuzgrGa9cK4bWmPDsMB2ud/ZS
rfH0nA/dltPBhK3kmQZTCMleUO+On4oTKGi8fFtAr69/XpBZG9TKMDv1vh7i5Mlt
VscrEq0OGs5q1tltL6hkI9aDoseBUlKny+sWoEXb3sQVsoKJZPndD4VNrZHUmOb7
g7K11uKojaxJJ7zg9S+TBI6ETU9y+SYkYjI7LccdDRLxNPB7kJxpTizL0g3ycVBS
IGsTomcaQz7XkNsCCONTdAQdlJVnDpYCkAZIBW9oL3hn3yRBCxiTSXc0XWi/mV0s
Y/2UVHcSjVIxixz3+fsxPIRP3rT0Bmf0z6xbYi2pDjrRWT3pOrr8zUuiF1UFHzH0
B/Wnv+jl0efjVAyDmXHdtlSviYO4r1j4s1p+/0wjnX69euY2Hy7om/jDzfwMsKec
a87tmXTu5Ql7YRsxAMeE80Y9gpglKvC1HaLTG3YDezvVX9p0Y3Q86HGDQvUpJyjy
OXlYcL+bERvjFKdKpN1Z9bTNDX+EtvurTBh9lvc2hhQHA+vqWRPsUmIElbHnqOrU
8rRJkwsDODfO+G9vj9+lv5wLaI9kK22wdppk6vS6txJQoWUgInU14VxKh9OpPu7H
jnCuUR98whzm/KWJF+47e8dK8AbjsyGIWW5w8PPSY4LOxTw09Gi95LL4quZGKqrP
e9kQTU6aDVcAEetsT9z2IGmBBPMAfAWI951GlWPFi919rdStd81jePRsD5caeyuh
8Fn5Dnzsl5ou9azY9ClOgiZkHEFs+fEZpEc/stCDZwzMIJeJoZ3WzRPuBczAAyWl
+DHhcv0x6Hh22N281H2FTe9CxDr7DItgsvG39O3QZF50dlBDs5DjnWLAUGJfiQTr
vv8h/CqWaT++eq8d4xSx2G3pFHICJYYiu9RJ2PL6kSLVhJP4r98/kNQGZm12d1JK
PCh/0pG7PY0xgfDGw70Vg/cVEs90xHtbMM9a9NalxHDnuouHrBhZQ9Kk6clgnE70
So/+vm3WZxXP9bSAiRpxep8gh2UY/qkbVlJXMDlIjOmPEPxvc2YhXXYuIC10ZdWt
wfreo6iNcGhu+cAV1CG9Wc2FrapDuclK5nrhvXNu6qBkn2fkGT6l8FUTHsMD9eXb
aE1+gfrwF6U8ycQTV6Bj8eU7/VJdcrZ73+Zb9S1CeHKu9gC2eTNjBb0qNnilBW00
9k402DVntGwCxc175kj2czNPWf2/aTSEUq111eGj8rycuN0zhSWw9JlYFwUGNegs
DBdA40ZlfhPHqpN9ay7RF9Q7RHRf8EBYKV0rlV6nB/l2OcUSmClbAJuAzA8zdeM7
fiuK2yUb061NFtgyLcCuhF6N5viTTkJoX1YmvPMswpr42d5bfNrAo22gxoL2viN1
YmTfqsfDNzAhslfziicvovYCiUsejvDirDNoU+yi2K+oN7DnPYwrG+rrSahOqg7Z
5rvzygnqZKe4qMUZLQ50v3isM577IbsiP6mbey9Rh1v1CZUWXYH0a1jTPcP6DzMf
JaHCm10J1RU/eJ/ZSYkQuNMLFR+QPrSiGGxjEmCpAwi4EoMNpuV0gmOs020BMmL3
VHZOTXuXMyCj5+GuSTwBjnckm5PBuixtxV+XOHH+eA/JaumFTYRexhweZ+pv2U29
Yz2UmGx1/G+0x3kNfJdpZLrygYhmlHy7rlB7nTxHFZfBoMo6aOQE5Dq6W+EhKEXg
WJRprXI4FF1E7Xfds0Enj7PJQYHP5ZgtayTBN1gDp40QI+7TLZjfvdyjIxE0HwDO
hJxPJLJwJsYp2lxh4l3NsONk1Wl58UrIXRPI5LUQZ5CfOeAi63ZLhSfuRJdXxqNL
MQdGVobh3wLGbLRLYu+gnb/2NNwI+MyGtCC8VjvN94THq3xRtDE61+okegsSmSkj
D125STo9UWVtIpSB5iVd6pO4nKlfH0wS/FnDXCaYvejzljnff1UwWD/X89URYFo6
mGcJwSpR4DwyI4hEwtRK7sqBEBAKR2l6CFd5mT3YIVSqeGF8tGnKW8m0Vrmfuw6e
8zuDHi4c22vaxZhO64AnMgbZe6Pzldh4alPpCcJlHVQ2FBH63XZEN378bUjsefy8
mdYbYYc1ebvMSs9RXkf3gRxseWoLYWl8l/alHSLbapQscbjfLyqCHLb1paq2X6lg
k8FMKmoemUe3f/TdJeO89cUNDDweyhkRHp9IqYWdFP5uGfWufPCD9x1KaWdV8ist
GWA/Mu7wKB43euu9zgu5M74zazvdwQMZKOALMEy9WkjLCB87QaOWaXSlMlgMfc+f
Qc2UyVWuxacO5x/QcVGwQ2dZO+y9j2P8ibczSAw7wrrfrb4poCp6rAmYP+uu2Ex+
c9GyNCL+3TVVob9DOAVLhcb49cPeT3Sk6aGTXJmW3NIqa6vUjsOJFZ1M3YaXRLxx
UgYCt6tCca46uCaqsEwihbAiKXNXVNQqQ47Fh/JhavFXfldQlKP7hssgdhh0Y0Do
QJ5SLjSaJIzdx5iryIYgQqmFQfv1zBhaxx1za0g0wnWbYDB4jFtggCHESTnx58/O
KTkxrP/fzewwChCubft0lIDko1QoKFDwK7xFz52CCnar9je0pH0LlTUwOW4ueGdI
4BPeGJqdy69KQtUcBNtpByTNqk61/vYJlMyiS+TTQDMGw5OyoCM97C7IRnL+Dvts
/QQsUA8iGUZQAchMUZohg5ZWDT6b+aGBiXYG0O0UjDBTqG1fmxRTKNnZNk+BJky+
7SjSndmn+Qqu5zT2aTCJKCDw3XCoNTpWC7xjAV7Mt7J8RGMR3J+j2/qpIpixO462
IRB9Mk7oQtVUScZkunHYnYyU7oUzVEkV3VUGzW5Uph6gU8n/avwZoDhyv2cXTNkd
dqvZX93YOkQduPghQ9s7URQXUpuM6XGTvAcz6v7vS7xLoquktJu1TNvKOLRXHuFE
mZO4Iz8VcRbkoH/Hlm9YOI5X0VhvEJKaScpvwToyZXPAsE2anovj4anoxk1v87aP
wzNjZtF4y+GEoMOZKsbMth1KEWPnXByrAMAk/2CRapElzhK7RoWngCBCsttDYW0Q
oBBgDKJ/ztZpjVcvmWkaskoyK/wM0tmd3X/Y0hoTKJ7Mc8+9pYHccElBicagjZe8
5aPuY6WARA2rm5/XPLpwBksLjzI46qq86nKgwMmnRAvqlYKrf1MIFxw1JBowe7GR
EJ/gJkYUABgQHaUQfpdxQ2+PXwh15VN9o+y1mV/86mIk2lcBUYlKWGm+9Uz9pS8O
M9TVN7GgVwro836KsdYycYdJwfsBKd42ogeYuMrSL4jkUG/CAJ3sotvxTkSziAeZ
FdU320iurXCVwNrQi87srE9QfjI3uxn7L9hsRHlNIvU0czZhyUgnLsoBuAcJY254
x9DzOKmJvbpaSwMNGgkq+mYnwLvkKx7CRAnNbTf4xu38EbNN+zrJqLyzSIsyY9bi
hU5eIo+Vf0Rm4LX3vdTYBTKTIQv+9FpyU1g9UNSdTLOO1717QQynXb0wBA1GneFk
Fkh20wQ8QxpG/d1dc2HrN+Yg+0QlWTu2Er1xgyhaAXeFtYKuO0Ep/C+d1ZrWJIjK
zaWHSpGpzGQVzT//Ct05akojWRxwIWh6q6wd4vwE8g5PBcP4p6aMa1ec4YtZM3DE
MMhTJGmJpgIlWw1Ytw/3Fm4fS1GvUEKCnxsoSQGctFr2yW1eUFKk6Nkf0CtvZD6P
JAf7YrUT22Gi0IwDw8bL2IBRgWRPXlGD1d8wLzZd7eM8uyIUREa8M5Tu3zN+3GyU
NKSHFxM1iyGZGZt9YXJAKYeDCtcQr3U4koIET34SegsQpHfYBfEzxnsK3lX6cd/Y
9eXNC8355hAq/6kBHPu2RyMJxrlXEftvDyS4mVTQ3f2AtYs82n3BsVfF+3NKDQrt
GkXP51E9o5nTFpa/mWVuHe1dFMRpMZKkZlfY1+wy5yTdbmpB0R477Wr/t4bqRYIl
XmOETp553U0AS1H4K5e9inzPg/HFFC/WNF2K92XrsGOYgfHYsXNHCt/jKEg5tTAu
Yn1226BTOe11saiALrszNFCdsznKDTAIZpVrBzXp+5tVRAApIBZ7uATjN+8XdLVY
nysKL9oi6I5n2wAvdztcRHLQTcESo4pXPaywtXY+ZcBrwuUIBUJRQnZa61jhL2PS
Tbyt+OTg8MpKOAnTheaco0pPQOB9CDpR7bxjLCuBy4hy2h6Uyrb/EqpH9J3joBNd
VRLuTMr1GcrO3FZXjxY/nRk6gZHSfSYjofF5nn8FxYW8jX3TTSxNsfi/n7O5wATy
JQ+rtDohI42HuzRL+pXvXHYu48eYukvg6xRIDu6PuT7ruTeJ1ARTY6TZ8wdCRsf0
iCDE5YHdgHlIPlnVTBnWmebYPC/iNFWW06MURQbA+XNZVgAM8Ylkq2qzSlLJuhlu
ySeUt6aGlavGJUJ73+LqdP68uiqIMKV9O9HI1O7tCU/RXDxHm2KBr89OqnxKPhi4
2MpGa4gerPSeHyBgVmH4dXZ2tPI3G35PuFac8fmOmqIyYLSxocWWamX/lnetOVqv
hIqySImpkulMFQHAW5KSBEVYHUpQBQ+AGMhshUBrISG48vcW4vqlhw8ius9WzIlG
IyvwmVpo8PrBkEG9YLgwF9xCWiVr6ecH0A2hPpGbJrGLLtDY6mVKkKS9cPdvLcV7
Wv9nvtku7qRfjXt2lKvuyitoR3f0pRDbj4Lqo7D6qe6gVYDJUzA9rHlRC3jQWpI+
94SXF2/6UHFyhBYwm2gojbaI2g9EnAqxtU+ZPP7UmBezSfVtWfT7f5Fx2P+QeQTG
h5OXHmmbUYmo4Ch9HCP1OQRUS1Y0+yeDZAo1+8bnwmZfEIX0UeWQS+8MWNAOlAUJ
efoxgyD2LQfQcCey/Htjivj14PR99qwQfnQKPgsZI8bDEZfLTtcE1e5ccgN3BESf
Wn7xheo2NTUAY8jQSAPCIGMdy4vW9bq6ZCnfRqmi2fC9qK+YTOHg/0NvGmk2dfwI
8xOPYmt3DT91Nk0Un0mBOzVc7owRl+r+JfZ0x5ih7zXt74Plz5fZlgI+FWyEaUyj
He/QCJx44vGC4nI7taPY/fgj6j5B68cwkh5Fwn4bYPLMnj/yg3L9ZiQ4PbuA9PRn
bHfIwMsnCckuGV8SBhTJ+wJ+agoQOMtozVw8sy6Q0NjsxscukJCrz0zm3WV1BAIp
ktKhrcInaDMslxBxV2BmJBWpCrf0kqiQC/YpRDSTzljWDOCI7neBGLZ+1yWIJHcd
sy7KEocyYsEOzYIiBcKJ7rb+UnyYY49l5J6izq1Ts/5soms3pgLGRlgTcUGEgn+K
ml3mZaJL9kv0jmNJdOUPbN9PoUqcZ4xcQlE8Shb79zl2cxVVVL8NmbrRGhQfMVSL
RT20Hd7dx5PGBZtzZublToQNK3CE9vf0A6ljpUwgkQwM9URppbT2gm4oF+7YweVJ
1LTWEzsMXSZFie5pmOYKyftRUcthviNq4TaP779/8gK30BoUfxK6PtxQA/U4Zs3w
7FAd/0b4yiKJPpyF7kVNcpD2Uryn5hy0sLtC778yYj8CqmoNTE+zlsvcDDZTDFOK
OubCmFWn7s5d7gE21NEN+DiHISmtTy3evEdp4xCxlxa4BvXZhdwH1cfc7uWpruyA
FGgkm2BNC3xUoO3KJoFf8h2B4qPPFBdIEMDxsjxPbVo45KC/UvKGfXzrjCqOWlae
U2d0EwNrA9BH5sFbacxpmn+NB0bk+419VvZNbGAcIuSl4hYTXiBR/z/y6ErzB/YR
1aDCR6xCXkC3hqlOumY6aV4ePOnu6Si/a8T5Ysqm1mFgmr0NwA6rELg85MvPizeS
NezEHCNziBq1I5P6mQBzoyPPULJI/9bR0G8thNUWmdk3Uim643Z/sNe6PZiGXu0F
W/1/9lPNFP0FPBt/vsDaMgO5loa+reSEiHhVLK8SXk+zk3vBNlKuxq2aUwYkWEqh
uEP9oxeHfjqSRQtt5QKLVSraWw1P7r5Raqkvi4XucBMlvCDOJqfJZQkS1hevE6MQ
+al0jxEIJyDra1ZFYTpHVoUFh1amluiE9i6GCmWJ6O3nr0vPRPHgG/Lf0/E2xNiE
eBVLPAzkzfIz273TNdc7hGb6owtKaMGYetlbkRVMcxhUANwT02sfUNdibNM/YPVb
Jh0h71lF+pk3ye94tONerIVRCxTCxvSxC5HJnV+Yd7hY1iHIqeT5QKUZ1QeRPNfk
sv9qFmD/vaFSHlMVcMd51nMQvU+g2/Wp0aEt2vYmkxJEtNnB738WNyHuOmLQR9Up
odHawsuyE0LTP3Ur1Tgut0oovGYu/uPJ6764zLhUF2oNZ3AMXpURJc+weamH9DFb
yW3IWV3eNfXquX/S9ZS+Ppsm4a2oS5fS5hEEzBUJ0vqpOwvdnIJ8G3hYf54EbQRs
qnVbl7ZwFuM1zG16RKSxfilFVhQhkoMyK8hZ8qEycl/e5Je62/LZ0i+yOd0U7iwu
Ns9C3NtrxeWdpXV23oyGIFV2bGNwWOE9eteWlwuVk31NBio5RPuVIz6rt8HyDJaa
gfwKp5I0WxhGiNK3o1rhovqjHJorsewH7pXr7dtNRSW8s1f0fLwv1Vru56fYmA71
2662pZDXZ2opZTrP3oWVI+lsTj/fA8ErTwa2ZXJ66HxRAonZ5iORSBA2YoBudPZN
o9ZBjPsRuLV7Mikuu0fOTBwKBncabeSxwduIsmY5y4dawK1w8+Aj87pMOhSzXftt
WGIYB9PnBAQIRnchSiv9w5MOunWrMu6pPWywCNQqCHfoSymfXGEtbvo69J04nlwK
7BbBefbWvypKbqy8mnsFwSm+I3DT8l0jLl59jpuajD5hiYl/pdQUEjgLRwkgNx1l
O67UpA+8qVjmcic81GiSLcuspqZV3QnsDXEJbXHBH96zC5nqsO91uEF4kaDUqfpb
8NOMFcOc2Cvm/gmbTeXek28BuShqTXCYR8Wp1l5vkerdrwDKIDAh4Ev3r2Ea0X5/
VCFHKq83NQv2PoQA45FziLrXQXsAa33yyAaHaorVXzX6wrQzVtic5DZanlnBI7w5
N71AkK1iY+AVIUF/sLxAaEIX4vyvMzku7AFfYqikWHiZkEtoAsDqvrQp/J6Diqx3
94U+w0BhvX9aP5+CZSU3ZZLRQ0k9pfl5C8s278obSiN2D1D7LW+PROXOqViN80Zr
PLRnPOWuy1bbZjUtS2V+o3WtSWCSaUCkJRRPUAkffQI/k3gdbSMAluoDoOxSPHmA
gwbQCQk0YIqwFY29KLwrvmt0AU1Zcgk7POaSrAiLzSHrkoQeJb+gWEzRPAnWZcYk
MEACr8Tt8OXDbPOryLwip7IDublxIzTAH/H898FF535Ze8UGG4wk23WE1eVK4Dkf
DzrP36W479JzrmUqlgXvH4IW2hurfyrud8HsBO6v61pEfhRkeu1HJGEV5OenwAkb
hYXRvq3yRgSdZPi5TqZbALl0yX6nVqAdxppH9JEyyRqMSdEuO3ZYwX+pOX1Klqux
onavza1IHWXEU2DxBpqGSyAXAAHS67ChZws/I9Adxzy/1zH5V36sdfjqLIloPA1L
c2iKzmiw5XuyOqrhefPH/BwwNxeN/M5j0Jop5VSR2TRsWtZN0UmLz3gi3THbOddJ
nMSDXa3UbdU0S/5yeZcZ+a/BSeyD38S/ApZEqHnEu8Yp+c6bDp7aWwjpFOdDNEhm
TKpjpAfeMWE1bs6pfhOcySwH96qOe5luoM7n32oGqewMCwyUm1knHCZCgTMpBAdW
Q48fiJCGiVlOoaZtzNF19urSlD3tzUdLKWjDG0ADaIlndshKQFB+GH83p2MqXivh
l2V4u9d/KK6R1vOorng6U2tFens52AJK6FDIixu11DIzuaKgzd12KvtSrhbtbhL+
Ch2nKsIb1XRcvRqmJWjXeNWh2JqgaaCOz+rWYoM3/EgbOTelfWh5cTONf49r/A81
eq+u9Aw4AGkBU2XpCf4H7ukLn2BvabU7ga91TPDQhdl6FfEGP/zN7/vHZ074SeRd
fmjg8VprnkEQw/hyogzandAWjIjgrs6jOMGfqKtYp7CPZ8MovQM5ItY3IUDi46Et
TBrJPrRzVCvVPt5kRB/+Rv0gXBbBMnu3xdWrnctQt2N1gAGrB9Uvqse1XW7XcqTg
zwGR5L277ct6DYxhCHDldNePQQ5Nm4Si7VwADwqzwgacC1GDxhWUswCkYo4DFwSQ
Wrmv2h1/K/SeLWp3cIf/iFFsmSPdb2ufPJESFE3MhsNJ6Eulgab5nOiprWvnRPvf
IE+ivzrM3J6MnM9r+JMQSKUNASQL5UNT0soLO3e745jqCB0jHa9u2GQyvB3aujaQ
FibvCBSSqB1iziaHtzaFGzAxp1KqTWgNe0vilSpVQTj7VTCiVb0ilhrtmF0NB/sn
NNn5A7f6E7Tm9Rux5MS4VIHo7au8KxrHS3mcpkeNl/JmLe+v0f7dioc/bH/cagZA
rwbaa2PJpOh9PS8zoRq/wmJcykAbwKnj2xEgyUYmlr+4K382VONLGpkfh/k6ACTK
ITz/1acHA/nqPzTIJJAgP6exdlM7W0fYapr651EfQTltCYt17u7SblUm6di0zx5Z
yrJK4a2tZnsEIvBiR22u3PmzFySkysfMxFrlQ5tb7OB/9SumdTHWQQfp0kblqaRZ
4QmCXRZpsYKuYbfQELD8TzkiDJzOs93Pk8C32iRytRtSNt1Uv/b87CyD9cZmJaMw
Qp493opyeebnCNgEHUUI8hawI87LjIAPJItqavcpU+ojH6A+IjQc438IXzxSr54c
SVZsASspNpmHVSPjjvR2HvKWqJu/ExUrYGS83YK6IWfBJzyYqOcJpqSsJPLk1tis
iBBL9dsZiwcBpdjL/+Q0x1eQAFJ0okR27m4pRBP/havw/IFHZC/1M9reIrD5X1Gl
KA+R/0XYtE27EqW24iMZqO/UfWxp1A7zC2l52H2eXa/r+Yv05BAn+jvX/4sZhAdV
bBTQKcozoMIu3feHwwfJDZDgR0RuXub+54XwIvJL/U1iPEja+VcyiTOomJs4ykfB
MWXtjiloZ1ZeYMQaw057cZuqXeAGaPDuhI7Kt2t0XalKX/KIuAVD2nRtLhZNWoWH
gsoCa7G5oFVk05ATEJk1tGMK5gDwrACBOY6R4pIiyXGPVQC5PqXth8o3M64C1sYc
J/180yThmpjBpVqE2PslGJKGnGAY/zFNCu6S0nhaKspa9ww346A5PLmUn4z3i8kx
b465NK+kM0SBpjNAbIZqaGbDxHI/Tk0HU+UAolrDVYSUI7xCa/3ImDssmZunNuTj
fWXxUjFDZQWcDWswJmrUg3As1Yb3qo8UkQDkdfZsuIRw76nsFnQZXOpWG3FyCIJh
bfpG12zDLTQzzwssYlgFrndwiGASrKaS5/25MaD4c9pvfal2h8aH6iRqIkrtMGew
ljVc9wonZEeEQg+oIaWX7jGB+jNxsXw51YkoLkb3L6b7YT27O9wNAqj0iZ/yuULT
mf8podjbmqWs4cYIVA1LU8yqWgS43hZ5431bKOnNeBEIzXogRUc4F1bGNTBgY7qx
TujeQI5YTLKXVPgbAP8D4zzrq3H5FD+pB5EgRHp9MLgINkamhR1QHyYHpClJEjsB
TnV2vtHBSXzoxToorDNZg65zadbviSBdYgXSrpKnoJfd2ckm6xeoNkAMvrq9/235
s54Bk6Rs+RgFjORlm5A5V5sYxcLcLxU8Ry4x2sWOLSf51TMm5bbaEnOioNq4eNtR
fuFh2FDfvPYJvirxF1cpIZLwrE0oCHnbozJQff3y4BEtdEVRcBrg5ne0BXGIE1Lr
JGl5UGOlNmHFhNBS04G+Roy8ew67kS8+uzpc1WIPvt2kRzZnjXLbbOQukXOfZGC7
E63hZDgimfA7XN80nin2BdUg7bSENpKNIfh9GMzO+Qf5YLIVi32UcIh2dCIDumks
dTL6iShLyrnz6QoE86kdG5K7c2sLbWo1CY/qF/+Qosh/SLF+5Ly5hwl3xmPrlxhG
Vbf8raH+4d+EmUpYG6Z9zuEk6DeqS5nA1+siLNS8YABgRN6aphyRdQGhU0JYNY2r
PUeli9aPpNKwkXMXngUvCtfJV4c69d4t3Geq4FSckkK/yr9jNx0K+jQ6xmYhqY+A
btcuD6m0NNSG41b2LfUJOnSmIWlJSEObMijfKP42z+EF3RH0fJSkdT50fC1rxnQg
QZjRay3SGV9vwotVCwmf9g/mrxN4op5jN321fDb7jWDT3wAZt2GtbUeDxYP3ZnFH
mn014kgofxe3mly4IQHIFdmunID4RnDNOILgevMXB+WKCQrLyriy5wN3LSDh3DQx
DYjuHl4qAC/xH6oa2LgjPGM2epIYbs4rSdENJZNtD4i3gvGaS5Z6kE9IMLZAi8Yz
BiVhkE99/MA5XjAAifJhgUG7SyFj+L55qD5VxzT/lJwdi8086LeOjIpuKcI5wspr
NJigzjg2AO9wAwavpUurTO4hxw9FzA9yU3jjeoOZUiAYVM200daiSK0u/7HOADoA
7qQSkti1Qy49vWpZT7AGcA/wJiekl2fi0LfJUKvn9J0yIrInColuwmp8QfnfaSqF
/S6Q3cEFHsRsglu4ikXL8atuADCF3QWQZ2ypLgOjPIT1diaZMn9JYJgTv8R97o95
FUc95CIo0T4Ep7iqHzgv0EK4KXm5ny2w6sD0RKONf1mjH09A9K3euqJg8mgEEDYx
FCD8ZRSW8UYDkwWuVqHu0EVpvuS5yfaCtMFLcOatdEuU8QvhYrimzAFZzYgvKf3X
QcPv5nxQjmLOedBG04zZVFFd+XXUUIO6lSC+p8F8XJztSK9SqUyqv4vZ+Z6tLwWq
FZvysYYbnQr2s7JEVJZAt2thJim1Udi7NbInOpopJ3ekIDFmbBL8xPmd60ndUXuR
CSNL8b3298CK7s9LI10Cc7xHAg4PI7k0SAgCVOXj5bZgJxFiRxXA43DygLthVYwy
JfKW60jkUke04hqvvaY+A5KH8w1akg6dfeZBRV49swgeuJ29OmR6YvLLI4ZriOAq
6T8XHuK9fQbR2klso+yoThtAWt8Gpp4ibg5Om28uP01rTGOHatHeDvOJH2PSpeMH
IqU80XYCQxNtE4/mVmx+CE1sfMYsywJxUQkj0rMG3AkduWAk0CwmMFPmMjsKX+DV
Rw4I6pG8VnuUAx6DoyGnTLKyFbcskD2nLG6obgigy67hr06XxQ+6lv+dRWgKO58Y
ul93UAdWIPWdrgiXZmP6l6HKlebb8j1pc//nuzKTKEc7G4FICazJo4/StXnt88ph
Yfr9tuLTdIsnYJIdNNzlQKVF88XX3ERpt73046ZytiV8ZDHuDjEpayXLhxlU+dIm
kSPd0TztKmeiR7zpQirs4U1C2q8NKnji8gU/b0kuJUvdowqN+AjKf3TIJebPh3qS
GvBFa+fZ0/0zBQ6Xr2k2q63gK+9ol5+TkbtyUd3iEQeFJaYgLUxZ+SY35ueqlv1z
3/YoKLGkw+Kz2G+ztCGvLkAfZaGwXrcZDIBY+Ss0WIutasZHjaJhLqZThvObtsEe
Ucx/Dv6Y0bXwhuMz+bjGTR76heC9t4Tvg2zXd29OuzoAEhbiTDJzbdXpLimMGf94
9Jf48AzXNwpTi9IotFd65RNoiag3CERqZo+HUq60PswJKa06UkWOjP7nCwdxR0Vf
ajfYhuHsGgcKgKghVUAhViWWYBGbxrs0n5YlRNwZOIdxyODwuslrfJlnFv97J7hK
TDvaAuEmSHcIQoWjGyQot3qhKWnT8WfWaNBYFVM6A/I7JcCHepvGwzF0JMGgh7Hk
0EWBZLtjReDFKmHwhye8AisacLZmyPHieciJCLCauVIBIe4nsr8CKb1V/9p2EQoc
Ytz4qx7mtd3G2wgBr8qmcVTxIO8OAG9Bar4281EF6NVVMNt1yXjUxG/aXssDh9kZ
F9R0kB8sIp7Dwv2yM69+vQNW/Z1NH/06fmaZEHIwPbuhWSU5gO/9/gMAbFz/OjAV
YYKBsAuK7n36VekEnDPkVdARq8NATayYh+1rSqlv+qP3VOkcuYSjF2E1wCFWEPa4
kU1RCL16jS+jmlshi2qwPpfZTrhcifjxEJAys/bzFJmPd5JWuLl/Zh5fknEOkkkq
IG2761hiZjkYqiq1kKjRe8jomsSvgcrixUAi0qDHnLMJZXHoZaWHBLq9MRrI67Po
p7IXmtVnZ6knIigYuN4Wlq5u5whUZSv/oiHdWwBIJiJhy3Z/E9WTTJL1rZAYnlaR
etsiVxtMB87kWdc7BlNMJcs64yuVO9gKJ54K2P4CKu3uYtO5ZyeKdEf+e+xJIenJ
MTmfOUYEZwE0m06Rkgf2lMI+ibCBn/oSF3tQxKJ7c8hA4WCVOCD57BL/Yez2Hwd2
Ycqq+VnIZ+w3VmkZxpzqGl7kVHOMhpgh8o/ZT4sHFrNnppm6xpnFMFwFKVhImPFI
PgONrz018cfJmLoSAbI+o58cfyzXnc8TP/j2ZLQrSm/TRfhX6mXbDJk7XfjzCZPY
DvUAcb4tjGs/yHeobt8s18TfKqYuNARW7bQkIQ/ZPgy4RuQZxvJvTqB3h9mnh282
kVT+g1ALyH/Q+9Nc6hASQn9cmtUwEx5DODtxFd0M8Wi4UBeR3/6dECzJLcUmCYVb
k8/3YPes+SqMmFGAv0KgstxZ7Uh1X89p3t9VZYuhjN/ZG+IeDL9WqrZdmzcu1EJa
V0Be6wWqYHAWpw2T3+9vq9/3ouSFxF3bsuLEWTjidZrqP0NEWpx/y5gS91WgOAH1
3++HCJSFlcPHrc8ndNnWwkDP2LE2mwvPV0zgv7LhvcI+E1QaBi7fPG/VJW/uel9d
30nn+IPX9qgRyQuj4XSCPrWRyqMweRQNagYcYaG0kINAn8P47EV6YdMa/bKuJA4D
kKWHVSxrAPjce8g+Soktbwk9vV9JHpDvDLrvf3axBLOS7qWTgcqSuOJt0iiuvXnO
j3oleRA8tG10vU9KCSsEeKl2Pi+AhI2RX1LCj6tk041USdf+PZgc3nfg/UCc9H1C
bBKyNnJztyZzzXPCiNhs6ZY3wm9QzeikDagbu3vsZgc/9UYUawmIgARcKfXs0HIG
Yq92AxlwRiIALnscuAIXNxZHvb1ENzUvvFojIr68blQP/17KVT9akO7eWY82LYBA
E5LSLO9kx8rK3wW4c3J2CYv4INrRDJF/nrMOcOUYRZiaifthVj2w85KOTeiw9VKZ
4u4IU2GD+i5Miim7tFjVgytaa0DfJ+ReWsJF6Ae9oTBvBZruO7ZoLd3FO++PPJ9C
oYc2ogpscUql0UA2n1RvBpoeefsl3CmrqOhju32POAoSAIm4Kvev1vCw8R1lrjTx
Vd6/0/lqBegTKVnV8BRdoaJ4i2EwYjSaVownZkhhMh7YRnN9q+AMmVAJ7vFa/XpU
2ZI9n+uD/dpyjqf2AfiTYA5OOmyulVgzXAA/KPDuNQEzCCmaAeb7MXXBXAd0qr1l
GjRvtETieoPuqZo+OR6RD35YqYVhXcNde6+H5PA8cXr5xdCclw1U+xDL05m+6Y+U
zhoslo1w2WIwPv2uLw7rg2ogdqobt9XtzVWPE3JVIZBHTAkpPVPrrKaQ5BpE1S9n
PXRoNpdJyfNieqiJ4jMIpfgNVzMqOYedVn5rheMoxoNpRhvPVQpKu9GJkuV/4rZO
W7WYW+rUdYDP3jnpt6sXknpJL6ehXjaRordGT0TciDCSYRVNltZlKvEn124VKTJk
uI1SS9KCqtwFDLidKKqEA1Gq1jffjx3GWq9lsLuRE4wimSAnZT/eTUroqTm1B3RZ
zRjRoc3XDGHSHjHz8hjehNCgyeL2Vg+KI50Vt2wzjApqwcuP4x+gDBN6NIToflkD
YbzUKPZlJAWdtb0O+kI+YgthPJIMzN5Dhf7wrTh9rNRaB45zWbfy3euM1ykinTJ2
lmv2TDCFipyYdRd2YqvunXZKuI3NLkLHHGvlm8g2ikrnBANNwIKHB+KzKH7ox9xw
GAKjCWVjU+juNEVTi3VKBupLmiFr+HiKnVFvovDYUangboIr7eRiLdQeY/+W8Tld
eNL14bfinBhRUzsY7tj1+v+2xwQDIHLoTpFYsoeOe76i8iGRI6EkD/pTonqi2+V8
ICXm+cc/v623gQMSRNldueIKpClfylb01hoVoJYLgGVRQX2TFTY4XjmA1w2e9bTz
QjpGeBlKAsodJqYdu3nequGFCRP+o0gtNfHsvqDBTE7XYg5tpSiaKSGmps/nCouy
F5qUDP9iwl0jddrrUvHZ16tZ3j1lbpzVdmtO8jGXxOikk/e5gRQtGW2krtuLO1gF
4acP5oa1pjEVTNI/l6Y04beGuvaZ41EbvsrQi/9wcF40JcBg8G3LhrEGODixyUs+
pxc84zBYfPVA49rlsBrFZMNeI5hI7wuXnLQHVz4t71ziN9Hq2iz3KBn7BgNrQHL7
pn1ZuNyBT4GN7kgALoyJ3w8KKDQqMiFcPUMzfYmG4C4E4ENp/2s2varTiqsBhJgN
NH3n4DlA04pnRksx8V522cIAaPu+W6feudNi/TlHynbXCf4lrDhEWW/tsyBan02B
IFR9Zxajw82vAVo7ulV6CGJdqspGAtr25Ndr17fq0NBvTFUmNjOeiCrPm1wJ7ZTD
iwg+zUR75afkz2Fp68j4DZoV7NDlXFYIwAgh1xSM1f6+8O7woIvNugCExcnJ0WG2
5VZJvuHUZbQahbEqcAr/ricgQRyFjnQoHZUtK4S2+b1z7aGdK9HhicNMFft34pfv
fFI+e9HqR0AE2A1q0I/0mLMKqQY1fBfX3ac9FxVwDHHCgWlQaxRoFzvYcHA6W4WQ
7FC2HSTap12gsnD7FnTgXH5Xtycu/ZTmWpcsYFsJKtW1Sr26ES3WCVAXYSBZDnUc
A5AHFjnltwwPyrvWkVdRMpv28dXCao3bTU0m+Qr0LL11wt8qkXATUwjhkGtAxImf
dknR1+PfQn2Z4S1LZ8rx0f6SSUqszNRFSentdS+YcT8vqPsQDwe50fO/+APcscDh
P0BlSIpp6SyUnvtS3lT4qG5+3eSW5JXbF0t60E9UawSmMjWl35cO+DdtjpMsNjAo
zw5s8Plxd8vmnNBuFc57qeubkYEygPtJ1bxgraQ/Nz4yzz91clmLNFpOA8EEd2Sv
9R53PeIooeSF+9KRX3ucbbw1TYCrJVlN6+9i7/V+Gfab2PtfwGd5LjODHQnL7+dW
Dfoc1XBGkujI6OrpEwmEr/ick2wfml1NOAr25H4ntjifIO7jnHwoIZW/l+7m8wQc
qCAfHPHSZWthBz80fDmjDXIA4rVAyu3T1n6zNJ4zjY3LsZ4k2ourTy+BdwhiJRbW
hr9CjAP1sxP9n+ruMzNTLTor/UTyT8yFsuiKpuuk9HhX1a1ItejjRtCByYSoBf1F
TBcJa6KTQWAsn/5uaqzIHLDIXM08k02z8DD+vJ+DWOKs3ukfPLL+ykR4WjpuLciw
b3T4g2/miu9jY2S0Ii5F13tuoVW+ZxXRlMv6KiNtQOZRm9GGx52y5cN9FRuTw1wY
Nv7FBdn+3UpQgM/vv+4kaOxNbPLyphTzmAk8DmhfpTGOhoL9WdYQRtR/fe88QHRd
CTP+Qcku4gHfbqiTHB1cYVUc2WxZj48JQvb/AjcSO79BVnfvFW0hefQrkE/o9DhT
rgvWF0DRZSX8yoI7RkapReQFsfAAvhXvMjdjVRrSv4QLIrnYxoazMvSjteBwwDz4
TFUte8mNe0dAg7pV3EeuugIiRs5eC4ihrnxoB1UKyfmgDnXNTgx+K6HAjfixPGZt
Mmojz+S62zpB3FjTTVUUpYr60BmQDQY/ecRluJgdYCNUI5QF2tslq7rfcdzp/Kh8
fv5t5d8pYIKI5CmoNdDvJVVwnsDcdcqp/KO1AToVoJnU7VqL/cU8/Xs8d4RlIfGa
3wKk3Z4YvHP6dCTI06uBmyAc+mb8RCkr5EFE9ZVsxewEIstrFX7OAr1Bfnd6s7vY
7wiLjamuQcWMGgWqB13tmis3mw07LkczOLR8RVT/bO1s2KGFOga3cwrBJCucukBW
N4HTnWRdGjuxIcHjRvNLdmi5EJ4NSxuVNP7x132kcgWEXDP/yqk+dGFC/HmzcDax
sFbLfCchNYRWVgb3icWrcaFjXjm+S3IpDCUQ8OxpHliwFDueOc9htitnaBN+1QTt
Ydh8w+KzROk/ybdA6RVWxg9yg3Uk7xiLJT2qhxYmNs2RghwVQ703gb0V5Wxkae4w
GYhtUGxi5zgN9DkY+K6B+B+TVr41i/q6/pErDtJK0zA4lD5H2mvkQnL/HdxeB3wC
TgBxjtrMipE0SiMnsMVTQ41DpXw2r/cq4yGX9AZ1Uwi1HjXirMmwDN+9dhGUrxuB
vgulS99w+t4Wwv6zbSRTXfLa+w/JKDlvlNNAVFUG8uVbUp07Xlufbm8GnGbo3Iq0
KasnmR4Y8igp5GjMXFyVuhlnMQ0vpEw/yU7UNSkDMVms/seXEuHW7HPbPNGTijZF
O708gGT8a68J+WcVBOMUmEPPZ2XDms/C+5Oud1TFjPgIuKxsWTfHizL8Kpq3E4ee
HJnkX+UJ+wyDpR9z//nu7jhZTC0Mqk2a3osz5TiSXBOw7pxRtj2SAj+n8e6GJx3C
KuXgF/NPTlCbPDwrZ6N985L2nr39FrnyddSFoPKQzzGFGxTIHDbaLB/Sug2WlmN3
aeKAFiL/YznNiOlQMM/vq7mZuu14umq9Iui/W66djBjMdF+it8NqZw0QT/T+EIvE
ei+a1PkedzlcOKC9AMMYFvtjbAIFFLb3+u95Pak6BnFanCqRgH52CZDstWiwOqgZ
73bAC8OysujrG1LEvLqfWNl5W574WF7vqnA26JsqGno5uliwtLkaJPm0/azR2pqr
Q987HqALz7tNwPl/VqMCr9fqTGz9U9ekaRKBGgAI2hm6n5Uh+F6Ox9lhG/wHO/eH
Fvk28xLMLMinjGcB01IJki66E+QHBpMElMTux43nUDLVtWe/GiLsMcTQ5AEmVd7Z
RdcQdi07jYb+9wci0YakLeIvV3fxf58K3HJbCiAtqkmb6aMNhHNkFgHZlYtreH8P
OvtvmwgUgoTL97M1S8DFGGTnMOVRM2sUqS3/EYuAvb00R3sf7dtnRHzkYG54JnCv
oz+eOd7Ta17N5miwlDrIFrfVaquoeUeQzb36mPTZjf9b2+ha7p4+JBkcuGHti1ZI
0IP/qIQsR8PBjdjtMAEMSfZg4SN6ei1Gk9bCQu9HKiEwWkGiIlYFAEEkZmhEZumB
F9vCgZ8Bv791A2fiRLNNQabCXyMRgew9QZGZjpfXuALQ+pDuKwiKBgJfcPiw2bTq
YABvRqZ8b4J+HEu/hlyyDvdOAwlqLGD1kjjxrYrSmPjTRakT9hTrQt9RtfgQYG09
1OLQOTQweXUzt0BhEm890uX8ooUdt3oosWvQ+UiL/xvzWt43OGi75dA1s+PnJQL3
0Fek4BV9svWl30KPQrYpcnZYheaD6zqqNpYfZaghQqm7+Zy3Lq3CqXqpdPHBsPnM
sWx5d7Pvf+Kk1MANXFIJZhfoL2m5/J/Q2WIqZUk3bWemQuH4qXvd0Ov4PMjvJQIq
88F3EX+dp3qRbmHTaGJNobakxj9AowADxg+fsT+8kV68Tyt/77OUlbZzjBEZRVSu
7LQsUbOrPS3QHEhkHFWglk+rF3qEanXdKrVo0+OPVqlOqbiqzJAKhW3MJnoH6XFp
ttTKPkd3h/W18F6pJyW9t+yiwdHQ2If6GsJFQNd+TtwZKDPaREfZUlqIONYySH93
HsVDjIQKXiOLc/PNFXjVp3IRF8j6ARb7/k+k9uX8syqh2+GMaGojhpwJUaxfiyWY
96QgIwg3r7dO0IgYYhO6hqNuxWbZNApHlyekddhddVqZGW46ckQh2AWDEh/tMVHj
Ia5Jo4mnr53hWOw3dD8GOJZbKrIThpYbsH2sJ/v+MK9MmA/SUa4Tt4+6S1KRMBSm
ZT1HNT39EvPsY0zYVlMfmPUqQaGze6M+476hvmel2MFlCPP5oymU7dyIpPleHhU0
uw8+C1b+awefZEmRgw52nlPjT8XCmcQX/OCQGASlOGEEmfYzo9SMfcOWZzRm/rNJ
jvgQo2aZMsCxJUAoF/FrWB1i/6tgyl79R/yrtnm2vW75YYSniS8p6OKG3X+VKi4F
8CTfTqsCL0EaBcmRYKNVJ7NmBYgnLON32mJfnwS8XhMoFR3o8fsUiUNJ6yfhELRY
DAn2Zk0mv1/FbXosJ+FdeSVVSuIPW91jDeN+XDvdFFqtGwK2v5LLq+EJ2wKtnSt5
20JFW/LqnXaJGxDroVhUIx1I4Z54RZd8vNbZZ2kBIARynwz1Qg7gwtcYplKUE3Gc
8MgIWXGpdEqXUjcOp/lgdrUBHgVTL3Io9vE4RyvGmJMD8TApiqaw22betwFCMt1b
i5qIuCQ3eptHL+/1EOzsYpGZXw1eJR1mJ3xqd8+kKn895nr7YVGHfIlkvxzssuFI
zgeaL0g8YGjztCdkD3+Y6clZft2e9UJcSw7LLZ7kljAqC+6brLrWjbzgpUpYMgga
yHWli2WXXDlxu7SqsB9gYb/SSUsHgU6Mxc9NYC3D3VAC976XCuHGga8nckD47Njd
juoBTXrY8cz4n+2um+dUolsyRbX6tMjgHGH69+AyTIe0bGZMJ2lrdnlK8+VHn6sI
EdhLDTga8pvg568RASSYgzgxXgryAwZCcfChcSN7IcARAFG+nqY8KzxJsfl4yurv
bETQvwxfVb53cOQOAVvTu8nqBaRSNyiMhLSwxouGGK3/flGP1fVGX4CNghfdFkx5
mS2UMo1NmlWZcWeWVJsLF5Mn/NzikxCZcX/x4NsZyxDsXvOUrVwtrNEZ9350ZJ+3
s7Ap1wb18DGNqeM5ScycKd6/d/dS0gee3uV3DPRgDhWncHmBVpuluF+r13ZPFhQN
wbigvW/92HZ4KD6SrKZfnqId0LqsRQdWjnOOTUWnYzxsRXL9Uirku55hJi7GVLyb
97QLxMgMXFLzgMQSahcMJ9/umkouJJdLRpKjHpXaYjzIfjexbS9met1kc6iMuCdG
EsBsgGBLxVJ5YTwydSw5EVHFNAYHKqE69ofa/A1U+a3rH4YFYpf8Z8bJw3+fNSi5
i/tYWZvJmmMkpO1MeF2v85/G3BSUgAd0FqQJVHdYyItJsjtQ90ffE5ZCDGfI1wQx
415XhxsliHDKcSPHdKyqK7AFSb66nCIsdh1u4WuQA0Wutlq1tyoMmriuRQTuF8Rk
Uh5EG3HG5EO/zhZJl8HjHELQoqLjSud+bcX2//djA9DvJAiUQY0Zg1sqxa01+sxn
05Be0UlZxwBXXmAI+tERX5u4i6yEm4OnsVzQWYeNDMk4FJ5iHYRG6kXeNSSA1rRu
QZNyrHWCIOlSuqshmHMuVMVKRzA28Mn1dS0X0kq4KAcfJPRIGTSYqv5Fhk2tFlh0
24oo9Me1iY/NZXL/frqmgtmMt2N45FDxGzbBSLbD4bV25yL5I9eVTFwpxOFR4ni7
SvxaloFWLCO42m3B8eyg81gPx5gse9HDhrEDnitPnvjFbOzfmI1x/L7eJlFgvRFv
anCQaYSqjBRw1FQqoAET+HTOX8GadwRs0FtFi/j6SAER1Cvhlw7s4xpCHjurRVxQ
YcwIvXu2BfF5m1dWMyDs1N9UYf9LaICVjZxYsM7NcJOC+2cpMHiNHOWMpT/8AkPS
ypbDtGVnW7sTl6F3z1p3seRzLUHYmYqXr1tx4jMxsKT8363A/8woW49RbNGTDLnn
Sz7AqR6s9cs9FDVczljD9cUYQoyBm4T/wZZ5yhixejAf7xTp5JBsCn0NQ3k57Wes
H+8VZTBMUH/n0pl5qcEeK8/G52f0b37cVkJNiMM/O9gpls2ADt3M+QSyAMwF9hBU
Azo0PCz07bbxQCM5oTK7miu/GxjvEckYM7mG6/n/TNiqg7z97mqFwUr2KDFCfIGm
6dEYFeyQbzNKuQP0PfX38vq6o8k6gW+wB5F8hjlF9Nf28Z0uspB335q+7TjYt0tJ
F2UTQYLEJEiopqVceppHPOKc0Gs7GM4ybuqALevmmt2Pw7Gdj/jMQSWbphEVVd9X
RHPBhZry8mglx0Diky5wRR53LUMaYteCPFokZSwBKQ8659PKezJnz98YyY/BZmXO
ne3mI/ZV+R845U2Q89AkEUFv9KCfQr+jHuOv+45GglsCFWzIcb5TWf1YRDwMtLAn
qlXKFKHzSfZTEzZZqiYGcFyYT/VeheXofgQ9wqAYczLIKStE2M/5t+bVFIX5t65B
UAUk3anVDpWOW/+ab0COdNxcYbNOd6dq+mF1iDRVIowhEAy6WuS3JzgXdVPwgPeD
sYbfV7iM9G1ns3K3EeMOfR89ELZlULVEBvtJ1Cnwj1n86iPer8WvBHw02/cgGfvs
6YiIPS4/cFvGnIyTXIvFA1N7MtCwN1EHq6j48VVziqQ7Gb6a19kNkbAfZYuQ7ewN
4URULfWC63hrbdqrRSJlO6713c/4tYERC+tw+Hzy6pO7wuWjdi5iABghWe6PTMTi
ZwAyMUzDEcsOZSwS2OYbVpqNHHVX92ZAUOB16GXquuejUxqcYPPKtiyK0mQbGGPU
Cvg1WpuFVin7UVuLQSQGaXggXrPUZ1zxo5swd1X8sKRg+YY0W4kTFMKS9uY8Xrv+
X9RGd5Aw1lCO9Y9p81PqJVsxMLvFoE8G48SR6MnPYnhLZVDvyGS3IHODVAK0kIwy
t4FbL3DbgzQFp/Yh9PFMF+LyrLYbIsffF5pFyVYiYfXYMo2IHyMX/onppYgz1utL
qnf4sC72QG9SqVYNfIAG+ezTz56y3KO+B7O1qYT9uPvVXgoQYCZgQH7STOXUAOxG
yuXl+Git/sAzuI7BshQT8tzOSlFa+VcZmY7G41zppwDaEczzgfAuaozm+CofoLWo
0FWmXZv0oLn2UdFslCA0rFiXZSZch768Gj+GarcuZXr35lIiFjrqHgR6St5VlhQV
4yBBPDbXd466chJ6DK6qR0wwCnu2X0OGAaeVvw8peBvph106gCOIGWZ/jqbI0dzY
Hn1TGEigsophirDsSF+bPz+iY8uYCPVEp2o4GLKnkNdfodV8DWAIbl78z3mQz5y+
z3T9JRcFUCXNue+rah20mNCUJ1LNWAU1zb2osPwi7l+EXraCZvl0lLhn+lDUgwhN
CB0kIxkHSCmT+I8czQfrIkJFrneoK68LZ5xI4Zr5+kEFmXrRmMTfLZWXtU5edg/I
TR9i4+V3pGhIXDC9JSMWkxmMzpUrbU7TcRUiCw0tUEv6f2xLlZF+xP20rvS7nDNc
es3g+A8oFCjVDcEYcDCPSBBXmDrls+1rUMdWxwoLXk8nf51Ttl+jMxeTn/7np3X9
reM++92Jxfteqp11KonNKkxKPduyQD7xL+QYhdWBwZujtetmct0gGu8QhM+XhexA
iu9HbZe742iwheFdQEok4iOYLjZhHig/W7XJPn+8rivwP39Zhh304DVutM7p6JaX
SqMVuq9EizggzIh7GQ6Z2JT4z8fVyUElK1Vy6FPToxFFuaBoh7d+6Mo9pG4bq+bn
L2V36BYEY3XFyKhyVmG9UK/zoXEbUVKnur/nYQWyS8/rdXXWZdXG+hhU0PlTUCkW
69eQcRFuTt7cYOLujYk6o067wUludnEbPQYjxpaV5lnwMHSMMlcmbtopUv16msfd
tSVUpAE1Dn2ax1nYkKU3+sy978W1oisC5wbZ0g1XFXIgS4UiFHGcoPsMMRepEWoW
YcTuxIXshz5rspIAG1Ro35iht75JdHMpvn6w1//Q0y7xKA0aL7a9E8fAPYskE/lh
flxRm1eOJmp39INxsMxnJW226SlUJ8hc5bap9LMu0MZS5hokhw1kWF3zM06xOtqT
v72lh4zfsck/Yo+WbNXg987OEge0kIWLuZb8AooPQCg3rzPsBm1DJqXiCr3l5Wvm
vORS9XK+YytEWzNlqTFnEYY05W6CfDco5McDk4PPxnUTY3unHMPq9BEEPjclagLM
cvVc/sneoQ5bDlyFxRaCOrxwcghmyNpFUJE7qrW1nPPN6rMO+BK7YwZxFSPn/qPS
Pxj5/CdRCLv2VxMKEqYKaIJR0NLrCpnZQmXoGxHUYNjpiRhJAE0HfunaFys+dSLL
QHPpNsynJ71dmI+S0+pZcBlKiHT5xw8VINYBDd7IQTU0bksqOWICeO6DEWfpyFa4
kSN/3oqXPrl+oQqFUEVA2YdkbMOPtkejxKWlV4l3LjdhaoIZDluLZYv0Hgr2rAQI
ko0P9tTsELtbxT/BoQ/iYByopuWIMxESV1amYLU+uqGoleUm8NCWeqKQ1Z8G0Aql
sxKM/b8mZd4HbZUgVKOzuavbOrdtrezPmJRsh/KHWl/NBQSATZzu2Lhoy70IH6ba
hrKecdziRONqB/EFcVTpYJwl3SIVZXrPOTequFvJumlJZEZGiId+URqfTyhXFGsR
401uOj7NA9NPqXAe5F8Thx5hjMYhoVNbiE1NirKsr9OwYZpcVwWnNvzwa4oj2lAi
vU3G3L7fd1eDj5Eij1WwJK3y7Ta0uL9NaTmwS4FTqbbxPmM18FjIHPkfGGc8Djlu
23HF4Hu6Rt6d6LiUzBgp94rn1G6wn2Jy2EpU9PGtc+alU3DpD6EwfrsveeMbhrwQ
WJ60mWR2yQHPnxOhY/jEw7cSZD3Bh74Ez779n1akkB261SqMjYPHxY5zxT7zSFrI
t0cWaQt30XMfGqPGPgTYiwuCnsGwuNq+w480KA+QQg1yBW8M1KZwWm9KYBiZJZIo
6kWkdF9wW+3qIQisq6pq26vlwiZAtA38+b5flTMEDBDFkmBblLCtpxhv/2yShNA5
inv55kFEHNuIubG8IfQ9He7CitqCG8il0dfNPJ8Co7mDCWOCbU+1XCAY0ym0q3pA
Yqv18pkdvfRoV6hGI0m3muY5x8cCqgj1zH05sFLPMWM2AM17TNcwlYxxmyPp0n15
wLY7ip2ncdaH5kkvPVkVtrggeQ3CfGRAmOTnYJbWCR+a6NX6jng2vqzwh0GwPPhl
JNNCpoeMF/n142vlyaqKjmP2HhJK77lWfpkzcy/N4us+6zDjF89bPaESRIBTAJtj
f98My+8Rqogx0rHhi7TTpsZbacUXRDceW3kA8097bf9gH/Ddo5oAbyePqwErskp3
7EuiaCW/0QVF+xmBu0j3Z0WuDagqqwwyq+QurzAS44AmkAmfzIFHC5F5aVh+xUpO
/ByKNZ/bv+H5WChqBuAA53eTfKvIpcPpn+DlUq8LxCE9O6Xa9kJyxxLBl2sW9u3q
8mp5CYbYsPkMo735h5zjoE61oT7S3FKjkCc09P7wP/wxG+kLpV+1BqNRmOXw+HBO
JIgnfOAxhD5W9/7rCkwHWxVgtOLxep5pF+z7j2YuHF0mMTYAISjsEv0K07D3GDZQ
AKLSf/gPpZobsVAjcd9QyU2hohqZgaooEw1fiYY8L3VOfdn56C/7Ow1tmZI8tVZL
68Hqm5DU0WMvhRngl/zbTAsutlmPAydnu+MhRNgu9mmKrDfFdE2+4xMdKYi43DiG
rFSPK3z6kuCuhgregvTQLysb5BhJaGsnQSzKtgwL5l36GZ+344U0Q3HaLfvySoaH
TOSnKRfoES2aUKN9GDWWYUctXVaLcCTGgeRIrvhaDyN36zet8Y5wqxSPDM/nuBBp
eYg2+5sgver7WVSm/kgGnC2OjGJJbp2AeGE/7Zwz6m/0DZB9EJ7uK3VAKM89bC0u
RL1q7Ty7c4qPZONJIieUsXX5MnKpihrW2tcAi/UWgqi40TDYVLYAYRANBXdXq5sm
jH3wkDkkZQJ7kwgfq0DZzjtHgkclmiiSLfbNQCttidun3wDesavmDBD/XfTeiRDk
ulRMFRfFUB4In0BSJO6Ty6Kx4LEMGaG1A9shwjKTbDcCO6bhK4R2ywGGiDpPumff
c1w4YV0spA6fIH8wBErmKouyKg97d5OR0k00T9fsd7MPxoNb/GnR6VJY0cE7GzjD
v4XP79YZ9aaNKw6A9To0wgVL2E2XBg1Oe652jspKW5LUTbdJNfWQkp2ZVMmbYw2J
weRaUqzSHAs+3smEmVLSYBBJpVOhh7qjSaQbJ92ddCqH4XPUvgjEIx05XFennuGa
rEVqLfTwlhqQc/oXRhLbOu5tpPxVrrsKOU55UGZEKMnP1P79HeCk2BwrrR/cIjsk
rwEVZ6z0xsBiof26yt4A+GkhFd2rXfQRhmKF25Gb0owZM/4lpMuybHirVKHbtx83
4NTIJ0u6Z8LPat78z1BEVDY1rIYZ+JacKbVRjTyfjRcpMWQXVCB6tyvMk00KMtHh
xK6QoRzZoQWhpD4MkhEEFtVh6Z4fyqYkd+KTbpAzyFlD+/UVzbZo9WzOiduk3KSw
tXFGqzpggkowZJkhWG7jZC5NTkrmWphkhFlExqFoQQvFf+kD6Se5TTSuHAoen3K8
IgDYuLn0w3Ja94LILZgwEeewNF1j61Asfy7PyEOyYb4t1OtOGSfDawqUCnqzv+Ae
sOfZ006CrBbLTCg3NrAKNKG9qegp0lfmlveCP5vM6ZW5i/0yLFvkSM8j8Q/zHL2C
OljROMjT7uYMyySIDFC3Cf/XuSqS8x+EWJT9LbiRsy8TP9zHCkk/pr50YpO6iykJ
CP+QYIcaLKZAW+kOTK/Xij6Da1CTJnZGYOaoblKPy+hhec1mvH2Jwn6RL9Lxq76k
of0mQ8OKGManKZUBcZndjV9tHMjllpbzZqvGMcawhD+kwI8D/q0eWu4S08Y24yTv
+2cguB+oW6ce7t09Zfy27SB8jF1LLS+fv+z33okblmAwkBt3GPdufu7pNMFpI5Fy
gwk9l3Sla72qOzWHDnhwqnik35YZR8fdmHo50/ACDIMQNCuD82SvOvUGI4SvNTIj
H7iV80s1jMgH2p3IMy9xFLXCMWcL8ECnturWVb2qo3Ga7bqc1lOK3g1ijvg4U5Oc
cTDkYrwuuej9nUTg/c6b4d/UL3aJY+js2+qVi2nhtqX4TSIj0tdgqUgMaH9ZWROZ
m0wjzKf0nHnhm9+mSxRGRjJOpqlbhDBHsA5JEH5Oh6kBBkArLlP76HWd98IiaKpt
2DfDt0QdK+eQVUzQJx4TyZlnZWPULjzghQlmiMrJLalGJ0Yma54Pp8x0/E2Z5VlX
9uEDD62FuNNmsfQl59ejemaXhUs9Z9P4+DvDSeLnVf6G/8h8sPrqgXA4N1r7Mnfr
Fel+2kIopjXZSBJcW0zOV2O9GMuxe28UfBYpqns+/PiIoOuU6MPPBcyxzQqQlC+n
eHJbkk+k+Dt0X5TjpemBFGoBRqkFJacftcMyJp43T9FVn8zqygcBi8HJsPHG/JDd
NZCLpNj3sBI89vSUGcqQYcaVEmFnbEu1WV02CVqUQaKsNjzY1jHfQoO4pa7vcLuW
UoO6HoUC1xpAsNS0djCY61mPR5Yww2H7Iowg1/jKeyMdxa9GR1x8iGYlmeXtKA1B
Bh2ey6Fnpe+FUriqU5lqGYFhUze9BVyizpblUStAOCobqJ6NckhyGtXUqhFA8Gax
Qo3PCQBH6vkzwkBoCUucyy+rYGPcZMlizNyf2+dAuoXwmism/sJGBGSLXwHAlVxt
gnPDmFah1P6dsXQPiq51vqqHR9fPRNuTrP5pmPOVDIeV4iKLzPZf+pie4g8H07DV
lWbiYhDOY05NHhpkx7H1QsRaqSd2+mMjsJ1LYOzYAGSBfXjMbDOcKC2g7thCL+PB
odibX5ryEUEcfqBU+IZ2TNwIhiRx+kqcPJ37QQeXNvlpIyj2HWiW0k3K/8Oe6rKK
AKqnBow8eagePuOlg+O/LWycQhUnwUdn99Pe/CvBIeX64tiC+wI6docec0dJxbmM
FcvsxSGLxEulUmsvyjPBAok5brmX48Ix6R9gog0jaMusapggl/+x9GG3owDii68Y
fx+r1PbFGxAhJwrrTLCfWjOSNFFnXkjCTC7oWtwX0fMxfi6UANkj5ZWhoZZL2Ikl
kOJywzNA/91bDFKdIh4ENBlGqfcq/Igk82Tlz8X/UcdksqilBSHIoqmXQV+juJA1
fmAKflZ60cJy8QtGXpighCc/3STa19k+xwMmmZLjcmAXey+DtqbdOxpclu4Oh/A1
0+WY71l+hKJ2Psk8vman6fP9dTjzhE2fS5D/C8+jBLo5JxdygdeOoW98dphRN/Hx
BAUgc86j4X/Vll+wivk6iqIo58tJ1FQFNlNkOcwkRZZl4jddc89uSg0seyZY6+rS
sCWK8yKCB7i93f/EhXtrUK/Qr51ofkQZqdO+7WyiVCfWy/7cCrvPntTGpZ49k8tE
Gn/N5OzwvmPqXbnS32M9+asLnsi2Q2umLGgdLa1vDHYOt+srnTCfjBRvNU27cLfr
/EcCHiZmTdf6WuK3cHLlR1wtMYb5CSt0irE4QPA364gXUrkFD/9E19Hz9Std7YoI
khH6bzVUyrVJjG3Sn3n2qB0lvgEgTGqMxyyC82oNyPa+msABW/FTi/nV1W3mxTyR
16AeKSBl5E8R9O6jegnwXj8xCRfF48AphMVsuPsu/j8glX7kuAUP4gS+DOYd0VdX
5XwYdYBae4XatA976k2V70XJeBWe2rt+TjnNbeb+LYIYTuPv97VIQyAQ8YQDAGpe
5P18iGO6i03B43UNdxg3kVFrjP2W/iOlXw2mSCEnC8EfXizVh8MXQkY5FWSMap8P
6tvIQH7rXnmKfdMlgdNS0Y8DAepWP7YvJNIkbIawJfxT3hcXx5bkOOFMNWzD0xPp
NqLwGxIvYCln/OO9QfXM5q2tSUGAVDdoVGegDzaMnr8H53s53THl3NNhVFaWKrsz
mjDikpEJtPgMRMtcdcA1ndp4wF38idkP09velvnAwfxZq6Ydw3sbiqrV07RPLrEe
M356Pv8X2TXY9oH1DqW4wIYQAxpK2j/I+DzwHSwsWZpoEwm4DD1qYxa5/+OfXKLZ
qNFhWKtjMTNKzK2UOCH18S4zO0dWBv62s5f5WC6Ac5BHo0IdqVQI0RxJ76HlOR0R
xw4xEzD79BNOLbtki3kdIAv1Z5EWGeHjsEyDJAqlHwHeNDVTY8lWTjoTAtVGXEMn
tloByq4MaalczE6Mk2BhyNpqw7F91VY1AWjlTQWKvyjtqVXAVRVUPLHqYNhnBpUI
gY4N92YSlPYWZ5zPks9ckJpRJzbxjFMv3pecdtpgN6s9lfhINVLPc4vEIr1tPEP1
/mJkXIdmc6RciQa61ftDtvyuqOecixcZS9S9CPLtEGomlTaIW5r84y+3Hyv5rYL5
kHGjcQ7pWjhg5kAxj+4NSUsfad0tK30yGFir+6zG5CZ+VAe2bTKptCRVaFXGmyhI
K70c+E13x8DCaJS9Uvo/4J3rChYcbHypqgCbUwwjB4VkGSseeJy0mgdP/jSIH8sY
6p41H79rA9Bszy1whcxMXPCymuPN/CEEqgtA5byKKkp0WA2OwhbuRpX1lyeUjTH4
V4gKTglYc6lba2GYkVhRvhPQIT9uUM7Er8yM9ICogMl0y1/C3PN1x/LMti/PxVJN
opJ5jOW38kWj7vwBOA1DtC25X50GgbljAAHaFxKne6/HyC9g9ZvE5jZdp8/oVquk
7mvE5AZoKwbemPSUDvbKic4KpCf5Jo6yQn1lLhshtQMx6fWMT8S+tFF+8uokg5gh
SJD+dAfU1c1tQ8j/bHbRcNW34LMJHAN93TUDsaRlfc46zco8DTdzYOSuDQ2EcfgY
8giIW7Yt15RksP6+YakfzX1cpdo+qmsSFKt7Z+5BBNB5ya/j/QxhGk5yP8QZWIj1
2Lgpcf6/nTPj1caFYPEU9biG6pRad/PWu48okstiiNTcXTYpN7VHh5Ts+ZVY3kKD
JO4lEyAZcHiYQR3Nu0WKBYvoqyJVMQzwrVqJO7UEnbAjALqQE2y1nBsymkXSL8bd
vIpg9VPHEpq8rdmg6FVhF69BUZW3TcW5EWlEIwqYBRxuPSe5oEYdNbk5mOvumhXP
nZyjHFMp91Yyzi3jUmZLN7BUpDvBWU010TR8Ngye8balrPF202NzbN4wkA6SViWC
8Iu1/0G5I5vVuk8ByIC/y7YVgKSPIjIIwikY/0gRyaX7cXe/RJBa8fiESSXhjJr0
KgRs23/U6Xq+E3Y1rAguO7mnUltE8qeZzsn75MeuQKwvMCwsWkqXRVFgT/pkubgg
qj+NEZ+h/uuhvKuLuMWkINtNRHA9Y1UH/w9Mld7VPpcqciKhGasRVlmPTwr5uw8c
XRsDnAcoVOzVrUZ/A+XDcItCQjvUsSHyXqTlE1qTXiPJnbck7taUyP+7DSEUWmRT
4DP7HkRAgAe3DrryCba7tE5nm1fN7zBe4D+LS3S2rAlVbJB/WTdVe4xFEIrgoX6i
K8o/n8rClz5lwVlCvILdlZthfYAK6p86EoVfB52saMmqR2eln7/Wp+upWuEPtsb0
6ZV/ISPRF0VsEEoqc1mAUJ8M8fp8Sg1S+mMDSZCoLbK9GdqinDGVRu88EScvCCvE
zQM2+599f/gP8rDdLsuVde1GKUwX3NiKujjSGp6BJCcqICQg9PsqezzLh5HPOpxT
YkkhmgHQ3spgtMoSuPZc2mOdVw+bod6mVdIannTbYnErapBedXIXU25r7Sdw7CKm
TibdPM7eUfHVAg04us7z/KCOtF1KktOMFwc6wwI/OvxDiolBYSoe/vq16DEKLh9e
ZJ7/Mx2yTQ9rlYPcN8p44hjWpntnkE+cAtrbSuw1Lxc1mqEAatldG2XXS5lFrPlF
7BfXEiYBTffx6StkaPdr4m2Cb9rZYMT3weInDWykn5sI4R91voEap7sdoSy8+/rO
4cd2/CivCmlKW2sLUBNEsaRQy2ASQRp3FBUmn4R9cWXlvX+aLaq7ez8iaHN9QUk1
9n4ZIqqZmj47zZ9CAbeKij7uSMnWUP2e+oi5YtmN7hpOJiinEht3BLPYpU1aOuuD
paDh7eOlLVCunrniZ71Qoo1hhqTIp1RTRGnWnezh5HL2KIWxqOblYOoCUyRQmk2X
dVHLf07gcd/X21QmunDAO7106q5cyJJCU/l5FVR+Bfi+dGneI2kBykBGwcVgr3Rw
QpUzoGPI07a5bVo7pSEyRmrT4I382MawpXwmJxBQcJspeUnTuxcarOvWDSJ7ruz5
7EOMNIM9DPUoykoKRGyhz7ubVFO7qBkQu59/KjR1pG05zM5BveFZv2zfwVYv1WLl
t/61PA6wT3b3gsbpo3hmBFpf6gfW/+dSHYcYU3CH4SfNcnuU1xqNEt/7dwE3m87I
xs3X6XkbHedvxcSWCSOCLPyrvNhuPGOI+C1Z5r6yhBwsLxOyCcecXQqVitlIZclt
E+xR9W9oYLx3ZFBMjWP1eSBFDQLcAkSMJDSVvNtOjRVCOWAnV+FAt+ed2xibnPq9
N9efHJC0fxCd1haLGrGoHTKiMt4pSxPg/sSQJKA9t52ljPuNMICLLohoLaEZ6SP+
dYcjcUSkoVePHDJ+OipX39tCFbSxQ9T1F8WK3F3gyDwvU5qojgL4jrLRp4fZRvO6
pTe7FafzYUl5pnCpp1rEKNq4hv8Osvpi9Q79jqVL/h5mKjB1z7DtZY/IJdnOiAvo
jorGZqJR5hodUEc1qt/fBQoNfu2fGzvtif6+Fl2ZR7wlZcZnD1uqEJNfJq0tpAbn
20YVfEngRQxqG7y8R/vsTo9FlAek55NAHIEtlBL4MrJSTP8i7SaM074oPggl2+H2
/+xbE4OtRaSyCH1dFUgi9SVPdenOwYAVuRYVFRU9EXOwtGau+ipdAXyX/qO/rFRv
WFMqfy7KZed/JURYjI7ahfXWZpAKbB6eoaYR68QHBrrQfWH8uMX+XYGAnFQUaLHA
8Xv+FnDeDXQTWR7Jm59w2M/kF6MQrug84Q3JN4mpai4OnysA+s7nsiYLavXxfBHn
BaPRrUgDU6awgD1MAPjw1Ze2K3CN916gKtoIaHeNK9v+/1T1DQmBrI4hrGtUlsZ2
nvDlrqjVoOAk3bhlautWczBM8hb6bJYqVvOnerCTgz0WdL2qTuauKoxAZBF2iGIB
QCAGfqykqhgOeU0x3xPIrqS5MPwrRAjGqe98R6T1W3F+q8kOUXwXQlFWoGMJh1Mj
R9rojSGlpS1m7Ke7UoU/tZ3xJGIA8zXzSrsvvBIXiRrRqtoFOrE5eQDX5GFE3CvK
nRX8FLP8V8GDKiYUzotcaSNUYxPPgo4TKi2LyaIvvBVICm7vXk9V556a1KRkja9D
5LJ7lREhGLx+7odFFoKJLROzJMAh2BxlTi0916APDJifbcLWJRS66apQzSx4V85E
mOwVkn6mzsPcV47sIgjeGh7Gv879BPP8YHwylnXV/xLdlTPZ5OSZznI5W0qH8hLm
hq4gn2JKlJWOkmC1G+FPvCEiO8hysTtJ17uQhSYc62yFvW1lIPb2MX204EEchSQW
2pYuMZOaq3lHxKFyBsFBKtPVGcpNKWJTVy5RvIxClNzwc1PsAMpHBotOooFvONN/
Zh3eh+G07eW5POAepEOuQsHGG/eAJ9HwcUcSXmvnbZnrQFfb0TiFZ7k72MD951PY
v3mBtZyfHWznerTus8n/GyP7qh56QkWfEHBPIv3feVaoivfBPinQN2jgI44pPfPE
9m5gOYIKhuUp42qnwMYbB+Haj3ihN+J7/l+a5U/mF3taWkFISADUVrWqVKHmqqqM
uUec84SP4BdEBdKyAmsFcMaguH/Qgfubt9Pn5fHwBq4+JsETsxi6QdN4+wtUp9al
7BB1k3c6tUFTElPeSK6b6z3trPOTGlhVXEYmsqIR5BRgn1H1SQzp8BJf8dj/SKFm
rry5Cmi7A3PENEfmgRcdnsgoeiwNg6fNt+PGr17YS0zSYRPpRbn4Z2lxaVjPwdtk
5+fYiW3g1Rs+PNmO0g+FC45ThpXyi0dHmRmHJZk4Y3TmrxYOa78qtb+HXXW82il3
7nwAM0DCHpqP6FyYDGLgsMZyQ+ez8M7S3iwbjLQunnjn6FJx3pjZwPPLEr4GTQ6j
UwKNMXH9ltBQy5bSL5C4RKZSGGPd0fy71QSnnKDbo+A0rLdaLJITz/PIQGAnaVWx
E2PID6kIf6lzXpsc53hf36CM8jHCq2QkvTzWWqE8oBnWC5FxI1e5ZWrWy/vbn/B8
YvywXACTuoQJrnma2JEknvzr+JPkLNaQRiPmfLK5mED3CK/+dw4ed3jo2lIPTh3b
jdjzAWtR8jxekfTyXGahdY3/yQJ2q9kwPKwHqzQHDK+g8iFWmL30iT1kPlpeeLc7
IulirCthB6bFH4Ri9M/MuFgEQJkh5+OnlFDxK7DQAkC10jsLpXBSDD//WykFJFRj
xwXpIrF23/JDfB/KFxAHPzXWF6bUV/04Hmr4Kt/oHN5lQADOAtoX9TXywAW36bzR
ukjDr9G2XtnMlI8x6c9wv+evqeBRiILYJmuXwOxZ/chS7x8ApVO3rV06ZCYNfawU
BmSRiHJf5jGOmoe4ZZDg2nsgFMqJovHAJkhLumJL+PXQcTloXZ0tMMhFiS4alZRl
i2s4HhUnDs9CSVxZLtauyawqgSNr6yORVmQcZ6giBPAQGPZGuoPY4eUna+CUzxV/
iz5OBw2gHd8s8sg/ngC9lGzZOcStIXKSrgT8RKDeuSpciLmd1rnb26kHzWg7roie
TebgOA1gh32CQW6PDmzm/JVSqk9GpCxXoxEmXKlGJp2KI3rHBb9s4OFKe2Cui3K8
vbC4IQf5vfNfWzcaX6QHDTfUy6t6JyBEuku6LuzsCroxXotOcuHz+GhuRRxe36C2
7uGhWl2qivK/A/EfPe7UhNOIkzjeH7et8tZxhKL7hJfeNxZit4yo9SkwkoHY5iNa
QqZT/lDaiWioayr6Rp8f1PuqTaT8b/NqHs4vEnbjB+0zGxuAHq9nQIlSni0Hi2wi
qsuzNrR3I3Y7TSuC0utRKFnKiAyWD4RBEmZSAW7Np65rScLUSOgR9XmcrmiKibXq
NBuOLjFNq33BscI/P0tvdP0+lUFI9xizXf6xaqgsjvgXmFxc+OlRsgb0YRiqr9ka
gpmX+K6LUUJyFJYW0fRB8p+eUDOGPuU/Si8OlzhozGFYvNS1SJvVVq6TYd16LfNn
FYJ0AjIoOhvDGVZEusk3GmNUIqyO6apTLTlcEy6iHaRJMWvhQrHkpHXOMB0VdkIr
OrY599r/fm2Zn9ixvz72LgwTzyUaD0OOCgocxnTJY7v4POJ5gbcOnos//mkF7e4b
1If3bUKJca8MQ62SGzYyCk8+WyPSrW2EX9KEFcI3GPN0kphDYqr7rVc/NGMwAhek
hKgBGjx5JWEALpdD8mqqatkMj7ay8jk2kMn1Wb5emjYCi4Q0sJLvdbSyCoUYALjz
9FCM8FYCijtp7Hodb7UjsEc6ruhDOZu/QTg8sHpi5QkMAkqVmT+ozF8hOSprjEOu
5db3nQsgDYOAIoyyUqSCGaUMxwqj2Yzoa5P6l/6+sLH1/mj+t69vSsiP845RWmrE
zOjbq9Dca53aSqkkyETiFkSxXT+PcxCWFG0LmnKy32upgwmAnkEjNuUcshqa8ItZ
WsVgr7IBkz47PpVcbH6LW1RYrH5HK/Zu82FlWCH1EgqC8oQldoGJq5HeCai3hSb6
EyMnbJmCMEIZ6fDt2M2aM8KGKR5jVnLyCA6L9sayR9JNwPGyKcIw+Lj59Tu5K2NA
/rQNCtNW8/Fy1XgKYP9FKsxf+iU3kjLJ7dYvd3uJvPSPNl95q+r5Ut8tEnz3Xjvm
nCUDef9kWHsGGHwYUlW/ru85s8VDBdOcMeM3Mp/yXdr6Tp3uvNVTesYCw0iaoaNx
g2qnXHJoXozg6OHs2qx0IjwBi6HOwKFE1Wo2dT4VXzPEwTJH3aqgfSzoL2JEPBSO
AZm/w+T+Xxgk0Gj/bCbkwvYr1XCJ32AjXWxZh+2PCzCTzO82zg8BpF2uIYq95YKG
mZpi4Rh6r1BL60CxzmP5wIwNikh3Wy03FsRgaW3M1C+F4nqVsQKbQwlAP0vm5n3G
avwRl8zpJuSp630Xqh8wSBLe4ywfx7Ne0Xm/9nwNyKrpTQ7bv/loSKZvCY8D0L5U
7bgoPbhJto+JS5FyaP5WGUG0sFNWLN2RwGi71uKv57qAd02Kxo73wrmixTBaWwqO
ntzMsb63kaJupGxA7okOSTM/Hmu+NVLl4Ba8vM7mX17ZZmR1/0e7w3sIbENEH1GC
ZdJW7jRXEYfWP9Shhx+V/ncydljbl+GWDhiWGbhshvf52m50mWwYmOhyqEPu3Ebr
VD2UMX3ljMhERUyI6q0nIpM69Dk3r/zVmUkrLCt95+mS5JjtAAXDusH+b4o0Zcu5
X78BUI1XLIOaRChLoPclZX64UJRKqr2oIYWUpdDZTpMzwUskyGr6+DSx8lvCnY1b
DFsXaiLaN4RQ5oDXNnA3QtWaXz827XNfrWqn2MIuwTlUW5kpi8z8GSsV7ODbT9qM
hwANwFFZ/Bwi2IO4IJNlxJIoBGs/ZNbXZWcIFPLEoOfEwQMvoLJN9LR315BXpPY4
4qz6Jenun+nAeiH83dIbd//XN3fYDCwiR+1U950SVd7x/dYSr6hAecohKA+qPDBz
In9G0iZvU4Kh3sLaPfGPMwM1n2f8dp46PnpmErgV1yYjd+FnX6j9JNP96D/5S8nR
LyCfagb16A0G0Vg13BmEkDNfht8gIs9oZYUYNAmMVOG21XwX3wjvQs8R8Q1QOiMn
RpPZqL0uqw3uFg1ZP58wXgR/Vg+Yo85wNlUTRAHY1fE7bJrmm0TQnHApk9547lH+
ZOxHQq3CZfbD7WAi6lSOJ1RVgPfTfDo+69ZygSEb0IWN6XC5DwBD3UuBGtFuDro3
s0RzqeWdg7JZ+qm/Rvksf1n0k8bn7X92mF0humaVKsIbTmQAjOO8oZkc8vhdcZnS
7bz/swa6/nFg3fJGjgJtbogQOcVCgIX5J+p4u3EDNGlMJsFf5uM22UBOVwN7kfqL
gVyw0wF7IIXoc9Fgbg/kG8WTntJ/ZM0V6SI3doa8I01asIKPP2xiVF3aSMTruiky
a8SojoOTKty3rNQWpC88qUUF7Um2uBgo/fqRA2NTJz4q0KSgqoqdD7INBRai7HJE
16F1h/UnqJ0/mcisOCfov9XdyjQy8MA9Nn5HYIUL7m3Hin80XUqFQ/R389Z64qtZ
iIIm0+XaDLbagq7jkihDViX4V80xLIlt5O8Ij8nB9gpKRw5QIKdACOhUSaRiEIHK
XYbbn6adLb5OFLopVax0HGST+r4oTLDYY0q7o0JimDAIZD11VbHnKg6os6N/24sH
NO7iUk7Q/7Gs/ly7M4KWD1GF8jH79RHi4KLi6beMK9oaSx5zxF0W3lTvcTuK47lI
iNllKjTvb0TIubVKoD1RD/IATD0TNZNLaD8RBwVJ9O3TLF8oUEUeNbOqLd3rE1YZ
0+vUFXWNvOnOmTh0F2kQPfc9dqsCe4hrwus5Y7VwSykWi4Z5VP/o/waxFJdxOAry
y3um8Hp2CokvPMqtYZ8jLTufKEup/bRLFyok/nAMq48LPyGRQpIJxoogXXC7oAy5
80b1nh4z9QQ+2nRLh87dMr3AF3hxYWqSs/Wh+NhvKyvJwPeYzT+l/YCgTCLq/Fjk
YHiNyRRLkNPknyk2gigh6aaZrT4IT7FvhLssMeNHo9LZc0fEzTAPxWP2kceuGOIQ
SAIBVLxjsk9Upto8WKxVaYyq1mCAWltNRmMTwmQMhGRbsw5y5opNdFLmZf/Djxhq
KbxcIVpQ/j8/kqbmqXyW1TmJocN7QjYbNWfVySgMhTlZxLZlpY4Iigrmh960GwTX
SEd3CrhXTIdE3LRtsnLtWEJeUT4dIy2tRS9eZcMpTa9VNV1GSeBZpKm0xy0yTHq2
upM07MO32QrjSQSMBiBA0VuYOj9MPjZyt7ax3yjvAkofzaRWhro6eaz1oY0ncjRJ
Pk8TIMGOZaLR0xLo/EhmsCJen3rFv5ilKQu0gqu7S9xTs0ZLoNd09ZT2Wt08IiqL
9rpCQr++9aaq/bIXC3LwsdFch9oo+j0FO6sxWhpd4dw6z2qpUuLY2tiqzWAXfFog
VKbWiME9VCnHzDD//feeyC4vzz6ysXFt18vX2EUBLemnqwi5GqbBvrqX00FxTCK5
mj5PljPOBXi1TtWCUEML3LsryBnPXBzgKsiA1M8gNR7ryalDJ+c/PRiXJYCnHOMK
C5EayY/8wymibBRrA+Ww5tGd1ESgIxNm55tXS5WpunjCJvlt0eMrsSN4W0i0hZ2J
82WgsAgmUJWc5qIip7UR/JmVLRsSksY8JHrnX9izgdLIXGgWANFyHBE8zijkiLW0
k5V1AdJcmmFVL9K7O/aUAJQjWif1u6ubLtIV9RqsEsukme4wCUvxhOXv+UL/or8O
LSxMLCqs090sz1/kXKhOUCh5/t1wmxozY84MFDEuHI5sDwlwRWpubc0CL+YOIh+q
saIrY2Y3E/PWuwBVXe1AaWLGwn+Lo+yV2wX5VaphjDbmBU1joqe6tc7GeSZUwYBp
N763Qn6AawwsU4zYwILKhHTOTmSuWmkxxFRD7+nUmHsro1ArOLxdoEDGHEJxOiFz
x4VFxFtjR3Qpih0D2RvisBXGlT0wZpbe13J9IPvjue7rYqbSl/caEosI6C3fovHb
XyMqpnPoRBcrGGXooTTyte23OO2eHMv53Wu8XxDLFj4Q3Brmv3dNtZJvSZLNV6KM
KB0zJ3fbqVJRRibwsJ2x1qGLTlVNivSEQQa2lIkPw3jh3oPMF+6bS7e2N2P2Dq8X
rgizFvMAT1FNAJL+ir/u8aaMn8qA4CeFw1IQEeUToOMe37RZFNOSTYdApPXWLREl
ooTwF67V+6z7p1o/5hQ81LlF5q/wgtRQusjiIqQvK0mM+ySYh4SAOtWehfInP3Bj
1yjr1mpUSuIK6RfiBPjE4+SdDD5omVm63cWDJHBcjI95hl+fSeAJiiVidDYLsv7H
JGkYBCGxS14V4FeWwOC3Ue5ihbZa7D9RksUJJhD2FCDd6dzHeMUj6POu+P8EyOxl
ApgHCn8tTdurkU9THFHQf03+txrFy8RoOKwWpGvHvElptSTcmbeOv82BBv/dJHQV
Z1svDxXsRfJyDuZn4hOvinovcYns5LoKVK6/W4IvPgIJmTzgZNU/Epml3y7FiSAl
P3iT4P4knGX1FAuMM7yKKAcMjhQPHZvhAh2Z+LkFrr/eMesp7P6kheYLYGqPRukx
Jbx6sbTq40dj/b4MSeJi4bfQGYVQrVy/MrNfWWih9VvJSstaGMFZmwaAD+l4j1G8
eqgfQPbWHLPq2knJa0QZWw9u9o29vAOwl0EQmSMnaUBf+HcxKA3PsFJVbmAt+H/K
FMX6FEs9GBFiNMDpdYgt3GPpG6KMfcFXPALfFRkJKMVcntv08Qg2LtJvJYj3ssxu
HzBT63U2yj8W0mHiL7pGgBH1eb5OrTzwyEfnStPEMx4si1g1NMRoNFwwfx4hFDD7
kvFXZXE+oS1Y4LKb3IypLGtArwfgK1I3uIuBg+SrDyn+rzl+VgieE5t6dUvzAKw+
DDYPn28Tx6HNz4DpsCEsT+LsbNYFatk8o7Xzvm1FegvNHANrN8KlWXAhZhDc/+k0
ofsBxAaasrLAqJ/48Pe/FxPFuc/Wg1hkhnAcFKURacKgf5BVudRh8Cmjb3g98Xsk
jscRM1t6M9USMrLAOuJyMFodUb4K9QV+C/2IBL+a3J+5GR49s0yMwcYcbFnbjCyC
hSNP8f0fTeTn+p9wJ1QS6MNt19Xi5XIr1ndZLFebl8MXCO8V5ljkKqcOE5g7HFvA
UxAFtd3YeVKLV8+/rAsADP2NOHJcMftbA1L9Di11v2fHHJDIIzRaBOrHYAOAO3Ys
KU08v/qy+iWRS7hc7XiKT1+ZfCRkTHDWwb0ahqgwjQGa0t2umrxMX5CzDzm+wegD
JmwbxwgtAqJXSwQl+jUrAel7gjlRX7OxSaP5GGmSamLrkZQfoGja8qdaT1MWyuKh
I845jdkN1918xb689nzftSSYnolsksZ/g2hvpc5wZcMWnQ0KSWY4nfqcIkwqKv6O
M68N9ETxFuEkHzG/YzPuJOB1tzF8NDa/KumH1lbBAjaN9RpgIk3lsFcv2gemR+kS
2XpRle9MblUqx8o5X2UihdQfDk6EQt68Y8sxLYYOwj0dju7HDLKysk75Ed7w3kX1
Nz6VNxQndmMdTskpDm8bBpMyW+bxCqBPgCmNJ2vH06d+Vdw85tJgEkuNJ7H/7TW8
UFOrV06lTMUyXaGoOgag4Dp3RAzSyILKNubUETmduS7BL7H5axx4I/W9EK1CNw2E
67ODpe4Ce2w5r7fxoXrO78m7V1ymAhU4ND0IeBlZnkmvfLntOe1kvj97Z79Lj23+
ulXtIlXwXTyFHqRw9C6KydtZPLqOBHnz1BNWK9n3VC3lGAwUM/+qSf7GP3gnPBrC
3Jgg1gBUcnj/ER0MXx/i3Sd95nJvvEpGbR27SSlufn9Cjr3CFKoMLw+yF4tjNxF6
U5hrF49kXdSuMjYste+AbnVbFbIt2sPxWtStCJsbZB7r8bzjMgOIdxTnysCVYmwG
eJrGUiguO9ie0ICkjo40wLGQ82msBNit2pZAwkgKaMH5146CMBd8EiKd4sngewW5
iCG4Jy3kHRSqm7UyQv5pyZn+1O3aF9AAzkAe6ZYPsxncbBsNUPtj3sP+aPFjhJGN
HVzGjcLnaG0Em/zcg+4n15clKOBPY9OAjgC0ETtWrq6yqG/N/RDqErluSCVFY1C3
H7ZMF/bk2b352oedTDE6WplbNdCZyghz1WNVxhKL9K1WO1isIejy4s60NSJmkc+L
ymw0QpwbfjTfvBWP4nDdcharYNxid1TV4cacFgNKr9oE5rQurHx9NJak9vpjXZ2Z
vlNUxxQUm3eeo0pP+ljWBoSWyv7M5D7KjmiigcYWb7iRzkIRM5qY+suCjFCU5jQb
Ipz4dceExCt3K7YVxV4L5731DoTViUMy5gOEMTZHj3sr9yoBcsbqvC3L0XDyN3rQ
48ZW0K12yZb0J27ASPSAdXG0QeEsDOXU6XFLRm+3JSBeZeuewNRrDm58scx5TelE
mW0Lvjb0t8ktC7nksdxOmBco4o4WcDpWsevY2AkYHV19MhPhFKlGQ/rRGnTXeqkc
y7pwocephiB7/k5jIgm9R+Yl6+lK/Ndk/DJyI/32np3fBXhJtIY3F0ZoaGCK8jYJ
mclNV5dmxKusruNz4Bo26TqMzDYPtDLHJQ5qwt/+Q4Z1ydFWeBEOjIkM7e1vGb/r
HHSF4cl8oAyM14f0dXTZTHNB8YXJAnL/+fv5ew194U5QznEMaJcDSun+HC3BDzDB
xTPv8K/aa0JqK1LR3M3fcrZxuuBjWwwBj4ZMAbO0pCh6rt88senqppimv44pXp2v
x3aL0xZVfHiX641FrKRMFwhUgaFhM9cYyIDytnf6AUfVxjIOCfBvodxHrVcCBdDW
45E3PDjAMhFq1XxYvJGJMt7Rb2rlqlwor7Nm9VhES9OpKYkzMQMWzm8BQXpvur6U
NkuihoKaskU8thHUTZw0zoInCHDz7apJ06vwmlSahZyT52sv/uGoNq4/sOhrjeJU
7PMd4L0EtxoGuqptNTynM27SZ0SrzNEm/OoIrv2yc1ITHxTaEwQ9dE3pX5rVMatS
DbeqIROkHqCJfyhQ5hTKXpCaJtJchn1psiRsBJ2rSw1LSQLBljdCPy6UlESRmrq6
cz2ZIctYhU35AaS7hXObNvOjbkMSdpu6+UlR5K43Zv76L95BAQgisoF2cAQ5nnwt
DHEHyCGT6Wm/vA6LsYZxE5g8Q7ZvfhTSM77G2FxoNJyR0xJ+gSPSRXOAR2yJS+H/
6n6aGjYhuuH6d1ppaEht6cXke4YDayvvEzKvr5rTlZfQcxfqxIDFfSrVlCuc02fZ
X8FQP/QXwGZLmZeQG+B6oXerM4CC9bKXBYl4PGq6bggptV9z0df4a/2yoo6Q1Lqu
cEVrWMU3dzWKZUzTwsoGwgVDfR78FnXWJPqnIffLqjoH7zWHf8LRk0gZpZC1CJJ9
aUszYCHI3REdXdM89V3PZj+1q30d9ijk84IwhP05EAzctV8+xqX93+c5+yC3MQb0
5gru+cg/1V4mu3xFE+H+QeamRqs0/dZjcd/AQFVePxkuMrqpcWCTyZQy+PwRtjJk
TXjIfiQwQZpE6/tsTxRGmR1ajXIpkCvOfAM7MkGAuMCRAc6LWyv7gBSw+AYF59KJ
8yiO601So9z1RRqFayHgN3fzucgqz55qMBFBzKgUmZ9FaRIuF9nyVs/rZch/dTaR
JRU/zKuTYseww2EP5PeromnO5qwleJBXYiYv5hrkY3+fKNeTvPMis7UpGOu9kOwt
XCImXZm4fcch1tjmSNj1ZZkm5ufMibTnOPQcvlY+EQmhPeHdyfOANvxlwecnMo7L
cr79euotPvv36btaCIL9g5WgGLFzByEwOAqxn4LgYj7FzVTVybguiN1HZtRXaXYd
NSV2fU+HQfQlYnQUcJl+KvaRhv3LtfrkWiaFdfdq8KBpWxexexf486HodPRMvXTA
syPhlVTv3aAtmIeGabGJvH+WDDP9x2+/MoZMrseJ02v2zaGYkloJqPyfX2mvFVOS
VTRoQhtufm/lWwQ9c+SrCBjvkkbm9hWyupVl2FiuArUeY3fy6wr60XNnkf4YFP+u
2kAkpHX9+RaRoVRzwZk1QgeIt8Vl4bWcQa7SFm/l/TrRcAIvDMRNbaCDiJJOQvuu
LzsK+95PI0JqlaSaNB8vhU9YpNCPIwxBwmhqpVhJKUQ//Bb5pqbVKg1l2GhycWug
K0Kg/PZXjGkNiXU76W8i7ZqEpQGe1a6+gwQxc6uUHY+uv9CoYCY5c9hLNqPurE5N
znkLNh8OBEafHRwW3ZzH8UuDOSUJpEwVU7rJjzbeFYebXEd5mp6LrOpn6S+9/v2b
oCzU82bg8v0VmtvKuqt9stjchBdNkZFxtVCXEO3OIkQ7k/DFRgs4SERt+ehC6bsA
iTu1zomuf7z2IO3qGesgBPfB1yuMGWho7ZeUCaGqKxMyvwbaNzqL6G8rTvDNt6fs
PbGjL/hXDO2qKpu7HTEaJ+IAeacDyFwBUcFtXLT8XIOeJ3HItNkjXUI2WWj5UUw9
q0Vmnk5DAyMxwum5AFRdtJX4ZorpP3HXoPJxHVoYsP4b988+mR4xQuCK0l1hRIJX
2cSTag2/Jx1+Ni2yozanAb3Ozw8IbTtgxKaTKVOL5MVXJ9eM5LBRalxM0HLejrba
vYj63HqL9f4m+p/fxMpilp7ogasOZq9/yFi4ZvUdGcZyz9M696i6FHM5tY+O8oZA
tDaBU5ukScuRaR2IZY4eWdTCcHrMBJ5XrAtvbaYtk3TVvrcqkh102P/DtYFgoVSz
bASWE+tnaHzQIJCdJEfM+Ovm8aggQmCkkO7ognd7HX/YWlaW2RJLa3Kuct6Ssg9e
w0s8i653eAOvS7ZqmjaRaYZhsp9t7NfQKuYqIcgg/qolInPC1pANfrYE824QLkCf
XV6e2tjse+8D07Yn2mBxReNS2IgXbeo+OKMDF+8+kN9D6wiActcWxy1OU69llu+n
qk2xj59CK7zqNCydLACvL32F3YFDoT5W8FEotsaPl94bAg+Ju8lTsS3slTyMXCfY
CrnlzjgODA4ZmpstuTKAmXAFPgP9fCvBjiUWYhDrSH/d31es4JXKHvdJXvZWuL6C
CPyRQJFATlJ/DvF6AOSj6do3yFFcGPVu9edmdvMFo+ugCAsBpcGUIzGU0aBZFgi4
3pDInedyUNHrmI3oxA8Kq0m71Eo5op4Xq8GcCtqC0mV0JGAyCQrnTXTIeJe5n2Wp
23OSQUYxVTK/LHLrZqGbcIh1E2deopv/f29k6CjgaPDBqa39dv9rSMFCOSnLYFa0
PpL7J0NNl2lK5O7Pv8t9Ow+p4BeiYgpimJ+NC6P96jDditOn+DWUKypIV7Jpq9sB
SEr2d0tox3cRTjWMCfEcxMkdwTEDfwHgIUjWAQ2kwS4H6yGNDQTdnJKWHCLzL9WN
iLbQ3P/poJCedf97M5zfy643QvZAyn9Q0XmnMJ+M0B04hZHM1q/ieG0ev9vzjCkK
0EilAR2bfLWa3Q+6hobBY20ySI5iax21cG9ppQQF4xwvsjyjbKgr5dN3uwCF0JXw
NPj/kW3cQY3WSzgZmuMOqfYIwxdkvwBqgnrAxZacEEay2Ta1LzuHCEt/Osmi00vs
20zbCYj9F+1Q3maKZ9JIVfnCZOE7FbvH1AEH9XUIbcheI5l8TanRE0C03QS0KDXS
a41fUw+zIiB+9kcBBSKcB1mK/Pdxb/nSQdv9PVvgLsjYGos5G3hXQZy01nN3d+ld
oUnwBq+JLhrX962ntZAmjzueHXaqomUKRegNZmbamcuMmyRJZ5ZLnzzMa7qdO/Pq
oNa6NAGBSFz6xlmooGCfUsqDMQqSYYTXwBVP6bwt0sqrgBMXp0ZJD2+xJx8FKXb5
LKH1I+UMAuvCR3DZeYVnXl6GSB6NHyEyotEgA4E+y8ksg4ngz4mI/398FGR30oHn
YL+LwxiepHw8pbny69gX/c9lGWIneAF3AtDLQZS007mdnw399sKS+cFob/ZSurMQ
Znfg2SQeFfmI8E5XnC6OmMCO6ye275RZFamxxWuQ5O6IxwbD41cD5YMn6ZXjtOMj
VL5OGJoKo2bzBLtrRYxBrPvHITvuEdQG+cJkmm8c14f/s0vUcdhpCC0uQ9EtoRrX
cYd5j8cifp7ZlFYsHvzaZd94pMWC4WjMC6TtBgBGxnyyl53a+xcjAVSNCjhWuJ42
USaHQpR9esjArZJTUGE3m3JGExXrrnmejsjeHwaduZzFLljrsl6Ip5za0w1glRfK
LMvgz1r4a9ir8kseNc/PR740bjnygdJ8EUt4Od24jHGHDeWJ9UH5ylLZEU3e7qGW
X5WXiVFPeSRZ7Mjq9Zd8k/uQdVj/XLp4ytMBqQQu9r/qrZz7zCllrZ07ZHV33iOi
Z4fj32aoLPgV2tE9SiBDXYDQzd46wMjxXwju+xy0QyQ6iWlNf9YFULkrVipNZaI5
6hBuIlp4qw2bcZeUzD82jD7LGQ1qC2BuqS/i2B5qwnGZ/XNC8kBZe0av6qe/maAB
lnFj/ThDS9Cl9QKCsRIpvtsBaoDw88YkdKAWra+E4Yz/KjHSoFvVRxeHnEsljlY/
izeAclo5hJfAQ6hGVO9CamcZHZixiFTT+gGHexS6cVc10FlkucsBLqoX6nVNCERJ
AXPry5Lwj0l3+GQfoafEpnpoAATlInqN3B+gKoj4qtnWqes6T+er0fvo3KA2yXtn
cvDn8t4w35psxN32HYaSIb+veXKFt/sfNZTPLhaq3bTWG5+SyTzlx7SQXEO2/PqC
Pff+wkqSvt7JdhajEBrl2M6xoi7u4F7YVkJaaGgpO6oSzKJSj3h7kUhZe7MlJFOo
7qzJXhSwr5Y1EdylqkcQsSv+FiMghowbbqzMPKwa/ZqCqS3KJ7ENmQFRrKBNcr7P
2Q2x6ciQae6ue+fha6J1sZ9Tpi+5XM+y5oy52qkraKe8qCP13LdB24+HxivnG9pQ
HAF/KZHl7nXhavO7gL2gmE79QhoYdlrY4mD0ScSnbRTa82xBWld+W7DahCF1gp1e
2ZuisQj0+0KHVNRbYsEr7sIT+2nVrNOTZg5h1o2JidAImnOzKbFKE35UIqbXqDiZ
A0+HxFDmAgMxpVZcbUJW3tzbvzl17NTqZfKSNJKGuTqCVimyygyBUwdlEfZyM21z
Ck9rXSSB9WJXkd+0DdBlIomhb6bCBt+aShI+f1bq3Q17fM6dtmYspP5dFWBOAJ1M
7Mg9IoujBJjTBF+cHwFsngOX9OcgEJmF9H73p62h4oK0Vq8mCqKbE7nrCbNgXskp
NgOPZQlLQcHK1cU5g/GkOiO2/P1OiP/lIxNNdP6BoPFxPJt1zy5nUF6DfOXgjlEg
+QIRVhmmxLyrJS9u2In66EK3Zt2f8z0Kp4XNSf0l5OjYUA8LAUkJ/8E6xC7qj8VK
7VpROQqD814GhboXGNAqOxVO122vis8Th/idzYc9HG4tnZWHxfSRST2ZQxKZjGkk
CXJUoLojhoXbItBq3+KW/MA/CtueQ3heMtWe7sDy7XYAU0OUnBJ5041wi+oWUQ46
IkWM8igm4UnaEdgRdU5trKLyGSk+4h1f2MPqIkrqexZhYkbu+wOCYlnhGd81tAnX
hFjpvltTXAaweN6gCu/pvLvZduNm5FmSEbuVu/V+3f6ls91Sfw9tfiPJDZ57ubNG
+HdKaVnprgqjTBt7nDpcjeZqgCZmPqtf3LgAs0v8hx2z6sWRZ8FFcYlZe4G2zxVP
g3H9x5lnLcnE6DwqNk2pRMiC0W3nSXE9NUC+zYm7OGx+0Q8cqFbsKhOGEgxdS7Oo
3Iu3BFaRUKEhWgZs5M0bFa9MYxsQ0nvUdX/RRReXp/MhcqY/5OhaGakJ2C6F7XiH
xx9DAxlsQtNYZq9EKWdBGZIHYBgrNSUZrc4XnXG2bROUW28hQYkDsLGVYIGFA4bD
j6/J98U4VnpxwiOAwrMN9dB1pjjUsK9+cM3rMX5GzDL7XnHtNWBzi3qpyi+HEZkL
dppU8yehaAbWTkgfo0Hv1yjFikd4wThimb2ZU1a4+PdUW5r+MQSI0N0cxSopv8uO
l5pfo/3sBziwMUGq9Uf6UnEX/h5o0vPkWwS+ulDzAStCK7d4r1FcPlPwO6eWQ+Hv
ev9FYD30U6rFN/cmbQt5uKdvkfDGDL178EBfNFOXXG4lJ3DXjMrb7YwQzv44K5OC
4T19EK6SBrSka3cdfglPHp1/Bowi19UVf9NVuQzcNgFDDgla5UahoCIXTpExkXje
JCw0s8KG2VDge6LoGh5ZqZrMiadonJdep5pN82COeBbJNNxBV5hheegQ+PRcb9J0
3FH/1k1FKQ9W+L0pTzeGRZmkEVbf2v8VOast+3QC6g/sZlktH2b5bUbfwBHz6rwa
Ghsky9GEygmBJ5j0BZXglOSOZaykxAxLsqDWEVxYHtglPgKec9EkeEhZJtAhU6S/
5yekPnb5yYoDbmgd44EMShzW4h2zMrLGX9lgThBqMiH1rXk3LfuUDvXVOFODusbo
ZeMfOBOrfUGRqSG43tgrVdPr4zDLhPaQraOaG70qwAt2+o3puubz7eZHNL2v9VpK
FddlZWH+EAwKequng24FMeeZ7GG4UFo6K9RHHBhcUndaw1aUA7dUPQDU2/wealSt
eWVSd37GHEjSy1Mjj++PR9YUpT6xNTrWHebHCkvbS55L64ZbXoAXoFzyWXix84fT
wFoFBQkDaONfnygrZRVcCCkxCvrEMuIkHf6cn1DGlEcyViHrn2yjKIdzt6SO9LY8
TWF/jKS2HdO5GfAQFNEsju+4oTzapGKuShLm0CBdtDWY7dHFEGxLikbaU668EwtF
ldVxpm2obdjGo0/nueXXbZv5SjGJbWRnZYGfVqILsBBNNEPlS5s0qsEYQKzWDhIG
bW1A5t/pDid7RqDqw/ibwr2jpdMpCk8dQ/iM6c+yMWFHLncFdd8uC+5pmVVrhh8w
1hQ7PtAJKihQYq9JlOY9b5fdm3dEeFG3j9y3KFG6+2EoOC1mmMq5A+niz6XOPa5L
/gVnAR6VmL/fNVe5CzM50iJNe9BJiSmFLrnjZCZlpOJCdrwLDCBWeaOQXjmqvF0t
Ow6cfEQCJC+KgDOTZVfrORx13RGxrUjUV0Sp/bPiR3mKuNqu7A0KH8+1n07kbhI8
G76qB1Q6tmAKgks6jC3K+JitbBuKOWz0cSvzwGqs6AJ+JRaUxJM2L5THhqc1QU2F
G0SZeePZ2ckBMKAEXebo2UcNZhXBSbJ1MfTrZziOS8Nd2JQpxlsmSv3pTDPSgW4L
XuCOqQbs+AiHLS97lfr5WUUBzsz/xbcuyvX5oDNE+0Hiv8sWWTV+pou4IT7muHJc
H77ZeHlLdD76L4X5fx0bIdNCfOxCjqS6L2NGnoGktZqW3LzvGvdQ8rkf1ZmV3AZ4
7JmxmkQ80JORVAopW5qo4jNJllMyf8xJJe5S7VCW4Hpk58Fftl+Y444epIYsFJ/X
+BjpzdgHbaVrmWNTXuDNN/zhCqLZiWoh9cLQDF4AnAgwN4d5ngZSpyszEHT6NuTQ
1XJq1EcDFKVQMdxiObz1XK8aUSIhIAs++2x6hdAsZ60g9rycelAiWY83foYv9ODk
A8vHfAU3TCeVYk4F+g7NqMgJ8k1YcttZDVU9sl16oMyGjzeszA6GlIdiAjn4kRgY
KTN2XlNhJzkgUcpokiw/H6NjHyycoS/iu4chENsOn7IoEKBLv8KdH3NsdTKHdh4+
v0BBzjh1VWrzAB12TXs4wFm8okzNoFAqYXbnC5YQMuOAe9V1zmkgPMYr/UC98cze
ef7uCM5DUen1Z3O1OlfvTgoTmm1ERZpMfDR3D8YeZc3L9tn0Gpc2Q29VWvih9WOF
FvnT+dJrVrXYFV/zCv1Knhu3rtYh4VTBIghC0gkbDsjCXA+64MnvG1xkdHn3mEOL
qHWRJxIJdiHd9oJOH2n73YYeNkxTb1yXdzrW4VbQNvhiRmZzuDxs484Sp8eg/jd0
S7b4tL+YDb48L18dtPjsDKWbyXQCb2ocWV2kr+XeuPj/b3LQ0/egz7F8CGyfYMEg
EIwxPJkCO553pnSTcyxseFjioUnlX6KOxsifqzRj2mat5bvewQkhCsVW9BFASQ3M
VvC37jzAkH8SNUrXOUfWw9xRVNQY74Zlf7StWQsUjjio168ehMzKij7tnxNCwYKy
XAR/UHxMqf5rXKxAKvHDIzYjXyxx3iGrJrGYijNuhA1TPkqy24G8yHvMP6LPnoZN
FpLo76BVIPDm4t3RBx1s1y+Df/HAhYT9a1LkVT/StwfMJUoKo2d3VAd+S8AaGejn
ilmLQ+P6+z1cLPLDnr0jRNRESGAJ9rUvQlYhRmTN6KBihuxDiGu6ScKRET5DssGy
vxIENnf9FYniGcMWNht3eJ5hL4cBbP82r+Ouyk/QFrZkgr/s/ngAbIidmddndzZE
I/QcLqBB8sFCFSefng0ZSlgA66ozKQZTsyLYQcf/ljvriVnrEiBgNbAL5iJ5h5w4
Xz4we6lOTO0cFFK8DViyz6TS/In+rT7RGZDf1Jifh8WtIMd+04RbQY5KRNqroYLw
Z+5jgoOAYYGHitn4PNtx6Z2/pC26vb6Y8a6pNaLvVSqjhlDpEuD18YdHqQ10RJaG
DWG6PagRZhwzgkvn1lFQRmCZWiX3ltseWRS5cBwPuW6k88jsQqd01QMghgqmkOZm
qsr5fiuIRq9aKEoMbBgWfATp/Lf3sLTPfRkKqWvQcIU+FT7T54tzehSaUYfK40gy
ayHsMkUgIz3McSGthLce86bcInys1kFfSKCWZJxDCvD+ckV75k0vGL2FIci/aAzc
8IKTQNnfMLtPpPkvSKm5aryFUUZxDZFout2+A+TWM5IbBPcn21jh6Vo3c/kH7WSp
IYvPYZCW20BFrfNdTbRBqx6OglMfeHxAgOfwKmaHs/CjU2MIjsrZyUW0CLi2zW5c
lDJcV70XJQiMQbVCP24SL6VtcocBDF+zgn6a/A52alZAYoGZK+C9KPDYwHzzq74+
d5v9DadmGXueTizf9LjPKKA0awndhGRG2auzMsDw9cROXsyKof6a9drwZeT8LYPu
Zo/oX0EuJHntCfgkfSusqihLJpEz1qrxRY706vmO7VjefnkVACvGcheOM8EHMFNA
lVNxltZBagrIOTQU/Mziv5/Vnk0TSCJ2e7tPooMcQZZuCcB8G502ANbkCZGKwIn5
dNxYQx9Lz6SX73gX94rZ4fDk0Cbr4oMCAOLTQHYFYB40kOFMrMjBTOcv+e856DI/
HzygAgVnWzMQ/UqInTwbawuqilLqkAEMi/mRBEr3B6Ju4prOL1q8SQ+rNEz+xY3U
X9j7XDtocpswlMJV8GjrRGxt59JFsh9M5eD0SUJaBPaVziIVZgkdDVmMp1bOOTeY
B6DK4U/5j6EE1urpGQGhBmmkkcZ8rxH7dng87gVv2jKvVY9DxDZ18g0yDi+a9+nB
RZWt9rVoiz8ENiyG5DpODoIS3BaMqdao7LauQvWYSCd6dMN6/GtESBSpvVF6L4Oh
2DY2/eZtfBh9XStCpTSUvI9sZ/smr9c4EZgMWx/seaCfiPvjFB7wGP62HXg1AaL4
CQdAcU9Jy+2d4SAqZ/cPvPeOfYc3w5UKqJZrrbxMEls/qUXUvJZJco4kpBnZaj6w
eezpeiBMQe+rwEjLdNRIwBSQmcQid6O8B6MBO3USdcfXlvgfGTDo6rQzzbqSH5Jo
KYY3ovdU+A9Y3ldy2eU4J9V+LdrJfM0VkMYw9AiO2u1mtd7SgMGmd4BA2rzxzgxK
9yY3XyUyFgKHw4+j9HWFEemkhX6Titw4l/q37TnzZTgBJE6NnURxEYImH1qygkdU
WpDn+xiyQc+PbpjGlWGXf539pmC6g5GLqvQn4n5UnEUv7mnEr0XCmHyM0vVLfptI
ShclVnmAp0unzeFVA1tk2p8a9SM+aDGuW7oAA99Yc5GmKIA4ptx31CwF3OFrud8L
HqRygyPP0MrUOofw0XiGZERFxHyHJREXBXMtIGrlzH/e4Lr/z8PX8oB6Mh0JFFnC
pvgTUt0OY5xnv9f26+AOf5hRSgVCa57cCQNgalzFIrebxPYefn3LGlIuyI/rTKVl
R+6d3BP6Tdzb9JLcgGwxeSsEhNnsuNdWSRzGqBA+vZDxi9m82np0+216CbhUSuf/
4mUgaV0DwdS1IWeoYFKqmbxCwWj2tLw4m3ejEGNT7KVI7t7o6C7KTDVUYZdP49HE
MZCCadmwWm8smW0SkH9znplpGOhe24cD4vKRilc7ECNmYs6wZlUgdJOaIlJ1idPB
l+PJFHTYlpzK6k+pJh1A5i0eHzf5qhK8EtVwxLaCh7zijeSZDjdz1zlAioJrda+/
7cSVIvk8JYuADobovh4+Dvd00ZDEl+3slSq4ln6MDwZKriDAie1sWYLl/21JpJDk
5FF9TrsbDFThRbw1xpOOqHBAx7v9pgAYj5dpBf8IrPpkUoE7K+yG6LmNK42TWVX5
O3HQGgr51RuOiXc00XwM1PLhNd3XmsfEdbWHkb5usk3u2gHydAlk9XJTmT1m2vht
a44tvxiuPiuMMFGW5aioGU6nUYxTKUwRjSs56EDHk2pOUNySYaU//cS8U6xOePTg
p50bkfeV8Nnz5YnFiTI3n2znqDtsoD3enZgId0NFdCgvQ2Ho+Fg94DsezsVCWA+H
z8jxS34gwc6cdNSzthcUglsZXi29FqwPXTm+0JGbGzWKUfviGumdqxfFErh1c8iK
vRljgB6GPv017OtZp+NdFD8LjbVd0fuWdPSPh1yFdxKs7vqr3DJpwHE6HmN1vcq8
s9W643DxJ5lzYrjHrsjqonKhvaJjwWVVhh2vb3lYJSuAzcjxliYhPt/x6LN6hSM4
iXimuR9ocvZLIS4HUAsd8QxM+ud8LH8AUyfMIH0XJEUQ7sv+sUncasXYNp89gspj
Uj26yS2c65ZAieZMpGrAZVLk7ccggMxrboBtu3A65uBN0yfegzUpXKhe9xYeTplt
Kx0y12Q7zC0kvQ9re9GQpmE7aj/LfTl6HEkwl+U9hVxfpDzuNnUJWkD45Z7Tuv8o
NnUYHbbRtpeOt/HBagU7Uvl8g0IwsUiFxNzfaowLvse8tlSGa39Yv11tXQa6V+l5
fVtH8/m8hfAo+s8ZBXdGCA1nJvBKpadqqx8bdFv7Fq8fOWgQJpLCekUlBybbJoQP
gfODFbJa8SMvEVudsfH9eX1jwtJKT1JL5qsN80kfcy60y1xFJg83feM+zOL8k+zp
+MmRm2NcI0Xi+ZqnBKcA7VL6/MXxciLcOonhqJItJtx87R9S6eGgnfvyEnmE1Z/s
HFZSRZcFULks83wrSqyhKz+RBhvSGGx3WEaURLp2gdVsbrFLb+2AQDdw6mUNa5fX
W/XSWKoIui3SwNp4ipdfdKF+I+cQJeZVj79t4cUntIQlcQ/MjXKX/OWyIU+p6Qvi
iesHKxblCjeQyemzxPsySmTLwQ1SLMajaGXFHOf3ms/1POoFRkX3OE8FBqZDopK8
wAmCxyXRCiPJKyooZFpVdOV7H0lU32QF85x9XBM16EF8ABKfWBQuLkF+MI6Qj3nY
h0I1czMpI0sqtJnPtytUIh4egv2GbzH9Iq7RUNypwxyPbqnsxGGnqJZiAuJ/q8MY
vurhH18dTHY8Oc+7XAOOpFT/bQ1C5ASUudTXWgHTzqPrDRNrSK+8UF/aMhowccbs
bFkZZ0Jh+T2Sjc/++wG8ZjG0fIN88qjBRhbZGp6sSt3tN2VDFvx5Is/hkEoo/SrC
CLrwtJITRMvTSvx994J/yFmjbGWok96aG4n9uUwiIRY0zG1WEok/wPKx+7YA+3OR
iw+BpveYp6mFR3ZpxZk+bblAQnqeCrvxRNAZ5ZZfP+ArQrf8DuDGOj23w8b79fwV
HBPuQIehPIuhBM/tfvZXAu+QaB0mVT7yJzMkv/4RcfvtDC7eVF76CDV8cdBSCbkq
deOf95eaOW4vIuxECLXLNedDZ36CnbbH9qii3A22HPbylMP25DliKIZbh+pqFb8S
EivlL+/f61oKOQAYl+V1AnrCRJSHoYZY0hK2wyfU/u6FuEdZwc+TPENkzc0PQ2gT
JqwYiDyINmmvNCJVh7rKJmI1mrKwyUgu5ex141yP0V9rnUtOVvr34firapaR4NqY
JYidIdkFARoAq4nltt9qGrAlRMRS25KqTXflKZ2XRISTgouZH6A/7OhvqgGm3EO1
4vXxqQV7JONzamVAjWDH40s+Nmj28XebaufiPbat6P7Pgsj/PJxw7i/EgTBZ2+B8
ADA4plwEDbVnELO3KYgKI3ZFaJwsC17A7vMOGKMRQc77IFTpvSpQuAzxMl7i1PBO
Xykj4nnIjv1yP69wO9zJvJwusTsIdUJXI1fn8IN8JmV9/Q3yp2ySLfRMZJxStsz2
5sLfA+8hpCO/Vvp/yNmhxdRDuqp7P8JO21R1GggE/fL9Tck3UUP7LvggeAs1bcX4
wYRxMOE362VQeIMQrHnyDKI4rdaJlY+M+KgkHIsq752lKDx8a6vFuhfppGvDU4cP
l6UCN9BJvJicC1sH6JM7TM0265W8uvfjvCTcGyGrc/ePzzPy+fyeJHcABh9Kfkgf
NDR/jx0Nl3REC2Cr2BW3QEs/8jbxUSbkBFYy83gP9YaRS0Si7jwxTGm6T4M/TnYQ
20jJhtBTD7Ytc5bnpI2H6+qxyb8WfLXjVPvlFER1AgO9qZNO4HXVctGdQ+bz/yXP
iD9YJKdbPaQVoD9FF8PEB9TpvkUZn+avChFxnORb8DA40PM8ittcQY3sATTi7rNy
AjHjE/eUTv+X27IhKZgXg8hBtrDgSUziv/65DtOYaF39AlmgR473GB7Y17KO9BCx
HfBnelYUofuYau0evPyuopLZXNVdnQ/S3repM4WmZcDjc0f9qw0HDh3m8Hj+24A/
MJUuk9L6l27SWkP4P5NHPHCGNpUh0paE6RW4Hc8oyPh6wXLfvogekzyeos5CRkh/
1DVpjldWccnffcG4i/0v4uPRjOdoF57RAiz1YrgSswrXltbreBPIsVo56kgF5kQW
x675pZAowJTRJpSJr0frJfxc8foqIHikOAQETR1WIRDwEYvHgbQ+Rl4o3PR+rM3S
jvf6T4KwPeNpyjP9k8dD1+4GLEMZUGbGSNsf15rnlk3hFlYO5oi34FtqxYt2Tf7I
zy9TkRQxtVp0JzAjanjsDtDZ7p0peVuJyccJTS9WedtYB6JcKIx8Ewl1e4BHkRpF
kXD5bpUXcMMpe52gSdCKSk3rT4kgN2atqebhwD3cJUuO9TzxW5Fyl8md+x6hD7Pd
N69Gy81c+74k/7Uf/fjEoZ1MwbkWRS3UNWaws7y+Wk4CyZO3Ngm5KJppQsc0yCcG
Gn3ZJXRJ/lXAysI3UGe4iZPjjCApKvhb5FYE4FpEPm+yeDqIKAdGFgtkf3NldPT+
q2Or5MW53uidVGUNfcwaXSar6QFIQgHdEhdp9SedKUqg85vZDc2bB5BUOQ4p59A4
e1hx5OYBsISwG0W5CZrn6mzoRMGKHjUcpbjdn8VcUOHF6i1N4Q5nsx/2U0Dxv3B1
dVPUPvKzzC7v49f15C9JEw1NRTvTfq35cnr0gKEo+l7IbkhQkbna/gjBPdJ6i5Gg
mAvb6m7jW6q+PkPmMbYavBQHHHlInsMgdjfIEF62ERIkPB3VlN+roLmnzgFZRM8V
pj2vOLYJUaJJPUvDcv4rp1RVThzKlsYfs/jKc7TduA+sg6/GULZwGutkJzrex9rA
TI9JljRWoOdcjahbOfNbtZfXDkQtzvSZ58BL2iwcIY7mxNr/3t+fwxYlLbNEnJI6
4Ez7vvmbBkbe5s7Q1Z8VEcipOuCkj3XcoCysqCW/EqYbGT9bH/4Tm2DxobS3bBHl
C6NrFSzHTedYN4noVj4bNhOGFLhMfgp2Di7sCV9iDhfWH2Es4ZVPL/frMITH+Fsj
VhTjEr/hV68XwbR5xHmT5rUbrvWYglJjDsGzTzwNtkfq/7iLt1s/jt1F0IHYv6C9
M5R6WZQnkrkbEm1HEJusbV2SpCcBCtJUG/rX0a1hnXGtu8tch7x5cezcFvCRf0xP
D6FgA9CGrnw+6GGLylWQdTMDDcmVHlKXAOJxlps/3CswjIoadMKYWDQKxLdH/T34
TOmOJti7GCq7WWdfLLM9BD86Ko/Zm26TzpbVVlO10Bl78HD0TouxR4H6h/X29ImI
ezwM4GHQDoEkDMUkZZl0yBSNbKDuMR6LfhvoBG/YKzrDO5UxBh/SrcB6qJBZL2FQ
jxq3Q470bgVzyRnS4aI6JAzgHrhh+fjqjJJ8S3RoU4UUzHHLGixT6xwiWFyvQDLZ
77cBHaMJm2TOh/9THenSgFsP4NtXL+93OaS4cXry2l6C5HbwKqoSv8l1kNazq0TC
doLTo+TUw64apxhRgHEOFZT6wJwSZ2neovfr/owlm/kbl9bivA5QDlgpD9advEQ1
mJ54xZVGgrIcUH+g/oDyaIDpgPbNiy18iBN5x0IN48z3iJQbEkzRYxwGk9QRzOqp
YpjG/T/v0vn4vumpVa8wU416ivMDhEu4new6i3nCove698FuJ0+6hJAmDZU3nf0C
2gpZwBUoouRWbBoOLqRbqKfztljh2pHNOZmW8tzccdSiznilAM/Gq3PGC/38Nw96
FZPsCziXD0JB/A0AbSBLFbL9k4XTAUJuPj25Lqcl8k2B34AQyucoqcNp8RHLqcjy
c0n+UO4J66rl2RTgXttPI/5hnv2QwcbEfWtvjXdgZeCtD3IT30Z12O6jKkhsoXvs
ZBxNUgscXp6Tdq7uxM4BxQDbEq43bVQRidtUk7dDygImrPUaG/qTL6qXfou0sHDr
yH9JU8nqFUOe9AVbHtW8yu5z4bgKymtSdPPyntalaqDdBhf3sZttgaOUtDAWJVKg
8kCqWaMDOK7UFC+CzPXqd4sJxh8aLTDEsIIo6LSBbxGPr18UbGlMziRcdv6DaRjW
Y7XeC7hAT2CyBPaF8lLASUDbbX+y+19tnLEZ7y3K49qDURjhEQalpGMNKSwwTXlB
cY1OaN/ewjfPfpPSw1r8117FiUXyW9b7WjQchZcEVYRJiFvZhxNxhX4/JCc/8t9a
yNxhMYEd1qWNLmnM8P1FqwiQS3YaCHzcXfbD71WcjRDG3Ii5RxwYsHCAGX0VR/MM
sqiSP4OLT0y9S7s2dssBeGzVC0ZVnMx7zkzU/nml8jXO0Tx3J9KCUIiK2ddb3/+W
d8PlqjCV9hBednupZLcDYx1JG9y1vCkouEtjJ2OiC6iQFxOaLTm+djf6Egl9G8Qc
pHTZgWlF1/XQHl8PXl/rFm+0sf7M3PRdnU84Ny71I3fjGb+CP9i+xmWxG0qttYn4
C1FX4Ggx50iegh1isOLEROoYr3Up41UkPZAR4JJLgjx89g+wJtwG9Ypq7DJ4t6WC
8K+FASB/No1bz6zcdndbGcwU9C0yyUSQh0nrLhV7OSrhg9irpAWp3zXXi5CxMsmF
nL10GhNBp1AJ/FZhJDM3gGbVro4kPm7VW9U1cB1A2pdMxDLfco8gEa3Q2OAMzGEK
bJZQ+9end562TfbOvZQLd0CVOfo6wts58Kc00rfxpq4Ht4uMuft0/PtV24RKd2lZ
E5MSBlG9GKnAIQE8Xf/7Efq+wDhIomWZDf1LGQQ4alraCJxSRKJ0ZHqGt1yNKiRy
evFiaezkTrqPy7vjF/jmS73i5YumOMqtVwcnWsvhKrld21xvhl356UBRDbi9HKH1
H7aeWZPA2ah2Yh/rROEZ+PBD6aT5BywivVVTkWYNRFjwbm/8ZhvE5pNykrllOF8d
DF1UqIqGhJAbGBUT9dqIC/hUFIbxRGH0BhNaGILc/hTPUPNHCiUmVjJd0SBwAYZH
Gi1aiHWO8V4xdG4Yj5iurj4h2UxKarfD9jdHSNH8SznOVwCqpAKn1+yDrO/GN8c0
tO4iziB1qetYPlwjB3igRC/ozI9COuToK6jQXF2tFwxoTYMzCMfsdT+4jNCY6+tO
xRxBtO9jHbMHau1raynHrL2oDhf6qGF8kkumwWBl1VJ+/uHOcCGsYNYjB8npqdPo
dCbPhXPig1vJG8yX8kdRntwjj3+NpU5mpmiRF7KakJDmJ+VXT/sV/cMt5uwDtAS3
+ARfRbYo9b9cFJkzbJMWKx8hUzR5zGZRqG8pIumdHYbwkpdkPOHezVt4u/nuMUAN
hFPqGNj3Ht7fO1Rla3zKMe4ZzGE8TGV14wLgcQ7ZPUbfhZCJxktQdy1N/7inajrN
rU1WRcWMwvyKoMXlaJMRapGG+weJu6FHI+KNpENwtVgAXHMcwpJ3VEkszLXumq7o
6UFYM/2Wc+D5P5GJIKSca1ei3qyTYtv11MbYhr2XrrYvIKAM0y9AwpoiaMr2BDdK
jnzq4Cy9T/tLZskKBkVW41Bnvn8DdNKWj14a/CMWBev5p0aQFiv4NQkl/nvXwkwa
JPDjr5pmGow/InZag4ipMkMqo15Zo4MTJvGlZ4uamSLci5NxfwOMWrheyp0VgqK9
hV5DguUNHk9dZQ+gZP0F1BDky4HUPd1zMC07DXaqwRnGdgOXj1fbX7RMEdkjOyJ1
QJLGMpNYM5T/9sKA6lUv4Jd91H0FFbPGouaqMvW44L8n/RU6Jtvfv8FaWp0TiQlh
7RMlcqZB8XZmensner8Pp8NhPsVYqJ/T11Skp0wWQuYOJUezoRFrzee//eqpsSFH
97HKprbdpZ07GtB84+0fSCB9qKhF5EBrvDuFBTpyFkFMhJmD43tITQrXPyc/EHFe
GK8Vtl27HrrUQIJLP/JRXE9Xiw8vtqyMkmPfwkem4c2PXlk9V/o64KyAFFHEazYT
FcgiAu7zaTSfCGrn1X4spWBwbML7L+5Lpndl5AEhvDBx5hYtd5xOKXNBMJV5+bae
LvGyywhSz5yg7qu0J4fAVnK5+9mVeN/OnvNj9gd8Jif49g8uJB8C6f0VuM1EIpSq
zc53zK1zxBKqR6lPxkxgUoS0T/xiq7t6pNYTpU+eqwOrrCWYgHmGhvx788DRuBSX
f0zfFteLsRheDzjpZYBiVgwUfR1BtlLX4UWrEH4AncPlEK12TCu0OxfhKUnY8+ZA
DxBfrYwL5cbNILiatdia+NJdcADtxtCl2tX44Y5c5lrhpqhOZgUfRHfQHLhNv7eo
0G2foead2rYspQfn9bS5cdFVSRqOi9b6HzSGKh4SZiGfovSrULgwFsMkDBaQQLGo
Yj0RM0DuMzGpZOFB9osRM3twIhUIVjpMs1On4fER8sJztr5kgWT2tBu/OMXw5tYE
88ggFzjMdt+dIdenjO2h9zmHvrwbv8ZbuTe++aflBI7kJxWZdaj9uuRThCPgg9ZW
uNwB7LK25RLAvGijdNJGzIwqRrusUe9mZQn01ze4czBOnV8cAc3tEleYd/sr56oy
Sj3bULHIdJvmsesE6pxMdBbmYZIimBaeQd/UPZSrKLzeZLEB7Nd20MJUYzVnNt+3
u1LxP3TGeHst4rDCjrk/2c/ZrE9g5A5yM9uy5g9GZ2FjqfylwoPu/X37HJoWHywn
Eslq1HqZga1RJU2AAJ+xEbE3AnYPm6YGfAQKHnie+4Wsi7YLyRfJz+gCNM7FweNE
FmnOGCuD+v/qjeIVcUaLZydpn34lUb9p8jumGP2UEyd/2Pp0wCCicQcDAUS4gnGO
6Vee+wE6YdqhM/+xnZme4vNU/7H6bVzB6Vw+T308ScKXGUCynZhHPo7A26/nAgFV
GMe8vwmXRgU5ZHLDqnIg6cn9NNQGxPWG66lYON++UPFlRO8CGb7YK6S4+K2qbppd
xWyHGf37wjyQxVZaW0vG0FprOF3AFTlUj5hL1eh0vUK+t6sVWCrZeVIVFzEoinEP
lY9Gx2K82Ft+6tgsI0j8qo6BFElnsjRAH/pGiblA4MzPxe9uoeHCCIrA1iahdg77
ybm3j9Q1jlKZMHMbWtxuh8NxpWqVfrbPezKhcqWvpAiQtcYzSgBPI0GkRqrcmcd9
NUK2YEuo36ah7b4HYyqtx1WNRuT8nE7/PKEaxJ2CHPGJVwY94FQQrjFcbqMIHNzP
HkWQZO2u8eQpMJKMVgdFbFjhq2Yh9dyLzQik37gadCDN02fojwmaZfFH0p/OJ5d0
7CrYTEz1pHJoZcL4oA0twU+W6XjGO57oVkjI3vPryEA4PJXNegixwUkAjnQA14/0
1VJn6SSalzuPl2pBlHprWc4YKdkWs+NOZMDqCQ/5rhwDcEeGHmsFhRJyoNOtRh9B
GHksGruGPkd7W+NQM2DUw3pHDkU/TlCDNBqV8e1Vjmnb9oVHCZW0p/GqHrJQp1DH
bosytxDEM6okL4Vn7wX9zwjp8egEF2M0Cy1nv3GnbkYoRBhOHVLB8QUlC6NPSDoT
3BpNzeS8H/BpsJPfzJtFPUmEfm4p7N/nBUIJQiYaxu5Qc7cnxi1g1j8zfADxBaid
sBMUhl6s6DG6zW3sZ/B+LNiLEssP2xkVAJe1S1Z7wU5jPZf9vBVC+upJ29ZVwf7z
glYczLL9UdvIEECmLse1H7ZQ2vODEmNsQ0po0Vb9/1nPPxwVThqktOU451xxL/y7
wJDdl1D3b5cToOOCU8lWWytxFOFD7iMF3HxbQu2PpOZ2NsmQ5dRBIPVOYfm3NPOo
Thyh7y8+UoGaXfH0A3ew3zKcJvjwWIoUC6UYl0EqXJLS608G3Iqi4USlb9hak1+L
27iV3DL2ixtRmSy2s88Z2xu3vx2XFtQplL9xj0JASnbwMdWToXWFWuTR9xRG4w70
L7puuJfEP+j138FMyTVshmpzEaaYClzIP1ES7OU8aeOTkOtoqzhTcXYTbi3YTcoj
ozFHqQYke96YWLP2Ijs0e1hEYFgWfTwyXB2OSg+eNmzVzp380yOgA9hRQDUC7qJp
wngLBeWOw5ZAYzlXP3GgCN5PDsBkJH+wu8YCFrWwK8VvJGFsOKglSE2jQZg4eeB0
O10jR1qIXnM1jfM0uIj6cmrcZeKNQaY+r5mywFZHUG1uEDq/sKaQnkMjWZGjpZKX
jJ+x/WMcrmG8ZdCfVohZY0103Hb3xtpux9R++zI0N1ZE8CQ3J3kHZCgnf8edlr4q
fOxz9uIQYTst1eKX3TT7BXib/Nml7tAK1NTw+TPlFD0EHSO23aVQ+786BWVGiv+c
1JnYaith7HjYc5Eqg8JTOZL7o0H3sX3woKgPU23jjL5+2mxf3BesFe69tcd4XrLh
7/vwyvx2kNaCYcSDoIKyZ+fyK3jTN/91lUJ+F+nMaDtd2FHP0srzQSwd3Dbb8C3u
IyqsHS+r8el46F4F+OAdpd+eSc2s01AWk/rU7vISe2xLX/YZVFFGRqFs1R8ydeM8
H8P8AJLVHzt2qah0n5UdhDPY4JdzANe4YOiiWXdFCL9M17Y/MQqNwdneajpY6chj
OXFFFk0i5Vn04UztJ8c4gNwfMXwty4auHiDRn7WwqSMK0l4xBy/h3XVb3YKZaTjb
7+Jv9B/bozzLpohdNcoJBfrcq8HZJwyZkRVUFgs7dYazXOAvOEBh8kNvkBfKzmU9
i4FLewlRT2zzPPXr+WgxfjmG9SK365AmpDk6efxPiTNDECRmS1c9M+PtCx1yHWET
Dcp22Q1AvlbPEUagMjlSRIDpAH9nqH1wCZqQ5x7vMtlc7nV2sb+5PwWDSk942OKc
JEwIEYBzpRUs4CO4JNNckRUxn4oH3uERG1odufIE5m2SfxRWkpMy1IXtQWkuurtz
I5ArE2OCGPFdqEeD93jkCHylC0tb3MW6zZ+g7LDcr3Ye29CmJepXtlTqK8EH/sw5
uNvF1kwk8mIgAjLVEV1blI5q3BJ/XmEIw00Gt1LL4B1CiA80ttERsgKjvzZPNUFD
iHnu4gbhjqajcPuIxn85XUdpTl6N0CCYnhj38uq8zaSF1qXyMrPjt+NGrTA0YRI0
NGYOv9doJXBSXaQtA7OP26NInCrS2shRonSqWnP1fVvHd4IXA2zCmA11BiGM36q1
+AkDps9kTiyWoRtwRFwyuy91f1l8JcLS6PZhlqMyqGXjxAgYO6PyXvo9dDfJhsh+
6T2/G7+a00vuFDkS/VQdGTmbRv3sWYSqExJC58k5Q7Xw4b3NI06N4dOFtZ87wM9X
aaBD8lEQduiWjRtE19Q+sIxrQQKIIyWMr4jCZO0stoFw+sYl0SdzwQvEUL4EkiOw
iY5lF12+apoMfHbsQx5CpweWJBoBVGHKVbd3+Z9EeyWb81SVXNI8nx/xy4bPRjpX
00t/wy5yDMniijfedyRGyezOGdOPoIUgHwpF2kAmN3wkpdtqWiLh9BkJQ0CvJXHH
zDoJ7YHYgIybZJr+jgkhzw8MANxnvJbwrd9qQmflMbyk9x9tw3glXBN9IH+/iJSS
hAePTA7EtI2v3IXLajRl/PnsqUc1jcMRh6SVkGn2oVXqjv47sKzy7U5vnnL9SzLl
fbknOCI2NHmp0ryzmDc4A1NAVBpvgmQy7xFf3g4yB3VqR+ej4cfYkAvZwoJY49aA
FXffESBbckZk2JkV0CoLvTgTTqbT81OyudlG4AFoMhlq7qEnSjSrasWPbh/OsSbE
zgaPO6cVBlJ+8ECZ56u9Eez9MzrQbjNIcbicuh/JPj6il3WDtDuG4eD8X4X7ovk5
8itkB6h8u2zj5G5vVTbDuz3fwcZHxrPU062gKxMKg3ypOXVB9+hSDaS93JCc6agC
mYfZvD0ljy9xH+GxdCE5RpvgwVov5Nm4dUhEDZ+VSbHq3KD5tlGAdhxaDkO2N1Ze
RuQBeVtyLsoj1QUP11LOUDM42dY/BAFeIM1m2aFfSYTj+yTMGXRe/4FpaFJOXTdF
IiSRFmXUfZn/bX25T82HJfPhQ0daU9TnRMtXOEEvvnkVjTo6ViENf1lFFmUkQyx5
gcE99LYOdP+3AjKeIXlj7coegP2um5jNWmhzmSsp/Z09SdGwyoqRO3yxK8guMSgA
4L+MJPYftTJGYS8Mz//2I80YTuBMZ4iEHMQXbVZ0PVCXtJdxI1hQuWTmzL9cdSyC
Lk0xbGdZE7tIpZhIHvhOQsCUgYEBPZxePOEhONweATxZ6OcezNmi+LWwc3DaZ8iT
dCcXQlpo3YI4Hh+UVsM1stDs3DT/79ccyy8O9cxqz2Cn0Pw72hdXnUrvEJMVoXmC
d9Dsph2jIucNZzxq7XrK5jTjJ8QBntHWtEtqDkckG1LSd03YvTm3ZIksbY0D4GCy
ig0EJIa0zUjOHmFp/jko7T7WFBo/58OEfKk73EJHyuKJMF7n2CwdeGuxJeTh/UgA
yS62w5iRfasGl9NskphRrtRaXWk9+8sWkGkoa0MlGXHOtUoHHUyAuibVpc0Y/o4I
P0Ho5dXFpHfirg8IV//vdtIB/G0eK6OYCcNn8Dk0YDiT7fAecN82DD/t8IqQlmSn
240lNRvp0gbitOuVNslfsOBFGv3bheikvof3cLqluOw2dDihbCDIl13i4u3IjsGw
1af7fMx+oYhMwyspuq8UTioOHuo5q7FESDNhihQcjS8GvPwQzLZAKf/tP+nYpX70
n15JjiKsnZombz42HygDh1Ve41FU8jltCqG0iVbBllWnm3LKTqW8InOXFXYAX0vM
Y2OzsMXkYVGKRaeWUns86Jh/f/BkS1j5Yalq4395yto463ElKNV1kNAqsqkaNuV5
ImMTiTgPF88fO0fZl/RfJPK2l/uw8zwzMdHIViYutjqM4J33/dEkzggEoab3EKbc
psS45Dms1ZKNVKo17Leg4l3avQsZeA0uHNIdPvs3Mdnfd2bfti8OQjYprzmngV8m
hdyI/xgMJ03eywY8VS4ZJgT1I04lNu2TvwVjQ926G5cBuetQFE3hzXIJ3lh0UIjG
ZJu8YD4idI3+OGpSmiHLC1bUipN7V71ZLNYI+vtSe7+Fu8J0wjzIPEFjdqKColtg
r2vK5lhZocIYsjzMoiZrMSWCPbJl7HWcyWZPh5amGSm5N/iQqT/PclOBwu2YTvBb
k8YYOLd5LIZzCEuJi3ltGakdI23MNfRB/nvBXxSiZ56UoJgnVp0QSd1L0izXtGSB
SuXC4ZK37p6qKqhleBvqafRVVuS4LgBfwMRLUwGkptzoilz+LQp7DMbx6O9LPYFp
wTGUjw5DcbTpX9/emTXI9ADAoldezF7BZEp2ajsWtvQPoLe3Qydwtu/vxmowKmjX
fcOduj8VxvbuWEPV4IsvZFByxXpPhfmLaK2QNXqAwa9Ec7iGLOkuQRNO7k6lEFEf
rRgbNfvMXHURNEzDNvZoXYatUaUFF48CPfMVKP7V3dGnQlKkx8teNnQjoLbcjBRX
ZyGArZI5Wahy68Qy4qwHUiVnN8AmQXUn3ESZT/1/XAXyITKk8WQObm4yPG+AgZOC
2zb0UDb7J/w28pd3/VUVU+1LSKFR9DRxXMyAe9G9tH5MtuiQUrbDCQyJK8Xns9Wl
PBHfGsqwudmdwn4XYZ2tbymRtEQfMLJw66E2EVDGlo4WWFuurqFywMmMOrLdfmN6
PWvptfoHQCF9doOv6zsvgQMBGXEWc5KTcHDCD9m0YwaqiIlhdv4wvF/pz1RlGjkT
qsDvRsw3Zz7udbzpsd7Eo7GXsmogvvwOwhmzrrj4YQrScFZK8MMzAOej24fQ1J76
Po3N8QkwMXUW/gVxuqoiQWtBlPdbY0plUx0sNhVl1zMwQCpGiJPq2YxgfBa5CS0h
m6NWOr5iOqX9/gJI91xxvRISTEp+H6ce1rmmSdeLV2vSA3BiwZdCeU/nProEdOBQ
MUBeQuCjkjowk7c6640YDX/pp0QNXUHDS/DxaiK9cQlAkjG8FUNcqTaH4KHLZCf5
cYcDG+4PTYwC6O/K3ToTwAesJfTpFK0vjj5hbdvDlcaXrBU63R9z2l7qoJ/LiCzb
rnY6686bdne+3Imu1D06m8N+7DdFq7wujX8KmofBMx8jF3FBj2HKpo9XLV0BBMzd
pYCdS53WiZ+x5LBW3Qlo5pIuTHbTbzLHDA7IYntT1L+Q6A9o2N2x7JEcIEPxmYtM
04BUlxLbjlnii1oKgq5WFVv/Yy0Jdx6aWBQUg7dNywLE1yCj8TmB6d6+QMAyyvda
gLKGYRiBKgWJDOSKAEXCxmXKkTqgb9CC2Gi+x1CRkDzFIpSbXIfhPrYBK55OO4WB
YRQzeYPXCLvgKYTEetM6eypn62MV8dD8XgQf7taFfDZ3WSovKyGuyquej9QopDu0
WbRwLjoqUc3d/XbImYPq5uWDNKcnsBY2TuVbgUmPBYwg4Jw/K91SxLW1OzSQT0gl
CWdR+l90kB9kopvodTY46OrxOMtUlcy++lYM8EWbb941gcJcuvNWUc79H3qvhRqP
t12pzdXmNV8KSpme5Q4DO1k/wt2BLma5adrNYGwJSeTbgxYL5NKE3G3xqFDylWfI
vggaymhVsxIc2M0SEbAMMAvePGzwrSjbdl0w8hz9PBryn2X3VWeOoWj44l0WAF8n
j5BVVcVYJnZMK/HG84cHyRYjoeJRaJrQ4X0/zIaaauW+G/eKoCi8yntIqBxkUvw1
LIHZrElsJb2+tGhpk+kzw66BrQeOLAfn4KIGIywEJGFvOMpIb/H2CfN4I8j0Xy+V
f8w9g9OTwJlLC9yl7aSqj1hSkDybXmueIgBSso6wII/Dn1sjYu4f76vBhvom1aSC
hZ7cEOj5ZNECSd7DA5dSQf82H+ijDZrpDqxk+LRBbRYdtV3VjIuOohYAE3s6gQqQ
C46ohUq/67EmfyWYpDshYiWwcYhJS/1YzH9zNIMQlvKab+LxhGafJKXmG3gROVm8
3sR9zrFdSz2NsrkJLZFSsABfxPGsUmaauf23LSIqdr5NbU6/GEd8hod7iZDf7lle
TAM8QLxDjzgZbKv56yaJ1XLVajcmDRSx5jsCM7aDyWxSQhvRhpPKxfz6idRacNpK
lJUcxXfcb7Eo5z5FRIbufj5to6Fh2oZeNEOs9MHvRqcjJaDa/KwjPxvpIFMZyU+g
NECy7jLurKCJjQybhcN/HPwethzIXWWUTQbsbJuFIZviX0rIcDDAeTgxiADB1obi
pToQhYmeLRITzsCG97A5yqJV/dqxy7nqIM64gNzNhiw7kxWT5zPvPQV+RZkwaPIj
0PsuanO8TDnt/kPW0VLEt9Z0i0e5/K/uVs/ysfAuWDFyOCWOZ2ysBFFkkWt/Ljl3
Qd+MGBgcgJnV/rs1PZZvkYnQ14PQhGUm+japH0x0b5OZmIzFdDur+J9BDx6urf47
hWY27CYeQB9+DGtssWTvg+mTitRGt8/bE4h+A0AGtVkPHNH6YuJQXYD2B9Y7KlDv
TGWJuPl57kAqYEjbUVcmgt9Mtme8/+MEn20+gTgLZ/PW2jrpn3QU+1QlkWkndJfZ
`protect END_PROTECTED
