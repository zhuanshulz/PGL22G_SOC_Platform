`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MROhhEhokt6Xj1GSAC8oiJk3yoUQHbtKCb/OHEUCWa+oIRsDkPRdIOA3gCuq2srD
hoRcKLx5oUHb9lWY5Eq1unxOoa60zCDXxbpCd67xDw+qJDqZXR7k9O4FRktwFpMe
0TkeyjSAGs/txUoalOa2MyLxV6C39Y5UjUd33EfoEA++NbgKQSy+DlPcW7ERkSUn
lV2U/ug9DfgCy/EG/O+PfeEd3EU2OEeNcQPuTWSQdAe+SxlxPisNTte8lLsCWqNU
jw2R0IahNirWzZWac8teEaSBbhsbJ6SBehsalWK7WINVWJoku1NF9tl6sGIuqlBd
n9hnhj/foUTSBDzmIbPV67n5/RSnBfxNA1+6JvddV7VKKkRzMk5xa4mMWfqKHe1x
7+ZzoKlnKV3t+NxWA8FqiXJayWp0n/1Wwor1kfd+dCm8xbMS7alO5b8+WIFMqHpq
BNLxZ44uIT81jtaV/v5eXDxjiLHBRP3KHKO10gZfSwno8yFlvT3WmJpYUTBHk9c9
m9GEYN4eitUMMFpkmW+h434xBJriFMIiUZIFZqU6rsmDxS8C5TmpEjZcufbuh6Y4
c4YnZJV30VPk//e101q6/YdKsSlacgGTFTnxZo381Ct1EE2j7oOZRo5XCYzkROnU
VcewqYukJyGqG68Exz3qbIApB82MWqM87fusWi+dRUJlGNOqKUYdWivedcLT2g40
8MXRkjK73nFd4oZ7a1ROAZOc2WQfY86NqRa8mrm3AczQjuye91iTYwWq8TsIWw+f
a+/lTW26QdmKWoP7hlIaIHFiN5/kcAaVSppLhhYUo8U53Agb2D59rEs+p+sMXKos
dyUa1Z12ULYVjxKwCD7pu2fJU0232vRzBqWigbR0DASS1y3Ttoth+RfQTfh01NhX
ORnNhGhzwcLNNicstAOl2Ax/geTKNv5PWLnOeYPE2lAQ8vPZQ+JmfMLru2MEdP5i
lA0y45oXBJWzA6Ar7zi2JZ290xPvjtx4IjRdY/TykUxVtiqbALzucsBU7fiV1rQc
3qtkHG3Fl/b5QvmSiI73ZAi6CScQFf2BmMEatMLQyLfCDo8/5jbiW3KKBFGbvFyV
sp7F8WRMA4JIj2ERPG7nu43EYLqHaJnq4N2pc7irpz/6RMcvi75+uLQPRwGW2qf6
N8BURYisIYk7YFYKL6+9dJqc90rtxpEDUECPlI63diywptDLAB4hn919F8o0lWtn
qX+hQr6oTeA+W5A0PjlWoSLE7WzMgt4aX3ddufHQDnsICQphYv6nHm3IJg29Zqod
E8J1nsLRsd47iYih2ooOorUr6jxn7p6vkO2hqVBzVsjz47h+9J5+l2PVghriDEaQ
OQE+LI7VECyOANhySrk3iP1jahdMXPttd7J1/+2kVcaQxTJhBkb38jHAdi+4IlKo
cASX0lUaT0FORbleKjzS9zXBRX+0Zib2BCFmmfXScyWVoz/1cKii/A8z2p//tpup
Db1B4dfLBVu9X7sEovGZ7oOMUCeoct0G/OsxvEBSTqWs98gyKv+NEvqUszn9airC
MtopjbZZpnYgCOu7N+UU415G8pviR5ebWFpEaCxL3by1qvdr6jjO8XkRD4bVML3r
ExjEEnAREU4WdhCf9e/8E3sQyJoqspb/oOTgKY4mKxj9N7bp5teSSUJxFmbuE9dA
B5ORcFTcqIgblGoNHjuYizDcooRe+rBpvEx7h4BkDMMpJFD3AQGKFk0k/iPYp9pF
sluJwmgdqGvwwYOJ49pCZvsFCQL3RUSWRWucmVw38SwoGpkf1Ndj+GQNr9k1fgMr
nnCK6NL1dlwcsc3giP05i/vJG7EwV0FInkGgdqwJKtcM9d71Xt1/4w+JBA9f2jtm
jMMjgOQfBtmkgzoGVciBelCKl2z/RJyvgB94/JR1oJfzjxLHNGpOQhIC+m7RIJ3q
8fuf/4MmCd6NZ92Xqh4FBlIYuUwkP7JKil3VlU9g9BZhiG0GVIABNGYQFUgjgV5X
6gIm/0e6/5rRuYmyb9hBSwUuIupxd2caGnw5hGuKA7lZFpZ85WXSe4Oi7iudOI5J
ZSjc613pzzzLxq0SNZyfss2J8PZsx2wD9CSbSM8x9Uwsm7l8ZM55KaMO2vtT61i0
dTVMNma1qyhuqo3n2AvPkATzJ+vur8r1458O/qP3bGUm2zt5iLaGQvle+Aq2LAbo
hTsA8k6uCpKPt00+pyxUqpsd2d88IDp+InsaA1jMXVx4XB7mV5zUwziW6Y6y+czT
eSIATg0x/HkGHaPJAHCHFHzmMknwvyjNyGB7s1ASi3RK3GnIzx1/4Yl+M0ZOqrZj
2jNxfi3w06XoWux+VZNo/WO6HzGu30kQDQew8IzEX/Nye1E20+Z/kmFb9ivNcp3g
zsRkLMSH2wrhb1WMp6FCzrU7ZT9pVY/QknRDqtzvKn6HvNiHu52/faLkWDzWTRQJ
JEsxmXtN81R8RCqL6IUXsb1c5i9JSOcGd1W49gAxEuQiL9tgY0gvljh5ji12mQSq
+xRRGt2Rs8+g+Xh5FyIDWWwqvJRmTYWjF1a0yZ8+q/jFrOEwde3n9cJMrQQFOMJJ
1fl2YS+1iNUdujLkQ3Bct7xWJirRoI0jQrL7SFHpE7IHinVrry3JulDDaixDJM3C
k+hp7SSoKb/bUBTNCAu1MGWtm3Un68HpcZkvVW+1z6LY1pdjtcPE8O9mKgcRihRB
QaS70AjUORrg1uGplEcC/fJOJArkz/eZHTiBZ48Z4NfW5X1rSu5wHEnozlWrrpwR
E/c91giasuOCWm6lmXcW8Ucwz7nNvv7U/si/fXbj/qz8T2gPvIOtRczrYPtezL/X
bBzEkAaIGnY6cYhbhJHKk2iQTqiV5v7qXJcH4a4/qs4auuKDeIEq/x2rQxQ1V9iQ
uYxXkq54SqG7ZwdBF0IXdeILI/iq2r/I48HYyfRBP26qX6D6fn5tRQvzofoqkv5d
n8XREPrTmdRAhAb/fy3D+KaoTcz61hF3uiIoTLbh2jgNbLhNVosfzV6xDOoxqfti
SsnxJSUp6ACVuv4MlBLbyHF0xqyFWGo4VAlT63Td/6xh/E9ol83HowyVA1qm7kMm
ILTQ7FLAs27NuJ9P+fTsMWuVzfGj91t20JNxczEMgbIkb/2pz29hhGn7BnrVsnjq
8u30BGgsbGlZhuNJ+gABM48AGzfoYJXAwLgWDwhgg70w39FipQ+9FB1YYH0AMeqg
JeoLXGEY2XkyB1x3MDJhGwTNhBPuosguELHmukl08JP/+/e/Aykz22OQtHDj12EJ
eXMa3kiQ5ifCTFx7tL5lfHUjY0AGlpN3/4QpKMBJbUbb1nnfQg3PYlJO4bRaa58q
+gsHwcP3FHbeG2kOX2WsMqey8giNhqnZLeNI4v37kty0gTEWanepsckWfaIxbDdS
B4Fa+e418N+MyhaUOGq2GHZwlhmUReg9mGwN+1F3dH0JvaI2vMbJMRZdaOIP4Sgy
whT5M7nBAYM8Wv6IN8WG8gZTo64DKFm6i2e2ENSatbn7J8EpMMBxurmWBrqK8etF
pecTIxMnZpXy+PayPZMaV0m0C3dg9SUz11ezfWxJSuxpURfB4O2a9NlmMVZjbFsR
ifrvs5g23o+EIKz9KWlDj1ZSDvm0KZ1YfvVptqBFSDr80+hVlVHKYdIA3POnZQbf
x9Q9wywUimabb0mQWsf277Hi+9C0xDy/1MkUJL78RtoXQF6FMlfrwFanVbmDwRzJ
dSJ8JAZ3e+q3oN86G7h91oY+lRfgTtKAcKe2aFBFWdAVIY1htQRzshufNNrfGzXL
h60JUS7EQwq1EP4JU3uOIVK6r7ZroA0GEoh/fwdjiQwJYjTlPdpXQfoJvFG4VztG
juWx/C1tcv2uHxSG6W3dGX9pxesyXHq8S/6lG8mx1VZuLnZaieaKnmobnkkSvjVS
9aAhw8m5A2Ts2BFb79vDLAteAH7euUmV7/7+I1ijhDXiRhUyoy7BaViCejs43urs
dV0jVTxHG/3ZyLsKzkj2CukbloEpdMokpQqyD3YAImPqMbz9oSYYpx8/9xW0M5hD
SxOer3fIz4ISq2+AUw4MpKPIZXBckg1nxMNMRx4atof5MmYQkBqzvd7uWYxOaj/h
F5c5KiwHgyx1qb/037ixsJ7oNlJh6nGA/8LL+aWP6/EodqruRhj0oKBDJVrZgtR7
ze5g1sYungZFCgft7sTSrIanlkbAwpje8AQnPGlzQWaLvy2tMlFdxEbjtzALVHQk
DHYYjbYUiaxMehHOKTu+Hwv0wf3tHKKQywxSmbUA+MsXEg0Cw3GMwIOE2WSzJAjp
ErHPWRlL6NbIjsTn6mmM0ZGAX1UoRom5cvZ1U2qRbt/5Hc1Ssj4D8BicyDDKa7OH
R5nLtsCqB43GCRm9vZ6rn3WBErsOSWTVI1+B8N4GFZt37nbPUlc0M8/Qa4IuuXJK
PGi+U2On2gi6PEAkHvix+4CoEykTnPVvTKoqd2YniQ5LXrOFdiydHUELD4wJAsCB
WAljejwUpp1GV5V1Kq9LVa0Ed7/nSqib2gsJUN7+yQz5nqcZg4DL8vi2tWawrLmE
vS/i9MEqFFMj4uKLpwcKsNgIDmVDFvfKeFw3bOu0y9QuxfXcL7OKYgpLnuL7msvE
c7yafJejoM5VXkFWEso5YIOB29C0Hg7A+8vilZ2CjxLWbmnroug+9AxktL6N3zkF
igm9aO6XJz6YtfcMcJzLRZuMHKzmLC8twwLWGbGsx1N/4atUv1rMQ/af04lTn9SE
HtQnW9HS7C52ZDjvOJDz3viuzjG/0ZA0o3I7RQI3bajXNxtf8vY7mruryD3piSqT
MaHOYSKcLqaaQ4PzIR4tlN05o/rXr/7D+BJMwYmLhUvMUvGCUPA1y5CZ+UZnb+jb
pnUfJt7b+WRHRybkIA1tTed7QGk9zPUmfZeOqazv9BAqR1hfEgslq4h3vP/0+x3V
iQRQIcD8e0el5f/wszvMPPEi7qL32FPf6lmE1IX6Towq4b58pPmKzy8gQgQsFeeJ
CnfTJhanA6hB8QSZhwFE4lPnVZCLiyMVf3yw/5g3a2yKclqjvm6wOwlhPh08iL3e
p5zDnYXEVdiR816dP9b0GRlYCGuj7irV4BjoqOJ9//91SKrKOaHM3nmTdZXX/3cW
7Vf1OYOqF8DiHV7fm/78k0A4yLKMKEbqzVjg3lFRDT/nHB9m58v0hAjkYX+Vw7Ld
GMjguQrBtfrqqbscKVWh03cpp5/AES6/7cWYlwm+Do29wCfK3UPcokb6awycslfk
iHtavHAvX9Mq9ALdQIXxBtOFu1FcNl6RSenYQlzRnuJd/sHhUjuolN4NExCyXXSY
QCT9biuc85GWQsdia/ixKMZe9R/RGuC3rw4D2N//7/SIVce6MWk5EWg00gHNqL7h
6FKbAvW5i/LVBl/lfeRfBBFzfpSjBdZT0Kyb/+Eszdvl1NKK1Cxl9XFEUNRPtKz3
4Lo1l++ry2GFxEqPmiTChKMaABuopPMc1V4nc8tungf+ifUDJIINJntI3UIoapBF
jjhsteRbxuvLcN8ojY+b80j3DnfUL+ftJdVL5t+9ivfDo3/CXmIEzOXhrZEMbtdT
Q6TpUeumeZaGnOXGPJXWLRw3zDLIrpPc2bBbktrwyGnoIMV590yUBp9NPVtuEiSL
VFLKE0RMg9QGC8viV4Rm2dqi+O+/DWYltd69cE2oI7lP1BqMbgH6nBiMV2y1eZTE
TLASHop9OMda0hgG27Q1ju8112r8mLzysRNHWnNNxHzGr0qAm+ShYrrUvItjZ00u
zC89E49lzFTRoxD7C9PmhHQD0lFY9wypWsA1yzHcWCebcR+M6mpTIkXujsViBIGv
wWUWjKIzIzniP6rtQdQKhLOgI6y9+Gnm9Iyhlki7Pgv4gYjB3MQZPL4QQLVCvWxy
TIHa3f1v20nnBPCEbAFnALQf/05cOOtrH7op4EBCrmoyKuiTBpvztxDYAbiCfi29
Zo7zWGVzrAtgyDA4XoUQ7w7IknrW47KFgVSkcxowVo662e3PWq32CkND/8Mz20uY
fHTPBXuVuU14qI80hxHE8PcPRF0Gs5xSmb2yfXZFNGrZSTzluVeEx86LwC1Ube8O
J8vftg47W/yItMUEAl0iix/PHYg2HrVMtgxLjDRVyds7vtguzyOl7twgGNXDM9eB
j1RZNzITiculql1S3caAKbADCvpFF0WLgqwUtGjd9PAwpJTLfST3pUArq5pWfjHR
6Cc38rFgCciyaoeHltZkE2FHtNdoXY1f4o/fAHT50ijPFBPiUIoswqMD0+UmGYYA
tjLzH/us1nEnlW/xTMN/uiC6IeDBu4PEotIM9fQeGm2kXBZNVmdr0Bh9defWoLF3
G8yoRgpTrq3YM0YkoBv1CxBolVcLbjSB0L657iwmwB+v9ad7OjQnPmvbBo/B4mvX
E3XWqlyFpUxOlEhxZAaITd0PJXkY5vrq5oNFehDBAw24KnfSqJedtW+U6Ncqfih2
njMQZaK8a5YB5ULOtPF6L2EpWF3z+Z3CtPLxEoCt2NXkt3Rfxu/BqFqaGTKIJEJN
/6u0dyYDI9VitqVvdFHmCXhnwjjTxIhqp42Hjt46GzlbdMqkxajdKNUAT6GVCt4g
YupNiwEzUh7qZwXSqLjeIdWNGffsnTio3seUNT2aCeojq6zokc5WkzS8Uro+xi3a
ewEFpUqZX2u9C2Wxw+E0oCWKt5wRETYn9IFu3ocHjnboA+BMQO82vWwccF2b+ccP
dcsdlgiSoB5fVoDLro/B3tzl+F3XSpxM81NO0iI0QGlAIMY2i6ZMmmjrLNcFowgN
HZuDWTsPqC9cOVxefUgoutNdIq435k0LlRWGZCK/Qno9szyQjaLYrrUBtPyh56QK
L9c/KAw6UG+aQDU0Vzbc0kgqlzkMM9nIE9ggPwI4Zmz1N5S85gdgowdmt9QqCTLQ
FL/MRz8ipkVVEmxjEAlYPEA5nPU3nguewnx9+7W5gwMv1Ct2dqMCh3+a+SlJtRzw
0gsh55RrHnFcIk9Sy8u/A3XJqtptWWPTM+/H9u/RQFQ5x1fYVtcqTbyiWEcEnOPb
YmYAVWFO4p0a0fad9HzcFFJnWgOgYZdvMu5aUKhekQVBvDc3mPCXsKGPitSNi7QU
f1PjZL/fpvOzHSsA8LCWPhUVTwHbi5aAF0GXqf4NEcXYzeTQ1k1hu1X9TvnL0c0G
zB6UCKrWbACZ/E8VQfI9lCGDCM//gxGIzuIYkHowVI0m2LlZ4hiuFgWWQJhGoMCb
nHWDs1JBZrF4q7yVDQyhp7rqN9LlDQ4ZNEadtrkM+lA75YZctFe7O1i1AsWY+OIB
AotetR63K2GRjkDcq8tITTnN62lea0Etq0g3PoTtjbG/9FFrm6WvLxcXS51lHgGA
bi08yZtvwGWDDP5423P3kM8KOh8Rfd4UpoKE0Z8u5ubvoyQ7BgcM9bAZNuYWzJSA
tnqb9wITSnEeVo22uNEF+CA0vjz48qc7Ln5XA9nOvo+QhMwdJAr9mnb2nxTH1dRl
9+pv1cqwE7HWilba1liMgWgv+ewjlZwW5RcU7+RXXB4GCclS8hW6KoyAQf4g6uou
5m2EB6hnJXhLSwCEZ98njcFPdgK+MwABWGdR+Gs4HdpvZLsZzDTLEAgK3MDUhaaR
Y02nDtQ0UWgINyscImciTfQLiGQTxBT6dQu0+R2hzK3f4eVXvcpb0+Smt4DVql0E
6C6N8s+oUGOIu+hU7IPHZRebUDttn6CMDTAhZFF4Fb+jXEmSTXIFkX1IrywzDsY3
fKwf1qT3jgerai4Hz2MGeOT6zqxG/eTLIopMewshPG4JaxN06yfSbVuSkg8LhB7B
QexvWXis2NZ88/As2EMLpcRL51YFERzWGtk0BM8eYVzvPHhTfM9U+SQ0/y2idnKq
RG2TNzha4oCEXUoPcJod9sc1ecjaDr4p2YYfF6KPPD3iBuFhki/CwP6Cid9/RwJy
0n2J+7jpRELdhIQ4piZuyNhaFeHj0uROFvKW5mZQq5WexQFHtyztTjOP9tUFLeNF
SGzBLZu9byc+aPGVO7tTsjY/caP3gmMBPhC91otStVqQzyrJU5S+ynrv1ZfHreox
DKy5A2kLr7VW8uIZmR65rjkHSPVdGfCDovQ8yOYC9UG9klpfwYejJblpqteXOyGf
4RwMsoMboLniItb/+rWeIC1YXBCTtYq4b2tU5ErqEkgf12D0I/bfjD4XAAZJo6i0
yvfkdq9U38I0FrdizgshsA==
`protect END_PROTECTED
