`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ctuNCKyhn1bGv6rrRe0c+2/ZNoQ7RTTKnLqt/BBIs4qe1wlmeBPtWbcegJjRlP8F
vCP4jkNyeBrEihijOyq9zbVsncfv8nl/9zUOKpLpFOO6u+9CUdEOX+zsFDvtxtWQ
7/dfKzmH8CkLG/+dpRL0iB43ozbP4x9tadi9QMRepY/16U64Nioh3Ej+oFMziV76
Eb2W0YQIE8kpMYOPhgj1XEZ8zlX9HrKzTxxjrhcBULws7tcF6cz6Trdnod0jAUG7
c7/HstZWYwWOKl005Vi7ivBLrnwJPzU/iVKw9bRZdsSyuiEBlhVJ0Vrz3Pwwi6Df
fvfNftyvJ7sv8z7MqHvdVpoEPhgl8sJvu878qaXrWToV1GdiW+79TzXVFWPzr+Hr
T1KODLW7Ca6fH9mSBn5FeVp/EZiQUp6U0tnrKao8Sw4ZRvGy2PSaZwONj3LOs7u0
1tHe2o0aJuRN2SFFBZJuzPlkLmOPhOtOTo6aYaxl3ZfvNn+rORHfd72Wj0UxoGnw
OH/EanESWKdES0kllwQ4AIpDDWYm0oCoO7/B9alWWQjjEP4BoV/JM3NrawDIjALy
RA84FC3+lRa8oi3hYv57nR2pAh//sLJ8YURk/xUDZTxK+LEbzPn2/qgPiF4pZ89h
68ZdDlzcam/+8xFqogbvWgkH5HzW7EfkTEM3Y7rX+ZkdxHkww07Vz5Z1Muw/PxFG
8lNMeyHVskAV83XIvsNzXMAevPMv20MlIv8/j99+N3I=
`protect END_PROTECTED
