`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ziCOdwixLQhfelF2WS6EU5TLXZB6mvzFyuFFS+ClydbhA3q6hxoX7kS4Xn7DQ4eE
PQ+3YCVIaGI4vjcbwsezpTqCCke2Zh4u2AtjVe8xCRDWXbW+iyn0N8KZ8aDNB1kX
9W9DzZJBxddzS4MEIAI7+WQ7dSnUccR17bHi9LLmNnBOTcBt3tOzYHhGw7tTdsWk
3U1Op8sgWAhxM6VacDdZct/3mmOXPkRH1ik9zN0LUSqaUJyD4EKrxFA0GhdBidd6
aqV+ZyRboKHSt0RbYh3SGIaOAuWJE2DEe6bEOPZ7CJX/2Pyqn06zHzX81lkwJREF
4dh9zeAfS9MF+/GKCYQBZAoDvpew1RccfXisG2YaTk2dCOoQuLD9HbczkY1YDNlE
PqWx1/51TDJImBUELj6pUlpL6ny7SSbQj8BpWC5ZW4l7+u8UcH2aJ9MQ8lFzlZoL
vuITvoQWi+ALmS6h6p9Urp0+AVwJHaHVyolJliXIelelqSUZDY10W+cifigL/yEg
Oiyp3IfHAvYew2JU/IqazHUBhMvrm/zoX4qnz9V95nGmeuN6GLiIv048UlZuObV+
xlXcQYlIwDQ5nDjSuCGmFhpHpPREx4wPddQFfjHNhX7V6rnpBUCN6SvYHqYZCzY/
ek/2kn2Lr+NSqvkqyhyO9n3AF/wDSfXo5/rC1JSkLp7lNzvNlP0hlCDEUnXB7JV6
Y9zqUYY7tNsVxhwEseb6s4MbQgP3cGogiNkIfJl9jdpBzMZUsGdDutXT+ocrux1r
cYRwETR5NntzVFZtJYB6zMcI5nbFvpn7XW6wCR8KBB9vMCAQjk+WUWRVU0KhG7em
wJpb1dJVKjjDLFefem/NTIH4CT66WqX1ZWqny8DAI7Qju+XaweifwQCcA2Y+ykf6
DtSI23YSnEo13Ha5Vu3qEEMB08T26qf8Zi8WeBGSsqf65tiKGY8D4m7L75jATcs+
Pw8E+n/osAD6YnzJlljKNg==
`protect END_PROTECTED
