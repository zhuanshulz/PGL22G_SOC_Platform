`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hwBhYZLgfFKKIF5WT7AjQjaitsMI5VqYc4SaSOYfzbQpyR9mJ4jaTAc0/FmQVtZg
paS6JQRUFI+CQB1QpL2RyDgqlUvlFL7osUqyl7wNwfenyiy5/JuzmooKxe5+iNDw
0B5d1Cxo50HqHtsqUgK5PVmz2+SnWctMpv9bO5JX8s5bSLcBYKFIA6lHwVsUh1xV
CRNLNpJIx45wohjaQcjC4k8Mg5vrnKWqN/p2ja4vhAz7tU0raclQTd89cmHD2P20
jrDYL3A1BP+Oz7/iL5RzUIInhyoEUt4aiodWRLbZqkoiMagWTUNG5LR6vKXzOrH5
91X6oqK6r9G+OWxxBYdVJJ959N6g1DnpS8iO33qLjn4bzBCTfJgDlKVaj2IdeFFt
bBo3s6Dkfpw96X6wIITKyNVTCKqqylQPkZGn3YcmwETePly/ffrd2mPGkdDfsSwl
wFVUCjq9dIRXGYuHfJgpvTL26utabPfbauJy3ZQ9u44RoGns3sRYtToRF3/2deBM
rnpnSiW7gCOEaXDZ2HpWOykVE+VSDzuqaeAPDYhoXow/DUeESxUCx5sfm8HYctG9
dVSl0xpbCeupH+v5slBF1pOjCmz6LUwKkjlzjpVV791n+FcQf9C+SKOZFRTr86lW
V++Lg8Pj15wDMuXvurkhSIX+9+oCxTqFBFZIepo4QjzL/j9xfEk2pN+NqZhK8c8I
IZKPPBD0iiEqpWLCNKGjQcKAAjGmYpL/g6Qsni3mfE5Qw2+eu44U0q8KoAitU20S
PDDukAghXJC2bI7fIs0Hy3TCMIMAgsF+t7WH9OiRFLxqq/fSLBuzVEBa1XS2jF8u
+tPjWyNsi+V3Tft8qHNT5uAkQdZcRlrT/S8zuBRVfCBULkRcOSHAEgna6oIV88KI
WEInhRhDpq5GNNTeorpJCGzYMySH4K98my5z68TMzLWZk/QP5J+Vgi2WM48jxEmN
0b8ZrIquz8NYS5mQ4ttojyUQna/6a/FlVTo8mcJTTzEJVjS4wfNYEJ/ihDNniv7x
0REaJAnc773PyZLcaa1kGXxNZPuGgzUQk1lp/IsrSHl1JBIE2OR0LCW3abe/ei2h
e+DpWVnL7CdsLl5jFX0wt4+tQ4vZga5CnPKj7p+KnhJk+yHALkZ6vSnwBxfJmvX5
W4Uvw5KS8umhe1pqyNW6Bh8LXgPhHXWTMRTHsw14yIiOEyNkolrFog57Az+7Q6qu
5k1D6Vk/nT93FjS2WeDPeLR5FLwhifYVkhBctVKJPuK/n3fD6Qss5aHk5gxdQ5Od
5sIkFdOVYUiFbdZj+/Y2WWLgd4MA1c5YgQnLrlfwXOg9CGY/eHk2KiOL+FCHQiTX
xuW461x4/EjOekHNWlGanY20Gc65N4drIQuHOGs1UoSdu+N5M3fVqk0l1ZOA4UQ+
60MmaFQZkqpcgsapIudcb3qEotp1rFH2dO/jORTU25y3DqGoLlug40D+CpWjt9PQ
RrHr8WGMDVsGXLshbDzWvND1/5SffldtB+Si/1RelkHPSYryIcbFyG6AYBev9FOb
feMxEi/jvCzGaceEgYGtnJON7tTwL73m2L9DFvPdmEOtYolWCZ5xyxJeP2MruFQz
WsdtgMJsfCKY+ypsUVKr6uZhhjS3z96uaO1BIBWkgUM2NUJqeAuVJIUY7KSf+YLA
IY1CNv3+yTkhpTJORnrEATtEMWtFMUT/JninbuXQRTGih4yDnHgE0UFJRdBZK7V1
/Tmg9lOYF7I33aJHBm/s9p8zbLotvGx2ryx/VXmOpPvARSKIdqUQoOMOpi8d4OqF
KBxWvfRYW9Hfy817oC/3cF9yiJmPeMegzsqX8FLQ/2lAPw5iWPWxxMrtzIHoUi5m
xPy40asLyyVwG7Z89J84T9XbkKEqy4PccApnVgxK2PbG6MErIYOTzgjuypi6eXvJ
LCGLJ42xjsvWM2S+wiiMzIDrA6qto2kI3yxVzUdtdzM=
`protect END_PROTECTED
