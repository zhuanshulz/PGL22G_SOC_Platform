`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GY+GHb+lKAji2xGNB7UseAdtzEO0ZKoB3gfdvDy3zVsg3AsI+hs6onsjyMeqrk6n
4XcgApX3qvuqw/t2b8btBPSRZmRZ7vbZ+JbS1SE1UyqMDiOKkqfpKjrLocIirdkX
6XRoVLNGI+pod0Qp7op+IK+HTLrkj0nbcoy7cbMkqdh8cYtQArM1W6dj4GCzE4iz
f/MhGjMVRCmsnYQXbHZd2dUeg0Jz+yO1t9iPFpFtz+g0TFLbMKO6RPm+zJBsQnlm
t4vX20KF4wifKzhp+Qi9mbd8ArCoyOB+UFzzgqjkc5O/ChMBWE4hZCJVA7lN0bIY
sTAxKr+9pviI3ibFgI83I98PO+l/97fI1LqY+sHWmtRVw9Ol6E0SBt2lQCZ+N+em
+qx3bDkUYjnN8FEBwBLjCtFR4gqgRy6DH2vFloYZO79PtakT6q58zw+3Zyn8D/Oa
kg3jjGVUaB5FD2JO62IyDWsxCPdTasPTheRKfMQ0+QBvbMVJMNTbyXyk3vNVRm6G
7fR/vQ1BsEGtNMo/vCcLUvUl0lvoMq2qX4ZW37frNv/vzKPw01fxLuMX2Ek1gclg
ubutJE7Ud412yW3dwnyjsL/KKwiO/bfrNlOFVg4RUvg2d3qzq7IIP7b0+ONL3akk
XC36pCksFno5vQwxv0kRXcSAVF8oBh6MNW+/bOD9uXkOh0BkVjyVC7M1CKW0skv1
oPZySZ81jvgm1NvoSBfnz4H1KUuQqo85JJo9dnQn8y3j6rgkIXKWxWTaMZo9EBY2
bioMno+nw+Gxt1N9jYqG7ZHecmhFSYlV/mEFQNINCrxZmoCkDTcvhWNwMYcM2mi6
0mCJx8hgmTM8j2eHEfDPFjqDDpytyMGOhSb5EdIiEYg=
`protect END_PROTECTED
