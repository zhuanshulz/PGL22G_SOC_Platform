`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NX4Ns56ea/h6lbXpC4W9vvfId9CjBjK7HM8bAyBK95WwInbQ9dapmoQOBn9tm0xK
EClrDNlCgiQoSSv2RvuZhqVy8htZz1gRsMIqPlUnXG+SRHa9gfenmp5syIPUF4aK
iNfQ6qOm69jDJzwNl/TgDIwNILMZNBeQMl8X8DxTQf/sfxJOh+nTDkqD5Aeszo7X
FJEbmLoqsqp8VOwDLI0LOi1wAzIZhbbu+izKJWKUmhjGwNXjMrYZhAWc0q3ej+KJ
RXFaZpip8PP0iOrEHJemm+/8GE8saNgD/hkSe6q0ePFAYRw4689hBBcyNsqbXxfZ
tF/wHzW38/IvZ15GS3RlN5PE9bqiwFoiYFdmnDqYptzFA/IYtVqqB0PT+UHjGUFL
HUabZQTPA+54bOR8RFlTIABsGZJXnJeBNKgLLAVD6OBIbEVTpbc9t2aoNgUatvoI
DSgOPC9bEMJ0fvZuOxFKlnv51IwX7TcvC08E2BkxlZqGSIaocez//63NKaoo/mF+
l7VYHSWCO+zDUh3ZeagheHW+ctB0+jGqjU6iKrBTplx0sdArePXxovWA4GZA/c99
sfAu0bFE1kx1gPH6at/mGWw2wOdOWob+bdR8E8TsmItgd9Y0LDwhytzFH8xpUzYK
gVx4PF+rGCwL0YdhdpUGJDQSj9E7FZkFoWCJZ48yp9Z3dWZ6tddkn/YfC46ZEeIg
3Ks9gBaZOc+iytVXVs7twUMs/OWg4M7403gx1Rh2Jr5HftJMy+PioyNyU8fNMFGj
/hycm607uT3qCdPtxzXqI4yDpC5nwIbGRmigeuG0m9C/JiXRv7r4SPjCZjsu6jtR
4oubKsmJ6+wK4YEmmBO6hNOXaWK4ewvVAeXpcadZCrlwTOEoihRcDgPMy9oAaJm3
xfrZFsqrTp235Y8oveN2ih/uqE6M+2/bTIy0VkLx7ARq9jhQkpId2hDd9CqKqsxF
V98TFghKegHV3RHfud6yLPyZ79F9PnpqhicmcJZWaZuJC6Ny8oBwbn3C1+lRARG/
RCQn7SrSWfGPEMmNXbi3FDdbPuIyoTyeZSLJsBQAM+9ddOBdfqmXlT3d6SBjB2Cw
Lp5hGnUkqGxg+gz3GIA6YGvyFIayYC5vmOYv8/qrv6AUNaV1fFxc8fYoQZW3qsvV
nwgi6o6Owc80Cc1VfKAdcTPqkfE/IJcy/tjZkGAqDMwNq2n8qgLwk8Wz/uvz71Lh
dHqaJUTsSyWNa6nUdOGEXRG+kSASNnnI01vFrYH7Wc8IbIvQ0KD63svMTH0oTV51
9zdje6dL1s6hAGtMJUEyeGmnTYJf8GiDiqebuGdIrNvCn6Afva0uxsUP9eL92xyD
`protect END_PROTECTED
