`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tVeJ7BrN8vsIg0ZsONx7JNA96y3x+to7nhFjPPVUpgKHLw+KyzHJIbwxeaoR5MY9
ThaY5wL05fmyStSN/m7xMhm2TKNSbbQ2BmwNbraQXq5JnMDDOKEEk44hmBf6R9px
/dQo52+jnv2ZKPvEYngkDuhon7v0qSJt5LmSbvrQOs7p8OEpMXkSip8ps8hE8xzb
r7mNS5JCyRviTTb8cbZ2ZOAOg/Jw2oeOUsUNnZahfQ3kcrifzxQAiNQ46U4SWWmB
3gA4Ko04nG5TxfRRBx2aaQ9aH5HtAZNuCohWtT+pQ+H9Y1GhN9xbV5h/25HA8Baj
LoTsrA55v+q1I9TFoo6niKt2yGL9vUHcVQeoUxjfGv1Wi5FAgYpowzpnBobbVVZ2
hx3jd8ypyCCibk4latg8PJov1M1Dmg2+mf7krtCKHHDWWvY52uojxWkHdyTH24LR
AedzMdEKmWdYCxcUgLoCtU6/WnwiimbucwIHnToPC4/ZLD3h9KKYBdfkQb7MIUNk
GWJ5Xf8HbrprF5aFtYeKO12Kff9SmcK10vcJBgDvcgqpx3iyG9KDWQGkx1PYV3TT
k3yZEzWQSAu299CIrUxdcSg/xMZic9LXNYkrJD+IGp+152DGvWCtK3Emmy8aXifH
MTdfSV4e4NGGxQnOqnTebXE8PAFcK5wH5NfryEaLz9vn+4lIA+0RFx+/WmuAYJbj
ZTfHqhvNhWQo//a3M6QaNsFunqjalmtg6y4yWdLM85OUXm+qISL5+Pn9rji00zgw
`protect END_PROTECTED
