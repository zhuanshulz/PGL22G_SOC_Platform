`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2X4Z5V0oedDCnjztshLmpsarqooJK/QmX4XMc/M5OjaKSxP9MG949Ub+cMtFvm1Z
TuwZIB3mAC5iQr6Xwy30P7Q07ZfJYB67wnSue0vcw6PqERrmyFAjKGDI1slxitFT
P5gHxSRu65m9EE+ZtE1dti4h7X1Ra0VBdOKboca/lkLC4JSU/zwAzluIMh6R2dgq
gq5sxR2v8Er6aF9cITsiJ8h5fdki2a6Z32RbAAkYzkEd9T49pG3P0tnXykLTBPX/
UN8Da13wjVcz6cRQATHSGfHtMfD3b/lPX3FllqYYjfpJsOzncuKnv8CUcNZ+MBPA
87TJDg4d+JyPmg4C+CrQDj1yOa7CPocNOIxxvrKGA+MIswLpMNJEfosK61liCgHv
rZcJGGC1QDcWO+mzreP4nkoQmV612LB5mkxuDUMVENm7PbIFEQiDtYGKxVylt/BQ
heKZRPONCHUQJ3Iqlbp1MVCXF3L8RyRfvJ1l4FpzQHOsA4JWLzVub+vSwGEzkGs+
n0raCtTK0fZumHcqVyhX/dzc94Cn9PjCRAN8r6X0yK7ihnuvyN6n4WOjM7TF5k7P
YvfsLZZZoCDZqvo9yvouj8j2ddb+SIlFWtQzrexXtJ2c3EQkXY2NmOhzWbh3NKhp
qGPTHBP0KFsALfqCLxWm+vDVUgtKcy0F/e/oXct3uUmq0b36Y/lm2kI6XE7KURxk
bnwno5SjZGa9mfLrIMIW6Q==
`protect END_PROTECTED
