`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UnYUS2WiUpPEiVmdaRiibpt/vUoFrpcdarPc8AFM/muLjBZXSo4B+jOk0alwbaVy
ND5M82Pqrmt/3m5a2zIx3MKFlHFPPre3UR1XOFTMVNYsc1aVPX6WgR8byIc5TV9S
HVc8I9Z5q0U7z6l+pni1kLWvA7q9KHFkLa/htkD7+shx63gkG69HGmV4ZbXAY0f2
G9T5/ITh2+8jfBTn/tnLgejx0CoD72787B3sJlqphqpGIGsNFMGiUIC9l7f5CVD7
qvFlMoWMB+ms62l4CwK4CG//aNrLJ9iGrnl9+zhycaAi1uHnEh1XZC6ukogp/F3y
grN92KoizUTg3LxB/ndd5k9KHJ7RPbGyp16CqDcoKy0c/+a0OBXVUxqdmSD6yKSi
4CfGYjr9/t5ntt9sqnNo1ehv9wx/e01zbqOpksl2PiNGjZh+NexLttr72VhzAB3+
TS3M+hXCdInmHa2yE9LMY4C/V44eV+pyqguwmehuWDyDRA/fI1fE7xdqpbIR600/
tvRUu+5VySP3SLp/GoBScBQmGfcxhMUysSQJLlTZSFiN39BjkVRL7/wtzzJyp6Lj
P7s+ocGdG85GMw+uzljnHg==
`protect END_PROTECTED
