`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
11IRw2+bIFmuXyzO9Zp7YQ0PfefJd+NtZ/KhBUqb+F2M6uVhDXAJSrp3t13/SScT
jHc3JJRl3NIGXIyJv1tYBa8RcGzA1aQj1OG7E0NsIEM6Ok6LUjyBWUUJ7Zl5h3en
UVOkcxlbXQoIAnwC7mEGBgea3JI/yolq6ypNa4/Y2cKxX9aBpWzxad82xxDnZq/3
uePZKPcMsYk7jphNWCl6zqaTaQmKbcV1bNSxE6e4gb1fHTqFM0ZEnlM1lvi5tKpS
E7EiWfi7Nwngtf+GRNBuEXsauLEtU1CkKa1hlbD+gxuG+gGZ/b+Fet8YCPNzaOle
SW/Fy+8xqGPesZSa1XIW1lFSZaIs/KB3N92bdKs1PqSaJ3cVg4v/pu3BejVv8fBX
G5YqwB5zm1aN7EWejDKRgBqILrhlP1FJfkscTHw5jru3UGU+w6ALgUkUlSOV+5w3
UCI+xWTN2L5VWgVfyOPeKukWdOqDEM0+gMutFcEGIlZaR2EVZhQvoYSyWx4GJP8Z
AH8IRauZsERKps0bZOSgFgDko6EAQ97kW0SwfhdMzQITs1aLoJhW+6vGZjeaqjoE
x7+ScOimwH5MVaLydHbqepZ1bbcs7AYz42SnHsAiucXwrByMZL40uLadqBLMC1zX
2oEtSxUoJ4Fx3sZATMJenesgnEYQgRenNcoRAGDWydAKCnT/1Tkdf5PJn5RDX7Ef
/7gKBIzh1jvRdcXIX9Eu2w==
`protect END_PROTECTED
