`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aUf4zafrSvF8yWyXubq0Eubls3n3E1Z9FtY9rf2QCSTQKmAi1VodOlqhGcB/iufp
BnkDKOJ9ke+UczROyHIn/VYpd6Wy25gxN8588gn5zXnqPfGy4GSyxx17x12u0KoS
3GftO/kga0O3zKWQy0wiyg5sX/2uMxKMinExyzWR+nSrJkf7orT5T0LnlFG1/edY
ygeCX1/qolPG9yPbHquJe302Y7XnpY5dC66GcIgNrZHQ8JRvWloanjgsUja5VnSb
rnvJfYJDBe//OB2fKWUvWlRc7b9Ur4N/03ETAbohFXL7U9Yp0jpt9t7QwWpyCW2L
bRLNdy3sINj83AuhKxha/AGVqJHLBZ/O9Mo+XtZM05WhJx4Wv5nDRAz6ikDXnsgd
0ggYxp83bC3VVGDVcdergRyd4CCBtx9kYRNOqQVqO6IxOUPiHVtgqjm9/igjK2W3
TFhpT9zKdVzISc8GHEQw+cBYzPobn1R+XLmOxPwu5z4r6AS9IOcDytrgp0dk+tUq
WmKnA5Z8GgKVT3M2si1gdIvTglQUzq0D8MzUOFId3tNq/GZa+S231k9Zdr+94XnT
MKkS6IuCqgPz+2uddBwDsiGqZSCHA1asx+YWGbU9XIMrSaAUYGSXF6H6Dy/LCL6C
zR7M+EtoZj33VJBiuFwEYGUbiHYAO38nkVtXId1w7uz2qFVxL3hCgp5WDIXT33L1
8clvwNn3BjUOmRY/CDziqtN7qG1zmAt5KRswnntcZBoXkM77Wsp/eCIdf6oxXGqP
nzhp/ow0C5+Y4WOwEX4aWvAvbtsNj66o0ZwcGVmRMkqohwLgCT/9dvoOlK68iMXD
5erVoCXIFCjck7t0lspWb3g0WEaP1OSwyZBmfDQdKjIASv3+yf8ZUO+5eL4I/OMl
sOInQAb1zmRWcenCpGM172B4KlrRCajYofI7AZWsY0pCFP+F3E12AfVf5g2VKILp
rwoCyak0CFG8jDN8+VolNxj0pBqPgZS+7hErN8TijvjvTkqwNlPz7D+QCuAO4FOt
ioG9RDdBxefHWCAA8EoO8yhS2k84VLCfzO0ctDJzZitdT/vYAcd3L5HI4yrG5ml8
6V7mfRIyLN0tZc8oFF12ZbDxzYLex5PRvRVwk+92qjMNK4uiOYK+1Pp7OgQsf4RA
bzmirkCwunx/SzsaZBFWYxbfKKkw6AdjpAsUzZYj0UyCV9ftIk/2WjSjZiNuNodT
qBWC453v6aYODVqReCp0H0esLQDaDnzqBTMi9BwiXY3YVp9eS37xbxogNK8TwS1C
wJzmGsmFV1rxDIZVl96MX8mZ2cMz5yIqZHmxRd2jdAGpOi+nKo0i7GD8SmPJyJ+V
tRj2xHNoyN3ZnjbAsKuJeQ==
`protect END_PROTECTED
