`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2DCJoG6W7cnnP1aEukaSKqTwXkg+aMxpVb9Ff2p0wXFWnL2VY0x+k4kr4FrD0RRW
u5mZOCzcOuEIOPSEWO2TiaDPgqNgNFKNTZaiywyU5wIYdfd+jzHkWhcZx6LfzInM
5TDQQoxyOGgDAoxt0VNyflHTQy1a+N6l9/HwUPxAbYKb+6s7IgrZoSp8Oq+SBWK5
kJ2rgJRGIJizMcOE/VMs1SQ/pHNge1W9Rq/6aPSPELxTlzSsK/goGyx3w6KAfwMA
A/XnakTU7Co2k6rzml8GvPbcn95KvuVR56ATojaEBF90fMdDEAm2Guavf5dBHrwd
Lv3QM1c535j6MHm0H43+wAswbW5KBR8nrEpeuby+EdwIHdwaYwEKNo6xStPRS3Tv
8Ld+/GMiHbpUP2QGmuzx98fEriCUvfYvVh+pRzNtl4SezGhYDRKlcJODjatuXSw2
1XS+KZrE/D/B0ILemvVVZPiIsSSyETlbIO3NZ95/ovMkfu3ktxIE2s3Rl66Fs0+f
pgOtsnjiMl4js//9bFAsvHrA58v4SP/e1ucYboSq7Lb6fOwQqd7fx2lDbk7WgsNf
nFmocFMTITZC7ELdXMxziSMxsgRpNcndF4c640cLHc3pcAzRGIjqfuOCUgVjSVF0
NAXQpgew3yyQXP5uCPbqUAbLy3Swm69LVNkbv1co+ypbuuovYpoYVYUIJLtdDTZS
`protect END_PROTECTED
