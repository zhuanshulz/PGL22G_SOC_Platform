`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q4TVeJ5g8pPAcuFhnbsBc2pdlwrNnL/PdXvU/VNc/4AEbiD19UeL23b1bY8nKRdS
YemZmthbOtTRGci5+fYX7N/5DeEiE3lG3tQouSkiLeTe8vHoC20Vj8FfG9arehTI
DrrQoXgoj1KYrR0sh8PistdpjB4J4LtIB7mZ8UqwkT6Lbpa99xEsfLTsZjYNX96Q
6PWg59Ss0LlaD2NPFbok2dtU4e01fxAAP5SOYxDRTP4mNk2tSSLtRsFO+khcXdv/
sMDzfTJxDEqyTXlhZSlML4iaiJGF4OBdkSdp0W7SUF2XvAiuAFOzc7AqjKHoNGJr
ltATofzoXtqTs3XZnPBc4r4loFgzVtYRRpL18iL21ydSDPF62MwfMxaytk7Xiheq
r5O9MB0/kVpeONpubt5eY+69hIMBQ6U2uwXoD51DZol2Y9IgTG3kPwjgf8bcTGko
aAYKzLD0CdeiYDyJ1x+7lLrAKt5dX+zCRdBOqV0q0PmxXCfTimIczB83Vd3T/YML
ePEo97UO50u7MAiuKVfDvZNgv/uwgtoKhYMilEnwG/8pGA4xILlHQcMFqe0kWqMs
yTvXnlehczXI4bv6iFipHTC7FQKq/yn7i0fitvjrqwM19E0FF6WsE6+YwmsKCxyZ
h9migUFUraoZxmUWObrh1v0atD9lp76m+M2WFK5dTPWlv6JTUE3F5ubCpJvuzkCv
ExiC1pL9qQUsnqFWPpAU9Fa/s4dbI2wOyv0OIe7E9263stc9CCx4anVEWyWp/TjL
LP9JMh7tue16UFZH56pQ2qj5rFmDAqjG2I9eU9LP4uFozqTOxoUxyAgq3PKKvI+S
4b2s1w9uWF0Ep1ghqg3outS7clmIoyurYnrSY0bSvIhaiW3XNECB7PGPhENsoGtw
WKnZg2b2sPrjy9+ZCFquPtlyPBML8qznCt1c8sTaLvc=
`protect END_PROTECTED
