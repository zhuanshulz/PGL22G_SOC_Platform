`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+64L7MZypgWX9zw2Y1uiZHIMbLqq2dX3jfzTI3fPahIn6g1lBmL1EqWpaSGzPkr/
c2GKZ+huLxhsoKifsyXMdWcGRhh2UlxqozwHZclFK5ZEDeGg6UvI0hw9Ab4FtBI4
nDeHZgVMvnSs9pkxHETYAEB3eQi91imD5qveS7hWFA1EZ3fGaCNRn5JZlzQCPQg3
i4WF1hsEz/keG+1KWRbDQh8/U550Dlv/upqKCl1SfKp7CJy13Ph+N2nLss0O5xYV
PHYbuKMiHWErPGPFg1gmTo9xWBq2VZ2kn/3GOQ0fPQ56Twc5WA+C+f3N+cXuECSd
hRprgCBFo4OSIXy9pkvOVnbRe3RWhuCHAuqlW0JWMpQNUyrQk1SfrQ1oFdS/nIUx
tGCS8afXh2LAai4KKlvSLPwBIVqcgmJC/NJtNHjB0qhqVVbIn0vZnT8YwrcFBQmb
avoCnj7cuNCRugfbVqUWDF6LbwpS6/W5sPiioROpfEtvrqU61WGmeLUHNxD3DE3Z
kde/pqn8gmx++FJ/Pi3CFtE7lsDUzJE7JQtAz8LokYTQ3iuoRUxfsmJjlNUDZeyP
VblOnkmGGQqvvIumcvG8GHejKtCYytWthR1GAYv0ke7qBVPK42Q9VmTADFs5N1Sh
yTOCTtKG9tilinigh/oOconmpnO7I95/wTjgw/4JAuTfqwt3Unq+n3dBVHkr//4k
PshJogFKpNCeXaSXrLgzXg==
`protect END_PROTECTED
