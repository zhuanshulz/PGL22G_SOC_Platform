`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RrbOnQululRcpNV6ef4TEYwhqkQEk7VrwiWo1DliGDMtM1AQKTqMl+XSPoJcoiEV
rxShMWzuDsM9jUls49WIREHQ9b8DId5UbBCb9zKfRCdQ1xdaeN2FvQMhw2f2nOJw
ooheAYEdY/yzUns/d5EoOpbkoh47K5FOaUU+AM5otSjARLv38fT7nCfr19CoePer
DmObyKvB9fXEhGxAGVehjArcbq1Ctz+fwICLsSXcVq9X1QJWLNBHO6t/92uvNk09
i4C5ap/6WQkwS6Mxn391O9dl8pff1cP1yLnLGJaxU+LKDCAym4yL4NbvC50D3JyQ
ICv9i7SNBSOH3rwRJPUembdKL3raCVh7P3PFqfQBeWX2SY1fAM7k4sLhkm2b6hGC
MYNS4meIRIOxkCBKj041lTqHNP/VSIBk3s+SFe7J+R4UktTMvSqSD+pyh2KW74/S
EQt8DUsJweLc2je4BPdc+uyg2rr3fVI7NSGzKCz1DqHqg/YsWEqNxV+JkTKNvWMq
/dZGjCNs3Nrk6/rmRbJvVK1xztso76AmmndtuTfzwQmDYVsaDPEY/npq0b/5njcr
8krwVAkq3DHr5lgA7vzBErIlLeSX/P0UnU5YsiPeTMfT4x4iXO1Ic3fAYGf2vzsj
j8BiXcVO5LO8bKtQ+ljYgQ4AJVI/0P92O+bHZfOIksDJKEeTktaMXiEFMSfZHUzA
jYaGj51AgE1xWzMJdLdHmnDwnpRcoLkEcNlQw9ZgI5/lYmXDDSgtSknrIj/HGgVD
gBMLIX37xRHnSJbNwQwzmvR1fI0WQcNYfDGpsR/8UPmYzkIXWNgPRI4icQHR/r6T
FfoFeHuIF4/SF3r/SC+B9eihBPBAxY0OijrnOByNWXl+zh8Gy8id5atEC4pCzcR0
NmGVg3Kqj7j0L2RP/B2bJc42B1eYLwUQqyxvC7WtjF8c5hCTG5pkQ8D32jJ2hoFq
HjMRZEtIZ0iLykmHRIoRSo6OW/J5tQxDwtTD/CIQN5dGx7LKsgY14tkycO2K/AWK
trJXYvFhktpDgwJawxOMvI7TJUUPtOLF2QsIZ3lOvAEkA9IrIjDcp0LkeaMwJgDj
N74YYzJXwZbkPPMtP69dk+BjGWaHS1yBnPtAeI+aqxczdmZQwCTZsw4u4vwPtVOV
w+WOS2QHLzTls18M/8FVTANeIH8fOutU1xcYyJJ3L/LEMt/iUMxXQr3khF68lb7x
8KrK8Wn26zKuPmV9hB/OXy9Ly2vlTxeff3KVYxFc2yi64upPKs3NNb0B0vjcBZwN
ZZhiQhEmg583O8T6udFRq50yaCJy+ChVHtH7KiyjDTscy3HtDvfw8ZKWbIrWp9BL
AhCiqiPk02pW4DdNWqwMnQWkdJy40DsvKw68+RucRgyWVC1BqqLkE6K8oKadQi1s
neOEQ3qaDGth8SnvdLzW7FlhBGr+8OWP6OwAEGNqU+6Ddx+Xxu0TouYFPgI6S+wZ
yPQhnEQ09YwhIn6xcs+UU8L8g+DzhmSkETU4qEq4JFcwBiIyEaUvkVzDz5lnObZD
ra2/XPsn/xWnla2byQHihK9pgPZgD8id8f9rA4knvb1n5YKPHZCTZShebi8wetGp
nOqR4rXCFdoZov4MAWqWR1HKeESegvUBUoiilDOmapw08Cl86PYZfFki1/paHlg+
Q7mt84oDETwB3iTICjQkctcZ1DUMEA+HyRrNgn9dKI6wMYv/nVCCPkZzKTW8Oj82
UM07zQXXKapttpJ1x+6nMAWKCDWUlJS0r4R6w1ogbQBqfus9u4u190wTDTs08syZ
v57rkUaQZCFD26UTOyqAtTD+vnYfQvqblGCgN+EL/CN2bEPI5SjaybPkhpEU96X6
YAQprYnliK6PwNg6HWf6YO8isGwoKIggFoN5G1YRUlPje1gS0V8e3HbmUEaLRWL1
cDjf7zkM3MisnmFcPjceIjaH7YVJRZCm6cBSO/IaMXccztHBvHb8bdAPD0qnZsof
uwIpD5vFHiIlb7slRj8F+mKev4yBiENN8IwtmxGOkXDo4c79jKA3szVGx8SLtXpt
I1NtvJ128dJFw8cG/AEAqoNTCEy+V7B0YasfHP76jVuVUaggYATbDUgH55/+zRqk
9OwXQcypWuxxrEZA/d0FU+r9q7MykZoLbIQh33GLQX780Xtna/BU9kkY/NcG6m9H
g4rMhEjKzSsowQjH6e9NSyA+zwa2Pkq1/Vr9gyjmxNg6HW9gw0Xbpj9CwO8LaFbj
VPCFn5pKMaQlaMf/mdoB+4Ia33etDtQkRwbT3KZEWTizLA1IcNRYLjdi7gPmfMCN
5azs3D3JPLyO4uthfq8Ks9qKHL7F3nvsB54EyaDqdblpHQATdYl5ZoGGZld1tmkQ
vPnsUXCunpgeDdecBqnOKadCD46IFmhd7V2+MNCI/6asWuQaKrz/YWoMzJhW6hci
fpeTEJC6lrNZCUw7HmU/k6TZGjvdOs5H4OOqniqGWFpciWRSQPfMqUPdsaLiZzn3
QfQQXZNVI5zdoS1FcxFK6Y4ZqxWXixgYNqngUcOn4tixu2xb63us14UY+gpFTq/C
BXjFmnGt40X1I6G0f37pk4TrbL8bQ9IygMZ//5zze2XiCXvcY84QnUlno4JwuRj3
eJsR9k6zZ5gXMNKpHfyVchH4UtCkz1nl3FUfhOYOSs6mkk24IK8SjfjQkwA1+1rA
IYhE7y6k+UTlLr1YfI4qSsyTzwBnx+g5jCnCGMTk/SXbyr6GZKCc3TET/cs9PEwU
13KkV+vKpQ6xGeLg0bfaQWq1Nj3N5wFpMZb6U4vO1OA=
`protect END_PROTECTED
