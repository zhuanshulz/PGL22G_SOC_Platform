`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3cKmz6U1dAyR4hZ8wPWRELKg1rhvCTnTguQrcOgAxA7Wz9igQEOxpMq+W0KoqnCa
JOLWWtsWES6R57WOgucTzJtAcwgOeyFj4QKkECVaiqq/lodnvbT5GT10QHcmZRoN
EFvb/9HLFUK/qW4BrmTPb4DlddbQ2WC0hHnM9nMrB3dppEU8TucBXb7d0g7I/XNu
GwLJwTcj0/koTpSrgx2PT/0oB4Rfmeet2seknw1lm0x6fTrROy2LQ0MQCFh83Aby
pccJRVm9jtiVIsPtqmMsVHg2SsEcx2DTcIHet2iFjvaJpPW/bdONPDSBjjFyOfnE
bfHUGR+2ZZ9d9dLhEz+oKLuhyqNAQn68ddTOtp4PYdkYCMCEcaBSQCSaXmqK4nFe
jmkp+Fb4XLA+AJkTlWDgyYqIyOSP3kaXsI1XiWMSf/RroZKBSOJCJwtuBLaTCuHY
13zVl36Ma2sgDMsmUCdFkdnq5AzfAefYa7PdIx5g8W8=
`protect END_PROTECTED
