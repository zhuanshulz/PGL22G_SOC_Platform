`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HG6gg1/KBI4y7Gr2rKh3xP1F+FxmAEZvDTEMgVC7O2HV1XgCytU43V+heE6g659G
C5lBr2lK+df7dhZMIOYiZv0/YNDjyLycxQDU41uBjaQ4sqIZpI6RIQYWDJftnHsz
Q/w5SX+CMw2wQAEjitpl3/lB3lv5JPfesztF9nxT1uQoe8rdn5XGXc2YaXPtDihG
J7NqatSXMXJvc1s0AARuLhGF0tZLWODn9B42D0k8GBcBA2Md2ltOJuTcACnEp3+U
cCjbElIPWBzFjD/XD+YyPMLP3aDGQEUh/ygOAU6EkLNlmxs9oBqeCzUqaUIZg7Cw
pQgaws0n3/xKRymF5aARlYroPYBPUSSspw6leDWDgMmNfpgpKLKsiHLxDClPb/i/
byxA1Qmwy2fGqmFBDpkO4RYLlPWIYbIB7FcmcH461xu8T3EPp6W2H3ER8r49xr7h
dDXG7Mv+Z7Sq/iUSfAsBCFadzHB4q0A9Kvh42M+1pyx8loN/eNGCDMrxH8F0vjfR
Wh4/+wDO++z/0KG/z6J1ITnfzu83MMe13C+7LwR+UcRIbZzm5vRRCHaTTfWVJGaO
fUf35qToMXDoUX/bF8o/htCk0/iMfEp0NauvRIj9BA5WvJyZoLCZimJ9Ze8zcnr1
pBKP6npQc6WcYypgHkGcfJ4Dx2Nk779N69NtbxS9PaVvH+l4yg25V5irntYNbOKV
lAzWVvhF/yyz+BuPsAp7weJsSIDaNmPKLNwzlTq3EkwLWOWphWVcRuNWVoE2KMSc
wII5nWSZ+MKJGir4NQRaDyLAXtn/mF2bcuXZVoBJAyVhT1bpHMjJDKK/v+QBrsPC
ve6v/GBsncy0O65wxpoSQtwsJPPK3BapyV6XtcVvEo3qrSZUjdtDyI2h0T8//X/Z
DN5tozXVl8WdNs7PeNJ4KksBf4ruFxGRzzz8OvdI9ESOMi6itqHicrnVThHmzIIo
aXQ9IoIeW5wnB8K1Z0UthTgPGCxNVPScLSKAkcNR4STWU/6VJKuF3NLQLWuYqYWR
ZYoE5bYJiI3pkoc/lhMzI31qsU1mpWrF8RWRs7gx1EK4/mxMGmy5zE55OeMeFLmh
npyDWSLkphieQ1ccZHZlH0ChblDRHYRFC9uAl0KRFzcOgNgp22AAVTGjsgcVD1M0
6lk1l0j/M/DhHW0JfYpYXky09JDjgY8+NBkWJSkRw4cI3mgUFs4t8A3Y/5iEhjhW
3BWwRL+o/FM/ItHG7QVSaSlrliQXcsVCd5n4pr1oR74=
`protect END_PROTECTED
