`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P2mqZrRI2o7hCmT8XodJUKq7JRNwkBS42o2Q2Rj0L/otKe5RQSzJKKs1a0eMKzF+
CzVcOMMVZpzNeexoRMjfCKd53QD2CNZ/unctcUB6M3J0NWDc6D1uMbO6V3oQvGRX
Jg5eereK5jLQHgkkjr9K9B5IvE4uvF5Gdz/NTR8avbLH2my9fjgtSopyV0qhy/7g
P/Ri8lkzv343GFqs+KkbMzIsTsWpSF+FQ/pVpYM5qnfho5OqHw8p92XvWw0DhhIB
5B4Tyb5zSKOHeUL1tLMcXFXe7Sp9NGFNMzfQh+YvoVp+TqX1klFr9VdI9Oj1B9aI
QVP+PsAu0U/KlMkOY1VGVLO6uNmhaMA59qgv0/xid9rXJgDu0yxh5xtQOc/o+FRO
2eLK7/hTh41hm75/IW7HSm/qLk35VrUcwF986flhuOtRciwfydzWyaCTGLEliMeg
u+W5Bj3Ru0TuKlbg7F6k+1kWhiCELQYTF0ndsuJ0js1ogYR2EXRFSGmJud+oM9zb
ZlJtLhCv5nDy5M4zS6eJom2YaBvKlKH9mzZVjsD/LWwCLeb+IhIWNBv83Vm2x1Gi
LpXQrRY+j7ZKZpU58B5VZeHbQmhyTy4gzamLuZLIZ02ep99llZx7ZuzBvmkiaEUs
X4xYKW4PQKAzImBOQhQq9g+lq53BaNGM4yySfJIt+iTSIftkaDQWKMNcPaub5FoI
ohV350aUkVjoav07Ku53XfMO4Sl/Ovdr/2UyAJbwD1QzJ37qDMfjQPQSXbPgE87s
gpLkBWNmPw+Yk+5Wugb0mwIcEwnl9QQ4fOOs01aCP73TxjdipLtBB2Yqjy3kD7dn
zGSeFTZQcfP6nqP4dFuLDWTWaTNis8g6b9FidSA/QJL8hb6+LI4lMZVG50nNwrir
AQTPfLpENFTwuGW7Hf0WGxPpCfNhYJm6qRcXMRCVjitlL/fCHcp61xxnzMe8OeVr
21qXxYGFhqQuVtVcI8dBt1CXaHIgvQcbTOq9y/ti5mfCtf+mQjlSUGkfsp728YSX
yPqDiYP+U2N1bfYyUw0FN0gkWD7Yxz3+4QIrEZt9bPxBOlfWMEHkbj66N5PlpnMk
6BAWdfj4DSor/o/OamUvfTnBjaCzyhh8/ZuxSy2IcchisIozKURO/fnA/SvIq/jS
1oNb9ZbfNNFCJxVFU7j0tl2BHxAGMBix6BxNkHoIvEo6JN0y4Ul9p9B86WhMw7GD
e1wbYoHx3hDAT5UdTobafqrPdp8XfXcw/MgqmWtUJYYOMv05IfuIuyvNHyH3zcf7
OhBiR3Ce12URyfdJ8jLMt6J4phEQ7817o8wQAR1X+8Oxkzbe9RPrR8VAmXEA7IWi
pj45hz10jMThg/qgDUmXVtzvwn/UxKKjb0zVAoCvATOPsj63unR1/T2fq8GVHgDg
p7nmyocjfdLUjyQZ8XTUq/SHSjFA0ZUIIqIF9+GBN/4e6S8v664XfwKChSMFM3Yq
sUa1R1pA8q+hnIcjuC3zTPxQkC024w/prBvuhWz3Y1nxGYBzEps3mmtPUUtab6cw
COJzleGl6+lGqIfGfIuYVXDELIDXcfbfV6EJzxWjNcuMBDLHwZYx3RMG1sU0wVKF
euXLERmH+rqFO9PrEZGH242f+DadDGcxRQS9unjwpXdnfcFtC1Vqp4WkU4YGqos5
vNpq9JYgwAc1oFNaVW0+ljcDeQSlRp/1TPWPx1IGTvyXjeXkw/8SpmBktrzrGAuY
GBQC37FXno16nXKxdYIYZs7XnmY06FnsLcq2KNg6pOuXr9mOJ2/D5YImTKoyxH3l
oPquQJDK6cnRlTd3WCvMJwwyTNQCL2w9xsdWqf63DlvV+ZPqG1o9YvptG9XFWMVI
LlRp4oa1o1cv1nIrXGaCSjSguJCNYovr/3XyPHBhQGtZgIKDDEfxFmLK2xtlYlfV
cpit8zZuYrLoLT7+Xr7W8NjYXDTWuPjNhicPR7E+mKD8CZR4qsA0+VI884X1uirG
fGsgUqhMu0bXu9dGbIvsIBXGa0IOWUiYPPZJYaWmSL1E9q6Eb0Uik07o42vovAkB
ZCLKeEp0bUL5oWMkfEkHeM+fx1o7WuDnSY8EJTDvW8ZK5JSYpbfNuJXb7jUnrXaa
RMvOJFCEQd+4MUQqxKCcjZ+tX+6t2q1a1pKq4ecdSylvamoFqstV+ms0oJngkuoF
STwQttl22jlq1mQEk3P9a9OEef3yoUH1Wi6f/RBYr3p9x5f5jA/jBNjUs3q1XkEa
qaCrnwJng4OVirz5dqM6Z7T5vH5DTjzlWp6gJ8gLx1Zjr7ZmqSnJonChF1pL53mB
XI7PhXMuTphXBX5avkDMskYfQwFSmzHNS3QrCUIjqBOrCrI87+ycAJpqpLJ0Ere4
XLYZ1CCeIfEOEO8py8nHw/XBkYykdsRB5vKpQ8d18pd/W9gSJLugTn3D+sguGujc
3xzc/vylKBUoO3vejc8FtPsACDqgjL973wIMDuhDoEDW2c5/3DbXC5dLzxITeXwj
OScWq+r18SwM3Kktv3IGM4OKX1EjbxecxOagWv8GmkqYKo0FAvU6vPSovCZSNdMK
zaWQUkj6pWU0XuHuCW2LYCASztnSGP8g4mGZiVA6vAfuV58TVBU2Bkz7+RT6lMFz
jPr27/WTqC0HIHeKWxr5oLnn9gQej/Q3t4csmmohhIVmzI3eoJ+Xng4I5zWET0Ae
wEJ1vsgk08IRBF6YLKlBBCOVzROmudm6QpkHO2Cc9ip9UsYKVcFfved5jLjJ5BUV
1aaY6FjLjGsPTUO58iNezzEytzdNAP3C84OTootqB9tii87eVtrbCPZOftkPKsMU
AczTQ6ulLhBT9Nmq6lU0cvEnI0rElEoAVWpvwSiIrdw/P5PHXi3qXAqVTiTwXFzB
k63aa8YPstE5YpsDoTEAe34rJKy5ne4PKKzgLGRO7Hp15DJ3Ov777dlsc4aV1E5B
wlyPVD41luSamiKnCMT4AYhD2+B46aPjY9m1L/HLU2z2VaA/z2mwnDPVqTBgDNxO
nHjC8g2nxCxKSkMZPQsAsyV2zyoK0heerHhXFfVZMfHJI0U/50cFXQv06Kw2osso
KsmyQFcVk9TCQYO3dYWapR5k+mIy+rDficpka/rltyJk+GC427ozpsn9Q9AT69gr
DsfVXOzPNeXgnF+5cztCRTq4eumNYnM8noPEZ84uRv/lvvPRJF7YTcK9fdeeclUp
14MXBFEmhp3SIYLVL1wFMvWUiEABrbUylFInTAf8waPSk+k/LMHggOogWura+HMU
yRc7JZwYHUSePaK4EBZcSAScd2Yizq+bJeQ2GuOtkHmg60QKqAnK4APg+gklSDco
IF4/WRUh+JkYVWYECNgTuV58JmiQmO4gJDAK9RvjM4A0rCFqhJV+MtusJcCvDH+k
KK7zkKxUKj+LTXYmsgi5Ub4wm74tquYehHrN+AB0Zq4QUNFqdlNeqd4LGRiXIBCK
8K7b2PHW40XaRvkChD8NZLgzfJTJsDxQONhn52ztLKA9d2ZkYMph42EXWa+NjM14
xfFSL29NdpJMW1tDtqR28fkrqupWQd+s1DCrrQDIE91N0AA3gpvVu4Kbl3miUSfm
v3RRwCjzE5oUmoQrN+MOkYm6jmCAM5NkIpYWVe5Sxytlik9G+MxqVgzWTdiCKwJv
tdeJr5vG9XCiY6FUi0b5BCtfL0qUZAUQoj1ji/h3ybHRhf2G6TVaa/u/3onc9kj3
BNsV5kp68I6ZWC6BzQMrEBweAXnAC1Qc8URFpPEwOeZoEL3ME/CfvlyYvcubBDVD
eAfUQjshfjpcZQVPKeoysmX8UQd6fHIofqqhObBUUUNQmaWEpo6nXA59hu254kmv
h+JGLgUhYZRhkeT7f5ESvhFy9dJF5UDrhbbS8tVtpgZe4z9x5mdQ2eNkrDaUrrQB
7xTFLOIBaRJsHPBW8CzCMH1VDQGwmLwf97gfR9SOySzIZOIpYj/+clQ7BD0mfeYm
EPwWBJgicGIdDQty+erMyGGCDA6PA7/kvJI8vrqC5aF0X9mQn6hTIfgkCJtPMpx+
oVaYxwGCEfG0W2MKwMHAHx1Wyk3NMo0eJUus+wwckcg6narH33roG78Ri4l//PW5
sN9vWnVdUF6ZJY+XMCoykgtBK5hveiC81rZhOWWGf9riP+F3dlkGQxH79QHDIdz5
3+xn9WdCASX8H+28nJWUft/Q89V1ICwvMwUJne5VKUK6nmUbKKhI4xA2dvLh+zuq
EjPUMJHDGfYypJvcOGE8e3QIuJnz7pJoBHYMLu7aJ3hRJccs4qkvnE0DsyUM1/ab
O8vioslbAUeaT1Jk7GzTaWXrSNFpXd+ScqdQ61BfmoYfS85NdM7+hbS0Z5ycthXJ
DEkjBfA1gY+yRHG9sUoNb+sNCfdVIeQw+aO5/1MSqu2vq2dWGpjbFvleHuvva5yF
mg3V2cc00w3mRld0/u5iwrP2hIMWexidGEZxSQg1IutmytJuHlV6XkO+4utFvkwZ
YT3iT9lx3I2bYwhbWNuy9rCdatzoR7Sf8+FnX/2D+XLTjITo/i3IDrTJPg4sD14e
TA6+X4Ipluaa0a/5nEkpCmomhBsI6bjgKSAQYdxmilaeZ6VSJTY2cxTam6T3eBMO
wTJyLNe0b7yK27B/Iw0FD+8HpY18/aVqSb9+o6fmvEc0iO1d4j51vdprTl3R5mYn
9ZHDHliVo8VqSxYnDypkYcR6dcUhF0w0CJ2I2aQGirHDjF3X0JNID+PjHcSQSWwh
3O5LI0jtBoip8SdzAfaUItSeoESZ/3uiWDyOB7i0BqbHYOADJDhnnL0TRrLc5tQV
2ob9eKMWKExJOhWXq8yfGj+XxLNEINwmIF3Whj5QA1kPbo0Dv1pnhXyV2fPaIK3c
tWhBeY4UNdHeQEqSQtnljSARPx1QxBR+WWRppv3+P767mvlM/CcKqGQavWaQpfOy
14vzIq1bkrpd5AYsLBZiRqPTXjfttlE3aGOowDXVipxl662veOAbsg3F1ppuD+l7
wUHIHzM/l4DdkaZWKZ1dCB9xDL2OhLXwwZJO1neLDRhh3nWbfP9EdZkokAIsERb+
lJzfiuOrZ5Q1WZ1nqA4Wzeyo6mfqkjnhTr5szIteT0VpXB++nT0CmQKSRb3zI9+N
dDsvFB8K327Wgo+e4xYIlfbkX1+8B0X1F04cJdryUrISoep1fFcQEXn6Iuxw+diW
ySKv1YKh1ArokFvSgQOi3lHdPMVG13U+AaPsmN2lmyZ6S5XLuLqKXt+yj3X0jjuY
pf8Fg3WeY2qi2JtLGW6zg5ZDQDnBlIM+I8DBXr259hVw0UIkSzm4ruMCysGQUBOq
N38+303WUwyyBKt33i7mMccTmN/LMtCRpPHsyY6vu/La0Hhd1b2DG2NEbu6ous1G
Y5yv1qgtTSPu2uZvupGtFu3x6CnPHSJ0ASLTFT/UdPCUIhLi5z10XnHtmxtELcJ8
LrNKsSzyhxNUToYRUwQ/fRF0B/i380QPD+VoE3SBlZ6xNLFGlurKmbBiI10tlg8U
7aPbBIqEBgnM9GnwkAonHrAql4trhxiVGFP8gW0uGMN64O8L/tEoV2vY9lhrXbHy
K8fhQo8nCcZO4vZo+f4zQnV3Acw225IO9cns2+pzXjZsD5vN6ZWI3goQucz8d7dj
KUTuKqYtbuwgAg4XYBAJJjMYty0W7I4kHI+D4RLdSrbRhFSDaHLAey1JVF+rj8Pu
R2ojz/6hV1BWDQ974E1jIdspl0K4mqfHDYqCP4+ngeohvZHPo8gwD3/X4cv9DE+6
SWdi0tqBlnV0MZzpnYsry3sPiWTWYveTOBZYgVXgY501HiGMnksfnIoq1UgrNPHQ
61DOIbgHLSJ8AFYevERLmBjBml7uwLr3mGIoXQEGfB4cnYov6AnUjkr6lcsNutcM
5jumTiZsgN9nLFH/GON6tHsIz0erXXuECn4kWmfcDQ0Xu36qXl0liPKmooyPLQ8F
LhaaqwVU4ums3ScmF/3yRbeGB4qnbjHYE1QP/4/7h61KxYh0HbR0tCt0sh0qw7G5
7sXqbXheRIDSmJbf8IMRDgQu7bkHmvkd4yyPF282YMW9dS4+jUct9Hs5WZlHyHKt
Ur/YHU0A+LLVKRJAAhgVY/G1V+ZHjEIkJ1UL1O0XSB62Y1UsvZlUfYDADiwmWw5M
rXGZfBLXNaO39T4IDmv0J6fpF28f1CX7lqWELXVHbdDBoQp4v+3Ig8TSYwYFjQct
GFSl+yGofJ/DCqtGmfLedT0/EMWrI90dgXVD+MoGbzykFxnJralPwnU3S2ICEwd9
d8Dbd8YzCdr5Y+GYgt8w17Su4UdnsYWAyCBOn7nJUoncGsh1pzGRU4FOGW9nSCkh
cgKO9dc7sD9NYkUS/vAOjyxj6iZCmN64KK4AmjL2ve1b6wtQENrJABIWkGYpd5kq
lUIwVT1wVxiUnlpkjnACLSH/wzfa4xHMWHpAcppT0emHzxMX+JQntnmh1iqKNKal
2M5N3oKJZxWZtpy62OnWuKpgLvKARRcx1LwVDWB3LVw14zldB1xBOQ7CMz7PBbHP
Un29Qe3Xq1P+jQ1WRyyZUCRdAZqD8FlIq8P8DFpaVnZB7rClnmH/jLzWpcBCTHTn
goKbsKZJ1c/yAsvV+NEEfl3cr3a2gCyDIAXZ7DcTvgJFZnW2x1oG84TPW2mPlnVb
DYi850p2k6sFfg8/lWkn13YpGbfsIFi/j/3yB1uznOAMNlKXa+tw/FAlrxNQo9rY
Us9+XXH6Ln75MvP2Cyp3arIboi7NTyhEM4PevvsGgDGKnPHVsrcAkvSj8hG/kjf7
vyK8irVn+bDjK6avkgCl9QKrBBqP1NB+JeOcu05LwUtySo6WF/EzS6nvmcUC65/K
r6ovyRBPH850qr2t+bGqVAbtkX1C78+RBOmbEWoNhy5BkgWqEC1MdnnvoD7j1deb
s4ciHcGXK5t7mAB4UpxV61u3gcngNJaagqjMu1O4EBqvWkIsq1yivSbIE6F4rJbM
hMTbejv2Wb+0tTwdyWe9exuIAx4po3c1qslTAREL0CfCo/MRC3nwj4pTrf5aHJiv
kK3lzP06+RhVkvWEB+5E+SZkUhzSTaaZ3Ag2lGLkg2odLBMEvF4rczU519eUOGHI
lOaSO7di4TJyjht0v3Ih6jyz3sdPt1ZrVhBiz+BdWGEddy9aoYGs+7CBkSbNltH9
1xU1Nj7YUdU+lQCJBGzbQ5yRQQA3tJz8UGDT8iNfOkFeazbCKCoPsHnWsMT6VelY
FOL8EdnQPXmLxIIkPWDdqw3QonZJeVPh4uRY12+memINvVJt7ghvIqfxfaKCZWuq
0pvI8APl/5KSiI3lcrTEXVhfG99m0XITOUauCWrSTjyXSUvADAyLv7zSNqEGyWSZ
Vcm26Gec4VjgWWCb/k+rDyHnwNPp5OYDf9AzYCc4R0lFFjiK2Buy5DRry16UlGDk
USWEKWqqDF04pa9+HCYebA4NpDr0jAtBedWd0mZTTubEvZ7tFTUPFN45Ti5GuB8f
3tdAX+aqmUOnb9EEbq1x1+yKCiEywtZNJWEHnRY0piOaOA2P2OFFdfby2JjfgT8H
H65ikN9u9VqOuHAokQpS8vHqGIJbErIYqcgsG1FdO2fn815YSdzP33vdUAiz71wF
CHZjHS06m30ktJrmjDpm0r6k9LXx/OsRNyWBcHqGx/9xrIu2rAGoe/V+u6ZieUJv
JCNftWoyqaSgZU+12Gd49HP46xj7vhDnZ7ECgr1snFT2TzAqSfaK7EKDtlxgA5ev
gWWl5wMLywdHk+5ma8SYsZamLW0wv+TAVZuGNv7PV8DknaYHW7C92/DOuW/egkOr
XzF3CXNMDS5BE1fHebW98Wv5rpw4dDV9edNArMAPB7peTXiLInXddyiFisHll+xh
SQhP1izlgD/v44uu9uPdeTttNNVU+vKgYxy8oXunDK5erMX8Ak3dH0pvvlkeGyMg
zIiOOLLSVGZfyjGpmXwr2p/KB+sxKukaeId76CR2vxDpX+cuSTWTNP4B70M+nwG9
UIV0JMyrqr3AAV5cn3t+KafMbcUzZemoCb7HpNthM5JF0Q3f5qUV4qaKprmK2SP5
v8ZjGWFiXFqJqXYCka/3u0V+UQbyKLdqPeKmxowE2JlItQuUQcNCFqleX20BpZmU
HeSaHP0VGCVV5BUo9SvXLSJD8WU3v1JTf86E6c+PI8b390A2lEGP2lfWTUk1YSHX
TGJaS1rLasfzKGhKBpVZcF2wIvnrmmGmILEsgPp/3tbMnhUTPKU7fUlOeNmq/uB4
zWvzAHGFrXw21CEsEm2XurcX0Yv5lbW6VRuMOn3F6witeJeHZJzePnxfjotQw9dM
SIETHLtLnDkViHhnErIfR6uki0r74ArLXDAtdRcLs7/AZvYBMvuaOWWGnF35MObU
hNel/9vDlugcibb+3c4OLZAQ57QLGtoVy/wQUutTb7VjvNYkpaY/Q5KeYVwFnMCy
GxWRLq+fpf0RF2OWBbKMUbKeE4QTIYfJJYV4a70bz87+bwpPfa0VD55ki2qU9hZT
RhOW9vNaN/E5hdOMg4bbH08+MqSSqE4/knjxXLuLmD3qQ9l2IOS3xPpxUTQf9txT
swZ1V8svKtKUjp5OjIOJdVnUfTlpVH4aA8saALH3TeamXF+A5LzIJ826Mo+ZSTXy
J9wmUbQ1pXm2yt10WsJO4r7eRWhPTgts9B64aCRHRikU2/qumBSap/XRgooZPhKj
JbyegCMjfo4zp54xXrImWPsLd0JNDIsRGn/Ob0sbhzG3ijWtMaRQlth/AfUTLmVF
NWHmhea7QJ1F/9FQAnKgE1DGEZmTNj6ixWArDtIpsDLxXqmzx5Vis/5Dar2qkx++
Zq4cYI9U9Dp1wErEsP1yjGDqG6mfZdM6Nnosef86SCwdDIcDL+C307RxbDnS/rI+
xdev3L9G/pBCTBfHBe1B9Xs6MgIxmyT9Aov3M8TwV0j3bJ3LyxZ0Xi+LLX5LTYkf
64Dri2abVFF150Nlt3GbE5WAF6nfHFVUiN1XVSv7mhEMLGyce9eOi4hf5vNPlpfF
vgFIRBiVCjAGzkSUwC6cCZ0s37PlkMktDUosoqghHV7beWaBi/eNaADeNu6kX/Ha
IS80TTyPSBzdJr4L1bDujN9meugAWGT/Ne7wK8pA5eZvkPhWEpwS+0VYBI5QFacO
ByC51JA6PUdOgFk7bAIBVpPigYiDHpCbw6eBsO5rLJMCFHMho+SSxRdsLeODkorx
9YSq9J2JjL9GRhjbyYgJ0FHe5BXQ6mUuruvZcnZI1J7YAynHDxzn2PykBEz42CDc
7Rti1uH6oWRD2o0NhwjPAYQjLBcOrDoT+gBMJ0bKxmvsQifCM5sxuReu9DZUWaZo
vCuPHk4Ld1k4RXNyuqxnD11FNEn9VT3UZWc3U4kr0fIAFjBfa5ZFGSrTpj+OfyIl
uUOuI4zu5CHVqw0z3WkAbIV+FeoWw3aDEc0aYJgpYva2bxQRWxXeT8psCh2qj1TT
yyh/9zD+2SzHFbreSLaY4WGUtNSAABv2IM9Yu+eFQJpA4E6uocBfrFLQ0801F/OH
HXudY+dVqjb+7SJ8XbSnD3M/pTJvfO8zfid9uNPmeCGhG5npLFNHn2TBcF+yenEW
wShJxjWb7DakI2Kejen+l7F0yKWxALrUM3D5zVChc5soWSR/H+mOSdJrNkgNt1gW
qLYITV8cvK6u6w9NF75u+z15oa0vjtbb5XdpKL0LkMucbmXy9PHplhECpHP6bM9e
iCeGiwvjyShFj5i8Oy/dPGHW5apWnbjnVaxn8Aef5RPWRlTkJtrFjaXTbJU7A34n
zfQKaBBO9i19jFpDh92wkyFLYOVD60X+tO2BFOL0f6SegCYIFEL7dlV2DlMm1TQ6
dhJsfEczThIfocVj5XJ+YT2JnKAqtYbS8yJl8/R12vvXMs+DYxuT62UcxdQGyDXL
1h9ZkNM+WVfhvB2qgOLd6ffggMQEC6HO9pTRfdfrrrvV9/yOUvzlE0ZJ4KpZUV5s
FUZ+ElSWJRhz13mr5jlYQ2yRYNiaGGz+s1uS0xfHklSYE1J5R2FpjyNYTQcvKVIk
+Hllx65xnB6Bz5bb8cVXpcyZdagawFD+k1XTaIYdGffCyJl6ovq5R3R1WQfDuB58
1e1ayKgVzab4wp/l+R289Cjb6L6L+aIfhlCY6gbIc3IciNerjC7HucwFpMMxupDF
9Jp3FeNUPCy9zev1kWFQXsYDZcV/kKh3k2D5/ulkrzu8g1uY9P6+jAN1xd8yjAGK
HQquTEBUionZ20Oc9AE50xspp0wDQ1NPgPAW+X7Co0fLp/Jdm7blMQROOYs8imdZ
cRSIIoaw/49tq+7I5GWuwH503A//qQUF3/HImlEbnMKiEpPMyGhblW+xU2hZ6vsh
lLQCf5wBSy2QVrU0S2kGdAHcBHlb/yNw4mtzG4F1g8NE/3oHOjrq/r9BZzYZ8hjX
OB4xROvZdsfnUdOhK8ZgBNKUeQ+E+9ill2EPYH43zLfQqmZAKsF8SxnguZzH7CTR
gR+96ibg2o6NCnQ0ZoXU99R+BO0lNRpdIpvKsHJB3Ik5ICWPMIgX9m9Ufe/8YE46
0RMEts62dWkxhmsuYfu4QcT0PmVoT+iru++7Rbg8MVctsyuctqGsBRvZ7VfXmN2G
sNcsYxLsTXd3cAlcrX41WAMTROXXKePMp7nto37fZS+Kz6UdrFZGDPqmUdP2aMWY
vRUlMNmmwQ3fvDAfdE5a1LpKDngzXlLIXpDwAzhf5i6heuMZt2eqq+lsHX3FfgFu
KY0ZcNW89ufn6VG4oU2dL2aeION8Sq5SniifVoF8anvQCgcpfNur7x4Kxe6GaXRI
vfKOHLhBgZ2KQccf90jONsWNDTsj6hTB1YOBLdUptU+c/MaU5zy0NzrhCqhmOROP
Hf7O4aYOh1K4I2IWfrFPa4Qfo9+S65/1bT0OrycnW5UdfkpZaOc3zYZsQr2IIA++
VpsnRz0KKk8rW2yFcJ1Goj6o7LVfMTFl5aYS/uodxUx8DTewH4uNjWcZDR2vXYT9
Lhm1tvMD1cH0jSlip32VCSQtQUD+BffzAWNWbcyFFQzzSEHb26PPDWfkldWu6acT
7H9G1ilVQJw/vBqNu4BR0OajYVnjxOmasEV7OulZPAiU2QH1xLOXwKFrKrLOJTZS
8EWaqs1hfM/uLtWU+zfMBR7OaHyf0p4qCSG6lhBwm3DkxJqse2FXeWk8fnHbihRM
Xr5E91RpBzjfslFy+6EAUjX1w6QG/qWEO8cYNswzJnJjJDyCTnPaWuWMDcmwlGqI
cdCZkLdHI2Z8iCHVBt3BdNzfsMYdrf9Gjm2yA6mR7+mJstlXPwmisNXxp1Xmkx2S
Vs1wjFauKWs3sFvU/9BGmprBxXl6ATGwMOmh/XnrlQQiUe6caT2/cOXRFN06NUxj
1L6JtsGBERuFyTH8aogOEXNAHCFAhMihTjy1F4vMM+Ab4uGiunYoSEcws6pDGnPo
nRaUN4X3MOaRRSR50PQxF0B/qdtU/PwHCnAITyLJuVlVfHHKUXn45R/rXOkJJUMN
KZQqyhVDUFQu7SO+L0XtIV+rYcu5tHpIeNMpP7ZF0FcV+cI4IODggyigafy5M6xT
1Vofi2RPTIKOGrJnx8M57hqrCk81hK2QXkmAwho+S3aXzZKhRf9QGltdeaVRz5BZ
EHJUgWiLsDRYLOfX6F6Rk9wRnMaXRU08npM2h0vPXSMKTZBkUacBgZNwE2jqtHYA
/vw9KnupL/PlgPZlcl2SKGTEB6SzIcxFJGq/KZ9PIVx1cZrDhCqgHwpnhn/QpsV4
ehbgR9eyaMDKV3/IBFoMQGeXTJxzkuV5YVxOaahgl02OOlIbIRswL+O5/YCIGT4t
+jrLFCO/+xJpFDpqnyLDDipv9+wYk+55dykm0b92OuD9UKuXJjmkYlBz54pAsAXj
Knv7x1AeSSv0kFNTw1WdmIrba5W9d9CKf8maubJXAjPHgrx8+f2mGEVpIYdu41na
5ujbQRSpDseSM1++shR3OX8dlAOqqftiKA5wmteEtbDDrqIajLl1/FneL5XXeAFt
MagxmVMmA9+vnw7g2HRTiG/iEI6SXzYj0+NTc0QxlyfIwQ6+RlhME5OLmnyIjA7q
zhbanja4na8DfQzXcL+C6ypEVbA3+4ysw9h5UQBk/SEAoTNgZJtUBrGEZsXLsFHd
8TaMKv+5+5I1jYk0t9rw/we1COgWYQeZPHWpZJuXwFSun7oo4VLahOtwZwuzlofh
Cvhgi9gIrvLqbKeVJaIqP0C1V8bNLDIQxArU9DWYTAlshSIkZXmjTAUKbQCCG+Mm
jsdhgxuvA6X2HfvImyvPIA0SV2Ej0AY275rwY3a7uL//TqnJxPRpz/psKcIdxYXg
UrOwNfii4mKU1NBfVBVn4GQ+0EcT6SHkTo0PMv/xB3GdfaXHAiH3GxdBub4cv/l5
SvBxak+Hi/sv7pf7H1DCIcQGkjMQOFmuo+7DJ0NUvRdFllmDvETijzDSFTO+pJS2
THT+wooCt+B4938qEcWrMWgL7sRoxjv00lBROJmfJzwSitYEycXwZoMjHIM1Qk/G
maABWvRjyos7l+8Uw/muDpkZJ1c08S7S8hDo/hXFNR3CJOpWt4yfYjaivpTeP6SR
+YbE2ie8NFUFfq/pJCZrKedX5osEIbeYwTwxJrqnWuLCinym2iniaiRJzoNg+Zvy
b88NYvWb6sHfoC3yT5lBvivcfY6WlZj0rDPhBc7BUna0TZYAQAxuYZohBVynQJ7c
muk+st2bVet433HHAMdwCcWuQdDxNSqlBNTuLT3LctsG6G6QNqDURyWSPXBPuh+K
3XBsg3RhCYCa+3GaKbtr4lJpWQKkw64rvQFc5W4L5Y0EyxtNnqGYAzJEf4W8bPMP
3m+h3YvK5HmJXgFQKFC/bSGAwKllgjKf7ho1pwkOPOxVDDGMA/FjpPTq1XXjvCRr
DceJzUh9pwqncO1n5spHXluCayFi2D+1vtB+tdtseyzvltsGWg9jncXj3Qymt5uV
6B/xNaLb3tOZo8OHL7IJscL7HRkz0RWyflaQT6oq8oJHHvt5JffU+r2raGVm51Im
2CtIGiM7FOnRxppsi/5mWxoo/0A0JiR/66EXTb/HvPDiStWOJAZUrqqISlAOOY8G
/gAnVSaiy76j+KXIB1dIq9k8Ir8z5qmlpJT16H0OJ/UuQw/Rgh2HvnYoAzQKf+aO
bTiDkHfuvo5Sc1Xv/VisQqiwUSiiaj4ScVrRsxdRB/O8wbrNNky68N8Ow2KYe3c6
bdwscLkp3rFdr5IXk7TMZkJVo+GkNYmyryc7s8jgGVw=
`protect END_PROTECTED
