`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WTr1yTfRyUiTQWza9jqHT10iIlSjYJAj9QJBLVqjrNXDxQet8pOnplBdyTs2IPZz
6W94ZqckL0HK5wgzUQ4J1pSfT68Ih4EOUmLtOAKkFJ9MHK3gKzuc2t/shKQjqUgD
88gS4It8taOKRk2740xOzBgOM/PHbc1Bgmt2qbTa26MOII/ThRKikeCW1YHK9P6f
XHos7ZXPINpV5TvNKw8gK8giK/9oiiVbLd8+LjgPZ1WlOuwsgvIF0+ITUJ4mJavW
spBVdBk3DwmbIU/R2nIX2ndKdrM6T/5Z0tY6FJJlZdcQoB8gMYR8VoHilD91gPsx
EOo5UZWJOP6FGpbNWx5Y8o9ePGdFt7QqvYaE4cRKj8M=
`protect END_PROTECTED
