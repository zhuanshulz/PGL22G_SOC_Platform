`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J8uOo2OWR0PqfRmuKo1resCyjML+4AuarNMs+ACVH5z4nY6mdANCkqfTXLEVK6HD
Hsdev+bu8wsecL4oVpwf+ZhAYSQ35VjqP5Mo+rLbm6gbxriJZ3Ay+9aR72OkiPuN
k0PYsFN+vWUyXL76BCZzUfMesFx3CCD2KqicICgRngirQ+Q5BkWg2hrO76jnGKEa
TJ/dMAx2cwpXgviciKCLFpbYtbjpNqWDJ/edqd76juds9I+EMyUovHaCOp+r0DZV
lA9L2ELgA7hZTuuckjwhrW7NpDvgTndaezzlQ/4An+sSGHDSa4rclqLQufO+SaVR
2bAcETkIEdkLotdilIApky7piqC4uF6fntXv2Q0gWWZ1yj7/lpefaBKkq9ZKNxaN
iOvc4xip/TqtmOWIQYDiPW3eC5elpDRokrcC52B8Q+JwPXRkoC5AG5+PLvZj0bVL
DQ1Y1U7YJOM8SSX0qsHc41YeLR09oZMrJ69eb347tKNks3gEchyfz+5MyeACbF4a
XxIHgvSlrK59gpnygiUBDwL3qVm4BjlmHWt4ZmglWo1hU9hXZXVPrHZNr3+d1bKC
8PtaZF14lBs7HfI2jcrkCWoB8mOPQODi3AITx1mrlh7M1p5n+8GYA/i25awpbVIS
f5T+b7f34uIiFloytRDMw211/oLTWSg4yg3FSJkQaIvRpBkhNsdKj9o+engi21xE
sJcelxvLAMcV1rRXe0TT/90pg8DO/HcxEY973lNFH5U9NTpGV1j2q0puQ/7Hu1Et
vzi863eYXGESTJbyJDacmvnqpH6qPw9J8XSHQl7Y0B5A/JndeZypDsQZO/BtDX4+
cPxUNrfg+LfsQNofBm7Y71Xn3vV9fEgICb236ayByYDYUY0McZipt61PUMdlcPhq
CKucFiL3j6b/+xrI73NvmU1ZSYoffEF0mZD9681iS5HxaOz8PB1UftblG2RK3hyC
PNZIGtWZmCORZVJpR6YjBdO1vtf7IgmVGngAuWQZ491B/ouQqxSIw0D1PItwxy5p
mkzJYBYN0xgXEGyZGSm5rMBTSnw85W0gBXTuTFPRay6gd6ig/b4pAfgNlW7KSafr
IyzqJL0mAmrJ3gJSxKPjc4Xsnn50XuImKX2a22l9n8B7SQlL4xduE9nKJj6MbHug
VqUWhdEWzr7LkJzdLcUwTtjvzWxgdtJop9SxHx48tCelaxgkc3LxKhxhNMv3tfzZ
MWDGzzSKXHqlqnq3Jf/Ua2Of0xZuaeGT9Itco0bCgRZMBOhV7q0OiOcgITQJM2M+
zQq34cEAqaIJWtVWcUJjFyKcXU8H0HsK4YW8CeRfbeEZ7+NzqlaF5oB0vQZLy6nG
0fCA+xttSjLZVhXX0efQQb0vxjSRiJ2VH/o4ts6JLfDKCMLhuI9dLg/459zRgZ3F
khZZSxK6XXM3GoWsLbnkKZ8eJEimcaw98yLtzlJhOjun0aa0oC5bL8RB4jNs/QGp
iLBXT/e7sv+K9bZcqsfOYdYARbI5DBizKQivCImrv+l6Xx41TJC3OO82iPxtDzG7
RHQZMv2T+cHUFibY7lCYWngEmZUqXLGE9dcKqhvRnCtpT01fiEbZSFDaDy3pc7VN
u5SGNEPGYw/WWuamO/O1sUaHkpRprsqSHnWVyIhcvPJ4WfxsIlzLkAv8sMULqQjR
/jlx1d0+u7LgO4gR0zqTSWqll7GiGJJXA7LSzFhA/hdyekHWH9nBSXPGso+LHlZb
DIVGvBw3vLGanYXkwZg9xA1wfY53MtxvoCYhRzdlhOlsJ/smO4ceJTo60CSxdG54
0YeKZuaqrcxzepZY1MF84nIwkJBt7x8UDokkNk7yHusd4ZNeQ0bOxB7gjziXkOjs
0jOqiZi4yKjuVBFZdFG9zXY1Oy4N2gGtgtHalS7gsXzzo3eD39Li60pJ8o4mV3Z6
vwxPoIuBcPV7vtvKIxq5ZIXHakmWRZAsBxnykFbn53dwEpYXYj2/dzxCxIdo3f6V
EoZGh4vNmzfVe5VgiHXww4Tw1v5rmAWIRapyuPtSDk0bqN+gTJRbvCPQ9Zl/Kohh
xL4dBirGN+c/Z5SdAbgwUM3a4RracJCaLkoe/jUnGsgYlXV5wUeaZ0wKo41+6IUm
Z9VkUdbQxAipbUvq3t+f/aH1JWv2AK4jb6WTk2GnqaeF/ORH6hAs9RGeNLbETTxT
/1xzxqHL0WH2tfGdlXzHLoTetBtonpRxnNVmy9NvdYgy9yUzYDLDNADKrj4h1gMg
MtYAI6f+3hh/RoFpEtiUfs6C4bhWUPJLKaY7pHJl6lytctkBD9fIY0lxsJTtfSxL
EkApCfct/EKS2b6Kt2Xal+1y/oOjY1lqdsVKHSLaUTOHZfMYSEnKlX51ICtST68R
svlo2fGtObZQBz/Ndh76p8JzHbueM1LvbiqyqB5gXtJZ8odWmXVYqzxI1+fYghSd
bouP3n9DrmslYS64/O4Ao+6mNRDp7pJAmCepU7bXZCY4xREPnwfw0ZqeSPH0tXOi
WjF7D5fGtF6vm0323LGlmYTs6Bz3V6pSR34pRW5BQeJIuRJv16EyL4du4gtA6fAj
dz5NDyTOdowZv8TFPdDbXJxVfjeG35sXhg7XhPSbVaGT0t86JL5wNwvuQubZ1Xs6
qudVghVdosegYuXbLkBmf0664QfPq5qmpGcgf5sdAlex+aV6mebaLFGg/Zj22n1Y
P4Mqn6k+EoVGHNlAcDssQFV0jkdEbIM9zw63HEf1t7c=
`protect END_PROTECTED
