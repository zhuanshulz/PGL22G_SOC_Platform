`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wmFa8mRdzIQMZXtFFY5aGZEjBIRbUYhqEBJBwqHzv8FZwSXyz8IetYJnrtnoONS0
MdfJ4XH4iPaJSCjpwmHvWDo44r5KzTCIN1FmRDmo4NKbsuQDdsT+cXrPy0Sc0OPH
b5EKLv4xALbZuWaCjFwUovj6NBPX5F6SNqROI6yK1wJTkmh1mNfRdI0MNGYrkuYy
N6ZvFT6R54JYgJwfLIjXkufxKtrgK0OjhngubybfFBXKpM+WJnFUwAJrA06yIjj2
bETxB1ra6qcPsSeRrKJiAnQsbMCJTr1CH/qYlB1cHI7OrDr/CN+2Vc0vvTfbTmOj
BsUaso6IvA2HGFJ1yb8IqKKesHcZ/udL1T2SiBsz8iFQRpTFqjWut23xbk9VgGCz
iWjkpdQXQbxneV3KJGD6gJat4tjdG5Enf+V7C9GGrdsQionQ6J774VeEj/7+IArg
yc1zka+Axkv5RsurXiYK+HXI9tHVhDdrjsAWWD0C9+z4EyD1Jps/A7EsDfHdQNL/
OnkFceOE49OcoQmU/epbKfhKDAlsbhYsG7VgagoUaIuf/LYVWY7bdqTwFocRJR0n
sX/8S5eDF3a7X+i3RqxBxBNchfnwCw/whQlYUyIUFRtbLpc9CHJ7x0aNbkt6cTLg
POphssefG3GmlpmkYDqo9pdt2BobVm8fTRY4SDvuUpBsp4yXECI455eYfJBHFLe6
ITLXjtyOg9Bk4IE7uVFE40849EGBfISW875YF1RVsrMHd7WCnIF1sMnsxfOBZWKt
V3coniL72s6lv7Bu38fG7D0wzfeUdzs5Tb6/UvuYqlNOxpr13+1N7nVUCIXekPnB
iIoH9shWF+YdSQLL8NB/4GRAalj5w8CUTPM43a8rorWfHdkmYbKyqxnN0ZkLR1cP
f4hSy0YD/ifyUDocbHcwhEa1Zyl7+8bpCRruaGOZWx7FUEJen83SkGZNNI8i5itq
HqcAj3/Ad0U1ShkjS6fWKJP9ZwUA7oi0WZQrWlht2ezSodUcbpAvNY2jEJHuy8Ca
X/QGripK0g7HgXooFTWjdT2CIQ+9Pbc7ehLgEsthiyRtDGvDHbGEiyPnBoybrrJb
frLUsbi+tBonR7TmGzPnbkojB13tOWtxODsWb1ZX1qJGLd02qhFZU2ZZkKlBC3RH
uMTTdnuBQuidpR8Sito4YdPWfmDNBTjM2iDFeAfDH/vSplZWUJh6pXQwJdL6XjKI
bLGNjXayrc0zk7zHd8exltEqIluOOI35RIRV229i84jSnl/4H4xxpDKsGytiFEo5
36Zr9P8csYASZFtDpknoJbIMRlgPMuTqWmiD9fyAaQgqkv4Xmu9iCbPj2zq8vv6o
xXMSwT3W44LwItCDHE6+W1Bc8WYL6rywS5i9IVUAqLBIo1OKJkLUSeBJeLP//yoF
ci9IQ37bA3M8S0Wf2p2pAJQ34CxHXrQ9Rki0/k4sL+mKRFqTOgx2uuTMpbAdpAb/
ywwjbTkXrUdfUn7vxjrB8N/Oppy0DgA+6KOVJdUOhouCN8LLvTUerZodeynQoMiP
y0RVvzj3rWPT1Ceeg8Pw8hhopiHjuebXqRnHBOonueeR5TqbEGbJ2L9nuiINqAq0
jI/0tsW1FTPaQJj7tGMVWi8ykLIbos58gWqDn5PD1p9OBnzR4QKWIWj8wRnV10EZ
WSq0zMYLE10HlNFIZECaq0XpR7k8IqfiK/sK6K1SZHdkTmG5vP6lK/4r3grDFi8/
8wEGi/59JH8Se8qUmURCXIaMcIzWu8qAkjzp8+kdk/XhEMoqFpKlem+dGkBN0Es+
kijINOc/jEfqP/ILS1V5kel+4qplxVe3vS4ACmJ14Mw9R2+dYYBSyx5nlMM3L7Gc
dfKKqe+X78U5JjPQJGuORfGZu8j+1nASSSZppSiB7VWAVKwl0o5Uq2LHuXTpTsuX
47Kc6M7tTYAmw+3PQQ9e0KG3pRvCvWXGr1dXGsK1cJN6oof+m95FSgT0Vt/RwQSe
0YIpSByAkZGXQTTzSvgTcCKg1IzQPRGZ/sVnNvWgkTHuLZAZv3XjAz/AmJEdjwqz
/pXtGnuqtLyj5eZHcvOBIsBllsGSEs/0ealOZWsLKs+6LP+6OkXGZMzClx8TGFQV
acvrS3aUi7Igd2gBDwadOzg3s7FrfZn4DxBbmejbug/8HIrgnUN7+gTE/rFOpP8P
iO7AZ3mTNIBw+55cvtcFZwLvzN+veVb1kNzqO4OJL7AAVBL61inH5fuUH/ye2nK+
hISHXFD46MrDM0SGPDxg4JD0cYiqVRS0X20wCfddsq3+3HQ0i4XPRs/oHxgmeyVi
7b+AD5U8YlZTxbUj4CdmnEGO/uc66i+3A9wZ0g0jiyXeQ6R0U2Aev3tgLTXZusxi
d5wpnulHucqGuGiIbSMYjDH2hJHgvfMNNm/ymjO2Km2EBwpY4ZvFgTIKBN+fOl3s
jh4HtY6HjWR/p9VgHDAuoa7NRW1GBfDvtilK/DvyCiuK10WMnPsBUSUE0lHxgY/W
027Yf4/7950V12aCrhKbfy13BAI1gT8WlvzKfL77ADWv4b0jr4MkIWZfdthy4/20
Npk+D4aWpMFRevY//vUmWKCXkO2KNhSRJZ7ce3K/0pq9d+/47OOqVD9KYayRM48F
UnwSf68YYp9hVhxzcL/iSflmQ0AGlPVvnToN4N7P4MhEPf1sKSJob8ekHTyT5egh
qtkzxkeekuyV4WUoGJ95DgbbbEFG6oMHKLsNDTNtwvFFWEJvNfhfOQ8J7Dhahxjg
QnLp4XMIXZe2ddos3GxdMvkCxd42kTE+r4l8En5vZdpR3aGunfS/RDqDr9JZapW3
1eokiUfFFpAV6DWzbIAOe+ytGCls9xwILEkS982qT1wWCDZ4WG59lTkSSHHWyVev
l/9fygIPUV04FBbcwWD7R6671nY/ERwd2dIlg28T4bs=
`protect END_PROTECTED
