`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Op1nTOyHcbQMEDIrYbbv0xOsgQsv0JcRaiATxyihYJLe7LOccd4m2Nuqpk7XhT4s
1UL+qHysPoLld/k8jGMzSVuBnYh3sOGdP/L/QMF4KANBQQ01DsetA85jC6zvGYZb
Q0XVivH6mqW+SS8RJb6B+nJDfpMxgZtaYW7I9z8qYxWsJBX93aZUV0XrnLBmNe6w
RwfTgOKBBe2g9auB/1ukDqopvJ40brTiFiN3qWDWIAaIFyxSO2knx11das7Vvy8A
8bBHJbjw/BBc+7paU8NIx3Y+GkRNif5Yb1MeUy0PQNDR2dWkMLm+G7zSKBFfDBeQ
5LHSEiFd0jGnReyNweBZ6/FRTmr6fqjYOSCactmiPcjN4FrOcXWkHMXl/tqjo1E7
5tlRf7l60AgKYwe8Jk/7ba398yVhDlbpHFKHHXQV/m3j2y82v229RR/jEP09FPu7
xyGkjC8uJB/F0MOV2TM4OyGNM5ZI0fO2rpB+Me1vaPaWRq5l6Qu7kdAN39zBL3fC
DRfXtn7egRo8FhVMcoBQ/rS17Rlwl++QE3cfapqSEO9tO6yKo/h8Py5MY59aDO1H
zpAmiRFNjUfE8tSgpgXK9+AQ3CFbiL8Ut3W0Yh2D7XyIVHjGGsiBJ1WSDmG4n0sK
5e467KKow3GA5RFhnHCl2uqSJ8ODrMVoaob1TksXn8Wgn11ssKPxb4nlpkagVcTN
ZR4wu3sg9H5aoIiTGzGraIl3UXVI6Q34iJkP2Fp7Hveb86ER6kc1WwEsd0inYtUe
USHm8v7DaeBDDBbIPQ+zqOYYMdIkOc4q3LftXIX2ymJPcfPm2QUP4oyVZzhsgHUH
ZGCqtJyniFZRSPkMCeGCc/HNSfk329FMgsbkTR8EJvBqB4bexot0Xew8hdMBTT8O
1LZFn1KbktVxBWBQnf6rkWTiQ+EDn9NDxTshAxsANR7HVaEdElfj1KgFHkgJLrEC
7zeD/Sn1B3J+rye2KCwM/nKJ2yf+subKM0AxVR+AgieZOzJeKMxk4z3JGUV75zA5
dwilHrLzmx/8uElh/DskvK1SLojgI2hmeesv8DP3aBaLW5C3b9bAEXO3H0VNJY9m
B624/XX4I48/Za+nF9cT1RcceH/ziqC6lqkG0gMudLA8JTPLqibW9i2ortaRZNR7
C9Ju4t7jrg5ryjkLOMN/DRYxeCMFNtZR/Bo+iENhbLciMo4L5a8yWWg7AC3qv1Gj
6jgToyOhK4oIK/pLEqVUDERtghEZvXK1zngwMoioprSL1FU2Sjc/npBp/cYpoFQa
qeXBwDnNao8xkM9YUSE8nnbIHtaFuSpPRSxfgF001Rc=
`protect END_PROTECTED
