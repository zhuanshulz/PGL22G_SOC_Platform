`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
84LJbn2JQIWnvu8N94uPl/wfQzCMWdVjGF1iH1qKx6kxb6cGn7XWU9AhXB43NxF4
qnZH2P95EWtFzY60D5cDKc5WvpeCmwwXI+/NQC9eqxMAMHBSw+6j9ONVCb97ypsH
G0Y4Y8LRnQbxpXA5ixd6sxueF4MLaetnTzXyIuwrHkTD/nYCAxa5zSTnDWMpHEGl
dvGqn3/HIB0oHhE4b0vgsf+owGMn/VJVmt6uHHi1ONARPrSOBrMjdFVaBalzVTNo
mrS0cJ4RM8Hkz6ZZp8/cKgRoTCaUyyADbiTSqK+MZR1Zi4SqW0e6Mnf3cN2PUB79
rufwDr4jKd1UPvd3KEU1vmkGpoo0KUn1pGWK8blJMtF03oBpanBkEBBqvDIWPSZB
GNce2fZQKeSoj3WmkaJ05Lc13KbpSopC8YJNe2tg1lS4Zh+3rvaKiObGAVczANOW
abb9Y8C+Wvk0duUbzZxq/aF2QB2tOLgh75N7kP075sb79HcasI9hWBlWkAA4cOVM
quTDKH/nBkYh/horJjEmd4feOwXYGb6NpsEa4X4kLS/gxUh92pzRDbo/jxlDl9iL
Y220hA0r6ahIu1OK/wo33Zv0ys6Y5Uh5O50XRrFuoqeHteDAq+ijEG5YM+d4AssM
zdokFpUWsvWYB62uo7UOPaExdaCjfYmZjeYFQxRcEhzqJRkU3539zcJnnOLMxPVu
UmK+nE+Z0ay/xr4xSX3BuFFWyL//T1jX/vCQ/dCzUpJwX6dL5APiVCdQQ04Cu683
`protect END_PROTECTED
