`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eq1PxWp4VLmbrq9vc9Ei9VXX0wcwYdBBMZRvaQ69o0v36sYNl6lkE7/mqO7Qtsd5
2bo0EJwR+d517ezQbnvd5XK86rsgugaKKXFhq25f4btOdHTyaWfzvtKJil9e4WEB
TN/mzCKsiskbW8APR4Cv5V2fz7cTfql8ca3FGq/yf27fuIJ6e1mbxQzjuI/ofTz0
4FcbGTWH1kMsLerP3o+M4V/m+B3aKWM9MbkeSEGn1UJoQfYmjpZaoGfQrlVS+jZg
0j7zbjsCfX4idmZBPtwqIqdGzP5Cfm1pGf5LqkM+uwEa6MiXeQCF03VdWkBRRwG9
qccVvxJrNfNVg5O6O8W6T25/Rh3SE3Fe2n/LvNNQHAWMDUb4iTqGmyvm2O2R8j6o
4uuRfB2rlXSLq5cs4y3RdWdQYvVKMstj2IC1owzYPYKzdn04MB6t2ovSno79xkJx
ozxo7Aeei/EaxanEJkwrMnzFsNV7SvTJtq4LW27WEkpYTgUjVyze8L8d8+yu13gS
btEFcYd5Lgk3ELA9KdZ7BQUGZ3fy/bkhAheEI9Ql8zLmNCMTu/799XSSBlh5CA+v
3c5PQhKzifEeu3n8MD+GLnTFroR7UOgtM9Y1Mnv2e4G9dFXCRE7fIWf49dLQPPs8
2zQ0ypx5f9ZZ0iYAyGUwVOHyD+OqqLURN8ip0XrodvxA1RL8c25gbnQDBKLkbw7x
T/tStzWEw1tbxWXx6h5WlcXMe4wfKNUu41Wwc/DgV0QsORY3+IyeCOCTkae1o7rj
51M6uFVmM/k/SPX4MR3ebN1a14qjWVOEhQjltdOciDb/Wpgci3KdanHGWF5HZXVz
xOLA1bqZYfeg+CxK/bqD6jvDnV4SNx3nOZ4yCdfETEO6Su1PKO0kHWe4OJHRlHBt
4KkFfC5VFUZti3H2NJ6jLV4ZVvKW75bbjMhlKSZ4+Qpcq1m/kvyHirth9eJmi7z8
jDuRQMnZDH3zMNrf+K8E1HrUvf1XLSxf1txaBhGhyVPkmfsnHDpeNKQGXT3SqLGk
u8zhIkx2wCy12iSJULI1cngi64MQfewf116caGrXAczuW4OjmBUFaQIcEZLFjlZQ
iJTW/hJQTqe90vG3daUWC7UlIuQrh++K9RwIV5ZrmThGg/MbVbUxd8wEgmHZnNDk
43q3H+lniwot7/TZMsGs7ECdtR/ThVWd9pt2vlXaSz1jRnxzhb6BfAYraiGoRVCZ
k5LNXy9sx9Pj5bKnizloCm4fkJ2rzYZLVRZ7gDg5ERY=
`protect END_PROTECTED
