`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
55USJTXlndzYtmG/EcMQxOVR/FubGwehQUDIqjDODZ7a8lQ/SqqE1b0wLuzXGVn6
ZHSxdTbf1mzAlVi6roAMlSTcKLQJVQ096ln0bAqAKk2RbcMpG42JIOz5h8fyzMnk
P1aTuQoRLPFuMP3vRwOL9TajzElIqV5RQeAAOVsULi0rmJUtsKxqmtoT1SwT4FMV
qpJXaPWqIQhOIB2YiUF+k6CkO8VrxdxGfWv5SNk4Ut71xN66gUE4vb/2nt7ZLnEq
ZxBp6uTkRetoHyCnXxaf5U+39Vd35qfTFh24KBWaH+/B3HoGafweaBWJek2vfdNG
qcvsamdeG2rxj95V9gUY6mHPE6VXyedE6kfnLoS7ebvQK6qKGHnrlTmPjHi9mEKn
`protect END_PROTECTED
