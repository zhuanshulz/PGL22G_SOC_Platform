`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/Brt8+R1KwdCNSujXA+9zItX8z9XxSxFhk0HIQaJZZZ6vCvMJCCbPfmfa/0mvQir
qE/PhqoK53gKGpJSPdsVrTrxU3HI8P0b825c9vZmeqKiz7i48701OkX7R3oh+mLm
TgWSNzDEeSHfJvay57CWAbkL0qNlOcGcAlg+Oox2/5XOxY3VtW6EncYNJAguLwKK
WAsFRPK+5LFCEOfVrdcAbIBVFJrDfG28SCRCtYh0xcqd8jChrbXro98jpyjxM9Q0
O7c6jfwPfXInzselfHN+VEHH+jnXZm75hU38kGJPuxuxdkAoke/1cjYu7ezP0iiZ
ntr7iA3CAgih6YdgXIPoR8pqX01diZTkTSidaX/0sXKsRi6y2CWvnAvQ0GdkwKz+
PeT7cRc0ysY4HgOxrKApnLNShHsJfGS9uo+Z8NHrgWRt7mnOkmWq/V3xk8VEtrBc
tX0pFUYdCd6sGM1urIFbZ5D+dflbFc/Wpy0Mk9e85FOCV+2UJMYEDKVpUKRQoMhr
fGBJ67hMwfgKrMrwFtwyTj+0m4Q9+tTg4td1+gHG5nSsQ0ETN1j/g3SCS2GDgxoE
ENaSWOW3tfFzd82QVw3jYurmT98LIPmWDtQP8c1uV93VLIPvyQbtz9tNh5StUf6h
7EzDUE77fd7taM6vMrqfgJjAKskXwiGNlKdLFOq8RedV+fSRvFn3UtuCDR/a9KeL
mgeGtQbWo9Jcdbh5xt3FOigjlhRpk1YQV2ybiRIyVCbghJ4UHe70qBvA58/JZdsk
CFH098dPU28pNwLLlOedf4+3o4a0egBzZYmh6muuBKIGuMHgDoL4+g9B8+YzHUUD
p6uDwcKcW/8l4+FBr3iv8FKOeEsffyBRdS9hqXqf8o2kqzOW/hhxOZjiv3EexBJZ
RSmdWsG7/1nZQqBsjxnnSQ==
`protect END_PROTECTED
