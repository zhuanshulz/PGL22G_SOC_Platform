`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UneXhDKXCxKjioaGnQ/+pNXkeABH69hstLS78cOBVaVKbJUDoVjwpo298KEVFh36
wx/YxJj1RfckQ2s7Mfffa6o8TSutf6Deho0sQjGB9n2jM3zJ0tNDZD7K4uWaCVnS
ZuVQVeLDfzKjBPigcIgjvOKlgeci+AJ1f42wfBAq8sShMAglNoPweYp7cCtuKkhk
OkHM+JhXgCTm9QoWgRQ/f50VcIyMtMnlLpvUZ2KCGLhSh4MuC1glX+BpIbyThl06
437xU4uKEILbbiB81MP+V1f6QonWZeyEVTjpwBXKahVVf7r9e3Xxeomf4QBHGJKf
0KLybiLPfHX5OvkSArMgPVD63mA46y7QOWbFCGEm4tTtwFIg/c5LQDJ0yfVqkzUr
oEJ+wuuZwWQgBYP0TDd1lU9bt+RY/JAuzX+pZrzEcPHd8aC9t9T273IoO5B8tM8+
kJcoo3hcsCSbzEiog49eHg==
`protect END_PROTECTED
