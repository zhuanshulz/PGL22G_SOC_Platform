`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RWUgA6PdY/Ou05XxHFmKwVM3oo7jpC4MdDJsaUfbfBY1cN14dD6EGrNQCMELILKf
Y+Ofa2AaKowefucTKeyiOmgJj04aj42kHo3kZnK0VF6P/EC/NYf1LOSw8R3YoiQ8
Ld6beRmOzW4XoKffHcL9+KBVgLMA92qKYntnosPg8uxiueEBtMP0zAUwA9rwzQvY
z1fEPNOh2SdvrVM5QdXyZddcQ717NByoOuZr7TIoBdA+uUXpYfo6UyOf58fqOAMR
6AsQsVN1lrzxTXLYc6f0AfhLLQVYDVu3D/CZD4l9D2mRXiZUOF7NvggQ7/HYv+5B
T3vbaA7lQoVoybIvEb/LNWCWnMaRsKDlsqWYsKzbY0E=
`protect END_PROTECTED
