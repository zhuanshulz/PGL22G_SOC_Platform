`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EP94aZ1yC4uFXDYoJ1WgTR1vQIONfrCCDcVSzM5x0aw3h4yKKwxh+4vPOsJMncO9
d/BV7DHbPTZrcEmjbc7R9KFhhwl3ZuLnDKGQGgWd6Fndb1Xe8pT0tjk6Cng6/O46
IEyfRKu15QHQwAfHgD1tySAC3wCti6bfmiL7BWO24lyKYQzuNfM2iiRC6DjkuJnM
EiR8vdholQifu8VS7gjnz4bkTFsK+arSeBhFozjFNQNr0iCbFHPf6ASN9xHQPGj6
mm0O97wfP53h324aF8iGn+sCws3tqQJWMyaI4puZ16psX2G479NdlXaTBkiJEhRX
Su9koDlaSxTJ+HRTIe9n7mf2ClWtbThBwtJ8MsRKcXzDWUBWA6y3STtJRV8V8VxN
j6ehKrsXti+wEl5qD3tNyKRiQazt34JD3e7HaAPS1wieeZEcOyL0RtWs//uzjgCB
R92PgPxOz9Jt4B4ZiJa96JG1aNtA37CGDOvotNMUN/aGd/1cQao1TcaZ+ox3jGBU
QcLXCcjllaP1eAr3+E6yBu9ZgSqwSqYRCPEmE2qVvYO/Y74WIWsskn1fW6NknvNV
2W5TzXEpfHf7e9i93fzaVE/aqy19Xu/37Ew74d3d8SxzAfg5mQoILLwdNU1JNGSe
7ja5SGP+B5Cpdt2Si8BBe223+4i5+QqVvVx/Yv8Ws2aMQ4sEAZse3RmXWKy5/foZ
55/8vWJ2ngaf5rqjbsjuWVXlJz5K/Vi/D2FpyBQsfeFULSRPy6CiqA5O+/zEDCYK
Y3/VjsXSDV8xz5BWnJ7IHBWvcJ6XhWcNWz7q5af7XYETg4w/gqS3npnBg+3xSv7F
UOGhghq4UPiykjx0aeZv8m/aak0RPBTRksU8sh2F0uNIf/OdzHaWNN77LMu/fQSp
foldFxXJne0Wj5lz21D3aPnEsi92nvLLg8PQPZE7Yw3j0crmsgn18Hqwj5iOVtr3
AZ8oPLEaAJ41rORejV2gydw7yvhQmHdKjzKiyjKr9WdI90tHxxdwO/rTR9mQwU9y
4HmdEv9G1mxqu9gzz6q2IojCzr0husZq5lU8rS0Nists9grBd7BysoESggP22kLH
DualE19xgUsZPAnj8nGwiB0EdlFy1GNeOnNMe3sXbRXGdF9DDK/ItqUfl4WYI9qT
zqpoYskyU4ogzDkbkuq54eSBWPTfiqulpxbpkTPR44fECvyXlIyLqZ7DwHBlNEC5
6wQfsMQDav2+H+nPoOdygZ4g9QbzUwKXMzmHyKQfvBmi3Ysrydr8K954mNYwo7wr
Jts6QA6q6zDUId/RFwxCd8uRbf7EsDV+h5WV+m6JZboRzkABKjvjAr1Pr+2YRcxh
w5r9NkAACdzyTwoxQhOdJ2br6V8MAMPMdOJ3X4B5Hb/1Ryg9s0n5otGQc559gu1X
W0EMzDNRohbDxNAWH4dWeD99RhPkqd+bi7iTEFY38O/9b3Y/c9Wu7oumZ5wTMM6W
hZexyAaVTxGUW1vtnc9trpxLNAGhu2N6E4dj+DFduBs2HUMgMrn2ybej6Ug2+bkc
yFbYXb2Q/lixIZCIUfaGqAHPozyW/SAIKjph9n7DaMZNXwmYS/J5NjnTfRZtUHli
6OllC9mfe0vticpXo0RfXpB3zdRboaQC3qB4AjI9zWEeHKvw4E9vqWxlfoEfSuZ6
x/2mg4XtIdQOPei9p9QY2AAxKNdMUU7Rm9mWN2rZ4lk90XirD8fPnEcUzK0PTRLt
v0KGROlG9o+iVebxUk6zeVMcCUmoLpMZifkst6WzUJmd/tDG45kN8UKWR6qrbaIQ
3pjJe+nTgWNOYxjmV+oZJWTTWU8iF1+Vm2YG36+KQEnjMbrJAKq5ErEKl47zoGuQ
IlLT5qHSJG55WWPawycT/QFPvfYZTqpV9OsC3MMfu4k90Pj2xBV8caiDKyMzz3+Z
aue5sOfTsTvRIlD8gURoOIG3H87AiCI4m90aNMR09ogKnwbpWElSdWx37PtyhJ18
ydTHiNAa8wBg7hZmAyjLjMWcOvDCTxHz+ksGzVJReHgh8JSAChzx8J5rIqf0tUSp
XcvXjR+WAERj4fzrbWppwGVogX01l6f72K2k3794H2Mf7Bs0LdtiEtCk4xhbP/NY
P0QQ+LvERh03dcB2g0Abch5yOWmyHfnGu7oS7J26Ea7bo2RPIaUHhA/nyHlMfOQU
V/ZOE3dqesgCtyJ7pqKrnqK+OtoHMDDEGEZmFd5cIu/fkVvX5FSTBRoOFaW+lguj
8ii8K83QujfYuf+e1zJ3Mn6j11ezutolLjsp2A0IdCwlk6CfrC/vfcfkF7S9dZZd
hJ/vmvPun4EpAT21TYEgTGbPelkHU8UNeoqBnw7DAyZsHoO7XFKFx8OF/hstOu6f
7mnF3n2twB/OlUQ6mc1bNbVxj+HX7ptq/JWZsBmor1gWnGXpLWFp/YdixYPcShRn
n9SeVx5nXJtneY29XHBfPrg2+iV7r3cwCLeI/hO9gBvqb9v9WJWJE8QsXNKAp2Ue
ZaUWkJwiw0LH/HKhptvucvbXrVXXnzNvT13he++0/SH8VHGgy/5u7zaS+Kcjifyt
neGTtcPw1UepWKLaP15jb3jW2kuauI+1VTBlGBixUw+Uq+4Ke/urYXujPl/1oHmX
Wr8dGmMtpXb6Lx4R0L86rjGjf2IyT8F8f46I7faXQ5GAXoc0ocKGvvfZ72E91YGR
Jxwjr878HUpN6OsQ71tQi8UJhgl0fwtGBkKFXfHftuUgoQ9t2V2C9PbnVAhBNQjL
n27KPxnmDDfP9A5ivsqa3ljfc8pm/0o2Bs2+9TNscnF2QPTZy/nrbPCuvrmPqMmZ
hZwissCLAqr+z09VcKqjmeeGDZEn9JAF64nvyBkGfOzkx96O4wA+B012+84XJY0l
`protect END_PROTECTED
