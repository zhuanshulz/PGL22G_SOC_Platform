`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y6ompQhMkcH7PyCubMFZWHVt9r4mzwxMfjLIwGURwVupq0zfwmmL+y4l97QZaqJ8
08zqoH3KPogiubVO3XVm6fC2/6coX8qg7JM9rgeuDxb4P6/LMmvGtfoN+9tJH55r
Qfv3+lMsJMvc7NPcE3WVePfDnDp2aZo0Er7qsElCUTIWRx9o9GhuJamPaeOaBcgg
nYImg7bHHxShXYz3US9TGNnkXsNdVkfVa/oNwUZR/duBWWaDOaXio8pr6uEG2ClM
R/Bxayokw0XTYkqIusdjoHgM4rtmJJAAhS9L8udX8BPqmPEH6y+EiF55hzwjeaxH
czhmC8gC8hC5GA01Zsvm+NjzV4y24xavyR0o5P4ETcM13KpZFnqSts1yBp9OXve9
+T8a68dUWHMoMPU3df5ygUHEoNn5/tQKPwfujGniZB9MVbBph1m7fOtOCbq0vkk+
O/rCzsgiYN7K6VXOs1ibcQn+lMngUr65Eg8pOYho3Ixzu/dpJ2d3EZtPgaOzv6XN
sdAEsAOMjAiyTaHODeOM2UFQTljop2Gw5lS0Gz4MMPe6Rkpj8DoigLNF6LY75rtT
FSYUMx6SFstMvHVO782Q0ZriPmpdnoztNpkr3Z4rl/2j+osVmhJQ8f8JOfS1pDsv
u09CwQ78x0h4AV35ml9WrdapIQwxHgrCbFaakHPOZKjINWAIh+rSLBmd/0gjPcz+
WWHhjEZ/ZimLi88lnDE8c8raK/8ehGpBPlvSBIz6Mj9i5X9znXFN39yH3PduSkJ9
+eRtfArqmHWMYSVTQy+GK09K/m1l0aqAq8GnPf+6bVy7KxIQBhlDLXB9pcRqs6rl
M+ccHUh/lsaFTvrfXiKaRBM32tknePH1NApNqmanUYG3T7wZe3sxq1Fv8jR5CM4i
`protect END_PROTECTED
