`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1BfcCUP6/SvoFf/GDUFiK2OcGVTlfTqFJlbuzw4OQR3eDemNzhqPo41BiE5kPsX/
J+Q/p5v0H6YNJjmw0wGRoUSKmOuS6xkaraNz/GjVyLS+YgQm937w+orPYIioVrsy
hiPYnXoR24o2sby6sDyUxeTBPFoilXP4V68sPpD7QG8sRE9ZBVR8do/OiaM7f1U9
fReJ18ywnff7OTGJa9X0i1NUgU5cWOEr2gLdULaJ5z/ArUIQaNoq/O/flXKFgaMO
lyZ689eoztQKqZ8tFxK0uVQlOs3AImDtXJPUVHJAxg0+mB4nwRFRIAAAIkdUTHCp
SbXcwU01HH0gkx2Jv+LRS1WECzbHYb5AaRtB0NRDapgAoX0InupqLAmB8PKhN9q7
5ZmRQekk73tuRR0nwXS/O5UscTEdSqtOsdMWsGKSnUjGcymwwmPRpj9vmSDMBKwD
88wQJPEkA8nRVwV8CxZCYwVnrlk0xfwPT+Dzx5wyS4Ji3/I9GyikV/JubU2wIhSq
t0tAVo1tkNq+qnnvicnYeOg5SwIowrL7h2AJsGxLYLHlwCsRA51SAkNbhXAojl3d
fFz5+3Wh+cxsu+6EG1GuWlqwtXkEki8HeVmK0JS8+8dHZrEpJN/N42L6GDfTuYh4
RiTez2PhpAZOnf2wbXXdSIGaSN+2HGQ9VlHfHrzkXciFj6Kp1ptUhIVuvZAIRGJ9
6dwTnBkzKOILUJbeh2c2IzprJXef5z5zL6PVBcE7WeKt/fZrQ+YwPcKiemD8vZz6
IopMfhiBTH7it9pwBEkX3PphEmgruTgzIq4TjhCs1q7hz8N3XmJmdpwiR2OCOwrk
Wyb4XLHguaYUAMl+Oo+7lBCSrvT3EYCghVLYYLKm8hgLVg6B2vuyywQoiAs1IP93
/7dVQ60t6AU5R7IpNbCUkJm6Nin95egyV82YVyErGe+/Gi7up3jWGJ1zrB0tvKrn
fRJuyIjUm+1okdr3zJX+ToqPRTmkHtVdzz9Gqe1V18xabGDL8QiLpZLUvWcaL0lV
l9gacLUgUWGS05mk9jtCmSBE5DqN0lUZo5Om7iuVvRkWhI4mQYURz5JlnkucvyT8
Oi4fVmtAO4NKozBx2degfpFOXTDtOsrt9X1sB2KO8yTvfoUq2c5hQ5a3bS5MU30J
`protect END_PROTECTED
