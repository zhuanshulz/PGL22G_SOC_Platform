`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4jPaE6lq6uaq9VXcwip1XJ3u+U77CNajU1bsw31vbOmA0b420JgZFpa3j5tWyDmd
ph5o8PN0JBWOdSd3YM36ZHxAWeNNMTDIaAYJBimQ8aE+/WwftssIkGQCU+3TnROJ
eI4QvtTrx+P5M9qKKvtkmp0h4TKYXivmPAZO5faqyD2smny1TTjmUzWl9OSrlQ0L
eCUpF6dHF1BVazgS8boNix5R09I0lBPGThe2+5A4nmAAtircwU9ZZejPUzVYKJg6
WDdTWUFX2rt/iomKfJuffbByt2f2fHKfaXsGij0if6rrWsaQ12WvbiA0LmgEsjR5
rHmm18DfQjUsH8RKI07Z6MdZbFY1KudRC1qLo2qTiXGGB4VGG2tk9q6UF/xzhFCZ
7Kt8Omr5HHuBcDBHiyVOlyg4fqudC4ZsvrLnkOxlveFZB5ULLi+P5jPs9VDZ5cIy
4TGpPmaHNdRjsAZhNQJQ/k5le7kA+wTMgEOLgHoP3LOL3B/gx4F5w8RZez1FPNzN
q836JH73QeSH68f5oUyffZrS34nNk3okb6AwhwzDXqQvCQhE/Z3dxc0E4WErZLtk
FIfSn2HvhAsmxAT7bcvmYVrQsMlq4RVaKN4psIlv9CLNHxMFAY4Un8Ro8nZAIatI
WhytPDitFS/BTegufsRaZN5djIhiQVw7pEpe0FBk2mkmyp6ZHO48FCSlWYxV1iBR
uDrLWaqGKy0+DIPZ+yXt1jsjugnIFst4BcTe16q8dzkgqoHpBsqlAMv2Os1xfrcY
FwUaA7wewAOF0WmgaXpHwBGJjEOTCev+5yAuI//77scPMmaPxB+29OIkKpq5F1hv
2HiwcorLZyNEJ9+AYC1sVPl3LVxLndnCaI1oUl+HqKh0iKqm8nJL82H0WuD5/OtK
CPtDEHVSRMUygDRgcO5PnULNlbUmh59Lvxv1lV18DOeooVtPOxuxUOSYCXCQw/ma
crLX7odqwpIYmYnNxhRrr4VgJHZecCdGNI0yvDRe+1lBNIxH99cocHlVVRJKSbv7
FynmrqnS7D9JoFHbzXqvxYdPK4h8BaDnPNByIapJNNxDSwdoDnSOEagyLSkXdPbx
E5zAeR5lHgi0wogu/tWV8TWy/RlBSUY9pA+BJ3AM3C75mWltAp55nbN9qMYVK4WA
ai/Pvw0IioN09LyACyb9ngkGLZO5VlR7399n8PSskFH9kWFEWBXn9FCt3g4f3bDi
2U7EuRz1rXsOi4AJ1naa5ebotxWV4R37GqJPHLr1XafWQ5zTDJ8c1pieptkbTP7M
KYsWwFUhaT/3BDzNe+yWkhg356iYajHZp1EjvcIHxIk07lzJvBOIU/vsrcMOUNBO
1VXF5C8lU2DnFMmj4dtA66Lt9R0ivw2ydkMHTyItzVIVy47nX/ormDNrJu7WdxQc
ThfUWPc1H6DS6DH6A5JBgwc7DIh5x9KKtVEsxFVuif8fNek2BQHmWMtVryEJYhhC
N7KEp9ImLOZugrAG/ShajVdyGx6yb00EJQ47r+2C1xemB8oF/AtSOkFt5QHfOg+j
RB9p6fOoTiRWYt7XNbkpDCdSnOE2WjJV7fqdC10gfiBS80vKER9II3a9IurTAfSX
t1BGeXSlX0hF0md2Ly2ve1MCpXfAF3bHmgn1YPoiJNz87e2pnxG36AvMejKftSTo
XCBmTyldCHZAz9QPklyAzHJ/2V/M1NhF+mdo2BpJBJDrUe98apn/t9/+9Qk9UkhI
KSGHkyHI+e1gWwnawE54ZtIvv6EEJwoSaWru2gg7RV26jxgp9TrhQw5rWczjzxqp
J07O8294oVAXcCEI0giXEYmEkjvXjMOy4HyOYk3VZ23EkaB8BhSgw4S7GIMgzUFH
ioWJOKfjlpVvZqzymHHE7AyOHfYmk91R5VfFJ3NIVAKsUKS+Re7VwNukN/lmIDLs
XmaDQObKdRz5JXeH70Kw9MPwN9WdqeN0UxM02VAyLAhu4KXDLmOFsxT4vNSX8ky/
AcfwGSet7Z2q2rQ3MIc9IMX8y2MZCmFCOIdSR7jbGICzxeLvlHoxfqPlsioNAz/5
dSdJJAMztAD9qWo2DYEvG5eXhamlyDZJo4Vs1aWhG028dlts1Cv0l6O0dAsxZBOL
dNi7BO5sYC9J+CtOp2fGQ0gRF4jjcLsMMD0wxZw59+xl/d9Xn8taqz1UBiC/EOBI
BNBO+zUPew7TPvoz8jvHbmzyGAdPgvubfVxPDa11ZijAq2WTBAeyYdKK7PVRSwus
T4y9jDXuasMv7VXn3hpU5vzsXa6RBYGPLuXTo0QhODRJ0EWburdQtIFe2i3ICA6k
b+pfPTp2HvXohEBc367/ZTpX+mDOCf1smWPCVU/Q+5PCDG9gnwjbOuZ9/BE70ju9
mGsnALjVyjkCzTWuNwoHbPG2dJJeaRX4QSNKoJxG+kkhq75Tj23NSBgN3jshj03n
HmEQ3OYm3AR1TFjWq8fudP1zmRXlJDDPNb2b/3asOmD3hbLCHGmW1GzNua3lagVp
BUNCeqLdMfsNW4pvJfA7iFqixdv31PlVKjchgYAYPr1eHJzpaLIYyxgFLEoLcBz7
s0zLWEydQq3Q81iNI8La01/ShWznNeeWjA6JP0SiNSXPpjhmDjOoys9rnjAntIY3
pCy+2/lrRQ8m3ph+b4yTyGPViaHB7XpbSPkpoHtnnpQggHj+8qudnzlTRquYLuhL
/gpG8B9i0/EveJ23HttC8M6bUr7oEKd6QEzUOh0Vf3OAJckUwfetx1gP44bJBncb
PUrnyJ1jrg2gzEI6IsmOaSTwLU9GgqJUs4ElBHmYnGwJqOi48TLDKZc7mnzEaqSy
NRdHpNPy5DwW4lI2UU/UNwIPEYV8xrpWm3U9mdHJ2MsncZI59+twEnfitBjA2ZFI
KXissKWanJYp1kl/1/wOiMRRx2is5YBbmuhyCY/brf/vFD0uUtaDu/DKO4gWHT4T
xASsIEIpWmCrt73cD3BOSBPlBwhMTiAyxkuE2GekRKx43EOOmKD63RMPWKbra5iT
nxaKyYpxO9jB+aHI5SdjTZi++SUlMWNaUSjT+ONHPgeUqQ7PDRVCmMAt/colqWlj
A+mdU/lYoAAfkEn+RX9kgAPUo63jec4mrjBL5sqPoRMh1zjFJO7udXQJX/VSDdMT
L0Rtm6/R8eB5weOL1mUZWlrIkk4sPU+UUSYkwSU6ShqGZkqyLCjgeB+/J0PRQ3WR
qwJzut06nqXcYgo9gHI/XOaZ2CIvXmpPwYrVayZ15e0WVSBN4BBNcYUEN97tMUPT
N0B1nQycONWhL7rAIMfKowWRQyTBwZOPO7XTW4ngE3Fcve7ydP5LW0MOTgnHSycE
/nKqkYnSuxxZKmJPp6WUe9wI6BVBJoHl+TfWJJCpcixxaGC3vf9hQ2vXA5Ce3NyT
Aa11NW1+rXM/fwGRO7xlO3roLaP9R2JFnAM3JpdGq1I1Ag4Ga4V6mQD6mH1fq85K
aq3DJ9SWrI3DDBgv51SJ29Vllc0EdVuDapSJwIXgP+EcgxFcRJdd3pCUx04BR43t
PxkC1I2mvmGKZtF8G+omk6zo2OluKlcfbVtWJdhIznbd9uOfISqdTysf5ZfwD6RP
UBF2G4Qhy17CbdkiYBiBGh9rmdwnHTmwcnK78ANDUuACHfgOjYPOgvoDXGjF4brO
ihMpkIv066oKT+riwaN6QpW/URO2wI8DzO+WAYYcPpxNNyB+RaRd6IieO4zoTqIx
gL74fqZPBxthlqplEpfxoUYCPxjlUrj5sYahVXfXOpWJnpY9M1toSXwk8lAd7e5v
fyihe2Tbc4VB4a2MVBj3S1Cm++q7BrctITcqkrI0ZWNjlV4cRykjSyW9iwRToEpS
3fD2jK2emxfva4VSEo2qWF3WEcxL0KrpaKzZh4v18xuGmHjttRdBRIuEJJbtdVtL
HtiNRHl0M6ybtMwsss/kQEbyPm7KNX4crcCts/FNPEavtKXJR51Q5jvnevYMFIjM
FwFNtMCIKaL7KMoOdo2xsKsMQWiw/1zZ1m8I9GGqaJykmsJEvq10UX8wNGbHu0hM
KOMalHsgi/DlOuyBDRdi8AtRWep4q+3jCfa49MIPbF6B1sAFvfnZBm7jY/wO4VeQ
R/DhvLEhrxD0hdaWKOmvou7/MaWs3oEP/9n7OJp4bT7dBkoPT5FvssMC+t0JyWNv
34XMiD1X68eRTBmh2t4Ms5ZyiaMtsOALjZO45PXbrWpf2lM3qz7C2NucGa5J5azn
OCxjOrdre/2sFtNv3gWb9BJ9OxgMA0WwjvftWdFu/N9zChp8L3jgMO+NT9cFhXV1
t5KJnDlXCeRrHekTcYcsWz7TQ+mA3OtQscf4T1X181feWRn9IEvB57MZqcBmKOif
+r/unnMoHtFAhZqbPeRCpRhoQ5RkvYb4bx/WE7+XmvwzjU+5ZsaC8HXLoilc2W0y
RrlycbShOCGt0XMUseS9AGeqc3zIyfK1W0220vyJWfpMFI8npAstAkNXHJgOvjJC
Dli7feEiTjVdFkxuh8B5jROsmhT02e5tbg2QE7HojH/9/PSaTvOTK94WuA7h7c8e
XwnR3gZew//Bl0BK03+OK0s/1EwFSSE0uQ+s+Fs/mXVsfMOf8rZix6cVN/xiSLLG
J5541hu//klZV/EeNOL2ShxjLBwBOOLMpIyRTvRNXkljRXOZk/wcfbmGUkT2okXt
vgVA9AYD71fMcAruaECbmIYNS543XWdaWiNdmMyu/pFmoKevvcd00XDMudrGfe7R
9UTiQ2D8AXvLV1yLFaROEGL94NsdpLqN9K/kY7Ix0wKlP3i+VUjPdzEaACuWplU7
3Qmvj1vbQxMl55hVxVxfmxc3SetzwVpcc4tidgEM1CdYZOz300IGBmXxYExcB21N
4w42DNIls4xkgtvER8s6QaRgFgj7gGIAHkgGQ2oe8asKiLPwmQS6K9qxVzldNMcS
d5Q12pIBec3EDDOu42EoOZ67TLQAtg6yoUFjekS/IG0OP4IzupeUP4cCoAjxttOf
weC5umB+u4F+MsM0keB8PItxBUqn0+hPO14U4WLQlPj7TR0F5Vlnd0VZFzXzGFyJ
7JQ8NmmT9j9xejquyFx0PavJ4t6qFf2by7yvxZ1QO+x9d6LfKRttxtDhbSUdZYSc
iX/OyE0V+00qLDXD2o2ZbqmvI21iD8wPPR/RuOHBWw7cKkUfV/un9mY86+/bNlfD
XgLhoLjZwgoh9IqsecTyFUlpbwFf6gZXXcvub2JHy/zt+qlKksixXKEg9s6Kx4nB
pOQazSegRYG1KjP/vydQrji980QlwaumHAV1atme2e8plOBUU+Xo6BKzWmxReafa
Hm6O8J5acl6VTUWCDd0+8l09MkWmdAzEnXwiYgD7LOkyu4n5CctH5wW2LTBPzrqe
YIF8FJZazTh/ickWp+N02ZQCudCOL6Grrw9p4VZQ/HHfr+Gc/6JHONzOwdymgBet
Ep44P0mS63QNGcvQWbykA5/N9R7j+kPdFqHDoTPG5QK/tVa87AppJv4e8PQtd95/
DtWI5qp1ip1DdKeO3X18r6N/S+/2MwF7eI87WkF7Ohq2ZDue0CN2UxFof2W1WLW0
MNuP6LpG3AgqEO2JoPBMwPvogV+EyKAirHnJyBEHJHwjsVJQprkKEdXxHwZ8q8PR
m3JCE3tM7EYDjQLN9StfZG7vtTkGug5CoPBEJSifvX3V4PRieXfqOvLq04Jrdawt
TwtlcKZXhsG+BpJownV8d4We7dvpNLu+v7P+1q/7f7woPwRec/74+pQQfPMDR6cF
J6xPuBRDYJOYscaNFZ31bO8kQ1D/B9GQ0m7Jo6BCfLeCr7SsdRsuof7yRl6jaHPJ
9kB8+pekDFxtVCr4QiCbp/PiQrqH2t+s2hNZ34GZ6tK4ddIUIdwKzqkZmvcfp8ba
vvN23q+3VL/pv+0Yriw2AZvZgvPjewUPJKu6rKWcz0Jo+GqhsNEFbooD9nl4gy8W
kX2P04EFGiWefXS+cvrwHcDtmUUaYgPeP7MysNB0b6H1vCe3SmAGqOmeJ2zIjD13
eIHqIjDjpOjSeDGar6tr6zsZXtZLkker9io1HPeT/BTgTPK1d0Al7kswmzZweQCl
E2Cy+xWL+3uiubM7uTSkEhsCbl8aeb+sb9/2x5bgsNjEqA1xLVcpAO65xIBS77Mp
/EyLjx6R8QqlBAEl8Mon2mmZd5gubTF96yyYphhemhqbXnaSytBVgXAy8PyA3ase
MYZ/AtZw/uo1PtgOQP8BhaN1cPh3OFIqsktNmsqgs67AvWnOfE2mWhCHhFLfuRMR
PbOsiiOi+TrcRVLdRYCtP2njo41eQCo0CWw682WITMw8xynvN4OfBS/M6QlP3igw
o75XmQ4nVckjU1CeVJzb9M3GuPhE0gpmYi44bpQbtHrUo8m982dmdSc2Ord4jYs/
hxAEDbONXt32OhY8XQIpZshq4FsNUSe2m6cKkm1n2JWyi8PNAg7i9CkBzg4XD3yf
8e9y70HWWSzcuk6CF9OWarjZYzqqA0L6yZ1c8wk8iY/BZ7DA1s16kfFWGjJTRCWl
EbwYPLCkAguZH8KalVquaCRv3aF+TP6VxvNLrbt6p9nsLBE52Ktsii4WjMoZYwsI
2IJgb1QWK7IIKd3Je6BU8wXafnL/ejeo1HpQ1/YnzNo1YFyVMzwA0POfVbNbsREH
MduIb7oTEsfNuMV686pLAE5JTFKmIqdYo390FaWRymCKP67U2lWcLLkuP83u3xnj
tdPVew0K0hvESteLvjVVrqSoqIRA9sUU80q/WjdIxlF6FaOVxLJDHIyWwDeP7A34
HjrSfaB6jzVF5zNn5+7gWwiDYiPP5SEtZQMA9K2z6DUZX56yYlsN7IDhT5XcjpPI
+XKOiIgQ3Gnsh+45AphpGF3JWGlGK7gzWzrAbhNpwBmWw/oS/OR4vGzsGRKJckT6
5FRLygc/49sVZ13JGwy4ytUvmgJv5U8v7l3qGcza09di7VAy8cV3gCjT9qawTPmG
a8yaCJMYPC28XNkuEnzZPyk/Cueb5vLzicePSTh/WgZKeUB1HpAx/C88GoTcvjmA
KImpxpuD4gUn7pPKM5EMjjxjSNTtiDtKb/6SBfM0EVRRvO7vyNCyej1WKPyTqDlR
B+1kMfDMbAswwsSA5k+NBQmf5sL6DTrXMKkfIZQqyZJIBUC/TZMBqx4DZJgIAquB
kueewhxM7zD18d/JPic5HxRs0AwzFBK1PwCSlYsc2D5uPS5KaTbpk01LbKPzDtsf
DNlhzW6ggDG3JRcR3FWToYcIyTLQJYVxkVlVTuaZ7ffNZozbVTsBEqx9p8u7C/Mi
KJ8P6L6m44/Sx2XvLpDHgD8P4IibEuduJ3g+GDF+mLJiuY8sOxFaCjthDlCpvrLt
GMzXDYnqJdBziguc4TMEaM9DYtS8EFdF07QSVWXF0JUg7tvXMyytWoKewt+ZhlhW
cxeIuLspovW7Oo7kUpplksPnOBtLqkWKm6rjcnZzm3/bjmgGbeYHokZfdzahzBMV
FDtz6Rsa7sq1TQifN/b+Ourm/8cWTxPqSGs6SLWl4jIW32HqtZx/QwSzlPmPTre4
2zkK/1ydqiBd447GgKfrkRJXeCdQgZzRceNi2Io5QRNK+g2xUvowxYFr0hykf6UF
d4p7UxRFWgDEABhN7f6MHPgo3YljdXJIESBnxW0LLudgyyEgq5D1R3r5UvHx/JAp
5GwrkcvD8tyY0w7IrWUaEPk5ZD7HeAA57GVUNMRwgyEi1OGFRxkMtMP/1AGgjShN
jRBMg+x9LJBgmotRoOMQSuKcSL04e2gwhy5IvbKXHuZRZzKJXZ3O+C8KLbrPG4Cw
tFY4kg4+hyds0ZPv7t0iaufHlE5sq56/upPMqWXkGXW6uzExHdPq5EWxHDJ3HVH0
APN8LOI1QLu9QkVPdOe6T01HkOY40ApqWr8He7B7FcWBo22/os3DvAmPExTi6pk3
RnTO0AxrbWJzPz+1XPY9FDTZQImvfzH6m8Hw7ZBXlun6WZhEEilAop5U+cI898Ug
FuO2jJpT/ILVc0qIqeW4Y29j7QnxQq6xR/AY2zUDchWkfK5FxiVnFfXFzxgtizLY
ubUS4wHWyKWm+aw52O5/t9pauozTq6xTPrycEqKP6FyN7nwH3wPl8WcxCOmVeSbP
xkixTYykDLPr7OhoScytOzxl/ZMzI3Ln+wEebcmD33CfJTzeFBX40sVz2sTGMBLr
RP+3Fp54Fm6POQMEW8FAKJieuS5vZKlaixjRcAq/CRROV/A0SdGsCGTvuPx0upgt
wysYCng0DKZtiDPTzdTMiQm4k6HKz+slwd0fzQMcL2BRnHWmLfrYZyF4jxDFzk7a
N2K+57OYW3EonyKs1MiwluxAhglzuvP/xDi5qE1N/iBR41JY7W9m770hikza6Vmx
dprsJhg8VwB7E3TNm+nxHJAvNONOWGNIQ2SjIMt1G/se+xiO08gZxggK9E0tVp+/
65PT7Ja+aURprYcAGjvMV3oNA+kiazD34OqKm8hzAgmqpVBn/MlPATH22zMK/cjD
4D220ic2BKq3MSzujqHFnA346EoCEf1Rqka2IP+yrZz7GPl8eK7AxjmoYgvPPZ6i
ySPA2Yx6p7RtUxU/1GXX4MUuHOczCKd8AfYgMvyeczGnt1BV59qDSTG4Mf/pgftq
nRmGj5hsXSEjxSfekPmuPKfPB+d5xbLQ+F9FV+rm9pZC9Mp+EkdglwixDFOqHnPw
yHzX/+Brz886691x5/6yjTsmh1zcG3jqPwnKZpYMHs+507AT+KvmJFagPZ7Hs072
iusqPZWEHdhmPLz704AOYbXJOh5ZNj3+FpDXNFLyhtYEBrQdsSHiB/hqudp/QfcD
t+cadCcwQPMFMYippaAAi9Oo4lDFLW3xUl5PICqp+XsbAaf5QPZJgc07hmDSBLmr
Bkv2EgeWoglErnu4Uo1B8fjYAp+MkBuGNPuYm8aIGzseXLSh4V2uOc45l4nNRzht
q2jGJzZ1TtyX0QG3SzK3LxzyxWSRAWeB3SgP0Px/5/ADVLj55tjzNPt3a3KIyOjz
DZIs0M+IW1RTHcBof0qdfBz8k2ZqgFyQUOnK3o8ZM9pOqUTCni4eeII2J0UBJaDy
MxSbSh/x+8Clujs7RisUbBIwc0KyvZa54rdGLvAsGXG4vqHObeGAnKuP7BEAT7fg
8HAdm8ZZqMewYpWjqeWVaOhzsaIS7YRRDmePQS1QkwEspVA03ikzz5XZ3ERLIugU
jh1JAolWszUIWOraG0emO5e6bMDf+poIp9BFVUOBublB+oOewfO61bv6v03wgBVj
r32IwFTPb84Ak9i4xASmNskzl6QTVHO6UEwyoRdqs2t5rdYnrzrP0bxNRFDe07KF
wQZUf9HDqU3Xu/sDwwjK0Y/MS1cPJqyH/B3mDHw6qWFTu+Wr3D/b0J8t+/qPGrWn
wrOXgDXroXPx18YBboslzViXoVr12YxJvBM2Mj08Q8QQAxW5+eXv+1YN2nzVfK1i
Ivcu6mo10gUijBEkyP6aB4RSaZ+v4tCBZP0bBfcuNNM2aSHyg0hZiqH0akqBQnGX
GNxCIj4vmiy+BsWRGrZ/N2YWskBcZv4ywa8HiE0ycZjOuG5PqZTAR3gS5CTbslDg
QQ7tioNaAMAnWA6t+Ob0Oa6S8t+Qtmb5NliBwwQOBrCgFxaOZTu/cITK4PxipTYa
2wlilyoSboYQMLCC4u8TTxzdI5+OS7tkiofPb0ZA+PHrtC0czBV/zbLu0pv8F3vj
diJaHvkbnOW3uWhrVAk5sLcc/CLpho/cxRqM6RnyKfeh5rEMg1ztHXZm23tW4Lzp
Nz7jRxsuZA/LTKPBUJswF3EHb6Rtesu0Lg+j1hV9f14KQvWJakzVs+5oVrC9No+J
ECdOSZrtzci0Hno0tWS+sKT/Sv3mV27jlrhca00uYqI=
`protect END_PROTECTED
