`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fF03QqycOSZvfNXDkB7BvzZk+ILB6gENrmiN2tUtVzo69qULV6g4HLq8U5iUN3s1
hJdn87m1puqHUltTddL6Moyuyx5UIoLMHLVO+NxLN54q1SVGzVxZq+L5u2i+GUbK
/SFeEb0+ELc1w+CRdgaIjm15StorY5A4x8jDGaz/rMJa6wuRSZGDMtUkhYTdxN0G
VKTAPp3F0iOxtDse38RKTFnMDNtCeepukCiu8uhgynMXd5pwQrcwGKZJu8RznDA8
k6Zc9AJZrCxfGqo2ymwclE7P2G2m1MAKlnIi/uQRzXpr4bIqPe/wIWD5w2kzMhH0
NFHA4aWUUVkkFCT869YQX7ttMiRZ8iWZWz/VlsMMPsgE7n2XcpPczoBQCSRXRp8W
2HH3/G24yb7vx2UMvQHa0JxzGjlT2QxbLIIMRYfJgrV3qdcOVOgp6YhYcQkD3gzw
WrsTRCMB76bnivrVPk+xACknIS4v3338pZsuDk6TuSBGZImxRbDORZeIt2gJ9nkY
0vt7grcPi2xrx6iCuSBxgGRQqlgqsEUgzKJ84V8TkebVnKVpVp1pnzBEbrDhhweR
9jyogp80Os4jYdThEtzrSDmlsQYM69hsBoqhtNl+1ZMN0hytmQG4f4DMLbxmLKUe
Ll0bJ6cyvSnN+v9vrv/NhEtC3ShJFaWvpFdnbreoFAnED32KOntdCb8liJ31BI5l
`protect END_PROTECTED
