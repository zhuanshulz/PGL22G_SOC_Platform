`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
waGUSs02TraboBXQEBan3IzwByCQIhnOr3vRjIyDF2zw/HxBPmrqg3/D3UsjIdBo
qfq7e1T3rUP3/HKlepRve2nDjQ161ZhD5eQ0SPhWVegQn0gWdIKC+ikTWWbk/pp+
HSEw1+fVla39Am75dMUP4IGI9d42NgGjrm1+aHaX2V2dTjdSgxfMd5+dVnND9Ue1
lGwiG36Cwgj2t35nFe3QBnI1FuSBdtrAYlT7fSQI92KAQ4ne6qbJ9Rr3UNZhhWE5
rJPyKdlZoYbx3TAk8x04DBj9AYS5Uinikz9w1RItuWH4lebMUVaB0jxHQ9UN7IjE
IKUXsEuemslHLKvpUNq+lSxVl2DSBT2zXbV0XRZWGN7AT/IiSk1je/1+OLFHABzk
wsLNigArOVIuWPnuziiTqZwLEH687VvPF+9njb5FjbsiPDKAVXvkzXDsAGkVhQLo
NqXN5SmZ1FLLGrW1I7Ca4twdFZFMcgY6JMQa1g53FVVItq374BtAgl8WBpbAwFK7
6gIOSVLE/rjj4N+SXwK6Qg==
`protect END_PROTECTED
