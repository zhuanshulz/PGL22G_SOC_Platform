`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
psVoQkQJ6JKbig73AYJTohOnTZ+4x2O6lGcuqp/2xWyUTsJrC18Tjoy88G1i1vNq
aUZ3zRTDMCccXi/+VjpfGSUq2R4vfG5DNaIWMZPVAYyrE7e35uajMHLR+I+TKR4N
RRBmDsPJGrqWeqYcxbizvKWcMl0NUVUALLsW11Ofty1/Vwf/onkXgMG3MEYn9tAW
H47JKQcks5KX4YWOb4S6EY+ceK/tX2jL6+gQD4geycqQfosw5cboAesGdnYdT3EN
W4a3dXbF6DyAh/lapJB1Ifx+B9p/ZXo/7t4iEf32VBkzZnVr9sZxjSpE5rPbJl01
8ZUpIv92EsEgs7PRMGNAprdtEYaT/xKcyOUyyW7JqIkfxqeCoIZqN/ltt0+CqnZo
j86luh5yOL3GFiGyDgyzn1lodt9C5sa8ku3Nx9OwFzptrlJuKd6QeIisLSnADflQ
4KLALXTni6oWUmB0DlV9M114wYxTg9YCvDR6tI/Y/47+qgv+Dcz8EF1qK4qAXGAr
XuuBTnmM9UUgYllqFyTmzb/aOXyURdG2JnmmHRinvOGcU68FdUqpYeHOn8Ilkmlw
/Ty/7AUS0PiV6Udin6xwNYzMCKHFQRQW6p4CBSf92r78Gp8sd8HFdymI9yeXaAJJ
/VMY/GHDwMGeEDhSC+ETAo7N3sRhsL5mq6rhnIJQh8cWvRnKvQNsDpiLHimTRMbo
gzm1kYWWB9keLi6XgArrox3D8F2WBb5IzlKzEgi9M9yyoplEtU0ClFMAzGDTU+38
jJoq4CxsMOYPWD+MTLssMkmersvZ+JnwGfaDisfXBpRI6iUDZ7YCc+M5qMbWTDdS
eWnwXhjD8PUvBPR2yXMUOQ==
`protect END_PROTECTED
