`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a6+paK2wSxO0p7KFesHCot6XzjHmXQGpTOFrJ48Fhly9i5P75X6lydZak3TSTTt1
+3+YDmpOQ2DdB88lLnwAWbTwzAycXc8Ry6D5iuoqQhcHZ1kn5mH/wfJCr8VCksZ7
wZ8cF9mXlRfBNYRXBE1vJt/bzv1/rxBf958mToT9sTciNVunnMx3AwOatCzh4wrh
mUqfVbXszNKQkX/79HAD6XV2+O6J4uNtSfztLrJhsj84r02MSznrIhg6nOylFRvD
aBd2psi1o2WcT8Nm5TmwweG9blntJR/cMEWqARG6iU1Rhy2n/0CWyHiCc6eCYWEd
yaLBEzuV3I7mugsbi89B6oIF2m7ZtrDPBgmE2U52Gus8r33YqYdhdoRhda+OOTEB
SI7Ee7pcPj450ryeLWOr97f2r7xzzf2+o3szJe36YVtYDSIWtyREQlCcy2jCTXim
BEfgHUYY+6DF2K6XpD6wS41DU93BK4J2dRtbVXMxY1PWdPONxMz2NUKuh7wysmMy
MmeIOQTM6W+yo98LjYnozZkCUBYD0U2+eOJiNCw9a8w7ym8kWVMDdbBTxR7PTk+t
CV7j5XaE+wl83IJbLC3RZ7H+9tFUaHcYGrpQdD4T1VNMfaI4vIkyy6FkqGwSh7/+
WODQFw8pFWQk80YFLv6O2mEnt05mMnO+sbb6EFcRalj5VBe78JIwzgYAvt5NRvwu
eXKcfS1TsE7IFvGZs1/AJESnQ0SHw1YKO1M/OFhi7RakMZo7XZO8ATSxu59+xoYf
Z5G0WZxyLe8BUX1jOKGmvrFO7EFFA5fmRqMT461o3k4NCq7cWCzRztPCxOk6ezVa
TjFBn2qadPjZxLxs7yy6ETTVyQj06byZ0n+2CmdPt0SR0mo2xylDXgrNYMyZyKdo
4xWiAgVpyWGJi7wlf0tLG6EIDQRnvK1i3cGfc8WRyp7LlINdil3hr4Ey3hQIWWgb
CGSidJAUpGtP2PnBg03++rbA+W7MMeSPYxOaOe/bJ/v17FGnqBQIRefqoPQB8tKl
T5hAWR8+Hv4J3St0xywRVhr9itB/j2VlD787r+EKEK3nKLS2XKRVgt8MZzt7BzXg
eck3qenBVi0OgFE2CqfXdMoLCZHGX3dghdLwYzBOaqPz4zexAdKXQxobzA3BKMvG
ZWOHydjleqihTM9DSJGXb5rEc0OXy2AU2iGr9JlDcOgCoSAJQVN1b4ia5ncECYzq
M6I7QNTvZcfv1abFPw2ZDVggVPS1QDTtRkR1HvpB4IMSlwnlummxU9SyZBc6RMhE
3vSZltHEV/7TgtRIGBjqetGGrG22p3EZPu6Jz1N2oAKp5ppmt+Kkeut94U4+ml/R
UO1f2OqPaQwCTx5ls7b9jXzjnyb2CQJa/uCJVyJP6baEJe7D88dGvZ6Y8+DEDtHD
ZiLn2NSCj4veHzoDUFIwWguVVajYCnou/XN1vnAD0ZX/ceGfmt7kJ++i4T+ia/Tx
B3hYGoYNhxgrD5eg8WOw85/tZ2lj8C/ain5T9foLzVg=
`protect END_PROTECTED
