`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cu+8q/ePyx5VfAcpxhB0zXA+qXyHIbK7VcO0Iyl5nyEem8ETjRaZdFG/0s+RYLSd
k6Z91Vl0x9UizLo6QF6jbTwOjcZubpl68B0uRR9rZXmn91lzXz2ZujD3HrPs4HUN
D6TUS3eZad9u+eVRsQ2Df+yvC0iQ6jKS5f6iWU1L1JkWjpq9wNVv/VT08w3H3j1F
vBOkfcQVUX1KjUAS85ioazcNZNSJ4OFhD+w8+UDlUpn/FipU9tYpoZiS+AltyeR5
1fYPioHzSe7EDIGpquuRftmEChc7dV4FHy98AA+lUPuxBAeL4VgIWJ8+dbPufn8L
wkk2r8kZYLW1tFoRuLDdQS4UjHdGr98nsf3Lojs/E3q1FjLQDMYvgUOcQ3QPxvZr
yhu9PR8UGc5Jffd4jgoj28oQ4wWvDOETrs15LjzrLpJGgxj1t4wNzJgPhJ+Llbrv
4D/QfhpSUTJ4RKbNR7ytJR2Efhp4xmOK9l0MnNchJhb3vkN2m4cEMk9DwJM8xePh
9BIBGjQZ2DFC/7MO+Z2Jl01yMd9GbxrxkWYOcK4vZOet+IXTgaY4Pt/7R+V02S66
EmUmFVTNrwbuy86mA914TEgmpjtWdYwGuo27N56LjGydKupZbv4wNE/UmCixohu6
91H3BJN0sWMnTju/gzkuad330OpyTwtvXnBr/5PlnVYItuRXZTqQn0ywlL0EvqAY
xY5SqEziLT9SJDAe0LOqUzq0SEz4kLFBuRGuVSsdSGyBxCiE0mdvCKQv51zUuK4U
WbWsllcMDuhyDrYdTiu1qw==
`protect END_PROTECTED
