`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YRhRABtCcCgM0h3olE+cM4abbSDL1iN5uS5ndy4zDryFexI17kM4ouyFAKCU8Olh
VHcXIdW6na6YHI0nW6WiTGLtyXgA9Dvusi5aJixWffPJkyjKW2aK+eJCbxbTnlqi
x5OSBqPuy0Rl4U9IFuBS7gKhkWvddciuSd/sK5NgcqiwjBb0HwejeNg0eRaMGcNo
/3TAgOoM/S/YpvyMxwUpD8mTx/XukxYex+zHMEJkW4wlhSO/QIwntkwIzbLxLC0d
Pkq7Z2n8hYM9HPYKnNQYSHRrpwpq5JW47zsTxyfjV9+pb2TzVrTrvZ/Rs2BrQ0hc
2CwialM/kEiYEVsIJCtaccJ7Cklazv05PIBL27LbIw2Zl3CaaGX1q+hG1x9I3uPT
j59Dm64GjfPo1x4mK5gO/l4p7kxgFSqdy+Sf8IAR4bO49lzXBDQZ94vkTooh+Ksc
DxUdtzOi3izVL/JNp38reNx4GgOz7n8fSJSrwXyZI6o+bwxgnIVoB5R/cyE7KF2J
VHxBzE4DgbosavRWr8WhCmqAjdmiAlKH5wpIkrDiiKyTH0q79tJa4QyjKvKFGb4O
USaha+Il4b4m4EEM96NrvEmKw9hwxVg3YhyXpEOYFT4SZd59Wja6jrYdCdyYF0Lp
gCemchXuY0LFsrllS39YF/lmTK6PL3OOTJv/CCub1gweo2kJzm06X03eccv1hwPD
VPJVTaBjPCllCcab6Y1Qac0bNbC2iyk/lMuFt9vrFBg6zmK8QnUKmUL1pXUFJ2tJ
XwFgo5CvqQE/WaPGf6mQ6tP6p3ea4x2EcHXSxm+4ZilMESoOOJvmzAxLKgGGefVl
SvuX7A9wZFJrkh/pb8e+VNDGxTooyE7rIxqD3t3L8hACHU0TmjME1333zxPpa4pt
Xi4YL7bpjzc89b4SUa0TZHL4Gbq9MldFx8mtin4x1Kq3i9znd1wGMReRnNk6mjRf
LMXW9JT3/nJ+HXvQrdKL3mScQ/X0kwO0TH0Ve97l0ABiuN11HD8FpNpKzB6TSwP4
BCm4X3U9ubHC2ERMxD5bkmuRbC7P8Un8M62KCliXmTqGWQSlfeju0cdnhwOZrlfH
TsOsvoMn3P75cjptQULtmIluQcUJWxdBXfARYGMdzXRKonw/7gI45oJKaCksV/ql
raFgZU1bLu4QT12KlnfpCauVi6wQ67LzDUynLfeaoWKp12nV4EFPChYBMPzVEBfQ
o0vzRlsW4eMfdsCy/ITQQNgR6LB9m+75FZF6gryEH1V0VDtJQOqp9JS/tlnZodpc
/i51ubEj9tHBi48Wa9zhfWL8XHvOgukynR7ZIVFIpPt//XeyV0jkGp6m3gEcNDUc
TrKEPni44XB40XhyrMkw1sCMtqv8kmu4Ec9y6w0c4UYfDh1PypkkxdSV0ojEh0TW
Bxy+kERJCyzp44gs90gH/qiuF5g2h+4/LFLKKWKSSNhLFazGDCooZE6QLWrsv6SW
ibn41nlgUuHd/A7BS6pGv9BZbkHpmuGQyfFDKQAhv1BkVduPLcOvrpmcrV1ALyfU
sVpgtO7fNjYL7wH2vlU3Bkkv9HQAA6W+cxgc7QwlsJK3iYbMff2N28u9x9CkPXaS
KBuI+75rbZL/Brjrun7/93dmmVvgvPc0zO6qGQkXwnjKLktIoKIB29N1s/nm9pBV
N9f4ePvDPGwXaOEdEYL8iHlHqUjevzUhKKg8NC19FS4s+kTCAkVxlPPlaYTKvzz9
NIfV72Yjyoum+6BgtnN3AzVWk4XHvCUb4WFjf3/MnDRfhW4GYPavU59QoOcOeqA2
rxemeJKIse75hPObzr0NMzvi7e+xLABP693eH6lWYuarvhY1bf+l+jWTK/7SVjlj
CLq4PeOhrprMsx4JneLP6KCnpaw3ziYYmvqrjAl7GloLrSsidN/O+v7yrDJvAo66
tT0jw77ei6D1BfaTaDBnOFswty5uRB6EstPu+8NZXkzIeeem4gW00iK7YyWWPXeg
ObqZTv64kx1dqx6IvjXB9993HnRSp+FV58GEYQdygiu+3HIbv7+n06shDJ8OeQDy
ljAUxfEWH6qUlumRg1JZIqCi5djkas+3ETokqh+W8OuO7pdF/gXaHVs73s4NUn1Z
JlrlFAksqLPG2kS9KBRSPRxgWmFennpj9xjs277MWTTb57K6CxT7lGw9VygyNPaB
+9FBi3W44FZIs7WhSM3o78hAjAo71VUvEl8hqUpqwticmCutywmPFbXd+e7Q1kAm
Xd3u92/NbjzYIyJ6RqE1+kECRxsEZnheqERKY9848BPFrR7fFA0yiywEo2eaUZJ3
qothmcLzcLLl99YSQBswUmo1/pYv5HvJfYpkXCqK04H/wGj5EyU+jh4Xt5sUt2KJ
27v1wMFNQ0v5W9BWK5boqLM8L3ZVuG3V8/wEzZn5yMmimx9HPyqYwefJo5KhATgF
4RyDSptangbYX1SZ7S3sdnzzWfBnTkcrOPzdCFKkBf8zztjJ/hHFGdKpPzKGlgmn
5fh1OZbF0sORobZeoU3jWPRYw1rjC3DxMcppnPjBfMCaKqKK+xrzhYwJs8FQWFgy
rfw52r9GCpaaIh9oA0f1KhAPMcl3H0bn8oroyzj9UbZ339tm6uAq762OLUteWiiG
0XKkyDb+q9VbXqpb1Q8Deq3t++U9rvzWuX4CXChpqCZ50Gj53vcobol5wKHSDSBz
iI89C56H7pwB4X3ADpXt3mnpCd4xOgmbEWpcXui73iQh7LLzvhqnrf4BPk9CyNn1
G6ldaR/eDg/+RRk6SJAoWJeQ4NRvglPvDVSgjY86Zax1N+tD0g+6ahjYvJo/Cr+h
Uzfhs1m+w73nBORzWIm83BAMchvfcGeNv6IciHRDl1EUMqH4cT9iF3XIt9ccwSe9
d5EnbWlNXXNuhb7ewbCST1GMzlZY7FwkKuOb8T0ep4UJ1HvOyqxh36PaP2+6md3J
foSqaXzGEeapDb0EtHm3HbtXcHuMkBqlWA5UEeR6ds9FSpEmXuKTfqL4RMKshuFE
3iQToAPPTPcc810rzciXratenqWPNIE6gh9przY/YxAosdQqjPcO8jZKq6mAaLvJ
efdVISJbq7N8CZbwdHnFv5b1lgv9wQlj3q5oVbQcAl9Wfe+6tSycr9K+8YHSyiz8
6DiJdF7i9D0Lh+ilhV2WUcfd4xMB5yKlMDDVqlaOStRb0C2PHzH/eZs6oJZ9of5M
D1U6cmUPzHE03ctfWzFLmqdLk75000WfjROFf7fIAtz6lRzGy/TJOsK1emIY0V39
V5FZVwwWHMH/lkNk/x+IGjfM8bk1XS+NKonPx+onjSN5Fx520AdSjTa69uz19VLY
CdLM3mXP76lj0RI9kGnXGN5xe5TEBw1hVb26unB8Y38pugn058vxInims0YWLmoD
8oC/NlgNaCq4IJIkeDrlH5dQBvMC+mVDQ4UfZ7KRztgI0De6syD4K3nmgqyNH02c
DxIzJmCs2Qo3IK7qub9nKCwPNxvUvICJRAnlVolKLPc5ToMIaAAy45uClxinUKC6
BzkvtqYBFZ5aOZw2S40oUmKXZu6nCe/nYK7BG1KmW+V+cibs0fGlpAMedMMXC3cG
zHXQmKz75dgvckUShk5xxVCrRTMEcQTb16NLq+oqiTufA6gkEeoU1dYfO4Tx7Poc
BqjYAbNL/JYg73NcDn4KwoqPFQ72dPc7mop9HGKBl27CCDHaiAV4HjbkZxZ6o6MM
5fx4tgbp3OXydPmg0TYkdEMZkO3XaCVysUao56HKAfgK5GjBhk0v5YkmVW8YDTmf
qEnLuRz/hF2clDSOSO7uL8TERCEHk4bG4vFxfaLc8vcECpNelVbFNmvv4vfNmxh1
muc8NsqgqzBpskWeMou567Kh2qz/n83ZVExEx5IysoAaQ+5l3z7itoEjMD1VH3mB
kSrI2KkTelhOaLjvbeRnRKVSlKbJOybxwp3Izdb7UdES30ntcnq/wFXlz9VcR79u
cdv6cegTHwggGHSX+4dDo0psXerc5xC/Nwek1+C6Z3hUua1fYn/1WH9708Z5QC9R
4kNgcXFTllRfF1VbJ7gvDeyiPGDQUPj++kBIEMYQFuXpi32Ywl8UgBCdPzal5k8i
1J2NzO8SOwrTmzoXnlaZ7FcFqMiT+1TZawpWs1IvAYpLpAAXUEbeuM3zboYWpHm8
o2RTkx3WvcW9L+RVa6C1YFo/H6B8yQOBxMum2DOFN5RJdW7KLqKtQgGNltxPbFFZ
mXBmiodDO5Zsy4dmQRPHd2k5EJmeXsaxU1Jv8BZbz3AjVDuMIREhg9F+jENpUd6c
psdi6wa/gX3TYGkOLjVOgeWdafLghvqlsGgs2xa6Bm4dV4CUC5uDbfdNik6mRPkJ
Dw/DUfDphAWs7KZflS4ygcOBpL2YpvJ7wzF5mq1o9xAL7LHpFIqoQzJgXuxFc4DJ
tqJ2MDOu3GWjNpZkXzj8NaB/AkyoUOu2ANdMXCxeczSPwztHvQwu/KhODO4eMnov
rjXhzZgeJq48SaOVEX6v3p2Hu24tWy26ydp9VeRcf5nkQ85Wg5e7IbJq+odiX20b
i6BpeQlfmcUVFh/Kh2polJ8hiQFgKE/c3Cp2H2AztQtq3fDT2ajh6UsFvBhEvmtL
s17PfVnDmmB39pIm7HevvTZxHxBZlYug2ImvaDyzIGprnYJuPUkEeiG33ptU7/pw
CehNcqTYlcqXsmim9tFC6BkKCwwXABH4EXYTcNbPV0jJs7tJ2MSnv/bOItR3iF+k
9ar0uUlq+vYnf6BG8t8LRdzH2y/RYzfrh041f5KfJYbwDz33eWjp0KVtR0HgV81c
9N5/6K95cf2akR1g1QaOdLaoHJl0X+6V53GCCjx0WD7in+6tV1m9x0/ghTCiizaw
Vv+qeGoLQBPCpKhGn9467Ektrt6JFTs53L86zSsqMm1/HdA8/HTFht6B6q9rw8LC
TTbbCWkfWkk8zK3sOy69z1psqngzOwXW7tVu+N4/hTIAs94akKp0K8ilwjEUAxPN
NnX0OrkaqQVib3Usqc+97HV/wnF6eJ5yhhrGDnd3+buEKhHmvLZFbtq97b3SyHHu
CtAJgRiquOr0s25vRFKWoVL11auNCcBTfehhcRmWzLOxzl/j3t80ZeRC9LxDJPAe
a4L33z2jBp2GrC0RDW0Hh1zNgPgesy1bOUFO19M80a4SXnmYMTETFV4rPq/p2IRK
gGQvf9mvd0ajELiv7RUP6XTHxlGqKWsMKxWHT5wAmW0CKet8A3z1M9TAicqrZBH9
Z+qCCnqTCYUrd7q3IQxZ0t4Fe6W1XAqdFmZk8CwHY+U1IMbfMFIPAUJIB9DKWDrW
oIzU0+/3uPpDAXzslDLItm1cJXkvVz7QeNvvepPNDo7vZSPmy6Jy72xJJmjlhRUY
nDTHHf+vIWKX0wJud/BvdB7X2RBz8SOeoq2WYeu6Ra3Y+1pzM/n5D2F8pUe+QNzX
iNTRq5TEsX8oNuwdcxY5fIYtDN74eYt3Qcms1vSTLydiRyR2ZguxEOLHxM0t3hEi
z/tqv1hYR/8iFW8wcaJM4w6n253h6DZGEITnUAVoZWLTi4j5mUuRM+r8e222p6DE
NZrRl0stj/kNT3oZuKePHgqQ1zAMIshRIvS2cF4ZS7PFJMUk5Y0bW5mpj2/FM4kT
1iL/3plgKtEYnerfQ/d86vp32zFYVfuafJDnK3jT+aZmCsaZfG2ouL2+MeNxOiki
/Py/4qtNKMLSeyyd/e77nUtS/34XG4K7wwH7S4CW+g3MvDu0Cq5V9YT3dxigzaQC
SFAUGYdqoCCNEiOF8CQc3XeXwQJ8AColwcgexlfrX9CiIQ0WwCpYsSMSB/Exc8rw
IbrAUPvhCjo5H0yldpTPbBopuHsae3yzUhD/GvAnUouUuwyXiZ+GNou+/kTtEsg7
MfadMVoN+VVbib6xJ1mKGWfgjd9ay+5MF3oEcdz9ymWUtLxDrxMH3QnK3W2X44/U
D5dOYkt2Zzpb/Lbrwf/NyZAUI5cj90aj9KzoJ6pR2aVX1Z+CLImz5ZLen6fMBS5Y
nLAzVsNDSlQJ8EnZFk9sXIg0j1Cl0s/aEt7F56bCezhRtz+JUyReERTqgDKZ3cYu
0kOGKAwKyiy1zJF0qsI9vDh6QwMHD2FQg2jvsopGtBmc1PiCO0edjZJRcXkqW1yM
jGRIuN0oI4zoCl24EAiGV8dgYhIevxngYPy/tqeGl0crj2yPl2YKF+oOBa9d3XQG
SKWJlj+BxyFne9gYTsGsPEf5aTNQmW6krqOBBoIZ2rwI9Xds5tZjxAqTfy10sEBE
NNSkGqzVC3Z3aVJFsHgDhNNKISPSvE4phmWzfmyUz7gbVgHXTQ1uRMoZHCQ1h9os
7GB7fgDitFZlICZKmvgH4rqrCGPM/0KlMPg7mCZ/CLaD87DFT6ZIQtjODe2n/EL4
oYq+B5B6UzXXSKJSS7r7buDp70Jz8iyHoo2aK5qSwMb+7woIjlO/zq7FWWcHvjgW
kRTiyZlF/flIhQ900ZEGRxcqZlEhu13/ngMHogycjrFukioRO1jtgmzsdzCjYpaI
Ot6oUyyr2CChEc1lLsInT6lMc13cAerSXbZskMV1vCDy6IN6CE6h1YsV1M9Mlfcx
S59gQ8Z/eUsAspUrkFYf9YYn+H2ScXMv1EDYydMocHB6BvtvYNIyVBUZjJ/ih/7i
Md8FUqgMqTDT9L+o12W1KL5m3fSwNEDc9JiIhv6i2LrdVchLRm7F/NiPd85T20J8
xaxzHhwM7IMq4LKPXWQ5EDkxnOok1+viEqukCTfAGZNmeq4lzq5Vx1Jih+YL+qKC
h/KgwIkg3FK3Fecz3oGmC2K8r5HH0RurWz8p0kYMvTOEXLPRl7ndIbutJdnUbEhY
DPNeK6HuvlEi+o2f8iAd6aIHi4tXRv0B30x1U8prlJLh4EcdGR5JGXVvPYGAXtMS
0qevVrwq00zeGOKBp1LvQD/uInRFheHT2Jm5U5DnYmcoz5XHFsqe0xv4nVr6qFz8
FOSJasAQjBdGtYuoExJlCmAImX/RPdbu/Nvywj2pCLaCVruQOKn6HfTYMKq5PNBx
1lucchvSOXIMYUxr5et8XU1hlLri2jcMJr3TqDO2IWhiL71otQCo8m2SucSjyu4s
PpntLtNo2Dt3smk3NBxm/bt38Q3IQeA9rdLu/IRere1AHCbnSTHddnnZToQI/J4+
TGlzi5h610bQFCwwDcIUrlTHebkq/GIHFwTWg5rI9Pqw8AHcncTFJPa1Ee1P5UHQ
bpbv69lM4QPkrFzZFXP3dabszzmMR01U11P3SV+KFI45BNKq8rnIIrlnyXCdu71K
rb2S8XOpKg7iziWo5uBXUlKTvoEnhhBn0l67N2bh/ZzSmDZzo2yZiB+wiR+/zQdn
OHDWu46lc/zDG7mzI8OBgivYnqgdp0l7bhu082BWTsBLuEaxpPzVu0/Be9RKOo5E
6/zmQYN0S+ToIpCMXpJ9RIXbGAoPbJvIQIGiklUcSYdNG2mha7t+Cb/bMZMOo04T
CphUMN3uFyPSbRW+LjbylEWRXzwongmbEhx/iKNnDVmTJgV0Z+8toJoGxXQbgrZ6
tAUSFj9LZXoMhDLTt4zLq9An6xZTkdkdQYiN69QeEBFNvTCMgZEV93IgPJbbd2mu
LQujYuytv4E9Wt8P/9RQb+ZmfiCpGJUfmg5lue1PCrAOcTzROwz1D6BcXiF04nRk
2iLwn8zhP2GV4D+rYmG79dFltnqwVZAC8ASaXzxYtp+Ka1P90d14/lDPtkhz8uCJ
64bnNcwVQTeQ63VcUbRUNOBJJAjywIt+lSeduBoY/+gIpcYfICh3kimHUgco+i4P
DDMV3uUBbatNf+9TLh0yOkaRMzJ2pBln3fI9LYPN7oYWp+TPCodHDNdAKVlJchuV
/ymHOSPwCnlC3V7ClzjYN/m2+Uk66pdmO+sbw7tnm79ACQpA9YmgenYNoVyMhy4Y
LYctoyupioEi8ipVF85igacILIJzwebOJVwjfUrGxAyuSOh9Dk3IojUzn4x+qJj2
8BoE+JHk6oONr0bsSYrScS9eMEKl0k7Zg9sRRjXgGhgalJMay2EstdUwrpHDWsdG
lkbeUjOXma2NNZ/VgpIP/Y8XXFSledWKWqSyhd1MPLa/dHSgtjCDFvtGmPf+LRJE
f0ndCFivg5Pz9/CrCyE8wScwI+FpJgvYOBm4UEqthvsqpNAET+kYiFQqdYx49bZK
49mElL4kwp6g18yd43QJRfMHggv2XfVdAd3OX2mPwE4x1n/Rb7L2LXNIWjMVTzEY
Q6DiCc4Q3GhmDTOnHv3li4l602d/Kt3LCCTe7i+Td4zoO9qJNj5PPnrnb4uMjCbU
bT9Wx2jNUA6mxaOLTBDeiU8dZFnNkCOuMKxcCERm9+r6nRwymiQXw8F7a1KYIpQr
YKuA78U0mags81Za5s3fUk6UhwoffB7BEAk62k51HWgBQEhNonAZPVTw8OPQXIqs
1m585IqFze1v988zmLJ/5A==
`protect END_PROTECTED
