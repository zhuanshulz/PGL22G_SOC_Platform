`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FQV+i+UJ1ns6/88iNqH2C4pOBfL7wJQegj7zLielpvcwMOrjto7aXfrqtPcVzOFg
I70hAdkI/lL5zc+0JH/tVG7Se9qHQNqlcWaJETG9Fnl/Wxitm1sut0zrpGZrXww/
oa+kLmyRwsuGptXUO3bWVzPmS9KzNZfh6yoCdukwdftpKM/iGybQRbZVafhW3vQ5
K47+LR6gTolpbKQEHsmr11srcNJgQoWfkP8F4l4uHXqs7eVpNy9GMzdXGBEFaOjP
yLumSkpS+QtWh5qGrI8s1P12Nj/h6IudhXePQ1KmniaCDxuiUTFs+58mD4++SZWq
ry+c0CiI+oJz6kFJJu77eP2+A75gJNT60dfMTsP1Q/sVWvSgaDhckdCVg5tb6equ
URdS6Wf7/qMPlM9bUnu0+IJ8XqUEDl1mUCoothojAbra/p5TX6m6nzCcqTuGfQVL
5Ks4xmU8oQzk4SwX42779wju7OJcZOIlYPbKNhylnaLhv5kiOqCqqrppkDrNZYdW
mJPGh4TSgIr51KwhwGKPI5C0Rva42Q8xe9ajlRXguBuXzRc8mXthpwRCQPBwMbe6
HWoV8ej/5NQDFihfKxL57hpmZLBRyleK/9SLB+IcLTimlou6T4h2xIBvs3eN/X1z
DxtJ70iFM3IR27V6xwyvnONMRGh7BgCNxKbLpzEk0QQcRu656T+BvRLp5KPQmbNM
pVC0y6w5h99pCyVL0ai95YcDiwuwriVmGviK8rishSGNyFhOjI5g29aIVWhf/KxV
tRrULTPXCo5y9Yq7ri8xEjih9ucE7UpzvOCQukGs4CdktZ677xJ8gOJTCTLtdPHt
YqthINpzuAb4+vIsVT2oxHDXEm02PBBhGtBFH3q1RGpysU2tkjQo8lim6UV8MddL
uFWjMbxBOvWvVWyn7acMSEJ8rYmH4v4H24e9IZT1liwbNC6sW5xaQ4DTTOICdjPb
CKV+LXy/xcIAUrXQa1Q0zA2X2HfmIM80dECQ5Ej//2Z1jg06rL0UjltPcg5kZAfp
a3Lks8bm7L1iNdfiN9cULKZcDwm6BrT0LxdF+kaULVLYT5EbODlenOs5FMV4Qhw5
VsRkw2GpjZHoKXDlfcJniZULlAKuvoyfu9OY7XVw4JSsFMqG+NODiiWcMQI9x6fI
f1LDA4Z2TOvvlWq1OVV7hiivIBrkR3I5p2fEkjBoceqQNC9jYxwGk3RzPmLlAdla
FHjxu+VZJz2ckY18wMA32pq0ekFe6PWUxkmxuOB8zq76Wkd98jZ8JpUVuSJLJ/ot
n58w9Y2s4FWfcXPrN2+HXglF5NAhsmWm+6Hy6GbNrS/ESZyGa6kHSZZmQkmmkZUU
2XI4soP1DMpBdOCGDcJyHpity39hH7nk4apT5B3e3wzfNnyDmpy+A84Pr7VXENXr
afZM4+u3YIK++khd56SksPLatixAz5Y2WrwD6mlLB/fgtgE2FQqmvRxJoNd3SxQx
TqbIAgGDkhEDFYNpPdZ8GA==
`protect END_PROTECTED
