`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mHtrpjoyU84AEkp5Kx3JVMGWRfQfa7+9rX1/Ry8w+bL9W/lGWwsXudEonwMP8cyt
EOawlYGvwTVd5sRgKbE/fWWWQaYI8a5/EBC/9CY7Gulb9XIrps8UOGqfo0K/5m1t
tN6Vp7zB1kFOYFuW0kLDsIyS5TxuU2ST+Fr/gZYfetateMWJ+WGl+5w82xv0+sYh
ZFHNv3eoUq6Mx4zW+xQiZLQDzv5qlOf6dKenARv4RLEYEo1hylxcEs5UlAUZBKQa
fmwsWheWH5Ynzq4UophQ8suzbsqnYhRbtRF4w7ynxw4JP0sOLUcLSKWOs9r4T3WQ
UuClUD3FNECQFcZ7noZfi8MwfxGN+52rXpJgQCd71qzJcwWdvDW0Jta3U7/8uayC
BTgRPe0ztiiRL2CgtXed3Gok2REO9OonzEKgE6QOF/7xTwxtLEEcuf73QvYxq/iQ
Ec0WnLMqUn/ZcnbSLjUrIntpN3kEEj4oprZwEb/qVKJ2CFH5mRcC/RbQPy/PO5zj
zbJrodCK/IyPxqZN2U22+2MJCd+m9N4tPLq05N07BcHPAMkXi1BEkClAwQug+wW3
ovpht2jrc2XMtGzWP0Xlx4PkF8QUIg3vjKMVhC9IwD0gfUtpqXERkZw6YJ1OBMij
A5lKmVyyUSUayACHCAT5URUjYoyr2aZLLLpGqbhVMQPqteT1Z0APId8rcXbVv1w8
wNcSLEAicWDrFG+qOphSntfgkWA4BQOM1fwHXwLUlm9HNd2ltfLBMnJoAVYS5TPb
nRfpfVHYVhBN6uxPW5L3EPKl9NUbpa1Hyka3cZUWMllNs51RU/lgsXdDwRUOThQ4
2jVPtddvyZTVkhg71/razRBRryX4sCJI89V/36Ni5izO5+qHEnSfvP5/4xclFSY6
AYP75QuEqNE393pdOX24tNcxM33pFQy2/akd5Ih/5PQeAw7+8i/DmqH+yzv/XuS9
t6cGRjJ53Ka4TPl3nzSPVj3+iTo3jcpSW/nIjTYiKvuOJuMm+vWRUUbOg47AggtE
flqXneyxzmdIu80GwflFnA==
`protect END_PROTECTED
