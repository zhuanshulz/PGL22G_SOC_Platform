`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+ON8HtriJNR227sIXqGZfsvypMvzdanQHU/QUzV+BZ+QcCN5HXkSrv883GD+/S3C
Sa7lnHejiiWecqB7aUVTs8UTZFAnV8VeuntZ7qKNKiklrtaooBEwAZW8tbzNq+OO
GfiBPWUlZ+y21lKd0XuTsqka856lsyIhWmLT30nRiT3RUZKLoqt/t2cgZGRck6hy
RiQ+P5cJMOstYU/QPnsG/ByKbpDkDgSWd9Uqp1cWtnj/b2WzkrBGk6wSDgoU7NoO
N3zPfRCGsK4ik4g67JzzQNGfVxnIi6gu+h+ICQlB+hUO80OxNvmlbNy+jWFxHjzP
PIP/SClzjO7VO5x7XUGMA7JQcCl+HO2NiQ4jL/Qp+x6OUSVyNWnWctdIkFYDCND5
6ZvbUcZiwc1lW4U10DdXrKi7b12P1jfnN/O6xGXxUrfOP4LpF1kPmlQc+8s8XS5W
RG48C5oGZUby4ExFtAChjkBE3Pc6t6TmbTzAU1KRwlhyjgT7h3yDuQmecMmWAUZ2
9dliHUX+t7YpAb3i3RQ5Sm4y/pU3lRCjtmiBS1FNPuiuqGl3OWxNw4PT3Pl+7Qdm
kp0o2cM7djaLpM5xBWtyNcZXX+yZTG/Tks3L/T3V/vFgjU72yOC7fxqyfeVCcvHy
pzgK6v5CgQa6nANcRGdnxuiq1PhgHoHndk1eo5mL+hSA1OHTDfsTekV4Tj60O4pr
dHF5m7FWsFXoul1NQlgx/2jmalA24gdLY3mFhJSof4DASjlX3wfTzg1FIR3X7WnH
pDQhIkFprHKsEsOZLUot5pGszvV0/C4o4Rk2se2JfX9+yX5WJGjg4DmgTs9RC6W3
XY0PoBoSb48RGb3NfJLKzA33rE5ugGSlfqSa+BnQyqcuDEGMIHCiDOUqrnrz8jcM
Z1OeOoANfOuqI26rYRgm2HrZYa3sDBt8tFd9lVWdmmMRff+zTBEldMpfJQN7o8Gj
F2cauyXBiQB1BWUCpl8YesuO2WzivxDdGC3uuuSu0G8=
`protect END_PROTECTED
