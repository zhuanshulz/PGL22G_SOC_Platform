`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GUq67pQ3xlAD6A/qIaZQ8PLoPKAKbAL80vD1ZrVrCYlTs85puyrWBPrTU19ONLtJ
cv9IHN0vjcP4LvNA3jgAZLgVxQobb+zBsPPQSGCPfJpPTg7efeSENrtjow0PMc7c
0BqKjb7aHm0Tkr7W/C8qYoL6RHz3dMi6AM/xMw+5bmsS8uNDIMIPhounjy0g1hsE
N60WTgUEr1Uw+DvBmnTJjMf5mDr9bwkZZ9hGBPgH0Meor090upUWDW6obeKLPspL
urgt2TvtcuGmm4t86JnnjFlvJQ8poiV487NvBKk709e7ZTUDJlf8e/BayBs1KDOu
ZRu/Ya+w8eOg8MKKQsP3Vsf8+43x+BurXHta0HBssHYr+ddhqCe+h/R/Km4OGBtE
AflyJtH227Cq7e5C+mRTU2YI1ML8j23/zqfk5SJbC7bb6/rYFVvz4nS5pIXc51dN
x/t9g5yk125fiqIUpgS+Wq2W0jfNRTyowFXx43gE5E6gr6uniYEzC8Ew9fHOPpln
SG/mgykqBZ6cIcKoXYdKQewxCR0mRA2Dle23cUe0XRyCPzz0Y8kFdrHdT5qFwqDA
sqlQvTgJSl2RJS5j9297oAo2ib0ycz29KXTIdST0bccdg7PqvfRedhealamWQiL4
Gfyey2jhjSMN1DvICTYotog95kTCQsXX2D63+s4j/vqC8aESKUVl3m5ofTVDQxCZ
tNxRqx4mFHWC/bivwW5lkAnaNsU8v6tE3B4iakzNKZ6IYVIrvjT33fgCAvJvoTZu
GLtqgHyqQVckWRv796S/j3emKw2IGg4w9GN5dlmsEb21NPrI/oIA+n0Mq7OIskDt
zp18vylO5hHkwGIWRn1S/dlG6nywvoAogRdadmvWP6WhDIgqr3Z3xdQ7G5SsAkSo
k3qy2YEsrvR9KexUPFBHzfMcC/wH9lWsLgoHtaebjLXjziBvwetpvJgUa+K8j8q4
AgsCtNc51L50pAYXD8ON+7D+wZ83Um//ZuFVZjkZyPDF6xFx1WkDO+PwcRDeTm1f
JfvaF+zdN8rJ/XGTtAkumQCp14dWKqg7KKW2BS+7dw9zRxAba9vIBw3RSBjXEXa6
0oTFXdnFalbxqzC1ad69kHqe816jCeHvWT/Q0VhiRD5/ljUnuAdimhzjRYKBG9nX
tJ77hQt/YmxHlESShuf1WhOA0gGKKpzFByaEwIuNiIeT+YC84KA9bpxDOxbtMyOe
m1NvEXzFGmt0hog00V4eyQz+IBRX2Vm4qkgh0/P9KpLPeIzds8H1CMZSBQygXyhT
2LduRel3hkX/UXvaW8XglC2nkjTQIz6CatCmdm1Fym8b+JzaQAlz76imrFlAqmLV
9pgiV6fo5lk3dqJ+WoHRHPi3HTpo9QPL7SSgptUR8Ev9WfSEZ4ZmyD12SeaqpULy
rZIwVL86JNlw0Ly9xL/vygOEaVxE9bB+pqq5QUXqpGKU6kPwgjVqaNlymtkYopdR
DemZOriFzNWHrMUwKfWGMkuKrJ1vcQuy8h+Yji3896HpbtMfVmbcF64rj2Y66iA4
7G2OSirOApqsLlIRdkX/q3ZDW7X9aaQ4tg+9kqN4Y+7FNJRoH+n+jOeRDIPZj2+M
zYufz9gjeEoKdsvXRZ5Eq0a0WqhegN/plicQVim0xJepMXQ/uxvMqTByWE4AINiD
CgEi659M4ZUGcX0GJDdUBZwtcHur+oszDTJU5fINU7BNx8hBDBm00Yfxp1t8sHnc
rUmyvsM0+1qyWSVZtdXZQtR71Hha/3xDvDfviJkNOb7WzHQNPEtbHi0DXS4aa8aM
njBVmtXoxJfLyzi7uY0BTtttIDMblc5Czw9W6Ty+kSvqainjGi3N/DBwKAu6AXY/
SmRxkGOMnvEM6J/BhNfLME4XW3KX0fj5ZwiL7MDpiyHUtdn9zxskcmbezxrdhA8s
JPy8OeraYXC1EaNt8IGxsQgtwW8hEkOiJetIbTYU0YEQhkOsaaoXOuH80E6vUrG5
vGtftqN/gxoRQ29P9Vw8i5Uea/S0oI/kQVoRoCS+lEYzZez9vUjD5fza0BnvYs8C
YnBeG9TrvRz6/vjHIObyDX0X0gPfye271FHdJ3HM+MNo/7lsvOv9H9ZJBxLNoQmI
tOuXdNyHg72vWkSMv/OGr3Hn6YCbbTMgNHo6hOhlrv1TMuk+n9I4OxoeG7TRLy+/
sfph8xJPSuKgTko86axKyqhTkzi03VqrR/DInw+KRar/3kNBMVQkFlJIFG915svf
MqmnHoEOedeb5bgVSOd45TlTYcuntQxJJYDPQ8JAApC0mfFERGmlnmkHf3I8j9Fv
OzEGAj4nJsnzufIIzIui3mlT2Lz5Gv3nswWbVmdT9GWe40r3Xx1azjGyHwpbKRz0
MM2TcJxDTVprcoUwqgmzBTlcKQSYhdnxR3ps5CVJmBPFJ/+YzoVMFT94yuaOLEf3
KXPnNL1wgpd/Y7zM5Thu36GeDgJ/WUkKQGusO/hbRleZVmlhnc1lWcbj+NzVCje1
I/tmNv07Z6/VXankl/NvTvTy2r2KfGoHexdwl5eFH3XEHoRpbBWFClxZ6FxVtBas
WpYyQfdmr9P5aGqbZ2ykn92ilqFRrOeZ9hNT79eg2YAfHVgj7lMW6bdC9W2wxpyE
zOUw8G43ho7yXJO2N5nTSC8UkOZMK1dj9zsXBDVaYBpxCno3se/B9ZTDBn4bVk8p
F7rI6zyRcY3OrHl4XxXYQ/L67eveG5TmNZ14nSKEyMZivfYa957QFQhxXOg443Ws
8yTJKxtea+9LitEAWkpK+gr4IW8ZydbAA/21TG5czRLGyxkFeSn+TX6UNxGn+bdB
k+n0TwZaZ/SJ+/Tx1587vu4PTHB9hBBVRV4ve3VXXtvSKAkPglwyWhwG+iRp+A1j
vNrEDydZOiiNQksJHo5Z6Avg21U0IoGrQAIm8sfFb3quJ2+xn4oKK4793DqFfUgB
LEHLLhlu3Z3QebVGo+RMuCWbthNfz4EGjpcVfb+Z+vAGRdrBKPh5EHVbV1oqDull
VtVW2Zv8FwbCjuQf3qizm74CZ7b0p0OEYzzJWe6WkPkxTg5yCCCze3mc+FaLKKRN
cwSspStjMqbsCTRpDWnJ1NqBoNftQjQx6bhmv9791kp0/zKfzi7PHLjlxuiAl92K
zZiUETFksLyhqdtZyIueA18Q1JfoFjw7g4/Z/5wlrLXkgf+yhIVbtSMicP67eAR7
AEXG8a9zcq7P9N7v6DGK6KJwVeHfBpuk+UK4Zr3kKA5WVf6bt5sdcHoZdGJeZcRe
+tqbZnsHaVXKG9ET3FpoNy+xi6fuj3eU28gyQtB6i+M06YMcaoULzsLq/rn53kjp
WgNm71uyVHPMWzKdPMg7EeQuvNfdrPryD/VCvyFj0b+eniTKpsEMYA1QtesRYOP0
odq4jKXe9u0JzD6SF5bvm2rjAMw+wCDOM7nh2sXW5j/j5eItAYs2z0b/FPo1S8xS
Lb5ovn3uNrGTS5bkv6VfnW7RlRgKYlBpOhfJT9Vq6o5hgXNZycI6KP3sJNFqbT2M
EGpKzZwALnJhVIQ9AAazMpWGkBXlY4s5ZmEqWPgaSVLOaNblTIVhLaheEF5Qhzq+
C6JVYboCk7VdoFRDVWgbEXg+tFrVfm6FZ5hvNMBllsBuwXBqRixbptIa1mYT1u8x
8kdxxInFArQqZnj7CrGsRnaAP5wCluxSn/qJbJ8/iZR4Y/zmBFIZS+anWvZeY4WK
CxYs/9eaZHMKfHi0PYQGd8YlMx6kCVDQhyV02PUdCBmmOaFil3JFIAiDwpq2/uCe
Da+a1kONaibTjZQTdaPopt8KGCIyUw9L5Dnsaa7KYsUtiWybhJXF3sJFXbtRl9UY
Yre+7JVKCp5Eg0S+0xnTvnIgHzOaQN0rFkTDLam5HMopazkxUDqJlIhDdyxOK+WP
k7K/KovNhPxBOJXGGJ1vKfLT2+Ckz/zkMyjcnWf4oDHZWKimAyoGlH7UhIyW4W01
/MbROMwgTBeRMJ2WdMXlM/E5HT7DlXfx7CBzrGLcZWUu4cophR+vfV3iyGNHJsOJ
ZzfwwRBmcI1goGzff/dpaCxhN6kiiI9P/2fqp2iHMiKNtkPYhsFrzzTdWrnDpYZE
ZOwK9zXabW6MkfxYmryPFv0kpFNv0HmNK5c2FsjLwRENGZcEzbHyB/NhyUgmTuPN
gKeVD5dTTUg1HKtz6xzIl/mxzFNyeLyjjOp1cdD3TCFSKrStkeqgjmUdJMzT60Yh
Grwvq/djC37XsH3igPqUA49U+AtpxEln6JPnjmxrup9OtbYwqfjOUTt/ugaRdZIR
LRwITIIJF+Okltn7hZ65ZHhbShimXIoH7/R1vjnSvjVEhcncYONz1WN9UhBBjI9n
noZqBobZwZY+Pm9HVvvk4nsixGOWiXMAOSgGIfiKJP5EBewPgXzmbLWpPPx8o69p
qxfe/O3qfYtSQAvmiD+Gq3fXn2TTyvcByPZ/1Y1A/uenwCsuIBXVGvzq5oqlyxpo
xlbRqf82VzdEBML2R5eolgpCaMIDWJnrUw0f85CAJ08POdSXMxxHAVFEcA5H5h55
LCDbQVkPGAZe2s6BoVymAFuS3ZnT3UlLOclFtM4LdmcOLitjkRkap67BoYooBhlz
3jtJkflG+PXqBzxPxbhHno4+xOsg3c3fZ/ri/xUuS39nUkWa8yjFEODKPiuB7Olh
Ayn1Nj3aBBQTyrgyu35QFV/maIqsXUAenG+tXHYMy4buUwyavGE0uekowPXDWRy3
/Qd54gQRR+BtaMtth565bm5EeLzhcWPR4XSANWt7AFig2FhHvN31ce7tWu4AVNkn
6ojdSIyMRPq+FqIJfyUhn2SRBtxgQmI8k/ELz62e/M3UPea7VAEvTnRpGgQ3nGNI
625h7vgELicEK7MPTqNjVxo8OCeBlpbulgxOvpVs+tJMRuHvpMVfKiYrSDzI3xol
uhz7O11jvGj+KO3Op4fVCm2946z+DAGcFJoWpuHpaQpSf2UOdZC1XI2aLGAQx68+
bybJu1RuhOTg5M2YdVCozvBLE/6PaBjamI+SGB4iyQdKLj90/PjApmur8TnSY4B7
Gx4FJTyH+bWn6y9ByTu6e5n1ZKkSsAy2Is2Kooq1j+26w+ryg01JaSIg8mrJvbb/
fgdGwE3ciG1Az7l1af0SVji2nUCguPGSK27Ami3gzz+zImTJApPgBOqgh0GtCDlq
LYoDtvmUExnm7QfBMP4yOKaliRL6qAD0m3Ci1d/EHjJuuT8N4NidJ03XCu3tP936
b9wjfi1cYtb1cOE9o3hiMZX/ZOeDEdc+DtXjHgxZTtRgo8Wa/TZb7nMpC4BUIPjW
GCFz/difxVt5z+fDA6UMziqYxLmuD1uojuVxBQm+qQwMGJg86XnrX88JGd0wfkDt
594suEb7iz8fN9ZWRTGh/ZWuhduOoMS+bJKYAbxs1NOUuxDIA1ghVx2ly7Q6Inkb
LgzeRMPDAUREk11hlLKhV3zO58O9OFcVaszFzDe8m92YK6rpHP3QicIZIjjgBIxt
/8CiACeN4ms0FMLcUuzjt6FbiK4rPV9zz9Byz9GhF2Mx+13hbLlNfxA2SNIqc6Ou
ArHvHskR9cWsRO3q9uL85ePuVvOl7UWOkDtxqP4QUWv6Q1oZ3OMR5K1kkoN9piaE
dstVfKczlVDSL5bUjv1GHxrc23oRx8iM5msLsj2vNuYlcyx+yxW7MuW4/xJZmQPo
9KFS1WdVoLYF7ASzr2+dOb3VsPwtkbCGJ5VaVt2b2j3Q9gJUn3bS+2rVp0weO+NJ
t3M3cHDWGXi588UMXvLtOuI9QzOmpbGVLCwhdBkiIyAIF0RfNlIBKDLmasvYfAiv
CnodgfVeLb21V709WSkqxHtInzHnmOVDwdsLZY+4Vj2RLNaaJX8DWJinIhiJas0b
t3+JnNYM/AZMBNqWbBr0V2w04+OIL2mjwGGfRC4Gu6D4UBSstSSU5t/OdR6jslpM
hvPwZdYl4J5eWxeavwQ+7vlSpR26HZSP3MfF/K6s8WClNl50eBZ6qLt4QECfLcNA
mAT38jxirl8IdtkZcWbO7UsuFvZ/ws3V7iGeM2ermaU28jTTCw0mySTwmsU6EuBR
2iM93WXpZK7GUvWXQxt6bAk1HkrQ49zoatGbrSbODiocZHBBf8HmXe6ORGK+xL5B
2Z2cLvi+/s7SFommBjjc4DuHmm5UXNFs7vu1V+nZIaEzpzCdjUxVT92is10mPC66
oLt1AAurVP7GisMpn6QgBbDRefKaGeyRqjncOfJwFjKH88//5hHqqqIRmNcjdbe6
EdVelnnnWQVhLlE3OVAFDn4/99J4pOETANildNsLEvEOl5H+E9kMOPVO/fVjG7Uv
M7nagx6yPtTiLK4GZZmNcM5LSaSsw7ocQpM0wFST7lcsWq2vjkWHUoxL+QofYIgN
3YlCzWfPAsAbbb41q1nc0IhYFjSvAyMlvZPOt24Cf6ZQLF7HGY78xe/m8kwkCNo5
Nsi10XeeMxZYu1r1lzdjha+CbdVP4NGu3INKLFiPT2khYNq22tDI9+7HCoxSwyEK
BqEch6Mg9+iKHzY/5lKGuWgUNoxvkWyBteqQZ0YXHaGarOJKkwFDerm+y5HErbbE
UHRBbQD8VdB4OQoPB5iqLi+9aZoBeSVUYg4iQXKqpq+SW7wJ8saI8xMt8yCsR46z
/mx+hv7sBh+tLOnLsRjBDLlaHev1LyEtzRW/tOgYsMUCw6Q+ovjWW7Tg4agO2xMl
SEg0ahkQRyqj9zR4/QhSUZZcd8uRdcdK8ZLxJQCGDYYIMWQYvVNai6dHR/0R3GDn
HffSan1giwAm/44dHEcGRGfdNPmaj1W6OmvCMUVjwqeZHA+Dy+b2a70hl2rE4p5W
YGmMqYat6kR9BHbM1S2URsyoIcbe0ZEikUfPdM473MsHd6FfaRePYb1a23FAMNwR
6Zzili17bXV2gtD34fVcajRnpUdzBaR2T7yi/VgIb7pn2q7R8gdBN+WRCKJYqkZH
gVqpwY8stFf8WDC+GPxEmA8CSp1vfNUkWfqU2iV2iQ9S2Y+xaWE0jhwDnRpMc+WT
XNrpMgQz+SdQ4s6EZ1v8V9YUWGTi1gSzpvvI4ptEoSiX1fEGdoYqIotqhvJwLowe
/SroahGycl3lE1KnahuRJhahrObI8jdv7GjZwuO+P1Gb7hiXKtTI3fV9FgTARDME
lnmXyOqUBIkStlbynagUi70W+UcqfjT7PwRpm3ChkUntpw/CgERKW/KPnd4RzVx5
Ehg0eoSuFgkFhmV0va06o0lz9G4sD0b0qjGeUmDhbHNAJBxN774XpOOhqPwIPfQd
/xORyErZPICdJFBtR/KGtkwP2HXtes3DOOpkiEAeNOWzfmJVdESff//ZbARnabSV
V1vAFtY1cwzArQjBLXMYBMXRBAAzW8Kixmjpav6boufRLIXg45YvIae+nlB4/9ND
K3EVTmgCvF0RJthXoUaIKvCdZGEZ5mTKgA5tNbOHo3NPw9qgRu9CWi0WnR3jnfeU
v54HO+ukUpwSS2tz2UE8+PZQ3nttZwcVUamP/GFGZNlkZhfO82Fe1vWMrj6q3VRp
/Zzt13xgWp/ixTC5CZPaPlcqxwd/X1HDtBnhvDaYdiAEZeeNrFSjCfmRgS1zRGEg
qDgFW+pJWD3f2qzKqBwb0xcjfF8fRwkiE+HTPsADraMlhPIkDS3vdGOjhd8+vcSK
aHdld+YH6Wo0u5kYJirIBOO/+7FkdyaL7S67ZawED31MORiS9pEOvY+ziN8ekMEr
Qm/Qkg+MYycSyRCc6VqoInBnN3Wgq11Ib82Tgw3AVvHKmxgLAv9YO0V8nGEl/AGi
Ej/ul+tGF8WI3tWDmjpXWDhFCvpkLI7jGifclpdje7X7hUt7W7u4NyOiTefqzCeS
7BPRGeFyqBsZhnDLW73sgZxuSh/uSNlhpQ/GysbMKiuFuT6nzCN2az4vibYF1iBV
UaSrjb9N2GCv13XK4KFgJX2LEUfauKf3zydLcAB0oF98+oFvActwFwZxE5R0rp6d
skvc+64FcJFp/Uf11bKvUALGfxtvTOEJUUD4tv1CD8Rufa9KOangpnwsNOyb/2ww
nID7fY1fL4M0lf+h60iBcnUdlElhxXq3Em9zquWmOJkl3WX1gTVsXe8wGFtjnopK
jlFVNwIWn6QehvjfTOiUulvvlAfSjAHZ5zGP8Ztl56dz1cRyehEBzIdxxiv1VxQm
OdG+f2XliKC09b7Xhs7+KY3lrZz2Eh3qra7Qd1Fi5JgJZNmlonX/OBYNTOsbcEB9
onvU75XkRJL0pPYfAja07VNWLBmFl+BeqFN05U+VC4yyG3R/ENIi0BhxsUbfP8gm
4tzlvY4gT+HkO99GewheRrU3Nb2MUiV2pYa1ZZQLsR+ZcZCicHL46i3f1OVjaQr6
eI284x/PlboanXrRWg5bQPHVYhuYeE43h06fmNgqZjndDcpqm/HfzO8i8bNXlhnu
87IIzr4c8V88KVKWAkzyxo+3FcyJ8bwSw6Uua56dzj7bOwKtEgknDiWS6r8YXvG2
JanL4ys//0n1AGtJne8aJHfeJaJPhxWXCvOorq2g5M9PV0grOh82beVSWTe3LGRX
YRE3kjFpJgCcsa/Ast0iUuQB8lV5BryUHjgsiBMTr4YCS81eiRZOJtc2pbhOoo2b
BDgjnRlPiAyvvClkR1v1N4bSIKw4Ck3C8LLgvQ3H6Q4+HwTSvw7L65aHRzfR2uXl
Hs4K6d1N+mx2PpaDb/GYUSEtO6MGVmGiJuA9XP0BvB35zeW0zSlOvqVnVSI6FVT4
0pYs2tERVN9woLAsmTc1cwRfrQpcGrw/MsCjWJrUx6BNpKIeLTCYj5mNIlGEEc9K
4P9QA45vwwPCpyQqcOp62XwUsEf69r0vn6AOhMrQR8g7eiAD+K2vv8JgoLInaApm
c7REe0ML87Ca9+/jX5BJxb+UaLkCMiL5MgLNJ7+5uCJ18nTbhhVHfqF0Mn7VXOR0
SIrbNEXAXcTT/UUBjCAMyk8odz8jL4fkBoXl+T77/0CDpZrkww8Y7aNrwQu4uOdP
Ok9tRHUDSUnOGnn0OCSLKPcdvDiQSM2bHLrKO4bPVfap37yGdTcxms0s4Ptd1Cur
5CG6en37sXQFYzHvVxPseyC5zqywUL/qlGPRj29s2Y51qCPSNIAF70nUfuXiIHAx
TvQbZh4SQdYZcVtn1AgEkCFgWZofwWWnoHQzIouOjXSRPMs7Wi0T16ECMmDiIeCL
d8hipApBZVQIUip/BkGa/2OazSQYXFu/S6k7t0eYAafHSNC0eXDDYSoAmZkQM//3
acldtkvQGI5CCQZG+l8WeEQFIBX7FjKQt5Xc+hcYwbuUB/YSrRQ1vgu3agsOCruV
m82Ddz/ZAJDdDRZu6jyWRw3gLvglTXSY0ip10iXIKybO8XioHct8TcpDzH5/UJr4
bPAA8CNNZ/hqcZ8VGxDKJwC+gj5KTrkCpvFAzXPMTXUK8Q9qYplX1rutiW68VqKr
3yBAa5gPN+nPcNrC3OJZ/8lG065iotzZMJVZXZan5/SpYXvNIIXlYJuyNpa0h/1b
9j8Qen1p61AhIx46jgDWDGtQttR5vVIdYaE0EGkYjQO7GPzqfME4Hmb0iVfScUxp
LQpCc/FEgGv/H9gdEF+7rbSmCeSqGmXAU/5s0sts5Uqq+DPblLHZoDP1nJpUND2w
t92Y82zi35c0hzziNwQRnw8QGcJ1GDPRrnngSZ5egIvq7oBoe5f0i7QxunBE8pN2
jeY5IfXIXvljcDORW27Due87BKP8Ox6Fj9L0Ri4igGhNsCB3wNri87fTesj2e5TS
gh0l8mT98nm3f/Ld2P44kjJk/zWYk7/omIbOhc0u1ItV9Oo52y60uC/KYlu/5P70
gRzaVEeUiI+CyNk172O+XkNk5zK4IbDVaf0/ca5WubCMpLQz1ecafWSVR3qi80Xn
TMGDAdO48ok7wviO8FIieg7Yix+vZYu4lV1qao+iAK1vnYXYHhkRq4KLd+6Eufnc
Iemn3Kjv19yvemux1K30/7Ml5D9z6bAWBvfQ4c7M5xZctG9bZDjrUjXdTNdWZo1T
TDzF4cn6gML+y3Bi1lnCa1NRcjEEE25tvB0D8YDTX2HcJC+rQ0nJ56X4gyQ2gCdl
Ma2wdN9DphWiVbYtVgPfje/kKGcTMA703riGh/PHul7p8s7VwkJj0riC3mh0u+YS
AdvxQCXH2ZIz6aRJ/tnrWuBcTM/R0a3ooqf4MWBxCbsoqoph8ZuReLlLyBm+w/ig
i/1g8HlT1Cl4rHJfSVq6Rz2kykabqcLv3EqgPPwI2whRhqkmFjBzjHi+xg9BCjEt
5aX60VC7OMsw3K07pk87ijZflfjmUEUxtSMsgADDcvlocRJX8aqbOK4KtV0MtWmB
5FWo5XYp99psvis+0H03z9AXddrnAXHF5UsFAN+bcyykI4NkLam9aUv025KCf6lf
uQCP7Ixa120ZtgrkQUyiAdkx8w/7o/ODbWt/9Z4Uj89k2Z3gLVUuosX6v8u4Khxj
0SDKJ2b1q0dNMxCz3mM0GN4mzxphje7d4RocmKSDiFP6hxN83i2YFqSMxMzh0SzY
hV8wpL45NN8aCGMweKbCMNgrpbK+yIDX3dFnD/aQ7CrCAvZ0mZF7c6qzziI6wSSY
HcTyXZt8TF1xzXgj2Mx9xSG/ujluNjcZYIj6c/EO6bVBk6hswnRGGCUm25N7SYBv
oHR0ZRdlfI2F23cka05ZZgToyVpHl93obpQLRt8KNsJvTF6Kl7HVZPGt/EV89dYA
HvEy/IqjE+cRffpvpywdchobN4vOyjzjzRaTMMtInoNGS2O8OxIQxwIpbwC6NdZn
3toCJlXyeRYnXp1tHXDJU4exZ+thraB5/ULl9bgDyIk9z70+2VYJu5xL2b7dzTFm
TtJETARAVQdg1wVD/1jYPy7pGoe2AnPRuEc1YPsdwLnHyyLFbzVCKdllpKS5DmIB
FjrC0Tz0Sz9+TyAztFZGZnhAzn9hHUz91q9JP8YLbc3dPtxsOADdUjOte7FQ+Mp8
wVmCoQPCAtMn6PxxZ6BZhZTMuccK4doE80D3IuowXri4dUm4CENzwRNecs1jRUg/
hAqbP5yBxrtO3xuKQJt3E4lfkNrOMu/LdfcPYdfwKzCZIqp5qkbkvifsDRe5Lcgo
SxPuNHT39opr696eVK/nBi0o+lS6sEIBv79aWiy//dhAnfggWGI1sr2jempb28nU
R47uCi0yvuvmiX2ti57IoDWzSWrkS+2VZMcb2qm5OSawYIgNb8Lok8QpJKZiJ5zH
/sCRjYK6nGOVAvYwp7WyTYN/HgXijHogmBPb+frdyVskAQMa45aO2gkuM9HYk6ym
PwhFfQMLxrWoDie7SUJITL4NUEM94EiM5ApGlGAsX4eHJ/+GpzvSVWzT1zp6RHr9
5MeQBBwXKBrSBhgCbZEaETHFBUgRvdbRSXAeZ+zbY0oGoShBCgeUIrq46yfSx0HU
1tPW6exr0tmCma4HaEiIAyaIxKg3ddEJTMUVEsSacYSxUfbkqxXu1IwCnVjHzOrz
jh9HQovfeB1AEVjzJbagAD6hNjNAeRgFrGLVHcG58tg/t7pnC/dcEsj56EVFcYUc
tM5O74rBAaFhTMSFQx0R/hX/mwPuWZ7Dki+y4ymG3DXPHftuEB38ZaZrInWHuNIZ
JZrzDe6LcGPcLd4FlDVqYFNtNOx65O9RRTf6M1nOQQZYbKRGioifjhuhvkaEfPeB
9V9r4Rlweba73fiNbdWKtNWINIMU86CjxwQ/bnEElF8zGsDDjCWfSe3nl1p8l/Ev
0UMyfUwLO9lDfWl276eUSQ==
`protect END_PROTECTED
