`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WQeOXLLcYlwHwqBjQ+kZr969JS7tUNvFKB5P2DTFWiV8U0NkZGM8FgkD9sJaQ61G
nhyCiNgecLZiIX/nLWDwuH0M6wgS0tpVVX1BmjcFBvbOUZuxklG/dOfW0O1cJNCH
B0TBycnyrXWRywdfv2axXM2HZW8g408nyUMNk9SSiBpQ09Vgo6OqgVbjhtrfROXE
BS4plalefH1bFF+j8A36Jb8A4zVdt3ttWC8URvd40jjs/PxxcuuFr53OcWzKB8Tv
Fpfb2lhtcGqw+3Nae6nHG0v/m3qlnvBKaz2k6qES/tci62xa8/aUDiTKV8Rn1f4Q
tVlT7RV+OZNPOvNefEcC06ac+z2mbfTBcjoSIhrRwSl04oXrrJ/hRdbEzS03luLo
vRYpq239ayaO9fFDeA82ZvtDzS1aGr49UHAcJfVEOD6dMfobOXgVv6WPC/0asOJq
ebDHw1B4JBk8uMfbHuiJuIMXnSQNJcYH6JocRpTI87iyfjNXAZ5ndMcuoxVWhBEH
se6Gs+BfwaZR2XVbyJg3YE6REtznLcWrNW8BbE2DHUtg471JvVnaF2mj95bhhx9g
qE8E9SBQclJNZjO7tBZejtJ6WaOE4EgBBUxnPWDEJPvtjEutI9EDVP7pfFjWn8hF
gNZrbQLXrV6CjcdhbJGGas4NQbBtF+n6YO5qYckKbYmWdLy9KTdT6IP5gU36utXl
yo1AlpyjTe4CxjVecWFGWe6iOptxoCfY0vSihFAP/sA27IX5p+J5MqI+sSeUUorU
XwSfxGLKXVpVPfjpj0Wgwx26C65eQBZXfmGnzDZSn2w3isgTYr6iv9W77NpbL0bB
IG78vi+wYgvMbG9tyLv02zPwhwr45HzGj2ElALbYhTQrCLvJp4pHv929dj20igB/
LtbAbJt1Pbtf89r33j2v+mqfPBj5SZLeacGrOqgiRZyWIVlR+oleOJo2VFBNimzk
Up4zBZzBuc+2YoS3mkECRVDurMSEDTMQ+/dKt1jvp0f4QI7+4r5lyQGTwjU6IgfF
XHhF8HslIJDbBHXPUTQ6FcF36up2UucIHLI9cnz2mD5oeRkCX2g26OFnbi9065na
4wUBc0w1t4HqStgzdBREmmLYoNTpgGZiUTfO4iWK89Lepgw5YmL2Uy2NJuaOyH/O
6DuA8krdeRuSWeVwIBn/S4CevPakPxzY4CIaHQbkbuAbT2asPC7cqW/TKeYYKSJK
iTDSYd8FQUeUZe8Hzv8os/9yFIUlIhZ09e9lGMsfhMLwFHJwuKhQ9nimgJUVP/EB
Qmui/pTrEjRzNnbvcKI+CJxzA1rIKJLbOB2Q/ACCxRM=
`protect END_PROTECTED
