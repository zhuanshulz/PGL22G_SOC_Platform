`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qwvrM/BGlFpOvJRQ+bnVQKuKCmA7ZY3jYPe5AQCtXjsP/0xwrCxnkI8INsdydpMv
HvuR38A5dehjmZ9S0kQPu6kM2qgkOLOtrU2MU01+2eoyeQJu2xplhIboxi1Jsk5E
FNCFB/2KwQsnZRK0cRczwKjqYtUMBrzzkMsqtFDbLRavKR5jyVD96IjtwxP12g5T
uQqJ07myL2EooA4eyqMO4vGJmY6RPclMN6BQWYy9meQFrmV0GcvJ+p2dmGN+8rxw
qHABl9X069W15+eWo8Hbo+mHyytvEzXPmLR3SYH4t6bYDZqzpj5XRAVoEe2H4tM1
IiwJ3fYQ4hyoNp0q/PdrK8P9IQspGewLJt27Zz+1GKDURnVXMqusme5GHT1NNWB2
cRYfKUGew5ipIecJcrhBVw1B3NI6n4y2lxfj34Or0C4l/yzq8thuzU/fWi+xUmar
HCn4f6vlXMRM1xXsRQKSOVuh3sjKHfh8/M7TGOxo9zAJ+cpEU3Xrezgz9QurMHTG
qVN/gdAQdqAlvprIx11B3Sx99SmRV8Gz32+7G/wYHCeAn2z4JHGNmR7tfFXPYqV4
/bmupd1YyzwwxEXHsYAgepcgbHWmPeEGcSWgUb/CLQ9tm3U9jloH0Qv/RfsHjxHO
or7o7uCWoOVXwVcBY/XUFsVb5PGuEcp2cKXJ8SZwFbENdI3un0PNQHS1BdEAWCRc
dD0IoVJDDeT0faWzccSF7wRmqBzqcCoicdzXIsVt5N2DVy5SV+tKREwX49uiIXhG
+652jN3Q7k1dE9Sh5wwSlHOCR2TL0q3mWGwhWRGy7wDCZfQwJsFYtrghn70Im5yz
VfqshbSkCryCdFzxj5wfkBo3fEGHI+3i8M+XaGtaM3bOVKTL6ghurkul4U0aWMEE
KWJo9NcMsNvxhyl7+FF9MKOqoUMGlnRT9n/OeuOwMIbXR66fVJtwvOmMosMomwFB
86wFBpnQNXOoiIAbAUaxUEdtCyGFNul4HIz65s0/6lQ+Vrx4mhORjgTOsU8+yXu6
MwJpuzfD/vMJDpEMf37t+FabTs6PXEqvf5ptMsfd8m+bYbDlTIgHrQvGWJS/lq5p
4buxR5yU/E/FyAP3iPoVRi5vhnvOGJcWYWod+v2radoPuGoQQrP2uE+EUP32RMAz
QMVYQX99RlS5sZYkjGMcyk/y6JgBhCjibERZ0qqCY/cJ8kxy5gbVdmU0wnyfjffr
0kR5zdNPkIra7nU3I8HWDiHfpxON0HzR51v+YMtiGGvc5diGyoLE4b8+OFFPsOG8
j8kvhdHOjjMoyggoy6zydZ22GI3LOuTa4UpH8hjrEdOCzoMIW6J1Tjfzdefd2ILX
SQwWMoVsIhDk81zVpIOn1I68jK2+7qux6tXAJLJoPIxLveK4rtaI8ioZlGvLuPMW
dXBGpoJkkENVm3aE/z21UUavY7UINxvW511Gehym0CvOo1/m15Xc7gKLKfBHwFc+
8y+tYw42Epl3PcduToGJ4dd/Eo4oeUzAVVXtYRSoqwqZkyIBvPskzPlC2tFAYWtt
tj4x6sya/tSGgNbEcgx58G+G3XpXHU32AQ8I7ScMWOYxWujPUaf4xpNkmgF5HfQ3
ytQANOlQvzCmJrb80eU1v7uzgFnO3uhw33FC9WTh+9TKCvtSnOX4X5vcqdP0GPR6
3H7+rYQeWHIk3sPKlxYoPq61cX7iUlZzY7sM3ZUMFEF8/sR9XsC+ldcf6+ce8Jkd
ohJWCTnOM561QoEvv3bwksTz3fhqwMScqbWg76bW2pAvDoM14b5qNpGNhmw4TmZC
WnTi+71M53ji68oT42k9VnWVZT/V8CzcRFoYRaDMl4UCh3jzo7Lr/QVWv9H/3cr/
8BUxNXrBZ9OHORfaqygTkC7AFFvYM5vYxDG9AZmUmIaqxSTO2r0K/CNAxrYx4mZ2
ONRm2Ze9lYekuct9tqi+kA+u3nKHW0uBSSOWLV57T6gA+t7agY3wUVG50bBXUht6
o2d0Si0364BR9sT4CqYknZDcSK8/c79vemDUtabk6HpnAUU4Q48peHXH0PwKe9Hi
ggGfZNxQvgsrGK8oirxgHYyT2V8DX4oRp6Sn1Kq6V9nWCVgHlHW9J8YNcRmBbfQx
9h+9QofS1v8fcKLvtdb+VPnqwlz9Fn/7+MZdkWFf9H0rRHexOylBWQ3Dcu8rvqnq
4hLXwlvdi3ULru+Ek+gHLMJXs96Lp+n05hqsoKyoI2IOjeNkgV/AuVwnxXGfcH0w
27smmv04CLPzk+/F02coCNrfaIo7givIfj/TG4nUsvkbnqdOzAaQnH/C9U3x2x/P
0SXMqP0wc9DKT5a/dLs2pTIOrYNSOSFh9nCUOOOLtluyzi9lurirRrwswv02oueo
zhnymHBl+O8ONgzAZaIDZi9QvUVRuN8CH6pYQ4CH+SiVhAnGlbQ8CyMo1Y8MA2nk
x73i/XMKSwoClTVhP6i79EmlMWhh/9MnGRRib+IRDNtUnFkF/+ansNzh9BcuZNmJ
7JAphOdU5t9wpD2XX1bSup04Z3C9AGaunuyruLuiYCtiAvJOfCRJubCNMUCFp5xw
ZZZHN+AO/wiZLPyEVf4SzrX12lJY5UBwe7Rf7gUrk7KnO0c5oKuMUSEMPeKESICP
9x4Ky2KDYqSrj+G44wyy+nJgx6T1SdXxRx3c5eJTB5PQ6kWgUSyKuG24ywVPzhf/
aIZhM1EVM2mb3Ww5Ko2Cce8yZV78Ar347XXM1wrvmC88aTTYa2/s5qklQIr/pvEC
OLL/M2bYxoLklR15vz7nkktyD+7AOy/aw0Wwb+y+DzAzJEKcA4XfmQvXQwg598JN
DaxRi0E4MnHRbxjJHoDNoecuFAq3hEcX3RVFADlYMqK3zzoXyjPPkHwMIlfE/Izm
kG9W4N4AArsArmpzgYqsm846wE8p6s1pKnKFVZOYN4Cdq665Z5935LCwUy4rqHWX
RmYjMAL9I/0JlMoY223C1vKcvSo35Z+Jf1sOeV6xaBrH7H8cFUsMEgfocIBQx0Ux
9yLcbQK/nN0wVLGeXj86C931ZL5RYlt5aHhhaAsJHjHINT0kMTwJ+01g/hXVCt+k
30AysCL/LVGLm6HyJVbiZSLf+rD0juA3eMJoNznCYZPFA4mTdBEIfk1xcnYqWSvm
KXVOE30e+F+TWJBD+vO38UiKwS8//zYlfR5ksU7b52w/yNuQU3aOaKhGm2QrI3Xl
fewSh344QTg6EhgvePJU2v5PaVrFCgqy3Fh+VUJ+EwDAqltTq9hL/U675DQy/3Mm
Ax9YrsXjLs4xHrmPt25iuBTuaClJM2fXs/JF1kaa1Bbo5KpnQTQhXIQiEfEBrimv
Ag2pBexjz771Z4AaQOPlwwQGvrdS+nEPfkn73J/bn4eX+gFe0698MzK245DRp6/h
TLeJRNL7ryT0zXzCmncFKL6Nw2HLIkj3R93JDdfo0GU2cMiCHwsjuk6AydX4JQB7
krNqBRKe0gztVFvCSeTOz+v1rdpmaIIc7in7XcNpDG0blzPjs2usiS6a1pkbeP19
PhtZB37AyWsL2pRtJ+MgQILeHfeuusWy+GUGBG3g08+IYHE8wRlVun+JYTRoKVju
cX6vrowYSFQJAh8Ptw+GPLutWqlEzVgUfHrRoLNsCsg0jX1o8AwpliyZ2SAtNezt
P5GaTP4/TgwnG/v1ppL2Ru4flFaC5lPdM/BjDz6YaAq90+dZ98WoccDbu8QHjfTh
szcEOhZXtL7DHF6GDz9NyNIT6rZ481PYjuIhWF4WDPfAiGXDQzF+fxQkRgHwK5gt
7PRlMdGVnL3VqfDH8jBqhGJsjpR6NJR0FXtUfFyTRZ+sL4S5yxdtCsgF8SVD8y5D
AlcRo4q0VkgZLmYD+fVG56+rvrNcPEPnQX7FXi6pevTbbxeLWvTdyJ9JQV3VbFZz
IgAxYeUitvM6kACXHkg+bYRPiTRRXM9x7H3q1vTdAQ+W9rSjTlKaB1tYm2ACwhzv
l9hCdPe4VKLS7V3V9Gy5yw==
`protect END_PROTECTED
