`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OysuaPakt95IFBNDXrQr4dqIDq83cMf+2oZmId+jXYQOI+yxgnYrCvR+CaBxBr81
LfJ0LcUj2ZCHRcXFQ2v2wStrQxVa/clAsnOmne2+xb/pQjR5qcSHKwuVPQUCTCyT
7a4clJ9XATrqmG1cvj9I5pfqAbvOfkeYcit8ig4ekhz0XbGhGoU22l1QNZLEYVe3
lZnlVUjaQgefkOHQmflmti9lDcYQNi38PZ2jDZ7iaI06YTLVgCkcC2Pa0t7qR8Xf
yG533OaICAurUihRwhiT/5NDxa9IstzHpt6g+pPn+oYlwWYlju13XLC6wf7hhG/8
lJKu174PhWBzznVjZnCDx8DemiKfWd3+vx5PG+KNkeRXqJuh3FMXciwaJCMzt5qC
LAW3BOPzkO3Er6tlNPMgnwtPDk0iq46E5t2/hYFIL1OXEms68izhgb0V8HkA6nqb
aWcRyyXjzvTEjj914sytIDC3EcqEhbG8g0V4xzvmPGtAG7ZDZ4EmRTCMV+p2Vtdf
z008JeTr7aefVuKvnVLuyR8YkmxY6dPMhLuAezVUmZrLzPP146SAkO6BEkgPelzd
QMjRkbLG7m7XT1fLNOCBCvCUPEolrnyfoUNYpYgvbM5SIGECXZ4IgH0UfZrB4jX8
4qknAYTzww21LuIYQ4YEgi4Ou4Qk8FBZMuaXoRok1aoLymXVlUr8HaXoyjw1CpiT
gJauWHrmXpdxXHj5bmwlTSEdKdNLzPSWa0DuPDsXCOtNPX7M9cbvEt5BibebHqyU
BNdvnMdCv97NkFnEJWNHdzizD2picvJE600YEZUZntjuWuVt/2PjI5GirFlOcw9B
wsd/CDEGDN9fWklCEI7xpbqzwvoj7gQ2dvqAh9NzkYDzpyi2jmGmYKpz2+rmKm9S
JzgxbivOuObRY5V+luqFeyX5zdxPEcpU6xo5vsUoXeD240hUAHi5wBlTQoxFuOz8
aZOKE56O/jW4zu6pSycG7xtwHoHetmcMjqkLyjRSLSZXTeaVX7fHZdz7xTiRJoK0
NDT70opc7ZxNWNeSwAApl91jCb2llMPu23Gwac77aQPu2r/CHCRxfuMtphIkq8Ud
ttaOvEqZ5tFMXzhL1ig6e9n5e2wd3Y+k7IVa4Ac+kN0UDLV9fIh75s/FcikQb+p9
RL/FjGUWFUWjU9tTdnHoPaEUhVgDNXPFw0zR9wqub5E4aV9rmbChoy1o8o+3qxPw
Wlygm6pWLChhKOPe6EbOcT90elK1+6Z1nTwMy4Wp1B/qwov7TWQws4zqGZXUy2Fm
4BPIYDOFDt+R0BXRx9TxQcD2mOfbYpKUOl+F9ECswBP0yoicix76GI3fxyhWJotc
uyrxVWR0jNtviL0q10a1htJWkuE+5xhK9MJTHKHYpXZHXABVIziWEU8MgAqelL1L
q7iWWo/KZXTeOSCA1a5uvBAXkPuWRkwwdoCRxTPryYF2pLk21/ZdPJrf0n7G/M1V
XLhvLTgPUL6fASfIjUDgiiWIQAVNu1R6sUNRnN2dArcKrWHOEEb1lq0eeee/K03k
ENXoNkOR1+vK0HcVPhbiQ4esTnxHRSLacdA2yiua8aniA0emYnnD2gOCBPOZBQeS
/j7pLFNSZoa//qs2zlq/yD6Fu24qkIh0k7kLaovCjX2N5AyY3HNPZmWka5WCLtzd
Wk0u0M+Eko3hMmdf8hz6G4K9l//YMiMQF0Y9KDa3FTAzIHtBqM0oBSnAO0nX+Yx8
`protect END_PROTECTED
