`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YtVg/cPYpIWESuAO50TxRryE5Zh0ZbY4KOF3LryE+3uFaUzJ/KxAUh4oDPA9DYoj
rANelbAfQvKoS6X10zFAhGifOgXZ+9yAv6m2GYeStsTQfGxNyYRmEGHvMfBswkYZ
kntYEzwsxHmSjuMkWZR5vMsxn172dyCbDwuz1WIDsH/Mf4VJ53+8E3Z+SI+RD8Ys
SEamlrXIbSQQ89s08SKr5vxPKC0l4lr14SUdCNBIj5iS9QEdXpRbNrCRpwR9xrul
7yz20SpwllH6yjIBsH+k6jg7SFa1i8QpTXtjqohAdbctlV3GUTfwUzEXTb7npAI1
EYYTDSj7o69Jm+xGtXFLkyVFzzfzSFNqmYRbjV3x6KE6ryM+8BATlvAvgMTakG3+
rBzB31rZXdTDkbclRiTSObSD19mzDL6Y4wuu64+LxjU=
`protect END_PROTECTED
