`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mrkdjXFxVNYDlXPt7Zbk52870O5TKVUdBcG01hszpSUJW/CkLcDMTVWmhNZZThwr
qp1Cxhn/zUy7qQF7bm+EGxhz6KMKMoplWV184/+xkoRaumM4LooTuKXWev3ImPM7
E2CtAtdrQjMwBCpKcclUHWx6FaXlxNSaQ2A4XMLJ66AKfA9M41XTHEuLfJ5aSI8B
Jcd5Q8jnm03SfCQ85J3PY+cSn6h51Xb1quTdHbFF3OkFvO4LItEavhtyTQoABl+r
NiHzN17iX2fyGVkBNDZB0Hq4CU+zrzJS51nhqbHHAKqbCLP1q5OGQdoOSwAs6z4J
kfZ6KBiZtyfPGZ+0p2asJqKB8yZ1YSWJnNWDPQV2BLGRsrVs+GkN74/lZmBv0Q8s
8zlfi+LSrk0AajivS33l6wQ6SgCIJoVpfCNZl2vjIilx2YAhjZ0jIzuw3GEKlYoH
ht9vhNRBfmauOminElURgmJwmLIurfTcz58DZ2/ow1VdDwqNsGSsMjf3yPWi2zQZ
PKCsn1yXCsMfuUlIKD6BVhyhbhyiRK2QsV/PJtMTXULQD1dvskXFwyXmqLRbLDuH
mQzcsy7Dibi1jUXQzobeanyX4V1RLjpE7QzcO7K9SUaK5IPwKzNmFAWq3HFBeGIv
smv3HRDTOxK88BgZpumcUYHZRriEkO4ALP6tvz7jUIq9OYZwAwY89CRKMEqsV4xS
x31znQ4VrGEueRlCkLqxxPGIK2REk05u1qBUS16LfPma4oB3VzS5VokYr1Q4va83
CsQZv1AEvTmBWfNGwHd2HpaO/zQyDNILZak2QTGc3vBGpypdq+088pi7s3nLLtJA
XXFVRjrrge0fdUX8L+FMeQ/fMV4FLdoXrgEocq0yJhKN7uYczRz9XhzQg3hgYx0C
OdZmWw7Gy9NT4WYmW4+J5wxfIRtX1iIfkwgbG4WbzOutba/x87g/pkKX4TI4/4BK
0XQ+DPzJSkiLYv1qjOF3eyLaYFRh/LU6FBSHCHURV4h7+HDSGmLiwVkYVUXZ8BFB
E1DmRtSu9S2aq6O8V7+Mi1L0G7cPXLeFL1v01zy5LdJQgbqL6XzLRlI36DIKIKEf
YGW/qMC2Jm3gGWARCz7+o0nbAIwZQcANsW+sOh/fzPmpc/ZA1xgsDX3FdMHhhjNB
5ss+eOAFMfBED+0MANEYWwUW7yKkU6CyVSxoNYxM/s38C6eOUsC2BquaSZZ5a8hc
5ySioNr6OSrgCU6gRFmvwk07ZZfi8cUQQbrEz0A6zmYfPvQQeQwJx/qov+nMLcnZ
4aWQwOCsWMn3LgnFCfdi/1zo1wRTuRnL0Oq5A8SzRfU0MlwG583HzE2rdzLDVbSo
qAZYM2O5UojwUypRpFuu2aAEMa+SA0sVRwNZa3YsBdNkQlUJ7J27KXxE8SMY27Sh
2XTvhgxu2VK+w11+6CYyMNoqZ1mAjQBYhFYzp4qsMdD9+l4AM88fdEDIOdPkjYSS
EthIKAc9EirhcRYP/Pu7wwsIQT0be+Q6u6nELoQJ3SUY2yR/6T7sSazM958k49bW
+gWPyxHX5kxqRiQPx2s/3wHml2l8fJEixnYafc+0dwR5t0zRrIIyQB4wX4xXyqpv
bPOI+vqHdELux8mZsBiSS3s6daiZkdVyI+ZpWEpZuulh67e8F8MkZbGB/41oDF0p
b2byVLcJgMx8hTPouR0TAcaa7199EBc5pOLCKz0/EoTctJEJLvyOIrbxb2YzZDDJ
/Q7igj/AfK518+nK59uveAAfRGJjjnM0D2F6DrtHepnC/yeWV/m8RNoLfxwW9+sh
vOiZKRJIHBILT7HLCMEKBrPKeJOy8i8p1vwqfrr17XJAWb7TdtnUst7kBPjhJV8+
Yr8HJ8XpNk+yrDPPTxJA8BwVB6n7ESHCiQ99GhzNrv/m76O86Ho/ECYgO0dpm8W3
z1IVzPIQYTLV9KM5kV75UBI7qw6m9QQEDowEkw+O2n9qKISrGTTwZTHBdgnElbDg
XFgOOI81FwCLCqvSzJSIuaKIKiN0MH8vA/0p56puhUvb2wIJ/fH7Osm+QKfuxp/o
UT3Flrv6IURWgqzTlvdRFllUKpBUdqYrWQdfZFifS/sgb0ZJv216NHd7ur3a1Hk+
xgHfQVNZUz273eB250pxUsP6WZ8dD2H0Kkc9/8AjGB9X6fJ7yP/sNNLN6UnVIQTB
om7mmKibq34xy1Hu3JNc8Cl8PpS4N0KHjXYmV0AKYrDdoKO9E8CVRiuYdqSdY0kx
G3tj37bBLuVUpmFmUcMgT1WxuaCJSAcDGozWuyhGICWFNEEDXwtSIKLrOL2ZI2au
Irj6r4MYs9E40OPxAAQGx/rRY3ee/eA5DKWnNhR24lcvMHaRufIaD8qO8RWiuB82
JVyWumqMqxX85xkKiI2BhvoEZXtV7aY5uZMQrR/bXXOtJn8fOrp+BivAvp/vgGmp
7w74ZlQ9YcNSh8031sSueYvHJQ5xYL7IbwGBoaO9Sh/YmUZeLN2yChnX0ZPblgWH
5BeyxAYntP+PR+7nYgmVQf6EYDEH6VNL3/Vlm8iq7kqPq5B1fXmx6qU5n5AzVJPr
ZoW5PKgofWZn63or5TOxL98K0t1lcVd/EuuSyhY33OyEasH+jdKuEuIcz+/FqLF2
OQO1W2Gx0S51+6GQCPEEHrp+sVHicsKHGD1SB9Z0xJq3o1SUHtXPyUR2TFXkx5dW
WyM+ExGqqKGyLAURn+B6pQT2L54pS71WKgbGuiwbhqijxDEsf6He1UALOhIoRXnu
Vv1SXcNJqocnU1TE0hEFZkAg5ctKuFgJvq50XnnEXqMux0rlvTqQZjwITHXP/XNy
NMScd2sOsPFAn0C9fZ2DhR0Dg2QVlTagA8qu3AnLyMR1qUkBG801KDFJVdKj40BS
jxGEHlD34hxffinY2UJ0JMMU9kQZj+RsUGh8KeZ2Mc1/85284fLPPZmL30msdPIs
XeR2tOPqhjkryJHrWpmr7B7NPjKkyQp5V/x9PnHOHuply0p/K68F3ljWYpmbVU8O
KnazNDTUFIiH8KzvQC70BaOYtRJI9GdXG+m/jO/h9zXeraG2XWq54uYM976sTuvG
1RhuPzcwsuf2JDp/8r5fC5uAmT/clQerbeacWjG/7rNLNxuOqzWAjqjEb+GiQ6hK
DArDh1VHZ0qg458ICNaVJbX2q9iBh01Kjb/mx51r6y/2BrFMX/bzD55sEyqzRfIZ
xYyDGun3KdvEwT8DgmeLK0E3nsqvxWxnzS2Krvm6aujIR4O/XHxW7vSzCEKZeOUh
FAE54HcbVJa7OyojsjwYt7c1oIgpStNTSeAND6Pu2C0kd4vZsrcFGE6fNAItLMYd
v//sGtom9CE7LbZnzk6XgOlVFfnoJHGqpD4NWIhMjhDRQmtOCjXhEuU+/yChQXB3
/kmHYkZUTCXKWC7134EXOlzYBpUzzYo8pPtI0zIFpm4ApM/fZn2iE+E9an3FGsqT
KXwYKvQ5PjLokXctuC2br2mK7Oh3Ce+/2psYhPeWl2gyOONAvLa0qQUwNlK1OLhO
daIll4Jy+qwWxHvThe/FaB+/dtompSJMUg8OhA0hjFfK+APCHUTDiIJ8/BVD7TsF
oIBDYvCYLwSnmCi1/sutgDTMMoTZByvYZELhT5vEez4qCGgDOBeXKNzG1pA5+t9t
HN4ts/UBTR5zHG3s/wF0abnpo6KpXn4nEY2S/4sH3fcgb5UiXdBAx7bURYi99dKt
53sql3/lMoloxUNrRHh8tI5/LxTu78DUxcJoHSQLJOxypxiBxH5bYuMGuBvaK831
b+8gsGOfkZkH2RRhWJV0yzK2fa/FIv/F2Vwyv6QyVJZekwG2qOYK2Dj8bJ6SLUt6
kO69jhSUo5idAGCC0xqphIHOzwkKfd2Q5u8sLGXNvrPCt5IevlHGyyb+zTr3mgra
TI00+iwfsrF0va0ywg2rqpDRbcFu3YyP4pBQdc+H5XVnEsq7RuM01yGTPSiSxaEq
QzGvnS93uQ/IHiDJrXhQfGawVnZyiETdBN98YYgjUK+HReTndzuE8+aTcm0GBGPz
7CyXJdvJYdWD9ygnuxohtjxx+40A7L7Ze17iFHuJfkahP7/L7bG1AcY7piDJIZ7n
tNGbQKLzXSWnnqxXycMkLyKUBqQ68fRqqZhlwZsRXmXYfAyqu4Cjuc67bnqA33B/
lJEz4rHSisrlVqgqGdoxSiSmYlO5Ctrhv/PvZtOxgczEjt13NDRZfjkIiMFcfU+g
e2QIMcMZfs0SK9AO5AkQAgq+QAoB6eUicXa2BU459zdLdl9HQzZzksgBJ7cw89Rv
2n6Q7/wjl2/QxHIZOFLKHkhgiEajEudB1714hd4DGAxAflT9GiUnjrEb22gNBoCf
jOKy8Hemuc6h1NHW+UiDls41iy8UxWUm5G2arn78RbSqrcQUe7VNlWTJrljtrDZg
ZG5MwzmbD4rsWLGfZePjpQXKOztNE8c5Mr+MvjWebR/nLlC1QMERHbnOn/Iiu82i
tzkTGexKaNxFScEKtByvA1gNF2xdKtS1xN4iZN/4Vssz7ecZzVKf09AaVE2KpwHi
hzbtPxi0PAxp83NLlogbeKN0IyPzks3K6AoT2CC88SxZ7g8waJnpL+Ym/u4HorB7
ixB/EwM+wrqnDcofC9WRoVc0iLJdt7vsDJhDu/MkoYJIcQiv3kCBEIEL8K9IR0jO
p6owckd5Gtal+sAk2b6Urr0PHExebxqRVK0zt5PpHk+UTdLq3w9Wn/h0h+OaDElM
FB4MI+E+uEnUrZql32sW0E5urc8J8zEZ9kNixk6ZZtFf9IGNrtmfja+XGj0Oui5j
h9MsBYOmoRE9ASmm1mxL9vzxnvCv+MuB+NrjRlYkEWlok5bozdMZRJr9LQ96n1tr
zK7h0rkGMUqMjQU0OuclI//I6vr8KymRFzcmV3YG3UzwwldBjUbVy30NTz+pfaDO
E7jazZcQPNslIXwaLE3gf6F6qVUXafJOMNsxFHDEcvWR1nN6apyGo7PyyiBrWV5b
74ma3kp+GbjL6KPXE9Vj6yCwrQnfLMsFQMyp1y4kmWDsKcli1g6/iWWAm7VbmKG0
4XsfrXpLzrs+GPhDHcl/x+v9379RPeePxcIWZnY+s8xOuvXmVkMeq9kTFfvLfOmc
Kz8M1MQQZ6QTGJQATsOz+ZMeeX9s/Go+EYWpivHyzsFYydGF6UvGYA8iRWKtnjGP
j0vlqi8IYOirSdWkWq4SKj6HMpJlmLVfxLqr+19FyFlJyGZf0ZxwIGDiWC+rEaza
AKyzeF39k4Zb167UlXTEPBZ4NgStn2BCVnePwqE/QHcS+bmmZu+ceHA7IFJkdD+c
EnOilPSZX2WlvT+X5wPSJMFLQdrmx9GYVlDj/F3nImkwFapkvQKpEmdXMw7PTZ7+
+I0deJlsqK/FuF3fBnT6zhS83co/DWd6e6U6gYzg2bQ/q/gV2MJrEaiEEuZgamLB
2qzqNfXvhSLRzh3HWQoCoth35+Lg6teJgcQVh+xOsXjvrkQgw+Bvq5lx13PZNolY
HF23RbQclpJrk62MGZXJHO5u8Ynbx93AuW2PIrdBszXUI5OZmSp+Yxvm58zoQSiz
IZE6QSTcxS7qF1dImgpqee1RIosl02JSe7IwTrPoVQr4YkTwBCJNPMIh0hJbQLyf
KDco9ukS6YsFN3hmtScq6EIr4mwzBIZwOV8RWKo7uoBdrMyFWv9roNcj1JVxgYU+
MVbb7ARSuQTfEVv3X108W/JCStQpOY7udHh/VjvvrX/0xSS65h8jw07tZF6ikX7m
BZA9PWDja5f5MJKvZq7b3Q2o9qwnA04zCfU1coMku2aTLVmYFB3C51mUqhsLU7nM
/Oer2BxPMCBKun7JDtqtP8vbr0dks60V7JeKCI70uk0SdY1dwqXMEffwlx9SMY7j
yJawxS0kNz5hnTCT+0y/1c3V0WM2BltKarclCNjmXIhbX3DzxraQAhIc2v7qEwv7
FI2CDSlOctxaP2LYH+Nvzfi9kMlifKya72iKupahr5GzGgIiHFNdbz+QXkRg/FgC
IaOQ3bZfrK5Td6cu9ItxXcbu/a3iEcpFl21d554NXqF5uiv2hHuf6f602XYO4jN+
QJ7Alacz7DhcKiM9no7VAT/6Zr8xXffmkCz5BdBtPYImeWTIVt3thxjZ3e3gus+T
Np1CJbJQUm3+w7Si1uzgqm1+fV+kxmmnMZtHQKvRp1c3Z/F3vMBlXlMBlWg7aPAM
LaWYosn/fs+0MautGRPvx+5dIcKy5+ItblpGOXohRHvKuXqNgA2oVNTFIIbn1Kab
87SmDtsKYgGWvOZ7nR+8A+jgDtMmbFNfZca8PPnIFw87cJMBPYZuFMooFj2tTieq
06d2yhvcni1tkJz3V3OzGTFX97UN3Unwfw6bvtxWIznh//apNG8nIO4P5ctk0Nsr
MmpoMyAGPFsrOdzKHR1g12XZ6edqrJqGJjG0/BjWDHII7/nXZvIWt7MDn+HtYAWQ
tF10R2eGtxKRaiz1WpzcqyfCe/yUDvxSOK0Uw//DSNCegsvAK/f9ak89rN0JqZkS
qMQA/JIRNZ3SbbQI94IBP2yyskETZ2QTioZdLPGsyBFT24S1sx20dL5ciN76O+Xz
ZbYXrQgfVxqGvC3FloxgayknPQGmU+wu+PY17rT0qj17tf2a8GUAsGOqyA7apge4
iBX7TpZHwjdEIUtQc/8gmU3WZNRM1YQ8znjLsNJy6moZI86bHu9r0K4WSznOg3kg
GIHbZY782lFKVBQhhNsI7SQEkaI3UUUxSOBNvX+ADLMdoGGRtFwSnNpt9C0q4gGX
AAYXCvELzprc+D00PhrOgFs8cLDjoFnMt28tcLKADcKbNfSyZjxTJZ8XtgJioSLH
cdO7ncOrJaa5GdJI16bEwV8HBC7T4pwUAtFIn4Jig3Rf87XTn18lqe9535UfW4zQ
tASwX64AW1etuzhaeEbA0Js80epePH1WGB6ALsiO38fXzhge0tcegZ0A3Lcgzboa
BB+dXjZePDb6wq7NijYo2JL9qpJVbYN5wX00rlAQVxdvKt4DmlN/sU/GmbcQA1Kk
LYh01JQA9tMjsKXjp6u4jYEOi2jYV9LXCXm14+Fb1KCE9cZdKCDNqYzCgB1aYRo+
79+CeSYh92Ufbn99H+aVYFN71UWazw79oDGyq/u2qbFxaDZ+TIE8E5TDmSHjJ7uo
BUV5D+qkg/MizxfazX9RYjDy5yee6za+8fwSUBxGWNwwF7MKbXLhwfGcQVc3Kq8a
GtInXMjR7BNFy3wav29afS07ZScmASSDmrz/cvHTCnb4bJhXiORuZPXv324jiU5Q
IgnSMrxuOCTYyikVWsqdyPy+m8b+nkL1vmihB54VJUqFeeS4+Tr8bT5fpWKYrw3V
qs3YRZeEn6yPKzHNQJ/hphONTBFynxV7Yoxl2DNFDwPWdSsYOMY1oKaHiEM5FjIR
BK3Nb4ZxfdW6HHEUMYUVtZePW3re+piK1SQ1qE9TBmCVS3RRtLvLWCd36S/6ZMEQ
iBx0l71iuP4zNssRB2mFIFi/6+lOhBo42fW8vX+HBfo7yArb8docJqoezj3fQTyc
abLx8EVjNOwyRxKq89HufhdF95XC9WzNwFiKorpFMITsSUrDvZafv9HcphWkGhZJ
0Ke7GsXGP8BUdfIxEbHs4FbnsP18PAxLPCciSX2d778stIPbzJrcRTUiGu+eR0VD
6FcrRedEUhFp4M4oVhJwklyGiq4/71+pfHUi5xsYhahkImWZ6eWi9dCSvJdnW3gI
9VzUz7Bv+bHU8XvSlHRUMuQ6f6E/R1EUJLlwj9pICMli+XhaIAGf2R7Cu0fhX3WM
VrK4OIySRokE+t2A2q6n2150Bzaqi16qdRH8qtn72YmoA2+MRSxU6V++9JtuMPPI
acU6ZCt2lJSMvCvxvglv92U1WOoY5BGBNB5HeRZ8kHvPYPe7JcuVQMK/TfUs28yD
C7/yucpobpBrjmuXr9Mvvyh3VUpnH4wWrkZ2NYg+pyxIM0OUSbjQ7cgtDr+uI7k9
inzl3qHmTjQBy+2H0ytqqn8crT+zlkdXUfczuLC6ROq/Bf+qVUaS71AoHKXmrcL1
Cd+WFRybn13NNrNbDdi/WBqFyl7b7HqSxQqldvNEQq+nSwL06XxKXdmYvFeuXitd
8lTBNlYAsPFh+lpYCh9JloPEBYylcygkJSHpzgRBaWo2eZQxNl7dzlOmpv32Z0zd
i+3Tk1sgLwKhdGNoWbf203RFDPsWcLPDj+NM6NvmX+a7ACGnyEYHxiuChviuAdyQ
ekrFrHrs+MS2x90V2a0xDW+/NUjS/wiiE6Nbt2YjaGMvJ1uEhGOobahr9fKRFIxW
fdwsxk+tB+xiUVd1TX/99RH7F+LY+qybwcEqyJ4VDK2Hq8DpN+yqyGFvP57N8kYA
6ON3KNWConeoEdmiHvaHJ3WFZ7W9PnHy2tzfsyu39H4O+kGYos/m8V9V4blURUWo
GrQgKzHBiVBONs+4JlfBEJtZgeuGkfbS9NQlsIdZpwCd701qjqljvM/q/2wDWrRC
bDfQ25P6iS5I2yuLZuaolKAyxC+JY3rWBtLSUcO3W71x7HBZ+AZu3XhvREJheIX3
42WNc0Cgyun4h2l98MtSQYFFoloQntDP0A988pjPSmdpRbMy6pIq6fnbR33dIPcA
bFSaRbgTscaWutzhiXDvwtj0ho9lqoKi8kPV3ef0xKnUHbFJ52ZRvBOe0s423ESB
xsXED4medETgPSAfYpbeckz036JoPiA+GM97OtSIh4NoDKshKZG4FfpuEiH2Ht/y
BPABdZ3iR8U4nrjwxBO7xU9g/d0Co3E+hTVFhoww2X2WdR2Pls4tUGa+A+iPN799
PQzqNOlGDqe7O8aPtgVep7JmTE17W8IqAusMNOUUs6fe1hbcwaxpfS+1G+ZeJ5Nq
ronfJwwc+9fGUiacNJo3fvAfdWuACl9rcCmOuhSVgRFG8ENsKI8ygkZJkRLZJsEP
D+YKwKDE5PpJo7ttJhG0ejJ3/FJGJELF73tndjnSRqviLKZLgKkCVClxfPIEuBV4
qgAAH7UM37FevTgbJptD7dYVkBKQXMuUR+ohk2DWtu3Drx7QyvrkHPc6CNxIYrvC
7VPfR+4fyD5HIEi/+0wiRRfNjbuPC/pt8qqyBQ01LeqMbOmveI+z66mnPgAAXTP5
vQhN+wrjGXuW3E5EsSeegaRtzHjljvIcJAOLbfGIGxYw8kypDnP7X+aGW0eFcKVh
RI2b2X8u/0EazB4IcGYAE7pDUL3lO1LDaxOMGUwiqbYeOStFaY5EUHHJ1jXLjhre
qPKp1XeyTJs/be+KNExJErXgWkgF+mNohimgW0ddf6NaNUkXXEJswTVmtpOQ8Ni0
rUjMQeYtFw8U0rKwkBiHKsoqvv8Lmgp58qK/tJAvlWchMOSNhxSlEibhDlEVK8hl
g78r4mU7GOWkJQ9rVy7vZMUxTac8o/m8YTF/Xm+bJKTouz6NdSGFRDJ5rnrXNYGo
ZdUayC2PeJW0RzrI9rx725prGl9dTbyikN/EKaqGdz85xNlwnOCfsD3eo+v3Bh8F
WSYPR/4COAAktw//g5VO90kM8xNcDqoFp3nlxxDRYjzqMTotVz8xbTZLw4Zdihf2
3ueAD+0KcpMy0VEqFkH+wLXyP+b+/VRn2ubo+YDOkQTb5QFfWzbeALZi0mmGis64
HjQxScgJRZ7IwcJPcjR1PmdN1RNDs9+0UOO/z2o9fOvjDhJ6LNF84u5v2twGf78h
LALDnojTaGuJjpzplEul9thmMGVtQ3d5qK7AdVLlY9RqAfmGF291JrxPC4T1jXgu
o4HEZFoW9N8p8G0/jmO5sQacdblc5hAR0racR+bSsFCIM4qRfKvzdetvi+RICKM6
u218U5/9g06gZcMEFJZQWIurx55DtuyfM4+KhvXbpOKhRkx0zrCvNFLiAa+dLojF
TzEJyTN3gegJLITWr5olzWHtDcvbJ2wqMn4TeWeiidak/JnkHffNFOblKgLf+A2u
RoKD8VCInNDl8zr2nXrHPd8aF0oRTvkko3oaeErYt9CoJ45tjnq2j585FXLTg0AZ
i7zd7fePSRhdfro/GEOVVHXh4mMjKL2I6XLN9D0quagw78fP62B4ZOe1SjQzOf8Q
jiHPcLqdTlCenSflm2lRF9hHrk7gKxMLuG4YQT2u+3s+wcfiv0gbrZ/lztgUOSxD
xOEZ8kXMhU4V5HZPQE8GBV90PERdQZ8PCV5Z+qQl94Z4mbfCVFb1qlJNUSsxeb5j
dunUENRiyKm+LpKPGmNVmHhrw0zNRWrITFNEEKoEza6epXtPSFqR2SFiuZl8KwAl
KjmW4hwhxBNN8vqlWL5rYsAuIHWkg7PiAaELSdvbyIzr7R6c4iOMJO6unCF6cbSN
Idxm9TQW3IFhNS2RxsfC5f1f91kFheem3KUjHQW66vTER3K9eN1GfsL+48xAczQ7
iM5rumQ+65gdSu2misvOjokTdW9RJscvtn/4SaBqV2kxCKeL2GmUA3zMJN85/3BH
5E8tEVDlbVLgm4RkMR5gWcP2FBblQC98kddo/USbvobsEQkPlMTBNoRR65d+oS7P
iY9Zx7yVPUqFcnfEtRZ98OnHpwYio6oPPfI+lamKpWO/lx71uVduULogGLLb9XNG
923MOyESPNTaayFH5l7KxhNuHgXA28RJVoXFpAgpY1StQGB3SWrqAXBWHgtYmLSt
284tEI7BhayE1CNPyLBAh3zs35oYVxnsWyVxyBIrALWbrgSEkZLhbjs1LSFe3ApV
A/KTK51Wzb37NzhcR2UugNvkePbQSnkeEGc5XN+tef3cTEP5WMk6Oh3sluebyckf
wRND1RReTV2op9xWPq+hls1zAVH+s0srmV/a2IfKMFNVPqn1CEr/pH+keCimtb+f
4hDOelCpwskX8UoaMMFY665RGNnkBZA/sy+P7ZNKhD7MEwBnoCDis2XQ8lRtVszG
+9x8vcdpcsPvdwOXXf27ZiyTtyjCSyvhZ8OS0Z19XjR2GUHNoQE+uP1nKdjmoT2w
NzdaNIwKKb6VtbbibFA6NI2lFvrFBn0FH2ACdTlEwJSYXqmGvd42G1tP+5VwDlTt
dNNrdPT2JBjQxs+28DHGYtH+JcjEEal9gqIjJA1z59v82tIXg/Z7KVQgXGTHrMzN
KUAGfQtVfcdNBT2BuDD/gcBK+1N2AcYiXvXJvquHKCAqpfRhu3ig+dPnsSDWcJkN
mVeNDUpPu1npkb0Ct4frvDVvm8KD/G4nMWdTmfsoNCrB44XiE/srfEiYKVO5AAXS
ZBh7+3GKaCetqMPIfQkVyjfgCCNCMCkOpUeYcEUWxhF6LeJAjDTJtC1P2Ncj3Sjv
EXQs9OBuVZq88iICv6CSZZ4LGx9q6hZv58aQaUV/5+6wKjUQpz+MjTiT5uvzyaFF
CXg9tv7Nj8DSjQ6sDdm8NT40R7l95xXvfLzTIuLPUP3W5xrgP3UAh5pougKg8SoI
By+8wUxEGqvFARNXSZ/1ePynhvkGrhDm69Ctpt8dD81Dek/RI0+027akKsnDL/Hp
eHDOlT9vQGsVzTvwoZG+/RsxbQu5mYYLCZ4S4qVtR9hUY7JfwtGeszri2mI6oPAE
jn4kMJ55W6rLUyPJ5pW4DpJ5dmsC1NvrmQwfJ9DgNDVgjW6wjXWBsQkCmhp+aeKq
FsjxeG+B/d2C6j7Byoupw+StiOYAE7RpY5JpYAPIFZr3O4gfKZLeu/sL4Ok76M/U
J9qIxf4/FwYlrlYjTDyvuRq+o7V04igaFbXbdS/IXDhlk6NfekN9iLoMc+d/kpXn
/DSPYBAZC4TuFfK1bQRTYlgLQRSaiFdeboNt21U/6V55aqMAKbnhJKH8ragT7bRI
iKGEFyISX98aLAXpPxDB/06mUMfxPbCuFgDF8eh/lPjc16W3HqyUWZC59/ZHwRX7
DbL4N48rmaITEKcxLoqScj5yUY6RWAMEP2hDdHXFGFg3oOCbTFCkcOaJmnQlj8hj
YVfRaRSx0l9thQwLYh6qjdaneN75DdStbuvRQLouCmD7wZbCW/fmOM0xEPNB3abH
k7FKsu4WNwKuHueoRopNOB+E7xwF7fPk68XVvIpnYox1OGABvkDSnLnpaRJ7iZ5k
SQ7oFM2+v/QLwwApCYnappSuuyktwtwInR5d4v75ctxWm0csfHY4ZV7hfkkIBmXo
JuPpD9Z2j+FfTbd5GfnAHL61nTJiU4mNOueBDx2oEVFkKk5gIgIcpTWPOyj9Bk5/
KWDAplckueInPImaLz1mb2aZKy3tgwT097z1FrCDbsoCVqcvlXilCB5SnAOg2Gv/
vIFr08qNYxp8dLl7EYmeO62/wZbpAgMFpj3FdmIT0tczxx/ZmwC/Og6uCZi/NiXp
n0T1rtHJjE/j2GnJBuRy0jzhiUoga/rlZfPUTgQEqSkzgw3gGeqDPp1dxEP8PvqD
aG3zd2RVrFD6na8iy51FiEP9LgQjTmfbAFEuVYVU4RJ74MpwV8TZRvDGmS3fWq4Y
pi8E/8FTevT0Ee5cqs/VxJc8A+/jseYKgaEanTBsoAnBo/trX0TvwcIWd61tf3M0
4i/eBcrhw+DQLL0Mx9Zy4kTFdHErh4pxv/pD9xlA1vwWB8IM518iI9UK+Pie0IfY
ilza/QxEYic5kWAkTZD7sSgmsK/3c1mwXARbKmYBFeKOlilgwTCV4AtxvAGIrn/w
xwLlnSXzEXgRmkPNM6E4OcZsAbLLxmQYferTdrIuH2lLCZCFIAS54fxAOlKWHieH
Y+yR9dlTuxnjdmD/wP1viM/iYis0sLqkt75CNkBradWvc9Ubpg6bERzXwl50uO6m
sX9n3ferGzA4GmGMnC7NBj3mFZj1ZUL9LXX9H5ta3eWGGW1YsdlSDO4O1AVwZPlU
ivBfs5ZOCTdtTjj1yc0YlOrZsFuEka/rtFwckIyLJ+pUB0db2rRPIGgh/eGmdtZP
HX/nUcqGiYtem8ZzEkwULzG0Licked4Nvkh/klJjRSAasSLD3PhPCI9Ow5LDvOzY
hiIyhoUD42KznaQW/eHep3jaDuD6Wmi7mcbiprcmJ6+CGoExH/nf+P85nZLTA4rr
Z1fG6COUz0kXdmxRXXJlSlkzeLbKJDH/7Pqbu8kpz6OcACceUYqo5765zB375YrC
3wEVVPS3qlXDAm8FiE4zUeivXY4cxVvrqxKPzurjQrdmyInigpPTozkg4IC2JSAy
QEjtBKLTtUpLj8Fz7vi9klwEuWDzzzuYqC8T2UKwxp+OtItYGuhzUnL5s3jyDI62
pgAl3xzX/ZoMYUqpXPFM2KNr1bWlA84rj/ljDR3VZK+5Fmf7aFHGTFkwEuskmYMJ
6TXSIzI3t1UquRWq0V5MSImg/k/XdHaKHYhBnS+ttl9pJAIinEsyvnNfLd7lZ5F+
jwDQeGfgaddkYw2q7bmzFbRLyIkU8X9WBRXS2YTBM18K83JZdiiA8ioUvoHUyyrC
5BIk+Kyi32elxWnVV+ntdc07qdlhcjEnfB1Id0NrT1BfUyEntYWH6evKckUmY98P
/ZJf9QH7ec6/3EKnSkNU1ouXJ8wmKXB3Xe/hsOtKpOE9wk3IasEmxMQppD/ZYqP4
qVZhpdL+bz4bJaAcFD8M6j6ejCVM7e8ilbXWQGOMDDPpSXhSSwrh5OrZkRYI0R0N
8RoWovmI8EZ1x+e9DI8vbMlfaq1LqF4wvQEy23cNrjXVAZfvPBY/RqB7TY4yaU6h
fzRsvErQQsFatlnvkrGJ56IQ1kwZKuL7an9GGI1zcM+RQkwpJhkB6A1cI1va1k6m
Gn2+C8I08KihG46XJareW972GsbScQt6EEF2c3mvFODR0UWuYteYht/KkH/CB8oB
qO50SrFaRXsiU3BFLcm3DWypRftdnpyEg9FQphfxmLa/q/rbnTZiSs3iPq5L0/j/
uYu0EYcuh3c9asUmpkTxU0epY04MrDcdrJM5AgWCrLOPBN/dZuLAOnvcDblLdtuh
aTsZFwUY9a6387sDcq0TsS3NHK9QNX0opPqgWExZ8EkUJTE2ERJYhst0qLxXPzQq
HQIlKW7F5KCRVrlybQpZgthl2+F8Gh/M2JH4OxQ6phXVYFvSXtQg1xdIXokhTBE7
dbtLPZtbghTt3d68qDzEUaobAkyBgNqeYkLBhhw4rJlkeGUFzneSTNGSnpAvhP8u
/gFi9psXqY2e8fhPTVodfzCLJW0tqhSHXJ8DQmetqfq3w72h7YiRRtjxmVJFDeeC
XrerDzDKw8pttRJTDzLrlhRpnkhQGXjK2RWWfrt4V1F2swKJ9D3brG00wt5lWI7o
SxGrNJmB0neCpRx7sR6ceTUdQvwMAhmPHrWsCArrMA49raapj0ehaU03XZ7jUy/B
I6reIt4UpUdptcWMN+EJp85LVdJ9kPGr/7mj335VWRt6+rsi4J1owiUiAofjLKAR
lu+3qqogCZraYSjfJwFtOjJeJCI0UA0EB8avSkywqO4vBjJ4mJqgclLCvVJieHAq
qaS7gAQA3b2uuGwawduZkGarBXralD2Bb+m78e1Z0CwOsCiTWoUmPBNJWcMIqvfh
sGOSo81nhTHp3X1mRCPS+FhxAaGx50MVxhuN1m1YMrv1YQW4fhi30+Ya/wKV9c9t
p4haJAfmmmnLsbwX2LySK9c0Zw2iGgUJqFWMnvRzwXGeVME4Wcp+b3kGWWa/curT
2vZbZ/lJmghIlg0QQoF0BdkSzxMOO92cn7S73WpdPABO5ZKYEsRdmN9bQEcVf/tz
uzSVPxmVclOVrPmpbz+G4ltC8q0KceoVZocszuGV2xdavHL3ZIV9z8/rpb+LK+JS
VIpFXKBB/mKBv9RMUhRMH0QuMwiPpxq+zzxXc9NCOxAeRjsG5tiLPVONCnN+vNaA
E3EMJ8wBr/QI6KYvNBbb3h0OCE0eaEdluQZmzk3Gkvg2JqNpnufVqrD2I5Opr1W7
DeUukFCmCJuCdZxvvKjFnr1tkfs2HDI9ORPrtOAZNxmg+xKfCQL4CShR3RVbmyw8
PkSrh9e0UquQHk0qjxT6hS6YVsg9SvIYCWDL2hKDGJ4k/YyLvo685KNPx3yhYgXU
tl4IrIe10w2HLR9//RasPLpk+1drqvGK2dPHb6SQDykdJ8P6apjOAOff/iYkn8gD
zIgsLaUYxOc2vDLwk5LsLvuq4HV0ZQ9HU0eD0g71O+F7hCzQSIkO+AZufvqGzxIm
WyU23jVfsnXYV4x90iL6p+SUmsUIT+QE1J5QoBAHjlR68/TYlR5F5TDEYlbc09Gs
Yhv46Q1ABersUn4q1aq7Sn1trKU3lBwO1rdjSc+0tnBpOVDQkmt8a3WsslqFLwJT
TY7d0qZoAtOGPr7uDt18b2dVp7+gPRBmwXIfotJZXQMSdWadbi6+5lKqug0gh0An
8Gm9T9XaQx8eII3Vkkirrl9eMg0rokAM4/BFLTIK9+UdGeATea2c3LzQrhRNXL1R
9CENiECD1TW7MbnLnodYfyO0huRlDfWghjalG6EVM8HaHCvfFdFgQF9j3z4BI2HC
R5pRdgmgF/fpUySwJgu4oElxxek5Y1l8n4tLydqEqZumcTKS5iyj3SNiVyF5xDqj
H+sk4f6hBQt2sW3PBxWDLwV56iKWo5DETB//VmpkX/o0sVKUYMPlokXL0WgAJ2nb
26bt4Ge8nlMmtu6iFM9qmq5I+SKET4ePmt0BJdNA2wF0D7++quLJdoZK14HeYLsR
+zAQz6ho8D5Bvw+g3vBYW+opnJhEIc0JkbHWdOvwXmaEuiTzaK4Io2f0L4kK9DPS
Nr+vjFdgVuh14kFLISx4dfXDl3XpT1GMu2lC3JpzCpfuMvG/aV18bqNT9LjjNCo4
IJJsBRTRNVtglT26iRvOtnG1CV9WKBuktXCQt/DVpnA9n3OhjOhXb6prdsU/uMWq
dwhj1G4y+CGWCbue86PfFHGmDVornowVLUN67iEF0qFVrTgV0tJcnerG5pVd2C7f
V9jU3KsgBVj/tik7PsIlnS79CLC26TClitkiA55F9311qnBkmKrlpySLPQMrjEe1
7J9x1NBUQjimDgvL1X69DK+E38SIkQuPlAOLycwp+T9ZKc1UsH2Ua5287vc6bmGO
kzK5IXQducuxS2xYQqWYtMsT/KQnNFpB3jHPiQoDePGJ7pwWfD4Bgbg86y23480j
ozl/8KmaOyyVpSWUOuOUDfbDEij98Z0dcOxy0KCGBooqwa/JlF0y/BN39W4ck+fE
u6Yc0jVxjMuK3PdCyj8Zq/ASW3WtxvXkG5nh+5F/FU+uFgBkxrdkPpy0I4enX9/D
RaCBGof6iWxFLxRG3T4SVt9tk5pIDBEZsTUKXIQU3sdLK+vB5P2ZUb3JIQ20+04u
4Ab5tVPHRIsiCuGzJEEMZNrvyEw/Z4LMMAtR+6fTAyrWRcXGNmh1MbBF+hLEbrPI
N/eRGIGo/4QeQm7VS/i47OUMyMjvD9lPKs3vL81JuI1N9C1Z55hXtQzQM/0Ove3C
YlZWEia6O4HlKtNuU4+7N0Enzwfyd694Ph7Rip2XFSA+FVfkcmr/E+TBFq7jLcTm
PC01Z9LOKFI1nkJLIq69H4m6BnVvshsEBOh15eGuRQMYNl11oiu5O+8FHu2HFSpH
G7WdxN/z9K6C65hHzHGegBW+vuqgalgJWeRRw0CZEU2yPm8RY0+HjHryXLw3u6eF
upL0WTaXJJ736vXwNBMVhTXHBPoJ8hCLm5H7tYtWzDdBKOEl1ljSvUibOZKxymQ+
idUnPsR9OLqyEZ62L4nmiYy6vIvCBrB8niNenGZaTbZlKICeDOUOsipGxfaWFb61
aH9KBjjJ16pPWO0xGJDKsgd6PPnL1Vo5xpMg6wjfhslYCkeQF4uJpLXHRnuM/Onq
50sgGK1iuxY8GPOC6YE08lEq4e0miNC8FBJaSe9BhlFBXvKBROv140+n8WhlFJU1
NtSHp0AV6MtiAOuVdrNAUpVMlog+BityJc4mBYDqdZcaTqTXe+PLLF3lGSp+WAGC
OfMjA8m90tlET1XlpewflHGGfczcCMdbhOZSHzeqWcPt3Y7Z/Z/sGAgWRnxBcpWt
LecDQAFYwZLH4ExD8ol3cnzodJ/MJeRT7BvnDwN+aGfuVgvfniUoBaYAOOiHvTfA
SeS3fQMOf5fYfmNx3qxirvs4MWxO6Z9QF7x+2xmLyaNMzy1x7O85fruyfGpHeeUO
geffOxjTAh7jWTj9j1zzx+rxVdHDr7ThEnbjyvMP6KZlU0qaCxrNe1WthEsO/XCu
Xr5kNiIqsbe/VjNdMA7jkCHg1wBtPtGPJRXW/gVza9fcx/l+0Z81/gCdo2B/iVna
44eJvFm+13NHKjO9o7OMueiyDQ/iQ+ORdap7GMlgT5oGwVVUKA0cNeKvemzpTqYL
pI/a1qtqsqBtd13sRUIX2d4t9T/2M13fNWrLE7dxgyOjoQ1y3QZoPhBtDG+BnmKN
WN0Tq9BzbjDuJvhy+ju53We0CMuvCZX8k/5nPpLTrKAVXx8QePNT98AI9SCee1+1
glDHzCavLsyxWZpv6ON0VIdDSXem0AHiLEdADkXFCWuqEpntOkA6nITppe/mfsnl
GRVt3+yl/pj3D6nv8dODq2acMEGGLK9RXIrWX6vNP4sb2tQdt3WhbZo4m2NNshoJ
CQiW/PCGjy/ibmD2f/jt/8YcTmCYwCPUWyIWGLOfhmu0dPeIm86QjUGcEgG44Cf1
GF/HE4xh3+hANkMfnLIu2ndDenDRkSyd+DArb9UypOVxZY60/N88uh0kme61UHjj
XGc2GtP/BdSFPcOe1PQAYlLuL2HsKjVUJgMWuLJxvjHmROh0wes8yFOBfKvNZtlX
+UR2gjRNS+od4X2H3K+bPECaFIn5mYRTg/4BmG+IHXXEvFbuxnnXyYuEhsEMRKpj
5jAyKyHAOjCOivH/xrretDN4yfQIQNPw+bGvmNnympFXEowCVIOWzHLqyGWgVMqQ
TD5YX+CztqHKjt9DY0i3awi0zaRA56yMW2y6hTcSd5DM/2IXR5zBwqNblCn3PAxi
B0NQWBQxeV8qLQ5dppIXoCtH50WZQJUOcJCyf3iS9b5pUhr/UJwiw+Ar94p7Ew8n
a3NOrdQ5x2Kjlc67s2y9VD6G6he7YNc4obNfMbNM8orf9pWLU5YUb8wnD6MTdl1G
Csuu5Bd8sG4gtVavGwlKCtNe3JsXFSzmMj+cwtrVKX5ceFZYK4keZDFsQlE7/Cz4
ISc7K/1W2M+QRAiLpVzlV1OP+3SODXTqOBjA7Lf6d3J8Ub1BgIyMFMAg41eu2yu2
GVOw8b4ktrssS5jsbNc4th2JGgKT+Sh/UTO5XX4+sk8OtkepqLyXFk5VMvPjdVuI
KRh/wVlBewJFkeDUHT5GGqvYD50JLxc8sv84lMFmOz7YpFv6t/7E/dOuDAFODoh/
TuSJjxuTcM3pZ2eAlOrcIkPxRMSVH4mbCg/gUefmrlqPVq3YEqZfnZQ/plhbK2bQ
rrbwmYKFthKZ5R0W1j9rPc7IBd2Ta2ofSA3335UhhC04sP3JLLS7yqE9S/vAGJkr
tWaZUhztiZxoZjV6WWFoZnRqtsrNDyhdgezX1BJIOroid3gBjckMXYBUdpJQ4fBU
N9GjbTN8ymRfZIHXfgGTTE9+IqB7tsYSgZ5aZaBilYdBAl1zw1rp6KTIgcH3WrOg
yJuMniuuJ6VcvJi50E3kdrgXsBCZUNFOi8gMAIYH4sZvZU7lrJ3Uf4odZe/aPlxM
X/JUJVhq3F3JhLaHQzHQ0nZNk39RPNFjIjcaOtnWjfBsVfamdBw7/3aeKLKrNspP
MExGaCO6xUWVyDzsp3D/oEzS9Bv7zp4UEHchZhQXWgG5bqnI5terJXPkrSyE5Sex
bHQ5tKSLWNqYLKF9WnZCDM9JkNglDY4MTcPEZn+GU0kZpXrOAb1j00dcJAW/MubG
2z0LW2DOpfxcY84VvPgtfuQ1yF9Kxd9MWjSHC3lt+Paw3BG//6vhK9+Q+1wBk1ff
dBSFHPos0h4bRLU1de1Zk48KUpj/BJJ1b6phU8JBzW92V77lvC8y6YiR+x2xqlao
mV9srD41biEJDG1dBD7mIEurThD+2y9nm7b8b2DMq1LFZScmlOfDgAjvaBaRyi93
OJWN9sZRJAmUVP6hZjG8Hmm70Xc+R9m6nftym97IRK3RvThr3GRw4BI3kdEBJLzc
hRxgbwI/+Yc7eCMN2pLCW5otIdalCEescRnv45m4IAJ7a/y2x8NCMMAn18CzjKsY
dLSBpXP6VquVsUTAqKsRmQL2s7XdbtlFUE13/HteA1yJGjVAhCQoNzuLtPQSjPJM
7Mo2vmbeVIF7uzjBryPbv1TUkLNijKTIevUIgY0n46Ywy6zaLgQEbY/ds2j+OviY
lNNb6MDfnaw409NSD55ezUY6O3imkBtB1o1UVwtiJKQt/a7/rKI4Twe2eMkHsj/G
FncgF2VX5dfX3MTqStm2NLXoNGVXZMX2sE7hz235z+JlR1UyeNl4fiGaUw3qf6d4
OyFhM52wOFqcC6f5gAY8yYLNxyG5DCMQ6Kh0AaUWcNnIqW4Kl7bR4QSldmhLbXWe
7apMSiva2loGbB8JGxQD/9RgbpfvemVi2/1wxNKFm6M9xEzQ3QlTgGES0TsrEN3G
IE7s6nvOZK0QcsLQbbU/vVTVu9wjPw+bxbYocP1jNobOCuyXyRXgXvQVeRKbY423
BSegFHtUqy0ThHteHPetxJewxrYPSseylXO/J7DkkygEkqkEGJDHpFfg/PFopCZR
iUd9pICxnLhB3dqeNxxN2nNoZd8s9n30qt8i9X+7ohFIFjPE0kMRR7iO3rMYVD5S
L2azKgrdizeq5Ye68NDO9hhmV2ZQqHZW6hZa1Zw6SiyGqb7oivlA8rFT7c9Pv1wv
7aIn1rpMumdK+VS/6S7giFFEmD5TF1mMqNGb3kT05Jjrc1yXRhNOMRt1dOQ9ne9W
9pHgPwDh2RZMOrIW2W1eCJcLsmfFBgKkV6Qyq0nzh+/nFCcx3MQt49qUbkGRr72K
QfYGdYjfmtEhBYt/5IxhOurYDxbXtzCKGQCpE/ABY4Hpv/L1pT8MEg38W7iPHU6R
1L98fipg2fZckMpejUTuPDzboxPxk5j3ZfTb242/g/7soox9L90cKhrKe48r8TeC
ZUVXYYmXL7KYpozhpa7TbiYjbrwv8QXNgTaM/zI4zNU9XdPqH9REsKAZ7iUPsw7Z
0CypEAPYSGTAFtjNYwIw73oFwV5SVv0a0hRVxHYlCiDPSrF4ETwpaxnV4dCLxaYi
GOyphY/KCjKVkfMuIcoptYO0mHgpVmwV/JF7gQvhxa07Oqe1aPlOt0mXj0LdwO4R
6usFzhkX7ZPGKtF/I+49XJAx2hxL4L4CL97JUhQolR0uAwfYLu7Gv+H13HAYfRXg
Qxutr6erfsLR7apz4kUBJtUtD2YJhUPPhq5GiLvzdsxjbw5Fn22soXsjKF95dxaJ
+GrmYZXGjsbDW8VEegqMvQGjevASTJiPHNXPyfu4Yz8kAgQhk8ASTJ3/O/hiL6rt
QR94hRrNXs5ZBa/SQi4ST+XJaIM65GXSIDdotSFPybD134O4Gyotm+Kf6DHcisbu
ZK/y3F3MaCsJndDHiGzjBMJDjuHA2h8WPOz1mmXbkK1L/P/y2dHi2HsfZp5ANaLD
igW0lYeAuYfqbYc60y2RBDZWxUKgTTTfPeJiADfK2j88fWRSXb/PADtS1KxUrZAg
viaOO7vTp6GCStzkQVq/UQsHfR2Ji4qNSVADiy2c1IYRdh0XEiRmrp7bHjDf4mMl
+7ljCoStWshOHQDAe2EErWLEJ1N5VjABLa8yGJve6zWRMD+tZCFAfTjuoxO3RolV
6UdIxiUHmA4cEju1dRFE9TkCv2FMx3/L58XrO3IDJjn9vyGNUl+U++7u7Sjw0pjr
tUYQcuuWS+zwE+wcaz4uWWnKv6MlZGW5VkrEObhywSq9TAuAD6Z7oeiDSLbKPboI
yWofqGYORDSylFyVuJJYT1eqrN5GswMhQoVzoMh11nF+jx0+U9foV00TTt0LJkfq
+l9dPWxPWNNSr+E/O+9zC5IXIS/56B5fd2cMB2tk13bsAS+AOcLnMLxPEKCKpANZ
S/avSUhTVgPZ4oRNixa3fu8O8x+nFi1FBRYdehpk0bTKA48KkLzURa9HAXokW6LT
VpYhH7B8Fu1Bm8TrsoCRThfCXjZPEo2n/iAWUkNa113CpsiuQ5dDdVMexwziOwyD
wsBf9I1R11G1H8yeri2EEBLAurR8heGHG4g5LncVZRj00oWbxUkOkknqIhJxbdQa
sjUshtxCjejjXdwi/r45DRJDJ0Oj/2a58RKvarmVawz/7ZI+DNWrrRmSR82t6bQ/
JMaFVvdyW3UEt8HW0IunHFQ1C7SvApFW7iMZJjx17/ovDGRNflKlOZZEGf/fpQLg
e28QjMLZl0uxd8OR73fOsqOe4i6Rt8ytncrutVlg7WXHyBzNUB2lQI3p9oA8sD0U
pLQIkj+zOTjNoMifKiaq5h5Mxd02utbp7PehksZT+cps4ctnIbdYrwawJZ0LpxxI
FXuVv1Vj8itT4DLp0E9bK1uv//vkTgBdbEwCNgYY9se7K1fr+tS7siyMSNxGR5aE
kr28pnMiT5rkph6VOI7MnWeESGKq2ZKNcutUF6VMilHZ5GaXXkkzzl/1bD6RQMIt
+OKR5fD0QDbIQBu7YZMREaCqq2QYcwJB8KyQCa0OmEsWDZI7s+3pG3Q9w64RDBkl
W0kZbBX5VnuMZ+/lWevE0RwWMhblA8tZ3mQAviyyeLMHRh4lLb9K+219ZRx21kW6
35r7GeuCS/sXE8eMlERCBfPqK2L31rrMHYAkYgLLrIhIBwpIAD5hv92by4y+Ajou
nRJv/AwHXbKwRpenOCnYcDtTq8RBMLeNqXtTbCIMyK5UDHav4Ia48uKSdpDF+yRw
OFt1izkrsb9V38w372iMRkM71xavyMAJ+giUx6qB8WsrrTHFD/14m97RGO8NH0Rx
eoPMwAqdhTIx1SJuA9BN87yX6wLQ1DS61aCDiVdNjeG6/95hSFky2hcwujTjd2QT
zXl2wU3jezjBysT+ATM6qnthg0M3Zd/L9sWQgs07LTgHAl4wIXHJRI44VR/qam8B
F3KRukLQGCRhQpMKQudWEK1A6Vg4nqWWeBCcOVdpZzL5neOiv01mZlyrjlXuhhYe
GYYY9zV2tSEqh0qAEDAkUou6WdedD2m6ySDBfhT/nIGqRC8dkR/hSMFfsou20fpU
nmmnO6I/yz2xVYmWqwHu4XJ+SCPANxlP/1Moko48cy6KLRXAE01uJZSuBPp3MmQT
tBhk3K4mvswChKoYWdFHun4bXMuiM5XD7Iddt8SN4/tWYtr1JRhJYyUXdv06tRGo
tTEfofumtLAB0B8be2+2/GljqULCYkVrod6+BUVMOXdDOm0Nu//MoLOzkSXZ0Wws
3GedImBUZCxCU+MxJS0sGh1TpNpWAIAVbydleYh8UA3NaajKad7gr0/Kn01dUxxh
rfdCyrUhic2V6drKNn8EQ3nL0GCyMzgMvevyxpi7n9tkTrqoucnmJAcBz1YR8BZr
Wrc78bqqjdfFzPXqVdSSGd1khEtiwB10PHCxwL8WDzYGuSzghf4e4IzVmpW1/2Ym
PKFGpCunhOmRDJRNOxGfWaMom/m1OHr7E4pcebtS14Oi+CNBQmF2b028HX43n37u
qC8UGX1K6Q8i/Mco+iI/K8w8nAvMv1Uy3/wi051zCAgg0bZLX8rCG5eUwSicZ11R
QxhIDFhLXDgB+yZiaDU2yW6nk1HG0m7+SlLc4WxM5+1/axxwrsrPQPnb6mfm6BT7
cxbqiofwIVn24vyMSOfhx34CtmxAg0joQ7JqNrcd9EBO6oxYY+HgL9uWHvqtF6Uh
sYX2FYp1TpAiEaAnUjPIPSJaj/Hx7EfhzREjHjXUDUfayEPqCiwmLi2U10hx9pp/
A0dyF2UzG2yzcwVXE//4cGgwZ1oR+O4dvlpfn9o2t6XRjI3dmiBFhWFGDg6OBLDW
67dHgI32MJ+HHBzwHQdAFX0Iv+iCvMS74mSHSeg9+g0d2/hly7MYE10ouRG/GPt9
OwMLrR7oo25WFiNRZ3eu1G8wViWh5+faR1fupCnWcJ3dCf25T0KiXy4qkt5UkUXs
IbchWDLQBUK9Z/XcyhyK8Z5VgcGBf+iToZvUWZjEMyQVwvQ2Z70qPz+o51QrwhyB
l8irCCaeKdTPWjsYLFR1ixyVHk49KQn2tvYFD6KxhQ6y6pwJow+PfgCTFo9OgV2F
Zf5IElDtdOvG97Rhs65iAqJ5GuuUz6Ti4FJXG1jh6JhDAeOoOdc6bFWOB7Cqx8ld
P4/mLOq7BjuPnoGEdPxMJoDqXQn2dPlYm5+ZlUSHycTNYllCvmd/TWPD70dctIr0
wtGBukjoONwZlTG0uTxaPy2KwkX1Vo+ZHRYPfrp5rboQ6g4PKt7QADzwGA0kBMxN
ciiUZYeSleqdeQ2DY+lK2PF/SHdBnAh1hT9gd8ZhaSOBgRooLT+LfOpCJln5gVtq
LNE3IAQ5DOG2LXBlm0wjawz886OxqehqJzPfTLry0fy7VIUBygJsnilLkLHihHIW
fv/74K7VcU9K2+jjl25NhA+8FzEMTeq8iCScP9rA2jype1xaqRI0ZFoojvupFnOL
tmkyKDjVdDYzCD+WoyRtLQ8rChl7uqZ1E2JcPtHPlc/5RLJYXtS/NrgMv7dCMl/T
GOQrifTxx7bgkFeOUSyCTpAioRuEjHqAL32zAilHgKKQffZQWgN0PbPUm4PY87p9
0aK+kUM5XvnfnU+C/P3EqrGLb2pN3c24SfEplpDthKIEvJvfOHbt7AE1Y2p/LgJY
fgQ0KgFR9wAwFbfg5qSvfgh/NOE1xVENN8MNSO3Ie++Rwca7hOuxkWTn9lc1nJmZ
I77+CI5N4LuHoRjlKrONxgK+x5X4aolw2YcnKttZ7RlHMQCOzFboMjUw9Ku2qiAW
TqTbd1LiIa25DZBu//NoiiWSb8By4qf3HAzunQUxe8aBRvttiAdSZaJDAigXhRT3
kQYTwVXu7Uk56fHKjjwbZdUro+0MId+MIeBc/wpVsQJydjUXPAFBDpwoZ1nF9wmc
9xW6fHlm+BjAOSBVvfAMQpdilrLvKTpgaxIwtG0tIbqrPJk+5ydS5LOrayMteNq/
ZZj6lbq5qpj1DhkIMbXEqViuDTi4JIyWDYSqLSpqEtny6Ho1+AAD6UNfhhMD08JW
lJai3iNUqP7F0V3LmYIh5FLK0qh9UBVUPWlDzekQjo7IGV09N7Z0xioaBqEtM/TA
iF3u00rgvrzYt+sFlgrM4JjeDdZXGe//DYQfDxOWfHA9Vhv0MAB+Jf+3CkB1D7Qz
vimUMnbUi0f6E6XikH8xdscwLr8gtPYVwu0tw6aZ6PZHTnwxvOsW/imwypsalpCI
g8tzeKaJk+rBGxHlWCOagQ4s42uQS+Hn7LYdAutzb2x1OWuh8p1zkX3XSAurR8c+
YK7oAagDqFFgxI8/Pr1gLX1FeVqJ//+QlPP3jzc9fCESacveK6pybxwkU7gOyLyV
V+STB3zdBzbgky3YJ9KWeEiwabxztDlOzb2zTcBTWffkOGqJWTfHNqS3Xyr4LdXn
o7D7ooeDXETuSjMitxXCBszrRHCyHVUa9GtTMSPsv0KBOk1wKklBGcG7MBPBFXqd
lwRL4zA1JbG3T8f3Ph3T3ae6Les22SDuyxa4Tc4hJXlYrJJvd+qj7AZKdCtXrJpw
IXAq2WcrNoJDLeVMhxmGMpU7ZTPe7sMZ6Gqe3nJJYS+40rZjK5IOtkoD5OgQPQOT
9VXRsZmiS2jhUGMDOdupRzt4ohozVWCE2GF/zS5uxqzyYU7AN97tKzyFD4p33PES
BpOabRBKsi/Nt46S1rd/mRCd+eTNEW93xuGIkR4PXdAMIVjPrLmnri3anPSZMiQw
gcaQ3DHF+t3dIqjuYiHgNJg9H8qxv2BfmN44mdZnhe0QyxwoXJEGJRDsK52Y35Gl
uicjTP+W95M5f5bkx4i8OPT+U0jDCSCyULIvGj76VLLHUbXA/56UY752e0XGxbdn
fIft0o9/66mZTc9VkHty4MgPImZ+URl7OjbxVlyT3K3L+s+WZMrbSppgurRnL1Co
DTAth7V7zqAo7Yja4MqUttweUxfYPO/yPNXAI11G8Pr6h/HQ3McCF/RzUW3I3OQn
t0pI7qi9e0t/Vpe3jGjtVDgku2BqsKNg2E+sHWnin+W0aXdv5wi3iH13k4Lr9oSX
6WsLRUgiI36EvKeHF3qCjyFqGgSX5A8xtZGtNrNrC3Qu8WtuWv3oKT9Y2mQ+xPHV
+6kZ1hUB666iscV57gkFFf8YZ5cQczymp8Gv038t/Gqwqqopo4HcGfTec0DtGSH0
ZRBAZfK5L0bPf6aj+hTBcLn7Q3aT/8Zr1Vp/wsGfNCjoTg+mJod/q1v1wU/czvWe
DsH7l59WLh5cggmnkUlAPV8sm1ERBFFz+XmOX9dR49ZnDhIkXekFYV/2Rrp6bM3r
u5uJk1KOfy4e/Cmzkbze2C8ZvI4fhEe32qOXJ1zKjIerC0Qt5qxc876x/7w0oMfm
PhlRxtlANt8/4IjT+2w+VpWiB62W5n/OUeYgJXqVuv3cuOP8U4vWrr3U3TGGyAAg
GYhOtbX83Gpm1fh4ysmgt5ACwYBXe/11vzt9P3zXSX2V7/oUpj/oDMI1qbUy7cqS
HhRm1B74mN+oEw0KEGg09ogdIIHIc6AB66ISlZS7FzV/Ty15Ijnnp1pONUXRmS6x
YiYfGDDPzK6BVZNWgACBVFu9kiwlQVMxQjHi8yxRPcJ28gHqAF8Ux5mqPF2f960n
xXIf9w4yaYA6RNYF920Ei1CdGMz2YG81lmvUxy4/maACQUFjw3dksRyaSDAxuQ9K
5ZRJNIpKtBtVHXekYOWtD8I+Fro+IZQED77FZoI6Nbv4MyyjWGx6OX6K7zGH9ZB8
hyjzMGo5s7rgCTpYxqPFEdfUDO1GsEzXk0GkJZDoJ9vKszMCO2wuWs8sZyq1euGk
uYAAoPyuQTc4zzbWWADOY6p+wFPMGzALplquAd9wf9jKNdVkIDderllpW8SvCnEO
KZevI+iO6D0VJQySpD/304giJPJLLxpu6L3aKcYsXztAJhNnThpSyr82/gmne4lo
iVRRpQoS1vti4kQolBvCLbTqdoJpVmWM1ojZKBjH0bIuQTSb73JeNlFxU5hUYNef
uDPnTgeIBi/V2cH4FTJOHUMwEYrAm5rBD1IWLYNODxLepk1JILk6jEyuj9aaXfN1
2AN3e6y0+XnLmu72Z39hoUxvC9uqP1PFzzfZerzxBP1J5GSoPyybp0eM7NzrFBHT
X9Pfcg6E8TU3Z92UTi7Q4asMa6O1zv40iUBq2A5A6J4p8ZYlq3CIC3z4Ms8XzuEF
+9b6LMS3R1SpRTEqS+HTflxRp+fJQRU5D/bPxS7K8f2jNFxzCUXrs3YPhPfWBifo
ue+PigOPkSHLhr/QYos1z6pvJEP8xmN4aWqndetjUTKP84aqg4/Tb6yA3F5SxNem
jTsRh+C3fMU9WoF7kN3WONwwsHl3ftG+CuR962VwyaliQ8eCgH0ijchhULhhuHGt
UT3WdhGT4RVCLxW/dOIBEBO3aPJwE7osUeL2TCPiyngWpeDxQV87LPQBxAUh9ZzR
0sOtH5dzRNwuMmtANPMUnyDwG15/VzENd2s3uFRp2FLIGEcLbBibWApKQMhoUo+m
NiqS+n6Xqar+U9WRHUjRwHiiNM3UDtXWz+xHf4q4mdslB/dCFCc/hS3uSnwg3Dvj
hdOaIGUvT5zBTTqdBkhH2WfjLjwhSBEwlg71wTqZ4SYz23XOwsoyuOGFCkXokRtf
W4AmvhLwR20cYWa7GgnJsRjGlr/7qdI2D6xcRfgske21X+OGV3vQNWSSUrKfedeQ
bmX5KVkRNv1GTd8UYfappD+EKNUaUkHu3mUn2au+ZnupjXp1ex+SuoLa44MYDdmN
WyfUxI7v60wn25LeuD79AgYa0qzR6nfMaG7Qd/f9RXGeHT3I7BsL8ia76g6kW66p
TsXJSfocgk/4wa9h4oXx1KoS6rH73udkN2yh33NiwsPvW2JxaelpY/fNsDnsoeZ6
2Kshwq+cwJ7D8I+nPe87owTci0nEA9gk8Qd8kGfM3fHPonCqIQphYQyEb5mIJWoi
FYUnUpv3NgaAc1k57tREhsV9a2ESzHCg+M8H15T9oFDZnEH/OnDX8uIIk4ZSlqpL
C3c5DwSA5KrwnBll8rFm0ydzvuWAIuHpo8IditX8IDzIAKTSFGYRDDryLowf1L72
OqDdr8WrTwyZ0dHifeOU5WGKAOmVbhB29VsIyzPbGiYJDPOc3zX0WaqS8CyK+jjl
Ub1fCt1MKuN3zAEctyZq20dw/d/MVhHBXUY/aSA/CdvUvZcq43RM+3enWkau338I
3RCIfgXt4uRIAuuhG4Wx4S3JBQMDR78vywE8+4ZEpWiZD2+7qyeg90lmH9nVBCDp
FD/8gHKaRroMYpmgf36CI5gKAmZh/Xa41I/u+fIvsyfLyeMTtMqtNCiEbc9+RcQW
OAytJMdgQrVYHZPcRgoklgWWFlK7YkVvJaRUX/n+IB2Qxni1ZJeD0VlFLU1ipdwr
tks0qcnOJG2ojFxwLm8pT/GxGMDGBFTl7xTrx73255vUS/s1llPLNVUxtSbkSJmk
8rJRMMs+6mnBOxrIm7xwjN3WKXVrlMzmaKAKjaRHVpiG0JqRpFCE53LE6rD4o2Ke
JvwziBEHesZ+i1J6ODukb8k7G3ymHPtc1YfWd7QjGyO7IDcKBfHloZPJHJ1xAvQJ
nmz72p5L2fCv6PGh5SGS7487hRrCg/9gTcJzLTYUAytwyT/fJdlSQCRLLDKHoyEo
ymCWgK7CPNEyhqRLLNYhtn+8rgwszFKvCf6kcBmPSCT3s8coXsZUAghJzO0SlihA
51Hl0MS2ilezNdZtJqVJ66rQ7BsvUkjBHxfSVM/CAbyyaZxYFlPks2pLm1fO5gIO
TcauWfTikLTpvQ5LcuGlmkGs9rL7gj509xl69rxGSVPRsk9o7s8M5qxqdzF13qDF
OmFxIPN+rUB1aS1LJS9833mBUx2keKpR3Xqcdr2oRaTISGVWbipnCPW/AjpvXfYP
xvBWQMf41j/nWh50He7jE/rprRBf8KVUb2pzAeb7CTO2b8WllQ5sw1amvvmtUD4h
dS5Yusf4zI5494hKoJygHf4wvBgZDmy4cMX3NRD+MgGwaIdrM4m20yD0l1IfyUXF
zslBVMV8ipfcbExr8/6zZ+ObYKvg5z3bOV6n7LDwNpgxv0gab/RL8clq9T1xyAap
n/Gum42XaZnalfVDKdmadsSeICmfahGI6DaQMAZujH8Cs5MSjafmiQqOXsppB2Ty
6Kc6srx8HU828VKR9FurWP5Uh0RTb2n1bjR4nLE3jlmKiS2BNvcUiwmhU+tywHxe
+aZLlnTYVXeTC3Ihh4Qf+PdIkxd0nOWO2+hVX+A52S1ySKpdLd86jJFfvqt6BC6m
fvSYOjxSRq9wnS8qEkJuUHPypV/Fc/f/s77p5PIHPI/hu63jMmxlocAG/AxpDVZE
7TfW8rk9iH6yDdebGjWGprRauuYCTtDou3zR4rERNNHcB2ZYhlCxxepdbMQ4riZC
4OsL+edrG2/0oYhI9pPCEh6eTUq8155nEKtQxey3nrWC5yhGnoeNa5O/O328lxgv
0Z1mIAajnUe4T58Ao5o0KF5licnmHGbHv9KBgTjXAaiDgUgv3zcfDIZNytLjf8jS
6cFNXjvfsY6HiO/Szz8o9NaYxYtFg3bODHJTnTXw00OaID9fSYvXh7BAJ3FoCaVl
tOrl4qHELZBs48mXOwNvWnPDCwOG4jBxExcUBvaLGhgcENTZuJAueC5fH+SN+GJa
gHPhcaAupQL4T51kDgQwwkPiPATEq4EhArAd3fN/ICuj7s1k6gxCxayiO3Vzfo1m
Qf/bczOTvMuDKPylW6q/Tjwi9gaX7/0kZO+5nVAKp1NFu1QFDpv1F8uVATSPUh7+
YBFFO6IR7b7fSkdqWkazBT25NeouuUj8HV9Q8fxkP4QsspD3t+FVRjucekMiZwv9
xxS+j6if10BbFXiiQkxpZsUPh+jw5N9mL2Ou+Hd0F/KNXDW6lVYEdebqQkxE8t4u
o4im5sAM+wbOCAFggFY05/otUTw6GWzMSRLy1HEO9tXYHcH2PCyplcF6XsXakMhf
apKW83iDKlqQmhjhtMhATpNUQM81lkAnfvKmNpN+ytbDoCxH1i7u1GMg07ltPoCp
NY/rA7CqY0RYJ+/TBJhvy8J0UN1M4Pu55yInuJRkH0WA0cj47HQgQnn8mUviMxB9
TM4eUZRJYf38EpuGV+MyzwJkalmkNuXgCNJ2yOOsWO5yweL7wn2TV++hqftfhowt
n1/x0oNGJWhTW5HqP24ZU8B/CzaABhZIFEvzDEJyNMsSe+PcBWAV+6nCR8mcgj1k
DvXVDwcFYrW1bGS1q8OdKjH3SBsDsUk7jWe7XcdwQl6IsCRXv0TmdabkYrhgvHoF
91ZF+4aNHet6tKHt/r69JzXc9Of3WKwOGjvq/+f4Y/Todeyft0NUg8IpDmj4h5X5
OfDxkthzyEeZBwMJKwv/+GqlpnrfUUZIXfb10UQSS9zRcyM4qC6wJbG89x8rEvmi
hTp21/KmD93Cx6iV3sRDqVTC3Zwfub5Z1C8/JD8uDxBZd81qtDbiYWMi/7UALpMx
rNCFE3huee5gxhmRpGRrUF1u3w0/H1XDxo33lux9R9iSqY7ZQnZgK9bqGT67s0d7
7ptwenz7IPYH6Z5NPI24GV60gEW2Dhww30hs/ocq0Ui3aYAJODna17qFQ2iARm2K
0pjFEIJtx5yqgV/8/2v0JnypUiQV1dvHhOsPGm8eCkncZkRO6hSAzYUe7ZIdAW2I
HUXyZICwSxbOphBph9DvYs4UAkH7xvjdyYaw1Y0vtVm9OLdMMH67SBkAKa19pCit
1UTuFWhQaeJIc4Gf00604LMMpoCOFjnziE0Tf1k8yVY8Jr07NAbzHeoeCzjBd6N0
AMNQNaW543MuPFx7zy6z45OXlLnLMoJPJ8dTiuGOslZHWrMCFlI1XAivvfg0TnI0
kmJ1B6SmAfm1zknUBRxVS6pSKp3j4oHSsPgFG5sxCzbKMQ5II3W2Tp2yf8tI2gtM
ptAWa3rgJawDBe/BdAjjZbm3Lf3vKNWv0BpUUcauqo2Ylu1RxeHD/Dio79m41gOB
G9nurZU7xsBMZ9hZI1SGYxjCqlxeXgOFQ/U1uREZFYUyr111zXazYX9XJo8zisFa
JtQBpKML76gt2rAHXYRcN2/KYnWjL6+dwoziBZh637eTUq5rw1NgFgxIDaV6GLtz
ua26UDzpvq4NFgoo6awuNnQtEGzP+3aDW2XFafa7Z9WF9mVvuhcPk7zWG7Bxp75V
Wbi8DHcNEKSq2FYjKlLL8yhiLv87D1jkPC1Jikpv9MHMgknm5ftuxyD7IYWP9nNp
zO/p8a0vO1oyfDUgx/SPMQ5g8gbzLzgIoH8Win5xxlxQ16Euo3Ce82EYvK1p1h+C
EA4XOzyBjvbZur8NvZFWkgqZ1f25W9qyNldIA/0rnBVoR0udxmaETmwZoqEb+b3s
dgJmiwVziW7EylaHAWaG0yMk2+b0Gp3nkMURXcJONqx1X7Av5n2nR5lbDQaohC8e
nwExpC14/3do0BSnZnVOuxlXo9W/rWfPeHRK8TSZweW9fm94Aw8dmu+w8hep/fFx
b30ZoP0/Jiglw/eM8pdUpvr7Onx8gIXq8bm8I+23UXz7prA7dGd0/XhkEMPIKJy4
msjqT88pg7EE/PoVSthVEdXw6L4oWdFp2zefBm/ZW7ZsTwh3CEBAcUYHgQuJorO0
5zYGhZaFaXpFV4PfN3TzStRVwrzoDmadCOqSYUsENiQMR2LuSn82uvr2j//66HX9
1XJiryBldr8+z3xWNHiyv0xd51y8FX6LjV1VorY9/2lnNXRLW5Ee0tElfaz+DY9F
mmJJJb3WPAQJH1I8XRUvKzieNcyMjwyA+UgCD7YsJzORVAdMGm8c5OiVoKJr0K1i
JKedRbmms1Hr4g2jjIFGaJ/GXJh7HsCPqm9QNQcbLm7Ogbe3otYp72sFPycBixE9
P7gAaiAH/EtnN78JlpwqPICN8HJsbZFRCppqJ5VB7W5pNoGlPPD4fcN7bbPM/HWT
4FjGBSDW4EBa5fKqCFzkAV+l5tTufa7zte7teIWsPa37QJAMLrPq6H09J6YJJDl1
jQOjw1dAspMxWiql1TSNk6HdM1+bCwDBAbha1YSDKrCNtotufvrzYUh+BhZY2Fmb
cr9nQv6sHVmg2HkwQ97X+zbUnPd6HxCIQ3OG/KcMTLJBbPC0+hvpysZlr7pTl/CB
mVMaTE1aByHJHEryrbCWDWUiFbvPMiamEMs3R/qiZpiCMfG8zqzchYQNujWz4jPx
k4mmhBQnaIP7bBr2/NB6/GOvoAV5P5h3wLHOCG3RFIJQLT1m50NJeHGheBmop86i
DUYyRhVowfqqZvHv55Py0wsAUPHeQE20xZCWDWkUiAoIF97ZQAxH0T5QEAlkA3Uo
XfFXBk9K9ARG+TodB0616xFxd3jy0YZzpQ7jb9WrKyDeHOIY4vMqm3lxJJAtXlQl
pGSjdbjRiM4g3cLdcABZXvTrU4GgHzD0grgG97MHqv+xmRm8h0PrugAIaqYfQvsP
S+LILqpUPh1Yf2nK2AjSMGnRe7kY7HKK9bZUQNmjlR24ls4AJze6UBkv2dqOk9g+
5UhRid9kHwPklD/N3WX0o5vUPuDuEsjOv3hpwkTFZ5FtikR8QmhRwhsJLAGInFx7
knV6Xxk4vdijj6Yl9Y4dEah7hIVjouUjS2aWgawqW7aqXqOB4yIy14viABiHIZb1
mhvVRMnD0xc1YaE5bs7Dp6hCEAn89B8a4UuMYumTkUS6Tn9/oOdAA1Pn9gftym/7
VLgrq0O5TKnoi5dKpyb08vkquNAdsbTwATA2mwpxDQk/+BMSm23vGCvb6hpOouow
bS0wgaDDX/PKHbuF3wveywa7tQbhNFDHBQAMO9PnV2tHXzvlFKRBMAINvcOzF3HL
Gga8bUm5tE0Obs1CvoQe7gnk9fq4cd458HqlQ/rRo7rHv2BLsGZpheLSjyl0jeZ+
JVnGa8nAiqbgDXGssCq7qNWoJNeGKpx9X9XBNtj3Q+aCKcti2CMAs26kXmODGoD6
qfOLD5M3q4WgD4Ej+ze/KhZJL4sFriQHtqng8oph9L147DAmi1vRKU9iFchpu/5a
CCUof6gwo3WXkBXsFcyK3JtFk1vyEqDB/nx8dhT2Wgb5ukb90DLDXvvtjXp3y7Pj
fP7/D/q2E553sWAlLhQqAWVXQd/yoMHqfIf6yIChHPTxOnGonI/mcyJyMKc4eQMX
vTNE7UtPNY+/LJNtiGyEUn9cQBc2Bw7YSlwCzPbJHyyuL1NK6QMz0uCMHu5wC0A5
e8ZJLw6kyu/FKqGXACuxze3+37HwwkZ3E4uaDxtjDpNnVC7YIJiPmzv39sCSzUpf
zjHb7MIkfE4dYpM2XeN/je4Hgp4kNTeyLqwAlbOYTr3RylF2pX575I3wH/BxOmXK
i56wr/0V4fU+pgxce4M+Z3OhkdFjXlcFDeke8PC4JPDwFaSq2+Lw+rRF1U8qVuJx
mvLRc8Sy+kRRqNE1Hj/1ofHJTkgN6UkT3JBefx84QtggHoD79m5ozUAqY7IqarlU
UckOh5JWs9SM9kwCqk67k/ryDZv/j/+51HzMQePkHC9YC68t7L8xRQq3LOm2og8e
5iGa7Q9SfNHlkvx/dsuL6lADU2slisrCTMcdOgNkrsxyHp4fr7wo8Q+1QcINdzph
3eYzjGWt6jgR2fkVFONV8AuT11NYCucviwMf8uFzToi0vWy/SH5dWLfxn8lqnRso
Q1KAOrsqAbxL6MYauBBVAuqoYumiclZ3+1FD6TdXPWKzyx1DiawlxKWnc56ydRhk
GQvbv3Cor7EkTvBcj+WW4bxtrXR20037c4YoZIZPWMBdbFMLQtn0yn/lBXjW+01m
enwIyJuxWN7kzZcSScC/gnHXCv5SvCjdTaEpMdHQFTW88mNAJ80PAFUkfSqL6AbU
k40niK4TUOAe+PY/eJZXv+kQu+01LphFaYhMBGlXs8Snl8vXDlthqdMnjjw0kdP/
peQKEVpFNBQBdf2TvaB0jaKVeu9eLQ8sY6kINPPoCdOXp7dbW7U4GiB/90sr8DgS
ix7G+VQQkNJ6Ky++o/vENLq9IwUpztwzg5U0KcQSM2eAkXsdvclGxxC5aTQA9v94
XzfqwfmX7Z2le9RJc3rAAUhytGEyD6oEZb822yBeTT+Awp4qW1yc5ZF4dz+/Q8us
YlENJOfWQLzVvdzBnQcwXck0Hbhf65UmzKE2TzDJMqJZzA5YRmT9uW9kxBIIpl0i
DY9HJxHx+ZvVqjLK1IQ1B+4mXcAPSCCInJEoJc+sPOTkSUQKSB3Bsp34AoDRaCjx
7jwo836rN0garl9rzzb2lgN8lqrYeYZzoY0UrqxNshPKTy4Px7GIqA2zKQJazvE3
KzAOFDQ3TpbHgim2mQT86ZFC79dA8eWS8Kns216g85BLBp31NW/HVV1W3BXJfIT4
EPIrb2/93XKX4BukT4hqqHSNyyqDR8hG/UTlVJxAEkylwuTYMJ6xsUPMpFpMLEVx
c+3jd/B7R/188HFrzkEC8HGmJ/+Vn7wHLWIUqbSdp8OPa2ZFkZEjJAjGkiKkI8OB
+HR02jLnvxVbRWM4j0+/z6G0ZqVnZGpmpN5qwYjaXERoho+uFtg7399CISIvYJIX
62VDBlrfFy9IamwKaDKnYhZiIO7Le2mAA6eZxPp5X0hfGx3sK7nszGD9R3YZfNe/
mEp5jmRfcxSVLuGI7f62WZqzcne2Ob2p6rkDtU4fTBflaqpOnrtzFFS+MHU2zg2d
/Ry+3Z/rOD5LOMzMC8F2RQGBVPdKqbGIK8lwoVndT8HrJjXb9hp09Pvk4z1rOHkr
jdMssKKduBRUqZmlqXRPPY/0YccspZBEdg8wZTUYPvccTv0ETdyz0rMacTQC0+A/
p5l1rWZA0MZLmjh2pzDJGncdydJmRdbFGKeLr6UWsfk/RS6K+6QxpkZrC/Nbpih6
9ZvTAZhCxf6zKlWEGqC0IOiUS20KqvaBBJPKODGjVV+OH7LuKmmZf4FxAxIpNN2Y
nEE10/uSzHo2oR1wfeV4KhGQSxfJqMp8p5ICelTQrXrTHhNJh7eiUskYRX2bPWqX
peb6pRoyr3aIB3RYwwoSMru5yF937aAowrGLAPeK4SU80LmuUiefBkexlrCWDf8/
UKVpcPeKGqv0+oukuWlypZQI7W2XT8ornwXncV1Sfdx/zJxAHpjB2CSalGU6cbaQ
CPiC4BEGjcszbprobmB0l+2kxxo35xYxN4Itg9AX2R1S6gFuThRa+WwtN9l89B/7
d0StID87eZDezcxzJrdLX5HTAJ8l3ObhEUNJOWofVqFt40JlkLwpahTgx7kj4h+z
XDIlqxa55rYfgU5u1dne1kZI1EZnxo13Ego8PzjJkwTfTY0gjFNKax9j/NRqnD7K
jwRmnQtbuI9gI2KDVuuGLetirci1DksPmoafuI1RQelyU24xF1oxVCEFL4ncwOIO
cw5JI0CcAk6tvQAKfQa4REJnsl8GKwQekcZE81aJkua3jx/L2n0PaJyE+iN+QlV1
hsaHVXrdudfs6aEIdl5zowR0oKKJJX6BVxZqRpnM7pWOPBF36CUxaE+K/lAqcq1B
prfkb3kQ0y42TMcKPAjiVjwQALbHTTRP7XK+CAwWh/QWEbc8XNyxIMIis+7Uq7gK
fTd8S40BJA97ZHfJAftwtHy/R+FbeUELJUelLpuETcfmcK5CsxoenjrEcrt8WisO
FMivR1ykKDFobX+bRsqSQc0ETpbvs9xiVxBU8PklamxUGxJG28fTNzjOIf5c2Wec
Cn0R8oeoxHRazBafczBFGUlCM2xhNXpV5wFHWOjIT6ldC4rqT8Ackq903sc7+Ntg
M/ZeGzN+twq6VX8LREqYFQh05hnDgzTA8atSvmfst7rn12pOGfOlASCV2uUOAG88
XtbeuLyCGEFSV3wxUUmw9qy5YfUXvSvU3cuSxKfJIDRfjEhbVReOEiv2KU+CydF6
E294pEK9dPC/+sg3vuElnXNg1tp0aDDDXNZG95jnv/2nk1Lv9w5dTdoKLxJOCBi0
E4s8uVgm2HA76J54sTCuyaUCgGhJ30Orvv07fTgMgRT9+wyjeR0YpaoyVi2iS3wg
/q2nNkLYa531T7mAolvME9Xs6Svq7wR9KWygHN8MVGDDTpfc7vru3YAiN1GMYRXD
OnqPk7J9ab7dld9n5RD8i7TOEvSMc1u2jdLDOVg9gnq12rOQbhdR6v8ddTND7B/0
vWBR0B38WhQmYzWXzgA4aF0DmvkAa2GVt4YyjCuIyT+HqovBatRMpHFonRbuTz5w
UBTTbqSqYqz4I0fHA2HgJr9Zbk91MBrQLTodIPS8m8ETULbgZxT3YlUOn1lVjb0q
kqlJUBXsFq3kQoOEIRjli9eAoDVD770BuYxLDtNPUDVX4xo0gjJJpu9iQ398VFK6
dx/uQKaNz4T14u0UtgG3w20aZXDJg1w+CSEUGv8c+oRER7uQYpL3eMCE2hismGmX
nbMN7+vI+ojNPAmp2T9fXQUDyrEVaL8Ro+YFSEhSBM3JAUuNvZ7RVSC4AfKnKjm8
JownthLczbHajyMv4dFoeas44c9sRg+OZnkHndLW/16Y4d56grh6yTKkVoQ+CxDO
+myM4H44HnB3PGn4FQFPM7YNnBut3dL1oP3eYCYT5K0R9nUPSwS0Rnp8Sib48cI+
HLIzAc1T2jj1kyPl6nVu/7HkJlG6LOcuuC5tqq0qPft5voqDC7PP1aAmjgoU6lEk
Zr7Ie0isTsBdXZKuLsIc+AQ/T2/S+tIZHEy5RWNofM3vMlc1ycb34zS9N0UrYhcH
tdUCXTsiItOlRCSIGuWnIs45epCJ9X45idSATPQDuddIvHBBHDSevcHI2m/59kHV
x9DEFhe+Z+6f8yMdUXpJ66WjEXJMW/eFs1YqZZ4jvUZX4+Yg8dVjC8IPv7AfMgrq
cXPvEfP2B6+deBSp2XdmOnkbpJ1MEA/r/qs2Xkp5lE2iI/vVi+vNF5tSukfk/Wej
cu6dlfrxTh8MzObDrM53x4M+SFh+1arEIQFe+06/YH99ueToASeXiSY5jTCYYMec
0k0AxrsXx2IFjfMvWY/4lhIFl+23Wt58CHch9BrCjfbub6wj3qy5XSuhCACrcFvz
sRTFsITznEcf2VfJq74ncQIaTv/P1aLSV6loK2Mn2O7wHWPgDgndd48t5sPLncom
v4LcLeJGMHfdc9470gdGsFjAK95vSwH1RsqdBRhoKvOa6RPds78rN5laY3VdVJwx
pcfRnUSVT8vq5gqfwrRLSqUoUvC/mDugz6wkpVzLLubIqcTb8FA5v7fnKp/CPm5d
g3aQXRxBN6JpbmdszYEmMFU7vnBaE8cFJ1xqXuoYh6SYLZpdMR8AHi+UJDKNF8zy
nd5qrM+WzI2e0Gdbgz4Vb/99myUYvrGsbRxLv9DvFjj/8C9ylLqmuV4ws2RI0VsL
MraeewDWaQKySSjEz/b82Mv+NUPyW2KmHFuO1ACWaB8Ymic7wgCU8rSXYG1cEScB
aGmalxGIyBq1AwyW3Kuqz3acMPwF1yMbrjODOUMAT5OLpIJjZcPSKrX5HKUxE1vx
9uZocONmI5XQ1D4vualcmzQLD0VtPauSKtTXwuzSxT7Kc4gduP3Cenw4awewO7uY
Y14xK297JMWzzGwcyhR4vR3/rkHcfu11MiEL/Up8AHeGGTpmTUR2LC/F99rP0KmT
Lm72WKBpKVzle9asQABO4qC5mkv1yatamGUolBkKGOVVccAdLBmeScjDquzeqAW9
sj9TThlyHrx1sV4xxug29IfO1Foibw2v48fznlrqHbPNHppG1MKFwCuPdnGNVQNh
sRDuFUSqXIlliGDP4H+C77CT+WfdVCpajZPGnW2SxAn0JDVCq32Vwqmr156K8wX1
WAUs84euevI36kNFpTXLFgiueLFnuIRgyVaYdhAVL+rL/UnXn4+yvBnF00jYYrJy
t4wPLlwvqNawZDrS7+Hd0iufXMeoZ3372IDUHavloTs69lNTMRtwV2hjwcn8e6Jc
YN4K+Wp9luzpngXrL75M4zZu9uvu5gyJYCdTlUp9mttlV16jICtPHpY7k/Kg+SVk
A1ODu4j0crMgSVYgIOo4f+S3MLGrFjeDTr6eaMgkO1MvOMS8QYVGsFJQ4mHBsdHh
sSjm/PNMlY7RQ0DssSFpYWagAiTfgE0nGlHMWShu2ILrE13/YARl/qfaOku4wp8M
pipT7eB3tM8joDnIgIXR69rZ90uwX5nrffkz1sN2wr/0pz0JgkKQutIkgUZ+96C5
iZ8wN0pRczauYnC3XwrP3ij2lMyD5miuHa2pfI4zmSDCH0x2BrclAFZFQ4p/zhC/
FskbDfTyJIOrSoezVqWti3iX4A/lTAnBJQQp/71QkpWHydXA83rZWjIM/yUvtLF1
nAZTGJt0M+yh9OiJnuwguTMGvjX3KFQK6wiWmOvXKo2iRChFpsTUHoF/WknxbdKR
qJj83GhVrdkVGesEbu5DlJ/BevKA7adECIWZ03tv/yXHa0iWhqSJdG6qrBXZEsVO
EmRquLA9h5IobrD5XVPQz6rigA3tEJeWwCJFFwnM4ZuQr6tB4nJxtKc4N+kZzg92
G1BbaKCwREI0/5/Ly44arojBG7Iz46KPr1m8z6yuprfKEwT5AE1bcEvXWz51Sbiz
NOjvICbNDab5gzess6hlf7wxr8rFdoy1/+RENi3W8xBgu0aY/e9CgM7jVbbrOfl2
urf1qMm5T1oATVMlfwh3YEobzmeRQtUlfcW2zz76/x96tl0gznMFc21B90pe4zGY
aipb9pWJTi5PhRbUJ4+XbVJ6ef7FROIMcEhYG6LNlSwCEWTImwWdGPBVXTW6MXd9
i/qVC4ea/XxcAiqD+W47EU4dyrWd73dssq02cPYw41h7ZXlJcHccOcJQawQ5nNOd
/vdKgT7juBBh+GeStyJ02n9luf1Gc8ZMXTNxZOG4e7HpoK+jr7J7iTaLE1dcszyg
2COGFcaydtBINmczcWd2JEgb9C1urlkp4k3jO5bpNp4d9YhyglRNNbaFkMdsDIJg
lsFuaVdkWLiN+tIMXKgq86Oyyhs86eJjZBAbzjpUfu1DB+D12CsmSPYUUvvy0CSM
cPLdDKORP/o5lj6FOCB4H2VnQiGSz+FnzULknVTmiuxFWBOWHlVd1maBecOWWH+O
Yt2KOrW1UDcmEn58OZNaazyCRD4vXOnIscmNbuaaodIwLUc2PD0vOG4U7YDLOpdy
ChySCGE9t2PTbIyVgLGT3D0UF1z0ANcshE2Ndw6MJHB28tBOAbkaKrNMOWeYZdhC
++xBW+ti6gtRVXyYFQxBJ+eUYsbw3QK84M9sbYioxjvBnJ7vDYh+HFEFm/fMfx4H
wnaWiSAkyTerjlHBLvJG3+SBCSBuBjq8YcUQ4UbrYXR9XG4QyASCgm4qCbay4fEd
eYtOoulZK16I5LzJKhZzMYrAkvCKSHHeRDzy6jPo91s4zyxrG8yts5uR+XY+c/do
83gqTWD0DeAII4zXCPui9msMqZkP4lmXJLs1tiDB9iiK/jiLHTJGttAxaMxL6T1s
qzY65OEg0chH117d4a6hFrtnVMeSRhLh4tHam0q0WR84zeqg52lQ5fxuLS0DW+ib
02tKKLLLr/8fz2TPmBEsMMpNZgQq7rHY3SZq7ULS57zJYm6xDYdXaJp2cGgizGbm
/FxHXlUApSZrjoMozlR/Tq5bQ6bOhfvNlPrI8LmY8v8v24H6fMX/fyfRs71j4sPA
ru22sduLzkOCptEBxBnZssLklEeLPRmF4qcklgENk13d8/ZO7Z2plwN69fZg3mdD
Xt+u3G5fGNG1K5NZhpi1cRzN2i4hGLWEYKjdDrwhBGUJawSX1Gyz3Be7XJjGXJKY
SD7Yy6j+H02t7cJJHY4DtsrIQAFD21YXbusGBxJC271Lmeat09Y8n99b+5Nt7C66
YjswbEYKMfGO+Lc87nQgMrMfZfaQZBjbTFr9IcBtb/GTfl2yiLMTTpD7DC4NYrCP
tCYdX6mPUqmqhNhknwdiyaYK156dWz562LQX7bIK3f7nkWXL8PrXL1TyP7O7qmqm
wVEBOhAROHsP0s1FRYc49clhPB8xTkBZJH7JqNgBV/YwvSChiNIh0O8wWK9/GlXk
vP4gtrNEx+5S6Ezwek4mHD0RovrCbAWLfLf6wiGDTttIsD1ZdQ03bBx4XstX5uQL
9azw+EjD+g3ls/ZdrGF/L69HWpcjVUgZigMKM9jtHhvyaAgLNTvOHocwqmSOBoE/
K1+tL/pmG5DJGfU9ZA3x7W75z8qhwLjHubKFVmcPDZMoFdzFXv4+9a8NXwj4AiFP
a7aMB1NhRPQBWMqiiLvbkg+Q+HisJ4ab+xNQEgnVx7oQ6L6PI/HkG7qJjAaePhC6
asdlfbJUeLP/igVCqCA6BP6ez0rCkNyJ4ujD4rJxSNLKz70Phi+N880zNdDGBKEx
JrSEy9uGqO8/Z5tne9p3reRtK74qbNgQUnTzDfP7hM19X6yMVDue6bS8gXWT5y8P
FkXNrjsnaSQtErmoXGDAj7wNG5j5pZITh3Y0KOCD1G3RVIHIYcldSXjmYuCLFXKB
vf3yD+guT5w83V4WPsztt0TW4cwEGB5KjpqTu/nx46fskxmMbYVUh7wcwXbCML+T
Mo3eNsv/SfoikJ39gs0x+HHJTD18rIqPG3i1l4FoRV9MoiOiUABz0u0bbaCt8sMX
GiSqHZl3yIMFO3qCvVr0LoxZAeaoyJmjifsCyDSyBUI95CP4mK8sMWoPDwpGXnpA
kO6SDueq4TpiUW5r3UYWiyjtqYbnfFJoV33erkS4xjYq5B8yo8sa03T14Rwjm9YT
A7xwgotijp71d2FSXn3Y8GdgKuOyXuEU4ANRzhwo2kGZsgy7j2AKQ9VVqdPq8rqJ
fXfnfNpVluI3feN4FPd6ZErVXOVthGvfmvj0dOJiDdBqBp+ewdvHDhaSJFxnbznp
tq8YumXc08cGNaAbHNsoaNcg1GJ/dXOzXbaqm4UresPDUzuKdpGb9LaKMC5qaQae
8H4+zo+aYRT17np3jNaHJ9HF1kf8uNGY5kddCoHYKLGp6gvHuA36j+XdBJDACU+r
f/CXtkDxC/FwvgfgfLU5dvT/UU2M4OcxrwV1NDGZJP/gwO2iB2830hI0tCGulTHX
t4WaORnCQwz98C6g/8CtG+QerFTHAVZV+wit845qlmzZx+QkNmqU0RKwGTH9DBj1
fTZbmgrDGOY8PPUwoFyrXJ2mLzxip9hBC4SQGgDPJMHkVnOrEWKsfjGTkSlVVhIJ
69X7ne42L1Nj2S2YN6BjBqNlcM2efE6gH5x7/6Wiu71II7n8XQNJgbKJTFSJwltY
3ruarlK5pM2sZ1ZQ+tysbwOPABZ2XZSKv9ObrscjkPVqR0AGUlS5wx3Oeu/ufDD3
+S6UYw0LmYuxapiXzzRJg5hng1qo15phcCCMNzBVvHExnzHNrpk6Ctxe7m1RXgFI
J0rlj5wTexNdWIS97m4cSEnz7U5v01YlE1hf5/1A9jL0/UiyjW3lLiy/VdmuSY4E
GeToQsB8oeQU/OVrJ1FGRWJFzW4dU77szA3EcZgcDsLZgK1J+3ZxGdPB9P9Za1Ds
QgGN4KRA2U//YtGZgZeAcLe0dXzwqAp4tUhgvj97cVFBifLCNkbmB0tJYtTWnZNx
BdJl7GycMKW8EvUZxbmM/h+RWukimJasuSPrZEVEWPAkCoEZMvABV0XwbJbpnUe4
eL71axYTXs4DOUVclbziJY6c2P9sD+EKaDobm1Q4zUqDaNSa9KUAMRkecKfPQcfW
gY1Idw/ymWMl3zgZlSUXqbPyCQD13/EAnxffE9VXPmq6VCEfJFPOF1aKJ3Jsz11a
Z9DI3ouor4R7GiBeVR6jHleRgl7FdM5wGh6FROvKeIAKPtyKb0GweZZ7mTzbxx8W
EXJ9aYlJyKWSVUK5uLqty2cd8yFGO2nfP1tvd0Y9pF7MeTTk7gjxLG22i0oC4onQ
SJlaf3TZ2zi7fq9b8u48IKvlEHuurgMm/35umuHdcCV+3OShfLYUi/s+dGZ5Z9AO
lhLxWZV7hvjE1J0r6cimD1SQ8qr1mqhowVGlE0QYFD5DM9rYsRyei/FR5w/bYb1V
Fpc/L1CRysekwmisVlT7Jzk8TOv4zWFS7FOUgP5dAyh43XsWV9scn0TsB6lo/NCo
JSuHK8/gOcpYSJyMbRa/WoZVZ7KEW8nWYQaaxkJDbzWOdax0v1xjSLHiMScH4dbJ
Clur1yYB3J7jlrkES0CEw5HGWutfdVwkDvkM2PHnhnDX0KIn4PVVAhBB5J5w7u25
TvBWcU6AjnvxW6QmkvG8a2acQi2R7C8Xz5yTyqFCvtlkipILRBykg3JJogmKGNls
0eS9lZzDYV1zmDW5/AJbZ4NXMKPTUEhdwxZsSJGoMXMgZWX7TltEszXFTSpEXgzc
Mn+CiTKZeDVMKIW5p4VHoq+uWpqth1I2OK8wwoXAC4qpH0nNf8qdwkb2cqN5MeAq
SG76mUPgg+BVpoylvbnONQXeQipi5Tgu2e7jZwkHXnzFiN7tqhU5aSNkVeFKJrtR
XW6akWTABsk0EY3//vo8CeFhk/ioOz9Mj/R2XIhJQ7jyyr/LYosQz5MaX9HtWyr1
3ULjgikMdWtiQjk/M5yg8AETbvbTtRxF58WES5e+nlngNPvlMNkscS/xCCfQXwfA
ARYm4U+V9eufSFnchppCqchfjJ/G+fXsvS4XzIMVC9bY8BB4xN+GDEzuqHFozt2t
blEHg+J+V2Tx7QEPVPaKnzG4+ANmjCIskIm/S5aOnYnm88r/cDL/9+pwqV6RB6mx
jLG4GxrIYuNV6sda00CgTGoP15ay8747yRGGxK4VmWTTRtEzgPsimHi+edv7CvSE
/a5z/tDVo1Dxf+EWhF2Y+mRDdhIKWg5hkYqry94Qoca2nK2fCX0D3lwwAG7ufBq4
ZO5uGCOwonuL3mTZl3J2Qx07ZdRC9R6W83uiI17fwQ/zEO9Vwv3Fp/tGD8oD0buJ
oJtGfNP20+/LoE5HVGGvDK66I6zRiCbo5vBaSbzLuVfq30LLt9YVeDSmwMaSWdmU
Sjb+QHS6d9EoRauoZDx0+7nvF1np8S4y/jQw96NzLC9o/B2QxwIWA65fGyFMBQqN
D9/xd6wg6m91OOta9Fe9Gtfuz/i4M023aWsQ7XuvCaRNLCQuYHPQ0jdODe6CEVa/
nUTfSXQLU9H9kwBmSTJcIvSnoEhWEe1W07973HMThD4BwxZV5hsHusLbABCbIjjl
3ZiJFwG4mc3CJ+jlib1IBGaRynZI+hqkDECzmBo3hC4T718XMy1py+hfR6i074If
yYkVTmHxRuxKrgPPhpf6TDIoOUwX+tVm8UViqdlitnngmVCSFHe7s2BeaRv6J2oU
pDEqkIQM/RN9oWyFcRWTe4qlIkjgrPeGdm20WzbRlj1gQitK7nTK1unNwglT7irx
QA1Qs1uOYAKZe4U1wbiruNtSim7Wf6+IbijIOg+qKemVugKeMEyjQrz5JwpMXvPg
xhOj4YYkStY6mwMxJSqrTtxHpJK3LuWdZucpkv8PFtP0ankFBIzqBXD6ejpdgmiN
mrMO8qUdpon0eeJkxlinHD9gFCVtncDW1E3+I9WjaGAUqfV5YRcZa8an+86Qqpge
2s1kuJ4plM70xb6tkCeDtWZb8LuXC/pnRPRxLF1Yjm5G6tTa2Xyjc5+JyUkEXK/p
DmPHNLDrsXATdXckdrZp3BtAT/0UoMD00hq0f0OqBctNYlnqI00guKm0YqtTnvyU
5cseNwNwtvibDSGdQ4FIqOh2CD2P9yS3OQ6N0+0gGMYooczjgXRmdkMFvHPtqdq1
oX7koPl0C4cGWOa/Qn+nu7UNYRnfQzDNInDzwgVe4DtFY49aKLaNfsqYvb1qay+z
elTsKxzZhLzU2uq082/O3AirymEMk8b+yGyG2GznRUgQfB+47w4dNRJW8C/miOHf
jnNXIJM6umgRHZBlhCvk8sXEZwObblKa/LNbtga5aUU8zUvS8JJ2eseOazzudDff
0W9gF0HfdGzbYPQosJIQ1OMxsVA8z2pxw6EuEomIpPzX2Hj7iJh31mC46lNy00zS
Ur/UIfPuE/FIViJeH0Hseoz/InL+5jWLpoqAvm3Sj2EADBWrJYWpCvSem5dDk2ik
T1gJXPK8WRZ5LlPwnQwB5+4Z5KfUX2m/Tl+0e4Jk0dQ1cA5cYZfK+f4uYGmJHnMI
W/E9ZZLANFjRlOGNuCvc3e3mUGFIPdp0QS7jc7v19Zqnc7KKi8Y94l3bQBcCW0XO
fYcrmv58P1k2R1aSA288onBHYZ29TKT8VZgIIHgzQfRkmV1/04lHLb1k1LMlJKtu
MrrKErNHA77x5TDfc9TPQ9l3lnQPxMppSfXJHH7U+yS6Ex3a+GAkx5PQNQfezZsD
2U+75mqO0jgY6csKlKq4JScOEDJ/fYcdVD/lfak0mkKogF6GkZAzXpv1UzbyokOU
RdAUkd9+s7py6AIV48m9PfEqaM3AHH+SfRzjKgpx5yuYW71Z/0fZgO2IQC2YxLUW
cDacLigBJNGd8IRm/KQNsyN3QFQI/rFl4pYZjndCiwg+w+5z8AjOqvQQjkVDUif1
EF4vSU00XysaRUCrdoXQc0i37MSl3ZSpZavM9hRfRUJuheJYlWTZ3ZEJ6OawpHv9
zW5hhA/zspN+jti2OmWrnmrcs/kDAnXt9WsuKxiiRiqK0mXK2t+SkaV+va8RVHKu
bqTAKm/GnKeOj7cRR6UQhjXgaBB+xr2SV2f5MuTkVf7uvDI1W7ciOM+wasPHH1Ck
LXc374QjjWHzKBxwVRsoaWgWmAqgZFmKboLvi705iDwHeYGZBV7dxJ7dU37DHn4j
JmdxsGcBWRQgKGH5jSaBIZqoN9cZw1O6RDbp1UK7XlixGtq25xkzhrEwsgQcGzFe
LX6PJsa06wAdk8HggVXh2cXGY40B7z7Jj9dtXlQV92/0icTrEBBxWdmGHviJMRAu
XkHsCEmkap237GpECJM5IxhuTAjNbggw5RzqjrjuhkSnYWBH3tWgUhT/+SrN6bZ0
XFtz8pUzVmEdTtFRZmvGEBIkFo1y3nRs5On5k155KIzOai0kvye4XGHLzxN4z1tZ
+7rsBmVCVBZRLGNtSColOJfXxpwCX74seUoUq+5ETjQY5PKRwJkHX91GFhAD/QaV
R+vyfkHciehbMoCv6EKCreMGvQh9v1sHI4amoSa/WylCKAi2AQqT9mYh6l4dTIis
9bqHKVRPurFNtIt3HcMJnmxbUvwasSQv9uWL1EeHt9eNPmoNYgZcNYSdE4GdgEqR
7txdn0bfOVlM8TWDp+VPcr59T3nbVI2ylsJwkq1P6RJGKgFm5NFhXLgoWOkKt+Nl
1PaYU0Pi6OxbngP4orJPiCe1P+GPJKncRgWCsj3l7zE5Xdof7UmOFRHEKqE4ldqa
eBY1mbQNqxLWb/CvoL3r4589lB+wzP+CzmupSDRsS+Ixi7OhYUgMbkW2PIF2pcSY
1RIZiAuEEvKBGu7ykXk39fzrguqY0PYSoqUebyFEkhDWt/k6HZhL1PjdPgYdjI3w
7CaUEbQ884OLegm9cBZWitzqHsRmznSEiLtf2Z4cXosH/5gGxZBvhYX8eAtwLa6P
YhxT2QRwKJQN4qoIRLOMbrN+epzwzh4lx3c3IUUCZNgQ1QBfEN1owaXVrOU5yk2/
k3mkC/+PXh2jCpV0P3bO0N1dCJJYZQhfTUZiUDZMMwfk3oIjYknEkhefryoIvZQm
dR4MekIDJKLe+aRy2q2pLb/yu8dXKSrvFuE7AeSce5uGcWbzXUdwMTYBxo++u0y5
A1YrraRtSK8T7EhkQ7kSaY3WQDykpSmx/5aoz2rqVv8OA0HwzWPsYnG6uQujuWW1
HsANa0vIfxWmnn03LzA77wkBx5gbRhUsXz+yNqumoQabjmRgpDuIJkL0/zP6XY9O
AWHGyAhnApZ2ylh7E7Ev+fKK4Bu/MNjcMmbKfHAMLBYsrE+Lc5TVG2vxbaPj07o8
Rdr91mIVmNjqQbgGzKwTSmX5O2RlmYHDG7PbyE0Q8b7UgnjhxAvgtrceNEEd8/BL
abWEgau44qt1KLl9TrFeLP5pS67fkq0W4VhzxAE6KjPzbXPUIlj6ixiCW8Y2y1yQ
I0RPtJMsPoZ88JvKvCGpB8tkZGcHXiYURJMKkRpGOIdF0eVh70CELFli36swUkut
LCanYBvA/jYeJzVRkEbJJ5X4agX4xun7a/Vwu2TB9KLZo1vQEgC712j+O1zzRS7m
O3yL44ZfAOtJogIFAc5hC2/Y75QBPjcw87HPw1/Fk+dxf3UzEgjqWHpFhVhbzfZC
o3kP6ov8bZKBFzaUQezSr+1BjfHwh+dmiq2B4JbB7iofqvpnPKI4WmJsZh39K9+W
F/kJ6E3gqTDMcTs3w9zH1aFbCb950FM86Xtdq1fHfOexQrDrizjcQkVXJq47b0wF
ugITfjqNSU2KivlqlEYdMOhs3HnQn0yxicWzaYEi70/RO3MLKVy4u7uDJ2itc/8A
Q77mb3esLw/A0RxVEfMbp/NKbdq3FF24ylFCELfM3RBamlB0ITwTEmrQo6tkvdgC
WIUzXQnafBtdKLUi7mtDVSByH4XNsiBiE9OKFcHMNnRb9e4PtPwQKX7aslhxHmAT
vkgWCV2ljgJlzIxT6fcJDrtuz0ylEb37KdF5EVgfcapZqxsFUyKG0zVd4u2+v1IG
cqJxj4Zf42l7WuywOWsUNct+4BSVrm6x5JkE31HcRbVbnXdVI+UqZhV0RzJA+iBf
PAoAbTw8E4fjMqF8j/KDCJARnB5l4vBKdQoW4vYCafMSF7k0iCpRgrYRUvaGURfO
TZWHTX8Dj5zWrsbbmit0/Hwy29V7rRMLaUcjPaBfGlYKgq6tXkxdGdn0KJ/Ve/hf
sxGRx2t3j8MHPkwH0wQrhOcaqe2F1N1kdKyjm2zDVbFcfO+OcMkYkMS5OwHetU7E
9JFVjFKOurPBwvzu9P7pN5pBcQZ3LkF73TcAltQ8i4nJAby47La173HPSXItXDtu
2DVDNgjaM1MWurR/6D99OVZ4KNXLFiV4+qR3H5bH8yP/+rSF/79io+JqVL4lAUgA
HeL/Vpp0OXR2Ve+6QyJayFRZsC1TkcqmERlNATbg9Z4pTppu+rPqFpkApfOXlfJi
E5FxPeFkKQil+lltj9XKsQO551b/UdmLtSZxxrG3wWFqMf6UbZqjovjjVINn6iPS
zxumpZfdqr28ja8gMQfoSxWfW/EJAorUD15o60XFG3ApfafWsUnEFoUEVwV1U2ho
zB7UmlIw7AOhCxl7uH1ORg3bOfNl2L0KNjEKQRxt2UUphSxNCg/Vk3hxbSzCwZJ3
VaNDyQuvN9ntD0Bxv0XHGSez2xLaM176B7RajZ6OPDRb3vGCNMSQAx9ZETYrVw2u
ogoYSHoP+rzkQNBV5GcaCXgSbooJAvjRtNTEfN+LUt+Rbk2hM85uPrss1Y9eKcbV
vm6oDPc98HtFKqqH+3iBodje0RM8Ow+bi7qdU3H56rkXX6Ok/EX/zK9MiaXiAUvK
oEJVArjsqYx3IjpzwVYoic1ddRMp8VCRwzunidEhKD9SKsOosSjQY9RWQyxce4Ui
Ds4hI3Ayat4E7Gv9wP1wX25TLG8T51UAHd8jvzHhRkyTwQXZCSDkcvgD+LeBt7D0
XhhIKFn+URNAy1X8nj1RRaFMzjIDmbZdRcsKFzKSeouSr2oxZ4t2yaPqshYzmPze
WWhue/mZfn0e8eJ31rmBCf55+pWghmIj126RQUfCqIowkdCeUIh2jZF8EwnavfRF
+sjesJPD5WJe2hnb+PapUwP7EVjUbBsOUbP8YzOXpoTEZMrSi0Zr1hr5MWCDqFP0
45VkJW6TefcxNHuw+2rKEG5rbtislLdp3Q7KYDn7TNGaHs0VCXflABMk6ojrw7Zi
zUiULtSiejfT1iPRfbzL6WhbD6irzMN6k0xm2uHC7JtBZ5IWIcGUIPE+Iw9FKNWa
feq5L8s+vaIVHZ5KC2a0FpXl3UYsLjXy8xtJp4LpX3/vU2+03/GSFeCJIFmCjesD
2XLfw58HirohCJNhMns5MgSMSx8hn4ntHh+/kSazQvqHJ8JStChBl++jaVsO3JDi
s9YYnvtlutBfEikcZfZZghR/b+jIOgnNjPenEHdd9VkaYMbwV1iwgGUbDGaQTX0z
XN85rApbI6XUwkJZTGlhgHlAGu492qYUfNDsW7fTFP4ORmNdt+T7gVA4DlTKNxJc
pGF7a1XP3BN0yZMbgwK1mcKDWM6ZJ1bIocK4HYQO0EnCJztPT1rewYgFdvUBNWdh
9YMQWaV9a2BiT9y4hOKZehIFmG6J/++kjeWaaK23uHKcJZdJj7Qz/9JCz49nxTcu
M5bn8+w67pcE4kO72J7TOTOQuAsucMICXBUKJteDWDZgyMFl06r5vwI4tRR8OCe+
Whm2KPcfkyYG/JFPfujQXdXAx5OMjjjlLxK/KK9ZScMjMhobYxCPllEt4lM8Xq5s
Pw9eoaSpCU7ch6AaMDpLZt/ZlcdDWcM/nVCtBY6gMKG+LrsfD3sqV1w5Cem8DVPk
f2MloaeJF6muepA0W/ybrBhvbBrCD3StG9UHo6wHMImgxVA6nyas9lwziD1E/J8M
8uDM+Rm36cRJj97c+tWkIFV3XkYaYJUYAHFQGwneDGSL0x80a5kYx/u0+4f9AVxJ
3y3cB/zOch19pkB8wzQ43vRdnXXL8ZsNrox8Y1cJGGwwlhnvWKEgvEyg1LpTpIWG
/A5yeI3ruP2Ok6nhE823GVFGQY5h+RsafdkzMMh43fpo6H/GACFDJ4AZQpoOzMfS
8y8duoV/BH7ZUovo6J3q/pgdHFNnod5f+QGDdzUbI6VKh//gLK4pz8fdJepsJb2d
/Aku1siKGuZc1DnfoK2Es/1WVS8f5UpQaRudhnlYOvIuaiVNHVOm/AEbWtYRC4iU
YWUnK1FrWhUpmfqYra+P+K+YXlUq0VyB4cb58+A0x9nleklvN2/iiza9M8HlOVn9
tW0QJr5wYxgNxxE3q6rtoEl2NeGRgZGjV4peqTirTrtoU0Rq/ZDwshu85MnoSx4b
reWvaNkY1XiedpQzoZft146V2VSzJ0ED31GpWQLpp3QrpGrxAfmWDOJ+03USf17U
o/+CXQVXqMmi8OIXmeLgTbtLAmC7LYfpAqremF8I4dWPz2cuEhxKc1W0UUM7eAqn
+aMnBcIjvfsd9XA0fGymLS6IB5U6RE2BzlSA5vH1Xc4f3S33RgxTtyi2UcmOB2Wi
d2FrdTm6jPf6MRWFTdl5JN8zqba3dmktuYIJ7SAkjRkHU1o85W5HAE37ncXZSC0w
bCxy+6OHbwMuGW+RyG72DsH4rqkr57UfHukwzSy0Wwnl+CssI3oZCsinLCB+cpRB
7kBDg5Xqe5Nu9rO/BCtAipKFCwWgqIfybZWsqu9P34TZ+6StB3gK4hdo/7ZKRdbz
k3BycSPOqjshtkwGueSK1+w6rRCSbg6BEA4tZv2L3kn9j/TbdOUTwOWoRugCKI0P
66tDyF5iJoKA1JsOEjYTrm35FM1iDEAQ0dwy3AWYIY03nTRYylA1RU2GV8hP4FL1
M+8sBP8s+DhhynTFU6l4yn6Acq4z2qs73lV9RGpX6dtGfiDn1Rd43lGMRd78hpom
vfM135DYGzWlxhCyGIQEq+jkd76l7MYuBf5JskRm4FZtgMkwMfkRN/KQe8jcwxY3
qaPpSKZcl0SaSt7u1fzCWztwMQ8SsArk/iet7rJ/Y46U2azyUOCK1etCsAzfZuRV
A0DhuJjQ6plqf/tT27jfB3sJXoQUF0u7mpbBGjXs1VBou3ktc0DSso/BTF7ap9kf
oP7tfisrIdlavf5f0vwluS0emP9AjqCfBtjA/HenaH/Au/IBplSmoNUqQZosDRef
j1BOK9DbMWFqeue8dA+83caORxqKYnCkCmQBJYBPEPTP8NdXXnIMmgCqulThj8kM
P51AImqDN8aZUtfwkLT79pEqWEh2ye9+EPVXelNROMs97r26ac8PKL+3BDVQ3AOX
JlTtL821kYD+X3mlrOBVK2C9Gux+ainVfWnppCODj6uQYhielNmpEfMgl+hkTaf2
vRIkXNHvR8DrFglovftP7KNylsxldBSibX/lmxT74th955O/W8s6IaXHUMx57p1a
aCwFHnaKyIUoyuivXQWYtqT63xxJWhyicIBXZNIZUZep+oPB78Mjhy6YTwbGeDC4
dgIJHzaVxuNoL7F0n4DV1Z/dNPySO1D0v55EsTY8Yxt1NyHV8MJ7hJ76mJpLfZD+
UlwvF6fo/R3ba4zPOnaP7jANM3R7xzTXCuffINCWqUw7FW8bthhAffr1TLaylAil
k4nyKyHLddRE0UFZ0RNayfMJIPBrax1W2wMqdo1eFX1n2wQX2sVFQcKpI7y2d+1u
u4DOCQG8XLFos+HgpEQ+2FITfNfM5nzlWG2E5wQslMTBKJLHVRd/SBxdKasapcbg
mkQlYRZ9Hn+4njQRECRZBdx2E2qa/DBiCJBjmEPVLD7WMTOkCKYTlja9VIFbZRt4
vwysGxcbRyuUikTvFAwfuImfLQJgYdTwzfQwRO0wRLu9VDBN8sz68TrVlq6JNQDy
nte0PLxiJoccE9pb6rSNtag6le8bMwxyQXnjNhjg+Cj0+2oMwD7pE7cw64YOGR4L
v+5daO/zSR2EhDu8+uM5cp890AgVl/KndS689T1F2NECVD0J0gtTduDSOUdI5tqs
BS10a3bMd93FhZzY31IBRrtYvR17O/CZvAlSnM7FUubUa7kVtGUbQhLxkHQrexrs
uz+JGnYSZNSIiva1ptisd42CVPGD9P88F5yrY3YXWt+BKX/cJIibvZpI0pHp9oqC
+eT49+c8RmGk+Zj7qy7aEHIVNJKmFwJTDqKToaLV8kQkuMn8AA34IWVY1EmUkaxN
CRsHvqLa9h+wRIwwKkXOxUfE/0alh6cQQdQ3YRbsrqFmlvBpixOz821rjICTY1o3
RHdOglmLguM17zWTiN4pNNkaDaWd9lES/mqbWJ1YcTyO27gSNRNTya9EWAp3c036
wwqG3RaPahV0BwSi2Rgen8nRljSh8DrHMgGLnX+7armeWKu9SbIDNUxCNmG8Q+Sz
kTDGVrDwERLASbCSz7OycRxHZXQgDKGks5/vEmJGEzwrNvPUpAufcRFMmjLvgb73
gdj+AviCQmJwT1xkM2MCqbOtbou8cWqaNUBD02/Fdr0SL0AJyd9bizhmsQwplfmL
gsfmy6gqvHgkYEyWVbwrtckoR7BNjQammbw+B17ZBCbiNBill95Fg1VtuA2L5bWO
wPYMCuQ2DYAxhCSIXAb4JCV87X28G39TBSXHmalD+s04BNA78qkfyA2wbeY0h94Z
oWUbf7eZ/XnWJp+/SnLzeYQZjPKHdegL07c8rOWzg3PzvSfcJHPJZ6XRwvkvLs0b
IQ9VaXVPzQeG1R+eKvnBLMQhZ4PCssldH8SAlp7cYQK2JhmdvXISozZty+7b0wk2
eVPlWaVzqIPbdN1R1VcBABqEvHVV2nIzEqVbADktffdnImdDiPbiMXD41eB3SO3t
rJQxqADtzfC/Ned6EQmTHM8GQJVwqmx7hgwI8eCtDaN04MMOqXJ0EKuaHDVLzIfU
hjHJqzCZDBytwOWCg/N34RoQN3uBuKbjiQbMm1XekvsalkBL/aEHBXsVoxGPgtG2
4g5TbJSY57T8UVJ3oDpdAAV0dAmuEfdEszeHSZ3OwPo3J2UgtykN33FSrpUlLXno
YzG7Jowp1MvwBLKNgsC/6biIIoFTsmcl7UdkEJ/kSzP5kK1E6CLbm2ES6heUsXXb
+V9nPV2qJiBtCIDFX0uYSL3KbxUegtHjkGtDX5niQ48U8KIDZE98u1Oe1v7jCB96
dQpR8MSaZYUeEoFPriUrNspJuX2HuRg5NA+N7unw4J3wbuuYR3W8wGlzyPfEwbwp
gndQ4rMedXnUil7Tj3F1gwJKx6US4X0Kj0WnoxfxCACvlhzwHbgiIv4QHmXAdae2
FjJozVOmYZXqdbyRVJi3P/S+CrMLY+fyXX3LJCeXO5QOCSUDZX+d+95L6S6AU6Jx
l+nQC9PG9yTOhAxiIKHHySEsB4l/+4pqcp8/81g3M9t79iA0ax14+c/Jog0YydfD
QnPQJKSfbY8lqBfBNCSOOSVKFKG3BnN3CWV4PzLamr6RPCzNb6CX2zwtiI5lCaI1
NXUKWEx4xPmKuv70fuTzTPv8drsXq3DdOsDIYzzUBQIbEzv8wHJHTmigdMmlm9uH
l3Wg7hzjD0dNwj26XKu7L2aHbNujTUPnmG6gLLZgAlP/nCaNsrvkcipTnWz6WaD7
g/FVkf79UC6h5fzDr6VsfDrglaYabcG47gZpLUFVuFV7fgkKqk5Z/E3XKdOMqh+d
ct4MjPGuI5+uy8JNWfiR0GKy0NeLHtjpIZzdC6I0YnAW14zJnNwKfVQhi8XYw393
LF8TprXmv44XxfpqXQO6hEBJRffQT2cIQUEHMD4Hr1QExYtDH9nC0NaGWs5nAI+r
O0jhIzTiOv0SxihJtOl7PY7o0SiMBiXPHmCfkp5nJXrR8eljhOqc1QgwzXHW/Ypu
WPiozgrSw/1JiAaYGk8YcThFF+q+aegM03ZC9Ijr8lScfzsaPGQyrnDK3U5Rb9mG
JC7pYk3poG0K1zQVS84GguiNiBXEyx3o0qaK+lKQ9yckupuxO8cOx1Ql3bJJA3Bl
GUQGufm/QqEZ6v3g4n9MEGWJsbyekPaDSSSYKxu1DE9bSE9I+u7gjyrh+HWSGTnl
ozc5lGyO2csOkuWkaasMNlkDhHgO8TGzyYtEJ/x801kh1sSAJOuReGKqwnj6sjcn
SwAgrGnZwzpOrvoC1ASR6L0H5MM6ZOV5vFdtKvll9DOaj7LqiHczvMy9bvtojgtJ
Fmo5hvPRUTlSxmzD9JK8t5DIGPRwJowajzOooRnYAebfpK5ThunGt5kjGkddMQZg
VwKsMT8YjROiLSIGDmBOmKimyqW4x0USQ/PVfAlDuLW0TPnZn1VNIOKkVuFdO2KT
Li0Y7WNhOvXTBvNpaA5cEAOwnjkeypncKyCE4nh2/BdabhHA2f5RO9NfmLFlUu8i
KXD5s9xkfwj16oq1e9EcZX0upsnOSKHqUpcgce+oP6IM+r0Haxxj/XHNVAHpmn9s
1NhXnAhSWu9joBuz6kLGAFTBYpr20YNnoXr4bBLDmbWZMJ4pq7wuK2DO5c8Q2DKE
A0E+tBEDsevEbnejW2IXvV6XLpiO88vjDM+l/pniS7rxy/ByyEBh0QPfC2hJOLRR
ngIsH/x+HjyjDT4Uhb7noV/IaC6fWZEoxKhZUQ4rqiwPVwNkQXBxMla9b+aMy6kR
KsP7nV0aReqSA0EM3tiuU65qx1t58KI80wrVgubbSbqLlFQHnuZU1EtG/icxwChD
9V+Zg00nOHgfSJ2v9SXdoRFZgXZYTSz9PiZ0p31MxmdM7MW2MlBpZJAXsDaF890o
11gdevYA0K+Be23qS/ZHw5I6PGlS7rpkfHnWdwQw3N0Vtw5SsDHy8qCsgktznJQR
/U0omtfGHw/LlLKOm2q8e4lfYMccpVB9XJ+lpebD/Q6chjhvcAaD2BODiK9sNOeB
mibt/f9cqpm2gbWKdgVcGWw3PTeygt9K2s5IzG7dVoRPj4FiRqIXVHeeXOWacIoS
RfhudqO6NHUZDmCjKOj20+FRpTz5gF7SNPyK7uXztJlKKiBXLnqKY+BCow4QNC1+
u6Rd3A2a2QpJuS29HVx3wKpnqDM1hVVg780h8D2WhwNv2KWoaAMhLusVUPTqN3Hx
GgYqYr3BnkVYI/ZnRnYLY650TTYUC64iSM97ttKl+aPkEUpZK8sB5xHaEHySfyGD
uuuqDWuaQ42LzR5ow0pQjQ08vpePVFpjwHI45FSP9aTjxk2QoStZbCS45fWO8KW0
thorTwqNwY+e6Q5ZKxFC8IghUnQiq+8fyNENFfsSAcjzDubkbGR0GtLrYiY5lGUP
gZxOZtqyOGEnBCK7qN026Lj/mHWJ3oQwPlBjyt/H4T701j34rVR7/2jI8F/CN20w
KimgeuqIEwoglNbIISlbO1Zra+NLF14cizWINJPnCUF0uBPpU5BTUMFlnFSWe6We
RhYYDGt8NRXc2xbXH9hMA5QSQZWUyv+oEQg+3xzIGLWPO6Qgc6SdESvKOiJT1eAl
B+mcc5k1vkOItUc9kk8AIcL9bflUTRY+IJJlWiPC74ZxQ1VfqNjKGu5sc6NKzjvx
GsWlMwU9mt+JRq9uU2ZaNIe6x7PbV9pxkquCUQ7cxuvfPVm1eheNKKNf7G6/y4qX
dmQgtBK8jKL2QHkjuiauY4RYqPXaDLipHVP4LkqHjuBqUIrO7knjgZt/mNencXfh
EZMT701+EffF3DPQVpynWnqSpH3KWFSIEOV63gp9r8yvGzY3RTIwso8FSg/qSvyi
9ZciyenQVQ8Sif6PkKVOv1C40CX3om6gzG/puAKn5bm87MdT8luqaOCya/4WH797
FhtRb84feH/NAIK1pX1mYfmcEMsCaMmjshB9ssp6yZjaFePdB3ZoEArqUxYIpobH
v9vht4gv+9boI+QiaJuqkPnMplmJaO7v0ZMsgQaH2YsrOU4NlQYJv1157tAZ1Mk/
KYaWnbrRHFqtDOluAamvQRbkCBoDIcyiF8b0wwelC0XK9f3mQELT4XcYqrLzxGk/
6sjA7pTLYaH2E7rwVDMMQ2yGYUxnyja4cUo53uXO0DQplXdt1TV0LjFu/q1Cv0RK
7bPxiWpUy+s+55ZIvW2/Zln1BpyjvznYJempmNu5NrfOPTpU51JFRQVRArcJxBxo
23Zra2Bac5lDu+MXSwlBSNBfe+hY0GLwLe11TFaE5A3fg3WqdTqfTIK/1oU8jhRc
QsLp5vM19fYQiSVO6lMvNdrSX3jzh50kMRpHJn5SYtW565bDVNWtdhAim4grbzZJ
+aoqjdFJ3Bxo7ayIPIFIDX23iwMNAnBI0crITN3b3UC/RI/J2oeOQkTea5gOJ8/4
TGo8D1RDqxGOH6PIOchN0u579ve4gSJkZyxBFaDzVmGPy3k4NLm961fLhMBXy61Q
udXWLJCKDlX0YEA0n3S6HnAvo9JCEP8Qn/pf48gd1zsxUe0Tq53GKcC7+xs+TYlH
/Azzqi0FooDg6csOBS4hH0yJ+eiQbYoUevMWw5nJ8PBEPaRk5uyrrcyaWicFbELm
w0BeWoYEFwkzYIVlOd8XlUqlQnfr6aExQBEwEh63SmwYzaHh67N37KNlQFIY6phV
2VGitEcGYkksn+u4Heb08I9f2U+83rHjVoROFfk8S3ANjMXrGwyNCEEpjUqZ22ly
pYFPgaDjGvqk0hadmsTXGMAhdKoqUcLq0m0nFuL+j+Q8CnJZTm0Jb3b+H31ssrom
qP4crzE/73PFgkTs2AzBzdiXF2apBmWlUAkXld+LkJmgylg+V9A8ihspyvqZB6Bd
LMyh1dturPR/sZXnAV9mPXBeBVz7+adjXyjGYxYxQvnKQJnCH6rfAXDDNTDbUrQZ
E4UvLbs5KYVYwgKnNIRPxD8c2fhm14yKeaTUB9T3g9iIHAMB1j5ZErvdt3NfBLJP
bnH8n9eyhHZgQw5A5bCeOvQEgBy/3ZpEjfmg8Qsd611JSLFH/7vv3JXEnKE+a9n/
Vj973Jm9B+BfBYoECOtgZ4JlKiZ0tXwXXibjkSqOslcvGcBgFZtT7ksXpHVCZoMc
X5XHfvv0wsTBlVZVwgl4uolzi7Qst+0PgX0FqDTCCFEh5XLZy+g7DOLNOP3rY5q2
e66CVcPghenpYXPn7DxSxdJf3QBCtjJup5XnqHeiiTZ8OpW9vlJYNoXD+o2YV1Jm
facvacLy6MeciT908euwitBkxudqMQ3LOoKHh9koQFmkYMKBdFZE2TcZXumK/T2H
fS37mD4Ojb3qZ1+PelplxGjylezrLKGCxtDMDunpKv4pPIrl9uSVrUqQjX/u7LKF
jZ2OMVvD2KODAR/bjgjlc2Tl5ArV0ueunwHOYWjOb241r035rXpcPbOHwYQsS68c
98e2A1XMcsv2jR3TmzNDWM+qljvS6tDm8eyNCXkRwEGdip2XtfafT0XKA8R5fHYi
Hs9EvY8V+ZMAEQfEMw7zR4eyiuWL7aYCoiQqSzLNtHN25Uih+/D7eUS/WUh+edYe
QQAqeq1BiIuhmM90YMCFLlhKKbvhdCtf1ifRO8/3V1aA++nkcVsbt4q34Tif9UgR
RrbfmUx4Zq5bAsMV3xb+xoL+GuVaxHV/ttG/ooKTBRSgR2P0PrSPLxx2c+asGunW
VNeTNftKDIRPBOO0+L93u5JiVtTKLCaiSlYrs3/oIiEa1c8ssKeucP3/YLWIg6F8
gtwFbzpRTXK84+iKHWiJz340ZP7GKyx+YRph5rTGgwTQkLJa9gCmdorCRBCki0iI
PRRRhYcsLt0mClbKz5/M6rcGGQXoJp5zo86gYIR0bHpo0iV1034mP+LYcrsuadS2
ljC/fYGgqNqPK2mEvQc0iCL3BjjMW0lGA9B1XZ9kizPdh8F3ct0GOlAsgcQ0f1fJ
OAljPexe5tzo9WdeKl/9WPyyTnHbPxDjxLHuotPcvB62vGxHUYrvTPKnlIRWIYyB
Kb1qlrJnSIM+4Pzt6AXGWYJbRVHm8ND9Ui9k0TqtW7m+ZJJN+efdaRh9Wi8hcgn0
4flM6Bq7lFUZrDFuh8XZq1JyxHYXgGym9Q5qxIPNtTdb1IqVIi7vcnZl8STnwSmX
u60dURW0aIoavvz8C+Oe+gbSGbKjQsH0HCcPkx8B0zcvSqzMlsPFg9iCQS7cltjE
N6Us8U8mcXd0YQ57jccOhKeXkZuSL2y9kvTdMkZJldmKV4pdobOf+MDlZOcE3aL8
nXZN+xylhy9ClLd/LJRoJjWFEf+1hAmdE8xleCXy24VMbmJjmKoNYYw89LbiULYF
j0r/z8lnImHofRlC4BATlWrfBLCkxvPUGZB4IBq8TyEOBlAKHQhysHqYQxtXxyIT
XgBAJI2IVXIn2hBVgfVtWi7ZwkiI4rxyrU9ojFp5T/3DGttiJ1Mc+jNdVBuSM7jQ
U4sZA5vt28IwQWMsf6GLHU+Pq6ta4/DG4i+ElZKb+LBQPwNekLTJRsvJYkDyVcSB
qiNzNW/4Mt5XGHD8DBIF3woOzrcDINSKdahiPvqHGSRWIv9Mni/kSakd9J4+ckUq
w12ZkMFDKrHMFqy3Q+JtcA+hf1X3Nwhvl9bXECUih2jNd9rK05r5H9BemLRk0MfI
6A6rjs0duRj4F2Ua+T+rj4XafFpTu7r/VGMm/fWEmJAat8wb1Wq6Kxu9UF53utml
vyCkZYk7lSDzgdM/g1z3xPhgZUvm2uD3ocGgerC1uFOimwYBULGTJlg8dvcPn+mu
twKJDZbcHmkEOaR/9xiQcpQSFCOr4goYtOI8wMhsT9+4ma6DC5HaGkgeDgvcDdoe
twJzR0MvzAkZVvionRHntO3KS7gn+3ER94jj+ZLefUOxyjlsNPryPbrUtss161nF
tpYbczk+P2ZyhfAqt1RBS2rpEXQ7YX/0Dkv9TWhgKHEiYU3ZIdvKlMLN/4/DsRQb
DNxBjgSeSvhLZ1GVYWpXEpJFOdd5nT8Wj3NjWmQLjuIIaER2AFjq3OToKSOOZajg
2NouFJbb9HAyMsOm3qNFcnagXHFtguYckxHNP/OAtPDUTB0lfflABajKO2HQ+mGt
NY0UT7ZgQtoeOEUEkwMwvbLNGie13hmsh360LtC0SXhpqUP1OoU98/DgJjSuf/Eb
qJTW2qYkSDUD+XAOUvmuvP+oUKKqc+5L+813GBbo5+0u8VTLrAkRQj7tG8AbyAVO
X5P8P35VQxbIFHDN1BLOa650uPfrb9WvtV5nwKl0aSwY9oOSYSs3+Jrny2Dyrh/y
3PUsuaxBEKnEKeWsHXsbc1sGk6YMshe5Da7qmwct+DLdERjNHUb3+8ra0Vl73f1Z
xz3tTJW+4RRCXBLcHdnQ6ZmjTMRLzE16uYQw+szWWTndBe95pti9qc9D48+t0AXf
lASSFneyI0Qpmebkqoi1p+tbKYW2J+oEMGDfDGizMAQx9l0sWN2r/uMXlJY9crGG
1nGeHbpcUT9ZpNFpdlzJVw89OF5kGyycWtw92cyB7VaDFdW6XrGwlVGmfGBVasvh
yjpDW0+AiMEJkQnPpNER59gt5ymtdnCuEh2DcWD7pCwUPdDeFrJVAUKBI6FL5Dm5
QXpsLwj9eUIAGzkROyyNjPtuBSq924OTCNUawXbPDvstaNGxzDVtcdoQB9oOpQfs
bjCv3+6mvOPJVSgs5NYuSUuA3zPRfdH9QwrjU5zHr8+VZFWiQ3tl7gVttfKVuwrf
EfYhr99nhG5G46I7oAFBG63n5KMOgKsnNi7m3K/FUynF+BJMH8yXeKAhh2b+diGI
pEzLTOzOcG8VB1cu6GvZi66+Gw49IBO08Fc51VIXAwsJqe0h/63SU+ZskiKDeyuG
3AWX79OmTQaXuidTxMI/AKYBg3U1+JNVZVF+S7UgKoK4UYDRMmqz2cjY1uGT09bo
xJlzReEvCahLQuTL5i3lT6WFfX6nTTRo+DVzHfWLcAefmH/CL15exfM1QBGK2pCn
5MGWfoL5iMGBj76rzm0CdKAb9BPTpHXHa7OGgfRPOSoCzOyGS0VsqVkmMJzeHUja
DQc6OUhqlWQx2vePMrEbzX8ql2KtUfNuXj449padc/BoLTDZ0Udl7tuN4dHY8Dqa
oYjqLMw/IzW0iumFjjy4gi2tt6bo/5QVnWMkzKSs5EVZOT/lmQBany64qsIEA2D/
5vlFnDz2k2oEdbxEppKm2W0BtqMokDZtv6pnkusj4yTe9fWPHdlWYEqgFzXrRGUR
Ynq3R8wrjMQzpgEDiMPyEUcM3ucCugnQJVTB1sw+TXUcAKH5JeLmD8Lmayl2g/Cd
Hr1p5S4RRrPAXovi3L/4Ep/+DEdzTLe30Umxu+G4xL737cgAUoPC4TUWc4fMtWDX
hcCLPqi6a3on9Go7eUPLabMFb8mp1ADdWRkOX5zasb+VrsMEfRR15Wk9uxpH+KEb
l4nlYwZPQsniSwmGplDamzOZVg98UjgdTkbHGRuRYux7f0YdDxqXFotFQHOo9IvZ
O4ojEPPmonu109DtdJyDkUn4OFVpu+5zZElWr+t6xVfufFO0UJ4XPApfJyh/N+U6
sq7XG3JQuPZP1c0DAot22rbNIUli6hA3oVNSk6pU9VGKT7pxOA+Au2jyuvrn/fio
707FqRcv+EG8ulhxk0U1nQCXLAOgMacAF6w0Lwb+UZp2XU2cFQLXaiNFJYS0R3bQ
bNgZgmoXpAgkMImWNmrI8VtfAhqUYy897mDzuzt1AmAElqA5/AgA6JnhxL0XShZS
gHbYaB7QqLhKPXPWiBGUw1hy0a6ga49o+cGaCDvusLXaBYg91UjoV51/YguU2UZZ
L/Kb+nWGa1+Oa9Tm6kRUkdlk+Ub0Vfa/8xFNt/gnaju9F1I9r/qyyB/2Fi3fqmb4
9bokqpr7fABilo7sqE7MBmB45kJeasi/YxMlCDr0LPvajVV8ZuHjwZFoWUMpTHE5
+SRoNKnxm3/aot4AL/XcC7mG6ArDWMkszeYUVF3tjQwLeZknyGcSKAcWh4g7mN5M
w/2aox7+leHdZe7tKwlsoFhe7jOecfnodQf7RbeQ+Bo8bXzkeR1cCzHhlPUaTcNN
feERDNZmeRonv0SCGeQ7Wr9SxfPVMFhCY8jGfYGBLDj2mOIrpByJ13BiLrmkNgDn
MQQte9VzMrw7Nz9oJlRrGED3ZbXsAFwj/pHW0OhIvAIjHP4Tl0QBS/RQ1WRWWNdN
Q/T0fr415b4MgM6zX/aOgfKgJykJgcN7OlxFdCd0GcJzIERCkG8R3mBG6omwY2wm
zTQiOee4zwQIOp3dLSFpJYk8hYdCvgKctawUKXSRkUGqgtooMSJfhDAAHDGQtttX
JyGHUec7jtLvE2rEkblMKbdXkOer8zk+CRQ74dZvDOfXe3GMP5rXw/AcB+XkQD1S
tuUVqGE8AfbeQecNbwMoXMLQ3T45nqQrk1GiWQL59/D7AjN/GjH6aTcrfldyDmLs
498/DCgpeSqiSNyFzdj64g9S5g8ojgAJvQJFvEcWTmLaLwAqHViWdtW7pnNqevNH
9JB8dWVxLR400CWRLa74rGSLt5Rhc6U6sssfq3fokVhUsiNI9F96UNgre3QaOqTO
KBIyOSm1UmthfYX1cMqbykqaV93xuJPXruTqcJ0l5MEj8IGGXszv9ZzQUL82Rw1B
9YmkWRrCLvWFpmBxj5DvUwvfjbzNOFP/OwMrbl9oL92M8FjtShVXAyJ6lddKcXeQ
zNbFb6eMfY4TPiL8p5wRicsFMqtj04DxiO6wzZ0tAFq4CThV0JkuOmpoINbiwscE
/HBjuAe0eTSv+olZbB/vZU+NzRpQYdewV0wQuVysgeaclVGWWAC9zCHVykHGNNux
Ya8IkAIt65d9g1EDfu+7c8haKm+32arwpqpE7b7dSL5n+l6RaqToaqJiCKvx/ExS
StJ0E7ZWosJ3cbAKwHAjMElyH4qL/oajUUWNr4pA4ZkxgWPa38cNowfpOndZ39CC
lGsdTQaC2+XepGHdG59Ru03NUpo4R6MfHHX8gp/39/VQdqDmu5ILFb+XiMGy7lPO
cpJio2Y3nS3J4IFqHPAf/GLVrlA1C0GHLWLtbGhSE/ECKe13qJfAVc9iVjQzLZdt
oHfYCAyTeZKUWr7+Y+pEKlSIV1SiKvhIg4bkUGPpcqN4mJCEtGYZndDkhEsF3HE2
KQitThWh/LbOVO5lDXyElnwc0QKeVQhaZJRSzAcymvWResrQQgLhUOox9hs8MFPx
bPVBPQNA+YSzI1ChqkRXgN3heSFp6DfJcRPr6rda8Klw+WWHw0x6FZz7Ivb5Gsq+
rMzmMWhXqlssSgeAARGCRWeSMSM1RB/Aw3YD7G5kmByKblRw7wiHwHXPMuxvEO7K
bx8Uj9SZ7ILzwEZqenXMyBJseBgMoKKTQJw2JfC56iJh1F02PdwSI7EIg6u5fUrM
sSklL951bJ1wmzQayXxtU39UC0GAvIo6fw+CSjkvQKAkUeRmf6dAn/JtqRxi+9+g
s/+PEgI8AgEJY7oyZrSuXL0oGbqVfXPrd1Z7P7rW7VPhBFB4Lr3Ik65qhJtyiCRV
f9kQDKpMRrMxabniLzktGWa97coCxDCiO8kfCaPYQ7V6FLGy7YsCFtt1PNgv8mdc
Y/VOqQGCt1Rj1fCSgd1j4mGhcgxw++qVLNOwp8MVLdxXGTjrxEgYq5BoFqi6N/FC
txpzZKXOtH61NhZyd+uLn87c28ZVhYf6Yq9f5Gf3fK4qJXxu+CuYIu/4Vt/qD4dR
5WuOY7J02suUqBlHwrNQWe1waZH7nkxNAFwPZSteQeUNg+9y3TLDfDkXBFSJ5HQV
G9/IQRAEIpuPKowrnM/a1yy6IoEJNOQgOVyU1Yd46/B/BNOm4ktNK1kK25sltsCF
KEjC8C31DKmKXrOUYFeYy8Th5KAaFzmT4GUVwY3YVFMTpI6bIbYlqe9XnhGgJed8
cPBi/8jVycG53+DLjiNPYwNf9GOQXsBd1wqWtHdkTQ99N3+YlL/4gEnOHZsBeXmd
8Se+yxLZ5OQu4LVa0hf59mntpfFY9Dg2vDUPoOUoL7g4yaGIDd5pqUN9v/+EvlQ7
1GvDmmxgw+8Hv1cf+FCRg9l4CgRUPL8gOXdH0OIcQ2wPedKs2ljKNnkT8BfEE4bi
caY4dLmoyiQsrxHQDANTXVdodpBAFYEW6NXs28E29338UOQY8ihzaMtTTtwzXrEZ
2IKSHlf2hHxZpOe+0y/VeF2d9XktfEHSup+fasBRhnydf75e0X/ChHXZtIoN7bOj
PkCjxxplIC3zhzl5KgdF5fP4YMaJ3tT/9U2yJjT8Am/tON8320QKWC1U5oKCyH2A
DeyDB9hDFb+GkagIemkonUJZTt+BVqEbeYXmEitURJkC0Y0xfrxe45DNBwBS9fan
2teywGJTRQAnOc0VDbTltXY27UsRgtkcr4yE48M7Yyd3FScVCSWnfKNLRvk9KUcQ
HIE2Of3bFcnl04jSnm8pilS7s1SoW+qEsGAD0Pgi4wRSZQbeTJSt1zmBlky14wDW
rkEbcfcwqd44KvoM7WYyayoAbSaCTgjB4p6OzUvm7i/QMvIO97knQpycMbHV/fxO
dxGdJC0+vafFQHfbyeR+P5sK5cE6ScnWSWcOc3gUX4v0HhsjzYjMJ92CqeefEaIK
9W95VPy/Dk1TfKkFR1I0G3kkfbOxdQydpI4vN93a1TkL4aENV8eSqHpzt0w2IkK5
D9Ez4idRC/3y4uGlWmCeuDmpGcp4/0qup6uZYIslY7vK4efWjqltjbVZlkl+8RAL
7etgXjyLgJO+Vk1Vrnjb6HBQ/HaurVyzDLYOxpohdUB8+OWgO3TUhqJnFySG6IYL
LY63Dfc7NMdvXgZOOXTpd6u1ODHOkUjt5jopEFiKk4pALyXmZlmfqWs4F/QgQbmZ
zdSyzjL109tWc/9F5xnRj/5Xv/RZhafu1CQGlC/W/xTJGZqdjaQlfakhfNsMQCv2
fc8eXXYudvYjCrKAspPPaWo67vrT/eTJtlUsWQZWzPG5XHMQWsV82gIqL3ONSVTr
jLGfebbmutYiaMZH47jPIFnmTyvV9twsbloGxP0u4lFPWCxECcZCo249FNZ1UVJG
OAlnNPfdDnarZzwPzkERk4btem2x7kshFSwPU0sWpkHnm+84CSG/CmEQ+vYUMBLG
91Gb66vkPOm0fusjES4RSNVdn7KupEzvpp7bKXn7CFtMomVdDmGg/uY7oqrp3Gnj
UB3WfbTisuv6kTtRQBaz8fVULyJPsgQYhsiE31aicmmFtbS/FRTzqV5ZI+KwudYb
+FfZLv99+k5bOZC9ODxk9ToqB6Z6mg9iQtYkVuWSj59wdxBeGI7f4igvjK7m5M6n
MeX/m0SGDnyCRMNd5oZZtxRAOjlDu5+atnNXbCvOi62atPQgE9wpNMHmLr+0o4uG
BMKcWeaKXdyghKlNWOItIMgqSXdOzXIHraR8aqJeUj+XtpfiZAd1NBe1P3E5cH9Z
rKigCWifEYn9XM+9X0XYnzhV0UmezOrF7PenJDl2IUkvTLJOd9t3JWlkImC2BV5y
jZ0XtwiEVK3rq+V7VANSks7qw3DuHoiYgP95SOvWkIXt5YmBleld+GQq2ppNGSV4
EgvfAg1M7lOn2mLmxYDVrI+teVWAjm58nPrOhoOoESlO8t2Zwor/HImCr6XnqNHC
uXoUZYNJQHcSdw+wRsw1BWBd1uCVb1lyZrv1ArhSIxzEogrSWEq5ZBMi1s1aKwNB
JvyjF5rwbahekuTN5FZZLjPoLeY6tjNoRv+ijJlKNlkooZdCUCdaQpJj71FxaSG4
iV8WNUemm/EoaMnF+dfxRwcHaSfD5PufxCgskwLTfWhrIDte5MKu9aQwqXnXsE9c
mfSQsATLJ9yc2q6z/CrVzSTyvwOiyih+Xvxfi3LssP1eEazo9rwjOpY3pUxm0RFS
zcAll39lE3Hp/f+h0ptP7tgNKX6onl65mBuuC2l4msBbv0FXN/jtBz4enhRx7xEZ
JRSONeQdK65cnjYdqXqtaucQznQPy8MMpaZtdh3uUdIz4AkkIYk7byd7W9hQKYC+
r6qMll9SGbF07KoHGjpIKxvtaBuA/8h3Quqet0bSVZllxyX6Z9VLt4x29G31JEVt
CeRE42wrCQmvJT7fMr2sVzyxHAxPsyZeUP6AZO1NpZOdUXTwU7enpR6mdKy/DW5h
hc3Tx2hjQBnBx8MWIPiz0yYSAUyQs+AS0zKHVtP0V0DTVhBQFdqQbNGxLP9UCS3A
HuEeGcGjmABciGazxDfLGLHDu7nbmYzEzDvY0MldV52YYpNynqoVbOL7T6vQs1hb
OICdGacYjYzfGJLAhtdcrw1V7xwEio+E094p8Rt3tuFzZN503vfeXj0SS1I+t1mF
Ad/WEr6KF0UBnv+fAyVBQTI+Gv0C0lPyLIYjFyniJxYmHBY8RHV5XNH5cI8/FfXE
VblhVhvmxyvSDyPEcAGBuUiGr12PQpvcRP29atfykeDSsSb2LziyqO0KBrF+N1T4
wVmGoZN8S2EjOU0iDjIrJcYnXPNkhI6c3NTlU71GqPyEeOxBHp0sGq6hGxNrLhRs
xOZdrJOP7yEU6Hnj+2vOErcggFQydNr0owxpWflXtTBLq6gl3lj6p+tbOQzJp2BI
dKZ2UCn6l6WtQh/GKai4OuR/ky6pxET2oR1AkiTuOmb5218ukjn7Gj2e56u61M6m
37TbcVoQ2cm9rIcXGFYRik7KAFLxyHCAb2th7o9LG7Fe+uDGSfN++UWFofqbZg16
fs+MfPi2rCQBJLLGqFY3uxnMzZLoWRUASgZb4++2wEll6GhtEFDK3gZb3DKFUy9k
p/z8gPSNM8Gli9ulJhhkAZ+BArM7fvU8PqcLT6tXrU4Oo9LUnz2NWTuIER8L5b3z
qEZGMUa5JpTLBRjVGWNZ/mSyYtGYmpZn5PFwbqNKJnH8dUm6a02mS6cK6T5voEzK
Rg6N3tHIQWJ47T9CkRSdhA0QpnxAdLAfwBzre/Qg8vXUbduOiYb/JdIy/uaWcxsV
LMwL+sSzi864uCpKAyiwEivn6CC3jxfQsRi1WvRPF/v5dPMkk9EipDjIXU98qrJU
lyuvwOnntnxt42cdHqI9TItY1JA5ZmElBWHDA0F+PKM6a4QxbIpuldfyRpoOsI+Y
eenhou4VUsR44qP2R/chavvak4jpDAjJVBZNvefoyIN+QTEKl923xCRFE16PJ6Ma
57freLkHGA8zRtxLAE7oP5HaZrjt3FY+VRlSM68t1I2/9PmI+yG63vwwF86vEoP2
zPt2i6WYXTgWZNhqY3198x5qr+Q3S+pxekVv01t9ImkaM2hYdAKIJfDSmvMNQ5JA
LIGqggVjn6Qv1tCISLK6nUKGitS+S3e+a0txBFFrfS+oAvOM13w3gJWetzoxQImB
tY47cyPxCDWBeBIqgo3OjVqap/r85/kN7H0lJPfpxPMfb+pEKwv3yTw0P1URtz5O
5hDUNkZX4Gg8Lkdk34yBcyEqLUck4E5RJ0bPOfw83+VtQS0WB4o8oVZ62/wWMJ4d
4UxwYfHcdgycal2Sc/l3W5H9qJc1yv1CUmKwqmp3MSwXkf0jA7vYvK11jRiT6vrW
cGvuEBId7Ouq42reQdb9MO8CKS9dEw2s7MuQBE5lzIPszCpV4WW+ykWJ/GX6bL1r
qQR5u06nepvFwOuMWuSmOb6CGxqh3BpLvjRYqE+6Gv+ZXEzJYJqJSjz5n48fwHpq
q6+CY3YVCvkGiWk4lFREaOZxKzw6zW3K0n7WyHbE+p7FjWfYYYD2HxQ0Dv6k9IqO
3E7//zNx/kZfeNESvqix588CwK1gxIbLXfcBhOoQkeI9DVRKz+riiYo+Yt6dMxWD
yAed/UttO4AocjgXRPocfAgZldy75oE7Gz68z1LzeXuFw1AFHHDl4CTd0tC/2WEG
jMgrX1RunaaoMzZFPknTHLBtUUYur6l+lpPdDPk5LAJ00vHfxDTnhKUBhYLkC0KC
HUEHvXMggERao8OIkjqUdLObJnIgC9vhF/nXr2eib90aQF4GdzzwoAqp+XEr1pT4
G4FMaUt4ubihkJba1qg8gbYi7EMtUSHLyPjHBKaDIrZ2CBj0FEXdeMLG103xthWi
uTn3YVU3S2yw2rxoFcO/J5vZOU0wXOYcnpwN1f9FbcaiYTJ/MhabBVQcgN46s1kv
sMnmLtjCJ9yvYiO8nFp3i1URd1LyOcrz4TxAuflKwyB3kiLxZg6gj7DqGEpC57YV
Hfjc7awRaLxMpIPAif8cUs/IEsoWFyN+r60RmA0sWV+jjZrGA45/QGP47LzoKvq7
OHyiA8jwzxzfePULJFmzzjUCIDZnoxlUPZGbtj4gTM9MfCZSYhavsw2sGvc6J6Ag
GsTJLg2sWfr0LRvsqpT1r9zPNMuu9+CcHMxrP+ZfCOHzrHMyX1U+e46SIXDrYk6c
AONmIredj9U6EFWbT9eu2xQBzyuJmEpFHlplH3ejpS+b7FblFgk/8EMBsMQUbVtK
/jfh/GN82qUvUVTuVzwGFrbpSggPPhGEULOEozGKrwvMBK1IYldVEhJUavufeHoG
NIQyiFh9mFukZsKGHib1+4pwFUcj3G8b25K9ptqLzLP8tc0aTpv14oez650A712Z
1EGwwgTjS3aNP8rb5l5fDCkcdbBMYxHy8TqLzjY/cHWFnj4mRYA9yvohaDsNp4bb
XbQ/ICxVnf60CEeTWGdx/GAvlGZ5CWuUmeT1O9bz2JL1Js8vi80SsmD2kvumOioU
yv3dvK6GAD99zRIiEGzH6YBupHxUTAX9BDuG28GTFayYtGes0YurDC6cE6f5cdbI
n4SQFelrRpBG7FUICH80nH4Q3UUb7SldxEauY4+GeOF9ELxYEjrxntBPljXkqW21
XZmlXuVINwxmW7jqXWx91TkrClFefAQwtIqfAvwNxHJSpt3dZTyXYGIOzwVaAagZ
pyhz6lPWc2bbYnLeDQXO5hb7gIAoKa+WSW98uWfPutPL2CGvw2Ospm0SqXXrJe+d
/cR6j0OhM0G01jVSWQ0aeqt3dCAnUMGX03V0JgRVQWo6e/uWCjNI5He0Vy8x1TbY
h9u5nD+e3m5mLdrTTjYV68CDshekJZV3h0jVq7UnuewddgNo1dxsC98hFkuMiqgw
MWhEm2z8RDX8xPz6y06mMybJ/fNBa/nMdkl970SsEBDxtMM5BEksQb8Te6iko3Eh
TbuTYmb0xLnNt0GcMqKuBBIWhdAa0BEvT5TXDxfOX5T+/Y1xdb7QjDU6yMWUbp4y
x6iZVuLR+eVhhsTvi4StJR5IM7CuX0vSpIQxH6bV0Ikb4FGbguhVnRqFYCFLHdvn
Q6BJRQzGB3lIqzFexvfWFlEZv/j4pUkgXPBOxGzsrIf9XSfNCfWWe1/eL7/XwtEB
PhKAHMxE54tc9X+By/A7gBOVv5djnl0cTGB/rcnosNS84SQKAd7uids3r+T/EdGS
wBBAVse4+gq6SJDyKxUCTC/90WAcQNi3wA1gDPV2cWIeKQ11Y6orrd3m1LV7UJt5
3XyHjU2W9UNcCgJn0EUS1ZjKVV+MzCWLNakqhLLd5FspU4OOgGxTKTCuH+KTr158
LtECb9CefLR8gcL/9G+mFW0V6esysDRdFp0IJlzVwcCYFLvaoOM8gcjWSukYKVTY
KYERprV1oqZEAlmESfb0PFKp1Rf4Wdn9Q6TEmmh4AwQaKzNfGmacVbLK5BThVsv7
znWIvKkr8lBFc7QMDv2gJPy2tE5R1nVlLtIJWx0IOsXdU50RFrtODWfrPGOnqaKl
vWIPAA9xiX+EqZ8QaMBJmpoWnyzgdRzR/rc+/7UIVuLFaduh+S4WlGl1Hx4m48jS
5WSbVPf0VuXnL5gCZGWl6SnMkavnw/YEejuCgBV4OHY0JGSMqjBXy1fO7clua9ff
tLgtrW963MLMMcBVMawOJSqsSjzQE3uP7i/t74C195H8vzXLuVevjs72RSMVYx45
/Z7qv2XFYII1xO1iW+Q0NAaHkdhtyBIDX0OVNm+f/Sv9MVA5LSGuv5X5W4NZTUjx
cCrFPP/5PWbkQv18NmaDvTR/g6HsyHEvw5tBDEb/NRloVzFOZHGBVYRwaOlyZg5B
j9xdAh4QGPBcN3BEtxA3Y0KHo7fJngQ36qIHVsKmYBNu5o/cXurRLGBBOQk+s35N
Iv+49dLPixfzbYCVTrchov9VzpP+XZ301ecRhI1mxhZq81cLiVw9DOZTemTSMDCv
BJZDwi+zSJI5NIx7ae9PB7Yx/onXiY0nBBw8AlpU1MOdEyFmXzvRxEmFoVMtMCRz
qRFpiFvsQRBNlpA7nkRO5qTO4FLZn4e/7K/BE+vuuA0fhRx5jK0tBOufWpiWbYlM
7S4vKrc6nbqvKMG0Lv0dVbF0IOKGUC6q158Va4moxW+lDQfTLBSF31E84TnIy+RA
9jtqMOChKtzUizYuiWabJrRwZOb7MA+zGU9E8sMgKV7AVjvlb41L2cCVD79n5E+E
G1/0eTpCLU7XCPm0yNv1pIOWio0t+swpKCT4ns0MyfjMu/finAFadHiUNyle0SGK
kpHfkgfrZawiMyyUg41ENDBLLY0ikjeYNjvnl7xuu3q7lypNTh3PRYt3Xg/yEtwi
uJ1fn7jqvSnTAyBFMaYoWtnsMJtBTs8Eah63b5BRoZFko+K9a9GxPaW5AqmOam90
zmeE7LD5owyN07G+9PsP6xqQ9rePH0hOSuQwBWPZAU2jQTkk21VtwY/85OENxAjP
JJlRzHmZqmt/4amLYSGb/B96XoLwxTDJdyv1QfRTUbBqwa4k4Vuv6vRNIxqtaP6K
wGAv2i79kjJfpQt7Uu4/SAVWZjvZm5F0jIJsy95QW5v8ctMzVjzzxeRo8LKKwEJb
XMKHWCnFySKsLSjoRiVRuN9JUMJUQ7nNWnlEUR3TYL76Tg4waEqyTMz1o9dFpHVd
vrTRcNGnApYnk1pqrEJcdtNMUaFUBZu+pSYdWAbdKKBC/xzhC3MEa2lsrGo1Hu+K
JxkB8InS2EawOUEbLPm/M9gh4t1vHb9BtBCsMukdpmsp1brFndpM3o2td8BZzeXi
RnzGGxf6mZnT7RbiAHfKHtIBAJkEvzDz1+U19WnKK2HqNkJ8ENcut+mJK+AhyMA/
NKIIjD3UTKF+CEGTHwjI5MSNPNJR6H5lJQ6BuIJ+lmlmCrd4ntrnixqx6AmhxJQV
2U59BbgdhRuJiZqia5TiHQP9Qo79azAdMmuuRpaM3E83j5qfvO8LgKUzPmbUYaxF
3d4MYo9qCzIdYRETiM8IUSn0aGHBrHgQQDgffne/EhI2xUKm3rfhZE3bHT7y9rgr
7VHBoskMhLf0x1ZFAWVwjugX13M+Xtp1yOxESJOGRHehOtmaD74rKmM3hD/4kq9o
t3GUULeJ/yK3TbAvhBaLB8yvdVUgZ8860P8sKzECR5dK5yu6SfXRwSibvt0qIMsJ
9PX0JF7+7kSL1YKFVkfY6kqBXOh3ZuEFaNuJRHJmiJ7W/imVaFYI1k2JS42GBVPW
pFLhSQxwoR/japiAJYJYyaw+IgNQv1hJIoFRKJPXEvzAm+L7CW7aSqbkVOQ5CtZg
VtfLF65IwXM/IEjUOVdQW+59s0aADBu463SUSw/cKTMEfaENBjMrBsI05AKCe4kT
kiuo+oGxMmHmwfZLJW9KFEbQVkRs11HbVlog2o92mgRIUmqFuKMdFP0KbN587+AN
Whx2CrJsguCBg/bKahAFHL4u2gwXZhs1eAAg8YC6QlVofo1pu7YjJJ7vqADK9qqg
rqiY4dvL2T4hXzLoEDB/RXcT4HpJ58596OAx9g6ayzyN4ZW/42Ggiml/F0yhfcK2
fSb82q9YkPP4G1Nt7Cl8HNNr7naviHhQpQn7oZRnDHC/05wxXCqIgaBticOJXIok
MjR8uLVPxu55R6cK4f0fG2oCpTelWt5+tpAn32K23LR6OsclnKa8xm0xCJbBn117
YRCCxxkzuSrJ6uyQx0cDXFSRQxU2bFfm9F3uZwy2d3rwLWHCT2UhuGzZ1mBUsKwb
i/mEQ+y1eBCf54aLL2/Dww9Eck8TM+FX1dUCiw4AA5SYaDG1z/pIwAlSHO6aljSu
BSbaZb4kyK+UbBCjeJaYbRU/pKiW6IgXMsBATcMnpxt85XNhFxoB1WFfw4FLtSdK
IPQgxq6eO4LYA2dsET8uN4Brfo4umtXkdd0vRyjtaXEBkyYeBZ0B68jFv6npZM9R
6gzi3kxMfhpSEEyR7/qhgMpkGn/a+sVV9OWkwPgpSkp7OxbG/z2kZOKuiXaQKEdw
2gq/qgk6ivXqgSB0T+1hVpKxqF0JOc3K8KGqH6itPH7fbGzWak1xYerCCJbziPDi
uaYHJb3a/LVpI01sY99T+3JumDUBA9+v8Qdvi0QY+UzpAc6XxGhRB2Tstk0ZLU+8
lbwGay0FednGkV0m02cujDNntrnTgPV+KBwtnk4mZeFzG7YRMjPtsiCetMphyZd5
YyqLPFa/qoy2YBkHVeg5DYwNepC/aNjmWRzSIx9qptViLvOi0LnImO2ytoQgdLss
f2QidIRYm7wh+PGwZYE+DKku6+7seIHx0gur/6C8oLyUShJ9B55SB9cnwpBPc9T4
pdz2NER8xceViKhoo293tDkzLGV90wJGZ8tQmosf9yxjG4vcWdk1fyDLsHbCPoaw
2/TdywA1w5EUDJRDZ9UojPrFJgT1wsPq72thFdn14QzxD5ECjgkM5pZzPPvBVt0a
f++t/T+v5+blm/Kjfd3QrySopahjCLLHgzJZxTaor3FyUrznouAjZQbLFTOy2xtT
pnl4sil4wbuc5BOU4bnC8ovDJ2xtBC93zTx+MTfC9Y4Bv35m2c4oIkqse+3P8Xpt
FKWtTMpLAFtcSDFl8SN3EneH5pAln3nldFKABQlZz5tav8md+4YhNyHcF1k8U2/v
0HCc1t3uBek30oVeBTaqf2s6EzByH3IHF0pC/+wSRSpBCK9KuQXKIXVv0KgvAxR7
fR+iLTHMMYD3YLYSUScfryTIaEeEiv2JW90YMadF3N+VjBLYWH/xeJMQm55U8Jx3
7/MF5EjLVzGSpBEanpZ2t0mZd1m9BREaJwEQN67PjRHQBTzouf1kJwsBgUNjN2/4
dIPQp5dO10/ddejbXst6w9pwo3OIBWAc6IHVVypknM572kgvHq+ad1Y57O9y4AGX
4CNiqW0BJ94EtrQ9kBGsW1NggsYFV8eD/xyTUddy8brtPC2lDE9Ryk9TfGZawtEj
lIyj3GjmZ5SpsVOO72qBS4ueLB8RApvoCFxLBttMuBMm0ts2oXyB8KHK/yZE3KDQ
6vuz1XRTnkPjSjY2bn/RaiExnUCVBDWaQlMzOBU3k55M3bqc1LxwJc2pVmWd3Dwb
it/XTU1fltXRJu9BYv1pcKD9YPwlpQIXCA5kKOgA13nX+dbUMbSgIK/LNjPbvdrn
ZlO21B/6ewSwlfAtMEiCmWiSqR6ltagj48ljUhmF/MGcTmeVaNm8OneNc1iJPiqW
ZbAz+CLleEnyZ5Jyx/nFdSPUg567liD6XMqrtHpfYbagSi8+3RQc1LOM4kgx/Bad
nKz+Im5AIm5O1GOcjIGhwAkcuAGiWi48UJ6X5Q55Mw+YWFBHp50oHG8te4bZkiqe
C6pxUhk8VdVeqEBd24A1d/kAJ8p31JaiecjgFZMZ8pWpGxe5PdRL+WJhtLVYWsdQ
SxNvCu7SWNxCmZP8HjTiNAIDz/a3m1t0C9F0Lx49l3XrAj31hIyj67bkGdmLDe4I
fKmilYqhkGyp1+ojyBZ8xCiJyfc6CpZvHmx+dTldI1e/+5NLCyNHYTXMiaTk4nZu
2bpbV6zZ/5Wa9rQjGVDG64FaUfb9UZwhdVps4ZvoWfbOMq8QhNZ6RGmyugkdq33O
ovcQVZm4U7p4Idt4Tui0uj4xeeLBcBh9xzr0VWj8zAjJztl3eOx74SCg9FNgyCH7
49ajvpNBZ+QQ9xNb8PxpyKTvxZNgKengKcI0Bgk8fZUgPNg247MwYBFCH2VmIYxv
VBcz84/Yq5dbbvla1kvQ18tgMnhfhgQTiq4bihh2CyVelaYge4ykiM7mWPgl9Xsf
QfWtmU0+VKW8nRjU7kQSuLOqC6MTl9IAGX4EpIMETiU9Fiswiyu5x4ewEgbfnNaY
i+BkepUfthQno7IM0MLfWUd3v07YZCf0WFs3rrAIj0x9GI0hfBCL7xoIfJb+7mnX
OmiSqA2T0Qi3Lk2AhP1gITEQ9e88TQu506i71k1wDn+2gDE4t+Clh/NBHDNMf41U
OUdFsrNlADKKuu7L8YjRHPr0joMaLZ8U58OQHPk9zLGfkUEJF+lbwK6oKzVif0Ht
RFReauu51esmDClA/cmlLsMHn9XvW5Z5aJEjEtYAqC95GZbpyzPH+NEvSsnrLyAL
ZdRwkJECxxaUPngksjo+pk4hHTb3+tRve2u5/0kBAurlMhG7GGyrHw1uIW+SUXQW
kmg4EFJeKV+rgRgwUgY+tfSDa3PHVCOVTn9+OvjL2Rts+Kk6KHXAxadKCkgJTehe
pdYct1b8vTeTgWQXfo3D8s4HZBVtPz5U1JE+f4pfOe10L33bF19f1H7Ww3tEwTlX
mgyiQ/99S0zfYg7H7MRAqBA+3YxVGXIH52ZRB0IB0tG0Wp/rZcIkM5P9iO8Zec5u
ibOiUBlPuewMmKx+Ta/xO8+xgas7QpezI3n/3p7Vqr7UwhMorOhLsNYo3rPqETzH
6otZdGh0AfdiPmOvJu6UF+SLSZ3DcI9zDG+phV/vd4A6mY/p6vb+assOqhSbSdoP
xLmSuORLpse2fIMFwvztrGmNumuWbvvxEhJOCMw4Tuw0GdDtEYAZqye2j6ZsMS9K
O1F30motdiF0UPp1th+UOtc+cc2emOQN59j1RGM+GyZCMYdXbCEQkOEsJWphJ3an
Y1Cv18glzWxbv2FmzL/g/sxz/K0kUpmzJwaCV2/ET8IRzjUn9sZhuKKLsHHmvm2w
b/gNSlUMC2AmBiIyfnWp+7K19xiqZaBEwTi80uUrunZ/JjbAkrdAVNIOxaMAffLf
xwFYdbMyr/wB1klZR42ESiHSHzHqmsfN7tS/UmgNZfPUpQb8JUkBj0txNCH4cHSn
BSDLfVj0dZYedU4a5FbUDxy99CSxqkHKD1uXFPF+8Nf2W5RvKZ2D7apvKrEZEpTm
kwE5Vnb2L+0RLLQ+f7jxVxb43dhAlqvKJEk0CDi6KPbSqdRzAkDOEMeklpyXr1zX
8wWbE7ASWKqUoEUO5CrKAIrIRZ6FTbGPZzuE9AfJnkaYR/PiBCWCHokdxnyVpDcZ
jNb4BfQCZVCzxtgn4mQKNDaVdJyME05HQjTbW9zmgkQCTwmU+So41b6Y0NX/WwyN
jiLNupcdRWHfLLxv7AbMkhn5fCemethSC81YUY3mGUUW6hkuWcJ1hI8MaiWEKRKP
WpO+Nm7k1Zpwi8RECZEzSQwUoLejKEq2Lg0Mid9LLQMQHsI3p/K4W3upRnQyfUcU
pLJu1wMQYmI0VnDee/mQkvIP4m+9qv/wnenV7YqXwQbcxeL0eSE6wsuSGUB6/x8r
ZKZT/C/Z4MReJn42bT6n+vu3AOVHQOK49xYbT+lZU/ZngY03Sequ3Uj5urVTJh9f
9WEc79I/+F/nZIj+mOsTaDeaBLtKE0/Zmqdd+mKq1N9onRDUlyGmt3/qja0UWK5S
2xZMMSmQH3QqFy7lGEvC4zz7Tx7DV3q7bXy2xiw/w44+x7sjBGsm5yIGv01OLTrr
LtrZGr1INvCa+R/VomNb+RF6M7MZrcg4ywy+sVpYh0zJYjWQifI+mP9Ozwg9MzJh
6Cywkdv8vp+/1KNW5UpzCpcBbAKJQcJa+QwY16f+qzLi5br0bjNNiQ9SmyVy9VDH
BltfhW00XYjE8ySM6uAGXIUUNBNzK6SqKCI5q6VrdUOqRtTij+ToYKL8xN/KnXH3
8xBRPlG9ZNYODEcDm2yYRDW1AffTCw7vdo8paPLXbcGDTK9zjmgCFTi00O6neHFp
9R/j9L481VQZHlijyhqjP80RYJmgDlbLMN0QL8o11grGwls8AgdMFSZOdDsvhkcT
Ezpmy9qH0dR+Srl275OJV2EsKqc2SO9nRGe0rhRmHTFbJJtaHpHYU2TiwLq57/Ic
7DI0dYWBCBKvHmS8HOcz/gqdcJWqIDKsX5+4SfExRKro7xsknIM2LjuHowMXz2Nq
C8ftHsARVDquJx/Ih+ERrqJD+KcbFKaeC7TNphiqD/TfxH2Iu7Kouf0Bz7T7Ivjn
5rA4+LK6Lo0LakGuipfPigusI7tXPheuc+MeLNKTKDgQHNs44djTwq0vQ5fmjRpY
wzntbIbSeImNeo6cIOXzvWtq0K9TK/YAuVXY6dxqwpGcq4BQL38Yc5QXy9ZwRm77
pNZQNBuksKZJBzfO/CNlVRnbgfGeUrpQ3oPuxg0JoJKAN01IViBoYcS5R9SbiCkY
pUswbnu/lJiU73FV7bnnJUfPRL+ui4J0Y+XNhvmTwDCmn0DqGrvDr2LoYXTHwj1U
ughIoPq+d5bv6/31lyYNc0AmjRreHKY1FeGsakxWKcWoCJhStoGkRk8Cu2wwPUne
vxWFbQSBuu70pM3fr4FXwvQxSwbyvL/L86CICW57viv9s6TqWZJbEGRIh+EZegso
OyI9QbQMCm/cgc1+1/LkaF4NaVnF+O2HUCYoPoQowjMK9G7rfH3fN6KwRfg4aXvw
2whbpBnCmQqKZ0T45h9XXmcxECrEucbJJMwwpQ1mYm5bJIze5V+Zd8VSJIRHugU3
+8rDIi69NsMVv0tV1KPpuq3xsszQO8MHZQHKf3JF0BszWoDS/ggccVIJuPQj3/rm
VbqS/F7qnpFeKPplFB049IrM4xdD10YguqBlD3w3HqBBnwtp+zZkgl9AggztVGxe
eheY7SCdGhakw+oNqJYwfvWCWCKZ45cCHiIR1N56JCMZ4tyZJFypAaXD9CGORpvy
NZ02NueO1tsEuEdtjkHUe2iZQtTYYCYMevfUE33S6p8JK5/8WQaMt3aC28WVEmO1
W85TqSIgU/eHF/RmQziY6B+CzC8rp2MXfYQN+gOxqmlFTn10l0Ey/j/9ir/tDvMU
GfpNKTXebLekHScdFMlKa4a00CFd3RBdfrR/tQFfGGjHBo9gOq76OPNA4BlgAImr
aAJNEK+n8PnelvbG7fc7n7LEgrJsuS055/h32jaZF31/ZmmaN8o/9RUcMu8Z6iGl
A3RvLUA57+FwNfm+nR+d/jbTH033K/EjjsHZoxphw/2Q7JkS8X3rUkO4zzCxqQXT
zAUFyzk6Ts/6/GZga1fbzC1e8q6ASBTa/8pGjmhScg5PZs2ARYCTFTPqZGz0WAJm
kgEeM3ZmEVhEfvFPVVO7xPbHwIqm/+hGLSxHqe9YI85uQKMMXkNcBHMAA1VSMSmn
//plghj0t6MsfU3QW0m6jnW0Mhv5J2IpxmDOZU/UWDPxoSQr+GmFOx2diqMwhUAk
PUuHJT5ADwBC3VNxG45h4U/K4WMn6EKFDzXtlmKJReUNhfmdPdsgaXpNt4nKXn8p
8LciV0s+YzwHgyt3hBWfJblndSr05rdgMN6pQpyUEndYaZhLAYQ5tWQdEBLN9tLb
NEzxyIJuVmKpHIaN66jwFLYFA/8acnjMINEuRw0oWFg9fk0lhHj5yPChP9g1zxWR
RXC/khCLyfrkQqmAgQqL833mGPVqEn+sfTkfCUeoFu2bocyGirgdBxcv6hhgESyC
BoDvuR68TFW0se5DZIX/pWkBOQ1mPlXtizMDWRO/eXlvJK/Y8+lCaktpCbmLP5/N
Tv3u2UZM9ZEPFAwf39nOfEBNILuoIHoaxwB66BHsqh50fC8bdvpa9Lc2VmkVqN0B
iqUE/PGDMCSGuv2smTP8rRUsK03LT/KKTYWV7p0YCaHDf9w8s31gFNzO0Ky15V9N
oVOgAhLmAJzC0IybztzwxhlCdwJi9zyUhW5QYSUEK4GZHdIdTyWs/z5htvzgmFMX
AUSivfiT/1bH+dib6GIIPwfV+Oousdk+8ORRydwBaOZWqXVUH3AN720ePy6TDy+G
Rvm697T9cbkqHCPra9Wn4mhfwd0PTuCmnqPmK1ybnTv7SOqenQbJ5Uvn2VJALkfU
eaQsMYD3WSLBTkmXPjeyVprPR17akRP65UvU7J2Af/8/kCQnnFyVlwWWjp4kl0wx
WCrnkuq6AVFJvgp9KldV9eg5IfJlQnPrbxqRpNYw4dvA0ajOt6orC3Bbk6bj6Z5J
f4tqviBEW9TJm6akzS7CmHwnx6RUtggnG55ubCiPn6bn6os9Kn1IxrAc/nw1qMLw
cZC/SLHmJatzT6znFcLz4WCYIa89NlxGvPUTpXS473VbPp781+CI9f7bwWhp35Dt
CDgl5YhwTDLYRsk8OcqJou1srDtN2gsUwuyoaTJXFzJvsQ8rlhaaZlo5p0J8BYci
Iv15jgs2RukeeM9wuVQj05HPInLiMtyicpEfT1UW8/7OHjaP+dILZptMWBt1N6Zb
78MCmGQHzVV7hNdC8i0qI9Xfw5Abki2zDHN290VsbhKtDeEfr2jPZPeNZi/+6t72
qszUA2OZkcfPYIPPTm1OqknstzGZUP1wnNL3fLe6FS2qXH54tjpDXvgn4pk2w6ay
8FLhQKM+YjCR6CJDcKSkI/JVg12zvW/oQ89sww7tUGeERffRvdDl5tbYPzqPB6Yn
ns/ch4y6u+K4+Y3ZxCfw35B/m1nhmubPmnkSIBis6nDHmEDXDVPzgn2veFN+vXuq
SXxpjvBPYgg0y3m3T2vxD0wPbQZuPoSdAvogVly90cWhZXTnbf4S+YWJ6rsXsmDB
2vXU27ziu4KI87yx45VzODOmNIjxP9ueczrZpYfO1+6Bg5hchbWFZldaS/QkTyU3
xlznVvuf8XTSbZjPDxcwE1PyWdZXrFjGiN1UiBsPb2jCg2PhFyqxCp33qldDCHV7
SJNN5s5wlaGcAqawS7X0sH5eqWFMw6bBseSR9cFWCLutNqJXUUFOZcTHRed785/v
ZHJWFvdMCys7PpAdlaXTAef3Ieq4waJY3YDYchVFq8UA/qnkrSZiVqyUJhm7DefV
cHI/jDEmArGdqHmv8oq3qPcn10TdhfqmAYX9sEoCOOw0AT3JOPkhMVKiuPU/Y+Lg
gSd7GeX+H4sXwnDOd6nGrJHViWK/0+mJlIoYE2QLwrnqqfGPDR3b5oNdWgKjeFbr
PBwfI2vyol9sAh48uKtSGog03/dS49Dc0I85SZtv/1kEJej5aA1qJhwiVnMBLMLI
r0/Paob5YFm8a1pvwr7ANyVUt3gWOp1JFGRAB2TOgd+lEl7ujVdyvZWym/h1TFRT
nNXRX0NIsnr6XzmnRc1Ljdrm0QoKu6/G/7hwFoVszh6jn/SxIhmiUZ0sbuodoQtU
YynQOJLTLX7U0CVq9D07bxwCpAp5/u/ThBg/KxlAvVri7GSsTEWKI9rjEC2xYXMq
1PpG8sz4y1K4zzfnXUNbVin95u6oHqvbFTjpyS8fnHUcNtaXp5gCEzDVtc1dPAuI
JS9iQJap+/Ud5tgR6P3GdbqEoiHWhdjz3CS3nYCJc3Hb2H/VreF1N7k/4E4kRtHR
OHG4Q/+1+QyedW8ADVlxtzYbKpLVoDKhTc8NB657L0WFcWiArEmpSj98K7zwSwd9
8ZF59W8eqGriSPg3IrUO25kqUI1WcWcb4xbfIKc2lMp+k2anZVbVc3yrQfmb3Mcd
fNCFW0kkEzDyU+Wf8HSUuia5CYWeR0sgcBsFkdRCdFw1sUgwDgHPQawcQWbzhvBx
l5eon7A2h3/tfbs8rfUZIdsWbKNO8AUXpXllI7H1S0t//9zI2L0JWpCli3aqExyo
tHzpSDqKIrKzNKCE2Jj1HJFBMG3tadXfuSVz9apE+Gr0UKt5RaYSKbYqqc49cyjJ
D6eDNanNMLXo+tzeUaxS5vM6peP9J826IUQe85iYcbGhBNLWqzjhEIcFwLuBx+BC
lFPjnHsNEN6k6hg63+lBxFAn7yHeE6Ouw2KaswmTGfzZksP7JuokInoESI8SW9az
kcXdJw579/nNgMKR1aJMCm0RMLLUFqarUjmSYrrMXLnTc36FUMAnkRqqlOrlysSJ
+uZBwobG3u1auAZCO8nXDxKnCzEQw/g69mzlMetGJhl/KvdcHSCJ5EPeiGVMr1ie
zMHz2cpYJOB/RIbH5aphk3VfqnteYkiKSh8vhr723OdHyaqb8sR6l7scnKWpufRn
X/c+EKjwX+oenl5Ac04on64WKW7PDiyd2Od4CEOWE2TX7eNzdwV9IKUXcYkCg3/Z
C1JTBR/h3eaiCOjhRrV3zOwFS9hPtN3brqxM0c+WiHLINEP76bCyj910sDFkGQrU
K0rEUpxDa3MCTW2GjMILXPLV8B6WPx/8d9qFRBGhsO/pm9m2PHxCcySlPi/d9q1/
TDi2/yWBaP9rBbRhyUjhf4x8JAQ4NhaOGYJD4fUOOj9SaW1puddaUJIIHGeLcYl3
QYwf+ABQRV4ILp5ehaiyuyt8sSyIzoSosRSHUixppfWQXdb/vXSfl9hKfGb6EBXa
lNCeyB/H9JKyZmTW061i8J3sc4Q7G2nnwBBYegOW/aE1pnacNwx7YKoPr1qgDkZU
p9R0jTg4SnPCOaXRs9Ls7BhD1BAae12Hk0SEFCiMr4/4J1tVaMJi3n/NrO3pKAC3
Ox/oYsVDQjL8isYIezdbVAxgADvinOImcEteNfXIjN2YU3kIF/krWGqSyp6FMX3R
omyTNo6bFuJbPDrStCKRporJyyu1awlK87CnecNECCXbODIqZ23y0/MjPFu5INXq
F5KnUUEv/6OHaNhl/b8nZwLlJ7tp1YHkayh3QtXnsUqfr9Jwp9QBgHY9kD2ptRoY
zz8w1HIJY1JEK4dY4qyhrOgjxRXYBo5jPPKhzxtcjcUooXBTly1a/2n6krg2DqYM
gJABQAGeL49hnz7KPo1HmRzcAlQi6/A3geVitcaDOrv3HCguq3PzQ2xPKtcRI8Wm
S3MIcrjhrUoyCIUphG4TswhvIO5xFM5sWx0FNN+anXANFPukdQCT9r0o1krVMZuz
VYVKXXsxW3kRNPngQCRup3GtDH0h7IlRWJ7L3wbqzLkV3moGtr9nTUu1yn1v7j7t
qtW88lj4HArHul6URTR4qcBg58CQcytWZkTXySbezlWHxP9p0l0XeUk05s5gjT6B
Wgyc5Hn8OGmsW5FEPiBcaBVGD6Zxuat2Sn8Q7uD6DnwB1FWwi933vg7MAn8j6FoN
O0CJf5oq523qRUIzWdAHa/PxjbDOJ4mHdaGZ1nY21vZzBV5wPbYW1eUqlwXywQNe
YQ98x33MpY0aIM0zI906biRugpuXe/vUhYt11Sy44QwFdXp9Tz3/CRZVu0WBaWmA
ywwVVKB7kivjO5hQBPycZHfHlu0PPuJmOzc8oexA7PnXBJ0lUN9uRi+PnOclvgf0
U1W8YrSYDnImFWyucIZhLDlzNE+HdJUeAKol7g8Wt2P0Gncdbx1FaXuWjVbT16R/
njfXcdjX0wth8YyDXxU3/dZJh/BT+yCi0Ouh9qtEOrVjkiHcXYZbksvcNfN65jMX
VNwOnSdE0wZaafFW+SzpZ3uX4ZshwPk+HcV76jqe9DUm69uRPczGFP9nlqERlLh/
CNOfmZ0f1116F26Me2GqHnNMvVUL10i3btb7uAnpHQEmvZA/36ro8+FkzaXvnObQ
l9k7pXcHIZHHRdqeWge7OvJ3m6xHun8TRfZA0vMuANWdxTI/v6u6sC52YGEPkA0j
Ud/FY2vf3DEFR7AtvHjX5iL12tMJi452s0bVbpUo3AQTefOodidM1hY/PMZ5xvYj
BjJG5AFmPrGTnZd4hBPA7QM+hGFH/uT/xtsY0SITjO6TFVQ4eCed5C307nxrSLq+
vGqLv9U90Ov+xWYbDHfr1KVNUJh0N1L7sMz7qq5FLph+4eOToFGmP9GD/Qqn7gZA
TffQlJNIuexxVUlUu6r5gfUtGQNRo+BbJ2uNZ1MF+gPCfRyiPY/YWNaUqEBiaAPw
uL6OQ/1ybZPENGchu+ToG7C5af90X7r44Mh+LPF10CoUt+GtoeyOlJGgJXP9DA11
f1Rpr1r1FJqI50nSjPqg5flSUcmKyFamRFlb3Vz28QTT2teNsp9hnCGJ0oEUNbdP
qHbPiA2BzRiN2mGuIT7FTYwOPRnk4Kil2VkvGRWcISbIm6zw3/kfgHeWVafr1j7+
kvTKXrKdKMbmYqiyNXozSyXSgWd7Oee49K0DTafX6to7kwbmj8sgTEcyiPOkN+E2
n0IsEtLNuEqKX2+S1mbL38Rx4cEwsoP+Cpj9pGcLHrW9w8cAggV2sFmuPc7FlzC5
NgPlJ5xf4vZodawSltkwNvjaFEI1GHygCAkUP+HrNqMFZgjwyEOm/EhEOqgbc9cz
bmxdX96N2rW9mr7zSjjl8ONE8dAJTjv3/mUXzl3ek6eto02/0bXVg8ajrB7neirc
T1x8v4+nHtQkpNdZLquBUhWBl+rwgUN9eM2VEza/W5g/EWiyiDL91yD8urVQo5Sw
ZeB/BNOgPy4WDa17ZiJW3lPkwlqD8gexWwqDSdX6dCTmYiOmKqP1qvXkAaBiqoZn
Ql5IOP00QT+K+MLUVWnPgrDG+9ZBUfVU15BLw+0EDnsx0Cp7tchYhkzXp00f5B/o
FBHGAu3D1cQ9fvdzNL2jJS0VKqHBZTgXFnjiXbssKffoIMLL+OuIEnRmKmcJhHJL
rYRhbyJbgTFdusRNWn6UDhQDvtVSMrZyjWkT22ymHBcn2Mswv6jimmbsuBZOLYEG
eYWUQ2jrZRxNO3fEbuYMkzkt0uGMsg2semSjlPe2koSDKpgK1QNQUXdjT/ci51xP
u8MRpNFqLuFRuZuaSG7CDqEfI7pC/zZRRAyNiCm720omuM+ACpPsxuq1VPLqg56/
upa8SAOmiN3Nfj53bKYYDZ5QrmSFsvj6PmW3E+gw1/J/WItWOPfLSkSjrzavthQB
v6gvk4ojJ0+qxteBp6zF2iPEtM9BwDSH1tC/ngE1RSztE25UCtVIPpQ9/W+OnQdA
1Vy0i2hbGoYkq0Ks09zEMMebweZjRFGXaGzJi04UZBHX8kNj9sqLX+8GvCAGs2IC
92lAaVr3OoRO54pt4tUUkBnVh6p85jFUptRglFByCv1khUbb9QJM+aAXHoG9vuNi
sYbHlWlSATkX5VzlZP8AySO4038L/uyvOpMvdlXVILTJ2dmr0AMv8K8nEhb8ZBBL
JYuhJJs7ZiCCVNWrvTI7d+DTtkNcb31281iEJ4vlgtq3P32PLTO54i4x3Q6MoB/+
dc+Xm9f6lwCmjoX4/hcYj7Zep5ynQor80OkAglna10KvyDPLlF3iUNajvekK/QBm
5NrmSkSw6I4I9wO6VaYceqmvbUfX+WyyA5LHng1QIAW6PK6eR6QWMaYfHeM7YlJM
GJj1I6QfDg6huY739aFJ9SH1bk2J4EBL5Xo7JMdNBb6OSTWShx3w/WbWut6/Pc4B
EM1Pa9+kK4XoLyzeHoXffCyq3aTkxkgColrHZwhWByZ9EX6sKW5OS1F5oPQj1zj3
xC29hR7A41Bi7M1SBd9aBlmOHKckaOoOAVCCufuF7znRYfkcwbSg1Su1kY5Wn6Ku
JtDE9IIkNPP+GIQDMyxaeY2ds2+BYJOPP8lP71D9X9pQ/xVUNfDVJXq7yP9GMXoP
+mjN/KOJTEXncfl4R8qswI3/Ol+mCwBGMNIj8qOlJR60J/DqoFgBWNQTH+7hiNEb
wD5Nbl7jCIryNiN7CV+5/99t3hPDU/RB+ZrwQ35gsbroFltZdHRnNmjx4fbcagDu
z3KZZrO6m9/9h64Ckyq67WRj4Wl//jJWdts1ceDwSv5tc59lg19gpN/IMGjVCTBi
9Qawlk8AejMcQ+QpD09LWY7rdNlbHH3NFwwiFRzPQl+yaIBZWWI6qCJS2/mILVUx
m7bafsKjTxoa91J71517IgLGtZAw1NMfuHpZ3Ovae2dSObS5vJrF9eOmQX6lQ2yT
QbQp45OT7gO29XqlYNnvDJXHKawWtsi1NIqJwxxAYqA/SMUS7l7J8bttPLzhG2n+
MjtpDqGYWHFPE7LKQBVm4XwY9bt9tWfB/sQgS3TwbTr5QpfwK+CsWy2Kvyhuu6sO
ABIthzAuMDoVdK8267rsZnJs9PH4imrRbOHXblq7Rz1PZ7NI2X056A2ay8lPDujP
w+1Hi09EQG8eMUgBeL5K7dCu4JXwVMu77Gelr+ilX1r+G4wxbyotx/3l9wuVoXGi
L9SuR5d/zPVdnBwLwWcCoTLrohNxznGdQKD+Lu+G5SYzmReXAb0YUPHw/ptqVq/J
/SdJ0o5QThFfCeB97GxnoGG9l4P1a33eilC1F4VetWIvCEB8UAqkes/DRmA8/55e
DPVVLEYgLNMn4/sB95OAsk8tu1/pchTOG/eoN0/UnyCQq+T5wxrOCKfvacqGWarh
+AnK0W5g7sfBqL7uwQF/T6zJdxbZKfysR0U35PSl+63BRQ6bO3od2LhUNcs2eq+g
WzZzQ+AUDMBYMM4eXl+hZsSxgscl+qXzwpoU0BzVhLvGuZ67uELBweI9JqgMf3uN
fsfD24DWXKlbDQohW7pi/VxorTynUse3E/IRIX29+gGeIO5uYxLLt4/4Xy3pk+jO
InoTE9RMjzEb9cg4JyBbsQKkWPVeJP4MPW7k7p+9BnZ7E2Y8mYUFombZElpii0XI
e7gHNcR795W5eNVezSFKZKU6l/mx+NaUAL24UtQYpMjn6gj5EXmQQgX8dNB74ki0
85iMiHJNzHnV9tkRCc1Ci2ROIfYMSGhNNp5TUuK1t7fC27GoqP+Bd0XQf/nxUut0
YJRaf/bSqCe7C9vvPumkfNrh84dKDIsh3vzkYP8YNLBnIr+RfK9Wg5h0Xg/uFnMp
O2a3+ftra69Ns6KJShGTjHr7j4HmTXGKJNEi6E3G4i7D1Bysuzj0U/3Mz48yGW4K
Su8/IF/a7tYNrLc2sIO3L7idHKIcp8Asw2BPZcHkkboU0djtVWbAspxI92ZeRU+a
pXz25FCkGyWysuiz8pNqE4BiU0c2T4u66OZZNsiwefv7IYPD0NuUGsGsF4yVLPQ+
zam2//Q6ink5zFAKnqmPi5sHmqDG8yYdRSl0Rlf9KyN9S8cmf155ZTLzwWvYAHmP
4aV7OOjj/NhLCk4mivNq3tXKKLhp9fTvilz2IeUOiJVBs38CdmNJ+BrMKruJTrH0
hm0vHafLMyOWSUjLlutIwgfXuzFe9RU8VIdmS/t4o5VmyrhRfL5bFh5OF2nWU4Fk
PuA3YgpfjuiASRAIQjqOCufadr7TcpYbQMt8BCAbcJ9CdDmmgms3ruhMRpuq1+ti
0o9Ha6pSPpwRaGehevZXHCUIa1JexY5KivbDAVoLO9VIO7Bih/vdbsRVg/dsD70O
T/LkMOlcF9C7AWLya0934UHtbKcm1GjbkfTsCqmuZFoZWdXPz2qek8+0tMSqOI7X
rfG2jBWQdnmbp+56V+7suYEqXXJUIQL1tbQdG35Qq6TVYlNyS2zK61VE7+lwctx8
wVAaga99cOYh8oY86bBrPkaamxgRj++trTmaOi2LvPZKufnz0yy6ltTFnJmFsDkX
298yqUooPItYU6AHm3WeAUOQPEIB4BK0QqribKszi2MsnT5s0rkuftU4CD4rJhYe
4b8m+AEHw6gxTKkt+JvvPyDD0ac1wZ81ZKCV9g6Sj5ajgyMRwI1sQIOu9d0bCgBs
qY6KPsT9qgPmz7+hvPPpXIq6A0GAxhCzHezzL8/i3KJPdWBb5lY8JvPGExsx9ppN
795eyB7VUZcminOxre9+8+rJAvGlYrisYxmt+mMfhX02zK566WbwQ/BifbmK26D0
tWT/IAXposeaYBfQhKSk9HP+3TvjVE87+rYx5RHk8nVPUazZpLdWQVW7r3LvVbJM
nUWQcQaCtwuDo9uHvvxq2S9ywQ+gWrffvjUYrmkv+Uxa8f127UjF6XrpgVRpb+aM
k3YMSrAXrbCSLNk7ZcvPaGkwY4DNiw+p0CcGZ9FVzZNPt1Ra/ZwMMLP2LC+rttGh
ybtwWsJZ3B2hz0jDgIvqXLllYtHPtUiwyj7gsfnQPzOEJTr0L01B0ZXhXosxI1qg
r6mVK7HYDWInUZZCb3jgfuuxWhobcxSttQBLWcjnRbnpK9ZKT8YRxx+M+aPRI2Z9
LG4Vm660jmci/w0MLJeIn5MrJMF/TMR+X60vbK6/4LYRcFlgw7ZLHqfnxqc2TTTh
SMbPhb309E4EoY73l3z3SEZxDL+MNJros9QPUfQYE6+1vvIwPZf5PZeQkNwStxsb
NKL6J67eXe7ePJHZsnhGUjQO8lYK7O2oR7Zp7NqcGOhWTmwWMVoUMEZIyPoxfieW
zMqFnhPFx5opoIw0Vf8IYqt1GMEy29A3iro33cwbcK48S6OZl7Jx0NVNWjnSrb1V
D5rdxpYslGeIIrgTQG4OhgpNw57Yre8o8VbgPRrkr0W39PRXcLWIJrmnWa7WpPDy
DSLJmtokJD65KPfVUneGpCsjVs5m32t6eJKVC/zybxCFmfwe2GNGZRVfLP95zX8a
fdaSl5IK1SSveLG/6E0S97wRVII0xz2cirIHeBiq4g+THKgwVd6eo7kLjDAXe9F4
vczdhU82ZzpFUuAVdqw8wa4ybdv1ChHKQowBIEx7tcu4HxMsorZl5nHPY0XZhSoh
s98kVHn61Ks3UGkYBgjbKQ9u+Os6+mxvUl3uKtq8D9n57sZpR+QHdb5qK1CyCCT7
Egea+IrzkvKqIcr1YDu0duWpVh9RwMCafmMZdWbtjtacemadIU3ax1ODjV31ILVG
8soSpZMJzdd0+9/c2/bSLwR7f1TXxDRMVABE9faatbDAkAkYg8oZ/9CbmhXgpLn1
iRK51u+Rl4dtssWGDoWlSk2lBYQ1xwajggnpsLZHO88e81TFaJCJSYYIGoaipGlV
LdXQa16SH3LC3PLHWb1y+/y8HTI5mzpAc93ZVpggNzQYtvtYCzmEiyFOKZDNUFba
EZqFq7gIsPbMiXSBnhc9nN9CGFu/taEIfBrsCCIZvhfa9auSBreh0rup5AfGaMLh
M4hxZc25y/TgdTO1ZnRsBOIevtfLiV4smc6GBc6541iGnWts+0oR+0Gsp8aZguje
zt5tpdYdSXW5zON3ypukl7WMp880Z+BUA4voAUx27jOd8vmeiTMvlrYTgbEbMUto
XICdXDK8uiSQeW8Bp4WNNWPJGMruNALlamECEpAH9eBZW5wo+tF3bcq3jt2LMS5S
mUzY09rlvl/LsPOx1FL9QY1rMrw+6BVO4U7YoSNGWqNxRiEnUZ3OqPgNvkQRnUBL
ENGpQUfvAUz/ZRNvycNXQdGJZwUP5OU2zyRV/rqOVXi1o5zkuJy0BJO3EvIfTiFh
jcm8dNb4Mwg46UyGMT+TGlXxPqTfLS6lvRSybOXIGGmewGoUBGXR9NJLj8o3q+kt
bTNUoGYjPRPM/fs1vFGQf4TPK5Cy6xSrayDu+SxckBzAmLyreW1Gh93NvnJ0mD1r
xvcOeJj9XMkapRII9bak9Yo54aUanXT2hBIPFtnPWhJZ8jV//Lwbovgx++eVTuVF
iCijClqWT8o6ZDf4G8oYvIM+fvoqoBhLtT/mXNdG0+VnQSmOVWaS/Rs8KaFmuUYy
IXBVlA9COpWBxG5o21whORrziLeACfU5kIgGm5FvCJ5p1Qo6jsvU1Lp3u7YP8B72
j2JanAAIJ6soKrR/5MVf2yr/aPdvqnZC0EVfG3X/cOS0Ib3h4FDm2AJkeElNzisa
6BQTztfej6PPesMxUfC+9nDU4PbX7BWeAWyxbDr2KXLvsG15Y5DsYJr34/0m3j1K
bbuywklpH1XULNCzXAUeb7D75A7LUBQpg+xfNlXTVgAgtApSyeSfUPdMH7PFokjn
VBpLv7YKaT2IC8Co2TarvpE9DMLZpC2BCEIZWCsTbSK6FIMTJ45K3tG4sdZN5rEZ
qohMJzntyVGoqDw3DJSiswqjx3pSubs26NoaOSGB5hejKemhlLC2Ovrw6wx7QSZz
CvtisRiR4neOvn9D5NS9m08dF/6nGgHssk/0EMSFMV5T8OHul4+O5X8RmYh9r7XU
mO/XWxM58UcxaN3FUL3MRFx9valjWsfDiHw05Zvmo3xl2EStDKpsib1mI/89LqHU
m1kK30aiDTf4mIlPNRDIJh/E8UWisaGXfvbpVQq0iQBIwrJjYvgOenIJXukotc0q
+zC+/PakNG63jUJH+w+Mu5d/9plvSCA96UB7oaQ71jYfM+TILlBQJp9LAThkICMZ
+yu90EFwjlVwGVRkve9O+p+PpIkzLhVY7JCf8JrDQ5hKMCsD8bit5P9agcpIVy+K
NwpPdjuNha6MYIUjdn4hwbCSrzyxWTQKvyUgGx/0dCSJ2/GKDRmELJk1yTIPQjXj
1eXSeIx1aUFBYFBk/j4VBCbadvrcKDF4RTklPn9/KGcmpxsm8TdUPCQbbWz5c+LI
GYCmMPM1cVMtT/spuCO44oBCU5Xa1XKx8uZi67zpI16GGEacM2bPdxsC5ojMGv75
SvEDPj3mffz77CWN0ENN6jf3ZUd/XhBoR2TG47H1+4pPL8EQgbHowMoDW0mhfkar
CtfEfIshPVW+TN5Bz3V9sgw7rJairBIwrDzM7ikxfavtJT3QtN7LWoV8/jLawknH
+IL6kpgm9cQpofUBwS3duG9WnZ+HlQcojqsyUneNgVDTEYzBw2HPpXZzuYHrLox6
lNzG3cOq0Zjtl2nrw/3oe2aJSiKg1wkXCP0yBApSu23NL5xLDh9P6NmPKcRmZ6Gc
+a83ACgoKU+ytgTTTb56nzkArSzlj1fy4n/Z6K3w+itOXzROCyW/nnKpxefyuwUa
jKCtC2/SrPvDgQVQBiaobfVH4jmIn6Zr6wDQGKqhfdeSLTAvWg4zPNOaPm+P3lnx
uQqQYDScmf7BiVWhjs1FjrS0/Cfigkii9gCIa7XeZsRafXYHCEFWBNkIKoh6zBL4
FhnaPgB0p5VllcY+y/Xv40qmJr6EnIuE8in8HerPG9YDjzYtkMFbn/3Gp5oj0UEC
DDaHFAS0SS687POg5kRs03dnJqz6lX5PhyusUSzva/tJcej+wjc6fpRRHofyHA6u
5N4z7f8z5RQkCeEEwQhZvWAyfOjwZxjEIq/gjDtY3/mBxNpbLpZ/SSSIZsySQWDI
JnU+ALAB5Mc5K3Xl1VvwT80Qj//kDp9VMpmyiR3c6PWcZC8GKEJQ7gmabKdvh5gC
6UtxwSDh57mPRrGlihihuqVMpgBCkhzADmvLnNjbV1f33b5KJEDlReZnaE6ntFuy
azvtSoDCOn/9WLoqC9vS4Bu6cIusFN3ob4lR0ZEe/eg220JThH/M9FXTFO1qbxAG
s7jdKOep5aEH1jbsQRzCYyudQ7OvQL/5ErI3opiIZOyf+vxHazbm66z2N2ppJk67
77SSGrRzPRXna6U2n/4xvxYQakd/2b6B0r3c8+tWriL2f7BagHEPcNcC0T6VMywo
W4nuVNOyv4ZpwBG9FcR6yQOGhSPhpXXlkVBzaZ2AR7TRrSBMGFp+OpViij6nmJfK
Uw3VibcYdyWGWSEbskurn1RkjrBnRsS8iXtGh+W7dPG4nb5jH+uDuQoBYIdxH57a
lnGvrI/z2DVIb6F6e6n8bFm0pKIhqmMpoOQlTCkHruxLtnRs7M7BYJSAxEB9Vluf
BKkqkw/rDFcWl1/2QoKvsN4hB4rLy4tTYZtc9VjB+UPVKjt2PN1JF9Tws3JKi6vl
klrLIs74+iMzmvA9ndfoafD6XJtTPhnizwLWaTYYiMctxynC6uiw8ncsPbE7X9gP
bovR+Ho03E5R2IFpxi4J9ZrbrWSbW+VxKREWf3Z757oCf1rRuMD4RZwTXA22oTeF
xix0gZZohoruzxxI9KFse6m6hwytc2ZmIVG6l+LYGofjt/tQnHxmFMRCAVG5SYmw
vvEERecFfI1maBHUYl7IYGP/qR6Bxl74fAhVIM4s2+tBIti2OdhhFflirZd/TPJ7
9EYcljC1VDC9wQoZXIL1X7c7eiyjK/bAuIDSlQlhwB0T/edtU5rOs2ygDAf/+ZRN
AEYbcsun+TssH4u/Q6xt81J0Y2ZhOJHZqVIKAYHffA3mGk0aTbVFoTO1uBUiAXJi
shxZ/SAXBdTmgcuhQAMexISbAg7s7aNeFslaJk1nZo3z+TYwRkOtpQ76aLxr4qnZ
SKezCJMDI7Dkw87LwJg6fgkf4cMBWmIkAEa/6DUFea1IKeMwUBPs3POyAH0a1kK3
+MFUExz+DhGE9AvCZ9uG2wR8IaQxmf+OYm6qAbf+EPmk6/JYvVbiAIW7drbzGjVz
qZ1DGZPuvpDyljvpbnwyfA37JnSTe42HQmmdeSFGUZ++gA59mGHh259ChnOulrgw
qCPG8vtXp7haQGYQHIoMHVo1EzIWQ8UbzcH7S9amN3px5xaNY5vuhnfD6PXOjrkz
3pD+P2+o/sq950IYCxELZKLr4O392HrOQii2ij9i04yGBGrCDp0FRRsWhwwI789T
3A81FBMkA7WSBdhJ2KLTfObSOgigHdKRlzPFIBUc/llIIrrs6fOQpM4fr3JaZ1rB
QFnQYD+16cV8qaMyEv6OriKTkuluQ9tQVz1o3t4iJPfUykoSShMEhRm5KMp8gsTo
SOsv8V5rGeqGXStrf+N+R+SOohksETP1Wnlb+mLSaqDi1Wo7UzvyO6ksfM4qlncJ
z2QLz9FtLlEnQhxpNUxRQ01TQRXH7z4KIVp8iGrvPl0Ey2fMqK6E12mjtk/cYZAk
EL1WFa2u2ernj+R4udo4JFBlujV4pF+cQ54+wPUv9bIM60uezLit3YkOS7kdYBdz
rGX6zMJ05vsQ3cr/MDSbPjnfpjfePkt2Xrbda5l8KFY6gu8qeE45J2J147gXOT3B
DhUJrnA3pfxj9BojBaqjjKpzFjNQPSfz6sDtBjmLV27cd0Bi/QhbLPRkEIP/IgsM
FD3fEBkUYH7fJzWkfXu91IRJQH/TPo13eC4ZPpgP7lSLHzNjety915Nu/7+giRwl
9m5kNcBTpY/QJjZoT6UQizsI8Spf16HZ83XgRMI2unv9c76hW7CK9K7gIeO98gz/
qKBv8E03RiXidsi2/MYy2QVmGFovqkjYKeQ2v4OAmKxrcmva32GCIe/vJgZqC5U7
DLn7LGIttBdFgrbbzX9EW62DndhkX982K5u6ZMcSUtcLBc3IiaCkVE3ONl6/pURD
43Y6IBe6n+tSGzHrfloUsGiq5svCDeKciiinH2DJY9okvmw9Qrb6PImVhC4V8Ds9
Xcd51yUYBeq6ZUQLSyCMbbujQYMrV7hb83Ynvu3s2ymfkcC5XLUuD01QQ6Az9rwQ
0MEIxxjSV6DiKnX5jwpp9oLs7Nyr5S2WzRLccon3J2eCFdRT/JGFneg7Z8uUIKz4
ZG/X82Lq+ulIKAxznNueME/IWHR0WTyQi0Bxilps0/WLcdMDkKrM3x8/uX0YuWsf
PUDzc2wWcOWTK/xxb0+IGnPM1HRm2ZYPj4yV/ikcCTn2KTm0au0CcCoaYFpLeRFO
sMWcXUglsktNioNfU9PYMn7TsD1iU3t6bBZP6OCJxRweCoAr8ehV2YliBWhKcvXf
e3jsWWIboaBw29PU2Zkj6RWDWBPwWQnN+Pst6QbcUHVum8Wll//lV1meglJ4U6Ny
lLoLe+2xsxh+cLTPJLQIOjpssr7ZO/abGaaTl1Gz7ROyiRNDXUVWNSNtPOdcVe2O
bIf3x2beooX6pwzbzbiRZMPGn6rV3QKSEjamAbR2/IbXNDrviOYXs7c65HWgiqXv
rE8IcltXptfxFeWn2oiOmg7w1fhLwraawCw6XbgkgZmwDpEPGWMsrdIro4Ryr+qj
0j2mBSVAtMSlacldwacJfGQ12jAjavSowfaxIA2enj8x0jXcNaRXRF45n59SF8y8
XEJ3GnpOI2+CJuVzxiody554E0XcxkOiWw11wYW02A8gohdm3kIv5EFwkyfcrUnN
37KmsBrGT1ojs1C7sIHikHh+1eByUOUcbVCHBD8S9qIJt4bfn2Kgams/RP0sevz/
P7QR4F23QKs1+oFqs/cB02sL8dOYLaJ0l1dlLpCFObBBa9xYQHM5pbrIj8tt+ESF
XSSInUqHsBGlPmyhjcyWQrNlBuz33redLR0fH/aUoR4y9W3Tjv7bONVxMamJdMXE
X6STkYGCvxzwQr3YfHvv3VU+VHgaKv99P/3aZP1xxc4iXSODedZ5hMVfSYqRoMFJ
gg1SWjf3NH3Scwv0KecmxTlb9BuDSpX+xAP0ZkKCbpjZGETzj7/8ex2rLhuECj/Z
FXUrnoDAtj2aGtHh3IF7+szw1uvCX/kjMoQV1WK6F6q5c3G4Io7KuqoxsV+STGVc
1a/zDm0YwOmgVSnoVWY+/9A7INVJ4SBflNLZONdrEzuybtughFmrr933r98AzPJf
fPL4gFDLmh0EBy2r6hv9ixtgGjiikugf3AnccsgRcCUs1LMUs6J32vtUizQOy/SF
2EZAWt6q0/Qh67KZ0YNwc5vYwemxOLE0czS+IzXfG0J783ZYDGYi1ZUhYlB3rfl9
Ug0gq71ZMfMDx3Ks6Ht7lmXK/pHZqr5EQdA1kA3YuFFyp2DIBWvK9iTUJB6WVuIo
tt8Dm5MnadcGK+ihSpqSeOFDzaBFpPGUJqhsbs3r5WZFfrCplEDaBnZbR/1kZqwR
sD28MncRHYGGpZHju073CsukhNtCvHeCq7YSj9rVr1yGdnF1JcOXjTA1VXlpLs1z
WT4jsnntcEvspeqyfLkzlff3uPJG0DJv8Tisar2mb4uYfwbGPOUFGPMg9qdy12+Y
x0+Y81Sp3HKPxsV7oSYLkoK2WXXKBPBDoB5Y0POHj1s1vNvv3rHNdUFCnsd9brTr
r/bnllPmGn8shdxtHsWzbDiH8mulcJHtCLwejnUpSa496Sf1Efw3LzCT2PSFkX6L
nNHfOb0cxA9/+rfYife1J06zqxTsM1RVVvsinRuh8RXQJg18+PBRXdL2Zmkse1eR
Z0/BpO3EMafK0PukX7gMjpwNyHxPtoAr8/rzvmgJaMi0PcY8P1yP9aSvvC2nXaly
1IgR3wT7ua/VYHerco/3gKhhNIRjRZjg3RGOu05DKuhMZ/DZZCEXQy+GLzqyOSpV
Uz1/HekyK8wsn8hCdKxwf9zjBmZbjEv4SViUPOb8b9SYZfTWwz+5OPIqqY8db7tP
sl6mLyVgGel2XJ4gmTivtPjs0ODRqGXN7RWQoGj224jSJGwBFAlhc3Fb6VYlQxVO
Vojj6V+JJiNhPS77SBslUEMK4z8IdMhKw6YUr9RKvMb7n4bN0kejJpFJYWiLCv82
DdA2qeAOXr0pxe9An2cRRIV6nVoHdP/JF7w24ioA9SAnBtAJ/SF2dRN+dRzhmqsA
uHb57CDrjS61bxKanGodnONSIjslaA4x1rJ/8pSjuuGAFA57aWPzggmcu1KlOnvh
XfTFg/E80vuzFuWtIJ2oqOq6Ls9N2TjziQetRbzqP1Or3kxJH38sU+sp/YyVE7Ud
K1fQwKdZI1LcemtWSvDRULe5HzBkfiOI6N9Y0bd1kMlNupnSgt4j3eCvZ69bj9vV
oQCRdZMr1CzbtSgc/MOFZInkQ/Pvx8PttZkqxzzpY34twHT89Ll0njYxpEi45ujI
4Xurm1FxXXlK7We8AeBtQunEDJnRb81Axhr4DBhincl4HWdFt1OBSmmrmxtdYh0x
cgEOSd6aZcopqOkYp+ut2hb8gs3kzXq8Ra8Jt55dYAZe1NB9+9j9xUIgYzEYYCZN
9NI2sHo8o++5c69BOn14ruzOxj3/aT8u3IRDrRvZ03uftbYf7PBpiHgZ8cS/ePin
fV5a810WeFKu9MwhNmlN4mQMIJD5wqJ4K5jRe2XMeGg/3n9AtvqzTeH2zajZpYdb
kcs90ETQ9srOfQLQgXZs4KQCZHF+wzLdqIaLYl1WjDhxn3BgJMW1uoR0aon8GbZy
dz9IMWD/tIaMud1IytSrFo+SXXeICFUaZEpnk7SHm9BRzfJ8ZkO8YRGXP0WKMKj8
jc7AivtgPL8kxScu/CxGImzM4Jx0vFu0CYMCHwziE80JqgYaXWyv5DifMZlzZ5/U
IHzfFfs2Byo7z7zTsqVixHkw4mLmsmwV8YgGHBOnZKGw6qW/4L9CBuddSNCHNXQH
7ZmCDakif0M8MiyjfQWHHKIYYz/l094Wb9nPVVrv9czm9l6Fhw6bk9iyoAuTwYDv
6fOivK+uw2668slg78V6PvXd/SUdg+EM+CsmOEMZWvizfQx1h8OG4qS/QDEwl6Bw
EgReHaWI5okJ6C1ixQJbIGOwOo21zJ1XsgWEHsuYKN6xL6oiSTK1oeBKx8dycJEh
FWA4RGVFRXXkQ9CP2iERWz+w0BcgJ3MBFKl16rIwH8h0ZHa/gj2txqKypXiTE57X
fkUGmzz+gAxHFCMEjP/9MSSwHUwyjtBiOhANg8RFs02KzWqkM6GVBfFYkfpHSFta
eBPwY7G24ny5a3QyqwEJkuEPQGyfhgIzmPvE/vIBALza8V4z5PyH43DldlL7GUjS
lQ/p4OjJ3RvWpLYoz+e2jy2A6USXTcSS77TJXnMP+8XMWRxsiZekVVDszp92S7j+
4fEiYSYFELBqdKxMYZjGcm9G0IdaCE7uCA1L9D/3R+YoLn5U9NwWyHD+/sGpR0Zf
sTLavW3RQGff43Bxm6FE9qtFTQ8vcANYrMOjHeytZYac0KrHpAz6abLGsPDjlFIB
ZxuOkVf/DFT9jYBm2OlYUKxQt7ryyPky2xf7GYanPQZep672N4DHy67trvT4/Srb
FKl8NuYZJSGWAWWbTa7hg5PcO6+FAirDrtK6tyKc0jzZl0tsVrFEAn+Qqfl3J91U
SB6RBfSKNwt+RQg0q0aSwYeOT7U40IS8WRusKcxUX47Si5jDYORvvAlxyAzh+e0M
SJy8JXbY+hByKEpUfX8MLKleTLZs4ADCSF4bmWarrWIbviPitVKLwNKshpAxDlVL
BU0Mm5rK5MxcOuCG1kYVx9wtAJT1VQfEckn0ysYMj0lVm5sWcOc9xHEd2nc9ufgK
uJC84xlJS3qsW/lcBq2MqC+4HydqzhtnVYR0ebXt0+Qff+b0913olwiDePiBWh1W
Y4Nh/vnkRM5pMpT84Hc5v4UP5ulXxM9GG/ZAY6dl05NdsfelnopsdbMF70sA6Had
iULCUks8U9w35FeXonTMBohUIufqkf4k43tg89IfZZ0jYTlzSFDtvDoZJlN4HgDd
bJEusm2+JTeT6CxpakNr83w3uXGJ0BQ0Th0EHxQOmq2lJTrFc8w1cXeSReizUnwr
XtNNElQ3MSShvbe7mRCdDbtq2G1Ki2nSpyb2NGOHef4nvETz0dFAoX4qOQzuupQy
AqlGxOOOWyqqXCrPLVKpVWLv0TfgL1RbKg7tqkIC/eENVnSbKjyg7GOyzdLRDJpZ
SY7gkhUUdUUlwS1GS9xSGmVEtqxd0N/zJX8kN11pAMHfaB+8LHNDPTxYHQL1rvgn
azRmAbagfb9IGcT+/moDomRhq+6/laeoD+DUqhc0Q3lMOlmxGVpgIrbF8gPxQj5S
yBDS0ZVN1FutqqFEsyeIzmEeEJPczkw6P56X87Qn4EgGnMC8D6ExVyq7L5ml3Fju
yGA8gc2dqE3PD3/VnuAVpWEUYc8Q+HxEc8iDH5qdBAb0+FjCNF9786/RVJUIMBPt
uf6vjNiZarZVVR6pHXq4OK898mCIkP7AYuUeabvzLgDjuStiDp49s152TaFuV5AE
6gusH9kq+8DH+v8gSCV30h/s/LkWZ1+3xhF43UmfXdDJY/d9H3cf2A2mYS/s8U3J
E+FuCo2Uo1+scHrPWp8k3+1s2R8xH1vKSdO5nzs+dg9lC7KQyaFw6PSZ7mnPfpjD
MduHDetpYMAB+QP197fLXPR5pu60UVOU/kgXeub+trsGHRbp7hlUciJYVjjgP2d5
ZtJw2GmAl/kfpnjeImSwNZiBI7AzKFQvdtZBxm/BmnEvpD5NlKW4qj5xg1uJDBlE
Wu23zNFZ/KdCJyX0vU+oWyl4mb840AcwNyFAeZH6s92Jm51odQuoWSzHp3OXZBUA
9GRcuzATsCzRYZT8lcxRtd9HgJ43wpHEl3HYBxGhZURxnotbS8DaBPEli15fTXEA
MolMW1Z4TZrm6n+pwQAoowLcFTSS3uh9ZaHz1l3HtxTNwIrjl4NU4dt0OvOYEfJz
Ftzoo2UMwHyK1ynSSYZI92lIkDf3LE3s2WpGcZdjMcZPpeKeA5zMV8yZMTpjVX+D
x4+1fmpdXX2yPMVi2XgdP+iHstBeUc489kruEoRwgvQmbL2Mrym2fMWokH8W5Iu4
MDrwyWVSuaOihrFnmcvehDlKDx7SNoTQ/csdz+q/y4yCBdTFE8mFByRgpDZH7jug
32IKRjDraIaoF/Oc5JAj/P6ojOpM61lQlEbwii6HszbwOVP+sNhm9fr7a3uNLlj+
+/DDx4mKuqDZqmyaDuKeXB65ee0iXmQCXyHCiqh1HB6gAMg6YzosWZseZdTz1LPy
hlca6/hamSTPHxdPsK3ggQmds2nwnxA8crcpYK8OF2FOT2SDLON7Mn8VFTFNPkUQ
Nr1+pVnx36w2UoZlXUeSbMRny57Hm00avp89z/IJfAJ+GIfQxumC4QT1+EXiBTHt
zO5zxoCPDX9MxQcV2uVZDX7RteN1Lw8LVuJ9DcRieyCCkhlFjvvLUfQu5Ul5Y4UL
5o7zulbHcUTu5JaMThXtZxwQd0NE4dO2tTITNdZlc8z5GMIYBS5bbQrnHd9TZPso
ZbcFv2fjssAJ9Py27DI2uHu9Z9bSoY+GwFBFvkrg9HSXdnCUlYOssxJCO39l5VIm
a9UBE1vaRpEuiiZJG0ZHvMo1aQpkLt6QaCdtPEdur9iC1QMmHaRbK1GBEs/Echb1
ujyN1VTNrKriRiimBl7bsoxM+xwHbHLfoZQTQ+nAksC1ftLcfNfZdQdVFebZZ+no
9XXd1tv5csqvy5M6ait0v/blpSo7OfMtCbA61380zuMCW5QcyIOhNqfTnJOKzo1R
yyYWCMr5VO588Q432Gj4L0PhROt7YxkzGzNjjfjiQI+WDiaZBXYtPqx4FCsP7pQY
3rhkY+hgmILuOvjVeKFeKsib7n2SbMqjxBKD9x2b4D/k/whAeQEbTfvzoWQ3Bm78
8saGJxXeSCVIaZn9p5zuuzpBJz5izqOyD+P84tChSSXcF9DwtP1anMbEGBCWnvAE
eVHnX423HtyDo6f1toRb8Ja3N14M9stNYz06A/MsiUt+9egF3LpWT8kiG83JZvrm
uzW55dUhyYCv2qH/m/KgH9l35udz6Ma0gBfOL43cgJTfwV6MM9L4fje2S7PCqYMC
Igwe8PUZOs4Ra+qviRz+5tUw/5C+/EVe5QKhYwmpW6DbOIEH3da8dTNGrLQ9qAjy
qHLT/x87UP8kW5hzp8Wp+F0WwAPM6Y++CvfieKi9/24Dld4weqh3MTfHSIvoZv+q
WRwVVhOmVb1gjCEaFkn22M43ilqnEthQlNwpmFR3bw9rUcI2LhV2oCIkfrtxo1eN
tcTqx6Xak4bNELiGoZB3rtXdiT0BTqK+I6cnwDsPfcxdfkUYL0Qh5b2nJqH8ViFl
rxnCueerXQMTfaEY13tIbdP2kB2ycGymGY6Knek6OUsWqjmlRjwrK1roqhOtm9i2
mZudQD/o3BjHlziwSqI92wzOil4zcuo4SnX+MV5wjP69NrZXijGwGi2byMDQHgoj
zQTc7nAZZQXOzkvQ83PEh2QLGhGfFNjBslPUDHc6ktsK/g2fua1kFlbxZCXKR/VC
2ko+mP6jyK1TLISMfAWW4Wt283tFuvdG4uGNcaUIjlcG5U01TM1uKR0BIs4BEj8M
E2HFLbTTBndDD2oSZKyXfjQ7E0O4z7Zr9u1jalIXOSlRMx8mpy0KAd/lAKUurztO
/35aAYt5n/Y+HaxOvAN8N4V6l1pr+hOMZnKge3bRqCqyKJn1/Esaw6vGvVyJ3Vfg
QrZhlWfNqlexWjFdRnojdLyn9alg7r8fUh/HIbpsIRB2IZeCYZswC1nuPo3OJ3GQ
Gnpo83D4SB6c6cJJtJvzHyAd9Tr4TOrvcZpU0qf3rhMh2oEonoBTzfnTtXFrxQub
PO2PESHK2acIvz3SdUCZrQjuU1o5Wk+67NFoqtgLtpwat0Q06AcafnDr+VVPnChc
S3KvHc9NepVfJWhLDUGESB7Vg7aPIrp0D9cMPoDqYXAqzpziJozJzqP9SftDF1sV
ahHPu3+37mgrPWazeHxhHzLy8kSZqALxD+C0/3lQ/0mlGJQ7ixtwM6XkmnsCfe96
mRd8C8t9I1eAjNgeqMb2oq4vNiIHii6d+MHWLh3u/GaUNn+inQaoWvPrQuImtuLA
capmkoysKIM1ctSx0PF+R8Niwr4zp4Ykmxi4QRqZ+w63w3wbABsQnuZsfpa48TFN
vaYbYFbAyZxe9zB+tRz0YMRGuIeTPRjdJkd+JoprFg0G6J/uYw85jaK+DRj+urbj
EY/ucp7uNRTbALF+74D5DWEaMUr3hCuifXxcXz/BHkUDUAM0ihbtLrXpssiWGx+y
H3p34Zv6Bvw7Se+nzmbyrNQsUBttmCGLQdlEjR/BlvhbuQsjl8LlBkhaM+qw0JPW
VLkx3zIAgfd1ZhkAr6t+81YK/de8G8Zmz98+fm0nsgHjxKgPhdC1VuTvt3uZA0GB
0we2th8gWG353uQa/+0M6h3BYCO9gXyC2yuTgKyAM5jJDmL4GnNrJNeMwfHxZb/D
hPtmv4Vmh73aV0NWrtNzipRl6iKQTJjmiwybxgvmnja9/9PRmtdtZ/F97vOLmQqr
K2r+0uxRFZb6Owbw17x7/naM4iF5WFkR3+1M7ocBDp2eOVNv6QFq5L4M/rBx+jOh
j+re8wPblBcpcM0Rr3FrBZEvUEhMNzflCkJGFBozn4BY6lOHp2GBXuj7bFCe7BsP
8XI3+ngWFSmh1+V7zdZUzAKdzffdO0Yigdl8F7/McL156yfqqIHUa6oszEAh228V
yDDLnN5xd5PKSvsjkahrkY+nSoVRp5UKSuSzY78/imbtexCyV4Dx7qlAiw/vJQ2u
oqQTAi2USdDMODPZESQlozfGEs7qPmyH77fjRZUQ9LXkUa8W53kxpQTaWzf5pIP4
Uf5dkya37GQe6iriRXTRD0f8BPHRjSrrmkb5tqZSU9eF4aQVKA7OANdVenRCbXwZ
qtOegCZnguR/TDnwZWz1AnTdSaAYSnoGHyIDyIEzMoEcfMNae5z2SbbgZrKQaqnW
1Ib46Jio3Dk6d4aLWLNsUspJip/mK3cWMC+2rWuewzPl8xn4SRCXaKoxAQIuZxQS
xxXRVUI6NdVV51WeWc86m12SIFjkjIIV+zhD7JC7+BsEuXiLIeq9VAFQewtG1eo0
1OX7L12ScQ8vXsumCVrYvXwlYNsK6GLONfy7MTuM/ti8dMpds8/ZhUN6SnmgkHU+
yGtaThQzcoqlzvTYkQenyP8IhM+JiL7PhTxZ+PFUTwP9QfegtJJ+7hL0tjzKiS1T
wGWTLp6/iIoJC3rRzENA/GfUEHBHaLieoT7891UvObDVAArbiOzWJT9IDHKXv8WX
2BwuZJflWLOCSZWd2P1r09zeSYaLEd/VQUoKCv18TF4Q5tjXHAW8OjW7HfOi3GZ8
XrWZKqxcFK65rsgixpIj7jFHA1tnBItiTpbd1YY/kFlnbpadNNZgK5rBqCSySzfR
AJeJm6tlXYPeha1va4AUYHQthsYo/UkERzPZPnm5Mn0baub+9uwXWlmuV4CnjXf+
kjAZ6cmFXH2Nr8tDdlCd5K3b56cHT0fbvLPQmFj0O8gJVZKqsZGc0GxMbU2knXU+
s5SpVzNHkWHXnk/lZTLhFc/nPfyxqmAs+bErbbomzbxM48hHHJVZs1iwrOwnMNb0
9n2+D+KRdDMNqF/c45wPJ2dXWhsxvGm7hI3ngCxMGnZ+IX6cKeGsYdLq3C4rqI1a
hup/+jiISiZTjVw1lHaEl/DJZN9UEycrI7bC6/SeS2Qq7S2aSGkcswHgp73OOZrO
qt0TEhslHjV2NWDoxynX59suLw/pw4LhTHWUFaYoGnd5I4pI8bS32MdMB6XQOjW8
AknhV1v7Wf9mVm2CGpm5AuihatxnLUBKzTDDNUKjEMFGt4Nnx3Cxgk2nsGs/VpPm
PLA/ZjWLwr8kSrTbK0kCdw851bQWyHEJQUkxYZkTS7iI/aTSKjeXx+Z9i/3Byv3A
tPV7jEGJrqfmV9dwn1ksI95Iji1yz4QgDHwnVYIGlDI9hBwmh4VVipmdtu7vgVf1
Xyap3d0xbV6AYbPqX3fdwAjQgPpOxfCWQug3GPFT56XtBCD6/oq2CR1F4itV5b5y
PG79yjJaOnV+JreCi+hoHTXgmg2J8oxL97UQxFTm3rPnlnOLNSbH8Ot6MOLMvFM2
HhoLWW4tVv2dmII1Vm1p2af12C/v8CwE0/be9AUubh2U1aiP9Nib5YYyP6cIWt/l
2D49WMECHUZvFqUxDqj+rrQKUWmFRflpVdPmBrXMGqWUqC2j/Zg6Y8VoBjr8AAtn
+qBXg4HRyVOWmxYGSkw9IK/o7xs9gH7SBp7GokCT4IvLgmYU2oxGMi5RZPmPCOWl
AQKbJubf7nYJNEXuzBiGPia4LFHVJtxLghIlV4rQ32sMjJed9paqZfQI9VR+8r2Q
H0z2DBSXr3aDZ81hLa/yrJt8Jmy++hVGK5k7s6FZd+5IUFbEdZCiWpUIC+vsTGxw
G2AlvjsjWA07reBzUGUVQmnFcTSQY/iLLtX8uWzsn5sCsZu8ZzvxxQYyULx4/yXg
fQQL4hc4RngbfkWSKxdtx3ypBV65UOPZxAseXQtq/gANE3WDMFRgkaKXp9F15pB/
sy9LEgj1XAws4oL2Lu14TeCMzdIYOn0MWjUD3jh3amKw0/CWT3oOL+5Bt0F/+NyG
W+3gc/0R+opE7mDgQInsxuxNfSA0rYAGIcZhNh7IDxco+iN63bRZbXrY8eObaYzp
TmRE61i7oYhhIR0cLCmb1fKYrngEBsDGyfB3pG3ioXXU0MrEIeS+u/8o+SmSnwJ7
+kaCosz7TRra1HJ2IpudaRBVOLoEfTZhiHzy4zovuu03BCmxVQKt8tsyAFbABMT2
LiCxpKBo9GHpOgJdCz4ZUdutQYol8UEb4pjJKsrHAIFwHe1ybpvrNZVUTUi9sgK9
z3n+df8zN9lSsmxWhobfBipFZKVjGRtNaW5grYvCBLxzeUzAk2L+zqj68y4Nmpv3
rXpeuoFzYIpL8FlT4dUOIH4mu3//0g9GKd51+BpGnEPF2C8VS30AAMYpTxY0oY2l
QDjMiVY2AZhe/ONFJI68cPsmdDTRy0xSorNd9p+PHwmeUBQc1bWI2SABiaD3dtku
fW+ZN7h3sb5fFFpcbRlClb0jhwYg+R3WIQjtEY7cM5yYJIvoTXrYic79RqbLJw2j
ZYEEmk9amReo9cHrAdRHLIFMZrjp+0B8BAEEpGpVlf81w36G/38Yc9+iXRFsjcUn
969XDloKIdbxinTossl8lFxurTd+bbAu7+lZyB5YyiyK90sIGMnMtfPunQtPGxi/
iGhAmMPkgzsnUQ8LzkONDLkoONATxnFqoyT/KJX+acwno8wqQmAVtWZxzE4niZq1
Zkz7IgkbR7jMXcNCWtGGzv90iyG5ePAt54x/uIXwu7JVE/vetclh5GmUhBv0QJi6
0qdMPSkA//xCfd2oHQyJW9CAhY330zCKelizOXyL+wW9uMxevJhxJBNxyfzNks56
m9hg9fhtdgGlge4c1HYV+Y0hBdQInTr0iVWBzg+o1EYyrej/vaPUN1n2lGGiKohN
xbM5vaDM0VwNawu2c/x7TyshyA/8NbZKbDHNrBWt00q8OWUHnuRc0rvSZiviYlaI
PIosuaLbdPwlAxk25TywE6Ztump5I2Sgy5vuRRzWTM393wEJnYIubFsfvosvKhv+
8/Ms4fYgT85mzf8SD+9jz0MnwpfdziqGXqnvQt7SLJ70Dho7QPvfMP7RZckniI4V
Tnf3fBJNAP1m9xwuefwJ/0rI70vaayq16P+Hkkz2H5io4CyTHd7cib/DTx8Bc1Oi
XDric6Dk42LBAbvW9KKKi1eaPFzmjaMrV4W5OMuQTyPAnDwVWNoGrKKYumfF/5fY
lkUd0gEnQOPrh2AKIzT0Lhp7psT3AgIrTNm0jvH5vuNYVqQDxE8LIOweOKQnq0cP
NeyQia9AmK3S3/WLPUR6u7U4c9gPMFINNwcqjPRqzvxw2dALLPZwcOUpX3ZcMN4n
QoFygnh9z45sKKUjB3fXjUNmk+W1Mf/cWQqXJL1/vcal7muj7x7FjzIiNDsW0syX
AXETNKzzL0YlyMIqtWSqbpNR2Fq3EJa8H4fqvf0fnrpkgV8ekk3rL/XgDG+a+E5g
EQqe/PfAf3brSQ3Ol+XbbWlSghoGOTADpJBQRToOlb5/GsUvVaKFw9GcEXZ1IxpX
ZQbHH/A/XkKcl5RSXT6Ia6DH8DbgxiCfs2dABcGynQf7kC9zqf0XcJIvM22iWfC8
PdREUoGJUUUOmzdi6AzdwyDTF1rXAVVFRxSaxHgX1JSm1AjX5xdSM5dfwD6HJ/6p
RDvv01+67BwfYcQq4w2/Jy6xoo/qIWHB/zqnPjhJdeFWbSq3FytvWYcfEOr7oDCE
hNT1GzPTzko60pfBBDM34WOHPsOMvapY7GAGeHKUszwFJTXCJ+84Mp1apn1ZceLI
a4ma/YmofydqtpQ1LjGxIkvp0SXZ8c2WW9pBdWjV018cFtWWGGzp3TWWMb+nZhR6
0RlHs4A2x7mtATNs7qpOCniY0a9nX3h4LgT7U114gp5emJ7uN4ln4clsy6/qJ0o8
NjVr5p7OaJIcbhiizJ7QvoWr6ueUIQaJAc0aQ0Si1ceLjZVsXfo9GMGycLFpgWQQ
vsZRu9QPOuhH42BPf/rUD+dElh4nNke5uXAuLeWE3Ltz0Roz7NHTwHMqIzpHXMh7
8pLgUWulApwxDwMVePXirDi77kO/z4sXr56Yk5lxUIuQBlzI195eQEWNFYL55Ul1
xSyGpahq1OPokxaroXECszhPXzoFXwQabeB+23ZbKt7Px8+fVOORiqJ0++JZGJr2
Auo8+vz9Dc06ljnP8OaVCr6ZVRpUFmAyhKg9258eIM1RNHyPcH9b6fIbs1xw9tc5
AyNbfw8yNtCDbMEmNers619iK3TWmp158NdYylrQfA1/p1phYDXOa0AvqVrhw7rY
OTrG4vFFJUU6nQFopyVJWWHcHfMwE9RYwOoASBK4TKux8JoElCYXW8880lADB7Q7
/qZdqUSsuNmiWlg/8jPncZ3QfWQHBo16/JUR74d7d5A2FI1iooysR7z4+or0JwTD
9Xs9BXT/CrIp/zm0XGmiP6Rc+rvgTsMfKo2DfjGFn1anD5g9jRwK6eNJLtDF1V5g
UKSkkrI5ucSpKfWGL7j4ta4jYmb23354KTlgnCY+Z9acVjS8uuUCU3rljdLuePM+
+stBgtMJ3zDJasithjBrc5Otz0hk3gKykZ9OkQHt4rebejz2PFWO30fAWnO3SRdL
ekI6OmD9Ca8QN2L6WL0pBscJHjDVoR00OYUVJubJh0cJr7AlIGPWqJXqtb2J/zbl
LIDpBPXr9zR1JZ1K9od3Cqb2WgSevXfXxZIjEokbMZAi4ANNv73n5sbvs6l2Fjgd
ph8Hj/746Vw5gNEKiSJMS2KXkqDDe/uzVZ7e1wyHS4TxCkE6ekTanmes979XSDpB
ZOwlo0KkZoxPDQKtCy/GhxZshGPfPGTfk4RYx4VX9XdNO+zBXoICYmyeHHr8DVRb
8B4as6OYvgd4SzSA0DyZhUxRSEHHl5K8OyGwtyWzj3ItkuVAlao7vx14REr3g2zU
5pdqMABgeSD+HvQneVlMF5hj6K1FC7pa0K9g7A3m/kCyRWsu3704iZt/Ppgq574p
AZSJr5hWilQrLYnqQjF4dvoptTUdC/wkyAhf25jWXntVPdOz763NKSlIOm5zsUXs
i9tkdKZ+LAg9wIuMx20sURhUeCUcfnhcXrWnN2kerQo+OeSPgBk+hPpPUwwiDzJu
MqpZi9mjaMHlBdYQ3Zi/CoaiCU5Z4KN1XOxulKwqiStH0dNNmcfmRyqaSIy1RNr3
U54xLF4uPxpOylOiqa10XYcHtEU06lbm+H/aC4xpnXQLIeEtQDeJz5GQegwifDiZ
Y0+3Dzg0R+sBFN15YjLqdW3GLHKVrq/uvuCghe/JSI/d8HhbGbHHoRTo/LvOpJGc
WHJJLAxKpt7BdFYIJHJPHsRyl9ELKqq2xeo3Rmi29LPGOQGQ9vF31RmT3rpzwaFr
/QkQAvnbP1EQey6jYuqXa+mF++lNP2ngyXceHhHbVVX3dj69imo6itGaWSgeyF2V
LDoIMzjNwmBrG+UH35B/+YQoRvVDCvmM0EEg6fjfdhgdFF85wUnMYHyrc1ffONQK
i/BB+Ys9XVf9h06eKanzjPJMboR/uqxyUuavA16mU4vdgfx3r+mSuehourUwb3n/
wZN+rewUPDFDbkmmaRH1ufJUxLbQdlR1yUdapPbvBpbzY9aq6D2h6hNRKJoZi0eI
HLALoOs6QjkIFBy3Xpj0P8p6j6Qv2L9Esp+0yx/+UIPHNszpF/sFSm52g2P4fbvh
4SYzWqZccYqd3vtkZapTiHxTuECP1SIVjzmsf68/b2hEtBjliSG7H9e64WctGStr
mHGkFMDP9wREpPyf4/4OB3b7aIzdMR8BTu7wrjzVyLROIp7+OA69NRK6Pxi3nE0l
VE2lwJNSShzZtwsEbDR7/hs+Mj9lN3FC85X5Ppt+M6UBqEZ9joiNtmWzoeK7HAAn
BUuWlo2cbGt1QgpGhwA4Zr2fmt8HRkHs034kdXcGJX6anul5rLEBGKAuDJx6clXB
r/wYizCwEAIURunH3OsFq6WdCgoWAT0tMxazeR25IA00MybvGuv2cSdVc3ZAMZcE
K/Ey8KRT/s+0q14BdUmq6VdXuKJk4l4ZbKHGpHEUb1RhvhANTmnGaWKn0GChDVNq
f6gSAcJJMhf1e5Y5tk+a12feWByv3+LfbNptdyPY9IPnmdr8roLQdYVGOqeA8FAs
clyR9eMFdEwcI+L303FHQsom8jaK5pqIyl9l1jhBZ3R1UFZXinAiY1FRoaCZxLzN
DBa0R23Lz1X4Q+9NKqW1w6/C6eJp/rh/OGO+bceAPmE0uueOvDSLaJm9DweXDNKK
iN1E9EuWM/KGTL5ga68RDM9yUmY5yX+ZX5RIgrEmA9YNyNon6gbBXbKJal5w96NL
rF6dL+yX6prgnsI1PlCJqe7fSo1+ReM5uXkBMmw3+/5gYPm0xXoHaE7UIvWjKrIr
z6+x+LBX3Jps9aN+6AkmbPBhXbbcOCOq/D3EWgT1lBk+jd4HCDeYnZKEKxE/MqQr
tLj2bLOmQNADGij315PXJEGnl53G6UWE1wiY3Dd+YhmD5x/yLuDlhTbphgW2RPp8
8iuaZIKj7+kUn1mvYsfGCLyGhqJAHeybieNIy9LSySkBqsKSBiFWhqcZyB7l0CWs
ATDqiTjnzqC012WvgWG4x6IrBBhKNxBhFmtEvpNRJGJifRcVjx3pf2T3z8z1Gu6t
KTa5C+KxxEMDFjdmz+olrl7oiq9hDcm9ayA2386Gj6x74ZSppzxPdKzy4Z+qL53J
ki5yLa2Nm/58hJjPZ+2a1BdqZ+M5/VX8Ue+jK44SKgmkkhFHlK/TGUb54dZ09CTP
imwovs8l1m/YJDJ/RwS57FxQ2ytSOKcIwwbseIUcQt0mv5NUS8MjaNvxYkFp97zV
5jhYh2RlUqRwgou853S7W5GWlZ8o78hN+tkbcLXTYWaQ+IOnQVtVs00LAYTeRq0e
dPpRPJjeYItb3PEsKOp9ejJomASYbLZqQxf3DIuh5lOOdlTKOo0RCh4ktsfO5WvE
bGpZffo3MqoUWDy/YkwZysz9LumrdcGPRASsmgAGUm+EALebYnp210RhyMGEo1cw
u10axZBrdSnzgMmTfrY1V01nfkgLhp5yPaiGmdEPkCbi5MT9v0oRQlo+Z0CPQqNl
wjo4ug36tY4QDJRMUl135DMGqpV3U1c+jp0CZWzwvI4gxCVP4q3V9IWITYVfhIip
ljYWYb2OMlXWlCxx9xk0M1YOW90XvTKsnCasuCdSFAca8Nh3HST7TbGSb4HHxhIJ
S11f+w8sYKXLtAFjilRSxXjfhLLM2K4u6ZE4sencILaIXiJA1nk0CzKw2jgyZStk
VWg1XnSE2a1tFJRLi3cFzJp98G5BM2z0u0g7foB4s2chr451VB9/TeStxNSOGLZo
ipO57DCeymzYQ2jvTXgU0y/jVUc87vRmNZNCw0DnFr6xtV+OoBaL6UpoKZ8FNuhO
cjCKZKMYUatdAAJqQ4CwhvGfO9thJhD5WpuY2G5CPRcdCxP2hamkUkqzUpV7JWcm
GzxjMdFCSJJu40YT0k94Z6y/xlJR7ZC32hGxIHTTsGsSFyS6+eeIBe92NcafwXpg
9b1/I9A9u0l4tr+yGFiSBQy1slK6nLcMjGLtSfSxiQDe5q0r2AXw1FoxM/o3USaV
1jl4LP/hvenrVOYOVFlalJf0RuLx51PfXokxkbqJzBp3YKvdLVt87Sb8ZRkcgwIP
5ABUmSumXY7Td+x3vgh4aUnSBBfRDiXU+NrjR8pJ+hb9aUA/jgGiC+gdBRU4hkTZ
VaYoupwXoXmb7h2JK8Itzgej2iG67r5cnbwODCLn5Q1SLQtzIJvRrj4waVEuEcZi
yS/zSyO09QFVF88fTg6zXEI5b0fELxff0+o+lkumLU/WfEU1YP1F89u0jOcnwnMW
I0qhZQ67JzUwRYNJM8ykLnrfi/QdrjGo3aAGMG2GOROWelU67SHXB/xMvWe/lFOT
rzeOn491ICYqexs1v99iunG4rRwy7augY4vWqblKqn76MoUTLqc8wCwg1bIveflt
4AX5HIVtkSO2lfyb5gR5KHtNcnJOeOOGiFpv+LOq2plGnPp1NEoxTMqs+RZzLZ2G
1XMHoSMk9YOC39yeSLtHuHryny06XsrMifNLGaYzHS4XOGPLwVvww76A/MTQpDIw
yajs/W0YhLVVhJf2LphTi4Obr0aYo2O/1jqsfysCx3SoniHFDRaMJ67hdivF+g3Z
q80ZuWeUEIoTLgI9TjRzNUqOyXVZGh/5CqZ3HRFhXEvtIyNleXPefHcsygsRnO3X
qO1DH2wtUZTis1aeut1uFrUje1ySG9Es96ZWAD6TNjILRvYvchjnpkctRoFx8QTn
+ABXe0I6TeeDslRnhTbThSbhweHzWUMyjHIU3RCTXKBjbnrZy44+v3CzE9L1SqFy
ikSEyinHC7HEOKDzL3wmlS2L9du2OMtuARuKgY+7+0JhrCdccLoFJvDj0Vd93R3b
8+2vXZf9vlNoYC75Xys/iFZK7nkp3aUoXSlsfDBHa61USI+DekM+L4IgXC4CYFyc
P3fTDMbkmUHjcd6lYgc0TrderW+5Tggw/bWB4QUZDTOSZ+HxDBQoeKB8GDneAxxC
t9ns7N5xOyQ95V2F0yS8OBzvI8nkTee5y2q1tJ8D9OybdabaUrfMy0wNOwcQgMe2
XSntQQngAk6z2aJLPOo0y3u9Y6jINcy729hmMgr/zWvwRvB77ofdufvq87LCbYV/
Ln5hodEauT35wIIqpduPWyfmcnu/7TgNqCNJUS4sy4eGoHZ8O+vfUnwzec49OPe0
dBUWgNJFeITYNEHCEv0CxTmpcBkdbHkAoTHDPrtRK9X7OJHkF4eE7ZARNPKImSVY
shE+teggaRAFE2p2Txpl5e9zxKQ6rcaW16OF+Bh0cg5bdnxJOvU92MzVAZALZLrE
gy8vQ5UgYtPp/7yQpioYFfaug/pnpiYhe6mEf0vjSrnGU/VsBKX5hlR4qNptQXUo
V9CtZrPRidb34KDLj4NDPzL7j9tFBsKtROLvLjvt4DjrQaIQcsSiTtViV9IsDwTv
ViKN4/yI0orSP/n0qG4hdOc9FwbXoU8svugZX1U87+J5QwEyvc9XgS5biTQOaHoT
lmlLM7UY1QA7ZW96h0ZKz/qIPX+N39u3X8Q37PZ6tDD16+SEsPNW0lVaj7bb30hs
3TokI05a3TTK1GjwICW3ciZkLqr5hjWnUHtPwiZQD//z4rvkri1a4I6Xqc0/FwBi
gXmoG5JrI9H47SOTIEheYjfOAlbDH9BQUsHMLvjdfozYZ1spou9xc47yv/WRCWmA
dtVDqOGQ2LLW1IZAygujHD1ji6HQMcKcXY03TVz20Y0IbaVqVlEfZHWn+XhdtJtU
TCxSms7zAZvdMLCDiS9MWv/p7IfVKkdMCLmJYJ9UezMQDr+Ug/627a7vX0Ib+qIn
PkIUv9l1BHPUeEC6++eisauZyGXiaG07EP65k5i8b0Lp30y4MkXwCDGAq9eoizzN
s9J6/zCxh1RKIzJ+DSaTnTI0DF2gz93mUfoJOzSaZQFM06FpnhUmXRqfbVSbY6x6
qdi5V7sTSuHlbMFAnD/0hawwVkm81IIW+ybifvWnLd8gpfz7gkU4oEIC3h0V0UeV
rDZlXt5vnsftwBOlE51Wy5a33zB5TUmBtECpAtUMNUlRCnlygeYt3/Yx3j/gnU7K
1yLkSRFPDn7c341L3Z7OuazCqu7yvGXzf0wycOhrHlXyqKygN9hy+FhYg/NdLKFA
7O3Q5VrCGlpZwWHSRs44XH/V1NyNKo6YyhyLkififN3P/1k5voG4/wRl8QmUHvDo
yYaDpdVkEOT//MC2NMM1luHZUMmL6cOdUYBvhMjdXGGn7dazVMudapH8JKTQTGxE
YuBiUWn+iLZ495kTdRemsXSFdFCDqWNKvKCWvRLM9w87j9roCmLLUfikEyf7gRBD
BqdM3b0MJTV18PuRaCZhpsnmJKSA+1rH675ERiO+AV9fEe/r5Wfc8aL4Xk5WHcpA
9NpOy4v2sZjknU/u7VGMO+Mkra6zJ/xKEJkuGGmCIXYA1tJMxGR9XG7H05iF0Im+
BFZn72dxbyljETWYSyQqtILWizqpvGbP1EY67JuxJpHVK2P3aNf6+eCnd5tSFaD/
HcZ9KDAkfNPqQiI9wqU/UwOhBHa1v4p3tqWO4HrsfbE1MxGPrYkc+yYOEXGEFhsy
MV+5s5qO4Xj4IeJsUWCMNhTwGm+Y2lIomvYAuyjT6rckTnpk+lwTN8E6ZpiqQxsq
mPITyHdHWPO9+C3TmbcFYlXCik9DO8FDKQXblTIGWunl3rS01jtyGlzOf+gr/G87
NuPGmTYbFyk9N7j8oD3lqNtdPbDJFf/DRJ26nc8IB/M/kAmLMI+tMRXMvrp6QoNU
hgVYHAK17EQN75U+1Axx+q5mQLRV32wdmgwtBUMz792j4rxdqBg77EZVH7nKMfnT
v+Qp15At1AZnRJLea5tKBB0z5rM4cmpbpnLxdHmF797H0j0qJUQ9BSfIP0zfpf/4
ypAGwu7D3IpQ1bOq4b8SFdV2TUYQfIbYCVrhVPXG8kj+Y7VqX1mX5VeohcGQrUH2
mSx9S4tR3NRIq1Ds5/IAOzA6VBJH4arJA3r8kJUsW1WJVGd/7jJ5S5GfgKputniz
kNZ2ZBDH/2F7rniXUuYhj+BDh62jF9T/Y33Z6fYbi7mHawl8y3h/7yzxfuXC31iP
rDDMT4qOxz+kDerBo19lx+Nx1l6Iu/d6YgTFzORELXtuMLXlGVylt7kxoQVDC2GS
mCv2rHggtVdGjNw/MlxfHWpuQxR5R6vDGucBw6zdFrJQTYvUENP9wkJx7cvccpX/
S/4Lzc6oRA9kheeR2LMOU+1dHJl3rtQ0l7Y/o755e5Q0XjucW8HY9F6EroeNkGqa
7ntQ149THi00B2G44/fuTsLpsJ8d+f4pFapnQrtnG3lK/OPoLUvblazOQiQfry54
/zRnXAS50ISJZTmURQDdcwuj6n0hYyEXbdzKLL3vCPIkIwjadvWTC4x1uGWDyS5V
ZtGwmxrATY6FUP/CZBqXk7uhmfEo+KkBHy+g3SXKfaIlE1HixW7RGqroAi6IXlCb
4TMy7sSPIlPkCuSpm22xqHhCLD3E2gHPnSntJRtqQlMsMpH0XceZI3X+E+pA3YQE
e3txvKhHrXsWyjmqwv86y5BQ3sx2NZVN1Fy/JwMszIkkEpe3mqbQjA4SU42BOYUR
m8r0AZiIwtECBo4KCgNsgP6w3ZWJ/aklcd5PYMnK70aOeP2dDud2P46PJZbhitsp
laF5zeg3InP0PqyBiS76iJvZB5tDLh0mhaY7qIgw+v2o2tLXj2qJ7ehGCRgq2TKg
hg48U1yLzq7IRAmALG+8jktK4jD2DL0ZwY2yCg2bZEMhoqnIJ+LU9epI0Lt4rfru
sQocLlnLYjTKBeYz6vUfpXJxzOD8cVE7sOSGZQq4coKrnrnOCZnM7foj1PVHHd/K
exNMuusw4KEgVoC/y16TaF1sblIwkg0DRstLEUkBD+pJUaXgyDuvO8Uu09oEGHSw
QhUTUtgUBR76yKW15h68Vys+toJ6knB59DRhhKYzvd8fBvd/1ZFWlyzHd5VbmUGA
hE+ymY0i8+g3cvXdprWWPV6Lh3/TWgqivaSAPbIOgAwBjX2e6oVOJl+ng0x6BxKv
njx8vgK9gzI10G1erM5Oz8hKVfaAZa/vjhkKkmoMNOA2Nh3lWvK+9Rl0LC/S7fNe
P/Nz0wsusnxoErN3YHvYMhGJPhG09IFdy0j42q2su0HNOzUudbhseuwq49wkIfrs
/qhAdCAF9cDU9JWFlxq6g9bdz9MD9ctSEFevpneBMZVZEsRFmGkuvJ5RRshQ3hEC
GvQVlLm7MV6y93wN7vknjNHBdE0y5hmMk335kQEJAHBGnPYVkhXohU+ayxJ3OMSU
al1nMPCv2AVNf8twlepL/hkZ59371AQRUrsIkbcknW66+G2TCZVAY+AyQPXTmihV
31PQsfNwE1GihSNV0fr8zzwVn8Q2oO8TJJga5jFnAfCuAz/im3ts+Eat6pAy31o+
4xgwsxzN8rHCe04aRreI9Pgzq67nNSTv6VeP/+PvlpZHPjR2rsmK2WK0yka4rNVc
FpYkZADua4Hth5mwsSIXc68GDX548KFzX0cy5EkOy3BPib+PG4OFA8uY8RH8EpMS
dcspM9KmuIs9F7ATciJj4heoMHmJ5+YHnYf4xeDSM9+6Z1y8DAtkHuxi5SXAnbrc
gX4IgM1m183yhVGFKbxGzJT75rAp3WT6K0LBbtJTPWlPVGxtS2VZtggOW2tbMNqL
bR3AlK8CcYaj1umBmeNk4UGEIPPQmmlVpAfWuxdtWVdiNzHHDDSG6oC2lFNIm71w
M7yH07e829oQZsQ/0g0+irLOpuxXLaLz9bO1J/mDP8sdRdKJjm+zrKft/799qIxb
WWrv5ph/K4S35nrTsneTzYrd983gjas4169Dqsaao+ak5Hl5se44f22xJvlBHdfB
5gBXY/SjWfD1cKkSb+slwDYClfHf42h6gWUXlcsCGxfFBrEC66xsB3N45M1IK3jB
VA7A7jbvp7K9S1gnCgDkzjC/Y20mKvxjNuTY9Bj8Pe2Ma/SVVWb+a8YG94l/vBvT
G50dqwrivzmTghBl/NW5fSaWAW0ybAzT+4ohhOywYtPKEk/EumejqLBp10q/J0PV
g70F8KP8irGWsMYrv3sFcrRGVNSjZdWTPwXiMZFLcGvmf5Ge41gF1Sa1Xb3+4jFY
FqH9b9l5IpH0bOYlicNfKrGO8NYp5Exv0hOYhpcLGTuiOWWsQV4vPLgfjA3iCxlG
N6U/Dr6DjWCFc/5onDCMzCCavAkXfOs7A5yS8eER0XcCogWznoHQLmyVNAPuUqCl
H5O5ww4N55ajT3n3SowHB5vBDpBjk5poFF6MciPT3GZGVAF+vJEW9GdefID8lEV8
OfS2HxygISVHn1NPJM9As09DdWz/FNBln7oLLpZ2+Fe8gTA8QrUbJ48CeH9+ow/P
ksdS1Rxt1Sfi6jeQEkYj6XTRnLgLOsxpk+qq01LnN+fEJkODEojPiR78T1js/U2D
z7ZJG3t3E0vXA9/FBv/WUmal+LsZ3vyaa223PJ2tmn/mEFo+PZMWHlAVaWIRU0si
AaWtHJLAGH3NctrAt+UnimOgV9MPo/5m5dFyazKWXk7YJ35X/wtUekeJVES+u7j+
fdXlZx/eQT55UgfchFKSrYFy7gKnNixe5324XW6PGF/H6fOFXlBtMZKavibLCtil
tbw4QS5A/zybcfmOuFKtUJKKQ6wGh72LyYxw2x2XmHoghtB4AZqonNdwZgUJAS1k
WihorgjFZGY1dur5iuHsMgKgKU+JbHTU8zVUoX3LDqRSpJqya49KXwqZQXE330zp
AsRIx4FBU/9wTcWeyuJLjGsVKzr+sW1m5p36XFtUzQ3/FWxOd7k/JKHeGDeAQRp4
CDCSITZiU989CrMo/+54Sgtlr098VFMOJ94IsKPVTzM09QFIM+genZIx7y7imdSg
zaYcRWNJHSBTPGqEqGttgf+rx0BE/0a5nlx5wBW7ykfgrZ4yzLH+yocnAqefnJ0X
F5WmuVIudxBrAYcNBcuwcKQOynVg2ZGxg4BAtJWyfCRCnwYxqHmpQRiRSSJKAo3E
SNOyfssejp+t6HdmFEUDghgEHYmOiI49dDNxomhJ/fX+197UnIcFJaV3ew8+6ln2
S6QaKijIsgOu6Fh513/S+CZ7HNy4ocdnSOdRt4c87YRcf1/+ZS8mCHqKIheHn4So
7Vidrib7uFvDOIoxG2FeAVnOrt5IgxsFw/WFE7lo2rGilPGxk2d+TO5em5ZWpWx2
G1nk7FNfjiLjisCs0z7eRvtJikzzXH++LT6PQlsdgD2I4Eh8FY3Z/gtYPoF2iDM9
hE+cM3MKBoKCNXfGCet2IJH5+GQBZZ9nuy7CveKVj00+FKGP7JgBt/dO/5L1uV3/
oIRRgsC5F+hIvX1cIG6GV2wmLwXtQdF/GFgkIy2NjCg58PglSKfkHB45x59YH2lv
ONpdyma8Ww9JJizyvuO/AYz4S5mFvZ24KJBNRNigNkgftvHrA5oYzI566pKoyCPj
zbxUDn70NUjGMhRlkqLf+NP6I3pYxiVb8YerDFi4eU6+Ojhp8547JanLj0Txu6qs
c2acrGvjU1XUsoJ4gBM9z1I8PgWn96l53b0GyBsfni4UCmO2SEHiMVcDulCVXwI2
BHATTczU4lKwiYatgc4XWykpgb+FNNLLzMV86i7//GkhyIW2av5UlDeVwjpzw0Dt
5IlJB1kDp8Jjh0hOpLv1JiVDYYwAsbSq0I33vM1oGt0q/xNLUc4Ib86yfAmca6qy
asiCppqjWEgdJZ7E96WzGpBMrWeyNjZWRM44iJeEQnxjCxm2jT+KiVWi/WicG/6V
u/cpifD+oVvugNDwwgJVk1+/dD6vXgt1bcUll9u3Tf18bSsSsX4LegXDrNtaNhFn
glhEMSGEeu14sAqHGC0aM9/cR6FxD1Z9JQdZ/VtHVlQZ7aCAUvkeD1ClANoR0b0d
Vx3Li13t7+/gyTWLNzVeIHD9r+QVaL8FyBI8EO4qoq7BZTap7yOicpdad2UhNezn
GGMe2k4RtakQJYtPwAxnyWRuDCPtkJVjq8FbXzqHDss+INqlQpFWX9UOgmHJzmSZ
wcY+s1U+bT7ul78bf85MHZcvubvsG9IRmZ3M7Mc2ld0h/OoyBIq/FQG4j6pfpXtq
+QBZGrufRFwqIOtIHFKEjdi/B9hRkiCwOeSEMC8w2yDGmKLrHOgcHS5LR1XNxm7u
ZpRZf2AdEJ9zSyu+lqRoAGkTWqDe3nx6y8DR3a21O7n+d2hDkov4+r4KKFVdVp40
p+LnAFw/aYlrkGJRcJ5V75OKkN+U5FItiqOlFUV0FGBw3nHOaeJr2depvID3rkHm
CSoVNn45xl6j2rIO2dH1K8lvZREKbItuGEW6QEzNVlHJLEfH86vDpcKMbPi3YRAi
WmEYNm5BB3nm57pkdQqyrsQDOwZhvH1WW6UN9wHLvXgdlI0ITnmMBd4m+abfZqMU
qR/bCGcx35JmXvusAobsOhACvOxURfCuh1/1EUdfT5XAX2Ob1heBTSAoCHxdbfRu
JYfNiyCCpKt0waBpo9AMUcO8Xx2NULT4cbREpNmdsPNCx8kdNwUpbYhdzFPfUiB2
lFjADAzxtm8DIXJlC/fBPMgW79YComSs1HxKqup8Gqu9JQ26fWEBVDKc6V6FCc8n
iGKs5AOK3Sc0K9SaEPEuJzJ3Ho0M7h7/wyGwIdXHZPFuJ+puGQ9GstTWj0uv+Jxu
8icBTRcoYYzqkh8Wp1CPeK2Mhhc2dVsNiYDfxfufjotTGiSsEOuwqut1fp+6LACt
kU/viT4I6PN5CnL4n3ldfvCXNtjQcIQD6tU73J5+Lqtft3raThQNIa157wsYg3pr
pscSlT6CrYa8gvTBY8nVmPHOGrzdcYlai6AGPlB2YgHiVNd6r53N+/AH3ZJtE9yD
N16CnGt055SuZS0JujMx75UngXWDFETPPpg8foS69VlpvqW7xZl3tC/05/96nDWw
wDF7k20MQWKYpUdIV6KHJK/YwDHliBVG8R5CMaN9VTxzJwRyAzL8wHFsx64ld1SX
FeInwx1mKEovgetdsBz0IFBt7QUbHnq6v0vojL9YSxYQuxW9kj1C7yW5GgitbHQA
lTnSUkMjrFYTBj5m914WF/5rVn5bF5wKY2ykH1s42epcmcyXfjAsLKNR5rTmLLc8
J+7Pe4Zr88Fcb7VT28oAXb8w3pCetQunhzxh22uUMuvtPgipAavWMCiWhG2JaBU0
0u/hxTSvCiLbZ/78c4O4qYkg6pk5hZt+kYCqRn+aEoKvqiSofScF8l04gftk8KDJ
fmIQkqNazif0goZp7gmPJjMRbNkXQ3DmVM6qrA8gfzuuk9yI2Hyp60S8eaInGatx
j8di2Meubqsu2R141rUDiTafsrj2aWXuWI/J2bdvhj/NJzwMU8XVA+kymE/ga34G
n8BN8cKQlAbJjWLDUidMnUozQ3YTuHqMrWdo74lMYFDjTIfeZ4TPtOMZ7P3F/Qid
3D4y9EBAst0IbhBmhvVw1k8ZFahi6OLVstZy61cNNdX/kFk8R04SI6xp0AYYGppE
LoksmVuK9B8E+T7kxhHFOly9Z5cyUSDK3Jd663bhr7got7NeoXMaKBWGBuo/L/K/
oDYrfdGZeHvraNqbB7sSnpFvfgSyZPrFsv5THrQFxW2+wZPeVdEmPHHG+M4sJ/+R
SLMshtnPN8lHun+Ny7H1TZcXHXoPFMdYRWhoe28mB2/O0TkPTSEqVN5HeakLSR2g
CkZBThYgVJnn/2WfXVOv46kjpGEJh9TccQow/S7twuvBs+9Koc5Lrvi76ziyoOEM
RXuEYcmZ4eYVZ0AT/zMuaW/jSgAjqfIoDKqszMMxvM8OZPi9ltLYtcGiJGyRZ647
Th+wVL+DxcNTAQ/Y3CXKXpO6N5xdGE1047EKGpnJXjOoB3V3484bR+JeTLnIyP0b
t6aji38tNxMwH38QvGmOkxHaWlL94IblwsczIjYBRyqfLQ2mUeITPs/8a3CNd1LR
EK/0kHFG9lCRK56t4PeHgUIgQB/ja8iTyF3x3ilaGGQY3NU0RBccchyODmlffj6w
2SNrutsFxbhRMFkaq9NVVE2clWk5nNj1N0vDlJXT0Fup4RwAV4unm4U30sK4K4Pg
/uYwn1bAwm+xCRWGAkBNHEZKiXtjS1kzx4FUP8zcT73EY4jDc9SBf8PBMfSrpCsZ
z1QTS/lCFiQDtsF8/8fWlx636rkm19uOM0sHAyrMqE5vAKdLNZfyVvl+1fNiPddN
mCLzGU9dSQXI5m1Pnpk7mdkLL4DneI7TQtJI75kIUzNGg7ghKeACFDpLQIRm+ucI
HuoMrZPqjCA0kjUlbMsYELVQm5niI9ZRUiMgWxSG7FN7gHfnWDHY2N3mgoR/WfF7
XJzXUzDUOyDs1YODufNjC9S45QjL3ADhzM7pHLwTM3UHTa1l4arSFfJsigNwQPjN
JtdzN95/f8w2aTGy0+SKd7E17+SifT8HY5RTfxJlzDwbei//1ueaCjThoj74HKV/
fq5bgDgSVVE/pilg/1KiZVkKf8qBIcrabvXoc4yM/JMk9WP0pQniMgL05gqgQ4VI
x+escOhpjDn6fIRgD546y2IefhMZqGl6IG90JXsbaPGOdckN1JWlpSNbWkFrmSQK
QqPJgm53E+A0ZSdCovBPL+07gu6tFNtxJOhurihtAj5qCt4cGhvhBbMvTMrWs1SO
qzkjN+F/yyMXseZapKK2T6fgIaBTaAzsyzDxQhD/uTh34m/giHHBrv95ukTowG+x
/5wy9rPXoFSlMQj/eoTh6gOPsC4j6fGe/JUFr4v9E0MJXUrlOSkOGeXTJigEfVod
hUvRfe1Wr1ASlMdETZewf58PMnkUkK+KX73SXmcuPskb1iJiXFzopBdRCvpzxwvH
n4BvsiRMMkwEUcwtUYvlKac/qQ9lxT42UC4mhgJ64dGYf1ZM/mmlwrtwnLfDefqV
/qlr6xoyp7KVeBO4W6XalNJVyUHGzr6BYSCRvcgJ/Zf0UyotrHaMWZlfdKGy9G7l
KPxQShcvqQ5VQEK1w1aRQx1OT4hS8tume4iFQfLgTrRgWpO1ah3ciQYbSzV11jnm
CJMyO7HAtAteWRovSNv/tmnzXmYcRQKsjcFBQ8rIK0tCatPrcVbmmjy5NK9SXPDc
aHTsw28BJa1d8v6qr46k704fk7LXcp/mubR0JOA61ovFjUNQZyfa3aRP89akHDAD
is0mFzwxX3dKoda4uvzBERRa/BIc9gQl05KfksGq203glQaMBPFEGg0RtkL8kfd0
gdk+iOSnWsLghr3oocW8r7qNoO+57kJ0puS1CbjTignuu4LG7lk2Af5HR7gMRAXd
dD30DTfszr5wxEPLMf9Pa/VG+XECjPgtHhLiPRPVDVs644YeMnmAl98Ce9Q/I74E
iLKF2G57Db5vCzmfpuPye71ZCPfIL4HRVIdXVKw3+91CIBWxL0quoVW+MNkp2QTL
IA4Y9rHFw6heItLq5TWCsuJpGOGMWpA++0VwrTHwxfWhRf41tK87Lo25IxzpH+GF
3KKr3nkm87WzDShg1mu/ObfYrG/k6duRi34bo+9vYiuQW1BN7n283+WU13N+GaQn
dNaVdCTyrFmg6gAD5hVGxhiCF8qD/UGbwmQBbGGzt+enJwjGV6lNEpD0JKQKfgln
2WBiVmR+I3hoIixvhmND3CqAgB4DJx3iq8TQQA8gqUWc2TTDO8CU1qCwrq5yXWe2
TUtA9SDp37Qx/O/DKpaSWL2Zmfd5IUpLPRtjQVpV5HvhVUmGJILIV3nfZuKaO2gx
mN4A94yP+OOA+eMqj8mpFM9JaqTbfhKcTeSydmcO48UE9vG5bJmzFoD3IYD21qfL
Voa1EfaXMznOQ3Nk99oyJWIlTA+dWF8NQqbxBtyd/PFvopooBa0Esjp1iKkcF11P
zV8Y8JqnUnYFK6wECPA35g9WK+7WTxl0ZaLZk91ue97XGqyC4c2p0XCP9khQlj1A
AQrS6xuTIIF0pT6q6i3R23g7EhXC6Q2/TiGXyHW/Oz84lj7BfKVabz91tF72T3un
93pJjSrZnH0Aq6XgUux+vNYEqzlVymLHRIdyionWIpMypF6bX0/ijNESEIWXIASV
bSvODTdEfh31B8q2lcxuhlkXmkxW4G3MOmrscLpnPrTdGgSPj48MKRWV6xRomxRd
hUke2zqdPKo4mdlEh153mpVRiRoXyWugujNMlP+iQp0DW4+o90MQ1jW2dLhxpd8V
XSuy7OnJ3W+SbDbuGKnGk19XKtT/MxW7ibOLvUGVTrIZJnKRxyCQNY5SLOwsK8Gz
9A1A6GzcNSxYW9zg1X7gj9ZUJj+ZrtsMRkei64FUg9EDtue3wD/A9UooVKJ6nFIi
gK1lUqbWAJ9GKAMxir1NRvBba9t8WzUuz77ItLJskhVZZhL3o2eWyMzReNaoOgZ1
aGmeEHpE4YJkUf7ACFaIgEw+7w/rWLJ/gWN6U8HGv6qncYNdtputMB0w0W6tqWcr
9w6bONkBG5SQJXWXn37gtgoh93aEeTgYd4ryt+L/U2iq0pcAX4uufr8fPTj0v15x
brQjtnVVUl+hNqae6USrfReWUkWMJ09qemSq4oeX4+p4SXv4S7AuwlWczXNgzXmy
zOFUkI9F4H4Adm2pBDqdJfNVfGVGiVRG9hi0LJaY+2/550Q2M1za5AV+soxvO9po
jdVU4nrfY73M22D0iGlvQhX35LY7Lj+3PXMj+I88uDuSAuFSH6On5bmg9365fJKB
IdD867AoS7ll1xixvRpOlkxf/nWxct2soNzyKLqwmp3+IYWuh+9Nb1d7NddNUm5R
E3u3nB1uDk425RFipiPPMildoC7hKjEX2QK2gyvDXLPrN+aMfhXunSoB2/TsB6r/
VqlVylSTsA17NofMJXw1eWQjvLGz9Q6+AgUJ6tp3JUyMpRh02BjnLU7Qm0huUZy3
p+s8V2rMx/h869MXnMTaHA6elJDee28Q75rnblBMRZ9u8IE3Y7T2dZZnwGdEUE03
qPztMaWQq6Rt4VVkox4t2t8zwwIqMDzv0lTGqtHQv0EGwNAFB/N+wCnOdbdlXJZo
HnDSjoxCDxesCCbGIlyM7YFM2nkuA2PIIitlPQzSwSbBBtOP3kL9U1o2SLT83I4q
nQx3U9HAoBsdCLc9FOulEAlYwJXUYS+MaqZ17+plnJ4XRC6QPyisK2AFuJUEN4oA
Bb5DA2jt92MODdx9JkkLzzmw2ZKh1TrU4K8EXvQ1dpUxDIb/+Aze5VhfEcn4mHCX
WqAuq3r55tBX+dIGfzV+hfobX75ZZ783aPwAiQbMXfrZBfYTr2WDJMUAOdl0vaaU
q2oZeUQkH7f22+nxPvGENjdermzA4gpvKAwV/xrWtu/eSfK5NHbbKmx2k4N6/pAX
knsSPtTiUQ8GXF7bzbXqzsMjSZGOdFNNihLtrMjJk9rM3VH48MoBulzxnTSYOyCx
UMMjR4V0jCzw0C9yvYumR0q68owwvGd06VQ6KoH7BxkUa96vAQDdHi3SccqDLp5L
2w435uSuIeYkY+aFzsfYclO+0aTzVu6cz5Q8oxZ8thP9zlhNqGrD9vfjVb7+RVhq
GoFq40vAxxrPAjyxO8D+YUKB6dhzgurKJmZJwhe1dHtVOCPKzMbggofzGyHGFVCg
vZxaW0cHloDj6aTZlcDVv4su20FscuLKY8XSM8NZNzYcmMSI5GVySfbKpdhkJoLe
UDSejhAElIQHcmuc3gQBnIplORJCaQL/TlRj42cA9HpAtjMbSmkANhcYRH/Jz4gU
1tI83vHFI6vqxn7zgiWzgAT2i4WIM+UnLgGjHeF0Vk6Sg/Ol4fZAmqWW/mI9jEk0
pIKlJhOYXVvhMRAOEuvTKfWbq+BrbjlJEXIwh2dRnx/oIB59wWqwOIYM/jhfq9Mk
fFRr7WDVgYyVX/rCYnLjuab/oezJQUTDRH2AHlm/Nu/1I2k2hUMtPhrwN5fRoPD+
Eqn4LsSJ2/r2IGUqbUyrv7qArdFWPsMcC19HxdoKYQ4idJLm/XtHELEIZuTIq4vw
XO+D+p82W3pDkWtcLvvNwbD93J01m4MxGWp81GyZd6UffXBHlNu3r/eMqLRD+WBZ
JNK0Hx/IaQW8B9CW35b7a+RsvtwCN9j58YCLTHCs9RXJbMc1UiTl934dt0bRnuaF
x0QwU/fotGsTr36vK87eFqt/V6PjfMr49xmlwIPiacuASA3KaPOkOMXab84kGGvl
eMSgA6z/rj4YKpXPv8MOseCFQH+zEuKXwVyEz9Fy9HbZDJrwQ9zUfSqn3WtFowPU
1fuIyfdLvPVvrB7CIrNta9DzhKtCd2hxyLxYMXCTLHyKcpUOLf2wZwL0Qha2WQWG
rEZ/znJUfrCOoreYtHc3l664Av/nYCN2jYwLMNBWi5QPgHeQpML3sEjPRBYEmfbh
mSf3TgV6sDIKYUfOpmTQhqCYNDj3s1m8FK6U6c3vnf0orBCzDtOxYRLhFIp3pxyG
rekRigdfejSYdDebvFVgq7f8RanuLBTEx2YQAbWKSjpAk8cKPq+iDHmC8kqNq36Y
kUR9WFEQhVa/ogevyMc5va98anzgi6X1DvkVRfGzszK9s8Hc9p2rl4NNwj5QSSBc
YMhgaUhhOBCAAvdYwCRuRnMvUaxfU1avMR5uU+AmM0eS5aeIvFFK2EpvHPbdqGhp
x2PNHBkkAgpJteBv56XI8rhxjlq4g+ZyPcjsOIvKChKjvBo4Yi6pPOxTgT09XaUj
JkTOq6qsUHA5Suzfv5Z+7MN3g32FwTjNZwOByuzy42c3EvVS7kCKJmOVV/BdlxuN
S27AtLFGl2oqOtxhNtw1+JYjGOYvZ/mRENPDwWQm4YHr2nFcchDylr/CkW6E/BdV
gr7e4S6f940hm9pWikVHa7++Iion+rRnafxe09HpmP0JMsrbDVXgS0JqoRhW9tZl
l190jUyO1VjFzCz7Qa0j7/qsaVcysyZzgej75jDjOgA4+EurAGDKanQ9Arx7i4RA
F/9ZLn0oNV8xguFCIbB/5r7TYZix83yNSb2avjrC+p9EiIc99whx50zz1S+jijyk
AhkYYxnbyM9PJBiL3US/kYSEuhjaJZEgYceJHst6hGv7Q3nkHIyxtOA/8+wE3+m3
IsAznX3jvjrtKkKHv7PAZfDpBRXV+jqMjiou0vQSBcHsMyoMSWrtMLAMhUDNLhB2
ERpv/BPUa6q3QMj4w5lu6hAU7GmO/KmhF8LgMi8iIAhgFwAa9Xh8972aPUjwaml/
3al2K1g8VK0ifOKEWFy0Z3T4DIyNwc0Leg99v0PbPqg5QJ0w5gvg022SU7kb03cD
iZu/SJch1Jcq3hFPyfWBHGemX5O7+LC80D4dTqMtCT3LCg6JeZvheATzuPR1MMjN
bp8zB4caJcWXDE/k/xgx5aab/y90q7cz64YK46x+haNTaFl7fqyLhVV4FeoBVOu3
GAlbcYzm+hv2v5w0hYqmzDmzP2kvfFzsyjiRHVVW1tUX/QFq/lEP2gFH6Nt+82Y0
Dv13JWPVwM/IH44unV8MBG5+vz/ID0U8k+YZL0gvT5vu6SYaZEh9EDs9ReClSbhU
jZ7C59mkgH7ZeJh9EelzUmt6bNOiV9ruubV9uGxSJQuLJ3MzeXi27mhF2PpoGk9G
i8dGYIDsrqJxraj1l8I6YdUk93KcVMUQ8BnTWmdXMJqUlQ2UFlKwV6uXMN7Ddz1p
uEkb+QRJwMg8Gl7BurkzRrl/bAtZliSV3nojNbtTHDPZs9hgTIevbeXeaEyMctU7
4KyZ+P/QwUTqNGj5BLJltwFlJiJ28/ucrLgCkZXByCVbLxCtP9WepZJylN3nWfpW
dofFGGeoeGmJ0SxPx9thPZNyCsMiW5BoM3eZK1QYfssV9XRRXNAmDDqaqSbnEw7e
mcSZ8nSi2lFccEWQJ5iHf22iZq0+i5oI8Me3qPUCY/jIkOd+Ks9G6n6MhEsxESU+
Bk1hr5xekkJYN6z1t56m6MfZCevCWmB98VacoFWes4sYZMbn3ghwwnI0mTDS5XSf
OEdQzSfYxqJjo18KGA4F7e0VSVJAqtO7dl7fSePZn3HR0qB8SUPhVUV0UCzo+QcN
UzltMCzDwldd5PmCARrOvypQWKD3H8dbJjvmY529DTG/2Kpe6sUuNE5P323tPm03
MDXgOyV+bAUXjN/Qtp/VzYenAUz5bpp42SYAq3AtVyWW2JYuD3wJ9Qjf3u+HvoLm
67Ufkb5kYoylUU5dP5KTAdlLP5pxqbww5ZAHo9uUrNOOv8/ecU7s/tAbBHheiM9g
gAwvtdrqKemKYzluHJ8AI7SxatIlwTlvccnBbPd8TDRMuVpoulyWEujjtI6W77Ip
aXtpO1xbvcsZAJgcdETvV5JzrsBwQ9Uw2/Vkn687qsxOag3LWMjZ8famt/ZQk0KD
aG8mQI/jpiIbMJP0s+ceknjq5oy6B0Btd9jsX42Pkf4ZB/kqpP6ZIpEU5IPqOshV
WckWhQaa8hhoJ/d3ADqFqgYQKiF/BuvbEWCOyyJo0+jCzQNUYdPkkl3Z9Qu/Y/d1
s2COHOpq5UuRqvHaMMeHRTVvdtPHTQTCTclfRuAbRtO0IUEvd1KGtj81ivCMrEuG
Ur8/JJOCpQoAM20vgZE3rX3L2NAvdAEIKrxrHuBMDcvb4VhdV2GTpIGgU7udH9xr
lh7D/hQucJwqNWxBEqqP+b0JJJ1g9RAoy6ML91GI3h/W+EEYfQrv2wUng1traxoP
t13a5uh5n/+4r4Yx88lxgqbtmbwf0bMAWApuYwr12sC0uEdU8G01Tpuudb5Adrd/
G50rgeX9iYiQpIzj6/IViuAx2zTemNW5r6PtQVuOoeRsQ1OQYUgT7T/T57VarbxF
y6dAqZ6eB8NDKgLx3u4tXH8tzcwNa3UaRMWht9fwzc0U6oTIg0Fuom3QuGg9q8Jb
ASfkI8+RJpvNq1XxRK5Ie1YPGweRxsxuAm3MXhnkNOvMsIs+4jhUC7udtbom8fwE
5DfIAouUo9XL//u72DCg5l+Vrk8DM4PQAtWFqZJMSfQMlTrjYz8Sjslz28qOCo2P
LaBp6VTOPUR3RdOodXoykw4A984TBDPd3zF+BpEf0nXQvZVHLVnY45UKj87y0Sst
/Zt1pq4JnkwTgZW/0uH+NC/y5dYacfAW2Fj3f1zHchqMGLKIkQVFmrgo9C3qdaUU
yWS2RhZBtKDvKDvl7h8aFJAojG8onNV7YIPW6lH1XH42nHmt7htDggiMkN//00eP
zilK8ZiknC0Hs1AUW/Cl4+bPRl2oixbdp6WeTJ88ASfuavNtNungNFMIxEiDDxjF
8+AKziwW6+iAvEIPx3mzpmxuwfIGbxLQ3/bOfprkI/ncIdo0ZrvCeSykJhm0C7r5
GsQAQ5v1lXkpbOZirWpnqo1JVOKnDIpp75sEtuuu3yUhQCRm4IdOSpRnim+Fie0Z
HA0a42go8EtKpkQEzZQ2J8h//36W4iBxT64f9oak1u0qoFXHo3dSeBS3qpoA3jvg
kat3812iLnu/aoMpTocoC6v+O9K3dR/GQCR6KWVf97lmouaTwGQHkhWc+OU+aVtV
ClV5aCG5oKyxkYg09+MKwiwTbQr/yi+GMm55WV474Q3UBxzjE/+N7AIZnwBFf0oL
jnMC/+OHOMOELpvQUSyNH93m4533eDxbMdi7xUTw+8IZ264/DS8q6cWkOIENjd42
tDsj6ZtX+xpSVcheiRC0CjwYfVnRdMeueSv6Drtu283wTLJZihpUXwdKjQoYARn4
+mtVvudVq7y2oQabnS5TFs5rUe2EX1dlBKbl4Dj3tW3mSd72Fxv2yG9ysW4xPLUm
J54Gjn3WMR7UV8YF9GbODUb45Wcir7Nqo67H9mubuzAhURwUAlaE6NETpWtTgd9W
LndnVQOYIeoHSFXQWzUcih+e2cCfdrDrnwFR+y+UFIbwkjd2stE9r3u3UEs8BtUO
9EirgnQ21hQTua59SIKayDjgESgs5vi84J6ijikDk1qT9CjRmJfBGZsrl2BP7IDb
Iyl7dxQvlXZK6zBMCrR52IgXZMWnbwHwXEMlD0famvg/iklKZaiNoA7k3QEnjdfM
/byRlSRtQ0mIWiB41DZ3qcB3fyKqmJHrJWRcn50b5wxBz5anE/1ufyhiafbtXyB2
wllG/5B8d+xYPdnV1veFGVGl5nGLEGp79k8shxCtkciXZUmmUzO7a066JZY5t3uF
J/bOkxXCUz5qbUh2VogQ4riLZccSeEQ1kvYpHm46A2zilmZGDVJvisVGk8AeHOEE
Q5cLTdMR5aEg25cA1WeTenMiX8ZfiYDpCIcxpBT0v8UVzZ82ratWTrLRoirBaUI8
IyP6Di7cdgGP+DK4xTjCOYEGphnDg0b+6uOeJ17AimyCxSSsT6Xf+QYCNZynrU/c
jfWIcpQbNPvOIhjKjNmt7JII6BwzJAV9nBegvBFF/NtJUx8YVHlGFVGWno3zAp6E
V97w+PI7A7JpBnKaSZwt0Wd6Znz8sL4tFlU/AeKgHkNQ7/D9MN4T1mcNYwYJkdXl
XSTKRqDoypPF/v7TvcwyMIjxbAenqRefs15rqj7ksZ9CWelZXGlsf39JoZlqXFzX
w2huwJQY6oUaVvyIxeAesk3qn8VDLrVn+XQ/JgBXH35pKplTbz12hV3KCqF3JQEb
qs8U/ZipKqFcebmkCvl94IaNrTe44yLyxroPNB2hJeLxEh+oAq/R2Y2ITsleF98o
Gwy2wm0+ksfAbvBiRbQ6EgaoT7BVRCC0+HFGBqN4bs/E1Wp5eblB0SAYjOLYJB3W
K+lhGkYSNR6Fal9ZKM7gZKFgKvLX4d1X8bOthuvp/hzgruO76jMYBAABNi/K/z9C
pHzwky6Vu9Czk6HpyqWfxRNXQ8N30DHRtHzxyxDzIa3RL2IH7SaVPnp3oijjyRGK
U8LV4AfVs3S+DbcMQ1/kv7AQE0cOP6q2w6bTTrhdbuWjMu7VyjYpjMAwoG8Dj2QT
jKwU+u0oD103kHfzM8h0HpJRHrxJ7KXOpc0xj1jRqhPt4G5InZJH9Kk5tF+0xbmN
YTPn+2q5SNxJO/VKIdR0lnRDtlytyEZYdCcRyhCPETv00pgIrNJrZ0NLpentupV/
Fnbhd4sOmPSBW+sOyDwTCKjsi7ELQXZaNCUFsJh2itnH+DtMDGPokIyc3Tqp2M1+
X4OIGwagVA7YEg7f7Qfh926TviyQymzwckHHh6dnfMNAt0asxFFhzdPxnNMfpLQp
1GSxTx1RNz70113kPbH5bnAMxKrYW8LNG6lMA2dXIYqx4kd3RAyygt9xRfeiRUXo
riSvwGYCHEv0iWPzVgp7eQubzK1evKcj98OG7sKF1IAJQx0YQSJWeuN0mkaXVsWL
EnYZmWLYz3tc4oPiRZvrE5XM1R3Qn/CSNpBU8cl91+Di5l0S/ICvY/gVZqLDnVNC
1kUTe4UndKZ+QAMLxPF8zCHzEci1TqLVsMXjwxA/JiyXTKrRS+C53qVahQ33UxM0
aOdCuu0TbvTiLCCYFdD9kM0zOpdOBPH5kcFutmGCrwbUCiDABrZGf2ip+B4PrVOu
aMb25E3LckjIIyOx3ZORnjpPQ/BZm0dmoXJ+zmhaSNlsA8oyGlnEsYYQIIQMDeit
8VLyZjoOG6lSkgelw5GNTGCszhOTxD/VF9YJunc6g9xh9mulTROdeh1S2XNZacZE
xEtf0+FyOuSowNF6wJuFFo7WTcpvfJ2EFotz0HR+TvqSUeQ8T1eYCXZlTaVKEVoj
Qg8WeZj42W3mt3R3WkTCry3rFVvpjqB5JRuUpEL228ekfx3GzRL/vJ40miRV9ykJ
fL38BxARHOzemnsecy/EhJFY6Q7gpd0hZVFN7amtkDgjhjQ28G/a3odd4RXwt8EO
3XIXcIuuN06JDZlZ2kPEsmBy5Bpog6NncbtVRP7pknNHMzZw3siAMZNSVDlMyh3J
IcbrYuE+Xmr67Bui9RWlxH4JDRnMyFpFb1YVRDtbF6pE/SccLQyhvy/w2pzQi/3y
dteTmJPI5Xxb12ZyO36FF1WShyhhe4M+fkL0V6ckzwLadrUQ0WUtGX3AL0sgjoXl
u0vE8KdQ0X8y/C64yyec6KwPDbIARIJkVeU1Ru7rwCq3EpCYuFYm58o5mnEtSoBN
XfvQwrMm9e33pdr9HV+N0MkbJ9SovI+N2CMuJrWl64Wpo+mtPYdOEueCfwsaRogF
X55YNncMepQEmG+UFSGN9QYVDJBK6wqcWSQbrff5r6sGFbXiwaGddMLHRV56xny/
xYiV7w10NMEcLQtU5EL4SvlyEofn0mkhdk/ORsebcMM9pIytgtIA4LYirFtk+vG+
L8JVHAnOEuZnLWu4u8p8msTKZrus0cx+WpKPBfKP417ECuYq+pr4npdnQmO/R9hx
Tsk3wRkc8nLwxSt1hjxPxPOITGPCN2DJNfmRkn4WIzfSHMZE/5fu9mCD9/Q/B1M/
YA+OLAciOinUCjwgzwqa2yOER72n61jjBmxdp7jw+6UNZ9gtuf9nq2iOkRkI3gor
J3cbfdx709dGR4A9LnJJwY7QaJEx1WG6DSFQQiT4NB58Zgih23/0TEf55RLs2Svm
ARIdg2HqXAtnp+fdNwHuc3HQIYajmGAUvxdltv+pM7RPYMiTkCbqo2T/YW45X0ub
4BtS09U2CDPTvYSIbNJquilhYkAKBSByyhEQlgArCPMG9b6OGmGjLEvgXuFxEDJn
htHo7ITkOjNtXGWblklsS3uDisotvqt4PvDE5Tr4HIeRucA9VQD9FRqkgJL4cPci
8DLjJXHZtnhWZLkS6d7nuJP2iRIYFXRUae3O9ld0sxLRPLkqlVQ5neqldsASCHca
2KRArMpE/zzAQg/VJOCbGxC0YbArMz741e4wBFKYXk/dfzWmrBET80jF5dIh7n73
YESu8NUobSJUc7lCxYE3X1Elfyw1J35W8qrhbdoUQerwsPcapPWK/PaoEeL/MF6Q
C9L6Yr5ImVLXA7loK181H12nbzPcoTqagSOHXXPuvilYbEI6HmyfQOYXvdoPzYtv
YsRTlUuYj8WEeTEjD5pGS2Mdh4+jU57r6WBcm5AcakJM54JdNvz4xTS+PyJIs/pS
piGVpe3TPKIdd499aVuElBQuIy+4rEuxOcLmhJ5IJz5WxPHQDOykxpE5C6mtgnRk
OXYql5YbwvOhzyNjz69sx+RVdaTLxz6AveJNBxAKB1fB5ZFoEx+MmPdT9e9IrEIl
wC50EA59tm7UKGD28o/McGZ6ievmeHh8HVeZ0F5Ron1DPPMpHwHWXZwOakfg9C1j
tEnNhNv+V0JvB+21EWmFUNFJ+pziFnCfRUuK8KsL/SDCnIuUb1sjl0QmIPVHncEg
jaoqEbIGcKt9OfhnWgKgYAX5iys8lxQP+CzfB2WOC+lXnNV1dO89TdE2NKWufjUY
V338y0yGxjziBTeb72sS7uq1H8v+a6gxnauKeBp3MEVvHFHRnghTjqAn0xKQOOEv
cfqF84X3SExanvqLMO0rsDQEmLnKZRXK+hhqVu4jIEhO20pfaLS3Z/swN2Nut7sK
bYHHLlr9R+41CxyRjeTxp+YY7+F5RMdClC7LodbIGfJ+0J6jytJOLrqRQV6PXfzB
HrFAfkHBVRyCZHhYcrbVarRde6GscmPztMQ9wfh2ZazfzcfmujDhPGzYWvWNcqVa
KABLtRbcc9ozG6JnC3XJODoGMNPzUi9cOMIqxf8yitskvb+59VNXPUbxvy+ila/e
zb0g5NIFd/DrlqJCO9D4w7XHOAbZTyBuHkt2k+e6qJ9b51GUo7Q2lSl4gF5sBr7w
96MGvhJHMxONzdVDj986veSsIZQYP1Edq0xibExZaOadXbe+MJxJQtIH67dfFFYy
tkkDpVfcTqHjPor3SvE1dZDptzbfgL/El0Wq8JiXYnEcpik8C3Gzo6BFRV9JwMOJ
XDyGMcX5S8rXeJrzo1SFw1PgOGJFwCF5K9VbnexAlt07CiHQop+v9/3ZWScHXII7
zK23TsJhp8RmwIQtrjnxQ3dBDJ0qUmTNRNnaA9bQKKkXkriI1DiCVdfNNSIfS92w
RUqeu3gmrkAkIpqF6UXJEUpRRX3w9+LbsjKacORBpz/NvMRfKK4t6Tm6d55L4D8V
aQrATCOsWWbPIewTswc42PCHklOHOQnwgw+EVRGRNtLpe4mbhK34OsJEOSxVYyz9
PRSy9dBMx5iPcZeo30Lxi2y3462mey2vNNAqtPweZLEsTF8DxvoAvvxMAyrM2SjS
20nJAiEWrAtk34rrwmcs2noQTWVMP60JSagE9dqHoelW5zWQx03bYRpB4PAYT62K
AFCgHXE5FBdBY71B2CftawVOyz0F2Jme3MXW9q1DU1VVfpZJAikJHkDRJmL4nXjZ
G6cQqLWmkDve0QKH5iXMl9pijrvwRBDj5/d3wZP3Uf5IaXzEBhfCid60ZP6olI+e
k7CscqP071Hewn9OUIktQKPR5OKgxFWB7fP4hVG2fnIsb+Bstqk7+f9AbyhHJPC9
dj5U482LRrtY4OLZmnJGkj1OvBRVhGVDzqH6qVjsTgW6WJHNBFEB2sfpFPPKZBK+
Mxpc+2HgOw7j8BPAjGiv11mi9xKBfsU2MrKsNgsEmyR5MFRlcb4UewjCf6fl1nNS
B4su/7NyfpmR5qt0jsZKPIqHdGMbLzS4ofmEiaIeFElPdZ1mSUw8pT927Az5q+hv
u9IY4rlRBjCEtl6lNoFv5hAQue2WU82iZTaYYCufrKI3ZxsoT5c6Jc2J+GfnUORB
2QXZepWjeqCXSrPr+e6KBKjpiCZU4p8xfEenh+bi3/cdj8cmtzCJeKVsX1dYpWCL
2ZGd2ac38uNouiCq/yp69u9xh/QjAUzAcXP4mhXed5p/Y5YaZR7p0Vi6YF+NffZG
jPVfu+4SxYJXlfsjbg4qDpdLLiOTnYDY3Mh0GXf7Gvoq6RsGRxuIdwsMnQm4GKbT
mJriIHvcIa+kkM9VBzQQ6WFrlWnAH8QCEaRWiRGMk085PNeHhLa6zkT5H4ShFD43
ODEOOCnCYkfIJ7rW9hcuNxFLGitGckmbk0W+bMo7xnqb0GUl0fFSIMh/RCFbd3U1
vlxE4hXv2xr7ZMegXprzvFrHAfIg4JceBs3yhvHGJK+8ydCAKjgBtm2W5tCCLBlp
zs8BAZTNkHH0jYEDvVyglejN59ZEVCjLkh0X0q8iU9WBxcf3AYWJwBdn7jmFuY1Y
GCcCDDwAQBsGENq6kO9hqcqauI7Vi7tBdJagcdfCFsfO38baZiSb7T67sEbtuwpz
N12iAfQuRVM11+7pb2lnB2ciZ0Kt4uwgDFBMaIow+r2GAlfScn8wLR61Dbwa41hU
MFHfZkhZwSfYvxN1Pgp1m7l5H8E+j1dM33W3zefY2VGc3WKEz3qDmxvJy+DiCSX8
/UY82W4/C8zTptIJx27b8yXtLx4h6HrsFfe9aB/82UAy12dqbDN6zFa7n0WDLSoU
6CbQNWwQxhPRK3CdjrjfB4vdrHTaGWuLs79igY9CpXMOLtGcQ5om+nq+JGLGWJ7q
ZwrshgHsMp9ixkSpKMUJnhMJOA1OyKaTv/UxwS9PbHE90GgC3iqj8DbxwbxClWIv
6Pne56aPc6WRLZBK8bTdm3RAZTHKp6VbC5J0NwkUf8k6gCB/hQeV5wT8Fx4YsuSL
lNexF/vx5Tttyb8F70fsiS12Lyuly8lP5Pnl3A+GB7wdk6ovVs6p2sg5YxB4GeZg
lixyPH7XaNGyVjX7rxoa0zv/ftuvtAu1t7Xz16b12YJAZiJCCpmJGU8ZLE/NMMUD
SjV4rfh261iaHLsATyH9/7tcVdEEI+IZVZKV2NIqfDnrH6bWzPaP+UEe44R5jPO3
pmQmX3BVOh1LHN1pbtdjrkFHys4rMTpffNdYH7x7Fv6p0KsZ0ZGQuV8DfF9lW7Be
YPsS9TxYq33LFh1aYPQXHysVS54jk36W3B/cJdOi3qiqGjdNKaco7ZzM6VGyA5HO
iVYGD6xexAvzRplFROTy3RwuEo1L18Q8yc97+yGv5yEd3JhMOJ2KCXAD3vyDXCE6
Kwl4pcngzP+CPsLIhaWGL/+jXt5WO0r0CfZ7xAJaheWaK8p4CMAWVKT6pNrJSbdq
TV+z+ih7VdBr6tBOJrCgvxN84jB/6ZEwpNohJWnZRVl77JVGEqaTFHxl8hGjpsh5
oac2LKyK++vk5UYeHtFWfakAogJ0OhQl1tlC5Xgroc5thJsLCzYhXlu6OkwW0jnS
ZuY/PFOoYIM98zt02IusQpD0ubJXhg68HaHpL50x7rzvwCp4ch+QXMQ3f+b//iuN
k8FAmQHxNGDkk9xPyDJPp+jmYOgSGKgdZNKVLDHtcRjSq4NjMhhUJASNC83qjiCx
SqnpCXds8uFLgHwtLS4PA6zQbIlpZi+BdDKSV7Q7APmaO2bxxDXnXVxR2Ne/uAFT
aojr1ncrfVgd2Ad6A1HB6Sz7Mn0KreAN6WIrYzHvu0RZvPw/JwFlwlgIz+UmhRv8
MmADgBEeyqPfBlVnZOBcfyjUrnfzyoe/Z/J7CYF/hqolZCuXyamR5rnLneMINEwv
nUJQYco4IamH9Rjmo9OAZ2fbZId1zirjB9W++04LUV9D5V1RM+0wpciukQFT7MI/
UDZNF4GGY6B4JJ1teVRF9ELuOIQtoaNbsYZjOom9xZzfu8obrkZ6pu959YO9nEL5
a1h6qAmleCV/ANp9JxBDW0ZiyNbgPEvdz7pylEKbUtFjjahVRwd9licD27OnMgWb
TX8Hkb+dfV2nWz3TSzyC9vroybdaaXRikqPQKMOnCMsmx88EAVL5h9QlH/qbtrKc
fjf+qKU0HvLC6zCRYvFVViRFdJM2vBJ3MKKnJ39Axxz8NytnVPrrVcRaNS9wBeSx
bPqEOEZS+26EKvgr6Xa8eHp7E3+NV2aO6gUuWz+JNRy9Yy3homNdtkCaKshZ5V6l
0DwsghlyrfZTBCoe8zpZnrluw6J4KgotC9DEXBPfCS1U9o4QUfWtRtTKeoZqXdkd
80usANoQuXznWU//OvZbficBQA6WV5Pt+BZikk/EsPEVrLcywDihYuM7BSwENxCy
VoS2AaV2p7R+2GvHjDTDBEVkAY+XhL92XAio6mrhvLz4BaxPQAwQUBgfE8J5lsOg
25jPUcQZHCL+SQQlXjG8xGCjNtvaIIxzKjNVH9ogzeVGFgZFy3gUsd4i7uI415k/
TnoL1vvr9nRaBDOdzSEOTT5/NOgESZKZI9NcWafhYJOkmoOy4VfBtQPg0hlfT3dR
WlvoxFaBT+JRo+OI2h0Rp25b3f8NDpTlDZk1W3Rqrx1Kjxq5VxQPcz0xHZ0iF3zL
dt8ng+1L3Z0J+kdNwqzVQFk2L+mii+QhGEHz6OUAsEH5w3EBkeSQup9PCEJcxnq6
XUQej4wpQahAkJeKnF4p8khzOlmb9/tSxPIIh6SE/giOZNdLV0E8nWAEcPygP6XP
l9XEpDV0Gs8CSbf2rfpqR8xpTmtW0LEgLPOEgu4gc8qq3aZwJhcPLdr64VEyjY5p
L93FMcC/7dDABRAiJYZQkPDDRZjqhfSaqEDQQUI2lmql7RTPB6Iw0zYu1YGXTxY9
+o1ORzp9itnQfh3UTND55hKow8TaUwQ+ZpL0vxNsYhi+PBOm7DS+xgWd9OacUnog
Rag2BIIpUODfWL+Yzi2liYp6L8C92XO2j2uvEVUJoB9josuVJs/lTMLiKbrA4/7C
vJB5J0uzOKlMo1tLH3ygTSLy6qXEVBV8YGWl7xbiJz6i3AUYFbvIhyrTDCe9Vsi+
a1Q3O4tcKEEt9R6Fjq9ETkPHYdy9q0vxmVaGxF8N4Y/gZAfOoqoPrHDs4Yu2Xv80
9fu2IQgXqtW0HIOi+cT/rIK4wDyxVDv9c22Ndeu5mRLGSJXDC9x6ql5sNZyxJu1H
IYCQxRjhGjj6NGGRg47FitexU9tFE9Dq2Xx0jglUFeL8ryVrx2bEpSFczTfbeSHp
PMyakgJCxBH/KRbCO0H7Ld3zyY21gdZmsbjxJjpnCp7/Nl8xa/3BgReJ6PO4n9HB
GzLm9+1qv6yJK9U+x2X5Mpy1N3tnCkMN48gGz23GO//J6AZnpKWivnHR6cim6DX2
qo3WAelv/JLkXjtriIFOncMYT8XME4FfYRlFu4aJiTYSiYbNP2JWf6EbhrWPwc8h
2SN8KG4X3xUynrpfO/v4rDEF8htjuTkmbIFHo0BALE57dYpOQifqOTZD9qQTB8Og
zZ7jbTFkwY3Ms6sEyZnrFMWDe5hqytstTOFImzI8n11anx+bb9FBqcopoJVDELiZ
OlFM8aLoYN2E1NoEc7uaAOslllT05QHjNQywsbR3I382Hb+yIhW0uxI65pUvoCpX
ok6wb/0lOlr78t2z9XVddHUXYoenCShchNayFs5sFekSmOu10APvdiUTsFsagmFv
tJgyKCZUcvOFebTOlGt3lh5qj/GHANmhL8bIh048OhkH+pBqUkcYL/UV9YPECXhp
9EMs3P4+1RjnhE1lu7wzWX1JFYe8HNS3VIqeYzjJbmRZW4yamUnVzy6zB86QRuny
9Rnju7ZPFv8Lo+gOUcEwZ2PT78Qzxzg+cUMBLJ7n19ZaOH/YrC4NHFkv305j35HO
2fb7zGIyyIDSUvnXlokZioq8zoOgoYztOJv6hCB1YEMR88xbWMSxtfAYVvWeVd3h
B9oXlk6MouMKrt65yA3nfJIFmRm9snhiFnEmyv6ODU+EiXeDlq8UHcsJnT1WErII
yQr5fjlxu0qQeKk9Hlh81tii9Nl1Z2UkqPp8qKJ4O09VaBTqyuzKoNahAN/ywiKa
GVRoXVmN0HFhjJ95T2tzwjbpcQm/aqhTewPS6X3DkMqhqBLQkQK9czCF8IgIGBty
UQw2VHZgfNav2JRgoTp7rqzzW9iE3hHOQG+kLtDpcn04Cw8RnRWQ4R/78Xo7kZMs
f6yeDBIf8Oyn74kalYrZgNp8Q8LnQ9coXU3sLaupZ6B3Y4Vpboz62invzgigpBXE
meq4UKr+3ZNBTsM18FTZrywo0KpUfrrRsiL8lrcipry1GP1LF2uFokFWaUfraI3/
Jd3/fCIqvRCuOqPxY5vrNs50CxjIFmNqRMXvm7/RRNp+mViRoKKjT3roD1zGW3N2
dWByVrXqrGFDWtX9SjQYJFWtk+AdEYBayiQaGtUmk82WcVCQq+OPt76ACTKz2DdO
1JHrj4ZtSwnKtdIujlvqDHEEcPBk1sFTXSdgoHwHAkQjKRFMeGL8KRNExElDVB+j
dsZfaeN3yFCXkqCn3XUJL2vriZLaiUDeKCZZ5F+29NYmRuqdcw3mcMS1grd2lNWq
Vc36NdJSzy7Rsi7pfFTA298GNqufofKZQ4SBtfgfDrePzpBhwJ0VhLL4jR3F3RcY
E2GSXiFoBdXl7oGNPPF6KkxlWSUQq2I9Bqie/uJP49oBADYP1Skl9NITKoduZ13H
pjh/qrJkiYKUzUiEwWnRFk6aNDR3nXR7+FivJZf9+DHEmL2IzSRFFkqh9L2D4YGn
SX8I5t7ks8S+sWCKCjsC++KdOldvBimp278jIFEscwtNp+7n80qNmp8KcjttNv5a
8QWt3Zlp4LqfNlBTLwcW76PX78XwMK03i9np1OvLubEG63Q2qXfkWPFcG0X2HBJ9
wljM5gp3SKRnhZgTMv7ywkHJE9eEswIqBjsVXYozEKIo1/RxP707V/D6YuCJ97Kk
WEEcWTDi3gxHjYyfRAtmtxIfEDJeM1xwDkubW5g/UUzHUh0KDt8w+Z0iQnpRXOtp
yxvgD1Hl7Nx8PuNtlJzaePI5QqcNaoVEscx+LyKQhORgriH6tFItupYrkKIMMjC4
ms+qnvosXLMI3lmLmOBLTR9yyZkDGRYL6geUH2uf3wl79iSV8eAOSoV7NORo4/+w
ZBp1vY08s2LpTKDPV/Qb2tZMMeaVW42w/UkbSLYRaOYCzUggi5aqUjwkFbvSM8Jx
Dg+mXWg4M7eQgECg+f+5o3z7PTigaPyJDRJ2gSm7yBwDSfdH4KfjWOM0xGW7S8En
OZJmxGMlwfASNHbj5+LnWKV/k9bIJQM5YXb2J+r1NI9MG+cXtRK8+4zUC28qzS2X
3Wj8o+ZzNmpV5TMB/65z3cDuTyHBhUPPY+DEKxpweMR+T5RIYFwEZ/SOI3+x0u+5
pU3XWi168Zpo84ynbPQXhK3VFDXGCg+aBRFyRcUh5EjtCM8tGSOUxzXTyZUeb00+
rAMiIgXg0u+LJGYSF/9etCBuXnEQSHvyGiGMOzNPnKpV0nJ6/ekYOLwkrDY8Q/Cz
+tG/M4I66SZ88AoB7xHQPa/VulBKYfqHKe2c6IQbxG0xdnmMICh1NtqwFJhk6mPB
Qp5md3GM2D5Ixj2NWPy1ywYLmrE65q68WnzvXJ8lN6pRDS3j8H1w2o/L4BggulB4
ijqQq1AdhHFcqIwOW4SnYZrIeB8LPZoc46YkTe18p+V78EclhmbN3Q18XIzGkNu7
WzAA8bcAddsyA5wpmveBp9gqxkxWHZit9MmPtB9QSBvgEEpOkJOYetutZc39Fk/O
W55+gtQhBRdjl7Dez8i/QQwyZYJh021yKjl/fFy4ZCThVRpKWAz8gbinaZ55sfv6
sgd/6ZrXkgr2o8HNg69sFO0owKRS4dub9sA0Kw9/PHlTvZui3n0RKY9m9LMad7Z+
Y9hVy5LLSythWfUhgSV1+r1OCQf4wqYBy76fyJAjNuYNTm+KsQZsOZWFqFXCaG0c
HfWke0iKWZUYszmlWaUeOKWtga5ir2YPUx6bi0ZrRRJL7phz2omKEOO+hOhEZo3y
633upJIG+nGdca2w4ttY2SdevMBAOKVjT1kKun6IEjCQ6R4HeJVsS1ZXtcpK54BA
nZhjWrpD91/EeQWlC4v7mmpA/EGGvRCEDQkgBz1G2qSJEWWJqxxkjSuAoOCwmJeP
ahWAMm8weAvuDmeDrPRPynDKP9m+n284kNlG8vV0Zr4H9E9s5SQNQASTkEcMLf1R
XerMcONlKsZI7en8F6RFTmKR2AdMb86INN17y7AePBoi3eyNCjJR9nzqJeeCD1Yw
/e5brhuSngKeCa7twSAHqKgB9Ltz9uNBTcB/jRvnHRCuveigYZ/OdkSKtyWgc36J
nxbTdO5sxVlnyIt03pgCtss+hJYNaxWiyKp+dipcoGN2WBoNtWp6VJGGy7hmGUwn
OalZyBHLJIHjaXUA/UGuCJ5fzSu299z8+83UM665m8dOw0DPGSh8+ly2XuZBSk+l
i6GcwBEgBVW3RMo+OPaUWcfLmzSolef0i671nd2hR6y2lnW+RMwNIWWu+NVyYLFW
NQ9VOpYKKIRSSkS3ProQ/GMj5Hdrtgc3mQFL1JoAKrNQ6FzYd3d17QWQrKrwuWiZ
ZhQAgwrk0AiHDlaa55gDeJOsqi+egxaDg6faNkxMhYCmMmIKjPbVRyEzXgCIFBPN
fFI8MO+Uf/EEJ5qg8AtqHD5awjN1nW5u1WM7Vu8VgDDwxoOkgjNfBsyhaPxOUGfu
/reaRZ27DrwQa/YEbIJGau69PXYO965Di41+hnSrnWw9wMoNEJWPNZ7qhdwNIEf0
NkQ7rSXLiOtL3t9ewiN5tO5/iA1r6QD2JZv+PfTbj89mVYjmz3lJj9lPEC4su2Ka
v5I5HGdTs2E1vrSMujwE4BmDVPF1cwk67pWdMOwvKXDVJdWsqy2kvci+pKb+DR6G
Jyb87KjJ+drCRlGdmbKa4YqNQt/zrL0jyHwYCOMVnynCYuKulJOHyXvuFJRzT3R9
Yvq1VsU1HbwKJBFgM6vKSLqwvcSPeDYmANSWmCSxvWieYMg3EsOe+ZmJ6OZLIDc2
tV+ZCZJliRPfcXMPur0ElVpYo6/0OSzPHnYS7beKMlN+Xt8xx7fwcAMFr0WZlJTG
JxAvmLmYcw/kuwXo1rbLTimc4dQvwu+wC9Mpsw09sZKrkCxgUUreTiAyQ7KoKyP5
W8P7Di3HJOCxUMErWmvt5dF5AF2repdtR+ciP9zWFCS/8ikgqcuTPcbCpHf0K7pa
fJK75mW18CUPzDMfuGvDxG0lrAvm2IkNJJPjoVvLib1xPCcCLrowWpkC0tuuYKYX
yeFjMaHMuzGlRYTJX4kr3J29pvQtXM2jbZe1PCm0lxQrb1ODNoUyNpYccUzVN6/K
6gAopbY0v0LpfIuVesFgmfiilprivRn8l6jps63TW366YA7R9vvLOFbxfmIlbauR
Pb5l6mS/PnukRHl9ZMBY1lxfpZeTImIakshy+dDul42WVkzhDiBrXELUf9B0Lc+B
iWQaPIDTB54oh1rzrn2NktRkbLy44gsiK6J85m2Mi11LlqsuRzwU/5ZMn8f8Zb1V
XnyNBEPMPVk4pesqqK/1J1fJgxZFsgqQiRf7PMGVOCGsBAW+yaw3olzHBrwo5qOg
aq8pz0jz1fuSfenKl43LhXKHz7zd6bEn1yvt7cYRwCCbdO+Zl98H+/GPkitiGQlq
lTxmSiB9gB/gPcCyQrpX3RLkP231HymKhev+uSl7TyAWFjMHQzL1sTQ9d60m09z2
dL6aLzAXoc3kcMrSkMLQD0OHVDju/7KDNsLT1jVsgs/2UDon2PLpPNMqmgjGgoI5
vW7ZONoS1ktevS56cfmWpecDXqYkfMEBayzx76fZ1i8ntGRjGdS92H48ZKLpXXpf
wvur6TfSyxvcWTe2lK+AhNA23qICzsywuhiQ1lUqVpKI5Wy2PEnW8qDxlSxARrLe
12LFisgKY4AGabHvPpBJzXCjXMcT0y1IRLvPYxpfofJ0w6z4xHEPLLqCpSEa+H3P
tUGc3fwaNuLYW/Aho0Z5wkUY3Awvzlq9E1N22E/D4f5nH7EueIa3GmuM90hYcUNb
rnN9c4u7ZcSFnUIb4ddPEs0V9xwk4qV3f6PCpIiwLKC6nynS1xWa8904e31IhfCZ
ctvvhoxs5vq+yEvVjKAHkumYPNDGeTL48JaKuuIjD2xkWHZcjxWzRJETktNC5GsV
U1+2on9GfFtC4c7rMeiAEgFge50qJTBThQytNU/xHmDJhgP2D1XMUh2WFm761lt4
yHJpm06XU8Qv2gh56pI7GS0LWlU6AnlH15tIDeRCwXzyX+RTxruPLnQw+QTNR+Bn
/kIIiOwlSwQt08+3AA8PaLe6i9mDwRVGhx104Mx01J+wmEg1T+cMJpnQ/XK8H2YG
TK8F5fLBKQQ8zZB3nWR7GPPsEPPCM4nxdZs1m5+MFb8GiH5SEIw3GPylcbBeYNjA
PctekNmRAzJwV97YU58K6cFr6Bt8jqCO5lq6puabSyiv0f0IELfTdEgvFJpuxs9l
HbgJf1KgKfxLAZHhrR/iV7uq7R8WmGYTbrIM2uMIxqy5Qx9kSKTt3tvKIqn+f1JU
Pbgl8A/RK5VAEoO9hWzTxbQaUVI9St+bGgbPRV1gHLQP1zZNj3bJSFjz7hnU3X7L
gb+nSwQ6BVMBxC7lr+vknsexR+uPWs/TfbY2X8w/Ik7Kh9XUrmq/o1F4myiVaqJ3
8FZJwVzQUtnl8jGcUpVEGV8njka7iTYFHkILxHU4+UNgu4KWVcyBYL02VtR3Pt6v
DlJRw9r19PmqxRLLDysYNlFCRhhe7MkpLJrOKYqztKXy6a0By/6+xoXxEA72PDEo
NIXf5WSpqXnQHX0aX1w74mXSSonjGaMYzNzngcPb9zlvCSEphOvCFiS+7RSUiUcw
ZS2Sbvauvf8kC/xTvAKS9ptAW+7PbGVwPr2O1ML0p9uunv1J6Da1MCrcRGektSvW
qVqnvaSLkR68HpTWa67Qn58pVbyWnkhltcRkI8t4AqT+FdGtoXBsme8WH8vi5A+m
8SEFO1Y6z32I3agBmS6p3SgsDaMlLe/p7W9m8t13cJRJrmuM6zdaPNqri/u7cI/P
wHsa6eGHOhizMaQVN7HJr1nDCue5hQv2Ja2EE4+QNeM/DxfXXWcsBnUqhXvQV6Vc
ytclACTXk4jw/gnBIx/SgLxtNuwMvC8wYscBtRvB2/rVuuX1gqVpzi6vpEtEnI7I
QcTm5ZGc9RW/OjTNCaOTrxkIVGx7s1F2SnPIcEaDYt5oxlRmnS3I4wRm+2NQoeOa
3TuWqeUPWBwqfX/aFvJfMyDeidP1aQvVXJQMHYkFLXTxepc/T4FRojq8LuF8d/c/
QpShl1jprlojaSFEbLJzX4mIaKq2A0YBZ2jw34RknAlZus/QAzCfeViax5goeXaa
KHDoFleXv6BEKhwbNHPH/f11b6iQV2C6oGqVvFSjIVVsdZXXJl7OVYoFgZT1oUgY
ZmF4a4gZF92UWUrSLrN9vik6CI+RZ56uBfzqbwYTDZvBpuEx0kXSIUbQvAKnMST5
fg81FSI0UBxowkxctOIrEwNLbvuHT6mv/biAzGywdntzDzMNeueJjhmwXc6vDYNd
/b7ArLaH4+IKEWA6JiiCNHX0ZLnVmWL7Ha+98RZDah8t+Dkn1E8n47zhBjbX/NK9
r6QDlxGmiY38p8c9DrAlvH6jcwQ7Pu51g5Pjyu73+13TherLzC11bNNu9FW7aGQd
E9z5K6QmPrnsoslGHD+7gTObyJYXIGMdAZQshFAkQtysfSTs/mFcjp9RO9pxTecF
eSYiZXrEY9UuXze5vSA1IS9Dyqhrr+5Ix4pEYDb/cP060e86T00rb1Gqo//23IAO
lk3Jj7qbW5XT/K+hLlIHRlSH/JRnv97PgkiFTHFAleGdOrAbHK1jMCCNzlDumVVg
tRup3jmIRHtfSGTP8PZ3933q0kwFRHco8LdBSAI1X9jgzC/NnWqALYQzAtrpEUSE
iCSZ5zTND5yyFMCfa5x/QPLs47MXWCRsq0eWf55xoIsX3yV+nvuuX6Byb24M6Ygz
QoavIZURb2MPXLDqr6GTPsLj4TOCN9zaOM6jYnIKhoQDwNOJopuvbhWbgLUb0WUa
wuKqpbhZCQCE1mQDjMQK/95n9BpSUnWoJTy2IKRgWMjExocG/aLDS0EClTSUGta9
XbM+Uz15Jl2qZe2pZ9iUxdkxBfxPPzlKELr/vTBWmxfKxQhxKN4vbTQoYaxI+phD
55sjNgQ4k8AAMZ0YlP1uaotj2m4KVhVycKNTKjh2yhPfN3aWWppVw9DqmUKlZPLv
Heg6cYoNL2iWxccM0fmSZZWPh1rEwKGDDH8Uh81O094quqZbAk/lU2EeKxX9UlS9
FUc4RvClUEHbWzYOWoSi89H7yRrFvTZ+W7Un+Kv0sbRlIeuak0bPoWP8B/8rAXvR
T+oDOWBtJhlKCUpr/9FfQInYJ9yGWWdy1Ra42+ctEeXcYrEyA9oaFtlhCaCrdo12
xltMry6NCaS8YcmROU1feJvv5MPvWMNITFO8pE5xe/mhHeTnOrqAvTvWBCXZNf0J
B0vqrA0qYCkJPK4JDokSussD5oeEzIqXxdiWO5xouAPHSqpOaS8pfrikqQGIzgY6
Ta598YZ6UtWzHU6WcAT34508NmUqsVJ8LnR8lcf8+knQwzVaYELqA7gAWBKYmDX9
L0GmEZvPUaew4EZG4y32sL9UIp+6FGQ+re4jEiwcqiuH1CvldfWi5oLt7+xIg3lR
VskwpB8/iv9g/aHsAFiOqLbiWPjCG283KFAXU4hASsqcb6MeGb+N+fJzK4yxsIVM
VWno6zVv4/w+LlRP3QBD4FQLJbc+C2ZgD0hI18ITZEWjIycp7CW9nWFGOLJ6/l/n
2kBT+yGC9uYT+TOAQF04CDyAI60QAUUoNdXlqvU6DQQj8h/XfYVakY3phmsKBytt
uMFB0xr/p2+3I/Cj9J9Eluq2oYasOg7WK1XAD7J3mZS9g5sbcLk/SRSgV+FmjCVM
rRKSDZUY6AreTSEce7YMA2JZ8rmwIw2fPZmNrbDtMc3C0GxWHZXSznYYIn1tPWTy
Kxob3ZBZ/2zjhb9J7wjQWfZvaAdmZzOt0RCBpL62jt+7xiJXxPynDFen8c5ea3EV
nq0XA38ofkY2oi/jeG96OsvAJ32kbuP5UR0UoJVSyeh6DFje7Ja4enVblm5joDsv
gyJg7hlusQ948Pi60Z1Qceu2nAgQxapuO9sZTxqIxLVtJcBbwKT+RiA0KqY9A0tf
RCY25NmyGAvJyGuPaWGtUbbWS9nZz+VLGVfK0MwUpGqGy9JjgVBL4/8oIAoNTS4+
HSwmxvgSwXwOSvECNpsi3KDKxT0BU6+EMcBTwjIShmw7FMzhTaD8h+MGyk0lR8pw
VS9gTuBHjbHbmhluB324C0oNZa3UDo0Ajrblck0xh9DigjrAJ8GXwENzA/KXbByI
qkGnFxnhtRUpRB/hKsGxmLW7xY+hgNyIld4jgxFD3N58Tt3ohUHz4hAEQIpHsiRH
KfLXY85LxnoWWNzmz2YDOYkKbnDRTguIjreIhHo77T5Rxy5giDMFBwmybgpGzwDW
/N4bWYGFTiP2wW0YaWKBZCBGU0F/kiKKLrrd0ghMnPYQtmBxiVw9TPRJMqwBToRL
n/KNXDPrjFHj+xwqSMsO8eANNQUsVPk0MjN6fzr4slEItM1PveNZJYACSPTyJeYE
aQui2gSsix2Fmo1WzTCRDxOp50pMczJhWdxSC5w12tsQ1llesKl4qXEcZVvuKRHu
Ab+R+jNnOdYd+x0S5gMAOGWokdyjw24f32X3325p5g9TrtGC2q3qwkXlNhPLyIFu
yEUyF0fbSKG9K32IXOqMizfuq7A7JuEXAOiAURzDhWZAtfyrB3rnJb7Cx0WFhyxb
MxuJWY5Myf5MwsEugdPqTZTPah3Jdv6K4Wekcftv5cab7XgAR3KHbnmB/CiL47QX
+GzY+ZTza/NRtu3ZLZ5SirV9WKNigJOg6EkWUtoPKoXtKWe5fLcSp2kOdWzj03kj
RLcjVWIRA8yRWWW588Y3Y1blBP1HOrbJyZ7Xizz19KMXV8i+xlYYXQmHi+vYBuDt
5R0A+JtSs0Jzl3iNbm0ks2cMfBhSHeyA1k4jH7OAwXZjEZ4siMrdiGjODuYLdONV
WPu/QO3wpkhKKbaB6Pi9VRbdQeCNgnvrsQICqIKvLNJrK96GnaqIUkItnsG1xfDg
NgWupKm0AvUSX/5CiP+ngTFtPKKn0ZHAx2dW36i28CXJ3gTgHmrAI7+RkrkINqU+
5WTd6twjy+v+4km41mjK2T9GIG0+QOzIzAKbICDWzsrHHj92E3hphlbzbnsRZf3e
yEPeuQhSJLvEkBTvdWrBsDqw5dyxs0wqAqUMmYcnGhEPOIz94K8zbxN7OKGww1xW
Vb7Tyg5TBhEB6HrCoIq9CdqomYZxT9DHQfy4HhW0IblXaGVypxcJgBxKzgO28Mt4
C0USqm/gEZcSOipg/QJZ7gtXysbChnpy+0W0Fz2ontl3thQjS4apT8Afvs2ZyRgT
jxpBR5lsw2+aluaf0idZYGjN4DP/ir8ZON4Oav18F6zyRYAmECAS6AUo9Va+QGaj
z6oFVYb+KIO77mmTxSXNy48S5oeGur0XGg7H0kpgDkoC02n/eotWUIYa5HBG7Ca3
1vqGollEgcPw9t/IIHI7ETxIzGiuIakdg/meiYC75FD2RuT+O/08oHy4ZbjBASr2
PmUzwPJFSoKATrgHuDVi8Q3vFzr8MaHgiU0g4hyS1cJUVm6e34G58v3pHqfM/I0f
9zw0AXHjW7VfaBg5CJRQtu8SV1d6ZURsdSgoD5Yy/JAeMD6jdOQxnmpvHta16EYZ
y5u4HptQFEUth9dNlJmKGNQZJLDx9yqKG/VtUtKVV/jVFGJ5UixC7TWX4Vm2yjQd
rJFwr6r1XDvFFMQe+z3WAs3QxTwt+WCO12wqGGzaCasvhn3U0P8TXMQBlTqiFIbt
A9UaV5RYSfqey0fCGzK0GvwaMI+lGUViWRCvc+bG6LGqx56JBLv9Fvv3Vg6Fan7B
s4BY1OiPf2LjW9GvpnhfseqP94XqTbaik0ZpYwUz2jTCmuIu7w1fWvm6MLKEC8So
JxsxSjnV+pI1vh9ukqHM8bn8gnRgQ9TXvuNfq3ujL917K6d/Ki41XKc/iueiYRUU
Pfh3D5lGYTuS1hEz13AUMC/hvzgS5GGbYjWpy25zecwg/H+X0nX2s6BIPhZVxYEJ
s40kjDbrLPapX55QeDu1bVtj3LbGby12LPDep7BQx1vTBJT55gdlSBeJUwwga7ZE
OAP+70b4g3VYvIWas+mGqIYB2DJpjXjzEOxnwqsNffd47wSQtlXalQwOaLd7bh7k
Xi8Q3QQNTrNw0gwrEejCXGfkYV3IjtwOEk8EaGxWUaMGmW3DSUiR4IxDFHAf5m+s
4ioLKbKT2aNTaGFksu4T6KTdsof7Jxo5wcAN354RmTkxAGBAKSD2h86YYvMh84P4
0CmEanchN3Rda8mLnTDHFa9V5sa8mKA06u4dSOdaAXGY0SwpP0xed5klZhcJP9Rr
5/ZLlFfHZoDfzyg257NRxdN1QwthOmh/Gghr8U8uMa9DdiVInLgDAW/2GzYG48lb
Zbbg28t6vgNhhbxKbesT0f5STV/GRc7UEyiHa0/9AulZS8a+saG+H6lk7azPJri2
4t/LFgl95CY+ptCyrHkL7b4ChHo320Muo0w/tb81VLALW0pZK6ClHqqdZNG2ibHK
dU+8xKxlkrMD+cs8n348AS9qcO9NOGVSHxvis1pDUoy5bVIsQQHQCHONyxIH+qgd
A2PsGzWwdt4eZhesIgJQQJz/20RovPzPh893EDCi8pmkZXEweXMGhcQDSHGc2yVw
jFlAjtjo22EErMtgtZ1GbOBBU0atZ7S9Kyd7xRRikQc0V3crll1vY7P9wuZo8PBC
AEWIeP8ZB6hmCWNmz/ogDF9VNJfzRVNmmymwkDmikETIZR+F3Qy8c+UoWs4cwZd7
mA1mh8FWOjvEWRU3qstgFyVNWYB0VdfbJ2Mg0BQ5L0lQUoriELNMEOQcIt3OXcod
s4NXfUcDgsfbc8m+xbLNRgzbVWpLZB1q39DVPOxHOmC1nbJfb+bvLrVuFewvNdCU
feehG6kiv9R9IbLblgHAlWx7u5ezYEzDdR9kXPE1oTrgIS8sv6jZtCDS9P61gXKu
t8S5YrQvsCGZIv/YGuIgwF4JZGk4FLkSfBLf51AL6EMoPydVoZuh1ZTqiAUvGx1j
gAGABpAsaLfNzbEyf7DwhQxnLyoIBfu/8Vl+kOwVZPGt73sOb3k434qYY14YT4qi
V2xFHDVmiHf2xR9IHO4XGzhCI67hi+F/fiLmZLj+xckyxvm6M/+AMqs3vmjNu/dP
nS4isnetko3tzkv4t8Cy6GypbVo2gVgpZWzC4XwEu6xnVRJVqgM7WyhAkX4wMdoN
QsX49p+BDPlz0RmWEJLZhSu1hQJqm6ewDC4zgoRL9HLlJHvI71c1o5cYpwXiH6jp
vhszponUSQ3AiYFKFSO1SWenAI05ujwU9L3N6i4BCR3/eDFHK3iuB8kC93JudsYm
J04rlLJnixhmfm/oszlt6vxA0lVP4mn4uGQ0iX8OIMp1OOKD6VZ4KmwP23717iR+
hOHD67LMF9fjmrlrtfzidl9G8AGJ/gWTCmSNc1um0u/7zEiYxTS5eMIpntSTG6yS
mF5NI5TvwCzQ30lEHmEspqG12iIYU5Ccp0DM0GUKTOrSdxQDCjvh4bJfqca8bdnC
4pVHzTTfJXAPUnNobEnKoy16rf35rKr1vSd349H8vZU56wI0nYoa2Nmn/aHc+ILp
EFW3+QCLXnXXhvZhzyuN/f6pQd4HbDI57GAf7kOD/8s3ROL9KYUPqOCc74O4pqio
rRUY+NSkjjg2ntNW/W6Bhx5GeR/KUvhwEwcetjm1nmxAdlkEiFWmXUuBJvsKponj
jTBqnaKps3zg8s177raVDFijYXMrJtc3xUxYMIuhNoFBI/leuVTi53GkZc2Q2aEz
IRz4r/XJwtSiXIhXLzYZgw5TSoHeMZrQuBEVDLyEUmFBqJcFY1sX7g7O7eMH6Xiq
ikvb3zR2b+qMHyZDA7G4wUCv8sBOrSqxVhW7mQL9mUUxHDssdOXNforcajB/Ha7C
7SRErxQVUBWeLMOvwJYUQ1GDvJ1jiLRI/CD9FhWjUAfcPZ0PI/ev5OMIkZso5vQu
dAMZDWZZ4odhQj4jRaGW2pvxkh9R2DNsBFqI8Zz4RpQBWYWNGlEzG7PDQClwrQgF
eRZm+sCe4bxF74/E8tU2gQcB3ndwdCZVKIYLSP4qTF+q17u+P2qw8ZplmEhgnAJx
DlvH5o5rqIz8SvWJUoSQWbad2TbF45qhx2DuMmSBWW64DfHewHB3KOn/BAnDYSBL
cqa2SffCsSoYF8/qO8munYiNcohhYZGZ9i7/RiiHQx5Ki+4j3Xlxml05Ynz6HU5B
1vhslm2rdeO4SP5b3o+2bPiitnnYjUWqliad+GZB6FfcPLSekUhezGTvOYDwdyUm
44BfaQ3GX54LinU8mdglrz1WT8ZU5bh3a68S71tLkGNTT/NPafTErWh/wvR86ub0
3cIAjPS3EaN83vkaa44BHSwINo/TTkvoHuX3IEatobaLfC8JdpV+owi7CKSU0lqP
k91fdTXEslusmbT3oYXisF1sS3IrlvK1Dck/ZVT6w59yBatQzD0sePhxY40eiEzE
13LVx05hHPja6NPHu8XBKcP5rrQrFkx96BSPcdiv5Ck9+DMnmElDAvZr5VkRr9Dn
Z5i7w5O3edAkPUh29n25nxcGfftt6H9OzaUKWQnocpE407Ehax/RX7xkipCbQ0+7
QBCyU45+y8bG/AxmTxzBszxhCCvAiqMwnXmZDbdIAPNcl31KUk08vf8rfpbGX29I
0nfTJNIrpj3HPgPzDEte/sflj86qf9LOAf8JVNMwhOzBzlFBO8xJRJEkgEbFEnKC
9aBYb6MpKo9VpP3dRFPWvn/Lt9/BylGRz4S+uNu9VDWCB56bfqPiLb1+xGU+dTJK
z9Gjod9WQtmZTo1EzhFdM7RzkUafFsdnKvhGYBICyzz3meq18+X0hUi+xQtExjAc
zPQ0179PB/r29NkDDS8sG5N8UWJBn4tTiFTW+X4p4FTkEtn5J5rO1ru+EyIKrh7i
bHOJlRJtLNXc4xpvY65b8dwRMSQvZn349Q1U564QtPT8Fy2q+9d5zvfsA4E2XGcS
qSZDtbSwKnQ9uBGGe7QG5A6SvTw6bC8gqe3ekhhcwt3wHrpKgT0BT5uLXSEbNI3T
qGr6thBcdrG6dGct/VQKoYwRAbdCpBqsIsyrej2vc+2iuFrrzQZxdN0fbZuxAScx
j0WqzowCx9XUbP3tEft8eJMGrtcw+9tme2pk0EzkAo29GnS39FmHX6RDfmMHRNBz
Mhe00UfxANfubKDgJkZAWhsxAo5isjbOasVIZRjwucQGxEs2khWM+QuWf/rAMMDe
Y2Y+xVL176tzxKXSTpPwdBt3VYoPgwy6bz4BFJotPJjpIlDj5NTLNeREpRwzAOxE
kJhj5z2trJcRzPjW6ztM1tdmwSjt+SgjSSGNzKX4OmTljU6IyT8SGuwDkzir+phz
te1oHJgIG4CcyYmTLglPEpbyltaDRKsGo6G6+PYtjxU44p3EYK9u+t+6Z+9MODYe
bumhU/cNOI/RQXtPQD++ZsqJoqjfoszrzlgKtxdh9lnJzIKZJ9iFrBKDw72tVl6E
AUbEM8cHe0eudfyF6XZifINFSM1T29/Q+YXQayXmQ1Dai44oMH+G7TqP6+DE8/vW
1QV5czEs8BSmEp9D8kqx2ux2RqkdFlEHSIUZHcJgp/69K28Ovj9zQwprHQs4/kaM
x5a95B0m1jT2hAvFz7jDAezv0HgOp/UJ8pI6M0rw0WkghWJ0b9nRor5PWVa2G79O
GOThPJUNGEWGAG8XGVsuBza6cWxYcZgqQKO5jQaeCRqGU3HnrwzTsXmCp9loK7u5
htcwtK+sVWaoPp+ZxNvOZhUXUmUcgRzqUejZjnl8lDuXy016EFlZu7RO7PP0XHut
7gqb9cYivd9byz2Tf07fAoxcoQTnBuNtfTo/rc9d1RRzME5CuU7FBQuaOANDWBA4
abGw+kOpBqsALahx3ZWsnCA4NEkks0vckVBfV/aaK0e3SKnIdP0Vudp4tyYGMqBR
cGywiYJ8VoKww10RwxnaDZzSOn1LZ50xpU8EnISnSryqFXCSQNv1jnH4dUppNevj
clgcRtnRBOpkxS9BqVdLvxwPCDMHp8R1+0MXeEm6R1SISJwxk151uCG/yW8/Glil
n+8BXtqZa53Pw76wJ3UHbgflOZVOqmmwZETHSC6eWn/pPs8DoEk/bZAe7Np9E6EL
5SWZ/emIfhJHBynG/EIF9B2OOqhq4SnOBc6EC4d8ZPAP/rXtHzdZB9gzZhfDSOnl
B1bNZXzNSG8dZv5IwX2F//aGceZSxgotfuYjS0DgM+8+gDEG/AemUOS5MJJVhhbY
OOxuZQIdCZfppsvaWUOjzRqbCNESId1KIN8XTesK7p8aWieL4RcotKlMyReo0meq
koL2C0KIVsicPYzGbrTmqa/jznh1N4uEil0tcs/W1O90Z0i0ctDMbXXlCBxhleOD
uJKDkn80PEwz3FC5XWj+xM2PvPQ60FgqhooPpaR7gZQSWF71PBmVmWmcVEu0R10v
ni9OgEX3liuGTJwc1q0/RbQ9ySAXbZLzxzmvyjoSmkqpEg9gEHJ5tFim6RM1hROm
laEv6efijndaFoFYrDYs7NNpBFoNg29osBIxYUeCHzSuhY7swyBekFi3JgJppnkD
urjBzYVvUanNnTaG55I2GliDELRAeLXIlh5TkAefDYJFP9GJ8dmVON+KNdvr9cqZ
Z7hOILpcZ8QMT9LJJ+FZqYnPXui8DN5mnfOxnz63j9U8TkUDBe+UBgkSC1nkmkka
sIyCUEvO2bS6fOu/qKn+8XQTL4zOLBW2vdA6eQtsVfkm6KjEXoE2Yr/Io92pN9cO
KHKNwiEFzjtvGEKyYVqs+UzihjJRv1KeGfXyuDPjuQmXvyxrkKTQvpHGMD9JnEGQ
g7jR0tjQyWV5Bf+AC+WGv0IBs5M+VJxLigZiJxYdMrZ5Z+esdTHsR+wjC9413Fg+
gkeLSHNDeqJuYvKg+vPXFy5Rs0nV9p627cigopev5rEMxMuvtmVVQh9fZL4Zq46r
B4llu8yCT7tmHw2fmS73CtQh4aX0yZDW7bU9JT3vUECIYDEI8QH+lAg9FSvdo9j0
6rrOkV/3QTKhaAWhtAmYorYQlaot+ymHm42Z5p3A10VyQ97saf4tEYeFOOj3cSw7
21r8mfwfO60iqNyBFqATsbNG5Wyvxfp+48qobxOwAUz1Ch3qA7OtFwSLTfJdHXaP
f3T/+wmiBXcfXTDNLAfAi1CvPnz6XszMfBvmhwqtHb6A5H9blf88nJIjCaDLaB+q
MVGQOta0P8v5pQxn0sTSWS1s2gdhsdl24YCvg7sPXb8nyOczfZMT2tMzhu8k2P6g
Q8StU4nExfjG8hZ3pB0oVZ7fKpht40F3eQSwORUfEMVeYcCG1LbHNYwHy4aZlV96
RnoJP3dDw00qSDZFciugtpeT8ZjTXDqf00TfrZy2RCiaN920sbfqdGGeAqVjviXz
kG+N1DGY9tRkBaCq8e3TzsJ4289JT1TSdGlyWdnUbphCTVvqtTIDGJco7445gGoP
sntXQW3yUtg65e/yS/hB3OCczAxcR5mUMOXupzRUXFrKTLpt98gRPXu8aJ29H27V
O7GAp9jIWGiGmXltNXiwADDOBCWdQ4NTNI/0wVKsTnf7MjPfdnRQut6jzYFe2kBa
1t2xZj06w9B+eiWbENK1o1Y6Mnz3abbh7fjfQTmgvScxbRd5/Cl4K/8V0SrK45jw
vh6zHrx7XvULwx35nduUGgwtc4PP+sNUkLzYDjfXZkZMEOng6CKskSIZ8YhrChA8
QNX1a4OOpzRaGuC+mgleKexnyEchSLrJeiTyJkgrCZf40GNA3siTL+sbfmWTj1oe
zJxoFRpoK0ignwnsDPsglX66t4oT67h3mxXZd1qqFa+CgtVocp0GIyZZQKC8pizt
XHIfBSHpsT3kWUE4SbHM/IROPOrodEl/T+iPU5bv7rD/b3Wrfk5BOjFNE4y5/Qxi
7nEId47Ez+1zm2ebk6mEZ7fTfN9YpamFub+OXhXTHYe0Lj6O+Mr70/pnf6+vxfQY
6XOojbewvrZQSIvDie1uMWy3/cQnTLkJ5fRKxMv0xTSNgRqTZ58rvu1MPOxVmdAg
HscHRuhzciGr7goZB1HA30J3c62yT1izLGMDaOsCwmGpDfKjdfSg/+iUNndE2beQ
xFljwc3txuAeGwzSVCROtz/u2n+oAi5stQh53dstWtUZn6YZ8lbJHabkyKBPOFhD
fxTcPkqrJkJR6mt9/OADuXuOdzeFoZFxAn/KM+uaet99lXktQgYFYIGFHK7Ixr0L
79mU0MU+hAFYq/hZynGVLP6G2MT8Vb4ZHLCVVPSrSXgZ0tSirngAChk9quefIisH
ZwN5grkyMgMtaDiPPpFhigGujr8m1sH+z3oP5Dom3KS8r4iOtKjKIOmsJ9J5izsF
meWVGc1ZZGMgRn/v5s0tWYbBCcN1jXcxOSnaRhy0qyPXwQJvxLRGdGFB8Ewdbt/u
VhYc4k60fST/bPfs1N1eQy6Uc+EsstIGhkHFIpCviuele3xQT+PVxkl26LjpmJZg
CxH474dIgl/igSNtdFs5jn6pG5gh6NXuvIgzec721sPhnGbnl2lYtOziSqCSjjvz
V552FRToST+Y38ogN5ffZ3Qy/6w/Aq34XwJWE+ZUFl2iJ1F0Q8kQt/zQWHp+GGCS
kG0D5lkhaaSiGHM/9GRShDd8k93rxjvnJ/BGdPjoBuogspvtfLFZkS5Erjea8ors
OmVcZLwpb02bsJ1aOaEdHNFj35NLk3T+diYpSQMCPPFhb0rcbBSD83uIaRo0z33t
Y4tZVi2X8mJrqo3Ozjn5QTv9mlNCO/DqgmRzIZ2OBIgYNwQM55+m+KTzjWu4/qGO
cSaKP90XNuw2cvEYwGW+LxXdLbfzrQzixUR9dtZPUImDH6PnLFXDQBvnosI0TY/R
0GwvGQa80nUcxitVOwXZlmVDkXxqXmUhH5cx4Ppfvf5ykhSS2SrssDnZrF3XIh8F
WVtg8l2Q4DnwC9Hi33wcxt5oJUWNJWcR+sIjCGLqN8PXpBCW13/I++isz6o3+TTN
N8ScQBnfzABNwGXphB7gEoF/kpKBi9dOtAJppX5+XMafZ4ep4Km3Xok6O/3pEXX0
SXvfrzqdeNvKvUVOzwtDajxjxCk92Sd+g1IEWjdTv81Tq8Sn0KnM8B/O/DNsNWRH
B1bSg9JyKVidhZCnq2SkBmV7hBsUe9XvBPhmVaQnX/A0SdBj5NbEzzdkRNQ8TVdJ
ctWMB5f5GiVycsGZpv9ZLbXGKBepQsQ8BBjXZZnDNnNjJw1wLC9QWJ6/id8SJcOl
p2UzWZ0n0UZn7b+wXVIvX8gufLsi6Rh7CM5rC1Ptrv5lKjKvI4yjRGs29kghQbxl
sy6uVVqKy1IGG/x7HMu7djVQylmntVXQmaqsKr9boj3eY1Y1MApJqrLm9ljZUl+D
eRGkFUofbI9kOf3ZW3mjlVD7lX6QT+LOmK8trRDpf44EN3kgXwRSpHUz46yMRzwR
YXWGmTzBmaLHqRTCLawWpRJ/phZjFK+4xyXoW5y2WReDtVfWZW7OaDVp68BRJ5b/
Np8s+5a+vmQQ8HzY3A9uEn5DAFiyG8A2G7tZSJRaVyvWQov1Y9DgwOTy9mwSKKql
g8NK/GGuzO9ntQwFCRaqcKqa/Fp44L7rzvjg7egJJ3UMIIFh9KN/ze4n5Mm5ve+z
NmEXnbP8wBUVhXmgiDDewferAr0GEK4RlF5Qty+D0g3vSG3NwR1Ap4aBbBccIbwr
bDvgZ4AcvoVQXCyXCXa7tOaktYOfE8LBkTRagztFUZEyZVIX+OF+GgfFOKCAWMfn
g7+t4m3m7hIsB0UuGaB6KA3CgPc4a+CiDyaKq3ByRkr/TmCizgx6mIWBCK5Moffa
OSrrP7rb7v/z3G0cmFLGL4erjTisDUaHTaVKUkNdr9X4okXQjF2x7vc9tYxRRWJ/
bNyr9hAt2670tsbnNsCZ2nLYSkrI+GbnLX8W9xzT8gOfZAVGSymIfxEx/ma6tT+x
x7B6uvccPV7yr77YMk55dKufWdxrMjlPLQhw8PlArfBPTxd97ONducBqqhZTyTH7
bYYmhDnHkGYpLNq7kzBN//qyeeQGzCvOFxlpRB0ev5MGXnzBI3Kz5dS5WsweTFy7
35zESO65Yg0kbozr+5VfVvLj7EAg6JvFmRWnApNU7z4ZqYqR0ExCsIOZmlPs8nxC
kAYO+Y1RHKGdae4CwwpJ0R5FKiU8OVvg7/5ISsJxA7QzJtBuIu7N0pKrFGMXcKJw
QyqQDqpQo3jE8tXb/iA9/LUVcHAMyweZWejsTYMmhrjxAjJXlZcQTeVLdSFe27We
w9gn+Pvmig9lhWt7YkqktdPEBM5pe/egp4NMQc33uOFJ3GXNgibJ1zQBBEXQXBOo
JRP3ei+vVUw3U8ODYeefdZwWgYK6qT7mJfvxEr6e1FYFyNyJPQQGaSbYl1Mska4b
NkiF74itvK1dVCI5b2KQcftAjRJ6G1GsdTAZB57z6c7VrMBzTWR/WH8etM0K2bd9
dMwXR5synld8Ih3jR5xu1OWFygui6g4B8bsthaDutO164pEuQ4DajCJb7vW6af1k
6sn7TdwLq3wIHjb1JXgjXs5NrY054O6zpTdBoWGQzWa7EyRRsk5comlCdNAd5A/+
3U+SLFHxf2TPdb5hmno6TQWv3mld1PN0t2g25aARVCcI4IJoFCwXRy9VeSyBFD7k
FUDv+N5+bIYfZrMUawOJtEvaPd0S+Zqxu7t0zshrbBlRkpCdpUYOfPpcR6kw42G4
Wp34sqwQLphq6qPk0oVx0SKjMTzK/7N+e8oa1nJ0XnJfd3r+2iCHjtwEyjwOLdy8
e/pTKgXfUbH3qBEBDYCsAR8MyNTO4ebmMnDSgQbN4gepzstg4s82tv/u/nsbNXGv
asdUfCjzIxjYJFXqmqEqv5hyn1NABoygcZY7LPtvM2ZHaoc07I055N/kOmUwCBqW
AvAO2s8SVACOzCN1whom0hhSpkYGksPSwEstWPIWZZQN3vH6krmyaUayM6JDkSJz
65iJ+H4ctEkOYx5HzFBgECebsbWW1llgN16pKFVaeAJNMUZzs8aneE5AXP4JZta0
15HX5Jf7ClaLgdZyY7rsMkcjMPuZ0a7u9iRTvKiX/JJnuVZ5A7/rSomaVTsuMEhN
JgzzzM3nCaCtxOursT2juZB+HuJHSFfdzb4CWbm6GVFtPPiuSegOa1iC7MZtmbF0
AiVTSQ1beNBVe4nk1C158X0mABqPtuJmZX44bLdGuNv5Qrbi8vCaahk0yiSUn9Jm
c5ViegjV14eG5RcnvoeIbTEadCHk8LhiHGDDqCIoPi+LEjQBwg8QvGaJSMu3Zx3W
73Y7H3LU7mDg3sNMVn1K0tTH9dAuL62706QlpLFNikobVTkn6gJIMvhwLsmW74Mw
bzmuQOjx6HPKig92/RgXrqE9xp9kYaUUhcywI0bMbCb9jak5/bayQFeh/xvSRD2i
3d74QtYRBa4t25Sdf602H4s0dkTlWgTOe6YSY0zELjF+5s6AVpw+Ov2dDkCkeL9n
h27sudHznNVed7QeP5YxBspVFfigT6a7HUgNbuDQGdz5qM7ogVyUruLwozgUkbR3
CpChISjf+tk9MUsRRkdfJwU5jjm0mbNBnlamokMOLzR97aHzYdDPY9jGUvgQ8cml
Gx3HDf8nePJ5UY1kLAhgl3mlfhnOWiceMUZNb88MToLwwDQqkqOzcuHDkbjsWdaf
iGLv9SGb911fJKEx9SD9wpLgBnLyQ18rJAK3KBuId9BD4YXj2zYSwmNtv/04A8j5
1rBujRaq2UWlmnFRVqUaME8kRgJmOS5wGt+5b47XUzSkJCr/uTvijqZC1XpCz4Fd
sbYwMGaXgtvy43j2tFIAVVyMjKVhPNyHcnYvvV5sIMcMoIFikZ1q+6lB265d3oEG
XhRAtzRQxPDFLjRuM+eW+yH1fwL1HBnLdQSz8SotjzlVyYkymIyUd1jE8ZydxMae
V3F+8xwFtPNTKRGw5/B/KABvaB1pZit301FkqUAopvzgkaiFMlt+AmjCwuvpqskM
tBD5nv2z8t3xBfMGG7Tm0S2XlPKhGtCP0e1Va6YENz0EqawbBG9ApTTisIYG/xyK
5Eh2QRs9RsQ4SgoyeXu25uld9sJa3RvMvLGymx3GrZHeVxs5Tq6U9L/8c2IFPj/5
nPubz+OUNfhS9azKl27TbxrwBHrlfiXHR2gImtNS/TtV1K0w6YfrdxE8uh/pRRwi
Q0eYy9XKAn5q0gw0lkpWWKEyHTUGK1G21IFWSbT4/9LraF8l3SZqwZgcVn75WJ1B
XEDomcWonzbYiGJPEqZqAHZ19nb2q3ooDTfQLfQHtyy+5KDJ/wynPjEoWY6a7J7m
m0/sLcyf1LpBGw2fb3c7xGhtOsV3pKhQ8WgWz1YXtN3DdcDQ7AztEp1n1dH8G9GZ
4QKy2BSN/N/U+3lCIyHpcdt6bBIXVZmKHLP+3vu45Lvf3EtOI3xAwpr6p0O8FSRZ
n2p/3XHdzdiZ/MCVkeD6n1nIiZR19N8peXssv2inVIJv65IxGpIzdg3EnHQ0Divr
TNnf5bJLwv2rLwp+lGNxKb34/Kt2qcJFDUw6xnX9k82315faBCtFCwcy/hzTOEdk
ZCOa95XXDXx/Z5Eqe+tG1kJuzkla1kfCkJxGC+BIDn4kzP6LUigSwJy++J2d3cHm
9CprB8fSZhpdwbp4VXVNbI4yyMIjiozOjefw7uftZomK3txuoDkkBiYSPZTFKqbV
lT7c/sVlZz7gJ7J4oEREOzwnNAa7KUvUoht8CICiW3x0HvNkEXmSfF4+6m0V+1hT
TnkjTN3Dlk1GwnpUWpE0BBC+FIrRdXXqkQ69qm6HOsm8oRg6f6OL1ryWWcYvQX+S
BJb6L02NVc52ZBPBYsrClCegSMqBoqObXK7QxzsxTCo15OOrHy0cWr/VU0br0OoE
qModHumov10zFpH5uYksYYFNu3B62bY/6WbsgxKUqEclKntte02s0gGGqvn9umBK
xfdxZQ6ticycVzjzxHoJR9Bg4QrKgMqRALk2q5nRykU6c218vXgQHgCzl6hgpucM
+nOy8izmo3qlTOcOj5HkWpR8Wr5kcC5LP9OXxCrQa4FZaXHx67f+esHmrH5T25UA
MJjZ7pHqdQOTbWtMyMx6DSRMjgAQOmayF1txldpaWq88fFEI4YUwDoyIhy/Ve+g1
pNOg4CgywqBihpn/FBpDupKD647LQL9FlOqCaA2GZIHI8bg/1PxlqGzMVMtxtyT9
SygGMGXmL0Y71lDmBZGLVIbCoeKHhILepuy5g1YllC0gFxXLOLDNdrQO+AIMrIKk
hUVSdlqMKJLWXYPHQ77Llzl8GcRTiNc/DY0wxeLWxULf+JvIka0c8lwxx+WKets5
5k7eqH9f9jgnEvTxRtZSF37vo9RTlMqoNhhHzYrxSxJDgX70vFMxT49XEZNSJPpV
eDlNxOxNuoWF28mpPGBitBsPy4MbcIu3vPhlFDcHFFkcY+H0nLM3hgFn7ZsZee11
g7nM2J4svWNWsiThaaggSPgE9yTpnYXjR10Sw3N6Ueb2l5DdaA5VPwd0cNntJ+FS
gcxDI0Cy8hOFsBM5tLv8Rw3eCiTdFMM6FHeV7Bkhem/+Snpy0IR92XuYF5T5v78o
i7oD7Y86JVj+AIYEPPbZO7vsf2wgkinn17S1PBvc731q7NnIwh4AliSrQO8SRWHV
6AI0cZgW5qVdhZymrY61AbKywiJxSDPXtQB96Vb8qTouRtso5T+bwnEdX9p8H8dQ
0BuLtS2xy/FA7vO6UYGfNmn6sCgO8EyrNcLGfuS4b+squq5XReFSQvLFxv3/8hqG
JuWybXRLs6DS0e0Ub2vR7DF+ilNhh6BNT8fWTF4NPzzSeXcuZyP84C+K/fMT+mBN
+VMIRw91E4O0aFNpLuZgUGa2xkwn/j3t1paxAe3GqP7rJt+q3Yb0Qj59cDMfVFWZ
2nFvWRKSf14pOmoWTONfgcSrVFy64A8W9KQU5xquf/ehH5GvN72ypbdfr7pDzEiI
gYwJlQoYYrgEQjOr+wSuh21o/+pzhl8pKEFOPjA85wCFTIpUS9/xzZWepqXT6RkL
USg+zoZG2aB3Vg9QO7YL/WGMFZyHKhw1h+HabPr53imo4SJRhKzeVO8A9FuRKOb9
bWaJbmf1spoVpcO/FAGZKCxlE+/VukdFG76loWNqzVCwZz5nhCfzVhaSWmO2c8H0
RsUP8Pt+Y2+SRt6Mk7rP5Q7+vCNN8WW5JSoln5iBJ1dGpNAQVsjU6QrPdg4DV/fz
gos515XxVXPbE0ABI4cuX8lfHYzr2UsERf3LNLquI9B5iZErrRfdVPU3bdJ/H15j
+RSkaZ9w4hKkolOyJn8CIM00gKgq6pnOFKtzIuuRy0OqgocCOHxAvFjeqrflDeuW
ugvrov1jhCVu19mJghjdlYNdyhUxwkqz2nQrWw3ecsvltKNzfKEjTWV/nnuyG2vg
BuQ4ImA4bs6RxKmrBa4S/zuxB10AmUmHupcirMyelNDEiTNbJMxXFjDbd/wFJuZc
LtUjWBP+g682FD2QBSavuS8pgZ3obClLbl2ceyQ4zBOfVt5vfjGkQ5ffdT7J9nVB
RbETYMtLmfEVXh+A7FY5CtxJk51wK/EhfU+2++F8l6jzFIiSmlDKGnnM4ysRt6cF
5GiIDvRvATnQ24mXL3DXua6Cr7DT2suxKcgOq+w3c9z9e8z0rbTWaUwmepnr0HKa
k1ypDC1wTvb7NCqnkuspb2JGFEvyiB4lhWxKaAEQeLHXsvyrIERvrC/XhqnLQBO8
UdBoKbnQ1tSS4M2jQjB1fH8DPIS9TW8iq8IKwNs98CU9KJhcNTYppAe9Pg78gmt8
ifQbptGiQO+E72CAtfF5pwTMQvsQJ8ItF8LRvbY0uBhSzALcdkKTctF/LLW2R6VQ
s6OJzkxcdQG7lhlG6Tv8LcW6Z8CfxOHS+mFK+yIubXy/hYfVnHgh63aWdh6JPtf+
ycVV97XGIiJNsYeBjjgjd7v+faUrq3AKg1pNCkeCPDAnBGybA1jiJN6yKhnqhYgw
Fj8QTpJs8Yr0TTdwJYOSjl6bzXo+DNk5rEPIrGpRBbV31iI18VY/mWoRkZPm8wDv
WXrs6Az/obUWl0F26geMWGKhw/YTSLRYuIiWNs7FleM+T1GLM8fYo9ttUnh0MCZb
jCA6bpqKj/lVDYVDITUqmNw2BP5yDcFaNBye04tyxt9aRTD4cExq0QkZ3czLZxxo
pY4ZCy6IEyzQnTC9C3Gcxo25wFew6wBAhIoVAy/C3gRb1hqiDdaya24AJNktt/H8
VNr4qB3EZjeyWRoNbLu1C/T4GZ2WJgAlg58IPL3l4NgcqdJEMIAKyuz/msrgLRwv
qQOyU8LHwTIbba6YOU772l4uBMPki/vkGj0DWpT+K85uuqmWrLjSaBU9qOucYrZS
rLkwyslYbom5rCtEqBn/4scwGwFuUXXjnCVT3e48MBkQzUAmNcJMgt3OSReHcg0z
dcxLsBcTG1R+yMMP25ioUQ3whmha3FgRjU2Nxz0wpIUWM7JmwXxgKjy8e837aon+
wN7Fl7yRsVWihA6ds5zKMl+L8ygIRswLME3l+EOSAg5Ii1n9/wTTApm4YR3dYnK5
s8vlE6ucUIvnIG1L5qtlk4GeCP9ZF1RVPyi2LaMj6xw3coTR9K30iqtCb7LBxmUs
6jnlcQ4E4ew0ReIyPjFVf6XUI1zSNaNyieRp3AGx22ZRag+UBuwrtvTRcfMmTV4c
Ii+by+GVLpewDV3WLmqYR3Jtb/vof7Y+dhwSl8+Gag36AiZrY6EO+kB53GPnNQpz
0Qjk9dQyaA4LkPAMlpv/XNBMNf0hxD+nziX/dR4I6GHR60ITWZJgoGNWh43Tzy/M
d3Zgv+SKVAz1SekWgJuJYH0+R2x9Bzo3jLeXQgfoEyrY1GkAMjmYnairhqRtC7Q5
cfPB/Z4vZBgwB9HoHq2IKHOQJ/XE3qLJjYCCo6bzjg8NJqje+nlZ2XipdQ9FAKae
atmTST23oOqsdTklVnKX4qAgealY6UPvUSHEyM2vlBw9DsOH7TqwSxzmiSvKkHJH
kVP4mXTIO4dA7QAoKyptx+BpwRHvR21siNaePvvVyy5mNenEuf4sov6vD9aivnjB
hrfHVL78nP4CHFR0qPmncYWoeiMgCJzbPsy6JS9dzRDxttJjhvckTYkmkAjpRmOk
QLfhHukIVBdYk0S/ivxWGa11vlKb+beiUFZuwU4pJiO9NFvcLad+62cfOZZXGjlV
gik+TtxPt2gDrB9iJ3aB+SXoj/OEjXpeP4mTayV95tDZXEpGU9mepjbMVHTkaRCO
zZtt3cgrWigsAgRme0JiYCmzxM3+Fk7E00w/EtBIFUmU26vnqpii4fjYoqWXkrym
dZrGWWkGjKqE42Ceiwd4eSMuIP14ESprniDmL27orHYSGkvbeFOjmpDxhr3sJ7n3
TNzpP1rSOhPE5O+W9YMjWDBdomGFHQUdrN/UpD+X4Ez9m0g6b/CPnhXReY9oz3qH
vATdgUZmBX1iaZp9YN+Ler1nSxrfAYuXNF3gtYgVfhr1xv/vAwI03ZoHMKqRxbO/
qdR9TzFIBGTy4CpJyHIt8HCsJr5q7XuXRYfpGMtQv1u6rih+JT0u9SjKzvvHL2y7
Z1SYhNmXQo862E5mwBJKeKQHdAd8LpN3e7gGQOkvO9BpPdYJve9sZ33CZb5V//tm
G9Fn3S5BY2Rj2pfbUxg0elQRFh7G2Qb2jO5K+1AFvRI7rMSqiSV3zz4Za4G1Q6nl
uSuA2wAKa3YLGUG/onJyArrVQ+omiTglH2jp4Kz6/2ewly0PXgEblbJCFcQhIDYT
bj1/ZUe87EIHEzBQmOlGZfffEMGznbnV0wzzAiWwfdKxXtWhUUfj9cBwfcjFtyz+
y89RO0WRgptlz/Faap9NDkeBxJquYrDdgfD8pj2Jl9fPHB2JpACDvVtNnGsgzptv
sSZa6F2ZcKt7OP5BrtCuZlXmc5L1n9PxtpHQg5Uwv3FwDtcGgSgHox0MxOYqlmeE
td29pMHeu+o4Ad6oTfLJ8LDwGb4EBPlatGpXu6oNmyVjvGZ+7/Tze/l5YLGb9xbx
J5MfqGkcUg5q57XVFBnpAAiyXG6KRfss1Ds6EY/5iS+Flpl0w+SUheMc4nCLkqLE
BllZw6DErhXoons+I/j/XiBGViPWr/VWjej2vVjz6w4tc58/GsQPy0jAhoFl+MjT
2DdZisEXjqYU3XHOG4vsq6e2DOAMvAS6yQNaYHH6IX7vGzuV/zEqO/cXVJjMItRy
fBEnabp/rNhGMCGJ9VgaJQ2EYnPyv5ZRPps+r/aqxu8JPadgVIcwgyWa9k8+7lsq
fVmPIbW8gX+V2aAf3TMbtxDAWPYZWWR+twiFxOgWj8T5acfb45cA/hza/d6YywoU
0G33VOOTCdaKVyddnViHhMb61yihL6eCn/tDZicT5M3Y1rziqn61VGKAjbOjN/V7
zOneodSwPcG75+mhpR7pM4Ew/uztGOD21fipx9dU0p2k7F0CgmI1O3VqZAwXV2Hn
gy9YhHXErnY2Pn6XMXtXdAHO8tR2vQUC9re7D+vMDd4ZYts9c1UDXItb1D4xZpIx
x3EeSq09oaROpqiwA4DCw+6dq+LkuJgYioH/TWJTpMXhnQtob+CYMiICW6C2hIaD
KMkLXfv6eoqRIWFCitqdIAwOP3LxHGnb723ewKPoWC4fR7HcVqAQtYmnNm3rXN+0
gsx5F7gScq6wE6uX4iJs/T2s0Cfyz7MLJ7fQgNGKuw0BpA7AEs3u5B9/QV9z893Y
pNs9RSGEVhZlgEC03TDPneNoCQg68BoQWJQZJ3tYrrKI+1KPrcQMPEHqFoq2A/Lg
kNPYYrgur8DTIfOR0M4pgFJXYnLkqfXNzdR6//1m00IT7JWD6XLcW9yIGCNP14SR
g8FW9UWizMFGVaOfTwLRQYLbxecGbFyChp7b2SAYfjhZxoDfl0OicAQMuS5YBS19
toXtnTi2V2nQspbjlTDl3UT/KuBSfiLPWCTDFEoYPKmQSt68FIdpUf/s1GwxxFT9
26ZqNxam8Cv0qpAxvbp9paXzkg0sdxbXUX1DQO4RmxOl5HL35OxqSIMssv6CGQ70
b9LkXM+75OW6Za0l1Jb7V3alZewBxNW9fj5O7jaAJvkuG0CTkuD4A5DqiVP0+lBg
HTkp2TFF3PVuKxqcSDVA21WYTPeSXCciUYSuPd282GKqYRvCtPLt/7ahXpe1PdSw
0nJXGIv03uoteo/iHGca9JiwcAxJNFqtZPsuepV67nGg8VAUMKnoeYC0Q5I8BgTX
0iHLYr8NJPDZDoXoxX/V8jHBFtczxU6DLY/dAATBzQ/9cCV7BvfFcBG0xDcF1akH
To+Puq0w15lizKGld1GJIn3sRDJrb+eFd0kalvJ1FmBpe+XnI7j2uj52GJ5FLbd4
b5E15s2eWDhOY6UwxnRflM9z5aTH6+cBVhfqIV4LfsaSvYP4lUoS29QEdKMDujL1
wG16Q4qHktYeSstn5LjCYVBbJDVhNBqgQ2PZ068/VOuJkoof+d+dlY5ORJ7zPQEO
HxZ20I7O39kyWhSeponnZ0FeHZzHzE3JixEx/VpIcLht1BuSuRszm7Otrrow1cWS
hDVnj/cScLzzVk73ll+4AiY7ZZo6332Og8f+hRYyrPgq9zUCqjas+pRSTGwAEQTz
1cF3qC+N8izHvFxtLLxxwTlBfbD/QBrbQUPu6rZQIbPdYcNcrwwRFm2I6gGEiBF+
2W+9uuJZ56VMzg/QFi1fxXOxMOrbq/slFXvrf1Z3SS2DBZqsaEVcc/Zve3O32yO3
Llk7/UnLvE55r8cr+z0/oiJVmLFgRAX5+z5Kc4baFt3LETXjtzY3Y9jghF0039Bm
uRVdzS/te3rexGLgDwo2VD+6VielCFczjhn/g9O3Aaqo/R6mprGCWVb9E0B4bZt5
i9pzWBzRXi7PtGFT3ipCWzuHEy0PdfIvRiQk/A/izAPimHO0sN2OCR6eSc2NX0Pb
Qjz38LZlIS/lA4fFsnwyAl7LOUIG5Spof4X5mFitxGeXQiY8goM6O4q/bel5jzk5
j7V/1n88eGkiQrfHyWTA1w+myeJ+0MaTCM87Lkh6d6tOKTz9B+6xqU3pVDKG2Ihd
Rr3AWmXah6Qforo2TaoDaDfqtZ7YTKywMzpKT4o7zMSG6TbQhYVa6zmhGBkVEVwV
+UaEyqVmQe/yWx6euCFid+6cqeIaq0br/uPeElgId/qY8OYZoqsspRyoNBJn5yXn
2XzGxHHhqU1fekiD2aGuipSYsMeD7mt9BPyHM5B7/eznonSWSlWD+QVylF4c750F
g1T7enp1Ap3CabN7EDvgbcTUiKIMC+p+zrbgllhRumfzq5/c6zPXVTZkGL/w8rLN
Gt+9zA1vO4FL1ahos9T3iZ6bmGMH/ez8WUagNqhwRgy4aQZKk6OUIKj2CWNm8C5O
lU6ISITXD8OFbzlzkfL3P+0L19PPaA/iv/yV8W3DQTbfbqrbF1ywNkibk3IYAITd
azo6oJBhY9lbc3IwPDd2CPMG4swOSL9Ui4VERSm70xhHGANvvrxwMhrS+Fx43Nfr
snmUQEeh9A4t4jJMoM3yEufbJgHZlIarH+3MCbOG4VZ5YDghr1DM+Gyku/RRbodV
/O2Kxq/7MKw2+tlwCtwAHHPr+RrJPJ2OQYV+FYZIQ22Xoig3oXI/JFHOhEEzU55W
bOw7V0Xy1miGX/puniF+zUuhA7NeMBYBF7fZrwqF4KRhQfA1jRnshp8k/4vfepGw
FseVnpYZCHI1KZQXpKYG+qXpivkWOER5JXEq1+Z6XlG+vs6BtO3WppUxMxhf5aPP
Tvj+vOZ01h8gVqbupS3mVBoEOLtZGpDUpgh3ozk83iZ9wVzi5pxst1vd90Bfqvkl
nay78QGDGQLogCoexjaWPercoXP45Rjgkb7r1sE8b3j84M7BooarBvTRQ3mSNt6a
c11BySp2AfOQU1hCl0S8n5fSNJwBo1fI6dh+x3/pMiEiH+UpasIgc5vjwZ5q6wjW
r5TCZVdkef0QKFXRRuS2HBTop9FYQnnUD9d4ISIlFfWCcs+gKVEnWHoH1Q341cpg
0A8eXnDuubZ0IeRdID0Wv80oIF3yEKDWxd4/K4j7QgVxCe34ywT2uD4lUyIVXxsr
JxEf7dhagDwPApuKBbXWyeJQC1hX7/h05ULxc67B6fUdZ0oHAGWv0ftOPirjY2Fi
ja59dy9tge81cJJFh4yziXK8IeZLWmdGENshXQP8RQN+kaHUyqOT9VhrRbUEz+p3
dJT2bYCRksBINLpOLzKx4YwRT6hZboWPzSdLtDQuTmlWmYndh3u2otnXiYj/6B6T
XjSBCWPuVb4oBjlmN5J17CiO9uroN2Ia49tKvtzjgMmm/zUxjQu7YFDjDodYixUb
DUgM+vndNdFhMA1mlJgdF4dfc7KLG7IDp6pnVTKDngIVfek2sUbcJQGddLI59r7f
FsOsBXHckX+ku88tkhiOB8PAtQS0u6bCoTBxUKA2w2LMlN2XvhIzj26bSFYVPUpA
cpWERQKDOyTUO4Kl069mW0XYKONRINNVqLveYp6LI+FHBHbmoq/hnqAC0ekCGYpr
ejEytwluvMAgoLbDW7+nOnUaAmMhaUpg4puLxnjZfdzjLpCMhMd3iTH2zGIH+UoP
LbN7jmsjLo4mo/+B3LuTqQ3RF0cBm8uhdFMkYqbswlmYdiGNFiW+dVz8zRrL3aJx
YYZZ30mTRtCNvkVNCT13udfqq1IY37pIPAd0eVOdaAFS1Ai8etelPnm3ltniHGQn
5pje0jgc5km1pcfy4xGy/ZdKirTEriuFP2Wu98kSHs45pai3kK5OXnYkiDzdl/ch
slhPTwGb/7UEFfa4N0qXqCPaLWSUUxZ/v9irkdG9c9SnVT57ZX6AaD+Tc0V/MLBb
od86wNaOZJENwUr2HppryMdw5fcLdnr9kmYH9UPQN0zpdGrao+Y/V3TJQZroHZX2
HaZq1ow2A/1DXkNA+nshFamKNfpOeX836N4rrV64UgXXIqWCq8ST6LxZ9LRXdYP2
mjN/L3p7/j8IBm9pKK07iruy1IMMSGh5tSie2ZUyOyMHxzTB/0is2O49U0EAUgZn
ynI5v/9+/D/0D6RO4mJbLgCboS9s5G8ur+QAYQN4Gex56HgvP1m1DuwCG9nkf0Sa
fXMu4alhF/c49hJ0YIVZ8ibbnrlh8jepujTuiQqxaLpkDbRO9IWMdbIO4VLMP0NU
EpbNH6nPiGeS/Ft/ITQBGI7KtT90arUueh/eU3Wwawhd0hbIizNZhHS6MFj84UXp
tfq5zdla8nOD2FvGpNz1RHbX4NggX45A/1gdCxottxd52jdTsUKxPyTFtc7AIbzD
FadJX4DJvHYpqCNIGz2uQ/krD0IgmMkZc64213FdvldpGZwo2zYb90N3NGIEGLs6
l7DBeRiz9DcKo30cO44LLQyebTKbkzr6vh+DIjIGIQpl2/RoUKV2wHS6ZpmwKmw2
71LBT8godTLZ7R8u0RAuzLwIi4BT9VvHSIThqIapEVghXTI9SokORPq29aDu7lS8
SjfpIvdCOpTk5cLfbgVYUUNSfuW+RlU0+CMqlIhKof2n3UwPiGnyFsoD2nTRtnX9
USodfSrkk34F34c1Hd9Yvb+pFHmK8Z3dZ3YYUsU8rggJD9jVbPpjDmBA3ZXBD3uy
8TYBSE+wK7OKPIHDHAU8d5iVjQbKghp4wlh8SmrbVaO9EtkOOpgUZxjwwkn2jgGT
XmwM2j4pLNhdEnPQ+QEUCqDHgon30o0td/nAmcAl1zmGLDqC99/eoph/N0daIOJy
SdHCYGkLWvSEt5xygGTyxA1E9zlYGylNzUa4NmHx+D0hkVzA3WQ8TItPZTkUljnO
jo+AhprlcDxiI2ACgBahE1hQ7AJumf64O9SHZPeAxXU+EF3LH1PxpeS/aFXSK61B
Bw27nByVfJsPKiesLNrL2EZ344WSTYSzALp7G8SMupivmVWC0UBQNWwhtxL0mIo8
WdW2zaWaETB4B96i+OA2wElc+Ub4oba5Amc7GgMVe2QoGz+0UvZCR158jeLW0AGP
wnvv9dS4eRO7xH4siKIPMQEHOt4ggg8ASV7i5I4orn17YsSRMYaVt5w3hd1ukLes
1Ottk1x+KWeqQqpHZ/K+egbPjlC+9SOEU6g0ucpcDoQej4RxcRBDet+Ib5WbGT5f
ceY6phTx3E6l4GBz5Iat6f3MKcmXbmzUYVlRsnphUPfghDPzOT6tQL8q8l5l4MAZ
ShX6bmOdrmciVqU4wi7mkDGiJt/PyjwHYvLgERmLHmUr+n4kDmnRdNsu6QH5Pq7B
B+vx0eu80ijs0yTw35rhlrbPv5upGEE1z3NdsQKxDwot2iAVUxQGELRA+woGWgKS
C0U5wQf3lGaZDsxk2u4rqgJQCgJO5T029uH9tPBSwI5Q+AUBuybfYz6/Fs/KgdAq
0F7jr4SwjWvWj1lQD4grQsQ2Ny3UjQ/KVPOy2Zq6VYOV09781Heuj0tDz4UjvI8G
kCnuZSdfanMY4/900ivalsA1Oozspxbu3OOPAtT6+Lpu3eFuE/IRpPiVu03yb2IY
YKv7Fwh2ZyYQtzBGzLAJabOQEpPi/Qo13t5oGE8K0UskQhPXVfAJNygABOZPMz5U
793qjwRw/amMAminl97iIItvp90nOS1Kye7dHsTwTqPAqTbbMsKO+XesjWL06t7+
14OZo+zuIvZcwUMmJ6poKEXopjIpHgd/dNOiUzFwzrqGw2d0hfLJVMJrkHeQtcnc
yrLpI0LzAxv+InQyhyC+Q6cXxIh3p7DbPjs2VsH+Toagca10TJuzEBr9XC/7J5h2
goDb3811oB6mrSJ6QAttBk7LEVqAVPrTfELfdIq4KOpA08wZmMPDW61Owm3wAdWB
Er3xWgDbjA0spIEz9o1prInxVsY05nUcI2DnKHIdZPemkwQutwBsNhYnx7IulL/p
Lae0jJKh7u7bNhFf3/Owr0lM6kTAEEwi5TWbZnZEFmNvpPOs3pi+aYw1apqevSlR
tAAJV8O4ZplO2FfOOmMY8XfUQG+zVFgiX98nOU6mbBt32hRfNZoMomBbRYySgw6J
Gs4BSBbZCSJsAzNDsByPTc13oMoZNsgH9M7Yf7VrfYL+BrDp/ul+u4BL93Usz2to
xtsLvAb+EJ55knp8chXLKoJW4JPyUyt67iRC3/qB+dc+C02lBAuLoToJVtAnwukJ
3j22FQIML99iCkM290/IKyY1hNEw2uHxJ3ETFPjfNDAaX+rGAaF11uj2XKBqtq9B
xiCx/ss1hyMs5ChlA7VVmXqQHMbN6po3pZ+2wN5WJFDwV9k9JaYHO8/7kFvwLhbG
KrtsQnAVAcP6NRQhHq1gwkFJONv7mIAQSS11vHtu1Cj6XcyNiGTiXgrHO1poywY3
Olmm78Pg6Sj6r84g/z5SmQF1AL14yie5/13g4uzYrDxKgcisXpRJCatothCqhFfg
ujKr172ExeSzEIpCTvS8XwSnmcUhArnuiaBYFHraePLOCr5IVU6B5KNoJFmub8N8
21KTv1vNUfj8sbyoND4Fes699lpAfB3wY8gmVemh8DOac/BbERHEZomxpZ5cQTPP
J/NrEyfg7+QnjrBMOvIO8XBkzdrhLLWnoSNo3an7nMGCpeNDF2jNpPfFFLHk2wHa
zYlzvhy7YlKj/umPaEJktfZ99t0kL7Zxs9aVMaiipjZTlt7/6A3Qoj9oM0T8p2IL
UrYfI1JMTtnjBIAoTZp/WDa01+WXaZN3CSUgcRzpxjGZolqzFjkXfW7TIFFPZNvF
48vf4izOJ631+BNUP9j12opQ9I3UwDKgulsw7lL6bMnj3Tk4jKmWSHU+FRXIdNPH
/NTIoY9u5a/tZzcbU5fPhq9vEmbBNlJ8vP8cqQeHE6wde17JiwmNAZUbhzaJE2MJ
0/SBlFKeT0tuOGs9sC2YyL3NYkDUrzZk0nf7nvCIwtqsm4ClMT760feKMDypIu8l
R+UDf30iVru4GDNwccDVV46Bf4baHqNXZuS0+wyupbIMYPY6JX78A705voeWWC9K
AojBnRCqbp15dmfDJWzJ3pQK8HVwlq/b3gfRA3AA2ubXDYSNqb71qu13JGy6r56H
j8rW6c/InqtzbnOX1IEzncRHdwKHTOUSejgPzRKTvBsdW05dQcLza0ox+ZF0Cn0X
wdMhP6d2iVdUUSfQOTQkvF4KXOZ8yaq/TeGu3y1vdDabQWI0SdhiyIEJIL8tMwzO
L2ZFJuxEDqIfHlC6559Ii2O7wPC1voZEDpbHISZghY+2TH9ANRhgKoCfQz58KP1h
hcW06f/OiuRmio3923TPHq6ALuggCB0OdGfw6kEbDZnrz76jUfnkUtiGDHtgzjBE
ktZMOIpWcPhI81rq5BFJJvqxTRvq+WskdbM/niUtimrNYbsNY1FbkdzbdBt00cYa
X1b9GoPYioSd/J7c/lN3oamrmhdqCybuUmf3EozY+6nObVI81GBahcakwQ/cLQqu
hU5389qqazs1cTaJHoEf5SLTtJV3uzYZyKuskak5H0u/iIf45G3A0l7Poqv3QVLI
UiWeYeUkcIAfMhDaD+ZMBFSozp4nv8ITKBYSTMJZAjgCrogYpeCDHDPL3V9RFkPu
B+e1nyqsU8qO5XA0ocNonuadaOFVZORzqHPOi4K+7fNS+e2ucgF0f8NXZeR1h1zj
k7Zp0wSug3c2FelsHFHA7rjyGtqHJY4kupNG4NoDPPM2kHzZ06GlO8EQGHreUUT1
llbG6A37z5jhutnJBx7Mc3NYT8LN6P9jF6KlYrTDuUA1WlqgKJwVI02/X2nIuP7+
LYD77GvTZ63NqQ1h9PEe2E3+P+I5lNP6wIZR5NV+PHno8s/xNgOo0JtgbsbSJgKq
vmNkG0a19vFI+9ynuSIJ/yB1FYli6aDVXllTQ1BDUniEMAMs+0GOoBpELG1+A0ho
OrChLWM13/6xvr5cgsfZrP9ataQI0/3fTSbk15lfyeaRKW/BxD9v5bUmX6UWDt1t
Nqj1SVJPLmepRzAXDuFXCerPjB7rotw8xsx/6iu6nAOdjiU4BGXsn2uiHgqybFCA
hQXKODCXEeqNZeMdXLFAqMVK1wOyBLkuf25lhzWGaXaPUIQly3c2177QjHRs0NCS
JtNAtqba5t9NeYXehrhAGsPTUxyjPuRtvF9r6V7p6BcYDnUPTPvUr856/Bago4Os
mAGf6Al4utK2rgOYlfxmNTnLowQoQYkq12EeuUXR9IaYE/+X1uLJ2Ap+/I3PfFkE
YP3j3n1cixu06+HUsL+E3Fn8Qk017dKzpEJB/z1M+vqviSLkZEqNPlR2VNHt62DI
T8LmH0Tet7k/yhLIm3rSpS4C4jF5JwKFRZCA3hRRF8Itq1d8GvzJIDulpMiOH8MO
/vSKUXW4JR2LCZ17+DR6DQs97lpkAexU9pg5jWLmkTXPg6eqbVruQZ0lZBB7b07N
dEZlYz47G76jEQWaUbv7p4tkqA6H1RcTvrQs5VynIct5121CN47eAPQ+hQcZH1u2
ZThzPL2N4sw+iVf03qV+LISO5Xc5cZnqy9KVuUcc+hwfji98Dg82KUjd+s0OwKzO
GD/Ya05rxZbZg0XfNYglSM8Kj7KX9+XbSuIWd7fFfiy9m1ylcnHN+vwqE6Cqd3vE
ZAIo3JBaRlSvLm67cXpAmDovN5qN05ljWLz42NxUpqjaUWe7oDWjogX4IQ+dMDfY
i6XRaySNunV7T3ftOFg94tRo1XRPwJIg4f071XwDdPHp1IjEEzZeJQi6F7YFebg4
pm2R93oMQSLgfk1E71zNRyTbv3cODFZx88exXMGK4ytDD0xrfknsGyg+VVuvPSof
PCPAuEPCSoRPNB6BCM+JgwDLkGzpTkIm9KGlaLed6D/j5c3PyoHyFpmLUOSJkgYb
dTOVF4FwJ2W0GKSrLhFuasMjCUZFDxaBvkSeB8VrO7P3+HuEnURWvwlT/pTl9xda
PJZjMzQBvHZDF7uxHZZ/MnyqubRZ4pS7r4JvuTKXY+r+Ha6KteJqjYKh1O4P9WMh
gG9ZPpaLv7mXqlnciZtrvRKsX9VD/HK33rPE4eZsqwvJW2HOkXXUVgbANgKW8q/C
+T+JGDrOlMT7AduUt7wwvzj3Cf+j7Z4oK7+PtEPbbIB7zbHqXCvONotyRiYPEnDK
wncQl/6m2HWBwYPSivZkViSB6Jof4wlp+Rljj3JnaogWnIUifkVwhCVzPPvhuAOm
zMB9mgkOtZMB0eKNNO7PRIgWLgKS1mj9Qxmq6uyflru+Xc+k3aIaKHhWscw+aa9W
J9+c5ktjquCeJxmqrgK59jV6gwtCjO1mA0LxuFhmRmy4vXgu6rEMOS+rj8G9ICBx
BU2Vru0TIRh/EOv8TzB1l8D5hTsTAPFyfng2F/CXq8uPZ7Nk0MMSjbqVZEipNzL4
nq17l53aO6FF9e64ulMvwTWKAluBh5ENn9ovQtXIB/nUYFO1myo9qVmG3hFXI9Ar
QZF96IpmTlCauzbxy646hETmgKEE0RInDygvyXH9oY3U9I9y7unmLz8ni6zuRZ+F
5IuAYyavEdyDci8UnJ3wgpSb5pdgBbb/VXAyP10U8Ws/PJRknR0/wGj/tW+AVSQI
3qatGHURAYa3cGVMTj/lWWf3fwg8oFD00kQLbxjpSPGqWmwJ4XQDtCIS3jTSJsIR
l8+8HZ+UeRIrTgbzBrc3eFHY1UVpYMPQ/l2IZ9dh8KgOflW3pE5z6+WIEXa92LEB
xoAcNrZ56fO+wjqWLScBxVLOGBEyvAwWWoO4eLrEl3TRnh9zX1hzJCG+qpdp5unb
gpEDoBEH+jCktEwC6sdCSCSOVjMevuqEcjfBlQNnOkKVxdzCSOYbWrmqCkDV5umu
ryF6DhyaTNWBlBg8F3b3YMYyfQa8JKIjeNER4ShigMq3SfcuCT37iJaUJfAUqWU+
SltPkBxHSb/QzjDp+Pcl2eu8vUABqUVLVq706FVZ/HeWkYQWPphwwAwiw1RD2MXa
XxD/Zqi3u+GjwOsQJNgNIb5X1IEk7eidlk20yxoerL0Tib2iTPQFAOHeQQs9sWAm
1IMgh5lMwpkwj0smCVuNdR3fI99mjSdKII5GChPpE+sK033AoA4Q82gbn429ej5q
snhBAmWMceBuOZpEi4xBNlGxEs+cu+w9HQj7eRdkel9ivMT17zUc/RDIij4162c4
dS63aedeTP2RwrFJrB1uBt7jDuEw3H/2T3kPY9HkNCqfR7Yw0HDBof4+2yztJTfW
CW5ZjvmsJIb8FiEE6/n9nYju43bFMVz9kb64ABapdwwMRTP6/6Z6Jp2VBbTO2PD8
DbZsjZ91O+L+Wi0Xshm70oJjNgwFHVscM8XEP9xdwsP8ee4mdDFsM6DJDFXVFxbV
UnkbDZxpVL/I44QQyFzcguqdpxK7l9KH5MqanH5xUh/hHqAicG/fQyCPEQerjUfs
0ilpKLglND8J4rdFon94blrCvfurkjVUKEgiuFuEiM0TIkp2Bi0bg4C9e8evDlsv
8g/ryoufQj6ntMAgcQ9LZPA1R/ylSUQD9N1nOpA04yshm/gz0PZX3j0ENWBmhPXT
dK2wTh/N9mMB01wns6PoDV8bxZsBPjCnm91FM2t549Khu9GYy4mn0CYjn77BjFbc
tx306vpLC5xGeB1FbaK7K11ixGY5AdpiopYm1tajWkfg+YgoeOL6754lM8eMpLEi
Eywx3+1FSvl7r1OlGTwW9nLALBx0H2EqrqWTl0HhZmB/VP2g0p2zTsLarxF8jl0x
Il2AbZLxPwgBFCXxHnl8siZVYqHyxhJczpIe3DsBALr1vqAKxIuf8+PE0QtW2fS4
CotBAM3u5cXUebJYz+mhxkNP/ad8eWwPlGZkHgAq8sYVZGJI93yRC24cCr7S0y3O
vmZYqkquRX+BjeWvK7vTtdij4cS06npwzDe7ygNwWldRtMc4ibUXoiG3wKg7LUNY
k4SYFeSmqp41QAT8CV5d0ZFkvN4rPli0gq2C8qXnmue9w4+mca5kl5PkPMPTGp4Z
YBlgJnqlSGA0Pvul0LPR90esX3X+Ddk75BCvw9U6+tQ7WI754f7/BOGqviszlp6M
ayBSBkRrDN5KFPNV/Oum4xFYlDJLVevtKAuwYDh975l6yOtxma+ZGJ/9Yw6IUR+B
zwTu8k9zqlKbUb6lyWDQT2+LLaqWnRn0DMl9pwNv8EFF1/KT02WTzvJL2UgmxrKk
XzO/Evgm+YWL9EVeN4mCcLMVaMzCPMc6nozXBBOg925rUThArQyj3OnQpHJHbxNb
bWVRVWsslMEOSBbsjAeET/TEjHjJaY0izN00boYSLDtElKFQ0Czv3COa8iqRxY/7
LhCTesY0MA9h/5HyVQp+ubhsrmlauUGRmY0KUoHWqDIdIaq2hfSh2Wxm0P4lr3zj
3+ETDxqfBJCKGe+8PIgiltgWn7VspgiK++P4DgrX/s8ZVb6NAV7XljObHyNp4v5X
rJckme0AbGRTFV6jH5zV8mKSCKvLh2qalTWRgkoT3UQNFSWqiPxMJNfjHxbmwd8F
6g/d1wMCMvz7uOrZTxxy47yo6ECngF/hXctIe3yN+8WpV210ZYp2qwgao+XtSoCD
UE9yUz8+wYgRK0w7eNtVfbG4XHTWRWy11hZkXJkdrtjWHrsVUnwLD2loDS5r9L8d
sQ5BS46Cl1raUCCNL6XXWWpuzqrPth9NglGQxoHFxa09T4sujDvClgFNpgtmRWNC
JEVvFjLL8rzzxqT34/rIfkEug0+Sl677n249DtlJQOhdtyzJYEAR6Ov/KjdWIViq
9kY9QoaAOG4AonkHx5S0LWR4kV4J/xvV2FlBx2hOgBzGsK+r0ueWGa63m3cU6ykv
f/d8CUsHXTNnPclO0QEAehRQHIXYi9moTLlQxkhhwqIId8lRYwyD8TYz8vgvuRr3
2tHADaZ7l8XudTeqZvpOp2zKEbSaD219jLKhjqRxEIjPSjp16Fv6qeCAaiNTJCOQ
pwxKhL2U1bB3qXyeEKoxQHZ0itHx9jq+3ONnHNPD1tFP3Unav3AMMudwJI1jGM2t
+JZJXUKL4tTnaDBIrb7MWYxfJS4sv+cNwzDkL7A+XBoZCmNCWBx1QsUZ3skc47SL
JG3K1M7rDKWNNpAMHmb//WptFoiQO2yioGb07DuZRIeTwsVaIhhCVLaNhFCaSlC7
Ihg1BEu0bce3F8c8Idxkcpqb8uH/ZX7cQJX7s4Y/f6M5H1JSMH4hiLZJrxkj37lv
8GtnjgEm0egX4zsg2xiHmxSFwHnyj6qAJZGFHbyAXgWGdhugSaUM6PlcTQl4Ty41
yiMLNNtw8c/loNy/XHAGIpebXj1+L259tODEoAvW6tGlP1H8iS7M5fb+tAhMSAbB
eJafXBlcGub+jVrAlo5cDeI3cNo6m8z7gViE43MNKD0SQS777CZU3XtRUxtbUr7/
NsF2wIxfssAW9Zo4ie+3yIRj5JgVodVpdBK8G+gdVxZeTiaFYb5KumaWTuF48JNd
BSH3++ujcNO2wSIVl6e5RzyVM2s2CdUbvCc0vZbUd0aMtVvByV7ejAq+lliZ3mK+
hQAK3eoirgUY7t+tXl1Xm4SgPgG6AKIzqqYwSDVgPMth/q600xnmIFpI+LK0hvNb
y9pYEbFikWN8xn+5bYsXXlVA/mtOERoCXqhyzgbetmhdN6xaf1JuhqehbMP706CC
lKytBRGBixG52Yvi3kJ33BfOEu2DGimxfjV6/r25sR5NtT8EHBVO7DxkrcaxMLdB
NqHAzbr8mZDzmXb4Y90/r3OIJ/xRBmo2Jw73/OHISjUPvy1gkZ8a0mwooC494IAi
sh6jmjUlIp2lu4Z+/3SBnqUKJ6LPKycx4tmh5n5MbARn0KmfbC+zWs2CThfJ+D/P
SsCnfgcXaESjcH14q4Pfn6celvvBjYi/L9MBVNVw2y1vvmqwZgfGwAXJAOokAI8m
keG0sfMhmBh4tscjavx/M6G7oTHDS2k/ZkMW+evgXn/+lZ+ESp3YjMbtJmgAOpKu
TpQw7U5Qk0CeMvkAGjKKd8Ik6ZtJVJM7yI9jUGQ4lVHqrq2pGGJJFrBC1piPX1VF
J4mTkLpgziC1e63WbYpMEoEsTsJFKy9+v3Bw4Qxgsj6tnYzaO7nCX3bb9kj4Z8Kl
My0gPkE0+xMN9+05h9sGAIzYwr0QfvqUZfeW2g0T59bCzjm1kHqSphD5zsVBbh6d
MoyFqXlrONZWHAPd3v0vsE6RaYdhCNydYz5Q84m1zfFYg9U7saMb33tJ+5lukX3X
j5PBlImNSW7xQ/M+ATvCkeC2BAWsnkeZxm/Pr9403wgzt0Ud86EVnLcc0XhRbMj+
dv4RaJWbxajSk695IpLGDGAKTeUAkwGKrTVBQDSy58jQrZTU5QZCgCeHCvs8skWz
e3AiPSqBT9oS0NLAEdyvgOCmKUo04T7IHAa8ikKyGrGbDbsggi1gCpVoBdeXOE49
QgWd0qwCtxrlese7NcLyNXi24951irz0PdFp9yMSnyt3y0gFCeKpcdpgtRAvEofS
dFq1mp0fp6nTcIzuFYT+/1XO+qNO8ia51WG6Co+1RFk5x6xkIYHMAu1sAjiEElLh
C678glt/KWOE5C96XfdtQd4tO8Q6obAjrN3f+LL1PpS6Gfjbl2STJSn/ahDlZrDp
19HkYKtIaIguo2yB7uEqYwPMtqCbm89Z9dFGUSbo3+DDNg1zGD81iTHpjyrTWn9y
3SPjV0/uonGuaK7TKLG4XthpqpwVQJz82HJhcZdbF3fDMAW1rkZsxm/kVaQrX1Re
kpLdQr0ZFULs5IOUHk8pK1xc67qri1JwGDM2fh9VTLqIGyhu9KgW+w/4owjLpYUO
Y/hk5hAK4AmLtIW2LT4Dnz7fQT6e1tekQ+qzs+1gn8R4qcK9FGlO/Bee0e7OBlSF
N/m7foMteg836Twheaz3lHt21l6QQRHqEZAkjbl9ob5eOhbFSzplUIfUUgciAkxH
D816PLLdUOVv8ydINPD9sUclLGz+lIpIFsGq9apvRic6FF6d9U5jDFfHZxnMM03q
KOuDHh3PVoiS5dCVBTfzTJos+CayVOtBiTR1LOfLjwwruTZbEld/XNogBs8GzjmC
Pdj7FA9PPe01qQlxsZ1BlfGEfHLPkbxrudnvZYclxLbzZNxgMsy8HVrhGyfOVv3a
26IzFI6yJ7vBOxDsHJMdykXPdvFaRBOkpx4pFG4N4NkBFsegd3CfKaamiWYgqOMw
3ooy6GWmH5RRcj7JyQ2Rizv6Q3Aip/AJHCkF2in0PD11ort993RtWjpuLk7h7IyS
iwfaDO1leQao38v5e4H8jYWdyGQF5U+hvtVr0znYCjktEDyAPpWGmiDRf0fYTIYm
259IIEopy4QC6gpl7K4xKH0a2SIBeNrmO98OfqF1MRvTLOemretjQthxB2yunt3t
gl6tFlz4+65qknus4/iZBa7qlqIwoGymWuWWwb4IXiSKVKJ9unBh/IwBmfa7Et3M
VmhYz38/3GiZSl/6blc7bNeGdygXaOsgcIEFCeXjJWc2VvaBItjE1SPbu+u/Uxp1
7JPuSU/Re5m5uYifLMohMVWsrd9P9B9yRKRwg5xgfb7wL/uSIdeJSKiSF1W1oSSX
D595DmeTQ+GKiRmxrwwsoqkU+gPd8bN6iAJ3pTlZi56rqhqppbs1IUxouqBemYAk
+juCrcg+cSO0hBTj1R5iqc4k9b66KdYzbBKY0IVL7QyzyhZABha+a1aLCtkJTn+n
kdFwVb9L6VvFnWYPdl6uT3ZuQwMYaVk8vMeTwgVyxYObaPNX27gdlL6hY8BBz+ao
lAsOV68MK5GJHqLjNLppC7v++creC+7bmFre7cfVWOFwfCHJBrmZ6qUE7yRogLG7
2lJF7d67mais5VCvglsNeOrwn33X7fTzaWl3GYFxH+YDmqWI/HJpVW3biEPtmV7u
Btbau6T63dqLwBsqkV7gSPQbj3Z5+e/p+8Wts/5VDXLlFi3MLBLUDBlXj0kV+Pmr
N7S9b6w3ORvE7cwd0p306SVQ4gNPrRhQtiMTX7fEf77/YjTtI4iBsdehyXfYC59d
3WcyJsUFMLR5DKrc5tOwjsKx7ir9vVsykWNfmvTUmbQQJDAvUrPWCrv8y1P26ozm
oosEbgFxpbnjhZN3JnyWjCPZh5T5Ekhl8fCS1UZkdZ66h3Grdc4LCtO3+FIDXOdE
elItHtQf7qBX1tmoS3O9eakKy7orv8Iy4F3ODYbNOAJ8mdXrT8+hsdZJdk/IRhgC
iBeUdC1fNS9gJWxTBRrkELFSu4fg6SWtaapNrjX3UqWybSUZH6bYVV1ngeWReyYI
xYDCx4Zt02G0bGTTMugzrNW1Ae43OgANAYKiBc5Ie9T2HWOS+D9OBY16wA2OSR4f
6dRKmkuQLh2ocWDW73T3fRpX4FXTnvjgV87I1QXYOT1jdpXOV4wtqewiMgpln3dK
xhJNP32LTh68WnONHHGKHnhTvyG0N8KXCXADjHHudb/2V7RPnNHzW8qC7pT8LQ/L
OrqddvtzMJCbopKFLicU+nVifdWbaUmGFQ6CzJwxPpWEP7q9BAsZneotG2oMRXna
ZUXsI8AP2IQjUbS8lRqOBV7Y2NXqaDjs20Yekq+bfcC7iWVXaqPMCBr0PFlFZcxl
r+zfINR50voHDdYESJIMs0WZ8AN35zdKcfzz2up5b1cVrj3JE2B3w5aETVCDbkc+
y+ANc84YRCteC6rS5CU0u5JBzaaRNASLU/97/bAXSrS54/fQqQdyf/0T6XfirJty
JgMt6+hv237GlEeT+VsVJfdb9pjWZEBBwT8CCdns+BXm02ndIYqMxyE3arBKJ1MD
6LgPhkX/9ZpRS0iOwO2SD2HpkHnmLcJA4C1QDv0xwTr+ob8dHP4cSoAuAB8eqclT
+ISAlcC1TWFY9c11Js2xHUDf2Cc5v3R2574Je0J5/1T4gpkcNc2tmrgzIJiMhuZe
cGuyRdyKoP5Q1klYsaR8p1562mT5RG8zIvgXlwyL+78bY4/mLY6TKTKJsDk5KctP
tIaHg3w9HnLAkgJLtAX0IZ9YIltmOz3ejxZAvG7GrO563LRHKiWlo3EGTArNYp+r
mcI8vMj2mIlz9V2k1IDLP96OUaNDo8s89ulMvSiKgTIzATgcNJ90O4j7wjDyehO/
XEBvGRPPeGjjEHgV2NVyU2UiYbJuR830f33Iia5s/TrWuiWOhpEwKXGHjVPG22eO
2y0IOfQtnWNN2eBcMuKlge5K9jd6H4BfHQhR93k8ocCQuviQYm3PcoxJhaz9nAjB
mFi259Usvxxt55U0Wa+n7FrDr7+0JrjMWXqoVH4qWJmRXw+BOrmU1ME0YMrfueNs
LxSzClSNZGxB0GV3YFGS6RBXfh76SSQua7s6iBr1S2pnJEPR5AIPkswuroY0Zmkm
zJ4v0ZyOF7mtVgTF5iWUZRdajGSRv8lus6IC+hbgz3E05qLa9SAIN04dC0jGGU4F
i8Ixj52SCsh/HA+Vgwe3EJEoUdBmJigMGYnp/wnWhN8sOy+ECFpZyE8VR5jOS9iL
yecsdzJKUWmvZQvgMf+vBsk0qVLv0fgn/4UcPLoaQyy/NATaDNsnLt4RITmf202D
34C/HMpaCE0DI0SFYbK++ml+R4yQKbMSw30xEjcfarkQuNZiNsTlNAMMybkMY9x6
bYqvDDHskBWtx3Y7uPSDpC+LrRGHgZ/xPR2ppuizO8mqa70eRrS4Q42KVNE63nts
F07CN2iz2w8vIVV4cxEn22epKohSeKd/4PLjf5NF5KdJDcfyOyXb9Kf//o5Obs7h
KzRT08F+biv4Ud+DeFsV91JrZ7Po/ecFce0R8uP+65w0nokouEoiXJHlepC05aAz
RpWYWSXfBL6Zb2VrYDpmpuhcdvKUsy/3XNnL0ff8vxnymRKL/YeZ0j+/wrxuvc/o
ruUyii5jkVDKXrxclYRumQj6kIC1J2IBSHbT4oqQvS45QZOP2rYDIKBvLZOAZIrd
BlbVW1lZ4VnPnvq57kgfNRcj2Ho32HfPFp/+yMkOCmWQuDjaONKBLvJoD0JTNTrU
+I5Y3vg+gyql6SPVyA0PRoW4ye4y0B4gmctFpbRS0DxooMgYo84jplcz0vG1xQ3F
Hxq06VzoAL6SdtpRPDNNNmctRd6bS0UzE7keK/d+mnmCehgcHsChosMBnANEcLwH
gtNk/c6Jfg2SLoQH7gklOpy3EQ+fm2BMv5MhRWDesaq4IvHVPROo+Njaiqu2KUkq
otz63BrM1m/LNTO+dDb3h6RRmS6hMCvFcuaRRxHvICAzpP6tv/qK9wEXfI6HObgP
J8K3h+VWaQGGnVJZOSVxIqoW3K314Bby2Fl64+KVVkp/+Qbm5HSt6AVqEJ37dqNN
6ZoWxCyDBXFsXOR8zThwdC6qU53fvkS5/4Nd41M5t9ejPP/Qumw79UGOWoUTGrxF
2K5+ZEngBKOonPMQOBXRcdA2wdQahRz9X5o4KcUydmDhlji2Ls6pBRrmkPOHysWe
eyq3Y5nqWAb71IoLagdbqb6sSDxQPEAhcGQhH/B6cB5T/FvNPdIw7hJ87PKlcxPm
BIyCs0tm3Zo9OgMgWf09fiJevskDN+NYzJjbCn/al26mLzYSTU47I8pDcY2UuKKC
ZVOJLY6z/r8eZ1dFqQQWVkF1UEZca/6dpypE8A4lKQsM1QSgwCQIDSW1vVzOyU8U
FXTBMFbfziW6PRRFzkUFF1ldp6BaD55CbpnqlcZrhYwm/aAjKql5L9057s/R01Vs
t070G3B+h5fV1NieehSgBh0lrgjV7CUWDC/cnETSbpMD1Ku5DQvCTLrYfEuQ/Pbk
IUa8csD9TejvKqpFpd1PXIsC1wYw1sq5hmRw7u/R3cxSHtifoMvV7rus8RPnZ9KM
FA1vafkj5okY6RXBXfZyjpdCXAEyy8/Y1iV9hh7pmgTOT9TfaCjNvlofT/al/2oz
YF31eH9MeL5cgvAq+w+5Mb9b1/HpurFgiqtRvOgiv8DA2recFqkS6QIzW3J80TjA
CNYsZkIJbdq+wHnwqrAC4J04adMzOQPlz2ik62VPJdzRe8A+aKpEXLkJ3PcL56L4
Bd6n6CRd3i2Xmq8VyGljjgfJISDeGElzQDrjh2VzEHvDapT35HeXsNreOwKiL5jy
w9GGiI2Ajsy1POfnpD1/DrEZjbfh+O8UTNz6olTfqSu5sc/T/5D52w1B79AI+IH/
XLVOgL7E++LdRBznuIabj/UeP6k4GNaJd9PTMdTHlszV2kuUgSwGzAYCBEQqYfJ5
VDiaiTPQ0xo0F3s/jSyo+GGB7Cq4Mi62DzxjAb08fcqtQVJrwlKxl5d0V6z8agBw
U5tBhYBS3gUPYgCcpCKTs02x7EtqNauBC03vxc2V6ILFCyJy73lUNmDHxHe6opB3
u/yWPVONIEwqtYXdUTnM9D+82rNXvI6Tx5VMxBoh5oaGtYqBNQvLZ2wozoRKj4a8
nDewSIVGLIdA/0Tzq+J77B8d6w+IYVKnFdKI4FcK/atukZaTwhVTifTb3AwmpboP
yX4KEcyhWjRn5wBf3LKJu95vqgYzxZwoC4txHASxLFb+3yhyQ0Cgxasf0Cn3e6yy
c3AerYzlAVhjeRfzvhJZpi52mv+7ch2MWWh3rOl787b9lmPhH6cGBwBGhkO0CeMT
7KL1EhlkZhL+hnB5u43rZfa6GPx9/ih0VKBM5NMxIB6+nHlxmnBFg7aRiX394W+s
geAiDA1mFSvXoZ4+ML9AC2+Uv/bkyUMzdIp1pisvucGm0eRM6rYcBS8Lb2oy0tJx
KztG+I3MAjHpTfxsF4Q22js67FpwJYAK4SMF9NWWefmEaSiLLtkazNHWSng6OahK
zvQXpbeagOMpHlRmS1k/LIzUGibOZszJcSnK5pf8soBtBGR8DDu2IvigRn1lFug6
pZAXVx50Xua6UWUeKQ/XfAZMxhuXzqyGyS6pttb1dZpJrtvXh3llgNO6lxIYlydl
KDEkgkuZX++EMOPIyARkOWKOIzisyZ9KpnaP7sKcLINMiLMmGYS0tjL1dhgPK4zn
Ftz12JcWjBy4g6A0OusfMHe2Q3sk58hQSARfPtqIbgYUGmSjqfvwrjuTJ2kLZRPT
Q6ddKJv7owwTvtfmTPuH6xcOMD50V3nCuhLfi0K07cBECuMBCgp9izmrVNZ4IGw4
J0nlZ5MWMKbnKZkFHunRodzRlqUz/64PwS23VxBx17hZVQujUOVujIfhetUXTaA2
ZyEfoiofI/lbECYR9NzhAFFwS6VjvkeO4zYckPyMPaHqeR1EXIq1NmdgYjRgDqBh
OX7sAzYXk3xEQyYQ3HAf/o/ightqMFzmnWDD9vt5hpJ9AUsYZXG+fUsAc6xLq7yD
CJ2xbxFsFcSvsrQUZWaFPItBs0AeRm6LhbmG2GOszIAEIxmyM6XZRYUxqPP5Bw90
yOe8CSHSIp2gRkfnScCP9hlBD9FgEo7Dwef9w+elxmAtrwiZRUTmkkUh9NT6mdFe
1ZNx7TLvrRcu9H821bTXM0FlxN2D54U/BM2hu+mko4AmOr1f6tcZk+zUOFsuQ9SK
KEUU1mDzufcQ3Iu1XlXKN+oLajhHPrjG+CnHmRXTwRttR6uW8OeW7RB/jAF39USV
hHK9owmr5sW+HmMgsMhUabBhug0YTT34pxLo5MtdE+wci2VTRCs7nmml5rxK8BdC
29v39SMM7krj3m3LAcA5C1jaq1iCnHAJaXLU5nKT/eRicGIWV0nlyzvt5JfC5kVz
RT9ENtH0mhxfrFqNZKTYVBxM07z3YfS8SwFem09sbVVs2YbFWzJKMAh5DL7ujSbM
DISJHkk9ya83cqRCNg5qiGdtIw3EMYjQQDqXy/IsLpxfEQmBkjgkbaacsOaOf/o6
+8L6L70JIVOmUmuaVg/8mnlvAlblzFXxhRtDzA2VMNsA1OHVFbjHE91Ds+YvFZ9u
7mCqrbrGNLZgOPfT5fAO/VlXuKr9Aw+Xtat1DXZjrnO3b/UKzGkEbsJsxLkpwRGy
AAgOWpEmsYIiFnCBWRyuNQfCS619C9oAR3c0KtUEEVip4Hclj5YP5/3UlcAqLHqK
RGsERJUpgodQjj7uk7PaHqCl0yKgbseo1EYwEV0q4fyzG7KyBvvSzQ20IZ8xxMbO
Q1ybm01LTr8XJvj1/UVwzFbRBfqrWItxkklB+fUzDsrHGvbWCP15yMDQYHtt88pU
vRSmPm2pOd1GUZQgbnHXmdQ6eIYgL1NNxmAH6F0yM0Jbxtxc5wLQJ/syxce9E8Hy
cRAgmPoCAeGqU+rEjFCIP+pFUukrurGR+WhkRInIDiE6dxJyyh2PU078f1lvXkUN
fYV5neNZ2Xz9vVQqAi87KDuC6fb91+S0BXX5e8QgRS4k4tLteOaIOmleqLH2Olmg
N0TT4eZ6ZM9fHKKmvoJxvgAYyRqAQJ1627z8Id1pLHfIoAO3/lbfkORvj/PgqUv9
wm424muidhD62Vbkjmy+msTmmTDqR6Wh4jtlN4ZLTrXH4/+391Av+5ZJr//Iig8d
2xHa9EuhcqxpHfXznLPX1cMe81avn6W81DjxU4KEvB2TomJV9BQyrX2kXyQLHVxT
oxsXrmX0Rp03nEJDE4dSbKVKQpKx8BqfgwrgQhnQspvDMv2elnMrATppThvruTms
w6708+MNAzRNQFPSlE/t225L+db4fl3Q7LgwOYS0mTRHR2DReczqKuhAR8CiT1kF
FOOSA/zAwzb1WX5EPFXkYJvX0im+XpKO16qvYlgMKOdgC+KNgDq+nlxO+NoAn8pB
yH3hpzPiXoxy7T/tIaW9CsoB47k1/ctycB/7zn4Ht9CJuMguM0wI3Rz/tAxwCJL5
DnZgQqasHgljznCcwhL79nqP/LX6GcA4Xgt3AhV0PhL7V3GojYWLq0+2rCBrOtcu
I1agXdqSmXg3jRpKtdVC0p76g8bhh61ZNWi1fnYpCbEca9PONposdXxrdD0SiJwe
JCrNoMdLaVlXWz7QLo2oGn5DQ/KCrn1Y4WtFf8KXusRpKGt+jvn6o3ZPiyzTBbwU
oIy5S3zCY8nVvDaDHtTpPxUuIV/hVA7MlymstWi9EMeKXBbtpNS8+Bo/ZUz0r9Os
J5gnEHAH2gW9AgUchMWJpuoyeQBW7oEu9xPA0DY5LQzT2BbuLhoCOpNd20x2vFL5
AttpIlN+NbTHABTpQuoipP/7vgYP0BsbjGPvbCWCSnq1pEhrxtI9zu5ed0OgUSSn
UWxONdYMeh0Z9mmNBfUvp2iXzPYGrE0JFlDQLpA7tw/QPtbXvQtNrH2mWWEBC2V9
WNmcGp8LsFhQWBuSo77gygG6/vEY1+Lr2jiD8DhnNHtcCuUc2muPDBT9G3WvMBpz
U7oIrZISNoG36IrlnZxLXBv5ZcQE4OoEGjDE1WCJhvXAvix1H4tIFCdorWY4eTaG
ynrTxdFJ94mDqcWrZp2OAH+RXcmoJdEcBPs95wUgS+Al/qY1hvFp+b3DenMZLJen
y7qHcxP3T1bKlw626IiSa4WzGG2CmiqOiCC5wMNGzAaNpLsAd/zTOruixSGHNefd
OYqbdAePmqaaGM9bmBkm0evicfsLurr9fQwILMwM/AMtPT+HBSF3Yf6TRt61lCrk
FOEjtw2Oyt5EqQ/V7jt8BGReUuq8oPHxXVXNTLqNx7yZwKiX4BRNbiNKE3IsN2Q9
p2QsnrH3wtY9pYDMehd2NYuWjNeBf9ZSVfriXxDqAoyrx8gc/rloBWtPXRkakIq2
2WLJiyhbw6Q5DoZcQo1nYhuiLcMFK4Ypf9HI1wdcaeDa6UgshNqfRIr1zhlnUG0u
NDqc6OiCwNf0TkiQi0moVy3VEu7mm770UnHFJzvQ8SQe6CWwdzfgFBg6ssnRqkED
Tsk2xcnFUWatGu7vS0J8wj5fWqEyINZY2025PPzbimBs2XPIUOm60ZkU54+RzCUq
ZA7p50rfILJS+FOSqriHkOq9qhd3s61gc8V4brrmsoJTZTyzEi/3CvjKBrqqIcKZ
tGFS8qyeECsZRekAFwn1sVG7XOwwNBIPugwdEsKW5LKSY+1HG7aB9esBLZW4C83T
04PTxJ63OKTyv2NcUrCt5kQHHEwN9qnpSg/+ZyPr5VAdZtxmXUyG5WebngubG5gP
n4v5YU0l3zy7LmzjglCVgP0JAnUbvB3RSljuqyQfe8+NTTZv8gegWM0ubPw7BbIK
sqVVEFSzTh21D7H9/+Ledeqts26mdvJfrLIqWi0cHG9H4AKH3El3gLgHq3Bd2t9I
1Pddw3ooyxfdIARLhmoJByBApCN74cxs+BS2db2oeUl7hCz0WJzA/UvZpcmeAAiW
g5UD48KGXcHL8ty1AaFbSzq6DUWx1eTBJQ0boocfeao+H0Net3u1Ys6Pt/l7RqWq
ZOq5bGQAHjzLPPtpOVoeMUebgJUifhnQNxu+t+NkCmLgiredN/J60YdWhEnQbqU1
iIPZZDxRD/aSC2Lg5qci7DDsFVt5TXtN4yp9WVURprJdPyHTi/Te3DVWNw2D3/jZ
m4xHrSH0uMogK5xgghryNNB0zLiAadcTnlJ1qHQGFVLTFnXU67zwoGImFS2+dYcT
Ze93keP2MMPXapQsdj4Wo7yJi8t5TKagz6xISGDgLvI9mqQVL+5s1Dl4hF/Ok19N
zSsnE08RlgnS7SLmaYOXYGJ+ctM2IlY7WB3HdcavJYLMtvpKYwKCKLJpCzoi+4pQ
anRLjHPC39Yy9SVOOQibS2BPU1JN8fcmZkOiQUTaQxKi5Z13vBYHK+WZ98fX3EWA
hYOGgmbNgn7iBnaQR1lUbgoCupNJJuVe+T7sFnYBMlhrET4faZzympbRviMubmiM
xkni4D3ldTchGDmrBcJlManQXAUMiZaCGcw6aoo1K03szDBjbGMvOlxfOgKUgUFu
vabFjgFE4LS8UickKc/eNk317kiR3f+hpKdMCzaM3wy30++mptt3kJQHXvMPoEZ1
ufYYke2XNu9ojJjOPyso/VAVNSuvZmxL6axEODYKlolcv7DwCZ/uTpMdbkb9mT3i
RFs8hxf0rgB8FW7NgIqV5Fsp1bmoT9sPs4HiU3dOjLcbWL0KRvBavwtudqTyVmY5
cO0yqPqmRV0yFGlC42t7h2kFlXa6hJ9VJiszYqITFVu681sGaCuzohPKDdN7J69h
InTgC6jP0kRVR78rLs/34l2gVTWCbr0orTC8p1CKbhvbuDvm+JbVGadvPa9bb+Vj
7XRMUhrlRGbE8KkouP6ksr1jT4ed0jixQfAmy+Y9CxKRLW2jtelEMB/zNIdmriyw
x1ogavoiQRWWKph6vskR1/0NFOXBbXgICg1pYChZJFZziGRE3csWOPuwd1XgYS88
ba85IiSLQfnpYpxRfAlosMqMU7gq3PvJeV5IgltiqiwMDHDwOajHA3lrmcvk8hVB
NuSR0ry0/twUWa2w7D3X9dJgQFdwyQJ9ZmcIglo4bWpw3cv7zwkVppMLILYbF7oL
Z/Kuqhabas5+G5N/aTHqtQ2SPP/7yJOi85ijxuvrVKDk4nDV/soYo07K5JXDlKve
Pd/E/4hpo+LQfjInacAUUfYUQ3yMJMxhtAqQRNzkUd9C+qN1GaUV2ZzNSTmYEqZI
U+RUjpwgQZGW104L7T9Vy7T3l9FCs9BUsBOwzO9cGOvnbSP4E32YBVpkoGU10kFK
SqSktrOqI4tjKjerF/OIoI4JSNfKfNK5SsYWCE4QHR/GJbL9uAFR9fkPBhwrvlet
16QFkQV7CDU7V6MRY6xXkXrlvP03b5ZimpKIjodU7w8yaWi4u3k7SSQygO8GrGua
fVUHjM4zzsMM8ZkGYkZQhSnCuEqv6ZZLGFu34PcO1XxqFSodpAGKZ75KqgTqtqHO
W2SjAvo7pDU303wG8pX6KopUt/jjPEHrYKxGS96RtyBYW2DY/mwic/RrCWXuy4fH
JJjeid2m+cKOj1M3pIBZpdlskBFwMti5V5yVjKDaT04uzQ03j2F84GgteVmtrYWI
zGvaUgrbp+5RO0c3uYBsqiZMdS1cWg5X8OQYvcfT6FNqLB4UfkqdW/jX2JDVAwSt
13KrsA2QfHuy44A/np72g+6JdZqkZeKQYop8UCDbHEgrKde7QJcXWJhQZp+4pfH4
fqs1bqyPceHHwJcU2iFrwABEogt1lwt4h28CloK+HybhhvZg8rEtwkrNtm8TdGPC
XVciDUMimvVqesxoai8raY+a5QPV6F+umpJyab4UJYgFH3kHHhxaWvaqO8duHFn7
aJlQZWgdmuMx4P7j1QAykpqXCoHU9Dkisq8Qk27H+h02fd+GMbVxLr/i86arcWO/
TZG5OV3wzXtV056OAiSvfEvFhDHxph6P8Oo3J7EI1MBwhulLbGckzMDAkGJCL9KZ
A16AQh4sG7OwNfr5l0R7uYkTRL8WtLZuYV9SCeKzZLqg3o5qkd1E3zl1GQVBvahA
cY08r9e0r1ZfmU3BqKGhg1HZmojsiCgbVQtOyZB7cf0MSkxB1NhXHDJ3CFmfxrhi
iodkTXKUR1w9QYAtp92oPiEPx/NBuifIr8opz9M2n0lGJQWRrJ9xK/lcZ0uhoQah
G7qA8PUJOSbrqXpoYgO2rlazwjxnVE4+HoRJ1B7xjd5hgf3FjxzdJ1jgZJFbW549
NE1Z/ibfFtHQBGKI12CGq4Bm8odSAT+Ox2dXHFCm6zwXbY1LtrT2S5zR2i0bdoj4
M6LUJh3mb9oRy5Bv1xwkqzqJMT8/DJ6RvRxPRCIBHrPaK/xUNzH9yETxobYGKgJy
MZvkBTZehb4hL0xQWA99fkfXfFWKEWOhpTE2WyJ/aADQF2fk2Ojxv9dkVDR3rVYh
R9/zhr6Zvs5a3/LV6Gse82o30eGu2TDm43sJW/4iFKZGXuYOTihkfB9Eofw5x2CJ
SX8bmQSx4dK8TShOjTSwdtjfx+xDFFd50ytPTHWhX91T0wMM/YYnRbNce/luq00D
xbAdpuAy5TbMpTb8IGENLzFPvEOiMttEHpGIxmoHWhwb9kiW5BiKTFf+6cQ0DW1c
RQGIsbVwyr12y6IadcRHu9uExdJs2TrcljUOJ0atq9vySF9nbD5lIEnRWQwKnBm+
wDWSTQCkv6UOSn9wuSU7Q67R5mR1WyVSWBgoBSe9Q4In3AV4NYpIEC9BkENcXVde
hS/djHg46izPvkWeH9d21ufvgChH2ibJHpwYZuukY859GZiIJQOrnBzlQ5JL1hR6
ocTwiN7rO3G2MW2mg7jGBQqKuQAVhr5E99xAQLnBsSJ15LZW9s3kI+6retDq7pCg
CKaNSSR3VCpoG9KRbZvrXQSdkML/aB/y7BdsTKT1vmrx7rEiVk2Thjdr5E7fq91V
u3DoBNGS/vnNchB+0gWJg29c5xkJ7lCIGyFMrFPw7hyIsCcU1ixLSh3LEHDgQ2Op
iDBJ14EE9c4g6snUqSJJ9z5WjXLCuynhWRsdUyLOutC3myN45IYcpUWHuN/ZhWvM
ILY3dlJagmCfKbK68MKR7SkSxsdnCp4BJNJALtR3MbpjblLioW61E9gpJQUs3uzF
12QTxxrfd+ibRnBX5WTFj7AEqricXuYZdax3Qqyl9kHQAHCRnTWXlSRR7M9rFv9Q
2OTvdf+ApxGV5xCK7Sicc0+IS9AcaJ3jmxp+t+wN4bhF4aUo2MG7mE9Vi1phQwLj
zgugrG33FrnXaFraUFlyNRdOSs7eT36jhZi8vzfP/g6E5eB5Pys8UAe825GvlIVn
L/zCu6zMkbG9A167pdR8hRv4Hh+mywZ8/VOJEdnSh09Np3QmmBny2oad07WlMK28
vgA3VGNPSKS717kjZguxAn9KR6x9RRsQrmj1vQ6FpomZLHmPLKUYox6d06Ke1kOL
hSypjD/UNxEJ2s84RV3N2yXjqnBAM0uwgKPYtw8a4LJdNYP0F77C8Il5OY6JmWs0
Fd5ir2dFij1Aj/wYxjq8Y9CPOmTGn3PUEbHiKSYZEDPewiza+xKqVF3DetKQfniJ
ZZXY2kC4tWwqCdYCN7FekhYsjtoDHLqzAyOfhpHlk/hhJ49IgAugS2XSJFfn4vI0
sKqDzuNOgL1jzoRiyJOMvG70E7waccAx9Ked05CxOSr+KMpePDmrSB9Sw/x07BSa
g1C65zctn8b6LzOKv5JABpcGa3f1LUzzS8+B6bWvap0UyUlWu/MCpXBMNVm68sL2
5IdiRzoGH4qkCxXOnDmBGGJlLxfCdr3EKfOiHgegpBgjkKfNvReup3uva64FO10U
HjbVfeaY/ngY9526noHSGx4T1YB6wXyWLuJpylnYDolou/tWvz2ZfFWBGcB8oV4f
7SIvbwvJbcTG38XiGS3MZ01ofvJ7T2eheE2Itl3zyQzGN37oRNy4i5hx0EMp8f8N
wN6TwZj1blScHKnkgC2+k5764wTOffYM6YkOPvok69XkPXGtC5eG1pySc/qyn+Dh
vb+WxU7imoApOLbNAF6+K2fb6IwLNbhrms2HiOwLf96fEf2rpKrZ6ghURPnCRPZL
anWwU3ra+n9VAaMRemVtW95YyLE9JGoKDuil+oHhgSxsvaMJjxPNCLW49aJFsm8f
uGVfOUPLGNs5XxXOEYyKNQa0fqts/+mUJpM4AyAQHjEm57gBG2MgA3qw/Ohk0kOp
KS38mJqI8xqM49O5q6it1O9GF9ZROZT05PIgRR+fy0Grw4OJAneICd7rPhd/Spiu
6N5ADjdV6+xiBCZ33UNuR3qHN6HZsEVHIlksNi3oPX+IbM+qDmxjY++Oanlk8mQV
nJdo1dnGgPozC5GYfEoJceDZwmK+z8bPDj/fyO9GoyrxDv6tNJKXfgjoj00pQQE+
gCIcuMPp5rLdX4HhwMvkfSiv50jo1kfhbR+A0QDhRB3Pi+hMB/KANEGNLGDoggUn
S8rg27/Bzv6r1Yqj3enIGK02ZXACvHDyeHsYjErbxKIthLfNPs24ZIafqcgPyqf3
Nh7xc/rI8XEePSEO+Z8o0+xoZuf+8HngEeTuC35MxupWLweysEg6XgK9XZY4EZeh
K3/RcSnOPakZPgEjhRgnE74kJ/rvZh/Xe1QuMYrwxuTIU/hdxaYPRxGsSPdh5n3Y
6ggEs5cn4DvOsea/9VBOrouuZj1zus1F7vqW5FZFUDQMCUoSTUiZ0Ybby/f4W9+1
GjAMdQMp4Tozh8qp7yvUlcvlSF27KmOsDcIu7dHPoryb7sT8VB2HRguLd2UNOi/i
AjTx94klsPRgGqA9uFrJtUDSjVgL/WDCU/MvsSlmOTqHGeeaWiyinDoil9HGEAS9
VlNVcytcdi+gVedNm8EkuUI7trF5b+cO6+VsCDeT/koFvGGsMpVsQv8pURnSnIip
eMCggSGdaRGm6np0Ump75uuvD8ur+me6HuzhsRxnS+Wy/Qk3wj9DMXP7ZvUPufzR
m6+zx7DvqI7HYnGGfjFe5P/BoJdODvRahs0VV4/tCTVtkgeF1ejAfn/H8llnvZ9V
PX5tOd/T7JcKgl333hJRNbKTzwyLTsUi1Wh8Xf91LNFCQI6Xj0YV/vgSvqiLZTkK
ZUC2K2ZoAieWFmHkKoWwfdRcuzd6YZ+MALyjli9XSW3VFXvXL0XieMvfji2CA62V
L6MtRc57xtRyappuLmVixCoesJVidQuCC4oFsXSVg3b33+jxiqmsss1ozXm9YR4U
e9ers2i9pxCnRrwSfDSHJeTXy/l9UBxOaJ+hLJYKhaXa5KO4tbr2hkRocr5vxCwe
dvYVg52xDSI9TNvhKYZOI/+IclXajZ/sqp0icoe+3y60ham988mdWjBRNO27QikO
YmV8ACiNZU3HY89Oewyhdaf1xJoIWvVsvwiWlOBpZ6FXOImXLhmPyDdEjQgVQo9p
iYoMExjnS8d3+NmNIm/+sLxl4ksDjUaowKYOvjs5J0Q+Rbu+4kJIKXwIoYWgsIMh
vDSn7mnHoXcVPSPgP5J74FQJhP1E434QW+MSKKg56nNdNLVrDcnEegPdjcCX+EqC
Vxfq87AZbixpF6roYniAqM6h3arqDWK7ZKihUwhFXOfCmbXejIog9P0b9D3ojpID
rlfcLyJ+vG2BLNAG/4wAAlgWUYXHlscRdiXmOXc/x6bozuekyw30++rMU89WlRtE
v6Xg7dhIHKSeNpmjgMYK1nlFyR9rogQqf+V9lxHDtBlMCo1GGDJcxdydOk0n9v0j
R69xCtfE6ftxukc1zHaCBLZO9Z2+O1u/hfjFWVKUmym/P06ASfYu+ezaQlInffSB
aynGIQY/v9bdMooDLWL2DUNnL6TOhHtT0yLhC9xkQaRRfEJLtOaDQ2c0e//RwyMB
c/GhZkXrz5Ov4Qo0PUXzvSUtcgj0ipjvMTnkVekW7HriW/yOY6b3sQIdltJIXyoF
mDxWjthPQGQzipkPPNBquaX8rZiYa0bO85wcnhlbikRlEOE2tsyVy7Gh9HkbIVrI
mJJhiUm1jDyL742OPoJd2btgsK+ozO5YqUBOjVaWkbeAKxgzNGPXI1AFOcPxYsx0
72Z3vIrezBHnGeRb5ODElfRyRpPWGdzbIy+zSoj8C5DQ4H+pp0S7LSphLosBCsIB
drN9Tb6YsGZYZFPnGRj0++2l4tnkZGsuy4R302Ofa6PT6FO4e98v66ya32/QU5E0
X60WWcpzSPwZrJiDANMC7JAGQVBfK4r8nxUfRY1/NBGh9o0n1G/NGpnymVk6SrUX
krCKRKHBupd7RQ5pbilWS2pCX3rIQ/le4Bt1vKyUo7GvpeNlXsZiYUJFJszEY3Q+
XuhQLIGm1zQI6CzpixRDJXIlH4gp4CsA2kbtmwULKZkAE3+JLeLiW+c/fOpAVYMD
B9yLIUigE0uDye9XmuihbRgO1YSUTrRqbALf05llLytKrAjmKOD2bd6eZZvIIk89
Ub35zgt0IWfcXcLau5qQ6eJnjaJ3nxQT/nUcmZXy+90du4gFImNy60wV4wAU2I0w
7PkHZjspPzxD4u7bnNpitQv6YEzfOKyV1LxUgO9Z5Cj1YC6f1eHO9PtT24wPOis9
iqxu/U6sjLwpwohQ1dpBnlGNKXWTQeZnsiFptEFIM/ZIKZT528fSMRbaWgZiZmr6
9eDdGvrs83LKrLRmFLmv6giw2L6LwXfkZqdvxb6rQy1nVnsMxg1GayePo7YPRDAH
IUzfEUw12CnOhf1/blYV8VX1OAfNzYwWLhBZHw4c2/O5zDKIYUOBmAn2ZcoxAm0Y
+6SXzStpDjlfUl7VbeMJQJCjN3PGmZhtgkzdMAqJrPFb/aSHnfH36+6LgrrSesk8
RUIMMGW431cRJU47xNlic3gOgE4pI5UKcRltb80BOlQUz9bBIQ1RsYypAbYy118m
nXhFjGENT4iUyagSikOlADaOAjewXuvDk1paSfsC7xX5U+5Q5F3ogg9LAXRPu+oq
ncC4fxrWEqhlTzAN2bDk6xLfu7Gb7TU7XFUlpqo4RHRN0iTlLHz/62G5aGsm79AH
Z0tziHRekDmGoMTmE4z4sYqKFutrLnjglUxJqiNsqm15siqbj9iBtM2zhqFtAV2O
xs7eUvbTmFMxoarqdwxJT/kN9sCgV88Nowkd+FGnWvGsf3IdN+XSerIyVJIxKQ6C
ablCFW4fT116n1d7jgMtLivwcQjT+h3i+XiBi+tBLA90c6E1OHu89vIAHg/6ikFq
OycVeAT5nukx9tcM5JYLAzsfu6Nv2cXsvvFiJZ49eQL5KizL9hB2RWbPT3Tz+s2W
HnJJBSBDfZUcyqPt1OU7BmyGLJn8qfCZ1YwTMpIDEs9vTt7vo4pvM9yJ86FtEugx
ZrtenFmGJjxrjTyMRmmxFQgD/3Rov4c8FuvSTXx8KS7Y0eNTi2OIoanEMpUFCK/+
TtCTtDO5cXrV2Bm5ktMM89AqgnwjeNbgALR/vU+bAPSeMqNGd10tJ+vg+oqQQyPY
USABGCxq5wbnWF1FO8rbsywEH9OKWpM8aUXPPAIZ19vHOXO/dI2Vbu1/npfP27HE
c9imqJ/UyQBpo/SjdAavJCzD23on7rbkKLDIs241SJ6EPKb4iIGVozY23qIjZA8k
59nESH19wPpMZjVrMnv2XPDfSYcQybwYCkkzfoXJyGn+Gvpy1Tr+7/C8TOmZn6Bu
vjr1v2J49z36CpSeXLwLOKWoA96D6mGxqvsYbDtYTR6xnuMhd91XpbtvrumSo0mw
WpK06xcEojpoBTTL3QL21rPHmfUNQSNbGP6cVf2Ihh/KE70XTFNlKjmW0DYGiYlC
8uMgbwPz7DeKZjOB/rY8NVEztY5u0Wpl6qWPVWEkju03Gk9wAbMmy1haWbV/mEdO
Ogh/vf1KLyHnxK4YFKRgVPLAMKBZwSRIL6NhOZLCg44p+NFCYH+ahoUuq7wy+4ch
L6zNUoehPd4DPplJZaetOizHQXjDIgPMFsjdQq6+M6vyYy+min6uXknqgEF/jrvs
q9HSzKK+M1KcxBT2t8tP3ljZyQnmXefCbpGAtMZwb8uyELm2GjMn/fLRqGFY+OxD
otZFG9O0HxAdQB0JY+zo4nq7apgJnkINtAZLsMY/xcvVAQTHE1JH9AVrYifFF10d
LL4QUw1O2WxJHoMBt1/93zg9ZbMYT+wyknmoaX33EUDdaMDJfg9tJoafBigBVyDz
B5DnMKOfVAG9Lz+3zLw2yw0W3o1hTwj6NuYgGzlvEajCLRHbrhoYNGP54Ld35EOA
aOWjL6tcIY/TmvtBeHH8bwoGsr0AJdFaHWy1+DjcTSpxdcCIb3nXQmNn1YcxSfSJ
h/o0mDAe30W9kVsXYAK27XFQXG/7ESo72ZvDlKUeXw3VHsVCvhvplWHf0/o52e3k
rZSELhjc+A+jsv5Eckr5Po0oYAz4UVq2R0E74V5T3B18rVAsdL4n08Yofd4lNUpL
Dd1MFY5kDGjf41TMx2lsUBFSte2n1/qsWiDtolQNTaslmmrmtGj2zVHQAD+UErrI
+28Pi2O67gAjE4iVnQWCHATeS5u83Iklaz/goKwnknHD7fOKRWsHM+LoJytRscQD
UsGSxyZ3hFcUXjDh904V8acSI2UWOi6t6PnHih9xBaCtvzLfKV6iiTYeXr/bf+Ll
sVGLB+oepd/Su7yfSoxxV2y4s9cIS6fXK2Wm/gyzt0v/RAQh3rUIgkAsWeMbzQsz
xttPE0NQOgUM8PmRz7Q93z49w6BH7lGg9yChj74noLLf6Jbh/rasWOPTC6VeYbIj
PiRFN5d/FocNyLbffX7zwNb0yYGiGzOt7HkwKNzMFdp4++uklNrLyIdl8vP4nDfW
My1On+fFz5P9kNB8LVGlcNjDj2GJYFNegeKfHxsw2auf9aqDgRHg9owYXo895FCv
qy62f50ts2+cZBdGXDkbTi33kDVvjhCDCumfNM3zf/1h0tTb9duyicK9BxfjJ1kW
8QYh6ioXhQV0gOFvD8/Y0E2CdKJgsZa17xr2dHx0z4aABdx9BdAJ1yRZVBtAkwWC
HQ6QRQb/Wq/cZTRrnHSJDAiELDBfrQoNukSq2ocw6SXdb7w3FCJdIlT42YBnScLh
OvsdUFXsDgSBBB8tN+uCOjTxbeipB0PYEzwSVxMcrTDDsxAon1HoWvtqLZr7sSzH
lHQ6i9CKZzjFs+Sc6h4Nxp1XOF3D0umjw8BMmF6EdVL9xKI55B0SCMX7yGJjaiFx
Spon3ncyq+JRIBk4cPP5V++FFlfGtpcaRdxgek1AD7puaWDidsshTiS/JVHKHovc
EbIgdL9S9MWXHe4RKk/RH2GsCu4soXRE+357xUgCspcjhqlxxsSjc5mJQt4hxoXC
lvj2E/Te7/ZPQ3ob9/U//b4fmUpGxvRijUvrNM7nBDFGfuGbDIU0uQFtAs7iL2Wv
U5+muKiH6nnbDMX3K7xW4lXRElSbOOik1twk4uTF7rBs6bpMBbH6H6lDaLV1saon
AEu8WFv+eZKBiK3277AW2BU+NJo11jPCiL/wr5K5LH4zKQjZJYmWPEYOnfvDHqtO
m/m9kIqxJTD7RXTpgvdW0s0vuInYlgQ71z81iCcBpnnWrXtF5aF1enGQEqOCWKcM
KB4+k+dkIFinYUCxWIlhLsieSYU1ZyjGFn1PIXBQF0g97LxuPdMrehE9FEjZ6pQR
Le/OkkMB2LX7mKlJb8AxOKZ6grm675q1o/6avPAexP/kTgjc4rI3icsbQtiZ9uAI
Mp/54sq+5ToiCv1zTEe0DBthTlbr9sfGqg6s+SM0Xl8msDnug2KUnciVtQ9gqW0P
hrjwtUsIVo3lX9ETxS82jNabCIVPo3OovR8UsdxzIFE0TG/h0ZwSA5hW25GxFv1N
Yn6OkUuXqbzQfEa4NSIbqUmkwrk1wh2AjiybAkqGluVexNSvSR1bGgzd+1xokIWL
aKVw4Rnpc5yVpHyXcWFQLBHhksKXfl16k1DcD7WCRoiux6zQ8kyECzplfSETMBv9
TJa6cQjXFX0OGsW2DRRouf8YJ8dEbFKpuTBrk5Jlwibqz0KuszEIXZfkcVFfOe2w
sTUHcu39fC+Kcy8QWzaJgK57A2yEW38y4e+bOIjfIUD6+SGqD1wk4nRP8OZTuf54
coHsUErhAFvzGaHR63DcMm4OM8WZp9f7wpmz+bPdxWiIT3uTFrjyzrwE3zQ+G9BB
SXHbqOHJbIZx/JdbCmcjqY+0QqGrXUWH5mw6OYh6RqmIXFsCYTrgPFMpgfRLOuJH
jB41S9fyojE6sngVT8cOhPy9AZOFVm+VshXegPp20RUvoAuWPcoHXYcRHtBDDpei
PNaQ5wuu5d995VR5dlpdi2g6PRys/uGEbCzmya6nDJw4iYCm/ZseRZY1g/gMFzyN
fOtgPZKhQHwKXiFV0rzhV8vBDpNu80jHzMhXjQUN9VbbufkC2rND4/iNr04SCq0o
CqTFIER64kdSEbnBkpKyEDYO8gRujCO4zpOfcHJIxUmJKK79C2cfXrQHqbRMym+l
LCluB7Yie0gvm+WWOajjMwCAxXWtqpcAQjdZcG0XV7W3G5NUKMLrP8rnFuhFpTjd
fVErU1QzuynKeiaWanPWAiDQtfpzUKP3OeEh/MA+OHY4AvSAwX5jvW159btDGFXA
FpS/CXEE0GKBbIA0Y59B5T3LFMx/V5AhwUtUvQU7lXhKymwmPtAEAU7qYTfFCqKO
ynsMf7hvSiAoaXSuUPMqAb6jmV7+ZTcqIxrleziFh43waFrpLkdi/mR6mjRV+8ez
tEQX/F4ic5XMGHT4qd6BpeQsG7ocpntWTTReF/hnopeXkvijpcbM6YLFAI8vbX4T
IUWzhLAq+RSDISakdNQoCgcmC/8mbG/S1UWby4yAJsvycNX8nyCsOlG2oEzUdPcz
iGYJsED6DrRaN0s7aM8WPtWJ3jxtbSwlhmVtFRH/7ShY9/u1F5aHpHspCjnSYBAo
MB2U2hwQ7ucaHpIm9mFB6q0Kf90Gw/UpwyrcuubwSt2G/ebi40ZxntXGLvF6+VNq
CqK4XhUbIvH74EzZo36lfT+bohB3sqmtrvELRjFk4nOtbzj+sdwC2k3oB/ay6ds7
QBuzOvMOCik1xgBhS0Baa8jcWvClPg08x2mZI8yasBHvfYwBegAoD82joabWOcRx
Cj9F5ZrEO/aTfb+cPK8VPyFWUd21MkIvyBQ2sfDKdCVavZcItGOLSx222zZfG48f
LjQ0jsSLUrgFk/b5rqRFXfqFwe8M7vVWzZPT3WdulK4PUcFWsUC8GHqWmSdLm0xC
jLXvnBvO+OQusF9zUhRV7kY5v/uHwsOEv9LBIa76Sxf9zaEqGAx7CXiNkgoGA0ar
U5ITSvFOp7kwwGBnqBLdDX85sBAyHzKNBsvCJWLaGXHx8pB0mb5dCJEYf6A97elx
J6oKD8MCkXDnkW546zB/o75d0RTIUzjrEKO7iUMOFrE8FqM7NaZZfy3B2SHzv+yb
HBZ/WJI8C8/593UMQWIbf5LvFW45E30IkQktWWiyflPw4rFrumOSboYH1Pg381Kk
srW52StU+PMoTcMIGKhB7SPyVhWCd2QOlFG0mKIC6ffpqnTmTXchwM2HFrkq3Vtk
fqg79A326vr5TDfCEmH57aweud6PeInq60Fi6J0XdirRPpz7iZyMqb20QX4RNRAj
4D1m7ACZbY/V/9K5V8g/lsSiXFFOCFGQ6mp2KbXe/E2Fse5uIoQN0UdR1wh/h436
/Ve/bbv+Gd0oBK91ZKiAgIuFbyYijDcn04jBpJwzgJM9UC+/gKCuDn/AKnrtFqP/
LS3EhFNU3mchL2lzwcBTOjMnFCOwz0HOAyGpk5ENduBzoZqo4CehsFWdQp1UrP1z
kmMJdjaEYSEHKb5SRa0K+PNPbX/PFJO6vYvJ4x88rlGhE7QYK5ZbaIkFQP6HWhZj
o2ZyTPUzMdkBiu4NuTGLxYcj/u0EGI/Ks9rRarXmWax3U0LMjfqu1HoZnAnSQ4M7
8WZMME44qyDEl47eAWM+rtk+D66PQ+34Z3vfdSwS837cLoYfqPhnAfSLhbLACWbx
dARuyJWgFVO419g5tP63orM6opb1OahUoKtQ3gepeutIf0bntq/wXF/LwXZlcjZw
VZkV2EW9FuMmTub8m2nhRPuOUPaUORL05OWT5ni+DRGQQuYAWoUuXXke8BqjQyIx
ctWLvpQCiVX9rALryx+p2kbzQ8S3S7XMm2sAgEVPjMqbIzlSxln7yALRjEgf4NJK
6fqzF+Sz1glNBK42w8/AnaBCf92V0Bni3WkYlhbeGz/BOYG5P4EF02iuAZMhNChn
oCuSKRzR+BVnTTXXr9mlJnGXxOkb4r7VrFZOjk30l1OcwuTuYYGuKFQeexGYCCQx
DnUyrTSzK0xn+TAAVTkAuepPIwgnBoizK0P1QeOuYMC9R+qlCyN79Dv8SVsRTynk
KIOQBaKu85+xrU727jZJrxMXzjqozFkYTGpPhz/5eNDKupya1li5vfngGMStAXQN
1f/RxF2QXaMOuW7mufy5b6kofUMJwcJQKS7hYFXYSV9OvVeerswQPbemCxu3Tfq2
ZzPI4hBZANfp3S0c16MWn45PtC/SNvMjxyMO19644ABTlL8D51XdXhwsyQrYAzMi
apjXUih47wETDR/xyMclmvGky5Xt5pDxnfVGIwUNQx4IaftebWBJgrhdFlrlsCq+
fuuGkbjdRWjElMzWryeBQ3nWjdmcfXslz5CWKRI4ri1Fz/F7wJaqgJZdsegtZ2z8
WCHJzcDovfw//fD6fvCK2JoSEO11IDcuK1qKZ5A0orgcfmmokn8DV6Qer4itBIdg
F/0x1qSi7hwTBs+0IddwBqTUpnPTZV5kyuH0/tQLluGw+6W2yzj1E4DsHI+uZ8SK
oDo8YQMn3KqlBpcMBEElNqUStZ0o9GJ2AbvW0iIYE6CdM4sS+q+l2cbhivbMYZ3Z
2fDZI60v9YQaRWs7yE+MFX01/I/wew8TXBaXq1ik5XMbrLZsAGfCg4mouVNy4uZo
c0t+4CsIpTIunQ/xOL6txOsOc6MeauPEhsqtcazBdYpQprv6ZlWRuDZPjUZtQjwp
LPBtbFXkN1eOzMj1xEVLhy1/EHLsxg79TUX2YZQjI0llqacDB0e8LBWJSrBkoP98
GEJINsZkhAHwU6xhHYulcY7TgxdLv/h+S3oBnnfd3I7aTLQcTvzFuPzp3vCkrVvM
eUkiK+JzYHUjJCbT5G0rrsuc2Iv5Pt/vNkFKo29DJHrupXy5djtK6h0QNAV/WvPz
5m4vLiNZg9PhsqwptwStoxVyxKFbm48y2iYkWp/RM5o933RXRJJS0dU3fVXAabCx
ubrqiH9eVtpFu8qO6s9CI6X6d+k68G9QpXKlYMJIVAnV9ihXLcIOJ2LX9/lyXAnx
3qV0WR3AJT6HnkUJedSb6ShZ7/X4uC7uWBN/eEA0WBzF3SLBnhsBN9z+eh+q3BzZ
cTkfjew2F9KcelOfSlfiAEJWiQn/lNlfoDlP3q7WLPaxsGkSrH2mCca+jrAPBoY8
tjnb07apQ1RSXCmr6T63QUK4zOhnDbOiqwbbwJ4Yhx77W+Wyimp8+fp1gzqM5CZ3
o/Bu2Wt9X/wQxLsdjAAjK8hhgLKSMJ9bSQh7j0JplfE2fLd42vT7M8SOiYYo2ZOr
q/rEihkiAIcfIpiFdvd/JSgBx+tGYdXz6mWS4oiSvC+basHIHI/jOitOCa3W6jW4
hfKoZdYGett7l0bTlsJQWUyvHsiBaWjqpHHPGfa2IsE0oxF2cRIsNlQqd3eCXEkY
s9vIeXXMk6cvxJ000W3KU0X/x3KAT8oQ4uSKp15bUHMQfAOvmR8IQOx6bl+Qw4Oz
mrjoRsZcjvUoRI0r/83vKARSQ7UbSk61LHozfuaHwsxVkSru7KZdbo6zhM6gNtK0
bvln8elbrkyTnT/oWpNEuOqkjJEoLpt1EmGkGSgOLFUXTbRi+mTRqT/PfevVZGBT
oP3MgaAmbgKbItdi0JQxpFAdigj14orzTKVLjKiciYR9Uf/FHeu4XvO9NjYCV7oU
wO6COWpvmBR3IhCTF2FpsSzFysvfD8li56YUA0GRdze3LO14QZJMkvVpbAW2NaDn
TGaegELYdAXBAxBoga86I8V/akYct6RXe6TuV4TF64oe4Cuak3X4nLpXo8lmFpkf
ZKdkBWujjwo/Oeh37zFd18Xmf/tUQCwqNHIRj5/rrtW6fukDzgMcy+A6DdWoeuiI
hGg+qnCke6f2LiHhM+V482DTT8wKxOgZj/jTRm/UNtXPB/71bjnrqjFuVpxO7OmB
GqK9rwAPF8tPkkrWuQUVwqKlDtnj63p9EPsPvfU9lCbhplKJeu4ICTds5rswG4Rm
bMGKO71roYfR6gLtiyr3uJJOw//OZt3Y0DY9f/GV/wDPsm0f+p4PDNAaCvuf2Yq4
tRaDsG/6e81AKfOhKs1VIPXMouaKRO0AYuesDd6sWCxhun2d8JbSFGvgabJl/XYH
coeummRl/80MAGho5hocbJIKivT8EdWYD+L1m/fIMb5sb5BvdK2JLZ4TEpGUNDyn
RdhwQ9eaPEB9YtE9QOO8xJ5ClBfOtB1X1p4snOI0evwozxrB8pQ7WUssly2fkem7
4+mD3ozvp6R/VMfe1u/ir8y0Op4cZOBnbxzjmdFyM8jwB4EMpjGjZsrJ6Psq6QcJ
6yXvwZ+3z0dN8yk9OIR8DD6c6842aO/Y7g2ud42g4AxwsMkppv2ouS6Co4tPlIFe
CvZpYyKZFjXDTtRiPefiJq3kv8/ACp+Hv7SVV9gvrCavm7lpkv5bo8Vi64gmeOgH
4EiNMS9iEod4AZ44BtyDwyLhvRaTi9OtWxApd3IT+m00p/BlR0kuiJ7IH0KtZIV7
B7FbPkah46tROPmgv3O2EjubvEyLLx+5NSiA3PkA8j71jiHlS20vRTUPdZsXbN+V
eGjyVQxqjguWutvVywygmo9eEn+oT3aW1LfbHDU5yM0LgWS8jEHoLfh/cO/l3Qdc
Uni7WUJoYE9aD5IUSiw0e3gZ7h1ty2CatuyKJ0RwiMBS+VcCpLPmmB2seDmrxHnd
u9uravoSUhRph2ELFZwmK3STMGlCQ2fRpcsxX90iYKvrtEvh5CXLBd8zVyB3VdUF
HF2df1dfC7C+zsDGlsujKLB5KoAbl92FAmINTRx8zKuX7s052r/Ac2YQOlA+Yi1J
S7Fewttqf3J32LFYSTRlCr+fX8/sN2DUyQ4WwB+Z3m7YZ2Zr9qrF739DacdI9V+C
tiZaGsTtco3ZQ4HlGwIwa9bhl/5C2xCB1xWyUOd91ioWPnKAbX4PRDlyEI/Fa+xT
4cDMjuuiT7YP68qN9nzozsYBaeVp3lpLu6iUUNPEIcu8lty0xHa8O8V5ReK1kQvj
n08v515s158XU5u3NZU0psDES04Lj+jDu4B1n2ns1rL+WmyjM/9Ekt++31Oot4X5
Y8qeYonlyAxEPFNS6+mST3Ug7mJ7o0spdzFRR4q3OMSFCA6JNgvthTpxIiwVg3mN
4BKtDyaiV0v2IDZwyZXAN2t4pS5X/sQWb37kCGUPtrmg5cQ4fNsxB+J8AgJST04n
eseYW+sPcKmxFV0h1Va45nO6vqfBUGjwcWtdnP1g/TTkVfEbOxEJyv5Y0rdaxGYB
OpOU064Pvc9W8Hppqn3JPZg6jiKaYOStHSqYreaRTcZuAcZ1VRMG+YrCfK/LrPgb
bvYxuFYRO1sBtnIAyxjwsTDdP4OJ1Sb/4Er2ecmsiixaa2MP6tCbcNbiKeW3BATy
fvR/JLzb5Y+nwq4agTR2pjFfNIIneQ3C4sNNF0uGtrCsnJ3P0fP6+iFuPe0rNYpa
PVkxtSTS/XKiTlKtD7L1fDTLCAsXyUqoFFlVZCawi+LGQLJfYvENWn4KSGexfpPT
dF8D74pmhpBd4BvmaH2JuFNJ3YgHVLqtGeR6LsUEQWpe6h7/uEcNpdqZBcgtu1UC
fC8rUDxm4He4cmjyaNfdDiLGI4iCJ+mZ7+xea8/SqNjnMZzEB6gxa1kTl6LnyQQ/
6T77pJw9gYY6urNCZIODzKvRdxHp9T/72onYadMP5RET1iNFed34G2EIhuugcYZb
2lJroxFE1f2bGiFEWTN9AHkj3RFH7LwbP/ktRzh6dly4BzyLgMXDaFtymlRZrisb
KTSI4eCmFIvxXBgHXw38sA1Vch4y0BA3NAVZt3VhogGzmWmtBKSqWYTYK5dcV46L
AAYDeJ7uWcCKPVlocF7r2UJIHDmkZLnSS+oOjspyPcTGevI9neiw9FpjYvl7ru3x
aKgnGLpNjhJEYQNcRdniI0xRsCYUpgsFTD29/ZxguqW/I0FbXJkX4gIGI/zPSsN9
TR6y60VMhPTziVXL/dcxu3lSAZjkUfQupewW3u61FPNNVwMO8p/GJWPb20f3iPRi
d2U3jtY8/kGprvAZh1NGaO5owq+EUJ8Kxgj++sTayOsaa6wn/xIKy4nqg3fcVh5V
tzv+iNrYvmH2xcm/cqEOu61mYReFj5nrpDUh6fBmA/RuHq+EcddCfejAi6iZp425
cbd8q9Kzd7+isvR9G6fRf+QYHOfXoMdI+dOUYktugXOAVKh1Th7Zkn+JgIpl7K/E
LQjza9pc0BO/77ZHwwbJw3+vruZsq2TVvOS//CPzVnqdoIxyfy9nAiWRj30YcunP
HxruKwnphrxxjygc46AvqbU4nJavzUNTPJ3P4We/uLSLSYT5Pmax3xyQ7PIep5+C
AjXtb2VsCAQiK1MNCcY//f1e0v4RdyaEGwqtjrTLBOJKa09eabjQet8YROHQEmqV
D8yf6bWLX186ft79zseAuSZA+JIOOMFzqWMeqvdXQTT3KgMJpJD3yUzKnK7PyvqB
TYLcPk2WkaNZeUu6VbcFfoAM4gY2MXpFwdvaoKqUlo1a9Naw7weN7tftvczzStrF
5ROR1z/gBgguarrYbuy854kYn4gJIvAW5U66jBCDjjCnirJwYV11aNFAwJT453CJ
OEZBK4PF+kYD3ICm1jydl7auL7wmhiG0dP2C5obeEFWqixPIFp9LmXt8k6QWs3Wl
WrBR2Dd9NNsfuTIAlEnhFfKOM9GBy/5fdilSECrLqv2lNJ57+DuEJ27pkvpMUXAB
HjhNy8iRrjV38xDJ8AarWpom6tdG+W5bcljK9oAZUD30DP2bKEXMivPTgCcZ2YAq
zFA/1nSCOtutUsSca6HtkQs+GiL8FZUEtz5AGnzOSHFjNTKo0AbdIMVO5D4v3nvm
iltBDjsDQJxOgO4nD+f2/Nebk3HJcARWFXxbS//VOupkI1RZ0kFUFMsQOKq0CLW3
Nzcxxob/T9nQcvtm8n424owr7l3zKBdlL5awYQ7bMY7QdgJX3BaxUihDo2Wa2AfC
DBpSNsqcCUFjD2bc3VOTZcXovZRJtnKhJ0DehsmXqS/ZguEv8NLvFsSxRp2qoFhO
2OVFqTNda5XvtnU1EDrAVQceRIzHUrreF6nztD8uaIsXyUqI6+fwAXV5VPH8uQ6U
I/lhMqA+qoIGRU3Yvc/7L9vJm4Ld5j3+TVovJXvolJhVJA+KtYpR4Ll2UZglxImU
P6C63z8SQAWXUsF2jrxlb1YxgzTu3RiHTF7ss6n4NtN6wvJT4UrS6wFoDY9AAwIs
ncLXI/vtV4oTWZJz41TOE0HHS1qgj1DzOpGizphasSy++vyHNAPRSt/HCVqGPBHg
Z7ZxBhI1H0ZxoB5rqGuQoKhEcBp2D7ZcAincK1iZRBgN/fsrKhoqOInutwgsBH/C
MoqR2s71J/QxkCRdj06YnE9zmMr3QIpXZ11nP30Rgw2X9TDOw+yxM2u8wm3u0CvK
0a50Y2FJ2bd1NXxl7pcWlu8C580pKh0oXEMLDsLB3QwEy68HUsiKgtMNCJ0MlQ6G
FvB4PWFoZWByhERSLFjxZKO0pBxRxvryVWosezxonoixD0fMFz3kBCkXl4QT32ji
9pwl9vuw7alwH3oGSFzfEvbU/JnV28sa6k7dFN3byO9snT67OMLiz7OTbTi9+G8a
ItjSkV0GqPSNhitbFgeZZ5DuDO6M44g4RvTV6PNdZQy+z5iBOBTNThrvGmAn0cvV
7F/fO0TCKql03mDciKkF7/Q1ch3+mO+ssJgD2KH9OLU82vwX2TPrOM8zyprlPxU9
aNKTFr0TJWwm3JmvrahbJFpqyenvGlBVw8Xl4dWAJqe6nQ8pYTZ0AZuAflInPsrG
IMUu8YGinU3fLKiqdqR+Yu8rUfVBuQuzdnSiH+LbAzBMER+Bec/QGVmce8n3p0Fp
7JgpBqMDlZBYUrdy094YBJHvCHvuYB7qShPBnCDFfH5QW8Xf410v/725vit/6TaW
Il+CSzOYRKguH864gPvewNwmUmIAalIlgszxDl8a2P6wYBB1mDPwN0w2oMmDVK2C
WrpvNb6ZGAPZzjagr3qaMw3+ViIR3qDYAIrDQ5ctzdoV8A/aHIREP+KCm0vpi541
ymbgz4SBoDl23vKUB3I3Jk+J4gIPGcyFr1oMKFiLdeHcFChLfVxygZ5hrBc58/zM
+EwRZWOGsOxw8ScMAMYAwvFLJqwN3cU9gvgMXlrAMpOgYmpsTfFoKR0Y/CKqsLl6
iN7vo9Cw+8Szg9IiJxKhpnCGyYmuSHv4meROaLHZoSZJLH5XmuhFH6mSo14/1HjH
3XHTZWqczGlRTWzEo8EW9sIhbz9jTuGudJkj+TpDNT/VrLaLTg3k5QDhiCno858+
lzZ06OKwZ+sVkFm8DYGF8tR/2v4J+xnCbog3GXpZ1RyOIMYeDSoZ3KfumpTAerr5
ouKZ48nJ3//g0IMK+48pa9MwaX10Sj+LKM1A0nOicolNg1ld+/bENEXH2xmqX/u+
EUvF1h1vR/N8X51lZlQ6eG7A+Jmuy6CkYx03n4sK1Jz385Au+2pLrNdCVj7nbRns
7IG12ac2CPlLTLg2tgRYztXyjrmVnvtVPnmgs6QtJJtk5CbAju/kI2Q1HQReyf1D
kSAuJNs2ZpQ0RlEI/5k6zS4LJ7PI+8emD3Xl1QUP+EecMYqcgvAWEF7ixt4iroag
gHGt9cHQrVFaCMolv3hFRqoCbLQoGipgBPI1TeN2M4XIeL0OZkItCsDAZJ6zHHwt
EnFLb0UGRskFknhy6aekXNohJfxji5j5a+Lu3SIr1MvKFlS46aQsDx49tnijmNXU
+smFNlWgIri6elfALPJxipERsj1S2AqzLL7WEZYLKQ7R9YRd1ERij+JVKgS7CTCc
G+mItFIfiQBsgHCvQy/aKepGEpbSRo4aSwzHqbGzIZjI59L32yVh9EXJefwvEE2o
b3yvP5ZKacTLb/JNbwHAAz2VuZHnJ4TfBByt9JsqGvDUVrmhl1z7CDVbkOWC75TJ
d4zxS+853kRIZ+GxTNvdTzW3HClF8j+7PYxehD/ibwJiCPuOCLzK54vNNkVTsmQs
SH5O5eQ497z5ezv8rNbsHcv/CpckJZVU+BmMMlNip6ce7TqLiDDLS41q4unCf3lF
UYNkXjmfBv4T3ZoghzBQGLCi1rrcm1skNFyeIJ+DaT23CcCm9L8Vh3iiPVBIlbwM
lBzG/SGtYhm1hdKGFGbgw+5NJKqNDF0BqJUIeWurermaVZeS2cKEjmR8M3Jgli8i
4DesjXvL4Hw0jSkehCyRjMcrblyww3wh/uEcVQ8AhQ9TIwfNR5g0wGkjFYhu4OeD
ZK78od3mM2+AXNmuQQ+Ft5O3jokpGSTEsPvIoLLZ1PfHTrhTaEU6E3KbKsZ/1QK+
Scz/Rk06IX1g6hW9MrmLEnVg78cFrbDt0VgT8NkQID96KkM7DVedBJP8Zi8g6YO/
Vev1C2aZZwRrmEgo6TOPtSmTEji0mW3Lve1DyDE/4utzw1aG8KKY4vIVqU67eMO8
+ae3hBCtPDWge0CXOmOUfHVbD3xliV8/TXu3cEnMGTmWuvS3zjn91IP0Jamc3VRn
5W37v8sUqc3nGHsmnSSDs9FU1y1QRjWQLVnDHmC0Z/IR7xmuI1wc2TRH4qtETVcY
AvPmg+2D5twDiSoUMc7ICukBIEVIkboGhxlCKj97LhOZfg8KvIHhWtE+OzQX0P7f
LDID8eHuGNOS6HrWpr/Vp4ACicpvDAqmODIY4vVevkePZIda2JBXWNcVVyqbKVq8
qH710SXl06T3EKnMtfgy4jYR44v/FJIyUakLxI1RW8929kfv9NvM5PETb6ijHO2W
j/8cxmLOdfyRiKmqFh4MSERkVYXzEAehjrmHwHJWIyU/YRus0E6HG3JB5AboZOSf
jNpzZfgoaxCW6WG2lkbyjkDyFEZl9+HyqdknYdJ09JDtcUkVN4/j9ovEaSy/Aaa7
pfnhjhCcw9dzwZgY4BQQswxGVWu+YlhjYGe7j43Q0MWsrTGymCK9w4S79Vt+TCXr
MPg5J4J9s0wsZ0TScT7FEzKqJrPkXKq5LjQamLJ8LcdXJmxIdM21ca81k2zDd38V
6NL5mxweg52+r0glUjLPbKeD7tsKNNT0yOqxOly9Y6WRY/Krmuyh7zda+dpPj1PT
FzUXSMb7NSCaUQGhVI8SiF7wi03GFCEe0hD0OQPLwEQ2PLzvN6p30V2eMu07aOnB
trNS/XfBlKky6wE6waGmEPptY5Bmm9XqDAurpE7oYCpUqxf+pJ4NFwRPs2y0JLtM
9MfRZsQVU8S5QKt/XILcp4DsFuFhbdmyxqKJGKI1rmAF0GBX1sBaJaXjFmQQvcEV
WYvMDlgVobOTwgx39GE94+MmERB1tzZQYSJfr2yqBNSMm+3lvoo2cncbeZuZVMCK
tszR8bkNwZ9IwksT6mtK1DFNVczX8YCnbvzBYNRhrtDPp6eMLMHgjvYbJDIoccqx
vQdbqMNfNVy7GrnQaPfjoSeBLUquR5Pz6IwRcLQHJc/zc/vslrIsmZf4E1SFRgTL
HzUSPF3pWJWNlsGca68lALmc3U6q6LyPVngEM8p99M77gnOa6pgcioBFV+stcFap
D9bStB3O5OoyID71nVGrY73VOI92VaLVLqBdbfeJQMeAxGcX+GypBS6oAM7Q7k9D
U/ZGZHET9crYjWHOpN/fdt7pcnQ3tF11cZsjjAsY5WtjW9AyVCIRyp7LmRSBeQzi
DqmmW4vwA3/kuzsaLzOOE0GSISg/U9ptPbWfJdbpRXI5rhsz29Zkvp1X0BR9ahfK
bZJNWwDc4zWy51MI2m99YWuq5JWRedoxbdrMSJBWtR5ZJJan4BtjGxEC6SfkVkfc
neJwvZrXtnJD3GHURDbVO8OaronG+4x0qhaLea8MUuP9/3wdHJpCkSW845ZbHCpe
SEWvPB0bevarWab0HmTkREmq4nND5ibnrAKX3uzX8BoPs+RdyWMBxvRwUFBTSMNu
95T2YWRPoBtrSSQbvPG8aaisU2Z1ADz10GGwvrjfHUPU52kLvpGZ+qI9+A9M2j8c
WjsxxbVTrw34koQVc9fGl8yJucsN6smXi8CcGouxZqdORlIrZcxeNy7Mj1O3qTrl
tFdc33GYYK1ocWR/OMLDKab/sMRpTz53U4NxF4Vzs9anEQy645HZGNVJIhtVNMSQ
FBE96K9mUSgBRjl0h3BuQO3HjQ6XvcD/EKAQhx+ltfS9w+N6k59pzpnwaC4A4F4a
GP7x3/9lskST6MXGisjyyA/GjgpJrjn7i+PnL/Myu9KcF2JxiL0Y3rg/0dp10ttU
1v5/OVv7aElSq4kz/hsNxpBW77IDZYl15I+KTZ1L0az4Xp+MzEc48XxkKVMKnXvA
zeE74gBng3imUaXpmt+BdaUx1WaZ2Rjz66ylbj0GvDGyAKOPr+s1PAlFFJwiIR7+
VWe6zeplIyly9rItD3c9PBi8AbjOBbIFxJ7U/PaNK9ooGTG2qqppgaE7cdi086pq
Bkm/PWtj81zh3WemfYHTdS4x7XVxAGMcGiPaBO6XkPhkUgvrohbQ5F2BFvw+rmkD
Zhjr+8Thpw0qscMQ7HsavJ+Y7hDdgsCUEg/y0ODMus6PkCE0MgTGlY4K4n3i+gPz
pj3989S4I47amXS7ZnOStJlI3NaAgmq4RbSa91/xUTaqKpf5x3wCS3CtPcDGNPkJ
KNKEXq82lQKrWyS9UBpl+a/k3X8gt7+znGCQdo0oOhdeNjP8lL2/Yo4+sfeLOiRH
Whnq89KV6s2MmjSo/IqARVV0YYcJsCmy8e/QK8URDuw00yMjXTcmXjD/a1f3++G1
jEsp3QFVJb/mqNTqepPc0NP0wdNGplDOKECYigYvOBg4KDY6PWMw7kLhdsps4cmQ
a1tYqZvi3bC2Kv0AfKfVfjAsITi0GNYtEuFNGJd7GwrsrUfHWb2RUq+AD8E5DzgN
CQlW/j0WztAmD+yDpKHFfzJ+6+B8K8J4z0QH7Uk/pmp+QLByBYZUZ5K+46ENGfRE
jCHGBO3w0Fp+RHhPNc+GeHmcp6sUgsEeQzdbQQTOOqCdyg2j1x5tWYJfzMUt+BdG
w1NRtVu8MggOEh0BK+OeY+m3nGnRgbCehuVZysbTlifWafbtBxYLOCUqamD5YDnz
ap+lVraJSbVE1HdfP/uIHUZvA5RR4lKn9Tk677TDuDhDoIsb0fs+nQv+TCFDi9v4
LzXb4pWGrltfuAiH3KOL9OogxsXpXxr1bNDWx+4AtCMqOTEWEPyR0+P/ayAZp/eN
jGYO+79uRBOVHr3mNPAmNc+U9calbu6yfNzTY+fcOO9Tyf+usdVWxbxtkAyVGAh2
WpsLKkr0rGBzrl7t/J+gjojvhR8+s2wXU9Hph5jlNe7GoieSqVkSiCGWBx2uxsDP
fvf4NFz4vw4maBIFxP3wUZ+J2JHgi8xJedXDq2NZewe0F3b85PzOufzS97JIDdA6
AzQAoBeZz4bsWkDm0IcP2otjEZeeMQOh8u583+omuPf3jF4+xipwGNa7hGRBTFkk
9XGWvHvcU4AWR4z0aEkq24d9reFTX3GRpnNPbsLFa/mXFZ1NgpJm4HsocOpg4PKG
6jVEjbYTib01NQ5w1g6FT+7rzWt83MEa0v1vU1cUMVOxo/7bsFC7lKsDqkTOXpC4
FZ2osNjrP8WV6FtiqKwk8YrJUrKEH6/CGqxgpl0gRdGwbJheCXZ3wK4w9LUPeg+e
TkTMb6RqqrEAXnLIaYhUkrzI4UwLlse/y9nhCrvMQGmdGLJ3GgvL6P3nPKBHJHEr
lpxjQQk9X0b9pK/tIwU+NVmGcFN4uIyOlN/T6fn30yyZD1UkTecFtF+QHkkyhgbk
lHKHRoZKgbuvj6zB2mqGxe6oIuAUkoiG2exV+T0l6Z+IwUr3aqxcY9jAlMWShsGo
YwJEStZR9uYeGoe9OF1+QeoPHrmccROhWxX3sDtP98PTALNKUt+FVc85aqPCo+k7
pzD/UnEt/TMq7asFnUnUZpHkrLdaGqyypf1dF08V5wBqPzbvHo2LmDHdkEp/+qwG
1KIYUdh/oPLMsHFcvccuqAL/Zq1UzOjWpoIABpjMqxEBSvUrtboiBrcAIO44eFVE
7ZIlkVfhwxU2LG3vgFJS2pJ8zWG6YPiStLXRfEQqXKpIIJvIzl6txivBHPV4XG0l
JCtOhNHRxC1vdrwkubkipwPO4V/CbRQ5mBRjrU83Lsyvz7Rue+4l1OL7R/HecRed
JcEf2bx4Ug6AhfKFb+Pg0uV1SIdUxTjt+EgQaWBX4qNqNQMm5ZGa+gmqrrQsBawr
IyoQHZxPDLucZn5eDckYKLVvKUa1E8UQJin9WtdVmXOAp2/mxsngYIrl5BJsBuiE
kwiMjrF3YcnRKeSHZwRXonFEN6lHFSBrCyDxUrzExanLmMwHcPBJYKgbRIbjYYuC
WWhNuKOksRYbLp5sCtI7D5ReAM3Sly6/sse/9wnIMGdxMO8uW840XlJG1GckELMp
OnpWYDbQrcAsQI5A5mIWfVltjaTdQpcr0CBMSDKYkhuqvuKfzzJo9tKsSUnC6T5z
D/QzEnc8rzzmmMSkQkzMl3TJgDmJFZ14ceaI1HREa/O3xokzI39ao4/PQy6m6ixm
Y0V4kKF7asuXPqSemLjC4qULsyvPkOpL6iBwfrY5+t9edBKLQ7F9+p0ueJh+MsDN
i/b8kcMtIGtUv3ylpOwSTHMHm/Dq5G/7g5Xm26sTm3xhov/9QZXAm6tB6Pm4Eriy
cHdJErYanfGV43xBUyabHGQJPYL9DB4p63gTqHRUYYh21Da05qsFqzc2cLtQIKyF
FXGHCY8AMkI2VmzJ4NJug95qnsCboTN7+XOImch7y4+VsYralYzKIo3KSewyVGz0
vCdqi4nqKUxVLQnQ6bnqDuzxAjOL/UrpbcyoN183ID7kLk5gIzL/TAuAJr6fZSq/
a0kKQXQHbh+0TIc0ECz06/A6UdlQdRdEXKxi0TJb3fj1WSMvXOJ535wOM59XfXIc
MDic/RgTQHx2j+pzG6XAOra5oCXSeFKnjAWVrKgGNyMSoVh8oRqJfQLyRe6A8iN/
Pn5zLMpVPuBFBZ1/rorX9XPqIXpMV8j8NKFzcFFXxp6M6psd1h1Z5E2iL1J872qV
jwPdCN53sflVwEgJT9zMbImLui/P3ynLx0Oe0RbH4hR9b7kzQEjxN3w9kUVwcDm0
7tHs+zmSaFdZiEVst52Kzty03gZN2lAnkG2LycgH7KLzUm/ReLU5hsBA3jxJ3PvO
zTGRI0LU1J3gVYSj04DJ4KL2HhnRiWUJfZ5op6sdN8dyFBvFbqZj3Oul2Zh1IQdZ
41BQ5awv8SXwSYq9WE1fG7WVrE+UlPgMYU7imPjzzW/HTZN9AZYXePlfuBTrpBSx
kveLQ56ul/uRJYDCWOQCTOu0+tp5DY8hxKSYSxEQ2uC4wqMxxzSmE7XJ5PjRg2Mf
w9BXWGvsF2GGM5BastTx+EYf1XNQV6dnhkWNfi/+dslWTVmBmoOYeD9hEKdH+qCF
hw6XOx8YgwD8DVqPzfhruKbh8aahzzlB0E0/VVUo8C6cM5jfItauxM5zUlZ/NSH/
iD/0/jvZTqPjA5cguPhYO3JMX4hciV+d5nJXikrQbOV3W8sg+SOco5L1fCwFzMo9
u1KX9hAQxcYRP8arKY7/caPzP9/wQN4sxSmQ+IATK6OVW2XRmjkiQWUeQI6xB38L
19XNofIP/nD1xpNyq1Zl/Aseik0maGVhuzd0qAnScVRx2xoQhRuAQlN8AdCJq0jC
wHYV9MRyQ0eBqJ9jFk3yKNpU1r4pJQ20Nkk/LRtSOxtB1DvL2EsJ33RP0OUU5ptJ
hJ5AxtwT4MAIlKU9kOCqB/AI55DQJ+DGE9G9pNp689R3douX94FfOLHbQX2d7IRa
lYEUUpAx72wjwqhG3gwccZsL/J3a9xgGuJB/PnjImUpWN58ctDfqGNAzq8HQCGgn
mADEwil6LNxh2eu9CXShxl35uPHhwrBaW8/cdsuQK2KRrDHF9o5Jw77nukz3f3WB
zVaD6K5L603SE/BqNevSyVplbIjbnH6wGJOLj1g4DFLLPsGHt00crL1ldZKGYRAr
4tjF7ryVvtHcbaffygmu82C6KjkzaBAqVO1Kzp0/YHvu33wwerVDvwDbvtFTuuef
6QEGtLzEXMD1orBbePlEwz0cYqBUd3uTxZD58cOh/cxzB41iZVM6/gPk2MDlBqvc
yWwLTiQmc/8Y5XlATfzQcJ4e2KsMhyzwvlx1aG0fawfvHin1Q6yt3ShazYguyZcq
w+uA/ef9YUCJMMyokt+tIGbFrJs2WBjR/RfgsjGc7FalHDkIGTLx6+fDcY1Qllw1
qdGY8cxNtOa7lqERoZqoHBZin1XC6F/9uhU1FKEBGu2B4ihYuShgnprcGSvrBF7I
xwRnUMEwm9B9j1H9k3vbFjfgnEsP9SH8DiTmVrkUswB2N/uZvkQtfGc9AAXHNY+5
XkZ3D5L5mjvBVZA5lURC8a/iJRxQFp8KJ4Yoa6QYplHZA17+RqvSjBVWFJl4SlyT
+IfYhlhXre2o+u1FgbBw94g+YyYAQlfM4gDzy7RGbEEippu07eKEdBFBJjmmIGn0
jd1x4WqT8lfcpZRKHJNpXg8NCF0OME48w7MAqViXuq79fjCQ3mi+2dsZS34XF4gN
YGNVQYHIjMCx6zUkHiJVRkl/PSs8buLBDdAOBbdqEHRqjwsandF3W96e7YL+oLG8
RPq0sYoMRP2TC/KsOdvnijaeGVGV1hYVHKnP9oiKzcuYkEJXHqufA47Omee3kp3z
prb89FSB7EvAK0GROJ1mFGGy9lRhU5SUWNkEA4xmFtB9JG5h7pOf5mAaH6IrN2cI
aTKa+Dw+aJNlrO8ClpA3zK4Bwb3SPZKUas71s5Y8ts7/W6lmuggWi7sqe7ObmZCj
Jb/03x4tC/cIpEg2ME3nNumgwVaiZtTRVdNJIhmF8q8hKljmS6288kXZsRwdxB9a
3oj8VQDy21Xq71tK3ZlfuMyxT+72ff7nVwUdOHMTtJX8aZAGW0YiZ2F9cb20qm2Z
/kG9J006CkiwqZCqkHtk2ddpc3/Rl0IR2+V0fy/rZSDlbxcfRp8+dImuQXIHgKsp
1Qz1kOTBvATJ1VMI8Y4+c8vjmtOUxQlTZWf6saBGDby1LeTtizsWjc7oMaQoSnAB
iQs0xFSUV4fes/kX89lGPlLau77Q8YRKkJ5/1bx5+X+GrbYphPLqenxyRxwN3w4N
68+ZIRlSoYEqtlJMOzxmPtN8q4iSPaiR09scgfXAunP0ZBU0YV72qTrfx2PU1RxW
58VeRwGS8PctyT4zanp2HxwsROLXl/F92Ukof0RqDg+05Ip64cEOuKWmTOaZtaLi
ZG0jld5TjZIsCgZMDruN8OaKMstX8+toeU7Sp3to5lqdxCJSvJM9OwhMcjbANpT6
vrfw6ObfccT5GsuwfGMFxsR9z0Am4TFyxlxIO+9WO1/aigszgnNzteumevdUy524
pIhRZ7T/xza2YXVErdIEJNnfOvzo6pt0ROPfjzYor8sCdvgy8RCCWqmNA//qDkNS
dEba37JbodkHLGs3m682KjlRhyU6AHQvvOPJfXJREW8xOB52IHlQjcXPakfwmnjF
kD78fcmihnVehTg4DqzVHUH/7qKPaL4dipIAVphXbjtvsKHdXErTao4y69RC2tdw
JesaRN+hsDelShdQ28QF0Z/VdGTuuwt5oJkf28aKN0kp6qKN4StllrT5EaPCJnBD
rFFlBANmN9B/ENS3DNkIH59j/AGoa/PKXJsnJEAXWkEFXP5wkIqwAXoLG0YRIqqp
YBWucqA5/j6nozX+JZCwU2AYA44E05/KFx5isEhsIwOES057/PiX3Nug63PXiFP6
8ZS9DbciDAeNNXUPfGbQ4temyBzcQQueK0C3wCwxMJx4sSGiBmRQ5PVGBxrZt7aR
3jbas8E2cppYgWAIiPsazWFoDwxhkwWQA959Y9lZKiMLZ8E6B2Gp4n3VPjUcHPM+
2aetZVkPdaMIcX8hv7yFflAapS1TtBO8jFipAYYlWV4U+ZzGRxHiVsD2Z/rcivs5
tmvecaVESicTHZdttsMn6VqD8eI2ahrOoMz1y6Zob5JZoqwIn2KLLsbk38OdMlJJ
KDPFs157TlXbuMGkiUe3aBhaVnMo2gIyc0I1mu/g4pwlOADMNyr27+NWPZquRTRi
/y0TMd67pkH8BNvp2mbJQfkKaFQnBajUG9gm+DkAQ+PmBG+fK53IUNqTj03LUkz8
xGsB755shiPfaD8l1c/9FdMPyy0Ylfg8LdRjt59h0EUSGey4lYCfxEka19bOKdST
gVK0irYnPU/Sdhcfo+q9wcvt1/6h2ezKi0FjwuZiwGX0X/QYxM6kb3SfmbZlfR2n
Kjhz1C8K+h3rRZllin/iRbCR7BreEQ9vgGFQik/rV9Rv0Ul3n9M1wnImM3q9IwVM
TQYcG4+k5VAyj9a5aUktR6+DM9gxyLQ9CfaZcB6AIUp6gfFksVhh7hcqc17Zb8hS
4BhPDow/5BYaHq5DrySYZgxHoxiC/epLykL3bu2DNAWrR79YTjsBECxsgCPmYXxt
BK63okjZ+WCECLxiavnAJRqHok9EHr2DZBjqo8PEyS6uOztuCFhgTDN1vLOVsc5E
CrwdycD6jCLQJWuW8k/j4Xru/prdSAoC4bebDWKD5XzwPefF4g+FxDi5mhZfn8E1
QJTM2O8ZVo4GbGMx/TyvtpQKVYzwEPnc07trOoGg0aHku/JtMOkLWQIhDnDZn8Bp
a2mHDjpgAvQ9l9MVlcUehQ5wID/juQaPG0JA6Oi4AQBcm8n2NZ9b+hBGXQaQJsO/
o8PgTXpiKMxASApPTSCoV8esNAk7mjef3kaI03DSXzj4C8eDnD7KTuuGyJw4e0yb
agO6g2Z293JRZ1rH2UbHyivG7fbnXAk+CmG8I3CDlzg2Uk8xTPDX6xhvZJSpPcvg
cZbU97/19Eu9Ce3if0iw1Dw41pJJEjK488c8OxLB3o6EooIJMmivWwxHzoTg6Es7
p0TkZiIsWswMnWQpv10h2Av8CkGWJQ7l34h1r8wUO6je8ddS8HOo69ZUR2LxIy9w
Utf5hm6JjIKM6oUo8RBL0MLx7pqy+x8wcATmeK87aZjN8m6AipDBDV7Elrp9jTAb
SzWK9iINeUOODUMY4bOJYqpwTAmqhEdhE8wpcJxjbXhWt42dEwX0HN1Bg3HIzyic
Dghz56RiUMLQsRg6q3zUgXysLx5LulPIuNxIS5S70irV4C/L7VoCQIUDsXuXWMM9
SKtHK0D0Y72b9mAWdyNddLZ7QinzUcE8Nb41YMllpuDkDfrKj99Lf8IDm1VWy8IS
iS4KI/Jm68O4SYTnPaZn6xYEWOB4hYQPHtziUGdc0JYFpoIkBaGszkXjNsQWUKlQ
P9gM2sQXg9BjnkZ8z+qUVVpUEjWzC/BZJqv4HIx2jV+2DLlehgL58f4KSKo5xiDh
o5GY7rUOswEaeV/8K8v7GLZVdLPhc/IsqG+NRr8mhs33YRT0HQ5Q8aSpu2SodSVb
rVSa2R7cIYGhQ9ZkFp2cbNbukk2MuAt9ggZ9L0rrDXCsKZHtQc+XrCq3MOw/V85s
QXPTQMVEMhUD7MWI/rA92Ld33GGNLV0Uc7NApCZreBIXUJRcIIxxZYV++NpnVIQp
ohFCN7+q0+uv/4HlAmlAT6yKml+vo2j3CAF7xESzh7P4kdlPOq9+p7R+lJHjZGY2
2YsnAnIBn/q52HySzhSYsSdtPnym54afPnHqM4PUa84IotcJYt5Z2kSVzLjRBKGP
Egt3fOIsqi0VqKSge/MzBwpmSX3r1XbRxyuVTY5LHB6ML3SHdPdyaloUjwWkVJsC
a528LTEqoik/aZgq6C6ReWmZ2zKV30Otc+1tqEp2jI1fsUzR/N+FYd08bpsq7CWI
btuhLgesaqVGOlpbBiXnlpB4NZahRJzsepYe6EZMMYepWy72G8BxY3glawdfdDuV
g7VSQpzcHfHR5983Bbv6oF/fQmkf3jCnQw7Ik2dTJ5tkjjDWlyy47uHvQRxl5+P1
Xsk+F8W0r1lVCJ7iF6aH3rMq03HuvKzYxJ6NW7ndk39601r54bYmnOs0h0AtU+//
C+6a4Ipe38shj5ViZerD+8HLbBoCAu4nBpsoSeDfxv47UdsC7OOY7U/L05evbxXK
KlWXivy0lRKc/WMHAHfNIYKxAnWPyh1FfTvnqlxF7k487h6zGl7F2UjkaCjsrNSu
L2H9KdZhaTEvCNC10LtcQNxwEGSOsbz38kPefXjSs4HJsZjw/F6CtXtolD4rPLKJ
i/UliJkLs1/snakRIx/2zExXfHxYeBAIwADfNTfm+7scscRrw7z3i0A1qd5LeNSN
I4u6wRrl+hikuHnyfemBVDA2cIc3UP/BZqXFCAidHnCKN4zWZLm8r2s5JR/FuHrZ
H8UnDrXnASQTG36bw7DbOPPnTC95PzlphxW3HG1x21CPHHGR7zFIKkjyv41NYrEM
IIBLBOHmPd9AZ4OfgLkC6AeWbiPy+S2eTOyQMP9O1U1un5tlX8s0IF0npGziil5b
YsJBnSDqGIqzaR75IiY4KDVNDyOPCmAT5C0nGnGOj4BSKim99hllFsuJKND0la44
CB6JktRFZxUQkP3UbJ9nYsRXiZcI5YK20Dqm8RLF/KnF6Zxg2NoVZvQQPZ/ioPxA
RHUsuii8XgEYoQUmTS3Sj1lk4QjbD/6P3NMs3URRsFk+c+nUBgXyIka5+cW+qZEU
sbtSoDL3Jx50mepIBcRT4cipLfEQQybhwo4qO9IZi50/gSmAiIna/CdPrrRDqhLZ
rM1MMKRgJB5cmRhd3EWlhBvaTZ/TeDo7oSw2F6rCK83F4w4T2dMB6EkG43mUyvUD
FVIs9pJKrSHItdzXslU7TkZbvV2i/Xy4zZz0aWJzkD2j3+yXvZj01/7/q/lJI0nM
n3mOMxZHUonFmUQbn5bnXBrNUCJQf/JWbdcKcC7qic1qg4cGUwrRJFhkP29Zw7cn
pVKsa0l2CjClqlrrT38sAMg3/eeo/29IStjlbK9E9Wk8kH+CbqRDg3BekpApS/sw
QLi9yzkCRPLR5dVy62bP9dSCN98wD8GlCLccVpbmDbtP1gHQZ3eX1fQ/K8Dc+K7M
4NLB+xKc4ANyeVjCrkbD0YZeN0e1LN/8tIF/1os4viF2aPU+lPxAYtZPm1qI8kki
LBlmXJ0J8M1MtzKTScq0X8CN9QW3/aJy4gAwg32laILpCEgyn9s07xC2TK8Ay0qJ
+Yt/bFDnsqudoPdr2Z/+5p+OAQfM3giSEr6N/vRd5XqKnuKWFHATwFsJvpooRc6a
PymjuvT7RTSmlNigKE325Hcs38cfVwiTVS2Wpvo1aMyyxnEbzYsma8dgRNUBka/8
48A3/NznUPUC6Bb+vppkV+FdbKm9dQD8AvvZZOoOed6xWGOGSkG7PuZCsdWsHAEj
Sf/8Cy+hCkZgINyC2O3VfyP8kVSx88iHXeUZTYnHHpWqefVHKsCRG6/GaGm9eLAI
WNOkJYJ10YON6Y37WABb4wy4FpfBIlO4pjC5Rot+LWjDCYTKaAgMKUEqNajMCBhZ
wQM4EXj1kRUtM84RiQthdtIl1p07v3fyiciRlYGbGWQgRrFeuwBriO7uhCeFZJEb
4UVQG+NlXR4rulaPPxGq7Y36P5lh7qPSUNC0xEP+5n9yRIKukbneZRlfZeosoNTQ
t1OBTyZ0XKJdNXcbQ2NtBtsRCS2YFKJmYWSgV4SFHLUxtFa2htJU3jdckVr6lPpK
DOB5SeJqoKo2mVCAcg2fpTwyqqbAKOKC5qd/NWYw9yc9Cv17nU7C5l/AN73t5tj3
UO4MAWL6CUYrdCdhxD0LMwx2Etw3slAINXp1hdNl5q0qN/wbk9IKi3rZO4dUqjf5
aqBjBCM+inkwVokFerHpK+zIY2zFGx6j1kxmQSGNKH9L4IElLFwtmjKzB1L7mrhF
lRAkDp2hZD0sS5FW+Lge4FtYAjMpGlN8Nvbw4kCJHlyGTrGvx1vgQtsglmXOvbyd
HyNie56yzeTUyd4QqXWrFrDNiflgw1e1QzLtteg0i1A3acfaKtSBzItq+ORdrLd/
4S2rigHsPqqBUkmPk/hwzClgoDU7qYYtpD5d/3+QPqBce/YX2DlZnh5D2rLFwYD3
0orQ0JOXhz380FNkrCm/XxHfn4qQXc4GQk2XO3dwKwTOZYtS6yHS/rq9jPwQShcG
acZhZ57UOBqDlDnDgehdCpVxPUGRX6TqeHHASm4kSNWqaNZTv1ryKQnSuSeX3yXh
gSyTF81pAaNpI4/9w3IcPibcNx2xlBMps/8OJplHFlUSvoW/0rvptMrLxLj5MXAU
l7yz9mQWigTA6iVCNPBeUjq18dTyyvZnq+u6bl4dZBKS8leuZHj065AkDtwBytlD
9zP7Eg7U/bHzrBptNPpaifysIIXYySdbxGUgvAPC3Lm6AXDIJ/+2TbKHAEsR/bh2
z89YOc+D0NOH0jim1JHbeSgjlQuvIvs5JnC4GugMUvBZ2tz+icdUhs09FOoR+cSh
3ipod+TEmRC2X76zEU3MiNjNkvqawbu4WkgNkGBoq7lh3XqALV6yQVwJJhXcCyYp
TfU8IshVjeec8YzzUS0vc6wmlhY77Fi3gpElIz7RcQczTFFiFHudF8M4jduhpfIg
cfd1DsJV5d2U7mQF5lxMXmiBivQeD+dhPMWidHhku6JhbrVut5+tFnprPaOqT7fs
aengJNnGnrya2gjvIqY54Fg0rVJdP/VFYa62GcJGih/vybZl2Cn5sj8vMWiz2ECe
Us95vXUap1R9n9CN7hDDMvWw+FqhkiEk72PjGaw0KGyrIjn2NmkWeOpvKUuDPAdu
syDte1qZdHNauEeKfCyvoNT5ZgYACg4w5tcvwdMIsHLXvosrj6bh4ew31n/FBeS1
l/yuIvqkgY8ShQ8eFZkXZybeL6KesNV6bJeUf6mkpwoERtsn7uA3rVuXQ530rPTv
c3j7lFvNmPIEVRpQRfhYEo3CA5jCe8df992l2WiUN59XaBd8HLN0kfvcYVywlxth
d3ApBQiGPrg+YdIqvX62CESg+XrRuInl+l+zHLVvtsQtJMqITt57skIt95G28vSR
eN4GjGM1ZzZ1L2aZDDAeq8+jve8exEzrx0NEndHwW6nrPMzpaJnIDeSPx96hvwVY
vp7NRdxvfchDaYde0GZijK4lQJk6xaXk7lbgMN+D69nFiYRrUh6QgZo1ULeSyrGA
F61oKcOYLs4ehj6SGiJec2fZIw+Dn9uM/anPc5GZ35kOpF7B1X0qMws3yOk9ajTs
IVTu52DAgtwA7QCiV6KaZJmiSa/pb4ufyTx0KOxfH+k1BoKsr1PxO6/Vns7HZMi5
XEwk0S55X+XRA69qms/MTuYgOieAmurgDMfxdBBz4KkX/PO8OKgSRTYZ/50gDkRN
IdPMO4EcQEGc5eeqyBC2yc09KBSSQIcTzDmfslkoPXgGEPzcAkl2GzuypqhzOlBA
76zaFWO9FoxQPvLbFWViJWV0YlcBiMnxy/mRg/9wKroYF5eBBxt1aOgS6Cduq8SN
aGeywJxcOG9Kg+aBW5yrWaeY0zAsdAO1ZaWPZe4qC53cSI1CweSiNZzLxuiTuZto
iNFTtj85ad8K+mdWGdEQWagkuEaEFYQaxeVYzebwdVjsF2fiOyGM0ZYAgqQsBE+V
/TWAEMPShmLbtw5VzYePd1CV4MR4tSQV8/MzDIQe88ZIxEQXjbk9yPDzJLOqnF2h
vFBHPewbEMl4H2oWdFCBzCW6ZKuv+4udTnh6/43f7lyqIUohKEIpbiiCbWIn+fqd
4bWdlEKcqnDlDUp3iu1ioNjqN/yObf5fu+TrHFsGRRd4j7lyjE4Vg5IfzC57qwNX
HYb9APsvNQ3k+0UeR4nxBu5K3uPbv/RmayBByIlqC+DXBtXg97xPMxwe9IuUPFZK
gka9FlNGpn6aND9tg24Cmlgnj0WppSUqmHhMSZ+Iy73gMaGHU+SRo03301L8BH8H
1saO4hOAPIb7GjBauh6paFsQgT2u0NvBQIoejy2wRGW7UTdVQDouuu4fVZBkgMcJ
scUdR9nqXed1y85BQkAacZbg2yWUHoM1qk4DJIvESlEn0ABgC9UgKDbYvp+fIeCm
Gbdqjrs5m/r2u3KYUWpVbIoybd+vlVOACRd3BbCE73JQ/F9abrZ+ssjUAXpGSifd
9tvluQriLEHr58XoJrbxnFGwzUGYeLsuLa4K7B0aXwqu9fESlr4nfN+ccQBLQcze
T1t8v4OHlsxb9gZPGloBojgT6uT22Ybiq3XKAGNWWDSNROdB5TQTB53H6PKhJMwN
/7CYZ9FDMvmmHtBViUNHRKGFP1A4iXhfmISjrO9ZmEqdz3FFWRRKTfyD6jmqNkH6
TQT4uoUNQVFBUvCoEtTBOxMKH0Yd3HIBQKAyiUDRcLjE1pBN/LH/UQuT5LoQhfPQ
PLpyQsUpdG1A3bm6Y+EpnOPficb4Xo6YcXwmviEGsLJNb1Ziwrr14ujTnup8a1qQ
mvogCbssZ2r9Sjt7+cTNlh3MHkrnIsf1mu+3YJDU7BB7Nt5clv4RT7HhnbV36yg/
mj/+Knv2R3ewS6SFNzTbj6kFx2B1bZXo+XFtPfYD2JN81am7PxVpgBdCKgVMZPXN
M/F+c8hIQDyyhsd6q17hI+SZycHWSJgf3HpkbqtC285mmmhSDJ3ujrQgtAJVuv1d
zsOAFLWodh8CQROyRI9cfo/RVu+aBVM1MBVy/phKrvTOpOZTpEiyCniWIIxEHD7u
t9UMWRf+1/kU0+NsIM7xnb+Nv/IsA09Zi0425Aw1GrktY8t9RIxZ4ulwi8ER9YLM
kfPT+TwsE+u0pMTrpJWomLl9Y0I843xnRui0Jw3dOzc3coG4pX4EZDAjQLYqW8j6
hAH2SqvzUrnm+UfQOl6CoL7iRIJkUgR9LcxSwJbRoa6KXPCO251rRw89bNDQyAzy
7L+gATedD4n5IPqXNuBTf/+vqms/Bf+pOEPGKWnl8+tTayuEUT4FJL89NnBoE0nx
/arRv9UXUfm0OytTbUmQ6pFei/orKzC1736uHWNVL0Rrn/twASbjq6YQ5M2gPYm7
unBc4Zhh6iDvHxweWQa34VWYIOvmNCOYmWCI4rHA+9QSTirhcsDPsyCEQfBv1nRw
ryfQimfNnMZGCMheOT0F+AafFoY+7Q3KaQ8oxB6+Us0Y0tjjAApkgI8p3slZ03Dj
AGsFRIVWgUgLEU22uGtd7KKrXx3u6BO7WRmBfbxaj2pzFfiBp6yinMPYaW+4Zk7n
OlrL+gMqN9dqnHuH38uR0DMeaXDz3wLUCF8OPMXw19R8mPJ15GoFH/t8t+O62E3n
uvlJ41R+6bdUYupp1C0qxPFKtg3AhmJUIwuAET29v1xn7bGmXqUqI5SJsi7WTU3T
kn7qAPnPg11dKKTyhnLvmnxVw0wXxRY+k2fQzA3NwpPgciNCGIP7b3ZF/ZJ6jm0D
LXNlsMKXHwLK1kkPjFm9PqfaaOuPVTQHXZeAXEWo2X/XlQ8V8jkIKiuZ0GCJ6lrM
qrRgC05RVZLyuL3z0BJpU5DPU+iRWO5w1SvI/wTAwj/cJDD5RbcI9TboIKo7kxaC
uHyUEsnuS3vTiCW1hnrX7wjOfKtKfECH3UehUiVHOSxy1IQPDCevpZdFn+qFzUhE
pCk2jWg8n99kpBf73841atKMIo4WL5/7ybsz5QhBWzBxt00ZbJlhWKN/MEejEfZh
lqZZwmRiijUMHUrWac0iaoGuYyX25+9QvPL8zqlgT7aXrRjUKPsh2hA8Hsps88Fw
DXwRepvSkIgJNxUMHe7a5HJ93wH2+ycXReMJl/9JWor9SZh86x266kYEY3EKTK0H
ZHWNoOlwxhHTqy0g/tfDrcrmvBCUJyx2xtyXZM85dCH94DyqeMUchXAZ6w8T86oO
3rh2/GLuTj+UiMCHlxpJD7sSYpmHn6eowWVEBsgIH7NzY18DfbAzgi3aOm6j6nMP
LTWgd75YfkbtDanLvLe5bTEPGqxkI0s4QlmQfCwPQAcdOTAEUcUwQMUd4bqYRWkA
wAlbsATcdVybVdbIgpqxf5CuX8XxyjM+hTFBHp71BKehPDEljvgCqQ2SGZf63+Wm
OZndUTqKh3ULmi7FRLUjpAKcxQh6sQOYzDrnuXTO8M4CqYzFwmr4VpS+Jmdnpgs6
DGnRJpUcmML5yd16HX6p9AHJ3f5FOjTy76oBng0eGdPuIJHMN0kCQlongcqIhRBT
L3u1da3Ig/mGl8PFQVQq/tetzQeaPjYlfy92i5OPXUHZvyI0Yx9BkwUzbnJ122Ql
bgFHTfUlQrmzEWf9cra9B2r54RLed7jirPBQa8xIzWaPCQ4OP6SUIHbCyM+tz9iK
fYiit0ZwFB4PEUp/t3xNSt2Nbe+imU0eB6ecTiAPtUuuVZmcWLG4byYEQFWKcj27
06IwFw0fG7O/RAHe0ybiGLvmykcQ7cEhx/WcfB76C1peUgeEbtGZ7DeRSoKPaGuN
VxXW9b3O9N8l/Uw5aWLME/jD6msCMHNY4pC+p4i35E1HKpEoTJTo4OAby4wlpUI8
JUzknXNqdH6psqpMpbQmTDgZyKh8ZfKI/icEaYoKQZAShHtShzTw5gEvUR9XcLrg
kGHfhPmJTf2WlNfxWQpgQs8OKCVH8sa8etWJ6njkBWtEcnt6myWbJLEepczkb/n6
sQ6wnOwFIwSgiGGmb2/fFXug32El6nfPDILGumgJY6rB5SxKOSJjAe3dFuvTuR68
ZiSKTJAt9rzXVWWTL+eSKY0M6pYDRRYEcHyxuKaAziNEVA6xYWwfWPoAul3Olwmk
cHS/skaoHc/bdZr2nL/VtY7ekaQ7l2Q9l5bTghLXAeYS0wuxdS2gVI6y0ax9Uk7g
NR3kcuKa8t8MCw6YTH5JtZlHk8iIH/EUIE0J+JrpJ6C7+FhgC4Y/kvmD9rIH22FC
cAR+iLJpdnSL0alWFrOKnFBQYedZUZDHMDpuhsQIp3rbE6mbaPtMRXpwSgKYBI+o
bWvqF600zyvqodT3cv34pHiW9D1Uvq41HKGKV2iFDJIANiKrGtscu+UZAoj2Az26
6HGlax9aH+FlNFM/zE8HQj3sy9ViHBNdE35hMIrXkmIfSLdNDR7DMjkVemW2mNfk
8SC57sqtZGZyjeGpSlNpWzrEguoIC2GY6CvPkbGrAqcitVY7MxWaSyh7InOnqrjZ
TkTZJh2GvU2ML9wkyhaNmsCZr1kHcdRaHmWj21M7Q+83Nokxt/RLCnPYOGkEjafG
W5N4ZA+jrT7hLtPkeTgB9qFrr6/ARRozinFbH0nc9d0kyDW08p+gnvKWTsAe8PZD
9+hR5xpkKZYTWmo7eeE/wd2YNhGgebSCO7so9lbUA37xYh9AsauMKyRQx38uMDLD
WAVPFSfVu3iaubDt3M5DIXU+SKHUvz0nE446HOlbYoBXNxQx6mADybk4mgt121cH
3CTxkDabnSFezHas7YYbpQ2FsFEGeNB753uY0JxHpPQ40+IOsVkNsPJ3oQ9ucUaG
BrNnCf2Ip+WLCQPV/Kx30/d6JPClW4usoYVc2A5l9yjYfz/zM5HE2DaTK+2Visbi
YB9J6IiMlcDIXn4XZ41k5XnvmdquxoJPk/Ond/3fbIhPUSufD96JXCtuFQ4f/Yxl
aH/R1OLnKarXPFlMk78axWMqM/nX7Dc96WKm+CUO1J+24MUvfOcqclqHyB3H2VsC
lJCAMOqO/NSBMr4ImH0KReTQVy566qZaqi3dQI17nA3XTla47nhQEhJhzqe6bKCE
GZFbbxZ9MWsEPzHCkxi/05Vq4VtowGBHrpZmjf6u0f6wentU0n1oPMKCXMUl1M9w
2hXeLLZJquYZLBW49fJWlBod5s7ZXiRjZJW2YFpMQod2u3Of4jks9/uowTPwb9CP
HfYvpaQQOW2GVwarNn2/cMhBBZFk/M0eLszfRGxZo//XUYYqn4fSz1RP/mNJIBWJ
aiin6lO4fRhb7P05JN3vU2PC4OBb3uvDUSFKghP+iih+B2Y2kJJQVVXkn4tVfhKt
thkBIewnSmKMSM5ubmA4dEspxmRbQjt+ipaSS5CfIUitBN/H+GFEFFUkcd+rNLp5
G2Sy6RnuEhz7hXrS/FOgiFPOMJ7eVESd3lFJ0daoF9y5MfelK93VI4P+uLALCuQ1
PRX9BN98F0cQfeeyEICBgTRowgwzaCcXzENz3lGrmS6bs2dVVsl0Hcaq/wDxaBTI
SC3SsVF7oqJcaVRgRDf028Sftz4MJqxSU/Qk8ODBYncP1EaJrO8BxAPZcOzzEC8Z
ekWtxGrB6Dim8ojbAvVgUl3jHspzmNbWvWJDno/5ViCTbQIAZhDFmiHquo25kMn/
LlpDf0sB2GEguw9MKlcPYfb2LcvDpsmfKrQSLdjNjzCgCWvQL4WOENXTgfPwW3dn
Rq6xKxN45vq+oCfnyYb1eNmLM9yDnLGRodizyvC6rJdKj/n+PFLpSIU1TJoRrWWe
rQ8Q/u6OklxEzuFtbQrRF9zEDp2WbAL+FJ+1uJ9eK7CjbQ8cFWWeXAYzfYgNHjYi
1W0y1IoGycqG23GTLrWyRFdo0qahXDGLybhW35/3v76XfP7ChagHDTSJ/YRxRhGG
PfSeL70RUZi+ThmUxZbDqCk2FKcCBsR7+WGietqI7vbaq8BA5BGS0y5S6UjyvaJL
L27/3b/g9TSPw1N6/QMrYmLGd8EDR7R+gyXFD1Hef082e+ixc3NbMJdbKh38zg2t
IXtCEt+5YRHaiWKjmpQQHMtkAFsnJ2ThsG+6hqXN3aVhx3HhWPZKL5hotS+lV+mi
fKiUCQ3LJSh1lFOIM/foS4GLa0qD+2XY3HlLFH94mWItNMdJEtyGk7HSGSWyWlaV
y0sF8+VPMYqjMe4NcrbGFTzqhNrLnVh/YBUzSajEEGnTA7LI28y1GAROjBohyVXt
K7xGVbDL6ODVWXewiI6ZtH9jvthm8G3s6JtQo9lcat0xIzdfzJvSKu4qo6BzJQFS
CAf5VuRChVD6VXC982n8SC2g1BKz47MMXJGhTGA0XEqsydCZ8rjBigVA6ESKJn9O
M1LXBwUH6aqorokc5BcrD4oTL3ChKkdGy7CrwMxHKoM2WW3uYatO3gXiaKlQ1Lte
EI/NibcgQb8ilqr3OpJwCd9EYhxlJIRe/EYOTRVSBtFPgyGwBp0tw6hj/9C935mI
PMcWCVNaszR3RfD7ojcoZXWYovxpY9LmwlfbZY0kpJWmWw+ry/sPSND/z7cpmzB0
swyEsfs2UfcKAKqrW33szentRiU8TZogc/uNbbT8UiMlNMSlrONFPjOXZ8Ex0xe5
YyLvO8QjV+WSTcqPiNx5x/JfbAr/oQd8fLLAOLTvswLJ4L/mc7PnUU86c+OpDbte
JAHnXS9rbp7249Uh7wcV0xOEdXnhlX7mFDBaDUxjXI20tCf+SeJuP1iEj4FHA/Zk
7Km567+T8PlfyvVEV3Vo0gC4FcvnUTwstplPUHpQ+FCFhSxtCW4K5c/PN3o5C0iO
pNCi4oHrLzsvPVqdDoatP6wfwskwGKPkpa+/Rl+JmucrD7zQ6aKrFKMALrteUv4s
sVqHlyiSL7FqHRdePsnzLARRAMhdNRKmXhff72QGQJiH3wHlyoyWEXlYm7LzcWFt
JmghUyK2+kyAKn2D3ETqsgDZdOyD5vrka7EXT+wNZ3GI+R7mD80ZlFRjIggt21Od
N+T3nQuJwFGLpRWzI36U7RQ82++Nhj/VR9nT9hPxAloSSO+TRpq/d18bPFMYqX7n
tAZBNYKgIGTCZk0UDo0iaM718Q2+pp34ubky3oTAyJ+PfBNVampcLnLbeiv/Gbcj
GkEi+WbeYH85KUezvb28gdk53FVPaidC070r3kebmMXZL3EF8GbqhTH8OF//5oVX
qXQlpIMWCiar6SxdmRA5Cr/7j2RoVZgQsm96PouuhHbyJSfpOjcFwEs1WCbQ79rK
K3Y+/smk8hEFe1AfftP1lZNXlENKCSOYqTPiIUKhem26jFgwhCUJ4gJNyEMJ9aLH
NKqboPbddIacd9/5m48QwKg9VN9MyG4J5ebl9i2wYsMJ8YciYDL/sQ09okK69hIY
hWMklSWgSYYOhm+bTI8ECIZFOe/mFvdshVrx+e6MOvn2yoXyzLwu3wIMO2K6BrfL
hxwH5LBTKZIFL0qM/ewG+jyJ1JCToMjjcz4mNVE/5uLIe1uI4LVhv8Ac9Dv4+mtg
LGZSs4qR7bblYVKj0OH3ZlDDYse+AeB93E6z7xJ9OgLhnj5P+4RR9ODMGGfNUQT1
68RYvs8utNowD9Er28Wr4j/LM1sh++TZwIe5pgamkkyzNumHhWvB+8i9bcuCDZAb
NQvUMTKhLq7K/ROWSs4WHT92j3/srS501k1GSCikmEWU7PxXoVe9TMeWg+6wne5k
qDg7eGHggRs1W0MR6mQO3JVF04a1QWF1vBTgrfb4A+Rsq203Xa1v9o8kjR9Lo/FB
t5CfSRMARCKBADepYby7doJGLZO3GFsCr0iyy9OF1xSph3cBzXfRoDX+dHS658WH
OEIgHgzupn8J1rUg4cNHjEGJ/BevWubLtaJlvi0tgbKNwYFXWg1Dem7LtSvxwcfo
`protect END_PROTECTED
