`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C4l+oxzrAnjIO49UrSm8q90b4OzzwppFDZYXGigIq0RDXLgvO32WZnqIyg2GqhSA
7LXu1V8J1DIZ14eJecucTY7RX8Hwi+EDor6OUNPbk/9cRe/YVgCxa1Hw7PaOlwYS
SgRtMzr7eUEJeJBcaf/DLEUHidOcwysBPUoNdEGJQtnWHq0JhspM9MDAlZyetx5I
+Q1SY1N6KmPd76XZ5YSjc4B5ft6rtC4Gma3RWhjQBax88AQGJOsAKrcGKc58rfxa
jfkH+JlkrZv95uilRX3g30W1N6B1MR+yweDSq65L2Y6yTRzuftwcTmpXjkQntEfu
Ezoqqkt5+S2jwoAlCKdhHX9+cHeA8fBf469PlwJb/2n/n1wkTFJHkSB++NMPJy9p
9RhKEi7h5x20h7myTXf4LjED4rDap4k5kosZWVYgS2UAxLmCngvFOmYSKAO2QRlW
UPlHMza/aEddKDJefe/iKGAGqQ0ioF9byJLl8fHkMCU49ktJqjdBA3jBhC6XFw8K
LSK5tq1b1K4dGvMhGV9w1/GMFbp5cB7O9DIrX3yza0UPRzZfiUaMuA96XXHuvz5d
wnaZF98AMpaVBOZggMDHY1VCmwS6lL2DR1STaCpaG/mpQ9W+xcscQq3+S3k9jZ9F
9JWtz05F5rrlUGFMiRv0PXSzcAfYJdm5c8IW6wooFu0naaVV5H+Btgj8XqU9hh1O
0fW+p97VX2Enh5qDUzd3fQjkX68BSnUhgCDNYqgEQS7TDJc4f1xt+E4GjDc7QD1J
T2R4aNPV9mnpkZWR5QdEA1747uD+J+KDiynTWJ/EKb9fl0fPaxqzMwahoUbOQkug
C+9s5kvq68iYp10A6n+N+/8PWTjfhHXwczaj1tQ2c2KrxIu8csLFbkw0NCgUf1zG
/f8mYCrY6dhACHhUirxdli3wCP1JgQriut3KhJS21baX7yKpuZBiXTLdXTpU3hUd
Vs8DjqU+N6V9ZcHZGQHSnJ0eIjwQRJSZI7qCiSf2H91tJaPUsFsPbLSeGmpCR6/4
zIYnOxOuopGv5IhF9oeIFS8duTkSflecxOaZhP8PQ9HCrqwkp/elSWi5GUe+gWil
ONdiijxhIroQ0FFxjvh5mMKOejH04XiACEnZX+lskMxSsRTqpGq7aNSuORWWq+5e
d5uYxWlWalaL0hRxXQmx5is6JaNv4F3dHoL5p/jzvn/KXPNDBJwdHh/qTZwwht6D
NbVQGGKXCiUgQsmAu+JAcGSi1f2d4kfFjFCynv1el4Q36GCX3Z2YeUEuTaCWhTVN
hb1aVUAumiwkWLDnGXkSu4DzyMXTCNrTLY9q1ymS/hmybtGAncTa+pSs3W4kyher
B28JFZG6wypvi/kv3VU73+liYIFx2zQ3N+6n6U9fkXv5WpFX5Dj89z9nOVziWnEE
Yr8PXrycIOrEqFGHygRlgbkUc0r8PAKbsKRvrv8qiowv7Wmqhn/xKjBdclboZlWJ
fZP3WZ9QiMove+hDv+wtjjSC4lsJLBn7vc6sXGiXB17WgPiAeXYh0z4kC7uYByc6
gcS2iqHJMvsQ/IgSrT2lOHBiH6WGOfwKknZ8lG/bw7LYHo0udOpVdLj7CtLZvHuD
DANpubffZT9SKuxpe5cuU2uIc0L8Y17KsZAA+6+nOMH9/Ti76/9kiKTUOhnhihiK
1Gs/fdqIJBARdS6XY1mtD6Bc8LgImfmMtP6nRsCFkIEhlJXQzvD39RouBw6BFxHh
yMyrY3TbFpJQ40mY+NrrE6CY7Q3/VJ7C0n5RH3USKyXe0WWzjVV5geK+Awy4uo8J
sWKMENrB+12WLmwQmqqkBOCEmypFpJ1dva+p2+lB8rBEc9OkbqLajE7tmHOCLoaz
6TeGkLMvJE25iw7Ca65v2o/ZlIFutBVGXQws0vxttvNTZeoe7fCSYIWAXj0Va48i
4vPP3YL8CCKTvC0Hgmi4K5cPB3wqQlXx+P+cz0mU2VfaGqDbKKmzETJ8CjwwnEd1
Z6bOYziVV8LD0OB1CMX0UVzmRSL5TtXAWbV7Nae3ecGjEARMQ3DrLqUOGpsDnesL
MM6tjW+jA297Tr3NEGnJT7zVwqJn1TiHWkAb9gWZuc2MvH47esrWGQI9IY3bbuBh
uqaQQe7RV7gKyp+zxV9ZQLqwAOFmIhossgwhAdvDBY4ci+lwxDQMKlATjL/FVgSB
6xDwkFiK1LojsoLtKgGEjZ8OiguORC9Ajm27nXSJtdoDo6auDJs41hK09YVfSuak
FsBDspxf05sN7WKoWGU28bDV4KvrR/0+tXYOhNjYO0BCAvh7Y7FW4KHeabkvUC+r
rsXVHzRmgcUZjWpEt2kSNOCm6wkeL0/kdULra9sDHMLb+ybFVQIR4er+07QDXXAZ
eRU0a1kqP9zbKllrjv++1zaCrpO9V1kGjizAS1kFxKJ9My33gPcWpdgZXepVt10S
w0nRz+d1hNsULZLIgkFA1+Z2qALsy6qLFt8AXj76/WQl+cVEhNqUkSgWfGgvwWsP
ruoj3NkDuEo9j522u14u4XdLlj8gtix2iTWJdsnyZKhqm16B/FdCLOyqAYfnaufZ
ebnwSqubSCIKGkoFOdQhGjFrLvvKkYgNICS3EtLx25NkW+qPwFotAWv12QKkVWZu
B/K6nBEX4qgj4sQdi/pJilvkxX3QM8/fTaYeblHYGpc6qUKS9sR6aU0xMPVGcaJR
UKiDhL4UxIVUvlxOA+aO7FSldUgeg0rN+3ykT7lN8DvoFnEdz4talbCuwSxydqMz
jD0ijVyAff1DodAHmLeA9uXELDhRe90DcB/mCDVmoMKFLKNIa5YfCz5Stlc0vfph
eU/jHl4p8tg9eCLjsmWoIcnW9TaG76TiFhGjC0Wc0J6pwjEL/i8WsHtotG/bzhGQ
o9lq3VS2T4Qpvd3co5MGS9RkK5T58U7qgPUmtXWhOB6EnUnS5di7GVbhevMTUDYR
DkgwTNJbUaqBGbXsbzC7xYiZz441c5RL4XN2X7txorv9GJU25nUYWaslDGsq/U2U
f564B9sjOhRkw5bB3x/jqYgHjOw+xGx2D20Er14Waojg444iCm9bA8rAPP3Ol2T1
qKjFefXlgFes0Ff9CfwuSFHH14JR0tfoa01vYkR3n+OMR5XH9kRrf8d97Izp5IZB
kXroxzi/wJxLniJdz/peVwRgJrAqBH2L0sDZAEcJQBO5rJB+g5JxM7F9M9A/msfb
aC+pOBHqUAe7i6hLbJJlaj19n8xveUOok9UtlYrU8WpZbI8qoolRR3RZ6f/Mh8tC
P7B8KCEmYWV9UKFVyt9j+3Frk/qbHg0gbWN1l5fAoyJ01QlLzl/F4tKA4SrbRZX0
BD5IJT0IfHtZDAmQfIh/bB4tPEH+qzZRLxQjgB+8bBWhgS1Bci9e+HoUKRJv3K3w
VbsWmQwUzRlySeC3hXElaAJnBh/srervYYz20oZhuXiTYTu+MgbfJWX6FBx0n+vI
s24RxOzFK9A4ShP3u+5fr1W8+z2kZAslxOWQYK10rQFd6zXIZu6bz/Tl99BPXspi
tyU3bkdCN7g4KCVP+/80Gde9WjEVVhVd0YnHhtmzZL8EM2fRq/kTeD5ch5pot578
FR18I17qlZxXTLGtTtN04ofhB1K81Wzb0Bc1PSTiEyugzMrTEXi0nXSyQtesOVwW
yxyeofLUtQKF20HfHPDwb39d6zUWQpfbHZ2Gx8KyQfVfa/r3lKJn794tu7Gq59Lq
p5SsTxytjAbr9vwU6un1lITIe2YBpkLvPmYyAGTlfdueGeACYWGixlTu1uQ6e/FG
1K8Q8M/aKwuuN0vAsEOvdrRwQzOW2vYf+YJIuhxbMjMIuL/NsblpeoBPl0vJoK9V
37In4RjjvdlwoaUPzXjikccFxC2OdxR42GOJv5e0wfgJcYWbFGz0oH7ZlStYMmzy
yGiKRvhE2qKp7yDCKY+cf1POs+HQCYIyXonsG+1Curd5ZeLQBroNpzFvmKjMjEtX
Dy+ZchGo7aLN2gWa2LDLJ/XF9aJY71rO8QjTPqo+NyNMH/mF4zMXKDqv7i1TvZSQ
z5NLxBI4O0MP+KSQysY+B9UOmd7BRk20DqbJhs2zsiU6BeAMUNEOI3PLSeJptaCK
XuiUdawr6g9nXbh+9LsFSqae9aukeAniynErZmjsTfLLxmx5iVjReZaEFVUvgr+9
zCrCLAb1JfnQKb1S/1fNqURqzrnSsgY9o5VRl2iIiFFZIJzzUxA/3A9J6X+1QdKs
3o2kJMRrWIY30gbh2ikuFdO26br2t7dfzM41zQJaW2CFU1MZcUbTzullTcpkRJoI
ryuPtEm0hyqX6RaxXs4Z7Yi2UK5gHoP5MtDLcd0pgllGWIz4pClTgXFqyZVqtqLK
fn3wlpo55El+GWlQsrNfmJAcmZ6CJIQYb92hjF+vMMDwQqK2hhUoSX0U1mWN6AMj
WxFzWHMBiyAhgsqnSTplfCf6FMs6mECUguikT4OMxWLY9PNGg8zrMyJ2yB9T0/Sb
UWtVZ+RIpDFk9ict3vKnpa7rp7RYHRosXJcWANaIF0t1XkEYSbQTLK/70SRjMVfu
KTvPopdjJg5Nh3kXmr2cu6wVXrducustE8pe7ylp7indnut8KeRqQ2W5y6cC9Afa
deOjFSadInE5QKYxHqfstLaI7rviiREClmeCT/afUBqtst1ToOLquUm+eUkkLvip
eJBJvy72oyDRCbX8t6G6isE8Oj+j7MvpQaeeDg2j7+8KedK1Sl56JSkTVZWX/0Ep
uRJXeIaa5mMNdg4AR4Ej7hVrdGqOtAv3EKTPWiOB6quLi5dVk98W3ifGEowW5scA
T1l/udUimN49uouXhB3xW06sGFCcf19Qgi87CRDACXcAx0YGX9uyHvmYeY9vwIMS
LmAOyafWN6QydjgAQwa+o0bVzIDiRhfYVUIQjWQOOMkf3gUySfML//WI5D8bv1Aa
Mbp5O2amSaQOdP54g9ZXJJvGREpnDgM9JxgqAGhPqOPN1x1R4zlIE95N1lPmh9nw
f/XujHNAkcgOdLCVw0W0iBYTiF2YXINxvxorKCBmD7z+nk9U4J2ST6pirURBoM3b
l89Y2G42KvZh6uyR/uZ2vZ0dTlXcypcBB2q1lp4UlAHjvQJaPL6eyLrU96LFI1Sc
PtD/qKYboZugWsIVj+yI+KTmmkan/c/yT9nIpjPBJgiRctB46mgCLzaRVCX+7OzQ
EtGXd5I4AcY2TO2Kjls+q9li71iReiPYrDjACHxTdFBmE3rlwuGfW/DfnSeH4Ydk
m1XcqUWS/DM7HSmY3fCLiijcuJR7mrkodt0ribq4SxwcIVZkloqJiWT6xU/oh0S9
xbWBXxiu7TVXms971QY2/Q5yrji/egPq96nnH/oy7Rixb2ECEIL0pGqpKOKOUU6x
VRkWTUpaDEykTGoW3UnakzWWHS6u5NaLtClM1ixbLAV0mk55kU3Kpg8+HbOl4jyU
rJ67N315Nv5nJDjNbNTgpqdmu4CXl2Bg0nAwJYlX3ncBQ968q5ukZjfRUuF7xmMw
79H1UAO9a8h18XtJpkCSwwsb1Gs7XWJzFPdz3QTJE4QGiDO4pR3jG5kITqbGll3J
qv1uzhcdlL2C9qQDBn6NNqcvT2glK3WJJ7o5N76OEqxWLMgF52zOejNGr6Y44vTg
Zq4hnXDhOsT3BQBWbrahzpwI7uQIcM6nKywNH1nc4hnrJEl1mOXJ3qMAUVjUh8Vr
946j8/j57lRHO9BHyf19SqTps5T9LTZhg4v5WT4CO3BQ7imIcF/l0Z5gKpfLPBkh
5qpKEsYvxWwC+eNinO36DUHx9SfCKcBy15dVhMzEKIk8BIeT/jylqyBdfAqR6D/H
MUSDCg15QJggfT390Ku9v010MkmpFLywgxGK7c2cF5Rtcnc+bGfQD0fnA8hH0Pir
5ZS0y0dDihOCNKiYN7sfwaIw958BnfsTsOqnpwSPCK4IC+QjxvkcXnxip+zQEErZ
33rAOFXqtXBkE5PDcFPBnhk/rYwd2KpdxXzj3ZBF1EvyUyYgwjAT6E8rM+lrvG3Y
KtH0OSY1V9JiK/j17qZjwyqLCkCxDfVlgoT5cfg5GYPlmvQOjORY1KP5MV1gIxFq
x1RcZsCMDgIcqhgMPHLXZc/MAPonKx00DDiUTdP7tU/H/CxDCuPJvbXIbK5ShVz4
lLC6UAFl+myQOoOKCDzFLHKKws2ETtoV7YFw1tBtouvHS8n6igB2Hv8oYsLftfMV
uQml5VqqY6gEqsSWjAZNUmg9AabZNjRTQFRjk2CYSt0/UX14qSP7sKrqzENBKIUb
GgkXKpwt6waFIx018o8DTE/95ge1a6OwYZvRVzetOayj/VZTwtO8D+x33zcLFKVC
apHj9gI4SIgMC0nSqyWtXyqGt3oJmIb2Aq3fZ6fzEQ3DySbkrzZJvTOLG/yCUCLU
ujQUbf3g/JVpGS0Pck/1An8skMEbHkqRyv5xFKfSyIJzLvZw95W5DhLGFy4Xaux5
f3GUVEp76t7MLdd2NPhBUujowpBqGCYdHqhNBr0l33FmC4vc+aTWjFvcYFmOU5Uk
4/WWO64rYmaTW3W2ZrHqTOwc9Kpf4cbPrFAhTX7z/pY2VxXDcE++SDfYkpPnCebM
34c+Gf0WmBStNgo3HqBV08HSZUsWmsXxMXN8R0O43sjKS3hDYiSebB9gzZuDocKD
wcJ0a9ERcqMnF1qArMOuWste5Ih+Aow0mhXogyhWwu8oZQEKjYa5qxHI3fReY9dU
mdps1p2Esnq+yft1GDv1gWbTG/gvGg1KUBlrTMsy1rLLQHSPqy+1RxSdpFW3UFt6
2aMRRAbpBqV+gg90PCdMlkI20Vur1bTjmsriDBt4ovVYAbXKuEVhlUgMbsxT3qzU
unYxwNQGsTPtmU6G2PPOrAXs4oMSzzFtibxab+461gTXh0BnuHuvC3vPKtRl2ThW
X3oJjS2UFpKmZc0Vh/19YbCiN8Ycgn5PeQPU9OIIn1zP1QodC34BJV3/dd0vXYnS
LHST4E90OrNBsJtJG5oTAalFFCj/j+qf/A5V3ePblz+xudUpvUwLbubg21A/hOCA
R09VIK8ylj0CHl6BauVCoH+tIT5OOyJxElqBnpL05R3X/MSQUIh2cK6kt4RKnZ0I
MYIjz59W4VMDjQgBJoXQf7U7jsASlCi2ErZh1Pr52/wtawl3JnSfYYDaSa2GbtdM
4PKmUah9UpjSKdd/k0hyykXjkCNlbHSSxECBDU7tk0WnrWp++DLwoV+nkma2wIeU
rtFsiDnn4Mq8jF5yxQaecC7AhgZYJyxa9mGJQ6TAExTu2LjonQgEhal3hxs3gF5v
uEUiRvL/jsc6ovw7v86FjbhFqWn95kZt/wUypWMoBkerZniRcKgqb1VRixyo58yX
9AJqgxwub/j/rItd0A3yQhB8CMITuiApwuMyvxtgxAKbT2+PKbthciLDNGJtmFnG
omPOz3lo+KJdPZdO90M+T2IHH2IyJXd1Acwt3pu+kViwuLtMpMb5wKduJMHVrp+2
Na+Rg6BIVLpR2RJFqltLSjTvLmLc4xplXutBvj5OYdfLEtL91NJu+sXO3yIpcafB
lGXDtrXWpzLKmGpCZPNi5qLC8AmQ/L9pOWE7UkxNYEgqOKCBtzjdyymcgAOEkGP+
jo0hRTAExzixCQZbwLxQf/SRXoPspYgAEoUVhhSF1E6omGpcajMLWJhzmogr20lu
sf5a6dZjGBGCGcMEvVkYNhAylV40xgg0XeOFdEfUhIE2HbhKLcUAjcbZooZtdK8p
PsLr0PQsdZtFUDVUm2F7bDBPhAYq6yRXuxUEJs+KYd15k7nE7heeulMOTiRfho6u
56obRA8tTK9uG/iWGMv5EMMxRnJCX4GsBReXx2Luegk9nsDAjgiyCElGibXPWxpE
YTCirdJ7ovoRWVYrzvMGb7VvsEbeG8W+CgLYbagblRttBupFiRjHFT6HAsygEpST
AAb9J7liP87J3vP+znkQG+EDuMtjgHc+MG5/gRccL6M5VpAfBrEjc3H5LxptoNM8
1bdSltYQBXXAuJrRJo2rvwHE+G71P2ocjB6OVqDfAk+/GFHWxh54OTz2jykTAP9k
BGejCPmjhzrlmHAIhDHw5322eplnHpUYYje1Ws/uf7t9LJHrAP+Atckd0II8M6ru
to9PY4oHHHPbe1vcUsjMPxOazigXjby7RXudUuF1WQ1hZNMuJWsxp1DjZLKA6tF7
KUweFM/TXhVan4JMA/gbxsTfyzhbGbUpvRm/q5gyaNfEW7LNB4F2vTsDU6pnpRvH
kTRYFtHu4jMIszEuL76d1f7BshrO5Uyg6gOv70qS70wT81zxL2gI7zM/1iCQU1xt
HyxMsRVMWu6wxSC1duMwv/YkJB5L4n1GEP9zl/TsczZ6Oq81FIUEws0ZC+MjI6+g
+ZwKvTX4QTerKLxifzMGXDfqL9I8JBfiFj1tJEV1NEGRYoj5SaFXAwowlIjwsOeI
4DKz0ULPwyAfNgEbRN+++ceqx6U7xALUxGDyytp6QD0bEJNAdxo2HEpM/onGYdnN
Ow6EcCZb1jX0PZFScNpzZNGx2v9bFNhmWy32hneGbzEbIctOiTbi3hrYVBYC7ltl
NEbTDSJQ1WRiIoXhQr7PL+1XwJd42lZM7d2tcLD5u1iH0YW3YgxLZhOMpVmSH8sS
ylS1mtHRTdOpdeEskc6UOxMt9CF2ne4DHqYBWKGOVXZnb5eJX3e5J2XTvLTgYxGC
9QXMs0gPTEwa6/6ODsuVTRJg6nIitmORgSkVPzMdORAYFkk6rnH2HgoY+SAAQ41g
SNFi035gsnYn0lGYuWhR0n8Y5xx4L2q+y7eoqv9kqejAv0tWkgjhNuTVQlz+UtG4
eUdoi7ixfFadrJh92gdf9mF+EJbmOfB4lEfXkh12iz/TgAXOUmWqjXbAaoioVFc/
v6aahkn2nCMyOkH06/p0l+4NIgsgkNl3X9FF7J2tGQv6IHZ4tMKo/WR0yD8k/SVk
SesMF43N96/X2IAs5ZhzxguKrc0BPSP72gAogGO3wqoTyF14Ooyofb8IBAHgySev
zqsxwRpwwbGuRCtun4t+x8mOlt7QocqvUEgv9iVPuF3JxtNkJTzfjcC6U7kRTx5w
KGX9+6dS/MaB8j6RHlYqj0+rvX8r+wGIaahpYLJz5JM+SnP9xz4BihHK0e7CpjEu
0UcQb/3FPTu/LqDYtMSRcBOVUhtVpS3eVP8IY5A+tkyms0Cyp6LYOuihiCh4t6+i
9Ipy6/ytOF9f6jUJf7ciusa7mDeYTOvcGKJ4qRpW2tOH+vZc3SBbzf9Bg+VCfurK
nn1jU54VUZko0W/rdNRfwCCumM5z9KGjijS7a/4EQKLwFJPyX6bJBcnyjht8uXst
gpoEOQuuh+rvnXIr97Q/OxR+ef1FpRv5iy/ttEmay6QDsJQ32XW1FYiTowvX2CMJ
xgyeByBE+MsoCpQOCX8DfSnKCdFpSAG9c4dP7t2WhqzAY3lnMUE2OaMvBvhqWNN7
R/sFMi9WSEiqzsV1KEwwFU0u1ZoGKDaPSA/Pc+Vn7CLFpCnuH6gsOiSbcKwAA6/U
b2WbTGAlgn5qpo7MOCie89HPzE3ZBmCyQCaM7fEYHCVOEtj7hX79gJFLgwvz2HCU
6Ta5+a9yPVNQT4GqN4jFE5FL7zjsi8/YcBxzgXbU9cGpTzpbpCMyh1Rzh9k5R2Qc
dtbuI0L3M2ve2NCbPlqa15XCF2FSzYCM2XK+FuzZzXmSuMMmic5GUUlbnVTJdGT8
ay7JejZlYjgkmNz1gdMhU1vHyrTZWAV4Tplb2xvxSQTAKCQDiScQs9EBz8fvCPwo
vJErS++215T0nXUGoC3MlpmclhZApDImV7NitIhawdVi/RSXszxJkpSoiZBYEUnV
z0yDaNDDbhzmlejnA5/2lVDubYMhhId4I1KfObzywp+1vteg/fbkZhgwP7VyWpww
pqn1pN4FpAJNyaksq+WnFZ5h9VzLnls5HuXdwXWH4ThcAk3UP2eC7AjMsFHD7zOM
yKYSwa3v90+qrXXgci/e/V2dXIZB+Hc5HSxJKcV7e+HZf+uEuzxWPZirG21aVDMB
gOdm+MprX7GeYu5R9fMzXGTutolY4aeglYWbhSXcOuh4jOUV9X9UHfRIxraNoyFO
H029Y8ybIfZ9KjuxY93c7YEeeiDt3yEAdWbQXOZTQooAHiWEi9t+aVuC1KWeYNDI
aMjpzf2Ob+f2sOj/IiPEz/btCq+NakvVS1HfLFyvaiDqE0TkVCAd/1mhETYOaoJQ
H1AAvwPKhVpMJVBS5NUTJkxEfPXIcJ5ouRDXsn2vUpXpBr1ToNcTuTWNR8q//mbS
ds3OU33a5/kqGV1VivpAEdJphcWp3mRa7El1S+gEkzGFi6RNdX0Az+NAG79nLDQl
+Yj7r8rRcgJFgKUdvP+DesHJ7PGHYtvGcovrFIqkgUNb4FefXbGzsCzQyCvao2iK
Z/W/08aim78B4l4EXWzWfOcnlZjiloJT3ce2ZHwYjpI2zkeso/t04jjWEV3KUcwk
tGVL0C2lh+29vwFNKVTs+oB2iFPfheCjuZflZaC/LRbHXVNdaVn/DvXOrroYBjwP
yzBNVQskdr5l3UahvDC+wxkqC3oGKcyOG5PPde5Kxepecb4K5r/1gBgrtrVTKUNJ
Fp9mcR3S17eqtJpJfsplSli58kLMf6ehRJX47FaCyEx4atYdfeCjQ/Qyu7NV5W24
BBx8/z+KGKBR265gbZgJjg6dK6KcaofE89Cn6a5iDnw6m0jBSSqPfo8GkgdGt1FX
yscxgVyh1BLu+dvGbv/XEJ0ZcgZA8uYOiCa/uyMu4cWfPgSP7Tr/6gUZZZORFzHf
iJLlYkNxIVUj9VhWle0aLh/luJM4jZNbakZGmhHZvzBqZbzNDwX5+JuvDwTn49CV
w9OGdTbu5sjbxJppvBtF6d/1ea2WuZK1kKR9v1hTncJVtcQMpP2Vx8DbNT4oolq8
WeO6e6Eppr8njGCg5ZHYD+kFm7TpU69XObjp7ozgyDUai83W7y9kixcGYwCPf+tm
saifTZmZcJCr51XqUOe+qF4ZKSCaKg570ZscmvUvvcb5Lp7jK4i0QGMuLvXuncmA
zI/vRLz+EsW21sA3U2Wi3Ue3WHBxjfeRCNS53f/mY1JB3plhst8Gh1ZpScHAAoPO
CS+vKbx8IVGZt1sy9gx0ca3+graGdXBsekt1Jit/MeaaA5leejKRYBUstnUAJrhA
cX6OMc3CLY1OWZlQvtvw7rqO54sNJlmSMFaD534ayKM8xqNdt0l47S40MuSLVZMm
heqHXfh6H0jbOeoPQPlzmLsTZ0/GwseyC33o8NcqgHKEU/hNRSLGFJUdCXma8Xzk
AzMKOackGms9zNge2I+LZAzh22bG/tgw/A5ofqBrNljI61y8bzjgI/pNcfwFn6sW
vnsmUgUav9+y4dnzBBTVNd9suBJgvgkWBLyX3GwzvxZ/C3jRbCJl5Rqx+fyHVBIj
1EQP4F8aKskLkBggkiwnHRscpCdVVVcoEezHewrgXM4kRXuU0XCsaMRxloZlyujj
cRMokjTFNbiv5qiEJWn05EMk3PawejtNgpwg3Wo6DsUMc5hFh9DbBok8D3WSiwWL
iXQ3MCpBqq2fowF5F5W5/YGuJ6pdvg5vh3vH5D73T3yLCvsIIdB65JDxYWWlRB7d
MPglBoaLFiQeOQqNWHMsGamMXmMWAdo1TvjL9yvqp9ddGQQkV+9f9PwSNEy6w6D6
UgCQKVaZIV6Q0c2F3WKs9E+BCNACd5IkcTm04wwpSEJ8tX8fCBfbQFVwv2tRWIGF
aOp/A0L140n5jwV28mrrh7yrr4arP+c3xczdvUJDMJx3L2PRyAP7GFvgiaUPS8P0
tgqigWhuuXcueY8eUJRSmOfg1PyAFW94ItwUAP/tOupjJ/nfhsSC6oSf8oyUuB7U
5CDIyrHurhiKBwfV/2iTGw4mRKKBWxZU7TesByIVIFF32h5tWJPaQL0yiKtum1u2
D5fsqOB2ASpVh6FsQ6tOVdQIIpXIAR6yneXIuen8RrBY6kp5+FYWYf8pm7d1ki/H
XvsKd08eKWSBjz4bHnKSLwXgGLuL8UAUjTj2NXKSize4WJEDCeYWhVyhl6yzkAwR
hBLY/KZasesTEpuN4r2LnASh9EmhCqm/G6cfoyLriQ4tTGVap2LN1/2iLhuhemk+
vuzmTVblr4PUXOe9P0+mTNa3q/GWALOKdbADe5j+N7Ej2eBBX/dPZWdeybXCmPd6
tThnWBTOFzcEsBMU9uYG2qunWS2OZhHQlYqd0NXtkBRpI5eseF6X+3Y7MfHMbyCi
4YrFJhLOK6PSCLKxg8+vjm2BPcUzU/qMHG7OZ6iDAVKIrFiMZQUPi/zkw699rJHU
ls7scMT4WijCDHaXRd0hdyqbZ4bqEad/1mhqnhjHGG8ITqL8RDXqNcTRn8Naei+Z
Duz8QVaOGTAmQQUp2sK4sc8121I63hJBzJKH4d35Pl3h1BpEd2u5TEvl7VttwWHS
2626gbhqQ5p1aI0xsUI19HK1QcE7MFYW/tCei8hqNsBDxXsQsAr5qZyJQh5eaBQw
UjZ0anzqGVdIhKq2HYTrI69Gjw2AK9WSy+qXSvH0L8mfTpeKMcKZi7YwCIcPny9K
l+QO1WWIYUNA+yx5vgW3O2U4afvHRRX0rqrGtWmOfPL4ir7TITob0UObSOM0/8Vw
Ugag7UL3zx7mBnbaZWby6D6eRH/1m/E63wKZP8u5u3qE2hX3du7On5nljyz6XcaL
ezZX8Mhg51+E8TMSCSPdx5w3BFI3EEv14iRN3CZ0yYerdkP29+VO17mGJfj+gVic
/5y/kcz8nMbkb73BJP+x29Bcyc/Aagt9xfR72cP1WtObhuy6GnJc9MxosGB70Zdx
HUBo6zBiaBHM2I2kYTBjhA8mLnWom88/zDDPEwheejFpz4HaqZWgcTH7f3taLPdE
XNBAhekaAa1N9Y6OF5YgH58P5aNhi2BAbZOw7H8I1Y+ROCQN9AFAJFNbAXM5h9fs
+ez42bWFt8IJj+pdpnfg1h7eX7gT3gsR5hGq0QID0sLd4v1vLRCt23M0+kRZK7k8
wGtXqmzMy9XPl38ehgSOi5n3bbxp320bhyZheePEB9P3iarNkTqQnkQ/Y47COCsj
IBD1j+u8gn96ePm4mzau17qLQc3SsCHynPYrS3bUrvX+xt4xmS/XIdcEH9PFs4zE
Jvd+rf/fWYSMQWcdc28kTnkql6KegdQquRlygWxA3tkuvMghyZTx0ipDXgAOAL69
fNhXNtuquSajioo8ZMN10Q==
`protect END_PROTECTED
