`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u++C0BAARnZYp0wki6fTd2Yop9vWM+JAYV+hGS61b2kmyTG1XHZirPA1hbsztKuO
me3BR5bki8Wa1RliKDKW7ZuKUFl/uNPWtwCwmoRYemXFd0GBMLaQAkm0GHGDpQZK
mFd+j0sB+wMhVKUGQdOWD/dEQE4BYtSGuepyCbE9mpqmSlLccD5R0XGcwEkVqQBT
4VUTCRcBPe5J6AwgTcofcrKC7/XbW+DT+vm6JW5bcWr8WaXSCHfCBre0Q9aVsPQj
uIwjoPmoY42KlGXJLVrcdPl2EdU9tIuXzXXdiO0rABzCGM7JpKWc4nU73OGB9R4Q
XVWopMM23E/r0ExvK55T7hpHk8zPBHQEU06h18ctxE9jCKop1nDgVSMF+qfclDfO
Zm0llRhbKFLRnys+Y35PAgq50WQ2/iot+46wgHksnSnCEk1L8JlKZa4+a4jIOal0
RuDYWtOqu4s+sKLoN+FIsqBNFMCFrkbk3BpMscnQincb3XkpOM8+G90NwHI9RKTg
EPdRri3NyL4NdZgd3SNJhLEp6rPTM5kch1VWo9qyJTi55iKjFGwvvfM70ekX6Ow4
vkKK5y5s5lC4qWn3MGq0MZG0c4I4ba+0Qya+dT6bnHVT6OFGH06mdD0iKw7B932k
1yllzO0hyKFgbd3pQds3yKLIqbTX1p/pTx0x38b1NDo+vz0MiPUX5EDIS85XnSmu
UxDziAlqKmr9W4M3Dz0S/fvRKNDmc7clcESDDtfbeoyNiJCZWfGnCD1g0YRbK2wR
vJU0FbDXSZTflJ2j+1ghUDtlRUXoY1L0OnG0ZFkCT+K8QDm0lElc4J/HwnLUxKWD
Gnaq5R7vCyStK3g38Q6YxfqYsMr1p/VgP9wuJiEJ93uBv5piKIhqUQ/4qciwM/Pc
5oDHUekCsfjQs8OU6dicmfTKLfBPiYrKxh9CXcqV7h0p+Eg8asnLiFAibyJJWdnL
iLjrGekX8p5ulehSP+RDSGnKx4vA99HSFU1sczj0NAi4wsVzRLqozVAZN+ZGbWpM
n87DlV+hTfru2TlQKCSMqvyrJ6KHGMnPfvLt8VKZr5lvN3x+NQTvsHXfV1eaLBQO
f02s9ezJHXpk8TA3LtQiOEzNsp21g1fYvbpw9Qkz7sSyoORAegV88sSaalT85oPk
Z5N4ZNutsICOlxwx++Yz76ULFdOdRL8TODWWuc+BOMG0g0QKwi266aan1AlVdpCd
Zlz3K33sCCSMat81h6Hp9eNidxFOp/a3tJ369XQscuanh7q/5AO1GHOLJr8dgXFI
15qAUzUYDQ1onxhoDwRtbjoObwu5JT4gQH2wxRKuOMU49Molwcb0LcwVCVSDuKm7
`protect END_PROTECTED
