`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MUVXyuEr4vg40RVBvNZX3eerWqrLJcRuxHzh9KdVu5VdPa3hen1ErAw+g5mFwtxd
/aoHtnW79qWe6bGXW4u6qZUzqzcYxHXD3tR8SwP6DO/HW26uKBB90fwpka3Qryvz
iW9OdcGcLFLk5UI8aRcWvC3M44ZBa5fiwbYBikdi5U5m3YMQ8TDJyTQrOotWk4m2
0Fl+BuyMyZto2qa3dQ3Izt6R0hwrzYbhCdAWNZ3TWrf2GSW+jyWJerxrhN2dAQ6j
+ui1SCjXxJvaQI3vppNCPmTD4+U2E2jOv/5iPO0UXld0NHUb+bKX8zI7ld3/8HDp
CftnN74Z4NHaBl6jL3BVfFBwoY/GyTvaBBPLiF8PcIr6XSHB/XrEjV/UDCt1xdOy
LWi8+xAzXp4zTd/vh2R+2F5kvx8vr7lPBh/DI+XqbFHEqEPCHeQBv0lxd/dTF93K
Jb+IpyOOsOHo22SHmPLi4glHJyU+pYKjP1qquVTaAlHSQWPa476/Gb/QiYV0Tp18
3nxHqEgz4vT8eGOfZkjPTDDlUxrFBPDxDFZxHtSIoxHxi5lfe6Mr9kD+wmZ+UF/J
SYoKwDq2SR5eVCWGXdLUhOEpdhbf6KFver+iwqLTWWkBPQ1fTUT/aeuv/hGLnHfu
WxjF3cwxfUHBgT7OnQIquT6KeyLZBWAKDeWvco5hc0AMBP8O2QIcgTPIdkuQxXje
`protect END_PROTECTED
