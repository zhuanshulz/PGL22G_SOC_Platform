`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xk0gAxOKfMhRhXQqx1GiDPItG5x7fFpYN2OFleOE4Ux2EbccbkeGlHJMhRWyjfBe
5EvMNJUkgmHcEWmk2tNwe5wK8XiLYlmj07Ywb2SjoE283EzJ6v5dZoJeok8N9ffj
Oy/ZHm12hOmdaGMuRlVFyc8t30IjJG0TX2vP7IPnB0460ATKvzi+UXit/dLyApNn
Gsxm2lmV59LYcNvXChMzomd7M5nkHbvT256jlgegqYe7t2Wo1ODPvw8qcOkhn/q4
g+HkVeu7pKtMyQqNmISBns3UJTdjvoeJOnxkjjVu2LF7KmSWhW300L/7AZ0yzcjI
n5TkowbB6sgcNHaOLgo+X66OE5J1o0q2fz7wYnWZLPXekBxt45V+3d0QOjrvs3p4
1T6kkAlE2BfxzuMvDRVucy9k0OpLVrrZygHHTh4KspqwvrOLaLO1xZ8oJhhZ7Bda
QgmGKZyGdSvftdL9Jl/JQVv9qV3X1QmeJPNRxnXk2xbx8k8lfsH02+xLaLLKJ8ct
OhUNf0mQsXQ98Po/IWO1mQnAm4UpH2ZmPQ76a01Hx3n6aVYLvUbJxhtkPS9dVipm
/44qZinUCZDiK8h/JsnP7ZPZvoKIe6fQ2/1r6+N/Rotgn3Q288+sjnATgDFgALU2
aj0lJ2ACqORMomF7Irk6p1ELTrnhpb5lNZkmwUdGeCKTr2TUR+5ISOztYFHahGcp
kPxijDae0opqCLiQURv6uAswaYfBzKlNKP12RfdtncCLcoAB5RRNTfpUhQN3oKEL
M+SVLYmRwuHK6XkDoHXlCObHd7Fn9r9MPo6Su0VDHI99dDRjqEc/Lbkn4H/cCVPh
PDPWP7oux+KDxAkEJG/3gCO7LWw3Qf+RTKZJ+RK8ouIk+fBPM9IP57nAoYQ2VGVs
mTrCPHhuRdD6g3Kdm3N+806F9CszmbEpLERws8zfwCuBnPlkli0QSMUddciTL3IC
xICB95V7N19rZEagBZ9bBg3xafjSPL9nLcdtq+M5NFQ=
`protect END_PROTECTED
