`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9KgnHucetg3OfPRg49ZjBpV8BEZ1hSIpRUXQDwahNAyR8NPoxw05WreHAby1oPgs
bHoovP75RX5xk8z+cXU8y99vgPtoxBmxaQCvS9uYaGTXgMQB8KRo1uU01nOIHnyR
L+o5GrGhMD8xy+e7+f6qr1c81xqPxF3j2bEJuiYMKrl4/CNqwO0mPVYrTNiDkWph
9Y8h2wCgtkzsO/JbJiYd96rMqjKYC80CBWNWgpkhmnphr0RDCNEGJUJNtMC42tN3
M/JiIgDZab2jdu6YcJAnXn/Dj6c3fXFysSMhLfV7ofCVuSanj83As+ueWADqbHF3
+Edq2im2wAPss9KtGk6DtNbVnV4ZVc36oVvKX4lF1mdGRDO/sdQm9LR/niaHP9uw
cfcDHDotfncxJPzOGbEzpPaF7KsvpDkgo7rDZNM7puSx9LGZ754iNtzFPX7yD1iv
2TLWD2C0ugB4jG8JLVGuKOg2V7AzbJLrr2sR5K3rAKQttdmutHHgHCOeC4sGJYwG
m8Pt3yVeAgIxdiP7mOpw+ic7ETzxzvEvCElRmp98Xd8=
`protect END_PROTECTED
