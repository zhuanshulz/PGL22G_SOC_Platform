`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mm8u2z+33h1w/zxzug2jE1h/UphmjLWh01E+W/9O8d0ziKr6k37A64MRrL+x6h1q
yrkgrNv3CR8Jd8ZjdfLtcWTtKGrE076yFDYd6sfMDoR+BX+nOYet7DGTWvCH+UdO
nGMAnXq7CE6Gd17UhRtoN8+mGeosQ8XpVs39xGpkdBc6qwb/MOTaBB1z6sKvHdIF
T0Ig508rkrn+y1wUPxA0O+1kFfClVpT4SISffeuKmOadG25iCovaBYlAf/S1tzpO
ZQMII1aDRK/g9BcsUnrCQjRpwbTzPbNLCekzkJ7E/z29XmVD7NIZ5dSUrJhfQMSu
3BXLgVXTQRFEvFn1rrVmuxdlojnnUmfqeOshIhD1K0atWaD4GDKxBlV1CAm0saxO
XzDxyl8cOqQI7OxvCfDSEmph722/qHPK8Q29ECgYDNI9IgGfp9bACXhLVSqUbWeC
lmNQ3d18zd2jivIMeRoujLsaz8N0qO9MedPj43yXSfVOL2xGYMG4qPvcCacXmCcz
1mTxCDXuwQrt5H63l2s1MqhqSKFCfFqSSbTkM6AGLC4Rma2ErOU37s/091dpzDzJ
fyr56mKH8nkz/t9zBttg2M1s9yevM/u6LDf/wejGPJplQh5X+cDKSdI+B3jVa9fy
g/SdWyK8/y4gR9CGxu8raiQc7Xx/18YVJDlO59gfZQCfsUaECtu5lsJF/ptZiA8E
USR1iMzntFvj1E07TQEB3XNbXrc025QekmDhdKGvuDI2cJbFFs68yGrToCH6/fsT
SIDWbjRsY5ll4aIiojQce+xcLr2PoIO7kFDqckoWmJ6G010VxA/gx/84nb3Zka99
ZY2dyZ6r7YwU79RW1aXrlkRCQPV7wVrMUlOJJ/gbwi9123SU2vq0o1jhRqUp46RZ
ekbIaHAADtlEL0L0zpvuSUHINZUk02zg2bJj+HV3TqDyJYrZzl78tBIITU6Q+NRA
V4yBa1VDlQnYQcvlUPtVNfQYaxetyF8orS/PDfdwPARrKFWQnCIHXMBeIwPboPmZ
DbJ5sVbtF5EYZatuVBs/pmOd3xOFDxOKZISAX/ARBMILrIN08ffVZub7qcvbNyiZ
mRpw9MX5xPXvZ3K0GejfgPR7al5+XGtx2rLTEZdXZkUyRqokL3HxXncTuZTJRpe2
9GDqezbesIMKwZWnocIEvTFkjm4PHBHt3qE9HjgaSafP60qzoi69uG5SNHI7Ja76
Ora4+AwEQqf1iqW7LjO8HvAZH1wGTvHqVh/yjGslYErlfaNRRU7+ZFFV7bYuBmrt
z2ycCBrCpXhSctvPcozoD6SBMesT9vx0o+x0snX6SdC6b3y0ggXIT7DWYOFaUIe6
VvFL8AMnb1ghbDPs2KwjtAETgArHJxk65ekyoW/rB64VT6RxR2wAhXqqP6g65b9q
bydgh+N6xRSosMIoTZp+92zw2Wna2webzsf5IgbG3kKzPhgPd+sv3UktqMidpSxS
pEyehTfqQrw0NLau48aZDP5IEtuGTBUOO1haO16rtHw8vOy6YiTM/d/GPzQ32G27
uhQabyVKd2samLr81V5L6JHN2fMNqaGHECj37A6tfAYztY9cNvhrM9U1y+r4Ak8n
Pbi555Z4ESa9VRYSzSdOIDKK7K8sddkqhV926PTHR6XWpwEudY54oY9QErBakHcy
opyunTaoYoScDvcC3E1JpZXO2eUivigIwY+pEfoP6JpH827u0Aa1njWehdhBG6k9
n91X02eL+OH44TT2WS1wiXfgXeT+xLxQV6jCumEtgWBNv0c+pYArCqS4ONBP5aUQ
OEdb7d6nKxpgEDyex3z0gdFi7ohxoOp2gAZM7fxviFNUn3RCfQQiXDC1WUV8Y439
/LSnAYnbUL3cYFat3BwV26Ws6/5PQprzLk5pSYHh8TeFy9+57V80v/+wuL7NImVl
zwyUiLJB5gW8ZjhI8zgvW2ao9tjgoZ40ue0j6iF+GMdz1JipJwiCfo5ljFw3OLZ1
ZN3mPvLXdsld991wrlWQ3mPb/GsjKHae3Cj6JmCTeMNYZQz/Ys/vXK3bNAQd9Qfb
zFKJkQMom1N4lF8co9PpoGyIU9nQyIJckq/KVIOW2lF+1kgIwK3Rmoi+sGEQsxij
uKpO79UnA4J8/Tj8kUYN6eTD4RPS1WeakuUZx/mDabmwr8Nn/JQaQKl/pmOCDD5Z
cZjKE8PK2rNuRuYis/yZFQ4fmaWG5K+p+NIaFITcAKqUAs06XVbIlCXxiArwj0XA
KPV4/G3UJ8/RPQt6wbjZ2nRhwSgfI08HvzL7NnMAtVY3zLIwvIgruOnyRXTJE+H5
gSPgl24wKkjnA1eHcAIm81/KTxkj2EnLKesYDLXWOrkwSVgvoDgrpsbn/c7cx/Fj
iN3MGH1+VCi29jXZ54IR3JNS7W3Hkk4NVkAWGqyllIQssXJvMn2FdCH+KS2QZwD+
ERWSbANFpMBm3b8T4IPBpcPo4HJXn8zINjjowz+tb0So8b0uyB8DHnjuahVV5GqH
pwjCfXULa+xcaRd099WDnizXbpavPrtUD40H/w9ojIkODrUz6FTY431GvKEOj5M1
6WAS/6CmthkZl/Vf9ndaAgMm0DBGGzAt2L4M49STTlOxQrHTktx1vW+kdYhRH+1I
KSJc/RZE1tEkkfN3y0UWEVRCZqvbrHSRkLBH2y/H1lnwNVhCHDNuSfbg7uIp/ESh
knHNzjJXLTlWki3KsKhfftQzjqvGmx38i01Bq1KJk3714dO4rQeWNCcK/gzSz10b
nSEmTrDHFoAWgtd90IhrynWqlavWcJl90SRbHSsQikBUIOnlpYzx4QRqFbpk3NvK
W/j7hiagPx7uoLtlbrUhBU2TLeiOEtFtPjJNq0V/8aKdStJ1RQbZflNSNme7vpOV
W4m3edS6MgV3ROtiOoywF4ZT/3kZPIdVj7yWFKDPt8NIaaAGldfkbm3q/kPXjLnX
/PepIPTUUiCaOSTEbuAQYvAObAE/Cob3TPVNTgtpORHW0tmtigNDFulQRKVzVNUl
7y/Q8O5kZEYScL2Rw1Lomw==
`protect END_PROTECTED
