`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eJWfZSavugWAEamiMI6jzP7uv84wiMkt2GPRmVIv4txuvbIPAKKpLzCwl7dvyWLU
sUKMJde46lHy512ZhMQz3aWPXFMKbhAHssULcPdbjuKfw4g66jz5DlF1D+BdG2Rc
2wmEKwLDjEtcBrezDaBJzKxrO1d5Otoh998+pwa3lDg7BiQ7z+zXSktMOFnvIP6U
JVvKs48y2FxVnAcncdN1ywWg9a196lQC7HckGSYriSt29BS7cDEXD20z77B3lwBz
EZHWqgTv8rl4+DN/ZZRHTo5+YdzLwtEoPby3Qr31jXwrk0RzTXSrRq2pgxu423QI
kRs1O1bEY7YlNWTWB0Xc1Mb9imQgawxwdi8pTH2Z2AdxsdxYKGz+RZHnOhSc8PyN
rOfRSWW7wwIfaMCB5UjtXOZ8OKQ8M04u0LhWg4FtxrnoFUyvnH2EqvxfBQ7vnwN6
hvpBlbDmSjpcjKMUzrJL+9A4ab4m7IK5NQ23JCGwGQjsBD1K1OqqtLorT+ApJdfX
7NxDkqGe7yFcgxfSRfNmkJTvMVvgxC9BNN8SprIV47l3VdZpScD+Z8wDoQGhrRD4
fDErT+EtG/XksoFUMNU7nfTf5PIDQg2lzbnLg+quYtFynRPnmlSqrjUTKKqnrMgJ
UE2vUbVvecmr+APAJXktWS7sLCiEhsfjQfdNiZokgwUVDN1KjXFtLOp+S9PKrNQF
eylQyZILMlIFOr8J+3xQUmoUbtvscIb8lqRva5iQTwtoXp7tUno0lUHPhXietToC
YesbFC3HToV6tZbY9NDUVZ13+GMNmdlePHBqc/l4kW5Y6k+ks/BtQbbbBlBz5NqQ
APPW5a6rliE5ePfJpe+w7cEpYHL6aS6FpfF6y3P30QW0QgqKzVEBeUelBL+tynel
ZEK689Twes/0/Qt86apxL+HT9nVofwZTQuy1A/JQAxlKkyQHh1NgnpUmWBNVRJE2
GFCrkbTDpAXxK1Lah+XhzodsFG3XunFn1f6bPW30fHj6eSw2y94JVCfosCihoin2
4ifTKvWbj4Ksee6aAZArnkUcYr+IsvIW9Gqsj3GdHYMJUCB/9T+/mBJvXF30JGHg
hYftlavV6dmivZAgS0aEWDPUu55E5zBFmlW1+EhPnQj1sQAwCKC9KuZtDBoxPVbH
uqcpyCetLXY7bkL8YJb+rrM0uU7kFuOXNjnU5N3xRjeriS9IOHs8Y+bA8Z/lyV9h
NogfXM592JQklIl3AR2NjUy9suytafe1r+xrmDMcTtLdQvevcL7wzp3N5n7nXAlK
zoImJPcH0d7731/6SPnB4bkYHBMh28oatI/NCH6q9W7I1b+DuwoAD/pQ8lO5lQPZ
PKPzQjwAT+MCveLfUbOM5mzL2rCBvOSMdZaGgl/oX6TdRHn7dRMhcbdnu//meuou
L/zAVxexRX5fs6b09YC6oTwalKJifd2rSZrzjgR1Vb8ZSydbKpFR/W3tx8ghD0iE
L+aTDRhnTrEAvms6woZyQIoH8a2MZojOtQWQcJpA82TAG03Q5ZeAcUKirrAvPeMA
CSHRCr11a5W3OEF0Zg3ze2fetQ71lMgeTk8wDWKbiXewnJoowCHgVeVW3kVlPwWj
v40bRZUgTLliekFpXACoLHBNa3WzEVgpLLhbA8JrnYfWj7quqjBVJ5SRLTqTzUoF
rcWirgu4HYlsMxSRuH4Ko04kTLLOa3u3OfVaI6dssLEEI6b4ZBhcvHqaUVFuUA43
LXBjUN3cIW6e0BFcrJNLnzYF3RvmEoGwy5OJKzEu1bs1dmDpYRRu0Z0DbG8xckPp
w5rF9mVoanvenkIkpAJdECsMlJI7fwcGxyHEJ+uOSO7feM3HwTRr5VAMthRB+fIk
FmuaaxNcxdE76gp3d6AbzYVXmkVUarc+BQDZV/p05r7lMqvMjtkuDpPKr085wgZ9
bc623jqldNCLCcuGItbt7OHiBwrJNc3ihMyPhIAVOQhEL8p7ICUlHRkiZ7Mepu4V
dl5mpcah2ts8ty+VZwHRMK7UryAg0B5maeqkRyEAVtYx1tAFhd+r1Aqoy2PpzTh7
dkxu8PVndITklGKNzhsSQV2jwlGlkOmF/9zW6xc67oilyHOHhvI9LamrxpclFkkr
IZFiShvfT0zaEHZa4ijwOFwPgHxxKcCyVZRNs/S7IsP0YF+EbvIY5QcvdHHrakqc
HyPF60kJgrnswtsO7dRQBJ9qsa6/UeUyMB0EfdhaUI2F8OsOc+2T+nfKXKWm6/cu
ycaDl1GxvdgzOWqSmVKqu3oP2JcKwJH0J9k1a9NyBl4U11aX+Pfbdfsu00CxKVtk
RgW9JekvHJhl8Uz0m6FVL20odODoGqASUSRbDw8+1im03RVucFF5OeiVUPOuyeZc
kj2OtDSGdQ6GyLqy6YLdnw==
`protect END_PROTECTED
