`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fzHbo9CjO3mZgf+e8M+oFMtJOJ0Z3OqDTPve+pPlQ6dJ032PCgHxzpf4wU1Wexsy
jX03ysba/tDihWUDPLf5O1a5NQjedVN/4/eaRcsyKgqwHG4UgrHkjU8WBQbvBuYK
CCtZ23JZ8q6J+VaXC3ajadJisEx/zy+Ju8Jek9qNNngyRqP+iF4B0FRkVPF+M/sg
NMitil0GcXeRMywg4Vh0OBTtW/y5vAlt6kiFMumsOHk93uSfuAVIXVe8rr7ICT4M
cL4gPQJ5FZeAmMVQFZoud9HO4GilPNsQthnP0aDsSjJ73XRzGitJQDD51VVT/pKN
qcvTGapQl7Opke1SL8TCdVa6A49r3vTqGX8XZjQW8YX7H+o8I2qrZLI1TmK5GNO6
VYRvCdH+5+QpInZur1dT/tw6kYGAfYpXz5b5OlW5ou6rklAvel0XqgCaVAZ7b1Fs
NCANjy8hkRwg5bWjRLOp/xXcs0qGP9qkgyHHYOUXAWgpYzpUirjwlgRDvj4pQ76Z
QqrSUJ9FKo/elfJGSWbYuaWoDei6qRDid27BJ0qTe6qfRT74aOiIlwV7gDGr+pJt
Jh1ha7prphW2eHEKs4lCQOt3Y7rCIHhTVZI/+wv80hAq0H0mtUVwCmFZrAKiYUz4
6hf7m1o6kJtmkYg20fPMeN5TzjCN2thDBFhxuLeouHQ/UhGRglIZi3RgqRtcq+9t
`protect END_PROTECTED
