`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XeqdUSrkfA5qUS52XRYsVG1kFVgnCPmbj7e7xaksmUFbbZM1aaKSTIEghgGpFzMX
kiUti5GNp8QweIOfS+fYa1CoLaCQJiCv0k+lbvtVfSHsQsNXmilM2fGf8WZy/z3X
txXTBzZJ9rknu3YSwPQzzV3JVbzgemXQwNjwxn713jNdZu2oSHtNpA/4gIbAVDIj
UDNAlIo+0DLr03g5yF1kzZpp5wbrp3sNK0+ZmMhH2p99MWu7IkRWyl95yvNwiIfi
LFRCie3cUF3ehneW1J2EkJYfQdE4Map1GciOxVlqHTslgdr8d5XjMErAspf28oev
NLxHkQ66Ulw6o92Sh2Jfz/W7HZTT2m5+/oNtjNEtpMFENg3xgC01V/WQ74v9D8XB
B87dNXvhPXRDXRwmGcBTVLT+BmcJSV1fL6maxKEyuexKtA/iqYa/lcc4mF4d2M4t
UK/tFYiiP6EnrdITslJNRPM1uwguTRfUgAsh9wT3WNnhDq+T3N5WRdmhtwEkfSwz
/zDhs2gPJ0Z7aSNDPncB13JTmOwpB0ufgPumXKYPCjXBUDxG3G25GsDVWhH/th51
ormPVKr+5AzzZ5g88MZsS6DH0SixU0VYtSEamJhueWAomDyrHr+URsY8aO06QCJK
h/URMdgpP0AaXtCv0LBMK3cKx8kZh2UOST04FycuDrcimHwflQIp3Ql8GWN4NIhH
+RwSc9/2bQut4+0L9kQs2GSoSZfAJffqZcKhc8c7RKoyEy9neYFJfj5ZDllB70c/
PfOvv4hKYp7hTW9565kEurUEzMoULY3TvNiSYmcMNzbVJaRKxJL4IQFw0ImawUJP
WpNMtEhXeqhjT2Kvl4urtWqWAOnFP6uTnuEoBE/+Gmyi6U4+2pvWat935D9PTVvx
rsp4OpqNjBdYc1/krweFPcUxp+4hZ1TqfJDPZ4zEdrBdaqazEmxNaz8Jsnu8upK4
HoW1XD9m+n8pgfNTeYDfwKve83rLcoUA8/dzw7BaD0Rh79hr+5rwt2tkXVcY0jXz
zuZ8ptxHToJyaXjQ6iwM9pCadloK+936M07V2x00LTj2LvdrgTktXCNdBvP6FD8W
Tl2cqj+vjVrhAhFxo2w5zbuTRfICBjtf+VVA01/P2Mqyxp9DD0NG0TzMnZz3EzC2
0pmllogYrPcN7vkdUvOuynEEBbe1vcHpv1WvasSCc/A6Q5/pkN++vjPwbVK2QgXf
jfQqn358nthZEPmk8M73l+qFKg1EIvZNAb4jJcQFJ9FRMG9EQ/uBTtx/qqoT9ICG
qnRNrbGMTXuHEZ/Ms6H5ZMJbMNRJJmxCXyyGLQSCDQdjLVAN0PmaTLlJE1FdyVbO
XsXYVbP4aQJtu8MVhTlPNl6PHraTcY/jEiiSffC76G3Ccy3gxaAo17egMrJ3Ut20
J/xOELZfy8e3iyJTD/qPKHBS8cAb+3ezajL7V2kHAiw01Djr4Oj8vrNdo9CDC4DE
Ioeb6Qt7otlkXE1qXcBHzx4/RfJNIOAtTsQZu9EdTw0=
`protect END_PROTECTED
