`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WEveYJvZokTlGDdc+bCkwNcQm2CxXSuFXyXvpXoGF5OfFAPcjhgCMJJ82fgHFpEu
dI1J7X65afUGKfXZHMGjL8LxlFmu204jNXNSpgJX+WgsRoodw8bX9XLjOHJ6SKaa
frpGeXxTzgXL1jL0a6gwF1DDxMUSNz1YKsR4s5sXiXu0FFYWQjwBQ42hko/sitAq
SAdLF1hWpIzCxoZ+gyPj7FI9/AdgmfJYnMviROnSPoZ7SrCeeDg9CTcQBBhlseRZ
lATrqxKsHztQLS/xyyJOP/Hk/HAw6Gf/Q9HtCOV1yTGe5e2macvqVUhSLLC3EsN8
0iYpeUJ8fANZBE6sO+t8gxndMjbJITAiZ//UbdsOlYJq+T/B4PwPumH76g/RcsU0
PD+f+EvD1cF5s8b1JqIMgA==
`protect END_PROTECTED
