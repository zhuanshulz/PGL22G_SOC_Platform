`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LFbP40h4BaTHvuBSb1JV03HnkqvNHNFVLDYclkFLd6x4zA2UTrIZ0Dz1tsOYvUK5
iHpKiRa/XBr1fpSZIk2pZtsu6g2W+sLLsjFqgN6hzHiJnu+Osy2gUgwiCau+Fy9q
kitRreIzvNh3PR8YBYPVlQhQf9VKH+a7pYOaze2wjOm37v5gWFHUkqv8KkwFkWu7
SyPxFe6b2zVcKJ41ushTDxamYQ62FiS2Hvl3AMMCLd9LiJBQ9yJEjJAHcto7f+FH
pMdO7W0RcCZpenZtQZLCi2P4AJChuL2mqBamzpso0odaSA3o6aB8C83+tyjq9Jvf
4WzE3u2pxs6SqSzULs4LxboCBpozBw1ecdcvjQmSsly+fsVL/uufZMsUEtnRx7Kq
zhR4UcmMHXYkm0L0S8XGvpznJT04JzcY6fJst5rvCeY6pl4rKsyYDH4VF0FdVadL
+j7tstGpgPt1H1QZvt/WPNTNd5tB5DbIUzqg5aGwRzPN0axc3w07eZAFkXEBibhG
pNwMgVMvR0IqlhJhIJo5cg==
`protect END_PROTECTED
