`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UCekniY3r7GvZrL4r3apbqP+Dr79adpM4oxPr13IEXKoYHO/Q+uS3iW6aQndyYth
Hct/tt50qXkS0CCFvayslwMAyss7MFqnirQ+03f/hIEgkpQXFPYFW6sIkQ7R7XEt
pDVxAE6KLLHcy4j44ZH09r1AamQy/lkBibzpwNb0Bn+uM8YAoVdjuMQndSzZzd/J
NLaTv8QrF+DsUBxLGp0xni3xsk5SCUErzr/VHiRvqKPQ3CICPO390knVTv8fJT7f
h5AXlGBL6gCJiL3dZm1QjRJ1fJH/pe0kCXNyQIZIfDJd7FS2kWZ3x2tQZwH5E/9K
ACTk+D37h00AydOL7QaS9301PpPcjnmxufWJdI7lF2M5tCU76NXy752XkAcKzPTO
Y5Bpj10/jly8bnc8M8PsKbv7ll96xQK8/GFiKe+gI4vB71hjsKyZymirleBKQOW9
xnnEv2XevHC+bedPHLKvgKweBGwqpxrfbpldjl7wpk+tkHJOFqZ3buCYQg3L/gsU
FU84GyeXq2sdixcLdv2bqulbT8tSk16CYrO9V41E3H2Ytg38GRXdTLvemGfftg8o
CKPRrpxSePZGuQOqu1IgAj75ZiR2tDM1Ng9Y44PTzpz+rlRjtZuR0QgF7KZEmTcP
pgoEBKjEvd6bKDCGmBARkAFsep2cHess03EXEobZkO53msT7LkO/msB5iEuwTsSy
sJIizcBf1Mj8uSKmxm5SnAF6AnA7Wu8xd0DIXdX59ZX2cZtNzQAtgA/1/0AdU8MD
rNXGqHoOO05ZUEQdZI92Yg==
`protect END_PROTECTED
