`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QcyTvKw5IPAnCAshMPF/WF43WUj7Pqewa3MB2zhr6QSrUVCeOAgqVTCf2wQcEtNY
+TwzYx51309YTz1NfCYq1FveCib9YqD3DcVcFB/An2c543f/TBznrAlU4MfuG9wh
FecW8NLWLL9w866f8WWQJ5N7tczUE3hcMQKo4GdDAUvkoybf/r8P2dAObRrXg1lZ
a4INAke1L8lG9uC9AmUcQU+yL2N+vaKDnLkCMU5cZpYnGH/A7cvpQmuV7qTSxFyo
KrD38UcySl5dT45zUzzZ8xGnXCYL1/PSuAB/h2cCId4urdE4w7oKagU9jYh7lysS
HBJLMN9/TSZTgOshRsKXbv+VUAOihmr9rjArz0dY4JOCGJiJw2tFS+dWlTPzg3/d
rpOyCmgRz15HFttt5sw7QTSX11oZ35Is6fWj8rLaMmKZyt0rUKbPVrBJ0HdYM7o1
Uhrs4z8ey815ouWzxwv+AO2jvsm+H6Q9vfWKFwyf/Tj7DvrQrwx5rDlV1+bbAG5J
YWjbyuuXj+lBZ4Rx2dYsGH31F1vV0WMfGJUvN1pijmH1R0jP4UTH4/Ha2wXXD8UY
vRjMY09SVBAwh+Ng3eYLAO5gga/xvb/0GfFEtgZI/uI=
`protect END_PROTECTED
