`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R0ii0321V47ZYFcAFsQZ/oXCUiNsZ7ZymmeLVjwBeUt9vawn6BFMBfzlqbEkT8fn
reCsmGYKuk8TK/4d58TUr4741OwWM2s/tNN/+4iiUlP8YziX859lzxLYe6cVrwYs
On4eFudK//L62vep4w1bDx0btS05Inz2dRl8gVGRgwDj5wdsOiK2D1UCpBOmj0UQ
GKz81iJ+1T+5jpXmPp5exCYKTSPDYi8FiHNsvPvpCaBc7cnK0LYWS1nLQdSm6XNx
AO1VpWkIWIfxH7CfSQxhCKZbe4qWwQbC47/L7mFAqZ9IWMoL/cOoR5k5523m9vJz
W89SjA85oA6NSeLGiGF0fTu9IeOSe/sTd7fiyEK2MhqoG8bsU3ZejdNyw+VD7gp8
Wm1Ml8zeFKY54tYR9Jv8j0yb7SAkY33ZDVvK1ZlSli6Mc36k8ye2aLShqahINo1D
7Ns11pVmHdZRdWWx9krb2BHp0Ix/jJU30Ri11OJwcgPddc41DPxp+fFJpMLjbuZb
/itVP1qEB86fWBx/K81wZVVOYvncQi7u6xrE+6iuYLg6kd/YV+rVl6g7eIioMRGp
9a3qUQaLxR2T8dny1uAKZAoteFCDc72ZSRVjYm9ZzsKRyICNybQsrealmxLPdsbg
FjnsHhznYqH+yxGy0PFhE06PckB1ZlbnyfUL0AFTs8j6BSdQG3pvu1wiUQx7oDHi
`protect END_PROTECTED
