`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JZrW1C5BHPRkVGl85jMIwVhhIYmDspTAm8MHtz7kwItA9T3gg56YV8u7dHOxtf3C
Iz4zRRuzrYvcjMhXe2cOoRZkU67fowV7cUhLjoBvJ4U1X95pNvfaUk9wxytE1WBB
tyRUycDPK0/JlAfz4/c04ZrSDTZmfER37oYC9pLQBpSDR/nNP4iD14O3dzUg32s9
H7LtyISpMtR7hBPmaKluOrWzNmsvUgAH6GliQHFhf+h7Ai7D5DmDEtoXGvLDkb7V
CIR+bHaZioeKSnjpE0KvYCz1SsjX0Ieb/i/ks1PJipiyDVupP0vJHpoX9terq8FX
+nTe0n6e+RzA2u+CHmsM8eu+XiyrZRYUfo54kFctAFdIVv5mww5XCZV+aIEJWSVl
10rOAeeQ2+rrTPe+aTz14ylDyTL8iN7q3Gtq9tRz0rvAUiOdga2/IQ1zRX3SU/7U
6Ui+TIDNYQvb7FgzFBfR5/px2MiUyzgrfHijmP6l+jQJQzIMsAmMIMVP6v6uOybd
RI8mGodh31x7crLH7Gzeq6urCmIw8dejHvZMWUlzaUBmckGXHRAuyGlGB1fSg4dn
1z/XLumlsVvpf6bjtknc/aguoreWePoCtCER9Ev+O9L4Eq8jUE2zvkdXlEaBef+F
MDi6UDZjkU0ecwNiltxQHrD3VyYOQME821ZVJDEeiDnWooFP0zc8CJhg3heqjGEH
Le5CN5qnB73XX829bEnndDrjcuw5BckfSpwKzUZpmINh6Nj4xdywN09pGZBtqFrQ
PFSIiZW8VqaH4scVEel+LTdFXcLizGVZNAlW82E3Uoo0N8CVxus9031OCfOtkJdt
ritS+cBTo4dQWPqzXHrMwR1Ou0WvYPGIijJlbsHgOcmg3MffwovOpsm3Chq27vhO
NdL67VkxSBE6Jza09kAf4g==
`protect END_PROTECTED
