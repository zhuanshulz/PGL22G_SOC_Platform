`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9+uxquaYCT1tQEhepwTZV4ptXmRPqzN1mnAxv/rW8tAMn2X4XydBobMKIhKVatn9
gaMTeTIyj7DVfxSV66rrF4S16CMb+/10Cc40hkQkAFh9q6nT80pay3ZUrI4CBmp5
jiWGSj6sx5JXIYkPCV5rtY9jQH8COToUJCwEaBQbvPZjQMOgItCOe7x3//ZoopMx
gtMJ37zhQLMD8wh9c41FPB/C7SWTQWSoDqR/i46UqmbCiaTepw0mgxaBAh57Hh6B
k6Gf2MCd7XKh3kvaSK+Dyv+C1duSScZYCiEpdgbtEkLOzELcDituzLaXn0rs+Ah0
7ahL0tlKNme7Bc/aMu0kFV/Lke+SeGgViUbrLy8oedBhn585Q8scC5rOV6p4zFD3
SCGgq1LKdSEOiz2UrfAQnyWtOHpp0yZKEZAyPKqRuvBnXyyctIol1NhqM6l9chRB
hby8tpwCEy/OUEd1MTz5f4qrvN6mm1/PUKyALReF7LJyIEw73SgOKw5Tn5TFqeyP
xg0/J5BOFPBtaRmgiMxR1toKUqGMUoseLBUGk9KkkI1pyylqATPehQP/5WsiMUab
C4g+wfEvAt00aEB3g051lcixcqui918Zj9PEAKzd3Y6ygEtqvoFEpoM5JOs5aCtt
NN+RaUKrYpYnVRAU3ERl3Ih8WCoaP93gTqNh9TVYugmwHuRyBY0ipI/Eiiis3cg0
VBJ9t2rY7AX51cDtkehNtyPA9PyicY4kYT0Zvg8OUV/lKYUMV40tr9pS6yXe6dyu
BhbdV5u8Otw9GwgM0zfnPwzsMmbEpI0WOnQw4+C8M0sNHW9UXxtCnBMFSMwFTKI+
O9JW1yA8pP2o0BTnEtWP7qzPu0IdHNN9Pt+GYtl69jEgDOo7blSLcl/s6t5zBIX4
bpbUk1qAiPks3aWHESrdaSQBVb/JSJfox/7/tZHTA4M1Cg2lz1gGVlaZF6pSci0p
37rjVmOHo1SKa2UDgYEM194TE/hFWTJGhD+CRRyClOombXMnZsyaxUI4VP1BiS8W
ySsLWEaPNDnPL+KGcCjcVH27DFe25TIHK19is6bom20rNh+clnkh8SQJa2zljG78
0a0Ik+AKhP+mF7Oy2SAoJN8dFDWTaNrkkcPVOqOrOtRGsrogE8ipMV6YwSvXR6J8
5oBOZD7XzTFcb6/jpjoWLhf44pO8QqGHbxX70nK/Cf1rEfN0MtOL9fIkmmF/VR3r
OwLZiMT0lF3JAxszfXGMdjRyLelhWVYUSw0mHxRuRgDJUNDECBbusmmRpkJdarkS
nlzScZqrGCL1OyNP55ac0q3Tm6+kWJ4Xyo/iM2CyqM2Qj8ntPDxy3hl8F4OLvSFX
FFKb0oAGEbf9jvJe9BRYOCnaHo5NV98UDcjGUZ/FbEvmTsEe7GoeRZUDiGQ2MqbH
kUoAynWrHRZsHB85voyuDkl6QVGk9qMG7meMJb5clOKPerHNiZptsBen5TNNK8zY
ELiOQcIbfoMHRzq2v++j2iIm6CAArUG1BJr2bad1ZIus/q8l0IPB4WG3tBaa1D0l
EJmE0dC26R3ap6aUEgfhUketa9mtJjG/qtPmxzA11kbsph0QQZkyw5b5T9378eIa
ghS+kMqf1DgZ76JHNWwruaFowWEu3H+fNkZujbHerZRrLUQLW0cKYB5v1uHHYuOb
/2j/UMRNpeHKlPMcuISf81+96F0aG4q+onE4pO8X0kk+7sxT+PBRpgNICZLCQh//
eHq+AdymSN4QZOFZIiXDoB9enroHVf70KEX2l7GBoVTVttLNegtZOf/CIFiW1VnN
Docyr0le2FPEhh9cYBI4NXWkCdRKYLHT3STCXhLHeb+c+YYRzWaoVDB7TomEi3RW
/S22coWGiGllEI0pRyDyZ+QL/BP4rOG5P9hqxaVBGyHvzvYm76hUkQJ3fYHhZ5Xj
AMyhk1aO++FL1BmlrOI4twD5sfeDcekegt0YjoxZESlmYmqIdnEJA271o4j/dHaU
HUUiMPXtIpZEM7izcLmAY+N2kwZ67LXyNacDoAYFubOHdKM6NQwEiF5wfKfF79mT
5VzFpDro5NIQZ3EnTSUj8M6cttHuhx85FyZNvlaHtrNzlFfAx6qWhzE3nV6XanUB
Y14Tywj24FT5APb6C5DhpmOa8SzdklfLaGIZrQbbCcuR3YM0ZbzTQj4K2RnkK1Ws
oui6C45BDqrSm34LFssTTaA//G+ijMOu/HWi3PDbAZ8ZqPuIK/zkWOeFiEOGH8GQ
YnZrpHCU0Vw/X0CLBh6THDRpXTCxx3acibVMkCF1ewhB9AOOczlBkU9PnbBwfqMt
y1ModkVXHcvh6kCy4Q1mQEdwj2rUX2aafct1C8s3nlOLHvi+gRpQ5Czjz3kcUVPP
omzk7sdzstq9TnPyRd0LU7fI5xwiAlGWJIeOJAHhbUsBA36m2kAiiPVWS6L7LwsP
ZBeX6qYrFoz9KfDsFc7oTEOkygdM66UUrrikjmhtrAHzMBLBIc6zMYmBt7xkKgqk
xje/Zs1/G4msApOTvZMnYeQYCUz7sINwZVLf371Wn39P1uIsQ84o4s/qDm71Nuu8
05n4Ai5Nm8lvCfzvsyHqBqrFERcEQ+8spmIhg1FV2hxWxMmGae220WvaF+7mu9zY
nJPer1Hho3V927h0Bp8ZpfchAMMfvDpdT36GIUgjfYVYd/oivC0aIIaXRH3wnrum
v5LT+Rj8gYNEx/KkIEvkz8bAXZFwXnT/NZYO0nNhL3G4fLYO7D9MD/Bqh0Xm1VxR
HK3krAYcdF8H+6tz5lLE819O9MaNdmLvvhmOdRfP3DnsUQFqacAZp9Nw3DsK377Y
3Re4HPZVWl2NuNmVlkgG0G18TSkyVTdJE7gHFD9HLQZbAqw/Ek2nj72L45Ete5qd
m5E+ENGJ3RQSMWdDYs1AymctMY3X6+cm/liVU7NK51UYxil7zhTkDHjlVEikqUWH
jjPxsBt6Btc2dvgb1Y15v7sP6A1bn3sCr6wb+nk7maKgkVQFHcSwWYnm2JWQeM4y
05LbMluq6QStztTU4EbpLqSCTn+qeWF5SOYflMJxr6nff6vq9aDJBswlk3/FvagO
0Qe8TOvl2f7PY/MHtlhajZ4zb/i2eawJw8X55FFSgIhW0EEnobyBCb60F3bQ8HBE
XgWbgiV30LhCIqK+r3iCOipJyVhpFYdNHZxFsiKUcYhOeJL/kSNvcElfEwUFtnrr
8wK972T3ICeiOh/wh8/nr4AQduKutVntP0OPb6gFIVo=
`protect END_PROTECTED
