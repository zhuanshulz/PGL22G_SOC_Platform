`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NdadTG/m0sMcVXyGF4LrwNbAioedOwGbRUFDy455Qd2nRl4x4rX9hjaC4KSETtGk
syZkt24ITof8kfQ4XapL5vZR5SAl6dUl45phsL8rsTJGQS9WF65mlK0yQmaDZLnL
zIHQUMnSB+QeowTnvrB2NaaTeMhqH2fROWcRQnFwzAZXjgJXnCojn2UDDlrPdelP
k+3UdYTaRoypqW/6O6/6qwtyR0JDk7CHB/xNo+jZPL7PiNolBSy77gDhWPZEv9tT
GYeT6g0F5tYR0GfiuS90+lTh4Ia5JaOEujYZcqYv7bd8sYXWpSztndUlpvl4xVkd
A3CQn2kChaFIDCiX/7pniV9deUgpjXeE/l6LbigGqJb7jcpjWMXvo/2foDkqcdDi
i7i9OlFOn2s2vVGYO34AJxTQlQQgQcKOjOF9LsHqbRrTIOBPvfrtcl/u0lFnYqL1
QzFZqPR4NCS1nQNdmG/fqmcDR88bwRfaTiWZUiHpHu2pm5eC1/knMub+0/2hIdmG
aHfmEPSyIHWVpr1yZsUh/eGFPw7P1BYovq6vmWtD71539vY0HoU+vSAS0S0WqG8m
/OVswkKcTCMuAkuqIxinGJ58jrSJKum+ZSds2KrUepQH2DWTPAGIxC6tEW84hqke
PTjGjJSNcetBgjl7eUCYI2kTNDr/th1gwS3h2ISnglBkx4R9uIy5410HqMnKdAfA
6TKZU7lbHN5Q5TrSwiCb5hJg95Da2NeKXvUpRaEHGicOz0Nur0haiNDa13MKiTaG
B+758kYj/jRU2NZuDQnApxDO+gr0exCDcAsLqc49t58NIw3FV76BG8M+mNAvlyC/
GlPTDmRmfE2Di30/IFptSxPcQrssLKbhGz3Duv3Xx+E+ND2H7F31oRWUXkpyWGL5
Ra9R7uNfN1bXWVbSKdF9qA==
`protect END_PROTECTED
