`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
thmtBTlAOjqnKfr8oramYItgsEwWBrwqbPPdJwaqTCIxEB7Qv5S4vlF6DE1lnDv0
5YExT9G3YECJqt2ksRAfBXCJwZyq79lVszIZvKHpWkAgsDV0gfom3PoO6v5bPKWY
z3jjDBa2GEIi26t4+wpxhF7GHPQUd+17cZae9JYWXbE/N/i5eVN+6EK51laTOY6u
TlnFUK9PIYiC6Yix8fzc2vJKCT72/WhpmA+BGcnGLAuma3CRrM3veBNXsZu/uqJJ
7piv+PmlY8tCdajrFge62j3pdZs3tTrnuxwKZq+xMdr7YDWy1xHbEQuNEZiIpff6
PXaKcLU7pizuBZYiQ6rRW2b1lhYVn6+rCkJAZ+2qUwNgzvFr+kHJcu5w4HSqPGWR
9+EH14hE+1FFwJ3UVnwB1vDMnkKKoLn5hk8WRrmGIteGCixStp6vPkurv6oyAAPu
IdbdJbdhDGkNVgmFb8GcDT5/VyaCaJH0zwrs+b4B09sGg7kiogxf/YDaa9pDDRHB
aFNnunz8+2imP/OfgPvd7XiyADfhTlrn6j4x6PJNtRs=
`protect END_PROTECTED
