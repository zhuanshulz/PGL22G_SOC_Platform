`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xOljhKIEMqWM0cbypVZpN1x9krcYOvq7N/xPF5Kr+9ZDKOqTmGg0JnyrqQONJz2F
vwzQmME4DmmbRp/bqAf4Wr4czLaW4lSq2RPYoRpY3sntkrITtlqwHw1pf86ZVY0H
UM8BLHfb6xzIPAyvXwNFYUok4UCXk+2sqAVL5monq6F9nTBi2f/YbAkrCP36Cq4a
lP6ohMKOwauZqksVoh6KCf1ZsP1b+fs4E2Yn4SnJcXz2esZm7f4WeAUo4jY+qhoN
eSMedXrWXdocQ+GrzscfNWWBtfd7bQy2PDIlvEmjVgFYEJ2eC/wF9bA8p38rq9re
vR3MugnLWtxtLW52KvSqULwkRd4GpiIhZWT111EQ6nnRMpZSjHWrp0QITpm4unM3
kfRXzrKuFzGSqtfm1zprawYf34qZRuNdDCKq6fr0dhck7IWsAu9NCMFYUMJZs0ag
COqWXSI+4BXlVuhTyKQkPuEMAkCMxqomRbqTS0kkeBISzwBgOli9qyd+ThINvMRl
KXj87T9nBgh/BIgiEQQY51jzOXfwHk+5N79aQb6tHd/6GYlQgqBbsaR3E2g66bkI
hW4OnCkkox8hOltRqMynt4KKSv7rPDHxc13QgHC6p/XfkNvVXj5jyO47OIZIsn6B
o9invjNrPF/QW5+/I6MhxJfpK+usk3koFVPdnupWzLO91AcIPVazCcLDTpVr+Nw5
rruwryI6UOAXovr3E9qHkHFJCVYSyauoXdAny+PRiUlZpR+Q8RsyWPeRPYc/g1W2
vSXg+DdiM+FV55OITWjymQIpcG9l3O2fQeyQVMiv9gozUf0d2y3Y3idzj6ReOXBm
c0BaqBXVpeyWZJLmcx7H4AxTMd78mAsEowhPJh8kpKlovxi+0HVz/Ckh+zjHHluP
akdG3SLDvXLzWzk4t5cfxrERdjIPouqVxU9clXXIoGE2G7KryE9Jg/qbMyeqKacx
Rgzcce12LRw2fp1d1n/B/w==
`protect END_PROTECTED
