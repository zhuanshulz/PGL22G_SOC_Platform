`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TFuZ8H9Hav/snQaofs168/9lZEttHsz63SWL1j4XpCWbfjInblYFQ9PLgw4rE/af
MGa+5xJcXWm95ujTCzp+1PeNoMexXLogs0D92pej3MqOvOkGuzX1rty4wjxHJPwa
Mo0I7GtG7yByw5SB4nBfybWKEEITW2WMsiG75ZpBrg8rcWHUL1PmcCI+k+v00tQd
n2q2oFzdGretPFHEEaNTlnW7Prel61/AgPkh6uyFuD3qNpFX8Ygc4neEZe7z8S4y
p0IZUrVTtNGis2+Gb34PQNZyEHMYnYF9Bl5BgCTppkLAEe1QbaWyvvfScLdLLFE+
mtawzaAA4Q1T/NNIuHLYUBCu3ANWBSK+pGqa5pq7W4MQgp6Rahs3ckTQ0FVKkFqB
mPYiRIxiXxeIM41h+mS08qGUFbmnLcRS1CSUZ5HMn1Be1uG6zbSIQeCw0pLRtjrq
YwM40SXJZHKifSNRsGEgd+SS/U9tCfmx75TGsSukRXer0s3OqxaU/FLgdfV5SS22
u3o9eaYVRPEpkGa1t1cMtCxuvRGhg+DQF+45wr5NqJNjD+OtK5QJaXW9p0piiUyV
ISV1WryVbvEl1XuWZEVvTAqf/x86qOS0r2mKoG7hhWd0zKtGkUcUo4JOx04bW/tc
P8qgW4iwTN0QeC+UlDLLEw22p4VHnNvkh/hvgE6iz5a3vuk7BD7wS0DOw85bKSv2
cIBXjEUagLSziAca/iXa5btxhqqc1DNxOw8omRyxmoasHs4cL3MdKIIQA44KCgPT
DFDVeO30dbOH8UfB4I077pmH5q4swsFkz7CMGEjAtolFF04cqeZ+Lmay43kzzV7k
hhuz26I1hHqhEHJrYLmSne8eBoi+5Pjlbbd4IEfkjRYr0KcD9270Ou6LQ1ivHsiG
rOvc52K3mmLAcJMHfgDQH6DL6BskBJksqhadoysHrknfjvLvDu9srlN8kOolE/Iw
akAllOOI0yhByVVJTDs8ieC00gC0lLARxBbHzESAGMSyS5RqfVCq5OyG7GWnArLN
RMRVwQzJA+77XXk9544ayLqsa15yhWC2eGfB/PawzT5m9uADUdgbUZAABleryLZQ
SprPEJg/g7+LIjW6FlbwbkCAz0GfvR+SW4NiF9smti4yJ5GDsNKt5LMLbsgYfFCb
Lho5K4LQgqMdh3mBeWlQHlYb91+uXXU2cePYTAQwYWPmOf5ioZAFIwSiNoyefT/3
0PAS1cZ2An/bQ4y3E/U91dPq6IINdvaHzJwZ20Iz/eAl+PPJf8S5jvsvSod+1Ahs
CeIGR1wAgZSYk7Dtcxoj2KTUEA1ewbodJXjQz4tZR7dM9MAzb7w7j8yD6AmgNoNM
ZeCa9pm0PjrOrp62wC01YlVuhpghXyk6cY9bfM1RleTVkON/IQoC+DdacH4jg8YK
nsK6p1KNIPqGktZgYTb268vcygKkqwBbupdEdnwfuIZDVQ3NmiKIt4l0eslyicvo
IVOUhOlb67w3P+OzbdBr3N7mT1b5Mxe7Wq6pQQc7ErtzA5tWIWuuPM9MIs+7BYQ0
QybDKSegKG/n3LjRlV1g/ZRCoOuyJXZ9taGWHWb/ahuMc+saV7+ZABxJ6RC6v5VA
15KLkiXBS8vOCgxeeETckBx8nP2aA48KhwE9lWHBP1tXQG42r9jW8Y7261jRx2j6
JibWTXL0+9wRU35a2kWZyJvHHYh9CHu3ObzDX8hYL6qqlkyMlRhSqvtwzg5oU8hn
w7809/lvxxdkda4BManDnjvf85QtK1/ewpUiSCMBHCo0Vknc62B4IfpbaUSXzy3z
R13LYTBbharIdKcTHkBCYSmTPRVYPvGnO8VU5dtii5BTG0Vn2o+Ek8pJZXR7ANQr
vpv89c9/aRybC5RYG7gd7uCq3DK7ftP519LpqxhXZOXPKzSlTEy6JHNdfRrRJhiu
QzWF5l+dgkVpLpDwZg0mE7Y5V0XCxyRGds/FIiHsl7B+BmaUXyEoWAxg9X08/Ep2
eOE4vgf4j6OBw0LJMZgCaHWF/NIAkhGXCEQw0o9QqLzcDGyaEEsaTN/IL0dpMRCk
JB8e4QOrDvo6VnRsK6GKHaz9NrqINdwNE65kkSPHBxtWxYCuyx+F3gr0N1WuArJ9
WXdZ5nPLQh2A+FRXQUmFc9xOshLKYOYE8AMI/Amm2XSJdPkHK4GIp7lA4jXZgNaM
isHMzzNUzzvPcE9rhX37dau3dEg7mFrdP1najgZjOYREBJgLNE4oDpIfLAhk7npG
A4T9px2oYMUujOhqjFeCiMeEU2C6iise3gZad9LBycwaDecXWFlul1RpB3ze+6du
Io2OEnPR5PYhgHE7hQoAWpTOCySpopUujIE8I8Lk3SIjxjolid4mGaoOawnlauyW
jWxZJtm+dSaiY9ziQAyy1EHdnz3+XBDUXLXOyldHh06i82+tFPk5YbWftAWlmGg9
l5Ud4EuCMwple9rxNEdzFLwrABGXEmJ9VgnQr3MTNWELioCvoZZ8yfbQIcOfLX8k
yv7Dehlh/OfM4W01ITIFhxVM+a0dv0tTdUH8La4u7nDDx/6pKGUbpJRZ6e9CoTes
BsvuLzjvqHu4rBKgipsk6uGGZUi6n2awDUmuSLELSlGSkkkzTKnxvXM+kibUyZH/
9TaeUjSbTj/2+xiDB8GCvEMGh8yH10F1qiWsDibXxqjrKL+k4fAXj7t/Ef1qo+RE
/U0ybANj3lAT9xx0AERszJdpodSUvZ4Ald/eik9iGBEVaSKW83Xz+LJdmePBv+Ew
U+me+DJ/68/9S4kmFjF7mq7Q3C4dZPh9IETYtJRRP7ydvIsSa1QAwtoJ5DVi1TtZ
wMrZGfk6Ayj/kQbZemA8IxHrK85UDJmIE0of5z0msoh0tJFRiOwG5Z/vi+x7czyU
gimdy1l++UGdYu0vtdDmxwS9m0PLsNNXeznrwxhtuyDlFmfZ0V3/jBEu9cS6IKpA
H60edsrZQ9whNksnGPZHwQ==
`protect END_PROTECTED
