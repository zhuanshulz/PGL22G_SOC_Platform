`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y3RMwj0H0zLyelX7XNTWzosijWS7HAvluvN42tqPJ4OPAynldkyBHENWieA8/FKh
+G7Jz0rqH8Qw+lSQnDvoxD2Kn6hn8Qq9MNzH4CarsiKYJPE3kzUCz+P5qvN9KtkD
qDNxDRHMlAci7ar203XA9zZ4xD+YUlwmpePjmc5I+nNYjEmXy4J6KqKmUoRRYdzR
puhOr2x4kT/DnRaIXqGQtjnt9hD/uLNPefqw6Yiuy5fe7LyZUss6FHdf46q3wjR4
AKmyJoWi7mxid0fy0+sZ0aVIsY0+4mTM1ReT6AyjV9gCHnNA5DAK4Nrc1Ew+7N5t
rm0eoYzfieCfE3+oZpzLB+xR78yIYZSdi7gfZwuH67LkfzrapZPvzSuQulnpUxUa
TBKGHYEOdBo97uPN7ZCUfRwjaE2fo1kl0G8Wzs2g39xysTLgpjSM5XrDVoTQbIGL
iQJ8q/QjQn/60xsp62EhKPxqaODiiKh45xG+T9Kbq3IRSTB5FUQIGC+COSfPSsdP
tGn/sNe3JFXFPvo3vDLTGzttu4knSAdt4jQO4jcxEPt0xtQIYWKumUSzwUjexLzU
zsleHJyDGqPgPWHq5G6CoZrEO7lquZq4z7+l22kFQvhFFxKopZOWR2/8CcS2YtpW
/DJCXihTGlDF31T1CprmmaUASWApT7e/Hbo3Gf8b+QbclcFrCuq9bbx1Qhm1hF+b
URsZvmTWRBln+X5X7p1Km3LlatNwpoaFCtf8GNW/RriW2iTZycS4psMmmjFHQl3/
L5/Wb/CDK93sAIYVTGZK2lDFaBfS54AhpnVb8ru7SH9cYrh9qb5CfizZueY2koy5
nt8JyEWGiVM22g+lHAu+gCRwXtjyx1JdnRJgSXtUYcleX2abw/tHBTaVWBU16ID/
5vhFYA0cBpxITv2jiMpGLOW0HLUQSwvLsVJShtnxade0MXkCGxx7pwKIw/OJn2Rn
GxdbBXD2XlLZzXheGzgesv6PjoPwvCvr40x6jPjP4aS1tgmHWxE2WWJhK1pl36v2
GH4i7sS9ACB2CVbXRgui8gFOt6G7fuuENsNGudHZE3jG6Lh6v7LVvkbJPFkU2eHr
w+cYiABa50URmoarvp2UX7zDVT5OYbkGphyVCV76AKGUuTRzF579rU6qCCM1EcvG
yIlIOGkSMP4wZXhwRvD9wN5hF3CXfQG5kaDGa9IBWde2iiQPhEXi8GPB2k/d1FM0
gK8S4IUiXfwvvgIUSxbw4cQfZJFhPBHi5qWJ35M+BXzUo3jBBU5CH4sPOQujBgL7
WaGXfyxQZADuqgZENXxoQvL2QjmEfU6+5yFAGyV4if454P16xx6JmayhVFNyXpKk
JcBhDjT2qOEn10Gi8h6P7yybwYCGmuWX3ofbhcrGPSm28VBDbHnVXGsuC9D7iRFT
tw3sjILyiH+2ikCrk+2szZjKzU5JjxK2GYMgfv+8XW2g0rr/Z5bmUmTxF+0bFSaQ
b6fz7HXJGXVGN4vh3rnfA83xydLY7g2ivMvCJ4vHgR5E8hQNwrODDIiKm1KMQQBm
hJA6E5Fp2gWfPHbuq9V3Zj4bAQ10YRqwPNFmCsTGnkdL0nQOLobMSDkC6rOz05ii
3AtNYE9Zi40plTChO7dPu3qgWQtwjSQzkDsPUXvlTh5tjWAzYHe6ezH30Oe2IMDY
4Oj2sRRoo43giU4amsYp1RQd8NAoqavbeqZ/P//+7BpWJoEgI1NCqOXIz13WlHG2
aNceY4JIVBAOoN2fJv5MhFcb6qarVEDLKEfZOHc9mlqKPDOT+qfH+2jLGvigwNUI
CTuz1kxLnoeXm6rMYp8Ye1BbcuroefJXdyovenalPvtxj9pETQ312BfGM8EV38hC
GlkYbNu80klnwH8oLyCNgl9itx55fyf+AiUhLkn7bj9D8Dwm9TlK72O0c08VUH5X
SSvgqJYLWbuk5zBmxMCDEg+ESq3ruBSIMZiZFLOfk/48GUTqp0kkoMue9Jo29JnR
V1Bof53u3EIGpPDy0mxXMEMqDPG122OvbosJHIlhrWs8Yc9DMyKB4jP8paSS2BjC
wYbAnVxK6q2bSkV2ZKPzoiUsbOFTv8cZ0GCWqHgpk5bWF/RmfwGE6maABudo2chn
eENwAPs7qVLS5Llczt2CMG55pRdTIHZFLb8oqThWWymfvDrZjuFUYQKKgZvCLOuj
B9hYFBuMh5/6Edvu3l+CAuu5ZNX0TDiN28UdD2DDQ5zPYz1pKIRhy5vdJoKq9TDX
3VNGoZ5x8Pec+fzoCCkC0g==
`protect END_PROTECTED
