`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3fcKgegeI3/fNjXibiOk1068S5LyMl7V2w62x2Y5tsK4g26YtCMSPWT3jp6OzBwv
f0L6vLx98xx6AfdDJjqjIQVp/8OKAFz1zPx8OgZMIkvPLtynlfIKVw7O/KDJfeQn
+REUW16N6MCq/hy44DzsTpawuimkTx5uSoSevh9PCfuh6W4DJP0YLyP8zkn5gkfi
/k+a95NHuqFZqowTOBaXBBMh0yL6/xoO24WHl0TvnJ2mow2hfId1Y9N3nsaL4zV2
gPlBG9CWXCv3N1nLVWtpSHwSx12i5K/orWeba7Yp9ksf7bUQQ1Vrtd740rnNBRMQ
DncI6lLMxp7zKX95fHBoiXTds1/Dy/X0raYD2/qP6kxas9txH7kUpDMQLf/Morwg
IOUqnSUXH+Q24OOoPXzQFcEY1WoI1J0rPEbi4i41o5puD6av2T9R1UHoepXJEmQR
J/WVapyVT/0NelA6ywbiinUPAYVmg9rppWXkDS9CW3P2Pyq6pylZGocI2DJRG87d
zBES1L55sTg3sbxnIbwWW4n56G943r75CrBB3G72pKJWNSV+G9s7w0hTtj55h+1M
/IzYBkBH6yF/LOi2Bm2dFiGKooA501H7DwoHCDPN7UGS6m381SmYJi7MQo/grFGH
h+zIR6oSQRyDzCf/1gSkoTYnxhSEe1FRHoD27nFiydhBhr0RBpfBynvPCTYkpgNt
/NGogeHYGwJPFmhGVlyffolzaTz5Nlb9hXYeWswy9c5WruVBQhP2HRQl0ptg2Dch
w+2Uun1dxYbrO+UJuI7s49Kbxq1smN1fbHWWje5hG5g3x5U/5ib2pOQU1vOwm/WN
Jz1W0i77KKbbY1h0CfliBcg8L2EInBdMaP3QUWDPbreuDHMnBMrDxXbW0TdwjDhs
27QtFuhA4aZmrHolgt8lIce1xnerMz+iKA8CjIGosT1+B9+u/JvMSU70+l3aWNHd
tX+CR7r+5gnzBEdle0bdB/2etKWEX9NNbmBBG9fF8RX1Cl7dMOWXf0AIwnImVxaw
`protect END_PROTECTED
