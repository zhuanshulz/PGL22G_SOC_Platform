`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jTmA1z+d7BW4UMOjGRZjKlOykdKmGdwpAwwWrp1BBJviggHM6hnTQ4gu1Lgusvn9
wiZ45lkk38cEQQ/gtDxHvtBVTqyhGQJ8TbRZ1AICknAjKzl53zRRKA44njNhzofX
cuXvfzxdJYN4eksDv8mA5VHHfYZIXg/bgNI450qPSXJsSkLdv6zzKe0Q0jgdqIOH
OkbsAuwlXkCz2rCzspXNcNTzz/QCm5ZP86KhDbvPS9t7hhwF6M4geI9vXeu1AxYx
SxEwkbBmgOWcELtXgM+SlFewaEgCOde9fo/mB7avTFKWINnIYKAg4d7XLGZTW+yA
ECZbm+F1IZATHfJWVD+Iz8uEWq59lPOmJ5tfAo6vvKHMQIGlhMouU1EZZ9DjvavX
/RDJh3VC1J/weCzutCSryhQ7h7KirenjL2doUR825BxgC9S2qx+afxzexRS65Wv/
8bVoTmrTJIcN1rDwbcB0kQ==
`protect END_PROTECTED
