`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9+zvmQJ1UUDL7ZMBdaAAYj9w60i+iGoiaiYSrlajLEE13BcJ4loTC0fcFRGswBlx
nQohCg/5GNWOO9wf02sXbp1GFhXxDUFpMzeJ4ciJapD+eWbW0Ia8MBfPT784WUWO
f1X/GnjCXtxlCkG4jOtnBO6xc7wJ5W/sbDRMfZ68x7i5aDy+dm2uPSa613wU7bR9
BcgdqjQRdrdiMyP0SUs7gbHYgcF5i6OLfkQu92OEF6ezS/UnyIOUx4LEmF/5vDyd
B2/O90mW2fs8jZKyvrRJkUMvXKEPZWAuQBzRua07tW+jlN2lv/CglRUY3MfEl5rC
1UAzdleQ0Ew7pPlKRVC4lR7qkusZ42V8cPtPvyKP8iSK9Q+jPYwltoe/5cQPalr9
fvNv6wVaKfQyoHsfmln2WfWDT4SNjggOJgzN67opzmI/pmNlV7tSsSHbpRDPwcMS
`protect END_PROTECTED
