`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+TdIPm29gcIcziF75oY5itnJW4aCtkIGxZsk0HHoAfL7n0G/i9ORkBWji6cvFwwk
3paixyOqUAL229Oa55ZYgNk1vTNbdaRIGiHYQVETowqYT/v9f/LpNIbGF29OrgS2
s/i59K1XB5hBlrorqYoYDl3DObAuinR1u2npEyFTnPAK7CgmO+4w4rei8nEmwY/p
IBYxxEqUZR7WO70tmslv+fO496yFseuM0NteeIvsUj4F7OaAYRS6dfdOw3pH1avN
luSmuBUKeK+12T0+SR6b1QUfDcZyHL9+yiK+4w3YuABIgqFgumKpsFm95PFmnkeQ
RKU0jSNNA/lTnv4bSW0QsvR4E9zcvVBmJCMpDZUuae0lY5/Baad91HMQ3ijdvPxA
R9BAJFFx5hMm5tCLHjv4inXNN6ERrHEkIoH9FfYHLbznPixYFcWmaQ9wEJRYQjX6
FIOSnKE8gUbrg1j6KC8NSBPf4LgRE2oTWs4ORh9sVR+SWoMiRvz1hRNZQFQCBghb
n4QYDArpxyQoHJ1QtP7GpCezmomai9/sDdOA0Csw8f7ApjNaoDf1UEXURmdZd6oN
oy2Ex8YabG7fFD88csbt9cYcLFshWE0RtbQxayqaB6iJQeKhsKHzJBdEMjMySYRP
Nl6a7wkc1qC/2OhAtrYrBcPhgM8l2j/Anqk0UogTzSqUiMeENlYzjfKQdJyywEeR
OFipRcCJWbluvHZDor9onvG8yrQ50KPimEasHcGdsLNWGXKfH6Dv2gjjB58TxQ+g
4dBisTTouvdYodaR2ldiAA==
`protect END_PROTECTED
