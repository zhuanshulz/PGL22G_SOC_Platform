`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Oh6ch0yKZDv6qwGmNGxbJ+YxVbeDvkOQjHtKBkR3br6ypTyPALJE9IYymuTut04C
wFVOip80aOUlMi4vVDyPjVD3cBVAhAD2Q8Zt49z944hwaL/M382jud9ViqRbnMcM
RThe7y4cRyarWZKQ8OMJ/arKC+e04voduka6Wynr5AgoG45Tus+kY9GCBjHqaEAA
CWOvc2R8ER9o3Jf1ToeA/kWFfS3bK6JN4CSaJEe1x1067461L3SF8vXU2J/X+49a
vUZUylOMTz2AJ+E6kqoc0GKZMxZFQGbBiTQfoIkyt4auhUmcI0/SCLx3x35j1HBW
0F9I0kVPqBr8ckW/FN709olRfL5BfDGSitJAZGTpNsYqUR/eOVgfIxh1Xm8+EBIw
dnnObvtGD/UIJ0EOQESyUz5qCYV8PN2doL3KiNKculejHD9MhCki3n1OoJnYEyeT
ye8+B0BlxXuikdO2nU7GwYr7YpxapTmSfjXCQPCVfH0JZWgNdHF2LFDjZiD86MtB
6H8eH3PNMxDNmWikWlM2g5flbhdTcMiI7OzL7My7CLM6TPH30gP8DvBhBUNubV3X
P0D6l301MMzTGrbH54GUtFTvqDi8zV3+dFftIG8Dmk23VOO52zRESrraizkjurzv
R5jdA/cm8Z7PbVfv+8IygpEmFjmM+CT+JrhmD6I4j4s2/HHdG7/WISBLlduyhubJ
NjeSfSDLCyN2AibCAUZFpGW3LWTvqLUwgNSBUFWwLZoPBmLBkwPYisn5HjfGZhIM
32+RuRey3LZcmE6PSR7i0VdFF6P3g7PecLhaF6lzLjoFDXCK+whN5Y3LIIgFUAWS
8FWB2X81V8s0n8G5f0REl9F88g+R3bboY+sU26NaBU0J+r06YDrjd1pFBBWps24x
UsNrAZ4ti/52j+LNeFZKqMIpOBWSSm1riHgSOEFDIcFEPv//MBTDwK1uYv6uBcAK
oiFj82/zmORo+4pED0+wsg7r6/5WtAImN5xwEQJJeJIwlLbT9fZsl4KQwL8zXQ03
axD/ROVDTgew4LhunPn7JH091HzBdW6mfAoansJk5H657/gnA4h0+9bAttIXCTV7
gzjDoLWVqBBXoBsN8PWiKA==
`protect END_PROTECTED
