`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BDpC0QTMnCSnoGqP6fMysulLpvskZUsF/oxgTS9DuNhSMZYCTIohLsU0TW08ZX9j
m6b/4+tyijw0Z8xle/1JirGQKe6xUE6osO7TgHmhEETDN234RXe5KFeyPglTcUf7
x5IM4UgASoRVV3MYB55h4O7rsKi/TUB9rOu4RWXk5ra9UKSjNm0eUG0JgYsNrhH7
KL3mrIO7yl8QsZRr8+QGL/NMH1/kynKkBqdq8NdzMkNr4dxiUcY7JXUDTNbRu/6X
fbwOEw56AdnxMOVuafaCVHQy59iBLM9yUV4lqFf8HDlGCOEknmxpCbPh6KXSh+wD
cX+PuBYdwhiHugF+zqvfIDz35EG3jSoBf1Z9SNDZhoSOocjF+FPQGvkdLgrAeSoc
x3/YAYOLRNaBkZ4Gu39X8XGGrU4JJGCSr8WSHhssBlAITz0O4jbiL7btfjfT93yt
S3tB1Q8W4PUWmyRNHzHOJLhgF0EVdPBjwqZyGO9ENuaG9eSVx+JnMg33E81m6ADr
lcXn93+Klq4cTMt822RJB+W8hwIwgofFCEnh05J8b7k3ISUq0NV0NKAS4351ooPw
y25kD1/5xnM3FWzm7hAaW4rFsAis6rRxianzITyLC+v38LceW2DZRwrqOnChrFTC
4CkGvqJ+UcRaM535jn+oA5zpADTgaukCz/r0eddsvyB70lBX1iEwQ/5c0VvyWxhX
`protect END_PROTECTED
