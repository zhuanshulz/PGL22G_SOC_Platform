`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DGSlwc1g/X6dU2VW/YA75JGTPQYf+ktYHiuwkjqITPW2fJqOQiihlYH2g0x51fyR
FYF4e1xNltcm3PUsCW2w6sl72LQidvuxsslogqbtIIpbF3HfwYsxJrraZt0pKPZ+
CsOIAZ/4QsOGLyV68yGs6bWXZLydvv3NtG+lHEwj+4GC/j7kECxD/0GMlsL0vnFK
zpvNY2SWqWhllklZa5dxJK4phK0TVvCSKN4oFbFC7T/FLqTEuI++xFW/7FO4F/CE
y8IpXHOd8W+1BjMWlNC8RY+yqeKYcLaa6DiqM0baIEnSO6/ZfMrxkTUF/SOheZP9
Hg4FJ5DxPS8AbI0YYkvtT0N+i8nizZEXnutMVhv3OpAdPKfBpPPaRyC9RCFK6Jrj
XvyUUutE2AxAo3mdkz3RrnuPM68myynVF9EItkC+gGC4FBGnigYCdFEPehqO7J2K
65kDefyiHmgP7bjqKtpDghLtQDi0IUFIbDRwTzvvpWgL33kJpzRUzLTt/98em+bh
b6XjhHnXSCLbiUIknbYLuOKwgs6hlUo4mOy14e39ut9/FZc+nGzfkziccjkt961U
35tSZrKD46cLrKmIJYQ82V1PO8JbKqbzzD2tinfnM1pJilemCUAIYrNKJgn9PzbI
vqiQgbGGo2SgFULNorGUGeJUHq1s8fuexoC0XLPKi0wBqyPdrWE3EqPNM/BEhgva
gEux+g61gBL0z+9Q+4Q7q42stAYtl3LtYcoANxyc3ciVF/JWqvYFW3/Hkc+x4Tw2
G6CznOBWCqeyA2RMqsY7FZ5upfjeY6C89BfGHjP8WK20Z+xRlDNAQpI2TA2ELbFB
e4S7CBah4VKUvWhSoGvt1Zf14GQsVVdSdrN724kr+lGrgjFP+rSlvJBaIfG+jHmy
aeYYZ6x+OrglvEm+QJAg4cHFQfAGWWPfW6fIfg/VeAz1whlLN/c7s3yJC9TJV3Ur
SoTFsJtCd/zoX7FnXXIf/vvlo8s99GOf7ZfzMF0GABHWonSwUn8dfBGs6N39UmK1
0BNWzbhoSrIFDn3TuRu1Z5chu+WlPLCjXIizM0ZeF/RqGMIR1czCx2a3DoypJlNC
sn/9qeVPOac0BztmtHR0ynxGzW68I7/a/QarFn8sRgmCcapoPlhdXO+iQmWtrgsc
0sbpRVa1BsVUlZByKbuy+g41X8POkf48LzHk1c2mELaSjghguFFa0OGuLkRFQdx/
fAmwcs1WBUY2LL27A91TZBblRtPfif7WFWSHkZDjBw8eXUOQ0RX++uBVFke/etZk
y942ZEy8/AMs25OVdlcsLDDXnw3vj79sDifuM+Mj6Lg4LXvJgTczkoG/tTpV1xwr
Dw4N7k0nxqLHg3kwaHdYBcwu/4IQBPenAnqLUBIdRQci/INTCHWn54Nn1R/gMa0N
/vsHf4bN/me7UkP5xGSJELdcbRabRTscP8CDzNyTdu0/l3lCyK6z4pIPiThUQQLK
Q1j9rBGjqE6DWn1D6ivTJUdzg9yGIQwTqUZs1gg4F7qI4DySlnnQlmYbbEPmNpC7
tveKamAauB799EEUsFLdHbuVK5TVn/Mpheg3V77+vEUIn65OlKjyvYPcF1vCvxed
stvHfGLwF8iYe9BOCw9FUo/pasei+CFfof9+y/3ug5eIA6XSXrPpKUUziFyd0Uda
YEp0x4heC8FbqWFe4x9MGkcb3XU9IJ0/GJfBd3XbQDZTd31G6zb5lHQXWDLGrR+e
ZsJiDyRuqPQolDeyIfONqhCvqnRpuFbk2uqP2NOBLlpzQw+WKkkno2uSA1bGTF5K
yxzyGuqW0yXY9v4nBRnuGchldygpZO110Z5MqZDZZ3Fc7Yzoq2G/BfyV+r+d7/SE
tLGMOOHiQDgXku29hhmowLpTT0c0dv0rfmNPm0Ewt06/8D9V1Dsu2u5weco/9UJ/
JrS5yL5tmp5OeDNztOdNZxr2okiB/1+S4qvIifKWyrtOIyeLl80luYTedbUpb69a
9EppS+GR7F3bybi/GvMnMMaqpOBAxeZkvBXh2fA7a93W5D2MI7oIkAQjDQyorkNm
H8UkFaN8HjQCuhQTbRl0oEG5AABoCcxLk38XH/2nbD7gXCFbhYcrqUNVi4wR7H6V
5/uygY44fNG3uO67n15/fCyf+wacA0U9tfELME4phGRSlMEgJztwCT1lx+SCtfAA
DFqZF+HyLC4FA4CsTneH6J/TDwrLe4hOPlhIQsZKwYuqt4upVFPjGr5CmGZ2b4md
0ZwCE1cSuwy8C4wIhM5iqdx+ssWY/J9HLx1PrRaaex5Gb2qmVV50JLg2JJetJbT9
Pd24JNyG28qfzYJQXMrZUnuogWaDKiQ78dXr1OvL0/VXb4mQe7m2mQaLG8kE5qrV
0KR1ifn0KcgATKDcj1SJYMZCjFZ+FFLAwKYW6ife9QoZEUZu9e+NA+SiORBXTpPE
CMnEuZa9hSolOWBa3FRXGGaNxL+zeiWGIMPxoPXe4MpZDnbZYkN/UNMJHFMofipD
G8a8F9RNSlYH37gR9VJ2ATAe+TOfPgczFYDjsPGz+FqKPwnSyxYFc6PYn8UebhaP
DSVu/Ao8zpBtzKC6/9qtgIoDoO1WT4pcSqyS7wNMH5M=
`protect END_PROTECTED
