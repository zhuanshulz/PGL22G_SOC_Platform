`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V5+LdzgwMzh6qKBxsVKLnDPolUWBjuxR2gyBdZ7mudaJoGopEhCesVNoGUp+g9uW
6fxLhuCauLa4iGxXNg860p4sMjt5qlrbCYTYLH4ZpWh00xjIErUdDFXXjrgb/Eyy
7Vxdcz7elR2eqao1625hj/JT9Tm8cU+D3SFwPC1TUrFuBpfrL5GvPCi9PA4beVRR
sLJHQCZJoEEGZ/4Ev79nqWGPeJD3bIzSpG53hD1h4z+AlYPDKF0+OcBzvj4SeJSn
FyzU03/F5+xfpqgvmy0s1rM7jvSxj/dpFyScD5dwEF4bnBE78rlwKpqiack1ihqZ
JCCQNDI7OjoYtf01Z3TaKeHGddggTaXUc39CpLEuWcHxoPoYiNYnDk+RS1fcpaw6
ANy6weQFRGR9g1lFK2kPRwFbumUwQi/V/eCPsSl8W1CA6TumrOQQ2zrwpjmB/Un3
sLIk75wPFAWioijz/XNs+VDjG4lD1a1Zn1b/g8s6sUL3AcLuC2lkTtZtvTeCQ39o
YFC3OEVxvIda12kc8tCgQXBXe+hp6ADei33isZkj96JkdBaVZIJUMZGyh/3IQE89
ruDl7ONczasJdWB9jcCCN9hsrfMeMlLQ2lNW4YpVH080ON4e8F+BvnYNoiaX2edf
H+AVHbfv76h2Cr6PBYtSGLNOCFstJ6UkyHXFmVeLLnPcPxYnOkUg8HohrbvXUR71
L2tQI9lToIOfpnaJROPzHr7Y39SgXNhPrgXgXdkhHkMojB0Cny3NiUs98lfe7pQ0
2PlNOl1b2cyegzUPDNsIxNIiqi44l+Qq5ugsIlQNndChVNFdIDr/XIWpX6zkEop4
RL3VtZD41secTeSSCaBSUzmhZDzZgx0L1e+ReqM+zUBdn58dYx/dlhT3EJJIoFNp
Sd2B5sCa7Gz9FjsMZSBPLrJ3nHPGQ2THHlmaZeX56RDlGjjupXMVHulUgKkQzAlG
wZeSkTjcxxMqHlY7IWauCj+s9T+0YQgWzZyNPTBUEpvrApDppOZS5MY92EIvWbap
59YAF4n8T3ZuFeKqQmbden5DyNsyq66QNdmqbVgbiQ0MNLOcdMnxawpmsjioNYVw
uSEEamXb1H46X6CH517wd6gzG9n+/hMrXGiPeBoYHBpj8CNfnsMvUHKlCkVvmiUz
vRs6IRkj2pxSzdVapILar54Q7T6HqCgYQWYe22mfCyI1TRDigTool+72gWpn8acM
P3ic8/K2uSo2EyiqhNEE9Loo0R9pFKF7kIJKtSmq27sCPBbe5U5xHU2Diii6h+aa
HwVR0qj5z/DgiaOGseM0HaQq5VtXRoTYM/4W/MZuiu2jQpkHXs+lhnA92zxnBjLO
+iaH3fE7lJW5jjJW7N+TbPK3ofc1b3R5RcPbWmEkN2DCPXi5wrq0M2fAN962VoYY
A1sUxraS41WksOuHaKOC27KEVzyj03zHM9gAO4P7a9jn/UZ1Z91Js71J12ajtRor
Do/UQqvxXglNUO5cGZcExkKXY+zXVNbQSmNsl4F5iNdPjMa8sF1u5fjTq6TPieph
xo3Zc+1aV4vOe55Xh/kBRpd4CpcxmzjAy1hunnaR3Oy9jJIvj8VqYYz3jc+4zhIs
mb82lofqjeGblv4cOi0cU5jVQiXZyBsw4hoa607DnW7Ah5gMwHHHpfdUsxEKbvzj
tD+d67J4eR6DfCQnYMixY+Grsx1ttd/6u4dk1qfNqw0KBRYjhrrc3uodfIpJjvG9
eOa4bvEuBDtBYCHgFgTzhKsPrVVdkAhohSUieWQM0hDiEbVv7Kx5nsXD0Ep9iGTM
UVkvjUsVNXwuhOl27PKbTfQEU095Q6VHVRspdA4lc/tyNUFPr05GU5M8V92TdEVO
FsX676wWPYl6jIinJm5JD545RUJ+R4A+HYUuVsRzDrOp1O9l9qkNNf3KQyaEpwaf
TwSh47aCMjTKn6Ejo/5hxj4pLitIs6ciYE746BXG/0Mrdm829j6FHdMVGMYvtFON
1ME6YJvfo4YRbdF2a0ygByNQznC4sdCYb6tqiNXrVGSEAqzY1CXkbRxyHGdtJNfI
zQxXF6YegqRnzlXYahbCqPpr7szpYHXUJxbQQa3gGnj+kg9iCdqp8/35r0XWi/vZ
cDrE7d4GKLql5CEVuHauQryAf2gldXai0SKhTtEL843QHwJbqWJLTzFrW/2XfIAf
KNp9fiQvCbZuo1/YdoAebH7CYzniAVe4yECeymOn8ImIolP+AdKUMXVHpVmPe20W
9M3HUUXvWxIpxCbIHywQjhGXktn1AUWjR4lgveRTPbRHDjJkEkThQnhjzahTE2be
NXoBeUVtrFTOicbalnJPXAXYOdcM6qLBThzpYbAE1pCi5HnPmmLEB8MP5MAmpvQw
2FXp1DacaD+S/6wBbNPKlE0YcHkk9t/ya+lqs2Rbiuaa0RkSsxDjR6YWynk27Mu/
SCiiNaXhPDTetFdzI7j6daP6afGceBwQYZ9gC/f54WGSp8q2fngx+idxsC6nRCD3
yYpKQf6jirpg/LHtzXCBmIZOZ6+qxY6yFNdF3nOWaO+UeTCUvsbtuB4Jtuqz4xpa
KHyabTmXSz0X5/PEoU1zhbiNutoGLUd2GPO0BxikBV80Ol+81HDepdsIrIug8+nt
aASrHM04kWu1/ejc+Hh+Y4nusV9Q0SW8gnp7GolRKvj5/YeOwsFtuC/wP720yh6X
qvtDK/6n5QG0h9mLMmfHwvEtnv4syOk1BZYH/3B6S57xdITlHHzoxCby9KzkCh7n
9antB/fnDN6KV20e1Q9HOCy/MFe8oR8w+Y+37Pvz1maDVN39GrJDqK8NiR18ygS2
pLAMjbR/Xp42uB8BjrrVjm4RakJERDNDW4qDJsTtd1+8usdySD5F9joVDRFABATj
ZY6gjDSOEocIgXfatebhsoYkO0S7oiZuztigKAkdVwxEj5o0OaIUEy1LxqdbLrqC
FGPsSI0bsEWOi2lEaC7QDk8N3dx6f+Q9gJDysVpIYn7yWIs9qtEfL2o0Rd+aJxv2
VG9YAxvINPsbPdowfqhNwMZUE7Z0XdDQv5sbs0WCrKSKeEbtPK8WUHdQVR6avqfl
chtZ6yho0XEsKrPX6e7+9kG2Eas2sbu3k/AiYO+jO00NNSDqilPy/cKeCQMVN6xH
RUrdLkIuu/7E28E/9XU40dLVlbbmGQ9aboVIs8152AIk0JQN2Z5Ghk8MzkTTj45z
mgOdwC+3nlvFJC1aquBnX6m3oJGjzoDCCyC/Sr/nSiprTuzhaDFFB+/XW+7+J2EH
hMrjznH0hP+zMFsufqDD5IYF5aQIRCDJOYbhll08ucb2ajmQDkM6/2B8e64Pyy84
URwWWtxYdof22ngcPXfwgjtNt/RnE7//YIFnhvKiB///2d3NZzxDOhyVZInBarey
L+bfj1eST75GK23HYHlr/eJVL1//c4MIUqOHyGSkYVtml/v9zUE5hKG+JePTXwlB
FN0sO0KbjGTGBxCJbumDB187jsZMuAGfeE0mzA8iN2mVLEqF6M1nafNDGApc5vKC
eigve2OjfXfvpufGw21jhW26PU84joLPPrIsBq4kYMMmB+IyGMsfhuFcAjUhlF39
KBcdUty9yDv39Tq9QUS54zPNRUnPHF9gMYvtmGOFGqcLhHMGmWYECEPoc8oOsNpR
WcgyMon83dW+OF5s5fkQFR5AfTgSCYmHBlbJHyWrBFskIY9m4ti0q6/8RE/kkSQq
hfxXK9oH9JUuxEQpOr1hADb8hO6pZvvPygHrvdOiOYj3hSEuFRcHAdwpZdmuRBxE
Mr+rJDzX0s6D7zttAFy7gb92Kqp8EBfT75Cs61JViIATwnEeWiJkE4ttpCaXfisJ
x/T+eMx2CNAOt+Yy7/NOXhCPQll1HvpJt5OIyzP8EWts7f0KziJI0JHpRwnz3W85
dzNE7kpgK2YQNQlCFK88oWaW/rKQJh5A4edp+mayZuyPNsKIb3hh+3QtLKqKBI0Q
IJhlR4p4b/R3g5rQZeRLSatk3vieS/LmU50zt4H4msUG+v0Mc+XGp74yFQ1Sc1MC
xJEc+HjOeh0XVLIMAX2HdD7fENV9nvPr+GXY7QgpT4iTLWXMNocjADuoe24kR8Fs
oZEoNTY3ud9uxRe2PDh7mEd5FozkOqSVbsuum7gEagBF32i+EUdZsLiD1Ux6Hh+P
2YlGYaojCOnEyDqHzaRKOlPgOSxnZxvbg22WbieB0xDso9Enscagez5lOUD+TOdt
uh2M6YNtPuOZKQlXLoTPVoYLET50hwykRlQ4MSAYbJmY8eXqaoP1BmI04V4rtqOt
wi2d8fBZRBtiWUkBVM2ZgXH46+BN5RsOrN9iO8go+2qHZSRHeX9jkYuzWp6NRsuJ
F+dQgjbDSv/NMd21xatSbGcEbYFVgTnZLY4jMd/iFluoWdTEyvg3llFUes3dJzQM
g32Ccty1aO5m+MRbjBdGdBLRpZDVpTjHHzmDA16iPoovJAmqQI4sX/n8TCykaM5L
9A0l4KXMs+P7j4lfMugSr4lFscr79NhHZmGh5U8MHJ3zXP7K356EL8xdxcw35lxk
wng5pl2n0xbrJ83ATABwczRfhZ8I+6Z6HzUaJvUfM453KYeYqp78cirbyUOEESKp
hg6+DDXynjCGUQ+sK4xtDuAsBxTBWy759w52YZkkpUwnCsYlCGH9COFyZ6i2lBNI
yQECjCN9dQat90KZDk+87gBjtIDGcP7VYvyIS8B6o7WQG6NthWscsNyU70RIrwUp
nnf9UyooItlLwfBxPu5ofUg4iZf7FAILH/GvDr9146HqiHlpjUZOlooX34tlaHDs
VEe2AKIiLwa+9q257d9uqsybNPgPm8o4HB6/FUWwiif/paBCqVYGmLJOsiRs3ppA
q9Ee+Vs2WwIpOcQyyEpji6k1zRQ1p8oiuj52ZkDJB9pXhyGhU9JA0eVKtUI56ypU
LuBdzwlGtGYEF4PBT18/u4qhacF2ah6YJ2rWDOTnOmJvdqwRQerABD+fYjSP3qfZ
XzwnRwUthh1KSO22c8zNnd7591LdKZhgqo0orUdoyH+A4Uk7/o+RLIf7nSNQUx55
f6vDZepQTG/Yf8As+dEHBOnziveYkLyTjdmymKXlgnq08MQj4s3m3nTauuIEkU6W
bV0eyL/AUnNTjk0686GZUL9irwneQJ8WnjTRNZ0jn+PKm2pr4xdPwLd8MVJVgy2m
XUvI8hr4vCmcOF1m5afCM/zo2K9jDgSziy/mXv/PakKTiatdl3PSQ2x6tJviVI1b
e/y3wKmMhJQ9v5PO7BvcmA2RRz/IvYMZJNXQ3GnyXor2S8Prm9Zqja4DhgscGTLi
fSnREqMTmSPiq8ynH14usAIGjC1Lb3IVvmREuSdQo3uzoUmJEclyqmV4ka3hmhO5
wAaLPepRUk3oXidCs9dwoM72QsAv3CB7UrWRls/a6ZopriWNdrRmCNtUyKHRwzRf
3lps0VegS1QXfC75ze5NC9/NJ7Qtt/oOmwN8i7PdqDegeXruslEFUcfHX751AlCC
iFDprUsD50HjMk1eiiJDm29tW6aj0l8oOzKFL7yEFDD8aSoPv5z8FN2YtRfNiA/y
bnMJwPVMUktXAPfwHOd+wTZOEAZ5t+Fvm/vcUHs+fSQvlj4IcKC2jhDrdrx7MNty
uoEsTEBSMk05qmMhpL5I0MxVb3rl/WYH2Z9I3DCvOQm4zZOz88Me7KdBP27c2LCY
2ZQjhC+Rf4vWWoIWw3RHkvTDQUVT8uQ70S3ddvsBeW+liFovBFeeZRcKpPWcy6DL
hyC3eQfKJ/zh1QZwmVguUt1mDjRLRIG7mw3J2cMEXopOinsaxLq5eGLgLMFGP5Bn
mHQ40eRHfV1dsKLLaRQq0h4XZ+v6jqXKBrVRCb+NmJihhlBxcZz0GmBtua9mWjPB
bztkpBMpknqKHUnSGrj378mEbYUFMjZUAn3cMmKthWzUS3ZwHeij9K2kxN4ODG7Q
vpOUigGcec6sKzYRCzYPFTW7rywNwEN+XmxrhXM8QYT+BKTKanyWP6tYbOrVpLy9
vDHSpXvUkTDwjgYQaM/363HZoRKiWrIEH49R4r/32cdZ4U+B/0eNFPJX4OL44S5Z
Erv5Li2wWo4xw1atwTV2CSqNB+GUjFWhaiaj/fUla9Jek7lPqguTQhYEwttSDGoY
qXCP6iK2p3Ki1+jlpGZ+sgP1oubCQImlMLmMO9lgcaYt60mpPmtm3337dPKh2xw5
PC0cZA0pzDliJjrhM2+1mzH9rTc1c22cD30lCmgouOcqUmqeg/+kDridSzEjyyuN
CGK54/wWnZtHqNWHG3GcTq3od49vXG/96vtE2DVMuIULNSFn1JoMVfXb32/3O+i0
4TWK418qZFegKyTPBZh/qWn1OzZbAloHVTXhBowM/7HEjBV1MGKLdQvF2WJiG1WU
erso/g+676M0urdsq1B4ZF9mYv10R+mQ997M/OVYs6d7d8EnKujFZE6CCfe15IIU
exJGyuYlVaflKnMCVFTm7q8ClJ9CjLKEphNVUGNH++grDMJo6bynD5svN2w4A1bM
CxLWddRNiATkERl8uBnCKdp/7TyStZPbRpWDKN4JvIm3bIBF4qjmODbppxP8qj8w
w9oNvogPet1MVugtopShEvaUBCyCKVBp9lW53dU8e0PswIxGGAEXiwVByGOi60ZU
sbMIWwMnmqaLQPkmddZQNc1jALXhvn/M/VyU+BFrF8gMwXoG03Dog9rItTBgXtFM
zAXH3dqFCi35lXt/T/l5t99lHwVb0IQ44TfIn2Ptl/DU4Gh9i7soeu3YTl8YshC0
Vxpqn5jNdZfwtUx5WM+OHf2+XHMon8l1LZS0I1HaG3UE4XteUGvrZd8f29Lqfn2H
SrB8TDKh1JbWRk0ucFk7XbjqDcpZM3YFVfGMO4ipl3U/yGxv+o6PggO2gjkzJG+A
oze4FUvnfy7oAzYb2jpfLCQG++iCfDOuUUrGduKvQdIL6YuPCHjjw7Frs9avxF4N
O+r0LCI1cHF8M7iCFGUlGiZRuQQNc5WXEhmf1M4SqUjhMcOwlDkrpF96L461nt4h
+6KP+j0A0DmADS4wnMplZvzJ8Kg10ybMGWUr1AIYb69dnxSe0VHbm2qvbDxxZdTF
WfMNFapEw4fACdGYgXR9nKETEzjr9bWt+8kNAZVdYR9oaq2cXwEcL0MVzRPQZ3+s
alo4rkV0VxuRCs6eYvX+BOtMwUNOkp7+6QPou2d0Ey12zmfS6FbKyW2c805zuYTH
HYmzYp8LHkTyG3H5zTgQ9k2Km17F66/28xCw9+TDPweA2hvJ84ffK9pzqsOsf9Ow
rsXzZNPJ5GxizG1j0LBnvVG69gYETDrBqEGNhCkB6dvISZPOmpIanFJXf0FtXWTE
JlQ7CeSWhqfbHPTkDPYiO/0848kwnPc1rOw0znQMCyhjGFWvq183YvaxzDE7PH0r
F/Mq2vGeS231n605YdEfAr/Y1eyqr3VoMZnFNWpsdFy3Q1Y0ktzBuRgvSWIXLsCc
5Wbmqstr4fpyDnqJGXxYMgLsxEdpFi9lytl7PNwa5CfcUQ5RcZk4Q6dDO4L5ExOv
8pIjBFNKuX+ynmo8W+CyKDLoBYttBrFSi6aeLJWXa2o5zKNFAep72Wlq+IIg70u+
FwaKn34kf95Osuffd2JFq1KgIcj1j7AP10smfCUGT21Mo+XxPTy0SmM5f0yMNWzY
XHmIogJ9/Oo9hBtFtp3BteW3u6UzcrSMXuPFdyRDSaB5sII7acCD7gYjeiNtOJ6j
Hj6BIbhIotA4yRC053Q1Qbec8+PFvpzIKpc5TUaEh1itV9xH3FmLgXlR6cmgR2V0
BiRjkPNM6PSLYXhnDKA8dzApblLRkTRimpgr8yKVSaO5/5JKk5ky9qsTCmgmoIN6
ap51Rkchegz5brc8TvcRs/BAxwA52havJPCk/CfnIu1lXEeoMoZ3OgideEPYp+2T
DL0FUZgxDYpNZmMpN/7aY/yyoDmOwY9gRmMpzgRmzpaRt+2orkyl6CM5OJJ8w6Z5
qNyMl0VtRox3WSO1nXUCT5s5T2ifxwYa/+iwQWeo+6RMVAkztY+pSs5vg6h2m2Ow
9btddp97xMTrZzRWxqcYGWGZ1Qvs8lLk7qF+HzTosN6+JgRzkxApbLP6nB4lHzKw
MqAUWBrDBeHkpsNVLN7HuANG3d77ngDlXrs7nMcRtwRuL5Z5faKa61pzyWMHycIT
G8GnFXoVy1ibkiGz+C2nRBdER6cMTxrZ8mXhYZK6s9+Pyv226rJWoN/uSxa0EXek
UXrNh3znKs3HCrm+E+GOwaq8sPTlblYafySenS0CNxqQgMxTFvsV1YLvb96om67u
lT/tvedu2eH/IABY7oXHvcsxg6uZmrJsxjRrVKJlzWGIEHzm4LtUT4HY5ezWEbp9
6aMffZRDDmnA9TSx7tmQfEgijhYvfNPMDXfTwR80mpHRmQtYgTlj0ckcevcttswW
UquaGrYaYr4kfEAtiJdoeFGpD9zYPKHEN+6rZtiCKYNAdKUng0pRjtD9mUfdP288
rYnPILgvof4gJqbUvkXGUnS9o3umiOMbSrnbW6S55a8699qO2/tprL/0eiGch6jm
Y2sPkjOdSZ/pGSiQCLC8rZsEpagRl0ofZkExr1JVpoIkVIzSg4NzZ4Sp7CaSPZhc
jBXDzmAUV8tr3Jnd+YW6d6yUYTvhFrl9M/HQ7HaEuWO0Hv1p7t/PH6GiqTNU7/bq
tm5d2SIohbAtmL5E02y79Ll2xPucvMqjElbx0X+5xquJXXicJXAVhaCVlgNCLbtU
c+VlyvjZsrnlzEfmyUclHCi2wyZP1jlap7V7RLR3u0qmWnyzZo8mZumgy6/vGSCY
bXwdBn0MCvJn4Esywg3GlyEkDtQe62dBvumLzv/GxmNN0SwTCCGMk7pMiWMSrUA0
IuB3sdtl3lyiLlaNUiO4g+Vbltrs987pcWnH6/1AZcyAPhMNomm3Ioc7kp6tKxA0
kGR/E7Ld/uHEu6bDZY6K1BWmUUzIRh8KfTahV6fO/7nI2DFyFMvxPPo9yXKv9Ur8
g2C9B5VAwAww+fBnJ3UHa24ia01tXRQlZKa1lseG2nbTAOZ4h29YbLktbIcbvhAT
+0SwTOZ3ASNpDbjlGUluIUxjevP14//uq5e4WjI67LKuEin0hLbqNbwVb7ZF3W5q
bbwe9xVIdODLQlSE66ZEGIHWWl8YQKIpkRDZGFCQHSLwLGp2rqiHufA9LIvNBFG2
BY/Z7rr44x/jLbCmXSnpI6eHjMXIVyRB+mgDi5Q4DbBlFQP+XnrAuscS2VxKBbBj
`protect END_PROTECTED
