`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xA9i91xUxvOfEyoeVWbwzN6UWzu0l7GBpKnLJLSo7yq1/13S7AOzoB+qodAnrIGG
dvsO8JZVGgWsuULI0eumcm1su5XP+VvCz8Km/c0SLnSxqF2/F6EQgAdQeAd1TpmS
OC2zczNjU8xVH9MSfiVnB+LOMZjvCHqkoQHnV3cLZsFGSkbzbvEGjxPFGZFEbPHI
aDttFo80Y8ga4E2Pdvaf17ItOOZRC18/WcPcMuNXiijigDf3eMPbIDzxTVHGxlrT
NG68AWd24iHkxAiP7tDtx+vF1B/dUnNJG27gy6DkDYkOqIUrZwIEQXUJUzzpTuh/
ZDvzwIb4uhWwj6SYncR8lCWP1sRCyCQvakRJwauj5lT64DVvXe/+4DdS/ecav9aX
+OtQiCphQuhaHcJyvw7LMGwcdRpz0yLyBuf660t+ROecBY2CebFloI0WuORN3V7p
`protect END_PROTECTED
