`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jX5pvWAdmEh246Nxj8Kxg0FcWsoyWUN+alvsjYzQLWhSEDQMr3Gyi2DoDiK11+Pg
23UW1wXi1d602xuVrqVV6o9s1IJmhhuadrao/MEN/M81cfI2NBlgY92Wi+z4A+ny
KCMCr+d1hqagEJAqZHK4VPlMa4k7tSYoFKGz4eavB2Y/ixFy20msWMzJPN/yzuAM
4WehDyeW+rdXXugFRSWruObzPsc2mjsmV9ivK2jUYDcYKtydQi/N7JzM2aY6G4yM
kt1SQlxs0BwwxF6gwx0wQFk9fVNTwqD45BMlBQNS+OkUB30lWxgf679pBOdfTywH
YLQBaRoh1QpA0tk99N2ESA==
`protect END_PROTECTED
