`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4Q5jdTiewMZb2RkGbr9z6ZLWrcxcw/Yx8RYSELiyZzw9miJcWNHyTztjd/mDCr0E
MDpdl9ESZvLkwi0dt8pD6XympMfcjwwAl/zT8SAaPSE+N88gDBc7H8B/VVMgOpA+
LnzUXORZEG3jFKejtyYOOOw6J4aiSSCWFaIbcXY3vZZWtYjfVmiQ8DCeBPxbza51
mxTqwLBbAXlPThnMzklbQgAf4fYvV7eu8q81nPbR8v8qIREZ4mez1slxKg1BDkeR
xdpdflVtYGdYX3UCZk1MuJQTz50vHaROUikDP8TFeOtQ5Tz3nfgDIMM/3hqLCKDn
kyx9DHDmq2hpsmpq0DutcPt9RxJu/vBqNq9C2Ea45H4=
`protect END_PROTECTED
