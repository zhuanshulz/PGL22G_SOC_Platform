`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SZXNoXzJwjHp98cm9vfoFQ2jqZUd8EWulS8IpRjVhRig765sEWNq+sgpo6Xbj63h
iqjXIrG36CRBtX2c3hJlBgOGO1v/IlAzMdJ9sUIVbkYx1CJjE6OWbwz8CyMQEwUs
usR7ikbG9RI4ddsww7uteXh1oWQ/uSnO4WT5jwLOXQiO3yOcpt1y4ke88Hb5gVr3
hEtQXd0v7QgR3ISt9XQIFuxpNXC3TSxJ9P0kCFIZ62xNUpl8M3TE/ER9YN7ZC3FQ
Q8dvm59sgRd+stkOToQub546s+CtfprehHVT3xlME+8km6WTan5P+XFdF4zARZKS
fqDKrwmmTdRmuCutsOIJf7xdlY+HRbjuaedftPazTVVODQYycVq1v8qGcRq7wvdC
xgEk50EuGcpv96HMIxxvZfpfW3XqctZzG/Nv7PHiuyAKeKH8+l0QkUNZZ2xaVB+b
8kp/s7YIZ0WS/iGDUR9wMA==
`protect END_PROTECTED
