`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PdlnyWCTADDl2B5KbBJGW68H0CApBrsiQDRIrMCbsLpounQmn2lMd1ZLpcw7/K2F
fgBOAn0wVYKvgm2AjBv6zb5L6kiQrxvNrFXyIhY72DUxudKqi0cYVxcV1QhupteY
QMFvz2o9sdseOYFnFzcBpbz0c0eVV99TyyOaLMXuFnVNXP0kfB05fMlY8ofbDErO
xxSFfNH8E369fnr5gUOXt9A4xgDsH/dDVfnbS0LFYoARSlm2AhsLTcaW2kj6R5q5
ZMPoSy7066pAyvVSAD0zZwWUcguaAZnylPtQVkSofAkYuJxsufaoJIL08AyhdiXM
alTmqsgln0mMPLt3fxhFY4ZvnHRRsP7HcF+EI/z11VP+QDBbr8xwN32oNNwb8Vx+
2IxUD20pOqBOAdv6BYL0y2LWwTmOxy66LadpMeWPo8rGN4+m6KWXmqhUSnaHHFwy
EoeAP1ceNKOXx/ususuJr7T4lg1lL4s9t4yAxtEzVQuXCI4Q/Tnh9jWPvjs5W4ME
tRXFqRncwt9nN7axLJf3rYN4CDqMzXtPVLACLNagKeyH2IvbNXIz3b3EW9UwgZOm
zDpuADQ1OJmaC4qm8kZ+o32n4UvrC8Eep5QhhrIpq8DNnCakoIOj27HJ4vWeRdaw
MrLnBbZYBs4lK4S73fJ5T6P8wR43bjxWswd8f0idzGS9jC+pnnjDWck7RpZgkWTV
eAoJg6AXiGdrr/FMIBC9oP12RQG7LYAu9Zk5IgLLT22WnTKBr/PP0yWkJruk8Cxb
`protect END_PROTECTED
