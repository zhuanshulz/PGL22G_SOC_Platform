`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z/LSmb1jRdn9rQMXckqpSD9kIf+KN6brpLELyX+2qVihd3dD1FCvPM9Kpy/C3cIz
xNgGVAHL1IAlOR3VR+RFcx/nxCLT0WuqLclLz7KBWl5VVwbv6fkl/JBu4vRkpdai
WHRqndhXBnQQvNTI+2rjo1ooSz2jNmhT7j8qBXZfhAT336WrJJqv1hMMNtgNZRO2
oZOjkMp1ReaEOKdfcBiACTQdOBYmca5Y9rmENe8aM30ugiPH3KDzlHGUsQC1GwaS
77B13nSyvT+5WFwxIDhhlC57dSc8/cwUIoVXJ4h39gjEJJhV16jg+HTYSqA7wdkF
dRQRlNwPzgtE481h26u8P+uiIwwE1jfddpzmDzeHoPKYI1yN5fnwKAVnNg2TULt3
FjFfhwsil6tOv+qMqYvllhTSE3fpy6IUFFJkZyDRSHqLpkRLjJtZsZ81JwEorvji
rIG9siPMfCY764muotfsYYhlB5dBd8z+6LsIQMeKMZtxWgc8VWsngjxazrSkefIU
uGk8N3jdd6l39R1iXf8GaTC23LIJy2VCkWu/qlq0zKb8vqupfT5Q+S5gABX2/R/G
g5FO7Gfm2PLygwLutHg5ct/IJdYatcT4Ly7IFG/GwIcSTSfTMSJmIaC5CrgkAtFg
HAA9GQYykxYcDt0aa4mJUHK30Kqa1KcsfllEdozw0Djn+E6Lw8qGL73hai+rTIkX
OhHGgKG0TAzZosVumBTw6pUFZKc9HyToPt9DZq11W2u3XQWWwh33JrFFO/yIOJ4j
mhmal6/UIWKaNRHFA5za4dMwp3EuyraSkT8tJkZK2eox7PD/xf9D80Vm/MPEdp2k
4ZAsXZ5/j5+Z7YjSZD0QIerhS7uaaI+nXxaaDNSIMvTw0xd2uDWO7C4BP++LgEZE
/WEkl8XyAU34a5h0fzaYZtykVjoqJwtGhC+N6kBzp7CWhncRGSeB/DkgI/ZP6p1f
WsrPoY74q8PiFZqSChuyggWIaagDTzw1cGUdB02cpIxf/ALGIMKntsgqohz78ddw
qTtb5QittvifDXaVjf/hWeyqhtfF1gq224E7grKbQZITNbrFp6PZCjoETiPHso4G
Cxpf0JlIUWdHqrrzzGr32qKQuhB07DiO40QaqP7ZWzIpy42FVCe4aAcIm8DLXwWg
Dws/LkQ6kazomY1XJx+Lbdu6XvI43kq0/9HxBOX8BBNO7XNz5lFPf7ko/aiZTQqd
gZWERtJSHw8l76r9xYtHpqDsnxNjz64tsUQPG72QtFmPvoX4WrRF7/d0n+5J+w/M
+nasRzoulxK123ehH8dqHkZ0T1GLLaaKX3yymv5ZBevBT8B3vZpEzKHf7grYbczd
VDbfhz8uuv4A/+bAfs8+l2UESlviRkVBd7lNlZ70CqBQ0UqrqM0tatwYIVls25fx
B2Pxp/8LCSTV/+DFpcdu0ZskqZ8OOE0wS996Q/rzwshVrv4/yHabQ/oXIbguCyCd
xstO/olY8T0/fthPpPA1hg==
`protect END_PROTECTED
