`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wRFJtMRDblCVBwleGGdsY7xSyitkviud5+aiHbfQ/a/Yd9R4Awl0riMfpiFTbgr5
QGzKd7gG5Pf/w9M+iZBls+lWpLuD6H5P3oBbstFrc4L3AXqmNCzdEkfnYhzuryqr
b9bHl4IJLWYPOdafF+Tgb0UWCCTsOg+sIueY26rnHGe04bSBfgS6oWWBqv8q9qqp
d0QyyemcBHtZmG21DHF7PiKMa0axLHJOqc0aUnU1ZfFR//dm+QbP6nU4BJz4RmO2
RkhLJgQE/UHzWYGPfHRQM05s3K+nvjER2c0NfvLO8XatgKG6ZehdQ97zBK5J4EGd
FvshDnyh5QabjwFbjhQm6N5qBS5UxDQ1qM+bBjyHxhtKxiVhHo+zFvmaEHVqIpBZ
HcU4lVe7fRPKom4hICWhXe12lDcK5sXHdAfmDsU/uMbr+L1WxYPVlR5iKhVxZY7y
OSVh4u2Yw5UFVwCkFoCpgZji2OhAIFA2xM50rB63Z5/Vz8JjFBkiNj8+j8Od2pMv
MGqtNsvzX3SXIz1njLHTRZuO4aXsYMyH5jJUFOykNxXQ4GlDMYD0l/AepzUULMH/
w5C9ZWWOoHCOT9mMNi83RHcVrw1ihZoD0YUE85M8Yis=
`protect END_PROTECTED
