`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9LfcYBgzQIhcdK+LFgA+3NCPiFklGzPEej3AnR13CmZ5s1PBWq5Azu5NRWc0rbLh
XmENrNQ0UydsZGscfKb7NAx3Xw3jpAC7ep6ChyO5Zeruv6R903s3yaVcRlP4jeq2
h3POVrEvIl2A0fctwiW8Xu1c1N1TvakCeayX7tarDXRa4r+1jQvVdqzR2RoXQ6VN
auMfS0P/xl0ZDezzutdDitrakTllpBuwJbQ80lw8TSYMO/IifxmF1JPHtBjYIRGy
GOZD6osaTOsLaLfhYz6b0Q==
`protect END_PROTECTED
