`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IghABYLzC4gqv+CoSvLWKka3hzh5knd901TxddokUTjcl7BcbhNaIdnoVkuMKys0
wpjhINKbA1aOxROrEftDzHD/jtyPetotrUESvIHUnx3URbE9MggkZKEf+9ABC7uH
G3NbY73verKUoMK4skPlmNHrB9wUJLZlMVmrh3VsqoZsVOFgppUrs3NX9VI85vxa
JOeIPsfIB7VE/jv91UVren3hNTrEd8GI0+0NPeWGwgZmBPy39ZfCGQD8bCYKR0TO
/ub/Yumb/MMc/GImh7hFtyluHwd1aVpE97jXWy8+q8SvrD93+51inHx0wpwU3vkO
aD+m3McsgZ/FG/PWR2FJ9BV+P6IRuGY1ffcQQugbHThiGyhxWzFEr24klLRFInvp
`protect END_PROTECTED
