`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kpKnZaAreyWzYmWuLktQAqUFYhpHTdk1vIdBVFIHJINT35oAnO5L4nQ4uMI+YrTa
u/gDsxod3tC/Gtgykk03LlA8UA5+yZ2AB3C1vChFLkWcsarkW3Rxug2tNHlKWZKH
R9nwDrW39wRu/iAuaLfMtc55878PeJ3pD/kGPcqWNTu28rlEfAERe/v9Rm6KJ2XJ
xcfqY+VZUCZ5WtPyS68QzoRpCqP12De/EijjCSpJxkS2DRql1fFSVAa0uwsJKktd
abu07T3sQ3GeouFSgsxJ0y7BZCcVeaDtnz7Dg5MpJa1ik7iA0idDE/joi6BQKIfg
SlASyPagwS/gztrUN7RT0cuiBmCYnm5+caG8pKFoVVz3N3z/vDMxvqOzbWF1IAOv
/q4NEs/4cexMnQcRJqNfrfmaa85hhYUB2CIXeiGfVfGvrjn/51IZ2WWaJeBo+QzW
qJEK/Z3Wxg51grpD7T5JFBQ2KU+LLask6x9K5eMlBOsGaEr0K+Rfn0+GeCz4w31i
GM/VttPTaSlDkr9gL2Vb2ZPJwGczV50ytzMaklyieaJVxnKeI9HGq2IrnPpYaqdI
+qM62NVJ66Bk9/q/grRAbzwbrg7Rk3Yj6gD4wD+SO8ooSY3Jn1+UgrboYqf4zJkR
qDc/wtVhHoev3EY9gn+x04+AqNFLutT4CImfIQGnmaF94v35x/s7MQex+lHI26A6
otRvAywLAR2+HluoFUrwNpiSbmfHISFfMLN5Uimm+RejQIYYXmdePi1LF9qSbLKi
zF2HCUMs/HsPX59wEpoKo6alOBnPXYgRJMf3Rt0xuFsmkK9xzO+Zyn6NWSR6oCuv
tbqArSOBQiei1DWTRMNhyuvHrTDhp7Gs9OnT5T+bggVFdUZKMXozBfm68oA5t5aJ
jpEAbGg9y1XyEcZpPnE3brMpo+0UZg3/gpYwoDj8FIg=
`protect END_PROTECTED
