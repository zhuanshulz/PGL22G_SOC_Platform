`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tk44b78IDY+nS5YlRIs15dpVUqZjbfFgBc64ssqZxlCcBg+8STJpFTWFUHug+RlI
hP0mEwYJ+JYuNNn4GMa9LJdbIUKRYbSBExsDQnR8L7iKjadz3eudM7/l08hZBB+F
10AJR+Q7fE3P538aHLXocuqN6lvXqYQSCGw3MePNqRve+iwUXVUexsWe/5LHJVv8
otxA4MhSuS7uO0ab+G8zyA2vN1SeoMC6lEzpVvacjBY249uRmTFLXZIXjUnxqNJe
VrM6djiZ8Bbv8jfR/c3Jky30ZiNbzxCJO7C5KbY2NhyPf+G5wmIpvNU1N0NCxuha
x+r6yNAmRdP3mNYw0c2n2v9rppKb179AoA5p+vu3oTegVdpHomJqS2uBoSsCEwSS
mYe4i123v6o0sy8g8E1KCYDmAqZXC5bcQdwfk3VGuwgFNH6v1GOTr2Phlx/nl4bB
5jRvS/XzSA24cYEhzVmPhUONGRKcLPJWPegiv/dQSEm2Tvl0RMKdjZl91kk67sT2
Fv6Ua8DkIAN03jmyeEw2v/mxaBofyyaEJPf/snyWPea1MwJIHLqIDNyd5qsVYdT6
dXRcmKp2zsl+SscGMjI0Lg==
`protect END_PROTECTED
