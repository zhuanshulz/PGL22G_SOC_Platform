`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gqtvQ3qJ648Rirab7XJoVA/qpsqnvwke908ljVHbdlcbSTePZ8XCUxPadCy1VKPL
Bl1eYOk0IczMsVuqkqgKKE7IWBfT5hY6fISRd/9PlZFJhuCOvhpwjQXtYyqmWsCc
h6cjICmup38zzD0is3tSu4vBcZn4zxShPSP2jjL3DLg+VRxbZmATpfHcQXNnP27K
Xgk3UURAYt60L6YjIJSigdFueMkZczGjgEBfgvftqwMKDDbc2DQqNr/Aj9BK2jEb
9v7As2Iq9DMRvERt/emmWiP13IRuXPhCQl8jCWSIH6jYrAbCFIxP2qWFcsSwmZE4
xOOA/M5zkZ81TO4Sb7rA7eBmM081RG7X6QfjYqcNTwg0EWfB3p+AjrUka+pB8/y7
d8d0jyhonADCVVmM9oR+l1IM/czB6cda6GvsI003J2qT25u4XTH0K0F6qtJrISm9
MX5L+pPPl6n2saVSLI5/af1PieWjv9T6YCwg4//DVXS39XgDIxo8Yk94yos1fhmn
Xn5+qC6AV66wqLMp8U3Eo15BproNHgfW+6oK9HRLNFELSb3vY4i9sSj1MUQmDD3J
26reGr32jpBAaXFfJo+LQ89w8yVH1M+AQ3Np0UutTaHePYlXFOAFLmwJl59a2kyt
kOlUIcswcznifJD9uISr99s/GoGVDir4hnECvwwxZ0Nig4axh032DWsrbnCPOLoq
+8Qd07jMfOTnqsAgHylC3iYIrxDevqTfdWlem9sb0yqZeIH2Zs7ODd78W8TUelpB
lpGWjbps29Bvw7j32nzZPcjfj0VjlZ8FauhHeo9XPLgmeKXRd2SONQsyEB2wW6Hb
KEGyxhxI43ZjLlBwBcywuBfPGXdZZ7bBg3Ibmx2sdL4c3RLTUKbzJrrPFBCt/OWr
o/WPCP/MsdQFuhTFcwait/chQwd8rD3VY0i4PB+1bKimC3HOEO4XPUZ5LhYVdbpu
NPq/+o9eiZ5lHSsAPxYmVWcjQ7lfGSuDHOdYeSrkysiaofhWa22RbCxrUhkzOHRZ
HEMVPQgmXEA+Sdw3VyczOQOKpatIHE6m95G6rBKWTzWJTQEizkMqQJodlgHUTCXh
jbLdravb5wsep6TOwyan5ad7jviqoFiKD40kpMPyaZKDUFrg7Yj+v863uJM5EaTr
VK8BZTCN5L03VvB82M9P+VA4R0BwyXIILT/8S9bu2EBZ5t896WAOB5uxLJq4V32f
agw5WMCFXLgRKt3cUUx09gbQIlxEVCE4w9WE+ztwpf6ykNOLYBtvbXHt0+6Y5OcR
dS5084KGPu4apsf1m6SyMQ==
`protect END_PROTECTED
