`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0sWwaHsYDEAahgSP+yCakU8nYu0mig3qEFfBk6+xj15F6EaT65uyeUoyg+OT/rwJ
clT11KO87nqGo6kx1KtK6KflOiwdqMO/+IYr5VJwBssGFP5pmilCx/22mwhffX+5
73OfN2+c5Dt/TODohiJ5xELZxMIDTbevZwLEWXEaZj4ssy38wJLbNeD5J5iA2F5i
yoeQo5ioZLGU8275gF7B07fKHXHqmYigyVzbDBLAquhNZvocMpwJzvJdjGUzGc2d
cQ/bjCEFY1lAtGurENyZa2XLHjRe3ckAXaO7VK/UvtP7LQQJsjyw20wItIsO9cO3
4w3z//1XRbBQU+4BLNC0qUdwpV9PO3YcE5HjtdkL4Yq/3fyVcP7iJ/kMqErhzm6L
VAikARXZKknw3AZop+ohJfkyQCwMAlQB7RD6KZZIZ7wIPorP6RPYIMIGTT3a5N8/
IP5ZASiCWsQr6qn3wfLA5w0xrTmxtj+E+MPrddVpPE6jHOn2RZBhWakNPSjZdyER
ekpAN5THZ5fNmJrUvlO7ukLonECm8QKJ0w6VHl9Z75hcoHzbK8nGmpSlCoxzbNdF
OxuvYt3NOORfxv3EHdaF8RZY7j1tghj/o/GhM1drzdYTL058c9MyC8jDg91OumbX
8Eop1C3SJUgdr6nF5kjTr6KJkPDTu/rGYEOXDmLpSty73LGU1ug5dO5yQTKlQGJA
9vT3Cx7UBunoQZb5YyTcZTTi3L5mJ6fveQfxS31W/cPxTT/0ZBeUj/yrxSseQPmu
2Rr1ME/Re1NOv0YslD0ZFNwNzXOkbdhantetge84TSu8Wp7GhLr2ldLHrK3UZ1ih
m1ZBl0Jms2p0QqE/K0evBNgUI76Qf8VCXETlThun0ujwyxZQTwz7IuEz2ZXMMrjH
z4fCeFUVln2G2XWdDUy1KJY87cJRXZGCHKG5e1Q6qs2+G+aYC5ZY1cG8a2IYh1c7
wmu9ianurSiofCnmDl9yHlMHR9NTsd1GylDbEF7U9vVmq1PwZf2IPVy302zcwzNx
yfIy0D0gXbr/7xRa5slr4Iy2VyCoY1XQGuSXOO5tcGMKhf/gtnRVKJsuTytIg+7u
lOs6YAkYLHBC+ZR7jLdyeFRS2Am2lFbn0cn/Q4c6MUYhCe5PCwhFIZLGghdFpwAH
FXjEmZnn9dN59/LEO8yB6AU8gF41fGjTUUUIypbtVE6jUSUZMgkkQ6b0FxA/vrLS
JHftNSFbUOcjpIuoaANxQ9om2c3w/uaTSjfSC92/dN7Lzty9F9A2oviD8fC8ktLJ
Y6eKhXLjVcLnxRlLvQ7UHC39/7jeSYBFJrxtfnUTIu/n5CTBNyeYijT+jxA+sX85
3ooEqB6rNleabR5BcBqM41WQUltRZEpXcuO09+MwAieKOWgjOrJgHa5h/tWzdYLP
hZ0Et2c/EaL7K7e06Klwldp+mlxDEQVuDvM7Dxt1i7W88Lx9cfcWoIqGgoVTx1GL
sSB0gucR1DTmLjsNItfUPVCsMmII8UMxS7OUmA14mz44jFNgnC+IvD6LVwWEja29
WJLUwlHP74X1ftDHWyPo7HcFMURLSIyxY+cf/jLphEqEpXXNPW3MUrr3YV30Z/Jx
9AY9t6J0gAZlToM06mQNyQ1jw3/D97ModKXZxBtKJhg=
`protect END_PROTECTED
