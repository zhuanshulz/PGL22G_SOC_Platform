`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vsq8mrdtwapPIKU1CulVvzYEhf5eYayJmNEyqp+wwQW2ZF/7SaxYFrhw3tF2rZL6
rjVYFg8QzMIfjXThbiIgaEBgUPg5gykPnV22vuxeIqdwcX/oa9Ufk3CtvuJTzwbT
mJbplNpUs2M0U0OStJzx99SkyS4jPCSwrS/vH1D4RCTr1g14SG+UxPJ57hUADToT
NaEIS6hVqzpm6QrLvzBzr0UBad+NIwC6dNkhA/51mZ1dEqt3hiStHbajCjh658K3
1HNpNJYMT0mk2v2an7sMLeFHQKcR6lfmY8M65ufClWkk6kXA5YSqo2K7UMjIqqZa
sSXCV49A3wIeg6zaSrtv+x4z4+uD3YsmsrO4eSGQAWDHIxKlJdXznA2g/dDf2Izg
73HLTi6uaT55/70MT42N7nqEO+lvug7Ijbewojq7mh+nmZdz2GClf5cksAqkubrz
J9eJxVaPldW7n9wZ1fdxtFm1EskIbqcMq0xaygXVUn1PgAGk6k8tA75/Gx68rKkc
625Afb2LI7pyuwCkixgqQLPWNJ4tQsq6L+XIpAOztNeYPqVfNd/1GnbteWZBUhAa
aEPE0F5deDAlcfHklztO/ZBWLdI69kGumEj7wyEK2M3WXvs316jnFZYn2VVg2GXG
`protect END_PROTECTED
