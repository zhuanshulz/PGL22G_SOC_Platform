`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rwliG8RDidhOxrG3xi9/4SdOw2iIOS0xUNgQCmaehcgdxAnhochxYC0HiGbDtG/Q
668Nvu1/ah3o4y6YGvfRLXlglHSqd5rz6Y3iJ0Az4tW2/My4ZEiF+YTsIj2GLBxi
PvGzJTGfxXa3sAYUkDkMCiugx7O3wTvVU5jWSqzTvl+ls3an0JgaNyDMgJewO54P
l4jci43kJX94Xh60zbu2B5XEK/i/vhvk4siRKSMmuJA7vdVZjCIFFPHEn2SbFwzd
8JJ3fbGp0WZIF1fTVnrEyFbK4mt6LE58fQw+nTEsUK28Kwy1mifLhIonwqydfW8u
78BXoZySJGrFTmYAwuhVeL7MSeBSS0+qXrrkUHYYegJB/AtC/OtHyG3OdG8HOKPn
MW0FfEoDfkqkvlBeMSY6K2bVU2a4C/Md9OYTKP0QfB2TuiTOxt5AY5sIiIWgCVsw
z0wx24IQdHDLORQkA/WKBrlUA/Sda4W/yLstNFm8GrFlUh71TQygeEG3NTASakqP
dy4z4uo1+nyqCrbTRye/Y6bOQKzsCI/eIEnVatluU+k97TococUJyzLe4nlxzOvN
9AVlD3mfLl5WGcCGe2P1JJmVfmGoPADczb3Pl2k8kZTkH4hCuRuTuf2T10H07Bdw
1E0xbBxvOEqy3NR/2UWNiR99v/MgigkWI9Ai7lHDDtWuYBv5xamkw3t1j/cz6V+P
kord+FzWLi53Ax5Zc3Fut0Pcg7afWLHbRdSZ0tXqjQ7eRjR8tvdleYSwmUsJ9qWg
YUent6vEWvo1+imSNC8e7XtF6/Vct7I5et4TVqMvNDai2M4mW3AkelczpfIopb+2
WBL6qfViAuGLMTjNXOs7wpTTmFRCC7fgBDOEsa0Eqg9NATDsVQEJXiCl2bjNl2vM
gEfIniCtEdjAhpMtoa70goRXW7Xu4ocd0MpmFIMAhWvUegDEmMkM8ePy5uOg5PsY
2+OGc1splG42/G1PZMWvts4btS4FW3bSa3baHeX+UBdzzSNhuUNWCH1GvCVML7h5
axM9FWbXFSfOdT39vxlggIBZuppqKzFAIwfGekECKl/JBxs7JFdVISWed4+PY9M8
ggs0MEh3I9wHTvey+PN2r58blrcB9RHNFfOzLo/FTEDnPAFXLJVKxvBN2yMGAyOf
qqonegNj9RSDDsFJ6TU3yV5O3eDqNvrYKgtOW7GnmRd8VR/bki7n9TzXWPUvUzhs
j7YEdh0/jhMDleowTBZ2i9kUEAfo534J2X+A956FhkjXwlkefoR9TG1KteP+0s2D
KHUx3dzTP2czYV6TiJE1sSVyYs5YWh+8DyOxIOglqqNppBdXvhSvSXGEdyVV7hOz
5ijYxPJpwomz8dot1/bXCRYs9MpT5vQ4d6JqtOp2EQUMGTpW4DQDi5FobDNsdwfR
/K1K8x35uKg1UvoMqIz2iHUjY49X8K6LY3Yv9kLcf5UImLnhLlRlcJvyNG8Sur91
DIYUWiDjJpgSpvGDK94q3Wh9hH1FfhZt/Wnn/UyKiGngHxMOT6arPh+wpwQoz7R/
dhJUlzPDd8CN46ioxkzqpwmhkPGhsp0JHjCcwrSaDT8OMjXFU7Fel9lDGVcp/5q2
L6TPblZcD8MAvC7SljZVAh/H4tsrEM8GeJ9OF5SdS9QOjtSK5FvT/W4a7UWiw9eG
W2XaK9QS/w3E+/RlhY3kJNw1yDZn4bPR5HwrLSaBGc49DyDwfPCVID0lyjm25WgA
qOlcDXzqk9/pS15vTCJeuww0UwieQMG7UHmQ9SQAaHK4D/0gN+qpJqLjm+oCKQS+
QRdnYIGfM4aMi/oXXvcCNah5J66YoKjBlw83+F2I0lH0rq9/mZALZwVyNpSnLSla
5hDkjIRf/UcVEhv3okPNjQ9Czgp7dPU399d0ty/g+/E8YtjyFJh9B/J5bmCZoZRu
8t/IEbBx8Kn5mseLPCGvGw==
`protect END_PROTECTED
