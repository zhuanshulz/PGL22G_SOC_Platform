`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JepcqBtEDVlEZhaQzT8gbPwQ9rzXADLxoLvndwvndMBlhjmtSmg2JJ+QNSWNzjKA
DPuW35iheF3xCyjSIkfd/DLpgLYZd7yUhqcqS8lMjis2BZDO0XIW7x4xJMzh26C2
+2iVelfMihmjVR1X6evbFaAVuZ1cnhGMgQvbMTOx65YHF5oo0EoCT+BPGErqAxRX
0UVNMDtObkZB6fj1qu2NxGx8ew6o0rmOCzXUAwHVm977k1UYZ6ERJHPO02yH6P1U
9tCVRWhcxIOtfvPTVlx8O6/HjqCHcKqCJdZKDLA7j4TufPPw1nhX8qg1IQvvTD9M
Qhiwvevocf1o9W7biBv2R41yVPIl6elAj9pRX0TjqcfJyIZeQwjBMMnGNRIp1up1
A06zDep+OE33wleWGvVHUm69oIaTzm4T3iJpkBWZAGyAM/EpewPBKd4CaYg8yyya
DTwNNsXrEnEnKp+9sr+p3Ymv5kzWSO4laLxGn/vWKhU+WUfp0XgD+lnNkDULXXUx
QURpTIoKNhc9tIlxIvPEd22dAUM7Sn+jj7Mwl3JJIAh13Y1JsIFUxp/DWLsLVX32
m7geqF/gtTIct7i3ZfE8VZyIhczdFty//unl33UYFe/Sgj5d0h9tuwdgyKexpwY3
zEm3RxosoMAKTcTdINrtMILqTk3UPozzSzWu5yH16FkT9JxENE79VD5ZT/P0X7dD
G5uSoNjDJRg9hJo+5T/7dvKQewQcL3hlXhflSRvMHplGIo2HLXdKqEJNvgvtu6zc
lGa3NyR3kkLm7efM6ERUxmc2Kt4tG4rZYZTFbWfcCXywcUM7xgEcvDP3fXpMB0N5
4ZLpj7snvaBeKhkKWh87dGqKxvBieuosbCiKTxyfv5TGCgU5M/0XI7YGlkRS/Qh2
Rn3BtphediHna6mtAxso15IF/voM1GJ1OA6hONqlL50Eq8N6jMwi+zq/o059G8fF
GJqzpCgLliFvVVCqPU/HZucN7mc3RN5MqYJ6+bvA3O1ioPaaZ/TTITBp+c0D5Yz0
Ilueow+5EYg187uuK9gYbpUP0K6Vwhrkd2ODerisnWpPYxEB+4CLweNpeMI4/9+n
M2HJyxG3M9jJEm36NEFZKy7XR1IQBSpAmpFKs+vPL3c=
`protect END_PROTECTED
