`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GNxkSny1m2R2B/2SHOEeenzK8opltz4FosoEXDEjEYsd7kgjluPZq+acnXC8u1P9
+pULsuVUn/NiAME1AkXbnmCid8UkbzqhSPN0/4GhLposAFrImufwzRtt1DpfTn3l
L9LRrxCa5QZvAUWzc/zsAPkT7cc0yO59tj7WCp5HJ5H881yncEif8H1HzyKZ5qXF
mT4uAELNhelWVVBBsteKhBHz3L2vkv9eC99rjDVw6iHEAiXpopOz7Ocay1Qdroko
cjyDr8wOj3FM+cq99Kzantq25bTYEqb7GH3QT5yGIkTmuZ+NHkx/YN6vWDr/HGtj
h+DvM45ILM91u6OqispIu2US3g8pOrJCZpDNxOdw4GwL5ttgo+wDo2WV2ft1P7+l
OqG+G/7RfE6RRHCSyhvulwoSs1QefOSn8haeB2YflZnjC35oU2V4T49zBJgYvORB
k461gXVTbEkvaopwXlOHoKganqCDbunoeqDo5jsVLSlwf3x8RtB66VA5hG5pE6Pl
j7srj3//iYX9Ysd6M4uRbsoMftOMTqzUtB+8CPdPw8F9lF7sG3nevH/AOkdOa4WJ
JgFtNkbHb6WpxKR78LodvDuA4DubjlSFt2rmP9eRHWF0M6qAaXPMYVyOm/bmHazq
esG7WNq31d/VXYvvsP0MQbiYwsUFI/BjXPiy0uNuTg99HTg8PPH36wQ+uPrR/tk9
jckLoqtc/Vcg0AjNbQ+BSVLXZkLe4Aop5+YUgi/ebTYIAaLb8JdjmTKou3lEZVNL
sC0UfnPNLBtHdH1mXdkGs1Lmif1b2aYCwN9jFpZ1B/kltnUIHsKojd82Rrq7P7Qa
5sflehiZmRKOu+npbzd3QF77/grH21IAMvtA7+uAx2Et2+iHcTf9oyESWT3BdiHj
S3R6E8LyEIp9885/Kh1KuCIZ83CR/xZJYZA5Fl9B+xa9Rs4jRRXBNKrSaMtr5TUq
Lrm/p4U7nzQAanfCZ5Uh/5Dpa/2U2KI+fIjh75AQ02CgFk0yPyctz5hBCEWQdVoW
52x4rZFcAdynp/EFcwv2Q/v4o0LOIx0oVbUQcPgukwBRm23O9AhuG1gHp5x7DVGw
xQs9ulTIgdzey5HU2YOddcMqdMd2Pvarn7jwStD24t/UIuv4bz9sfmSFXVwuK84u
bberwrUYXoHaSe9OmdJttw8ir7+aAnaB9D00fjJ29YL3zZz3SknxI6X8O449Gddp
RtODV2nxgQsLapzr0DSDfXFsIarNb42IICV8iMdvYG2p0HFwhrr8JWF23GbOEns1
Xj4nnd9v4poxqFTMCJZDOYVBogRmBsXwhiKJdQ1Q/cYS63/fV2NsowtRI7tFtiG6
5vlPbo3YR1Gwg1siP836QL9Yk8XoXr16EV1nbIgzSCvHgyD29hG0G9ioR1jxVxYI
5JGltGXd+RY3hn57C+TND2JhNChsTsP0T4VVcRbZJEmDL0TvGHT4IwtVKIe2fVmT
OgTiqQ2IsZrUQKC1fwOLFuaLzb/vi9RWtf3rZlipPtu8E1gPKB7powy76r13SV+A
ZBVQ96pErppWqqx5Lqd8I5XMZhVlxHHi/K1e9Ok94Isxbsnl7QhEgDpDGuCZCaZI
mpScqnde18VgBHUFCxSiB0c3o9Rtf0pXUAkQui1na1aRc5ELxS9ZNyJb4kw8yKet
u0hVjWnXbSXvfc9MWtl1LGMWmNVxKN7cswzYWWLzAOzromkVvhVs3PjIhwvroqke
eI0mhihWHV/SqZaVgOsxkz0o+2IMO1tB8D9HxMyTu2IKyC2Rg9bqHMqvAGPNgS2h
YbBLXAuY6PhXNfM1S/mVNSZaUqnPfXf1s1KjOwtjrVsJ/xngLdxW0FpDnMhS6haw
BKMeKR1gOKhP98UrP0hl/5ujGZ63yOe8Ajyz50rlmMSROgIjMlu9XQD8VXd3Ra+7
yAspngDLSP3qinapRYhBgt6SfWMdvBWSODkIwM7I7+mwgj7/YbGmKvQewLsIvnVe
b5l4y0vNRMqH/J3KAs5/udqoXa353bGXmtKl9Eme6ICy/vHvco5rorOo/RlSf/BO
Nw5qyvtfZZrPBiA5kHRSaF8a+1v3pmt2lWWD33RYZhnvB1hVQtg84X1oZkOpWfm2
xlV/SlydsdGUHf4TDtavzRWahFHBiSbb8PU/rg2MkAjAM6nIWMZ6wa8mNqtKbU7m
CvbEdE7TCl+M6Nt6RC/YsSdGC8vZ0S8N9b0Bldq+68K+X6ADMG2dRT+z5oC70Rx2
ydMtPKX0IkBx16Y0CvN36mw3BDePDwVYnEmgvJQOyAZ23eTjlMonz7isr1NN8ogS
pHtzEtF/lQqW6eOf5ZQDFdjUYf7IrSJUNrr8BKTZrZ+P3JSp8SEFEh89AyD9euzf
v3UHvSLAOhmKXQ/sp5pKEYgS6Rl/YN3nZO4UC7Y64jWg06Nn38AJUKy8SnpvYCHv
075bwMhGvBKvKXXzXjuFlHolxhZQmJDQvX6YlXB/0W6cE729U8c17sXMxnxiu7Cj
rt3BzLlwuWEA3b0AqGreo7vRx150RTDo3DUvhSIRwpWSXK2B88+fjF0Kw+WQ+ayd
NbrWeXAeMHDl680RVn42Kn+K7nY8h0QAHAPGB5Fv8M8d7EfIYpWY3cFz28aZwoO+
y4V7hh+17jFIrCde/MJDVGDKXMKagTj0i3Ihmz9/XnvLUhjZVlrJlMKuRvhuZXAU
ulE1wxCcsrcETPNJ3/212ZVPKSyHwiG32nHSZkwgZmkaVGS+1i7p4+Ver7R15jjs
QzJmXs2uHmG0p2TRl/xcViD2C5/En7HUkYOVvxsmGUJDbPMCpJeHJB/9CywVV9ut
F8srIDyTNSOyacV0YkB0FpRZusYEJ3L3sJNYqtH56T5f8RmG6QWppVdgQf2/C3qk
jGrRdSfypbKceS6MuE35dOgTH6peD2YyOkxSIHQRdV5s58v8E3myQpNxNvm5hXcu
CH2/zdLKgN2qmVHhY6oE5EN5izy6mnTg7e+5EkeNvEMu9qT1I/62Q4tW/s8T1aBW
PJeQa1kjLGpbtoASEB02uctQowyF0S6OtB97eAvG+tQ9+I6r5k2L5XtQJE4+OhJc
eRPsx8VadyIHs/7shvwGGwQyI4QJYFbjM7iOAUdrRw/o7HR3y+rsoCS4ED6vTdkL
JXrLBJCr6/vgOQsiTgXzGcZGlPw7GbpD1pEyONtblwm1/7ZHYg6ikjl6HcGCv728
lV0Bafqzcu1BwNarR9Haxi2w85DJ47wuBugGAU3KKsBYCN/zLw+kUu+S56+6r9FJ
Hu01iubd7Iqhq+XpEmz2Lu6ouPcwmTpUhB7uMh1gGJ2r1yrqeYU87T2wtRz+pq5w
c1VeoARvkxOfMcaCyYVpNv6CnO0eG+XoKcMjtybkXwyfdozE6/7sKov62dfmlacZ
H4Xb9Op11HVAy7WJlpD3qWsPOsDb+f2LwwBbGu3JVbsgRee/WxCn5QOGSiNkyEqB
wtwfM68OgL+w/J/IQw2KTMs8sL9gisLi+fJ6uGZzFavO+8MpM0Es0CY1gfwP6N/o
VdfbwyfKBxi7ibuKwWPThShJwd9vGdAC9T+8O9rYGJTtyvfJYOCSEmAkopo8DjRl
C9Yxsm4ukZLu4o6lWw7d31pGMwIUXTVhaLP5ncgRymBEQyfCNfd66lXLsnSTXkR6
oBycc+S4uo6suD+s7bztrGFrmNWWw6pF+TtOzIewo9Dl9fcpyqhjs/Rb35EqRZMs
+0NexdXQ0WVsDu+8ir1nEB7N9jZF0b1I6DKdryEhAeRF4EkazMoHMlgxB0Tj/W5h
aSYcZwCGuUAAgwKtiNbw/4YKc3rsqvtyFep8jpPdhZ12pIKzrYR+I1K2lU/9NGTZ
whtnJpYtsAAUCkmKuJPS90srgHV2L+hgxfME+TYA1YukisvhEwF/qnM7SAMEstK/
nM/leC+fBwuXe5B1eMnwwzBYnlZKVgxv5T3Qfy6CRRr2hPXVP+Lj4hP7Qh9qPpsJ
XnTaKl2xt5iRVwHRmMqTcJcaclUSLaxgyA9bniZiYiRm1Do3v3FM74zDyrtF9KYQ
9u5Ow0FK4Urv5Iq6kpiWhnnGldp1iEDKhoo3dt0ecwOk8UH/YGYfLzz4Og1U8We2
EEAv58CcjWv4ACAAIb6JlQ0CetG1RJmXuGeRhFRConwtS+0ON4SoQRGXq+LVtqjz
Ognh5Qh5U3Zby/7SDEIwho8C/w323AFpoG5yqdQs1yeBEzZKcuQfvz1dEkOu2nHY
45cZTkxgRZ76ieXmCxSpg/dkoxLi1h904f78y/5pkP+HmRoB+EUpx+xFZGb5dlG6
U7sSg0Pmkkp4nm9fn+lGuYn0VwOh/WRZBmqlzMAgpuVn2ypA4tbHnDgRcPj172Gk
dJhjoslMzaVHlaKEP+AnxW7iM7HRCdF7znyBrKrMOPcAuhYNckeg73gwFW4QG2Wr
WOMEX4i7QFrujBtVyoQe8UJiTUDmy8SiF7l2nd7qr5WODFx4/Tyq/jn3vB+s4SAm
Px+CWNe0Bnq0do6B+62kKculTM213IOQGe2a26lvBQMiQH42ZKovdBuI3NhiUn7z
zxZKieAUPnpLVPhGeRIv2m4JiVVJLfZYTYa9RRPQ5jYQwbrtPEKejNGDb3ie51Du
2xAngkWAxHycuah2RPjZMcXjyOmM2QpW73NNxfLTSrNWXDaDHjSPP0rPpYSHoBPy
/yw+g2aIH5QFXll4oV5xNsTqntNPSe4l3ghn0L6yS91GFiO+LjE4EoiIhsKuBl2q
7XFZb/Jb5AHAwIRGhl3c9q0IedWGN17Km5iUuMbyBHtYgsGDN9HmetGvyDg2+vv4
nP44I1NYGcRlMFT72JLY76ePUFCFMmWIOMazR3VUJ5iq+svOU39nNgsJcUkcrycW
vxeJsnh8P/ugg7JeZxI8rCXdTZPzQWfAVsgFIVeVcdSRcYgVRTe6MvcvZgiHVyiO
HFY/AApaZ05pUBhVP7CPKWGLYfI8t/K0JYjEiVCH11FIUiPosF82G6dqrIUrMIvl
DJS4+SjsxbkWlpT9a+qRayzPhaxiURNZ1fjyhJJrvTE9aAFLdS8EMwFgErC9E1VW
w8hxu7VHZlQddSaTlidy9cmr+TvYGYWVdmmPrBJuBr/Iv0nkxWcdzWuwFChm4QI1
u6opJODVQyj6YuR7l8o1T5XeX/eNTjzOmU9uuNeeMijxpaCytcWWc92I1lpUsdsz
8VJIkv1ELe2w0V1dWYkdfkzwksJkRRAkw05o1p5dR9BIrNdCtVqjJuQqTVh8iIZX
tmP4TDGJaG9H0t8zxxYzzFUC9tiqsepIuauQI+ZyXTRzIu91ci+Q4jY4Clp6yy5r
W0op8Z8QrvF0RAchclD5z3aD3Dx/+mFE4x7yzViAQW/Krxc0FrF3+d7AB1hWl0Rs
PkvXeBD62krW2qJ8ylzDrT0LZvOtCnJm3d+J8F4eyYbKHzMDh1AoCyBsrrIW01vl
tyMGLOUkr6g5P3wFLeY27B5NMFCvRZej8AYshEoDxX5toa1epzK/rrKKsbgzbYNx
e7HA2/YvTT8PtGfMluSMi6I0RxB452GBFY8HLy/59O79j1MtjgZwCmVQzan2MUI8
YTbYNoSEeNjIQmUbRK1X+JMlveurwcPL9U6McLoTqbm297wGa4IUKaCyS7xlQX0k
Cn6rmJPZuBpolaXCNGkucWrwWqTBrc4KAeVg/6qGhs2sSran91+NfANM6l4nuJOw
tVBBs9+4/xC45kWJUvFIfXEmrCc6y2NgLUueYeZwdPLtx/iUGKmYffl208vfQCfb
+PjGYwOWUhaonvVHsuAyKPsgcVIjD9Ol0Vat2JDmVK/j/1MN/ItUSuxJjEkaBV+x
elgXLdYhqnONHIS890CcIyfgz0+lAS3YH/Z8yR2rC21itR3UN0YKGDmb498KXD11
h/Z3m8L/OtcG2hnQmRVQhzIxNJ6E3g8mzApSr1UuDgSVHGFo4qpkRMDrNfvqORJT
7iqsGdhQt0vao5JkQ8XDwNDTAuhzQy+pJpBsKhofh++EZnjhjVF0MIk1XkD3P1Ks
uGd6pq1Ks2BNAvUt8Ab8FHym01IP8iZHJElUIYUf2UP/Ficr5DFbHO67141lLnO+
aKArXinY325BhqG7NhKueFrWrtEBSeTIWc+0sSx5bOq2fPJ13rt56L5NNtKXNBTa
4cQl7kdu1km/jNO7+TRama49xhq7G3NpKyOwSHIaIZ9c5D9vfkWB7qTO4pBZ71b8
t5XUh9vJNYZUVlpRoN5kCIgvIjvRCYLKjdIZpSxZHu9ZwK2CVQabY0vH/a7bjqEj
gSgKO8uwPKctgls6jvUILUjSrFEdXVmFO1JT7NJtAkW9tqbSMRDFOAQ/C2Mnb6sa
9jY/nzPa0IWu22hYfLQqknMuvmfGv4C5xdkb8IAJmNID0VZg04XL2VboIkgncScd
70VDQbseF9eG46lP5H4u7eClZzDQ3lQYBDHsTLeB6veXvkxmOqd0K7f4wnvJAgMJ
1XWzP4vWFN5DQXuexZ51i+befrr1r3ACkjBvj2TSM5IlunTh2WgvTSJVT+jG30kZ
7jczqmEfitZKvQUfX9Xb5PtX3pc0YIcJR9Ebi2P/VqhO0RYEeJWdzVtbLm5rQ+3Q
ZsxwvvyPlB8MfEVOA3nYaHjW0s5Px/sFbq4fdL6OLPuQOg3FuubDHZSNDNUnPBKW
HZkc6jMz6sEd6N28S+eWGy6qJODpQItJ7ywjWm8/xZjhD2LZYJU5/8FQ9LdwXFAB
cVRWZUpBxSPEFwn5Vl0oNg23xpjyWBjiS7lNCQ0hIQ4UDQ61k/WHjaLkekxFViR/
lCNidyJKumAq93ugZbP1yXUacJYV1Jlf0/5erKzS8gVg1FkHdiE37GlBLeqCKrth
5Pr/9KVZc/Wy/bMhgihs4cSSfMlm/JXpEX+w7bIYM+jPpueELSHGX6S7SWAgsJME
1Ay+j5uASe5yWIbtYZwnPLdI9DdSrm09zWNZBaVrav8qZn8pREwXrYWZfiVAgpY+
CF0dbYOr7La1pWVEnVcjFWj0iZHvFJsbRhbdW0B47lWtol8LzQy8aFsLLpw8rpHp
gSruriOWQq3ATxi3fn8KCEUcnqZlhuW5IoLM8wwC7PKQerftP5wc7s40uoFxw03f
/A4Xtc1HaqwcxselioK8cuW59TmQHn2t1Xk4HEVgLkkQAksOjnUj/0BnD5q6gqyk
miMAq/QG6qFE9s3TG8oGWCqQn0qDNSRg0x8Odnkyj0SlT4X3iKsKLjDshf1mXI/J
Zlb5+P516SeFjtPCsqycIhW6e+/UfW1PF8r4ZcvhPLDkVg9fgYgyGQSrJBRZBs7F
JarID2P4Qww1kVX8spYO/PrwjuQLGQ9o7/p/+fQRDrLs70tyQz9piXZyJSJ4neKN
7hbfsLwwrfzzCfmn9b32frADGy+9G0poY2/bKFFCFRDIZgUC55KOn4UJk+HT0oLi
R3np6bR5dlYjpJfQxKyAXUiKsCA+HjjlbsIx2KhhsaKsCQ1F0Y+h/dmSAocXIT3H
PUGhanqjl+OYkGKJ9EU8LaBJK7/f1RuRKz9IRQFR1dmSrgEvpBLqDUGZXbI5MsCZ
bGZh7aHbiZMqXiB7BUMQx/tCCbpqTcLIQ8Ec1m0Nr0HOi1N8SaQ3cnGRBswNK/08
i5kjSo1y/qVTAhcomcPzW1h17yxhlEtcUDRTHDLuroVNZJIYDRKSqXtcmaJmc9NE
Wqv110OD52yzFVYMReEGyRPmgUDAUw4idHL0ci1ZPgziQIjtVjvSbr8kbgr0VVFR
/S/EhaStKwj/GmnpM50+hTMSETBZBCnua4pEz7khtmAvVlt3e2rkMXCHDS9Ipbk9
3cangHPUs2mjotmKGCLo4rDEJebStbb14viJJ4zlqWJNHB+L5Pbb2/+7jFUPSSgY
H/18c5+VSwe00fGfXrGD/v9uIqS5ZTscJAUOfh06kkrFWpTRSGv2kMVXs4G2/Nrw
ahPLix2tFi5yV0EmBzrZiH1TU+hutJ7/tpHTn6ASNjtz6tnldsD+QT2I+ebeXNVU
YZQ751wSNwNqlWP1+3UJghn1FOD1lGRIEUKOTel4qIeYJCznU+f9Cn8+3UEjxzbd
Rlj+Px2FEcsxas+Mt9epY1FhbCOjNDWP3jkm66fhLxUuO/S/sr9DDGJG3AbVMwuI
iq8W56sBAjoOBv+zLQkAnVUAS1UBGrVTDsTtJ/JosnArXSWuwJlCpP66Ya9ko0fN
eQPukq4EUFFc+0wazfuv0AABHOvYmFuhlw4Tju4Td/h+t8IxncZv53XvjKanBFtq
3qHUaimroSE/snQxwcaddR8UGqCn8zxSg3tCgPk1Ij/QX7UhSQJzuQbUfyZPz5nW
9xZ2JbUmCmwukYbNY5nMs4ohBub7bKoRjtlMZOUi3ro4wyWB66sqSCDdZtWIqMCP
gi9smFojewjwIpA2FgoyRmylFeETQNTsUCkqFrzxGlLtNSN/azW4O2dj26ZcrVIZ
RpDrWWkjekqOd2ePd/wjTDnMTpbJm7iLNfVlr5NNPOQAIpV1DgUvxdmF9EtjKcYD
ab/swjr78X0fRRu/IQwAY8WnPzILhzkmIALOuY7GflcwKCaVFaRu8qI1aA3zsuv9
iQOsnaESDB+R9ieDD+PCweMkQwSqvpsLq82OAQmd0zH5MyEW5RhlFZeX7rlBw6y4
FEJp77xiBk45jlXvmeNsFhn/JrPTZ8JOf+bf1GIQutoiYMN3osnwQ1OpY/TAY4e0
bDqqHUzKnSGmhid+W9/pyMb7ZEeK8mfdH1HJoWfbXFQvWFpMQdq0rVSuAChozTie
WHc6OPXq0SejXUqUd+HKqvSAM28ZPiQmjxNF9VEzd7j4uB+ynDh7gicTryGprKNq
ZcjPalXYB4Edo6AzQW2s1RvdfvpevC1ay1oMI1dLjRMloXdXLrKiTyTGgwOjp8pW
esMuscBBBEoCaQpQ0fJdNgLzTMqOKGvyWtRPwM8TB2HDhMf1ITp30sO82XSKpeZ/
JrU3kJXfQwBdhpfCa34F5bfdu9Px9UfV9gqhO8okYm1UCqBUod3MpRn2Yoa2nwij
OnD9fvpk6+j7VrYKTzHFRu6hNh6Wt/nXT5x/kkVVbbkI/2lLw1nrc74VY82jK3KJ
5mTRae9Oxe9uT4FJorOFH4McgcUBZ2zx4DiSicG5Rj1jWQaSfecyWjlpGoI4f4g2
Voe9Op8bjl4hPYeep7I0arhgKKH3x6YWuHsdngIShtTOLaT+MbPu1ugj8c/jqEBH
XKb0c+9lPFjPXhBLUOsCBNVJmBH8h9aIwQIGTvkgDq1hd4UOsqYVkSryRmyR+MT9
tT18CxCOuPYUq1Dik+4gnQqP3sJIMhogvEM8celR/pj7uEF3xlhz0Qoi1OhIqE/P
eevooW2PDfvjDMZcc6duyw+RXP4cUf0dSVYAzgZJVnHHXH20jDZKIzUZaI2t8zh0
R8juHaKzgbLKhmjpae9wDwZCA4u1SgGynHvVrLVXh8PAMcRhdxITuDTbyuyk62FM
XWrsewfL1jmJYOpo4Nwhe+IoBEC+HK/9aqhQCZHDLW2i/2BoohxQXdYy3M1heYrc
fhFhSl5SBzoii3yfbh/0Pmf/hyNaOq4iQc94qCxpHjzyC2y5EdgluB7pAy4dhnmu
vwIurplGSmvYWP7tonFFmwt8h4uXmRwLAraInGSaItoWuGnJaV2irc5gKgrjaCfj
WjAr9ciI9I2qgwP1DJw2DVPoS7qoTmmG980wTwqqMPj+f88VSZQGInPXNT1FUAMS
/e8yTYfXnjVsuxwWJwqSZ+m79u8OHjD+Gz+Kxfz3B9+cnWWty0EICVSOW+K3MhOP
M5g4yFmwNFCUbvPVeq23d+c8jZk4U0njMAYakhuC1MKRzH05686NDD2meRi6zic7
rm4sp0i/Kv85ueV4HQuLl64UcJiaJeiUzP1bEUgja29LycqL3Z0wRfv/sXOOgSsy
TT0VQ1+mkTquCMPa33BpOtPPaSNliavoMz6RJkJ7VMQ9patLi2uX5JBn9B4RTNE2
IKvn0lBx5XKGS5X15s/ImYh3IBDbBn8QGCQd79aJw/fNTXPoMsvVoWRMvtoGBfIb
4Etjp4PSAtoF/LoZtJyUdnWrxxUkkf/jxguPCaH0trEVEbAay/gqrEAB3pBrZBvJ
DpYv5dVu+9aHjquJHvi6SD37E3aKbMblki90JwMb+XT2WAAqFVFd2sotEs0Od6OG
ZFM3ulC3/XH3zgXaEv6tyTz+RW1MNiqxM0Ui10MFZyPhhBnMB7HBJL3jd6EVZ53W
1Ko0pKEKliYGNJlxX+bzmfJx3Hk7ALS13U2JfDTo9+P9gTJIlnn0+xIFIQDvkBqX
d0kfnMVUgYMPYL0Tw8gfvtdJ23rRndYP6PGnsMNnDGtdzklTAf9x86zch1YCqzWr
57r5AK/iTmdfJwWydDZbu2vgTTRdHvoZM164DKHhHO6sdmHHsykoTsDc+AB/jQIz
3tnypN3ZGhTt5/lhzytYXH0++qjMjio82cBA8ao8ADysNkQ1wFxRvEQHao27AmDX
DUN0RkddeHK0erYXs37nYDNQcRo2tnceD+9OsWY2aHGx1r8BARjqijG2ZjuQyw2B
eoWjhMReAV3wNjqJ4d3tyUyfGdfdE3sqcQHUntEl+XmLzxL/8Klcr88HM0JK4bwD
CvQmboeYJQ887BnGsSlkDhMXry+ftNHoQH9PPPIVoWC5pzTZDNwBE8758jVzR1IP
+7JXw1qtkvJwrGV02aN7Iipzki4zIIrIh8HwHqjFjf5rn5A+xldh947o5L1xon7x
soF8xuqArKhdedIY6dVTI/pw+SvFaWU8/1/1jlPeuhdF/8LHx+bsAmPsnQCc48zc
z7fizlbWC9c8BiEUTxIfmlm/KYmyQ2V32FYs6uK4SVdcc2eRlHDC0CXQRNp8IR9t
wQcj4RpJ2xppeN93pmNF0TfjCMwW3BeHeWuGF9cZkiEapON8ra0ysoQazui2vIIV
e1oZNThU9eGiFz6X3qksJm6BBYhvOqkuvn4VBowIGuKXSOkE4548NPbcyJwUyaPi
QJVths6xVFj4+iHQJY64q3+j+4WEgLVwdlz7cWHwmGHZ8BZII9DOtsUtWgfc5Omp
Q6I0UTHQJ4UjaqX914Xy+wxmXEB2UsATEl16svDVFn4josdqBnByaBj55cnwer/L
CFCeI9RgcKDD7m/RuhTA1yFGbYzX5ivNNXs/wezJL4KAkGCugCjfeAoAlucJRRLn
U8JgOJwZhkmqbDiP445wQrGd6z/b8m1/VNxNsqa2qRFCgxfgCyyNght5EWUe/dmH
rMXmHbELTJgUFLPRS9T04+YL21wunrU9Kk5/FLNGN5rrB1L1CiyJpx3AkY4nY2pu
pa3JKsP+DBoJNdLi/YsUwCnpX47WYo6E9XseeriWkPHO4k6xswAQ5AXcR5YOBFlT
WWxPC9X3v2EImdSnNsDr9lY4I7o9FqeYl6D6UhdReCvObLJR6vIy1IKtI500CEW8
awR5H1kYW17lVRdRl0jHkcFZC0UmMT7qC4XYEees5xdsFZo1EHs35tQuF/1mDy4t
ekE1vPMjmyNndFr2eJDvN+VusDFN1w6/g23q8eEyBA7yAysPTMqJV06ickGkiEN7
a/ToNiyUzS8ekXznPm49vGtyWnq8XXKfAcHX6Hh4S+peJqMaX22NjgflFJ/uflER
pHZ9T5dkzirBa24jEk1biw17ZVCtTyMiK7eEJc1wdlOLiZw0+nIlrJIgd+nXztbV
AvM2i0kFdWyfU9VbC8JL/8F6cwOHOuiuhIUYl+2LHRqfKtoN9TR+BvIWg13LZ8Jq
T1o4ccJOqHEP5iAhjqY7Q7QPjRIf3e4QkdxKhB7a/k3x8hKQjs2iXpUoLzYF583R
fOS9Kz0hovMo7e+Zsz6Sv81tGgznOqMzPFANly0NoCeXYhODuH2gWPGK85ulOm5a
pTxVbwYIRZ938g92PlpLZyEGoeqWvTaOSLh31tEklz7eAzvg0fxYTa35/BKaJrkq
q+caYVZTpMwZV0fU2eq2tGrY516eh2fODS/gIf14ZhffVFa5KsGJVXyz7vyxcFBC
qFRfCsZgz+y9SMN33xvMGOeP9dKn0jrFd+1j/n23UfSHSv/i47VhmCpsy1DRrVtO
QRY373bSPhl7amugTJdOAp4bXD8HbUovVmNVF2p4rUHQUsclPO6d7Qo9cXXx1aet
Uf7eqrhu8UnqfLaDjRZqHfk/3dQY+mepRl6X9E3UJMw+d2ogSXQfwPpQl3jGHIdB
mSrpfk2yQOSSwfiaebZuy2BKnHobWciRWXypsUfsp6Gqs052622wTvPxqPXJZXdj
BcftjJh4NWMtYcqOEwaFgOhUEcckU+3lI30h1oNIJVD+nZsm2EaL4ppwojU66MXQ
Z7CXWlufPgxoe6pt6Kng9CCN0aSUDweaaB23UEuKN2M6Gj9m1eNT32DjxMNkiP1e
yJa6jEb7EtuHxIySxnmp73do569YYko3ND65IQ0hyPrOnNzqYyV8rt9QIecER7JE
alaatEyO1jHsYFHT8L2jDoaWFNRiiYywGu0u69grcK6TDYqWNhnPLlYfsBIhnAli
ig21R46DkD74rYhFltNfG+awm19bJ1+OIueHjPMbCKuif7vxtjkP0+FNYf/lPx72
qa8MckGkhIx3Gw9IvGBSnQ+L0KcXvzIeeYIyfs8YzAYx5YODwCHfli3buVeXcS4Q
Voz9cuNuzkrmMkWmCFcXEtxTt7VHLdV2zGjJczgWblEQyis4nHaCm3XSFtQBtepd
lGA488xYh3fe6ol7XDEPpcIns11ZkqPkxF05Bs0aBukSry1E2fYEEl1d6qoxnvEY
614A/cqvN+ZbYG+HoGKap6dSBUXHI3ToUE6yuAkmUyWA2O30ogMx/xvqRGe2rhqt
quShoEKioK+fL8+pMRyb/BAfkGdUziE3V2Srztfuz/4rErLZF6uRVtvJsgqjRmZm
sbgcDVKyZo0yb/Kaae6NTDZi6NccRgdgLBcdhhp/aqXMBfJhKo4qLanuqvHPCu5W
UiF88gTGKtMH7VS78cjOFAVPVpKQbGPDDETeuBylBZoeopm8Ux/39CAReBEgmQFp
jFpzS2ce+4uNK6eh7XaLByw7yWJQodFrRhvM5MRKAdDofCzuQDSNPsHN7Nb/+kmy
pgoOBrXZJiDl3upIRaZ/RCfXIpfeviNscTXqOEqxm+T2lG4a2yOzX9dD8B3W4mI1
HdlC2XpEsuz0Fyk8ZWrdO3vRRsQIMfljSQ8YiS/9h8GToedEpcGxMqkglDfnsbC1
kerN8kdpsBOcjmXQbb2Y7791ZE74Evl6W7bYXPP/cfT0fUJ4/4Om1Yv5eoy8n+K1
zbp1i2RiIRKGD3+IjOJ3LmcdRwdBkETZ2x4jo+2JMxYbDSxrn0ui9w6iG7TQFkA3
nfFSg3p3HH98tPP0S03D97isYB0qZNVqX8QEZJaNdK8WN0fv0G0elXWXZNF02e/t
Ub0WII6bFceNAbdtnKJLukGC0EvTc52T7gxACjHWAD1bOo5eJrgJzqjI1lZvy53/
0rPlyNLkXQfC3U1sfWUzxVjY8jQSpSFvjyP95TNL2flNbNpRflUSgoBE0ytcQQWS
GgeC8OqYdY68nUPWS4fW4nzWt6Thk6eEQZHfGqb3XJ+hatG5eccK2qyUGXeGVaC7
bxZ0xFBZYbbHglMGv+cJGf/WmV9p87OYcnPrjeUalshJGKdbjXYD9HopfuVcVuV5
/Bbgyfe4vxjvRThTf9wgJKz8ZODn04yOIjQjyOjcdMlLO5vMHZ3fWzqRmdMUzQKt
U2hG6Bka2jr08q+79aIfFY4tcKmEHOAQNXPef7CrdxqOPFcJLB3oydumPQDuzuvs
1LmTA9IhqxPupELa6Wfeo68jUQ9UECW8+oZHtGNgmz9TS1zKceWYiSTT8NKpBqJ/
0sESRVsVoCrjqK9jwYbR4Uic3p3omOc63xhP93jBu3zQ4Ua3yiNziribLW59JT0k
hsvlp4XxtUlrVChsonkgo72Ihtd8agaQn1mX5OLExFfIszb0Njp5Mu4vz2Akwyx3
mbCd3vK/hOCe+yPT41LGxAMz5dPqSlm0a4Eoe95TaOGZbRf+ljMTiYdCv66ch86O
/F51wP24S1fbkrozqNXDugLLLWX3qJHKyijkh0Uh1s9jGmZDqiSoEGIpdn/Gev8F
kEUV/Kq4XASCl27QLdQVrEeBozuvCORzfwKhzx7iPYtyKl2URpqqdWLW9+9sKDFY
mlCPIypkufslXatbIFdPARYYLai17THkXPXRNSDLeD3LAX8bP6cPKxV8PNv9+F1/
422Nir3vgZ/+98q+2vh/3jHNRbpFwA+rV81HR6NyCEKyCtbiNpKkG4NaP94E1/T5
NJ8VmrvRKYTKO+mZStIF6GU1qddm9ARFIQj8BusLsmBQ0YmSOLryYGoyiKOnTyZ0
VKZMkiI/XKjFh5npqlZlT78OKqm2z08Ag49AHPMCWcnoP+0nSnOQHX8XknrjU4RC
XByl6ubKl/jQtFgSypAN2g1XM9+v2cdH8TJpW0s91TC8Q3bmKux8OftKqsaWrCZk
Yn9PYSMtcF07Mr20RtHNPuK9zlmEzSiQqW+vE2JdafVYN0Dzq1O/Q++mr5mCFx9m
dsLzSiXg4HQcqd55sKGpNmpUgRkQM15aJ/zBRRifS6soHTQN5Kc5RB+ew+nIzmOA
XFJ+kkKY+pOXhhQzIQnV4BYJRQAPhtXW6/utKd5Flv2ho3qWkqpk8puN96d8sZOk
OHdX6EF+yT04/LI66uf9S46QVxlWDQ3Q6gfuFQkjBLE0SFL51K/7sMwjwoDCCBhc
4c0DdlZ4kfvwwsTFiqi/2UV2AkeQvGACaDLYJgSz4DZiW5gfur8mwK2C2/Wt36i7
5dXESuRWqN/Xr16iR7hXd4XMc7eEWSH/m9xUN+IxF0LBKtPPo8/6k0OLFGNUkNCk
wBlnPv4kP8D8XvPlLzD2ksfTJ7I7E1B0EvtOMl/SlPXtGch5Cu823stk7oGRiJDO
Mb/BCSjN9Vxepm1UjoHHkCInWPLfn1+Ho/1uTF9m/QLhiZUqpi04D3JMxCgQh5dQ
KreMJFQ82dHT4JPs6xCkTL/Sq/8uRAed/SEY+0j7U2XiV7DxG2JgK1dwImxUrV9K
GXn5Wvv8p1l9AmPWYDEj1gkEayfiXRhCTsnOj67uamb9eO8p3Z+nlOo1zZSeLTGu
Vh/FXr9ctWIjB9B6o2BEUURsZiRBcAldrqzZCRB2dZGl86O2hRbuPgKsOEcHk06U
hTkajnYiSljy/2KdSsljyPAKnPPjyEzzZlgmFWSHex7TPPT5pVSxFIIILqSwQuLH
HXU8H9U7s/kVBOg/vf/G4SUSdYJm0wPo9KlwRVWc+fOXDTX7tkn8M8PfeLCAv4lK
esg68GC1dCnkzrpt5l/BLLjRj2XtI5E+rHG0jE2FFcImVgLiJas1LTNGoawWoglm
PvQ0wE9ClSgeLUnH3JSCFiNSCv51yaWCRLcelIAMZB2l+zIya4gQD+DTvVSPn2bt
WQSFQMMyHS7zIXSYfGsr5HkiGgEz3l/B3iZDRt5DUu5662g521wirEf+7tueHXIU
lozZX/XMDIB99n1czp0XWyAf4VYI35gBp2NmEgK3KHrGPtFgVyy06pqGiEdXqJTh
si2mh/ZOvRs3BwtW4z0dX9uA9QbAQP51LEJ9iW0kmDpgZJdCHk7XDINSinzFih4y
lphZJBu9Yn56f8LejTxSU1y+mzaen9AGXO2vH/gT+j+HzHUY/fMF8TEE6hKdPClK
gLoMR7QdCxp2Rw0UHp27HPqDN1eu8mbKA8A01ap39U2Dr3Ugd98aqn0Ji0Pv0uBc
Tj81HT2LqBPI65SB2dvtA76BMpWKYuA/iDpjkoCT/oA1xsL2QYwYHlDKhf8r5Z1Z
+uv++GLoFuuCAXuYMPE9nNiFfm17VUSe9xDbbCPWzh1u5eWLbrOnTeW9fxHofrPt
tz9Jx3ImgDWYnvqACgQV+N1bSYopaGZcajuGkCJ7fEVJenJbVcpOiQ98PUUlBi0A
X9bXNx1Q4cUGI+nld/MSBDvV4IjTghGKGKlZUTkeRGbVqSG+9XO2gS8bdHEwf+oY
tIl31U2VB7St0ovEDpOeOYNZXoade4wWUlX/tGlykL5E1mc60BnFVjMuplbhZ/S+
6CgJf6yAXaaHuevaTfR4KSX7eIcknQkxyysCsJOBHDHDyJXZg74/scQG0LTL2pQh
P7msB9HAzSlN7GeKDP3xQQlDMZyNzmNWNJ0wiVieVZLlzi0em1+TK5Wo3EMbKT1B
3P24Y/StTqRwAUTB9jKwE7bxHeaXJE22yWqlv4TkVFb/2KNztSoLrDdqyABQL9LO
YxRVRZ6tmtrF6NYUY12EoLscGlvU/fYLX2YWnUscWgHk2xI1L7CStv35o8p9hucY
jW3Sxj6Ap6ck+EOA0GdKXq3VCjQwxTccaWsw+FESzaa70N09aMxvvXe1eUWuNC8m
5G3cH6Pn6B0nG5rWEZLepnd2z1Ejw0MiSx6tIEhf2NceByeWrxYUfAzlT+rw0pqN
jKumMyu3DbtNpOh8mgEhZcjyPIAWUA9Jurksj0BFHUC4kkSf+E+sreRhB+cWccko
KVZkRko0KDilGCM4lGbwXUzgf7MfPtYFsJoyqe3j5lVW16iLd+Jv01vpdJeNI58N
otWNNG0fwo1b3o8lxhBmUoOtkmLdWRUf8dhHp/xlbzD1olmbv04Lv+39dIhPiWRF
N3xEiEXYuvL2jbuWaSLAsLE0y6BruvDzLo6YI7VUUPQdsjrozvdZupYVTkeO1GuF
O6Dr2W19x6R0TJtGd2V5yEVa3oyvn0ui0Dz9Kif32H3U1OmezR2FWd/+6zpM5UVU
TgCgF4KxXPW7GmJ2r0aTGDEWw0r4+evVoNRhScM5CoZPW65C76zKIabsC9kbs776
VpE0LL8ZwJIE4ub1QN4+i3p7xXVXRbNyB2R9nM9NFbtGXlifW1udx9FeNLE/pSXj
B6/QNbwtCODSdR9hTrVW++mstFydjQIOvcM2AKM40o440icZ6tKFwEqw1txbrKh3
m5ejs+1zsLVLhTUuWQpQlTNN1Ylx6Ujift3TNm8lZa94FxLjON90wq/cCSMeERvN
94/pShm8qWG103Uh7IMkpqDnDSbd0qFXQ8fFmDQlMzobZvBT6bm7PAMwSx1IWCm5
QHd/FbJoyJDxtwPhVVUAgAurXehQv08zLGVnahWBgFrCSSFS8PuSAtp1r2UbOyHB
4J761Gc33Gf0USAZSsayfhyL4kGjdjo8X/idLb4SN6pRA1BFDV7JLVkuezNmpyuA
QTDixFhzMwe7nPpWe3FY/rO/bDTl+oXuT1RfvnRQxZB+wd6DJlIQBnzIf/GlNhkb
xouO6KdLkeNCmmLQzmHDen0ABfKd3w9JH2Kr7wlpMSJSJBktTfbXo+CH4IMmaemA
i9pIKREUTeddy7fx9VNEKvS7/ziUviFsBizFhupsGQMsvot3p6J193zL0mTuPKDi
2hYp9xe4uyNcBpV5YrX/u1JnBqU9hESxuB7KeMyEmJWQLJIbh7/93K+5GfseWuTu
1SdO2RAD7Ppo4dLvRi4r4TOlp5O7jspNXp2JROD/mmaKftfrqXXNA9Zif6mbs2zy
RwBs2HIUZkmcSMHjXbWsyrdZGKlHK8esXoFQChGOxGvjc8IlcuQfG3iU5XoztMu+
vbZYk/u9AUppiX8wY9I0j7mxpMzUl8Wa82nvm4dUcHEpRr2WoUSS1lDNjsbwBJcf
7bp13roU4JtcxrSRwriH7yfyw++VUll0De97HFv9dGyL1jm9aEE08YlhUVHe8JWh
8S35kLSv0bPHSHTwrYyKGoRao1vocZEQPmjEq63kFs+FsMOCewl6P92JgDYpbPjh
YkU5sZWcOszMCTY9mT0eGzpAP1a5nFSRJnVloe4KnjGqBaqHU24EP4hq+xi8X83H
mrvniE+9zlvxO+yZ8LBbb7VNr8c0NylX4i9PY75bRAHBWeTouaJmICakO5Uw27KA
rAauTlVM4qisLsq7hkN5qKJc81jWZ6oNeVn6Zu4y4egYBtriiiVPYhsKtWi/pSd8
4FEo9ISBJsZNXUeviNuton/zPgVQzN0y04b13OVcE++lSHYitBlYGNhcHOTpypoB
op9HPsNpoq+or9vMzy+icp+V8aeBZ/NDHRXw38qOAu3HgGYaavPgitE+mzzYBLkg
Je2Lpc/USpPJb2I7vpJkrDro+kqNhrMgAFV8EOvPn129PwwZHRJ/ofLYhdN0DYcn
8BT7cukYM5aYEUm03F327ET6qwszXntJ+cce0EGwon/2M/QYTd42B8MhsPIg2Koq
lAB15SFAIjQUN3b+PEINVpk4pMDzfz9EYF0wU3gc7PCtVS3AWrxXr/Mp+ttS6uPg
iDADx9kYf0o+uLOLDCYmPkfEtlzW+P1k8iqQY+g6oAlx8vdUqChsr9LoFJfgLvBZ
trZgw/driPfbNWKtzTxgMGbW7todICwIOIyGwATsgRV20BXRkwVX74fZtXz3Eofu
9oMEWjYFc08eLRzsZi+UcTLnX+659VlNpZ2ONflMV9+0BEWgLF2MwiIcAa6yG8pB
/gNukbTj+owGU+n+677KQqtuBvhj4z2y5t+0FjkWojgkL4n5xP0wL2Y6ZxXRJWQv
jegSm9feQ/PVSCVX5gQwPUosSutqGnrLYvcg5JFA7F8FeNsP/UfMWhSuxTAnrDN1
EJ4z32dFHvohBa8AJuR/C+anr0DTyxhnzBIRqmTTa4HKy/gIzP0T08DfXJkVpqLL
ITy0TAH/cAMqf0mPNqpfnrzwHsK0IyWRg5QrcvG8BErzrfZkG2vhLxCHBVOpyiDl
PbO5EDoR/74TPkrn7UiY31PIWHyocSOdU71OadA/JFzbH/v/o5GdUAvg4Vn+NBAm
0qGsC5Rwv1GB7ASmxggQAJT5DU5ps3WFUNHTrNxkoWQT+Au7jeIHLskh3BQCT0E3
BKfayYJJJeyMC3DUhkYd8v21cIvqjd7jf/vaSLgvVLNGKw1iSoEyLmZemZdpvWvf
4GLK4+fo2l5vnPgkaqpOw4sDbkyfY5bb6NIg+xcHx8Hro2jMSeW7WoPkQQhF6Dpg
DhZEdeLMIa/8u/LVDOWJJr55a1ILqrfKUr1nypehB6tWJOgCtw10JCvYQ84+SfDs
EDrG1kFfcDULQG7ZI+1lD2eKME/VyCLyPLUToCP0R5gs9tUG3H8yiqthyyqjOzyM
GETQVyZ4UiEsIw0CzWr9/2YfhI8JYDmTvfMIYjohaK7en5NkLJyzcBRSJzCinyUP
0gBot4kVaBpL03UF9eTbNByQmWpX+Uie9eEc09lbW7lF2EivYRiQWSLOMqQpYcqu
FdYzUtnKmxV9he4thxN2UgHQLmBjf2Rs5aBreGe3gBS3iS8dewgIMEODDqlccw2J
qObzG/B0Jw2cDjAM0g+pfaQBP5XbJpUUSqm0983QtI9Kbdf6y5VSLZV9rDoKMeob
p/HSF3q7z1+dVrlcH3FNuA7zjQR860pSZs4inS35u6iv7wR1UGnM2YkPFsrpnfJB
8+5V6zR90TBEZ8IfqQ4p1sieqsgtTJTgD3x5TnpN4scJo1ytgIbxo/Q7K6fT3QE6
Bt+X2HDY+n9V2MeHFliNtXx+zftFj/sEyQOuL2k/gpk+69xkPrnm1sESeo002gbz
tmcAWiV+h5t380qU3hXERloqo9ofBgKiPUb5FyXgGmoBptQH079N7tj5mGHFimE0
d0HvC6hZcawtLws0hfrNIwhTAJivTa5mcWETGgtbw5ZTJG+y25rGh4l5+7YnVUL5
TyAQfjEJJ8CVsuY9nbT68PqRGbfZr3GNp81Wszj4Kh/lm9r5+qcf/aDh7Z/47wm2
lLeQQA9Bsfwog4JS8C7J/dKYkjbF20P6A1xsZ3EfMqt2oX3jXEX9q3nFYFX1yG71
QNWnUHoHpwHlC3syo33MZnNiJPClkDX8XlWiGM+G8XT8p7gd3mxoiHjICY50+AA5
2YorFYulKW24xCqWDwxPVCEP/lEQl4L5xY6T58zkWb6i0Xsj0an57v5PGslsG+oY
pG1iBKExch/OZersul9AeQAuEF2Ui2QNHHvb6Ys3OmkVn/+Ut9DPZ9p8Nefqy36n
yUsIadP4lS61N+U21H17kAveLbP6xHElKo5KMOxz5Xg64Mn0U2WJLRW1JT1XVmH/
3sJRYBcLQvrHAbhEB+Fj6DA13w8TggqLL2i2VPGspaAIAOCSk41W0JX4E3B6SAbj
kGERYcma9PaWeN981ydcRAku7EPne1rMXDHPoI74G9vBchW73TOECPOGdboek60j
vZLVYmUkPkZ/6Zzcl1bCAgfAFtbMf/oJTEfrb5aOy2reGrCen4mccC7dG2AHehlu
ri/mjFpLqevX+FGIIuvuFgSqCdsOzlBH0w6qu+f4jojid53VO+s6mqJPFIMrOOlX
59PqomfDpknjN41KMaod4ytW+a0W/9hwu/F0mTGjfAhr8FPH3gGJEjRzWsof6B0J
yHGIoeJjGGgw7QX/1XDUxlNu/q+EU/6sftEi8cqFBWneV6nVlNdQ20oKvneQfJxa
9eMh8/p9PIYZv0D0avRq6FbNmyXWPECZs+x5ilLsl/mhLARl+8POSLxPtEQYYAnX
9X/NUjm/sZDZRnpdwZi9Ac7COVDfKLbwK2WD3p/1+UbptjVCq4D6jAhMOHIdRsWz
1+5J6mIlnMuQRKz/Sn+dGwEEqU81fVkD6Qu3myKi7ViPKoia8TBgytk/xdiRNd5e
GB11WNocuvVbh0I96Te8XOmUTk+Ks0Go6Nr/A5xyoI2dmBIGpDvKgI90Rvc7jUqh
fL/dNBbkFr3E6pe/O2VxWzTJ8YWOXyzkKRogKQC435329y6n7yYz5XNAt9a6D4lN
LDrscpu3wi0lYaFftrWFx9LJLBI7qcMaKAAs4pv+JKRWJ1dUoI3QQBpQjIYN7tL6
nbVWk7T6b1PJQl5cugOoyBpC7xZMadSWDAVg6NqiNqufdCTtpJEGVvwUMpGPbvl8
quNUSa7rcNjoopbMHjqdtE2ONUYi8ACS7JNdxJQ+ctFQqfM2EVcEM3YtLSE8P5mZ
LPpTtXWYPARWSpLcNsU+sE/WYdzC4SeAERx5bsDsbIQHCEgVm+LhV/UAuuIuT9A3
0tt2epExbcncwrjTfBl4g8QVy6vSuG1fTQwZDhNuf7lQ5CsTO6gm/yVrGIaXf4qn
vCq799ygkMfsSUr8reFHHzv6gW1CrORGaD15HZaod3xC4S1doRCK7jO5JXIkaryv
WmUNMGfgSGOYjvFrnFa/RQRR6rkLE1eTSB7PH5gX685aluFIQOlars+hL0IB5zsW
bSHZGYEh9B19JM7kz60qsmbGkMvT3WMyuKq6KJfYHExhsjh7kVcQZaMoKEEUg0ji
UQHsP/yMkTgEjFqxphETKY6KRmMfebVKYXenOHPNv0k2kXl6uaSybXTsPCnwYmgI
vM396jLiBDvQ0UVA0HvLw4c3IQqe6T+4fIJHCTAnX47HWk392eMpX1879N+SeVMH
Vb8L4Mh3cD7F5LeOUYRwVOamMp5x6yagapdOGKcnfKJutlK2HtwtvKunZrBfkb2L
0Fqha/lRprq78mTQE3I55E5lryaIQb8JTKzwtal9Xqi7EGhnBZKvvlVR6Kia//EX
WkXxFtGdvHgO8IUudDVgdxGVqlLipYyRTTqPvPsYlWXV0HOL8nLar+PSMW0wY/07
pLIFVBWklC3m01mwpPwxoiI8e0vcVrce5psxTGuulgTeHi2snhWaWKzHHf+cBBFA
g7dX5Twsikbh1xPXUBw8KZYdcHPxA564OcuaKWRJ4a5E9AFdJ39tsexyzFQ7dBwh
vLtcjlt/ymPX5PhDcm+JVyOfPU4OhXsZ9O3kqtfdHAfJYMcDLMYb5TdoFKjbzQVN
Sn6ULW10X6OUa6z5RuQK9G6eHhI9x088rwg1Jeqk3ABTrT3VkYPGwQLRtF8ehUba
wLuqu7lV+whQbTt3wKuM6MrfNInIV7RQ4/Z1+XE95fYCvjKAhZJm/Co9ydzkffxy
1pzAWUKiRs2k4PvyIDWP521wtqmj94pnL/00olVF/yvx6EnocEU/V6Cx1hTNgD3P
dbgJi53mJDrvCo3p51/jL3XpgC4wVItQ1Jj5CxQrdQ0q4a7btroj7HMw9KwK3j3r
nhAzv/4+54unw4VAEgyfZ0mX7k3o3rRYT42SPy6E8lpYODxU3ECg2OPAwku92Eii
hLPjzMeIDn6ExgifcCpGYlULBxda3hvCKkDvstG0GBnBp1s/wngmd+6koIfH8AMi
Fcn4YAGoWdwNzfmJKouAP2puz2BsMupPLdOUlwvWX1hW95NAEtwOKZkSFj1r5LgH
wPBhixd8GA8kIjYPyXQMfit62pbZJcwS2VnyHnXusqqu94tuTDW5gPhCpBWpDuA0
eCHldZ8zUM9ZXOAerq+CBSDIf5/PUXrqvVAHOzOrao4qnk8vIW4QzUONOmQz2F0y
tS32GaI8PGgmliCDcxZ2Yog1ZuBeLVvLjVtJIdOBuI0KqoxNbkHuxkHfclaA2qBX
9wB17FHJoziRfPxF8unUtwjSiN7RLdfz6EptqOl1KATsSPd44J8SydGxDlGGtsGi
UZJLV7cgw/XxpD9Rbp4Hs9GDAVD514UV22oMu8E3+4sdEYITyhJIPio7cmULhBGp
MzQVwc8ylWBVdAk3zmkapEZfQZmXsid78KRAEzftUSZz/0ugcSLmly0d6+W9Zp0Q
mTE2ZNik1Rtepu96CvehBEjVjrMiMbXVdkLP6LWkTvP2dmC8G/A1VEjmbOkAhDy5
aJ5O1LEWqAVCL6uICYP0ljVXgNtR9zlLUZOsmWsDkKrHLUGbixxA95bF6zCnByVg
pZTrn8OAC72RV93BoxI6KcbE83jZlI2mDstpbzHkz6kGO8Tu2AeM8Ea+gE/TQzeB
bBCHQpHSzit3UYG6xuGv6p4NsuNv9NDlf++nKr+we7q8C2XIO8n7arBICxs42Gvx
Oesu+x4F3FCg5En8+ihl7kizVJAgo3PYTp+GSLwEqTXc7s/yy+CiBe01rCzjpLmZ
HvHyZo0/jbd+McEst1GMpWeDPRR16OJ/ou59oUZN0BnMr03g+jdrlEDNWREpw/ls
trNdlWDK5/l1bQOkcXB6dA5ZJXmQNtJeCHyEZe39gSun8oi/jzl07+eYi3OgvzgN
UsBC9Y2L29fTOOtEJlZ6satSFZ4ArTzXNkEijA9sBPHlyHvlJ6gjPNUmnLIpOAD6
55M7ZWYf+xP3KekWyzzTk8ItC65vXJ/aiOj6fzcVNGemNhhKiIFKezw35zwPLkoU
HdoQkv1YKhQXUKthiUscWTCBxgmoKlDLoLc66blt21iMRB2qbcwLfRMPzhUj4ul1
k2myWPNxb1QrSWozpOnIRIgu0z+2bZ18aLZYN7fCXi2ln7uoFQEvNGbzIakv9SL5
1obmtSAYhDirij52ga5HBkX9T7so/HcUbhlVsXPP9E2Yj5d+hxKlrabDmSsJAbqu
Yx4rayvTR8S0x6SgEqs3hdyci/cJihrsho1YRzH18MtevFxMqZe/iE3g1joqan+P
gmvHvWj2hRs+a1HuKI+p4VoTmhnPcxAvSJzBtZr7LyBzUARIsFlxzDyfFnHln6O2
Nm/tJYCfdEWnvPa6At7Nl/M6UqHPmurvcha/yx5NaTSmN5JRfp1PC8zcv53jn5EU
xd0z8FKeMDtK99BPQfOR4pyR1WSKrV/mI72wN1Z3ZI3RfAzFpceJrZt3E1aL+Ic0
tz4EXNuP58CPBCYtCtKQduE3Pr9n6l6vVkDRSwCN09sra4QebvRu4j8Tuuh3FGRo
gqnHjuxN9q701xUlMoCAtXNWNDa9YDzbODNx/4Z8PWZCu6eolzElEcd+8DZrV7Nu
XHlhdqdjDkZ9QrHvcwZLKhOuJcwkgRoZ9mH722G2PEkpsgq6+uz77FX4F+SRa16p
lU1b6vkTh5ktU9sEhxIniPPdcZvL22gbli0hDZIVDLjgd7i3kdH9dLD4513QpQc7
yF/qppuPpVjBfwLqMoqWK7LU7PzIVrnwwPL0sJmhrIM4IUmg6411JMWKz0QIWZ6/
uCoD24RA639bj4P4nPsZzsDohYHx/DwuzvRpEVS6GcFh9b1MIKo3nGMzCZ5QhUGu
zoBwPZV3iIpgmtpsPxIkHXwNCps9XlInVZHBKHywLzyg7jXpCC19apuhiq+ZHQD5
kVgji8A4qG2UUhrGqIwYT4fvI4zK3qmv/QYM7wQpnmvkaqwvz06d5Qg13Eb7NJBe
ViW3Rbj1GyGjF1YzybYr2pTjP7+K3vtjROJSnfU244XBChwmvpgbfpa/mIZB8C7p
FtiKCMZp/vJulhnpmqkQ2mz+qwG/bECE22x0SYtrNFcLopWK7+Hg4AykdYaylI3P
JaCiAJJ1bR2m4ZryXzTWdHH0PkW9N7jTqZShqWPKjJU8rEX26nBLK5jJl0lQ1H9e
JKLG+S4nBtra9uUka/q+HHZL62tAwyFlRAIxtyWMLSh8eDqa36iWKAu0eFu2YpSD
5awLmu5RFWVCZLIsIy3xcTjAgwXkb25ToJuKHlvLGHAbYtON8vcqm2OxH6W6R6Tf
rjSQqI4wE/ZoLPUfEHL40/l1YVr48FQ8hNebuIuSntcEWEiSL47BRIV8cncLx+0K
v0bbTE0AGwR6Lg1q6eABo2UGPDCuJ3xsX3YgXt8Ev7S5uWqF8WiO6lr8rutPOG8R
Hy+8KYcl6wGJDBcmtMn7md2TjjlPH9CT0orfBzYgHEMO9wGo71zI7dQAPQH9VNxb
wayvkyF1+MKEy/3hCAWcaTrvHfmjKO4/RYsa/okGPjKR5PKCmVpU9vE+9/kWrQIL
AWNpEy9zp+7SyPfp9FPDFyd20NyHNdI5on+nItbRxnRhW3dB6sKYmjQuKeMxHtHg
uiJBUsAlTGi+VN67ZXGtEPYWMSaY10Gwxj/s9ih/JO2W8ClG7jG+3D1eMggVSBWq
re1ZKeE1t8t4IKwVxcOVixmJnYMo0En5VHNiSGJIXMel1ghx/Y0KtME2aqll77U/
ZQbgIBal/6xQuv++9qkNWKxf1TiqTeqLSxTP3jm5SXPt+nFR+8Mp78GS5IqjtONq
bczSWOPR4izNmAxVqPUBNPbKNkokEUhKdqCtzo8N/vnetB6m57raMi0+z29OhtAK
oY2ZUyAclgwNXwLGFoiBAyRqRU3ae6Bt3RLVMsOxvJ6FzKNuPQBydLUau3hWiunT
htw8kJU/YO9QTgSoG81riWickw9VfuMGVmYvQ72g3AphQhm3bZ2yYETmT7lynbzN
IWf72tIS5JS4kGWo2Jim41tpAdU85W8jf1sVkaWCWcjRf0eh4BVqW3CZejbIpvC1
II0VmaiwUvWgrk/CSwfMaDsvMtzmNhQ9DiuKToOuYWf/arIw0CQDF03HCe9GmCU+
mLys4bDI1ziXgHb+yYCCaUDMH7q4UHhDjw6nMC6icy1xE9dgLwbpLmJTT2pXN7wQ
S0AfFfvwCdmWO5FXuim4Igj/IMM3Sj2aVGVyytC9UHBIgV8XcryUhtcvtYJ5/EKv
3gD3xMSntVHLVaVehIkJ90kVLEDZ4RtheCS6qmRLdXTn8CYCSdJ+q6TN9FbOXL94
gJLNCtUg0kAATbxq8+DuLL84SOYbJduUX13jPQChgjGBlezjUMyXxUy/Wv43Qacb
LYL9i/r1PHz6ohNhlwvKL62y3bO41j0VY7xkEQmH9kX/9ryBLOhmkcfHlnb3/Yhf
Gb4FxEJwB+jwfTF72aLJEQ/uKzoVkfVTkISIAlvIvewftyPUGTCvLRNCCChNt9AT
5IzkENYrZ6QgwSIk85ktvdkOHvp4G6zvD41CIgjUFXfVNcLQKjBiBBP0dJVLJVmK
2myIljkDIWI9KsdKUDLZKGX1gp2h5PBpAEUJT1dh6BzD8fa1EUt1kab67qAA0XD0
dJRNGxwUJcHhoG0+LatpE2HcLrrxAUBJDwR1GqRFoz2pwYStytanKwZC1YWstr8N
sYvNy7qWpXpXEEx5CeoE3Aq/zDPb1BfgR2feRvy9S/SkKEYX95p3XYPDIouvNEWo
AliHo2yXCH+Dudv4w6PATi/uaXFWoIHY9ciHlcr9yNlaxY26XbSjjNMTi6Tq16kx
v6rYzYSnpzxxMYg2+44EPiGPN3jYJ8mSOJ7aVLDNrKc8gfpVnPndNyVy5iAH+yiF
5UKFyxrEB9lDKHtu5wEC6MvL4wLp4Hfsc5Rikv3m2cYo4cjjKqF9u/9eAkoBxDrd
3gqUX6NNgz/DwoSVdRzzZXPKbSA4EoVQBmwSQ1KhISym5BfZG3Egj1SQ9CvL50HQ
EXXME57pkan9FMaObvSoQ4Y3D3vnYy/JrDE9xtmkIJyJgsN/fPlaXf1vJi6X15Ge
qY0VxCol98SylMciIAKtCKy3f2wJtoUthJ0j4+eIvu7hxh7ueWMw9xd6aATtOMnJ
/F4MtBvqAEBjNICogG26cUxphCZs2YcqRFcyK/OukFUIw5a40WGOG1NhYdXRFi7h
zKtNdF/s1BpZWp3zCXQL8tQc8uNniSWc4uu6k+b5Q951LNsfxBDvIaaGTrekBwb0
KE8KIeAJDiSAE1KWMQCtDh3aw8n1gNznOo02VUX5NM0A4MM1uCSvSKl6KMvXbUd4
4CyjgXsSXIQWPIlOGtQpTLvgxa/xhODO6cswp4JCLxFqHG5o7dufsbwUXq1ST3Ez
magY+888U9EBTrUhxGlSU/XoCYpcawtisLa+0vKI+L7l6BU4btzK50X8tMTLhrvL
KzI94ZA65NbEeTe7L9XHbeqU0g4rUIXQHHB+t3rChAp3HwBCZQXLLZ2WDBJ/fB67
7raxTCaUmJZr/Eeiy7dIKuusTs3XPvCiQeTQj43YPmDrgQepoBplZGqdgOr7AYCw
/ZYwnC/YdUGcxRsIWUyqn1I48IZ4eVVTYxrlVA0nWTQXOdlnL+l17xzDKvuDpe30
CmFwu5iyX3dZnAPcJWOmBpiiOhOOz869zC2sYrNI/RDHjQcfgTmefBr3x0/sYO6V
Vg+a9O9HHTAgQ3JmtG+JD1Hg96eJ2/qoLUJJl4zNrFWqKK6izu0+qN7CGoaJewPn
KZf/CUVdhgH+V5vDhFv7wiam8JXNtJDU+UZOrvgM62oEP0F4MGDqU11vbx13MVk5
MbUBh+vOw1uQM1++IFtKMmKX5bbUBVo9ZhHV/My85UIdMWRk2JvzyVo/HQ0MDJ7G
896w6r4ZDvg5kKAkf3VpaYigFjgs+FXqhBnYneXryf0rdAWQZMQ0942QG2kQCLtr
5/S1osovmQrZV7KT606byf1afKiUR6gPn8V7XcQGNJVjrX0li8/RHr1nJwpPx4Tp
KYg3NVXwpz4w59ipf/+ZWo+7tDFqKXfWDQxMn9OTNXDxwxZUibUyI8dJK0RDz2rT
NVJFV7G/aEHZJq4mr5GWwUT7EON1WjlddSbbj3g0D3Vd7r4x1aIaLq/tUnpbaf7Y
++C79bxPjhZRYdKydHDC+wCm1N0rmFdij3+PQWnDQWZtbjxsGInqjpFHXjRv70Vo
ShP4lX+8hrJBk7KgtMyR4rUhrt9+B8KMe1df2V9QbraP8yxuOvOj9EXKfeorMYq9
tyM60Df+GuEyBxVuBOOILCOHd2e8cOuoWthQNEn9K3ggoxw9v7rSuQqhz4IQnnGz
ZRKxxjRmXpScFH4LwTtPgN2y7vybZ0Te9MzYfKAaC/dJhbueK+AXHTIJIXMmxtFj
ofLgrzxrYgECbMwModA/otkBBiXgwXwMmtiAm14v1nHJcAkJMCNQMhos9gmfpX50
tUNfcQHpncJ5uKa83HbW7iQjfuO5x0Q901gePjYqd4PRgE4WB9Q6CR6WSX5LK2cV
9siWK4oc2Wg5p+tHfqiTcJ/UgRn3t0Gev0kkz8ApImdhJ83EWyuH7xwzrqmFIY2r
5zFi77TGwP8Oq2fMbg+QwBB20IKcu0Nm9lPEqyjp3If13sLSQniIXv6mLe9VA1AC
tKhoAhOv7TtZXvSAYFzt01p2OjD1NE59INgxgfNFG8MdwBBRoa1XsztEnUb2X6iY
50VfxECsGzTCRe9cyGI48KWz1Oj5Z+sSFGBob6pV5kK6w0nvumQBf2o+MmEXd8El
JTzGJtyHI54e92FHsZisHyyRez2qLEnWOyPAtNSz+LOsZ3oatp00Xc/Z8EMC9dq3
d/VciMJ5vpXGThFBaw38yOGEzP9Gw6pdxsEBndSWK+oWNqh7ukFJOkkhgZeWF5Jp
kDYugf+1Gm1exOb/mM6Q901U0bsKjNeaEHFreBTSMPaSx0qbOBLlu7cKNE7YQ7il
qPwHvuyuZRzfKROVxMYl0KO802zGgQPKC/2BvYteCJolbnYd72g3wZ20jWcxVjw+
l7DNV1ariCb6dVw/tfrkeXQo/ykwvq5Xn1yuUUH7MdizuR7i6LFd2m6dQj2FcTlR
TFYPX0X8Lg3KYsF1uOOCIqmd5JIhqmOtIDJBYkGDIADuNWkzEZvCZmxYNOy8MHSg
/suxc5rhrvLRWE7yMoByYPPyDVlu7PS2dl3x2vE3Ua6xHjEbIY325jICR9SwIe3F
PUnlkLTOTcL2Aeri0uHEY5CZWR5sZKCzXOE3jw7V6/Tx4UufT7de8v/blsuE6Gyo
w90krLHxaUHhGBfV/Cf9P4OnjHBaRdUAfiTghPBoMZtEmSS+/nb8lSJGcRKMdGjF
eybrhzgvPlM7Y8T46iMNT/ON+/8mVPA54cdwyglVS7BmLKpXjIfxFk5wke0Z3/sk
zDeO1B+Bu6rbe2fGTmGllQzTxKp5ZVCh0g/dQRoYcBc3dstVnhAIVEnXh2K2SP0T
KLQ3CfCMTXC++cUVVsppuEdKxHcX52CnO6a+ulG5pqjw8aZ+f+IQzsptZ4uxoeoH
3RNs9WdwWSi+7QApOGB3kzZ076MrTt1Y1SlUlF+fshgUHdmQD076hB4kRirXXEUP
JbHrIu6isjQHsP+lgu14JhHoxh6pQ/wxYM4GbmUhbylZqXHifbWVkMxC0CZxIM9c
p9R3iNaOFWBdag3qs3A9fAe1m5ThdekgTjlXSQEeFgc1UAbflgXy8g5ZHlZYdQFM
FeIq1rMgFcOTe0Biv2d29qCzBiPX5jPcwluRvRXnzbcShcM4uNnPQiYkx/i6zqzP
RP0oggXQSOSqDJ9YH+lu6+7p2buuUIwbRGYsf6s3AJGLj/katcdOumSqAC8kQ9O4
4Cqvnj30Xojm8+eq2MC2Dh420hSGxQtkQPsmfOSSR5Nlrrgw7Mi0BaMblGVmgVhx
sxJ/dKr6iQLTZMn4sSXmuW0zXnkz5GVm/E7/zfyHt0GOq7T7xvKfWs4ZLVc2KCSG
YE4eb/7v5mJp6aF9bb9ToQGWyEgCwtX0bu883Q4FaP7d5i1h+HNqN+fMlZrYSY8E
vMEjGfpnORlZgJdemyeWdHLUXdb1Y4ex1522zL2/E+NXn8gQEzae8exQ8zhySD/a
bjG12GOn3A9Q3+4eYRAKBu/eCZFvA6fnWj20Z+TRNPxTg0o99NFuv4MTLsLUKxQa
YgF5R57Akd7eewINyKALzPiQUbJgtWKzNgeVBF4X4l/0NB5CCPSwKM++WSrjN2U5
mQ6mJuq62jZcGIRx+xBDupm3TKLMwwWnsuQRzRvqXaDvkf3CwePIp9+LF+jQxeMG
JFDd/yD6sKto5j+4h2tQLLSRiV8MFbDQllTYoamoAi4yJOYvtqUp7aXzKJlKB6ke
vqb3l/itiZIenOdsVAF/Ig+H1f7Pn6N+Awb3C9YkQ2hVgMBBLOjT4rm38GMqu/Di
CXJ20dNFU+WXBymKjSVFPNYQDShAtoHsYWFIcTz/81MdZMdsedd51eq5mrpsfvip
i3IBDfZZunNjJWMXxoV2SWGjCkjLLPOhca02gfZAVRYy+vEzGd6k/NxaZphJCZvg
u8Gi3+2jJh5Dj1yUvqb9ZzpiS8sCpTEIaOK9tO3xLIZYDEb4ixpxK9NOXC5dXmyh
7z5naETDulCA7EBuKgKOJ7n05+sYpydDkxsNiDE7APF2MSst8hSczA0wW2c78laZ
oiCEyer41HCSCRMtIruNcM8sVwW5gCMW4hfRyhQPU9ZHRqGM61UVTMRPoSfmfDTF
euMrGtT84faJTwUiTt4GpS1g2khbkhuyl2yPQbvm3PwiNvPugNHwMeRpM6z8Fgud
HyPO4lr2L5v/aFGKtzU4uyzInu3Q6Vphgxhj30lMqP6jr8ICgn0RC4P1su2EelKa
NlW9wmMTM37XkvM9ewbFYqpKiEZ0DEOq8HamtCsx1u6Kli0KLGl++y5NqAqrMIqB
QFqwfVu2u442I6z0Xbr1u6MtwA/8SQIzRPTY/LtvD2jjPapIXCJHm6FVBaC5Y+G+
JkoId4LLfT9dgeYsj0v8RNn/2xBhFsIOP0eSoexk+uf02qlgDS3L4e0LMxIF0CfK
gaODwhAjsu9vle2y5I5PzUICvMXBXLuCG4upRryKXRMlPV6BWgVtnLajwFHemJWP
o96guMo6sCs27GWqp++5k3l3IVdC6CQZW+LwLCsZLqdf+Ow3RTq/bF4h73EeRFT2
cZvo47ByE0BE4VwiYbLoQVFJYeJkoyidjkzjoCWVwEAPcwQJyvv51ePfKRZ9t1oq
Xr3uwExnBFLL4APVCWnkA0cEtpN0RmzPtFCs4IE/4c+kZKMxtqspwZW6lDuoZm2d
ANB7RiynTe9la08cnKilodewA9HCTdNQElAr2tBuEVBla9ZAKVfkG3QsWW7eMg7Y
oUABBfXEU97TtoV+g+LoZ5qllCFVWJdmF23M8Iqo9qPK1il87de4Cv4UmnS7ht4f
hUZknHeKY4uhPuszIAPrJY8Wlem+jom2g7O8SZjXsD2++wtvymAkjezPqqL9AoeD
ImYCNlQsewRpeQRSgtawJGUdXA7ynp/+XVlGpllv7xAaOo9Z+a9CmoDkvxF8TTii
Wnt6yClSr2SqiqUIv7WVYyo7ZgjOhrTiAjShhbC3BT2dRjwNiEvz9gprXGeUVIas
p3Vy6T/9/a5pW1bHrRBGWhzDXbOiAaOmkwMUP77qOyORuBDsjJc5hOFL0j/3lkrJ
rISZryCafNNG1OPFCsf0G/+P4oGKK3ACD28z7GhNEpwTjfqlI7GZqwsAXBHICfGy
vsM8QFUZB6Euj6PwB7Z0/NMC88QpBPF2xhpgs6ypdVDh4bDzSd385cpRanLjZ6w5
ycrUpITchFxrlqAeRf2Nu+QWJiZqcnElbrKtB8Im1El3IyMgJvl0ix5eQvNEorkF
RdgdjX6cYWAXbOZmCWaNyrByhShFELvmP+jeYIwawJ/KB7SX1kSncOKhaDBTl0RS
9ORwgQ1Ngl4UsJqL+/UAsPHrfuOdb8jKEsEtqeo7n+5dUDFvbejXl6CEgn0w6mg8
ZVb34zNXB0yZLqJFbCx+5kUgFbAHnKQOqLcZ3lwy1McU0NgODYsZ71uWM6ZJvIe+
DYvJwME95K8isAiIvOke3BqtfiEaV+8wttHFiRevWq61z1GN+DpuwjTOHgW+nku7
QKmOMpkw1sxIMz4QOpax2CB4A3UHf2VRyXsoSjAtflJ2woEV0i9krDMBsGWYkjYs
Wl7L3pEmSkVJT90nBSB0i8zQrt5LX5Gd0iaAAIaCtgwstQaS/aSPT8XijqoyWd4b
M4jq2pTMccpMvdP5gkYGHNAITFomUecqpB+PEbD4/dno/1LCZg4F9Otrhd+ZFy//
3VZVcSHpQ0SuS7zpTkSSO+ay67u30bGZ9uO/U2jTx/+ZY3508m75MI1iPJ/sOuGZ
tjeBapWtQDoqRaBl/B2X0ZYW+5BBY1hlrE/CMGGNGKkHXSTkcXu5p/8CTM4dmLk3
PsLOA9T83bGKsJEJo8HyqP9fTHYKIZgQQZ+jkjqNQAovDreMAB6b9hNWnBLsBO6D
14Hc7gukAaLKCYp4YD81AefAtEPlTxrU+FZ2YVPbwEnq4Jxdu/nBL3dRl57jKma2
80jlBOtCNplJfr7djWiCkbxqJEHJCLg1G5JmuCYdgt/N7s/aIzvrwIg3PhWuLIkw
SvbeW9xa90TOUUMJhvnNm6yYqz40aih8v2NOm/zvb2mVY/WBU/BEtWUsjFD6Foan
U5cZD5aM27cYuDjnDMU9peHeEFu0mGXPDbPtFfy7MoLPiRSWhs60TL8Oj2iF6zjT
XRU3jqFyD2Bhvj3mJTIhdfydb5CGutNzF2BpIvsf988hDKKkgrB9+oG0Gnh3GAa0
4dC4GAqx75xecJbtWu6hbDbJNZCRpjmaSdi2R1QsYCcLGdhCcm6niZq72pKVPGnJ
7zn9ppqDqS9bjkGopyRPcvgHGgCFUqqbtF9c0VWz7jpdVuG8NAuN8n6hCi1Bl21W
PcEcQRjH1E5r7lTpuXwt2IEOzNq+WKgy+uF1s7lMazc+ANh9mAgvBsAjFWrvBYmn
cq9HfBdarN49y0+uUx8XuT1vkNV93plNxBszDVnDEmW7QPo9AorK+TrWDyp3bJjZ
8K82hQ9aHLr+fXPBqIX9dotv9YlUkeWHUQ/EPFIN4kvwJ/88aEQG0KCjQxkX3Cgz
rnGrx/8GIf7XNm9+c6AeN5OBVQ+GuAjSPevEjDRmOgJnRNVmGnKrHzsihzDIeg1A
gQgMwAX5o48MHMsaZEymQRZuLIB39gBdcTjP0emtg6a5euiVpmSodcmUofujrrW4
C4iVWFazl0SC5oQ6DTy9Qwlb94+lsoxA2rmsWnGs2XApYGtEUZQpKDPaLne13mGh
rvRnwKaHhJhcvbY9gDmGaE4e22amadeVOXbVe0opkFFvqm7zZJKzCrRrsOOkReFo
XC50Tc1vb/ezn0XshUI3HSR0vkn/wGQas0SJf9DIcGcOfETzbRgfLWvMIP+ypzQz
LqN3eWzIPDGo91sszIFvqMXxbrBV3v9jSowUhIkmKCE+dTdSADHhZZxfiuq6XVd5
pHiAgv6jQ9qsFMyXleAw/VxHvW9xpRw019Z3j2s+56RMIC/7ysAOMPIHckwfjocg
Fyic5ricGcAOxAdBc9BwP0u7RFMA+LYU0sgtDJSNP/MbDjvD60FBM+NUBSr6Sbgh
W3aVj0UoXINuqm+9aprCR+E3t2XDCfLvkLyysc8jzSlxDxM+N3Ru+NxLd95QIRnZ
TAwmMwb33HI2xnDU9Vq2SZqzPLzUuXD+uq11RyfQYxfwjbW4o9mn+yiNH/OtC8yW
tG9EdQ4HPeOkQsDi9hJb56q3yaTluY9/VkcJUeOeo4nYXK2qm5eY0P62FctQ0lQG
bdyXHc4lAddTp89KFvw5FDgnHSa41brCc+YxVq4dP1re7GsI1Nx+tkZbVLYPsor3
jUfMj+269yUT3XS3ZYnwEcYCrIjh/FP+n70lwXBpq7+aGt7dJ2sdY0u79Py2i2Sa
CQAmcsD8ISzwSO6M/1L+92lb9Z/hfT7KgvjgRV/Si+tUxjqmwGYYYIuout5i/ZNZ
ODtV2FpdFP0Cr3eMckiuxTp0yJKlFabY3culFxRUXP1TWAKiR1p4rpeG5wiqCXdb
MMFKaGTG0IhYyvqzid8QHLPi4OD/TZAKxctsUEldLG7P1AKLaVKgbdKesOa6VNzt
p1Vw7kqF4bcSq9oXYk19DSqOxU6kpsRp+lR4q7bg/HegEbgfDLZHMz9FQwODLKsH
M22+FhKFH3JLpy+e2zOIYHg5Bx/JogN3OtrlYr/1Srq1YY+Kym5MXUvvvztYFhqE
ODcUkg7XqzE7l5zVQLD0E1TaCJcnu4pXAXcBitZvHckkYRUtFjxfqUdv+IErc87f
mDgb7oOK85gbxmUoriH7nA6iS16CXMaLFIjVw9+eJ0ljcqgtBd6oTQIvO6tuxwEk
68SwnA3FS2d3fSpjLfqalRdrgJRxRZ2lZKc5VByWsIEvihxeYBXz0l632lv7jXFE
yJr9o+ldkVmR4aIFttdJcV5vokQ443cnO95AxCyiPRP9RU9Oa1g4lh0YgGUyLUBQ
WSSgasCihn3g8Blualy256ZSGRxl4gIlDiHQrWK05JGmXrp6OwkDCcCOlx3m301L
vXGQE3uCli+CwRZ+LKTCVOsfl9LuAJ7H1mnrYWOEgHFYCBmfT1EIQoh2VjNH+7No
gYRTmUXR6HEu4XSJbZqCMgZFzYY8+42X5GqQbkK1voXWhF34vBSCxv3ygwdGxuli
JeEG/OCz5lRbe7ngysNdgB2Wr6ZoCbKZgseVfVK9oxNJ85BCqEGQqIvYOdVJERBR
aHbvdKQg7lCVsEuqWO6hHWjY1LMsGu5ewbHCfFwpl+5J8jslsfSCwNoz/tVtfEiO
eh7ovuUzRwIcLchOgNKNvXCLaDZE1Df7QFZXC5FFLtDPqDIhYBsWsEkWf9gynBkx
2MlCABH7RWLapmPJQQguPleOb8i3rWCn6lC4yZSMqD6aLvH7tfop02CEK3Y3MQcI
xFxleJt9tnObjIYgn5WvOTVt69LQD2TOuK/yfGNipS7p+FNQZ9sQV6T1XOVsqg3v
4scd0SfAJeeH7LsOBEwW6HZbEH1G8rwme/A/A6RW/HrjMLIW7xgoPXHFrBZUmzoG
0V82j6FrbT8Zjgh7R09M6JyxzrElhZo6+E7mcxoQFolD3hT7IK5OHZx2m9/WM2Tr
dmTyqiSG3GYrmGBp2bD2U8/vvGrs/eAXQVw8FrFCHdgWp3XwK4kqOg9CTqxDYEXa
ESK5sRGcTTtdJG9HQQwlARd3ukOh7OUjzNyvHOmNqUQM7PslU6T1G6oGl7Iohr2d
LDyOfSLNZJ9Q7B6XeMaMKZigdehE3jfKNsHhgzEcLpV2v6vYad2Uk/t29GzkFdSt
63WJX9yHzHorb+W7UL8XLnfRfKfufC2AGA3MFzVkMlEthKz6zNBgB913KDUkDZxL
VWCAp6qOHhzl08d20WsKNVsxRV+8mQpx0qD4cwO4UqY4zEvrMdaZbTJtjFE4AFMM
Ifyo7lL833Y44IJZJaV5iFYHjanCbHWzduxu+4vYK9/TR6y9q8OMDGqdHNv48G7+
nOCz+8yzL1QDGQQOjHoYyb/FeuvLrPwsdBw8gJ3lDqo/gB84pS3aisx80XItXa5R
M66WXPmNjGJ0Em9Gmb3WYnNCnfvpxjvwFHQf+p45CT44mjGCpO0rbE+awJ0W40IY
s9vMFnuzPUfIiCD0tvdi4nATQoJ1YRElc55QldBytt2SF4DooT7WwOIDA0mNVfl4
stjMydV+I7Ab3Tc1g3aF1PBGkARqBzvy+/ywmn+y4e0nEkkgM0ttZURQ6t3eGrYO
1da2MhBcpJ+etU5rSa7tjaySy/dOnCSXohE7OLN5OQC2pcuER3Ira5Yk7rcM9DC1
k7fzEtx4hsgDjJOelAAkuMDFZiYidpX1PbtY5e8+8869hRzCGJBeuP0zi3dCM6/v
xDhpJAiKFAjWBx/+jYvc7P5RKNZGtpuqkumGHUpFKkf00Z4PkfI8G8+8uQJdoWrg
e/irEZxWpMiwrxfdNnb5AKd4/p4CSbK3ipaytyo5w/9T7q0ig9UglSKvrfhdfyhc
OEWmSAMygkWM8QHwuvRzLmDKtLjEt0YXbtrAbQoRwRRxHqsccZ3qGgocL07qzt5e
vq5U3GYZAhJSS51bg63g2GXUyq2Z+RByDPX+/v4DC/R6ZsARwK5fG8XG4atl2FpK
P7NRt6gsrcJOOOMSpl/wxmlkUJLN20DWNMrq6FlcLGrr6fbxAygmnFU6d0xRLq9T
h2J3+FpBKd0Z8eV719bkfqKpNUON1FZvqO5UhgNuGekQOCv7oSnjTmFhsmD059AG
Gqn41zMrFr2mf9cA/C2wkIO4WhF1QYqAfMnMimJvVLFcoyxtoKRat8jcKGA5xIyq
lzzRhGlLHzmSh+j/MMNysBhIsSCktKDLmvH9PjvMkcEpy9JaYrQWBZuiQL3/5iEo
OvTMATUaMrwCiUVu5AmNIhwssDe1CUERsC/CHIJlQ3iJilIDSAQGVdXP5mzXyCh9
qXlgV0Mr1M+kU4eCLdgamibpQQeVvCKGnJrO+B5P3rKecyQicvwmQHuNFea7iQV+
NnY2OabCA/is+r/awtBMyOAj0Obp/ZrlQIbXtiG9CTnwXXqgESHgZZeVU1lYsx91
9j3tGf0ft/UJp24rgpsG26hlXj/Tvx+cdgEqZvlelBb/i5m5gUF2ZNNYgeTN1xq1
MbNJWN0zpJkDTCRlpBzf7odL35H1drAzK/hcmyex+DzC7uXfj2dBYvbMl52Mmqdy
J8k9Nw5Qtn0g9rCUxANlQugRdWr9W0nLuPqz1UmWB+Wmhi44to72C1lOU2OwTnYd
WmpXTuayhd8REcLxMjaitFEnx8gYo1Yj+E9nfGyZkl5R9pvjx8prUIZfJfZtRPPL
HvMLQqbAGtUkFWdA/51AAgMHqqaXazLJzNn4nvF5P8icLwCCiBFhS2m0VDjbk1Rj
Rn/Wqj7BjMSeM56xzQMawNcTSkyqZ39LFkrOM47Wzpko1jztqnVcGc1wnGJfjq/j
Wnz7vuYd1Akp4p4QTch2B23ZVlR5zq19hUZpOfrgJFlZTi/s216oHPteA3gCd9LX
LFwqFjN9J925baLbM/yk0gzt9SiJzR+GQq9NJvmvefofsx6/ID1YQOyBXID96wUx
6LPEnosCvQUn/zsnaZBq0cm3c/vd45jPNlBrmw7kejECHkoLf1S7AYR9Vp2qo+i4
raa/TUM+sly8hslPsCHoT9mSnLswVFHyCiG+IC0KrD011ko9ZObJYjQKwCvfXQ64
s37N/hpfvKZzy4w9BoBC2z2WmYaeEgXQ/KUWqT6b20hmR4depwwVqohTKvVJrNEj
yAdiRFthSZjHkxeWG46hMvqRryW2uov+CTaxImnbJSdDHjb+CsXuoeL36imtZX31
YtMv3chlM8KyI9b5YH0Fm0WgczDtJ4Xum0rrSzvP4O9Aobmdr4IDv/BhZEGlHpGo
J5BmfnG+r7YO4N/07Gl5pif9BpU+VUA2qMFVCNw70dNc+K8VS/OmEQMcv3+JfdfO
O1XMmNO3Zo3AAOzzn3ZOv/dePpM+nIAH+5vB7hfSlIPQEZtPCrmoY7lcQ0FY4wdr
9YiBPBV1FI8StaUd4EZzBmH7SOXoClZknvejzlHuvT3VGbmKqqmFXDDSCwg4iprU
KKu01iB2xiFFivqvR+9z9PlkYzS8TqO++z1RkGTSyctsYegh/79+uxsNOK8gdqGX
ZBkdsVTsnGsMDXuTTWaWtZwuB109SQhEiLaFExNOhcK1kygnKZBeeMQeeEBJhrvl
TbZPdxcsdiQS3csG0wu6OnN2iUROiLBAMH4G9CSnhW/VO2GpAY00UqSta4m6fmQ0
QbCpqsD3YN+FvSghYRkn18j198l23ZzzjbTXta9Xmck8EbtiatZmR4IUO4ZOeWIB
gDNtnlkezVfgb6K80IbWm2QF0peYRM1+9EwQKHZTv57B2M4wGvW7UZCM178aFvam
3HO0lRdLeA5g7QQsn9wlqxsdUgmTDjTRM3JCdCtchvvwRwKyGp4pcpkK/PUFv8Un
xW8wAhi7Wqlxcj3ZmMJUI2TpEqpEyHGbFjwvdQ2ffDYBbt6Q/7mEDjX2fR+u86pf
AGMTCBjJ2w8nzO0YjauHk+CF1bFsaQeRhfZaungpowudihtpvOXUmA9na1xSYiwI
Hoxg6v2QdlsYLCbgNjVBpaG3f+NXjNgv5M8sNOityyxoeVR2eYH4Coef7g/Mr1vu
tlRCoclh4/FM12lxSPYHneyfr0koAoaXh3M9NeVo3o+ysLWHhSZ0HvRbzPjmyIcV
+P2MyBdzM3MWtZGwF789woWqeWIZcnVsCj7k1d8V5B0cW3nQoW5iPfKTJPyu0oJZ
b/qHUoKjhdxY8QW155ZDQI4vrr+Syj3/CqMtfqm7ANqDBzvH6mS7clAkxYFEKfZG
zww5xzZaCHsGFBNq/rXo3fyE0jtJ3mCFaE+9oGyqUU70KO6ecZ204ZHCot97o+xD
p8/ysi0twl1XpkvTTUBkN1K3atS2m55K+nSwrFplklrpo8kREvFqsWR9yQBm0Eqo
hfhrQ+OyKq3Qe2hukLkn/HXtTofVUo9D3IXSV1gZh5LviSsaEAj8HzVF1/sFkNxE
28KFZKVu1mRrpwqfY5wSrXU9BWn8jS4v7fdGrBL9KbXebqd7R2vudHtiyYOH+LKa
MnszGqbHQs0ABcATobjohPavaLTOEET1p3398+pO6i2feIyW3tsfQ1hyK0tIE2UD
iq5yku8qAQKwRfStbLJ/NkL0tHkPEllU7HwiMGoowzO6kTGDn2fsb8q5IFurT65+
CCGW4fZaou7eFjeSaH7MKdKsyM5R7+wTDbuYf1H4T3A+OLnLmcXieku0+hs3juNq
Q3sheiuzDq6IgGCdodt9ZxkKDX36IOsLDyKYUthw2p90tG+Uf57HAOYP4aaGLHaa
OwIjJ7XptV68KoXpdMMxa69hR+rx0s4uBGaiNeGnmw8CpYKX8Hbn0fyI8Y4bgP59
nT4+rh3209bpyDsoSzIHa0SEPm58K1r942bWgUVaaQ23PoZsomxLkQPMx4p1qEjF
kWUkZ7yAPkcYTHIOEAWxbtsfbQb+Dz0CP2a8XiMQTtCsdoEEU43hlRW4P0Gdevmn
RUOb2SdH/M/J4NwI6E9pnhBZGerwLJtgfY3qq7bjueGmOtDL0XFScx3/zRIq5rpD
nOfRpkNvU7xBcwtO3yE8TnRUaP46UL0kLGVFPEOvMTFn7kaIeulslfVTg6DWn904
Xcu1arrSddxbuw39dnZG7EnSdpIUwjfIXDU45Fmbk7lm1U1FOFdcWqXC+HB4eMgL
N6dOiPO1piOfE5SCR70G+tewFrtS+CQ5MsQLgi8kZTOURP9piKc7YtHRoDdKeZfe
Nbsa7yuIO+O6BtIAWWOKhuC1Ek/6VGQmEHSjbatMhtPEjUEarrrzT5uMt4ZqhPzB
+ua6emBlaIhQngXdgZOHEDQ4Z0GggjAEu/biFgeabM2EPYRLhlTShzrX1Spsr74a
nOd0XJX6TbpV1BHMgiBF8fVgdliqjNqIC6TvYHOR3pCgbBAAdTQeAveARvlDp9fu
obTwtcNzS3cRB2GQWEuR33ZAirte7PmUTb5ffEITdond8n0u15HIFlaJgzHgzxS9
8S2cvb0r8k31PQMgnJCqGAj9btCAsRTrEf7NdVKE6GZSwH6A7BXq9/7Z32djHsfA
AscSBkjEf/V8tu/I0euVthi1cU8sCEZuh2QM3Ck4mEILryhA0+c/wXSKaamqP/UM
Y3OWAjrveNJXZ+QC3UknWhax5OM3MyZXPjoi8mp3hH5SjH++vedTiSwYGG1upcAe
GY4nfX/NUe4OmG1CRunXoQW3h0M/gbxnzesg0Dzvru8k4WlU6hWyI0txBLgzYS2q
K50GId4gT0TXg6k4n4BmbDZD5VdwTWER7hFM6y+yVLAmUrzlLBNl4Gmz/pi+n5D2
I0py8t7sMKXkYzwyUINKU1kIaeAGLx0BvuSx8egsl6ldWRHdTmwZHXZz08n314SU
RCP2cjfXTd1lfXcJ/aMjxi/CwErHpU2SagrVl4pL3MKoBE4KrCzTjXEU2loGNawW
EVyDmMFcjK3nKSLWaYk0yqPsof58Bt6wP6gEeXA8Kf9SkRCB3cmlgaNz0cu7SDHI
vPr48hShrHFomPAwbKM7Lw5okIdw4g1CmKRhWthKJKujcdOZbAr/Rcgc97Q8CDYt
tTmP3DQYtIwogdF2hb+AVdHmv2EaqlDUZsHwlDcJZwNgh69Q6UHmoqUo3EqX6Jbz
5ZRRjicaZzMwiGiRuvFepG+VLvyh39B6RsGX9gRrDV0pQcZoxYj1d2ktBxiTjt4m
GK3jNyWf3sbFYBe0rUePCZFR2Ze1omydi+MImRGjvPEm/CvNsyIUFO1I8pkJR8nf
F+IyN1L5aOH1/eZ07yQIa/rXh0KiVi7WKYQXliGfBmc1niPz28Ra3/sHsa8fPb9m
HHt44rjSxDsVdFSt0sc0PtpTtdBG9NlZNhb97VUeBBdWvpcRoqBlgESyZLbV+iGB
ld/XNN4BRX8qkzXGiBrzwImw/SSHtO+y6AvBvEjX+sP6x4iXKjrwnNQGtOu3rKel
UQP+To7WEaI1+rB6vX6+cjJoQSoaKAtb1NAcgJIDpzrky+Z3mYFI6oq6AMHJUUsw
MaGdvFKkuWcwVoT6U66EnebHSNgMNFCqn59qglToJy0J9uFTDNAblyqIjgNgXEKB
THVXrYlUJSw8mJQ7ap0AruKCcZ+5zMc5/UcoHQJsZPMmRiuT1YI9MBW1W5eIfUxa
yvNcZ0SDi6A7fUEPsXgvB/qGwiTFmanrTqd1SC9YCjrM5eZydw7sle/zxNUKhTbU
++18mSwIyHD595J1+nNHn2qmTEnFEspcEnykF/beD4AoSal77aeC6PZQJ7ewPVhC
mrd7wW2QEQxZ86OawFuVIt16QaVtURnTpz0RAfVvXObjQcJSksE65A9AlvFTeojk
CkB9RRCo37Le8rKhIX9WcZgen4fU5N0M7nGnsaL+2hvooHUQIfLz0cq5cQZy28eU
sMFFd4hNZApaE1Wla30p4H8/lvFKK/NJ/k9MK9GTpjgPs2zocUHktoDJfhUTbQLF
TmS1MUXoUMvo/0eZum2I2BtoDVSuLbx6NHdckzprDsE7mk5JNdghJ2AHv6fWQmZe
639N68/iX8lYMwt6sgi8rmvB8kSiGUGIXw2H+Vq/Oa9R18TKlSVsgkNumjlRx2+4
jj3MsuEwYhJ+N/kycehl9e+u1s6hESa5Om1ZLdeG+LTNBzCWXkMjm7r9MT1QwW8c
X8eJb+nVIyfBg0cGfC/7idC5VJef6LGFB8X7gpfVcC7102MFg5Wx07pV7V+SyHXC
hgAKuLcSQED2K+gb4Gx9xDIEKlseq5VGKCrzhqruB6dlbMqwqd5SDGq2PE9XDENS
Hc0pB/DJsDuXdikMwwEyED9PuC6ImOPHnXNKX4QXuMMH2jo1cOtvFcDpmdrHZlIF
RO47ahKMQJ+kjj9jPDBeglpPn5UmU4FvOTV4rngpyzwOszKy6abT5By5NE7Fvpco
n3mjvQVDfDqN2CGOUUcnRFVGRYYLles8arfLmfyZy4hD3IGuGomhvjhi2uHkN2aL
sOWstv8hgkU0EoZh+onzn24daN+lXCjs8wdbmnjfh/tcT4m0vZews7BLq6qKzZPN
7ole8+5pA62DvXfKE085FVff/z4kI+tQ9ZeZd1Il/TOC7jytpL1NlK+INTviCJaS
MVP8QewYmaQO/3/OLL3aECR1jQCYkVEMkahOemS9vTGuUC9JbFa9YLQheZuuJ1L+
hEaMmHw3ZW86rtl5C9n0pHo8/Dnb6HS8RIdrFMNS/V3e/pPz3dzXk2PNTpt1yOjN
ETrNxqEL0JSw2qFUYBtB/cbg1pJRPq+NLhEim1xGuSrkrTxPJNNuq5lezjE3l//h
ifYuD6wWXEmXJVne3sgU77hKlotanNIMLkkLj722p7RjUjmIy4eK+valTgzlWeDN
NbPxKQ+hE0CvRIvmLgNzTzSTXED/VeRzK4r2v5d2s9k9brxt9K7CEGXbC7jRTAzV
fhyUuKNRj57sQNxwfKKIStVuz8PjZvLcVoJzvE6Xes3lZi7nnUNlF27OZoxsq7v8
wU1vYqDqJT/4qlB0/Q/zRYL7VHiKHl6ayom+WOy1pGam5z/qv9jLodcWuWFPvi0F
PnBtexcjUngjCqYEftcaxZFzeoqz6a5DwCvadmpmnaqQytGgLB4a+4dGsQWBkThD
YzkIj6kWF/5wAog2IjL18GwdTooGcxWnSNDQxr9IaHIFxsc1RxvccP6mlQKiJ3Kb
xwInx9SzozV3p0QNN6aKHyPeEw6pbmeA5x/Ks0mhK64p4oC8xKAqqwlxqA1SyCuP
zGIWnH9Vk6wbwMotpcKfRq2PnVVgfP4v8MbP6jKmbHstxFvh92aOoKxYoSbGnybp
2aPMUzJWwwAVGhkheNKKsJU4w5XrSxnswD7vYJoD3kqraog2qjTn8W+pNeOGrGBq
a5ET+KNGKJsuKY2uX/+yc5r5ywMJ2dTPI7zcgJZvYX1dkhCXEeg2dnAYgsUqmY50
7Rq+UNMgfVBWcgIs1gh3J1XZv94Hsei2rVOjeM4Cocjbh0RCmThp7pYv27zgG3JS
wRgaGjj4Syh5kxC0qCCTth8Av2M146iHA+24awTAwQHtLkg+GEZ+8XBxZbNo0Wn8
qES7JDadrC6IXtlKzV09Bwcm3iNQZLDitGFH7nsQv92ML5kEPZ44uvOmamc3KcT8
/g44gEX7xwf4TxZh+den70N53L2VFMuu4+9gW9v31LcHbdyKOhin7ygHZVnSt58c
VAmeZLJaqlVt9RbFceR10uQdWGfGdabefYurAc+qFvXaEBGCdQdyLnwrkuFBe9D8
SI6YxGfGvii9kV6TC0pRBKZ7Ue/CKTAAQHQwKcVzzxklx2I96woZ7PvH2yAA8sbx
9p4qDC7HJhxbcmbiCLp7GenZWG5uYoSBxk142TgDp++zEPcpo9GzIfnz0TWmgBrm
ptvbsY2In6I+wEE6LEDvPHs0baejAvg/M4FDManbmLLZyAx8S6mGpKTLDiXjfaU4
htFgVdUc9FoAp5+gdRCFeID8XIPbssNBE5jNm7fDKdrXBh7hJW2u58fYMl+6wEMQ
4nCkI9EHIiZvndI6qL9Frfxb/+oNJcB/GC3hVtFrLN5sGjICQkaZxg2HKgCcbh3m
mI0w0pQcQbDTcyhKfDsOrAdwxX/lNI7/d4g9tpSNUOSXHO2TvYmWRmkylXjKCZ+C
jXVc328MbZ+wfAQtnD/55OTT4qVNO9lZ1lJtpHzNXTh0VGnNBTvpDKQMxGPr2sg/
6Ay1Dm5PAwrcTd7ynRwK9IXcnKb74VQJqoF2TzE+VGtWVbxeKRkqyPbthNObrU/P
Fwd4GyfbEidg0sskNvbJBvlsvdu7rsfjFVk2InpyV4kOubDKR3x/iQwlhpsjDgdm
au4SUjhJn+E9jk0LDTFhbA2u0JndyN0BAzVc3pTqKy+L5KGO+ar96hyJseEyjWKb
gjzsf6RCs9S8Rjs/RprofrwAtXZ/k1+iHmN4QNrYyVGZPg1Cun0dg1UvA/ezcVB+
WULWJZIHqq1y96VAefWcYiqk8Fg+BiH1kT3ptVziBtlybGI4NLGshp03Y8ivEyel
77Z1NtpewsLpcIAPms8O19LIYsy+CqRwM8MIBgEz6vteJ+g8E85jQ9PUR83gr2bx
TlHfUAxk45H2Usbjam57v+uMxSe2aEij6mHnP4VM1kMoShaRMgDO4R/lpR+1drgF
VfDZJAcqZgDNB/bSVT4lO+PcsLBWVeFTEwvdts1+KhVbkRllo4KA7YUvXvbsZqYX
/iMm6OGNZeLNohteGVojK5QmSf9rn/NJRfLWqopBFujW3p+jmD8wlKDBVi2+3/cF
3eFDgJhjS3fXRJrriJeVy/DJrrslxS87TX1YHfdlCxdOxEKmi9dRybamo/2vfffI
/51R5uOHkjSxFgkhKbcJFx8achzFaDqmCjIose1dMzEZaidCIKiunUMVQ6EAcLJw
y58O2nvVHBg7/h0wj39rO8PrSyIPhBSkouIET5rVyCalLknv35bCpZctJ10PbwHr
AOqapyo7Zj2Do8i3ZifxIoHYkwwme6v2rMtPZj0vn0Rdj0LphiRTp37zIznn+j9q
XoyvEbrevPL/ic+QbA5SrC2iF1Wxt0+ymkxGKaru4LVHpFQ6BXkFgfvO5EzC5eaw
A4sJsQPOeedP3POR/efNMMQskIXBSsLJ+asXpYOp3amTTQLyWPg1KheyvhZWeA1R
T2Qg7eNwC+q32IpHxett4j2WzMUPcd4yBEA1mjMmhRjUV6JH8aW/CBorjvb8quH7
t3xvw4NfxrZm5bhIBEtyYQbRAVP11jL8QQclLELtVlXNmDD0dqONSTT8E08duUh+
lBNgZQbNcBXp+7Tyf7TJzRkgrXCkVC0DA7WR58majax4Z9JLJZRz1iw4FrbN8nXk
SWyixIjJibnZa3s9wuXUpTrd/KUWUBj+mhBGheWnETQQLkC9ruErvnij8486v0EB
BdrlEN2z5Osryqbb4Xuy5eePQlJHR/l4lX1dIC+4SyePp+vNnvu8TPrPleUIz++g
aoN+K5v8xLtOyGdvZ2yeFavh/Ah4kfzq5YitbpGKjvmr3QjGpabifcJ3JxeRuMyV
0wcAnSqz/dJOE2Us0BLcZt2jbVuGZV4CCXV7tCikA5J27nzrxitNOgsBdMV4b/iQ
8t0lbKszYQRksIS5o7GAxgbQ6WF6zsadFPVb5cKycAQUnt0czp+RRIzjhBrzEkK8
SxetqeVgxHBwj7TjrWQkv3yTdM9PXBFXPsX8+LDE6T3rJzmXnYw199FDdWW78TcP
MTIroOXhyZpplERYE8uJBwmQ2TVBXQvarIMoBvvll5ghEtyYyjjoGA9n/fIb+GYr
hxTfpKGLIkz6UQIkjC0Zfr55JAvxGAiXv5Eb/W96rXCkhvHZizehLFrJSemIJeVi
lXRKaNYm/uf6I+1FFnfPn7iJQZX95WjwuTY2b9d+d3fF8VpE4y4G7eh2fIFws1Yf
F7SVZl1FpTOYQbutHzyyz3bs5Hc4nVrUeFKkYGLooWusKQvi7a1Q5CX9MwVdTbRq
6OF/o5oeCsqnN4Q53rPUG+u5di5rM8ig36eDaipSvRwL9vcyuzPv+hHhgMcJBtJm
Ut4gGhGOThzQev3v3yD3dGqcUyQ+jKDCQxrB2NB8jjI8eErxx/cvCnMgCpQTy4Vr
CWTQgSfY7ZcdJhqrOrMd+hUjiIXVhCKMeW8fPkLC0NHgJ9Wzmj85Z1r3wd6Ma5IH
xkjf5BlboU5c2fGBdmVhRA5PSI6oLaMaX3KKNHrJtcJyEfTqnXF6ekoWBkZ5sdxs
QZgPN7Ivgit6rtTIBHLnUY3WMd0RidkCeY+3k14DEJp0+uz/ftYyoTpxE8ftQfLE
CL61kES/44n6yQLtO0mcnTZpaauuqeoVavMmK0FTVGmKvrD/j4E5JLPEFPdXUdFE
IeTXJq1xwUYetYb0SdS/Uy8lxpSUhI364X0n6yRBKoeZSZEnJvDUIs8A+Rr7NmRW
FAjlgrHJd2/Ayq9g5N5ziVZ0TzWXyehGZzbwU7fE4oAeoPOwyMmURB5ZilSgbD8X
7XrYlNgqhHcoYvTuKeatLgx6B4fdaEaZ2zQ7VWIejGJi0DEBqU9MX+hq2n2Nt/hY
Kh4QTqnrhUlWyHGTtkoCKV7tJhR2WumBwMr2cMIjXwZFf+DgdD/UOs/GTnsC8WJk
U99rx0iMtOw5FoXE8R4E2Rno72gGVnzCRt1ofINc9jsnJ2aU/MhbGaQSErE0Q+32
6Mwnfgq7/qTf+dPaxYTLMigF7DjbrUEGoCGe3TQ7jvX5V6+m8QVOgrWdeMB+rI1j
RC4T09zQPARW6m+XrPhi0cFmZ8cn4QPbnJ9XYHlQoz7fzH1O8DGDcDHfsancY1DW
vC7PZ3QkWK+U1QO160D0y0RD0CZrfuFIo9K4qnwr2Uz3ojjUcUYrHQN0FpxcIREp
vmWDz9YPdaDs4OzCgKIhZy9zHnByTpar3ViTPffH39Ma0gMfVmonZfiu3YoenFsW
v5Z9SpTzxFJL3lCPPwvISo1h/ZRcmI6hHcZqbvTCYRHhxEo9QvbYsGNGAi8sY7WL
p8f7b9QTkB+h1xgBkVlSKdjiAp7I8KDQUxDdFINRGUlU/Pymoa284Jjcpo5xtdmv
eDQu6/63HsC1KND8QxTTtX6+kIs6Tj/k1qL0QwgPOd3vmGP2Sa8o4wqZmDHog5SP
8xVBhkbEkC935j/N3lAxVVdh/jwTIzSu2/5RVHEHrObSQK/1a/RII0UwybttZGrm
ptXg/tbdR9Dsk1zMnKVUmuPLdE++UWoFAO6mA1Jw9beBKIrLm/uYCmeA2b6VN8c0
Vn7OPbJDIM2fuphfzoUezJ1QwKt/HM7NV+BJjzmgHHCgArpTKYSfE+6KxUiVp31H
6QAfBFRYEQoGlbXpuwhFobfUZVA/12YX2BNBsVGHEA0DiMUQ/+YK8nLSmj0GZYDE
xkyQ9x2NlyxPzw9oeTYVJxEdyGyIyWIWiLTFMLGbK9BYNqhbjxoy+aNPsJHIpiW7
2UBRgdRQ5O1q32jgH0EymQ3L8JXF3bs/X3Uk2H2axWBqPN5ctYeWm7euFMkAjFHf
nzhZPgNbqZ5YbmdWphIpzOWaSukxnsvYB37Z21+4B3i0NPraVQWF0JRZAO2pPSrP
6pxGm0YmareRTa0YXAioX0F7/xRJHEIdIWLik8iPTeqen3OahHH5waEnZBdBs53b
ZicBemKPrcz0o8G6Ev6wpagKx6kEryAUjQGqHVBRipLBrm4Lh4rGvNp4BjnehYYz
/VOVFBH3E64xBKMwgiDVwX6CPsQ0rUZQUBOOA0uJlxFerW0YYpxXLiv2umQBSvjy
P3C13uoRLEgQtmP5UzaAOvsyLsL6PgRc5PWcTKTwefRP2lQ/Keq9xraUiC7X4K/O
8MC6o3BcIHIT3VnxbtfURTmNXpcNULwAu5sL0qJ+vwr5JRuY6JMnt6z4d09tR32L
IU7EIvYnV15ZXHMDWeW4YNF27mz7ZEQ2pAtQn1vnlr/X6RX8c+xHHQ0vrg714g6j
w5qp6CFdbvBClJSxhRb4jGWPMAyQndcc5/tE1hAHeFC2FTRe0+3RnrfYFvNfoKYq
WVfo8PxG2faGuu7cBmaUTEUlH4onw6oJli6oEptDFsNscV35CMrgxOTfhqEtJ0pO
L0OfrlHl2X0pQ14bPJuZBnpUaQ9kLNvbH1t2OKtyY8KW+sf8PCZaU5zraVfqqQU0
INuG+/yv/AHD/S4jeTkwMtTCFIkDLFpCtI6cfxLx3DQnzu2ZEzP1EV2eEtatr2S6
rGtv1GZXjnyZfquOFA4lQdRTMOZnKfHSSjbvqpDqQYf9GtDC7BjNiueMG9U8xlf/
DQAwBbie9B3+LV7S6/0UgcLAHh6AcA6kjbVvcQwIBPJ2K7xcJ5GgztR6B2DuIcjx
o87AnhCSEWFBiILGcbEHm+oI5KxFttRj96qetFKY4HgFk4TXaUFArmF7t+3IdFXo
+S094PaDpDYrsGIUIfzdWIjKh8p3mNic0nzbD8GJ1A99Qu3P4oZ2aPrZ+UNGP78F
xjoNAMK9ScYDpdXaqHgp9rRJJ+ePXd+o0Z1SwlYrg3aaoUQ2eYrUyTwOhtD/wVdM
JHCq0F62wCf3pNUYxZxiiMl/gLGibLEXzOHEZVZpu+2L6lr0/4wkaSD6SxcBaXhO
B+5HdqzZexgi0ehtajOtbxJjq2+Zi/gu8S5OrwaQlm8OlD5zMD8mecjwJGez7nuh
YvXU5BmCDU4E3ZNdffg5IWkihYnqSFXu7cvjT5vw0rvY25AWf2FkF2KQfBJArvb9
kPlYeyZVtAW56ILw41ywnjOWH3nDoE+tEnC849xN+f7tGr7ghPDVa+0GTjvyUnzh
l6AiydkbghfKgfZzK3950F0Fmvx4eYJyZVo37T4KuklNMLN1ie2McV+U8o2mwmWA
Ds8x1xGooFqsB3n7lwFsAq1QG96Y5Pfae+7PlRb0/yIetIlnNX157i44NLl40IZw
fA3y8sbHMCsWsNwqLQ6HpNRoylQsa0hFqnO/GxADJml8GYs333KGsNsSw669TsQ6
8vTx4UoEmK90T9DK6ZJ2xvUTi2QxTVN9gLA+LiR4rij45zb4JhvJom1LeHpLxF7p
Z6ikwswc7U4XapE/C1EsI9v5nkUTkOLMeTyAJrAxknVc+BP+JNRmPEJ9TKy/m0/3
6d9m4Dn7lt7TxNUQU8TtUtWmVBVUaegE7wxyNtoUHFZgXXsi8Je8DEdg6nkQbEfo
7AdzdzgJn2u5g99Ry+DDU1UZzTIwvWDXKKsjAmXL4NCHPCkAlMVJ/Fobw3KEtH/h
1pI3mr7THNK41GeMC9NT2rSNmVxfqD1jb5zMk9p1gMSJopNEnSwGu4kr8Ran/Q84
BfOl4alr4brO8imnJWI6q5KZ6KfU1YUC0E+s7NcXfLUI1NpIN1ld4c03vS1GXmtM
L7jEuxMhUT6qMrMzPvnUxc/N5C1AwxYD2ZYS9R+3L/E/nXVp6T9G/WnmVfzCVR5t
72Q5CKCf4b5++0X0hcJ7DBgIkPhaUTolxIAC/G3UzIpPv/zaomgHMapzahEkyYZ1
sNtN4/2ZoWWeuH7EMxGtjUQzSxTrx68w36D6wEHYAzkihhnbO0TrCQr6ZV5MRBbu
JDM6TfV/O/NlEPBqmf+WgSK/L07ENpUoXJIM71+Xa5n7aXfSRc6za/MkVKcwqLU4
NzlxBTC92glTf2wx3a7R1e9xbniDtZ38V/NOzgqL2pb+V6k8VL+1WFscv1alD0Cv
oO5m1TgpGNFP0yXQkq7ygwNizc3/IxmXgFfeWjyAlR52Aiue4BYQK16Ufv8HGhQT
v5VU+yc3yE9GxnYlmxzCeTx/IbCUkJpc3b0jffpTPSqfUVQcjqpceHKLHbV8AV9H
8STgJLVTy+zc4pbCnOtENnF6zTzEMELYQeBDdYDe15LFuNvgCf0RSeIFjFc5QtlP
OOlNjDuut5WbPCoJoEvMX26gOFY6/SIRkyfx/YT/ciE2ONt3T7mQ5NrEopNuC/55
0SfjxHrSbLqizgZ5GvsBiN9MIsmzYzCNUc/BM5XYN42bMDBjhJ6keLL5Al93xfpT
t9sWwokVh8uhZR2sl0a8Nte2RDFDmBoBJFvphqRU88xi4/bt0AX8IlkTGDTfLxaZ
xzQPeZq/S4EZ+eL/ekZO8DUGyyblfOe8ueG0PTpC9fUM7JYLJkw4laE6BAOnCKkH
tQIMUstC35n5Bx0UA4T6igsKtHuagDeWjpfNrqIewOL4qHgKrcRr7gwczeqD7cjn
A/7t7eP9jGfWQ53Esfpz2kbnDkZO5mLz25fccHvMM9UeYuXIJ2w4xFrNuV4iDDxG
btJhvvO7VakmrXAg4AaSWBQYId6nrkUr+VSDw/Ad3e2NF4Ox8X8fs3jI0Yyh275q
IPFVG83IuHogh4f9pf6O4EvIZY45/wlPsNI6RFNAPXD/4kKAVEI+ikdfSLbtCZsF
Y1umb298ATJ6LQlTPyJhPtyH36C0hfF+RS6b+N+49FisOWbKctIlB/p+qXo5U/tQ
mF0LRc04bt+YFkTkNYiAZMvbLKNXMn1CW3dILqBsm4805RiWpis/tkt5QixXTR54
Qm1K5z6Vtx5lXCjDcAwvT0+2B0tCLES6dTWDgHe57uPOtt3Ec0LDoh5euGZ7dxo2
BVXg/mxYU1wcs2yCKWvo3S7knQ6raIFsUymTo6KXozpz511+cG8quSYYlGgeQunO
YnCA/AFRYQwAuwnNbF/KPtxPGOT7kWr1+Fc6MKthrok91iAlKRiJwJE+THvt1E4v
ApJzxFboOLWgiaMb89BcD9lC8CU2fTFva8+LxYPrujRgAYCZCwFyTQNfdW+7YAGH
+w5D9EGXfhEcDNayak81iKOA5S/KTaF/9E/p8PclUCdqmToHk7ZVO0ZgPqHdxD1p
PkHgFys2608ASFYHdwLhbLX1AKUUOz8caDAcmBY9aGtz1DgJmPsatZAl5HXumpBc
nBd7rVvNP8Dw40Y7IgJtPB+r+GAUBtUqdUP/HGij7AHJluVUHUVzzR+XePjbySWv
nJ0V64qdN3P02IfUePhyFcUlylY2VzXwi5QqDze1l+NulacfLmInHR8k6DC4xbwM
6RZJrqXSGG+vCjIMPCs9bIAGrXQouOP8YuGXfTaopb+H24KMFzEKLE7b0o6elC5l
KwBmE8TjbAoMzLRnp29JX34UCawUjepHFpaRCv9RtWffLTHLWLjpT4R4Feku4WXU
O+84kRt9bRvsoK+/KpOxqG9mFKmsrxXAROPl4biE+t35TM62SXQox46ga6oi2e7S
EkbElyaxv5SG4hSCexea+360/RP5eBInLt6fM7ylc3M7vvn8UbK8hKpRuqpouUGR
uZXJ6w7XHxIHb1b3+uaimlWft1RFByxcZSPiKWufpzhkrATK86KGNZEiC4i6NwP7
L4L1MIGAo3kMRLACutzJK/mk71FjM/S5gD04bD9ZIOeYQ9M/2KqTWLYEO2O3MPbH
UvnC61ujjTzPbPDibR8niWGIfGUjNvyTjMMGuBH6QiG364HwKxm49PgFQZkzJumk
8Gy5GVy6fMWv23IDqguTetrb594kHIogv/zN/pCTl1gJEFQZNfZtkVSI3P0gMYyh
Ndlc4LhuJuOFBCen1ELms9isrhGa+P+J9tRyRibyuIDKwPUKBaaCLlBUlGJGpmaW
KOCseVGZUoJlNOCF73sDRuPl1zE+/Mvzk8a/o769i5Sx8U0O569deWabgPLeFwlM
m08ExwDf0s++BhJ9ulQd1bJNkB2gyMoY32k7vD/lD4acnsieU95dhz2W5zI93klr
LsUhp6UxuNWh9JlQFDVQRxCeyweNGlKV7zZqjz0iPwL1yu64frHN/ia0XPoYQcSA
B8mSi4antQu5REhsEVqYrYSY6p1B5VnavJW01htOaFwYL8kHmek6CMufxFme5VAG
IYE0o8mw+5iuehmIT5B1nP8pAUsShOAh1g8ngT/xSDMn0Waa6a2cyhXfnwDIeVKB
bOJLKETY3S1YzT9eIED+t/eeweUMMzF13t5faOZNpp1YU5jDYE2rKuSPWOcpePSg
Sa1VEsMpco8HKRstdDq07a/D/A8eDYbMzHThz93BI0udmmncfsrJ8cYXtaC3/Wnd
ZcA1v+/6Jg5dzPbe3kSURnappEmoSdji8yhir+Fmd314ZJqpmcVkJL6OyB++aiMG
gtlmrC7X7u2/jmaLLYPMq4+mzfDzHmbWvz6IbszqSAz2yjL+2rPSkQWDRvVsm52k
fyZ+lqsZdPNBuCRIC7OBEMsZulJ1xv7uja6FNprJsaWkwIxUhubertsvj4AEgY+g
I3AzIJJgDF2v4sai3YBiNUKY3ZO0Nh5XB5A7+RBkOOfd6zCddnn6FL2yYUSvgHw3
V+uA2Ut3e549T1PIjJdiQ504mDeBKblJZ272TdEY56QwlOLJ0sij3uAJvIwmw58K
BTyXDG7Uo2j8Cn+VbvWBPYKZQdcvYhocphSXExeV3mDGiYqTiKG4ZzXO5R07qLUF
RLrJk0Tqo2ChjXsdYpqf5x5FISVR6/z5HRqzsXqIfVw79Kfaq0L7BNjuNwUhT86I
EPOeRQYs85DhUVnl7E6uKdUyz38jgVslGqZQehfaD07yyx+bjplUP2NWEeloNxfL
LcyEYvbY3xhpydkJWgQrIRzTYd6cC/ClkaaBKeye01vhtSdRO95XNypIvkhxE9T2
0Nh1+Uuo5vK96q0II15tHxe03LjpKqNdxh7bcef9+SkCR05Iq4wU/m3mg+lKZC3F
OVmdGun0nzlO+4BX+gH/0KwHP7ehBqd2P+rD7JKxsnwUY1wuqnkStM49rMjq04RF
9Hb1nuUPD4jl/WLYD9fYxbrMm4iAD2qAIQFGCVC9fLiG/0xl7l/jTQYqYpZQkfEw
08boSvxqtqHuB0hegtoO/ipdk78R7NQKGlQIwqgZzTwmu/Ab3JeZ1qTW+8Yr/2YS
9ZaWKG0/sQc0SKuGyIOzj/KpTsL/U/9QkLNctMNvbjcOB310VLhK8It4nJBHtw2G
qc3Ft2Qbf6u1a/lSUuA+1gyyRGTQ1m2QV1gid2NaQRp3fPzXyKtKAk/hjSJ6twBO
0klIZ8dX8dv4lLYc+7xXlg+B/gPVFQ7IrKIi2zciubDccZmQYnlk6/Z9f+I2wNP0
odFyRCqm1KiEkeXzCKSH6+kX9tTxR1Zy+sgccjg7egz8Q34F54sdDolx58StBMLL
PUfbqu8fMc3Y+A1qllzYDzke+eeIB7Yo6amDT2ZxhWcPxtLEkpnFVDQIQ+fBXDTj
fJ4CfT5NY1IQF4JrwYxS5bhe7ehtX/b9UKgcaOJAu52sZWORjajzL5w9rxiOnOaA
KeJ7awLRPJ8M7ftJM9xdJAcJBC60jIrh3dI5bi7/V6NFxJy4zkODTLmeoiv1EK50
3a5Qf/21zgsbHdHSGm8g/m6C/+EJEUk7DlLIItdqmU03gPNG+rCwMBsGlXSQ9nth
L/GW2n4UZna0yuhhUUOUkD7AtFAoM1HmctBNRdUMyVMfvUmG0rTHr/U0imY9tCuu
OBDmqvU2KU1RFdG7joI2uDw3mS1AEP4lzDiNbpCBrxv8H0DHJXstt01fHl7py89B
NSyq5cOTghaaERCrPTFiYahsppF27IZlBLjMS569COmwbqS7L/y2pIYP1oOjOFsL
/p1v6ujhvFr/j8HCsm30F4s4taBpf1X4fsI1chIQ4bv0I8daQ62wGYCxVm9xDIme
Wc1efib4IC+VzeahFmYBtYc0uUVT6gVjL3Jv8ArrNm2PGktBJjPxdupfcMQAkK8g
QJAVQC93g6MVNoHiSoDe0IsEYv7VM0OnnOJfmcLDkR0K2jZk2NhTC2MNERX7L+xZ
+17v8+KoKa1NnZyfrqhAWObsANYdiN3tegMnu243DTFwRIHGn3QC/j+xoN8UkaaU
P7UGglWTgD0YiPI+AWQm7MC1WVLhnswmfdpAg0lb8bT/SpkT6tk8GiA0ZoYMRlm7
rZK6oA0sG5i4J5R1id7VRtJQigHty6ZSSp/uxZSYJu20MjJTak9l6qoP6qCGc9Ps
L00nI8SCenEd+/klVEK7NIJBq+TpbOpl3A5QWS2xTj3V9jmkN+C0wkotK9GcdWEj
egudPXR1ELeL/N9RNWQrDYVzMpsKb0ekEyJFwtST3EIVHbek76bOpKiIb1wkWw5i
JynT1ttLzbroqWWX6zTJ9ae2cwHZqAqttLHaaQLA1+EqVk9tFlgFVpkuI5iGFrmg
n9p9Goi/jKeKo6VygF7EV+9sac8b1dJTizsTmtH4VrsVe6k2pMFvEHTVgK8uySBH
ulquQqQfae8nyV6kco0KFhCg1xA5P7VL3gZEoJCOupZT4ZWQO2UnYU6If5l9wD37
ck4uDPaoX8dUvnzJdIG0/HE/RKx8OOfVLlodibRQ5lzHLcTf1d2EHiqlcbbn/ntw
GXNczQMz+Uio59Bo3TVCZsnUObjfCRkfcHW+Ehq+DjklfQcMNqCS727mjDBgNPzy
9g3Ausb50Fk3HUIWpT0rJBcGxjiOu2kEBet3mr/MICw=
`protect END_PROTECTED
