`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H5ajKHvTJVTbwZJ+0yoO9zv8M/BosTO7YOboXt2q5/AkllHvVJfZqYVzCzCYiWsA
XcwH30SppF+ZWhznKvpY5U2YgPHwIBxI06zqA1kPUuA7/7HJgX6pKilKNnyEGlYa
p3Oa3xsGmiM3CtF5HxMOW9HsAd/o83bXcKrknnmfX9YdLAhuXBEHnmpelWXlB+fu
+IacC41jsUmeGCal/T/7XinQiFUlHGDRBrNYUILlUH6aCWY3rcvX1WrhfVLfspaz
YqE88Uc0gQDQbp7wdDLnpc487l4ToMuCpPAT5zcBacxqLJlIpltwed5okxBkx8bd
2C3TqoJuY68nuX3SvV6voY3i/j+TS2cFo/YiHqnL0K6G7bXTyQmL8hAFe1z5Xf4l
1BoEwwp62wOa8UplHwUW3e0DN4/5tdxzndR7cyCNzBrFgdRtsiptqvH+InSyA2zY
xriWsaWjJU7JcEy5FEWDaKjSl65n3GHwrTU+MJkqTUf4CpD8iklk+/AtlsDZDXGQ
6ZONaJWVOKGPk8OtMRrGHuDkM9M4aLnVqrhbQFGNQHlllBzsWW8hrLUsvA74KRZL
wxPq6Cfncjx2nWaKy6N6ntogQdnaMDF3RjoyxkU5w2HTy8hrWGOqBLGPCcT2MqFP
ac7cuCVwYkMgWpEXwQqL+RLpR2nfHaMeddpzjFpNuL43Y/t8QuF9KZ2VEooliOe9
tPsA5zDQ+1IGX8+pZe5jdor7wd0Ub48PxX12gSFrEgz9gp7WPkP/d93uAP/xoaOf
OnIFLWVgtNESJxfdhkZGkrZCa5NMrw1qKSSKi5SDi5To34lR79R53Xu+2cZ1DV6m
2qjmVBH7EpyWLi6sAo80GXHP+vyt/tQmtDUD9MCYbwsFd0/jVtbHJ08bTqfwo5Go
cb7chhP4EAxLMu3KUBCa7VTWCq7z2nef1u1mJlXvQ79SQ9e1Ov4r4FDeNrXbYsHB
TxF+EDyTzgjcfN8LKURvJ4mQMjNxUro1GsIkLv8/G4X1VHKcszqYmFI0wpLNdfBz
tVgsWhjNZbS1YXTuFEGluIeDTe/jKPU3/G5OcnzAwhwM+k/PvWpxWIhDF4W/42g1
f+C5a1scMIs2R9b6jUGVjdJw8suuiIdsmGt51CFdmxvvAx1Bl7vnu6ouw+4bmwc7
GSqoHEnAcPrlTsAlWSvYwtIjK2KkzR6N1xpK3woMlYbXhRrsroVRXClYL6vtRAEG
MJ2UupZadI0szAx8JqTr6Eid7ZQc55jUIsht63TS0/LHTjdf27DnHPPrB4gazV6I
bxp0G0P6r69ja6GG7TLZSeY1DokMtDvKOatcUAfYiKPTbZLvIktlnWHUcOPxy8n6
JLtkP/7D35YEK97OeGOi5wVmLn3d9/g5K12zeiT4sto9B3UMjyXjN5kUc6KJLWBJ
HgIfpOjlDli4j9L/DUpipBwxaHmge7kRjGsLvdIOl2v3WjIZkRgBP3njvoWvVnee
w0TuplTQ0oiQoobQmnevG4TgHiiOekU3fg83mvDf69qrSbQv9f1rPmCrCXffix0b
NM27RTKJ5lKVBosCIhAHuTeJBu9cQ9H0PLzA6uBllE3ov04GndG6/1SWKlzWfaPV
fud6zMD0kEfWTUSNl/ypNvTLPiMwfl83XHvc3Xz6VQDg0r8rd8dwgDkPiXU7PXcE
tkwnG3Mj/AcXNX2G0ltXDLqxLr3nEJIHveB22LkN+STek0BrVhf0hkU33WEhoDYR
LuvEBmHZECNm6TqcUIAy7Nxt2e1mmMlMjjjU+mQXH76h57RPH6lbbN51WPdazwCA
R/n0ovNZcUhzWPHCGyZULvWbvMwvRrE6m0TrJ4sQ1+/CqiHzmg21E9SVUvouMWda
+k3+RZ7he2AOsCzB/O2/+sTx1H4N2lTmNKYY9L5aMlLuaNNE7nFXDafMiQIt+h+X
3csLPd945LTK0lqi0Ptkib6o+R0HlOY8Ia776a6TxZUhE6HOC2vF0KBBlwTm9kW1
rcjtaHtO9U4Ljbm2TAcY7xLmixZO3OWmHRElzL5Zr5EMF/DTsw1KuE0+Dab2CgJI
8gJonFURqV/+heHj+BRTlopCfXpwmNG1BQ4kyJD9w6xGjQxV6SCOArAUf5Fx7/N0
5D0eFsi9s4Fgm7ibgGUvS1GN+Vp7GNIzG/c4PZrbc35psbJ5IIW2+MwIOOvhdbf4
l4XwzsbAkhyK6NrCzvxPPw5D/r56m6D75ZJEs/koBTV3VaUDr/j2h8mBu/6BXo1A
zX2Uqzwo9UHx20af81KDLqmNOHHUCzPu8sHsRir0+JNoHznMd2ZQWlCwHKXSGe0H
J3xuZ719ojf7Sc6Vth0DADSFEh6ceI6ubep9v0Sg1XAJRISEAYuMqBkoPde8Zsh2
5lP+dY8eJK/D0Om2PkAPVlQyoipZuVQMz5LmrEOvpgY0/UFcrvntm6zqqaZDHUFQ
XHWJx2nVnoCQXKF6bCZO4sDYWoEE92g8wjcLuHP7OwGU7Ptena+aCdnlRZMEpHGo
I4j6ChVRylF7oG2A0MIUQuNpgADFP3arr1pwyIOrp5GlYgqpkRqCiwvN+ZUln79C
hEo7aXT3M98tynIg1BfatAsAsD0STX6pk27+Qd28q4sSQzst05hIZ95IoRsngDEK
zooWkShvBIi8qh34amyuIM7ArLGNDV6EBLKzz4D3oYJP6nUn2rnS9qI329mmn/ya
YLGzGQTu0GRYl2Bgs49FOpu8Cz/NduiEcZsabMEQTbT2AMEcHcrT7+ud4KTyxewt
fIaEUvFHRLfs84caGhQTEBxB/5C+i0Xt3nfm1wQrRQL9D4BCUKAaYkvA5fdtBuUX
nNs1/gl5ciGwyonVowmj8iJz8h+woonS15AshV3BMZXy8MnO9kF6BUnrNVie8SFH
2zpLq/EZgHzFTGNlQRyeyO+u32APskVwDNkBnhHqGkxXEQ6wtX5EHpgvpIb/l1/L
tSVI6U1pTmZu8RTqJSx8SdRkjQ1WcDfDUhFC9kNfzH+QpmvWy+t9oV3eRHCxWxMU
nwuOap09YwYlOcNw7VOEKRBrZCDuafZMFqR6L/KdH9Cxc6uQ6obM//CO0R3YWirt
3ns8DSLK+3734T3sS4Poo2+ybMYoexeEaX5me1Cx41kvvgOrDaHeku2iYGOK9fyv
DoEENCZfqBBdGxQf235fXimIBnCYxrMMBFwX1aUD5WL/C5CFA13Acj2C/ImSvIuf
ptMuWHsM1X1FJ6iWRuMoHocktuIygOkTulYqV2KYSR+XZPU0Rv3MMB59tD3Ng44f
YKEoPL9cPiIoubPb5L6qj5+m04K0tZjLjtNZJ2BcmDcdQdZ184l+5KWH8oDUogcI
2Fp76uzhCm9tFAJdaUTWD77ahONEOkqL3sAHKJBpjs0d5H/IpixsoUBqolIjsUX0
6dpYCqa96RQFaWn9WQY6A5a0eaS12oYYcsyz8u1N5PGPzc8FO1sA1yTe9/7f8BFy
8vzSUXdL1z8w7ZrD644smxPRuPaJeWHYpmH2iJmxvd4ZeDca7+0jMxU6yuDClZ3D
qBLLijUb7qyj1emFhnA3wjv2TEgWW+NnaiG5rVovGwhmdAiwKIKLpeEsL7D4P7nd
UzObY0zwIpzMAmWYFeM89kmUh8pJcTvia91i+YwCQIq241X0jxNynJaUxSmD+5En
RUCnlg5k1gZskWKkk8czjvGwf8H8IHC3J+tVGHmM2LfQTurDeCKlPWJVpNG4JcZl
ZITLETy/HY/IkmOIvX+EY/lr5T4EhqIEw664ShVS2UqCaEX0E+pBKg8Cs3k5tMRm
GoyC9R6vSK+tOWeqLx6d7qXmdycOjYwW93pLSxXRjXiivwnP+1pYInP/yM7CpHk5
irT2leTAiNhcqBuF/NdkVJOo92Hr6AQQLx9sI3gcP6QYEhGiPaoEcbKZj7byWbiL
Yl/7f7/I9xWV0HMexaNpzpxeWwWxnTJKT6gNh/Wf6PK/cakacqJ7fXhe5bjg7/sk
YxcL2d7vNGWLulO2098F4ZCpF7PlyCpF1+Oq1LNj5TbkXE4Fcxm7zQRI2qY6LKbB
8bnD9aNGNyWcssl/ZmTgjMgYRyG9RQ8tArXV2/GJ6ywBDkbMIF0QyF82DG8eEtL+
wSAonSkhKU6c87nxelgkoAA0coFWTyKMSpQ8fM0cq52InNO5bk75rXVLnnMOsTnF
NGcNp7YSuLkyppA5rGynm+jQbjMFzz3Dai0XnIuGbCYwM7FH88Nd7OAqgwtZKalO
4H2JE6Q7InhPgrNkXPKwieuWgXtP3U+ppwsJ9NktgDrWWO1Szp/DOpboNo/Ib+D8
V9AOZKunZIISm5bLkUSzePBldgQR6MgCC3lczTj8jFZTC33HOA/xNmhbwcJBQVf2
13ngZSZ706AXrgD8KUAEdNMPlgK2bT3q6B2Dq4tYzL2ZqPIAw9+aKJwK6gr/MAcy
EkcEHksi/xe1zMuC57iIcI+loUeBCw63N7/mgkkuHMXHmpBXsBLaEiJiFdcKPllI
68j02Hgz63k9nJZZAVZaD1bM+Rh5CBmFOvi/LXdmsJ/6tIMqh02NJZB2BTxl471R
ExIHCnWbYcmoZgw7FoswNuQjIx3HHg/rJLSPHL6BzX9bXL0xLja6fbVcbx2MQcVK
wJtNe1UM+lsLEJu4CFQVTNnPnp6SUTjB4jApl26M93U9m1VvPg9Lbx8XkRruoOz9
`protect END_PROTECTED
