`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UothPf0baMTSeFOZxo0Y19k3sPyJ5p9Av1E8rhuT5kxYKaiW2qrUcqid7A0OpPPc
r/7mJ7Wb3lo9f0uHAX3srGGWG9VxOyNeXikx4TgywZ2ycFbnPBQEAqqDJvMvYG7z
32t+IZs1F8OPjlaYuY6PmusYouqu1lCx3xT0lEKyWHwPELIIbJyCjRS9etn8mod7
PmMjpqcWOT4fm0IfcNUYJY/5nOnINbX6/PZjYwerbmrFftEtKayQWE8SxMQ+xni6
HxmpqjIaLEzrcAakkZQm49VIP7EBStMDRVdIXDXmpfE/T6GHE3Ir0zYoJj1et9R8
IOz67SO+XdCrIMee6fng5Y/1Q7ob9cV1C+dQLGS+IV6WF2lgsPT9B1t+Z8uxCQUb
qjuJlOypOf9P5+oVKo40g5VdRr6ekZVJI2WuYJ7BdMgDuQRq+bwcmz05JXo4Ci8D
so0ERwJdSIGDyLo4uEQ4G+n5psnDdfV6gKpcpjTbMBIHprfim6xXUhfk8ODz7ISE
cfEtDXQK1+cxmPQRwbME3Iv6g7bKsaEKFeeril51bh6y25PT3moFET1YnlowBqT5
DFeHnGYMll362bPOvR81y+0C8q+xaUHXy+Nas/t5quy54QmYbTAzLzvHXvRf+/zs
SDB69qNQwzElST2FRSC1gnbA3QWMrrbtj/973y0aQScqxSQntSSwIJC1dsxwWpFs
N0K4ZG+LW9+4vk1h7qEzJAYOFzoEb4aeOb8WLLaf9aDP0VraJpCPs+xiCVb1osxP
HEoPFRMsflGpHFH+OqlWAmz7etsIQt6+BIYcxQU7i1y2hVoRYbJQap0aQ48C9BpJ
fiO9mx0noB5G9iFxHK+kvUTM68v9Vj8XK/PH+OwQmK0WZcukcygYAfqxHOo7J48T
+uWusr8EL74XzRzA1LEzUZp1akzMI+oA9HI7hLztr/dPvbb1Qdc5TgtI+xBpGsus
p02I6+ZuU6v4QFxEqzax+X9i1nCicgT9wy7YdDEYTpQK4BEmq0vqV+GQwP8XHVy0
41glrRy3b3Cwl36b01fvEtJBKioGdtv/lyu00pccXjQ3/H3FNzncO2sfDS6GTgnl
+dyD/kB8tD/aQI4HXSK7AjnePWpg+VPf3Rwja0rwG1yNDJ7hXVLok0MtRD8lJ9Ch
6NRSWI8srDO5mxc2JY287H5L++5rW0vi/LHsi5sTxmanW+LQ3cBow9HPsu2KgMLp
cpJ9Cw0J33y6ObZvfd2V3ZeEixwlWQwN2ojKCBHQguJXzD6gIakDwMykmQ5YE8Og
Bf+fGvwWosvyCoqvNEaozQvRoQSdJjEha2vVJTLFxydmrvLDkNcu4Zx5GWw4E/of
Qd9Ef/0+sR3pJEDW+0kIQ1TAiZeQWoQCczsvy+RSEzzyHwKXYMzLMmRKXbdy/xPO
0IY4eoKTEVr92wUbUSgw3tQK/XtwXbcV6fNtNoxXJx1LRX7eBrsxFglw0RqVRkux
zV4H7Tg3ZpwC2c3kIPT81c6pcdjVtif8IJt2Y8dq6JXXtI6ip6yEs4Yweip2vWMn
Ki3wyjTbQzKpGW976lzy3NdrBbiD7RCm5v+D1SbzxPTzEr/bd6MzG17J40UDnDjI
FULuPBe+0jP7QJFbzv406zVnWvmSJ/dbsF60Bza+DAcG7yndllIA2zzSfn1+UISy
ZinXF0Ai6/zsOYrQJWOApTWNu9cvg8sGx+d/xRxrTCrLh4mvDTixt2ymIHghdZJB
muuKCfmrjsNro/wD3juJSkkG62iKGYxnKcuJTGfJSpfaC8sSeMnBkAFT3V1n8+tm
CyJC+1BJijsMYOULFqSCwKeXThq8aDrs0pe9DDp2M9w/NPkxCypIJe/+ORN5QI+v
Ud4Vg5GosRn6QK+RvTj0eLGjEmhBwLGW+2GiFQbsF11FAyZGisxdjoGd8Mri+F0y
ZBfDKWIZtA/rk6PPSQXmx0IeexWHW5QYAO4nbyEplAZOxHQQ4LFoqqGoghTWsYO2
PlwcAeNjuLLDZ9ewjvji6PqIpKdplI1HiYdzd++LaGaAndUujP/dQ6g/Nw1ppZ0i
`protect END_PROTECTED
