`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cLX1BzfsQzSnDesN+VA6tHtlJry3IiSrju5d/KOrn2I/yFyUzfOdyTFWVRBAVYy9
ei8Dg6kjI9Fsm14hYEqMh7k8k5nt+aqFWTImg4grXAMgI5ss6JLJpP+gZ0DjJPot
LjJSTAMdmZMtIet503PHLkAhn6RZ+f+Zhfli5SAt7GfL3KgSB80tODiykDZLtTVd
hCWq2ShfjC+OoY+DtFEizPpNtnJvPK3uwyT4pjilL0TCzeYXpiRum1D+KldZMC7S
cjoVkMKfS/3lQotdUXuLlcZ94wEBjmpcp8jzM3/b//0zznAQz5hU9XF+8eMd63g2
2mBaR42UX5RZRXWbzfiFiWoXXUv/JBVRpgHIhYiySSaOQLI7dxDtstD9Y/qcOntY
dUlo3PfQDF6Fp0CXzvXlvXQzbGZrU6yucU39L13leb6tL8CUOKqdq7igZ9xbVG6+
lL4N6D5eAPc7AKkmTO0/BjU4Ec8LZdZh1toxpDXRcAW7jc5GWxTTSwHB6eFPAM0j
QfFEgHkud/bIyHLuAav+SkQ3nZ+R9FBj3aqEdtnXwbU5SdaJlOFimGiQ1FNKjUcQ
ZOQQxwHVSFd0Qs7oNU/M2QmRDAxMK6Tm52tdjfydzIv037ED7bAEwv/yIZufDe24
gKZvRtTfPthAyFMg8uTTYW8AAd01ZqV7pLxeV6AhQCpRU5dAzAjOgJMK5L1z2wan
hp84DPyndPgXyHIIiRKZfTGMeYp02Pc2nUyAOKVza6vNpWq/Ny4T0hvBGWwQQl9D
A9pPN1Ir/FDWCpSXU9JvmMHlwXij2H42ffQq+6c964cV7SF4r9b3QFAmZJE3mrYo
KIEJCbtA2HssuIOWNr6V2alzQMUpER9CDf1OyZIk58Y3WdbxSkQ1M3FxmkiGUD9a
1Vk/M5TbZyFcXMFLJzlhW2v1EuPJjpttD6gUufDi7niAi6qy7leqpnDyNq0nWB7K
uhR7lYsc3AA4QexVYmSUGgc/m/v1ckLne5XQhikNEvV13mJ4okS1Lm5rDQWtDFRp
SI/yRfNExX9Yta/YtjgmdVvwGbD0QIVOwZCz+NE1NiyCaTs5L/uZur1O6NX6pQP5
t3uJoRbcHxwA9wnj09FWPlKZHPi2ZuvW6tq47b7Q9ALKFiGSvLUZK/U/f2mKAA70
uvpcovDPNglA4hbzAn7/UWOtWdFkmSKOZ442SmI8LfmXIEWMLElvJYIMwyrNrGVl
iN29zokKoaCan5bkKskh69SvkYRM7V3JAsw93K68brGGp9Rr3ZqDVTLmZXwDBSf2
jakigGUhvvMqdRx8ZeZhT2rVbQCizVqHaQFaPEj3Z8J4C4cjCSEmzgfZDSTIb3MT
qpYQ9+fmW3WRfGtsyms1n6Ksmvej5HhPoiaB9JHzB01/MQWG6s+b+AiQraAAyYzp
Twwm2RLNVw478ams3WrD4sTyn8kUCv8/1H03Oc+eThasw/reZfO/F+WHm3vQsjUa
2XgQyapf1pesw2GKlkmxRFOWydzML5dGK/Cjk2Qd81vMfZgdrq/MPo7GaN0XEjnh
uBD078X9pzO89JwkPClACIY2ss0WDMoCYFliI9swbs9KdyNnMJ0CiiGfHNynjWtQ
B3iAgY4K6jfDtCDhiiQQyABvtsfT6LTN4UmztlHNISlRmYfCBjNiB4ozN646vUQd
6n/IM9qUyNDKsv2V2e45kDipHlX/Fm/7a8HBDVeRNuk2+ygnyaBaZlaH7QpEJZyr
KVtNfycUjUlzNT79VbjMnwWoYOchCI8tXXZSndqL2MHeg1hV4nGqw/Xtf9jREuIv
CNCnQh718Mtict9qLeHUmiopotYQWt7Mdayp1ehmaGyrPlX+Nng/l+OdGAkDVgUx
3cgTQi7Vji8IzQfWnmXhvY9CU8A9vegX1Di3HS4PvM8IY92dv/osNcQoBtIAfZYt
ia6HvUXLjZ7FNetODsRLzWTQWm2PPcSuJ+FdZwP9Ufk12ZyZRz6zBQpYzYxdOUN7
Skhm53GwnHEwmJULigHkQ84XQrmSgLzjwlZtgIpsTYQhZUv4Aj1NNjrawNowd3gK
QtdoVimwotMwegaiGr9p+fpYGAzzuyrRev9MTzS4tTr0VNuVS772MlgWjSgglLbi
BcqlzmyariXqNwa4FZoSGx+iIAs2lsomCkAqDYJoyLjXeBI4i8x0yi9IWKKWiZA3
deyvOssdpiJ/e0TbOx6TY3qTPo2JQRJurvKdo8zuJBQ0H1leKxiNergJp4Trziau
iOqPHg2Jyp6QeBOQcBN129RTEUtYe2bLgNhOLCYf5qzkInYC/nYWiOEKJnE0vPzC
ROsPcl0bYl7SawhrjWZR93I4c/lnSa0sTcYGoFJNPXcHLklZvOxlBgMr2L1yRo/I
yEMZ+/5qM9wfWZnWLeRZZR9nRI9Eoy6z62hjSUVydaf07Gf1IoWcyPq1afAjJ1OT
dUV+cOq+v/560NCw2rb3AGy2aJkk59kPScKlRIDLrSUCqOPzIIXjCHmMkFP2tLdt
QB0bHeGAntTM5tuqZJQK6YzC23z88bipCX9R/h00U6W/1PoSZMpPD/kmGUWMPTaP
EQFEj3XNbBHt/DQ6C5VAWsOD+Rb+c2RDz2c+1Crc0ZBXqCvpz+5DMNJwMSlGeYdA
WOuMhJ9upoAEajl40QJvZ2j5lkJ7RWS3lIBzijZsd4OLh/ApJCDOO4HGuz7EUGXJ
NdfLLlTNXKYAl+74emwL4kTu61fJS0N6DwSEzO1qNk3rLElequEmrFUM6h6I/qJx
iB8AUpGzDQiZmxlyQDwwurKPbzrp6jePNJlBOEh34mXjkswUez0zl2HRQ3BLpKpC
7jtTwnP9KlZXWmeHq3cgU77IINlfJsF/JKZvnXohwBZUXsSyWWX7AcV13CrnVdEH
7ZbztTHGpgvXYnJyBTKAGHMG/IKG6xHP+ugP0PWFHjCd3MBSnLP2MTtffL71dM8j
+yftYTiVJ5kk/U3E0yaRI/FGd69Z39SEw2agh3rVzYd+lCMhLSEjO1R5LeTje2r5
IJagBXUhZ3rVzuFfROwns6iTZu5r4dVYocF+Y9GFHgmi8ecW4fr+ES/lMt5Y6Zyq
aHlZ1pNSXbK/QgjD+J/M/7jd0YKMHhEkpJpivYbtNnJySoX5H8AhoVNezsFs9Ws8
efoUj69A1GojY2RLx4AWctrD5UovgZWqfDJbFD1ONCLjTP4siZ8fQwQxv2Jbp8de
3S89q8HUxUNGCQ48sTlLUaXQzBoBn1u654PBQ60puUCD7EehcSaJZnwqlhUfZruZ
zG6mP8mRTHnNFgbdeWDGVwhFRE3Kaslvs7yQJoAFtyRfYsqgoEXoVVbtf3pqHLU8
xt2EuK3hTmJprsljULB6Gz0N8xPRsWOlLW8iD1hxxz9Vu07HQ9DyW6AWgKknnWzl
9KV3pycIDBTWgeZJ7rEE2w==
`protect END_PROTECTED
