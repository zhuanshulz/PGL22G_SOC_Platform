`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2tZECgMz6RVJtfbBHW7pYOZ9xzNFcloHeAV77W4whq++v7p7pZirLLE8ikL4nTlh
qI1c7qzusTJ5HoCyyVJuO7NhU2+XwLrQ4re0ec2yqUXd9UBwYtAABIZZJiBlF+ab
RrBHYhzVkp1Fp8t6+EZfBKb1FQ7LKLsiqS2QAmD0im56vf8sNEBOWyjHxpu2zDzb
AGNcOGG3Zdfyb73MuYQjR9PBqAuhCJvEYPNpL3Wx5MGlNB71fnIhj7vevuOV4rNW
A7BzC2pRPH8aZIS3wvC5jOV7YnNJmdXynrhET71EDQIsVkzR3xpkdUGtNXoPT9/F
GjApKYawYGHZbDTcWxqMkBIiZtDKG6JvqpD8zqvqtXw53ntUziX8B65xSfWwtr0o
NQP403NG0u9KehRz6q2JnOs0vXHXudsd89d46lHcbI5vrptEAhn3fqsSKwjeAt8W
UXtZ5uKqmqB27KwQg7slh/icL0+772oIRliUInho4Goy8TZMHH0Ob6vdNO4RVuhh
1lk3I7il7IBWyR9roDW17A==
`protect END_PROTECTED
