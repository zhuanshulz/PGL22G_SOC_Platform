`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SQetTfuv1TUAJHBXgVZiB36i8oBCXeICHygSfECmRc4pDZ1pMTCpg3vrTlOeLE0t
TBPwyQbKM3h/CaHP1fh9PGyU2A3v3U4wSnz1nTMR6nhjkUBVzp8wZVUgZGZpXRll
3gWQlNgOyeTLeQ6v91x3PXgk6N/pHctZ3G+wJH67zKfnO+z9JvSnRR/GOYlVJIqn
B9I6S013yJmtGaqz1EIn6uTfPatGiqC+Bx6IMGrzYtCdCuzveizQqELPpdt9ZTNU
yhAw0Ut5vNC2cp71M5CRH3ChXAL1OsdIjipYOo5S2yVZzZqNcxfw8ZhqqrOS/TYN
UYvOdXWj1kwSM6n7S4a0uY1l2N73bnG7nn6Rb23ZEAqIkLayzU7UCdWd6nTUcGaH
GQFknEQsueIjBo7u9lMBQy3iODIuLhYQxC7W12xlryRTtPyDpv4KRKuPCfMM4q6E
6qYhTwtKsAxncajQwG2VjJe6DnocNx3kLz2sSEYf7ITMLfZKZUOiP4ZL22nWAPWB
W8/cmctuYffWz/FAJgUh5sqskHIP7hSzWD2TGEjGP0MyzkiUMr561ZWjRAmwxwbW
wd71YSsY+O3dsIXOpyAynwg1si5IuUNlPzVzA857INL8/h0IqZJ5sTSsrSGY1Hw6
zefMlVzJUQOiDOccHQ5dmEsJ+UySCD3LeIx7TdjvOd4K7kQkfEq+3dTyZ9eYLDbE
p83VjZdCN8v+5bZNA/cPf2hJ+hxTSOB0FAwThnFh8aCcjSUcPJnkPYn8WTBGIrki
IArZcnGW0fpJIVFRBbeLsWkAlnbx8TvAh5LVrUl9e1AejUt9cMIHvIHgHLAYyzLU
zHrXwyAJ30MmAgkWacrle8Gyj++6YfcwFadUboeErp4V5fLk38yKwKtNAXof5b1a
`protect END_PROTECTED
