`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w3mUs2v3mQj5JxtNvaoN++V4/gooG91T1+7rL7R3rEfKg7DXpm+26tgAZO4+iO3C
DP1N+i7/qjRzJInkwNYj7mD+7eB7F4b65yvUGzq85+FNSAUI1r4VmrJzFiCgN9zR
zJjcQLfAthYIMFHAEoflelq/ZGJZlQnCl7oy8Glry8/YVs3WyPB1WBD7rKzGy8G6
TX1+Eg0hQw96W43ykJh5J7ulAusZUHdkOQwdSZufi28R6DC+3+uIQYiJuhSicS5I
KIDL5r6lWJOWLt5gqnkRTfOMakxduvxBee827tNeqnYOPQInVWa9ecWpKGUkXHIh
QFf1m6mG5ayzIdA84YQihC9nsv3iZNn6MFFYfe4fJOALnyNrPtrQVZXlMLl/LjCe
oRNVUbHGn5JRkNC+UNKhDOMON9bvMnh5JwJdSLMir+fFvHG2y/N3liqXn9epIPTr
XREEIlDeGflQwquUT/XDIN9fieSYDIA2LI+ahKGQ1XElw6XKqQYU4ciABMDxi/GF
INay1Akzl6teRuMwCTwpNCe8MvCVH0DGw4Cr/ct+utlZaUy/vLVGfOR4wEaqGVtW
XYkMs7QLNO1tV4zulhP18SwIbIV568nVWT3OaMNkEuSOpY8H+eSRJfgdRhhZnZ1N
APoaEmdxxUeJXuiq90EJZPZ69TmgdrOZXA8kV2siYoSFbIqPzNDZg0lkA+aiPjC7
P0hTq+fSEysyQwpxeVxxJarJzNpxXBUEnZlO+MaBkuCmtTlhVmzRCqnVviIjYxYU
1rGAFhcPjMaowbsYsxKKKJmS3T/9g0xbw18p1yEm/Qva6P4lw1EKNKLVVh9XBGl5
YaRN5X8CMLBM1DWGgjArLe4V5MyFCxJNOMmuN0fTc5WS49nFARG7JE+hEiBsXxdH
2NOysZbWA8PGnvxKPij6M6wFdyTdL5FkXWUHLVcGRYyicUiSa3KB0He2LmnhadO4
T38Ig1DMqlHOg6fO+No4YPVNsB36rE4XLHU/SI3saQkrfw2wEPMkKiiNFM2Ir+vX
6EJycNCyDTbz/PBYemAywAykSyZB1OhM84wUJ70CWIlfoD8IdScCtUDs31EeYE7j
05oCaATNDJxano7MULDXhw==
`protect END_PROTECTED
