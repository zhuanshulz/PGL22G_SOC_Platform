`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vpLMnmHUqQjyddo/ciBwmpJwrut6DJHi4WPkUeDNirDIZE0r6akPoDrRmSZQoyfJ
aCP9qgnxaz01N1+EU4CB9qRzseQJKJvh/sc3UCrKa0hQUSzypUX6aNPlweCTKINl
0uYgLdFcc9bdd+J6/39BCWVvOStnMsqVgXkFC7E5qPC8+CJAnmPFqoDIyJM4Jt9n
8kSdZL7wNLyx7wcQTbut4QYfhMM2CXLc+JgvT1K8QhPFuMLDeVjaRmWVeDnuUUud
M6DVQr59Hb5PhY1veCPaxuTFvU7qBogqHioSFsLfU+nrpArg1BbWafiBxsz4TTpa
shO2phsw7RckT1qrc2oETC9lghgWCd8/K2nTKbBhr/aJcI+HOsSe725lSt9nyuZg
UmR6CKzhsmmWbTMi/yMscUHn+62OuLCQ4+n863hyqhwchfei4uvV7CVI2FKYJ+6y
Ts6+wSJKHAMVdaNE0Ipo1Fb9hQOQmQyUKWWKYwF33oLUaqnNVT58CSho5Vi0ueVs
Ql9xjo9aMqm4NtgkyeB/txbM3jdqMyr2UVZlFfO6aR95TAZIVe1IDkYgZEEj3GPH
6jsdLfEtcokBB4jqx84fz0by9/rVJqKgkCGajbcu4Cqwa2/cA88O0Ei3oIYcuSwS
FReWMvfxjaKlFzTGC8nnF58x4kq5t9qRsHjabZe12o7tZvmSbB9alVeucuH3NqB9
NYmtSj9XUKpf66CL7mnci7PiR0xYTtqcwJBjNaNO0D81sikaXpOiHNkRlRa/FfCQ
HviHNhBXu2h2SW/e8M5CflMjsPsTj/PrtgXFi5nBrpR4Hme0DBVBA35cZRgfx0og
fvEWNqayh+yv1EFGcffB9Nwzw2BzZcQARHo0TjXLQZMmV72c1X8ipcb0qQSsEWhR
3WXYIyDOxYNKyybiMFW+fLYLA4PLcO6UUD33rh9Vy3jJt2ljk8Akk89sWn4KF1XZ
emo63hWsUGUUDR/i73niwMM3rE/J1VCLLGRFe9HHROfx+kknHlsQZBOhV20o476I
ucoXqrt/4PWHcbJUzKaOR7+RyH6dW1DO5WAEgIqZK5NiJXNnWd52lNgAM80LaIo5
mUP3cdXGeWY9Rc6hyOzQXxwnenEwCX0fSoeS4Y6YxtBkbgTEw9CgjfRyXkJ/9W8b
0HetPzPrgQK0D9+IzCd4mqJzNaSu7cB6LEOaxioVpUyG/u+fZkzbVeNT/3a3IInm
aDPqbLk9vm/h2k2SLXAEuoPSe/B0UsxpE99EiO5DZFM4Qmkt+pX8TkAXtykXQ40f
j+OYz3At49mVjFXPk+l8K8piYlLTXdqOxUg9Xzwy8QdgufS0hD3m8p7oNrfz9G5s
Y82lFnaBI5hcGjzF1dWKD5jdSkL9gSvJ1RdorYCilLlUQTtn8eax0/wMVxAXnIBY
wztxkE1sFUXM3aMtOhSehuHYDeZDO3k3tFAUnjKCN/aS6qdJwTBEIj1PheepEcl3
EPp3kayZY7agJzO1cRmGDLNMqaQp5pXPY9kWlSeQz5vv+2nmR5gnjyxmYASIBdZ+
oBnM91orY67ouZOI0/21JwZtcqKlSIFJfULqa666Cv4jVe+LXABQXamiaQt8q8xH
sC885f2AVK7fjh5GYELhoZLBSwqtzsg8ZBCUQn6EcWAkcghilmTcxhHWqJQDbHmk
5NxyR9SSYTGiU7UPYJfXGQ693Uowbr73T6DxAysYrGtysy2dE/dv7pz8lJr3Becq
V+f/e/LLyp+PjyxHGKCqrscwBHQI8dRn1aoPyC/bo+MxRmH08tiof2wGB77m/J0j
SyiVcYxmp9PNkzng6mti2YcDk4OFJvF9kLDEwiHTdXT2Zn/Xpn2ipepwS5guE13U
qaoPhvYX181ZI0mMc59/+yYz6rUM84V/w9G8rPZq9/Gx9UiSeJfq8xtcUwwbWhpw
fzMqS3mFsd1CLswzzfFhvrNtw1vM51i/eDZPBAPpc2rP73A2VmIx2IASf56l7daH
azJdO28zBuZD0Egu318DROBObbsS72o4pKLomNpoCx6wrL9I6pQsSwXTX99EgGJr
2wG2Sv9Zvx8+G8SuZrj/0u4bXMbvzdPfn4ivmetJLk1chYuW/Tc1rSLVGUR+NHvX
24NhrtvAzZB8O+LtRxo49pdQ/gysF4/gNCUw/iTOoMD7EFvb58Ruh+1ndSS3iysr
ICqczhAtA4HYfP5Bt+r+Bu7jcGARbccVeqOdjL/Pv80hHEpdFnmFDD1ebqqNJYS2
8ZHxKyCdlKJtHSDbIZGxOqslmLdwOCGDgE1Q6+zNYtWrolYSpx99b/wZcraoMEsl
zc4Zb5HnPaJYUE1v7cUS/p82ninE/tpIBb7EiHBRmYoXkB7YX8qkvhKPN1HjDzez
lOYhEhtnUXoi0gOTR85sOo1eW//bIcvx9J5wnEZikk+gEj2JY9simLh4e+H5Hup6
6ZQw9+5NIQLJ5jjsihHWKc8W+zXxoA4qUbMps6dhVliY3K7/gSAfKYH810Z32hye
DttW6+5+ZlwjVbmmSnsTZ6SRaYyBr4+YaIzwJZyjAxcHTsW/iCIR2Twa9ftu0bxR
zNNx4EXPJ13fkAvwSTo2AmrrYkRE5Zad9kJIp3o+F58xSyibg9SfT+bds5s1g468
bj/7YigpPd1TPhQgOB1/LIvqhfuT6CdgrA3vxw4VEOJKSi8I5rMHkzXMcOtITrtP
Q3r4sb5hs/f62XWec0Zs4qjU1Ppo7k3DBBGAkvfzWYwFRGMPVoAufFN6CGTuraU2
MdR1WjjmbQFhb3nmIpM+dWUE/b+TbdN0DYCIGUt4M+962htOWA2IhxUnJysfbz/t
pBQ1QXVK2PiXWONER9bu4xge9riaaNNGq6J/L571PHh55JuPBftvCcMOwBzQQC2P
432ehDEQk8+PBeU7ZAElHVZ9nOE8E1bT3y17LUUT1xgMqieIncBYvTdthR8dY/HX
E0YiVbOEaTerulm4MDVEqrLjwsHO3UJFRTo6ehR/ZO+KGG9V02bE7mU7ffD7xEkO
r9mCMOB2a1bGPbDI+W6tfHov1gY2r9WDr0YXN2b8BIM/C8GDHCHaIgr6/JtYR5SQ
Vsz6dmG08ef0yk1arQYkYMqs6BKR8hYL6ZGEIfsINuj8dB82bq8eZLHwKb966Xv/
O8uIg45fqgxguMJeaG+2doVAq/G1yfNkpImEjptxaeMto5+sY2tEtoocUFVaLEFf
3ljBrr6vxPpLNbg50O1M+Xmo1/DgebQ/MZZz9joQb0iqV69BPYTDnT13XGUTm+Q8
j74xfKzGIKftIy+JzhaosPa+EmyJQYN0mo7/LzpiYoo0/8NnnPkY9mVCHplDRZQM
ZSLtd5pZ5Nrn01Ps2SSMB9BbN8ZvPu3jyxto26AiCLw616UM5bblFxyGkwF4RZvi
sUU3oFy4bgEpdJX8o+GNb49snxyofXDZ6FruxRKJwnyjAUR5awhQYv+CeROyPZvy
6cXRTLNGRFamFkNyJrNX8H3Yh7RD0TJRaWoSyl0c57Fn4IbgWv4OLxmG5E/aWSRb
A6+zKLjrkFh60dAEX8Oo915a2GyOla9MfYWf8fJCdmbBxcCZJaHMlEI1rswVjp63
Mu8DaGSycCIoa1VVk55pt7RAbXqIutvAySx3lYLB+SizxgqE5yEjApLRC9dKKFuS
ar65h0EeEOzUxwfPHBfHfLsfgjSks+ncHkhVE4i7Yq6rngqjPTyHw3FhIJffUH6w
fs5ViLxHll499ECzTNAiNArcvXyT5i8egWz2f1ktpwTJSMubtKgoEqMYY3rrDOea
bf+r8Fqi4YKtLF2I7wxbUR9UVtJ10DQWcLJhya9hv1rrFmwqI371I3EkrKbATkI5
9zKkkpolS03Oce9ie+5LEoOi8k5crYBVCcFxmPiz0JuC+33UUBEkIHGXDaBonKpc
7b4SPiGzZCauem6sDq/5vi9JC3Poz+qGY2t/G5lngzFAjiYbLPqp6z1yYvp6o+uW
2EWalZ/kt1wxoM1d7wY5naoFSX3eEjPNM9lQLC55xiJ8XloBVknqCEabyukis1+E
WbnH+v2oAJ/HKuhzLDOPtvlCoa92ouZIAk52A1Z8973pZ2lK/I7eMaXzmeHi7aIN
kkUezSt2M5C20zKtud+75T53VMRuDUkWNBFOT3AfPrJmDqrni4+p1vMCaTbkLbZ/
ljEcEJDWBExGFlDXL8KDgUREDdlCLBoqBgZQTZQdTkgXOwOc1rfe0vB52ZWXS2QQ
95TAJVbVJaxv6v6xuUB6Htu+bOiDO8AlKucDErKKo54d+bHUKLXL1zIZHx0bcgi1
86wWwnlaWzcNut/UdJApqO1SwD7m9JwS5MbYyOFrs2HRShLPKOFRbxTpPkzjOnLB
MernL7RTj6XdzpufeB23zt77lbmDWjL6VLXhZ48MhNxI3uUKoBbSAhLYm5Eew+EE
Np6EuH64VbnqwJhsGozs1NFJdtsx/+ozw5aE5PjVkFJvcVtVnfdXRqH2iHzM5Me/
Gneubdjw2F1hmNsmU1a7eRzB6TqJ7rHddxjt+feFadWvUIyY5/HfwlEWSm/hnYLY
O24g+6cZ20VoFr+//gMfCwSWlxIxwlyQlag5hyfmVKzoXDFM+6nvd9PXlkQcp8nM
EzVeiJ2PBpue5qDZDsbrM19zAOy5w09atGZPBd4czjFRzLSvSfh8jOevGJsgcLKO
PB3ElEyefaP9PBk9WIKlYXjxVxo7bxNmsihFJFj3Wem6n7Dk0ku4ucKS0a4TI/t5
5yLtdDPQoJ6zn/+9KI08tBY8xhnc+S61QBrV0M+X3gpY94ah8h9Oda366g2rI7Jg
Rk3/CHECxWt5iae/ggOF1hijohT/bE1buuOei34fAiMAR14w1wmUooTDT8QFrwuF
5PF4dQ5DK+JCLp3BDU4/XzCknLunn9WX8ZaC3BPeLXqMHcu+cfA/3ln3XNuBc5aN
cslJ6hg8FJHXG+0Q38r9ygaBtdlq9CfwJ8jQN9ymTTsjw7PeBuRbvAX8cd5k2OP0
5vTUWKOG19qMtSiK9kXns5mX2tvPZatyxqF9fDRtk+uVvNbBsnCXdg2sbwGHjj6T
GsCh+WdvgVxjyj8v372sD56pZq7zTPuHiizZK7obLX6pWdecdA3vnGgU3uOzNvrl
kCdVXais/sVr9iTHKi7vwj6zmHC7NXiMMrUbnxlFw600rlTg6b1s9ARPVtx1sjhn
NZzaIkSiqUZtka/FLYeUWR9hEzK6p472m9/SN9cMlf0Sv2a631sKPm4CSY+XL0oF
v6gsxN3suOMoLbRv8rnfXXzY4ys5IY3cVgZBOlAC5+Y6SN/kGXPyFtuCDFPpvQ10
3xvlYRF3/EmHW2UOMGFj8uE13wWqlM5sgIhO4GhD4qKR+Wpjpl/PRZsthlA30Aef
X+wEKg40SetzgWfG9Xe6JQdi/ozYfMihvKEVYzbI5bVR1jUG4jO36asnM8fJpl1o
iswbm0aGO7NOH5C2XvtITAUaa0xdvfrDkTOxVpmyPGb8kOsyJLIO80f5Me/7CZZE
zT5fWFtRHN0+jx70c4prklC1tkEABMf62TN0PIldFYc1a5iyVpq13JVW2WnlyntQ
xo1j7/O4NLq8CesjNF/20uFO51GT0078swXfDt6P8uZhDZlgUozdQLsG7DUGtEfK
LaxJWFw0+sp2eC+6keee6Ke40GCu78IiHBqGc8I2HSyrvXUvqWicbR0x05EO5M6h
Wv/Yv5W96h/j+2MLBbCpkHpkqVqC7lxAYCBmvihAyryeGOdyYkNoCU+Px6GBBP1Z
S1X0UEJZdnAKe4vtyyW6MoT42rBzTZuuhrS8z5LG4Ls/qfGptal0aCWJBE/FS1A6
AF1dlqMtokd2gi9bS9BxylIzEhHyOb3QjdcDgVeNn+Rb2V6viixu+yHVun0mu2Tz
+5RyzPMSlFm+BLnd93zewu7AqIW5DnYq1059rshtm6UaKuOxB7xzHS5j8m1Gg6H4
/QpbYUBFEdBjNuxE3KrmpBiwb+dQTQ8l/SjBbsSZ9yIyPuji0w9982/qH8Stj1XQ
F0maQeniqFE2KpP6uMAmFVaql2OAqYkc1z9Gj2Mo9MujAukGEBwzsTqvF8i6cTOp
AItHdyNTrKzJrVlkj8dxGlS/YSQ3Yzm8bGYSBBEa3sHEF1bbOTYrsybUAUS46bkG
gHuQ4NDx9nEhpe1GrKYHXmJiS+WyznDVseruFMSBMHOzYfWHYE3KBX1PY0cyXDBa
5nZfH5nelpeb3BB8NP8M/9f9rg9+XYp0p1+A0bG8ieD4+sXSk7ZBrRat4EZ6nvfp
xM5t31OIoBtHISLqcNq77I3DKbaAVcgL15ttY/e3va573xET27f+r8GAt2zOqlmo
MTOOZ24GccQugSynYv41ocHd9ayhmNZIXP/MRtQ7q5VNdNIaSLijlUu4eCFXEcP6
V+AtPTxE8E7ojguEJn6j16FbuvmSXOWLL0e3dljKSDRusgLKcEWDvkL3HeC3Vvmm
DclxzB634TsB9zQt0W13vPWM7WcArlrd44HljcR/9HbnsNlf6I9BnjHCClly+vhY
THRSQO6kSBsgJmoejyoXgge9EfhwFE2oBq527buVeFZQ/lTgnnN9YHvbJGkUHkJc
hftCxz/kHZE3a5ajbu8jyqd7+3VPw/PaeE3KA7w9/SitjWpfv0AouhJvjlltNej8
yJmlcFwukcPVALWw626GvQDWufHley/mdhpgMLDwiNfG8tfQnDJ7ySu4RE7NbFpa
VaQuKT3pjnuSc6ndHQG4abWrgBYuF3ezLOe/FgHOs624BRzuvmtI+Wrra3dwtgHI
CpwV3Q/tw0QJsnP5SuRNGJxs6jg4K8YpGKfFnLcTcXqByjyKipz+3eb6l7F0qFs3
RQci5icMd0N35BJxtsAbwVcx1uMujDdNFaBAjdenEi9pslcSUgW5+e5tQ2CWMXQd
YaQG5lDC51Bzc4n4brACQOa/i64GDDqBQpR4Fg3vvFU0HQnEGj8XEMuKolZxPP9q
8gQUpsoum1kQamOfX1AuvYecEl5lO8XMHzL8Cd2IqqfJGDC5DETqH7XpXx0pKNHx
NKPT34jgOaRUOcoOshCo7RyHDp7wEPkFJDCFLn7N23UolUI7GXO1MT9cpWTqZa66
DWqQG/p/iPDiMKUuqkPg97lRu+M61APnTxpjIHC5HGOhibDXbXLTmX2gq+mtWS4B
q4Ud33lGsX4DT4gpc5vyCbBp+eToeMnYaWs6N2+NApApCVxv8WfT38DwVJxgMAR/
gDZ5nqeYU9jPsq3s+88MUnNyDa9zjynHNjtk5Am4WYpkP5anvuiRhXYpdI0+/1EV
Ex1PdJseIWma+KeB5TAmsjCciF28eS8sfAYRdQH8seUe8h2x0QqPMF3845i01nCz
Q3HuAJ9B/ScbGLTXXz0p4L5ad1483imLlWy2Pf70hCKlgv+WhkEZLLuEUlBU65Wp
J72V3EHOTLunnvhh6uenauwtoXutpfaTbkf3pzipEmkMfe7GVyjrZABfO4PNsLYF
VCfVwnN0zactWokKc57IaZ3WP8mExND7TSYwVHvU0aSSkhjfDVJdv0rtKJbxOR6I
mpQA7oq2Osi+/Mkga4q3zzEqXPYMJAby/nhwmK5OlGuWOd96PCKNzRuEjBejMWHi
81j4TWJfniaVccYDVR2t0n1ffaN02lXbWOAncZPWZlSFvNX8sWVENWQ70zozGheH
5uctTN68VliBtY1zQmKjOb7RqmDTlpxwgeNswnE7GSl+2BlNxXehx0qmSsKZDBPb
iWJ/g95ip5qYXCeZDF+wtvVHMj1Wv0tsqAIhTC6XL/zEeQpAAXBNSTTj9BvD9fvd
Jg4hrlgk6+1MQWwmtYnja4jylOGZYBfc3Mao+azlj5Gw05URvxE6DUlgs/2X6/gv
9wdltEJ6wydq4uUIjR7uJzU2ThpzHBWfohyybRTd4nLAkMli754b65y1+XF/doAJ
nTAjbgJke7cNMO2tyAxNDyrx7FggA6LXkGtxIQ53U9vULQX5oajXFTxHEdgcE3Do
a3sW/b0tG+E8piaBV6J4l8KRPUU+BuauYkeSMq3jm0Jpf8vuD7BEFk40+rY2nrqN
v4oxoBrjzjYmT+Ixaxql869PbVqAa6o4rHqS/2g1XWY+Gxo7b9BPsaeKS8s/QyJC
VV03P/tL8tQJLbY1HYN+fHWF+jWHkFTePPVKoi5tYpfZnKr2ZoCQz3Dv8bAIkndG
K9/kBxUCZsoeMYjuRKkePqLSWA79GPEgYuTH+U6fOH/3IUVHZ5v4hfjh+NodKyno
ThuoFS70Qp1lXF7EMgkRo+OG0a9Y6lp1phyzfe61pUb5vYUYyFGx7HjzFUjWHefi
1bV4Keoeyrh8C6/yMwHODJODwtdNYGyn3pJTV0nqCLlkKIThSr2p13GxpB1rx1A9
6NnxA1sry22SQexNNjGTsCNrYp5CSV+Ro3HdlUMcI99EJPlNsEZMw+nCoFyyvcJ6
9U1IaTQNLswQix3w/iQMW3ABc+MS8jdh1TY+sKeNOp9ZLbf9FzMXoHjPiVQVT71S
/r1MGBbPzqkTdm6IMOAMP68dS0EWS1w8e4Vnf5FkaU+zQLLZwcsVwBPnHyIjRdva
VUFDlWVJc1BUGabpETYDcq7JeO6FyLjWTHZLoP3ihcv6q3kYnU9byw/r+eGimf72
YEWYZ2gvBnIX8k/VoHcuHvDCFOFp2ZL0R0Jq/hfGaLQ3UEn+DQmp8kBOqdIBewM9
K3kXmTJ4IEHhv5ercM6exY2BgmSfDF9r4kkTU1xMKP+lowRtj/nK2V4j8v7XjtSp
KkvuLk5Th4G+e2OMtDJNPcPHnspmr2ZWBp/+/7Zar0clBZ2yZwQ+ZP5w+lE/uLrX
xdJxTp+kz9BbV/sa5/eqBYLuIL30yjkv60LYZOU54CcdO0a0HG36dzevjsidh46+
WqqKsmOCEQlsfAu8DgGIKdTSJD27XZRfU/U49yaKBs9fiBdqXFBIABWD3mFclAwS
QEbaL5BX3iSiyCQr5GESvPrmR3WatSQHH8wP2IR9f1JwnUx15lO98695yHdYzgUq
+gjeO74qk/ixnQWZDz2kfPjg+bi9ITH4pYd9GwYDKUgBqGN4JKfJvTyoQ5AgOxCB
W0T4tL5hte0qoK7M139CW3Sd9/vzhFgVQiNq6wBVOJmmK4TocnwPFnib6yILSFeb
ICEfIj64Yf5gLD/Jkb0f1CgXGtGF4Nk+sy1s+NYQuKR7WfMxlrcbpinFmLto5i4S
/bT7Hl9zWkkl5w56qIQ4CWO9VFXSo8yGVnY+UvnUu75A//X92cUFngkg5lzo+LI5
4fRUbtrGynopZEyxkRRWFfG181B9Roum4wUvA9k5uoMlJj6yiD6VC60QxN1fxdts
h24oFhyJ0NChFt2bcZHPD62Ou3wTIq5poIJDCLmvEfJ6gCMUdBy1jmvV0LeDjcCc
zx2uu+Q6zUFXiH2BQdm8pKZs9rIjwgI5tD9OdTJ3JYqPN5nfcwYOoYbZY9fQxfmc
kkKV5TB8NrDTCjjWuU+4ECRC0pvfpgwuERF/GgML0dkj/xjIqpuonxDEHwebuVuJ
3kfKWnmoynvetrDoF31uGxbBLfHS8qh8cHBq2eKcY9DN8ISswuDqNtSF0KEwp4Hb
sXRCDgGsA8YPnIFJTM44hCMcl8l/B2FIXdimdG2MGVwvpYQdxlLIb8qJe5env3k3
Vogu6zYoX+W70hHrM1ooCq78KSYFgGM/6bjJN6bUd1V0/75bVAmby5oLsDOL0GQ2
u7yPm58M9w4AjI7r4EoSXqcBD2gNo3uo6u6LROxsnrZJdT/t+6fkaznt1Pd4rGC6
fyC1uX7ws7tSb5hgCGO2YshvtupNhS/XttsGN4WbUzA=
`protect END_PROTECTED
