`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MWx1+vldCScre57HoKK0gkHQdcWIjPpEsfdpm+rDSqB1nC7zW6Gfw8rOdW81jSNY
FHLS7+PjmegiHRBX7b2cIvpazQIe5m0b9YW6Fld1YduqFCd0j9CKhJmhRDP40och
RRjNs+inC0CPZ77slgr6HDIKjZYUtiQFlMrpG6YA8wXckbZYi13F4asPINh7F73y
ZNAL9cCH6iweRrEZkpyC9EI4gn/V8PNoxxz5LhCzbMEgMyP/ZDWBEZkBujYoLlZB
xPX+sjdTW5PCRYidd0fE4gFBYB1eT/UdhjFS9fYeh8tDkxg1rdo5wISxazVLY6py
YyXMY0QKozfXrI9Iv9lULKUmirrlUxhRH58i+BIRhRof1KDz/gRleh5fxaBjVU20
l/I8xlnjUr7iJ2ZOLYMDDtNJ7FdJ7/GWOl2GXGZkMn+oxlbz11xXw8iJY9cZLOHf
pMMob7LmIC2UeieD2EUB5d1MHL3jL+fbCmqXajrUGVdaESjjTEogxBimZnkXaE8n
WWDt6c+O7COs7ww3WCnL1yRb/EhaZnZfV4DnFxikL0YmskzQXPZ+DJIf/hYDB8iY
HJeyeq158hcVQoATXXsHxzcyNf4STCTI05y0I/SK+Zh+Ropl1syqEtU2Z6wbFfyt
EzWj76i80HFqsW2p7hvf+hezVcE3CAZQYXXCDRtnO4tj499Ftv9/SOmRaVrRlWgW
Zw5vp/Uie1dJQCFTOb7Rr3AOIW5ganf+dbOxhKOOI397m6iT6phffP1hBCXh2EDg
ZTpj9Z5+xrfchk9CxgMI244g5a3MZLXbKh/ob5F9aKJo+dWNOc3ktvyCqHcp5R5i
lTi3f8MXkinUWtuxWxa5HFraUNgp2ObaxEdycyGA9bXyjvHQYE1lgHjpfSYs0Uk0
dTA0F8e2f/mKUGhfO3wTbD2DnLQNBhHudmOWEQUY4B/vxwg+xdUnkL7+8lDSpMU2
OKQANsrKa7p4Dis6BTQX7UldRhNunqB4651mmyRAJ9ycCTAQiWynC2p+DgRzAFOW
Ol0gpP33cVf+hjGNeFEnjl6281XwfLqJY44dHSsEcXwJu6vGRyqw2BOnvSB09HGE
Kgy4Ewd+r5SHP2dXjaUbICEysE8ppe56gOs1n6RkFzdp1VfAwcchAaldypovI1mR
FBcniuCyN6Lzx26ghwr/txcglJ9lj36eXCv2gPfKk2XL4eMAUFxbNbDyGABMuQBc
exP9/upyZBq0PH0gkXlA3IhK4ULeTzQWOPn1i28bX/ubJH6C6lHsxfvgtmtc1Bqs
APnZ2j4cb96v5pS55xsX7TSg4iu+c0eeSpN9oWbJqdtqF1XoiDOAI3WFZs6unMpU
xlIJDwwNlJmbhl2qEZQ42ixLBxUBz8qGpb8iQhmhxOoQvxy6SmWQbcHfr7VwUtLG
N8z72bMiQsy0iFOUYu1uV8ZV0uRtmi7UHZPWl8tLabV6M4wCk9r8o9rrRxrEiZyp
DkSvgxjzMzO171aMMfNqUSBVvpFhEcXDEAzk5wOiJeYpfVI9uFl0JmoCz82T6c5a
AoPqx9BGPFv9e3Sp/SjZQBXG3R01i6yNCIlM48vBb7ysQVtIqVIBQeWBbk8x9qAH
0eufDM0y3aeQmErFoSvo541cRBnNKxTLqSMxX7wtlDYuCiMuVla+LvRtPWOaoyPs
tqDaVgnGf6WJn/FxUIQBB1/NRD7quSBegCq6ahC5u45eaUUv0uhRGOYXrq3hD8Bc
sV4Ky29JBKRtvDjXapeL/Bqiz2vMfg0b1ur8Z8lzANaExjrjsEqYbzLXwl5IJatq
lbux3U3pVlfXZogAkW3hranz76rqV8yBF971dsXra7EGKcV+/MBFQKqaEuA8IiRh
sPCU4VnReWheB9e8MPN0vI112L5FfihpjDJkEw9Xr3cuhyyEumE7Ltm0EjzQBXyE
IVWEWgovQ1c3fgqhRew7YILKssMGbURtLhMm5sEI//3DnAgO3B1WWJ3qD5sMTDC0
pWaN2s+WlqipFotbAhj6Gy27Nnpo0IfJ8Oq8gFq0ljL/ES2UMgBCLBfbViGsYTyj
rQsXg7Fl+jhepvshaiM2t1fCZZbiAwo6G4QMv4j93qCJ7g9qaWiu/wpgxhCtGk3s
feMZA7YO2hSVhKCN/EU83qVEW3NedGC6zBsqy3U3ObuqiOxBukmg/lWgZM6i0cIJ
3TmjfGMB3ujpD2fbIGDfKP+fqCS9TqICU/urECRagry0TYiGxJNuQHljnMkGDC0Z
lHhgYR5OBmjtyNrcswudRWSUT8AJOscBGuipiL7t4s5KDBcBJFcGTWXFtjDKz9fY
W19hrZrWolMqjdKqZZORLTLO+45z0cNyTdh9T8iRIClTrLxU0Jpd57xdrAjJIV/k
cfMAHWTq/m2uvvgtUkQ6h8cx9YRfmDD2WXMnw7ZZl/Bw9FgPWVdo0ICETFPWnZeb
oE/11e6Q55US6Ev0kVxALrzekyP5F2ichuThd9HWwhcn2ERlV8NDEBLmMSVpsob/
jfO8y/oAkJg9NdgvGBS8M0YA/ltDDZAGgSMwR+2mJ5n+VCUuoBX2jCewZ4nn5Wez
23uLmCij5Gzl8j7Z8/HepVGYTYLXwkcnP6Ni5/91TwzE/QiciViZOnOdElf9nwTN
WsJDjIZMhBGyNEip4BWyahKpOS3WawoqVnBBuZHAUfGYXrlnOzxLHymA76PxRNis
OO/GZh1zZy8Bu+uu998rptq0eyeWDN4H0R4LJSiNhOZWJNlYExKYadUHf3DMbHRV
8J3AJfRmcT5FWq7mBz5dRWCblEqz/lAYz9jWfMojvVGoxGmo96Ub4vRBWFhKjCm4
4IdBYf/J+a6wgaZDv9mconDFXVl+nV85MOx+rgMGj4Hrr/QPvFzXWY3ztY8VQxaZ
ZBfNPUN6fKQCWk0A2aTICrtXpaYsdirblpnahgEWkmrLMnGymOQLYEeJn4Ze56zZ
Z/kaatMYTIP0jskyTqQ5K7iHzVbW/Lx2UjPZc3MxtE4I3csz8MX3jOovNAoRRJz2
O6R8wdTGfCk2CwC++2e3Nzd6SuH+Kw9XBT/Z7/YA7B0eFqmNEWq0KMQUZ+w2fVe9
izD94qHYm0N7cs7cSisGxA==
`protect END_PROTECTED
