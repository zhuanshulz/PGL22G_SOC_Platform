`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eqET2qsXjjKz9QA0cyLW7hErQlirh60KdigcHEmWXObP26jwKRvLasL37XpQeNuh
/I1YE6fc8mrdquHYe1KEwxpnoF4X615ErkPXvnjWT7ad7KrYB6JQoFr2v6v+Pyc8
7sFd/iNkdWVMurKeEJHuWn1OIm/fw1X3ykloM0XVN6TIit6D24gr368HfZhiBECB
LnjOTz0SVOY8QyD33tDexCavnWFjujklEfbiHJ3nOi9zj8+FgmEI9K+jMRNwX7G5
rE9Lgv225iv/ppZXu3tSfDbQAlqOf4liAxVYMjyYDQ8f6aGV47ZmiP3bmyui0F61
+HQpOI9oGY8IRdKkZSnVOs/wiKJTqSBFloM4P/DCGHyZrQcmzcWo6CEO+Us6+F58
RYdUr9mTXawy+Rej4zFe6VpMO3Fi2pzFqXy1tw8eXTINdpIVzgZLuYCvEuIa3EFR
s1PIMZJG8OmZF1+vl4aX/Fo9MdKezV/MBfH2JAAnXE9jZHffPEg6C7Sieglmj2ec
gZ6C0XNcr+Ye3+WTGD5syzLN+GbMfDXelHJJyP0NpxAm2NuXTaKQi5WC1TsFQTJb
SIf/b3zQUb8b9sal3U9nAqGHLUNCOXGB5H69fG9L45CHfVvSiAU8E61pdiLhfOjo
T48PeeJCPSjstsTuheH50yxFYLSO9yHMKVq4dwvgZhkF18JLcHlN86qewD1RAx1y
/HWkuTQjeBT3TXPOmWLqqbLjbN9bsym4SVySzI1IBZFp6eQwmAkJyXqwamZchIbz
JrynRsIvlTPpMzJVABkqf8E2rEBFS7/RXW0yqn9fR8Kecf31KZY7GzZFMC3xfo3G
+k6Sp4kNKHXV1bVWuA4kn11ZI/4e77sHHDjc7lQlXyyi/yzHnHermubKCC37p9h/
OZaVCzxPKBTpmZG0iZLgT4nT63Mm0d3nx2CB+IOLiAK4fCODRnDLyBvhsQUs/DC4
eTWuUjI/TfXi1EzwkImnZdBwJrd3D5Lomrm3uHT/CzN8xCsfS4nJfQ2Hl31M/eaA
sJ8+Gsp70/CYd2ThlsgxLYS2wsthNKXW3u+0QGXTOJoab7Uu/rcnQUcgS/ULyWXy
OEOBhk5+Ssb5DlGj1H7ofB0U/068dxMkjdwS0T2hePj1x79wxEXNn1nWinPKwJcf
zAXjKG//yyMgbYfktzHAOjF3w2OklSmEpT9WiBqakVgkEAoJj5LlL0ZlDVLrj0Tp
LKK/AlFPo46+Z2tMMW3YPkV7VYhQysfgw+4oUKwQaYDjSbFlKF++xFUb6Ig/C5rc
iqCVmUaoBO/x1liAzoNLaEqeJbuUOypOFFjIu0GMeyjuxVXNKKUyN8zORajtvcmt
/kjbSF91etGnwt1Fd0+ibHRNV/Eq4rtrNelcd3GdgfJhdZf1I0TTJ7SMBgFwbio+
OM5UgoxEjqhQBccwRvD43/ImE69cUlKVLBgzF0Qkf6P0u+z/HuUsx/nnV+xSga4I
AI8o4kwwgUqwuPQ/3oO7thQLAdnL4N7XvXQUocdemvu+LdULti0TPT4FQwZx+nl3
EeSFiZnEIgAl6Re3lTluwULVKjpipbvTvEUAqQquW1PTJ/Xzsxd2PeaCsbNyPG4T
edwZU0UgEPSf3NTtOxcD+BspBAMoKn29oo4/Sn4Qtlx/tChquXHNXrOB9J1iF6eH
PonOhApQXsKvDFdcl09kGAvi8O0Pb/wLy5wJRkJY+QOyN44caTPXNLPNXL0ghDvK
vlXF3eA7cI7EJH8y8goNJkj5qABYhwTzFTcWXuFSfpFeDklm9MzSNyQsyvoRnsSv
qH27n8LglhBNfcZ1aUp46HOJqaPL2HmE18PEUO8kAfrw/MBqw2F3aAW98q1+pDyy
9PAjCIVFvDCsxAY9jAGUAVYr1Gmv83qos90cRTgtU4pr5Y3sOhT9XJrJbR7q9cW1
+A6P+/oT+zyrk4fvJl4mXcyC6LlELAMWcvZ4/ow5t1cfCwVgGuRNaGMjGCIMDA7Q
RPTFhbI4ZEsssFbaDqheno8PK7nie73X5hfQmikKmwLmBPKKN7XYBoYSprJfQHev
M3EzKfQTH4M06q3wfKxATqPHyxb8yRitz4r6bgypD7dUQUD9yRk1hx8m5SNJNUVe
XIfmY7FG/ca8zs/Mzv31x/8llN5fvCDxzD61Sz6yhH0eYLqAvTOAX5Cl4Yr5Jk0X
bS4Ao6N+LxZuzK2oPynUAHJaDo56o6TNuxPxer83LNk=
`protect END_PROTECTED
