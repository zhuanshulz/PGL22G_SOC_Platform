`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NNVagA2m+WXu9ThkcwT22nj9TkTBhZTcE9jkGQRUWUhfQPlCP17/m+Umaa9T2Hxp
hXlnrujXBpeD0FJFKJSPfrnCIu5Ne3ylxOE+AgBej9FesFKJg95JB/XXISdKNXum
Q0frMaH+OJXHnNbySAihy9vDjhsfYf65LsVfFS5RPz0Xtj6q/46xyVvYpaGs1LKp
l77LYwo2B3RlcBcHB3YhMKJhQlAd1skK+vuI9VhXdfWT+HqkYTiWqHnWCskDLieH
/zy0Oc7/mtATKrGGwQ2om7Ud30S+Kr0Tdut2xQ2HN6pDvckTpBftn/tXQZMzbLEP
ocoN7hXuJ9H7Q6cMn2rDeYPwjQh9iXNxlhA1K0PIxMTa5IUISbjg+XTUvfax3IQT
Eb6JUREMNKUBTpA3HHkCr00uJY0vB0pfgOJt1HrFLWqU4ciWgy7U/bagM9ty8inM
N1WPJ31/DR0Ik86TbajdajhaC92Pg3OaiHdNxoUZwXyo86HEKmKEXBy+U1NfGSav
awEYh8CVmwkpE4o3EZDSuh7NUBSgEYLccaJZgHJHHoG2fyoH9I3iubCHSkudqDR1
8XQhXBxeeu3QZPsHVHwZlRk0RN9jSiauRsQRl1PQ8DhdO0PMITPrF5iN0Nx9hXzE
L7wtxjVVKOp3RU1VORg5tc6VHnL9sdb2iXokoU4t/PFquss1OjVuzsnJwd7KR0U1
9Vpb++RwHa8ZFoUI/LaGJwD+7TsGS9HtjgT0ZWWYm1ZZ895opukk502uTLv9n23m
XT4xM6/LT5SNwJx0sN7G6htFPye1LqhKv/+Q5hAqKS3PgTZIsvnv2OkInTv6aOsC
IriILirM7JCHM5plDUwbI3UFjMMNZPF+rT9sCSSXlZhKmt42vSfe/tLyrPiA0ORM
vUyQg0p96k7EfdOqOi92S1trmJ1w2ohaWARbhO7lZTkxM/j27F/4d29i8IIt/Rak
/kHEP4Q0AXFmrxAzgY+TGIbRjDmkbQDC/JkECF11p2fiS5IVPyaiKHS/3umffesw
vdP/xYGK+xoKZgOuWqK/Hvrhh1qReTP2xQPPCK0AeaVm1x4tcHWY2drchzo7z/vC
my42ngqt2btoqkQEbt8UA46jj7H8Y4TP1skvP0whIKucrfWVEruQSOmhGRo4gTpm
Wjh7rbi/u9f7iyivxaTaIwb97Y9fdXF6f4xDfAiG2PqckFKfejwtNE2AuoTf5VJQ
kQNTlcAKJZtGooDh8icrDfvIC649+4c5A+tEGhPjG3u/QX2DpBh7UGeTThx+tM2W
mP4C6JSV3+EUYv7vxGMa4l0T3ibh0aKtv+73A9Dn0zBAXtQm4vO7XeD+ywF/024v
`protect END_PROTECTED
