`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dmeO71sNtJ7Q4sOnbnK6ybBD9SxiujLvAF72pG9yofkDU5g9yMlsX0MLJoXK0yMd
f22L+25PYAlBDBZwQzmwGGJtjfWIS0RCobC6utKGuot7f34SHkiqfOCLWn0vAPa1
7Gr39uWg8zYinhh0HEoGzugj3pvB/RcPjN7CQvoWHTJcVNjdV602/hUkDCftayzo
TwNI2sBlP2VdlXw5VAo82j+T+8f2TNReYnZPYG38PdvYjwjujKfQHZbRMdNtoCJy
CBzRa4PaAPMbXuRNopL3ZiCYLHCUqmBGb6zh+ZiZqo+SoJJErQvHSiwvHbkzOiKp
HHdUq3m717FHlhnVmJObGSAxzDLBgodW6F3G3ULu+snHwf7OUHgqM+BuZL7Gi3y9
/E435oiW4dm/WR0UpVNVBa0L9o5JEYuD6mWzAqnTNArN15kh5Lfem1UUCqFvxf6w
gNhkhN3QF5FMVi6k3V+HMLfqn284eimoMMnPrkhRt4+hsIeGUj/DMFfeVJ2up8d4
1/W7ykPAunXAa8vDCryu4ESrS2/D8YYKKr+ZqsOzGtyXIMgXt7rs6g994OuziRLU
ZhkfusD5HNClglo00PohytYQcdtAjJZls7mLAmw4gmU4IBKhzHUt1p1trk7+TWGs
kunEZZRKR60l9hbOP1K3D1+k+8EMNl4ik2v6y85xr/C3kC1jhJsD6x3JS+/CJZ9X
lSzR6LT2SILDAwsMi8ziDcCkCyDIdJUgJOoL9Om6P7OMacTkUL3VrG69T8R6NgUr
5fAEIkUzMZjotKHYU5r4yW5GgsOQnq5c1NWUXqIzjmICsto5Y5OKJoyVdbzXB06J
jlqSyx5BK5VozCWEf9ELOmpDCfDYg+sAuRRdkQiWS+19PObrUgcNtQzZy3HgKKNm
QCIr/Ax4mnVg277sf1hNY+p1UFV2I2bAQrb2shq+lHx/9CFRiN3f1CrDU/XnPmKW
ELSI8YzKVt35ok93Q1zJl6OIplZK0a2p9jYj4sY6X2+0UBUPqkvq5tYoIx3lTvZQ
5W3zaC+5rFuweyNvGEFvEie8sGKsKAUgmcdM1QJqrVA16AJHfOHzBcvpzhBweTLe
NwpsQFHmivqwWnFNlE2Yk0eSXp/Y713uyMQHGzP9uUI18UYHu7f0jGwZRCXgwcsO
0teuAOi3+e9EJVhsmI9nrMTvvWvNfD9crLpgGtwAc3B7SKzqhiFGhr1rDmSwSHGW
gtepgTOQw9mnkSiOhCnCGF9C38vsshvhB2I7SQPcIEDhG4aYHcQ+dw1wooOjCtUe
c2Z3Mnv+kyQH9V/3BdmA/uMxTu1cibKO38YS1m4+2++PtVB+0/xBEXkTXg5bhTL1
`protect END_PROTECTED
