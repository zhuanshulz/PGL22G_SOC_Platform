`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j452pxXcZ76eK1iTzVbgyKe98D4yUq4y9kLIW3b1uAhDEFZzI5JdOiJLRrnT64hI
aTQOW11ejV637yMX6UQbzFVQUt0746ySRVC0qHqW7ZjO4Ed6Q3kXi0clVVVbfoqk
2Hjrb31HysULb0JOzEl8E/UmJle7GceW7GFrwCfwy+MWb0dRhOtgFFCmgZ74P/jF
W46dQpX8TFYu5EqCyOCcs4qE4JADuvsI8P8E//bJ4q++Wk9IP9snrDHSBnHKYJAv
mhOwM1uSytkiaGV1WLCQsr1T3S62CVnoNYnYIP/2XbNgnGmkDC9lRsy81LmcTN8D
VYvXRZlWSw8/+WyN7R5mkYJvf9U5aegLmzqrZ9TTaSZufmqUmh8EDU1Q4IvyLgTb
bRcGFPTmwLWmHgJbIeqC5xSCZisMSlcAW8C79Ikx4poJ+6HHzrqGem5/FcSzV4WA
1dRoalRTOn8VE7qsJcSDKA==
`protect END_PROTECTED
