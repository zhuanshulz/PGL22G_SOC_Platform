`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m1Mqjx4WPkwOLaA8LqV10V0xqzztCe6Bf+ul7PcpboXIdcHzVyeQii7tgivuIMJx
bd+b9Ngswd+qx3AoM6O5ie4RXLORPV3dRREr5LZYdkJ/t4b+JbWDRg8Sur87EWym
S9HsmL2Ogy+dVeI0m4XBY99AeyRmEIu/5nCxK/nRMK7dy+YGTgJEWkabF/gtSqMB
1bmQmVquYSotkIThBhB5EgSmDJ2EJJAyd7m4YxDY72aIr8eJZN3klD2xmVcnjqz4
bPqMwt4xGhKaEDJ7an8VOY46JdB681N5VZ437xiH31sYNhT+UmBy1sNmOO78Mt1P
k9f67UMwsmzRDgjIuLWNMxJDGTt30xfdP2m+ACsi+cYhWUdjc07hCd+AJR+9G026
IOrrjFEm/bxphc3+VlxWqdiYkptO8C6AiUuCbfidTU/on6InEShN/RvbacpSiVa1
0tD4KRnkdPSkeKijComq9TRQfnCKmZ8h+3g/Pic5F+yCptpHAAaCIcEEMpwNj/dl
At9AY8ycaLb+f9o6RzmJpGwVkCQyEO/p1mOtWMadKf8ozps3XNMP9Ifb9jrzptB0
L7UT1YN404t/6TkSkr08UJx6iHt4gXWHHwHp3tJhE9WqUipDv2Yr6dxKVWjG+1TD
x5mCFCOSnSq+2fWVXwL/MJ9FVr6p2bCli7l/jxYC9tmMUvaRUxBrRjXnqNEVjUqJ
uy/1mOA/yw+a5f3Ul45qmmR1Z4usCCUGG44z+1Ec9hJwvSRW8zmaXBCls9kghODX
zdiqjibPGIjU2QnsrnLWj+JFLAke4Fc4iJXfouteysrdVrkViiIW+4J5udyJGrV6
o93UkaI+r9gGJha4Y0ZBVhA0k2C2rQA3R4pWbVpbhSHGbl3rB0Z+ZuDH/xUtwa5u
ZVV6b//TRRzVAV77Z3DUHggjLBbjwYVzRfuOKSw/m1MZX1RtiBK0dEg19wDJ0Zg5
ThECjCcFxwinhU5SoM9byiCyDoSdZsForOq1kBC8zNWjt7tl+dF/ZFN0UHW3rJEo
k1FKG4SMtkDRZfKPdNTxrIGtvVCppofnEIftRqgfx/gla2/7Xh8UFmUgPV/qPf3c
L+3OvhkT4Tq6tyyRj5Tm7KhcyR3sDoNQAksU+UMNWMiS/A2354MvtIMA3qKKk5ft
lmbNpXnpgTSBPb5M0dbmCAiQxVa8rV3PssjRcZ/J1rCgSt2Pj6C2FxNMEodR28vs
zuEeXfbnnGfJmjumrKyYrDfSTkPY3sBhjEsqnsnMVWKWPboRiaC39mlYW8sz6FmS
VL/H7KfrGYVaQRdBxiNwUEX7UzQ+DH00fVJj8YM/Uv6UjdOtRjYF3EIppXISmm+C
r3eNg4mnIZhbyICDhBwL+xm8SZGB8VtGfQYNh/Am76dFRHoVXphkaGjvv05wnitl
Gf5xI0AQn7oceebaztCOq8SYf47X8F32mjYVpRsPBz3D+uRJYvAd2mssmeZXCQPc
VZt6z6YiiRKFwBK86udzPmfkl7gLbfuOmD1p2NOZNNLnQCZdUYRY1KcIvhfVDmZc
VMIFxwDDMSc1Dd8xX/3R2I52Pce6X5b7SfgtOSFZV+/iM6eltZF5dtGFdbL0Sp2o
FTcA9TLp6Xdq4U0aWeRvyO16sSDwEEwu48lw/0w8/mz1uK8QGjm+qs8zQbI84D2H
l172hbd665VzA3C+u6GQ+UFN5I4fYbv32mvSJSMyanBaZ7cf1YcKOPZqqtmqIDCQ
pRaoe0DsGzCTkDdGZJCC2X6Sj+4eR8kfAn+UFhEZ1HdWE7k/rj7Q7hHz5PcqB29r
LAF/fu6u/oFfrmAeG+LGXx3RwYoZ+9cK2DFm1Pfe2TeWBw/vdiwBnFh3e7FWH2Yi
ROw7WrmLZ43U03g/JNUL3mPkcVlbIXBohP2K5LGVpS5mdqIFsKZ/yW6gvDSIHFnI
Oc1SYDKSN8DuELuoBnk0jyr4VwFSHsLM9g6CmCN2lWoJpS5ttCqYtQABhd1+sqqk
IJstzv+6k4oPcwRLvhnzqnujUKHBJpvG7vQTfzcBnLEYqP+txF6yFZV3rh4/6i/I
AklKPpRHgaZWqDMq3iO8t3x1is3D5yiRUHskrJjYnN4ZbshMNMG42vH3EURvQcqc
hocKMkh8eqdUzPTHQ6wWAwxzSSx5hH9q4g6WHbdfILYKGJ0GA+JIxy1ofBHZM2VP
0S0UWqTd/eI8cf+sZ3jiBvI1fInUu1xYj+53Q7vNNO0aFw/46wzpDwYBPcMWPbPu
5wxDZuii/R2zfSQhPkIxZEVw7DMuzSG8r7aycQYfFIoteI6mdDq4frF0YouucDrY
FdsLYYmQkIETRCE+Ra7LxWWU9DzHeFXFvYW0DDFF2q7CpRTowCqz6PUmeGZ99ckF
mGa5K3ETrPGT8rh6luR9EqMNLIxaOFpogVfi2C+6yDlTrPokt+yrwktIgL/JKeBJ
1dKHqMopxNKTU9/NVsstO9pjPxMYpwq6+qc2ImAWoiMQp8vJw+buRh6Spp3FEws0
YuUPmdvPzfpyI2+vxfIgPQwnyftZPmuUyVmCqa8fMRGEBndgQcOIBSRZ+sGY2qGx
9uk6ROecgpJCthVvb+g6sYyfa+NhOg1wqWIdLRi1ow1Hrmbkvg+ZxThBgjohh4Vx
0q0SH9g+Rf5dfo/aLU5qgg==
`protect END_PROTECTED
