`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nveSEldD1dYhIvFal5k2fh7TWJCtJqDBc1K8J+UwIQ3uqKjDaTeTbZOszVyGPPdC
Amrdhs090Ybx9ccDcvOiAtaGrYBsgiakqVXbBimfzTKINkccoaituMsm8vw7sRoa
h4eRybwEKds46p/NB0P7T5CJmz98PQg/Ygf4nHPiJnQrnRRaUYgvhb7zAph6qZAO
kWelP8vgfrU9l72/B6wXYY8YlODr589q3H3OmHBbcvxHueSVMaaDAb5migOErdmW
N9Y+r/PwRlGwvZo9jDsjLiRbPSzTR+KTr5F+0EG6NYIjDDzHLFi6a9Xm6dAs0Sjk
7aQ22rxpancfqOh3DMrjAiyATu9BFAL2Z0xYkyfg7tgg+gkcvzysy3EocoFtE9wQ
hnrHvp62OIlctzvQJnbWk+FlE4696i2I2hPxn6jOqbW+FBRihvKam40SPXISBBnC
Gky8GtX734hvJ3bBZ9I+gRVBn96ixpLNuAfJMATr80TPlRSMDAWXMOVxFAJ5uDL2
wiZJavwV+3UqYWynMFFiVyyJ1tJ0zfvsP1/0nRxL4yNYrnxca8GKxSkl/uAaWCdR
KuRQB+iaIXXd+qzIUAk2lXrmDG0hzXSAA/Vlya8ZWKDycYeTLJ4FLCPx1Hm1NrLn
AnGm1X+OnqnGY+ysZL4/mFAt18kDcrMhAsSN1mU+4oNHyodknmcJDbnBybyFHWD4
IuZ8A53YoOghVdoL07mWssg7JK8kmsUHvZxv1vWXt04FTkWaoLgCUgn4BpbISEUf
xb9VWXT1B3sU+WxLDWV6xAchRuGlRcDvIv5D1NuYjRY641W1lVn4Xrr0mcpBp+n9
t85xEjqG3gKS9JMGUAZEBr4i1ucnvLQmZ4oJq6/bCJT739w8OXsuCu9wDsUxaTme
w2qHtbFKeqFOJ39DOSXjx7QrN/R1KWqoyWesXKzlstL9pf1FP6wcd6nHOfubl4Gt
USA+frQOPnfLFyIpjU9pkrZ4/GaNNU1kpaJ5yDK1eOzg4J4GgEQtCXLWOn+Qv/gv
izcJR1oNLrC+u1GBPzcaZfYG/ZDoXUQfdPdrDw54vO3InskkGUYwzCVzo65aggoj
uiiNnqe+F54vw3vWcUQwKuzNgjQg6mQGhjbkv/Ygfcke9+o5wLoen+HpMPCs1wZO
`protect END_PROTECTED
