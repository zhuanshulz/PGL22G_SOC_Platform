`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zltdYYbRYDkumb1g5y2JWsD0/EbwgK1dvi6c1BpoxkzBvYtnhp003Pe9XkPVJZIN
oWpJ88U6AO9StpRybUotT2Hp43ZPgyeJkUuG8SwQjAQXE9hRqMqJ67WUP7yw/NKL
Ue0GMrR9JUlv6F0XSgaMKxGYa3f3SWEot8OjeX2tFyauBUeiDA94ntkRvWXIK/ec
BI6jnb/gxgrUNTzX4+wtOBl25lEdV4ZF/2MmA1+JLByDc8Fk2EcJeqSpDdDnjv6p
6OBtqSo0Qe1L0dQolNBEDlQwWdhgR3azq5ob952GQPqEA75w7iRofo1OOam0aHUO
aSwbY+kBTHy4o+OXzISN4w5LE4TgwgwvltzhxcIFmCDZg1WEQGzwpW4ES80aNjaI
tnF3HaGte5SqoLDrx+S0lUBEik57De2yTeZp9gDafGLqFGp6zh98HQYwtfdgnNfQ
5e3g1fY5+E91bmnQARjdeopgNTh5lviEkaLrL8ey+6MaRlDR+YimOnL5GWt8oHR/
x5CDDjVbS5Tfx/OXgWOQtzeMgGhBgXKy3vpN9jGV5mWbRyLowbkIILaN3PuUwY26
lbJIvRm5zPYk/gyp3POXO7fxRAcyKpGZ+Wrs7K25ICxJBIpH12dmMDP9auk7afWC
vyXGgMbV6XgJpO25JaEN4UxNH8aazi3rbKIxT9oPipo2FQPN9osrJNJ349cnFn2P
mKMHpgo+qgr7pM1kNHzg1SeIB9v9nsmTsV/wKcieu4We96H/4hvZYC2l5FYjB++s
r0iRkhaqAk0uRECwHI4XwPzoENvOcOl27GUVKWQBxrP1lumWQ5dBrMwkiFRpq/ep
/4Qz2sWJ1iY3+/RTvrLXVFT+7tpMNK+jRAGlMDg/EqOWxCwum7GZzwDcOtFjkr6A
XQ4ppdoYO6BA/MsLbafx4JAitgMJphcLqKnzXf9613TGt06IoBwKDW+HuqbqM+d1
RJRI9zLcbEB5JcyyBsJhypP6i0ZLGiRxzHrtBcHsLtuohTcxY1vHdo3qDopYx/3k
smsJDkfRoKYKb3XJHgEsn+z3wze8Y3wRlF+ssQN+BcUECcKz8KOLuOTz8WE4dnTA
9WjtsHncY1rB5/Lx9ea7oDaeERIecoWREF+m4PRm+3TGZHpzaqfaQ36k4Htw57HV
0n6ThqkK+MKCZAIXqxQLp+JdhR8yuIGSMv9em22cj5bCBpTiq7OUeSyyYLXIXZMi
B4QCwkdDsrHXuyY0KtRhIw+WmSCcEZKMoOojqeqzDMu1kgdS0MY8IUSWR/FD3PSa
uQTVg8kLi+WgFaNBhvigitRkoWn+BGLzw7eMzwklo86LjhZbY9OFjfurLu+PqOh8
viBXCe4gt2yv2C4IkRY8saY50q99IlBXCyR0rdDnzj6v2JE+lmKjaMIp4DN9bdow
J/tD4BiYiS2J7DONpU4VYrlt6DWJ/VEWQKsC9ghgTf9HxrjaAnNfny81ruNO6Z3i
AMi6Ea5bFd//fACS/lNXXpOXCrC8NsZSIrR4HRvRstTmmXJI+5+sby3gwN4JvTlv
INDFexjAjGUmKOZvu0flg1zppGnk7FF6Jo0Gsxeb9coh+820t9CRr7DwquOY28Ct
TbeOu2atk0gftrXD5sRQjjn0BRvxaYUoBPgzeeJDhR84i0OhVZwbU8++RJfJN48A
xrQ2uuFvua1wUH/3f9Aa8P5EvyCWp1bDXaTH2mDTuJc+A8ZN3hgjNCCnGYHeDE1j
2Jxmb1qi4wd7E181nZtOohTMYdHCeOIPFfk79lpIh3EdDyNm4X/mEit/LoTh13Aq
IBxqS73LhUJf8820wfSrU7VOlXG/6XkEL3XJFmosa272o9fPCtLz3w/5XZeWGSck
10uxyEFGxN6jdxINcuAwVc4aNDzoCQTpWfYfYfJIjQJDB0O8TkmIRGJA/9WWhnLT
UQnZvVcpsXcz3PJLYOX/pcXkpbNxdR5Ts8qmsaRAWBjzgBymLDZYeHwV/TP1LmP+
+6B2No24SoJQ1kuAwb375ks49JR5k9LQUFwA2V90ni8ZM+e65fvnj4xgr/IkVp4J
/5PodJM494M4D+cixiqTxxpHIl+frwhtpUqgjkIFX5jZAIO2ehVIJR63woPnEo65
flXDqShQVQ/Na3ku0cJAh7xUoWxpw+BbQ+0AuD0yny2UjUCHFB/chQMIOagdjMzi
WGN5iuIoK3tTv7qpNfSTobgv25kF/cuEuucf/cfIkP2CbeVnjnTmTW08a54WBzeE
U75paNa8BhMwWfMzTfBKb7heOVBCUQOSKT/F8VgNLwx7dBc7zz6DYeRd+QAB+J09
QZJpoigNM0XohKSyL+BGoKIOLtMgrVkEdASNm+VYdghhAlI9xhgpb3EQBiy3KERI
L3bHQiZWy0v/YuBXoDlNfMpnnJmqzLN6AmhRgUHJgfcIlfTl0Ut3qZHRGAI45IFJ
kbMLetnA006bHuWl3xT7Esy7FK1iwSQTgGpJ7IaKS3P4t11zzCZdc/kw7GlE0fCr
e0C3JDUEhgWA7DCDhSrXUTp+UjLgoIPLRSVLjz/MntmMD5nBkE++ro1HucVBa9iX
xSqChwZODMU36MuPqkPw9YjMn+hVghObRL/X6KGcjeg+cAaPq91OZxFr7pBzaXR+
yv7/UQsnPXwrY/c4Ff08K7e9dlFbnyNzN4YnBA0SGY2qCypMWsf61Tvo62z1r+Ng
oQ3ug+ApiE3e65FMpXrDESEs9XsToYp0DReu0czkTX1JzoJ/PYl8RJqrApxtwCRb
ALSNJs6AL++wvjuCC+WssxCOMR/rtt6xHyttKu3rfRzB2+W4zfmzoSn1tkemzgCT
Sf0zostdeNyEdgiQxIlS5Id8z+OAwHbBwJW/EtCYylnHNnr7aVNSl2YL/9fqnYJn
8oe8kEjNPv3NcoXW0OHpujixJ5YUCONn7ETjG6rch01ik3sAwRiM2bDX4ARWrDGA
DzGMu+4U7Hv1e9DyDIF02BD6iR0I4mm2gDcxcMlj7SIABQBQLkyDhBG049YA6mo1
otWXnDiOI9kqaZHPG7V8G3uf2ae8hBpv1a+EFWkUEg6gPbIVy9yx0zX40IVbubHU
b8bHWXudXE1HARCHwG7DjwVZZYTjtuESi91YQDF5W/ahx2wafbkBWYpEJiA7Ahwp
WGodIhVK8vY2NVXrZ7eiyMyetrfhRzy3zK5dnr2NEEY8rIOSpulIP492mF4R54an
pcgQhg1Um+vhczivbq/io03MFeKY2otpZDxIg+tq1T8ow88ISVMloCT2j2Joo4tH
bElRiILSvUXy148WurLKSV6BLIEXtgw8Wb2hkntCkD+ZzoJzbaIs0X3FldwTeawd
t6dc36sztKiNErECvaL4pWh876ZtGfm3U29hUv3S3sANmTVy2Z4Yj5VZuv81Xmkw
Prp385koC45J+nEhvM7rLQS0lKz/SOgU+f51PCOuaZcc9TsjmJsmJyH4cVyY6vcI
nmF5G1ADtWdicbBvc1VuW4hLhDxal8i0U4VIOo/PcaJU9hKZrA7fgdZFifkXPBW9
+lRdfcIj3qOsXMZo5RSM+5sPppZuC8bJixjBmdhcQ+4CWeM1HPrV/KN7pKp9MlzW
K9zWMhid20g6JTDRzVkC8o4gnUQy/r+tXK1RA5CO/Y4JAetmaeSEQfwEYXZ/MMZ6
d2alpPwoW572avmbd7M/TD7+X4+veatr6Ha/uTKATZM8GogbHHkD/uijAf5dy4bE
TuWFN0OINkz4/y1BJpNBzqerldS+oBOEOVMy+AW8OD1K1j17SRBim/pwwJEKN/zY
hQNChOhHdgVmwArtPKaWzDU46v+2xRD5AG670dF43NBffjd8IhMs0u1nS8vyASmO
fO71tE/8pqmSmmA+MDEr7tV+NxETF7gOt59UUlZ+6WsgUlN96CtkBPrmcXxhYeKr
ouDBsSwekBMFbOY8MGY4Oysr3hgOWI4WNYRuOOrqZYIWfVQ/Wi+7nAQut9qclugR
NH/MOO9X1x5MlUaR1BD4airb37nbqTHhxvstA60oK90+jxSDUBvSsDnK36EYee75
8hJSTNIVZEPp6c76LdjDFmHlJ5A5fVA0AZzfk3WUO3x633BtBun3b8k3eHkHpaHE
5uNvz3mUsjioFgpvlVFuO+ZTbp/Y0C0O2g0bXUXG6bJ46k2JSSVy9LGkzG9sgGV8
940eylxPwi6DYICJiV5X9d1sZS1r36t5LeYh1ITh9jug9u5WBSgcgxc/pK4k7M0D
kTdbnrCcIo1TGeLp/KbiOIWfgLB0yyGhCxJJY11InxwX8dkWyUhNw1cOQ07YMtPF
8Pgfay7dpu9mvGWSiimgniCP1ZznrU6ODX60ISmfoZbTNFk8fEWRzrlub6wKvA8P
mZs/MCh4bdTsXQC+i7a+vKQCAjk/AgGNybsTbMsUojOVYTrTqPs27LlPnwQm8zUi
ikvH93niOe/e6V4vS5ZuudQ8goUSEXrzCLvHOSA2EcnZWPwvUMpsI0zl1311j2sf
K6kaXWC0oKVtWUIzrJnvf/IFQHK81RM6RpmwzKVBWZbQYcMxXA7tjSUpbzS6IHrE
omm+UIjtrm8Hh4IRk1ocuLfoCcvHASQoXmmv778dbDq4lTq0ZS+qRct3mHLKiqpK
IVeV880pCJFBE1MLyiKEyxkDdC4FntRWDR2pEmk6pbzlF8bF/i1uSLFtg9GM0vSr
bYGeeSGsMeKTnGSFMv1aFpceyz7XHgRvo3OhW0E5tl53tNDn7jX0vfWP30jrce89
kdNXA4k95o8SyU0tMQ6waBryNN4qH5HQLqQJWQAEQdrO5nYqlMJW9dXBBxKJh+iz
w7ntFPYNonR1QD7uFtgURM5kbvh/XQpgV55brNnGsZsQF6okHZ8y8dztSTQoA+j7
ymG/YOAjf+GiuCLobwic3dr+32mH4Z74o4FbZhcBY6+E9Cbj0frZ0ILuA699C90v
U/j5sYYYSNJIYQCyr1Db2oDhO3ZNZxI2LM7Q1Wu9GjwRwj3BL7ylyv6OW+5ZfN8H
KXVsRHIsbGH4FJxaHBE7CA/NiFtDCIE6aFfza0XYznj/R81uYSuTFQgLJBVp8+tv
6MqAkmPLUCSolu7D/r/cEO2quBhm3Cu3MEW81vzMUpKdLtg5ITci420miwKjtXif
s9LSMU2mZvfb1ChzFF81bHb7vq28n32q8yhxoYWkjeEXylP8QFmr/feYCUybkTw0
PZiwS2Kt/sKUr7w6q7Q6c0NyB/2AN8ba3LKgMTWDIN0m28quhi0P/y3R7S/9i4bm
3p7Js2BGRZOY3EPy+byITd1AjbHXjmRa4bRM+XKMn7qMX0GB5ToyBb6Hr2CWmNqI
J7MWYsygTWxxesRaxluRurkUu73Rr9U3KM974IMQ5leQLHsvgeJbH+sf9vByE4dS
0QJfgsR+i3FktJ8VzM57Wb8+wTtz5vHp1aLAH96chEkDGX9Bkd7DBlKu2x7z5Y3m
rMU3WUd8vN82bQL4+HbGuyEbmYys8dY7KpmMbIAB77gdiMr6zFVgV5ZuWirGM4xr
qa2uV2dHggxkoEPcoGfZwGR01VZWeRUhCRz3Ub5R20K5TSDBxq76Ogh5ppX5vM7a
4B7xrnDIMip7/Deo9Dw5M7IF1go7bA5t+ke5dsAzyqReXV8yJYRGAu2eP2pohUE+
vUUgM081dQIs3b+FLLe7XWadygC5WV10mffcOdJAv5NxTXorEWOgKfZXwf7AVBhI
FEQyaqMfF4zs6cBLMoFkcP76Jx5nrI8joT/tMsDcQjUvoByNAgXvbRHlL67OwJ5w
3VGzBy5fb6L1HrXy9ysTIKS15yv0J2RuMhw1TUyhebpvs+v2y2ghXM3yTZMX0lX7
TpRq94m48NJ+y5zVmYwIlrfdFEyBxJ4uKmKb5jZaNR7cMWDY9ZUHxbaiXeGpfN+P
/m2AQMTY3zm0U/i1k3VoSH6ZmyDvIoIvS6vJhLD2ZigkJj+EwHqmV77r+ABMVX3w
yZkq6nOFpRrWHDSLCrDC5Tu7YqmUhVpSBNV6IapCH4AelRYdISmT1f8t+JNlsXSJ
ALeARsYbB0UHSbyHqlt5znEfWRBth6s95pvgMssJAljrpgWfOPjiht49iqX5Zb3d
cl+GfxnotMEfe37BwhmY83asj5xqBRnlR/f6IaeXeIdtZbLsPOhHpqonrQ/6oo15
gMil2PxZPNAdeFpbmS19Zq2+k2jFUgmIrduct5j0lOrDRB8aW8xon2/XBsvbYnup
/EXhQLz5n2KT+KdUXr7Qjw95G3QFaX5ZYIEaZKiS8a6IMEHPQM85Pj/llAvywI0N
FP4vFiVMP3VMSjNCH77deE7iLqqHglsF5+jgoO9nZQXOq/suDtabAOhLKBrLZoD4
`protect END_PROTECTED
