`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FYw4MhTTFIEhkLWZ7sQ8Y7pmqilDYtjkgUlOGylpPQjPelfzgRszTVVDbH4BCibD
i+LAOJpPmykonsDMZneKhPrS5uMYc3qOF34l7TBA0Q30ngRswv09+PJaA0olpS5a
+RtIuCNvd+yAOaEWZPFobYXQxEu75EhkTQuIxMeOB8qiEPD3AZp32GT+P+vQEePi
CkMFnxWwHVB1sxJRVXI42h6ESN3pCEi4BRm4Z6G7W7rDKLn4G2haJZxY191fhS+p
xnuWif6EUrJBh3Ve7ULgag==
`protect END_PROTECTED
