`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OPyJnjsKCQezlunNEKg6HCvW8+Z2wivwpPGxASBIccdzTMLzRHXecYW83IJNaL09
e5f5pEIor9zmQkWReRK0MK5bMdoOe/zhDdKgMp4O2N1Y+/XPD8z0WBAkRf95efkA
a6FIeytU+WPpjHs8kjh9lTYMK5yWLRkjoYjQ3jEwLf+UQNliJfEl5wjZBVABs0cA
6b/xp39MXEMmVFQ/BQulGCXs1Tl+ZcQ/dQRietk3c7tyoLsiHilQGbF0wEUNId5K
eFW2YHwshe4JJLh+FoPGkQCzbFBwOUqPXhwKq0UCtiU=
`protect END_PROTECTED
