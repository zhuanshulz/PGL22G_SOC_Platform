`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NcGzJnpUncIyBeSVg+HPx5rosq8rjg23bRD0iXmzX4SdFgrMyEXuTQyjxo6X2K3B
9rzXKtjfBeuUzAv/xQ2k3gptnRprAHi2GUrz5ql/CU1eLSO35zUBw/xPMdJ7kqV+
CFA35v5juM4yma7O2c9Hz4TssjDCflYBIAt8Q+aEEBx+O7OB64AZprsV40woZvLh
38jAV0hDqyutDAjteUV2bnhxYOSJs48w0WLwymcfsiinjs3T0Iau5+kzONTMd/9w
JoN0dYZeCQdTItjplpggXkWKovPi+X2B7SAxXnTeR+OOYPMWp2ET64Vm582mfXLX
f0JQiN63aaI+tjNNBINi7LkqA/ZEDkP2D95+app4RYuz4R1ZgrCCEx5aEPWSJwzV
um/D+W+Q2HpSzIIEsZRgO8zFcMLutcMb6JlJfU5zpFN9EdhgtvCZdP4e700C4qyt
p/AlNx3TllEIhTm5aB6CeUcKqUwSgD99pJT2m2CBGjYwMn+zs+BkZY8JDeN+jCUo
XLTHQ1b2n9cQza7KTq6TQJvocuWsCngEJoaiazOlqedSLf34TIdxxQdxCi9s7X2B
6Z/EqpcNy9v3zgA/alc8GhZSw9nZXXipifL54N2viX3pUhdCuLWY7PQA6vZ53Br3
VzLQaNCTrTEP8TaYn0uSXbypEDtudMwPuOuINxU3TOnW9n38Vhfbfm/2trjvgoKR
`protect END_PROTECTED
