`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZxkWYPCVwI8cIaHK58NznJ6iJHiKQBvE+Y1ivpDy9KOeCly3HrAQeuNwZ5aSVkh5
ImpEtKKfOjDnlIqcg5QPILhQb56GEXUFZvxjv99Q0ubQ09Hrf5A73ZQgvMKEXMO/
SyRl1EEFdwXAHp+txmm8BJ3Lxvy2FIdssVc52Zfv6SJTaAEkZzTPAY3QFHpy7nHF
eDWVvPHIjlWC9ODFH9aiqOkKLz6Bo+6mcBzZ0AYN7r+AROwrfU5p95ADnZoLU4Jy
QEIys7DUkFHTAwqYBAzLXCMbeR2zKI0z5Z4BAMrJKsIBgMx1pwAHCms99mc2z3x3
Tx6rRuajFHh6RL7mp56S9jM3+HohTFMugxYIrqzkl8Zm4va4StfYmfPyaWk5exOS
B+iGGqfuxug0EO4YlxjSd2XXDWLygXOMku7Z2ttwLXcvM6zKF9Hum9rqwNLRGJSm
uYvaJrAYemXaTx9+4qcxRQAGp9qlsInpgTf5oc/+cts=
`protect END_PROTECTED
