`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bTADeQpPK4bBqeFKtWqMu/nokBJPLNOAfKWdDAcjWN9/W4NgohuXWgHvcJUWWdTG
mrMyGT6IQbVjw9WSav0f5PuAem0uAEAxsRGd7mquCFRjwuM/uEHxcratk+hGT970
xWh1ZUunN6IRMICdIyHZSqM8C2nCD84h5VzfPbpnsTzaTWhxHqdY7uFiE6yaFVXv
gyr2Z7c/Mil1tcORY/Gd+mZ8J/eys5ldGVIeQ04kiR2ibS1KCd0a0hFN4k8TFAC6
KNE2pVUV5rOQMZFmeZUH+7nGs43rrYZqE/BDy967dVCLMisOaR3IDdmSTFlUO1kI
geiPZDzEvSRQ/CBWwqKDY2yH0l4jPJkyn3YwLz76JQrlBCic1uuhdRFH9OuzagZp
K5LHq88ndNXxJVT3+ppHKYxzL4/wXfFnouEUCPMT1XImeQMvzCsM+XO2FhBfRaRC
IBScH7vmFvaRRtZDjos4k08/1WtXWZ6KcDuCpM+rRT63i/uU63q/nmst7g4Kvpka
vxA3AcKebm6cfxl05+2iwLDqv392GfBRJwyLiuWMzogZd84S6/5h0IQ6sJYqu0I+
9qwY+mwiQj+AQ841Vivxt2ktUHPAnGyEKscuMNL7GWXTTxZ/HW+Ksc5HxkTW25ig
iZb71fDVwuZjDP79r6WOfqNHv4g1ojMK68pOP2Acn7NbpgwaFJUkHUFETi95ba/0
QsArlannNF52aqc2ud95TBIIjR/RPSpFka2EDYaTxM3XY/jytjX66Hj6h+HjBZyz
w3VvYpsS3XXEy4EjKrPoIoRgCK4snssnWQMuIlB8FQ4BlC7cV/Oe6nAl5gW7ZojW
SrOmSlSa4PKligF2qTHW8tO9LBP3AOotn4znzIXTfJ6fAEf+5xk/40mG4gdI0yX9
KzLrwWE6pQf3cTZvZ0toxnPQE7ckU2AChcdUoTgE9EiYWGm84Ohf4E3TCepFd0ii
04JZG+jw+U3Gy1igtRBRk20QvXgXecelYMvnVQy9Chmv2kdjKmXTPTmBLOb0yQPl
fZvxAILXZnKGzNk+e7IHz4IUKKhwap/T771J9lHj/h0V/IfcmIVHEDBto49gzafR
So+7ni+OcI5/v9uh/gGA2Vx7B+fcetWjtx0d444UInZ58FeUPU2h4JFsFXrWU6Kg
f6Bk7FkjY1t1taAFYlStd1AWiEMKjIKHokIwX/eQDl5wdsyNMzNcZJTV3lNln6hg
4Wpq+qRSSV9/pG1KNBuNaKwegD1S5+Qa7E3GS55p5jKgQnpLEhE9JllLWS1+L+uQ
91e5YqgN5klC9F6m9X+9fdl+kySnYxoM5mmQ+vLlI3NhsMgJb8UID+/6lXAU6Da3
MG5ieywAtH/Yenxto5RrFUc+XsmkdSZkWbWFJXjlatoBBXEcFgDTWukt8wiZqW8L
yusuQNCFWCPUMSWT+5tppMpL1UH/THx8s07uJlgYYaH9ttUb1yx8s4ihPJJQ2vGM
/KATO6/3zaygEa59MEIkqooi+XDu8daRwM/0hMdCAiEu2o0BBxZMCX++IgFP+FzQ
2Tbc9Mi2x84t3GxeI7GkzGWXDgaRdR5lRRvta6szMGkaS5rZoSm8252WunWYcDHT
GWQOB2f3y3qucYw/1k5xOC/jVPyqZhAuy0J/NiR8RCM5uNp7X08EL1SjA/VgbtEv
fbGwbJDMUSh6OVBFamiOLOY4DaM5aSESBxDYzUzlUaBF34OmVVnVeBUzfyEXFRiI
QfEFiLp3c5HxujtC6lcoj7Pi399zNYxJb4JIQvMNX7TKoXbYUqo+k67Ve+21Sykr
UYrithaxVQbVTqQrLTws9pD8pMvo/uneaxDCCKCpsOuy9p9th6LHOgck1v+2dn6N
M47rGtKSFwG+1Bj8tGZ02sRlz2NKwDCDagk5q0XJ0Vaj+BngLYznRt/HEH8S0VK9
oWbS3MPXXEW9Hp6QXXGMGjuCSv46ve/0aVodWTtrNRqaeK0uAT13kKhatqQbjkee
f8xKvt6DQ+bpDPwC3dtP6QRBxf77M/EMYEm911qVJ3oFtK60sBW/YeOFl88W4qd2
hQ/N7Ae2NMbXG152M/ve/fBzWSEca307tMt07sug1nooXMXNQEy9ZVKMqlzewCWu
Omlt6uXWf3NpJ9lPrQrzhYkwGrH7OVr13uhFvBTOR00RqyZnVgziBFhC0VX4oNgE
tjX/tRlRlteelSO93ojrhIijZfWLk8k8+b/TDlTul6evU1kkq5N3JXQoDN3VVoQV
PuhIJSGOxJR/9DMRgLqK/S4oABuViU1ftPgyBzMlT55QCO19Vmqw4NQP/ktyadmj
kscWKWkFyUZmqc/9X5AubJjBF1pRp6AQUi78CfqbSg2atWZFiw8Pjk+Byo2FNt/P
CxoQgBAXBsZBLqCtRv2Fs9ZBCj1OiNvdSjlUbmePbFPfs+pSClaVF/Q/gQ6crHRJ
4w3ifYcg9MLRVg5c1WFs9Nbil03cGky15CQVfgRniKxJkBNr/Z5gNbEH1u6wvHkO
sVMyIfgrptF/+c51ub4kFwtzMal8jaGlP2PFtk0jl+/1+LEj0k3QG8AmHfIhnFiF
WdrCqDU3K+VQG9MuuUBRrQo9/95I/A4c5VeXtqF47fRobEWEsGy7XwYXfnMYCWC3
`protect END_PROTECTED
