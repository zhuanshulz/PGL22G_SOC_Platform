`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mvqPnnfWPQsRlBMOQp98BIfH4xGuLmm4g0aINLEVf/7qfhKLJ223twHdDflytf5W
aF1VLiIfJ4paKKKQVTvAn5CQCn4ivMjZUwnQz6SOzFT92pZ95yTOvQ3biTANM9P9
w+mUWF94XdX3VUGlXx7j4/DE+cqTav6zlOgPUk4HGrue7nKpQtUJjxbAjQ5LoCFc
KTrUTwr5UROcrw/djob1a7d6wJQ1FTYHEI8XEBSBdYiwcDnw9Ml4Pu8auusyrrc1
c+NajUTBoMu3y7YYR4pLBRi5Uk1edg/DZsNoKBQxo7YvpcxbHv2e9nHXgVhHMNNU
XmEFNI58frzPQg+s7ByY5hP/sbW93X/PkKgmMIUJ0OKLoBQSnbKa5yyRKcOhytfO
Y8LAuPEbBZJBI4yB1atyzmJuaQ3UGMSJ8vbVwUYvHST5PYEXjQpXsdpx5Yi0IBs9
4OxBu7pSxi8nHoPEwNVxf/jW8AJqQqiXranHesufMkPVgS2JY2xjg2wCsP3B3gSu
YAkysRUbGhADvgYbjG756hw7gTUxbwHdOlZ+xgGIJgTwH9c3JDB6fHg1Z85xlieI
2n1xH1SDQTrSZ7qL4xKU/qF6Eu9kH6sUBM3yPmUHl+8tU7mLExXsQDGSX3lRdUUh
RuNuHsdf2FmSj8WsFmjXgb5d9W2N+8G8wOJS3fX0fbTyFE7pixGJ3iKPr7VsnFCe
3gJnqHGI8WpitPGlAsX1/pnrMWGimLPXiDpg+e8TVkMomkoF31+WG5ykNmGM0YAV
+f9FNFy+g6eERt+cq0wVtheivUdM0L8Hkhe5ujWAEKPI9rkjbTYQQIGxrOoiT02S
QY/mn7L/7VMihg/40wlyl4Wk6By+MPpDWNghJ6XCFOIUJbUfiSQ1QECRmIjLmtPQ
`protect END_PROTECTED
