`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l/PoTTq0BgW9F8eQhxalgcT6sjREL9ztBgSoCZY9lmpIQnac8N4Qr6uF8WqzoCMJ
UGFZ9KWSHPzXlC6ep2/zoLqA8arUjRJxVQdaOYK2dxGc7e6obsbihaqfBPwMmdmb
An4OqXjkhBY9s3bIaWrQrlvqySqCpofeMGWu063lVJylX6dHv+MXjMtbTeY+ybhd
Jmmy/uySWYM8h+ZmJ+YNVbkCcg8tNrjCsxAf3srapg7P04mIqVDK0E0zWAClySLp
dGnyQxBYtfowxkRuba28kwwiY6/5aSvL105uC3iu+yaVlac5Or6h23T3XpoC8Z9t
cx8CM+l36dYsQOEBWWES6ah2k6N/KCaBrJKmHiBtZHbZ3IKun5VRyRinWvJgkZrd
QXWjYqiGF0KUxU+0wVsal5ICnvosjPaxA2YpbrpMzi7gNrjwfTqSroHeDdt2B+H+
`protect END_PROTECTED
