`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1Dk/eQ5NBfZfr4jFpe9hIrM0pp0eghyozl+VbiCtlvJqXRKfQgaQGNpmSaRn04zl
nv+5x20I9jDuWR5fz++nIigdCwXaSWD7+L0lj4/TbkPxFGuPRrcNpZr/a6NL9Y9W
uK7l5mz7l7ygGs+fr7XgS2VGQUY2pnzbJM7sayyjVD77Xo7WoAPCzvqb3xtoau5G
Dc39AGdvItygI1kf/cyVHxWjDGTNI0A+BwbaYCJksunCKcxbWqurq2p3WIgEUEyp
uKmMXWjUqu1vDUdiF9g+KYr63RKfX0l9UCTjo3Y/tVFCmonnAASxjWmeLx6oE8/Q
Q7ADvt7m6kdLN3nABxZOnbObPROFuJ79RBhSv1elvFaO9sf2fzX6d8dLAcAuMU49
i9CXUtc6wqCtEX1iCyHw4pbz8s1/eTuEV5d6OUWY+bwzKWCL4DZBS7ilgm/EW02B
uz4gyJDXwJDagMqQLDlnwK8RIez4ZsIrsLvOUHm9jwKGxYQvA2ETbCSUe6Ei6Efy
TV4dLFk9k+t1+OVXHNJStg==
`protect END_PROTECTED
