`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6wh9p7G7NXfR3zuHrIo33I+uoZNm1DnOluHk1xLtueQfRZNKAnssihmuIyR127zp
9vh0ENhhG6BqDqVdFPiz/U/KXbHg7EvTBt9yOzUTY9lZXHDbNbUUiZ+wzjC3kne8
vErZwICvHNG5BlaAvseJGK2O7mBShyDROsMLjWAs5YVORFzM+QsOk4D1OwqVjXsb
wSN0iWBT6V0pXdDVsvzhzYZVT7ttuOGhaTtgvheluM6ZBSE8N5FhsRBcj2BfAV9F
77SrUifBvApc8lw8y+IhMrtfw3WWDqfkN2mlPE+X2J1ECznaAm+E6YJIFSZpKVRU
cZANPNiMwRNkStf6278179N6wxsYKhXBYVf+cbU8MjfAhRONQQWsF9oUrp+ItSJ8
4YICSOobs3aEsCkU+0Lf7apNYut3skM9a8hsJHX6AV6EBN7BEeZOVISk9xT2paGA
xdZ9Zm6KUnufDnPGi4exI3ZDWjouGb8Bdbqq3bMjMztQ3nIuFVrNSfI7W40TuTpW
xe0LEG9T5VRoFv9zG22EeESJ6z4W2FdMz9MOFBn9G78puWhA7u4Rzx9KV8HZGBbn
DZsuEB00PKbsglnW7u9UIlHtyvoev3fo8pTPCZs3AwvX6TQgc7JfFnP1xyT+Clyz
HqzCy6256pDzE3Cm5PkjkThsvX9KYvzlbr3EfYY3BzhyjW4200fiWSjq057Zlq/d
BVgevqKDXcsp+6X/NvwgS0Cm2mXIWZOmOb5P58TiOeqwoCAMeqm83ePRwEIL8xp2
er0ZUfRRIfChoklxFlw4ivMd2BGW3/FvS24PO7jgmug=
`protect END_PROTECTED
