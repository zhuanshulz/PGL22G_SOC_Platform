`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AdMc57e5t98j2hpYoV7DXYkqYgnzRdZJmAPDE33E4JqdxZlN8Yy2eFk7GyL7T6MR
5WkUl2n6GPI22q6gsWExp0dS1vNlyEz4D+O29VCpBrxRCO0kD7GpiY4poUM9OfIf
9VfV1IW4OA3R7QcavHOm/zbPrsRGpKnQ4hra7W9iej3nDDjarS55gg/ovcqYjLR0
/Vw2B8Mw8ZUpa8pMj3u3maBbvCdRsdt/cRdAgwQDcMgaUjhUHEUEW+U4UGbP1knW
X3cvbw5WSvHlJwP3SEyk4sWBpYI1qGcRVCzkCR0umjAXNE6nzhImt0DAceMQiE7e
zF+LovL3zppZ+pkVuVw/fdYyi4wo9QJxb2mUbcNOghdtphB+Tvxde7hJ3oFZ0L3b
ISjM4PT/6nnlGxIdKwMA6A==
`protect END_PROTECTED
