`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zpWVUCol5zRBSZ0qB2+1aCPx7VkXaSih0VAfH4wJ+PxogwyPFY2Yp1lT5TzPAPmk
zn+34cjt9SvdgD+xA0cdbTuyVucNgdVrrqx4k2P6OGs+zErsz4vRJIdoYDz1isBg
rjdM3nHIzzMeAo2xKwecptcesCOt/ff2qwhqKhYM9rgOAxeN18TTq8oluUWGKjSS
NRNGclWJwUCV+lx6ubtB1p8n5Lk+y57X4bdKFT2SUkex7TNtFrFqXFZ23j1sHWPD
D84EI4NICsmEISzWS+zlq0aJjYExFsejXNt+8K2Jpz3DR+jfj3AQUyla7Cpvkopv
Zrfiyz7Jf9YeWqcBZO0JVZ5Ws7rxOPmn1jUpaGQOwahNUBpBSJENGvGpIY6YD7Eo
kJJMcXUeloXjNbH5hrKqNRhHZYj6Oz5lu2Y3YRMZaR0=
`protect END_PROTECTED
