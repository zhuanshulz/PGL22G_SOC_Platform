`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JZzA15VbHFthlhr3Y4MSnPG8ItCavMx6lamI3cDEcfxTRE+CXEQDaj86Oi0TyXZF
+Fx1f6rdYfQsVlKVa7fOEkzpAp4X9vW60y71PEy+YCI5ius+HdikYByLe0Q9GAkd
UyYF42k0h8C9AgPRPGtcH2ZmlIHBG7l4yBPOfmD/v/RAGN2FgO1TV9ODmt33/qGi
KuGXPMix9KqNz0i5ec7Y4dEAOZlJIGanmzUuK7tYEuZJfgNn6EQ373VcohQpWG0s
OPe3JD63aYALxamZjV4ZpvY/q3+qhuNmujZdownj35oPoSDviUIVIdK0eJw8RDeW
oityzTJiwobtbjznMU3wF3RV8x127nfJwn1ozu8HElYlp7Oj6JKlA18XeLxrsTuA
DD6V1aTEspVQoF3nNu5bJA==
`protect END_PROTECTED
