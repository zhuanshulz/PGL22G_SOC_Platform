`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aBnzLog/kEy7+oJv3MASxqfXAFphdt0Jq/3wYfIQuN0UlZG1MkynRN80oZlwnOMR
lqldOosaiugS9FBSQPa1EnnHw2e1VaH0zSP0KNlHVT71UTFIzCSpOvc6mHpe53Vn
T8Tttd1qwsJdFI/QySRxWSJMMEP5B81vmjyO7oJ4ibl7pn+nsRISAjdMGqH5BuEz
WUlCobdD6ftgGxWgwfrQOvWpo6QMYGEgGISImhDTfAbB62XVSYgkJHIT4Lq2R6Jt
9BjuUtW93bxrYWka/sPn9fimS694Vs8zaptwLkCHAzm7dEhZ7L3nxjyuPM2SPh/4
I69nK/iWFg50ms9CbTSMWCmKl8USIni28SSlt4ed335Oei6kiN+MB8Bn1IhC6RHa
`protect END_PROTECTED
