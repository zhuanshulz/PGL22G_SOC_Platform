`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
90ZYldowCFYbeatOt6E1zilTZKwtPtnlGhH4eR/v+eLwNqWaSlC08tPmVLILz2s7
UQThY6gl8JYbqmK+k2FqQO90jfYAQdVQ3gl0gJeyoB4b+uqdLErRzuxYvEbhlTHW
lEC9shZGZGO9FUafr6tafk5bmXql4oA86wY46X8l8+9imPYdVrMyKlk+MHONl24O
5+kFl8Ljr7riFK3zBeogaKLVsOOxQGyRsiSYsG4deODD0a8CHbCGakpptjmtnPfp
bp+LiYRjljzkWmqYaaAi65HnfJtaGuA4CpjC2qPgJ0WQ5yc7MkhOI4awq/IYXLBX
f0hFgZUg2JuOx/frP8waN6qmR9dV8A9bxzwZ5sn09XL+ddNAxIDh729LdmYc1B+u
5oxTd5q98FhgkNcutJI2yD4pBOWP4ZGecESrnxEMQ8rmCgHV6XHQ2p/8BXhAJBHM
w3yqhDlE9mIbvzGkHNCD6gWIg4S8I46gOyEbY+ErVk/0cSIznGy9lgaFI9IdFOWy
Rze/By9/Ujyv+IHKO7RJAaixOTL+kA3+55Dtx0Ipi4inDvnW54FYUtBQWNrWmR6s
wIw17kXzKNxll0OLQjw9UITszBHgHY+SxGFrV21+CRaC5liUR9eN6y0AfBpq5NHH
4ad5vO4qRt6IoytFfklMzPsiIS4hYSxcjy7qczdPkMpp5XHcwT5gx9/18hNDHgC/
bEOrx3gHU6+M1wht1vxB3QIKB7AA/L8G1r7KwzBTejXAFw0BFurWRnpBENX5qDqS
jp1qcsgamVHP39RRyUePCn7cR16/82go35kocOMx4SsXa2Iwpp5Rvl3j2/Pc5/zk
vLVIrZhpXMVoGvJ+kpajZHZq/q73VIVc/jFyydPb+U4uxlhR7BiKKW0brTRjmZco
C4vF58uHJjp0LBiIKSz5ubCf0+SSiPZ4SrWoZwqE3VMHuKupFkfrMocVP9E1DWDg
exNcXlPfMkfVxxUN38m/0lti8YXUWvMMJl5YoKPwAgvXsapby0JaS97wGg0g/cRt
f9jAeQEN7bzXV9DDxfeJCjms6dhKYZqAhf1dBQ3faLsaPjFW9cTke1Vaes7wKIbS
qF1REzLBDVnkjw60AQesrYF2wO4sohS5NbeRFGo1V5DByZz3XIjon4J1gyyymEr6
iPp8m6jDOr70iSEEzDpBv8TURS/hPEGnCvOlhLKpQgfD9k1DDcET5LVrm/0dXz0b
oG04jBUboIV8GGwqTA9ohW+R1zDvjgJmaMLd1e4OO14EUtolUTaUSraFpizEkHgf
w/KEHksiISACWfC12fJVgDTeIRCqAb04UXv8z2pBiHIArR2YjIwh4w04DVu/BMUV
sNm3r0d0qtSAWQm0iX+tRauZj2fQxzyi1qvLo4Rx0IqRMS2KqbVBGzQJpjl7mQCc
a0i7eTKmhTAOU67NOfoOg3w04tObeqHcaran5HzSq+grcn14TBcPG9/ANPQN7U8e
1IGslxv7MULpQeiAnrNeSas30FuIajEa//yx8307El1I55/rDLN8cBY3LlR5Ay2H
fJ6ptEw1VVeRFWAS7+QOPSUXbWpEEjgsv91bFozBxtWTj98itVX7YYIe1X/H7TXW
aZkcUCWnA6qzLysYQGkpMSkYLL0WAScEDqOAjXYjO29AbWQ26U6YnckTdZMC2YnM
cCeAv0J65qe5vR2vcid2rrp2f7jFfSfA02sL+jm9o90rK/IFu0+V21KWefsWKTe/
PxO8DEiZD3cgsyEttuuZEs38OnXL7ArUdFXrlSjh2zUQ8X93ZwzDAplIQp77q0rw
LHt6Dv7I3x7DLN4QToPzYE2zdxug1QK5jAgUZEE4ClA8PdIRsbxxW6EdQ+q8aLXS
W+VeQCxQM8ORPAQIMlGRY/5ca8yrLMlijSgAR1XI1e9hXKzbs9NVfxIbQRGfprfv
jaWInpl4+OpeiHaduvzH6Uk3cevM7wErKkTbug1yfKPPEHpou6lWDXhvydYheKAG
VpQIA2EFhSQOCPASKSnSjV1fvZnwHI/rAGrxqiIlubayXrxIaCaPvpxnz5QXZo9Z
vXA0M2DAuSNVVqR8JL5bP3vdtOXmO3wAFiTJMWbPlrM=
`protect END_PROTECTED
