`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w6b9PdeyF6fCYgbANQ4ZI0HkgQQOGNleBlX8aJqN5TTrQtfN2KOTjemTwWnA1qbD
VwmAG0wS8VM6vlEhrNQqLGw1h+SQt6iG0PW2u9aflLfve92//V4w7kXY888F3kBx
ihWlqYdsBIXf7HksiVDaCaiBmNexz4H2DW5A+7DzUvnC49ckmFVREY9Dd05NO/6G
G9f6HXPALItclJ4z8hL2FQXOXCE9VoHKGWNOwPnYBcAV+vLKcuoux6J6RNEiFapX
8kIYfrsDA3Wvli37uJe3aFQKLj3lyeimE5ppGDBZF0iwaHpNeK8+NhASdGXbwCAU
px1zPMbpeJyJR//Egp4W/c4Uj3u2D3Nisr+YuypuhhgBkiPaFdw6aQi+t4beH97Y
eLKXe/OD0QoRb1q4R6f/7uXukeeVrxXWTx/OeGi2cdt2l+KsFrMtbN6iTBnGNnCj
4rEIz7HPWkRxLBZrA45w/2CZrmINp2OalNKmJOsKUpkwIcGigkF3vn/CMS2wapF2
B7TZvy+CAbKl1BhoVPogAabjsyAMoOvqVKlJRZmDXU3+kXHFZE5JaYpzbYAmUURS
ly/laNavu7UH/ER1OPO/MMx7p6UPuGdsepK5o1WnAVGCVM+ofS8a+Ie/s6d6CsKf
SVDRdzdH3JGEvuH+/Abn75xXXtfkNx2A7d1JkJzTtAWEIe4ms762c9biU4S7KskI
HeF2R/xssbTB5t9F1KOcfQjYTMfgBre9NSd5lb3y2WC3lBcQ8iyAWnHKT4Lu4yi6
4Ub2lhuINkyO2kNDIwoKaiDOjuXzDqsrPH1NJEubNS7RNlHYdAlq5lZDLIa1WneI
`protect END_PROTECTED
