`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GzUjucXivmwFspdCWU6AhCicwLNENVyt5lgV+iEsgSfyZrlhRrFI0lm8I0HLEdLi
4C59nKKUWg7eFTR42tU3xwcFC8UDCWuFC3u0ey1b7kMkglKu9cqmnU+x6aD6+/aw
uSfDx2kF6/0zgp8JLaEI12vTRYArSEgPC0nkMSpIz32OOeFpC3kxFmjXRhW0Qxva
S1+SRLriL1WVC3NciVNVRicmC6kq8wAIRbmzBujBWZTe15Q/Mo70OmBnw1fvqnDz
pchykxKujn2c5fbm+XFOKrGHgBMxjT0X/4+AChmo4GTjtKn2bEhmZxPZ+Jl9Vhmd
nMnw+Y3qjgSLx+dsH0f06nNU2IloAEIrHT5iRdZ6rjrOXISB8hLuH6AGQjc+m9CC
7pkld4DQP8n4Jt6QQrUUOnacxZwkbsKKxUlvFo+Xhb37gjnAYFWptxcx2wGH5wMC
REbQu1/iHPoeFW0kZ+UCEPndm7jHC/Sm65+KGFgFMirWqKAO0ETVqthdazDsQy42
i0F1H5K6M3b3nvUF4D5zv5qBJDaJQsQIGDXlYGfin9uvb52+NoGu+HNBMuBigKX8
`protect END_PROTECTED
