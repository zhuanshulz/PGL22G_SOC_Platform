`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CsexnJq6EajMIHrFJefOG0484/4D4s084NfN8ni/NaGYBS1SrOG7442Sp0g9WqAs
j61/fpD+QN1bwPC6r4dQh08NLA2upiJ7JJ5pfm5AS344ScbbJhuuCsR39k3e7LiY
GdLnvdVlyfr4xPAzJ63ZZUmGTVv9SpPosM1JZdQAjflVXQvZh2Z3V7RXBZVzCdf2
W5tQYeeZXunY1OPwqvyQ1I0XrbSYdJgNkIPYCX/W0fSr/3jHoT4EW/SNoEHIN0Lk
MaQ3Qj+l/8vxY+sKim/jZGR+8n7oeL8PbQHquq0juOHGA8y8Mdy4aeW9yJuEm2fP
9/laT44owC8LYtrdT4VsYB3ekzigoRAnKfGQ9YSz0mhUpIi72uvQ691QRcKndmOJ
+KY3Ivf748hnJupyD+uf3fXHH7t0ZdqCmnJapJm3Pbk6zUqFG3iAM51dU7NZXwjE
JMBKMgO18nDwzCJKMkvRCCH1FoGPo4FXoI/RHY00wPVVR0o3PGJ0DGLU7Ooce/Zg
zetoCwcSwQh6Z0vhhmzFxinoEWK+1xH7pb0ytCPwisIfcQa4BcXiDPSlBZo/PRv5
ocybLGWTrsTekUmD77oLAK1UJKk8ToQEI1yHYrf0u8Yx/hO2Q7rJi9/DUwUrzz6y
eZRXTgau86PBMxJEAuN0c0ar9ZHv0XBEgWacJJOUtw3yetV+ZeXMepS/Wuuxcyab
lcXOG983gxgJLUTSbjW///1rziAwIAHACpZXMmVYLLDWVsW8FMAra2fTP7DVLixS
oTuSbMwRSuBtVdYr5MiNcv5r2hPJ2WRm0yAJhRFIqgQajjBXKBojPhRnwlwG8evc
FOGeMDrpgoCfsqKO8e3IzHIjf/n6hwmMBSGJOhrZkWeWYNlTGl/jd5L4dMhZgyBa
SJYXMFsYfcsGun7wYhqqXi+dVgmtByTq5hV3v90i/vpGDmNjEhlUAKEecExtvsS/
LFR/q900JpoEhnI8jYMeYLLiV9ngiUReD3Q+WEt8ingf5qk4N6H4oQL4abmQFuCS
ZCBCn7mBU3K25C3Mnnd0CSOmNnvui4FSudbC3zK52fsberDodL4lOaOiiWTM3KYm
+IMmZxIAia+/8HaPfWYFwYd3YqfWYiokBmZeL6XaQ9VR+fDHO3ROcs7Ib2H7j7RS
TaRhKfZswpGGecBS2e9DMcaeaoA8TLZ8PpZuy90ocXrt5ov0yUdNdmgx68XYUEtT
fl5wRmsVRoi2zx7iC4HvNRzIq+0lsqGRSayki5S+6TpBncDhp4vKLOVRLWnDzPxf
SM0lpp8gjpsOW+BEqI2FmfF6+vfRnoqxZzL6KaRcMwK3E/mVURg2tXY10libIgzB
mLMZIxSoojZAU4LgRDPz51zckXMaliToZdDFC3p/dfWLbKLJ6GkURQ1uvQ8IAThh
gopD5H3NGnLRXrR7fGjoNKvA6tVVWeCGsEa/kq/gSIS57N/uKW2efUJAYZ8rHU8v
XMvDL+jydhagvjm3eyYfSW8UEpDrk0glLKxVBVcWGrHVE+jWxvvOQ3LBuomP6HjP
vW1xn8CMAndEypn9U+PqN2wtB8IszxLw6Gim56RI/K39duZt9nRM2T8L2I4VZs4X
`protect END_PROTECTED
