`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VHrnkkLWL2cpk//SaylJ/HXXsLwy0LrrtvmhkreyBzhvF6gWaYIQARlH84VWcdTj
o4I9dGri7PvN2rF1zZPQMLor6ZdPX5c7hqzViCNQKmZNhPRKLKVxt96a0bjFn50b
naDRI8RkEBljujqxYj4MHOqsqf3zIeOXjDrwpvbfClz7N/E9k1Sz6qhQ3zQCUCRL
to6PTmw3JnpDMay3n7/4ty9v5rSqyoTWLbT5R8zKTMuOMNwmB9J3srXugaXXA6oW
TiJ58u4sKaw3YnjsmNSByy+vMMpKhihwte0zPf7g/TlCbxdE0TpCoohmfFzL3l62
+K+9GVwc3i2dVYTSpsWct9aN9z2KRyBk+p9IVz4cQ3RNk4oOQ7z+uLuAFsPyiGDA
eKnq38Ma+sDMoFdJKdQa07v0hpQwrO/4GbYCJx8g9bNdxqKgu4QTHqNHmba/6rDp
0GhD7vd7hLv+AyKXETrnjKAvmhdeA+B1vc3hwTYVwa6NEVgQiuzbSBReefFfU3fA
pnpzKfnh/UhS7iEcXZ/wRXbWnXohD7pFjBmAB/r1/GwO4kSxzOf85Y1D7tjUBEYa
XYSs1AnKLA9I6uZ1QVmev44riZ3Ys2P8XcVRCdJMsofjAnZSBFCEz03xYqPMNNqH
jpCI1anJRaKj/Ko8uhMrBHYQ/H+s+/GMZS/48IwlHvMtBrt154djsqlTHpGkHOMq
0kgbD0lyWc/tZ2yrfB2mxIZv2qqDWauBpMCsJpVO609stEKb2ljejL5c3zxyS1tF
ukUTn6dbD26s3Ux7KVa0IL+yAvC4dnSE0Oa7zY1SWrSKx8jfPlMwNsaFnHAAAcBE
8yN2jp0lce15v46nICIKsdGg9isirCp3DsNjdLT8Ta8GDIgWNFNYdnsEC/VrwtqM
qeZP08+lDwtMArMK5iy8o/Nsx+VF7Ia53QZFvozIu4ep2f96F2hOBFjmV0csvLmr
PlRnZ2C89i64XEOWpw4jY+WXDmkF9qm2DvS59qCCDIvtWuube1clvsv6KQRj+os9
ZZNnrbwRnQ4O+Cm8l2gNBhp9iyN2VO01srkcGc3m87aKNQmdqGvtmOnmRhPh7Avz
0B5Vd7e4eJQOl1Uz1zq/cN2glmvIBFCrtNEwuxieibDujbiW6O8LqeN3d5VYK7cn
b9JRCB5ej2tzdRYDh/Mm4iND+eZk4pwq6gR5VeyVb/tcZK6QGJqB6HShlTYmO2bq
BugoBs+9ATVMUd69UqXvPuR4Bu+oVqJNX9vYr+nH+5uWuUsaQoF3Xv/n0rWhBhSc
v7JinvPR2FVnYN9hJisKMbP1yBDYcfpb2nBwHusn6NJF+8on/gkBdbZnJKsZfYlq
Zpw6jKTIVZfdP+SRoej7Seucge0AKdWkdnXJKWPyAxMlGJcEYRqgRLxE7D+2ez6i
VKOgZvdqd41efBlQVLje+PGzYk7Gk84Drx4vSFES5absQVI0fYjddLH6yPlKrGjs
`protect END_PROTECTED
