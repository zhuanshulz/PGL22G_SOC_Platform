`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PxZQ5yDHUpbH5ukQ03duieyEepbTYOncdS386Lw1kW4DDzrvhZd/41ghYO5eiopZ
NEgT4MWKr0QfUJr0+u4/YUjrC0Wgu9p1PXCetDj72J27Wz8MMW1liPRVkANsUmkX
5zkNs+DY2bwJpm7cDAnkxpwtbm7I4B0C31eJqlBVNPRToXMCokbmYutjpP04BqEl
vmNoOfzGs9J+HY7ycwIqKZKekteb1Z6TjnI4nh5ahkBz1z5HvqUsS3dS03EzI3OT
0Ilh+xHN6BNGRsPZPZ0WlRTmIY/j9Yeae+SyIdei2g1fT+15p+f8xYWr+8cSOwe+
rwwYcI6ApZu48I6gvvUxMYRxyNVfHM2/LL/HcAwnZczUyUHH7o+iraEBiAk6tp3Z
Y//fmUZsc7jNBUCHp/HFMk89jR/BiA1ukBnmVCCodO2gxz34tCeXYstJeEy99f8q
ih/PSLfW/s6UT7an1IRQJTTMZo3PvsDrfEZSyT/hAe5DSW1cG2Dj9pZuIGBR93/7
mFSsmERaXrhvgHaD0Ig64gbahsU4OIAsIj0Ika1flXpzvDCKLts1PdOSDrZnI1V/
WU6BVz6tqOCot4bmxknrQbmjtqjM0jDOAtmjYQ7qA0gYH6mrLQnTnILHmTPnBdk3
U85Iyse118+NjVb/+Z6V6ITYsCwj8gt/ZscHgAJFH4A221BmIOAyHKIpWcIjQQGy
KHAQSV9T3VIGuMOwV9NSmNyn9+aHJFw5xsdTFz30wsYuJEClBicQ43/LBZnbyYMI
CuCs+oK44xlA/QtPc8rTegndlP0yt/AHaQJTZNKFVWfLixehXYHELobhbg5ZC48U
qrKacxfWoLEoL5BUDNUM6cex2PIW/TrRdl+YWT2AT5Cbds7RzPFyJgeC/SxW/BLv
Nshav7jlL0jW1SgKJ3Z+vj44h8tl9o2vxiv8+9aD1qDiWDmrSPqYmE0zjezpZktK
JEiWk9PM4kAjd2UKz6jZEVFGAiWBvXqrYC0gRPaClnHuYfdyD0RRkr6MiPxHudrx
uvVKTg8EXg4VTkXRYQ6TssGp1riiQABNg2lz/YS5oAfTwovwZ1wWSDiCZmv3dXs8
ACiKUALCwViMO4FJ+bNQCCZANlgWEUPY6CUTX22lDMpLKXmSMQExXU+VMSh5HtG+
KeFSpthyAvjLiDKIyZIhrmiAxgChtEnewTmoTHfudA2QvzVhjGYERC0vFlvi9D+3
xK1l/g9tLdculWSGIofR+AGUmMrJ1wZ0/gT7sVFdpTyjdS8Z/xKH3Q1W60zcCmMJ
2V/e7DdZccyXvJivn1MKDvqICEBBV6E1TB23f43zKYheJS04JvDJrvWRfUSiEAcf
cfT2G2qsAOCFPBeVO5QuyB3X7tK58NSHi4FH1ZnO302KxkYWdIkWMDDnfQyhyQ8Q
Xesq9YNR+KxSBv5VCaNWZyAAW7bmqHt6RK/elDZJ7g4hXSMTlZjPjZAfxQyGp2LE
KlpzPuR1ZJG5XkJ6lY05E53tkWwAE83j74itVQlF+tJq2b3L93fhb7fwVEMiWiNU
ZrWvO1zQkxSHgfKE25STViGLtz0//4jNYHp8TnYXhFOkJ9Sr6aXkITNc5y/E89go
hen2wfwi951+FnBBULFjQWZiheQIxYdeQCT53SaRdbemQK8mRPwl5PD0AHwQkv/X
feg3eO0SgWbAmJRdnHqUzVJkB8DodpVcP9wqS04wQqrvtZSMF//RRNR3lPyQ1Cdd
4YNlpGB6Y7wbySaTErOrX5jXmSgl67+PAyEheYGobJQKon9XfGGRSbC/+VknB2qw
Bkzu1OD7hoiyWT5J7FTyzHrWOCErCOFbP2v4G3ZvyJ3HpdFj5BMowBXy3KMITcq8
LnXR5VcVMDuYBpq8rI45iy75yZxNEKgV/a+d366Ol1bTcGa3CYf59Ihbgi/9hlBx
gQTi2SSQxELNGpFL4x8MHlqiLTG8lZINC9p2ydjqwePW5HtEFUXuSlM9RL4VOccb
kRwJi/kLzLxB2JOQAj0oaae+E8u//NZHBLLZ/nPUfZiCNZJ9jjIpmzDcPCY4rk7T
19Bk/9ieMBfmiX+eolY0IalSrrPHgGRhurwPO/dvlUgWBtyZF+yVG+M8ykDTbrt3
Bu8/fiz7sowiUNNyzDWLl7tJlmsLyr+szLTmLxyujyV2Rf0O9BYNAwH55018+xSF
jioZClafoeJC2dc2CGIxp86pZU49KAQML9sFG95Dj8bP8KoE/LkftcGrHsmC5u7t
PbbxuEmrOi+1vP+rEYccqeEtQV0WorgN//lc/8QN6f+eumCU4TBe1FnSyXCyIIqJ
x6z3aIrsYdYeBJy8r64Un1uT6XDFIuB/GkjhVQy0gT02pPrOBOyemMbUnFJKb52y
YVmFRtxnWYc0cyH7BH0Yag==
`protect END_PROTECTED
