`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cpfgH9SoxuEK22HwEj4vWh+toqloeXFdeulILm12c/9pdsGQGFhKOxCvLeOuCH7l
ZhazBU00H+3rbmK0oARakusYgsanDmLzT8O8Dnw0j1pujL7rjPwygU0qOBTmscqy
F4FMw1LvGDa69aht+Rsxyj4vrwzWsI1eRwe5Yzzpb0KdfXwW3ig+CgRU9Q/YXfbt
AUXPmxmsKalLaSmzjBvzFFAg53ccLCjR3/oDIu/64JMsO82gOk5aGNSJsBm+vkjh
fWKAgRkp+ygocqGWHTDbYo8x6HWtCXTqaGjJ1s5DwL4kQwx5Tw6I2pcdnipoHbqt
ntO2i2o/o6QW89NhNhQWsXJiYBgfOKV64khKlka7NGxTeX+OiofCMO2MY0TG6Ari
vwIwqIO6DjjtbfubGvfvddTDCax/qgrVeSj7BSnNv2zWWm80AAzgIa8JmqLbQgXm
VlZzwxSCu1lflMjKYD0H3DsKVY2QedacSskVpcSnLRuP5gq2YyBaU+wM927fVhxw
U36B/oUyr9PMEx95+4pSnl52kPUU6J+06Gmdbyy12UraIw6WmQ+ASZ1r1TFq25j9
iqMda3dBmbL/G4+pU2ArM+j9GADBc3wZys/lgDWk2ut3OoxY3edtf1+7AqGd6b8G
JJLWtqG6EraYMwsqqHCgB9t4MuN5a2CPbPxbtG4dFJ31eS627fmZ70cleyTgeXl+
tcZaswCckDDO+ewQ9xGUYZNjHmMRmb2Sa0Yaebo/jwCfbsfOjhKPWHUZeJS78aS9
qbbI9ljmQqnCSp2895Y57wvjPeILcEpQKXXwuTqGqNBvDSgVcBMkqlt+wLfJBdw3
udnwaF4xaGX+qXH69/9kP9oLLs8GaZ9GI2UR34A1yf2k1OG/UsqcaADgayvkRu93
k4cdABzIPBysUZvxJ06ZxFW6myYoYKiX0OHynVQMl2zXeOaKPJbgoFZJ7NBMAgzG
+Q/aRrce2mlBiJ2ofpNF7Z7Il1VrtdfXKCzhBsJvHSY7lem9pILgsb1PQrQovCQA
AqGBAQfgXBU/03rMVbgiIHP/1xKU6RaPVmtiGLCFwZszkW0eD+wFs4vPq4jHpFeQ
9RmHDcy4eMtNMRenBB10pO7VHBmHMfW+RMXw+dTZ7GBeT6PVTHz+XJV7L3bxyZYj
3/5vR7dta3YDQYD7rGLlUr/myxiaA+HKweDPc5VH6SNch0lhYT211WfJ8cDu1c7m
LcwqZ4s5s1t26rqK85eI26nJSz0Euw4axf46LvPu0xwO+qrt2RzVfec60lx5xA6C
/WHA2g5gRrJoVdh54Jaw+K7eE0VFOQpzSF93uQ/7zAeucOe3e7XbSnA9sjSLySc9
zuqUQreKP5NmAl10Wui9D3uaK+Q53FCXCpAYnpvMkGL+2V481ttZgKU1AP/5b7Uw
unScoFN3mvu/Q831lM9qBm684XdPwE7J9lzVoScr+My98q0qbrpCabAdfO/yeZ1G
Qy7pE8vbUb6DqoExgDGw8562bwrdds5s9G0VF2FRPQDuXoXIIxy9QPUBS3hbpH/J
pObGC8QQNImIHEBDbVcOX+iVKcF6+OgvawnY5P7smyjo28Oh5ue6CgFajqbfwu80
N+EB4pB9Qq0mB9ktHIU97A1xNwjQ8Y/opXcfwDC9XFZzOLt3aqcsQU3ioUjMisNs
SuigumdkPqfjh9UCMO7J8CJexQ4L4dfKZWFpL+QPCEhXOi8pQSdtNA7uJ0XqN7iY
kfvi+f8c83l0UOETJ2UhATyE925U8F3jBhv2zBAcGCpmkgeSoQzJtMiRTgcLp6mm
URcWXhnK6W88leCEIbSj3EfyvFZIKNzDfH2/iqia3W8dboYe9Y+Y1a2X3gim8/TV
M5CpsJ1upAmLrGrjt9gFMeLQgbU9fxQV6xt+PcTzY9Gsk3jieIgAMuP/Rxy9H0xo
7Glw6w/AL1GoGRDs8orZ1mvHr0qig0tMZ6LH/yi0hGpqHTHLWLkx6T0XzVUyZqc2
+5qgnp4jtajxC7zVX1E/S/t/mjEocqt2BJUoYgQhhuoRtCGhTk/w33SmFZqUteg4
AqA8IQxOUXnt65jGp8KNI+03+WqtTk1pvcgSEyu2qr6zB/zSC+6tpWx2gxkIrwd2
LXKQQFzGCMWgB5DyTcFgqUR6z8p+V1eSn8Vpx4gHOu9KpTVLPAXjt/Ajq0Ji69z2
BlasKVmXbO1fsV90PLa5QZ3+9HmOLK19iuZiXFuZv74fcM/CD3LaShRrbzJKc7iq
5CpANyh5/pFXof40VRXfWyT2WrXTvM1+meSGN0elKF3/t+kojPBy/sNkuDRUcDwn
QWhak8wcPUG3uNW0HmnQy35qCyacVHzTJVYkadlu4gyryxWImUBjTMMdcC/1YFOR
OGQe35rCrk1vokvHRftnkEqWQWZ2nT/pH82GKmpwZaSTn2hxDFF41S55PYsH33d+
LHEIfekiJ+4bNjD31ahv8FB6frn1Udaz7cWh7UI7Ueua3Df7kCCNYDMQF60RV69p
/i/hPBI+0esdn+/bgXrfD56FAfWgZv/XYuxOiCIfj9jSik4l/P83ScFcSppExUly
QWTlF72EqwqRJ/vh8kNhye18pfBDmgRyzqbXdRtifuJhONhLaWUbrKgQQZLix2cx
zNGF976CzO0/66cdgmr/hoqm+G0DAUL6U362rOW7N0mKE4nYuBTkr2SvAurfXbBw
CJGjtx8Ea2qzSehfDOLKlgrHldhtSeDD7KKD9erHFoTH0vgnA7jZ1Ad0GzwaTZOZ
3CSCruE+3PR4fwotA1BqmgrS6b4hvKPi89ILLP/byZcMDkJfhJ3it7MfdRKGf3im
swZgHGc1jqtysEqVSSjWKVLUgndCvJKp/1FTCIbyLwMr/RbXM6kc1HJi/ft/A/KU
WxQb70GlVyZUtOptv8sOwtA5Fw/VCg/Prr3F0dnD4nPu7L8LfeqHxMvho4cbhfpu
bHIJZBHZxxwLCfBxre0nO3bIG7yoXBJLONU6KPgiRUqBWhjatqyaipeHrTnyKrKA
ITpT2fFLMYRUVVurAzrfY6BwcQTx+jUdY3Aiyi5st+glIhkmV/BrL600SBdXvzZA
SfgURYZ99kexKv310shVqrIJLzCijNggllIHb0DJ/iXoc8mYfITbiQbfBsXWZAHK
vfmuqQzU4dHcJpz0gMouTzRlG9ntvXok7GzwxYjXlK8GpISAUdsGbxxNcd5BhK6d
zP6eaN0avuBZ9UYcrjeiQZGYieHJcvuYoEQUGWCoELalIi5yb8SErgTJAsnGAB/T
pgYCKhJNea+ht1cCO/NDrla51m37V/Pg28nD0PXJd3XxVxkV0XDRfN/+HqRO9lvK
cXgmCcA2LSEpoMAD/q713BFJISwjtCZCOy29K07RVvd5eiHA1xvAvCV6ZEEE53tM
ZAj9kf3Ga93mQJhZiZtRdv99gVKW/HEb6/zFHIFiYG0r87TA3zk1JuKyaYfPfWVg
7bhGwl2QgVa/71G1waPGIIJWcD8IIWVjG6A1fS+CXM4hQUAmeL05ZBiXJOJAU2rn
KxvRAmbv0DCZ5bYe9vPoxvFVX2ScbbBrrnqtgtWur87jslxkpXwTB9TAuhWpN2vV
ZU9uCtNb1qdoKWs2/+IuVabGkef0gkU5/KR2fYQW38p4I6jJCo6tG2bsLpuANH7j
cCb/HZuYlLdvQvBqfw6vSmkc2ci+yLqziGOGuuk4qQ5uip1+uu7uD2dBpDF5IUwf
G+k/Le/U+yDM+Fl48GMEDiPDcPkWAqUe3N9sgp6E8OvLgdAnXtH1Pn+2oG3W7w1x
+faO+AKYJpriybYfBnbMS1/yoTYi5O3g/WewKnwSccxb+vNgH4htGgB9Ry68IFT1
/VduYwE4bVEYJj2b4shY7oUrMsUxyh4MOePZcTZyVictFHeb4hepp3Kw9Fb35KOi
j2yDyrthCTz/gOvCvMz7p8PCN0M8mjlOMnq9qVzAS2FD1qRLKjya9RaFzxj2KDzr
B/GEXTfJxfKCPVbuTFxtfHYDTv/1GGSmfbYmZrs7lU1OldIVRE8rQhuYwINdw/rg
o2WMQ7zKMNjju6+nXYPYdfg7jWFA9jVOTFrp4j8HCbYzsX51t7s48xN05yi8mSQe
D7Ktmzd/7RBPZuGVlLwSSPCtRsrlWNCCJR3f1t6BKXtHu3LdQBWPD8OkPIeBTBQT
fhEbBaUj3upM4Y7p/y5m4hBbBeJRhQu03LN7OIX69vw0HXbbcI5NxAp/fuw7nQdm
LLAJXlX5U+WQk80Lt88oenCaKQFZ33GYRoq+QEX+VcVkuQkmv69V2XFSqj2j/C9L
e/yUqUTl2885XGicTcIkSr7uyzECtDVt7iTs3VBbh97zTkoWuqc/DaZMvHnu3A7h
FHVRyX5qXZfQDpMLEI1/PKT/ViUp0eIGsFWPcMYyhd3pccN86LxZ1RMWMLFNkEPu
ZmJSB4WHPPffdhe8CBss7pNC8XcLEtnhbxTmhTwhZWShh5QhOWOKR5QuiQ4SjF1y
+ahYdA1WqX8/u/HD8XB5AgJKhJTN8F56/zraDwEkjP2u2YgpA7d7RSvsnf4fe9g4
a5s0MQAmMIQ4YVcrnZ83FpJuQae7nQL8nGagqFX/uElKl/wlv7Q3pK2vumJG+1L6
oqyJIPdzYADa0dDVncADXz/wLO9wPQH2X+8/BLE2Rz0YurwMiMpEPkiNABikrAiO
bMhndv4R84s2bXixE5If4MwsnPeLkanmMgy2caafQIipnb2RDRc4+P333LhKiuOh
ieepZU7pihGCP0R+JmgLyrvs7hW3BWMg31whBspyk6UNvpSWtWz4t2AqqWBLP4tt
WjIqNJ2JGZK9tFHMJDt7aGRC3y+0Eech2A6piTIGAQCHzYISm9Ttl6VwnLh2PjKG
EgSalBDLV5QOcfuUlhgThvPYyHW6DwImovqqLen6rP4Ebq1/dVO9/NdIyn7r9YTm
RLN7lKagQy5LWHRCuvhF1Rayfe2EzRKP7QsRn1Q0lslZu9qDnsPis9z8souR3aS3
hr1dcx0EtwyG2n3ub9lGzk6UuY5JjQCC0ZD5M/T+e0kb2bv4jBhU0/OM1CeCwK8P
FY/SxP8ZjmV9Lr6Hs7BVCzj+gjnIFT5x9XwuSvhh5iOTvuO2NMvv0ALm4E68tknC
d1MGYZmW6rh5b3OzEn1W5xXUb1+sP+/CVC9lyI/H2J1Hd43Fpbidk/3huP7ut604
HXI8+li74+QmYFyIAFAAUEiz8RkevOYiGhfmCGBAmzGlKtQP8hrqdi6R/dVP2h+u
H9TB0ku8EOiN2DGWoFE0Iy6dS4LrARuqh1Vb0KMw44tu9EMMZOns56SwIeCgyBbl
JNhj66Hrxrdz1TU5H4mhGc409z8w7jgL2vB/ft+UUQlaTJJRCPgQcWg+/rUuVVnH
T7mc6vkL74q9U6mv07XowNr0V1zpUzh9yfk0CutfDTOcdrgS3+5Bzs2Iol2qSDk5
3DVfGHekBRkhMah4YflpiFsre+GniDvaah9+n1MEN2mvPJo8KrRQTfPpMulif47A
32oNQfPW8Y04+MDWtfa3+9DlBEZB7hkvHlpvXynNBEG9YkFmGxr+/baS0oPGf9BB
XgGvuOBOOa8oGVpkZbddVPhEJWjwh1gokQsNpu6hmh7FOp4Ch15NGyZVALqm71v9
YD6CXv+Hiwd7z0Vqf13dYYSDzevSE0CM94biEwX+VFfJHYS5XwvNf3p+vGXbwxD1
+RGfSwC5BE/oqUlbWht0dZZxqQEtkQaFZoFb1oB0d0PPZZLJrYRVQPXWtqVLIXhs
iBPsTA8Ed8a5APFN7whkfrYHFc9oZTUbkA8/+0FJE2tHABszDW5Ym2gFakig8KHB
byfK2PITl9VHF+s6M0wHhhEEzxZRJ3Sb5KeZP7FYczyRZ5B2WPkklmo6zJr+dMbo
GqqFT2vvHyueE89EskL7pp9QHP0erISy3Pi3HgKJT3lksVRuqzusCcgjBzE570Mw
xEawa961eD88zJ7L0KFAEMGIiWg0+XDIh2qU2nVOo5lixklu+yf8p3fesWLVmfB/
rgQ5W6dWjgl3OAvQMNwXpfCjsbRj2DGk968hb6stySuqW7gUbm7Iz1wiriv8GQkN
GJzFce2UcEpwgiYV5CHPz9tG87vG1dUmTnSfa4s7Jw0m+T30OjW7R4djLO/Z2J0N
Pi+1JPsriN2naN/8sa9iORGJ4HBhetfCTycWeL4teciznufQuQhPeh5Gs2VWLgKk
hvA9cbOR0I5iQUUlIcGmGHbeLvUDACScEJj06joS/TLGu6NNLWcuzlLGgFPrAd0p
mY8V8fgQI3WVgsYT8odIPYOnuD15QPQS+Q4TVnFowM3/JLQqftxva3QxBeJKK+JB
IwCIT1CbdZguC8lByfSjGMbLGhD/0K9SK3ITcXGsSb9Faf9osqYatEihIlL8RK4F
6aJTmttrhsjgR+zpW3BprQBtI3PvRfeoIw+Mowjy6Vdentj/U0u+ZcnGfoJBUy9m
jQthcDURNthemWMJ9yk8oawJcEczNjB5sgexJWQYFYsjYQuvcpzhi4rBI1q9mqGi
DOSG/K4tLTIenIAINaLkx75VQsSMX//v3RI1i7Rh1+jNkes76PxDXNyQxFN8bkH1
P1g8DzL+dJbQ72FCijk/rjhCsMo/Gn9Dm0bh/VW0gX3sCRMGcVBHEABChoLUEpRr
BY6mtyw67xmAWZX38JDBdTXGIbFAQKOUtYAYNK8FKzka63nY66KIIiPgbC3vf8Uk
mwb7Pz+9mIEos5wJEv90ppM4zhXXHd0LLyFi0ZzIgBeSg/ZLP7Dzg02WsT2RCt7P
EFYuGzjpnwzvxsiXNThWME8sCPagqs4UkxgqVX0cwOyHBIA6OfNEDzvYid6V+ROR
HX8pTSa0BbQrYzFxu0tH943cNMANCp9UTKDjkiSj5HS63MBw/vsujgQ0KsX7BI9l
mEmOrmOcXqBEH9TDyNYHwg==
`protect END_PROTECTED
