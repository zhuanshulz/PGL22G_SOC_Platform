`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HGVti38ByrbsjLH8iBJRM1AJC13sFC73LJxwegv0zQDOmrw3psooNWdHMKy3KotW
SvLzztkhPSzmtdlKt4DUP/X8QVrufFSEfcthusjcm6xSIZRXSORPrvVHx/zPSMzk
euDI1FS8IE8sT42K1sfh0LiQ6IHzxO3LYph3yWHWMMNm4bKvG4WIcfxuw9SnGKqs
sfeP9gDbRyGY2pVVb0wsUCj4M+xsGYXYxBDAoCw5qgMoAmpb/6DiAZQUYiW11jn7
1iXvN9FjKlfxzq6fXGgM1MZqu59GWNX6xAWBVVG2omTs97DhFlKH/pSnDmhFYF05
TXz1lVitG+hKXVoWVPdkzTJ0HUgPaWIH/VQ/uoN0vQlVEHaPPP59l1S7Z6MDGp8s
F8WgqQkqpIXlydWeq2fLmLXeNY4tMg032KzsvNFID60P2iFcmDgr9o+E6qJlsji5
xMpBHsNsM5+cCcepH/CuvZQr5nNiRQ3+YXLRLF9kekSA85ZAVnFSpVdeaZwQk4+f
91mgQ70YCOGBcP4MIAnIm+N7SAJQQQJ6JHHw9zKWmLgpYLiyaDSm90GHkRc3xulI
7/ZlMcN4XDuN/WJAJcUDKaYqrXPQ9Wp5GSWXaQGYHOPyEcsbArHV31QfrnO9jFBz
Fg0+OGKxxxIwe7a2M4mSJj6fuv1MIH+TCngbfqSGzte8nTI//cQGobA90yPoleOi
Go0wyfHurcoU06jAZzvoGx+yLIgZHSR8tFyEevJ6QnkIYy/pCHhHs5IYG9feUyoP
97j1GoQWHqR8bHBYefmAdyl/pVpT6SkjbJjDr97UEUL6emdBBiLO+HuKTzWGjrAW
tNooXrBVXqi/ERbvXAE5nHmdHsFkvFtfzAWtXGiE8sg1ME9ltfDabmFM/KltG+em
zPOEsHssd+yhfM5wQ7zfEdfqaE9J46FcY0QDkIgTldK0aUp2/EWfOBw5cZFrt5Zq
enp2SeR4oM2UI4zxL7/aWjOawtZs+l2XcooISmSwR2DuwHCzBYxc/ZpW0mjVWWW7
QQKvf+pO3salBhRGtAljCHyX0zcSx5OP8Prd05NY9acL+lqSV1s3l/JAI1CM99sd
lSW7bcT5KRo6hzLC0r1j7OzbDh4F9oQwjAT0UTZBvq/Vc+Ll2tVCpYBfVNDKeDR+
H6JgJgKL/vu3a0T9IUFF5jx8MyfoTNxf7NNN7E/ciyLiW5wgXWvRxIsZjUxYFFoN
NcBKlr9X5zEWJTemKKWHdkVSLroDkkfUHdkojeG+dLRf4HorgsYNjrLm6AZL+GqE
M5QUKw5N+2Bqj57vKbMWgjc2/wJ6OJJ28ik5GwPu9tzxTX64JLCW9r9somjShBBC
xWZ+EhAFWtfTG/V9f4b5Fl26O50hE76ru4RAbxdN6FMuzu5UHbEjfZTT3kyWyEDq
NmoUcqThNBtcVtpdTXAoMvOhz9IJj+xE7Grhvb5L4NBQC0f6CZT8TkU0SYPqTS93
eTgT6wglye1Nf+LYjaGnjPze+kRKa/d/GASD8APcSRHHCYY/6Nablgot9nwvelQh
zNPL2TyXkJPd6Qkr4W4hhPsTmiWUWbldIEuZNqypojWYbaWJimM3REQDHih5U0ys
Pa5kCkkTaIC4v7O9tDVZoB24NAOJpDIN45C+7j1bi718lIDwQ3O+dTQzpT/Oxwuk
hitY+p0Ku+2cIrXqU6ku+MFzamFxlC4a3p2PjwdTFrMfKpGhmxTI+oLRoNDvOIu1
B3VK00Uy68qinDAWeTDbppibEIsZjDoGMSm8DnC8snHxH2otK2bT2Q0kwqRfg9Z0
1iD7g1H70CUX/RkkVEm+m1D79/VxpVyurL9OEeBSElPEYVhsDcRUHK/jFYNSoSm1
Eflgot1aTfkL/IjDr0hM+VZSq+9MDDjChUHySHi3odUe6sixSwvivAmJBy3orrYt
KMCmBK/LaUpKpKgghEIt4jTTQzIR9ECzdvDiD+Rs5d0RGg8i2+RRu4N7hxLJgM93
Vd2c4ZG0H5CLG6Iqg1MNsyvn6bwyu9R6FNNQM5Rl8AdsELSJ0PedmNL+k8UObWvH
ymLVIsVgsbbpkbjfE5n680liUseklk6plcpbY6BNbqy6+XYasAuoOIDvKZzgQhxX
pK/qZjGdh8YaXvWgau8CBcM6uAQECfMD4GgPNB1P0KX+XyMSOi3T+aDfFhxtSfKg
a3Yggk/xSHAzDrK6V5U8CrxOCv3sq6YBHbADDZ6S5PV+tvPuDn9Vs0PsR4igZ5Cj
BU/k2zF1k/pCzk47qyp4zvsAXDlNa0mUuZDZrTE7AXQtexH9LRFeUa9XAu4pgn6t
2SFWad8Sd+p0QGGu+RjVOisd4I9DRrS86oRisss+xiXPe4zIEbTgKUUFnU27ScLg
U7bNJjBIPuHz+aMpQadth1jUYhXRS8DgS4c8jBpnK5MFUnIaNkrZUByUTCGJsZvn
/VCXdIecl8pPAJuB3GSNVBNp91AfzxA1+m3ncEWMSiDWQEf2Z9/GWs4jnbm4+R5V
U/d1BhMZUKmy6Di24s/NIJTvb3voWQ99ERFAxJ3GZO2ZWZQ38b51qE6ypKYX+yrh
zxRB5kE4Sa2Mm245KYYq3B8dljgoFyyosjWv8qxGC3Ue9aZd4OoL1ttbqvoy4iMm
N5sgrvKIduljsBtmAG6ALUcMXhUu1VKOU9mb8LWkWygM1BsST1XD0GjF6ZAeh5ZM
i6RPT+KLdZ4mZ+KmgDQehfcHkOZRy6D03ZG37Fo+LAJlw68tlPqL/6KLLrLHCqFt
0Mm74+ATmwGXRxHatmX7qw33cH9rMGAtfT/cdntFhpNPUX96688chcNTWEuR0iKw
mP5mApLizbSJp/xC/z1VGPq4BFWd0RZ6ce2ZVwNL0SaW4sAZ1hGJmSHqY6mabpRb
XBOaEgD/Lku8ibfXPErz2XJdQXhQ2cwlIGfGlpkb9RNNYi1brbpaBsDtanC+cG8h
qdnSRq60lwLAcPWeOHvvis/99veNZiY+hwptwcBaj3kxBVpjv9XMHbkOkolbvdvL
kbOXYc/4u86xo0a1qJNbb8pCP82HPLs6nBGM2t+Xg8CVT6QGLtMuKN8s1M4EoF8d
g/Ri2q8j6sl180U7lCprmYqupdZvJPv9NUBdWh1/GIHsO3qvrlNheu46lGwbnLPU
nMGTsrZ+46JJumxcd7/pDCcrw/eqy/6ozlMus+bTE+UYh/hgaknWSajXCHDFNumv
w0TX2QhcDYy9DbLn+hi0oGPC+DFLvVbzKf2HCxOar58UoHR0XT0HHhw6R5rqZAKs
FAnRHFMkIuA3JAcpojmmL7/4JIkcEBiaPXumdQRnORuV2FeAa8ZWAaraRv3KDAOE
RTruvsa2TJpjpD95vGn2mPdXTTdvXCwGSJH1v/SrqGVXlF8aCTOgbUhVTfAqi950
B8RqvtDUAEigZizOpFRjSOpV2TlXSvO7AkLX9bo1PCI7aMm/JnR1eOGVl4jUE6lY
+rhVqZl+JFcmI8aSRIzOqGfnmajpGbW+LGGzveeoO+XxBSz9GPSlB+RlRv3l9KPq
Swi3ncVL4w3FxWXM1GvNysI/VpOhNaV3YCJwVXkUYBs20xWjeBddHvuWNdXPhAll
TyiLXT1/dFSSbqoc6PyUuuhlVYGDcV9qEEW/pXWBkh9UtRJrsEzOBxFtebyH0+1+
OlIcLyNCeOHR5F3jvExoAj0Z+TPq59XHaXu25PHU9omf+iRyGDYMdO/pmPf0jgYd
pXLe3MwyKlrHNJQGs/NlDTesLQAUSr5hPNSOUIaKXqEdwI4ydQhkfZ4ZbniOYYoT
O7knatAJzs3N2rrbk0OMXzysZdkBW8YBGheyLDQlWhxxRvKUNTT6GMTyjY2QlRHR
kv05LERXsBMfAO6I6P763sW0qCkjx9zi3TYtvpELwAES9RqPt+HLwZ1ySTOOHAaL
vNriwSrB6oyRVVwkYqPYZTQg5YDOS7Z47MUeapSojmZGdTbbr40wjvK/lFjuGH9i
G9oEdtKiYUTvAxCfPNxOyLByNJymptEIIa4m1tLl5pE/Mp03YrOmGrAVBe1MG8l0
nw0E2+trWP3dt3MqUk0Kia70KXjD4wWesOpfkCMBs5XuVcvergoYriXPb0df0YU9
tLdnTa0mnyC8UQkPbTI1HY7ykFQEYa5/euFgNb1KiWWWvWrBfB5iyMeT7T0pItgv
hoCuQCKD89Uq1fLZvyrqdAdsEodVDtKJ6KGmN9VhpjxFBca9eHe8o2b8wWqH78v8
xkJ8FmDFUB6jXDPRgK15QKqp0OGbZ1BrtLdbahAnUsvwpz3O9LkH4qHtwmtTaQL0
qNsXF+ywXidO7nwFyrlxw9UP+mbMz0E0pRWzRRSAK8vA2whlgXoOt23H3IFzr2yo
uTX1nE33OjomZpcdOzifHmjJqmWixGupLY3yAh3LxtTIqsTfcjP9fHu8mVsLKSO4
pOA5fhZIJW/vJvudKeuWWZQwl4QKRipkFqPMlBnfxtj26yKcuUyJZzFiL/3AhDlQ
Qyid5E3uIYmU7VrOjqBJz5lAOprVK060hNH50qtAa72WHYwABoNsuOmONCGxpFSJ
YH68KrHGjnqSTf63+sx7IuzPMXDGjXt6ZW7B3iD/Z3TPpOZtElzPKQ3ZWAiiTPA1
16VSvprir3DeLZQGAu6CGqeFCE+KuiiJTkY3khPDusUDxX50lnFn4RVv5P5dz/oh
hrm6MlTwV68xBcUrnd5Epfa9PHhdSoMp/kZzluzNYd0gDJiEdLAvST9dIG/ahfY7
PAkSSiWMK4AHMFrAFbEeaLrOneYZItawPSYcLm+eNLPjygSXK497nqN3Co34EKpc
mRTGW44odQv3H0VeL8GWUqsiOCdQOXFqWv9+dQin56O93e6Yq+lkDPSfZFP45D7E
cS54PHTxOdgIek+BixTVztdi/VWL/kcrAbJa8fJeN9uvdgv2K+dizOjkBE7BHbvz
aujYrMdCxxUPqMXqLp2lL9eyzez6oJAFLm7uImHNTt9Xyh/WxJ371ywDWqiGOKYc
PWIYm0mM5P62DN7hcLA1M7pyO8CIRv11IiDjPVcrhNlD1qzz5l8BtX+HKZ/e+E0y
Dsr7eDGvfmHHHFibsy4eiDzhPSa0GyNudBrE+yASsGK7wI1gNGcgQn0VZgk2/jub
ia46UjNV8ktVyU5ZiJC1ntEpPbVvl0eljOJocCxNe2H87066fGY+m5MaVnmIzPrz
MrvKSQnbtK9xIQr1JPkNLEqQz8fYAZt1XT7XPmdf4WQtxxpc4cIkBn3DlAYEp//r
SJ4My3Dh7SSMmbR84xdncupPXo9jIwuHlVLwWcmSTToSbYkr7tFIf/es+16yoSAQ
qZDzMi1rNb05rCyqnhTS8g==
`protect END_PROTECTED
