`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
55fHMfDEirA6tGeN1x98NWoJpQwOje0RYPRdL69i/AaC824IHwcUL3Dym2MHAB6W
Hcy58+7GHRM8sQ9bsK0Y+atl9r4Rr+DFPxT5a5kqJhnHbC5mAriUW4hhfY2QjPW7
suZV75ulgu222Y5rrtRi/GZZLNnZjn1sMWjFIaGyaw3JD4Crora2jM21vKGpAF28
vrIhwaHYh8BZ4aRf9BBIKdqMkn84Vp4DJeZ55T8FSTIKJTZo1hneI+1x4PhcB0g+
4IlesXBc03Shr2ueaNdJrpj4WPEzsvFCmi+tTXG2XViuBpEBXx1CMqNZHvMnWb+z
F1UrKRUJUdbNO6bOjqaaj8JTKmPODitEPT+j/DHo1oC+2+m8cs2O0KHES2LjQj4i
fC9yBrE3JyKZoClGo4FkFkN2HqRpqY1yex69y/Pq2HY2ltIJg6jgXs7tXi4kSv04
DWNjbnJjUhX71Svp70GLW91zu5sfMLguD6CLGsCcXlpQzfPrqWMvqz9dt6Nj15Ls
WwpbI9iLC4jtBTa9xvsbIfTJPBbtKRBRxyxTZ45F0crLcQ+9gQvwLMUjdYiiWfLx
doIBdJieoxZ7PjgZQMJVZ51JZ/MeRAMEh7i3+4JsKY1VwINPtze5iTWrE9XwtSyp
Z7ZXJQ1+JjCTGAZLH3ulniYNSybYhE6WQFJB8uAOXWxh6uVXRP0kSBS6DGewoS2l
YIlWEM34BjcmrZj2gjdM5c8HQcb1/R2R4mEzcuQN2zdOFSr3+MuIZv42V7AxSGIp
efUC/Y26MwF/LmVCdCpGq6AUKDf8GJEUflkmnrPBAVmA3RmSg7RZrQ5Mef+uQnTQ
QU8nhwePU/0zHllT2mrXLqzR+pC2kJSP9R9DGwHCa3Q9YQTg2TTqaQR5a1uP7qq7
cD7CjHMcYasQPcqk7V2MfLwJYxs4sQcJP2GhZm3nqjA32WppX2s4CQHLm/DBFWK+
ykm/QYCpeSIt0Wmo+ODRnM/To13T2Cdr8jynFsMkFVqt51CeSTaCVrmTaWrAO5Pm
`protect END_PROTECTED
