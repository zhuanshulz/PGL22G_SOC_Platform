`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4SycShZNtdugF8Aa0QSe+Ej7Q1q3AHjMkf6d4kZMT/r+wvzMefPcGztfWHSPsnLx
jjWLD1nXgLlftk7MDB2XXtL5yIQyfpyuHPpkq418p6aUaH3NJM+ehDh2+1g0cAtU
ige5O54lMCyu+50Z2iLQLw/FvJUqj78DkP0unMMtJah52kKbdGqNUycguhZg4rvH
UCQ2EHLGtpx7/d1/rvRtTC2BwCpaGOKeIBnXwnh6kLSx0WiD/9m74ep1wsOWcgLQ
d45inPdfTE16QvTI62wF8r20bLIkflI8L8AmLzsimYy+WHMmAOmoJUFAT9d4MJ5f
lV9M4xvHY1DAWtMVrbMfGNgxvTkVIRrgwLU6R0bvstlUaPl78v54y73G8C7bIhdB
42zWjlgPSBAJ7doHyG6zK/7k81UmfDSfHlDekYNjrpiKojbjyYjj0qAytkkL16DJ
/m2oJAMGZ+dKQhMdmSkqX8s9CSC/cHNUH+Fx13zueF+zUwGNi48U5zlu2XDNtaPF
WMjbOsfGroh1IknIzCySvNkfKI4eMDPZnjgTX1kWmvB73KJRVVXIW3WZoy7K8VFj
+hOmfqqCi9Zf7JKqT2G/Qg==
`protect END_PROTECTED
