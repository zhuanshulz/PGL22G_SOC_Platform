`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5Cqmm1PP5uK46YS/ExRoT4CeLS40HbxrfJmPsUhzXz0YHZbcH9QWA9j1SySLBYYR
/q/xucuOJU9gBiJxvkM4AwNxPta0gFu/hBi4E7InuoU8GIVwVV/1DIJc8FmRehEi
sIKhZyGFLPC8qxgBIGip1WnaSIhRgg2HEwQ7VhnQeBcHYDQx4RRbxtVEaEDa0K+V
CNfhSC70i5gVkUOYwcQgWqGe/65krSWpNLFPLx+50pT3tx5YUIEqQre2tIeJn/R4
iXWHjtFZVXD9IkqI2XURJrjKC6l6SH2xqm1NgQ7XGgJI722qcgEyRwNyzGN2dBY6
KTdC8kmWGujwHRRU1xZljY0MRo4EDOgdVDCq04E9HAqxcESE0Mnp6ZkRPZi+RKmi
9D2y9nIvXMZft/8llOrWgoPv+LSb1D+63b7abKK+wRjHmD/way54pkHoeVG4eS/p
7C/ODpb7o4PXGN4tHFOPaTVPb5tP+JdkYjm1HuP9mbwp7BGF5gWSdzjlk689sgBY
NotY35Bzitlv5Ign2EU/p2JVn1KOjaPdG81BbN6ooTrA2Olx5VMllTdwNBvDH3uU
Pij6GdffK4XqD+rsIDgYBS/Qx85m0bGAle0oqdnZ/iu2fbOqN4GgsjrylNs1igvQ
Wb3eafmbvQV+gbXZS9wsmbTylmn3UwsQkCLf2Ni5CPuGTDgztmUaOeFkRs+ZYgvz
iDdFpTNg5gQiTur7NhGQ3pM+ktMQS6WFo557hOqMmYlyHCrjiJCUpagWBExv9/Ie
GL7jiMGUumxtevONcLB+Wu3r/0hT+4nZfX1hEoKPGXl99/mFwrWiwHWyhkKzkZvF
`protect END_PROTECTED
