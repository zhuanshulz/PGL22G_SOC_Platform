`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pu8fFqdg0pb5yI9qfWyMPMzVPMAywxDmhjVakF8hx9oZdEgG9vMMgbDfa8wNXzdq
Ew1Go2ySFXNEk24GOmGqnikt2wjeS4y9ZQ/0US16Ggyvs1tj/UNApMD2jQ2Y101R
FV9A0soHNVe26fOdsADUD9DdjWqXUuNxWL7rSaysCV2ENmqpUX1IerCMMaaCKjIr
ehAj1oi3sdcdi8ZkKD/5yhsySuGU822whxxkexn0FNCKCGxoqSbxq2rYstzgyMsK
W+ddsgxGBhqixcUum3OP3aBZFV1okoaSytWYiiFfhWewViAfA10B3WDOM6Io09xs
BqNbymH4qLSv/tfrJ0xFaHawVKUcGVHMpgwsNwCGWDnrZXJRSqAhy6WlTXnw085y
DZXKw8a1sxIcAR4SCVB8IW3b2cxNoxbBBHFTA6f/1rdSEARZB8tw6UXT/wopd7cX
aAoUvvvUXKeYynuIwwzS4K1+YS+xELl8F8jc8HY4KaVhKXx/pSfqWJgi3aNPgEpJ
TA3TyNNzCfhoNvwyv5lVe0Luow+OXthYBECO4PREizsB8uOsjoEYxRptqWI/fim7
tqm7hF/6SwZMbgNCEU6w9oJD9jkQtMrIMatP7M7ccIKnMkLwdi4/o5rB7QFUBBxA
EbsvhkRvNO47OPsd6+7e8D89MpZE3kp7zppuid2PqgHuvt6gt6LzPjeS2HZq+0sS
iAmVgRY84dWZM0psPYqmfk0JxMDmoT6HaGcPg+Bfr99+TmB3kF9kjcN1E0PyIWiB
pQqzTxKydT+NK0F62AH/fsfsiQc25osBwVaFWnL18vSTFVfwnoo5NhzQNmcRSReM
9poh+2APcSrC51DfPw7Um9UWADuskFnd29FmioxfaTrGXjfQhTXZiImUaklTLPIr
yuj4jd6vCfgz3pCLUxbngNDNy9lJmWbLZl9tC8CAhn/iqyAgajnmnpd1bf6yVgpd
brJqopOyJP5I8eehkDG4gZT1ck6W/uQ7I6tEB1DVLPaFyCqbCAQmPLJJWd73l5ej
OqKR0nv4WNrB9sNqLAuULl8QNWQ30xQuGpwPwaAxt2eDupoN9dLyy6BznGl6yav2
`protect END_PROTECTED
