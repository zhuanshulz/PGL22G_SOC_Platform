`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ol99FBAEiPNPM2qS9sbwLtWvvOO0O/VzFKxYOpxYaWsuZLd9i5+nRRti+8kUCMN6
PN51xX2vp6I1K3unaW7gXgW0uWv8mIToGxkxdaeJIRpIDWLo0pP5fZSGjJdBdQlG
F81MgZuIZNTlT4k4JtujYwTmICGFI6T0S/9IHQraWrsC//5Ie0vCqFFLIIrVQex2
qux8hieVEAANG9fMS5+fklLlBk+e/iAK1CQWWMATZ8jWi5vsfHPs6x1owXjlJV1w
BBZrEd4yWh/5fQkx7pULSysO/D3IZ7PdQswxTcaquWrk+leNUg1JKOp2ssCfmtLx
tsKDE2sOnG1aCDOmnyrNcgVFIPV/kyb0QrqNL0UkEtGRAuZV4nMNEUXMKOhZrK7F
tiYBqcJ8jJ2PVlL7OedWBK5TNoclqVnxST++rrQL8kDxzUhcBqzQqUvHtwSahsbj
UUjRSx4JR6vVUchebhWQkXIYmr+svA3jUnEoaaOlU/xtEwFv8mzVVVLJdyINOET7
gBI2s1OiDdDFCEQ1+2c9aFHQNEMkYKsnmkWSclXN+vrRYaKE7mnKTjvXweNdbrmI
eJaZrQwTsh9rzFAq9eITV1vsWNgmiNeNTqXbx0yv7oDznEUEQ2kB0dj5qFSikh7Q
IBREHOYbgvEVvyOVqBw/hG8kmVjtOTBJyC5R4hUpZHWEZXDKEWzQ0Mbp0gSJoJbl
y5Whxsub2s7gqUwrszIFsKCmI6jRFLS/iI5OpM1xOZUHQz3jT14pMO4xYs+Gjv4k
Gx3P1Kze4PR/wOSLBx6sQGQKktpxrvabM+M4tWotXSo68GQ0D10efY51zVcz4Qpg
VK3p1kKxagDq+3keBkSuoMYLw0t+AF2jnzH+XoeJMPNub2WNBR2FAMuGBp4huj3X
DkXFxMbEKoG88jch/KHIvjwKpOKh+HFXso2M/mkMKrVwwiTGR4eWOeQxO4HfwxzU
BDQFOyZ+7uGTyk5XrPe32/sVWylu+0FYKdjWx3TkLGQXKZr2tJpuVvsBWAeuoHMj
dJ93lfy77F/8D7J9ZpvN8e6jD2HjlvX+RX9xhnSlE852UMecdjxLcV/5m3PaX6o2
a14nz0yMlxhkB/evUr+vjkQiwyRsjMm0F5Ht+2fkWLiDl0JDmZhrFtwhcyDBfzOl
+jHVnpSDv3ZuR3lX/2AuoFcEUywGNjosSPqkKBfCUgRHFY0VP+VRSpRo2t/C1QY1
LJUl8Bsuo9aSYNxTjrVbe1nXvKSLY05OEabaxNejov+S8Zmoo3QMOsMypzeY1gjV
Qqch4oSvM+LoZerJ/Aoq+4Lkvs29TNalwYxdrYbLsbdBUqelFXceHwaFk+rqs3+/
H0jwRjYK4sE5EXeymWkCTghFJidg4+D/7P600iOyLGGO6Yd4L/R8fPRVaLclNbRD
GaI6D081xXILsXfoomxDIOdhVm7wwtx8k4haTWl64Sgag/kdtqOWdkxjHjd7bwfL
9wtnJsPFslDyUtyUWbNy/M5A3ty64c3jH8Fz/ZY3l9Lqx5y8SKH9kddiyVkh8bIr
8YHm+RbJ0uq1flVY3VGLMLi5kbY5i9oXlbYgIBEbXha61muVtq0t0DuX7ZbCd1dT
h7zmiWD/1amH3FdIA7+8TiOGC4Y5X0JPwUAq+pnVxF/hCXJE1DrwlkAzFxMvb7cK
dK3dMr3WUaSIVDFaJJK3FSiHiRsN33nU4ELJxGBzQorBa6MyJyDjyBx8W6dw/9G2
j3FZs4LPZNJZ6fltCVUXNYroagu0Ogf371KS1AtsWbRlP8sjWHKotOBMu0xLaVhX
3Jg/ynZlP/rGiL43MjdIPmeFcuWMEi/NC8QB9JgGPlLXmIID3r9PEBz95YY3+0KR
Ymn72PzcG6qBygkxpSOaVaSOFDahvoInxwAizjnuotMe8+cypNAT84QnG4L2JN5Y
MJe91vfr2YnJX5Ej+X8S48QgcS4l5eTiEi+jGl5dFZjGoSk0XjScm+JlU9OQCdNz
7W9prnRldYzqxHymFVEzYlWjFhJuz6CmXh/1/mY+tQ+r/fPANLyahpwhNdTkdzH8
`protect END_PROTECTED
