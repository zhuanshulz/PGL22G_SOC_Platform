`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C86nO85LAApQXcvDk1YdQfg6Klv7JEysmyossFAgIn734iJMnBeMO96QJIZ7/oRe
2DodCrPJqukgQROrGexlos4gcS7nsiSAHx3O1bLCULUsWhPmbmPD/jgpMQ836DVH
fTzyp/4mo/29PvlVmi8oEDxgrYysLXDBnEVZhyQv4UuEqnCoGKvN2CaSX5Ytm+6R
UUMwQ2Lrjo7FFACtaXjHarLpm1Unydc2L0TyYwjE8RBDBGRtmuyHZIVWZLGji3Pk
1wa822Aebhbxo+RmoyRCxD7jnSBoivrqtB+Vt5bF/Xfo1OibQ+1/HwBPxOAdbSFo
`protect END_PROTECTED
