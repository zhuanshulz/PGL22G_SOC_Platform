`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fjE4Ajg1sMOMGSTjp0pRgtn/Qd/sE/6Sz/g0xm++bcYe36QIPByQ5/HEQNpCf4pz
706xblLUNOtw50xiyA1btoz8ZbLV1ojaeUL+teatx9gmh+TZjVnOB7PQgAbEgQRF
O3ucY61nHKBV1b4LTpBwUSHIl7jMWzDJ5XfK/0FQhX1WGxjbOESMxdXr/MfCEBeR
1ay1rZ40LvPwGzNPpq/nBrA1C/NtbbdvqvvNsZ5uMa3tu5/sv0hhC0Os/KwlPPAO
R7MbKvlMaUYf0wr8QNxfDMzrvfCzN0AMxEyQRlQef+j6qOBfMqqLrjCg0pQM9SLw
kI2B9dAavh5e9MZKcJ9i4APOzlRlYw5n4JiK758LiAOffC7wpNqMh3GRXUF8PKRn
ECUHHgkMC+BStQJvUCv67YKckOXWLHxygs6kOuNFvv7r+NWsAhSEb1//97SchQC1
TLDNoZ1rxSSZ3gsJeFY2Xg==
`protect END_PROTECTED
