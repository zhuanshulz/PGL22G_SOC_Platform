`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WLJSGAInTC07X7CsPLKivqr8ctg25jjnE4OTvPEedZ/mEGYnY+WMtii1n1qnOEFV
m1msYqIST3ogBLlLGKNxKwQf5ZKeOIq0eR4U4uXMvmBbMNv9N+pE10DNdXC4Dz7y
OWN569O8tQ0z9rAUo8BirL3CN8nm6rDd6Bnt6yE2cfvjOtrr5Ui4AYxQkfimcVHa
ts7JW3II3aWIXzLD6yaagt6TTULpDfYFgiwjLhQGniZPx9ecQyiBrR59feXue4Hn
tS+8bDxgDGX1S8ctmlRgBm00McvObI1L6O261mLNuTU=
`protect END_PROTECTED
