`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7CpJYm9sWD06meMf85TPAqw73Ynh0Wbdke6+7MDms6ORMOOrF3xaNkEaQH4R2q+1
jkvoQCge7HxhuE43PSZPYCdOoFwY7q1aTFSEliBexmR0v++qzg7sUyC+MwSRz/CK
3O2GqRJqGdgX4gkvpqlWVlLtvH+GrBYzvU5pzUWTeEMxXn0hPq9W1lkp/jpWi3QD
UpScyHMJMBt2ElO6hXfjFi1U7wU4YkAW2sajqpvNSkB2zLyftSAkbnpXcKqEroDT
+UnL6nwZwISg7TSQXK7nB70OyjYF6gh8Um3H0PAxm9nuBy4mnMGZC9ljWRSyV4nj
Xp7O9BYNJukVgkgEUx2H5MVWmNC9g3QzHCLzGm/Nugyfui7NtQtbjH1Bli7wpBTn
oHiSmeBymLzJHXslN4MQadaD36kMWJJpK0CIvUKpYciCpwczBZK2ygLKY9Js94co
n5LjLL5BqPi12mvJ4w93xAddxmmrJvQ0h6AzyDxlgB54bP9qTCyslM3DTdkWzj/+
f3gOUqq4Pd1e+NvL4EMWmBjWWN17Nu14328GKrkjJaPEEVFroLl22/wuoKgl6ZSB
y6uOzCsmWLaPep4j1haJL4FzM+CRSFlTGBjxs6YptSwvdgNXJEd3TEPYrYu/Y625
ogYofjqC52I0/drXUlckTmARYOza+j44SolETW8zDRVWdKNbEk2p1J4embIipD6g
icKFgJh0qs0U+FArX4SRtfOJagSRvxc4bpwynmbxyuFlEFHkKTyX4Eo0SaIAegOA
DY6FBqsf7pIP+B1GbFK4v5XizUevqg14sVedXqWH08ukGrjZO8+tNXoQw++kHgfW
FaraYcc3MxIUAN53deijBPLNxuJFCLZolwvVJGJNRzDoGzEjSZzgdfV2f+L5/yOl
2Pd2AH3TfVBwkcg/g6MDA5EaZDhgiXpyuNqnYCorZt+8R24BZKUGqyl8rQlGfF2/
53FF7Sr6rWaa+whJ7qxbVuPxil2HDjNsi2+sIDynY3rK35efzY5rbbgX8exL7RUk
GD6j+Jkpc03bpKaswfoFOOXSb23+bsVN5G8nypBobyT/4v6jeDVOLoFLRmCsUrnJ
oS8HeYnB7fv9+/83UDI7oOnM6XJ+xdPXdGowsD7F8ZCZhUL51LrOgH61aTrh3HK0
nNyiVqxTFypU7cQ0rGvyBZCs8clXLfu4uErZeGionMTTMudAgcv44p73qAvOQYe2
UVvyE0Kt4W9rFwXyYZe40BUHRo9BnxNNgoGBAa3jyjPx8yr8+1uNvp3rQqp6XvVG
+d/ehiCJ2ev9in7qjeF2I61ca/lOxHeWLz4JmP8TmK5lFuXV4XClqVeYu/Es1cw4
49L+bEjXKtiSOSVVlLQtreQRhWUrCEMk+z0cVac02DHpenrCkkzJbsRLY8QbaIlG
t9S73oOueHWPBY5uuHopEq+GCAkmonW5S1ZaitwwU8H7PPP4z0m0wR7UQHVixYZS
UkQPDi3E062KUiiuXSkgYM+H1DAt66H07n3Oc7Ewsj4pe7K4rAP0y/TffZUCA7Iu
VD0KegCsDK7Mcf5OlZBIoutRj5paOve32eP35XHWl0Uot7BcDd5JVBqcCG1xOMRJ
Wg1MbQoNSk3AjhqKrF3rDqqdWEfMeRdFEOpUCNDccHf7ifQ8iMJhZ5IOupWizl8E
0w9Al9lfeQUZ7z0X9Y3DLDv88MLSViEV/HdLqaXiCfmwVHzM1NgugQGTH03GuNdX
7CYl3WCLJ0AmY4udRl9JfzX0/C9GWm8VUxhXEfAjGHVznutKdVb51ML+AOfXrl07
QNaEMfNjQCMUAod2EKnadOohM1BWdGwpek1TZFmHQhmgLjTyESM8GZU1PRlSIrz2
bXnExifPvHmYsluH8Dq8FVjzHE+560VjLnczoqhYGwAaDwFW1kI98H+nwwHANAaX
Bty3sO9Sn/NJulUqeACacOPBdXMqOKxXMjvB/He9Kw8uE2lxMvCClhsTwISM4NmM
AXfKWeOE+CiNV5ysSK0IaXA09yhbTBBHLet/0tntkHYamUanoff803u18Dg6VRXc
O3TpLibgFJ3Ma4Od89T8NptiL+d97bcZQy5L90tUATg2vInP7WHgHZ8JCcsHNcAJ
rWsOKaN119+ryHNEi/P8Qy5x1jXYvWCo7/Vhli85wpUj/eKv5Rn0HZpzELZpkBzq
Ig6SdINZz4ROOHhJdu3MeCLZRgOsE7iVXb10tfY83nkttnlNN7KDG0WZoPLvJIXh
29h1KAZQBBZ5JvsZ9aOCRD1f9O6cgNoZovUbV5vQUrHQpxwapnvagrvd+LEz8HWD
qVnxsOoQmZHcPKmOWL1WRrffN0NVsd+Pydw1gcLzdORXV1eYlBH3JwXMm1T/pOQ/
LT1WzczDuHCaDzABRJU0EtdwcpqQfrCX8ld4mv5q1LKKGHpGtTZGW2g69zufQXu3
LcJvwN3HY8VC2M/G8cHHtRDblRldm7fvIUSP7RvXDFdBRrQLT+6VJVnDK5EN0UG2
+tSCDu31+S1M/pznTYVLx+jR7stkF9UHHJadrMsv0yrF8gLlMoFEct8lVAWsV5td
EEBcl8Bpw5ltcr/gxctXY/cH7yj8m7JLtYI3MU9SzHq9CQLBsxt7tO+/YSp5gbrM
b+KqbzBEa12g8jcVGr8NRvpURRdpnz50/mF6nD7850Eoh5q4ois5ylDdNG8rb9nq
VOvvVlryvzhgw/tRCljXBw==
`protect END_PROTECTED
