`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0OeFkwO79vA2KSK4GcHfLlQBXk8D3mqo8K9Nxgweg2qkmkN2+PWxXRp1epLnWen3
q4kOIHQDOKZ9Gpgcfjzvr4Y7craYpNqcAMXmttnzwtmXzxfQLyqKlGNT4tnqLLHg
BGX/PmcYe0Mi1CdsPm6hyd/eBx0pX4n44YlQb7GnelVZlh4+fzEXzk1Qe5tMGtRJ
lg8oWCcCgKNIbBY2dcsfKIW19Nl2Y0n5oWxh/6GhvdxxcabiSLkRn6RM0259lSds
8bbONhZwK/HSl41+INaUEcCnP4KBJySDN5wGnGvZ/UwFsHsxTT+w+LX/z4akdK+i
5nilKDCjETerWMf7HdA+XTMD2HWQW/R0NvVK8c3S6zBQlyhsthzN0RJhl0tCuqgv
zOJ0EZAJE1KZVBQWWL3EKGOX6es0KVlXBV57OUFt2tLbg+oPVXLKBPclXCXPjcZn
fSGnazPOJgJblEV02FQ3+yZJ5YisDBKVNnwllRZ4s+Y3xRHagIqY5pqiJtxM9roV
Lv/hiO72xgTyPwnupfR33nWX+1jYftpf69XebwBi12KQgxVamqx0dWlnZGHaizx/
nVnE1RWku1yIx9zOA+xOPXWrdhCWv7bHGWEUkDbMnRVLLCtAnMhAq3flWGMhERtV
`protect END_PROTECTED
