`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YjSFVHn/DMs6ne6XzJTKEcHp0Twhw2e6dm0X0BrfLI5FJ1HeMsv+u9yPlkyBAYBp
s/+IVPfot7cXfxEOrKYnkzHuyVo7iDYUdeSmYoaKdh1z5/UBm4wPKVWzApeHQRRu
AjaacA7WMDcpP0SAf8V+xNQG5/lHK0PiF/CiWE6lcxAjGeUVWQc5Vxhn7ESi0rZn
Lmt5dM0N8cmpfL8pjAF22ZB/50MhSDq0Kqvv2QSa0wC8WJlPzXbwL97WKGxeK9/j
gYwS96DY0ftRQ5YiASZMsXE/ilaL3K7cdjVMyddTixV4CRUk/wd7He95Sj4lB1fm
0ReWqZ+IeRhOyoFXes5x97PX0vKJk/MdTAZJZdi69lsweRM/xVtQTvzxtlsHWfVa
yMrtdKezhcP+ki2oKD6r66G2fw772xV89rin5/mwmizc60eN0+pAhCyg6UyZdy/Q
ViH76NFuM43J9upKXiVOCM4K+ayHxWdZ5bALzC/Nou2dddt8b6g+ldN08d0nvyoe
NQy3Ysv6l33iYyhqMgRYbLcPzigGxYjqmtQwhWa3BV2qWqyE5PTFKmpZZE20JrYt
vBo60ZPtHHmfH7gv+B3qpxDkZoYC1th6pWlxIW2pMPAW86SNdRP63zUiqtP+B8Hu
frQLpix3OsxdTXSklO9SRBvGgAHc0IuryXSJx5s1QLRwbWDFI02mf7x/vfardgQe
moiiYgXS62UoLIPQEdW4ingzEubDGGKrtLc8zBepd/gnFnUEaoUsgiyBVttpnM54
PiDdJuWZYGwwfqpkN2Akp1b8j7JetTniYZ38kjlXi+LpLHpf5J1lXuc1ntD5irYz
rhwlNwNPn+YzvhL+kWFG2b8ygDWsnRRnvTXsxLAy1uekEsdTWgm2bdWShrgBixWY
4oAuK/Zq1auz5eHxKHimTFYDSm2EK4Vw88Aj/d4GJIDLoIfrivVsUw9h/soobNKe
xVOFioSSn4ZHISRX4CSVoDkCjDF78Bmwe5eq7Z841pE6fUCaUI2b/jEK8VJTlivD
nbDgoBuc83dNmZ/UCUNav7LggrFQtgZKH/ssYa5TaoOJ3sQ8O3znh6kbvAGmg6YU
WEVS7IHWehn2/QqeJbxOK6U/JpXNtfTPE0WuxG6Cn8Bo66WQPd44DHBgspxO/8j4
7J63DC8Hwk082ufXBUTmph21g/w+pag4kRJupq2idwelrKedYQsX4Pc9vtpln+Yx
6vd2bd1W8gZDQM2JI7AqgXmXbkLMAIPYyiTdkdlLpJTrLbazMG9cx+lpEoyI1v3Y
YFh05B28fGc0cHRsMwj5cMhp2gVVBS4FCcO0bbg/70vMaw3bgGNSpA8vqrscD7WY
4qflE7CfdSJZYmeGRc01gkzRQuOPVIN8n+YJaX/6KQp06RKoGSE3347GxZYAizWF
wKkZXB1Swy0aKvwIHIcsenhtxiZh89wTlc1Heq25doWd8PbDmghWbyRPCG451zUO
fukCZSXsbMEB2DOZdWeW+R1kYzwbwbEBgaYRdrGO0coMDxExksAHjFVcknAwcPKb
G01wTgc34wh4Q7l2CQeUfw6gqn9jvXKeu8+jV5dKi6TdVQyqs0roPzLB6Dley5ks
Ctc1up4dYXdesg4vnzrkFDbPPKT8IwLlOxy92exFqN26DF5qC3RLJVBaFmwBk1e8
d+2SXEs2fGtyQaIBPQiTzlXFwih7Jp1ey41+n3ty/2VWM6vkzwbh0A6JPIWOuPNf
yDEWZ7CBgrT9eZ8PNFOTZRl+v9F9g+EqIGMnFSReJOLPah4YG4UmD+NEMQPmZLit
6P6GEXioPUXzrKfdGrugnk+iZe9q49fVhXVeCOhrxDWFgVhdNrbRgFlShfErLNGN
`protect END_PROTECTED
