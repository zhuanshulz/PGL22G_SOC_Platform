`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vkhuw6wh0CAqXoNHibTFrQTzM1ranOmNZUeGNLs3pR1Kh60cCFC638kZWeauXexz
zQiIukwA4jFbxRmX0mNgpzgF5pLY5pSeEh8JCmu3VEtQTyveA2Ka5h7FXeXKeBXq
O1tFmgvGL/QBxB/ZWTk6kmS6+yYuVcfEimbd6X/JiSDPA1miI8nMjnybdIJUur8a
A5/CAUzj6yPrOQ+narIIp/+jq1CO8Mp3bqkhNT+RqXpnnet4UwHCGjbDSAWToge7
wcNao5OsDtWeWogeYf1yKtrXxMuTuhRTzgzwphb8bWoqecnCcxvPrpe0tnV2VwOi
ZdRfgtj8JGXqbX/MEcHDxtEqNiqL42a22Q4XgnFLHfmvqr/U35yCx4aN5HDR6DLi
BFiP9FA2fN4eHpjDuzZz0f0cABlZJb2bJaZmQUbhMv2V+n8RKH+ki7gO9WhvWoDk
AKPFI2gP3R3QMSv6i9NFEwmaCMFab87j+UVmaZkkJC9hbvL+zSfpPpOgd//QMymR
MVEXVRhtl1/idsxyJhORQ6JHkzDc6KtmTmKzCw02XbXO3ON1nj0vs8b1T8Edydfa
We53BxyvPK0Hvd2L51G6eg==
`protect END_PROTECTED
