`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VF6vGmb3QvTx5mNVxGEe5FINcoVUwe5QmcCVQLlsVdZbJEhxqxS3d8H52GYUPAIW
QF/O4GR0ORyXHvAVjKPzqLH2OUWNsI/fhxUX9D8MuRN4T/qmH9f47PRpQ/r/A2a3
BAqnGQfJTD1LlkbJdKipU2iAmNB2F8iAKcdvWWycYXR5QXSixFe6r8H5pvMP1MNl
o040r07qb5XtWfTFvYBCgdBobiisb5U/RG10vHH6o2AQVXH6iBczzkA96+1qQ4MH
wy7+USc1Id05agZcTaZg2UVGcSjchrG3sSXKRSvgFu+L/UXTdU/RE05IFDpFyYbe
nqm9zSLBixkQZaU1Kh81OE62j9wWqo+6jZPgahl3w5c5JIzm/2wUTPWT7+0FOMbv
bqEok4+robIyUgScYfDOLKjxL6H4dCOt6DqIp8+bfMnRQaceb1mCTGS6j5GV1o2/
DeI6VfRdPhi5s7xPflh1gcf36S8Qx9/HkZSdLb/QDGLLSWb4z0QII82i/47k+Bbc
gsAL51ztix4bxzPFrnTcbfl6BImcoObf2kn1KMGkYQAHKQYor7ybyrGs20Rl33OZ
rltCDGZ5PF5rZZylCHeCdjoT+cjQ4fUlRou3yTfrsE+2FjWLF1mJkRHvaXa28UXG
7OvxLQnlvgfpQR9L0MBZpZ4hNsUNdGogmHIKqkkh8Fbea49YI9UoAeB+E0owwovj
pl23/6cOxAoQYnnx1Ged76nKXcZK9oZwKduPZ4q7gYPO+2EVONjGarpzk1wxo383
VKKZNiP0JF3ZoA0Cniu7br+3FyC06Sz2PfnN2dtizCynaUr9N6aObTizQ0FkQlfq
vDA+h6yJZ+Wd0cAgs/H9XDwNqeh1P549EOXMUs5skKGFQrhmrL6ZlYkOA0jELOfJ
ndVoZaenXhe60sykk09tfxiRhbS5ebMlNhtgNMGWCddZ9/IZs79KuD/T8R6j7zpp
joIoWtxGmUdBGeTiwANkwaWLSFVxsQylCl8rM87TxKQ9rSoqyIY94KaFsMhl/rjn
bd/4eSS4+CN9Zj7T68cy/hqluteQOoLJAZu2jY6IVUbWxLkvebsuW9oUb1v2YutN
VZFKSsFbQ4NK11de5C9AdSE+SvHRaV329y9Rbdq30GWGsf6wmi4KwmU4id/Avyxf
GvTTfqC1CIfpprbxKFnk3qR+cDU8wwK8qXyHy7xw+QRsE8Odmv2xQZWj06houDX8
FtkPxTYJW2hHs0Ity5Od3DmlvvG9AnUggYa8X5bKLRy0kB+Jm6JtHWbJfU6GZhsc
8vK92MjFkKkKqyWW9rTwRCpypO1hmOXPoPIVMbZqnbQCh/plV5s1VPQ4oP7AdxOc
7ntijYoFqdyBWXCx12JUjNIq29gldLkowh8XgrIB+Ph/RT9fVx52nc0nT9XSWmZV
3VhIb5wS8LjcJMV4+u/lQuivPXEOhA1S5yGA/w1QrZCi+he6uLEDeg2vZ5AqYMQf
GbiB9RrtOzVkuwx7xLXp8uZZGCrNrZBUYbp245mB4BiNK94/tDGcusArU9tluNPb
Qi40YUmroC1UkopT8rL6x3TSjInZSkFfVD5zDLnhfqGqWP5wBIwedBWjwpSSPHx+
7oXVnW9cj9azku7GakDLZkvS6mj21UIrpDIUjUxo8WJNyLD0eHKlEEZjIIZ6fJ3v
tSP+GE4osDE9kIa7mt1KedIzciRPfAHYoC+07exyrb7IROcs2CnnxOxe2S0jD5Y8
gq5owOu87HMieafDeIiqXdSimZKK7xDXZlHJZmVRrNsymN2hXW9oMnOF1wF6GE+W
c5pdyvLwYUxY3hmgJognmticxAIAgcJqlLbil8BfnfWYZ9Y9513c2AtwufS9B3yB
fayxi012AGypsPaCTuhJwbyNJOyOAFLWHHOGcg7OPT6ARR8YLt1aWNhZCNLhrhm/
TZIxxO+u8Vh+wTHvHtLoOU7RyX8ayCUt5SkWDc+/LNNCBtCk8EbYE/ZuJASDn1qZ
h7NudTVGjj+2NhC0VbIPvuhzJ1cAHmkqfO8VjggSSnyOQ+SGjYcq5BdMT+JOrI1T
SyrkAwOGICP5DU47Vv+/+jf4HD5OxTKDQzAobkds4DR0o7FVZlsxthE7gfxXZOCr
WTpCJlnoagxkYCgtqBRHXjHaZxT8RnS2eB+RtIblv9umW825IbbnwbPSTZi920f5
i+xghbVgeeZhnyIeTwZRvPtuMQhzEWIdLbOQKS65xVyjrehkRa9qTwrW0NvbnDYN
T6YN4qrqKqKAIZucyml/Y1hVOj+jHHqrWJUZcROB1VyrOGX7KgdOG5R7Gor6Loup
gz8SEX1pVnDXZHSRqelmsaDzUkf9tbq14lu/TV8XdcRIHgrZO0hrfK6aOp6OexjU
`protect END_PROTECTED
