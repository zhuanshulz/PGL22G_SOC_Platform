`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/OCzqI9Un+7q4zNLj5bTYXgaj4DXk6qZGLwpUbDWErpYZo6HiH7O5v0DCMOjPb2F
GRs2D0bg9t+tnbUtlUbGdPByC54cOJhKC1DvT7ubg3Wb4rbMb9NhPrAwhDVbWtSV
5g3SeS2u7XcBlG3zhdjqaFL4Jwu5HcYqHtkDz7IydA56ZqztJz0RvaSi+qyT9yM7
H396VopKnGdRC3aRR9kppAiBNAA92T0kpGdthbOTBP7onnylxs+f9cagtNTWna3a
XEHvMOLPc8Sz5SxDzmEQ+K8wN4MJyQI9oqewaRx3wuJUuO71xm1lw8Ekz6vC2Ges
8hXhCXY+LHi5N0I2okllcxFs3vRQTLrsX9SAGq0Yqp3EMe1mcWjIIvdrzo6M4yPK
vHDzOmvnlbmD6LawQUDBkgv8tsyHTCHPsdLG6SDIgFQJIEUTWI7f8auD9P9PRFh6
CdtcC2MjnEYc91jvr34WLFp0V/kVtHBcBCxq4XmT93Z7zmljNp/jTWSdbehnAaqG
f6MwHigy2QaxuM+79ohq+Y60eJNDuyQq5lA93p5mYRxIoFEoxuKTjFYle9sJDd1V
yCcg8nZZTVCX3leyLx6x4CCf/JPzA5j8FR3wYKK+y9DiuvZsdbfoWKs3bQfeRGo9
`protect END_PROTECTED
