`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zdxKLsFfQ9aQruSsq5PknbyXo30HcD3xaLCx8qjzLkgFu2t9YRg0sUJvY19DvJ7U
b7qEGejg4zkzY9T9uceEC85q4ONGqORXCabUrrZ13YYZBVlG5x9ckzszjGgiUNuz
DdNrzfSWZezNR8XAaC8ZALDDwxCSxefqGLSZfAZR0VEsnpSz6xPvCeAu0ERJE9Ib
KNBaC80NJfig27VIZ2qQ4kWScTMEAYoyBpSMHNKG0UkanJn3/4aG3yRdwZGqZNRM
sSp2upR71QJNdIX5/jbVEVM6kNGa/sA7EVnZ3qJbPLHohVlmr5upYgTfgDjXbDQn
iHiZmjik59c8rr73nxOhOY7EawvEIoT3pA9Mao4FKyTGBIzdKooP0nednyEMCLsP
cgrHr4NjqahZsAgZDiXDv+GfYbtbddD3g5rsnMmQs2o0p38hTuXfu2RmwXwmSaUM
4Dp9gYVypa/ys23ULFo1c3OjrotiFIzOd7WLrobmXJhE+5TbPrv+z/AVFtiqcz9n
PnRzYelnB/PQ+FEVAYW1kE+7Aj9lNlB/iP26GU98Xh64SBtTKmf5LwRh6in6vVre
43ovm6WxjxRk9CU06QvG/wcL7hUToqdPgy9xjgMVfPh6ElLP8vYlPyuGwJN6QOyB
3NdCUKfR9Evpht7nZdrkZdKBgPmGqAmAKZUOQ9a2wRxEzT+B7sZquc40bBnelYol
sHYigFB75IpWSikbQP6eFw26ruM21lEzrlND6pjjIha89/WjzQfDexTEXov5e9Yp
I+4yMkJt2FvT+aH4GCv+gq5ehAK/fcjGVAfOT4t4hsarkmWyluCdl1hbmoYyycYz
xIA+MmjBZ7D0eQD5Y8Aj53kRpUFK4XEQB0E+qZB87B/n2t/147T82rb3SNda1aET
3wjdgVICLhkASf/+Q1rr8jPmOexk2H773WVYzDZHCWZaNzMZnl8dhpepBHySd8t2
cqUFS//8RR8uQpDPZ1HkpIKebE03fnrXOmXiGQrjsS4vrY42fYqDoJzrbaabHukA
yWnxwNR9yyDrboh0bZwlQl5Xa6zdMBUqoJjI2iMlKu0O5VQvj8ii1DflS4NMkMQS
nRATJ3ftZ+440849h8mFT00Mmqcml6WanIZTTk5r+DdsJ3LJz+VXyq2Y8yHMc7At
UpSRrJZQgBt8YOZjk2lxZKURZPzctrCI3ZQ1rofvjc8KfUWnEzWhnQdtnEn1PHaN
3Qa+wYPYNh/fLo5okRh2IxSsR2EnSbHI4PTaqO6FQI/8OmyR/3esfq2JOLCEZtaE
K/Q1wozlFQcjWDQvES3/ziLXs/wwzRI3JnB2aXzL3dzkB1YFHX/wfU2NEJnhbNr6
iviVNXBGCYoriVJf5VUJLUMWYKkQDm6xSReqAX4nt9Et2A9rd4a4IuDheNvfeK7y
cx1POFWYC1fYCnFEYREK3VVzNgzJWEPiqt/PjpeDuvla3WP94f+1QGMUPM83Q1tU
iNaLGeksMx1t+STLZX8YYs5bqf+Ryuqm8mImJz0RZQ+38IozgWnBj9LfyHwm20EX
K8agRlDwn53C3cGNuReHE0u5kAdKZ4G3VH78p1nXekTm2bLqHuCeu+vcscRMlJdW
yk+YtSV6NLtZRDP9PY5c0M2Ckq9BNGeBzJKR0AiaPEP5M/UuwwPYnc3u0H/LlRy5
AQDf5otwxeyYGqnyCCIgKj6/zbbUCbQhc/N9rKepIWcu7gWDVPDICGeA35wl9I2U
TynMFzYQgHNcsJpFIJxJxUxLeJzkcRrTyH2dUQ3FHe/OHnnPAF+qlLe8yLWkF9A6
4OejvxFz+kRGnr79gHSL6p47/dBJa13XEM4qW/FxHgucXMlSK9m7jRKDBUqFYKmp
pIhY5tGJUpxppYqAnO5yhvKPs4xhjQjeC4RT9L/GAwaUVI4RMNlmZdVbjyOWE5hY
zqdCh8cukF3FPfS9tOLk33y8E8U2zu04Z6B/VjofRZ4YOkuHYhk0UQLcmTUQeZwi
x6FNFhEh3770MI3hTfFAvURzClz+XjcVDFk2XcV5BgmP2YbXe02MzSf6N489A83a
oNJ5BwVELGDLDYcQn92NVM7ZejITwxNCGQ72mIuThI08vGXX7CxUaPrVInpmIOGS
qwfzlJnAKAzB5a7xQCz9gq1sYnCvjaQcW73H5Fo467Px43e3SyAHqpcKFmGtzz/C
/HoMc6suE3nxGpffkIyj0VJPxxZa5PcxjNG+4n+bmC6IcADBIKqFVITaEDisy5h2
o2v6SjR52umGuOc53H95P7pibAalksIbrtk8OcM+wRRhLDF1FrQBLJ9SheXJyhSi
511KNWtKOQItNgF4NmL+BD8zytapoYsj3a+Ctv9pH7PdbL4JaPGuue4TWLAZFg68
xalm8/atCVJiFRURXQyuCbZBgET1dVEYlrnbzeEPHLmheNF5Y/NWFxdyciZ7HNqz
S/dBgtgiuJlrOdO8REjoJqyYCP1SQ2Zxols/abQtxJm3LdcGzJUGSL20Z5dHOJpa
eRPzLb/Yz3/DfyFhvL5dxCNH4Gucs1ETcxBNFySTaFeSFWMT8FFqShlUbCy4NXX8
Cvh1RDcCBwsYSEgLTXPplszgkXyVf+TNMME2P2JSjkDlBmKdZ2MWEWkcgFPUX09r
FxQnozxrPINlHTJYttCuj9Z4qtG+oCcroVpa/bjnskGSGzGxKX5HaARADsqntQj2
Hi5xaYzRY+MMmD8F6uqQMu/9avqxqCMtWae2a/gI0UMEtK4Mvs+aWLjz6OirRZXq
j8ABeoLx53CWO+mWfnULAc01n2rVsGuTfCPn/14z3FWLh7ZHIxHdN78zsqDIkYYQ
qKyEQ95KJHerQjQSJgH37Zyzj2wvWJePkCORfs6pjudANZboi+DI7uDbqMNr6fXg
TpWvjQRK+q08fVeoT80+N6+C4qoYk6MpNN6do3dJjE2iece8DuzpbfHYqAdu6XdK
Mo8QGhKQrkG1+Qp8uFajKeGfqTMPqNiuiNB0aWIV4Cl4t0cXif1kLHrMoRpA4SI9
5MaoaqYr4I57JnBQFHVeOSBbj1hyB5K8+wtd2SiZUkrVRGma1RFnjsHK1SIFJeeG
xdDtJr6uf82YJa8fcOmcsASVybUQSFBROgTjHubiP8NCtF3CPH8YGE3ZZx0d5U1u
mpIGNUXYPupj5dmWOw56aZcR88VB0KSuR8fG/MHYthK2Et1PgKpPWCS3P9T8GuQS
Allk3yRCXIzPdNeFuzJHaFMms+esVKnv821TEL5kKO9acw8y01gd1JCjAxsrUnGV
jiJr0LpqJsWNlomYD8O/KOCJ2NUH0ybH8iDDnlbqgmupDroyreHbBGaygejs/I/d
oG3OAdqsKOOI+0y2yaVcYxc3v2os0eoV3idREEGk56LbsGFiAeUop79hivlMOXKh
EBkFK98aWcURWqQibt/DMNomA6bolwBkd6MJ8JBA7j92609HlTYHzUBW2i3CX/+u
f24PxA78B30ltvHu2/0u9K42l//ZRbo8GeX5aXgo8Z4xDh6isR28BzDcQ2/LTZag
EVNzj9oroQsq7MvB5uW8bffdGVPuMwGHeHYLC+/gXilaDxv1eQ2YmJv+dwrquW2l
pnsanLeK1ni392df1PoLeWZnFWJqLViyD8lAVe8Vp6Ae9aqthOcC8bjHFkVJGzui
cq/IyDF/y2nZLZWXMGYKP5ogwLYevHzlmnXGXvfDPQESyTopyn2A8SPfGgbKUsPe
0WZMZfKaUS62EvREdRmDXJG4sEBJxA9lSwwmMFJ+WNfFzTFw7qIGULuMGNKGOJ41
b+hNsNFvAkdi3HlhyhD+BshWJWn7KhBXeal/DKpWA8cSkDJv8siB9k1oC3O4stVe
oXEOwtaPNfONpkrx4n+d0clbyDVvOZSS7inzD82AJz12mjFaWVPyzBnMnByGz4vN
Dc/ZPA/HvJnubkOc3DOWGsx6i8lukOqD8+OZhE8yZ6HNzO6L+AtucDM7Id2zKxz4
QstpxbPXMr+qlc/zqu1xHx6sXlkfBUTQ3f0e1/wPwYDtf9YrkCGDN4BHlf/3CpoL
U5fm09FgbR0rZha09vhAN/W7RyRTLaFlxmIj0wZFMS3LgKWbp70o7YbR1LoGZW3D
PtqI7ccqq60plfIv8jt/2pzEmXZJP9PUL5FYddWUY40bkUBa0cLK4XEtXvgQ2tTK
v4Ed5ht/mXTH8Jcr/E+uBxAhw7bBN2IUaL6PITUoB6vGQxKywCKCgcnMaCgVWf66
ZepsuAiK4ak269gNciNsy1jJ8b7crxhgWMOnIny22vvR5xbUh7v5YIVFyLwHw/rp
dONt05Hrq4YZlAMwPc2HBfROtqOKMPEeKhIsdBOhF4/akrBTaaUE6YLoptcD1cMQ
xRRkRqOL0aoAWIVrLmsmvIpfQZ8krXOjFpK7MQNJNMTDgJ9l7X4J33Zxw5QtPAU/
QL7SWYl0DL23wj9GEWxvgg7idx02x4HDuiY9eWayLC668y6b5dmGdcjbJ9pra+IU
0EIDGhpv/akwbC+NOO5sEnYtwDa7uxRcHuXFKuT3UlyTfNu4mPpOHK26cVCctNh6
ThwvFcibBXy4YtoUj5W29rOjeOxN4IslwAJb6tHcSGg0mL1ASNx8sEIxMwgVpgFd
lXd/FLLkIYm/gELRr8z5Aho3iNmLIZiQmACG40azyHFaCnuqmHaXocrnY5ntOKmb
c8dvKlOTmThb44WMOAkuGm0dyaMVtlfld25VHepedYGN8IZZEqSMWD9xmBvCA8Z6
RO11k/pKWbO570RWGLfPlBqQydrK1bKjR/09Kj4Kj5sC7KiQxPEHE8hnb6O4s2eZ
sRbRMX2uxkPDjlwHwsF8cgg7yzgpIuwJDBesN6wHx/J0qcP9cQy1xzs6nlt0MxQ/
eTUcp0d3ET1RL/QdRU3isb9aXihqWztwhAQUMehNDOu7akZcPvUx+5tV6RIU4zky
8OwyvYxZF9Ye4Kn5VMUzU5SxPWq46Js36vOIu4nCEj73NTP4MLD9+S/3IMqGkyL0
akQ9t1Wx1X0y7I8/BPYZG3M1sEPENanG6CUNliWHLgcpylrSp0J352wW+NFD4gy3
UZg8OEAp9nThO1Z2kotUP4o7TUEXVrT/DLTS5/tMh4GfNCAfAkMsoIXIH+KsWHIi
qdrnYBbFjzDSdOAMyEiAuRlfcg2hbNmw2CR7wFP2IP/3sdawGQIG/MWAmgafuzSq
Rhch8tSeO/u5UeJw/PBVS76DSbN5CyzNCEbLfk9quzmF8d+6rBRA5QcMX+aS3/93
5ZCXkbAXpJHLQo7GJI/JHieG4iZ0YGKU88CRz7yuOuA7oa49RrohcedUR+DS7a9u
O4x/7I9lK2AYL9iYuuhHvoRuE977L3Z98ZjpHC/5E2+4P1p7HHwGSZPw0fcB1BaT
+Ndiulo8pSTTnHkDLEd81Tb2lPcp70Src1FZQNdYndxv1MakhVHzRT8XvaQipuNo
raCbdDJrgUCm0FH4vrgWx2etZu5FwGF/2wXQnjgW8Z/19DBEo7vBBygiM2IRhIL7
fP//Jecz5wX9sSStTWL1rEqd++NE7L0KDxT9Db/8t0VWLtIxj8luJhewOzjNeVRl
2G/yqONAm+GjYeWyaWOYKL6ZSHDoDLiftX3VfiCKM8olcsxMRHPLYsw7yX9lQJt/
wy6+9RgVSNuGe1kF2tMaGAMllxucej2c33eVQKuXi/faW9PzMrei6TODU5LnVFcJ
M3ncux6107Lzx0lz6Ap+NqzJ76k9MYtgCJUiVy9stnugUSwRLYRc4PSOo/bM1DFV
sQUuMErdu9PjUQzBvjsoMtIPhMsy9GVsET3TK/O3FG6uqCWmj9wg+hfrUC7scWdc
eaPF7h8q6Ai5FGUTIpbEBQg95eQ0KlJDaZluOMir9thEkeWCmD9YlEQlbvy+shPi
u/krEhpWhlnFCva2egUJy0mZCB9LL8snZafNDzjlsIxX0n5M9SGHR2D7ji326QVD
k0RRKLhPDFG4NSgwI5bnEhu4DrodZDMajXSco1pTKoXuE4WWb+2MDQuXBiKp/3cy
dA7vZVjxcucTdbS66iN1uxXUIwvsbTWk6GEZF1Iqxd0lT+7JDw1zJUZLtkBglJnn
TX6lJCEkLB4OrUZSkvuXfM0sByicqznBg4I7qNp8rkjSEAgdK/VWjMvMJ2wZK4Od
jwjPqBLbK5106RJCdouoli9BComGCgHPVaoKop7bBoZBbEIHywjC+FL20B/xbwd4
bTKAVP82Gen4YGOO88fK0BXdI/vvWedYQsHeXF8eQSrRdVKCacZ9LSIgmOcHLM/X
UOuzlCc4qdKvsotQuU0OM0mNtAdlDO3OIUvPTWj/ZMIfyNJQL2am4r+R+Dv6pkht
9fUpTfHsASZbQr3ootRAfpKeSDCq/KbUOYeEuXLnQkqnUgTS3fatF2MVYcfQ+XmN
Q4xDBiL5hRqMdHlZJkV5wNmGbu0i1ZrdKagkTDfSQOP02W3K+5dCOOG2P6U+IvVa
Yk8PKPB88ZaE5yQLH2qqSo+nxF3BFVSTKE6IkuYw4ZeCWQY049+nQm4YNms4bf8g
frAzIQMhERwdOrcsyWNXzDv11aVyD3ycd/CEqf17cz35RLKq79R4VZBGjt0TKmwX
qtROzfcc70RxIQ3gE7G9LmTvlKVN/wr1l4BJMGHhPSIASDkz9sQ2Niq1tIl8SwLh
0oHBnljKeMPn4PZJpICD2jUdrhf5XnAPSLOizU8hiW6gCtqnWVjYtn3mntEHNEPz
lDi6Okkb6kAlyUv8YA67UiG7LmwRR99eyqeUaWWYHj2YcyaWs2IuaaG4nM5dOinO
D76zye+hnnD2CcQL0uaRvVkagorwDU71IN70uaeuELy3/OVXJEBGbL3fyqPxAiQV
W6v3x25PjgfhEXWlmcxM7jKzs9aXbUq4bK7mQsFGUPO+mt2OFUaFJVDH2drs53Gx
kEcblPkI/Fg07y7v8PWhGcm2RC0ABGi5wzlpbOYxcjABZtBEw/f6hCcbHKtCnFy1
pBsre75aj0CQhLZaQK5Ke3obYZ0Nz8Y+QhEydd4y00NS8BxPMALARmYtxo1Vwlmp
4q5rzBI30ZnlwHU7adnBspVdP0lh8NIyqBZpiGmbPa6AbD3l5Yl4Yd+wDmu5VOnF
XfL/BG2ViQRkmZajClS2fxUqGZ0Kaif8o9Uiw2hBI/bkaFk+UYfrZfN/9lOTQ07L
Te/EawTys2I2qVC4QxpZMsFzo2gukphZdzotQ19cdyCoUHri9OeB9a6Egou+zf5H
GIPfaFo2Crm8emHY/722E49BSaH8PuIpgg34+kLFUBjpE2w5ss9HCbc62CZ3XJRl
71acgLQfSPIEroKgT+Bu2KW7QSudCAlftCdWRBus3JXHqQ5/7Rx8MPwYQbiLSv2e
Hq4tdT/qSTjYfiGufhsars169nDbOHQqJ8ij+X4g1aU+iAKPSdgYWzgIowuJlIqx
daulmGXURsttGT9pycUvOCFPAgd7vBHsHFCj3t+PMfSHtjr9cnHm58UAuzIYfIyD
iEQWUwL6ccuFe7WwXB/1beV/hE6bW9Tv76hUapHRXmlpcoPkLH4697zXQTRidSj1
Re5CPErAHDzRAEj5bGwe/yKA+7lu1V/9SPXSg8QnTF1HUfOOcJv7eiAY669JobTE
s2Ff3iz3UiE4yv0StKpK3FRTBdVMwKlXQExS6yuhdidzjS9KuuMqu8wLrDL35tqE
8cEOwKgW09362RQ/6G6nsjRRCWHPnlr/SvNdSTknPFBbMcbCfrIi1bJJ77MECSiv
ayOl50bIeb5u2w2JGC2/4l/2xztvXZEzcVch5fh/0lwGeBG9G9Dmbt6fJGJwSK+a
EqeadWksK/6YVSNEQlJCV/l+wwPoArrJyTryqRFYsS49VmWVPg2EAGPLXXOmaew4
uJS+ilsLVUXdDdN4Vr1S5QknYGFSPVIZsAC590nVyu5Xi3kKJUNOwAKTttZdyGA5
g530m2YzdK4VV8sZJIgk4OsjXAZPZw83dTIWpdgJqmerG2E5h5KW+q7ry2pzlAb5
Ae6UY3XUY/7CQ7WxQfBm8HFj3cV3Nic4hETAyoFqPBhYmdKfshtsVOt9CL/O7Sqn
hmqBZwNADejE/CFCGIRW6UtcRjoa78dXwd0rziM6fYeUsx8fWEc7fh3XCal7AYiS
AfBKC6H5H/78895tDe+fe1BTzy7Kvq/AeIp6E5X2bO3R6RR3rSjLupQHge2TQy7D
VzMAlQtqid81Y8nIAJKPvDEkqJvivODmcaLnI3djNRDravsSLp3LQkRjD4ctNCXM
/CT4jverPpI5RItKMSoJtQuA2rwyOddS1MwrN8MGWASlLWrlvDNbm8MV1RuI6ZHS
EaXqYt9GSgSFmUSsYtiFtGQoV6HDcEmmiQ9kwx9zpijANTlqpHikzxPpxEeIFvM4
eqEczLqCn0CWhVhLFeRMjn/gPv3/7S/VW+eS7QoNFwVyi7vt2FR5EILp2T6LLBTj
jaKXLm84X3BH/BdtmCl5XL70y07A6fk6JIs4Ar8Y9vEVgrxqbHNNWeKE/1y+6VW8
rH6XwtuBkUpPEJC3vVaNMGEU7/qqF4BsZRq8PJlvhSYMR5U3iZpyrcNP9y7XK1Nq
nL8s9Z7gtQ4fvhtfE7Z/LKsy4GHGFPr40WAtSU5koLA0b1u/FMExSeAe66UCK4BA
/0SYqeufZNnSH8hwSQi8GhXHzt8853gw92tNe45IfdboZn+lCM0XH1EHAQ3BjWSn
j7o2clGVAMhvwiOVvgH+Rm805O9nkdZFFbXNLfuuzzcDyulZPua1bVQQZpueMKcE
2PKp1ZOh37tQT1/KKDouCYmVu+66d5d/Yh0V6H51PjhXcOuzZp9DvXlUx9jcQ2GE
UoKO26Y0434iw6OTY5ooEbFV3/lFOVbt65wXq5S4WXeg76iCSyabIWtRCqFKn6Ad
4uRVlJAsgbICUA8CQHl0s9WlMIn4iDWY+SbFSXYrjEKn3jwl1UMnap208Wu+QaWO
zMlRsomb6DQ9AGAZ68I8w8zKszZfESBRIfqMdd9EAmDvaxAK4znY/lZf7W6BzFwB
YT0bnFGMpLtfVxS0yzdYib5a2bRTUeH0Y+KDeeAh+Kwpv3AZsuxr88D9HOW9tEId
qLQuEGSK0Em9BR/MHnaH6MoMjcKAMi3QuJSPzvne+/IrT/afJv1DWq90Qwn9dp6m
iXbwdJkHjw1eztZ9Wi58hyT8pEuirLVfJdC5KEHwA+mAL4Td9DHbn9DUdsD9ITfg
EK6zQNnH7r9eUHJw+i7Jq/vxTaiNqh9pbwF7Rw6PFnOjvxYOrizACPqilEN3wBhW
czs/zy/LXEAzJ9njIVXjCEBOfk47SvCxGOHewY5+zG/d+1CJBPUebMAKFpjMa5yN
Rijco3N70JbjJ17/4d97lXJ5CtnzfBWvODH+FqC/rcWrKamoEleylx+//aKaaoBs
z1372hZ38iO0STGdt9NJwsBLG4MLEsPonAdbgSs+kwuq9i0joi2TCHnjwh0E8mLA
TqEDpnEjtoxZB+9ShqyAZV39cwXAOkEMHZyIPq+az9g1g6tdcj7CjBSO4oyVt0Oz
iTMCwq2UiMgoPWoqEH2zT4ky/Z3GlXi2zUehCvjtSYYe/d0et1yG7NB3oTPMqzJ4
Y6DBaWCvvSRmJIIPBL1V7fwOMT5DozVplgdFHZh621oa7fkuAY3WfCWe1YX6wsdq
dHq8TsQU34ffDQ97HxJ34KF6ImDG0TiUCBjEk5N8KAxMc2gSeE6r59MRzxWj5rFz
gC/GPmXymer00vZEeyUwVaO4EyzHAPNzvUG99SSSe6F+2ili4Mraeij+sUF7CPZz
SfhxIB6Qd37ywu8oGREPEgPNeR1wsrE6++Y2ECTfU85NyrNvafHca+9h5RbI2jFQ
DcN7F6EU/g1PaH7FOyDqSUdbrtotifomlfvj2TPZU9f8Rd1DGxaamLgYGSUouHPo
d38SLS9/cZsHBOxRyG4pC+6GEZYM/EEdihzVeg+QKBFyK8bbIF1i7ZxqyuiocEmj
Gsrtr6sbbrtauoN4raVcWbsNhvOfO/FM+49zRhFuU49InjnJ8gcVeAeTn7skOSag
9861y6+6XjYxaqYP9GxU0Mju8LMsoG5kcJE2suFjmbX8PRD4eOyGyeZZkY3iF6FP
6bULhQdiMfUY2ePNxGy2gQva5bSWv34C3T4NWVlBzgUs28RtL8ovVIuOT7QZabpk
QbCME8kIHXHzDSFgtQIAljsSG7tCEFB1ocM6Zj1sS9ofkYnDzdnclw1Xk9w2tSe+
QGA7g4G0y4RZCecXWDJ+A/psLsQznMJ++cYDMe1VMMHQzU+kAzDVqdYfYBQR/ZOU
YG6xrufoTuKf7n5mlfCo7F7VCTN+GLrQJKX5spWqfhXX8k+k2vbFEIIuSnNIYbsX
j6npjbpY2funkD4YA23T9nSGfFS58TOmRDEKLs8Bts8F9TE9KgeJZqTpoZtJbeS2
o7hWj+0cxbvF09MTVHTp44PKjIo7iqHWCNdQ2DirjLCzOq+GEFM+RzAVorrmtCQi
Kqt4pZ+t73zUD4jVRJeaSoHIaf5AIWoqRAHgNDTAjRLhXX66vVlGmhVDi40iLrdw
eaTkef47Y2xD1CtgI7rRFS2Ym5HdVdbLlpNyNeEGOn0fpH1sksjvAWSVBSsSgTR5
iObIAoHnjWqZOWIgzl2tfAL11ViQRQLDJGy2ouO7+JQJc9TZPI74pN9wDRo/AymM
EjzpvkxWryNOd83mlVvwHqWpLuPWgzUZwWRuaBp1Rsqw6WLd2kp7JaTjjAJjuFC4
51DOb6gRwiVE5zt/Cl3/fXNz5oiRo9jOVxheZcZAmA/RTW8Iup2Y/PI90X25yHJ2
L7wX73lzx40eUTbeMu3UkOeknYfhwhe7y8BMVThPGVAfGGMShpSRWlZDgUc20s3j
ONhTWJGBN943Ujwfk2cQpaOS3Dd4kcNshPXmF0r3kablHCEamz1wUUlSmIxWnNrD
9D8ieUoOdAOxNcao09CYS8912dYPOtSgR3cSKOyPDh2gzeChaHUvD/UkEguHSikt
Qp8KQyHij38BUyGhkgiTjNEK8wIihpAY4Lu3Gmw7Uqf5qqHHxdBtIG6JPq56AOCJ
eu9hghJTxl6wPgnh3OfTBKTChsUTcL+sskpWIe9r+sqIfwBdjJcCwsgP4vhNamq7
R33pJ6mOPGiwjHSv2POFnrh5wp2vrBitZnHQrB+wq3AFZthrZFqsxqMBnFY/4sgZ
tKxzn/GxTwZYJvD19Pk2F6gmNOFPEAQPwGqZ6pJqdl93TuDPMFYPp5k00DuxsD7u
BaGGmsweGYyi1zCpsdqS/Ylfn3f0+IDtZnIP8cB21+2+zrv94rsNXeFlHT+fVHLt
IAtFPFtsdemV42mlKjTGUogpjFi9gueqpyzcKYgam00y7W/oLUis1JrE+r/s4hsU
jSMvqpqm8EacH50Drm74U/WPmUE0TPAtflQ1P2bGHEina/9uJHNcbWX8R6iFIFrO
phkakg98aRS9TVy8W5pxurIpokC//o3MWCvx5FTrQW8xT7U5dENhZHfihr1pzMky
VxjNgeCXQf8GNdbxgiWBEcb83mR104cymelvclq2NzcKm9VNYpXcSO2oo+8XIIIk
m1uGRSdJUOAo89cxypxOf99lhfH4PYnjEyhPxEGGa8ehrpNK0Ll4amcruPsjensT
ueH5WEPMTgXxi761bGI0bGgO6s9ip4oSNrFvvnLxMy/9RpiXULC7tl4Hhadim5Dz
+Ws1OgqnsdaVOxdPs17hLDnGXFFAAl3oaMoJli6i3lTYMtwJlhtVSJmtU5WzHwHZ
WHJ72+ziMK8zflKL/6TtF2cHulb80Ll9boYCDl56PzsBfrxXHtmwyKZAy3P8A2ON
Ra1f0uzzdE6ti8nls3FFAOZP9Z9mq6ERC6pwZdPaKbijoBZbTmxRdL0+li8wOOdQ
BCFj2RaO8KWWbENxnTq4q5LJjfvoe83lka8M3w9a3t+uQYjPCp1iwFxJtQCw1QBE
FQtLkEznppDc2gH4y2WcedLF9nQxNPxh1F9BPSqLUtquG5HL2L7GvFcxBsCK2N0E
5FIptTK0SvupDpYy9Fsi5UgQj55DtrVKcXc7QNHlKyAjDdZQAbqgxMNEzPualB6Q
Mgh3Wrabl4RgxvtmHHccwZzhetjH9nWR5caD1ZOJi06nMPKgbDH9VZSFj1mt7uyU
7VLwzcvHWV0Ym8AmhmLczeD7Ke/izw8TdKy5CadXVqaFUtGnqiWLlbZnfQa1iIgX
VhxRSduzqlWuSdBewGPK7MucexeVFDybSWtV0Wod+mh307bf1Yo+ODiu55QbV+gJ
LVsoPq0YiCgXjqTN9FS6q5361wrju+D9qKUKYmQ1FhzZ32gtu6CLtZyLjdfD7Pzz
IGpAGxXAqLhEeKhfeZ9pcLKvTOWuV9+UxFW208/2hIyDo2f605MPQ5LLJQD+lZnr
izLhG5Fia6nB6E3j6SiQmr8WwVqqGXqXcRurEEmI1wSJOO/xLA/Og7gdG8XbSAvo
9blvDxG9g/3GgYUkvr1uSp0SOmzFqT2039LO1z4+DRlKtdv+pp84U9LPrnhg47Jd
3/HWOCA+lLWVCzpvnG8Kklbck1TYARJ4XJM4Wx28RiWGPtkPtssK0osSnwvjEXle
hr8HDfQxiVi3Q3PtFJAXxQK1mrSr6ee6y9un6/3JXHtxfTPrQNTMb9NMNuGzVmGF
PMc/Uv1Qd4BWyljBiNmCPBhMOl43ObPiccGYCsq2hzlNQIvB9nrGBhWbHjqjD/AI
FqJXeDIh5gfjllUV/8YpuqAoK6q8Vx8P1TylNMAjOhw=
`protect END_PROTECTED
