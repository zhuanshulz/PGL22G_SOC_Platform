`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
73+TtgyjZsGZZKKTDj4UdcLIhZ2Ud0uzKERZLPdAA4D24dBqxOUY1bDgHJ+TPiqJ
KyB1zSMsjw0xRe3Zuo3d2zJvSWA+C7bXe/NYnOFNHi/A3T8fPJNxk3dqqw953Pyq
k5GpFMj1h3b/VKBqwv0+xnJjv5xGI7SdwL2nVvFhHi6TVTjOimg/yQYxdXlvz5It
1dvtc/UtREZXc7NLJdxcx1RlIMfkMXqt9urwxj1diGhQAMT5GxesLbwjAJw4fFHv
NyvbFNTbI8Q9XB9RkbdyGBvORMZDWa5dsAxMfrqg9Go=
`protect END_PROTECTED
