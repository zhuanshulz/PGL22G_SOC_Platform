`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z3EVyTKI/sf7iiK+e/b/iG7NyD/hK13lV/k7S2XMSvf7mQBxgiOowjEb9LNYS0cq
jXS9cD3A1/wlHDmKfs57QzKyhqh/yelrWAOaca3HBWhn/F+A7kQDJF9m8t/bRixN
zqIcXlgEH3tIJYyp2jwicLg4L+/Q/5JJr3pKw4fuewxkJ80AfvBt86qhAOzMGyd0
zejt4W+GMkmybq7nn6hRcENLnDMbQgO6q1X/GF85tOrg9HHmRofG/yec2KyaUYdo
Med05ydYaydIbfuUnkc7dQQYPUWH2LO5M7YlZcPyLCTBs4exs1etXo0a62+zcepg
KB5vJ4Hs04prenON/7tmx7EPkgpIkohlK1Z0KPCcG5d3Hg0z9idHlnbqGIU9ZK1S
aDn5U08LTes3aYVkyybUhUg+/R38QrFmlnnfMGzsKFJXKn1j5jbihiFalNMR2xQu
csWq1B03oZatzmiEnc0KBXGgQB6UMw2QdreZN4IhxnpjNaJAj5nl6S8OdPbwbk0Z
OjzrYYKssNOtGOFASXoJZMZugeJYaiL4IDL0eYIn4MQSzKi3US6k0IC9XZmfFV/b
ch5wlciRALwl8fWW2BOL1hwfTU1KhhgBwXdFAqmfq5BndrQILaAiD5rMOBmWfp9Q
drd1wMTktZiWZWB+3nlCTvyxl5ffxRG3i+vfPA9jbLSZNfj478A0yOZ5sZWu9SsS
fdZSYA4FQ4aZrPiiOY+kCJCV9nx4V6XEPXVr7Kf8o6tqvWQAFD7Rtm1fXngOa3La
3VZzT4NJxXrj+V7z5hVZxihgcdQuU0hpmsEM1qRV9gFl962bDdXtXxxYysfSlISw
Y3Apw2BT508r59UL8Xq+Eyed3hQseH2wFtVdBTD9zILrKt+OiNKvMrG1AuuPAFXJ
`protect END_PROTECTED
