`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jWuqNgx+o7uhORlYI0KtupXBCA1So+hRdQu8UAgZB2Zhmkrvu6VU/K27GRn1cUGo
GJB0H3ZK56tAD3o34ZKEsGt3T3d+CD+mD2GXFfkgerhope+NQgepUvU4QA44VClP
sacqPfAbbzFIxGQegv6yHvWww0xQwrt1jklzqEbR0zd5EClon379f+6eCb4cJTfu
LCSCQYSJmbtrgmCT9jDW3P5EgQpalxFhWutIF0NZigZsRO/7LAurLqn07Be2U9CF
y+/jVoIHdC/9Dp9ZoL69l9D8hV1Lcm/tj1IP3OBifn4Yz8k7lgcRodR0NvWIDOZ+
EVrFxmtOWH3HsK1GAfVtl9S7+rdO2jlCsDl8Mv4bPmaezzYPHQm2dXkjwE3B7WDG
TRgGK4e/gq/cvvcR3hWSfcNhDD606v+793MdN9EaiDA35Mq6OgdbS0pPz1+NeHbc
aBQEghFPgiIn0aOaNxDIDlJAsByMjWpY5iPNWYz3SzJqyodDsxM2VkXCjDX+duNi
lgw6rtrzVpr/4EmueFkPi0fsmihLPQvbegqzY3agBrOzx5v1duGwvI0A8qtFMLS2
np0xs3zKAkp83bDUn/HBpRdv/v/89aFeI291xNhQIbF/Vq7JzuInY4CufKmpZg1z
8+NcQEtz5zNNN+Gja8zOkiCHwgb9Ke9y2oXoekZ/+pSjH/vFT12YKMC5C37+6K+N
/U78DsuSAHkxLjW5d5TR7nfieRTYke/hhAPy0CaI5Zy+UMGSZeBP4rGxfK8pNB+/
MlKlnnng6CzMarFNYoh8jOTTyBVDPki/5C5vt0aQ4EnKpANkMJE49xJtQlZSgKHz
gAMLCRg0Jybaadg2Ko8nx576Y+C3O4jXzAISn7kkOYxHWf5dOZUZl00HYM9jOtmM
w/cT84MCBAnBuvxF5XM6hkwWVcCjuQR32jsIEqe6NJCPtd0+pzfRURe89H2zdBe3
A+DVDZidZNDSQrdbFxsXi04KWTu+8X8MrNGRiJ9A9QXwUTMo3SkCP6EktLeYmd9K
/5UexPiD6I/BYcFDTvl2XV+UX8/iGU8I1IBomVZJjLbVD/iLYCclxl4AA3o5HYuC
Evnfu5f6FLAU8kCnRpoxxe1JaqUE/EqfI3nJy3ss8VuaNBzIRTFx8j1RrDm4wmz8
Q7XD9FC0jfh9/tqKz041pbZoRlI/TXWgD6R1NqHaRH67pBcoMHDRvYUVTcvlYSXG
gykLB40pp3hXt5zf4/Bbu5lwNCZDUIuyAoCoDeKaEuMFkTHyfTUCn+OUnJWYawf8
uiVV/lf7uvne2zlc1ji2c2IQDgVsIycIq7UShNm5fAzKlrYPk0u/xaH3y2UBsBr+
8oja2zm5qjDKmO/GLI9b5KbC1lXDIlPf1nuP8/3Sr7Wk2+Esg21/SmuFmEBlez5w
fmck0IZS1AVixTbUVrhZmXt3YCkfuTV4tIDDsqoBsaHUhbch4avCsIAMQnrRcAau
5CKglV79YEMGl/UC2x6rz7suXYluFuePlvwnEGDdmIBpqo73LGMlcibuoEE6diEb
2dcUwqN4PemCPwg4f0BDcRHboVJm8sY2DSNznbuRq07xWWiwlmtvSRTDj7E6V+2K
9K/YFpsHKd+3CBjg1lMmgA1Kwu4Cf6smp1h3HqF7+lcyTUzI+4RAzw7/0vK0cu2Q
SUSq5ynS6UlY0uagXPuV3cn68O8GBS4sKbMpvskyNulqga/idAypXq8UjCQy+luO
MXIxUrK735Wf8JTKMi6sp6jilmMveNozvmywAxCO0xV+w7Vaqg3+JStuAgqBYK9c
SSTrsahrBBJZAd3HTK1mNVbD0Ybd/S449EX/WUp+IDk1PRVAnLnnBeNHTj6wNPcj
3nnAKx2hBOjyrMoG6jWYr3oigif8WDt86GZAzBHintbVJF2na3AdbjQDk2m+AGcz
cPuqh7eXRz7M71GpZqF2By1fh+yG3dUKkIaQjQLsJHt649vHwuDboY0XvkG1iJI9
ouPXySpov2uUZSk9nefthWZuHhclj3PHR7DIH3aopZkUc4RL3qMqbHAAdM7M2u4O
ybKEKbLwxYg9lCvIIfwo+zgv92IzJjHVMcGi2To9HJspThOE8lbyYKEc7PvF8kBd
UxslCCJTCrjEg38sVWUVezJFX5dAEBtpjC6Xh6eah+a1/oh7UooO1rMj5u2zhP3w
NThD2xg7gEOvyo4EtgtDW+7OJLli19XhLzvSHwDWcTxVEjZ4GSyi+Fe6WVws71AK
4ZME6h7Cao5a0verCH9g7GKGCEILLuMxNPIC9d/Ivj28WlGQAtxLtd/l3cbeUlhF
1ouQ4LvJyssoTwM00GKJeAK3+qEg4HZgRpyvJeT8StYDpUJlMpva4RYBv44tTvm5
gXgg96BltyURttf9XiykNymROOJ35xPvkoLlhMluzfSbHUah//vAUpxZvt59piHk
3LfUpFizvHQO1ePLt7PNogJu4UB+tmd6eovx67VoDe6Waid+zz3hAIbSv5LdyZes
WpgDreW/T4bbaWNO7sYtgFO4O/mR4n4eLC/zw/Yc9/55faTlhsriGIzO/RoDy93H
f8zcIC7a5SrtHdbC4BNvGA3BLqC0R4e/p+RudZD2ReEqpVZhYsjBARygTr+C60HE
T2smy4Xtw2fbYLE2hZKt5j7zXVuBhJt1BFIDEwzzjn+BUqBlctyOW6DBuY/n7nMc
wYq2ZfRKaHNd6ODWmnvbQPSxsA8uh9L/+BICG/QwHF6xohnpVyHCcjdfSRl/r7vR
LBxuHxmaqurKWp13jqUpTe2M83d6137I+A+hLURrv//Vb3Cj3XfQT0LwVXDSaFK+
/v80aeYQhCuFTVPn9yiZJDEAtC3VwiW8z6/lZTJbYyRWcHnWQNA7EvyUussLORVo
HExhKJQDzE2YfS7WLCMMOyc1NEmo+RF5bcwk5Hf0TzE15uodFHEOD/zb00h0pdKu
0O1AsrD2ZdPTY16N29LGMOM/P6uC8veaMsXjTHYu09PXKuRZxnuZjE/fB2Y/QYFE
QIqxJW0KkvsAcoNCSCxM8spqq4pd/11eYvpvF6kzBlskDJ/nxVj/H9g5yZrwcGyQ
mcefVxezJ7RxPwVYX6oJEpMgooowuSdZ6oEw42l0aUr5AaEfR9tcWMxHPT0OEIIS
rQwD9Ay8At7s3QnVoULXjpIgufo+QEoK9T0T3lSB+oAvpIaJ7CwJFilqLMMEqKQE
jnEolgjQMCnzawExmn07+NDFWt3PABTiwD0CfnbKyuhRVHFWLRxErxYG1iP6ySnb
eHImgpL/XWrq60XkD885b5pj1IUkf87YfcE6EIYl2Nll9PVj/fz4LcdDv3zYBo3g
EXs/sKnogNwsgneHCMxJTOrf8mshzUC4R6jJArLyagvBnsoxHLxMVevjth8Q7iJZ
IKuAhSXES7xD/BV7dR003cckiFkWos8pVuZUWnvbCjWAOXhKMqBtNuBPNveSR/Vd
yv1nlzC8XnJ94ofCyidQZ70GLpyAzK/hl8soXNiKU1eOLXNrGhv+eMuAhyAXfqLh
JpxXsn6t8M4INzi+IS7TBVqF9hcDlmOrmB0zTnyoAMb7STiTUw3kF9NgUN8GXqKc
XnocS4N+aqusn3h//kE+Sh4DweJp1hlo/dHzFN7ZO3NIRC4d6iduHadb7RHwzISZ
B+zEhVS0eaQasI5fyBZjL+1F4xcAw7qaep1nG4Q+hokp0aEkbQX5YuXj/YxeB4JV
W2CGub8SfXCBm5eC5AfVn8/oQIo5AsgNCsTQymD/grNhujBlrtBScO0TqB7y57if
oF29lOuDjvJVkwJEOTN2R3UsckmJojF3VETDcj9Mj2+TthiFhjqUB6auczKvk/uG
iwfMhuQKuOM21e2vED/G43rXnqOqKeWyPqTx3xYR25d8oerKepjem2p7r/D72MRY
I1QiQZKR7LTWox/Tk+/juLQ0PLx4b7FNVH9499jTlKcD+pEWRflatvG0s9z8890B
2FJfSO5qmvXqax9DZw2tz9p2iGPZNj/TisgRABrN48rluiaSaGcE1R27j4r55vyp
lIvQVLkM4NqZd3tByGeXy8AAZz0UXwXPNNnQtbDYPUgHce+baxbe6UViuVWegN3P
QkbQmziM+I2hX0SDCkobzdUjtfXl0/qux8YC+LBvGLf8i5HTgBv88i2ZEhSGAkSy
XJXijMqHxrExQnjpZERV9yzOh/oaYb79Xc6Vqz9LR5R+eZ4W4OpIcEJkEmeZkqdL
xmKTQTzFOlEata4y49E28YgfANPJclTCP0pLiJTXILhO+ykCWSb+GLAUDnKAo/9y
03uJ8mKhzZKQpF/JvgTqKJUjpMGY5Ze9BkAgxMk79Uqe2yvfOxEUyq0WXTdXJw5I
y+CcewL/9GP+W3VHiMDqHtYNw/hdi85WkbpT95Zp1C7uVMpofS/HCBBef3WmduxC
QvgTLZhwnKX/rgL11vebddt6OvHi2FPLNVfPZZY/B5r1lS/ICO6oOJPPbiJMWVYo
3QFbIYolJRFKcJ/S7/qzeg0UdDWCuaVpFOc5x9r/ujY7KSKUkGDNAV3upEOWoNoA
QSbyvZVlgOSTHN/a6j5eIO23WFB9QQQGsKVrbZrIRmy1wyOh9iFM6LkCONvZcymU
KhSxMT9tVF+f7Bwwtvoq6NX/UMSx+MGu/EqJb49XlNJJUM95UR32wru20feJjfMI
PuapRYsusw4DyCZtocJacIbyjYn47wicwHNR7Gsc3AusRguekxxQQfUtx/07ICpM
DZ3whfzo8u0fcNMQAs5yedAQdTn02gk4IVC+SUqqdFrtyzYF+ZAQ/4Ognhv7MyUk
pzd6lDfnNZqdkUXbjw/KAVFxNXlYmN1B4n/RHcbrBQDExZQLfQrrYM2WqJzpA6m0
4iWCx0xDpywBDFnkDR4FLdd4hzHiOGgZhcAfaOJH4ekqeMyZ310iT3YJwwINMS3a
6bgO9+BCPJDedXDR7YjgUrribSLDD/x+um33evVf9dQAvKcDSm8IHrZMBYnoIHO3
To05gn5McdY+j79Y06Tf0EPMo0HQFSIOjTR22PbkvfDziSC5blKafEjIW4/Ek7ey
+Rh35+YI3/+SgQI5jI2pS7ew+n7+TNwIO8uG7jD+zKcb4lVOUChghKvTOLk+xlhf
yWOJND5iERD9bhOodNNjKvm5eVaUhML8vteVuWM3WEE3Nx4s1/Y4vj2MTdNNBkbd
V6bi0iFqOmT6Yok5SBJmfwwmtkrONRgdkVwHC8krcedCiaIosZrYtOeWYhq4PsAU
jo/fPuf+TxwC/1dYlmUM+0kkh4s1oIUkx0C5i2LJodxoozMYSfLHhHrxVcifH/dY
XFZb60GIYOlz0x0YpTeeTVBwpzeo5zQSM+ovBMyLbecXmkgfI1mnK2N1caHcl5Wc
XdBxAvUDg5PCDulERQWDCCdkNV6RMLW4oPjNDnYWvdAWHI6ccT8C4nGtF2YfJ5Ta
PXiJMZLvyE2/I/zC+x4pXJJSeHiR5dqFopdtfP74tCJX+sQ4ZAK1JQ7RcUVTE1wL
MvQ1ausHlGHkADwU1R2hWU9+ybligzLNH3c7GGpK9tkdnbMso/u7bBwbeAZAnzSN
oax6TbHNeJi5adNWnAhUzIQxuskEsLvOlvFaDcSRcR/xZ7bkmBzlk6IG4MFU0HKH
uVaOTgTyQlmg5XRCXGUQ31fXAJVubH6Enp1h8a1MfGQ2bcjES5rZPgfGZba+xZQW
cEyS9086NrlNox+L2baEO/SulsrJ+MrvxXq5b7HJ83GYSXhCxXf21Y1xJpFt1VRi
g6K4ShZyGV+KDtBd/lB1BR1AHWXqFwe/F/EsQyEPAM+CotAhaS/F1yKJN2F9myOC
jTS3nDzFM1ByFK3TsycWBW6rMpFF64RlvOraPdewlFmh9IYfHu4l13AaArEfcijJ
c6YM5SiPTl504U++SZ90hmkc/gCo4GOfc4+AAW4FokPVgAA1ECjzVDFttec5aM/M
hlVFtqBL8ySs4QyiE94zcf+6j314rS6mMZgARbkcEGuVbaFK1WbYtVys/Are0oB5
AIfKox1QGwzrJtIuN1z5hupNPkB59JV4P/re3tJUui7w2t2SQRGKG59ECkOak0Fe
HAjRg2pPZQJIwEOsnBjIMjPV3Rqxvk47izOEbk6H4DFwRofaEzGYSTzW5eKDkaDx
FFbY85eYCUdWqx/a4Vruj9qLNeA8ovY7Lf94WeMOPKRSfpQrbViEZQw7VOmVT7ki
YtL7XYGx2FeHBXKJH1pkoKE+qzPj/YOauYRROHE6IbDXdCQaOBy7dRnawOpYdeEf
Q+G5ZpRUBCvcykv4rlSJRWoHMdmewu7ORG0k6hxa8VchJyT0GbStdDGiEOH4YciZ
vDdFr3M5pFlvhD780ds7INhVM0Y/Z+vM67CJrYvyyBCZB9XNJgpDqZEJQEpL88zF
KHPiU06I8VlCpDxrnqrEmOjp0qK7rIM3PXG/UT5lSEIBKBgIoH71kgsYFCqRiF58
j828/KK5JwpuOB9bv8Mj0dgkwV55vCREW66pgNZ2aJ6B/rhBbgUPtD1C6K3PJa1s
FXfXnqsjsS+dw7RIhyatUTLZd1z5PjNXIZSl67VS7ZKkLqUkNKaA5CmdG4JX+bbr
4DgfwaOUVCJftAV0n867s5AXdEZWwNAxnexvgSYZ22asmV+Hq0i9BHmhh+xV4Jn5
Dhvmls33Uk2F9q/otbNH8FvcmS9UadoKzoWfoUAjMPYFqFQcIC4PXZiehNSKa/D5
2VgHeuRL92n2QRJ8v+BnDSCjqqkaYdYpU3N4dCP/ubhYax/j/EzazD7gC1oMcMwX
Uh5ldT49pXelN+aI/4M4S5N+LqEk0cQa/tCUXdwFZxB2UPp+AiysoEebltFx8/OE
JF+UEpq58OkGD/Gs8LrgC7WKBfukvgg/JgUzLftLV0RanoImbPQysUZABKmYBOpx
ZGtFanuxvMEXscei9488YZKC+4qCnxztRKK8/cI3D0A5AMGKxxOAP0G6aIa17rQS
tHHyp/6YG51uArmLegdMlGZul9tgB0cHDKRgZe3/HWbFpdkWE+BCRpsIhX0W6T26
1hvQuxuvtp9m5IwqbBe2OEFLs/nh4NX3Ra4/gCJv9ThBP0+/AILXqXl5iO1GWNEi
Fjd8eaMRNGbSzAmoiQJ+FMPHi5UXlJ/qCyAA2AERqj7vuPoD1d6HLsop7qb3yySR
syv2cyFFRRG+PRv7asOoxB8wJGNs1X7b4HkwyvQEjeTtUrcQ3ZZoAT2JS+sFVnIz
WS89DRsXEerkS2ONDsgBCNfIm0bbuSauEL3AZZv9sg2+mmGEZPqdFzAaja9BPF2x
2tBy5KCdjGvMg7wxKCHsxKX8X57/jRYOt2G59OpaudsmadWn+Gp7sS+QVxAmO9h+
BoIoi4y36U/bl8T0qyFDcYnEoVrPcdtj5rpY0ADpRQGbvCmiWb5FC7ETpSbU0p7I
T4VMa2iYz4Wws+7iXvdoxRPWb1SnflMeY78mb4vgkjwE8FAQ7bK2KUK04NP13U2T
gZURwSrn33kBRZospDValCLxbtd0SGq6y54mi2JbE9y3gqjUuiZWCy5Fxyj9+O7T
Q+7w9Ofilv81BsVfORtp+WfvzNXBf1uSb3rO+rIQLH4/7EZyi/jVAbcJUVkZQgkk
T76QmCBhyqAGy3ho/GRvnlZZe4XfZcmpKhn1EJnrUBsOuWcvMLgnhK/rqToi+x6X
JXlyW0VSLy9jzaj8+j5jHFrXlZWOKEWEiFk3BGa6ua/R67m2KTjeK1eEJg1+PN7t
A2WAagt3yMOQoqxV+sI7kLkaJ0JYdPle2ALazp0v4FJHtifFfRhTg3zE5rEAFHo0
woTxk7VrKdW4yE18GakFxXxB5uFNM1nmRl8EQkfZA25f1qvbGJHBzCa1Ox32NAl6
tn3k3SjRomOmKZgS4FN+8NMgp4DUkGU7lowRDlC/sYs33lqHrN71yntMfiw6W1yu
S9ArQWKOGyCJscNnWvzXzDRcrswN1OZtZYOTB1c4sROhA1qvhLuXo6hoN3AvrLDs
bluxzg8pWzl/N8oLK9USfdCzbQjIvpZgTZour6zLoQnHQDeBpWfgyV4EO7BTggWT
dtQ2dHimXc/qTn0wa1rZ7894CIQTxc9qfeCtGRdDyqJSiawNE7mgvMjaD10VQQJk
B8Qjb24c0/jY3tMUa23WEAzMYZkC2Eo3AVr5YkMAb4yyg2aJdA7pkkmyarujDfex
wyvGuIgyqemzed4mIv4ZEGqC+Mq9zds5IM7JGm/9k6OWjrFr/SBjLfAKG+X4k7oi
hmJjl+kzbzgKj9SFvI34CyWORhK9skGrT+KjUOOoP+nGWEKLb+KQrGQPvDCy5Ld4
Mt2YPkhAni0E30Dx0+N2YzpK1Tswug3a3WLyu1cUi6PsQBf3HcXuBKHUQGnbievE
12I8FSk4T77sfe/y33bmwYSV8lgEN/PnHaLDZoTPsxwjhFoIGLb9UWAnerYam1pc
8LFfikoz28T7ad3ZJ1+7VDX5Q48w0QXenIxgKt/n6sHCiRN+ZFChjhO99TTFR7aK
1AcO6ypGqtyAZMZbcXrflahP52tLLuAi78pyNZ3dIr3OT3wz60GzOUURt1S5kVC7
lHpKP7lrRXeROH48eswyzNtkPN0y+Ir9Hmrancprv0L6c9H07mgmITuj9npvz8ot
l8CveHSnVRAWQgw/erzpcRaNITJUG1GgeLSlviw4jHnEKrkGst49B5ksoR7mFqUS
43YaIjG7WpbvQOT35RmrPau/QcI9i60qWFngYDQiaPejpB093GrofynVQIs+dPv9
ePpeufY7sBdp8UkCO0pzJFZbBxY30s205T3p6hz5I9PgmOqiLhuPj8QMn0HU7i53
GDSGKmSmlAzwO/9alNUpnDvhiy1VPaj33itj2gZRHv2oHs0+WpO3/6ZGS17d+hMa
mzBDMfLpAMdfRbuFGmcs7dwVWCDr+J8DHmdxx5lDHh0=
`protect END_PROTECTED
