`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PIavs4bh7P/A6LMxvt+Lw5QBkSC61yzmaSn0sHfelAf5oKEA+psZyKts0bfOKyMM
vljYwokSzIhCV6B/HUqms9g1GQW2lNY0nrhtM3kdebC8oLf3+/oVNTeMSnOPeZFm
jXtNKxJiMv5sIFl2TIXtDBGpkzDrJe0MmYtp1O4biPNsPBrjNH/GmEoa0fdsahrz
fyX3tUbvp9vVQ75cKQYkhP80zmaeoAYVuhJZTCSk7BAd22Z3oAVigtBzUIVogvlq
wvpNKgg6Pbzo+Jf+0CwtgUKVJrYzIetv3amla4bY+RpZ3hrZ1PSlDnJ73676VTOp
IRHoooofVBWzkOlufZv6HnwM6VF2K5YGkaeB1zkQX9MOxDI2KbK7WlqJNF5qgmSK
l+Zpdi6YR+zkyMcVwz8bLsjdk0TfNRB0kybHN6gaKMmY2OuF0qhbv99ef457z58Z
oPk5CHpBCmE0XHCB+FtaN2TbyEO6SrEOhuK+z4hlXvnr0IWHxlPEi8MjoerR8vKk
TOgsc2j3g0kUN+rmfZkDC3Kn5AW/QdnrAHUy7BEfVM5Lx++NLKfB1e3MRxDcoNoD
qIL7QO6RJTw2QW483NNHRXWifZV3Vita5TFAu4M55ZbxvifKVpnamA85QwbqdrfT
pb/RZAf2TYJ3x3TltISSbOTtnGL/05TnpsEqEsNjSYN8/dRvET3kl43Hy0CUym3A
yzlyuKeHXxkH/onZhr5+nORKbFoAwc8EhdDZxGHnEHQ=
`protect END_PROTECTED
