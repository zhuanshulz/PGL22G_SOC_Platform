`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rLvBj8dd5gZePoK9Ci9c/GNmMuo5lFi4nxgYFv9NoR4aTOEfrqAsKRFlh29O6Jzo
+WqFG8c3E4hKUeyCZdU00MEbZQEhK38zzta1QGjvzRdy9VjeWg/2V27Hk6dQP6ox
aW/pyLNDXC/WsG/4MuMMWHo6JXBe1V6UoqcUySt1FKC+kqCU3J1sYNuR426flUJI
KQvfAhfuqYmPgHUW5F2R3cXFeFvMpiMhnDjdUdgYbCyEwBYQWQ2hb6BSCz2UuzZN
sMHnbkP9acrp93GclPsftPVn91TPijula61Yiyf2bT93+LIUeVCKGZTiOj61BQpy
YQSas7rheDbutBWEwY+IRDFRKpkXObOHrRCcodpm6arfJtPAikQVq15tn3DaSGWp
EAld1bxvcV52Ea9w+sP+yYYkFum/x2AhZvojFwv2CB78zokvb77u/xRMHT7nsQFY
Rrl/S5NpXROztmwEXT/iQJAkf5YUmMCsdDMRdhIV5v4IJl0KXsECLZlar6JSxCQo
XKXqzvd5i74Fwb9wZOeB8wIINh7ziqbB5Yv+v7N/pjfwJJnEvHRH9ZBRxjQ7PYG8
Sqp/gJs3pCvyBPyODt19DDWku7QVUGeX1OkvadrXZzya73N+Rk+D6ACwfF56jbcD
CG6f4oU3BrLNwBHRIdrHffapQKD8XycVKP5/y3LUrqSealKKPG7I+bDpO0j4f9Dd
gIDcBm0JcPvIZHv97Lny+tp4o8w+2oouexiJ5nY/bCU7fL/iNEhlvLsspy/aUCNo
ocbOq7YzDnBgb2aKrQO1EwIAA/oYQQrI/wnvOIvoQdI=
`protect END_PROTECTED
