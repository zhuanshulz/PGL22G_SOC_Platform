`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XrypzpxaiJ8b561AJYGhArzwcXpxZRuwHaS4/Te+VJSr++RnjIzhfjZb9zVdEV6N
pxYz0UY77fJ+XPjCB70JS26wApcdSce31Q4R8OYeoGlnkOyaaSxmEkAEnMMNqMht
ejpw3+qvKn6vJz/oBx5hS/46Cbe4VAg9h9zhd0SVZP8+liB+BGPI4OTaDfDHRbT2
qgYnuzAbFyaFZoRD0nwns77z9uSmfqp+MCVK0mCG38NdD7Fm3IGL+4PUsXZEiERu
qkVGNo94KwNtr0ndyS4aRvpebFnssBVHeBGQfdaeYPFADvn6/uAixOvWJ8tBZ6FR
gAFBD9WcdYXeGmsHR6uwRyI0x6/4D0xdYZoOr+DyxHWpr7KlUgMT762uitWir36C
Kh4S8lDkQVmHyvykZoW83d56JT4qUBkZQz4t1Qve6xyOyvHTfNIfmgN8Wn4224jS
TsoxM9TbGbtl49tjGc7H+o+5Rn6u1DryNUgqBJkn4Q24fKOAj0TPsOeW5PVcBH/G
UB8VTQ9JcXoe4EDsIquoEs4Lh7lf41o//DdHQ0U3tT43y8QVo5Wga4ZbEzCest3a
36VHjnD6norDj0EFDhmLfsPuLLMHOEM4JGmaNpIJ7REBFiftK48exHF2tvvpep5I
2zdW67J7im4yqu5znpzlMRD1MGyQrHczpAL9LPeh7A1OJaChCZgk9+vy7Fj1Ul4y
x95yt1lGOcp9hW+G26BpupXCEmuqniSp72xhVHiFp71ZbbuydHbFwBzjRoXw1zy8
wC+1jvxAltIzyLf2AG+niGN4KVKrdnnHbEZ60VtjYIsYXsIoUY2Yk9ky4UVGCrQu
4fcUZchQbgup3UH6BnbhXBYi9DtEc7woUzME0JHtGM2tLcySpfnF1CEJGrAvmXl1
RI4vhYCMjD4nxroQ/WtwyR64vUNLr1XL8BvHVCMcIrZusjg0AmivkuK5nDSNae7p
/wbyTSqVdMpaH1MIVAMpqrRmWo95Jar3nj9pmc4RbUAMzm/wROEkQdJ9QHPEzxD9
5gqBX0cRpihdeS6Hejja07CxXQa7ur7wAHhMKbFqxIlppo8Z2q51Jis1c9gUSvcR
It6DjDlulRWEhnUO3+Moej0jU37xL5og8jn3LFMgxtynVPY0YLw4pH9szRwRnyRX
Go2uQWZbVyvXeSw6bdvjTJ4Mk21G4Rra6Z1Oe7DcNk1udWRCcAXWsj92HeMjwiin
SOODPj6cJuRdyg+Fx1PU9uWnO41NTPBlBbt/EAUkYnz++7GyavZpMZC5wW/PHC87
IR5Qm6RGgawf+gDuKnn4T+rPJt7H4HwsP5ulYT+qpUXy6cevm6RENcJ7lX9bLNhi
epifTuACICs1bp2wTK5ykciDIrIpl/QufmeM+8QrXz1VwYpa0liKwR06LrjOiwYj
/Dlx+APLbf/lc8NJHyO+CO3aBNd3ndq3GOnMDqgD2Mv3MVHpLbpYpwa274nZs/f6
hno1DQpg1fSZFtA7IZsudrtIS9OvS8mgs1rcVfQEorsR3jTLxTH1MXYDDHHi8TAZ
enyb+Qm2/qzLJ24BCHJDwmub8bGfPoMC/1U7cQOQXfR8JTJpygvZFnQyVB5oEIhp
FF1HPfM0r/CgBd6O+85f963wSq327nHL+hQvZbUzbkD1irL2//ip2S1XGsnDSwBd
7bYs+GblOIIdphgffTvRVuoSPKQYPFYammnZpCUdn+o35Hx+D7PX8QFOYHfIa+VR
I43EpxI8mT57dnNcdYUTsBRr5pymhCaJEWibrj5iTeNMeb2XPAyJmHbLPtQuGHpo
VC8kG0Qok8GlPZWITfXwXemGrdxrQLEOmmoCjfuhvyowVpAfDGmkIpGYSLUsNSIF
nKu1t3g1uzTkPMoPCjVDfAEeUtG7fOq2Du7Qq+88scxctaNDBz9hZobwSnFOAfnS
1NDpjnXK7ym+j7+w8nWhfXND7xSwUAnPX6K6KuP5dnL5MBkW8kkyKLS2e0Lvpplo
LeJEY0AcptSQ72uyG8k1ozUqFx6hfAzh5eySaflPV4Pz65WGCYWlUiT+OkB3eSYJ
WiNlgckzfA/YK3qUvynoKbb66yTCNGn8vEBTtHWIE8iY4b89Qq0J10ExgEI5BQy3
nymiiUWcs/BZQe3NDwNxi1PL+DpYDDRIzaunVfdkrTZgHCeBqCHIv8AshettILf5
WjJwuOkWksgaVttrg1W7RiJhuMSxVqVWdhoJML2D8X+zY0lgKLnolXwu8z01UKSd
Tb7K1co4O46BFfA9haPxMsQJ7aHKenFo4TICM9oxuPbCyUHvNFzb13HZG5UrdY7J
NoAf5VIOgJ1D8ybhE0NpS8x10l1VjmUgkanPgm9t5nBFg59y159d8jdQE9XUxe+j
B1tKGL1kkFrWd8lPcDLqqp36eI01YPByicJXlH+y2TxA5zXcRmlhry5Bliw9i+++
z5oLSnpxdIXBXjX8kg+fQNj1p5lLa+SWG1zrqXHYO5OlVJpVu4RveIlgK38+5rBj
/bdDyDgcCTSPQT9KGIR4QD89Ltn1vJ2E3COGw7nK7tzWyaRb1+Eewl7t0L2vd9I7
g8DbKKgQ1uxYlpwgy3VWc4veB6MVcN+lFuxdJAH1/suL9Kf2DZdp02KUqz9o2E/k
RYYbrTigUyWVY1bCIFpgggYtn+M9/2Ll2zEVewN08xgYh3KazvaK8/gTEhImNMUF
w1Ud4VbxIMN3wyHgGYapazZ42w0YYQ6ivwZehB3uiwq5pb5Sz/pQ0iZzJsn3zGR0
4Kc6RBx0yAKQC64yNsE9VZFDIDX4lqMbg7stzy2bAnp/GP7ExH+ELsUxqeI3r3LS
ZlXmdN0ZcJ6uqNOTVawPvtN8NRJdybQkmYyzuWzfV/8cwu+FZYGDKWmsT5ydrb88
HWlFcF/uX1G4t2S9fSTHDh/fPX4ZNf8tKi06dKyYhlk=
`protect END_PROTECTED
