`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8vsXQOpTbCx59s9wJ1WzNzKCu2epKKOOnAC5y2eGYena5XjAxYMLo7zyOO0q8tXW
EwDGuEh038w9DSiV/aiirqCUoPY//xtB1aQhQYfluhUwRs8QJE5jM132KWEB9F25
6x+jkRE4JOdL5My+4umxFRWkM+eTRBT6rZJuOVHGrZX4SqN+Y93X7cuu1MgQvPO4
eWIySrJf1Bjm31304bF6JSYHLy6yITLIIEwvydbiSSpKYtdEAuIplkQS64MpGh8k
vWGiSOqkJ+zd+CLTeHSJAtOd6cU1rYSXada5gR7D5zd9UaDzWOTS0S1vC8SdpsTC
vCYD6W9hnNkf34Q5Laj9E1/i+ckytMM/tN3jjdIRyWOMr1nxhY1iHhX8Xsqi9TM3
UlJS/svvwr9eMIyif5UZjld7Bg08tnKPizmCQ2bvRGWgCBWPTDyVryz1QyFqG0Rq
d26NQ3JSqsqhZm9K4mT/CQ==
`protect END_PROTECTED
