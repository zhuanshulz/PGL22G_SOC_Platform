`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kAmjqw7eQyipuyoZg+NqHnZ8R3Ifmo7+1O2VGRdm5slOl4JbWscDs2gn11lKvdd/
j8rfuVvRhzk5wnGsLGnqhS9NHjDc2ftuhKoIEFu6sfJ9EoPEZz9YsR9xwIW2Wepk
s5EVJvdRZmcwjv8B9BbiJgek7cJJaUCMjUErLSyqOgD1JzJX2Udm9XHKCXGZ88SI
U7NG5UdCzVsvOs/cF5knrk/1pitvgAQPhcBENQTrAcYH+BFfVLd4uSn8Wkw4w5Z+
Z4dFhv2oVSb+545lPCwrStMh7xa7fxPlxjDegtqhZT9bopvoBf38KAGOE44TDDHQ
GlwOQA0E9EWfKwTpELq0o1qBzFzAo8heFch8Otfz/vpbViQBupLVitRqHkh74TWB
wg7BJSTUWpjuRt9H5slSt7tSRXDlQytqdz51MZVtGLN+zI8fymcZLYdouR4JxlLe
0ND6XggvzVImOxMcPN1009yhF661y8h/3iMWTVj3+Ms=
`protect END_PROTECTED
