`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zHWz9liTbqaOus+RrXKmkcc9C2i3PvwqiiQIpJoqPq4hIbaRyULpPpAcdsll8C9U
Iyf1eRx7lJdPZCuhyHLOC/cWBBo7gfVwAtHBOmXFCffWMM+Ns6LdhsbkXJrnEgos
FXfNLWmo+2ulyD6f/rf0u1UR2VUbhHzd1ODdD+fr2kzxyWQWCvobeed2OgKDWE2x
FZeWmueh+sqG7LFs8EANy+vmoXQWGdtJvTfrFBsCgIrBlEGljrOv03oHr4Sp/djM
xXTLMVq1fUlJ+Q9LOoF6W3ctxTNOEQ+t42MSsdJuBkbF8gKJnds69lVjtk6+aA1T
5f4JdqINQpvJULmY0z1ck6+7os5YQVj98K/f+4DdI7I/wrpEff84Nl14sa1IJHWa
9NVOl53vnMegJpMUR63WkaNcdLgYUD0p5UN0CWR3VV6XH9z7HyLsE/EddVxfImYO
pKledIcOcliJv8hxCbcTtmp5HDg/YVBLgKpk+DAr8OkG//YpOGP9c+Ls+mx4YIJ0
3frcr4MjsuKYVnPp6jToM0jvRkYoytjhSBXC1/yvct1GwdozoAfSCpUFN2MkdrC6
wuHly2FXvIVwPxc738lBQRQHmXui6Mw8eMbg3NAnPG0T+HEtUtRp01z56dxUsvED
3Q4znyx6yQZY5JChwiRkiklZ0eOZeeP1O1av/MY6HND38ko6fdNwj2MRO53TRe9f
XB0oDn9kb3eaFBRScrgoRmqzmzd2vi3GSM2H/Vro87EAs2XJfScEIxjixWPCm0zG
czItjgvLr/yxxgEiXK1O+W/iqf/qhw7e++2Y6Wkl875eHzrfxgdUhvlntjUz1gAj
XLDaxEVN0Yxy6hMqsnYNvexV5HNlGUUno121HYcIOl/9jjF8/Owr3bhIQiPFyGM1
pw9xGS5KNiCbor3YqNnZrZsG+rONHCT6ZEyn3gIhMbotMhcmcWrYk9FVo3vm9zLh
0qTDDmom+o6zeKebIQvPU19/AHXPX9h8gsEz0dJ2UgwDG3r+FD9KsSqMS7STv4p3
CegK3Kke37vram0cW6U3HZX4yOwxkQp8lNWY+G4UCFyk5ay5+YlCxMnTIQbu6KZo
TD17UPnKjOs7yz5tbDKfeZKYbKODQk0taHgozYfvHYJ/AtOMCDhj4nJQUcBZXLtr
eQhxBgFu+4EwcxTrr8nPPRLH/CIcjhL5qvWH+Vb6JGh8dNUJ3rR4doZLIKUjmHq3
gcIpkUIycYVD//EII0szlCiA33WWE9eGXslHNADAZH8o3rWl6kGxXutLcG12gb9r
sQ4mXSSvEgaGKq1RvjcZE/oJLaCq9e7xCzQeYPdAvwQrklBHdzNxsZCl7S0BxaKB
29NOT3lBV+EjGa4pR88pifkTTG7+3SHCfzC/3PT9ooaKpmA3S3PTL2w/9asWwRDq
EfV6pIP270P+QYpeypuRr7m6MqcqjWaz6aE7yUamu161MgVSYv8Ec/z+OY1T1ioe
lfPBP3TTFmFezJiVpzZicrLYN7dWrW5DRsf0YqnKVlWQuP0iJFUGCEEL1R4baLq/
o7bDAnbVEUWKjwf8HZDkYvx+rn+ffPNQoVwrm8RT6t6jPVdU9fCUiAXB+H3ENp+T
HLzNAyG/NchLoOthgK5WDdwu6DWl90NXBLQ1KP4d1YgUELvYuefesKoA3UChaD4M
iMfSYDWUyBwAJTGqq5EXqBXajxxkcRMpUuWivjIWtQ+Gzdb/pN8BPlvHD/cBuNYD
2tgGgcNiGg+QnOj0eEYBz7cdDO8ET7fo6MbLVhvMysVBf/D7Bw34WX9AOdx/IWxx
Fe/2ccZVWApto+7FjEK+mX+UMaw94ahNiuwlNz6zkLAWr9voJhKognV2YweSdbEa
b6tiwIqDgy6xEv3IqR2yE6eCPXJCYSwjvpXO7CYtxpm9dyDKwUIxrWnyIh5I/dH8
+hyvRr5kwJ8xNFklkW00kUkONb6OP9yafFWnjoO9vqX3311a7HbT9gJ0YO7msvk3
XRWhA7IYKG/HtREd5SUSiXalTYexjWux3p/FA0phLNaalL90u3imyo5OCLvVM/Mv
HB6P/qFWHQfgmGHbW8xPRn5XPkB4xFPYPXCL+4fB8v69TTsX6dY3UshmZlQWy/Rg
2JZr8d4fdvVRHf068s0M6uRKZ9ZAD7AlZnPXOEAM64XJ0PxPV0+DQCnDfsFh3clQ
1rtTTun6XJOzF0PpZg3BTa9wuc5Eod7G2ha1ATVGkovtFn34os4av+epLmjrL2HN
Othrs+5cB1mj96+Ffr9VcSPSF5vs36kCBXdfoTlLImUa9pTu5eUnnEKML7yf2Yrv
vNH93YGfpQ47vXXAmkjcIOsdVz5oeLwZ2McHluU0uCz934Rikaz02v4c9Z1W1yHf
kot/EnuPA7uaxAledvfdRCHpPINO9UJgt2QTuz5PoNXVYmm/DrTBMkaFSQMO45Zx
z5gO4IhXtCT+dlqmQsjdRp/UPieQyR/mYSAHEwF/EbPI1ob1BUR8qHlTTP+rKMCt
EMadNxEnJj/t0Z3N9ZehOYHvWX5MGlrkIY4WK83j6aTAnSFefXsLwqWI/4Kd2VZA
DywKRZfHCYmQekIeori6EBPQK+cVV8tsMmW95UWohAC05X6pFDJ2R6Rk3uKz59ec
3qofl7au9ldn8VJaQeRIeTQsL/dO+yWc5q/8Dbh1SoCNgcsEWi588A4pNtf8KnGk
BjP+iy0QDcs50MO1izoadi0ja6HyK0DqC7LkCqQsciBrtqUETgxi+24224Dn+A4v
rOENyOnUOHUgTHTZmzcjHEXqjWl0yWiXHRmcJcs2vlTAc72Y/VbzlhNQEFhTnJ0n
lR8ItST795gyc0LljNstu2jUfP635lkPfcRgV6sqzmpjIhdmQ2FleJVMMMGtWtq0
uWbfiAhG4mD+xgUGWhYvoOj9JWZfSDRKDDvZGhCz3OBThD3RYMfJIXmm+pndyyGE
WRt1/DtJvyYgfWgrfnKcA7LlrAS5PeulFxj3Gwd6IDm6l0qJoRIBc7d/Uif/1wGX
A72YxDnUn3OLt+AzPPe3Y6y9e7GjilrnIqdkiORSSEkarb0uRF+ePwD8zBqiUr3h
sOraoa9fxUkmusnRtZolb+JXaeT6wiYH/nM3kvkl+WQnuh8Fl2NKAZf/U88v08yj
YegyY23yimQclYpz0hLhk0OtXDSf69JXrt/XlhE3X05vmuwAqLxINRPu/isDGKm7
DV7tl5qixl4bJ+fJvvhe0Zzc4LkX1uhuwAeuUe3S3Srnivt/8Xet8fOlUQYdkD4O
YBLRw4CZ3yJ8eijuDIcwd424P//PUvFAWagvQaPeXHFg6p9Xsl/TzOsIhMa4brRO
xzTKGOswiOyj5+PbT0eiu1UwPIrk/7HZed1gyjmzCUj+hWFvzvOwEYdbnnNnCu9Y
6QAbjWQiOan7Ri5TH9r/r3ncsBBleq8bpbnqdWH04pp/9WLxXyQSJprpJeBR+7CR
BPUgLLFjCp1plvlSeC3wvXkifM9wCBZAWoxo6mzh8H0n6FYr9sr0WAYVNlT2sDr2
qeGJAtv2iFCfTWyITSBWkl405enYgp088xaSbIEMnrcbxjAkCeopeZRAGFIKlPLE
5dRp5QRd5ntTfio4HdL7NNS275Jdbqd/3Cth/gybyKfPoGp/jE+fCuWD6bNOIHAp
AzUx7NK2AaillrIIAUhHqEcUhcytUG8ZBf3L+7zsnnXn7UnfzCWZjDuyYEdtBOK+
SFPRuLORPFGKi0U92pJGwFQvjtOiqMX1L+bB6w7z+yRa/C7p1hhfgSDzj8KMTQEM
0k0g6LiP7hpUfpTcy9TCKXPYGDzNjRBwd2Ay/Mq9aV0HABsgqIDH/Gce2ph55Z9M
hKvC73YgXjgj7k/llBIdE5fPf5/D5Knwuid7VHe/SL4xTGBQjzR5xnUbRnscR7tG
HDlWTnE7ZEfTw/fdiEulDrr9IQsAUK45IItDXC4EfG70nZxSICbhEirjJe18iHpg
WCRCYEYtLhUZ76ZabW/qLW5rArycCdKfa13RFr4uDxS+y59BLzKGKJftp5m5xjrc
OuRyOpjkyG+8OB68jvQkmZoZiYoXQm4YQhreyZMU/9nQciTUl+Qj3e0MtfJWmkYl
l7dXbna9bxA4iurWlKdQPTzdNOAYW/ZXVEO2oZyV/zMTDJQ8/Cxu2905NQG7NrGy
K/zs7W8Zi4HeYoMbiVC/KxZRQXWXHlQj4AIanIsBTRl6dEtYqWvoz8wqmGLsuyD9
6/hxCTUXKniKeuo1zIfsPv7pnDppOR2J7QnmSZ6E8OfBIoMsWT0QeXUSw+jxxwvx
9FozO6YC6JtykWuH+EF3bP5dLW/6f0yA4WfJFzKODqFpVJtQF6CdyH+9zTlB2j+2
godPsA3WFY4bePsa+lto61v0R2OdEGGh46bDWU6n0zV7KIT0UnNoo/TVW8mTkaA7
OiZsH2BfhgYmCmCbSI9Mz8nXqamXowgt1zTkiAlxiTJjpyq8nqPlBGhQ0gu4krYZ
aPMtU+Eg+2LluRPHVSuNw4fIdAhP4rbGMtTSC4EtAPMbl9mIH1RkKxFkt14ed1n9
Hk9PMQVw8yuJkJtZaDteS7DBm6gXTtmkmb17Xju5097FdszaF670iQHrXwIf9cdY
IpTKiv5MtBPC/JGdoSoV2q5b7YEApyIRdiiFcaGp50EqGp3UXBVmVqytSMt1dUKf
i44vupNRsL1vrU/mrXCKcCYSMn4zipMGVjfyCu4KXUOMe0aAT3Cl/P2yymA9rf9z
1nSTaB1JJHFEAINEvpQdJPD85veox9nKKjQM9tEKTgrKXQdj4I+aLPDRvzMgstEa
D4xxiUJMUfzYI/XOuB0pCkaSbpInb/m5Tx1ajHk6yR0f9COzuP2aG/nP81RRT6lo
x9joQpzjAu1Lo/P2S8bibpsMDSvoUkiH1ohKBCA+zdahnLXF2JRTGoOZOkVhdWcA
/OWkeX7Xkd758GS6cXTYlLkwWG9LuV5YfHZ0PzCuoyzvKy4H5BAwFq+DJns5GpmA
RGcETPdJ/aaggPXXlLSO+HrmHIKu0daGWMedpmbEIYtgB+85t7/ugbngPN3V1aqx
0oQLW6d29EGnUO79era4cskeP1WNJcur4rXRARDyusHQYaCMuvIxiUwN5Mpy5FR6
c1OO9stjXC9iZsVgzudZyW1b/9o1TEOkhVNDD3LiyEQoydZzF1a5eGJcAWPk8N+A
KMgN9k+8PK4S6wHgYg0FFT2uC2VPn+JtXq2IXscNPF2zbcmyxjNPc0gYwpiGhuxG
nF367adH3sMkIEzBuJE8U3nZBjYfIbvVcf6Qsjn5NAPquHIaOK/KKLmM3ew8dD8b
pvuTnaVEpUbFTs91lgreCPpUg0QlPcbTvOBrc5sgCDLTBA1OBbGwXOuboKxt1ER2
cKNDCHGbs/Y/FcDXpmvZYOapwrKRVddf+Q4wkN0XgbsRw4WHrZaE7KZRszq2/8xZ
NDPjwaEV4aaWzHRHwscda25jBAqvcLCKE9bPl/SDVpv8e/7+YIhMNAf3HAQi8s96
dq1ckTJmQdsSbOjvgD0eEHqL36V8jUw603q5GxY5+ZJOjQ2nAB8Zt0pOGkyeegvu
p9zzIJKB2YoJB5XaQCWF+s9KFRJmqCiaJWf4usvSF3VQnKxXmjJpgBKkZd/YxPUv
7toH9XeoQKE8JYh5p7yw2mnuYORxkNP3egUEGFan2RcBGFPfCQMSCF0yN6V9AxGJ
XoVQ37X69t7Ltgyr9zzHv+P0FeGuKsQfygO36g6lSw1WOOUOF6aoW48DhkBZ6uK5
oHW7wfu+fBUHRt/u8xu26GUBZ2YIljydCzupHPi80S/0hKB9K4PLCNcBomYfhg2F
e2cs5G1Vkl8AFnFWd8oOhBEFayQ6DJBvYR3a3fTcq+xPLAifNhBh+yePVqdtVx6D
RXgHKVrb1QA62QQ8uC3DU4nU6UqFJkofbHni3hgWnLk61VA+Oo7rxTQYSPVrexEa
IkB+aec0hQNofUH+LnoFB+zMTCh+s+VIbrLU23WyqCZqntLXtFg0vthvPputQKpW
XG01exstNd7O6jLnjwXfzqJ1yhDryYBqVqjA1Pl/gbXyYAQDUdMZv/098mgbvKBP
tGXE5KeDwVeKWsVV/uZwDBD0BzK8insRjlU7ZCP8MPgU6fDOG9S7mYzjM2r0mM3x
Qy8RExpR1nxUFB0riZxtavAJRRgHbZNkHq7P5C4Fkeq2iW00PQGKqCNrXfZga8En
mlUrcdmPHL5PArBtDpd/F3i/nXoeNBLeyWk2GVoFlzjNMh87DiVdLq99OXlHR+6E
WfWx5iLkBiDFt1JS5L1iv6XKn2KprH42ZZZINzo9p6qHankpuPLVpmlsWjDXdacM
WCntYyFfoJG/ZiHdsvAhJm2TDmom0G/i14fpivdZi+lwfNIcSnaqITLPaYyUMZB7
/yS5qloLI3aqAEd7B43GgGQXUzzU3jYVYgRAf0oTCduaanBY8jUMGNZTpvbTBHGx
aJwry/z5y5OiXVgt59AS7yLonVHt6imEUD4D6tPYabmlfsWlSz8shw7tGN9dVEg9
uVxTmCLNmvcW+/PdNdAni0bVwGs6h0D7rMf35Y/m9AcgHkBvZZVAEiVwqPPTRw/b
YdDmPHOzcLpz840qsk1a8Jg3P9Vuo66xJa3qjC2CUnZEzvYJHs2c4M9GJ7a/sk9f
cLsSPaOKsfCHOW2U1xo2nzkaj1Sg6R5Qk4UXGBqsODj+IUWWAgsqlFrOPYhPjJW+
RSUcZQco+YPliVSNu1+T2cIHQR6qBb2UrRTW495TnIeOxN8A5pJaHPCH14dQE11E
UYy45P1r6GBDtRPTv3RyLBoHOmfJsSApWwStMgMUZkDTKrXQQ70czPIhqqsa7twQ
i1PDitqtd1nzZRD4gS/TviOKHFKvbIoB+ZJwxAFyQiKFinQxdNteFWLTfO3eOmq0
TqSJUsDYhITAJ5Pnf3JKq6m5tJHlz/pYmrdlsDs2SK/eCWFW6S4y/g+S5H3XYJjS
ga2kkdrHNqYZ4ixJ+nKa+HoGJQS0uYOrEYgFPAR8ugDi6xu/ig+ARDts2Di6phYa
lB1TAAoGfkqUx8vMBFWw4iqo73DqjK1H5nhQat/JKH0ECSNAgzgY4VuEgGZ/ldB7
C1W9jF1g17xODvfWIqFwD9lyOuN66q/Os7y664/JlXBbPDwd2o9D9a+0o9RF/a1M
U0QduY802bq5QSwlMlvCXnQCoiG92ersFtwEDW4gTaUuNk/nRTv2jbKio2WFUbG9
xsggdY6tSkZt7Zex6cEN6wA4PnutoyHEvVyD19fNOcVtauCg/6c72qBVsdOYYxrD
CTe+RNGwVqsBunbeSABaIdXFXFT67PMXo7tsD9jxCWT46PNLX47+pOV7bjE0Xktk
KYWvfnLFMAwx6PcZcpZS3B9drxaHLHfHwUc5j2WDiJwMkg7cxf28B61eOt5mf8J2
9OEUxrR2hkmmZNH5HO3NrDE3qqeuJk+TJ7fk/HClewrB2VhwzQZ2n9QvUKTBEoDI
xWkzAV2xPRbrHonCHFyWuLzD4DueyP29j7vTIii0/GN9j1Z6P6OGt4xInJAjJOl+
H3drXhRLvbmpRwErNub7pJEGG3jBxGyg3RDghuGibroI7SAEXQCw5e5tVkbMajtD
G7Smfdv+Q0Si6tQdBiXDz35Hv1pN0LHlfx6PBy4OmVHns4c3GGNa0r7XDd5EyWfy
rCUfP7Kv1XovEg2VWjfx78lJ5oQ1RbdJ1APUKzIbufOJMec7dAfxECZlMWbWy+f5
U2m10lh8yu4CytJY6dq7w/gpHhdsDjegNN03QhkkGPBkcWEtC7czrAfhQyOk9yEL
UH3FqG4B1ffYHQu6I0lt0vesmLTh2OWHb2L1aDjQA9gK5M/CHxwsceynAPDu1GlI
RmBYtiTkQJXLP90vTtfjXNVJoWFvCmXL7pQctKmTW1BkGbOqeLb+u+P+cissCXUh
PJRDSIxszlmUUbz1uYXIXKaI+/icdXsUbKBvDwsYNQKO5tDZROoUeO7h+BDkJt4R
z30V7MSPdOw1MfsMX/+rSWKMvh3zfuqbOPhccE1xeq2Y4MKS6luCCy99luZI9Vs9
+U9th84oSjVPyCPnI9kh+rix/l5bo4Gt09WA/NJvJ2zQj/k0Cbrtm8xYUjEC1Zgp
7kvg1xN8Hr27/QrqoGURrkyNkjfFvWzfqPG+cy+8RQz80/UBdFMvzRWo4i8t6esp
T0qcjZDuL7UqiPg8UOn6X9tDpjwebF9Oky/naCflWLzV2eaFtVTlm14CU8Tg2d2+
ftcQUffoWNRGqxER4p2Y9u9UJafzTPPtkPGrOpRpvQX7zua6/BMAOktoqluCnJSL
QPvWDfDUPO2QE/vBAjn2fA8hzw++Y3pJPHaCI/Sd3e1ZPaprGduQHZADMvqP5WFR
FcHURMQhUkmkCCSCJlTFjaAvd9huY4EMy1ztCOoH4ODpNCwg/LujWKY5cGlc+qoZ
b1vWE71Q3ca/KNnECR2nuhOENlM+DjTVKvpAN/N1JBAkG64N/B0uYQTHuKQs7xtx
YFYUmuRN2dDpo1iJfZ3V4yGP8laOSAOSVA2rT/AoVpuN4jUzLYsX7OzvuLgG3Mv4
IZEFIH0kOJ3tggxPB5ybVvuEScEODrpzX6XoGFAOipiRrIToKVQRg5x5yF6BhjVX
NmwOfWksbJKxhP6dSw+jBRaNSSwMl7ikatO5uPvzRt416ymUnVvlMw/t4/Z0h9sw
CYabOTNMJEgkO2ztR3+NIIBbkd6KSy2clDvV8FUFS1Gi+G83N3Gcc57uprqcH0P7
YazUW5cBA7qzBdcYPjwn5XNyHjHCOo+nhOs3k7v1aQ96InRxB5FC9RTwclzuhJsh
C4/5Sx5MzJSNV+kLIdO/LOKZiDIXwnBCN1tv6YweXSP5ie9HL4EONcZrqFFUSM2F
deYBeeCv7erbRBJXc55Mzu7TpsbYB5oWPTx8InBtf0pzX8roGAc/9xIgt2rS5Vun
ER4ZUaF1s5p3/OZ4JfZ6e9OOPzX/L+W32I04cn+utJ4Pm8JRIQ93ixiaTv5m+1So
VuS+w7LYxHdL+LVT9fl57pKRK/3ORkR3yHyeew8QD3z3Y1Ki0am78fY7qWT5GYHL
AYqBC4CpKk6n6M/Hi6TyKVLvGXAB+r8BQQXKE1J91ur7T/NifqatS3gwpAmpZzPk
9WTJ10d/VYSxwmdl2h+n/OJmZE+XjhQd/YouAC313ZC7ri1kpzz4m9xWcOJkGnGT
08w8Gyj/EtOAWkN7diSqirbWa10xMy3OQmhJoGWeFEGtH7BKnYBDJDTkESowi/HR
n45WI2s7FoMv/sLzq/Ns4gUr/YR6TOM4od3pzYrdEi/F+I/0cs42XnhOMZf5bxMD
DSckB8RIkxnDThJveD6kgElvacwIraIM1f7tXo4Dzpq8hHJddTxfSaQQp6eHK39w
jZrnid3y2kGtDQMwaaY7Tgc+9nsBcG7T4zPLh2xhgrEVnDuA9M5kJmfxsNJbJcHA
gshHLCUoWEwHgJ2M628H6+6aWfBxuKXOSjw2fCTN4NL/5cYUroJZDZS3vARhp/Wu
qcr68M7S/nOJ/BnjzASqy45j8HC8llCHM+2G5k2eUMcDl/pnTbSx/UUC6qH5/SaE
U3GaOhaMFv6HnspBSIusrH09p8Qf6bV+R9cwTw1vrcuFv5vw85mmRSukadEgsnGq
WlTLX0pBOFGI4YFznoXSK7PWQpGw7AY/Fqo968LY6oocSJMWj9/WeudjGjlQComu
diNGZ+RWjXMkJvNnqhZGhOIz538ZCjrP3jUbxDp+uGsHICuf/DTfQiJHZf4Z4i0M
uWH5DiHsmYOjjIdgHqDHszxiULCYOiBP6Fvlvre7DvWL5iL6qgew1S+HIgo4X2MK
KWbT0d3eXMo/n8AoZqj0CbX6oKWxxIp4LLJmuvSBESRBcHfRuoEdQKGsCw91pToE
G2ewBQ8gCpiK0xdwgiKniZzO6hBdPkRYrt+l1uvOJPHqIV20Y9yKxCfB0OANIqwQ
iYqmH5pFbB3D7VjBXzrf3MREQCWtGCNq2sEnOMyBPEACPKTzGU4CUZEawNa8HCBw
Jpqyo1uewulJzgxFiLtQ2pCMwy5mS4wDpvVjRmNPN9POhr1y+Or8eOkFvt458mVa
cA9f6znu4mVQYkfvlVvWILeIPhOmtmCpmT+QmNt72siu5R2yg7diIxdSZJ4gofak
PhScYUN0UZ0yFsZtaYL572j/U+ADwmp0qJ0RaMek6rhwq5/EpxwMQJzookgF/+RE
oVbNWzDsY1LE+L9izByq1SPaXmqeaHnq4LzovI5BexmiGQjJ8IUDUIGWzoeHh1xZ
CpUvm5xztdGpvOyPBKcaPeZ5PBUkCijpvH++zCB2+wOQz1B5N7+BKgGdE+NGQrKl
uO/VB8DPCjxwlYF0fjewTolTUrFM2Ec4ZBI+IdgRqAxMrwW6ayO/oUx/bi3WQCXz
sRQmxPed7xJRHLENVL8Shmk4VMVSLAUnpLlz4bjd9GI8lckcixwxQtGGGo+RA4gQ
OJlpG+hVxcalTeUkSusBkHz+zPhmASwauvHz2Ej9utpl8so2+7flofGxfJbcFWvw
bMgdi1pexqt5IupNqO5LWBXc3Bxcmjil2wHnNhDuRBMC2HT0RRE3A502qFG4lb4+
m5QIrT6O3B5f1+uOPO3D5HuWMu1MSYzhdgqWXGhn1uj3SySc41TDKTmX/ymSdh1U
NCJKPCwDs8vgGKr/Yah+6yDHudATdFRlwvYRMZ0zu3BDlTKaFvqHJP1ojEwry5Lq
X03YPtO7be02xci6DvAT0P5HdRDptAlvT81NsLnr1KllDvmTYDF0SMYsZ+z86SDR
ZSsw5Ye9bCgXqUtLTGBKb0cyXQBJ6rRQvpXXHtvR8gaRRmHMOLcyMUBG2fC0OCmz
0ej6cxQAdVTi670N3Xl9r75yBBWrFxaFhfhqAvGos8FJPNE1xmn/PjZbLJNMsuEw
RaBXpovwv8HEaFCak+duMyHZKg2PqneXkRaQU1Hy7D1HLj2m/YciXqomN/XNeOBs
Qcy4637E5jNR5woPFOlrC34G5teJXNlq86dNhPdAzDlgb/3HaKM1nlSQz+OGvyJ0
xtG+CSELFBQCdUFngsWnvjUsutRzP5FZZwY+yZOgwxYAyRdSPd4a2cxrV7SVguOp
Ki1SIn+09p0b+2xTbG3yPSL8eSwBdxiWnWl+1wkjbll0j51PtX428NtYz47xSFm7
vuz+8BbChjaiTEetC4FnsXR/ZpYlD/1ptVlP05ebgYYxVIsiQrggS3NPOFxwl9Nw
08M35EPtVJQqCxp0r+SBZbPRvFATac7HXaCj0oCDiju766XuP916YMkHdY/hqu0W
qvvFa6HoU0a8gVtDrgoaIo+BRpn+Plp8O96aU+cU1Hbq5A4NaH0S08h2VAoIscNG
U95z2hy3wPQ1eQRQtSL5GN8/42BzW6LNI+qcRpU2Hz10296CrjFrPtqHCNtzX2el
deYaTzIAOrevKksBFX9tr/AIKG6EMV1HoCa8HEvgdiPioycLceojtZMvgUSFrg63
n5TtpIZ0Ry0NS7gE0N9GwuLxNz15JWyNdVpgrSjuZiEYOENov93VngVsE5bQ4ZdQ
CI6qa3vJrMJzArIkTRFR/1oK8HUh+FtXiI0GwGgkk74/RjcBPnwnb4n/Xi7T2xzU
A+L0UveNUXLYtn0dO2HRuyhe+DU3xYBbM0sLhZXprDP1nqWimjGoiTp8vL9KoWau
1D+43FAspU+cv65Sy/r2NsDflGWufaFM4i7gAo2ekhHtWQjPXwRFr2NlUzw8sxUq
pH/a2FknuvaQJ8swayT4oOt5W7sJfRmFUW7isMvLxGYQYtuP87xrrXzIsENj5NAF
z16/Oq0Lb5zOVq84K+jqAjhYMykLJNfNPEBpBfbzZ+q5qRDuKvNHyGO5gVXcPv0G
llMcDpTdJoHz5hIF/C7kAUVynqXcbildAzt2OcZKPfwIoAFG+U52OGwb9wauJvO5
B2U2gM7Sj4YNkluGBNns5aeNAGtv6mt/SfSUeM2GCnDufE+r2dwdSJ3E2guRsEaz
RL4jLmUnuKmCfyfuiNb9ohILOcvCfzv2rr+kF+MynZNxhAYSjNLk/U8g+liGKH4F
cUeoOIqz6gESYV+7Xe0+T5DdiB95U6YQO4sfq5UzznMdKfW2NCCJ/eSAoUHIVkW5
WcK+WoJ9ZMxCXXOX3rr9nhxg7FrZCxXKuPNrKCm+iZAHyJsL17Q8vixU4TcbT3uE
e7NSr3xUomhQPFv6dV8VBDTGCOaYoLl+NBHXktIyS6WEHeZysIq/3BktvwvEst9F
8yfdT2LdxUfUZahX0EIn34nBwiQHJaB3ZdgZ2edRE+AwlqYmjJSmSsEuGhbENWas
Z/PHBADommxllV8vagLnY6YFiVXQ7XfRtUSxZIsyIdE4PcOwd1DAZFILLZ+rlxM4
XumGBJYh/dYTmKd1sbZqLoenlE1JLKFBfaucUUeL2QWx4hB7B9wOdQ4ihZiH2VVz
YAGAZOCFQvEtjkrKLIB4YfZs0zS3TUHsh/zZHJcov+4V7fQVg2VGGqsyT1Hq31lS
PpGxxYjUlfSQnxOpMrYFZWIVi1WNMTwT7tF8ls0AwD/dP7vcWh+v28yJzKmDzmmk
Dj/pSQbv8A7aIDnkf+s1BRx13tvBjDpqDbjlgoPDHwZwHguBDfteSW4h57zgfICs
DiCEPZ+W/HCjjWHlGlOyIM51jiecFc9vWPXUVo2/Ovs2okThSJMGR4CmumSclt6U
fWXJIKF/2XnDiR8HRoQWw9GQAqD550qq9zaMFGbKUfVJbfMAOBHVVou3VeURiwMt
hMIHFUiDUqPgm0bZaBLZuX2eDhKSS0pbugInGknCB+rrbyXXu2gUVwMGIvpiqi0Q
RqXC2e/Nan/Sn6oE55xtQXaPAsgw15g/xrY+RAs0jGh3VzzO8hBV5/NVN8MB2IFj
Zw7N2zTIpnTy9y8ffItMPsVvAYlJ8ldPVmceEBMiaPIYqq8Zo5KtD0luFYDUl7iW
lNqE7QDF0otLIcYIuG29dm94NpCPsbq947wGdjz65oSujAnXsAFHhmKKgxb95KAM
wRoTbKVsmgxM88zBMoxrE82TxT0K/VE/640vz82NJTdYVRhyQF+b9ffXvZ4OHNN2
xAw8IU7HmVRsmQsHwRGwPYkDPil3XyFHnRrrqIkbgIaOMRYuhf+gPTZ+lsnR8J5A
xIxDLDVUOGroOhh/+dRC4WkzlaqUz0NPxFskc5sv7etsFdwBQ5wd3DTi+j4yN8Tr
gNTQC5iTbSv17BzTDhU3dQ==
`protect END_PROTECTED
