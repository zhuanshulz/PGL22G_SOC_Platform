`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4JqUnSjM8qMBEhvnf30tYaQhZKrGoeK7F4VwFJdJKX7p0GT/+vBBQfTegOcguWtv
SUZbZxgYScn4xur66b9mXGRbCQb+7u7vVv1tKoBh/ev6KU7kTxM6IricG6xAoQFP
txxJOjA4A9Tk/8ySWBuIjYKVrrPRSl0/HoaioeTPUH1Ahd5oA3uQztBzXmlzNqiV
Z1dw8RCfBABv5jimrzf75r/USA4LC/vdAwsCK/TE8M6a5k5EZn+jF3RRX/3bmykj
R1yDDZYWIOh91XCvvgQCWg==
`protect END_PROTECTED
