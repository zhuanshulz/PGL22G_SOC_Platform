`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
erKO4q0p4SnSY6dGzOSbSjC30LxD1e7uxUoXjcDAu3vOTkoMzP5MDnDufRuTuwv5
tNXPZImEYyI6DUt2g3d3N/sMVuMOkDGz7MxmyRrKssdwr6vImOWm3fUUbQQ6dcJC
tH/Jh1llto2ijpfqWulAZMKp1aR/YqGcmc9CGaI2RYscPd0JguCKkCXBKnq2Z+zG
KuPDJWk0a6h+I5bzpnQs626CdblSr2zVF0OIHbyZZqV946QWFMtLOrC6ofV9KFcd
sCn0q+4/IDTW6IEKWDJVVL3YGyYjVbgZdrva4ibcBMhTDhVcb5svk1WRUDYVtfyL
rpEMNj7wkjHIVBcCQUVDFMVMJGby0bSQf/Hrr07uWJmmpLtqKuJmozTNGr2bflEP
Y5/mYPA807eTtDpdTJnmctOHlm+DX7Mkkwc1SdGd9K5qleFbeU2gmIyW/vEPeWmU
TefLqIB7V2xOzPWHhgra1Mtaa4K1mcTlKAh0bdw0+C63POUwOtIqxtelrfeY3pFa
G3vTIR+0eSUKl1Ip+mwzuEjhOzSxp6CBV2YOzkz2wXGemIkMO/blG7V/XFH4fpKk
UfwQMs8fxbklkQaHDn2byJsocbPJTT9hVW3Ih34izPyZ4BBotWbhlqyn4rV054o5
KYf1T9/VtjRL6URyt4bj5T98y4UGjijcmz3dkkUkqxEN3xQJAVQsQVasD/LUmrfa
TPnX2H0P3+kL6x+gVd5dHvCnMZGI1qFO7y0OnuZmyJRkAYsPSQjpZL1SqxQ0hYh7
18aaz4ETgAtOxvnp7OAh5P3QtAYN4AcNdlf+SNSVCyZVU16/WsreBv90lo5PGoj4
Wa0kmAe6LJJasjpqzcsclu6q/DCTKTVrH9Lbl+rBlMdjH4RTFcqYJAsuzuul/lie
WeJ1vA3K6yWIiQ0f+S2WkofBmLuDXB3qANdc1S1PZhKQWYAEsGwKylbJidYRqBgx
9aWUIl18XDxoNR37eCBBdQ9wDy7WyUSVSi54RR3jkKBANSsiELwOeW+r7ijVR1pp
wWSseVjLm2rjpe87vaNq2eOQ9tENGArb9MUwyY1z+L5i/3zeo8LyIdHu5rtnb+Do
V29kXjIV4qYBorN5iVEL9+2p4flh/SMCCKr4EMVyD7Wu5ouFCKQcjGWOtOFHM+CV
sstEL+8c9YYEoCmnc/o8KnNo/B63khFAmdJtml8ofXKSuqVodUskKhPU4rd5P5zH
j9moZv+zt2IBohlpRQklQQce+xFBNih2FXQ4fAxVLvwdJza+YKliwCd+kJqt1/cI
K+LEeoF3IPZ8ZpxSY0fPKn5UXNiQT2+yEVmkdwMewOnNgs5zdzhBAT8JIh0C66Dy
OnInsG97L4Je/IuaQB0V1bjA/gSH1xDnH/H2UOQixHP/QvYtrZq+ok9Ab67VUi5W
vDnWmqaLYhgAyejCiG9bA/gfa3L/j+c0d3cA/A2L5xCjmMEpHwDI/qS68ihg1ipf
98IL5i9aAnZMrZNfAxbzWSMMo3riVGM25MlnUizSSdmAAuGLNP1j4+rHDvOctxWn
1hL6HT2aJrMxJW/bzgvEf8th82phIywt4m/PhaJqWXqNAIMYc7vcwvybaeWrSFJo
KjAsD1PYVrmJg7fPii6ug5w8rRQhQtxgsoK7Fy0CSD1sp813782KPZnVYBqpwRNE
LfMJ3VfLFGyQqb6n0o3lQg716sAYn9uvxWZ9M5auwSqD5m34IRbMoVSKY5HOZEEp
xO2lUi0ntn04cb8CkF0K0pyoI2CADeOlsDwhasuHcAWQEm5Vsg6ijuqLcNtU6Fm1
Piqfk8knC6c9p6+BXCcjO6pfYIsm6ZhbuI53CEfT5KZQjdBy8+JKxO19fkrjhlbh
0KxJOU77XfkSw8/bTmIhM8pPzjWA2OB6bPMTNUCxGFVBy1N2erUF9ijgihou9iQm
Ww17fWW62dTeeJZgX8t/CkwXdgKH4pvFxxcxrBsSq4/8JpUyAYIeO9JNYdB2xBsf
JzpVeQC4iFgblJ9Q4mIvitmilgMnCLX4s9mtj5khvzsa5uyuefN6PEda3U3ZAz3W
r4hXbF1DxtIstooQ8xRyIH7Cyh7BxGfiUnxKB3dJIi35xU0wvIcXiPoozTwaykK2
IY1ogyvnv2FdAoqYhyARRI9fWKhxbPcYeMjgVJLhwtzL43PHHrqN0GzxxOXa9fTu
pO8YY15KCnD3Y9/HTrrHZInmzw7TE41y6l+OhgvvlhBGQ9vt3HIq2JZj29YfRCmp
mhAp7+eOieLnwnhhlO+zXN9WoucRsWlfd+Z+yBRLbpooVhNT+w1JtNLVEcEsww3e
Uzk4rLuKdcWjJeAlKUqHlPeCm8ZesAliSKzzSeTZ1misotW3WYQv2nnRFIu4k32T
dNsG9imsu4m9kk3b0vj2dm8y590ggjIfw4PYa/TG30pspUrvoMTU7vyHxitI3IZ5
RBSm23dBFPT3rET+55HywRaEise/JkEFr105GJTOXfBw3nshvmpBFyy9Nm6+MxV1
tbu1fZZR6Pcd+qPXzAW+Nkc6wwHlbaU6LFZBBrSHS7cQlcXaH6YY2ZtXP2ifCsE2
3bcU8RptC50INbErwdvrkU0jNs7C664fR7aOIQz6zXrZ/4DGV4H9S4gHw+VpUZOq
A/1Kbi2Z1GYd/TePA60UcA+wgopb07HraB2/Qz1ZMK7nPR7e72dGpE2h2DQlO63K
UoipGYHswupie+WUMA/vX7Dfpn2dMZo8MlL94OjmJJ6gsX+wRl0ulhjm/wkgZyM2
LsKqcYIJa4JtzQXLiRkpNFpo7EkFPx4YBbRyqAG3GS+1LW2St1iDhzlDl8xtJepw
cXvchHnGIRATdcTWKtiV5PZuKTfI91jXJFZPaPjbaYqYsx6SRwTQVjxu6gBJSJB+
ZWVbE02SpdfLpYmGfontsMrrILGTzQSmDeqhfiPRJrtj8apKzUvi/V4RJXzn7xWA
zrNzsV4SqHeE59QjuXKOzVlc27D2/8mv6NBEWCS2iTE3xLGvwIfGlGSRaESdSIwS
SW18FZxJRqkduwLi199io1VgZufZOiHTAQkBvytuVUOKMbKM3UXd0Q6Xw/Hgyc+e
0+XZc7/XPjhkpwOzLNDJDHpQcWILjSwH4h12E8SnPaUJz+faN0kNzOsik4V+fM9V
E/4VHtNBMIBlwkAanf5REBd03cpI/LNArjXU1b/rgjxPsejXXoK3QKG0WQEAp5yq
A0gmjf3kj8wFRIvyLnWIFLoKkZg3ViledBbz1BNO0fYlfCV62qAXhQoKns/rvNh1
0nSk45nZuHOJ6QbCBysJPWC3jNxvwsoVjgCty2/P/0cINRzbyWQhlBPRjw+1KMOD
cKhOs41GX69owpn6Revnw4qmI6wiDg9A6mQ4pHdrv73d2RUrOsmHzz/sFmlv11Ey
7rZdfh0Me6SMSgG2VNBPfDAMGiufFMVQKLHkkEhLJ+AKC7lZoB3BF1P3d2xiyTAw
0mXG5hQKneP96u7y5ena2t7WnoIuM5sIdPw4naswN8BXsuAlpboeNm2YE5y3tH70
UooCDaxSA/Q0i/mUT9843IGcrHGxdqrgGMetbQ5g4S3CMxWhuHBdR7s7Qmh2XO3X
70uv0XtT4co5RfQdmR7TIIRSdMClGrICaGQoRXRzcsKMVAyNljfsvV4njiVGDuS/
EvqKrwMq4RbDdmPO181yaDhR/R2sI4ekMSB3Ess8YbJfYibqvHKZuoRShmOP2WZg
5wvVqm5P1VrMbPmpPZ71SsTypWDunxe+8Hd5/4vFMmnlNHwc/J3ZISob6TwqUzF8
/9KcP3+b5YpdZ0dGqNzpgvnuE/dJNsIxww+nrLE4jZ18rq5MQSpE2g82zPCfOql1
lGS3NhxE5bK96/tn2kxTY6z3FM9YYAK4dJHdTj2syD4D0773NeP6ZNnhWS9gCiWg
nAdjtAOh9EeDXrIHpQSQ9zqQi+qS4JRbwGRk43+8BK7/F6u3N1De2Cq0vUOdsqkg
JskcChDxxE+1quDvi5dhR42tR6n4GoW0bjF1dkX5mnsr+NjNEE0E+CFnsJ9MzXD1
KnznBGAM0NpNjVa/MACYipHm9hmWACGtdnP4Lqioasw2mQ7+zVU9FR0vGPL2Hnrm
qcsMHwMgEv9HcKGE+b3PGwDdPW1TSGLbbXjbiUMpEkbVCw5z3Ii9Z7WrQFSPuPXm
+IrLu2VYuj0AYIHHhSAJad4RFte3yjVv2WoGRLrTk7EB1w45POz5ZV1wHwldU5Et
tME6NfL79su9fVnS//c44d3YIeYnX2Zm7yTWpvoOiqbGDBHiGEY8lokXGCATN81j
kCSeYP0v9P7R/mqUNUZs3tl3GUYwDBidEblVMjVRFtOkfmlnfxvsxPtQdEnTxMj3
eNnc6hE+Dscs/ERFNcH4Urr1NZXwb4jWR9VyCu6KSlffU3dFFH1vqf8VpEoKspzZ
c244S1EnzsxATmQADv4hkfozz3CDyN0mUVut6S51lMJvU4gNgL81LccxqMaGF36O
00zYcc4W5QCHD3nl4m7hV5U8k5T+a348LJSUEQPw8Xibueg3mRkJFK8j7n8QqncP
b+vj+Eoq4WTAHu7/Cd4X3pI8HWO38Fy4TUxratAbfKXHmC22DkZ9saHhqhELrEZR
1MGpHa/fZNzR0Y/G72Vj+MspP9KH4LJSua4iKclEQm0UzzQzcxVUsU6Hda4kle6M
jbSv8cSJZMnZffFYt9bG2Z7/IQ2bcnzzv6GvjJD8sOloaxoWJLrYyglkxTzO4k73
AdCZYOvZFv5WEvOmuhRyTOPFXrssS7GKI1lZ7DKY92kSgrGGt4L9rJ+wFPBTB7dr
ZcTDHGOmWU6zxYmfWd4RbX4J/LpAz4CoV/PIdIN0zoukCwcisKOXvTrVAfazMOZA
m4uT2OdxNmZd9zmrYNKU3WSNBvRxzHsLlklS/OVnWLt9zKGXK9T+iYOI58Yaz/Xe
3+tLueEhlQwC7oRHZQ4200hr/OZ9DVuJXfOFZVKm489yez+2OxFEEItgaKuVfq4c
Cb/Yskcx8P5m4A4A+qwIzGbd371HmZMXoNA+VRSDnLOzpQieBvZ3N9aruVxDLsl3
1OL8Lh0RXOCX7z+R1A6RcK7FQLiWk2K1SHWJrOVGV9F1V1VyubLCThu6ZZ7UA6Oi
AOjwds4IV08rr1B2JOPbUkje/59hvou3kG10qZgHv1FtoDlno2mfKFvQrZIYpfiM
XJdaj+GR302U/RM9VTFlTT1whVNMNARBNa4Y/ng1Pgdu/2C/CNzgSvpg0nUCLGLB
OaNFZz1+1iLGIVX7ejqV6U832tiJI/bU4ru1Zqdmr3Pk0wqkMsF032tsdSfijpEf
iSl3UTey3rMLoGrW+zabETu35hprCws7K4G5CUWEzL1jwwiMKW52PXRIvmIaFs0i
74qdNoodBMBYpT/o55I76ppKzue34mfO0mSJD5mM5j7Npn9JIaCdt/1d3DPAPund
tP9IJ6TX6aIRD63d5J9Dbgm9FNNzapSq927BD77RFNXCsuO0kg3+3Ny8OIG3FG14
1L8PWxxA7hFgPJ3pBCcvXRKzwJcoNWQe5+RbBjtR4Uy5MBQUW5Q5roXvS9AX2fCn
`protect END_PROTECTED
