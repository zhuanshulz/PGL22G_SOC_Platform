`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vUAHILf0ClT+2/G8x17yC+gdfoOVSFG/KGLBhObOWhCdzWPe1n9nRX3id/Hr6L1L
EsgpJPZjEIkB/tf7h/g4e3M7Up+5aXJdENY6nXqHhZmY2c7b8VAU9VCDvlc67QhB
MfF4f+w4tl8+h/PhJ/6AyWKHK4rBRm54xwNMKwULKkkpPwxBp0zaJWOOzEp8VbF8
g8RPTfEdn1uvXkab3AsPgrcZTuHEhylW3kDU9TWDMegEAryis7YBCvJwkTxi83mh
OKgzlds7uTzncxZjkdUyBWzV9RG28CHWd/N1LCWMvzQTIKPP8lAmYysLUa4x3O7w
vz7A55Jw9SwKh7PaaY3Tfapm0AwlMyE9YRBQNbnUJLbPYCATYcAIDPmRiTGZm6jw
audauV52pgwvS/mmg0OSfnFsmHZQlx3w1HXtwDN8+om+sB/JIJydVuOfRLoUOhY3
dknPiM6a5C3HJDERFbR69DG0sOr2kWEZDWio05PD+x/kK0+qWwlxHCWl5cHbDqLv
22MlJDtHQkUoAqVV3FnL7+pctfojKqqQvp619xsJq95E2EpVwTtdfFkA8e+obI4v
33p9cyYQjNQt54o4A0kN1FO14dsNe3eGEbpPqOmgDl70rdB8JFXLxgXMj++E5VbU
1cBfcwLjre5+4vGTLsxFDHjn6rMpM1dTvkLbZ8ajWA/3YHj++9JKCmXr5xWSCFtT
O/wq+sjTBJRLpW00eVKLBbbpO600IJqCDT4iemu5jXSGK81gXbBHxI/xevbw9DmL
fRnYuzLsoSlLiuYidsw//XQEKPx9/klBUY7wn5e0D80CLV2W34J7/jO97MihKW4M
G3Kt4gvdEtfa0aaxS6jFRdSo8H8/GGz6/ntsiOd1D1c8Sci2XcncBIupY6jBY6ZJ
TDcGadgijRuTUIDUwVxUNeUtBl0yAfaRsIlfcKWiHytksCeRr/JqBmeSXN5j0i3C
WRKkWXz49GR6iWtAau5wA/qliM+aQV9uOK8CTvdYwIVelTwGy/1BMnTTcw+lyNTO
HTtZGavOZt+xo/xjZRqHh3DwxCN2WBP4tT5lDL1S4nNJrZp9JwgFe8517YsW8WC7
UQD/mQhng/3J2p9PUG5ZbofbFgAWzyPppefyjtLRRExsJehA5X1Tf11Fw6iMOkR1
GRg5HsDksyMVr8CgQHqLOuQQvG3dhNw4rb3BxIO96DSuByG8LgRbzM6EqRc5OwvG
MTNygCeaDFqmWRjTEhLNWddwKrJsx82LYenQlA+XVyOS8UiOCXZg0mPx/No0Go/a
LM8/+ep60FwojFp1b8u06dHf+Mcfxf24t0AyOdAiE8r/3t6DEa+pcwknMhFlhCF9
i02NAZpRRjM77cbnmoJkJvsm4rFFLoiQrH+r5l/1/AZqNgoaq5xTcMdkWFnONOi8
MFGNKJDJSjcvgXIOGtlSxQv5uQEu+Y6Vmq1wzBw+xWYDXtkJwBi+m9Qm61goAJZL
27dFV5rk21TuVKhGl8tveCeGM70P0caS61bhvOGEr6LvjmjTM1lGFcj0tmliMnyF
cYtEEGgrCW7UHmIgKgX8vTvlAGyeUbYjewsOW0RvTKGl6XizPsDmtPZyuW2dhLYj
hY/VvJ1/2uzFs6JkSt0sWK2nXoVwJM2umdrJMckQ4nh9aeH+lzE18H4d6N59apZk
PnP2VsNZvdRm05edp6zQd0S4iQtyTKKxzI/pICRhV1CdbfEI9IBIYIiAsLG57orT
K3fc2npNCHGZa04tZibi8WoaRcGueUXGKuchxTJtJBn+QAoBw4BYC9+PWRZdDFHl
ko/oIm8LTIhAFOzm4pDv2kKUOpOCcBCK4M0lTuXDRlRB532BGCw7djWT3+emGRmN
H2302d5lIWT0IaNq6ukQ32g26DrRPQVhtKE6TOs527Aq5AHp54O5oPRzrRhHMAZ5
r7gfjBIbb3G5WPI7Ugj+aqlHg28V8UAQuCCWeFGJ+LGJKMFK9xff47Qa/bRWHDhb
mKmAMD0FH00bso2t3u0YFX/g9oX63Le6Azr0EgEHBVg/mZqk3QXfNdrRGS8geVDT
R4AX9feIvdP2InFRgZrGjtq6UecWchqT6F5IGzFxzS2wjOYVHYWT25KsCWl9HZ5L
QsmpKeKSDIzCCGSeM+wjnksJKcwUE0igDTUfdZn3MHMqjHsRbgSv1j0DiN8a9j99
nvoGE2QCfLaDzrgDDx4w+7oOajzsWqc25HrmQdLlxT1u0cEzzTptSE8rFIOLILlk
Wr0Nr/ihiZRhd/+OtTqo5apTb+YvVdBA+UGmhFg60Mx31RToHCEqbw/rahJ1vrVT
HICkv8q4VZmQZoJ5vkXSAmgiwCXmDaP6l7x4aRCz2GmnFV8r0sRwNbnEJCsqdWul
d/fxdn/+sX0vmpJPjw5Qe+GC4iiadHDJUJVgFIwEFl1hJn6ox5m3Tu6sKv89jt9L
n41sL5MmUqr7D3bu6+jLLqLfvd9eyQAIMv3EsbrVfdjgjjvUYZWMeV4bqbAIy36G
8FUhgi49GcyNFoP42JYHs4SWMBlzM+3GutKOYZMKNuRPU4WeE2xCLueM5BToBeTZ
quY7qfmUh/0nB3A0blC8LkX+CyUe8JL6vSJopJKBhmoPMXxqmarf2EjfyJ6xTlKa
O7AgNezFjU0kOpja5ORKGmHXxdhbgFyR1va0lYSx8dxSGhKxMyiBiAskb3tj2Jow
GLGJ5koAq0uAk+unU7IYGySNcZta6pDh1OweIx6sjgBnGMwuk1sgur+D+x1RRsB0
XlspIJQBRuWbGYJ3QT0/W7i5wXbcCVM/EUSedvFtXx9pkgGkvhVVXOXqWaI45rsr
nOEbDxel7HAO2EPQFZzkSbZaD2yeqFB4jxdK/Nx61tvmYLn6fyk4a+8W6JCahsau
UzriwDF7w/eosrd9Ju7YwsmE4kQttMYUf7/TMpBldw3TChVqjPFJxEjKwyaZjJTu
B/jTX+r7zzn0KZKjXyrPQuOTJE1v8gSFsp5ulo+C6+NGuET4FtCtqX+3/o6TSSW5
gUzFCJhUp7KmO9EaM5ztmy7UdRgyNb21TVFE5MN4E+rEy9bYxTMFVIKCwV6UJ9la
XPXu/pA1U9WGk9rH3i9+JpOy7hoEZezBdaURaUc2V6QtPzgk43OKXx4WxXfJvxr3
kTmz1LpcRITth9y4S6c3dcZb/Y65QIIHOdo802Vz2cRK8bSoJIdXeW/PiPrXQMuX
K0yyRbJghJ0cnZ0qaoWh7cS8Oa71R3U5Pg1oxcZJNx/1ehgTt5WgkYZEPqn9o8L4
VsE5XNvzYaxE2T2X0hSMp0jQCFnQ5081dLBxqTvK4gpg6HIaPNPQ/6j8Als09s0f
GK5V1f8ryti/C7+Wr+2LKkGmRFJXcTsvXAUA2CEJKOqw3bWA3vElQSdlYuYD+1Go
AiuDQwWg1mmmQNYF+2FOzmV7wSUUMR2bXDd7nWKqqOFEHO280Azzx3LpmgEgNmez
dGZ4UaTxVlbefXXHvgatvA7XY/Yy/96DUEQrhEpsW/Wcf6F7Gw0w9S7wo/3TD42B
nZFskfvuewMahbIBKTMiitn6E4hETWkeWSt3azOu4NA14wkEaPjf22TFkCTtSmkq
pgCGytf4ldG9tJTGrUMt/JsGxokB9Ca2SY7DAzzeqLKyxGWShvKhBAEMWeTRW77x
GBspUsTrFGd22eg8t59TsIR9JWzlNigMltaov1w9/TJd/qHi7xYOAPbNz4E23of6
rsQKIC6PSCvow2XSRufKM92GnXMuQ9lEowr/IQ93kAyzXKYmebnaZZbuPRvWYni9
vHJNJlBIQDcG0tBLS+5kUAUME4n17tFZgWdRfvPIdfoWdB1tVJwuJufCz+8W0/HB
RAnMaCtG6R7q0E/PkZEsCV7OIDyRvZw2LunI1VLB6hL/jkcnXJ44XNiR1j0OMAEy
OIxwwflR4BpTkJYy64OWFxEvJyok9/AyA8onN+bayjgQyNYt6aI+zFrSH94FyDcO
gMfBDBeW2RWEwrzDustMdwU1V6+LnNSQonQyKtgWw+cIce3pA/NYZxUJaMjCd6aa
DMLuy6y+7aYWr7AOGyekP9PfC96BqUTtIL5Ii3UxDlOVIVudbceXOaa1Dzdqkdvo
I+LxdMaMAMaXfFoaehf1UNxhtl2ZAYiUnY+9M0+EZU+Dgflohi9JLkpqyhO/tjbR
RIA7UXyTGbfOf0d+ob+HIxBX7y1qKMN8NVCHLf+lcHbFRcDZhRM1SOoSFlad5fHU
AeP9pPhyyCGHMdjhinpMygcmoeS9k6ptdPQnIXX/Bd3cGH77oM30V0odvxxAJkgX
X+XS6PDNSM6GKA+qe/IT0NmMqYDI2EP08To53a5W+pVDiyLDwAa+OHbvni+leeJJ
h1+JXEAvErENURpSGU0+1jlIU1hKMMYPWefwJpLqoP8D3bv0teCmShrVjL8XCewd
k8qgAd4oPmDfQzhAgDkd5Ry5BbJwfqUNpwWCf6Rs2cPQ8+cpjhw4nTOlrRWKW+8Z
OYERm8XA/Stm4SZs6UKdj8Knqhkwtc/dXBGeVTTyjKCpJpiHUMyV8530cKNv8H6X
IgX9VK0eu8UmcmS4z2Ynldhpys9aRPNkvzyxMiMxqeFQij+iKnnzp6Yf2S5ZMs5R
Up4e9espmBsdLCorRB6XUR3RbtP7UjscDtGDfoc2M5JZ9mpKxq0ApUXlATCzrB0j
5dDflitRrs4MtZuApQAf3Ce19+7Jwki87diIQFcs/mU=
`protect END_PROTECTED
