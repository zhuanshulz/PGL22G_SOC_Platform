`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xd/wfQ/RlPc4N47OdCZkyGMtGBpwuQL42feueSeQeC6EN91xjcvZyBtOoC+YB7L3
ahxJ41xjmaVNhdFYOLA2j0mfltnqaU2Sa1dq+8/ByEhQMDsHa/Yl/+F2sD2Cjedh
pTjMoBqiIPNvQJIGvC1Akxmw+RVzimdBWQnZEqfljK8lFBC50/bArScO/wo4YGwq
6g/FCA7rMgp7EeTmdiXQteT0iUOB92RjuAbWyJpPje5WsGfEgGWOgyMV1l608bQu
U0OSROVoOqSzI0ckwRzaDezsx1OA4ckd2qETlnWsnyt9/Coh85d8h1Fqkkd7Aqzy
WFlPwtdBF5nC5KXexHftj/DXGBDuQmhNT5A7ZP76YRtI0aAfTnoJSRF5LstYEfjg
b/lI4/fGU1zu5GJOLzPsxkEZG1s7coRN03+9cKuu0Vhnh6mKWTft2gH8AGmeJfLp
3k4NgId3UXM3gNYJDwM8xa3CxG2EzLsg5eLVc+EuPiZJbPKh3qPheVharfvfH3jo
1/10m2Fwy4jH4zCWcL4sx3Q+xKIV1rf9RhUbtc9BMzC1PJ8mirWh2xOcUdNA7bAk
EUDP3dos38jnpLFFGS5dBw==
`protect END_PROTECTED
