`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sYzrCh7y51pRJ0gh+2RU472LUVenpXZhEEfEVagiUKKnC8cl0YDNAM+wU6eACW+K
IWGzCb/X120vBr8gcp7hI8j66PI2El9YALpqMoe+rHG7GSt2/VQ/DbWCB7plO5ub
53m6gVczuzOEm/Dx6cpqqqFJWj72xwXZlem19i+ugVPJmFOYQBVrDEKRnDYviTi/
6LYuNR3yVmoJmPtoG6b8j9Czc3+CfhJw3/vq7GPKA0rcLDteAjD1JpjO897hlu6a
CFSpC5+nIgPAr8/BQMV0wFn7LWOQ8G2RLgarc/kVbXLgMm+9vmzJgtR/IWyiSg71
AowrbgnSBu7vwnsBhcwsmdGg6UdHpD758vEFbMETcVeMYVMgk/YgmPS9x6FAi05j
4FsDjpZ/zWLmu/2Kw11ObYUrCDTOvwTRY6y0Cq8U8ad32Y8ZjdYKv7y0Ogs/5NwV
Vj5+vNSGH0uDjq6LpIUi9aV8I4TPoOkTdQDbFfj5pGHEbmttq6Itc4EqpZEKdglT
`protect END_PROTECTED
