`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DAYXpgg+furuFmYz+rayPvDS4lwXudzml+CcMxeizMh6DjrcEXbVybUvDuMv/7he
EEFqEVldl33GlC+UsremPVWbSVF+edalPbfudqxEW17mboFMITjAzf96toDUB5b7
YcPpT7dJyoLDp4Pjr2godVt9H0j6Gf6QVg+Q/AMb6tx/Hu+Rx+H1cH1YKlMJMzfY
PQgllSse7ko58X26uByQfzv3aE24p9/+5Q4WF2gyUpU=
`protect END_PROTECTED
