`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SLsLEAl2upURH0UbtfdaICi8gK77PrPwOK7Ai23k1e7cGqRfX74GvHBBBTxg99ka
lH4P9+poM+JwRmsLoA+ZrF0jC7iY9TxU59qtBVzUZZnDrrvK3qYpTJSs3ddYz5ay
V+tzhn8cTmnmSXdoPey1Gd5t9Z+7G7mOAQ6x+BP+J+hZI/0YDamjWpQT1gUO1+10
GhRQJH6qCaUhK6h0IJ326udErLXgPKwuJXkQc5+ndcFp5gHFahEoTMP/D3UYQWVV
k+YNxnkDf2299nSJ3FjqJOoY4Ek4BZ9D8ai+I33CKVt2CsOekaeZuxjEvgJAEv3q
rJN55MUCtRS7R7rkDkNLWrGEpybzu/5vHsbkpkdcisqWfBpELdaHaTNQY1pWXORW
MM9Wv/8HPv73PUEIsy3aj7nRxp394vlWBuK8F8I9dgP/UXbwZJBPVeIRGHnuPQ+E
N2+XrF5z9hhuuZgV/waqA4aSd36T9sn1TLCuONEIzWuhEFB6tqhyZcqFKXfV+AGU
dstXi01ogKRHAKJvC5vkJrJYUPwY68ersy6fm6RIkcxi9pMdyxnfRZt1LqYfkDwd
k61tJ44do8NycTgB2725rag9Jn+kKKjrz0EWZgWPopIfolfsmLUG2bv8/kylIVFT
3mCULGyIga6Cc/igo63WHIEkzecaKn3FTJcZLvJwoqbY9GTAKNSXGAhFnAuB9dNB
FikaDLI5pHNcchz3f2OBVsS7qzPLBY/oAF4rZIHHUcF+a+LCH4EaWlAsbRKmPmjs
l8tGeDPRne5kvao5VA/h4QZilcq7dBB/ZWJxiQrBkXjg4zLe5OwuhKBS28z+2GYt
5Y72toE96MYgO6gx7A8/MXZf8JVixl8bX4jw4/WEDaeOm5+QteBoXy8NcQrtzSza
MKMUVdRFoPhLI8Xt7wP+w2bKR38IdJUX371MG2e26j8JbGvZcIsSbX9Iu5xjvKv7
1ilDT42A5KxaREOfZ/iUpzGvIGFplQNIh4kz/1IgFO19X61ZduafkPV4DMCoDMJA
82aR/hLqsXbMFUkEHILGJqU0Pu8mQr2qZ6diLtdDqvD3zr/sDlhSTUK/+qOUvDlg
ED19rcmemKoFbJ0DWCDwBEEDogCGoEBh7oaWaipfVma2TEioLCQtrvOh5TOZH93N
YlGHfEYSME9W4X9WgfkvanvEyg8/d2gK5uykDWNzoy8LQVyDZFWI4YzNHxMsBvT0
muo7mv9SPu4WpnsGikE/hWLhO6KNGn9dV3H5XJgEc939jB8P8mYc3fEjquiO8hlj
OMW+R2sivYGI3R3oFC1ju58FqR4oJmLsQwyRSgbz/Vywsyzcd+ZGnjyq/ShNOfZI
94zm89InLNbL63JK02jXniHW48/zlZQmCa7DbjpGoYBIzSBUXNeGifJOaHgLLiSG
fs8z4cOKkZwzYTpiIol0dYERo3uCPbLvJ3h7XUEIsVntvdOjra7nMfoLEze2Vg+G
rRNmTij7/KY4fhDNk3UIiGbaByrGviQUM496oS3826CSJJdzo5kBHYTiUPRaYm+Z
w5jmxTU5FgH4PxNWSCWrE9AJ301Bna0axW0JxnyyQWV6iLJp2NSCNyzzNXGtKhuC
MWbnl9j2vdDRl3YA4N/w+H4gSMKR0/DUJ0NEUD+zZyos3JwQu2HMpIxNjDgIQfzi
gCE1exPs0pnPHlZgNkqH51D+kDqn4bhZkrppdQ5mxAcXyQ1BMPRewHGH4THj+HoO
vg9PuhxKAtXC6jWMzFqkgbaerdaaDoFUL4ibkSB0VSO6Tee1gjbnqjardlfDBs4H
wX7WiNRI9jEVkAniCwzys7kUcBOgr8N0LuG1NecDmPiO2ysp2E27CRoKnkItdRHF
k5Qy0Ox+egSTX1x0Q2r9Rq5xryZ8OKdpRLymKwvWCvpPwNwYl1ULH6UqxKMh8JG9
DDq0nq2OtoFTsbfh/TrkmOW58L1In9UkzXOjrCE2NO+fYjOfyXv4HHrI5JuZd1ia
cCqRxL9gaIy8yIgGWgud9Zbp8BdlotMVWsNygcCgZZXv4T6HkyXMnQ3josmCDvJ5
EyaLYydb7OfNXn1gWcW5kMocOkjK8QR6ZyWHOw7w/kQh7upL+X9Oe/M5AtRu+/t2
63+W9uDNjKusY6hqXC07vQOfViFsw+PhHylA550pLil8yFIUkYOLU6iigVYSm+Dc
0paqwIsvBwD+d/Wf4Adshw2w1YpdP9eVFbai7dC+krfUIf/CmCBXi0AjUKMzdklP
RjxYde2nfDF+0N6NXM5w52Qcp6txi8PeCK6uyBVfie4Zhgznrb0wQzJ8MIO9ScDq
MgESWiM+2vmLZpqLBBTf6kWXcL93/czomRr4c0ZGq3t78DjBgSNOQDdu8YqocGVv
MgtABe/gqXZvcF0gCdD/2WPb1CZRnwyZjxEeP0Z4O/ZK+gRjmFwpXqcVQXe58nIP
W8w7OD5ceZ9aj7sKgkAQwPOM35kO3zzruvidnAj8pD095Zqsyt5/vtLdC3DJOh3P
p/mBC5WKlUfIwCknF1SvckzwWI6LG2kvsQd/tDAuYTxqp/ii/liQV3WI2jOUI4DW
MKU6tJ/dXNXifylAOq5uR1j6JEV/mL7QLaBboqvKgWnI7qkOJMWlxSj2NgGSUGHZ
VrziT36xp71eKW6TALTO051nIeR9c3uM2LLNRhi3q4hYdCGgz7XrRzIBhcMQmw5Y
y57SmlRI5pED4Cw98uYyjrnTxO1JEdVmS35sppnvG9qKuFr+M/9Nebc84JSMzDqq
Gnu1bMZ7FajPgTzWsRbIl2kDc9gQ8DTOk2Zuit8AZvTgs+/d7fzZDPBec04MsuRj
bdCD0BRpi/lScqJVoI9YqXElRIQ0cMIgdVcYXujlojkZWpYEdF22NyQwRfBVHMll
aw4hXQ94NPOfrcai1KcX1m++Ovs+XvUkcjddJDTxJN0AgAaQlg/8Hp4EXxqplxxu
bcZEgLy6kMwyZdYlV3uf+XuRxRLOf7eoDHyzJy3s1ZLC9nSOalieqyPtcSSZFU6N
wXI4UD7GF3h+GNDZOeY0l8VFvRLTvsU05teCWOZ4z5G64ZhXLENN9EqvrqmXHoZl
Przy5fT6JPUtkNvzZ9+wR6sZkLdXG2cQAS6Fm+1jd3AXHEd8Nh3HWLChyQsua9sJ
6LX3nOzaurEF935DEU0Xq5KKtkOo1DYrM5IIwPHSKIERcBCuF556SCmDHguRj2Vn
1KS2MXQtHe+C7NeuzJJd6J1pT/E322mNrcOqSHgfHenV5T2mhUFxYU3cdoPLPhG8
hUdV6QBYakN+0UbaXoTzHgHUkEMP2aZLJ8+c94KQ9SL44kSHYUK5T37EGmCubCzc
uDmsuT+me1LKCZQfxBsyHl6kBdkKlsNUo2++d2xmovp0qW3yk6cSvv9UKkNFYwXS
JOqqRisy/4rpJVMMV2zeumqR9NAK/tBYzLMOd72WC2an5GUAM78z8eNxqk3DdEmw
mi81Y72nxQra7dUjsTAb1rs65xkIpCH3OuLua3Nf5tt4kv68VYlJkHtsMJWFsXbS
9ilSbgMKe6FUIRbe/8rzrGRUCvAPvTB20bBgWO9Fv5tgBGesmT8sVci3NFMSj4MG
6PoCEukw1kq3690o4+uLstSi5NYKNTU0oMduOUcAA8D9IOb9KsgJ4E9epDsoiQf3
dBap9L1xeB/ZDtD1u1NG/gRuqcXO3vNe1F0hJ2O20GgEFOPG+d1iXrhIdEoQBdGy
BXWupFuA2XRBpN+iYlmqfZNOca4XFrO5ffSXEehys0KyIRA+oSZWf46hVXmFJ7U4
50ihCEdM5y+M0ebm9OLNG68SW++SSgi33i3LhL3VFAHG8ujSIPvKqkeE7/WRq0r7
v23HmDICUs1J4pmgRQ0A75T76meVpjWd0Rd8PF5R/y2iy4EcoKmItfIgIoZFZBgl
wYiDOoqWl0cD+AfZnrAsX9Z1Xy+Atdht6oyv8On1rKy1oJs2dSFPt2JAaxHFfeen
F3IJoQFBN7P5zGL0Y+WAMYUwuZze3KS2GpIhWm6wS8oHRbNffawCUy2HGHTy8w0S
rLxvoZbjBWbHHtUUM6KgWwub0E8wfhGCPRvrri5h5IEsBZkRNavWY941geZ0EKh5
p/y3zH40AMXQf1gmyIbP+2QekMoY3Ub+YbSNw3FvouEtLZclQ2qPsS26W3PMRrMp
NRyQreb10FomHInMoN6JT48q5t2ErwKbO/nRAfOMkRYXE9UU/94hh4KtU59sO+Xt
PV8ksK3jXmEGlJD773UwsZ2prso0KLgZZ5MrEmg/v6VDsO03qgYXe1ORFYzAAohS
ZoxeeZhbnUKbRsDL7jXcfxjMp9TijqSiv+k1mBaBNkLB/bE3v+jsDa3v0yIz8nIZ
HOAxVvm1guPEEyoWP0xGJHbuwVPEF+BHKx8moUlzuqblnFA+hFqreVrg0xIqJvgm
zeZb02JNcVHprR8kXb0n716F2/O8yKGhbg+MwDC+uVUJrUudOyW3YKPBE5g3IwzG
/+zyBxjucicdaJqM2ZcjIFpT94yovyQyNgkB148vJrjuhkmZ9IuJMAexO9+By7UX
bYNyaiZ6qoamdQbxJ3HaxjXNvtl8miCKmLe45SInmKoPu/l3XGqQ8qKCQnsFpvSw
iWVRSRZbctnBfe43YCVBvDGbr7hsTB9bKEA2WHs4FihwUgc/lY21uYS+48uTrNXo
Oi0TiW1c+gTBqMyRrfyu/24qTeN3+yMwLUVeWNiDODB8bUrVN6d6tdRpA446GMS5
6x8XcW9WAMe0j/wt10qqRykjPMIBkTHXVIwmsU9owxboMNx/A+pRa+yXFgqegysy
+PNMTaXEQjPvThdn93keb0VC+eucSTQXG2N47cNj97c95+CH0uqoVIDoVpka5hRL
QiA4JaxJAme/DLYkUG3szDI1EdRMgefKc7QRIdEVTiKXn56aPVaAnDv4KgH0H9nA
F18vfaej/noHqXSszqEZ3DwJvMLCmSW16d28SiB3LHD+ZBu4Gx3wIf8KpVN+oXmD
snxuCNmz9By48fp3fQl3xAajNV1NCX8hqB9FmtRw5fZ5WWTdjeyQSEnu3Pj+Dbnw
q3QuYqcAW41QQ6EZvZcRJT5wbrFztFS/VIl9owHR+cuyHc5+E2BNpob+l27Qo3Na
oqsztvD6+AgBxZ78i66v6QL52YR5CBUli6zvdxm/cW4D+YphdzDfQxICz+HMWjgP
yf/aGavRA30HGXwS45Tfpwsd6HgVkhFh2+heNNub7ETEfLD55anKbzw8GclyI2Hp
+jTx3BSZZB0eCDOaGX1OLQ8EfLL4x6pQox+iYXakS5JtfPn+NeRVaLLWfi4Ajzab
L5E1gKYRmulhLgCb8vbFEqe8I04jsbcMe0NqhXY5dYl0XgDJlBsO5ShnP+xjQSS7
7Vapva3qTuxdU+B3Q3FoJ/mQupUBlJhZ04WEH12c6V2VRbBy4R3Ex4EGmriO0kLY
AOrQ+4M4UdvaKrK9oTjmel35W3vBVvaz0wcT/r16bvwbgzg1tL7jYSn4mzV9qw+N
heSHKAIh0W/+gJ9eCTEWV+ssMWZmWZx/pSomJjLa5QISNSgsLoi4akbjWtwuQr8+
5AWE0i7/zKwIY85yxhr/lLudNsG/o3xDwlwgR6p8gpgM998LBiA2EmXr2FOS/cFD
DMq7J9hwPnmFFuH+64/FDNY+7rVtAlPiLorVXai7PetkQmDtxDta106Cj2vZUkRW
p7JbuAswfVNZUn/z4aNWLMEOkF6TWVi4zBsfgjC3QIEtUHJMt/1VIicziPDs4xIR
+JDKhT1CrooS+95tD2rMDI+3kFKN5ZVO7tg5iY5xRPwi4GJST9PCNhD4mGx3K40C
ewUYY3bQTNoHKW1xNfTvzd67qPQHuRWvkz9Uf72CAYMkntUUKId99k4NYdMSmeEF
YU1dzKcFDxR5o+WZSgJOVwsFjaadqSX7guVL39Y1Gcu210HMGBzHZM0taf3dk3fy
vsfNrFRuAsf/2dA0/HLYjA3mrBc88HlFmWOSXq5kqIaRu6xS/CTnLXPDQLpQbGpx
yYOzgSKFNZVirTe39mXtnd/oDL3QOhpGy/nWwkBp4NH6I4X/K7jYiVZGlv/iwAZr
qtFtzHN+Ihp1A4ZiUEitPvXNerT13fN9HBg8ftkhoKlEQqUYKzJ3QJT788fhZbSR
+8dhIOM1LZnMHsRchJzGVvDirdxa6u+fxkzU6OqrRQAhQseQPBu41oBlXkN+AUx0
lOjQcZcSt/OLBftnMCgEXuc8fVep4wFyviWyvjz2nu4A4fJ17mB9Jm7iZ535HTqX
8jLmTqiy9CejDlPfFxfPikZRnbgepoo84hD3eMRpMZJr+/jM/jCJHT5zBCZbcUUh
0YqY372aILYI1ev/ujD1NBxowcNr2Rp7xlaPybtnLJN5XJUdDTG3PR3dRt9Cl8hp
n5xSD6ZkqWNxn3S6csvMJcmWrkBunjzLWSP4NCow/rxDSTN73agJKqcEku46dyCc
IF/j5J6qwoUCMGoQlAFx1VRwW3bp3voA5avftdORPzco0sxs398COZ8F3ar8i7Mb
07vKt8b4espTwTUyZ/dmv335J/nGeAAatCOk0hp2fHj/ndl0r42KyzKhSa27mjsX
KQ8gZ+EsKmp/H/BkdNGN61Z0n0cyT5d3VYKmmCiqQOz/nZaAxkkEpsBvRcK5jxr3
SHVu6VtofCMqwmZYbCo7jy20sFoGuSZi4BgZL6tqhcqP+DFGxWciVkvFFb4Qxv+l
z2OfPyEg1LmMIahm6ge2pnvwp0YrgDHqZBUstTfO/Oj+xG97rf9StkYmCjPjFqd2
Y7BPLJHns4XNnAbwjyhTHkkEJ3HBTttR7tTvW7foVrRn22l4bQkpnuiZBLKVq7s3
z/FRTLYmhY6cc19cp6L8LbNmAJytGd9ca/cvwDhm0KZrMnrVUjXOmPLTZfYPMNG6
WEs6arRAafMorMgm1yrzPFzXoDD5OMsoSr3B6sctPW+XOXtD2lScFqAdy6LeN7Og
WqMLcn3kbKMOs2QDmApc+0Q+HrjU7WAGIZ5GYyA5bBtPBq3HMM5QdyrLaSH/hLTZ
/hZMLtBoY6y5xcjnaQ3wM1EifD2AH7Jh8oE7F2IWTN/g7jZhO2aSlmP002vS/S0K
AHoEaQnrWA3hZOVzfqg343MHeXwgq+7cIQZtAnc3YSgmpenCUqd3A+FrMRVz1qnp
gHYM6OT11pRHlsIH1X8k4fWQWi1F+ufYXTX3/7LOupl6JO6oPekkV7kC8u25wA3t
Nb7Wam6PMtq7f3J5G4uXljrHllxTrCIHAsbWIL7T1phBRjuIAq9tZzb+qy1voGkH
OkBzHt3Xg/Rkt6Ilw6oRFSGeZFKxdqDdXk3k/Da9sUqK3eSL8JEl9j+NfHV8BUik
xAgUnx3GB0SbxQE6LnKZjnyCoDSr1swYNnrEvNbMrWuW42r97SBFAgx9B5TkmdH2
cTCuX34RCl6U5KEhqxPrmhgtnWh3T+b3+c79oJyZZQ0PFb2AZgmXvWN8YqrVuo7b
kfONazqZkktR+y5j0gf/qKlJauqaCwPVeECnozaCELYlv7ITdE0LTR1/8ZmVNIpR
Ct0jcAX5L4TnPbhLdlpG5HMoEFSsPCRuFcdmaBwWzhe1Eky5xlhBP9G2zc01GVAx
8qECJKjfb9XnsV5X5MOPcQk4ldHhFCxdeHoNNA71APdAjbeacRWJFt2bbOVejWlJ
4SfdBGKd+DuqTrjURyUPzr087W0+rIQyskNnHXUmgFFuIO3DfYJw9BXGkovBvfwk
2YbM8ZUa/osKNyaSoup1DnfYPuyJma4WS17o7di2LlSnC0LxQ16xFRil13YVqax4
RKrVFzG1DNHtS/iFY/kwtwxuj3VXALd/mGNVdYCEtdo=
`protect END_PROTECTED
