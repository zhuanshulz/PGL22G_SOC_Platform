`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uY5nBqjtT1khuYdg3t9obpDE+q9CT7oDn5tIH5shIjTdtC5O3UZfrcDO8iEl5cSo
oCsfUGVJiwYmYrJswo3mXZPbgmyuxRa60GiOl8qw+CJ30lVC/diUcfWgXkEr9T15
+zVQZBdwFvVAzAKkMHhy9VmQKfvX8xKp4x3ddAHY+zTkw2kyZv9/xzJFk39eRJlR
H3IRo99nLlUj5LlcRJXaaPn3LS79LuD+iTGH5mGi4ReoheLFvjMTPuMpBIF+XLAz
ZdslJ5rzxALlrhEshVn7JNXyjFziMqQzOMroTAO8szOYgI2smrbnheAeP6QVHs99
zCVOe4XVpNcWSMCXOmevzMIz+B4FnUdzDP5LXWq9mUeJgVR46SCU6RL16aogPGO4
gjQpMIMLZphSjZMnrM0QkXHsp2kzb2WVyXV1ypjByHJoY8ZfWS713qWd4WcuQ+3J
VXQQLq/O3H3oRlkZPO1lsgmfm0v2W08pgNcNK2tHiHjLliHIgmnYJ+ffBXaPEdFQ
Wirgl2cuRyyTqLeOUzgt1bmkvwcACK3VT5jfZW3XW3a07UMXqRFGUMneqYRvvl2t
eASH1zb2CnmgpbNdvru02A==
`protect END_PROTECTED
