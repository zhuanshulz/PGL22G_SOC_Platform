`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
drI/E7LcVHyXfc0r8S7Rv+lUPAoBT+Y/10C8BEb3TIuaMHXnq7wMWJwhPezsb2Ms
jSv90Vbhh8CM88hRktR3XOI0/NeZ1kr6wrREamki6j1F60UmFUecvV+ZmmRbJNoZ
qZgsIt6niAU9M/C06MNU66hOy2dGPwuINJeMVb6FNZB/s/VCIdPQhcJ4PgieXaKt
itCeOjka3tUHVbwOfQTtHkmcHj9EN8K9IDgeuo0xa0pKf+qBx5+up+eQvfqtQc/6
7XqWHMAdXW4MgtEimSo7KliHeJqBPowwjnKTaqtJnXQwa85BAulW2eJkuUyCe3QG
Lbw6juZmsoCwgSnXtd8CyVbh58VdrGbT2MKXY7A857aEm0oCavGSKlgNFva5DEqI
NSqfE6Ltc/Z/nq9xStX41QSlu0YVEk7/sD5p7oCnzyKF0ojRbbRxux8KsWIrMe+f
R9eW52THdpXbbthu8dIeVvhbp14YerjYOneUcz/t77W4C7kHYgygTysFnuswAtV2
irTCfthJiZ9qVl+dT3DOG3ZXR2WkMdkk//Ss8gqExs0IeMSoMMK33OCZcte65X6W
r4kehc6KgpyHbtT1qeuCL4ytan/lFHnUF+BXyDSbPGKkon7sQViIUS4gqzNGdL/+
Ri0JcuFbPikl1yY5vDFClJ7y3QTPNsAOwvTLyaCQH3jsHHZnCBJR4nxY9i6lzR9v
DVakHWQhIDJhXJUNqhNwzBTweDEoYfq1Ev6XzMkLOuJ2qr4CbFVnrtFLns4jf/uu
dM9gWk4gtBI5t9E8M6+Q8Nx3wM3JTUzHc+uXwUIpX1OZ7zDzerop4EGbEcFZ+6RL
DnDC2cbZ6++KSvQgvn0zJpNVQNhpYgNVEnAU0g/edXHk99yW7kNQP15K43m6Sywg
86TfWuIMjrqu452r4qvz1UbWRCxY9Awnt5xPPgmH9KixYhA1FgVJhXzC5toePrWA
nkK+AHbNIIG+qNwqqwVmO19/hGyxa8IFJFGmLib42MN7sfYQ7+uU+VxNb9rA19a9
Ky6cwc2cLx4gXCiX7S5e9++LYl43kHwPppEhnWIw5sI2TmFOJNJEUt83KXtbTM1N
beho4RLB0YU6sXQE5vuVMatouO74UFNZh3RFLk6LoCoJpuiGwSIYu6KcfT/zgij8
KuYHyugO7DWqfvqYIoMQ1U2LRUMBqnLca/TiEte7TLlicL38XT9RTvV/Ns61VYzs
UpE3GyraiRKsVxUvENU92gglkMS35IkRMApG+snRk7azuhYnPin+N+zQCOmAJp9T
oFxDH6I9AX8un9pyceuXAj1uOxzg5i5UvCGPYnF1ptBvafh7ZsAbxoZU1UoBDc6m
6AmAryckdl4xNcHAiAE6DCZGmoqSFjIglK6W7bkLfmAePOwInlHjuGEUKzf79y4G
JUSnWfNNCyrEOU0dspg2toGeXASKZz9Lcb3aGfRsUum4msOMzUVSae+RBQeBk4ft
VC/ticu9iysRCEXYXe4uyiqZ+rn3LFUmE585rHvXwVQvue26GNzPQLv2C9QkjeAf
3Y6/ipcfPHvr6enIfwjDClroQhSAPay5pYzZeOn+KPZnJ7g1Jw7KHa76wd8Bli/H
ek5GOb/lPwWt49B4S9Ab+trMY2LgCIsZfgM9bUSUwWY83NzYjo6jprn6CNqdwCqw
GPqe8XGheHIz0ANn11mzYwADsuuScmHt78ePGTu5mC2m0nmnEbB+51iGTfL3t/JF
kF2qbiL3/Z5iG/sE1YKAAh6CVbopFmNkyHlCmMz0V69TrcCISV9Q7kUrKnVQIR24
DVEKrwoIiXrC8zQalxxYaRMgBV+l+LQEr1tcOdjTlMnduZqshCdtrlSRPkfxwib7
ocsu2A7zXjzm7Fk9f11DDB2b8tqIOV0qYVmAp/Xic+qrrOPi+YRrKzB2haazHfh/
yh08vKSOk9v51GalpshDHsyBxVq+dl2JPaA8DwEc0G7ZrDpI3UoXBoWjxEQYkjWc
1rTsG+f1StfRRJrLrZ/0zYvIhyvnnZy6ncnQNRzDR4tZ4EXwlyvjWWwu5YCZ/aqO
KssmJF0ms2qWpTo62Iz+Ycb4EHjftlZCD9CX+130J5tzDaKyzC340JOueHsQQYNj
1oFl2dM9WYjStaPlwCWQh0ZDP9p6Ig9oYTiBgy9DUknS2qvIAl1sBiCsjYyKPsfU
ojl6KZFeUp7SXbuEZUUXkvDEgS+/xIYWHJpX4hYl/R9Y9o7MDIsfKQtUOgD2nzZI
M9WZ9F68lt4KLoTv15BC1g19JK62QH5duTd8OJEnjciIWjj7YK6U5OIMekWItJPX
/jy6ktUT7HON0IZkc+yj0pXoYAQ8oZqp6qzEDX5jzLI3+gOdX7ZXw2sQua5YiMMX
7pMmitaHT/0ldpOumuUxS80tQXQ6UEti9P40yqBJ4cKeONuVB3lQkQbhCiptQwM+
dEdFtrlCUeIkOZOgUf8vkE+ZvnObvtsK/GvuCONkjHIS7xdZy6rAtkr/OGAEhkFM
JgHEi55wuS4UEKL84Z9gaKt0dRZpcLYKj/A1vv9puTtE5Si6L0cX6KklowuLuOVo
bnINyzeo8LyeNT2jOPJIT5rKeyFjJVfqYOK4V2SIh4blUgR1ybQSkA9IHQwNGLAS
vggGfyjn1RR/sXgWOJsqRjmq4y3JkmlPlFCKMcDGR2uPmKVG9kSat+hslCcUY1Ps
wXhIgC35IwgnVQxDzOZhfG/h9wQimw/EMd8Jvf1KAqivyET562woHWK6AY5QcLiH
XObocSLtYgWLVTFBZudbMRAQVW8pje+4BWYDB3iqzXhW5eQORgS9LRsK+kNvc7Gx
cxfs1oapL3t7PtH7/jJGHIYiAaNOzSVkmsJAR1XfCXFCXOJI6uxuy7NguMA3OWAp
VK32n25rN/4DZQDLa2y4+Y7Ky4d7/Q/Nmdn61x0dXv54Ejp7g0yywNYQDGoHWFWi
7gVBCi9Cwpbmm/t5gxVDrcFHhN5MzcRB5fAoNWOpS2AO5FKAV8lu+IKacx4ENjKB
UR8tMMzA3FfqA5cw3kjjNb1AYBT6vfmuA4IQXPayCJdhm/licqxrMKU4sZ7dX/SD
jZMk4iTpdTzhyeLDj1e0hMjpp+KgBd+a0c3DkHz7AIqV3kD0M6y/6W1M6i8myPeR
cUieTGd7f4Q1foeWQnUdh6pmNfoJ52clF2RG0wFuFpKCUVKFr5tNNxlAgCCALHcz
RIsDUTiMDf+q1tvt5ExvEnYbhCpojzCxUXDtMpi98ZdYGOUu6oxHgYTyjq+bdMah
dNgembfqD9P/nIEwq/8be+csaWG+cESmvA8rdeTgaf+QYBD/cRGoJnvmsflWHZnu
sSkqz9Ffjla6WtoBIMr0DAoIvmueHWnNYx7TPSK0jkCAwELGOxWR6TStufdYEqIL
7Z3P7Jv1YyAxnoQzD2nE0mk8HQ/3DlezYj+5gYryyHSWpBOVTY0ifFwGUfViUo+p
WvJBDKTs5duN6HDU1Uuz2XSBhdkfzq1biq4tDLdPqq8LKx6hDh3LHSDwfaAt+Jda
XhhDJ8byuGSgYAj1tT/QXPH4E18RGmy9vErRB1a8zFbLtUACBiEpexfTCdSq4HVM
OvSx28Uur9aTPsDFmRNBh9XcSPgATOvydk/BqExD0vAzTOwms+S5QrUlPM6lwmwq
Oy2eOSvoI2s4L7e57eLa0Hm+dguYFL4oufQhR9H8BjWNEcZo488kEZxzV5Jsckss
veNvh8ylohFduKlvd/N0lNJnw/hZKYz/cBSEXu/vlUIKstUkLjJpYnMYYMFhfg6Y
BELMwDjJGDfq8zrpRiGv9tr+bLa/BJ7SyjnljfyPeES4bHPHbHlBhZWpkp1Hn2AF
76CcVC2yO7ME8zR+U+lCE8XhiMAeG/VMHv20vMuMjmGf8vfdQNIN8XoGk8S3FC3a
17R3NknYolpwkAywsUvmChUo4dBRVUpgoyJgPc1vzpD87Z4O2dsYkEoqx8YEXFAO
BTQT3fgwnXyUcQyUAgv/1ftqH6dHVsUuIaqHMJ92D28Q12qY9mE1Dj8Te6H4e3Rr
D8NYRhl5/RImf1BjhXdHGhnrCVpy6WlI6zyzheDvVbU1XUhyZS/zID+3FcCmsteB
JxCxkQ2CmWJZ+7GoAjaCRuE8hXfpPqAbSeFOvigUrwLVc/EcCK20C+65RTDBd3KN
gcvCWP1u6pVAqroSiPOXPtk1OZBvJ/Mb5i4x9i3tgcejlEeYK6dbkB/wJmTDGjhF
28FhL2zx5+GNKw+YMvmoJso6iXakkSeMhXUC6o6KuFQ=
`protect END_PROTECTED
