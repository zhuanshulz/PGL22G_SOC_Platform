`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uhcRRfYIXqeK5RY5Ttwz3NjYguFgQUjaMoMlPzxSuhpLxwA2eUlRw9vVLEirDGRl
KTC8T0cmRQRliMTe/e76aKpHJDOpHHZEEadrvGCRANoyDoRr2NnIGZqqmFGhTwbP
1yW+BsicVB0Aiba8Uewcww0x+JmAGBsXy4B+btOyOSuuc7izNsB4fgKQQOQiT4vJ
RucbyxG2K/pbc17JMqrZSbeePKTdootd6RH503WzQ9hELYr5X+TtIWyj84tupF3z
Uh9N26e+qyc4FcL8rCd5rRwCZGuRGeiJChlebTfac07Jgp4nPzSAO/75vvOaD2W8
aZ9mN3jH3uLZwD9Mkz0qpptvHCW7FeVZjibPVOCq2vwva7K//llFI8gl3tNVrNqp
D6fSfdeLfi8ZCOK/MC5F4LjMLuNkkn1zhDI+rhpsX93zX1+EGt+lSUQcAhs+1hr6
9zEZuj2BwJbEuA3iRScuNX3k33/+VfjPcav8dbSVd9ts8tO/X8o9MQqyeTekhZP7
Qn8IIXGuX0SXs9gd9QXQaGQe8vDzXv5JPgn5nhP6NP8nVkQ+LnzKjOM7JNmVKGxz
mi0hI+xXGM/b6mz+69QW6zXaeDzn3Z4EO4IdjYex9n23x2t8yNeRtY4Y5LKdUHfv
Ym3PSAnyVv9PSuICEzIAv6YSrgczFTs8lO3HA3ldJfX0NH109JwwnH/iUZHAcpwO
PL2jDYXCrqaSd+TLZLt1A2yMlMYwPAufioCMQjc48mKwlDDAzvqjkjrsUWJtuFSF
MKJwE2KNeuBOq34LdanmypOyLYWKU1APNIO6knlqRryAppbJ91Ih+Cxza4xeDyNv
`protect END_PROTECTED
