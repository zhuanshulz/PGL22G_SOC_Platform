`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PpaWM8ftKAMnZPWx5yOLTfw4sxdlzqnt53LTj7AAi5i5Asp/fgZ0ymuI3HbwFXDS
cuYkvw+hiI4e2YK8PeTGobyW4HDjPkiTGc0IPP+VrOtmwV0J8/nriBMAUGkvv/DZ
vD43+7ZpnnDSUUdVVUTUFjAnmVAmX8pj8qYFK+mqelqbvOuUFSdOVTYtu9ipt67q
pl8R9KyZMXlBHqM88OeI0DGWfKAyxMJOKX5ZUf4IF+X7pxTvhQTfT4ROEYN8JCuc
lofE7l1GgKYNS0HYal3eCHolBnQWbyTWpI8uGSmiBN9E6+N0rrrdLWV19opsDWxT
FYo+blSKc/r93vsk9M5KgC2criEiqYSNJUcGrlssNcjWxt4l3KaWMQKxoVTLAhb8
zUiCWfWyLPwln8+eExsCIVHci9Tfqn4vn6qvVefjJ2Og+iRQX/nkOXiUkRBz8Q9A
aEB0sakR02+pHJeGCUVbZMzd9r91lyvEkM6ELrz11cz5QgqgGaFtS07ApSuBnOe7
hecIneKi9uYhLeELy1KMkiFIiF309oju0awjLi097VtFOBdqD1xWO8J+LMQPwpSK
QswsUbbYBGxQinU7OF3ynrpqs5d9IlAo1hv+Rcu6ilrTWToqldrWZ3My12eH4Hmw
m+R06yYy9STcV+tHZl7lG3zhzPDpNkbKZwQ77lEy+49uTkbyWY0/OZ5BKFkb81WX
2PQq3ygf3HWzUTbHDCVuLo3jAm4lERxrl3GbVNpF4CQhjecaKDbkjOMR8J5Z6hR9
ROaKJl+QdbxQkXxDG4+RtWZJziCnrqzX7JLFv2ZOKZGM8Ao+7/fjORetE5rtfuYT
BjyR89Td9dfmDGwoy20M4rPv6vg0Q9tfmzReMRTo8qKdK1/LxuhnfUr88vt++V/N
7fWT/NURqsFBeRR1SG0Hsa659NAT4N6UJcG9Bp8XeZEB+SYnzOAlop6bgb1AEno0
EzA+gmrXrs5fI0g1pw4lk6qRf93/Ktq9qCjB+i40fXw6LM7ssbelFjObq20gxBsr
kEGCaFSV1KR10nFJsq/S2sPjsZw9BwcfUtSVF3Uw1CW4WBdWhXk6lXnTJd5Q/KFL
1ItBSrjCa8odjMb0N0+1JeNVumWo4vQmO+zieCBSoIHKmvHSRQz2ghTr8s3I/0CP
OuWRTpNiMxX0hdZCbXRQ1XHIpsKM/qpEBJAff16mZ8DuLA4TpVTmwQb3zjfxOHLE
UIjXruRPkjUsNuQ7OJgmMMTF2H5dT5RzWY9EuDfDr13PtZ/cPqFirb7e/0Dmirz2
itEgnLCYJLAIgobjYc6v9+O09AnGhSrSB7GObHqnwS1YLHU9QimgaBbfIt6BxpN5
vLVpd1QuN1byR0dMFZYA3KkdA84F9tA2yD7pozqRlC6vDtPWLi6Iai+5SWPeRlMp
KydEwgMNmA/fPlbBX4lrsiAES69tdn1WiP1CnA6Vpcd3P7ThmcF6Lio0rdC/vaH+
UE4CQa7arbvtg8CvEoW1SfFYObhDZqlIXUelSj8qnseVUWgJ7+/4FTkq+q+wUL3X
nwqSgbbBxicWK/DPKgrfquOY3ERntctRmr/wrkTn5QTZ+fhQ+OcE0H0bkTZzErl7
bvqB7aJCCq1ZYGV1NwgTnmbwRbcv11WL1pCkp97ljLckhl+4K7kakpNyf2ryhvzr
QbZ2kfGAl456UQn/n5WA+7pRgYs/97PwrDobuuxkVe4XSceN0cneSbFeJX5SKp/r
dhJc3cAIsc/AcE3uL9U4QaFcEIw4ytIBf7650VuZi6OPvtyKL0c6h2sDTDGvK2Ss
eljJEPFLgfxnXmYMA2gZNSDWoz4tovxaXeKHbWXtCsRYj8Vto6a+lubMEeZu2sI4
VDsDt9p4ceyJfBTRc92zipuk4iuDqcBBIQbpS1eteizafrYSC0f6y7TU4Qv3sRCn
FOysnN+7DwU2/7X/iEcOrK0zzLC0dvfKOA2KKxWqhlr6aoO7IW8bgUh9YLRSRd7K
HUIdg//7ZMJPKg/IM+eZXuCz03j1rs1zYZvqNSqx9eTo5DsNdInTNlYYnzkqajj/
0ubJV2jv9x87pabx/kAhnI+nBD/POLMN3oXd7nhxCZhny340Rxd2aXIzkyzGQ28y
q5eLwka6d9+/JtijIQlpg8tzRsCARjp7uY0EXX4OFVvWT40ypbKjYgzEtZ8DCVlm
L/dTJ3ACbiz500sBSVxhevYHRzmf+ajj4Mp1dg9/4QGRpbxsb/X2tPgoi1DS/6Jt
MX+Iq3JfGMSbcPxfjpz93zN5OqkPRxFtDBXZtL0AQuJi+vNe/yLgSEnoIpaLdIku
twyjSY+Lej7unIfp3OMqyqIiB2sTS2dIp7XmraC70uB8t+Qt8PFWaIO/wP+6hCFJ
EIRCtuH3rmJxdxP2/HZ9q9T0Gzfsfi3nWf7MZuigqz9uxgpnFiCtRgJBYbFQG5WT
F7meT3fmERPO+G2Wp4YQsaT0cgYJO5mZcbbGTwCTuvefLnNT25wZ1aI2f7n2oa8V
zNVllo+OikCpcygt+yQWDLAR6fTF6eeqVgwaoV8qxg64q3ZBuyFam6hbX6lk9HHO
0/zDeSA7XYLpCKGkF/ygV1CZJtSHWLBiCsbhlPP2ImE7K6kyc9YbqVhHmDcdUkVo
EGOsUsVos+z4EyzPGCJ20qlYNo6mHrYF7txLrCXCUU1stTI7SlCYk364WV7j5E+2
TRV8l6JPoAg+gRSmIp+nZfFFo2TIPI0SDGplmarG4C8GxSfH6yxvX793Ei6nrlKE
qDwhtOJadsHNnUXAjO+AViA+xCWFNptETx07dTLRnXMSszPMAvNSBySqXJfYiykB
DmOH0AfOiP7F1B9sxFb4DrcO+caguNSLyhDvL8RtFx1Gt3Xb/AZnLTa7t6lwx9VA
6iv5ojBRbG4dw3//Ch8LdcA8YjGfZIUNja/1tiHaEDroVKrzwuPoJUzxIl9HmYha
uSBXLLwpe+Oi/zZIk0oHGDdqKwjO8ywPHJf+Jhy3mFQMkysrRe9MZ0gNkJFCL5Gl
12BLcRjGGq3G6HDSOHZwocQEDhs90gnmsIx4NYDD+raTsdYXajH1DlSUsSwiKHNA
zvirKZvuzDO6phWD3uLf8f+QZneV3cgVBbgZTIIiScL387jYo4pazWKtHq/NRXWj
3O3NEi8/P3W9FfOFKPqbwB5/L5Xsxz+Pz0z9cnbdXq9DHkNEy8OmMq8nyiL8k9Tx
sVZivBLWgJVlIIxPeei2jSTOLzyn8jf0e/9rU31tYUnJw52lzmGIlu52zppN6oBF
3oDmkKSP8GUjVF5Dy43EBe0gk4qWGMiyuMbb7Qoy3LEo2A0jNPDF9fTF3WWVIKqA
SQfwflLUiO1E+YDjvxujCHrxa1NZMfv2GzSoPFxfD5SpCs90bFlHKRS7SYj+2FK2
BgAz3NE2D53KBLYE99wDeGV6P7Zi+6s9OUYucFMkXCshhBdyQ8uFkViZPGabB/Jh
bt/Qe/Bhv/D3VkG2+Wt52M6ww9e0L7MSo0Z3DIWMyqrrQRHSReu61OIs3Z4AGP+7
0GEnZ/SBGiqgB+dg6lgHUI+FPjA17lp6wWtitFARcslC1PQVJw749qWLhiLiit7o
LCqwbsP9EmHq3NUh/bmh3V3tBiSTxF28UkZvTBjfw3JDx8wKFkKqyQQgT7d8q8jB
Rq3X+AmcAWuEH32/uRwxVq4+32cQyjp6768fKEjXGPymw4Pgrs5RzXEUtiTqG0qM
fZUNyxMfvXDSvGar0CU+4jV2htzauc5OMbj+xG4lKmi2Iphlp3D5qM17Ro1BWnNq
6qOVcQEp4reif6ruUuaIFdTfD4aLqSfUzhAeYkGy8oLsE5CnViIwEhkUt20xKsRl
jNJpIuMGwv4zcWbWXvv4tWj/w4+kM4DJ+dS8dMZWwBtZhuXqf9mXTTHIc83SymyQ
j2iF04DrjuA1cCYuMS/YvTvHQ1pCLlpOcf/2ZYd4Mc/6sgSHot/CFfvGhQpJaUAD
CZxBRJuIMoChXKDaVayN1fjOXEXcxbBk3DaXqrBI9pTthTlxSG4d8ToPt9gMnLos
hSNGNa+rBnib02Y6P77kVpt3FZPpGH/IIKKlk95hHnyw33zi/+wdAxHVjvXCA9Ex
BYgYZpofKfc17LQhbci0j6yfSTJCn14/wYxSqhfjBzuMKdZ7IriIhWfBr7DgFLm1
ycqLdcmJ4JesbHr1A4zygZvZtts80jOCkzObGSmS5++q6vEXc7gBylhwuVhBN7br
KT655rPQU06XqmcopjL1xeMl1oAudau0XktZm//jXVDQip/mr5lhpyFuQAZNY2cD
YkO2RsWF1pCrUuRUY2E5sw6wJlLYcJX+j6FnEvnM41tXhUAsLrhUVErDd7W9UuDK
7O6s70ke8wifLxu+o3decJTwDsmJi3yl0/x3vceWKYIriAGldGvscFKLPYGgceyM
27EWcHWuJ0Y9MquotbSfwil81txpvjzCrgRvVhho1kiP9vBAL4NEihN44OJOgRUc
TaMH9nqBdfL9hH58qh3CRBvOrk+evSlrkkim2PpukWNxSr1n1qK14dkgc3MiMGCt
+i7JMte2RXFTGfv94rFPYtsWv3dNyX1nNPJmvS8exxAhN3SNbszP45hO4ezDXJlw
U8ohhdhTOOY+CakHDpcBKiL2xHqINbxRGg4DyAVDqPUkIvNwO6lv3Huh115KXLQN
BamdpgFRi3FTjW1CIciBQD0MF7CRsRtuIUjEqvJjhuOZR8CxQeUp5iWSlcJo27mA
6Q2toUVE8WDut6Ic8GHTo8BaPcMnK2E4hAZb5BTAfqkFoajcAFi8dehQVJP0X7aF
jEyJMwCDPAlKk1/8ySmj6RuBDpfxnmBZ0xDg8KyoPbHU/kbGMNr1UYwKogkcAYbI
wbak37VfuPb0pHD2P4aouc8Iv6lSSdMtks/PLVMuiQvK8MFGxjFKhqvaO9ylPfU6
Ckoqongl2Kj21eTk3UCorJCN0UM7yzSXa9OhGxaKSlMOknyK2BT0a+bNopIG669I
tdPjn4y7IrcU3dR4NsXlJZKga42Ofu1QepTDod/rC9Ze1l+zwN58C4DKO4uAj771
m0SBE/X2ng13pkw/qL0yutwpYOv2rc6vRjJNf2tot/TbHWcXHBXyglLpkvBTrFE5
mL2T4AZNnlbxHtTTGRS5t+JKm5ZTVRFL7Y0onLldfxeA8VyQrpEgVn2+kLxwCfos
D7f4HzDX23yHBgf0rBhMOgdDqJvAxA8pt8YuqvkAwiCbsBdiYKypZMeJQvXYOxyX
Mirwxo5PRvvwiEksOTXPNBbbjauK5HOuS+Yiz+m7Y3S5KxA1z4JmtDD6Zfi8lkJD
lzcjkczcacBGmiUDTADO2B7I+Tug9yaZos/vavVuriCBaDsjhpF2eIrB5oWHq+YK
isGWWrUkZZBnXvnLyx9svEpTerWJ+qfLDyDyo60dVEVwHP3KfU3cnP8gxSxajqOm
6TV4lfTrP6cxBr40Not0tPh/WhIPqjFVFUPWggZVg528pbzNmGP5POj6d145ZyHj
7vMhsf/S/HtvKhZM43uU6RGkhoEYrrZ1Ofz5vtIXiBkq9vkMpqPnD2M02hAXeGmj
6249/q6WkQB2RfG6HAiVpXm3RuzKbWUM5zmC/02xH9ic66EWvhe5R5UppCc4vvAi
HqKaqmD15rNsdL/ByUl7/gDDm52qnjsxPosULVY7Ad0qwKZSf9qPNot9/TUFnvwf
5u1U7WVbL95ng+Xz/QSpaq4WNeBNeOzLbls3xRoSB+KX7QaEvefHw4OKQt+qt4/c
GnxnGuJA5SnaAXDDnizGEuVsapdhZIDcYtzfMzopi/VzB8PfZDWog3YQQf83wya6
D1KR9ahdg4KRscs+gFk8tHetpq7FZ7cvpCiSYi9It+HsFVeBptBYCWqN/Tz/qrUW
H7WVSGsZgVEBgGS7jmdF5rH/TNMd5iCtN380BKgH9komvAlsR2aVxLZ4Pzy2IFhT
TjhHUgO0xfH4BXVul1+hZllYZGglp/wIlZSIHn5utf/zcDlGRp3XBOeJygYo+96z
7Avo7ZeeXXEMV9wxpiFaB0idfJdewxQzKE/RCTbGve5L+lQ5pRn/T6hA236W1RcR
cnubsokDUpRw5Qgc7neFXAYrtxyZ5EHkzEO7k4DXN5N7kU8ULKPYgpkU8dYi37AX
ah7aFdxcx8bN0YUEXdKdQVIDoL3WbQcqZpb4lQ9T47Flfiwrq2u4d2ue6bScQ4UJ
24cQSD/bhNMDGPCdkM7EjOrwUh0KXWvjRWB9Lrh5r/LAABhuEnKssK1Vkk0kXuTJ
iQHKeScZmwMRyQcprWppxs0DSBWXA/TtdQF3FTNXhgpT3bV9vNPAaKIQ8ZQBu4++
JRFXExfcrtDLzf6GipVLyU5LD4iFaPtFu0So+zHb4VTt+9dqXvVxXBbL3nIs+0y1
w8armp5P+0tubW2JIZ7ZmkEJBv+ezDqwXkUcfYmXKm3CsCHT2s8bWbwTh67U3kyy
D/q7M+0+Vx2cG6xkI7ajiMrETh2kHoF2hNE6BZDJ+wZKhUDB9FxH+glJWDVverpf
zATmFJS1XqPYnHLXLXEICcLVRjGv2US9W+cSomhY3hZI0trtex93QPnVA8mq8v3C
W4cav5dIvuF147urRdPUG1t9ryxqaChWt23Dul9MBYYMWj9kI5WDjNluTA+wDiXV
howV9HDDshOL+Ctack/pofgPVm1KxstWMKZI9qU8iVfBMaFWfGr/X3/AyLofD1YU
KTE7/58q2eAbKMdiV8e5XvKCzh7XOawvQqdHOkWene8GFgeGZTBR1gHKWMd/VtNi
UxUbWTmgJVGqWMrT94nM0SVuiqqL6D3Hoj/xPknBFBgn+GSFNfCNnb1+GtkLU49n
m3P0Ge4+MnT7BH70h5392brrYSXpVr9UPjQz5MU0NHXIlWPse3NxpEF0/B55IYQL
zd8faC05nX7TwBPZ3EG21Crvp4kvP9eNwrRjjiVDUbmaSyN6sE+qx7cMEr0g/Kb/
disbtB2rHXqr3tOJD5VAHUXO//fdA8reLdiwslhNyX+TtB3BzmFI4fFp1Zl7otvj
HgTQa62GvzLwktwXcuC5Cl6rf9TWOcH1L5dRtIkGz83OZuf6ocWGyy/Oaz36wdw2
aRT6j6mhKb00LvhiEIfbBcKHwE3Xo8HnTT2aonUIMKHt0uJo3UhGwfw2m+SEIgXC
ltgs/yrjYxlNzT4xxNiBeL87PAEZ/YynOFcS71qRCMNxFzXg//K9bzbQ4Jo4VD1e
gy8Jf8YLgK7PrvNHceI98w7TNHs4p0sZHUPHRBBSCLb9HppIKRjia47L4vwyCBYR
kHMEjL9zQSe0PZNvLIS98dp5/vRsVHiQb04/U1w7HtrxWkLGApcpdYi9ncnSud6m
FcANSXsA1GXdhdRoi88BlMmeOAoFBJB3XVYuFR+NV7XiFihWQ6DLPoMNsxAAp2Qn
8toRoSJXd8goxMqmTBc1dNakIADKZXxepvN28+cXwgnub21sRxl7pSpPKtT2KqKx
d/eYvk9exXPVPn/xv5PEHsTuOw2Jy77U70pML2BD48OyQuGxx13fByhvL/CjRtlU
Mx6WRrk14kYbetLC18iI6s3ykETdvNbvhm6QuPRNIjANMM1O4qb/VW+VDTLMcZRp
YGVGZJ1RSwnrC1eK4ZBZDKon+F+aToaRYKwdbmvYKr1d5TPoHhXqHL91akrDHfOw
+H1JNg4T83Ef8fdEBa8H2be3I5DviXpV9hrNnWFdlQi7+ZAWdY+ijOq+oyViv/Yj
GnVW1TMENjZtS3OrV/bUEr8ZHEGXoloDyrYYSIzo6LFL5E7032WxEd1V5gbHwqoO
V+CKeg4uxVcF2t+0J2KFBSxA9ovz7nTPFuObVXzt0mLbWYs3Iklz08yeWBX4KFjd
n+dIWlBA9xk4wnbBL8J1/RKldsI9TnORB3JrBfo3UPWnD8AJF6iyAVBkSXtqOUS2
pfQrFcNHhPkwdrsg4hW3ci1OexiD1oRg79Yoi1ONYQaRmceajQBWFX+OEXjOLZPf
y2ipNyHIpbukC6cfxoiGYkd94UXPFCG+SGGIay82Ztd/3/yDr9/mXWOf8wtlMbqs
FMwZEcZRlAMJi3lmzGogQsjxsNo0+wDzxIpFiQ0Kp0j+IkoNUhFSMvVmUfic6eIq
Ho1TAZmZnuAOcvtVRTR1Kd6po0XnMkXSarFr3FKAx6cqvPdITJaUD/8yhxLDmxev
JejPKS4hIbgWMV7Kq86Nrzb46bz0XIBZzYZfvr3Faccufi1WAR4mpNKPc5AHLUvX
qQqN7B3YgGkVYmCEX1bcaV5WiUXkz8SXu2e6uegh6FslOYBnw6kvlytsfM1z6lDM
h3jSpZmNez/YGAoDDfuzjpUm8VE2B9NWk6SnkpZCnBCmfP/xWTXPcfgKkMIjEnNs
Bzp66DMpWCpebjtN/7tiiIFBdCj//JjfUYyQju4HAB3VTu5Y7EA6gChBpCseKANx
FmBmusnwtzQZKAfuatMK0J0YQL2NGscfNzpOFAa4svTl1JF2/R61X6hSsvBVk7I6
xZAYwN+cuJFNXcBT9O6k4YiVAXn1PDjNTIEg6V7nnOiP132D5vM08mnBaUPiYk7T
fft22CtTjxlPY6wkzMx8YUEKJ4KLhvWINMqmpUWJcVLOWNq8ht78HHxg2psO4VFj
u8SNhGvRi22oUVXo5jqKCg6Z2KWasflGWcvO1o7BeKuE4E7RGL+KhYkajSwQBTFp
L+EDLtne/LDHtH1NU+bUfNGqnN7pdMRSXam+yxg4Xx/DMhmU4imBhxPHMW8yKaPC
uWjf1kOXNdK+UaAaWWYpgp9HReErJI9wnx5prW8pqTRfZPi5zwKaessK0z97ZdrY
5vJVgsrqlaIMEl40BcmxWqyDqceBg275JfX46IEfZJ6bAKnHQNukwhD5hV3PSz35
pdl6P+uljDYI57vZ755JrSVCuT4o3bbDBYJ2dkdLf2DNmbMVnitVPey/Bh+T/wjV
1+zsqHZErIM7Vti/tKsm7L4wZCSwKU2iPctqwLqfEng6B0pyh5+b4Kztv+0/3Piw
Pu/kGCONZMnoP/LP4Onne/Ix/FTHwP35gVcOWD9lIa2IB1Y5lAolLjm8BMhbWfd2
UCQzc6WrFHBze+FlmBkAcoR174G5Ugdwd20TwjeKyYXHM2FkkNBgExpvrAAB4DrJ
AiGUJiXm0kR3vArBqKbMUmQPCxjfW+H5tOjzewxC/U9khR/OQXbV74iUM7SKa7DH
i+mVRqW/2FzSY/mzgRDNLaXw+Fe8u3NsicH+yyZE4SnIq2qLGuhofSbbgpYuJ7gx
5XGtAYNKpMFzyG1Cg/ltYEBXuaARKY1DcWMiv4y+j2rFgjnE1m1riiG32qdNVneM
g1klQGOsXLimQreMZXgbD3YACXY9npB5cHGcb5yOLYCGtkarQS2ba7LfOKtjkV19
pKxsnWdK1CnTq9gopB7w6DIyVXgNspsX+yq3n+JeiJ4jV9AcMWqrkaGM1L4gEdcO
b0/YAcrwIpvUu4gNFy4X7kX1k8MhDqDggnoyA836aSp6ew4OzuEp0wF/GZGc+oum
b0P5Ha00iZMlmwRpdRBg9YzHRPPj8oiL4imDPtaBNqCb03ETNZvwQq+NA7st02wT
Bqhofep9rLryU2ktfrCTWLBSsOPk7JIwPejIYq6GzOszrKXaoS2xH660M1MNXUA2
M8g5VERah6Zsy+KJ9UXDeABCmPp9d/4r4AsN0oT2uqGS8L7KNADTQym9z9kpwcAg
cntl3LqIZiNZV+Yk/PtIADX8OdT/N8Q4afjju5hy8lqgPLvvUcIg6YDukm2KR4hl
q6loPo3BQy7pduG9DCZh0nLulEK+rKe+kwoUcxjlKv2h/MPE2TJKRVfs06o3Suek
BE+Wn7qMHujW9K/L2z2yk0e/5G5yP7W88Okw6Gk1RDVyG4GiuLeql+wMseTJSsBI
1DDdFWTJ0GmoTZUBZQ7R2RarY7XWBU7LRdeFCZsC5NRlJNjvulpJ4WbLDO8F5TJf
+uj8pyRXDA7zcc6yKbDjdXI5A5sHTXDIWDVTQ1x9mhVU8cwnw4dLy3UoienUiFpr
KVXLo0AZWxLzXAuATOoKoV3KE8Z0AJoM7jLCmMId+voUvl+OsyJHyztZMCB1Yz+b
1Jl/ail9bJ4hrQ044YFVs9T/vCU1KE7MdNBvpK7FKAvS9zMXHFezcItJHXcNtwZD
OjXtPf2sCV9NZruZtIkdznvJhaypAbwM/+4keNiBsHY7k0WtoMqKutpSDtiTxmyJ
RXEW3VRXRivZgTD49sz86gipUoXeXw7kM4lZzWg7Bxr9NQEjFxKximutS+u4T456
rfeT+CyHY//JdJ9SPkJ+pHVPX0jzrVjm74myORCJ+SDTayLkeoHhtvUTZI9v2Oja
w4mFjPYLgKokttrMXR/+pgWc9q4NIcID1zzLBmlaijMeEn1kARlHvsk6wzKsZSx6
FUwnxt4JM1z6pM9BKkhtV5rOIFB1x9hVANrxfCeCFMowoi6xflPfsvOWkdvGyy0H
6VyoVKfYMtaa5a3WmT/0YY1yLZ2VKgH3qrUEZTIj0RpEb0w8X1Sc6p69zloy+Dm2
4tq15JTwUoc20u/1bzcT7HRCmhImKx/UPB8BX0x4krfUGqQ7rZV/vtMmRPsq5SIw
bFbezrW7jukIvEa2oBdlBQlnePCFdWypwgBNnaGfYiqMbECfDPQAWnn44yQCJg5t
WPCYKP7tbIik0QzfoG+V3/0Ko6yRnOc4DuhpEJoLuiWpbfBAisc24VqALHtY6X6F
3OkbHDXiKtkUY0s60kjJMK5rrPW1SMDxvBYMlkBkpc4MKevknWN3+orbCJDF9jWx
PIZAPiHfnXjeCWtBrdyXKolNqu+Hnq/W7kooJCkRo06Q9An1e1Hxc8IRfqgJUYNp
L8IS7PEsyX7TJsMZRgjSsGaa8RxbRj28gkL31VTvyPG53gPPSe0WmfjivRgdNNge
eS7i1mOuZPD/zeD2QDLpZOMY6nOVa8hRqj3NVvpGQOnpWhmWP9E8cjGNIbSFgXkq
QKpLVuBDtPdDPIKDU1584LunP2AMgX58gqBbZLnOLe0XSJhTUW4wgQygRzEo4Zsn
C9IJ3eKbJtVgVkNWXjBTOvLXlP6gCUbuDD9824MCrIsUqVidfpdZJFFv9tLO4m86
IYZP3vVnRE3hTCWgBYexFKCJjgjoqOh2RxYwhUonpZLNbMujexFUlUGI9XQ5KF0e
Ls3mI7oeXo4LAW6zR6OzLeqEVhOraN/Q6YinoGbKuVqnWD2JPrXye0PisHH/xjvr
HxE5aUfFIj6B2gaVJEMbupL+doohqwMrbZT/UmkYkt9hKyw8NpMHiGDiGrBR7ODu
rl3onvwSriv0ZgkgwPu57DMhhPhIh3/3qHZr4S4KSUSS1e52G1OlHu3A499PntSd
Js4Olrsc+XgGez80CmqlA4FDhbpP3PY3vlNU2SNcC7yLCK3wQZGVHebUUHzx1zOw
/SiigQcogG6CrSxrSJb7ce/kxxjnmHvsu9FMXMZIeOpxU4Xi2OeP/eu1D83bRCPc
3VGOPRoSYdM39EZ4Yj7MPJQBWf3pwuxSP2kAKBg31xIsEwPXI6asudVlBCK1F8/6
B21hx6kiJPAWRZPHT3JliwAgZ0E8/7QpzVC9dI29bTV/xKlUlPhye6PfGU/5KgDh
wTsAXOQZCt6p1HAO75jmSwOv3oyI50da48ojYTqUCnymtSp/QCtTypIQ3Ve1DR0R
C37uV7QzYivO5+RmMZDImpdeNL57osccmU8sQqsvEWAPUM0OmqGGxDJO3rhVboIF
Gmxy5FtG1zwVIciJwt+IJ/yumioBXeKpQpXlM8OTxmE9GP2JKNXA9BlsSn2T3jMS
lDlt5DwKV5WCsaci5qRMCHahtdSRw446T3g/pIy4t5txDtEuChDgwOc7FQe/g6aQ
OGARdvCvF5veutnyv3DPTah/uw/z6bklCxSkOju58PxDF1CJo1NMrfkZDNyufa0K
TGdZngvF6WwawwoNRFz+R+GwzGnX2m5M26qKKskTmXDKLO1ibCD5oWIFXcWPEQrk
mCyHvWPD2ltfk4Q2C9wVCLge6nyh3kenm0q3D1HNjlPdl5I437r3iYFNlVPa/jyV
1cL75Jq6oBbpmUzTNz9dljFdBx9ZnMKCU7npsaq42NBUUZHbYmZpWglZcBvLG5Nd
1esjMcPGIcTdA5poaiV1fZ0SwjhLYP7VKkkObBLGBtZJq93s9sx3T60+60I9tyhp
DlMOWX6HFBVRtcIUXm2hJqrqoPLcbiRejl6O6oNO9QnS3ri4L9yk5sslAmzY5x8D
yFTOatowk9645A600QhFQ+PVO1jPh88nYbynRuHVRWMvNNqCNlBqNQhT0sApIx6f
zF56y8B8Gs9fPWBX+ShOXOi2b7AMK/M5wBqXfbUecHUD3AL0y5pBHsG8UzKN11m6
MAQpORB9GHzRmJd9oP4mdt4nwglmF16HsGPUciN28Y3O6ytHo7rYK4TkL6pXdzRO
pRpLW/UF7ATOxUXLeEP5ghLF/Jn61d25xHfkSRzNwy8w3OyHIvtX1b/A1m7tFZO9
7pKJqjbpc4RSiwLlQE7AwGTizK56Ml3MSMKjA2HU/JnMxtAa5X+p4Gf17oZXjyQZ
IYWgA9hz9H+qZSpLe6C8D5q/X7Y6y+zQ9towjRbwttMdrczyDd7JpbOZqTXqS7il
ml+iE9z8px0/n1yJ0tm4pZUcbeqpm6ayIiQUawyr6+fh3XAvwqJfNmNwU3QSRrX+
z7HAA5Yg53dBLUk8YrzqnIVedhxkiiU4pGeWCmSwef2dxBFmNMPODP+qW7rKX+ND
tNXummHpoCrxTJn+joExLJeZiX109D78NmKvwRFXvMfMvVPGmGQ08/PFEkIIQ6gH
uPIVEc/hmmOUDmw8UA9xTS/J2Sh5fi9AIW6fljXz7yYn8s1+QEaIcpyc/Z66gea6
C84qK2D1F1GK3qYS7lzdZdITEoeORrHvhisaKYVNqBfxSXRDrbPSB1lPnz+Febsx
GunDEHP7aHPcZWJV+QhGojoo6mQVVfhOuUJMRyNFOq3Cwwwm9JUAuF2lrAA2/ivd
kuRGvWTFpLz2jZkEowKcWlF4vkG1eWYG+M7DaoVXWOxLqBUvO2y9ckm4qH0qZ85X
fCpV8acjcfWkH9nUMjDlePkcITiU/nhjI/gvxqG5aGLSDDDUXrMiOoXoo13ObXeO
EnNxgW/7fcWhnDZLxAwlhz6H2i/k8vVFm4Iijma68g9PiGq4DS9DUEXXc5kO/CJn
PsTupp8d37Kw9lNrMkHCzqkGm2KOTQgKYzg6Sym293RvEf/62b3KOOxg/P8peIic
6k5AiXFNKouYGBHrd08z4FdLJkR6okSvkO4a6BsJFoFkaDvH5xA8ZgZ9fdheIsRh
ZogWzPqaF6G8Rfq2dwPBmYaENxsufzDaSqhsP1km5XXB7TMMvB0olsW10bAguIVo
mv/ScswQ25uBFH+XwgqdAq0BwPyFC4aLaItDRV0p7vC5qdIAUdIYviqBTp0ljJCo
I0N2oovKX8gew9UT/BwBdaYi9KHE/Nt6t3sHEI46nUf+lCMG+y869Auoq9N4JQGr
b3BpzMRQLVeKOIUYO80UIW83+52XTVxORR9FpA1feJUjv/F06PlzXZB8ZB3Ib81f
gvmHtmIgnxMQTIWSKW6aul/KWWmfvOYA2BF4sI9GmNzRdUsJg9FOj7sCqYfO/nBB
vyuk7UByQHODqdXBnkEXOtl32nwi82lFLXyvSlmWhXbW06POYadLJW1aHT4Noym0
/g/VOUa2QLi3cXVA7PpNPS+KDGAQPShXsOEWK0RhGdUgx0shCVT8wog3GxqKQVJI
kQkVKihYUrnHTehwYH0MXKfz6DCz6rcQJhfvcmammdhxfdQZLZnCq9kYVpBnJotF
TwEK6JqMDscHyiou/0t4X5JwV79CSPgMYwYhnU/JrU7jZXXvadByc/NRawpODKH1
c1CNs1S2ns1ehVGfPhXPeKQVrevFq6wmG1q8nnO545MLVLqZKmicS+duzjDWUu3l
jYj2jw3IY6HaNpH1djWqipQTioGw5fzYgoPcuj+h0e185st8BaRplt78BYG2mn9E
HVQgN16VResrk01AwOnjaMdZgloY4/zAXqriMhQWjZA7yNIod+u4UEcN0nskz02G
AFUadPvKrG4aMIPKIX918osF4HrXQDDxz/IZQ9/ZH98xNQl4k0oLpYDImswgENPz
i/t52c2WIhq17nidVePFjI5t67Z8nlatloi2XQS24WgGR6+wYTxO5uuiic0yXHNC
oAXCvwmzFf19jmxcoXzrd2QicgzTEPwWcCzKquMNInpYAw0Mm2Q7Mxxsf2bd8WJU
2z9xMSfZcIZjl+PSQyq76effrP9kI/1xo5hUYFSqbWmcBRIlwKjnAdhDLgi211je
jGtBlyJwqRJYNVKVuV+wN+QPY0DymKA88qqU4x00A1sxEyfuCGOI14O59rXTI9Xc
eqAXCde+920anGi3m7jZT3/70M56wQDyyxXjTelp93nTpx62Sblfn7cdS94hteHB
fmYCcjzYEAZQoi2R20rbObF+gFLYoeHbhyUHtV5BsV9LFWGs+n0UBfM4WJP9I9Yc
bqMV43uaQCIQFDOelxZcS1iLP0ut6qivtnAWLxi7IwLiVg9aoEHXxeHn95CqEXOW
5g6HxVzxJkiUCNhe2m77CICbpeVh4zkDYnhD0cotJ6LPo1GqDRKw74VEnKwZxx9D
Dwc4iF6hM4AU9FMb+ckJv8UGic8a2dLmEqtd4I7IzRwv86gu//X8GQJxNzC6u2kc
3jJewG2kzaWm+QqgD0ADgswViUf18p3YcEg0RNwi73EITHTkAxDNNsvre3EH88PW
8Vm1A0wfqFmhiDZxEZYD+O5AM1cqh1Oa6xW+aWpgSO59LhtslIfbTasbno5edAhT
5neLQYUouwBAlffCVakEKzJG7Ha6Jd8pdIlCvDzSyccAGAk6DysOGYW8l9ltRZjt
iQiHM+xmx00iafPC08NThDkLyEI+bLiVyb3IH+vwESfOZR8ke2X3TKOTjL+YvDPr
pPNc6T4JY7asvTIqGwvi7E5c6HsBJMsA9IS2VIt5MW3DfRA3wXBUfsxh2IDwbPDw
e3nFCbIsOHnazuTHTiBE3JrgiA3IQ2GbWzDPBqkq9i0ZZQypc7QMyC2JCYsVSpyQ
HDJ/yHZX6L74N9ZnUs/d6a8MSp+H8e3tZ9+ygnkW7bxK0uU0PRBfZCUSmwy+Jwo7
/yLtF2f9PZDz9z/2sq/J3oGlJyHCOrSQJrvk1F+xhkSQOH7RfF0GOXNCXywnhGt8
3GgJM/Ug8Lx8vNlcJUg5ioehnaAUuHoUhl+7W4I1rF5OyVxmAakINfVeRsg2wgGA
h9vHYyf+oDyfNTFNDHj69Ymd1Ok0h8XWBOkgOy9Gh2f97xZ6rc8fIdy7KeuceITP
DzD+eYubGJRfvxCbD4ZNZi/9SOR4HQ5UOIZBw2H+34LXYd9KnWNqfiizcc8i1Ueo
qJa3Ej+ater0GzqUiorkI5nNFyQXEdKfa81FycI1umLhGksGrHPJDDp8fOF9EsM7
LR4kqADtHsxDsi+XbHUUfL56LSqmeSQmz5DBqBRFnzSaMOQ3cKAXF9IBYAmunlE9
C7S0KjD9ITf3RSneQi6Nl8SQ3lHpfPUD83Dl/P7gcEG2Hd0Bb/gxeJdC4BHotgyM
WiPtNywNpe3Yrgz05O6qP2FQJxTgp2xdHa9Ghzd6wl5O7HewmJA2rrTHrU7fkajs
fuS8DSf4NMEbXMhWfGDvN9jxsBECB7H2tzGzHyopUALdP7vR2NzpqI4AfC1Z2B+L
4A8IHmnQzCrRGRtmWxX2YG0QlLlytvhr5dzi3JR2v9OXQO5392ZgMIXTCJiOlAGv
lN4mJXa716jj/UPtA7N+ehssPLAShIf6dMZqnnsrv2RJ0nZMXFhddlFN5U3Fb5V/
wPSgUUSQ9rlUAv3obxURGvEPKOXhtCGkeaFfES52j0E3G2dbIMre7NLTGPx8K/4i
XoPkJWCVqo1JRCz/f75JPBEFXX7mnfm/l4rzakZ02iqPcCbKzNiguToERcXgeN6g
45NN047mOjR8kJ7UG7uRN+KVzmGWXiNprwUOzkpjtfOAqKnN+mLKMpo5c1TWOy56
YC2ePNKfvPRQco2yriQz3oJXHnAijoynq68Lb4uLZqLwE+zS1VC73xa8+PfInwOK
67isVqB31B5sRWR+TqaKk1lRoeSVF6mSVXwqUbHHV5pQ31CPKE47ZIUbZE0kYv3x
mQzkStRAPLYMSNuphkhVJUgaouMNRCeFjut8/jfliNwqkSbE0cRJI4zj20+ndwjr
DJMdkzo2ZG1xef67jjI5gj0ZoeBDjzdTTadd8EQ1VkvaBdck5FHiH8a8+oKIXcRJ
LtAbLBcS8tXznrljaINn0/VlUh42AaV8yzB2vEqOdHQdcVYqDASmAjJfCCknUE8M
RxVZyBKTvtlHJCZAk+eUX5jDOdNvg+DD3oU+DdH13TE26Hw7JCROJiYCqv/pYILw
jBJkuUHjLANltiOntQRzFVLLRdIgfzY05ivZ4gkyrp/UVL8mbldfiocbuQ0BAVd+
rNvObyFAT4OO4BcJCWUGODQradGlzfnfggpz4LDaY//Fw8Ooqh9/7vb9QiWoBK3d
sXpK6TNvBssmDY3SXr+WjMj22LKRL6+Z8N1+ksvSC9Y5L3EdZNMzlKuzjmXQ9DZ4
W4tR3qbyfWepTqvFEPd9WM5Rw4XAiUVEfbJuzIBESC1dh48U+KxpTB61rRH4Ax9+
KG7PQVy2HuhfgOuJPnSKGFnB9Z2B1+N5X2wfsuLqKeArdAwGCbWLWwlyAuqWF3i3
vpbkj7EsiVh0zQfZK4t9hG1iGjjVj4SWX8z9cnPBBo1RZme1CfecD8RAR7P13hXd
5zmi8hNAoJPXK64gN3Xv+D31FJE+Jv043YgdZnKbtu/LlPHPqmka366/DWNOCziU
IICBxbhI1QD42fqZhN8IEsCHmbx1VIg6MMsq5ml1/3LHq92WLu0wBn74ZU2wWwx4
ofe3vbA/WlRP67TdySRggjEQLEVWfkWaPtJIHsYFOu2DwslG19kpFPHu9G04M5Ke
C1Cy3d+TKnbW7OwPCqohkip+pF7e3RyvWyKacGO8m7tIldYoEWMofuuWyvJm91EE
t4bxMUHIP5brVd1kiMNq8RRFeeAMUPf7BI90QA0+poZ0vKc52We2L/xQujoZvNM0
lQJftG9MS9+Ip+ZQHDYmforF7kPe9EA6HTEw+drlAJOYibSC5X4uk9moBjW6Hhyx
5TxjMNILikxSO8HOTIKP7JBxsakOkKNKsBiF8PkaW5TWIn3kBX5vCP4Mzl3rdDuA
8SGn3KDLSY+n9qBdZP43Rjc/Q7+/CwrhLomTQJMHySPUdj/zfD6zglRGeIUEpSh/
PIUp4jWHZpgcoA824qYzNu45suKh0exvudCqI8VNZoM+izQfVa0xV7yihdJTD7hj
XXRS5nE25ydcuM2DsXeSjjLFDPN1i995ESsV9jb5VQdqqRfFkn1pDYeUxTc7CAIZ
G08uyH6jJ4i1gNlHPR0X9C1WXuJi94IhZPS4ECdiyjK0x0+ImBMu55+jK7Vyhr4F
ghCY0kEgQmKlBtzVorxXcq8oBpE/yeI6WATXQOkfEr+6ZzBEOoU4H2WHh71Hq+yg
bCf4MaAuIsoryRz0iMHUSy3CYGXiopjG8xrR4AxLOD3uNnizSmw90kKyRCFxC5oQ
EiahUD9qzC7YAx/LVQc1FSjh7dZDusjRJg64VOGEHb04iDgLQf9LL2QRuszgAMTi
ByzKr+dOwo/+cvlez9xfzkx1IdT3incKdCpLVHPn3eb6A4C4BBppsFuVwxcKCc+1
E9mUxTWZBhImu9fU45lq4wy9h/pCdSyDOkCT8+1hNDkhw2ZzSJU2/j8CNXr1JghB
cqNDPqxfUc2NEZlw80a+6VyUtUogQ9O3nZt2I1GUb+6muNqShsr8sVvr0a4OVQFs
+OakzFIAE0dOm2yZaVWQwWP1eJMza6qE74k44lGMEo1uMtD0qoucCpanKBn3KBjL
h2sSbQzdzuPhKqNqx65u7pN46WvbC0PNUkA59wVxHDy+2/QXp+VJkWSmoJKLdaHm
kyMIN8w0BGz+AFvh02Oc5SCbjFHfqqHtIbbza66py8WGbKayCx+dNKOoN63hmldm
a/Oh6a1Ru9POi0TlnWd+RPQPWfaGbNyEecDtzetJFWZY931sWQB3P68hIYE/Gpx+
eGwc+ZB/ppeJWQmt1kcvRSjj29Xh0rS6bBehJanryf10SPONOuoFNAjrLDY3C3nJ
is5zcguKo4JseOAGSWmxZKGHhHrphv4qMuGFbJIucSaMO7A8Rn4QfxQ4VSv6X//X
3GRFqzCyjFmin5J6PeMd9SSOSmZgbuORVjQ4QltTQ9Qc30Bzkm7tNYy9bmw0xEBK
l5BJcyGVUVwZdxWivbdIjX8V/v1lc7YSfhj8Yo5bmupz7zCx/J9H46W9878A8tFg
zElMQjO1wVkCTybJf5rFRN+5l1SjS0sBe0NVLK84T0qM/a8RIaGRsU9Qbhr8CZSM
jCO+c7PaSwxrZJyiEAstlAK3lJDI31v8DGPdxKe4zR4WJX1QvYFBlysrnrHBOf5e
1kHjkBjWWvZoxg4farAWo3+/Kw/cFKnZhCN1zeTtt/aPpPyiglaA6rdYNJo6qCv7
kq4v60IkzJV3KgTtSDapAxqpl+MnYqKDymfOioGTtgmEbWvQd1yAcI07RfRDgTPV
aVNSMtw+oE2eeTLZUVPG8DTFiHE1WCHA8SMXyeH0kBiiab2+hnTzeiyGQ01KCjAl
CJ6nxS7qz76bv1t2TFvOd9cLGr9tbI9cowXggxZvdJBvBDG5i6WxZxEJg1fIBcz9
1441nrrlZM8zVOsbQqtMRyLcEwC2FJjJMH+Yk+jhjMzxJQuUcKlGumV59vPiO5uo
DnqsCuLGiykzyt1vGq8yeUWKALrXA8n0UzJm25IW3K7R2Su0Rbez9KRnCNivY7XT
KdC1HchgAZNRXScCxGcEN3fr42e78Drdys2DeQgKLxseClhhV6JeYjDq2Dge1tA1
m6hegIaeUhAF3YXM+tdlfOs/KO9BPoh9JAsukq+C4FWCvxg32cRhStjC77jdzAQw
OW/6equMAfPBtl5R1J+fzFAR7qq86708+ehPwcOOUDSE29p/wzW1nnPDoyW150l/
cWL9GJzOYcdSiH1tXEkNWk0hFSC4eFccuaZDV/e6tfkPGZyrQFYFOOOMeQL0OGyY
CI83L6+/cNeS3878aSJv7dZOs1O8z/YtsrO3GDyOS88a5MTl64kIm0tgE2+L34Rp
AcueN+/5/c/PrMHM+CouR/MiZx4egSf5Chjkz5yqCln3kqieylLQb0qCuIegTpF2
lTqrAHXGgp4gP7m3RDDHipnEFrwg6OFjZoBuhtp2tK0w6GlKinFUdt4CjwHD1H+a
vBbfifaQgLQq0a3AjwaC1q6r8Rl476Tmrc46G6gQSP2DYFbimAZu7C61aQpqyF+7
p44CgnlufwzsrFKWC0MMKqlVJF873gtpfWMM1QhrblUe0NPvhmdYPZ8lrHgBIA+Z
0Z+7SbUALN+V9SjG8CA4Id5BJbfji72VrWqJlVqXn/Hqtw9KznsWCWaeod6LfxHq
hVUgBdP6JspC2GXrqS9CCb7OpdoxKbZCgiIy4zoLZNLIcxgO5eAu99IwEBQW9GXT
19rWjydRH9m+n4iy6ktEEj0+3KkxRFPhcPyeqjnepxW/yZrmxWnI4HJIQNzxY2oo
wBfVsGDLZRerRHZxov+AfuVH0k/6MaNl+WucxSIfiz04g1VR/c8aUJoZiX/izHtK
XpmmXpQ3f0tWtSQgYXLTKfdLx44jLwfMGEMDnbu0EJRe/eTnMDHnEb2uybfPHVYE
fMoJQ7jUz8T80dUkRcO+YbBXKCW+xwpnhHUJOa0BAhod0xoQ66Aot6HPDDhLHVFK
lyI9jmt5un8sFZag5o5EjLruNAjH9G6BRAkeGw9CY3CZMAy8gR9K6RidQnGPxG9h
dcdQ9qEIFB4vpvCsvgb78OR2nrchcb1W1aMprMU8TQxAUNm3oYP3aousYPSYqb+l
JxWsIdMRN7tmjbxuC4z12bVw4IwdCcK558UxHgHLlb6lidwvI9MtWL+tcm28xsay
zDuzuKpT9lKjt6+QRs6G6+t87MjjGvWYr4TU8zZzf+NcfE3d8lRvb4h1q2Fuqcio
VwBjB+uIe3urbju06UzyxUjWUIWLbgF1vZmLJzvWgr2c7Wd/04kZ9xLtTIg3MbH3
8cs9WHWTygjZMZ9rKRBlSIO63um1GkU+NzDVwULw4QOtkXIUnSLtu3yS7+30oJ6S
P8MacezcDrPs7s8haESP/XzE3oPkPYfqCk3TVVCw9/mtQsLUr3OUOYJgvRRak2fD
cfkftcYxpZNCUuWXn/ucY+ttlsP7gMZMobwHGUt7lXyaWNMlo/aBVyfQeCq+xUDG
nTuAT8wKWS7lMiEVVy58ObiqbuIZVbliNDK3USX8hvpdP8SbCS/6mnu8+aNcAX2a
/TDbt25yAT3lvUNhMLW+qiF4+AIYV7iffgvjpfSJCvdNDNsn13utUArd1ErRPHKP
O2PBGfCnonWwwCzpYFYUlWwYKC73uiFhAji9oi26DjZAHqVqa3n0eBM6GDnbWSxR
01NbUl9IMbYQ9vr+GupJKo7YVROcGpbBol9XxHdd7wxQCvgq8qbfcTfxxOUuC7Oq
FUJy292vZWDrETxSr/dLxSSip96sIscpD8CMAO7hoFSrP9FBiclrRpk2ty9j3Rpz
pMuFj/605/eWHfGwpY4FXlNNrjq5ZKs4wjS3nARu9+kJjnFocm/iq2lcBWJUPjLp
Ot+cP0oKZOmePcq6CaQU2IEGuZQemrUEVHEbXY7xf00WNnF8KDFR/2JLOTd5Qu6c
syJeF7l86GzVJ28r1bRaQVt9gwXOgTJCbKyleg5N8tn9PCo1AOu8q1T5ZWZ0DpEE
icBcfebtU05sTi04NJk487azFzrCMcdj6w6RgV1v/QkJ1x67qwS8Hwp3uK0Y8cyA
OrRihLPkStEmOpKxC59kxiyg0eGL0qAcvhgkAbZYSqi8QY1e5WEC/uqTOuGeJH2t
GNLEpvb+LLz8NPYZKrN6oCpumbllVMm6sx05i27F5N/NS7p6+aWVX/6aEVSGoVRQ
0JUODUj8zvd9+CDiYCsMtvK++l8m/GgBEYBjJ/9qZ1w94KHG3CIGGNEedfMHa/Es
Uc1O6yJ0ridegdb5VSaY9hUau5wFoMtn7m8HTSI4AXjUrLoL0M71MIrB07Rtli6t
+iIAoOXTKRSEdFMJAD1cOUeApjjL5mGIdX+iC9uSi0srGUx05gJjVAZpAExZTv/U
Rwnw4z/DiScr0MVChKuxCAI4MreW6XHFip6lS+EiSK1q+WjncmO9Mn3J7aV7e9ff
Y3qv0/V6Ngc/ogXHJ/L4ovDaP7HGR2aqTEcGc9KZfJho+SeOa0RIF0f2utJFGOc9
wdzqHFgGs3fq/tUKIUYOR1skrqKdpLU5sHSgUV9VWmvPcusNvEWK1DoKV5XkfiPn
n3OaXrH3kC6c3sJAuAvG5i2Wl8AHJXcHeaaVMVIavpcqj/Ea0EkeqFnMhwE9I5AK
X6Ha19doXg++BbaHkQj2uNAGeISnC0E4ouhilmcHfO1jhKfXDXiMXFKCCf7KHyfy
dsGM97k11cE/dpn+AhxWzloXmQaa6GFlFhG00eJkQGMXS2xHHzY9hEJmWJUD8Rq+
G7m8RBXYzt9uk/flwMgkrY8rDZ5eJ8/ShfhZs71e972x9cj5482s5hpb3K4Ul9/0
hoRTczqoBviYVSojezmmZkwHxukdqZ9MqiHD6eAjLcmXGPwBdPH34OqYEl+s8RDR
BwHyp/zT8UnqDjIE+j03bKwSONkkqXt7MLXwWA7/gccU56x4ciMDh76ljPn/Bj0s
dwK75cazYtMA2hEnzEj6CSJ+Mhbem7iDN949LNYUxyRaM2NzWr7unfCj6trf7Go4
Sj6NvucNFwiHrArbYsfO+fYQ5bQSfIj+pAoHDqB5QnbHQ1cMMl8HoFYe2BnPQ1fW
mD2Ss7tbRT3HZczZRsZwpMeT2Yovu9rB06Ls+qs8N+4bEkL0YM5eqMOBAspKXhXA
caPGci1V+B6UmiYGJUMK8d3lV2Bu+cu9fMHaDQHJvD0jiiZtLFgN+8KgOiCESrwC
YcJZYXByM4tbRCrmozad4gfHVHuz9BJPsG7OPBmopQBT+MIknlRNnR4dFGaTyKMU
OmfdEjaR7BzociVg0LaVHhIl+K3RzGntWb07XTQamlZUPxTNye349vPXnMtStaWQ
O3GKX9mBJqm7xJRumNqv6UX2dV2cgCjbqC/xhh26HRuZAOZl0vk402bsBOdtrUT7
+6o5E8c51m0nv4myrhU2A+Zoq31sCXZ4nP5TL06c7cQV8eXUfhmxv1kJx76zZTWc
LI+ZoIBjuMycqUmfYq1Iy62+364lFCjxEq85layhB0+uSI9yVwjmPuM7zhiN69ro
`protect END_PROTECTED
