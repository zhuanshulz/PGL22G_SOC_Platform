`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/srX85zl2npBTAWDe/rcHfq2orL/NGXW3N5N+t9SgbLJICZ3Hsp/V/cCHU8Xv9dw
ihKGGNdhtc0qLFz3ayjimBdSJEl9v4lap3bOqzuVdA/X6xRUtGhWlaAaAHbzQ1Le
9ayvW1K+SKZg0uorAKJdncj6tAgvliDXdF3Lnvtv5t2iYyEpwXsHKKKBhl/uvqJk
ul/Ytav0pawXN9qNcdgNBTrBlnaF7VlKnqtHfs7QopdOkPAgveydySFa3joWlRna
9EAMBcCVOcAX0pwOYukx+lMC4J43144MD1PDZ91kmaQB9FAS2sGE3actOt86WOZT
zta6Eok3ui3OROPHbMkOJxsOf12jLYXYWL3R0UX+3Uv1MPPzDZjVPlB36unww66F
bzf6RgN94iO857ZH/LjEFCcmThkLApz/+sQ+BNDKN6bg3D5k2MXAF8SD59DqQVOX
SxNz3Dz69lgSLRjQY0WUOxGUxGT2e0E+n//5/dHbPXajPIy6dzLdNu7UPVm0l2fq
ZNgOLE3/9J9ZiJSsQ9fMUI5WlKDYEjm1GnQFHsGCfEKvAdJbJN6qUQzVtR9hQwja
j3TcVcJonLKeQ6d37N58VGsBPpFRI4GP4QYuWHbrewfG7+484idjKbqvJ/xgkrWD
kbmkJ5d/FEUakf1Rn1aOa0lRwgWVax+Lz8Ryssvr9AnTk6Kk6Lk7CWrc6pnCbpP3
DWzADmMC4tP3vay+kVs1dI4+8AMjXNEq9fZ3Eluv5QYdtGC7TvB7rivg7EI9AOJQ
HhluitGFaktgh2iHkTQn/j1IXF12d62jEnKCL52nG5m2qDcEWLpKOOUVSeGjAw0+
qBcxyPwUiI43hbx64wjaN8aJSIo/c6IFcVXCACy6+zFLDFIJg6CyZyy+oL/vqyge
Vd3b4nCeorEwalVZpaGOFe8GRc19FdZdx2I2wTeuEaA+IUXhQJR5qGf6uSd0Xbz4
0Bu/WZDGecGJrHlnrqbdpNgC6Bg0awg3SNAbxd4oaMUxdi9WqG4zbn+YOO7we+I1
DHgU34lggCWcNafC9+CatlWQlxLUMxdrS6oUMGwfSr0/eHZ8k6HifemsfXAoesN9
PwBWGIaL/2xpjpM/Mn7wWWRAhI9P8KkBBRr012yy6pmMOFuWj0+RFexnhFnIMpSg
RklQdDo0guA9ZvQ3HzRKF5tYeDq41q0OlWUya5G6pY9zcfeCedta+q7xvZkYX4It
KCEWF4+6zihJ2Kc2XUNyDCDERD3Foga1hZP1DIRis1Xa2OMhsAuV5kxaCu5ox9A5
IPJgU7Fofe0v5vE+FfQU2aYQ3jnt+jfUkN3ctft9H5akXqJ4vx+4DJ2ZPHZn2gaS
xZg6uvVUQakqBdndQjSX62Bf4ZhQx8OVgXdcFl3YbIO4jbe+DkcUOQrtZxtHZpYV
3m0PEkbSuiGeYWIecBHIaOmGVVLawcD+XeK1NGxKmQTDa9/b0Q534NIx10C4ZXci
rKgs5UCF6rP97TjUypnTosHhv18J312DJMFoqvF017aq+Yd9/l67dhzs/zUYGyXO
X71LH1g8XP7l2kAPzm6I2Ultg2EWVf3fMXEMEAm7quRitcjyZyacLrUZBlXbhabp
TpxM/m1xxfFWmDb6iQjATiWfpYkawk3qL1EkZzvc5Us+1C33soFVAkQ4tYcv6YVh
Ul4C42upZaztrjQ+SNgLSeo/ryUkEe/PXuRlb+atYw4KgHDqQfyYLDklOZBQx8hI
TwSAWX3RL/6JrMuTiMIufREoG1tBVmbq3VPVMWZ34vk5GLsjy9CMzkNyAGHkZV1+
l+EebKx+s1ryB5C2Ajgi8V5CMAXmWs9/XbDJ5hzReZuc+OWC6c8EdmyVJOcjRjJI
wdiKCIeEmt2+/hNaX79zp2zpSwtX3MXaNeHpAG/zKp+UdbGFoy30kuLoumE0Ps0+
3kS/QBBF17VAzKAbRKLt0eAnCb/X3n8MQ9ipVubl/yHlxvUHudL9F7eOV9nDC7S+
7931qsDSHYaF1LAoVpIT9abNvaM2HdKSdUe3czG/jvG1IhqbEWd6z2shw8xSfCGx
Hl7RoN3hVZDEP6XVf1oamwu8wntuHgdhDuXIoH/wHqOLJE/Hx3vM9s/OWjM454D2
dBDI5xwuQyaYVzPW2jndOcYc9zKS+YUUCntElMvOkMziw9Mc6dtzldrdfX794X1s
E0Wi/uEc5a7UaS1L0KU1amZCEcmnljDNB0/6ks4m7dYbKX9/fuYvNpAabYXlghcu
Gi/+wN93Pht6lObz9FU2tjVkgWnELBfZwYquUwmgBWnqQP6gE/ioLXIApwPRrhf6
x2WyVURW1PwmiyqrJaRZ/WCTWQafH14WbJd2iGHHRXrANsjnar1tD+PkzEdB6kO9
PPtzB+xRy6gVEcaOi3m62K7CAMmzH8uhxhNAdY+df0kLE3bOjOzpdMfjaDMZ31Ov
t4sINcBN/kP26ZMiABwI9rVdTClXkGdbYr8syiLpYtskJUALtetoCqybVMlmCTDb
ryokTLXeM01Yi42TsztDlmri9LpDli9hvo2CgQvMnjsTHhjmCRQjhiKiA8R4Bg+X
vUoDfUg0jaSmjoInOw2ITkP9BAmM48+xSlYNEvwVToIlps4rqfVYfYNWNIz/NZAy
R/oWdxSfIziVCq0GzBzFunWRVDIAmx3m/skmcqRdBqFUxH8HpfZwHsusQAmGshy4
SlZ3U2rZ9kMOM5CP6gJX7Z+kqXrIqSk/aWD/KAQJvv4GcQe1ZwHR24wwHaMRnLTh
rGMk47/5pzbeoxCgph+mIUKV7IEvHm4/KCNdGm4Qu8Z3V56czM9M44PAyy2N6Wxw
N1enEFHNZgBbZW46Me5RpnxzDu1GqF9NjKNCjzBlIk3CiPyynT6g/VE3rtGSdB40
YZ9chOCi62YgRp8ywe3QVSbM00JQSSHyD0rGMilDIqKXSNILFxChyzjUsMuaLVGx
YCbzxJfCmceGTeBfEZKLuyRjg5dqHj5gf4tOAY+lGwAOpWe6Kz1tPFA4tCrwglMl
qdosMXEweIcBPVVGtF9mWZDpEteKbBz/BeocwS3KxB5C1tMOGx+hUCavio72nf//
iInvUGXi5QcYIC4viNt1UTVhJwsEIUbwmZt2EFxlv7UJmmiQ97lDndrIbrXU+x0e
3PG2DdELW99MJvOjtBjcFRTkZqx+npxF2pT/yWM/otHYW0bMHvXLL9FDh4BhSQX9
4m87M6yHwCZMFjRaFKabQOzPbs6waqvlqDDb/oa1fpNEIcgX5CrCpM40cuxXoqpn
fmAoA6qkqxFkyihBfm//s4G1v7C2GinEWqKgoIYOZzDq9xO248l8sFQAgk8VJa+Y
xy8p54Y7ZUwx7wjsuJ1g50pHRaSAtkCrXq3bXK5HSmiiskIopxcpESzia1X88bsJ
QcYrNWa3IQHhTNOtzXAB5ikuubW5w6GyhzDTZ5UHmfAhAH9o5IceEM3gfEDB2dE+
KSHgNc6bUtiIu7J90OZbQRbkvxPSmJUpf++EdGkYfDAksE+K0oAWuw2tKEOkCnIf
nrzBoCL2WaaPlZULYBOwwE/NGcs0rhZWDEq/jrh5g8acWP4p6lU7IfuDBaEXrYHS
NOcDd602q+SVBYi5Oe82ezbnYoWUxhpu3Rlcgr23Ka0HtEbj51p4uDd1UM7EapRW
rmZpCKwL7f3Ib2LuwC+6VH/tCaaD/2I2khqMEbyJFi06RfY80kR1OBPko3zjQ9P5
bm+vO6iYuD9zJQGOOGpUYP2JX6dML8AeFpSfG87SPkj7u3NOnXk0iMsCCGWfyNKf
cusbM8BH5uw+khJN1R2OM2KXn65RZHcjYKkKXzxlfuNmhpDKWzF31m+VIjP5JEx1
G+16u9pho3cTvbymRArsywqYZuOZFfZn0z3ER1pkpgJk/kZhSdF9qHZBHDT26Ug9
7Lw1cY02p2omXkcV0sPLGst0p+7fsaKcz6NWA2/7LVWX9MvJ55p5dG/6dDybNOod
Yg1zYf/iv2fTvzI8p9XQy8w8oEvDI9eGtDC+4Hsow3VJdHbcHZReqtUK4MbHrEPK
+lhPO7pmCarsav3AHZyV8k4qHuoSf1vNea3zSJYAMm4NhcgyJTiRoVi2dSLIL1P0
aytUl7ArMfcvwkkxIk5klSxRLra/nVKvjkwPYfxYdUwm0YIW6RqB7IRQZ0L26N1t
1NLAOj0XhKohICJuT6nmicDKE6Zcl/XxiyHBGTv1kAJ/XddIf7XqgZZgOQro6M+9
43vHPB5x+B/x9szCEX5FYPIMM13ljJI/0O4NNCg7vC74y4o9dZ/niRxletwYIiHo
ye6/wZaQbAS1VSqDZjI7iyUB73IhBsfcE7zSOUXBgG8q4Zc1jw0+jNRfaU8R9rP/
Iy93selG+iSNvoVsRthxbfPtRL8kX738s1O2j7hyhSr2YP9G+AR61G3dyWOVkOrM
PeldAyBuhSOrvyfwCzb6JgzLgX97gqLxlvYKqj/qb1j7aFDsjaBA5ApULoyUb7rC
wnSgWJqKkTgEIqbScLDGK6GB8+VFat5ofg6lwKzpiEGpJVHA5JwR65WqKLIpCQOa
KAP0R5zevrws7DUMEMDmHOFg19SIJXpRlG+GWMiZnvGdyOIJXsmxjEHbOtPKg4vl
BkBX68MzH9DdobmxV+nnupINka7Y1fNFL+c5EC4yCe1dV98zHNNxjkUaAh6kz89a
GVE1hsFX78SlXWuf/P4QdWJAsVTmd5wHAFaEfQg19Pso/Gsj8VIntXM8txbYiF1D
QgfAaEj39xjYMN7wrFK/GrkGwZAuEiN2M12HjL5ibHJ4eEvK+FoYKRE5yTO/xqRI
6shvNG3oE+WDkAYVV3IQoDz7z1GO+QCiDjg/OXeqT3T090k8wuarcskGIsgkHRC8
/7DydtwWErKGrWElxGUl6q1Y4BfKyf8o5DcwDr9/gpht2llqq8JbBc5U6SgJ1pvg
9PTcp8LuXad7EV/Od+X0P5jma6P9FFGK9j/l4o4axUaAenpjdXae+dLSRq1+Hsaq
HjnrQmcAmaYhpvwQdZHoCKVhpyXxIVUDNK539t2RnvZatmnsKZUCLqRYfdbug1Dx
/wNqFVtjeU4c/27oB3TBsO48YaJctbrsY75DYpZNwhGM1WPz3VzY6DrosPVKMh8B
j1imf5y2kY3d43tv+eCIdDWL3dWtY6hu7GHX810hcwmZ+ljRbaLLgrNI0YU5sTm7
eKaRcBC8zq4wbZkum+PhR/bDxV678CDPELeoxWZu0X/Hy1eyLogT0haFjaL+OTOB
4CFaA/i03QSXeTPFjVQcOIB5P8dCrU9yt4+r4C4oQTKP2ryEssXBSgA2u0Am7wjJ
ipGF+76CoevuF6Hr7VDo4vTVOkqArnI/0lCwtXxxbUoLatt8B0nHnmIdw/rdkKX8
1nMFgjTuAMnpkcMfwdz4TNhTWTYzwyofLdRkbgE4FdUUv39AKkxrOY1aaylMpSEL
Q2U0k1MyxFzyA8YL4sDIacdHJUAPh/3aQcqU0QcWtMyCFrXi17sbme4QXw6cxyRo
EX6HQfNy5BbHZoZGKhTYgqa8Zi8J1W+KZoGlErKO7qBgh4Nsu+gq2WMl4p0FkRlf
LiGLu3x5l9KnqylrXNFVwQYGDfvX4dLWHbKgNSRq8W1rQe9G2pR84Sdbf3q1TMr2
Zsq+Lhb3JJHGw7yCqch1q963zdI+9IgwIRJYayhAb3ZhS3odlfgONSBx4aSW6fM7
RZE/59xt6Ow1t/RjE8vh+QVjZrkplPRCtz86Cqa+pKV0t7uyvCGHLuuCvQ0IZ1+u
gR7CGIyyga79lYwqsgy63FDlMjggQDlM2te+yweKdLC3j3LCrZfLHKhRWK/gQmB0
3DD99fhc9NFfGb9KZXHqejj7qaee/FIfhJBrwnuA44bcSvKQCtG+KUGWNc5CBr/J
MraT+lSx6KMBysgjyDGO6Lk41OKXSF/HWdy8MmQb2jL4WfHr7khn1ujBGoQbv2qm
IsRJ8x37aOGyhVbFCjCHL88S0yjgbfWvDHdqjkjlYMpLmw/PPfl5SK8CBNV0OION
7XVle0JD95DRvARGZVBQ8bSGWmPiX2fJ/p/6n8AMd1K9d4nzy3WI2sNQ5sLuyDX9
G+O/kzANmkH6KGyuVQbn4uGhzDznc1s/g1OZlgvTXvJ91BLaR3RmyEKlsLFm/gsN
F8yxCIKULyPHdhzp70Gp8ujjx1vrQH51YSsojhZnor+8Wk9nppjHZTH2fmO13hWc
RKu1KB6VACIL3tCGEDJh/BUjg+rryovapR1j10zw+NrJWND3eJKf4m29TII4zt43
ISYu6EDnbqK58I9SQlnpZsIcddKSRe4/OYEToagbsPF/ETbDKFmakdRbfiXxNH3k
wuKIZUSuRLrWzHWfxiBIhHNUa0YIsiRs5/qCXbgEhaHoyyGV3a7Nk/QYWZ4KwDei
RsApKjh5ogBScT6h+tTpved6PTIM7HNbsyrSE3LVDJ4NowQe2P7Ti2V0ZaBhxswj
Heohguo/pJDMBYoF8irWvo9jkKrJ6+VxX3qekqEU1yqfMJ4kVl1K9m3kxTyuF5KM
5jerdxrnqX01GKSy7CwAe9y1CyV8Gtg8fTacVCbp++vsNTOnjWhtR3gbnivDi5zh
60icHiS64PRT6YqgQJQfZ73kYHTv/oVF2jDOtxKl7vipGY5bYdIQuFawjBUDTLD9
aJ4g/e9nsDqtpYtdxvEvS4wXdpQ5WnCgQS0f1MmDpFJXfCeCkTiVw2nUyMKg18X8
q9FoToQ6KdhRCD7OfUkPlbPHz3sLhVuiRBxPZhGocF7yqItGZyl3RLgE3DFHBJfl
+AgqgPOMB2n5Vp/EJE7UvcmgkT7aBhG23Pl/fG9JYBwJx+IWD90KNxaMCt8UQVDF
BqQgozh5/9OncOfSz4X9eS5Q7x1to1gSHtcgbomqUqWP/R4/xkrHv4DG+mQAK+b3
HmcfxuTR//Ny660oLn3DGl6RiTo0DCrnWR1ygq47Bt8n40wRUQzw7xZssgONomcZ
lTqLDIzYwSiiTG7Ahb+TZDQJQ3UN+ljaXA/WDFPCuQHZpxtBoOiT+NpX4pdDPSS+
95OekySfjO9moo/BUwA0NgnEA/6sNKupkhRKIZslke9jCpbkVtFL91T521dkWrVK
C3unxK7l+pgQmhZjtJuGd863YdbVARVkAHyjZaEGEoi5rAgOruMbnVlIr4OhnsK0
4SIqJIXfOA3uP0+ARbI343PAHxfwLcPpN7ZKaGi6pBZ4UfrhHdnj8UwgjmAW56jw
pW2rLaSVcLQBrbJBfj9IBX9A/F8CM1OgSbS2yRm4lJhb0dbESuPrHRiEDWs9cNJ2
bi0acCsoig85DfMftkrTcQp/BeDSEZJAx683ju8jAM3uMR+f6StnE3wZXL36uhqv
xaJiQG3z/u87eBGv6jg4ngN+DHeq8YtheOqk6LjfIRHFBHa1iVowL2A5WpvNgTKH
CCmH54gHuArAhyiVCrEqKXLzdYiMKhgl9OMBCmMl1qHMSvfewhIqFSUqOlf/Alg9
5zs08D7lLrZSRpKDASDLMeeVDNl8DpsgGQb0YiVN1iv7drs0YfyTpqw5vZDxCGIJ
9KXATOQCjxEW8JsU/D8TePYNcb4gCLPbvV0jJERNxpU2I2MNT7GnRV4oRKYbI7Aw
Yrt/0KvmwRJ18QNRKtk9PCCY1Fut47VvEeZ681OXhP19Gsbr67YJJyRvwNVkFf/I
pZWhIgmRi5FrSPSX9E7vBppPIe0+S4I7ceFaPcDuZIo35bI6ejjUxLjLnN9O9Inf
DUX+DRdsyEFVl0WIh1pwVi64mVt+dy+17R7rBuSm0GgjE6rC3Rf/Ryw0+BZOgj6h
eM6foqx26Om8VIY7+l/PzqvVQaHWkMapgNthy+DTzeDVPA36by2zqYxOdVp4m2R3
Qmo7FEqOovLF6I+238jP2DyWwsg8two921LzekaV0sTF+fGbR5bt3K7qEXs4MI9I
JqmXQMgot3BCf97sTdtBBzH/PrHXCR9EijEinayAoI2kYf6AN4fpbmO0ZLrhXGsY
q97KFhn7pAiSIz1ohQeQqUip3OYKCac13HEntfT1nl6oYjJSbqcamdgtHn4czRUZ
jHC/XUu79ueXTZv2kCXvWXbCXrlIot1htD9w8717d3PBRIJlTL/APzptir6QS2sX
PWuRE2WBV7NbSdXAqHGMwkd3UGRiJfunvE3dxBzBTlOhb+OXBrpEsm6lhYnnOE2H
VKP69w3rVLjCL8QitM3NWg==
`protect END_PROTECTED
