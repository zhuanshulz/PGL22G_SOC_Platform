`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cODPYOUC6fxGIAplQTwIsYiCCzVf/pXb+E88rqTn6M/Ib4X4g+rLEQeecuRir3E3
R6Fm3PQo2dr4OGOHtIt36Bh15YXDvVJhFpzkautFAmZvM0hbWoI4HTqUn+5Ab1TN
PE94WG+Uud54vnc3Pru3N4enTiDiNfcXyn9odintq50dW5pn61q6gexJZ1a/JYSQ
0jnvyp8E9hH0q8nx+cMbWP4o/RbvPGLfsBpI166ZP6YGaa/S6duXEqbCH8n3Z1ME
skHAevW60dgKlOEfTpqEvSRb39IKdP9HYJrrAvirCtdZz9Rvbw60L/qKmqnDxhHk
wdN19YmVTfwmU/UvSHbxMQen0AEl40avmIIzYs//7ZPeiWkFla8V0xF4Ye6fzkgn
61cLzrduKGcQt6L00C+nWXmPCtWmHlCCDiXGMEP+uJmbzLK4e4T0tucyn6X5Ppn9
MzoU2/D839TnOH2m0FrEp86wJ8bLYmLxDjIWWNuBEPmoZRgT14sI1/Yf0OoqG0sQ
domPHPK+56o1s0TeNUZzMc0rdvJ0xi4SMxl8tr3RqpfCbv46Y0YicLdUHGNzGGtT
WmJRK/XvQl1sCcAJR3JG1NeTjqR0/mmNEjQzJuBFNeUuBvp0mrh3IaNqYqYiAvkz
zyftXkTXDlnr5KN5JkL437OyfP2AZowo/2o8ABS9/E/vZNjC0FN4pP/O6KqoTTFr
CAD69CPJjY3Bs/gAGSylxjfs8LaaUmgZa7UIqURe00tCdwP/wMj4lnbMJZE1OB2K
gfKDHOaSrAOePf2mekvEzXT1KXjRxKr89j/V4izR0auBiv3/T0uf18QPPrwFl32o
HWQRBGBw4QtUdt57KNObFRpVd36dddBD5lUjEaXVhlxQZu2oR1819kBjIgHexfxC
ruhxxtl2qkdHVE+5HER6uggZED9FYmZHaUBrZ/7XGUFIxKjMWD5RAR8UZZlo0aYW
z3X/J6M2D8mpqHOlXCQGjkeXo/+JEvPstqLCJUMoP8WGyarHdxigMZEowzPagz6O
jlBE7aYFWHmdCZt5FCwBiCtFp5NEVAqJ6kSBGFBxX26kNMwIuK07JJcTVgJscT8P
awl9Zd3QNVUZ1kkcSc/YPtWatgeuo9XXWzQLfyadB1+IY4OuO7RVGfrrbF5pK/Tz
9PgFlfgJ7jTcqcvH0xKBTn8o5aSzWq031+CK+GiO5+HEBL+4/u4V5YsGFk6iPp5Y
FQ5iLHm5ra7yAj9c/vCr5VDII3HKiPGNWt3Ns9nDqs2+AMHfaCIys3rHNAkDqgoo
oDGCDv8FWIrbXf4XtZSgs9EqPqXXTdhgQUzukYhoBgFJZdgyVI1O9OaKkEZj8aqd
ncuMERSsrtHsnibdfdTUlmlgrJ3Z/GG0yrfpsAlQokNZpK9f42PTnp4avkFXi6gc
diCpbaxFPSEwWShXCWgDEmHViw3GsME3CW3rwfjLowfI70WerXTRASgmAI4JRP3P
jlqUxT/LzXC6wCAcrOxF7ZIUlfv4PBrYnXJak+Sz6QYvOU2TvE94mF1mRFI2IwDu
18KeClCfI/P1C+8YvqLfgBr4EqGFPd7DzX/lq0g0bcxCr+aNj4RJ+KS2L0fclwhw
Y4gVX5JB6Y9VtUI5MN1OJ5MQObmTxZjcaZ4RdqXOfxVGYg1RQhEgWkRsqNsozuoe
6qfv4Y23fy1DBxVxot3o/1RA9QgiDxNjWGUENAeAb5/yJgMaIuluBIShWY5QKUS+
d8kM15pLDD8nihARQ9MzRTyHwm9CWbFYn9GDhuE4/KQ1LySoEaOfCg7pjfSi5mf7
yZjvIQgHrdJu4wLXIpdPR/nqeTYOlfd88XyA2ApbVyJmUqvxLzDJLaWIIUVH0Zuk
w4Xyv+qTT2kuGgi+nzDfIoN+LkXO+SGcCYhVxZEjPK7/N5640u8MhgggfqFy+tj5
r+2o7rKxzSnuM3lkeI2IJmQTCsLaaygFDc+gGaKnzExqqeiOxL4b0zyWswa+xzup
k/PQcLkJjnRU/JbbcdbbqQtmqzBDdeeo+SmZHp+gckBBtmJlVLzA1bks4B8GjZsO
DOH59zFQdI+NHBFLCCytN6kVHQYngx1ILNmkMepl67hmsz/hOardnens/XP0umPI
3Ae0mgVpMsVGZpCcUf+5DCYOFKWL/9uZJW6UuqgZumqMM8HGFNHFif3469wGAwnS
S446sK9UQwcDZKMflcN9TYVCbaXFlSRNLZmeJHk8nqiXZaHXdH6dssby3/e7oH55
5iMcs8loEG9OaKjIYQhCCKmao1AkqVTY+5AT/ioFgDU/FzFORv/A2lzAkEBF8uZO
R6N7Pocb09NWs3BHOzuBv00GUdyOfHm/LE4O/jOA37K7fPUDrBUonfxC3f5GED6q
3HJQ7lBtf4ABO3PU6UJkE4uodlXlkKdVYPaOnWKE3YPkMoJNeE4XM1V5zyUnjEqj
QEgrWFtcweLjZiFBxXykjSkAmi4jLJ2cDy+lPEBXWKhhShqeCiSy6IfH/1ef1V5V
xJxiBbal8BNXt4jbKgWnJ/mMvBZpxsXTJ4gfWl/lLbLwUSgul8QMIae81IYGu8me
n1y/hzQc52lsdl72Q/OEJbkvnJyNQ7CcQTtdanVJ7vDv7p5Rw30h7lsYJ8iSxpWf
XrsIxz1MgeBC8NiV+5o19a4tuZG85rQOWVsmP3dtI1fSSvguDnNGzZx16hIQjOTM
AdU3mLQ4YXG4fyu//ZOrc7qmqGAmfRZFfUW1CBw9OrjDlzWedJliqO9Wpv+aI3nV
CNoH7QEYGzZUl/QcgvS3lgzaClcWo/GpT1OxtlpseaHmj2SEoJV8Mu0KypgzBhoM
JWyQnRL/lSb7aAe0GnMRrEAcztvMHB3dv2JFpx8rkJwH8Lq+0WFDe7PTA3ENkIOr
qh/FcnNmNE3BUr+xIsFpD4dEKolLVpytX/kjJvG31ivs+V6Ee0I2O5cuQvpHZ0Vd
FKxdGh6Lf4sYryFkLBhnCEgaEL//eLmx8aeoTE1OPrzBlnv81wy6Z6BD+AADtstH
Lu8u8ttxSmWmFZ7macD2gCfdMGSXUrtMAWPsSldz3+ODQ9njL5Wwx5d/fEpFLA97
n+28mSU66v4F4Mx10Io6OBMjjoU1r0ES/nxJJvRQyo+YoTxScvRfxs0gSGUMLl9/
8i86lEBK424n2MVaqjwbfTsqtFfxHYLLDrOhlSDyt3mRpEtDtL+OnE6qSzpKDYcF
sUsgn+Iw9PqUGoSrfkINIXmVWbsZwQHLWBUxCDobVL1Y7Ncr7GiJhaP6bLlvq4vO
c9k7D4NGR4NcpzFWOSB1DSOpM/8GdrScI5uX3EJl3HN3xs+AiVc2A/hKmbug9qxS
sgoy4uTPHg0NKZEyfxU/k80ZK3cKtth3iZhl2IrFw7dTzLLcW2Zk9A/L9NY+ltku
AHHdc4QqB6e24YPC6EBML6znb9yIcUb8v81+SYmnvBfbSgcjcQwd+Jt3wARRRzna
3kZuFmCs1V/NZyKyjxOT33ZJJBnbmtUL95tSVrtYsnfno/qx9AUonClhka0HzTg6
I/+eIf01Wn1trTKjsXz3Ljw/i0o5B1DAi8RO5lWZ0od2Tz6ml1EV3XVqmin5knjh
eB2WEXynib6t2v8S6FJKkRWEDFG33mleBy3ITGmCs4OTRhVlGhU8FYfY+QcMrjBn
5GpSjy2BaYf4+Uc1pp+mt7qmovbzAAoHJPk6UgMyihaR2rtqxfpPkCSvZ95GTwYv
Gugov1bw8khG3xE8Bx3fF8Rj7UyeZQMwIc8Yntlc/8LKF9+RQMGCDf7vq0LVuKwp
BgGqBnEZ7eQGa/+mMqOl7dhXNAufWL52V6PRZrcc1DDTon8nybs1nqpHbzTC/Fw3
X6GVmL6wvJ0gWxWQ08v5RXlXtD6v7t7hw8gO/pyp+G4EDlIToOnC2u03elKK8Sx6
Up8pSk4QBZ7HX018HhL0Z7VvCoQeQaMIr5/An15kmH54PCEWWXhwvIroc6nwdI/9
9FytdNheqHP+wUP7ivIzBFVaDLawPxwIqWp4z+giPRDOPi6JlVPbun3aJlf1OBsS
GIYE3+QokJUclfKeUZNKXvbZjb18WEb560fpn1BWK45Q8sLErgoK1qk3PLgSRzF9
Tp0VaNsOVx6XwGID80r1vNdR8a1fEGK9RUO0ucRfrknQH4rz1/KF5fiPfdDI11ua
H+H3WTjnXBNXfHtg7EMAAohTNovTFQO+5VS60DvGjgdfoyl836UFYwf0dDgWB7Wj
LV/tEklW2O3im3HoCkj2Ssybs+HMXYw/uwq5uxl+5Jxym0u1LXcZwHjjRwTCkLVg
Y3ssdvJkpLHvaj/0TSBmkYqWsXeQJDDRcfOQrD/qdjV4eN0h0t7tgE2jk0eorJjz
BeaP/sZRon70b5nxE1zOiA38+RxHWvwxk7ygywoeY2qNKXPwr/2vJdrMuoEO1mh0
PcwAiDabz2W5F4vsm5MJg4bvYOFz9K49jW45WP9gDVK+g7kww1BfaAx9o2ZdTBii
lZRb1RM4QpDAY79xgYFBQdY71PpldVG8KMEI5vAelkyh3cSdKS1MUOnNmoc5fGxG
Sx/+AAOKElcEXgMXTApWEcxTNWm/D4lLdvLh+9GiNon5AqpTKQHCVNXNalpPSLv5
B977PVfDCVrjgOChdLEwQdwmKYnNP3QITb+8B9eRspNEbFnmrekb/LIwBw2yVaBL
trGdTnOBCwfVm1ZhJE228ZPj8tMIrMh8e6tVy9YcQ7EeYffzW8SlPZ9iPkeEzIc7
DQTz5QIsfiog95U18vum08Sp3xSnyEnWIaVN0Y22VOTHFzuE32InMDx5i/jYFB2F
KNXRXdYcHWPEDTinTlKtsqr6OGGHsIBYorbHws/7XHAnWgOZofS8r5AhXRjn9yhh
gRDO+WLds1SHs3k36K+k4l4v0jZ55gyqhrwwY0vSryfkDrsliWtZTqYz4EUd29Ip
7a5VVDglYTb7ibbOAP2MZb3TGEj9MTZlu7Qf0ylIgNuO9b+J8sCSUP2YRKM0kbz0
0g3CqoL1H9OUCJxd7P2eg7YSn3w29ctkSkkhlLq3vaCkEJQ8MCkIIM8migNxaUA1
fUPXRx76r3EoGAAe6yYaLR3+gCAWbSinExWOrS28MPHL9G+46SkTNOHgCoQ7PGDX
yJQDqhzm+/lKNnnN2r8eW9dV0s80uuOsWHM/ucccdKxCBePYz2WLmLLWDGA/HiUW
kS5febUXm7TCM1B5RMydNg2+XPFUnkiAvKdvI4BsNflCZzttg/IHUrRqOfbSi+as
BTPXUVClnae0/B6tBTo0sekFJDWS7vmx9d294Y25u1cVOKGoQIe3rN87qQdW4Hik
qpPPzxt/4SeUCeUuFbcFRKdipPFxr6sZU4/cSE7NM9T4IO1bVasNSpgYjMGf6Lqt
ubMz48zjHke6LZyM45wOMNvtYONlnak+h1gLbSUDawdEMPy8Q9u+hb9Z6OCBabnk
k4YJIdz3Ub7kg0Ia4evaABp6QxXpKqKTs9/5fftM4rGJhmdAYsujy8AFKpOherDM
yt5yUl2D86ZKLNgBD4zu9WTF6L/XP3x7OcDEcOyZ9xnr3/QHvWViz61Wn4DKH6tg
/DZL9XtAVutv/8dbd1sLoAYL5CziVhfQuAEBMYvqN2H2LJuIcpPuKzEA8BUXhwDn
sObXBQQ0GJxL8dQ+BPRh6Ckn1IDJT4Uurasv4ie3I6hFicUARJ6FcuZjsXeRoVqN
rNHu0HWN8/SLn8Ae2tCjXTe1Di8oblGraoAW6j7ZBg/8mRWyx++OKXfc9uidjMHo
gfFoIGXjQp6S4CSLUA+uqnoGpSrJfU5CF8iO12th0JoLLftwYeu2UA8PDIRec3ka
2KPSZwme0HX7TPK9AEl9tE2/uGN5dQXpNm3aPYFNCg7hO7WpBZjBt5S3GQMet+45
LFSWjK+UacYlKmeooiKTyf7GB0hcgLlwSq/IrTFGBEUFPj/tjh2iF2OT5uS/DYZU
72ehAP0I4GI+3i/Sc0vhK3HpFnwozQ9MI/FE7BVqUpOqKEL8sQE4EHC68mt5KrIx
d/q/THp838bOYQIvdDSTcuVZ7WEBcUdT3Rs5OrANR8Eygl7XN+DXEuEf+W/TBUgN
xVtHGhVfC9jowJQFhO1ezXuk25aa74taGRrzLTD1Ws9lG0Sy01q0nf1BSYAiwdEa
0edOJ8CKeXfWSHFWfIY42R2WfJimIoGuU0kX3AE8rNtLXtgSObWVyHR3n68Femeh
MvPJvKDu6pBUzgEW30X6nVl35I8GvfbpgMaQU7UiP5/xgVMGPJg7hGKk9tnjzhkT
ZTxwSJUJV9YqR7418kGbQTqe+vxdSuuZwydzyES8IoqZd6F8FPncB+H2Y7w0kRh6
Ex+GUegp3Sxsh/5OhYIuutUEwh8HwO2taEsJXI1s1t0f05yyB6s+05kAo51FbxDN
ydg1nSDSz3EUjc9ojqv5sfYIbGUuicWXOBefXv/laSIgxk8YME2UzEWUzv+5QZig
QiI7egZJ/f8GLeCUJL+XSSX4FoIdfD4PfFAKCqsUNonyVYjDWc+DxwtG8QWKrURi
RBK9uoFnXX3DRMFPlj6K0NmmDCdB7FIg/cLEVF6VZaZUczwPFJlgUchYr3dFMiA5
pm5v69Kxg7teHvk/bGTl8dFnOZPHqJoPzlt5hbFGclFU9TmeWCQKQEjc3pEuQ2ek
CAJqK/8mkJ2YzwI7DTFGexfC1WL0UEdch3VXzGyoonDLTC6JcBdYooAY+J/JOFeF
nJ6cs4t0EWTmF7lfnbjmESm0DVeE3GVBcmX3nSu/AzGQIQtF6BbjtWFGjd68yES+
o4QL9TaU1KO4BCeaO2DNb8Bv8SFNJ5rqQ4ZuYpnaf/oWw7NCUFCpVD8leAbDOycK
MKLMVzxnRJh5NphApe9RzZ+FzdI+0ZojdexyX9wK+4NsCl2yyIxHmol5GYJtOD/5
WlDRO7DzbzpkfkeFvrSMyhN2X6vXvxdrbOAyNB6As04/SKTloOKRFWcZ4ZLXR5b2
McUfzQuVOQO/sJVLH2Ahb9NiDo9TiSINcUy/im+i7QfZ70sqmGKeKx3V2m50wPbT
0hZlWNF6vn4KfWaq4FFx+Og7rDR6axVtTEwHZ7p/vecbxa/GpN9ubB1vGcpt3HQB
4Kwt4XIqhat42+ck3wY5mn7MIOsZpPjIBtX0j8doQHb41zepPgE7XHCJexUtGc8P
5wu8Do1jTRR6B2oOptgf01Sf5rndkwQoX5/VKh9q5Igte0kuxHjeab0qGaZsDkkd
VQvMAkv+4mAiFdOHlq+w7CvEh0p7FWmPM8gV1+l0Oc+tTzWexxd1Ek7mE4HwVwF4
ExCiJr8FJwxEfPTs5SJjmOjFutvWd2okAyP3Iadfc1zVgG2dxDkzUD09C0lXtYFA
6Uz715CHK3jyPsathjTygc3HNrLTcEIbohM53uk3H6tTk9xhXxplS+WjE/mNsH2m
/cZGdYXtqJZSfbLAlPMU7s49VR7O0RhGU5EmAyE2rzgoYG1K/qfFRiCQN7OMKXj9
uVOQq7lxu6tURglFS6Nlc0CFu1bzVhwBnmzPvx0L/axm1i91+gDhSrOqcUsffD/R
4HeexE+RvfNIITYAaBqYHLNApR5q3izX3fc1LtaOxJQbZ3ZqWlJroWJBz2UokPqi
kVEBZ/IcQ4iRNhbjWLCMwz6/pH8F4/h1I6386xEV0ADqsGZkQjSr3ED3X/RaweQR
y15xeHmE5zgp39EoIcN3brx8qpnQeol19MOPS6cfv8oCfZQSV5XpxWXbj67p2wJt
adyWA7faIF+/Za+0bOFWxwu1sqkVF0y8dozR2b8Sc2f00kosa+kGauX5It4B0N0K
hUAg5Y3zaRZp7oEjWAsCWZnoEC9Wjo+pJ1qWxMw4GribEflO7gLKNQnV3uvahhn8
tRgzQaEQ6QlWjEPJQpaFd7Kjd3mVh/uoNA6cO2YlYI7YO1TwlIg+7Y4vH7H/E79M
kAg1OVmH5clxr11V8YZxUKTiqQyOHfe8H+WiDkXJ/rRJA20lbHbSFf8mFsr2cFXo
EhXDgl9/01gRn69ivjK/Ew6esHfJ8uLV1PO2VDOA8fVVMqjTdY+O3rCv1B/E0EKJ
C0Cza5oR/DN0fFM5/Nj0/FXk+muXMjdnxn5T4Y8DyRBUqbrfyl/bWI78qeaTwB/t
xtIma1VR0S1BClZWVJJ5Bhy2ETQpSMV01TVE4ok60PSHshxIX+VByI1yJIf+ydTt
4FL3txa9U7gyC4jVbsj2XWsVvJMGs9hztaW/kZJ+kwFsGJ5ew2vg5tQYr6Qj+p88
DZHmF0MSAuztDpU4ThsfrQA9pTKwyn7Jvxp0UdEXEDOmX5hsJTdBKDBlpeugDpke
niD3tZe0XbTTaWkwik1/Dn6TL15WvJ5qHZuIIpnJYp9QoG1qPUc8emO9JcvwjaXv
RyZvvw1l+M845i1gdatYxIWvFnWMgc96wz0N3FCvsbp68BDmhm85Il9ZwpjhGJtL
babdorgx8GhkIaZyctif3rInPAzNdV2HBMrlMvMZs/hZWZeFN6C7vYreL1Dn2OsC
/NYaoWjmwDd8xSm8ilaSZA+id/KJxUcPl4aTB4BrWnPcwBXyN4r46EU4nBF0CkWs
73+zuNu099H2NZVog/9IW984JNIhytrOI1j27VYAxIKJ0t25xIEitA3PKax0EjNW
dtaNebPcOKNKEFTOK8jTTTGFXYreT62B7D5DdFb82Aw19HCbtgmHhvYvBqRf3JH/
NdRJhezimGDkDvrqO5Y+k8GU3PhF1ja/UVXjz8XPOHy1Xt640nqXYGfLAQbEDLx5
ZTiSQYLjr4cG8uiWLb8CjqkAcbcCyIO5vuBPCXPZw0A0hm30rbHQAv5FOj7zN/In
vNdN/QhlWUTEN75xSF4Kh0nh23/pRqU5c1C7WUTGKY6I8DIROpg9lRU6fLz8LIK8
/suR8Vvgae2RRMiqr01cunDbEvdj2iAW3mBMA1+vBA5mkIIf8+vENvFHpPdZD5gu
maAaHfQkH2+54ZZ6WaqBTt+mkM0XAz2YDznphqr4WxNuovZrIlrkfQega4FVT/Dk
5iWXqz1UevVrlFRYSz6roA2QFyLRNSIk6C9no6AS3ALlug9Jv9J68bp4XJFAJWNb
IFDROUJh3neTAIVlIZcu+T6aF8Qw8JJXdYqOm30jVJlCWPVgIHPl1gVUMcqHVVF6
sPwuOWRrph1tfnDvdjIuZuHfCLH101lQa6XHZ7XxoeVbhKHIwfQ/YOcnZdbHPP8j
rtWxWKU93mvAceUXQGjGDsNkr8SMR+iCDeGcUzynOUEw7zIOHj1tC+PZsmKFpCQt
MOCzmtphtKWZNckhO0a7Pnz4PfqpX19fRSVcki4g90T47Sdijd6XO/DcLOkRKHR3
vL8ydVXJgZbavLfLOM5yoistBvITWsqSfDj0IS6RWY/2thDSLAHDUcIyt7oQWECX
fsf6SIc5c9Mt6WA9moPTELD5MyEqaENco+XcoufqDfDSGyQ0Nfg6ijrKMjSnThVL
0W771YFHi3+o4lcCZTkznfCqltZJ9+Xv36ADXB6yXf+04gqKUap1JM+IxEuHAjLy
IrfSkBpAZE018Z4TXab/O4ipRQIGjfuNPn2Ag7ErB3ZkoQ/TYQSJEZ6OxMacFtRV
Wo5tFdRl6TS0StQzgNxbRTzMoXtk07dKPq9mlRZj6o+DHM+q93YnaUiChAAmX3Jj
OjVLS3ql5CXlqy24w4mCrQuOOaVMwgb3+wOLrN6EHmbduVQfIlFFQQGxVrmifb4G
bwGTfegxU0Uo2AVXLHIRhK+K8DMP3j3/bUmf4zlwG00XCW9eEA+ED7bR6hLm+kB/
T3B0p1o3h3C5tr7e0eHkBlLu57+SrCiRhI/bS6IaGge+nCsmwDKa0Z8z+b1coMSG
846kDCpykNMQqHP5dXBbVsjGid7S7M7zDx6WkUaD6FiQZCMYpCo4g8qBW0Ntb97/
ODunQ1Zru0NOoLhO6XLdcwyRP7i8Wn8s9MNF3+7oTAdU1GDOmbDLQfLaD4dvqYze
feMm1W4cRAd8xrHFtPi51QJYwDhPUOHPrnRFgtpTms1u/P0YGZ969pMx53wcC7bb
KBfLemCGVOpvrLT+MbXdCxVRvDvS1rJHKOnw15HECNCl4dvGsRxLm7e88w7Tq95y
nmDmNfU9SMRnGoinLfLRl7lsW/Q6XB4g6RTi8sAexq8sF67z0JZ79e47fqhNOptE
x+VlNJsOUdj6gSJATj7dCpke8rrfea2m2kuMd4ypECcKpNybt3pYnU2Klqubl2uY
Mc6eHrK2DoJDRX6WuJr17/WEkHSfYZcwTk6vIoYLYhYYLs95qTra8afghhV+TDHx
aDKaDs12eSg30mNgz5qqTkeOAUU7oEHLP6FffuRrabTXaPZiWCkf4NhXy7Wlj8J+
TQf33zcZ22K/eQT8KGf/aScJGwxdTEFZFq72w6rwtqHBSizQ5z280WWy8dIwQdP+
EfvPfeo3QlsWNJ3Uyby+DVpz1aAnxP7mq95u/fYOT924mmx6Uk/LjfNdaSVzasdp
I8yjCkNEwd1vpzjYbi0u5neUN6UkZKfq/+afMYcU3WC7goRG/eVhIyveS/Zsklc8
8UGXhjTnRhzUudcmetHCnx0FALglDFsDc+kwZrK7hge9cBBq8go7ngTyPWdAxupf
NPf1orJwODGFGp11NCoqFXM/WhBXHihpk0i63vmxSUz693AIz7DQK8VKnQxHyOa5
vfxHx/XxfEwAPkxU8V4hgRjECQ1hPbcXP6/GT/zpnbDLZyzzWtImGk4V1sTJp4jk
hoS6f32hQsC7+Wteca4QS2rlZyLoUi8DljY31z+wPP3wYt06FV18idY9zJv9wqyV
YPALEz6RcIZXxTXdo/3aWhiGN+Y7wiI7N0tvQwZv4T2q91DR5ru3xAxv6yBemEiY
5CSbrWDd/9aq7ovms0F783XDB613nKmkZDXLgLb/UNVclckAHInK5BoVu+gC4HTZ
QuWUUScKuDHI+T5CRvqw/9Ycnx8kxzi+cV37rPf+MYT5FFFfeyg9BJzQ0anfwT2/
5HPSOZiNF00q7bneuzPIiDjWIhlL2OkxHvW8xNdJ55a07Uqih8Hnv6LEb+yVF9oW
7ScYjifRQtQZcakguxLihuIdarxn2iF1uUfj0LG+GxVHROWL+3utoRN/uuhS+g5W
9FlSqwC/uP4rybwB4R/xfMTXLx/u+MMSXcYMA6ctKa4wdrIz1sy+6vXtHcgPU3cx
pwKy/ErIGGId3Rr0h4C2ZlXqo2AF9LGxrnQRH43hglyPC+78E82Fm6PNCVpTyhli
bRUh0r0zYt1iG9cWChDvsdiMWays4V023PNOl/Kt/17EJiRRRNTexH3NuZJROz0V
IkkG1bJ0KiSnE79dss5OG4QzZyGUIMaOp5cCNR+/vIqEb68ghnX/PQFoRU1BhFdC
HTSchVJGc/mM/X6KRtsZtdWshCxZHWV9oq5teAJb+iHLbU2kclyhB5eJjgggVanV
cIyIQ5wAtORQ4dKoVrdqlsQCDvWh3dBDtk0L1+oSCCgxxTGlVdwx7xyT8MT4MhlY
MpZgSZQ8O8fw/jRVguQdhuk6lpqGf2iHuNAYZo6KtJg7Bcmbn/yZITiVXa6XwCGy
quHDvbuipEkMOwXU18fb8CabmzxdvNNhPXHd1b05wJagyXjTYsFmz7Aq//VltgHG
SeBj3JJy0zGgPUyrtAgfe1NgbtGj8CmdS9DT/QaI44OacSUoTU8i3dgnZ5H0WuOp
T9wrX1/5jjka8N2To4tydWfN+3hwsFNuiqzsdTsNwT6P+6yFT98btTSfFU4t98oM
6P5NdJ2MCcXbJYHPTdNIk8OwINIgqrCVv4gaqUpwsSR3Gwzrt5gSDYkQA4hUJL5f
FPPLLCtc91agxeR8eaPuk8MAZBa37DXx74Nn/upHu7tEE/23bFCOaaJF/3YUvgUf
HrbO2BVFBUot8lV4xM7Jd4KZzKB3W1Cq+pyGZeOClIS+rlHttboDhR6KpBzrQHTv
TwEShtItqPCnghWvbEglEBTsUZA4BcB3pD/1ZPbC3osEyZ6/u4lvzoMdy+YWAlD9
Vm8PIEBwbK4L+QMYsY4pI6EEDKbN/TbvNUvxdrSBPCM9fotfVE38u5RwdDO4f8lF
cQJO6Q9DzNeLTfGgPMEIxj3MTz+9DwdbnmQUjRm4B8uLraLt+FTdttXxgY8558T5
rkefsImnczwouLvEAuNpTAX/5CGFAdJAx1p77v14VvFCPIz9KSGC2ug3+e7isGfz
HSi6qp6HL3fPhsHmGRTSVbBlXPN7vjd2olMOgsRND1us+yDVT+et2S3YWCCRcBbb
NY23QjHWYEb4TP85wq6M1gH2JHsNLr2uhPz4p43YgwL5MF9lh1hv38XD8+rGQ7Oy
a/+KSu+Sw0004fKfIlCcAaMXAAGksl690ehWL9c6N6XgA8uf/MBPnOBssG9uQEuM
eTE/Rt4e0cXSNrmOy/dIyV/ZtlAIeITuhsmzmxAO0yedhAYNyUyI1evx/8eQC1Aa
efcmEhFe+DMzSS/kJ4mB11o227KElrP5zv3TK1692bliiU6K54O6iIk00rUXypui
dXOME/o4C/kH91Y9ReK7JlwH/wOtL6chTxuewgEPuevQnZ5Mhytu4UVFhOhdzP+E
+ryivxoyKOQnxRGgPSmpI0w/msTV42OQkzFM5xeg00mBQbUmw0caQpsGrq/8mV+o
S5o94jP8lFbt9IiBNiwSQtqR7AsREX5MxJUOy96in607gaAJV67x2OLHvfbW4XBn
1xoYLW4FW++59mYU2HoRBhDXlNZcLMMWYfz7AlP71kNPvD7U3iHV0NQR+f6LR3Ng
n590/pn5YjIiwhLkbBc/mFhkt4En5n+8cHKAiFWmCIn+GIwQNvYrGVX5FGnqDUJd
C114ty7t+l620q3+60KOn9j7Ra+nC1JTLp2rbBwGJ5Pd0UB1g0hG5saPQj7WcRPX
Y+V5xdIpml8Fobh6KGulVtVUwO2iQWEKFK/6RmfPTcM0FwsjE6JLZwKJWlartAqz
MTtb0NdjD1YyBaKxP7kWT775BtgmBbvj+aMArQtQ4V5uX/U5iD0Vo1Jw7zxgJqKK
fkWWm9iRVsQ8dKNvd6831itA/Ml/bvjUzog7+Z/8iDq07nnB7vHGZt1o+7+j5hEL
zb/1BH/EvyYJ5ii8FJey6wL4HOk6CXHaLX2vO9T/KzisjSVbcuQJSy64yNHX/XIu
K4RuhXYlOT1Ez0Cl167v9vQsNqmvU8MKBeNLNJjV/Yj9RNk2TZbWWcS6mcwoJXyJ
FxeETHV+0942gSAHRKVzHkuNRTwF0z/lfUbNM9LyOMbgf3loYQ11lFJ6P8zN03v8
iiVmoseGacTLztRAixe7Lzxj42FL2JvvV/Nnktxmh8VZ5j8I8WAa7WnUjzAaHcZR
CCEm1zLGDkM4vda3bq3vspKGkD5ZlpOosNyzcMx1YEacju/qxgAYieNCgahj4IUM
J9FKfi/p6UCdm48nK3/2gB52ZS6wXofAES8kEy8CrIa1jHkk7euPHlgHcW65wcvi
rv0nOCvdc0DB0DuIimlETMLIFIhsR8AwRlvCYICZWSWTN0yLys1fH0PpMjVVn/oB
fkAHwAXKQAvue5FATaINZ5BXOroAvqPy+kTnw+JnHw4hQFXeFPQpYKeQ/+Km2Txi
Hns4PUGnImyT0yHUbwMqN56TRJZk9kjydTr2r3vGLvthOCexoFXZ5luW9cRpu5iV
mRDyRY8K7pPKk1qHCfFcbJ1bQTwYB8XSEPcd8WDvSQZqD87Z0PC+EVdJ9VDntq5d
JxNr7NEFdx9RqyZ/qnejbC9zY8nc4KlwiE0AVDBuc7Fp+T5SAIOWRNN2/kwM+oO1
pCUm1POCUApyg1TyuD02tYEpcHwiJaysRznDFGNMwLmu6saOuR50Gl+1g8WCcTJv
eKulT1XETWcEyaCba3RiVLPansv62LPfT1kXV7yFNHdFxGsJ6ex0uzBgUMtm/sZ1
VrFfXAm8lJI6z9o9D+6ZMiYfhhQZ8kAzBBQ/yJQLEPb9BJ5CZ2qnMFPrmzoHtTjk
A4B2tFbwQTOMDO4RvabQ9aYNvlAoAIOCItkR2GZrMC6plz6XeKcLw9ihVIhZY8CJ
M+6J9fcXQsYsWR4X8raf90+zOoAHYRzWQ2Gq8HAMuNC8Mdnz5IBJZwh+jnPyOwnL
0MAZsWoYSa1KsgfIzdv4e+EN+0STHcgYzk3QLTwEh7R0Z/ilSO7nnguz/+JkUs4O
0VNgoxImESb5xyQnk1kSz8M9Ym1FR80pdsDvGyOvCPc6XrOG+Mkki7El+60n5lZC
RKnV0T8J7Davs9vdqkpkWSlggpJC4SFpAbXwoy731PD5Fv4raKGZ17kzS7lZ0k6C
fy2Tt68NE7aIQRalNg1PbQUQoblYjPsobHHJTIfOiPFjQnAzKYr6/us7S8i/ZDBI
Z9zweUDVGQmJJmrHIt4KkG/wp3Te/r2h9DFKSQ44dlvXns084vg49YsGc3Mdcx+i
kpwmH0wxKJ8/xOD4+Rilnqwavr1kJ7JaHsNkdKCKuntycmgq+LIy1Qni64wOsOES
HiiueOKxap3KtIeauGrw6LbJM9qNK1RMNT4DcFy9Cz4wpiHxoEEx5FIk/Qswt0xt
mPZBQZd2uN9UA2aSDObi9cPkHajaBT7GxdInJdZRLbHLenl8Zb5JqIZi+9w164fD
c2ZCMrRjRNTrQQLAoa2wVNI+f1/RavFI1/k721SR7mA0ClL5e8Sv5AmaR0xU3EHi
5JZlqmrkV0qOZ7u0vhJb2nMvZ65fFWOYNZJMEPly/ysC7pafDbqgZE3u/NdvEPTn
R9Vyt3fiqdDYaIIzwbOOEs0KrIYUHzDz3pafJs0D2uyie3AFCe4IqTzNZWhQLoct
5W2E4LEU309+hURcFH6bXQ/+SF7SGJYXwLqk9UGplrjLsihvprEtXWh1gCdExzqB
pflF1/NwTu5s+zDksYb9aDXh5r7m5momzZ6D2lhtqW+sbx7JWs1Gaem1PiVpVfH5
ufraLHhP1waqE+nTduUMs881fBuQyPeldlRqPaS26W5ATzIT+W3v+/I6cjslWv6A
gGMOWK58+4KGgDwldVNGP16fSNxWLOacqDmiqxgQYdyzdNUMKJSPggS5S4AdfhXm
SY7UlHQrMoCghsn0CYI041OOe/RuErioJebyv/yG27XMs4z213IoQYQ1QDOOwiaB
g0YINbzivWtgGT5AN2BhylfwqCjptNU8rWh3OjPzjrB79nfyifqPeUbIroEu5GtN
lMgDsbxzHAFAPVk9AmO/AIZd85Jb0ZykDGHaqlZoUPE43HvJhh04+8o9rji6fRex
RaZ1KsfFJhmtdWWitTFX41gqxOWBhInOC8nOEN8WYjrWrA8hYadd0t5NF2a6ohuD
wJSnIYwL1FuBOmPuW5tkRHOOUDXz/nMgspw+K1JwRAQX5hJVRCNVGCYoFGtloG/T
qFnXHVbfzGkIHEVLoDncJCBqgrp3fcsS7IkWy9r6qa5Oh/TEAYLGJVxQ7rs7X3lG
GStTjSqmgz6R9MZ+vWm0snxklg9XmSlL86DiM+MjqUZRrsHCDMsuBK4okimefKlE
DkGTTXpXTqjansxBqE6wcE5CxvlWUZrGHiJXLwc2oww4RRjZNWbRTogsYAk63DV6
obyEdIn4Q7l07nKRUw4zXrNMMv6G2soW+pZCT1tQRhdx9aM0hvjqZV2sLd6YwHBe
GZAqhkgCEoYyH82wg3hSDqCUAgkOEu2v+c9jfNLjDQhM6mxZfuvVDi77VkRUsliV
vf/53su5n5yVz722PaN52Jepk4qS5jbJNv31zlddwQto5tal2xDN8WxJvhamiryM
GnLuwGnWBQ7S6o4K9SZDPgx2BIN6ZPBJcPRKdi+RMNEnESYSMquYkTs9D22PjmlM
2+Sp7qJEmjr5Uy9CCVg95RCqz8EwBlLcEp0O519rmtgRGdthI1UGWzWeBQRfwAVF
D0KLoxFTI/17VqlTYx9EUjmD/xZyDUGvUOQlekI8nuahi92gXms+1dY6XaUd4m9m
h3m6RQ+YArP0frfJCC9HRFGU6M8MVeDYlZomxrDjgJGay3rkj8/eENDIrCXXMira
UdVSZ09Rn00gSam2N+ZhHaWKwty00tB24PnGhkMxBLVDfsuYHJawVgFl3aNKOenE
QOiOyxkuc/as7n4FWeL2QsBpg3bOE7arWyMVmGCRJKDKe95wyG3QHrsagljsRzcM
BJ2anu5/1kP9c+H/Sof0EkeAiTfwqSqR/3e0T1nWee8/h62O2BzfCLJfBV3SZ99D
IKhBF7UKEPWu1qDyzZD88jj1oZSLfDc8rx4Z17BvO0WwMCtvBmcso3+cQUQnJiM2
eXJOui465+yOgaxuN9dQe/HRLRNjImhk3DWg+9pBN6JaMefhKAf3j0FzdYtMGMlc
k1R7oRt5o1uze29eAzeTCPY+4Jg2L1Xj9dJ29wED1cQhhkM6kpzyLetCW7cj2qnp
qoiIL/q7cPzQsulsdw1GsBuOzYDVONMVAId18Nc8WZnqTA6IvyOk/xIOhzd3KHEi
eh2usd8FnRpr040XU4HprNgYkgL3dd2wuJu9qAatXXHVt7vg9nwJjl618xn5w/Ni
5gd2htScATThkGnwH8n4xZNluD+gFMrx5bIYhSohne4n+UucVQZQudaKGNBK2/TY
l0f7UaVGQs0yQZ7RcU7ydsZrDY6ZswM4iXCZ3+F3ZXfWm8g/2CVn5qIt6GT3cxsr
hQ7xPAd1lYQTrWyPnWP7wwz9M5dE6JM7TgnlPcgJ79pdi+o00ImkJVMfRhxkM6C7
Bo1BbrnxCOQdwMeUSSBaFGPCNgqvipmalN8cfcDXFaCVYwxulCXAY40+ocLDxc5o
6icCyZaBASLUFya5JMpHaYH/DqpymO0BRRa+LwA2deRslXVYazq7iA+Yp7Yt09A/
1xbDRVNO8CgWMRV72SSyw4zVn1lsKjnuzXc60KfZTbkf6wUQQJIjdSBRwmysY0VO
PfvRrFmU+OwCxBxSOlx1XECG40eNTohj+Mvnw9GilCHqIEQASqPUzAqu5yfRUpBe
t5/YqNm3rcIuCuQ1W/SmyV1wWrykVXkpUvbd59LoyJPNcKxmg0TtdKz4zmaiKPyv
38tlh6w5k6EZVx5YT4P0P4NMDCxIGA0MHPYvRJomdFkaPkcbFnnH9zQLLZwZHy+P
E3/6juwNPSqhn1Hw3zF0/AlsIx975OGucBMVjc6g9D064wOL8D2lncebT/hzXbZT
I5RJRXHZM+E+pHFaLyYVBXYz0wRY8428EKmWC4qTofxa1ichVenfwziY3733HYBz
N2ZgKyCwIqUM/GCgied9C5F3ZTFqDVTTKfXcavO+UB4Q2dT15vmvn6CMrbhyRi2Z
d+Z40tyrEsPhR/eCYXR7rG2ivrBhlK8D2JGF54rZGSacy3icgwOoSHu3ari2MwUL
4LoaXjk7BIQBpwISwmKiufmyWX/hmFYvTiEKF5dvlYrY4J3D24X5TqmzIB4PHEPZ
i4NWEYGBdqolpSgbqaH/yma8YLvFoIXH61KhcTg0qbhvItYdy8gcNTbz01J/CQZK
h78k6ZrVhWCouO6L5LR20cE7iXo2x6c0IUGeCc2jv11EkSDIWNvKW/R+W9/+UyCX
8i9W9hOFeauzHIRzCBkJsSCdMApvCYrvDL+O01RjSif32EBlBobw/d+/jZmRIOyh
Kqy7DcMI1igt6QC+OiP0W6IxWKuvuyFbaYUa8VStzJ1IZqrqEST4xWQo16zslAmC
FUKRHVE4YXDxFp/0X6dfIOD30sBXADEVIN0fw6qNgqEfCNz6sNCWLT1gH+GrcT6o
itmjHaihCwK71LMy2xaFAFZf7rhEKv64jQViS42RtcWMexVzbzDKBZ7gFL6+y/Kf
ddYkD0msILk7oTAGoe/2RLuHWdmPxNrNL6nBv2QN6ksKzO79+o8gknP5aoRPNoZ7
hIq1Zr2PETLI3CTxo/Ag1WBc9jNGptGzjHeiLVMR4JrFI5knIrFkmISfn/MPVRem
vUbZogfOSi2fFwdNptA56bduxUkGFVmGmd6kFoCYBhoiBbNBbK2zlQtMkT4sDnCV
8sSVux+9ke6PPBxeAwOdM2rodvu9mdbrD3WdmGF8xqn/57Q2QfX3U3TT/ivgEAXd
RLB/E+0CnVNdKHusowyIPBGTYMHWrHRlHLzm/vLjZ1ziYqnvoPfupTvr0PK2WcvC
9zmgan0rlJ1uNlpwYxHbD3d1DwKxQC9vxDhgfykwlt/32NEoIWiGZUhtfKFrL3qf
PJeu+AXql/YrlpFYOQpbgBLWaeYlQm06uh5Fszsh+AXtC+QoemHNJu1heBf/YA0M
RGDvuiNooQ/vKALq+2Tm2IqJ1D6Hl7UiEFGyFj9G+/CM6Ddrk8aAeRpEV4R/6ze3
9foyl1KMTQ7VXc7mLMAWee1HB4o2PswwMAuEI9u0WdKfMKAxF/+OEp8LNL7by0CD
QO6vU/zwwrTXj2gxfY8UH44hEzDJnJ9ATg8V2NJzDzLsfEri/cschUou7oo1HBHE
znIlghIgybPftsvNIuBREYR+lCze/L4/xukCRG4teu/vJgtt8zmEZ+mULms+xfJB
mLctIA/KbUUx/Q6w0lp35tTcm8dLToDIvvL2ZtwM4w8f5aRSCmQ6daaa6IAbKxuz
vbFTSF8s4fjvM1IzthxT4aipVWrIktuFyopIy04oyYTNxAem1Zc0DyYzLZo7HqPB
XDQcsriKzSQP+oONt93dOdBi+/bIQhC1sp9GyI+guJn7W0xaAB2U86ons39GRbQc
1FeK1fNeE+kDt5dXPswOIq2pCsetSyobTBJ9k3F9hHLhbKSVy9vGX+T2vq+Os8X0
pKLQfitDQhw2FziJF71gFViAOqlf/NmP2MuwmvyVCG3JgTyviBEmY1aZgoJzotZH
w6vla/QPiymdrFO/WwO4O+wC8xaB1Qh/2QHTTOXAsbxCiiAG4wA2gOxQQkEOn3p9
mtva1lmsoW00Oz+XQLKjPXfNahNkweq9Ueww2eOCGgt66YZvHra40OSfzL5ukgyd
X48aGoVfSifp0gR5yUDKVuX38Aank6oT0PUZUegjO8i0CVV7Xx3VDewcJ6APmAsP
sfgKSA5P6zYl5/3GPgdbRRfGIL86rycDouAKo0R3SuRsJ58uaYBiZ2CWYjO2sllH
lPO85BC4Bb6DIFI2CDgYUzVZUuvrfTGmNPFdRPPWJz2o2wqkzOKOfNuBLvTwVzJV
t262D2CPAX45ne92i/4OKU0rG/od5yuHukMfv3CIP+Wt0k2/8ZSrC5Oy8ng2+TT7
Kh5sa5ORKsy3WxzWKGa5HT6+5iyYYLrEf5vG7OHS13piHyY+nqHKh8o8T1qRa7Ex
PiILWz8RyRZ/fpuILw79+YJJA7+j9tUp1lVq/6jBWKG1LJx2uEQj6KhsLlWvMN04
MAX7CqiXYy6IoCiMKdze7+Qhtypr+6OvfwwBR2qii1cZdE0vffXYGa0IXf4Kg423
XpsnH7HZzLgF6ifOVVsuoJ9sBPwThTfx9+Vy0Nib2SAF0+Oiav9mULP5DJYGQvud
3Ao8P5zNSYUThBDSSGUTRK0GXFfRe+ESNFQIfbiDrwpYi0/g0fmqExJ4PPHnIBaA
bLrnvWWiCSSvJ4cwBS8K/jaIn4Kp3fWLGdIKOZCsD9nnOvHWEFqdKcXA5imTll7o
y5LaPjVLbc7OtMR9LrK8MYGIrKHjtPUkOF6gnHB+AMjbc0tYGuaXGBGg/h8phqg5
dv8YfuB6itqgQq5HiRYX+oNn9mkC9uj48CMxkdnzxjrw9TXCDpyp0Fq0RS13QZpg
FMYUAKyxSXUKjjp8PSEBhTKwAi9IQK575KPqeyfjQY2JYU2l092Qj4sfIHky/CLl
s3vffEjRvwmaS5zkeDzA5hWXrFyUfzmGIR9lRvKQgqNw7J7FY8jtaEH9jipTFqWs
eRxot6MG5vKdg9NHRw7N7yP2HA/DQepfKNd5fvrs18Fn+bfKFyPuqSjIWmZlYuq7
77e0ocEF0Rzq7g58OiKKWP+QlgsneDHiNXbTSyFcXtRyxBqT1JUXNthyKGA78/Bm
TtU7b7ZWcDmRrN0cfkjmDLz+MOVI+b3MYDTQWH1u0Q/OpgffjyroZiqbYnXDoplC
MgsTjG3yjLL6ltmbfThdrqTOcrfFW8eF4QtFSIJcTWcNx0Cr2Oa3fB2esKmdNeyz
j8dy00Ay4S71WRjHUj+pXLRUkOi0dpdWFFjsVrOnhyhqJp2Q6VpVvTf1apaLYaFS
tmwUk6wOB+/Ti5i2vNvQnWlHGbATtS9t1YD5ky/ZvMs8NpqnVAQqlW6yovxIOo38
jgDeB4VPI5H1t2A0vJP1KmwTUN5PsIPbJd+J581PE79YDOAoMZ72CxWNX2r/wYrH
9AA/3hwr/gqtKKFWjHci0IiI/5dFWtViK1spihSkIWdU5sPpGnQB4neBZTMgD0TX
8b1Ftg/g90Lf0uLHZRRlJ6Ihj1pt7QRLK1wp+PLNnNQ6KDe5j6tA0bgE/fXHyKxt
RTqI/WIk+HmTLjKyr4BqPQbF8v7ba1rfS1XtoOIStYWoduVVBHdlZeJsFNcm93VA
hfm/In1qN+Lq5mPhPcnsFLl3EKlTJaMurmQ4fe0nzR5RayiaxypWo+wvYuFAvlle
Kp/2iR4zVCQpUO0q07rzvE36QI2qe5+KzD94J14HdFhiSU2tArRzMIngj9BScT+o
wHVg9eiHxgUqZuVBKyj//e+6Fl4A+Su5WfASguvuWoNOqDSSJwe7m+G9m4GOKYUl
jD4hF82o/3rM7rXUcSCjwYXi94vnXi7HEx4iFrZGaHnL+b65T3O4h0TcwsDSdV79
o4kJH+zfCZzrWoC36kNNQcb3nW8eyFZUj05KJxW5QPOQ4Na0mS5JM5k7HBjT4QbH
2V/Db00JXzeR4P9yR4GerAHKM/0lJZFy7lqR/IdgEL9RRgEfDMQt67NZB+H1W1Ud
gauQxFUXHZ5BFOnOqG2BfSakr/SUSumJBajgXXQYo66XEqrA6mIRwyeLp4D1tgco
KIGYL1igpNTORUUWN0tWqBBsm4vyLPChhv9NjrIej6JvCV0/7iEVBwYjX57PWXOG
2jQk4KpWbe+KgVltnXA0o30sEEGNQOd+63YglC7+EX3rng4a+qoQC3I5ptLT8jBW
c1sn7Ouyi9Yqp+H6xn5OE3IYjC/5Fw1es2+EvZl2f3yC8pT83iUdV9++oz+iLZyB
SBoN7q75qIQJyoKbMerFkL0SX8ZX66kGu0hYuf5kmxBpNPQK4XBhTJp/+3MGwCge
13rCX9gZC9+DcYMb4f3U/dg/vXuAe89d6GORffU691WzCg31EE3xgW8XQ3ghFxdN
Ky8lNhZ3Unlbf30hn7U8VS+gE8wCiDTa9V1S0F8IPptgS8PEX3CalNrn4Ak7uzSG
gWkrUZBkBfIzjwKSWgm5mqmTmI2mAXnl/is7SbOWVQ6UJ4EOcNVqQTdYs2QHltXC
NBX1z4SCWrQHr9NJYBga5lYwlYgyxVehN0Xg/AjZtj7lCsfUYKvRlPUVOTT5yNPi
4RkdmeWajONE8DtylvmKyfTJ2qrR3Cs5dfqh3HdCZ61qqUghoq85Sa5Bn8/Q7n+T
Gf9r87PHJZKoGfJQk3Srrn0T3TXQdt0XRZqoYvksxnbIwopXJKRJMEUErfrkCw/5
Goy6j9tyfPf1t0yBasg21VMeUSPgt25yPNuAbPB4bJ5BqRG6/rD5RtGYwVuCP7w2
bgD0za+Gq1Tu7wEHaJQbs9bPIJnkGzgmgh6ZVCVfBTnqVdgOQFeHJmGLlalB+jk9
NRvb8XEgC9DTzuGB0RiPxN6PpV7KNZBhlMY4m/1L5mrzS+Jg1AF2UY6rj9+QIBen
QApo3r8x3kpUBYymOAWGyJz3FXpXQOqveX1vkFCK/KmMhdOTm4+txTqYcZIpEY+f
HO0uHLWEcbosBvufGFatrVehgyfv37IKLW8H/esmVl3zNz2qClS/za6NWQFC7Nrk
uzjwq1UNl+wvy0j7ezKURIxq06/Od9lI78rTIkWbgawOr7FyFemle4p2sbQ20YU+
3jeFTz6dENyHVJ02cpteogTP8bB3X78p4pk0Doty2oRtqEVnM2CaYyYRTZqzYVbS
yvYnAUnUQSzrdKtJ0sQCTRWr2m+6fPN07+ClnHfvia/P6FYx44YYVPgNHDOu+P5S
mK+AdYysdJPluGqXMJ/fCCbdSnFBuHDQ4IL0wAwr0m39zVEFLklty/dcZG2HrL0n
s7hB5v6pi3fDYyRhSZRLK7hUMcGUdDaNiMP2qRvmOqX5L7mdPqqTdOCG+ZFbZk1r
EgX4kVHcTOIqSi7F0kD1JxWStMEhg8KUW61/LaYDhskXahFnpDlILinJbAkAG1Io
3du0p+LYAiWmd3J2LV0Lvd2QVFbt8X0VZbHreuDwy/Q45vWzSvuBE915L3OGOzNu
kZNoSZlZlCLeAclRC/p8bXRTuoc/WMfs3GU2mvvgm3gMpokINd6imFDOGXBN9pAw
xjZFCVdyWozpqZo6thGLB+iP5t2d6gBmkMThe2n2tPL9hqWSuuJlHA5jA7WqVYMk
2gQTYMjCq3i25VgkniH4DDz3F+TNOwf+xrveX/qoa0lTsdy4OuBr8oPO2Rz/w+e2
0RIEaIA5wVbXI4xgTja5RCcsAudCmuQb/8L1rtdE4XS/Y07MNxdL/tZvj7Oh/Q5b
Xya5c37GMSK+2R7sauFaiCMQj7dgVloThsxTEkBdMIDVEHDpwr1Lt8WsV7ExL6WG
WDu04VMTebiK6fWde0ygc59yvzgd8pOUWrtYxKBbLpXIAvVDX476SNk9NhRy8aJl
fGyeZBJZwzJjxvv10GPpbK2Qno6C4/L0hceXbnRGYVW0xywHt4bfTXLWtrurlDJw
NrX2XtfaZZhHDwcBnaWc7YO6HPe/r8lmP3c+Wr7y6PBrgpPmymGvE8gj5BqXAyoI
0OOWaW2iuZNLD/OHwac+UzCn9R5gRqsUH+4GjAvF/HDg/3BvPZdTK5R4R6rg6Hyg
+e/dYQzcQoq288ETgyUDTbv7XUltttOP9ePoSFCBB74w53me9K2vYIx/wmyONtQf
y6CU0v1bEjBF4k3tWIgCGjNRWy2wOg+/hoki8GotAu0DQ5CdQ84iA54BRRW7h5E6
GW9b9YfVtmqqxfTJDFj1+Ba40/cCZalLfu93kXLxa3zNGVmrzTI9tpUpiP14yU7D
trfo4CiXTy0ycKKN2JSlNg0mCmbSZzLLoaSTjKLME9CbW+SYGxQnUgbn+5x9bMbE
V6IJR+J2xEFwQhZzN6hBqHdpDhYpflG7v5ngfyvTN08a6ucQKCj/gvZXZAljqU7k
dYG5Zkvq+Q3jV0y8BFJ1hbjctRtB3a+3TU8ZWEnfSRKkhFNf/nWsI4QYoqM+EDoC
htHIQrouuTg6VOLVIaROq4v0ZwMK6moIiXUddXvfdw/qNh1UEvKiztIEOL/pGaVN
4W3NeeoorEADv07tIwAjzRDzzmcbeWJm+l8RkzoM6dxS7xcJMKCv/TDqP2w9SEUl
udE7qzzlv42JZ29DL6MZ/QxtSAZJH06H3Yx2D/0gwBFOALkSE3PVGK0gGn9EmRgz
xmaScoy+gG6E2w50x8un2lPgFpuXKnVMwNHdfOS5oytj0ibQaQuDsrIU8ytpZjs/
w2xwd5TsE00bR2NiyVSeYIk7tiK3kgIfBkQHP9UU4CDUXDT0PNCIB7q0+1m/WiMm
ssUhLlE6V9YgLOnqwNKr+67PD7fymeEyuJ22H2E5JufZCMl26z4fVmH6EwI4+VIp
xbdFglkf6DeC7ZWR91QJIZfGtiBVDclPbfdhhWuYqOmQ6JD/bi1BgQULy7nlJuVK
mtS+DRF5pfol5x1BbFA2XuvxbP5Pp27V9/NfL+k7y8ngZCIcPQAO1OmQSns6uK56
ycTQ3aEzSS9rmSkUrjZAlD59JHqTIAfaHBznJR4icNvo4M9KpzB1wUM7fIi8zJBT
vq8ajqyxsRS/wdhriNxsZ7osbHafwUiTKdupwTA9QJJMh2NI375MZMBviOwJqot0
h4QMv1Za0XXS/nazdwvP9ElOQrgarb10guN2S6CXC2nxjjujACs2yAnuwUlW6XJK
JcLPhZ/djl6bXYEQLNsQVUtG3YUvpEc9S+Be3rVlxx2Ta/RG3LV3JVEcX4q5I0ir
kcR8nnJxcMuYqEQb5t3Se/mgAiXGz4qznamHJ/sKKeo7b4+n3+ivx18qv3PkfEMr
SRqCxhOwuOAPHqvDhwtVSLNsSwtOCuS6L31niMNZWlEK/COzZjBfYbiAH9aqmnCT
gkpoxOJLZYvlGoTyhZW2lfdIELlg24y2p5IvciapQs5IdPRNphOuLh/V0Lu10Mqh
iId9UAZuzoZy7n0b1/Z/eBHj5zT9gtuPN+sc5hQ4hZCrHtz8LS/HyGcQj8hWM6FX
PyJTDuur5phym7aXON19jhD8EwLAlG3HfCtiLXc7F4f/QCdtE9j7ccRbUO9tWWWg
xTXtWnciz9VhBVrbMi5VbXMq0t3s4L20gqo5GnXooryqF7Tp0+5wzxXZ8n5ORNmO
EdDSMajqINeOVDCH56l3uu70QkJhWHl/2sMXBGqUOWmAlDwTzzyJUiMm3iTNWqeO
AmyOp8wHq2SS5rvM8cW6BgdAEnW5KWSoq2FMXwYv8YiNMEISrXP1azqPBh3nJ1GZ
26HoFrdSUWIMwdLqo9hwA2Cai0LKZ0Xm1KCileLAsl/1wdttbRkTaiI5hWlXtLhu
Nn1ctTCKNOZRqaJVgpzO4mxXnN5qzbBbA1Cb4HFa6kdCDeb7yuyyw7c8AKC1lY2e
tmydbPMyKef8MWzBhLGLfn+3odxeQrHrOj0NMQlbtV0Pk4VBLTltGev2r0nkQwip
fNx0eO0fZ09Km2RPN2dYufhNgB0j23/BQvhciKRjtmGXSXxd9BCf2yCmhTF10UiZ
O/7Id01AE/Zj3RM2vJyxYsovrlmU98t1/Ep4RgdASbCMGpShTYzuV8XxbpOf7/AE
zyJdY8xg6U+c4odfXGhVSi0YyK+pqAhZs92uSt+3MGk7CXqv+pheu1DXhbBpXWvS
/aEcDx44rs15AqkeenIm+DCT1191Rfo+/kMQPsvMRjHkuVw2/vbiCQifAB2JihEs
4TAV1HBfpTH//+m13VLdAFeNgRMcEjQY8wJOG5aoW0W1ap5Qa9quBBUNQtk50hcx
fehUZ8rcC7Dkmu171+DMm+ljLJPaCE1pC7/MS2qbqRw=
`protect END_PROTECTED
