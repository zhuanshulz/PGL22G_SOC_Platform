`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qmOJR7h9yI4wdvxRtzUsLI+htU4F3gRiB1Aw61tzE1kl4dCNMrx94rojBOzIsE4u
OBB+m14aTH7DIVQjLV3QX6xn30LZv3cQMH+sx6IHxensl6CdfFOqNiLWSsPx9F7D
r7BvUqqO69+uiVYv18mTjDd/sf5lkGFPlklB1Nb23/yHWAMmxlpHrDiRYy9MdefP
dcmEvQVdKeQenvQZtk/21Kk0Z3MJymNguNrE+iXRBNEzMzSadFFF8FYevk+7/idW
1vy8NKqwte28nrJmDFkFBVAVA97IDCPQCzER1SHIZptGMnxM8rvqGDv1fCIyMwmg
P3a6E62hgcHsBpXLwkH2fz1ZxsSSo1BHgq241ztRDgI68SZ4TuExSbQF1FDVGisW
IZ/RA4QHgAnOOSnlPIpLbg==
`protect END_PROTECTED
