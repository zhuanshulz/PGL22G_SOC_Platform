`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kaC73/F3oC2twRjbjv6orAXA5t33xzA82foqCgeaQAfaGaBkW4mu5J5Ibf3JVzk2
ki5E82U+OhVhrw7s6y5Lpu028Yoblvk7rWHeUlqN5NRSx5WjhS4x979sHVJjWRCK
d8qtieamUbL9loTVgrp02QnYd+DNmFCctSmNZVks1ArEED9+/XuiAGAF6DrvEd0X
d9O+Hv+bRNfpAgxBLETSNgRSrynm9FJkXMAVhFCK+3ZGo+NltNicw6KmI52xOi0B
GcYtSO8ttlQwhS5aaw25hEFo7so75AqMceLnDyaJHPQtiALUyGBIPPPb/RACWGRx
BVm0Hiyw5XWfSkPXVLw7b8DGfx9y88E/BD6hkpuFHnis62sYYi6L+IPpSJZFSrBs
F31jmlC2vKLLB0QjutlC6ObGrekO38VJY7Cto85ImqjD4lpSixikUN+OjAZhZat3
oI4oBrLrw3taxzPSLml/gVK+OzHntCCKI+kj4yZ8ICKZ3EX8mM+ZE1kE4DGQLaEp
9w3ZotOiCDxrnfwOBIuRlkBqtikpqn302E2SllnwpR3vI+sTC0I9Mg9IGnWCIby/
3n5EHeDRPRi/Gf6XuD1Nqw1O/OFaOEUpBApn+xU39X9ub/uOETDdwm8Y9L+lUOxc
KZWyw6wpQsVF7ZGcRADl6WXB3rMerCQP8ZOBys9ZCBnOaEdK1h8ScfozfJ9yeuIy
dFsLAkOTgp07zXFkNsmXUyGAynH1vb6ekp+3bQV+YSVXYnhINC7TwkQqhqZg+GeS
ub3t7Y70/43a5vB+0QQJvQy0ymuutfM7buWAv2ia7h68Ui8krRwUFtjK5Cr4BUQS
ffA01uHF0cndNSn/KK0Idczf6QgMXymsWGn9sfkWhFUgGp7bqYzRweggeCUBdX+p
W1yOYjIFl+XJ5iYc0wCcCZdC5aKgBP/ep28q9xag7+6RtbRQjNszVJj2Jjzfb3Xg
K2j58Kzgu2j5ZKLGZcYoSFEjcP1Ri0OZ3C6ZGYYnqGyU5MJLbe/eLnDWP/kiOUpY
SoRl0GW3t50xSzofpmrNbeA/vULdQIdP6WyproKE4SfPcjdtnUSbgtj5RXzqXA8M
hUKGMJZPg8e4DlbA2VKucfiQ70NnDq5jLqEU29cFJlUMaVjABPPc+O5F/vt13yPt
zldmD66MqkpzCv3AF6eAEbOkar1p3pQzwtJQ3y9i4dcYON+YbntqtGxmtdmVvz2s
5ujWB/+SUwiJWkk5yH5j9MLjd0h0IP4refMMkzH70jYwDz9SoeyCM/UA51XuewQ5
AB3zZHvTEWD1Y8HD22qNay9wNpJwLH0yZlVlu3hg/qRSgkFNBIyk9cJQuRVF2Era
TngRH/qHRGNfA0MFMvVebj3hg1mQLaVNNMwp1HbF8V+DM/Xv0m8XLPTnk7yU73ei
ifinObVfqi6ixK3J2fmafC8S/33d/VAiQ3zxkn8QsXt2lvYCx9lGo5MKjzOrNgNr
9kvUc9tQIVjrorzDcdD8q01pP2egcvvwEjcLohDUN5CrBE+0hIok1/Hf6Urfe+gz
p65cwG0CBros7tQ0FrGq4VoFz2PmhHedS19DBEFIQv75XPZd8gCxhKrBgm3VvNG5
Ixm1GWP+WKyTV/lkpz6Y4vbg/XN0hRdCkDe/nt3u8WlPjVYm1yAh9DZ3KwipC4D4
GWOOSEYvAcBupFaidHqd9jADn4BWXRxjcofUIVTeGzSPWqQtJiNGCV/SczBZ+ADy
Me7mnYGrC81iLYVZbiiyo3OA8/qJ33Z18Fwxl90uR8lmub7dwmyY4Zn9ImzGeGBr
PgyupDp2UZfwh273nTYQpSx1bQiPfTdFe7KUYVurpQXGuiNC4XXlZOT4fVAUD/JY
g06rcQY89Kj+b7H/PuKBx1d51PKG7+0BT1fu8iUDu4eWoVBRiIlbwZoreOZPcqVx
qZ4O6xUk5lVmZbLC+EAiiSHLMXf+keIDWqKx8TakLldkbGH+2DRXJzfDmw/BJ3jj
zpI2yhynpoO+/DPfS/QIufsJ6mlESwhoSVIb7YRcNMlHO7F5OZwTdiYyU08OX/A1
YaRm2QclnM5VlJE6xI0sObMEBsCZaYnimYnU4xT6iekyCweUO/amKjK6w7wexKwh
ahX8vDAX171aWQU0cYr9IMAEmxYUFytZzBvwYyt+9+5RrAcyvAJbCiiCRAcEhVtJ
n3qi1TeKkyI8AGKA4UQFrtbG5Nkijlr7vZJQaYXvV9T7mE//bNiPfmYYTVbvgbkq
5n1nqDu2qs69EWKPe9yFmjA6uVbG/U8uZwTNlRYLo20=
`protect END_PROTECTED
