`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t8T3X1lOjBX2GWsTk7ukPTP3LXwcKR4uIOIx3vpw3bWcO1fmmFZaFuYuV2lMRDY1
cEuyVuR9hs5WNi9nrZbQJXp8q8Yl6+1IQO2hgPOJvse2b0E2jZPGtWQXVU9YRG8e
Aw6pUkXoTp6fR5khj1Cw051R4EBy1/wpFaj5qv2jRUBtZfdVPj8GjSNdBJxuiu6z
k6WXrCxm8hYprDlwBVogdsXsedGBsdHtWXH22kDEon10B133VnjJuvwToQ6QNkC5
rjkAQ14Np4d9/i7KpQlw1FSQg3Sb9qr25YZPtc9lTO21EcUePTwBvs9U36WXZOap
N8lIIa7A3Z0U0wGXtvAJVSW2IWLp4D6/jNj5hSeQ1RWdL4YjF9G/IsukBFdp3QmM
mFP+NV666ceR39dRIcGy4bWo1oFNqLCx/Ym/CqXkO1RKW5vYpCtk/+O9CoUL/5uK
RuySW2W41MrxO4qOQ+OhzydMrnWx/gr9+N5PIxcLFryxjX6hleMwVTPg73DR/T2n
bag5Ph+aTavTQgNBmXmmIKrvhgNY1airLcd/KPCeMMI=
`protect END_PROTECTED
