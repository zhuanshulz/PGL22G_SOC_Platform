`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
irEBlQeW+0rM0XA+U3JPkTJvPQnItB86n/CcQsf9odvSK5VA/DPQtStgaC59ICjv
udFSwzDF9nZXakgGEJEHzs/26TaQ3pXKzFipJ6tNnitR0HvxQTQrG5MOWmjE9UqQ
OK+wIqf7YSWASyQZR1w1BLTnEJ12SDuXvmp4z0E2vDke5kivnTO0dDYKaoGsI0XW
stpeFmNh+nx6TOMFioMvEz8B8xtd8HLES9KFon8ZrFLargFBWOZN5imUwi4d36HA
ZvQsAmIJoo4JPXZWkJ7TbyLWdiBI4aO6S5A4sltyyV+LTZKjAGDUi5VxXS2s63V8
rSmX6NLWPnSNxNpYj4UAnI8vdHBpH/wUTdKCdq2YyAO5mTMtDv8cZY6Lmq2jcUCV
TmpBfY5T9lff/d1ofckduhYNTwOPLbpXLaZ/myQ7TrrIuExbrHb5PmZkCq3NwzD/
LpcltHbH97tehXMg52zKDijHALvgADNd0FaVHorU4pIHCMJe5ACVZkPqS2inAeDy
04j9EOrYYHDDXtRp23DfP+Lhx9+lYXZacL2F48vfbmKxG1Nbs74q95F6GmHMvYgq
3zx730Cr1nJm7A1Tur4AJUBrk8zAZBz4zAoln9+2UULwmvGJtTiUszljrEfRkb+s
Nle1HTeT2Tvr1HPebDjY4Ea2Eq2Nq2JFd5ilX+CndpMINzJ+hd1WEI6RBqOzjnWN
9UUFreToywtTlbuFFFKqLz6KF1mCLmb4FfN772fPgaawVz9Avemdkz3kgH1SYDtz
j8vvUJAu4VvCHr1QQb9ZeisXT7kHRCd1TblBNjjkvxecP87IbMwOdCZFFbdW+jEb
FWI9+dWjPkb6YpXOsMpYSDyKQ2l0SL4AePqBKFvdD97XRoExFs8aJTM1Y0Bu5xb/
zoFqiJ+DjPCS8ritYYCVuWyR5H0+ScSqH4vEp3BWvhoq5hozQSsOEHAg7Jttd7tR
qwsUskOf86OLqOI/9B57G9B47IutGnkMHzFsKkv2SApdY3ybfTcx3V5Di7xG9imf
BNcGUQFuCepLzsJyDOevNywMzsRINyEYPkRJRNI8Gr4lkKzZmPr+uqtFXh58y6TB
bV1LVpa8U3xI6vlEu2VCy9MlQShR1Vu4XYbhHFjRMGWz9rTUh2oGjkUpvn6pAW0u
GW5UICF2LhSq4Mca47sHZAe4J6lZ2PK/um+kapK79WZ39j/ZQ1zuJi7VhUaYKIBI
73i9bEfNOC0bMlKp08yVQhHzVJq2qdviMMuQ/iaaVqN4GWDeoLWt2wVYxFgykU1T
88QjXHTa37gAYQLmLRuibYQhMye9uoOLER5z/yOPkE5FYVcZTDC3opDxxWUltju+
iGJ7uJ+VJ87LLnonPU4FLHQCTU31YHzsLpq1vyRXGDRd2QFA7mT0aPidiysud9VB
XQwjQo7WD8Waj27CvBq9sBxpF81LrM+DjXQ5zUV2GFPWeSvr1tOV/T+W6lBMSkph
6SyXUbNJcZjQ7P5lFyDL3nW5ym0SiHSb/ePiHn+D7I+hYuzTXCoU1q0/RJSXC62e
ZyIU5XUC/C9xIX3RO20Yepfo68KFOy5nq3HTGmAnw9r29z8JgvigJrk5mzQCX2h4
1gF70PCuwfyJMsWNujk2YA8o772v59rRGgpupZXuTxkqhF7G5IlKXOwmwIIZjsee
CvkZdQzXo8ub6qNMbV9JUu7QJTynL7iRE+ABqCmbJRJsojdSCv/Hsr8Hr0c4AtVO
imvnr8k+FwKocaVCjfpgAeRDelYGdocMuoZbJ3uj84ry1RjB0/7M2wnh5O+9xWrl
AHmW+byJ1gIgEV9adUoqhz7AVCNssAN8zRm47As8QidyNuToO21aPiT0nUbYxInq
SZu59+MV/c5/6Qx3bxPI3ODqrXcp7EYFdQST9tvRjNwf6rw9KmQcQ4xUgT2ffb36
Xx6JKHvQe8ATCPDcy599iAW2CjPhwFQG7yu+vKVvqL6x6Bvs1LmVhH8tK4nx6MFK
uNwEWVtDh5Sdx+4lj6rLbfUkZ9L1z2k9zVenpOfJkpzVbr6cZjzDEzMgXEBWzcMU
BFbIdROqkTDNkU0IgcQNfjXThd7bO/Cw+m9LTt0aSMG9Wcr6nmAaHx4nl+vJ8x7u
pS4/cVajle7NlThE2v2GjcxVQYHI4lLc11T0rmXkInknomh0UEY9iQ+AIj6XlC2r
6Z7bQVNXvfCKnqvOAxHCsc/pmUKWrlwXBTjFQnDQvsoWo2LfyQq67oWibvyY1NYx
Ke/qC4VjdLv40O52xmjWJUSCwUnOfuWRIucZwBRu7DTrd3UbCMA3wnvwD8H2Kln0
dLV9SwBmlWBd+jY4mLPiWvXwCWKzbmQTxuyHOt6p/NNDpIx5CGCbpN/bYL39W+Fx
29xyggY8Ut8NoeUPAIVRfD/aBqlTzxBub2fVUbnXxVxmHMuFSDzP12b143y0ECmr
W1/QX9fyE5Mxy3IxJgdfZPwKdhFSsQYCDAaKa8NXticxBUR9pZt4PvDLHfVRsGCf
wnSGxXvM/xGW+Y2zJDCrU5k0PSdkNH6KiBfkE0ZI/7nl7cAbgq1HeFCGkuy8+rk9
DY3jiXFv++FSAD1KOTcJQaQsgZrJ2lvYfEiFQSHUVVuIhsfw8qrisUK7T6+E/F0X
rQQZYbxWwJ31CJihaoJgfJboFZq83p2Qic2SJZ4iXeJfEneMmapjdId6A8Ep57ZH
7sB3xfVHas9ZBYrlwgt+tqO++BM6mQiUISRF3EVXT22XBq3kPxdL69nuY1OX3kOy
AS+7RviuVbXaskGNJYS6TerX7WFFZmjw+OnbResFLJb60WEUNoapKycZ/bTgIDVC
oePossYr9gbzW7Mi1EamuJth2PwMA5MmYsQJJ56suwC1STuNwvPP0oOoWM5yf0lX
aEeROGeqzNoj3KJzpZqt6SOVj5A/qe7vL8RB0Qi+CqUpboQGiqtbzH0EMIAQCAs7
uwRG46dHJUg4vKvmax23N2Q+9/xOZVslHR07jk6nmIqnlBTYnvRK1Go22XfZQJbX
4nY+LBckhOOwVe+wgQTRlSLN5SpwsKSVP1w9LcYh0Db5I0F5S0m3rT0f9Tl5EYBY
pu4vPAtP3jpV/Zt22dyhf4qbQm2FGflKvfjiubJ6tOkPTGmSxynd5pHRzSp7x2r4
ycnlv2vIz4jGNRJzJTvoaFSLd1qOFo+833BGD6T0TBHT0THkY+x//9ZBpoRTnUTK
C5jxJusyTXWEqBq+CIOirvaU5P0V6iDaDwGsK/PXwurSz+yInWjQg3jsI7YR3Txm
ofKiTZ5pXWMKyGEZe7/d0JT1oT2px0Jxadbvo7EFMy1/ZVCxF56apTnZzmq8dcBX
u6KJWByFjk0pWjpw+/P01rUEVeC0haQKHViUxaSj4T9geqyG8onQTHMnCtQ7b/a/
VdxCIMNp4mfCseMqnKWMioYX5nsSZmHL+hJ4yXOmPBLzfcALSichRbgXB8SoeoxR
lExGcoOooLzxZ/rHpH6T/MmIEWmGM6WDKhUQqheqXoBH7KUZf3QglFA8a7f8OLIV
yvWi/DTUnm7U4PdUqpAdxTpFktknAyvRngycWE1anbMjQSTMQ5XQ/4gChl0BZSV+
U/g+RfhmSLc9NNTiv+HQfbw+fHMi9I0b64oV9IiPF4n5AS/4DsMin/Xfe2xdxC9u
sdltAyPnTan+jUKIWRc25Me0ghsn9IqptCP+sMdEfFzkRdPrJz73OvfZtNi6aKSX
HNEjIeeiwo7xdSTigKsFhCE0+zNLlcMVpxKEBHPRO/Bfq6bcvClFNdMsaN6uYOW0
6mLxAje/6v/C97W0yPpmuP7nKkatrPi6pkIr5f6b85dyyP7ooVIX4ydjpDJlxUbj
kimBGw7UKmFkWXMb72pvaaR1/2cjYp64759/fzgfJ0tVDiV7syFRXguDJPAec6jX
qxh5U8V+2Vtcq/+G6EbO9F2fore/QzGJOhbzyJqTUQ74bEC+S0Qpki+XoWjgf5V8
HvQvzDtoWVs0rDxZJdkePQvMNuRgagpMj3BFMp48KYxoipC+QdvbUWiIiH7HcxpT
ismRpH+bIERtzct5IiPruMkJjBLoSsxrDnXs+Cc3wFzHDbvjKAzFf62NflQEIaZJ
4RwecIpDRguhi1LdftRBGJiWofI0xncReII0hg5zR+ERwlvVoN1Sdo8kiWXi8oea
diGjesOaADDq1c5jzdtg3DmsE3Jh70e/Rny9iYbGodyidyrrC1e55OSsMJ4o0Gdl
C/XRMv76luYXBwFDxlQjOr3MG8Ul4X2mqsc1EzOv5NCiiR3c1OQn6Kv1DbNV/4lf
pmPj1ZHyxWNzdqM3jS4Qcz7ZxNa2wkACo9k7mZI4lsy2OeEVEDNmsiALzX9WQlnp
n/2RaW+7ls198hBitnnrjVxca9F8TgIMdc7MZ2t6YS1pPQk1GKoaRArxwhkwly0C
jVcKASg40tCTw4pYjBXnbsPFKdH1ATbma+UhNiJwzWymT1WlnQP37ikgekzOudpx
QnRg3R4kBH/C+eplJa6ozortjo4nwWAtubuyr7UdXvoXm3VBRhb5PKXNPJtUmx9N
Fyy6pftFG26fVUdT3O3DxQTIiIlt1Au3RVXS552WNv+78Ok6O7M8xf0CL6Io4Uaw
1rIbXoZWi2JbHx3+5g3CzJ6Lr9WuT40PonPnC50h0stX5T493GkChiAKPlBcZbVq
bIl5KHOZxjPvUq06eUuaf8+ahoO2XaX9a1eZW8J8cvMYm+OVaOjb6vvaKd2XihvM
LVhPq846Lun00Ayt3dOjzhSdLHtDmpNUd1QMQ+cMvpSvHTFeMjIVAxvlZINwVZjX
OXE+ryAp4vDdYRYM8Kp5N/kQQDfISI54ac2rKsbPU+BARzhbwPjejJAd5G/Hd+De
X84yT6cF/1b8P8ruaOxCsaXBC1djH4VxuLx+OL6PXlBX20yXLshHtiXhQsQrc6CG
wJWTkF46FObfZI1UKNqHGtiwSjpacd4SBnyfxlV8kZMPieGchtJrAYL3rvSa0eKe
2e3e9eSX/j0KJ+IJGl57xWy1Kmd3kxvxx9T6Q45WIkZgBl5rn7SR7dygnxQ2lfzT
VNzlkKOhuAAhen4vRS6MSInyILzeMpauWGLIKTZmErJ7WEzM5NpTnUZF4Z+QmCUr
Br5NK8SqfQ00PRykU2hWIoPPalD9gU6S8JeZ4M3hw6C9kUM4ZOmI4Q3CriBfwDQQ
pcKfNkQPpWGwbtBB6IwDWzz7NW8lNMsoqhi+nJuN2pYb6AsstqpzIOpBf0DtxOQV
P5kBtB+pAoB7c0PbAuv6PADIAjXxf39zIDugHw7dgwP9hAh7VDGwBmVhxt1Yu/SW
7by/oIO6N4e8rRiMplPuG8R+mhTRi/IiHus6oCcxsRGp107ZsahMOV+S2XItyaE8
7vPBKjD0nOC4vc86sURIGdojuwq+7sEoXwg1GHBa8AFZBQpjfDL8LQXHRFSJRaeE
URG225GyPyQtx2wbLH9dHew8KR3Ni2Ro7ovb8lYI+dIMJ7k7FL1l8dAl5owixW9t
2J8myDlffvJa4WHO3NarV1zsEtguhqQigZvrOvbuToDvSuZE3/k/+ZMeFGww7q/O
96xsfRlWB60pi/ebVR6GYm6kJloDN5NZaBiWVduiyobTu/HnwYUH0zpgQVW59vyM
/AS6EdEl7ANkDxuEqjTc6WMsADx8v+W29ddtu/Ach7YprlKN11ta4/vslLC22TVm
oUxwycyeFWovER/7/WigZJHHIrktKTVUgp9gw7NKacmUpux95Gn4c19FrLLBEquH
69DmnXgG8yJUI6P+hd+f0aNDXGalFr0Zh/tdmhv0My4VZ568RHineP4H9FN8gLyM
oRv0i9mnGsIBjUwpfiqz1sd4lo2stUQDHwdRq91RJDCTH1fTwXJc/jXiAXQbzWru
AXB4U1xJE1fpj5GwmNNE9j4Qdm4zAUX6tPS6ZURdSfN2qaGGscJ935nRmEDnRd/E
KRDe8Qar3ROBQGij07UqIpKxyuQWPZpWkny8JRVRmJZBBB++T7n27f06bTIGobz9
UKwSKKnAU5ghVnNQJsesJ6zxeTqZz7KHBgqZ8NgV+hfx4UFH1d9p++++CZiohlDU
B/nB69MVm4Fy18jkpp2xYM6aQWxVm1rxjCaqrAT9SMlUiAC0Rr0r3Hb8Csm+UvtW
vM+u0cQI3cUrzopKqTLsZwc8bMP6ubP4VSyrY1Ag9nQ5fhonxBn0TS/LeUHYTCVK
jkSzR1N8urMf1O5WT/xUFJJWmHOYsK4rHEfRk15ppS2c0T4h88/Er4jqk5u8M6qK
nEbgKXT/5MrbXxCqCSnouiTvk9SL2z02YzievTXEO8dxJBf+i0MYj7b6VjjUtdUz
sW3i43uqA/XMq72NkYEiWJOfNR6vFFjZpHY8FR/cVAZHr/G8tYYZpl1MTGnl3+7B
pve/xwom+XcMxIMBDI8LyAMSU6K3hmys91cS1h626d+PzdjxELJh9IOAP8QpPKJB
PBul01SxhiyhTQZf0RNYWDZPXdo/y3Dm9Wo1JxhrQ0I3fvZl6BVUuA7ec/8h1HW5
EBGImVi5YB9lMW+5lYOuv84EvHzkWAwdmyTjthSal5M9M/dHoZAGp6bUFTi5deHP
WVlD5AAVIBVB0mBEei91mKBZxhpsZBnSMUYVDgJIwKR5CvK32I0znnx/hHDS4XK5
2TZG+lDnecSxJoK7fsnYh9jEXPUaUGPQOPwnFTZjugxSoyFbKmh6pi/s9V6pDFDk
bDHLirQnbQA3r43hEAJA7pHQs+K/XF2hdmk/WZbfZFO1xoQ9Dv4jPcaXargWf8wu
m9etDyXuLe4jDKAYyoBvT5Kty/y2Ll5QO/WAeMLtktvgUxQr0GKNvvWDP2wOQx6t
sdfFR27iEcI28U+S6/1NAjRTmM1yOMeeasu/AjFRXIjtoqf3ueZYE22mVULye1kI
nCh+WAJR+D1C4EEnv6Oi6Bn0eYugyM1qDTNls2pY0xGO2rVdFAppt6yrFPzrZaK2
J6wwCNUzzmJ1sm911096RcwiIqVYwbGHjTnm+xr//ap/A5cjmfxNDp9Tbr5C9Opm
72/xd9QFN5QIvqrQNg5+Twv3GnBAEMEWAPYpNFtAn+bnKDzBrdLgn/XEAn0uM80n
7ucxbdg+EyGkOh+7u4cDaYNIHRrUkh5BcuAcs3b1Xa9M9x5R6rzcqu2cBIIKWigo
1EBKatG5HM5ZGecxKvotz0oeXhsbm92Z2Zbrbk0RjGGgSihqPFkOw/SJzFcLmQtZ
6yWTb4c/Jv1TYKD+e6DjMqkUD9yQ4j16sHglTNhOJ7yDyZA4UX2eWoBgGXwmhPqy
8I1HnuWFvP/n/UufTL+ZelS6A27HHaT/qfJBz6n0VcWCyMMM2HwRbfV5CyRk82Qd
dmEAgaYQDnEXQkj5H3XPJMrJJAntQDOe5QjKOTli5skCZ5XPeTekzqC6rjOUVml6
Ofp6U57emoy0MjeJigdrB61ASkHSvkeygk45yG/r4sooLvNs2J2EinaLSK8Sqo76
ia7FP7jg3hojL6kdvxQT/VXoiccqYr8NvL1XOcQgmoSnJcskyECWVJNpuSy0+Nkm
LaL09z1Zwj5kltMdfqS+l1djLP/+Xz6cpgyI3Tbq+JKPOOZRX8xip/bMg7ej5Djv
R5zau1KBiFxWF8WvmC9ZuiBBzm2O6mOaOgv/7Ujtqy4toMiwPdiMFABMONMZGO/w
zsOhejGSPqOBJ5UeVoppTc+nRLkja7nxQG6gPfBL6h7NTtBhn8NG0wPqE7NG3GzP
oHAFqKaq5bt5B4e828gRY0FY4se0fnUx8zBF2xntKO7ly0MQyz6aLqyG7lop+P69
s4eotfRdSg8fNV6HL4gD3n1c3ZeIi6W3dP4E+zeezXgHgX+ZYx35zvq8Cv8huF+Y
Snw37YelKZStW1fJDi4cGmNnbmaPUxUp1US3+qI5RxszxSAsxoP/lIGEdjuBDTv1
nNL18SSR9yAZlQlB1VEffPO5+OnJABanHIM6CyUVJJ9/VoDd1bDe87A8u3EJGeGI
25zU7Rr/dwaU/szTkfOgO4bIY6B2fjHORf6ySC32h+4+Z+JVauQEExVClulsF6JF
Kp91ttXNOCN8kXFmBPS/3Tt8XJ0pCmywssOn1svaIGoaC7KDX87zlkFMydDxLN9D
sISdwhhCBcrFE0jK+zj3+rPDsVlZ4eMEYzh5XxBhAhrLwLyTQQVFyV7bZWxtS5s+
8Z5H2CsF8UVmgsekDTG6YzJX3MgXogW1D5SNrBQWXg6DiZ6WPdaZ8CPDLL3/l7Cm
Qre/2wKwDHeOnqZBw/mR3XQT1pFGCsE9EWvArtb02kSVzkYlSWMy9xCnnPa1qFt2
T8yNfFN7HZENpQlTbOmpFsRoVTwc+3Ru/MdhFKn9PxvnrD2rYWR9eEq7hpZDhZjV
MjYsSts9Wa75TYkrG+505zKOZ4u77JBxbCY5EJ81acdX83sMwTErWjM2sJvuqvGM
25X8R2Mp8FZ6H6g+iktBEMk6gNYHED4V4Ehsppx64XqMxR7OZor2eLR5KYSr5nE2
+NiplMiDoPe4G34r6ljSHDUgmk7kO1sv5aBpTh7jb7CIMdWC09NI+mga1JmZ0VIF
Vrh9bvgsETzQ0F4KW9WMG0XatOAksIyglGCH75H8Iixf8L/jYgTqrxvOOE4hLcF7
5O1gNhPNbzC4VRhi2EXl4ZAezQ7SAz802LxxuqiyCt2GQaz6KNbivLNvRD54pcq3
4dnfB4LjrWJctNzQnj6TZXKDpA7Iszw76MLJfMhYOn6ZKU53PYsdi0bRdbnrwYHR
MDt3YQEpU2QdsCMrhIHC9XLAIFedCTQU67xi9jgbA1BS/bBDyfEXyunZ30otpfmI
yFaxMnSxzfeumlLQixJCFR731uubt064WqqaXZFiwmPaox/eBvnL9rdjL0DxmUWp
g15eLhfpZwRHahdRruccCDFS7SG/jKVY/HUbskQhFEYDAJFHy1STEZeCYgRFf5fT
+E6oCJ7+IABcbM0khX6pSY/9x9zA612JboyS6+hhh7v7SY/lmmsHhwnpQV807Xp+
i3Oj7LJNrdtBB1s3cKaqdH5y9S3g4F2Y06EjBf4mgdn0xWapro8rZvSrRVYr/5kU
fRliZSj/A0eCt1ft4YY9Iby1o85kGiB85CsLFcMid2m6aYb9AK/x4MbPCxhMdJJa
TCc1uNfgRGVURFk6iHKOkxKwmIEzTOulsAIO49tuba5NFXwWCVmi3VMVC5/AXKes
i5Uqom8WzOBTIS+69DfPhefMcGRZvL9Dy+VRGKQH18J/EL0NH0y/xsjQbGP8Q4qJ
ujY3OXvxziF7biGORqfT0Cx+2n6/0+SIXeVVzgD1ve9bHcxSSJD8CS28p58pBRxY
qae/pZvA08N3bHWOUrKuqFdiamDLc+2Js+drroh2PoYgfle1nNtk/3TzqeseMQjx
vCGmB19fp90AW1x7UGsx09ODFb5YZmA5suSxu44/DiTtI8mMWnJ2J30qit1MA4Ob
fnHirTZAiezDOeo6q2EQmRXWzb8sLQOG6LZHqxLSNxASaVr1JDv7p42X+/M2SD5Y
+B3UZVISc6GYGd75m1Rxut4zsi2ZOzHFZqyh97gppHd4u5Fw0lx/DfZkAjMwfx42
WK5oK+B8W+WL6aQtEQQmpQoF0BBbmPdx88udl9n9CK6cGX3AzZWBl2D0eKdo+ZZI
h7H2lz/ER5w4lW0wY1JOlj12D8klet424egkO43CG+fqnmCHJScPzwiAc2X3l6k8
Y+nY9tFWgplzezKm1B84cQOJK6WPEcJkifpWgmKnAR/G4JK5+gMs9KXNE85AABDp
TyaZAubuah4IljpW5Dl30Y8HunTUdls1gxAuPQxHwvx1QVoUgqhUf6HhOC5yT4VF
dGDB5CnSfpsdAempVbc/VVPBf2377LznRfnHxRGRCiWHKOQr1DEYkZ31OVcU8obX
78DbhfoBSFfPA9AScVXqY1jWKGeE2GXjuu8OPfxBGsXSb+ofwcJn1UXvaj+lQ0z0
SntwLQCjuWpHk51JwvcUUc0E94klIq6Bm7RMnJe99XCs21/u5YSIuU/kC2JMRqdw
ACywdm6JYgZfTf0hhGSiXU+RHrltCBABxcMeGIkVkJshJeTMGpXnt2FiuJ43cOZ4
VBxNz8ZmxO8CKr/ZEbVw1AK87OhKn8XzkV07xwh/+xC8WQF9ICoYVlT2SWT1tZwp
SzrJ+oE/8BdMZXAjDID+8+yX3JAOdi09t7ctMqxxUxmkUtIVwiBSZPT6t5N/86TM
S6Fx5q8zsWpYnNxZ7HDs9dnqIPiLbDcjoAsRO9cQWi9oZNmGZJwo0ym69BG5BCio
RPIZtEMcE7yhr9lchSZanYbOuxXGodL3Vg3bcJRxmC5hzC+c0nDe0x4tcQK26/PX
Vl7ZA87yHXT4mc/SFbpXJPelxspQ2QKxjhr+GXuGM2Li4eFtgYLenUcA1nDft3fC
KhbM5wasoRooWhLH5CH69M5Kng45COGjrwxBp6NjsOL7ofJPI0jz0dDzPGMCxKqr
ftiRp33VT6WLp7lpg+7FFx5qjUrFx2Lhq1SJ6eMieN4BDoKm2Vq9citQLTUN9Hvu
4ONLzOLx3JJnp68NjfD7T1ZS3JfQR17X7i6pUyAGGaaCwktft4m7gI7l4boXl+CH
xdhp0Zt6xQM3O6mXSiglz6TP78tWQDElc8n2G7OJRmAO0skrrfeyR4zkUgnIznYe
4dVvehuSVJTx8IGJ3wUBpnW+qn0A1Q+cooNAGuYY1P3Lyj2p7JmzxwsyP3CxU0hR
XKvXd/FHNC+1UC9EQDiAmhBJjsDGKT2w7YoqDFszibWI5N25JphPnXdM3B6+FQSH
SHb/bLgKiz7s9ygKX/9x1yoARGLDqq+Fw8wTDXZSKXtpmAH8x53/vLe1xalWT5Nk
kskCL0MIU6vKOFV0ZpQh4LGPaaXQ6tGbTcSSiiBN6NQdzkPYpPDkVyb37cj2RGgM
NHItfhe+5wgiJDh5G1Prw/2OFxz8GdZb2rWWpdsz+2c1DfmlCr6Haa5mKejpsIjW
0TTN6MeBCUH8bZPWZDG2ok1iHHpmuRtye5mlMOWjzG0pQSYls+tqal6POXguttyI
c7iPSTPDAm6Y15gL05A+vnbxMUe3P4ZxRZCsDCz9PiKTku8cLZYILUL+GtwKjJRK
EuFzim307EF29o3igrZIARyJbQPGTqChnOIyPkJ0x+nHRjQgyPuYm5vRTR3sJ4p/
fV3Q2ggGF31R519yp96tVVgU27ZE7WKIXb21iWlLR3qpi6semDV6cjoN8APkI7Iy
ymgGLEbRlohmwqaxF4nw6Bz8yS84gMDC656q3Vbe9v534AJmsZyuZG5rdMdAgqsT
0jZvIgPRSS2GC3rVJZ9vZ01ZRC6kkRPkfsWdPCWTY/lA7/3P8UQaFG1JBndhW3L+
fQZtYTGcpRQUyseChr1Kem+E6JTzk/1nWVM1IbBHGdR5T7+C2i1aBx7dcH4GU0kz
0du1DKRQB2OzIM74t5bUklX8uMRqjyOw7i9OVbhD6+b5ALTrU1JaAyeqoHSRYCt9
1cMQxXbzpMmfbpxDVQIuUKjXFOETXcjCfkoQ721XbWDG+cUS6uejC47jurv1eETM
caCSCiktCVRHzkwJjJMFRwS2YeKJuHDuK1TQodehUPDoswXS12pssGN84fekNkIN
ehXTshb3S2OomjCxd1z0knlrcpspFyN01MC7la4vtx9wkhK+WXGY4DPfdSkj68v3
CFRb9hdwcPB4sYiQ8uu5NIgBGByawZce2+s0rw6DRhjIWTPMncPQCz3wQaGySGOX
ihODiwboSpMNT/1VM1aMkfmHZlWNhDxj5wMdhW2i1KbIPqyYmEqByq/pxrMd/uf3
KV9sNOAjB93QmXmQb8kkzV49x70Gk0lc16SROMJEgFHUyYRJ+Q0SwSC0rfEhckwd
ZqGLoc5sRPHwNRTqeuSqfKmGH+F9o2MKA8QVGTDVelcXCOu2fXkM7ms2vxFU+bdp
Z+CLbRhydnbBm6D0LIGZAGdlXL5hGJMJnK+erq7J1nasXLwobOhxFbvL8Zgvd0Ko
kCaev586SlEFfhaMKOTqr06Oqn2sAlzcUrksClHp6BHnP9KWOX2uJEIYQFMCXhxj
/bQrtfRWHQh9wuaElyenoKGAUJar+EEJNEVTAaLI/OFzKn1nEZR9QqT6jjIYLWN3
PM+7OsdeRC6zTf9z6gEr+d3oZws4ZDUy7WMC89+JMuFm/9cPWznIs2FtuCf/bOyj
Rd1tcqai1NgCE8RlCwPIbuTzq/I62dTlhwRCtC3IN4WKr9cBaGJzrVbVXSBo0bkd
wD801abo7PPYaAQNSYd2COUUzKeFHwlX4Om2RZsIDe0RNNHtIlCIgs/dJ7D3UMk+
B5MK7Xbn1NwasIEiNlel130YQe5hNRJ4gVoZKpnq35R09QdbjxBJEpqaWGjzm+L5
EISI8kJ+t/AFIPYyWUkw+2WKsBHj8+4DZhTuVANqvrK0YBg2NrVeZefD6ZdrZ7Ba
QuQ/MD6OSk/l2GbIc6wSbPJk+8e2zy/vCy25GY9JehEN05tQ0+0YHB9E3CSj4wlD
gFpn/meXjqTe65Va6mgBCE9dYRz2IL/oMPou78UWea0YgPlPLUD+aCaE0qtui4tG
YucbWlVNvcjxjghorZyg5WErf0qwi/Nmc5gJwz0HvPzypvOKSfTEo7RE5YNwjWuk
oaprCWsgwhQb5gzR5p6V3ZgATkt3o0NM6ks7c1rxi9qWfSok6laklhckVDeisfM4
sn5DpFCiqk8jukXPc2uA9w==
`protect END_PROTECTED
