`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dgrFOo4qc98YBuRdEYkldq5h1HJqoarYKy6f2ogzYgcp3pxZSVxvxHskGFuFdLqf
Pq61doVzKVTGABd/1/4DbyX/mxbgp9czXGt/2BXGYLzAGcpZbyBINF+2BQwysISl
AADaNkVXeAyDmgqJXx+teQQePkTD3kA9WP6Dz6trI27UW3veuBs5vGHDh/qy1l81
CjsaTJbSXiNIGN1oEOXhKhq2Up8zK2hXhmSPDL7pQlhNWObOaeLExTzTiEggRx0g
aliUj3e1aGHvkDGqNePe0MY1XlSmJyDtfytePZqqfGra43ODi25xbAWy9FGbrn3Z
1k+QhSnXshPjvhZER5HUX/wDA8sSHCsSGuSAZ+3XHPJBJa/qDlj2ELUnfJQ5xd7P
AE5opEXX/OU50+eCPk1Va5PNCNY3ln81UMBQejfhKwktIwY6IVHYW6pqWKJC2MZD
sg8P6LBNcHCfr/MSEPZqf22CgoKeHh2MPnNumvYEfv6ZRHe7I5ceTP3dGXn29Y0m
cmTQHYdfGeegaxwkbttGoNrS4LIH9d9Y+Qr6X+4SB90Erq4+wpLMdJrYGpW3bETZ
jcGYI+F3x9baopdx2Z6R1r5rWd0obM5ys2yYKUP6xosQu9msYv7Zlz/yZPKsXaBN
pV/+dtXubxEqhqi/nSR+wEFqH+bRJskYCmJzxY9OzqrJXESoQeqRRi0EO4Dt8aQY
`protect END_PROTECTED
