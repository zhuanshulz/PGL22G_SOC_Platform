`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gxbw4r7H+vDAFUujURCPaoXedlPQZQ6a+wrO4qpgp6CQGuWX5TBAghD0XtDzQ8r8
QafG43DL1pNRO77uKvIbeeuXWtzqnbSD7MnWc2lSkV7BZLzK3v5QrGxba5Xe3PKE
86sMh923on/K5EyKNN/RSGWMfgu8dUED9YyUpTEUzw8MkChXiXimTZYtf300g3aT
L333JPpFDKEp4gUKHTcmy7f/6Q09G8Xz+2/2/pMm/N6C9ezDNd0TPKnUGWbx3AYX
1wzcgdjpewOX3BnJ90b8+GIEUGGpUCfUjYK3LU1kca5OZL+YMaMUOtALTlcE0192
mkeIH6wrtSVcjCRr6OfPgh3QdenlmSNEmlkPoVgGsw8o0Y3yZ82hTTpnR+smi69T
pLgUkW4/zgN4WggnbGb2LZUR73leTOpkwebzOuaT3I9PbMUNvXiSzbU2aXXkioFh
FwpsPunQfmEwHkwgokXTxyelw5PPhWqKA1a3E0cgOedk2xAcGSIkW2evPHOihNcd
8TvXJflBYqp+3iyKHphvW4dlTCqbhgpAziNHbBkKJrYBGEknGZFjciWy47OeWdAl
3a15/G+rP+pqnbn6SIH8pGbaQudnXXq5JsRNseZPvCOk9utITD5h89jLh1HMBgoo
uXLIOCfTFoKQdGtVEiZFSxnGHkThc7XTzJajO8Dxnr++rrhLO/PHXhLHwy5gc7tH
qpNx+Mf06fzL4hT+eMHPZulvDOO5cyatJueGdMzwgGHdYGdAcscCJ80gD0FC0Mac
Uo2RkqhDPo+/kSjbc1BCGiDqZ9mW+T/P6q1NHYI1SN+w20C3kjx3zK6h0eNdVlI3
WXfzZgj0u/2YNjL1V6eq94O5SLDaeWhC4g0oi4vs8mrcYiQOHExXWrgRX6PDQ6B2
aekbikiGNKZ9xjaj1LQw3obT1/ObxjupxOVlwbUwffkZOx7Wx50soEC1v1MbCxYx
jh1gIjU/fVdhP0W5eJ5eNZaRbfuWjXWZJdh9wQjou5AcRNg17oSMc9YoLt67JpYm
aMiaxjlWBqEbLaJoGTbSl7qrBjzMGVLv0au3tfJNPmdiEiCTJwBpij0CaWo/X5VV
X6o0I0Uo/oX0wjXEUJm9DVOS1ZvfPe2gxD4EGyUj1lwiKCbLY1ZtD7EK/seyPcux
4l2CgH7CFzH4kixXwSfJcUr4UwcRO7q0rUiYz89gzx5aIpw2u/twLnAiX7QdfQqM
KkixMJ7GAfc5S1ZoHotg1eV2KzEFM86J0B97R82ARt8U19XWJ5AQNus/wG5UecVn
rWNU342DU0lp+Sr0qnxsu18vDnk39KBP12vBr7ZImhFaUs1ggyhzLX+5u3ItRYff
XcBRzLEe141ISSDy/hsssJUSFZLGw1+Qpnm6cmuW5j3O6sg4NOnlv+1bH3wKeaMU
Pw4PaMlng1yzkgGffkVhTM+zNe7H5ptnNEls2qxHmbnPiKGWYnzxy17eS6XyG3BU
6q0cdqeG9OFSsWxxFV+SnbIjopfx6kCzBZ4ShtiS2XL9aUXZZ7svSC07SBnqNxnQ
QoRCIVrhvvIvq3PZJzNpVgU6hqyC9tPzqm+uXX1maKgnoOoO96ZVFuCvLBYL74th
Qj5aupb5L2udmvpniSqpXpjR7wr78fsE2eDzEyHdiuY=
`protect END_PROTECTED
