`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CufHYd+DNgF31dX0irzLNyLv3oxp0c3RsHvvLQrcDG7sbDjlW0sVe/jXfSntqTRm
N+evMCbBF8AzI4i4UtLqbeyY/J1aoMj037Gr8oQvyV7ni2J3TOy48fsPs6m/mz2g
faYPErF3OMLDTTuBxiLgzfCwVQ4sD0eE9fLdXG/5a2g7257cnnzZRq64KEparUVQ
CobOethr8ThyU5UN3cW0lZP3HWU2GdywvSdAVr0IV7RxXvdwo+ob/2rl3epNJPK2
YnmKivn5S1DjxpzRya5VZURe9J2VehcD9mOiN9rphuMi2pJApKod8xw4PRdAr7dj
yuMPl/Df86VBAWpLJcTMygqGFf0ky3Y+ZhkXI93He+LHZDuer+vzZkBJ46oKV/dS
BAgxe6FTx/vZSCDgbUxru0j5+Sb+YMZbGs7vIDOp6/oFdSfY3vWvILeEUXu06JpZ
LfoGhwa6rKtraTtBDtz26Ve+sQp7ahz4r5lfTBe/g350g9LMWY2elpAoREKRR2B3
bCtRWx/4FLPrlTYlvSGM4EHJheODDOLtxcxhwDJXhB6YJ4Nqsz/zdaf794zRjdQk
Yv/et73OHQzw7ipXt9GbQlQTxBOdRtKEXgPEnsYbVt7mCqIUfimSlAZaIRpn3n+J
hqA/jXOa577GU0ALu8rF0A==
`protect END_PROTECTED
