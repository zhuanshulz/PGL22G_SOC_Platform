`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PEW+0wWV10e35hmmMjojhlCM02n0ZRtzUofjWnHx5CAAhlv+YGkzqdmMWrg1C3w5
AK5lq60s9M+knfQ62O9aWNKHBpgrCUZ+KM3RR76BN7d0wQ47jdSBLRiX0I069XoL
bKwR+zqOw/M2OPH2jnz98HNxNh48QiELJVIEShOe6KUtKDtYjhpc/5u1eYF4fxp2
JGazKQJDdW2ZDlQIzcoYri31HnIZCgPXSTDAaP9W1zVnQqObZjbHCd+y1ouCKfmw
iGNI6orw0hoGWHRHH14dV6Q9C9ylW4xGuu+hQT697Ql1LCQNGYkax9LeRDKGY5SA
QssIWYbama/4j9Ouhqi1doYJvYFE1qYLlkizYkmRM/tjyenuHEo4Gpf/V0+E4fBF
zhXxuhO0beuE5gF5eRj9jeXIyyBBzQH/CwQ6Y5Me+r4=
`protect END_PROTECTED
