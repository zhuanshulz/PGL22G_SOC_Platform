`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aYLGwEceGXg9Sm2kCxfFwmA6+iINCxODDKDUn67JkrIbzo4aqa+1klxEsRqNPbGa
NUgd/Z7MpMtFiFQ/SXYNiuNrabcOH4nzP4eNmRpJLdLV+Wbj845TnX2LGAq617Kj
hRt9zKyb/dgSWoKKbbXrsUrHCeU+vJc6HnVHwVlZJfqXRuBSSi9n9NIbpkaYln1B
z5tR88UvRnh+xgEtCND1FEth1JNTNRrRkU9SK8QD7GXHrK7xVssNUxlb49+iltQE
mmOhZYXr+NgQ0EIq9ssWw9fUskyabB6fyrg7UF2iIMk49lnqlTQhaTmsQzlRRe7W
3zsMCQIpygjOduMrUMFNF5LdpJpLeNdrCJOKaGWx8MFpZoqNfbaM08KbIruETycl
6ujbe4dDlD2Wrb/fDaT7hRFmf8sTHfYMmRGQWDzRpVynbs09JLYBZe1lCppwv1eX
+IF3ESB/d4Hy0ioNUJ9c4ehUcRqJYiIyu8KM7Loor9Ts1B9GbnCcyR3N4IuwM5ZU
vKsYzERrhgIhCSEvav3tOvci7lnbc78YVi906YGMxVaphC2ti8U4cmKRInvaAjkI
BmIcdt4U9J5z87Fs76c8VdkXRjvETMEJsAFV93hMSV3WLAwvr3ODoRlJG9talUBN
aT1teAXZLhkgNM/Uc+lO+5/C6WjmvjjaeOykoM9dzwOjepeeNTgnlC101aspWWn2
b+pM99JdHbNQBXb2HYjxjLsuvOFxnoCFDLq1RQavWM4NZFtKFkXG8BB9PGgpIsgH
+xagh3ROR8mpQi+ziLvOzMCeiW7P0OOcdo4LBo4xqtVAkCiIqQ6BlnF57e3iW4N0
e2Jc5yE/sAttaMbJElqm6I8oXZ7xbIfb5MpGzxYtLJz2pfuDZoLgGqM5sQomUIO5
HbldWbjhk9fjZf2Cug5ZFGawFTvpNtVlR0cNAI06SOGaIUgdVGOk7Y9jfX7Ev4+t
jTsZANelEVr6GFpVYb9Og4Jbd9ezlEId0XHUdl6HcMkEGkqzBbOjgn7qD+kQGvo9
cbbduZlytVUTkAR2QJu8nctv9Bnvvjj+NyUVk/iu8ZWAdklIUQfZfXqvwbaQ/N0+
PQJup5O02nVWZvtnFRjNui1IUUdQVtcaeyL+WVaJUT4JTB1eJHuFOW3+mNaywfNn
2i8fb3QodP030y504gEDOEMiO1BabFMTYD+iWwknwqZtWh+PQCvY4dZTxLNyCzqA
LwnYEBtFsCta4AJQs8X6hqzf23JfRhiLtr61sFrAwXSXN2DrCNY1aStkayDXp4wG
FzvGAkVX43ILyrcUXQWP2g5LGNdxWDZ302+y/y2NN3fzw8SH61mz+EEjbt9ECqXN
g/uDx8lFWUq4wT4XDDYRrxdFx3/zLUyK20dUm6XlVA12vpJnqA6TaaC6Wf74knvh
gjXeIxpuEdY8Ijouf0weI5ZIXxHBx8Et+HqjLTTY3IGKgWHwPR98N/XWMNDKNkat
2Wc4T7x+MjbNbJEU6of2DJnq31Z3K4GPDo50D53x1XnECwEbQTPOVp3JUKSJxBO6
qbsAZCqtDHRzbyQV/1cyH8h8WD+gPJbbf5WC19tEsonPVIt+GPS/E2PrGfmsgpQU
t07uCEPhoorcwromuBF1szCNEIIljKiui+loIaaoZPO18eaIg2e7L8EMqX6Z9NnO
yspdgzo1HgB9g3NVOFIzyBYS6xigwfvBT5OlmrrdbLNNn7GRpnY1N6bBwrP9+skL
N/Qaa7l7rvcfn/uXtFEnkXvkBCbQEhjBXfChDVaHkpjdyttUSwY4oFXLERvgPRdB
EYqTgeuhCdPNNzrPzChTAaJEbkMGOGOdnWivFEt9+t8bGdwlNAHspRlvVB2BF6Qr
PixrOKZFHgmRtB4pxjFDbetp/6/8Oq66wGlNgXEMegEo3BJMpjOK4sd022rWeTeM
1SdB7MsudSGGrCO2dWbVnpgGmOk5TfQxP+xeMbb2VmMHyPBFp5OemAy2TboBXyAp
/2GHQNTJ9WMq4ghmQQdd4wm3wJaRRdVD+7/5pQnLhmFrt6+H3OjCjwg7TqK++dSe
FTdHaejHWliZfeljXTGeWSQCRkdW+dgt3zcdBvqqxA/k24E+B6zTtVd70LdTsh2e
bkXEZJIzXM1EEH1DGEqj4qkYDJYDf5ZMJuVaCsc/bd9jFCTjdW6PKEqQFpB3FAkw
6v0TvO/t9EUVXtbIWHj3OqEQG5WXcHEqEhZQCuh+frIAFqTz8hMOME35vFI+7qQW
NnneMInAw9UPMLG1+9urBE0nITq3oeknAAA5XytNHZCxKlcOgKWkMZ/Y6gmdJ6rH
tlggxLENgJLj8UD1ont5YPTh0rGKrs5zdVvQ3ot5cAI=
`protect END_PROTECTED
