`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zahDlp5EyxsXUfiS83oZkrMqhR6Zye+TJMahQLk+bTrXy+/gNpECNJzx8kZXoWrF
9YmBEjtuSwE6svnDUe289Nho5uxG3DG3k1EaQP5CuPxQvE+VYoSMo0iPQTMn/DTG
I+L0dS8mVoM8XDUQ0hn20o0YOQcTjPExm9opZMljm+Q1oJEvASlrqwwFFc7wDme7
l1t+8aqMUwgUrXlhCuVIdic+saHlvPd4ajgXpnaB5PBS60iTv7Qf50vXrABKQvBV
nzB0U6gOl7v9APX9lPTj9MzPsnVzIjpWHOWuFjNfjPuMsmnF6MEZQQGAoOnDcanq
mSPPxAnbWyrh0PbB06QFzJkzpvUvWu0ZMqGU4pp/nB/E0g1F0jzJ/G77TkXx+OsB
Qc/SbzqI+efUO7+wsjBCsGiDIJN8aE2x5hinTkENsK0+fk3utE2+u5L9R+WAKAgP
B1xQKO7i8v7oW54k/YQf886Mg1VgtE6ZiK6N4MR4ZqiepsS7H7M/DWwwfdtwoRpt
80ut8J0cDuVsToAmhgjUiEphpuaPhhgFTCFJ6/AVoMDdMzaVcJhaTWERR2JimMzj
sPQ5W3ynW5ZmBXABMYO/vg==
`protect END_PROTECTED
