`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KSG+17yutop3lmjOpM2VIwrXexbpIicKL+F26DM7Oz5bTa3VkzqepJmosKigccRh
3s7AbyIDZ15NL9PquoI1bHq4a7pNwoPtJ4XhtLnZDKd5lTp6QfmM0HOb3St7JWWD
SrmzS8a++Z6mYGlKUAYBSnhscAaYeDpgrfSTOeA5QdSP3pqBhGyEfxrY56SQ5PIE
esKRGJAg6gpbyrXpcmbrCd0SGiRQQHJ7I6z/lfs2B+fE72JTUWfCC8aNhBxctwhe
KeJ07Un0/ENgc7jkYHtfWRUBkR629v1/z6w5LzLHNO3zaoNzoR1tLzPNCLg3gVS5
jyNOvSnGKVENoobeqkzCTlT+ysLA9QGgUcDH7FxvmX9g9/rWAAxyI8NCpDlZYxvF
sPq/wRmSBh2y8awb3X6RaKeiqw5y/2uyiOEQo6bpZx8YvElhBzrfcVp2oj9Bibfm
VZckOn/7vMLnNEAB6rD+p7XA1ctMVSm8Ftlq6YUZ+Tkqvyz/4JMnIrJgZL5eYvFw
X2GzGoDjt6wpgUDsiF/97Y/xevQI1DXzM9/ssBWKb9+NWsB7LcqdKXyS/LKiuKJ5
Y9s970NbPaUkBSZRrZpgSaZ85V1hTANiuUwPE58OB8lmnVgaLQ5i0tfb6hBcMReG
3m7JlhUxtARoa/67d6xO48JP/pLVRDGTpdMMeJk5HY7hfNgmNGjWaZZVYukkAdTi
IYqlWCGy7/qdLg82EX9yNWLde3MuvpBzxzVwvhdcz1s=
`protect END_PROTECTED
