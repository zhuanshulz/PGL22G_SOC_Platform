`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cDilJFteIIh3f9rRRzaWO2xESaVeAcoCfw9/XcM/x1X3HQVHPr58Ovw/WTv0svkF
F642hmT2PkkFCqYXAd//r+Nrw2g1gnwM0v6lBkuOqZ1CdXqiMKrFI0f9V74BigoA
KyqjSfj3q68kkUuxz0ZL1SWKM6YQLsGIit464w43VOOMtRQOwrMSH0hIq1uLKJq8
NIV7t2aCOYtIubywBMcHtQaA/PsYwNu3S8Y0+YyoGdnHW+Nx23HZThmZNh103rDe
/bMfUcs1TPJ9FIM6qxcakVKIZF/cIhqiMSqu/oJI/OrTG9pVu85gnF+ehqo3LoMt
b1blbPizyMKzKcrMlMmy9EOE/jBefooP0rI92Sw+4/GlEbWP509MUo4Bxdw6jPSb
LJK33tLphapL4FLMpEMipQHlEQQb7PRQjEg/CQql9JpBYWgIvPzpe2AwCZgo/oFU
sebdIVFSbl/alBVmyaoeGb1GmAAbT2ScV/FmP8/8nZ3MBY2oumQd9LKy+zk5dQXJ
/01+7qq3IXvck3jEViUmSBCV5j7LDYKPKHcl7GG0bmZLQs5Mirqoe33La0ZlTyiS
rqPEslB47WLozmbt5uBCzyivUEok/XJ0xIK33uCao1arfCFTJCI4Z0ioQC6SeN3r
dX2GrLr1Pg3LnNq2nZe0uZ1Ay7lFYf9TIi7IGIW6P6hlkv/pEZxlhn6MPN7VmpBp
fBT4mmz2hddPTFbV3jyW09UF+YqV8+azo01QJaWkZNrg/JkZRem2pVNBLGMJYnbD
9eUREd0w4RPvRb9tRRdhZLoyT6nZ2BvHbVaMaV0f/8sFOpCMU9YBWJw6z0N8Q1mM
+DSSr57XY/uVZaWIZ8MxYnrl92kglLoC9BjNUxO+4W5/8b9+erthKSE0GmpN1JOC
7o6meHE6FZBC49SQiCwkp/fqSxvQWSUyGsQ274vMGMDsMaMnGQpCtbjKdol5QFaC
Nq0DITpz4gIzikOTq8t9L/kHkHeqzEotmLTEJMAABTZOUJtZAg/iIngVzSuSEvSQ
QYYpP1ctIApaqkLGGybM8uxi2e0JbSDFRFN0SpGFyFoLGbw3qOdZ4mhHZcA2TVop
UzzOV43tEVbQZoMnhBrX/8nV+x0NyVkn5fyyo58qmbMK1RnCjRt/pPZLuSE07M6c
lgF7O6NkePSE565+R4er/Zgs2Fl13xR4RL37eIMcIZAoVtwH3HA+V/MKXuBL1mqk
4J4VaEUPyKHjKFY4tIl1irkYRPMVBXQtE0YaSahZpaZR79gUrGhWAdDj7oUKhTTq
j3/BhDahbdpOzQS07h00q1cE6/PiLPYHjKHPzzDrt5SfetCpKTuH1BXQ5+Hpa0te
jGckAIcZAGyzttS30lodiVkmeNJIIxMaDv4AIN4Ux0d7xSjBZex1H/hI/DOke8Qt
AoXBfWSD7TP8YUwhxIz/oMvSo4aUgiBVIE2cL5dHfmRzcC+7BA3LjdGl94h4JIc/
dPqBOmTHtq7qGRtxKyLfEDvigcYvOLULL3KqEixQ89Xdk5lvsU6le5qLbhfjtRHm
KvaNsKy7IkvBdYzg8fFFxQ2gOCJloQg6k4JXBGSw8CIAbzA5SXI5qrWLJGKbA2Ip
opgWkUoAThftBzwxxTuIG6E7weitqMLFGMlPRROVHVnh6xv5g1uTJBEoWRiikPRW
dn44yX0YQgbx4dSj6+p20UpYUXz6lbApL0awQCLz/1QulfRqXlNcMIXJPSltDM73
1z6PGEeOSeZC5JEXE73sUGhwSLELfdEqEEiXcTo7ZJFv1yB3Qwo7I9JZfK0Ed1ye
p8lE9KQsXfbHeZWMb7xHt6hOKh0hAXEqqKSYxe1w1uC5/0B0HbXvMlVnvYizcvj/
bf5f15HW5WgxgBXsW/VJo2a5MqzPBrc2NPc9YAYSoto85KdOIM3Tkppy7s7L74eZ
R1yBGBLAldTBBOXzj584LLGxHHyOfb6lJv+0ThFozF5fC7zDlOXhRwhokrWzM7Jh
PlfG7vXtGKWF6AJ3O+Ag5qF99Q4iZRxQjmILtPv6zIWK44dnHrfs3tSqsAIDSbQD
7SgF+WeTdbOrk1dVoWjJ5jw+a89YmrDmBWhX6Y2u2vUhlKf8HQ7SyLbMpbvwMJgC
V/mqScjsefMjYwWIicmRX7iXMZqEG+l0WXDEfdIUplsRjMiOJEAbVl51TgBVzG1D
owU5EiENA7ocxE+Vd+4Ar0O0CSyNhZ1eIs9apbxFZS7LkKQ2rSClGlPQe0y8l7fN
Ut8irWUmZGsXK9UeSI/BPve+F2MfPeVLC3Im6eNeyDyHupWapJKIoa5xQNHLhf0p
LS7OaCRPIrrXWBNYbNuh04MRtmNicM3vLIL96IQqO2XbiM2uLcyyPqoDXwghglfN
UN13T7OLsGUJbL8owlNh1CSlTJJsYJlQRKDbJ9GfEff81lWe7hIWKRjbJTD3xglO
s2o4iLv7I0xqsL+jS/QSUI+dYBXNFHn2+oaWHSK/kAswXKsnyPhVo/CEzMcYo2z3
ircHzLZUkAciezk/BqAagJgbyzrWttc4LRaXippqeGII4w9H47nCwTvDx7U+kfNR
cpNZ8J0WVzslcJ/Zuz7C22p5z6/cS/LfflMQ+LbYbunBwdbjYgldKdOe9qMvZn18
CV35ZHZwSqEadjJzS+9PNpoTDOEBpNeHrXA/bXSgZd37o7aYOzoosXzKQgKBGin1
4rN/HPE2inoIQ+uJskehpqwklNGRfzR5oLhmB3YSXLHKBLJXtsRefovBE2gaMxsN
kj3EjR+kPqf/9beCxSlcy7a3tnaOuFXyKtNd46uBCJUgPs+TCtHpuoyPlKfZRs5N
Ck1eH917pw4yyrGJpL4tIfID3/qRRVEkAfIvbtLxhDCiNPebFz+i8EUAeV5t7zNZ
S/Y3m7np0PIuUncfZIKWwkD4rS5UnjDFsj+64Y1gn4egUzzJchgqQ5YZkRWp69kj
vwIz64qxEnKBrWRpzwF2vVnxQxUGEMWVRD2UM3+g+FvE3nmfnKhWwvwkpUNlrMJg
M09e8SfRmJ4Rs0TOcObHjU9idkzX24A9t4ZZMkwY8AQvy1uWsJxkcBYcUhSHXmuo
tPfmNh+kenlczcRfYMx54SU8TZoQMQobyxGkUO2Vi0VBOV39z6eIKgcTJeMuoEI3
aQnvbk5qklCQd8KhhZq5SmoJhr/S4X/ij5iKOk1HlKqrzNXga9oS4Xca4P6E/tNY
B3p/XLav72KSzoPi2LQcxFFRzlu8rO8Ak9AYnc83EiHqSRJ88RTN/FJ0jCHwbOy7
Rt97FWTXqyPpXhnlcP2cEbsaUi4N7u0TSy3nbdKa2VL1opY1Ve4N4b/VkIU9poVf
RArpKzyyzuOOG9qoIWm5tUgTji1S2a6lAidL8xsJ0bJogV9cNpclOuQ8JYFirtSg
2UDlwsN+Lee43/gSxDE/DRhL0OIP8SV88UliDMPGefbCtaEtyU6X4AObCXujStJz
uGltCgnwEn+m14ZWz5ls0GXIGVlXZpXOQl1F2C0RuwU8rBUIyqMrsSsrMwrgcsAn
KqoDSynbW7RnSwpJNVS7o0D/y53jcAODdO1L3TTjIwaadB2Y0LlMPTfb2/gcO5jD
RK2BA+/Jburghw+mnnI17qkjJXIYaKNFmmrui+tNMnEUKXIBbYeUY7Fj8jTA7sPA
OtMr3/brfF6Mq4L+987MZ6KM0y8+0vpQ1TNc3zLJEWGMordzCd9g2zsk0QqYnJ45
ath3XygcuJ6uLsa8nkLVAfM8qIwMaH55DBHiyLjrjebl6EnEvvxLbkkN9vGIRPqE
j54vIOoNCY0zWY9vkzx1v2fDsnmO/TcRPQiRv6FzeAzTazb95amTKNR8HS5e/9ap
OXRG0rWpAnyBkADRVzfChfvn95qfpkwXW3cmXOryANS2Df3mrBErDLlRgB2YFJBq
Gf1uuXNApQMcEdWwzT4kjozUlzrpwuFEJEUdCFsx29r4ypvnR4tgNYfKS/VsKM0g
m8lh8vyfpgDCnSKZ0kBtvxpmv5JGGQyL8hDNwtyrjNHWx0cF6XIoykb2cnkhOtP+
IQN+Y/CbjxslPX35JhOxX15Gba8nchMEI/UDFWmwZlmL1ScTYjVNLl07wnUd7lrc
d/DBH927TXqthzOqHOQ4Sw==
`protect END_PROTECTED
