`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ltIYZnA3ji17cnm810Sq8ECT4lTriRpe4BcQNP3n9q0X/ceJb9iKAbDqq7muIYCO
Qhs3DUM3oivTlAQdLIp6p+GanEsjda6KyYFcAE3sD9eeAr2SckSJ+OdT3x20RCWM
+z4H1F6vDYtKK7hup0FLcmFiTvObMSrvfMeD6e7KGBOYdGLr06ussHhfz+eJOlim
yMcrEYW8vtSFlOhl7avcLrYyi8O39/suQbol8n9D1liumkuTMBGZFDUlGrq3n93J
ID3IBOGK6HahcQrHoPasBiJDcnBYgkmT9GG4RvimNzcCk3sjDb1l0SaQ/lrU5kX3
E54UFRV/HY0izplG0w+J4aQANGN/an3PK3Yla7W0O0ILuXeebxAY5RVTXPOQqcyf
nU2v+XVpeVvlLk8fjwy/YPbqzjtNT8SWk33TxKjyxaAwAW32DsQNspyVb3sM+JY8
BwypZBDS9gFw3yLWcAjkOsFc/Ls26N+FiO+jvL8aQyH52n9jB6aC9QtvAFBRz3Eg
hDE1EHUsp/itkhisYpDkZw==
`protect END_PROTECTED
