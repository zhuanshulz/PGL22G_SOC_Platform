`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SHIBVgYtnSMoVHrCRo747SzEQrbtYoOtV9sv6GkrgGD2nS27eeM7m95ni+EUZMlP
QPxCEORKALfV5SLnHGqYHzUBnUMG0uqouMYIbvk1/Y3Uun8qvQ+LMjNrysS64da2
8k8rYJcI0b3GI0gC1os9kfmlkD9JAx/Ry5jU/2y8wbuzSp4wn9NM1XLQasQgl7OT
0y7Pnm5jAVqDRQqG13Pvplsu1BkWdUjaJvWWRwWvZQSzk1ggKJfzgt20q3cTFg8n
fk3QMmlEzmH08c7LzC0PP7AJ/OCDO9FXklGBY6WtowhjDn/ICy0hKOrE8Gt8KYoE
f6sP2bO6WIhT1UnEDtPc9jFYhVlOlYyAghJPNYEH8l63trqyh95cqLA4nPD2kXg3
CUDjfNBUmkfA3XRwoiMZ2ipTodV7zlrjO3Cne0AikTPV5KdfW+VeTaBszu7AiaRp
U4bzjMcl0wE57OCy7YRRSedDqm8wnvE9QFeuBBIPw/hQrMUiBhqwAq6hh19HYNDF
qxkTyjOqrdsh4eJd1dIDO4w8Skp47qn9/aNMklBesNyi5hiTBSlWTvqWmfb9fxzc
VaI7dVQMcsgKnXVREbwxxOSlolyhTf/vDwEFgnAVe3l3xf0c7UORDcnZqX+Qqi8s
/TJXZt4Ai32vfWBj4a9KJffaYGYw74Qr4u1piDq7Tt9pVAQTysAKL0OtDL79GMAi
W8u+biI7iZ7RsgiqcX7EzP/BlssuU/BaTiyekr+OqBPQvXphdpfRbyFHW6Bdp5gB
d3kk50zmuGnOr8V7Om+t+5CISIG53a+JVq+8Q9Xx/Ann7cReW6yOnTqesJngGfdP
xeKniv5mRWMHp34KBOEwCWN27DPcLLQ+cgwhCB0Uvdkr4bxSVTDYumSJWX02PdaH
tV9/rZmr61jEp8NfcNu73KVnF5gvE3dcAZO0F4xc94daUk2T1cBlDuLCTLP6wXm0
0mTBSN0aXeH/G35GlFzQNtlFVPKMptQk0P9RB8ol5IskLyu+Vqlb2u7851eSX/KC
PWUYACVMjBjwT6zDNlGjQGtZ8Z13erJnVpHDIQdhR9o=
`protect END_PROTECTED
