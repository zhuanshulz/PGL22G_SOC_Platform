`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/oR9vEw1CM5B7LRKZqnGg6D6EuZ0PFHzys6jTtlfNLntaYg9DpjRHSMCvMQUvY3H
M0/kMfKGk3sAkWlbWV//oHWgAnsuf1foast++aT1f2uoEGHSR9ZmsVXOGFprChbc
LajDKHjCBR5xmjSQpo5LGvYgAFXl6XxBp3Wn8qoEQsiyifWPgH32IcamGSvEdbHm
2aj2M8O8+uWEIwWZSyvY6t4zyObYT7UGrfBTDSxMI1O/zJWu+k/V/uEMj1tAUDQw
IiS7Xh4dIY0wG5yoKjlr57Xb/Wn1cgqHc+Ap/W1SYbfc5qU9XScUMaJS4QnvDeSW
2zWoFpD62Jdydhy0OLcIiA0XsgEWOWtg76DhYh9nhwxZjGp6hokbzCYlSNpYqpIh
ORXnebanRdwCttAnLqS2LlMYa4HaePv/O6DO4h63WYv1JBi4gs2FaVKFOkscjOor
GG7yXa6YyMPJeoUhJjG3tvynPN9MEoi4lYWY+96AnpzW7rbppxyO+Ri0mFLoBCCJ
pO+yH30DgEvEtGOPQHpOLMzGb3O1qaYSUIUHKkRlvA3iEzZ0r/hjxoAeKntkZOpw
gzWPE3+1bvtIw5/SshMvd4gzbegN0HwD7XsllTcLM3YFE5SWg5/b2mlEa9z1I2Nl
HGrlz5noB+Qhs0EXNovxis64WU2F1TDs7YXO4rhiMs36aSpSduGl02iwR56pqLoI
vCUZ25lWU62FjZijOP8xtZ4m5zqd33kxfQ5bHgdqI0TcQyVfJJ8rooLAeL2PheH4
boxMEMi3nFQ6Ze25zKRBKxAvLgkeCjHsg1YuRFoQb8ljlxpwAGZ58kZM6REKxbrR
W7bfL6kpzSTxbPZRdteJaNH70RUr+IkDr3YHw8WL8wwHaZf87QO/pzDS6SyHdHDe
CsP2W8bGBe9wm0VSte9yfjqEiIrzU3VyYzttCZdJjtUoBQBeEVIbt4TxH4700Uw+
zN2gz5fOK/r1Jj7TSt7NVSp132Bv4okecsE47ZbYNeptIU7GQBsq02SG1DK8gKrm
4AUiNgBwuQaZ5fqH6dxkdxknnRqWY1wK2UjVmk0wSC02AH2TM0DvdRgpf31VkuEA
Mu6uh46JkOx2pJ1gDMZ/e0pqJ/YQKjGfg6WI398jSWOPku8eELyGKS8eV8v7z6/R
O5bZv2qQZSHwHF+2bts7wkM0Rx/OwwzF3u8oIymFDQY4xu6hDYV4DJ9YXiTccsp4
4MwU+gwbgMZbJeyyv/25LLFq5lqcqP/9nflEXm2hLEk5Y4xg5X0D+yG0D6OiP684
vGvZcmJGJCvQDK+Lm8cdK0SQ0TnfOvK0CaM/M4mQTLB6K3yikhJEfkUisUbu1Rr8
YffREPfgwMT/VAfbzb8IxFHjal4abfbAtPpYJ8s46gHvQ/UmjzfiohD0quWPyvJA
u88MSXbPrLIHO4GAg3vsQevSIOdoqZYy8YmFSZD8YOk2f5Jv4vYGthKzXoOz3H1v
X1gkkawTqkIDeZzs1UzTalwJrCESqgkZJzopgQFozhrBoozFry3yQEF7QULinRgO
05zDKWdonagKfUqZe/0NDlPAJ3rMfDshoR5oKauo7tA/tX72mdtjK8jMUjPBr6mc
gnO3G7Uovy/sc63rJkIUWbt+Jn1AJfdmR/O9iIh2yl11hH6GEtg+xpADE3eZY7ov
HifRn/m7oPSsFhTT0DMUb8B0D/dW6vYAL9w/7VVt5kG4KtX8IeK+mDGW/FZjhRw0
Y0Jima6mRebw9P2YC3ayhaOC90bkVNJeRwlxyDJ/8uSJS5G55NFo2KNRImIMfgQM
fomse/WVYNrt6LLlLa1xdm6CRiQywbCP6xBYhgTLtjcNBIQOocMMcyze4766U03e
g84wboGOZ8RSM9PdYFyoz/5XGq9VrfQKw400EzfzDkC4LDsM21rPJvoVQLrbqxoN
22/MXnD1PpvvBWJjPlfDbjFsTQOywhR3W9gS4BHJzAPQ2pyifRXVbG7FNlu5xBZk
PP/8h2n1XCbMV8pvrk/SDk6+evrx640EUsOhetRM+/nsyx9APryY7/JgPSyIDNxo
34UIjlsNJQImZZcHtKLi/WS+cHCHI6ipfcz2opOt9IrdaAc/EzuT2o4c71AkLcho
HGIPe8bpdwyK2hlfWbjePZN5ma9ZSb31jbuyXSLi3w33s5w6H8Q0mzHTp5z39j2q
vlqxzBY4j7o/B8o0GPHNFFfLoRMELO/u5lT/nTtNjm70hYUTRgVv6EpiOwPTZx9o
7Ft4TiaUBAKbPpVD9QAwz6as7jEwmEsDCsHLtoyQMI1vAbn9IeCKa4IROu0o+qL3
C2hXlYCJ9chcGeYPhv5fNz0PH5DfnLmtazvnQfpc+3wD3rgf8YxyiqRFfGH82kq5
8h+5g8MbNE9dUpPu4YOhM1Q543/RfsARsIQA/FCqM8hZTDe09OsJzHCIpuFLwR3J
7DzDnxsq8Or2FZFG8VkCtvffNDVVSIbRozAbPk2ZbwZB0NqIIyxlKph/MrBTORez
Z9gu3lIZPCLypu89Wy3lnyFWAsoJXdekDdM9uFDMFOfCTTGBxfKdfYjcRXGqSm4n
a4H0uor6LTEY8FULZ+WnxygtTac03OWT8azLFeJ+NO4SudXlYyOvODsAU9+yeCjX
YVlR8Mf4Xtg05rnzgfVJi1e6Oujsy/zVBGHQdxC/5m2a0mtPQZ9gPxW1+iAzouWI
6XKf2PSQoZCuo6WjYiDXaIwqUoVCOpgypzTLzBqledoxwq7fc8BzCyu73Mw75wQ2
+s/T7/7e+ChmHQeKiSbVPGU3K1y7YR/bIqa0z6yERsqB1mEDAJCMz5Pvuk9SV1Cc
d6mixzvib5rsEMHNLxmPwBPejH4ys/WARHkkdwJ4vG9j+0n5gh63tZWevWDSA/2g
Q+1A7afmS5mQTtptdx539QW76TUYv1k3lTQt/c49dCvvm6qNxZpEQsuO2EC8O3bz
njIiAgqL7ETFUZ/HkeCzJMNNGg28ebM9YURWuLN44rbFpsM01fjgxt7CD0eHIfI4
wkYzYvhDvgL8B/wUzQBFx91spqyKPb8I4Yic98aWqZnDjm+2AIJkx0LAvI12N1jD
gXKIPlzRIHbPam4Msb1zVNUfoKFPqeKNYXkLgqzNQriDtcM3KN9xKHZlYwwIc4cm
71mZBFA0UyzY4zJp1ijHdHQAH1tg3MMMRVcT3MXfi1dF4PAgAP7RffAnKpE+8+Se
hkqaXUDT4S7DrDVUseJQb80g3xZsKz5lLAGIaD9sJKJ9oJfCWjzhvKCSzfbiYbcX
lbwzrAoUj9+pe8NBnc19P+xOvd0ETPnsYzTJfI/xopUn9BQg+ulQw17oA075mZud
SFDDbH+ZVSbTR8cN/WbG+wCE/1+hyp4C6ElEz4S0mmZhEz8ypqDvL2EinPdzkGny
rCC1YtYsoE4+7DJoeRj1MY9JZ6TKExARRYiDxANzherHnLSUowUdw4U1n/Gxfon9
BZTylCHTLfPuufS+3dGkz7ltKKnV+JGwlwI7zrX6S7T5MqTXyqXOhAk2clhWaXAO
aaHh4hX7UBzUCtjv86jGBHJZgfbt48GREcESu0+RaRaPwic4HOH+gvLUzrNMy/Xw
IZj1PpNQLxibPGw/HyuUL4A34Nx1hzTThZ9oFeMTidTanlBg8imum3jFdk+zCpfk
DjYeajcRNMbg4aFuVYqMDjb2sk7nEzsoxV2FqDrIjB8M9aTEi/JSi//xsa/Vah0k
lYSUJjHJrKPhvnE+MnS0G2619vruuT4YRe7+QBNa4FHgIiZuIba8xlWbUeypP1/f
p2S1jciv8Owa8bCTDi0alCmZvyzKbGcXXRGeqQEm6PPO52ZMyuXsAsU0JfR1zdpX
b82eSYnJC4JjV/ZzdH4JRQ886J9H+K9qDae9Gt6677fg68jQC5LMG8SoN/ULQDz8
gyA5iIOizDhCKfih1NMq5sBTVMciV3KR/gbLaZgHwvImNu1rbbh9jdvOtTPdljnR
A24PhVoSr1JrH1Ixd4dk3uc1MS2QNacT6js7ddJeFbCMfCf71sm0rSL2HlmDmml0
6lABtvxtmQLfh83EJ+3nOPYKH8bcMc7FUErbUJP3AhIhdlyGPtH71nZj43tAZFag
N8Ghx6Uueno4bDsamCjAvMysbbcFXxLxK0S2VkmmmjDmmzFaVQ2+Ac0GhBeUL8On
hSEVBtss7wPMQuj0bbuja4HJ5T2pbZWlPIfl18uktUd8vt1bVYkO4WHk+LUkKfu6
xx0Ge1v4E8s20rmV7NDlaovDqNCaf71PtziUgNG6t1w8KrzUPIc/jWEekR/iMF3e
D68roqBGKrvVr3Vl8ux5VxcKfa4q09bOc4qgZOJDjPpJOu2F7YsFrqdS2pCK1ynp
xwFKPQ9V+F9Fz/orLzjDB8NZsTfoeP/D3O0/qsEyjWDbd3Z9I7KKWKt/Kw9AM7Qo
lYYabz0LyLBJmRFY/3/F9qkQWwQVqqPMmFAfvXvV5+hH/qBxRJa3BrAnx1tvPGNg
A2+fP/WrzP7Q0slpSOPkaeWbLPUDAVG1uEaNJ02nJDqorjXDneNG0HCqfOHK9JwF
8oird19QXkYtJFKPhgI5Bv6/cT67FdcjmWYaLeIRVdjmHCh6Hbq9s4ASp2yGkwNm
7DuCLbeQYJUd1MIr0PdBncb5C+6Evde/3ZJ4shZDpjLKPpU9TrBZh6PGF2niPlQQ
w4xbJ8OASEst6jocAp76Va/ZeE4y4RtTZG4cYDl1L720n5NiwH49VZsHUlP/07XI
0efRa5+5ojluAuOK8yxZJLFE/ZSNAaDRLdQU5N/Jy8E=
`protect END_PROTECTED
