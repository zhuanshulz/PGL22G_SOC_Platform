`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z/IqzshLfEKJMEH4reD+67b5KdiC6PQiDMHJGFRoF9gg0UvuIP95evjJQTIXpUnx
sgR0tyasvDDfbAalk7ahDfTDGtaDQQDh6zdI45CpgeSK+dx9naZwii5HuXsaqhBw
UoTmxYSOnJugO/sHc+WN6FnDgudWuxh1UCcIBH0PvY+I4cKyw9aiFYVHDW520Nrl
CyA3vrQ4nJuXHrXTza+Uk9a8V3H5YJQl8jdYe4Gww7mipjrAsCiwiw5oPPreHA8h
KmfAubUJDvDKAGsCpEkmH6ou5qAtZKwYy6UDrIl/7MXZgm/VuEmtJgAUY7E+khWp
hPnqsWou/6mIEo37PQrGSv7QJzQNem8PulKwYfxiZmBDzIBzrmj0RB9P3tZjYMQ1
/WAyjpYBS8cbMQsApGBmpEDWeGZYnRMtiJ27zCcKlD+0uqsHXDv4GWQIfazAM49v
JNyVWR3JWyavNyiYlFe1UEy51HSly5CTl7tKfwdMslP6MBrWdXn2XsF8haQsKy16
SeDq5vBdCGMaweKyqjLM6zNGEqOz5k+UKRU3jGTEsN6fcDFXjCjtkVxzKdsD0wXX
RMq7P9eJPbne3iORlnYKBMxy5qji14zHJlqw5wJytrOPLrqmubTzw4bBhBzxC2e2
QTAS5XiM8HVsqSfHLvzpRo4fqF5sThZyHTWcZvIIwNpJGt24KUYIPJd7cfNDFLOE
as183Ft4+6OUnUpmb6O1hKbRQVrLV0NqhXRquEvc4dWExp45oHD35uvI/7H7kxlK
fA5SbeqTAGkZSAKiSO++/NdWFhmRx8Bl/tS1WnM2nj+kuQIWQTGBc3CUTqVQKbc/
VrR9nwS4GuNQNi0Ci41cNd3FX59WmTlDVdhSft1z4Ue0nW/SlctfQOqbvwnwMwHE
5ODi5sZgK2LU0Jpe5DAb/YOW12gC9tFCxM7g3m0BatY15GC/xF64gAD17MpXZIKv
Y2TGzXnUcl3jVTatAyQvqbmhGGprXd95GIMyGU2E/la2o/ZReviMmlWXB3KJycRf
GnXZ5rE6y9Y732tfhk47QW9lRBUF5Z40qULvtjSupdmDPtRZjN0fCz16zmis+bN1
8PVmaOayj7c+jnHyyo7BfeR1mGEcl3Ne9tMR2N5c0Vpo2ZPYa4+j3BSIkJpz26YT
E7y+m2E5t1hwxIM0s4hkRhO9DuK7ah8pqDwo/XrGOzuxHW0zfKAMfBwY4OTJed9m
Lo7unMyEODVku4mDO3kJ8Sn/Yj42Oxvh4bC9RtHzH4EgtvHc290e1dW6jnzqMblb
u9TTTRAOCw8/So1d1m3lMDRMEqg1mhKitSydmNlhmldCSOmCeKM/prPj9piu4WGs
yyzwKZPzrnM4Rk78XFVCd42GeUlXGy59qnOgFS3b+RjfhLVcK/9LTPgFh0m6MRS+
kePT+sPSrJVu9Z0RjOi3+ZszCy62xQ6Ft1IiNUU5aN9Gu7kPRKQXxTyDKXezi8OQ
iPVSKguQZOdyPsl08ilFUvOQ+nzTBMt5AXhor5EDF/BxXVcPYN2fZujP0J+Tdssg
rrrMkIYYVtxN/S6WRnoBSbJtDNa6x+xfJQuEPMva+9+cb30JoeYd5pcL+r9nK9RX
C0ATNhuLWx7Ch2xKD772N1WvGyU6yjsjWyVbFMoogVbYgG3g14mizmKryya5auQr
rHa9WmYp8sVJY6EOR5iPInDvxSKfRlxU3y9FBgCGb74BTLhEKDn0IZRhBUamgRzg
JAO5QpX/5iC/12Ull6lXWWG9oK/4MIGx3dlV1II9buS9rBk6FpWu9fYn9mR5JQ9J
7tic/wTd7iovaYjIgDOag/u7YyKg2gjf/3cZv8l/9zd9k7DoyA/jSw17dQ8fBBbm
h3Kz1zHp0GMe26v3mGNV3ZrLGxd06hpZws2aRiqvGMtgTEX7YV+9DmXn8ivrk98t
hKhL5pLvQQiPFx2CjmVlae0+557A4/4D1f23McjpXBHlEwSjrWJh7lfKngQSZFv+
Kb/nmroflba1dWyGc9tZC8JbozZ6j0Uzi1jEpu4XrEmCpkPGQiBmZNlIxNC/j1uV
xZqSc8uBQwQe051guNVNMbxvYKchWmI7kY1nrvhzL/Ss20DxioCUo5hQ/GICtL9j
57NGUy1IgU0CPWrNVJ0D98WvzZx4ZJV+uzVNbbcQUdvH7ryVB+6bYEX+rIDDHSsZ
LWmXOCbSx6LnycbZHsQ/cgTBhFBJBcAfOP8uX+yvCTlWsokZ1s3S5jpBWSTk1og8
NYy4oQ7AIU8NSLaqgD/e9s1eGs/cwPSCWwSECfRp0WEb9XUqroLUavK4Y6IN/EkL
MtzaBnnO9VIffKA4pxkJUjDmvsEUWAoS15xRl0fNoi1HQFfoX3y1yx5Ermgv1zrg
w+zz/gWFid24BrZqsOt4n3HJd/aUkgmALkoYICqZNmDpMIyUn9CBLPkaXF4tq711
skfqtIZuYEOkbpsbuNyh8HdU8XMdohExJbWMH9/Z9Nfrnl9OKfTANv431kks2Nlr
+pihvrcrtM/BpKicNhRD1cf28VkyuY1TBh2otFYOBZt5atN9oCn5PGbmUMMJF0Bc
A30somnerRfOr5AxfQtdigXH3nHzzT/dWBojv4iSFHybTmkMTO1xgwxe6Iy1mTC2
jG8HifKdVJyV1qTB2i2iV7c9kIi8f3S/pnIjjQv2Bkag4iGQwYK0ZnXNqtShOpIG
n9DL4Pdmrono8w6KD8lZ3hSBgimegKceI+k5ULnv0rmNIUmRQ62YRiYHipUvOM41
XtZsBd5zA21LkNUgTjB1HmxVJsBVojQ07feH9dybLbZu2mkOfJLQI2GvZpcXIIgc
9ttPkBNz6q5kDyVj1yoK3Nx0zmtrlxn7/Xa3tREqCyy/03WNSI+mZ2dOsNjDiSiw
`protect END_PROTECTED
