`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NiJjLc+K5mipzcMOEpCGJII6Hcbe0eRUzjNZvSajYoqY5i6hHd7ULESwlaaHz7Mm
9EoP9He5p3XNQxTSB7x/SHzd2yM0yBsLuEaSE7dMREwuu0hGsRwW9Ia3hNHx8H8h
2RVJjIcLlm+SqUyOKf8bHiAKfegi4uu59GNfVamiz4yDHBSpInjwQtgScAvgqKax
vxusGx192o6upNtfD76tOoCTKDi1fse0B5RFWJdKNA0kwyAPD9pZ1+2fPW2PJwpx
ecNjxP28uHJAhWm5w9kGb/5UYeuRbz7Df1n70b7K+tOa+V3m8RSeBNsESgT4oDSG
GcC5QHor9DAsAIGIbkKXlNnuz9/0pAT0DymOK+hzLzkqYaQuuqBkFzz+bSJi4MQh
LYKF19viSOodhNFWOPOF0c9Sav8qBypqhTzCBzGzOorrRfCJFl3no+gAoApS8/aG
5iMlZGnedSwXV8TLEpsIu5bCxdQaM3mSrXciQ+FXFKBTvEBuv2nD3OTnFMUdFfl6
upIkBxNftS9PXyBr66+GMqPWApKileK085iTtsMj2lqdtx5jPOlFJkqNAKvNMWr3
fIZyIOLU3HOzYknvUs4Fq5d0JJ0f7+MqmT5JkXJ2iwltU8OH4yOeU/ozNc1cCPOw
1JNDZjX8lxKRFf0iVtmIu1hIkhiwYK2U8Ieu57xOd21WUaQkyOZfQNSbRF+Vr0Ue
vnFBCpL6icAwaW3k8ds5fb9b2EbHN8uBuo2bo3WGI77R6TMKK+I2Ea1OKWGvqbFK
LuzpVKUZ7PSTNpIhzUnRb7jaSXQyG6tYQoOt5opX19VpBH31NdXnnyMMkE+UxYXq
YYq/TtWoKLD9BrzEtjZ4YwyZg75O7hp7i9tt3V+Ti2J62gTYkq7N3k4oJdhzdpU5
UwTic2DVIT5OM5yQzOBa9VD5g54dnsg7zMQn8blHrR29G2j4JMacHN41KSOE0IkJ
S0DhNnsrA051hToBItNjAUfjPaf0xo3LTDJLQzqhbunyATsZlTaJRRksTuX8VcUN
XDftZ2WTL2PoaWY3JmEYCZqZhy9p9higMZXs4EdQ0vY+OIC4MN2OOiIcEgqhGl+0
ZN3iq6Q186iW1fc40HvEketQnGAAhTthBfL0uw79hM6hEzpQsc8+4JdGLorvh2u5
R8aNre45rdgHVKuX4fJuFkaPk4vv/pBZ/CNkZGSJS59FuPs4jsa8d6ozkTkKUWDF
UOI2Su+RrhM0A/+9rD3zN1/kpbMRkXr/8N8yFe7Kzu6Fub1cPS9r5sS58PAhMqx1
HYQCYUtOZePhEctnxJXe2w==
`protect END_PROTECTED
