`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VNVtXm5j+e6yrs7W0aNfqByQmBgpsrM5/d+TM2XihM48bu5r8lNwFcQL7LPBYB1R
vACTvDya+zDbKpxngX1mMXUEHt5boObvsOCCVQh7AZDeuLckFTd3q4WrDX/q5QHS
NanLz1YgeEpTGJ0ZicpbPvLf/MTw8+J5f+w/EfXh4Of6Xl7bKpYAUV3X6GX8QIe+
MbYKZ4vKpev1ibUlJ5oPldjQAXYbHqjOTiuto/S3yP36J7W0iPkqG8Z6Pdax8hCa
tu6jJzu9LX4EHrQa7kX4ghu0h97SA4QMuE3cY7gEnsbRE6sGvo8x70JLe0nxSSyu
od069Q5q1Kqnq+bqo1wKQ7G2Q1Sz5uHsV/9wzOCuWW5dEnKqZY0FxAkDQ0iinvom
/hbcIw4TvsE/Au4BeQ2qjFy025UTCsMHvC/4/PfmiMOVfCWN27cpkuZZaNDOWcbF
XFJjHAmMYzU2ajGsD7TMCAmedqX2f+HoO9QMyxEX25VE0GONYAe2RvzeY0WU51MG
peSpE6oULkOr4CXYJoTCsYaNe9/8y9In7iG9xllsuyEcHq5cHMm2PR2jwwxa0Gjh
V+FmSk7Ti2AaId0wRYdOzPiQTR+StH+uX2DBDDUTbk2Z5zuOmTg7kxg0cDKrafij
8XypAZtDpeAL0RuIHcEKcar+guEhMxgkFGmXZeICapCGWKJxZtkncW0ZA/3CQvb9
wybejUXR7yb0q5R3ov0mh46BZvpI7a2852EbIkzDQHQjNtzbizdi3t40g115b5T4
c11LpChPlHrossXe5tYQZNAnQ2Cfqsx2LLNDr5ICJrom2tCwHAnk9sPvP7/f5InE
EeD5xfUIzKXITu0l3QWfAMdHXnTzNiqd49v1v1NID4QjjPc3efAXOjUfWa/nYL/f
VXHl3AHcwscF98xbVFL6T0UYrENmF3biJu3Ex4BN4P8Vs8dah2do5J7CcvAk9lUj
ZSWk1niNTXjRfuisCVV5ZefkHRJnbHFaqWvc2Lh8Bx8NSfcnALq9/0axres004qn
z/bldf3Ku3DnIMcFJcBppCpeC1fnwqbm6tQop4OaT4gboOjgv/M/7af0h7e5AOsm
hV8DThkhcV1Qzz9vGBExHKPgofVZPT5nlAi7GtmWp9kCIoy2ymayFlDOQnltE8fZ
ORvIKji0m+qcbzEaT3Oa96xqP4O52fyLf7K/7BOsaVeLsfFjP1xuaMW4WG1lx2p1
Nm2edZQ6cHt2qIWQvNmmIGgZ/0a5AsXa5Avtn4e6+0NnlSRZAOjvUS8PBVYkeBrx
H3ton1l+1RonHEuh3hEAOOAOyuyQCfudABrAMCtKHMpqoGLeS3YKqA8WtIZFJNAk
Dj1ow2C66v+wxyUpo1Gu7OR6STJ0VgvfgGb7/gAVEjbJgeSQNEJMvWrFQXcuBY+L
Pm05LvjqQ5OhEPF7MjQCSFmVzBabEtSffclcZ2DH9zsazWBbMYfNOoQMwaYMgbGR
12l9bw9Jy2Xn9U3jODUSo+9RckugPJqbc9BtOVYBrZRJvR+9ed4PLEnvqshk0AXR
cTdwYBPYDCis1fiTqBgYzR0CcSNlMxvVpt/lpl9Ld+K4rnX2XJv4LJwqP11lKn/K
hbof4ZSbsDC+Il6fU6Lzfd3W6nGUzUFkEn00amMu+bKbC99RTVkIL7dSnACgqjZu
YAZnVtGPRmywQzPOEKr4xitLuaFn+iXi9y4Fmt2ORZC3RXmEi69h3G6pPlg6I8+4
Ff4qnUwgn/oGQy4QAbGxQbxN1WrjYFvXyj+FSdM1m8JEyNeWDt0VD6YlzfEHILCM
AkPteNmuY2pkOw86J+OtTvaUD2inkNlkCinB4lz9es3tSpA2QKFyVzZibo6B7MsY
W4EggWadIfo9nltrkh+hgR5l5yrkMDbNqkWfWuwuQv4zSiWqa57JfhmLP5Np4QU/
ziUkcA+mZeLdbcXTUm5F+AE7nTeGGc6e9P2IO0+tAi/Dh94leUsZzsXgm20Gkjni
XemqFRRD7LdQDShMqbAM4ep1bNMQMm02jl5c9PM+/zv/IYEOlmWvpCaUcUPR29nf
ghDbGr9wBeG4PKT/OWWLCvV4ZYKMDmFIxg2n4Ee6g5RAbh24hob08D9wHAtG+8yH
vq+PqwSUCBpVBLhxMiY64kzH+JmdXzGQR/vGXOTaESMhvpHMvBhL0zMrg6DS5r8j
qovcRWfW0p1T1g+cbWYJh678VNRyZ/woSPYUECu/YKU24V+2oBc8a94uBn6Ieijz
eu/Dg0W6Cjxz+jLFDYTr60wn8rLimZgwIdJtMpUW+7FO0sLtQbh8hvMIqnTUghMe
woUmOWgMPkbNsY8/+43Q0HIH3JT+ufNU03mRxuC7AgnBLzhZ5u0aVtdnaumPZ/+B
3MxtlbsxTkB4XnI91MYK7ae1JrvJWKw8JUyCdNLQmuYZGRaw/RCHz7qiidAkjqNR
S+e083Scmf4Uh5FzzmCCJK6GJsmbix7K2V34zEpsjzgXcyfxeJc6i8XzPj9l4X19
RcpAepVfrCcJdh0lUdAcLDoQcYVbVV34SKJMze4BY9l/pyQuc71kNrbcaizD7CLN
fW6DkXC4nGYswsG/UlILpEgl5WfiaR2ZFTe3D0pz3hbdI2JnjAH+GeEVdH7cItqu
NnnajCuq9sWYSa2YSOeX+wR5wyUZuqJQiZS36otfySnBOFhd0u6W2dmb8aCBzrDA
GpaeutVAxY1wjU0XP+/1Vo3QfL2/N/g4o64NqBhhL1jmNkDEMMuBA3iiSB5UAL+t
3UYRs9zMhoa62AfqA7x4OLQSUbqwXmPabWHAQU3wAu2xCMl9aW5555Lah9ZobxQZ
4kTxckxeh7J1/AxTjyT/sxTbNO+HDiz/zFJo/ol8N4OWPe23Vf1pfwwX9vT6RqRg
QCEfhYHJnTuJF82qB/sEJAJMg5xI4rNql5cSGRuTdz1EVzdTtQ3xwbWHkqn0WvJJ
BfLgn/DZ4hX7fOpE0Uy/Cr9RVwa7bfpOkWmkQpwflCgRqECuOp9dN70xOiTxvmUB
Gu7c5wpt/btHHRyVBlYmopxnVieW0U6sE28mLeiI0J08e9beETVQqXnaEq35qxlU
GuFoqTccVcLOvic0CMYzuJ18ZJsdoZlwIljxiYvs8w3UyKpui/gl/6y+JpZqNQFq
Y/U8bHXfnLOWhBJAj6iRoLI9XZhOy1C7aYk75h/L9S6QVBlaoVjHN1uGu0FHNKko
3X5+dxcdeRZ8Gor9kq/ES2GRgl3boLx8zvD/l3/oGmg70OeuVft2JipXoD27af+G
oBQG48BKZvLpADxReEuKiFxRyp+DtfuOsuRleOZiNfwnHRGa+rSJoOuKtWKRQLjV
NrTy+V4ikojmuEPw62fh57R8lbizHR9/I66fOfw9kSIKNoJhgNwPWK9efqfvRMUH
oCTB4X066mPDa2GNxbnBUH+EAyO2aGamFbWSNypAmPjXbCJsYAQFpsYSE6I4Z0L4
Br4YedzuaakLTwgwD1dg1K2Povdah2rJlYAgW3DP/y0LBzfGG42xc8ViGBx30fSa
cMM6Dla+fOCJpRZjCdc0QOlI+1rtRi+zEWs1ZxsNP8byVsZ5sARWJhQPoyAYToOW
q+KxT4B2MqJ102UoAN8aGnBd4l6GgrIlUoWY23Myb+Y2pcqqwfp14NPOX9PO69na
mBJEl5NjjH6BjQPyPhxR+mShDeSwC3YY3dIp/E3R7xaD8570DaZijxNA4O/3AeTZ
cmyjaloIkSwnvCuOzUS2ONQ00P9vgGs2CXxtB3BuLSe89SM7J7Bb0L3CH4Xq4zId
zdB63Y9EKHhAdbRNHBKknH4ZL8dyU4Vblc1fIDet5cZ/u+WOWIaFAW65wqOsWfGf
1rgpSz+nWU49yIjOVMMQEJsUxXR+JbBiFZMS5iS+VlY136D+QqV9BmyRZINOTGpN
BtU514Hv8Ud2WvF0GXuNdG+Kw8V2VXojbcI3g+MsgnGxmjEo1ZeFx8AN1DPgdWit
DODn3OVPbv02HkWffcC4pAFKXtY/1AUUVcc17WBLhOuwd8QRnbbTSwkTsZ/dl4WU
Wvffykz08zzj69G3WddcFwrZwP1EyV6X/g3dPdI/OXQe2WoTkox0Xb1olKK/rmUz
82kqtc83Pd2DhvwS5xSE4hPz25KrwXXV4Hi/0ZURGyXN+Fc2BrShSRoD+b88JHxP
+KSdZWVzcYtzOD2RNnpWFDGLVbZZRrsxwe9tFdtx5VMy2eGd1ODHhbHGSO8K38Ax
dXTSYnJxsTNpu/77D3chPowHgnhZMylNsd5NWakTDmAhOReRUizr13Wbheb2iNfU
9Ev6j/cG1r90s1hcXj/ZNb0LkYRxew5nnXPTaqT2GrxYEHL3KWd4IeLYdXg5nkFT
QCRRnSQPHL52TNFSgEUXdfMgl+9OpR80TTOTgc8P92rVKJGsGhEgebOQZb8sXjED
v0QqW/T8gIJveQ6XnHl0Kk6q6PksVayuxGb/18HICNGoJrKI9ZcEBrvRrnSVc6If
WNZYDPMJRZrjBCJuJr3U9FOcOinbeY7M6WSzfHR8R6Dep0BvqZnl/9llBYliIwaQ
+KAy1Xz+9ogxii23vyevkCUMG9hXl3WnAmq+ICEeIPZsaF5TPsTHgOx27qttbW41
SXe/C+dM5RgCrawTOhy40qBUI8yYkW49JMtiFH+fqkacF6a8XsU/ENPo8WMCfuwl
/U1iuDq2qG+9q+D1rHbkj70kBH5FJhLvIrBVpBoYWv1rSvwB4ybahrua0vWo4sgX
rs/00XOgLNd+w93dohprLh7yVVmBfiMoq+470GClXIEAfDaFx8CENks/cVBQ5QtE
3YPvID4WzKBB8QaRSU1NQeMpGWtUG3xeGuFy4LfC0iN0FHQ10hhFkukuBdP77CNw
/lTIJw0QpYcXuB1eyB6JeeZjdAlV03zUrrfoEwM7Z6XnVg5/oh7OJvmWd/7OwUl3
KzWAG34GaI7/HGopKCZCOUxrpvx4Tu7gaH7oPqoL7vhfBgDNlIcCWXknzkRCBInq
3g5gz7ONSk6XZUCCfggDgVH29ZUxojDA87jqpGXRTE724cB7t1lmLb9vnwGdHwep
ESyc5Qbfat20DVgBda8svRrlxkoB/gbTaWCOEAvxvenkWUyszOeqi37bmUcbDqqt
PsTr5BlEkfI5P+Ntrmn7uBBD29IPlF5lXBAyXa2fMhiomeheRa8b6s54NGxw2LSg
cPSGGT4mhpCSD2KQswy8S7nMmIYTh14qgPmH5d6WaVm9caPh6zXkvQTIBHSbSX1W
7yzKHEOD7rpKwNRMM+vWgP6gMmQft1MHhim2BKVrNKHw0uylRFo6uBpY3pg+azAK
AQNVxc34GK2epauS+pv0A/YT+sgLj3ufoJ/ucrQPSITguqG09/pnmAgS+HyFC6xA
sDjF/P+rKf0x59wPwlrnwMSTZocUugO4TxraTqabnym++pQ3scr7QufUWSE5AUgv
ZkZjtWsoiz8CJo+7RhM2SttSa+vjxZETC25zZMmHRLLSyXVU/193okqJKkdHZtmZ
Tdih0nZt7PcrQoUWgT7hd9rIml1ZQRfldhXRdqwALlrKsgiIZyK7W35WNaIIF2ac
QLuKIad/MVPDOFM7ZBUvB//2RapmLsJq420crDZSzgEq3ofvXktpHewxuqXRMhru
FxZBgGtBf3twNQqHIkjNexMJSv7TcSIuL2bIQmIUJGDqhUxe7AkZmEaxB3TrsoOw
+mBp79lfQZHD3/o1wg5yxQvcUIh1pjikbsyAzH1Ywhhp6o66dSdcqJCpPHq+ztiD
XMlZV3um/wZYuQNyg/Zmh4DgSZRaoXgODasNfDjO6IDZik4T7LHeVq4I1m5PjnSB
dphS/o13hYHbzTTqLjKc4ZLuMcspWzAZTN1NXnum/n0NN1Di2FP1F8mmpXNaTW8E
9bbVcq4K6W3x2kozMyQr0wmwxxqXohymNXsH8m0/xpoMEwkAUZc2yRtBVZF+kb2v
AgvnXxKeGs2nFmjkSnFKnzMw+6pp/wbH6mGl55Y2jfvF/tSwMPKrNng9yJxnUvU/
608FjIkLRDn4UZ7sU0Vu57Ui62R34O7LyUuJVpFEaoSuZJ2f4lODYqT07zLHd4US
9QMn/VC358fSgCiM+Z2hCHqNOw5CIjxOY96o3fMOVIqvoagk2KMIZ//GloGQCsRE
VcFbmqKm1k4utgK9lTR/gQJQcO5dnFO3nXNqE6/VenFzfRAZAjOMKNIOHP7GuxZi
0naQLqy1FB3JZ74/OyXaDc0BKw/QNJ9Wz0TGiaCVeuEhttoH3Nhv0vYqBpbNPhNX
FD2/dDh/Kdrkumq2xdFoOSlTHR84vTxYSIaKBfQWiFxSPFF5AVuwwBtxVp7GTojl
LFEe4Rij0dImHB2n1G4HlzxJoHVKN7JTvD3zxMeh/NyHSRLXYVtyyAhBY8guh90e
vsLQvkfVD5vjMo9BkEluXz4nfopEIULKHRtN1PI8EVX88nnLavcyZMZtaPIhjZJE
l2PrMZg9rq2prEL492/FOMBjOzSoeaBYBLYwLo/z+l6g9FiEu9MjoC4FnvoEXPwc
qcckuOfJVVeCcY8fuNJOU66kMDO+hI4uwfM5e9FrAK5dCh0hcQOd1zyd5bku5ZLi
amkARV7hX2dVwmHPx7OeoRiu00KN0CfJpo0B3WjqLfW89PkRKOORego4MOsYAZCG
w+NMeKPDg6uaYWpkPn7HAaTn9uTj0CttL/d8BpIT5RanyTzsoyAOwWl54Y4hJanY
FTdd4dyGRxEwr9JtnXUFQZrJC3CdoWFepGgTSKZc4lwmES6gAjJpOAoW1oS+zbx7
mr8NTZpkco9fhpWX61ZtQGHYEYB7XUBmrAByzfIE/j/ZIBAZ1UTjdqSfNm7kdOPy
DHH+mqpuNPs/tradjlCQcetGm2yQtCjKWIgX+5Ogslz+BkIzQ1J26Fgx8qeoZC9M
xuXA0DAewKjf+z2Wa0b7KkC2N6YXA0S1psQahXRShodeJzsgknED2hJl7wBKspu2
eL63zOv06tWrIuoiY8fFVCDc0iMO0lbOE8YKaCPwU/VkaB0YpUCOLFTl7OyQdv3j
YZVSm4eywfVzkaODY82GIdJ3xvDZmm7c6/hnpuOs8khrviFsk/BNSsj90IZkpgF5
kNFwOwcXQ6APTTJ/+fJ+zWK3i1HlNzuaoNVIRo9K/058kST+7DaD7GmswyW0Hf2L
X6pKbUScpl+/RhbTHeGTRmYsubpCiXdmnQdMuirxGx6xdi8Fnmt6pgw3E5pyHdaW
spNZn3qO5u6Rq9ToU7wL+Lv2Lg9jo2by7ZyOdm6Dkxt7gA5Gq0hpP90CIMkQL7TQ
2Pb2/Q63D+X0lFrb/pur1hgqr+JyiM7mrnkAW0meCgzDEJMv2/JVF55kC/3/ljCw
NyGvF6qn8suwYvU0sweF0kO08/v1nUjOTJXBH0tYTyexD0bSQivwUCErGjBnsCQ/
azz1mBEFNZLc4wORS33DQm1RcIhyCgMV5hNFIb0yk70eK/eQyj6BAnr3MRcAW/Af
BBeyNDzm605UYxsjJ5UgDxjqJ4SProiPmhb4IVnp0ekmQYLdye1aur0LxiSiZNpJ
0hSBMKEbPGb/pC2D/UmuXkLLrjNqbIzAqQrFrq1zIQ5uhO9f5pwAiZZT+QurfdGI
+tAMpRxvLkP8tow++WDhoYBCzpB8RnuZKuGO4a3nH9r59JSyi2isUZyvXxDyaBlO
CJUtGJYn8sRGAdCNtH2iZ1IHnUP/wrX+ANQl+b/4SyDNAZhbQmywUmafXKqNsOkG
E5gjj/usX03cjd+t/VvIZWAxWHQoJjc298S3rN+xw6TlktjzZO596jItZg8wypom
X1oFQQ2sjkWe386pZU7jjOQy2EnP/wDp1VakAxZ/nPsHrmdp8911te78drZFzCOh
kuczlSh0PTUVALMLxQvlOPXGeBdAmoRsad8j0ToXJKhxNrxayFcQOni/9ztA1HTi
jw2TNsNOED0zsAHnhy2uRy5CpAJDq6tn0zNoswrp9ludZQAJKxu3+9MevBZcg4BY
R7Zp2C7nBh9LblDaguXz/XFil/mXNEqpsOQzt4icvWQPZqyBknp8uUZkxmxlWiMH
kQHh5VL0o7fmOqkuiZzdfm1wh1xJjDnvz4bdjLJWPLj55e+ggzUGfuvyVlI9mYlL
1gWUs3DHtvKm0m9Ts2Z9Ym24yBYF3oIKKVqNv+k9nqk7TxxbZekZYOdC53/9szjJ
WGRyiSclPa2eNxsA83JXYK1D2D044KdKnSGyehsWpJ8FUlkZSVs9pcAEEC7wRZDD
W4F/PX6qRuOSH72rQysksBws8G+1/R/2572JdCGnEIAUNKvHsuNlmAObVQ/1k6KR
0nATnAnxlF2owwjvWCnAT6vP0+2GqyT0xF//ut9YePj7ey1XkRNWFDr3yG+M+1f9
HQdGJjW58WWcSuWFEzqpKTtS1OMMmEKgkJ62vOAMCDMHRKy6H9JsnQWFXktmmEEs
r9XMk8bbnXEqL3jxmGmRNvTVwNfMx6Tq3H+pCeKUSgsq8To3+hyAv3CdFcnh/R1f
LR9Ez8Gc9dRrkyHHMB98SggVGEmZSmNuJfEjT4LM05UfMuJ0yTm0oTu1RtbvuC8h
IcS9tEEbqDEyplnsgTGOZYGkedljI4zNJsyBhNhBz1lojl+jo4AYFfA32eNJUfrw
FaHNxI331CrSdB71GTyXkKkDKDEcd0cxyYXHQM0WBGeVjAijKZdd1OPu1EvL94+I
sW0PZzvHCRchuONZHDMI8+53UOe782o7JZPFdB7ju6jeCfBEZw4tg3wDpO65EuYD
26qUfvFLL/jv4sqOgFmfrn8iVCl4Bvqvl/GgK8IFjuySQZ/fRFhj2rxI9Ba8DhiY
ig9Bu/J4BhSwAyn4uxABrQClpa3OjhVWtcj+INTGf3HNAJs5GnFDKRHWhsCdj4J1
RgVMQfgNcrccI2ZWGGhoX0r15KIi/q3N4xUlJqBz0DacGkRkpQWFbqZMb/DEvTUg
zZAsCuzFV9RFMAPDmPB+ck+6Q8L/zhPDdAy//xiMp6cxA/syPOlA/PIGjThn8fDl
X8j5AqpqcQsON6h1WA5tKGMmlMTRs61VaT5uw6zDK4UBSjSIvScV3sWwjOvxNy/G
ficU3CJdnZwL4kAhJ/oIcpxnzBAeejwQO+Z9hEEJZygPx38Y6N2j6yAYXzoTWA3B
sNEnoznF27/zsdr/g3BVGB2qiiWzdFHJACNPYH/rBEGwg6nAXdcPjxbwD12I5k9j
dH1bPx+oTRtA0coGbUpO++fb+jAdv8G5XQAzOoP44q5E0azWC/eh9Ykp+wNBoTSn
U8lwSSWASwCCv0C0YenAw3/aL8OSY/xlO7P7RMW1kEAHi1QnP0i0I9x1UVGtYLf3
qx67Za7Xyx/SjX+rll5erXMAc1HEzURjH28Tw6U3E9MS1Yjcd3hPDDn6e6pvrehk
5FngpARdH66/2csIKl+CWVE/g8ohMtjDxYLeDXQNkDrRICgLW/A2wQTUKW0UnXXT
ayWJjKU044ugb5MvgnmfLcOjSMj9tsHa4CX1lrAlpJUzgWnru+XuuRaLh5aASSNb
V2tLerK4YLzprcJaEWxPqhlp3tIvsdKNz5YuDZTcnYjpzN3PyxZyICjLj6OMH56I
OQ6iC260QHwM3Xo3bXOphd6IFmFTZR2fN76+Sjumu7VNlgRLOYHvY2TsqnuHIb0F
hJYzkzXzx/LN+xL0IVzzPOKIFGOjgfhmmg60g30YhE6p5OBeO37udJVQerwYZF2b
v7BghqQbzE/0ImyNS+S/Afq5DvpraEwYeB+fLzZ6/jzQimD5p0nqIM/3xSGaWcWt
vjn2/gtBCk7nkhb4ydJugQ+iAm/+NTrpjO1ihIwB1TZovLjE7G9OokqfO55DvX0Y
Rbdl7Uw9bJdT0cj6eikja7cEor8EwBsis3qgp1tY+KxfTR7dvQ+gfTNfWevbiHU2
pB7GtmDGiC4VQWBXmwhmWfttExpetWpNQg+0biKOIostGZsJKGZZgBJI7cqV77dv
qccLaGoZJ1DpR2NZoy5lfWgMl1cN1If5bDl/nqMeXooodJ227pCHyT183HoC8bBV
7dcTJsbStNlD//u7weyvqYuy+dv7ZvyH9ohCbjKUwqFq6TfrmM3Xy3rnpnfhdDCA
4oEktZF7A2ypyNwy2XYh6qpLeQy1ebJMTg3VsAVzjK+qiAWLcsA2732YjCoE3/at
vWTRiZweIQ9oNfAdaPHv9aeQsdRv5h6yQRu1qGl8vcI11p5oMbJ8U1WSQQLfrCog
Sq3flIjd6R/KDM+DPhKCFw3ZAd7bEdR/XcR4Qn3J97BKTUQAx4dx4HwkVsHsgjUB
wBU6NXATlcELjblFg05JTSJzORppPFOapmPgoUtOELg6A2vQJNzwGYJyv6WV1yH/
saCC1m0S1a47QzhylgfaiyRqjW813qS5kBEDZ9QEG14Us3DXMlPgi0x6mzT7CwNA
EUq4OPy1hLvnJqNYu74grE0H8HXbH0ecr6d9l88ql+qhGLv3wrVvPL9RjoDmtVov
YzlWjfnAnccAZzJ+zsB1ZocKOu+RDQdqjzON+vh6RdMKynLCSGgOh+ouQkUV4rSF
B43tHMWk46suSaIpeJJQwzSJEpvzYsgHAMmO7pFsgabhMvrzEOdQwoSjQdFlS+5t
1/uJa0WHyHFTlz+1PyxRAZUooBZ26p89tcqDU8nb93gy9j8pPe00gLE+GdQnIeT/
XXUS4YAmqKQ/xHbu+Ca7q59ncE8u49kmP18ImTRz1NZdSvi5Jh7KDj9OwJvPdmhr
gNnw4+qWVTIe1OxZoWj2hDe6xPHP/kO5VMMAN6lyGBJa3UBeRIU2ptAjSK+hRzLx
byWbpS+S5o49yLTtMKaSqXiyXdsVbw05WNJghO/IFMeAAtmrilZUKpDyMRDmTEep
5PWrPfWNWE7HRgNoAdbrIWmSmg4MO28IFNPDcyik3eTqBlXcV/ehjyq8gbgPn/bR
32yUFkEgEP/ZHZ0UhdpulPoSDjKyPXa0XZLsJf2QqYLHDz3uGg7VBgY3a6KbiGcb
++Zl3SBMJobvB6AmDAjwKEwGkCrRq4apcQheOnTyuGsDcrq/56npfu9Wlw3aLJJR
yXtpAJEuekfR9fxOMr39FUfgzuUy7rLljk1WnLLPONipE8/COXM7p/LLVsV6xriK
EY6aESnp1UaY+KoSCaBsgCIhFs6GXE4VWxT29HwKdbOI0Rik4tfA4Qr7mxihBxG0
ND+io9P1kHoDrTPbGxIV2QKNK3lSb8lvbDw1xbknVkrqZmbL3GhqLnBrNsNFiBSO
zLMtlp3yOJuyXXvtsupyn7xqsrt0btfBVrQFyuPiuzeKp4H+1YOQgKgu/SbYg+8S
19TMWYl+PYPHgeZuF0CY+ZfJLd8YqA+Tcp/KMBldwNMKRxtdWUjTj83qSU+ue3p/
GaIW0NDF0rbY2amxnHwyxkDtJj2fVOmR3gsa8W4qwNkSxCyX1VpOug/wJxdSymHI
vefuldT/7gv12q4/75v3DMzoun9JyzZO5JWr5UvkqB6G9KPN3EwEI1kwppD4j6w6
BsuKwHpxyGBeUkLUPhNv7irnsbuX4UjTLUxXrAQUNIj1eEwQopomYf/juLAS/Wro
v80l/2RrE6AMwaCZ8syGuEnl8iqejh3Lzx9UjBmjxTvps5xV+yR51m25z5uvxH22
SfpR2qKnq5oT8b/9YgZr1tCCiC7GcMcm5BIvADqtUv0QGJfe+RM2K5neuYHpcNbV
3rpJpvleNVYz9zzChpabKq83eHXK4lfDN/mw39wbxga1ySLMhyBUsk1YdsKQUCnd
jjqClyHCWto41+NgnlOXHPqg5yWd5kO8skctg1kRj5d+RhQC3nAcLTt6JYDem7oT
Lik5tngpV3xjN82KXRE+x2Euu3pOFy9B0pKuptUf67khX8Pt8TYTNuZur7k76Fmk
GFID9eRKSBcTD8R2YfiRyCLMcUWNkvDeluYZi1uwcy8YzZz8U9K1ssFgewavdNjc
hg+TFgbM0CYNkadHsFqZzGvU2irJdfYzVHCH0SEOYlB1RedQGD1AGa7TWH3hpZys
7Vg6qhHdog49VRVONhuSPSpGjeIOzh0EyI8nuRnY22fckXCh7zeYdNH5FNj5QE3y
MDGHwaWdjhWoRI/v9fr5k+3+WoGs1BCkELd11b/q6N47FF8NMpWG7psdwMSvprEQ
km7+lljPyfMG1wqU2/M/oi+o0fsC+Jjl31SlMVn04Bn8jyAjpm3DLaqkI3s1cIA/
f/VIGpJA5Alkeq8OCkw1lOYJmUCGRB2A8v3mBFuTHkCv06FhRtT/ywfrCzXhj1+4
+qfImFzWH4GQ6YJN7UjguBCmYrGcqR0XliVeYXDp2lPDR7NPx3dgxoGivnXkF04Q
wL44Va+xv3wp7GnIc8dqONz3R4M3SrjgwmtyiD2w5l1VhWolvUsi7XqQZvOJvZ0t
Z4vizNZL9ZsNbAacey63yCkSfCk44Rj/VchzrTf4H3omKriqD+tTo1lZmL5ATzXn
Xqg3dqAg5/o0zf0BXxy5qHjmMmSmBk/Zy0n2sCqgFFWt6eFfMADfKKEY33gi6/t0
V9K7sk35A0yLmf83Ao5UyQmu34IGJTVlSHvjMYkq08P7RpG2HlEi9tUAUIHu9Y+y
NU2EC7044o9ye9DhOuGp8JiC2JH9dJzVAvGeevaaww7NwPa3/uLFB+b5MbYkwkIb
OeuQHDX25ym1WCFSpxjN84c8gumnOj6Eo1sNuz/S/SQ+B474g5dP5Bo1W5M8e8JF
2wjGM5wsmAsIdcvUkFUgkYZcgGr9cRbXBmGMRJiq67mYEEgeUd3UhynEKm5NB4tT
oZJzF4ulpmR4PXuoMGP4nxq4YqaDSdWqjUzC6aIJZDdOw0mL4lFadDES2WFwvImC
imJ6ipboPzvLoiyRoxtcQ7uGQzlw+BQQm1u5xXqhhwc4VVF55nqaCMXuDbPny9dk
Cbq3QYRpucTmtQ8NIb7U6wEApnfQoM8tkR+AWpmJoTFdCu+MMT78P32B9xd9f1T1
zzOKLGaKqKYK9RW8nNPvmMrxPZ7Nu3OU3SbUvuBb8WPGVQ283aqsCdIMAdwWRKi7
OMEbacPPoNjU/0aArUPlK0YJUmseFSL5ZULTImjOsVdUuUuRDC780aYFkuIqj81x
B5QDbmFD3ZZ1VirMvyut6TX+OvSG0BTGKUEBp0iVGLsrO66+p/g1NRXVu87qPdHX
9kaF/I83+gAkR0vwc2WMdX8MDn7JfYu40Hnq/5WAPrvYKgd6jqwcQrDZLMRCR6gA
R+EFGk5ZsoroedNL3FE15AV83BPqt5wjoJdcEUcG2eo/SE8NYu/p+hcbh9ToUccG
0TG1ivCo+85S+Tw1QmEPUnxsfAgVVjXEgtjfaaN2qNVnN+3LlMOUv49vMG9vFUuw
268OMKnGL06ZCMCtNMNx2CNqPSH4e0N5TBN2sqQYzLtGhr8U2YLFbKEwqlHy4Hmu
fssTnls0rA96nTlPzFvrKLPmR7e3sJ7xuG05bPFd2lpcyOHB2OXs7JfxynMjNdPH
sh7QkOi/eppM3CL+o7i6OBH8T4e0n+0fyVI6CDLxFHPaKGA24DlZe6t7jaa0lwQI
KMt/sjs9r0Xb8sVNrt7GSHe9fa4wEfaIsuSsWLOtHyQV1uU9AmHrfCHzB3/V+XWT
FJuFBZN9JKjHIqhDlBHT5UZC0mZglRUxr5jWKczYNd7WJKwfI2E1owzl34x8JwHO
DoNoIPIMRG3MA3Q5fH9SdO1QFYXzPDVkphl+0PA2BWw+DCwiErPx9gQLdD5+X+wV
atXBDfvuw+pkw0njqLDzDtlbDwakTdJO4IV4M+Vzkh6C6mdEW9+hZYnYz7hGnk9d
okSgAcXkUGQXMOvnTFNoQBJlXcMTitsJ2hWqEi/rNHyLfi141irQjgg8BTt9ljzd
3T4St1uTkEYE1cHOTMmGWv7Vv+MTT28eyrr9fXd10M4VS5prXrCi0038cvCh8FGD
J4Nk+RU/PWwT7nCcYf/+lIfsoaL/nPyRUZwfzLx/Qxd+OxuL8A48/f/uOoz2vgcw
pmQHBPSxxgsZot/ROtkaqlAN2kVaM+tDM2A3WCGAIvuGUToOKN1dHwLQH2J6R6cj
+qgTDKOKcjksbP1v3bF3P2oYHCZQH6uFWSgDoNBy/HensqBOEfhnNqJAvuBlyY4b
MFpEtp763JSkxbYddhIaXWiB6jlodXaMj+W7VY6AEJR196MWQMxQKch8DOJK90mU
qVXyhNrN2uKRiFjsQN25NQnkG+uiaB3kT0g0Csu1YCpLXxJeg/88u5RSUz2Jwjc0
uj/QJo8neABv6Qy4FXzF8gmNntlDkyHeRphhHvBmw/eD57GIpUXUjupvMwlEV5Ty
Wwl6EEl+RxkOOv5FBbfHvGFzOdlj8k2aC6CNkHgSFpgy0dXXaI4B42Q1oEaGZbbU
kJ3CiipFkMh1Pt23PJyvJnJJIZ0XQFggnuwdmMTUsjxox/83gxpM4lpw77XjjP2g
6lqumfgHGJCGAAmt0G343zHh60ijT5gAsBZGo5292UvjacaCHKfjurjUei/L0wBX
Qzwzvatz3hq1+32QWrQDKbneXa4z/MRgu2CkIgVz291gqjzB4nJtzyxU7DOzMusH
+mWyT9X9Hy8/wpeUiAV52D2AdO0aVvjrHv9l7VJx0EUtSMvyDi6gnCWDV26GyBxH
WijgUHoihHChm5WlO32XqLkQdST7m+5F5bNKCzpHOLguHqD4PW3xu8xicOBzzFBH
o+JaKGdfXbwxNc03rGpXO6kwGe+sfVJPYnFCukzdMtx1NgIxNmuTHQUdydUiH6Fn
SrcLjWlaNFg5GglG6uHpkq+fen743bfYp2f4GoLcGuruwRUKQ9AEHSRO/Rhe6W3X
PXMsiHpTEXw5wX8qRUjdwbti+yvC2zJWDNZRTn8+uxFNEogr7eNac34pUmdKtUqZ
4G8thLU/DG6stUQ2F4xd2DY0oSnq8gS9g/de50WbdfaYc82m8pSsS+rbhuJdg4wX
IoOcia+lROkK7u9Q0XJlgOjfbBbbitBhRSCe46CLDObmypDwW75X1ZGG3Qb46/hp
+cyulbmIDRssiFceUdnMqqQpnkeC9r5K0fDZxxDkNvJXn715XVGFdVlhAzP+Sz2w
5WhlO3RzlQl5KQ2bN6Vj/m2P1IS3v6RNKGyI4JDYz14BImVk44hO7plr0MuEHtUO
YH3jsI50D3bB9PS61k07vMf3E2J7tmBbwJpboSzUOE3wwekXjVBHH29r16NPzjLX
ER/ze3V4fpRxORpWa/X2QWwHdB3V/pdHgy/wvujqxogk0FGaQyybN34zPeNJEGYt
dhAnbVvJHF3OJj9z6jBwXpnawRjk7vNmMY48ouJq1gYOwhF6aPYRUgpvAUg37Kab
c2Lbr/kIuudEqbE+k6wyVjmWyvsD0CqiyWmhjT8IRM8P8+1fRPoBw2xEJE0LHjrR
LqL7MWhXgZlVVXomdD38WerYdeEOooJ5eBylHeAvejkPqdLzzqCMaSefMRMYXlix
Z6TdWUp5H/nnICBKsKGW1zWiZG+7A6IkbCbNB3WxlMfsj5ou22PPxyvR5ftWoqZL
oDy2bzK51rYUfcrFfrIwRZw8UxCEdpvIy5BpprpqlRSlekE33397NNnq8VogXejc
kUzL5QEAfs2bGB2OgLe2SCzw/dv6PN7y3j8pWQNaDTfsrS1kC+RTME16qeTZGEKZ
cn24K3b6Amz9DATSE+kCY7r+3YzOE4q7MpXUuhLJ4sjcXvf14u1mvGcsaA7Cbcfi
UvJAl97o2Nt1aez9V5KdT+AVFYyivc7GY8KKSE/67E2uIJBR3oVpXpju5U/0aLrL
q7gZ0gJUCcSgZYDTx5yURjqkakY5IPeV/HmvVnGe+UcpoIT2GDrcbZm3S4kVAlmK
jbPNaGIP5+lCwfkYGQgh5FE18O3X6WKcJ2w/OBD/tPT46ByfpQkkd+b/RHsBDBEK
JBh6obUz8FQjpK9BwkUI//9AVWw/SS9+2TOzW1Pb6PHjXVuExwZ1b7AkWMiqdYKC
b7TXdVLLagLvc8RD8JVSVQFABMTIdHg6i4kWGop+pRiSjGxGWjmkuG4KT1BI4O2Z
eMHli4h3vfTQE3PVFkPh03Um3J+6eICTkjXJYfqD+gOLBiNMHImt85c6nWS7ie/A
3/GAiddYIQE7cyOzDRjhfT2hhbvC0od7kPRugOv42Wn7Oh2Y7MYBeHgZhA0IQTpH
y5Hr/CIpulJXfK0VQUNfeoKso1xuVI3LapJ/uQMuZB5vWFFrEL38haGS7iBQeEHB
KOc5VRuu4xFhT5RKeT3oK6pvAadDoELP2PQDQa65EYEQ+SLstj5j3tBnkzNjZg5x
T9B3+WFntf6JjACVlXwerIbELfUnun61g8Pi1kvCHrecErqlTSj6yVLYy4dauyhv
MU9Ri26ljTfijtmoVWP02PodRg/vBauWZQ/b6DeivsIu4NSPK36r2K44Y2H7fLNi
snwt4bc1jm+85mSe86lK+amrtHRwbKb64i55peSBn9Q+z2yssNRkp70ZS/bGfhL0
b21+R+EhtSPlgrdIRYnTgc7dJRpGwN/N7K/ScMGhz/3Ythq3yF7I4rYWXwFGsyHS
qWJ0Ck/4VuwxMgjZgWHfijxUmBqchcaGD1eKa7ad8z8lZadd5QvufFjyjEVnibCf
0FdsagLBadTb3A5nRdoOVy2PySvBoWfz7I+D8naO99Q/ulTm0O0Ku2UCVxdlcfGM
T6fPXlsixyebiC9SYrdCYBBfTe9RaeeqqB+3RFvwBiUoGtomY681h9s79xluMPIX
vuW3QtRz9vGLtIBrWo4k1jfI8sUB7G1xEvVNz+/8SiaOBlkxAhtR96e1pUOWcB0n
Dqrn3adfSMQEksNk2E5Y7S39HK2yyb+jDRgy1ejYNLHacLaeCm8nK58966TV1QDT
TOlH4MFufyLvYMpIbp9tGwwYrA6fwE98cubNZ6RSpOwAWRMAXgdC7YYopmp5Upp+
1fi66wlNFHbjXsIjBlp2UvMkLsae/x5wLEN035ePYT0L3iQ1KG3x3OaYwMrLrJm0
8mTQxoRiuHfZqSyBunM1VoZLpwQxIOc0Xh/RV2D400XiAZkyf8a32xUq9C8rVdu3
9BhiaEg6OFdjiKHpWmzNQ8Y7O1Va1tKFV9G/VgtUeCTcOhKh++b813OP7vW04Kqx
2d1JlwnFWHPEBejffRVa3y20tOQD33idEV9a7kBndt4/XH67V3IXdnPB4+KbaFQ3
ICDf8pL3gIEmQjZjmripgQY6aByFEeS0Dj5NdiQPxSHcYaMnPKQeg5F9oX5am/ql
r5XJCHTo1+wr40OLLKyEEsXQUltnPQpJJvcrlD/BTGbK5o6M5HLQ86r3JFobmsR3
FphpvW4yb2VIU4OmXgXgLlnjYJDm+VEZW5bwJN9ZKM9tGgaZ/kx5nk9xmEMIwCmC
vXivCY7OYID69CQko6igp9VEaA/9pTp2DcURrsIu77xT9yXbKrOBdXCOZqdjWzbc
trS2z+aKMWFpG9CNHIEEiGvbkcGDodztemOKxR6NqEU/LCjPyF0MC129Oc6IPZV0
7Euv+E9CfGdVr0j5i49bGW6JU9dhSmcE8QpR6vkKlSuPYGU45HOiVMt08Am72Q/r
bNn4ZL0dtWOszTLQIfAeDbl5UZex3fHFmt02FYThaIVtWL2d3xMJQTBt3o8y+y9u
Arvz6gua2daqbT6wafRpTPYeazdeE91/TCRPDRAQ99LSaKQhC2VXar61cbRvtpg8
j0o/zLCYUaYjfV2odzufbzGjeLfbUnksQuKnXaRaufy3CYuVCeIXd55NIsnjKntZ
LNFnMoBff+MWIJMZXx1yHUp5aicS+iGS6BZvZD6kDSOmqfj/UzhkG0GqkSID6HRU
qThi0KZGYjw6DAha1gF8cAlTZAr94713qXx+dYQcMWD31XqBX10Zp0F1VLem7N+O
JbpQvXxOXqik3QAYeA9or7fc+VrzZTEdBUUnHUV7xg5dfO9fJLV4gmvrAM8NU2mK
mDZHT8lNzlnawzft2mbMVq7jR6aiMBU2mmatmoolKmhUeDZ6norWpREYXkkXVunQ
ng2GM5B0q/ZWfh36XHZVT0/18ZeuWXKjPcaRri4S20uC/KqiEn+wPcR/h2lNhyWh
mVMYPoUX0OgDblDbT2rQE/4xP81icutiyXZp66tdZyTg5h3vG0tVg1Et13znnIaB
ESifsss/PM3KmoTW/ZnWhqaN9VmDB9rrmCDyISn9GO7hLEUxBV7WfdwrbNTEK+qO
yllb6/bm5NnW0XAvjeeLXLZbZ7xJaDcMpPS0Eh7CFs6rFKQqHB1oIQxqO66DVrXE
ynEDjp3j8Al+ABNZhgoAeL1y/zvP1ru+gJaBtHgZFLkmwT2+JyEoBz2rJ+F+fUP3
bWUYq2d22f5gXk3tS3Q+4VlYLLp39h+sEc6ZkDtRQMsWc++RSUeRvJrXGm1BiAGh
QeAEZqSR2ecsc9PDFA2wwj3HTOJ/YVwV3GNxhifSUClY1o3FS3Rjr+dC13l59x9G
QcP0YwwhNX7ppsyC28ChGZARZ6+mEodJHWRJGV2Pfrc08nFBQW+0OqxeLcni2yhm
YICkgFW7CNHIx3wxzhqEJsYdMpVady3gvxWY27jWIzH/tb+558Yg+4fXr4UPPVde
3ggZNlq1R+BsMQZ8FSuyOjOdo0qF59DmI3u2G+0z55xlzN1wjg4elwMiH4BV+dz7
JrLnc5yDeR4UN4dX0kvha9hI00Uc9+QXlY7Ad5X10vMxHbxmC0VWA6D12XEcrxyb
tarnhV1EkNm1RYNthhXbfY/dr6fj5KF/KGlY2jcAU44iHvJq9fNvSS7lXdO41AYP
IDMadMXn696b02hZMYGTpx1R82Y6Yv5CMfEtKJgAEOt5AuhWtLCEegSJ/psUDwsH
a6TOSGVP2PKWmZ/zt+FB4Gp1H5yDiwLcqbtPo0iM4F0PAgMRVrpReB6kyxfGMyLa
ymmbj4LVOG6FIbAUpvWejJXeWZH/FvJn3aNMvxnS0oY1ZKUiGdPprFzPfuubyWpB
HccxkLWY7L3lPWZbe3fh9MvTTj+5Se0TrwKodNCHkhnkIB1TC/S9wwkeLgLEhpLW
bZOrodTzvo2/N08yhcsvlYB2mrrg7pyJn9UOx0Mcz5yoFkHK6KNo+L+gTZeL8B3/
AY83rIP7k5RVSfkfv3hihOQj3vxIQmeVgnGLxtGe3vdLO11VY8Z8WrsNETgWGLxL
w2oGXznHyraO86ndUwXoE3cKL/9/1YwIz8IN8dWmheq7UtqVDxkwyoS/y/VMtFup
BBamG9GBN07/bFXWlLtbtH7creM8O2XCL0jezbRcxf5AAsLQ2TaXh8gz51MET6p/
cnUmXA2wbpK+D4wKuw8QVqEKaATw1FevVzJRy5UXdvLpA/j9Np/ZW1fUi3ZJOoLJ
1OY9zleevrOZnGX385nx8w46Y+30ue3AKqa7jXa43mrU8oCsJrqI1di1NL25V+bQ
cOFdnKhYZqErpOZMaRmcHVf0eZ+pYF4RhlfZzLX+pRYNLPx2JXC3EKKyT0FNyybS
9qjWGhV/ag2MfcynogWHXf7+jV+epfrLrRdWgRBheUcevmEI4Y3Znpl0QeLO7Bdx
hWaZae+ws+RajeHi1i9VDhUG4gYakd3ATJknCm2alidj/pKzubozUfQbaSvoX44m
L2Du0auRGcnisW4FPgAXFeooYQ8NxOXLzK+K+Ah8S0PW1mxuulEibn9MDYvzfXWp
1tCtAJj9LcKOI3dZZ3rvpME24oFqVduMI/eZLyH+ZtFRfAMeg/zhn5fciPUqBgsj
a3ZFRpPyWhcqkSHVq0ZtjADlC8x+p2129cfM24ML5xPe/sMb2qgmL2pJElKQ6F1m
qsPvubIkZwUbgCcJ/CVIaPzD+d9xlllG8PtSk1OAm90fXuXfucEIngfCPuuknzK7
6cuqFsv0C7WsEwcFN83UWZu1Xi82pd6+CzTt37l6xXCtmXgR2iv+3zQXLndtUFUx
3xn43ORRmTAGadZZQCcixh0SR8gTs2SBglfQnbxVm4KxLi4irTh/XhTCd2vZiFMs
U4s7lv5Bxk0Lo71ar/MFC+ky/txC17tqk9TXSUYeqNOrpzhIIO2OC/NB2W6PMmKP
NEvY9ODw+RyvchlFSjbiVz7Nmma/PhUJKROxJYWYakPF0OAwl7Raik7IKebmUml1
U304J0CMKXRnw5oHaxHksVZHFJfO+lXM9+XaUzLpAyHgU6c/LV+nkxk51pnwPaS5
Ta4es7HIbR27wofk+/kISZyqhXfp/OBzraA0JjmD6LCVYCoejuwynA26+KA2+hea
Pr9Gnzevpq3uAPnvSoHd5/4da/y0NvuEcBWjFbtvbHAT+wyu5qudrllNPWQVP2a8
OJcHBBO7hbFX2q4Z/jvQvkLDf6qMOo3X9qh7R25eAfqbUZi6gsWW1TSe+ZbsCboB
Rpk/Mj8iegR8uUP9X4asvECH94v+CUDCb/gmgmb5nCL7jOffNggPDyMGfNvRGA4p
S4I9S390gdxB9vB+9ZdY8zICOZ4NM6cCj+lJxxlOUf4thUEYSzcYPWHAjyCfAngh
GUjdGT2Claq+aESlt+0q76qhSa7txaiAwdKEYBo+LcvFgOg4uf3VxO4VwmPra7b2
KdWkaLLonYXRs6otyQf68xNL+t10rHWAvVXIWxsQ0ECtKfnQsXhBbX2cMLsGswWi
1a2ueub4BBxeAqQaxOsajOdW1CQj4uWoAD3JMpBOpFBoSQ98k2mPJP0fqDw9ZyYS
yuY5zbI5Mi913ZIpCP41hxvV/Byi4PK8qOmA2JcyXfFafmss2YjYS95eVzdG4pcA
HI8J+qCw1kRlw/H9FjUHK9L84qr7ahkS32VCgJi2HClQlp2tvoAMrcXvAjs8YXSk
Mu8a5Xdx/ecYZ0CFtqNWXA1/xZAqtnysecigUAkc6zroS0bgKSWLrndfIzsNWV2S
J639sALIx2FAmdwZfQjjMYjUg9jVMiXsRUfg4fnjoIEYAvokMPNO3YaUKRToiXvm
ctROVTWtcu7A6LjIHueV0hPv/+Lm9UFIStZ9ytZ7p42+hPpcQZxLk47m09prgN2w
D38bmb5Jf8ctceiMNxB7JMmmMkbcSeMds+vQiSmSQlIPF2uqCG3jjVRt4D6SY1hF
1HzZxVCu6uIiuufX+w/f/eOBAqvbO/gerpPT6YuDOE3PVBP/+1EUJHgurVljE41j
cH7+0jTxhCRIksNt9wlyYcgfQhjmLRxE5EjAqHKo8MeeYFAoLasPRqo3z3dAvJnY
giFISVkH7sGTu8xmP7Q2Tlv5nxTcOx2eAS7UEA5eqF9ca5L8Kfw5zwrO3J+A99MN
382VsPs8zwuQM0YxrGvJpkc7IZJgY2lsxBnNoEfh4WS4fFTVAOxB/k9faeGSpXeT
0ekCsf5mV3xOUd7/HEL78PK8A5jEeJOvAnABdYT68fE8Eku464IWb1zqxA+IPgQ7
KWpEMB2JnzscdSjVc6hrBLcNFXApajLNKr9FjPL1pNkb+3Jtfv5mpfHjU9jocxYC
RPnqTYrCdrleUuqVUf0GNEpkx3KyOCOkPrSwCtj43W++oNYndkXIiAe29tSow1rg
BfJAUbJIhFaxpKXGZSY+Dogh7nQANlwrCtb+me66VFUli1Yyd4iZEtV/ehrM8Osk
yRg0zYMf6ewQoKiXslSnqTGdlrqaadzDc2NBt9texnbNlN3fSM7B1tDvHdIQDPKZ
toWO3wkSeeCL4S8Rjg6vdvVLzGz63p38LOzPe2cGFlTaLWkTiLYNquxQDFJMQ6Zh
TQQMEV6vlP9+lxHBSXDNnwNW6zT567Dd19R4wngKvKJCUvE5/ziDMNZ2n/g/Bja9
HUYorrQDLmO01ob0ss5qZy0C1MlYkQORmbGX2dUj5By2GLrWdWSFej59ZPARqV/K
1C5p7s5DhcVDsO3VTVIK2LF/zTd7wZZCxPQ4Ys4PrGTfvn3PFl1cR8Hz56Toyx5q
+GTbfb+3tSs2QMO3Xnv+x0SGVtqI2D1caY62oU+Gs/h+tM/fgaGcJx5LUYXYnTEK
hYx+UPpaROQR9M8qcXm2mM13USa324soLAbfN17sO9cyY+NLhIVAgjvoZ3JXgk9E
gU8j0jXvjwtmgFwQuWc0ICPIiegKmrxTwV/8A0RpI5jd77KQrvxh/BJBkkl0ojGK
JeK7txva3FBNR1Z99IJ0roc9XghVZGCMnArt8Y+VpMzIfemA7KbYla35jaHuwo8a
YeuPtc+4cRlA0Yui33iLPi/UgpmKUM4ANjcWVGRJ+pnBW4uVmlP4IqqbvA1sZCU7
rk614cu9yXPUTjnOEaeSymcCmG2XFjQ9C5zUdH0EP+GCk4UxktpQ4gZhCpN3fGkQ
/1l6tkvmV0wLF2r3mN+BoendGKmLxXJ4IjH5ML8RSyL+48t67g14pYSxDTpd1nfo
UfNvZHO5E/n8iy79hf+AnAAuTTRmN/8TxrIIzcyL2ZsvL0w324ZyZl+rvZFZoQrD
Ifl++94jNvIaavAcFxVnfdOx5gXxHylFzZdYULWvzXqHP5w8eActjsrqnj1TgUlE
Moed/nhe6qOenLfgDwAq836VGRyQNYE7l3eBYHsHTUC94mMog00qmneX36lh2bD5
Z31Yn2Mmx4y4xCjByUJEXKTKaFFvvra4ExcTHknc03uRO8xzH47oSF18Btu938xS
AmTHzEIDxFjDdm88TghPI5G72B6SP8X0Zz1FiLcA3LcejkX9lCX6ceAV/6cmYtZK
8u8PCpcV0PlRiXOHKdgEcn5J4kgSKgT0lLhHYDXvYoQPHhViHHDc4NBB4SRrLlpk
k9T2QeJkkkEBgrpTuvcUHemAOrGig3yJbJATRrLPLXbRgs2kcmqXQXNQvgMuJayn
agHIsPo2bsZn+coj3+svbull0DGiTqZXOFnlXkQ7nbwTZL02OWzr5QNZfyxceamy
FXaWim0BuN2NW0k8e9pPiYXtjYLIMX4iXDI0wayKK+1DC0xGR3V4US1hWs8590SY
q/G82XyoRDn7YDjVrOA6KN+fr/u++1VhLSl/8Ynn4bjwxcxJT8WkLxAtrNtdJI+Y
a4S2aMJ8/NhZfMPJWRxbAntbk5SADebygDHcpj2+bmH1uSfvUFGY0b2aBEaQ5aYg
GM9nWvj48UIZShkBX52HizSw7SBdhHtgYbMHA7XZ011DOt6F42iKzPWqE7feKK2+
+g6xji3MuFOHPSQVJi4yaPCPH6bXCyxsK7Ponvk1t5eCjO0i1w6AfiRD0aKdh0BD
dq1/+SBaTk/Y+Gf959genSjI95VRjjimYeVnoAzzbCf7Qw9JyiOiqua8/mxvhJI5
lj31qg1vXkDZP8vCZFcEcwIZ0dYohHtTkOM/0o3NvDYcP1UUIYbIy5oD8D5rvxGM
erLf5zZ5/FFjOaE3CrpjwFCgKkY3eyvz0Qo2nOwdQ4NCN0XiIIdVa1wofcOlrxMr
S45Mh290e3JSxiAP4kyR7e7aI+dAj24yq4Slo4okzGff9pFVGxvfSIK9jw37r+bb
Shw63wguPLMibISHuIRbou2rpadHr8c9ykPoHc8Iki9YK2wBq8Nh8OkuXcwkD0l4
H0J2/nE154qa91/83xdC1FC5MT0VPYYpT7Zta/9YUOZCHtNZ4LmRGjTEy6IRd6so
zXTOhZTuW+ied2YnG2yABRw/NFHVdc1aWC19t25K4JB9QMKd3bkX8X2GUxRPkA8A
ZL5n5/GJO/ePZLM54Ajy5eRBqeAsFzSzh4BC+EpqwO/VVye8FgOt5l1Mgo11TEM8
2pPQm4Q7wny2NNVBNjx70J0Q1+Zm0721Cw4YwmeFyo2nhKKl1VL+n3cDQYN35MSt
O45blcVT887EFJ20IpxbYqQdWGh8KbRZWlqatDSj6N52q91sQehYD1S/tifTZVvT
3yYosmFKa/MQQC/4LenTDHsXCfifUeNunWCVFy+Wr+7ppnm8K3UenjYirgRYb+ar
nj7a21qQtPLvoSKNZbb1TrrhafQ6LHoelO7SdgIp4SbApCn9qMNRkPKq8vKqOAfj
X7JvXsN4A9WlKS0JzTFa57mNnC3xudESGy/FjqPOh0xBqbT9H0lU004IFmvLCAem
4RwtfgBARB4a6J7iIs41jlmQL0YaSQStNQ5A0GY5M6Dw+9nxF0QBi2xyxgjFKIaH
SM8osDgZBgJtmKrvAKuOOUOv1bHoHYVNd1NleocU/AzweFAAFfH6spsJRCAroQLM
aedtm7TlSKlbsgg8tY0/oTYHp3pBb8VAYqepamPq1PNWhv+Ruqf3nHy3cZm13Xl1
KRxwV/OMsG/Wg3cZD+KnuSVZXvaR7vP0xcdHSOP0mCttsBMTsW1nQKlAmcZjAKzW
TWTEVaZU/7xAQix2RBWiTEITu3sjits9+HfoKm0nYt5ii9o8JkicvoA5/mzXxeJw
y5HiSrctOR11ZDPN+uuqHwWcuq6KgTjT4+5N8RMM44AodO+90rYCt2sGMUvmM8Ch
aHxFvaA0vDYyhOWXdD5ydGXuK8AZgikKhJCZCHkHHcpOXgB+cojCqrCRVah/xoA0
YLPGrGs5O9RC2lbQu9tjt3sUpaXglhbtKW8WWWcrj4aaGZ6MgV0dMFV3f92BQTpc
99QmoYkvVfFeIshYCVxnlPrX3FiFTJLCfu70THblWQXj/IAOtmjGteAeIkMTvG8k
jCNl/7zj9FA2+B1otKfsz6B/A/1MW+fTcsvsQjIfS1ALChL48rv6xG46072koVl/
pVlcqBCIQ8/KlQAWEHAg8g0LwG2S7uSpQiNGdRy6AykKSYY441y67epxoFy//YAr
F9xgeIpNFb1yK6sziVI8Nt5vdr+a7s90LSmNy545KX56v0QeM95e7n7/XRZcgbYN
vLsqS72AapCt7TxBwx322V4cndbYGDTQUVa2N6EE+9HG7VTsfEP8k0+ygMZER/vx
x3MW4zaKZ8DToxp8ueh//ugHRgwiJP3Gg5goUrO46Xt+T9Lit5jxvUOmOsSIsF8n
ZFYiMgLp7UEQrcFR4QykjptCmy2XzKJ22U6EADuCAnsS2gJwyzuEPFhFjwQKM6mY
4/OSgb+m5zoF1vKjfCf2y/HUWJDVZjQ0cOBacGy5mvZUd2iHmKA4ZoeQ4F8Bb5vV
w0fXYCcvJshQ+YVAwNB0OFAFr0OKCqfiNhO5ApOG4HHfchCy33UGBtpQsovavXRK
VjZo0bH8KM6JqayUtBHiRCPaI5olrwtz3QK2qhAs9VeoM5e/NqGaCdHFZEA/c8XE
5citLzmr4BUGG+1RZ7KXGQ8toK4L0P1PbI7oQT/mHV4onJoqCPLFNvHZIFZ0eAtw
/Yl5soi9TCpnZSpgk2v0U5jaMyrqR4neYIgu08LNnflRpus0Uy2o19sOtFTPMtXW
dxldA6gj0RjVfoIlOnA2tluVLPFc57giT9SkPh0fpp9WTm+pFdlq6FL5kbl9qSlV
UHipXZHjCe5bojYwwBByib+f+xMOuzUMf1STsbgY5dgmB1ICidMOnMsjWB8Vb8ir
U/jjbR6kkhFA0YvA+gUjxs1zrNMDLzQAttkkNGlr6AZNesqa0d1/lzPWNNEAv+lq
+d3fvW0reFxI7cyTdpKfC9JGEvFwKhm9ivDjHreAKPb+ZZF5YFJ+KFkITNMfHRad
8e1wt7D4+QQRyjYBXk7TSWMdMtlIrlj14E9g7LcmgBlfJ9kiNgPo/MsqZnCGY5nJ
G/4R04I6rF2Bv6pzBUEHBsprpNPQRhirD8X7Ltue/g+ccKf0cHclpuSd1wzPVfkR
EHsJxFOxNxRBFCoFMG8m1flnrkyA0+G6gMSssz260FA1q48nMLt0hnIGbkaMSw0H
MQl0ezCh8Edgd2rAhLiMYKGXfDNUgHZlI4tH3xs7koUy0WE+gD1R1xhWxDojnhn4
lD+AlHWUFDxA5Su9JeupZgUo2MCTV3rVHZQNP/dPrOYBg04B3oId8ZdTAo+oxyTJ
TipwzKRgcvuggN4XyJQIGPzq3lgkPjPO/TApGM6QMQV8pCUlgsCqbmp3FFw22gkP
no/kO2UaYYS4jXnkM9BM07iB/+n8XqFkF9wluqFbwrg7Oo+ijoDGjy1nT8tP/0df
lxuKUo6t8U8he3bfGgSuk2hC+/0/Axr5JbmgUqFKMWU0x3uf8EwBI1AgKDjbeI8p
IEV8goD66K9nSnR4e6Kp1pR3cOcTMg3T4szCtWM/053eVlYtSM9S+IGij0U0f9G9
sR8mRcXtksceg8yhbK2Q4LF/diSq5u8sMZfsOKjUyvMgGaaLppmqQynY6Vc8BCpf
J+7u6EwnM8+WZomMnt0M/hwLYfS21m5++2zz5p5nbuWOqRSx/aY6ZSOONi5JwbN7
JJSw2TDTV7/1d7TXpRjyI/tyI+VAk9u3Ajm4ki2MwRTTzGCeFfiu/TAl1CLGlsnk
6dC9sG6YFXFfZM/mu3tqWpkLAb+uBhboaHC35WKAGOnZzWz65sNOqUgJOoVh3r8i
qUenCHfwTRVms1UVJY4/O/IN0EA1+oIb7N60bSi6Tmzq6qHgt5C2Kmwr4+vQeSAD
vViDjaTktW6o2jE39AlNMKc0jHD7EcjbVbF3Vmvn7rUqqE1pt1fEFt+b0WFiMzZD
oogjKVAPN4/MDvmyQikB4gaeHzjs28hu6keV6W6ZtfISre5rlGEDk4Nu/esgWetX
3bTf2OxRDEhIzzTTT8fzdiBRONwwiFwgQneMZqylx9Dxc2X1StbAnfmFN4qt+JvY
i9BAbX2tszTG+wjUc1bEeyoklIrQNnARVFHhA4X1GJ66nECWCJZSfhYYMHerA5So
Tjlh88YGWWqcmf1XD2YflXIo73/svryltlTZWVkwmdvmUjwIPh5pcu7RhkRpzQuN
m/IxMVRc+wLZWR47ZH//N2B36a42f+PkPpuMQGdSkXMY2lbx6LiNYnoQWHLrDPC/
7YOn8nrjelYN6XA7C2d1IDuPxiGvMUqZsNiGnbAZNrW3YO/oHdjnUD9QzYboJMAV
Me31duvdOmGSP4P0IgSqGMVbccKZ0LPM/uj9WizIZeEVgQAAqbA0/qiIgvHsr1ms
ShXxSI/v8xHvAP6/8OXh/RmFGw5A+76GOZF11xOQgJk3shb4Wb7quLkN6X4/vELx
gZzlaul1bUCWSienHt711QspqPwNqoYzG8GjM1Vh/rh6P4R1MImdaHBM5UgJiQqH
wPU6vUWLP+6PJPQEILEwtb6Nf3O8oTowst3CWz3ICSr6/ehLy5Yu9Dpc+wfwahA6
L8p/34aUyBuab8QcPc37R4aOTHqX0VQn0pVOdr9d9/B1jIyPLTBwaitAChZ5CMSE
rihTHcpnHra8fPDpaaK1KLM17jV+xsjlCNFa+XKY9xJo2xXMHO6l3V4N2yUm3GNd
V6Y1dE4TS8VyEgrnoh03SARrDugkXL2rUgBOysVL+9M75FRlpxvZp/1PVim0ib2q
oJuWoutKYQuHPS2sEH9GYmtjlqUEQkHChtmol84O4uNgOHpBAdiz+tUx8JCA9SMc
dAMUXb9XVjm59PxqtuTIdVt2kYTnZ5/X9JRO+K4H0aN26GbTq1h7HXd0dKsvihaE
YdGKl6YKiSYK8HRfdltXwsmIKtcX7PM0FM+keFzI5IAI+WNO9k7aA/2i6GrzWuUV
tv0SsWo/HbsN1aw4MmhExAGEQ+hJruGcFeVah2zq+R3ECv2CCN/vL5pBwB+alicj
x70DL/laSqjVSPrSz0fHfS+7c5M9TUDriZWDv/BoPmMOl7vnXHq4gL1MnpQoxX5G
fCdtH6rSLJhmV7qe7War5p/x802t8qm71EaWNQlQr4qP8bJc+mlXLgVjJvH2vQhW
QJRl0pAEeahr7sJ+R3Y3woEtyZn6vbTVAOUQxd7LxfY7ahaYo3LAj+ShYeQ4j2zt
MQUPnVXMdAcwEYS2TyxgufrtS/VTe6MASSIJsSHQMMnpb1pQnFXQ03UH73NNe2lI
/AggSjT8C1Fur+DrGBrUsckCXfK1hzyMkV9d7Hl+8Ym+bMW+c7/PrhH8Yhoefc4x
7I9QqnNVW7chiu4MVeuKBaodT9TD/UEOUOELC4hFXU/3UFIUnEedccw47LMcxvy3
4fthhtbpTxFKaiN/OvpKRVVQ/CdbHvx6f0g3AgIx9SsXctekPobRoZTH3VNbJNOG
vuAgs5qFoxNmK2WxEOIXNMsURObuLoQ8vJb7x7tj28XzOexapHvwV5PH9A/LQ21Q
l92OKf2UuLSSn+TMGdWTHoAVGobXAtTN/q293WiQRd+PV61IPyeGLSYA15/rQvV4
j1kSIRWk4m+cKRqd69FFmo2HaClqd669oWueaakWxeRaD7gedN0Rqp9TTvNS2vmq
Y0bSel3lQHtH63c6fIW4VDM/0vurIztTXzyPwgW5gBZnhdeOpI1z2APxhGVMA2US
XuG9OzR0KKg1fUv2LldClF3rzcMdGBrfReyn7mye+1/2EGL8VwNr1hseHLHBVLtp
uOtyuFaN87Y9iuIJLqu6Yk4sO8b3+flFWY9B9O+NCchtpC8WnNbbydqpsxZhZ/qY
GM0hfc89zIU9bzFPzIt6Q6ukeqXBgzFksAoxZE3n2nKYcEmS3czdV4zrx0vFSiTw
RHEPepH++YVwcbV2I0aX7ZF9EZ/gWfL3ITXRZIWV1jQo/AZ26gIhBFzc9ryLQTWR
x4u0OCSaB9qR66jEPFJ6WgvYvoB5zSufChTdXPDGU3uP94DwYexK9bwckvBgygFp
QRa4rLOK0yc2Aa1tz81b06n5XP/5C/kW7KaL77yxc/s7JB2ck9Y77JcSplMLt/tt
7Txwc3AKGfKTEC1PbBtdlG8r17DGdjDjqwi3plXQzXcH56ake+XTK2JO+/qGfeGj
92yPc+sS4Qbksrl7TWCe2XLqhCq/atrWzZdE4V52z5Bg+tYZsy+/fdC/Kd9bUmSz
bNZxB0gqAOAWk+dZlnoAzZFUZJJPddsnjB0/I2n5okVsWeVgJYajOfcJjKJ1lJSH
P7d6Qlxh900IJMvLYph2MDMO90tYlOpqslDc/sVHI1YudgLXMSCHZuSmp0mz1P8w
f1c/VgzHJqUB1iPaNQD9/VTa19WsgTLOXA3g3SP8VX8ssrnlfCAr+VemKLRVLFPw
czbaC8RZGgVWlS1D3UlgIFcqTWao9e3mzR9qElSxKHWzVs5scQNGx8k2Cyg628Qq
3Hc5CJEt/LNv0skUe5+StBNVw41jGxzeB8nxwtvRZLyqVEFEXhOOpQlIafGSHWIG
l9Irf2xJslnRrSD6KZIkoCFEkTnr4rPN2kLwrj37iofnVtbuzHUgoNBPw15vYb9z
ZOv4fIpWtNVBUcinUhxxXBCGppnzUKiOv+7dJaJ9n/Zr+Q3T4f8so1Sjbftri2ej
JprNNwxtRhoxpeIdqfpe98fTvQY99XftabzxTAGuPhAdtsnMMSM7LgYh9ThWJ6B4
WN/miF5vQUngui4oj3Z2RaeHiE3k831tnymW32ETFl4PVHDeCiotqhMkFUH+R0O0
1mnQnTiO5W4jmTQyd5ImqJr8bQJVolxewo6yIgrsFr1OKW5mnU0BSlxi7iJ04PTE
nwE+0SIiX+cmnVbNRU5dHMX7hEVhdlLstmL6Kzh/wpVZDQ4ZnRf5nb2x3SUARjWi
LumIBh7IbwmXabmMk/6QYxtaOSCEoWiTCUr2azw0NdSgPaBfTrPc2ZqlkZP4bx39
8VCpcdHpUIgtF54UT8ZZ1rfWR/6149xmryrA+zTe4iLGNnVrWz3LAxhM7neeI5Bi
RQezj5Km/7hbTyE3tYtB+mjeIn5SlGwd2Gb9pFDkh6443ffCwtTMklDu7YWEl/tN
9ev/Rsz66dVHPP47j3GIOpof+HImRNVChxoCOVSTzyHamdRpNEZtrtdpPD3fviKF
0JrDee7DCgmVjUxM5slP6A+MeZVON12GwOet4y8Vk3WqXbhNfH3rX8K2NIlpZn8S
wtJa2RAzIhUgjl8FA8SKFPn3HGDebObmDqEEoFEIY6FRGE5QMnpLJuS8c9sIADMe
yJIhRoz5zCwVg+lP8ZjJtZ9v1zHxr4LzCJvfoARI+2m6jtf2s2rzYOBmrL6aZFar
fqzeLn9eoxfuyfHPP30uSPtD+a7bcel20JOdh9/p22nPtfxYhEOTvLfNRCYpt1K6
nZE0rBUHrjB55xtIs86+ByCmIjUcGLxQxGVM80Ic9mcC5VVMFoIBfcbxcv8i2EIs
MexM+oiJXuEg7NFNIAPdLXiwH5FBpjPJ4c3tg5iXvgNyLrRuu/vU4/xlLsbk96En
7y6ZCHHAD/yfN1DKQbi+lMv/Op4utvTgYLvBABEnpfkB2py3Dwx+CirrGkGZKPw2
waoN9cKU0C1K58x7eQ5/Clwqc2JBEwrGuW3Y4MRI8GUaGE/D5Y9cjbd2MpWDjRwx
vRpXMOlZoP/4Lt9AiThBkFrXMZoeVj3Nplg1nMcPhZFm4mN4KXNwtLiQ5XdtVwht
7Fn+dxDgnbDszg+fqO9dJob2iVRUyhJjXTyB7P7Ol9+MKIAS2wg3bw7BWwAmZQkE
Xopbu65fAmYqgY3xwH/a8wDXtwFofRfLxsk2lBFkWqhz4jclxdJYa4ci2loC7Cht
MoVsZX8pnqJ2/W5EfaezzO5dexxaSAAcKNGLeofYMYM1vBqd33GKdnGn1hJvvBF7
6VRCtuT1lVoCjFwkwzn/bMDQ3F1phCydWEsFJZ9eIyhkIvHkqHWIScTXfP9gd8Nn
ZIv9T9neiMNeyiX5FGPZ2e9lyv+L9EFDRu7aNkULaBAJ57t7FyfWw760Dr1ZbziU
518pFzqLnbKk/dlQ8EZ9oCexAgAutHDfdFsh/PTy3JEKHjJwz065tsk/3g0DeG1y
D6QUQFX0rwnLQlTwGVM0rmyQ5eQny07Wss1Bihl+QL0GJIZxOEaQU8a1RxVcTd1Z
mwuO238chdpafVdFsE4UTeE+EeITwDpR3Xa1fremMTupRYlCzB7Yy5LDEXDsFr2c
rTOznRRbORBkBQgN8tdGmektJjTXczCVEEAYko4racvKNdOtULJFc0/HIlNFaT7z
Z/ULoKHCP6FnIiT1mq6fVxOTRS+5ZXdGo2fwl2S9/00XPc5l/wXiVk76hgxK8khc
DoVNkyDrhtJEBxIqVa+UYW1eHl9D7H9A9CU3wPiGt4CKEIeGkRdkHRs+gLWRfS32
mHIAbr3y/kwb4RpeJM2m5a5ocSbqR/hdwNIvaJ7WHVvl/bfWXHyKBhmvMYEe4qFu
ldNZziHZBS/Q/TsRadgGIto2nomaqRjvUsfteXyJBOApcK1xtyx8dKWtYylCYLqR
T1J8OgSoBP9+7w6un0d2Cy0D1zVKPUCMZ7gUM6Y5uiB3O3f83lgZgO47OlHMQhjV
Hlae7F/0K7u8zMjv12/RBQe3VdcGKL9U8PrM8Ee0MCEJdgMDHFC4UCkZsqlNE7DO
+ToNEz8Jy/f2i6dScLA0BW4dRsXDg4P3XtPAi9kPgubwLAH0Ld0HDWQBCGpm8V0u
D5BPVTA0FVJN3y7k3fISLl439MavggumW/Hj9PxZzNMmwf2aicqmbD50X8hln+Gf
FsKNxGykWCSgFf3xGcMJVefchBhboYtRWp+ujUfuY1fX3cfMQ74/TviBvhPWpqQM
LXWS1fNPqJjtNYDpS7Gyhdk2nMc+YuVwW3qamz91rwT2bvIpZIK6PquxoZewGJre
JD/l0KqjwBuDFQVE/b2leHU8U5/F2rXbex7MSEhm6hM5gLMqpusWQhhBpajEIn2V
2IBDyEH9Forw0BtQM1J4uQfefFd/hd+CSLT4Vj+YmnLqI7jMtbtGgzxr1aZipHqY
ckmeA1dKvwgm3U2CkOJ71+zZdF8RbMsn63pnPCBVI0bQw0SrdBeijp0XzMoGWSHq
nmObZIzM36synFku47UQAQoM1VhIVCgTpjFLvRYjaDhUdPESFK/HUq4sE6/vs7Xw
xKRjnavVocLhXxIYdQcJrPXiNhJuovZW1+jfOcvRRb4jJaJFRjgTMRMLEOfzcxgC
UhTBuuEFpUo/5sOeoVNMfTehVGalbQZ4IXfLeMH7bQBSi1RQoLosKNqPgUlfSRcs
sE2iqwvxR7EWilNgK8ca1AC1ruuE/mrMX+6KXAIKXMcO37cRKA4AN4nWLMbJNzKK
9dg1BE1tEN550mgcRjdAeQTOKZ+Nu9iuIxnZoRfOVPfc9+sVXYE9nYcLnLMXsdIe
NoyNBr5QrHvZOLA5xzmzMJgSvjVuKfbLWArEd0e0GqFtnOvq9LZTgG6UsATyTerR
uE4o32F4xU0OZb7PBCJ45RAIS5d84IlAm++CX+LF4prhr5Gosc1qWEJG612fVi15
`protect END_PROTECTED
