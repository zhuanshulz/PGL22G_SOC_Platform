`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CgUx7GdJpCVjH+jCwEA12HpsgeU/jUCT7/qKdlZl40uKucOARgOrOQ3vytax2RtQ
2jOZlvf2xI7RMSqKZD9yJ2ORaK/MhcSEfgkfJ4XM3Vy9p2cdqUni3d1j8Ri0QR1m
sMrXPGEC6W1/dt+tdXE351fjlMcOhQK59bbhcvqSLvBRNrBrDiv5Ysd/1nWJLWbf
ZOcBZb0AzlxZenmKIvAQ9IafoQDB+K+b31zUHPNwreFkAvcP+brSfzvAnh4RH+IP
kqeeJP613/29MLiSYrwGbNslGbIjaHl33vy/NN2aw0SU4M6nIekqp9QMG9C264ml
WHLJoRuvr21bLnDuPKKkW7bohHw/YGo4hslqhFZkQyp0r4TtyXUN4W9O/pLzYXGk
RhHqp8BtM5VKepg3jWJlEBW6Je8E+DTwB8gNHkSHOY23EOSsL0/yf+E1OWE1NsfU
Kv4YlWQnOTL3T1c2aJiLQe+rmc3dezyBdRTQx/3XVDQg72y0ydlLazBcXeIRsgq4
s6Z6+4kvCIr95eBXZh/cWTUJXvGz4MtIZPrPdQW8GII0bQimJ9ej5kNutju/1jAF
DArkkh5FHQIwFnolpKsnhHXmxTLqGSE4g3rHKJiqa4QRz5dXU+ZKVuorxmxWUXM3
TY4Oj5oti9Xmq5DmhHl0SFR2pKRAkidmC65Th/bY2GjrqXoWtxk1ft9REa0f1aZl
qEDBl1sXP3sHf2dSJGSLpuoDRhMSrCHpT9xaHO3oSieU0iQPEOgop1IY2dgEUtM5
6dREH1zpEF2jAd6IPUso12xLtP2EtAE8VZZJJO0/HFerC7D0xskOiftfZZh49AoX
FAOGJUlxp7j1eDEjfBdfoOKS1N5yXoZvrWdWLuCFGofbcl6iJXXcv2uCUOx9HZz9
HItHCHGmdz/jMyTGfwFOVpjSzsbxYvyJ4deD14X2X1tInkann1b8/Ua8zWPF+EuP
4a2u3zBCBtqUZXzMIjJET+nMNJsjSLdTX/s/9H8ZeREMIFnywnMZOpXASzNMaB+Y
uft562+DLyt5WAJiLFoycyZFRXbcn80YHqOXX41RhNmdSXHHA0F+sfKYvbMpbl2C
TdulfMkGOfAIAlW5j6bgsYKbmI/tV/M0RdbR4BEhzhvp6uKvVRzD2gp7+aA/3a6K
+ULrTp27rw0poIt2BWLW7pyfjuxRgXImj7EyUyo56LhfDxpT1TEjrdfikF6TOsFW
yLPmIxQJ1EJ2REjteHssXQzUH2OZ9SZNOrrgpoU9SESnAO7kNityUmhmUexwd3Jk
di9bJnpuryPh5mLD0NHMqjKWOagECw7eXXfPRKQxyBprstrTVvudvRqA88yUtJlt
p5N6AzNqtHahxWFzVmpWbdzdfwE3Q5ysRQ/urGt/HBkbuEHITldqhB1rUtztLZ/W
K9AhJmpYbhYYBUs4OzH98Inlhpu4sfg7rHzz1brxvYAKOt5KQGsF2XkAtKHojd8V
TQ9HCZNsIEOPmGSrWtIi8BqVG7Gtc6ysbXYn2brxfeSQ7xQPIBi2Fit5VQu/PpET
PtuzrpsUQYxiR/33LjIvAZRmFBeJpbKS9Ad8lOzPl+au3QUFfC7EDBoDpJEqjAfU
PRsZQ8U/gHnk8YZC7RpRWj2BO5lJZfBm5QCsC5Mct29dL9vVyeYUP3pTtQgcuo1V
kNbNvJmDSSHM0zisd6F5RudwfWcjO9IYG9b5x4sjtCQvJm3f+3lGrGnhNxtyEk1Q
bO2J9OJN8PAoRyYFNNtIuXp7rCANbi1K6kD0Mr7orDD7b31CG0w8UTSgLEJhGnl6
YThygDUIZxv/nIhp2o0fKITuQW4wCuxCWkxZqF00JOXV4YG7CfaHBlV+opk0yqQs
C7e7dea/L/TUXXGUT7zOCfWLwzF8q4LYq2FcFPL9SdbfaOQMoag0x7Zj7dUWkZEk
Lcet97M4aseUbBtEi+UFcwIXGg5vMZfZcw9w+fjDFWM4msO67DK99qEnmJZaHj6j
9o5zyh3aqM8hGTrgrhfh+LcfAkCHCikd7nbQv1jIonOJKqIwelTzQGvBryJyq87H
RnzZ5gJ/wLY3lhHm8Ji3sNkmXlamkbE0jd8ricHDXHkNJqvfOUoKJepX0RRIIkKP
uTa80/9UkJY2YhARPnfQbR9ub38RC5xLEwTE2xD7VAg=
`protect END_PROTECTED
