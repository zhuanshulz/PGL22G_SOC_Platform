`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qnb9GGpbPKG4LSwn95XOj6cQW33gsPHdI7yapo/H3DQcwShpLdouG33qJxbGIe+b
SzvR4BBBJe2t93Tj89nBizKYwr73ye6YY8Uk37VXpaPhjPqMzWrVfTd+hQ42Btzz
LGxFKGEZfKp6mkAUgiS8je/Em2qQcq3hlhOxXYUjUviqD2DBFUiMn3l/7XiR+SeE
V/0OcFjSLSDRrOkS0nFtMdLrc2Y7yBLYyXctlKqmFcEIQvg1WrvGHf9EuYtUUONo
rmDs9l46QewfV30/LYFzg3/Edk4QQQZ1deII5pjpsNeQ4A8/elW6EjCe2j5gEOII
iNHKqdbrL1ZdR+RBi5ijit5gZ0OwyNKpJZ04bTtdVV8dbOO80qaboUqnsoFe22rt
djKQ4Wfr2Oa8Irvy2mkds8Ngkz0AX9R6gZCYWgKiQEZRQmnpwicJZwEGCWS0CF0k
avfJk72FIkZ1tsDHfGz3pb7xBMBhh5mT0jgcirXYGMkfzoqBIhN8fboMAp0nd5WQ
sgDTskZwq0dVWF8i6B6Vy20twt697bcxTo3T3TP8sn81TUVJ0TO3hP+c6BQjCXc3
H4nIuhqLCELhWzf/Q0W9odIiOtNw5u83y3BCSNdRO3Z9wuFMalMYA3Dio0c8b3s/
8Cf12P76aSu3b5BpHcWBgZwsTS1qJFz3j9nzerFxNg9BkW8B5XAJzenJunPhKNuj
LBLZkTQ7GJ8EWblJPv4lWpa9npbsxxL85qho4ylHo5IkF0ctbpAy3vSeeetDjtKW
6rnW+nsenM7/10J0+5AiRGXvx8UsHjXPzKd1J7+dv2eXx1LFoDwOv94imIXoe/J7
gAr88s77cCIXoEisL/A86+giA3siNZoBl1HWZgC9QLa2INhb9UZ/J82uQFtfoiPc
a67Evhnmyct6zPGLqkc1CWNSwq39sqJ8tgXzKQDamQvNgZi6M/oxtT6pxrJ70hWz
DYT1VbrmetON0cOQRGBAd94CPWyJ6Sh4Vl3vOPDQywchiDeoHIZkuDCakA6BwyZd
TDCl1NaR/Lp+Joo5wDB6KttACEmWmOqqni57IyoC+YQgoRKMbzB0hjZSGQLsV+6N
CKFujXYkESZ98ENSSJH7pN+erSINmfqQIGdFmbuNHviwfdK73CyNlEPsysNWNsWU
8OEkn5wy/bMjWLLx4ZAZjiW1j4isewhFcZ4lHg04wFqwWdFPz0jOemdNW8Yn6mrA
6D854xDDdOzPoTArV7e6S5ih/bBMuXjWdkr2I6yLBY9PYqNhf0/NvgVLBABmnYNx
UF4N9PL6IqgNSvKK/qfO6yZ4PgjxPYvrR6B6HVlw9w+uKrywk8Th6uR486lIaz+k
pwOdXfcx2DeVgW9//aP/I8w/9e5nUgRnKklpPKgTVt53AYwPH/R0P16ne6RXJJo4
b75+SyaL+lnu/EugZPwTRVtImYlFz9rVEvvJYFWhuxo3Og+BH8P9ai90FoTj4bEz
73d/nt7t4laY8vdy6YHJp2RS2M2XRiZK1uSsXLjhRqIkrOockCG6tjvz6h/Jw96Z
bvkOdgBDmKhnw0qggnrSGltzrthaiI47SUh/9l9uhg/5Sp3TqTEly1ENmnFA74kp
OzdzosJHfeauURiYuWkQfDpCD/BnzGGd1MVWAaiMpIGMqMdBljswobpQTZA0yNye
gJiBaHMz9hS5lIBclUBlu7cawYMbSzBvDuPqSnyIYX8g9/CGcZZ3DB+BSBbNW3Zz
ZYH9m0ehiNDKeHguKpkZiiDxLymOefQi8Yh3buDAHJzZ821su8g34LUjCn45/txB
GRUGCHPAlwTNUHTdZ/5nEkugZkis3xXJ6WHtHVbl4JKuLUpJnnixflvRUTkZyIvX
h1tJw5H/Q8oHzB9uDo8pY0rYAglL0FvdFAnMoEB/vPcpxBMIzO7Uev61bzWiKNVv
ZCvS7DXsYTZCYfZQd5DiR+4j6YKqt0foA0QoasGO4XydpTF4BclrjJjlR2rIvSjZ
xoroSUtv0/MyHc0RjaAarnJZyxx6lc6dbiaDlkubinY7xqkuiZ4MXRWJ7neE2DKk
hgQbumaSYzvemhxlgcHBRzZD44TCvU/MvP3DenXqvr8bLoT7XboMYGVel7ic9yH5
KbPVYBtvGMKuCjuYjH8CdWaqq2QAFCtvCAzYzPGemJG+vCej+G2SAAP42/Gch8bQ
+d2VNgj3BovpcbDZqlhB2tr635XSuKRCJTN/8uQN42ukMpPE90tRzz8rNUdeLLih
URD5Yshe8RdQykCdmln2f28A3HfPKxAuq25W6u0DmX5guTEc5tuEkFmH/mKEQ0ib
IUDjH/LhTv83DQh2l6UH/dSuafeh+xhpK93mYEPJi3tjPojiUbRCEVSqbD5l4I99
2iK7LIPXGztIrS6QZgd75SNuubAbmfmwErV/ltVp4+KU1nN4JDUpxDBMwSGsga22
+qrVZHsMbfn2mkSskULyqWU25PCk5wzVDSFPRzdW7BmvsjW4CJfO/2r7sihycXPF
ihABwE8bwlkANj/Xb+R7YHNjX8m7xLmqq1YDuN84fpkS5n3QFh3H4vRNoFwHlIu7
pcpoILOKzZwAntwVyg7NphEHGKTda2t3MFJZJGcvf7hQticZTYsf+VJXAkPp0YQd
lgCmuxBG75Jo1TAHZM/z4Ygd7Z4An4epjZAnNs7TZyuCSxQ3hZPd+4zeBnq4D/2D
pitZrdpA67h8AbhtJtvMvbgRr+IQ/dAN2T4tY4yfFzRs5LNbLDn7B7byTzBHJ3nV
E/9MLRAUzpVdcO2ol+eu6uMen1qJf0eJWANtMe0vMBgBRwZ6tjVOYSofbh2g8GO1
lVupMiqepydaTKl2QSxzIGnpVJXcY4kAZtvocH3X+35M+IOZSy6ofbXIUG4fwC6D
lYHlzCui4GQeaO4KfuEtaDRddnqyvhfPWW818KVBknOF4SzF8+bPNZM+vh6DuIW2
ntu+f0wSR7n9HkhL3/9Q6lg1BrS6BZWDm6f6hZL2qPuGAkzacyyypR9kSpknxsB8
1QQ30OYZCs8czpE13iJlVPsbZynENnbHFWz8uGOvzZ1ygweRqwI68LW6vyaO0Oak
ufloQotARVSWHPoLxJ6eBi/WMYi/ym/+bkSrxK0QxNGOs2uClkP/tGyI8kk6GIv7
miWaX8qME8w7r0rflVbTZIMev/1g2qRRwgkjaQxJN4GFgYPrdGL0QSeAKRJbC8ua
DU922DnW7Er0Qbu6pmrujZ+mwnC4nNBor1mae+T+7w+M5T8UMA/cTEyz+A2wCPbp
XPQVH0jEWzsvISjIziTl+9FLCVglw7uly448hcF6HsBn4zIwJSV93j8Yt3cLfo6z
zMttqT9VR194hNfQwDpmm95hpJANhClGAmDigSRevxrFOJHHpXslEi59FsLyU1aq
rNbSz2glG4s0MB3mr5uETMm9O4oHkfm2Jy7EpueARZgV8eo9XbylNVsXBmmlLn49
uLSPEa5WqYJRcY3l1n/EoFW8kgC8fwalKei3DibcT7U7ajyVldKV3v1l94p6MxAZ
tXXRojqyPz7fmGqpagdRYKIS65wEBWsHIEdcvbhJhsMrwHlKJZh74KJz3NdZ1nBA
i5+xCQNPJjde9HaPY+mbKLwCjrHWvUiKUi7zBnXFD+lT3C3geu4+GtZxgFID9mJN
xFBXMvSrXoBz/E6/PBMwVD2IMee7HGD2wOCMZzUKaxz7AzoQDfgmjohNAeSashus
S+uVJzGVn7Uc2A1BFeV20Xf8KOmJCnaRSUmcO3gaGgZTrt9uUl14zfE3in896t60
5ewrPbZiir/U7xXg+UF8aEvuHvN0tq8XtaIOXKoL/dAze964QlQqbJewRkmri4vH
lLQ9sx5icN3LjP8Nw7eLK9RI4OzQ/iJmE/GNp3L5GwpypeNbVL0D5/wJy2AZ9mXh
QdoqX3VNdrfF2wWUUMi0HhIptIvyzTxGtdMjR3biAp7cnpowAhJXl0/LbfajE45w
3sTIoATb0IAKsmUqWxxdKYaO/NRnjYfh3zExUw4Eve68r3CAp76fHt7zoBsKl2NG
xDTzrE7XVI9GpsBWX2pKujA5voUcXot8brP4ZWDTAphtWsLvDa+WumxrB8One+du
aGAELr4wX6dllKy1KMdCOtSC3qrp0cR8LvAxvyrh8D4ls9bvLcP0Mx/kt9+ZRTjJ
bEFP0laCPdgBXlGCfrmEDovR8s+gtscwkmN7TTQqJL66NSNfiRbeI1xPmM9LYCbX
Epl+U71hZVnb+6dk3gIO5EQuqNGUzsloA1ksajpJfrHoPsvmBgU2o743O1o1X4MR
s7SRNeE1VnVDUpOwAMYR/NwzGCNd6sQvWxxy++VM7mQkylkcLkNl+BgU85TIWyjA
OoSfYkmLucE42XncqSByzqCtTDeIov0SDSrIhe40dTg6QkIpEdbXtpYFp0NiqrbQ
oFNpBNIWtz32XsEd4mdksNeczfHDmduwQwEMd44BXPBoyFlhay+7w0oTSo4D7A6L
qpVje/g6LaueRhYZmmIS1dHG+DgrpWR12hM1LnOT2f23zblgxmQOrQfp5a7oCIJz
d2iQFK2aLxgaGHj3WaVLIJ0GXK1K5XL1hD52/CLiK++wB60tcH7Irnf2byIKY/g+
oRtYY5/h3M4fowBftHEEx8YeM0Ao0s4TZYt8WFNzRTD0t/7hY0qoQMEbIfa9ZI5b
XEn2aTm862xuv7oM5jj+WRyBE8rduUCky7x5/GylMDMwXed8Wup85L/iRBxuMwmG
Jj4AjUA6vw74phPYOIQu5ieAtApYj3DnuR+YNR/AMQ9tIthJpXtWFvqUH8LS9AEj
6qJj3+/aeZV2mq7i/azTSFnX14USj6U5LFjY5vSDvcFT8RDPN3myrNvy6cBPjLOJ
yTpvW12sblPViI4+3ZG5vaDoIQdMfHpLXipSovyuGklA68yMIwDjjWgFfsxy0MPg
S4m/X28FrYQTILfJWS9oQcyYGMipxkTxsk6ZXaQy7wRIi1odf1xTyWeftlaiod+L
3FGUSsxCDhjMXtQ3aZO/kQ7wXrx832M9sFUDiv+Wmrs4G5xsoyufOW4keoaoiGlD
LIR86Nhk+V2trMoIH3SKUwZpUMQlYWvZrj4OVHTS02F0Ob9m76Lozh2LRlr0CEnJ
an7Ct2AVBPodquT1tQkkTFM0ebMOdoss4SCXPL8arl4OVAK3xSHpAe6a4QWtNsYF
8TWzSAi3rRrQjVK3PZerynCH7d2b5dubqiJC3xGyv6Or63egLsPuLlAA9kEQdMom
r0tUd3I3GNC/vYFHo4uejw==
`protect END_PROTECTED
