`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XGenYgxQuR82erCR8w4YPl9E+lnbaRKB3OHuKVnGyp2HemzDSoARFBXBn75wsG6S
D/SiaMRwRz6z+MFL7c5vDjT19KkQWR4VLzV3MsNU5cd/2t0OI8+P3UP3L7AbPw4o
7nKoe2AQW2FGNVbAanxoDVwZO06QsOmM8xpi9mFv/L7vOA7qh6ZqYAX+2ij+oZ50
/cslz8UBZZ1XNfWQKPSGDEuA8ySaBSIUYEMrLohRHBiboznUd1T+Lz2Is0U0hCqY
ylauO1lIpNxmlnsYiuhv6bBV9VCDdAs6EsSFj7hnWMVzUeWXhiPM8dpPCxnD+8QF
WYGgiDQlp5lMfgkfPXq00qUVfj22IeYWYKOuWIztvd7EqqlGp6rSME/S3lPP3q8w
Iq8Mk5VU/NfEHg/1/ckuLOTas2syMI9KnCr7dbETsnttpa/qNzUk7Bu+1gMAVYI1
6f4QkvnMI8WSecmUiOFPqb1Lljbv9a2cyDOAukwBp6bNHq04XsLK2Z3IWQypSPhN
FQyw96d/ewZAKr3wd0tv5NZLUHlEK4PhLOutFH68mQpIhwtDh61BuyzFVjb3Ndiy
qhgayrCLmh5e3iHJFDJoOP4xw8kiTQ9sLbbjmo2myMZhTMPJCUD1Be8udw4brTI/
I4wH/lh3JD5DohbdGHeFAURcX9uCfp3lw1MVgM2igi3KdBlK4cdulyZbMYlWsItj
MRHkFsgCXAn80zY+ZjzeglVYgqKg+CL50AkmUZ4OGhECULe2FUfwGJF8HvGB1j2m
OgcDvpEWWViyL/8eW2H6jHkkPOp8a5RnRte8qsOa9od79oPG19UIeqLoiGbSw3EH
Opa3UEy0Yw+t/+EF1vLOCbOohOoPAGpNw6g8NBUlLaY=
`protect END_PROTECTED
