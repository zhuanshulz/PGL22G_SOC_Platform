`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
80w6VJwysuVfFPfyfdeF6bzyseEhM8Rl5ucarLsmZEp12tI15pC1IKKrcnWiy7Zm
KJBbAuQPWkrC3Tifr+XqRSFJ95378YEAXq8bpZyS813tt0OHZYfDzjqz+X9SqRAM
ewvlyYnjbdQ7OQ4X/tiNAIKB0xpWsMEFEulmpIpl0hp0FLAL/NyHSNlR5kXFvER3
7yIicjBpMsJ3cizG3KrksTJWxOZBz8EwgeNYmVp4O7GvVg2x4QdRM6MuOz+glNVr
Zi1gQ6+8/5LUaiuduPoGd4+RSKMEDSE8ibeDsEhDHl6nfeMxCbmI0j2i04pGtIp+
Z+c3d8ssPP2oofAZX1Ky6f6/2HU3MYQZjUUXCVVA4QMqzvxLwftGgthd8+3IxXRl
7jBW7v70Ol+5tB4fGPCCC92hLFCyylk1bUHSM4jxRl8XxhiQdFnaphe2yxWvVAkw
Fmnc5tQgwTbcW/eRpvwZBvvItcUSPKGrWVjvTVAYlJb9N6fZ7ie5BWoaBwyzDdQy
7lD0zVH7uM4aXG34mjYo6n9mqdxpLN2sPRDnvU13hU4DRbYuI9yL0c4x/2wo5ePD
FZSrZGfNQGqcquFy5TjlYMnpZlEDmN1PBjXqgheHR1J1KBEcllhml0XDrwxu7D6f
KRDbzziMAheGgOEb9BJulEDTTm38pR9y3LUtdnmoiGXvu76gQ751uOfN9fcoEndp
4Glzq5ztTJA+DJrWeyrovkzxei7Ze/6rlUauebWpybmJdMlMicfLb0aNxzpmEI4b
J+jPpFIBFzpf398nrpN/bqRhiaimBbZucLw+lxuUGKgQAeNqwLDf4z6imdgTV7Co
SEUBIS9PJtKFVHga76W3GJYHoOBtXE0Gnb+BfzvPz7e4toSoa0QWJdv26izJjmOH
clFrpYvi4TEf4GcVZujnGa397725Uq6a6nEn+rcES5x4bcvgZ1jZZU7eOwgbg79X
dpZdMsoKlQgEAWt5zfkJ7gzzlHvHVKQIXWSv+BlFssTHMetSQI5kNK5jSpZK1gLL
DioGNK6gE4TVmneDqbf43axnN9hAkTx73HKEdf0ghaAufrLP697UNOxjv7H+Qvad
0z9GjJVC2g2nYIwOX+SabERVRdBAb4iWUQzrTYPs5ijHjrdsX3XGCOJ14y4Y0SnT
QHPDuGq3gHxAnmGbarU1yqgPBomCn+eiAP3gEl+44PHfBWJYA84ZpR272ldOn63w
2XkxQ43oD6/xQhh2jcJe2JWcxGG/PxbBkoVaGMIEbuUVe7oUJ9X5RltSkbEdEqkV
kF2s1+l9dpGfyQKUct+cGWfUUHSTxsVzOpyuTzJL8Wm8LqRaUbzMaGw38I8cHDw1
WtIMgrnxvGpIsqpnN+53oy/XlfmgMv/x30s/MPU/2FMJm/RFHTvUR/ecFegg4rDX
20iuMnFjiMe7jMrBdOmrTCLfApYIx5hiG7cl/tduNWvpW3+GEJFhKEQbEqiu9JN7
4h5B77/oWo+UulrM1uBvqa7ngIigAC1vnsBQoxF7KIgkzd02rGtwFfdqG5SOUZsn
RXtHZb1s17BWrZLBpiHHDQH4nJasXoyA1YxF7t1oLgxcXMKku4RUauPkCPMlR849
hyUVbMfVAnFYLiZi07sjTB8wKogKaVX9cBH8uViQbDOPOSISVmEWs8PxTBD+FSNL
chsJDhC7pLF2DJPe3bDOvOl+hmmCS0gQkzXRQa75a0HLxNdDayXAekQUK76U22Ph
9EE5m6y6vbSOD06TX70hpIzMaB5ay4PAFafEefvgKIWZmcCszpkzrog2QjFf7QLI
CiQsdW5MUFfkbkanu3G1OGuptb12xKRMlRL89Edi0/TmM6n0yEIjIG2fmZIGvk7U
o+P8cy4G87rrFr8N5wS0dyFgnUgBBtfVv8PqgQLfzH2cLIy1GOuJ6q8eRX1azQr+
yUbF1n+7kZRiVkRcLC4kt2dDx9IpFOEhob0GaAzd7+zjSJM00gaHmXdu8yF7+aNE
ddUJqZ/4O6BPpr0tgFuFVtv3AzowjjuOCrplPz3VHMLo4If0COmhSd4djepdc1nO
L8Muwz2tFRWx+Cmf7HtL/FFfyYxSLSA0wvQNvk2kNVj0Q+RADV8JnBo/6s4/BwJn
Nyf8jkugvra4isFV7doqk3MLS+Tpx9Xpd4n61wf1KBYcCdsv/lgXaqknAc7arsCY
VDhboFOlMcQ1SOI2n4TJruk5JPEBAAd4DrjOj9yb2zz5lFAEmTex19miC/BGdwo6
f2tcytHgTG0z+8+oZ1MzussgBduqqe6tVd/Y60WOmQlWZHaQlHBTJUtZPwL+m7I+
m4+UsX2OQ9iBhPh+symGccDlthWGe4a4DJbIVrvt7LGOSYeWQTCjGAPLzMrOUOTc
iAUf3NX2yqk2GjAVE/W7iF6XLnqWp4CpbNjZheJE89foWNw6ysyCfUqkON9zHuu8
0wMkZtrbg9Yxlh7Tz4KrgUqdRDMtNdbORPXFCXXs4GBZ/rYFTSFTU5e0obl59oLb
wKf6aFZCcqUbDtEw73bZ6uza3cNySskak3WBsTGzIJqSSQHlIIVFPRACb+vmMK9g
YSskL8shWtEttqIo0LNIGP7yt1unhrtsn4UnoqltKNZrzpEdk3XMYUjMTB/WC4tf
a2bL3Cx3Nu7w5vp0Ajr87bkvU3K9TogU+xG+/0Mk9KKTgnuFS3MNBfyIMZelVFQ5
SMyIZTc3pnrsBjnhrkOSghFcvVNRXICxqPaJ0HiPMM5rZaaUDht/PRJGQCLO3hO4
BzaDkM3XrtFIJI+juej7MYx2rrh8SXtkEM7llmbAwJFxO9XypwQkRanP/8+2QlFR
52r608K3sk2U1P3Gj5bfi5kiapNC8vfuZTefj7wNWAnAUuu9Qzoc7PezT4exISOf
OKBiY02pOumk36wORf/WCLVSOEIBoW4ctrI9kaKFXZ+82xWVE7BXvh0ZcJGYvo+T
`protect END_PROTECTED
