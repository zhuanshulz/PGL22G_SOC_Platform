`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8UYhjLX4mJgqH8oAFJxyXzFl2EgNU2vAYrslI7x4SpdWKxgU6cdirECYyogsW109
CJvVsVC5SLRMXSRBOlwLFWxcd1ML0p4ju47JzissUEaHbGKD9Sacm1D5sChkgnEH
ygDAGMfn7P+vRvMX7S/IpEjhlGC4J7Q922W6hM5nveXjpW2KDcHSd6laeCielYQO
OOlXYME+HPZO5NN2EGLEuss3yIiw4ompkoSYpp0qxlzk8BhEDlM8NmCFyAFk1mzs
3yxIy5BYfmKKsetD+UZYGS6nmQDHSAbMIlcIw0WpL1jvZoZ6ElzYhYSjPBjwN5LS
Fapfw2JUX/xIZIiL1J23dbiKBU7AErZScC1BQkZmMGh7D4WScQE5Gx6xO3R3ZRiZ
d2anfehUPhQQ0HY14vphmw==
`protect END_PROTECTED
