`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
83vkHFd1e7sjA8YvsuHqFB7pJDoM9OSvqHaxeW6jf3wLKrRP+uQHQ/aN/FJ1rBzI
JvDnoih9wbkf7cFEI5lbwv/YSfCh0hJQMLCgUcVQIJEFXgdzVFxlFxHnhkfZO0g4
Q6059UxfOEgJvkh6qv237+QkQfi1TM56zLCsAEZoCWr1O1o0y4TfVldfN5UALHMs
WoCdv7XeMJKjyFxxihyp+xdcGFAPm3v57azd0p9eUPXFIYxr8vtKKmSzyjNo7f9N
C6de21LYzarzoUBzArY/whUVEds2WSEXkw1DCBm11yhZLZt1DxYPCQlJJqr/iEp6
fpcp30WpqaHx0K73B5Jq69qHQfYuEjf54BgejRVB3p+RNkwjyMxyx8teXqlCW6yg
JRBtrFRiL+281WZh9vDde55uLn9FGUClU4rcsaYHisgC7QFuHjPleeLPTR9tXgq2
UVod1gru1LVAIj0zPm0+O2JGKCykVDBEMVWo/9UA6K0nbySZ14+B5aCU9D27Q5qm
WlghuUla9dPiTHyRqYwicXCbrBOp/QnDgSgvGJJ5LFSi/EAoUiOYTgZznZdwQke8
p7ap5J9TE7T51YTqDJDjcvVyms0Jk2494crDL6gGMxyDn53UFJ8OrFOPDrmFNPN1
rdUoOcGIJIKwqmIss2iD5aukbDtFtBiNE2am261hca10UXxJlNnpRO8uaEiyotTP
r4LyCHhoFl+4IVZHU3DmDMLtpjDwIROBBcBa28m+Lgd4BVWVGSdNMpDahQc368Oi
F39cYEKmSIX10bks1LaMtaR8lVd1Ih87cw+lylP7EAThnNeyeN6wunIByPv9Yhon
/OSrvLFC7qVVPSb/1P+EfSRVTtsQYXNDytQCfNfXUXMvvkg00l7DP6JCOIvi4DCf
/zRiGSx6ggQkDarIoAq91R+Zfnc+BEy/0ke+qnrYORTluGU9501aVpvEhLvLaPKO
FnjzhmpGiNxgnDygZo9pvy8X5QYMV/gypnMaq19fMQi+1wiQYsXUWtYrr8OwUX78
QeKAsuJXtsJut73XnGJxZGeH4su2CXroKEsDZjBu8HKMKEkjQB3oG1gtxPQbncGg
8J1JoeTYDRHiNlZR24VAFeUYQELMgmX8wbPFbjF/2pt7cmKPW6+bPLwx+pL1y9FL
quEhBbyvfh1FMz04esAT4nLJG41UZyCb06yZRsRhmySuluvr6Ov3763EHP44GH8c
zvoJT7lAP7zNb+6eSDIxuz7kiZfl2uHi8vNAiAPwbzNyrNFXMiZieF7RBwm8LDfq
`protect END_PROTECTED
