`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QxmsObKJGZ3DRmwTXe/DD4HtKvPyGxXjqyVaQMsa9av3iTWpmnlsF79GMiHXByGz
SIcxzHijojaEA1UhLwYkIaByj1/zvQQ9ejohYOr1KUnRu6aYi3xaohnHZrRxtcZu
kNCIIhK159S6HJU3imB9MT47D1pCjUpvSSI0amOvXFeBOwLCO4JKx/tUSj75K1lH
zKVfqM6/sLHDa/uNEVgFUujfotdl+rG7aR5PnGB0QQw7TK+K86nBECghIh/wR1Q6
8/4/Zz0vUGFKARqa10m5lS/QHZBvVJbQhbEpvDpJcQRadt/PBR3HlLDnGmtCrMn0
JIaazW2rF1ORVxm5qg9lYYZmIFCP++D5HN2fWGcA2Nu59FSkP6ut8RMoFCk5kgp6
3JnKCq1apiTJX4t/lDu/T3VeLKjBL4/0ugD/41SxpZS2mkgaPI7ZyGF0uPt6pMvv
rU/AP2KvLz0TL1EYfeXwP8QkFyuzit+rIVnGOojz/V/0p/8S6R/vUce6eMGqTToe
y6vXgQm6duow8rsWOpKTLRQ/Qp3+pBrmLi1Hzlm48OW82WB0LWoB9SCL5VZruXjt
dx236zsiQIRkZUaDKeWziXiI3iEuKoAKXFAO1WW1gATOtiQ086Aej7szLDRSw8Ad
FYvwAxfgyhC5q/Mk7768sbVXxTyH5TlsuZv5oK1lYsQornkYFcBHTpGK/aggRwMW
tILCLTzKIGO8oIxgJbThWVzLVK1HnlJdaje7NTDACvTuzG39h/09wkcxy/BNGcje
4J3E+5/OXcw/Gdjx5YRoCSRV6tt9z82p1NDheX/05arNgoU3lBQ2g6/NFnuvmekx
mEzqMywFxyd0y+sJw4QucBjHtNsExZUagTikXr9i+eG6UipzHvaWPMkOpHclhTel
cJ2O0tZv4sz88vPzu+RO1tohbf2NhklpT5wkE1LxeGV1/wGaO2uOJHSRLuFs0yul
OUgaBATSzFb5hI0ePpXbQw==
`protect END_PROTECTED
