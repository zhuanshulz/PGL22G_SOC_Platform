`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uGTPHCNKEBBLuysVWfxAgTNhsE0aBHEzCiFfTBEe5XBxsJ96NPOFFHYs3mDol4oQ
Bz/8jAlF1EA7Wy20+qL5bhK0nrSvyLIgrkJLc39D8SRxOr5lthDew2Mxygznt2RV
W+ZtXZ2CEfB5rVUNJBM7vMKJS4rAsElpLsITJpTP0jkwiNv+P91GCUj76RvDOv7T
i6aWjOThk+hf9f5Jaw7qaxMysHFwjAXWJwsufsPR/FTnmP3FbwuetZKIRCF4XY3V
ub+logDy8oOR3DrW5JQHoLj56++Kby2l7EXgkEMpe9h/KPIrIdZV3ntF9BJn+ldR
eokeQB1d0HJtrbV/e9UjQOniSL3WQpvjSEH3oGKhcTwmYW7Op6dBkgvybDBvX3B5
i4fBBFi8YMYCVk5HYl/KkxUIaVUVUUDRgG9SZFUumqE=
`protect END_PROTECTED
