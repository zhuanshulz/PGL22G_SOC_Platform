`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
27jn+JpVpuqO13vLQMk1g+fM+4MB9P4oKth1Ei1RkO7+DRKoHDsNwzeRsKU3Envn
/aDj7pC/4zKDFvxd29TIV2EwosV3UamjICGtQR181UOvYe67cfua+Eu7zTWF5mUP
D1ibgCCzC/ZkMDgnUtuxive31fr2y8dHLNkPWEolqlFL93T4y5WgqZuMLQUt5dz6
1N1iXny42YIqbZVEUrKlzyDy5ipCsXxsCi+8rhy+kw4rtTJ4HAH1emFRxll9q3ea
qCGOMfC5bcrPb1Sz5e81I29FqGUY5zC2sw6y7a31rWFWS9BsLz+c2kLEJiPsM7ZW
GfvbiCfzkDLdPntH++TN2p+imTE0JGntPox89p+DEF1KBWf66Vp3AIB25otSiNpk
`protect END_PROTECTED
