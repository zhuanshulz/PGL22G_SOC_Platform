library verilog;
use verilog.vl_types.all;
entity V_DDRC is
    port(
        SRB_CORE_CLK    : in     vl_logic;
        CORE_DDRC_CORE_CLK: in     vl_logic;
        CORE_DDRC_RST   : in     vl_logic;
        ARESET_0        : in     vl_logic;
        ACLK_0          : in     vl_logic;
        AWID_0          : in     vl_logic_vector(7 downto 0);
        AWADDR_0        : in     vl_logic_vector(31 downto 0);
        AWLEN_0         : in     vl_logic_vector(7 downto 0);
        AWSIZE_0        : in     vl_logic_vector(2 downto 0);
        AWBURST_0       : in     vl_logic_vector(1 downto 0);
        AWLOCK_0        : in     vl_logic;
        AWVALID_0       : in     vl_logic;
        AWREADY_0       : out    vl_logic;
        AWURGENT_0      : in     vl_logic;
        AWPOISON_0      : in     vl_logic;
        WDATA_0         : in     vl_logic_vector(127 downto 0);
        WSTRB_0         : in     vl_logic_vector(15 downto 0);
        WLAST_0         : in     vl_logic;
        WVALID_0        : in     vl_logic;
        WREADY_0        : out    vl_logic;
        BID_0           : out    vl_logic_vector(7 downto 0);
        BRESP_0         : out    vl_logic_vector(1 downto 0);
        BVALID_0        : out    vl_logic;
        BREADY_0        : in     vl_logic;
        ARID_0          : in     vl_logic_vector(7 downto 0);
        ARADDR_0        : in     vl_logic_vector(31 downto 0);
        ARLEN_0         : in     vl_logic_vector(7 downto 0);
        ARSIZE_0        : in     vl_logic_vector(2 downto 0);
        ARBURST_0       : in     vl_logic_vector(1 downto 0);
        ARLOCK_0        : in     vl_logic;
        ARVALID_0       : in     vl_logic;
        ARREADY_0       : out    vl_logic;
        ARPOISON_0      : in     vl_logic;
        RID_0           : out    vl_logic_vector(7 downto 0);
        RDATA_0         : out    vl_logic_vector(127 downto 0);
        RRESP_0         : out    vl_logic_vector(1 downto 0);
        RLAST_0         : out    vl_logic;
        RVALID_0        : out    vl_logic;
        RREADY_0        : in     vl_logic;
        ARURGENT_0      : in     vl_logic;
        RAQ_PUSH_0      : out    vl_logic;
        RAQ_SPLIT_0     : out    vl_logic;
        WAQ_PUSH_0      : out    vl_logic;
        WAQ_SPLIT_0     : out    vl_logic;
        ARESET_1        : in     vl_logic;
        ACLK_1          : in     vl_logic;
        AWID_1          : in     vl_logic_vector(7 downto 0);
        AWADDR_1        : in     vl_logic_vector(31 downto 0);
        AWLEN_1         : in     vl_logic_vector(7 downto 0);
        AWSIZE_1        : in     vl_logic_vector(2 downto 0);
        AWBURST_1       : in     vl_logic_vector(1 downto 0);
        AWLOCK_1        : in     vl_logic;
        AWVALID_1       : in     vl_logic;
        AWREADY_1       : out    vl_logic;
        AWURGENT_1      : in     vl_logic;
        AWPOISON_1      : in     vl_logic;
        WDATA_1         : in     vl_logic_vector(63 downto 0);
        WSTRB_1         : in     vl_logic_vector(7 downto 0);
        WLAST_1         : in     vl_logic;
        WVALID_1        : in     vl_logic;
        WREADY_1        : out    vl_logic;
        BID_1           : out    vl_logic_vector(7 downto 0);
        BRESP_1         : out    vl_logic_vector(1 downto 0);
        BVALID_1        : out    vl_logic;
        BREADY_1        : in     vl_logic;
        ARID_1          : in     vl_logic_vector(7 downto 0);
        ARADDR_1        : in     vl_logic_vector(31 downto 0);
        ARLEN_1         : in     vl_logic_vector(7 downto 0);
        ARSIZE_1        : in     vl_logic_vector(2 downto 0);
        ARBURST_1       : in     vl_logic_vector(1 downto 0);
        ARLOCK_1        : in     vl_logic;
        ARVALID_1       : in     vl_logic;
        ARREADY_1       : out    vl_logic;
        ARPOISON_1      : in     vl_logic;
        RID_1           : out    vl_logic_vector(7 downto 0);
        RDATA_1         : out    vl_logic_vector(63 downto 0);
        RRESP_1         : out    vl_logic_vector(1 downto 0);
        RLAST_1         : out    vl_logic;
        RVALID_1        : out    vl_logic;
        RREADY_1        : in     vl_logic;
        ARURGENT_1      : in     vl_logic;
        RAQ_PUSH_1      : out    vl_logic;
        RAQ_SPLIT_1     : out    vl_logic;
        WAQ_PUSH_1      : out    vl_logic;
        WAQ_SPLIT_1     : out    vl_logic;
        ARESET_2        : in     vl_logic;
        ACLK_2          : in     vl_logic;
        AWID_2          : in     vl_logic_vector(7 downto 0);
        AWADDR_2        : in     vl_logic_vector(31 downto 0);
        AWLEN_2         : in     vl_logic_vector(7 downto 0);
        AWSIZE_2        : in     vl_logic_vector(2 downto 0);
        AWBURST_2       : in     vl_logic_vector(1 downto 0);
        AWLOCK_2        : in     vl_logic;
        AWVALID_2       : in     vl_logic;
        AWREADY_2       : out    vl_logic;
        AWURGENT_2      : in     vl_logic;
        AWPOISON_2      : in     vl_logic;
        WDATA_2         : in     vl_logic_vector(63 downto 0);
        WSTRB_2         : in     vl_logic_vector(7 downto 0);
        WLAST_2         : in     vl_logic;
        WVALID_2        : in     vl_logic;
        WREADY_2        : out    vl_logic;
        BID_2           : out    vl_logic_vector(7 downto 0);
        BRESP_2         : out    vl_logic_vector(1 downto 0);
        BVALID_2        : out    vl_logic;
        BREADY_2        : in     vl_logic;
        ARID_2          : in     vl_logic_vector(7 downto 0);
        ARADDR_2        : in     vl_logic_vector(31 downto 0);
        ARLEN_2         : in     vl_logic_vector(7 downto 0);
        ARSIZE_2        : in     vl_logic_vector(2 downto 0);
        ARBURST_2       : in     vl_logic_vector(1 downto 0);
        ARLOCK_2        : in     vl_logic;
        ARVALID_2       : in     vl_logic;
        ARREADY_2       : out    vl_logic;
        ARPOISON_2      : in     vl_logic;
        RID_2           : out    vl_logic_vector(7 downto 0);
        RDATA_2         : out    vl_logic_vector(63 downto 0);
        RRESP_2         : out    vl_logic_vector(1 downto 0);
        RLAST_2         : out    vl_logic;
        RVALID_2        : out    vl_logic;
        RREADY_2        : in     vl_logic;
        ARURGENT_2      : in     vl_logic;
        RAQ_PUSH_2      : out    vl_logic;
        RAQ_SPLIT_2     : out    vl_logic;
        WAQ_PUSH_2      : out    vl_logic;
        WAQ_SPLIT_2     : out    vl_logic;
        AWQOS_0         : in     vl_logic_vector(3 downto 0);
        ARQOS_0         : in     vl_logic_vector(3 downto 0);
        AWQOS_1         : in     vl_logic_vector(3 downto 0);
        ARQOS_1         : in     vl_logic_vector(3 downto 0);
        AWQOS_2         : in     vl_logic_vector(3 downto 0);
        ARQOS_2         : in     vl_logic_vector(3 downto 0);
        CSYSREQ_0       : in     vl_logic;
        CSYSACK_0       : out    vl_logic;
        CACTIVE_0       : out    vl_logic;
        CSYSREQ_1       : in     vl_logic;
        CSYSACK_1       : out    vl_logic;
        CACTIVE_1       : out    vl_logic;
        CSYSREQ_2       : in     vl_logic;
        CSYSACK_2       : out    vl_logic;
        CACTIVE_2       : out    vl_logic;
        CSYSREQ_DDRC    : in     vl_logic;
        CSYSACK_DDRC    : out    vl_logic;
        CACTIVE_DDRC    : out    vl_logic;
        PA_RMASK        : in     vl_logic_vector(2 downto 0);
        PA_WMASK        : in     vl_logic_vector(2 downto 0);
        DFI_ADDRESS     : out    vl_logic_vector(31 downto 0);
        DFI_BANK        : out    vl_logic_vector(5 downto 0);
        DFI_CAS_N       : out    vl_logic_vector(1 downto 0);
        DFI_RAS_N       : out    vl_logic_vector(1 downto 0);
        DFI_WE_N        : out    vl_logic_vector(1 downto 0);
        DFI_CKE         : out    vl_logic_vector(1 downto 0);
        DFI_CS          : out    vl_logic_vector(1 downto 0);
        DFI_ODT         : out    vl_logic_vector(1 downto 0);
        DFI_RESET_N     : out    vl_logic_vector(1 downto 0);
        DFI_WRDATA      : out    vl_logic_vector(63 downto 0);
        DFI_WRDATA_MASK : out    vl_logic_vector(7 downto 0);
        DFI_WRDATA_EN   : out    vl_logic_vector(3 downto 0);
        DFI_RDDATA      : in     vl_logic_vector(63 downto 0);
        DFI_RDDATA_EN   : out    vl_logic_vector(3 downto 0);
        DFI_RDDATA_VALID: in     vl_logic_vector(3 downto 0);
        DFI_CTRLUPD_ACK : in     vl_logic;
        DFI_CTRLUPD_REQ : out    vl_logic;
        DFI_DRAM_CLK_DISABLE: out    vl_logic;
        DFI_INIT_COMPLETE: in     vl_logic;
        DFI_INIT_START  : out    vl_logic;
        DFI_FREQUENCY   : out    vl_logic_vector(4 downto 0);
        DFI_PHYUPD_REQ  : in     vl_logic;
        DFI_PHYUPD_TYPE : in     vl_logic_vector(1 downto 0);
        DFI_PHYUPD_ACK  : out    vl_logic;
        DFI_LP_REQ      : out    vl_logic;
        DFI_LP_WAKEUP   : out    vl_logic_vector(3 downto 0);
        DFI_LP_ACK      : in     vl_logic;
        PCLK            : in     vl_logic;
        PRESET          : in     vl_logic;
        PADDR           : in     vl_logic_vector(11 downto 0);
        PWDATA          : in     vl_logic_vector(31 downto 0);
        PWRITE          : in     vl_logic;
        PSEL            : in     vl_logic;
        PENABLE         : in     vl_logic;
        PREADY          : out    vl_logic;
        PRDATA          : out    vl_logic_vector(31 downto 0);
        PSLVERR         : out    vl_logic;
        AWPOISON_INTR_2 : out    vl_logic;
        ARPOISON_INTR_2 : out    vl_logic;
        AWPOISON_INTR_1 : out    vl_logic;
        ARPOISON_INTR_1 : out    vl_logic;
        AWPOISON_INTR_0 : out    vl_logic;
        ARPOISON_INTR_0 : out    vl_logic;
        RAQ_WCOUNT_0    : out    vl_logic_vector(2 downto 0);
        RAQ_POP_0       : out    vl_logic;
        WAQ_WCOUNT_0    : out    vl_logic_vector(2 downto 0);
        WAQ_POP_0       : out    vl_logic;
        RAQ_WCOUNT_1    : out    vl_logic_vector(2 downto 0);
        RAQ_POP_1       : out    vl_logic;
        WAQ_WCOUNT_1    : out    vl_logic_vector(2 downto 0);
        WAQ_POP_1       : out    vl_logic;
        RAQ_WCOUNT_2    : out    vl_logic_vector(2 downto 0);
        RAQ_POP_2       : out    vl_logic;
        WAQ_WCOUNT_2    : out    vl_logic_vector(2 downto 0);
        WAQ_POP_2       : out    vl_logic;
        STAT_DDRC_REG_SELFREF_TYPE: out    vl_logic_vector(1 downto 0);
        PERF_HIF_RD_OR_WR: out    vl_logic;
        PERF_HIF_WR     : out    vl_logic;
        PERF_HIF_RD     : out    vl_logic;
        PERF_HIF_RMW    : out    vl_logic;
        PERF_HIF_HI_PRI_RD: out    vl_logic;
        PERF_DFI_WR_DATA_CYCLES: out    vl_logic;
        PERF_DFI_RD_DATA_CYCLES: out    vl_logic;
        PERF_HPR_XACT_WHEN_CRITICAL: out    vl_logic;
        PERF_LPR_XACT_WHEN_CRITICAL: out    vl_logic;
        PERF_WR_XACT_WHEN_CRITICAL: out    vl_logic;
        PERF_OP_IS_ACTIVATE: out    vl_logic;
        PERF_OP_IS_RD_OR_WR: out    vl_logic;
        PERF_OP_IS_RD_ACTIVATE: out    vl_logic;
        PERF_OP_IS_RD   : out    vl_logic;
        PERF_OP_IS_WR   : out    vl_logic;
        PERF_OP_IS_PRECHARGE: out    vl_logic;
        PERF_PRECHARGE_FOR_RDWR: out    vl_logic;
        PERF_PRECHARGE_FOR_OTHER: out    vl_logic;
        PERF_RDWR_TRANSITIONS: out    vl_logic;
        PERF_WRITE_COMBINE: out    vl_logic;
        PERF_WAR_HAZARD : out    vl_logic;
        PERF_RAW_HAZARD : out    vl_logic;
        PERF_WAW_HAZARD : out    vl_logic;
        PERF_OP_IS_ENTER_SELFREF: out    vl_logic;
        PERF_OP_IS_ENTER_POWERDOWN: out    vl_logic;
        PERF_OP_IS_ENTER_DEEPPOWERDOWN: out    vl_logic;
        PERF_SELFREF_MODE: out    vl_logic;
        PERF_OP_IS_REFRESH: out    vl_logic;
        PERF_OP_IS_LOAD_MODE: out    vl_logic;
        PERF_OP_IS_ZQCL : out    vl_logic;
        PERF_OP_IS_ZQCS : out    vl_logic;
        PERF_BANK       : out    vl_logic_vector(2 downto 0);
        PERF_HPR_REQ_WITH_NOCREDIT: out    vl_logic;
        PERF_LPR_REQ_WITH_NOCREDIT: out    vl_logic;
        LPR_CREDIT_CNT  : out    vl_logic_vector(6 downto 0);
        HPR_CREDIT_CNT  : out    vl_logic_vector(6 downto 0);
        WR_CREDIT_CNT   : out    vl_logic_vector(6 downto 0);
        SCANMODE_N      : in     vl_logic;
        SCAN_RESET      : in     vl_logic;
        SCAN_EN         : in     vl_logic;
        RESTART_H       : out    vl_logic;
        TST_DONE        : out    vl_logic;
        DIAG_CLK        : in     vl_logic;
        FAIL_H          : out    vl_logic;
        HOLD_L          : in     vl_logic;
        DEBUGZ          : in     vl_logic;
        DIAG_SCAN_OUT   : out    vl_logic;
        TEST_H          : in     vl_logic;
        BIST_CLK        : in     vl_logic;
        RST_L           : in     vl_logic
    );
end V_DDRC;
