`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2nruY3OZubDbRWVzGLxpyoFSIIMvUsNdhOqPHQXSzUJ5UgmW1iou8ipIsmwliJUq
9d9BcZ1wvQXvtjPcHkcfctRV85teKVBUYuC8PJnVA1AOSpjnsEkJPoyHTKGEa0sl
8jTaqoCk9A8XbbjrOiok5+7gBob14thVPjiVtc1Y/AVhkRnFRGuNVQIZP6nxIQqf
Dt60ZUT14+BL81wUAsGdJOQJzmKot2lNwcZZRKjwrp+gtowAB9mb/dlHh48M5aFc
vqZkpLHrddf7576mDWS3IfgU2UEG+GSMOr/w22A/f1igm/z3RX4ICa9uJfG1Hd0k
fm5kig3sydihWO1MrRd+z7J6hzqZxZeXPF5QG37mb7yRo8QZ1Jkyl0vEiys6h6/K
VXk0zAz1WaoCK15t6c3qqNuYmqAQVZ4jS6w7cHgCY3CCroefStk+QOPhAbopTXHi
CSS1iPcHXRvMO3tn0PAk7h4Tr0d9AoBdxygg2wSPXYugMZg4iejtKxL0ytTI+5AJ
CD2fVygSVT4yFIqfjfAscoe3bQ7xkeiF5Dd53VsbGu+xi2MX2ibZ7JN/zX7Hxnag
nrrHcqpQp/3zlVrBZK0MHKAmc1Hmf5z+aySZK9w39MZK8STyxIWMaCJYJnsYCsW4
0MuEB+ZI7UZdWboLTbSKkcHbFhE7rwSvLE63KhY0IsEKBN2e51dNxnZPDkf1wkCW
sP/Ao/8eWQp4hZ9aMcoAVp/8nf/3+K+31yZZZlEJGPW9NiDeTLZ6mxQ4ixbUuQXl
gOcioA+/+sb/qeZlGXUJ71Hy530Yv9UVB0EtpBMiq2PGMNoaeGhWfVgDb9UTLyt4
p2olYbf4B+G0PoTOcSb2UYXkvM+wPdWvs6L1Qle2OKDVPbC6QHXBx5Gz/7UzR22C
BYqbSrg0wiwJV1NbQ8ymD08Gror5QZ8AitLslrHs5K/LoMNNm9lgP8fe7UnHwJjE
ydaZvgvzNO8WDxzkrDiEai23Xau6V9lmcpHebCxx5VAyTuO5rV9/zNWAcZub05Fq
hXQHXcDr1HPZ0dKOmL9duOpUXFFolP9E2BrCdDrmW0zs/2z4R0Y66QirSEmyshmN
7Jy4LLkDIIta0gw+Mfs4g1z+iiEe6mjwvQcyGdx/jNfwem/WuUGkl/YcKIUczOg3
kFLktl1cuGm7NmRFcFinRB2f7G/7m/7CU6oAQWloJJprKGQV2n9C36Iqs+o03OaA
Tz0lbj1b7/3FKw03MeBEpP1voE20RUar9DwL6/4ZQac=
`protect END_PROTECTED
