`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a0eVwsJ1/HaOUpxiNQloaZWp4UGm83Dy4TiUFi++hZ1JpsA1KlNwryDhmNbuURgB
9chUe5Re/MMMJRWY83HsSvaV0+Rp4IK3C9KzMMbdoFTUwtO0owIxeLo7D9kPzG77
3cEwH7ggYPmPOeCideFBXLiznnotvR7WWcKHCcfiPLnXmoAC7DW3iEnuKID6OBtY
Yk06eVTbx64QoMF5twKveI1dxUGP4WwwIFBHKr7i4uWX9h/p6Sq0PNrEjCcPYs9R
6R6zQT5bNoR16kEAscs4MyBYu5jP0+6cu9B3a4nHWKh3KxaI67+jUTK/6dsTn4Hw
ns1wTyRV+oZQQUM/5+0DoFaANvB6CAa6EjoQeqy9LqAPC+xHDpmUFep2MX4J/Asb
wAnmN4qAV1CXiNwWCKgLT6IXpqd4pV+KTLdNL9fHoxk3FUrd1FXK8O1j4NUgzNY6
12BRG/A4mSuIUv91VAte9SkQhdDCaee+OTWfsyS+mMzc8rM8hCKD49uf7ttthXLl
jDQ+LIUmiQYbyWzQFCvXcwwB/kBpKJpMLrr6LOpsEQ9VPesW7sv/DnWAiBo3lEI/
Gr+PVuXbXYuiEkjEtWqylJ+nHK7ruVnvoWcoIMYtOSiZuPjAPao7DTIjECAsBeVz
eKGUILy0SMY5RAjQs4hz2k34PZA3g2hzsa+oPqhErAozArQC4QDOIMVRzuhD+KkY
Aw0KcOczxDDgi2qnrklEr0hRSve7IO63opdCL1Z32aUn5Kjdgn88q8nv4BqHgvdZ
u1BDRtouoRrXPwBSxSWDH2msQhMJvfhG2j2tg+/lB6htZbyXa8bcSilPHlHntIXF
WsWYvO/1PgZvR6W+BcIuqicdLUfUJ1GuKi8HUBXkMmQSdH91AnqN8eSf8Un9rTGf
CSR9Uu39ICoY6sjpUxAGKbWWUqkpLNP7YVI7XXB4TGuvDGk5aMJnu9aKpfntIKTg
oWztuwJTWr7bQCCoHkAdxjMhChUgaUfLf8RLzLoc5es/hVLsJ+l79OAGTiNbcBFm
liPunOwnKTcuqzxykn+Ak5Y/6UtpBwUkPDL7wv3b7t1c3kdHz7GGEI5Zoe7c3q5U
wZ4h5DJ4x9p4alawVezshk2ev0SNSosxPgNT05cXtylA9ZnZlgiVZq5biGAhZSUs
ZAW+lXH/lufUuGBMezM+dLFHpwBNVvItTBs20WQUOIa0tJ9DGFCb06lRvp4TRNHN
qqGfJ8gKz5qkOfzVNiWzKApmqvHOOFCggpxG2iHQ7kU4x/tX+zgS9IZi470gAC1I
SRq7mmrq7wMcnqyjeNqB6mWNz0J/Vey+tVzaaRkBOxaETieRIFzpHwC4iZ9KM4xw
veQ3YJX4FkaFxwBOOABBQ2BRn0IYNrxaFJL9ejHeS8+1a9Q0M30MIpOgiO7RmO9E
3Crz63MXSkPd4Oqp6pTdZ3FyOd2gVmsGlekE+bNtPVBaShNhXzSWTR/KOfBH5b6E
`protect END_PROTECTED
