`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jR7Nn9SvfnWhAT2KuJnj+zLehE1NYNGciPIzO4rI56RRNCAoDkGWnoavL8wpYuZI
BSpJ3T8qzB2sOh6Sg+pjgJRWUsw97mZzoB4DzaUi/Y5Cz4W6w52FBg0HGwmAqBDJ
nTOJWtERzxucVzwh456IM73m680/3P3FLefsr1KXqDezEZs/TNweZqPEY5e7Hg/F
NEVqGk5x0QQozmIkrSfPLGjRcs5/XCVEG2fWBH4SDQabRELSYVPb/EAacgjcYhMd
VwU5+XCc3Gd5VIgq86/GTUMSdd2+1PfDlBjZUSl5RTdjbzgUH1YPiEDhTZ75OxZ+
1oLAu40qXpAETGGvfb+TzNlczzv6yC3MdIRhEy0ir6dvdCyyOlCujKowrHOmfj0r
WL4H+RB6hSOCGg6wa2Pn/HTZkwt/0lXaV2ZxZhQfidHbuM0XSnAbvKRE/tr4jfr+
rnP0WHRadcUG4FgtTq/hQLBdkLGAmJzSf0hLs+6/o1JfhgfEtqB92OvBdqNQIDc4
Fyc+zKzUL6xJtkRiWpRwJkUbS+ZSSJuwaDCGSbqm4OJQLw8Dv5ykKTxQ2O9K5E6D
LeQLhtudTkPP4k+VLoLHgr692eC120GHJhfIGES6ywikOun0SJr8CGn5wppBNpgu
OsF0tJbO26e3uLXpa0ZHjbAkRqTFeFt1B1d99Kql2zlcsd7lnBHfAfS+dcSkdVQ1
9flv3j3DgUYRC8ICGLWG0JNAFYHdzZZy4k3Ks3yLcIyAFBQq9qz4KE9gz0VP3eab
CecvVOMh34tyCJv557N0+iM1dG3NRaJHxexDa7whNZgpcZCWd0tcK6xBU/eJPrqI
ZntgpXG9T3I2ExHenKXmZKQFTrZNw07TzvKKs2pQbQJ4JxEgaUasCThLb+4I0o6Y
UeAaGkh2d6pTkdzgM7KdALT3kjDYhot3YxGnt3B92wtAcggwIbDctSNecbonhFcM
Oj2U3ervDrKk7eugvKm2/SmPz/LVasF1Hx83dRTJI2n4lT5rfYfL3ebCPCSundRF
FnIC81OgLzTO1AgS3Mojjk1JLjxC9XSLi9qMgFvHYFdh2Lr7QOzVDl761KATPwHE
zPe+3VoqP8jNU/X+moy4G7H52ApxeGoIf6GazyXCjTAxH32uBWHQEC0Nc3vgtdJd
KfQYwFHLOZTZJpLmAIqrUI3uy1ItqGrIzIwWdbcA68Drd8a4AgSybXSRwHLTMzPl
XDf3BQ9NooAF1m6kE8qMjIuavWKd3IwCt79BDK+QMOeaQhKFn/xX+ligNof1uL51
D97ojk3XfVyTWsWuPDg5upDDhxLYbf+S5yw9SE+/1ODT4ZUwtTa0UhFd7e7uud8R
+zWUMPRConOV3wMd8mqmNKHdtw8vAfmcMDBPpBhh4sHD4c+RBvlyC3dgn9r/QJLW
YsQGKRD0/fPA4Ca634SphhMdcBOSYygox/WPSnaF57rXDRnnQA5fh2f332hQeuyY
O9tquDCOW1x6hjMa3S++YoTQUHFdTYUfJOaHXTKnTVbIRpIp6s/f/yfAdpYZWJoC
lt4l7N3FR8uduN1FlGk5xweneBKrsVhMoC4cpHnonR0Mg/QZog3P+lwbD2zMayJH
rJ3u5UX4lHXhYzLTT7gKRvEdHXgY49RxpyaszKk8ugRuOVmXquDgk8ypO+3OnDjB
nz94b+AcADAL6IUU6VpcQclzUKNWpvX/J2QhlRMQOl8A6N82eOV/ZRHCiN1JXSxD
XbvhYlVWN8p8uUqb+GSRPEJc5B4wKRa2ZIqPPgnrty+f2wWuZWrYOBXIRpFjwnVq
lb9wi0+eeG40fiVM8yRBISO1g+s86plC07MR+X9ahFkW+CP4Sc2cDCUjcYRnxT4O
iNv3daGgV+WaLOshx0GO7kFBOtRusB0Ce4rGrabtKxqnC8Qi8jSCPouXGVMgIP2C
EWynBCUZABuEf5X/avZoFB8Xoi8xbUniuzkjBs2Q/q/lg2T36xkNLzMzn8yOy7MQ
pw1LYNZp3yImkQP7lZXZskTtCH/w1kWmQz48yiLX5a5i0cTJJPjkG+c/H/US50HG
vNpmM74Ks8zvzLdoWNQdfH3ct+PegalpiJ8yXMw9uBEFuzHp84F9EtPwk87r3zrE
MhRTlvRg/zQURMO23UgxqUPBM0UMdGY4WyJsj3xC7G0Ogc9jdr0IaphaybAOGMbG
n2xKMGqgmxOv0eYgUfm3i4eyMoL89h5ZMOpUBQi1OWCHLgiy/PmSm3WW9B6cl/ta
ddkAkcBXPF2lLhCobHR+pfLFKIiHxhnNSfZZLacuKCNS7X6K+KY4oefQ1xwC7oqm
sl/R2j64hqjPqQDnFn3pDASHrG2LOEOknQ3GBUzA5zCNygc5qtzvu6dqrjJ67r3J
ur/tipq54Hj6pZryJf42o5H51+tfIQwkRFnowGdMYZwjLlKXH8ZrFMjkDs5NdJ2f
BorBjefWuJkdfc1CktcnKX3FS1EMDSLuu0KJ4lmpwMZrWRrv+AzhHTOBnCRsQDeo
qZrIVgvkBamt3Mk/b+bpmhDtBJN6BMeizMcbXD7Lo2Zo6vD2oGcWWU/dgnLKcnJw
X3mtfr6MKbu/dlrwrin1Yd+bmm/+cders3CkfWlST7oKQTa/q7og/lYyuhA+52ZE
19ujDMhk0sV++jaNdyodbqT7JRH8S+76bALeNHylYj3mWGDAV9oBiIGgXKomVsm0
icz1y+XfJDwYszPAVQgpwmkKT2tkNiBB5qpQI5KrV/bWp9H4kG4ZHumTzQhAEiHX
1PmEUqFnxKAc0/y4Fd0yMs31nBRv60nuuRX010D16+vYKvtjJcCyvouliJj68b+W
o+jEusY1AWOOwgTScxPCDZ57YK9oXKhWl6FraOP45EVYAeRFRbbczVNQ9GPxUKQC
Vl8sWKyLhsr3NnPw2my5LHtlQuTFNdvbOAIJvLMCDqL5Sk4nCGxH4ExwHg6FeqIy
LX01YwrqDqxhaIxYRDc+29w/EBVIWt7lv6I8hOAoybAiu+Xi9+YiLkbpBPUq0um2
TWx9LY4zjXShQTIVRHhkksZaGFCIDtjcyI2ZsuINBZfMfkG+RhkB5pKkmC+TDJDQ
31gg+uNcJksel8YpKhDi5f3TrfAMqaT7S4LPbiEMlUfnDBzFAzdoEqUxsavVJTKl
Fu52RQDGaU9lhpEFZDMDdeTUnkbwvs0UTbryK/LnQE96el24SkeKsh3YfJLsQD76
Z7lEVODpaaDlFmJLWs5bTbsQtFOsW2WQe+kLIVtbJc42PJBM3niIUOaRTFNbsp4i
UrUYlX6lfBroMN+o0IanuR358cdVprpOzfWubTPPZrquSR2RQ8h/UD1I7oCTdjxg
+3aeT4kqt9Fdzbm6RdcuPw4LDzIwAsUIz/fawZUvYXynUYV7POTME6PGo2Pd5nv5
3QmqXis3OTX0qyXJKTdOmBPDbSJtdkUCyXT8Lky5lC19I0uL2MU7H+Xx4Ywe/ELx
8DcD98OPByX095c+cx3IgzCHyz0tRq9SnTeI7z3FZ4oK7vYQY9KHiwxsSG17vNMs
vtqxJO6HfTnpU04BIV06OtTiYDx9GfN+e3CV76vSaBDUeLsKr6XzBkL6ikVj2zKL
6doOHV96a2GA1m5inlZK6j7rFph2Uur4AiRuaYD8nMD3DNnYTMEnfWwSFoV4qBOt
Z5BCXfszs3Pw9EDilo+FS/MYN9bcpPNck25cnQ9uK0oG+3l2jdB9nPLT8OG/t3bn
fSdaG8gDQW/D3XX2hNQSmybs63dSVziDsqOCL+WXokRuL9rQIqVTjq2csiGVR26O
NZ0gQa5ED2KRq7O6tbqIM6q8VGbxBBPazd1HCxzDAw0Tzwpr8CnAsN0X3dlJ1CzP
HWH39TqulDeKBYFW4oI+J5qwKYik87L0i6U+TTm4MTYIL2raGLnsygpExUhD9Wh7
dqjzR4gWMay2qwLq+fznunZdwIqO4VHzo8KAONuf578P9159JPQMsZG9eFnAY4vG
5TPq63IWupN4BNrjD75YJmtsD64eMC+M8vjfb0LCGL6FTl2zvS2PADcJNerl7gyH
d098Uu7NawlZ9qX6XIR4E6SKDnQ0UTVW1aNpkT+D5SrYrgp4JPG6tFd5bd1ibhpN
4tzAEUpcS1fhaOJ6KgcZ4lr+ZRDDXwoeZgcf9lvMlYjQuX4J2RC3LFNuzlEAURhT
GMDAQLIB0qAlg/Zm5LsYP/ROId8vF/UP6fb7rhHAdwQCU2EAB9Zlq93ZLFmyigJs
u0CpmmKdRgmVK7ihaVhSp6YtR47wRvzaM5Okn0/0GMyEuT5wH50fBf1gYNBzjFog
r7KpRA+P9KNrYuGXQgVRXD0qBrhe6rSQmHQfYznRkmsBmNlXlf++CGGeRAOXdq5K
VH9EA2lDcEot6MNx2pRCBbqFSbBMp45YpLLZnP6JAfhDaBqonCRv1JF+x2yF7+Hy
qAs++cv8tSPCRxy/Ji3r3YuBhjbxZOMuw6vhg9W8qO+PtRWFringYOIa5HKeY/ZE
vLqrmp3cxssezWaQMCOJsWKBW50osjUGZGudzL4ALa2kTu4dTHg8HR+gur2dVO/r
edGC9wx1hPz3A0g4xxnO1EYRQrPnWYRDvqhP2xovRGo=
`protect END_PROTECTED
