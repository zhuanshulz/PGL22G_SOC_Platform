`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oxrQxY8ffFcZW4z77+neyiaeXgVO5lRmiqtG9zP/DY/sZdLlHhky1h471s98OQlN
NhwLN6ylNiw9W8Zp/Q8joNFWrVluHAOwdc0FShgxNQA05A9z4683arGFAKGHjg1S
2ykXASZk8ih7FA6EzPQlynmGj8kE2J4s3nXRb1LakBZcTa6FOQyzqXvBgI3YheW+
51w0moMhEz/ujudArGjb+fgWk1LHNk5vOgN2Kriy+gfHAADEYlXekmzH2d5k3l7y
2FGFfoP06Sw+uiaRjSbIeF8Y5ul7gAP6cIHCPL8aJr90yxZodcsbDK1GNtyZbDgt
HuIGNr5rK6YAbHxQdFHMOAOd4cQYIS33n6G9L9kRfHUZLSwtuPGAVeMH7HBp+ooQ
y+CLi5+3FyG5Kc5Tsc4geCDD4Cq1jO3XPq2xMjfPDrpFHcFhaZAYF7P68uIaBdwk
0B3ipk+L20DQ9BBYn5wkB6YptQ6A8MmqLh/1nT1eg9DKzO3ev1cv1cmPCJMV2c6t
VokiXofVoIT5jnBfcJ4rrXOifY8WvXtJrim/uMRznoKJHk0ba/ty2TO2yJH13Y6l
73ccYKNCiIacmUVaPuGFokzx4xQb3WPXjTrIj7F8gT5Z7e3qHP/ii+KNJN906/2f
sOvLqrPE3Cs05aL8TN5pS+U0UJ1y8q8o7HjIWHzljM8nJP7KrwCj/TV4nhM0A6XT
qxMCtIQP03I2tw2GNBSHLN4VepS/Hhphcjy7GWfqXlv+avh6SktAh1ZwHBG+trVc
BSFifWvVM0dd9PJhwcyknR1CJAMGouajhRNL2S0EuTreBdKcbgHYXzsUbTKllJsA
16LW4HY28a2SjQLv1QF6NSoPCBhlzS2qGtpBfwRBuBiiXH5l38y9GDtVJoX5nM6z
DKdk/GErHKPbysyqHNjAsI+F9L4VSyKazZSndAYXHX3utH83x3ltYJ3Gd8N1AaTI
94iuxO7Xmvyb8tQ7t5qWMYEJs1hkYB3HrU/0kp/rK4yiEVUe3ntIvHlLH1uz4PTu
wnPDTAx4Ep0/XD0F4Q5ya5W7vcvOUrgp1Jp5fR5+StrcTRG5DGYT33CHLzxmgtCR
Fyl1LYlH+PrjqWW1V/r8mKlRrr8jyswPqjxfh7YtFyS9WpNj8deHEs/YeH58SJZR
mwM6/DXPrgKC1/rzMKe3VxxGOtRWKuq1UUT775TgACRCBE3NIB/Zuix3bQms7kiE
LmSHWOFLywfps/03dlbRAPW7hXpELs9I3yt/rgs+d5pqg1iWjJK7reG5UDlIZJf2
lTKtONgJkXM/jrtwldoj3QpE8YE60lhFb10/Rg+OLP6kiufngHoR0se98tyzd6iU
Lp6czVC1yzjs2mm6COsHD2fX2T6ghZjJdY10dFL2nX9fDPTdkhehnfmepbRwEWcR
sxgx13utTRGzgUdNJ7x1ezeOyXwtk9Uo7FTIMk9J4DtwCXuNxPgBfDy4pMJFUJd6
KAquw5Og5WB3Zg5A81gjMy8K4nmjZu+hxDgMiCUsW8wp9LwF+pHQ7XhMiGKWymHt
3YzQBFHrcf0v74h9g38Bxw4SMnT3GxXz62cvb2hajjjYyFhXdLL32B+lTSgU5RFk
p1CXiXB3xZSrOPD262iglsQ0OuP2BtvI2g2SdUTa+9dMw8YnLH35xQIgJjFT2RgS
o3QoveTdsOaoZzVU2I9C92+he6aHD7rfPq/rlTWTQK9dkvQFy7uoOE3oaUbyWgqc
2Gd2inqwaEeReBID/NzDX7wTVbnh46n+2V6MaZ7V3c8+3OQwYi0xLAUZ7kKjlzGv
`protect END_PROTECTED
