`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J87oClCNRF7kzfkmBcXbqhas/s1+S6GtlUqBZSSFvHOD8yO8JJtrfifBoXczWicb
4goVafwKH+arGLXvzHnIqoF7jwENeLit7Kub7lilrVeix4g+6xQxT0TRmcTMwnoD
Qldeia6Ktqmni0BbhXgmB+X7DwRh5NY6as1D2CU2MlIOBOC9CQbBwgXBxHLhG94v
or3SIY7UnQX0H49kFLezLgOjgJEm/Z2k2xicSsAIg/emyOjxbEA4yYb0xxkAcu9E
MNJzrjvLgbAH3e25QKvUzZ3KUZpwZp29VLx4VN3YVzmq/G+NbcpyCgYwPoCJu5iT
xSskyW2YKO5eytrkgZLAo3U5kqbiIYGfvtmyzAVkXR8qcOeaf7R/By5Unl8Q6Mtg
BGlxNa3VHfMRcwE5cNghbGqM58VryRAaU/FLNDSK+jsac/zV2dy2ERFU35ki/I7/
RfIRyY0eQxpSDEzEWp49T6PPouqBlGNeKa2hIcVjZjYFJAtNMX6kiXXKk86wyoNw
/eLgDKGrsyQ5MH8wqSs5ww8NevCF+aiNTl3nMIIomy2rm2Ic0E2U9CL/uOmCIgLT
uebA+3DTnlWaOqcQbgDaAS6p1ivd8D9z2N++8tP+MVGWcnm8z+OrVDtgpn12W2s/
ok/cfAGLiENxY2z71SPBrIrl5n/7eGYVFSjoMMMd6Jy8ItuG5GIDzoLA+Z+pKGGA
nVDwLC7znqI6918++9d6dt7I9FWJMP1YTDYI3djxkt4koecBJ6hlEh2vCfTpN6qE
iKYIMRR/rouGWi14IaG1vpw2ULid1mNz2Z41RvLLMeBepejBqfkfxS0I53XeHg7f
`protect END_PROTECTED
