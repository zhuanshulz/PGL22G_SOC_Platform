`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a+kBb+djz2DshXu8FCdSD+STrNF4iMonH6axv8VFBqdC/XEiw+2JHeRVEZHK5KTr
5BIUz/nJKd44pRhTW38g8kq3FjoXR+GoCfajcg2pKPvUDDwFmX7zYik0QaBBBukU
jWpS//dUDcWc+Z4fsCrYdXqV7tUFMYl8TRZBPSDqpiUChAwDEMc4Y32/N3gjiW28
c/11iWha9Kdrg96DDt59HPz/K1MFahCwdlGogDUOXShwa36ZP0a8ZSXQQeJkIY+j
zOMaVd6hnfxjTc3DVGjPrdCs30OXSOOV1T5MKauVMyFnG6Y7YrzlNPGyKLGicJcV
MtWw47++N0bDlg03//ucfjBPP4FqG2FxuV0BpyuHLzBUXENXu757G+DpR0/0j15A
jcT1iRllgmcV3v+MN3xCtjsnTbeIWgMIFGE1z0lAvdSShtdIR0MpINyWH3PT/H9D
r9cSK+U+ZFzqC7L3EmPaM8GNcpKN233sZpr9jDSkD7qW4iG9g6zPELTTmyL36Fo8
2wsLCU3gK/ttIlLH1r57uMCFvtEW0y24nyrAZ0rRiYKc1U7LrmWc/nFaWM4mv2z3
fO8auHGsk6hIq6AcykHYXInMQQzs2xFrojnW2e+To6booxITZHoj0M/ibr16zW46
LQIBU7FNH2NJiFi7bmeMKgGZPCNCthK7evr7pFiakG24ZSVTOnW6Au4+NlzSFH11
HjF+UBw9iaTtdUOcJuw9XMEqbmV+CfYgblGHSVTRflB9Ml1IUbpr0GE/yS36TNTi
mQ5XvYQaqjjUpegABYbJDIi5LM6QdfjOg8Xque0w+XgCnhys+YglhmE4PMotXIiL
Gd3po0AqkbEJR9/VP/qq0CxjlKuGpEqVJ5ytlrcITlVZt5CEDdrpYd9Xzgva4FpF
Um4NECCiAxOlK8WQkJmk3zcaQF3qFVVfUshvJZWdOYw2Ija/4x7BYNH/po9mNPxi
/XmSTN+ovGfC08mB/7go7+SRtGd2AzdCrrS0RK0DOwQ9a2D/6TFN/gXD2Pv/tjpq
VT9uEpDBDU35kUiOHWdBkat1cibyZmuJiXCYZZo8s8rRKSORUuvlrdEKqqNLazF3
HCwDXRzkZRM6R6h0AgAhtGziWcGE49apfc5BAwXmjn/pyxN2dDSumZhjv9vn1pwU
+eQa9bkVi0lKmuG4/DrQinCJUC9gSbz99W9Vn6oum5iGgq/DXoONAyr8voG+pbus
cAgkQvH2XVbdA4AzTlwWUX1ckliQUsM+3n0iIu7jcXktcm99TCA0MSdgrwjRDkqr
kXdGqwwLhxoiqAdrApn1GaPlkMybTXqrBG5+gxMxdLUCeDWoFBq926zH1PX5NtOP
lV30T883bGJ72+OeEnaJehGxo2jzLtt5VD4+0zHz2V1xDFNaeBVKtBKDI3eE3cUn
+gfiIt1NBxdN3FqfxiFmG2ixepE6u4Y6v5kDqBZB6GBxlZyPagLjjCk3W+QucXnD
U/LFYwbyVV6xnMNUDGn0kNJrARghJ2EJ/93dlQzWRGfoUlXRteYocf8SlT4GGRXh
wcBZMYP+wV9p+NcIZRGGf4DD2oVKIyvmxwWWQokLQ0u2A4Cy6YuI6TLQEJurqiIC
AuC/cIiqhSVEa+n3Z1dczuRzRi0vx1YMQIqyU1pvIHDJ/ML0ZnPtPdz1kIcpic1j
0OgnojiBbR4dmdTsyIv6qSlVyOmENx953ePCL7VKUi1/4wBWUAu/yERDWHA5C3zC
X2k3CBdGfOu1SZ45l3Fgj9Db6IOmPpNBNZ0r86ASj2IXJqHtiMtoEb6erU/Ts4SW
6c6yFeH1BivMjd7yUDBV5wiK9WC/XhTv9zhTyHE/ukpiFlrHcZDC/ECo+t0JMvya
91dNe+8KTWO6Zv2DF0GO2IcA9qPXkmrJJDmCeeHh1jiKueVN9ZSAFIVMb4POJHH0
bPMhhczamqxoNjHNVaDtXoHFLHpqa4Mjpyn8l4/7RfWHHihgOU72JfF1sgeP0D4x
U2s1xzVK3Y9yzy7uowvaGo98mkjp8MaPg58OJGtRgsIufW3BykAXrcld//xRrtHw
8L6DDfm9HbcELl3kQLboSsTSWpBVDmhPAEfzRwCowXsUTa7HH/UA0ZZWbzhREzLz
IYSexPp/SpqD8mAyoifQRoQpp4HQFWIXz98tajNLypzrpFyX1cotRy07dkgGzo6t
xo2zIcLs1o29Ll5ajlj6ayr3QKHFB2KYb8BxHzDkHmIIhjR+aOQ0LGsZS2dfMHMM
1fGjDcVfbVPbAxBpXvQnjdpTIsuUnSg4T77H3+VsgB4sjuzEsaqBfAqMDqQMdAxX
JknJX8JqN8H8pL5mr4ZLMujvGRxdotTlpQPwLWnsK3zwAcwNqN0YKW/cnU8i+EX/
qbNM24IjaFN3DZBgyc4wjPwhlloJC/W77U8Xn8wGyZAoKixwbVAyzFU18D8NXdnp
rvuHD0mFMZBASVlh24tAtyGyZA/ccAJn3X3C/N+0HbDFBGPk05Uw5mufmdn7OFML
km7eUXhBIIRT32VkJQmxDpYopMILhu+k0U92cs0LpShcWIqAqs9geNG7haQOCUfM
M0kEALzhVeyHoPccKj3UnuSU3goy728jdo4MowsGwn68DHDiQwbu6NuQL/z57H3e
Vkzn0T3b3iqbx7eZGHxLd/ltls6wuawFzHZ2BlXLMsH8X6cEZIsvhefW4vAcZG2w
4kIjT5Q3m7F20ML0VFDlYAV2frj5dg6N3QQtBA80cmRpNOSrlLED+9nr1Ancmisv
NNKZQzQq/Cfz05COXzj9V0Phi4KvTKfnYSZSd49Zq2vl8JWbd9ppRZORU6q+StKA
gPuLl3Ivg/8zaunh1SFHU5DY5SUO2j81T7Arw8iW6JKM6mqFK9YZUtt2uk5iPVnS
fUjE/8AbGXEPix88JkbXpEPNzNFglNoiveJUU5QAC2LdmNDR1RJYg+Z5BMdzYK6Z
ktnGoKZA/pECcHenSc8v9g5JZThIyHSwZbQtSqPMG4ROenN0hKQgsn7EMh9lXU+L
NZ/TVOiydIbhQpzWFnodcK6CK2sXG1KZhLd9e965zrB8cpoaiSWDQur147xE6bIb
6pBuSqgTRhI87KL+itNKaVo0wep+pC/N6jERIhKaP9KprGeqtBW7iHfjQvWXQkM2
oZ7SyM9Sop67GnK6CJKSCFYFD2hn9rOAgWHKkxgb2KSJeRz4MNSPri9kpikJ5xDC
MhZjGNUwFyYq3Jtdm29Vvn7UMyLgU82qnuFwUnpwrTkQXbBM08OdfiQ2eCTLPkDS
jj9tabRUzGraXK/Sbd/vN9VXP1zWRraXZbHzqX9tRuQKZ36aV/TUzbyueZrS+Q+q
XEqwwVIKlPtr2I2G3QMfpUvWaRg61tgd0wWkVhwEaXnquRSi3bmxGmTG9JzpV2P0
qSKTSQaWiBOwtb7nv53tdAjPSMBRBPGUQZHR+m463Ru6TtUCOyyppU7IkB9WTJXy
6BCuCuFufPnhTr2uaIL2GvnuSxxmYK8b31rLB76mwU8wqSSJ9KGB9kkFwKH3tauP
QG4/ku6EdJn7w9yv2V79n+gQr/8AqiGJq0G3SfA5TIX97ZAhBAxwzS83UaB4OJMR
IV1CJ1w4Oov8lzCrj9Q4NFqYlyCOOyspJTZwBEFgerW14juwc0hftY8LWb8tR+6U
`protect END_PROTECTED
