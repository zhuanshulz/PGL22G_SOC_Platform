`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E6xPpXnOxNdTZ89d+ouzBT1uI3WmR42PPZgj63PVZSt4wovQLPBFuR+Ikg0MC5ul
DKnopF6ovwioxMlAMEv2Laicmk0EETH5J9IKtiacD59gGPuW7KgdBm+dtBXcO2cd
3/sD/L7DPIvmQcXRs/jYVWeI1vpC1NwsIluAOGUrmiguUtpXjkM9+YlrGA9AyinW
mEDIj+3PB3p5b7lk39nzLXngqJF3+Y4IX9TW/8AZPnju1MuI/5Ai/vdkSFW1ps1u
c16zq56EjHXX36RrP9kpZmzxA16UTxLIYhUCq1+oN0XG0TsCe0tKGkvtSb0eVwyA
6PWgCDqObACBFMwj2q6Qk/jQ1LHia8O92PaqcHh4yv+vLsVMY2RoqFQ9l6NuZdp3
r9Q8GI4Vuy7YIgznzLcis8iHkdIMOR28wqLpfR0JG6iMOAtDu5/oFgtMxiyc6rKU
FVENGrqAZ5I9GVUP3+v9Me8zXGaGKQVyE/w20RG2fb/OcBQGkxi/mbtaVb7tvNwX
+wQsZkZSCfdspRGk6lfUV+NXxVKzamoeIhJlVLoSSrM3wL+8HpmCv9ppyulT9+QL
q3lutSbZLjwzt8HXU+cl7Cl1Q3w9VWXiIMK+4Xv3dQtvWnT8UOTZZy9tMBzISDZp
dKVWu9IromPjtesnMMyORgCDW7Xg6wxtQ6jKeVxSZ5qhYbj09xOuqMVfK6JBIWhT
HdNLJdhhswREp0xCEHqUd+5x/sTdCJH4K4lXY8cyXCiKd0+Am1aSPd+CeQwajJhJ
9sUnRRFfl15IipVCsgeqktH/LwVLuZEkhEcrFR6CTKbBeZyXOrkAGduicU1eDE3A
T1sFYiUFnVCje6IHOrioK8UYb2noIcojOrgy7luTnbkCCu31x9b5Olv6kApG8/5K
cDaTuFYQRZQyZA6ggjFev0ljtrUqHgrQYowBwX6RBtV/uCxOBgb01J7Ee+Uc1qXO
+eUJBxoff1iIwvheQWsYQ0nCc4adI7sibMXR3iMyuVudI2gsUHjmXG+06NqQgDmD
Ph4rSLNdzeDrWxYucX/9G1gHHxz+0QcN/T4KkNlPMavH+b57r0lJf8KLfT0cUzGg
b+qQ3vTGeDkzZCY2u4zJ7T0UMs8E/cSAQ183u+qjoz8LZ6FL6iGXyraE9xANtGp+
TsfI30vbxepVH1irSzyESDbfNhMTiECD5vCOt5KINgdUiWwP1jCEKebB5Kz6ZOqj
Y26tUASod1UWZQL/JlAnrQikKgupqqqVu5T5rhPSB8NR/K/DC2XPBnEePz5xN5Tf
OaXH/ktJcqgoDFscPf5UvuqIkJwc/8f/yO/Qcaopu9eReznLGeFlQ1xNRhAFxvUi
v6aohG5r1BiUIb+GyeNND9ldxUQMYnUP8I39LGygYfjpDjyI9Ls0m/3e7O/qqFyf
xUcnjNX6jy/QVOPCabJhgB5FCXkMauVx3bZ+A1meTX0nGvvODYGnmmvY1LwQonWT
Z6eUX/f/JFZ9v5IwPYzUQog/61Uo6SPq2mvwjgDxSI+G6CuYdb70voEjN647Qjxs
uUqKRGEz0QElcChQfQ0PWH3OiKgA87YqykOwMvtuGA4=
`protect END_PROTECTED
