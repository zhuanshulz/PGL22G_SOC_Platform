`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cNAXNJsN4bje714LfHOp2bZGP7TcAyb8iFN552XnwGLpB7h8QPfzoeCsUaaIGwzZ
ve075+j6MRcZEJ75fzAmwFPPtloH+HUY8fCznQ6D6IBYEhcoXFDnsuDVRJEFMNOO
FaSUsiGSPN0xOkAOdm/WtF4suCeL0wTDeQtnY0KMlX04NyDOuIGrV4lX2YSlyL/S
vdc5sX02CAvvDLEQS9uhIM6sj7gOwqRHFfqZJ+3Dwq1Gc3VjJCdWAsU6xKTIZtFR
z3pYv4u5Xd40gLrs8Ukoogett14YF0n4/ti8gggbi5ALVC861yW31d83cFEGZc/2
NTshJJDzLsewZz9EsCJppV5HJrZQAOoy75BuVWpkjF1zkb6d9cYJtdwux4yyb18e
b6JS1/LUJlZxR2iHFSrzky3gJ8yTrnqqtpBHvZzlre3rHV1iL4xOqHtITwgu766o
wcUY/zY2PmhiMRMWgKjJGDN74VGnRb5gL3byibnWqQOb/c1ViJWtpeC0PPhVS/dJ
B5u1vics10TdiqZuHYxBFzRujOkOf0ohVt7O12ZGxi4yCpiRszw+o4CPD60KQug7
slwWWshXBmZltsgTWiBJOzK7i1RwLM20DYxZW5JjLGV00MgB+Rl1ZgIaICdLvBYW
xGlIMt/DXhHRUYR7Ky+BfxlOaSvj7MXiG7/QxMtdGARTix1nfYbxHEkA8J62K0jN
h2TfQoLu0+HCpyl3WgQobj0tASh8op1IEwvIkMDdag91eyaeOwcHG5yceNUuwwmB
mpGhryLg7OkG3FrABrA51k7Vd3Jwo49gXhfH05M8SlaoxAyQqyPbI1Dvbdg7xMCi
vpgIHnUA9XkLoepjRSBnKKfdrGfUFv6N4pjVY+34Lsyg4F/AaQwpsN1khC9xg0Eo
EKRRysn7QP4+glTH9nSddNzzUNxlqgl6ywoYUKwQAf9hTxVjMBJq+9qrRkXX3uIj
iJzK3ujpUe8y25dubek6V1B8rmTDfURr0q7cZOP8PsevF35mgIqTr3d2gq8XbNt/
wYzDXHVUx4hw1vShTlg0OPeyDZfmqXox+n/YMXiCKcqcZ2QFlh4EIx6kkilWKf4T
sQVKdPk/gg8i1ZjYuoLxhZmq51CVTBZwPyxa5jPPxdBmk6Ydl+a1LRlwMinMJFEX
Rrl5fnQddIruWdGKZWqj471cQOUEyNBE1mdUuAc0X3YlXfx5saas21I2LvrXYYbS
hPba0XniTaK2rjVg7RZJsu2/460yVnXe9Y5dhI/i8Z28uqNoXpMKt3PrZhUDJ23Z
re+GEh9f6mCsN/kws1n3DOxw3LAC54miitdHEXRmNXzNsrenrX8iV097JZs8V1sX
ceHYLIkt4LW49X6G5Npy5fnJf5UeyFyvplwAr4GUy0y+onpOw40TpY23ytZSQA7W
1nYdecE68Is6Rf24UHATHYeHur4jpyqyziwctm2nTqg=
`protect END_PROTECTED
