library verilog;
use verilog.vl_types.all;
entity INT_PREADD_MULTACC is
    generic(
        GRS_EN          : string  := "FALSE";
        SYNC_RST        : string  := "FALSE";
        INREG_EN        : string  := "FALSE";
        PREREG_EN       : string  := "FALSE";
        PIPEREG_EN      : string  := "FALSE";
        ACCUMADDSUB_OP  : integer := 0;
        DYN_OP_SEL      : integer := 1;
        ASIZE           : integer := 9;
        BSIZE           : integer := 8;
        PSIZE           : integer := 32;
        MASK            : vl_logic_vector;
        DYN_ACC_INIT    : integer := 0;
        ACC_INIT_VALUE  : vl_logic_vector;
        SC_PSE_A        : vl_logic_vector;
        SC_PSE_B        : vl_logic_vector;
        SC_PSE_C        : vl_logic_vector;
        PREADD_EN       : integer := 1
    );
    port(
        CE              : in     vl_logic;
        RST             : in     vl_logic;
        CLK             : in     vl_logic;
        A               : in     vl_logic_vector;
        B               : in     vl_logic_vector;
        A_SIGNED        : in     vl_logic;
        B_SIGNED        : in     vl_logic;
        C_SIGNED        : in     vl_logic;
        C               : in     vl_logic_vector;
        PREADDSUB       : in     vl_logic;
        ACCUM_INIT      : in     vl_logic_vector;
        ACCUMADDSUB     : in     vl_logic;
        RELOAD          : in     vl_logic;
        P               : out    vl_logic_vector;
        OVER            : out    vl_logic;
        UNDER           : out    vl_logic;
        R               : out    vl_logic_vector
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of GRS_EN : constant is 1;
    attribute mti_svvh_generic_type of SYNC_RST : constant is 1;
    attribute mti_svvh_generic_type of INREG_EN : constant is 1;
    attribute mti_svvh_generic_type of PREREG_EN : constant is 1;
    attribute mti_svvh_generic_type of PIPEREG_EN : constant is 1;
    attribute mti_svvh_generic_type of ACCUMADDSUB_OP : constant is 1;
    attribute mti_svvh_generic_type of DYN_OP_SEL : constant is 1;
    attribute mti_svvh_generic_type of ASIZE : constant is 2;
    attribute mti_svvh_generic_type of BSIZE : constant is 2;
    attribute mti_svvh_generic_type of PSIZE : constant is 2;
    attribute mti_svvh_generic_type of MASK : constant is 4;
    attribute mti_svvh_generic_type of DYN_ACC_INIT : constant is 1;
    attribute mti_svvh_generic_type of ACC_INIT_VALUE : constant is 4;
    attribute mti_svvh_generic_type of SC_PSE_A : constant is 4;
    attribute mti_svvh_generic_type of SC_PSE_B : constant is 4;
    attribute mti_svvh_generic_type of SC_PSE_C : constant is 4;
    attribute mti_svvh_generic_type of PREADD_EN : constant is 2;
end INT_PREADD_MULTACC;
