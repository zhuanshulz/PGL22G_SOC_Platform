`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LPmyBKc/P7GYSMInzK/PyVqhfgkFrnymA0pi/MIPRN5TB8KIbCYjwQKpSQMobrTU
PXT3t+Y6eT7o3LjbGtrVg85esinFCXDFfhlxlGKRkOESuG4eDdLNLzb8ghROax15
aYuW1PDZtEfyE1p3pHJzT+ThtfVM40tu5qKQUd6iDrgSy3rpgH/IsA02fdomVcHG
IdZ38cXJNwEVVR3ZDjgovF+DPqNDm7b2j4dBkWmMKTsf8JRTeoV2x9IkAucetrxX
+vTfIgzHBKSivmaI/gI6bVGijZ/nuyeUp4LYb0BR63D1M66JRQXZgyKtx5K5nYn6
/p8Q0JAllwbWmbgFyGvaUzJGzD/h7McmR/6S3I4EnZJLxj8Vt0Mvgv2/D4g23z47
03SUb9medtIz7xua6fEPoNDaqwG6rrpFBChNO7bLWywUvqIvJdJ6pSumuuUvM5+W
`protect END_PROTECTED
