`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pVCG71NHzMXjcUAkKZZ1S1d5wimDtvpRS34yacO6Jq0xgHyG1+h9wsrlcwxij5UH
puJXwcLckVI+I8sB7vN5EwHKX6eG2gRiYHO8wnc7OHvatzym3/FB7ea4Kcp2lPvI
t06Qb3xm+UzCdHyC+sokyh7u6NDlYJJ540vtzIKv1LCEzpLAUQGMV2kX2XHJforL
VY4dU0jUOK+qmkkxClegvKELZyDXXNCTlN5mUZN1Aygj1cTHlTicwz3bidV8Zx5x
1hQm9INZN39Y6shYXU3WSEqMZW1N7Ux4mhrW7aXJyIjuv24eOOFvQXNjTyGk+d0u
251oBQyiXrA2sayRudaaiCwSIEa/pkLjmNYCq82z87L/dRRyoZ+RW/O/LiINkCUe
fgP4vBeJFiIA+RgiDNieTKaxH15Z0MCh+Xeuye/K8ft2WN/g3WZrvBWNqZyzZ7hu
H7QW+uMT5T2/G2KcEMxKaWS2WX6xYEO7Xm9ORzqgMXaW5PsTXcaqqGAqr4m6PD+E
2SWbBG8oW6Kc6mbNfdfpkyAGAGr/Mf4sX5LsweukPl/xSbYKSJFlLNZiyHo+aVNx
zOxtra1yF7n5199W7fda8mtQu/XofAMFazn7Le2IwohM0uFdSCbbjzbRODUgJDvR
R7NC1HxKKlSYX1o1xrVACO6v76QREeu/VgJ9sc0LVqfpRiCbWnlyx8KgdsS/qwWo
ciuGxm8GIm7YJ+E4yMHKFFKPalqYc4dPEdhMjnRE1PANfWYAF68PoIblNbtDM+rz
uUmx98KLhlFkczbgR+cDlYwtDnl/A3Io/RC9ypEquxwuQ9BSPRrgT0Rg2XtFkp2b
/sYnz0BTBB+KBJnVYwHn6cOazcoF1nU+8i3yvUdgIGh223sSRaRhB9V6nhRdvbbb
glc6Jr3Oj24X8580JeWwSBSMTCnPmNSDoobSUhBdvl2fUD9ZiXGCTzQDCu3MS2wS
/VogJhNNdlEXu9DqTK0FbErX5+W7Urtknli2q2Np8y4VgEBeVyZpcyQWoOidvRx8
fGtjnuzeqUgcTZr4vm9UG62hWQOx7hYRgcUVy5Vke4Z1F6O8KamVF3E0loL0eeem
X/jdr/kK6KOYMntDfruakacJHZt5NceGHOLN4hiyZU0KgGu8uf4KikUcsmwkRwbg
oTMV4A12auaVIGbENS3xUsJYNwAlzVtWaGyNIqaTjiw2bAwgQxLCKltk+HxuorYo
sPNbmBOcpcX5A1QDmNSo7vqnkq+/fawH7k04F3l4Ls+G5RHzfNq2GJRLL6Je00Mr
Kkbv2/ayjxWsjhowQVvuZozTSqRBd7gMvPnkFEmG8ZHrIfQBpYOQLuWyqzdcnnGF
COdDKWbiOGrx3VLQRptkfmaRpthgI6mIP2t4TzvMODlZAvqOaJlF+kSgSyzQEHRu
aevCCBIHrHjoDCGl52Fi2NsiMtv5nokhf9u82vzmpvqeM7UXOYtZcjz+wIbIT2DR
xmzo9MLLbCVStdwfwZrMyNhFjLTQQkAI7EOLipVmrAggrpzjXnLkmaeGRcOpVxIX
aEp1/xFN9SHorwUYJQUIrjeA/yYLyMdqOVgH6g31f7p2h+y9pFBkgqatSZcRTeY/
sKWJVLB+eKL9XxzFMIGlEiaUNVm/6BMHLWCjOyuhbde0OJz4NxjXnXlZI0gnBwYP
38GhfpF89Y1CPIyUFtyU54FLtaORU9szJ56lc5lUaLLr0zGJq8TUBX6LUzmTYyC7
cSJURt02CUxBz7+82rfFZd4sUhIdDId7k1SUX25qDyy1k0mLiqDk+yVafnRezDdK
oVcR5gfgd+/OzNg8NXHkz5P36micAVQzRXTsPotZ3inLDo6jhiByIN6h36w/p7Oq
EmSWmIpJRoSmj4ksxrSuEUL3UmTgVJnt3/A3xPy28/h/jZHxC6X0qPDRm3XyoWv4
UI2wptiwqrJBtscrt/qYKwvEFT8OMaaxWKcOStuNh1w=
`protect END_PROTECTED
