`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PKv95VEKb14s2Op1WEmcf4QKcYZht8jY3bWs9aPuGCaVZVi9NUIv5UrNsZvEFY6m
V4GfHR9d8TKq/pQL7pEvYzJDvzllpiW+msSlgavpARp7Mu785zlu590irXF0DAUE
7tSp+XoCWlMJ1TZzzCxUcMYrYRTI4cLt+Ka3tnL9nJMaRwitHCPCxa8tL/34Acce
EkTS4+5JRrje25gcGR6KYyke60GQ1aAQ7ApNJ201G/Y0/zP7ZQIlDAc7jujhCGNJ
WQgF0zKSOqmCeQiikQwG7+hGc1dojV135RjZctSOgai7Mo6EZZV935XU0ETZuuN5
CedjbCKMtNpEGQCuubdUh9PGUZUAcwntmPy/AmLTLLunCf4LNqIK7bVbuJWwhm97
7skn2dF5hsENDQ4L7tVcNY9iTenlp6IjKqUOj125elRkMneKiJhdzjcjSvvYGPIr
Vi48sBN/61ntYIbuwmVKnLaD2xqCImuELEhXMGrxCywoKnvUMf2+hz+8OdIVMI54
5+w905324t+wIb/SQOTiiwUQEmHZgI1w+DzgMBtAH/4ZreBekb5QEnSe7hILANho
MgVKeXPzPbhGZWZJxQz4qq+N5VjhF7914+bpZyQRQ2pSKPeuOCKkNvGa/ACDmigY
dqn4bn+QzHBH4GJAqR9VnPif9HHhxIuRBczUPQNRcliQtK1n9QpMtEm22P2N3uGR
1QzvIvQkgl3QSz8YGx0dj8PBWQQmgKMHtV6H/IuHGMisYQRHxkB/0moMMWT1e/iw
VVLUXw/FaSN6MS5a8cR/4GggW0xmuENF4cTsfbh7O9gprRCG9jYDx5kCqWJrV8F/
jVP3Yi0/E16GDqywRYh9CRHo1h7KhzxB3poxxQmDWbWMYjrcw+MDB3GNnk6JLyNv
4RI7K35ZHivjRUpYYnh9uJSmr1upKjt14wLi9yoQMtD6yTK53xQiXTEvANsNRJJB
RjtL7lMjbRexLb/lG95eK0ZFtEPm4+897oDdNgN90Mu5MTPJ+mW6JxpoATu8tuFM
xADiPpt5s+D4g36jPw9wd3XtKuxS93HPbfbuighkpF8m5gNN6oCfZ3mJG8TEngxk
zZLldV7E4yJsWsVgbRR3WBrtduy3VBsmyWOB8utqNctf91mPsf2gtinxuHLQjX8p
YvQGVQnKmoqrSa1728MYJiIdzBJ+nj7D2Aq2QYKYavxxWpnJ09PTxlX3AN7STR6C
WJk0tgm7FFHEjV3DUAN5sumQdx/IUFXx8xqHO8dCzxplNzvHESOeAahAulnai4b9
KEenLf+aCtofsUr6MUaY0vLX8S+MAcPPoe6jVl/Fx1tZnA/nO5c7KgrpZnQv+K87
UeiM836P4TrI9AJEyNglZjQ8wcWCNkiN6ok0L6zrMi4wQS++Wt11C/fK9nKpAGKy
tOs35L9QDdi92tM/RmYG5+dK0hYcsZ3mE4aDyJdIbnDPqmR/XyAPpOYcwnScMeZD
zIDNTolWqSe1qVPzCISa7nnrYmIpPYN/NBGnu0efZC9jdxFFWm5NvMls8Dvk4xHy
gwhZ0JiyYABs8XT+dD5VditKS5yikpq6gB9N6H5vX/U+p8qEDR8g0aEmaKxBYTsu
49SYBDduRTBAn3PF2/GCF5t5TFMljv4yjREO01Lwg/6BGFvXKyGWji7m6bok9I84
AglRp3kx/dY7G0wsij5p8UHln2nE4438LRm0P4gaSJ/MWLvNTsdWEW2AmC0NjHOy
QuLnHKWWGLJxaGzdfLMqlYmf4YdNQ9t8TIpFJnz7P1EDAz/O12fwO+8RoyrnY0DI
jfjPpOJCjr0bjQTiKxiiIWoQVrNL5+vKmpX4LlZZnQixQms4duzWOWiFB5yzXWvH
Rog5VrpWO79gU9Xd6wF2q5bQxakbGjEZyZ/qKldA5t5m32F23UbNNDUILTIfCyQX
+NfeYibM/akNcB+7GcbmDQ==
`protect END_PROTECTED
