`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0wzFe6mZFAcOFpSq07gt7ONlYXQqH+AXVQOCDXDgucb9LPK2yAX5gsj1Hy1faVGq
/LXOgxDA0iCQ0/Nzmah/eUOj06c8c0cD2G8Zh5d8c+k16MP89m4pdqVAXaspjR2f
eR3IUeFGm7D6yicuCMWN0DjOwqfvjv59eRoarIaEg2ZF/NHP9hrhflxoYv5+fGlk
RWpe/5L/YCiJ2liwLUIzYNdjGYlXM0Qb/wj3+HBUkg0ZHV2UpJ1eazO4kNyHQ5Wg
+DhjNha9cMLxFvZynNBsVp9h8pwj/hLfTAEQcqroGFYHJqF3JmMPY9vPOedexi6e
AJeUzc+TYRzQcWilIpS6E6UlCxw1ThRtjzvCilR7OBrmJI0HDY8RvWWdlsOK6kKL
sAJOr9939fBEROvWCqHb1bKUP5fpxarjyMj6DiOaM7w8zS2BrQCLrXKnwJPXyUVE
4xS1M4l4d6LQfvEVzqJd+rs14hy7FoTx+BN3OwHjelBFuoDKXfiDmo7vPrJnwTVW
8xisPfz7Q4fVmVdDjg1/DfNdk5fEZK0HyQjGpTXVkmyB//3OCb/BnJLJ/wW/mWAp
NAxtIoD1Ge0k7dPW+C6ERojUJBpcHSsCZ4xdGd8gzIG9/gfDqAi6v6PT46Rt0ivc
iyWgiddtfCUnHJFGZ25umlMeUHxUGQe6rJILo8//J7I=
`protect END_PROTECTED
