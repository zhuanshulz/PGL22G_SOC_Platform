`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9w/tY+Nyr49CZW/FEllkXRCAAPkknWAJysx3XktSWN1a81ArkwoZdzcGZeC2RKnn
gYHO1t8SbqANvZNuftrcKvszYKtYWkihRzhvlPXJfdLC2OmjnM62h79B+bOXuNRS
RDrL/0PcnWT6pa5e2fVRNjkEPsT/X/OfsVOH22KN51RlVgXxb1EMRAe9e59Nwcd2
S/9yZ2tcgPju5u9yC5DCJAzdZLa/aL1nPQbTDa6FJoL3z6UCA5XUG7ORv1Z0ThQ8
JJz9sLukWfHMQDnEQUPJk2MUB00Gx9sBURnAK+fpCUff9kd6ulKkhwE2FNOJyqhK
ybUi5mXfXXmkS7wMOgoXRMJAYeTsfE1jAB1Ln8Xy45ObcMOFG+P59D9TOHBXO2Kx
KHbT4BOTwsBbJ5dATmDsbAq3WzPcmE612yNWMrVuWfr+o9tRXR89uM8vnFPptEde
`protect END_PROTECTED
