`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WQYrcLihyamUpNG+cE1HWvhqbiLJ9ATYHu+B7c2fk8GOLhtiv7WSVkLDN3DH/OS/
XQuWyklkfJmPM4OSK3MKqJarwg74mSITPCIzq8Udp+3l9BxDiDDTID13gAH4wy/l
klxuVAPB0hWxuup//S4rOzx8uLc1r197q0lpQY5JksNCZOVjjhdgJ5ujfkZAPIzc
9yqEzeORH3QLu5BiUBozStFTS4JnAFPnMbw1UgJtoVK20Y/9PwLG1qDicOYBSv+g
5JIAEQuLlHRcbUeF4ZaiE5yl0PXCLhdBW8FWt4A3Jic1UnPoRWgT9l3gtpBeXOwl
inTUWHKIxy5gNPhDDRNnV6dstwdusAA8bKrhFatAjsavGKphd+v8j8NR9BiBv12U
71skgI1fYHRZCLEcR1IwHffrv3YA4ApHMxZmYUm9OWLT5ZQOfNdzvW/nokUM150B
dVcsLfUeFrmGWLxJfcLEcMParRQH24n37A9t6c18NT++v8oggorF4AN0cZ1XmiBo
GyewfI60be+4hy4ESSAjh0h8tbfRza8J7flTo5pECbBs+ly36YQjckWmIOVgYVAH
H3pYg++cMaGMS6bA+QdO4pUe2L8iMliza9CWW06wLmKPsqIJv32TIjWYwpHgh7LP
jJrVz/vVW6Fz+3PdFwUOhlhVEo80JdEChCGsoda8yA0sWQLEIHSowPBGtCDqrb8W
fqPVJcsuMogymqIZFYSfnTgeyJYMDdVlFgCMqei4Ev8iHJkEB6CnUigNcbe7igJQ
x1IPpKYpPW59eQbx1EiQOZGPzqFbMRYNKkE4ffqFu1MzslgMxEYr2oRnL2KkvZGf
H/0UtIZzUw0wcXtY3pC6vBqZKsmbY9UiqjZKediWmnQtXs+t+HNqyP69Ikn1kzQf
vmTMCchuWHTVWkZuH83qtIat3Vyk/zAuawbQHo7wJGhCHurelkckjGq4xHMDXGuz
RqD4Ry6bqcBba0gQj67QU9ilMQgJHYmJt3PdJVXM26tXJuf81WclTXUkCCoq/BFg
U3QEGe7ekJ+RR5xZ+v4LwCNtZBa3WP4OkchVytnDnQk9AUeBXfL1fjpNUkS1MhEe
KzrXeXuPmGlGYky2nFIK+QHPE5bbr90dJfs4C7yR04o6zQ+ORorqUZ3wlYPldJVH
Qz1Xxc/G76J2NAsIXvCsUT9X5qlX2gZGGUaTTbgtk6hOePUhUdALbcoBWej5TwKT
kvM0GyDutvrNzCJrEVfpAjgnKVrCgWpPuxUHM0q0OiqxDoOcWfIHHJRWOD8ekInP
HIs6mRcVw0CmYkqE1xTTMOlMDlPhCaT9bASa/JmhfzSUQZ9XATJrPpbDaWm6Z1pG
VqdEHUm5sq2Vj//y2KwEkq8WnSfoPpSHVp1UN6cf58z0U8M/7nbxBm190Ca3hPCm
Di8M+KsWYfWvIs1i3dyIhdLxFMmfJmxp9QAqPIgM/B0TVdzpNeZ2pC6+ekmsgGQV
AgkzXwwibm3tBCaje58WaYQndHbb8107ZPVF1jlq6DuC9bo+ykM3A+zYLaoWiiz0
sAnuUKqrLNAPD/hxpsLB7ntCFwesGAMVPy2ZIyvCIv0yeM5xvGv9mMoW78wDSwgB
14p1B5N7M6weIEKoo1Y2iH/f4xsiV1dgmasfX8H833ySBeqUR/h+h1ksQ/9Vcg6D
tAdqHGB63QOdO442gxa6QiF32Eu3KUJSwExv9bE9pvbkf21nnXA5UQZXOl+wk9Dl
ywP5GP2+Xz2fVhIReSPotxC+ann0Nx85AjG8X78JeR6P+QgprJpCidpx0VQb0Toy
DC9goiGh3ZTQjHRt+QvrQlV6llPPjuAZYFdedv9P8bS9mM3Md41hkBrgGv5EMfVA
LDJ2QpqMcrEjZuchGDvcIjXCnQMlTzF+Vb6PDfHg2oATQkIqPKHrGJXk4SXHzrnZ
z6MaPQA1eN/WodotrIahgsK77e/0h9IHxDzYL268OuVw8Y5lMhioGHDme0Da33Yw
U5FmMFcZ8BCpI/+cK8RCptG4y8fIuXLgMFDbqlY9gN2c958OvcyyDAEddkGr4H+I
Qj6/yjzkfRvucYkFJVkJ9oYXg+wHWxh/7MeAmuzwxPSfVqU1U4ohMc9vPlaT7W8q
l9Jta1zOCPAGPm045RkPXH0kpejhvFHXZM0BiHBY+/zTikA9y07icRR1OA9aZE9z
AUEptv7toa/1YlLwAqax0rx9q9wlpokI4P0Y82eX1Sgmq3cYg0jzUhkoitzZhdN3
+Hy+77NRJFBc5D+KifqD+183pTiEnfYUAdtZMcGgAzpK/tViYj2Gbzx6JeNBkDoK
Nrk9u6GEPYtyOQAIHQBfwwzZ6EFmoV24OvWg7qcT0vUOnt1aFh/oihwQBmKzuF3R
q20cNfogWSe6cCpbWSeD5SiFxDlaCST5/nk/71PBsFD7zzgjhzVKfU1XOdV/18xo
Ft3bavmNbWMJEdSgR4dA72WkZXOcajgOqIeloYXzobM8t3tJzJSPLa5/5OWP+BHP
8wKwOCYt+DewENIutE+kteIr9EXl/XxPHvGdU/PXR8jqz61li6RrtfVX99XYgmRW
8AEJFIruMwOcxHVQ3MGiFWnc5Q6Nf9++0LphvI01LbdqiD/1I6+SgG9BpuS2GMeA
2m27GkiNwE9BftgQyW1hzHVq3yvmZFrGZSlIUKzSRDI1zjA2IBDlCfuI2EI7wijJ
UAG7Nh5w9+3cIR0eOIbbakwkZHNuvpo05+mmCjnMmF9SV53XQpWjtrDPhJMWF2Ee
hXLXMnCALT49+PgWwZ599EN6S9NO7dCftGFg0cSODTiNBORbF5GEU7r8VNEgOkcd
ElDzgGgN5JVFqm7L0x0mYoHKgUqjZyoeZOWg4BbuFaAe+ZbOimDQq4h2D1ZXkh35
bzDw1sWCcxRZO9QNzQYMClRmUcQoaXoEMlNITYeuGtnSJLq+H3OL3nzhndLXOT6E
/wJrYqwzYE9NUVw/DUjjo4J4sDgS2Spypo0aPwf7+3w0WMYpHbbeuZvW43zjFpsX
hW9i2usqPdts58nf8vH9UvKkNvE7Zer/VsgoeZjmI1QuLmwW6vmKIXotznHMk3cf
ItnTyfxqYBBNgs/1Q2oXWT+oKWlzph7oW3f8ZNcfdLFICoP0WErMkjvdmjwhDABr
dx9YfHjkjNUACvxKn6kaKtIGY8w6DshCYX+UdE7XtOKPnGXy1NylDrhQ7PqKvJqH
c8ihI07/dukshW0+W6/8GTuJOBwmLMuoYmIrEIhZmSnObwP/7c6ARs+u9h2aLTZA
fluWpWv+mhcsGDY1MgSX+jhtZ9LqUUbyjqNrVwailvOwwuNPXURmdOVyaX+VJ0h3
TlnZHZ3Bovt/3AiFbPuqXfL6mdFmOYJZHrXxBdJeZYhCyvtzpT8tNqCQaFEq7MZr
XKBf6r3CeIj0rIjC1LCGTmJ3vljX09ZN1+LvrlhRiR4VSKuNRD58PTjgkk8+UBBT
/3bmzILz1e5MhweNSvVIBhujm5Ys4ts5EzXivbmm2Vg=
`protect END_PROTECTED
