`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kGfamSFRUVZsQzWll5BTDH185NMG02sobrW9S5Bb3KAY1saum+Jadxl7C8l2E0Qw
GfAokwrsTd4WJ4hypIs+aRfDsbzhBNlYEL5RgXQ+WCZ+cmV1bR+couOJ4gTgMZlb
WQypczzmE6s66If6nvhZa3VkcEUgk6ZARzgjXJuoxL43xlkFOiKhnnIQW4HNdJBJ
cTHTt0KUEwOaRHiAhr9D9Amcr9DNM/8aI0y77OgDVT9mfaczQJ6bap3qAH+as+8g
8OxLJiYaAPv+g4RQqqkwYfW/9ZGDoxj0wkQTAftoVr+9wRnjEq/cHJPF8oKFqCp6
1dJBHOVis2BtcMgyIzNQvjpSJ0LctB0/YrgFpjAIw2iTMBbOZDk2z0PoA9M2LZmS
X3gID/x7MoHgcHxXKmr6leNj+savbsjM9zScuk669pqvggYh6soT3gUvN6LdN1iw
p3nUX6KoiGAEQlTRZ7M8duMGM7InGoqpLMf5RSTB3em7torAuBzNER40OwsnFpVk
ZzyMSR2gzpD5vPoij7c+CVcdqHKpu58/Nt7LB8auKDu6x3KIC7AhF1sae+3lmMdZ
DKV+W990R0ecg0pPF3Qx+nMVY4fVrVmKQXquADl9d7IYW64gTafWvIYTbbochigE
sZuiKAdRdyFKJADg+TEcev1AWJvVwEe91aP0LC5kgnfLXUsQxD9dxFxJkTaCVTwz
Xw2QS+uCCYEagbAxKutk5JHuSsZjihl4xp/SmQaz10cRnrQo62YciH8ZWV8YfdlJ
YCC977b2p4eUqnblLXa7GgETq9SqvC70wjP96FxLrnkZ7NU+8SJsVNoY38Rb2B9K
UArnCxf8ZUkgyVzKVPdkVImyuPqDUJMGuFqIsjVgn36CXBZPxIvTMRSOOzvSU549
g3blQtgHRenKiatGrs7c2sOcdpwAIoy5nh4hEHGNdYU/rAaVQcTOAao8elV3Wtkd
339va4MhC06+KXzjTECNHiHSKylN/L8e/Z8gzDbuXc9Ms//W1rKXt7qebasuW2F8
mgxFDbP632+Q0go8QM1q0WXSUCbzm7rGZh2wMhlTerFvWQkXCJdKpqc9JXERTWCt
Jn1Qt5uxffFYa6crCFeeXz4OF762slxZtRXCkytmN1I2ORBAysoDo61X5w9iqsqW
vlMUg+YLli96Kaw2SeiAJWY4EBvqbdUr48NS0pS0mTbvQpnvQot+jYiA1Dj/KwhZ
th4146A1sOrlYQGxsIOCgyZMfpg+l91fqc+HL0gYsuMiXLpXjOWnXkMXXQtYijDz
x+6avgxEgYixul/m4G/GuwWxfgDscdEksV4KtYFptMM7YJTrdzkP1DSZmog3JXRH
KXybEXhzeEqKZDqsusgcY1czvQnLbHtY3KH66Z3uZwmGXz0frKgAtAf5ka5T4wCJ
cyu3+mz8m8crB6H2zu5gcsGTF2Cd5NbLEcJD+cJVvm6yC2G9oPhzOp88kcN4IrN5
vv7s5AekNPw8ZV/gq1PS4IhJK1Lrf6/WQIccVzzSqebBd/DlS9fYnhDTWNlTcIS5
1mgDk5kW4B0iDSIKeG7BNFjDo/wRSaLnuoOEXvNL6qjkopdKyKyFTphUyGLYy0OL
KjmKDV4e9yLhbfoPD0ctIVHWCz3TBmQ3ot3/Tz95LAvBODKbS2vwTxIP+VNOgHCw
goIlQ018pVepmXDphoMsZIas7bnCGggjHx0LnXVfLzjLj3ZYjsegAV4Pq9XdT9YM
hL9MthIhya1f5azO8YqzMUQd6SZjygnhz0+tkVTiBYxd/x1laBKN7+khy5tLpqDS
0Q0qxg+IcWYegVfhakdwqVl4CkNEkMsUFu9qQOmPbDfQGsQkw7Qszhk3c6VGjD40
2wdaeNizDbu5UTKu0mHquoyxDLCDAkKkKRF67No/HjIiSA2VpJeBOcbIo3cKe0bB
hRadBanEdMbS+qi/MdQoVwGqtpZClb2rcrz4D36X8g2Steo+lZ+x92Tf7lL2FuK0
1MaYp1/9ueLJX0Mq97Lmuw==
`protect END_PROTECTED
