`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RklVGJ0MQIh98If/BgN5OXBeth1tIapn3D3gtqJ60MI4zL9foW4OH3LQTgFLDG17
spvlvtuD8dTBHv+nwMOGqb16UPzRYDtsPHC4QbOTXrC5OHXKDrfU1P8+ji92Nbc8
suFRP1NhVzwPniF2j2Wv5oC9ZOaCBCOdjbOsPLJFtHbXc3pC477afFcfef7t3r3O
5uW+E2cSe+o49nwyfzuF4Dg/FM6OM7S9sEhdhdSaJ/DjIGaJyDh4Ng7crez6hbHi
w1FpQYFe/ns7o3PvZgI62pgyJebO2GUztis/TY5IiSSLSPLUrWi1pTEQklW3TrHJ
J9tujS4Np+CWWkLPwmBxAr1zdqOrSeAw8HBBU0fjQLMXRbZk9o4MrR2HBArKBngD
IJNi2s5K8jtrLjguvJOWxgNHMNIFLz5pLkZk2qZt58B55MnUNsrcfUUoRsCsFnaT
`protect END_PROTECTED
