`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/33dxPliQp2oBmVtZdLPKj5wiJiB1IXCcrFjfnFdyAFA47RmGmvICpH7nJY0im4z
GlD9GjpQWmrlAx91KMLGu5YiGcH/pObOuQJH6TN5LuNeM1pyxd6JFAaWycHekSWS
3UOQhnihXt4IbxbDBd/isfrOjVe8fz7rmRLZCb7YVPCzpX3INip55vabKBtugf5m
VFYlF5SlGeyBrBgRErjp3R9tSEjS4NDEBVEHoyGu47+3RMLJl/gZSoofCwaKOyDh
VSBmtB0Rql7A7O9wJtD2nuD2040PUaT3SU/0uhkJe2HXMse7l55a4N3H1SDB3d8H
bw+stNMBTn3tqRov97KX6OQ8NN6uVRn9vpUCZ8TQleYbMKkkpJv+5qeF2lVeawIG
Lq7lLU0Q4n/BKG1rwlPpt7aK2bhs5XzYgAT2HombLRsFAC3gzWDKW4Fd1WmPKZTN
GrlLCpx6FImH46V6XafPAnKfwL+fyAzdJmE+MLkCTAnnIRuMGWrKlyrGac3xFGdh
ZTmVV3GaPulnTkVLzRbk+CHBG0fo7XF2zLVQlAvQijTJ+xojM2MY/jgPS43utDYf
HpjdK75npJlej0Z4otlHXwKqmyFsy3L1scz8lQl7pGGaXvLCFd5cUkeRl2yuFpY3
EUmWAD6eClt5Nt9qQfbmPg32iwHWl1ERMPPKxXuzGy+hyw+uXpas99WRC7SrU6oS
NCdoCQ0SE5C1E7Mh73h3xgEo895AqZnKzHaFWlWV+IOSjnCunewyanXDfxSV46vw
pbtbhJ+7fSXSOpIRMWfXvJJk+kFyL8u/sO+JBkxcbOAWobilmWEMK4zqso7wcGJE
qvPhJygiZzIRBACWxu5hJSUIam2iTtaN2Aa8cKfBC69tf5ID+hPUjxUK97LLy1tC
SntJEJAv6NwfHShSdqZNHJ6h5WLMu8+fwI3rDtg79lnGCaITmLnw/wdbFSJlO4Wl
vAir4oH5i/un/E+Hjo+HydhUBre95gF3h19zrs6z/AQ+37R7f1X+xBm56iPdYQCg
WvZ3KiK6TYIvKgl1uKMXcd5MYJzXfHnW87rtWDQoOUt0jfLix9Ir0OsuxV064B0t
XIuBe23uiK44cGnOWOUhXRy0fi99h0FZAAa1qBMtHfGmzasph+EiwIKmLLn7Dql3
TzUpwkn/NqJ8XpAPK1wWZ2NlhOklVx6OLggX5ZV4RsME4d0Ok+nm6n/Rs4iKkUNl
S4EbyZyfYVfYma3OuP3FZwIMMHjKXgMAxOUh0yFyfr1MjYACQms5hrLNhiWAwzgS
Q+yT33J0yNp2/jyZL9GzSy2VtyRsCdhA7ytkZx1YO3/8z/02NDOypx+vXIDju8I7
L2v3DSw90yI8XtM+b2sv9PKBNe4/nmae8jyJ7uphPQ9/snjCnqWQzjOcd7ZF4L8P
eQmDB+ZJGDwdVvaaNOpT6W0VMtdICYyUU21QwqUGOgOvUaS1z608JTZJE4It3OCS
kb+OyDs28jWIGq3h2EZdAZr/1r/JcRSnamC9qO5qKgPtH15zXBdE4gMlCpR6INCk
XoWxw7AVkYPLpSinlrq2TlBh0Tl0WvxmxiLn17A5ktKEvOxTJInV76jZsrN2Skqo
myW6bs1IA+8QEFZHfk/arkmVSMopyA73qVFcD1rewIdSCUGbvr9cJym0x8URrlUK
2hr4X3ZUqnQnN519Ht9r06cOpKk6c13NPp5WqI+MAt7pMKg/bkiYSNyYtwQ8U27j
vgjUWsjQwuA7GMeHf/0sQQIeJ0wqemC0Wsv6qcAxXa0=
`protect END_PROTECTED
