`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TkJjshQvWGvdxCunpeVOO6RrHDkCT14frU8Bv/NcCreP7YT44b+FfL6RCfLgzKzw
HQ2LCik5s281YcsFoZNbBsh4NSJhbGssYYrg8IyK51bXijvgLfgObBaI6DWjq+8u
5TrdFBB0/6wI2xhdJtA8k6rY57/rjtgphK85Z7pbj3VnHvMkLSGyxMCnyuNE4fkz
xu1kgR4Hjo96i3InRxPGWSriJ7pF/ClADCTLGH2qcO334L8RyMLCViBQPP1jWruE
DMj7UZw79dZCEjQ+EKnlsPbodC//63WwKF7He3jrs9x9KiH3W1jb4Q/30qXIt6y2
65XJcVDcsI9ZvCzdRJVl2WyMhzDQYZ+mz30UlZYzhoK/qIyDXCgQhcRNOb95+ASR
uvovceTyquhyfXbKIB/Tf9hFukyqQHD4cxVjHjaQwWCmEG+VwnHwO7hiewIneAxu
vYqFYMQWS3ml4mkNB3bBV4wMvaK9o4QK8AOPmxGIOCodnLmqxlCDKVAm+PJ8ijcB
TM4k3UrrlJMK1nS82IH4m8b7+70N9Rld27cZI+k7fkcOEFxMfkFLnWh1VGq+Jb2T
4fEk1KAIJSQuXwwadOXsBok8lyOZzeIHq0rQ8QofGu5T5YYJDB+Yruualn/cG4ql
D/iU+8nZ7ebstLgysPoIVk7sN2aTdbNp9qxRy7BenqWkOHJ5lXyD2QkOEoIWjTrj
oPbL4hjl8t/OIm3sbUBm2w==
`protect END_PROTECTED
