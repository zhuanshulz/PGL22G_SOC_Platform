`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
238fD38vBMN17kGQR5YCf3TIDumr2Y/iYdglEBxXAaDgC23KBon+6GZVMD+/qZ0W
wXfw8cZCDaXeEVmIRVyH2RF9sJXnxHw8q/mMHEUWtMc03/KTE0cU05b/dHQ07J0d
TesF06RFHBWvx0Hcx+lJKG+sHSNMBt+7235phaIGXoJne3DMaEW318t+YS5iN6HO
9rnTOidVpLgMgv0UiGIK3TEJbGIDs0TTQ5t/T/PhU93JCiK+uPnD9CCI4k9Qxl2p
CCLKWFi447CCY4TOpUvWjK6eZcbyeZI1ppFi3jhMspOEf+wp+2MvYi1PZ0Jxzos6
aO5JZLRNv9jMaMMga4ktDTU9YfgZKM3HhzgKpGpxPuQCnyePS7aBd5zqJhP6joEX
ghX9OXw3EPSidumeY6XKRehd1v3rWJKyn6DrosLM6a3K+SVSqozXwsu2CMAIq+vK
ceR1+uK/168ONmAadYtv3iMkyrBsQfKW+BgPj3wZBNJPGI/qukX2tRAB/mQ9rq0V
o//zK1YXWRB2c/leG05OzSamLa+87PUEKkuHkJCroq4Qpm1bUu47uRVsJapAVRLR
0eNRCwSr7nt+pYBYy2DWk/AsK4IBI9ikFhwLz4ltiY2roDcuP2XcyTVYbOUFC8m6
OUBhS7Bj/xPQHT9koWFLI1gAEwZ/XLv5rT60W5xA+3PVpI940sWsswzT3rH7qnze
jxEUsV0VTy9ZonFl3bD/fMnD+8+UjUXo5ufs734xOeNIfEdDNvR3sUonkwBa5vjr
4o0oxJg3X5Yg9M64ax8L4IQQvfuxINhhByx7b5yXy4bPGfQxfc7JHIb5vE6r8ebr
8WMohBtIQ5+r/ogL/hocf97Tvcb2p33kkAlWP1sYAf28hLPXqKkZO5GFVKNVmfGX
r64XhT/KcUhH1bOiC2XqdpBiOs9k3QMxPKzsOTJWWwAQGePIAGq5ShA+8l6v8rIJ
bvyDUIvOWbRIEpGTW4MUzg==
`protect END_PROTECTED
