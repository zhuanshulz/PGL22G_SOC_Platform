`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uddU33xAcwojBftV1X4g1uSUrglS8ezD5UPZtf7gNfPwjKGBKnsJlnFajzUjSBNs
NszHieut4hD5snAi/uU/0Ck+GWtcAp08F71BhUgMAPfpY/+SABX9Wni4F0qTdcea
tSY2ffZeltj6ycdQqOCAfNoz1YC2cbGFEGgneLJKgQWVV6OyWN9frTMNwY4xoYiN
CIwJ4cGwPM94NR0sSC1kb0mFBcLE9pGDcCMwlEPJTDIVB6BGhdsQTF62CWBa3UYk
x71P5Dw/jG5hUlT/6R84hQjrNLjV32xXRTEHktPRDowIFQiKPQQjGw7xTKWJK+hV
/0evPeiULoqg2Jf8lDjVA+f6mUhaifsuLUtmNssrRiwJ1k1vDWjL/t7+7EQnggKJ
KKPAAR4KMqqEUKKRVPTmXRvQgSynFZbj33Ln2qbdJo3NqLwF7ydr3WnVjP9gBI4B
`protect END_PROTECTED
