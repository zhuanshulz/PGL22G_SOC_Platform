`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qvOxUPpHInSBS/ReDCbTfZI2eWu3LFNqVR82qUU+eYGdW2VF+F/vywR9hnsc5fAu
JJGBTDkKzENPmTpwV0r+R/8Ry5nvmg270ksrSLIcLt6m0ZKUYvwSHoVVsacciXRw
lY8ogs0o+N9y8+0ic2DFMZiWA6phl2QClSq/VmcSEcUH/9wgshzEVov/uwhzxS66
YXNfeYFdwSFu6Ze+GhRg5sc+s5UczvxMEPUi7IiT4JyqwEFYoS+bcsfsnyixaGe1
0F0qygbBLocRg1w3S3oC++3RAmVke8xxNt32nEH+bcx6UIf6FpwY/GQjXMZ3XyNV
hw18F9NtPxOTd2KiogSzu6KkP8AuP2+jDKHh3DR4F8E3KfSkWVDwtIpT+l2/mCiu
VFstb+s1YcsawwqYqJbJ3ZAWE2Wf+RpQ051Czezu+sfThcaNnDBeXRjKv8NWL4C5
SggbnG48LHTyCAtrAOHjEMaMY64zdDNRCMk3FzLRcBIj1xhDLEqJt28MqEc+wJg9
69zJ6AC67k/zVSiRV4sA0myCsO4um4W9aQ/4N4zQ8hnvswFRIPm4moHMY4JPiyFL
No3E4iW+Ub3wi8rnlTpsnA==
`protect END_PROTECTED
