`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7oABMjfiSpRZc0ywDp2UzMg6vpJhQ2U0Yq5KCMnKS4DBwiwrsDw9DHhLRN9P5tJU
Qls+T5jH3d2m4wnSgDJVLi/kz9jujrX4q76GIOSn9QBkf/PgcCq7KQkXyAsyXonK
KIbq6t8Qf92K1IcjsticZCRxc1EVPB1wAgIkzUz6/fC9JBr4bGfbAa9GxMWEntgP
u08lcyISveubWbqp0qHnSuXIuHzVHRqEc99FaltZwl8wFbnyvtJsHS8giEbzQAtZ
4nJB2R2AMflJdsfhxt6dU/eQianX3LQRO/PFLyDkB863QFlqy9Dtphgcu8jjUNr9
Wl2ITWwH8ZgnFncUfaTlsg==
`protect END_PROTECTED
