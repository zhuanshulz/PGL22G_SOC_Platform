`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iQ4qJAucVQCLIhwdFP2DC3Heh8XDiED2Pf+aMm4pGJ5zW7Ed750AXpBwki6A1fZi
8FzrB28nzChwImLJ0BggP/jIVBq63i5P0FPn4OKe4B2YPLDHE72uDgEwEnUMrfPQ
JMpCm9HiEC8XLl1OVHTUQle1fTl7um6yTnVDhHdkVolEEnkWQ/5bllptEvtHry61
dyf3++cFsPS4aX66XKNiAwqwrdiqtZgdEIsSeDLpliPY+BT3OYyyVPJAsvCewxQx
JheQs52M4rw8TSrv0LHrGMhOFePB0IvUhtPxz5keu0+jCI1VUoId/AYk/iPOl6ES
4yv2WyDsrgS/pSibM1DUHNONM602KXndxAtqBWSCeeworES//NfyYscuX2XaTV+H
+xnFSp6q+SlYrXbULz1SynrhRjiz45tOz1Mb7eQYNff+zgbCSNbzpukIZvTuTfx8
XsoqZKCZOp0ZdKX5q3Fl7kNBzpoRej5Zb7PCNFbx1hNdjzq+xFyva8SFq6N6eKC0
keipiOLWEj7ODIh+HEqdSgcUvljNFLvMO3fJnUdvgM0=
`protect END_PROTECTED
