`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1Tgz6sy7NymMLWS3LL8AhfxSHTp6mQLnglzqDbsCcNUE/ji+WfOKt/W5Smu7ISf/
UQTMpeQJ+LPU7z8m8VFBN3soRJViI8Syh/VZMpMkmNSSiiaisx+6ujq++wLtw/ho
kxpGe/tYdjodYRwO8qzrIOt9Vc+4jWmfcyHY0gdcJfby7RL0NFxcQ2wKA3xnJuf8
7VCTMDs+R2D0m/O1Jk7XMCvIUbcgykUg7FzTM/AK9zAM76W6sfti0PTjlWkNeHzT
BJG4Ke8ZiZkp9EF+flhKqtmlyOFNmgwWgVp196Dx4AszDsmLxuCExk3PsbqKr2PN
Jth8tAnjvMHO9GQrXsdP5E8Ft1QH18LKkItc9o1YWQt9Sg/npwHlMfMVhXMZio8K
zNZC+QQDqkSrAAq6Bfft7Ygv2x4rdGC/ykCpR8aTzp2bB25MY91OAcRbTUc/qj07
t/smV8egJMp+wZWmxaRDNTYusnNICLTjEyCGM86Vdj6uDw9JX4lvTEbw41xW7nAI
yKdjFmTUoilj+9eGlBfcGKQKKISVXD9IoqrNsucVq6tt4goV4gL8OHgUTN4GTcPF
RctfrTfG7vhSH+VGyVXgGwVcoOv9F8nhHChOUUXJGOsg6YJBOq4TE0H2sVuwqtMG
hZMlm0DwNJ2836Hz3t0zk9y7bAt/t5u26RX1DQ6QfmVp4owZR6P1RgF4VKZ5WgCR
t0GUptMOano9D/OpPn7BZp1wZdYUJDzLZiD3MPIMwhHZyArybGyPOZ8ZzNZdBfe2
v5/7hVZWhOpU+6zktz9FKpewoh+TWSTAb5N5LP/EM1OgIEFOstrf8n7ZgvSg1BA2
qa53SGagCSoMLLmoslcpXJ3ccl0bnPXM/K3svElGpWoHy74YW7TSKfY6PB4P89Q6
Q5YV3qCJH7/edR/ziTrKpbrAq8hr0IGMWSkufRlGXWuQiAaJo+dexBDwULKyFnju
L1ZDutIF9oBof+i4LiEWariqYQl71hXWM+vmsxIc9+7YE6gVXX/IJsXkQCQoZZPG
tzFFjrpTgU/qMsXzx9vIrQKWCuDJbbfWcb5EMfhUcaQ0VlrAMCWdlTbWMYnpEa8L
OEmxoZZ3f3I5QNgx5VqqKvnUndlF6JhytBQX7Bv3sAcNlHAIbiV1fo2xdTHn9M9y
3f29mrpOvXItEupf68sdkJyWjH0QybGUqx6HdTm/vwj2n3Lpv4JoBt9c+OoBQbdp
XxJR0G2X/g0ACElla3lClubGx+cJIb2Yf5eILbvEnWzX72R0uDTLhtBpx0Yhb/6N
o+nkLySVx9fh78UkFbzKUnYvYrqD7RD7jH5rAdLgIlI50wvyoDE9ULxosvgwNJJJ
pscdcsrcJ+hEkX2s7XsFADmD03eC+yXXncJhp4/5dgfOL5yPC4bS40LWVJwh3qqS
XQot/HNyb4T5InEzWo5TyvOi2ZB/eTNx5B4YdxH85C+VlkR8UxljmzaYnyljS3Uw
0W7eu9v9q6w/pZhUYjIk413e2HoId3Q61V4TXOZjP2ttIkqBR6ElDMrYvqq1Gwn3
1yFD+BH1+h4O/Rc+vE9Jx4HjKm/gdDDUMrhe3mGzAaL6n4CQGo6HdbzZDLWtr7pO
xeqznn1GUXwh5TmUdP2O76u91jRiu/ocOzXKgua79fNLHjboQ9CLkeKIiuDpgvwv
ueU2/ieZHwkQzUzEivBRgiRk167iasuvmYJpFaIg+fL30F2M1/bEArbHax/5XHV+
06IJz1CyPmUnUHowO+BdQXyQrL/zpuu5hX1GtMxhfrPLlT0DnCH+3Ep5tZy+GsRd
+J5rRUwZM9X0xViw5MfrDMXsH1e9sIZafh+Q+dDfLvsyL1yPoBFOVdVBtVomPTO2
JhpL3ByWNuCRZLtA5vLL/IK8mhCFZjU4j8v1lRPjedTGMHUDEAnbIcn0mMc1QLe6
nRW3YzoDmiedWEa+lYEYV/xOajU2zgHrzmzSZ8YuaB56JZs6X4XVgKo4ZFw4HXI4
5Z7tq/785uxUGFXgtkSbAlNMcoSe2+Ia7JqvJ55aTu7U3G2vBclwiSM0XwZGt5Pv
WeXyfE2kagUEnnHpfsvlUTUOPmFCZXYRlb53hheEZuSVy6yoUvG4Z+CMR9Y8M/2z
X29o33USIah14AG6kjlcETqdpOVsvD8+/6RRzNURe6m8Dw1pGFZKUv/fE7Dhb7m6
8KCI0xvIVkp1fjAyvA0IskzTL4HcgxU3RmEH16n7sp/zgarLv71Kdl+UJPThKek7
TWZioZTgqQLFhIO4CzXjA7Xd7omF+W8WHpzkl0U4drugk6nfeJlNPxwEdWoey9MG
TAUYNlQOlQlnLzGiOCsr7YEcow3Z8/APaDOSANh+lUcYYqKwGO5odMJy+xDEcWi+
O1hkpy4MyG+bh4bHwY1JAZe+8aohuE0GyXGdcPWKR9lDEp5i9GUMHA9ktu9depBw
XzZeVgTa+gzhZN4LwBlZz4yxqK4SNmkg9OJV30wnxZraN/bU3taoBn9wqFur3zPY
c27P7m46FOiV7CPr1vv+l/hc9+E97CYen/+fVwbwg/xXRgnQBd4bHQTjZZ/rnV0O
Prmhmyi1id8pI78XOiBEztyeBiS6O03htxpWNpdR6sogwQ7OTHET82f190bYINgN
o1r4aLeVX12zBrCk/3MliHW9u9ORHWcb25C3RqFwnpVZgWJ5b3H6CBqadkNqQDSX
AF5tbtccQXZaQZfi/IQhcr0nNKyIshSkkP8M+KqcVMoJiEQ+8qEOA/FipiAVVvG3
eatn+dRwiJUkT3ErFDLFu+GvA8ET5s6uRCCuX8vOg2AYLSe1ogp1OflhfnAAw6XZ
b862XBRF6cVjeXS9QW0Fbs05Aw9LuPsYT3ZOds1x1fN2sHct1XiZWvCwwVt1R4oC
3gVgnJcE9DELUnIo3kgvd2DBZMN/x2gGpU4SM+UlwnhoIesvRajtgXI3VIltk+UP
C7yevU/QPrJRDARtTMo0qjmXsOrgzYC1FNqvijomT9+EmpbAVpxE0Vr6VMllpv1g
A4nJ8nG36ayFPbgMfy67szaJEj/SPvWcmJPG9rw68WmSHsRSDN3zAYcyi6CalOsW
Ed87lPZUXRVhq75f+TUpfCcUQoSH0aCGWomfNyxV/Nkypn3hPVRy5wpvzGwtbKcj
`protect END_PROTECTED
