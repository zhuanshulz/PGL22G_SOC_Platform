`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qNLiyjHBkFMHSg5GcNpx/ZpA8KODsVQKxNzY9b5lzmShVQGtNKjS/QBhTU1YQf48
C08stC2wJKjYa4eIVkBQXUMk2BuUXb09oEBOqRkTR0UqVY8DnGPaH4kalRAEGtdg
WkCOSroQRBDME9k8r3ikk6cGnWARvJ+NOYrLx9ZCzPaeC8Xufc8DT85u9SY355gk
ot2OMsvwTXIfhPXgeOaoxDOeit0IpH3xjItMI/sLtwIPrg5Of8G0Iy1WE93GpqtY
HS9sHw9P9Bhdm/Qr0nTUAezXFqBprJ6SaSxG4gwNZz1WLYMsTPaLwl2sX/a3O1Rf
N8sQaTiCuL7Dn4uJNVAVB6c2Zj5KULFNXHx/mDMzmwn7nYMFw7FbHLDgndiDCYR4
hgO2O3QNueZKkfobjjClH6at5vvb080PnH5XnKDI2cYsVvF6akUe6g27r6TTTgNI
NAqw+dxpAXMhtSbuy9Jpu0JArvbp9Q6Q3yl49GDn353/lP1BKHxl9y2aZfcNBBLU
CDPpuVyK+NaZq8L+eyffuh3lzFCdfchnYQiJLTCYng0OuWfL8U+u7mv6LnVza4Ki
iXT3RF5IAmNmXadnv1lQlo7IXoG7Wr0z8kqsI5MOtcjB847sNkXChK3c0/X7ZH0r
wBi37J6mx5IZhQOIi6YLcjCvlgDVFlbi447A3VNWLvuXf6WVjgHNYdujyDOsLmt5
`protect END_PROTECTED
