`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5KuLIVm5Xn0jw5XrLFeiMKdS0c28ewkF+jwS469/u+VFH6QCd5+NmKIT+8Ff/7Pb
Md58KF0EArbuiD/JxxFJU9cL2ALx+mHf7NrimTYwUecNcZm0y4wcK+4HtaKs4F8+
o0nZBUeoHGvDXVROlLSunJTdnZv/++zK6UPfOGinM2zX678L/1+GkIyIuoU64zQb
6OtlPd1Jec5lCtpQumJtlTpslXCFhXQunF5PBDCndlVV8c0MoP5l9rDHtAslIU4m
cw2vPYm+4sqvAUioCMlHIHY0Y3HZHwKGkyw725Chf3UlVTw6LT9jz/Lq/zaXL1cg
hBcWd1VBoM10P3i0q5hAup5ePf38C19TlLYVGQzfQ+wTdAuXEZWPYHFmI7NnZw06
LMxXRV67+yK2NKeGKZoE2JokCH7rlS1hcFTh6+KxpdEoVv0vPABuKf+XQv+0bSgB
gmO98ia2E/Krnw3A8m9BhB7WizuxotVqX4eCAW+47pGDmkyvgZHJ36JHZrmIwOCH
7tJF3lG+7wBlKx/KxIDLGy45CWA7W8qET+C+26iaEgmbLlDG8gPPRAhodkzTArRx
SBI3f76f4BLIeoipkOFyMtZPbonjTzMxRZpl1DKuzNY+Jyu7fd/Ij6xmHpIi1hA6
cqxX3fQK2Hro1TRXC2JIMdLBYARlt4TascF58Ob1Jjz0oRFupztLmZxmbe4YjttV
G3NerRzZWuaINdJHq1lGezr4+mX3w6Oc5XhpukEE0SWWOkvRsr1vgr0IH1INdLak
HhaQBA6WbGrducWsTlNlGnYv8aW6k8hFSvEk5FQVmRHY8DNFbQE9kJngWfCW6WoI
I/gptJ6qkS3EjF39EqMnIgZlzll4iBEWaXO5xs1rALVykS6dqgKvHpHJAt8i5rnl
L1WM5PP5MlXu/NzXjkW8uw3i0BIy/AQa7fhwjXryvFOHAAgs17MWeDiFldcnNHdt
DS1Lc/GHq/sg3NEyqDjBRIOopVxFTsMqYNKsop5ai+SEmBRa4i8EojbvDSglybAQ
DZCg7DL91FU5jh8gVRmfOUjRALJvyT3v3IYRnKJsafujZCKSimMvIPwifQueY6Zc
GvFyesZdAGPSHM67WpGrAVpUKSMk38RNpgFGJnPwmZvE8s0yYyjLKOb/Yqh5wUVM
3ynRmUrDhkGXlwbktRpBIXMKA5FzOsxuRZ1uay6xsv9onnoH/3r1pOeWnOkILD6z
/fWApWqAp28qSeeWbPL+Nn9oISa0XyF8BGctNW+1pbXedK3BfS2S22///2uZqW8r
n07+AQgZzsQgB3B3VUfWf7jINUb0vmgqdPpWZRiyA3BMjnz9Zoh8BlQ+NlBnjQUI
e74w5Xil29fBuOdlcM0fGopgqZmEhhiJhmCVbUZ70+jg9TzNFK4uRVAvqEEDGNFJ
Q6PeDhZgwUVKXLISoTXbVGDW1J9vEA3ovfE1u4PQ4G5RPVbuovcK0zK9ptJATe29
308KsejXEFwAITUAKqmLjAPkZGry+VFGPPHHNEFoRf0Z1eHpkgyI/v9eFw5wati3
S8PpGH5LbCymShjP4q40djBQaZVzKrxshqwjqu0jxtem9SBQ7UORIBoqUvSQN/68
408sIg/yrkoCwlt1UhsHeG6CE+O75QshGET9JyCPGSn/C4POcpI1KQTVi777y0Vl
QTqadb1owaMMX76lHSc8EA3Ug0mKtxAjazQuRBIzyIGENz6PJLSRdn80L9PC6HFp
5UZ3OTuVekpzHAMjLyuBI3lKBd6bklynXCWGswgDrsKW+4BNl461AiVQxnettnju
OXo4KKOgjVPjNUYDE//A08JUprf6vwDJlpva6GcY9YvZFbTFtdVaBdRe5ZKz7nA/
R4KfgWDhiWtioTAfIGmuGP2Y9fltkBjtWwFwNChwd449hIVvkrjUn6DeRsxsZqSP
suphudxU7l69PLmR9hFco3zxLexSOoDJrqVwZ2evakW6K2MwT2cGrCA5cCWJK8dQ
DBxhgkreT09BdJvFuyPLQThYN9xPHX5Wo6JCvFyv2myobAKruTkRBebj28oFGs+4
o9KfcuruC9GoLfM96QbjBN7JwI9iKxq9U8gPegfN6DR5TMJpOpKa9FwZntGNSvLM
RdvF9Oy7qpcD7aHc9lW91SAe3e8tjGBTErWCSJyDXNDK450n+RZ4aD+fbYN6j1Hr
fkQoSc27QjVC23YT5WSV0Di3rdRiD4qFQSl9OR+pGsQeB1AUV3glsCjfcTMHaxxD
pqIWpl+cVHgJSJ8j9L/8LSr6dB0TpDUQap5qvAPnaoLNv+9r9IfCcofHi85s5p15
T5W2tqpOnMJE1Ab2C8vuTUWUmdNM7oipxI/JRULka2AwUXsy563sFXicWkDyyj/R
t2zjPq80lLVmfbtLDyVAYc9VoeOHoFL5XcKgTlnzRrEQ/OGnB8zYZ7xsouvl22S7
lL0AkWc8bUMRAGioqNMiB8e74X3VTGVdWtIZVtosWwODwgR2vp0/x272w+bo/fs+
9XaIJb3UMA6fmpsDDBQ0CkB2EY/J8koa5acVQjM7Qgu6VeSr22lTFHfyKEi9AYfa
Kyk6fsvd0bTs4X0wh+I56OoN+dLA29ckEAODGUdI6falhlkPeDsgq5n2cf0X7w0l
0Yj6sgyyXWHF/+92cUfZcVEr/1xCGOtiMLkCCWd43X4EhykhEksX3CsO7A+Q/VfT
HzDRSPunMxl9KjRjakw88Qjikuf+2q1C6Z01LuDZolNK+s6SU2AirDWAcbAGF3pX
Bq6L5PrZAEzsMOwXou9Gu/l2uwdaEFHIuBShH/Qo9h9xSpe2b0Gc8mF2wGn84jPO
Ua3oS45uxBZxvwlAucLAdEMLtc3EoudaFP84kLtjVXP/7hBg3elveOaCmA1vlIjp
J/TsyfOEJmKt7pZ/OqoqyYRCISN2snpPHxGI26ayMKvikzoDIKLglclxlp+4Jwyo
K0iltSqBit7itvMzNepk4XOkbEhC8nKhgOtJrjIloFsRV2UO2S6Cj4xFkeYUgcrB
Bzh9QKIx4WpDdgd7l81lBd4bJttIBBhlGMxgYnCuFX5xQbKvYW1Ov/EpDAoqTYTw
hQ9h+PN7SfwHexYCf0FY5pwgkmA/KgshPLGNzDtKZITD9WYJW6nfIv0ATBrsfAn4
wqFeEkjlqCh0SW/VZXYljXhzv1wYb0ooaVJYpfGeoZFyc2lrQPTjcz2nMeVOtk/M
PEi67NCzufVqr2+WWmwyDkNg6FiXAVy3mX4rFM37S1PF8BKY6nE0EK4kGx/rPr1w
orwkxuuRRnLJo4RnPQquSwp6J/glxfNFqkmRORc1pR5n2DsCA4GB34cdAxm4ZBgH
6dF+99oIu9j0MqrocufVrCAiVZ9JxGXPGgRa7pZHDGEoR4HFLLFGoe5YFZck49lP
8ztbu3JTFQAlYO429xozr79rl5TvC69OO8AJhcB3D57/uZlOQ3WZaeYTKK/j5Cl8
+cxwtZskV7nLhX/Fq6Ilek8QXq4Et5GbFsL22Jdn3I9kKz0aLavkADOZ4m+XE8sZ
MP5c+Jj7RLo3PgagA45cxzdiUanUY85pYv/UbtXGi4KOB3PyYLAXVB75FzsLG5vZ
Nve1kQZnLKKEnKQ3wDK78WU97/vFSsGAjJrFxcHCcCn5uLDgyID32wqvNqQethE1
q7AEi/V9sd5EnrW9OHWalbzT/eFL9nIL+DJt5Wun7lCvNw1QgjHWDLmBp1YtSQYS
LRmuv3aO9Zl5T5QijVn9RP88KnRjuN3SgjIBFxWHThrZROyNdABQMYRg7h1/uFNB
IKixTNlS4iQrnFVPIy33J6enoITYvosuE1Qxm7DQS3SrUHvMB9eAqjUJe1sHHn8/
juJuAhR9Z/yIhU/qUoTWLTxBqISGMF8eV11sQQ8uCv699nCLniaqukUyj8goxaJI
4Q3fcJratM4ZPlSUoNdmar+9uyL+BB+OX7dr9cjJwA6O42Yv+WGHFCMdBV3kfxGo
OH4dZ2sG4c2HDdolJNR3Q+YOrqXVQBviEbACwVFq+1ZOm/dq8yGGRA/WbjTSWrPs
IQgL7dCPa4xPUEkDyJse7Z4/1Qjza0+pqgAoFrwO/bvx7zRhisDgY/oGby7W8+kX
4jnhSTJS+q6SMoelv7oFGaVe2MWVzjnjMqylyzoTvW+R7Vjfv1GMP7HtV3z5jfex
e7fxccWa9Ly/nxppiRE+ujFHE6yDuKF9CNHbwNoyjrO+0CbheiAtGfdLy7BCWj+F
OLC6CN717SXgJKUTlQOAIG8sAAmWy6KoyCOhJKSo+EOoMEPzR9oBAqVybBq7INCo
2DRVjXHuKK/8Bzm6C2pgBNu3P1o4LPRTymr4jqh3IfrJOGPeyQuvvB608Lu4NIxw
Tq/O9YL6I4JvSQrm84+HskimTsowZdM0VwGR/oqnS/plukZTp/efjNxBfyJX12Wl
+TCGTZHn1Xm6RoWFFGpdaY/zvfx5QqEwmly5I6Jq5iUvY0VDPi/APMVr+8tqLZmV
sA8XSOoAuq8S14OahgVouTGA3ftRKCQ1alcqQa5nSukU4MGWXwLgiHeBfIxmyR7Y
cNt5jRrKyfHuYQBxoEffrtymOihkyFEdKu+CPEp2GBIbuljAqGdDvV5nRtDbwZ/I
Dj9yAV7YGX2RgR6Gwrhejk+m4cdBTx1wk1IuSuUKPp8ZJjKCrU/GGJjJnRgNTNi3
KMe72y82N5LIaQ+iAPromsR/oJYw/vmFZ+V5k+iwtzJd4Ng/GqyK9x9DfrQB8FU0
d8G+CvcPX2HYfXjlMetARQcR+nWecHYHvOddjiak3l8euHTOOijmhZAP4tvmNdww
il8N+JHk77DnngL2n5bLrKPKGTvFQgIDVGpeJQCDvJpDPzOCCAk9jWf+ypDxmNJM
8YKohIvqXwk8IViESAunBZ9p9kW6+KpveMrtziMDYeVpY07TIKAFakYxP8yEwg8M
E7H6yhK0CWAkIkB9KphcYt9gaJecebH+/dkfl3j6xOzuJ2kvY4Ur8lk5Pi6Z1gp4
PPwTLP/udRjDpk3kwS002KiBgi/tLrmCFaN4g7Ecppo0zfjNvQFAyuWoTeWFNQ4h
3GuJ6K6qUC9qhYlXZPFuHMuM1tjCVtuYnXeh/4+RiWBdDHMVhCnUvMUqeV1J3jtE
mbh4z8zyWKqM7GBvpWCQnZp1vzer7JZnb64jYWBWTRzC5j3aKpy3+CUC0+NxAYkL
tkto7CB1MhqpsUHuaN8KpA0lmzLAk4si0McluWI3SH3Z8pzs1vEhzjRRp0Kiz5HS
4atHv60JFt3jXwHswiR1s2jrR2yp+/BfuWO8LA2+lP/Bz6yX7yLqFHD/4BQZqJr0
FAxLutDxSzqqjCK3AEEIMx168WYHofThY13np7Zn8uy/LXamKNAkGHUK399NTHFs
tjSyFt8NXglPEfF7WmacGhsg2nUddY9eeI8TUpgPG9KVVehgd/cwGhlMm2DwRVt4
H1LZ7MLq1C5KjWtK99qehJobcnmg5v5+k/oRmqjzou9tKWox+RUDxFrDQ6bYtLGy
`protect END_PROTECTED
