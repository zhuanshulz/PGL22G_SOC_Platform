`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vey18kXCg17osZo8M5wRSKrLgnEzqUToWEoaM7b5ijiCf5JA1WHgvFbvIEv3B3P0
T5sC8iZeXi6AYLkKRkp/iaq8c+GHy+TYr0yusVkHl9Gim4H4jj+h/UPNAYJlpzOh
k/Q6xoHgBODQ4EVa74jeN9LxrSEnsbehMalQtBmszwjcpJNnWan3Jgok4DPWmkZ9
wkDFFopV9QYoeRxq3aMd6vbqLcBM6rijmGJaQRiDuv6UML+yRN0Dz9V3rGo2a+Rh
Tp8Y9l+zhyGQJRdZl1yJp1wYcj2ummj5C9yyIaFnxTQ23NVBdZG8/HIIpYdPB283
c2QpNwrYqfb6DPAMofJape2W3yiIKwWl5DeXoQiD8jHr9w83lAGvdg7M5UWMFoFY
Gak7o1EdBYWd8wlLbSot6uXlAkKbY0+f2TLLEDv6FCQySJOiIqBG147MYSuhcIpw
rEkGk4GCmvZyTmHmGoetbbWryVDRaIEJ0Mfeoi1J8au88h9ymhVnJ8wQ/CNEJxNA
CvhGaC0lYKnhzZszL0n7MeZmAVHlL8rzhtCVBQcNr3nc+7IPOfC70I12quYEk6hC
cc6eLKZvl8uePo4u706dXL6jjAM2JgwrntstsYIkwwsFjV+jybLpn1ijVgIHCX31
aPn4c4gn2US8nvmkzPIow3oaqOfCPF27pHLuVtOcsuw+gucoGUF6/avqipQpMw1P
YEo3TbKQfN15xdqtuR7kzw==
`protect END_PROTECTED
