`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
asjRQuHim84j/tTYj8VxD/fwENrkAhbMqq3hNzWxe/Q4S+cLGkkgjFzKiC3UYPfq
GPk73Drr7R+MPKkAOmZloZqdNaquSqpLZhywxvOIZlcqZbIPf2c1Q97EpX/UnWIX
JZc1u5ck30Jk7Pha3w8sKN7mT8NMnlBbKgLcGC3AwouQQLpaxhMe2jFJuR4WBPZO
STRVO+vzAAfZ3d66pB0+ngK2cbUA+NcQUA0fTvDSNoPdXoDJzol9PlpksXD83CNl
215GsMjK15thu3ir2wsRVjD309nj9yCdvROaT27cE9GEYb8mdwgMCk/M4msMjzWE
Fdu6WhSZfXJLOfbTb+T3wh/cYtguruhZ6lJlC+zM1q1l2mD/05Hf1hMKChq3SSJK
L1502HVHqKL7JWfWxnrVfuqev4GwsktZJmJoY/2UjIz7DwqbNLTYJPWz+I2O+h2D
oe/p/2u0WzxtDVx/mvxuEKme8FCYL+i0++Z7YR+kuId8ifL58Q70Qrfw1vH1v75y
MLM+i9v5gvv87Qa1EWVy3+LWPo2hu+kr4TNDuPieSSfcSj+XdmJahdwyyXpvvEtd
dpVNJf3tCexe1uhh45/AcxfvsrVdPcix7q3v2GcRLpqFVlE+sTFey9e3q2UmZGQV
CboFIWIBOqn3wF2h4rVUG1huLJIzBAQKLc+hxNjyYaIrH9PYN2VCv9vWmeFX4Md9
UNRuxhvXBvWVX2Nw74lH3OJkuf93rtqEfih0bkSFotNbZf9S8ZzawZdiuRqzPgcJ
w4EyRoOPUP8YUzQAugfg4gGv1WMoXZcURkzZO9uDiU/dy4lXT7WMsiDQt2bROCR/
Un5JhWTv4aPBsobsC1cVo9TdcXX0zTFCV5FCsDcqbmsFF0APp6N7+It2Nnvu+a/F
Ua8aX1TagH8WRjHJRP7+76WlFkGQenVbw5X1W+3ijXxSxA5uygp7y/a/nV0oWRhQ
J5/Pq4D1Vxyndz081QkI0YcQgPfWzvufEcwtLW0AJCOv+1iwZ3IU3OkBrtf6izO8
AQe/PKTkOTnpntgJQm2Je/t5x45JhOWtDJxLVMigZhzDrkChCEpZRPF6vIgaAH3C
+bjSwrj8T7ueZVC7ArS2hEHlzOn2qZOnK9IfSJv9Chq4CR0ng55HjcAnogUzhgJ5
`protect END_PROTECTED
