`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
maaAPvZrNM9c4+ILrWwfcnTuUZL6eoui0vJHCVVUPkep8vw7GasSZPDq6mMjxXDH
S53gNsx7MnfAEdFXDLeB4zse4fdtZ3FeOLg1wz+7+5BuhthaKcDcG1y7LU7I+Qwc
jyf86v5+Y4NXqzWRhODI6ingmg59vA+r1sGhuCB3jyuA0VrDKea7Hf7BjEiVGEr+
ZwyiQFqKZYJkjkAOqVizNhiFnwcdp+QFbRSK2h3RGeK9IsiakyoeCJiXR7svZ+rQ
2eD/WXM9DLiHoznKF3Sr3XdQJ9Q27gejZPpij4/+UctJBZGpY9icxjxBV/ZLntb1
/yFXmZZCCZ3+m1fmAz0J9CJfvBHjV84JnypX2/gBovYloIDsduShlvLSTpY0wPh+
D5487Xy5ucQ0LXFaegV60CNdQbS0qVEGcc8OOpzTJqH+1CPY762CgpbeVMIftNT0
glu3+qZH+o7c9XiM08s0djBd4nOBq04d9gFx0n8NvD1X0aJ5thMMHH77OGtE5P8X
bOAZYVUcnCiJs/YRmjHURnwNH6TlWpi6ImLCDdnaMsOvF4RxNKdZ+7kZy6s15gcg
xksPyXXqV1wcBl7A6GiaVQ==
`protect END_PROTECTED
