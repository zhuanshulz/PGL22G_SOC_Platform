`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2kCpYlTur/pVJ4GSozMtqYCXF9ih1sfvHKo/toApCnfNpPgDhLCAuMDvxyIZ3wzT
WPFbWHhjOTfvTDgLPyc9rD3U+9eslzYEVSEqNnrdymAJyVfFFpMi2bP//KtqRnI2
o0xmZj4hA2jvhORXjIB5OfNjy86DqiT8FtwTJut4i2IQ+hMZsSYtuXD7kdddfcVV
1R5Yj287iT1tFNdYIW45GfOq3tccFQSLcbPPZ26mxPkDjt+HzFYxiNiAFJzXgIEq
g7GMh+NJXcdJIMPWGT/b9+2+WztBLRcIss9jhHrhdOpGWoWHOoSj8Lr3Tg1AV/Ob
SZHHPPvggNgo/chcqyB9+Hm6iDPiQKJ9ZIg+S4yAm2T8Je1BfAft0TBKc3MONBkL
OqKydEh/6TfWDbLnUR97HF3q+a87BpJkT4nMITLPmR3Gqb5T6FfnDLBqaqZxcXkk
QsYUkSsyA/t1iXH3aoRgQVuMhacom8NRZX8jWTj/7HevwuY8ZyNpmYPapVMiMNPp
AIQMHgLJrtTkKmRzWmRUJztBU25e2CzC+pnOsitsOMtN2mLeiCBhrI/5tWG6BFV5
tq0iuSeU/mctIGu7Xlc79yy5rPiwCl+vj8h9WMnz60ClkwBBJiX4oXiRX2VBQPId
uiu8/WRgX/ZNciaq6KIi69YOaaLZpfUvPGW1pMi0I0++4O6oxEeTAL6aAP9hPcmY
iCqH8yY+Fb5zKmfIGTAjUyyLFFxbGQ+WZVIT/5u2t2AfcAolKKrLetBcl9+Yjv6W
mHlmEdMiEMx0KYgla+p2bVtiLaAduLKC0h16h8BELH8+II2sq5s0kuPGaFG5m3qw
NmASHVJkqVADal9hsJoYRCSrfixmm/t4q0Q+9fReMdi5ZGRlPCGrQUCDQXEBq15g
okpOdKJ6i182yB9k1f4xi7YmbQ34h6bv78Mr85/R3yvWniID5JgJIUqIrVnTbCmL
y+rbhmjVGqEqucXIaHzJGB49ry4sdvXkjF8zdOVgU8Mt/oQqK3rVEbKiVFxasXW1
i9xvWll4JRU28W/Eq/+8BS2LXFJNzFbqzmaZ59GQYAikqIlfLsTF8Tp0iNoxkBgH
2TlGUrNIpj2R++SxtUqjauOGHbT0Is0FvDjEdA7qfcUutjBVvyYAflIzgWYvGv+r
oAa8x9AJCea7Tpo7wcCsf0+2fE8rCDwld1zq4W/uOxx/QvkSvoGfpuJQlnNEyo6t
l28IiaAgHVAm3vGHoSdj5LOyxWqqSV9+NceDDue8vZpxccj1F2ZSy7KAQ0DoyWzT
tuV2sOsMA7f5/558orokjEcRV+Mkl+TpATBoBrQU0dZHD8YTFU+jTV9FUCKnKRwb
Cgt59RUQvLP7UYik6l2mMWsZkzbvYDbB/esk97wG91uZX0fsCJMY8qg6wy2lcTVr
kyV7kicZkE7SeEXsxMlW1dtvQKbi+TrULeJOs1bhwK07N1l7P0Toy2V5vRvbB+8n
Dt8GNwyWxu+7/pLSn6d8tSByDBFVNDko+JFO6DVmjFCRC49DXLvbS45wFDTLabHr
edOPZl7n9hWNrhPm473+VXclyqMG25OqGgrVLY51CGl1Eaq/THpA2rDRIzfyKt/4
ywRd1MNZ4PJiKj6ANpahQLMRIP9fkCIqpi6ol9YOjRntar4QFAmuVqxbiPHemzX2
FfJWisI6XFIm62a7si+pxBLlSkFKCdTcNKju3wGBGuhoOo1k9JAPffk3+MCX555s
QqSYjavgU9b/6LTg/OoLYNaY8ey5j0VKCIAZLQcZ67jgX1JgAE4HHpDlBrYIk68Z
4SuDwPpsTTMRctg3YmY2a+ktykfFUMRyCeUYPZOdURqNn0xtFoMd/Z5b2GlonwvV
hiYoHgVA1hd8Y/JVxpQoSkpmr+zxcbwclLh8WMRxDRJblKMMDXpL5pXGTSxSRDeb
rlxWx3w1RiqX2KAquY+6Bv2e/iBGvwds3qy3aQxb+MhVB6NXafkA5PW/y3X5F9E6
Q2GEvlM9kisWZNry0JWU1Z2b8D5xr90mLBgrel7VnhEJxnY/h5qqM+nhBgIAsRIJ
49tdnlDF6VGefLTTpRvjsg==
`protect END_PROTECTED
