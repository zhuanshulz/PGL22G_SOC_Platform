`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FrYzHHoCQWGIYrvopo+0Oo4DQcv+PrhGw7G04H5AaSTRSM98ROs/CX8znG+0L0Aj
d+DUeLFEVDck5b1qtTN7p0Asl6Zpr5rwI3EAvG6u2HMgw34580PVzjZieNjJKx2y
BoS4jG6WT7vInCNL6nQgnc8Ezkcr6eA198sH5f1LvgUdYaFWqOMxaKPVWxsb0wCR
ZAlhftU66yrqFUVOot2kJPVZMOqpP0zyw2v4uNZ6G1WTkXMtMP2MLRQwh5iFd9lz
HfmRjtIqAEchG8c6ZsxF+VzAXst+yaZNDrfh4PMEWc2cLEkb5dvjKJpCM3W85l8U
Ukto9pVf5rOzMNJlPTA7GOkADvKBOZqTr2e3QuqYHuSXl7+3Lh+fz64jcZDjXRt1
mbFaREDq2xpPDkrGGA4VtRuCwSVanCEbfmKX85aOMcFGrxl70k84GHr+n0jjB8e5
83p01qsu4upqeW7t0KFcaVFelHc1/UrJDym8eqPPdHV69f3zvFIgWrnGQ5LDx0CZ
luoFDXjnGfN6pX1WpdJAZWuN9C9zTVJ+mem80VLyTlegYKAWR05Oxz5+otkqbY3Q
aQ20XNahD0yWfXr2o3Sm12jv4CvggKSvu5oyF48UruSzKBXWyH/BDfRGWKHNB+E9
KVp+IzVDQbB/KWBR++K8OA==
`protect END_PROTECTED
