`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9L0Jd85bCNqVSq1FfnbHSEH7P2sWj5fiPTeY9eZsTIOoTCuDlkrnBS2CKq+qoudQ
RaE9B0xRwM101CgOSlty57d8TY7+oJpxUVp6J9rEpBkZDGcz0Aku+ouXZ/pThjqJ
2e1Hbdea5vqNumVF6SYqSrRZLnZSl5oLEBkjSopm6cNhGgX1F5nFb/Vxac9dhVmb
iv2LIqX/m7fefAea476IBYrI2gegMEbMTDpjlW8j4EURGExzro16I1e9S3Imfl/K
4kVlAIPMpqivL4eNxjq6YtIVCSkNeFVj/lmTQXTk8jLN9FFhhgTlei7n4jeSI3Zg
9tKhMH8krYnZ1hBvs3/QLg==
`protect END_PROTECTED
