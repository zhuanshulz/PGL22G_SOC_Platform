`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wj57u98ph2ynzZqlw7dHdmBN7A/9gsZCYTsMUJD5uzylM43dKB4kB0ZHK1U83n1u
dGsF29DiYu0Tn9RT3ZkR5Fc1nbclzM5lt/E+JJsbz79KZYBqF1TbMqa0w+dLveri
AIN0NMxtTL3XKEWVxYfVf1iwzavMUdPFLR3T3eInklk0+KKbNE77OBZ6zTlpAH9d
Ooj2e+YZXzjhJr39hvl7FAZNBT2bYP0sBrWJo0+vDiPKVjI1Cct2HKYvnqYgTkMJ
Y1WwmP47qMYbkgS81Ls/qJxonS26MZwfxATjMH9UhHPsNOScIxd+8XJ3SjGSYXxC
AXkb+xcxkjG8h+0dr0oNy2jlg7Or92A/YkKyS2Y0N/FG50u8OkeMT/i7vAVv9bL4
MK27H1naqW0J/r1qtf8gNHOm+1s4ObiUqNIuDIUkDgNdF50OqFnhjSJEOSUCl/TU
RyqSPlFQFWZRZto1HkNqa8knNoIjuaKoawwWEUMX6v11gxzUNoKAs178LKg0UmtQ
d40PoWr5l6HIjKyo5+MzTb5p/G+QyxJwg2oaX0FwtcCz6l8Qf6BErsIwPOrX0SdG
pBtXasttRBvnCR7vCky8R91c1CuTOGkhF59LYSFl34euS2qVQ7Ac0YjZ9cRHELgI
yIWZ/eOJPLeG9qVvlhUcieaw1j68rX8+uGGT/vVp7aLv00lDX4GaimUbePVRCvty
7stKmjpSTIl5LC+fDghyG+AWlb6/8F1K9IV+z5+EmCPBsPWKIoOZM5fTfNZkhhp/
Mara4tAx/bOJ4BIxtYTWHAM7uXbfCyqHP2D3cEJNgXINkOWxtUF0oNTQeP/HgPLp
/F1lQF5VG2xoDumxvM1N6jiWkCc0sML+DlUD5zAos5dh25D98MQxz/M0DFYjWNJG
l0zkM/Wpz6Camfj3HimW7lvFd7Vk97zt5OYKA1fQOYLgkH32iJdd/qCdYmIg1QyZ
fvlS+2vjmfrznOeGyVzwKS5C+LikaZNus3wvQravEZS5qRKowNayk5/OX9PfWIw3
34ROacZyiI+xlUzznl2S4QDZRnwe57f38POe5DDFWuGefsGf5ivUuGHmvqt0jUHF
`protect END_PROTECTED
