`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D4yqdFsrkGKd9Zr+VH+DPmEWsvqicHP8W3ov+MaTY9GyPMe7kBeTh7ej94DPsr1x
UJlu+X7gUzVoKEI2uiwHfbgFkTCsuz2ay7bXeOde5ca05R++SFPy4Bj4745uy9ds
Qm2xWW5qGNrza6mt2G0Ud8V4wh3vO89+3gRyH5TZnGz8ripZTm4nUEetgBac9S5q
mr4pQlb7M7IGy/6qR8hsO09pHN5TWfo7dxvTTVfnqVHSZxpS9gGHxxv8F4vfewTk
iYVqjsWSqzvIbRqBo4Me5+rzCtwIkneZwXR53gGLuqI5trFVYVnAaghHKEVXlyI5
LJooSXL/cjhIJkWMTzKdjSAm3/mrIZg9NaqyosRumhRMLtOjEvMyFpnqUHp+ltDE
4o5AXfJvRhBiycrPGHIBhbviGM3y3mfKAMhqywd9vsLFjoOoYk1BEJ/vyrFVKISG
gRsMAVDF+xtIxVt/UPf9LPu0OLQA0xfNTtLwoqHaIYq295RCOhqBHp4nun0Xu9YA
LR5lUtjxgdUCEqyL1j0r7yWecNeuN3NV6g5wWoog0Zu1zg97YUyFNOgXM+bfg5eO
QRSiHw1fuJ+bK+dBfU/Y7UiJZRxbuOS/F6BHLKMAUSbZfN06ElTb63QOS/Yyocxa
ZApOZn9wZiwMO1d4BOr6JKbV7ANMNpXWCqLFwcBOAZepyfyVaitWsGPaKSeEYON2
OCV72D+f049EJZq3FRxmWg+jiEukXLIO1iXU7gnboQlycWQ9jKXUJwjVJPnpATUh
STJGhJbNt5RAuDj0Em66qCOBy4fTc6vScCunUo//+NzK90uRxE5MeXXMMxZIkIa5
Cz6CI/cwjto872YF+b/kp+Qa/tCEoK6H/MPT38cZVRAO4Jzuf9Nl1r7Ah3J+Fuzh
CozYHQs0qmaryqSgv25rpoHjvn9anIKrd0H+y02mrYw0QGny/q2waGVqzRwZSCRR
8Uh996R7N9+pUa4MzpquvopqbFmqcwBE8/tT/0S4n2CJ3f3AqeXsazoZ710i9uEq
rEPZq4JEa+aaA0B6gkycNh5jCyqF9+0lqpacbOwF4CT7OmydMmDsY35sgI4c2Z1H
62ziVsyPJFXi1AWUNmiFhrOiy9yopA4tKPmXcpiYgr3ETfkb2R1izZpfTP7LIU++
Vz66kJB+FWyLs34nhTjcktxnfqgzDwVCQ/G8jfQYs9Zizp3QMDeqUzhiuicp3qiR
Hta6ZxeT6G2XFVH4NhsSMHJ4S4WgPImHkB1V6ir1sogjSLWpTkOiOgTiR5LSYgeX
q1MwyYDbBrJp7XU+s1pvGNQ3HJF3j9AIaeSC7rf/A31Sp3EqDPm0P0y2I9ZWsTmu
yzPflqH3OhVYmrrEvvq07SEeuoU0plFVcagvEh4hpO8=
`protect END_PROTECTED
