`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FqByHZ+9UMGLrYO1lErBKveURPVWwA0wD255p9TP4wk4mVUx1F7opkTqs1HKbxEx
c1Lsc6zRsHnz9vu1XH+0W4udLLBY5Nh4URNcn5zhPJ2UsB/cgM/ozRh9MsAC8tDd
IoI815KMsY5DghhdyD7A2WRXcD/qm5UTCU1EJK/TDkEFqtaNvXzfW6JaDaEOwl25
jCJFM7ic7MWkefDQUtMb5f6I5Br0ox4Aje7DnqWXT6QiOleI7kZK02dVU0Xuj7A/
+gtnMTDaWorXKAtXXYS0i6PzYHc3WIB4GoRE8HP/pmbAmSbD8TPGBF7sfqI1bJhe
AowhLT9zHYuyieXEJZqFpwcHZqqw+Hl+fVfQOkHfEHm0HzSIpmsFMM/yn6v/O50m
iZ2qkLsMa/ZETGpi0L4Jbor8ZC13U4iz8tfCAcwtyDyiNstmuKq0lQ3OroDSdDLK
dKsreRiMwr9ixi4JIpqSLMfLf/QD7JgLG/vAAsn7YO3n45sBEirfV6rfE0APMaAI
p/LgIJSjm7P952P0+NU36ZnYUNr250JdaPOrabyv60iZG/q3hh0NP/OmmzHB6Y10
vUJ7KM3ANVzGNLA8gyrRYUi2c/wiBTwZFyVrtX1HVQTOTKvVZDaP2mMLWkGqx+Ef
leomFOQ7RoQTilsf2XGb8KNti8jstbMBjjUFOMHT9/LPQmzC4AJysGiIu3nlKKUq
R+Krxd7FOhg2e2rEucncOg==
`protect END_PROTECTED
