`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BYqgDLiNVJcqyKlIIm/TK13vMsH+N39nbRtMSWPvKKZNtGJDEQ9/f5qK33MEbqSr
Ecdjj61nPAfsm1iuOGXQyJCeTfwYzWrZWhhkOy/G4QVze0bdT8QOEhgYC9aYqobt
5QgncwV5Uy9Rm0druQO7cGjejib2dkCpDoy+Eo11svuMangAU1foUVIpzuc17w4N
Xld96865q8BUTZGufrNhByJV56KOZa1d+oLabaHX5e6AStQrt/NNE/g2vkZV+wH2
Gx5GLZ7sLY2XxykW4k7TZX11QPmCLZwUk4M4ZU0u0eUtse4FL+ds5xFG5eTX/6u0
QkCoeQ5fAHZ4mlztT+uDAOoBAft53LwstqX1kGN+WrDxXKkHspmCBU6Q7vS3WidI
YkSt6HGbMnJ65/aIbDZhYpGDd/phNnWq9pDJvX19G1pgqYkPmj5WTWtzZiVtbVpe
WsDpoW1p7G3hEP7Qmhe24xZn70WRfKPSAgJ+Ukk7XaIuh7cR3LSyP68yDtTkYeBl
9bhPRZY9t0Gn0rKc/Ts+pHo2cgwBw/zhQ6qEyR8IUTQ2qW4daDx9HHalgmzpnO4V
7pkoJWCaRJf6vvOMo9GNSNwm4OWbeD36nxsoFAEI5GdeEhE/WUTOOASNqy5dT0yI
WWhwd9p1/tFUSvde2CPd6Q==
`protect END_PROTECTED
