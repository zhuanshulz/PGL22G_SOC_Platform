`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QXYC2qq0vnFtsJOvf7IucfW+EKWjBJ0FQo1AgIPYt6u2A4GHX7RqaKXHqwDzSGiR
g1j3pwSbjWNkfnT9PCneT8YN36jB3fxnn7uJHBhizBMim7WhjU1AZwOXjbsoiLBK
AmI8v3GAVE0Ya9xAhTuScGfwQRoH9MjVAa4IQcqjFQOyMXzGZPBW/7g4AfGM4d2v
vwYt0vOWc5ZSSsuiR+PcOjXfkGFUV2worvCYM6x9l0r/PW9AKmyWImGcTjfDR9R2
8uBfxZFu4qVX4RnfnR5+k5g+H5IfPsGT6FGuXj1BY1AcJFadc05uuqx5l+LVlVdC
dAl8whY1pjTwHzehKSmmlk+IbjuhdyHaViFrn2q2XEom3E1KH6dWr8a/RtwpTcP4
24idYdloMKWtzbU6/ogmhpIkz4hHpft8Q5ecvlRMzaLTouQBo5n0Bv7UbrHIovhA
DEGuOQmp8i0ohykTppCZtRiuQNLvgCv9xeO8VZ6mMGYu4bB1nA0YcZqFLKRisjXV
a0+IuybZaWingqkMw5wg2Q7o7ady2rzYztdFpjZKeSF+f7XmxeFMgjv4vdk1cyb5
Eh4G1nm7AJcRc6qZLpWMyLMRBkcsejnHU1XJ7b4S9UymXR7kuNwNtLSVZ66AvGqY
aYwaiSy8pWSXez7YpHbz3N2wwk1d7CBOJP3/gk8p38s+3oUBKTWHrdC51F77t4mk
cIBzViH3hJ2FX0IWeLnTuxjGzFHuvDsKTHYWKEdmsjOiB+wlN0ZWdx8QebX0E5/a
wz4jRq+gP1yRiSayvqA6B3AFc2LhS+H5ouKmLgVK/kLFnCpmzHg7KOEea4lrom9K
D+BwnCCqEZ4x8HZqy3b4xwi9zi4SvbL9WWFluIbZNVgRxdFmgDB3kqi7eC0dge6+
5FG+8MFLC4STk73WaEU6lR615DEVLp8Tyuh9hTe0UjN0+GkCKhRW8ouJcC3eb6HZ
TRZeOZgWeYK5pvqeR6VVxfYWEPGxF8eyyw5G9JT3StACiFawMJXAurkRJGdt+VhN
VB1CSmlg3ANdBxk4SV99TID1HM18ccasXCA1JyWTVdVnxNv4yl+fowOnn5Y12H/7
jN8p6Z/JhFcM65Y8qXRe1VvEpGfYBZBl2NkT01DWjBoOO0APqVRdrdk+sEWLNBFL
HqUqC4CBcvQ+CNHQWTM+4Imia3Gmws1xUX1BQ6Zhqce5IO+MS+uVDlxXzpg6OZ7m
cjqpzIhh4s+gkMtEBTgRWIw3uQfSnHFV2O2jkiymbuRfibNwBwIJzo7+Hdqrikoy
RRQK78qLRWgoHNdMPuB7zr/NZoUcZjq5nsQhk1zwqjUPYfc+DCCTYa/hvbaRSbGd
IQ53TYXQ3CokJQJSOvGkL9F200HEZmhXfxh08rvlxDmcUuEbjrq1OhFaQibPh8GS
lRQ7V5GSGc9hQ6fGf7AZXlwljwXIOik5Ai4STutiBsWNi/8e6sfOg0bP6JxVkMtW
XA/dZEUKUH1eyXNlyWmFmbQOf7ZJc2WDMFRK7hKOTsZRGoT9KDKTHv+ngjsyeTSi
yDdjroHJMLt7JaU8ZKZgsEbOuY5ShkAawB0xfGwB51NPWrX4nkE9c+sCZ1uA/UvX
cm2L5J8IGNGnFrRkk/KoKmOjOllXh6/66y/cr81sfYEXDtOoECSp/woY3S/j07CG
O4A6T4qc2Q6sY1BZpe2u4IxnBu1t6qyIz8MArUNuu1kGKjnJ5U7KKop5o7CAfRb9
a3EiA09PLoMjxAg6gDMhkU2/ZfqvtYmw4C4DLjp5+tPd68NynK0sSn2LWsfH1sXv
pzXYZpb6zFaSn5zVOxGUmjURFks7Wae0Hm8cayvlrqaACy6R4hVyGU9Lct8EKIoF
f+I5I20jw7E13DaAkSYSPbR7CAbeSV5b7VPbS6el3sY0xB2KED7N0WbV7aUN71d2
x59e/MTgg/oQ8M7JdLNO6JY1e2zKUu8xDuI86XSui8qt1yLiy9KKsrizabpmImOM
s1auEkUEbv2F7U0vj1iv2Y9Md8TKCPLYHv+R00Us+U8dXlw7XxF0Y1p0QMlPYBZe
5cCUW/ghHJbrA0K2mel36udFHwyt3hEGfeCBRiRqZVztAT/jMiTGm5EkY12H+vMI
sf5NF5CLgP3ziRmUGD4WxoTLPsjEUGCa94Twr3zfJBkPT4uf1YbyvjSkf0bJSWId
xk6akNDT7DaBIVdb7YfhB03XxXOHiLSsBoj33mLwH8l3VkaHt0PFIh2zYkfzcjuz
yGFefEEorlDE6SLJQpRb/91YRqJQ8iu7IJowYl3lA8cwRT4E+XpSzH1UuPwPwiyS
hp+MJx/IZ9blJTkuyD9QkVA+hrmTonhhfju66cW/gcNSOaDXQvJNGx9RfGqNHYQC
GAL1xyFJwzZxquGcnpPMziCjpYgVKeHgLFE1H50BQCCynoEdI5fQMFg0qB4fWBic
NczdTIFfyL1wRzL8FsR0LpFe8op5o2QAFd+7aF5hn32fo/VRx+mNP70rP2nMWELH
MNRRy+4Act1tGHlsIzJlL/EiJHeDuAA/NHMMalHJM2IL+Gp2ei80GJ68grS1Ur60
TjQ+ZyUvdWkhPKoA3iyg3j6ZSVHJUhSt55qCZ7ur84QSgDLfSISjee9WIAFCsMrU
7C+9j7PeQQEYp8s0DFNu9Ud7KA6kaz/1tU+tNTxCQSz5M8mX1fVGmQSbppFETvWy
4Xtji6J6ObByvNGlSX1iVCM6I5hv1c7Mamz9F0AxOxjHAjaEb1D46ccC7g3OPc+V
mRXzapcPzJgm+/LRFJtV7Comn1aE/8YFAE9p8FOC806ErvjXQC+R4z8npRYNTxpl
rMkWiIShnw9rCm3KqLccJR8pnjX7FLSlOFtKVQG+3ZchMShfgqj5wO3FMfQdYj4M
Pdc2uUacNRaDyfjZxWqjEITdBb5bnbGnOwmd4ZazJO6+tf491pYZ9h2oXBjVEL7+
ZmLc/9y9bHeNiakSoJD+LlJmVsNjOJqRsnLpirK4w1o7k8Cuqyir3NY2NED99zY2
FxyRkDLKoByFI1K1VfasBoWwMLXk2CDLpU2l5YvkWfFPRQZwjh0lMn65mP599jqb
At2+zVWx96euQ0yojdoVE1+VNxW7NFmBckdyi5SQmVZ/5fHcH8IjNxDfTQq2nPK+
HGB/NAqwEAuQ6aqqkO6KzC46EnXF5OsWGuv4M5lbf4KHfrTsOgUlbzaQDffJ07/J
BoctVMPt/mvdBAWBFDeDrGf0sw2FnuivCA17avXePbeN2uh8T4c2vafViV1IihRr
4SvJf2K0cyZE96FQRELh+P8IdPNtwGzyk6vlUC37fKzg3Z9MC0TLrKaFzOBo7E0l
3uKRM2KMelWHbvVhnurvxhr7ZHSKdb0hgzrE/bNZg8WvnPQqIs+iMvsbaZb5Z84f
ZheBWl7i6bD3R8y481mNoX0MiXplDra7sNkXOOB831/CqQMh7DkEkJhbLqJRSc4f
gObNb92hEutrSK5PuvMOpSJPdjnMWlu0/G08Edr+5w8KmdhdneZNGuCIoQ44qBTW
Hftro6gHGXFmAvN0qcWCOhdiAE0AI5pHmav0GiLnHC0Qn8PnY8aoGIsiGFWqo9YJ
A+izyFJTf+V2kK73vyfbydFvSx2rZy2ZXyE0nKAymCASxORuwzc56eJmZsUqZSk0
aRourdyxg8gVR63ri94NkSD2JefL6I88wTGknHOK31v9ImmPYivY4BGyvYIqBRrl
zCerzUq546QlbNzDETkwIIYctqguKvGt4iJZ6n9tKXWdpYsnbq/s3owAx0klEM5d
zHeDtzzl8N3GVXY8VgK62Fy5nu1yx38ej0fod2N8vkKR74TWs8NOdoD09CII03Yw
eaN4P8J7yHHwJeUuLkyjkTpzU5XvLcQjqExu7Lcz4mYrQLQTuVQFxJS1hoTEODzf
EZ4XawkNaVGtl33y2dzocXwSznHowzypfcMeEiZ8D9W4F6PVXL3q400xlH/CYtos
vNi/R+HVa1nApnUEwmEIaMXgq8Y8akFqBMVNs1TQsm5eWGX9CjXcg6v96TnmwHge
BKjVJy5+ItywGjbfvFcElwqYToXYb6ICFeYmzIvAqaKMwJMZR69ZXcUpNeavw7q8
W0B71/enVVrv656lWn+L1Zw1bttWhXizXpXEP9K/4/LEII9IEAZOpJ0nGCY+zVRp
GzF6pdiheUh7APWsG2Cm7UvXV6b8eUMxL7v9xVEtEqA71Lwiy1S1iWKp1EJiAMSC
MUj27HqQmAX5QN8CyiljZ1HtYl5JPIVX3ssXwi1VbNPlqYAwU5DjEsgD6P0Gkgcu
0pgsIdge2esHXXmd2BqLFfLxwKNMlc6vHai1Mx5TPmtWxsOiMPGswi1tcCy7j8Wq
pPg4n6jyqtERiLlmIsVv19cdRnjAjUaZIo8jo/oUlYW1kwtX2op83uXXQ1sSNXsi
odDNvW0NWj/uos+/WOblbmWpHpxVxRjII9WJA9OSrMRwkCGeKc9XCN6BSZwlxE0I
WPvgYrwQzQstmFuKb88YE6Wku3qzFMnw1CqIPjrn5b41nXs0vreADpoLuLCDZT5X
1LuK6Rv5YyWMx7dVXU/PIncujoTD/sRqsZXznUCTX9PND/P9dJWGygf5iGSQSyyv
b+0EpYpNmg5Wx9x6AYdJ/PMC8BqSC6Duz0HCks1y9gJ8McPVrl9hHZPo4dsgLCBp
pI0Ba/vWKrlExrn1JpH4njreIjs4TU6Q9f148Q5g01bhO5GKfaJkW2RDPDbLjtnQ
R/iAa8qfo9De+F6PbwOan9Q8VxFr4hpXrihBpAxiXuldz/l+C4wenj3jr3Tit/u3
3kwZxUJ7JVDrRH45yBWsuY7P3YgAMryePFSODeZplTDLlYtSeJQ6vdNFu7Fn718U
5wiOpZmkf/Wq0PQy1HelxZVvD5sQQAmcLxC36Ckg1yLCqty3lOMyp42FyMKKEbdi
FNuIhBrXWpLzmMTOcZr7GDHjQ1LkrEoy+92HxYV3Yy8MZV33lzf+Yq9fwoO8OvQ2
aAo+NkipUNIAP5qqPmawdowzZK6W7H/ZtFBvxuehWCAG485vsBQafyWPyeYi8LDI
LC7hWQ6fxtnv4T2H1QvJ5yapNfsk1ov4Cu9M4HRWBZcR4y1SEdhlN18VKr+eFvet
ZiaWTNqcZjcK09XtyM+IC+6GPt98fQXnFjbLqkd/iEfibM8C718KaxVpBIMSQbKp
wZoZRTtwdPapME3VlW3KeOMQhB0l4Z+fgHYiWdhAx5E0aENgGgTFpTsmRkJCJM7F
lMPOfQfVhtB8dgZyz7t1kUD3Fpg7G2fsxkQ+D6Ks5JKi6C/JDM6dJGnaDatAxAoH
RQ2IY+CDjONU2acJYyym/ibT7w7AE8Ogc78TfZgXk9dUSyhGTiAkQo+UHXb6eUXT
zHsmHGu2FRw3lqYk5vpmoOoUfxmcnMBOr5xFbwDK064R8RJIWOKr2XjVJq9HiyCQ
HomxTo+HWHKBVfHbb9++YUwbVdM013w4bdH3RHKCe/4FDR6QZjtGguS5nMry9BK2
BM+b+Jdsb9FNCy4Vgzc44l4R0HcQ10WVz5bD1YqEoUfxACUv7gSgoOWvqDdNBqfa
8k/R1LJLB3wCStZ9zoK+Io3tWDsNc0rb8yhRwDaM44JPPiY7SsHz4z/a4BbcT7VU
TCgRFWcTYA++u5TJVtpIunskozoJkTgUVQ8PG8xXlvxTiG0y3ySE1s65kkUEAtHL
90xaPRk84GZo5CzeYKAydkcsVg3/S1VWufX58+4XnoTIOUogqcnnBOjA+nA7Bxcc
vbs4uFo/hszfHcgSCrqWCM19At/XOlHo9h1KyrYITiChMPbzyQixuTRExI3ayMJ3
p5VF43fmZUvGYoeUW+c9uIizjkLf/X9h3R+h/ds0Ba8/8Um9tNI9Sv72K96+sMEN
wqXjp2aK2IKUI8iIuN/e14vC8wilqrIOl1QJ14FaliR4McmaEmPC9+ZCXrzearu1
1twNzHoK9BFn+jQY6f07IVMx39sj1c+HEQHW+SqdwQAI+XzK/WSVjP0UZL0cjv1q
MPjd56mhWRhp+euJIoJwEpjU8dpwlIIL2T684DTIBqNt4vGWsjeJEWwzlPPvnRj1
q0OgrpXmKKWeYfhUTRZ7/zBkxgnOfpcq5CtwZvyMtziMohd159ub5CTO2rivkmNn
7PQls9C1AwhYcBYt50ZOOrdoh5/9af23p2N207DezmJzjhM1CCeUHy39rSbal849
o1vbqqAVw3FZmVrLLo0WU8yLJpApTvewofjPNNHhzOm4TStWLoqflmqQ98XM1E01
Hl+HN0OWNLV6nPe8nhtlRt34IOBJcQWd5vWiEkzrtzM6Kq4v6FRwJ28nGvrWGMHh
1c54+i78K3pyPFk1nP/gMew7+YhF+sXyYfkpry0wwnp2QDEFf50ygIAA152o1TO/
JV38bOq+hrpTJUJyVkfhrIame/pI1w9aVvol8IcU/X0zPkRod6Jjnp5eol3aHvuA
+NPxVYhII0AJZ3CQ31dzyLJA33T0mvIsc6nAn1pQJXasV+ZWQXfT/mcH0Vfi/V9+
w8QP+jWPcbjcBFR6Ibi/r7iXEbJ6on8d93FdfsAmzxQ8OgzIcitvgmolTZ6X0//P
WlAKc6LNUxVaBT/2x0WSUyJryhV5nyhN74ULYzDRGsTm/PxPsuquw+bMNC3QeF7e
3aNE64mvIFZ5Y8XT/FmbuZoaR9Tetz/scESoYr81GAVPfxgpLkmz/2+1hTG9rhbw
+AOa+QFaUVgHPzOHq2ypnd0OPo0njG6+dTIDIRS2SvbRfY7nfB5nOagmzt6itIvv
RZhR07loNH5MgjyEY/UlZt5+k/ozEw2TDn5ZYF1FpWlkYUQR9RJ3Rygod/WXjfAx
ldA6IpElzsaiPCav+L8JFCeb4+mruquqO4ZeVPHheDPwVg7783zzgV0bQYYGBoOk
aQCWgF09bL5gDS42kjurdj5Sm9/N7m/IHMRrGsimRN+Jm661sAH1RJbrYlWvGOwo
1Rof6XQmDF4SYzuLx44uBIpayvqbdVbMeRuMoLes6pRTNlpI7yApj1gtgZdoqp7v
gpaV7hn3k+KoxPQohIBfZGoXozPWVL3ZN3eu1uX+vFiAObJkupO4az1+criNKI/j
putMBQHnZbhH1SHA4XdZflB5BezmKCmqk1dOOKJSN2HjjZ3G9uv6XCQ/PMTAUDz9
ujPVwtb4LKd9pqPRXItyFL8jv+phvNVwwdAT5nTNvEni+y6TrBFr+yhUknWJaXYr
OQC9ZKQjCP1u1pOcZslvtOcPVBsj9QvcwGg5n0XYktHIEL+66PpaR/iVDzRBNmL7
vmS+o8DX5wSkfXsLvzASIC5L3Vwo9bUnPmXxP8yTlPIGPloPH4+Ek9YbhpRjvT/r
c1r6LnXzFLYrfV34NCFxl6H3qNmLHxZssPL9HLCY3Z77WaHFq23nO3ml6/Qafb+D
NqKIPfCUPSUw2qrZvnqmCjOTOWJPlH6SDCfQErf4EnXtwijY8EUZJ12OH9l8ZrmP
74i0LnaALRvAzv6HNc1cm7NFB3JPYFKHi/AuKa3A+3Cypb/MEJc1Xu3N6LvZJvhw
T426c/C81ND3PBT5G3lh8741HiaSdAtO12FMRSWh/+DkZwsabiImymhfII4MI2dw
xX42LLjIAi13WXazTYkXISn+ZzfFGRcx2FJKTaQuF1TLFaWnp252RMI6nm9VJlnl
xG1HiFzd8oZ3ihVMVQK6SD/mrR1F1YREk5476VkRxQHskajKzE8O+pBKc1Gq4iOx
4cPWsZK/vWuBhWf/SZQ9Jz7L8mWoB8oTV8f2Xp5SM7PNShJPJkaA/eKBAMUrCm82
1Y8j3kgsa/j9oeH0wxudErkoRWmNmAUXWdkjfd65uN8ftDPqDiqNVRvR5PwtFs6L
bM+QoI0ihay6ar+sBd1GJK2zj5TY72haKauXohwacjxcurBwWfd+Mgom+cW4HsqX
KlnfljM8bdHI5xeK9VJ/QNbzx2kKX5ZRUkzzaYEDOMU37u4j6qmJOgJGBIbJXN9S
SbiLm2ChncolSxSv883QobUzjEfvQSyvD70nL/wfHRC8N0pmUNZX3kOE2rb2U2rs
lErS/G3U11wDP+9A/pvnPIbrTZDrcbzYghnJkWYfKr5TzaW7GyZftz6C/nNGRJF8
GXBTpzmhjZ0SNiQITC4Wa4Olj6o8GmC8MLEWXV6GO2fhce6LU5n1r9Lmh2iru1Ow
koJAfyhQApr5tjqSpw0pO+szN7Z5h2JUDbYUJDR0XL3e+ToYcxaLIy4Pu30eyKy/
UauBVOrjQFlSzJ9V1NAPCM9T3SYLZHxcu1uDNp19E/nI6ZbEShUCvOf7kWHx9IR8
KC4kOvP0vu6hLd67YzMBffFChRsIFWmIJpltyVN2aYWJI4uQV4N5gjQ0rYHSBE9A
p2Uv1NbBv2hHP1+EhNNl9e3eJZ0HVrNlStFBLKpa+KkrgXI2hT9J7goEHrqDliIe
kQeToaYjhdKWaLWbH7yC68Z/gWuoIDwg4PwWeADe646AmQIXXRNKQD1euKB+8Es7
enrVxwBQG9fLwfVFTXlcHC7hRmvM7h6jGdempl9zd0MZPUV7OE3gO9wTCF6w56DE
WFBcyWzp7pyD2E2FT71k2vF2TJNSHq0q/Oh0V5GGcDoZOsrr9ndE0E38WLQ/aVJq
YURjAkc/+y8esmPP8hZFXHnk3pjw1BvOBt8uzkO90gTgVnCpZRgca4t1AfCuzIvG
waDCYe0f29LnpQDew7YPUe1YUeEWTePSztc3QBVzYmCgW+KC8rHoBqdtQ/ZaarJD
d8+H3Aoh2qFJlPdr8eRqnn+CZhnJ+XT2Sw5mUn8aqW7EiZWggM/wG/RHGlJJR/uT
IjZR4SCRGFQSesDyGhV0jywhrwOFAt9lbP42C0DHDBEnKA9qsSq0RIsQiHK5ys3h
Ps4dZZbPQIxpqGIxoSX9V5fWD8wxZbLYXrvz+5LRXnbBOQXsoQUhEUmJwDFnY4AB
IRuen4d5fWzlD5i5iaGT6d2f6cmQlzIn/OJpDiBQzgUWQfilhWKwu2rzPLevDXW6
808HGJs1h7en5TfDPpYEMI0Tzx1XssLSCLihE4PnAxRyyaI8q4KwrpgtkkVXGLKT
89YlhENotdDp6afxC1Kz1kTjCEPN/DOriFR2LuUdQjByFPdC0Gcj6Rhk+zg2g+49
5smqh5niLFDmsZ3agEI/11Mth+IrkfZg70Z2tuJiYI3ZIPpiZutsGzPh6RGbqOWo
k32gjFDh+S1iVL6j29ZCveK1wfbQ5oSwxD6Ouq3D5kzaMhjlMNihfiv0J2tk7VB/
VC7SC4LVsAI90GHPaiX2wg0krp5b9E3P7H5HSO1qDwyn2NJKnf2ZoNQMnLZfHu8j
CQFTskM3KbR74qGMvh18VoM/6dHem9qAGLPoL7hUNUGuydlEXmjnC2PMC67nB9mU
q1HkygR7xy6W1pP7iTtY5DtOlP59bTjmwHmCXrq0fjdvy2b+O3ELd4XBDYiuK6Ru
FTF9Mmv6IKvIELD4OklW6zOtubgGKtYYqYMKfY7fv7VXKHkZTbTgM3rSB/lBGA10
i4MmCZH62EMRUlEcHuXDris7zzQYOjyHSNJKKWtfOwCyoClkNbUrsnSfTZ4wmYTd
T11jZRvlXf7h3S+RJiBNhUg6eLBFYCYCfdKcSwF6DP3RNOI9KzFAZHwwCWLk761a
BWcL9UUNZit6AgLxNTfFwRrEbVVDTEgUEr+qZbKxwERM/y8xkf3gMm7WWNbUM/ML
/OQ/SStObO6sYmmg7/OglZRq7+7Al+vpC/J64qns/HyCw0BlYFWr6TA4ArY0EAAF
+EbRqEWRYfaPzg3F8suXM/X6kpq7zE8QEbLGZqTCHAPDDQJj2jB/hqkxePZRIz1p
YyEcWooBiC0EnGAu7O7ZgyV4+9Rdq8WQkGM9lOvsoQNV/AVFj4D7JNuuRPFYuHzt
WYWInUBNCOpparZUGWR0tyfUAaBtg+DJnBc+u2Sjli4aTbIehSyF5FzB+cO8rVZ0
vYzVz60ECOfnZKMa8EuLqY0TU5ERH/hIfEo/D0wG34Okhy3AzTBCPfn5e1nPNSg4
wOMueVt0yWr14zpOUgiexUOOgHI6LsVnUc6ylDmucIWim3wXdccvNsTrABvXVSKs
EsNVZfcXF+FHlLXwOID+bMig2tzD+ZD6lVKRMz8nHr2lwxV+gGyCyZmEQIrw1nCb
luXoKo2Q0bp7ImnaIL2iIEhlJ2BeFNDb9gEi4ESX0wBfs58516hT7H54BYdqO44P
Xd6Evj50Og981QARprO+hel/Q8J2TIYeDcq8Izelodxcz52FgqANAv6GsQUyEP0I
RpHGDo7sRQ2EgE/U5YsbEeV+EbBdBulMMfQYyCkmZnsv4heA7FfzDZkIpX4+AXkF
k7WAP5TPmvs/2WGTzGTDvYF+eef4zX9m+CeuxV1n3wrSy3q9BhqmHq89KOyV0qzU
Eh3qoJczH+i/hi6OVs2ZHpAwwNhvhnPmlIhnszsIeghEIr4E3iBXv9oXaAob/M/J
g9Cod3O4qIDdDTReVWyyGEimhrCmkr7CHs5kcCX56sylQ5WnUxG/bbLfR8UKvvL0
L3kYGvI/lLvHmh9d5NJ71VTXbCl/julfxHL1iR2ZPZI6a63RAOhHWUNQNzKsWc9C
pffrTYj6Ji38jVgNUZQHmakwDoUrIsz5gm+cfHx+n3ES+6g4mbPkauC7rB9RVgLm
4uJpTCtprh2P/QrG3GXUQYnAc88Edv6jqgoBo8onIGy+kzi1JBxUr1hg/WW6+TFV
OSojAFbv+V3DpIAahr3fBvctBP/6JGOBjf32AQt6R1mIZf8QHlZ6GNEEq0svwagW
gsE/ELv1F3jSw2z17xA3GRUaRhiqdbSwZVPo9lPl6wizDUdqwEpWTQC39BHaVw8U
ZhNr2Ci1xw1/sSbOv6r4KGU00QLDmMq2ZPMqx+s9/8W1LvSUEXhRZGkg126oVIz/
VEKr7tLGxFITumUkMBuI6j921oPJMbNPnrBLeVhcfHA5+sNZF/temtQUF6Yd3ayp
inKtM2Zbv0SeWG0KDvjTzPNl8D2i29SVrKwLBDyCNMHVbbkCLfCyjyBl9UU7OW6+
1TbmXYuLC9hTC3io5GIssOqInoffVnEwluGNR3cEkRr+KZWxXH0+Fg/CMNuyN9g3
ucIjayA7Mo5yarDNq60Ou8Av1eCjjHptzQDKrrvX7T9FnsNvEQQwWlcIFP4gL42M
BFUjilZHjqJXrBytN74oiivKL4NtgT3cWGhfgbsmMynDnrNZu/Z+2gUAJz0OSMw+
hTfzNbxt76dLKGYDv0dTG/fl8FBY9hcejZgkRwaSQbV+WA5iVK+R/8yIskF8wLSD
71pedTIGPPxT6Lk87v2i9XenMduvzLSpCiC+8z46uFrMxtXEkbTJY0+qvm1OhDHY
5qWJQtIfdnrimFNEjD/f78hc8PhprhzYPuqYE3mHpIvskoe/68Fs4TC9JvClLs6J
pkBdOR6qSU/MP4gdinPMMFT7YzQRPzSWAMoJZID/Zvsi9csfQC6RuGGcwUjwlO6b
DbH4OSpm/+JGHdbGc1SKNyMODyvl8wATWUZgDIYCitff9nf38R/Qq8LD/AeFjy/r
fIYOGkI57CQz1NywtrQdX6zzVM1+d64WQaA76zhEZ4CR/FafMBUw9veY8QEi2fzK
Tt/rJFo9oWhqVQ56sOnZ5ZlqbhcgoKE+1yk2uUfRNDzhQr/GV5/FmTF6R9uB5BbM
DQuyqGmUMyrHMy5mZ+xX2rQZMNwCB4YjlOi+J2Bvef0RjVUJY0Wtho6Ef/Lqgjmm
ZvK40jpnHIfUeKscEQyS/JxEDyd/gp+wompmdO6/R26+utbVvyDjEuTI/RzgRkHj
e+TxtswAJWjr6D+6JoTrkc8FGVG30tC67Ot84n9FO/LMPdFcejpwtU1yXfeh6TGD
B5Q4XGtwZkONheUxE1Cisa1iFpu3E5MTVWZK+1JIlxpz0faPlMqCr8cA0E1k2rx+
Y2PzmYzjKq7vqTtzFLrmGdVw6eScNaj6SYxP7Izndww3sa4G4xddrXLXHhe4fGB1
zZBGLMU9O+LHHytL+4rcjozVMtSNBssGPbm2CBHIsXYeWL3ICvlxBLyeE5XZGEZ6
X6LP0KVp61j9Mi8ly8xlEpUmKdn1ClgWMFbGNMo/cvAsJ6rzqDQxlgzNFRltfJHK
ArTGKR1HSx1DquZ8RbLX+0MQ9VQWrRCBLZ7kgwr7MSKYRcoKXwJPHVIg4cLtjWzK
NSQ9PzjPZ+DZbGltTGnvUm1Ju42DE/Q3pLkBZD64lvYLjFd2R7XgpILtpt4iEBD7
Si5jMmUz1yhvhIqkbI5AafN6hDLyDn8SZlRsx4KlqPT/Bbx3k6idN+jhngRC+fvR
3uZn55nJvNDiPXr+iDgcUTBWcepYK4/xAIaJ2i0k1KWRX2nHcIhM2fyheXawq1qn
3y0mh2pZ0tYLqh4xMFJ9HmgZApA/aTA9QWo0fM3kzjtq6POrCJe2dPtjNNO8GQJy
/F1mAyNzpbJTzHf22+w4bFQo6U6MhlJ+W4mb5gmScuVR1KUlYqYEY0T6kq/NqexC
/rSefnKIt4sE+PcB2FFCJQ==
`protect END_PROTECTED
