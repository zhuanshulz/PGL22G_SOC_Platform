`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ml11vJEi1ucwCTKlU3xITXv+r+XFmQ2zoP0+8GPkpMPTQce+I2N7/0fo6rNhFUdL
zvQEMyrDzqSIeM4gWqaRG6/TDAgWmNqpJkvHrTd+aOwnQGtvkBBo/Py4HvZ4b918
23KLK0k9hMCfiYPcP/5yCeT/w+daTZrH5VpkJop3z4fWvOZk4Y9ZlxvZ15udnoMI
w+Pw2QI4tu7mJ1vaBzXC4wsE9tv9QtJV5qCgHxDe2xS9H1e38xoxl8fKmsy/NYdU
ao5gBYrwEzYeg/mqpXNcRIeuRrarrfNRSc3BqbGji/6Itw82fgbEP3/v6usEPH3G
r861uH9fo445yY0kbRO4vQ==
`protect END_PROTECTED
