`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bWiYxovZI5u7mp1lxzXCb1UOZv0wA2YYrfgzmmQWNOJM/vacIdw4hxEWIElHqnLk
HkFuJqC9nl9wN42IDQ6JoRbhJYotSQkE6wMiyFyMFPh3NO7daWHDn3Nh4DvO8dFJ
z9rrcrDm8kETlKAt17nOkgiD95ETZEQzVUFpNB1bdyyxusL7XtfeDyWU8MJ4UMQe
k/NkskCZHs4j50aBsMjBlTKg0kEr+pNbDVsLuB6GT4J2zW0r1WVbmgzt15KDrKyw
YbsoZfUbgYHzr1R3mZCardrxjSPAVLSupJWM7rLqe81ctfY8pmo6Qyh2C/tzYhMM
wwhEHqvQqmOcVxAXEuIHzyPwVqA2RP1PkVhCHcGYym8S+P7qqEX2lo+0xYKiszh3
a0I2QQUjC+C+3OfL0aaWOhxBwBOaQK7UhHFDwQgyJqDHU1wUSgy41gFVZ+7wuHaz
SNAjKP0NEIg0K6rq28FF0qRyQzjKVPzT4DjKOkWr4CE6zDA3ybS1OS1CXlcOY40k
g/rTJbYkVnwDEilxNToqZdZd/8glQLv+fWMzJJd6OlU=
`protect END_PROTECTED
