`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3kUEmZdoOezAyCiTjKSCOPq4u+dOCTPbQJ2oChFZ2b/OWDezpw840GDxAlrqKsdx
/WJjf9G9kz50O8XaHSqw0AtVYdziD3qcq5kRBnyMVGT0gpjYi1bMWOwUO4p1Zpbk
J5a2wE5F5PrWqpw5YrzKhtZenzgD7kNDgkgRzBbAE/NsBuFGvaJ7NH4/F7Swr6Lv
DlnvJOCj+Xc3JFEI+mwisyx2Tz1bJ2yV48aT0PACV7Q8sfOvGsBXVMoQQWFc0urr
gJNOa1pbpXStKINxTKRRg0LiiK1azAuT17P4r076NehVSY1S3Moe3l+ngFukBV2b
OM+JLQ3ONHd2S550BXgjH/siBRp1/N3+76YwiQHYNVoB6wdOqrT2gvkbWqqkPnTM
BRuS1hupovIbihQxuJPp6V8ta8+5h01raTPxBZyMS0Kqz9emyt2CUcWDVNRX0rYe
rwUcYAqBjSTuslEj/9vXzgD8PcGhTAIz607bOJR3R3HXjNJPTArman174mSP4ICv
hV8Kd7qiaIipTSPW9PDEY3xVL0HEt5wbby507ZJp42bGSxiGWFiydwdtrnxGarnT
MfXWItfxAC51nN7TX9ThPCt/a5FLltYmlFcoVmF7UlLbeZx0TQ4lXjas4dSF23Wg
sAkw1ZLcjIL3yXCyy/9E99wARoCtMp+TjXfYkKJYPxHvl+YEGKN0U15ceq2TuSUy
/jgNOkxk7Ow5336RWrGPUb/jqoqt61Nyqs2Tcbo3hgQTMEx+/++19HZAvN5TQ1Oq
TXuVqPScSH0xwLpzi1OpYmckN0al04KsA2iAJW9gZLCwUARqsVpa37qr9xdBGuBe
KmkE/YxYpSFuHp32aIhJXUEGdlDCMRAva0iyjd9UERL5zQwHPvooHu/uAiHiXTMD
Xhd+XwnPatOieE9kwX2gKHGz5kxmVzSprRMLdKaE0K4f32nFl8as2dDnJ6Q5LOuj
0rL3hwW0j9BF4DGlVk15IgvzBYraWM0QyGxHYa23cQpWpG61E6OA8ELlH3zmJ2/6
WZAyihd69JmSuW7wX3i0oTtHFWuN+lZCOTkM1w9/G3Q889otw09x0bH7HptTN3n+
d74IQrExqT5QGFbnJnmwahhsYz5qrzzRScTcDB40SeH9fYLOnVHP1QvYhXFOiHoy
c0kfxLmv15k5waVJ/fe3tryIoAlMR9t63xHEEY24fXUznfJ3urFjdEXsGHVcNLCs
AduCaR+bIYWfgv95sLumZzmZ42hS1zY0Vr9lEpGDyPAKTz55UOdN5IaAC6Pr4PcQ
idRfZmR/Lc8CfmTFGpeDbnMKz1Tfvt9RS2KZ8y1+SSmtuS5c0+1cAGNfJ4pT7pqW
ajwCBJRSIYz4yF8pyR3TLguo0217Nx9y3anqcavJJzXLOTuOGvRmYNHcSEHLbhSu
DR9hz9LmFWYc5db9CfiWbFkUJbzBF2gP7PmUqO53kDEJ54iVqQaWVJNTlVZkrpzt
WMUt1y2VUzpZ1t2hY8Os8LVXBFRWB4Xyz5FFr34oT0A3SyC/vqk/0P/J8i/XkaST
HQDnnCA+/oYbuimCzeRRWEjHM4jPeacLaCJdkkOtV4aZ4L6gOVrZTOC4JW5LlJsy
P7029/WFlSOsHNDC2DqV4DjknYlinyo7zpvWImP0voihNTQZ33HvT7xuH8r5L5L9
8rGQBZynd1pq3hWdLlFYFjMO59rWysa/y63Rq+Hjnr43deUl3rsYtY89gWVE5TNe
hj0e8pjSZMsb+bmsTqKRaEKP8ve3ph/+00MUC4ZGCv7LAZrXg37Z8AoMARDuWkgN
G8PhRZUcNTFx892VclaN3f9PYOqaeh+fBGPp9Bc3Qlhk18MKG3jDS2pvePlCAbhs
qKTgIq3ZLyI4A8zKFw2cmnHMUMPcz/9cmnoFX9c7/RJjd+BwgewiLJd2fMREbHeP
4gnC/SshgFLhqcdMBtQSjqjAL1k2X4QtfAGQX0BBn0yQhmFHekBC9xqwrmJIb0GH
QQRrGpg+AMJD89wPmsChXcgpdhor8UuaTfW0FG9ggjTsEqcI8kscSB0Nw+tA5iNE
j5jszR481ag4etdpiAPsw3K2fWvHNB7bohwH8WUc2I+IymYEZJetuhcvGDlTIPyS
mNftD3Yjcc1oZb2/S2p9eE7WxEHSGSIU0dpgiuMyZp94nJXVohcgvvdhinUfd8fg
cjQQlwZfVhM6K5NC8pwaKi4Gc7SIrjle4A0Rsf2CBOdwWQoHDWLdmJNgUt7u/CDr
IZp/zycKOqAQN/zLgGh7M2NI0L2bl6n2T+QreNHD0oV81/uRkTsqM9k+eHnlH4ml
p2yFAjml4ycWf6+YGhgSRFqFynzzsjtoB25NOZpVuhxqfKqOf0bioSgiG3Yn2qR9
CJoMe4hgop0zQh85RWE+EUs8Ak8WFCYpIBmav80nLdfKptViryw7G2s5R+U3Ra5A
6TddDgxkODEabRAlQC1P5FYq1C8Neld87X2JZsqFxffUa7lsCi9pkcXbLvIoKydG
QvzVn7xWjocFBfRG6tIN3f8sZv8113CX9TPHRj/uI6ibx+0kthzubeO5qKLAaOvG
/y0OZJUo+mxAZbWMvJJIVxmsAxlRF8kUBNFyfG/f8S4TX+xwNvheLYzzqLdf9jNg
3ICkejwioPJ2HekReCouk9e39t/sgkOf7ZqD/wOaSApo4NLPm31j1gxhwqWU0HMh
xdPAF5GTSOiNGLV2MsovFQSE8ZE9u4SEdd5wTU8VhuSg633RFzJtmJZ3liDz5V2c
UHyXqWJEh/MSQpkVTVk6bpnB/9TKUXyBiSvYpygnFrRCw/+sRH5+EDOEvaRxNRYH
4+9Z2b6Ew8KImLKT2XMWSmYtIcUCeWSP/Pc8Ff7MV5h0TjQjVf83GcDZCc68C3ZZ
XRKDABXGnngMPYqhMPBFvEqhlRo1RZinuQ1G0I6MKfKmPdwRtbwsbl6p7AvDj0AK
WsifwDqx/qExSc0vIJ0GV5Q4j5jpG7YGBvOJkJ9Mt/h8sbCn9XIHrqBYt0kq7vJt
g3dmztFtTFOwU3tq0LWVuajID8gzp5wIJMpIbJl8e7Y3UpLX2zm3nhxmKYDdm+y8
dk+g/qaqzDE7tLl5N6gSrZ8k0HATgXAfKFeMA+2Sn/OPPN4C8h4IzUKgEBA98z1C
nGHGq8uX95SOjRXCrAbAgirfdayTHM4VShswSByf3o6glcuXvY6zzjJmZCzrscPR
e682jhN0qC7g8HGXHi2hm6I3svaypClL7W6gZBm0QX61h9SVYrCPbUwhuGGA1Pje
Ni38lrBv7AvwfUeAo2L3tl99R3hqGylFDL7/b02iwycE+B86ALW4PmIviAjptn71
OqmKlku9ih3IKl9z4tNjK8Ao0WrMikE8BI4rh59GoHvRlvmjRtp0LrHrNubiZiN6
3hTAwysT8jYl+9+Bq1LEAQDgosQ3lR0gNY5WG65thckuBd2qDIDu3qJb8FB4jGdg
W1O116058Lg9IqXwnaT3KqvCfV6n7NoruPrkin34wL+aSuf2IXu5qkP+mI+2vQSc
WRJUz/CQWboJEqWvp/W1d//V7TJa8BtUxFAKlnZ9eZA8z31t78R80/WTwMRQDCZj
M1RL7+4yD84Nkb9SNVH7gfbEXmRnFYJ8VUtws3fkH0exvVJ928i3Vceid5yrFCB5
K8IN2ZVmTBUYh2B+LeMiDJCQjz69gkNbVqwqwDhUjVYGWqh7Qzpt6lGQ6ErFnCSi
T8TVnJjn1KF5Qx0rL2i1Ipt9/w3ZkdBkfATC66FJ/HCNumO+W685td5MLs4F3mfN
oYqJ6x6uJnClkZZEIgj8EQag54lXDIKY9FnKL22WF71CaP3tkfystZk/NRgwGp2w
fwp1k9oUwzGnf/GUS3pDloN5LiTLVuGD/bJqSiM2YX4EU2fr83G+9896AjFuXwh6
wUEplDdMvdWgpPQphz02ta3N3KN0+g1WGgCt3ddFYesqnFBLrf58hL0RsGAb+av8
moMYfMfT9HEkvf0ru5dZpsTZfgKDqM+1FBHz4nLwFAiZ5xXHtQJV5QEd14fzXECO
lztqB0GOMztmOT+ubSs8NWduYiGiTPtUi/Q7oXX5HMxCozpk+/QKKyo5AP+MP1bL
1y/bb0hPg3X77mtG7qj1K+vhxIiFoIgQcHbnP2h00MRDuTXyBVqWObHRwPSQpUsd
zHQeWwU1TtiDkwECadQlgEkldCl87OmDSRONxmaSqUK66un6DC6rK9Zay5tovydN
u2BNZcGNrmtzHPM9mmEphgpIH+s4o9rYrqJN3YvJ+6rb44bXj7XCY+xk8g0W60bb
48pzXZfztcjh2lRVioSlEZiNuQl7iS4NW9JGL+MmwPuqjpx+sSuJHWxxz+GNfY1n
WHZZD5E149P3HcN/4ZxiNyiNE5lSsM+FmwzJVD/LBcw2zW03+J5wbfphrArzaJRO
YlVZFlEwXIRq/7aPqVGextrYRDDL/igJwPcuJSE8/NI82WfIHUckYzJ66BcJVP24
xZb1k0m3eoXBBzjnp1b9YONM9ua2VrkWMBsQQq4vKY6u2kBEFBLGXVnJp6yV/VnD
VtUVmLSiU8Kyh9IW72chj2+A+/TaCL0QvToVYOaHPSS2PL3FStzQ42FTM65wflog
KnyLzYEkYgNWBvCf0U9EHciLUdJAAiPibIx0gDtoKxj42Pq0JpBJLubtS0wCu5ia
IKLLkAUx/VOsvtOCfkJV6r4GlNnNTWwcC07J6qJ1nkNIoum67UqcmH7miaK1KZOX
lGiAmUjhGJHgb9sYmyvC5nzxH+eGd+Nw8rzG5cMbdhOWVryLcYFhve++0czqSeZj
xSvKfAr5+f8yb6U5oJFLIIJlyHtPg46UISCIZOc4DMx7SVqlnZpCyqo2ZAIwwkHM
xJDYCijUsGSxX/cQsVra+VWwEBhjiWyDYf9I9DOAgEhc2fxKBV6uoCE4D40wjrlI
B7xbeKxhyaPhwBnqa+Z7wSmZaYCa5MXu+nEL8ENg5Ezrk/F+s0Qu03hsUV7vjGRL
3aKp2t12ZOWmKh1XOo7c2ys2Jp0F6lf8W3ASE2UXyr7vHhOKpIXlQnvYViJcAnsy
+Wogh4VA0akyUUAdgNkW0WmHbwBjixm1l17Z4o/rcyEGJhYxZI9StuxCSlpuSsfI
+tPa4c6jc5sqqRbdZuPERPJ4vCCNsD2/hcbCM9OZ0eIYZjwu4aHR1DcvFJJdQpcr
Avg9hOsg49UKMgfVk+VGmLYZ7gc5VrNPZx+ZDC3OHPnJHb0X/clueun886vZq1VV
pkPBYL2Bl0bSU6yRhacfxrv9+0h49AjMA9FG3krATC/qKDN2lYgTUKRu5U+uaLr/
l7yBhWY+3q4omYhjxGdWDOay4OoNjlu46ZY4sd4wsHwdpT+pseQUrvCiD4hSFCHe
3AvxbIj4RYG3sHWVZZPKGFwcd49duw9Qo8ytwywUHTf9GFeLFRlQj0vxXhlmOGX+
IqTsP1I7ty9TyjzLsK4n0A==
`protect END_PROTECTED
