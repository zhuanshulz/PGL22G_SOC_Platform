`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VTsm8osy5ObEl97eB3Fw4879htqQ9mFBT+xVtVMaH/EWG6ic69Fmvo4s2o+QeJM4
S9VC4DilViBqGr4xjInVeT06yHSyMqyAASmaAEzS5PBRFruPRH6vr8qiyw3RNm2q
bDKZ7SWQNR9hMtDjiq6yhr0Q5K7ZDRGFqzkhn4c3j1nANFaShY9i8dWXsTQ4kGm3
pUh9H73enjDowHmt5xYIq0sJvnen93fumVSk7yz/4FGqfMeKqsOtrQIFV+2OrMdk
V1ABpwLivQcygRRrbKYK+6SW8YltMsRLvhWwFUMameV86exeEpUlFVSioAqtlGLI
MrF6ezfWM2k6QdbPmcLbBJLIOSxkHvXs/pCf3I444mQynnAWxkwzSOFU5KmVu710
IxfCCMo/q4+Zsxq1TCrKdeg7BrVWzrEdvfZl2HyumGOUFhan7xLAE0wHy7GiPFns
oAeI6LZQPPItWNBkg4HZd6ZovTHjsUzYubtjUCs8JIgkXWY14iQcQRTaTdbempXH
1EA91SPLDDPgji93Wa8o4+bAvfb3jyd5K2Pt+06RxwBPffxq+HpRyppCxpIbV6yz
0J2ABVZ96516rIiWefEImqQ11ylktGsHq8JDxHZi3+OWjgUQguPqp57mHFiDJZTp
TyQa+gXoH5wR2HNYrn4akU0t41SR6SWD+LhFX/E8BJJdg3tKElwTs2c+B0vGJ1Pt
Fpn4q8Oyhsc2EbYrM1Ty0QiNCL4mVe7aKcKJ/idki2K3LKd4kef8jRdESVJ3kHKF
7x+fAJ3VadvxQiC2K5l/jk3wqJGmOKl98G38KxLnDLDdUIZNmu4yAXgd/12EtDKA
RLHTUPsQm/tVm46kB911HIl2ANO2Lp3GUKduwVWaFIEFaue3co30fHjqVGtcl1SB
auxN9pueGRUOM5lUzh0Yjg01xoklK9RnN4ZXoeuoXZKoKL5OvXRLDUZwlaL/AnNg
sIhtXZ9h+MF/KIL58H3GNHpXryQV8K8e2NN9xfB/6ghoNAlmsOqnUMAgYMAG/6zO
E1+2Iu/4n1p7YZUKvxRiCOXFlK3PMgGx17U0n/pnZY0kmLy2Ok2oV6iGDly6fj/o
`protect END_PROTECTED
