`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eG87Tx8o/It3vrQUgczr4ziEwSDyGeMWXq/XgZ4aA67Rz4MKhg2vPncCq/X7nrD/
rQmYx74KoFMWRTJs/gqdZnR/UZ7bMb8YSZzVjxwpUyZic1jQ5Epc4hIix1WYMKn+
i15LWlLQ83cjncuQ6WplkCd3Ej8cJnn3JBuJvypT3zpwBlFuhPIT45/i2WhTIhjI
G2dkjzXHVAxXTgENyu0m1MnIZ0FNvPNpXQDaIaiOYCn0g0iO2Y1Wdd5NJgiFwbfW
pmmvxnCDVssXibWFgPTfOOXistVZrDAZb8DkJU+NBx54aprUOSezBlzkyH9/MEno
8QvQ0EPp2uG17wfWUjgP8vofatCas8tLeOt//BCqI3JyieB7WaJfGwI1T71lWPx/
lmgRw+wO6TD3aAel/zOvXUiBd92f0O2wb8RAENLIkB73nEyOrYckEA9SDozIoZtB
Ri/dGmNkVIH16sCH5+1CtPblMu1GL0tgHK8xOjQOqGFMChVAInkZ/jY0vKk/Lik+
vhvrarYbWHaVcsqzkHsJtUlWV+yI6FIAIe/ZzwxZQ9TlV/1yUUW4iQj0kI748pIp
B4TE23y5FKBQCKatGmyo9mq7afmycHoQLHORPbfs+sIwjRd3wE/g9OrYei03ARao
DoUAJNp6P69KOWP2D7KwTP/WejjVG1pGdDmEUbsQX6i74Gj1myhnhsFEvXKixDNC
qFnAhRhl62jt72CvKmnUSTM1nHNeJSYz61xEf3t4+QljTcjTz5xYdJuMflpCQh5C
`protect END_PROTECTED
