`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eiEMCulV+lIrUUg5QfnGvu65vRTmQY/f7OJ0v7rjYpuwXTZNutVMWvTZjs/Ru2Di
u/q0ALALQaYIPf1e5ZOw/RCsPrFD2HsDBHyRz/ETyNFZaObLvfuPZ2xN0k/FgaKj
JJ+3NtEh3vJZqHDh2lGoadgZNlbZi4rBvPzFLwBlAnI+askJOYhLBgSN01A+Lx0Q
ryuAIdhQXt4vJg9I88RWuC1t8RdsesGIHyX9iNcO4nDuiCuaM/XIQI6RvIfn0PBp
kbmikomOJbwILReM66AjwCkKoZNgha1ahjP2oZ0IyjtYCmlhin0USpacW4d3ExvG
YEWFy5WRsoUDMnpwC+YEwDJ4+8Tj9Fg32NuVCf8ryPyOr6ZrrszMc3rFIUR+Aleg
1p0PKrjnN9RRVSjO/5Jq0XHmQVpECaDVmiTTBLpczLUaLemjY4sicnHP+CPkbF21
4UAFPiP2y7qVkCOB9UEp7CrdlpFV0Sh5g5I/99j8QmvMRTXHhHU4k44gpyhZCZBZ
tloJ53sbghqVQBORGaTNpFR5u/G9Zs15GV8XwyWHnTqPE/zx0JCws4UHM+PI4qfa
QUNf/I9JoVP5gsYvzJewCf6eOdOIQUOnuZ72t9wP/YU0+qMo6/gSqzLCbYinDwL1
NCOwKJixyjWZj595kaqiJ0+HnoZWClWY4hnAM1AgQ9dR7jPeOnxT/wlpofpKQG5+
lSczj+xNXFpANlOiR7DNBvjSgSLsNWeCybtxQ24dnPip08BirbX/BNznbPCxb5kx
B46nDyXZV400XnCFBBvgthWrTW3Qkljt+hDr1it5UoESKCaUF4l+s+fpjnkrce7C
Yk78b2Ek5acFzsWdUz0GuRIl0FRjCODy3QQ8QEKOd8QMhqyqY0EtG+EAArC5issy
AvIR0OWfoslQcpuog20gB3NiyLQ0pW1KIdAaRxmV2e3AM7YUt6CW7cc1ru9YQWe9
4LbQo00mzOrEvqPJJlfbErEsAPye3YAwm5QFuC0o03k5G4wGfzUjKVwzpP9X8GOn
E/gGQ4r4NI1rMOueiGrPv1LCMumSxhcAlKf3NzL1cz0fVWT3WEUI84d6hSq4UDOw
1k8l5ZCxxriJCKmPzlItU8kiHZnHyJmYivFZhR8XX7h+oJCosjLhQjw5BZnT59kW
hvkvY71oYxFJJStgXMe+MgHlDALC53cZWdfaIwjdFrp1l1qrJ4/Eq0dPiEV0sA67
DoZmIjy3ZvkBte/7aAAdNg==
`protect END_PROTECTED
