`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PqZmlF9x3vqSEhx1D/Z8ZTawL+4m2kjvfyp/oKFG4KAWYNJnTIQmQLA0wxX5ngvF
5yOqQDg9twdQZWmbISXGo0AtuhHi7ohicyeu8FukWZtwsVWhQ6U1hFNeu0yJumh1
tAb7jnaAqF210J0Sy8TMMlM+QbyewJT2NF+9W8qDof8Ee+L3k++egoXKqgWdoNbi
jMBEclf/kEAsxA0tWWaGvHwt7am3OKW9MrEZi7m7gMjXXO7MGvf4WNwUtJZfGnOb
LcVHKeZRq2tcAtHHe6H2ST6MyAW2meRUEYB/gh7e5dJTuRGEVqMZRvqVMNdZakTL
iIV1roB/KFB2ECtOc/SUO+bijbm5frZ8ZrcfycaVI2Yd3grsim3caQ774LvdOHLS
FRXavbZlVAyIW+V4+5DDSa1eDe5fEZSaj5oVkH5LEIfTbv4UjbXKK3hAaoyIxdMX
jhD6f587xxwN9TRa6UmP9QIwQPoUmDRpXjnYTDy5aqNaTheKHndwAMoAwVooL6qE
3EQAFyinUJKEMNXv7GJzedJ8tn4lt0XTPCJ20m9AuHLRMnTSjkhwwwMLiXzY8Vxv
WYRZEpSMtCA+rf8xmSjC1W5GSJVMw8tSdOT+IyzS93FQq59GqNS/aBp0dEMaAIG9
6jZO6eFGEcExvx+X4DkKavqmOHeAWfuPvMiGMf/rk744w3e2NQ1AVus28w91xUDG
Yhq1J9iQEbfF3ZwIn/VS7300SXMjnextSuCaD0H6yfo09cxs5pIg6m/ykN3CncY4
Z95lWjLcSXC8mQ4Bmx5rhX7JUfLmvf3baLQEdH3PcGDgZkyBzITKlVAMMlVfFjW3
3qt+V2Md+XEYjfUdXi8KPNTp9z9wUcPdzMArC7nhBT9YKZvoGWZQeQZAGmVVakrY
dOd6qmoUEmQh441RTmjzUX1yUoJpRJDIvLxM1ceclY3zCiKUQbNKVeC6GkX7kWBm
pC9jj8FFu2DJ/RjaRzzI0d6Z5aNP6/LeSKPIlZI8EIpg8NJMwd5PhUdGLCbmAQgW
Wu897L7PayyxI177GXUOsTWCWA5MHi/WB1L1JU8EpWRYrRmPMAwz4ODjuzxoHAHZ
zkkiud+kkLl8FaDi67FIArJedVUc/P/TEkZ8Xyf8Kf65SYxCA7JJEJGfY5NM4M4S
Cv4iu++YEEsLYfYKjatfNToNcAv2+vZQU8wDF34TIv7YFnqXXMpQmPPxjJ5vezPw
pKxRXBUWZtDHddHrAOSO2sFkO4eH9Q9b9R3DoslrdDoRgwiOT67VK9BQ7Glk/l+D
6frH0kCx2Plv+EMOb94oBgJU2a2tB6F9cA3Ijxm+jkAhUaYTte1e5Rf7gI7Sq88C
hX7TYSidTVcKnbHYfP7L1l1RDk3ekd+7jikNTcnGGWHZxZ5OAjE9yIEmGRX5VJ5T
Z0IKio91PgewnsF6hiFDgB6dcCy3oqdCi7J4DwpBScagW+G746kF5TU/lA7Tss4F
3xbnseFpclaJMEK87hwAokObii0oAvSMgI91fur08qPzza8AuzqH1NDFu/Gt2XwA
A78WmWnLT6Qnih7Sd11Qsp0iRK3XRZQlJe3thJtHYqC245OLTs5XFyvHFGIfoM7I
0Ngtsf7fy6a6Ag+i6QRVC0ufFxMPY14w11jMSjCoC4xbXPOMAGJOnfIWEJSeG9kp
NrlX31fQS1McZeS5JqeLedy1K0+p/3bXtOW/x4/TphYDy7fqeOdWxjRNzcfZVDP8
4Lves/gxaVoL5+7z0RA2gI7Kyovb+Z+CY5czj+/8reJeEz0KTVrVoFAJrkzVZtIv
1dz0T49DwGfrrz6jskd944JMCi6id+tT88pAGJap/4RfV77V+y5TtN7CWxlM30i7
eagCNMiPFk3xZ/PqOy2aNEtiRIZn4u3B/uebJUg9JloSlQE9YO/ecza2sQPMOy2p
DjQ5XQsek5vKYKzu/95ezG3NBUzOuS2zhlS46Ft5ryfRzN1gsk+NwVFmytULK0DJ
8KnDJkF2DZBfju8m4rbsVkmRBQhuYaoXP3FEYlGm71sDll4lfYpksnB1QUhxOLkt
5sR0tf58f6Aqc4qqUg3ZsN8gbaSu/iyNNdzKwfIOhziXUPXKLFEqgSaBgvOQrEVM
Y+wYfbViM2oM9rlmx8vFjBgtsnkT9BvErJQcmL5LLtEwjxKutmjyzHwBBSiW2kWy
DxvQ8YJ1it/SkJ5gzlS2WMPAZTp0TptQG73QFd4i/AQ=
`protect END_PROTECTED
