`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qsxh45OJ9YsDC0Lh1QdQeq5PNJ8aKqV6LUxn+7WVSV6Y6gbJEEdXuGgJPZ0QVdHK
PbxB62W9+Msa7rlBdzBfesVk05O8MamkoJej/WuGccsUEuRG3irXxtDkl7c8Oi3o
FhJEX09hqZG34pnctYA+AewGOcgpGLgfys3h7KP18fAAZbgBK3qKYPiPQJ9tAY/O
GF1+GsGtDEA8p53LhrY1t6hO/OS0js2h41hYC3K6foaE6gWyywyCfwaQqc9hHac+
lo984PjO5Ts14CombOvjR2s++v10ehIENYTbp2Ca2OIp3iyi0bJNephTwljgPNut
bcageYWxNjpPwhI/qyfHQO3Ywk6AAp8fVNTNnnKx3kunx/7pYR/BaKtNcFryTEf1
Ety0xbQ3Z47U8MqkShORu9WNuakCA0/oUa4e6t0u3b7jaerzZGg7XKt6LMWsrTV8
qmNdW7JKIaYGGJlHxcTgRhPEeByaPnJi8EhW2+TlYxMCW2XJUcyoX1n4ASRizbWN
Ce5EpwrQ5N2jQMUe94Vukrbh3IiuzBqxfunDWELlQp6myYj3Xu4rmFmgmZTjbvAz
iFLyoO6XLKcnvQi5XlbDCyWTG37B7q04s0DI0CRoe4bXpfia4TNUPlVC+IiPQsbX
`protect END_PROTECTED
