`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XnpxWej9oo1xRsKdGs3C1ycYWtfCtAxzhzHPhqTONNvDgoUJo1rc6PNochp8jORI
pOc5X6D6N78B3wWz50pFp4IoTS7FLakMFty091eSX1X4QzbFKYSvUyV0VAaLgo1C
YU2I7W0xOJAKFGcrR44J4SoVZjkQprQUTT2aS4dHtPLnwNCX5XOGP8JN3izx97pY
E3iGFk3XFbZdnSoFOWSi/RLL9NKvP8+WmGFCKJJUL+o3tU9egJeN27OSTUUiGb2s
QxLrGlxpjOYCFKJh7uYZUCollsfCEfnl52FQk+yus/kCAUoR9TXR/qy3eNpqw86q
uDgHFeSOoiCcNppkcqVJMg3sjRYsghn+jnZ0mZQGCvVezngJa6BzVtFu/xv+C4xi
3bDwsJT0f9dzr6/4L937T5ir4xXnwc0vqb+xg8eNEcLfzyngN09oxTAJ2cSZOhQF
zas7XmFnGaB2xngmp8NhunjydN3ajkaZ7MDMAv7WQPyfmkSdU3czA3Py3YlEVmUL
GLtXZQB5stoKfekPttq8+euFkozycX9jrTG70Md0oCtxcruZbXsxr534Ba2ffPsy
XGgA65IL6UiocJZoplks14x2BmnzH0aLrr5JFYry3VyX/SP9qqiXuQ7tsXJESVji
iYsv833nYe6bxwa7w78kvLqE5Gx6Ck0g3mz6BOcIGr6z8gCaf6r6xa11C/Egh7gT
Crdqxr8esB1bi3hcIWwbgMgZV7sjAjQazk+850KB5OtYmnYlch5pWgR17487gk8x
Ik4E87e8H3gpiMl1iZS0aBPsXsphICUIPQrcfdOW/WxzO+QXCq/xgL1VuwpdSTnM
BviQFEmaxoQZotE5zNBlSSOA8+oVAJbu6D1yr9/U84rzb7huu94kNQe7mdpoZBgy
X6eT0bi73NgmEiqfzo9vKFKwpQxQ0jCUM7ZMqt8qavS+cp/mPJ/MbBAkEKL4rSJw
f9uYJqca/wG6zG5PDcyoDDmqNvK1/HoDksnGdAIOdUmtpkfvSKsaPcMJiymaBUll
UH7P/TBhSlA/O2OEQNBIs2Qa2H6MFGjxu33F/4YSGxpUpTrcEq/BH53E11DkMc1e
Xn95CODhH8A4mR9V6pegeUXDrUoYRLjfEp3j2r5Z0DF5VFas0j9mLWrO0xbO/Cfi
RUikb/YqbPVPIWMzoLU7K3FnNjuaNtipjRiCTEbKLyGJ7I96DwvsyzRYqiaFeqQg
TgSs+eeWj7jp4VyDFx4jx+wRVCUA8GdMQ82H7E8BPRicWQwa/IZreGcwnd4EbvGi
Q35ifjhHBepBd6UQVZt9pLfGyT/JcKiBregZ9W63E353RLY+1JORviKJtWJLzSZB
Up6BrLn8a7hxEKtp3f4cI0x0FtxuBSuqXHbcxGfh7nZzp8xxYbTEwZuqgpaYX2Lu
cIbi/KAF25oXE1iL7hh625qwTANDsAfMge98WKyAUorMIRnU3ILDWvECHHNKfX8c
BHUFZZTYLYhu1fnyYlkjhf/zwUh8CXzIISg1BhB9GxE82xvXQJQAplmh9bFaU3RI
qIP8LOu++FE6doExmkrq5H6rkUOVk0Aa8skVHEwJ0lbCNZmyMEemlJTLxnhAVQcz
85+hPdkmzNAy8Q+njkTIY6b6jdjWdNRcSxgnMu1xOZHjyZ4eBUO+tQYb1Vr9xCBP
H3Qh1aGoY+IjmGFxDKF5+f0ElbSGae1emcR4couAoUdBtXyMzj84oIDbmPdjMep3
77OA9TO/NGPN5fnV+wJUSFK9K2zX0RktldK4YcsVolExFerrY0FGD4rgnJ9KDueR
rOAJ7BkokpvlEMaJIsf/2JILy47rkXkWdV343k1wGv1zwpBIOGD/6czEzL9av/EC
Qb+Xilsw7Z/ds8NbUNrTuJoC23X5BOegCcB1+4ypOa95CT96iszarL42xTddXLse
HNyHK603IywX9lZbi4EGI8I2V9pKWKbLCcHL759+cSVyQ1q6juxxP0ePGLeFOKdn
DtRC3Kte8r1gHgfDWMavhTWqxbXwQM6B3hQcAx6tj5VzeultJ41E2fuLO++6XSAM
Gkf8zl/DhMJiB9z12fG3Y623pAvBdoZjry5UBtOWkkAIIyV8bycMoXuIeu2qz7+F
NB6BL9KeC1+ETxdEyXk9tB97n3I2cEOTog7F3PAk7eDea08mdneVZJ7ob1zMTRjo
6/P9pM5gwnNWnqVzS8W7Nd/cSsg194c48W0G0J+5n2zfC5QOILgl7nBH0n2ITRiI
E6psjB3N943HF3FGk+U90eTQ1zLyq9HZl5QBkSEaltyh1kMRVYi+vR3HpCHA1xWn
fq7P3D2YyJN5dbgWLc8HFBp3KKY90gz7cJRZNU/mnZpLgKC97Ja9xl1iPUEsy46P
Q+d04twxkqdKw6GREuYjuD0gb5au7uVYNpx83xJpN2h1qEZ6P8zJ79BQ+WxjhBKW
+VrXKh5yiUgq8Q24uEe+dqMyTggyYZ879T4fH4k5srGuL7i3PUlWApIuZKHbZ8gO
uGXz/Mmp88PE4bCkmhCFB45516gnyQ+gbXESEGU3j2Lda5Bj9KcgyiKwD+1Pi1Hd
238fuce1Hq7VcMnPksdjbMH1bTuoF3yeT00XfI8tnjzUVrpYkCc2cdh0MetFRy01
RROgVs1BBi/TavPeHmneVjjyx8c9U4mUS0xwDYeyDkaTxWJPlou1uok52kXaieFj
kwt+ziQFuJZ4QB9ema3bvFJjha4YiBBHHIpgTP6uTdmzA66M085WMXUDA9Z8RCWw
pfc14sNSf4OrkKGIcecYGPTuD+7alW2ydCZZuPQ1kG+Xap7lVMr/K+AFlXlMuXYb
dzsDJNUs3nMFyjoj5kaEYHwzcEE3K1RZIm0Mos+FWBmE3IcH1Cg13IsPaUbWNPAs
mjUdOjWmH93LC7q91fCpUzp1BZOdStGSowzQmrjXuk0lgLFvfCPGfaz3Fi66wuIT
UgifNKs+bCgZOxNW0KFb0SNMtX4M+/tWazR145Wm7UXHViL+TpS5+4XIjns6Cbt0
4YZmypREGqT2Hkv2Fgveeq1Lp1mwBiJL9WVKv9Vm3209Ph6qWs8yT+Wyfv8HIihO
xOAL5kg1q5nhFswVafzfaAvCZIPMx0SwKh4aSrL26sdhtX5zUsNinrvTgfvROybg
PRpnzUY1iBO40yifGj+7WoguyWFo81Zq6KdM11tyfsPUIbkTVd0dcXY48N3e2FoF
5H7heCfT8apmmDnRqeBa59Z6T45bZFs9Y6IAQNeW3VqQ88b2RfADKuPh0/VQLrFv
YVKvfnDEMuWb7m+ZN4SfAAQTZWhf7trfGZs/8teKNtSA0OCxfQCryC16dPOWITJg
CII2T02OpCUHowvJmVn0SIulVkAPQyCjO0eeAMA2CssCZelX6twNI9OrfVtw20fa
XU7niMvZEWA/2G+EFDRVNQaDlOhy6MAoJt0kuxwse4GgVeG9ykOCIbAl6kyDj25C
CHzYwVq20Go+ZUXK+pvqBaWFmVP5QRyhwq9IKtzooqmOJ2HAXTb9nyAhnSsfmPV4
2ioNtEK+2zqDv5nsLMX7k37pk8wnO4rj+HxqUhJFOSSidKkmW08tdFDLRI4CUtGm
o4L8TKUpvLiEyvJqnIVAPjOB+Ygbszy9H3lkQ/PCHwMdzTr6VtO5JDirUJKZfYKZ
viH7nExTJJX5MJ/6ynBTu7pj5xB7dX6CWVnkZEkW+kEg6LcRSv7fFNzTjiaa2Ndj
QqeCDCL4W2S6YeYdF42KtOuQp7WHxk0wYu88f0ci/j1eZnjnIEsoMoD2DXoNTrR/
pTF482QzjJWFbXW8CnhHanY6fL8xNQgSQLPDNyhUGVqRdVpquZAc9ASSC9XaNbIj
v2o2Jg/NTj0qprmEgz1sOafWdvcIa3DoVJDcpzt4nhK8w8HM7qyC87QnWDmofctj
ZYyxGsLY8nrxAQmI5PMXqmn2lRMF4F9D1q3LpKmBsvA9kKyBWhTN2nA3orncJHAb
Zsuv117bpp3Lr9LH/rD7PCRlcqDQlG4offWzLg5/8Tr/NQJpN+RKVxdDQ9/94NPl
a0HXgIEOZrkYdT0ZwxSZmVAqJ/vZQ1dpmA1C/Bl5mrxgPfE48/SrRcVfSKzpX+F4
fWhuKcZLJ2T7bgjjXBBpl74pdCWBlmPjHwTYBbUnU1i3TJ1UFw8cwYo4Vtvf74BB
5GmqBESbGTdIAJqRwf012eyjudDww34AZ1cdUTN8pZyNUXjsmFbnWKq0CFgEXJ25
Co8y1dsJYVEodoPyMIsz4WbBdjlveDhLF/hQXs7VWnNJzLqAREnbcDj0d2IcDLIO
orgHX48lXqdc26TeHSLrXZtQsMim17y6o28tOpafOSphCj2/S3NsGH4LrEuSSje7
QR8CqZeVC5firRqpLS7dLA5IA60P6VT80Uhl9aVoSdmyh/BxhFheK+H7LiwhP8qo
ipAOB2LhILaLN2g/jwWiaSV7mkgmCyFWE0BdjCz68fWOWtMWxldba1HEojxmbEo5
zFV7z0MRHnUHWqsHIGs3Sh0c3jKxN2zOjqPJws9l1AHIFDdEETcmt99h0+ZfyjHl
OqFEA63XL/C/9VJJtvAtjLz/j7FZHnhk2N3PRi5wXoUHhqnMAJ+WBeNRaSh9MvcB
ASvFbfGvydOBkXWLIhaqCsfzHkgOFzNW4Hno35CVKvMxZNS6ejfehWLMGbmTi8ah
cK2zSp9Gy6SzKybGrkw3/cyM0HC/sg76/2sOm9/DAUvjACNNradJJ2xpvS1wkaQY
HHM6vGY1jcf8pDtrEkjxuR7Nh71bRxT186TNXYaSeCzT8vH1XjzEir6X8VM4iygw
e3jpZg6mSk2Cc5RM7MGGNRmxsvOcRKQKnEkZ72sibzCyurCzuvfm4Cd9qiZe8rKZ
aMGuBLhCNj8WNIWOXfBtvnPEImlPCpmjumNh9ReUeKpw515s1BoCxZy1MJlVfIsq
aHzoqk8xqEBIJXLo88nSkFphvL6nBvmddY0tH2V80yH0lUyOH6WriMl9SY/1DpEr
4EfrMQ6SCS7JvDO0h6UVqCK0waym3Gnf7rBPU8DcaCmcsVMTrNL+JybTpJq8g57Q
Dn5icPQb7oc1lbwOK+iErDbQzQR0HIwmYr+1oOB/5z13dQLlh+tq/KQ2/t3iZIby
5bGKMstwglQBycE8V8XSBs3CE1W9pA1BuFl+7Sl4MK3UBjpbOxf7cC/SXOs9rPKR
kq1gSP4YOvCcADE8DOslzt7vciaMTAX0ap0wz+hD+LXs38d8TglHXn5C5gPW3+1o
J8axkwvl6ua6jVfzjl52sZ9uuWDYz0LVLrXEo0U/ieqlxxKmY9H43r9u7IcYgEvV
eO1Tcroo0FO5/SbpubD6KbkFB7jxtwvFD5O3yeYQsHuRJ1eMZfcid2xw0y4ItLfx
CKW3hUEN6F9u+EVWp3z7R4lfFZiKA915A+G3Cn13Z8nEx5prBur1mTQiw+naUJnR
6XUnCpEezeVWOcM0VBoPqjqytASUk+sOxakGLZYCThqf6d8Tkd9gZUroSrLyHBnA
TFowT3emWWfaYESdYeRs+16ivVHT8RKIbTYK4V7d1CIXfMN4iCFLflTz1ufMApwt
qRGOI3kB1b5OpA57v+22dNbAFq+2bs/OaubpJcs4ljgVQv32aD57XVtuNDgFpze0
tgeym2tAj5QzXfQW61M/C9nwnOE8NTxOeCKg8w9AgVA/DaF4GupwW1LRAKVuBGJC
Eg0kjSHatvy3jTWCEIWNtTGYrADoBSf0SdDhrX7+cKxmoxHwLvtqdWquuPOySsan
6hrISMxPtDUeyHYXOJMk5nIf/ZOsjVUfjrPzCarljgpMd0XSq4aSrGuxy4uZh2FA
xO6nLCnZtQP/iGtNfaWl5VInExUFPPS6alGjGD3s2bZg+EeQPJip6bF6M3rd4E/d
sZNBh4qvij1hzL6kSOewviYJcr060dVSIcDwQcb+sGFYUyhbpZ9TkiKhQT7OGJ5w
0cwxaqcPlqVMguKTaWrWEgSDubdeka3LCb5VVrwPPydLRZPSkR4XCbu1zCkmvkg1
42/WmVzSeLP+cLRB1MmA4yigRIf2L+zBY5AVq/fwrnjPHJKelWp9/X2YtuMBjDDN
9880Ln+y4DxHiyRfmDlGwoxqj89MuKy8i2K0zYMz+MW4HyLCzYw1yDUDu+5ea9zT
S5mcxqDavZxKUWcaOS3x/d+AJbmKjoDE0U3Y3Ic5y/qKpmqmBlIWHev+PQ+YkcuP
VFKzFd2Ql5fnsfhVu+PZ7kyM3Fq26fu9Crccq5TVo8Z1YYs4csgKU1Gg/3jPiiBh
Zy/b0c11Nv78X4QTrTbQao2fhS6EC0f+ilYFHLb82ZNSDKv63xBGLopF4tKlNzoT
PolkMDvMQynxPRT+BlpxffME6i5FBGaKg4f7m5pI/2jeFPqFRK0uR2lR5/iCu3PB
/VIQvlNLOVLdN9NA97fP6ZVpVKJY4tXM9D6Pj+yqPQGBn+eKgbMSPY9pxTqtkXmq
A2E0wmHB61cBgkHerWNywAVufWknJZCDHfVSOuXOVClEe2GZE+k6XGzMiWhtTJgr
3Smmx3qajBAYzFD71zZU4MYW83NOwhJ5UqAgb7JHMbTBNbNsuEh8an9xjpB+DFXY
d9jhVTvG5qy8yKdIjSpowcSJNKoBQSsKQoHxQixPs8RXU4nGOCi9XPu82lh5pSeU
1kEbaMUjIqHfRSQ2pkDS8GXcEMbYi/mDAx8f2jG0PGph4w1lmA114JVm/dkqL1Be
i2FqRB6UGDqYawBpeJvGtx4wacTKsVNdFUYnaW4NwJKEIZanHtdlMVBaeZT7+a1t
oR/GddNHOsoGDlymTZl9R0QMnm2+S5q9vobotn7p1EJX92WdcaaZJeTm23XgRgWd
ninewnvIoAwFZvmDRMplfALIVBhYu26klEoBMaMH3+uhhihda4IvTuWuozFesupc
kuwISJxxp6non6KGcTTdUUVtZFF48xiNK54Xcj8pC8vXeuxK6OloMXxw0sUzpYd9
8ockqla8L1dQMq8uUsjmYS7fX1FoGQ9awYZ1O0QtTHA=
`protect END_PROTECTED
