`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w3IxSBBjmPfnLzRcCdOIS9rZr74LA1gjVS8LetxpxoEprb7I5IANeM6hXxzglqNC
+MAzKfGWBr3ixjnDbeGtdyQ6dNBkcGSwnciXfm9SgeqjXIFS/p0nIce/JdiFdOpv
WVnA4noc3Xw8ZoRzgp345RW7PW57Q81c2LOO4Ilu2dzaVAdaHYjGR5inT7pZgnKc
dnDDV3V3qnbaJ9vJzPSOEGAEaHIdBAEaYJoEVb8nIywkVQX8RwB9XdlkAE0t3m95
G+lwUMU9rEr9OpnYco07V8AflQpvrF4YCu7umdVcdDES6csw3XuCc5PddP6IjdYe
NsGRpfJ9Jxhu4gI7f9S87McY7VtXm1KEytyXlaF73d3QdC3A7SBAmFKPOO9XQop6
LbMoNKv6yYnCJL6M8Kf6smrIwLXnhgA8lWJmWvgrPSYl9FHs1ncBS51oTTjIHa98
xRM/Q/abUOEU6+tV3ehnye2ND+x4dtIf6yIyu+f5OzQfKCHXfdDBt5hTvezQPNt4
hq7XgEv0x/7aqCBz0l2r3K3tyhU5bL3A5wa8ZZqKASlYbUL5cn5+vgGmHLBsO2qD
HuLZN6781UTMddGfafTnaWcRq2Wen08Yz1Ym4B76NTWAJPLN+822Wl08G3NECzec
TPlC8X+UwQb8nl5+Zs1FbWJjPSVOKGESK+V6P3iuF8HhI9SoHW13hW+XzFLyyYU4
z8o1H2UBxVUS3csN4oft/3cZwFIFlYsX0c0gI5/YMgnQZCqaOqU5bDav5/J4OSSA
R7K63CGfQB2varhcU0rQzXkKsr7Xxx3HrqbqCo69sghQJxlsF+SlYBW/8GXm0Lly
v+ekKGXkH9cRak1w4cKpzQ9II51AFxlZPv9/PDf472gXUfs8FXiUN+71M57XtIHL
MQyDBFZXC7eUr6lCvKJ6NXL33AAUXY22xW9FC49Z/zzdozZ6hAZoLqDw/fwbQmYX
d2ovLC3AyHSV3Uh/00Iz0yxURwWl5TyLUsjWUBO4/8RbXJnPcFiHUMqDvMqFWUa/
m/X3v0ohEBH8XFwyUI/6rrqyMGtbwr7WsMIUp4+Aum5UDqRDd+vdZLA3NAns5ibQ
Eh3r/JvPuc7XZ6G0njdHxCXgnoOB25NKDT/XbYMkfBVy7Z81EX5CnmYb4wC984Zr
qHZuF5rkEIxfVy56/Xt2FszTpg1ZuB3ufwCUKs/tUtBpTr5WN9j/JSRpGroq9j87
QVEQJOTVAOz72XgR5/sLBqlO6sgUVvuCNz3EmIGWz7ON0AZXsMqazDoQQCoDyR8a
oiwPn6JTqW1bAuqUX2ED+dGBgzMNSVjctSPkfmXH09bJOex39lYPBmvFv0hAQApV
KNz33WHS26m7WMeYq5kcXw8/Npj/ccH9J1MPV5saVXT/kuYCK9WvSDx6hbF4DatS
Gx5C8jrFbeVksq/kSM49Bx72JbS/1BZWSW56SZjvyPJrVSerN6Ol/cQEnc/afrlh
fQOBwHVrvo/KCwKaXF7A+w54tX/ias/GQ6uCdJASR2EMS7pFpH2kNOEZd/UFoXIk
6lbo4mXryHevUymHCAwc+VVgrwCJuksu15gCdz0eKpKyHi5YcNmlwoqA8dkwrTFN
13+p3hKxI0dx8UpOPU6AGx1p5o4YLR5X44DJmP8gw7kUB0EjTPgGpfC4SWZqhfg8
ZM/tR3gf/qvQvMibw9tgkeDS1rr6oy04XAdkNWKBd9OLfZYtMTSzEJ600Xg0T4bF
8/FydYMEH8s5P5T2AimOww==
`protect END_PROTECTED
