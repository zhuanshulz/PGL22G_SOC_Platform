`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rcymoA+kPkK0nczgSge4WShwbq/PbSHPJHFfWPoMRDlrGEXEcKs9W45L2jOKjI2b
C0TV+u7PpVxRp90uSULd/FOeBdeEhSAgmDUQ8Oxh9HbX+Lzo8KPZo/WAso9f6H9p
Lk4/DHoCkzIvg0e2KUCt4KU77DcXwdtVyiTfWKOSB/cIKgfwAcI37u7nfZxiffni
t3/ol92JL4TpJrl8IrnSyguDgKYPqww6PkQ+75BJC3ZElTHW3babWEHz/3MKqJGd
wphRs95/lYJQ/gmNYqPiCwijStsBsUbdUG34p6+XJPqwnoqsoedrgX2uRZygc2/F
ET9On7lA/adtt4PqCSSlHUmXPCjHbZkc0iABd0ViXryzijf+ZuymGL6R4iN2Ezbp
6VEPvqGhzJ1SwaBcRlHl30+7jfNBIRZCuIbGlc/GCqioznstgP81PTWg+EW+QwdN
QECeBI2KyFnvywEx0eJnaaI1R5cdPOH18TX+LHZzEmpro+5GeIiVUFV2oCJLd4yq
QjmPDimc6yhlmYtDh7g7oo44/FKLO+2RgkTauX7UESEEsinqwkCXpLa5qZnzrmqS
OpGjROJxPSPCaypNFddyyZmNOZoxd1IA8JlRlVSDeP64WVDklzjdhkYIecaF1h8w
i+eKAhODDP1LRRBE16SIqyH+roRy7prNNlOGtkN0pYE92FxxiljKm0oJ0C9emvID
tJCfyHQAHcxHc4znXV61j2Z8KkJLo6uEMkagOkJCteuhltCfNIxDyZw5S5MVly6S
+BOzuVOHkAT5j7XViVWzm2uARSf0Zpc/uRtFSHpQRA/fC752CcsNoNVD/5ywEf87
YF0qbaVLOM4DprUcv/DElYBRGRB7CqJuYPLueLMFXox6h96TZxtXxzkPJX5m4QFV
EKQnNBL2bBAEZSELHB5RNzPDkVCh88oze9c9kropV3soEaMXGrpXoaWFFfNVltF9
Tvj8Tf91n21RloVH8n3q5oE2UovaZZlo3MZBU6xbmyDFhQdca4X1fhcbDXbQiqiY
Wbsue+sCP/z7OfpwFQwF6w==
`protect END_PROTECTED
