`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i1+bt9C/Gky6HM6S4ZqU4CwzKtGLxZ8PDOXvXkVlSpSWUdquFU0MpLcFSe0v0IGd
tSiNc+eHHVYUw0VbW8gM2rv3j3O+EXLztx1WZk85YTmxQcalAZigVYHcgWoYHaI3
b+cctTGG3iCH5tjj4AkAe6ZsWhNfUkkfAGcuDJf3962/iWzXB9CG+tJqlZth6dn3
JHkZAe+13AxHeKBu6Aj/OG5J/LqoW2JObIWMRAus4wXEBI7o87lqmvWn/TsOWHwC
mxfRB4cL6/IvZ+g2MQe33zIpDU/QHnQJXaSN+pUqUgJZtwQ+zzKbHt/5NM1DlYxt
/QvDjUzbROop/Xq+aJLc9rJmTJJ0svo0iIit5e1GJll49DrhWW6PVL4JaqyYUNtN
QGfCPgMpZPDH8Ton2045d5uGBBAv6lvVF4H+NjgtGJJlAUniO3/y/DiKvfYbXEHo
UKEmyl+qvLS/oRuIGbvrLRHtEjCY0+5WuZ1r/NrDJdE9fue8JsQa9RhLvfZEIq/A
RSagg8/P20q51muNyosObPuSlMr+/iOUgl0rd+EzbnmVwCCV62LfQD2nR/lurH1k
K7mgZEy5I9W3RC9d5aDC3FUWiNcr3+F9j5tNwKGzuX8tXj+U2GcYvIw0hF09KmN6
L4E+K5Dg6gYbPzOJxzKtsA==
`protect END_PROTECTED
