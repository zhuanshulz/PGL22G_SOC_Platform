`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
51BK5PH6q2JqpPL6r6bICHMUgYCuMGTgiX0qOgj5vzng+VeyC/IViK8uZ7nWcRSV
ZUDvS7bzaxQ8gd+rsKgvBeGNzhi2n2mo3fLwrzn4enCBTGvsgQiZRyIVg75/xNwc
R/Zof0SDtoYUiKpp6Kon9B8mP8ssh5bVbnxLTE/yiUvFAniyn8OkLLFFBhNP1Pht
oJPIfpts4hmaC06Fs6ES6F3J0KBXBanAn05hmLErMJqSCPWSM9rWINX/CrL0vWlC
LDNhdftsnzlrnSkIc2JxGTwXuerw6uf1aQGlDlbrXsk3pmJkOL6aBlIN6hcQ5bly
jr52exviQGf7xCeGi0M5cGte/pWQpny2QdwMkp0aKH20yoczpLUyd3lHPo4ERP0s
gW/CT7CjfMTNdsLGktltbePSnHZCp/BsisEPKDuGJLqgIeZIXqSDrLIr/c62QPwa
oKiWsLaABd6qNgNroLgNIqQad/pf3unHtNa0VY5IwudRAlSyn06MbZQN0w/9ua5e
PmZI1L52LAD1y2MLbP0z2jJiDaZw6+JOAYrjY1w4hT0e/hA645EiCM52b/7EuA0F
z5mNnPG4oLMdLy7hjVVjK2PcWrZV/jhMnXNkEPio8QoSzJXhv2PzKud9CIOfaZbI
IUhEFnVrFxo6OWfplc2WxDHQPiscxhNYvYVUGGfvji8jPrv1IjNVXbXLYcm66yxO
7ILA4yqcsQHNpX7CWWvdvBbRA+vf9BzWYFLT0hf0lkkh50iAqomVSm9IUpNm56H2
dVIONlxAXzZefvk96k2PkgCy5MxhHi8zQKap1prjxdD7LC76gHTW0TsZFMqDIomt
Qak1IXbaH4BXhOoDdMoS73ST1SEA5jKN5isi4Y1v9uNC4pmSPJyoWA1EZyJqPQnH
A/V8qM77BGslWEY9NsOPzIEWcdiPJCz0DCh2Eb69SfgL/tx1AwreXOnteWyiV5br
hSXfE+TUfj4CNhjyEmJTerWqCYFemxrtEfd1RLc6k1wv152hf5FrC4EsD1uKma7A
qwduv6wsOhgnX8rEAXvPLbs3ETyge+kfTj1ACgEOcUKpFq3BWuAfeJ0/v8tJ8zIF
gJrKnEhC77toyteRh2L///qE3+tEV6/FBLIxjTfLRTX8Pddvx8QWlQcSe+P1z/tx
JkYLXldFjArSJX27G8FPxToEmq8IRj896shPlMYsOSaHUcLBRIsiz+6LrZFVwy9A
PdNa3a7GU3O/jECgRWa8T3iWmGY28zOultgmpoh+C3XzRzYCFnCpFk0q4D0U1qxs
M2Ui/7yZh4h6P+3WU9mrCDbe7dYH+Xaijh37Q4T8WJrdyveGQ9/5VYdBOQeJkk6k
KVEIxuH8ah3m06nfWeGCrvyBc3DDrInZe3tz7M+7AnMwRbODQuKI34DCeE/HUgmI
GeLGyA/RDz5ug1PhCAGkrU4v9goloC6CHitPe54oUeOxUfISM526bE1N7saLln1U
2Nm4PLTn/B+WQDREWoEPc+NdSziona0oItYvRgvfBfreV/NSspFZX7c71hQ77abc
ruI3HvMfYvgjVHifFmOHQh6PHF1uRQZT7ad3GTegFrTQJWr5/942FYv+Eei0nwNX
McA7XLJdqb/I84MgP8eQUyEmV9C3OaTlgPislCFjZJj/m+RQtIwEzc2tTqjAGXwU
+wl/EuC8R+OITHtu01wkEZCGHajxKAyU+sk+mMGFyiHpjRuyPcvx7EsjactC7OfI
Xv8qvg0Z+EVHXW8soQJtEu8l/FfvEgyzepNf9bxIMw4+y73BGWnV1paF6M5YgXOA
mnThwIfewUXCzSS4ZFUB9fOgSo7UQ2pIoukjOvVoGGYHK2Zld63PYvEqxTssJE3H
m4y7Scbn9FvirPh62hAH2yy3lpq2OfRbSykh0uJuEGT8aoD1IFaqV1tY9V0SeKye
GJxt7fil4gj5It8yNUKtuJTMbWi1Cj3OWxM4fbvzuCJKoR/3Svt9jaT9GEwXYWDd
avEVRgNzhwUaOR+G3BilahTrpDiepTVr0kOCGDqG4ul4r4T/2c9YcMKHR+spDuSx
vuJkTaDuACmbfvqLyLgKeYv8/o15xCaj8VXcwvrlZ5/S9rBVLTH3/fJN2CEujplP
pboxgmnlUntoqWcY6FsVDU/AmTGPJQq3Ygc55hnF6qzC//BXOgz6Drs2Rfqy9f0u
uX3kym3vu44sqMuXj23Jcbfh1cOusM5Z5yB4peenTERWeGp9PSMg4gnxmGci+Gww
kF8EH/nAmYdKwTEVFH2CM+lMkqRA6Lk+TZayriM6e/q1YkvmuSO+ddwa7pBVcQRT
NmYsv9usIQbeWAyshOud3ZXFuUmb3Fcr22C9ig6Cz+KBKUqJTxkLdHNMZIc3iiWI
iUm5RkN4pZxT0DV31pQNceeomd3gv8h4malDk8MjTsRjhqaRxJKzls+QBGM8RAsO
mWi41xCTWhFy/5rWiLdllb3H5xEN0OYsOkzKR+x8QMVyo8Oh1PC7uNMkDP88RdNg
hL7oFiWsFJFjbuEIpwQ3LaC9Yzg1+bq8greCIoAIhBMvXvXo7XRxkdGjt4yhR+av
Es3y4Q7oF7XSi5nh+pG+/jg0tSs6TaLpN7G+X75KJ/Y3H2Xrl5IfFU4VIFGEI7O1
bEmkqgd649AemQ/DV4Y6LxcaYM9I7j5dZtPRAlKkqL5YQb5SnpxlJ0ELjz/H5EGJ
ffmc95lpfh1tZQE45MNenZ8IOoZX0+fw4dIWLvyEyrKnbIfuRIDgNQMoIm6Hoek2
U/Y1emodBbH9QpcWXJ7LzwlKCYKbpMc+3OdSeJAL90Q45uiZnhZ6DN4KKdtbfaFQ
QrvRwcwAGSGll7AsthAeV9SNQjoaQry0cfxAMvFknv7FnCjVY5gGRvkOFv0+M1Bk
1+OqIeX1HXzALnwWqcEpqBaEdcdIXT6Scrlrbyf+zjI1pDW2tyNvRGjAyFl2ghfF
lbuKxFo2ZGxR0VkM8BXbyCPSPO6F1LZSjTHMwj/pKl/TP2MiVxvJuQiNo3YKqIdG
1WVtVuCCi3U1WVwG0ppBHTQw9BvFHOP+S4L6ciN+guP32qPpqZzDh4GP5sfyPCiv
eJ+qqWuio7PEv29GSvIfZX4V7ZifWcEo8AjHr3+MpsvpGs9Ikt3EOOsq/Hs6/Rqs
eTuy73rIZok5aou1p5a8QycH9rkJoDG9ZjMJlEW9Obrez+jLKaqMgYzlnXxU5mTl
npjID4Wpr8N4SXFXNNMEiIHXVlaCqmBDcOFHHgI01hxvdBrA9ooWJqOsslAaHoVY
ev+rU10rN78ueyzj/6wjS7Cadjad9iaTuqsTNlWr0sIMRJ2PkwAJKA5A4x7DIFo0
oZ3fcHwiQBdV+PgHkfpG49o7JniCLBH1bPqwdLHLIj9kj7GeijaiPatAFZ5ZgHca
bVrnGVtpRGEH/i0Z2WbvnOpO/ui/0IV+hObxIBMjof3SPFezdDeHaBoJA5dxzAez
99Sis4xvIXxJN9fkTzmqxle+0NngwKwYe1K/eN9hwCAWHbVZoiW+xr/a0J2+Dhgb
GSfBgsgBKPGRNb262ELdJxRT6NJeyOu/eRUi4M4GrZMDzjLFAXEmnQysQW3MqszP
SPjdFuUoSNrpdO/jgbuLTJz26J9Bvl2Rb6ZqEvOqTBGl359uKgoHA64Da6pUvynb
`protect END_PROTECTED
