`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jD5jAd4GDKxyPRzyNOIOJkDxS2Y3tmTDcGG9TifGXoH0tkFaaAEM1IBdD2Zv01ke
PR2nie41keXAtgX5+k4rbpJCX++zJekhVz7VTbgNkWHiAMUH1typJF02pdGTGwkj
9xxB8FgFLCaDrqOI6ptbtR2vYJY/oISK6NuQ1BaR7RHXL0hDbw5UGDsID4whwYsZ
VpS0IsrS7REOU+iQZ3Del4ahzxrP10BDK/A+iUQ/lwbMHAnl2UGbb3hQLTnAgIVU
hnQBxcDHCPk6IrlIZvqfvgsSQm/TNJkCJTrC963ozDNihXv1t+wlPUY8ajJXlRTo
wNt39G63NSFRB7ezZwcS65mKhw58I6sjzMJWrfoJbDbq39OyR0zDHVwccvs4dwxy
RZ9vRToobifRtBWoGfNFHcTf9afehAx+N9LYpduni0Ll7ugBRphPE78AGtwp7c6y
3g323psivkv5gJSoP2z3ep555kPPhlUelxpW6xvQ/dGFk1xGgVXCg0HYIEQcbuI5
W92C3UH/z13VsZlUhZt5wCBRCw7E5ifl1uThv8QN+ey7oTUslG9rxMHLMNVJX+VN
7Jn+uUOqMemT9uZVxCGnmLV88Ueq8++J/iGyduq1dU1YNQFMpRN/wdubiC6xlj2B
o4QWVoTAFbAH4RjCTdiXmSoxGCH5TPZrtiSqI1yBGYldCB1R+JkTg+ufFgFx9NaN
BO/BuF9iV6qjjHAURREt/VXHm8val8mcF2gzvb94h5InO0YIubiVpcE7QDUG0NBO
p4Hxrq5awSKwuNF1FitfylxEKM/ncX/g0zvbGtpKHLIYx0R/Ri6XevAEQPtskKT3
CaJBQb7+FgRCe49krzFLQRSzUftMVvYo9UYxmwY5oyIO0cKdDvhZjl/iiePqXQ1R
LEUDTvECJ1y7u1AbK+QgjslId8qN8XIdCZ49TMYFoT5iJlC4eisewdRZmztQZ9Dy
LiFwMB7a7HEEiEO95JG+uZ8xY8smWUAxFo1kHzXZ74mm08gX4FgRnYE8oBDTiDr0
pys6KdQdCtVZxTqErcg65NtyMJROfSgda+onmzOft4AFN+ZwoqMVMTl0rTBKXAd/
VMSUTN4kfOpdRl+vKLKdMuXNrCJFXNksylp8aKCsmQj8MTTa7xWFThEPJYOsN/Lj
STsyw6NH+WaOqptWWYWn6reUzSy7MaO4x8ijJtZjp6y23fQ5b9c5dQMPzr+gCjUQ
MKP9bed9MSxMh+b0KUVbI/3dQqiwHGEqqn7SeBnVFLTlmr504Eq/Rk5j5b06aPOM
CtobTp1xo9EDg4mxo6Wz7XkOtU6GaMm0ZjeepbBxZponoCqx8ak5+phHE0PlXfRT
7Ay2KaEamtKR3pEhxf+jOQwfmG62cUygWBcUIvfK+RxkQDyncaxzUukDaXUSC2lU
wIHQCIcD8/0MaG2mQw0oSI65ZGMvAUKPaaO4JIFUxoLybr94NQYFuIX9udBcTc/z
x8egCcEgpvE0IEaryYvgwKc3l2fzxQXHYpJ4puGPsE6x99ALkVFwfs0Uc8cX3lp+
/fiBM3I73ObXl5TtPK4BZd44PC9rOkNlchUdXhvejishtLpTQHXHEmMgdbwpgKCi
xhVCP1g/Hy0YPs3oxScW7sRLBydgco72BvuXC7zWnSBofQe5OK4GQTcNdJJus2YO
OePTgJZfnobRGbZGcqZRdnJRUDPSu+f+gm92gAoXmeIHENpK/Bdovx/HjsKGA4a7
DYzg6gXiwQH7OVE50zZsPH9+Yw8wRkAi8AgR/dUyzR8LuR4L8gjYjlj7Oly4KKim
RmxefyYLSlnb6oMtyz2zMlm1CNNlNgX5ZSdXS3aJM7g=
`protect END_PROTECTED
