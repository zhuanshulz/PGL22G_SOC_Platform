`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I2iE2WSDeLqCFuRJStG9CAx7b4UB48cy8/X6IJnXuj50Xl2kJAA12kH4V24NMEpD
FpK3i6c9G0HO2qXsurdmvwcvhCeXatcQ8c8S+jp++WV11TB4hCXJ/lmBfAEGy3Xp
xpzrmqA0OJMw233SfwrG+KJxJrKeSsyDiY9FUdcGUj4YUOO7w76L7ZDrshkNf9x7
/Ud1tLuosKFSKyXhZLY4djX2/iV+BvnbM4Sy3ETnwGYiFCtMJs2QjW9CyA7mxSJJ
45yoLkSAnNJFFwxQirIQwEUGFQ0ot4NGPeWBP1IU1H9P4Beyzmpl5bpLu1ypNZ65
d8MLfxmqyt227/unSDRxUVigNvwNBJ6CT9Gq+8MgeX+d/aMeKQBw0Jynk/6nnJK2
13F1rvgwB1lpANuLvzGDQeg14YdIakMFtH4RAu32eY/8pidjUN7d2b6hSlZke18D
fCXTdqh9Q+MsHhP4sxnUhYNJmCmFfTDKX+WOp85XsBUrZDRp0WteGXld1hOjGeag
NcnuhLNwqnSyzb4ntciagbr3OcJENrFFNaKMeT/FzN/RBKIpI0i2l85FfWJhtNq/
b7IiZ10Q91Yu2Fi5xIrDxW+VsCvUge9pN0M8X8ntmjFhhRn6aNaa+KqC+Cqa3CJz
5WFZYPmX13zqV2ZC9mew3XAqTjJRea9eXJpNDlyBpwVjCLrn/5k7heY1BG9DtDX+
+3WJ3M2+dQa3s3RALp8VMH8X1/nrg1lwCDlxHR5OWe9njDTHRZeYCTq+pumqXCsq
O91AUH1AztBsrckPUyA99owpZqljzEws/7Hk3dVF4+g8Iq3575VXtl4yn3ODkY6w
2+0XULjAnukIw4ivaiSIRePwI7T1kcjbItFAlGnxFBFd3vWqn9FtT2/DlxDgKrsZ
IHyNT6s5e++UdZh3IGVwT4yTmk/ApYjf/hibDvpKBZYj4GKaaFyiOBq2keVlH3Ln
/VHrCheINjAMpD8Fm+AxH/EbZZGaKiCtvV9tJciyws6kmoLd2Kno5pKzdMjwadmP
`protect END_PROTECTED
