`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p407hE5iiejrOFpQHNd7kUJm3tyc2MXCaoyqciwAusZUmDIV7SMOPYagkfgTdS39
s26uYysDzsyIOPRYkN897Ep7uW2QutXVwBM5pxqCvd0HfZPklFX+2zQysftCd9go
pB6sl9mcZbuZFa5Ie1Ul0SM0csAfi003n0fBBCEqvP841ikkTcFgSTXrCIY1/8Bn
Sv7Fa3Xb9JZERj05R0XT4+rBa7bn4xKPWVffxRlbh5F4dwdO3Jmdksgm1igRCn/y
U+luvCdkNRyDshim+C/bC/991ywxxJAtSgfcT+kVf57HMEDyamvs2O0dYGq5/C3O
NpbUKrvsr/2p5nuBu0ibHrSl4YBlBzV7yt1/7PG1kwGj5rqIyNOMOtJI4n6hTMXl
Q0aYq0SDpSObY3GSADFZ18HyuC1leWYQ4HRa4kXiOoamoClQmB+cJZiOUkNkoEBV
`protect END_PROTECTED
