`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pYvAxWkDVwPkSYXRakHyy49d42ikkLm8wdhfwhB4xLm1YuCUaf7MYhDEDJBr+osf
gbYGW7r3T/OmpexyNMkgUuxMkh2VG+U+c3QDvB0Xz/UNDXRbAzAqLE17E86V8/+t
O8dy+7X1b7umtb8uY+SowFDlvcXnw0IOrp/+axHSWOLhFon+Dr7g+ZEJnILmmt3V
2OCgOG3laMgFXFVGvtH619Lu0BuwxYtQc+ZWUWRIygSM6nGIF98lnYvLnhYWR5t/
w4iDf/smQdGswRaCeuUeADh4E5quiLiWmqfDsTk/QfdVhZn0A+8Vtgow1yJXpxpw
VHmHSUeMuFQDK+x/VZWSgsz0ZJwQ/rzjB2Uk5PJ8/ZJLscLOX4bpVMAfSNAB+9D4
+XLCKrvdMSH/NxBPLw2RDeSqg4tbMEHN3tIGge3Nzow=
`protect END_PROTECTED
