`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j6+rzTzv7dpwp9peycKhJgnD9xxZaETH6fMHmRP5UItg0EDM66MwDJm5S2LijNww
Ht3UYHI8U8kC3nHOh54wN2Nf2WymHax6Xz3GiEYiKEHsSYCksCa5HIsHG3Uc/07z
vrh0x4Osg7rAfiWCayGtgKjpbry11V14Jn4hCxKr5X7KTMqPIz8dDrcpSPp6HLT7
SKTVpghyRgf4ifl4hlj5dzZBaRXHnNmELFucMz+J7sQBHgj3xn+1W0mc8+y2Epoc
cYYUbyPAmV1rAHa2Tik8QBefn8HPUuPS1jt87gC3WJMe5BuCC3jyCD6TfjwPcFig
Hdxcx/4UfB/Us1eI/TDGddml89rnXX0KgI4+BYLIU8tsCYiNzX+qmSwH51shd11w
`protect END_PROTECTED
