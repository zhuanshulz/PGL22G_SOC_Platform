`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uJy6yssCKfFzRBBV36L2DmBZmbzGGUT+Bn3Zw89go5orkB8C83jh7fgiqTVYsf+c
NihMu2AIxAtBY1pOi5f5ghnKvL+D0ezaXecXIogEfKqklY/9EpQ7wC8Cc6Hbhfhh
/fjQrcfYfAiPYch6AAFHbGyxr9HFRAnxxtO5pHmsCP5gFPZJ74x82O2rb6FyjOtd
31CxAPD0Hd7iyOtqAdrAEl9DUddouHhCsL2T3mLH+vQpMRnZ1O877r/jo6r4vTK2
KabtjQFgjrmimDRERgNlJyGE2NCZLQC4eHs//EnUXj5HMMcGbH8JhKfZVvRYgA7x
SjriaiYASZc37tnaDXPCXojuyIZ7OB+iCWsBccQa3RfqyYW5whDDKa+peiKXIfRn
55kINc6IAPgbVGc94VRckYHstCaCDmMI2Vx4Faop4jPHHtsvvUAAPvSEq4YCUTAT
HIGWy3hzJzWa5hrzdg+iTv8QxlagsobjP1vwGLFGLVI=
`protect END_PROTECTED
