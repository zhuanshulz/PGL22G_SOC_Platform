`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nNK+cPb6KyjpKu7x3IGRcqWZ03U52v4OQ4Mqx1GyAg5nuKwpZUDIi080qmUBSAzn
8+X+74k7M+JCV+y3x6oogrdtqFBwr0VLYj+tvGLejYojEm6kQ8keKKH8M7N0TaSe
dt8Eobhr71Kc5VD1U8RztvnqABBmOn1waKUcZa7vLENYmD9qUu58GIdivbGfR/RN
3525DohG/JgfmyxmIiZzmExKMU1QU6AAAwn+A97tpS15M1IQIrcTYR6FQKYKrHEB
BqExxBPV0KukRV6jMNmpooQiWj6jsz+fzg5KdT92v73j2uHNC4Ggj353kdYcu1Ww
b9a4sncsTejsQ6rs1TIwBd091hP73iDFq3zEk07YG/v9Ez+BByBGvvDAP3lu6RTC
ZVosR8aAMKWNFc/wDmzTp1++tTJNIwcI91aqIdo1omDySO+7ao3ucrXsxGqz+LnC
dDcA3upRM1lSSzbKKGVCPXMp0iHOqieIy6K8KFPo5rur3Coj1ZL0yAc+AKocKETY
t/KY8Jq4sGTdsACFbO6CoHmicxSKXNa6DwRevtrn6eZbT9qLCG1PsC/K35NUt7Tv
f6b7TPDImtz50aNZQCnFGm6M1jUAILKrn5G3D+9ghTmVdX7Avs4aKKmqgqZuWnQV
`protect END_PROTECTED
