`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ybWGrav9QVY8/CrCkwiaMwGl9po0icRUe0h0HhT2mdmE9U8dWuKhMxKNEgcrpfW7
ZFpW6Cgdp/tH5Y6fDcgbJzho7LgwDynjAG4S15SWkBdk3MKdHw9SxKQKDX+C4lay
XdjFOp9zSljwjJiHPcl4Sv98gQTQHogWru7oN4GPs58i8GazO799hgTPyjwtCeXu
9IB/QY40ojGAcxQftHAmG69GM6UAb6bfBC9oqHcQjYieuhSFc5yDbPHZEculKbjJ
dMSHHvKXlcfukDXivMuBbGU97sJ3p+AbURrP8LqDmzaHbjWCLWS/IgmHQ3pHVsaL
gIXJZ54etSyypNjpaCEFcHzkpqWsxzVb26Q59COIoqxApNODIwFD06LwOcjXe+K+
yc1fPY54E024OTyCUD/ZOdj9PKqHLrtIksWSeR8B8TVgSbvemT9fNKnWLi5vu9/+
yluLKClW8RgZ++kjn9Ct5U2XntMHRcru5g85NhjXdPb/q4jnB4nypxHTFohTXi5G
a6HUI/7a8t+df12oX3r6VwkAs0OtXv2fuGjGCYQhW42rky4tQs04rq+QDK1UhBc6
NtP8200X4d4WugkUCmlHv4bOcFOyxaVrIp/XppgHYu24xuDnEVsin8GW/vICJZTU
Sy8THwgb5YFyVeeb+l9Ha3oCH4ExK4AoO4neWmi7GB9MWkU2REwEJspLTk+05Txt
BaaYK6yhQeCUoqRPb1RYje81/m8z9Ysp86p1wbQeFyZhDoUvr6YDCevxQyVUKq0U
ZKFIQZdWsLvDUsWoZ7o8myreYediZpyXzeoL7b0zxDlqIoAVMhpX/+xuBKcmL9PV
lXhREprBgWEbgpR+ofxdhf86eg3Vp9WQQHMj+n3jUFKB/yh0S1oeUfXt2fWc/Gnx
/3wB4W8w/rrPqdV0Tm8BFJGv+SoJD78yOTzyyGTZUFsvEwHyYxDJKzFiDRDqHIjD
HJ6Bm4m1Po4MPbBODHIBjyOQozf3TZiXKfRBBr9S0WIhLeg8p1g+HNUJZRXnfIxz
hxy13fFmuhaG0W8lN7Xz4zbCvVx3gKrn2BJGGeAARqXryf6zbgOqPIeC3nyZ0P3V
VmnUorfmozgyQBrZJLxaEZRgAkJqPIybBhUGUA7jjW/gnBSWbPYrw2izbb/pMH0E
DykQ/KUUXbQMU0o/O3BovLOTiYvOoOaP3z70mvZXLxhjd6Wf3PGroIa6NQ8pX9Kb
CThMbFsB5Nw1M9NG0s3e2fcRNUoQqkQtXn/7tEpKBpyA8IdSNF8oeuvs+7Z+/UiY
sdRsLoed4vEeb3iDBLIbVTQNz4MctNun4gz3YI3Ceav7mHUNX1n50vAV/1arrcq4
wAn8SkFLL33+/9v5lvuMqgpSxZHu6cYhBYOqC7kSRfFWmjuUYrBnxgNsBHKRkvXj
gd0oDM4q+8FDdznNe+skI7h4OXYfF8eeSRjzmLsaGc0J4Ofv/AA0T8bxmHUqD5Z1
nzZTK4AHicUYh03DjcWhHHQzaW/ZUzhTKQV3NBgkXa+JcTCWFZVNXi31wV3aveJk
cHBViWFrFwb8/IK/DCTzhVuEKYFqRMQ4o4mzoaW/dwz5AuRkKjMSnt1SMMsNCmUa
McRzoAjgGRLMkXypF+KztbFJS4fKgtzG2mvJ5z93I8E5kfB+C/e11pL2liXQyqH5
IYZXbLVwU/5jIqP5eoHlWjLm47ZA/aLshhW1bikfeQKZnnxrHor9Ww+9Jhs26gvZ
I7ctb+gtrgZoLgruvhB1/GiaCCriFwWMZ3w+mVx9aQcpE+Usyvzr9r+oDSe/o+Uc
j+hS9EeyzmwX3D7DL2VECMoSR8w/KLJHvaKDJn26Lod0nlhVjzObTE5JxDmdTWzo
b7AzboQQNHnEQFHYbgN81KZPkKZXqPLRAmqQnchsOKanAO5F+blNLMV3YaeY/jb7
As5NbrymzR2uWYPYMKFCBBxykS26CagOn77U3HzgjVDFdHPvZTHdWGVqth4UqdF1
CcXRIgFUMVQMDnuDEkGXMMmfLw+b9h6mYrX/mRYFAJ1K8H4lVJEZLTyaLNXY5inM
lNvqGkE7QuCCHDDDPkBjJaHPPl7pNOPS560xPaLGefCu4oPTlWDCAxT6ljxEri5Y
144SuRSTv2QuLvUBxSXa1iidJ1/Z729cKv1apdSGHoFSVDZbYZ9Py0PsWJeE3YZx
5T+hZIUpMkObOLO81xXDoAHMAmMo942TBh1sqiSqK+cmkyCOcOZBjHVAw1dLT60u
8Az8DKfzJp8qkj3HniIcdLLpVNt0MeY94HFi158yxEB6OCHh7IyK/gq+3P9Eghq3
cS6YvfFnJKV8iAZn+Sq4jMQZpYRVGhARaF66hvg6DOfsNiI2aTMMTbD3K0sTen/p
Ocix29oDyysr6qJNNTh2Pjb82K7gGgLA8F8CAj1LqJhmOnO5BYoPQUC29h0y5zTu
iG9X4Bigv0oQQw3qhxON6woQiKokDcKE55gimG8l9S22VHKmxuBd9a0uDGkVNgC+
Ix6x8S0L4v4rHInU31dT7o+oepmip4nFX3bf52SxckwNgF7riLwHlmlBy3NSldpP
PY0oIdWXX50Nf1i+gI2thfD5cpDiYTghMbQmC2Rq3YzT4NmWIE4C7W9P34Tm2ZF0
6u+glLhgGlVzAY5A7bjiXDT7NpEaDLtXxn3cCaht5Jm/HWODJ9o/ujWKSwBkWhgP
QS0Y/tbbzptdcbsIIEOsoV4UD+t00MgaL2Q4B1bc9Y/47lM/8lEk0/ygKy0KCwsJ
ThkOTbtR1HCR8tJoZ1DtTiya2NgmK9XRAlcNYrFBAVEwPCEXr7K/+ULj+O5vT5Dh
Q7L6cUUchgfy8163Ig0ZOloTdyV+LbzU+MK429uuTDufxfdFR6PET8SeVC+N0SOn
mT8PJ6SWyHWZPd+v6ZO3bxh/EoxRuSxEavZ4ub0qa6YkesohPj/uvkpMjeN65dhK
qDS5xK57bgliug3FlpJ3PzJm0OGIb091Ci6cREOiRFp9i0T/yy3PRiGdz6ScuJ1E
3Cd/UaBW4E1BML4iq8G8+M77KUIuV5B/5u69TGPehLVgkMUjoXaPWw+9jCwuvZEb
1lPVnvdpJNBYR/Pw2JibX5KCRFvpESaBu7avp8pqyg0GGfXrRccDtsLoQtYxU/gF
IL8p0MAm+XjFK6ozV4APQCGyr/gxjDGASQ+mouKDAR7jZ5rv1d4n1aNRYlpdcOAk
/sw4YdQa0YGWQqJ7qCYZNR+K5JAC6D27M+3Rlv9i/LDKaqi2uSqamRKgH0bDII4u
S5oZqFYXdSUFqCibZrPtP34hq+SnTJD76pKXF0ozseMG9Dwz++rKHL9+rrPospR4
6y3nOWv/pQCba6w4EJq7LPIoRq21gMu8mLwzt+emr9/WoTmiB7JQIDL37fzVvODt
YHneTsMyZohs+dpThdgni4N9NlZQg+mo9nGC1BrqLp0k7hIMVr+lvUvJFHujdZt7
piacl7KTs3dsIrANOBL0I3SBNjTygjM2ufMACEUIOsmR9Dd3n7poOaqaNRozG4dv
yAeBVYiqnGuxwLhK0MGyTpPiLrRRGoTrmgG0rWwr98VvVCOf4mEPTe6K49CYfPi3
Kjl64QqaNGwLeu49eoNJBX+2M6XGBMiYQSOIRFBN3OfgHv9BSrb9iyG9cc+ETuM+
Qza3/75PucW52fcPijOPdznaxIWZHnAb/XmIU8cVwp0X3bN832KLxrwMKk2euNDg
PKzgz2N4T5ENm2SaA5Lu5my2AW49gYEeQxGH0WaDlL98pyW8IsnxuqbbFeHuILH8
YH7/43fG3BsuEM/3erSqAvPSEftPGRxBIMt/gF6fnXd1fZo7+Ga65hmuiCWWxGlN
v3oX6VskrmzPTNvYToqWQN1BOSszQwfNjv0HGQsWw1mFQMHUboWZdGdpHfiCOwYY
CxuTwIh2AACU9/EVeekJlcryZqJrifrO91sjyG4ePxjkQQ29o//GFQMciF7Jin4N
lphDT1Aa/iHZ60pIHC/D1+ME8o+X9dvKEfgIXvmi/44wZ08N2cyuHQuhBxrrUyYR
U5eoVWWOG/3it8J2a/zLaPVO2UhvATgRZClxXlnqzhKgke+Y8aozjPUuD0L1+BzI
WTTFPuk5wL2+ezTOzPEp1ZFYcQVnqoAw/SfL/DE4/0ve9hX26o7BKVO9odynDXHV
2UuLE9XqipLndunaRpmxq2sIGe2g0bw8OxVPWaDraZQAqRZwxWmfL56Lt8+YZueM
2+QV3B/nv5o01RQh1hx8ZvKWzlszLL3ha/+wqHVwRjfV5t66jDWiRtGnbrWOO+qv
3YzX0kKxgtnbJEUlnuE269ZljMEC7hwQY0xDtpgu2GO9JFz4FVDr/zBqawUfXXsv
mn73htbkzbShqWGXgFlcfGLxVbPnc+onrOhjIpr2fE+9C3raeEHboZmC3XJb3fje
lgfQ7BY9SLjWkZZ0DySl4ITZGUi1S8x0u9voo1v6QI0XGa2xVtlNmtJUGrsNErvM
vDHBM2oW6z2aQomyzfZC3GLhoBEB3JTK/py8VT7iA/ifPf4WAEx2vh9idI5iF1eU
Hv8R3Q9JzCgfflkUg4fLTWDuXKi+1APjbkC4U265I3uZgo4opG6ltMmJ4VlTY2BB
ZeTbmxC0IsUZLasramSspRCu8Zfr9SNFSJFBrb2y665XnKUThCuayOAUrJKHlWm1
hRp9R1haN8OswWF2l560SfdLR6AmxsKtQ2bg9FMa5gbN9EuyU9kOKTzhGwbmO/29
ieOVu6S8lselPXg2HYOc+PxE74NBRrfCzoh+/3ZBRuGyJhDqcrbirHspnb60lh/p
X3fAqbzcwzlardE0XIqm/j2DPAoy0bwHH/ar+yXayY4VDD99BEEFykLNQXAGd8ms
HubpY736tPwGAEE2Jz0VsTVvY4BPmS0aEdeHXPpJDIHtKAa2MhrKpCLXSU6ExRIm
M7Okbn58OO5SsSMW/n2jZOb3+wz/fJoEdnh9m66nOITEiFOx5Bu74v/JsNPomat4
spw9Ahs6AvV0U73JcQGWIwIhPWfcumBWsqB1G5+ltGez5EtNpVsZO/NsaVLwxlfv
ei0ayBey6kYZlV2rcO2KbuCvHz2nxGpBLEyX10MQytfPq6jIXtbOMyzVRx3gtNG0
WeDr6Nsjbjr/uEdJKJa0lSO0jS87rqO9mBHukcYj7NHQwQINc7GUtXCsQQXSwVNR
IyUci7cVVTbY4PninEGzwpItaamhFDvglxItMjoKib4xfk7czzx6LbMfFBsQii+K
03F/vu6Ecu7XCVVUsiYjjKNudQVUPbubU+33pbAhSxyoGN1tLiRp5ib2P4lhYH7y
Knfu2jTTN6hjwHTPWuNM18k68YLE+o/VPUJpx88wmyIiYvSuNKb+Jk1a5PX+iAyJ
zV02iAONnAGYpHdVIDxP8bkdThdi3xhsBb8L6aIMPRXGMzx4aBQYGglFruEERsQW
JFomBSk7WDvS8ifGowptox3wsFJMnv0vjAUAmp1uuuF4XPPkddgPqbIWoxlzLhp3
rO7DKKdYp9iUmi7ZF//6aM9pwEIuJs4gWYr9u4Sp9TEywdeHAl8ooAFRCzL9DchP
cJFj6VWZsa/PRwn7v7bVjd29KOWOOcZeduEvw3Bj2N/x0r5eL+R096EVEUGkvhsw
YYqE+eoN7/fsE/tQJyTxyu9Tv0hgkAKaRcYa/KB9ZD2PQgNzoZPRUrClRbe/xCVD
56FVC3YOTdpc7iwOBs4+fI6zOz+nRoVMFFviPodTza36WJRZdRxTjohmsQU8pZgY
MRTMOlHV06wsahs6srEWnTrZe48SaZPjigri4JVYd6E5bEYSyqNlG68xUjf07lIn
qLqXK6sOKYmZ1Z/ZUCKMd62iCgqUrwOidDqvruItXX9CoB2lBGdGpF/3dky4OLEw
BNhoPGmPGa4UkHOvv/50QAuPrsGOZl9PQScfb9JeDiALQbA/Rvg5CEa1j3Zk1LB6
xg+SZhbLsUERbzp64mAuKN3xPJaedlj5w1eFxzXnrWGK49lZoGwT6yKP3nj+pJ2B
dBx0lPX8Bf6f98Nb0fh1UuuTQeHjYL5YJVKXFbmhi5LNIZgq+veTFBVFrtuaxAd/
oFWtLiSixRhIqYyMhUZ7jt2oDhTCP/7OVqlMeR5ybhtQAGNa5pAE2pXZGkIyKNQf
mpFEfK95D5tk0UCU/MbkLF+YL3ZgI24aARud8F73QYT3JggDSlzivXrzQ8vy5X+G
d3QukYMlkgnG5UYhnWvdZiHvo01+lgfdlfbzZzVStKhq2iBywZYwR11qOva26UEV
suDcP3mVl7niaqBoIIymEJpsdGl01zZOmptVhp8FVE9KFI++j4SBUtxyLFJN+YUi
UwYfQE/a8KqjgNpZVL1p0M7gK3WmAX94riYLbZXrhLplh5bXOPYcmdPpWxmC93Oc
JMQxT05LqcTZIqP2y3Ak/0q7XjSD2oONNOHPx3BN07SQ28Xzvv9c6j894/5BWVjH
dbxiXrKdVpCyKh8ARQwHkYJ7bqzbN9ycr4i7S5MdUlO2YOpOzkA9XdbX8pf8RzY+
w8TQT8SWzgE0buVb7DyAllLmVjbythKSBfFsYBbdmAcgdVkfB9m9SblMN5W75FOw
2QYJGymPlJzg3f2cM1V5XixBL/w7uVF6+OfetiOwZ/SYsiH6cCxHf9Bfv/WoAQ0r
VRe0W9tfoPZF8/QsQta6BibmkGRED+y/UV8XoREB4EyiIMfBbg9zgYodCQnqHl1U
wktgvJoLt3dC7dQ0hCZgis9WfhyAgkwD5jNsI3Uru0Ny24SNpB3ox8qmgYGc0G+2
WUGOU//u5jpVHBu280bhyb9sDQyejKJxiZGqZIkT98WToIg7spDAWLZQul3F4zYG
s6RG/0Xhw/24qVPHeFTWUc7b0D7phoNzU0Ar85ZF3DHgS3MZgsOkx6Hqrd++1fvU
Wk+eS2L/lJ2B1SjZdcUN+4l2+BcmjvTxjQbyfCUDN+5dHpuWD0Q5+APL3AT/AK4h
nq2gXER7n8hSRve3+JFFcpeqQK6uqJxlYDRzlMQBhpNCDr8IbA7+7Q+1kt17ChTL
xaTNhjSZ8Uvg5mlkzliMibIiFOMdFm57mx1z9t8MYAYVWDFY/ujkNMwq0dMRgqTU
VVx3sNU58MzUyf5syxFUF/l7/CYoVfnODTYG8P4H2uZrXoCGGa7ETVgtsExrP5bM
EJR1tIxJo0VCaiFhZfUsg6dYnn2H62manhRuRFnm9LTGGywC9hsL8Omk304r0imz
Wi25SsDTqHOF2gdPlwGQVTTgIJYZtZZifZXkmVYSmeddetoAWbfaQ2ayxOr2fPC6
7WoWoUy83mIk6iUCvFKXJA==
`protect END_PROTECTED
