`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N4bixPXLG3YTKSTt6weMWQdgTQq9sPRJdhhq6kxgIqZblvUGJRYruT3cS6zbzIOH
/MtwZw+rIPDjdjB8oVjRHSWFTp9MseqDJvFcDaI2CULfQrpaNMhs1fSclqxYq1iZ
qg9d7irpgXBTfpt9fWHdOYnmZstwxytMyvYxp106Vi+zDf9Fta1jbuugNkwE2Pb3
SATLTL66xSa/FzbfCFlLzdGmbclVY5hrDT1Q826u36rW5h51ZjHhkddiUiL4PZyJ
r28O7tGAe3JaFsf6wFfrUw==
`protect END_PROTECTED
