`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uBPkf1AMPVpC12/fqvArwVk+qA2/EH5CjBFRGxDnN5dl+FIwYhsJGMMdkvI9PlF7
xb4wo1JsfvErMkOgjPtt7PthflHbs7sL/O13GBkI58d6UbZdBlPg35JmiHdOqR/t
/ddBYw7OCEKh39n4aNQPPxOyeJ0ldlHtLgQhAidQZNI98yt2v2GLVSbhR2QrZhLP
Fuqu+RE8u1S9dXbMqXYBftXAd3RL5Ef//WhItM/eAjez2Rar/7Grl4jqWQrkDYRV
FrYsqz56dxBy0oDzJyFwjSdQaEOy7rwAV1MNGOrNWcktSgleaD1+P1zumxiiGVxZ
o3S62USH7r21RVdFcGHx8FtOW4UQfd6Lo4YhRmyx3xpZz4Lspk8kEzXijMsVVofX
naVowKzohzWvsi6p+Ry5oCkU/jCb1f4Hj2usDir+U55LNNIWdP6df59tSXPURLQF
w+koC/FhP7e6hntXdfzwdRhoW4VRYtcswPPPWHSBs4IcZJGRhen+q/uA9GKmJWQA
217GKkFFosFt4I730lNsza58Ge2Ws9mC30iaKjoHD6s0gVBIu0fbUAdlh7u9ISb2
e7sKdXWcxjV9klKsJL8kvns2toTYPwnzKG40JL1tIlKOV8kdUWRyhB2ZSCk6XoCD
EtOqUtyVlvRh2VVuV8CCZDOA1+T/EEY/Dlnkg8w6CpTaDW8+dHIlSk+XPHTFWLzk
gCm52xi3dkQ5phHkQMtUrFy8vrhIol47p70JXfxmPXLIES8AH/+tutE+Hdr6o7RS
5i6ndnSPg1vd4FK82SIYz6ONK3/mYvT+Q4JlYcbGvRM/7YwtzgaogUNc7sqJUtTo
qBWtm0SB/4ZiA8QL9CiJsagUil1Szv932Dlt1JZ/5KFDulAgwATVC+Mb55SyT7Po
efcWwzQfgRBRK5xeWvzVcZCJ1Dy8HfePHCHMGI1QNbOC/tqF7jxyLgUMPLqiR26R
hOl6otIYlqHvuvnFr8ns1kd93H+E/6Q+/xvGijVBfx+txuu88uznJ7bAi1rLwQmL
O5a9/JICwL5xYjUKu1tO1tuANUgygh6gYixFZeSbO5S77QXrAkz17ru7cpQBI37x
VpZCLAcqypDjZnUit+w2iU8bgDkP52Kjk0Zkd2G/fB+qwFxVfLM34XnGOQ3wtlSG
KItd3WjL1n5w2jIg+h+N4I3mOZ0XqA5awLsS06n9Ym9rr9Z7moNde0U8GMb2X+1e
nwnGjE6tA4L2hWp6RCv7tsNWVgrTWJ87e54wcA3PM6My3mH25Zok3aFXLHfKJATT
Bi1uXtwcss2eIMrprs96KilsAH80k5z3nd9EHtiC9eW0TBM7Xnsjw7aDOoW7dbnp
ihisj+vH9GcIXwVWhYujKrH0Hc7Zw4Qx56mB+Emp6qzeQ9YaRNZ0FE6YDAtAao4C
7vsk+mvs3+heywK3fnwAtvfzrmmEW7EEvmGWBQp3qeEVeepQE8Dy7dlSy8ejl1R6
ilIzXRBVIukiVf04zgpRlu0q9wyJlo/0Hdhgdnn2q5bJZwj/AJJXTIk46LmiHAOF
GbhqNY6dxutRIvm5d1YdgIM4qBVMETq2EUmXuJrc3rSYQKHYKcmRqYx/WKZnIYuj
WHyLDXIboItw+PrIBw/pLUJklrfgqKWn9jgDCHY8JsgihH6mmGvtjPq6yKtk0njD
8hnAC8UeWk8ij7Nkyr2065RufM5chdkr7sLCyyRInxcYx1PWXEd6fOWxeuyP0E0O
mwPB/w7MnMRCHvMsu/f8BPd2ZIYGv5dJU3gYASrOBvy1/2Kej3aOzjGUdoGersz5
2d6mUtNSJOckk2JZg3Cp7ABMFMAFR7BbZPiWfoDOIeIeV3MvxvihBSID9T2Pr11Z
jXrKRi999XCqqfSCb/cUFXesizgKJ/VUy9N8zSz3chG2sTDNuTcn6nFfn/CQhl1+
2vOaQNxM2IGwA1ZovtC8rMX9foNmSB0PJUapek5Oz6aJo6/h+fRk/vLodVLTGdhf
1rwuZaZPqP68yxFQTTg+OQAFkMaBr6uCDUG85XWt6kvczwaOiDELrsCRtHyt1ABR
JOHk0WtqlpsVtHKMhg5IHdxFjb0P6bKnVt82SVOB4Kc8iVZIJ2KlQxZOhncFZ1aS
mtGLNX43Y52xVaPi+1lORC+foNi4ddtVq9PtN3QT2mdMgMAyo0PYouq0CBEXfEYa
isNiuKsp0azRd7YaCXUAlOMUmnjBlxXFZeigUDMl0oXmfTTQ1tMDjmBa1O0qy9XV
D8DGPvlSa1gPdkt25T9ESJyIu3KEgrYYwi2UAe/PCMtBhmcRkxh6nUCXdykVsU3C
+TQg50cinw3ICkS6KT8fs3cLEWxCpp3tDKToS5SzOK+xdI/bDD/XzJ/ycFtiHzIb
qOzaa4ypw3lNBquq3rhIgtLUFFLx8Fy3NUPAZ3rNj1xBcUY6e0dVhid7KWxUJzeu
GDSF0p+HMYhT9O/BMtaPaHElkFihoL/X0QjJDHHqIr5aLyuG8dHsh2SScHVUpdsP
TvUx2itfLQ63/mjbqIt4r+2sWadZGo6g5rXEbQYlZewI/BD4X9+/hP0B1wcdCA1s
8wC2I/WlNB/xdMYRlbKoH1w/wPgdrjLST8RtztVRsRYisS/XigCD1LP107S7vuS0
LyLY1z7TTpTecUNq3SQME4mTcsjCmajmZY3ROIf8KGs3HQxWgbFLAlz+qzjjSwvj
P/JqxmER+HFyf5jsAeVQDGEREwNsFV8uLf2BZH0vNQhruPVNe661Dveehxu+TXuq
cpX33Pn01zIZgYitt5w9+MSdKsbfnwjUHY0btVwNnxT5gUKtr2zWq3MGf/+jZFCX
nY5drM+4XvW1l/Y3Y6eIaIkyMZwBbkpFSe3oW6EyITfhNASU/+yAKjT7VqAtl51m
voEUIm3Y7EzR9oZZ9b+Nyw==
`protect END_PROTECTED
