`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+a89WmyDC3GsyAlWl8B3HhMpEOY4pcwz1/RFh2xrP4Zw7YBjVFcSL+2OH4qtwzpL
4eQuNAFqstkV16jschVw/yJC+t8tE8wwsTCml0S5RwY2EBpLZ6cLhID9bf5jhKzI
hkSb4pbzPtgfoaBql/SHrZgKZG61ktDKnOlIF7LTfupo8IS8CjCW2FiifnlQ8++1
E0Xa/U9DkWOV/VVXgahWcz1lOOdYR6hzMEMb7LHTV+yQWqzin+XYX6WMUoN+rlmd
T4Xk8cYnKFDo7RVHRHsnPi5CVNkhlCuRMPWe7gVtqlPDHEwpWbkNIv/V6L+jtqU7
Z4P730Vaxqg/FHS87Gmi1+0J9dIWnos4fIq5q7QSogz40cZQmoMuUFI9eUNsCziA
LnBZK1XZefDuTjoYoUJhZiwdB28Ron+L1b2ZfD+rmvbye3vF2CTO31tc621lF2A2
XWt6+7V0Yxt/nZODbNQG53FehqAoXfUnAulmPvTVBjRoW2Ul7B6NLA2ZzrUOWe1o
o1ei0LnDOda2i6g9Yu9It24DbPEZT0iKFCT+PO+foaBbVSzhJP04F5MoZNvyYovZ
sLmrubMmrz8DhEUyQsnbIvMFRijYE5QUCsOfxMvEuWEVBVuImnOQ14Vd6BsyVUbE
gGqiyGQPsubFqWsYMTbd7w+Ub70qaCEGjbuEDDLE6TO36By2+NdS7TQ9XIz96OrA
+IlkeoU+wK/LHdLSKZYHqR6Su8ankWmHIhqk9WXynw5XkoicqvMd8L0cfRLs6Bjt
Q1CbQdlh+1rQBPAvzOwZxF0G6Z7hWavSrxyo+bVhFnVFzaXcLAWNLUYSZrvVHslS
qtLGaFz7+z6rIaJaB8qFzVRJFZDzsoJoa7mHLZRhcZetwTrApT90Cx2S4P6l+nwv
v9NooJJlz5PtbXtcIewhRKx+EGF19bOClpR2TsY6ieSfqNFCJ2WwJ24+vvxznCK1
EBVeVLMrJRJcPJzYHX71POxj3GqnBqlmM2P81LZI3x0xaXFzKtVkJThGN5Z7+Laj
c49mH//fqeUE4rSm2Lkz5ArxwWzAeK4cx/4C0LfuVjBg9nNmy8s4tC3EtJQj2Dpn
pqrksOLwdRUmTWK3Ln0liVr7YQ6IM1sOWjQ1sc3LNpO4fXRek44h8N1gaEuVcVZF
amYp6RZBhI6HK/1uD0Xtrc/kFO1j2AdkHfYWy5T+S8GScP1ZclJA7lCxA8MVS0iL
VTNCx36nQgrWuMKjCLcIBbvRHs0S3vVlGl6PtxuiNuFJiY85KxenOU5NvteFUCnb
ukpTdn3HI9XEa9j6RhuoIa+FVclQnD7/hQqTK2TXDlYXDFSFAX/WZr2tFnc6V4rC
O1eUFVxqY7Me3Fcs64dYn3WFdV3OmO32yDixda1mi3zitZ2r60W6BHcWnXoZQYvp
sCzNXNvedti6pXaOOeHURuzI5HXFxss/2QABvhg5ppU4K63sBN4m+zaa0FvnFDTK
MxzWbY3bHBICrQh3i8pkf21bVHKEJkK9K9WpupxbBN9978WtVspSJZB68Yi6bA6A
/o5sVo3yrL/ziXq5Ve/wYAHCNRplup46ZFOEimmt7OM5x5vCrfwmL3INmeGkPpt7
ni+aOI571lMK3EfyjGmjB/Q3S30A2vEnE11FgMukX3UpTxq3T5EBbFfrcxqKdxkq
I5HYcP9o+y3VhOLqktr0FDt57gVNR3WBR4lhnuda1+9voJ6epFIKOlPFVWwAG1eH
iCIPeTJPHKBs4jUcIG5HGymRWQi2YzECJGyYt7txBwRfOJwh1bApZlgck+FZm8AP
ei3DOuU8hCvF+gFCjY1Hn1ETboVfH9uHoTQvz1e/SH61v5HpVOydDEw79uc59qqF
gVfiher2buSwXoGvWhlUJaYwMA0tFfRMEFd/XM83V3YK+pjPGWLtJ22NbLYOnpFg
+d38NMgFp/Gny0H7PQfHRTOhzeMATjrthomByTvwAL4+cCL+nFAlFBoZAJuUZLMK
xBq7sZR5QVsfe6FfTIbRlbOSe4UzazzNohT3PZHaHkRIzwtxv1wCCm1Swak4+tRn
SHCPZ5giXHdhQ7LVZ4eKg5QmflaSt/2rjKb2zD69O9IPHSswdO0NCdpJclI6tnVY
A1cr1/+QZh4hTef/eZf03qm60Qjd2WLwsKpbE5fxXteesXgb9TBMvs4w2vmg3Xvz
n5BmOVIaF//vcz8EEGWg2BQdW7pK3gMsNE104bG434zMgwnWXI/1gBry/x5G7cbK
oJaroEf1aHO2c/BE2M0uB2zbQfc6oLMyIMUfvquHb8Sq1DJuDBjzPjvtG7mBJpPy
k1tijS8Aq/xTryrwz6+2CLnTEHj4rfRrw1EiqiJ4SC9NN+3eS8HHFwcHEnDg7Jv+
aRD5Ko1GKwGhsiYhbWKfNABR3ViHH5nshDAfvl0uiJF3E8aw1pwtzjEW693Tssuu
w/83yzmEDBHRKdL23qjJyK+bADNsLUriT4W1V9QmQStQZpcdxQ5SeJB9MJaeuXlO
AF0HsH1liBmKbSjNEbfFkTnrr+1GBbfhaZW1dmk1uWYjQO0sr56Z9wXe2BwCB1Oq
BSZDeMkdeiRjKXElbMpq29PiRt9iFq8DZkWaQt6eJPirdrn5mBUqWdadOFDYGpYv
WBzyKaquMLXDlkNvaGK2HiuduSSY0R50qwx4k6AgBmgJK6lPcsAuhH9KhJSytBQY
DuKdDdt4hYV5fSL3JNxUQsUSNLjnd3i/SU2/hj2RU/50AwfDoryOrsIXsFXfKz4r
dKptUWj+4HVbnprXW8k39EVMrO9zX9wUEEpv8Zd0bET79eikcxSRhGjVoqXbS/xj
kD2SL9Zxn77KfADKkyC/lfNFJx0yLJS2A1YcdbRluWZc9mKKIMV7mkOAa9T+GtjV
n/NNAzFiWonGFsAm7GUsUPCNd2MMjaLu+7PjYs4ZWmDI4qpSd29ifWLnzLOmJJDB
HSmnBe/InEORSV1vctHq/Q==
`protect END_PROTECTED
