`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4HEcB0Cu72C/rKyb+5HgpEe00SWi42Sq+ew8/FABxUsFVa+9W8JbirsxKzlnq0Yp
9SatMMAgENud/YVvv8jOa8gubs6ygcM2znj0x6D+s7/GV94fWmEkKlUymCMfN4zG
lrif6LHJ0pAhMQ5Hc8ljTX4IXDtnXZq4kDFucMFhlkh5SyHjEc9V2AdwPIhgA1Gv
9lg+Pm5inrM2CzYW2/Llr0CyKmSK5A6dRpQv9faDLWZzYRyXDBxawLWZCREwxo2j
BKmLztomvrms3dttE7sZ+REUq2ae4DabVNqEU0yFeQwq3PVuRofHke8DbppDX0eO
mZ4o6XtU9bkpkN6CKoHARmRBrL1xYfpqOpSBxh0zM2FIZQI9N0lswBZ4C7gNmFpH
utfCXfauee9rrtnFFWO3RQYkXZgB5j2PEqjfX/HzfF8qzHlewTu0m4XsQECxJ7cO
4VUpBiwS8mjPKeCWqQ4gPh6h0sUJLOvtKxYHDt+I1nF+f+TcDAIf1u/WzdCtDlOp
mIDy+/M3F3OQft/8XN7Y2UToxPLyEcNbTFN2Aa/p47LecQupHo0LFQl40q8w5UoM
DPxA86xB7ewt+oECQJIwbEN3oojdAinBHlpJmo7mXNUgynnzJe1oSRskJJfbeBJZ
z0FMI4I/sGE6+uNOSMMI7XNmLARcvdmd90lnL6RlfZUng5Xj2BOFEVk1xL2SkOAy
7+9ZtzkPkRveLrnOJ1dVbRlw5LtwRLTGNfXlJvY4ybQK8neNHCaFCMP8T54ZKkqm
FGfNqWmXizHMnGV3b4W+Ls0pJVVGvcEYuTuGxjOlwPgxwqR8CEf4SiOFHmnBZeJi
K3ol0xQsaNjSvDLgLq45azbL/cUfnF/0LmlfeT34DGpBEPQQI5nYGOC5KrCzpvR8
nahLN3HNK7k9rsWu0zJRk8JcZxSRLvsAR7ijgVBpwYTlUoDvDtpefxltml5QMxDu
uvTnvK+meVBmV/cpqdIueRDvV348QHR14diCiAQrXsu2UDmJwfSayky5twyqb8D2
dTmO/qrTZrv/RZZLUvQlAtVQJhvQsPtNVubzoSD0Lxws7XYcyXr08dVFtHBqmqnG
1lbrm1uxOY0xtdqeuHjF5TDFR/yVM5QEnnujUlC45l9oGq+Efz3ugyeLsUG5EWZy
ecsMyt41c+dOIdYX24CxKcDf1576kJ1xnmYw9mjv1J6gFsnFTOXmG6D/PzmL/gJo
kfElyUKrqH6dP9RQk7YCGNpRWH3bmTuOAZ2Pz4ofN3cQ3x7YK22aaKLPP+t0xpCd
nPC+cQSVMluFyEFKxkCLQM+TbOvEouwGuz3MMMARzlaoy75EQcAJRP9F/0SID0EP
EWKD8BWUlkSnkxRt2PDE5pePzstNZfxFOXkN1AMO+7agV6GNnhQ7/mI5etZfz7iY
LRGORjeA9miAWjxSakjf+92fIrq5eLJKGVt62F1ziTNQzWjY4zwoyY4JgkeN1N0R
0c81j43DXyg3tT2jcYkAu+FrMC/WVEIcCBxNBj/fvFRQk5aq2qo4cVYhdhxv/PWd
kt32SKumXoyPAcIVOuOKy8aOsDSMXad+Qf879yLBNkGDtFS6/ybd94xBJjsvfNtQ
4TVJsjTCXucWHIpoUspY7rQJUAib55HKbNIFKZmXPAi3sDyha3P+FsLFlvKgOfrd
S2qey2YcE7XVL1mBINuWAnWTcmI5p1QngWu0kqP8zgcvQ6yGiiM5UWGPl9xuEYXg
qGV2ifNnGn52QLGG6dml3FD3goclWPfQ2W1O9DOhGl5O9B25g8YaOWhcEL1IA9Qq
6G5ag6D/Qs0y6cLwiM2V6ZyJqzpxXUCVNyyaxVzoT9LX5CBqaHOPJQ5wgHmthq+M
RRoj4+rQBdK4u25lTnpHXMPB7BUqOGOA7lfxq3vljcGXDPS9k27SIGRqXZTc/4i2
OMboa8V5fXowJGtWi7OYfjXEWbHTyPKJfU5ql54Y/taK/GteVNSmNeRfXXcN4TLj
SEGx3TR1Q4SK8roXmaBYh4fZ868WdLfGXK46bdMws4cqVwAzcjzTrZiYalCpiNEH
PONF1lV388EnelA50tMns4TGMRYhaUVkGI72Y8/gqXNjS/8kXa4/SOyap02VsiPI
s9rYfk72sGuGe9wBiJ14PeIiWmi9I9Sro5sycOAFUD/ZX8/BkKTO8vhyd7yYdgK5
e+xqRDKdas8YuSzEYJbqLRjw4tr6IyuLJviO9bpy1xB5EWa6XTZFGEjnjHhKKlOO
Dye3GVjNOuYc/djy8Oed86nWGWjAfkl6lCZ5n5SKLrl7ccZqmdMmyAkTdSo52VLt
Kk7pzFL7ihfi0X0bISjm9ehmOmz4/HCnPBx8G1ncbpc5jvKo1IM7dqWWqGJpdkPT
yN1F4lKBK+5mRKGKaWKoWUm5uEjtnNVCNT30y2xBeLNIasAqYnADYwW4vPLcxX1W
94iR1/cDdG/A8OCOpcVX03Ix4WL0Y9pVSgNgXvJWmasxU2j3trwMNR+fBa4gII63
/L2vJ40S4VE9U4MmJbQ03oc8kzyKGa2OAXkEnCEYy8OkXl+/JbP8tppYmqgRMcma
z/zfrY55W7hAeXw46tjNd8avYG3hhIKZlAdlUEMsyROarfsT9qnSadWJyYNMHPkF
l0Z8jkfacGgoydXBoVWvvG/qXjK6nuDubqisJvQkxKYvWD7cmex5gjQolNtXBW9C
qW4bYJXMSq+BxcM8g1DGm/YDS47LaOF00sKzbRBhKdd7gfDrojIXvZNFgdfvyoBz
GE3WdElDyVeh1fJ5hGmeAw==
`protect END_PROTECTED
