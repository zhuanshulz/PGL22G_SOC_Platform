`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VmEisjI4QaH8IdCectUZaZm8zMmoX1AV77D88WdUvUdU0g0VoIjkp0QhyfCrjq4x
ousI/ua2wZ+0kB3zmdaoJfko2C+8eJDuGoYat/vVphBFdlI6LBrcCt/q6ZXh+0Cx
1P2Vg+y4ZjYmaYyVmMfSL+uGaczjzLhsvFh8FdlbFIsTQHfEHV1VdbGCvHpHYNQm
JikBbMsFp/qLqQlSnnjOd71gI8IgLm3T5o/Es/UCj17mR9tUTvcuJVy5bNabnRHI
gkZFlVJgRiQZcP8QPhrxqsO70wSMb+fw4tkqIc8ZIlFs1whgkwNvjymZqaqjnlcc
btv/pWXRVZ3E78Mx5W1NOIbscP/0qUxFAEPD2KH5w91I5DuiP0l8QXQ9F8SM2ER6
z/xiDYncYJJj3AdC2qfN2pVe+IVWB8QAdX6jnzdvF2LiXTLzN8djQCEkuuZ9u9CJ
XfjK/7uRI5AGUvJ2EbsjTumwmLpkJcBkZFpiut+iUT1XSCtWdkqCnghclwYWc6Ac
8H0w3eWad//CLCcMCfZMCn3uOFlfcVY8JpugIYxU95cDUKlSkvA+5t9YBgskyXZj
4tkQcSM4M3J6UNcXpMO50w==
`protect END_PROTECTED
