`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KRaWpInTknJEYAXEsgVgSQEMlEbafvBe94eIaGEk7ncfqz0Vc7JEYyrJU9Q5ysig
WbHPscPcTMgAsBwwRkrQjBeo2owpzXcxDqRBgMlEFenJ3k9+lRiulIH3cRN7rLZ/
EE89DZGVJR9KTuyeiThsSBPB5HCsL6l9S4YEhECqVJMIkyLyb9yvQQ9y/LgejiTt
nNtGBt+dFwii8Jj1Nj+rhqLgi6znL5ns5MpFEjL6yR/t2o00bHqhvPUP/eDbjUEW
iKdG2hXcgWuIVSefSuaSaA6Ksk550Xf5bUkjRdXCHk7ttOQGXbm9OwaYF0B8fUZb
Fd1lZn2XzGvyXaMazy6vnX1jhxBV+XR0wvJpEs9SxFiw4mPCqZ+f2AxOkK6Zbo/+
zVeRRtlcya+SfyUBRHJZlp589Ns0ltromQsz2H0Zl+YGNHalLBxcLkKSCIzov7zB
UFZzFT0tCSB9REs8Hm61NesDcvLkjyNndOh/as1Cps6urXk7pFbf9eEXsY7CNTVT
zvC5FLQNtHfFVLyjpsFj4txQdf9Via4x4x5mVql+XnV3vlfmTuS+OLyBmKgX2sDb
hDfmte8nF1b1aJwqb57GDfEkmkD36wR/Y7gl8e65o7X92L5yzASljqgR/Rf94jPG
pJ/tEZlZKi7cAu6VEtpuNbs/rl2yBLXynIUqqP8QRKwd+c+LeFMmCuaqmYRlXqHD
sa7RlKXXQMkL9uB1847tmaFcPpRZm6ageX0x8i2XaZ1JiFHyTOj07sgJQHOd34bp
cugfvQa9MQB82cAJ4/doUnA25sm8Y7ZjfvrRvQFIWRnMH2LVLnKzvybgaP09CaSd
f1nt8w60EzuLX8KlceIx42/waAEFQlauRIWXEt6/BVWGoIrTLIJ6ncI5fvXE6sAZ
B8TA36RM2FR15KencKTxLQ==
`protect END_PROTECTED
