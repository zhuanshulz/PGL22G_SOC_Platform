`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KgF7leJp+KhLpJRxjl1JIEQfNcyPlHH/SdqhPlrddf8OCvJEYvdT+8t8qOFKpe77
rysnofgcittBhv8ELubNCgeboHyUPJBORMMUs4lWzztz8oqbyJiqt1MgI+KoYqIy
x18AD/B5n4roiQzvgruWUndKeU/bLQyLwE/nOA7grxYyXPZyPitEGFFD6TTt363b
pVqhPashhdun99f0P2RhWqZEZGXC0KpZF4oY71P4kgN1n6MQ1Aw1hjMam4EZNfll
LHHLdQ00DTBrtHXFSJ+6icjBhZv+78lfXXnJrEfc6FFWF+/s56iiwgG6kUix07tt
GhrYQalNcY9oQIWg2iu4XLxc2aPNUk2xgW9sf883wvMWssNNGkANGKlGOBTRYWuz
64nqOpxprK5RNafHJELTnAbv9JJ7X0gGDYxA8Xa54eeMtpWvV08n5L+rLmRof68T
LEVPwUz3AWy6Q8vYzAG+cr9YdKgOlj/921s/Y55aWdQ/vL0Vn3jlm5iqVsGFhnhx
5NInOB0Lrl1TU3QpnopDxhM/rvZU5hU5qCci8tuPz9zO1ghKozIX+gZnpYys30Dy
qzGn9afh1Aw+IY3Bzh0Ub8HJ8DXi1kxqVqAcMOxr4Bxclc1AaGRizwPPlucYQmKJ
oUuNqAQJyYka2EH1EFUK3excf6tLGEVjsd2j9eHJWgFxXhVXna4u2BPd/Sqjf89M
8otjqA/Kn/5yjYdVEUsH84OOfsVGIzm9HVOZgXH7LPeN7LHP9+oS21eqM5k3Jf3D
A7XvX9oby0k32ChTEQcjEaxi8j426cfvwCKFzAcuQNY1Wv8/mD9f+UA+Qgy3DBdQ
lGZNb4d8sgD3MCogOX5jQ4C1i9hpg/l33pUmFNhwC/qRMxitdLfDjfeKTBvlMMGf
Zgl/93j8H20vSHhO5QobFX0rP2dJ7/pMqnzy+bzMOwOnRU2x1Y+wl2EWd89MOJKB
rMx/1MdNaeBmcheZTuZXx2tjIUwSa7BVwGEn/G69GwrEBJ8s61Zx7nPQamg4WqiS
eL8qAttbz8E5eT+p45sV8yUDneTolRODmFkbYIqx9oRz3IqzIjUqJJ4eCwOFxTV1
fsmRm41SCAG0al4oMJr/0Z6xXu3q73ZYe9WLh6BqmG2p+nJfD6fYe39INiww6z79
Gk2ny1RNOXGjZUSIOcQS+RRfR8RuJdXAO0TCegxwnIC+d9VciE7vYuihoBrF4CbF
y4B1PVszL0EApGkS9Qt+c9RHgcaLHSpR8eZZUA2Vk805x5AeEVtaQLb/tCoRjb5Y
VnF3VQm2nAp1Sg0dcSHS1brIiDrEL6ufvH5mwqcz00nAa4YMFxLhYgKx2+F0pIZt
F3ahACqVpRiO6yVMoTDrXVgAIBTp3dWfeWz5tYH7Sn7Wk6zhelMCf87VtZhNJsHd
dRfZF+DZ1IqbXzWyiwfhUGcb2EQjrUwfgqExYCJk0yxJRv6fVvRcXqaaBNTprz71
mVCU6MsAf+1betWH7+LsPjOrgV4Ww3z/wniRqlrsPmtqmhzjaItajZvyIwCK3ChO
VkDGIOyI830l28w/lJXnFd+jyT0fUMSzgxgQ7DcBsw8gWTHpDdJCfl4ppudSQTml
TdW89YrZ6lqYglGFNlqj5QCKq5pIn9vJKgUg9+UxiIwpNQ2KCpnnVA0J2FZp5GPN
Gby4/qiR9HNkph040bbFIgYC8aY+A7Y7eEzgHcK7yNkQ8qXsnosAd8CIQoj3uDsv
lEL8A4nOqLOwUEa6SDK72+p4Flr3IOA5vYo8Y79z6ghCccQTiEbznrgSJbBp+GAf
uosxzQEs9K/A8OZoRXS7VKbTkl9bEBWk3Xn0WyhO+aaAQa6uGdQSLwxo2+qua4xe
oqxShE3ZeTIVQpVTakqAgdKa16QWgV0J68tJUTJSUaNNqLYfAcNe1kqjh7zhVhoH
FUUkUbMtE8R4nvhm5ELl2eMyGsZ4MNm5g6wg/sv41ad+YUHT4eRg5ev3lF6rXUNa
FQaYMJ1so8mNxyuHv7YY1IUbGGE2tEaeaO4djASva89ecu6D+9DS4T0cINBde5Ee
3tOABW1jCceMID6hPs82wzsaep5BBU9faT1Jeqg4hekd+wnXAMOzWeCYU6dfP9NT
vMAot/OQAjlQ4yxtupLsH2SI2m2eFmusLWId+H2BLwONH+CWerMmVJE/m6r1YBQ3
JjZwj9wDy8RBJlJwe+2uS/djjMaJlwg+vBlmr5IRyWDv2KFWF0As2xyIK/JwDNC6
ayfv+CCOBksnvINPcRY5paRD03CV3FMayBYq7kgYFu6976WU1uJh/eufOqqUyG6c
MqJ+gNpwDdFjN2MMaTtwnJnQnj0NH9BRm+pN2W2TfvEdp7ZiTehmfl39671xCTk+
W+AugcuGzEvwtbDySSaVfyDTWzisuZ0RIJ4d6js7wZZLD9OTp1j++GjOTM+Z9uWx
RL/dhV8Y71xo0tpR1g1AFO0r81dlF4aFBHypoqvxGTNsUXTbUcsq/gnKzlKNvG0H
EJwjT7+TBR10s2BqJa0n8ZQElV0d19Sn8yCicMrCscJ98CoKMlY3AV4TwnRC3AjI
UoPJzSaOI+DlbIIFVhTc83tR+Q79grsrvR1mKuyf3LIA7OdLMFNWrM0yOdm3SvQw
6cuCY96LqHT53WxJLeiAh++e2yGEeOohkYnXYv2yevPdi+BwmDBiv4bpQVPcNofq
5yDfC1vbcsxETaCr2BNApYlavfEGQBdUBPh4/xumLOiHj1z71lgrFU6hepbp8LT9
dXNGZ+zVpp7cJF+rjatsa+KRM6JJvqs/bUsUcJme1MvkRiUvTx8XwQ4GxdSB+/Wu
d223oRnjjWleR0bNtqXK8Y+WWKx+rEGmVcpJ+WrDFYYmeoAOUrb4Hjakf2jOmxMR
ejjLvmhSqUoLOy+o24YiqHcsLjXg2JbhRyUXPRcZxc4VlEt4/X0JxxrtFayhQrvm
oYf0+QcX3QySeuw7F1tkxE27wNZpTKXXC+79hvpEML64LZXz2PUWydkFZsUdFRdG
M8WljihMX03JVP7WvW/h3+n45x2tZE68n82fh9p1dJMeYOB1L76nDS+wws1/OjSa
TEKDFchd0q9Yb7FqzUzbMDhVWbi4ExpLQrlO3MRZDdmtRB/OQ/YL4mST2D/A4c5v
guy6qRfmt5S//rxkCprj7M0VYdHM+VpbKmJKsDWCq3ejOhoglLJuFrS5jYiFcGt5
LEFEh6uBTe4ZPow/Uj+LOX7AvfR/JnUA6re0fIG/fuWqYKrzZ2233waHuzOnL27Y
UESmb1htYzS9LTtGyEdW0iXqmaNyE7PZj1Ey5zTerVdlqtORJnEw9jPoBu+o2S1E
GelXT7PmHkKBDJdCSNQdNsrPYY5sjH6i4jIInSfB6gO3xLPGNt7Mjl0bIKYWPOgd
3KMIgsiMDZmUh5UjUaGYe4tUHnCzFX6yJESUwqZiNaRMdQVfI2q+ZqvOIoTN1LXA
XuWO69J/mQD7RbXnHsRh561qmHQQ52cyKydsC9wnZZ9q197tJggbW4CcQwiCGbv5
`protect END_PROTECTED
