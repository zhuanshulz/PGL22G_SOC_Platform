`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wZnqItakilFYRCgg73vT1g/mmH0ffzZ5bdTxI1rYl0/g/AT3RWOjtSLcs14LLauA
ZY2nWXWADpP29Vwlg2tC70RIfb0FigwDGx1rCIYjAUQH6wqnKrrKlJDkfFGmysrb
QsdUXJJMM+D5sXFL2TieM0nWmp8hu8LqY7euQjQzNSbswp/NyEF/6YThjgGlJmmA
ju9ZLHGq1/kObz+VmHjwlxNnGPTlmwJRy5Fhi27+PTAzxIkHQ4oH5z4MaZ9WQm3y
mMyEp8FtnUODD8w8dHKxV+9/xJ9t7arPXn9s08Spy1Z0dgFTGCSApsfioQrjG5nf
uJVRk0zCtmsc+KrWxoyFOFhahIgfwRZOgNg9/KEkduQgpqnAJdawPQyh1oet+cLa
806Fjq2Dw3SsXlzDgjo24Dp7Ooif46savu8lfHds4ePOjO4Zx7EhnTmlQNdvaAzt
1JDoMqBasy5KJ5cw+xD7jYqtPir+Xr4CRDPW2qJEGvodMix/CEOHZzbSsutEvnUF
/XGlH5aIsBbZBk+eZ8nfSw==
`protect END_PROTECTED
