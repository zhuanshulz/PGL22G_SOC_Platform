`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zg5/4HZu4rqM2VaLnoFx63IcYzINB6T9cjeMAZgM+bNY9DOVZOqkUs3OA5tmRSAO
ArG7MHPwooFMe3Hj9Neyat4LLjWc77dg0AdkG6ksbc+NlVq2onJk+08Zf5phhWew
5EIZcp51uSLxfIpTIwaQ/+yInlcPydGRcbfVJJPbqtltyp3dRrrUpdIifS5+RG2T
caZokcFZP/gSjcrZrPyskq8i5OoQop9l3duYgYFN6EamQZ9/cyLKpc4eWWvtkQe7
xAad3NJYM4QfS1liX5o+TCwSKl3tDqHHGEj6QRXy+x27ym28qPF0tmknKQ7W7upK
QZ8pq0S7ya9PPk/lTTDMsGi42i7LiAAQ8seinu+EX1MCDnKEFGlvVb9v/AVb0VyG
QcxTQL/DWdGANq9qEBwtPKSjmZRxvlZcsY4i8UdpD8nlLeKCmTzBzel12or/e3KM
fyJlF7a69hTm465MWY1CUZG5DA8LS1CDhWzmpjEBv3jmtj2xOKOwUs+PenKNlYK6
aBfIzVEzqG5KE3c+MLcfyoCxo+9Tpg6i6JNP9njzkpZ/O5DmAgJ2F2IOmHMN0dRN
Q3rwyRkKlzE9CIkYBBTKvI4AVpHzI8/Jw66tcJy/3pd42+XVQuoUvzlkwLV+AdAS
BzsqEkKfC9q6G+GGtjp83G60kHkuWfqs27aTANO5KYw=
`protect END_PROTECTED
