library verilog;
use verilog.vl_types.all;
entity GTP_PLL is
    generic(
        CLKIN_FREQ      : string  := "50MHZ";
        DYNAMIC_CLKIN_EN: string  := "FALSE";
        CLKIN_SSEL      : vl_logic := Hi0;
        DYNAMIC_RATIOI_EN: string  := "FALSE";
        STATIC_RATIOI   : integer := 1;
        DYNAMIC_RATIOF_EN: string  := "FALSE";
        STATIC_RATIOF   : integer := 1;
        DYNAMIC_RATIO_EN: string  := "FALSE";
        STATIC_RATIO    : integer := 2;
        CLKOUT2_SEL     : integer := 2;
        DYNAMIC_RATIO2_EN: string  := "FALSE";
        STATIC_RATIO2   : integer := 2;
        CLKOUT3_SEL     : integer := 2;
        DYNAMIC_RATIO3_EN: string  := "FALSE";
        STATIC_RATIO3   : integer := 2;
        CLKOUT4_SEL     : integer := 2;
        DYNAMIC_RATIO4_EN: string  := "FALSE";
        STATIC_RATIO4   : integer := 2;
        INTERNAL_FB     : string  := "CLKOUT0";
        EXTERNAL_FB     : string  := "DISABLE";
        BANDWIDTH       : string  := "OPTIMIZED";
        DYNAMIC_DUPS1_EN: string  := "FALSE";
        STATIC_DUTY1    : integer := 8;
        STATIC_PHASE1   : integer := 0;
        DYNAMIC_DUPS2_EN: string  := "FALSE";
        STATIC_DUTY2    : integer := 8;
        STATIC_PHASE2   : integer := 0;
        DYNAMIC_DUPS3_EN: string  := "FALSE";
        STATIC_DUTY3    : integer := 8;
        STATIC_PHASE3   : integer := 0;
        DYNAMIC_DUPS4_EN: string  := "FALSE";
        STATIC_DUTY4    : integer := 8;
        STATIC_PHASE4   : integer := 0;
        CLKOUT0_SYN_EN  : string  := "TRUE";
        CLKOUT1_SYN_EN  : string  := "FALSE";
        CLKOUT2_SYN_EN  : string  := "FALSE";
        CLKOUT3_SYN_EN  : string  := "FALSE";
        CLKOUT4_SYN_EN  : string  := "FALSE";
        RST_INNER_EN    : string  := "TRUE";
        RSTIDIV_EN      : string  := "TRUE";
        RSTODIV_EN      : string  := "TRUE";
        CLKOUT3_DIV125_M: integer := 1;
        CLKOUT3_DIV125_N: integer := 1;
        CLKOUT4_DIV32BIT_K: integer := 1000
    );
    port(
        CLKOUT0         : out    vl_logic;
        CLKOUT1         : out    vl_logic;
        CLKOUT2         : out    vl_logic;
        CLKOUT3         : out    vl_logic;
        CLKOUT4         : out    vl_logic;
        LOCK            : out    vl_logic;
        CLKIN1          : in     vl_logic;
        CLKIN2          : in     vl_logic;
        CLKIN_DSEL      : in     vl_logic;
        CLKFB           : in     vl_logic;
        CLKOUT0_SYN     : in     vl_logic;
        CLKOUT1_SYN     : in     vl_logic;
        CLKOUT2_SYN     : in     vl_logic;
        CLKOUT3_SYN     : in     vl_logic;
        CLKOUT4_SYN     : in     vl_logic;
        RATIOI          : in     vl_logic_vector(5 downto 0);
        RATIOF          : in     vl_logic_vector(5 downto 0);
        RATIO           : in     vl_logic_vector(5 downto 0);
        RATIO2          : in     vl_logic_vector(5 downto 0);
        RATIO3          : in     vl_logic_vector(5 downto 0);
        RATIO4          : in     vl_logic_vector(5 downto 0);
        DUTY1           : in     vl_logic_vector(3 downto 0);
        DUTY2           : in     vl_logic_vector(3 downto 0);
        DUTY3           : in     vl_logic_vector(3 downto 0);
        DUTY4           : in     vl_logic_vector(3 downto 0);
        PHASE1          : in     vl_logic_vector(3 downto 0);
        PHASE2          : in     vl_logic_vector(3 downto 0);
        PHASE3          : in     vl_logic_vector(3 downto 0);
        PHASE4          : in     vl_logic_vector(3 downto 0);
        PLL_PWD         : in     vl_logic;
        RST             : in     vl_logic;
        RSTIDIV         : in     vl_logic;
        RSTODIV         : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of CLKIN_FREQ : constant is 1;
    attribute mti_svvh_generic_type of DYNAMIC_CLKIN_EN : constant is 1;
    attribute mti_svvh_generic_type of CLKIN_SSEL : constant is 1;
    attribute mti_svvh_generic_type of DYNAMIC_RATIOI_EN : constant is 1;
    attribute mti_svvh_generic_type of STATIC_RATIOI : constant is 2;
    attribute mti_svvh_generic_type of DYNAMIC_RATIOF_EN : constant is 1;
    attribute mti_svvh_generic_type of STATIC_RATIOF : constant is 2;
    attribute mti_svvh_generic_type of DYNAMIC_RATIO_EN : constant is 1;
    attribute mti_svvh_generic_type of STATIC_RATIO : constant is 2;
    attribute mti_svvh_generic_type of CLKOUT2_SEL : constant is 2;
    attribute mti_svvh_generic_type of DYNAMIC_RATIO2_EN : constant is 1;
    attribute mti_svvh_generic_type of STATIC_RATIO2 : constant is 2;
    attribute mti_svvh_generic_type of CLKOUT3_SEL : constant is 2;
    attribute mti_svvh_generic_type of DYNAMIC_RATIO3_EN : constant is 1;
    attribute mti_svvh_generic_type of STATIC_RATIO3 : constant is 2;
    attribute mti_svvh_generic_type of CLKOUT4_SEL : constant is 2;
    attribute mti_svvh_generic_type of DYNAMIC_RATIO4_EN : constant is 1;
    attribute mti_svvh_generic_type of STATIC_RATIO4 : constant is 2;
    attribute mti_svvh_generic_type of INTERNAL_FB : constant is 1;
    attribute mti_svvh_generic_type of EXTERNAL_FB : constant is 1;
    attribute mti_svvh_generic_type of BANDWIDTH : constant is 1;
    attribute mti_svvh_generic_type of DYNAMIC_DUPS1_EN : constant is 1;
    attribute mti_svvh_generic_type of STATIC_DUTY1 : constant is 2;
    attribute mti_svvh_generic_type of STATIC_PHASE1 : constant is 2;
    attribute mti_svvh_generic_type of DYNAMIC_DUPS2_EN : constant is 1;
    attribute mti_svvh_generic_type of STATIC_DUTY2 : constant is 2;
    attribute mti_svvh_generic_type of STATIC_PHASE2 : constant is 2;
    attribute mti_svvh_generic_type of DYNAMIC_DUPS3_EN : constant is 1;
    attribute mti_svvh_generic_type of STATIC_DUTY3 : constant is 2;
    attribute mti_svvh_generic_type of STATIC_PHASE3 : constant is 2;
    attribute mti_svvh_generic_type of DYNAMIC_DUPS4_EN : constant is 1;
    attribute mti_svvh_generic_type of STATIC_DUTY4 : constant is 2;
    attribute mti_svvh_generic_type of STATIC_PHASE4 : constant is 2;
    attribute mti_svvh_generic_type of CLKOUT0_SYN_EN : constant is 1;
    attribute mti_svvh_generic_type of CLKOUT1_SYN_EN : constant is 1;
    attribute mti_svvh_generic_type of CLKOUT2_SYN_EN : constant is 1;
    attribute mti_svvh_generic_type of CLKOUT3_SYN_EN : constant is 1;
    attribute mti_svvh_generic_type of CLKOUT4_SYN_EN : constant is 1;
    attribute mti_svvh_generic_type of RST_INNER_EN : constant is 1;
    attribute mti_svvh_generic_type of RSTIDIV_EN : constant is 1;
    attribute mti_svvh_generic_type of RSTODIV_EN : constant is 1;
    attribute mti_svvh_generic_type of CLKOUT3_DIV125_M : constant is 2;
    attribute mti_svvh_generic_type of CLKOUT3_DIV125_N : constant is 2;
    attribute mti_svvh_generic_type of CLKOUT4_DIV32BIT_K : constant is 1;
end GTP_PLL;
