`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZjjBiW66JEam07cOZFoOb9+IvFkqRsKB1aDvcRT85LTwvpd2nZvameOCbii7W9+P
KMssENUMJ/ODZhb/gj3nq0N/VZP8k4uMhVTt5AqjOOfrhKZsC8WeeUVkjIIFCfQK
QjbDIsaElMCLEWFt3r1edjz+YE+mFd/JNdCzfSK8lpAplU9Gje03srznskONt8Dv
I7XxshB+CAsEjWubmRN2vOMCCBzRzgpf4O4Q6wEE6cj1aATrGNyANja6CqGw+rGE
`protect END_PROTECTED
