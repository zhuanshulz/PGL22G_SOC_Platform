`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xEQmBT3PmPK4xXXvVerfWa8wvl5iqnVbt26Ih+0ysiNrPj5a5iYfQnmF4mb8C7RA
cQihUyQD4q7FGPV3tOEo1ATA1CFY0qIPWaPeDYoI3KIvlj5TkYQuS0ISeCBI1c7q
I0oe4J4pW12/sQZ1ZQX+AaBJoRBjl3tTrMh4uy7ufy5O8Yq7OwOPSO1qHTm4FUTj
E1Txny3x6pW1FMS6MOjvb8AvlC5NRfvtKuYB9NJkC8EbuEs0KbuOMSK8B741govA
f1oW/ffVDocQBtnKnexUJGO76IYRGFn/ahVm03OBUnpPu1jUrSfGOFUoRiOMjL6m
XhMjirUbbW/67HgE8y5zT0HwAon57MyT8sEDpqt3uhUF6bU1oCIVGmzYX7sjk+1o
GHrBO2h6WakbGi6moIm8phbYL6Lfg43FLwoFKTJKoXmmTn8JgMfq6Zdvplw1cs1m
3EqMi43arFKkKM9Flm4mo1LUBUcwh/r69tirxlaTAFlPrsaUP+Ckt9/R47LqCeEX
zcgEDpX4I9pVfxIQ/YNZ/0BILw28fejXl8AhYrpmnn+TK+8uSTDmGGZO5uFqfdJt
Iw7bsG2NFon0rILlN/kE/7pyKP6F7gZKQ2rBDZMwT5PW2iJiM0fknj9KWEqS9Wn1
z3LlbCnqkvJE/iDgEZ83jrjt5q2ybATcYWy7I5z1OtPPDl+nScIMhRpxeXj/d2PX
I/nbMv9lcXMttRQoYihpszP20d0knuRcmyis+uCpt+FTmedVj9ukjdmyKr/JDG4v
bncu9EwUhmze2k3EkDEGGy8VdwXBrh3piVEwQTgTCr93YDKpN9yYyEOQ5jbqQrWI
CDi5NyEYxB1ShKNGPTdkoQ==
`protect END_PROTECTED
