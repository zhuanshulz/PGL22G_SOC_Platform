`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S2C7qteyU9Ibhlo/NRHHPqgyq0G4gtZ5RT6yx9tx4ySzhXsLl1hr7dQw8cQhbV8i
ktyh9EPou2khfQ4ldY18IC2CZsxt4im2y8Y5SA8zNqAQ1l6DU/BkjfZegjiKbmOV
HeWpj8APMMrxYiMmifCGLRTWMxAvKjkI9naQFPJF8rPGgujoc43XBU00GYGC1cb3
smGEZXl6vX5gxVpV71h6FoTPX5YmLPTS7gHQCFDdhQlN0VD+J2kJpafB6FN2QhTf
FvaK/FlKSBv/fnmtTJWzQzOcC2jcPeIKYbEKZv0FYNQxduyq7+ytwAUTu12p5g2j
7tkeTp/NcFx/3QHhEm1K2YJaHDUKJ4bY4mcF3592CsJ5J9Z3nxAinyEPj0Jp2FQ+
NoaZnb5jqEFbTy+ORm50EwHvnmk5WV2bA+vOoWW8vgLuq3is0Ds5FKrUPYQRuCN6
AGRBWFnEF5UrpNPLAoz4JPwkJjk5p83SFZ1PcOxePG/GDQiqZ4JiWs4kEjr2HJms
iqiLfqtiRnFuKtvpIX5Ba0Y26HBqiQ3MWZs8gtQZ+WcuT3d2cFiw/CsB2nOaxZf7
qf0JPEL+DzF365tr7j2DRyfcFmKtFP9zlgMz2WBTRuLwItCqecB7p+ZNCvvnHto2
/GCWNXSpxbgGdujVLBnkEZCkbJOuw9HmYkhrvMjq7MrjSBRrZ4EXLIHiK/4NUvQh
9oYeMsWbzfaMi7V8gVzVWI6tMGeryl3h9y7OTHlOorhIFQdwjjNsaqTmRJdfTr1M
O7Vz4UzmvtFmAQPNuYl/Ghk2LvJcWyueWEw/xfgX62V5tJZP9SIE4y+IHpweN+OB
JTLeEGn78v58+YuazEQ6lDXAVO5eY8iZQGOzIbuXCPnugEX2u63yyk70TJaHWVvO
`protect END_PROTECTED
