`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SXzAqpAG9Fjcfbtzu3r89Thf3eTBfijPdOKX8Z6QOy1nKc09WMK5umtzD8W+9dhp
pRRzKYXUSCUOh3Hz0E9PgXmKSzU8TaqV8K5tshQ9ilYpWpP9ba4Bwtvm62/VK55i
JPwoPJJ1COinJhQ6e65XUDdFNtTJlOlinW/GZsGrNbyXlsiXIAXjXvTSM04/8vW8
c/mSbXtbarclBi6i4WuzNFzus+fOpp6TGRFIzZK+GOKEa4heRFsGUxSL9zkB9Yba
LC655deIvLYTdK8N5QpBCgpQo8THoL0J51+tpQ7yq3qYHLpvTBqF2ZIqhVe1n+MF
bJeOekG2ekLhp0N3YOfrF+0QuJNJmgSIX2EMsomCHpYCheK4Pc6NdResKrTunxQ1
XV0nlJzN2VcZwQz8CbIn9G4CrT52wbrPYp/+SUmZ6ftaITHzxUBeLm2J2qJHD/np
/dY6xDypiERVReM34mZPkeshfTZwAA/FISJfmCq7XlzCaMuUyb1cDQjXm2kSjPdd
R62EGisQTEO20VdDNByXXPzjqU+vc3LTh+ft9Bn5wqI=
`protect END_PROTECTED
