`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p567Tkyk+YTNfCG90GzqbaPOjvW/7X0zUxPFxyzeu3nWV8ZVYWrzE2F7wfRwWRai
7ZqFR4YERjBH76pTMovlkovTY9xNTMP8MMD2ujOKrKEadnHIU+/VnhmMFmQDU2Ki
bN015I3+8nrYKdCDM+iE9mW735zKHlXiVYJqJ93tmVJauwOgocWRzin5DS0D2mox
q4czQvGxVnERLd3X82M3LYSY7hoJjamSWVFXtygX+FOU7Hc7CNNSGwsORxq2J2bM
kX6EThwZdHex/AnthK6wpt/6M+b22g+JEMrIFsqL9Uu/xABIeH1H4wIjMldaVdxN
Qqrl4OJPL3d8FdPt/FYSmVBPXmwpDcTdgm6muimrnZ4vo/3rE/I7EpPabceBnuyA
J6loz9tu3f0PxO3dImwb11oJHh1dJjQ3SqKyrV1QnWYf3ThGi+8Uzn11obw2dHsX
srKcZjIzxLPutYHj6CO0awCqyyxBLZ5P8qn5wu/kLDIZVurS6BQt6CDSlStYKtxi
lytqGyiVOSzwchbSAZfOcGC9ediiU3ltZFVEdBUHAvb1ESX8q/MyNvYGEmKBDiQ2
wg3RBR15fFdBJ5DbXFryoL4onQPZYIEyxGpRNAxVUtkAfkpVArKSMFF7cGU9NI8N
g6cVcGJk2P8ls+ZFe07YUCGfh8iJjacWomdTFiLigT6+Tdjn4y1sFFoFwPR0nLkd
w12zVxI8Y9/M26NaWnNaov3ODzyIGYmBJr5hs0l8jLm+t3FDdbjkcd/1EOH4pDeG
kvCIzbwtjs76LUFFqDJop2qVN2O8vGAe0J73MfMu4OwL92qoMCgOT3EjfbK8Pknf
bwmXzMbyWArb2hWAwF58MGXCWrxhkT2ycD1CoZKUkZtGDmZEJxwk0aF/FYpl0yex
otSMA9OOTn65/x2hgRNHm1P2++SoKTU8FRKUZZZ+OeTMDK9QMxTunngdNbxB+bIc
xfc+s8EVmltJ/Gmx2Ao62RicpxfowlFaT0O6m07jYaaTF5X1YP/2TiTSqN4AqwDZ
XqNKLKI11Z04Q55531OI80G1bhyf2uwF8h8tWlZCA8BZS2l+6M9PQl5SjS4QeqiG
zak9yVUAcdV7VaEiTOMHHKumC1rSP3khiRHEsQC7zfucfQUIXNYPHJHvlDNw8VtN
8IlnWiutq2pZS8juNGiltQvlPjq+S4WSKoDf+MLkVMZEh25tao72StTEEhUbPBSO
RrSNWzCShHSfeuD1oCXlsOBFVES38U2y904G6eS5Abi4uEb+hRa2BIABQIKppMDY
GyvTnJUbDec2y+Zdg6x3QB4Gi9pmLJ1g9OKmPHFJRPeyz1c26w4Y0Sr5c2ftpWXK
fJTsFQOJ0zKsXZugaO2mJ8VQFOS9hp8s+EWWsQc+J01JUKPk9CNEwOaxRuVtsfvi
XJh1IRVsLcGOOdeGxlCuwpCTmEZ+9Qz6NJewEPhpaRqrZtpdPGmVOSJcHdCOvm6e
glufsiClyLPvn+Ih8x7dD0IdR0j/U/AlFw8mg1POi2CYWznCzd7up9aL3Cs6Ufjo
+00ywA3qkH1gLxkIBJzyKRiv+iAzZPS8lzhaDF+xITGj8HKpXgUZmiQVGQT8KKaA
s9pB1ttivUayiWANPtdPSNsDEwFUPkd9Pn1VdqvTNZjNmB4znK8B+QXUcidbwAG3
p3nlDRoyQa/2YcfamaTx/wtkVdHvtMDeKzGhFib6D2+igKZQqokmyzCCHhzgI4sM
mYJJ6AliZhTtCtMyTeb5l9R9V4C1jTiG9yMHb364E3/+vNljhiq3GmvqVcnOmRl/
w387Bt3/x2U7K+y5DwXnCBHB864UoQi5gUBUjrDV1OmzRfAVew9AdWIlAcIzYl6m
qnDkZbFDESpn7FekGP+KcT1Up/FfpQcEkUOiXXP5obbXCcq+9qIeMWFR2IU2sC5U
Seu9IkChf+DGYjsevBtN6sN7ehBkX/l4ejxm3PuQDpd87BRbILxJ+SHYJ6ZmgU1l
8c4dfzGfc3687DPApZX4525xmCf/gexdh81e90BnUTU/vzAU9lP8jCL3azGaWyIb
PV91mCwSUYnrWVgVic3hK5SlS36eHVkGtpRgeX5EaMgwjoxJ8xW3BkXjQyyxkeeh
4K9PPBe5hwtsOXVfKVBHQ7slpbZaa0+hWJMxBRHbziSzilF509Ha5y5FciebFli3
Sti4ZoDhwIjLjsr32pCU4iDlVZp6ynC/jChK9/0tE0O6DIGIbvrf2zYSbbCbXDNJ
vEOAmWgGGuuuBJa4kuayH8Jf3dZDiPHH4CVIclyvN1eWTlIkVvm82yTWKTotYC5L
MMV4GbWO59mX6PsG/KZWGEoE3rxh5pw63p3O3XE4zpXxLPF8u++xZ3Q/hL7Lz8nX
D3CdOa8SGqa7/e/3bdhvRC43pr/JJ0CI9wxAdNQrnCPENo2x2bIKTjHqkjnPxOqf
yACH4As9qRz3EMuTpSQojqiqfqwYGGko+xVCF/tHOHEOFsRuyF2yzwsFMXFg7qi1
3orefPu1PDOHUdok/BPqAWTfcE7v6IdC4lOfJINoO0XqWhDslSxL0v5OIDW2/f0t
x0rQ+29Q95zFtshplVB+3qRkGDIj+KCbywzDBH85hqANCv7Q1Qtv5XXLvcWD/Kxe
+o/HqFWRZ825wjER4CQ+lFPlWee2I5vmpifEifZZiME157nMJiSFQwpyedJF72nL
i3wiOf5sOPgTtAzPfiZip3YJ5JCQFrAn3z+GMRj9lAZJU1I8MWqThxixL7forPCs
pXzmnTMPvgW+AghMKDtCR+UXRkYKmvi/D94OXwkZ2NpAc6xFGDJ65DKbG26+CuMh
w/3S2A9ET5OD2I9cf7q2W/t0JWZg7DIEaqd96gCfuqBk6pd4yW/cvjsJGuiC/GoF
Y4/NA9RQyRWOs4GX4BfYi48Jn2Fo8NIDry+79fJLMIFZA1sVVsBV+2vyBTxLbrIZ
Zxc9zuiGNFT9Y6q/Ldefv16Zg+BjsRNi6W5m9maxAMMggIjFK3U/p+W02jcCL851
rfGsJKwt4FI+MMCLZmSbjmJ9fA33TnNd+uqY2ouQ37Mie8xrurN9kQ4nTLMWXx1s
FEXIVv5RoWz7wjlzA+hGejMb/+qDHcC/ozdiN6W7TuI9KzHpqRzSAvrMEw0J89M4
YIAW6CFfHE//VEcet7MzhttysRDQdbFjv45PLZDR0prPeDjcyCu7RVtu/W90Qflt
jGxVRlCOhupmzb/8hOqIoaZ3S5R4ASlxj6Xzpn2jxflpTgpucVotj3fl6hmMX1x2
LnCSA8nJpzO4iT9QFsRnJrcvqVwrevHjKT0l80I0QjQ1d8baN59ZRKGbsjCKw7Ib
AD7cq1VytNZHWUUdU7e86qWvYox/i9ll4glbvJb8l7ZfWtDq7lKF4lbxKlNdZZPR
K653NB70NNBp/ybWuHdfv6S1k67R+X96EoC87mun9RU+W2yLY2RHFwEgbdc7Y2Ua
+VbZ8tk8QqYtLx2b8EsRNTppTMWhw+PM5QctSb9NcxpTmwAQ+mG9owo1SeBQZfsU
3g5q7F/3MXJcWDejjg6NSlzpPhXlV2cAyVG/TcEw8EA9VxRZt35GWvtheQcEMT34
oB8YKoJOd3GQzzqwGmjtvQZYq5geZETtGUT1og4PmJ2p0qaq2mUBC8znhydNdMqw
taqHM8+TIOkJA9QF6YeLjRP0J9SYrXSrDjvpAqYlfARC1OpEFswATjHe55i7gRVb
+VobNl9VRROOqKMBJSl8BI4AuscnYLPGo8GpSTGskBCRF5weXTdVceWkhACQIKPy
qFv2xBoEx0tFINxcGVVRZZIu6TVEruAGrhNBQzItl1PsAB1ra2W1UmgXan98P4Iw
`protect END_PROTECTED
