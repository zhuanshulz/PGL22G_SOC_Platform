`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pI5XMaDzbm+5u+3VSFlWPdeKyItQCxTnB9/TtO4F8eBJhm0KeIg0cqgrLmHQGvXU
AL8xzC8T6xtlGbXQ9OykIRqX/NLS0AhXIEfRo20w7Vy/t9Ei24P+Tr9GNsmsJqbF
tPYSP2W7AQboAH+uKOZd6EvhUiCI2o9qwBng4OFivLWP8y3Xue0xTP91aB7A/vKa
6x+i65PymQ/UKKma3YVOwd0argTBrMp+jAbxzoggLELjrfkBJrLpggpEb1Dqd4RN
4ObJSAedlDdzGY7lJTHqpYC3nWCrxpbOhW5nBG5Ir+tomAUUvNX4o5L+Cmq6JTIP
FnXirCCKBcBL2TIBTL77hkXyqNs2Lgj4KYq8uYsuyAkSl7MIFLSimremljimfYxg
dB/qGaYNwAwLZmCdvgsbJWskBSf7Y6znQnsAUowVX0shndJxS6x9nM9f2XTJGmeT
nYutrRUvp+joajIvCGvtSiUtG0UKg8ed2cFp6oR2MYInCOFh1ZuOu6dYOadJa0kF
LbNOe3639Swi51pvVLjcfwFQAMzbb36ub7gE31wiQudSN///ZSqM1YTDB+8HHnMa
OEaZG5ZrPLNZKyHHHn2ZhkHOBTXr1O2ICj0vxfgJjXr8ZldxkXjhSSw8bbH9cXdJ
ISfmPAIx4hDXL083C67BAk8S4wOdliatZTpgqbPDWx2L1hd0DIp7OyLAOfkZMxcT
MWfJ3XBxLhuZTxs420uWWCEriYORDR37tMGsUhzKqCQHYFxvy6nfN1SQDJhNRP3x
3rKCanBISsUuyQsAIGV39nxnAfcDej2pr1oq0S2VN2KuQicPxOERjTyKkxYXfzVi
9OUCKCVbQcL0o5J2PzxYedQ78UMypTVvyE/x8oCpTQOS+g8FtPogYuV32XD46rgl
QuaaB5MMI4Oj0DoPIqduAZpYgudkl5kJlnSkijFnjCQ=
`protect END_PROTECTED
