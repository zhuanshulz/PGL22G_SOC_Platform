`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zSUJOUeP8RP5cU3ExyBdPivBKVflz4cbrFfUv3GyodtjGbG18fWKdgHzG1ak3c5d
o2vHpfpHOoxjNByMAGjPcFTICggsq10xKGePFNxOuyM2Q01tZtvY2NI5QUEO2ia7
nycZRQzC6fny1eAusVcBoLzpDSALsprh19sJ9npzY4RftBKsGz4m2yhKW98SLofV
OeGdVYKOpDfH7ERfcIxF+q/aZKvA9exUVgknI2b0288l9YfyW99EkXCYCoZfE/hf
RW81XrAE9/D0nUSody4aJaQhxhR26BOfly6qf2RWVZnFA6FTA7C1yUVpmXPsY3lS
CseZ4ZS20n3OcfdxXZ1EEbbTRUnKJP7ihKaeOHW24uFv5XFFzoQxKELfeB7QWbqj
wUZCPfWdoij+Da4M+57h5ssw/kfG9vLdDB+NBqqoQ+9Eki335LVZ3BQnFUhU/Cvj
k7YQz31zHL0Ln4oWGVX0zfy4ZDyl19Uv/lZ3VWhwfjbwvg84WH6/9mWiB0hNhKm0
IuWTZ73VPkt3UaIPDHIzQRWYCqZUlJppytKzy4EULZ8n/+THbfBZhSagsEr419pe
3e63UfzeNwdyBmgX5VnnPG/ZMMxT+QfKg07YNRsYBK8trUYYVQyWAxIXtFjrHv6/
JpEytl74qUnG5vlBMgENfUButJSKSuQpasK5ykeTf5VxFojIrJc/QQ40sMh+5Tcs
ToRfDFN9DEa8MpHN8oWoJteTAJfJ5Qc0py6IQa5FWkfYPfgd4MV1qvo69RbeIjZz
pjAA5QqHeDKk6Xy7akdCsE8jkJ3HMRYcqkC0urtQQOHv/UrI02M6J2BwMJDROppr
jYwYF6ChGe1gwiHk1Vdj6OSC5z7iWMgwr+G359JbKJ1HabrAaYmrxFWUWilABlO7
zCB9Kk8V2Q9bU2YbIby/OwqWDepFCopf+ZIDp+8fY5WXGC3wUsSZSgEowxK50Ecb
vxgDa1BNdvuVXaOKBAPlMpcamefRJHw22xLOZT2J3+4qY3n3rbaVbXZQ63tjCuIp
qDzAB9MAv+D3fp/Y/4ukgEo4eCg9EL6yabm5WdhFOyhkv24OpdwDWdueDHXDuelh
3t9vdSJ+tJzPiUkxcvFfBGhJ5Hz8e4QsbnTtvsdgwNooaT+J2CH8/rFrp4gozIrP
EJnpR2vUkaXGiZYYQNUZZPCY3ckikL7TBgwpl6UDEHIKQIMii0UCiMGb2F8uuNZt
heI21f11osg8sJ6zSB6Ihy8Fh9yBUFU3qEtp7KgcBKbjtV7iKx8UVVLQwl1bQOy7
ItbacSO6usGWAQzPgZF4BnzLhyKyACP1KjKXAlBeXvbv8Ms6cykp5GPhKam2rXJ6
EF6PVNz42j1RgBlcAYScjUOCss9t5uZ4AeEtfKN8UDApx+M5KRTzc+vuHQl79mfK
BBGLFbMf3qXiyR8/ORLie+MkMPaOYJ3wrkE2KEpZMatq0UHXf3I5jryJsg6e+c5W
`protect END_PROTECTED
