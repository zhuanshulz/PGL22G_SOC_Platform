`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
meSOpb4k9Gr9OnI6MJXgLQqNoG8oBECKtjI0v9ob9V6V22h4UNtIWlBc91paFuXu
P76MJmUASYc9dzgMNOkiZKjnvpSyoDfIbq52HYb+7UlLmqIGokIABkVr9l5rWf/o
v4Nu7IqWDuFWloU3nw+rel+7GbslE6Mg6lSgQavsKjhRyfpywWGtNix8gYNJCfZ+
1wVQF/Q4y3Aig71sTX+RUJI/s9uHgtPF0ZpIU90ikN4DyMiiQR92EgjYdgY6zfeN
f6zOy4Dbz0oNfre/qbwX0D/mXGYVQ3+qihyuxn2rC3L5rBCNqRkMk9GzqUrDOYqy
Mu1PLyxdHv42Jx4NNEH1QrZWLuRkY/gXohF9g0gLroQ5rRNW1cJOrpoJJQTD5+NF
0SKIOrypFU3Sf4tKBFEiTZLaWwrZDZIqmwLo0N3jZCl2rLqGAHurTpROcFxUZR84
2ppIOZeqm3UWvG9IMU9hzu0BTrDe9cUceyF8cOP+pLW76axxKb5dAOLAw/wb5LS1
XjfbASGdyfwZAey3UDQv6dh+D1hHdvOpvT6b9+8zEYer2kvRCPOYMrdPg88jX7Zm
XUs1mtl2cW09LaSSf+lwdrb3qMnFN+pTOFEPPhDPnk7+Y6sgLH0yp8OUi5W3BVte
xHKjuElDjbBDyOsYDS2FmFk9TX92/XxTFE6FfGsS9FdDQgm+kxCMvMnC/L67WYyc
Xvifirps8t5PXe0A/f19JhVTBIZBFDAzB5F2YaafE3/0zI8OM+J0yOHcFvvrUCKe
t8a/agYK4yXbr27NDikBi5VIe+Kxk6c6NWvYGdJ5HJr03WQMubH6G/i3qROyCo3d
0UZQb0cyWq9bizu7lXOer60fMI1feNvDZQ3+UyzMchHsJxOuckFe6h7yJr4Wd1uq
Ph7VcaxBOjtml5rX5w/5peLJkXsG4RUvk3L0vyhdVIw9bXxa8M/K477CuRDdhCXI
czhMPV2RtgOuZX7LBr9avvCjTwQ2ZxibTUUhic+x6iFe1UonPaRt1m/xCcxi6S5U
uLoXgBN8RWDcXDc9HG+c8tSflK90XcW5qGUJH20251HHt8Hclvc2g+lYgYHCV3/7
yrRym8Z7sJRF6jOUi3GzqTV4MlNiMDILWla7B8Itnttngj8LgWIeESEc+U9EE1Qz
bW+VNC/JobVkNbknCN9aC3IyRONJDBJeUE60lW1TaWWWMedm+rnh9RJ8CQQA/ah5
7dW0wz6coacC1EIjQbmY23+UYE/mAmlUZhgONWKfdnX3TinPMS5orPaq8JOEBNo/
8iOogFna4cdM0RXLt/jZGPrbtJ8cnhOxitQK8DQzCJ+jE+M35ruAJMO9ySZU3HvR
NXP916s3poWFJAVB2eMkUs8iZYCDWrfZ7WQDnZpGg8Xu+KxX8L6P0Mgrv/RyuwuD
nFv3Kj6/L89Sss5HZrUjC72RVP/EbQEWNBiFdflJ9M86YR1CdMRabj1H4yyt1CsH
bqDdL/UJ1FM7aS2AbPX+cwP7qDSR0VGusaqQv/4zF2gr9ODohhc45BfsFwgFJGCk
seiKv9GU994BI2EMVFLi8B9+gdfYTdLFu72LC52eRmbRtDI0wCl/Va9zmwv68LY7
ygI4MY2gYultDRICTESNrUkEhBkkute76grH0YcBg48NU3TZYOS2FcKjGkuLCq9Z
vn9bW9io8UGy1ddd6xQMj2JTZVjZROXYelyM35sP/sDbzCLNOgQL2njaYOAT96JO
scAPwD6EY5EpsgABFmHfT2XQ+Rk7+UfLlmuv0DPx20d+wJy4lttIUCZ4Rq0hbIeG
PtKPaNNwubxX5cvy+FRUdx2PWylYPobzDnfqXXLV1moMV7G36Cue1GQuVyaNodut
VYt1DNM1/dab+iF2F8Ehz6j7pgiU0WQxF8p4YunEQdviidKNH+WUKYxWrZaRHR+V
lqitbRtGMA9mWcooQGfoARMyLCLhMGL3H5Y+lMqzml1I7cI2LBbwDt9+67Qt5Ih7
9fV4jSfSsQNY47OPbx799mIxrbaSVQS70VB4SkJCP6E9slWxgC8uGkbp/+mgRci4
T/WVateJhYRTENW4Z84fg3vI6KwFwXgfKeVvrxBbIvgOtcfgyaYyRcze7W67kGNb
Vo/VpvcS009RZDb6Fxnb9DrL9c0DAIjh3FAm1JHCCKpWXnUsP9b+lDdsV0XMOGAi
pxfpivHg1rtx2YPbpRF4XIoEKf0tY86FBAJyltBuCuB5RBfnA1pWVvQBSE+uhUyU
CIOYKKyADTPP33vdUSnbmZAfDvk07+8NapAscS4dQgb1co/U7dRQSTEt9EEYkXxD
4Qs8NhVAHLEAoKFbCjQNoCnix1oEn84cfo2/ur2hgZz4VaUY5KgRBx0rdHbHq5WY
fcOPh7PYoRTsHEzXMyjv1He9AAof3S92YUAsuZq9zDeFcreXwzAlFRAJk/vNlTsR
uCKytH4+GZecnA8t9RCalESBkyQbHMBiTugQUhnP2BhBL9JA/q5WPe84g7H4v+Ew
0qLWsU/1APvPOZbz0xEyLd+TI+B6OUtx4kOSxRQj/YFEhKZ9jB6txRz6cCZTaMLR
QZ0qJVSP/92F2lQjhCa7VbCJ+QDvW1ZkZTOjpYwsNwfOIXG4KvnM8O4xBnmvQvei
UyYBp5El8NZcMQLy4o4y4u8NWmHHuAsuBIQo9uQQ9hcs4b2Wg7dl7IW1c7GQvkRQ
6DGf3M7F4aDwn06xnU7koWIprkA6KcA8kCfVB3fcIZ2il4GLoSExXFsGdn1Tv/nq
HNgs9EzmfqNYvfSs83mfaU5LmBPjtVUYeuXYkaVQVEX1kf2IVtoxOIIv13FYRcR+
qcLzc3Cxt/JHMOHZ+g0lu6mSEkA0L+45ZlZDu9tlolzUcs7bq0OP++Vm2JvRnpOm
KYDYgrVZ6AkNaiBZsLD79Y/rJkaTlln/LNg3WI7LlABGEbPil6hdd94l3aZ6E0KU
CETG6gNB273zzvQQvAlJs6Q+nNNZI4f2y1SmjYYi4f4uCUFSwsmK9UTwL/24wbi/
IVDfqto7e4gsSErNiuKiCKhSi2P7Htka7MqZ+FBa87ZcDru237Lq/2OUwsUdzkf6
3g0XMB6qzAxFgLgn7p01nZ8YeEAlzljIucgBD7PhffV3VamgWyx431fzAB+Xd4U6
9YoUeEDODfqhKFMKmOOcAdj2lPPInAeTN4WMwsg3Xn0mghvNdxCOlbB8G40Z25IZ
pXwiqR9dEiMeMg5KU+HXCb6ZmV1WIw3gaHPcCtj1RjM8TLnDrXrW0KecXAvhZ384
u86UjLEeKb3Yg3ixh2Oia5LcWsv27xThTI/wt4cPQy2zVN9ziTWk2DGHIEVPSi4h
FS4OST66P41mRQjylzsCzdgCMHaZ66+n62f4Ianmxm1VgVubIpQotOmFNwg6nEFy
U/Mdoy64LF4zLuCIfkYnssyVEiFBoKSVb8pg20mpa3VnbJ2rKKwnRjL/KLjOeVNo
a0NFsESSZqgZEcfJRX4bdu9ZpXexikhOBBWIu2HUcsjir656Zr3cEg+m9xLK1WGr
Q/tKz1nonpoLtfImYEapWZUXbruRp4OHUliR7C5py5Blm8jZEY/6jxXvFHhU8M1x
k2DkgzWejW7IGWvGjMwXYp8tRMd3JPuyo0taoyJgik5meP2VhHKcbsh+2TF2f5zF
Nhe0M6OXtDnRZzRV5CX/S8xs60aHMRjGlUNUPsjgFwSu3fuJlDTYOwiuBG87riRm
NqQgzgqd6dbyTDTT7Pgsyxs046aiu1XECsRMdDcoAijD0mn3byE25UILnNKa9nx3
AZ95P4HjMvyVM+Rr2IFAmYwCOyBdK3AN/R2m1tjj6wR62iEfeEZHLcxQ68gemWfd
dAj5KMp2lM4VV+k4XbZF/rxpOlcvXiYu7cQGIjLIRBMacYn/y3Se0rFj1CthL4Om
P0bubCKsPBTay98t1WlGwC6iPafTBkuY3PEWsztJOvWqLIhctg4dCZCq9XLTwpBV
/EHGwFdcaSYnhjrYr4QFCGn+4yYlUYmu8rYbc8+4Ez70mht2HwbytuLxi9rf4UDP
mhXYSeypJZJ1nufZTMpFcxGclcJNeZwPYtr0eQUC+Si2ud4436Enkdm7yyCYyVQT
ZWj9QLL6g30yGpV3UdcfMKXqOfsMgRX4KL5ggetvM1Kle7/F8jfuPxZLyGVg58sV
k3XlYbA2bwdh9IkzjPX2Gc1BMc2MCLWQwVLjR8rubYaxzXxI4Z9rimaDMao1KsSO
Pt2VfL4J/MFsMrNml+wX+m85KE5q4ZbdY/U3Yk5WIQbgsX/vQ6rQqTSWAJfM1ehX
Z6NSQfxOj2R/qqV2JOJzKu0/JpaxXDB44hBD2o4JX0rPnPcXePJXwcoUBVzt8QLI
Jh839gjR0HJo4R9GhWKqe0BrcESXJYe4RB+ZrlIaxZf3d8OAeMQZOmWR3qu54jxT
96Iw716kEFYAr8u/8B/CUeq6KDNh6S1exQJLTF00XwP8P0I3fHOxyk260N1HAgAq
FWRNRsq+uDqJThWuG94bwjWSEq765jHG2Kq/KPphNvaSi9Aol/97KNg3MJOxsyZ8
LGwpCoHUCH2iUGq+KNJeBaTO/pQ3svgaqWPH6B5obYA=
`protect END_PROTECTED
