`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PKoS4v/KsbjX0/zalSWdYXJIt6AxJhA+SbuIWA+XohvRcm/nEkf0i9PcGOfOm/O7
o62fdokqXKGrrTxIVhRN1gi9L5e4iIhcirRJWB5FvoxApW6lPiaaZEpBi/meV/2x
6o6ZAPhqFGfPBIljhWo8/tuq/+WCnmXWc+xvE5m1HijFqw6rdBTKPDq1aavPW/GF
qfdsr+iVdekBlAm1LnP7SF0w9NBlhWhQHw4vclsYB79eHO5OElaVkjvp7FgtkmCX
wOl5N02Y19uPwO/UvqPP3iDSZ3ec4S5aIUS/tHBK34/V6fu0rGoqhCHeNT8cIU9w
lIHnKZjI+oF7b7Ha1Y4d9VIDDNKku5ra7y1kA1PRdsoCFwmyEVxzIGBASNlTOiuj
l8iML7uarfih7S01yT/vzWtps+e5duUVy9puMMAQUZG9fGEqk3P1ZUsZGZMaKsiS
ZEUqihe9TlcxHldHRYnBhtzWxrNkOCkq61e2Vfpb7p5k5U5yOx67PFXp/SGJgAcH
XpR9ij5L1yHuqrOHte7Q5Z+OPbf4pCIOJMnJKJ9qX75rmiY9U/EsuVgWVckGLY3x
ENut4SNg0eZzFACHdIF8t/RZR0KmyU1ddvlUD3vMfkOCAsNgjsdB/XxONEH2Qpez
3F2whL0v91APwvLfjCc+Evtz1E5PKkBCurdxaQji7cd1eHsb7F9pej8h20/p6ENf
fubQKpdrROpNkhOzgsGJ2+jr3xRs3BaB+5KukOqhG7gE6SoI+nf1IwdpeMIrHD+M
wA9Uwl/dWfKjORzJh5ATiNIPhAb+euTK+V6vD00T8k2v1AB1PMBaES0Myg1LMkZB
UMI+rVj/afsd6eip67ORDWpJKcpA3ptjLeUYLX4aLpC8zMD+PqZ0YnVHFzZXF3Ot
xnYlxRXGH8yucpBoJQ9buojlR+8YK373UpGfltxHqa6r8QRoi6BmrFgv5zfm8WiH
BTUIXki45112dXmFCfuvINqnRnG1rK97zhTzQodumQup+bOsy+CUQeNzczPuYV8y
KSfBruk9gWsjZxcf75fd8656CV+ysCk99NVOacSwAwPbRFyW8EfaGYA568E99DXQ
gHO19k6agrnKfg08NFYSVBycrTo4+uGCaMzxLuxL4roxsuo/Kpy/gpwsLO77wg6w
z1D1yn9nKdbG+tHGhFJp8Ogk+cpQEUZgsyJnLHPiHIjcZahRj+kUV9c3U9AAcIKB
CmM8NneaRAf4z4clvrYr8xsc6uOpDM/bVq0ZHC4LtzTvOywIKi/Yh8fsfBarV1e6
Uy3AEllr19+R1256q/O1nKmpufmXKTL0HC9WsIUHmO+aRmU/mWcwhz17ArlJm/03
TUVBxNbvpuvYpJ4g70AFLwdE3V4pG02Mh27TO24QMS1ytsGMx4YIYC5pnVAE4t/w
mAS6WxR/jI3L0Z3r5OTo9POLAoxAcAXmGov/7SLorzZ/OpjCwBcRRipVVGhKnIk5
BoHjLmFhA+argQ/H7uvkqcQCBPBH6CsYKc1GA4rkBOQDshLs250a7qCfUufvTyZv
Ulp0Dd+HKCv6EHJyHZ1S9f4b8zDlaG8/qSvPYoNlJm5S4q0Rwrxx4Of5u5FCXnsE
jdxVdSHzW8NMe/gosH5YYmZ2Utc6RPVkb5dcAqgiA2tzVsX4JMHukspYpAgkal9D
QlgHPOpg2PkOnLS+ytKVPLdn8KCzjKL2W5M757FX4NKWGLs0dRN8GsNXsKvFcs2O
nO2GIy7qTwpKvYZb765gAb7kBok9UhKg/pUYVNn8v1DxVzMH0d9Ss/rOUeAH34ef
URl57yc6lmgYQ+blou3xZ7vKIgT4KHBozsyKo14zR73zadVUJef+rgJRd/GTybN4
+szY9wf6AUPZTTQTKoc8Dsn9d6dYojQhUMzTnZSgEoYUmkdNR4YuUSrg/ufepZbJ
FTSTZNbwWi0nZWDHUntDN6WNDIxv88LnWblhzJIyyItutO2e1DHqCudAsbFDKZRm
nd5pyWBnvEjoApUHRyvPhbwB4gCD5X+qdZOx1x0oUX3V3xOQS8WyFkikRqxI1GjN
jVF4L43sCO2lGiJq/fu0A81RAnpJUUgjf5JlTja6leWnglkrB9UMpIi2CMc5oLbs
d1woPEu1O3kiH1EOW+xCEZrPSG9jhnEMagOgrtqXTrekXLYGq2WFjX/mCNFq66IG
7sv14A+w1A/pPFU+8mKbq7+1wVLXtepYeb8bmA5L7kvyfjGF9pKXobqiltZL356c
cNiWDFX/tDzZCwv03HjDU77NoSIwy51BRDfgi+BDGUHBxlmY+b34scbfuhFlDwJF
VJbqtefuovHZk6CGD52x0ainBsag1k6E0vWBHQjy/fb+cqvOtSDH4gzb9HcNCnEh
wSROvZN9CBrrQ8dv0ry8jODTk/nbj0cT6D/v/iEt5hDZCnbLpvprbSEzCJ8Jb9Va
QWeRfdfn34X5g1d7MLXDbo5u67rMaURL7dUAwogXKm9G/Nr0iwpcrxIf4pygHjYy
gGFFcO99+cbuxlraE10P+w9NnQHEKJ+yFPgOE8B9moYtM5/6G9gLrEnliE16ADRf
2UrsMCs80hmLC2BEB2L0ZFRADhxkSouQ5oU+CXfnNgz1Rrp7yDqZrDYTDq4Rk1kW
vhmtdBlUeY9AM+9Jg1PHm+oEyT1As3LUaTrgzak9cviW0FJ/L5kx6Lfbzjlbtn0K
3BvRu9jKRMNMZ9CTrQqtFNV9MHpSWowT1UZmheTQbeYwgLVE02oBEtLnH6JD6bTS
S9kZholbe+F2hEqLJ1Zr6Q2eCuUvs5IIWcf4Q/j+VKL+IHcYJmLp2FquuYdh77kt
zwoFlVY1ThoXejMJMN3EVOS1KzIUbp6lS8TmhD+1o0DR+nibi3hshHlk+jGnER0W
LtKvDlA0vU+jgNJOnJ03xlYKXHVf5g4VNy+3QOZL5ZYbtKkZF0N3nBkUrodKBXMJ
7ELS71qx3FVFk8w+G1QqKmmyDC7MDq5YQJNDRGUrleHmfxX9ixkMsEf8BriVnKdi
4vLyyQHD0YGLCVa0NrnqMGjvUWQbHLXaoL5Nbf442pcAS4JUWDH5sFebhLJMT6kJ
F/HDUz4oEEQO9GL4OtyCWBaXwfm54Izfd4yjOMlwx2NajUiNwRVU1aCjCuLUMfd6
8vIWN2vh0LWZqoEuZRt2t+7nAlO4oQwsP+PnaX/yW8D3/1iAjowGk36/bEvv+9ht
3VbX7Bpw5R27jzGd8WIvEZwcaBmKQ+tQmIzcBuPbdHHeI3WZCRv9Ub/4Y0oJpnr0
uA+EwvZjMQBt8/esY7euPq9ra2/Y9ViiTQoEO0EWybcEbc+QN5zzBumD5rUsIWgG
F2WJ25jDmEh1iIHI/8GwCi9SpiG71koJbJ1W5RtYC3B/ncbIxZ+pi2aH/Np3L3nm
DHTziVH0r36iPkC03jD1yAl9K20BW/oigJBlK28cAQd437umLyVZMLlw8vZjz7Af
Q6toJGYGUqBvx32dQR9u9N46+6Kmao4EDPqtAXOwvB4XiDaHXLtInG3hmvmEJ5L/
3wqEdvbVXdRpngmhd+TcNu/KWgg7Mh8V28Z7Mi63mwwpkSE9kx1EaaHFEXr8S0Ta
2xGFSus9oNOeHhDmKq3Ek+EsEUFJwLyLYXA0I7GqRFxK4icJUuXylA7uJvM7RMy5
G/a9FQD9B8PnKLoahnu9gDktNq7TEbmNA/IMjdUrE6mw6ji2b7uIHyzxu3EYFVhb
hM6HbRYfOULGyzwcg9eM/QB63eSdaB8totZ5lpPXgfWk6KoUkgOaODxwZNEUJjbK
65KWCZuWOPg9mzQjZDpgfTzAYO+LeTzpKtG/hyZ1yv1PTy0//00spgu4jJOla9Dt
0d0D8TovXrc+7utyi4AFTy3IgERob0fcB8KxCbjk+NQKfizmqBeqIz3TH135Pqio
E0uAD5q/9l8xnKTiva9sglzPQ0W5El1hq3risJZKbAe9EYbl5gWitwJFJ2F/RlBj
XE9dWayQr6Pk5RZBcSD27PvNC/fO57WyUKPdDX9TSIOBnefkgET8erdjgePZGh0v
51QNrOiWAonU9smZ8VbeZqTuP1F0Gl+2fuTOmZwg3ZsF+IyCBpSIHubpj0gmjEoD
I0lnOCCW+XI/FO+Afm1ayL2Mi/GF9upZeG1yFvr0HMS6BroCEmw1AieEoMXT7V/v
4lN+235sNNg9Pn94svqzhS2thsbX8QNV08sVdn6/Sm0khEel1GMSyTYGpNO3Da2b
e36c0d8V4ZV8odZ25VOeb8hStwiEXh0BslfnJU3bRMca+Fy5acgnsHxeVwJuWb7i
JJswfAMT43TWBXJJ/lV8unFL16U+J6n5FC/Q0auJBJeRkkDRfJBnpdWqZd8tCHfp
VT/+ARWWnnPMzHANtfK4vZuW9a689SRfYLmK1vaHWu/ISazDRW9J/I7ZSLyLfUZI
W2aiAvFK0YmV/Rp5HrD5TL5xWkOpMURYzTkLpe0NuSu0SqYnGRxCZzQ1KT1q4gBO
VL5gnLK/DxA39NnsvdD5pO8alL7hjJX4ZpcY38VQ/JacXCHoZR7LNuYXnp4dB1XP
aPDc8443NPFYER+N1l4IVimb6gR3cu7yIUiMeILw9fbJ4WU4iPZCq3Stdz6n+nBA
6XQm1E61n6Ywi9w391ZhE5AAQygimTh97hUcOgPRYBmbbZ6k6/GBLoolMAGQKsAO
1yP1lM6CJ+Y+nHqyp/GFMZIK3SwRdo9AqlpHyvwJkZsZqRCFB60yFhjJc1UIBewe
G0ZVvIlgq/bV/WFcDhZEdtstFPUJ9oY4zOWk84NqUiaGDo2lvZXWFMeqzgQkgcD7
aIKlKrBlJoEXTizFEjOYkxpWt3/MopyaLPGTP43f9CtmuIolzWLCMdS49xwF5Ngu
J0icGE+0b5hAZU1ui8HXU1b2aF3+Smo9UOQGr/SR9jI240deatc+ZVNdnAKpO5JO
N8KquBE0La9eeYSJ189MJdnoVQ9GnrPcq0NzXMYFuKG3F5PYk9Yc5zRwKxIaTh9I
cTwZLretTjspXCTGvWvLqDNawf+hXpP8OJdUwZA1aST1/AgwDb7OjN+6seidkgaj
DHn+B9+/SkJngsVRyMzMsmdfQd+8fZ82kMsCtyM4LqVTrzjid6gwpYZ98mBIKZQ1
jLpxSjEz6TL8jRCWAoLjHQ4X0uql1BV5p8Zp1x/dfl+rHtiNrWOQ6720gUdiBttX
rhQg36yibLCCUdotNyDGOQ==
`protect END_PROTECTED
