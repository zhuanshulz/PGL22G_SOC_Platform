`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u3BeNyvKO/XFoSOPWqWPDEXwaaNtfbAot0FzQZ9visrIJh6L6bgQk7HuviTNQNWH
DRYHqu5AXnAojZhabLxZ+az9GpGWzq8wugoWbPNnk7YrBz3RitrfIg6j/SzvbfsN
kJF4D08VNPQ57fN2DviJndsGHyBfIfw1s/VRkKWAkMNDWVZM33KNqec5MVGKuJZs
Cbg8oJLWKYXbFkg1ZRYrfttSkDwOQYl3a7zNcX3M7CV236XUUqvouT2V1eQyWLFY
XkVTeCq/5VwQa1iE816OwnNd0C5lXSclXa09uhuAH9ajsPXdzhZHaawDdIHcv6C1
20JUnsxtLILzwAG6NdOZZGDlCPHtABLoUvtXO/TtE5m9jNy2QKJv5t6srMX+2mIN
45QHrtqni2Rqk2nlddMEX+Fy7QBN4wjowTr0iqD3DD/CyLL6awVwUZu4n4TkxrpK
NZF62AVuExq74KH7FJ6O5DFFtXzkfPu6qMV86uXdjA5yL7lh/06JXBpUJvp1w7QL
EE1e93odepvVcnh6qtD60M/pvvSBlalvfCNfDxuKuek0H9zQgx/FqmgKLwzu/xas
`protect END_PROTECTED
