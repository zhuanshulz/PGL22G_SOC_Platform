`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CFXfte7Mo33uVSTeDfb7ic7/OBDBqUyvwcs6HPcTwOOElyftWbaxQnj+jJ8HN/uZ
v5U10v68Cd1uXylouFeeUx5ktew868FIzmBbtP8jACEkCD62UEMMSGqnA5qdHWp0
Aicad9A5SN0JRwkwMy46NOKDsHJg44mHJqxG+6++m+c3lis6E5EKHHvS4n3ckNFl
RyGdDFn4bxPqTTVEVSqQ+UITGto+a6+hahkRKt3kUSZ7WwPNJYFvnzzAO+ZHXyE8
XVPqzHY8LFxdtVyzhcXnNsINDVFMKhZflIuhXH8HqB9ffUh/x30r1lJmElZuW091
yGkhSDJVjjX+Gha91+6JWR7nJnXo7AkrIPUCT95pFQPk1/+E6q0xN6tKuQzEs4z7
SlppSX41JoDJahjg6dmeG5YxWZwmfk9uPD8CZlEayJzQQgz8/G5iZIgW64PD2492
7/07uLSyBxZPqMfAapoH+E17NTx82DaRCQtBMhvPZqmaF/bXzLck7dYrkDzyMy8e
`protect END_PROTECTED
