`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gA7zPHHafxAY++xc9vkc9iq99n/AkAQytNk/wMVMj+HOHA5WwXMg73ygt1HJR3Kn
U1BG0GNCNEa0EvbLZuGzzbJab5eCqBu34cizk4PevoPG1ep2+2lf3AvyTHeq8Mhp
Q1t4vJ7uHOHFK809obVhpgRSnckb0AhOoPxybI03QoGlBwSl8WFZqwBHTHObjsH/
7+oPUll3AVfo0rmRbski/KJHs7BDOw4/NRrqwSmR3QJiU8+v21RID5fmWsspFoqp
Ori7gTH0yFpsjhf8PiZpDWQvBMjkiJf0t4PSu5YBj8mWDVYXw4TW4o+J8+aVAPWP
dtaOK7YUqMhbHrc9Hht4QBG7Fch4pC+Utjhl1r0rA8KNhNhxPycKphjj2jRdr20F
6mb/k+4+ncP1hv2eIhSbF+P7hp9x1qULOTm6isIONMWupajnfluAPLNUsOmZIrqZ
Ja6PebyU7Izy5t2COA7L8xXTadcxFu1T5W8P5LXmqYCvuNiC4uu6PWyYvni6KcXb
xHvZkCcB65UijjiIdyMG4yzuviqfAI1cbzTlpdZacPldrEY3dSOqEKcfWu9I6S01
9QMa8v9PauVRn+q8OTWA8+KA1c0y6Mx0R9EPg58Wjdg=
`protect END_PROTECTED
