`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DPSnKDZdN56l16SmmNhsSFCXhT49GpoSuxks22lul/b3Gnh2oi6F8WUz80Nnz3mm
tSHpYGqzqzh2P+kAQS3IrYfVM4H4HzWVIA7VjghETkXAMg38olfTrj454L38ZYPH
TdT/WmW1BuSxICkZgIXk2mzGbujRT++tivE0/97RFqAiEI0GcZzUxh9dAqp5W7iP
LY8yJLDfd6jbJic4WU7IMrAMg8MLBZHAiFxzHDULyx8GGyCYPvmllXrz2PiMvDbd
zPHpC8WKS22CqmAjjIpP2TxRzZWfXUc25yeQ3g5AvVsIeKH/WTPQXYkPZ/ekCoPT
JG5v4bPwtdqizi/sPU84j0Fc8K+3n3CPoChgcFRdm+A8RyHCx9BO/t96dZFd17f2
XxuB3GDEZBixrSH/Aw31KupMn/8ZoKq/HfEWlobiH24CihXWFWhQkG0kUfVeSpOQ
dcCw4sJptNbi8fzP0rcE5qNRJSrtPR1iP09mx6T1iQbSPHD9WKDlJavvELxdjVH0
N2+yfy4JC0fS2jpw8p19/MfV+5lKAuTEzjnTI+riIMJKj2bvf+ThyARO1A+e4BNt
oQLynM2AZ+rLG4t0TBGI+zB9jmuj9CHgJ6zh0HIRYPdIERzaSKOMFREBDdbpfTGQ
cT8KeJs6VGtFGrNvX9ovd8D4Bk1lh7qlgNdP4o1uo50/JheZ3hSithU3Kl14qsue
QTYWYHcKyw8UQOza8C1bGScYMHm/UWqFToQLKLwf37+LI06N4ro2MtRienWO9e1n
2fIaXbwjQOmxMetb2PFnpjsyrlT7SRXzlttqCS0zDzaRdrAwa5W5a5OlMrdAp2TN
jBeMNszTRSdlL8v74OlWRdelWeoPDy581eaJET4WYDMnwlqaL2R0c1WyskXk7QTT
`protect END_PROTECTED
