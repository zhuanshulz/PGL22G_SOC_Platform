`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t94uHYjSGNAzuLHv6B4RkopfSOItjrPULCOXTOii6x7Os3ldJ221Pb20ZzJvLcJY
niXspZE+9vVfCfoM7ygqCunlFD6lwZD2cQgXmu/+LGWKMDmtH+0PsoyvWvIQNZw4
dAZ7qo7ktkbbnmMauvh1ZCTUDzMzR3Cv2YcsiRVbau99WAbxEVwAGtpaKskY+yEO
SomfYDVrqFuPhUCW3YfylnGrzDSoYuzB3ptil2zdpiJtSMJlH7Sht4eqHhDHJYii
e3jv6l83UeImp2pcETSMXxSZlv4D6b8qrBJm1l7ja0yrFhtXX5xOWsyof/PMoyDc
RMb1y7VHwwJpDSvsXo9wmtkpJRD6TMh4TYtoV8ng7g78j35+GQAvHaZeFyDAFU3p
a4KI3KjPNw5DpQAJhdKkbENFJch+IG7aGjYccAhDw2DkkIBQKstt3HW8QeRMLYOX
unaaweiFr8srEL0HTrLrgz0HfEEnPcF6F+J1aeRBG8TyT0W6JIRK/Ebd992yS7va
Cg2E2Y/dfKhkL/DV0tsaye19L9FkhPq9Kk1KBcK0UjrLqc1fQxs+TjntUf3fIZJD
n2Y6js8ZDZJybF48ksxWMPj3Zuzy+sUS/55qal45eWvQdc94ee5lgK0kA5CRtfW6
ByWIzEq4KMAYKYnNXFigAu+Qcz7xic4NUSxyQ2LvwTfnH3OackuzmDINRqr8CfbT
RWB3z2sYq2/SOFPKKGSyQ0kTiA0KQQzyO3mbZD6DQULcWYUuTqPwNqI/TA6P/k31
3s1G+tff+6yOx7cfPyEa2thm977Ta2UFly8y6N7iSeG06TPlM8rQUb6ni33D+j27
HsB8zCXAKunx+ze7O8LrLvQbhDtUf4ZUsrxBYl37czECfxZVu7up47A8afzezOF+
aA8rcZtZyYzmr/uY81DNfbJ8dGYT/JnQ7joI/WU8q3pZmq7tZgaA7Xt49qUzLzXq
WpRoE/9EI5n25zj3r1maWfK1kxXr0N4fWFeMtG8KxnnpBgfZgpTw03Pdu0htmQw2
3IWgAUhUzKNxtPLEJ9EJ3Ptqc33170zSbfVrBSsOf/qBoFLPtS3H51AzPtxtvd9r
6r6VsJ+D62yLoBRRSIrNbShmxfU+wPucSFHHiUHi65Xb9Us1a1NoAmdsJ2lMLqEk
dOy6VeAMGGnNRWj293Euoi4AJVMfqoTBzzH85raSPOgPCZ4X84MzD9mOydry+Bqw
43yctHcBoxWdx+R0mTiP4XxX9DPOC0rkoCsAbq+CtG0+cGwCa95tt24SUvF78+eX
v7BTrlntvWv+3gNYvb0IM9/cC+3hv/paNa3JNHr8azoKZec2MWf+PB+0+3+JiAfj
E3c0gh+UeXFVB7asR2Ui7AV5pOxriiCKNAYzqUqi0pqIoMy5TK2I7Fthi48ygiNC
5nSIYP8vH94sX7MRkrxnWuKGXdcebYLHOEMwnvRhEFZY4G9IFPN9YBecb7rcq0WO
ijj/tcm9lRCXqViSAbK8t2YOxd1RzPQsMUILgFIpgHpFHE1Qy1JpXLmfNJjpRGVt
oJuguGcpvadjQywj9X8BzytlifFcEOwkf32X4W2GCTwP/LHsQQxFdJRULLx4+2B3
NrSI3h7FwAQ+wCPVhZCjATz9yP8VzQQSQO9USdsJAD6C2VNvWwq4JlbLAM1hsHhl
rpnmKk9kdqOZFcOoknwLRgTdvMRROw9nRU/xjJBow1RvQ5+qZRPMVKuqoa61zTfa
hiokAzlGsiZANOH3AFinevXYZ7fKvx6rNB7TVVkM9IGUKB152tRatqhxCwB2xb5o
hywel2/vdeBiCwvJYsfCVJ0RgUftnNcM1fjdhqNYxgnIX07F6Zf+n+TOohA/n79k
6w9VIdp5Ma8Er3GWEv3UiMnLmWcVd7GcigFkqY9V9Paaz+H5g3ITSrQe1+8UXGyr
J06wxarOThyvgoJUOk8el3WaQcsUvTZX8cX2IqIPaC/0+FpDWzg0hYZoFQlhZ/3x
X4SL6qpyA8amLZPITiesQu2riCCew7o8VloL7JBOuGnmOOknI+mYg/wpMVyVXKiJ
xrTUK8f51KF63tr8Y0Hxaelj46V4s6jqLB2xk6gsHtjicX864JBlgwkhZwIS0LlW
vgeuJpegwOfm9oNeQo/1NE/EN6lVaJT6pwmX3ulRRrt+9CtXzNI09V0InqgwmaDX
w8zp4HOTaBIMtn9bLsiBEw4exAD8vXoZYVy2vsjfxuTC94gquFzmiCIsMCT3WOOD
M8Q3fSMD3VYjsvfgd/RKor/4PzUeOdm5JFqdQfU7g9z/Ghk0u9lHHJ8P8TU3ygfw
hmW9a1cAXdVcop9b3kNSFskZniaHVc2sgyBzeLVHka8kkj4/re1+VoxIkqkmJG9U
zhIjoLjob+Xloa8/1s/OqgrJPeqRl6WDnlNUkqqZKwaKDA+Nu361y1a0RWegZ6k9
JDJ4igOFxaFw2bOIlfxLdmqIes5xPJsq3Gn+3076wTZA+c/xgSci/FbSqpQ3b4XN
ablQXDVaLaxX3lJtQnXW/F1BXyyeNr+gIGAEftS7CptRn8j1X4LN+2XXny+cRtAM
kiJFJMiZJ+YxKGojAWzQQhP3xzFpLagewp5TQN7NcAgnFFk1EuuOzJZpS+ukyOu3
NsJIaznZXSQCKnQYePPspCfqAtr6/eKcWJ4WCv4RlZ0DhuQlrwcHkLGzip0k4IUJ
xpsXToxTOh1hWRvmip5ECYOOGscCJ8shVnFGqSYRHePFfLsQ0oskhrPlDEPRcfIe
rRo/VULWm05MVdzRovqaeFwHtOHVHsj9YgA3i9yfG8R/FCHdZXVUQj1ZDVok3MuJ
7mboj9ckc1G4A1KcoRodUwdmVCHS2dT31zt+A2+X7qxB/h2J0+WC3r7tUZNae+o2
triOh+73M7wLizXd3Okn3zv1z6UFkUbZd1TsonWkcczOn1jvmICoragpxMkGDi+u
gDeSImeQDEYV/lBiW3Oo8Q4lHSlKmZkRws6el798oVDdPxM/Joh1lb+0WSF9Ej/X
S3i+gGC6ZCXjPjVaiXt/HhrO0wwU840KApa5URYTmgy9J7815zr6Sm5GMXE7ktOc
ga4hwCDVBTxDxJr9Xke65Lpj02INSbelYvteNRlvsV399XKKpdoDSdysngqZPMs3
rlOiGJ7134EZ4vEJ6sDrL5qGhu5Si6BMdB2LbznaRXvP+OJLIRZLsIBKayHHUBUG
o0j8Pp/mV/r7glGxq1VOZFD4WxMH/AUS/lB1Sav5hejL4UlG0RwhebgjrXfX+2V8
urJDnqi1SN6uuMJHVk6arbyV/CA2d8NcwGUg1Wm+2a7PUniDHdYZkD41oLdttLJ0
YqEGKdL+J+SwcH4eJrjcKcorh7WYDFTjsfnzGaq0OZudSj1PdpRqFBcI2GECkopK
tkGnoCHBo57+5ip3HZUbqNNaywBVmz6YUulycdubpcN+IrpProMxcXfNEjd0RtWB
22k9g8Y4fxtp5rklK7UqW5/GHb7IwPmSS5x+AvU56RaIqvMNSko/+qNClpnhbaeB
m0x6loAfk0AEUuhhnYrXkwQ92tfj/G8wbKEvBEsbsNLIpLyd74+MmKElQBSJPyGh
hsgyeCtWRbKatHJ7IWI6AbPkKITEEylEMquy1bEU2Lk3RaLmWIkKz69NnqRyhkso
tvcD4y+54Wr63rcbbEATVtjHy5GV1/+hQEb4seuLBGeA5gkEnj/54JLrhkKTbPaz
sjabLqDS9NRzx9tsDalwy73zZ1np38E+oU+rLgYqkgJvEjJESTc0aER4DzDXMonF
8O2nuHwudF5JfIuF/EL6mtuNZiUF4GstrG9gfXvGiWu21YNtfy9amPJHgs1VhBCe
8XulY7aqFdOMY+kgkds1wMGfRkSwVgBUX41wrLOcH271YcaMgAmLorh7xqgixblc
Z6UjUlMH7lSCIR2l7awTBYEDd/LbrxR8ynOQ8dvCHzflxryt7NRWTAZpljwX2PWy
w/i+r3FEzpU5lS9D9W8S8zSdutywJpD1Ij4459BmpvzCT2trK63g1MFv20I3ke2P
RgAM+TbTcHxp+vMyDNQellGnPQgQSNQrpWg3zMxAhCNkEkprBwvntYyvlDHIqP2j
VYTajWx8zUq1JbiyM9D5HLPeK6alyNg08v2kvJVS/VQK5sgeaVpwqd2xh4E2eowa
IUZTrbeiyneJE56v0ep+OmUqn/dmntt5lOFA3gfIZVWez2cpzq16WxrWBQRlCYms
SiNdqSa5HXILVjJ+I64+98L1r1w3Bf/ie1IL5NYtTlHy7a4H5+s+QqZ2aufsuTxK
lKGhMWIZFmbGthjuOSXcQEbp7jIk/3glsc0knHZKawDkj6WOLYASsziQNw7lhMF5
rvm49gEwriPaaSmf+5zWg35NsTX+Em0CWWlPicA394aEgOcWvIeUiYgEbglp1mID
OKrS5KwgrTkJ5pKJaoRZQGvx9aFbMPnVzjuJDW6aVLHIcrkUXMzh/vhXoO9sOChZ
98mGscdffhd275TeS0wJ/rVG+ON+F+QNiVK2xpilVoRziBRnvGVq43VvKE15cuj3
0EhC6uxBxhcllN/ByR/xY+URWDobOEHP3vwgedIq/eWe6DBFRJLK32FVljB0bycF
ZRv0iXU3pQ9tkgNps6IyTG9upLAffm1RRO98sDHoTy4p5FkPbF86Tmn7hMlB29Bq
3QP81lCKa+/+GcqrtFYmV7tFUZL7KED0RtWzlQRSkFg/MIEwG8idVDxoiAbW97vs
UoSMKhH5zFFJ/HWAviwtZ6rAX7xMypEEmVgeitE2LtJO4K6/k0uW/jzCVw7HOMcw
uy8MESXQ8dF3ovV6hmiQzCD4bcGZj50ibpFch5CBY5zTaPoV/IbePflJ/E2cTSLU
p1vQu23tWYnMbrMwuyjFbQJQXET5cyi2vgcYyAa+LmwlzbEnuZ6XCUP+VeMx151N
Glae5sVhh+VoiRTMgV69tWqbgWyhNVcX8mVGjfZRt9g8jk/hLdPCw02ECvNSlBKR
FatdqhYHJC9ad9JqE4xYU9HoVSAWk4tKDQPOxJAcWjexs795NtQS4L6wYuYJMr96
cerczbL7FebEUBOaVmOA2zeHPEFH0oaeE9Nb+f4L4pe7IDt3jHABIhoIlJclrr/Z
fIYtHCYlRM/lUstGrRhoYzlbFj1AQ4p3Q3s/c3DJ5TcmDz1dVcsTe8/ylx0w7SST
i0Lzh67guHFLn6E4eqQM6mUUpr7ub4DNhlGYJjYH/9qZKxSY7af8xn/lLIsldHkO
qELWXd6Xj/uk/BNTzs9nRGVgQQuF+5uwprTeF9nr08rIizLPYCFhffMHbTZEHrvC
TK9j8UGCdRr91bKMHPuA34Pv7jo+4yXlsy6E5OAwTmjJeXby6lksmXnkKt0QXGv3
Monc4EoGA6Ig5BUGv5e925EYDupMM988PH5bhPCQ2vFXo2JpntCvLlT/SC3hg/+5
9gYFYHjW/aCpLainSS11AFaC4jSEOSoyN5Pa9tfPDV9umdJqB9swQaudGJ2WGK7v
u8gIoGhM1SxajyI+wVqLlIJBu4WXAJbuitZ4I3N5K7J+0rXy+AMT9FZ1t2S8xPkR
bOLC27b4f4t/EvFpfyHOfF6Pf5SGhAA/6/wdkGhGSMGf5KJQgdHh76ii1y/bQVG+
70O/lAHp95b7e90lzeBYuJKAxJ/qauOaWX06NFWZVtKpfMph2+etamTkVqHN9TVF
KxBCMM5CiIY8gmTe1ZlJzjRtfoZeDOFE9vheZMMX9lvFsn2EORSVG07prepvamjT
6FcYr8isItfPPooPyDv6fksJ5I41aB0SWMhx07fhqseAPwvxfSfn8xouG3lTSu9i
iGqxmgoHi6KhZ63qnxki7FojAdK1hjVA7JtyEHhUFZMbvroHvhnVLdmcQSkyNcbf
Ne46KWeEmVb4hDsGLDQ3QMGxNMv7ZmpwiwdyY1rW/wPApTdp4flAapiQ3Qn1J6mE
eMchV7JUPtBIRxCRu40K4FcgyThAVof55hg9NS5Vi8nltWUmxstqdg+wwfQHGnUG
2xmkRrOmMFy+rPu0h7Icpspli1ZM+AUmX+p6zrqvcChlO2BTnvFjlIFe84Q1RS8d
qOfLnhoL89T/0ZIQOLqQhryS/+zKnxknNCiOGw+l/b7XkhXEbb0xD626OWgTNpU8
r0UpK79ngnRzg2h18O9AhXV7xljdQuxo5d+go5XCzWHOe9GoiqJhRF/zszSLMvBp
ddkOuREZoNAb6yjxka6Ut0xb/N1lk4zKOXBU76VrdxqOYAdeJKxndDjH4Huhtt1f
aEsUKTXnMUdqTrlHACYNTde58C10DFHGFVNDZwFRDHW59Uw/p8nXXnii2UhpycSj
hRNVuLKTrtf8qh8V6VPmkDhzO5g4PieDds1vpCaGnAJOSpKap+6cPZGr/4ra/5ZR
9HKuuiPY7Veg504NUrz6mU0lncMjyGw1ylIMnhPtt2dAWtGO65rOzZSWGgz2dEf1
dJIoqRHMBbFErcayaUaxpFlqbmp0AE2Hp+Wn31GUbRMbDCyQleF6HNvHz1JdMQLH
wIycx/h9rdLw1zVa7IM19cZxIPsMGLlA1SK9SkVzzIDzrsFsD/zhNQqTeTLfjcFA
OLoFrReh6BPNUa7OPgzYgUqoFrECGx17nbWWBXaCa/clOsb2et56N2BnBCENMXwM
8/L/BzQWBRRDclMPhpWVsmD4tjzJBjhuKAjHy8hRDR6e1DfhqqRsQ2uFdJ9MGnyq
426hxP7N3uyF6dhmog2kXNGqisRJ8h/fkfYkeAk1OsgPDiTVcSGatqGFLY7gab/x
q3P79DSaWxCd22fRam6EZbptTDweBYfDN0uBf5Imwv+CHDzKGKV50vQhY2U4kBhh
MJKlAamgW8J+Z5DkcUUwc4aB7N5QaNHXPtTdkWTPAFSmNa1tzUec7xR1OXXcOhyh
3G+WTkTGDEhWkAeMau0R/XH0O21NIpjZAmhhsasb4dX3NXis8+HqiD/DmzEJkY1s
+yx+g04KcYJAvjj9DXwIvHwNKjMZiMHvBa3nd9NfLTNuyEfW1F5AanY6iRWpsd4V
I6OCS1nFSAk8A1Mcr4gAwfMzbWq2qAFp8R8pLMG9HCZqz2xXatT0V8ObJoNCBcvl
7D2th95W6FpXlJRW1/H+KOvNwlfZfuLcvzJVYcjupdwoDpXiyO9a02OavNKJxFfy
apRAlzbVNpGrEOzHqzI9fxDmthrnO6QLGxkPpG+u2M8gt53rud24O/8CU98GHN0U
6/ZRlVdZKjfRgHbxHtvApDc9z5mfBnVpe2g63w9EzCqP9HzoX7byFrcCEJE2ZGsg
kZtaxas0Zt6p4youl1GX5M6mQ11Gr/GOvLj8bD78Se9Z0W2hcYTjB9CsWdL5pO2d
UotnjPqLQ2Y6T9wQiWvfv5bLa02uoYdcxd3LoV0FBGiCf/KBjxGnBPz8CMt/rjZE
4pk/7phm4GcJkGVAex8CUyvaX0UvcDd7px0g30wQxI4dKH7LHkDyR0oyASfMmJth
oXjL3q+/kGMyEKpmpFCPKWXE+Bw8EwKruaxNr0cYa4Y8qzl5s5ur6jG7SaSgqcA1
4wcRGgYF3+PChrp42iNVajqrlSlvtZEU0l8fx1MrbL9X1JzG/Yvjx4d8Wp4KT7B6
1LTHBH7NBEAzMID/t3lhBlkRrd2127rfzcb3hNwMwHaXOQriP6oVrI70e263NSd+
YxQ3J3a3GFUA/6XgBkyzNj2bQJe5FASIDmqkR/Jv1yMqrIqGs3Af3mACvF15OLGx
hUvxRHk4eWeSAWriVvRS04PbRSFtZ01LdgbDEMGF30lf61ehnyaHZZoPzgMoqW4u
kiddyDdCYnKqIu4NQ8YTm4hATxNaC0vufN3bXJYD8tmwGvzcaAFnHJeTg/tfsz8G
ZR5owMUpawx6Mf0ZqGE/YJazCkNq7FiaTSv4F0uFU62ralUPqx7XJnF993VGFiXZ
ieSIrxjOhhslNIgHZ7GI50jBmfh9R5ul5f8jHNlt+KpBdlwiYz4ZZanN6lYDSoGB
vXbhBf0FAD4wLVdYLzG3Quv170MLBkjfQl9LNtH1wm/TFRY57jJHZgv1MKvf0Gdl
oKeRwiqEj65F8Tbf7sgf1U5pHqabR5C3Z3FSxZkcqW1XgSKNTJFJKLUsX+GGJrNx
i6NqIdWLK64hk/LpHs74ZcNbbQiKCja52JAfQ1wVsjEuKPS7XVGnmF2mlLx6Dkv8
RD6pgQ5nMUFmzFdeeTQnEqGZymEbOvgSCkah0UhxjbXMY+sfzyOSNOE3qDMw1Smh
EwV8WNHsz8YblMoHb5s0nF60o9ImvVPVrzNmWQ5pnv2guL71EHFoUcmZnyJ7LbLK
VGMXapnWKIpslZexCyXuF/hTa5o+cNeRSV25NAcnnI3/cmdsTqw+gAO2N2NlVQpF
BvgvMkgDZNEsvr8owv+X3FGEzuJtIolFjDDTUqVLuXoDxci+yWmGw0yrLukJeF3C
CTaky3xfUU0scjhISTD5KvogBdeuNdif7WVV9NCdTHqhfvbpqVKE9Lb/HkpDioW1
1h9B2A93wxLu/J9tSE8RcuK80NzyrcgRIcoqyn08OFR2eHD1k7udwmxlLG2vTFQf
C0+qHm+eJq0FJFhmuzTMoHoaOpDh6RzNii7x38riKrryZF6htHnlCj7Ky5XrkglO
108P27wWrUUVuWb/Qg1p9C6g9t3fMDdBMbyaTetcoxkSW11VLB7S+NHD9NhW/nZ1
hogQ2G8b6QZQQHorpN7ofFdAgY7M5VO2BqFqrExkrD3P1pAGb9FUmo+r5dlnqzwL
7OjfcXoqDF6SYsMSdg7kC/KP3mEb6jO8XJbGlzu6RWg2ALCe8744a0uGjNQ3xUzM
CGvjv+7t4pbOjylECUf8RoJJNryhVWur7t+rv2puFweP/I6HxduoEjDq+G9i4CCu
0ABy5NAfbww6JlU4fc7oePRwrTEGLS1JoQ7rVbxamHSU11xlC5p+8rHVLVSfkNmf
BgQqDTK9iTpxjCK9R1oMWzHQrrJnhUaSM38C6/YV+P+9bW/1eiv1DwZaj6AZZOn8
yOszxQhCrTwYf7MyGnv2dW5prK3X153m9JK7o74p0hqEUlPQv7+D8wYZ3liPBQv2
4W1vcSTh4RUMuiy9o/GccOgFxEX5by+JvctSWlV1p68Q9TiBJNISR0A4BxBfzUHW
iJv2/mImE5lluKXzMiTTFa53MV5Pth+Aaxeg3KhjYDfh6NWlCaQZWcPIBjqk0Qng
0LRjBpL5UVHdcCoYdw5woHXjk8U7Cq7NyTON3m4XRlB6W6RWeUR3pJcB71hnHvAw
Xi4FHH5gQT6f/vxpaAhszmuuYA1DcSnGkBuLTTKHME3PthoTbrA+tVCVTWo95XNd
cT6qu3Q/LCDrmPYOFBr4Zz/sQMS6upVPQKFjAK3fO8/oFladv8E/J/xKQOCnaEpW
X/7h6ULq4t62CQlRhkTSBA+Yk7GFKUybyJp2znhV21fqEW+vuIs5dPDn9pN1q0Hg
lhQeqK0uN0uWUQBabSKvf760G2XWp8QUF2xKhY6Qr7BddP1EhL0n1GhJ1M4EmXLB
OPnstPDG2O4aUItLKNZvABDPSH3v+YeGJKoPyJ+30z1jiNuDtUUi4ZLFqtS6rRrA
NQpmcwcI1KJ0sQlLv59CV4Pw4YQZDQyKRMKQw7ENzTz7cttoFa1/lvAm5GRXkqz3
TJuRsoreOIsjotrk6AhcSdU7LsbK9DJJ/Ho6gkvJBpYwv1Ng0rODy2XQIntJrZLZ
OvDKmi76yaO+JgHeZVP/onfQhnYSa/Qk0FImmzlD81T22bJlZ8+s5rvID8X5O1Lu
nANRhi3bLzJBBjz9TceKzeAwx8DnMuQoa3qk/pcQZ4Si1F9GBYclcxgNrGx8mTiy
r4FlNiMfVuY1uE3W06D3P/Bz7gGjy1F2fGdwTGGFDr1YWqKD0QZ1vIFn0aYUEAI3
RezHnFOtKKig7RyNY6fT+H0jMu+qy7jM2IDlfUXC8EzSa765bdhGIR4ICO6vKYAt
HvlWkMuYN16R9l7bZ/LsD+/vNqZVxMcdfqx4dtS5suK82Q02uwg/eGiVBxUHzT+Y
1SRcrF7ZscTscm6+UXMcqYHETrbNehREWwz7FO3IeOcyrRblLylao5K6yYZ/yRx1
UlBhV6xvDCC22st1QDS0D6iCQnES6M7U2nRucv37+ICr17yLA77FVMIRwnpMS1oh
ydmEoGQsfZSlSr06FA9Vqi8TYKD2kS00VuKTRCkKKg7HHMM3Jhib3kmR5Bh8HrAs
lJD+UCWgNDKHTRsdvzVPaCrgu02owTLvRIB7PR3R//9VSzyjLcFGqchKR8ONiYMs
9wzTNuvmGn17rtRICfcwlbx6EVRKBvFRnUCNFBoHc81OHUBe4SPfc+p3wx5PMCBu
Ah8Zp8fTUF3s9CxLkj/oXu2n3MoPl1+Q9gS2P2hRgz3SdLQzaEJ56ErDYx4VxXmL
ymr73/1yZ4WAmxqf9JmnpKNnxbL1LO0aEf88qAAgosdV9+PigSdCvhMDwfBfCW+u
MfN0qLczID2gOKA0hQ9ZctcmtqTfZRv5VDGPXUZEtkDKWFeJg3TnQPN6zm4JlMqA
Ypiik5FHBBA7JHJcIYA3XO/2OHCUdMm1qIF0GHF0o1t0Jkf9UIqfyldyxgPZleQB
dycKwtX+7lb44K3qOV+lKwYWc9KMnNXhvvo9gRZ6Z/nXJJOP78ymeC26bObi52ID
kF66xgUN1Mdj/GYXGqB+ugjbC9jr48Fv7ShuyNeGM45q2Ekxqusvj0DZNH+Izdtu
qNpEiZwufBH0e6cjF0KLSZe/Tiq1j+pugbo1aygyvQvT295q3ul/NHSv6PLOupKa
EL40/quJe3WK3edIJlTxSwj5IU7Z62DQvNWneXx+jWTRHAJe/2rcDVdXeZ43Ysmp
zW+3ds6ACmKGmf50PpcQlF0Dv5GDO9nNKUcX+ZMe7LbW0DlJ0JVShUKF0+FTWB5H
b64RGAqP1SzSlrenlbxD+bFwZpIP34GBfgBQ7snalA07UBwNAL1pwiRAThq95nmT
WzQ+d5JYmV7pEXjMgFEywXVRHakFfCzu6UWvfcgjJ2XUUanqptJ5Tw+mwKyNP8mr
GNL7Aa6B4EfFNO364aBgsqnXyl1i9ChhfjudLe7gAlJShcivL9GNjB2f0a/6cozl
kuFFTxEF8HjSnr6G/2pEr6OjoCVDj7A08Yx1tiuYHTk3RKxJtyLexxOzYL9aYZk4
K4pTHNbsV2+G+ef4mm49LD0vZHvdr+A54eo1itRIZy3EQnY4u+FKVBjkqHEsTmmU
HjDG06t8MoWpdV91vioEl2rHGP17pf5BnJOsXzWo4kachMx7zmaQHl0poQ5U7KYw
hPi1IR4ylndLK7kxytCGXlrYMyHjmvV5Bfe12M8g65VsK35MY62XJODMn36H5koh
HM2TGXQdpDEGoGDKNCptfncNbD+NV/tEvzw1PnX34Rn2M/CcmtUA32M4E6xJC23O
0LxtlH+/QrSWsSFqdMw/Pt+TBuAUSXHtIZ1PkpNdyEhVOi+GUPO3vUChH0XFIOLR
2p8QW+AzrewSyqwUfwBt4+D0yuoHtZtFbZtTmHMD0/8UO+L/zJAaBWBcg7NnSNz4
CfvdyKeJi6N08Ka7NN0ufiaGvGsR4I7gv8MaO7pkkayGsmZ2HH9arlGOm+R47CBy
8aFYfOVdr8SBU32YEQzO4fm36LaCghK/2jXQ3bWD3tud+LrVtdLY4dbxX95YwDkB
rPx6Clc5SKBa3lYGs5inTkeZLQBdIUTZsoqcTlnBBINF/qYbZLdhuuSjsINxp0Uj
BtYaviH19r+Xb+AyndsEy7AkNMAD+RgcU/0m8w4GXH6j4mAzrFY87s4R7+lkP59h
v7E46aja0lVaEET5gSJGiV2s5UauxV3iE3fD5JJPu8SNDfPRIOWfpElXeb355KBy
2s9iKCXCz1E4t4xiT07Iulu9K3d/HVrXEcM0moSjQO5/hLiACB+2Ik+bEdQixS1U
mCqH/Ve/40v/Jxedv8UqNmSXhLZ4pKQSO9PzX+DT3lXPT18waJMWXARCe3orPCm2
mnKPlAnR8pWBfX6rMAQIQSEmYKMBpkQRcRlnFvWEvTqRYo6ZUdNb+9+iOZko6IZf
DQPyQgDv6uhHQqAGT9yonHYlsgrxoPJjlaiCrl78wvBHi1pqeUBvPorZkIaZd2DD
/0W7aFgl8opuKeTs0T8RJa8woIH9j75gqSdJgHs9QeG6r7sHFvmDMhd4U3arBxzZ
qAKNxh+zHs8qKwUGHdsFCr+XM/qO57rVA85N8PfUPAmwAmBcyyXKDfUvxnmKPvKW
JoSEPxZUROhvN1RqaEWlkX3EMHVeV6MCv4DfsJREqqIksmaImXCRwBJ8VakUjGW9
xaKjyJ+uSRTyQgkVYoJobaSE5jSkNfIkK3a8VP0p3KAyFSD1rVcPU2NO9ZO0o2aP
5iHPMbam2owzo4EpEZMkRt+GxGp5c6SHTqtHmcQRlvmQAK+ngTnsDgl57xdp90lO
WoJ3LJJlmqika+QU2dZk0ExdODc9+3yBiwQ6fFQ1N3UO/phyz//kYQQQf3/ssddq
aXcTPIAstfT+Sf7b40+8cqFCosmopiAgUyww+F4nAFsaCxGn6NqopLJU6uF1ml+T
AePmcepzAeg797Pk+onck3tqOavzJVE3Nz06JeUsb05s839CRhejxljz0CoB0d7V
U7Xe/us4a3O3q2CH8GHN2tQdKXf7TLU4XDnKQQrHftZ7WrHUkJ3KryDrbTeDyMru
Rpdr4O1yNgWFgiCk2y4UXkVFvi3WSLTka93VQUZTexBE4yWp5Ry2YHZkvV6s9rms
O2YRJeQBgExvdawP2bU3OQq1VVLurP/slsSU/lpBPMGzRC9XInN0bzrUlpDnkJNc
KvP08gTlDgwZzO0qZBgn6eFL6P1PhbBSjzkV2Re4CToXDd9lXSXulUGekdDdB1NZ
hgMZWqrzDP/JTFZlkf+997zU5QEesvohyEYjr1BuCUwt5WLi0gBqwWAis+65+3TS
nz3RCRFd19v+T+fnoeotpiYlSLgJbO1ij4OMLmapO5Okw3Sc8aoc3EozSj3kMQJL
SKQ5AENd9RmwepLXrQkbWoZCyytb0S1HVdMNEC5GNSdL3PiPoEWdfagQWuG/On4T
+7cg/AYspeW1kBSrya95K4FmG66GheneFfarCN405pk22gDdmYLLOskM9rJPiBQv
sevri1vLNH+bFySnQD9zlO+oA0QptisQL5gLcq61gufRSx4qya3UwBurTLpHVNq6
+TuOLZMww5cTY35XFpWHfugz/Tbh+18VTkmV9ilxiUvCBUdyJhqoDV8myl1DyE48
TsOVGvYKeyOB6i38P/fdOi+hr6GPo1+SJfiJPHvcqAULga3vLcyjlFSPsYC/utMu
kyt9dcWb1zZ1s75if0is/5zyhEgue9sze8LcYO53tfqoVJhKWYoxAEXaPb2c+yot
vIOooFZML18Alog2KW00DWM3qL7BCGes/FaZ2JT7N6uwP5EE5USUAjVrEP7mUN3M
aKGAY7F7qVrbTLruZ4ZQ94Gz9BMFCzCpcQJhdVogey3z7lIeT4Ib71WUIvBFsU6Z
wIA+9PDKMwEyQ7RmhhxUW0ZG0P05yuyTtRZWrD1CcdmNb4/QJdShLOzkYpdH4AHm
+RNjmHSCicuG6lQXsnJh3LOYCYSG9//+q4Iwq8iUWXXiEoeJYVPuZCxGGMj8vKhx
QDQLAPiF/Wt1LGTxRB7GBY0xlqd5deGsMPYhgJA1ldLbcrdJ6P4kK0eE8ceMS1G2
wCQVXd3eqEW70kYKlLcQmXFUe80WFPULqbAYn07gIOxD8jKRgyEa9wKdrmV8KqYm
R5bIb9tMahnl+g8UvtcARlIMhS1kiDPF/tTy07EVttVAolFjW5jN3crhtLLjcKd9
iIBzea+90vPvkGaCcLosAjUsXsS53ITOa0H3h76cSzeLCRdKK/90FYpfAAXfJphT
Ap1mwPxmjErK9JeEkWSQfCgEd8K8XWfiQHV7BuyvhQ4UkFdb0DgxCdCNiE9Vyjvh
7GsjXL1nBILCLHYe+fHTfv1jhkOxzBLFRvVLku3aU1cyhGd2xJjRzVcBLkYHgWa7
DcC4x9C/zrZ687qwyp4wnHeR8J7MLVUN9QgLd6yAVrUDuDRL1Np9/5VeWxmVHe0F
HP5T/oeYm94dBiL/jnc3w+OOnwzjPqQUM8qKYDjJk+TWuX2I6wng53OZW2K7GD5K
FeT9k+FSUc2v5CVXba5USzs6IMn+ARWXXNPZDRtcgw8JNtOLhTN0VSi/GIhIvsIC
YWkvzwRacFxc/IhNyAbzSfQ7FRjV667/CkSzaBTDRi6Mx/6dGzlbbrMid5dIA38b
+GpdrWkDuwYnkUqKYaEJdgyMULAiEf52k67sqpebxrjeQzug3Y8m+j0ws8Uq50m/
2lEC77c328ey14ixrCSn6WO0Zr3pr5daHl91ubvMFndbqxzatZLpSh7W6FCFapmK
Lqg+9coUBmiNkmKGQq1rJnGj+pKoTYFlAtQxcbYaqcLorhPiFuaFY/dxwRaxCcQf
v3P35Kp7bvkKNRzhe3rRW07H+Jt0rfl7vV0yWIJmy0rsJr6V7zG23v0Reh4uSaNG
j3hw7nCHumQFq6UoP/FUjWQS3gd51LgBbULlwBqwho8d+VS3gej4VLhL4DjKDcPl
aO5UX2T4j4sVwjpX05/3XOMcU5JL6QvNY8v9XDu4HZr1twlCLuecNgpTlm/Q9Lju
K0BCMYJt4iJZT6+gBvFQ4y8paBjOQcZlyTd2vFLZMdR2fRrA9oMbuGkFq7GvyCa3
zccgdm0JdfUZ0NKhaOy1rps8Sj7y7MDa0/Tq0o+dM7C99shUrJQT1T7NpQ3DLMJ2
NE+LnY3lVNC/EvtVkilVD2rpiv+xGiZbpvpz+BKbz70aViOwtY+94qQJ6hv3J902
pAPhXhXODjQo1VxBazAgoE80wuA0/od1uJ+/CYAtIlkF3uUzP1ugJkhU8xVVsDBP
KOU2OMs8H9FzPLzJMxdf7PVZ2UnBfMXHoNoBatKnURk8vDXBWYYpm0Ct/AHeCau0
n+Ot/Idh/eIrjmxebswF1NhQ+bGUdYA0p0PwoAORK20=
`protect END_PROTECTED
