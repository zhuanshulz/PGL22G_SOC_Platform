`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uf7Doq8U23rhQ9AQQmHJVRifocAq1y5QoTgaa96m0/JfEcqROMNcoONGqsClAsxi
7g10FmFwEb9/tUxuYVK5JudbTN+5SHe/lbgTCyiz0g1fsgGbGGQkLVCG5iECVk3T
wjSj2p8iUdJ9BdgLYgVrsWMGPQ+spsHrsA+UkMinxqHF88ujNg1ACPoSOtHGwSff
u/9wYmL/bItAXA0/q/gHxbBA8jAv56BaArOv6GQg0Wjt5MSvZXU7ZFfMmd1VqdtE
RlKaDhyFpr60qt3JtmuJZW0X/m05HndH1L31WFuPiaecKYiG5Rya6wAd37nXDPUr
HKs+ll/Mx+Y7mfns9IoaGw6L49tReiErC3STgMvrt1UfXnicY7xZUxgu41g7QnwW
eYmHFJbScj8WZA5dI38MItR+Nn0rA+ECClSPPdcFbBKafmnZkjuxMXHkzkB1B6Nt
cppqG0D54exLqC9Ohb9t7IiL8xXSh0ATf5u0AiMg9RXncda5W4G+cMubALJQiKI5
GPI4pvk+eDB79C9B7hrmYug6r9EvUk6J3sH/KpzGKKisVmJeBkBZFbjAW0zPcPkF
+2aYbeCC8LHnWFLgcLYOqtFxQteH5ygcU5x8Vgl6Vir+B6bF6xT6slWsq4f/akNn
IbOJdGPwZChPU0hAjzO2m5VkezBbpvB80+PnXQELMcC209PWnge+13wCKH4IyUHb
1BynMuEV/E2FvUkp+2U5F7Svct5tpsinSw6qTUxIB+Q5i5Sv2UjwCdBEatrHFO+X
rMnw72yAVDfPRbWVQTBamMWB6wwhUZclQQbXF3o1dqwHgPLlcDXlKGRF2TN7l52+
82ai6jRyNrE7P5ujlCCwQLiBA5cGcfKjM3d5t2i1cap8zks+SRr187e3sNxi/0aI
qxxyJ4FHFVlVwaWYugtpiycUcGgL3hCeP6NhX1V+mYaMbcFnEBTAj8+QOye0OtCC
yttgykvhXls3UXwGZQCX2jDC7rCRR1mJx8OkYEkO5+x9yINpV1OZrYi4rlJZU9rP
vTTHWr9Z7QVgntEFML8GFvIcK8rRYHz8X5HLmeWDMCEZKGTK6pJ3mnPM81JnsrfS
zwB48C1XYydYNKIgZio2oTH0u4WCZnUykjlHrP+LPupeCPa1QKiZlYbX5R+aduii
KaCqlCq/xo5MtGuoZKK+noUCvumpa1OJ3+7t8BHZENiXeeRJbXzAlDIFCQU6VP/T
lpjELIbS9DJC0nVz6FsIBQnh3Guz3s0RpXNaqDZ6mfY=
`protect END_PROTECTED
