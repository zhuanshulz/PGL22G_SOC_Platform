`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eshC8C9/PVC+S6ZXwiRaGSAY/41OGMM4EELnr7kZlrmdSSPCTSwAfoxx+DadL5lP
72jsurbeJ80tWHAABPbaH90PyLjBIe9m9X3CASYmPVjmLM31bJysH8ni8zRtv/os
SUEpSl1S2xWmsPHfo/j0meUP3vZeQsot+N72kP8KSIaCkg9M22yWgtfD4g4vYFzm
K1yL5DT9j9KUAzCkSIrPaCriq0vBc1ZzhGnQNKhS8pqEcebQJwvAJ+O1j8+k22kr
QXgOAkXecp7kuApeajcmcJla+KiVJjBydSB4OV/Cn/B1YirwAfVLgdCgLZzkfWlq
/fmCnc8gMwdUidp1WtEYVU9nkux76bgLg8QyAZ5oPTFKXDLCNmutTtHoMgv7/YBs
j9EYZ6JVfOBjEIgJhuu7SLflQSbsqOXDFCCWWT9TVr6zyceadfTRYWo7al3cOTPG
+uq5eO1NPJ+MXw1KrReTnhPpsWOiyxxzW1cEnGgjJJFUks8ze0TVOGSrAvYKeeau
mBU37VC2zlz5T89Dm4T4ORwmQAj8KaZ2+lOctvFqRME48jp1XfZ1g2TFFzaFssFY
OmlsV7LRwTHNTFrMhAu3PDANnRl/Ckdoncta2LW+dNQ=
`protect END_PROTECTED
