`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5rsMPoqY4CIgV8yMJVucdCo1MEHhT/HKlujlPyNvfDLMLExkJGZF6pBHpOY+Uohf
0MYsZN1Bt86JuOc9T/ka81IjbtTxcy4nY/H/QOXEMiI1yc4glshi8NkNu7Fh55RD
CtDTlHzrxZ0Jbi/NaQ/lsoSEBzWS4wC6/8k3TIZ3eSZBGb5KQr/kuZekd5IATFqg
t9BPxPwLzbkEJMLJCjM5/sD9ZEHmdv6zb64k925uBSfqB7FiQ/cil3eA5fJyM1yf
q76orjXOae/SgitVQ9UEeDuvMTBFNZnZblB2BiLB2JOLAI+s2e1eHlDq1j5SLh8F
eweJyw3GllDaK7C9prPCxVTPFKwLQ+kQXEFieZpp8FtoggsuE+XmbtVsNMYimYl3
jr6gdIqB6c0XVPOmYjVqee5SsPN0Kp1FHCGdTuzPqUoE7TVl7rn4GZsiTkgNJzHe
YmCpDyyHrMNDrtx6qbGn1kPqRjnJT7NE8QcBvb+aBlLKrIiFOt/K0L1JSkcjAbMP
X0uEMPkfsQotQ8/zoW2DhSLJGVmnMl7h4UpTTvntQWUa05AYZf86Yh7VhEV2/vC0
eGwYsmf9Jh9j+IsyVWtdsWXYVYmhjcrR142KUDK3gL+9lIJqmU8BEw55i07Jnzvj
NaWkUXLJ891m1ymn0ikxsJU3c17RFxhbv+fXCw4PCKCRsh3N4TVRosm1toxjQRtb
YQExhkFIEDA+W6nDJKMa9A1Hm21WvffCR0r5ztWyOwuHduvjI4xkaQ1+N7+L0Bte
CqdxzzX8n8QOIYgwu6uR6TbbTsuOFirEeH/5URHNzcp8u+jYA5Ue9bcOJqU+rxN/
qA6giRJV3OzB5bx+6dJzM5O2ihPdjRyHAEGAhVdhSa2S0fTt07oGzvAB6mSbXkko
jj8irRZFB6LZNM3Jo+1EFg==
`protect END_PROTECTED
