`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tgn6tILWehPPofRMV1NQ0xEnXPyNdIpAWxDOXvpHiADloN7gnRX1WWnbR/H+tseZ
1B3bW9rC/vvFOMnODDu+ISUKLMPSYKWY0KU+SIu+LBVMXnxgooblm3G6F1+rc1WO
m5daVU0Si7nbUiPAQb/WSvywaRYTa15gZX6uR0mIIljPu8aQw8GIzbp3/myuZtdW
XNYKCeRAHWftOQovQxFJmRqL9KVdZNf+0MxS98sXnApMah9kS8AMbEo+de99n8yK
u2AJTpm0mtAsSxy7AcoQm2bqiyiL9Fw/0lH8AsHnujHTnf4jSspgP84+IknxAwBo
1M+mDkAS4voGQ/3pZnTALbXlD/9DA5mZgr8wH2T0yuMF4QEg1awNLtl6X1DBJQaJ
4fkoGjjuo51Fw3y2rydgnbu3TGQA4mLxg4Rvj3TYGiF/O8hTR7zDfmieG1cIlbeR
WoEO2MhBO/RnBsWPGUBVOny7ZyID4zTjJuSt5lnuvi6u3jRM4y+O9ga9ztGtgMfI
gEe+Ib5raXSM8Jms1guTg2HEtjksiTC6JWaBPvnE9q2WB3dnMnupgFtEBnx7ckOm
S7hlD5jnbtqX4Uxhy7m6KCnnUmyR8tgZtoXcDbLrppGbfraVBZndocukuoHmQ933
0FE7eusr+moP6WDqZcr2nXiSLOtZehOwlwBYH8JZ6lCxeAwgacZS2c9eX9ZC+Vu+
rS8kwzPQoREZig9bDPJ6GgnG0fq+zjl5hcY01kc6BWR0infOHHxmlF2qCoAezRog
Q4fjfQBQWE8Ui+mQjYG3emc7SNAx1ovJJhgdD0e4qSdi7jenA6XOLaYMWag3Ahwd
JHV659bQ8irmw7p1SZW/wVyNyYgc0Bjb82LLFhWjOJ35bso/3hptfaNWd0cEdblb
XVM6ghj37dBMMAqeJFQfW4PpqZ+NcfkSO7TicnYkDt+4eJvhp6Y5zKytlCy/gATF
Dp4aSZxog2Z7TM1F86qhh7OCRkHUe+hJtdbs1f0S/06Bk4IzxPFRsEmNaHJzW2uA
IzjJ4gnq2zN475DcZr03LvhYaPBPfCGGph14AL7Uk1NVTlZD/qL+434mqpws8uLJ
sixn07tL/RWpaDH5l7RInKVb3NtelIheW2sGr5Ukxv/PDXiimu/v4xub4puXzymm
/RQgC7QpKdWvOQhG4NkuBkkCQKc3fyB99416A4vGWglZNwJvmezvkHS1kOmqoWNZ
HOVFZFIZKRp5zGSA4ZCYRtIBZUJmBT4SuRQ94qkqBLETm+Rsgk6o7LmoZwukT/J2
4bIoXc3yCxzWCzsGMLBTqcuS/ZPZc+f8dyAshttkliyBa8xhkWR73XUGNlLVibcn
VNSb+PNQlUjvQCs1FmpForl4ALmfhT+T3GPj6YCCWFl2aTJ7e8V4mMfjm0gKbsRe
hFxkN9PtNSo5NwIHtKE98hBZvLaEkARENRIBrDptCe6k6lblgnoLL/xz0oYuPZOR
OQ4/5VscUeyCfCIuk4/DEXxH7NQ/mEhvWXLMIn0z5J7Ek8XOC3tsEzv4FP2Bv9NH
ykO3l9f7PNR/pv9eHlTD7B2oUy9Ii5ioQH4KH+z1qAlS7HAEBgA1+65AVTchJ5eu
2g5JCnnXtQonuEUBgFtyUN31FKlmHrFZTVX2mxeu5ZaDFL3uROgOf6QiXiHe0gDO
0FTCShgVS7dgUju8BWxbTw+xgcyw8WmmJXJq6qh+6O+47FXGABjoBnd7OIXvuQTP
1EufxERUe652K+8V0M7hXPBYW3w7AwW+5+a4EButvjekLoUysgVcJf4IfVjXKaod
uXVkK6BydH6zYxttq5GQkTrgLC91HpjO8lQQoDuI53fArMaDJZl/us16uuEHcbWE
a454/DDXP8DMgDHqTQ6sANhscUmUAbxaOAdrJUtNIAg7eBywJ34i9amZcBzP3GLm
XbHrgkD5iftd49Wss6IUEIUQz7GJgX+tn1U3cnD7YlT2AK9A2l3jfjUJWMQPYQIY
hlLw705DELGFJVmpIJ2+5QMaU6tIo6BbGtQg025+aOaTJxfC8oEL5owIe+Fz3841
hGAECn7Az6zKOGNTB1lzviRKjS1Rc3fQeiS89cfWJ8r8B3t3VpFn+i3mpWfb+/lz
v4ulLoNsdCkUrvtrphgGwAMQe71HnQoPtCPp2dDHIcdECxVKxPauZ+vid4+JUSUH
F7VdLk/2rpUUVIQ38f0ncDZLwDJxuPzuO7GD/NNw+p4+CULk9FLeRTaIHybKe803
rGd+2bq4QaoNzCizrGMxQE9wnG96RFags87kZq6unXGcMbu6TKxm46wsaNmS0xv/
9RIYOiESehUH1SvoB7Lggeku1UMdYVdyv5B7Ci3dBm9k6qEmy66CdQsPa2t+lbm/
1CfwyNQ2S3CcydkYogsdg6d0EHmCA8seu0GQdaMd/KSAB401Ienzx0q3AdwqVc/A
I/sWuJvFkDI93CBSgWdjPBZBZ44xB6qLmQpV77t4l9umvM1dgFppeUhU5UQV7vMy
fO+049qhNojyRM9cTASobyWWIoU/04X+2QejglIdT4dIkHC6CtXgFh+ab4zuRIlz
5GPEsZaDgee9gflja5naaOW27oh7PkIwneX4AkZMNlq10zrksSy2Io1e/ZuplpHi
gF5AFaSCp7REyXr+rH20zKgs+npaAaxirHUE67KEz5aS9HamjBFMIA9ftVYCA97/
5eKp2PPT2yoYbjZbPq7ztqA02qAPqUc71JSUqUZ7Z7apo02xf/pNm7FBboJcN6jl
WW3LPeFPkXInIXYHl+wboWnNlABONO5XqfaqZTvRnH8I5luLxecqh3w9+nCIfa0N
9z7xrM96KJ4idOJlulR/6BMlPRLnlhzKJd3Ut7jVHE+mCW6oOabXaW7JZkJK183a
SQfvEggELCfI8lfl7hcn1vEHF6kTaYa9OhfwSyhSTqKHAXiIVNuGv4Vyl5f9LwR7
Oapdk+O/Hrw3TtcyDqsFlR/G5qabATe3bt/QIpZuiy+jLx2mutFFyrsDQ5kAzRX+
rN6h760c1sAh76xg9pT2Lkqr38+mOgtKbBVUuCCmEvoprqk7uxId/wp+TjKQUPxv
lKsb5QA54cSq0y+5hWZKSnNtMX2HlbGfyMN5sHahmQ4A+MyhJGvuf/TkqN/9x6kj
Fv9UIaU5qyDfu+tFcICy0o3kinv271hItg8z/Yk5aUGwWxY/2FkpGJ2YU1JR81Y7
y39O5Cid/HBfc49R4dqfjETtnb5UV1xeEOwTQPcjW3XnADI0tTwqeWCgbNuyCaEq
rH/O3EkUiOj7hMvg/b46A6wlx5xYfqpLByKqJmuFDbpymdFdEtEd2YO0/a4KJVG2
7npoAoYEwLAA5VPYBiR2ApT5k4sV7gYdKxSEtadCiWPr7S/yuVL3JeaJVeo847OA
mXJHrbUMOPZcnz0AH8sUGoHDNCDxnNAMVdS5PFT4oboLfPbca31VbV3MYG72y/kr
axYC6kUyRupld8gmRS6nAspBqYThB2MIgQ634TYaLmH7ZAuJCASSDuEpeF+lnNZA
PWHBjYA/v8+cUsP96S1PHzSforJ19BH5GJNnJr/ywutCFhwpZlu1TGRwNXntlR7B
7/lDgJ5yERQKVcZ3RuSIHjdVq3Bw50elv47YGi0fzOWFXGeg6Gt6nv+y8hM5/DX9
uMQ5n3mKrLxvfFUgdvuREww7rLmXpagSoo8Xng0N38sVVAUT0Olj+fvK4CoEvSwE
182inKdCfTJzLSd1vQFJQhdIpYrcusEfg/71KuIVUzOkzdSCRZKcmk6GO/w3zRGh
bK2CGWGnCStCLmuGev+Am3lc7MuZCtUa9jM2pzobKJ3QkXKv5z32GbCNaLbvQ/r5
aoXJQc5UiY9NIFYUnUfHV73W7K0Z36v9qmxRguZBbKbCnIohuR0QjqxX6D7dKCc5
EFIi7AmCetxOMPuvh6mt8HsZVohPK/HrCWI1DBEaqbTpgm/RVu10GmzBi9DdjEe2
sOFVzcBIj9zqt9bCXtiuk9YcJacKNyv3O6UpJZJJh7SUbUW93Odsf2KWjucDKUke
k1bx1TPiemi7rE0p98rmIbboIg+FYh42jpomURx1zc+8Q/ssh66rXTbLw5ydR7MM
p7wgoL1mqg+9fOsslgsvM3KFWX+u9YabHAEpkoWkNtfrJ84LSHQMykuFtwixTKrR
m8zK6XjLdmksu3KnryRQG30RHd0/EBMrpR46IqCspQ320Ngcs7KFuaoqCSdFPnzP
8cjXZjEcP7LU8zoH6NbTKK9i65pVtPP3w60BUOSGvDUtSvOfNQDMMHhI3za7IBaA
4lW+8SygOfy9HHApnbAJ6v/76bz46nNJCk9ma9b46AYo3WcWoe/DwDlqVqdON096
nSgbDL0EivFlbXFDuiMWm2l1IkOcgO8qJsQcn8AqEq0086P0UW8Xk9X9J5WgbOBH
LbL1PRZ6CO1Dlvj7KRjKWO4F5cGMdfw6DlRQa1SH64kJnQ63gC9zXA1WIxPQo4hl
g+UCdwPexk6slYZOAOIkPsxMFKNEBUetVwq+puctrS2PlMXzCrFfJi/LwZ7tNrsB
C56g64gBKgXa5jXxxyzUfRtwkW6I6XEGnl0X08WwETbOWdLB51zbHO7y+Az3HbSz
zJcmndP67sS7QpwUVSzO+joEuBK0Ta8HfEA9x8AmiIXSUJOI9enuBoEt9FhJfItq
/bP65/Ngu3K7ieSYpYUIB8p0C493zFs+YjrKgX93lXflW1fkWtaowtazQjRTc9FC
XhbyzODbEoApqUkdGXWFav9BxxSrUn/dzVWrMe57wNd6vCGDzap60eSjQOVNPdl6
RNP/9FzV2faJKzm/h+pTTNfzLPiJ9J96v8ZvgKFesk9ADWkynvDYN6s6zuzVRYh3
WYBrPNk0Qp4VmH/HeC8WgLayP9yV43g2GqANhxythOKJ3oakd6n9wCVXN3AP9M7l
snC5ic2sqMt+9IzU4KxwiSlJl6gozZuHAuiNwFIk7JJd5gXsHy0SO64iy4Q68+lE
zRGa/6FidXX7AP0BW5dnmNpiKfMOgtxXpxublM9c+AatfetsAOplYA2rF3WoZumh
qHmgz6DLaOE0ywoCBPhCdr4Qua25wp0cKcCPbaYRlgjOcnbrR1KSxM1wOhRQL7iy
kxWQtGKqQ529G6d6eFAhphqgXqZBvwvu0sbKV57JFZU+vWdoGI1hNWs/XnP1Hn4N
uKt9qE4p0BauDQUCnfAfMw54FfecMn3JCK9nxC1zrEXn2ah32g7E/yUGMMIAYrK8
V80xGufH/R89LZdJIUNpL3mkSxtnONTzocP22xyhaETnCyrfluE55e289VVgwoMD
JfHFx9zeXmMdK9cm+G/CNg8QHG2ad4UziFSK5X+MV4Odz8vBrdpgtuwaVX7Cmv0r
iAHdUR/ga2+ZhkbVmPxryMlFh5B6RfoTLE+RCdui9lcqzl46qAxUwJZVhlBhdeEk
4thLZlUl/AJfPVsbrC87jYhw4MnD4qMZ42RUulOHJj8yq/xMKmSr+e6+6PuThKVB
lSnbSABu6HXPsLhyPeiBpQN73HPwsDY5rMuojikyLQZ4DREJfpv7qaQ21pC06uvd
fW5PIUDOt5KwGd3mxsKar5My1tMT7gm73LbRb3+gSqRrdzXmf0fV0FVYZoPN2aB5
v1QfQy/dFIPn52at3oG70y1X/QjMkCgeFT3JFisXn5Qvc4P653mcqS8TGfUVm1AW
/W50n3zmq7t9JvTVKu96d5mkRiqVnacNMCDU7xu4+IPRy67ZcgKxXC/R6MfYb5Cm
yb6aI5hI8upzej1A6l60tw+egYydNgXgl2Hsjwu52kCnivZ60p+nYh/Oq1Tn8I6h
iw0yJ+q1kN6Fp0t4uuU//ZHmQgd8mDnVJkNgNbZ0wnVeBad8v6R4dlYISMz0P/+I
hwjn7vYMM8hSrQoQeu6Xn9RxlOMh7JERH01ROemA7Xc2B5p551EHly42skwfOsPJ
3DxXyguf+DVigthB55S2Jm/SjJXVhU2DEleQIEub7rhfkNmixryXJCfK7BzSncaU
0kRjiNehvifrJGvvRI8rfROGpHkCh5f+VZ0w7XkBiDr8f1TqNsVpkm8+fLXvj4J6
+mRqsc8LUyCdUEMQ2Grr4avbB8M01NVPiyeCJ1IjhKHWPdP+WZYDVMaYuljsreMv
rxDuhSUL9sWhLWRfyFE+AeAeOyhpryUIEQgDUkueS0dPuRsocYiz6UEZ7uA2NWuo
TWQMqfuW+CfdonQj/dX/FPC388uCHHd1GDbCGUVHxVW55ruh0CtadXnqCUUhFhlP
PY2eVUNowGz1YzLGVh8joyJmmjUsJ4qMiQwav5nvZ3ttB5owzYHLqGMGets1hbhB
jw5qnxOEg4muXllKSr7jzsqAbbkWBJ1ZcmMLNemF7YCY1m//vtLw0LY9CQOq3TRg
yYi/r7VKwJfbuUBhytvvcYGnC0IYC5X/EHng5TxNnRQjE2ZAePsEU7N8Xf9qgLUU
nwXqV1Q4nNtn7iqOTgzpn3pXjS3Z7vP40D0TeWmsg+OvJ3ftWCq8eq8hb4fwvIZG
gYKoteaigzTZ54d0pBkYdQH9sed4GrKzFVsqKhZ4hSx3kVxV5Fcb0nD5oxZdGH7Z
dx75vUCW+2MmfML9NirPjeDWaO5vQzG4ypq+2ba8lXiAZZcXwpEN5fOnfQAJTeCY
fmYTUADongFkcsjOBjtzlcLUJDWSXST0pAU6WHoWfJKOhQTQg6dhDE1GO0XVMoxX
5n+oFMIJ9kM+Ab+OgYr9ae0i0TV0GraO456Om0hn6yOScTWPGr6JFu5s4RPAEqgW
z0akanc53nlHCkdwjWsa1sXy7k7/DadgftP94Fi95F8=
`protect END_PROTECTED
