`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tij2AfCyU5KIho51y7D7cGAfWX6ceJAAeITbNVaW64KxUWLWYkU2wcFQsoWHPFUI
+u8QHef5FORVgp1qgehftIUKk5xPwE8yHFfHj0wpXDKlCw4rUBlHnew9o1zDo82A
P1ZYm6HOXUv9ms2FWzP7VYSGY54+w5TRRAfin0gwx/x8cZZqLHVElVHhHA7onsbI
zm8YZgGqceMSu5tWyXhxuDSKfnFLHJRk3M3/OQeldL093m6qBgWx8GvpYyK8gLeu
n4UWC37iUVXIWxCAQ4+VDYdKkVg2YNDBDXyrFQDJd63G8VBmkwJ0O+/hMHmYiH5a
CpLGeBzbhhlCx/2ViBPjL+DSl74ptZfka4bD34aquYFit7S2yg/beRn9cgMaBmCo
23+fcVZEP3VZ+7dWuIG1iwcPVtOKwnSx2qF2ywvllEmRV76dz0NUMAmoJg64SvmX
y9bWCAqd98dDQ4XXaOQ1ITYSFLXJiXxf/1qJw2yK0D4X/Lh6x+91mo5B8pAq4R+O
VGtw4xki+XTk/tkb2iqucwGgQq1Qrra3luvdgCQBpB/sejAYg61SO72+AlCPInJo
xro1LiKgByt8UKp3H0H+Y4vZkw2VePw3chI9IrnDYOggrov29H6P1j4DEgrk9GTf
kBtNuxcQikAZ/D9UfhnRq/K0tFqYWZQWO5fmVDEkZ/Eg9ltDMDsl818zAIr0Iyd4
1HySd2aT8Bl8DP7t/tHMPoi6XcUFBwj18OqfGvT+/TPfPnPTBmNBnIERsOkucWSd
XNOECZ0hQNwpwCVN0VG0EBeTG+CCaJKbxGEZvnoKfCxEGZYUbhTaHauFjC8PoZAS
jtUjnf9xiGZ7g+GABZv9+Kg5Q9xqvDAy7Gz8VXUfZbWJePScquLRjdZS5iXSsyyj
beC8ibmDxqlwP0GcPW3Xd839co2yPMF7Lbh2nr/uhGuYrDFk3+31x/e914WNdZ2w
/6rB658xzL7A6YG8gyQl5lRkhiJ1ssqvLmG0iZ9jiWAi78yrPs4LpUJqc8KF8wUF
w9VGUflgZ+mdulzzl543VQBBcC9lggxblACA+tEbJjz2E/WcKgIP7lXIOaTjPKSO
wIaJMGhd7NfOTbzizcGdB8/HK7h3C+uD29YrEusUhvgUxHLYod0MtVHIov00WjAB
9fR2QEsG3clQSSVtKJA44C+mSA4d8bg7K4s8UyTj/jAOwimxdq/rB2eceXGI9596
JjlaCDY6p+ds/GYReikYvW0JhD9EzQMlQ69KvReyWFRkiAzU99263HlLUhhfpTNI
EakBpGTkBfG0p5PtN7FzY2EF2ZOJuN/hF70Yr46P7UMnUe4MXz52ZJdZKs/BHgwP
Pz//nd0DMkFZ/ziQ6vjvZARfjc8eTBQ9O6qR2WqXfnkHPH4HZnEI0e0lCt3qAsLH
hvswry3wztWwe3Ckgifc5G4mIRGgDeOAnYYzKjHVONJE9X7tbTnAJjqwjCDZI5iB
oa+V4gO7JJHYw5j/LvVF72CTX77zB92CB9S296RLqQOCY67qsn+i8Q1OVdBnxLkJ
s1NTHfXkW/3yUYMnnQVwdIkfPO/+jauOx2kpLz0e/1VmctHx1WNtuLM5Ig+b/KkX
H3QkDV4cwDkHZpsfBFON/XtIZKzx37Gypw99va9YLIuLZXutGu0CskayzXZbBwTY
TxA9wAipgH+qmadkHYLK9ej2tQ6sYP6sxddmf303snWI6SKmMcvJ73zN6+QfGUwa
EZ5fNdlnLUcmMc8/hmKQsONBNhUtojOPvQDXrFdjb5u9FgXPm4wfpS8MIfJ7JuKS
6mZUueeE5bLiOWF1W92GXh+kWow04KzRW3rg2VBOH3HEEVjWNcBcYnJ03df7tAwI
JAc0Yi3EeUi/DSTbR9RFaiw2NDF4YljXanNF/u8S8+lNt8hy1iGguzx9w6MbTCig
DM+jEUE2sIU5l2tSuoB+FCKAR/KfqP2+60iZKsYxGpEYnJ+oy8RCvLhj0MmH/vGq
c9DlldlrDGp4j2OPHMhjX+pzkjNcGUBYSAA44Xnz0572eh9hP6w9h1wHEyl4fd1b
8542o+fHQvDOGEQO+wCHKMUPelSmsNCvsnxMaALcoRAkrvPbakkobQElrA6fXMts
Pl3T64Oc1RutnZ2iMuz24C7NJBWqaR8DgLBidjc3HJ8uBx6BGqNmzuL3+iSXH7Ox
xQ0cKzaIrGn7+WSSzkDUDg3B9Iv4BiPEtzg8Nk2utNkS63ZjGib2d7tYtLj7YYM8
C9SWW9njylZ2uplc91C24rIXL1r8weOoNYZyCeDcN1/OcfxjcIrB5OsXLYR40Ius
aBd+u3jEuSba99OpnOYGT84DzGsuC0cF3eHZiT2FpvTat+FkBHfShZTki7zEAT0o
Nx7JD2xUT6RSPicYLN7jatQeBvql7+uUy2+DB3VUlF27+mCZRDD7Y2OwvxnhO76i
MZew3j4cyTsOxXPdVD1U3W5XC+UjfoovVD7tpI///+WHc3Ly/vtaa5eNOGOZ9V7J
EMcIEcnuDuI29q0hmd81DxcPDU3SybogNLLktbi4y9GUH2CSkeuf9JKlxKgt3Jai
A9l1CXnZq9B3nLMNgaIQy8IaSZf4sJWj/OVJjkn4dbcFprGGaE4Dk5RS0laGshhT
QsgyZGrjGghTbM8Fm4jLxDlIS4fwXdg3b67s2uZoWgELFRqkAdZoS8GyRTFJICzz
M+Z5HWWtTRa13/AC6YgQSTTp+K1ujjwVxd7TyGlQ/hqYLTKbCsIRAqVkUqrg5Igb
rZdfcP57spHkJ/goIxg66oTb7IeVPBeZG2os9F82npU2TKhkIEL/v0YvHubgbUFr
TV809AhL36t314WnyMdnxSUWb67P4ilSlU82CYP7Y0lTBRipUqxknbUhX9z25q0S
KnLz63E+fiRn0+BcghMlGWAn53D83RvdgTI+9nlZZ/jcXCTESL/acWgb7kRjODHE
DoXGAMWXl5tmm7Qj5X4DRE1tEVPaMmhEWrTmVcRutIBSLALVMlg/hF1LJckvo7m1
PyXDqk3hfGRZqec9ncfnUJAMV3MYnh5tIy88eGxag+n9cjXn4n6jYm8cb1abvBWF
XPu6SdjJop6zzf3Iam+mfQQSK9oGoGUqWOha8l3x9UMm0JsGXAgXq/1NLbhcue3K
sLoEcnsALy78ZunCKhDltSWMFgBwReZ7b4dkwPjo2CX82FmzTHEx1X9nf5c+R9DH
f7WaEbISX2ZZnrLEldQLHJjx4hbWyn1CTn2Chs6qmMcN93RCOLqNvCl6I1Gb/Mvx
fpnf9n3s74vEa6EgYRmOFfjVjpISffdj3Qz4EmmhkwXlg4T+qC3uP4a6CMCmczSR
o16/4Fp8u6XSe3wx+j+2BBZH4lwF3h9dOV8+AUqzBcM0Gv2kEawURhato7ydAMlm
rER1VOoZYJirLAC9vJFOSzGQ2K/ji5eq7a1jWXIqpTO8IMEqv3PCN9HrCGHdxmCx
/hRerYeGg+rSXOhTppjMxLlNJLBI2Y/npQOxmal2WIWuliMvIvALEaj1IEnbEZUt
o22ay8j+IuIl6AyKgsD9OTyVvsj3qZQACzSdNoaZJ4k03ptZ549XXHzwvSmvgTjj
piJW9WjK32TRwYHEAtzuM4Vu1K4ssfXFoxvkiieAymeez1lZMyQcv6+JyayFRTni
0dcX1XqNwvFHN3STNiacI2m8yd3f6X+5G7KoruAOP6fySEm9R+5ZrNBbvKu8Jkt5
yCevhKAHUTvirm6SUwj8Ksems8wCjqJvD+riFgLR+8I=
`protect END_PROTECTED
