`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dFoB5IclOfdpUKl6kkCQfZNcOsnG1GkD2rV4jxfmqDQ0Djf0e9v7gnhOX5Yn1Y71
cGDZ8HL88j5EZXPgWiR2Y/liLv2e0N8Dt3v0OHmoZZTe4GphMaDZngU0yvTW4yBz
46m3M217AhbohIxaU6Me6HYwBlsXK9yEyEZjt1zSPyVGIF+91Zt81YE0/Lu3P+iB
2i2bBclmk06C2vL+IP33x5UqwrV5uRbZ8mQA3ci4c+SJkaayfOlGbj8k1HY7x7/+
60CN4XfxP2MmlfEQgftdUC0FJZlOV30C7qDk1DxLDFF5tKJiOYPISILtnjvswQv/
1v4aXSe0wKrNhvAKZwmMUtEXKfvV4Tm07LdB0NTfcQvAgARzFn1lrY9yrMJBjBSq
haek2sOBNrAWx8NnrumkB+1VGu6zJSnwXI9y3ynZU5z0gsGX9dAnYbYDNCZwtbSo
XpOa+eo3cwrAI24s4yFcF7T/6MA0anSmrzBVJgcz/f3OJsxLj4tbx22PwUt/5TSa
NbTR9wdVgZFVTcmDHLvHvtVdZMTtAfPn7hY8bVNTAOkrVSwU92ktOJL8tE60eceb
CuWPBxpG48bUDWcUrpdUWMUbZiidRiG9UH3JY7vLpWiqhrkNjdVeL9kWl9Wgl7mi
s27ISe64Qinx/YQ37AETHdF27Ba2kHqjkF2dwGwWybcFmGGh5L59GflU7L6sKhTK
yMKIatFggkWaEYgo0MF/34EIyN88wq4pGyQhJnRg5TSaqFu/phQVJQ6RKERUR36Q
TYGYf6LadcAJtNvObpBQ6lGHXyv7hKgr/Mkwa2220LM=
`protect END_PROTECTED
