`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IivqJfEk3MlcpWitK1alhqBGfTk3dRthOG2EJFatEDtCZbPPwyWmljCWDLhHyRDN
4p3bZ9sTI9sthub5hbjTFnYleNSLTCNUKwc8+AnbKanToySPITZa+IKhRTlYhaB6
pkRm1dj2cbBLSfhqV00gusCkJ6r/oeNe4Chhx3fdCIDrfJetQ6JG6Wh0izSh1+z2
FAI2HyuJVSRf5EbIYKYn/Z+KLVszfSkiZ8iwFZZClsLbrN1wC0qCWF//HG+U3WgR
/SAslQyPkxZhvnYoX6WsoBj9qOvDE6e5NCGNUNUgEiITWS58tSGpwYu5edLobdho
aOjp8Srr7LwZK9sJieyr9g6jIJmWtuppbagxaX8+K5rdde8V1CrrNQNQRtgdAdms
a7X7h9lmYtvhFKYQry1DDKLhfTfaxkaH55vlFyTSfaKAgRCFYLtWVnVbIzUHo6u7
Dhf7evDqD5mNazg2U+6KbtCgzdbRu4Cg6ZY4AdqPqjp9B3m+C/yGaNM+HZivQMOZ
rb3fKuNs8B3PT6D39pIc+W2VCE3wx/acoATqzK01hl5304VpdPpbVxXgHmRswFia
7jng4PtGPVYCVyn2BzlgYx9Jy2NCDbqnQOV2OLXkwJmnZKDVhvvbrs2okdLO+nh2
mGPLr7pe9Hwwdx1p3Ss7MrXiABlj1upX2Kn2f/t7OWJvR3orw2377FpsdgtdA79e
VFX3T1oseojrM7RTjtM8SAXeH5sSdgk3eQ5GvITruFnxY7CZlNaWp26JveZGBphL
g9COCADPxgVcNL/sSAsaCYfxiV5sPVU1Dm4cbYRT46xAKfUpdtu0O6qiQlq/jk9H
6HXeMKw5+YjzH3z3je7QKCzhNoH70vCriz8jmjPl2xNvvb3xPO3PiLvS/VjMNy+X
HsHBTwo5rHUNkTCF7QVNrMoBEoBOYm9wSLpUBHrGDR0VullS3AQQCkwlDNHR6R2m
uK195p0auP+UcN34ncSXSNa9I0YhhrJxBI7UZDJVSYlOhLj9wEQoIjfc96QppGnc
/eTv2qKoc056mHata2WLhKgbF/Kr0CwtmUeYHoI/iVjmu1xabIgghiA7XJyZ8b3Y
A2nKttCodvOcSw6lHPcw4PBRmuE4BuB/nqxdQqyviPh4IBHvE1uhj2E7+Xp+/4nr
5Eyl/Aswyu0csSiBdkkJWvs2wSniWzDB9VBWgZ9Y01sFcuaksTMX5J2KqdsSrhJA
4j5ENXP561wZz295VqaGbe+UzOHQZwVmU1ljgTxE45Mgnsb7jaBcLndkK1D4d77J
+w5QLplWWFcc3izFApNNAlwViD8/hFpn6S+zPAC0It36rGMSl4nZSASomwjEoGkG
HsR5JouxpNRuNXPjAJ2WugQeNUkf/PsaMnEKJqSc/ckC8rkLnjxggo8T7/mxm3Rz
2smJ3tk5amM3Q1CJ3yph9G+bM6j+V04OHulb0hL598pTGQD0D2tWC6+L0h4Z4Ub8
N0bcQvLmZDA2tomIz3l1yFzv9fi7tqnQg0rGW0ZMzdjLuCPeJfVj4dVyhPWSAli8
Vzu/ZYrMWqSzGzgwj8QQwCxnmIaDzBAAiZcGT/1zwMCFp86q6m1vnvWF9T3LjJOY
E66T5DkMBK6wG7kcv7+d1ASIiHzuLs9QIeUy3ZrITOAtKHW1foY3IrLMwkNdO316
fREnGqZROOpLJNZ6Jb66YDDYIDfoEBvNfhRk+vLi99M2ApadLeAZJ1LZkmmM3r9B
UDdcfFXXURgsJ8VRfywi+vMrJDJcBRcch5zUXvUQUhf+NPZ7omUlik1c70020j+Q
8T+ywcPxTC6QiwMXBBZHqJwsEV2LTBGdjIrIM9U3MCtc5BIJHFopUPjR61dZsTf5
BmXEqQP05Pa60GJCsqQQizYlrfYzSwp3liUYUCg5NMyTm9Fx9FfSBt7Cn1WGCx5v
asQnNU1LvE16WMc38dKCmAFxVOWUGoF0MQsEekXbWhXu5l8r+TJsEF2mcO8d1Zid
C2+sj4Fms9TvlSuJrRwdj8NKwg0j/t+NYIuEGPm43Rj2FIKtxr9CdBDhtXZlGQ6e
M/rb0q7bTJsvIQL/855QlBlDgLYkt/quXD+jXoQZyzE4AI7z4O7DvsPacqUFoAww
yjYIioimOGdyNlda07I7ZUoDVi0LTaY+jZDWGE+/QqIkJOzb8Jf/wAaL6XCF/+04
mA1owGg5cFXHe0VlzZZvTlIuhpNg2D3gWmvMpcUtkf9ivkm9o39L3asFgECaz5u2
hszrsLG/3IIKW5LU0L4z+wx4EiydbXQ0WlTvl3Bo8iJqwlpU4wepEIUTkH+czI8h
3EJADIJYWdQIy/+d/GIZL0JzqkuZBFAiBBtcFk8vstc/t+KAdjB3eafA6AR6AmkC
xdE3GNBaCAmLYaLNvIZtJQ==
`protect END_PROTECTED
