`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0aAesNqC4WuRdPVr0GSy14FK0PGFmXWnHEvy8vUNM3Q5DqHx58175cWUMw+TlF6g
i8nizsLNgMBCPRCcSPkGxlFrdmB2U/JFo68XAg9lCHsFk7Fhe8vxGXrJa/10aPqW
4aqEMqAUm7jnmsAprb2cKy6wA8eUrWP3AqPwQRZsrvP9czgpRUwRjjMHQ4XFpr+x
reACmyhSOLaYnPnq5PV3s/75XEDb8zlfYxaMFZbcw+EKDL+LYtCi5M4Fuf82snCJ
C0aIjl0tZBZaQKDeJegE3IGcgFzo1RB5FgTOsr33yZmTMlR16c0emJLn6OUkS7Uc
ULIWTTLAOsRwkz6RsW7V1ZbsAtCiI9X06UZEGvgZV5X7I3h5S/m3ZOwLB1k/rlJ5
S5yHTGY+JTyqBfW+rhY1OjO1th9WR9QGO3zrIHBtVNSsinUAkZ25UCpNq8tpRxaK
+kQ6uY2PA7cylIwLe/uIG1yA9k9ifKZ9Fg8eQYpOKZ3SUBeFfdERVI1gGTqeqomO
7n11KNyDJr5rVe0QAtuGQrZwQ7tmDIRhHkCKmDLR5PKWIvGlRip6GGY0mBjRYmiM
sxoMR5b8hu05aw8RkEiLjWARsiuhGB1rU+Na+/OAwFi5npjOE+vhWgZdgfSz/ztM
DcXqVe4XNcYudyzm9LWxMi/ttxK7ikgXXBpMVCSQT3AUF9vYcu7KfpEkc4yyLgT+
1fqHZ+TWJ281T8L/7gKXzw==
`protect END_PROTECTED
