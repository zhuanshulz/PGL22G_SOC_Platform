`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
czRTpPh60WfjyPgLVgxGfxxQpjCjyhiQPEE8HuCwygBVzeN0kK+5kOFE5Q6jz4bv
xsW3vDbHwDmH3jd+rUvZpfarws+W5FBfCH8Bk0RsxZ0fc4swKUQ+Pr5YMIfOB+98
pI4wx56sAtiPiDhBkIPiKCN+LCc+hu/exzOKFHZD0WD5jIf9lRspwOcRCpLBvdBe
uBR+HVu/R4BlZpk0Keiv0jFne+kfE0co35BQNGwtRLFAVsPnQvkyH9IAhjmoh3BL
kjvC0MWFyF/Fm8Tb6+A/FEcjzWKkFSjSsCU7OCy66Lsz3v4RyA2d8+3N3XGBbeeW
0P9XOmf25q/XR/Fdf62XAw==
`protect END_PROTECTED
