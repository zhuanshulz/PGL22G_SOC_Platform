`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qeepO5DFo9zJ7iUW9SeLyxNPv4L0MysLRB6aXgSItHqlbZf9Xtagl8AQcbksJwZW
yWlaIcX+GGe2nFISZ2hDHvW6hDrjfgSGU6DxH7ZrOsv0LEM5PNRt2ZH2crO95chE
F4tU8Ac0sy/vVVSLflZwENYhCzA9FQE79xT0JuDhKGAjJO1nFhy5L3wCZsRXyqPI
zhO1dlv1tSwH7XgyJCeapM0q/NRif4kOl/h19YrLV7hZngABI2h3Q+uFmSHlKvKs
za1cieDzyNHF5Kg6Xz3T5Pj0kDIY1hxlNYKtEaX7YVoTlYBxmlvoh+QD/2HqkBvl
P2BaM+jBjJhnBaNTrhP/7mw8oElyXzBIyvi7Fe3CMHg1PRPw1utj8/FxuCHEFSy9
fil5ONzJyF/YYT2zwViN34i/CcqMzJ4W2DI8Q2GCpgsE27+ltZ86aX1XIrTA0sWD
VOdiUPPNin3oZpGGQkI039AHv1g8uUQ1GOUHiVWcHDcPPkO6gDFyT0rYrUnI8JuY
gSvp9ngaoB4rBDJNc8txbsbieOxwMRqolpTTkwTsy6CZkoIJUaQMA2Xf/WKgWxKK
VeNtDAkmOOTUoJVjQTipChDLk8jjhvTriMesgO8PRNlsgKTo6OIe0An71hA7+ZPw
vNE1MW2OR4ARE9eDQoJst9BVS8BL47YJfKcA9I+nJ+9mcyo7UIreYu0/1XXXliDF
jxgXTlpcO7PtvrA+3jVN/dE+wjRhNFtPwcNrzrEERrFERmrigXcTVqx5i86zOphB
H+X81LVG0PculrG+PHJ090EPT59FhLD37hUxuFZomAGt/7Qx3gjct+ORepEOwblh
ypa/BtHeDlaG8yBpCWkXdKcfyud5vtDzJtibpOt4yZctHAKdc6PK86Hkc7iS7gpQ
o53QXzljZ4iMxO+kYxymQHtSE3Vtyd7ytZVCgXmj8jOh4PzDCGqUCAB+EBm0ZhmJ
e4naBU4/5BMAfbmdeR8vPYayxsgTbofEYkXb7IiMHtC+8sb/QXME7f2zjaHRR2VY
H+dcuznNrr8TbnVJJqdMrDAXcT+C8jbQdqSi5WxairnRnQoccVQ0CQrJ0Yw/MQ1+
TIZ0lfJAV+nJDC3UwD9E1PHtTYY6lDuw8AjJrblGhL7x8uou0I39U/WyjujFoDg5
zt8TaEbVIoTZ+QqGYiRagbb1c/Jzy7V89Vv8iSB/EXzCf2ikGmwY6viSsVgJ0r/l
u/fgjJe/4qwuRjt0ZBy3rTCTnIWop6W5ohjayyOXzJohOqyRVcbbwVGPwN78OZNZ
WogoUpkYpmj9jJ3Y5Q6qK2IvQpHnRGLMkDBtzNY2PJvprBLlgJR0veRlru41j8lX
nyX9wmXEZ+Epi9eeykB0bRXPnP/S5Ap7/tqlKLfpOIXW8a5HKrx86Exhp5lmVs29
e7bol/EluY8mR98GVTVgWWsRy9Lf8K8HMTNTKSYsvrafjkZ0puta0U/zbDtNNg+O
Ohv/FXxY+ZOhOvZwJ//XFtxUcRTgs3MCa7LBSlCaTTAHGeeoJKjOHm+ZfNV51EW2
IWBh/cTeyb+VyzVUwY+y3iIS9vZdEaLJHDKCSIGPSTZubV9+05K9u2cXx2phpiBM
rD03OFKiIj1oHy7VbHujYctFGbIkU/UkPqCW2/97E/jDZ3ToypE+QOLy0U4lTZbP
c0W46j7OFjQG2LY2c3hW4O/arWUlF35w1IOBXpw5NXmD5eH0YAe1poSl23eJaMUA
l9uCNcFW3zvr4XV1LtmfKtEg6PINQm7ix+Odw61aAEPmbIK+O0uVL+C5btJteYK3
omiaNP40kcN2S0Ff05Sf9edtmyJDwI9kKcOkHoy96TRj3U8PTsVdtHMxAGbYOiGF
OApyLeEoA8yPUqm5utFNNEP3Reg4rGHb0eYYFlzhsYDKb8lEdlbScGXbF/Rv/nje
VVpWeGlLzaXB146FdgemJlMxcq0Bqruf+L/QP4k/ci7L2jdXgwt9CcpTVPAlkl6X
gAhfxFbeMNws+Z8VQ68Q7foVB1uCRM1OMa4ThpcLUgHDFd0iZP2RCRZRpPAAjLQh
mbxaTacGZDp99QN7JKIICe6+YXyu7VXDfgPOR2tSqDUoShHIszr7V4EeVTF8ylhd
Bi+OFfhpWmJxaybDMBoZxC2on6pyU+eBufEDqwXbOP1wXkDg3RfmBXpuaMd0vSVh
ZpnG9dDFOZ7oc8HI457e+MjbDxPPu+ozeg3eP0lSI1gK1ecRQIrVe59wldWuKcRn
pvhy/Hy6XJN7UTSIEbWj/IrdYmpJjexsQh7rOdKN0X70UJ1vRhUvBYCJNrt9IkYU
PIJf73yZ+2ZC6HwiLquWA3WyexKU6w/X1fUEKjO8XqD4Kt7SdKvBY+5NlJtUGsqs
X3+lKf57rvLTxDQ8vsTMEblV9AEWjCoRDkuLzD1KDo9gEbeAYJG1D5aEMHhoIXVA
wLXf3jMB0Rb+r3PODEwHtiIrKREBTSGOvqo+pkQ3ZTnvy2Wsu0d0IEh5nDBaSOU3
cHik8W+ETLNCLsURNK5lwiNPiNzc33Nv6GBYkmIu06uboZz/Ph5d18uH8c+vgtlX
Qg2w/TopQO3cu7kj6zjxMl/CX1rkqcH0cJ2mLAEcC7N9ewrc5FiXRy8AGQk2qhcA
cwu09C5O7Cuts03aG/+IHPUhtUozlDY8XGHQCFq4054dVfhEGmInbJc1AGTyZDzJ
Yl5sr/tgbY2TU+oEIToqN1a8Wdh4hgnE96zfFxh4fELf1Vy0eIVUo2Ws99vZg0nk
ev5LYaeEOHJ0qJTUsmg2qA7GHHoQJINIMBlBrT0ZXVcIVsI4cjVINg8FxcAENUnO
DqkxpFFBK5eux10CeTe81+YM4FR35NS3y5NKKPMXD5+5+DqCrr0at+cw91zpqKl+
sYo65Eqt1L6QO+UFlBPFnnQrmwtDXSfsevBt+YngGfGbywNTJiQRD5YOlbUY3W6g
M7RyLT8TP+FgEvLriilfaCuF5OLN4Q0afmuk3AiVhCrNjhJEh1Oj03V2yfWQxE2f
TyRt3npbReSBtKfELJ6IoMXxg+qe07ulilFUXVa4pnK49TESkaz8aas43CjdWfP0
aQ/jj/yzHUekBnnAhMnOKECTQcJOVlcBTHKQNo7FDkkzfDu3f0iIW+2iLGSrmqq1
twPgBuPJbnA45jXJ39PEFbRZmN76CXTVMSQMhAPlg6ph3ybeMsE/Eb78FgIuzHRt
BAscPdy1fyOdTacIHsxKw0PXMfDg3SZSu/0O9KFIV+KtxuMpFjaRTXM9wHFptFq3
ICNtDyp4oQO3Div2ysK+QyFoqPFuKYGZXtyQCFAeSs6+do5HA+XJ/s05IgGr/gQv
Q04DbvWiRRys+waWwlLNpPFMTfCkqN9CH02Kv3U3BNxHrt4S6AAcGVJcwP1QpOwi
r1TIYCJVEGK10pidjPWmd0sfDRj/01tG7ktlse+3yb60T46oAQZakzUpvD1hs1Tw
IqW5A1ruPsjI3AgPkSh7O/3QYAFEBaqN6BaCyVswMaL759OZbj6cEQyeNN4SV2iD
bBKXY7EIGv/IrHaX45dqTD9ydAXYRQzc0HmkYWATic9124aBQH/AWFEn8LfToexD
B9VjY0YExLXx2f4OUHRkfrQZEYg3V5fak6Mc/M4iV9mEwRQnYhEEKn/EvlLbuPhK
awJTFfB+aPqvnzlTAzJwgK8wu3eMUBTfx1/v6wy9JZ6EiKzEyTf36gaibZJHsGSb
+TKOelT2uOE8pM1UJxhR0pQnvwPbpRZZBilCLYmPXK1sofx8oaC5aDId9MJ9NN6H
N4NC+q6If292vCK0eEzvqeCNI8PneDDML7jUZ7nYA83IvUyt4pEvfyA7Nn3BmBlu
3OiJZ/ttzKE6HhnB3BZcQY4XLpDXNdAYVFwqC4j6NAfjJO+sdhXjoplhIfLfbj3b
7EFD0DxdScafoaNR4EfNO7Ii4gfr3t/lYht9mbVTsNOMDiCQ9dWh0WzGVyqYjsZQ
vDI9q8HjTFTTv7f23u7dNavDQYtquK8B8IsGn5VNboqvhGVJNcymyhyg1KY/Z+/T
K27NimKS9zwEw1C/2Op2gHb5g4/22mBfx75oI6M513lB9WY+aBJ/2Di3SpZZutMQ
CPL7GZBCbMIIAfyxQui0dw==
`protect END_PROTECTED
