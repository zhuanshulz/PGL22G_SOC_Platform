`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1of3oNaPVQSAWiDEdCzqjJr3L7Fhbvqp3cu7aIGBV/Mmho4LF1CUlLxFHgNogQ5l
bXJPx0EFRgpfZ4Bscl4u8yTqsECcjgjp+YYZ8eLB/L0SuvzZmKXmlXGW2k42oLBr
2wtijQQgtSkcp9QKFOagqTI6/B0yBWkEtP2ej8UHRfGl24sjL3vDn+jNaQMGeKOE
OnLHz6TttX+cpxHkT1c9zR9jrAUUsakc/iZ61nNFerlPvjxw6fhpP7woWU9wAR0I
WWgj7IdspXeDQt/77Nnxez+x5gKE25rXea7zxRzQ9SSmO8svsXMTqr+KHClnyNYR
OHnaUrpSAscePRl5podg9S9baCGWd8oaYJsYn3rPYLDVDQ3AszObUjjiZ7ArVaEn
bymK29anS58jimu1ii8gVQ==
`protect END_PROTECTED
