`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YH33nGuGAjr6hzeQYCi+i8rTvTL31oAlLjIL62lhCQJ1EBEeHSPREl1IoWnHEjua
pa8S2e+m8c9Ll6hyR5dFY4D26npcq4EL0NNG7x19iO+mF2ZQ+9pPhAnnD8opF3i9
co++l5Dm3SdoPJljRtQQykTU06BNVujMrY9WfG75OzQ7OgeKQBw1Exh7W0EqiLCd
GeBLB8DpSAOEiHb5OIfN9oDiacf5PtEuIilPATYo92WnHesrW3g1l3c4p8zOYlG3
xJoKIEG2Efhm81Fh0TMbOLuNomRrr+PhvmGBp1vHfBqX0eeDncGaa2kfxMNgP/2p
RSZhnp0kRThu3uxU/t+H9yXHxqy2zwyPaPXanCoFqkaOtpMUaySLgWj3dBofVZ1n
hDNyU58DMF7noPSimJnuJvYtg4ZxGFuXXh1FFVg9j23PsljISToU+5RBmbTPKxWq
1MEujrmuJ8CQ7Nnrye8b4i739/q8+PB8h4bh0yXoaPVJYXKuy6a5vf1uvqCGxpWb
JZAm/4LDvKiuEQX/z5+u+ECun4r5PxAEn4VLI34mR52E0t26irJea79jVXDftQrH
mzaDEHDUgulCYavr8eTr+Q3l3EgHMFGqMK1lZsLI9T88M/w82x9owysg6wv5oiw9
ey6ks+eguUir0PEOafXbJXQ8YxwnOWUEbVd19HiCpffVH8HKICRFGfNgHp3UAtyc
`protect END_PROTECTED
