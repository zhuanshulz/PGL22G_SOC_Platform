`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8MF3aWO/8m30l94SkObbsq2mGP7RxAQ3MXuj+Rbwhq/kEHEqt6WilPd1y17J0nqC
LvjzNwIYxU+SSv2RCkX35WoxsjDS71YokrEF/p8A0EM+csVIlVv7K8lFwGET49F/
Ec08cRMj9ipqj1K/yVaA0GOZCBwxTaXUYW5G3IKvq2ntffCVAhjI3S73jQb0vxMt
S0OEcOOesW47kS3yUzXZmKHEoGDBGp1SOlIflklhjhijT5DrablXNHtx7Wjb7O7X
dXLXxVRQNqJSGEj7fbuQsEBnhybAsDrkR3cIptO2x44XJ+omQdAPrIkXNg5gRoW4
PTOc4TKPpTkwJuvzyZvuFeQJfWAAnLo8iS6si9tl6CkMBpk5SsraosJWJd4NIcyW
Ld6PB5L5c7PuYTeUqvMhZi+ijobtXuw1OtUJ2AptGVSe4slilT0p5XMNZKon4Enj
j+qKB3pX0GvWOK3RDPnfdTlffD49Duiqzt1JxyFFsP4uC2D042UKU4SC1wJntKda
48SN7CUAVXGOKC9ooAtn/KUO9B9gYiHHENstflJO4yXIFIfHjmo76rSpp6k2fmtr
MtN7azem3xxzhiOGwOk7OSwUWv/vjdM85lfG35cnsUg7Q1WzlgWnuexmn8ji8Pos
gAjCYfbiOJ0YT7u1EMwK2Rtvq87ld6bT7THF7ieDs9susgEiT5/ifLLAOpLrgxgV
fkkAnRciwSGCHp8HAjDCotcEehqCkBlEihp9Ki1SKqtJyVzlc5mYU6E6D3mOdGuI
UAPkFc1/JY5KfGqImoNpHfU6mAYMIV5cHIwWsj5l1AZ2Mddv1z6zwTWyJ3pKs7H/
X/i0Nnj9CXJjcoOyS8EMNj+Kgv1spHPcx4aTnqogvNCbGeQiGVgJVRVOmKDtjdi6
F5TvMyYCHk/LGrXuOXtMUzO3I1vfkXvGbL40Yo0aUJ/h26Q4I3pH/j5z7oykBrXx
6Ac+L5NKQsxRvparNVa7CucX24XWBcdThmnjGyVO7v1SYgZng3TDB6Yj00qsyDgO
W3i0LrYcrPVMKZkT3Yxx2BcuwKgfnmuM6BpXtOYQOyaBwidd2oStXiWnym75T0to
BZoAnzgRV9cl0J78wg6kvPzNDSFSDz93nvz2Ivqy+WvI8+wJQikRBG3SUTmNkI7f
em0fsCOT9YsCzWL1/wVGcxrIfsqN3Z6H4Adjhhbl2hNcN7waq+ZK8+Wt9y/FVjjP
238KjaL8jlXf8mvgM+97jXDzmlEST1sVR3DnmTLuhfQQWnlGtpxiOr11WWmp/sDG
acdQz4DbaNndv91N+T3LvA58q6p3hU+kMpnS6W75YZmnOFq2aifFiGHdNt16beWu
d5zAurvTY6exlcxNBH0v/QYom6DjtFbAXYzxwi9IlrNKoM1nfxWSAbE+gqJ88NYC
kuxDOX5jqxFsHuDD59e4iJsFKueYQlxDfkOGxBggGyANkR1PmDNaLA52zIdbwxVA
PZOiOCW6I7PH1CpLUX+qjpgfk/bjcP8VmrciZEtTC2jEXvJmWB0XhAt5J1bM9kLb
/JGEF+WGu9EO66z/6nsfAJ5XMxHvtS8g2cynf7ZX47lRlRGYnboYHAJD7180LhG2
NlzLxhyqmLeZzoM2W/HXSXy0rN/pXWcfXstyjwUHjTOZjEMjVEdeg46KP4nutT93
wJe712kUt2MUsob0Ju4QdcaKFqcTX6HlyXErj4+UWff2k0CLzjtfF7+AiKcoDMFx
a1J/wlXYEap43UI/OU4bSsrdKhCkbFwtIDN0lYy9yCNmM6Zov457fRlaELezkb1x
GLREQo+b2mFARtkGTgeNSWgwxGUdgCqTLFAgl6oJsjzBNpRZjeJJTrksDlMBrL8J
jPbFtLx4rWPqiNVxzGrvj2u5ftIwkl4HXBnOmVm7waIu8Jf5O7T7rYNKu4XXyDj0
/Q+wnG4FbQp4ZtwZeI1T/u7LLVvlsyKeXzzNnj8VNtqP+LL4z+Q9HNmOT7QGLhEx
jdg09c9YeurCKuFhaQW2w6j5DOI/P55hBPrLx1eJjAcOnUB0oz3qOjuqO722akIF
VV6NIXu20Yy2lcKftD76T/RGs+umv/+jj6xoe+8xIu2ruc4R4DoNGm7E/4oEMOel
lrZdvRKp6OvTh03CAcYmJ7cM7Ya3e7RS4X9wt50mStwC90jO57KimpD1NPj56RPV
Nmz+Xt1ynFnxhFlZJ4cmfUMwEwypjr4Yw/wjS1MnsX1KUpN1sHndNq85KgR7pb5F
fUKFr0FLT2vlAsFRwritSIL8hvYo1lJo9doS5s2c6ona5Fx4AQA7tHCLYZ/mGd1h
JaTYV4nbRR69c80MDkWRcPgnhnfMfKk0fH84hDzHgYNyKzmWL2dygzSCnj4Xij26
quEa07BH0yLpfjwxMROPuchTKtWkv+p8qkzR4eSmWz/4yOZTpdycFQ0o3SC64P6m
qNRk4bW0RhMdLsw7XPhx8/kItZOBxjzlsProUGART4VNkVl/9TAkJ2Z3WRjkvdYv
prKQBzy3Jg0DVQ7thhyChAI1RINODWJe6O5dE4+xUBF4bL6hW1cXxnse/SMhtE2M
1WTN1LkNNK/ZSzvWfINZ/T4h48iz9FC4WivNFIhw3kuZnoR9Y6TN1cyjgcqp6DXM
IGQ7oznmYW42LKQliy5krW1SkPS+5NUsu50JrS12XocLf+isTIsM2Dzw/OveEd5t
Q9QWb8CXiSzuujaduIWrsZb8SUerAVP1x3W0Ji9/GZ9YiUM2bGagFZ8A741fUTJE
clZargDy1XWqwYW5HBxwL4KVVmBfOD6j2V3NPSXFYU/2GJ/lYlnHT3D9oBYxyszB
/ffCcNgADCucBMgpIWpjB186CaFADPjQg0gF6CDDv2/aeHiKtG6OoFoThhSW6Jwn
Mp0zLD0p5T4qpn5Xp2gTaJiXvlBdP5Nr5rlk/0AyyRPcvN1FKluOwnmerhSFbPXF
xqK+/PngUAYFI+FdBr7GgWxlQVdGUdPH+cRKeNuG6mqoJXiUvY8K/42J4y3TYrNx
Vy+cUlxKyVdZUIx5RZAl/qm7toBbMwgt2ya175BORNvOtQK5eawAWBdF7D6FnPZr
tDQAY3KlJgeE4S/KIWofxPmWUBZS0DXUiokMT60xph71l1PvO/k3UPBqFxJnemxU
TvoiUf/QaUrkMjM0iIjDEZnDwy82Ad/iJ4BxuR7WPgLiQuLucZeEofMq1cXvM6eS
P7bh3V57iTx3phmZfehvIs5/ZE7lNOuQHGCJpHYB7H2xfgTdgLVNNjmDlyM8Rab+
SISgY52CGQHMwYObQTAC7tyLwbO0N6C+lko+k/c5/iGVoRI/xRzcxj+Rnn+I0blX
nPFHGF/uOsAiN1K/3HdhI7KoDQ5rebM0METGmnpwOf1FK7mPUXZ9pe8owkMLMdta
nA7QoTAMX09JywM4HWjbyQ+jQgqtzwU6LbIhRo9DXM4=
`protect END_PROTECTED
