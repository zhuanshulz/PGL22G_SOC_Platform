`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NYwp2gtH6mg3S1buW/aHW6JuTDqBl83QPG0cI26HVxvwhSmQwzKKbbXHDhpFQ2mn
h9MZ8IQDeiTDX9/BoryhVT46UsLKfASYXa7yxJqizFtGINzNrPuBgkGs2zSkwhHm
KQAtOCItnFh2fK3Lnpm1xKPnxEa8FGKFTDGtPYVLfPoCR9fw1y3AXQdfFVgMt27g
R3bmXEBmGWKFSdWRtJ2iCJq7nW50cPDT8uanKzTtPkEr/l7jet1NWtGDYIV33Ek8
ksnU/1lLaWnA0t3JT4meJtS5ntoM9G0HDPionPwFTwPsBzRV/x8mCNrmhISn3Rcg
WRLFLM6/Ma5NMGXFxZ2jNnzb2wW7fh+Ex8dgPM4lzfYQl7UXs6gWPsfMql+Prp1u
ehXHF5ev9+3yP1/jS8eOZ6URD9l7FTaLcEN3ZjfZDQ6llCe3oQt28o+QNO6f6gfT
FuUYiX+P6jCUDsS1kszwll+2IW6B6Inhc/N2v+FIG2lVOibq13j5b7g3gteMder6
vckE3lfyy0VMcWXiee095mG5vsNWfBXdfEwZqtzlAnCQSu+7n8RnhabQl75Hw4Rl
cH5Krhwt8g9WZKKRfwRz8uEh6Yka3BRHCdxRIA7kDiJIxMSo2pkNms2A2riW4boX
LjXFzht3cM36m64CVGsn1Z+lHG0mEgKalY+mpKfpYiLLb6ST2+d937mO9cAntl7R
icJVgvmL7frK3yhQym3G8oHhQWFsxUcK8b7H+OoP6NVm0biuEWuJI7UE5uZc9Itd
FnDMn3FFVGn+D5MlnGJMdIODQBCfAhACGAXMwng6ZgmCKbdoQWziyg0QDEgDF/RQ
cj0A+yEWjbPS+oZm42Xp6v7o//VknSQs1R+tKTFwqic=
`protect END_PROTECTED
