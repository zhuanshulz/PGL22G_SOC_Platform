`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
beu3jSeQr9nSMrqdRnDKJ42nf1ZMGsNGXH6GAfYVrR6n18WeQIDYu0WclnOJAqcZ
yYfuFuRm5InoDiTfLHZKakh9o4nFquSlFRpVYj71QAxELEjelvH2zW26Chr9s5sF
BAG4eyOIPzgwQHkKLIYjzQB1xTS1o+PUJD3AXPrK56U9Kbl1eN/qYSs+9eFWXGrD
sVgsZA5uT3S5vCDfoui9VWLjXx5UI/h5sf8Df1IM8p1zzor6hRn3DWvDanJTyHmS
JVVk/4j6Xr/hUw2suUUltx5j16lkm+Xi2MtqDIlo2mQrL9B9tQctq88Rlr04mZ4v
eV7Gpq5cQd9wBCQiOVCMZwwXxAzK/rqAM+0b1l0yeRr8HtQinELYX2U1lk983bZb
aX2ACjJPuaQ465jRuEzGjs62od2JNtrS5k0ibef6DWtv7SZIXceg0b1JYNb/wopo
+ivTKgIemOVt04bbjHfZRyVFUAsi75RNmXFtAqnzeRQkqsZwCKvEjuJlC3Xir477
f1bVM0QSeLmPbQAcUQhkYkO2R4KxeQ95aEPAokdYbgDr2XdLP6yFLGCODDtsuREf
XqD+sKJ+6z3Drz0hR6ZvxqM+vtQcrls9Bf4gwS4/OAX/W2gO3ornpJPOV9MJNEtX
VzUpynWT3DRRB18I2dGZLMQfhf1ZH4mTS2CsqkphUr6QkjXRXfsYv51F09SWRgVz
wIYtWBOrUn1GtTMeegVRw73tnlwh8AOn9o6er7qlvFdMapl57DZFS1AaTTxVF61D
wIrB1cDZsceXffWxtkumAF1dn4ll8HtBHjBbScKZK6SIo6BP+hK8BH7t+3Q3uNa1
`protect END_PROTECTED
