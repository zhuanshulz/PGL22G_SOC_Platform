`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
55LnZDjwi7gEWZKia+4Lxm7n/Giu7UBSPqPfLnraGDZgg9hhfkGTrw7hsJ15iIzj
sV7AJ3VLNJKLaa3GdpdQSaOVUvvebKDs6amwfhR/rRqaxZSCKKYUVCbow73t58mO
2PKIEKOPU0c91jxgLlSfHjHMTuvf44tmldmn4qPYQd0iK66tqgAvOnESwxJbjPqu
PhKK1a1lh1exliNWaDjgjngO8sHGszTR/TN6zB0ftSkbvk+VR5yyreTIEKd6f08O
1PwapNYXzfDhNedkpy4upWy89kDVAhS3V4xC1tOCDGkCFG6M9c8d9Ozkg5qEfoVT
+pgcpF38wFVvOZDUuyuxdwpP5BYAXMDx2RLPchfo0tX9O0U3+cAmGnzssbVkX/M3
NN9FEAqsqbmlzedpQ4a3U8WgynirOj1Y+ekQnumQ0hc5quQsJgx1BGZU0puFDWmD
dFfVDcDjubic53m7DTSHAZMzfOxoQD3f1ZraRQ2lE+w2eCbF2SyhXFETBKfWuka8
rVQXncTedqw2U/MFPIiLlOWyExcNJwDVAV+kJ9XmZKStlJZ1ybMwGtlPxI6eCFO5
sie0a39gpI6knY/hLerQl/iKNj+7mVfpeerO83mLTBXI/4dCFN1HLazB6/oePN+p
+Tl7m1XXrdMtf7FsA91w8g==
`protect END_PROTECTED
