`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
THgQ8vFA9xWMyS3JTw20yfuMpoYujTSvxyslwCGnwPpnTBYaSjGmMM3Bb70KF2aa
1Wy/ikGTUcKqtGLG3J/Gf3cbcxqJ7xOOeOZUmty+ZwAJZ7caa1VefVXn83LkyPZB
LYkcAcKzoMRAjewy084qmyo52QaKo1mypTvHLnrpRPKWFHJ0nr3B5Xap/Y2805GW
+OL0y9CqAxAQrEwhv0AKT6334yj+91dAF/CVE+sTQu+CAT9OTjzVAEPVg1BOEH/8
Ol3N/p8pcY1NNkZHQI/GaeqVG7tBJ8RPR1aU6koCCfzKD2U4Go0sUs5vNOIhgNYG
6LL2rHq78TkXfHanA9Xf7eYZrjIo+B8rRz7b+v+giI8RO03W9CCE0Bz1gzlEPINj
6VJtDIzaeoly1/ZJRDus7TMyfemeljMnAubN5kQgezOWOal02PPo/Hr0p+sCozcP
PpaMnoXC+1HWUPHFsOyTTYgoschq5ByYyQqrdfmHDNL9y4YPQ8SgckRpwaPoYH8A
CHTadGmnSb97z6uEfAAceATjC0dDQXjf3vrd3ZURqti1/BOMDJeE8vgJ4mpq/9Sj
+hz5sTO27gVb2DljlDh26owUN/cnKDqd5Hqwn2dflOSqeE85ZIUQnjKYpKMBH45E
7HtMM3TBNjNG9nxLJKTdPRP7bMITZ7zlLwdTDOr5c7kUqgVhG48+9SevhDU/2jfP
ouBD314Z6OU5llWJzyn/8VkE6OX2bbM4hAPGUGPyA9jb4PzpP4U7crUrzJqaWQNP
id5I1ucqmBtnxxVYuy5pzqIvH3xvuFBm+Bwi1V8/YfiEyw65A1012BUvh4Q194Jo
rch1enHQMhmtYM8louuyNVSzxPnQ+Wmt7Y6cy754uDndtgaE6sXbiwDWDGYDJutf
4IQDh11h5NY3c1V1x1ftGKl4VVEu7PY/nThmD1ofRr5AjivS0cD9IR4Y/aX8HjnP
Df9aEQuMdl8ulqiuPqHzgq+Q+LfJkaZopqvmd2LAO8uYdbpQ5/L2QY0dDvCPN1G4
OP40IhI9KOoZz0fiNwf0S+I62EleLbJPNr312WP49K6AwUXszngMbcEZqEGtNIKc
N2vrp8eiXYjuY8Ba4IMQvonVj/q/8bbOcV1dlqazEBWbeyfqb9Xtq5iYZKea418v
bgehcY4uE+Hbh116aPqVWDNYD4TccSijoGAVz5iHEGZJ45U3UUyyuTYWgJ58PyAY
xRZRPfkwAU38f96jKn6B6dpwVYVZ9jEcUTONhnK8kMAtiHN1bx1q1FlA4pXwCgbO
05/1GPmmKEcLbRMwKTxqu6lobid+gBCVpt0br/DApOcI5BHbp8sgns0HcPg1reQg
otpsifxCtzla21kHhCo1rA+bmE96e1w/+2+3TwLPCB0gYajz/SJrtqkk0cvJNt/o
RiCtwWQ57WDJrdm7wGwkWC3COxMZHFonbNa/3efzfaHWJul89CiBBfSKRNzY7VGn
QJK2myFITnm2cOA3kH+nQMA0kGAcGsE4X0/L5xOWwe4mgPouGapFHciyZfuwXiOL
4MHAlKy95B1WaOiVz4Ex3LREBPjSTRKrxPV7axA53GtRSc2yFoLVtdxkM6Qn+6Oo
Tc2n6x2SJniodb3IZcYGAoJ5UPsPZXQoMSV34O+W2c/dJ7SU1rH8LJlaz8m+UdHm
2M29ymaAu6+DnrHPlY3BZ2qLo82jlIzLItmR+x2+lLQlP1IdVdJpSMXmJPuRfWYd
LintRgMzABapUVMGTDYxWwOgaWH32a6qntbEYwdbfiECKoV7gjdkAktHbm5Wx86U
d0kBoYCGP/O1htk0OWEpZMe8tVNW/KoXrShLXYq+I/KMeMFPyKFHPsoPT1vgFi/A
pL3ewSbvuWe4FF0VrYRHr1n9Tqtff9pP1da3d3h72dzGqVkCal5Gfkwndk1EHsJ4
/O1qf2Tl0iqR91LBfldLTliDygsIaaD/jNsRUEnADUrcgzqCmlw/N/KWs5fHULLY
epNj4rLVJefFjLp7D0NVMuilOzgWyPavAYQNZnaLQRcXjJyH65RkRkFqKGZwy8Sk
juyUS3w+nrSIig1F3MFM255wPBY83gdsYABqIJYAYPCjvcHI3UPnS6SJrnH6WJC6
D7fshHQgsVdHbStFl1tQDkUZSTQQ7674GLHw5YxBhAxUuFcLOoCtvt9Ng5rHIhlD
rhmMomonTlJpVNjgujS5CPB/Vqdg96Chp1aZxHuCJ/IPrUu4RRbMRlL7ZzCvRpPt
bHm29qjubbAWxJDpzKOUPS592DVXc759dcd9rY9B10RelDLOnMMtslDS3EaUkhVN
Ew8kyJvqd1ldKzRAyeJUUJKLbgFQoFBVW2LMdWDLUcTH3u3VjzzlGR1wBu7/5wvV
hCKj+os1fgg5EiB7SIWoA/XiidcikMg2OqFTFXXNjR9pMEZwLDdqlzh2bEqzI026
6aEhnYFTeZcpSedU9ztcNAquVK51BDz3ueYVdP5rxwHgNGgqqxe7kD20EZRRXk/j
pCPknbKmBG7/hNM94P5oaiyR/eSPIUxQqe4QacUPYRILroOMhgrt0iFvIaaTiaaU
9x5ozzbb73p5hqxl8Dc3OCQ96qkJdrVfs11524zILcSNUludq05hE4a6Rn6yzrQ8
jCh3yDsKFaKW4VWU08FNiK/jj/hWNQx0E+gYn+4BfcaI1MwpajQV2f9NGZyNr6Z3
tb9ADl+KjPDS0v/DIAUhfolFhXx8Yg9aO5r4/a4vBSsDjT5aoOMvTqYn1g2xpRwd
lD7MNYEwgaUA6DfKK62sBueVlqei7/F2Y1EoREGHraaLrYvXnTsRahH5vC6iK4PZ
VyjqZomUWkogYioBkaSpTCUlDeZJalYgf84VxVYY1WpwspUbVrc2g/Gh1zSoLF55
saXEZtYHkmBwZdOV/mzwUzr2MM+Rtz4DC7jqHn0zO4UkZkzUUYL4ofC1Yt2aKBf5
gTdUiRPG3erDBEIYmx2IuZjwfQIPP9x29h5N4XaDMeZUNzys2WzuDPqKsX3nCmYH
XcnCqEKe85PInNSluS98IbG+s2OiUgzOjP7vTxLcKntk0bbBm3kNloSU/19twBQS
84z3hjmVMdpiJfir3ytGbKeAVlJHw4ZaqB7kZV/e8RBbRSTeQ63yWY/zzdXesFq8
tkZBnyMOtmbTE01wIxxq7oDtYDGIhyhl40i+JUenLcxaKdxcbwk7Tk9uxDAvsPU0
qFkqkX1f5OY707dYsG+UJSiZd4FstZrlN9sSLp8dyMc5PYMKWulFuZ+sTKlyPAxR
wUZHciPp8vVMfGUZJmJ1PasCZCs8YbAhCvNwVdRvynmpP+oBCXpEYR1LVgoAeccL
ZJ1XdZM5rPnwyIl8/oWaI6yb3tTZBuqjNwfmwTwjHTuhFS45ErF3A1pPVsc+K4sz
4cceVRJ4K/imlT8x/BZf4uRS3Yz+k9RGDK9PTi47f/9xgtNYmGQnqZrBUOrxhvOb
vM45wzgQ1FrL3NKTSXovWG8J/HR1UIQcJpYGS3GIF7MJ/T2ICO53vZ3Y/iU0jJTr
U/pXW6uCzaT7RhX2Ovi2j1ybmmX9c3yAlhpO13B7UHpvgF02x9EE4EVTUOF6qISu
7rj2vAmcSCdnX9IgRf5FIyYFOz67gqtEPy6DuULYsX0okkn+owHTEuykw01JmABi
tuAiPDfxf5unKJwmvbmqgEUrFIDa5pQ3yKFvjuSvhNIUpqSP0K4izuMmofrmIhK8
xfldJYfgUtYRZodaAQmxguIFubDPHi3lDmFQXp/FjGJKEelKp/KPQRqgdf5ob3PA
nUmzWFtnwjclM5FKz/wdiuU9f5sXdP4o0eXc7CkIKRBuD8ieM2589RSvzpsDCtvo
RZKdtlMa/PpDVGjlOtWnPRX6Xc0ZEd4yllcRady/bmYNuNTEVvsUKXd2Aqof/Af3
lUP+PyammeCAcFGo9NSsIrJyD4Q29Z30R8cWsfa8HYN1mIj52f7gr8nKthD2w0sz
RENkAnYscW0YnOLCN+Y6rZaUrH5QCAGfr4OW0AicY576+JGIcXOC54QLruTjJngJ
ccYp6gFmzToMZtWTC+78rS0a0hyj1nntinl9lVzqfwHkpNeXhzYDU1Yv1KrkMRiN
p7G6SQM38he2PMbGGwmvGSIJ0Oi4Z6G5mFYcxeRTkde6pppQ69Bi//OMn4CGI20+
piX/y7ooeCwMUSTvZrAJ3voIN73XsIIlmNt/Iyzb/B/RqSp/0bpoBzFlKF+O935F
fUJFymVzqapPZQp2uE0F/qAvqhDErIQ/D7iVz1HErbxfvee7ymmgnTTC9NsRWZGA
nmy5Hs9qr6MSNAd2Vttn/g/hrCKLzfcl5N9bPuDJ2b8I0JHFIsL5ZOjC+YiG9X9r
ati+9rddr6X1XhhPGMCe91pIzG5HpM+7J83Vt8/GcF1BFso6TQh620ZLwLQhomPT
vkw/xv5qgeHlrIV/AdPqqg==
`protect END_PROTECTED
