`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+N5BbagBp7InA6UmT+/DpbCs3qxvx/UESV3AIQFe+BdEqedN4VKaa6uu36PkeCIh
yY6pBJgYuerldE3PghFzKUlftkzTOfI14jpjFubM8I3l6OSQfa8UCGl8kX1V23CL
ic70qmgmpeSF9JMLq0KOY/DGseSekLmJ9k2hfvmuPEiP2swOVQqrDl5AeACLrQIO
bUN3qZmqUTJKARa1UsGHMhDgh9HG0ML1CvUUSqCL5v5k253nqPqi6+KCq1avt58Y
swjvHaGKSGgdEgDhUvXbAnfuF1xO6njxyHUq5B5bDPxjGUPOSeOPM3S5EsU7LT0q
kFCTylhtb1DTf67EKvM68JZZ0HpR7Q1qu9uwcnhw/N4N40WBZITfGcH4kP4GYEl/
GeUE227Pma+oGG56AqCu7IstukJw/X5L5e7XhaqdVyYMrZRsL2xn9p+wYlwQ+mYK
z6t+rA4wBhCV+3aOrehghsTi+IZFdC0r+cQFQZyvI9EaLtvScKRUDcb0/ee8MyW5
n3Qvqe274ZKW2EDlbWWL/3E9yXIj1s4P18myzymo3MSuStpDJbw60ENAzH+ADDBH
SRvsMVOw7iWSLjrT3ALrRBTBxc7Q4tcGHXJjxPKVNOvrXrhwqccHBbjqbKWQjmZR
qKeNd0HxeobcLG6BChTJuJKNWU9/ku0RESH611bYyEs5roh2K/J3316V0hw2H37m
TM2bl2y0YrzWFOHWYVPXRBcEJdtkQkoudbcdPAPZlIM00MHXMGBeZNnN/SqtTJe9
Vznc69FS/d4eQO6Ainkm/60aGUri/rF/yaN1lA/YloWnVc4w3tGxspWZEUx4/hDZ
ZJdfuWIcQvjKsTGENkCbAylzrIqoEBkyqH/Bx9FeC0N3kbnJMKgu0zUHMhQ00C01
FUES2a+0XhSc9+rcCW0gx+ir2QNS1RWNHSdw478nxGTpqZ2mI75mD75njAE2jseg
FzHk0pUOFd5YXKN4UWjGiMw15jhGEWAh4pJ7p055EL+048zCv54gEZu/cFmSPvJc
bt8KeqtyqVbwaY+sLM/BQdcEGpCk8jTNheaS8UAgJI2HDS3w7I0V7RXHVitWCJEi
8FLkw9y7tnxkY9l89CS52pfDsaZ8xRf+3IEmGKDdC8n19IcuZmNogIj7ggZf9o2X
VQVKB0ashx+0/+Z4MHNUTxKGbXDAA5dTBHspwAhXqIRahwQwv7KPc7/lSC1klGcP
o8KihnoJMGrIBSK+1xSueA==
`protect END_PROTECTED
