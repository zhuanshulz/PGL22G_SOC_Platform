`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WvJ/9zDJEO1GXTMXbBmembkIY8K652rIjsZnpgV3Kd9SP+oUq8zqloLGTxqf4DK6
UtH6pWM4R83uvhfZcEfdtdgNi2ACJxqjBPGUIhivM7Q6XfiGv0yD/9fAVBdoEt3c
7oEvXwsYK7tKFB39NF9Q/wBm+jwikzgqhkn4jTK9Z2PTbo1/X7Y18rpNDJhnFKXY
IU4FgAIWXLAFqXDYXlwJbn2XOAM/MsS/Dgb/zKg2ex3VgkvZgbG50Og3oxjnCPw+
rPE8Qu+OcDaQtcB3O1NsakTEGc2IqlKBoaKYSeij3NiAyJ+tvrCmCPUb5C9s09YF
w6aLasWSkhJdHv8YUJ9rCmIB0xgMySBjCG3eI4kia7oO+LPEADPEfOPZ7rbqDEXj
JhCFQDDKSBWPavXf0gXeVcQBv1bc7FXVjSWI858K3YSuf82imhnPEs1oi3fpMo4k
OtbHKOZw2sEE+7idayKQLA==
`protect END_PROTECTED
