`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2l/EbGQFiVUbcOrvLndYh+hctVPACmcZ5Ie1YYO7TEmVHjcf+iZ7bk/uMs1nHNT4
4tvwSdG3imN8ZAJDs/+ZZnYdPfWPEjfYFvnvplqNyOIZAFFZpE4aOetI/VQV8pPz
1vQbvvJQVXVDdXLqeyYGatgESgeGyEzhEzy66O1yNPTDVS/U2oCf0EYXx6xH5+m2
mKn+B1wcqjGr1M7wvDkXv7YpG2aJy5lKyEqjIujS0gevAy+ao1ajdTvHYskvsW+1
gK8DDRr4LVX4tUtlOWUqGxBAiB53MVo2Ui30bWrqdZhtsSvSZ3UERk5kPVbM+Tfq
PE5kZweh6a896neP9u9xVnZWfUBZWV4BBxwTW3lW0JHOpdrW1NvTfu1Rru9uVH8b
8+gdQ2+qXduW9rtR6W0hrg==
`protect END_PROTECTED
