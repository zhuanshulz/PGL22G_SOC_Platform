`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bANeKvTdrmIIX0PwKDVOnlcPNr/f7mz2GSBkLfxFd4CsuHkriB5/NXpmkN35jToR
z9+X87YUBQptuO5/xlVfc5kTv60clWwfRH1XITnt2D+71KA+YM3vCQxwrKaM+Q5Z
oyBHwl71UC5MckdMwTzvbSW/9u7ZsSuVxqiu83WK6zY4aU424J2ciRes8ho4I92H
8ecfBd6jnDpkiRpQF2lO0erb8Y536CQBKJ7qNGjykNyoaTfmne8zqZBVEVkG0hWF
i0/DEOzgwzxESsRH5EVSSwqbObXI0FN6nahdbswmexY9DGKMkjXrNMevDa2DvKKJ
OS+4nvuxdofBPXtfrj0uZRMLUu0gJZwtGXIvEO5IqQXWWO7yhrIDcnzrzP4WDfKm
2tzTPKHYfABjqszceHIcD9G6a3pH1zq5iGoazqTRKrQ=
`protect END_PROTECTED
