`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yJlsBgnapJbjkTpHc+AMtKDQ8d/iaPJZGAvdJX/5Z3Ex29QUlaaXwks9of5I3nqp
y0rBN8pElb2oMw/VflterRGEfrNcdVnVRJRN8Njpczj0jLsmnVDB4ju+1R68mJAS
2VrhLwQF2a1h2mU6CI0MIUfSsaf09I1+293Ubz9mXX+LTpbETGfbRAV52N2NFnYv
1m3XFQB+EcFnSMDUIPFJtiP1xaWpHi+YIEVYES/BcRNz+B9T+bgnuzuHbMGwYG83
ewrQg1LHkupkvHWLh8PgsclYYaPJG200bWihbU3U4d5v6l05wkLlMeiZRNeQTPLn
fc86mw6VfZO5jjYMIv4N7YHlThpj0a7Rhj9FRKbFFix7ZHeKuFEWy70Y9ONa4iBv
EI5/b3xq3PYgl4SgTqzK1TjB0VuiaG+9qsh0igODsBYK/7LTXqEFxEXvkqXWyYZP
peCGXXNNN4FPHDdoIrCMYfHJvBdCqa2eqs/TKTMDEyjAcpO4xkpcN4gHyn++fpQ8
JSiCOaaIxG1eiiN7SgqpzbxGncNblP/XGIvmbLTVwpJPQV/kNeOXv/Erxzg+8xgD
aAuzMfCq708taQcJFjPzK7rELbtKMb+tKsO2Drn1Hs75W6G7cJftw04b5CqFkMUR
IX3HLnbEMDxLkQtvwStLUcV7DwjLYf6b4dHeb8CuEKQ=
`protect END_PROTECTED
