`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3odokvcpyY5xBkKF6O3dBR/9610Ww25EEzWQKiufQtCs40AO2JbdhUEBj3eqv2cH
uRUGPxJFyjnTURt4R/ZbCYLEutKZyf505TrJsnZq3jiLYJT2nS/JeOGDQjmgLSco
IqzNO3ughImAqVsTJEZMRlfFQqOuEqgeWvkWk033uZn/UqWFDxu80bE3Id09sktF
QSv0cUt/O8jcfN6j0Yfq6qS8MZRunIdW5OUTNumNzkObzlJST+fuhfJbBwRUbFyb
Nclnvy/LW6z3MV39qZ8AET0yXRrW5+z7/n5WyutLpuC4UPdegSmShoFMvj1LMTR6
pxYoVTPrt8FnuoycZoh1KhfBgcqCkRUwRaKXIZFAJ5Qoz+fErDifqx7Qa2BBMWhm
Sv3gNsrPYGQ02vGnaeco5TSSvV5/qDsJeTA3vf4O8V5hu3MgnUdsj+gG63X4KnTG
09j+qOb6Prt6n7C2/VGO2LCuPkgU4T428AbYWQ83fmryKUsqUtNb36T5uK16nsZ/
`protect END_PROTECTED
