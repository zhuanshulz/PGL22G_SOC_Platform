`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cOP6gU+56/eT9aubMvXPAk/vT5LcL0wnSej7jO4nclF4B/FwbE5s8ZmX3D0ymg4g
bsfypan5fXvG/SdkYW55jdRdORbogADG0sIgmIyTxruuS6iYM2xpmt1+IAp2Ji5c
VogKOzgFyVBeEPPOR+9tlhYgO/1g13AK6zegTEeaSLmP7X+iQcca0P6EH0JeYq34
RDcCoQE2k1wsH3uf+s4JwXcvI11zFE06of52Go8DWXIHOdc+bSfcDwzwRe+A8EVU
taEGxspPwkSpmA+WTY69JH1ZyBF47+RijaAK/ASHAuAVkTlaY9y0gUJqzSRxLm4E
Bfhlb628WtsZtmYjIXr2RC1hzdpIVWn8JkWKlSYOA1cIqLFyWbnC00tuiAhTgUDw
FsgKYHk7tD5NgMcBy2Y65PCl33MSTS7LjDh4S2s02EkWWMLN3W2RdxDWNrci6d30
137oQ3AYt7KMtAtWHVvzzx6c3AyDX3P5cqcPHePXK7/KFTOWmGRobkgXZaLupmTy
wYyXwXJdoIp3SOH61NPytwMtbxJ0Noonfre4qXPKMuvWxJfNcvZWpbwFjD5RDIYn
OT4m1u60+Ru92hUuL4Ck9wrUqQC3BFOzjdmSUKWDDo2+pH+HBTxvG7GlXQb//Kdo
BNbuMOQNxebnj5Lys1Uy+uuIl5qsS2zXxZQB7e1RBejdeGkR8mBuidRhhaq0vfLq
1qyRsNT+NsoOqO/nOrs+DrYb1NhIuYZSA9ykA2xGJWyOHSgqhYHnAXU12JLYBSIY
0bx3RTEJnzIzZQpNlsBcOeLl46uhFNi8m2840a3VzPDxKGHG0CuPXZO4DGg1Nwn6
1ZlNYCm2ksxSTjVhY5JOTsTt3DzHW/tuA0TZlWe9HxOTsg5IJTRDTj2kez+6/2Gv
ODUUmdAMoAuXIgbJk20QIITTwvmiRjs0c0H+sHbsPZH7TNyQrW2zSzg8ksBbfYcn
z/Jj9h1479IaWIOwfujYe9VfCramjqxo1jsR7204j7EtJIYScuS+262a3Wxj25ij
aq6rkUkxxhoq2LfMJZsOaQzw9ZY5NVqDV2/ScWWluMVl0KZ/W/KpH2ajS2rmVKjm
HhTg9gr2v269YxJbR4uJQ1pYP2XhdAOBz3dBFPrISVo6cmXmpXbGm1ge888qkPL2
G4xVsDtBJHRYZXIrERY492hNjFNvbmHuxrV4snzIf63JbeKDiaH/pQtUswMa/552
VFg2rkCVlW4QJ2CoOSmmd73jNydzroe4q8+grLQf1c/LR0FJbsQoOrwHj4KAtvmo
xJLA650pv3mzlItcV6XSzQBTbk3WuR1akosfDysTC0ekXt0l0moT5YLDxhd4xU6+
TJqksjyb0xGQmvIsKs8LMie1y38LIVCgwSmcZqleCJjsxpXsvRCe/QWKTGomhd4Q
oUGdoIjyeKdu+nEDxgC0iCERkQMNidJiteZWQeH877TEpDF0xoViLXynEGEvBkLb
d50Wl7Ip7ZS3Xiwvn+QcK1lnJ0eNkH1NZYN87gMOBMUBveihVce7/Sf7CfHSgeWO
V55g4gvzSGrVj6AlN/xTCaVOrIKnj6ChcJX93WNbNZVVxC5S0c4wxdabAW40kmDY
AA+Y/MwCBZWPwQutp4W/RvRorbPTLjbDYziIjFrQJkjFF27+Oi+JBdx07uJzIj9g
9yrob8luG5tVkwsZfBCIUdf/4wixYNY1ijmO/n5KNu6GL+U2kE3mtPGMp3F1V/m/
jZ2X8rJpY+uJyKXXyaYjtylF/1wE7mS+K8C04wGJLfUQy51iVtgcEhx1vrMf/Vdt
`protect END_PROTECTED
