`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SevOv1kE/N8BcvJkkKNSaFi4Tv7kGbpGzG+1iCgiQZJsHJC3IsfMDYDg00cZKHbp
PTyMgcDl2TrlpoPqLuV1kS+ylGbpHY2TnAUspfwAREB0O4ZJIVTdidoCslJil4sd
+h3q7NjEAQ4jsUnm8j8nTPUDay8/x4z4Iyniw9VUXLkc1GEqjSFupOvyZhtY3X/L
XgL3bABSpzmmja1jrA5DQaIWk53qDoHPxg3nXR7jBFymeKA8t2aeHnpUce/goCC6
Xe5P9lcBh+MeHqD8SPaxegzx4V4/JAxRFDa85kSjLtbSxX8lBhm7sYjXEJbC9CE1
gtqgNEABR3ui1+nDLhxTxjX+4itneWXp1NjGarC42NQ7+vQ2eI5sQLzkZKUHHBHR
IhbucodNNa3yjhd+NkcuRXDHF4EwZ8+vsoS9xbV33etcKZEEajAkRWcCNcy2vSUf
k+OjI3P27iCyZza5O7Vk85yC2nw6AHLD4wwXY1ISAq2Iwy9Vt9nzowaGqbvP73uW
Q6krk9y1wkYHGgYtLE/JJIKf9RQ6U6WaWZNaOhwkBdDwiDWSCZCeSvnha/ZcOngP
M6v3kyDB9x892txVBslZt0bQsNKaTnlK2M+6Qv6agVLPIyNYsIr8TwYC06MoN7+H
qcq8SFDkXUKet3X0spQ46vxUZNS54jbAIFwT/g8o+aQHdtO2tXwydh4/n3EcpPXK
kpPlDbZhuElVveRtDcTN+QPgBmkHvA6ipBKEEZUFb07bCHlU5fZWAVdCOkquko1H
5vAIkfqplZvCP9vZDSHXiwd5eKiqPyBtrLuvzWK/L3pnDKSFqQDgPmnactO8V4W2
sUF7SDu6G3SOStncivt9Bjc/xkeVKT59r6CMFhEDVfhgrhzXcfttbYeCdw2SHe/G
diCSCikGeXdbEloaQXxEVAfkKdpSQp2tgH9KpFBGjYrFFahKyDRb/O0pDDnajmeG
sC1R628CElI11cZ35KL1c+F6FLfWzGMEOc33Zu6TAPfOWw8dx8wn7QMFO8uUxAin
DVnXiuekwQkaUMuany+xRSUFfVF14tA+Ka3xb4xQ9a1Gokz2FE25+9+YSPFNXBxB
ZmmccEmu7tzJRunnVacgu6yH2uX+IrKhGHYy+aMF0MX1XR57u2fIb/CDbvOKF0jl
x83KGcv0PxL7UTCPdNK+YzIIidk7/wW7XOniIp2pqxbj42Vgau1t6NfnEsFIplU+
R0Q1GWaJxfyfO5N79g96AJC+TSoNvvkdSCkif7IMM3Tq9k3W8XodgRnzSFDJ16BQ
hSz+Fy8f3dtSVbzX2MlikJac8AkXKyV0KSm4sPpo8SJCMdkkdUGLVsxteTTdGJVM
L8hmsBpt1fStxQiY5yuDmw/MeEAGVgB1r4c4S+Lrav+CB8JoQpc4lhvP7SQgaEkT
S1JfqKoxFX74zuBfL7iU/p8f0JYHDeJNw+1N/MKBIsrkpUil8QY+wTuYoka74a/g
I2e7OHsG0nbngZMxBcePJCN8bzy6TDcOh5Bu4Q2l9CX111dQAHeiOnUpLV04dumU
5IbvTAXQ18a1eX1RkH9QsQ21lYdTohDGOSiSbOQCsaYURoTVAzQSjMozqkaCxqnE
iBIEAKyuR2QaSwbxZ7IDDnwGxAbMehp3JfJZzENregryBF+DJ4SjdRmaH1KM8Td5
VB/3GvV1cWqKW7bO9ofcC94FBc06k+uDGkTPfgcpwZarTtxKmE9e+aqgEV8eTnlE
pIbX7q++DNMkXSGzKCcSRaFqjPmLe6I6O7h9Rx6iMz8O7rBpXp+qaO5wocKybey1
M/ChubSud/NDa8z37zfh8NGf8S/bl/lccRO6SYMEIxasjFEmt2mlb6UAYK4/Lblu
DTpIDnHzCtVyDIUP2cyYTwPTO9asd+AYo1r9PcLprlpgezczEVZ6TbqP5mD5qRVe
FMCZH5Pr2dHEwkbnY1hzZNYgEBs71GkrrcyRx0XXHPk=
`protect END_PROTECTED
