`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DAge5nROHysrs63z+k1v/AhTOtzwKUKUjBo3/EMMs/+Gwbzot707MaXJ6PqQ7xod
HTTHsOcKm5QgOUowuOgIGrH+tW0PLldJRqyYsC5AOwmbrWY5MZJO++cGjIpRiA4r
bfuWS/oi7sj0xtElljEGqIyAffLNVZmNdm3SN4l3qWR4fWYslNS0A/3DY7ihqKxO
O+xwcit2zveyAM3j3sOg3X0Hpizctzvgu6E8V8P29LXg4/OCSL3L9xjDhAl2D10H
0rxT40KPupA9Qk85WnYSLmWWOshkBVD85/5WfJXWomYyGPsdirdkowW0fieuPXHU
Ba4EI2RT1UqCNVLU6KAN8jNY/xwuhB6iCbpM9Pbh57cGUP2A0Xk0s0BHTXnIZbbP
owMBV2S1VnoBjgTWF0B0Hbj9APQjkDPxSXTLdvM/y8zz3JBs4HLxREPjQioZfX1f
GDpfev0gR005UU4Y7dlq87HGX0/RehSfItHJGuYfRHyBRcj9IV6V221CzW9rk+Dw
rU//G9Q2sBPTieH5rnDa4kAWf4s5N77NgTinKhWjyOVVZh934OV+0hbdrJZe+cOR
tgJVO3SqHv2tLf0f8XC0phdoj+5iN7N5jjG4IuJWvL5a3HxYDiFeTRA4EkYZ4RVB
qSzvUwn3YKByn8Kp/CnvaPl+fRBIBY1U1UVD8uU7oFqJS6tztpJt3xO6fp4k3Qih
IqN5B3tOxYzew8vy7usW1CRtW8DgkrCUHn85NuMXdG8=
`protect END_PROTECTED
