`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
03I2O5fMnIGA4AvXgdjLo5IqDwFLoLCNLmmfL1xKv+JjBahaQSm/LQgqGB/m6Fsg
cOQ2+vM8/cHyGY9DHZM3GFtTpZC+im36J9/0xpsDMQgFiwid5q0rKm/Xyh2gzB9Z
JPo/BvENAYOrW86oukpB5rcY3UyuB43YkG3jCX59JC5KnTJHYneM5xxTfbK0eD4p
nKIvKuhZwTC2LAM9FpsyD3a7mnCUqnoWVbazgT2L/oSi1SgVJTfnS0dEYSYaBFmC
HsXf6dhOOEIW50KuMvmX1ju5VUEpC4FClheBt89sTRnAh1R/hcz2v2u782pNCDsF
Zu9TiQ7UELWEdZ08kzw027ASxEIOuHfFT4kTnxjT1mHPOvxBo9GrAJllAYC3PLXw
JDbwVafL4bZhvubDxiOOpwEQeHWlkYQm1lU2pxkVW+C+zdtbF2TL0hf66mfcruUa
k1KhwE0QJXnI22GNaeByXvfcfDsUkU95dJWfUMVmEY10zfhV+FAFEc7p5JZRHZ/9
T0+IPxY7qc2/bZc5ZVhT9LI9wkM1XuTYwZkX/C6YH7hF0vDGPIaQMxCv46fiMHHQ
wxu/94SbrNuUa7KG4XGx/HziHIPPS/4L18eOoYGNFTFH8QLMJo3gwZVxMtIQoAlS
gXjh8Llg3AfLToCb1xkm1US6lIFvfLoaLECk49fMT2gl0JWOCQg7sBUIgoV3FWJY
D4blVIfkMCA2yqz/3vx45sURgN34s8RY03MHMYTtrsSEXz22jz60A1hSy5qlgHZd
O5TD035lCfQbIcKE26d8/8nO0GxY5T8Nm9IK/Rd8i97lfb+3PvZhMojrj0ULahQp
eVbmpWm2sE5jBlaYNeKbWbDSPUS5CzILQYFTX8cnTxSrO91eLA5Xa0X1Dbk1Utm4
HhuF7pCTaQwFIoyASzAfuUnQ3fURcDepfb/5cihQXpdkQKWjPOpvMJGYkpZlJ/OW
lhbJtMIMgsDBq2lpMv/frCtJaoqvL3f0kR9V2z5VXZEqcdknt377yhFZVVFwWU5X
afKocuLtHyqKYZdOlx710PIFRLmq6PGCXc+Wh42i8IEM7aYeWYkAdbaRopsEJlhk
WcrdZriTQ8uSLiCm7gqymRlNDMkXQ7Qf5b3KGEl8vAXe7+k2lm/znyaLjegaVxB4
mD8+Xz+cmh13lY4NeCmFL2WaPQ8wSlpM4WaFvJkZk1E0g23hEoTMGOeloKCK1ceq
fIAfet2Ej0A48FRCnC+JaClEh1blcJZ1JNrjU4PZYAbaqkvf0Q59FYvg/G4AgyL2
Lbi8fpd4KT9VDPEMpmNNNdTzrr8Po1B9q3kObu83UoWPFcPKzzw3cnG97hWjC0zd
cJyE9uqSgTo+0ABh5g/5hg1EciGIAslGxJATVq9cvDuoT2AkIn2tDZ3RpEiPA6GR
RY+lPLtJkD+veHlgXAar5ctQ5TV8TRTvLBkhgmoqHTFsBYSCDkW/bjSSYZXUJcGo
3EVJjXNc64tqxRCQcnjzHpWySXrNb4oQ6Ivi8ldZejqZbjDPa0I/bxlK/SWecUhB
0o9A3uSheJIS/gSqtDjtZqyjXSsPwGBbwypz7/QcIzjg6VHyQtSNuy8NjydVDJc8
hiuR3nxfkedd/hicqw/TiKRXTCXNX1bI7r96DhYHysPYKVQb0BT9IB+XawwiG9hO
L+jgquRgJCwM8tLC25708vq1uAUdHkQj5WuqPaxKGZJxSM5NwjAqJ1+a/iPf3ul/
5oQwOSVxEqDRBErHJXek+JJn6KPIJXOmdnPAQAqRID5YsF9QU4f2mcOCfX98ZeDA
Y9voB68cs6eQWr0fPYGPtnQTV6sTaqyV8BXHXE+WQoUb30QLJJ4mqrhhAolALzF1
u/Y1gf2XScaI3odm1PaqWAXRO+5uOpP909fpHKp6Gizrrw4pSD9BlRSKL047osUm
lSMdP1KVe5swtjT5rlhNzyA1Zf9BbeNsWe93E+UaJ13wjUjAE7odes2uBkxGoXVB
h4oW5sj0BGN9UsIpaAUhg/j0rwqYqlFduXl0kNLEWFzBaINOu8h5o/pgpVZtrCE/
uWvZt4LsRPLuh/E9kZdtdas198TyX4+r7PtN2DAY/ePdlS61PwB09UgM05lUghX/
ydxpC2iM0cIew+xgCytCxvUk9JvY2Jrpad6UvxuhgJGFTFgvqRRXHtOhKA2w8a5h
MTu+jQqyVyrk6yxmVDeiAU7y78j/94tfAVcHhzFDR/CfzaD2c7GN05HyODmQj5gR
aT3TMz/SWeE5ste4xQCnTBfzxu1bALwmiwvQzojkAzLHrkfZDQZg90HqX6xt+UD3
e266kWoYMZ1sODvvq2+lJg8eaoM9tF09eDAoYPtcaOuakSLcI8fkt2D95euTzc92
ODy/EJ2qHph5eoFf69yX+vbVj7tWyuexRLNmTh7tYUxjQX+ddZUWfR854BhI/Opj
N2tp2mKiZ/RmWUa4EPlPo4GSygaKSCWBB7HftStB407RtoWEtxy/ZERomy1HBo+8
fDi6T4cczwUbpYoe0e9SaXTFpPqfZxlEfQj4CgDYb1B1DnpcC1IfRNfvkR3BzLKO
+sEnuRuYN61iiTMDWbhxVVMuaRvD9tEqMrr1qr/ghTPCKwaHamcjnHicdKD5fKKl
DORUhA22QTfgU000y84ez0/IAQiDNT7VWDDe/eXIPpNNSysq0SbomYNyus2GDII4
4P9QFTCqlXQ3sjmKaRdJyAJHCADKnUqsx/Y0DETgSyvsLD5CK5JqKfqd8ZgqkXJu
n6sA85KXfBO8AXLaIpUeYA==
`protect END_PROTECTED
