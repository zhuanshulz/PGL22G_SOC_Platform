`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0BENHBqIVvYmoYav6ds6NODcQYJ7hBVBToBhNI2j+6DJRZCHTMlYPDsWSKmWE83Q
dPtr0i+p/ZxfneRv0sSq58lZLCCXE7rAR+Ngm6S31Lpgk877BPWH0Dvadw+ar/Hy
zzQU09xC5AUIa0Z/zDTUSR5icKaJlY9iyvOLL4SLzrpoB9OTksD9pJbLUBQ+j0P3
M/55JGBjxNBQzsGHn23tmkc/kFcyDl6E4cHsPm2p71X+UxgPPfX2xU7Pwpd7yNxO
J9RI8H0rn0f6k2uQhjCczBfFAMJ40x1RhhfuO2v9kPVGEBtM4S8yVF1GOuO+dIVJ
cedclDXyd8bxOKDC9VQ8UB2eG6zuJgzodg0vB2I0pZFdYiSJZ06ejk7H2CucYHIQ
LM+rAI+KvF+7mW2QECsWVP3IuB1SuZJluJmmyDETaHdtlN6b1A3pm2utMWcKxNKg
IaS2vPPl5II/xTNAsJvYA4QJIQLdcrroxnCvCmzsarzSij0WuKIvcr/5NRDNcfzC
yXHKvF5MQcpGeNf9hBewYt1AfIJRm3RyOkm3ptfU/csKYM61mKavxRnPlpnyDG65
DyKQeQiViBqkvHVwrbNy8Nw1uaPUatRt1k7vJX1/LttrpnGDfmM84ODpKMNGtPas
5YzldddlFmLrhoQEoUDFjdEl/QsBRyudnU7bAwpnjmarvvQV8BipFiYhmoMzSs8O
KMK+MdwDUzwkCCCdQoCIc4mmhuFlPf9dqBXofd2ADq/LLWozfWPeeL+cNLPw1CiT
GVM6khs5mx5oNzhmV/nEVCnmI2L/kXWaNSSQABje9/LUcuc0L6Y0Wvcc5wFZP6EY
wXU5NLXBoMuAm5NnE33FmbcYiF9dhuv9TRujmh4iRwK2B9ufzzCi6ZbO3gTTfzY4
z6qvdr04rV7np+MMiQi9Lie+ISVTObDIGEWrIb4aKo7u+brTAGJW8GGyHlQ5bUMJ
WuHOuqdKCwvLUOZF8+shOReMM3YbpEcOshwhJomez034Y7GYUjOieyxQO1tVgtGj
I4scbj56e7sbD5WdcfLlDscJuVt9Ls25JE60B+el2Ig=
`protect END_PROTECTED
