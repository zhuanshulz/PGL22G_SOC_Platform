`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v0HV3eDYITzMvVlh8Fpg0MUwd6jsq974GAS3wpjr9o4jKBhjJ0OShOo2TyYdCL8g
ScAjVEM8dOxAPc2RNA4QqWRSX/VRr9kaUYxzpVLzetR+imXhq6TagzVcobWQp0uB
avdlvg8aNloKHFaCykVZ+m5Qi1FCbK+TxN4IfWmCDBHQvpi2KShuPwPllzVYZfRk
+zKvlv0YKBWmckheFSavXmBPT1bGFEzvzuQsMEe4m6Gmh3iXTtt1O4zzB61nxwPO
Es8Rynt3xo+SFYsnt8OqWCqqer9Vm9KeuZoIHo4f9BiWWSs4NjlEBbOl6ZlaODfj
vItezQIpGsSlBM92EnS5U24ILXjV8r1nzpHnt7vCIXifmmP2vjFmEUKSqcZTEqlq
Krpo6nXbpaVQ2VL6bTE34g==
`protect END_PROTECTED
