`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ny5ywX0Hfh9EiHcIJO6zDkZqZ+Bk6qsrQM1hTdPFLC7wGEpUR+t5n/kWi5IEr752
/XPJf2ekjFTY6nGJayBREwctJkiIoEJ9bAkHbTejR0a7rnORfJwG+8nZ/VDr2dOq
42JMkcuu7ccYaP9pmu09WBxBB26i3mhIeoedSQU7s0nXv4S1g0DDn8v7CO6l3ruU
KkQTl06DBM/sin8v1IHpod3lDO5P2Trblppeqxkceb5So8gkEyG34D4sNEHUdPyr
RUWFGsacaWJa1gvQPdDUg7ckSzmcYArk0yDtIFtt9pGm9jXDrSwcD7rtm4A8zL+j
Cn9JSJ3EEaEn+wpTxGu4Lxl1yAhovqJJs7d6gsFVkt5mT7l0Abw8h9WneBQsB/Ly
P6yjF2loMrQlqFc65TXnCg223mHjmdT4kzQNMcDT10SAoIh4w9D/S4TcHA4VEp4M
Gk/kphlOeS/gYD3vF4MmzE9wNKd8rJRg9KK/dvPdsDnPG8cyQdtx4OdfffsoRdEY
LUnXGY6rh78g78tP7GI+N5+TWo5Yy3WX8yv2uJSdQ869nAhHilkuj3s5LZlJTvDL
0y+3F/spNZvkFyxhW7Zkdw==
`protect END_PROTECTED
