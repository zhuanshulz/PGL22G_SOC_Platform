`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7Cb0bHVWekDBiz+jttkjEuyqwSPO1eOpBd5OzmuXVXO+pmGGcY0RTB/oYWYmVVqG
rSXcOPxRywzfaWo+EFP7fnVdEE6Rt2tniD34ilQl7W8jPVwnZAC5LuabuaDEc70V
FekXWE83eZP70b3geKaZ4YygW4eYK5IRJvLqkl1S0xd0lz6osR9Fv8JHDmvkvQKc
0fvAArcUo9if/O+3YUNKqMO16QS5t6sOVgt3bwm/rUADW2bKtSCku8jb0PCoNEbO
vf7GxgIL88HtfCf1ckURXlQnEgVEUEqRc7Ci+XMpVFPg5xMM9KbM9d1syKP6AClj
O7C+NMedfltG+OZUOJf7YRemJ70RyhylLI3DjYapxKVeN1Kxhgyvy59B2ebm+HZX
vTMHAK1hMmpQ5fe2DXjti7I3OQDvFzShth9ILZM65u63oD9mOj0liQhrPVe/jWBz
6aI1LBcNgIBlPz3tgKYhP7bnxlLExdq8B8UXOK8u6sy/sXfGUrzIWsLOJQiISKUw
1ICdFS81Cngce1lwAb3NFoCoANMZ6HLZvHqUFSlj1kB+fYQtEn+eGsB0FgHr8glB
FWrMsA8j7YfT+YDAqhegCzcB21UD1L4zm7G+XhwAvqsL/w7extp9wPh8i9981gRT
5qKHUXfNiZVi2xkxjDK/8KNpjTe3xcChX5myuLXIm3WsIpKpwaU+jQqjHdgBu3ne
JkTuI30lCpgjhYI+rnebQ6iLUTRbSzHiCjCBUKIX5zUHx0hfRVARyll4vAe87HHR
zUMcbYv/eD4BTp+3Bp/ngOqxDTiL8AMvEjW6Uwg5TafwHAPjeJU+IZaY6D9wUSf2
QpdJDmTlwRA7PY/adgnaykt/Al4ysxmcNuadLNfbKci6L3QmT7kkv7mtpJLUjegx
rs3eaykeR1x/EFLwYzzFioTnKWmBTDXNCe2V6aR8d3MoG8dxp0gjL8YLjTnHnrIK
MKRIRX7O4dNLJqV0mkgT0AH6Ht3Wcn3ALtbnFGAAdzy7TAuE3+Gx+hJfXrhij5yV
FqIKEJgvkClN4OmLpIohjCyRWxTkHNuZ7g9nMfL5eofWh7CaUDq/8wAqJeUsM51S
IFcSDFToeU8kMXyLiuzBtXt1J8JRBvPhCOwLQr4Tmm/V7p6s6t2MX+MTdDKWT2s7
SaMbSJ0A6SbSiXCSjZR7OzMe4L9OLR7neZS6+Iyim+UuEg6R8b268z363VOswGox
0B0MzN1vocjaE530WL1G0NAdP2op4GeDvwSVd8DWHNi7FTXnnhXho+/6639migKh
xyL5EqP2vZujzcj0qEhpMEYxgm6olOVJb6VEFBqKyiAW0NCHJDpBdqTs3vTiSYEe
geSsbYI6cD0PQgHtWwNGc/pQvNZ3Ptu064puJ5bVGm2q9z16+BWwQBUK7bW5++SJ
tvRY44ZEVF8mKwwipdPZ7XUqsP7N3XJgxIIGwiEqqm0CcwrEd6hQK43hZlBAnM2o
UgE4SZQcp72ZMnIGgaHRuUU/m7jVHM12Mij0jg/P9Ft+7C+E5mRPzR7DEoNOO4nr
3npeY0wsAOrL5PYxcAsD8gCZWL5he7R1BzrnnCvGbPf0Na8xyoiSfg1tqRHDYo6Q
oq67EbJiXos8IccIg7kRqmoYLHXnfzJ+OygV/Uc/S6A1STZJJzy3NL1yjVIoAdLB
vHtxyrYnKd9uOegMw5cKWewXSZHZ2QvWb2eO7efqwRANQC0LagMr8Kla69xC84Nl
dlwFHd3nSMSJRX7zTV5kgBXhuk8B6LeOCwbEB5itCvf51zMyeGeEbWAiQFkckSTy
JTD4VcDwlkQfu14feuMvezMfQxFNsU386Zjm6EgndSReMJpmjKRMeNx3kQ5I7W7S
sP+dWQKE/fCC2NBMsrwIA2E/T7uSl33hvB1Ex4YQ9OOFVpHqnO2MKKmU/57lQQSp
ktoLOgpt+A7j4dQR4DWxv11L1JwzdE9/znC9ukDqsZdeggVM86PYgVMNvkIh3J8L
RBNhrlCsLRmp58gYwlJOfTIil7QIkkfH21qXSa4NvNa70guJyU7AvmGo+H3UsJve
NK8YqUFjZuF6DpClLnFqoAhv6Ar0dmETc8fd0naRS0emXUzIfFvFeAxVuKMIcS1p
3WJQwliP8Pc3FjYDuXAR/23JFinr26t/HkLRdcIcTf0TQHTUOl+eUcFYFppkJN0N
dGqR4T0570ANC4xP0OJiwfFvJWFrw/bVyoOr/pyqwICwTUab/lnTwm+25a0jSZkC
cpzWfJ9zXTlKeGiG2vRgMhELDzJYL3UQuIr4rLvMvpIGZ0udJ2cpWxeU1X58puXS
z1VxUCJeAyVqO9yWC+fzmTn9juuKfiyW+i5Usz4VokPa0SQMK3GVGp2lYZVCkUhK
upX05S3wZsS06c4/eS/O6QgzrqyNi3Nh0M4DHI0rOfAz7usyecdIYqtAxclOy3f+
Lr8XDtM5zDlQAaS8KmHwBS/8J6IVuG+o5X9aUBoqmQPgGWGSP4osJ5diFD1aaFjG
Iju2/LtWmkagms5h0MOUrN0aE0yzUSpAkE2wlBAEzf4h6eIx2cwOlF5h+Tc+Dhaw
A64El1VB/dC40TvYy3vNzThwYWU3qIXmHLER6WyNcaf1ygbtN7etB1bS+WFN+Wh0
`protect END_PROTECTED
