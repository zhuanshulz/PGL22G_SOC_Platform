`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j/k8mkO/3Qh4Fdp4DjEauKISHnqvYccdlAk4Ex5tqvX0MH0WwMb3CPZ28Qq4zllt
l25RjoaoeyRUnTbRBeoH3IE7qjRUNMYmQJoaRsfMXu87TALxO6CMGksYHWWeCVg9
SZvxKD2ot8gfiyWLja0QBCBxmtuPn3CL6Ts4aTlQSt1uAXJaWmEsHOnlj80zClP6
3hAnt530/1/kmn69+5iXkz70IBBD9mBLUZU99jH57kVONOnDyJkfL3kyuiQcvXgj
6ERxKXZtg07J7h3jtw65eL5EozWNZ0NzMOhxXchs5WLKSFiP7e16sQcpW6SoH3DY
75Qn4QoCDuRy5GxFS76yGxWEdNC644Daw4+wCQpcK5M6HGkTR/ls9cr6x2b3YmtK
V0GEDJimXdOMoHz/JrZlQmHkjMQO0wvbkBQAqZEiFfkTYCvsreq81ZCLOgRFq//s
zwSNuPCYLz2GU/v/8da+K+/z8vWAUaviXXuKG9+AFGyFRRpsP3vpG9FGzCB9GJdW
otuLLVm1FKKnDodZLXTNj+PptUULiyfwsouFh4EVFubXUhVLr9tNeFOEHeiyoi8H
GeJzqULTbuXER3DGEXscDT66Wt6pGD1UDf90klWp+qZSMmfI01xzJ9KChCWO4PpR
b8TLc0sW1O+f1nx2r087vhV6nLU4J0I8wHpPwq4NEN+1mHCDk1xuhiab6jALYzkO
xE+TPNb/PAYDVKobEWj5N+X1xeIhiK4VrkWsnNXYy3NAEbNoC663Nmiz3HlRBL77
7p2TEeh76jJCgbUl/SEi07ekr7fXAxSmT3lP36HcdfpsF+of43wfn7T8HbIUgWdx
/OQZmE3h6l5QnrGBL11hPanlxQrZmaCZCMwK3SDv7CCL+go0Gs1hZ7beT6EaEJ9l
UKanb9TxS5mOBSWatWnstEo/lbJ//AiMZEV/Qjv+Kr8bwHV4xDATHxqFnnFszigy
LgDRILKdvIOkMKH1lPx4fA==
`protect END_PROTECTED
