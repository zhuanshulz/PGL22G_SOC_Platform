`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sUpCBivb0GfzyungrE4CG9zTsZzhg7/ym/SWzn1voQFuN4To+gT15IQLPWguU77Y
iIPiTywqdkzosHxTVLwc0oiUVz2fVko2jEqsTkyCEB4kxEAzzrmaCeP1WTozfrJ6
OjJDz04TUpMkLyNLzQSTHLetgIRcyDvPeIuOHwpq1W0IJDZBteLszDzWyDlVOi2u
BuBJoNe+oSaF6s8Y7d/S4389cEFEdatRZS9BIUKb705+cz8EgsDOngVtWZQPzkhr
iyio5WJ2Fj0b+zTyEX4LnownZOPARrX12Cuoxg+YEk3+lJTrAcH5C3kmELjxIY08
juvNlERXVtewQEhETTnqKJ0eLWwb2Ytr31bfLLWmgg0v4OmJHMUYdIiAVG9JClfn
8g4Ds1Ld1n76AqRzDcf5Y7d0JuShNCLCY+xknWab22bUqT2Kn4K5fTTPsNRjdWNK
vF9BYzi0EE+rdq9Dr1wwBDOtF3vql8NmCSO5lOJbUj/tq69P6PFfCNqrBhczTaj/
78twJVJQLiUYalP9+9Ay2FyedDgXz0Q6UHJ+kjsZ4CoDqpiI0usbuvDNBk7WWtLW
n1qHKlXpXB8a3xh9cjALtPvL8kWYZiebxLxxYhO6FjzU+i/g+A7BYi75061XcVCs
OiAS3MuEcTyY/EwfB3wkGPHnwY+G1vBPJUH/pVBWP75+Zwx7dN7HGt9aBmAnMrTv
YjQviOoK4i1+GeZWSfjI8t6ByTC5skrX5Cd2exG9mNfzQVWb4xgxxcY6CEWxPl3x
NwbtPy6r2YQ+OkXDIsVMAp7R8A6gFtScchsktCtkl8hirKTBD8CS+B+8gpfpWSa/
TiA3axEtSPH/VKUTpqCbY5dG4LdRpTXsuBvUfEeeC97YqxV+T0qrcKlDLej5w1nA
37igIfv/3cF5wOldf3eytT9dj0hE31ga3Fpd4XZtsF7iFx9AUlHeJPoac0vwJIoE
Iwc6agi7aYdxmLrXzAr7jZ1mLWHZNIzq2mPVuHO8Sd2AFDwSQgoehaYmrBmMSW1M
Dmz9+I0BMQnaWcqd2By9F3dmdJIX8nPAGy3ufi3Vu0HT31APw2Gk8rG17PD8AQ/I
r99cAGzGJCeCuNsFZZGB9CYubnnhXN2befQ8mrOYih13stQPrY+FWXab342Hh1/A
2uF74ZScIg18/NXYYbSXJu2O1BuVgK3GbnMf0sxCKkqfw3wZ2l+PccK8zSjuYiUl
vH7t+TWu8CVPk6pkU2t+H2FxyKNHn65qaFC0Gd8kEHS5e6KYnq8QCAZqc95Bxa8i
SgF+H/mQ8LV4PBRzce42M1hF8BsjCwsyb8bw/BojtN28VD7Gvkw7X2XzsHywbEAO
wgZxy5+nYtMzhwYjcKTvFqJZlL3NIPJJw19b6OdvaaUHxgtLPn2VOaQr8OfSveLW
vNYe1i0vUucX03JbU12nPRMSHRZLLFNQ341LLXJMPDLIQTvZYtiH54ZfG81YGsLV
7TTWQh4dwKmMhVzZtoNcajtCZMimojTxI244WYPXMrvsMWjt8H0InWI+rKKDI9vM
FTJBX+gXBobp5hZXnuvjLZy4CdlDMXQXetDexVc1Z9WPg5jsqq4NoZwV5uHpybgR
9YW9jUxAzbYW+jfsJbKKe7p6qgJo/9dAXSYQ/yq4a/6GJaN6s5s9BZ3Slna+pzX1
Qgrj9bK/FFlRFQUqYZR7MKJ2NOC09ORRQYTw4LdXXdrH8kX3+BTzloLx5rwTQBWV
s0N67+yUmBF462gLzs8B304wIBkhF/LEzbYZJeiCS2e7iauFBFXb+aSSWqzVuz7k
2Y4RhjfFdH283P/lJwNfV5cqRwVQ3JatOtwE0aMVnab4n0Jw7xelWO7deViSThJM
nXrtN0QzHQ0q62ZIfJDgn8MEr9mfj0Sgx5uIa9RcaJZTRe04K+m2TMfofFccMf4Y
8QH+7xgrw+j4RFfAqeX6lrR6WnqkcxbyRHElvJGA2Em57CwmlMB0x9tsP1Tj+H4g
CoU5yRRSMjjzIuAXlCwEL83FadjCv1pNRVwc+ci0auVsyldOA1oRWhQdwDkj2UvB
OlxKa4/hge2tNsDVwPZMBehTL+Cl0KFDa0UBCLBQ9xFEW2J3aw0jW37TLGEJkKzp
CvcEy9z9B4K9rn+PO+po1CYvCe6S2ymcsXjyucJ1iXjS36t+1ZxI0FqbcF5z0e+F
T1YNlU4bgcwDPdbxUlOjf83KJVOhB5NjH7bvCHZs4ByuJhFcAUtzMxB+0rcLGw+j
vHOqs5rBG1BOrQDKSRyvKZAZVB3NfjRw/Bc4MIU+NO/y0ScHyXWucjW5XELA6hGP
G8kzp9+oVClHqJn8qS1qLSkY84c1chNRUamEj1WWOZruBfgAhmZzGy0P6jVQEY+H
TX9WUqyzUrtpTFOibdcSd8vkOQnITo/EmDC7UUN9Q3Vh4WvRiULyPM+73vAk/wWq
IGjmFMJ3qC16MTQp1IvCdfoThFisb6kPSEhw33a6HZBFn7qPBgXRfsww+XN/+S8q
IBBP/MxLj9sKAUMj74uw1EjDawB/VDpkiUwYevkeut9Wl6nwQOpTGGdEKU6ev+ad
+6WUAhgLu8NGeNH6tO5bwbi4t5kvpJOdTQdWxctAp6P+YnZczlwaWVzC07uICXvE
zLndFR+b6EZI3F+lwZAMRIIsBthZsX/JXjondPq7ca8JQ+Hlfi3rqpKIT5A5GVV7
eBcn0sr6gFAlejrF1E05YMQektrt1uE5BEZlWSSxASjOVPMCQYcyW69DJI63MIvw
5PP2OG+BOHwACyRU9Lzp23Ijf83umzmm0B2u1nj7mUm44XxjJrtJNMU6fDinLBuo
qQt3buXaM/v1DLG7ffJ2LG5Hrs2ZdxwdD0uFBxTJfV9yQW+JwxrDnZMqZ81QoHIT
Tb1gUoJeTCuvgkj/iJQg3bO5C08nq5orH36ADDLTl1zCI1dAOEBlC2SPci2XIWOf
grzpXA91vkg+q9rjbgkPijz0Z8WmE3bGhLxkA2Z5+B0dFMalyU3vSNe3uxUGRdy0
x+jjFGwGbukOncthK3Xq5guuFPritAl1cnd2V0XHdeVIU+Mx9mSlALiSXE2e4YBx
feGEbYkWzUe8o4kHO6qTc4nLY5lf1WRDqHcR5vU2rATK8I4oVhLa4zQv/zgY0JXe
vPwKquchbmRXoIp8/NwlZlQR2Qh5dJr2CjFi9XojTBenCLDcYyESLz3n5qCGuIQA
dgfGpufouoE3VwnKuNccPXs9Wp4a4g/i5oIowVr8ps8KdUS5ZN1xiYphREtUriuO
vn5wlopW73sgwSat8j4KIzIBt5SlnMpsAHK/cGBWmzCIYKYajrXcISHZez35SHXB
NVoiLC6t4FBMqgcPtsQwyW69WE/cpGCrl8F+gUD3nzEV/5SODL0Lc+qxhylQg+ZM
Be1/ZJ4buijB9GHAOSLkD++3QwZMH4DpJqxq2flZmGgWdsId/hD9q1bZoVKgqTcI
RxYRjkLGfAW3FFHjEA0jPXVAJztUVMOqFXsaM9giv+Eg2JXoZyW3Ylm+A8a1/Tm2
xyXbertBeKekSFaXdUtFAXJ0pNmMF20yp9lxEsFi6I5RctW6gYea975Y5SNCkl5d
WKDei4sT6Me/MvUdOg0cvn0MlytQiLNGNsSFrJdd8sxxHBsCMJe31BVdYWXw/Dbe
GWohHg7kvZ1EQlaohs83JtJWLofjHC1io8ED+5hg4L4Qm6fSmhpbyNrd8mItzLhv
QIF7/iRyGc33ld04bY1A//ql3ZFvDsEOLhyY14an07/JKDXbT0MfMTWJUI+Fe1P9
bk8236mRPtZQad2oP2TKuilwXVdnhKsjQjdSYqyi09NNP6B+TrrKnya+tUrH+iAU
852enJfildLIBtM9j2qyyvqlUl8RBZ2KmvaJIiKY/Ir+qT2Dgwwok42tPPkkEKF9
9s1UU0DF4ddztJIy7gTDJ234fFwWhj/WW/b4jKzVCXl8xclFd672b6ZhFQJCUakV
bT7HlmUttoLoEKSF4z97AH2limsDPc+59mQBQzEhn33Rm2iyEQWJs2AOAT16uYbR
0IxX7jOLdOZRvI/wdMh7uWUnWAmoD+JGoMheW145u9fpCrr+UbDvcOfAvH58w2Lp
zZvuA8Ff6ByKzntF/UQA+ZuXSR/GIdl6iL2NsX9RsEPU5IDv91BCqwmYjBYBYD74
qHC2PMsQQ/d4J43brS/x6Gab8tV1jR5sUrjBm5fs8281PxAnSAn+RSdwpa51iG7V
b8frZCldftmTMd1xHIAetfXmZMunuT5afgxtI1uN/iDKzbRM94RTxJn7Zss6efB2
JiSlyZ/w5eUNWG2V4QDAjDgSUPPzDjTpx7WZy+L8tm4N5c0PyjsD8FwRB2NgRSCY
kMxOQhgPVbgZAdB9Y9aqDBaEHR9bc8vuF0iquZQfARd2TxQexHce0AlO+xX8cdA8
VJiDipo1I1ObcvOVm0FQHRIYbkE7Kc/Wr1InWDdH17MWTKceS62Nm20uDUuQDM0h
ET4aKp4Wwl2C4R79xkp54//33JoJ1EPtXZ0VumQsqpB1tbnWR7z9ssv4bO2bsuLm
oOLhyWtF5vu2OJbUIxeAX1dL4pCqzgU3i0JsjN6cWyMsyry+R9FPxVHKWubq6El0
coedP4LymR2WuVCd+4iWc8+YVpwWqfX/+SMlI7/jTHhj9KuTv2iiApYw8VdRI8wv
9DzTSZvwIqqtoohhezuEI2RLdwzhHb0nyC7dzTq1ODotaGEAi2HNtrjZi0QXcZX7
fdWEDpNTiu1kvKMkBV4hMkU9GDBHIfvPc9L+ofIMcvRrxaBGQwWB+bBeCwGSGADh
LKr3aRiqKM3v1smm2aQ0T7FcR/CbQKkRVjJp6DDeSBk91oNz0NOUmeJSLaRE2jy2
72snINecvyPuvcZ6gWpesEQi2Fy3tJnvd+AHj7CSylnJXzomAxiTT9ngkpxEcP8d
Om9C7cIdJokuVxllCLqgtZC0nNYNDAg6GCNeBDgAwAr3qnvzx3KI+LoPhEkhZNH6
0lXaf5m35eIUjbAO/GwSJ4o/6M6o9E1dqJ7ZdH0n1qsyLsG1ddhaM+pdvQF6PyG0
X/aLG4tJg3mK6I5Q0oaNCjb/0qrM2BMQf+AeWQ51Pp14ZnX2/sa2uRFkNjQD4+VS
+vWwsU6WX4ZWDusJ6FCLSSt5En+Hzv7fgb+I1LRdRgg3d9p46UJ0e17JmImuh7df
4ECWj+bcZsVb9WgCFu3aQn7f9EGdvTr3SvyPuMZzu+DTNAS/Tr+AjcADq/LVXNyG
/ZUHpRA9U6Psm4e90A6QZynMZ3pC2n+Q5dORbL3TVbpsAECeFlv7DvGZIhkQOXS4
pjR+QMpz2nwLKWam/hLo4ZE8uIWWqBbM1Xwn1Ec2QAB6v55X3vLl+YDgjt0s1upq
cOZVTmO7q77Xg5QIqgH+hPQaCbPN2rHDfPAi6zbw8ElJvkjfJLCPq7XtrRbZ9WG2
pMxG0YaTE+d5qL6CElhsuumLPSAkH1TpQXm3bQ9WGVi9NfHK6Jg/4juK6z/8bqD4
shGFJFl3wIEXxq5S4WuPElKt4QssKEhYBLWWN2s6cOV5kKtOg66A+lGR9oIvAbJt
MLH3YiDfGeqfJrT48qkyZxXnsdFf/2RwmBUdlj9IPQN3tItVnc9i1fnn1VgwiEqr
jRUQS7ExZeI+XZiA1GTaRPUOhxPOd+wqyK5DnFPSdtIDHPYS9a9iv3+05BMGstID
yisU2mLW7sNh8y5JDsTVA2ER0I6SKAZaSVk0Z86H5x24mBuBfznkv+wBRgD/L5DA
Ia0Iaxse+ve1VDC4HRaeXVUe0NxW3hBrqoR3meBvauVbMU8EvUL9gnjfHAPB86ha
W/knPYuPvqYXwpBhsgyJtRo4cr/lPI8kNG1u1VYbFMPsIIU0315Xc7Bd6CwINl2y
Z7x1Q8v4yA9y6oacchS23ydUcXArAtvhBitvryIDePnbWB+5m4/Q8OhQ3yUBOvmu
7eAxZb1+mGAeqtbGika0vR3V99AyLambzOTPpQCqQ0rDuyT1ahPbSkQQ8ETviW9Y
gtyGciRdNQQk1OilqQJLD2pNHf+iFlkvyOdrH68qBCyn3Z0OqpTehJvc0XPoS8Z4
yxCPBx3jjZLDf+99yxL1Ri/3nY3cTH3H4Lg8fwp6YOMfUXc3MrOP79m26C5IkCvS
CIIoSSCeEE6zvMPfL+291M0rMFtKOrqx+6ALAK9B1L6dnfQSoal0rr+lPuAwC+Nt
/3T5RcI9fnlzSa+XizUFhS1aOjFvnW9EuaU9698is1T3jw0M7yjj4WkMGCUX+bES
M8MGTvGPbBdcRJMXt7umNRRhTBjpgwEnEUhVdY06JcSg+fUf6jv2MJNiTH+mqWhP
yiEor8iRNeLPBzhWtKdo4WY+BsWm6kYaqdM7gtYbClrYItCcb264yM3PVVLdi3u8
Ndb6ydTrpwvNK7DpAOgIiGS6LOtKLflcTvcnfFQVb0AExR8/I8TaCQMvz3VYuTG+
IO8iaAvs1851l3R6NruwpaO56Pt5y09VgWtN7h+IJq4XN47Xobf9y2ee+dUxNNN9
B/d2o/mV12NhZBOJGWVXcoQdNhkA3ECfa/zcvE0u8vkHk6aFyKZxUweILqKfNsUM
YikCl8+KXltReJ+G9afuu6VazSJB+lAsKwf58VSFHV70uHcaSyYBTz/eG8OeKmEp
ob2lZfQEmYQFFAKyXl/g5pW53T5GvN+cheMfeYyjRXK1nnFVg0BCund62B4CvFRj
0RSa5mnEN9FkOAfkPkoWnGgw+YkiwSl3Mb9vNGJ04pXPb7LowVKVpxQ0qMJ6VzJp
vDpT4WTNGV8YXNWkvLpRdTZ/WztKif8mSnm9IuEK2TkOTBfPALDP2a0w0DVcDP5k
HZGa7MxfxOZcoIL9FDpT5giHrobHDs8Suo5AxkTN4um+m4uNrDK4jL10jXjpgobR
E1A/x6sEAWdYTBzE44QpoZUu6uzyda3yZU36Ql9N/i67KQIAr5xI173BbjNGqT65
u1QL9OlNU6xbXEZ+OVRtSPGxrkye4JwhRob7RJeSDgUbmY6zdpj0z2PmDIxgFd43
gOltami33tBkJiXNfLha+75GTGfHN8+1EM9Uz3ntUjqiIyzjXV/K5GRHPjgRbSFB
hsujH52aB60HsgUizYAqzFhAsQYXUOe9nATWOIbwWXHYhboudN+Y0vAWqHJFTIJx
KDJJCEC3ZEIF/6BK40pZKcFSffp56uAUCKyuGZps3KxC9kRk7Pr9HoLTwGix8q7w
KxllqCmVvRUbEnTpXzjZvdyen7g+rMh9ADUMpsat6dbpeMIbtDv6WBAZRrIFn+vC
vbaqhzlCFOfpK9qKthZE6Vhkot5uJ/7glBfsk6MxfTFyM9C4P4u5zlrN3Ar35wn8
UO15HrtFlFKny80L4DlMbl0v+d3UYq2hWPCH0CCrF/QPuPmy4y9r040xc3Sg6jni
rRl9VbuYiRmPwPlvDmWZee4wlxiij3l3uq9umEuHmJTB5fWLVWKBPZjCUfgKhmNe
PhsyN3Iei5x7qbjD8RpkJ3Zaigd5FYyHeIywhi956Iyomws5CfVR2jYvMXwbAqFs
ezSQaaapezEbY6fx9CJdqdVWIIOYlMcHkUuJlaEbhRRnJxZsSRk9WHM38IyTTMWc
hOu0CoqP2KqchBSdSmTwzg==
`protect END_PROTECTED
