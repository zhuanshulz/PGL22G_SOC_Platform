`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9bZg8SQVSXyBKBdkfOv+soErFlU7Uh66pPu3jLJMWLj1e1LtNgeW30JWfJMXF7XZ
u3YLWOAt3BGp9avtwUd0OgN0ilpfenyaZY/WG4O5RkY6DQOZ+iEOA3NMgu9X5+nu
4+8r4mYMfkQtc2DahoX/9o7oo1R01bdexlx02tyZ+8Hw48xO7xWb6dbX7NLxNOl4
XCaMPgU9+tBv4DOZUd47zb6srgNKxOCCArbwrcFp2L8EOQHfcQFHUyHXQzSqKGjB
Yow8M8epoeg4gak8Ngw2HYk70h+3kZGbLY7gnVo1BJ3Tja1O+6/qY6YnyqY+nIAY
`protect END_PROTECTED
