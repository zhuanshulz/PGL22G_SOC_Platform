`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bz6UaxfC7uo2FkV5vA2sBh8BJiL5wht6gv3dQZmDrl1A1rqolradHL9phakSkBhb
ZJnXaerGzfIVtpTQYzSgxSxawk/QawqsXTC3uQM4fZAYtbQuEVkD6FkIqMsOiWgL
wAYPY3qrAYTMJRqLmjT69Qd0LJalv2Cx7rybyvJp/sR0SK3n1wCV4+ks0rcWsy0P
BLEP7JicxlXj2JNOkwuMDXppkqvzck5k9M7OuDdhcyxGePRhjMy/ETMXMkUQkz37
pyba1ImjfhsJWM87Ghzj6gC44CZB/tTy7GthOUCK/cIN8Y+ckdYfVNSljvBOiEQC
HZk8sk4EnFZ+6etQlUu757d99THrNak+ubViITjK/XqFha+BHLACyGq0zv+QsyCX
u32aNGxFXYpJHh0qtQ1tbXIq8pZs6LER/WzCN+kqb/uzGkpw8Vl4J5ycN+AieRTG
dEkbwzFwFPqq/BYchLxrg5/eEog1A1hqcxGhyzHC1/Gzp/Ujyq5qGYAARTZQLEpG
xZR+D5hrQ3uhHRRN5jZAjRvVlhT4qbYY2ySOKhNdvUvRU+OZ5Mu2Bm+/bif5rLCC
IFNlkIQVKeJbI5l95FMjoCFSWxMWNa8+e50XtRXNCP29yOTgai31ArtsT067nNUx
Ps8IOgDbuEFPVYTwoaedhlQUbOu6v/0r4c9/bt3aQSPrMdi25Y9ayPdxNFJarhg8
t3dULQbRUT7wuP3cpGO5rQiYD43tEj0o8mhvcPMExTtdilRUGpSeFtspO3G3LLal
OjP8jzkRuEUr+7Cc0/IM0yuNy5AlUoGkJKGqQTM0JP9ZBJsMFbSrLpBY1a3JHw4f
2kTrGBQinjl+jtc/S8ZYkcM7IgKBNJ2wQ32vKbL9m6CtmNHDAN8LgqDGwbj80deB
MCND7LuSaXR/dG8Mb8j4LyEtVtqVs2Wc7wI6fYE08Gd2WRSpOQUJK2Glah0AKn65
yNQOdpDzq/Iei2zR0DeDxmLfhwi93Y8taV/tUiz51bDGL0+o8qaw+zZTI3RwNB3j
xw5DogT5KdhAUpElvvDJwEmBB20WZy1pn4qdNjlSDyFAwbJcGj8cyVQwqG+6A9ll
7t79F49V4lq87JXCw6+aVp8Lfre7D/8/JeEuK18OnXnXiqKbvtHbdzZZR+SmdhQ2
8OG0wwf+bihIm2cTkUuTgP3sQsHAFmiZfa5oIIFj7qo7rYEXE5V5+zHi4bCE81sa
SKS3SHvhYOE3XViBwKVBrZcq7jG0mDdnmL/3kJlMqB/0vuvory84Ek3CR2msB/wz
DTeSfEZhk6dx8Q3Lm9ixsuW9KwLzjKLPOs7O5Ss0JJIVamTg5kCtZRXUS+OEkZnR
H9ttWSORL+OIa3NHJ73mbOdQyrCyDB3w4ynWMlM4Mk89lByxLaYXnqlbeEaXjHIz
wZaM1ic8rJbNk2rg3X6HpMrnv55m5dspbRkTnw5US8jLYvD+1M1IVHY/8NwgI7bb
rhmFABr/lQoigG1RkuA7upHDS+FCDwt1izFNNJJTC8fgsqDzXEW7BN4KkVIvOH9G
irLbIsHGf3EUQuzzviqrgnvkc+cLDdr3W79vUsI2FHAPLN6KkxsGto4I9dbbI1+1
MwE73UcrbS1ZBq5ALZP7vjOsKYP//lFn7u47m0AwJ59ilCRY2FrgFA9AFVlMfxfJ
Gt5E7pI8uo9ZN+d9OqfjDncTCtDLsVSKYLyVP+v2F3UThy0lyzgSAnb1PA9g5GCc
8CyoeEvflvzMIJPwpKSl/+g9oHWxfeteexK5KZ1V+/QK+MoqM//TxbHZfpPMB2fQ
fhn+9OxyH2FY2+KxMPLBRUlPyJADuqi2B+R6bUmA3QJ2j7WGml3qPE+AO1aP35Jy
iRUVRJHxC9++Q48ToCSjDffSGhc/PI3LGtaz0WmIlMWRj9erVircYMDQrVE2yL6g
Yd+rt7oeIhwGT8bm5k3Jc5IwOmIOnFjA75+OSPiKMfLSzM2Fb9E2BxY0mKDC6rYR
JQNNNeR0JkMF2eL8XeqOXd4XwUZRHSD9yMhwz+ZomQVsr0P5pjMPiYowbac6lclO
93uI6C2eHP61ciiTMwuicICIbmnBBxt+YKMyN/gsIS6YlNpUzvPGbvRVmPuiJAeQ
fSwZeLQEVPXnGc4RJ/jCtdrUjP18yIRE82pJrjdkhc0Nza6kZLynjFyb7Ebr+YIN
oo1CsBIkAugydSRrLvMXMeK3dRmTYu20hxHUk4+oZ3Y5u6xX5WFpywv4exjnucYe
ZhukEwrW1MeXqP01ebJwm4ifGKCtnLpCP5LWPWiN171Z6la0d/aiEO071BDmvXeY
RgSHWaB3iQh3VuibALdVdvkocDVZp30clS2QFd4dodcXpPt7Ph5hgyctalO6OVbQ
1lPAkdsSgoES9Eb4jGbI1rbN2jcnZkV7YXJVA/9KySFnavH1uG8tdOwRU3U3Fn83
dYs5hG4bShj1K3d9jOcSVVsLck1g3XmBulk/makZKSKqNQQgBPzUFBvtvAjzNjpF
plYfkQTDgRDx6sN1NgO7iTRH2XlwX4xIIdzi4Zr+E2YqlkNbpoweBBLNRdB7KuUt
KzAMwbXsrp+ntgiTz676dK8jxmfV380EcxF/sO8dXPFqOAK5ix8AW30wQhBK53LH
2xnfi5q1x/hqotniUN6Z/BZjz2BNYk3nUENAT4szGL/W0bmJWosMJGggp4wbN87T
kdiFExH86W8IsNiXDMHViYjJlN7hDdbvuHdmdsgUZQBWwcLT/8mut1LP9jGrArzm
Prhj26bm5unwvamMg+UU4jvRcGj12Q8FwvWAZxisKDTrHgsoHBnjyScj3odpWAKN
6lGOIErMZu8sflLxJIu2Tik+QiALxu7D2kOrek8+1PziZnK4KJliXsz77GLsetaI
KX+Vzs3S/mtU7kJKKkXxTUJGFJzV9FHEE0zOX2c2lrbfD7mpRl7+GHDb8Sj4ucut
YPHlwTbyJW/sAD0UaiQifDMpTn180Aofq0z4nmuWwJm+puwwk2i22UorY1cl/7rp
wcJnjxIYnApuyML9Kjelvq0zoV1xYdlGJKz/aN3Jc4Hqgk4CQgjKvHacfwUHWu+Q
pnBp85mubf4+f+ryYAiH7/bMYLCJ/6FEtxXQ5PVq1VACd1wiZ1SBzd2vcSF9q2UE
pcDisUxGNn8DefSnlbb3u51yZPlKEH6QYj5zAN9WIl37AL63WNIS6PZEMucH2nfa
gdpqmcrPLs3eAJnn/6pdQj8ocbNQyID/6Xd1HfnW5kW86kqpsW2jYt95S7ZLNCHr
DJpD7Du3PirMQFCRXAtQ4IJhY0VVacmYlkn8toxntplT25wEUeH/TFsSGfSqBQYY
GptdBe+VllBfgRN2wH1Uru256fxaV5OJNayycC+IBw/KmQNGqHGsuw3g2NbdbiBm
gdElPO0xUdpT0JWGPV4P1UzgmHABaP4R4nCBrK42QijOj3YpfbqwZk7/IVJ2hta6
3Aef2KFF5NTsFe7fykhwqNBL9+lclMnKan/x/I9Gh5veAaAhKsMlLeHXYxOzHbdM
9RewRWGdMuWuhtByHL6is3EMWR1yOu581kTAzIL9HmU68SdlADWHxsCpj+4LZaOQ
q/sn0ZN7msyZjOl9wrTRIlKcQL0mlZ2Rw55XC3GRiFCn8rt5Tnxmyw1Un2mv+kCG
5yr27sjyy6bUgzOvuPVYXXKytn4dAt8dkImiRl3RHB8ONM3s0m/LDBbnOXVOs7ly
dNV5GAQJNLCNsxM0MPbfyz3caq4WQqOXDGqQx3OwSsni9PFnVskXhyLOeYIUoaWR
haACfjk0uRNccp/RizpG1J95aHm8zzsKuNOPyP4j9K/ZxoYtAOaQRNUAA7ywZTix
3D0Ar57kkLSiWrHunEYBz87DHItiL53O82ZubGmWZYlS6saFiiWmmXtAjoAuzwmI
INW4gaJg7se35yehm6ARbcIx2SnacyW/IS1VRTQT9iEl/8Kc+Z1zJ1q+JTJv9UZ0
aD2yYePwoR32ER8r2zVCqmCq9Y1sn5SWS9E3SHI6ca9mHv2PRX7kPiBwBkTLDH5U
W7Ai6KznxzgYohmmcES2tQrIWHam1sUjBIhekWDmNqN8mQGH/VWsbWfcRfcnla9G
sgU3XfVVGbLuwJj/IDXeoaHIm/9PGX8HUJr1T5/LFM4yj8OSa7AQ3KK8ckCS4HO9
2hhYJ4KgtdtuH6PbRGUHJJiT7a9EM4jSGnX8cnyu4rlPhgH2kCZkq2VV5UtXh2FW
m8P0LvvxINvNablIEPMmR1yFpSVSgYFoTCHLrP7nw1SD3a1HsiXIwEBoAb/k4rOJ
1uQQr9N2qJOu0kYjjD3Se3uqZLdQ77ETo10UQ6fKHM1Fu2kHQyEh/TCip82/EWFr
07KDNorl1iLUAJuVmpZcosOLp6IX6LjeJDPZ3WcsN7BXDxkv660U9Gj3tcqODH+j
DLdjONpFRhwTeiRTwu3PyEPg9F/Gfkl53RXquq1IJ+yFTTniSBs8ZI7E0N06ivaD
UTQJyOZSgXVvvUk07EUEKYhWR9KtJsa8CDm0gMFRQ6DHTzZJ1DT3/d1xCrYo17qA
RNTvdFKIpgeqABkkzFNaCdtSh0xO1iuojwg+CCTXHCbnWII78e/ojmVBTYtLgrB8
bBP3vFmzdjBWp6TjXQI424NyvKJXbtS4Br1sXfLD6R58Sc5gdW32c3dlECE4BYfd
EGW6foYjizfAkyQ2KuISHpY3psiaAXhqAfqq6GXnJO84K37cMPkEY5oDdrfgYiQ0
McTGk1qAWlVzW+MGl/9ot7oP33dDVM0hAObDp7mWNPR1IHDJE94KeM/lSuWXNLEi
Mf7u2oMcYwrsBsHaTTtS7X+S7LOz94eo/GBi72vm4BfACfuaIylsKfwBoCPbqQdp
0ngnH+U8Dh5ARPZLdoG8h4r60mPblTCgBdmIXEas75RLrjFUAu8UNf73ogDxJ63g
xdtMUIlfwOeCSWWiUb4uxlRl1dUjd86qnPHG3oqsv6eFlI/NYWu6ULkvdZu1q5fy
4BRDUz9cvWYQ+HWaeKwdLlVAFssiyDexLv0trJXbQ3dB8wAV8LzsWzqBtOTASVZG
8NCcbmeHU63bdkGmjrL938tTTJknaNUlvV5hMZQCb5FF3FmfXB9k6b0PjN0z+4V7
HSiVc2oUx+CgWFmqCaYx0bDmp2yoZ0MyNYE0u8LyCLaNiR/2XmL4iDv2F1gdb4KW
hCII9IJ560lcM9wpYNPVIzCCd09/MHXcRir/D4F/IEYbqWIQiuv17NBLY/mbTHEd
BNZQo65stCeYPnJ1Oo7TvORfDh+bTspJVzVqV1cHGqeb2mbf0hsbvdbCDuYL58qO
2vhs1SvPKbsUIhOKl5nUDA77yuTjdJYF7mfS3Fiuaorw00jpx1Cf6UAWE3r4RmbW
YZBst/Z7h0ygdwHzHvFO2G46vKtXzDZ2uHWqV9wQ+Bax+G89/a9S8/0EGDpSm8qs
WmFhZut0B7d35aNIuPS60zrLilISij6NQ4rQxaAEGOKeFUca6Gcx2pjl0CDCIOXI
uzaGJ6MwrukubnZCLqA6XmIsETYCLITftgxttk9LBTF4/z/J0Hju2raJGvknN2kf
5FYvjOvRucWzrzS5ED0xF9mkf/HYLFnjujfr/VrBEQ9GUQWfFgGB02ZYmCnE6593
XagbwyKhIIgoo698toZhITrnFbN8A/GOwqOCMCswnr16fTIQ7VOO6HReEm76LJRQ
TgPWNo7YarRMgkd8uDGw66lrjOrTn+1K2r373P8dO0f5+LNld0KmfZzfqyia2Ett
4zGE/k2LphWCo76+/gTFqMVn7PF2Ro/jO39yTsCQJBDebewDzx8RtIA42Vv56af0
V9KAWQZ3S6/WLdnKmfR4CA6sIrYfdhCwehFsCl2JhWZqbBNL1solrhgBMKgFqDBU
zGxuWVjHvBXVZYbg3ejPqggnIyiYx2E4wS9tg7STZpBULZ0SbpSqbJ+t3UmFzBbb
uSglj324/Dnux6mGSo5EtTRhH7/8EJ4dteMiRZoxRIQhGeXPa7JsjLV2HfyhIvOs
8ABN5wmSZ0G3kEmeJC8b2xN1UcgzxOqgUbPECQaab0t3f+MRo90ogzCBH+fBxgP2
j5i0s/EJhs2insEuKc3X/vSURedYxFxcinW6jRCyObFtzcZpediaI1rvyVgf9is7
x/UD23a/zlnDKNQniyRNh+MTzSQYLq/UzfIoPt4j8iWV19GNe7sfmZtd4Ye8mFHa
OKGGApftWYMxCQ8BdcRlh6G1OoH72pOKRb4khQzR3y0G5+75h9eS4cYcy+GHG9zd
lKOI+7D65M2nzFKvQngGITTC8ezjDoHoyUJ2fMPNpbHUG4xToCj688VCxFf9AMCw
pVBMZj+XZ04/vU8WRerer/yJiEZHBppAkquQzUeZgHaKNy99Tdf8KJFoy3qyRO2J
qe3XQ++yDw/k2b/ATJrHZwCNZ59mgpJnyUN2Q5m93t1wQ8nC7BnPt/UmtDFarDqt
NlGfhCBRMXzK1IBrO6cV7dnnddH/1DA9m98+syyvmIrHijWlcgEY+JgduSja6w9q
hX0hQ666b92hTAzsN4Jt2eds/LdmfM7ZV4VFdPhg5TqUf7uweXMS/JotIoGYgS+D
kpPSsBhFh8h/e8cQA32UpA8fD67hf7MUqSeW1HqJlKw56L81OIi+OGc8xlOGYTZu
R9GVoOwnrcluLt9r9d0zI9QDpqJ9fhwc88CbIW/MZxhtWWqMtVjMQ5yX4qhabT4e
CzpwvlePjjxEAF0l2gIdrqDR5DJTDp6wEfXMvw1LMrKIwCJ9OxWHc9SyoCfl1xvZ
pwCNbWk3I3ngsxmxErnLwPoplk5n1DB1RIuhvE3n4c8q8r2w2YdmgYbf00cocSEb
OeKyLrhnIhyVZveq9Rl3jW/z2VW23HoU2T2RYXslBZlLpqQlRt4eV7WoyU49CMiK
2cF116Qq6j6DE7FNzkrYJKSgPE18niGpWC8E9PX/LyQIEQlUy+0vxkrNbOcPjbGJ
GKDGabT3IbmAlM03mMSQf9ASGf5AWzT5Sg425XKj87g4b/yeIg1qsyb3TjGnEUdK
S0sUneHBnldEc9GGxI4GqNlyL7LXMjntnQou/odaaIOOdKWaxJq9WJ8pU0QvHtSb
KevhOWNxeBl/fUWBeSkiRYnHutBQYzkDUjPDDGpxx97eRQNjBfPZ9VkA2o7bifiA
ZszLm+nNhAJVWqMEBjZvHGn70c5sg7PXOiEMKnBmFtlhoqckkWLq1LBcN6dkD41C
RG9LSYfTggmSiv5lKobaLGPJ5bpYq2xCmPKoKOpRrdtf7rOQ3aEx00Rd76/ow1H6
vi6NGiCEHhQiEfb8iJ9BTTSjobOtizSXum+pTM0vFFRuR0UPklLi8czzgwIFiihQ
34NxbX1CQyKNtsGgz+x46wjsxnIkht+rGbv5izJzwtC5S3QfJRVOma3j0E5JnWlA
/m10fAE4il1ZUoD3Woj89eI2laZ3lWTNoxGK9iAEwDK9nDmCtQgrpaIGP52yOGjT
0nSR35hmPqLwt5+/SiHhaWFuh4uNxf+r6IxDj5rU9U9O62Gz66biTnUXcc9xEJqh
vFMl2eX+xy2RCoxwmBnbYPTpTqsCZrC3MeRsQ7Sf6FypnD2kYuu9g9BvUOQqQXaU
79oBh3+wGH0sQcSyPkuiCRPlECsB44gjINeAULdIBeSYKWQTUtGRTc7zVSe68od9
fqAB+Pe2vJCAnj04m95rYDGKgJf3FCDWAGZWAL92piKUcWS/DAcpsMCt5x81ksF1
zIEeJSaRGMIIUySNs/R10ZYFDV4AijI1jbOWkY9I87z7h3r6Tb8iBIIw83PRJw9U
XwpyQ2TR+AQi7ekhirhSBrt3vqY1qKauc0Mm9/gG8zCRRRwVVqWNB9Pu4Nx73LA0
RHVkw59sLdsaTFeFJ6Ny1NcyopTxGY7saSJcBQ+frAcjfeiB6Z0Jwy4kwIrJpp7w
IZ1SVCVp9FlViKiF+4x0QPGPjJoTmi2E8voMPQEBe+p8bcDA9zHN8sFMNLYyUGRO
qPJReOBgM8N2hpxGwtS2gN9HaJMIkPhypPq+LCaxztF8KVBMNi1R1h4m3uKhvRm9
OS/S5NebU28Prlk363ihdk5UMICwf01I4ZlS3srinC+qGa5LllyGQ019UcXiuP14
m9Phc6gZoTU33oyCWf4P1/KoRJJgvyMzlduW3PMGJwDFiQqJPKw76/J/W6uZEsc/
+3JjiOx5oWaN9fzOGy8uNs+WVktXFVngeN032EtCAp2Ec1SzOxdqHM8T8gcrBVC9
6NbflMBKRyhumTzwhFuqJ+gl1FxJVXuWQxIzZHw8YpW0ZdNCQuYL3TQeFrMGWKUt
Q0WvFp+SkQfPo6eqIzGliyV+J9hDgq/pp51JgYXoRzmdtc+Gdz8SjUAFt76VLCjB
T6gitTpzn5Q4VPgQYFCarSfKz3OW5O/sfJW1X0y83Xwp/FrQzQ5a3bS1o/x0XSan
Em1YGOY8SO+sidHvtRhglRFtu5SZUcXmh1dHmG9RCBYnuHDSBteBl9g5l07rQhLW
AIoATQLs/ccqlk/KS96CeYYG5xgFIx5EfTMcjmIZc88Hle8buxgRn3ue3m/sH2oY
v0/3HOfTj2XbGTi5Gv9dd3uPeWZTgHMtMZTnXcEkDv6H+lMwMpFr+8eYaK4KVggm
oHi8itnfJ/3usrvKOoPfyfON2WmKMGAOTaJVloYq5pf7ptDyhRpHKYrexk3zNYQ0
Rax05nCEeYpq0UoW1qWF/WvMoZa32PZpRL23ol3Ga3H8T9KpANUbda/PvqsEUIl5
ZwYUcvPwm11Lxh/ysXpMneOW6Yq28VSsHaOPlmfNPaRAP+n2Eg3xrCmSyKFvCsea
QX4rBLppDWrCEyxNyEZeECtUMKCfwfYwB81pVZ7VZEXGXzz620DJFd/NVBnFEmQz
056R/3TWo9/wkEmVNnc/J1Fg6gL7PtdVh+aVC95ZVsR4QUp82qsd5cLOG+Nptc/Z
zCfUQcQaQU5vCnPfY9B//rBiSxsggwzCiTJfbAkvVg4cKnmJ6+obXAKOJ9kPx+wX
jaSCUyrRF0YLLKEvBjUPUwWnCKTmnEhhRezrA7yia4pAETINMNt5TwGjI371TMBy
nZeKHP77AhQcUpOPMDZJzDrDgUGh1xa5ypdudqbKxmBSg/31obP4rzp9p+Ira4t4
PFKVpfUTBr/n5CO+NzzoJF3e364exBbRWp7rqdTMOj6CLReOtJqcE2Ai06lSqKmD
JgNdiyVhLedxThU8Mw2yc5yYBOS0ItMGIDqiLrKAcSm5dAfuAZ/2/4/ahHKZRne7
Yor7KSD+LbKjHd+Xm77Z0Rf/QYHnQIm8ljEhfpGCm5Tlafj/d9TzpOhaHcoXLdBN
/qq09eHAzDRF9EAO4+FNvJSpNVROCnuEd5+CZpQSIS4aVxHPPs8KAtb4/h+NpVlU
6vGb7FNj1FAUWjPhXG538AxPOeRPvcdBkLUaNawP3oQmIWnJffp+JU14UnfJwom8
pxXDios7xR4F0bTFKKXo5yDBWjNR2Md+/hX9EPNW5SYCbOjj2rMHwSg+Ee+2bAGt
chWH0lhSYttasMVkelCOW+tvSoZtnyFQnlaDQ8DkWA7AeTgqJ1OBMyxt34ee199K
hAl9mpCGWEsXDJlIoG1MNsNjVHReRmqBB7jkRG5l5xkxfPP8LJkOKun8d0a46iZM
6TVDhYLMJ98lExgFNr4Awk69TRv503C9EQrIg8q9xWEdkZRvT+cVz2/839bvyc7x
8f58QBRS1aVn9x9TEAOvHDWeOoc12rwfL/rn8V1A6vjU7GypISyYHhCu88BDoUjp
Wg0ej5sxSCUYTQwoBw9j1PXinsxKeIvJgvGXQyjS/aa68jfky2jddq3f83y3oFNt
Y7GMFOXtIs0qtw99tFjhQ0+jz3iFNHOMrNols6iiZmBuFll2S64vmNrQzvMwaOhw
HHILobE302w9eOktlZq4fRQaYEqIMVq/Pa5MmD2ymEMPkEUdjm1b9kUZ+5a4jXZV
+qm391MUO9ID2KSEi1QYIH0nM9YBt8kiqUjj1y2v18qqYELM0gcc4dOfptSoR3Tk
NskMHJvsk8CDHWVaAMLcgC3ek3qhXCDrA7Tg99mWEARWjIy3/bil0sE4bl6aLa3I
kyE7eIKAJK8tcUKmMi+IapffvHbSuumlPoW0dr+S/1Swj38SlZ+iTAF0QYUxoeQQ
xvlipo6Jjc3QN1zS+d6EIKUUrL1CR9EJvjK0/wEdIGM4lGJbrgozNtXKdojJ3eNe
q7qyn5YNgYl/bhgx0E+PgNPxyjsxg5F7e3xIVbiosTVeuOKhSuYU8HpHGvVBWLSD
CCl054MthbHvUqeIglL7qhyD3OkrI+qZxpqSS8CnZnnRqwQtOXvF89j/Ctl5PeoC
OCrONFfLpR/0+6qvL/vDq0TjtDtuuvIb0Qkfn7RYlR0PZW64wO2vlHM3NZzWCaKe
C4RXL72iGY10OSJLCVyCUxNWpeATWxEStntjSLkiipta6OpJ77BN/6bRQR+qxSK2
WRvJ3FsW17wVLrf1sEDxTCdvJCzsKxqPpITzjB4luHVJ/BhcQrFogbjkUtldfU4z
IXANWivOasNiiik/0gO205yXChU2PZWv/YTPKFG9J9zJXWGqY6MCaWvc3D5u6vSJ
/5TXY4QDhtgQ8osQu6G8vbjZM49+nqR9fesAhp9xZbnpxlcn9k81Pv3kNXEecsQs
p1k41deZvg8D4bPOaU1k8rDsBckdBJYxPJEz1LJm320C6LiHcSlgUuZECmYPmNhA
Ofxf4PrH+IXbdqpLEpnqBkmmxcXIuV7l7eiitSfQPzlZ5MmyKYesB/fg4cWK64vm
bol473TGA7n7tEeE3p2oqaGhY0Xuwyhp36jY5NLQSOhAiVY5Gd/eFZsH0+cTV+P6
zK1hYPNNNMT9Cao9MefqPvV/HNCvLzmNWHkxq2mEDlWLmvEZ9RxqwL2Ug4S8XG0D
YW4TCVyidfL0yy83yQxve8E234BcAdkn208RvWLY5GNECrtoF3PeEIitPeqQh375
OuyMqMnhUfmabLRr6VextwCGUiOSv5ZO+sfGV01e1r3zRz5TJaQDZIO4eIEwPNzF
HtwNu3th1mOOP7Z4mUGk1qIU4ADZ8RqYiKJo7srpF47Q6GLIgiHTw8wkj3UY6c5o
krp1xeUV3Z2s7U0RSet7Oinqloz8dn/oJZj3GFD+5OYNHaSSikWf0mcya0+E91T/
7SBYoo1bXu4rl/TNd8vxd7c/SjnAl5qtq2UHlIqX7XqdmJ41t3CXXvQJvJGYVInv
myy5hmoyot1pGGBhR+DP07pA6q/doGm/XNoaF48HWTYgpFxX178eDdkxWDnc0MrE
S0HDePPT9fmreRd4JAYK2LJ58vch3+ts+M9mzLFs0PVCUa9k/1TvNsAz9g5oAKiq
aK/Dj/Yg+d/LOK4xID0V+waiIh0NP5yvUzj8nvTXWkSlDOIaI2YU9xklNcrU1NmB
936oods8iM2KSvzev5O/iDA6rQJs3SXatD7Mqp/RIfcwIbZyZ1Y79rJANVz3A9GB
yDrz2rSYwHrDOcINoyUIaYQNKOOvRaX6ixBtqLCrbBrr3MnIvQuSn/koQvrSI4WO
tjyb+mAAPgTJBab4oRymNV7Tnr+VVYEopQR/oo/z4Jgoxn6PpqM4OHIP82882FL4
3aL/0Trfb7viqOIVBpNFRL9aGhOQjg34jxjJyymhFcy8cn2EXpfcX83mNJpD3KTN
/G8lhG8G2qV/KrK3cXN2BF0AFtCKPYgkmVyPwzXnTAYKymOwH2x+anoI5DJPtZVQ
WNlybPwXg5QNnKwk2p3II/yNQbpLchrXYIR52ShF88Zziy/jE2sIpTQR4OouVLfh
ySWwhyVyPeOlSFNLv7x81pn6orrwrQi7WvrAJrQAjnlPlA224yHHGkbSzbUcTuWq
9cJoPZ/xLBqLHJ+46QYzh7u25kWgdF8HKQscjA/E3P+TwojfjWol/eP+lGsfuUze
17DrzT0aZzy2LwOzcdXQ2YRY2Jl1wxyjt+YBYXlpj/ZpRtU5unVKDKE8ucaXew6T
PxdRWFovmwIUMzSslOwuQ6uJtAACAgbUfLzg0MXr8KamQzl6DKQTWUoQVq0g7QZO
rpj/P6unlpbWSkWqCZFmBCzGoysGjxuHH9JMzNst4lIub9sgLtqImbp8N4gu0rkz
NFfHmYmAPMp2F3YvYwDpetnGdYySr2ciYlPk2fQSgrBESmfAXC3HDnzeh0aM9HoX
bipI9z5jedsg6YaE0stFF3jA1zXyubP3vn8IShNnDXVCwQBBcr6y6rftCWoPlIN3
9RCSfmiiMjTui+1ps9UTR/xL63Rn58DXT/s6dUL2gFWW5u16UA/G0lfpWrTi2yT1
gcq9f2GOVdNJOp0pfHGLkF4GJnQADeu3R8dOc1GnFwIJiy9f4Zx+Q2OvedATIniJ
8LOhoL6AjMRpuCOTBwGAExifcJbCpvBBoWaBvIbPquaJPllLi7coZm1z4f4gidby
BK3CQshto8cb3RvrHhgeWOtpzimpXKZu9/dsLbraN5RrIm7gBEL0FrrKk58H4qGY
`protect END_PROTECTED
