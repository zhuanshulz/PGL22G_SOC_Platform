`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iz4KLB0L3E6K0B9sLN4ACJCwFPHQJO1AoqP+phIc7v66oMukGraqyzhOuvuB45k5
ur+u6OXFc8+AohCd70skHafEw1J9+RHrnW9EJ54YDY5sSVbJNDvyh0o7YaK+fJfC
zBAOUU2emprsyY8CjeX98Lq0kBOklkh1wZx7/sP9uKKgqcmSo9FZiHl78Qg2AV3O
uTZ9/p3VGswP1NmRPMwAcDDA5gVJh2KbyOY1VfmWB+m1K08g4t4wg6x2aNdeShwC
fOxscDlPIpZiF2HzI5DgRdEFH8pF0MhHRIosXirxKMtfqopuLZFmxk63QU1BmNyW
EVnXaDQ1eneTerwCYReH/KR08DsPt7Fh14bV3p30GJpBC57Ki5m5qp7Fxl8oS+RJ
hvd7bteS9w6Y8RDl3NtmJyLwEU+Ex5yKTsoaaL3PdquOepdaLXs7RpU6/rmxKsiG
Pqy5Y6YQBuBCfU+ohjFN1pxbml4h36gO8AbEMsVYjyBWZQMSfXyzjAGdJPMSXApG
ryZHXGMJpngwaoic2pM5rv0ZlCsEcJ44QGXE4VznqueuLFNh4BUK5wfq1XQlB6Jf
y4Az/Gmn7zFfLA+b45DHDlFyB9DsemaJGH47b0oIc3aoZ0N0h+B9aFJpCD94cvjS
VRH9osPac2/Wt3A9p1UNoOfbUbp7Vk4+txjfE+EV5IRFWbC1Wf3LNdU9Kjz0IQTa
uJDv3bjdAqVRH6VCGgcNhpnRGYgeCQiidJR2bLmvPovS3pNuDCj0smtCHDaioxE4
jOgd92AfHobW6LbG4M3sT9F0Db4nSuFd2XWVQT9N5MuunruyGS3qf3zMIG4SaMJc
rtFQaBOyb6ZzPsL/I6oMcdwmz4pCUhOkfc5KS6b24ETmyTowXzTRcZcEJ5DaC914
ilGncjft/jSvdsUBaFPE7f4aMSqrA1mRtu/IekNz9UzSZFEpRautj29e/u037qrK
+bYhQgpzB3arSbRLmnBJZHyQzw1cRm0C27UGo6TSa1PnKDYT6y6C2p9HuanwdQzI
93UimGKXBzAmIgKTk+d8OH4lWzFdmDAx5EbwO13VEiR2QxQzMOZNUf9J10TqTzCd
D0IFeO4wG/nd3mTnYmFuH1WuJo4CMuZgmv1F89eBhLIxgcADevq/6N8YfGpshScO
FJTf9DAl+LpCFyFx/kr8rsimHAl8Dy1CHa7HrFgnT5d8mNIx3MhnTXua6i1XVFn+
BCMLdafjn53TNso2geBTtikBuXVNwYQ9tziWvRYZJpm06v7QAUY9aIS3y4OIMrC0
nBp72XgAl8LrEU6uDXahrSclLVOCS3hr2feZ9QHfnc1t9eULSIX8ll6N6L+htmnU
7MPcQm9T1Mfgt9R4NRHXJc7Gm90H2X3mwNkokijFm+pK8ftiQMekmz6dFxgbPf/c
0l2qU5fuao/T/m+T+ZPi4y72YPbZMdLynCI2Sqx7znx9XWF23vc57yB1UB7Bf7EK
vfVVzMZaSHjk1HFc9mbeqahPLfFyjzqEkOeEEPWbHA83yA7LMW6TPYT9gIwP+q1E
IJDd1ePIw5cTsykmV8eZelLmEDDyrCLiZ+vJJIF1sn0g4MFXtaREarQPzpuBNcRD
OQ8D95z3If4D1h4/JpVAQK0af1ysZtVyaRjITWwjgA66LLs/3Z4VdAXkUDH2LsUD
Ys1u6NmECsi+ws+Jpu9rsWgSioQEGBbUFd2CoHDniEQqfWupJVRXAjH6x5t6Ro+K
LSpVPcOUdDxGzeSh1L/En9bDkHuY4IQTgy/rnhya3vwqW1CP+gW5oZliAwy1L4Q1
3KyRrcISckUbbQecMlFu9dL4DcoAGgWz1p0Bt+GO+8CFTcD2zrwEKaDkr2ZH1aCm
jJyAolL5X8ODHpDpRWh5rllVoOriiedR52N+/JUlimaaXD57XbN343aNfK3y9Xg3
na4dqgO1uPR7G7V2deYnYr+Q/aQDvExw6EwpKyyh4wuiNei8i7/iYBl7vTIq9Nos
n/ow3DMWlJ579Lgvon2fvj157Dcg8rWCxBQY4AU7uLv3RpuW/Y+yIR+EzbccHEQT
xRrWSYN7oklpkhHb5URk4ssfV1YUJ+VFxsckj4psyBlOknH1uSS4MB2leenbGYi6
depsVk3BAcyvcxDuaqJA0OQ7oqdSzfixNKN2KWjgPyoNkuwr10WIeRcxQkzbC6vK
1vWQ7yQdi86G0Ni4YanneV8eev9x/VgXCNKpMsSq6bOQC1niT4WRsu7qBO9X3cSJ
m3Nkt9bSAZIs2jM9x2T0OaYO87YznCuDYb4xex+Ll9J4t7AYieV1Jb55dTQnmQPh
CKRXuTIOTm5cAVSLiBNYMLeBX93qaYaeDD3jU1WMtkcruVGbJz+SNCdMX0rfR9/X
wXbcBn+piaBueej3zpOB/CFQGh9PN2/s9/KQJTDy5+bc16Wzdhrat/+uwIozsmrb
DZV0fxW9JAa/Qxzwb5fr3rozgvpdX/jgono2ru624DhtCbMTiXQ8amDui/ePMqfS
ZJUpgfScHQW4gOjVfTdSqFx3O/FBuNHBN3xbwD221PlhfhX25qP27Rtg8WS/NFHP
yChvYAgOBWyyC3QOjYAPUKGCJwFHgOyuUgmzEPjvaU36aoChJdPbvvH5iUDVBmrh
UuhCNcsvZ5sDY8yiK4qPsP/kXGXUKhmAWppzEYGI+CA5mzINYBpqmORiCy15oQ2c
T1CrWtT6MICCqzk3CZ2nu9sbTwTmsLFpTec06EeDinyYPVt+2AWUeo4sSu6Zy0LI
kstpsmwii8Zr9kLcEfSFP+dk8qZVBYOfxTLcFepEcpPMmQdxA0CWaMR0hrA9PLrE
M1Owyk4Gm5NylwaAbP655OzkfEcDQFgfyNA15akoa0QefKJxf6LMpJFUrjy6mpuR
EMN/aUriwDEWQYpZbT0JDhjdW7ydvk7viwQs6Rzl8OxbQAOpHeHi4rxuUjhznHzv
M5hevz+86SOkmOljdrLZNkQfmpIXLibP24GORW17RPjING6IGPBlbJN66WgmwbzW
YfRwkOTGFFc2vLg5/CE44j0e+KeMP7b+l5nUSXNh7en3fKpuXqzDauvugRFWvVik
NxGv+zjU0C+2IUQNYCXdyP5c8vPAfH0+EQxDApT+z1UawJd7WA8FuLSK2u8kKmBK
x2ODEjz7iM6gamK12F7jSJ+JBJIYpqpiCNl5DDnhTWm+lAZ4zwZQaGgSHe0O/C8C
6N9MGtoC26S+UYzmPOmszHyn2EzTQwfOvND9w7+N99UcfjYkAZjVN6lkEjDVIhhi
kH57MaSLCjowa5pP4VF/N+aR6Dwx6wlZV5nfXnLbZFsf+w4CQRoaVkDSw/UmGhTY
2GGVb8JTmJxvCD1WS4QyQ7FbRUzkVzhDgZ3Ci30/+Vau0YCijZBN6fQWfyGR5ujH
hbfCOxrwT6WSrE8Aa/uI+HZCb1DcyvSNJtkOltVcvqKHDm/8fOk0uy6zX8EF1iln
Uxv0aFwM2zan8alopVaz05lF1jIGPW6VrShRe2MFC9ks2J5UZRbu187/DKcCz2F7
cHmip7J3BonyuxduyLEQoKoThkibVzys34LPbp381QjR5jXxdvAD3IuPe2FOs2zK
sru05IlNx6ohRdUemCKT+K+ZTxh+fmIL4Kgli5KlBvDAZjgo5SNer+nkVrZJ4y3V
4zATIcaeQCrTMLzDdImILl0ehNMsp9A9Lo+B8ZssRtwuF4tFPI+Q5sOYAtTe73Hd
GURuL7ay9rmE0KzpHKWsVJBjWYTcpddu5nOEXCH/kT5rCSjnoPZajVcNxHJjxKnl
S/uGs+2RzEHlLN7dFiTCQOXc0l3GhCpmGrAtLYhFj4qNCSHCGn2BBD1WviC7Kkap
JNpIBpKXr6ZXa11xd0XdMznvPiE1M7w9KiPO4pv54KRI596qS52Xwr+e6JQmWHuY
712dfoo6Z1vJKNX3iIzf8iSZ81RJ47MM6SXuykT/JDQJHDxg6XWEZa/GvVijYb2T
1DYfd+WSOq2f843rnv93YOY7ntb7FArM1GVHR3IBnYKKJ13N7T/DB7iuU+GYtU/J
NHyRLCpDgHhcRTKQTLfTAcHKEw1jtc3uzmdwGLZJadG1CCbRc658AwUw6j6Xi3f4
9Aq/VwrNReBr1hxEd83204nytJoCeTWwQ8Nndwa5PlhEy9ORHlTq7CqcZjnxo70s
VhXkwrhgsezklkmrcAOXQbCWKmO+tgL3k3JUnOlp1bTIqL7Lo2HXvWOkcVB6cxTl
nYLCZFOKes3W5x+qAZV+kpP/55zuF3f5qFknnyJr/wKyhzKFp9JFyAcUMT2DdbLl
5s0zTGKTJxFQAqVqTByyjJ8GiO61MSmqYMNqLKIrB4UySeOdLP9yl0/AmuRNrM7Z
/VyimFRX24bzWZxc1UtuRmOjEE4Lg9VchQxGfss2rpGrnlw+hwVu8KeS6oy9XuNj
eRd5ZvUOK4aLPEbJaUuva2/tsX//9zFsoyD49oPXHDGyFYkYq1tG2qPUfdOXhQcm
tAsdtZ8QfYUFZrinme5mfDGt3/NZYSFNunj5tVPDrrU=
`protect END_PROTECTED
