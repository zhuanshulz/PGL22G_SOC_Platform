`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kVMCmdnwMbWhtGj6TZgoylo7t3QVNTwws/4JAyHG8GbmOj+UCchJqj2YK3jICKBb
+sDjo8mqHcHIPhnbRDXlu26h3vymTGAKwTMhHN2RWLiWLV//oEXy3m9sOObzY/eJ
VFhIcnnDSsq6pFBWel/qDVfPR7IUCsNDHBegL9aKOEblUQCMwwIdphN/L4JI3P0b
6Y8CnWrx6+J3FroqVWNyzu1ASu23ehk6doVmT5yrVy6MT9TbDaofLvSdJa2RelsC
gx67XvOIYTFsLjAYQiaNvtffmj0T2544v3NidAE08Xx8p1AYAwixiKQr0QVH0r32
WyoldJwwhoSLQcOS2/nkIerzV8Fua4lv8/F3WDFw6UeEglVqyNUejljM7a15KfPT
qfsNwpLT8YrQ1FEQndLfncaPvgI5wjeM5MYrolQKUW/gfMEllPTad/XMnh8DcEBF
UKK86sE265WKEITW05ZDmA5+6/MxGjUJFD74sotQ0drSYn8Kn8XoqDqn1wSSdoih
v1d6EmM2QU5VtwqQmbrkcsi22YJFgq2tnNhQE93H4ruyMcLtHkxQXaTi5QsF9Yu+
RGhCmCaVFGT85hiCWEvjFvQSH8F9zQB8+xQ6rpAQJ/bbOsP/rggKRrUWtqyWJiJ+
kytvHHwOf05jtRm08ecc1UQaK6f5ECte0QYwHSIPjboTySpX8+9l0GOF4fpnWLtZ
mwd3ZFdSie2jlz/eyIhQKdLDrbJN9+xSnCeYsPbExib43DJj5WheT7dClm49t+aW
e64xfTXZG9VEqPK33NzO6zPg2eJA4o23DTxZmsVTTB3yJhbZIYn1pOwPO8vb/enf
t/BlSzy859YVO4MhuQzhJdQwXMcCv0HivOIykHauOBpoXgshjhUkCVMwSOPuvBlm
YAZ1CPk15sH6yKjRiMhqAHhmngkl3TdXSZXx6xluQaSZBXQAVXPdWAqE7mqkIK1u
aynXDT2fF52kCDTbgSFLo2m5WjgcE7WmIRhVjIapb6IaxSQmLqP8kFHufKx8T+CB
4WZw0bX1ZSoLbi2rgGAhIl1Dj1dLFdR1DdAaAfTlIbtg8OflK3DyFoLvCQ6sNMp5
MjFdF5bbcX0d1VjdKcHS4CeNTwgzPwgGHHowsDI+V24EcmHOonhhW3OoqreNcnUo
jPeahqvQa/JTKghYNf8RuuTaosdwhvKwhMnO9CurntxbOA8W9fejZwX7G2a5uFUZ
ER3U0VmXESl4Gkd6qwCYqZgD/p1pxac6norquXLzv7EN1+6HNwqfJOpC3VN7G/pp
tl2l7XXQ4/+MGmv20vh/MLS9kGXpf0ckfl4TS5cruiLQguvDV1CE2B0qGdRuOW0r
6MzXthKBloKJIZlJ4PMpTToreOOG2e8yiVPHNDH2MSD6Rb77LIUlcPIMaeyyMJKW
Quqmtwu6VzNcP2BS46rUgSdyuNR9sNNVyr0LAHHMSPcJ10gFRDt5hD2vdligOH5p
T6SLle1in0ZeVf7ztQdtGUUWkWu9b5UuefK5vQSxS6E=
`protect END_PROTECTED
