`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SHNRQxc1wzvi5Q+j5TqxJHpGvozhUFn8KjL9zgn9Xe7uAg7sbTu8eDOEwFYheL/B
jJRprjZqGGxsJ5e84CJiI5YbIxxJCNhmnnEO5ikerW2g21cOI0EFjKUYqZO4V0Ut
oel+5zKPp75/B/xZ/vnej3Bt/HATnRbfimQlum6kMwqtDa1ZHoDNxDpt8sa6EeDe
FVq+4oaqwZUV5ORxI+eiMFmupTDD8Q+ldpMO5nJu8qTE4KalQXKqKkZifToZYfFD
trLxOirMqaJIFjTTPoWLN5KPj7QJRd2atHhyXOSrEF7BFCppoQWhwyKCxB1KwJ1p
R9+bY9TQNpZ3diNpCTLQlYj/L95H4lveh6USruQ1tXlBWSDm5zJRIk4X/byQZU5x
6ohy4DexgmUFhobzxwPQaDgmZFhGl80SJR0p2FfF1jgKWGPl6B95TcX593fz/yeJ
9vJqPdE+aLcZg2Vie59fabYuNIBzNPpc4SBwa4CsJqtlSMqe/omXlGRUilf8ywxB
EgS3ZQuKjoQmbx0FAuHeyFZHDbFUZzplrew3IJ34qdbJqTFxRI5cfIkLwWB9WAIn
DYmSzkmTUlJj2Tp6GPbmBT3hOcGmswtFL80CN/epJ8EDBfK0dc/iiNsZVzcpVFJR
1ePGpxFoY2jfwIAzSGn/DIiH2ivVQwGrTyIL6367BflXBolMb6vkubcc9x/PdWtZ
gpFoT130qadJyTiexMNBGABxhQfDevJu1PZSeuqkvvkQYOkDV7OrUzJGFJIR736T
AfnUuhq50hpQimSueqawet4S3L1nPdtF8nuZLPHOiCuXZV7X8S2To5l7bSIlp6H8
aZT0DLOODlhSdtl+vQS6PFcYbWxKTygswrKsXDX8SaMaM8ZLVnaT2Wf9Na9QGzAo
6+GcA5RN1kDtDvX+6GGQj8XjNVibklCeSQExrUPGoDHlZ/pTNiCrU00slETy3tVT
T/2+puYweMxNqF7iy87GbXmj9bia3Kj2JaM3RmlxTUzyyo5ezr0Cgb1Q8ShiD6/R
gtI1jEnhtft2XKxUsxenmFc79cfZMbmUM/3ISP8W23ZD+s486vmBaTA4JIFWf7pr
sSkjy0TxRs5MCYoRedFqXCRvE3j2v/B5UECkZR9d2hP/R1VLWGn2ifYCVas2lzUX
CbGtCwqoFuVJsu67PHJTVoXdNOg8AHp5M0drxB4NVSwjHwUG61B4y5ipcKntIkJU
j6gOb1STqZSREIqZXB5/w6RvvsSX3iNJNHVlBsq3au0a5+KWdR/zJ7KLzA5HPD8b
yQtLNkiruCUlN25uS80wIyhrGw3qFdKw0s80rYEmkuAYnJzyW/Kdzq8S4VFwW3fL
LkaFTxIpwIrgyu7nDehTBVW66X8gfuEjlvFoYU6RhLTRUDuOdY1TdxyOMnja12I4
vFwF9hdb4TvR8q8+6xcck3XIWr+82YnanTeQ2LaO0F+vwJq6IaWC8JxBGCJBTdZ6
+zmWFSlM151eq8znHj6d/8GHpi/eOQibd0/P8Zbpt7nxi0YdWGCgVov93yx+aALw
GmXGJ4fshgwENwp1OmtU7FGBMrSdbjHbimSAI1+L9VMCWd35tGU4w1ldHYN/UgnU
q9UkQzfENH/91VqkpEZNvqETr4GjYSapvotYIoMQE60tlGw0JblMwAE1DJJn5RAH
o8sPWj3j3wkgEgH4j9D9nvNr2hUaoSLvRzBwG6O6eTUaa863lwOX6CUy/ihs6bdL
atanzeTkbCsw1Y0eDMQbwhPopLyNJ4KqsBReyomqZrDrSdk/4LLIE/jIxCQqe9gN
yRFbOWHk00rosr4JpzPQPOLe6xM3bD408JwUPHkD17WIajjEBGYatUcbO4j1f9zT
Lw3KePuwQF4UA3C/rvsMh+qOKbZ7NPYDLPS0qt9fRWxx7sOfMdrOCX+0RmkrA8eF
vzKyzh9KICMu6oRBf5L63xPzwKofPomzNGow4dHVcuWIfB/IwX1t472OFAkDJ1Ka
Qpl5uboZRmCrO0R1J5/ZtdinUhbjSOVlfHrkPIHLV5xzpdj6H96pgXVFcrTJs8kC
8SZNJeBbEzoRreAONfJFbiU0TIU8ODfPakh3nzNWiUHLko9ZqaHG+YJowoZNmkWX
Z8oCsD0+y6pzEukxaB9kBranK16RkWnv73jU6TA+hSTFCs3lwYML5STLko+xy8M5
NNSwKuAyddhM0FebsJOF0IwRYoDumZZb+YmwYG4e7K9AYi3DKhm2gEBHeWsEF+rW
0ewc1HLS6TopvlAmAAMgnmnYXGEildmXjH/wgOWKs6gMmShN9sNfaZGPJipHyfac
vvRvbRJ4Q8UcMtkPbXiBUn5vVtJrhu1eIn0KAZPQFNNH+3mg/wF3+0cDzKxx7Xgt
7brfgPUbMHY/lsjHa5P4gaXYjteQRSD3RciyPgCdcIE0hGY6MtQXhpf52Y/hk/gj
lrsyPiy/Kbn3liMFNUgb/q9acRCrlPPzkCSM4Be1kBXvuGjQKzsNcdxIraEEdkSR
Q2WYby/yYMAEzwLuLVM0xRU2mPphdFSRYWcs/E0nBDktKXGsEXY8Q/IwsuVYiJIX
n1NoE16iD5O3Oh6SVKt/vALo4Fwm+u8JHEhJbEOIcFUHT5bXYQZg7NfmrRjCS3D/
ZvCyrVWVFrs4Edd/Z97yH1se2xEcPj7m0TZ/8Gau6BxG8vU8GzTFNiRcA5MemnJY
nQDeksGTSd1z+8/6BPjpXfvp9+es+kdpP1116l+RkGzIjQ7scOExy7oyu/aJ31Hi
N7Z8MKOn1P5ToeG/4zF6A+4CLELkgPRKSRDLFmCEmO1eRL2N00J6GB+HXYHPIY/U
PhztrnsnFeCfq5tisl4seVtMpdLT9h6DxoR5vbd4d/xhGuvcOczlnefzsBu/wsGL
oPOuF88ETz2Gi8wovJch9lBLhe8jqNbJ3hsbPmvUTBQ57R6H4rmItwQeHuyaoCF6
j4Q23xP/0wPGjZyxQwgemse9C5J++alPJTn+YvmaYJMhqhK68GxoRR+McTy4rLvK
/lDc85hMB/DQjbtBzfqXIgKdSfU14S6DQ33SpnG2iS7/NKijsJYu2hH3E7SSw01o
/9q6+v2eJP5Z915B9tBm94W0A8BMpy8cdLhr4jxdyjyxrL7UusspGulIEmPbWMHu
NXSP3jGO1DkbCxvRo+zbEzOUR58+KxuRxL3r1TMga5mrqaeHS9ARc2b3Vthe1do8
KHpbAjIhhaaRsUGT89zbTuAU6ZgzXKN+MuojwnI63AG+UpUVtHvs9jMj3jEX8Rx1
+TGecRpb6DQSafKz7uM8cncEYWOrahpcrtPbTsE43Z+eiupiBscniikasEF9IDXx
FUjFZX4udqP1GC7mt2ZoyV/Ee+ZQZp0LiC2omuqvF/EFdpLL2laAX4Ws7KT/5XsR
gKvSo+HPCjF8FfJJ+/W8qzgV0YCgEk7vAwWUX6m3hMB5/fF7jB8ZH3BBb43KD+Xb
Zgk0h8SLXuBK+9vh39CI2QRNtprVpb6xLmYsi8/3bR/6vuG4SwWfXa2LEtf4R6hd
Uewd8nlsHg3jNkgjrg7EM7tFaIbcbwB0XYPyHuASDGhnRKnq90gcqLCR9Q/Mxel9
GvDh4Rz2eS+ZTctcgmu4xlQXNpJaP9OhcaMRb8PzWuEQSXwsMAyLRLDCXAT+N1xl
yEvlbXbxcopGRJUfV+qo6CIwKmBkzKbOIDy8i7p1hGbJNQ+Fcp0pJrq9H/dgLnXH
gvSKkfarE5LWRC7/Duhmf3nvgxiYzSJjNNtelpgvAm16F/eoc81s7yfy5H0CMhNP
Qd5eI6A69plJahLv6DgZ+vK86WQqBW3IKsFVWVcMQQSOtpqLDFaEHQHGVjhYBk23
QvNmy8mkLL4+LQP+cWl/PGyAikN1z3tkSgcBNbN4ZZc1aGlVHAR0HJtcqTc0X4Qe
4ixHFUE5KkJgIqqXGqHONS9PhNiKdZeOX/CMfPUC74Vn3N9DOZLKVz4rlH1fafmc
PZKOBGgPxq9Sj9N//a2ByMsdA8TzRXj9PhVI/2Yt0sXpVx0JoecgC0WKtszcyRUy
81iwFbj9010fTOPtGrOoOJJef+RQ5OnJcNNc+ZjOCG1uHMtSCiJDK2oZdYc+q50A
EMXlaRvC8w7abKBTvVX/jF+AN8wTV+IamOgX4s7bMgi4vnlw1OKs83BbQ4hNB29N
dJ2LOUJU4ucFcfK8DJaIV/llFLP4wWXQG++kTwp4j4Aqx6NgSpjfk/vuvTZgDcoU
HaRVbtqW7/00ophBaR4M3i72UFCz7aZi7NFQ/YE4lOOziM2XLb2xIMEZNOZGwAEl
Gbj3EtAAC+dX1r747XkwffeEESQZoNG7lKD2IEFFoQChB2jJexUnFjC2d8IUOomg
RBHvQoNhsB/B9WK/98T/IU6USisBcj18RB+b5jw9vT14EtRL/0KkwmNFGDmFxQXr
pTpPdCEnkl3f+38c9QeGdvwrQCUU1hf7Oq24mJLzYZcqlwlbhErxr07GaTS23B3r
MzUw9EiNP+B9xNzTBSSXgP+8z00t5B8wkHOP1s482r5FNwYzinCQcZsklIA347pg
fL8tUpJNRod5fgfx+KvDiDztNQs4ZqIKZ6Z/t33RaBBa6pozic3Z2k23jqarlZBZ
DTvPa1rrpkX2c1JNTHzJHt0svVhnjGuiWZ8i+p19MVHJ78Qp6fQTZp/wHjKbKcbB
28f9NQr8wIzP5efdIrzXWkbS+lXYzesmTuu724NQiRYo6iJqERqadI3VcJuQj/Fr
PJj+Gk5Fo7u1QXk395Y29pUfBt8TM33nVVXrbNBafQv0uyayGiYc2H7NmlMpgHSf
7Xl6gTGhvw98dVfZG+YxHPpV48NtYB5qoIYtpPeoo8tZlwzK2Auio53xTPNy+vPX
Pga5jQ4L6BR+ave74+IZu/jSlvV1ter9hACi3TU4wJUc/9Z/3lDaavTknzehA1Ks
R7fMOfBAW2lGB6mRFp6ciSvGlv2Aq1UZY+xVnG3Aw0CoI6EGNqGn8E2Audq2dG82
ZtC2kPbgl7wtr05fgwPb5A2E6WtBTmDHB4WBRn3OsAhQYcIi36cZ+QZsmkcmhhfU
uRA1tEix2wIKHgzDVQhovqrKF+QcyFuz22LltQviM9H43RbC+ejsQ0PTVzJ066nW
d/Mk5h/HZROwXn+O1I5RmpdliPYDiv6WAwpl7objCMwEauu0E7UxjCT4bf7CYtKb
IV9jRGMOqK/WWayBKZkFa86mGwzJTaUbONzm71VlxCEErRve/QHwovX7CL17nV5E
wVJnOn75o899D9lLOuEXJbV2Qis3UKg+hz1DjurOvrCUdjXcpXfVWE+R5aPVH7E3
TG65oP/G0xLixKiaL0vlx8N3I7c32LGv8UritdEuMQgDic55MAZK83FMiwNGajRH
0zLF0ukEyFEWXOE++dOce0NzbIW05cPJeod1hlVrvzPx9kzTuEeyvGdN+0JOpk2B
bELtcc6Iy1pjCA62uRjlOCxhdI4DHA1Uglst5AMTprVClZkQjzfwstSo3nFGVYV/
hylTn87cn5xeIbpjjKgvDPgEIushkF3clZ2t/l1t+6HMfsuj6ZcJ3RABj5WZ2NMu
SDnwXTnSHiz5WFiPNd6n+xiiEeFgVQhNiSr7L/tv3772pNl8BTxypVkH0dNIwFVD
G0eKRSsveICqoZgSY0VN/Nlh9bm1AolRRQyQCCqfV9utspyHd+M6528rOtg67pof
ACn21eS5Sqkl+KHv4cjILjywvBP/bpi6nb2+llzMef3cqjkglgS3MH3wumgmWrL3
uk1GEh1Iw6mlaLjiAtK/+FJ7CaLA0yB/Qi55vFAmkzD0cv/hiKZrjqgzY3nPpT4N
Gw9caZGT4a8KRr9CwQzp/sU2o4h4y9QItA8TeEeIzvE1aYFR0DCphLxjnY5EuR66
Cah6tlZpukZudV/Ip0Aq8M89fPRItroDb7LjTATzrrB+g2QxPgNl4KhOOfEE/yo/
BOg0C7aLcynZd2aNDFyt8zHdaSWdpK9YUVogvCsmhfEBrKX9GjNexvMaAtrcY01g
EUkBpz+9PSsqiijJ7OPFPg87/EWwzSMmuvxMANPLvBbEX4XXAPfIUD7UkPL8vud8
0BGv3NdFHR40BuWm3rYWv9yklBTZTgXhuEw905QFGW9HmxF6TUc3VRwHS8UhpL8d
E6RDNhDPuga+Orap0tqapP3vfP4y44tb5Zgbfq/mbkhwkmi8H10y4GSnJeF2SmDe
F8EqZT+WfqzSy4I5zTxq0zk8Pj9Uex24J32aZiinpN5p3OugmQMujf9BdNCD3jJn
sy5JOXQv9PEG+XMFb4NhrX2d4L9IUsrFtjvJmatrpu/8dWB10TnkMCSqc21HCxkN
`protect END_PROTECTED
