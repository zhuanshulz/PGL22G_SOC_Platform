`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R03S+pwNovYr+DHa5W8ax/p6AZlh+mVbZr/HDbeUcA91Sz3QGtF6QMPBLxxb8881
GWF7/BMtndpAzse7ldLRORiBykkWcXlKuuBpgkdrl3EyOKp1qxpzHBKW5jkMYxy/
K/W2cr9CtwOLAJeEMfWlMJbg63P1+1aBl4VfiLoRBzBYEJsnX60D8Aj9yehzB4zQ
PG61UV1GjbNbKVK28TYbFw04p4v/N3j2w/Psz3/thxWSCq3t5GI8Fod3R5DIKgpg
qFymg2GLkJ5TJUPjrnV0eUNmE3/ItVAzFQ3AmeqYMtvRhiZMlEY0ff7aBA7SDvvw
JjqzpG/qCNxaEzP3Y3ADpDIf16lVBC+vlWgbaNfj1CnyeJmB2TaPSe3ymDpSgngA
0oGPY41XNIqVlZBQVd8ltmANwYq0BBXMSgiwDUB/7cnosfpVRyOufvITXU5P7EQ5
xkZCC9OKxRrZz25XgzX9e3pjEfMBRP3OT6ArK6uZjfeoVsQO0XrnJtk63p0YuXp8
qQoP4PmpIXmxkFqhMHF3q8zrZkybrsQE9MyBNCuy7/gr3afB1GGAH5Z0g3lR7CgV
83GBp8m8vtII1Tz5vRAD5nuoVKKx2K3yNhDX03y0g7OqxKsxY7xjbEvIpFTlZ6Tu
T7a7iBpvK7MojcHt6QycPdt4tLsNixj7FqmuzvYgPtgB5Hu2P49AhKd+0NAi6aC0
Wu/+sgfk/PDGjJv8ejQ7DJx+pi4jdDvPfjfVPQb4dOJLu1UinZAT5mxOzAiV4Mnh
XXSfaEbbONWHXtnWiKPj3OxZNUvZE5THGpHWSA6aAXOzJcw9EF7Nzqd6+JegM8YA
+gnhpAJOJWFbeR6Hr7iaCnNkvM0mfCPYcycQ8n4rlzs6FZspaktIyqrYD3YriomW
TPJDy425QZd6FuV5IRi8wrqq4n0PPzyEmsXGFJ2HnA4FoMOp2YyANjORWLc7YbTO
i588UfrjcQ4zPTn2ToVMtPDVPdPQ54wMt1J1YSEC1HKnAcH954AGcovuJyb5O/sl
KzepGP6Z153Kt+Hnhvph3l4p2e9XOUVdpb4Jvp/r+GXtpxGI8+ejjCz5rLlYA7Xo
xlH6yi+a5yZwWsDhynWbFwShRSWNRep9/5n41bp0KduDiqyRWD/lzG+umu7x/XtG
jQpY0SkQqbidLg3hEwItM93OK7mmHdy2fVcXQx/wSNHZ+AXV298bHO9ZgnetHE9f
Sdsj4ODz4AC5grIz7d8ZWlYeNm3gYiRMtqcMgWwsCmVxwOOoPD4DC3iZw5Cra8RA
EZxsU365SqSBBbaHIzr2LOEbNAD/MHeP5H6vI7v2YH+RcoSBb6jxdr+FvJ5XLAh9
2u0HgJcuraeUedsnKj8J6f+aSExUb5Uh1/Ki7MLi/FC8M7oQCA5D4kmNzKAJRGCs
vlu44VLYOdqlbQZC1ynZXEcxLDINTpFPiw2f7/V9QGE4iPtBlYH63xiQQLv0MfLJ
r+fbHhFntzMqKWaOZ7DSWSQiqAB742NhS1ZT1BiJkVEZEEm78YDDIMHSIK2xaIo0
x4CJcc9hbXcIKWYDAF6wseAHvw7pqr6Tsm2FPzYT4vJ3rUwqDxqx2NMZKk5ffYw/
aooa7nwe1t9WNVSP6+vKY0orTEtQH5LKSWLzf0KZSkfmIRV3dz90ymi7JFj/Rth0
mIoomjEqsNEFYgow41z9BGbC0c+LR9yUT2pCAFja7WgIQ26OJ1tHFngJwznkfdtO
lpVO6OEr3Iugn4IoqTV7iMeBikU9gjpTlf94/a9KT7iI0iwbMxEhn5x6QtiF8oLD
mwGYuRlMlOyJcYV22GvBmiymG/af54A4RybTxlwpUbpgUAYdSBMR2liETViQtYYJ
g0p7OuyMtOKQZaqy6YQ0B3X7kWdpBpTqgutf7wpkN7272bxLsdM3K5VxpM/0852z
SZJjHzE7BS/gqfzR6qu7VwM+2GGV9QBuWDbmOUTTLuEkKlVsUILQI8yIr0lV26EW
tPDPJs+yDieJlx7ed+wugJLy4iIaVbL5wMrztHRSBuZO7ruAIeHdryb3E6xfiVq+
y6+Ms00YM0MTTLIC34dCO65hpGtJ8dz4ZcnU18ZKR0e01Znwi28EZDzmQmp2tff3
AIAFdaorVV0BDuAlyplFmfxb5kNCzV/Y3YuYemVO8Q2x6vrTd13eC3wT5rO5IZFx
y5AC9f5hcO0PC9aJZY2SAbro2x1yj0p+VhTuzDAo4Oxlo8QfqNhy/IRdRGVr1qxm
mqUZvO+zW/7zF1W5ko2j+XGgK99YDQI1RBalovJC/jxT/kRCncmU7dGHPBv32uuG
f/CcaUxNFCK4xp2AZXndplXT2spKOMluS4LuzQDacBoZOSSKTdCYfGK5dC7uHl04
EI6JnnHSo/ioOym0n/ECNT6IfruWYca94EVxJRKlLRlIyn7fLfvY0Fs8z/CfM0iw
lgKcgJPqmutLGRUnYYzTxRqUaKm5c2y9NI/K2vkTMbFot4QzCbbvLwClhwGHsSrB
FHmFWaBnrI/eiJBf++uLGH3+YVAhPXxuXtKRcmAvvCHeFI9J4sJckZR3lHAZAPIz
6U+kdBtsQpOiVwFMfK6sdhfJBe1Ht0SakPnfnLIsZJsMIQKGKQiEiaCm/Au+GSZm
pRS2pe0ZnUu3DXHuq26E2A==
`protect END_PROTECTED
