`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
coJMTjinZWMSgJfAKTW6lpn1bdrsOH0ay80t/5PcHB6a6Skaqk1xjAftRvmdNgfu
z04B81SJrS9JGvG0vp+6xSQgZT6MZkaCXvZp7a7HNH61Nw0WbVyo+d72abyGQZiL
LsPrOecMSghGbzS1NE+zJQ7DpQhnHfMRIQhf1agsAhVp0iofKeBlkgAhyGfqYlRt
cc9ga39tmw59+PWjjjTIM2dEUE+bp7DZZ9IhvYG3efEGw5+VUrSJu09DJfjJFfix
esgEmZdLsUPXXfD1YRkSzh2e6JwG28h4vruFdjUptLWlu0C8CXhfTyoYrrVc3A/T
e8+fiRPhHtHTY6xpB8PEpOgVNaMqz3tHzG6JZAVjMVJ0fmTFvCFkblrUjl/540KZ
sxLP1NgQKcR7QbgR4Lmw2fITjgnA6bWIG6/KaQpma2VeWeSU6ZZDiwO9EgGToF4w
vd0GBxBZOn5fXV+BzQPakkqxi9S2tf5XJjYTlX1+YTWEiRqSbOKJ8YdTZctX3GyM
wRobGX11973ZMtbqAa1Gyw==
`protect END_PROTECTED
