`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KX5B8XTp5FoTNdST17cEFhYS1fwtER/Y/jIamkk8h07sLZtVVJ2gksEbgDNbdHmq
Lm0mcwfKFYqcRfnsrL/O5LyD7G9qKU65U39+8IeIi5e03VnEh2fy5rAsrQa51jXT
l7Ul2a9E2WN6sDUIvssCebE6fRfDUEajoufRVMTfMflvsaMUaEWrz9C+/MCNQLwZ
H5WuSJNrVfUHrqjUCUSAYvXATx/SAcu0f0RzoSDs0bF9KerGpSIm5EirIhFkhTaS
f+abPKEOIIteCMIJntDaMJW0GqPAQx4ugaU4SVKAltzSRnnT8tgKokeiyqnbzc5D
HO6IhWlSfZVdj3hy2jdap/dDBDCRQImBzlvD3xfEF0hnSlM4Gnj4eHXdWfvLpIjm
+F1DGiEYBbjnqP9998B0lbsNXC8IDMf3wHwPOLuH/LU=
`protect END_PROTECTED
