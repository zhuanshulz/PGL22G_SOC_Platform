`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
55hU3iTrIkW+kukCo1FtQBFKZ+T3PBJN+jLAjpkJ7O0q5Vs6Gols2bzEjfyn5VJ/
DgV6t8epHLk4UrNSpKkXyxl5UtCq41E5f6eNHuMo1TqLeR4GKF8SgS8YvUQ2PSl3
HhrVdjjO7HiM6eD8/fsCqabhyWkMnMfCOTfWN9SkP0qHAWVQXiFJWgZL2q8PjUBx
LLCUx93e2A7t2yQ8G/WfJadOSmPsa7tBnA9ypUz/h1ZhYaeAtPQQdCQo9kYq5+Fl
/OifR4Q5YgHaEY1hkVuX3Kn/uZUmLDZEUg4ZTN0jOdtYI6pUbh7w2s7rlmVdDvij
zYkYv3S/teJXOt2szzJTgO2DVsHT356SjIM5e+qrdnqYtcIglAAG919IdVEq5vVK
D7c8DBSL9bdRvJ8Ma6/qrlT0e9cbZKRBuykMLfTxETHPAbksqi18VZO0p91PMCBU
o4hsaD2uUdSeh9up9NQbxjFM6WXYBwD/oekQbInXdaOhX2rsMjMqR+vp+FpVK3tj
mGQ9pfyY4WY9q5IAI5cf0Q6JrJz3dUBI9d3DaSc6tj7P62Dn1tti1i+JzOHaCXlD
tkKa3V5mp6AwlHUJD1i1Rf1nQtCP+k/He6l4rOjBRShct6Eyvryk54mBrZcJTtye
S5PUy0+Oq79vRV5smZXhUCKw50J9Kc90uxiKXDS5Dde49yFlmntgxs+STzVvumrA
n/3e3u7nvGaxiFeuLybDwTWsrb1pHm0BfD0oFB66n4FoSgWsJeHkti2pasnGagha
2NXvpdqnXO/r28JMoI3lTbG2zlGo4sfmCHFqWUORyHeusgP5PHM4D/YkJSZTP/SP
Cfz/dBC1Xjfo0IarAA0dJhzryRQLNdrljdxgGHJfKb+mOBv/BBduR/51YyjFDJYB
jwhurR1fYecQ3pD7E02yxk7b2YYadXWDmUezY2ovlcmnnGQaiV+ZHBMfgqsVj2vg
yj1+VH5obyXBiaW1GX8kAhlB+CZ/yOz1YTUbMBicS0j928eg8Gu1WBVhpxJuJ9Gm
ZN9WK04+Wc2KY41o89/DlkdOnUWmaWk7zuiyaPZDt4J/5IzQog4ohlZLA69sHlcQ
THPbSviuCk14+OOMgbDgPrMRjJlD0CB91jGNhWm5e5pazoXOlQOiLA+JbnCsdAcR
yh9HzQCkQ17ucCpbutYxgLc73VYT3oTKZWDuh4QCQ+zDrgvAyvNqZMQFbfreMtgE
P8iWtCYyXm5wQlLNbFmWLMhFQcXigysSGI6JHpFlwJaO3jlYXwf7NUNPb6oMpg8f
NOCjHADjoRTIpfsT7BbmRV2UooXNcXhVPvsAHOjxiY/EV3IPwD/XxsJHMFVrg255
D5LL5x51NCxg0Dw4cAHKJHasPO1AKs6Ca25XxaUYvvkEXJH3YzGxNO2I39lm0TbM
SL0mlOjT6BsB+/V+J+H2PUE3nP+rdJoF+bz2k2npVDI=
`protect END_PROTECTED
