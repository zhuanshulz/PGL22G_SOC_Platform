`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E3eYY2CWURHi+94/UwH4Jilgf9HNDXLBD36WuDwWDE+vgqCs1j6ik+ZoqkTe6Qnv
QQjdYgdyn1gbx6k3YSOuUyRMdkaKoXEJqlhNk80YCUzzSwNxprV4hzR2E7o0HQs4
GAPELQ+qNTkaoTEwpkbBUz6LJk+fuStXdZ9bRda2x8YwnxGtAibqc/H7JXtaDM2Z
zeWO3C7bJn2wTjYvovRTrDonyKajV49KwpK/mRuaeQUf8aBGJJYFOeAyzpADZj4O
0Xr5/tEoO2eioGe0y8GIjq+XFL9DfJQccpZzqqjy+dP/gAV8+0hBEfMo08zHmF3Y
7VAQAG8/D1wWM477oc1y1zbD1EcOlzcNjZE74qScClk2dkQQZ4n1peliZJJvjssa
nlwVHrA080/23lxLEw4AgoXd7/NdLQBL84f5sWPeFhY5NvMEuDkhJq1OuzN+CIAA
929/LDDlkePeluPTmnUrwdNaOrWLjRpllInvDjm9/QpjsU4aljo0hpPNv60LDUl1
G30sTMJ+dUjj1ihapne/hx05YJFmxlbz0FgsYsnDFXxP/OmJ/zAbwe+cZHhCIdNA
eo+65UXAnL3h+bzitNiGTsmJw2EBUT/0y5qTKdpsaOnSIEPgDusSl1tCmeWdG+N1
`protect END_PROTECTED
