`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r6nsV3QHk4WtVezwkhpjKP72HLuvSsSNyGYOHEslQK3HNPY1mjLvxus/pqC1CmT+
a1A18c4g3kJJze3fWqRzk0sXCVZG5dskz+taTYogH2FlSxylVnuetVGg+x5dGKeR
AndR9lpsE5DpHjdkxEHEpgMwgY59Fwsgv4i2+nbRf/nlE7UR+vhhw4dq4T5Vq0ma
LlSOsTUgXrfde7/l7jg4uED0prbM8mj9CulW86wRlC0NyOCRmZCwPR8rprMsnWtm
e02JmG5Mql0b0FlLagzzwgwdbqNlkxJyZONe+7vFoLRocnrto1isuQW+jeEmQ4W/
n2FAY0lbvVnW+uiq/fSdXjZnWzgMTdNpjW5V39ykChLtHdjl2HRWisWbJ3QawfnB
ClbVNp6wkH7hN4v4H4mVsHMwKfkjuiNcZqWn8WgQMLCv+I1SaKqDYbSojghpYFnT
2HRwgABXylijeh2q65nK9kPogOS0cN33Ci4zejCHyN5WJqyDmgalc3sqJsDztxeW
/NjHUKjz/MmfPX29aDa68ynTS01n+TwA0FeI/Ct0MdBEOUB6ejpTkqapYIGdkv25
UIsFflFpVbYxI80oXVt4OVxhpGdcsEdN1P09ReBq4p6U9xHwKwwtifXqrjvcTG5f
GIqaLNPrYlxI+FeUOhGSfnqc/hflUqUW8uuG4K89yhVKdbPyaPmRPERybzBHpfTt
PLAN6Zve2YV7Y6OT8PK9P/bmHv1d2HOsP9jDI3LvLymAoeJ6KFSVEgutsyesQujh
O425eE029Q8qDpjPBWRkbg==
`protect END_PROTECTED
