`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bwZELzMaHKuqFbEG6masIfey4A1ae7WRskbv1DPM5mMMgGMKA079SlFcYGeWideh
fgqRaYuKZEfZvqrFzxZKIf9rNY/QIjCiJIHc/cYX7rKBaW+uWxNaZcnb/ojjpTEP
zyeJ8m+gjxKAokq0q1jHAm3g1xwRgZtyzCsDFjsssljihIsvJIiIgpjD6PUfBDMt
MlcEYD+vWkMCfO4N4eHMVSrFfMUXWrNkho+WI8D+AsTaR9x7I1kEs1SyQKrzX7cr
fF/frGRJatEzqInq8lKXvPHW2LcVCsP9Hlnbs+Sv6jF5WtV+22uLgD2ftRGEt+Gl
tvJQ+j7tJhWUdEVzbtpQve6wOmEKsVr7OGR/anpzpS6XlEblTisCo2Ppk3MOkzRN
x+0nUQDMc5j96sDlep6PhkdIZzFU5WFDuG8vvIaJFEcj9Pq+KCceLHSjPpTVgcUP
R9SfE8tKeLHnYkI5kuJ1Bnv5U3tAzDULqzaJHjDbVgjq1j3w0pmKsBZ7hslbvNiO
5QXZbLo4uXvIqp/F6R7B93mMvxTOHpVsxRpP1R3xae2fRGlVc1h8EjOd54jGKLbK
PpeECGWi2k3qP3XK64Gglg==
`protect END_PROTECTED
