`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OlU/yY3yGwzGNbCSpJ0sUNft2ljecug+tFeOhYU+SlmfNVlxyXiDh4rS/X8XM/yJ
ATbFNSGjJ7gVDVTi69c+jCu3E0MUsCMMypydFzQRdQqP8huK5linvYVXCgPhOKpy
JVZ85N9DyzjWP4e4/R/NlGJl4FRuc6UD5jl07zSOn50g6CYh5oJdabGiixmssx6W
2FicQvwhm1q9iaBYCtusecW/4LY9Z5pI3FGuHcNScDoj8JipWrRQBUVkBlwuaGqv
MUhUdRmgI0eU8QJNhaucTPjePLyGqCUx25AAjg8Itsf9yhJihZsLhpGqrRFe+LQZ
U0tEXDw/No8j3N26qt7JEcJxWdcwkrsOXzXh7MoWEByvLwhSGNW2CRC3k8tzn1Jn
xpKgWTIqiEHVyc1ZpXlzm4EJU9Ph7e4H4fWoqHiY+YzGDhSHNyV9AiusisAjD9X7
E802V5VnQnugXESMXnL0r97f1rDBvQs1C6oo1uSSx0Mv4koEqB+5nVguz7Ujcdes
T4jUY58WVkyrYbAYb1JJaxiEEaHHkUVTgPAjlPnCsKkotjdt9g5g4GvQ9nHzpBsr
l8e3pnKkBlGfgX1nHUbOXQ==
`protect END_PROTECTED
