`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qnHzc1o1OYB2Q6xhaI8sJm/8gXpy5LHT9PiTIiFzF7vX62T/o2MQgQE4aTYNkVUw
QC12onL+4nPG/phoR27huNS2G5fVKuZm9Vid4vQoAIBwfvqx62qP3aDqF35M+0pT
yFvKBJOJJ93tdkj+53oAHDRBqPypGakZrvdwE10EZx0j6Wi7g0j3VaLkewhtS72r
ab2yWQLyNUX6fvLn8y6DLF1rJzryzJiEZoeN7bH7LM0NvrHwceOGZ9BcZAuYtI7O
ez5BHXH4fsRDzGwvrrYeltiB5lGQ3n4+LopsPBLGZR0wnbKThCTT6sE/Z7a4i/Wd
UY/xPbWjAvcSMlK+pKvuajblKAek0IwPXOz6zlvafuNYH9zsC5tcGHd9382aUyJc
mjBZmqftU/z4lScBwUMBsyyyS53PKVEfpqP3vNXFnyOmlrsBWPViFx8r0XQEdmK9
e5t4j25PlY3p0ZcOA1sHLL5XW5m+D6e9mepcckwlK4XHUZhxDheBlYJKAXqpEBZI
j83JNrTlO4Ej/aEucIMI0rKGGAx/J2NhFxzqtwuzn6NbguHGUUzgEc5RFlt7U8gv
4Y6Ld+UWqjTZSpVNO4bV7Bx1ED+1Ft1p1WDCpaTlet37qksUffV9G1D5GEIXHJ7u
AO0a9cVxqRfvPPv2kXsp7GI78j8uB1dSwWlG4NlFu6xfaHq45GaVJbSTQLaechul
lLiUGMoZu16386syOEGNWEJd3c0CXf4hTB7EQIYdGSE5rkoHaO5Ozdgzh2bR8SAT
2SrRbK7dTJ2mRxlcyn7xY2vNBioG5TMtE3s+t7SSGYTc8jZVoJHK3Py26ER1nPrI
pazb0EWuNv+4S9GKBBCpI+56lOSFLICbS4uexqv05d2cgGcXDxIPEqFWN0fjvPkn
`protect END_PROTECTED
