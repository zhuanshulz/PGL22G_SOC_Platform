`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5JeQScl9tZf86xJy3tgEsrHyScyZrwSeIKy2f1TYBjZiUbkVNzSN1KWUMnlboahW
CLTYnaWvzxyTL6u5ghbPPKosQtESk7SulxFTfxJ81BzhQwtcMtha8c+vp7AWwczE
NkVX8GrFFjVwWQgO5flnHrIOzYKuaLi9cO0fn9yKsq/bfKZAl1qjPfXpw1uqJ2Uh
U426lytkp7dDJDKNV6KmNM7uQ4+BVD/IuXbIdP8Kqa+Y9IjqwmuT79B+CyQ9WKIX
6inpR+Fbpmv6G1DuU0CObTnd06KAmIU5QkIXmfOblfDmY0gBA615i8rSKzaF4vsG
V99Lk1gxcmSKgeUwtoPX7I6mQdJiiiZSTTjorD/kbCbO6WO8iBjFxz9xhOYHuqJ7
cGxQmdQyRnYEbGWZM0ymq3TW7+1ALEh6IwMVD57ErwKkyVB5HfyRM4joKTIpG10p
Svr1llzo1YHpzFX0TgR4ZSLJF2Us80aKR9pjRaZ/d/g2vNtFiP32URsYvlC0TvT4
3SJ7McxExYjsSejwz2vRdTIKL+ZBOPm1kSXGAh8T1y2UY5JVSkgyhf6gMUxvsfeW
aXgRSvsT3byc/GbC8Zo67A==
`protect END_PROTECTED
