`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NSMUMHbD+6PbAtHCYqEgl1IklS98ts/hWX0ceiZ7dkDn8+f8qo+z6+ATSci7xEol
hVw/u6zy23KhBZAd3gfi9SKeBhBbLXzUmKv/+EdDfTYGAPGZvFblr5sbYCSXPseY
LVXX1HtPFUIIsdS3mzFOdnzuNnUdpPiThVIW6FshX8uGiduKQcZXzE6ZK+LxSSjD
fZt0IW8yo9CFmcZLwUe6mzDwTk4enDDVfODevIDos95H2Q8SahcAxnJfWH9Nj0Tu
FxhLVBpebnZuhfgJckLwUL/DY76ze6tBNhaDn4aenFnGXXSoioRisq7yromoEpeo
PPX/08+aD5qP9X8zEZBsaCYT//5BlUWHa0m4xo7eUOhfw6fgj3e5fn5RTwW3CuBA
TdjshvZfpXh+Aae/ko3fI7/8SwE+H4heyfWm0OCUDb3uAIOgZmgr3MorYdS8Z+46
EQ3eaBykFAHXlwJRfqOkAfr25Q7Q2rtZKc4mMNtAnCAGuuO6UhJwrnvqIrpC3VqK
DM+pR11c0j1V1We2esTs9UhUyDggZVDNTaQUkEdgO3HSrZaQI8v5QsZH9yvk45dK
qXqlany3EJPMWXVEfKOqPoJy+dNYbaXJX7dRor+mK2Y=
`protect END_PROTECTED
