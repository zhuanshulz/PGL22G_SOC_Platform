`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F5SBZSBaIGI3BLrtzPi7V5eyR6TsYTMA6a5VngbdZ246/OabmHroHClgPZSpEnOU
udVPp4z/A5uH0dmiREPN0owdmJvTZ1BYc1mW18+03yw5ILZbDqRgDWdT98CuSBax
/PgvvYi3pk/C+yMjyS/98Case54ibT6YrvpFkWOTrux5CMF9178eygpwQM5nvYmx
U6ajgVc5zL9xPfZnFu8WNUi+R97g42IQHvSEDCe4BM1wF0timCP3pIJLqV4obaTR
H3gN+Vrxv5KXDhG7hPb9l4bA5iHimTR46e4zcyop1B18bqND7rZJBLm4Ool4GLX4
prhAVnnJm8DrbJothqizBrf4HDqPVJugT1JnVkfxVGxAkzlZ9xh7/XR7CLUzTN+R
lbhQSyXs7WwhgYe4+mQny77twy/0BKxKvEPXznj4gPf4A/uvEIzsgWkilfEsYebr
GC5TJAUQfAQisbviQi7sM6ccjHI4cRVPOxmCUVk+ImpS84OnwZxjg7TXRV3mKJAh
QnApyh7FQWWFI78YJ8ZOnh/L9MADIrilUyReDNN7e7LEdzyFu3xifPUvff4zNYzV
`protect END_PROTECTED
