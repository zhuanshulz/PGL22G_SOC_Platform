`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KQwl5LquxyUpYuYa+55/UEspFlKbYYmmZeVZxW4s4MWnnZv/GldeY5Yn9jCQUf0h
6n1vz2zbDc/Oysb8K4r6SxpmwgNj8HCSGwoBnDR2ytRvnI/d8m8OAlsJY+ooDakw
QsQoICNA4sTV19VCNjvGmiZen17AbOjMC5K7tcCu1lvbRiRitrvhAEabvFG0AjvG
fFrQwI80YtyLho3ttFOdrRSWoR5Sd8wt32qdig+wqqQvBocKxrnOtKSi1CuP2XUm
fqL5Ftjh38spdajD2wgDUFbcEqWt9VzT+l7YwDc81Vye8bZ/0cxh5aaylSEh0Ryx
Py2SF6ETzQOBgsszaBHVdBY62Zjn4IdUlP84kT9m5zYGRJ13zadvhFRbEXFIkxji
qlWeSGM3iS5VRxwugKJggwr/oPbgQDDwROBpcJ8VsuNwxsyZB+Imfz5c3PCOwy01
bN4htXRaX4Andu+KrARjzw==
`protect END_PROTECTED
