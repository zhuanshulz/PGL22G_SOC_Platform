`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8ygByB85e8KYPqTBI44h8KbsN0P9WUEn9HYgjm12aqyCCM/ib5LsAkkeElXakwo0
oBU0CMjKVCdpO9tBn+82S7bhYyTG0bfjuJZD/OXT9mEdRxAgXWOdsajXt7S4HwLW
3cXSZKjZVVKql6tuA2nmU3HS38LM49AmyHjYSwSddpYpgzk6ogECqWZcuytp+yBa
UfKjWqVBscdcljohVeTp1EFwPOkcVcHEOrmXnQVG7ScvLvLdRwT6pI9bs4QOjo29
j143e0m3fHDTcKzJu7iazR1PrYdt4eTXwWp2hRbb5/cOfU3xhAZQ8kklsjaPOaDJ
H0hL44hQ5fx7YwOrA1zvH1E5vxTdGpWhT8pFyaWAnyWkMeWSTZqYnF3dXiXGbKFX
WXw83zhtk2UL1j/34L09qys41JW3svrpX/Apdl9E1MLEHz9sx9qy1YIqa5YmU58M
g41Ubb3QedJdFj6zZs/cMglbnl/mOLq0k6hib1AW4Dz6JfPVOeYnCNFXmwAormv0
s3Shn5xWfJBfN1eVS2ED+Rp6UzIcHiPA3fha5umRUDo/idXe/gYHNHTVUlskl3Lb
I2iaJkhciKY4J/44rQHYZrlTuP5p1ZE8SV6pVgu8/9G7HtYUVEpoDXoJzU0hts4T
`protect END_PROTECTED
