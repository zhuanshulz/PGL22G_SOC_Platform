`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ytho6FlpCTXQQ+hoLwHY6nyyrrvmI88vzkj31u8/X4P+sECqyuxDJFA2X2ypNeeF
aouImnCuN9qh8+DhKGFMNsTf5ymUi1eZJLwU5+zXdNrDodtOhumugZi6KBx06q1m
/7cAJq2yJ1SMO3CYQkNGD6sSkDwHn1+Qri25dz9/6XvyFFUq2SyQTkXp4aQ5voqK
zuSV/oXYuQfsRwQkIYVC8XT3SKudxvSQjgsvK3v+WEk/ULRxNwrNuP8QCnFr7frm
FE3L/gZw9F3ju87q0evi/60vAO9RftcH1ZO+DsrgmERGlwKkfT0quFNY0H59pvsZ
9lYQNdGFRU5fKp+rbUCnK6SpLE1ahdtc2TkH7Uolj/JPoI6WEouf8UBLq58bZAMq
6u9Q568PaE4F4iFX1iBk49NcvO1BKVdk+SFVUSFChepET01SfE6ODmJUp9s/EH54
RfsbL448nGXYREXkxFbgK1Mc7bgshln7fcJ2AfqWHppWVYaCb+9obn/bu1c5WItr
`protect END_PROTECTED
