`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ycXBMOdW/qkVrB4VnB7EupoZNhBUG5IK5lmo48O43GkiFNfBke1k5x57+9EkIeoZ
vJSICrGl4lCB27VldLERggbrtLZU5SkXqPQKQV3DxV3RQkrPh/2IHF0E5jm27d85
frWcSLmNI2NdsX3VWOl/wfWqQOeijlHtdqc52oVAKaRj/N9OcsGw+XwJ0VQDVDch
z2bMz5CC7+6CvUAJUdJRgchqaU4yHSwaoG8XiolHVbFBGjktmY+xaktYDMvfKOq+
wvuV0QizgmauUcTLHfIg+juQdqdHPduRFfbfWRcIefqgLCeuAHWjG4h8GBpvzXdB
SPfSfA4JzQcY6B9+tftWVIYCRvzbJ/g7LX3w9YFAnLFICmhUXimPRktVw4cDSNVT
GldXBTnrTYTFu244nXvoFZK4ykGZkLahORS69qt0Ff2W0UMweq+BWqysXiuyWDq4
5AmWEb2vchWjOjJYh1XmhhVCfYICre9OF8ryF2e+yNvHIjqJBjN/4+4AJhY5MYhg
KNYmHRFv7jZzCMQsL3JcBz3kaRYHaKTRi60RoE+CzemjVNiLnFKRV4VXW6NBdLuK
MUDpTlxI8gi1RTMSkjuVNuip55NyY7gyVWqbiU4SaOxEMbuv6qdpDAycERqmiN7b
4i3TPk5wRZPD7PppQF71s3BmGstEn76wiXV+d0+1SPy0Vw8bbUvHifl8Hru5avk/
8+UdxZex+Lf3J8A4Gqel6UHljke5PQMi2TMZSEJXD5pVje+EoDJVw8/uak6NrKJk
R1/6ledIu4bPlGgiYKzzPpuoV41Tt9aMAgxY5vBGefJP4/eSD7LeV5Mb/pcjK1N6
wRnS2DcLbdXsZlUCvtD8XQ==
`protect END_PROTECTED
