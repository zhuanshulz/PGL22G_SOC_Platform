`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7V2odYH714gfRQC/V6Yqve12izVm1bU3n6wdb4tPtac0arpfHe0f2XOfd8ZWjni3
ZhVKz3IB6Ok4oFjLThJ0nIgG194zAf9BXBMnDwp3YwNxODVG/e42BdAH8fUM0H5W
QMAX5KrPaUYfNWnAOJmqJICmJ/B61j9fIStcj7RtB7Z23M+CIUYs2TLAsG0diMu2
l/Bbz38Rc/ouRBI5Vzjop+QqEmOaUtsSxCmix6En3Gv4KzwHt6XYLMyWOpFzUS/P
2G9xanYGT/mjvWhCoXymDFGYWu+baA8lzrt5O0TXi+a6ru6g594/h1kQ4QWwURn0
dmCAC1TQxUbC0VEGwQ++tTOg3SXRtdUVDrkhCUMrMeU5VmWdHltpjnbO3rBZk5uL
7eKEL7+rJ4mi0rJBIHvEQmCtkKKHFb82mixL2ZgoZD8ZpvZnkk865EfQYYfZAASF
zUxUvPrcPCFgnBJ+njd6tvyeVWjH+mQq5LMkCSJ6vJdy4Tg9FtqPbg0kc8dofNTg
MyzIdLdgGO2J+QSVfSSI1z7q0Od1m1y6bic9WvBdKrTxrHuB5WOQv9hFbWL/8h+K
MERD8btiOFlOpbBPtWGXt9TLfTe85fahw/JHaaOOa/k4R1ld+6+J5pXfxCWOxfdw
KhjyeljJ8dtykkn5hnSJ/9NB+rBok3NaDx56pbVUQm+cNBEJlcSg1dqToNPYvK4y
K+R/+d6qpzCcf67ZnTyQbzpPeKSEEZMi+StPdaeRlYfBWXpMX+cC9qnK9yvbmegS
WyWfT4jaa2A0XM+bVyeFl4rPT5dQwol7lN9lh46B9u/65bHswxM9risf2j3P7MVN
Ef7aKkM65NvqSljw1rp7/Fjy7z6axT3h/ILqFgA+9l6ZS8ctWrVU3EnynDwL3peo
zZh2x55dgVsPU4QpiICIPRkfTTxMg5therklJfbppbXMHI6VKkU4dGZd96tVo0gi
pnUUehg1qTbS96kV1T8qWbWTB01M1lLcCz22dk/wtrgv89aB3ZFNeUHalo08SkTB
fGsMe6R2hb1y2ik9m22q/anjVBiys4TiFnSnAooIWwsWt3Zy41sw9R6RnRTfuTJ1
8PCD2Zy+CEaylXxAYr32BMDhhKeJCSWG1hb3P9N47rvKNDBABMR1m55H6rGt9sFb
M+QQy7jZuepGtET7TsAXgA==
`protect END_PROTECTED
