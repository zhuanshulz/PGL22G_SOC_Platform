`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HMrjgLZ/fFKGzeTj6QWgFSepgJauCLgPFpwoc/f6ti4GpjtWOKktz5fawKvaXADt
zd1J2pZ2xuz1ZczrfFC9Gi59yndc6Nn3nK27AL6o6+z2Tloe7/aM4IEmgPrmFJz3
5PNXZX9DFFMguoBLvuAcTyszMFWVGG3hRfNSriaGWr7oYtwqG2EALbLldjcR0V6a
uNF/Uq0QtIej6Vd91oTY/B1L4Dmy8dMZWsDZHrqMydQMAK0bj/9g2PGavzzlAAqx
1P12Luy+jTvmST0ob0eV5qX46/A6ji6/z67WNIUX0Twwjqz9DTPsWzAbY7UCGsA3
52oiD95GVGTfyPzS6bHyCioapPdSMqXvFLI9ei5NpvfJEaf4123+jU7zW1n4REg+
fx5qW6aJvwhiSkOOkdcDIv1z4qRvwRYAOYruFCEiBcfw4txnRCqrcaywSDa8vm7C
BALLy5WjTSw5j0HLsXvfKnah7IUpq8ld/OtBzSA9ieTPEkrFIsnx7HxqsTE5MCZt
No0F5mKjPqqnjQsn9Dvang==
`protect END_PROTECTED
