`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uQ/WPgyX99T4bDijG7RtuRgVT3HG4xCR1g63OkPGA/+RDy+veav6ZTgUYI9zLVxj
/JyvIGy+q+BSVWxjpKQT9rw3dO7ZF/sn+NUJ+WyUZSAmqyq4ri9lc/ScosvuCHto
L5e7oT7gwwXaekdZq2K5+k/ZAX9PoIaTu+9zpP3xt9KCHD0z2pGs+HFIUEoJCLRS
Mg3ACK2wJpeviPosJNSGC+Zt63b6Wj8DU8Fit7wPNBhRcnvPDDqIVagfpW/QjxFj
jrZmcxA2JjR613h5Vvyy3VO0dvsJ5j7PRIO1/41VNHW8j0OYILFDPKs5peu26jup
`protect END_PROTECTED
