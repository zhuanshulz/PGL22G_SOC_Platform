`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
byAW2i0/SKB8DJKgZlufo3ZNhS6EnTmTR92HlrCPHcuBlrTPtIliZ8YRoVVSVKgF
BslK+wWpVgR8GklVY1WOIThg8IgdNCcpoydjydXsItxP2uP2EBBIZ45VTC3GC456
Knt9BBEHvR0Cf+ts5xjpH9R5+IkRXFuiZ3fWKGWieMQxbqw0moxZAFG1Dnt6MhoC
4XdBfdWa1MyPvyN0K7ASsdwrbLoQus1UM5Z1TxXCiPs4fJ7cXXGOEM3a/0JI+Kcq
aHWOUQWgV6ATjCLwHMYOaChtzyRVIrkSyZmottaesYAyiuVzNO5uJJeML8nm090r
EnjmjctUhgaTgkZAuFD5i8lAyl2GDi20sJiP7WfFHBVwqI0yjTy6pBjRx7xMamKa
yq8kVISflL+h+mOtUHx+IvdPALsI3NhG9uVNcj8j6VZuf/Dcekul8fpwSI4klSuy
KX6r+Ew4jud0GaJmxUp4Q1HH+XjKIFGA2I9gf4lkiC7pfJ3HuHVNerV02xstY/XO
w8BN6rWUwG6/l0TdJGft+pkvxYvfZJfmEHuAnOzFGV8QpczOXu65/+tMsKVKtfDF
mU/q9hd7/DY2JbCp4o4WhcRWYv7If6IoUBpzT5r5BFRS3jgNGAlDE/+uHohGm+t2
ZxOEXhZvP3TAb9d5V2OGYsbW8EhZ9kJYcFBFIYDzfOrNy5jC72K1jijt69peJG37
4gK0FT5ZW1R+xxGprZDmgqFt+0G8pLOvay1C1yv4gp4zKI4RJhHW7kk9evgcbSMN
oUs8FKGN1fncjM/WyeD36K+Avybu8nJqAax4c8IlLoQ4Pu2OucuN5aLQA++u5793
wrHA2OfagCNXFhtmOHJq5HkaicyEYNzfphGKLgA19hLkQl7ueUioHBA3y5Lc4oVM
2DSttpqe8JWs8wj/hRqyR7ThaNcSbSg9RBwGv5Mhu7jbJGDxWHUgjpX7O1UsRx3Y
yi3ziXi5ltZO42892N7LsYHhCuypLoVHkkV+CEnKKJdu7jYU3JkJOeH1JGOPJinn
7bAPO96IWWQMukmd3n4Qo1bWOW0/hbhTvUEH4Uyu4Xxuyr1q9tQdB5wPdHHygBC0
uNMpVNsI9E/zdo/Ul1tWgY+nP9lV8jD8X1VIZbVL6PZFmbPx5oXS/A8FRpg3vca6
DXmJedG8pvsIi0ZsTTt/yh/m04eHpj+w5yNP4pr1VzBKTm3yF+1UdEQ3k/+Kxhls
hGudqyDACzUBJMHunct/b/z3amVHGZqx1H9RiBKRc88jJQQhgldFaL+8rvjgBgnM
5VibqPVJvKb8pzenyRPLfkYVdMdBqnh6oW6JSlmtpjJNPgXs+Fp0gciv8M7jFsA2
9zrPiC4SqxEVoapdY+hUJrcf5M59FumypQM6YAFezzdTMk8YHg0wkp8O90LUI4hY
74jrwbJFZqH0bbRPXV4dD5R4jefbm9ruX7xOVwOTrwNrv8qiOXO3qBY5OJyJuBaC
L2J8RP12uP/uo9+a12PxfGwyGcaZEWfZGP4m+/D4MT4yvHnijUokp1ZCQNGeACh6
xdYYJovj9ZP8ZadDYz4Cs3zmCXK20d9rm6JJ1omZ2VSOVW0crRzCL/ubBdo3AY8y
YqlFp7n0pffXYeXPNpAE4k41kykifCMKnafZWx6hAByBntIhHNWtpMbpJfcWt7SC
793R0wlsZ49V4o0BRE2tm4pTeGuVKvjhAv/NFAwIPAB7irwIWdhRqpvHseXlp0v5
2vaZqxJPPhz2bjfRyHau0mZzXd/i6AQ4nKQCA5O4hDOEbwfu+5eRtFRDdiKOOOtr
Cow4CTOJzSOGyVK4F4NPje7wsB86vrc6ibVxCs6BRuoluxMRoMPBll0yTXpyPcIj
q3pEH/OZdf7dUJHLBWpj6nrefvI17hICWL0+FQSGn8q7TAmRMzSjjL2ESwjyzpWb
IZjvHgvPnij0boFNlVyXZq7i0VRVxcvcVxeKcFgqguN41Xvc1rghVhzsOsWP+Om/
98Tvajp02yLBEWNCIejsDulCnmnSYnlKTY/ZoGcujja9GGRHuDcMlSpbSdZha0DO
PrEZHFcvGROrMAC1ud+kB2r7f8X2R0HYeK55MWm7q/8S1zAzRhe2qXUci/L+frwC
NsbKF2T4PEPljKwVfbIITuvSyDKHnoZlk9ry54sqOExdndzNmpSp3j+j5mZgaPjr
fMzu52z2JetpYK7SYCSNsVq0IdLomBEfCHh5VXdxiseeUIjb0izUFnV8GRCTUUmn
MkmracRBedfb2p5+1UU4XX2AuMdA8gkTD78kmGcSBK24n/glhyvxZci4SK4g4kvo
aRdzirWGPKlA1ywRLcZVIbhj3y1MgH3mf/6lGkBDfSynUPY6VrcwuxO3IFc+oy2B
NMmUPPna5d09Pq1iCxxLWkecuzzlzf66OTYC3ClKvgU2tetIbCY2HD0i0CDwtf1m
g0Qvx4XWLCTYlDk7qNDXhpzrgVGQMDY0A6ftHdFUziYmEX5FQkccLHim5yeb8Pxp
06foQudQS8o4pWCMLv25yYmy1ZbW5aK2uDvMxpOdTeJa1d8eb6ixB0IeFfJ44BXb
I4zEXbD079beiZhZLVIfssO10sqr7p3U5F1fMSgNI2p6aOE97Fe6uPnnr48v/h01
X3cjz6I7rFNVUO3tRRUBNm9gkEIxyhRQPP0ZnuddOv73zc4UBwu54xwMB6mQn1VP
Or11TAurDlvuy3C98ym29D/G32+ZiNmyNjzuC4tp6FNCliG95CBYBw5p/MLlRUVW
SzOOPo5GVZBi3ZST8Vkgo0+uhaYAwGfJnjjLILP0IhYNdZJvbPDBXIxqVMbPOJVI
yQamqfYPevourRXZsNRNbYtKFRZCZjgB2Ff6gcDFnsglh01FH2AObU9U5qKi6p44
kJ3S97auMmxSbAFnNjXXWhHfB9ybS/7xqSSe0cbeXSah4uXOh0iJnMgKAELK3PoM
fCKDPr09zwX0Tu+z5SGt20urB7YxQw6v/IJ3/5VXd9cqj4qDEKlNzlA6eOHITeu8
WDtHzwMXCuF+lrxZCLn0vJas/49aRMcjfwmE/ZUxJ/6TUhzLTfwrxtZLaH/H2ySD
WlMgxGfmOV3jRL5Ap61E0GYGpztH0pA2Zd/MJnUZ9MCT0zVT37MwQJLIz1h/0E6b
AgQYiq6qs59rwSwkeupLt/ffvh5yLCWYnOCHeWTgHt9eG7IY8BZtKVY6hwxqdrLz
opISQ1P+jkJ1QpxhN0nJhZV6IDNAj+UB5bqvj/2oJDd0Q1BbXaxmi3pJ8cv1ysQB
axpfn8dW3qQ0y/uK2ikdpxI6A5k3DxEAvrMnug/JjhjhsDkk8o0OVmLQksKAaMkn
WwU9Tn4g6n2S8hABnz/IzRSdvwYC95URQBN/2AMkc5xWIg5t2T5wgyJMK7pQYWhd
GBB4JVqc0xzFZ+oKNL7oEbd2EJcSXtfNg/KmtPVdNhweSwjnjKQEMemZcuXd9Fm5
RVIGng25aPPzpvSno4mMu7M+8a0gaXp1/aX1kCn1HEYFGeJY5ymmhwsC/PMk5RiG
hE4gsRT0PKnaCWYPn2s64Oj7C8fxDGwEHdIfHZxi3ym0kfNWVtj26KtEfWeK3xFC
K5IhMNcrhJnPCOL1k4EPUQv0IFac3wLhaca/Jh03NN3Jg0Q4hZjp9KnMxO/+s6xt
RH4zhpmaTFqItsuasc6SXyHN9/u5sefsV1PyicckCgil8aAObsmlfXxaf/mEelmC
5nqTAAEB+lYanG5KnQH/4Q5y9y8kf4eodZWAKr7titNDE1JuxDshNLEcbtwky3k/
oK+LMgxsdvO0lCmVDrfNfnhwteIeocj+QpGfg4Jqt9B6AMvbWFNMj96mRr5ly+4B
+Yt232NAGjhS6Yre6k3Lzhed7tSi4XZEwQoWN3nWuqvU0GHuSKLKBEDPRozRZAPR
c1VcBS8dnecgVkQm1ZnoMjpO8ru2cOYReBwEc4xsxifvqMRgQZdtEUj8hzomHU+v
32/I0tUhkc2MXQsdk3qOlDVBnaBdB0gW2WKpYq1mnB8=
`protect END_PROTECTED
