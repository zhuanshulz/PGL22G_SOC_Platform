`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I152YGSciwdPBB0f2MzkicQSFThxrqew7cXdqWSdFFUQd60GekrxruOhbSg81SRS
rHmfz3FO0ny6WCOOUQpXLriQJxo9kYJpiXWc/LOaJNXN9W1SstEzJITQZoAYihGL
/11grTogcnGlI+ohk4csLVBw2b6hIWp/jcYusVXncfC/iqR+uGnRcxHXuaATqExu
E0raN6q3lnUlIUfALPQgJR2hAJDfRYo+6fk2DMv0lDn3LG7ixzuZ23cjLXjcPgJH
dpfsUh5ljQ/22msdTPoFoqKwIzvHbqUFJk/oPU6Y7lAL0VnWASbLa2NTEegt4KTB
CDeQ6Rl4Tc5KxF0+a0D+Dtk/7BO5vgvvVmXQBMkhwhWra2S2Krm2g+SGCkVEvo8v
vlUM4+n6wkn+sHu2r64qsVSgI/wBBYndgJPJskqXvICPTeGmtydx8fLpw33Gn4OA
WP40wgkzZNttS7jLi8T3Om/qJA8oTjaPFFAKmx3xLUrTyjKuc6tN5lPHJN81aNgo
B2tir5GCZ9Q1ZHA74kX4OnGUfQnK+wG5vQBx75aS70WPx74aesh6GysuEy9nx3xu
QXvBFWQKrYWWatUq7bTfzDkk4ioE5w/TKcJccoTe45xSeKi7kGdbfVlHjI4Hd3Eh
Kvmt2FCqC8os4/btrRSnu3vsdXSwpaRSQ7Tgh1TCOgtf+eAgVqI5PuTYCQo9Rz/3
qXG7vwbHbYDTQqZjkm/G4rUDots5XI8DQ7H1zC1YgK9q5Jia/iUDBKAaAWlQu6BQ
juj+hdUcSF8Q0dYh9ZzYXe1zaSjHkXX1RIW8fbbq/HdFPJQz5s+hJTFY9UuCPMCv
2RG2EvNTq/ILlutZaXWUQZhfqvEZFedPhQQcmFmiWk4x/BEEn1M6PXMGvGU06x4V
`protect END_PROTECTED
