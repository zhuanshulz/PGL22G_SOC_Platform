`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YLFxeJpf8Q8sktOqvcgJuJ2D/q75PjS3hp3h0wMygT2imlViAcZ8w3v7bzrcT48F
GP21sEUZQoNMp3V7ulpvGdoPr0qbTRu/sUAs1/N9vCRbYF0Xab+oE4wzkzUXOsTm
GEc7dYWtorLIQyn2khZdLMf0gTLbAClwODzA7fYYOqMcQMrBTyfiXqN2czYVDKFu
2VZjMLazMb24Y2dyfKU0Rwo9EIu597xkW2NLM/zaRX8TLBDp4U7lY3B5Y4gStkRB
AXoUN3MlwWMuhxs3tlmUt+3J1YDhvXVoi0D44jLPuY96r8+sKdVlwvj41xlQ2SXG
M9KXoA/M5VK4i1iO1ACb+QwmT1WyrOcLDeZuR9aM0TvVBig43hKmh461PXhQf1LM
oU9tZYIpS4MIUxFVoXGMQicvgtpp+0eM4l5DL4FyXA2w8wRxgHCZGTRBO+Sjtp5i
7O3h/OJPUVAFnVURGbU+v2bTTXAi+K+20YDi7eN+Ngyz/rJUWH5lr+KeCCSN+MJw
TORTs6L7o0vcs1kHCiHuYzit1sxdfRVb4AShzmHwH9p0+6DAjugDXCE8x9/61gRl
gJRrkFGBXlasn6QA0NKSBe20CQeZsLjpXoPC/d6CrcvnTCLo3RWF1JYLFIBG/hn7
avDDAlZReL0/kqQL4Jppzvz9azPYBVgKLpqIipXGg2GW89HUOkLCe24sXBo3EMjb
Z20QCeA2bmJ7j6WGjNCdfGoaHPhmO6Q6ymivhxe30oW/0VH1OLRlX7Jp0btyE/ZX
1wwml+3/hgSIC0P4nKaAUmzdn9BhQZL9vOl4lIZMVFOlZH1d9XEGHCfb2Qw2ZtSX
UkluVCRk5FxoHEkI4U7ja0hK1jn4kLy9z4Cr3YO27r9qxN/Jo/2Yg+b4oq4+upIR
Ww/n1xsJdZsYmfHRsMrwHGKRPYieZ4HguKRwsVHqdcEZz5BO96HtcwEPZLT4r9V7
8RRbUkC8IfF5sYbJcKxFadiT4DHGwO9E0B02z3/BtmqAqgFeOoIaz4+2KnIfAt5a
YmMPj1N5nVGXbKGB6gRbDftG8uWlEwc3rJoBreFueiTIfXX5UeU2JfE9XQJll1A1
IsWl9pxj6JW67bRfeiQRoz5gBiCiu22TVt9dVh3gKReE0BCplfppeUZ6mpOh602S
UdaELtteqkl4I2scT3Tw5xoosCwn9yiv3k/bETzO0LQ2bF3dca+7tq297YkTYkqO
Dd0fDqptydDQX6ZhS6VnJZ1jFWHLvhFfM4HI5/4yNPApkQQNa0mMDDkCJcq0dXY4
gMUMOA4eRShocgSsEvS0EIXTG5eip/w4RwiaoFZOUQq3gZx4iFWWzxexi5RA3yU7
gdvlPo4GL2/hwWf/2VQ84aOVTSyBMjwxwvJgj/89zEPbznhIE3z/H/OMOVOeWsSu
i20M2hlPWrervsqTzzxR8s0JwfSxfjDi4Jl7EJKSfP5c1RzK/NxSbGB8Mpe8Hqn7
GeP6yPzJqgzAH3tdgNJyrwqQQHYkKqX1l2OjwuTE0EMimNGihnTsSiGwGwml0eDa
0YdiUiJR3dqtLwlKOIShkscICtfcTCkDUWGuofIZuNcDa0rZicBfw/xqlhwX5FYG
gthgvHJwaNiP//zttUibdqFuv+cNqtHhSaJ67MRCnoPUVSroL/11bVylyVPu/UUd
HhsTPyQhhVKCM710k6bif3acn1wEMdU0ZPNAvJ/xj1ncRl6ZuRiwjv4B9QXWuTi8
gyStleyOIDCui2SO1FrxxvMY61FPjy98uQp9osigpdaDSxhDBwhraN+ose9MR3yN
UAyPxyGQFBFTDcUaPKS17ZbtR9bD0XqG6OQIFvzJcSaCMsDCS0O/ly4Gcqkqbvpu
+5N64Lw5uB5ULDmfhThl3RwQbbJmvY2TGllef9e6G+gyvUtrxPbx7uZVR4mJyHJF
E0AMNTtc7Vij/VPGmlzT9b533AhdebGTxuJlp0fYF6iIBDjXkzo6t99fCtRAIIT3
wEYi4o0PyJfd0n3i2xWxYKyVtZmkL7pRwz0RaCs3vOmDS1gkVNSTZY4qLWM0UIQU
Lv96wglJjplF5LlhQyGzSFzYJV4h0RC/bUB7N/B3WWR/mygBfMiNjcZC3pAOeXg1
fEkpfdiaT2PVhtyTCBeD63Ry0re1aE04D9EepA9I5quqkF1sw1yrER7QOIQghpnB
Pas8ifYYUkT3akM7QXnn95ynGpR9xaEnA61p2mCqUe6UAaugd1gABeMda3iVKgso
Rk4txPL3QDc2OpxDwVG3Cj9/fd/PfvfVUWZzCb9LQkC4PZ2PHeQGEsRD9xIPxWW3
oSHhseyqBr9yCdaJXY8Z1vwLbjFVvXQn1nZwxfBP38jSW5/07p4FQRlun/Ak2jHS
eijGKsUDVDM7QNo+QuIVrrTgZdvFz/fKU4aizvJ8OHzBDQ0tJIFHzN0j6VwnTZnb
wqgs1V2PmAWJBn31S2vl7H10Tk6Xeask/HnQ8+axJH4zKT/JugB0HbfVQHBnHbAz
j1wv/CETa8tUWQSmHsLzf/hHswUx/g89EDUTdAKs3Xb/TP3It+B98jbHK+nuO0Os
5GdsoYDCPwVnSuxc514eOkb2W4iP8hn/pYKdOUqlwcPtXp3VYcP3yZOtxjPDOTyf
qTPVcKRCCQu93XJUwydj8Q==
`protect END_PROTECTED
