`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7RW3HdlhYUcsohBh4ENICV5wGHRfQBFIiMj4r4809e9TYcNojYTsCCa5Br9WaEWu
0klxAcSKLYyP6S5koiyZgYwxN9Px+Sb8/xW4GI8hyXuouTdr/LaZqzldlohngNqd
Kp7lfmgf9K/Rands6curLc4dKBapWK/nq8ZG0SqQUnKmtTZLdcDdp+L9q3/oBhuP
IAnrWNUvtSLUk3xkxzbQU8T78ts3/jQtscjGH6EYxkYDjg3MfT5/G8p/QCjtqIGj
Ax3bG2mHTz5jvB4cT2uZeOBZfUa3u4hK5jmw+N1FrHuCMO7XJacBGw8gnqGLgJhv
8WkqvMno+YxMgnXCOb2UlLyApHZZoIhEjfEQMhNACxecK9Hb7lDZXCLev1DE9T+9
wd/BHZZs9Oq4JAteMvDpsk5CBjCssTvcbzKqQ2XUFjfi6NOQ4g8zj5Cn4YGXraV3
gZYf4P891Dz8sI9Ztn1vPhKV0s5lzYwdUai9lEP1nOBmecN0kVjlceqPXnfFJ5Wz
wBavksFWSOtjJR/V0CT7+d+2m7RhB4Caz2GgLaaiWrpiztOrG+G7wA4gb7Ftf0ja
d/r9sdp0in+9H1mxQSsCGZwZ37ThQIGZeRlRJEYGh0g8K+rMZMG+2DzYR3nUrJ1y
O3n26h86NcgxGNn6V8jpzZai1DJ4nXNcf2EoUr1tauduXY74Xn3rybjHbGTg3GYo
A1A/ZRXh3ml/+vTM8v7cdkNYEDMK3Nqo5/J6r5MwINbnlB1ZNLz6lEpySrOhveUJ
E5FfeFNzldjnwBRb46kr7/iGfKHLqxo6CCGEl/eA4L4rtG6icoK9/OWoEfH62pLA
vkKOUHM/c+kL8mJ2Os3M4Ab5PubM67IrwLbOmsdgQHhX0zDsnekIWJAAkIvLmLtj
NMJJdm45QdtQr1Q7zq3+Q4eGgAuQxWI+u4SMATy4O+b9SAYF7uiSbeA8BxS1OWGo
o4lNsIzJ15/THGSxsaeEyA==
`protect END_PROTECTED
