`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VnCsn/pxa4RNZRkHvbtgUhJYlIK0P7qytPg6SAT20KNNt2RtDHKQvHSgP1WTPxNr
+4PPY7ZHWE0CPhv8RLtu0ptAU0QX+ab1BJ3RhcLwlP7FgW8Hd0g9QrDTd8ETD8mz
PqQyDTaO6wWqDEPATmzi7LwOkyN+2QvNf7cyaf/ABx+Do+eknPkgnWleREh6zTN4
ExMErdqXV/YxQiOU5RObky04B2x2C6vLgRp1vvYWZ3LR2/dXomiPuQwg95trWkZ7
BGnCvIN/dvTtJlHbqv/18tx4tSxHPQPiEjBs2qNbIxGZZ9k6Pd2xJi7D0lhmfD8W
evspK0JB2QZCrNivregj2afoThLmEatf887Bd/wzw0+sLS+KSUAoXGyC+k6ygLyU
7jUaqMuz2TbrY63Vw19cA6SPKkKBcSnRJmQjLgQRO4mAhykMC75OpwsZWphB6K3q
08ajUdPe/s5GYtsYqhsY9FPbKbDCK3ZfzyPAXiuNMimhwdGrE6X3LpRSsIyF8UF+
X4hHOei4UKPjWhf7szoW2W4dEWY2QUL5yUzjFHSv7Y4IK+1v13K1O+fogsd3fIa/
ATA7sED/njNTIKbjC8LC5KEqg5+Ez1nK+SuYGyiUJOe8oTkvcpSotdQ8IdH8LgUw
odXf6SsEQgjA6LpHlfRHSwhVYmYxJcWmkJ5Rmmy/Qjewr7xzqJYwH29bTqpUkpBv
8bR+sTUYx3vquLgxiMs1EZ7AFTWN0Vw7ZHTkblT94TGQflXuP+EenvxrQ0RD+FB7
Ts4j22ghscBhTg2eGT8o2iSiHQPtw7c/GeaHpqIFjJguATbZu0VfOg4uOUeBuj3o
glTNL5f4HzLYq8AfRSbG1zcXieL/VTin+vY8PW3Ix1CyYjS042h/Htx8AR8W0U4h
OdKGRLVgYhHp8WEY0j9f3HuphKX4m6rzh5ox4BbLVOM=
`protect END_PROTECTED
