`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5SnM4SWr4k/znuLi6ASqNACiwp3qMu/lZog16Ed/P6A0i0G0dFmVOCZIgBcL/lVb
2ICyWrIcXZb7saOwMqJ9yQhdKyvwBZYKA2pYrzSTnF1s3qIgmYlOHZZIFGbgcjQ+
sof7T8MC3m+kXuGXVIuHjJomzP/dLm56vtt43YGN0tgxHgkM9WW0rxj0TdakdaIv
4bZ9EFjpkcsxUssU1Uk3yWCnBYcaekUBdwDGW9aJtCBdNxMt65iVrdZ+qUUveSYS
QFwHcb5x0xlsY7vjFyX3IXkqLmSyG6jACtn6822MqGMynCr6vm/M42+spXrOVDMf
WVf8xCy6DB4OVaLuDQ68FBRwts5T0ZgBGKGLKNFBE0kURvO/ITO/IMmiXYkVkAqR
dLxTtRkJ4JrnMGaqJKfttuWtNgWad7DbgO+hM+kQDkLvizlvb6DTTLD62CVGJsXB
l01dRSjyzgNsE6hdYk/8GKhQ+mf5v5VZVee/ydxHSBA1lJmIYHbDnz2kqrLUYnix
QoauqOT82N9oB/SCXFY1+gcKnkpqi59LbcpslkbGyJQXgkCizLLvDAyP5B5lPBn+
jXQ4ZtRSBHRTQaPVNAVRQOaB+LiH+V+RyMQQY56pOEC7G9sYKS2IU1gh4JkiYI3F
lvCtyZMWaq6ej7dWUeyR82w3BLJTxfA0TriRcHjjWcRZeUDaE4tG93oOi+rYl8Yy
0IL6ukBHLsciGVihkbHRVF+iXSEQH1LLBlwVEhWB2swjNy9uBTWoQ57+oClUUZ3T
hhJTKbMZ8HMqWuNzYF5OQ5NTWRU5ctfMm+JLkyS52Gg7yBRzPl0IZUTqPNT2TspR
wRoxApnZ7xrNQNUjEtiTNSqYhqzIAmdkYsT/N8ua7js13iK3+e1NZmTw98EOCvrG
hmqDkF6Koo4GHHRavS6+Nqoe+oIs/VEFwyR8fgRgrOMvGq9TzKV7zGbRvBdFISnQ
WJmZAwduRH/S5Fhqg6BbYY57t3EcGH9tWoPJ/y3fSl318VRv0cEKR5RsGcOD4IuH
pYpBeJG0DS3XbbN6lqZ3oyAb3VHRGHKeXvGgon/2Yk5S2jZflvudjB2oeAmhpnqA
kEP2+lsLXj2c7INv8YGcTc9YOm+iYBA+w9ex4+Wfbsoqql9PT7SRzFRq1ykO8XD5
CRjm6xNCeWXhhsZHB1SMR41W33K7uBPaiVI+8dsJQqPb+YGc2epoCdEHCl0R9mqK
EsjAA704ZUbyIiC1X0vGSX5hp5eh3f3p+OGf+SsJfjBkl/9zpm3mKVScRhbUcBz7
WLDBg5MtGwdbO9pybqxoxfKfvclLmB+6snQwQvmJk7bO2cs9hHKxWHTWDj2RmZWK
jAqXxzIU8ev3dvuUPl1ucqZcPEkK40wVhoQSsoibVxu+DRIktQiaarNN2CvZ6DEm
lnEPlluIuNDPEiBkjLVsArI8UYl0DAiwd57DyVRnWqJpNHxD23j4DakCaono8PEP
ZDd/49Z72cMn+halLJzYTene6WA8s1v7ryj+22yWxu+CfsDA7gnf8xt3id44NcPq
2uh32T/B3L5l1UA/Iujkm7kHZn1TcYKi2LF1aqLdjo0XrJZu+ipA1Wn6Bw9yjjRL
ZeVUesuW/V+m5CKwnDyIAsrhyBPGFma0sGC2IhF3aBPr2YsCmVZtrpnr/VDmHpiw
GnkjrWB6iqEyN1TAXGjRSs8g2oS6Hnj3FLF6DorphNrMpOWQTbGy+uuMfjWyy+Pq
YniifR1Ol3k4J9ONn9ASnbrIaBxkXvKMOM4fm6M2I+9rw+nc/05Jm2AOxijWxKQt
`protect END_PROTECTED
