`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mryhfson/RGpGMu9HJqN3MiBVm1XqScrglAg5nQAuniXLu2dArhY9HOci7haCKGs
BGR7p5VZmfNKpP/8VWm+j+Xp5ZjBN9JMPCt0Ey6jp5AJV5jj/YvoJr4N7LT8USwy
GI4fh6oHvYcMM+a9/W1HvcVW9uEb7vgQa8VF/Xl2m14j1VV3KHg/h3ENxhe6Dauh
m1CO2L5XRu/ObgrltxEtmP55iVBbL1CNoODO6hote1UgaWDmvCRnG9k5Uf/N+pOC
9QgSNu6YoOplAhYkrL6UpLiNKFPKiAEU/z2p8eteRtWSrO/90qVQ9DicIqpZyZxu
BtX7onihhEk2ftPkVdXCI/0jSmLIBFjFLzdZyII6vPRK94Tg7BJmDUVBSnk3LvxZ
6rANp/TjQtuk1qyW29A83X/UbA52stPd/cSTv92jEpj9Ua79XmTN7ujjRDgvT2PX
PCtgFXOIToIKa/5jDAyNuHRhG1gGT//jUd8RvRIY96i31lKxhTkSeyafnqvE2UfK
epzXUZ2sPsKUkggoqHivgCYlMGogO8dyAK6yyzAKoFYYvb5C00iJyKclb3GIRxWV
zQnoinyvdth9P6PtMSgEhR6J0nuH+BxOEY9lK0uUw6MAd0vjgJBxMcc9SNPmrJ7z
rEuHzxXMZSOKsKCr7dmBOQ==
`protect END_PROTECTED
