`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QvcJ7LU7OKwh68zoErbMpSlA6SfMz3hE0q6RRr+X6j/q+59jrzRRiLLZZWoIB8u0
MDXmzDBgx8R2c/jShAWGOFPXTEda6eriIkmOuP95P07T/UGdoKGdR4dFg1gsfv4q
eihqCztqXW7xwSnhZFQ97fm/OndTsiKiVSyyFPTXkeQTsDcyn0L81ImfFixdzm00
6zpV/qu/L6bekLLq7H7qECJxLj/nOD+/pgce+Gu1vixe1G/zZCsTeAPzdjHrxG9D
n4IVwIWscSisI8ppYqvCeDm4RYxM25NaPDuDNc0NI1bxGhK1OAwfIi8MltFtPFhs
y+gMOyBQCHJ8l9sxnBQvZg==
`protect END_PROTECTED
