`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d/CZ5kt8W1OtPkUIDDwKRJflI9fnDur45W1HKqyrpaOURaW+PAI3eDR5gRwRPc40
I6XKG0YjsrSlKWsAQkNE4Ls4TyhEbjb+bSfuKs3SNWorJDGqSNMe4iGaS9E4hFRn
lb1vd01QWkk5se+9hihsqW+n1W7jHE1u4SPAw48bQWJwJvrfmgXHSoFJaoTPg60E
ZX1vrrX7OiHESXdcLaLufHKqQuI3Qn80TDRe5PZHTRSYs6q8UFFGfMpqjeLEu/Gi
ficZXCxBcyK2zuXgy6fA/CjFK4Dx/YhZPCQo23XaKa1txJXe12sHK+63yBBWgake
FjuDPN8WsBkJ3MbJdrfMSbQTZiEkW+6UwNqnhijA/fc0XRyGAdbv3YCSrYY3Wt0V
0BwWvE9Nnc9DRrZOvRhEyoi0srH9MseVR0WFhsZC1fl5v6i1i7ZkyeM+nSymdjrs
z4H6pOE4ZAGvF2WqxKsiEumGl0sbRiw0T9kR9XNoZ7GtBsX9irfmFGbWKGcVVoxA
/ZrjNCzmUT61xsa1ZdCyQJ2FEdewJTgzf0aPy4UYooDq437Nwp2Of3wdQX3U7YKg
j6SfopH8oCrcVlS/8fAvdeii/XqEHHqOidJoS4Li7E+GDgjRmy5FCZfclujdBCqd
IE4HLE3cRvzzcC4XDbJHXBNvI+yFPe56rHW5CJ5PsGOF7nb8jSMBnGHkPecn0OCR
/0KYDnl5eFZfFvuoZOF6WViM+6CcWZdxsWztHyUtfQ5MGZU4QUztqB4GmyRqwuWo
DebZg6pGA6sd6gK02uki9QZv5P4Bd/rVE2D3q65zlMKGCXTasB8vY2th8z0I51W4
mxLJmf5O+rm3E1OvYMKb7aXu37FoSkR/4ilt2c8tNVJ/vT8iqj6sya56X+QjyWQ4
6QG/4HGRRcf8OBtWfqeCXUvlBR3CQTEzsIsCSsAEEzg6kX0TwVEa/mHED0jsHABZ
mr+eb0sgyhxpXxLROIo2gcB0Kfe/bs2haDWhu4VHDPh7v/V2iPtKGK3vYWYyGM+h
3ms7JKI4GZDvINr2a/mAGRER+gQvG48CtfuoWYpSq88+gQJBAv4PlfnDnoDsUI6z
646grdCsUkU+cyUb1FguAs/SJId5oz5dxtWfga0DhNeUHHElyv2UzJaYnOpEgyfZ
l/9HVXGna2oeyaaNIXMm1sDIprd/wOaPHPeQca9PGuAs8aiNrxzsLQ0+Wsv8i5oR
ClpZgMKS8Z1E20dFBJPG7RiDTALDsRfvJTxw6XJC16uSniEfBZzvfUMtWdoFRGwy
Uq+yoHag4uSlUQOPtNmNpIshzphLetnVVpubio754tXNcPuNrf4eMiKaeGKU3xHY
YXuLbFlxI5VZDwNySQWbP19U8UitIzcaoepaYZmnfgrMr1a+Knwkn+viFxvi7Enm
wGnM+TY5rnAt5aONd2255EKkuYT2Om8N6918ofsaKL4aeIK21VZLeE4Qmdm9gXP4
7ki4Yp4riogjE5VFjzo7H/IaFP+yQEakrYHzAuBaHI5I1K3MD+YOS9SVwBpDE9kA
YFwCSJqAZHnsAa49kDjlfnXtbNmTpbqxzTJNAfD6wP8v9njVFdaG7rSUGLGirnTU
BU++JUzrLSaZX+e7s72P1XMOip2iVSqeAm6bTfESqx5JrstpxLClmP0pv9gWT/pX
zb+Y/Dp3ZE0MO2kOxMTqd+uJiHh42VMz0c/lQ6oQv0v2XE0UKB+HbeQrL13DvSfi
ZoBUyPQhrHzTs6/g2USgYjoFyksXv8T90gH9VNpfk1AKCGiPIuoe/F9WDK1cyynZ
kWRjwJnL5l0Y7Aq2UxjiloBz8LwGLtVFt+bR1Ih6rglCAWRKKV8MCIGxpkyL/4ir
pTtwIkHrMYTUvOfIq46kBitcYxs2Aoz51Y022UE8tDcWaj/L6qPDkViupeLqKMoD
uo0xXOcjUkR8q0hj/11i3YVFcR8tkeXN+lJOZBLXIEZ20kPiEqqH1yCES6xt30Hd
JuaSYDjFZQ/Hq0vcJRxFkQC3OdMQLrzoBl9J3khAUReDlTGc/V47H1mtJMQXRPWX
Kdq7PB59FMMrhlgTc3v2MZ0VbQDqsCM0d9mqPwHOQGY+DpjWyzrBREjPESGJw828
R+nHeloJEOC7VTO4pFhV3ULxAvh7VoRKpKcbnZC3MKVEhf2GODEWsx3I7DKUE2yP
VpJRKnmu9ZBYWCi7gtJwa3kYYA/3RjF5IULtdu6W144gHSm8zaMrkkA/MmO+KNWh
PW0Ti1H+HoP96imGY9kW1E+B+89tG+k87lVoBFKIzmJtmbnF9h80ngoRhHBGJ/HV
qr/VJew8YWcOJq2Z1mCjWf+9ZZ3fr3idL1GNXO1itsCYe0QHKKw+qoheCer/HKTw
5Rr5g4E/La0D03nt4XE837RvC9myO55PGMDmiBF4NJlYAO1naOGbTxx26UMN3dqF
kBXvEe2EycDCfjXhWBz5N0HSRG2TcgqSsjVW1+/E3WVrfDlrB4htvUmMrUIRESMA
GhrBrVH4APPl+K+ufpilZ7bOie4VU6f5T29tpXPEUCja6YsPnNWJVzvtjlv+BxV1
hzBrz5HJnwIEDIpd0RLAC/wP/27pEIRCYYU7A/UI4ryT05X7UWdiFpnFQB8hVkxa
wMWBp3SVzAP2zFk239CFz6LIrD/6Eq66lZz+hxEjyO6cwIOmKuhyYy2D2sBKkjzF
BTaSKGCEhqnk8Oqd4vXbMJESnIXZyBiSMg6hHm1RLX2RW/O2pvagbIHyJtj/bDuU
q5dzKyd3lNiE016JzbmpFLxKj4IHVOEAwJIsRNxJSBNa4NWpx0TM1SmQ4xA0ESpB
+vD5keyrfEbz/SKV8W50EhY8uqAsBHiW1MKrvKeZ9RrmSxR6/B0EJPKhWq3nbnmc
Hzx5Kn0kagMerXyQ8Z/rjFQimrNWbBKrHfnK2JUOAFaqvcFVzgpc8BEInQhnZP3H
OVUpaYXWMlGORHhR0WVaNZWpZsXMA44ClMHVTh7WjUQN9cBcrQQwnlCWR62vA1Cn
AqhTX1okLvqxABj0KgJTsO1/EL4ZLbNxf9UY31qdDN5v6JUGeGpQjQuBtTGAkmns
ZgOFN1BWJ2UwsXgyFJYqTUCIj8PzJS/7oiCJsbe5SSSOhecjgow8Kwh9kL0qPoDq
LMpAheqEIM+1EoRcLVcb1OMjydTUU2UipmIpnQvSlWyp0lKVuUH6CjmPUXjyEIJX
bg2qExKuw+wJxks2uErpea+io5Ng4gxBYqcYYjklVeLYB8rEyn9W2pFTrYh++jn/
xvFdmSTEm0CqcvOOxvXZhxPCKFKpCLTKhrncAlFkh9YyeMQwRB6avJKpPlaXP+cp
j0SYOamPP7moCFeqdgSSTygyf+OV3zA44cllARn96TcCOSZi2FpcjVc1lHR9nA5E
HJ2Mi8kxgWrRikYJnDKqqTZDcIvymYAvIa8pDd6qO/Fo8tT8VxtZLc/ur297yf6v
Y24AYzO9MjHUiLuZHOQjW+XByfjPtVNG5WlgDwIpQDf9Ogw0hAoewNhXmG0YJU7N
Qf7RD2rlQM7nHVumJwrCo3qEECJQIIqeFDPvJH+vKLKwHfsZx7AIeJBORV/b/V7s
bWHZ1n+ARBAM2xA/DNEQlvVAjiCZTGBhnvbrbpDLWbPzvdMxoD9cA4sAmPPGmc2u
mdpc+OLfPsr+07D18d0KDp39XRH/PAyojiiMRzf6Zra22FpuCUBqcSljoYGh+m1V
4z6a1DYRVhWOEo+g+0i7gBdt6pHBUyYCtxBnTq/VdHqgH/FhgYuZ78pezFUq4hop
V4oX6r8cczLdeSKy8Wnm/eve3kq5AuovQzJgVd1slJ7JBxiN3ROCqtCcC2xzXeck
PF1QojA2i9PVGNaNYHE8tQAiWiEfFvoQYXyFLivTDV35lXE3KG6mIvL9iaNp2Htx
RfSgBIRpB1gCzPB/4SbapCzh8TEfVSxFL5bqPyYTR2K/wF7UPPCxA4sEzr9UTA63
kJs1wpXFh8iMWJZOuLB5fbq8i6R6lR7DQLYEtpfqB9upZYssgssANDirhkqEq9Ak
1zC5aWHcNk0xsQruRIFxe0Ras0vCo67tjndmLuZH0Z5hIk9yrA3vNTyJv4IDMMMS
h4FWXcFiOJRXcT9hL5engObKH15R1tw3oIa9NmEY9JnL/rksqp7nIgWQip2EChCD
AzS1sAXoDuKNJOOP8iCicMyfeF/BhuIuon+4Z/rbeCwEh+VzzYDQiKa8ojsKp1yN
cNccmPeQjhPsB6cKNdBgWFi3tkWjiQbgMml/s6oYal9YcNAeo10/Jaxm1rmKEWjv
NPnZFK5B9NIbzrIBSVvLmPXBRRNQUxTuJCNsbJtOHHqjITDfcogPwJ+KvhSC1NqJ
iMEKnq5mgqm841MpW7pfui0A42exOvfre8ur9Afvh7ZaArDGwJEOxLS7kmGso3lE
Fdqba799UPo7Mcr+S0hQZuuc9bb7VFb6t1TEnSw0U24+Q5K5DlAqxRggQKGVfDAV
nNQPzo2zNW1InD/SYPrEy8MsaC5eMBj/RRS54qJRSESrjUHI7AdpE6idNBfr/C4d
1zuCf3LjCuOVga8LSPDPnAu1B++A0AJGdJHt5Dc9JNo=
`protect END_PROTECTED
