`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PYzuW+ja8VFYjqjhNo+mYPrg0hHjn7D2jLqkcx0cPgUV2zOrPBuFacE+5c4sZ/NN
DDYd5XjTYm6z1JjN/eytFimLwQTYtTTfKJcmO8NnG5cYgbo0Lij/uTBoXWYNBR+Q
cEP60Ume4IZ8F5W4ZRlGDwsgP52QJctJR+N3d7yDHGXLQdL5lyG7naGSheWGUy25
xHPvFyBc/6FV9vyuhiPkbxXG8+3k0ZNMKE1JYFt6Q7I5VvP0KaYz3mNcWTZtB0yg
vPyAZw8O3y0Gt2eYp5JqCcrcRvaAg1J3ANfBjKNgE2VYyGLMUBliCMKIulIPUOVO
5sD4okuaHTBTGFa3mXeXDANcaijc/rOdvuxJ4nnFffvNsj3k9p4F7FO7PiiGfCYA
LzhoTCp/SLSvvzpqchKr6FQxEEU/l0QYTXB6mx0Zn6p2Y8BteGS7QBGhcc3TlIDp
MNHB+xO4vnI7jrgHACwoo1KtEQ904LBz8lAH54jF6r5k+xvn+Ol/Dsy6UCnHEQtj
k+ws//DfAYDD32pKFLy8q7nUDiLI3LqGZnZNeg7eQGLyNOlgdqPpYrqGoXV8Zcvg
`protect END_PROTECTED
