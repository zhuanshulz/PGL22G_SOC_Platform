`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2kqPXkUvFwk81mqNMhWcUSM/MS1BixiUxN0zB1/97OP49CyfRbNYEZnh/gmXLAgi
ogXE+jiYXKr0M0Ki10vcAzJTcV4L0MwGwvoOUmdC27wmipGLpNKGWKDWSeAj7nYD
NY5QZFXNjAhoPrtct2XGwGgeBsMnKg75zzo+X+gTns39dPeefsGOkoEwugFX+vKF
kkEmHw9Z3eXfvKISMrCaAAI5zyjZxmV/cOg0VUcPzlu/zE2au39JAw6t+Oqq1BJT
ZXG0Kaw1ZfrfqjRsyCHizmuRkXTmp4Xum9UMfvZNsC32fEvWaORBwuOy56giu41j
O04R//bCTSkHsrRTtvHVW+4qgJvQqjBCCuaE+dstpADUNMdNjHTyFai+0KhZXYIw
LlQd7PNyWmRQwC1FKN1kHNPJ9IdXP/fv8XaAdKUh4WBnd5syYBF1q0yyshldm7K1
02QmXqoasjw3Yc4GtfKyyQ5zXYNElY8hrZYa2OIicjU8PK7xdrqfO0viVmnbjcF2
trklRyaZcIxDr4HkY7wzYoITPC6jd/GEdEMDa10q9/8AtFbFVjGjpM9L0nzoFbaL
mmUK9hTsQ3JlPlLF+E2tIcXt4lGf/E3qstYoeUiFaFciLSDtPT/hSC3AzYfBSg2o
dGJ1CXH5Wu9wv86521g/rQFAs9BLWkd5Dl+G4VR7YlaXgzfM/HzXY7+7gAIwY2+c
M8J8sh4KJeAzJiYXHHp2MrjEimFn/7HPQbEKgkR3GBMOwwVpmKFdsfYRQ18/SBmd
uZFVPao/wece9JMVilCCILcVlA6KvtbS413m57yVcp6l0trgK1f3MG4xtFhY2id5
k9REjL1y0iaVvTCPANlCTzm4G9dyiSlQTSklCjGi2n9rxKFrCWjwGHsb7yzI92TA
m16hbYhmppY+5YhJG8pVmIY+6oL/A6yHW1EWx6mkOK+naoNe1ektgMqUZq2qD5uH
/w5YyhxJQ+DFFqcQjCHj4V6ug1htqE2CljaODSgWqrNOj0e1GaCjm3/3KzjZqvgu
gSNqwUE18BOjhvhDjHZ7BZwyXc4nChn+QjAvFl2P8agVdeeIleMcMVbdtIgY5RSs
mI1LCFC7HOXPyETIVnL4CHnliDPgucZQCSYQL9u7L2fUQrWZDZdgC79EpbN/2B3H
yrES/Oc6hUQhohlMC51Ids2XL6YJ4T2jpCUZ+wwrd5UpVi1Pxg//1AVOUmo+FCOB
vuQLe1zH+lcSEPLbHgvH5dMCr602U70nRrA57hVEzVwuSDt87/KMrVpaCvQL7jwa
DeE9F+I3ggDguKKOTjHS5etjruQCf1khEAf1Un8z89PhO4XPtlTert2jjrsnrRUG
gzwKxc6Wl2cMH24rF5pd3x+fbEVJ+3/vdY/bB4k6jhAy58+bugbK2283mBNjDYPR
OrCOS6fesAowmHpMyIM232hZhmyEPc2OgNnfO5LpH0iImebwZdu9CQy0xgamf2PM
ckAyd2n4XKA/XvRjJ5bF/KkbjQCUW+HKxFVGumIboupfi3q6DOOd0jMjhaDzeEO3
JD6e7QdHterFP0KQferHTob5DcpDLQZ+qKFEZHBuaoW6JAfXgZfczm+cf6ge9Yn4
x4kddIWOlsE54cI4911lVPsc9SB+SsjhV07tsbjIs+FvJqVXmGGpZH4OxlhX26+f
a8i0KdxODrhJAmkqoV4L4K9LcG6vOMRAyhVBmSbAbHL2uNkAbOw4P0o7FBrZAotu
6PuhpTXHrQlKfIQTJhVHnRDFB4w35ESwZRnbQZOejvMQq+XBGWzGNnab8JV6Qii3
NDBre6ra3O/kd+Fd41rC2h+oky4Et9AM8dULRUyxXALrGBCA2bOyQUtEzTBgKqa7
oYUH6NjHastpm7RuuUC3YKiPCmUvNl9C6CzrEQaNl9fFqdJOTg7uhl680AFSDl7H
evCuwfNfyXMcRkJIftWW0BlKmzNRzfvXXLmsmV4hUhveM4wOzyqgRfpBXaBrRLUP
WCxErAfdjpfHP6uRW0tYh/y/2Ia+fii0bOIjOXzmJhIy6sQe336lWnFD2dTiN6W3
5AKrjoR/FOZFM2qcD1nShGXpor84auncxqa3akNGPZ6aiYH4wkqGRuufnLaNv/3+
lR34bBjSnq0NdFYyfR5ggOM5U7lKGJf6mHAlPrEXXzL4UYSLujmHtXmItmTpPZgD
VZ0hdpIpe2yxZEbYTGQqqsrd40grR0+jSasNjxKVsX5Oe1I8fCEvomSi34JA6JJR
535cUkmic9DkkqyB1UlsaevZkFYn0W/P65DiPQUI4QrACVTHKBxx+jCFA8eC7zkg
5NdpBkD7GOcFq6xThj+/plvQOa+gZUTWmeaiTA/NPb9zIFeDAcshwYPntzJUavdp
cjUMrg7hYQf6uUUpkv1Hwss/h8Vco5JMnYexJ+lA8+sb7K1yFgWibprNc5WSLb/w
/zpdNv2EKKPLFygB4JKk95QrlnklsB8E5LfC0kXOk0O8SVpfi8dFGz6qduAfu5XP
pegzdBA2gsyvEp4oir9QHTvwf/IClU3P3ccWb9XyBhYrMJd7wKWBreIArgeVvYmc
m2PFodgJlTqddUwzMrs5eLVnwUOHI2Mm9ejHgI3bLzs8ccxTg4i3YfqRO6p0FhWb
uU5P+VUgML/nYNQM1rVDxSgQHdgMyrUdHNypJGD1VjTVXTvbgmSnZYbqsmqBSdyh
POoOjPvfxmwLzIG+OgjkclN+PP1EFo0oXIpSPTK4nxruVpsO5qymo7yXhpRgN3JG
/K+DXCti1iuN4iy9BySbdDOR0LVON5Vzbvy8EIl0snn2CtMkuTEyDiVvt4Mrr2pq
v+pTYBel36Bs9x8aL3UJ/+mqw0f1bmgB/usbcokBYEdpj+OXi9XnYEEUe4OBg0Eu
vY22p0ntseCW/UIoVEFG27/P/QdvxYzqP8ac3HZf0krEsYLmv12BMuRWQEKaE06f
vmBrgYT/6Hr29p+9krAO61QPoyElm/mMwGKknNTDu8JBLfSNYqRMNAGk1GbhpdiK
P9+Lmwp4g47AOf9QXRLc5q8cBFWk+yFp8K4qtbRw4k/Wor/MEmARxs3tQsYZ4+GD
DgDGTiN325AnhPoKRP+9P/RPWyt8VWVUHEm6ln5yPfwbGAiPmKPGZXZ7a5a+A9ZU
3GwRCQ96DGliNMJdABsw45qc+2XX44UT+bXl7QXXxwpJOJoK8QtsAEtTDZCpkJy4
1LB1e6lLAvnqMlgiMvrcFesAg6fmcEKkwwvW79NCHFFubMcw8zAZKRcim3+yzteM
2MUQUHRX9oj5S3dg8rorpYUal7gpBNTyopa104O96Y2RRPzUHuXP0KpyfNDJGCv+
0OQrIAG+UAk1XAEEmY8RkveUffG2YX/aBD/dko5XlLes+C6YA3q5lCFCLs0nBW5U
GVPboZlDCwYRCyvyeyM2RZRrNJu+TL7H8X9RK9fXE6RuPUWn09vupwESzlnSJ/Lb
5+rWSUwo9QsJy4Hg40k3RQa9D/dLGexwRTo+KS1urE9ofQq9m0nqu5H9a8/b66UI
aqUyelljNAnm2pMtziX0yiEXS8yqz32fD6bX/PChym8E9F5pIxRnvWabaKVpC6Zl
NXpOUJHHluycJbJMWhPRDg9C5Lwg66mMRzlXmcX7gzXqjOxK4fokZezr/TzBU6Wa
ceJTj9tZ/yDTaItGiMVIXaasXE5FIGWCeZwxWYObJFq+I+V+l3XdEomBWyyXP07i
R2FMOeU3SBCSMei80W4yU1EcGKy3j5Ewap6aIm8ZFF0bS24FuNlYG0S79kRBtgsQ
EJHIZi9haHP83aPw4L/X5FG2sxDMdvq0cISptPFom8IzmeMFNDLmvdCQjfkyv+mx
NCUpKZFZHFRa6k8/h0l1NoI9k+ecP6gt3PKTZ+FimAanFIJ+vskFusuLqqBxYgX4
hhYb/+d6oYkmvOyYPoZoK0+8CUIaPik/tq8A4rO9jQ0A+eKUgf5TgPYwpF4tfCL3
AcFicwlD42RIacyqYHuM7K6K0MBZIAUN+PEBahmacCCZmxkZFlRx1FoYMCCBNJq2
Vyx6VkeEpQrMQKV2ywt/+UKarrExai8sD/A7w6zPqVrcqHUny774WXn67ncNSGZ5
3bc1IcN/nUMvaCmIO1h1QwJJ+XkTcsKSJS2UQVqB9fTM8h2pE9aklGv/Gv8gBPd9
43aes7Zmjsvw778OwEmgp1MWmw8wpJuDyKAZaxZuf98GBI3vvrOSV/QyYZ2Aqxbl
ZhNvvYXQVERrePpHxFj3LL+uy7WPVcGv99xyYrrrhqlyruRCvjR3Z8Qr6BmoXdPf
O9SYqsjdW0oFvqR2T9h+Wz3OQV5lqxBevdjCU9zr3SXqllS3wXM7cx5uRcwsCcva
xVIMcbMsbbG2Zh04+7Kln5pfdEFliBe0CGg1ez5UM+HP4sM/cPNcqvqCNfzjd+RW
u8Wh0U/+UrTZOkjuQjdq3oq8Xzl4UN6hM5jFZQy7KvFC+MJqpsBCzdX8w+ia946C
GO1onIiizW6fNLEi4hLw87VBn+eZET7OIUs4HB1CjtHOP/B0upeReBzOZUshtTEZ
/Q2HLW+bKrF8ZAaqpLDX00mDneavTWCnl1kRY059k4F1fhIRssDrNDJsEBXpunKw
leqSMEkewZtVhF5r3/nPilfgT/u/QeMMp48metdJ5gws1vcyiJGcFdImVUiViAQd
K2c1wdt8OlWoL6YTCqRMF1n1JPcvOS+9RIX0HfDCUrY0FJtqwlWbJkZqggNa2Q4Q
W0qYyMOh35DqI6Rc5DYZY0ligz8sejkAPyuH6TCvwdfm02R1IXyw6NixPYBh3i9T
Pe8Oadfq2z58nXjoCWf2moGPaRbikAxftl6yMylvCus7l4NzrkyeEEkL+tglFdRy
zqS4TXWfBVExysTRNVaPDOHHBBWKdq+0Ozekj4oGloN3U/sck1WTy8dkvGilzpHE
GwGLukRHrHHBBOiJNH+lcqSDACO7z9pJtYf9YZCYwKo2n3YjKzC4ACWy0QMGwS4D
XV1Q0LeD1LK2VxiHzQs8tf/4X2kvtMoXCAhkbCaeGU31W1gukXneGfE03C93eELD
1rfS+u9YL0//HhPWE9drF7DId/deO/IVbNVZ5CB09IvMTs7m8mOJ5O0oa8NBaSTQ
KNunU1dU/b27FXMKoZgaQ/brPyLjiVfJ7gYK3T19eoTERoW9uJ0SYHDwNqkQmebl
2QogBdMG4bA9LP2sj0ZHqfCzqWxMgI0HAq8OK7vDe2tGxsUv7haE8bWiodIC5+Qt
hxmc5z1Lqnvnu8n4Cvh9OA7KgvAcBEWQNTMhPqEQ6iFsMYw+QXOuUYKtZEPrf35+
QnQU8OJ5Y+sKcCODNGmK5WFX5txKG55ISw18AZdUx39ddz5Lx1vabSZwD43+c+te
SWX06QMYt+UraJiIj0h6rZogiQOfLlQqdzElPF3W9GcaG3IdyEAlPtiENM+N1f1l
IM51DJlw+BnKawWxFwQCZtjtlbHPaTnEHc49rWgJAsyCLWM+sOjGtSLNrLv/WelT
p/WPpQQdb20tRoR5moGo9qFoaYCDjmNTI/B59XBSoZ5+7G4d4reFNyz4Aj6YyR8j
s8rXgMO/yQm3hnsRoBdboArNEbPe7dLfj/tEMI46U3e/SeJ8k3CLAS2+0/URNKWl
Oaf8+dj1KGgb4reg4UsTc8i00Hq+1v/0K2TREXneOABTctA6SJylrrm2zx5vjn+b
F4t2fQn/vpak06idc0nTNWkY/KuXIMktJIpyLo1ddpBSbMRPqC0pW7pv7c0gslee
3+qvXSFE6Rav9qIOq5kZa0OFQTshO+unxyGBWed3BZEpl/Y9rnvolOYRyDBObnSV
CcffZ5yFcsHumaV2U2uaHKlwqtZzg4gcnPzKILsbCZagTlhM3ZFM6P4cdcM4Pz3t
LiVgnKsU4Pk11wcUrwSDn+kOZ8G7hlOjUZJcZACFnK299VNBKfEKanvLReLCcZvW
MSKB3mkziqDOdtyAsd4x0YST4G/xNKhP5bA8zJXi/dLTFKw49XG3JfGnsc1xSbJB
c6m8kHwBC1XMbPNG3MkPLSNuzbiH89Ii/Bk0deWUFlF7Nsz7UvpMRskBKjage2c9
fiGQRZRLo3qG4K6sp8vEhz0N5NwbNE4ug1xvmGVbX5XRARP0dolXui3JRVlg9T5Q
R1m3/3piUckv9AJqwhZag6R9WhBqLuUUxikCFKEmFS6D1j3YY4ittFbSw/kvWdra
+uy+ecAEPP1Scv2VzpM0RastRBrwADRM1wGUfjNLQRx4P9o+Y1RoF2vynP92GnFQ
Z13uqzVXc7MuAtEcnicNMLFNxE+pRgDoSP6yYotX1jn+K/fNDxoirjab5oOP+m+W
YCRicEGTWEOB6w6ZK9f2LgwQ4NkwSQaGON9gJY6WvAmQpxyXmCQR0dJWeqXDqTOd
kTNGqVxL6zBlNKbhE3TyjseQVEm/uR8lTXeguU4hQbar2SO2o5EQKoIqfw/FvoS4
MZuSbazc1h1cwUJiOxSi92nSTxhpsP8CABdoTyEUFs2g1q1z4jhNUldZiK9SH7tX
NZhwtl93TIXBRGN3b5uIixSaItX4VBfrJSJNjjbyn7IRgjUM0EhWs8F23i2oxIWn
BIKzPouSj3CGOANr8DHlaGXAVn4oXeAVYW+4/AEompzdaFcfTJMVMj1nDiBpXZFz
N3oY6N3WS4Khr1qbV3x0xc13eJLnSohUVEzZdxFDgU4CVCwfBAOZ93Pzhl0DIzr3
nK63ZK330QyDCsuq2Yflzrx6KUAFjneK0wQHODiHs9pJeJOKwaj8F4Ivx6lOfs0N
d6Bw7rN6kgIWqw2eY4J8xi7G2WBxtbNNsVe5c6yG0EWGW6xuwNaViwNlyMGz/+7U
Uy38lr2H9hk70I8zKmvBlG7F2im+9sZ/eVVkLgtWgYLeX26aOfKRkeOIQhnqovjS
Z/3oq1cT9jtyNGP1ZPaMQoFGQvPLIKqKQvos6TVzxDJRCwjZuOFHpfcRJVlHNd6F
ESZuzeygJBJXJ1S6mT1mPR4wzj68FZZCxmqLMt+w0tNvAC97qKTiWI1KzrWya5VA
ZpE2M+CMqWfR/7YGH/NkZGW0vv4Ai56pLJSJAit0X7xUP1B14V9fpp+9MmjSfa/L
d+QeemOUsKrK3pjJLFYoqi91swniGwMcFStjf22l3ib84Nag86P+L+nKKsLJ7z2L
qPcMuyOzBxlPGCHC4hlW1DdtJ5tzPtJgej3PnQVAK0F9bCRN/7OvNrqKlIc3GGH+
oh0TOFPexNhWoonos3asoTmdVkaGr1sRJHdtyuW7r2VrJiY3CTuBkj5+8dxYGxsG
pY3kA3khWdh5vHDWZm3Pr3ASbFdx0XgPw2OZmKDjRKerCWf1cabICKMXCRRhihww
wUBBBe237gp0G1Ead/Ej0wG2UAD67S3FeTHjDGFoRhInLSfTQuNN2Zz3edl52rHd
5v4ygO+zZT+ZRat1M1Zd6zZ9HuURkRViFmYuftpIWdu8EjR/mOplwKewC8A6T0q6
RYhuRWe5j0eqmyjb+72ypapldytYr/K/w98mrZvciaUDFSaqz7bv1G+q1AE4JPk1
g+lEOPz1SAZ5WL0mdk4TC229HQi4f9bBCzZRL4+k+Vj56GlH4qmxx/1nCk9N32ux
4k/Qb9/btfH1IwmlKk5huPKQPRQexiTg+PZBt68L0950kklcVI63/YhfeOXG+oHb
sK1jMSAhX2L1gQ2x3i286A+W1NjndqMy05PUMT0U2z9w1nhWU3i2Z2Mji0JnmLZ6
L5noNmsuecnl6NBBFFQGg+YzOAW1pymn7eTZXRQXqwI5X1wEfqyrknq8TybH0pBd
Egc9Gg3JZ2pC3v5AXRCc5tsRixoztidYm1eRbRftVLtqsSUKTKK0OhZcYuxjyP4v
4tQw8PFEGujYeKvJow41xapM05FALevYYlAiPwK0YzLyeRs0BKO7gcxJco9c2VQ9
rR/qqLnofSz35a5hbvByEJLqL76TAC0Xr3zYPDnIsfuCFh+y3ZTXhy/6qQke9+TU
GDMPZZqiYcv5l9WdrX+Qm8v2YEkvEiqDXMKB1+el1FZa9POBXM1gi5gfLEcnCXm/
V9N1ccQYQCzgGGPA6CLtF4pvo3sthUML9c9sDT4OBsP3uGD92JfjxCv67ZPrH5qa
YzaKBJda1C4q2ECK+DzKb5nRJWUseCr63GQjjDB9vLZIrUn/YtP/gv3XdbXKRHlq
0SBQoxeydOnj2VR2kJpXkqTNY5uAZsJMlpOEvAeYXWSOIx5wXsjMrKXTXFM90bwn
ltwzcuFN4Y6n4P6UmUqf23MbfcQQv/PVtHes67RyGM6xdxxX1UsMNgM9I5+xHzRG
praUarZqwfnxk3PI3i90DRMh4jsjePhuQd6JZZBtW9l5KNHabxJW+FGpfdGXSOU8
6FF8LGzOcWUYnVZ279t0d0OgD6L8Bj2AIax2t99yPwGQKJePap+5uTcytbTIOaDO
Wf4olb8JlyVFS0GDUy3bkHHqAiEv5hlvGOHSdHe5FB19jNXxmreB89VTFlkxdk3R
3Tmv0JsfqEcDHhdp/HflL7BVz+LoAiG0k4kD/icnp28KdL87Hr3dKJB1HLexGgTy
hHnWdC28wweNlOTL1JEjXFWlELePbZC+hmHYL7OFBAkdFIrO9nJxHCT5ubFYYUE1
RRIhYQUYe0t3mxZfHShDj5TpxGXmrfBBWwQKT94rH/4wf9+PUD9nq1ly3W8tlhwl
wjIG5lama7YrlFzT75naBgCTBVnjpZB9J+xMcFS0/Kz4Nh+hyyxCZ1YZXACMlYyn
+itf1RKw/+wx8H6nj0OguELxfRD+ZbOqpL3bB1i0ln7xuEZ8wJ+xmLO2GHTWq7zY
/rCtWhmhHCE3kSRWyLa4flFeA3MGmFA7E0+ZoQkUSmZ4cbd5AQegbTAeyY4FdYUy
XmJzXoRAmuMqTFMzq2hlUINXjj2Ag2v5H92+G3fPGznznJp/5iLsMM+b8RJDH23+
/6ypEPn+vuUlWTIVPF1wq/dtD3SJMisQxLCALBicJtfoO46GbXu1GWwSmMW92dob
2gTKdZgetrusyqnyNSsi0UmRTnY9jkBr9awq7K04W0uDPeH2vPjYEx6enzKEgK6K
4s+id+TdkODFcRXAPomN0OPOoP3pMg77u6SHvL8LzITLwsJmg4oBEIaMdpFXMRCB
flg3f8TAgXDkYktCzQDQXkZCKzYrBZCRgIHNwf/7/FQ7i8HS3KDn8s4rUKqBBp6M
0/ai+usnLuXP5lZIFHLKMW5zBKqAZEIDtm0tssJ4z52DV1iDXGVqfO5M829PMS5T
HGLnITO+sK/vbHuN0+CshUgJfZwVE730vzLPFf8AF3UdVFNceHF6xcAM5UnjFek4
gqs2tZ5Iu+OB8H3Svy6Ri1UpErTIHCFvgTNP//03DDLK6oIzcu0MseZ3k9e5HxlM
vcUpNB/W7OwbkjcwWsrvhZJcEKIsHvTwHx3W/h+tiQcxPadantsYe+M1UTJnMK9I
HUCsYlmBIVi1hUZ9q58NI9CfVyeVWZlkKDoCst8+KkwYAPtFgzUWKu3+xutOFQjC
wtzOfzD97pe9fXQuxanR6s0kxCtcig/ikPnf8DmtOrrfBXHPDH8g/ofw245EkV1P
9wzonsN6sdfFWo1NRnKh+QnLiurlM1AFyx6RiDyuSCbm5kJPDXm9pdyCTN9EkTM+
JF7mWcHHFwn+Pl+jLjjvO+VUppLlO0DER8YX2rHw3nUYogC98/NcsyzTt4Nu46gt
VcnnmgZJLnDwq7WvNIRUIx8HObZG+dPTHrSExVS4ujNnLkH4OnJMJQ7pqt/J8ybX
aptNg385L1R/qB7tgK6X3KHRUqAvsLH3ihemkllLR3KyDvUrmy0KOn6b19J3ektD
3EFIcElEDC14OnRmkSo9Oz2XJ8sQ1AI+aA0mFpRxYr9/Df8J/y0mcZpl8Vjf+cN2
cfwDR8TGk7SNHt0gG2reEIc0SSrKYqNvCsU6zBMBljA=
`protect END_PROTECTED
