`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
swwljLkZuhgeHn7Pbd+7PthVAkHpIXn3heBVqyNiHhHhp8Fs6rMvWvxXLMsmsn7E
XYkJqKlNRfOsRdRTm2wrQxlfgPyJ2oOUOVnViNQ9CkpWp8HwlugHZGoRCMV2drQy
em+cYHX7q+UfGbBhpHfUY4hg5OXhLH1DJ6Fmz0q4gyy1sQy0yHjGu4My9x8oSOUD
rhRdgSO61oFR0fWDlJ3AlW5Vb9t8bLiMJg3Ij8+IE27vB8t5gT8E18gILGMEnX0+
9IJUmqQEE9Ra/iO0h2OJqoAlCwHD+Z7iyhsrxyZXQrH3P9lk6v1LFKunD2lAzFii
N90Uo2OWWJ9cIl0w0Mxlq4ble6mJyb0PODoAgMQcgzeUpArqeNQOjamBOLGKXAVi
8jg2UrF6vNuQtoEcv39WwMShmqQtBo2rhQitOrEVrVVJkCFukw4/jYzLRhu/egxa
GSCSqHU6hah5sBcCHUEdJRFvkwNceZ+AwGGAuQxUEKVwf1sxucRMRIDrGNh+/UL1
sDbauFGT1dTV9XTAf/IG99cQK7UM1mKDnULyfBLEtNGJA0Cuz8GpgUDGarU1tMm8
A485ubXiAvINmEwySWQkFcu35SUJb84ftZfIm+3uOXVEE4X7PAiNjCFWqz8OwM1m
+j9gqq6cSSkjoRNEzDSmoVm3GLyHqz+1y8/coJZC9MkMOq/syszN0Q+jpUZ+Twpt
r6ziKP98PnqmPj/tW0pBezFKf0xK9++redXfIQYV5eJDk9tg5wCO5A77rqkS40xc
7SUZhXpDFRCPpGZvvacdwjFQNtiacU/L5q6UYK7iJl69jhNFsZGwF3nQRjqjGR7o
zYjQy4Asg37p7O5RmmreRQ==
`protect END_PROTECTED
