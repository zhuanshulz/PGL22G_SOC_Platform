`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XKrPQQkebD/AgnDvF9zIfcB4VUBvQOjU1/wJqFJ5NptWNnWfEuReDv+hBOH+xSd1
/oyFlk5xuuBB8kYx4freHcldRTOaGnqrnfGW54FhNBEj0QqrMw7eEu1FXtf247Md
UU4Lu0pXt+ego0+fRizXn7qQGnSBEUlUp8w1dYM8q6TN0VnUyIBdm262/ndhPwTF
1mwMJp15ajBmEYgBlrMa9hn8ZJHU5xu8ThkPCT1bpUoqNXuqXaKPHBCc72z7+ZOz
8pFlii7WDz+p+i0Aqpy6h2GRf5OQF0ctciGMX10S86mFjTxyaJDGAbpZRYKz8LfZ
H5c7ypiW6TJlzB67f0Cj8NKEmROBjt0puN0pPDD9LIHVBg1JFbgCIqMhkY05Rt3E
P69A0BeiU5NEpKBklCEshjmQiXKgTPLomKnV9NAivy5DlyakGcrIJPc6vvIaiN38
4FTspFbobp6TISFog9kr6T5wVGWO2BmgnJzoPi9T6iPSEjpNAj65c367LW2cKSKn
ke4xZCWRUNHRZKfV5ypCy0//EAjb6sr1GL/j5xSb7swnMaRoMhCuFMC2W2LLiffL
11dfiGzM+Wl7Cv1M21lNqw==
`protect END_PROTECTED
