`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mHR6TLGEljUzkhh2KeitdalpON+e4S44czNJYmHnlhgYp3GtyV8nUWk5mq2SXxv7
fTMuwnkExaEN3ri1QiyZjGx0bsMdOKesYVRFCyzudBkZvfppU0F06NGHVpoXE0k9
VJBYmBpl7HQqO3GFKr9wbd7aQDDk0rEyId436OnifJmE4e+LoGvA8P6xHAL2Xlic
Jooj7H8aRBHepcEzxXWDHn6+c6pyNG2H6gH5lXoyd6Mn9iE98xllrYCa7AEuVK7M
ztRrzn/nqhYdUE60L3I7Toz4OPoe0WRWeWUtiJ6ytWxmfn8/aZ7nXlkobX4Knm8E
rrH5kEbywLUwmsAMhtpIkN0IXBNp9IYKliFS63tKvzXo6xekJFMu49frsJlQdn2c
YwEgGIVZGgmE8QknxFWnSwVFzYW+DcRdVloNGhbNG46mfwJwkzKd+m9pPbB9OEYC
`protect END_PROTECTED
