`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vXtXU8c+RdzucPLfwj8sH54JeBhckO3zFQ+C3PQFEQivkAgky8WJbeG8lu44zeku
xUehFpy3zUAPtR28dsKCyc0YVExzhX5Lsd07kMNcpQBucPdRhvSfjG7viYYWREDd
EAhsFFjKIfGbi5Kcg2mLXQJNIfxr9MrsDrAjKLazyRQ18somu01qtOrVzcMtbS0Z
PhBhBVVeyNF0IHkpIcP1pbRWsA6KmUYuqgdqsqOeusIwwCXbiAD3n57HIqcIxZ1p
0D4sXp+dxndcEXwaSb1ae19po2z9xu6vcZQrBvvbdoN55yNdlVDUXBjVjzmgqzgh
Hdgddb2gzlW5ls8go6avscdx9i8NuEVowJdXci1PH6XWbGpDF3HKKxBfj26L1Um5
5jmma2mPPE2g4Seb8pNv26c5yLn42+g8jTH/Hh2An6IASjGM0e7NrC9U5oxLu7dZ
yd29N6J6nJv4GW6zcdk65j1v7TCKEDe25k4DPhKoXwSx8agWW4LuWJS1KSxwGwz2
zqqxmmyZ5RYW+/ktjtAZylgsuELOjxP30nfMW5KtOHBWsqRgjn5tFtjrJb0id9T4
SeK7bFMV2E9ZZIA3t/d4aMHWWSbArdHoxzDAsMJxf1zKALc0aZp3qACTzrwl3/0D
zZJqqrurpLhXbFy5lbp9Gdf4ZlU51+FVtHKvKVzjGhX5GkfC406t/19OB4fpD8xl
T0s1JANgJ6UvKNZwYm78XuEEQkOzdbkJXXnasLicZ3KcI9IRBCta6AyxZiid+Dp3
CjPtcDGGz0X5N5ka7nI55g==
`protect END_PROTECTED
