`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m/dFnov0/agM3MOnetLOZlJ+Nm5YTMq6fd+Csf/VA0hOQSxKZUUbJaeOvozL2kDD
ZLtq0jBhz34iPsqGOIcXiKabe5Rv90ASNykDncUiFA5pJA3qAWiF8qtnZFkPR8hZ
EL8Y+zV8oPy8DR50pb336rKJmSO57SxIR02UbSynZnnCI6ai3HBOzUnEzr2ZmE8M
bYioIKM0Niuj/iVDm2e5ei3hu1Dm2M6xqal+TBYlRQz+hHOLr8S9J6J0g5meIT5J
vDA17wp45VE6i/xoDO6J4G4KEyua0N2DC91W9qhp+SOJ5r3hMI+3SsnuGfYjdTAo
T2HJzfEtn/a7Ljs2z1L/u8nisUj38o/l7FkfZorzlAYjudA7HfsfQumLJV84gjt7
SLPkG/WI1ZuJBn+8GNR1IIdmMA/4x/Ig6BOnPZIyMx9FGiENoNrZWWjabLynM20q
JFLQksuwGTNBTOB4PAVhac/gyApKjb44WVgAi212xzAaOIZ1lKIIA3DOiVf0oELg
SRHY3Ljz+ZgZAbDSQ1u4q8UfvgpEnUuN9R4xmwwRlnuLYLmFaEq4TsH1pz9X6nXv
B2NdKgokQFLwXtG6lGjmXYdNm8AxJGoLG4cvh4St7Jw=
`protect END_PROTECTED
