`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NI3pGM1h0hXUOBcrhEkeQvXBlnTKusqJSpZWZUl0fIYzFmTRCo4/6bQxqy2/tqeQ
HBWoss3Mw1uSyR1cWaVGetz+Gxc0deNVFd/Q6a0kRzxqLXKjkfBQZ4F+pyO3FGKi
tUPbkNz7cy8ISCXMM2jg083Q6ibItMsTYLI575FJX4YpMe2uQdyAInrmRXyTkI+Q
csVO4zTbKYotfDSW2opYjeILRJcCfVlQ09ouN/4Pzmpz2CMkgCLlp+eli5+BSXIU
8g0tUS7bteIY3kCfLUqj+3ysBqa0vK0b0NjeVodM0WSHOOEa1kdmsbQeyLvH4Llc
mTK/EKcFo9iorDzpBwpF1sKIHIgdoTyEsFTaSrgTxx3a8yH0Xvu0G23xmFWXyW5T
DedCkaKbbuGzZObY2l4wl17RGJCAj2VjUels8C7Kp9VBxkemaVlmtQFozXD4Sn4D
098twbbR/s8Dw3R8p7gOMVQgh1rS58OUWweIDoxXh/eiLfI/wf7g+pNdOe2NwRHB
8bLZHVxS0Dah/qExj5HR+dlERLGvgNOTwt5ICcYmloegR3oNPg0OQOtwCe8qwCWX
KmJ3ZIDyevyzxZScY4Z0ocTUUUQ4nyO3CTW8IiN5ld3v4db0y4goAqL2N6zLAhGv
D9a8XUhM3ZR0+fAQmVj6xxbnfDA2/01PIG3zIy/Gu0VOD/8vPr297UzmBqVaJKvq
D6GXrlZyAzmASsonZid5lWDNHHgJQTudd++P2qJ0XgIAinbmaASfsgrihnb+hJUe
vuRfPm/1lQlynjmTxDw7ZwxWkFQbiLRRfC94h6Sck88thaWBhJVx3bxPNJ7LxXuo
CL2ocTzTYRFxZMcLVkeCpjdD3+rEo4C5cj1RPD8/+HlnBvjrTRGoq7sLwo/nVGft
BPUCXSDMvlFMak1+EvFyoEzJlzZKtNkG+tRDlTyPM84XlsQwh4DMa+0OmsJGKC0c
pVtSD7HjjRy9jpIRqR8EL7dW4uuoju2fjtJ0aLtRLIWZr7gRwOk0ykd+0co/0ycN
TayuTZPBsdQH4Kekc+0Iwb9FCXLIlEVoFXUY2S+8klq/QzEG8v4+j6kfevy+SJzk
iUjAOsXd6tiW2WltOY3AgniRotOxVOzCoNZj16r5z4k8faUAebxgJFf+bKhxlV97
rZtG5Y50SqXF1Wfp6ysYaOgl7kOesc9u+1aC9PaUlOnZbmk6Wqo7ZOKezcxHANx5
Enr0rm2CYB4axCkNIJanhxBuTfTKy4n46an9RJMnUgsB5fzG+LwuJtSCzSbLmO2Z
eSdLsvKsDiKruyoIvuFj83CDa8EJux5V+tQrbQbDnk+pKLYNHQb/WPQ2z7+3/UoV
YPX+u6zy1k58isrbTEie1CueBIOCkiLxBuoe935S/YS6lBGWBbJJNCLPDU/Rj9Ta
d7QHygg2d4XJba5e5LqRpdG9gtd/FPecKSuc+glxHWz391jQrdOQ6P68/qjhjRK9
9MzxmSEJ1qjqzwvo+qiQUUVZSnjPkJFCzPYXciPHtlHQmjyf1Qdu0EJacw0pGsiv
rLAgCjpNPc9ag+8wStt1UwpZE6qEYyzqfmWuNB1vAbLK5e9eWoPcrisPtuemWoVY
wjaY72ESBPlqet3nfEf9/7uih5KWbGhTB+LC21VpivORezCcVsg0UTGbwkcuD5O8
nhixhURolnjH0xifzANq4XPPncjzGOtsCz74m38PXQUClJDFvY4HQkHpf7bcdXND
yRzQ2csYB3zilTzvNXuptJakniFa83P66AcYhr9jWHjQrIRkJToU2OTqcd8dpufS
Fc75qTMU/1OaqNyMkZsTx9A+8aUY7c5p7EslekflAMqiJQH9foRUZNBhO3urha2t
jlURJbj3sDH3BWBeNgezr3XYtv2b1zEdcoWQ/EqfHPtQHMiRInAMWRCABIgf8/3Y
+WvVK5+7HvZUntV6or8BjLTRt0+w3by+5aZSFUH0O8TV+aTuSusI94pHtfPpNV8o
TE33O1Gq2OB5XZSlMWkOHkmqhTtgHrk1kbFE9aToycjUUX8DJJTPX4/wgDaseKqL
8UaxeurAjRbBq6GJNJb3AnEmL6WnGeEZpb6fMcqyWbbLVCNwsQEMYZCtK0BmGI9l
euhXbFYHqyL6eyoqClweo7N1ir8FU63K4bItGYp+HTY=
`protect END_PROTECTED
