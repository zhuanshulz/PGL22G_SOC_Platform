`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PhSkKh4KHq44YzTpyYtJGFT2aApNHTGK+ePEh7d9oSveTpT43SjKuBXjApIwWkuO
D7/6rgudvSQiBtnxEAejG0+WzndkCV0TBElfwFWYWJeDnWpAHKNX+CrTPOvJQMpi
olpVB34yYtAVUfsPEudObXw2CTnrwjC7mJ1+DyPa0eYzcs9Xk07pJVeBPjnoVpDb
iW227i4+U6QyZ5rdeSkT+vjc8LsP9pEPnZQs89RGCLfQs5M/m7U0IX/klKNmIh7D
YbwGxPlTPKB/+XqAnfoJisy5C9VrAik0K7Y+R0Wan+tep1vZKFgF7hkMfe7pfsFZ
AsERXl63GGZq+FMh67puqd55msGrq4QhrJgB880w+9V8ZMe2quc17WqtZE58ywFM
UMeij64MzPOh49JAYwxutQ==
`protect END_PROTECTED
