`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xs0cMWrpzt+fC5a2/rCbPEJjRBmCPqjlv/0Oy/2KjrUAnvTL9R9ACHDc8jaksBls
4ZFwqogtuisM61qM80/hp6KHhCGvA2spnpaQ2paF+NdwR+WEpq1Xyjr7t1xubZRQ
gtfSnHD3o7gyARIiif775f/AsZRebJqaNsX+gg8zj0XxP0oLaYK0Fdj4pMNGcZO+
IaG5mzFUbl4R173lzE3l1EJG1bacY/Wox1mcgvN3uSKtkpSI8CJS4UTz0jGTcnlS
wdi1TMVFAkXv2iF+Q38FwNaUPk2UHFXPOuEpnebyHoqlNbFmWkp21DDXVWsRTnml
nZdqLIbePLVYjnCORUXqySSdonavKeFxxSInUAseQtBE7umQaAAquH5aMiUOtJA0
Q8o9SmbRrF9xL2QAE3GoZewVUmQaTbawodu7vHRnwW+3hVjXSsjceNv8tcANoAII
90pJ1JYBP9I3B7G/8ThKINOEUBgoM/YsGyJFjbqalbltjfCbL//SVR2dPcuhg1Bl
PQM4RvEP9M0STRdKX0HlHiL0qZbseAX8yNwDEt/GuDqaI+Gb97S1dQB8BTLnjfAw
D/YyUf2/VTdDZOYjonHcFlBj+BUbobMjV0AJ09gID4iGJLePdSq3mpUDkSuD0T2A
IC+mnzRPLxGq3HtdKML5aTLq/nLOGEfIyCNz0+/w7LM=
`protect END_PROTECTED
