`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MmgpsJBq8B+6p+fGMTRlc4thLpNeWb5rOuQ/vaCPG6RMy4aoGSNWLIHI3NcOtWEb
Qz6xWIZyy0Je2ct8ZdsO6YjrwbVgxZTdlo72N2RpNGLh7/Ao8Uvl83HeImllnGkZ
NbRTaUJ+OgyaTHnlPJGQ8laaX+9yVXzqzYvqGh7uMtz99lnyV3pl41R5AYPNRhJ0
I4BDYhInx4fTJcd4fIAXFaAjlH+TyYERtNw3dR4Wj7vZeRAjyokDwZnXE0B64oCM
rRyM0Qm6+aS8Is1WkUMnqVKUFTidrd+8bdJL5uO8IWs7Zu36ng/qiZSCPvgztLjg
`protect END_PROTECTED
