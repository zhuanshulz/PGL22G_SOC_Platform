`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zPGTpJbgxOc8bbpJ4qhB7ULQp1hO1+gZqvf+4lTMCHpB3I3alZUL/Me5XkO+cOhp
4hIX1m1Va5lTafEXVQYj+TICNHLXSpK1wRBfJgkQBXZ29Fgqtj9fwUftvbozybvj
xx3zoSsX3Ajv83/TMeOoUSE3VRTaGbZmvPJHjMFKAVFP7k6wcguTPGux3csmy8pV
sNlw5S8r/2uWSp+TgaZoviHaXyoMwK9yOnuELXmsDKk229JC1aN7binRjNuAiHyI
wDvxRY2gXcC1G9r6sJz9F7Aj9qaNUZ2TvRPRerF9/JVmzdKNsUFSBHCEOfPB0Lzi
xM0Ao5nqdA1OGXU7Low36ckzbKtqJKMMcSkhxKj3SAeD+vXSwRDsYvruI1cTws6s
d2DEtiRkx9SwUVd9AvsU/55yCJueMmEZhFREFZnBbppiZlec2BU7J2waFGgZfcDJ
ENpFr3C+Tjb7giVbIEsrUZCrfDrFIqAsdA7bJSPDIqrg2IzgHWM08X0zIl/2mNDy
WJQ3YJ28qdcH3viaXpvCD8XU4eQSsEbsuk2F29Y3o/NjT8sbtQHfEBra7A0nX6Tw
UoSpGHOK89UQ3b0pRaI0DtdiywdzBgH/mc4R9cH9qmRyQjm9WbmmGPwhzWCOhOlO
143A9B7viXDYX/G/KzC4ZgXBX1Nrl66OBrjDaEP6IdAV4sk2+dfII0mkUpx8zsof
ESjYgEHiajm5QyxD4YTXdvoa+yjJ+dLmSxkvAY9N8lkJTYxpj3Zvw+zxI7AC0Mx3
7fZGr0DusAIORT6hqxa2Gwgdtdhkjr5lxBZ5doy9pfB4M7RFU231NSlkhvBC7fHc
P3XQQrn5tiMFa+BvCDooQAisPggG2v0u4QrYAOaaiLOQ72Vq1q52vB61X95PeG2J
yAiqX0b62NTgYq5tt6k3WH+wdmIEv9ytvx4rCGbCllao9oB6exedNtWxhNZKQwk5
sJK03mlUKlawV+c3VCLxvYaClaL1s5GwiJvpoksIoEMoi6gQGthYWuyhNWtUcinZ
870mQVOE5n0s3f99xsqlH83wN/f/upICQVgDJRA2X+Kukbx6xgFkIPJNS8WOSMPs
gIFkRQPYBAQyJWi1k9s+ya+Irh+Drn4Cb1eAf7VoxGOo4+YyhUphr9SHJpwVtvXz
s6N92B9xrVkvcecgiZqPucykflCmBusdoWZ82ck7rJ6DQ7Wmun0eZCjXG2B720kN
ConUijKhkI9n8sCodshP7gNuw57+SOz+o+020RPfheqjB2KUwgi2P0Zc6cs74Y4A
jAoSOZPq57zjwTakZx+vKjD/wOXIPpXby0q6Q6rFrQMbULwzohET5+5EfILu2IZV
`protect END_PROTECTED
