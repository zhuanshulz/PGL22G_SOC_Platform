`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x+RUGfLPtr0yyNtA0Dyt91U41Bz1TqUIIckTJTN0H/1HyqW+rvAcw1z2U3ukYKG3
88NyGI6KG9AeAreGiyek2hSEvK8SdETL9PTtD1dUGRGTGirR+pg7EkqteoZjOq+9
WT4cIFWPqbsGgOiFeom8+a9qlDwp+svriJUhEPNoLz26fY2kDe9bWweYuWB03Gfr
lxlVx3154DiGyLYi0wMzDjtx9nMNgW4Ue2+fiD3/yYmZorepGUqbh0KqhHydXvKo
0fQVijan60TMrsReCV/8G5WjzeWoepkdDMenhDpPVO286D8H3d0G0dvnXjtdIbxK
PQN2nU53waHCZhEDSTHXgDp0aSxc0iCgE9THY+mn2B13MtjA2gfEIQywfp5SrcQi
QpfghX/1PfohxzOLI6cJFuKyUqRd1dTiSqX5Lg0vJNQIRUIFsdZtDsFxU0492E3i
Jmb2NG9lRgmH1r+8R8gU5QWRWdgndSQzmRIvY9XdIWukiPcRUiZbC16ODYvj2uWg
szQKQo8y8Spm7Hwvv6dxpXEH4IaGsena2SCwfZg3qD8L8WDg0nQufTHuGnZWBt2B
xzETdIdTjc1JbQCP3oGnxSJU4glu3YMzK51dDFJhEoj6rN5I3YcCDNYA8kzQylnO
8NJBs8sZ4KiOtABiMpWMBAe5oNc0fBIxZdMViKfgbtf+vNcrm5NcMsJdYDjB5zg+
zc335wc8YYqTEjN40m1ihYTPfMRd6pcnMtuwxnSpHiWsSVwQLYPOnKM8b3xthVT/
pdiTBLKTSeymS0lmagFhB2ECX2NYQ3Dtc2fi7OFVvAgaxzKYSZHiG+5bbz4hxBFg
EldufN3xDWFcKmhe0mTaVTgxW/l9tFI874kZnbhgpqEUaBzc4zEX8vj9YLtjjjFy
hgtv1RTCgkH0Y3uoDyOMCPTfB/v3rZ1oj/n2z5nQJHrgW0fwL6qjyHMqT3QBLYBw
R5xabROgHpW/tEoPndMeHiQ9PQzTNWmqjA50bdGle1TS/yoj39e7s+pxmwdgT9nS
GafSbzJHbjZuNj4Jmwu/68LmHCpgPPFpYCG+7FK2yXOTsO0dRuNaJbI3WhJrc50w
UqenPUPIEPatOmmiBOyrcgpxKaAdRscRUpIDU5TGEgf1fuG57NX/DMctQJYsj2by
jkHYjRtV1HuodzOIBdHrNxwFCoj9M7DGvz0cEVTR1Dsp0dOE7TjVU90CzNENzJ4S
IMoTDO50b2aMUc6ScxLgF+VgUdDYPk4cieKeBnBQZExemApzwX1IgW3ogUzFc361
rUrNMuilAVBcKGsuKoabSNqZsV4ZeajHdehcM3xVgrB1Q0+o/xBXyHiY1XiQ9t1M
J1b5E0+L8u18yM6QLeDSEEtvVsUy6wRUkp7g5oqYnxZuKvUVRsl0+HM3/GZePgwJ
7NdOgbaes2laxKeaO8bBkJf04mwuW59WzX1WKiosF4YAO1O8/Df7WPXA2noqet4h
0+Rf1dh99tyDWob5XGFaheAK8ry/QTYHdC2IrLTA+UNtwxjiNNbxLrPmWrGyMA0r
xwn/kK7KwT6UowFJrkM29DDOk/wSJTTuks8dcz7c5TFQG1XVFxFGmATxWJl2yjXH
MOX7b7qq49jEuFC7MXoVnemM9GtnMtUMcu8LWV/ORCLV8KRhNWSUoy5vGWhHDzrU
8WKyz+wrchhG6bIprUIBURiW0a2HecQg/H04Mn6oObWEHj6HADfe+xSIJO3OtMmf
AibpMTKa2j4p/+FxrjXvtpLslTeJeenHH3BcUACY9cW38lYhV5J+1tQpfLIowMbm
3IpQlI9aalcXoB7xdS8ZgQnu3SnGCiXaZpP6C4arVKn3r2S9kXlziwm5MmiSajuO
mZau291OwIHKhDUQd88UjKXXbpCDY703PrD5lMzocv5bYu1JaSfQRdfTE7vzYPPp
A8yQwKfFcZ34nftW9n4gTrCL7AZKfappe8/WZ3hz/6uz3CoSvZOQe6JXGuJ8fZQJ
zlP+SJKywHKKrkQ88v8zaVYhwsFlkoiGtO6rbg+uKEjg0dn0QckyiBWOherVF02n
fqmntIca56Dw5fcUuyXh87xI6IG8TPR0uI0PIGrqAdgWmuYIB55zKCca+arBE6mn
1gnWPQr/ddh+dwfE6VnHLFfI7yPpp6eRwlcd5mXenEmDwacJbHVQ+9Qi2/VsVqk1
4JYS1hpgfcetS0Q006cD/gHygdeRoUH5kHh/A8+toxTrEK7dgUpkiWXTxtSNAyJD
16ot6W+yssa6vzDQXROhKLJgUi9Bw6f7WNwbG3eML09keZnw03JLgCAdonYjpBOe
gdHP1W7Eyn+vEcO4yUZpKuUtRrOXhmFZfmjux3P48rnBAYhu8IBM3B/S4iSfbVjI
G0be1CN6EjnTzAnMCwzf/deHGNuwATyStbDvL5273lSvpwQicycscwH+piL+6HPv
4/lQH+yJWrYEuHsZrxfArnz7XurRWI3flC3nLUqF6+Jt8q/0HI9iYR7MuMe9RXwB
ndey1CZuMkdusmnhKeiAfDeRV81Hd2ZU7a5NE5REjiRQaji8pzX0gYlzYIOgr1Q2
eF6HgPEx8JMp1TaPM9G8Bbn42eUMJqtjisJyCmdA32nz8s18zqcTvLqUllnH7DVN
0seSeVU1a53+mAoCcw+A6o37CDUN06dZ6J1sxVQZw2ZXGWmfv07SoAXkAzR6/u4h
gde4ziz4dGSOWIEnfWukvd1oSvTFjIPH4SX0TEGOfm/25GUfnqjuXv4Dim3Wb9Im
ExFlZOepqgMtsRzFurmHj3u1934T43Cn5Ks0Yb+YdrexSA15y6q0CUdZhGux+U0X
24LJQkYlJRaJzG0al/1NoZGgr6zTj3S4kHtN4Y7/7watRWCwWhMI+Xc+D4rYyqeJ
hPWChleh0DYb6UOmBcZLW48uWIh0N4WsInIm0ewWuqG3trdJR5onclMUg78cYjGp
Qfi6DtoKkT+znKvL4+XxsMg73Q5HWR/g0NDfuargiw24nS+EyNLHZbx7XuMHWrV8
ouw15HKFfwH7jLedcwpmhZMC2DQgt2UjrPXbF9bzZZGIsKXPuunBu/vN9FkJN9CJ
tLv46EhfXKDP8MULysx14EDh0rUoxd4PjMVXQTt00V+Hn1uxJrg3mmr1GklG+rF9
fi6ix+u6PDk90CP+dRBrJXkftXi+OC9t6zWRpi6oOz0cZysDXyvq4GQ8vG7BPRTs
6/FDsLjarykiOAWkAniHvfn8JaxWlG5EuamiUZvYG0K90FEcadnEX6+vWVAUrP47
HgepqawYj13JiuhSfa6EWdkGamAzyp8HKR/ak8N9m/+2bRcFD+gU/BSPk+g681mP
eT7Bm0F2AJ3ohOghoWQ/PLiiP1QHeREzGz1rhrezFYfluCb8aQMayUWqs79t6E71
5utzE1Wsl1WQwqLPPWJ3ax1gFgf4V+RJmo8Ch3lrEkr9jn1OQrEbNSA8yHvnxjOb
z1aib01gB/3oCs4hVBUFRXTfnXT7k2ICgOoQdpwQixEUl2w3DUEJCbvqjUJIA6Iz
vSEfu9iQGgt+ZP+QjX1k4HxQSqeW14NP5ahUusL+ZyfndAfCvpuawoRbk6CfXODl
rYHXtAzV5s/+USAnfABAB6trCNGJG3shRe5FR+aEc026P5+Wvj2TE/WnVN5Du376
D3l13u5TN4k6lLVYy+jx9MEenal5RXLnxGafFVnxAHSmwfqQXQ/9A4QZ1RIRJfH5
h7nAdSrXM8fnF61IltXrt3WA0u6hjG5mfDnkF1QcJnL06OubVFAPnC9g/vxrE+hw
izMzSq2C+H0R8S5MlTeQsDihGp+bK/LDEwPdUiw4NeQocl0zVXdJ8UhajUAu15QE
enMgzS8J8ACt13GdHv4RUu/JBwWMljuQWXnPtzORzcAUJaYvS3jvFx4O1XFoekvd
YDwvD2yUp5iOyb+4S/EjB3wb9TmGZGujtJooHtVr3zFzgPRmM81kPVT9W90FVepk
si8DqlN3uF9UdajJyEETQKfFBR/fpWymDcyFQ63Hsglk6w2QFDjmUyYBUryubg+M
rEw22BrdxVF1Ti6dgStbQk7UOxUWd32NIwQ/IVNsmH84MZuQwph5PR36ZlIZEUcS
dj4T0HYA8s0LGcsgcTTCl/hPUK/2aZ/SCPKUV2xW+KzKK6g647XxWufntXHj/KLF
zwN+yjtm+bHVIid49i5DsswtsdfkKAvNIPoTe7gK3f9MJKEMcbTwHiZaKrq/E87/
mCyR/F+NSCrdZf1tNyIOxafwd9lBaAkSrGTZCYe1bv2RON9t/S5e3QX9vVWeKHIk
qjPPwRFDE/Yjb4LEoWTswEvSWPLnLJ/BlAEjqdcgf7pXGpgadclOvdlk/rNnuyVH
T5wHjttQsiWZDKd/c+XUhhYYXxrRkZh4atYGfWKhOKrkS38Bf93kTJJPedrVym89
hWhLuUAu+OasRiHgC8eLWKJd0sExwv8XdE1Ei3HS+P6AO6aMCW+Rs/xVbG5KmjV9
Oty2F38cx6Rh1ryO8GYWW9gye+fCBFXq+j1T8W7EPdGg34WqcCe7XeEtg4IEyBPI
DvxoZ9YsIvdfCvnKfMr3C3JTGO3SVJS5RVh6qJEYYLT9Ri0nDdwecw5jte6xskFj
PqDFbdJcDe2kux5ugpCbEyXI0RcgrudWHtEpxyN8JAqYdjKxM5xH/IHrpltA3hbZ
AuAYapWUW3SPhMoINMfaYO6wrdSLuoKjP73AsWAf1RAAZsuyjon0eKXLrQPNb5vS
zF7v1Gbq5q/fwyU8Obq1KFoZftNmvc8XRAuC1Xs03BAo/g6uEzinar4FiPD7H/XW
w6qbZzxwxksx1i5wTKdofEluYPOXLj1VAYRiOF8UAxKHCDmZMotnR9M+Tq0TSQne
Kcq4cNPJONOIVzSFZ0195qzy81fZo7Jq41YjCIiX9ZMhJMN6nrcjMAMlfL+bhFKp
lmqq9fQBmiFwXVNIHL69jrGV8qhr3vuhfmfgria9TOb7FuHKMNzhXLIDaBL93yyg
nmWwTPoS4g8/UlkZnDIlLKBeaSwdkErLoeIENB84zRp9mAM0igcJr5Aj3LPmzhcU
KsarLmDH2G+nyhlsZVFmrDm8Ei+BxsAvD9kNFQ/ZybxeqPfBlE+KrWwiE1FIR6+2
uXUox5RJABvEcNzl3pa4xKu7igGoJWAlu90UFi8t0aMU2XrPQ36QpTAqHcWy5zDD
f3yz4bLl7HasSyd2Ra3afpa+qcSCz128m2KrqRzp8mwcSpjnaY0qghHvxj0rXwNe
3A+F+K3upXDlkLJ/YglhzWaG/GcaapfeWTPSLn7qYTGWF4zCDj2uT6PXqYu+d5YA
CeZYjgDs1So1JEOgTW+Sj5TzbffoXjgDpfSyRXiQJnTpQ64PG66E4EsIQaYOg61r
28DNPGO5aTR3eGrzGqb4xspGsA65K/nTA+B/4GQxQssc5pMWAvZhuOKnOjWxhAEy
O5f45hs4btxgumbxhzm/IeZ0ONrZ6z3iDbANSytjngn1HQxL8hI89+mlYMGoqjhI
GLJ199frrNm3y86hYMZY9+m94dPMm/JFpNgrVZjM/hDbBu3k/hPl2uVJKKClQOEV
6EinDBg3r+wWZC7pL0Tx4YlXSfffmzQHDMsqT5ucEcxXh6wfaANfsnqMAiPjaq9q
6VEkG+/1MdIfSjRQ3ezWJ1a520ndP5Nf+ZQbZjYGZX5zZ19YDDwaUDTPw/nzShr1
ZUG47WCkEJmR0mnA3Wda808r3Tna3BPXptSICovy7JPLW3Tqouumji/Bn0h71JZP
JUkNvnEFBbIYGam2ZOFUvvonPMuX+vRkmV/wTFShFytlBVf02n2k3t2rrPJyhF2u
/pVfHC+Q8T86AtHGm/E5Ai/m5Z9C9zpJINtlfNHwSKeXY5pZJUpXvp5D2lqR45+L
PSXATeIzrUbCBOowM8k2xxGDHzRNzMJIMVOxbQn9IVBAhO44Vfwy29dgZvT68PLu
P7XOtTFKg2Zj9YQ8XPCr0O9PR21E9jOffMT3c4lIr+C8qX9KIf4Kp6L4JAqI3ndG
wfF66lRHdjuMqHwfJJ/c9bM0rCWay2NDthnzzukzGCy2cBayO86rlS+Ti6d+Q+3d
Lfd5P1ZCuiMFkHQHDftmVakFqSrOAmcol90SOAr6qDWLu00ZTrnIkRbriQLZJGxZ
X5xMjZIGZHPoDvfuvxgYXeZb4krLZjB5dtaHXpKTxO4EcfFw5BbpNpecbZjSLzpp
eq8uYCMi/o2PXqsmbfqZ9rgCUOaD+D9cBByUX427PK9A5LleBeH8CgD6vrkG1B6G
hoVwxGpmx31ezQ+jEtf9z1Y0w1iw0n+mr2BTGr8O9WMhQOtWWxVKxn10f+uEIc/Z
8jeWQ9XYUDcEX3mfnXUAisNt2YckHbajOGxDUr50KbP6ERvkmPeUL6CrT1NEhp1W
V3fyA1OztTOo1QZxJk/K+ozes8uPiZXs5hPY/51REFO8bxo4olc+Pfx9oqUblt0R
Efto6ELPLmK7budTEApx5yZTMM2d37whHldnJlFjzLnbKaw07+mmOIDMlPrDzFL5
sp7En2PS500KtF0A6PvI0gZzU0v5LQSblAIgJFsuZzqkcKSnMsXyP0COh+2MBc09
6MkaLoTV9CfuHmLyStFVuMmXXHTgW0y9ISNEEjdImZp2it5tZcW+dlVVIUuFRZof
TcPpyvMrvOxZPUBjoKRZ8ruRbZy3+hc/fxA7aEUNljeW1spbNCIbrUTS7kAr8nAs
SAFco6X3pYlGnqcn68N3nxPZ9W0PJnr/yR29YxxIkdX/TdhQIXeMDWW/hboa6LxB
7qSGd8Nim1hDV+jNgx7ME/sSrV6OYRtU2hylE59l+A0QHegn+MUq1q2/SpYUY2YG
3TrJGlb79h4B+cXHwBtDrfCVyqNNSQtSy94QHWvjDHufa1023JgLqRBB5E2XwMvc
Tngg8b4bbV1Jloce102Q2vQl7om6f3cphOBtJ44sAXHA4YWger3Gvdvz67ibYg1G
k0wIG2VTBqmATmy22d9sLfzP1eFZ20TOJWcXpewUdgBX/BzVymiD129bbhJ6q1sX
s7NIRbnfx6/YRVMeDf6eq6vIP1ULvkkrbI0vRcmaCTgkw1IwsuXs9tqrAFeZzMSd
ZeQeC9T2A0RFui1SflbXN94GdeAbENi4SN5OLNqpSApGgjOug5brbEMtyKP2NgBo
kZ/YZKw0ID9H5n471szWLibGtgYUBoIHL0eyAi4ziPSzlybP8Pcdx8ejG2BT/o5t
LcCF/HGCh9T8UO3MyLx1BnbeAy/74RX6Zh5O1Hy+/Hz/I6w6NzSs3bOiLmyKq1I/
sQ37jxb6ppyrbF0Rf6fODD8tShg0/sNyl7ZdOX9drmlv2kAqW23LD9sq6QNwxiet
V+LarHPeh3dYBKFp8H0pV8rkOUdvquh31LRTlyjP94ROFDnLxFRh6V7GfGmwugG3
v3f+H8fkJT54EbRu24n0Tt8Xvl+pYyAOWOARUE4Kvkkris1OqtUt1j0Oy0hEtpz/
5Xq48NlYWEbm8M9VjLVMqNaUJ9/x3iaSRfB6ZgSeOjv0t0KdIGziPv61jPU+/HDm
5bZGvtciWDJ0xRnDGo4SveQi8PKhPzUJa600dVarefbLheuD1y1A5U6b7adtbDRM
SoEGwAZxqJ/L9UmSApsP/iGV9DuizNDTylZeqD/RRJbIuDO7JV/R5IS3SD7MEKRH
R9RwpzSaWn0TZs3vKIgSTbGrSReEqw2KH9t/60U+bV4yGmvaWrxVxeaBbznCFQdV
ZmU+GenxUKKq46B1eqdc8YEtsbBkMeuiVD3AuWVpua0OqcSIsttCqTi6rGIV/yua
AOnjV9LfGr6OqJ6K2eJiimFnd4Exo5113RgqOu4cVMHq0O20eEcLir6QRTY1UvOG
wcRoKqPzijUC0wYPQwAvwrqo6/BRzcmOL4i5rdM12QobNqdf/sWpfzQpFsjcaES3
D/bt33UB0QU8MtUk12ASsFqruahDttR+GdZdzOxU7dZY7uuLlW3Nljx7eZORRa5x
FstIxQ+gLG4YNYV8xTyKIcSAyCNERmcs31jD3adp6dZ9PefIWpWER+RcdHiTMuQa
9izrCfUFT26tqgw/VJIxZ9we3l1igFZ/iHWhu6dU0wyPA1g/wi0bqsgv5x6U+lF3
RWeQEWyynYNfi8KHXHMs5i8gFiL7P6yzKA++lznhvGiRUjKMCsdZDUOfB1rIEWu5
XwD6vLrX473T0lJFmwd3l9Ici3FzvfSy5QN3WQ4/Qb4xKDLA23BU1PGr9rupuSCZ
r4vCEXMPzy0ZOFh9RoLsxnKHfn22NhWA4AzmrzbFt6DDKvactyXTy/tYzrrMrts1
zgXavif2CrgpAU00pKfCfd7UaTpHdblRVA2gAz7tv0u1BK5xayJAs7cVKsPZTPFR
ab4Ml5ikCXfQTeOKuc2CtGEd+HvOmNrWD2AMUpDPYwpNBlY6C+VKsbe7JaKFsIeB
RVFxG2kimoO5ESR3YZQGZULGA7xU0QmsJuRlqtSuRY8pnksFPijneaMOBlQMpmO6
qzvGJBqhO490IRKYcFraQ9RpnD/wG9EuSK2HfpvZE8godhW3LqbcjYlvMHIjZUVV
6INkr8759agAAFkFRdBJHPe7KOMywLqtY9n9fG+W1dd2kHhQMIMHql6LZk4WMu2L
+u6rfXCt3S2X7ajsKRJBlgp8+yW4p/pS/aybrqbhly61TgD6URe47FAO6M8HSZ8K
ZVtTAMx62NCrZPvXlEonofI/Fo3Qsr6U714T6iTLYfYxhhG2i5nKIyaOs5fgoUnh
9lZHUxD3bStz9uxFekg1R3KCUHWWlOyLXKcP7I4Jr/OBMTAVMxIbVIiaMjoIzYll
4dhVLbI07zpDbNwP5B6Bt/d06NgCc1si4DmC0AAD6zPz8O7mrGZy1PAeSfrujvwz
Ovv5oslr/1cL8kUrtGZAo/lcl0pwU5TNQzm8/OuTfv9gPN+0e1//SLmbsLDfhCZi
tQE0Ubr7iuCVe3YBjY3qQl3NbuVs+V84i1TMBxc50LjdG7fvMC1H/n9u9a3SiSKN
w61MsD77mCJ83V0ncorhWuCnZjCyecRurcx8Nxu2/+sdt8Rss7rGt01xwJeggLQb
fENzK+H3stQWgrhTG0dkNCOexTfG2qBieJ17JwfO2pQlXANExN1PDKxLOHmKkzM3
LPuEpBNmfkXUq/JgVs4vcUWM5VaK152k6rLxCzYQco+hH8ueFcphQin79OYIAIIE
J0vgLE7ofaA9XyvZVrPVoDcn4dNkVPoqoyg9eZLaCUyNAnj8ugDd+SJRColJarsZ
QBPBOicFGpiwDVissIpgRcQOI0ZZTZkOV7Sw66ZAES9bvUgPXV8wDSvb+yvrKbra
hhw/D157ksU+Pks6weXkHCrNNaF3j4zPjcn9DWzx07MR6AkfArsEaE/Nup98+tac
8XOBc5JZUDgWqT3J8Xawdgdm1G9TAztJzUGkvMEON1SQmbBfIrul/ffpNVpAqYm2
LGBquweWxuqlLGk/T5ip4Hgeql6Zewt6Zka+t7xwjsZyYiaFkWcDGN3eJo71/0x+
metLqTLFSoE8P2FnKfiE/eN5bjtrigxQ2536QGveuHWO88RQGh0omfycJKWz2hnf
WvRyJw/TP+nH1dN5vpUMog9TMi1nK12M563jsBhYFNsbc6UPyvEDu4jFHij0Vd3O
5WYjiRXpLBUhTgyeqZ7IuCX3opvC9iX3wEjn/4LcZoqVIYpo4IMHOZincU7BzPZn
RaDacqdW8htyFR3GGuBNMCWuMtjiecXO4n3JskaBUX+l8aLgg+wq0lx+7JsdlEuX
t+mAJn/RGHrgh4eJz+j8sinJV3hgXoJ67+fGHL9m77VJlA+VKstExvJs2e5rLn5t
sBPdSrQpQ+29gQJIr7ASBanq4XNDQ85Yhzl78+4RlI6P2/tTViGJJSpAP5KxWMGs
oppfIhxjBQmnNK6o0LaOnj7M4lGJV7IQb0lqMohAovfB7JoqR65M3n8UC87weYUi
EQmsLpIZ5xECWSryVyK5G03TH1khVZ3AjM9dULTpZqCsWNFXH4lge5SnI5DMgdVR
reSUQ35NrO4w7LUVZo9NONJvUtU4RJKryJ1UEKU17EiYbKoTS0BkMuxUHE+0U8vm
cUpQJiypYuWh4sTNRXWom56e66VCyMwOKPYKmgWbF6cNtrv60boRKfZ9p2SuhC5H
BZnVDSkHto03vE9XsnA8Fb2tO2s8xARQU7YKMmT5w6fUe/7zIDK7i+HU5I3wJe3L
B5JX3NZFsdPy7FXNQQJBGA+S53JHtLwXnJhsWrjpxfXQ0TAA+nSCeDVWeJ3i/5HD
LXxGYbc+obe2DZfaHm76DppKjjQW0pXCXWRAv0FdH4ejJONXmA+ObRofb7JF8EcU
kL66OZf8HEEuVZcGo7u8iBTRPey/fRGv0wCILxLufiC5ftClfSyBMTsW8iRTRJFa
UlROSw6RWgOMSnLbeh4iPHGhp7wEfoLUyAV0MI3YeOUFIzk6vPfSpoODYXBW22yk
1hK3jWzRnHnZg0P5zYReFOnslnzfNvcFK1YaXx+xrrPzxMh7Hfc8Cxou8YV2k3QG
ShU0JOfXjAngHk3jjhyMOKFpIW7dj5OVrgnI5eVLe/HR79zWxn7QpNv6S6IHp+aJ
`protect END_PROTECTED
