`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sbvLYBgJV6zEQjhObLOlkOeJIpMFkz5EqLOjIOe9sEuJxkw8Gk8oL3J9NabsBySE
Y+S87AMv+vRel/WfBqu1qw5vp+i61cYRAimqOFY+0PsMwM+1MHkStmE/mUW0fe4Q
FrITpV2A0jUcceUfR8qjXwMznULk2iWqUrAhR0El96PV1ReiAkOghssrzfhC2hs6
xIbFJxnIngWLb+uJfOitJ4Tb2ciOTAlxHP3bRfQpNcwduboqvdJbe4h6ocEYbCQG
MW5RKR1NWhJx5hpgdFWf4I1ladcwem0nv3Q1sjMW6AWa9VAeqFtIItp0ZHtOAZoP
OC/7uIkyT/l/oLvw8YhnTntEiVjMGpRD55bUush03aqybLMNZLtY02vgaVpyPOQx
O+XHsZDt+v7xjJudVmQdBwZysQ+AtSOZ/IunTdje2VAZHZLZYJ2MCMIjDLSoHWRr
WhNoPh+swasTln3qpRpY2ZrxJ6ORoPHe5+s/CVeqHEYIIsSIv1zXJZE7C3sBbNLQ
zzB2iBRzQ4Lpf7LvU9xxq/w/p1tKMT0MtW+6RCOi+t8eHlY2/POBw2OEskyXEZiE
mSkj2dhjtn9xwVsDLOeI4L83fCcsG0jtiN9AgjwRD2fqs8dvaXsDbw2l91C4PlTA
0kjUTvom4WTydjM01fD0WlgXByZaHa0Amf8iZpvVCZx8IrLyRp+H+giQE7vhSOC3
YFGDqY4/vbeTNGIswX7wkSusY070+uwc04ELpBymy+6A19G5n6IPInlTPXi4s/xt
jfsU4/Kv96AYEDo6bizCub4kyZljRRDzOlNU5NivIAFvL+/KZ9iOf7MhQRIn1tjR
cImW+mSLCqvS+gOK1E0823bUx+zrae/xs3rVbFH0eubaQP0axiS9zDo3/B8sVHbq
s3LRR9dCciKu9e838Hx8/3nEJCcwGN3VRe9/Z8ywLImhSuwbDjvDu+woJbkys3xV
9ELJqSDFm/mwivHCmF7qy9w+ZECjVZM/BxcbdTlxYFRk70i0saDwZqE85E1ad3Hk
Y8O4PW1+ABGF5Vee0AtRk/+XZiafPkU7qU855FPuwcxpI9VDDXa84NDmMSRswB5b
sgX7t/NY/YurPQve2yvFvPbJHan9kECEPZaNJogWqI80gBspRKqI2CruPHmUd8oX
+Pprcv5yk6bh11LpjLKzoX5Ome0WT78cMVuMPfqH9wLZBwjKJ+HxWe+jNoZBY4+7
3tfhSeeSp02j2tl5mfcCo6+qrjv3YXn7h3zCrpozh7hN2GjX2nNg9Zy/sTSZOvLo
454SCha4TyOSVmqxf3y/GXWSmFQ4bFmNqoTjFTkazZalqDwp5yrPc0Y2myqEVrsO
ZyggeauQrgyOcmipye1353Q5VV/eJrX9VIbE8saQZFw5yw/pRd6kM2Dsvq8GVbc8
ujj6wDLW6WyvRtZv4ymR9OI6gSZKsXRclDJa7D/2hpaBeipKTv1WMLrUPbBgkdL6
fSp79qGyjR/2BKSdCEEaJBSnjsBnXxehIY2qVoVXl6nP4cNOrTwvbtHHVkMWORD9
a9HFd9hWorZ4ertl7IhsogAmF4u+YJX1eg3kjkH28X8NVLNekD/JPBNhqXcu1+7T
+x2668iFv99sDtAmzZBItochZchPfTaLKEl0FbMs/hHvzhXG5R5JzoaMZYZ+Eyz0
aSIUr3KsxbW1vwm9XitUIdH0aaNYLCrpDCzxUPrhAs3OEz7hlMJaxqr1LpAtxSIk
Zk/y8BOFEGDIoLXEO5P64FNYMS3jyxOiNEy15ybeZmt2vnKoONE+wFDRW2hFIXv5
g/CN8VO3oZ//hmwwuNq0NCef2ehuFz1rm6AEfXHgJK3TH09SeGvg4EB7MaWnDyna
IWh4RXOwOxvHlHD+GYtKhClVRprIMYlkwC3qjLQMvCMxMXMKj1a3phn/35RusjSW
NKIB5AyK3XAiNjfIg+5+JhsS2TE6D9mhJ9pjn1y8wd/XzFKmF5ssxA6P7XgjNsdZ
7ttW+wHIZlw+Z2sI/3QI5JUPPtBKyWuQ5JUzgkv4OyA8dMZToeutNfMJrLSlyqJS
ZJSXgxGQrIdAngMsRr/TDeUBJnBm9VcJ/ssxPaGT5XLBpIt39r3z2hCVKEhoC/ks
s6GDhT535LO2RV8QgphCAi4dRd0UBeU/NsWJI5/rtGNCNieC3go8JhlQmUKp9lI5
K1i0TCVdSZM+F3Sob0pgl0rhDEw5qcdvQCQZsMlRPCiK22A1njxEKHYBmZxpnkpY
SIzyJme7xjae58HDsHKmOrNzxkyg9xhh9OjbkN9w3/gk8W+UvTGSXjBiAQFBRccW
JFqJ/Pinlvij/HbmU3jefpycKoxpK3Rrk3wuwOfvLIq+qMvHf+UhwKx78Ler/VyB
/8Az2K3nsEe7u2wbZrnaWVLWCqfIb62qj5SRoeNBxTPGqzNF4Mx6cwqY+qGBDMaW
Rmq6IAUT3tZGPw/7FicBCQ9v35lnLEUHs93tEY20JeJcTt5g84U6lXx/8ned31ZQ
8z6g6XcYLamkXwFKX2RDLLsWVNpjVVVAQK4BB5L6ClTQUcCe5IRrn1c+6Vzbc5c7
1nSVxPmKyDh+ICQEd1edooZBEzHr7OxfKaYYFmcDq6bT/3KtExeatpp7nSuAD6o3
OBefaowm8DDRG/SSsmQ3rajuezXIdTuV7xmaqoYaZex4nFS07UXJl3x0RZPfwJtd
uGq6FQHjFgY4rOxop6R3WHfnZ3yGwRV88rGuaYGFlQ3aM32PrzA5kd87TlQXccfp
iPwhvxuoh15ItbRAYwVAtnfLpPYgO8jbpp9d/Vtrw9Xe6Vy8+JJ7JAoHmNfmdtuY
orCqBZ9hbqPvoGaMMLsutRx5pam1waHjmuU/BgNgDMr2bol9qU9sKVO01jekz3yk
xdDK2BDNPtTpCogd5AmeMdZxZg1v5/lHb3BlkGOMRDXV+yl3ARxEFu7KPhUOL2or
6BKw8370YCFyFE3gvTjDgIKgZU8eJc7KXMJc4gvEwzZRlxmqmpQKGK5m4+UxKjLs
sUJKoJ2XkKLzpPaTAfGJ3Q/URjKgYxgHKtW2L5FD8WbWGKskl0SrhoKQgptC4VaW
ScgWSvc6Mxu0Wl8zgyPKUFs9+N3AnXTShkEEZVrmKBWA2QIGEX0MapsSwoFJZyZ7
Kca0ANOQezbiS+u2KUByME3pBBy8ErsSO2CKyYJSNrMV9OExDsoxGy1z2zddQUql
LSLvsDcIpwprDFthXBrTJOQgkJtl/pQ3fQoCyeUuNoY4arcld5ayaLdmEPgm0Iz/
IMrlH6ADAFWOovNh5kIzjRqpyJl95PAxkghXd8SJcfgNAPhflSMTO7m+GX37fd53
9PebphPFY2pbG/uHJ07eOreWrqN2TluYlpdVQP0MiaXBaaUayp4DIiX32SGeGUrZ
cln+up02DEyvkyq7uYGAxKJT2rdfuCIk0SAyWLGU50/6kPvrGWl0N8CbBO5UhIOT
NCmtUx/t3rDaB1qyFAonOWHD/B72vGT0vDVUOzzLOJGngPaWGpdaR04tKkFkPgvt
IpjFZ9E1OdzeGGFxZTr5htDzJTujb7q4y30k5z10r1SdGEdjVwF04b1sJoOG8s8p
mAMkzjugBBb1Baf5vzOYuARLUPvwwSLJiUvD4OkYZzke5Obj6Y97EIMFRSUUiYr+
z67Hi39rRsxS5s+rlXZ3N8I4+Ieo9f8hk0LI2D0Df+LPsQrOZIlpiY4OftR01zoh
tG1Vcgyq9uvWKBresqmLNRC1ro8saL5LtTPPP1YvH4bMr3h2OkLcdrwzagKaEfn4
qMlUq7U1tHxa737gBo8YOPZvPJDb3+epnt0fECDRoy11k5xE/wwnP85FWGPNPfsV
pRxhEPI/hFzRHVkqw7vUCQa3ElvVdPswde8JQzgmM1XBkNTe/PJvxgNTWb/sFqNy
6XfNt59+TntQ23VEEiOpoIEa9D4St6BRI3g1k02GPpenWJ4z6Fmd8PIuGsOggysJ
Pffv99XG3M6bJOgqxrWqh3zYPRejY9ceIlqVE8tdWQbaoXQ1kLPr7PAl+lQ/q3kW
SyES+vlEK4/wLOdTzukQPC9/nIaUFgQNpwsee0U7pOJ81BI6TRwFZt5erKDbh90h
qRV4iX6dWDOhVR1dJ+O0oMgVyNdpkbr5RCELXFF1febuOR8wKiRfVpN73T+NnQQn
N2lcnwVr9O9Wzpm4wmZlwAMEhHhpMaWtQfuFVrcT/UJaG6ADpnArjQmZdIli8Pl6
szTfUJD8ms55wv1JMfrFmxTxhKgG9VD1ibghpSAX5r5dF3Dti5xyxWXztaqGCrVF
jn2iyclTxEHCeATVufEXRT88NlBwbQ0O+QIUBn5WzHPXWPjqv9sciPzAIgEVpFBR
Bc2TPa/7j2RQdVve5k6F5qt70M59WtDU9ssEU3Bet76ij/KtBBvE6+FbUHi3fW8g
8P6gKVzu2skq2tEHFkplIawiyB7+A6tWKncxRqaN3kEFtpon+JtfBzRZs1BU6jl7
HdBLgXTgtDO4ayh62wNJ0g9pT2LQ1JVpIbj3VZKRoYs3PLSK836pCK18GhxdQi4L
ELx88kMP74w4K4bDe3cEWWyJninWDTJvsvixN8tIr2rZ3WQnIXu62Wp2RGHjOpi0
Nr6F2IjJl8ozRp1NQXxHdCW08uXVFN3Fd9BQiIhut543D+aw9MxGQXClDBBtKc3D
srhp8SttWLxey9+cKC/Ad4+Z9x0GJpe7TyLCKmnC8WDLyKuptaEQLwHkUk3AtsOO
GD4/2suL6OuXqsZ+W3t0bwlXXKz/25c9Uov+poDGK1atw9BL7IIq1vanMvRjbibb
qOBYnmZBzohKBir/dWPU8ilDLLd4wUYQ8QvD4ZAHZGB5gT6LkH5WMPRJfERilWp3
5t/A/HJTW/7R/ZVb8w7zScoSorBLaxDJYcHkxxslHlvghLVRZXiBUhzXswBp/m/i
C1AUTkCCRlx/kuGTJr+1Hz8i2NyYBr7jHJ/JWXFy/GW6wBdWE6dThWPGf4qQQp/e
X7OSwHqvbATrJxwWR3+z5NQHJj0pvN9U7IhBfQ4EtApmjdTRzJXC3PsOXZ1ZRjSc
4ZJ2lBFMstlyI9WnXjzbyc1FrLk2gKq29wBDOdnyJqLPoCMJU0uRoGemp6LLylIY
5f2q4AU7310s7qTTWj/BrQ7Y8f8LMc/L1lbzcDMKMU/DR/jrkD/7vpfvLYc4OhsM
E9a7AEjg5Vv0aezAweoAYfnlSKAw12gscI10SGvwtF1FRTVhFwufM8e+Qq9WOS5b
saaqAhd7C86GWOwKDvamiYChgfM5yrOIme1fWNFdihMn5K0WCVnIYAfxj5ICOOza
Xp+H7NDQ0/jet4fE1Ze6FM+mOI+qXMVJvxx9X5KLMXZIk/X2tQkCzp0e8CS049z/
iksX3k09vzBNhbiyDXu2hVz+wEBbGF/H55y4CjEe6sxmsbRnZY/AZk7ecBT9+eD2
LuSKgxJJ2bBZsicNWBK6NK71ngLQ6sZMetauPIy6guLbaSRk2P/s0CgWzsaRhUDi
nr0ZO4hdo/iR67MmeObHL1ePkI9OXb2zaH89s/Mr0vQ2tIev07BRNG9e+foYAygE
YYOpAJzOKeVJCDS6RFST5I7URW2fm7ZSjOcuxlqJ7Ocsb+N9KfhtVymsW6yz3vIi
ue69R6XDVqKOzJzCuYmS2H34mI24tR2N46f3hnwh9dHxSa3duDunF4sinmKlSqHH
5IbIgtqzfDalGMGVXqvr+nVZXc8TRt0iDnAspbY29ZwbdWA8aW6qOmNPFoyn+E1r
FcHXRx4bz146q52JwbykWJJs0e24C3ge7G1Scha6J/VbZ6srvHLHEAJ92Gn2mZkm
JPbDid0BOXZGA7InsESeVW8wawC6Obbh2VkF1WZxAXRzplY3e/79+KieXzERubE3
A/L3ZRHjysfrJYs7Z7DSjfq8QDv9+dUsG41C+519xB3YdKxkyyhziBoIh4LNuXT9
JaMewxs0cC2j/eGml96TJIZ9agLwR/AiGFek2WUkJIJTIXBqxJS1qEcxDvONYR03
Uqv5M+vwG8oRJl3Kve6DbuAMVa3nibm2+2O2jmXpeerdULKPVAxIDnAPH+MohibA
QrBf2qt/2tiM+7qKCQXpkRKkWibuHvnMY24OoS+U3E9XbnVHxedHZNSrnu3pK21f
VbQdJ4nUA2uBWl89n6SQIFJEK5ogeUpBAmX2a++3cCZCFZuhWBgZP5BJ71veaHQw
qhSfoKcVfSqdylDFBtXEXGFSpWDPRDOgm2juLg7WRZSdsBA3912RYu4I8eggdxYi
5ag/mxrWJoVXR5DkgrXMgyQTTbNwFCm6Fvx6pRAljAOMTbob25bi86ra6l7m0lYH
EPonLPldHgog/Zkmy4i7W58ZdQNRT+jh4y46t0FJBngIZKdtRNk9aFiHudS3tJs1
TJg5AT6YoMbt62u1YjWqHhnaBNiP/iX84PdE6QKYyHTtlu33YDPfFSYF4GV2NWp2
WLaPKY5tSTDpdC59gRsLrISHwQbljDPSoeB8Rg25RCSowD9OGkXRhyY8rItBHtQ8
0sqQsuO194/BU5wh7xu+Yo1R6w6puIOtY0hZKty/vn/3LE5d+0CPw706ox6ZPUTj
UG4R/7ybr8Kte2tlBaZjQgcDwEBbypLM0zycVH2aUWrGBKBQ2kGlQdC9wLNDMBrP
BkVJlbexNWxRYGXMg+S+vIxGKJ8S1hOEBPUxGVu+i+jKkd4yWSAmGqDhxLbVZTG7
vp4gmaLuaHCjTTD5pus9Gm1XkfuCon2jBvIr3SuRsQa7fhz752sqf1i/d/kOg77X
kYxVeMwpy5cByHl6A64tuggSZiKBuysglBfkFhQesQMk94y4bLxC72L4sd71LuHn
GPNXjpg9vvtEB8dK5z3g7afmcRWbf/vvG0NNdLyYToxXlN/gfz3jcu5G/Sq/i6Zz
Oc7wVRQLUOaDWDfCvNMA9t2/YFM7moKCt/K7SsLSppA5EalLA6dspg6ADN3NJ1gx
tGJh/Hx1OEhqV24yQ5Jxws6HqsmdhVJ/gHr+s5oq1aaRyqtbMd3a/3hR/85mSFIx
/mHJHk383hFsS2sOjKfgdtfRNbenKPlnGJp1Pm5gxUpNUyyKRyInpn82q0kyIL0S
fQ5m0wTq2v/DOW7hqhz9RmAiqJfW0EHvXJ1MvEAIiqV3wS2p7OIntPi+lYKsS3AB
WZWv4LQbcZq+f68F2SqUqRmJtM0lFQ1YlLxfNB+9tltcZkBHiYInEJ+XcqHnj5EV
dJXl8dza8iOUwlws8ONp8rT8/W0yfdohniwIYXOUTLPD99/FcE8snwhIqG4bR+qo
tOZ0SyejywKhF1dFV3Ge/YEXKVHrhlGudGDqQxeSFb04ZOa50SKFWagL8a2Is0xJ
KpNb0YwAEMevLlSDVaMDMSgT73paaxCWgFvQwbLSE5annnR3jEctkC06alK1LP7X
ZMJC8L+OVDhDWyiJ3ZcDSWAR9peqQNRm/IqxA/S3iCexsTREgeZH2b2mrwbMpAXX
JqQJAoUxQxMLybqQJHMliGRvwc5vPu+IvsR3nI7ZxwshcislHNIKajhOpd3icJv8
R1Bc9AroIF2WMxK3fvOB9Fp1nRFAZK7G1sixD50NYcnZ9f9Pz3M0hFGBIr/zrQVk
3fcZbI8bxZNcs15CLrbwCTBajgIs8qM/UNto7kvOSW2wSRO4B7E5BMFDKNkbQJhT
AQE9IKKlmjD/TaX2Qn+LDnmdUw89c7FQhukYtC7wV1v0f7gpw6n1Z0nH6qreuQ2T
JWNz8EjZPAiESDm1FaY6dX4YK6jrbrPj/jyk8Wr96em/W0PKIfIA9witaaItl62G
AI0RgmCVMvpZ0ne5DtgD4/hcW3RwskaUOhr6ZhrNypbqBprgAQ1BBbdN0TXkUJEu
0zWkVb5VPOTWgTY4r2hkUUkszNCnB0C6ukcVZwK+k5Alps3SVe311W4gIJ26C0N2
NTypAFbNYM+SlgzHB91491YKuTDficXPIjK+WLPDm4zYK1X5JP3ZkMz8P/wxcX5y
B8F9zBf2x4OwWHOnm2Da3Mh75quzrFYC7pGZja5NQ1TYj6cRDEq3iv74aYtOkM3w
6d5SLPHC1HeQqqmvdxz3+eVEanSiu0blL1G1xdSJwB0SNGQUs6M2XH+F0ro4D4Ne
zsbD4+Gw4uXeMwBgQRSxpLorqB9GJF8x96T21H+7laqVsGasFb49VUE7a1lud09p
hXQubpmU3X+xcjpkiWSaXBTFYoL5XA+8gxvE51amD6rQ76+dpGHotTzV8xalINT1
jIrk7BNq7Ngf3dMg07oG58X0CvyjgZM1CjSDXUwJJhaXYoQBTYdbFaYt+5+gCl4k
ADGH9q/b3J07c+ElIYvziTpqkJzMNVwJ/tIsovy7sn1+5YoaANELZMSf3rAGPlCO
J8pZISZudHolTvAiymwkJ3gETrbOjmof/dMwRyHpMN9zcDbozJimEMnfydaTF9fW
RtOdEOPc9bn7O1YUULxzX3YHUbi3SOkgT/UDryn+I1i5ONtl7954xJcsaf4ENEOU
1/8QD2PhnQnLK9YBmJeQnHjsb/OY2cxgasLtGRscVWmvFy8Lsx2ADkV0F0UaQCVt
u4fu9U7dlcpvGkQUdpsxD2r/fOcdbKOwsuOqUV+PdEeltiA0v2G46/PYbr8g0r4P
dEw78neUC37O+/+B6MzGKE2X3SCOOgiCzNt7K6rNQJvWMfH2ydUGdeeGcsvvJ5cI
MFxmM/KrpVNAaJTqnew5NqjhBuQT70VN9ynyZsruiiEYMbNiQGxr+r1mSFCA9A3R
5FhSiIprTHeCkgX5gNIXim+MUzuTBurpw1xwADy2nPpFYzriJ64dbGTdcH0CwBq6
grBMxOicupc5Sa9V5jYlNo4q+2jRtHMpx7G0xOy72VujZLCh8+PJg+FghQz8Dqy0
Kka3AVfBGMtUMmSi2ySlQfCck9rYs7nUiFtNyxAAh7Wy3chU/qXeD+BhzhjiYHva
hZ7ZccseEj1VuJnqayWBGiGkWa0DiV+xiPrM7gEFRUfuicPxrdIT+JQhhCgaMr4h
NNGSicUKhyefQpr3BRzPZuxw5KQSdgmn3MOH6mMV8hhsoCqc+24GkEJmzF3uNs/x
MURw3a2thZNXpQlLEhB3KsdMmeGzUog9oqctUhkjQZ2UHwc3LfSex/9+NsMY9t05
ABK2pHSj0Btf5ZcYdd6JESz9dReNpOLrRPJsYc0wokATGf8+3Jo+0Thec+R6u9YC
DVsiz3sMa+jtXdQO0w2vttz1bkefTgMdcZzM8uAIRpBzflHYJZYDRbFzxCvwjo9k
3Sv9+MA7JVfn5fw7Aiarlz+EpKS4pnIinCIAWYsS1CFebc9qZXuSmefTXI6uHlM9
xi14XVfEA5ci6dnD1JCkjw37bL1diBz/GB7BmpnqjH32lQ5+432f8dkJfGYu9qHX
+llPeS7L6icIKTzwRhEztxXdIgGgDVPksvWbTKCQhbj11RUMiV+v2VVwD0bDri5U
fD6/qkxouGUKKt/LQFVDhoz2SC2ilL730u16r8ctYQs6Yksd8ZHmqZ1XxtFo3pnN
pastIa1B2Un9u3F2aXy5vJ30hZmmowmXECFQ8oZDJUUx3OAf0pmwlsxxQ/dqNQwF
B8uqK4HLX+7VhM+7xSafDTeU8dO0kqZU4PrhyGvafliLke0axAWYOsOSywotEVN0
pJWYd1KmMsosiyW4nsdChmf+lLau6pEJgdBDHCPbBKZD8rGXhPZGJ0YBmiBbcRBE
uViOXMBIX187Mws+SKrRkl2ky2LvykTjNGVMXcw8cwhnqDtXKjF6O4V0ZxVUl+FZ
3aMsndA2wM17ZuKUZstWD6FoGocqiPAu7CMBoahC4yiyFH9cWDyb8KqACGL8XAel
0Y3UQN+N7q8VBatzj228C8p3/EJaPm2Gd+g6uX8GMXo/4Og5qoMJG3x9FRS4oWY7
GCKVpna2PDFS0M3hwmYjShkGG/DK/vjccJlyZyBqDDJQcvTQAAfih8GkNXDGm80G
BcxaDeITK/yi6uY4a47FXtrbA+2rmVuW3Mk88VDEUwpwRxH15iq+ah5zN36G25+d
at5UZIYpOi3LmeaOY7DgVRqglVjGoLduU/xi24YcV8mRk+JF0wWrk8UDebhG6hG8
ceyTj1F6Q6JGazi3LJMfxYOH3ZpJXN2/tZtoX0kYKjgyLvFvBs2TBAFz1/qqjhwX
FJZ0M5tp/jsV2H1iQeG33DLJWh3Cq8x+Q5nDFC3M4WUeFip+7uNgcsHJ0aVugVPt
JUH71kmAPIYMY11uwE4DW3qeAmvvbSI30+CPhYo4oj/hssAtnwC/ggiRww6Dpmiu
DGRw+akG8ZkNoD0ytso11mDDFzn/K2R16UIao7YoWVUeWaCHxzOAHCHQao3uNO8J
PXmH1uVYIqhkI/i/8yPzkb/t6olBIRUcnvMorSTy9+ZqCsbkuJL7RwfjzwfQI/xc
7hDPsxNQnFnvi+DPdIvYghWq9BjIicS3B9G+VVnPpesna80uh11nZWs4DkuaBZJQ
5dywiOwUjXYs+eMtScD63Y/D1aewjA9IvpAFWd3TMXUZH/rfG5/sduwMLDIcEM60
T4f3zyEchYSno6Dq/73vGTj8IM4eqsZLZK5EXXTM3Ys1HqJGGHHm+DgYI4oTHMKQ
Psj9MJGrc8bUzUJxjiZgP6J7ZmBDpXtX1PQQwOrz1Q5eGiskD4UQVyfYB4j4RkKs
w9JMzNXtt49sl+gfdBMTMyVmR4u0HoWV05abHKLiIpPgkRqCmZbnH5NMEu5Uur2d
3pxAi4rK0D9o89XcMgaC6RAnMEEEY4Q8pgjdheGemXd0BMZ+stdvEL2VqAGssr65
Sf2AznrIvALHke/dDdRtlf7k1wBiV328Bdqc1OGbviIoi7x5xAxOKqqKT8xkX+YQ
In4dRTqxjrStGmvHg3gIz0rCUmdzO7AvqExvjBrUEYDXfZhbwxAqcp5OKmgfJIS0
gX/WeczYB838Hd6NX+c+5FOQUr+lZdpver7496BFaCO1v6f3ptP1Wo6qUsSwp726
s5Aw1pZU7lN2OwMAI37kseAR1jPzqscsCN2TX5bllUVQscThpTCKzLES+ngWa+FB
9vdmG45cEqZfaZ5mIlHqj7CXNIZ8yXIqQDP8gauHxON4g8TiAgKb/5Xklsyl4Wjv
Z3Lhx1Unx/QfOn7Inln/qw+oXkYumrviEWZWEI45tHQU3uDhOiweb9JfWJMYjslE
+0r9N4tdDmZPrdHH61mF5U47eoZpD7TJA5ygBERbs4bAEgvV3DCt6MfT6oMRWqh7
xFd9pXetayA9IS4TyKJKjOyPeaMluPEB2T5SKvhSujI6CZSgRgiAtUf4ZndvCbBo
X0uGXiQiByr0WMwKRzF3n87Z22UtMICVdV/ivvUSPYj2b7EgaEvmyyaLtymL8gGv
2mmMPJVWzZ+1iRlAQ+FfhGSUo8bm9cG6ob275b8nbo9PRlfwTkG6XZt14kjEmeLg
0gSu/h/Tp9NpOQ8df00SINIUx8URHyBN8VVjwsd6RUZ2dJ6Eb0g4PeXt0wrnovKR
iT+J5PM1BEvoKusY0n5P1IjemhnlcrAAZ0pCvCr+ga12sx0LFvh0z0vR+oWuE67A
FnXSqUNnrTcafOleJUSFcF5/THs5b/IwRHQ5c1fuhwicgS0LqWccz0X54+RyTp57
ocgq2sOvFiYXkGr3pv499t8EpaETgIhUX7Er+/xk+vU+3hMGxysWk9Gffr9LgeNy
yQKp5kbHfAJr+jYw+t4ywUA31whc+wsdOxJuo276eCQ=
`protect END_PROTECTED
