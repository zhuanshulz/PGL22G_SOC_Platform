`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nKpeFFGrsD+udlo41pZCzW2eq+yy1l2g6+iOO0RqEQvvpxxrLd2u1a4UsefVk/JT
vfMMBaRExlMrdMMOqiT20+rUaHczOSje5B2E0WEncWsy5z6b5EgTipieKqmtoOxl
pIQC6Ehc1C9xpoRnkKfiPF4TO/hyq4C5LfwaZpE9SIRDYLaYeydOVw73JL59GFrk
/1G6X/ChdgtnPozJZGXMR0EjrBHnTDPo24n1X12WvaHEfWxpallddRX5Oa3s8dXJ
ZAlVZ+5tyh8Q2gjM4SdrZWAbvEgw8a4tknPeE0buDlU=
`protect END_PROTECTED
