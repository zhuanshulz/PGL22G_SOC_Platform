`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2/9Whjfn5wZ7ydF5tA6DMQqjzQgPgbD6s81iODypfBGD8hNasQuX/yDDMbCAZxU/
ICSkQK2tVUNXgYho+eZvKqnHYNeQ2P5/qFayi99EnrnafTDfxCvKnRcsjDZdm5uJ
mRKvT1LG5dPTtj4uabShesObFIl5008i7pnJ7r7/0dphGEhFW5Xw4E7PYU9eHhdP
FHVs9qTtJ+rYHsPOHLyHHD/bTqn5GSpfzonHXyvLjcggjwqTMeE5Q5vjbm3EGL1d
UV4NF5c4rHCwAk/j5w/QU5OzBLR9BOR1nNWxgbg6OhRuBV6Va8uCZuoL4VOsb0zK
BopObFHjOrY9ayRczKiOBI8N8YO9z4xPfVFkhRS/aco3hFxA92EzsGHF1wppJe10
r/6g72LHZ0NEcUyeYy3aWJUQ1jGlvNxmR4RICkZvb25afonWce24ehPB2qXDfVOU
RdN/rV3aCzhSOUnLyM9b0GJO1fdQYeDsU2x0CFwptSDJIOwg4KODA88Q/2e5tQkq
EL78dAaBhosFaCpIxezNFP3Q+F/R182YH/dH6JVVt85LLZ3eUst7V/o2JYv3z/PY
WlFw09K3ugLxF7TOOSq2WBPb8Oge9uErVvIxoKb0xav7EDlVNxLjVD0DyDBR23uw
SuvlRzJ27B04Bbh5pfqdfNYRtcCtHDKqTnUxvTGoGIj7C3cIrIv5x9YY3IMs+JMY
AQpHHPehgqGdCqXTCIyuTXULmJG6i9TY0jAMMuo14NJVitrSjz1KH8LkBDxN2CBg
YqSb8k0yB+JPZDXDGs5xEvPGbsDBT3+zpZolnQcq5txWfOmR91APZArd9o5ovNxX
VvhRQMOrGFYhF5Hbvfr03FiNJTPvpTCMd02cG7TJgNs2O2bWhYbJej9oh6r1BvyS
wOYWmPAUpCedgTHEDLawn7mxdLvnFz/C5jHiZofe8kW7qI82XrwOP7SJtqEa05D3
0kXd7X662H6WzTpvON8AMh34k5Mr596hsY9uVpqrfBKOlUqJBuKSnCrism8womB6
n9PVbCnn6l9vt1DmC493joTeIozW5Y2c4ojwkhU49y5CORty5B7DlpzfT1GUs8F5
U00JJLy4S58Ovun/H8CZqtob8gO0N7QGOXDbS8mhNBw167jT5605L4kiOcdq/ry8
oYTyXuMr56Jn63uc3YnqyuEZWGnUX4uBPSKSa06CxYA52GZHAy7GKUD9MPDJ7ref
fJnyY3sN3ejKEaz2Ayk0qWLe1wuZA3QmKa7ps7hhCZA2w3bGAXscdN0zaYmpT0q1
HGOieGnJnygp8DFKWNVsbw==
`protect END_PROTECTED
