`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kmEXNHlAnxN7PhxzBEz6G6xwgb0p5dqXNbSwjettpm7hKGYClmjp7GEk6QGz0nb0
aCeEUi0o1+mQIyYFuH5MnRSzfBSEtDNQ/nZ1yqLdFMw1CkE5J1rPMhfITvoW67l7
gsxKtv8gTDstJNQOnyvbtw4913KPrSp1Ce5kKnTMFPfSBU6HHRtDu526c1jiulCw
a9BvdJKXo4qf7Fu0fCkFGTEE1qAvyadE+XrLSkgRLyf3nW35YuQ95j4sqPQ31hYn
jCAHVqTdWTdkbjbBXYlMoiPZY/3sloXL2O7YyoZkFwyDTtsvlCjKdhRAoXb3ia82
uRCrnnA8Q/Sq3T/y1966STJWcOZZb+tCaC3mGW5BPM8QFPkNFjfmo8bsBFmuccLc
GXVeQqusxnZLCuyZJG9sNpJra8/pqkNyxmNrfTJPntg=
`protect END_PROTECTED
