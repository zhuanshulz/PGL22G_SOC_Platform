`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZZ5+3pAOCmj4bbwqWeOdbqyzyPiX4Om4Uq1bu9UgugQJNGl6gpndQGid3BwXvkcv
pEHflH5ENblfAn+861tuMbVCVjjytBRZFypNA7uIWA8G38R/ft+rKNbzZhiZfnsp
NwJ5Q3x8NwZRpwz0WPGqwdRNkGiBaPcGx8b4I2GSb7FgEG2egi14pFAuk9sSZySN
0Uv43E7mP0bsq2ijTsRTKhuSv+84yB2B3U9ERp5RdXVi5XuqY0uMhyoJ8+PfhU2x
EuonP/SjerxXFrlqepwJuV8haZ8AoTTrbV0BWDTSTiqYerfFtwtaVIIEFdVd/Zk0
49STDM6oaNBQpXKZwZ1ly9euHAQ9h5J9TWx2jkSnUw0C508w7GVD8ZF/IuDqMuIb
fJAW0Fwt70qqc/xb/hIYS3Mh9Gg89aVwmFlGpOqBp22dXcM/LnmfRlaHQz2O8LmZ
vtW9Jke7Zg2aI9nn4tmvLIoNqibu9eZRaJFF0o/Lt+R+ugQedEyIyCH3iXPF7MPA
4Mo4bossWsLRMjXH6X515FIcScPf+w7NPQnTzbPMfxrR4KDE6jfmPSLw9xUgLZbg
oSeig+ULanJCMkwFLpzOzZeSsArbG/5dLJ5baDJUpVa8euf4PHduuagG2XVq3sEK
mS4waSmlvfR2pBf8cf04e2S4oFFBTcYp57mVWACr03+a0K6OimBpbM/MMKEqvUee
Bc+afd789V5JQoeFHM+F7zvhr8r6KyG4O29ptv9Pc/09brnzhMCsUsZS3K5SXG6G
+p8iayCAC6gIpmTMZnWCUIaNYcRme8sQqyxvQbMnrBdDQF99kVdm6J+QGJ0p11cs
wxE4228zU7HefXJvYBennlQrD/GPVK9Fw8YHSF7Pbk/DpzSixa/oZi/IznW3beII
YTXrfn0QybeNDz1aMWjz1VTMrFaTTMzCRuC2m2H4nrs2teZVto0XaCYlyA6CE4Ds
+pcUsyCmc/0CDHP/rPZg+k1YhVd1CKisniZERo/oZ/6aLaKdApwudQ9tAU4tzaZp
sW4s1oF+C8RsOHTMPgXSmXBDV7WoXbFZPTax0HZEes6cWjtHebCntLSpBa20rxCv
uP0qEVhh0TPola60TDUVBR8j5da4IVXURFq2SkOEBj0rLKFGz+XaYnOYSgQh0/xN
AatmBFQqGj7+WHlYlxemBuodjIAYEpdDuK5rmFDOO4sbmbBctxfCilHDGvghtgW6
tVIsentNl5Bq+dxCssARwEvat6uCDhC9F4mJ9LeEvGWMoy53AzDT0glOZrAVfNyD
3Co82aVNKUE5GDzG/c3UwY/hoQQHmgT+6hFSXqsqbi+B2tTvSuXdOlnZjIGdKAW2
7EkCfaR3s/tF+a4n+HiTg0Tjg7Njh+nAzLzpwX6coKfXJtUxUyV605BO77JGJw1D
fOwUU4EUdkEdRX+va6X2d+n1iLXfBygSPdcG+OnehrAoMZLWJ04rbl4ryyAY7MC5
DgHVFAQqOJdrOu7prrndU/PxGPR9d9df9iBbM7NXvsbGwr/oFvInVbW4MT9Y3x6t
Y10pWtPbav7XqRC/YyIVCIx8ofQFzabte2u2MFMr9kiNsQvFBsl7m7SqazY6IAqx
4aj6Q7eR/z95xH7KFicC5JTPi7lj0zIxbspHyAbcwanuzFWNYdMy3Q+5yNgPIdbv
I3UknnhYhsagCPzZc0yor3Aez3nRaHLKBtgvDhVozfbTC4k0hlJ3SCibQkAw8mTY
v8apA7LIKRNW8ALSHjqw8QVbCvU4Xq0r8YvqYkAS2C7NimeWWr7kzrwLe+6euhgR
yC9BiUofZlzqjQ39wmOPJmv8qkko9pmbj/UVgPpK6najCrNRWSOzgYtVO4jBagBY
4fZpxYP1KXpDZunjA7QVt+IFP2C3xOk6kr7b4OOQX8a/qrCzlqrGYL3hrKEryCWJ
5LwNnSIY83AgmJ9OmbOcIoyN4ligrR6YEFiJHA7Kr9ox2ser+oP8p+CJDyFIQOps
ewkHFKdUCmd9j68YFNfbz6vmriV4AW2CTMkzHNC4C2TqSQl7qHEyngOZsMfH23Fp
NrMPXpIjoU8vZwlpdqkrGxcz/xNE7a95jrZJShGthdVldLPF8o/mqUESogT900Ji
ySiPLpQ5fRETcMvCWfOjNQIE8lrUUZIzTqPrFmztxiNWtPfbY3PYDL+6RID2nGO5
UY4GvMg+i6MJObJq4oF8nNu0MmDLZ8Sgfd0b2RaetceUlYiXMJavdmwg19ak3nHZ
7DwDXShBLVurFzPjSrGIKTAsR6JEFc5ByrUjnpf09g/MLYyc0qyMj9e6zmgCdhE3
gQwjHbwxWZCTwNQG+WiWNKhjtq0klLTrTrIg9QPMfFborkNd80h97rhstsb2sx02
BkdSGstFlemZMy38winKWYCmssJ7J2XeooZa1yMNrgQI26mrn0Zv/K1gS9NNt1+U
7PE1F7nPpZ9qDRaNQJzs+nD1PYTImFabdx+n7wRCrGgWMCX3AD+sAvhECn+ruOBt
FbHcWq6dZAXPrQGkZ0wPeGg2X4MQMpZ2sSz0vhpk6snP9YFiuGxkMyAbjkGtl9aW
G06oMlno0EIr8ONcVGL5jAVpNOeTfPAOdxSMYkpfo+RwcJNx/jtyC5Y2iDE4Cmc3
BJVvjwmFks8qOCnlcD86RT6sYWVGOvYwPS8dvqx0UYBQDiAvhQTpA3yWZBD9pjlh
LmBLr8a0kgLBAZO7oyFyZG7z+vHkP/EPeoK9RVDN39VNW8EsDONJQyYJj/ebPi0u
lV9ZMXTji3BsRh2asSs++ZaaOPFFk41g7WAcNcBYkNz51Ep4M9VizjfcGPYTf8z6
jNlDXvjgGPcN2Zskd5Gy5WIvCuY84YE1MKczA8icKc9XGxWDpLdfoqIjK/cwDNp5
3v9XDhvwLswMwZjTP2W09reLCkyGmmCHabRJtz6KLmH+JsALdmoQt+EhMi3fX5LN
+dud1xjXrSlgMG1Db+O/r67MY8q0oO/dbsO9U88UZTXs/heK8xaljPqxi+KaOOuB
m+mYCFGjPhVDLUcHUgiUvknnrQlRHSQKvlcAbkRuIw1ebzoubMA0FmmEddwOPmlY
n3l+2baNOLFAbNqasma4ULEq0620KKa2xN1hHrcqdqMorkzwzzjqEjbOokCRI/yt
7lBMFN9v2TbJgycW/C87B7NiB6sxsx5ODe0UOxVBkYW2fnTK4qlOT4v3ZUIOV2Ok
CmHV0A0Au0gKC4d5mMQ7e6QY+ZteJR7DsBffpBrwIhy5WrDaXMQjCgcDeuriWSwv
+fbOYWPhMcEWDOE4WuYNM3hijObg/ETnwdhUvTPh/X9GWa353YIJlY3RziG4mQWq
EL+ZFJ0aCxpGM5e2jvborvy84UsR6SKdbS4ocLouESp7TjVC6rXNEPy7kS/gmNwe
kxKYueeZtY7OCoh/5nq6IwrjshhplUcG7r0XggDCwd/KuR812UDFYrKcO8dd69yz
wt1OZ1yVCsAhOUU9/NOrYY4W2SbJPV2o4rpA6ef8Ob3+yZXPcQRFDMCHHMWpTuvX
DLEWOW/TCF4zwAgrjlbrPLM+Hys4GYJ0mLhZXoGspVw8u8vd5dh6bYdAVR6A+F6T
mbQGkhVXXXfC0VtzwxesFqHpfbSrgel2qPnRWZyVSSvmIc7+z8Djb8TX3bkp1dj/
xRsWpx4y2ZOAAuUC7CsQiAET+L4BwcUlf7ZcLGSLpBMjR4rTv7wFV1MVQLp1hkA9
r63rRD0GVpQiEyx8p5vcuIrP3LP+YkgEnTv7G8OCFumvcgdKOBcJutfEjUL6/zeo
Ln50nG5w1q5lK5JbhzS0Hp/6NOY55XkKxSyh+oF5Nmnb8NKygRerAgrTpQK2XzEi
E2CrIJFVk7PkDMzQC2vZnUzf/mBB+UG2H4bVaGhdFA6COCTBTeWxnBPbKu194Eto
1M+7dAJcEAJI3m2C+yJj+MQBX17b0trLtqTu+atlVjbaje0h2xTD7rQr/GCCPEFf
hR1QX4DOeDhovXV/riwrL6a/fS9QYU1YpA4XWKIGTodGtz2/DdHNok9AXhvJCHYb
QMjfNwF0YKz4YlDLtztFHPboXCOVF62r3XJs3Qc6icLyb1kcO1i9IH5uDF0ggscW
l8LeYpNOczfj6E5sDldN4WvX98jvNuPy6RmcKDUhvVmSLi3UR1byyoaaal03zao+
hkPMOIzkYxAwyUuNJxi3cixHxJMKlzEhhQgS8yveGJNkNTZm6a7DEGGwS7INIdZo
dsKt7FLGwpkVznf3OhVayAXIX4NSqkp2lcVuiHUh4OAkJWSB5qWMbF/PMJ5YMhXf
PMcfsADoMAVrSIc6rrtGgj9SObhWbZchAlbnryiccZSYbaZW2J4N3EdRo2CmTfEw
Uet+8cSRhYIG7P9FQcWGxCjsh6kTEcGyD4E/MglbiwUn9DHz+GtGULLmSl0q/EKm
FxjYyjk4gKZoWo3M2ch2sMJWI8MTrmheB7BjNu3oBOZXVhNm6NzMdXk/BJPaMMBZ
5VFHzuGHrs6KT6BieMOTghC8ysf5xU3RxvcaNt/F1FOHrKdyFqMb/EwIG0GoAAgh
04w5Z292186lF2TMrEofV0WgFcyG3w8ByfyZWCYb8VKrRtREpe1czCpvqclGWcK+
IFg1h4qXnjCLlCasVKgwWWXK0lj3ZUuKBizJSPQeq8D2LXIqZgN9kg6vIpOrHg0b
2f08qVtVy4TtJail8Ow8RV0KoHr6qEsmGRzPaJ61I48gFI11lKJ16ERahKCpcl2e
TJaURDaUydnO4KaK9Fa3ssOZkYNJLepQnx6jj+vHJOIgV+HrRzFDx1wBIbTNLhW6
9IqxaZxeXyAwLQreFL7Hs1naYruVjMfUzvE4fkvCOpqMc74FX5Wz4skDAoTHOBbE
TogJVJoVcrjUcmsC8QMGNoRhGeuWH6emO8sOQah0uFoipCUUhY9pgTj+GS9TXOxD
a1427Jl3adoakOQLuawuXYFmhe4S167JnE2QzBLtbX9huHEqoJEPyHkdLm0CD5I/
GMn+s2t74aRnKCj+gg4AK6kl8IGyo4rBLXDpRMsJdPgNAtdJQzlXCTQcoY3QvnIB
nHcPl9Rz5dx0xTuqgRrvCukhkpdmexZ1uQFIvjPCJ18yw88J7ea1JeCx9i3rXBle
DM2uqh53ce15g8lnWZ01FTP9PpSCPpEe9GLv1wKHgZg9BuhOy8xt4j+ZE9E6xsDC
u0fI4U68K4R5DGZ7jV6D5urRJdR1Dj1AVuJxHSjCmPoCDA3BL38053zV9D5BQcKZ
sda7uSjEg3ZMTH30oKJz9TzP87+GhodnFX7Ahqp5HV4qLwoYeE1IG/5nO3bZiJk9
nyGbrvvIRd1IA7kzHxBBIcAsEsdykqwxcujDCIUu1HGbPQcw/rxp2XASSrQWr+M6
TyA3b/BqD7lGBK4ubvA+yqUFf8/iTLbOrN2srKTHwUm2MGRE1ByOztbmZv3B2nFg
mhRkYBLKNIGCkgKz9KWiNcLKi/Kl0jNVC15NafI0zTO2aRq3SIjiLs4IEBOAc8yS
nkAIolRpZQk4Wp0qF1f7UVTj33Ny6cJbVymYSF87fL2+NI73Unm3C91SfbN0dDAs
TxGTmU+PfGPpI81xU3/rAkFdodyXGElMA9w2ALOoyvxMpMtYDAAtME5Xv8z/J7JG
M1EaUNfbujjFEMqcQWml7/PehBmPZdlHT7OdmK+2fXrt5dRUc4+Ni41venxJmJV/
NRk4B2bMJmLPeigXuBnsqwfEmgPeodxpkij9aGKsiDOHhhFdBXtXtk+yGzu0hytx
Wd89BfoCLtKo2uS9uk5NJdPFvX08L1TUDkme4m+kpNcV/9Gt9hLIqIehoMI+1p/X
4lTN26HstpZ5zrlVbw7XsAM7RxwR9Kd9GLTtWuMVFYifmuyCaUf66aqkYJ+K3Dgk
73aqoZBuIJC0NIoSTfXBjZOD1tbMYhD0fowTXFAYw3Mi0yJd/Xyw1eFxoRrjYwpX
g96wtB7O3eZ7gL5GLI0Mp4R4pJLR1Vd+RE1Zg4lXF0G38Ps9S/NHI7OOX68+jN43
gv49LmGtp9NPJncRj//KIJJ4IdJ4G8PWZFfF/6alnTTlqwE4BPKbJyiysK7UA/SU
3Xt1JNqKCoPv1+1qBQ25/HMPXSivlDc7WP9N2/HE3JVKbng5Z+8S7PBDMepB2kJQ
0l6tDtTvujQAXaLkrFku1uzTEwGZcb+JQbwVq+QK8dtNWA/vuxAnqEFGnnR6SGDJ
7du3jo5I4E6WI07K50LfXBFO5m6dYUrztcRgYF1PSR12FqFooYtCSfh2r/YYu03d
8TSUJXrD74zjow6Dzp4t4UQE4Nq9eQWTqujuRfw4I94E8QrZsEyLDwkAwzvq0kYh
sB9TIwqKb24Ciow6Q6ZeIf6G7ZaTD0ilDf45+9wiTewAQN/dw4SeeQwkadiSM9IL
fOq/TmUI1GnXscHn+dAWK00tJm+Yfb5oFiLD23DstnRH+0R0jV6JBSjpgLpEMgSd
1KX9Q76N0RSL48Yef+GeSBWSp8b51E6RaPrzusF8UNiIA4jvAY8njNdK66pu+DFh
//7Y371XdpIrc72kHSAmTvYd/RR5aRcZ2q5hWsUR3Foe0ehyhGijQhDzEFMpwCdj
qnUpgB2e42LCh73hi1AMFZ8klRYBBDBz8iWllhwej6tr0edYMd4xj/EEE7LQIu1w
DyhdYGufbAOW2gBomnRP6srHWx8RQLhfDVogAhqz9dNnCMD9xExg++BseWiQnGju
GySGXb6Ip8CjJWrQF/1Zd4zErY1kVZkK8cETpN/PeWhv9y/SNyyeg7LyXIRHA2Rl
0hb7NweUfk0uLwQVQcUx41w2RiDRvySMaL+11od+fjNCGzqG2C3BkB7U7PpQ0LLX
WTsrv9LUvpViGA8QgTlMFKpXWOmmvJyo1QDhqGvDN1IYC1OmbTsIT4vHTnvreKGA
3otRSRuTokhDyNpH+nOD6S9vQ/7weTH6NXiYTNjbRWedCCPQZL7CVmvItDPRuaue
zKPWaQb6S70Xe0i5rfxxdKsxjC7BjPVYaxP2O9cuXhK+sbqgkmfdvGqMvFzolx6m
Xim2mCFUz5M+4uHge47JZVVmX7UhRu/QsblVPneeYAVto5BLxRv37Xyss6rCd6mx
qjami+OUtVS3+iTEk20wkgiX12ypuuaww6qN79HbHkprQEgczb0h5Rs+QCzXxcqB
0iDsj5ARGZMvQZYYCoX0eJFYAIfJ6yk/3DjYZjVRTMq/IGtKz6cvAJqq+1r8wM5L
moxkynW5slghDQnSH+ITWC79SVLgOfuQ3frq3HoIFhZXNL+cqDxypRUUPJ7rKWEK
NwrULEqEOGsrXiFLf8dVcqcFnANng9STD7pm1KHWrrYrL3LnkgIOX18KFFJ7zr9V
Qwt1xxilzDIo6ZmKKhsKtYGAZEJKjAduWkAZoxx08M9H2zBrhO2WDmzHvLy9guTy
JXGpSi9ByErBwn1vsOg5EgTSJOPtBseZ/Ec02bmM+yk28TZKF8/0lUHom5B2+1qb
bmqNKQMFPz7t4xWlsuokJs7XO/5JVo3mAABhdvmFszkDvFw/6Pwl8nYjb6+fqFe/
ujDJfuuTUXQhwzomBfvuGeVIzvFPxMPbDk43Uj4c4grlJiw5pCjE9YBy8mR+oe+i
DCVyR1AKjlIGpYyqaDEEgfuI+8aXU9cJbWv+WwkZfwIZPjCm9Do9KXSDCrQ67YV9
zPvOboqrAdVQGwNDzYm/Rw+rWS3N4pZf/nTaKU/tX/c8uFK51HslwDEj/7lfVhlw
fLrKPCPWT8VZKmUiBnNDILKw3Y+oRT1UiMAFaSSUqybq/wDNBG9rBA6saVp4LwVD
LAswLvAO/1tRqsW9h02UlGYUOJmwd+2wCWlFhRXr3kBbKdpRQOaZffMT3JKMEsS9
Gw+o7b11RZcdK97zpzEttj1nK4NRPKHPkxbleB3mdhFUi2Wfwwg6gkteVmkyn2rs
ZBfG6GzPCr7iwrs4uQ/P6bj/hcWgl9PcHjgqsF2datt9EnJLijg3o0OBLehB3iAi
peQkchigrKn5mHyxoyslln/pRAyoqReG0xri/HI6O9nBQm375xv6bHFzrY8hb67d
4qSfKFT5uPvIKH5kR1Gj991ouOm42EykZvztmTNJU+O+fajKe3fsGVTSbKCrPtjg
JR2WqO6bUqk1BSVt2NGO81Og2NiyfssEC7bDjn5eJXxPtXCZH6JRS/1E10dVjp0X
pq77EUAhRYpu3SFekEBZBycKSO+wK2TuZhBHxPJZqXqo1Qitk3rkei0VlXzLR5Z4
RB8Tj4FIomuP0CbPuTqHdPkJuUDb3vAEdFmMMVCC0gV0nDQ6CJx06GSgmdrPJagV
brwiUZJaiek/+Slw9pwb5PssW4j0Gb9S9e/SJ9qOcmsQvcwGruRunNp+QhBczYbC
sq5FIYGTI3z6TrFz50hLUAXEpvew86LkhrnvtnQt44qFqI1pYT1cKfubyUZkW5NI
AJgEzpPsrTHUqs+9bNE12wuaaPRt/ksqDe6n5RAoyi7aQkMr1i9D9nZhovWwVicE
JpA9fB8sz0aeLQ9NOlhg1o9fT6QhGSLpg78a9wRisVFfMU2cO9K1y/wqxidFy6m1
iHytu4lf7hETLpIQifhk9HKUGOqJGcCmE6GqeYz/rTW4OskCbjoSt6ylvJM/vvgh
UBEobrAxoUQ5GxFqLf3xz8o1QllmwAlOJwnWl8Y9FLNZWknIglkMTl3uj1VTovAB
FknrzLydcSY2QJWBr71s9nm3/HBpnHUev1zGBYs8z+HasoiGZUVLJttcNdCZGW6D
3Zsa4M3ECAJOlEjZBULFCHDc0gPzAOlA/G5e226zcaT58S88SwQcBkqfhlxWjoMx
EJkZH/t2Wq0CM7DAudtVXuYVo6zyQLwUJNltBYjtqn/u5Sm6hPGr5ZtmKZ2ib5xE
j31rq2FuAK8weGN+29/Sn7nKQmyUhZx6W+ll6fjIYQ7x7bT7UGVFlLsB7FjE7vAC
3VWmtglp16CM6LEvL0j2RHzzy0GxmvBMQYVd49gqAWw3+WNqja3nhNa5Dx2z3Htw
TTwRJwLzaebpndxKiWeuPhkljIWZZuwoFSk8V+NSsQ9qYpQXF4yRNryPcEDta4/G
vO96dJDvMhfrGdAIbzjjobBiQ4L3TuG2pM8gp8wPwQ95IPrpsqA7Dy3591mpbJBo
Wr2l4MB4/86s0Vn1YyHNRZ31jc4UScBp0lGyE+KAWULxiFM97wcpJaB+MaNfTIwo
cyOExEPd0KlkXcjlL8sqNC2yXXwZaJOY2V0H7AQ5gsLu8U4d3ZqFtuHx9AKVe6UL
jKJpqj1F80eIYG/47/4mBf1TG/yTKmRp3Kneaz9BXWBX6UVBV1N+ChhCFSlQp4SQ
35EewCBOLd2SyEPHWbK76vH8pbmidT5sh7Tw48hjFmTNU+lk6HV0j9i/6OSACYeW
vImBQCjd4dhiduRxXzdynN14FEHMLWcKYiTXBHcBV1ubFmVrK05CMBUiGpuEpG48
eqqOqMxHi+q7pP/cI0D8HzrqaaELVKYEphCbAthOFsfiNr2pFqT8bxGVXyjKdVvc
VPbe0t0ry3hFgATlCtmlCUf4UE6OhcYbSjEVYmDUXblRim3TmMZGN9Qi9PvUyXN4
0/LHlClO63xSfRXC7ojY8P6DhNul1NslK8N3dcjI/ZXk4IuDted/Q9cDIfoocmtj
ItVqry7IXTjnVH7Dl/KXK3tlaJWWdcb/td7P4OEp8nvWZu0DigXjaLxOx/MrLe3r
oTFaqmElNvBMLOoi9slfnHbTt8W2LXrrIWh4n6VxFDF1rhxWuJr+TkVi02uehD0r
Xkd1tmqIhbzaHfOp9lDWJ/oceQEa1McCZw3geX0dfG5YsUmmmpzE9ffZtUSjLizL
Sno9pip0f8SGl05GdH9XVqtpV9QsstKARVCzR6Iawq4KLXWb8+QH+DZEqgiaaRRp
x/2Pxs1Ar/7h32s+WB9fvY06w5wATaUNijygAGyzJPnobMzJJFtuLbP/eBKaNhPO
jVA1GsHYcm+CCPcV0seynfh6jzgWVRuubDcThZdXGSQyBeUvXGxwcC7ACGqW5Flw
wUgpbTgf/AmK90eOUJ2C2p5Re6PG3PqhzKhbWs9WA4x/e9ZSSzscAIR4OkUD8CSc
Dt3udxUUQ//yF5yS11rLc8ZL+7k4DszPAVxWBBR2EeVSCrd2KhhoSNdSkfumJnUW
JY8TD8JaujI56d3IBHzOncql42P8RnbTjLPk6W8bjHOWF47Wsz0iDA791WiXHlLU
8wjPa/kZ5Hw8Y8rvUEy+n/di8v857c8D9O1IeCSq5XeBqCHZNbxE7EMZ3sltDwcc
qnqfPjIbEQFr69GBStj7B63RmVAh3lKOfx9Ws4rilWQEMVRZe9EQiWpIVAOJ8yAU
M1J7ZoYNDD2Cz5wWa4H8LHXkBtFf4ExGkRt8Izq78XncCYYxbvTjyXZQ7HgWCdZQ
6Rfk1b3f2T0ObLSQGcnk7u0iWWHC7kCovaJZjUG0IpE+lxfJTKYVGX5n9y7twxem
ALc+u5C7Sc24nYcmtyLvU6Mu8eRfKe+97lytvl02l7NiTM+GFUaU41g/jZtWby8o
5kMEFnZeVs6FQiZfVstsmvVlECTXS4yANRnqh6py87AcVHHUj3gRzpCRFg+v/F6P
eNL6DLx0WNLmPeKx2gBOP/0cDfC5St8Y7DRdZlpRbzITl5DjwpilPSvAisz/YofH
6Vg0SIWJV2EoKX/4tqrFoYlk3uZj2U3Qnp2lrsC5ZDCtQrg0v6RM2NNWuH6aWp/H
e23qN7X9gB7Y1YmvAgFmwTCZSThgnYnmo2C0J05t/7YbpBb3fzwcOg3Zi75voXYd
tPS6EYavKfiaPn/Uy5yh/cv/cP4dZboLpxKJTGCJbhS3XJ+PEVU80dJIn2QPRerv
HA2MxqGt7vKEu6hR/RubayW4o9tFcuwsmYBUeY3zUHCbZDzSKrCk+fyylanSof7q
MhZ9y0sMBG6nH/2nJJADLh1id6R0izy50IhyHMejE+gB6R5LXWkiP5II7pGSoOml
gPRPE7TeBFRQLBFGn7vFJkM+Wo0/HMTWd6GcnwDtRwlrSUlPSksMkodL+DEJ9yRD
Y38UNDRU1gjs+hF/O5yuxr6TJ95HK0WGuF/xXCU+DKcBjn237DPFs4sHFKhfjDXT
eoe18Kc4NEh/tTM5nL0n+LiZXDmeeeE6pQndYelC1RlX7OrWn2YQ4fBGRr6uc1jo
IKAxqcm1oRyuUl/CV3YdhIeuL6RlT3aojV7feZypmFIBPMVWtdsUqu8VycP9Hrrx
/RNlO64pObAgQeOyXesj9Z39d7ufKUagUqj2XEFOnKmvRsMT+UQzcrH0OUU6gonC
UYyFrSeJxo3bChITTLkjkX+tsyh77vUV6HsJxtG2UiHBTgjeATrzWwjXa8hehVlg
AnATb5KbFU6DGDObiOiM4m8okBwXNdfKU89WWO8DQyZZnx5nk91iYEkp3ISl5FQW
1RzlKF8njhe/h7IRoavKEazD3zmRW8aWGlQ6lC8gtqwlk4NAYjBJqr4g5yzlv9Ln
OiYBdSTXjum1+RHi1yI7LIgImvjCoOrHXpk8uXgh/OH4r1xuO8htmfFbNKF8bUvw
jrKNED2EvH3+yQz84EiALRPO4t8JsRyAoIJDzOUAwmW9sSOAufeCuA1bjLm346Z5
ukLJjbUggMut2J85h7qHQOGIRINh04bEzKc59q/ujFf04VEzNSttBsjN/JY3hxwD
vSvgXf2vq/BOgH0jAkKT2bWbt0mxxuYrrX6P4ROMyR6xULuQuADc4Vox1Gv+gXvI
Qobevp6Jl5yO+19bS5p+AoDmyz/Nv1/qJFnYlN+YeO+1Oz1WmzgsabfD6UO3nz/K
TRWx945/3PJQ6qFUcH72mcI2DsX6wbOptkCWScVWk1KC3znkXJrcHFOYMfDmOSf6
/oMH00kH2+iPQBwbkx1xY7Mjwflbmj+aBY2BXuZpnEe0VyMDLfJWsW85yEiS/1pW
6FkXXm8CNqTf5hQbs1ov05Owi/RoG+I7Cfk6zmcnsck1RkRIaew0epaLz+ZMdyr8
Dc2Aw/Y4zeiAxWrES9oKE70N3jvKLF/+rA7rnIV58UplRpzWRbhaOOL8WcCGoMui
TNUUMB4Y6adAs3ggbRkBGGElnqRjOGtIl1VuLm4CEZy5kxgRpuFM4a/eMIMlgVel
2SRsegqPzEddovxdVpsN0ZDg7S2xZZBkk4lyJRx5xb81Qc6JlrHJAZ6Z1XRtjat+
hLHwSBqicuXjcsuZ+iCzOjaeSmvZFDktlvFEQ+uMQRgNwO2WFC5DirgEiB2+jsit
D1gIP+oe8yypDyadQjNv6qptbqCtmjR+nthlewuIhLUkKPU9ToMV5of2mME1rX2/
hWoXwYUVnSeUlldjiGecB+GNmzfpCBCkeFv2B7TL5FOW/gpy5lIlzdiCy9oxSjfH
GdmQHrEcbtX60jLgqnXyUPY/Qcs5A4T1Q+NEUsCSW7Ffhttm8dR0BMYUy/CnNJJv
Yhr+Zjxh+EHtmGKm87aQVsSKUXXgJBjFX7Ap/3VT0PqXUyayFzzkWN2CNIdBMXFn
9H/qckP+Uy5kb8cetno05VO67k2n12Fp2EKsvI+hplfO2gAizjK6BVSNijS5z0Ba
pYs5VPN16WcKbsoU7BbbbsnWzkdU2/j03q00+EaZO2fIpuPqTMJonN/ZpNnor7ue
IgiGurWwS2HHv6W/0gn1PgiJf9Z+qvMt/zwzV31Ydo4SQCmmeHPLWt0g46juwo0I
OO2JQazdRaXZjZhBT5x+Pr02cUupIqjb83J/cj6oQZL7R70YGc8EYTUNy4g3gKUg
IQTuvfyr6gJUkF4L6sGiR7um02h/7ndlp4VuO0TL6GEax9cSX+qnsWCwbhkPHEaA
HVmeHM1VVRv4pd4rZB0m7AyMJKJFEVyqJ0MFzhAMQEeaRfy4gfKbwEj2OmjSi7mI
C02Zcj3nx/P8SfSq2PGqbSwgn5AN5h30NvVvbAuDJImVQDiAn0gfqCClW3afMr+C
wgwD+eXPt+tPPs+MalTy/b6Z3emwc3pIRU/yMZWwr7077QVb6CcRULVQqMX6QY07
gz0ntdZB2u9pCEvtZdAQ7iO8xYVxEQEYIO9y7M13avPLmklrpQd1pC8p40gzxLzs
gUPlu8CjKWD81tyu6fuxmKbhzUHDHSxwfZI4HXq57a+1WgiIwCRVuUS0CSq+wAth
DTUQ3o/tMybJq4Ec7iPn7OdPTsXtgB3/RTdrdNg7fRBf0FjYevwkMCTtJRKJ2jkJ
WWXqDUUDcYgFc6rHCpDV5tPhievbr9rNZEehYwAB6TkRp1y6NX+YmrSJN/MK2AAx
V9Jqm3Fv04LmOXTwlFWMbU2Vz/+xsdOI9/c5gkwvRgfBSSLDoNZ7cOmrRk/fjV+z
T3RN0/r1EGd9K1wUUTEivJe3949FBoFAiX9MtevBee4u1XZh9MGXoKVylAPTkt00
KLDzct5nyrclaOrWRbm0oSK4UBUy5sUq9cpRrpf0HjAhFAROmudKFsmSUK1dhnPm
+dhUkyI5+B6ELW2QWWrnKDgBZYwWPMCH2zBNHr06e09n32m1yJwwAZmtiDgZUeBh
eEGQLOIOg1MylsaF9QO2chyprnCwKZJ6+9aMg1sBYj6qltH3CaKNT0HNZ49BMB6n
oGVxlcRIq1yzLAd7wVDsI+NjlCy+TvqX69subld1d6B08X075Is/C6+3QUB8pqIS
GdGAUtRAtREJpHfEkaBkb9kwfZ8gAVojamrXgeIfs1tlbyagX82dKgOfF09VAgWc
CgSfHif2be0+qbFIydDxbj5R5pZiFuQ97iDFVZx78m2Rzm33lEaX5CScudUn50Yn
fUQgoOl+rUd41gWClJIf4AuM6wp+WPvgn5qx1nezzCGiNovmhpCQONbfW5U52pSF
PEZh6m58bF937jsQ2ovOIKn747D9Pw4Lv756ER78WC4n0VAuql56lP516w3rxbNd
/oyVWkVKUGkEIuNQaKVCEGAKdUZ5PTE/jViEiuUE0rITMjVqDQyondRaFzX+oqei
kf17ASm9+fpXSSwfMRBH+q/+K/m4EQXZCU+jXMdoaPH6pETepRkVDF4DWgh/51G0
YftOFbBv6w9wIFsor2IsxLRJtLfh1i9+3qh2HtQ/NpKcCOMYJYfV0AnoVEzphoRf
fuZErmWunsUtbbYuIgY35j9COXuP5/Qpq+CEpW2mkr6JjyefFeW+WCNULqHgwVQf
YfI3TNIhrjCDUhgOLhOvZiQ9zDGsUEV2Kc/VG0WQR834zyJkqQmVYMubgdNKt660
qI0ms2oLmjs2CblR2ViHMHb58ucWCKGhw1LjDH7laKL9TLizbg+ElW7vRxtT6HWs
hP/qu1pgZBSriL76gEO8CsSyTeshf3FrZPOxxoAmxHijkFQni9algEg+c263ZhGw
UA1AI1XWDn/kMYbq3IoZJlZUDaTPoIQhNTph5xvlYeYid90j6CAbYGXLRKeKJ8+x
rVGgdeXkgcIwE5fiCVVLt0zBKqVkckbFHQiMtBuQyUn0A+u7fvfHAjjjvZw7vAKD
Nvm/8WblLXLxK6lW+XB/j2D3URZGeo18/2Tb1OXlUHZIUin9vYCnfNlaI6lPCtBD
cWe3GqUAncHXcJV7Sh4n1qwNnpfpmybn5TRPnsmb0uYkN6RPhqj4NanlmvcOJdky
q8iuhvZ0yJUkcJnTCrf2jaROSRS+OwcwRmYhuWj7aWwAWLe6pYByW29jP1bJuVDS
qR1bqWjKLQxs2PmiS4VI8t2+t4lDQbLTYuJGQ2Aviehll1Sp3ogmgKrzG9LJnMg5
12LlI8hHres7FgWfKTAw7d5MUYGEVfHW7m0W7xNdQWjDD9zQOEjdVxMq9n8RFo6f
AHfP3LWaEKQisQdnp21WlMpC7ZY9VfnXSfJInkMGLK8BgmOy74DLSFR7D8s2xOjF
cg7U9Ck10TcfNRAk4YM4b/vWl3ptsOpitNxsFzg5/RliZxmL4qsnNdWZBKzQt/nD
C3QxQNwCmhBiIDo93K7Mrcs+dUn5/EqGHM476AvRO1f8aG/X2AOM6+oId4jX2XBX
vfRgQyzTs85DxLpRo+OYybF+SBbiQqEigFF18+GJPAr/LiTo/XB3gDUrxRHNkXUd
3wRIUgILqHz57fNKtdFpU/S9A411y/Ay6qR3gW0THJpIAOLJXLvJmOESx7c30DlB
nm6ry7uBZzol+MNyF8yKrcMZSgu9bfFhb0z3R250Jewli8FpFAyfchcNCCryofmu
cj3yC5ZNmDka5dIYI0Zqh0p7l9UH/+6FqFlqbsRsdtmbXQSMRloiYr8HgoiIeScZ
Oud2VW51NOotAMpzENuozK+WkrDsWLfE8n50oLghKaUwkHWaFuuBKPWigPs8Lrn9
Mks1mZpWW9267/BIypDtBHxhx+JAuKoF5MfSdXy2RfTBvSA+RK1ixMkU+NrZ0T87
N5Qv/0wES3k1sN/8nxnryfqS55+MgU++2tgUyGDQrO1ylEJh+NvRuszsf581hS7r
yyuKdvJAEFU8caj+w+Kh6WSM5KnXVaSLvTFZ6WgFd+qAyvqAwJmp/NrETCtg1e1u
7PaugK9wmAO+1EPUCfnVQwwj2L/LZmZPVVw7H9ti6XXrNLiw8U3AxRjbgqdjyhQO
cclQ7Xt5rkmYdtgPsrklGb8CSckbf9SkBcH8ks847l8XsXzarlNfFSbOsQkD4i/4
UolC739+2vRqmwcEz1afyUdLKesekri/9/ro1Miivw4TxSOQESsk/K+JFEnK/Cr7
rgqOgGnrpeV0iwgPupfqb/l6DluMdCbdQvWkGcannAuKAU/U90PbIqV8yhqyoS1P
LH//IayJeXNyuMEO2L5BL3xXCU69njn4BzdsAFi/9965VorDyyMUGoLIOmaNnp2W
2zb8cOh3VkErW0W8zhUW6D+LKssuovMYFeeSM+tdvp/u6rNOzBnQ6ZwH7B7XSmL1
pmQIgSQ8qiYQqhUF1E1gJ1cLjFlQEyXIjDrjBop8Hpj4nJ2uLw2AAyt8u1EMMWV0
PSQZaV6SczqOkmDKdIOQQwsmuy0Pw09ZJBs5KHQrFr0iNg9BFsrEpKbKirL7WFzR
TGqREjYji8DCTWCA7G17hPoDzjd+YqQZAta2pNrWcc779AxmQrIQkJPJ8XmftPfT
gFe8d9QVkJb0uBrEl9dgi2huAVSau6xFqPQTUvSzX7ifWNdnxmy6zhCgxQHE8CvO
D15llNbv/24vvoDyQP5mcRtC5kiGjDMkK2BF7XyFvx2YRGP8W/Wdpczz2AKnI8oI
n2oWVbxK5EVig3Qdoe/Z/lpV34rn5GSAU/hrLaAktoKS+ZUN7SAymLqOtRPjCpJs
/y/M3pB6POJv08ai8v20V34CTW4RSwYEs/FfLB3Q43e1W4dc3NI6vFDvDVCy4CjB
1X6Tpo8aTFVfcHlZ8rE5lYkOy6ucZQFA9TYzuZPyKajYP1Pm3px1KohkVRI/f8x+
KiuU/koMGcstlxMhM1QPpx26PWY5kSm/YiRaYpD0DRkNur2wmAJW8b51Wot6w+xj
kh+RYtZDSD6C2R7T32DAz89/B3DpFEA8LpgTVwqkllRCieTSXx7As3U4qfAbUWdw
otcoMmlLinrRD2q+TfxcAbVEKwVj0Asgy7IIkAama/n6np+JX1mOEriv8tKjenbk
rIMXlde+GwAqnbOdeWEyOFGtbKPocWZunpVJUBID2eo/DBX/6H8EmoIQOQ5E5oif
r+E5beRqjI8fR0yIUz6M5DrEEcfAYdgJNC00/QKS+A4FMnAR+HxGsiF/M8DUrOJ9
zdIdc6S7Po6ksKR4oTNJhVs7FCl2tRwAuj7fO/MkllwTOk3hljvqk+ksIYwxtDfH
BgCeWqfcy2yTLcD+J7t5b5iSUQb+IBv3vbPhITNCIpUKMwLPyAfs3XhypDOvwrEw
b8fjcAxntWLND6isXr685BVxdtJJrVcOTk1ml4poyQafvCv2DAcQRdAKJluI0dsn
PG3+dQxry8EhzVQp/NNWy/ItYZJwLGwonWY33UrJETB9e0apHY2J34Tivw/1xZkA
25lZgfXHzsMVGY65qWAy7hH1n/0VgxV3TnqT4ophM+7Vw5d8cvyv10Pxk7XI4IeC
aWll+tBwamIaEYZM+tnx59Tc2V5XWFNTKMw8T6bjwoJ6GnW9oIvwLp/Le58J5G+v
TXPcp+Ybi2d+0jGOWqR9IjyCaSIiNfPx8aFAWjrvmuqxU67B/OkKycR4D7ffvLMs
bNnp3dZBKAGF5ZudRDUCeVh6TQxzalN/xCPKK3AJf5gYsH4j8SUxt0uxAuAKJkLQ
kzU96oZC2at6PfVMNs2IbnByJr77wGZ+TN2fkZ2BY3LEJ1xD3oizyub+N9mGsDer
FFslatMGPpxtbr6WAXsj1kFSKnZW1o4ltd5AdOL8COMm+qUO4rUXHe9FDuiR/KAT
zggzjBsaXZFhYLIGjA9tFGQacBATywouHp2XVmvCTQr7NxolXxIddEWd6yMpycnF
58Ajw2i+Y8YVGCbU2f5MuNKoh/RYN8A6aHaZ1trnCKJIjX6aXZMbOYIfR3TGfIuV
wl+mmRyDo0tupzNuVUQ5AgLJuOx8kPKBaqys+kWC1lV6XXKZDLNGNnsimWVuJAgs
l90gse/UsB8GpvReBB4R5T2l6/j15OfMRoi1aNNpxaC5+9/X8Z55dYbnIy6hrrea
OmzC5guDeenTF3KqJjxxOPwS+glMzNlDGC4Dt6g+pj6IY4xig+/lkH6hVAApAiYY
qb5VIJwnsjJnVlrXB2BgVI1tvgueqMDGiC04imYqtspQMpSrQdKq03tlscxkwTc0
JfaJ+0j8E982Oav92K875VCcR1RMIgbVLS/gy8Z5JUtjzYhz2yKJIWhh6WsFYQIb
RUcuyYCAVhn02YoqqGxBzgF1fgnJcmOoXySSKgdoxoA0x22CFWmUsrUBJHvi887I
CR/RT5Jor1J7qSrCI9UKGfLtC+DpajkPmbP8AhPhdQFY2e+eJjqUK1meeHBnWygw
IrTrymXQSgLC98bBKzZKOR3/3gA0CKZ1r6vrYlqQqIK4jWJ66Qn9MeLCyaA03yp9
Mn5Dx8KeOqgBELOiU4SxffqPtbyzssLkumSSfgMOB4Te42kjajZn6Np4iXxADsVx
w9DWpkBwyVPUmvJPOx02+qS1jh7ixSzzqKL3O5p8IMniKyYD0JjjU4NRuyz1IJHH
dfv+DlmzhSH1lGAJgYr4S7e7tSa6EsyTtFZWuSrSkDGkAuztnIrrFLDejM+F7cz8
b4knZJQtWB2IClQbSCf9cOqyBJ0LCQjX36+dC1p+NspSmkSAXGyRnO0qLz6ZsHvD
YOCNnxJPzhXlrmP7OcKQKOgml88A6KmrNv4finheDQRYOl2w6YiC1XVbSrox3ZlT
gQr2H4UGncF+EPL7TgVa+ZQcDu+YpsOSBqMPMRCvmkH7niexd3Us7yCJlHbqnXvs
IhiSD6uGFReNkzRHwUj3/++bH1noaxXFKoW0w2HVMrcVai9PodtVxNY4y40q+LQq
uXk343mG9kRk2MQnMSwMHELQAKehkUCAlKKfp626Kj2vF0J2+KwF1YPCcoNI2SnI
cGiSWreweuhT7UuXVsLGZ8W15GOSTd9Ito19OV7f4SN1cW6KHPUN8nXCsPiQxGFs
q1dWMdMJtIGOr0kZfVKplJO/qim4ys/T9LMqHB6aZcca65Gbua2SDcYAJOfF8XNh
Mi2/Tcx4s3tsJdxWFmW/7CpidwzTwdg1N+WzbhP+1oD6p9f8rY8xLRHjggLXeOD2
5ErxVdeXoba8B60staZNtHtbCc1ogiobPakN4bFed90xaskTBA8PXTyvunFIBWF/
Kyp02i7QE6ClPQohbGORVV45p6CM8S+2DWHlxaxK3KFnml6Tk0o9d0TLdshs8SUF
sslZCA9qDf7M+I+9Q+OwzL4cYCbV1BelMawrQXIFJletzUWq9OXS6gK1gdjhUxYq
q85vquEQKcoaJVyy3ya9J8ua3J+ySym+IlPyD3mpZzcrQpZzjap7/3Sb02j9UlUL
ZMyj5lGZsllBoy47fPJF5dSJU9pvsP0roBuAOmr9PvdCrBlYJ+PpiADg22GfNDcG
c68GJWkS35f8inl5w8kYpJXN73v298U9GClw9aiLlCy/Bt2CL+2PmbFc08zN7LWk
Ug2Psf9QP/eBu0pSy5rlpdHxXEgAfhoHzAEcVfoWOeD05Dw7nHpOYreK2489X9J0
df//iSOPdm8lca4XEWjMLFTLFuUOqLDM69WxgRo3xdqw0/OVSclGyn9f+N8ACNsh
J/0qWlBMrFULo96QWx/emCWNSndeh2YwhZze0IhQcbR9bfDZyC0kxAV8GhITippH
e1ZV6rQiHffKVGWvBFspn+qK9ezN6A48a+31SAk96t06+L3fAFob9AO1l1qG1LVQ
QX2bftcUcmQJALL6t8yzJxTvElVdjngz23EpGM2zV2q27wTYEgO/y86uHVHHkpPW
Yd0f/F0F+rDZwoXEBlc73fJpxOmfT5KUP8nC97DXGmxb9fjaqB6DueVTKpfmuyOW
4vu6Q+h67idvWsBXhQtuhsIGsiqswxuiLGLfcVAaieXHwczFzcNLMGQ7rcF74qmx
+csM3HGM0EGrTDi+Xiz5n3q2HA66eDdpkjEBRaM7yyWdk2wxwVmfzm/0ZtfjpUen
FRp2Pxw/XDedDSNJDbWsJJmO/NywpCc6SGj6dfGj1GH0r4fvJ/VrgZSGy4CHGUTq
nQfEdj2XTn0R/JCKDCTkvrlYmj+H94dWdHaX04rlQs/r8afr/VofS0t3KhU37B2f
ClUmweIbr0rZAbMX0v5pwfsA/MFNh2Mj0+x3h8laEy7vAK/iCl7BE4mhdLCLs6VS
Z7GTyWVcZDdVK6lCke2p/UtxY487Sur7ATKd5T3jPGXVYaNo4tqGzlGMvc+SAXPT
OImTI6D190SUqIGp5NnkBhYGnJcxPsjn2EpoLSUGdcf0Yk7uPgkA4S+nKJZSuOHN
O64wyR4yRU3MJ5q58AwtnZcKITc33SV5xjOUMZXYzYPIgTulrvubpLb3z4yISbUJ
8bMP06Wrm0zwWXKkz7w3I8Hb4RQOH2fnb/jlaGY/hukMgRAf4lHAoBSv3Zz7M0bR
FvZQ6K+lM9vR8D7OU5PfKKh/t2n8A1KFzfbzzMvGEf+cGmiDPcMflBz7Onwg0Q6m
lcwmVjepWWliM3iswKH5iCc+uhOpijOtqOBCvQLj1Wa+VSEfLUpAYPqZod8ucdSZ
QtSbjhEOa1gj+FdIYZq3WK5i+2wtqAuw/y037hvn1pmAdjWayrbi7esTPNhxz9Uy
WwmSb6afTnj8MY4RYdn4pv5a5GJ8oqLQOO6g7WVPxPJJ0gL8NJxPH/uAQnQzlx1Y
KJnRki/OoYyJJy5YSgBdAOVWlORVNsFI5rnDvxlgfQ+ag+ySL/szGIVMEtE1Csi3
OZn25EIpVCAR89R5yCjoG9D5bY1xJzU0rl6b1vp9+JYSZw5T7+5VtAiDbNSo2gAT
pKWsZIJeQYOMVmMamX9/kBJSZ3zSPZDdE2soky8UlflpTNpFUBMO4yrsOGlG9Mfw
TmIoqPeu7lnfIrxll+/KJh+jkeF9X0Qn34MNig9KjKD1qsZPSjVEV84VACqmU/8s
uEys0K+wQ+dP5y6lZrO0+CkNNBANCdTxcqONLUseg+gvXNYKES04J0oUduc0tjoh
sdXBDAFkTZCasvW66WuXK7KZEl9h4+WA+8zBHqt3vYm5JCF39e9FMjjhST06Djtr
l95jewc65bYgsX3vvijvywODRd4qSREeSF7fq2engBf44rtSyK1WfBlzIjk1GlPD
kd7g+UYblv4EFWNd2Z9IguVf10TH+1Wrc5antZP1oNFFTSNe8Wbjqdpy2wf8Uh5D
DQXee43/g5Hc5ppRGRVfTBjLU0s1aLYHHeZt4h/xoDRtcIAxurqanydDxRn2crUa
FOfX11NeHDvtDgqMREMjJ8o/U403yMnXvple6/dq/Vd9oufFU3RJZMiOoTDFL004
P6qlpkvjadICClVWaw+lYbeB+s+R96h47e2BuJZY7ovWKunnEnINawBKnmXH6Bdy
Am6rGIF+aKjWCjJT3iHFZbkq0MuY+tYqxFxQBqZXnovW4tmyslVeczQCIK0zSKze
XV+GdrphONewmSSjaN+kVFAaRbFUkaU4QjtRXFMT/khloMqaO8UR9GnxRrlqmbHc
By7pGkau0TFn3hWVqHUtmdc0kSc2H1llmZkq25SHG08aK1nRmHWkL2/qM85SEYvh
M75cQ4WFfXToJpDWP0NFin9bKnBwfHkPM/XVJ7+WLmMNB/liXjHe8nSCKIT/DC/v
onrSVj6hbEHwn1EGkoLnAl0j6Ce91n/6OoW7MrWchpUz/S9PGHz9PSV9gMfWE78q
/CXmr/xzdQ+PV8Y6tQl45xrtR6RAXlxiQo/1bjlO4Rffng7cofQPNDIWJatLGdyE
RskXzPH3atFzwCGBpXxGnYaN5GTcgP4SGEu5yTk8a8s7LwZNkmwwHcs+9Q4Vz0ba
2vPVe2o/VZ/NMdf/nHBK6mJRs0/shS6l2r6mVOJhEd4DFIqBwLRNCA64nQXgYZ3N
haF+NXWOet4gdYxQ79xYioa0Q4kk2EnkhSXk/M4i0WtWS7g5+JfgqUx2U82oD/5R
bCbMuV2hvKkCdSEMcO3dTgtMZVNaSVj145hnR5lKJcS+U6An9bKBf1Y4X9zWlbvj
s3q7xL5y3qXn62cBsfoTUR/TRaD1pyQPwJkPlxwQjtD60ye5u21TiFl8vJ0YcrAN
wgJhWFD/FNgRaksIXhVJhFwpSsVmr4b4TWDa3U4NDg0qneoD9Dn/oS3j4TXSPV3a
rtFua6oU1TsGqTErFMmfynCwDLlR/kDczLef9XNZSLbPfweTr8RcVQQolDoobx7P
RWa4t9II8dgcf18K6YuxsbIFmm0/2lwE4ImEY3qwPiNulhX4QZ+3GMJOwdRydin2
+dDwJUtnMd8Sko2CxsCOov9IDhfZ5zGWEVS+nwZpo21Ja+GvPQrvuPOeH8m+MCSo
c08yxW0h5MlPlPfaMQteeeWjeSfCffQEMKGPXwGyqbgOURhazAXwb1PfFSeLtYKL
YhcDpzWsqn57Ok7ig3wGqBR32Fvopq/OHGsOZX9EwtiatOCHNltPLcR1YwWwpTkd
++kbLW8u68VIvKYHttmLrMsvTj+HyQYcAgBh+oGgiRDhkC+EZo48uWdGmIIDkRaD
7lCdaMg2ZUXNHBuTwPPR9qHDj9TPBBp68H8NVQZMeFpS5KGYoSjGQFwBr0UQnkA9
gB3JstvX3lliE7BtxlFXAjXdciWNn7p96A+I92/Gn+pRtO3P6zcUa2W/x+xCyork
qbtpNVANFsTwut2j/KCy9WDQ7DTlK4AshpCepJ6Yb+t33nGMzCeOe/johjBg0q8i
GJ4OAWkwYNd9Z+guCikMa6NAQPkoEUh4vxZj+misxMW4bYTKd32z01fFSJMYLDip
lLuYnoEe13kDXwM/5jLiWKKPrlJEKYYT8nKjh6832YtkObYYRTtaINoPQ7YYXGgb
3Ck1BgNW4FTt9etfTtF18vLhPYugSPdMNoDnWKf0lJvggITlojthErucdw4zXogn
fMttDYfCPPTayWehWXPfyX+i/ppjbcgiwHRTn1W0A08D4SKdmD343ZbE5vfidqTI
GKpFe1i9vf1Ta/e5+Y6N5erAXZjjB93YRp3JFVNdBo18zpkiZZVMUC5+PS3n05KM
/hT487MwpZoTPKp9PVWPV6Y3Z7oNXGNj6QEXquEvOhsHLcMBq/5yHENqupMPSl96
5Pvz3L0acfmYYkd4nW1IXJiRAJIBfn9f4VhAZ5UoB1UfZ190mKd1OoqefGoHNlkL
JLBU4cxhyba/bTpjgRzX2ixxFd6VwAaHt4fTNw5ngGKDWGpZhRsA59mETBuFfYOV
VVu5VBs9v1p1bH+pxJMS7Sn0mx/ZYnMexi5TutwyVgnSzw2IcOyEjB7lJIE2WuPU
ZnNnOwp1h1Rb7XpGKquew3OfP+3e/OSotO2GfaDbPx2xTiUqiS7HsB+7aEcuC0uU
uUlonf2lR2G6/aJLM0aZ71WXjJO9V108nooXdyUmUR+aXFJIm97ZuSMINMMINyDM
AeWfP49NiN1Zh3a+VxA1uv0j3zSs3jvWgI+p8LPP84h8AA52+AhPFrX9Vfy7oZlJ
KkVfGLgLmrO00HSPI+wGnUtMEqvldPtjAbYrCSzgJO7QxOGg/PJg9jQaHVD/AGG/
uAYcUJdUrLv7Dxn+fJWwZ5uqTZgzfRgg05aT834IjF/7KPpyj25J97Uh3RniTw3P
umPfhyzsWvmDG51rAHUM9Uc/ubAp4IYeYM1jGBo7LC6NIFrKYmV7yvCRCn5gdFF/
mLgPf/qh38NHNEc8K22MS53R0fWy814Lqer7lYKdn+0bAhdHDEuP52R5C7oOXT8m
6MZzRFZutEWY+ZTkC1CiDNW8N3ZJBBjnEA4DZdaV//gDj7/4xz8wzAMMesmZmsqj
s1h7eSZHiwBtCAAUZQ0BNl2Z8KlY1LBxM/VJzPP3XK7pNvyUcVBIumreOXXmmJBO
9abx16t94ArYScPxQob3O596xf/oEKUocG67xViukADwxXMIBgmPhWzjwAmrHITU
P8QDAXFkfapzwm8DCPoJQBL+TJmzpV0D6Vhj4mnQ8jTFK0rISEOGNa1kqA9ORg8m
Owg/XA2q2E6Zv+XUThzfUbsWdNrxJX2OW2r45vzVzQzaKrOltyDhPat7Ul8Hfd7a
YfPZUBSRVoiOkYAxIVAjxj5qmDCr0BPe5rfLLGEqZFl20h6jTLs7DupgX/P6wBbO
UysWV/Hm/7V+McGumR5i9PiFkc0GTWqBMreFQ7NddwJw/FPbKDlAXagaM2CHs40p
WJZnW17mbkWwJxRx9svis0GUeVy1H+QcnuttgUKrwYOItTUX5GHATsRQXb0Q5xvj
sRJyV1k52Adx2MoYPgiRId0/K7UaUUBvs4psi/9XomOkHWEePfD8OwopnKLclZlp
6ps9po6WzkqBXQ0SSTAz22+i/Jv8jmUc3tswWxfGakbQyer5OVOueaX8xginXah9
CDXviAAF+EmsP1Wra3gV19aa8O4enA+YXpPwZrK1wWl+i1qw+P/pxMJ3S4rvWfwr
1+KbgqOtG5jujRqgPcFfSG0rvGWqefwgXI8A5atqov6+IEalL8Gh56ruzlEQvumY
ZzmTsrcC5zq+e82MZWRhdhB4tgGrFnBNmMkdD5rvl8RVfFm8FEg+pAe/XeaXPIwb
hfnNuiAIXoogxW9PETdeW1BGNT3WW3fhl1Smhsjc7Ko8REpMrOP2WkLqbIV7qkoc
u06xbvahvNMjhDQvQ2v8eMhOPGTSwV7nQFeiyk7ZGzHfJgg9NcUHpxW0RovNfcdT
vMSioabkKGtNOWQydRGywjEncNJ3U7HQURgWeFpnpUcLLJuhRzR5RcWqZrIldwTp
fD5oh2vTH757jT416DcVGO00GyO1gp5BBC+aKsL9ap28B1P+h8+6xtXkXonCeLY3
A4Mf+6cDufJaF1TciSoW6eKGkbOrmvbDh4WLYvJAn/HpHOMOd74IjjkozujFemzx
2oG8gTpiRi9CLPp3f+9Vx+rcG2kQ1tLk40VE5AV/FpQf3T/IJU1yaMbe3W9L8n4N
AqHVqKbhyaOtQBGZO8KlmLgUb9Rl98ZpLCyWQpk/1CIrIXAy6x1VBmzL1aQLAbFj
XNVtLFVn4L8UJ3yIacXnvkQXcCME2/2t+72ja5Q3YPsyY7t5QUf0KVak9YKafSlB
c3MmCFvwBJXFtZHthWmZlAXNLIKUAoB+sIE6R8kSDH156z6aSBnDXJXB7lFz6lxJ
9vDpDuq91j3BS9CGgrUD5GGPk6KqQp14afVFK+AXslV6zY4Xr6RiNI4Y1TEcxn1w
nx3t4g2unQMofDEd51K2YznTQRAGsl6dGc4jni9d3DurBaENQ+kbENkFFhVNpCD3
CDyuKhoo6fpc0HGTpDlWeqV0of9iF3zys15zHHUl9TBXfBJ18OEFbYPvIlzUAGiX
9LK4Ke//KVi7gmAhfnRg2qMTxQBh04dMiigp3jdRMd9RRujV2Btz7eYEufAWwU/g
vDyqdwZbzDfh6ic1ftH/iaOOsiCg69XahXkzhOPV1m/M3nlwaKF3vz0Lo0j51jVj
WgKhwnH1MCBWu7JYNXDlSoFpiPP4jNuC3zGNq15mN+dStUzy3Q9KUBv5+SVj3awO
FAVievqgMjGyhC+l/r4wfypok5E9TZSUHVbPyjVg2XvO8XKhZvBblk/R7HOVUxm0
x+25e4R4dSHVpoXcgWH1DUgXfNtANkJbK9wWpFgVnN+roJszPfwBfghoplTpbtP7
L+DWpQJBvHF4Abia6/q3zmXqzK5PGS2ZoNNac+UlysCoBu9fcMmYr5U1xUO5rE9k
P+dFlCluija4EXnWrEi81664OiNz5SLlfcPE/oKGg5MXMm23Rs1FjdlzIjABeei4
fKNfbbkqCdhfU/SvcLOmKrt8cZX/VEYf2Oya8AzJx3jKvubtXwYC5+lGYsViJlSW
y3M1sddceWQyFxt45HusvZ9ahH57/VpUQcH8tJPOzIHD+I4Ijbk7cjYYmZN9iv10
BTVa5gYmDuFojMB6Q6cRDsTFAatLG58J2Zodt06TcPLJbDAKRk4IP6Vjl4/H3vWp
3divvY+GSZ1lG7jXTwXh5dGTOtpA1kfL37go5tXQco9d7/AXOAKtH0wawth7QXKg
lWacozWPzUSnXK4nSNiu9izNqXi0JqRFCR4c/N9P9WpHQqgs6pZnqsMf/BZFuhdr
n+IIRWur9r4cyPgHAFNnPjy/kLXxJdPeofEv9bfX3VeSzZloCAPzWrfTw6oziYyW
c07+BjojEO0jLd99oWnuG24C9OHT0TyZZAu6hZNYQWJ2gtsjcyYRDJUhgcG6BHGx
Kbnlh23D8hbjxeSkswRyrBCQmV2fw15WgjlnSxftwPDSMqVCsXV3By6lookRbSYB
RsLxLRXSoVOb0+HMFucQCGpGpWSioQkR5l0ISogoad5Za+GuBDSBakuLpGdVr9uS
cCYZ2qTvS/4YbFuBrPj/BwXn1stALaSr78dVjhfcPa6o+DA24ixfJ43unfD+01ON
Q9m7YssrBpKXtNmyj5qmNbEGpkrSJFf6TwIgR1X29guah0SHQkHH7B72lguVwc4K
++ny+A8moL1wBsTnUiwLSgzhYAZxKTqWN0BMEWQk4BhYr3ScWIgJS/5ZI4nj7/PE
As56sSZVmgBhqETVmnnWssw2oMdSvbshFOR6xEZTDJa0Zf7eDzcLBsghi2rnIg09
Y7/g2HtHiVSiFSZtipOLyOivnGTDDdbL+YbsyOaqtmkmuwV0vHS9zDsy51fj9wzO
n5qNJEPkrVqts3V2MHpw1j+yD/aGrB+5eJ2Pm4ANksj6ozUXfimRUeOC+GZkHQcW
g/oLL8ajeGseA4qBsnS6iFrF8gWx0dnOqgOatnQemKKwO0Mo1Z7tSDnH5hHZM4Er
fnhFMhxdgw0/FUdPYVUYQvOJuyP22h476LsWwdBUDBxpykt1VIMbtBhe8HIIjkK9
usMrYSx5Qx/KxtM7cOERm/18B8PxbI7fs80xZhCmXLO49XjWYMpB/l+LAjfAEPzX
kF6aWxpJPQx+GHTc59rKaEUNoTsrXo0/MXTuTCIgxdTAqzFNU05+cAhXPttX480G
t2v0+QAqI6ILj8kARbJSjLhX5qwKEaS6Y8AgLRtVBr5OyJ3gBM+TmOXzhx+B9vZu
5kGyiamey5pVlWke4exSqlJd7aPx0aXFrAaSQdiMMJYLIKL3AYw38qen4E3/aSbC
EbFYU+/zNlZ9lm3l2Ztp8y/mihKYKRIMapBduR5WgvrJmEFAgL47Jx6x/FZb8G/U
mAhnv/vnRNSDVZPVhLiAMzq/qGvNWLjUEE1yn/0hWxXNR9k4LHHlryraMJ9Z11XF
XRo7COJUqJO6VVm+lLAjZkoMn9I5lvro1TMqswyTsED9P2EDi2yBQSfzitTI7HT/
WI+NwIc3SkhxSHPIJgOnePIgmEZLf7igNRUjb/trQ31AkT9HumRpZa09ZsYNidpb
L/OiMKKXiIBTh3jSX+pm3k2a33zWGU00/ZrMxuT6LC6WPVW2ADp9rIg5dUX/Qt+L
CJTTtSuNcwwhe83M1J7hF3rwhJeGJq18TDByTHA6e7jv6M54tNxBM2XdYNhcRJUc
JUfeWdHwMWCFd6qXK/w9SbQiiQqJP1AX5Vj8Vs66NgzwjQZBxerNdCilWLGtTkZj
In9BGsi+Qod5JauD9TSAHdGx6OzgCPy93Oi0EcnBY2d6gGOlE6++IahpaGXSc9ru
4Ozik5mITJ2TPW0w4Mk2nhEIh2rTd9g2Q4NM7hJQ+anmyJX1iw2fnbvdiqNXT7Ct
oyHdG2DV+aAiGsgH2WNqLnLpRPqoxnrbwQsQtCib1/dtEnsNmTlXcOZ8xLudd8HB
BXDOB1sB6/dIEGohn0IVNjO08kldJutuyg/C8Cy6PddW1ZDVw4RqYCR6roVEqWgB
hst3j/odss+g75Bg0ghlgsjE9go71qry/jkGOphxwXq5TCoL/kcs9T45/t7xQ6mr
rbiV20LDn52S2FtzB50rieyhAMIS83lLvp6gH8KSBaH9nw5l/+B9S84Qa1d8LP8L
JvByI96ecfXw019pwFyLt6TEu5/U1cCHNbvjKBl8zAiUp1uOhYHE8xMNBB5m+dSJ
Ru99GoZe6v3/6HhkoVgtJbLOyxupRl+qxTSzuN7Xyzqh4zkNLEROeRDlDH40gNfm
57KGiUWcbng982NXW/u8ogS+nS4OUYubPqH1H7KWRdztsrWksAHwpx4vEJY3uheb
LR7g6okcLbImgfYXLL+GcxcMFHTs52xgChxtdvDX/osvGBz4jPEAUB9XW9l59ei7
t2eC0AzGGsfR+EJOdRF1ikQlSgBi2ppO6KSrWt5f68K/cqngrgCdkToE77JZqvMO
GBxRlBttarA8FkdsvCGr2GUZsfSTiJFpqNKLJ4/lKnSS27k4iU2Tn5XhB04VzagN
0dh/Q+nL+gsoBXeNq94+7bCzR4orFMc/rT2hAyHgusjKyht8wv+APUrod+mRkn96
+zZK2y16JHRAFABAUw4RMRbM3hdWsLaQlFzxWGCuoTRxfLPMPVgLN5yTXMK/5Xle
ltLHVktbyX3gk4q4vGOPVugVsHamXYcyxM4vM9LWy4+ileMZvCGAs43YVq3lbdaQ
SrC/yU83fS8x3hbT8XmD9YlvBEBIgKYKTHwTtduCfvuazmhlFCG9iXkh4OF9K7t/
lfq7b+TuC4DUsEu4JDxirH+Mmyd3uQZczjMq4ToGt7KVF1bjbIv+Z1wTzW+1sPhQ
piRJRYAGxiyy7lSwvgkJ5mArGqMXXGaPv89UNRzWjJ3u4SPUPHPSGsvWn+WKWKtO
UE2wGYE5hf6/TgjSFwn2N4nKx8pN1ORjL0PkhuV5hK1Rx3gNzhmW/ULviyRTJO70
eu6J2u+gTyv+eRTRTWkyVxi7eMl4tUEw8lhHKAh1eesZOm9gev+iEXVPjgaCXGJn
BC39YVRT9sle8wE7d6DHg+NbHfmELa843fr8hrRNb5/MgQL+FJniAmA5zM0XCmNX
/klM/Iz36PLb4hhdidAl4tYrIYIUegQN4QzgivxDUOnqxLT24VJiiG1xGusXzKj1
Wwvge7CyBkd5MzuvO8TPsYchP3ZdvDWOu2tt7QbHrbS1ocoi0LUXdYQnpZsy3Hn2
RCdlF9JuEZdCtNzh8A7RPb8la2YbDLuI9KY2T9RhqcddjNpfRJ2Pk/UhQym4fSBm
u7cgfMhA8O+S1JvKoNKaPyrHVl/3iOC2pCek0ui0JSO7ZJMSoNKeEg89bXxV3AIY
mQnz1ChijX1wRMM5l2Frs4jOua9ZDRH/WNIwOvINpPV0tDOBwA3VGkCFXSYrlwWh
STveuS5mO5wy45hhlgR/qB5ZqNTQX2N/8SyBCphZLDRbrM2DxnnHpo9g1Jpv5KeN
g8I2Abzeg3rfRTjuxeVq6oo8bv8vz1FEY/Ys2WPej+3f0ooSqkHzqrNOpR2dLQTw
sTfD+SyAQIHkfXBS6X02fPyqhmFACD4VcCE8ahjZoj0R58TOXA02R6ztocTr989k
gEQ0hJ4/NsQBKOiDQicdZPapXmVdjLdLjKOye5NrDeh8z4MzPxbmPHk6EYHBvppQ
NlY7VNykzWwc/SGv9W7ELy9ZO1AIK/eTZ5vEhk11vHTlE1OERf4McEJ9xtnSBeRG
RyLVP2TjdpIozpaVj0fWMxvxrbqLtcXCTHAj45Wphb3CE1wUjvlRGb18CUZHXPuX
BM+Hg1kBmjB9UTyNKkSBjVAOgUo/tZB+y9LNL+t88MnGZdQ15BBClHvr8z+pP8Ny
ph57V36wgRX9WJIr7cu/64Cc9MLzZxVa6uLQgCy6yDNAAF4vKRk0rOTZzXm8dsnQ
l+SPqg1WLVWGSxoaF0lIEx4ogWiQBR5VZ8TC8PF8RTVw/tKwOOAP0pwGWHgBFDoK
A18Vbi1XsYi2VrPtf1qCXUh5FTEqENsi1GXL3ZEat5XfKVqat3DtgUkJKoeaTn96
Isih2635ZhK5aEXAi0bmltWqH1Ga7leYOOTPl3ptlnEDPiaRZA55bDznPj9LbXXu
L6tTpVggXorSwgJIXsB4u0zSEbrZLaeuSrBthGSdIqV48BPJOOgS4a61lfvkgAvP
ZFPhJHpdf954kcS0ebeaAFwa4ZAMcra88QfTAz9vTKs/JVyANhxRfn4R+3E0k+/T
34ssnBL3aRMY45XnUeD2+dHLwoTeuH+nABeLia4gHUfv/l86bT02db3EEM12S67B
83xFGUFWxWbDbEnPLO3J+Az5mv2NLReQ2cL2AGEf3BH6R549CNeduSvdS4eMrySw
1hX/ZEGn7ABrGYTM0qRmO39Ef01QlNqYICk96nn2b8vZfqGQzQXygPc7No9DktWV
ybh1lU0NRy94SxOFwx5NMIHh9ZaviJMWY35IP3PMpdZeYicvh0ydGLhsCVPWgjl9
JCJrwrSHwGswbCdG2jSdYXYixT71ZI/gBS4jL0749ugpDpZaZ9dNx7htTY5a1T8X
3RLEqx7xAoqRlt4dYdP62Fsn8ZevaluEdfkE5jQWa8SkF4dIMuwIvTZCHlTLMxpo
CMeFsbJmZYzSly+PNNeHWe1Qi0+bf6YszYxiA04Txhu6D7gYGhJ/5GqhJANXItS7
VGZlfFchuks1n1M7Q1mvdNlOgTCtPTl2g1nM4xJHz1Ti08yedxORZisGeup0pqyL
LoDHKY+ZYKiQwhiHRCPg4RHN02af573o+4GPuY3vWggxoNUBcqerxOA2S2PuOYMj
C7egaEVIbxVz4/d/Ja2lydqY+U9InrOq2obuhN7rL+vcjWsYuO4Jb76E2VBdCPT0
Xkn+iqo7APq4+i2LW5C8wuYFWkfqD3FaJwlnVJ0yRNppC8m+4w8TYGfx5+bKTUnC
A6W19RFJmagcP4j+/01zoRpgJdP/+u7pyGuFK+GampnO9+Z5WAXgdSzOaeRVpQu8
BH0zSV3eMM+HbZSVnplrmO+IyJ2ZCpDvC9gvLta6wY39w0H6KO4CYE2YI/mloGYH
8aATfuMq6xnzGErRcFMi8UjkaRpgl7LAYBch4AEujdmxwl1bTvGMTay8YwRHY/Ar
NnBK3UTV4rgVqB+8435/rYMbnxBIuwu3KTIWNlzjLAKlsQDuZldMK4MDhBYWybJV
EY3kAFlsa2PMtdzZ/VMTePCFFRg6dZ0bxpsA7r9XDOaGFryVKmEczLBMcfTLviSC
KuNu/H6BSZPnTWF8tCbjBRpCR2txlCx9WY/B9zIK0HFWwgll3MCfijCYVC3z4u7l
/P/7oLzU6nQDaypm4g5HvyYk5RKTgEdXrG+OuPBhC4l55gfLp1guSMuyzWUeOYya
7jtmLlYwTyz43MOlHGoKS4s5K95bmo8KGBLIF2HDjMdtzqShh/mh4w/KSIUF2vK+
E5Omz4PX6S8+wmPBFAiJDXO1w6YoHG/jckSjjSHVgG+HwD1Cc6iY6cziZtTBOnqu
46nEnjKA0eleTj8gs6aWu8NbiB+xXh9FUSp5FCIfZAhtpcsDy27RVx0ae6Hm6Fdb
7Xhr9a976RQDhccrkI5ns3B3LzMfEc+6xpVoonIs9FkojXwNUXkxRW0LxQ6SC4WD
3MZVpXnlmJ21MXfnHCnGDspt44KfKN+J8TjLfqxRVMtMLdRllUjXHppZ3H1pQyUi
oUHWgFs7SmclXDlfNU+jqhMXQWjiGO4BklrpGpdYEN71vwOq6oZMslB/CW6r1j4v
H/0NWJfCm0lSi2/Dz/FlWas1PtdEE+lt4+XNM3o+4rXbzKCCm+M/qyREmg6xqfW6
VnzrH6l6/9KuK5llMiOtXauifp9+AQCxHqJCbX6yNEcB4jpXJhX8tV3vJG/xF9Ta
WrprIY+bTDGEv10k54X6PiEHi9HvpBmtoPy81hd6u7ikKs5q7Zuy2Z+ROkgE3W11
b2bBpHEI2r8tLO6PiPmJ8UlLSg3fj8ZCoPxKjXIEK67mPBELSYYNAdA9Og5GrZeT
w5Bd9kv59cPRykAC+jlszSFU5hNj1G649KsMeo0z6K3qYlbB3IbBAlhRNSiCU+rn
KFIVLqs+15Eo5sAREbat2TmIhqhHZVuhmMOC6KbHsp8E2nwsgpn2OWh9S8Gs0yRY
mH/wnGmAuKcLzYd0X/dqzNgkIXQMT8fJvsFZuGUE1M2F54shudMoNjzQ99k58RLI
JA1EhCUWdtFB3NibU5F8kJdb6vHw3w6aBmtPZ/0WIh0uO6m1YxQKoqtxxkOZOSUI
qFat8HMem23AscIkPPdOzEl/AyNtoNAl3AhnYa1D53TINbk4hs7Z8F2C8URj8Gxt
P4boOA0CuVk4EP5VdCoK+BHNUcILsddBB2dHdOQuO+8ddva+mPL6oaNQMSr+Dp28
Kmq0ZV+SsSGjGRtK/q1GMPFrCw0or0+AC3Q3sEus7HzVOQ/n7SJuVytoh9A8qOGA
vFiTFWlv0NswJWqjXqB/p7XO63kRRNDpbqpOUTHggiMdHoC33uc9ptwsr6dRDjwp
i7XodKoblZyJOyK3/Byu/KhOqLtxr/kTG0PDIi+eJylOyMh4M7Mtmx7N9RGAjYgp
9NLOL1bve6PoeBtGhyfJdHDphei+8OYfJGQTwyb9gMckhRWjjjNRaxjCHDxaqSWF
dgMdcP2S1qbjwM865Y1lCrHlR089TTg1NuRSW5kQgM0IoUc1KlV4WjrbCFd5aYCh
thMgEN4aaCgrQGsE1kUHXjgm8Gn1UdSfZ1yaPtWQz20r/bsYOLx26y0+m09Q1t4l
lcKED11J2dwNtrj6ucBfT72jWDhnZRGhbGzl4RLGIrnE/PVPzVSnRYJp0v3U4EfK
CDK/mWiTK/kTDlue81xVtq1VYq06Mp6OZl0fwCfFr6jau+ofQz/uYrfjOl25b6Pk
QjtEnttIsf4vhZNOf88P0xFZZkxWnHpEiw03CHTGGCB987Knh8Ji0s5Tsbs+L4dp
2tbqh4tWICEehbdL0XDfnyvVpdgJGNWYP203J5fBXkQTo5IM5vH+IiEe7tmVTlR7
Nzx6fWaiqCdFBvSL9n1mUWNh1omj/6TWl4tdOeq2iFA45Kd4wzV8S+Wj0C8Et/YK
zYQ0z/ALg9Yy2yzHTQz2XgFx6cLxDSeATrLqL0hiRTv1iogVvJAvxTV+YcHUiGOH
G6zxHdGXv21sKS6IPAA1H2a6G1LKjZf27XtAnFvo0vdUgyn22LqYCBJsxmd/ILxj
H6Rhr0TceznCiuyTBPkpotxTMwYjA9L6LFDE4AMXyR57GFg2USv9TycSVhOFm+oP
mXNj7QNqXzLxgL9tIFMHwotRcDjLauMbsDWPj96idE1VU4ekKbS/6f24e2ghy9xR
uHck2oCWkNz9TadX7oeFTETtjcRTY+H75HMBOTd+WmjKAv91/xx+0WXe32oaGGrC
`protect END_PROTECTED
