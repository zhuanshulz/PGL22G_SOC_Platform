`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2XYsYXLk+6SpjZWIMzftfUilJMM2Jo7P0bKC8xZ51T7vggNksXXTic93fKiH3rNS
jAWlA177TTeOk4mWpZiXDYIkPYKwsDLmdH/j9D8Y3xQNc/0WdQ5G8KhESGK8sF66
WgglLRU/ZD7/hk9NIV43QR6Lz5ueBBevwUnUyj0q4L6ZH1UB4+nbhPunIZZTXyUW
PhL1JKrzt7ibMcSozQWaCeF6SdylAhQmZeMRpQBfXHysQxKpe/UqEuA4eAzKoMgA
GnSJq0lcam+aDsl4TxnrG8XcJG7IDYXLlC4NJOUlk58XsDR6XAoIvVYJ0f5LN+aK
bfrezcM1JfxWMmlWJiRo0wbgkyt99zVvj+vb6ectnKQV8D48lUE0vmkz/JeZM9Fb
NqzOC81HROLVzkSnZfC39l566dYTWQHtM0E5tCMcAdYgq51lDZJgsdhnZAT4UZQW
noJNME+XtiqiRaTLtayyyE/u4cwNd3nybfwmIiVbouFNeC3e9mjuvS7+sdVdMGOc
VnKCL9cX/HVzA5mpdk/NE+dQhapWwW2DGxerRoS/rGkks1MS3SgCZLSBmnoyLHFk
QXE0HNvGpxl6T0sT1H4ERK4cXnlskYaB6l9zzrBK7eQXhozDSoGIOH8CG+yzq3qB
1hm4g+zOfrNz3jmvPC9IWkzGvJFIL3iMtx/tiF8JtFwqDxk4b1xrm0MsN8GeaRw9
tNh2HleDnuSFfo/z6ZJaLcSkIxdJyQhW3HqL15GHawyUz3szd7FKcJw95tInOX7h
4/+EPBp3KytZ2z6dVyOU0J7NJKhtSGtwZSxdyfZeO3ePk3DPakTZAcaqtQpL59uD
5QrydFq/hKNX9dhgUmb1/IxRToPeUiKAs/ldEqLn5GsZcvTZdgMvm/xGUYZ4hwJi
9Yva5XwcwHyeeYeZKubGFVHea50fyJOpzT95WOxrVplRIKRpZ+PjwMUciBPwwzJj
mB11nSOA5BS+xU6citOegZroPv3EDic03BXqtEL7/REYTBdsAfNboFfY7mLVOo9X
dXFcT9vKJZxDxli/rMPcilC1yogPAKN3ZW/eBc6OjZjG/2WRhlIzWTUc93/L60P/
hI3cNffBUz4PBtRZUTadxkVxVADOfnjb8ITk4SdIhy//xSMNBkm5yB2RISjhlXRo
1cW8i5eFuc+mShr8gEvvpUYaRmMVT1+ecCQl78A/zZLIWaQZ2FBlRuK59tAFTKhV
7JYILaRA6lNt0J26oqLCOeExGJu24pfh94P1oEOBpbLBN9u22jnNik5X87RhGKgs
a2hiHyDyYU/FO2J4I8zZneaPDjmNk9jgYCZy2kREC6zxx4fGGUZPlSegBf8N4r6R
/rEbDLfOIEDHNpkhtMkIC21VsrlqqlIPEp7WIzGBPTPMTBgGjRGXNHWKFndOrYKd
f+cMzR4aKhDgH6FXu6lRNYDMfk3hz0wgnY2GSKRrJM+SD4pyof0bPLe41cGsIHG4
DH9SZO9v5/POCLIWZKhYxQ==
`protect END_PROTECTED
