`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tt8URNIBdRazeJfeiMBvtfRcrCFLx95/sBxig2Gb3aqezoU/6nXx+IfUF+RYj/Ms
mee/rycRunkQ+komqVC/5eZ0KXBCYr1IvWxLEVnyCWEOcTWzjkA5Y5F1tRLOC54u
xFbKn5I4ZHq2CjzpA2WKOkisoPV7zZ9NfwkaiCaK+Sj5m1gQit4sonxq1QHfu1V7
dFN6nVmLfKa26AIYY4N/suqgK+yYgWWQqCHQRy/2HbXPSyGqky4pYIowrBAZrjAC
lwlyN20kOhHB9hjYqRS0K2PlrcVMoJI0RJsVtnR1qDBi2scR2OGz9tZdjH2xw25D
baCGq5/+AciAOaDb7HMj1Nd28wkyJgFVnQG6L+YCpHQINChHWwKs2oPKC7XzsOzs
CyR5F1sIGTVqYFieFqz6Cl5NYEM95E5yr7rwA7ip35ztTLmkQP69Nm/ckATe8PE/
2zJnknOlbCpy1cx05m6qcJ/+hrTlf2Ug1TLG+CmXs+Wbd7rYQd3OOZlw39zao9WB
p5UCOYsDU2rGBB5zo/I74Z00S4jXmzYc0uRVW8FHxfvbv65dd26KViAftJuFk4rq
18Emy8Acv86JeuDmQuTjb10a1/CAygwHdVO7y82YgfUjXzUmV54tMh4yrhKBLEbr
AvjxZ9LJ44ESpvA9V1+i0jCCuSCPAN99g7ewJ6u+lT2jpWLV4JPmOJIWRZMAp79C
1Uigw6Np2yasy2OpU/q2Mh+EulDEHReGEleegi+LOyyWqmsgwX3NKim4gLyxwUGf
Lg0HFVpOTYAfB/YpuOgmrVHTAGdg808dfgJo/24xhgOsLEh9CA7rd05Pl+VF1B/W
bPcwhCnCuC5g0UbQM6Hmj2tqjHVAmbm1cNPqJ2A753FlVyZ5A6UUSBbw3M+TtDd0
+f4MR2BQB10mR5Oa7Fr5d+gGhyR+PwYPtvJ/i0/VOXs0babxZoDJhw4a4vY1J6oF
H55vO2co5od3dtcR090fW7QMK7SuxI3JRi43NkFgpjArZULAeMKQMk6RyZC+KYeT
ysTOcizz+2F344vdD3+DrelXLtK/E9mW3Gzj/4RtladiWLCcvOj4bSawMwSZX2V+
sxw9DEPzlsxo5OZI5lGSC/4LToIeMrpiB34vO6/82xMXU2q07MNvnZ/jYYlEhtuG
c5wRhpC4B30LJNmZvy9Xf3wGVEOxOkZn8sXyklli2hid4SUsmkM9hI0Omjv5T6FI
zVpp9lwPa5u44H8x1mS0dXzRF8ayHkg2ila+App233fLsS9E/YzHk3GDLwlWxOLR
`protect END_PROTECTED
