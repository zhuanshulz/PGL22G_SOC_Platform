`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G5jFxB3EFr+qEb6PfXdfFLADvfFqFOO4oR2B4zkMkMd+AHbWeW/CxmqlusWFDWHf
FsnnDDzpgTr3cWCXeWqBJh07Zy6Js24CH39ICqRxr5OkdDx1Zy71qdWPA0LJLSjh
zhxLmbi/HkOd0fLeUWIH9evm5JqFRF2oaP46WzOBFXzVZJQLXCDO4WAubf2LXL5l
/axetywXZ3t2P2ABxNQJ7R+7yz7bYzxVmkh94ABD/focpmxUK9lBT1rkeNOLeVsd
EuzqJht1LOhX+ONWFlf3yIjzS8zgv0V2L7b2ezmYAFe1PkPlNyhiDYsUs2Oxf6pt
bwLzSSkokA1K/Kgt/1JHtjrnJR4oS6o/fPV/vOmNtWxLgUVH3zr8h5HdmegYK+0u
r2Kp33yDwZFUPqslRlW7ApL4RRA1+m+FYF9QEdWLkKd3Y7cRpxQtj42ZoU3MWZp1
4xVUCgYm0OXL8W2Liz+CTygy2w/F7VlDW/+Dn0qevL00A7ZM7CVwArbdpoPXwoNX
FNx4XgI18fvOqXZi6LVyAwPfv982PVMeLh7JeBaFILIfQKswO3MwAh2nskzErlPX
ZvnnxcQ6RGgKqhEv2EOwOfPqn+qZ9Gjs2jvPL4bBk5ckozthYtl572bD9u18nwRB
DHf10GIohmEYdWRutc2/rI6OI/dXCr2ADpLtD9VTZ1S3CL39KnGo75XDFsaXPdDn
tSCyY3jfK6KHq1RW/cwfR9I0d577OKraBJ6DJ/LkWi3/BpPlUlao2SxItiSquMFd
AqnJJQ5ArSzJQ4XF51e+QBtmRlipujnQn3DLq6VamiccsYHFds8EZQLkiQbU+FZC
+UhZ3uUfcigk0t1pjn5SwVzwFAuGKDhZ58zmdj/SQEMtGZX/uyv45CW/Qauq0Qag
c/bmDbDwMtaKgdSCUP3VRi5iN8YYyF1jEKA6YuD4NtVPF/3iJfMUVGgse5ds2bt2
G63N5A//TMYH8hR9fr2SfdUp8TEjvFVqfjtgZtAlGI7OwL0X6iKBYxrCfTbJvOG5
Ej8E7nC5oSxeGr2H8CXqGkPECqZB2KNZ0hZFW5sfBqmhazCC7+xX2DWpYMLC7Z2I
PLMycc8wDCEM46cY0JxQNcI4sGuf9bgBn9twgWsbclw=
`protect END_PROTECTED
