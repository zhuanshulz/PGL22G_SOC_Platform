`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AwZLbIavZeG00ExXfQZAtu0uLCgmhgksOs/eL103W7LzIWG4msPq0Tjs+h4MJ5xL
61LJV50Luja84tw9WPYYOFbnmhLaYRMBXZ3nAaTtXqidETy4eqPr3Uox9I7VMsHV
3jAKGBQrlOG4Rj1sYkWDMvKuHimtv4+O+BIGvOj74E35NcmAf1qYK0UB48LmGx/8
j1cdfdxjdoOpzXMD+2otXzGN0jMxmkB8SNnwFkkWmlGbr2jx6gZLwZZ4Ua9dQfEE
u4cfgQPDSii2SMlBkoGncARKDeHLacFN54J2eVWV5WdX9sqX9IdswlxCW+3WxESu
i2koplFAYrl2sCwSI8FYEsOFI7gyinQ6WHgOctJqDUomvpRU5AvyILHhupb+Op+k
nprd2uLtr2vBIyZaookjayn8njhw32+zk7KbtZs9vSjt7U5gkCOdaWXQrLLKqNzQ
pC/Sgq7XlBDPGXGILDb4pS2haIAnYVXESzMfjwzY8TKbYvb0Dd/Tjs0V5QWruvb0
OvuYUZIvlZkiZtjx5IyXY1We66oegx6Xar96fbDTQBWgT4oulZAUowLfBdWgYnAn
42/qIliCXbUhmRUPpkKuqR3RKwY5w2E8jwQIoVQESTJQNXlYl1p4E244/cufVzam
Rs5cIWs/kB164yn57Bi72oWmjvI8W472+6wV04mcfACsNQmLOLG7b0nV9iA8jAOR
4jTL0E7ckOx1zqVetPUGjJLWS2dATZ0QC9+a+Hz7Rdhl18RYOtt1z88xxPf02T5f
U1E3Uu3VR3M9dUA/T2opvWKE2WYfjSj21IOVxzDZh19JBkzyhgqIsoWIyGP8Cgq7
7IHM1rhNn9mnOTyNT7ijn+fH1ifP8aD7bGk3xDW7S/zMAg5iHMqv1+3nWvmgVIaN
fRibnPV3frGiWU1FJozxoVlLmRgUOxt2wDJI7f92GGwPDl4yrMVXB5FFtewessPx
tqhYepUQRGLeLQqzjYAwYyAF9eH82VpprmQpIlZmA465Gq+02bvzcnCuxgmveNGp
0pIBOnCBrPPJY+gSRSZMAj8K5hEHfXqUuaCwZbLc1YFvf+bORR2J8W46Ei/oPDJ7
GGBZ9P2Bc9xZv+xjBbHWc61NLtDs2XClYh+Dw/l40EUeZVXp76hDBahAHVp9eWET
nLRrMdAiBNoCAMvfRt9ZE92kljJBeP4y015GeNDqfkhvAi38kng8xS7twZJ/e7zA
10a3GtiRyQ/men1okQGXkd/ka/PSb+OwrO3U/rk+6h2KM22t7bzmI7QzEluVTgJg
`protect END_PROTECTED
