`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qf/2wm8Wz1ugp4f6nzlcjp1KNl+L1WpuMP/eiFRaKt4GaEfVCdKoClBRKvM1kiAP
yZG+Il6q3orxaSwQmgGd9Oux3aDWO/BAQ8fsy9k5U2mhXqrsZGIBMAe15r+bOjSh
4PmE0XYuRX8keaYDLBrd1rDHdNYAtt4c3rqnuSi454fTWU3wpIoES5x7/ILSGGI7
VtcWmU2O3tpordQuoIeehQSKBXQyyOzVRH6E8jl/EL2tmEbftaO90ZcDkuIkymB5
0KXeHeUHFIe2OlIs54qSw5QsOvbTAk/b8Z39NHrdkx0R4OBcBHNeBYDx2E6qZLwQ
W3ym1rTbtmXk23U5ztrpN658rmkI7g6/kkgaRGZYJmibQ2b+KgY/yzMj+eoV9piX
leiGwClDd/gOrjA+qdljqGyhA5BZLBvBec2F9HbtsDEG8MdHDgNhz1CxWxRmt9Pf
raNR/FeDf5tQlAdLQVOdQmeFJnr1S3xIxhWuUFWRG30eFGIQokRwTW2i5tmwjc3W
DYHWian5iE04Hvl3CSwsMw+KZZ70O/BwfcczpU6H4OqUjfiJBWiP9pTHv/Uh17Qd
UX9jQ1w5oabuURKfZTopgAoUZVnpK9KHBFb1NQyaPrzAEE5RiQbzdFPLuES/mhIU
D3BO3THPgZvT5Kpe1ypxX0BqpugWb2huDtnVTPRCXIZI9zS5ZCgIgnCcqDVSgq5a
5Nbv8hiWtGAkiip1qEMkVCv6bp+qPvzYeF01xoFNQ1E0/A6ELGC86qOTNYxjhrqm
2N8Rlsll/UUbgn1KN6hiLGwvsowIlfc4Fatzqh8TPssiFNBJkec9HNxLyTxu53Ih
7mt2onME8wlqoslkJIElYEYiuyMvVpuqVwgx3RhQxYdRlFV7qQ+DSwgVlvI5QAS3
Qafu+kUXahks8jLV0xwz0nA2g+ZW5NH7aTiTOfDAKAZ9vtq0mIvzxvbIcAweN5kc
xd4QNIhVZeQWJhhqoKzbxcXuQUldMBvOZJqcbCqK2yc+Ep6wOzOx5Ik+/keeCKq0
9cUGC8o+ik1n1u9Qats+HQh+xfhJHfwa2PyyFJsf5JFBrWXvlObEl52Emcz/GxeM
9ZHMQt0lA4vqkh7TOST4INmuJGjXA3LcfjRdSQ6+1VLC/iZbYeQUdhx3EOHI6AGx
wt/8SThi5eSN6KpCSm8QmQ2v/VY/TuQ5Ur24eadZfja5XN12DZk1uU1a9bJyxUX9
Yv8gnYGsGgJnWasTGT3VxwEF+fgWDzUCxVoK48v2ZyGOGOQvbJD4UMhcw1+D2wf8
aY6p2yuVAtkYknLV/Jz0LFWmIzx4Tha1oG9pXVCYFhuiWm+js3ZMTmSgvQAjAtAt
t3W4J5n9VWX1Xt8+T3tgf9yjaQdN7qyd3tEG7CN8KD+3I8PdaQKLT6p1SIGAwARw
EgwRls26zzTIbgDtVA1XLL4HOwd2m0+NzKUo61COzC9R7FEu6aIbYpEnw9sFooV1
TbwIc3Bs9oyWg3E48L5oBtYpQUwepbhFoMXC6eDACMJLr9xC9vJ6Y+GtHHgnOXJU
cdU643YtUC9xV4GjlppD2sL6tgWXcsXmEN/4jbElGi+8KD5iu/vdpXwHbSHM2BYf
R52rkupVPQI45Co6cpcc/6s5SmsdCbj7ZlDDLACBe7yV512hEq6ENqCoYIFd2FRt
PS2K+SGATm0wJf1gl474ZQS7TwhOxwT41UtouyqyWPhsPKvXThoziXMbbjMNM/fo
JeOHwdozEs8qS5lfnIX4i7cWIFHE3mde5gW2vGbOrK1eoyAjRDROMGy62SCxkFQD
UIG1tbODLn6KGLjOsofggOFrl6rfLb11PM3zdnMmRL30rSk0XtkFXPywiKSVMxbF
o8xPvCocPSqt4y8i1misQFZS7NSqDGnzvrEzqDMHoOk73jYne2Gt2rjCP1A0iOtR
wCM6G3fawFtSHHJ0AdzQGj6A+tbynfrTmQ9ioXBR7yLimn6UQwNcjn73PWa0J3XE
w1SuaOvhqfcYodHQ5CkMzzoyKottWJvaAWRttvDNslWLCsCL3XWbYjV14YS8GUrp
Rf39Kg2L5TcLFFVyKwHS2qymIRYsk1fF308vnt9NOiVDQwK8FL01j1V0xV/4jcWQ
hk8hb4HkAiv77B4pm3CFWZahBNGDqC05/Oz9s5KoyGrgEY6mzlaCX/+2r7xjPr7W
Ts3qxu0maUJq8owHcsxgtAqT0VnfijKTrcCocyFy1GjCrBe4TzspCUtILb3mye1F
IwFpb8AYwUmkfvpMp7A2b739kgZmpc0YEy06l8P8skkPFjxmKWUq6LuMVAw1Gf6G
xpY390WG1rLsFbQhk4iGeWMg87dnn2D3437W+hI/rYenP78jthvA6vOQXOlZqdK7
JAo+9LRscj/jmqWTGWXHJHDQIFKRsQt9P/56V7GcekhHC1zuUomxON69iuDi9sSL
61YNyiGVLQhpedEUijswCIGAtrV4kvWFyTK8jpHrHyedo9BRRkNcOyGTiYAuhqoy
DhhVhahIfTBUos3ZcCc9JqfQ5vROJTvTAzv6S/aEd6SSEa6U0OZ2zbeMdvy+q3eG
AE7ytLL4JqQ/Lpv/JJVjnJl9Jg9w9fUxVfr2MbN85T0OeFGbHDJSwSeZSpE25rzU
RnSoOUy36mlrC8hwGyAQwRB5mYZljaTklEC4iLd72sYbJZeQoGRq6+zZcw4ojUv+
I/4jOGgVzNN3yE0T42CqpfJ1UnP9WqYRzR62Dz9U4yY=
`protect END_PROTECTED
