`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IU6UYvN935HTR0wV/iGyD1p3ddAQng5zzvJi5N2SUvFPtm4DYy3LpSv7Uh1U3TKn
9iLBj3wk7nvEJNc1D+zhN834CArmkwJ3jvfwV3M85/qvkY2Fibm71SqnLEto87Bb
AS0ypFneKDWLD2voCljcv2lvIxI9t6z2bIg7vd2ETlL7jam55pmjcqTDioPT1kx4
GebC/uRPiRSQ4caezooRY7DUMKm8bJeWr3AZTdqp/ioLPCD0HMUPQC6Bare5RGxS
Ojgvtw1cTyyYUIO5akCDxZiKC2beNBe0fFS2u3/GzcZ7Zznr+YpLP8FNkBTEXTOO
K0RyNI4j4NVhIuds873Guk119lf97QcZawBZBI15LjNDM3umD2r/9QnxpbFxiLth
qdC338LZMUjeNu5TLSg1cWlxUkeSuc/SsQTaCwkFwZuHyDu8tE+944vWDri+ozSp
L2A1hQXwUW2EU6cZ+1FxsqWo6NdiLWPeA5AOds8mKHlE5t3Ej3lcym6osmrNoRRG
YIBGHUjo97BRGq2oejkR3Kz4/ZvONA9d12wOSQIMc2Hvucdp8Pr2ofVPCYTAScFW
uQxl8h81PoGxfCSxvhUSkAzq0qe9IxB5167krN3qdY1n78QeJjtG95WTqo+Sfzb9
OiKZrSVd+j76jm+V+m/K/5QlcFJIiFvxUDQjMw1USm4Q0g/XltAtkGYH/EReZN23
`protect END_PROTECTED
