`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qjcr8jvBy+gtMOixHgY7unHBA3PbVRjUAC6w8AEEI1nsjk6XScIrB6twLLxfVyWb
tSrrRzJznCglHktmczoW6Dh1YLbUW16dz2MTf0wFHeOCpkg28FFOSCtUsWI18IAq
h3nmuWsP0a/aTCpFsS+Wj1PJIhcWLlp5fMH0CFrPZBnCAHPArxrymfeyoMcCCf5R
aMxpb6Ze6/L2kOMWpNVThl0X9405EMYvfcHLL5hTRikxu2V2CwjzvN6c4bvyoIAq
GalfOBguagpKsR+Cv+ZXK2kgqPw87H5ZScj3TkNZwtzXP59cs8cUvvg6GL5hBsjw
gFDaiCSiwJuzdtia9iXcltSlt9q5cbEG5rBtcOK4LkJcD2LDo/S6Fpm/m2wk+ZgW
4bEGVratknbapSJFMc8tufeiHvgL3DsC+/tcqYNcp//MxYDfP2gJKkupTsR2FZ3L
NMfJZeoSMCBsdfsRnZhUdEDaUzQRYVDkK9xsGVGdEHAzYGsW8vlSWTRC4toBesQT
71+Zhi9nNz1qxlY31jnfaU1Dh7pgKwRWOS9cW7qTXhZnmk1GWe0nbBxo7YCqFJfZ
koQMHkK+wjg8ZubN2K6mmNtUC56Zsef7rB3idgVCQVccLpDDbv+U1DmSeeomsniO
Y5sEcaPX+D+cY4ySGdc6Nf74hTEv7Sn2xMyoQxXdTJT+qkU2Mne2OQ4NVQUconYk
UAGhJqHbVnZaukbFQ2ZoYTPQtMGXdT6w2txSgcGWbgTeuQPKJnbWY618mrrt3Xew
zaU4aQrId0LBPHEWqNPg2Ytp3PWs6JyaIBiafZvE91zbDM8wZcZvE8+XwG8y4Jay
rtW6tSNcRuj7n1r89EBZ6AUDRrPgi6zLBsn0akXjUtdQniUycV4NUJfwBACUiIRe
SDcJHCay69HpNSNYMfu7Bq4aMexBKiohqXuc4tYLXONAleV1FzftyUVBV0cd3kd5
zUjQLkE9nxOfOvRq/8lHP72ufaaNJ0o6tCB6SPwRxTs/UCk6Ify4KfMe21UHXA5H
5y7u9TLYaCJr9ULLnOUxNg==
`protect END_PROTECTED
