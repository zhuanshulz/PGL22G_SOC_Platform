`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bXuyMpTmpmoPsrUN4eKNZ0I+1zuh6WfeJtIY4CXN457LHm31I4NHeWJzJb+gqYUt
dc0QmmjlycLd9TcZ4IsVNNCyBATuyfhPiQ2N3BgHxCWjBqzjx+BenGy+cKz/YKcq
nwSpK8Ts2Ll6RCrP5GpWQ68hqzn7Cnbk/Oysskzll5rAGLPaPX1Egn940qwMS/0n
7n9tmdaSa/FYJ7jXFneTygP19RqvUIJefFy4bZSn/oOa4jDPx4PAehYpB1tdCeSP
hcOASZpY0aRYxU/VbS+9gFDRyRucoKfaSAUr6Zwe6ll3sZyGTP+/PgR1Oe4YKDni
+2D+1HDKt85TTxWX4sT4RK3bxBAhIfCtWbSarYEyAxFObp+TAUotaXMOrCit2L19
2advJgq2d7MyHValR/WYPLZrkZf1Nxj1JXhir2L6W9z9JTCMOKJgWoDgqG0O/BxY
IdTU+yhIMrEYH3sqAtucDC28un+4Zv0hR1aw4LS+Fr2I7hXaucAEmluXDU2AD6co
YZQiMbetx83I4o3T8FVf8SpPfBsrTnYd7lV3R2qDarH5ObG1FM3OsuNldzF2hsCV
tQEYKHu/uQmv+XTJCzPHS5BcmYuVlrEnWGcsi6lXzy39rwNGbYvHhtr97nNmeVeh
iuT6OfkCnrQ3f9dH/2RiNQOv7LNS+12xAMmAc34QiTYWYeEDiImG7oxnzEt7FjVg
ELeg9uNe2Xu2pqlpj2X6rkJPXPAzJvWGEexq6qq2xNZr2UpvJ1anim6DE51uC7Cd
k76aVA9cYqxDA2lIq9nu4+302VkVu+zMNd9qCgIMTglJMrkUJanF264qtrGH3KMr
Piha9r49jRVyL4AYuH5DgFTjzQLg/n9Ilc4oVVzRVgICyHLQ8qCcRfaYdQLGIVab
YuNbnNIj026XcVmVc6ynSZgmxLhzUx4M8UDfjhh+CHZjulyY+k93j4Q/vJQ1EhKr
x0Z8XtkgC77HrFffqeVBR7DUXjBTOYAtDgdtqCAmzc0R3iTzpm2fpJWeUC81ucN8
uc82szCFc1WWBpGpk9d5Ww4c0T4d/z9xkBxj79rizoHpD3lJI8MD8a2knK/4dCEa
AcOM7aNYa5W1w539K/x8iENy/ayOqj+fruDN/sYciKj10xN75fAr4PJn9STZy3aU
yCdZxLe6YsmuoaAUSK5+cniH/mqWXuJia9//5w8rALcn2U9+y/6QEBWh9pjJHk/H
rPFk7Q6+3cYCbgzXuBmHIkDQGZjYI8f/hKoRdZ4xewhKO6rnVyNRnuYn+ZakSfBx
k8CtooXboZKOprO9IbTS4ls/PHGFn75Bsn1Ki0oZiyWZgrztPIYR3dpougQIA/7t
eUoJL60JSBdbohtU37kxlk+ExhUNJJAGVIbd2vdrAYbp2Co+PxO352k5ZjMuEiUn
IHgcJE+GpDOKGAr7G3D1Cl3GdlQo0LxY+DG9iymEqY4Y2mQ03VLNk7mkX+jk8f2D
D6cYFJRuMBFiOtQXAL1leIH2b2hIukBdIj72IkRsMqQkhYQaY9x4P3wpV8Cg/3qA
QGAwhuM6o+C3suU1SR0zSZdvpbQqdfxgJ1Yz1yugQ0WoH3IVwVP7EvZ/9Y6glL4q
HqwZterMMD4FBlPnhOd732pYligY7Op0Ifw31jnucQX8iZnrMRhq0s/usVh7GzwC
X48tdefxvNhEI7A1Y+cLeDcHMOCHThMtVX2DPqF1U8CMFLmWGVhwUBu2y6slTRLt
daDPGMrEbgv/+JsPrKn7I6Yq7wOenLYHmb3YArhoQuUCO61Jgr6Lc3XuqhuLDgmv
8+/bs4Zo6WXI6iq6XkceTOQTqxAi2nMMDoPpXhRmdqofRLBDQdgtcjhTvvR50Ur+
/sFrGuirns4znY91K0lT1R23AQIfjDyvICT12lGK3rNiLKP4ZtSafBPyPikh6QUt
e69viOiE55otSwTrY/Z1dRX5DukQr0r4aks4bBjSA7rMumzEVMsW6ukoc6CLM1rm
xzfa5QKdlXWC1ISK7iJlyCYybWQRX3NtnukIkSBcABApLIraYizmI34SREoNyowN
JeyvSl6NqtV+k6XiFsd6xeqhfpCllAG6Fe64K5lKDzhxTzk0tUqE51x/rvbQORSg
qEF/WeCck2Lqr0P9NFDV/AQKmJwY56RLPo5BDXeKLLJeMrRBAV6SYeWIP5AlM2Aw
h1dOJof0LDn/CJAp2XVyzVIGXdun3wvFmW2+/6O85fTtdTW/R2dnM9dNcSvpHOoF
A3OkozO52roMBnJIChaTMGlxhh50BKwFIuOUhC/dUG1j+VdVGmhct0xtmGwyVPUC
jWyTdi+Y1iWyBGxeKjT+DxLsiUZ06hB8vGyD7Xc89Ub+hJKS/Z3o8Pfm1vXQLnz8
qsGe+RTQ2vGItsPVKjDPjJ3mH9ueEv38yA6B4s1alR/EqUvhcNLIbOvGfG0RqXvN
Svtlxygg2ngqiN8XEBJOrJjMAYkOBMMOw94Ff6zFZVKditKK2jCVFvGSaWXVXvoh
repeUHXn2/AGuJQnnPpJjtf3DeYtFsxz3PtH6NLnJvYUBrk0jExDz6gTcNjDW4fZ
NA8pd4Eh9VAodBjnTcEUiGgcFdd353pThhzZZyDmQgWEHT9uQtkq7E6mr9umJvlw
/KsOJQ3+LOFR7vgk6Hr2TvFzhH6K7CPucgJiHTqjOwy4+ZSzxVOuM6+/LqV2AE/J
JrRjUiPnB8MmZodGfKJk39yjaV5fQCaB6bDU0UraajGzvTOCltitBrjL3B4dPa6x
ZHSu9UtMYQIG3A01EXKLMNdp6HQkaZB60AclrUoFqtWgvJepv7jsUE5KfiNApeAe
IGH7TzcjCUQjV6QxplpKzAmVPjV65mPzS9CVPmQGdACkr9WCtBUIVSKeU4+Q9/OC
D2KMydQ65xI3aIQBk2TynbZJ09ZtjINoVjiUFdVQ52l8iLHxK/SgMQGXCUkhNJ/3
8cjpMhFS+XH0L9Lyb0VPB0vuixLTx3nQUUWXbOhCrXexavdzgAIZToNTSbL7Cv4g
Yw74WmeMEd7YaKBQWn+7j2QmYfljs/q0KHN4BdTAJJMrjJ8zHxuF0sX2fbIOF1RZ
nLK11S1DcUBtPfZ0dTzg31PnJQuUhKcJvhsk7AROWI/8vadZwSKKOyyn/3FY6+0y
gsMpfnvY+MqPFmbJvbW1I53ejkvk7DpnWCgTxFnUg24dB7oBtMsH3XXovm30GuRN
2LHWJdtm5lfyGHa3BMac/npKR4vM8Mz6HJh4XkqiHrHvbAlLS4F5boUJK2EOejsB
v73slJgMxu5gLPrnacln6DF0JS/RIxlhEWbptMbuuXp4jYbnae4/5QfZwFREmAE8
jp8xxxxHdAHZjyjkeG00AovsqU7CH6ZVbavewNV2C5b1tI7RdDU72rqEptYViTMA
RE3gTw8I3kvU7LF3Qvv3Ni9KhohbMaFXVj1T3ykybmruPeHrluN0kCj0vFMdP3e0
ACwtL2x4lj8T4hfgggRkSk9nasD6CsuEwrqcly4UyKt+zjJOzTBSI/2CeunP4mBJ
Nj8qdj1JfZfXsT+7Lv6W1UGkitiYUr3z8rtMkT5TdHQT4Zu8GbXqejB1MKawDo89
ntKqIla8/lCz35lbR+xVXcrZhgetnVkZnzHnDgar/iFydttSytR5c8580cXXI6MC
it7PhPF4un7d2skEKo5BNKnb3cvo79hwDBTf+mcAv17CUOS1rxvL3+Qgx0i9tML3
GHcQi4RJfQv2zo4qO/bvrdrs+wnqK/o9y1ku1HhLTfolR7w8DI76r8rSufAqH6/0
evID6nj/WUoN9LfhA20wIi4KqyXykNs3huUZTT4Vyj2llGhNIj3IlAJDOP/vw3tP
OyQqqby3NqQkT6ovfNYJ2HJxzQ6gbUS9LXYGdKdVpb3eNhMDDdi5z1zmfZs5tMDd
b0zoqGZeVG8aPEof4ScdA437RRlWv1xs19iM/5nz/kZ/o1uZJjFGvDdAJAEuwmfk
`protect END_PROTECTED
