`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fOsR5pjWrefyHV6a0ExveGYBrXWegKxDP868e8+wOkaeP7a9TRentnu3s8D72mPb
OHEwBH6VKascUKiiiUrSFT+J7N9EBO/F6BOaEaYEzOBptPp9lNmd2hAERBe+ci79
MTUOY39z8q/4/pRC60wWyuQocry+2LjsP866d3aHh9SfXJZuMKSydwUM+jZn5XE7
K8mPxHtm+h3fD27lEmHFWMrExgwkcSd1WIlejsQyPA9V9s/CtF2mK3qR6LzBnImJ
hToFY88XPNJPKJ+8kkXgc8i96PZeA05gzIkvGXovpN1Bosg4Di/2io3q6yuzcFkN
`protect END_PROTECTED
