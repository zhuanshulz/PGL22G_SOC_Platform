`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D7X7xhUoam0VhmIb+pz0cBgTY1BOXSWV3sDldWfST71NcHK3xF/KY8O0w8gCf301
lJZg2Ax4W8sfAyCTXHcKFOoSeDQCWvyunF5PKY10s4xfzbZQjLPhMOIbUXikmpk8
ckHvncWbkLDIYLI3NrK9UXZoQWgyGcIxrY9hGzmKyrvhkqCZOflPT+iMwDHS5WVH
NKa/akJUvFrE0gKxTC7CSME3KMrTlAYS1QRjn6q2CYpa5d34QnCybaJ8IF1FqHGA
ONU9LOfNVsQ+p8ItBMunm7T1JZkLtkopr1QfIwW5CJwGav/6mrtapfnyoHvI6JJ8
8e8ITEvXpiaaXekqvjc4T64WzfnW4Q44lkuxMkom+TDT7k/kbQ7FaUi9pwBQ7SaL
9UTl76AntMkErQ/zZXly+IDzT+2CGL9fThgNuRxenQ8j0sZjPdbGI3997GPgW+3C
gCbDym4ggAGvUmhFkftS7xP5hXCFY2AFaj+/DMz28LYACVBc8mB0RQHEDQL6GFqn
C5MxZggY4TSzZjeb5YtPAwka/QlRG2BQPwPPz5+KKyhaCt0HMmtgt9GwDvlEwJ+n
Xu47g+7rrfDiLVicHx5S3nAHyjEuqQlAfKmhkkDCdQVdNPIr+PeIXFPqumnqJHeR
IeeguYVX/hKZPggoi/PC46jKDrOkcDk6ghDgehGQLwdOESrjcYhW7zovFgVS+YK+
Dxbv0FrqJNz32RljaYXanZ1405l0hb+Tty2M1voNPOTwRrlzbKWaPHwOp8lNLL3d
4xy40suwvqW1X0bTo/pd5/9XUNYhIQfTBR2hUmtLhwywGsHZ5keT2IGTjHW5J07W
lsRKsRDq8rCWu6xFNsyT6PYhD2cj6zKshdTeHxxo16aRk5vbt2PGwduDO15R0780
+lse8EConwN7BfN2zcro+T77DrhbsiQO9wQ70pLAmwB3XoR/iwN9YuEgNCpcxjbd
29/coevcdPhrh+yXBAIVRHsLxWJ2bMRluhWfOL0D97nz2n0JyDmnpNdnM2aTEEuz
OoMVnAimqPFIxXynuHU0/J5Hza5FAsMkmoSq+tg4FNTvl51hDfQJWv1JD1fsn4Q9
dvAfK+pHF4J+27w11J+yUJMBoRCn5GZ6Mu9IfrgWjlRj8M9T9jsl9chwoD4I8Xi9
d9S3mWMsW4PWsl4OvsR3yjvEaopxv6yzVkIQGnnYHOamubfEyuCt6jnlzhr7q562
z37nyB0T44MJhNZjrs+qXfd77Mt3DJI4zTGtMyf3WwQ3ZxaTxQdVjJugpqVAd66A
ewcs2A3Cipm2eQa9EPlARRLIOE29rv+d05gyW4R906FQZwxrfcfCvppN/ZQzSvZE
dSVn2Ls8SR5m7epx1UrnsIZfMxpjOXZa4CNHNa8+uNRzbE1I0DHWx2ADzFCSwXx5
52Kuq3w2b5E5O/RERDFj4E7HDt79NCsPex6ESfPCr9DUtVOk4HoR8zZ/QP8KvZ5I
/BRJsIeCgfVAWPhHNTQPGQvkwHK1sE+K6qIj6oN2kaVNoFwb1hq+Gskd9B0thxmc
s2FR5hY4G/5SyXGyqDL959p6Nic6XuNDFHc42g1FR1RFsx7yJIh9pSs4Hj+NkvGO
nPBtXY74RPyJWgTFtB3UlC3AMqdmtx8cGEjKq34GY1pXLqgKkINVHv3QDTfe6/Gl
KsLLCqsvlhAA87yjd+tD8KvXmrsIQBQkiunS2xIxJuRx6dPaV9wGN9CsYrJHd+bb
lnkryXn5BeWI9nh+upU0umJHJDlCTMsJ2fObxBuMexBhx+FHs3qIwNgPOuDZc7tO
HDQi1SDo4V34r1w0xs8tU40SCNVSGcwUh53N7f007ZZAu2hlvGlV2LUy7IgO3TPh
ob1DqnA/emY72Cr4Xd1n/Ujon8hSzI7GtpMRyYviHUO82zs0BsfuesJrFJh6S1by
nWCAtYNBvr330MIjumJ6XRg68nyKjNQY9aQsO3i1xTQo1tmhrxTrf+do1yGYpBJZ
XxTp+hBPaEZkiJBvxOZFue5tZgwnU35DBm03JyEtNvkM9xo0TbeWwGGrgnZAgajR
Byj+0FOs/LylhlDhaKTVoZUe3yqZS6zWf2jTNUClp95PWb1yo+0r44HP6EqOc7Jx
3mdvB+EeTtj0bKpRasNorYm2mN3NSGg8wGPW8Ngpb7hJI1hgHHugsdhCSelZ8Swg
IeZcAyvflvZ6W2u504VeoQjme/Idj6q/n95dCVk7w9d7tTPBlB63EY0xbYMpb9t0
fMY3ba1fimYeUSs13eUPpw3mKODNWARoonJmunpblwW2hEISre5DZWqBemKiPKKe
N2Xjij+MOrnnuoiHhPoGRxPfpI5eFI8KAtOY8fP7qBl7RBg9E7sgF1Kr2ZifRkQe
ElwO7y9fbapCp8zlaYL5QwW/2a/Sthsf/MznFWDrUYMJMJ+Jm+q8a42NquGqWoMt
PCas3vxdCudry+0XjhMYE3bTwYo4syjbxWYrYhN+bEBcPugoiXuzmAjwar01N5k0
7IxnVhdJHjSzbxfmIqi/MHd5dbwXyX0k4g6VtO0cLBdzyIkq2iZprIvbgeW6KBS8
0GfiPIGbDCMNCnWFyCwZuIPIRb7ghm7hUg6JMGqPGd0zhy/CTwxqqOIhQml7mujA
kFRak7ZnP2KN4YmZr5Na6JEl9BxmtAth7Pdl2bG6JP+6DtPJrFrqvPXCZ6vuVytC
PVhA8wPgodUwaI7kEtSTThz96o1fOS8e/4m48O48mpQoxlfDZidEw6zipPuGw0qa
nsWP4hsH2uy4Mo3lGzYBtE6NgygNgSD3VU105Ow7OZl3vzOF23gFEIrhYd141Tao
evRWWNPUVTdQxLjz5efztknYMoJkZuUorMsUltuEkqwADNJcxOtYskZXyAbOlf3Z
eg8jPLIEKKXXBTslp07IWYpbwb9jSByQP6Dh6UiMT4jn0hI29u4C+PRTtGQAzg2/
njHIYiCkdK5gzkGc69X/1GLKArr9FdEilc+1TvcW9z6wxqPqCEqBE7U35Qua5+Rk
8FdLrdyUn04U/dJaF+8YRbK4zuaXmSHPxnDgVwlu3BIrWKL02dyDuZMbjcidcGNL
qb5KNUzDZxn/k0F9xzI/xnQhtz9HFNDM7t2RxBYUc4iQutD2tLooAJTrSFDpfTqf
HKVXdmmJ4lkm2WI/w3bcH0sBjsZpg3kdhldqnThmmpeKj7F/3kHJAsQhYP08m+YW
EqkKhn7VB472fg36kAXXwduJmHSDokQ2ts0W8+s4NCBTtPko4MGJdTS+5f7Ow0u+
S0z5SvKV/nV2UbKsdnn26SK6b6YUVvMDH7kP1PKu9up/F28rUCD7c/c/mowDPrYz
90NuAN2P95t7iMZLVaJAA3jjeLUwbxT8+OgQt4Qj9Jt2OM8f5N/7nvAzJgOvdlKk
KSbJYl9NNeoJeM8IJJS3A3DL+Jo6xQoF98z5yQveGg5v3ITR4Ak0qSkW1xydthYy
KcJUNClqPNtQMULa1u1LhpmXCT/LaLv7HFxNkfpztIZu4lpRQV3vgLIcRqy/Cy0H
8bYlwbPpwa3PCjRBG36QK3zLNNSIrrnVbTvCAqZ3q0CA+EA9yGmIA4H2RGdsnJSp
FTKPc9U2A7OBE72En1lxLbWTsmQNpcQJQFi2L2Th/iROG8YVykm2OhD7+t8b/Ssj
8l74UfZAETaryNG0IqZJAY+5jvYRqJf0TxbYsDLrCpIZREfqdcf7qtWwLvW63AUY
Z0VVTBA+14LSIL2oElaJn4y/IXtd40IHAad4SIvRJTTH0hiIsjGv7eixEyb2OroZ
s/IuYpPDnlPFiAlp/4G5ytk+dCrH0blrv2j2x6+23Wi1uNDWJvG0IlPQueHGiLK5
pQWec64qQQ0NvvTf62eLO9oS4cTLhT5H7nvYp7UkthH45JAiyjhZIwsVhIadk27O
yk+cYjWaqUVZpEiQpaOiguAYNL4tHGLwUOtJaCEKljTzegOcbhcN1BEM9qedHwvv
7znxU9p0G/XZMc62x/2GDr7tM94KnilLcEMk7qWOQKYvYecUE7RAC5tqFWGmFhAP
YZtAhEfSMifVlF+fLUAfXDgta9jUOP/h6Ymv0y1x3R2f6gqXPdF1qwzpKZ5aytIH
8C/h414i0imACSGpE0aN/Wxx+uiyGMIbg8G0AlyP/GI1GoJrv6d0byyl9lfmNVkO
mrK9J0taQd1b3D6Tc4ls+S5SkPCBA7NJlZUPNnx0buxyf0hwZ03jgPcjeItOS7sh
K4fXPmYk1xByIKKvSHzdNyxoO981jIG6eFU+gIt84WArKsLohrV26LcwOSmhlawH
cKeudS0r9BYa7FW9Sj4X/DLG+LYcyUC/qZcZHctCzyMqLJEFPftqlyrF8EYgktL7
DLBx/CnAs4QkRK2gCx7mWEvcXDuSQ9l9WHuZE14gi6mpy4nOMg76Xd0wzeskbtNO
cI122htnk+VG3gLfetJ7gD1a5PwjI9AuppiNTjVIQdH7rTOXmiMTyhQIDKjk7C9u
+G9XsGeertC0SNOp9Fh1pK8d38+FblA0CBwFWZ8LPuDS1YYyQEI0SeHS7jnDj06M
nmWLKvFPS/cqOfkZkosMI7+zzbRAlmZLrBnRiIxAIN/26ElBRalqbLj7O4hq0ESu
ShTsGo3j/bTcfx7rh6B8P1Nbz+DN3U58SluS5xvM2ienngcEvIOo9KJKw1GLcxSD
3c7IoKKZlIAhb35RN+uXYoK+Oae7M/+tEnIJp1QHAfj2W+ZXa2xxJ/IckX1p5csh
mXXD/JAOtZHPqqLaak+8kqNp8pVQnllhAOsclCflLQKOQ6KDF2ujMs7icf5ftSrZ
ucabRqMdMd8zl2D/AflCOoc7KYxusNnf1biAcCcb8XQKEdqf6Q1oL7upaY7ISyUe
D0nOQHJpxMPA34gFlepSyALjOXFuE8QU+kdMfhbo7JCsIvO396O0a5PAilvLZ2ve
JyVQ51IXCVtWqNZUmqhA+Q9g+rZdEbl73ibqK6i//z+cVxum+9pKkaELnH3wCI9S
lVtg8NPBvGkiTYSjD/7eoYLlj2D5hnXnAO7NKUO8RDs=
`protect END_PROTECTED
