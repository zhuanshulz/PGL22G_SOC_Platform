`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u5mXOuXbtK7tYmoZwLITjNZ2Br/S0qyC7Yiz75vrwcbbOm69bf63rL1lxFegLL4t
V0jeFW8SxjUcUR8nh8gvGeUZNSqZ0Ecr5iG4wkaeihds8InVuUwSfVxfKyB+1I7s
p1XMow/zswmzHvpvrFXaGpe1duOC+6f9BDXbU6GQo4Pxz23UtGUICebrrYnVan6L
w9sjxgtJtZhvnjKWHh2rkDQpFFI7DZifJKvDGP1OMPv5YxAquu1Ip0KkR2ZnFRi5
0dsaACokDxFJLyiY3sNutMg6dj8eVpvlrnNytlgaopjiOzdmwewlepL5w1eb3BFC
2QUPEn0teSBUkUWhE41lEaPFsqDrqnEhwTFWDh9kILdqI0Qv5p8BBqYii0MQj8y3
39bi+XVjc+CMcyGnuA0A262MJ4oW3LVkd1h6ZI/VB3zN99tyfj0Kni8rzAe+jDuO
BL55LAQRF1zl9mLZTlPxDtAq5wxTKnUME3mKFTJT450=
`protect END_PROTECTED
