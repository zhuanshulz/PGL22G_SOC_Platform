`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x7JU0vC1XnJ/CZIwYWHHcZ2G5rllNcEAnPlPm97zQFobOlzxlosudK9+lLreYgv9
cM+CwKJD5g4nMgTHM0sYdGwbgcIvZlX1xi1DqGglWp9r60sSbyodZhqFzrGWYASJ
NWATbmSmBl+oa1VLafs4oLYYsO/asg7jYSNZE8n5oEhSNgdqz936ATZL04j7nPBC
eHobqSq3Hr/9oEUUMw/wxULzDNhqdefgNuIJtMGC6FneOpQQ6ZeOG5iSr2oeu54R
7T7c+bVn0Gpyy2IghAW8GAd14prjTPVJXfFyy8bedz+Z2xfONFH82R91p56WNzSx
D0TLPV9Gi49fgGcQSz+uRO7nliMG0Ani8km1GrBOCuDyEj1Trii0In5VF9lZVfgC
NQGRhInbztzhrAYPVDtk+KXbVVyldFss86H0fWtCLvTAG4Ff4bJjjdTodM1wqI4P
WvdbTEuB/jCCbSsH/lbqNMYyoeI9T3IXWdYS86tkvTp5bkKE5C1s9Z+UVYhThBpK
zuqk/9yhDpu+Gwzj2azLMVOnTQMtOzURRb5Kb/6u0HJ1ZbYAsKgH1y4i+Vwbg3PA
EiybM+DwJVO0yQSoGej+C28UKux4MRzpJz9mH4t/2kg=
`protect END_PROTECTED
