`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FuFmJLC7w5mD6JEF7YjXsidASDpimRSYS13M7dPImnjT9xwjw2e32wvjyDAR65PH
KZuyMJYp5NWIvxhXh8kvklqz9zo3DPMS94GQucCp3zS/ipPY00LlUJcuwAYtzpO1
UKxN5BTgRJagF2Y+Fj8+ELk1LFcsm41DEMozPENo9q8VRxAUQymVG39+34U8cqkJ
zzEJevLbyG8n1QYlCz0enMzjsg/4C4d3+Do6fdC+44Vk9awPhyIh8Zgo7mK8XRWM
IvxABFNzi+3npHwIAQEmWZ+l/9kFaMjgirNzaY6RX21JZ0TChyWCDLixMJaXgIGZ
5XsN8KMw/bm1Dl+JEXzONaHrpOkKYfuoQKLkm0njUa2k19J1CzstCxAaQ9dKwQ4J
tUwSqyTqbGXZB5kY3uMNk/2qO3tjp0E1tYg7owB5+Bq/frKDkh7bE91BLW+OSpHR
F3b2VpWBrN2d4tfAJoWlNwwXUXa5YJNd1kBs6DZvvPT+CT113d6mOz8PW+h8VO80
724Zmf4RFUFRgacIjcpDg/rtz4G6GQgC3Eot4mQPLdYKuMvnzzFYIqpiqaUcpAk/
f8B24l4a0sv1C5dL3Kq4KA==
`protect END_PROTECTED
