`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sGF/1aIEysiiKIOSQ05t7dtCrczqtZU+LQk3R3vRM7eBs2T+3WxNPjY+d/dX9ugQ
a5AWCxVCYHlI7EbQpVy6yWFQCjt8WBMlnWqZh4r2LKjlp+rIM4veqKkf2mLwb9fp
RxjInV0RTW545wJuJLE3VtxTAE6usCT1lUW6HJ4mhXTHnQKiHDLG52P+GJ4sor3n
de2CcN3C8I80IVPLn7qqbj2ejuvcdaxZ4sxLGxAPCPK5fMtrzXwUkq70PDBWWqxA
dlZjedjuyGa1LKisgGGeD146dKSokdYlVJ7Y9B8nkf1MU4p7cKCBRZu7PEGejoyh
DKaTonJebYVZFdChN8ud2ZhR+eYwbYBBxe6HfGNsNED1YI7D6cVZLoKS6uprCRdX
saTra5UTuRaybcomILZz1fp0AmRm0FCvssnkF74RoGHVhVO0WX5leY3/ODVRFrjB
o45ir7rJGl1mpjoVhriASXiwh+Re3ppHwoBAeWH30VDN9cQti5CntlhqMl+qsTXP
IT1H6YXLkPnPO7kjppKIhksF3l15kZarWU8yxZNS7wfqeV5nU0c2q6dQNArpiLa2
RDh5FkcUEOYO78qL5n9uoHlcyYGR8/QXJY24lJmqxd8KGr7XYumuwlJZ6ut9JoWi
hZOnIZiu9HtpzIYuj8CW8WBiK4Zm24+WJ6bOCfcgCHroebvPrqIjolP38yekty5h
iaOAAnzr1r7OnJMU1QDPA/XzQCic9EWEJ+CUQ649PXTAwXa62+vl87C0t6x0TPpH
YIjv2ITmv8jVXM3dt45a+dUBj4PT2x3wUkP5uXS5FbnC5vrATFiEPOH3+uyHTWNm
L8iVkUHmNly6C3Ui5XEcb4OuExsNFhe+aP/9OgVfbh0WzYykawHJlgrDmoYJ3vhk
wo/MkaUPfV92LaJ1uqMwbQ==
`protect END_PROTECTED
