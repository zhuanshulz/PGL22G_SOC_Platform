`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4ob4DIcPAEqrUzyoUvl4GSY2p1K3U67tktYNiuP37JNEvuPDskHn3uQosT3LNUvM
DDGgr2XfsjsU60Z8iTlrsImKFHQ+GB/xsCv05VAYZfnANj6MvIE6h/U6wJNiiV2C
7nf7Jm0DlwQYQbzNuxpTNC9R5W5kf9L8XJms4kuSluZXUmM+9bKTWq8N/gJx5nn4
VJmXbSyMU4Rj880pfHwGFV+Jx3+q0aCpR7A/H9mBzioLvfQItAUVTWemBsRyowIV
Ad0D7ixJJHFPmje3zLCVqdGZAfqipAgUuH5/4OMdTkbO2icq3JNYYLJGcjmBCSP5
h2Ec8Oz0QI7G4t6cl3AAr0OOtXfjhn86eZ0n1134xY36c8b80CESFrf99ObfCs6q
nTBvFB7h0Z5pN2Zwfrwyqf5Fy9gctYqQpqr51NCt+K8Nn2+dXUflUnLd0BWX7R6h
ToKExvVZww+Lk64xktVXZPenuZD2Is5mdGfUaRsGCBrKP0HPvEdRK0EnKTcS8mlU
GNiKew61vRCAznRfo+P9NQRqt9UDoEVWYUE/J5QpQAEwj51aRJK6MFHjicMidS1W
tN3q8WnkdFZf5kCgfZ7tRn/YoVqFKqbCxDSqi8C25cnqsFHpfbUvAOD8UN+3dm/z
e41ChbUc6jd0P7JJRzY10FvRn2L5GSaQ65kG/es54sIIINrl2dCWexU5dM+JR0Uj
l7YOn8WG0xGc5h0ZpEyvrvwNUNud01a5GO9MUrMORBJpXQOPrsPiY0anWvJfXrVh
`protect END_PROTECTED
