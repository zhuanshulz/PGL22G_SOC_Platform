`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5/66ggHZYSsc0bdIgo15Hx0JYBbD8U2X6MiG1p2AD0UurbIRTc1CxF+j+iHP7ay+
k0SK547A2SRb1PqN9Yrwd5Yo0OX2ABtSs8MMP7Mx38A6pJHs+DAjm4GvCw/f3loy
vtiqiHgM7LpZ4aDzW5jK9YmGQyLPPEQr6vRRWk0DHbhM0BeYAaUSoiUJaV8rK653
j5MtctZpO4dnVmHZOxRnmAv2T9ICzHCoPN615TTshP81ebO1iuMiAU3j7KAZv6/E
KBR7T7yHMS4yq05oGdD5bSl194dSGrs9ra7KIMZhVEuJPBH1wdZhbZOn8lkHW+mD
8yorefaZPCcTnsLDywB6M/QWdSfLq9P5FWSsRt7iVoD4gj6zrzQVV8iZQkDsBXNe
NdsFpCG/4DjdLcpVnUumsYzdBI6xob2tdz7JXZGxRhInqQsSPf4DzCQqZLQZphj0
VJ83lVLUakbJRUBXEDGVYduVQFYOURJe27/Kmh/06y8vRfychx3zBATu5UZ11hkj
hyL71NmKX6MGiRzUOvs4QT7zpQaqMMeMQkAFo1hAp+kMpbf+hIpPptOF3TmS0YNZ
9nxNMfrZJqbi4PpGUMZSlTds8aSuSjJYQW7Tt9qZeHYd4Lx3/8Nl1du9BNqMPdFo
qLoXcd8OYpen45WBbkER3vcHEeF/MLTkFEa5MKMfN5Bl6ucvTNI+RuP+3R/QeD/g
9uo3psc5ERVyT+WDOtPbFD3aK3JB3tYOj94tRVXVagKmZbrfdOnLWN0LtymtDCyY
dxlX1JjQH8LJ95b2B4Sw0LIm+J+JcVw6sjqQANvXk1UmhkpNw/6DK0NXAXsO1vie
tnVdyjOEz2lCfuxPJ0NX6QPoNEygUboSEmBP206PINbblpjAp0C3YP7DgKrIIftI
f7laOuhW+lFjbyFoK2DEqxuJ7NqAXzhTmzb9VXEf+f8OtRek08YQrDE9nnms3nkc
zxRRYu8gmzfs2xypb/MTyidwxMj1AQsLeC5qdtnKTuyTMtAAJSKfqzyavZtBO+n4
pd2lDisuzK19QL2vnux4I4hsFwUi0aOVRrupIaA2zIy87GW5knbqxhjgUmK2YFdC
zTx+UfFtC1q9eA/zP6BUeD8Ys0NSEcdkKyO9UDnSjSvOppdmbWsfBpx1dGy3XQnD
LncVvfKttd6qyW60wHYKUqiZpDda7UjlNpu2E76PbsgPq5GcpYrN+fsrYE9JdyLL
lQKXhvqyfSIzieC4lmqQUtmHNdDff6NfcUcYmHQV02GmUvjFglzYt3Eq9SLco9Gg
sADYz0sGwSEjJK4hSTJ52bQ5oRckgFATHmhVsgWfpml+BJVLFVR8uqWR3pvRsx65
dIFwBMH8CetEvdhlvgJ/17Wkfax314h0yOD3y/5eLQ/H6emjgZb/wD3nTpHWqRm0
0kC4pFYqCvSf4HgNTI04nXt/pR8ltUuDFRumPuOtMtTvHv7AK6ebUXPVro4YLIam
T5PmfFUTlYactFKeTffvqnsTz59d66oCZyEXNRxOKlAjndZJ0sO7r+uge4ggW1y7
+GRp4IIMi4qQJPb5szlYAMKeMEqpQGirbTesoOCFXmslDqyXLedWixpGK/ZBfCyl
NpAtUmTesc20uIsW+4jQAvbbYBbTF4MRuu06mZEHDO8rHERJ77yIYjRVEw6o2V5k
XlveSquZGIBR5jpPIQ8Ebj3+7Yit7Lb93hsgnqvW5rgLfn7ryP4zWEp/JtpaNlj1
NYiD/V9jVkysVz+BXjLUpxbm6AYT4Sru8mReC9j/hH/NlYaOFecfjbryaC4k+Tp2
ovEuc9yLnxO46hBWmRCVr41JrHFY2zAJ0+s3SIRKvm01vJj2eijT54EuXwpDOLmA
j5ZM6URkUXRkA7eRXAmnd8D2PSDgn2qsgbiyi+KNMQZEuB/aO3bWwzmOkawWs9jW
S1MjZhY/ilQ4SudARPDIUh/qfp23U5aq7PMiZAjCVmVt7L75pgNHaOJPq5e3kVcx
khAalTTNcTO7i6+qn9irFtX+RDlezhSOTSkdKDu4r0mVsj+eTJ8wb0wWCKwkoVnv
bvnS/9hq8sW3Kt03JPSLMfGv5Gj6EJ+F7Rg7cphBchAgmhTF/Pu+opJ3Pw+KvR88
jmoeMv9J/fULd2/ki9kFsQePGHVcjDMzY6jQ+ZW31Rc/EhOk6SWKVgmna3U3nBEW
/a+Q357YRNDE5dRYH99U28BO8lb5n1mrDI+vcyg8YDBnJE3vYLmN4qdcSkmSpsMr
+DAHC4s3hxkgEw3aeyOAXz4qXG2nMVN5rT4F8E/2o/gDJo8j0U8eT6sz2svWJI5L
P2VtyItUTk72UPoqacdo7fuv3WYTh8gpQ7nAnoZ9ewyM2LWB995/nrM7ug5glndX
bnZ2zp4ukZHvGQgnG4rlxEDPd8COBU9EzmiQS1kEzRBksn60mZXmxBz1/TYL3eCa
ws3+8lpv6jMMk2/jgCxJlDWEw5KtwkeW1cJvaGAdfcgo7pWRVsl65+dTmwmFhK6T
nLh5YKT2hq8Swrb4YP/HZFRsptjW0EnxtytCW/A4nsh/sp9uRl0pYuumdXvhdB5U
VeymQqwwDKv+qCeQLZaUO5gLh44HCtGNfzwWAXCLpMQOLD7uRg8OgmKCja6xM/Dr
GHSrRVqFfqNzIuC/rk3sVK6zQN3bFrqsEwvfHQkntCmaWxg2/IZ6ztLOPLWxYXl4
cTA9NZmEe0AjSq6T+afk5+rk9zgzEuNHtkA8k7uUY1UnfbqbWwbIREoXXRBdwYXS
lr2ZUuWPFJkg1maapi4MFeR/Ku9COFbbHli4eMnB2kxo1l/DNQ8zkcgMLfgi5/AW
3VClVjJMVuP1VDu37/2qAgXcFT3j768mGpypL7QXrYG844mE7lto23xUUkpUo8AD
b+pJWLBVFkPTZlb95ehIbLkM8qUrmkjEp4FPeq1uSxk7VqLyZuh3arEr7UALQKbq
0BH9gqNg2zvxCmXlEF7dUCY9NcVE7B3hUGSukim1rydFUyEgnACKnERnphHa2+8D
Np//rI+aBiIWql3DfobfRUFqPenos/BtVfzGYf7cKT2vx5uLmHOmZBbCK5XUkDr1
sd/A1rJJMvbYmlbP0hX30z4nNX+nYAnrDDz/a1a7SQB/PmaFh6tNhDhNPhK6v1Sy
yFzbNc1hl9Y7/e6I5XOt8918ICvi62+5IKyPPw0o6lhEd1aDhE78Y13yoHIBhb2u
Blq929tT6fdDmPvJLKpGK5eoBEjJwMTXbrlXklBG6KBkfhRhcghjsbI0p2gr/EHf
Q5lUoRk6FUeMjzSoz8VLyQ4DwV2SGP+UdG5x6qEZX12srk5EdEOXQHXpitg2gQdF
rPN7dsNa6HITizyZ2/S8tQdeCOHsjn02lWucK1rUOAu5NUkzmHuxCzSLnIz1H1Pl
ScEm4AShBKLoS9LM/iz8CP4Nj9xAizWzFCkGUp/8WECIenUtoTezxmd1OnVcVuW5
PgZUdFsgIVBaXcy9Q414fHp0NhwMRV6x4IBixMP+KgaXbgYgGS9ls+pm4hFdz5AM
XRpg18ucoEAWHKojORl+ZQ==
`protect END_PROTECTED
