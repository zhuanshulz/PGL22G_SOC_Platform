`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VNqYVVyWAHvntZBt4nxKjJ5iSCWTRfrSxTgnCgtOP6K9X0tjh5CSPw/bd/v51tUt
IR8UuUL+rBRpeIL0Ez7qsnQcMQLBrtqGK5eNCeujrXUf5SiAlphS0yAzt19zjVSU
wALv9MAUB+ZwDdRG/BmwamkLS1+bmxzHXFvk09df3y7dpg7rODwvmRcwAsOFA/GH
sA86kv6lxj9TEhq1Kgv880cLSh0hnrDmDc22OcYoy4A8BWm5Fr5gZ0TnoEq2UH7m
Ka8yXCuMlgUsDG9aTcsTPxUtOHehC7pZ8TNkxVKCpAQXX2JqiIxfdcR7ZhwMPaDE
1nHZyEQGRS9iVfH27vFcr2JZCPlD7VLqm6l9EWXlZ+xR723o1c8OrjAS+NhVrX1K
nc9kInbqWiTB3AlCTBSubDjX2HlI/Fg8Vtu3VOcUCBGf7tVYE8Fe97JM8W4efUqg
OWlmwS2vd8S/VJQ9zgh1OrpYi+iVWniwxlw4h1dhHlqzlmUA0C6j2wMvy6UyXZ2s
vjOla1g56MPPtXiwiQXu0w==
`protect END_PROTECTED
