`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
26fJOmry8p8fvHf4KLzuaMBXFmRyybH955LfJqTg7vuXnkkctQ6/tzcLg0qULf7N
TD7+9gO8ctdRT66In0gRQt03+HMQhfjx7HyH8Tx4WZFPC8VzZtXruIKX5XYU4mh/
olvNTFLGpCBXK1/eSgWk4+GTAm3Pomp0WXc7JAnJtyiEpN/fYkueAb6QVL2hC+Bq
Eu3fSihjYQUeo8jW8C7nvW393BzqEaJKj50ggb89FbNITHs/niiv7jdGxQGSp7LX
uGJyFBZ4Vp0hYiHR6SMvX5+Jx1OBHowGoAUwzQdS2kgKehCeHHSfzG/83CcLjBAB
Z9mojHdFDTY9u8bQFkDo/Y31CsYOYQi1ySoGygQiQrI=
`protect END_PROTECTED
