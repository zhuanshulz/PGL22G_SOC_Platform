`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KDWa19Sq0UmhSJHZJ80QZ1QAq1sY1+P/k2R/IcE+VPsF2ZkkB6SwRlMJPCuz+GY5
sI7ckl6eILsEULiozP/5NE02hSLXMUAB+ir1etmX0QQ5q9A9e6YVfZ5TD9f0PKbw
grwdD4CcGKtkQIeuOa4zQIk6wJTce0bb3cJnRmzOtbbIeHL9Pct73LrX8HijuDI1
kp8XTABWDMpjk2S3gNzP/watpRI/P4LsyRv+JJ1x2d3sVxv4UCgSz7mhMmWgWssZ
ITD+3urLD2A97wSZ8vqNlg==
`protect END_PROTECTED
