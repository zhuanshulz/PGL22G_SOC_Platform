`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dSEyixAuqQ6hMYPYBa2QVUf4OxyWdLhw+rPvW0tLA/4LNHMr9B5VBS+UP7MjvQ5G
L/RQ4f+eErwB3hxzmOe2qoY5eRRp3w9gre9mCCJ1M5GkLB2KaV8Q0GStiuIi1Owj
1v7FfEuvdddPgBZtWPqpJqH+/2TNbOjLp84O11+9aj4GsO5NAnQ9ptjLRZyOqYB6
ZGX6fL6CBdSHhy/wgmfN4KgcxDT4UOyOrAktpsZa0/I+0um35phUcqz1Y/NqWCqS
xIvFVLjbGevNQQmuqxxvPMadalL3k7v7gn09Ba5BiCjW9GC8wbl5g247hQax71Wj
w4tfSrPIUg5eewpPJxzshDIb9TcxZrw/8vWpKymw7M53+H/TM0TLcijSgdh+bN7z
8DbmZz7MrhaBUtdxqMgNYEXXLn5bNjr0DZc99ZTWdbocvGOozWC/PCy+z4eOonQd
j2KLQD1mpQ4ASq1TOcV1j4UtXwCi6IwR8+n0XD5s/uvy9dFz4EKift8BJuKil5Un
To3nhkXpTFQyXu/W7QvPToktaf7uxD4mWHxqwo8orEhYIPO20slI22hzREjcTRb5
BcFQDgQBetVYpGuGEqbU+b6dVR7wIUSqDLGMtl2Hgf4DeI8jxepLfyuQ4cUEN6yo
dRbAwwRZPh5i/xj81SiYbukamEZnJHMJD2JpNZ0l63cumUPhYHLzZ4/UL4I70d8X
D0csaEcFPXPrUKkgssA4eFmI7gLzK51iEf6nh6ele4S6eSA6JXiDulguUbP+fLJY
wq2Psz+iuKkXuYuS/RCbCGL/wmUUmva9EpfcJG9oL63S3wkCP/8IcnGHvV8Z2Tlp
Nq85oe0aOZ3GpQHKMA6Dzrk4pklzxGWlPmttNlChh3EkWVP7Pkrned+Zb15TYSDB
OYgADLlhtugHOBsjGzF8eygL1+aBz34g3nX7YhCAHCM1pIG6gLZkvYCy+0Qf0Med
eoIMb7s+WHBLMl4kR07PolyzWrkMqCZ5YOjRcwxRdxvDrU3BiJsGEysR0EpBWkrj
Nz9TVDS/iuQkvCmTdS0aDQ==
`protect END_PROTECTED
