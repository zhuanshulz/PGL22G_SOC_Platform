`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LMKuvQo7ZQzBRQbE5zXSfs6GOQV93qaOSPhEM3U2nkDQWqYq7bTREGoqZDU0yj6H
ufH2ELc/xcxsWEHk96ke1v3hwo3oL6cImo2XsZiSaYrKpn+4nKHTZNyOQZ1q8PcU
8a+VXkr72s8v4pgUC3RU1xPQOrYQd+bImEoAvy0wO8LlN751lZGpQAAZlf9n1XC8
J3kuSXi1SgUmgG8WiA1g7I4285W4lQbAPd3OcNRqqAaos81xBjn9iUudXR1PuU7W
g+eqpHCgd1jWzxVc5AOHixtGfis3S0R8MzNYp0V+jPIFXm8SKtEBd32e8RC47OC9
LJCClDAmHriWKT4cgECtAUF7bzrSCSy7rSm0JOTLLUz0pRjXwJyozG+Fpnrozndu
qCxDNGuL9sc8++OdPwXTE/ksUdR00GCRzmWKQqKi6eWqH0GcfZFAZ7MuAWK+EG7y
HQ0DB/le+mUaW4Rxu6uyVXN/46SnBoJI8dA34bJiJkrIlWQEcr35Tq6aD2qO4qQG
8stzh6PYruL3qdutbxiTY6XxNj8/g+Tn+duI0ZZSi27wEZfmtmVEa50wD/KwcLLb
Kh803JK+yeLEzkAaJmQ3s+D1n4/lb5zAs9ceX3fC+ffgxMt15t/WICCEfARO2d3V
JSavXQalNhNe8cHSmpE9LE1Uqi0EoJ8svwBowPvOFgthRxVQXfPzbXr/yGzTo7ga
hIMn/5u/cj22Gapw4RRNaAeZxboEvyNSMBXt0Pi+YUETQMeJRz8OBucXxs8u3G7b
RNYAcMf0KYJJEXPnZQ+423cv3jX/JQi2tP3NsyZs7E4us0sHLPw/lLJiVFczhRQ1
ihhKIIfwr3ZHpxOokLa9CcqlK81Zdu+t2JuIiXZkZ1LI7UWLFsQP77PH3411thSW
y57O1R2rI8RQcMlhq2JLTp/KKPhXHuWCZeu8u+saeDX664B32xN1DXF4mfLPDOTS
vBk3+RgqkLgLGx0XdwPrP+oLGS6bhTYjPr+pncbuSIY8+lewa2iWnQikUXriDg6W
WF9MIHmisgalwZFC4BA35i9KbdYRsH1RiC3Y87hLu4mT4/UdQZ7W35fAbu18kzrJ
hQlGmg6TN1ggInwsQ8NTR0Q0M4UVNsyqnu1GkNlo/E5Nos96JejMwcNXPHCNqSMM
CydK3FLioRC0CZpDDXg/TA==
`protect END_PROTECTED
