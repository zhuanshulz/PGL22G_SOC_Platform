`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p9ON9dTMxQra0eSUottKf7Go7FTUYooan0EBL6ODKvf/E4htL063UXlYdp/di2w1
5HRltHYa8zvHEE6ijb/H4NaDG4rb8xxGnbW+iYBCaGfWrtgnkLZhXkzexR9OKh08
JYScR+AO8rlTh1SzMbq7sHlghBxntqhEZDLSuz6VlvUUucLwOfVkfAMrNJvdePCP
LHjLXn1zHwAkcf0PYe/f92cs4pRGfbMpQXcOzQ/PszqgGclylTuav/PKts4DPR23
fG/O2UGLM6RkHhvIXyRaBAdw5/B1I32UexgqonY1E7whzT88rGfmV3DRwc0DT5Xo
gfCWeX85kvmV3HSGQ/kJNgzTAY5746p7Jks1Kb9NJtUSaGStqlybdSanZx/aU9qZ
7RhEwHfSethPNukUqU6ZTz4m9VhUDwGjKXjDebMjijlM8c/EbOnb4VKYZ8N2ZtRA
8WJtb7PywI/fWdoTqrxldp2UOCBye5ynUnTeco+z2Qras75uo/JZU1GNivXH17ob
WSLCkBo5G+uGe5I2KbOsvWqwSWx3/9FoRuRrHovdTl+Mv8Ok/8U9g6MXGhxEaGjN
wczWCh4nlqysyeaC88tYvc6wcQYdmdBbx//4q/9l6fjY8IpaP2pnC6JFgUQs9NW6
2VwRmhkEImLSobupG4C0R97BbPZXC5Vq+tqEhD51ter7fxOTok/INHDwcQBhzWmB
9Sl9tGkQaaVUYM3rqPfVW8Xtp2uN+LUzbqRy1uOX/sU2O/+F1ZvWntf7Sdnu2yV4
WyIaNm7f7smOfvVzpDEkqkthN8h+JQjQ7OBJ4bpy6D+8TWJngBkT0t5lNJtW136B
NpD+hrpGqQg312H6uu1AYMVT2Cf8iSv210H+FVO8/Q7GBm7KPNQ1Q0pB08bWLs42
MXSr0zQbzT0FysT3eBpC6M/ztM4Gm/vO3qxPVluUZmtbO/7bEWvVHaSN7oaqQYk8
GS9V3tZ4HKoHO0jjre3XVegmqsK/AGeKzZw0mBz6EYNLMHraxEMzjZ5EKcxRacmG
i7fAj5f7TvLnW6KC1D2uiDFQR8VbdpmHf3+moMAmoPMUbkFOadWkd4Q926OeGDDq
PEB5y6nEkBYMNWZ2bgb1b17NILHzM56Me0pz0O30dzr7LKgta6i8BDp1ezlebpGK
y3RQ657tAqb9tJ81/hLy+l/BEZgU3tUXagauM1H20N41P9t6Jrp51cWsVVawVR8e
xgQBSpIZDL/gKwEF+LLQRYvrarbKzuJOk+ZArT4CVSzBtRIB05CJj0GOoyYnEngk
Ntd7vFepwapU7FdkC+/y4/JqWLwSi0hj+4dosc2B88WdYYQEzD1+4cL4A6BW6VMt
EbR0kgUVGO6niDQSfBSrx3EO2ifJEcdwmkVg/jipTnbSxMNzzqfZ6EgwlkiOF+Js
iyBhpi3VU15LQbcZ61SKgbWZT5PBgaekkIWwMFWJA9NxYBF+m+PnvGg2wRr+pv0z
UPeLikZ8Ho0L48+s2G4HFaS4KjiBPgqPp9By6IvWmayO2ROm76gYZBj5cGzntTK+
u/Hwat9UL1NbnOt4uhTnSAQh3Pqvf7QemJGBdQkV+322g4Bp4Er5Kq8brt+u7J4N
QtgomQKwpPMgmxvsg6FNNRww0L+dTHMllKfo6Iihx9w8UH3LBvq5NqlvtjCpbf91
7BbrMTEcNht2vTrbF3QWASfw8NY9+Hu/uIF6W17h2tgwzKQOPD6o8nnABLxNy1H2
WBuxrydWx9b9/c8Zj2Lx0vHxo07E7SaugFausk6CwGt99Blc1QAAf7NJgIBUmKc1
MXJL4LUKTfzwv3yUp6YSwxfYGOWxBq89GZ0qNUYcuacYXdplLnVLd1469l3siKKZ
j4x/FrywV6ivkCc4c0cyfXtWWKXXlzgEkUp50sNLnjBcmof90+rK7zkwzHfxI56D
B67K2n1DP+qiiK5t026ysgJy8f2TxpoillKrdvyfhvU/Qh4E33MVBG9vhV+0Nou2
VG46npUMw0W152NaTkS9aBRmG6XeBolnEEAM3fM63ohvPDaISzqIGCf4HK79hPcQ
YGeT9LyC8RlGKKKbJczi+4J7rzn5HJzHcaQfzaqwhiWZcWXWPj6UyCNx7ibGuf+U
dyZqIQSydPVIuIJ70TcMoBo/jq/pl2K2Z4tFcfO1fwe2qESmq9hlZuGZHoTQY5i3
GFaxY3A8vVMLrnhge1zvquOqw0tRX6ldMbROyVzyAMiZKCwI5DSacSH+gHILJ7uM
9Q5IvOGF3i0wtENSy2pnuU/0eG2U2NtUj9becSPdy7j6MXnxtpSBU4OUXGFK8opx
rYpIQ0zKVWdE9nziVTEERdkuRO94gF3Zxln5E9Qhed3uepS5LILND5aywFkDrebS
ixvPMbBxml6irA4zg5ElZ75Oi1qxsW0n+UkTVlHpmSN8LMjLX/RKvilQLaG9zv7A
WWddM35XF+IIpw/axcwEBi4Qq76RmKmJlojCdFuJ9hp7lL5QavqQI2W1tQj/n/BF
12teodse9MFx+quF8yyvex5h9TDwQ56HA1RQEZejEvu3qXFqCr0GemWoCQQiL8ut
5ks0ocP0YzOW1dqx8ES9zPhJ0H6XreGFxGs4aqSWjdjlCOwvLT9OH00ytFxvptvl
/KOMakpCxoMIXSJipZOIlK3M8oJ/Hv+bbxShCSY0jKmzBBsRiP0q11x5zxStkI3w
fhBLMmQiidToQo6m2mIgQlycq93SA0+MeGPYWfwZIYGq+V5E4N+eNGbb8K/fIlSI
zabKt9ny+kypKcH5BZUhGvTMrMbwV4r9GMD+0z1RholcBSVNzyaPDrpnjxmPQLWB
VN3Zcsc91N/u48k3PXprKJbN/lrPN9MLPNJcn4IqGRZ/zAoDSeSZ8Ulz4gwMUuMw
sivXpiEHlQH41aB8XTg+ex0/MeMO11ZE8elmjIxfFWGADDknPlJ7sAaP51gpdtVa
S/ISXLWr2ZSxdgnxBC6GRbs6Ean7y7iCOb6u4jdXLmZaUlugYw1LNTPJmdf/h5TA
d2TG/6aoYHfJIEebn6b687nM+aQTvM/LbyBLQBa8tWbxm8aW7bnuRefxh4rVyCMI
jpiDc82P6saSampciocxTGpxSUr+zPMWPCnMRrg4Kp7zmyW2s/17hAvFEuRPP/hZ
jifrJf8j8dbFgBwCUKuVHNQQfFlZ65vHyLFH0vWxhtd9kFoe/jbKrli8QAsgei3g
L/vE4W9a/UmVJYNGHjkWvcmy7aBhhCvAziCrZxN7o6tx1S0Ac0vQoDYlRBh3X1Md
N+TW85PXIVQRKnYUXHOg5Lkf3YoieVS05Ca0QNig0u9w52gWb+UXaD+YqQvQl06Z
l9YqU74tioJDY11z38z8wA==
`protect END_PROTECTED
