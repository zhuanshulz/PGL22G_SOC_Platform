`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V6Dhg0k69LT7JrmRzTh6JDD0D5fG7/fFYWcFY3KoURqE65QtJLMTr4TdkfiS4mMi
TbWDxMLkJ7s8UoFqQQSxPqEPlGsSYszx8X/qXfrUiIygVZUKkaqhglaxGdEwzi6O
ZMAfBnxgOmDGT7Z/Wj15lELy1oRWtoNMwejKx6dgFTgZpL/XpgtLOvlpGCjj+s6j
rxVBW4Z5aDsO+04Dk8pdZsBft1Ay8ckg1eWp5FC91jDxe2VEgmArUNFqoEH+1eV7
bSYmqjrhff9l1EOjTLtOyAqoHATsT/XMRK3H7QI/aeQdwgnWHEXknPMgSFGqy43l
Gn0VewSiigQH+jr9BXHlG/RzF/zKS1KGPYJs4HPoPh8+2/wlE8X05epx90GqY5ZX
dvyfpCWTt0S8j6FVXflVYNel2WfM645Pk1uksueI+8rAEg/1UcM4des0SMH3zFyY
/+770S5tZQ/oI+yBsCj1XTNKDkDPz+mURUS+rMCqwiwGafj5mPHP/vAE2xcu27wh
`protect END_PROTECTED
