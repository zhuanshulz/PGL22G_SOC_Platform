`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4HI7N9d/Yu0MMF09C/M1PTfa1KteprQ3URvmYmUCpv4gkpIqpNZHHDuh623ckiE7
h6twqX3OHcb0M056DCAYELC/PYFib3E1dDcLPhcStGrSYAI6QFJyAjzpf4meWZHS
eoK49db/I7RRNmBOHfBdxR3vXme8ywaC6oMSW+r+bDrfbhc8EUTQeRscza8Xx7zV
FkvAcgW7S0ET09CeRJvRHjTuNKIvDQiAxl7JJr6M6O59ADU5n15CPBfPdnbqK2ld
/Qr/GpoCaR9GD+4hm0P+qjgusVkLGfmZgP+KPMzwLAqLnsYqPF68fMZOfWbUoT45
1tOCmkqlz3ZxavkiynaBYc0E39XZf/gaEWWxZDnzZeESaBM3LFiF0uku6QsFWgLU
868+EYHQyTARoQlFYE7k5BMmVDi/xGP9nvD2/g5tv3yd2wb303aNK469AMNkH6HO
E5w2Kbd00mTaNQmdaksOudh4AmabgXj0NAIWHNSzc8h+v4RfT/NqYc44JTyouc80
sa9qjbJsT6w4mzjYxl9Ss9PwVy7fSFIcdZ0DWmtvSEGySVpxYzcU761O6NvK93fA
fBPWJFwQ8Yg+oitGf8u7tbZT09avlFz+65+19tTFdCPglWXFnyV/mfC77u4VXJ6S
szRIVt/AJzsoRoguDqEZUyDev1xDZ3mRX55mylIEGl/HGcFqRuD4ILU9g9MvDizQ
34sU+4kxCT41FeIcgNVuJLTp1wJvp4Z0/nK+GxfDvlngGasibjenEd7trmp6p3BL
s8Q77Vlh5D4z8BfGBoMh2JZ/zETUkTVo5Ngl8vF06nAEIdEoXIQXGaA9wD0DJ8mT
f994eMapO91nOxFyMprGJB6HBMiYhzC4DG0aiTmr/+Ptpxb2Kr4/4n5WMrLr2dg0
Rj9nQthBtKT+7jwGHm8eazDhlZQ2uW+fqcjdw37ZvRO4y1oIVNVS4SnE8BTHUFg9
2kGm7bKQhvfNbB1BQvOCQYeirZ4KWrl0q4TOY7P7CEozJ0c+EIrRlcvMdHmy9zqJ
EprOhZq+SM1BZ3bU4lX1PFfEzafJ9qEQbMzXjbMoASMBdH1TFpaS/3kLGHbBRIGC
euJ/zXzs+271Zp+7pQUGZHRMKvQ8ZwtdG5FOt+9bJ6KmR/uUvSPVSCQtHAbjLIhQ
1CXpBO4Y5DO0biqbin03Uz9m2PM7B4Zi+XbxLclRCwDdGbOn0m6wWlr1lpxHdCHY
HbvCTP43AqA083bOW9j2tFsd8wtHdHVwvt532XXa/hzQwtJdwtxlCPw/jdcIQ8N7
qyrKxGr3Cq7zVEO66BVWt2jlCNt3BP07/bFQyVxT/jI4VueWxxIYowJBJVM1Hi1v
kEk5TKdk+vUVi3mSILMrK5djQcXsOYJpQjN6k0r6ibzRBvgWNqXoo8C1q4rhZr1F
0R3Wj6yQygthkvAPGQHoo3n6J6B2LmXpNZ/8uIkFBziGnhny6EPKwXFvtWQ7Cjuq
CSNfOYeaIg97EKSmXakQmNhyZ5SwMbbWEWBSPJm+mguD7YfsqGrgzNDj6TMlF4if
UvSyU9SxoNyOGxdrhHX7v7BDGGc1vcVyoUeqj0i8vujIWl4R3d+UYSWbf/RjcbKn
KRRXEX80V2gyVrcnNjpamLkH3FQC86jO53Y94eSAKBe7JonkZO+03F7IV1eA6k8l
5L5PhWiZLLfnGHZGO/UTGxGFPfkb08mzZ0irvpd/PWl2dVtpT7X08a3a3m+aYvUN
UNCNeIg5MAi2Kwy7gaEmOrb+yC7XtBbN5Ne3mUxvsMmPxiAoqAL+iwK2kUyOiJLC
ZMaINIUSwqb5Vz2uswhXgM+AA5qweXnnFjV9/YQOFrMzn2fJGoR+37SZUMnKD8nT
`protect END_PROTECTED
