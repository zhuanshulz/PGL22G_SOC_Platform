`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0mhCFVRFRwnTzywMn7NytBvBExnEM2Rm9oJv2MYTb21LXocR9cSt+ML9xcMbFvXa
LSvNimwEiQ4o5w8YnYCmWEuIDK2S9ly2ivwqsL0HkfT9vWik7irBPLPWFjPE/Qj1
ja2XlQXkK6Vq0HVmJDktjCwc1hpQw/b+6vT7K/W01T20QrH/bCqMKrrthMtUC/SQ
voSGA8wLz3bp5KnMehAZ6gEMtsjpqZ2yl59ptfuvo2EfDPF2G+k01kZDdjUqHu29
gsKWeOIJ7ywVdJ4VSqLSY0HiUN6vCMaP0NWPz7N80DTEbXtKmi3aEg+wwltThK9N
rz5sNwih4SAPFK3qi02scl1Ysl2zTAMNKMJd8geLVfZYyKggmK+oucP+5yChwv0I
e04WIrEewahVztzL7/FL/UqIud9CMhc6f2A19gePaMh2VhKJx2VQ66igs5BKkL7o
yTGpFC5bKoYY8g30pFTHowIoui/71oQ9icFUSmEtG9pDUVByAg00uutDtJAsU7Gl
xgng7lsHMg/KxEs5JALjjc1qvWUtyiJPWwJQU/Spn8yrBDWeiBCxNwoMhQ2/InwO
9TGQUXv8tHe78eciBB8Odl/5GxNAPIpjHP6IsNWI85Ccu9grqUD5Lh8n9cALai5D
T5YMUji6QJTK2J/EgWperC2Vgn9L8onaYzSJemDdiURt1PSkVKX+8F6xiK+OFqe9
139YCbhsqq/tmNX3V/OIWft6/K1qQoJSkUFa4VVbUxhTmwDca3wVTT1egawFNKL9
/DYhlO6+4g3+IXsTG9s/KO6TyqhzoVoasvJUrP1THneFer8RYq8LdKTjl0Kt6Dy0
pVYLZEG7l2rBa2wGRlyvtgTo2RwgoaIHDz1aJeDDPWfycCaHGihMhlEF9OZoyMkx
BET3GQCKViLRfJaUhmZBXupNsl7xvItOgR5Wf4Ncw6r56k5mHqo63rSmc+SwZx/O
xzurkB129z8AyR8KrEhepRQN/bsZz04W3df5fKK6R1XHcn2MtJNnjVE177lFUhzS
KxoX7IlzL7UmAfLFM3BdOVTqstMqMHpx3t8LWgZn8+oPQFOGcNhqNukM8iLO4emY
`protect END_PROTECTED
