`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
98GlTmw/QVlVYrL/0iSkb+Ozc1U+GZWHMIIJ8FqEH7UQBqbUeKwVCa4l299H0lni
8Jb2efbV4VrC3sHjt/VbqBZCSSexUWh0iqzC7mYRSXFgYYkvDxD0Q7udPu3z8YyL
55TR7DQdBt3/QCbGOMlBj1YllqamHmwk/2wP5ad+MmRy5FFNRVDMviKdw69LSZcX
RTUAcDZEOqlCWeQQ+k4A2J6Ej3bxVquDRn8jvPq1oiKuJK9KW2QslvU2VIbfHz5m
kdZD7ifx3fmX3V73dyj4MU3xEuDcvoNPTjmSaB4UBd8=
`protect END_PROTECTED
