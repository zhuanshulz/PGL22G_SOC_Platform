`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MXh3PJLeyHf4rOX0ajJSpBEgtJ6/bgbC9bEoG2wUg/vaHrDBCEl0/XfM9ZZxLVts
WioS6nBN6Z7cdLsjs5gQAxdLmwQuPPctStPkT3b06T0pqpPcTknE7qlRtvkTaNl3
aKlv1ij2luzttkDVCndJYCUSK1p05MJ980rz/pwHpcsrfPG5n1tjnzwqqXqNly7n
l+F9TBmmrH6bDGTDx+5/ixPU6Pt4b9u32nY17gAtIisrYImfB77URNeO8o/npt5M
96H9gK+wJFBgq4zc7ZNAaiHdHVVeVVjbE5KiUSDhQBw6gl7TPeMCuj0GCHx6otDC
C7lgve+wVxVIwdALzV78XXnqQghAhgZWLiH9dnYGNc2UpUTYMBAkY67+wagmF37b
Mn8L9K6Z33LJArSWa9c5KgA22BNYx70E7kabsdvOUgCOavcrvniRTGzCFnQMXGU4
xK1ydILZetvlwkVhqt700xCEwtNqk97hlYQWWVbEjobGSJ8Hwe+JOpSiEQ2Cyt2s
Y02qxGGZmwSADe6H0hdf+/CQvZF+JCUL7yyrhl1Z6GAyg8z+i+F3+OUrc8Uj+Bgt
QifrmrGD1wQ5RCovG/Rj9kIoHT/CHG5Y4iDWYHjzlxqcD10IyDch5PnffX7FiYya
PRIcNOtUs/cmPUqBD9y+2nHfiy8tArk8R9FSlWeXEl4VqQcK9AmUfFrT4gCg1CXx
IsK70nBUopiDIpMtPw0lXPxop0INgOLJmfGSCHc17J0DAPscqLhFgD5S8z5n0ABt
QngWBJsyjgluvDIuy7mjoRKP+S67nQvcYlBWJIGxTakB1Vpp3qJWw4FiF+DoS7bq
sLpbNiAjonGQ0YRiVvM7Jnx+5rIWr3Isp4W8WQPOZvMWHXiBVUWokG+3GpMX+TSF
v+0G02rUOxDGcBZABHd5VQnVnsDROnblF7GDGMiRbz5jcgOvpqDswXpDYkTwe0/U
5kJ0kA2aO1iev6/hWa6sBLP4YyB+1PoVkyrT5mMb9uSsd45qZESItVxYWkFWbAqE
pn+TDbIg9UzLLfR9WxPTFF2mbUew6TgJxNx22dQI53S77mkcr3VWyZH+Ogevl4sB
3HwDaSZtNL3d6Cnsxt3+3i4EKy+T1vk7tiq82cVYWGHU4z0S6GAn+zSlsUUHqAy6
IiPDfGRTgfnsQngskJZLBd+hTkkc04jfsn+iyRkk+cJFYJwGYdxK/SR/PTUQDU7J
qb41dEEKqZx3uy/l3cyWzFFhcyGTHfffeHgKssY4Z85x21FLpXz20C//hVIHaaOW
qsW90DxK5mdrBY4T0wvVg62mIxX0ncSUjYISOnLg6e5DmDD3YFoKLCLJwgR7FwHv
KEN72P++zvemnCHKsmE2avtAEOYTsoH0MT08jGeQc34Cl+tM2SY2iKN/RpuhczgZ
/QQWDEkJ1rw4gt2VIaujjdcmfviocN4my697Nhb0//12LXjYnW5yfus3xOtUg7gk
bd66p6mj6KQ+A3w1gJmoY28F1b3Yn21Y5bDrzyrurm6UDdTddg2d0p3U+dzQR0zZ
kbVt+qzfcerlQemOuohI+kI6C60J0zRbG/XZqQ3iE//H3S9WoiKw0edwn6Z5GIjB
riKqLKV3G+LdoJQwLKJw19ELojvCAJul6ZwFqIU+nK8o5ox2R129OWx9OJYOsHRi
1OIZ4FCQDYrQhfGbEjWsS+N7eG8P0zWZEJeGMziInuRm2EqwOmhF1FX1GtUYZ1bF
veZJ3BVcAbb40a2dzmQMisH6H/w0FD2+Qbjf2N7jGkU7Q/HOS7exuZu+NCBnMFuL
I01so79S5YwNen3IqVpIRDnU8514BoEdMX6KxJ5cSHwu+GPtE8UsVgS2dRGu89yP
lyYOx0vsLOB4scXxFimAxaWBgjZP+BYQoI1MyEP2GRdeMPhXDypJD03QbRZfd4Ci
Q1F1ZgUMOUWMcMjVk1yv0aojJQeC4HNVP5Et4I7ocdmg7BCn/qXzDM/3UAwKXtXs
1/37Ft0BxivBOMLUzmxdP/LOjIfL6BumRIp/T/9KhfoUmvoDHOR3+xvMHUYD2i3Z
WWbvWWqU/GPiYciR0oaB6pVwu9YyENg50/s4JJCklPvnCIVCGfV9wUPlEGAzYNa4
rJxECMWT0OqbVmYoFkc/5BUEPtP0qtVPwmRn2B7H4sGrcLNz5iQOTmP4yo74rD0X
17H4SMYYK4U/LtgP0fTufO6JgGysbrZoMiqFJe+PKc/TdAV6gUuxCogyCYhg2oEL
OzVTgMux6ozdwe7QrfF7Kv9vBx2BMDeXrg/5RUw5V/pfSIXZ3BKmzcMDbFtESTO/
XrxShf2EMQXSazheBh2jRmpe56D8Hn1xxrsOlEc4wbSgJYFj3/f5SgzATOL5bLS9
Quyu9kU494s9K1FQ+JPL9H7ruUYtwFQTkCO+nTlEd2AObaFLBhvAOO7p8/EogmL1
ILklJEnuducuRQRAld4AlTNGv41mP46CvYCjPpXiyfSaWo8hBJs/2XOM/8LS3tg7
OlkgFeFuSqdVXJv8BvylbKdAdulo+kYSKDKp1NQbMqtIDY/s4uaE/rDJ1VDCkp7W
f2agf7298pA3DxLMMAxcBBcEomy4pZWPkK8HEbnc9+GmvcVaz9jFmm47MDvsHsRl
k8kbjqwDosq+36MUIIs0NpfSwZygKr5wdEIu8AtHvzdxPgQOPnCPabaAIBmkOSyT
ZryNOtBV0w0s/niFJr1AoMKYnF+UlxKfdr5qSxrAqN8v8h7oMT7LAKJm38eF2rYe
+1JUaVgHBBM1F/gw71PBjP2Z6LUuEZp0caaEjoEkRs9UILayVuf3crQZE2dObDtD
ipRd3B+6Sc2H9wqOtYbmUwzp6QjJS9tArx9lAYV34TCdsM6d5aV5vYGEoOErXCvc
VPKj/3y3RPHO4Cflda5ibG7l8reV2yEyrVvaj7cLn+MlcKHrLb/6YlhjyT7Ix5Bg
ojuz7+mtJ1mSXs8tJG8MIz/DhD5e5Uxz41S2FwxJV+01jm78JmVE1Ekey61mOn0s
oXdrUgOMSKkHLZIdkIpQah9mnHCzJ4RotujWaC2e/NOKTzEtDEJlZVBMCcxWGzVv
IITmc4/z3DqfT6RU7r9rvUAcrznQ08+dYSYXFSB9GS7l0jFLQAxDHe3yh7xGgApW
rMJhCEnGb68alBhml2G7KWIGhC+Knuq66xm8739pmrNgFa6XEd6W0yAkUim8qVY6
I26gL1T3095KszMAqFnS71pzw2TDToaxdE1RV1hKeWn77fPEb0ZgIUX+F0AStwkJ
TDcNdR2+PWOv2DR6YUFiTM/+A1qxlLmdbeCIP1WmIW6PEZpG19B5CNX+OgVxDcmJ
npnEIiVCEKWtreevcz6SMluk8e5wCTtrSan4fhk+rEeXgOQ1PcW5EGbvJ85ieWDE
aOeZLxa678bQBVJJtNVp/omcGXg5iJ7K3X4WRrFjpIpaTnLNX6vrLfyJLy/3ullX
iVaUX6S62aORN9Q4cwxqke9332L5sNs+5YdNpg5zCHbZWx6HLtHQWS9qG7knIZUT
w0q80rIRbrgqT6nQ3SIjLR5+oOB6bQC/5MSh1VeHqAc8SBoSp0g623Wl0FPdm3zb
wfyhgnonNW9Bgy5e20XACJr6ZCgqy5LACcvyUQKB5Yb14XZs1H2uomMzfviXQtXS
sCYokjnp3n8hpyD0wDFJdqDEas0fDL2wLxMo2DqQ7JADWanEmqvbHqdlCdrJDVW8
QkI5gTfUXo4VWmdBThN84OIZ5t7lCPU0ng2Vb0EnaJ9Jf/sw65rfLQrJjeV1RYF2
jcLWhkVGNKzIZk2Ln9UkybRXOERxbBrGp16NuCVyFdsMaJ9wYCHnx84APYwBNBGS
OVQBFJyzD0cVDp8zzjleWF4X2IrocPSJdjGm/H3/ZULE1u/MuKsYuT0CUawVagao
t6qqhiNpGAX+k0EMxpRu8rIQH852FZgL6XhazlLio6zN4dOiS1E7FMMWB6CajucX
nEbtb9VFsTboUIa5VFWQy2kEiwfeldui7pwWDxSFSMlgzJAiSGjs9Pjf5tjENium
/l0BVC8b2SNbIbfk2Xhi1Wj4fhH+ri4TFoT6havKYr35pZXeuMfREGppzOQNq9qE
Z2cgswAzaN5qbE3TE+dbEfc+ktKHbk7ZIgVhjZXvVFucSVc9lacE2omwORc5VLgk
XhE8s/vxy/rKZbCQMOT485iPf4cdZreljqR0PbsSV0rIfgOocwH4OagZQ4aeilgb
252kY/XpLPkzp1byRLNOtqly8267a94BbrnZkWeIAug+wq8D3H898YiUMSjDwxyl
8I5ts2Wlr1UveSE1PzIYDK//khLic6fJavkWvrR8lthDqvUfitSGHjA2v+MgOFgn
zquvfF+sGgDgAaLlsTn8jzbKIZc3kNTX/0LRS52Ut79SbeIwYokefU6CO7iBpkOx
3d5R1yrEeUGfG9tEmYwcaVPJyXSuVMYg/3dGCV0MwF6udDRsW2IWB4tVcKAZN6cX
uj+pf6cnXGp8V4/32hYCOfFDnofq6JfKwOACMmL9P/HpiZlzmsaJc/MCSoxuKzzw
1ODF67W1Md4+TcAUmPszMRkq+HqUqJv0kcxa77k/SfRU/OMUODZ+/fkS93xEYEIp
JLYpPgFeHTXY16kWEDCCKk8iuOuvYrvmfRqaBtRBAiopbFcXhl+XjpDSK44ynPy4
6+dm8x4WIHxDz4UBmmrXUfFABRPgthqvdhsVezYEgHaLuzA9kXxJR8cKaMg/i3HY
4pi4PH9J27Eghtj/BeFLi9+yLR5Xso46ANF7V2HYWNWiSYfHT335xP+t+4dCCtbB
/ZAdXb2ytveRBYv+PFfkcdadHlXpASvkWXjHyawX64pmsKepHdjCLMtM0YxbYuAO
7gVKkCpIkgiIzkPy2LP06vaHXSGExkNvgczI7MZsVKhtAvHGFoDGaDI3j/lA608K
L0iOoQaGsyUFtVqemt7VemYsXBuBBnnyHrHzwA93DP0sZ7UvvRA5vSWqasrT6qBL
`protect END_PROTECTED
