`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z1ZklWNUopJ8FiID/no4dnrk+wZGVVHkOu8OlmpM7+VbwyLDfmX6MVXa1xsCFjTi
Doz7vM41Iuk0MQxmyieNTzetWfQ83orUcsTrBh8dxIoapItIEFxkLP1xQcFOGVft
fDerSt7GXuKddWmi93ftGvmANJrCSnwLg8d76rAA5HnoKzNCPzJjgqZsQONdF0pc
/1UKzWT8LZ3n1Ur58wkzknJyN+FQD1aPpXzjXPgBByy2kTEJArBTwjcE1UDsAGOF
YjAJdpaISLZA2HgYoMTvsWSY1ehVYlgYnw5y3Rt1OFSCjTHnwoRC4a2lEYIwwwYs
Dj5CTGKQ8O//LYOGz8cI0kWV6gDE9bSYerTj8CT/oSttNUgXCEZShjFjbDlulBpY
`protect END_PROTECTED
