`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/kjJDlSfciqrtvLIgoH00ZwjmNanKT5IurRJ1RBcvwISW4EwaU8nlB4RKe0qMQ1c
2HOWUOu83mJzP9cf45aXRFwU9wPhFvSL9rpAa/Q/jUePYFBbix1rZ92COmx4Khee
rse0g8Jsznjs54TWP7aNhOCxmJDp/0Xix9lN5T6FIiNqeXZDZH88x/Dz8WpUHXgk
ZPpC4ANhKpl72/Z4K4QgdgY6T/dk/tswmsuRI1XMvkSTFJcRUh/HSd4++Qe3pjD+
WYJWt2H3ydJ2P8uZoJNyyFbWeFRIZTLFTWJnOAVwjTEG2lN/uUhp9+LCm9i4y00R
PJmcCLZX1W9keslYWANhze0Mo4zOtPGMpmyJQd+bhlLpB9dWb44dMh7rju1QAGds
CTVydKWhkVMOgg6thWXRclC+IgI4MGa0qeEs3EEHWr/EKJXaBsH/iyVlc7y+WoGe
2vzcrzgVCW0K96K23pVNTYzxLQkWsiYNkj7OiSmEU/cVgtOyJ0yqZLK/thho0/nv
Fl9bQIg4LJ843x/2FeQ/FcAnwpG2bwPYYmK0ZpS1h4Q7BWcPBXXX5vz/C1DLH/E1
oMvTCxhSTml0phOV5cqH6tVMIoAHpOSRL/MW+616mMORuStWClWCQrjS0gxWJcN/
wm1HYtOiLiLnkkiG7ZOJ1udv7EbEZry3YbeV524+pONjejIIqLhfKb5Zj1wNRd2b
gk7VRYdxSxUA3e7JFyiGxqzqAv0WUfYE7ira33cXI7jhy4Ft7ULH5+Ht/6Xno5Y4
tZGu20C2HIhb53M41I1EMog+/TN3fDThzYqTdJp+vQfSftkouYaeK4M5Qef3c4Fp
0DyP3IsNZOn8s4z0uilponTyjLXt5UzYa95+bZu1NHhX0xAWNJn010kCDyVV7Dmo
MM0nMCxMAEt5QV4GKdzKN2MhNqt2VfxKWdqwqumif3yv5yQwDM/TWiCQQb3uRlPf
APiwSE4exZvjxKqaswH/RYN54IuYnBZaLG/s7iVxRLRueT24UZSC9TtwicqlO+Se
mmcn6eNoFgwYbytLs6pLVV/Vw0OyL090/DiRX0bx2VWiVV5SI2hlSZML3mQw54+H
GzjbCl9fec4BDc607SDSdr5K8gi5/WYYyZ2SmZsuMUiranrOMlxijRjKiS99reCP
q9ZeehtuzAGdjthhdbTd+Dy4zUfd8+rR+nTfYoC9FLWqJvPOoEnrNNc8tPfJtx5e
YHKunIU23NZs7hzPPq8iyan2zS7GoqG3SOpGiTQvxjvRe4UTrHEjFLvuyJW0zLve
5piPzB/FE4/hoMaYLHMPpg==
`protect END_PROTECTED
