`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tJUbmXVbt+QcxwUXgPx17EhDSfP90IkMQm4wosYX5RF1R8/yjFD9Vu1VNevQpyeg
S9Q8D1QdCuSl6uK/9XbZQBt3NVW14G/wjJ0DsubThgiwixAKMMKo6jO/loECHP5m
YxjFJKPseY28PV0sEtVphvSQ2eIFCWVGjb2Rby1BOgQuH+Qw1HqQPmsrAnFx2Yre
+aNFRb/+BE3DOYpzgENS/EmqGxMjtpgTWSQWCs/O+MPOGVEsg9mqhFa/F+7xC9ry
aMFDJSUui75KJRLr7uZR6B6NfEeOBnUButIoqK5/8n8L+hgJp+bvp/kZOFG86mux
2PJ+qGQS0TVwL1/41iBZr9AfDVoaEK5o2y/WBxEIN2Bx9WgXnCRzTrluuxtbxF41
uk7jBSr80XPcOU1CnTrTQD1oAeRovkO3EJjfY7O5cABetKdlyZ24YLuKdQry6SJ4
nUmyNRGmRVG1+IjRurfofc7/21nP+V20hv5JzPkps7X5bAMM0qwcei7UGDcaQPsf
d57SLciUCW4lMBminK/wBrt44c//OGquXN1LKaFUGQ8pWrR5j7p0o2msbqOAphJ/
MRs9QyT6mFqkzmX5eC0QZ/WWKbl1aLP3SzY7SX41hGp+E9CA+nVv1g66C528vOya
wt0Ae+ane8KEyu+kCvdhbORcwdvIRUKgdm3ZQzvUvaDtzA3+fqTXgCDKCTZoezz7
BLnoeiRr+/vBNH8UQYxL4Y5fw7lsGNU2BuIe/MNjlf4ezM7CjBKTXkpO0etyTu4n
i15AVschkEBCq+V+X4GVlQQuhp/U9u9XiKzz2vC9xcWAFT6nCUCJG887mJl4BV6E
TlUMnzqFnH5TJ+E44HxHRACIFwFmf5FJKxzDAR7+eLe3EtCkNoWkJKauHUKrWFJk
MTAdc6dL+RsjaMRvfj/ZqCxwlt/qULleit+V2+O9hFA=
`protect END_PROTECTED
