`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HY+jX+3VT/qGgi1k51Fw2BUhNFrQLbm6fHpTFJaslpg7TUD1wiUYeaiVU/HwKZ81
eQttqEMbx0oYNICb7wiBdrMRjPCDxiClpx72HB8IPwhXU5z4eHgPp/qAABFhDlik
wqLXzNofToBJ2OZ9bPSy7TojsXmJgqA03JDugZSQ8Ne/99vJlu1POvEaNsJTNq56
Byb+1qUIEIpJoxEBfeudSl613uNWzMFwl6LaKbPygYC7TSt2OSPp544SLJVTggCd
bfcpp7NW64cJa7wk/vkbjWwNRsZU+ONXvwBbcvReTj6Tlu9+hId2K7EE3A/TEYgy
CcKlvLguM0cuW0O8mBJ4YYW1iqmWx5X5OP3WQUtl7OoQHX0rj+y2LpwMno4HSXee
pwH3AIru6Ewrmsktr5rzea0qkc7C3C0r5/0E9rMk1Ad/qtJOqv7yXmPRoXog/80E
+QNx6kSgmGL6LSDkhQAar/F0GTdGLFC5y44P9uS7aX9DmEXl4SNwwfvXXxP5cnLV
r4scehl8fmWXCGnlBj9MWCFV1Dum/0lOMAo8iAgrL/1o4QFphmibL3p7Svwj+RuH
BMM4OjPxVG1osDHPv5dLYfw2AvRG5X5TUKAi0mTQLpGXzi/kQ/KiV+lRTl0K0Fq8
GBolhZMt0ChoEnaFbUMCuzPTQbIQsk0jFEkAqSxvxFwWsCZQpCJKFfdIROrcO7J1
zHLS/xvNx7lnr28e1PrIr3b1aaJCm37pwlBBbsiVuIsxpfEiVeXTAkB9F5cY5z87
2ngE4iz7bLwN6nHNUbxmxcf5boDHoCcqLOkWUnc5mWsyQLJM14tlapROphVLZyKx
P2jepBt3NtVs57RxHah1QSwr86O/h3Iq7LDZRDXqbhqYvtLiUIz4FkSgEiG6d3Ip
IxstKvYlmVDYyt5scHpGX8uJ0cRyb59I27Mj2LCus2jIbtSU8pHzpW+Lx3kjmsIZ
E2ay3HIbbqmmRqa+sD74s22MDTK8ZuTLLfwScMqXBnnvDeQyCPLvYfnVS/qbxgAI
t6+ilvHLaJewo8zPnaUBPO0imyVFvLGymIKH9LL5fkGnGskrB1DQakCjl1V5rmCC
FcK8WmwsOlzLiKRkA+YixYKzWWK8xrK65fy9TcgP9L8k4MYKc85Es5DMHqhaVp7z
NKF65hkSSf95qhu7OJO22rfRKzzwwEbae1nR/TyL9b23AkpDeDDBUcgYCh0im0u+
iheJDIg4+jJTye4C/6zdfaBgv55V/3ZdLCUvPh6D/+ud0R0fB3uNew5wyfam6gUE
2jdzVl9JAfQeAax4mesva/0LtryAnxBiCkKG3qXKr3eUBhHtvZl52BhgIZo5vTCa
sKROfMf4KfXkl4RysMvm5lopiRGrtbf694+kI33jSo7qxoWoFe37Ttj/22uS0dBY
jwq9r4MJr/kBIiDBqKf0mZn4AlGLqroVPnmQDXhpBrvj3iu0V3gmEYFvS8Hpk1Bx
wKcrPjlzesFlIh5IHx/GeS5CzNPri8Wat4ak3MU8BMoQGmY2k4ta4LQyuobaA8NL
VewLEP+TJnb/1lrKi7p/Ia08hzhsCWecD/lEP4cZbYKy2nyV00f3smruAA2dfaX+
Aw9Kv+FpbvjsgaH+QrU5pTNPBIK9DyxEew/QekS31CgRl/pEka6YHvFrAM3FjD0H
Jnng7lDGgCM3mPH0K6XCfDsRTwCkBcBypf4X5X9fj4B/VxjbFZP92FxmKdZJTt0e
SmOeUrExn7+/kmTGQPldPD/FHPnj10nythcfSOIKur9ROpeArbjwuhJ+MqD5a8GC
gzLCrbU0hDnkQJQC41z/1erMqlT2pywifbq4tMnBk3Bdot1vJhS6TJoIMsE0rTkx
eHUuC9dUDHkioOfH0GF182Ed1LCwuqEtek9eZerlsp2ab5B6VA35FKvjHF4bg9uD
jwUmSkbTqSzhDngpR/jcP0JBLUdfRnJXk5BOk9ILj7yBZwNm8q8d97/Koiu4Hvet
pTCwErq7PWRwl9t8rtqmr3CEl0EXYbYzWxa/uhaQctnGe58C2oY824/aDrkmmqLn
SWUmbyoh5OK/xf27j8BtHsBQCFqDLiS1qCCMXzC6TmtL85Fk3ijvwImLqtRAGCh7
OvhqB5ABnAVgrTd1bz5jLKbG6LM2+EQ8H+rN9HnrEyAmDBtwTn3cXQKJnbW2EuwU
suLNcZlIRdj1oejjcvD4bylp4PqNn7wWILjGMcqrDpaQd3ekdo4+nnrR2qQFmIrA
35O4uDN+6bSaxVyvAcgwjfxToMpIzLp2rSHSWp85nq0khI8C/dCfPxzv2RPDHlia
z92InyY/2rfSeCYudHulbuEJiebJJ9Z8A5kfaCNNlIpG5D8EqGfYvYkZUd1IBpi1
m8rbAaRQK8W/lt5cHG8LgtzQy6bs+xX7ctyT1fPczFMXR7seaTe0JYYQBTSNEyCB
46FibCmbyA945RW9eeb4VqDUmTcexhmXZMU6mFFtb6kDbvfKORlr6rcnX7HX9PNU
+Eza+v801im2EBI9NinzLJCzc0tFbj9HHiwJ/vXtKcFxyBpjeENRWoEOJLCT8FwK
BM3aBiPg2fD0N2aTnEcJyaxtsdhh0JmR6U0I4uNYqfou0qgonONNHz7/TSEs1bwU
/Y2MQoRWSAnReuoArl4R8Mhux1DHIJ27GLltHW9LEiVGPQh9mMTzkPoAbYRvvpor
VeDnWBNYEvz0HhjkUcx2iTGX4SiguJ2mutHQRxjE1c0FTP6B2ywnZWgoIxn0dCca
PcOjFAMqf83Zi9ta3gZpw1HGFb6/1EPNwMZYKRua33NxOv9VG86iw62l8f7qYti3
foM5IUZMvhyy93/Qmaj+VhcBqVRB7jbWY8w0hDC3rBf91PSVxpxA9VuTDNCPD/45
SV2RmGjjw+h385U7qpDQo+JwCxmbpsFDeMAXxgtnRvoN7eruKrdFNZUR96VIytfu
1kEwBM7xRIryftOyvuoHPRQKMQzkOHO/QfSgyu6LzB2g3ioMCIEAkmS61tuitBY3
fCEyNxNTvkQPQOTv3DgvyzYLr4PH5B76FqycNyei9u51rkBzRMyFGN/QkaFPFHcS
hUUOs7dhmuAimecah/zfDsbdmCeIDzmL/E/GNaj8ClkETGAZA2qLzX8VAfrcCybW
satZ9sQaxx4iHUP/i9huJRA+qUjBcW4R+ea0OCM4SMn6lgtrfyd4u9M1zzEWvxqf
dgeDaQNQlCme2UTTmMgTSFdjGXfwzB9+TqvuTPYMRqoR98um07WIoDVlKPjqVMYP
HrRaVwYOF6XqrVHFkTaYtPKqru/FDGjqHU6XNlwI1mf/Ch5dxZxiAoqVLjeVTlHE
jWy4eIQ6wucGgSeWsnVoSMGkaoLH4sxD215fzazyX1goiITGjsEKTl7Np5Aiia/h
k27f5gMfAbKeq7Vwfl9LrHi4/T01r23YhQ84IrdL+Mk6poS8XnoybrKm3xjcp2C0
dot/TDMbBRIU+GxUQM1O0UX1S29VB46vAxTxI0XYNlUmrowtEjBU+3OWhfvfkEY0
QAjFLarsFKNqKGUbcdS8sVtIEsrxTkB+7sTLHornFgScwvfHa6ygsHnvCCgVUw7Q
5/CngdpNprdI/19bgJylGOn8khrdm86ExVLq3B+r5I83subhx0icO+Jti1DMIzKp
8EYDJLA7aZKPLyKDebbO5IaxD4nEvKe6It7J+6oVc8ia/5bUcB6p78I2MjcrmLL+
zv0Eb0s/JlKaN+CelEJBcbI/k1tekqu9uGf2bnCb+3Q/Nn79DYly+MYwNj+o7G8L
UC9B03EKph9zHcPeOoXHj92+3uumA/P1gZnGH+m6pRRrJXUqFuTuP0eSnThqV+LS
etppG8Btxe0Zctdy/xI7zH/j9QrhWVLyUzvi1Yq4R9jDcwhsq8hB1dKJhDQfSYhA
EiHCLZ3iOaZkwlaXpTaBRKkCR8XJG3U9EMir/D4PZLzH3hbhFZmYuyZeOCyRWnk9
HsExCiRAdaCC8w5enGzrs28JVeC1dejtD+zZ/c1SxRFExzXWsMSfwdzqh97F5HBb
ZEO0nvbvJTmbmFOHu+n/HxV1BbhpcCVBtwLsZPGDeWqHZS6XynbBY0b3jFDiEYes
agdyzlH0z7TuOxQlgzCGPxPe5VNi2ZaWl8BeqL9ft+lrfxzbTYU/MviIoZnjqxVs
hG4H89AixNK07CloowYw+HZKlmW0ATwSmdW7zpdVIQe0rk+AVHcnUJ2Wqj4ruiMV
aatrOsgstxgakBATwaLjs8le7lnQHvHZbl6af/triKGJj0mgTbty2FQOyn2u5shV
KvYgKDlm3sroIv72+k/hPOW6VATP4dXzgCNhu0dsjGi2fB2yyTfPqgUqkyf5kwyc
Vg+6H+9cpOGj5g7mg9V7/G5pjNBJWRxSdHgyEB0nuTL4E59y/dZjiHWx5nBW5baS
+x2M6WlOuAandCNXCVxUfnxA372PZIo5Jycplg0cZCP6lFsbqzdo93XviDCJFNkc
2H7PytnEdgJvemhYBGbWif5WxAzyQSWWh/34455AVUp+KxNcMeyQUPRdBp8xLAEz
cfwjETM6+1zlyHjt2l6rTmPTc9PwpUEmAS/5YOt5PSj+qCJGJVFyGakFXX8WZ6EE
+JcFM1Rcg9YE38q9oi+wzbUed4y8oLtp6402cqVCyLotlfwMpeM/Lw1hehLodsHb
1475ZlbPdj6SeAoREhfbo7Glulk44JtTFpG4tS4BnZaWN73swRENf0WjeXDKoI9J
4iU5Kdonua1eJ5JVPhydNeb0v4e+LCo+JmJwBmJMqeLFSxvk0NVwzopovpPs0oIO
q67FdATNbooWhUhRE7PrOIAxbZlfhGy3KIwxFnAOQMEHbOgByMmSz64j6iTybXbx
+0hOgXhof3WjK3BSWUa+/JtjCbz2XADwRKNhQ19IHCyg84WncE0UceUuuff5g5GT
4SH5UNWouuIhOGI8r9HULaFoyxjdgABR0gd8faYFCQCFzUYGDIIq7LkmUMv76QeY
fA8KwVsEH6g/SrdFYewWqK20l0VvHTPb1XnpPqLknY2ld1jTpJaEIzgXWeEli0t2
YfMVUjlApKaBpLLnL1dggJcFFOjipfe9d2yfjgsJt+lklvZUoMLC5mfCEKTcjMKH
0Wp7oIZ+w/5Sk5jvcu0ZJx6aLeQ/wsE1TwqBA6b/Q5cGT4gTBXo1uOsHqjLd5kD0
HJg9fo8SuwZwkEIB6EQILUScK0ZZodmHiuWDMhonYIWQaMElZ9FLNq7GR3It2irZ
3pmmjlpYH2ojpvj+lyT/fdguvzxZuZlKmMkRzWlhbjFLOMPqMYpkLIKQpmEy3XVs
zEhPdvegaHre4wgOXfgdRK6NpwHlWwphCKpvinL/kGDBKJb/G9Fhm97dfF/DSs7x
qYGqVbqmHrUFeVjUGtrBu5YKMM8EwKApuKZbBe7KgtTArguIxRdc4uJeL+6LMzGQ
qW8fN5JdYOX0om9LzFI0K7Mt5MoIS4sObRRvNDPhu2VF28dNasRaM5ykJvHH0klK
Hp1NQWk+SWTUSoz4yHvqDpK6ZF/VAPP73KSpas5d4uvsVDUFQVV4Z2rB6JRQaEtn
sQsKcbL0zJHpgymv40IB4kjUVbjyQWSFentcxlTkMMmRn9gFnG+R8K51ziDbcoVj
Cxf34p6rLvVHZphk8oJg6HVSH/Z7HB3fiTFBmH60cglsxcAtOxMb13q44AX8B8RC
WOKbu6bX3fwWMUgD/w4RI5rvIhls1Guwl5FQzzrNYV1zfCJ+ZEq3O8a6fq11FG7W
8yut95Rv8OnJ/KaV1i4ONx6LIPjVs0qz46alONEfPynVybSkTl1o4T2bgAbqXegT
kJjKIe1tMqvDxkEbzJXQHaZddCnD/hjLz5Ods38uzuCKb4baPjclnPcxJeYXcfxz
ldV7ER5sJ+4l6XE1ln1XRsjYrghZDDPnfwHWma5S6EPYVmVs4smJit5BwmxaD6EP
UpzYHWlYifMTq80Rfn4faqUlgEiJaqCLx20wWZRahayjqg1fD5vP8Yz2m7jppbh2
7K8BTte1g1JzBYayX+EO+E8SVhbiU21Wyej6nTueXVja0zChJLeah8y0tvRH66cU
tBY1ShvaOcqXpA3rrtszvkpz94JzCKZKwlv2riDM3++QiEWBEcdP+EM8Z7oWmwqh
KtMyzI1svagO1+aywAMzBo4k3YZ8kuOVq01fam7XeBJysfRMEb+2Sd3vlbgrBeNp
lhsFaixE4nJXbJh/JW1Xn9lSCQj7dEeugyhTaH5F7ifS2xvsNdsdkhE7JzB+lwp/
MktQe3poS2Rf5shC7W29WUeLEWdQn7rCkfeo62zt1eULau9Bm9pCG2UwnVKL+qCK
rdytyXYDHl5V6ecvemkRg8yGIpK2JojiidZl1Eda39a4fpukLtRP8eBrLDl1Tewh
Eki3+crgs27kR7K6en2Tjy3tYLMNhAzKdUtaRMYtEtPy3RWDp3FDJGQZvGwCDnYj
3gNZlUFPyVHnIEBqFh80rnf8ciA/cVgdAyLCGIZB57uOI1VFfUPxyhOVPkicCxLf
LREv+CKf0Q6yYOftDaSwfkm0E3W8KboZXzHzfyDshyyzGXISuJZ5GxiwP5TzaoJR
7K0rxnoilaArOCCuU/MRZ8tmtBwtr6yJ/PjzJr9tQ7jFeWy42SCgTNJ3v7O2RKJM
sws9diAqXwjJNErMHagC+9oedDVyOCVBDBlNV3QRCkjpcI521x9MKjuhEJ77cLbO
CuO6EHY0bJ+T4KsUqwwZFl1Adq6Z5XKeAgVehj7vEcnMtMEzMauWeAqefKCWDY6M
WQmHdm5slZo8XxesaJ6w97pl/Kgs6+Pbc/zgVR5tOhGdxMHtLzznd5ZXzj6GM2cE
iwSX1oPnPvrjeBYJugn2RzB3k4QJ69iKfd+o7bZdlHNOefKCGhiAPCl0FRloNxCq
pzQgv6Xm9adzbEkvQUZaF07XYu0YVdG6YcV5ehlBpBHDkSWna28K+GklyR5ftse7
JI9QMQkYsrKHoQERoFsueZvQfqgYXrFIUDIh8H5tDFFU418ApHSz3lD3XoovvvUU
bmZiU257AHk1g7nq3Kh+LPpDX0TzIeb2U/jWSOKoNfKtuGGPsHtHKeJ4m0pahizV
de+GuePqLxa12m6oRCxvbHT2pULnIPr4Eke28UAwBcN0ONgJ9nTS3ALU0hrRtSuw
cybTSUW7J6s9F6wUjIXPQQWRIIEkk1vXPvSui/Z/rFFahjeovgIA1FhV/BN04MD9
gx1knvGCKTY4O6J6rgvaAOlFTzXUrSghCm1DoOg6qB4Ox+qNfUO2g0Qw1pY4BA3b
C5YPca56Lf0JhshRtwLSQCJ6osWfMCj2DOFCqOKTqByApl1GpXpxxMNKU9A2JuBK
cVuuyghf95oX4j90lNKVR1Z8tLG6XidcN6abkDopdD1XA8NtpKq1BjvaLHXGoQmz
3fqQSTkKt6uUvi6j2+2v4lfv7T+C6NYwwSJfG+dphTkkeoign4c0pItucTbQS32J
lgfY0Iq4S7rwjnV3myuimTN1bi9XIXd0sRlcc6AbweuvssCET+VW0VkhkA1VYsr7
7zwnuXUm4Z210fhuy/BCgV4VFvycnRAiQaQqylB71IrFJenWCDKc0ngNz9WyAcCY
OwfCvCBjc9ou9qd2pRta4Jou9agW0bebucxim1GOTZ5qdIMhFONaSrmVi0EmZHPe
AWNXhQ5+HIe/aU6zOfSBGQJIPYaKMz1Ps007hpe7SGoSe1Xn80BNo+/N7I46fYLL
M4vXxsoQXjc8oJEVAXT44zx6uybTTM2jTSKi9qOeoHIGe8JcBb9hwrKlEK7/XBfG
yINce2Gi8+DjZAi/OY/mqvGnp+2cdCAW7YD5/Iob2bem4Zi9CtVj4tMap5Tgan7A
OjJRg11tqn2hv6FQjgv75G42tQ321TrpyCbywjcItKPJn/00tUvWyl6aYgttFifE
8B8fV3DApeDTZ2V58Ogy0yCR25elxdwqykzsbYmSnW9DlFvpH8nDH8WdpbwtUamg
m2Q7/frXvBWW6xzcOiTzxrgtixKbkuNqoHi0Z0TroeOjB2uETcINLoB2uTFOUru+
veqS+v09QdHEjmThjTc4BUHI5WofDrz5kGnBr9Nc3bPC8EJFUwn3WFZXFZ/26IPO
nQ+HM+1sl/Jg9qx4b7xOJP3GeIcZSc+BGLNSgqquMM6EnKFeRLvlyoXlPOE91Cdx
E3WFvF8vlMMxvr/hCyk6zREMQMqp0HottVIA8/yAZ84NkPy5SpDnAfS2wY1+pxJA
biEtnhKPVkaAyNi9UuwL+m7cAn9LDeA80T1h0WBNQGQpFmsLdK4gBrHn2csxLR+S
sDuE3Y3s+4cWuVHg+ohJK5tWmmkI4cuGw2ArgjT9Za3EWKwcDEt8DdAE/C+9/g1h
uRxFW0wghPrT7YJaUovZKHZ/REPFxzfqA9T4tJ/E8G1VaQKqOJuo6jPR64OgYcGC
7umL9FlzokOldz8M7h/IoUxLZY7yU6TpK8+XYsEqJ2b2t0ahh9diMARMQQe2DZyU
z95Y75M0gvEMk2nTNbImSwJUZ8aYg8OEFkYwwdaQEpU783xba5kYNQ6Pgbfbqjv3
43Hiz8jB2okLvPGQ4x8fdQodjqc8qpJWMe2DZkMUc7AYPv+gK7Pe8Bzp0oP/Xwb7
gYSlSJk20Ezmhd3FKcPQ798a4J0kwjIE8hp91LUgKlNFpxpvCLWQm+6z2GFEYEYk
t+2eMhheuBRdsrEgZNk8wxl3tmkGJoi58Ga0Y7qcNvTvcayPkq4W47TllTXL1UXo
4hXLDBeg35nTqtyBAEFM1emrsCCOsiqIf8Y9ZBlv239Gx9SmdVktzGPL/zz9xNhd
781ht5J925LvjJVZW2Roi0nrIn6yeKMSiQVkeglYG9d4PGkA/TG+IIC4mb9X678b
QY1Ou+RXbX6UeurW/6/JN7EcgF8vW7hD6dr2/pDeyNxNRzQeoKRK3iOzto6kGpMD
sAzKJtfTbpiclh43I9eBa8hKwKgKxSUCdNXhrhAa/XmI35/ffkt4yvcMIrqB7C4h
XMsxWiLp5y08bo8H3OSOn4jINw31mP+iI2s+bQj3QUZvMi7p8yz805btRNJC0m8P
aS2eLO1kIqUUBGsvXKn0V8MpJ3zI58FGjkDwBPkf8YVwD7reNoillj+oUbTSFYRz
X9HU4ktsB/lDzcW+Fyx4oBaChUlzytg9RtVhi1FIepHhL3y1kq59RZAOwYl83heG
3sSxXI7PyzE5ern5mj1ERTsYaQti+A4CJGS8iD6QUNIkM5WSguqooajwUVSykKYo
/p2l4vch2vXCYsVCgeo2WjsmSwMjZtQzQhVD1N4O2ifMcE/7bdl5rczaYTmp9IJE
GMpNnC6pBJH/UvPgU9etZq5i5NjvBeweB7pOPMIuqQVAo11iM95a0JC7eFRR/dQc
5ganbmg95LvaVnfkvL+m3VHWPEn0ISE7kAC2tFDJe5+QvvyltQpIqazIZqovkaqT
mItTav3peswrrPM2W/NDwvPzOcX8rWAoxcc8iEZGdPrSu2+1VCCtQ7H+ETZCroPe
rjkQqJhvMxIiWjGPy39fSh+PBvtGPXh6tym1b5Q3PnshxuCdwuDjKVfRBXtvafQ8
iwiGssBA5eQceNEs2OaA9QbHd+x+7797Uy0wuznyS2TNxIjiqME2H8Bx3arvftGf
O2AN34bkznkPobxlZyOGxz/4tUOF7MAh2nEED3Bt9odxtIr4DY/lSOwG2Gd59izG
9ZCQ+X2pU4jIc7kWVsJUUeW6PywpkXfFdSgibGpl2C3p6SWt95lanT80aoRBMZsN
gTUMGt+BfnKnq6D7ep5lp1phOkHR0jgCK3UDMB257ChtWk3CkH2ou/9jRUJIYg8b
Qh3/E4un0CQk/4lm6UISOWlIs4IzKUsXDr7qJBI1cmZAT0kgu3V+9lRAxLqpX02U
35mXeEYwczJNXRACRF0PsM67WxsWFBngOgSww/yWxSOVv1As1sr0uUJjtFf1sMJc
m8lMTF+4QPitMHZ9L+yEzobXy/+GW9mwkoADtyRQDO1uo/muxoplAy9awbuQEyHN
OzhxNLOF36nzuZaNOkkbXZUEFUvAgPHe91ob+hQLycHnfn+gpqS9M848peTDa7Rm
OcNVgT8fW/C1Kf9B8W25du9aAlL+Ls86OvLjpv7o2iKO8kAssRTP1nQrn+H+V3uF
ksgP6TtAjfTOQ8nSXxwXT4EnO8s3yce7LuyV75RBJ8kWcILgrCsM8uXn+5t9wOqT
0bKchrsPiT7AtprIwEVhZOMMWZ3mPduIeNy9QwyUbOMt1Bzlgsh2YZ9LmbDmofIU
pEq3D0bRietmyD2mDTz36eH5wK9p60JQr82wi1kD5CZWrB5YFEJS27CmsW0JnTot
ugcrd/ifiA6R0uaZNclLw836UtlBE+TZtsoe21rIozOe05SfAQqqQa2f2VwvejdP
HZxW9jNVzsncn4A9arm6jy5wGx0wCsWSZ9r864yK4/xBNAhf5P4KzAmdYeTAS9vV
M9/KqxMaDEEoW6iZZkchNkbpovbq4Rz+6U3EpeUl9gLgfyfeFmwhBWqHKw3ABGEz
GNOSH8hy1BF4BdMqbDmUBDxwv5AJSU9z5MXqPIiHdnViLPurie6BKPEuu1/4GgNJ
wzPRm0JYODqghJ3tql0RDDquZJ+m7cB8KFrhEePVyV3MbiNVEBm4TSYbWR7/1S4/
Nv0w06NFwlENaZXoLHj2kU7sLn99qNPsBtz64RXOL2lDXDZbrKRxsS3juBp6NRwG
dfmjZK/BxJD9w0nFTslrLbidPJOpINcjmVfQL21Y0tM+PdABE2iS2mjY5HZnvb17
q1RlKNL2jcLQIdJ1b1Ia6suKcNl2oxZ6WiiZhDvZBmKl2b6b4/nxLvbe8F6FQQ8w
tYRjZq0oPXHsriJ+n8OnzjU2nAox21W2RVjrOwEg/jkcMNWM/zPOp1nMSGDHGyHg
ffk82xSVqxN/iaJbwNuvqXSOuq2xIFlKY34KXS/piZRMWTAPAdayuet4YhWla6Y9
dWbnxRrsFIThr6uxw9llPsgrDZMm0kqczu/ORvBw/b8fT8ROwQ715bV+FYX7ufu+
4aW7wO1c7RPew9ixBvsSV2MIszO9iYsxYNI+yoszNc22WfkK0dPHgzXsqm5phc3Z
sDioPSQxTu98tmp4YIzOrDKUNb7dpDXrXVsghMGAXjiTZIlZfq4lGFudyf51BVN2
0Aw66Mv4pnyUn2GlTiIfqvNDUNQwCrHOZYSw2TC3ySZ5PRCk22jOovli3hD6jaSZ
HKBmtV5Xo57UBaL/QSc3J2xGC7zhXObVpmYLrAHCDSRIiYOb6PHnXy46fzdyJdPH
I9DBvJrHY3DxImsVT9QgkINjYF0lD1oBaqbjEgIXCTakT4V4WCFIhMXPaWeZqeev
lCQfg7M6YjLqueyqUc3LmVF1iHxr3VvY5mEcd+0zeBlqblAeZ7jc/HUMJgQLAy7I
1ONxBVGUEX1MkoQJCQGJU+B4ckdRw2jIFWZDM+TVMwvHkjx594fe1qRNmK9nQG0K
I34ZQdqh22m+ncK5TWEhM9tSlqtv9H6iAmH1gSJ0aumjxJ0iUyDWXHFm5VoPe1yZ
OEJr1TeD1Fqwyq3vu2YwYMevgU5qdIVoU6oManBY5wSNqUB9ZWi6ThDbkB31USCT
4i0FKod9FHWTyU4uavNR6MdeCa6KbHDqeByBdTfTmjeK8WrNvjCxqYhmJHIcjLe8
4Qkl6TBqJNboVC160+OHVhWqfzsyoARqGswBAa/QMc19rGae5rE33GHZky3UAv+K
wHy3dytvmJAWaAPSUfnMiByEAFzxQ88z+YOsj1szMt76f2a/gGLEqUSzNUoT63j4
QDFHmxmQ8Y2us7cfHt56ud0TjUGT48dHxXbloj3LOeRcn/n6cp+xlrAP2kFmR4jX
toxvuLFaFGthzE0WLOcCow++RJGOXgD0nKTe8iy+9mht9t22H519zjNplwDfP/JN
VoGHyKJTF/U4sTVB7dO8i0AMuf+N4jxPSoX7GYGhJ+bvoKiUbHxvoODKl38AXHaC
wP8Kk/ga6SioxlVJ5dDIUTFO/kzF9PVB78yEzua19TDOVJ8FfrPSzdThavFeMKRP
ij+O2B6LlNHqnG8RVoQLMBHop+WMlJzC3mqQPLryFad2cRbYy1X2YCy3btBF6ovu
a6IZGrZufN/DA0I/FGjd93ZD7S3pvvQMS7mnmawy/1Wxr7fp/bxYhxuh+O5QQ509
ihMkoYbYJVDS6pCHrDJ3UmWcHKzZqIagj7Zd0Ii34LPQzcsE+cz8IKMUpMVB8vOS
bazQbcDnbJL3T0jYEGy+g1VL5fW/SD48SAsXQdgPz3AroYl2sg9g+dQc4nwNCLn8
MnWSav65IZqSM92VKoRfJ+K6YWTRO6qTqGKcboXaZAsyKkFaM/SF/O4OYDfK+/A1
gFfE+sfbD6x/hH7Jv2KqBlddhS3lXrKExkrloGt9/dhpXbJ+UltS0Tb8K/Ae3xRF
igWxZMmD2TU/tMLvwYKVcfjFAvL5pMP+Y0CLa1czWBK8UGaqlrmTADRHR4MVSwK0
CIa6RPz+uasnQCDKvhT0XtYSk8PV3BtW93QozVlLx95iBCo/MU4F4EAbTH1XxuNY
oO2j0EV+oRS6oo36vrk1PY84xmTqorJW8THIGYFjLnyb34JYkyhHpW2/IvYejl7Q
vWULRXionTIrwy1ACIUihjkm/4RG7qYUuINjpGtg5ODdJzfPesv3+IZjLm+xZQoK
z1nsTmdPIDzDqZd0qQKVV4iEXHiMoFyrYHnF5tp0RuTZy7hXF760KWCSFENJg0TK
+CkjWQSkPyKZF5GnEA3/q2mtklI4RqJQ0Ubyjunui91MI5iAmLcT9cgX3rtSMrFY
qBnXmCeUsEUFvUbcqfwhtaPXITtRxC13RRNyEU/vChlQyvlqENCGuA/4UD+NltIi
UuOdtAxDTY03qdZx0e8DN2yO6uYEOT8qbe9A3AToY1TuDeCW8iAuBgnIE8y+4z11
qxsg6vNPWupDWkoEBB4qsj/ntVBcAAuIbLfFUCytR4nfsMvXf1ivk4Y/c+2t620V
j6xTDPl1p9nSm5kDdvjLY9Y2SPP+yjPU+jRLXXvAsGkKernOVVA0MfFctMgThw9Y
Oq7uVyWcZ4rTjboaNSxypJI6bPMqVYJWZ241NReNzII04rEOIuXpyt8lM2C64q11
+Ck3XJTKTUbsfJ6Yk6VFmnbb/sjjP+Yh4xOAYuZ0hlwozw69wrDgnf3Q0gAy6nE+
cGoS39NboPXpiThiTEuP4sVg5JBrZ3ZP8BL/9gG3qBVYuFLi4uixRLynpoV6RL89
Mmv8cvTGugPTf3MrJlrjqy4583ZNwLwYViS+g5vkyLXLSrT9i7Kp87HkYYDCGNtl
TEiIK7+3BSGnVKaPzDhgGqEg9ffVm19B1WAL0VNdWdfWMlIJ9ni+m9KP5Oq6lIDJ
03zKDwLoBk2NKH8JEiX5xhUrtwRa3HvaE3mN8/gT34HPSEkP3EI8iRFnYOiOt2MW
UTDv2K3gs491ATGphoswdNLq9TdOap7NqPeFQfPFXyqEkgcVEOoXG9WUBct1VT0U
lp/5TY/A+RIe9XKL3ibuxWvokD9XPrAGsCLeuESFq6TtCUuo2g9LvKfBflhRZDbR
yHfttlrbV8jPCxjR9J8UqEfLx+xthx3CLpqML5cXim/8AiXdIPQAPqjTb5W+oMl2
khTJeolj5ECXEuhQvG+raKPQ5XNt4UXlM14eZo8EBvEb8TL74ikMBlZUN9PnaMWX
QiPeNr8AgYL9LpJOmdaIP6EqXhcbACPzQ61zi690w3ZgpjCDFpApyAAXJnWMLW45
K4ONTXM3nn6QVzuq2EGuRB6foUKZoW3MqMCfs0Kjikcu5KlcMQNGP67m+64IVDZP
l9rwXEOHi9uhtfGo2SEyqkeCd0KPPWv7W2BYbv5oeGU6coFizQEVkkmOQpeI233K
kNcX6uXo6/8rknN0Ba2AkQOTg676wOVW2Y3eMaSCeksIs5fLFkBa1eKFKE8cAl+V
DhEnBFJ93w3/4oBT5kYsBhegz0omcGwa8LtkguDjKrziU0ycP+ncJlAlXPxdCojZ
6T94H3T3017BN634JMR8mEhRegdBM5x/wsVRccOgBG1QhIKUj5FpylZhvLI0E5H9
bbv2kn3P44pwQ4198CArykf2zNkoxFPv7fc9KztqKHPGppJ0zrORLLVPo2s12OPu
qu+9OW1WJUePuEDiGkYBNAcCUtq8LsKNpBkxZWbOqWYye8O8g97HB6bJ5XxNsNWL
Kx12XWnDNNfcWdzfwTP64vyXdTa1ZtWqfelBmktfpkL59c/SismIeg8/aWCyXYx/
XWZkguBKkOKNkLG+YjcAc6T9w3KXFjHCbSNwhKM29LXJCCj6jjSGVgAbBb8pyo3h
qwbPrh2iIulroDk/8zHl2pE93hHms6krCZXOOc6w3H9HlwYX1/e/Ws5RkAsV/CUK
QIniSQJY1IR1IpwiWxHM1A6MnE+zsGKYHQUey6wNma7nZruFvu0TBNyLzfsOTgcG
MONDTPeGnpBfmvLsPJxugn2y5j3QONWsEIF71Fw/6UYCx4VC2l2qVbTOY5wBPtaC
2/VnFEt69Z6QjuSUnSQNuTzeJjEna29Yc3vvR5bTaNJgyPyrz7AGGbuQWLmJxG5Z
+ispPt+bDxfWFURrrUsrClHBZFPU3Tr5YiiFO4+LcFnRdYj66rmH8bUPZANmlewy
KjuOezYPeLMzBKkVUkvPSgbT2Dy3DPkXkysQZmdOelGF6l9kyaYId+nHhubVV6KI
D9CjUAWTGd5mUU+bzH2D0jvTBFgLEBBWvL4cV8z1huniJH0oZkvbKLutIMMHEzb1
dhVAEW6ukkUukg5t3uPVnfhfMyaJHtgRcBZJV/nqI0RKpnAZ+fLVFTOR5WAzWOru
8I+e64wY6VrTq8VkR/WoS5X+h0t04/PaLwY/SQuhNLgBUgLU6PAs/L4wTza1i5dG
4i0ECeqoQ7Kd72ZuZ7taEULXjx80GTSKF/u+VsJ2DlUxBEUBAjkkmbSEaeqwOVUs
zqAldVtSICDtWp0AyrBEtUJLQLanzFb0Zbwi6GdZmhsCJGAXnO5utG1WTYMluHih
cBvJ5HsAIorlRPYvkun16iy2eQBwpe5pXA0UgYJoF0rLuG8sIPzlWmmmTsWX+7As
FlH89QUo9H9LPYbGRsYHJ1IeX88ZM7wozbQYDNCeihTusfgXr9UsDgM3Z9Zdfb+G
MgOSqtKGY2M4LSYvosy0WoL1TnTtj3yNRtKzAOkzU1QLAWnvtpR3/UPqnplMiDGm
YAA4McJ/xrbgQx9nX7f0DdIuOJpkCDmC7Na3VsFbrX55U2tzkVYkDMidOURfWo6f
eUAHxP9vFGZUBML3HSFzxs7LtB/qq/XLwAgI1++fcMnqy9uJOSjKJfkbje9vL113
SLBtsIKGkODFO9VzK868F7Vp/o3yXru4Wi0sU7xyDXuHJI4rbjOsDIW+YVpgCYaK
z42D9qdCrGJEK2ACBq7vtW6IvUcrRMWGgvpZpv9iW2gYWVba2qu0mT7YydoBrtyD
5wIjtjZ3gzhHiI75F38r8rAvTHP3kU2/W2EI5alC+ve+f/pIOONeYAgBIR62C7Yf
xOuHQKS/w7uw5hQ39yMwP9BBRkTrfIIVZWNuN4xOwY/07Qre2FdcLrKNU+rlz5Gg
j6AG7sXjeVKqouqEfOx72De6DRpMJ2LwG0NfxEGKnfuODxGyUYJfBFlwuYEq6dSr
BXN00BFBVQxvtTXZjPwyKYMO32gu6xodIYwEBretPs8y1cZNvywhL78Ibk211eXo
nuASyjE6cv9CylT5UzL+6ZJ95vvUy+q1PAnYsGqFw9MDBs+yKJxzQnFJcN4nDDPu
c/Dq3LhMyfIh32aau1VIr2xZAgsjEoHqG1fsfDx+F3OdZ88HMhseMroqF36s4f54
Oa2Z6sDrRNK0EuGjQ71fwu82xuYZcUHEK/6MkB5tQwQXRvGTEntSjPHUUZP7DVSh
bsVI7uXlRUh9IhT7uo00Cy3dnIxl9BpQtQlcdmKS9Uc+x9xI+7cuIDdsDdKFYl5l
if6NsmTq8Towe8bD4cVU0CNvSRiLJqOmjbGNzaB0+1P8eILoQ+Vo0IwHz/IL+5r6
PG9rZv1N0kudTnyscDV93TWdo3AkX/hT3sGIYWeKdZaTfd0fzHKNStcVrwDBJ+mI
4jX1BmrmUovohbFRHXFLyMcUceRwVw8QurUffvytufbVVozLQY67+tKbpgX6/qOH
HlSqNbI5LxS/0EHBfGjEDmo4YtdRjEMpKQI6oiR7RsffpKorAD570tqjSd+R7iPf
XFPMZAWB79w/DiU+hgC4hj5DEF3rCkelgh7BUlTBeM1l1/Hgn57MxoxmzHU1chzb
4L0d8pNnKwNBtwPJy0vvPTcPzm0EqPkOPL2B6/+76UclD63v5ty48FtIX16cVJmV
Sf9kt3GVWGoikdHkmuRQD1Dw7QnqovZ7s+wDAngMcdpDarUSUS7t4m5yJ2fsmb3t
1Y9Z3s9R/hF7LoVf2ejZs1D146lV2voPIpYm3dHwENmpg6LvpbTPQyRf1inK6xvn
s0zJX5exuYUlwfD6hod+emyJboEudAtu1RjwAWub00yoDNPGMcvZwaTpOlThr1fE
g3h8JiIWHE8cWKb0NSCVOniLJY4GkqNtmK438xngegEH736L6WprBsBLjGfY0Jda
eCveA0bYddSZU9KwARbhyj8W5yG4d++5xXz62LDJx9fP+cRNVv1GDdVX6P78GBP/
B8HNPCLLZNPQoF9/6AM46WyXI0OuPVH9SxPK0qFKhQkP/3TbC/dKYT5ApEAnDGpL
ZL4atY5ZfaJ2cuM0Xl/eGR6gj9itpjeQWNShFevtqRjdjifkygljRb2h2IUU6gkP
0iSmwfJq064UyaK6NO8MDzlbChK2cd6TuJz2VHQd5E7aaoOtIWzFy86FYvFrK0Us
`protect END_PROTECTED
