`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6wU000R025eJyYUSMdBu53sZuHx2KzC1luGhnyMdRrUE4vq6ZgpNEcAhWOCi2jtn
TUHToUbbCSJ4UjMWcXqzXs9NqcYZ7Dk+6SGh9potTTJH3Qea62coA0dxHBH7rTiU
F2Hmb2cRenL+UQRRKNFAZrOmERGLtvhGA1MQp24JzW+818Hp1Xi7ZbM3RrB3Z33V
GUHru6oMs+io7zo353tz2I21jbGsRx9IEgU/NnBVfvDc2XCbSaMoGTx5YvCPSWaX
/jZUnGaTQr0elIY7NTb3LVIx2HpZnM3bk/b6lLGfQejz5MNa0kjgjds/FeGcZsIg
PTmueW0j/hnMm6ULq3qTHn34f9/hQEWfBnicwZGdwMIJS1pWeNvkgw7YLy7z/UKh
o00hYntFrGB6/347BR/pPIUr8SpvGHsLHrbYwLz8VeaVCoff1ZdO8mn6KpXo/T7+
Vbbqlqmou5Vd/WNuz824UEhS9AlFLL/2UemUleonlPztmVzCT1J7/XBr0hTM+LdY
J/Zgt6hm7Fgm+3uRO1+dmFztMpUDCCANBu8sri47rwz7xzjcAIGjNzF/YQObK1zo
eXf/hp8dIZeF9uxc9IEF35dCSYjwdUxCJpyWBnFwzX36dXTyImP1vFGdWqXURte9
De5S2sQyv4bkZOjJNAjPCZO9REC5IEdZopw6Hmp3s3b8bb+f5LHXCrL7+wmU5r9J
2TJxhSFUM++ANn6zWwxsJ175afwW5b8xxjExptBLm4xMEif4axSBvfoOVbEnMSst
1zxP9y/5p417K5IVovU56j8GRK7aSEthTs0kn47XsS34E2fwcYEWHzFdl5Jv31xs
yQTIjEzbIsM4OHG5bjIC2IiZv0zup1U3efzYmyVrqBSjkc8s7Nr7M9arIaMVUBJQ
vnSiiRmz0py1PsvtjImAYQ==
`protect END_PROTECTED
