`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hXnYYtV8qsGJLpaMubjqBDyGGlPSwI0HqMpR6UW2BV63U9VHFhWq7k8oFkDCACb3
ZbIdjxj4UO7/J5Jfxi/fDVy6ote8nnqFG5/pyoEpfDXyYEnA1sycYHMaHrYQGrMs
NknbL8N9mRmrZ120LtzAtvfdEfHqFA/cRO7ARKlyCq2SnciLZbecQ/zUMglT0Phu
2Coa7IpD0ZjkmQk/bHY7AJDUmYhSRTDDxVeI116W4HL3O+VySZWfTDR0qeKLTT+A
jwPwCt0ahg1Jw9F3xg10fizryOdQdMuiWN0XLYHdr3R0Gu29Mg1HJ2Vpk7S4LRnQ
tgTFg0zg4winB57Cpzo8uq1G1lndxgdT6nJpKiIvR/2z0uBk/lUcNikLMYnQEB8R
AZbv+9JDE9pj8+y/9UFgQLigQDJcPm559QgTDODxEnrm5z0YgaFS6Ztsh2WaLfS4
omt1VWEP+fjL11OCDk9LZM1kFSbqGQOEyTZbDYcZDA/aKaREh9EtVENIYx/+acHc
Dn4IADQIsM8zrfU4uF7dsqyb30hOfACMzNljO31BYzXlX3gwx9aPc2HjiQQMTe9T
HTUaS/zxs2T5qxxHMmDGt4h6xZ0pveWxsSViS/RGcKpr954zn5ztquzbfBGqaWxO
0U/m+M6OGIm+jMLnt8CpZmkKY1GLIOrp/kMTmi78ihzs24zXLLk9VHdN6G0ujoox
yISBUo1Gp5fkQpWBnKSoltbyBAjcnLI3bENGy/ZZ1g9FoPd4cdAVfeIDzPxDZfGf
2EueDPoy/PJsGXG/ZAXWr/ITGqtoLdtPIm1y2HWB1TjIpI91lp7ETKympB3BZfxC
`protect END_PROTECTED
