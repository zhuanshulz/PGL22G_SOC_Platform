`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TjUlBOXbrFSG/1hX4duwdqil5fctwApYQItveBghGDlSuYz1DIOlquNe5yRV63Ae
UzfgSUBkp4SNwj03BaI+dozfeh/rhZ4Wz/U3942waH/GdWstUoJ4nZ04QR/DGDlD
jwZ50vdsaviyIG7UUBlajtmh+ND2y7I51E13gXsUUS3lUjzLF4Si16gTpWooFEjy
4aBcA5DTwFTmKkU33Q6ll3B43JPNFniZhMNdXaMZ9Lgr1oDZ2PxWBJoaAelE1RFQ
RoFhNT20etl0JQZyN19KD52oD7Ke4t6Xu33PKzmnkhLzxBDON2maEOfvpxdPYKBE
1uWHNTG8qosi2VLyJcetFYS2PU1JXxFwnBYiZ3mwU1af7m5vW1lZP+PZ2e6GlHhM
tBn8WXJqnnIWTCH+ICA96LNIsKu41nrAzFIHkWza+VAp/sLzksXd4svDAIuMwcps
rs06XaYaVw3CXdxDWRPB/A==
`protect END_PROTECTED
