`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ddd55sLJ9SNtHY88ubUD/lP0Fy/A02MBmSwbJYs4UnMh0hbn+wgAqKcfshEqSLXl
LwENMwzmPLc64yWLG9t37n+BEpbs8HMy20NJiJRiJyKP4sjNGvv9GMWZUFD3PwXW
r2N/mHa6n3UPr8vtTGeYjrMcXm6EIXf5m/KrfyzxEku55Jw3/sNQEfh41zGT18gg
9FIxZ9NnupzqCSXeS1cL8wfYdsKf9L8euAFi15yj/QcjdK8xqc9UNMsZXCUd6PxZ
sA1T7qp9imFtVPtIdqw2CK9g4VFyYm7FTFbAHjqPu4S4fHk1rh0LOBoH/yCw0Vfb
qnet+pHCBqq5dTtL7tsRt0ALiaTby5BzDi8l+HUGqpgdyaNkDVaKQy2UIxD/zEQb
A8LfKQuy3GGh8VY8vlEvMw+QBZAkMdLhsN25v6UndEtXNlHIy0ncywEwcimA2TmS
tdrJpjLDuPdVp4QhfK1WjDalKxpCN+CYwGLeDW931dwPp6MrYUHPcJLLqRWKEAmm
oEcOzQaRUU4S5V3X5mApxXOQeD6GjtCI+fLGkuuKVMJpgd2qrrFuQHC9XcOphyyz
/JeT5rKG04lgnSBBdieVWXPNj6QYEQeAdTbuqj0XDqPflkWKo7Z0OLb6qnrJEClo
dWGtMN3ycA3MArsks50i/G+qgLVy2Htv5MCvzMlp+1CSQBJWLJ8N8CO3Ly9UhKZB
Du6Scc3PgyyVh978fGIC5QHO6GwDUCgr6im/RJyR5iU7ZS2XKhdMuJQYtUtom0XM
gK5s6gtb1O6uMm402lx5N4M5+KhW8Hx+HWo06oAOFIKFXnL+W5d9ZtVzQAfJ+diX
Zzkin16jMafkiOnfExyMtf8ds1NkhDzH8EqHfFsho3gHBhr1wIitGHdJBmVsZj6J
fc2AqjjY6p5XYi2Ncf+xXoCI0pQHYomwlaEGT/kJ0Lg7KoXR7++pzI1EeqMTsWCG
Wa3kYtFUz0xLPuRTz2O3cz40GSJtV4V24ecc3vSdek9gc/O+UBNwj9WQBBPs6UC2
atZUDOvux3wUFJIX9lKlYPDYnX5jISq6swbijBrMV5TpsGK4YNtjidlanJgWpzkK
UK8c58JN0w/8mrsWZdAS/Pi9HmGvYgIxJS9yR/r7lqdODyiBybmPw/LtUL1oY1xH
zWGYNxJV3TDiGC9g+fo/EG6QR79RZDUY1pQ+LanSAmtee2ybLStTyIcuScKDaRok
`protect END_PROTECTED
