`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8K8uvSKaVIzvsstV6NymYQtI5BxFKDreae79M+/C1GJp5NcvPn3QlwFx55Z6RLOi
8tqeUwIFCyN5U1w1bgIXYPSrKepjMnztEADY4boAkfTYHL5v8L+BWbsQpc1gae6o
Kh/Xr+be9HPrjioGxdGiQUpBZd+jFiol8GpleYwAqFFauBfJiNlzkfcaQUT1CPAW
yFD5Vlg1bey/yp9TMy0o1JmYcZwYTd8mEJ5Q4IkKNWQoQ1LLGU0fbciE4+o79zyi
0BCgE8Sref3GGqzrn2llONvsjB8rNTMYGCa1Jt1JDyYRQn/LWhPuCvsgBBHOMvCm
ALGmRRA/c33pPpRpsxZEOT9WJvysQjzxvU0EL2VVnb8vboZN4kzwhPC7Cab+xsEC
iXHJuvkJF2xawRrZN+pOKGDjkEu9Z9G7Mk2RwMJS7T+i5HehFDlPJB0rLlNrVpHM
u0tmiYysB1j/009RgJU5DuCsl9QO6sS7k11AVfjN4KkpzXrk/rnnziDlso+1pPj/
VBzkyD2tdpkHeBMlv57mVwupUTjZiWgzbgm0QJvBwgxm3OyOS+CVhVhA65vMLogx
kboeYhCYx1OBZfQmcFH5UyHfgSz2PpVqCZgLzXjAH2a3c224JMmzQbxwY8nrsPH+
YzA2RA18sI3qBbIw0T17BPLsyxDio3uNOUmCYAYJlbNqCyOL1R8QvtPUZNMnrheq
QQ8UD5Afpwvdn0VYMnzQE17zFk9JPQGSk7hCEZMUDlEMOnL+1pSqbFB7ld9xZ+JD
UDaO+fS91DmtQIhjs2CSGpgkKikv1MPx5ypxLU+4EUT7Fihy9yJ7Yh6G13TrD8aX
cCNQU1Fc+/lhKlviSm5vLRcugj1k6Q+RknhAq/qvvgf6o1VRKf4VmVVErpX1Igzi
1dwdl63MWTACjniKKsf/rPcd0z0rkbBJeXI/BDWd3xM=
`protect END_PROTECTED
