`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ek2pYbMXHJ9BWAeMIMUsnbTDCNN+rdgFCeG4wcgPg7SI7PpYlvzdxAF5PF5vjN/F
EJEAtNLsmtpuYS/jPrIBJqfRPgz277CfZsiyfuW3e9RAG6b9WRdD8Ee+AVKIVTXq
CLlMN1NQqHT5YK7998G5C928z9995RKgkODcTa4zg8pDyTLxcAYay2gPd/KklYPf
pRuFHM62cVwmkZRgH8OZiGpBP4IYuT9Xs/85mpnv4I0os8eg5JOc1SPw4u/5+fOL
P+Afej2MJP4UFusM4r965dqARjKr0nTFe7cZyFC5VBLUFdRoG3NGLXp7WS84HWFH
b+v7DstWuirga/tIWw7jCocZyNWtCa6cLok9gd1K3XTanfcRd3aMFdt/dPG8Hbr0
3FZpA9CUgzG27EHIi6JSByNf4R8SKrhTFBhi+6HHdI0=
`protect END_PROTECTED
