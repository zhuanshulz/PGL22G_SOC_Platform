`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kErkJBd8cIDUGe0hPnPUkAkY0IPVPgNTEVTBrlj2OzTK8/xUIigBvy7Hw2qbvsRa
eqCEwXedB8g+FSWRXLWChUzLyC+DOwgUHhKTvVIQIOlzSiWdR8wdbV7lkRZESb7O
N4ZqXhxMg9CLKBrHc6x9SBPHKWbFd+UWpraakOu7suK7wXrZ6EwgRMZ71cK7XQXU
zaVsuXZL4bJJ1NAc1ET4GQtC/YdbH0qqR0uPgoB4cSDL+65VrFgFF6eMMjyifqV9
2Pv+3MIcAVzh2EaTNlWA5g==
`protect END_PROTECTED
