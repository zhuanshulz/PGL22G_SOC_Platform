`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
unJMfpWh7UY58nDOrm+9AttRwb0Vv/pDDOgkygudoS184+YtUzPPO/Ko4FuMg8XD
X6ufLLWHK4zeo5QwUEvX8GTPwN1yI5/snA77flKPuiZ3r9iaF0vB1TJg+R8DE3Ce
K5hjeEfgj9VBFTTNjzW0Irp59WyTwe1Y8hkqY0Q0SadRKJh2Uj2OCezMTGQF7fwA
uZtuFUEDvS56Lf51VYWgs81YRlZnp/fWh5Pq1ubGzfan8L32d7/OBOb1BHNg6lD1
CS+f8bEaDQb41OViOYGLdHPa1b4B6T6YYp/SRla1TFV/ydvhdPOVFVeKRFDOxEyR
ikl3AEw5UD/bHDNWHDpx+hjIj+Najcu27kPN00DVSoIDkrY7xS2MlHbQUn2gUC7C
ZBiDmcC/xxJIHHkw6AGrlih/o2nw+zflG7w30pvA7TD9+KvmuDqEzHiq7/i/ijQd
u8YJ2UUgD5iYwHGRMFVt52J9dRoomgm0CDWaUMHTBu6HtdjVWm7QpSa4Frm5fDAY
2XICoSuo3xGz3u4MbC9QUtnOLAXX61a8w0Oft1PKBStpfspwmlpiIKQLvTsomdEH
z52ioglf5W+QMIzeerpHRSaJvAGLFyQ8XpyiPJnmyac/a7vuL5oTSyx5cbWOaJI1
/r6Ne7xWI6bAjrp92iE2trp464uRziDbNqbgjL7u3crNHowQv/3w1p8Ai3hzS4M6
kbLm3xeW8hA1kUov5hQTQlf7Qg3sB9r+z29/R+ngxO8yZ17vDMVJF8dZsdZA7PYm
JmJ+BV7fIlBltr40nlRJ8J+HKZFF3vx46lCJnQ4LIRA+Bq7EEQZ2mu1rFaGRokMF
`protect END_PROTECTED
