`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MkBJ7wfLd7DVtZDDQCvBpvUSw22VpT5TbHLO8hSY2UomS1GayXwqR4eFKoPYOibY
W6HVEzo4zjXgvIBWOtCtBGEVb8WTydMnby3ApfBY62FtC45RTopDaNP91nOq0S0Y
Gop3F0rsJR2fVyYt5Hj387COqQc54DMceLpZ2qjdPdKvICI/ZYKm7ZChet5R1I+b
iw6n+wGolsN6wOeyXDiyqbLEdh9SbYaGjuJ5v6wrV0gig6fdOOCCODxkOL0wxdrD
cdSQZJJDvoM05LmHLyx+Oq/QhvPpkBe8z7tFxTYK1zY70zUQCz2yOX5+TxLsz/Ed
JH+AROyaCWypIWn/ICLoQq+lUDS5IAMltNLNuJ2ZEA2hnQha4UmcSwWVebSdGOkv
GsSPuj8w41SUDTUt1lS1EoclIEzZsCdbItGG/QKPpZ7P8QtGXyunWZfhJFAYIAgZ
6gdNo2qcoou2jp9No1UcQ52Qr+XruumX2IKpISn9F1h49IHkf2xS/ZTW/4JQshTP
NSi2D+LQW5GkvHhwkzB/66Ws7H8+8PmK5kbaQHYstdd3FbRfghlRACdIVOGHeo3J
E3URcLyhzxIS1HjFis+sAdQ6Y8HjluX/9M4kY/npRldQA1FYf53sEFbRVu2/sGjv
+S+AK28bT8OUi94cH5yi+rjixGIlEFj6EyhQJ/IySdltDL2rC9GgS9zHZiVdCpCu
IkVmOAnUQUQFuhcEpmfdIYh+aWcBh06/vr9P5fJ9lF6grHnLCjrUmzNHsj82ZPch
n/lES0Pthqa6chYG1DLM81HXYMXgBL0onXMSWv47TWi3CpULdY2WgFRGKMLJWvQS
LM9oB/lmCrLpNdQxxNKqP9aIy+cBskZ1f7lnG52NGX4=
`protect END_PROTECTED
