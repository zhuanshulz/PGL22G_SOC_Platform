`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pk0V14FlEjtlibv3Sq6KnQ6sLyJNgxgSeeSPLt+U/eF5gLVwkpa0lo9gbv5Lz/rn
wY1GGDHjSbmHxlZ2qmhExwBshe0vKvBDeQuB9BkQe8M5zGQJMBO1lhvAfXvoeD7h
d6uSTZQFH5AvzI92BUofL+BCdurMO7eIQ2K447fDyNArSgtpozzqI4LtZ/QULRPS
ogPHxr4T6DHyvULx6tQiRG1IC+nAO/lLUe2em2tj94gVH2knWuWcXbudBPT3mC1D
tpb0ndmHZOsLGV5y0TwayU9cDb5tB0/pyS0YxoINRW0pTE2eSf0l9yDq7OZpnUM+
gDyqyoEktvfxfcCYRhpk61kR882x4GcMJVD+Ok2DofNWAS8/mREPBEG1YoMRHT/3
0k5jfv6ZWt+2DaX5iUJq6wdeUXKFCchQxKRsO+zPiKR9dxLZiRpb/zYYwuAe00bD
FZZa0Ppt9XZ+4voOnWdXxXaRlNVQ3twazRlX1lQ2iTbXyQ3Apglgi3Plq1N0E9kj
qqJsFYJ3pCbwuJjjYwXrkjJpBeWyjqhGTLoy3j+Stqt/mS6OPrPall2CHhcem0FB
sdtT1gw9UH5BrM1jg7hpkOJurWEltlmIbX9IQUnvrd3bhowQHhjval8bL4QMR0RZ
cyRe7vvSSmIW2EaMbclC0JJB6cSDxX44MKlDYxyFnfKxP+guHHlIH1BM3m6HUhQl
DS9+iVMVMGnrT6WSirGMpFl39f48zKSXGiCTp4/pXGtnvC9Crteym3XIxF6iTfc2
t8aEAtvomUaYNCguXFaFdg==
`protect END_PROTECTED
