`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Dppi22+BAy58XX+VqV1tAcUqBkfjr6mY1CRfJizDss7qTNtk4HsmcCo8CjSRZIEQ
ZAzHLghUFUy3L1nReK4RISs9ozhcGM+8R1YfhYYM52EXyR/N21ww9tCJL4wQdL5t
yREQXn2JUIrKk2gQcNjw+yVzAsy19QlQgFtWSG1EqhcrHwuKMnowFCDTR/VXp7yc
BkiUoLYJN6YYOCW0N8DvVFxRd6KsSoClIxBBGRA/rS9W8YxRbfrmU6KoczsXYBt/
utUN6kA1tBtIi21oBHh3MOVHeZKdOb2rKmWz1M25n1GFuNJ99yNDebXrkwx8IuHo
JUvAF/A7nCEKhTrxbP8YL8QLPWLUDd76fvufGgJMiZjJz2JanHXOEee9auSo9Mcc
iH9x2DXQ2/5dIC8e0HpMPVqg7tW+W7LSZFcANnjwZc59WubaRWcQ0ct9OEO+2OUs
4OE37E453IlnzzM3qB9KcwF/wtSax797SJZ2pxe2AqA57etfjCjK+DOuiUeO/3/w
n37snZNor58Nn1pJ3nLj5HbqVtr/AeHNBp48qLZNB+vLb6NX43a98BSSc9ggwfcO
43SS8tLKZkemlRRy7QaGfR9vEazoUyO7H2AnEc8zYYFZ84U7jdagIk+Gr2AM7QXF
86BnSo9nUPmRCWm6NVICsUeDtLATUMZ8FDhiIL8bkpzx7ahJCihYBEQBGri38u+0
yvohNsFeLB9tK8Arx0kJWXVIfwCndqVNLRs5A8svO2j0OpSQ4qRrHElw/EsEJEKI
gIUoCQA6AVPtpZ+EAMLm7s4rjoVBzteBC2NEopZYGRwiFDTC/Kd3nhy9EQSafynJ
LaGgKyZ4vwHA08IB7iHDEAbxylVFGHU4UgFF1+KROhIsKxMZALamgYLqlD8si2+J
`protect END_PROTECTED
