`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mYjfmDrz2fYyhSquHR01obqMOBNffmmWmJ/vNju/BAPd+0J3HY2jcCA+WNdTegqX
d1TbIIVPMTkSvQIvqASF5Fp+gAcaVkz/jqsJW/h5eYL81ntSHBOiSHq0ytIeaFaG
xVX84ZBbhsX9ETIHA2nGaoUfnB+rCl3SKx/FyWLFlnKyPOSLvxDAAzKz2LIi//6H
MMXAPHeO2cJXGIGLllQDeD2agqZSfJyjuYuHRZRLppclO5lk3/dFybjl4GrNMogg
v/Cj5iEis5imCdRV3ageO35CplvzL0YZEk1eETTld+aSUO/su1C1z3QN3O/ZA0Do
S4c7p8yIZFLpKjJFFWi070cmEWDtzxla9Qbry/vNRXk9wp8Gzoh3t4VZ/fHjNT1X
AAv6HA5YWgNMP8gQCb0WPqcu1IM6bxb7QST6BQJ9sqvXka9AJRfk683XZv2vKhB0
zI3lHZzaH1oew1q15ac0kaW8q5A7BVbo31Z0u20ILM7GmU30ONqZEEFu6+f9rahs
3c+jMeR+aVTWHwloU3FSCEe5viWzLl1FkDGdEzAd33Qzs4DiP/5j+UnkKIQGfBo1
lwH+xiNytaWDnztnGMHCO9E9MVZIMjIkyuLN4BlhrrXWqW6PPwygU9lVlrt4b6YN
e+jG/ijbxkY87AAX8ob7HnXELGG2UQuUvBdMzVkogSmYgRg9fU/9uN208B/f4FbE
iEkBsNa0s8eASaRtNnngnJZxvtW/q0OzXztn0ylg+GCpa8z4P9+oxTKOLVI9FKkd
VBC5EQlJ5nV+e68c++JI6bO0z0lRAD0vj1yq9XmV6/wmAKI0LFsGMlNVLJoxhCWB
6Rw1brMPGqjEV2zXFHCvV1is6P17fXJClqG2cdABMtE5Y+85XzOZnpBSNK11ZYXT
bg27kMmNCp4PjacgoAfs+PdL4Wwu/NAFunuKKTl6n+F/xM5mir4twj5lf26wsGga
uOz591Yu7xjSN9SMtL+Bpt2LZ43Zl5xygNCnj9WI+RjvNb/7MyVwFoLKM6EAT1//
jbCsekTtGFK9uvvmYzmq1kiGdRWpRBgDgbrGxdM2Zf2W6aC8+lMcPhkIexoqnBtr
dH2d0YcO17grDemEpRFCE5PaiVYjPL7+VTQKGWJmT8uHgbfUGPVkQ+damRA0EwoH
ASfgAkwo0EhM5tpH5H8EtHylow7GdGriCwYpEbJXPw+iM7eQ08uU0hI9eRRhwbjd
synYna/tdUuf3gANDoMUrg==
`protect END_PROTECTED
