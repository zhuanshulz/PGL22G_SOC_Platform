`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
051O248NfkFgay/zp3nkFpgGtQlQqWFtwu9Dm0F6mfmSi0BBiKCmRrDox1N2F6Y1
8lGxKuutTgoSFHeSblIBTuOJlWB5rFHkcqPpZVjzFPa11UgLUTq/IJ1+NdzbZGa+
OeLQdgkwPANoVLFK/hlILFXDlgygn4LG4GMAg0LSatUZPCe2XYNdrSglIeiJdYpn
kkN8NAK79bMLyKAQsFwEbkUtH2vCVPjKfuA2KH6Z5SHYISPSuOEjKPJt22fc5EN6
C9wKXrvhfR4IU+C2FZPH0mEd6dnlVlnHCO+ZzZAf8P7mnVHdQ9z+7fc2JVBrg2Mn
ASGIIQTq/hYoiZn2GUupcpDdfFx24Q35cT9/eht8RIntp1nFuIMdFUrLAjocQucB
K0ohsdJLk6GPbcgxCl6pCj9gz65Lurc+cz3uKoYdpsE+0aCO+Vfm1gEK4raVLiwQ
/mkIUHNDpMjLV0OlloJ3oYqKUV7vibFqQtUyPjLSLlATfoGL9kOk67pu9FPx0HHx
lI8XBmCiyM31qvB1fgdVhrju+m/xP1HKvDO5qiqsYd+jgVcs0xK/r+DfBNv6es5N
ExZhXFnKR2vX58CrmzUDsw6E9hnm99i5tHRwU/5+3bU9ajr2aO9wogE0IvQMNgCR
ph9r8A+RhdyIGW9i60UtOl9woVPUHR5aT0Y1M7fg6YIJ5Yp8FJ20Z7qBOPXHEM6G
J2XwxJOV2MNRAjWGFOtmG3QCTS6T+iqgX18DfNTqf24F4FHd0b9JEy6U9KS1Kpch
Jc5tGjHgWoTzoat+BWSGw8TeZEkH9l5v6ACBF49tttgpbygclJgKqXpY4S3oIGbj
T6qUjuVcdTL/D/8IijiLVLV9tvsdu6w2JXzEoAMT2TNZnxwE6MJq1cwevvUrH3LB
2eNwYa88NzQFLBIM9MrMW6L66u0tjyuEZ9ZaP+SAjbxMLlAUN9iE+FsYq/HNkOGk
n47yiRHPf7Sxtd8RXVKvzqEKEHJ2/IUy6RmjyRHoDvaYQ0gTRZw6wQXaJBTMGk2f
aqnaPO4N0K6AUtvKOrvzid5pJ1nAqpwrN9ofmouM8JTc4iOM6eT+dH1LFFT2noz2
vRz0an0wKvx1MSK1p6Bx4WIVwisiJHiB5JZrBZ7eG9ZRE8LRJWG/1F7ax6Ma4AkB
TyAFBZMQhgF/Ly97LSOblTnQ4YPdOloDZ7h/e4RAnQ1ztcgKLEp9yvl05/Nv1LK9
cRyN68d5rW7+dNpyCo750SMP3neUqgjca2PzJzQLf8DViJXAdHchXnlB9jQcdcV/
yq6s2JnqR3p910tCKrq5sz1gMsQKV7lSUj+oOusO1819msnsvprn/+kbyeSsrHVO
OPaRcb8iLgEC+d1MCMOmVVHBi022Z+sKgcqlkjzR6bA6WpW+wmqNBDYP7/dMTBT+
dP2peZBXrim10DH9W9BknK1rTinaU++pjhycfuWW3qfWgTkeekRQ8JkdUs7Rfbjq
qj6ZHITWwHHjyaJBgVpXPXh4YIeA3hpjnv3JFEED2gnVhyPDtifPaftnCLI2jHaY
kCCGwCqSePTnBFzCmtjN+msBm1b4ttgsDhYtHyLVoSzAv2IIeZt5/R/Zd7D+099l
TJHQ5RdxF27hUnfhujBatnN/a5qghS7LDD1LgqnrBwkIcvax9D4bp8ODKhYvTT/8
DlECdu4e78qsIJXXaoMg+fXi7q2WOGS8j6esMm8dE5yFz8whHBI4qhJ5d5zUzu8b
tK4DqhCE2xWguIzfWIRluXyVKjTgRFbbdBswxUbc/0dwFVtAHXVufHobxwLXkrb3
xN9ciYGZN1HEZlzUnxLHuKPTXTZsBMNdz7r4ji49fGxo0f1A4ip0+Lib9WgEqXpo
huN12TZK38nWPQl1i+4knhDDsJZTqbYeJMaIQaMwYTzh6fnh3gwnJwJ4uQRcZ5UD
iRrbIEcWTGyCdiGS8UW6mhQVij9mXwAfzkhSy998xXfCluedN+34K+IOKLXGkzWi
QJ71a6XX1MMEZ1tU6MfasCjg5qsRq5MXf1uX7aAFDVuBPl9jg4MUjdIH8gI7oVgQ
shvEMruqTgQg3qnUw8ubjuYvieVUpohwTR5qKwindzsvbHS6VLWiyQFHYdwRhLrJ
fo0PqYpNPoicHlK0Oj9pQbRyaBMmOPAMljGvbdBGnJkMSpcrp2dqrIkwwm1NBlWS
XX9AsBfpU6Emljk9sbSInTSkZeW4WnZF0Z0WNSDRTz3JQxeHEnakqqSvm0JFmHyK
+0TyFeqf5qPdwRnLl21unmcypkKeoQ7zINFSqK6dVN7xJiTwVURSkRokpliHketM
s/eCjVRS9MjBy8mjjwilfb30CWu8R/HL+oAuNqL8pX9bD5w3R1KGRXAqpavpHPPu
48O88d6s2GoBBpJJ1m4o7w+XTADoC8n56IutANtlYLKnnLAIQ+YTJS1YxGCcfIvc
vVgq+o8CU4iz4IDubWTbExt7KdeQ58pboHC6XH8YgNYQa8CBL4MEcCMqzaUX121S
3UStkeL4nzu2qEo8q/CKHO9iPt37myRzQ+X0GGtSs6CNdsBf46iIYPGG2y04L/Uu
NkGIOyzmfJYooZ1yxj6JUBWXm9VnKEkuTmTKawoEfcDU04T7cWHHjkEBOCeYwGCU
JyoHRgY1/HsJkTVM1qBOgkFxKXsnwhBhWrzt5vwJVcqUeq/PEH0/h9pQbP1WMRxP
st58h2mkG/Lqy3zU1H7oOXt0+YSINn3scz30qXbbBbqhiQaR46TV4449rQX3C3zI
cXol7AHQEzqGTcIuu/mRZSqsgwe2ofuECV55Ec20142G0w8330MPsWORoJpTvSKb
S9wq4hZqMq5lAaWvlPU1+otUwOujsMqfBDxgY7BgMqxPMucM1z0cKJ9CfUOHoOpX
RjZ4wlsjZH3UhIqN1woLfbESFUFigbXFtAthouBbGtgLje9Ry7T1EWERdCGaDFKP
fKVrsGNEzZn06VX26AIrzzrZDLLcDdMSsDsnk5aRRrlmoIX6KY0NWDXHij9FuM+1
F/VyVrDRmLdQVWYMkElvOeBaIm1rsa6e0qksh9hxHiUnUrjzq0/1elCyiIMyzCrI
o7KkvCG39g5xKinO7R4NlQJPWju2bFykcIqy9/9gnaOXKaY2MQxwAkoz5JfTM3dN
dozqen8p46gPtMSj7i3nqAfpP6o4IxsaGrXYE9Tnz9YpfB3KmnkGbGCA+v+Q57a4
1G8NYGyA93clCLeRLJtmgFZP/piRY9oM4fQETTCvocevGpYH8hVcxhqEEBvcZF7k
F5vcqnTC+BpLQ8UQ5pNrHgWmh7oRfz8/pGqBgp1ePHzR68/FWmV7BjVdHy09Rbt7
B0d47MzXbBRho40O0EpcA58gErqrVjfe0CwE24O+2eTU0pBasEN5ITHPGfbVASkY
uXDp55zgIuiCinDfIHU+Rn/UeHVucugizXCmUX2de3Vw+tg2utPo4BUS82LMBJ3A
CXLKwDWAxwAsJDDfgiA9cVF79LsMLrqX6mCOa6K/yeNTcunLGQbEh7q/Lij4+EKc
rkLHpJGRUfrP14kQLETvO6cx2NpLWhVhJq/7ucirZNgjkZGF/qY+DqZSxJmd4fFK
9OFKowRcwmYbh14P7XT6pz+kdOxKruzyT9fXIIzk8Y07VJqUDp5NJc3cV6HpDPGw
5DXyfiZ6RK6yfO3aPeqAnqGDXaTYU96VJj+gao2UGo9c+91PXZf/7yf7jJQrazly
/p/Xyn2ES5jlqwpiVC56uBtrO973yMFt/dR65eZQw/0c8K7NYcKcrXceYcA6UUNs
bMNAAedzHBy+N6x6OKm3K1NzWmZppZghBX3zdjWSkB9S23JsVWiMPnEuHvH1nT4O
m+nFZOHZo6VC0aivgUJgZQO+tW9erTbWVk055ZisVDGDH/5FKmpQUnbEZkQ9E+d/
FBTYYSQGWx+5bHhFx5SCdh20MTSJG39G7KTICn1kSjp+RJdUmkaHna5crwnaVdSp
REXIPK/95vdkwytXLGrodd3vK+ZeZgSFwWLpXcOU665PWszbcnj3IkjRdY9vZsza
fBh0cMmjuLRL1zb8fOXhKzE/v35jhxvdK/ayCJ4CzBgAZ9Mwm8tcWm5CDgXm07jm
XdoCEKahLep6fC0E17J70u5+iHcKw6WKJzoMU7XTejS1SHdxahdAS3cs30tpRxpr
BPHQ224PeAXsEDN8HkYSthQKa6hVb227pnlHtozQOss9yeiGh+f4N/elGQ5pezRL
g3uhxJzfPIOr2cVehIc4Er0fLsT5cPgqW4Nd1CZw9wMZomdWK+bNIQjLNnPqRwqx
vEE4Rc06l1UcK9Of9pl+Jm52lJamFR6/tVY59us6jIcnexV51/0Cekip+kAq5Fep
UOXZZHe7+yFGSXHDL4hJvkzKRXtioS/UWzIN9VONZna1eSwygfbQ53O2BBWekJg4
yXYmbXULr8d/4uHnokMbVYyrRwfpLUwfho8IL5+y+NfoEeuzgB/1DbN1utEGe41o
QNpgeBxD2+C7ucyH+nwWp6pjVF7WKONd9ukCoJC95OAJR1HDNgch3Tkp/9uh+Igh
hL4I+2qozSvjZLHo2gbGFrCkGMN5RLgnPOwquax35485ZlndYQM27cN0R8YSdL/i
tG/8tfx14CbfWNURreny3W9tapFXx+jex7Y9/BrL8f76HrNf3Itgu3LaFQfkb0pp
/HaYvTMJzWR5YDM1Tn0LbHh/DSGN/bYzaMS6zeJCRhFBkEi/RPhiXjxi7EsZOXxk
LqDouOajor2OwIH7OcOIlU8hLKRHA0CvahDF4dww2Pz+J4Xgn1hIGDF0t3N+nPYQ
d84nzULqSGdhp1WHIDpeA9e1CNAFFmf0nekee8yuW3CFq1VSulAQ9qyuCoFbdw7G
a+mffLzF3cDyIz4zw4LfzHmvJ4H5sIwCpkb34lARHO4AjAuR+PDgz5BtuJSRsI74
pesp/hv4NcG59kbHjTASY/J7zFQTAimlC2MOWol/zsxRB5/kzeWFHoPZyjA1e/po
iWAU4+2rAJ1MHkeI2/tNc1gYeF85lwGRO5tgkEPhGFzpsmUFJXOuy9FWG/v4plVv
zYR/lVgtuouI2xNhgzrRTGIDJpQefiym1koKaCAQq6rmFT8qkYr3cxQwK6lt/juw
rr1xsc+PvG5mfA/SFYRkLelbUawhWiu+Ix1EUBZP/v8Hg3QsGxxTy20s/S1qVWCm
i3qEtOFaedpyxQthO7zn/synxKnPTkeyr40+K3MHlUfZyB+rwQOsuHNQXrTklJmk
amDMOuZqwyFhcn21hdIT5CO+SdhLIS8wLyhvJmwzHn7eCTfRbt/siK0fGXex2JMq
9AizPZ5NsgUofVwINPxaqywfRQkNJry5K83oNEFYOJ5nCPCi3eA4wKZ5csGzC9/Z
xQhOIMM1ubva7zaGhKejW1buU00JrB+yYfACBmmjj5Rg93gboK9XRnWSPqR1fh/Z
BAodqGl6V2xmsVmB9oRjJb1OWBi85t5ZJQOaablIH2F2mQaXFmiPwsDk+YAdNaTb
JEoRy9uB9MQkNlB0ziB+ZSvxm/bh7gh4HCKnC5q7RufYT39oLx+A8+RKKqAnLVPN
9AIvY+pOW4RuPZOpDusvvgc94xgFbpEHKSRrgSEmLYxrw4r6clJxP9L5koeB2oio
Yg1QI2VHMH5jI4AP4EkBi68xpOgtyJXPR5lr2bP22ycfzUnlbXkxGFtWi2gbYQTL
U2CRP/KtwaBp8dgbpVCoi8OcoAekrYnbfcXTtgxFar5//MBY+mTS0M9iQtI2n410
MAxwBRXp3aIvlpGXkYkkx2UgvTmjzeEhiD2pCd9LSsEE0ZXUXWBCOiokkGpBQWqp
klSMCrMgp4TET+7FjCbTRmlq1X9ewYfBhan6gpr796UDsq0H6gOCnqiXxgtsqmke
INT3humj4tVqu5r71xctY53Sbg3It7CNLwqbiS/XWTn9POB2iSmttfVzCcjTe1Fh
me0r/1Vh09ODOKZ/rf/daQHrsRP1GyXOCh84GspbMnV1RSLHCsKwUX0nW9PKxt3T
y6Z61vsvoD1jNglb8CGcHIsWLZi4Ipk8s6lIfmKv4wRW3aclIr1K7JaBXgYFVvEe
s8bYYey/McMV1/3MO63nM5hCLN2iBnv+dlDGbgWYYex+Qg6CMfp6hONUILz0ElBL
t6eYbfWBkjyDMamZ43vNSdinTW/ULGpn0/9GFFAAp0TxYDqNXiWrko8AbBFWGnUu
sgZ7+RrRgycb4yIcuyRm/sjiun3Kf8yYWWbeJuiR2EMqyXpKjTAd9a9LStJxv253
tEI+5VWd6FRxMkX5gxM4Ed15PnEsGxFk3pxmZBu7MbFCxz+sggxbteLJe1MmNT2e
dsHF8aiob6c249BinPfDQ/fTBKVgDxp4pna4cz9nQFavWRtbcjhlyyqvxYLCu5S7
TJebTI+vTX5coiRLWoea2hkdVggfy1ZBSA2cqxEvY8IWTUy1zLrGyY0GCslVrAu4
NUoBaSHEMacnI3KUfNygyNwRib0OcHQQNdzjKRSlEpu2eCbeemVpEYaKxSkCl8iY
RNppAAHVt0AMQcORrCMmmTD+wkNLaum4CfYo51RXc1ZzrHcA8wdIr0ytrV9PTINT
Yjsa9jjVbWne90xYTAwjlCO5iiyQC/qZ4yXsRmRe7OL4J7x0dZpoObS5/+pUf6fX
djfga3RapV+uOPGbunDWP3vD83MPWooWt3g2I2GD74jktUHIfOtMBDEPxXcmQRlq
pfKAlPiSIsyBx8OlRW6CM6pN9KCS8yvgTiWuddJzmLvoiKTbsVaFw/SDnCnSWNUn
ZNibY9e0cvXOj0IrAfFvHCnA4fkKBhcN25/Etvrv71RibH/QYGuqKS3TwtFjN6Tu
wtdUNsReZNJjU9rLRJ3jhmjeiLo4VpvdIClw9f+KCToxoMmDMg4zq0NiB9fN8FPq
q2orM31IV3d7JYM4xG5blVperfeqcbn+vfVY8vogDD0y/1TCtGNBPXMIDp4GT5kv
6KeyDa4vFTgCIN9KeEnZvDAlAo9XMA9XBIbzc3Q3VxOc8HYmC0qn+sS/QK1OEkjc
M2Hfofg4IRYV0jZ1yOKZhNVACTzmQiJ7aGtQfSIq8h+G/lTz92s6CilLZkaP5YgU
/DBGGRNfG46X3cqHqWqyEjKG+ASawkO6LaKtMBsD+HsHAWLaWBaY7L6C+vq+xJF4
S+v4iqBbcxf4cS3+aPzElhmn7JCciNQDwVA3hrhi1h1LQS1oq6J0+8qNf1RNZFUc
uSDwNIEvSGYV8KGMF0nqNVTa1lg26kTcdtf3csp0gxAzZBc2O7JgAM02HFhJfvz4
xWvbtIsMOQIcX87niy5eBBgX74KkCjKpmI4uuUxh1IsHYeG1VOYMZqph4i9EDqxb
1R5Cfy4VkLOiEYZp0nTfDDLSzUrJK9VWs/y/dFwdxluB3xZPR/SLe0JZme89m1H0
4Aae3ATASMORfMC7K1r1nXIbVNOdtCewBAZpxWklnm0s2iKFAFcLbi7oybK4l6mS
/aGSmQVOdLMX9874UAq2ZRN6tO6spWSdjb3WUF92V46S4ODxyGEoomQvIFpwrHPq
bXhY4cIJ5QxHaPj9YnOh0m2Zc+1IKEOyu8wrJiMqX403LmbHR3ni71brXq9yCZYB
O+wt3ZNR2espKU0UbL9UDp+HEboq3/5NWPCbq9EYkWjiIlJ9AgnuouwamJ1hY/Zu
0sU5eMzhwi18N4IE7aIUgXtCZnlqa8pFSAJACOTqdUBswqLE7I7L5NrigpbeFDlt
tp/fUJJcRlCw9cGkzJ9DlNlBfooHo7nsXeNV+z2TtL3EVC+zQkI+Xjq97uopoCCH
wacC8f9+QM5kRKMk1jgY2ONlCzw3S99kYPlP5fBrp5wbw/qz2RpsiItIQBBzbqKT
1mRMAfEafJQ765BRot+gYTpZG5OtDrbQ0CCr6WlqmyprnPi7ThP+9zFtAxPwtMUP
Hx82k7ctJuGzGHd9BfXSGWfhLxTdfGpxX5D7N/hr3FSigtbqzJqfUmxAX17Dkxvb
OSIcIgWSYuP/Q2oHUGqGNonZP4lOHXguTH5TkOfgTz65xyiFr8iVo2yFqaYg2B/x
ko9I8+1k8vXea1RCZGrS70j+wnr83QP3TTkc9YMGfbIoRXUkBwbA495qUstRoNQ+
ivxtNDvaacGzZ96hStwMThafzMM1NXW9+Ttit8rWm3DfNL0e1vI9kwbH1IbfPsuM
/uAcDIiGmvJs01JQZ0siCHBI685eB5M5qdcrFl6QNOknwHnMHi9B/oGzMP0fCyzL
LydDwUe03x84FV5YopvBg5SgiBQlQV6wfnM3ZwIN2RGGzmueI/kVjmb2Z92j8tJG
ycVkID389mwxKhIlCQLyq7tUFGeom0nuIQjAh4URYkAKmId8ckT5/fqLa2Pn+Ndt
qB88etpicPdAq3B3NOkGfH3LGQ4FF23nTRLEJgPOSasinvRgFsuJo57VKg52APDf
bQl38D6owW84gu64S9i5WiWHmF6JdpkvN532hjpQfNQX/ciH8EvQd2xcg7sJy5ZV
G0mDfxsZ8lrW2vBN2UuDGW/85Gn9OO07PDhLhq9gZg+ys31vxPGwCSpPASKTxOhW
NNcypWRkMrDZQ64IQg7C8Rc2xM/6Zh8bc9ijkWFL8UFL+zazNBe/zNVTQNgiBDBB
4yFtH/nNiFixoje0iF+XJycRby5ysUux91j+C0YU+DF4Z4xZEfbdTL6+bQ7J2wRK
+ETitJEubS13oYj+PMeZkxWZhZuWiMM9sJZUH+hGtKSham6NGv6u2yqRmi2A6qrj
Fi4tv/WHzdye6tUuHxOzuu5Vv3OpUrfBw4vrGjiqyRc7R6HDeIozwjAr0IfUZoWB
FAD3SLgRO2fVVUyPI50SgZE1CeBTOO+FGn7CGs88s9EBLOA6c4YdhgqC3R98zUDz
u3/Oc72JUQF2xLDmLNyHDQ==
`protect END_PROTECTED
