`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EdPrAQ7BNwINP7xubTISa4to8XOZ8/Y/BuTZBoNo0bSVekCdWFUKru56fIt0LKA5
QPn+z9ZUS8GD5lik5EKe1g+AI6lKTEf0ND6ySZg+3+b9C1Kt5ACvn6uVhv+5vAJU
CXTdOuNaC+/vc3NAF9P5QR9RBTJxvXi7YdjrfbAmzY7d1J749geN/L3yh9dsP1kf
dqOFJfCrhcxedE3WGBEQ88pSnft41eOmm4TwNL7C+IPE9B6sAxFB6g/Zmbg+vFms
`protect END_PROTECTED
