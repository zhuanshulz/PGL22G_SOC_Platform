`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PipGYKUILuQmDdjMTXiEip9Mohbnhmf0vS8OodbW0dD3C+CpoEkHwtZjjJx7Z690
R4Ag4CKwTszf/3tBqrIob46D67IdGttTtZbjS5DcznKhRuwfEdbtyTyQ1yJxq9N4
WHkv0QNjxXhKIgcIYuPHN5RyPwnLfPh4L7lUis6bIjaHo8mR/hTscHatu0XMFYIj
diwN3cBIBNDNppKl2lcN4eU2No+0G7W97XvtzJ6qNJFimbfWjJ5rvcYShMpg7NHk
oEQ0bBWtMxpKzXc3eme5Yb3gYNMkpmrzTh6eIQB/1v9krTqJuYAQAdPCEdJnp899
HXeLHSMBnsZtlULG8aG4HXETKIXyAd1h6yPsBywmCFDv5MjvM8byppmYOjXvZQWB
UoM2AWbPKitMdRn6itG1v7e602FkH/uulvC+Yrkx82YuSZaeU33DBVgTB1qTbjMB
bPWzXdAytt5C+vWdz/XzV9+Rv3flbsWSCQxZFLuAVKa7A00S1qT8lqoLjpiFSycw
wZf2D5Izz/ppaOzVdiM2gcmzoiobIBBNZlVShdattSyi+n2niYar1TjSETa0xLP+
WXvNHgFT6l3kHHgHuIhNme8GOUCcShSwY0Bz8PSHm8u/zJUxs3MvaASmZhn88fi+
HRYFf/mNP7tdMNnSQsyehZHCzRS809aEhCehS3K8QJHWtQqW8AiyB8vcIfJi5DXM
NuTAYBeZJjL2rxLDZXDiMUgMVqX1qMYbQBMk30YOw7Lk7/9qhk8j+kFpgFbCpiUy
FXJI5I8nVNyXP6OZ0pwaWsIZHTZ3wAMD1dcR6rexkXkV6M/niX1Epw3lrkYZH2Pd
4k5iVZLAhgQBFdGU9PDW87jR1znsgM80jKbLG4vfrNNoRssWfZLfJ13GYDwx26HP
dQn8KSkEN+yqiCTLpHHtsjlXCz09vu9BSLpgC1yTsNZFTYiz/LDogv++LpTRgbZs
PBcJidGd54IjzSacqLi0J+hCR8STNFj4uuWNZ3v9JpBKyTfsWx/44N3zxka/9FY1
Hcq2hs3GNSDeVf1xRi2A6Fxw1Sp2v0RRVWvE+oOOZ5ZYrFGHZY3oqBTdVu61uOyD
KjASnjUGDF5H8CCgLfDcYwrBto/0wFmOPiLA7shRLQsfXX6ynrjLWHLdDcPq7Tur
PmfVGDHDKj3T7cTdNkzWSVszfKS+QfrrVRRA6OpAmUYhZsa+mpTFanHKCLl/K192
qaSRFVQsVJtxBEPOIVSy9dqSuAocFZdI+B/p8oqOM0cbu/R80czj0CTfgHV+OdDP
hD6FPGOZayE1VWbpQs3dP65Oqzriba432+nio5rBvQ3BURA98U+rOEH/TZA98OQ6
Q0g1Bhy3bB8WiZLfiX/6vmU0aV8pBtH7eLmCVu6oBmTBokY/2xwQEHb17XwEWKBp
aamMl/Gc364xxkIwjDIxRQQ8MAehkYCCdODwowbxitPVUmUc1bHpPV8qScFvm2uw
Noyt3I/kSSenu5p7+qLbgLN6/MU0kjr6yh/ICHGmeqtI2U35frrUnI9R6rBjqNKJ
KCun72BHcDbHaQdd8/NGz+JLdzJFPRpv+YgePJGXzzVZcgqxmkOV/UJfftJKukMu
OwKTgjRZWyQmEbi+lE/pvP+E5drDqgScz/2qnaATrme8buRFdRKUQKUiXoTwBYhD
Io3POflr2LHnBapw1uxVG5YReWhYj0VVWpDNhZN6OQRCFt76PYXdzYZKSSuBIf6Q
PU9catEmoHC2dx3FnjZZDobNm9gxmspnI82+75NJ6W3mawWMm/MfxGl9msRreIBC
tvfgZ9ejuKjT3S+SpeCQDXtBoBhWNNaMWB8RP1kvLO6azjFzqeSY9iqSrGLaV00K
xMk/xpjdIxLHaeME9q/bckA2LBxsPv20NpXUYpE6fRojJggd+HXRLTWBGmyC69qX
3GR0GbWo5qguJ/mjtIPVrRU83af/8x4HSIMS5O9ToS/MzcNpTYXxBuUUI4zNMGgh
oIh7kdPjtZe9P3L0/3cDqtcOE25aUJlDg0gnN+h5aXduyP0y4PA0sySJdY5Gsnom
16Ou4dp48mAqJW5/+p0jqzLXIQlcHGskKtTsG9poHYMKO9zZKK79+LBL245bbbBV
RT8B8Dc72Vd1cf/l93Ij8HFQ3S4Ff0W+W9Sj/1r1bQNAfpbAxyIhcXguEq5bJgpN
b+rQOT9oxkYl27zdQDl3LFZCTr38Dn6rd+fbn31ehb9s7ugG7sJlBrxVSQOIfDnV
xcvW+MVogPw3i0YSwBVRVNV4HFp0QprOkiYh8iIi0FfbG3LeI2btSDtf8FvzNJDS
SouVpuJc5GF6oO0Ql4vlwtaXwNCyeWdnPkUgc3FeyYL5jAXAh9YgTLyCcTd9J3N5
v9Jo/cqdDd9tpZbfH15llrdGvchTUttEhhb/0Eag/NmZHdIMr/PZZPq0E51FDjww
7+Rcw8Jv57yqCl3T6W9IjbC2CRmMCpzsGOqgVZPkl3fbRzMJPZ+zTUvl99T7V43w
83roSfZzm5GX0YXilyLODu2UtdnNMlAw+MRodpm0MzsNlck+cYtsWFDRkbouCAg/
QPZ6NI9aNnap897ss0fYx4muo4n0vT7EqkkSk1E4XpZOPAXj+iwLP9O8eUyrsiZ1
6kkVMYHHqdirY/UXU461X0zvvSyaejW3gpLXu2Eju1Pm8U2WtSo2j34m38xkmneC
Ba5p5UA8Fit+EBwuYtVmxKEDD0E0bh63BltRtzzAI+wDu9yjM0o+huAr10gUTRZL
gPsXM3TE+nNyYhetZwOgJaRwxyTk01yePvU/ezD5yKKvAPdhmnEA6bBNWwbxM9Z3
gi3mF4FWMD58iDnw2wZDYFEjeLUwt9Nfky4ZCbh7m+jDn4qt37HifxWNkM97b8hx
kXL1WEkyNQvjhAqowx55c3Hju24G1J6XWTzc8vzqY9sivzS9c55fb8yowsT0Y2WM
cgnK0vtdwSuFaUl3XOJIjKr07+j5g1gSbeRkK25Dg6vZLuAhuUeL+osHGVKHL+xl
+ia4ozMOUxZB35jd0ykm3bs3Sbbp/0ONOFgpM/L7MCqmQO2XblDty2uN3Ccd/TK5
JKtd01Vu7C8B6FwYUfpXORmxjxA05QfygJLWONReOjMUVS2Gt/re0f/1I94bBa06
NOyJVk1Px5PhFg8+Ct0f7a+/cLMcK3rP8i0TvmY1WZeKLtMUn5ZAQhX0vvQoejRb
Axi71q3WX6LHr4S86ADy3SRTmVCRFtJH1sXFtvCJ7eBHk7MfzcfjupNHTSOpxil8
EPmr7D0pMK0abCRxdo4g+GjYxmyTD8hveV+Vab6HI1k9SIQWGawkZwq4vrge1X9B
jg4HrRxvTXSYwx+lvEhatCXpkcO+X5zh+nezvM1utAr5jJbQ1qgc3EL0wWZUZCCW
BkUxYvADFWlYMKSvEBk4niTBp+8YMRfCV3cMsLGqRws=
`protect END_PROTECTED
