`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qzCixEpNjKAjMLxwvlk2zWm4BifBMk4o55sH4r7x/LIAQeLVrgDlSHeirw7CqiDJ
HJN8ftow0jtDwWuZG4aTcHXEv03Ecel8oMpoSa0dDguS0ZRd/9PTagLnnJYozepi
dC6r5kAZjWC8eEMfGvN0A85PWnOWbNFQ/sIOTePd5H6xPiReKW21QKztB1nXZ/Zo
3IxCv9AKkpu3Xeq6T4E0ilTv/Nosbh2XrmZHLROxCxql5ZDr/xH4qa9XbWipXD31
SyiEzHLLlr48XBlh7/WUmqrPIcaccUj1LSF2SHzqfEn0i9512bgLDSsHMXy7pynw
xJ/XT5v2LnihYnqjHoV0MRQELKGX5aLVA6SVzV7HbKuKflJBEVxOqz9klqAamgVS
dZ2nvzUY2xOJjbc/eELV8JB732Fi7qYtVS43vySiW+0pMczrv872uqZ5Mu7OQkx3
vGqLi2flz7AyGzGstN3VuiLuLqftjw04/89DgA7w1GDXl0ozUehGUtzh1sYeX/Fj
N38n65NHF6LwI9gIzTsYmYRCLTmDhFbYI0exP9RyFaJJqLCr8tymcWtUzfXiFg+E
KyOFTncQy175it0binOM6Gc0KXgoYOl2h8bgn/zL0Abvvn8Fh0h4anZAv6xXRROG
3rXDqc8JYUG9/PFLkG6Po1FBEzj6d+mzwvUFWVIyzB7Td4SGYd2gE7vJeM930ulH
32A/BJ4qaz07FVlmTpM5NvAhTXcQz2HPMPFBWjaI358aflK7PTfJso4K1bYfQ61c
QbvRi8BKIhiKoE5Nm8oFmmdMru4go2EpMOmImay33WDq8BFQoPuGAMyw2vnTd3nm
7B0+0lXAlr4vzjsIovMOdodCRwQ0mTYifMAe6iBvtwnlRWYxAuVTZMUDOsUTbakj
H1cM0cDdD2j0a7zaY0fUu/DcTQCghjEKCOUghpaNhl8Beo+8eD2/WexKi6hI2Aip
V3XVCjJ51fVhoy4TdwNbo/521eOxgaPBQmai3h/iQucetZXFr0s365vgOpCCA9aY
usanyxgAZZRXNpg+Ue3jZ3J59lQPmjSk6GtiCBtk8c+Vj2VLXBZ4i1FGWXpz59xE
utGNslGUJRg/2e7SyW/q+kPQiq8u5jubvRjVBjACzPmO8xbkshZgA0iVpQmBzpAl
0IEggcdrqdGa+2aJkpvDtMzOe629kQFE9h36hh+Gshe9qnkxzZYRmIdtNOFKSX/p
W9fUUdDyLWVCqSXKASJ2JWRTz3OGEMQ79EnmN8Btsp1HLHRm/TREoPQO2qNCBVMa
3x5Qcv4fQqvMCWVW5k8jowF4MVY309Eig3WjydnatttWJf4T5PVPip41+GDXgpfu
4MZVi2ChWeanblt7fduRHNesVQoG4YCsKMaRJZ6lwWUMA8a/g4gmpdsgzGHDVFEL
JtY0qymIILEF2yIiy2mUjiIdG3cG/pqwggUiO9oLA9TmXzGgeMj++Snyb8dWALGK
ty4Cth/UCF+WhKPfmbSyeHiRXfo1b8DPuAYKFgzfCJGdCklANTwOySRhdJUsKwqb
8+qSCmKg6v+d84teOInQsoNv2p3prJxPdQhdv1je5dfb2lekfncJaqtmeeeBx0d8
RX+05Pduxh3nCtXhFTjI07wR4h7zIRUWpd/Kr3AP6/+q3V/OYUTWGUPakgyMnLoL
IHQe6zOgm6QEqy5G+Jxut+x7dM1zcA5izcu4l5IU1hnIqcxJ0IiHgJ2wJYAvwThY
+uFLmLw7C47dxUOsI1saVexp9gRs1hENsAV+tvnIXJg5Fh+QbBvUicay/FD7GJa+
`protect END_PROTECTED
