`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sEU8jgKD97GxE6o9MEhNxSl5GhWXW76XtozV3Otuuw3sio9oLnnt7Ap1pCGzSYsw
EDOfOQZEDJgTjHjcRbWcqHfDO7FmlFYiP/xi04s3AjjpwdnzvCtFby1t2HTITy16
2FAxSYnwVlT+ttsrpezPfnabsLa5ywhD4hp/8S+vyyrBIgIIL30mQgS5vYywG0jm
DMIcXUsrBlF/GKZpSAvA2QxjfNOfOTeSYmAUfjk6zIHrfHsGzXqPCvz7gzQaLOXs
7XEy9eGgDFlr3TdrMPQevJF1ckDudodLyEPuIf7SHH0z7MX2WtycwbGTikX6OMN4
kXLVUVyZPh9heFgWvC4zXjHvK6u+XyY9x9/UbgKZ1KzxwivCYPWeh5qGD2McAUeC
ZVeyQzGHY2PmLPcElcwNpIOg1HCChqrU0qbQm3BxvByoSwyo7TQ3qV21mtOC8TXk
Y7cjke/VJ+enltESeP/FLhm9dDI2j/7QFLYuT71/pIEc6sIh460WGuHItpLy4Z9G
QWhJaZaqwNVXuRgh94/apyKbKmfKbwVaDO1RE48T3aylujuJnJOkoYA52Pio/PPK
AJ5xNcJ4P9TX8ScNqerDZPysdkxdPbUv6BRYE+MgzZeW0LQ0f2htEZ7JsFHbYypM
iqiXOQDvm9dKUhSC/Hj60wErcNtm1JccKKdX5YyGgn97jH1w2evhopMkauQfdLCs
c4lkR6dV54fqRdTsy39wlQFO9nESjEmZ5XwwWxolL2z6b8Vj3Hd5LW3nB0UjkNxn
PlEnr6obka7UXYtvhbohpfz6+b6px0XnUkzU8obFNLInHlrbncEB5hVW/LJ6UHPf
tRiOna5jgoaTTb2j9R4s9unArTjLSXzx9Xne7eLUWjNNmqmRd23nEQLHfVKBH5ad
qhciA56x18fcbpyd63lCQTHzuvXK0Jyr88pOImGy+LR+y4U32aQUpuDozL9xsU/0
g8+vqD4dCJsSoVRT6b2OeGgGG4qaQm8FIQg3RVZiXxM=
`protect END_PROTECTED
