`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sK6+17c/pkTzcYSLfyDivvecfLJWiXATBRIyro4MBVCQ83MLbDf1iLERgwWqBK8C
qmKHM/ozX9q1qPJS0moYeh7HUCNLZRfu5JYLtlIQwItAU3HpKg+IviKQdSPYfiyW
5JZ2ytRvpLIjleeePkCaS1+2G71CJvSNVyZnxG1vJ94f47TJSQhQOlkhMo7O75q/
I5fo4ChlMVaFtcRGm6VRbDgXfNiQYMvMnKYohNF/OIJpR6+k8dfGGU5W3klyUWyc
cbaatp37/WylyqAGI7u1CF7jVat6sBFNHmm0J5wIrmK+ke61aJYNpAwr34lJJd1q
7VoT1nkOPWM55oG+Ym8rZu9TE+sx34ixVq9pJCHQSkTyUuNh04LxsOtit92F2Vl8
1Y1dFqdf1xl6UyDLfSnAM9ezKVvTnpDJUCDErcyIggB3PQ90+HypGkgsZ1M4VwwK
5i9Rap5IsTYT20B9dboGj7Gp4x3uNf9DDuH4YvXjV0fAlc7YgXbIBCSQALaDF2oB
kCG4Iu+bhyjvSqruCfSZcUCOmPWPmwEwI3YcMwTZCJN+jmka4M7aK/WzqKcNpA9I
x34tg1riWw6f6V+gmJVzu5n5PGQiEbuuWt8RisuLanmhnkNsZEaCzo+B6afwdqfm
A1icTyWmXrhjtskuQNumGa3N6JEEf+oqLMBCbyqeO0gsDgnUsTk42A8i4ghgbsqO
3frKpFWYlvoaIvk78ZgPy8ilhiLOzYhKxMjZg431vA+q1RQKJsyixZ7Ajo7POrJi
RrQ/gIQl8bOgMQ/Bt9g2l4BFOII0d9NrloI7VJdkml7qdHkgEdZQe+YVy5csajtt
7iM2BYiiTdG99Drrcn5z7Qwc2jBWnBXcnHI7pEgt/9LMUsOze2nqk3+S4B4vf7m6
fWsB6/51OzTHmYMJpEilj3uAPQ5xDgbfkHc05Z3+ZVYP10AQ/BDR5ku1x97fyxpC
0wYxBkSEtQWCpKrg8QSw6r57v7JON0E4nmSioan/geAi0lFHNo366BPyA64iYkdD
GTczeHG6z217JtGr8DtubcXDnngYW2nFyne/exILaTbBBWg5LYFzxGcezdCCYIca
ZURvyOmzpJMgc69EiZ5Jj4TTnC5A7a0fDoy8ZEyL+swzAdzeO2+kU5ZyGMu03F3V
i/dQpmwiJ3qwIvqBeXja6CT4nyJPRMTMKiOcamYvdZVGvhkAeaud8Chj9OjvMMbY
b1Loex2XsAsKEzB2AgJEOJqCLEu816ZMDuxZAtOo/ul6N7UXtLURuZ3BoM9nVwMk
Ol41UdJwZKPMeKBNtB2mVAiDMYoAbTSVNM1yi63Lljh4ksUiU4rq+Cp5l77Slbln
iwNxlWbCUBeksNMQg+Ow7LH+2sdJ1rVpjheS8iXstAT9ZH/BqpxN7kf6daK9kIuf
tfPskBSk/jtMCWQ/+MLeGoei3hC11GIV2j59H5WKZ++CG89MuIQooFY8tCmQXMMR
xfPV7HTOlds1j/slFTBGfmCu+lBxJskXq/JA5tYtf8c=
`protect END_PROTECTED
