`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mr6gXk08ORnijBsop2idfgckuSqvS5onFwSFNftsOiKjjFMQEIssRgvOZMEJFO/o
zqwBUMy/3zGjv37eUJ1wakOulajmjxn+xyXloyerkQhqd3pv2wGIb81dbKCnov9m
X/zrAnObm3P8gSE+POeoZkvRUJojTQK+PXiqQX1W4iiJlOHyyguFsl019ckc1ODw
Sz/f2wdLJUvTnGWKIbPgiM4llYCaNqXY0WjoPy0VmU/mASB/h73qV13v56eOySb6
Cs123Q/70TR6tNUJkEdtsKuAcJguRjPWpPPcfqjt3E4kd85BNGStkxRVlnOeMwp6
qYVW4g93OZoHzaUqKGbRYIf8kGrQm/1og6SPKoe0T6v1n5M94TQlrJVsgc33p3hA
FYE4BEHA/31oRnuICJIsXAJDJ/8/j4Nsy0jCXPnoGGsmV7Damy/DTlINUSJZzzsd
K3Wr9x+wuoqJG8cCDTOf1ee9mc/XBbxn1BMGnamzRo4oUI9rokxKLFb1X0nnHB2f
KQrnWgL7NLoFp/AaUpiLNLxhOGSWZUmaXsOzGqeGQOWsA7xT3Mj4iStlHEaIGZQ/
smygaLjYDGCWJt/K6aHn3We0krheFGCL6dtkXKilPt5cD8IwOcQsvuGlxdxLEnIv
8jFL/Vgxzu+P7l2iuavNxO0aVVzBa/ne6AdI4SUEwwllBQvKhqvn08KpByFh6EEv
sUTovkMxyF8aGQKCqNgKaFwo/ThGcH0QkCnHpUKKVjygASVyCibsu3iTpV1unx8o
FgBuExOzeA23f5EKDttPzMzBA0pSrDGLyqBcFI9Gq5oQntgs4EIggVVm0Hbdcpfp
GVI4rfUsJ4CA1V75bhoIhl9DGdZZBkNu2Dy7qq1RHdRnuoiFB6Looi7b3rH/znkr
OxamduHYSYgGX8XL1mnvHxda8+bzNILqu6NQ8MM2XLxAHvyL8Qo8ufTpUjN1USBO
8EZNUouw8s3hMHEEmw1PlS0WqWmWiR74roLZ/VS1qoN6heKNxZ51/SOcTPs0F04x
2emOsbCW9Prnv+RTOpRGs0rEHl0G5Ztr9mZQUbZFTgonHsTnMzzF5YJ6Hib9YS1t
9rFxJySSFJWf+TrsukRtlqt0VTTUTVXPIfY4em2VElMFAjcSHCSBQ1weohU5Iebs
4pe9onu+l+mcatMMy8h43zSXQwStYqR+ZGZ2tIkE7y74RxsUQtbXrkSxB0jyQCvo
UWTinTB3ptReZyUIm87PF5JM8MIG1ZuDkfELWLBM6ai0VW7PpW6pFFMLpGvQE5nP
8V2M9dZ3gNb0hIxwD9noC6oTG0OEAYnqUU9qTvOCi5NXcEywdV71kYn4g0Y7SxC/
/iqFzLxXTUmH8f1GHXwnsxp3ROlXxm6Vb5cx6Vtj9RfqEuUGqCw1vNjcA0pcNZSH
tpvI85MskMW7byOj4s1xGH0h9eeNRmgCZuQvhVxtXOxfIeFnS0ZL1xdg9uaXEdBM
RJCrfp2iHoom8DNj6drVGtnrSAoe0zZVWKvaUayXaLxwxMDcUE9HfPoqKL0S/RXv
ZX6N6GlhtpB+NbSgTRNTRtLXJwNWCo2X27TiQZ2KZ/NIHpW4auX2nZ52/a6c2qST
/mhmFK+Vb7xTHRg8kRTIsq3nBKHIssT4SyLuIHJft3a3smmX9aKRujMIF+qDDA+I
qTF/uELUZwnaQtAh9K9Cy/pLyDRoSKQRs7Jx2448mj2oWead3GoZWB+LYrnqog6c
tBenapGtwcspMLP4ZPy4vfthknBT9nqscgaRVJHLTiUy3QUcgvgzp0wys7VU5tWL
ZS6Y0mxxGyVkBsW9BlxPR5pmJx5yY4IZI8T3EvpvQRlS8Zy63DpmLYIeBoHUEL7f
5hOw9WTlUJzHxF2HnMCxilN4Bd6hlGTfrpcO5vI0qZP98nsTM4Tqrt4vnIbUrlTV
kf47Qs+ImdJdpa/W2vbGM2hH1QWVVIhQRevELShpeBUqtQOV7zorjf6e3tOsp1o0
EmNpV41NdlNi7ozNrS9xqVKwwj3Q1d2CQpl/unY9lRDV1lMdWs/+2AvewSSetuzC
1gJ+TbLh0Y1MZqG2ongL4GwL+3y0epGxcqRK/rx2bu5Jgz3Ms3hZmbUKHMXbyGuI
l1bRpIV8+H2AMfoM7IHjUHenMCi9PNnsuokGlG9MMf5KxDuj8BY0RFoiuMeG0nbh
ecX+Zx779HuS/jYnkXn7bvGB/YE+/NmppARXUTFCCk+01GUBLBGyyCX3YsyzGgAF
mfoidj+WdpUvUK5A2YAkVKR6bUPCnk7ihksQYsGUXOiVPJEAVUtjuJ93fCjN9Y9W
mmoh9C2SN92eeCRnr8EBCvutD28RAtD2oDGyPIWqsUzrz+Pa5Tx6S9fzkDxx3W5Y
bsRIyPPje+pUyGom36dFbKr8sxPx25PjFANZoL2aK0sK9fjhegLhkqFwqQGtkiSm
o8fVBGQnR6maz0NvU+HgorQ5y+a45NbDuvCYGW10mREcxrnHnInxgiFhDe3emsP4
OcxzmCSvNqR5zQID/cZvZ3dSsHsPxTRL/h/zPYOeByx9LF4t8rPUc/r3tbFbznE+
eN7VoyxTip+bHKnvvv6T/VAqlW5ZaXPgnsIN5Irjt20lQYk1gPvqyIEhURhcWPVa
579hVGV4tsjWLOWVl7BsrkPB3ZaN3doCVNqgoyKURblXSCm9up8xsOhjKM2pNCQ5
CqP0odhhgKTUBxQ3YswgnjxNbRwdpUKStGHq8boUJqqETJAQwmuZgcktZpF3LkY1
Aqvzx8D0x2DvrDNhrgXFFrmsEfUWQnybzlW8HMlAE2mxcZuYnkieQWEL0sufrKdd
SiSRFk5Ti6p9rWkUX6uu0cKC/279uJQIPUbmBUJd0rvpkW+78PaPkpQLBd8fOWhG
M0boGcwBe18fQQDAwL4/oYyjbA5g7rWLTrZ3LDQK18uV0LbFmTQoKO+ZdfHbnkKb
JXnI7cAv+DyHvJG9L9l6rIkYNros7UObrG3KS939Ep4MiEBMVUIH4ESEmwwPUhlo
b66nOvKOSlb/+TJ9jPledvhtNxCswlzVVghmempEzZaqrH4bWWGDAYY3H7pvR7TG
O4RvBNrH1El3KK5e+m0mcMX5IEKtKs9Yk9Q+0gRUscTVGDqUn0ZYFiy8QFKcKbdu
r/aufHIgjzQKNSxKHVktGmDLtkTe429DFxwjRzC5fU1LjXW+ttO/q3T+AY6u56+L
NIt4Bfzisz7wQa0hhW70P72KozMxjyfm5yaSB5cNzJPSE8nm/hnel1XSr3a0nKxg
1WGiNhLFakOp7KFYo2mm3DBbq1RdYzVvLui5zfyW7eWOgkKIsQG6IawOsT/HGtvo
w/aZGNSFRjrjHaLvJPhw4ZrJewt3b0QeG5t7MGl99DD1uPge7Cw+fRDNGOUZPBlK
QsdDkyZfOAxhOpkLZmRQblTMsACNHW0fTp6I4ZYpX5tuZLi3N5cmHdO0wJYMHKIi
QYfUAZgaeTRp1HcZhUuuopAXJ00+8s/dbw3Ol7hGPY+oC1wYvTlB2BTNArflmXzL
Ib0ugnOGesAnWXQAkFXQlIu+ebQEeLLIFAhaD8Q5R3aXMOpukU6gMHFAFTEHklcR
9s9zybGsBBdzlzf9adPv+BtG8qQ66Ixgoo8aH+aXl0PXEtddhLT34IVncoeun05j
9wVNQEHyQU3eglL7KJwJN0nZX1Xeia5BcWdXZhHxG75YSwuqc1VEtouRLFK39USH
5OuaJFHAkmVWu336OfexzgpohnAUgMGO7r6qN0MmL2JoaI8UBLDCRHK4kM/S/oze
gs85plbo2m3FlgSyjJDN76bcjbc3wWI2aXqWQLJMEPg+ItLpqeOk0VOA8Waf3SA9
PjvnNpitT/3MmdIdHxA1ydkp9Txy+shAHs95piRrIL2YAOUVK4jssXfdex9oWSOD
r5qcpf/BziRR8Uaa4zDgSP+/sEoUlbXKOIJA9gsykiRkxtytFoIyonqPkeMY1lzE
1tjJQPqFQCSfCWsxK/T85aUFPL2hM8RFuai/MxTND9CxhOfWqb5A2dARActcrpIF
jujiuDsgzjY3IDPybGQdlAIlrM5KaxKNXcBCZXIbjE+K5KCUqQVIKkDjJCwuPj7I
`protect END_PROTECTED
