`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K0Mgd2U6msLf5ptkjeXdLC41T3NC/NZL6sqajBkkP+l05kNfezE4gAr2xGOahQiX
DBc6dmLlIX3zzd7hMLcPObuhZ34BE8gwCX0PzUjkBT4PruMIwJ0biz9jc5ffA7+F
mexInSKor5m1FH1mvh2yZ2sKy4id+mBVAn+q7qEBgj5knhgblff1O6ncVmrq2hz4
5VP8+tVpVD5Z3AJpvVYAg7+D7py+rY3Zxe/z33NSODqzVJc1mPQVDvf+9yGhXZVj
xwYple0g77vvk0xe1A3v3/ndE1zdlogsmoJmjAss05xvofy/+pvKhh1GOAO8Ysbn
/Sa1U9ldAe6z38r3v5FosOteoBc8XQNo9bmlN2d/5WE4kR39rLH0cPxsSYDBcXg+
K9oDmyXxiOn4ByaPf/Jr+6SNOvuzhZt74QlKyD1bDlPwSCW0IktJhnSVIq/rkzl4
xOdp4LA2tOBhYZ2pOlyzne6MnwbamFJP1FxOm95LDXGNocbdumcQl2MGu/rTOog+
K2R/x5bF2uMwEWqu6B19EEk2gUqLN7q24rzJpMjuR+ixSb+HGxfE0PKtVJDHO0NS
nElfoEpycpZuQ5HbXgtuZSZpaf7PJGCYh4d2MamKLQKaPd80CwavXhKqJ/m7sOU4
8SIp/tj7tu+b6mvLCjbPMbtru72cmXS7cKPSy9Kz9DEvflY0lTe5q4NBlbszzBmh
32PnlSfksNPcYlwP/ah03W/bkpcpK2vGd7vwz0nRiAOGaO53twOa9QX6+YMJy4hR
WNEdkttaYezgwH9j3yRk3pDTHO4ZAr2ceZdNCQZq/6624uEO6ws5fKzbyWhdLRQY
EC27nz5omDsL3sStMud118hhIGlrP+3lSfL87byLJTFLNFrrSBzWZfo+0iedRjQ6
V6vC0L1gvteFMAhYgg5vu7DOV+SftW6+cUwMtLfFpjkpBw2rbW8ZZs6OGhlNyZbU
KJggB/d17Rv+7U64WOuVKcpWKjatfrS1EdFuQY4KZdP6sh3npB3REaYt8viIY3Su
rm1lJ1/LS/jtwRoUD5vc8u7gIWxqkuvNjiprR2je/FAd6UE7qO6tnPxfeygmgEUp
C1CBE/OKDUf0ps9BXEVbje87zm8WBrf8RbbLN3TqwY/mu5YXBxbZFhVom/ZY6ch3
TnjCLVZtt3aUBnRAx9aoO9Xt7isgkaDhG5JCR4rWfrJK+pqxPVNlYXrDv2AgnmLb
G9MJT5Z2KbVA/IOM3XXTxnLdb6M5YupjL2J29ggq0MsccPL14wIockw8Jj1+s1M6
f4d5Ob/WplF6VHwaNb1+Cv2p5ie4Q+YHaVqZW7WacbCXYyWDAUPAuRw0XRLNpfv9
vTC+ThCN5jSoCtZ7WgwVUS2efkAqNtsHDbPwUanhn54=
`protect END_PROTECTED
