`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PtQAF2tqkRukY2I9WpHF4d0UXEsqLtTahZRhMJ0tTIMyPMZhPseUIzvRSUb1TNO6
6HZmbOlZdxRsjWB+bFTsYpMW81gIVzP4Wk30N0ATOENOlDN3ouK6howmZF4BNtIK
k2N+ivgvxsY+2I1rGUbd7Q==
`protect END_PROTECTED
