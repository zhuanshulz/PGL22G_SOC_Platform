`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ycJFR+yhLnwvH4JLPcR0B4tiDmV6auK9Y/tR8MUOKWDIzOFrsVW0/9r1t7thEH+e
Z9E2kR2e6zUid06A3KHHBgPM51tDGlFBd+YDCUkcKj1g+eFxJJI1LKGJ2zUXwE4u
dbHEl6cjgYA65Df2KRM7TF2oTy//qXPewcDjt4tUZyNJdqODnGDey644FbeHk1i2
SUjm3+PlrJdyUnn8XNYjO8ThyXJ5B8DBixHtCRsqRHUlkX1cZi8glhTCVUaRq3pi
hx2HooeLSkznRYRFjhbmwQ==
`protect END_PROTECTED
