`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NDAaS4UShLOWSF/UMRYTt7MJ1wfdIfS8pJi4EzZxfghJyjbEgWyWkWKWtmna3yq4
me96oCZJ5zFLJGgen4V5WJRudrTk+rUNtkYybm8KCqjqqxVbBknFLlZ/P4CBWMFS
jmuXhZ0p50lHp07yotvP9rDz/6Lq9TgdC85OqY+ZatZi3uc+sqsz6Aif8c5vsBz6
EnPpP9LRd2DxBpki1UM/qneylhbWCZ2awE1kX+cL1a+bWfbqQp0PzZVejSts3iko
nHbegH0nr+mD0HJWEnmaVpSo0TXeTmuHBGzMN425p58+I48dZ4nlQsxB8oqY8TbZ
UpwlvSBXBDKn3Md53dvIjbqTVKAbbSLR4JBlhTcU8eaXUbuQyZ4Dx2RdGtdnBDCx
n4QrJVMJ+72E+JQKJeVBkwi91mAMLDmiJWX7MsNCKhHK6x+GFzdKOtrNnFXbyQDT
/MIhK6jqZKv1xPk5XXwCTsSeDhliQp5w1RfM6sWK2y+CWdoj5d6xf46PsXoV8/v6
EorDujF2WDnP2sD6SglQ2jPciYsA4e56v71LO+W3fG5Cwth7uyLm8xV54nACqro2
e2aX2po/C/A3zbvYoeRl0Pbj5ecem3pQUr3s44TKJba+2zPCyIE/3EMZKP2FeQeL
4e4ct9CfmcX8K1vBR8SDhgv/OpMe5v04wAKGjjjDozDQikqUA/FANFkp6kflzud+
HPKnrVP8qL/duUEu/qSvUmFGwo1Okli/58VcXXfLVdh8QXK8dGFXSwPf7lZqtb5E
Z4K22meCuJDCfXU7sE1CMidJnzWEYdrc5tL5uzPj7v4tWhpWLPC3B9DyQBb1NX6o
vCl7dBvwBV26KBVWuonVo1Yl1yiFYfMMeFe5bdXkaoVpc4KC23KvlpbueFRpioxJ
ZMUc8dPJiGqzrwa87U3xt4b0Ob/RG48u0rM64XDUIaxY9Tx2B6iV8F/eK50PMEei
9XXWI41NeweI66zMMc0eF1bLPJa2cdH9dcJ9uUWCR8nfubp+lCJhsTx1riBM1v+s
hMINdkrBHbNuX5MtuWha28wKObJMzUW0Q8fdOVNYoo4RW0cUdhqGKvZWoocmFJEF
6A1YvhpZcDhz+7J3OV5Xtg==
`protect END_PROTECTED
