`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t9bUk/JovDc2DHmhzruxPvkAEW32uyFd3Qtdfd9tV15oq5X7rlX4RfmpX3YaPBV/
J0Xktsu8QtnFnIFsb+m9OJ6GywfQvY92hsQu8AXc/wEjMGJIoJe0ITQ6aF43Zjqg
dsqFyRWH3cQvLXOqDP/B7+CVje20rDyUbwbi79v8jFisfEwq/U+k/ZeeBuPMP8vS
7weIkEQi0aXOc+SqfYrWOYaUDjsL5e8DrkcCNOpA8Y0khmqvif623woLt4FonU0X
dTt8pUG/4APRBAHtAFgLcx06CV1SXBSBc5JF9KBkMoGDupOaz8dMtdTL8EADtDX7
NMdI/sDxnGA9GuKKMuWwhV7MxwAa819cq2sXqrRCce3TYbziwmcPIObJv3gntQf/
rwZuGg02hModhBXCMt8vc1lr0anywCxvUytqeCzveAsL73RWSAKFjuqJuQ76zz5+
oi8INuCdumG2r6J66kt7qN2ORRZ2HbqqTqAU+n9wDLwmiPwfZDj/MQr9wNVxeczL
0Oy8MbxvHUEuIuKAC4v5tiJhBWDG5LHR51ngT9ykUOU5sR4b/UKum2PIXBSk82i5
DwWOg5gfbl9jEBU0GdeCdJZEJybTBbIZAoYGwkC0hWOdNAR67EhiQp7ryrNi+AWU
rI8hvk9kv4BshgOeqImPJZxtNDM8elusDUxYyQwyevZ3/P+DgoviXWEBWaA56wpb
DL3LN3Z7Qi8hCLREbh+r0ZomC4x44A055VPfaZCzAA5fhbfpKvIBPu+/TIOsAD7/
BED+ciI84cwIN7gx7FNo5Q==
`protect END_PROTECTED
