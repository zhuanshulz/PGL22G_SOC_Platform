`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8dn2RlEcA7U+3jGp5GqqGwHrL6fy+unMnFSQewAQf69jW0269n9EhsQ3Z4HYB2xR
7FPVpdDVZ2TccP2lf7sOO85ebvG8Umi+FEbR9kdHyVgybMe4iFAYE3Iuo5lYpoT5
Sp9nOygXA4Mz+PCiUsfnu9B7GmIaSylYPC4unMZ9L+DaPbdQ77roSTPJyc9tfKWu
ahdmu66ehIZpOrgihMwhnNAX0L+iPNwpZXTBgVaQG+y+Y89ZXNMfkmWvc4b4Tp0l
X7IcLx3QY6SYG9VzTiqEEQcScMU6cny8jRRdaHlzfhv9WUU5gcC0/acoJgGfq8P1
zNPAUX81rONMCZhMXqTKHDZTPb1h31dytkvFXAORmhI+ZIv7xyMu4+tp3FIz7JKO
rKTM64aq8oADY5BBXL1fX1B+NyQ9dmss22V0NpqgqH0r/vsiDs84azsz0RrxmO8r
PYzpOsyQE+oQ6arvDS5KtVZVd2ezreNw1pi/8SQmyNfPl/H8aC58F/w2qu+7Ft2U
KZWMozmYfUtg7l+8XJc9PdvoH5tFWR02ml0+uqXSKeNGw3LJq4GB6VnpKwQdHEU0
XSzHuRqRNIM3+zLZ7GbfByNjFFbq9dHRBTE7H69Bmo9wO50qLa3ZarfyNrQ5RIjj
54zlE/QeX1xs7SfGMa+zFkAFHUlxfHfgP2gIHzufow0Ubg2mkzXm4ONvVuHF6CEp
4V8VI0Rw6xbBraW+oKM4e7kZ0Ln6WoEbvvBlHUl81HJ22dRYgGIbrw8kdVQMGhef
amI1kQGn448kmlnKASLg8mr/I7qdXq6lY1jGAnGE3rub/c/BG8jb8Iql21f97Bcr
nH0AgUOkyGcC0mtNiYLVMpiw6MHmJb3M6Xzhf+j5wizfnLXDOg+QHbOqiIYr0JwE
BxqlmQpWr0zE1YldehYJje11eAJptuRBaV/1DbasBqLxk5EdtZ6EDEkCeKYrTqG7
Y6IaOrPbHa17gZ+hKV1yaXNjMu1i2SU+oMPFhUN7yLt+AyuCDS+sBo6sGJgN3CpE
R8IRd22DM/u+EjqL1fCDN2gf3oczlqTvuVgQtG6HmEg3K0D4Mx3Kf+PX1FfzXksT
DM+qWoi6WYTPJsk67EHfVCM81rewSuEBiSlL9drXTmelYmuHPMEz7zKUUfSPVeWS
oAjkslGKYYfbK5jFMx8v9YETbSmIIyFsuJqsFN5o4frXU5+vkxaslI+uCbikZYNC
exbsjrdGTCJUV6O3dOprBqfIwkA2nfj8lXL8OQMajNWUtwbD5pKoicrstxaJQQ+/
KvBEC8DrTaKR6Nobm0zI1kK6w27plcHG7fwVcHTnu30BtfG25pqtQEF+w3/WbD6J
T7ix5+WYJjPCWTRmE98Pw7/4LdFgMAIDH6gWapvrrAx6EyQQdWFDJHV6v2VwSvkR
pfQ3zyti22Dx6dfX0j4fPbRF29qRcwqcj27rLYh4usETqArjT8KiCr+9ieLp8U67
n6487fpt+IGF/VGVngVN1SwJ8roW4o2ShfiUwJpQxrZOYB+vbGR25/wdwBMKSEuW
JKL/caF/hpD6PR1aI03MCMDPHjzAGtWb8VnM314TzCmyHaxCOiVs3eEh9V1gssya
k1q52tf/Qq67ZE+yElc5an2gUx9pLN0jWH07n7A4cIIUkqnQ1wlkERfuzCRuoyqm
Dnnj4Y4aMlbeK0WakKS3Ni4+XiR/XeorHTQx2lucW03I9BjY1X3+f199PuD2qvRZ
r7OUYDEhr+TTHhHLUaLZWovwK2UFoVmvIklunu9mqpQy2ARB7GRTEgLTrONrwjgJ
z1s6WTQtuo+5ydwnQunjtgFVJO9fS653Bthpq5mQjltFRUF8to9ZYS++pBzgSri0
rTKmDy7D+0nrZLokkYW++GOnhb3N5XlsVQ0WPQYH1OH8KTusojYV1QbRIh7JNpx2
lfV4jQuFQPX2jDNCQ2ABSx28HgNVkfA+UusZES1U5y0FN3dAWRMflVc/97U0bW8/
m6T5iwaeQrG6Swmz9nHZn5b+ZXXu6kFXlXFZYzP8o3dmjDV+ko+JMOO5Maay0J8D
UHKgclWOD3h/46NSH05k79jhY4oxn1FYTf9WGbLanPnFqo7cvBFuQH2RHDkWoteN
3lAvJajkWFFB5Qw2P/Qk3HHo+bzf1OwpyfIY4TxbKQkPp/W3rSTuQ658AuhFb/6P
o6Nw2v0eYDF8U4KUcC/3wqi48/k64WWE0RAaZ19PaMIgNBcdvAYaiiwreQHAoqzm
1MpG7IWPe63yzpoaSZLuaqjL1Bwvl2HsElDH3jmvhtrCTdqEO3Pc4/j0ttnhg7V+
edtSS+Zs4fJRANQggK0FY4sQV41ghCS1bGaIM/XLDhCBTJptUubu975aq4308K5t
bKYVQcv/wgf2aXdBBsFZhDw2kUv5d5njqxWIgRu6oJCvDw3w1hO2uJXjOry7ZUOY
0W9kXHsSCavKecwLCSPW+cB0GIWk3tiAl955Bo4KByWWOksh506Y4GFVEVEKL92S
hsXT2/1O1Ay6pubZ2vMBrKH9mEUv2M2kSHS/AVWLVpOtKU+59ywUGfHeNzbMzQtH
aqwPbwCq4j533m7D4n0+3URmkCjujwbiQYVY/2tfmfIzZ2FVOgISo1VFwftIJLwf
KAXSqV+ecB1cux8Nj+7h11lCeXjjtHP3wbFx6GYmrdgbf+ViaPA1MpsyTrd+EO7R
vGWaPoWZ67OliLoIhOQslFoInLvRpVggm3fjVgWQV1Lb2B5+Xe6Mcc+DpmEaIXcI
TBrUyOzxsbGPGYibRuiugLHm9q7COAXHpu1uk8KTYjOGr57RU1+NR8OuYZ8hWdIB
u30Uc/ArBxC1b/xwVpvFx9l2/oRSP/4dC7pcqtssnrOBh+o3J7A+e36qr73PIQVz
5Dyy9jK1a5/7SCp4yNrq9mtDhk7HEUc3n2SJ1h0UHktbaGF7XYSjDw+C8j+Z1u3C
orJHOmrx+fH8ApSpDGF9KNXh4nF5uvdIWl/XhE6sOC/xh5C1AU++fxXap5TI8CRy
0zHhw3ugFgv4qrGmWhINRLBbWaWjZvBK29iIDaSK381MdpFHmJMiDCJCAUn1LVu1
qDt9TLU+11YhUD6kDOnKopM9eQyms8f+jdPvs0VlM7qmDAOEvj4cyjz7wGzM1CVY
Z/2WXYTuDnHtMZATAirbEIl9v8qMycSVAVJRcYNlFxD0fe5HVox7Vg28t9bIagj1
zKkxDBAojeLwwtQQYVbTn6faMkj42yT0L8nMVNEicWRPVzSgpjpeehrdiYJQnP8L
4hoJEr6I20HwA0AIhisR8myhaa37mrBL86xpTobSXSbsD6uNBh8XkeAAIVx3NlA3
PeodvWrHUIYXdbNRwKuMTY2s5D/PYitGLV4aAqXOvUNCrLdybDC99cDwEev6yPnY
t36XXBM3eRwij6rJudsbrqWmo2/h2nLqX3QUZCSGnPbX3XBhGlLaglViZh3vis+4
g6y65cJt5Q8Taz5M4z8yHZlFvroWIDhA8MAOGO9JC3dskiz9NgWW1OiqT1+zjgmr
a5rM5B0se4x6nF3ihlr3jfWEFx5XzS3HaRvzEugWgP6G2Hw2+ugNrRTamBZsA439
tRI3o+S6yyPzVi2QnV2HhIc6F0ldPmgMWvgWPUQ0aytej33B0ojPN7OX2LppMHIz
YYyze0JCovVX2AIWSiZb8U7sN/SvrOgdmQJlZL/ol7LL336E0SIufBpfsltXvecy
2e83U3YKcHm62gEX8Pb2zKrKToP3eLVsU/GG8JjJxR9E3BDDCOaWj+xxAGQpbf39
5efXP6I1oIkJxxomKYol5r4eLVowLVmdsS9vJ87cMpoD8GxxPnKm9BBEkEbanTl0
hIJrdk/c7gJ+20B5nW07xcGxK2fCrdKBQP5F3KDpVbVGc6LFqlsUlSR9wEtpwLgK
nZY+ntHToHVzkb7BrQW0EYigeRhQx7HB5odPWvJoR7xOgsU/9C5E+lT6CMwMLWOJ
ShzkuSXxl1LwEYQ6+Yyfyx8UjhspilaksEcQHAPUu7ppD8hTN8/ng8UUUbXIFu0b
51EEdv2p100YvTzJczMtF+uSj4+pUPV+B2sfclUwj9wX2H4uy7lMIx3ZWD03uUBi
EVqhWQgYTR3b5hPfhx615Db01/Tf+kosfdbrPw3Ae75G5D3swQc3r22PLw9VNS6R
woi+ysTp7wqS9fFzlHz28KD03ZdrZ8pLYtlyek0HJC9klwxm3Y7OoCuLaraFb6Wv
1+SBPaTuH8w3bOGqJUGaD6Cm5tj9lDQDuCOuNnsRkdAPDs5FDcC79cAC4ct3he8u
GeZqPsVbbtET8AXu537sbhY1ed4pzndZzb+EAmpn1ndgk5WbvgUE8OGGYhYaTCVz
tFDSkeTWAYvc3NxKBEvYDL6K7rfVlKIE6FKSPUuO4TdOLTOVhzK7VAYAh4r1QadF
Aoy2l2ow8epotzpn0qThm8i5kedplt7vj+7830dN3YNFQHNNaHsKIZ+KuTPXIWjF
wetLKp6SSaPj450FFTa6FGQVOmu2VhTM5EWrQ5ukWyBebswMZh125x/W/n+FFOaT
JLYQDQHf+hV360XRhCsThQ4Aj2tO7wSrnajw8B+yR1ywXMOuLiLz50enMCC59vRG
Md3UC8MLB/v+dZeo92ZBYJYajY+isNPOV/pDizYMLEgVZqlrAzrRSEPpb9eOz69q
PD/arERVHjI1frGCGv8YnjJKrfvm8Oc2SRfyj842MDb938Z6rYPbhBPrjngB3cwF
4YABICXw2x095pto/SYzWHgmNM5VLoKr385OZRCG9Ewu57o6cGhVhji6E+vtfd/g
F1c7TQ4c/I2FdsyJYB2cN9A+DlMtGqiHuctY46f/54blAvD536R+73GUAAtBLxR9
+6EnC5dNMxd8k3rHJ/2NP7CyTxPLBMzNcMzeNGXKt7m4rQ08OWrA9f9YgFjm4yBy
O7KfMryVZ1rJwHFMqKvh7L258eFP+vXin3CPJKu1At4TfqgbBQQyZ/SzQgGuNoUy
ucjxJttRWGQXD0voOBjT/7XW4E2iUDNw52hpN5XV4M3qBJoQUYH+/tqJp6rEhmR9
K+MtdpU5rRKNGhS18Tl+zbDsfC6Ft6IP9VhZxjXkFoMbOUWobnu+efq+5k+bhszZ
/SGdotHyQxHidqnvzqf1YGxqWVGLmE1fu5cb458gwoTSYV6heSsUL4jOw11Te3Gw
yXwhqzAS7qGn/IgelKOeI5mBLkZIRNUHjqlfenOvlMfe5ipCBaCI+zbLmNvgXENU
LJT2NGp01+sIDYkbgLhPwTmc8dxIKArEBiz46y/NhrcvlfGWZfgdpqQG3QprS6Nl
gfASPC7+jON+2Es7e0Hmt3yyWvjyWWA83l3YSh2XrRiXWzGHq3hPqmSoB0NejNJ+
5lKGdX8wrTcCmJktCvCdr6MvGTJKGAemPP4EnTzEaiUgVvkirrODdUlKO8P63Zk0
PXbKbxr3BqUKlwUy4vYyMXSLERN351L7wWQY+fctL3tQIbaEi0XmYAgsqn+qs3W3
Wlqny0rL1b7sA+GEE+O8sNLTBHlSH5KHyEKg4dTfZOvxZQ8Qxcq4ugsVLT8k9zuh
WdrmpH552nZ0ZmmuYxynVfsuNoW9doBPBU9RUVp3BRomzhxuMCDM7hPOZtAyMuyz
9QN/ZfBmaKv5BDZmR9XdcYaTGkNGJIxiC6M1Z823Z4dLH+GMhDxEuOVVYaecnxfN
1Uy3diwsLVfSATqNdg91e1t7UdXpPVC1enWleaU6tc8AteaM4slcgU7g1dfkXcUB
z1/8Urkqh5Xjw+RSHUStIO96ZbR18pGjj6bWTu8axtz3CvYIBI9n+rUIQpzrutgn
33PmReCaV0+jTfLeFddUoVLoLsTLt37AO8T2K73LDKLVlt1lx3RsXepHsNA17Jl9
/7uGkPm7W8Sf5IRmdt2eYRNZ+WXI5EDUMpR09ubjXOgWgVKi2snnNoo825ZvhkhU
HnOxGByf+a+d3pzrYlKFmo+D+9KouaeD+A6r/6xTeQKw1kxCf0sDJlqiQkLGbsmW
I3VheaM7XRlc3fJaPMNrEX0sceiDu5Dp3gXREpAxYKkGKcNYtMWm0z9vxvPgH5JR
z92jnNOGPIcThEAO/mYA4PwfKhZPf4xjakFLVd0T6fOS41+W5uWES0yluz7Nhr4p
hSgiCyz2DG6pWJTjCvvOCQiOkQkCE/Na0sVqzpYxufNhv1glJisCVGnr/b1txIfc
sBJgBBT4cZr+FAchXUpDotTiZWAyhXaofeqvIJkCEodHXSdb2PZ2YHYPU/7+jQlr
ZFl1IoTe/yg1wE/Y+TLpKWy2/GvlaTtg9REtnutJibLr6pZGsaMDn9q8mG7LFmBg
BiLdIbg66EMctmeakXKIsUkCfZjOVj++mJwtIVKUb6M+KAtEAlVwo8EaY81TU+WL
+pYwoia6IF5ZuZs8DKpwapKyDYPak8j23mI6lKIxqAE+0a0GXhYTvXHHS0x4lYt+
zCK3gZsszCrHwFk0bLknS2+poj72C3j39atAlWeWrB3F8j2a5s6z9MrH/OUR5vCJ
RzC4dsMN3wU7NW0pwnbIMNICKRfwKk6PD9CQ2sY0h/6Y9D6ojafrl/JYmVFFOEvN
Klds/yUhWOCD8B8Ey/1j+L3Kqz3/9KwtOMzbfpvJ2RdYfLFGv1hukxaiqrOKeZyn
cnjXK/y3b0EcycAcG3CA9n5J8aySdmbwQLn7JBCHfuqUsNtxcKUR2SrtdXare20A
vUI/nGU2y9Oen6POSn0YpaI+L+BYUj9GVHASUdliEMRqUND0lJUjl15prUUtzIaH
IKDAnjF92eShE+UPbJ0opAHRWEGA1lvehIxu3rhqqY8BTagpRK6EgVSL1sqc6PVx
M1TO4C2hdN/tHCgvOvHQA3sSWqDv2avPffU2hSX7V+w6NMMerdqu5/3wJfYpjCKc
IRXcEEd1sWygVCknYjKeBOkQUh+YTSqOnNpnSw3/2twmy9i2HVcSEnmnHzMt8vjS
XT6mjcG2RvB4i4mWCOJS2QVWCNbDx4wTYGSK+aDHyvbiyRYoWaauwFjp5vcaA03M
fGHKXT+c5VKN+bmJrbtVa8yN2jn1KXs+szCKeqkZW0uoIEDcZ2l5d4lyBCE1bOGG
AF+4HpH8CPpgN3hjxUYFDdR2nT1rJiLpAGgLjULLR2ScKVoP/P4pIV/6QSNqQmSl
jkXEc3CpqaqO15gYVDvVR4hXDIote4QW+03wTYjnCTy8ycuNsZATc5wYSM6gwNEU
xJJFnTMoGOofBkfbFhQ8Y5mkg3Y1Lp40MoQpCHynRvM7GNqlWLW/eUJcf/HuP4tu
ilEL55XOqsyDSC76IgB2JVu0MNg2UcGbBNLr4KarcnpkkHV/jFzjzIOJaEc5GyV5
Dkc6mpEQ4d0wF74z3cdy5feO9kROyNebOjib/DJx4NHAJMI6+lO2epuJZ4TcSfj1
WGsfpDiBurmpcFbCKWeJ5p8UkIN2akYW7AX3NmfvdH7V1uyJqe1W9RPhZAHsU2D3
9vkaRiBpSTPfldDNXCb2X5EZSs7uX2zf/DjCbgxuuZrpKEvvViOLKBu0457vLk1b
2liMNj8ZxAiIaAIM4YmB1tPCVAPUQ2oJ8tXBW72RYmwh366ot+r9quzigSi/Wcst
FJnHIIyzIeKmc0OIodyfgP3yb5NLI5IAoezg/eyMWB+aZuzuXcvhSJPX/wvP3nO8
YMyag+AfrfzDOP6gKgWodOlFiFwM0tkKwKUXT9P8MfL94papBhjNaWHYE0XM2ld8
iB9qqQFm+hEkS+5S/kGEPOkLE9HgMSaJpI2hmACyU7qqJcZVvXuRZse968WxvhLb
+mekItVoNjm5pN7gXtSfH30uxRYNTejnhe3bOXCd+3VOQEh9k/x8nci5igaqQkty
pRshEVkx3CJEl9PiyE37lHSkgSVH9+6c54lC+qbmDwyGNERB1AYqRxELZmmEPuOF
Vw+rYYjz3fsaDOYTPbRipKds3EkYQ6VAZva0S+pI2kSRWHdVWmq4IcjHoXq4Lekz
4YpPafCgdS6OOgMCS5laQ+10AOE6k4GW7ASLX+p9Ad+2nNnzB7MHvOFQOk3ruymV
vvAJvmV9nzIzclX6bnx/iD6w1Nx9UaH7GedqjUv8wZCxBcJNWuHW7/8gvqwC1Y8w
LZAS0IxZPJoO3TfgWM8th1mb2bbbdyH1UKa54lihtyNgANHfnguNRQdMqQwYyWDP
hMGG7isiTrDtt+FcscGeLoWUFE0yZUipYiwTwBNLXca0RmXv9M3mpe9gVU9hsfUy
W26UgybCesIXHd0KV+PAEtT9rsadDSgYHyr3+fbaQfEbFXA7Tw/mOY2xKwVXPr/m
1t61knBB8OANQGZZlKPPDoX6vMyFNP2KtlnK4aRCW5TGBqaKKZ397GM7yjNZwbme
cQP5MjZGxJ9jso4EWnj/xXFuc5k5csbNb+/Hp4vTOjOQfP5atLQuPVdgNIb2iNZo
F1nKAkM+nJssS+JpQ8ywAaMFkayN67HXtzsDLl0YdL4jpd3gAnSq/eCNYwZ3E6zX
g1Vi2n6P5ni0pts3HupKStOENA+W/tQuOtsoq6VSDotzRckmc1X1jomQ82KwcZ+c
RR7C8je90AwuKf40jCO+wyZ0HylARWq/gHxEkFxgjkm4I3KnmsuMzY0zUzBgD3nL
A4vsL1FmAJYT4aZVpE/nmZbvyp2k/MEzW3KrxEUPEl4ExAqaTWwUgtWAMyr39vbZ
BeuHu4RYaEsij5Hx6ZLR4kcK8r/z9RWozGSyJKnmvB011LGabsl0ILvceCTObDXu
maK4A/iERyYKu6SYWBEIRTh8NuFHRwgcFhLnTUmAP73RFM6IJOPyjxlaIeM63WTh
kVRi7POeHebKa2OrBPXMbLRqtaek5LUgbMe0GMKjfbuP4zA5Xxf+WaXqCiuNHD0z
uGzCKJdfDDh4cS3LWSFuLwFP0Q+Ae1Mst9NHoZU2kniGEVg8PO//ynY23YOeOR3k
2tk5S0WYtCvvG3FuJjhRNszIWNIHqctXQcPvxZCstX67BN+eD+qtqfxBQkAeQGLW
fH6BRPdLUAw3PISKqee1Ye26ObbfOW6lKskiQCZevxSBpR+B9joWqsajSUkSglyQ
O9HcoIWhl8uEr/hl1kBwvNxAYF5tx9vXrDPXBpaqyx860kZxvfU+Pie5fsffrdvi
Frxvgsg7R2SEYy3pDtg6ieoBgbat3NBdlQXIKv45Q4rspz2mqvABxsOcgIHoLNXm
MOztcf/DH5BTmg95P4maKlK0aW8pdr1VTfME+224mCKsS51ED+cEFHLf/Vb8a01d
RS7lcXuWu1Vv3dpf9WdEMi9Pve/2gSsRUihHTaglEqDFjndlX52ogGtINuNVtYCN
+SyrhAZD/NH1FPYoNWOCy+qsUfwEtJSyX4slmfa8JgV0YlqMgU56ZsefEei8zteX
d4sUisYpjFc4dJk0F7w5Fr/ZSglCrUZTguC6l1EM6BKjvkZfvDySG6tKOgyZdg8y
K3WtdihMimWg6GllFfGg1pngp1xntA7GXh2vwizGeRrhtzIVoyQqy/La120r2Jbn
XNNYiZoJjRrsGUJ6IG+jzKr6L79sgvda8yxzJNyPw78BxzfAwCf5NQfCvqq9wpvp
myUE/ysVsyafqKyvH6M5u0uOmCy0a3ebWBEUWWKnH6OLWgyA4EfySXsAiXDqKpQK
EUKIPtwF9DRMEWndgtaG6mffvzsE/EeutYRqfDO9RMKJsXb5oSI+2QOO9BQxJpSU
Mjs0TOH8f7v9KWvIlodDinycTjmWcqDPUQ8xgMpwIrmV0loqtV+KKKICeQQhG6EI
c0gUSXY0zxosqnEUot4L16atd5DEx3ZscQMzrZ1qZeka1yFBuZOKMfM7NvnJsF9M
ay3kZaNiCMgo7HcyyClN8TbQtcKo52c3O6IT9TPSK5/lsDtm3ysDuIJWmfXAlEIN
OJfS94ZiPQbiKhUO/FeafC+Vln4vLkWWyUGocorQh6VsyluBF8NOSD55bOa0cfmO
wK90fQHRYiQWY5wPfzVD5Lghdq3wznl7ghSztvZPaSMxIVktqeNWZrc3Ho4oY1pu
lnumGsG83hbx6jdWIXYX6512BCsexF1b2emWQ5ueGAtlDBCE3ufIg6pF9zl6ETSj
RXn9XIJLQcWLb4AWhuuagyBeh4eWkz6mbmIOMFv8W2jE4y9vQHvU9nIiFC/wC5Rc
7/wYkYlbP3mpep6hNYAa44SY8633DJ7xfEZiTc/MNr4vkZ/3KPCHCCuWRERZgKJ3
Sy82TTNNAuhqucd35VvtFnH01bcpYyYUlJdIyC3Lx4VP1cnMjPcxtH18+CaCQlKM
d3XDhq3a2P8wgD9NV97KpRd20fTO1PLmfyGpCg9Aflo9KIJM4JbDuy7gxJ14i8kH
t5M0LvdYmi134XtcwcndnhTUKyIZUAOO48MFY1p/Ki5nHa4MOCfETcBRliqFSYdt
DcYceLAiALXXsGi+AVGZ+47gTmSBzP2ueyn9Kpwg8t8Q2iEn+tCygIwnhiNj4mnQ
c4O5a4vXQlzrKTjvdqvY212DO0xjdv0hZnFj9QheAW8bg8nupu4iHAMoVxqjsTTg
Ie5i7ELLZJ9wfblpMkx/pltBda1IEBFS2nXNtsjkQXRBlaCRS/3YC8qj1E9jgLHu
gDGwgNTR1tq4daFIuyuLdW8l+XI2ksnA5Ak2dmI5w/ZMK62ra3EEsU+tOUG6Z41T
owiOgSx9OwOTsBoZbOJ9ZuW+TAAqXkKr1RT5cgvfIX7Q++vQ715bMm+LV+NfD0jA
GYbnqJoVcAhQfiRiOz1jNdrNovS4tnReGPacwPWhUR8uQU4QnGDPUV3V/gnB7wtz
kLmbD3TIrdx9bYP08BsGfw9CH/kDxggKrhzpbx675aXaaM1CpEtF3uw2Vk2nhT55
oR8WEkYgaLUHP6rUi3Fago1mnis5kN2WQrXZhhmMyDHf4d3FCCfWDur4rFJBV6C9
0lJLYEE8z3MYTvAGdRssl3rBniZBJmaXKxo/m4e2KjEB5yO5ESQ1SkceLPuSJVJe
OaqUyqH/QDY9c/OJZPC4E6Xot7SDtGItfFs045DAQtOb+X/zgasn1hyd9iA1NuAy
4mG6VXGSzQPRQGteC+uCFTKomZww/eMjsqBSQSXHNJ89B4DD++EiVClw/quj/mp0
dbq+OV88b1hv3awnI8A++d6kTf8Hl3HJPhYoafNYeO4IJ1GBGJpTW8lRZaygKBra
7SWdkiTNcuS3i5WOgPZvWl1O3VCviJ+ETpzWyaaDxp53XGgPc1bYPopb9OkyBeDf
EYkkuSwZZ8CvQQYvtj8aG3kuaw8xStGr9Ud3n4ctCHF0QglaLJr8x6dX2szWiFrK
52ZCmkKuyMTwsaL0141MTfY9z9Bji1SMzR05XN9bdA/9uuakwLyeihF9WSA+AvZ5
4KGQYtbmKTTahLK7OsYtLsDleKavP3P/KzjwN+OmPuGw5SnoBAujDJFW4TiK1rtr
ukfQ9WfocDH9IKnN065WIQ78Wxv5juXGZjzf5IYT2yh0Kc8UMAJ9MGEnmxYN4QW1
1Rg77dyUe8HaAJrxxQ85Heb0YN9SDg+sRHX9ez7I62x9Ixb2rdZ7UQbJIdj+zpW7
RiTI7c90+rAMyXmDhgBkxP0c5Sei743c9a+510EHFdu5FIYMdiduHPO/GEBDJxVF
G8jDVaT6fIcGreqO1ZtawwX9+mgGgxB6l9tHmNJvCuARuiuUxooo8N9WurdM+/Dd
run8cBbFKf6+71ENcZbnN1jAzM/SK4jSC4EQiTzDZrOEgKxbYDZw0ONc+iMYgCoc
HiYlE0QQZ23vzffwAvCe5nwidg8e+pGzBVmjszwt7sl0Ior4I5Cwm9jop44LKInD
oVUkM+PWmKtjwAdmrsVyvU7fIs9//ByUUOGW72UTxl3w08NFRPZTi0luhYNuXpjA
YnFGLtNME1yRL8/Z1KDzCfhN0x4iyZ77SPeB+fv3S/uoTLJtReNiabggiWH8eSmo
mEtyyrEJGhU2NCtAFfUuXTsphXTiWCSJU6mXDxQgzH/kVkKx7NHvBAw846wQSj+8
PoRVV2z43+P3Bchx9wLDR1UO/NYhk63XIAVwlOOYwhVVlJdI97INJlKUuAW/0bQ4
RvRALTfr4R9qT35eXkxszPPdy8l0GljMhvTBU8nIR4mQjXrf0X6B1rCQukrrTKBp
WQ9iY4G8uRjrvbPukjxXnSB/9WHMrsvroB+9Fv51UY6IpCBa9ds2C5ZJyxi/m8Uz
KedOhTcUulNC1qJYwWtBqcOYbyo2xT2i/uHiKPBk7buVb3c+AokYU0Xvqw8KaUaJ
0EqpEVPJMZ7qFDGmnlTDgxc7ByaGELiFTul/x1WoruxyW8nwmj4exKLZD+OblFgQ
AKVMTGF+NIa7TCxCPhCU0rF0/Q+dstwnDQGbuyDHin6X8zqXUyYnD+dXs98Jaw73
byN5itMKI7V+SGWPTz3Hx9RQTjbXk/3N/vaGRMBw2tDkz1lQ4xoPE2hI6MiFw0M+
yPYRXxfvLgzER+8L21WjnwPmVWSORJBZaugqzPGcwOT4VaqBVELg79p4ONq8x3g1
5PGTIoqPweT7RoqESN2cFWXWL+lrX3ucfH3BV0P5+nFqwUGQP/JY5XIid1X2+c2r
dn4ALudMIsVQfPUpk131j3z8j2RDjRJncf3GBBVe6dm2vRiqT+QzF0tsDj4PC8YE
VhxFvzrY2x2LjdxAOPURNU/KHX36zfD5CgkyYAl/wAFoTNCqLulVpytsGRzLKNYl
mjPe8xwWuDmOjun1xZCDusddfWOuc5dOBqWEVgWwg99+nd98vvIoyzH4SVtNmkKv
6oA5lSTTh28liUZNymJNqlB622IGrA/gdYnU/rpya1bR9Al4H1DxI0DaDymp8vJH
RgJCOSSFAFud5F0c2GwP4+VjjHPPswl1AixU6hVY3OGudeOYRanOgAZ5/8hoMXba
888g7g0vVIjo9fuhrlsDELK14Ha8jvjR/pi2DpIlsKwhIqdCTumm4x/0zMbuiufN
gRV1ZoIeEWAziO3qpB4//T/OpqDwHqEtFCXveo4sWnd6jF4Ah93kd84LHq+W7y4t
mGl/tT7auaNF9Xi39l/RfVRY+3Dk4HlFgxx6FO3INtCVz0CN470QRtT0s57/obzk
9yvl34kbiuudm15uYLSMyBVZymtQVSQAKeXr11oTu4cv2tWfQMZllWPG0QJY+u+0
v+AbfgQliRzJTJqHavGRVKuXCjcbiWO5aGFR34zwFrMwbA2d88Bv9Quiig1wSh6I
u93P3H53+sxsr2oMROeBSlPFVb/pkQb3T+cyLhJE8LoLateFo/xyaY6R+LuEeuZX
7iYoVErhkNU8SbvMjizRERtXmkmlXr/TE3u3QkdRaRNI7gtzlomCwmT5YkXKogQy
/HxIz9mJlHnWQD9tCJnVYbaq1hud3umg1TIv7m1CxYC4Q2HSW2RVSWQ1YQD8PUYf
C0e2dQZqVzJJ8gXY0EZwqegOStFYl4UYtkRC0UUGNYUl+mhHSPlzpBvAdcYf336r
kjLCEZTBg3AQje+ymsPcSlEArtZ8/TO0iaHuhZ1a18C+KcpuYP0blU3KaMNy1oCP
JudXCbCwZImvgRwgFsZ3FW9B9IR1h7/SHyhjRcs4Utel3D8o8+FJInkVbkgUkxtk
t0HI5MIYcxPaHtaSuWVQEKNY3jke/ctNHmqYxMvdhGgCTMUy0QlbiuQ2Uqa4wqRH
CQjKU3Nr8jLRd7IlxGkuIAFttIX4zvC3s6IIwxNkq8v10XytQOcbxqrq3qBCoSug
jdCaxhKDYj06IsP2vF/6K/tFu7Al3PhSxN5sVT9YgOMfbKlMT2sMfT5kZALpBbxd
0TJeGzj0o875x8IQGLTnvi/hb0ddmsuvzEwrhCeHIfW/K+E213+NdJbGH1EWgNBv
WHoW2i3TdEZeNbR8ra3sG8rzSO+V+b2b+y6uL5QCJvmZytHroBEyMAjqDcoaJ4c5
9W0J8D3XlsjPGqMl8Ux1Vo3rNq5XMUVRK2bNpS2co/FHwAAIrxe1BfXEbTXQwyCV
80I4BaXKU3Kn1WTfLBARGCUfRg4OgKahx5nMyzRqwpeaNE/qHt0wIcrI4Z52paEl
BKHIYAA/wEo/MitvfLdrOJh7HExG6obm5EGrNkjR5yVwx9YmwSJu0VH0hYfy/8c1
+q84fD1M+0vw6IQvLhbQ84FbAJ4IX9GQO+JQ6u68EME2nwUYz4KsROerayC8zR/0
Xfrrcuy1TNcw9mXDrtJuBCoEJbQw8VYnHWD11f5WSbabo0efLWdfgXjprRmHvqLe
G1xsVQliPm/g1UyTX5VQuf45hChrLmjNwtsF17xqpDNzUosEeOkbT8g7DL6FtV6L
WeCfyB7iIestYolvmXiZDP8OuFnCP7hQu9NQnKO2/17erFmARsqHWx1mTzjZ/N+e
1nm0qK1wMwOaoF3ez++KUeFMYwSdcQwOqtth76wNB2zApM/6AL/XwVEvFMHAOsjl
L8l91Ymw1is6YBR0weT8aUJXTNTWd4npmkBdi7arHf++VEaN/wieJ60Lw4iJhSCn
gC93MrSKu/E0XH91ebe2joCaf2MgGlTi6e9MY9/oMqUDBSpM5FDJy0+hJXuWBWyc
4xw9N1eHOiTrwwpxdD0p+sHD1oshdOdc5FZMy4ciAOrz9cXWmfXox9jOGy+MI2b1
WeZqnu1XNk6+DVyE44Sy0RNalOoKCB/OKJnTwDEROTw4RoBAj+QSMGQ0EqXLawVT
3GrCmOjoUSfSN3oFJ/BrRwRTSK9USpUazgs6qQDKxAoHtmhlKWXV3RUvbDv3SKYo
mv5/2apgT0tR/mdOpnI0ojX95CNkPofNLZcyWHG+oWNf+NsPLcXdLm/0CFJ6yQLg
8wpYZm6vt+txUS2GUZ9/4YHw8WpeUQbuD2nX2jfFenmp4ObC+DVF4rm4k9OBtovo
YEwwQ8CXNkzziIAVguIVnyBk9YiEZ5FXllkOiOsWbIwSxTUuXCj2CPxLuJ6nAxdc
z+3dUEUiJkTHKYTYbhA9wHYztwcK6ucfkpF3Zv72tGk4UrWzSbFRbAPgJo4jG4Bz
JZo+TVjRzImyXXqyIkN5d4as+IP1qIOuGngviqGEfLjMj0ebc2ukMKna+1XlA8V3
1I8wQkMkh8QB8zwgT7j7uexpDyHdITebQjTynE0XNifssqXUuH7Vr9fhPV//bG+4
VGbj2g8lDx0i9/JSNg8J292c+CSuke6986FaLc06peoB/etg77WN0fMXGp+4FOuh
coQewkFraPOBAeHOn8bYYGpOdyI18EeZ2dk19erf8VCjBfAl1hrS5vdUVwAxVqeQ
0gnx4QYe+d9Ybsl7TDkQBcUfETFjP9pHt7hZh3K5C0amTJ30biZdYsRw35O6dtRX
KsH3OrTWFbt2eo8XCPFtpeUKJSJmqybD5P/5udswHD7CGEzzQLw8H4lBr7jGiftZ
yQLCV6+v+zvqu+0V32rurfjSWMEg6CglYtuFlPPNnfBHibK5u5Dbp9nSbMaeX5Uv
QnZxCIa7ecYs4mb0JWnYA/52OJx+qD7LYIquSeeFej/2kBMwnSGmNOyNfv7I8e4g
/rXpo3uB5JOSURp6nhtpWFOCfztKaQ/XH9c23FbmiwyVl3QVf82ibEe57ZhGx9fH
EBlm0BbdclrjD3H7urTndAneaY8ZYcKXZd4qm7oQKbCHUyvK5V8Zjn3WV/n9fGAg
fHnSWHjPvOM9Q1xmDahoe2msZO4fbaZT+4LuVGKOzx6uXJIICSz3DyENqsedKUgj
vgffslmdavbi+UILAdqTRGuVQw63262jhFvyCRA42PW2dquiYutDnEc8Th8xMxWS
DtuDKBwjegBwqDXWMJGZAFn5eAcKIwYurybvBIt8WZjmXPunHhk2j2+9ZaQLbeSM
wDB6VeHTCxyjgiOug8pLLtX9dVXPD1Fni8yqaHLl/3ytGKi+6cfrsSv5eNtK4CRY
dCqeZ7TWv8g3W1L8av+LFA/cuzJIaMnnWtW63W0/fYlN8mdcy0ct9mqX+Db32NJc
t7AJhU8wu/a9ZwJEiYvDBD2vSJ/pU4eiSp1HWB4tOt+8H5gsVZcok4X94g+q/NhU
sT4Nif0IOkDalFsRVUkJ2q4hnS0BFfx7M/F0U1qlH439xLDDnZAMNEdzFrbxIPTd
cib8fLzGTNWVdk/2KpUWxeyAQ7aKZDR4YH/hWXQPZb23GcrfIcBktkYRGho1r2bQ
zYqLJHeGLLQSEo8dHCucVpO+of+jkZYXJbPtS7f+PBeZ2y8HYfncevkZe2gbHSlF
zZFSVhKmA5LMsBI7kkCbYEqxMFpiLIuq0YYKwzUB9b+XYnZtIb6trAszB3UODAFx
e0UP2jrgTeEkK8JD7kmrvgzmPMr7FJ7D6+SlUkb6V3zNjMaFPQ5sjkbufHgeB3Pu
0wBNmleskoVaXrygg5T+Db5PfqhXS5kfchw8B/TPMPoTRYG/7Hmy4UJ2BjhAINYG
jgC9UXxEOhOxWQhaO6PmcZw7ef8h2l/rCs3GfghRpq/HbbDVai8VrLz99AgVPFvR
w+4m23EuOOY91KUjiS9GlYFvA+R6Qq5SA1bBC5ggFakW1yPK7vkXUx/N/eBWRMBT
E6i9EfMj9pyZbZtaaUcFI9a19s6k3Gn1AR3iByuG+RQIAd9k9q4YVXUXPMJ3WAgP
h/bQLc95sqiypMCnbiqVpBDog2WRX4adhdrfe7nY6mqIMbfl4rYKbJ5Wdp74T6Xz
QNzWS1p0tlUX48B7KF+IKsiDkOU2qHElWOGiNtgv5R0mgsJmIR32a953VorTI+Y8
Mkv1HgfDR3FNxBAl6Dl4uM8QFNxeyO/9BKZum/IEdfE2XElVvnQ6vGy6/yv0dRJO
7RFecHI+NUt4mzbIUSPHhdWl7gTypAnBk/+PVVuDqTnyR6iIJF8WnXlpSghwCyHi
4i9VvrdCxSR68s/VegKWo0wGtQYm74iC+brzjnE+mOIN9wrwOc18KHqat3PA3onu
kqGNwCy71VlzutCQyr7EkH/9dUPeb6gZ1UzhAEuTObJjShi4+AdLrvHdiMw7EmkA
bEK15xCG4suBxjpbk4D/PyqB2hGMY8honkQ19I2qFFfGb94qSmqOfCu3hjreO92Z
MhznIp2kM/saExCiiAD/7TiqDYF4yGyTt3cneegQuRA0daBtX1Ioc6C6qDs4P2y/
ETewnE/dt8YCCPZXo/dnhlyZJSoyg6IEnXl9OM8zNFGrZ2qQndlqLoVezdyr+sxK
AsgbPfzL5VY4sgjToxx+YShOCOyP68KgVZ00jLvh0WWgeKqYMmGu7aKezPmA9K89
mLHv2cbahtr3XHdBdm6a/Aaq3/K5LURae23lPjkIjaMKCnaKAPjHr9A0PQvvYWO9
hZEvRtCc/t7ZPUPvtjmnBiEf4S9DhkjRMeY42BQxkQrJfcdyGPkaDmvf5W5yg4GM
+5eR0rswuKb7j6kVtrq8FKmXOOBhJIkknLVvmuMonrerf1gVODh2Y9GfqUgd6plC
XSgwKL3KuEypkMHMrHXjY9asFSd+ErMW+enBgvWihCStXOALtFeTTWk2+eAyiOhv
ZJtOEsj5/cX9tVbQJJ4YQ5YJDPTdII6ROHTiMzrZp2ntgnUEPxxhYMy6BP0Iy23T
4N4TB1k1MNC5KqNnNyoIKzjacUMdRjz+ERvRi3nu4wDyj+vbG2p4uw042cdiB3yz
Vf3lyU2qdpoZJCNqhw0z2ED7N/Sy8X7srJFv39YIeMWWbSlWIDs1pr6E3v0sfF5t
JJZTabMg+Cf4xbhdSFFBbpJnqq3GaZTELXsgtG6PAyGD5C1a90ZYcSXMlu06d4j7
b+ixnzTYs540qDJ65bXbUq5LDmXulR5AOwVluIkrVTD68AfFRrYGKIEoyRZL4nZ4
WUPoNGqCUNf4z8gMv/k3o2ZXzbiIDyHmEYJvJPsy3dLH8P/SVZUoidp9eqzCknzW
PDF7qSDhJq4lAJXiaC8xgUWpHsthgIpUVkEBKkVX6nCO6lvV1z10dIXsXzbLWElT
J0QfI7o5L+iXcQKw5NlYFCaGCegUaCduDeR7llVIJjtFj4q3UkTNZ0Vatzv0B8U1
XpED9Eqdacb/c9C45eQMfACQO0PmQsIu879RwP8d4z0BgIXfcWgu+Zlo2kot7fz3
mHN+lsDozwI84CIabWWkqfMMN+dqo9rvXdtY9/DHZ141q4rhy/j86OFy6ER+cVvI
7qeQjHG683NzqZ0c4KehbJ/53+Iqfqrf3S6RkgcHE6G3vRJgsIzjDwhpUR6cw8JQ
xgpwDN9Cnvm736XMO4P6/aouytMBkwndIv6DPKBR8Ki4WoSQ/g28YeHlUkH5159W
3yPzaJ1kDrhUN6Rs3+ARbQCo7FSeZ9ZxgWKCSLBNlRjJ0PU1YtJCLa85CnCb6bMm
Bvd/ihPHZaP5KUzO25iJLZFCsakaopSGYk9RpQx0IomBWXw2D3u1CFFAK7N/ioTf
kAORL5dsu/XBZJzSyijaYvwh6myYOFRm300Gwr7n1GXf00lz2YBVaOWp8YjzqLug
8et9biT3Q5/H/NBaYhxqHVyjqiMLJ8M+3ZV7IvrwjI0MDczTjYR6otDVzER6aLoC
XlDttyN4uNqu0CPEQVVVv1+ky6lfUK5Rc5VXAbGu3lxmaLhZoH1+svBapJWM1MGh
8mlEVTVV82pP2yd8Z5L9byjHlTTYXUNbzRg6BHXEa//hFI0utu2UAvjtYdf5etUj
BNag+JIlkFkseRtcPF9n+SNN29DMjQ3li5y55mt9/djT1lcQ7Ijs/Qha5sMH5kSi
c+SUOsjMgr504uvZuPwZ/4cc5uqKVAVZc12CGNdIRDv8lzW++f8MbWMPxbutvF7n
HulZvK6bWCXAnHJoYbaP5xkDTUVAnyCdhF8v4ZbKJ2U8lYMcC2l82P/xJPG5WsbA
YSpRS8Bu/Qyokv/OdmJOZ0PG+mzQX8htCmfVDHlC1SudLwrhDxKRTGr02EeMPBXK
cTYqZshCSDJ1uJImuHA0Eq5q6tRnm4XQo957loaNESP5YeCmWxFsNLksTJHO1XCZ
ozv5t5mcteE6rz1S3rL3hMkqIiyYSWLvv77E1kH4oMX4MgB0ST6Kx7kVjT0a0JHp
94k61Vyq3StF6nMvo/a0EYZmT+OYHGuJYlwUEfDcQn5JB1kkchvKBJHHOfQHauyy
4KWCpIJvwWSZT28OdghqJZlHl7CQp86NKwwTlsNL9H9pI5mijt00Afy53aZ9s3g/
eIHpZ8kAXI7VqhmjeCffpNyWNkxulsWguTgtM97t153aK/oS9TQT8W+Hy09fLcuv
XBZt7ICy9BwAUPktWZxlrTxt/vRqmSLALiBzgEYoKSx3gIibmhPs1iGKBBk2jRIM
bQ6tsTzM+ns1DVNqB9+IJ2aycuboVYN+CjjnVc2bhsY3TqGCIM0EaxQKNjD3mvqg
wwRtTnX400D9s5tcC6tREQHbctvwgODspE7vVn/PMXNLATHaiBqjY4s7C/qaJJhU
Qaf5GK+bWQorlyTBbywsi5bbEYMRFmsdlcPprMjgRGCOHVdPVmpf1ZlcBLfRN2Ho
xNfNaur11mekfWNQcq66NXZ1GA2PbryhKSpnLkxjeJxLI8LKARDtxUk7HrAe5eVN
xm4tmJue2UlkpVH+YDSA2gAsNC12cg5qwmRojJ414moOe4C9aqFFDd4H4YjbwH/i
M/9flL6D48SZFZGVp473Y82H4j+QbkmoV2cBmx1o/wxEdAht3rMjSWt2V+yi1LSp
Hzj+FdNPzd7ike2jKLw+sN/E3xge0cTIkinPlT9tNMLWkRXfbQYojimc8yETM/zg
Z93m/8vO9Jv1ON68vJsQYfbvcujM7e28ZoerBAAWcj3SRPGwptkoxQLqJiD7z10P
PKlgeHgkwyxsyR/vBbZ9nl7+EGE+bt2UE2qpAHso9NQ8qxUpnaik8RsFSQiXPYk1
+QAqLql81nfejra/7L9pZoPx1vtldQ6Ms1SRCA7NYMvC6l4hKkfE7bGxwc5NEu+h
A2dWRjYXzxmG5wR6yCSIOh9kIsxC6VIWTN254Ak8p6/mDEKoPQfQjRG8/jAEp+0/
zi0V/zw+k9FAbGjtL7JryTcMjIpomn5J5LPmaEqwhayN1jPjwCYWSEBet3EmPaq8
+I7GrKSMBPJQ+MyCI7sd7S4w/yG6JQ7QH3BwQXsFYGW5Xzi6nUDz1n5JYOrZ+YoX
5Alw2ehQ9wko5tU7t7BXvcv8TSFEhhSZ8mpSpX/oFYcF2E90SWhmGBTo+PVaFopG
5nsgXoSAuXgLp5Kc6//6vK4FWjrk1SfEwsCtyYkDLBFbcWpYoyHhqT0eI8AbuNFp
AB859mMJAEzN4AlEQvmiz8mY1i79V7r/lHZbUBvdUpsMoq7dilca8Qkusq8Ui8qT
Z28Oum02DyKzUeNuDds8VxXxbDRf12wqOHAAzD7eyE7T9egKVeJu/whef75WfbOi
GF7Z3Aym6aUqb2AVupiA2DffWC5UJ74y7K/InF8iM1N8jt5CQhTiMjl+FNBA0hoS
USQMESXFeiPi8yyyZJhsnkCZ5HnJbQAsgXQuy3jGfLSO8fwvUk0EvlB9N5KvxZdl
op6PSrEazf2UV2UCLv/a06UMkQ4HyB9ZsRw57sUOK0V9ITv48r/Tw/ompJ2ATTvT
wml39QwjzVdSveWvpuVnKLUlok9ZK1LcSYry4qowXQeuiTcEP7dJ3oULIAA+UZA5
6B0Kn1d/r0sZ6Jn9EUdQk0BvECKIj2YAQXoRIc4IUU1cDwNUsDVCDWYtbtFDQLJU
FclK9Rn1HTruEQ+hYAA7fUidDTi0E32c5Van0GDqnJWvcu6Rc93tXybMUM/3D1ce
MD7oDTIrzlC4NNbgW3flaOcPEJoDVqHqVC0QYg/6W1Y+Nu+muGGshbzR5l8EMteI
4uuJfdNjovToLBQW/NTkyB0EgViOEkDBXn1a7/EUSh8ftPOM3fIefirN+rN6Keuh
HuNlPRVfglVwB1pB5qg+j8GyLIaN3nFJgmccxHasyHZZUisIhtn0HkFkSa/sP6Ya
Vv6lo0YCnj29qfqDPEs0B8KZUDc7tNN+T854aToi9MKcnq0HAB/bu4am0e4qN6+B
vsBOLOtl1XRXb00qPcrLe1lOMrhzurG3uKCfy7gxg//IOu4uDqVrrPReL9cVi6wf
ni3WytSZloV/FaOSYCEA7IWUgnC0WR5ek4QlOe1PU2Sk7taR6CTVhNs6tDbUkA85
gKGV1gwf5HU+pPpM/TM1wc4q9FiTE0Dfz3f5wPgFOZn3EB5UgFJNyVuq8GJtiMgD
cP57ylrozBN+8T8eJR71fVVp3bqG89kIrz1z4fnJliCcm6VTmM1mloHmp2tqI4Xe
R78IISB8UMRA0EjPxaAdhBYTrKiktmUGAprVoEFF2vwVdQxqkodSAzUzCcuPEjLF
vL+vgs1PDVO4QgNdjS0r4Ewf/9QmhUAHN3RInuAc1DI4VqQT9mCJ/kBndaDFcDk3
NzguOy8HyHwQ21VcaJbNYraAPZixu8wY8NsEYwd7eTO5y85u5VU44ADVdgGkmtzv
RmsfDspcP/OKzghWZ0/Z3PlSzMaT6Bc5YPElZgKYiN+9e1hmpKo8wLKudVJ2gvzL
JiaSZKe3bhUHd0Ti2uwSTKhOvd7pNYoHq+f4Hjhojt1adax09FfEIsdtLYhqWx1c
FPExhWVqWz+A42DWF8SQw3HLcp+bI4v9qO5GNROp9CYYL/QDQU1WiJf/c/PxsjiT
4T0PYlZgLHkR9GBoBLHgxAA94sMBtGiA5VoWEtZXzzU7vfcEyTl8HvUjwAYKf55i
WTZdm0fVlN/CVVWtNDoq5pno4oijAhpB9EIBOsHKJ2y4N99hRZYINRPyPQ2Em1ih
EfaXRDlpH3ZNiF/Cy/nmIKfUVhrAe5mOqKaniCV8DjnsnQZLudFDmRX5+nS3AMCq
4iErKe794RgV4oLfsdFBbsioo4Tgmv9CSscxw9173FARpf86FbvZJwubydmpOPv7
82bWwpMIPBUzxpIdtNRseuBSxePWp+eTqqoJHWwJ1XiPlNHGDdvYGjuO1i/6jHO1
4e3FfiNQ/w1es31UJlVJCRC2b5otASpUUII89QuQyDW9afv6WgzopRdcvfeHGYgE
HjTy6P2OjowVrTWIgOV8DnWUfCZE+nBOh3HpYnrqZ6Tz+s4tDFd1PeiSiN4dxANl
GRt7h8wXUa7hgh6hNzhkWpdfuBT5Npiu2cA/pIv1cHyGEhWMliqgOSJgLy6ZcmlX
AbPl1uZ1lIharqaGGl6JmekwNieBvCzm8rVAo4wWCkrAk5TdVNnMiDgrY3JgQrRw
EJkCxvTW2gby4kRCthDK6iF1UrD8Gl5dU4HQnFYtlCu29BFPWTlcpuMuRvZN74kx
SqZL7saYsLyWqJP9hoq+R9y8siqg6s5cinbOS9vWfmRogjyCDQ4oTCcSsgqc8ymo
gvfdkXttR3fuT/2TvJjH5sAQIFtHP+JmEbXjUXrPF3tneJmQ4LmuZ0NmNN1jOcnm
nr+2Nix5qslA0NBsbU9tyEeg6az9uUtInqipoCd8LYk=
`protect END_PROTECTED
