`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bwyglp+mt42w05jDYbXFC/lRT14//GfvXU+QknDnebbpXrN4EShQD0ZmszCYu9Nb
r6uCVtOgZnZdxHtnkyVvzuQSqYiixgxF8aIAjn7Zc00CUo8mNCzvrhYHk6FUtY1V
2W1erQPi+f05vSK5Hrix8dT+A2TqQeiuSQGHqBPYCo906SwZRDOcw8BBsWZFdeux
ouDCNQ49SeCwkFJCwyLOoe3m3bCtKsxt6seA7ohEqKTuBuAxO9Rk2m8xZfHwrW6A
3qYP9Tn6FyVgc9xuTcGJZzQmn+qA4in1O89wFPJH9AphQ9LXPtGMVczI7pMiQ6Q7
Qvcx10KwnBBRUNOCPmbKwAYLiIjgzr2gg2ISbxJiMqryS7Qp5xz7U679beGI1WPa
TfDvs+mN7MpaQ0lmU0/YsA==
`protect END_PROTECTED
