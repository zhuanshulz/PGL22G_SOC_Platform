`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qu7zlnVr7+TUKwfo/MxvSs8NBsPCM06CW7o4RkGeQ/ioe4SBLxRdi/PX6ouLg4qy
9pmVeRTetoaNfrz/x9ZhHys1boYUpbSWNJKIeBrU1//b/1yfJhsqijxvkn/RLbPz
V57Hb2OXhQ1VX2Oi88KmRMtzICBl/TvbVRMeY5tl9yZwtzJSdyts+ya1ntJ4renU
7K4/M/DRXsVFCWfsYb74Yx5jK/xt2h8VB9C60MK7U2TIl3Rudy89dh6gi3TQTf3n
Tht9tFzGpll7rLr3RCEg3KZ20x3tm4O8ad5MCDZVJ81jLW3vaAaP1RvbHARs4XBe
ZzzvnoCwFcqZD03WqUwBFXaXbSTo/X7AvYoTdYXjW5jZrsfU0FUAxgPwnRSEVkCh
Z+SnkfLaOM5+WYtRXg/vNwpUrH9JNTqoMiLBkunp9FrBK6O7SMwXkRFt4BZMCd5a
tWvwYjco/wgauSkIg7FHXoaxklJ4n3l8NhAKd6do6rWRYm4D7LVq5XTNJlgK8i9h
cV2ObQ99vWy73GCRtCKLfoAupK+SsNVcSncxRwiyErxh6wRU0XnJLqeNxX8GSuFs
nfdpLKYFbfnWjaRwZXGrARPmie9/ouxh42SuhbAghtEyPp/q5unfEcRkrmww5EFn
XMbrWmtwwEIVG93tx2jZXRDdwp8q6RpyNZvCAds74AEdPBJZjL5oZt+fb31roG3E
Cusj+pZp1u0F7yx31AeKHeT8DfQ3WQPLDUfLJKyRvgSJMrtD6rcxdQbezy0zE1rd
8cXKaQI+ABvY3UFDZYM0QHjefcNGwwrAqLT7XEeFdtmNDyxFf0X6cu/SbTQYOd+4
Vta1xXBceqYPvopDfaXwyQm46J70ogMufBMhj5Jld/9TliXZ4dPHMnbpyh0cATrI
q0WSDCAMwuzg/t8In5m81oO3MPBz0Y4sVxSluRmYGl2QXOOzMGOQeFpll2lFJvbC
VahMv8Uhk84uiKkhVIFHN0lI3ZXXV03sDaY+N8UCu015/3UxCjcfQBDpFC0B6xx5
VXxmO77kb2dqyHccBmq4QjS0BIf9960HpqfKJi/ij9jUEyZsFahmCcE+2djvckZ/
wQh0C02ZYjY6Jk/4CIwVzhRi1npABPODAfqYup4J0++ViHJd+JW/bbxpnQIt5sUM
8sDS+UN5J6HImItA0/7VQW2qMU6qBm/bROZLUMAjSpi/RUUsnNu+wEAZTmKMLF8U
iUf4EEbv1FqWkoV6P7bQRmr7B1qoSUWB2a91rSpGskmaHybsI/iIvs08EHRFzyTY
WFUPjPomtalrVcc2gu390EEhg0QVxQDfH0GTx5GDRaAFR1XWqSOQBkbyxvAviNOv
2w9qnOhuZwYjtmgCERpgoCqRMk2ChGHnjuXtsfrAiZljn5qvF2vOfhGWgE8sGF0z
vUkH9XEXassC0WX0nd6TG7LJwIFSzys9B5Og67lvxeA6OKuDbCigF1A3OXQSjM5a
001/xmjK4kE7/LOiokUvit2ruYz9zp7JXJdwnSviYZMxgi5Fluewq40g/ffhc5A7
LhLtLBDwEr+efFZrLd+QPw33ErRFqRwRlgkk8z4TCrojvQ33vkrAo0aUQj0Ud4nM
3l8udHgiGr3Hf2fl2k1S8nQa1GAKxBCq3M4tdbTnm5f77Hm1md86cD4VtKzW4CnL
aeTGIZEi72BZOU4ESU301RA8swLTp9R1tkwaZgyf2TYaQi4bBbbm5DibMSCh3K+Y
0Ks317KR3tKutkzZHDzmR7R34t64/2f4mGxLJYJZ1QvPKZp1nv9bHWlZqL1ecaw0
TZ/q3HM96wpvA1viQfQA5eRqF2hr8s5/zzb1l6BQxdEciD/35VRaj4duGjGqC9CR
kn5s0E8/rq4D5vjbWwQlNpPS2DWOZbZkZpXfaFtFqpygibGzJx7dAkluZNuilJVy
KfS8U+vRHY7EDX2CYQDLe6k1uz0fbNn1WRoiPqcUv7uLZrJERgq7hLKcWrMGUm8/
604R3lGfgEEmocyAaf6Vg5pOSCEzcL+5EWk8c4OmQLucgUpwJx5qqW51rjMjXEJ+
m178lLB0J1uzl2vz4LTFbYgifGq7K+UAIFLktUYCTHCodK3qIw7H3OkSIv6x8jHJ
SsOygCgObkSfDReQniLvnp4/UN1i2eMFyzWqpPnMPJlfcQjRPYGXNWE3IarCDOnh
a4RD45qKpLbdek0J8QogyfVi46Q8tgNUuXYyzGrh25XQkPVBspSM7jAe8n8QbEN5
A4fxZrM1H0/IE6o+STIFyA==
`protect END_PROTECTED
