`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mVe8XjJEr22yKoTrwGvjRqYo4PvfO/PKWPGiLEWXQZh8TIX+EC6acpmu8U4304+o
KVLYnIts7UtJq9Vcj/As6xryMigTUgvUJJAz0CkbEceLQOjU+6ReMxlWtwD+RdDU
d2PDQcZL2Jen0kNUP5Dp/jmvi7AkbrYbc0AqDFpKLCFncNTI412AnoHkb/2+D8A7
N1qfRwC2eHUO8YqNUOzRuFg9FD7Y6eEV46OZdjzVt7uWlL6K2Z3rFJFv/pSOinqg
8pKsqBrH3teUhmLJPdjkL7/sg2gyvWSSWKcJtRd6f2oonVJBHvKRVXou6qV9Qj9p
uDlxN4XaGTeoSdSJIp4V0JqLTRJ01m9W1pwR689YHSGf55DZVqlLyMWCIbt8tIPq
2BLVYt86U0Nr6XADGYljjG/sQwrRvOteS3NMikTGyVSyA4KqZHEsX6LDFRTofFoQ
LXYvidVChaBba09mFcixcewNxBD7phZ9VwCCbkOsjcq2G4jaKj3tO89QHohG/OVV
ref4CgHzPJAutQBH1IxZ1j88n78gzmf5ck0tQD2AeRxYBam698JrRwFp5LMpL6VA
mq8sNvaJlYJ5HhgflXBP8RYejL3P3rzIyiBqWvaZWZ/syK9eufYmXQH8r0i2In59
thAvzTN56Zas3bQhKvLbSx7zPSgj/UOJ36jrfc1St9sJmNdurIwXSoak6ye8lS+q
BCYpQBC402bWtuvrXtq3veDU4hEG4jtoghHlR6+4X8eXKmTDAPicKQ4NaPtRZBaA
zOoRkMBkD8KkpRWzjbJyLFJFMDd9QfTqBwwzNcpcQEoUvn75PubIBKz/0k8JVoSS
acZIPjArTiuKeepTzmhYSTLwRxO50SJ37ZCogQcojZrFAxvNoy2cV1Ks1YQQyFQs
Xl6oSeivxoSB9guzsXA8GzEOnx7I2pgQ85Np7+R2TwbDxjsAjB3Iln9tg1Wg1gdN
Mu2BXWc4r3Dci63ttQ0Ad2v+reILi048nUWLZg/b2iSlV2dukcZu5mKbKpmLP0Km
9SFw/hmlm6bHS4IR1DXrGg11VMDDjL9MZDYWUu0AwE8OLmZsKTvuTakNrslknBrh
FYz41y6WfpbUl5lARyJibTVuA1DgedzhP7gqQDDslce7FSgnOcfrNJF5k8ZJLu0m
1nFBRUdsUBeyhNo/PaU+3L7qmL846a7c+k3cQbSaEMs2ncXipJZnXJTfPl6BI8ON
gt4NfaljzadkPewANnn8ig==
`protect END_PROTECTED
