`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
39GkoF7/4eb8OJXHZxvrcU6x5JKQQbOpwgN4p0/zkpWwtzAEg0d+78VO5M8SvMjr
lrmQDsV63e1cMI65eIX5PKELIx4OaWH8GvjoTqfJeBYs/ztDQTSXr5hWDU528PjB
HNcJqs2pX4ec1BMq7n/cWHUiecVFRxlL97WRYFAnRtrefhPwyTT/5gCeoshMxr4j
wtlnNcJ21rQoeJgCSgn4F45dqu9jzrc1Ec53p8A7XGUvcIiGGoB17AQXUQGNJuSY
2jiUl2NaAGeOCQsG7fBAmgbuCpgT33xcvUPP0pGdvPteIJUURdIuhDgsenVNW3iV
etNLMa7lpygQMliUIK3ePlgDgC1VvTi4RS/klu7QKllCb9cSs+wXZg2havtq3UH/
a/ltj4sj9aqFHnMQtzc0CxAei1Wgq7A6llisWuOEFz+weFabjGLuLfYg1zeN4By6
b0GHIPP8nklhQUmEFF5Zv86iporpAc2l12J5gbFHN3HPm3EbzU+1jXR/tuyWDk1o
reud4Lhc/XS+Gyzmx/hcgSFYV/uiHPqMfoZKsKPVW6+cYI3VhWVfZ2PVra6ld0GS
/zFIGJjlwGMUq/WSj0vVb6SD4MAQ++aVRP+lm9eqa9c=
`protect END_PROTECTED
