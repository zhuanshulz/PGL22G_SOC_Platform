`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vvfw8rG0uv3y3WbOfeVOPaBHiCE4nUVWcC+j0Ol/pxxD8YyjYzTE3N8snrBF6pOU
P6POcFJoJsskJd+8YuTPnu09XHAKCDRI/2Wjs4X8MMZrFgtVjk824LXlM4VbK1K3
LMZpU6/Kbyg3KLBf1nAJJCNaYD+gQZOhS4dPfWzXmvbtXTDuavt+4GbrCiYJ4cLG
KnHn8+x9AQGJB6HBqV2ywHtYCzRsIQDFnpOqbnEndcekLTV6fr7UxrmewpM9ctR9
QFvw+eSQEzM4G2JIQkQ1QazE9GOL6gfR4Bkn9rVL4z2+Vpb3+ryd/bVPL+CEBR8s
Obxk4nVvVRjuJqBR31jfCztseUETFReEnqTsLVq6P/yGq1bLqsE3l2iCc5nkUUY6
qcfUG8cWRcjk6XtauvglQXgmcCAY3KGiHY+v2nLCyJ/ILmToXFC9USCsPDjyyf7k
QvlDiBEO59aLgq1O9eNUDUhd5awB/FtZAGOw/4fBr7Xv2jZXFCVI9xzYyDl8gCBk
yzMdlaNksmEvHuimAVUbXljnRw8jdS5kcjMYQLyCxRiNw/1r7mdhNK98vyAQZR1K
WntzBjrmomCcDcz4LqpdrdERaoBlmBeB/eadccCVfDS0sWNIOEEJRLE8rnNYSovz
tuqhYgVcRxClYcFjZag/+Syk2pZn3l+iVXLS9J33O6ciNibB3NlVrDJZYw2HCTsT
LP3ekmeBAo22oJSo5/wFY0Z1ng43REL87ZQZkiM+HAZ85BccuZE/oAnV2lNhImIf
Gs58Pi72H+rKr8C03/cXJH1K0ZsDXfvZi2GjxATBBgYHrwM+TtvwG1v4M7MoxWnx
rGmO7/S+R837/VlE6qjpJRORtUbdi3Zsj6SWjoEyT5sUB9NaK8h673ES4KXqGtf4
iDcW2RtyWHauebxH8O4M3qWHn7vq05QeZbrkz2H/BUQ5GMWXeX6FDE8x1IH1FTnB
/9/XFP0NPYFuVJJEzNKeKDyy8qt5heIl/IcG0wCuqArSpbCe5PbaW0zir8Epj9b9
waTjoxQhsdqB0zqUnCMfuv7nJC9/F+pVpSAx65pR9ALC153OmKS2fsm8Z5XtIvZJ
nKWOBJaa8wRbVuI+cBlj1ErFpWWndTBs3EbT0ORAexV4PSc4llTRFIUNwHrwALMZ
0AOe4pcnxXYmsTOIz9j4UIlMFRxGEQz2LRlGcqcFaJ1RNwSRYRxU9ax8ri4ZW/x8
qgl7pkIvq/QNB6uKFS7LwzCTXw6Z/jP9+QWjRfcNE4E=
`protect END_PROTECTED
