`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MHqwGu/vQySoyJ0Xqh69Gd/rhlW9ZT3ixAWcsafYV4cMTKyjzrxA8Sto1pxN5+N5
XTLJfKY0Ahtt4XfeL5T6pXzW3f05pYenaRRcTGmZ7NJoNK71fx5U4qFsHNWSJEz/
xp5zRrPe1EwfITYdn9gXsvAA+eMqKu5vbD1sv6HYAYqAA1PhKFzbzZ6nEVwVdUsb
HUNuShnB5f/YaER0UxbBc01sEZks0IBYPisOEqBYcyXfGF8qIuM4nySHyRiZr1W+
mMlPsBF+HjnZWRVZ+DcOGS9zVFZAQOOekUCj+pcy5Tz9lXGBFJM7aqZK69d7OLYK
qz5+W9J8pg9qVYSPBmhMbDg/5+6zKQLdK0DnNLPwgXJZioz/FfOE9OICSaYdPI+C
prfe93cAcuCtpO3m1LOm8qieXnZCQFhTSSkM2Awf4uVFFpHPdn8DDIh4oiEHeeq6
kBdS3GNfWOyyEaAk7TL09GU3II25qMr9bc++f0hDlDTlNAOj7c/yg/ZLayhTS5oi
iwDDGZ0JFtFtfq0jXUZdrOIE0s7Kl/2NO5cN3Xq8bMkrdA7fUbrOBLNJhV/2h1+K
HPs0xpWLxujsEny1dGLqaSsbE5kov6+sMG8on3Vx4PlXVbnlIYdh4oWLw5nN/yBL
mWFyjA1JiT1r5Ji6nHSPj4vEQYB62MyLKN3//CFcIMcxE2K7v6cRhuLqY/O7Bzdy
2XzxcGXuI6ZaAPxaVBrHftFnPkF4Y9jZdxRqqrX5Bgs1lOigxcfAWrzAgulJiPO8
v85FKRMtBvcTqAmYi4o1DgXNxH0ozmbs7JJM6uYdf5AX/GZi8aZFfBAoeVa56BlD
UuQmHhFUiiIt5aHDJRvVEOEZR4mwXLD9VI6hzszD32yjFiw/y4essVdPneo5W1tG
6pXLN/b2soRlehdgWolxacvzSkmcgaGisHS0oeHhyUUpseJABRlVP9MH4ul3jlu7
x9kyo7kMH5FRBo9rlzvzDzfMNj15ORu8nBWZ2Ykxs8mg/3dmyJlfOlVAGe6Qpzme
tLcLs/oNLNguguSpQCKT3keed2fMb7q0rMsDSWTILkltQh79yrjZKWuzOULxahZT
rELYW8JQ3X21zQs1KxGsbg+kaUn16PbABm9cnmrohmx+ypsVlxa1sxo3jEqCsLXH
/zqPz6xmYlYMNIbkARgXlSUiKEOlQMID63HvBiyGKZEBD7R6ZfWlhwV97MxtB8bi
pGVNXWU5lS4DqKVn+rmNkj78NhrACiPGdnK0RJIq91ox9EEGEAqO7YtI/9yPrGAG
ZCbdC/vQB6qhfeacDDJ/kUaZ+D+Un2N/MX8S7dazFvEyhB5EesRDUrY9GKvi7T7R
BClFjCfcYC+QeyCaUuIMtDatqEqR5KCtmCHd/jUrdvfdwCifiX+h7hagriLlXcqn
UKGUMquQIz0qDO+iiVgMDJ7ucquZVa5B7EmmHLuWqDflMjjpzGBNYWoKY12Utgjt
pDTWuWn78csNs2c7TaiCkm9VEQ+t18RuYtHMoo6EtY0j5zqecDrdeq0K1BDzhRmX
Z9Xks0j662MWU9/ItdrRkEVoSI+OlfAERpKeQxY5JWz3s65TNnUhT1cZzeaNfUXF
ezyEsisse+nKH35MjcGgvcHgO2nEV+2WIJxxsb2MHRuWyjRU06LcFiF7zYSedzD/
+Z3V2LjuFYbj8Gvqm754NMmWdQCaPlcUbjKTGCkPg8ENYZWx3+Aevt1BarZYzlFe
kzlre1igRPA+HIDf/x0cOk/iXmpEmD//CSIYiLh6prNV6WRwJbyIcqc5nmrP2PW2
uDXUmXxjLpfVzaaetcF93Z1T2rOmS078wOeDRzmLr1gbUo4FDy4k8k6mAssAMWdK
OBRIoiu9nzSNCLdnjUP57Cx5fUnv52YZBFQ58HzaerEe0O6W9zDxxAmi0JZBtvoH
yvC0CNxgdZ1KLJDlahKdeC+kSOjzK1GuEHFNqEampIP0/nAxf/zqp1/mjOlf8qrM
vqLQzOFSuyvvhUOFx7189zr5aU78x8v333SYmOiV3TCJeFBCiJP5uaIYauxoyE8N
omIzE09jnQKxyUeUpNDuEHixjvERBioN4vj0U1Gh4bJoOpiJm+xbe0+Ze/5psYYi
ixcZcEF1OFgU1fZik0mLU2XowW0RGHH3zlrzKi/27CDvJoF1aJT3Pte3v68MXAOD
Zu9/mi7mRpsYDzW6uY/MT2t28ybcZNngGGas5s9acE2F0Jb5WEmL9lsZuPhKwPEm
edhzB06TK/louiThjRKUdDRAyVQ2Lvc4eQl+Vev04Gc1XDYmtSl6dJN+hGhbK7sD
Be3yoczpfb0f7FAa2tmliY9ltmLccNziLY+LbSWYDp5yBrYm5s34ZBaFYZsXfyFu
38VU5FPaDhdAL75X3ZrJ9B42NW/8eAG/QEzQ0iLinsUt4Y70KTyjik28SfHNuhj6
zr4WsUm/TSQKzSkBDWW66Qnvd8qUnTQh3OgsstWy1hlRAuZbRg5plwhQe1ofSTUO
KXnUd44UqukoS0tvbCinTlZoBq09lh9w4hu07pcmyvmIVFDQgsmT4mgFQWpAtEW0
1Gn7o6IV59vph385zbYO1bzisi8ADP+3Iz5ar/aPzuBP3VV9XPmN/1YMvnwO/xPI
PuSh+WRrmcoKaJjaCMHfsZNIAArDntj290axP0Sav+OQ5qggPy2WJS66lmBaOQyI
/2DjEDR5xmLdPPmhliHOq9LEhAgJc5URCyTO6jLLVSVB6MY/xix/I2vPL7a8TlkH
56gsf6PGJ2XwZuqnIPX/DRoqz5mwdh36z21ysW3C9Q0PJML2Gd7lIP1ALE3ToWgK
eoQS63BKWl1esuH1Ju9Pf/SL08ETMtWRajfZK+gbD7qY6mHDcW8Vg9eAF/6mPQ4n
dhxwPfyOkLK2o5q/Iwk7W6vJ9xoXUbqG9fZi35i75OvaZI0jdDVEJPPs7s10nRfo
OTzPEs3UijbUcAPfLfqadNA8ZWrq0ZcMK1p0WAlKWgjSAYParPtQZVQ7hDPOoRY0
ba1tnP2zJ2QID/DBt7X/8ZWYmfR7uQ7SqmGuKk7vYgRZMtG72LSVa5KpK1p5aCuZ
c87nvRsBE4MmkmM/mODCB35pU7Uei5fMfgM7bn3DNPvBVGDbQN9UXIjvqtuD+Ek/
DxE+JxLLkm+0bZP2MVb+Asig+zZewUwfY19T/F14IfwIHwBiuKtHjK9D/a8iItiI
Yk8+dt2qOKtsbq5p7TlWE6t5TG6Lt5EvxTSfQ2UgqrG2VTWfFL4aHXyXtnA2ThXv
SbJbBoQRGKrhdf6JKxgM6gpTtN8tnpM60l6JnNp2vyz7CZPdpHhGuVkL+nXMp7Lc
V2MXgxmpk5gxm9ZIGKQ3R5ywyqI3uAxMINP+1rLLziQQvfVVKpZizgmjapFNtvdK
i5UweNfD0NCWc8TSbK0n5F4cdO6Q0x0dOjKFyJRQUYh9rtsNQT1dIH6Ax00pyh6B
X6f2y+b2lMewd6qNfJ8vik2Qs+UxvC5GUgEBtITZ8iTKfsOkZ0MAl4mmua0CPJr6
TLsh6KyKyIM8nYBpMAI0mT7mS639Cxj6xViS6rV37a9L4MGIRoeT8piKS7ERC3TY
hZ/fH/jaaug1objwqtw0uGj28Gh8XUvyl+RF73vANUQdaL8ISQUM0ZoewmzlVX/b
BE10oOhp5/Gd/e+/vbIZNF0bqYrQHWLUZAx8RUE/QrwpAxzl93/Krd4U1EJHGRAo
nsyqh6PbXxUokD0NpoDngWxBLwEHUhwaEHI3jBtwFF9wKGhzZRqH3hc57WG7XH+m
4dfP3/T8NGzOltcDappTFUm/97pus9EQwGTBioLJv8vYXwr1ZU7ZxvMPZwMJLp5z
nHlI8phmWflBNm/7yYY8xZ36PoHS+SVcelD7XOytX7BYXPJA92ovb9DhLBLkk0du
j0Bg7xCenI83Cbb68C/bhDMcJxgLX60USz6nmZPycd2jBze6XWW3fVp9AC5BP92i
cpgo7udoeoV9PFy+/L+MygSgOb/qXYWWHDicBNSJljPCR/mKA/mfRhva2gWZre2s
mL7uVfsDoNoqN41dVpp9WVLpwrVd9deN8JDSNmXvL6gcDkJp6WnfQuO+S6GGXW7l
j4KhSgyLdssWqNpn9HxZEpJCEj2kL+k+LuRVUdLsO6Pxalmtr5IzB4GeO59+YAg9
U1ZmoRyODl3UfBqKXVBL4iL3k7uccroNpIteR9+9Vs3iO6Cs9k41mlTefktz/vLO
BzOlOb9R3J6HnBKyrmtAvdVpkYY1cEiS6lyT5phL+/0CZH8cU7h0cxJ9O4WPSLTc
/3yf2r6DpziUuPQ0UdJ6wXDKrcdB8aSBAl3RXTMfQkIK0Ul6xmD72zRF7RVpD6VY
3IMAdxlNhJe5fo5VmmhMifgN+lrKc0WQ5URgYiLCh44zvdd1qQvYOjsth8U4FSHB
mGf9G4aVYZsFIATxhOksthPUdgHTdE8qmWYXAuNA8QefO1ZNkCS+jkIVyTcAOTQS
Jpm3b7P2eI1Xg4dPmrhc9O0nTltGJcDmXHbwTxvvf5dmY20vC6qeVjE+5w/OnTSr
y2fZVDc2A6LHdUcZjz9m0oA5XOXdaKRXUmCYBRtBNAKBKMFCeSDmsYrJ9aLfJ+Rt
p8ovRtde47BJHc/PKXkWNwN3t2R5QDc6QVCQoZieB66hv4bPAx1RKj0oUYu3qtPJ
Rr7L3mHu7L6+avqXADQ5yJkcvx+jZRvW0w6AnwdK0lmbLYBJ3OV2xzQVfmd/tw/H
wSr5XcqutZpQraZwnL6X4a5Nh1PFLe3Pfs5pd1M8z6DK5nZP25uE5J6m4h9IWAdX
00mHrkBlSD7S1bJ7bxGAuGUgxGY0RH692IcLY1J1ASPk1G3/ovk6wBTliG5styrc
0YP9sDiFnBy1t63QYYT//0wQgIHYlfHDtb/A5wm+JRMXTc2H0Diep9Q0howKXDkQ
NX5xgY7oywCKoksKtJySmxh9cZROOT/Ukw4Py1MO7w3kbHAy1oa5ZTeC8KpL/S7k
GebuzkFLqS+CbNrC1mSDoWgJ7gzCIPMqZbBl2O+1T3pEd7XV3utjBoWL+oIKUKuy
GzjZGazdYAONHXAGw7Fdix3swmuln9REB1CutuInYgIqcn10W3HFTyNuYHK5xXKI
0wNI3G5+wIReSHajfmBSxkSVlTX1eLfZFLtp6aFoNZmme7kNultcIzQeMDMgr+eZ
LXg0JkvdUeuqfNZnnWc3+GN+foDLxERab4dV9RhxGBLGZpsCvAGNVJAxZIhVB5ba
2It95jh7nMNJhoUewiyTWxCct6U8/BaGJ6dQ/vyt8Ibtn4qUWeZRwFGgTZKvJB3h
8P7GAduP/CPJUwQsdjr+x+1YJQ+P8CrcQ/gEP/Bpumw=
`protect END_PROTECTED
