`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Pt+7K6ytW+ZmqfACA0c+TR/vD201ceE3QZia2+WfySDJRYHF6BSpgZrfVfBxK9Og
eQ5GJ+JeXEFh1hS81KCmYHPakEJJmwGCCp1ZcAUPgFZcRxbGs3qLknxy6nHpM8Wx
Tjn4lDl5qYXuvKF9QrTQFvzBPAskLTh7l0cE7CG3951ePZGWhP3jnIVGKAAR++bh
75QlTWgnSVOMkrAGcoOy+088UlfsTVaOx3NrWNPWiAtdjAwGIvCcsGbSol2P0ZW0
M1JNxA1zFF+molw8k8M3x5kOYNQOk+fJHYRTVVH8XyXnyZX1x9a2uib+JjQj0h5o
6RGa7eLXMP5H8LcfX4kd21o8UwMoz6nHimwiSZEGNYDxz35S10YwTV2gutHL3P5m
6VbyOqchDl2kFJAJUlHOfQLaCkJzsg1x3gYm/wbRV8z3KTEGTKBqkcyDBGEkgHcQ
Cr0NFLGGg9w5QEUq0xRDh0Q1aHVRohEJ0xx7sTw4NmHMlOdXynE1EtDh4V+VuqYv
RY6l2XpxeQu5INDvHDUz+Zam9TsPxGWEwYkou7Qb32sMa8oSUWv5YQoge+tefr0E
1Nrj3LU3QTH0i+mX3HVLnIbBTI8ZxmbxCSWhLUZKLUxTAKUNJlI2MLvWbQrPGJ+n
Phn/6pHYb1tK4aPExp6rxXnPbCcXgfcPss0OesGX1xWsV8TM2Vm5M8Ki9igYo/yL
SmBO+iAj/7/GjNn5/Il0iJBGlg8C6hcRSqJ0m/XOSch4jjrgpvDOVy9E7mJiOcnr
qpuOjKNOhBIFzr0uC2/9Bft8A/06yEbLqU/d+M3ntCJhaBuhSBdUJgAVorvSxDhn
WZYzok+Ujq9RUMvF5bImZcgUJf9qlZBgBklIYivwPcZ0Cn888JObtJpVD6joOZuN
`protect END_PROTECTED
