`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rqck/A8Fx84NghiEywuLMg3vC2vBzT1p5gk5kGheKncEPONNsED3xkMl+eBjcxKD
dNVPIES5O699z73g2m+L1Hk2mbKB5RJE2ajqihVRmCOfpwggKQCq9itvOg9vtB4K
gAOGeD+X0DxjN+IKlqhtw7ZYfsNfz5mqqZt/V1DecfEWQGtC36RcowoMR84i0I2J
5aOvxgflTCnA3fIXazdrDEb8rjm8GqLukaDRACMLlT1FAlrNoPcThkWtPkddrbqt
egQ1qoNg4npimsaF54ei4Ya3Wk7JusecqUFnd68X/kh7uKDKinbEVUxd/dFHm4ec
NjS1ovB42ThQirNGAogZd0DyPB6ULKXxRFG+/iPzhsIo8gylhENUy7aig9jGrrBm
wW+EKpF9ZJ5bAtuYAI6SYzpVW9ailZBh9NaXpya8P+645kNiGZvhdHmT7BNLS8jA
v60dxKa0cz8twhHKviVD652UAtFYCyQewo+KnKN76t8WW7XnpH0wRLa/N/8tJI5a
oKkSNyYVxtRRbE+wSg4fXfY+6/AKE+iuOXg+CSGTrXGjinYBpVrHQcBLKWfNCPMM
fNb9Sczu1ykUSjNDEDN/AA==
`protect END_PROTECTED
