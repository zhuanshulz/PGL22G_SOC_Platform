`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oeyx51OTPpRWHP9AZ/oTH65bIOPD7K+vDBkCaQxMvBQPUKOQHxXMp8nLmYoGto1j
hgzANhdmXY2wkdGdESkuxjQTn3bo810RZeAzZdA7zgHV0YY2sa7gN1SW6bXOG/xc
Rn8jXqXvHtePN/nN4rBulRzPw+IjX2XVeKbORfUG29wHD0Ofs9u7XsAqMIGgpcgt
8StlMzlo0jFS99CqBiyQMzqRR3JfgaCUG696DtEGKjiNgOIZyGWrXLlod9gEqng3
jRBbg/liiGjzgs3DVkhMBwtokzSgr4TDJVlxkpiKUi7Oi8qkszZSNFj+2zVktJ+I
eG7E86VKMinqL0E4ha4MZDmm5Ju/uyMfAnQkBnQWeDnaR4vUTFZiX2d1kMa18Rg5
nAeiM61oDPGqJKvdce7uQTNgLoYNfCncN13MD6PeCmPrTQwNdQW1wBX+mdUrXp0X
aifXnFMWkUCRF58d7VskiI8u2qxs3H30J+gLtJOjIGg4tQpHnGfKC7bS9ZadcxsW
hPBlrGIZPTRzjw0hFppKU6NNMpBuYGEKc3qvusl5UVFogIn/fJbWkr4O5Rw/Qwlx
9eg90n9GzHDZYsVzwXNtWWcLQiTFESHSvrvbCqLfWJqzZYJsU4Pqd/K9mJ8CTP6F
O2pg+cwVB84cyo2yaBuLpUxwNH1qPeop2ugq9lcWzYXfKCaGKrT/GTy0Hd3OWCuY
QmjRIiktjTygsxHNWOqopsrte6zn9Dzz2n9RwnGDRiRvCvnGzEK6aNrPu4PajUVS
diXuDv4IW11uw6//PdSP40tjqZ8KXQEODBxOtabKLpRiT1WGhi+CgpJ/vxIz6fPQ
/9H0apB39m4sHE4R87AWgOOsrh3Kh7+yIoyKpvSZmGeuu/wP526W3BBwh7VqSRM7
BEOUUAkPjiURBlT3KGZH3mthUgVkgZKTJpZBBiQ3PDYaehasgXm4W/yHuaAc/Bwh
Zk11vROzOJjgyACvTf8Kv0MPmZ7W49v+8ezbjtkY/epFAp3ZPpUqK+6AxzLUgH++
CycQjinm5z+9YgBMJIGumjYIdVtt6mT9Lzlp+Ekeu6RS6H+0DSPaLjxloqMl8g1o
G1sV8u0yyowtiMXbN2C7PAElI+4kqzh2zugYrxlA46qDFOswGKFAXgLGB5pS7iar
bhJxvCN7hdLwbl1YYOl/qwAQx4fVOC5j6t4MkrAfVpZ205tasm4SNRi+S9gnAfHK
bJ/J2IHCKmCxadAqO1UMzPftjOLkGeov4X2aK06dCPU9ICAofj3k1wj0XE3liYPN
FJhFPyxix6ki79VGpBQ6PPAe4V3zCJGvz7dd2uGFmn0jSfH5h7jPMjDJdTJSYQND
Mv3+/ovdmgNFqGni+95UTovWpYpIek/oxavdVhTpN9xwmuwNrm8SEIDOrzSKIy1o
o45vat9cmW7OLrvfjfG9N/v8xGTLuSsV07lAqxihMD1fJjZhC7ij5W+Dao0fMMQB
`protect END_PROTECTED
