`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gA3jV6LLTIzfFMNYQRVofrYtp36IvVufycVw4L+ZFv9Dg1NfWiQXqtgwxbBIZNx2
bcbsvhX+0E0jhBun31FGUuuoIYnCqEshBTZQJLnyUI1jGF+NZ7v3Xf+J34j84XIr
dhVCFOFl8xFUpmYVt+r00/kKp39ySfW/8v2NYKhV1Ol7Qs5BQjM0sRFZcO2XYaWl
1muXMtKET2ld8Tyat9m7SwuQJZwrmvZz1eE4pwZrqQluHiUOqSv9Aj8+9TctlcQ2
kBYbcsbZ7q0vehwYJ1kvPn7mpOtAFf1kywUySu8pY3nNnqojmKwPue0gfqxrym08
98ENl96jjUOa43Ntj8Lvto1setvteqNzFmmLVSpHpOPwbAxy8Vn0pc1ZfbVx1JMO
UWUQ0uwWquMYuvFFVXmEgAZ4fBLoEKS/KCuf6L3TJOLZsOQaj1GryWJbzcuMfZf1
Oh2f1EDDrTZoNS0qAY7gelMjDaVzmtZlzei6m54ms56D2ucNZeLQIrOnz+5cVkCS
YfBvNznAlpsgyJlEP0lXxFF/t0+oIIeB7MxGWL+bcWPMXTUOOFVhwaRJaeZ9hVsh
JdZoIbv6Y6TNQnRE91yRDgHR68Ain2mSHXAiCyluRL2zgFQwEr1lFBd10xn8Y6eF
m4pVAzF0WR0Os3DdcNf76U18t10WsNpmbaqf8ULTyMdFYNZcUHdOyh9tXmULfrDK
+OI9dachltlUAZO7dR6AJz/qsxibQSbkvxEH/bz6KgMvbzKa5g9WtQhjSphWHbgV
hmzDiSU2F6R4qhhZVtbCjdgqqUXg8KFNRva7a0Z+5rlhtEHtwxX1K86QGvmNvSJl
8k+upIlLPCXi90+UdfCGVSW5ICTgN3IK4EDJwMzybFnd6pmYHuoJ2wQk5JG/9Czn
wbq58A+ev+4vd+wxq6CbnWehxD6mPbyCrWW2TjVGeQw3IkQIsDVeEEZLwqTRcvHX
znJFajFw+GAhdq7WMstt8B8enAnTSBeUeSIBPE6KfLhIiUmIlubhLD8c3cxTCuyI
tXxw0sTap05XB7i7/apLyuDq1zGEq1bk2IUNKPOu5yIoaXJNp3bIqry4mEUeYD6f
7Q9tll8pJ7wef3VnwMg6qY7/EZN8udsIwJ1KTHHPB6BldLnl8gSETZyuhI407zYX
8PfkbSlkwTiU+vuazbwOnMGRy51TTy3FYRiuSgae7ItZ+BbnuiE1qHGAs29k7Vp1
`protect END_PROTECTED
