`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6TNcZZDYla7faJZyw3a7QRTvgNJZsPWg56IHSHyGnKYloWYy72eIHS1F/YTSsJn/
Wz7vI1TWUEdDHOtSMG3ZtvRVGrEBYXcWun+Yrjt7y7mJl4glTbnoZhfcDXm+Nt0W
6vUCrvVCQK0hbndpQ71TLJjLBR3hyZC3zawDn545SNx3QELhH4ZpS0lAnbfvG0e4
CL8mclEsvqkgLeFJ2tCZtba14h7mCPEfvqaRxMPBL02NQ58qlJheII70oiXUIN+S
8oZR3j78B6N+qON/4MuUY073sebN+0vum1BvzHQPg+X1VGVFnRk39pyjA6kTWzjN
i1TVdLnJIPbKs1IYdO7w/ru+oYw1SGtZa81Xo5ZKG2ymu41cJxilNH0gV8GyXe17
5j9nZkd+Vm/JZOUOW1+3NAVVEEt7E5HwxkMPqXEMol0=
`protect END_PROTECTED
