`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8KTsuUMMKDPFpjHsAgs8WqP8rWUjNc7eKlw6s4iyezw5+dglWCXZQ/z3EVdsfbUd
jlC4uNxo1WDcIYgfoIVTudq+a3KDjeRzvAIE7hzDgerIkJiao1ucEWtropJKoiBL
HKjpzZZlwW9sPJu+zcHFYsZLwXLYBhEC1L/AZUqPr9cZqLOl39q3cbnXacOEfgWa
koRd2mlRny1V13f64+Sqy31Cmp11RlX8oO7Mk9spVhcBg1kcXXPBCXmSqeVI0DtX
8GouF7/vQeOTIqeucE5oWEMtaUhR8/cj6DIKblaLhZIfpkSf0SkUaAGcKeBLJ2r+
ZWJaI2Z22RwGMJ1+CNqQq12tuZTT4A2MF4eI2ex98JHMhEp2X2zQuI6+XvQcY7kV
NEKn8hj/lCd8P15NffJ+71Vbfx/Jaz+GyGyENJEUYc/rZbzu34B9c5N5B+oQmoT9
G6l53VuD6xsXV1WdqZYtBBFNi9Z1JW1Tz4yKAlhV48ItYqlogP/yo9kXQHewefn7
4abDVTbhL65GFgXv/NFH2RBSFbAMAbVLiHJCmc2gH8s=
`protect END_PROTECTED
