`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9Sv2EUuOsn8p1z0rQRk9E2GlRCPlVe97cwlbpfKrBJ/hoU5TpP8lnUe94EEFOmX8
VYijhwtgA7y26VN0SBUrqnjX2MFeVNNGoqyr3o2DBqzPN1kwIwRHsWlgzgXK0Q5C
2+VZ1oykYCGmVvjItrQiA/m0tqC4hP19UeblTtRAj8LlNahTtDDm5xlpDp/ER8gc
Ln6HQOsHW6lwJtQJdV0XjQ3Ci65pyYTchBHqBQPTVqoEiCLk5CgAkiMMZzFFr8bH
9kMrJGDzVr56tdFtwuFnmsut4HTHfBdetv/nQ6NBQdIMatxTqBxlJb498n/becWK
eS0KIxruN7q5JJfz6rLDNGgucM/RNH3kj4sxHV7HT1ZOOyHAvusi4IoqsHv2R1mB
OFudIyA3oDz0pccsO/84b9+0ZiVCqoMviHcx6JLjo+fZO3o+mfG+pUbj7Q4EK80F
+8DPCYaynqa93KTGJv3mkvW0a51nQrj/vo3XPyHJ2eDuV48P9tX33/wAppycETzu
Dk9VdHHSk4EDskVhu8VZWmgFC4z0NfDR7Vhr1aXFv+Qc50ZQi1mqscocoutaO2Sa
IVnTLhfXwS9T6iH9DPtrlaxxUwtJLYWZKUa5rdbREpzdyQ/283SMtw64da90oZ5W
4cszdS4tZCCH8Vxn56pzfY1P+kWpTS1wli+EbYKVderZkiVmuf63DMq5c5/tpNpN
8v6sOPJzuy/VRdSj3fsE+MP8FMUeA9tngCHmR7TYGqW5WJS+ZQNahhcpnk2Yk2rD
hwX4FZH2Rvwsh3oNBUnXc+GxO8L3ANF60ewzo7o5SaYutpowzOB4+2uvGkZ3mZFd
cOIrfb5e9C4N0rA8jKmKXu+f/HouQSdP3P5dbD8jFPvmHmfmq4+sXOeYCMSm6tBV
8IPPeo72cC7y7wEfh5qEGV7khcyhrdeggLRU78zt3H53YwCBkfi8co0pH2rmJnMI
8j1oJ9wwjHQOt5Xn0J8Nvq7QPKJ3tUnv7Ax+jYNoO9lEcw5qZsPcYjeXYrDVS5+U
PLjWK4fekz0Po0Nsuo8aMvatPZVd+NnvGQESuh3FT9PUZTWg8wSZFTj38QWSNOyj
hHRe0iQpcKKx86iGV/gaxq0p4rNjDmcBJklVqTttT8ndFb2FBDqv/M4mlix+J/HC
DFAVk34yZJM/FU57NOanqztVDcf6YzVTYPmiQyHAo79Repy5EYubD7aQ3EKqplSt
yjsLkYeBisFNFQszAf6KrMkgqBe85RYPXz44XnJh0YcpoVHuOgGrtx6SWjQgY/do
RRAceNSs8MEvGkZdCSBQTOY07xc1ihIe+0wc8om1RA23HPLdZnjGo0g+AwtaUrc5
/iwC0XwNlM8Ph2FAJVP0k65i0aZwXlVURMQdA7NSgAI=
`protect END_PROTECTED
