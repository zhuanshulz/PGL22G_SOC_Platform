`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SmEs4MXS1FsOcTBYVAid/LG6Vhdh5z8iAZsRnpjrilCCuG6Nod+2G8YXytpXCxQ+
B6EHXdSC99mcW/hGdd2Z3uZGpttxHPH1PUHoqtyEUD04t3DaBZivIHNGDOCDi+K4
x/9hLv4IQGcM0fb9J6mS5C0hcSTjdJSeeHMWWyLdOIDFmcPQZGskO0JkBCmBEDiE
K3OPC7Gqw3RqbyqfeNyO6TJYDAwDJvBS+d+9SwD3tixTXsT4HWutb8AguCJ6T+xv
UnbIQ6KmSK+rFggArfeIdq8QCtJ722Dnb9a77kZgptOL0bkKrkcViYxke9KBlDAq
Kw7iZIprdQnE9SK/CjcFWfxAWmZFseA+JjrusnXJnEN5k4NEiOSv2j4eyb+H86Ss
tCMKZTW3IcRI7NUU45yAq8nZooSc7qI+VxRMeyovL2iDVvXCtrFtiT1uzrC7VvR0
3ZvdHMZyn/UX+/xTlJjMtw9YifQTB5Rsc8JPx7v9g/BUToV41WzBglJcVNaUuKXE
fbabG3/3ACDcG7+4/fRPtnTYESm6h1dTgoXiToftUBkDVRY4tF4qJ+zqFTCaTiMo
w10Ifg/ArhSCyGXtY4FCjK4BJ67E/IKN1MJjShDX06Npja8Ltkf2NeiDP4cQyv2W
1wHJ8WqLrOsDCNutRadukWQXl/isb+vglBevGXm/Sxs5/KeN6FEf0rYLQSwPGWeH
RCuuAP7zYa/KOkyH66Cm+p+2XagcLvdRmN7hOMmsrzeReMmr5dC+Lv+mScU+et15
dbYYIVmnRWkxpXH7ED2pFdhJaE/q9fZrCDi5EftpVINk7t60iOGUPYSQUb3Kalzo
/L3AYj7rEepTgR1XM6IUWv+LluUsjPUbjPed8v4qf1ROT7uqXizEhqDioVDTfwy8
RTkCZyD9fjK6pmaYWf4E67DQIGx9jtMDIssABh7AnAcYppSpsasInLkeiZEyJzxu
nb66x+oIo81v55p1E57ryTBiL5NjhtawaUesGLdmbh5LaI+P18l54Utp+GukRYmY
xFHy7I+LMpU98E+MP+UPCDrRMXXFIDoZEbiLbsoaqZhp0BxtTMlucLlEAwqF6UHk
iDKg8FbT+2RIo6PLuzeYFp9bVYPoM+3oxnN24FWwXkE=
`protect END_PROTECTED
