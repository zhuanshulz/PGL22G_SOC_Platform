`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BiQPExg6P6Q0OyN4Ta7VRGcjjjq773VaGY7/O805s2czGdnMADREpltv7hHniuoX
UPmsbszvmmYEEnC3s46wh9qqKq/C5tkSNV0RFYLdqOAoElhUhR6XU5DDdknNCKWl
B07qrhWHUN/H7d6oI0aNCuLnnqD2+hqSy8JGviRbDCjeYsMKRuNQWqFxgiWk4AwQ
rvv9RE4dYPWRjK2PIKZh/jQkyOUGfbueW+hKetXGSD1GyrpDHNuFNbHxIE8CiPdr
rfje0lWvEC6i6u3HrGv2Yfg7SeFLuyVnzM8WUvwiBPQYGBvkIvCpMVnTvNOIsSgg
tNNwVOMTIWfDDzySMFlD4Kc9VJPWHpDnVANkPhj+8bVXeYdLbQ/YVnxnFwWysTr7
62OteHfSRdOvQDMsW7kb1g==
`protect END_PROTECTED
