`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bWY70q5r7cPglw/Fh30otfSdjL15AwSHUccZtXZzhjSu4Xe0DzI0udu/ReVDNwYi
t49+n56fc9qiE6tMX/2akKFPOJ1+pTN6slfohTIFnLt6YZ4CxBoWldk+OQAFgh83
Bsl8JyC65mQabr/aJWSfrcRZRhYJ3DQ3G8l3fMB7BLUPelfqbFdNHNKjGZe3YnZ1
BNeLNIQZeKt3tKWvHikA+0UEXXSXvGCq7BzsrDWdGzxTeeQm4NCdoJlWjcAbwAeZ
MN8kChU3Vj912BDPHvYeyxo/Ps9ZTRXDHyvvrg4Hb3CscWZvw2trkpIRUpROYztJ
HJDuJlMRAH366IZpVCWY5XMPElKZ8fRa9utU/zKVyMTD/lE2pDRM3rtierLKu2/N
COkiy5K9S9y5nqnzVoWvdVAGdCrFinZj3T2abDqkJSRhdzRx6A3PAUGYTCSg/s11
XVFjKOfNw7wjfiITs5e/+IPcXD+gtYkHwDJ1jbGg3KzfcKPXn1zUjSTeJGY7wod1
Nu9zAXq3OMKmiRAfhSvdFf5W/scUZ3YwmbdDvlav39Oo0wlKrhxfxT5HVE5Sr/jb
oxje/V0FbAr4sB7T12LM6ry04KCzVKRNGU+d580cwDa7+tdm1dzFRlME0RoYUQwY
w7Ibu01pjHjec4/CmKTBJL0plc2jxaLpXa4Iyi6mpy9zMF95WnOgOUi/Lbq6P8Df
mUPiUYeSdix0ketu881nETOZ0YHtFYG3N4uumT0L5s49xjl8gvtyrWT4eLIs6bP+
GXfpMxDyk85escbgJNWLfeizTxhf+Ssk3JUn2VO89Aa2kKAk9Zw2AQegzfpdp8pw
B9yltSuSilmowgAGM9CEwdDDclXlaMUSueihHZu8sgqYs0T4iXnfcLP7gVV2qs59
nnsWs0suSptE4YkyZ+HKOSNBhn87sSInJOoGI31XmGpyrmaG6HoysAKfkjcDdM2y
ZHsKcxDbefB5Zd0omBWsyCUXbkz1onlcvC5Sr9v3kzGImILPvbcAJm9pMeWzwtwO
JvytTu+1F5xDFOXg6Ngnwc7HjoMiL0gDNIq/6xtTegH/Wyh9T/O27eWVTTAmsVld
eQlVpXvJ6GhoKEUPg6sMNmMdERBj2RRjrfOpv+H0xZ06qX/jsgTvVcka2cbq5MSD
TfY5TKPJix063/llNtlHuMhxTbEvL9aey3Q5fKlyN8rK4TzS++Qmb99+CIXBDFSP
Z/pYq94aEP049yl9v+PAMrG1dWlbzHgm1/4MfGgXFWStv1ZY0UyB7PO2UHFEvjAv
8kJpstpV1xKiW2g+lqNQYQDySfLiuKNUzpsqqvaF6dU4IxpWRRquJ29to9Kt7Cnb
gnMhbB7L3+wdKDTQZVjjx5yY7ZtKM8YzQ6juH0JGsNC2IlXH0xVxszGM8JeXTsPs
bpKBuSrXQvxlXB1Jv6tpAtxUR5XkbKCIJq0o+CQFXP7Z3qiTPIMABfLjsU6cwMGG
FieKdPXu713gt9JMS+TgOxykdlhUvrsEkRJZRz2q0oE4EFywaZAavkyMWkPF0Rac
8nnZIS5+O/wI8aNwQ+asH5V9rAJLB5d3/qXuxWoXFc0+coLPjmj28/uI56BnQxwg
G1dlmk8RaQC7Qsqfcl9BbGTJXYKsKyKiO01DWokadZ3a+oIPYQFWX6Z4kEpsOah2
Y+Z77byYpmQOIgtBlqutTk95ZLJBaD1yoCKa7Zn1F0M2X6PCg2MudgWfJM9KN3ZP
kQhCfXAEHaKEpi46yw4vnb2FXwFKgT1p36EdHP3/4uTmFTZUMvmUUJcwT37B1MiZ
NCMqYye9PsMUwgp/SGoEnNQc7yT6yLIz9ADr12vU3/AEW7M9weK+8khDibd5uIx0
OfmcCkoWYtFBKIRe+gGB2uqhFc+QP3Z9ZAZf/z9gHYBpUPJin+eil7xfxORKJYXd
A+k6bR+eL5ubH37nPqQkiIiGORz17hGLc2NnGSodnUSHD7rOEjOZ7OXI2MBKhw1V
KPEsY4YwZiZpL5ZDPwwujH/H/dLdKg0bgwnpEpnjTacWHP5fzMRh1jzHEnzevh90
bghmxopRpBohgRKeuV4+nJAxQxPad8g3gXtuVr+oQ0xIO/+Gt1ASXdJs99KcMGsb
l4TegGRiRJB3Ajm/AkiThF+oshWFFgAYs2B14uIm2AUkmr+omTF4gnBCezxYQxtI
EvZsGontkXcKbWcqn+RlPsgLJ/OOIwV1vo+fMbkjz2bV3PYwAexWOmawzzu5Lbd2
qjDsgGsQ/SJ9wVU2kZh22lGXW0ir/W2X8C4i8XGK7Tl62ZhqqLkMnVXKK5z3n1rX
JAUp5NS8rv/08elqmDZ44LGss97xIjqi/E037uCVdeWDzJW6iHtIbxn8cbBlomKy
JAbCDn+tbrCnkcWK5HpROD/3NJw5vMQ6VjyAHG8V07M=
`protect END_PROTECTED
