`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iOqrGW5L2MpD9xL375owC+mkfcatLS1MrEpsjOJ8JSlR4qzNCmTG3D4NmKtAc3do
8os6o7nRuaSHZXSguZ/mJajOyi8hQpB8EJRTX9z3ywqgMWUTe4mhDw/M7z77K6Zz
CzBL46lvyU9frxC3XZ8UpQHE/jJZE/dPRXtorjTNxI8WPF8ZluzC1HaA3S+9lTuz
8rCdkXOhKSULAnSpk4gvqcEPdFiPTF70uOqdxDUIxmEP9y4O5lRyVxMbV8W2K4lW
JHCAh8VuciSxEJ8bJdgqT2RR/WFj7kJwSeOcF3uMP/ouus0YKqeFy5XXrkJngfiW
ZsRPGVQkXhINRzL/Q5qUNjSbIpcL3X4pULstQ61sgck12Jy6TteNj0jY1yxI0glW
eM1emMcOXAkYrcN8/4JmUJxVkQipk1Cj0sNdV/fVepw755n6m5VA2WgzdoUH3nBQ
tCjUOW74orWlGenSf2N+pjNkbana11AvA+hWTRs1TPoGCQVeJkM+Xvt1sMsxqi2/
hmHecdERsPNIu6VnijFHu6LPPNTHwPI2C3jmRDARSL18atHPIfFVTV7wAQgX1KAq
t58UaPpjpVhzyJHNpj6A93nUD+BW0ZOHvo5QntEVKBRIveCmNqQXsXE7zLOnuRls
FUczHi2OlAB1fCafs0vis4paslYynGVEudMFxSiCaPFLx16TyiSU3342QLHtgSdg
No6kTvtPTmMPeehxlbbI8skfXyEVD/QdVSiqvGHZNzyAB3zeXV/gvp/YGFLzNISB
Bkv8kRDUDIZNkQ6VpPoFsAJAnLdLx+2QRmQYAfmt5X8vdY8r81/JOHdi+cEcLiIc
V9RqI47Euhb7g1dS2gXqRu1RIujEn0rrdC+ItedjLpwtYHfL2FTvXpuf7Y0lmcfv
Uu7EZ/SVqxJmgjtL2iAF28U7QPPbm+nCLB16d6BYnfjZeK0vIBCpS5Z7wW3JqcZ5
4d5vEMwPFBQ2nBt7Wsk7+bTtrPvzkGC36Ez75wl1fMDwe/jkEHAIcGr97+k95lHL
4cvXXs6Iw7XJU5upjhcedw3z2azc3+Li8OQRtYDgB2mXXe0ou4omUItociQYzt1P
ip/aCcAOapz1RbGMmFzTIIKjkH5Y7JFD8y76aI+G+rfw6LVF0IaqofbAs0cyMJN2
8qb3iQB/EA5murlLEd7ZrGRSdnGK/lCRdUVkxRfhql0j7sg/KgQBfH1V2XGXNuJD
SapYPSATlAAfhHiIJMEJoeWL8iaDWzCkO8HO575vYafZfvyk9huhgH5RXLMn2owR
uOA/bJB3disRI0Is6oMnQ6v4x55YZmA7B2xIWqbsyQZ57J2Nc7LWA8HdMtmymLLA
dWhOrBPgzt4fOg9vC682Q7bkqzIFFDz6R8aYoReoFc6W2yTT7P94poBPWSxDimoB
xo7ZOS4G+A1hOaziNoT3HocH3Nf+1P1cX16iHn6qMyJc+oiCvhgDmX76IHGQuT3n
1uyx2gjfal09HOo9Vn6bzsdSGsA6iQcXRyOMfDQMS9oouAOPJ8Oa5tIHHVU8DUwZ
VmpKLciojVBePl0L2V3OZcrjoJDXE1YaG1Pk8QhIXb6z24qnkCJp3XSdVUdf8Wml
KdcE/oW4MX/QWNbqkKsMWRBseQ6E6awFwHeaXMc4TyZP1iRKgSx5A+gXFE1YIgAX
FKPMU//SPAz+hm9EF+C3jN9fsHA3LDDaK3Wq22dUe1xvQXmRj441ICS1lot8S1ey
qUfgVmiT/iU9x9XTV/ENGR0qJr7Pt/ugw00R/kqLl5KTiPPGNfmkT8Z0q3FY9qsK
3rFo72N35Zs4W7GhoRPUaVI2PaiyAOALN5yWyvAWa+9TAnYXFNYhlph+RXy7enmz
ruB4BcaMevW50fCjSiHf4e9JGMnyGvzV3UVq+KKqvcaKyXaP9fXg7ASHGHAV+05+
W1v+6EX0cKBGuNID91x8LcXnAp50ovalHHu8/UbC06qM1VhsHf4cy6np74GzIAvj
YZ4lucEXwvjXt0UJyQrSys9OJq9arzDXixvb6Uw6VdS5szTgLNyx/DUjXjGttDmx
JhaE+6J96+bW+/ONGpATvzBtm3eWyTKPpa+cUpiy2sFJPZWSpd6zYueub9lGv7yI
jCEpwCutSieGYTsLtgYf/gd5KVulv2xosWHM7vSxtx1anjhYWLqTlrdjwuu5Beop
aWpnlxHqcpRYiSvtM8/2KoSrBq8jCB93xAqiWvjt3olq+iNdm+8R+Av/8Jv7nMxX
q0jG3/mzEZenxv5esspOCPUWis2cmyVCFjcMivGpm+ioIG2zPLKmGqQNq70mmyeI
y2Q1Ra3wdejYqIDDK2J5TxaMroNutwrjWwbFrkAwmLRu4gvmuX/i9It7RvQ1uBl9
ek31vxqYBq4oLwCiOoSjaiJ+WyJMUy2EzbGfu+SqjDphrRLuxn9fNYy6CnIOZJa2
`protect END_PROTECTED
