library verilog;
use verilog.vl_types.all;
entity APM_H_UNIT_POST is
    generic(
        CLK_OR          : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CE_OR           : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        RST_OR          : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        SYNC_OR         : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        OR_BYP          : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        RTI             : vl_logic_vector(0 to 63) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        SEL_SAB_CR27    : vl_logic := Hi0;
        SEL_SAB_CR59    : vl_logic := Hi0;
        M9_MODE         : vl_logic := Hi0;
        M27_MODE        : vl_logic := Hi0;
        SC_ALUEN        : vl_logic := Hi0;
        FLAG_EN         : vl_logic := Hi0;
        CR64_SAB        : vl_logic := Hi0;
        SIGN_SELIR      : vl_logic_vector(0 to 1) := (Hi0, Hi0);
        TERNARY         : vl_logic := Hi0;
        MASK01          : vl_logic_vector(0 to 64) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        MASKPAT         : vl_logic_vector(0 to 63) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        MCPAT           : vl_logic_vector(0 to 63) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        MASKPATSEL      : vl_logic := Hi0;
        MCPATSEL        : vl_logic := Hi0;
        CSIGN_EXT       : vl_logic := Hi0;
        CSIGN_PRE       : vl_logic := Hi0;
        SEL_SYO         : vl_logic := Hi0;
        SEL_SZO         : vl_logic := Hi0;
        OR2CASCADE_EN   : vl_logic := Hi0
    );
    port(
        GRS             : in     vl_logic;
        CLK             : in     vl_logic_vector(3 downto 0);
        CE              : in     vl_logic_vector(3 downto 0);
        RST             : in     vl_logic_vector(3 downto 0);
        CPI             : in     vl_logic_vector(64 downto 0);
        CPI_SIGNED      : in     vl_logic;
        CYO             : in     vl_logic_vector(26 downto 0);
        CYO_SIGNED      : in     vl_logic;
        CZO             : in     vl_logic_vector(26 downto 0);
        CZO_SIGNED      : in     vl_logic;
        asign_ext0      : in     vl_logic_vector(1 downto 0);
        bsign_ext0      : in     vl_logic_vector(1 downto 0);
        asign_ext2      : in     vl_logic_vector(1 downto 0);
        bsign_ext2      : in     vl_logic_vector(1 downto 0);
        ar              : in     vl_logic_vector(35 downto 0);
        br              : in     vl_logic_vector(35 downto 0);
        cr              : in     vl_logic_vector(63 downto 0);
        mult_a          : in     vl_logic_vector(45 downto 0);
        mult_b          : in     vl_logic_vector(36 downto 0);
        post_op         : in     vl_logic_vector(10 downto 0);
        CPO             : out    vl_logic_vector(64 downto 0);
        CPO_SIGNED      : out    vl_logic;
        DPO             : out    vl_logic_vector(73 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of CLK_OR : constant is 1;
    attribute mti_svvh_generic_type of CE_OR : constant is 1;
    attribute mti_svvh_generic_type of RST_OR : constant is 1;
    attribute mti_svvh_generic_type of SYNC_OR : constant is 1;
    attribute mti_svvh_generic_type of OR_BYP : constant is 1;
    attribute mti_svvh_generic_type of RTI : constant is 1;
    attribute mti_svvh_generic_type of SEL_SAB_CR27 : constant is 1;
    attribute mti_svvh_generic_type of SEL_SAB_CR59 : constant is 1;
    attribute mti_svvh_generic_type of M9_MODE : constant is 1;
    attribute mti_svvh_generic_type of M27_MODE : constant is 1;
    attribute mti_svvh_generic_type of SC_ALUEN : constant is 1;
    attribute mti_svvh_generic_type of FLAG_EN : constant is 1;
    attribute mti_svvh_generic_type of CR64_SAB : constant is 1;
    attribute mti_svvh_generic_type of SIGN_SELIR : constant is 1;
    attribute mti_svvh_generic_type of TERNARY : constant is 1;
    attribute mti_svvh_generic_type of MASK01 : constant is 1;
    attribute mti_svvh_generic_type of MASKPAT : constant is 1;
    attribute mti_svvh_generic_type of MCPAT : constant is 1;
    attribute mti_svvh_generic_type of MASKPATSEL : constant is 1;
    attribute mti_svvh_generic_type of MCPATSEL : constant is 1;
    attribute mti_svvh_generic_type of CSIGN_EXT : constant is 1;
    attribute mti_svvh_generic_type of CSIGN_PRE : constant is 1;
    attribute mti_svvh_generic_type of SEL_SYO : constant is 1;
    attribute mti_svvh_generic_type of SEL_SZO : constant is 1;
    attribute mti_svvh_generic_type of OR2CASCADE_EN : constant is 1;
end APM_H_UNIT_POST;
