`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kl8SVR+wUQyzJIbFbzTvqenxy86EfPcRWwcodvjaAMsQvm9sZ4IhwujgGW9scvZI
x8bizjwaTbU2+rJ4jyuGT2t6NJtenFV78ewCt/ZDAgriSbpiGQfvlSTk84gm+xuf
aVx2KJ9ncHI4MDa6UCgVZqMakal03EmG3akCSjQiaIxqjdlG6lMXnul0BRU3XUOj
Ml6CQhfU88TnbW7ou0wd0d8r1i8hTWldyTHz/3acA8qPUM+Fee0GtoFNF/sLPncC
QqoCXkb5RuxWM/ZQg7BMvMT85SYp+pdNTCjZHQGwRpUfQekoXECsBegk5uCO2Zyt
5s1D8CndPAdtsl8v74Pim4Zfx+9GtohLNt2xm1MEAVVmRdFBanlFGcff/raRZIbU
ExI9XZee0BVTKSnONp9pr/dLsV8/datvyGc4J6o6VTjq4yxysaurV0rCwLpZBCyi
A4ZnLoHJLt4pPcF8qbk03pXZonoAMccDgSEMFOVg3flqwgh5dufShPsTpS+1O9ra
6JfXXJ0qu1v/1s0Gf0A7rsa8eVRBOPozQUrom7qLP98Z69iBcVmsOsj3sKMEngxf
oUZlar+/Sl+0DLjrqGjqOtnfeKIgmPxXPMoCBuUwf/bawVCkWxdroh882X/WyxUf
Mu1vCViV0cLUCf9rCWMxWPoNn2SIqdedimOqdi14kLxnMofnRuy9u+mDDSbE8L11
3lzj1ae48RKEFuUxjUG3l3pXNYKzg2HasJdR1hTIIfxHapFK7BmRBtV9vdmPDUNA
/AXuVLjiGd8oD4BGkM99vDEfMBFkb1CC7PpKKevvN4DMwIlXMwphJPADijdKjw64
MBTvIxN6HjdvJo8KwVggUgpnsJejkDoxPPRAhYkaUTrL7a02Iz+cUpqv6Jt67Dc3
gxJ6fEeDKbtj5yaN8wShw7/RjYFPGMYPNCxUKITP9NmHeRfV2gbiUmInZh6wTEG0
HvmeZLcLEixToK225vWN8yfYAhp8PninENvNCQk4EQyuOVgXj3RGPrdpgl6zyexW
wdBeMWI1S2JQNi1C7IMb9CkdhHNeF3ez9FPxkVSyYDSOiHK0Jte1DfDqaGBqerE3
PCf2FvE14ZLJjGSOoEAYIG5usvj1FEvP8/atvE5NJ06yfPbxSIKLzCCeT6etRFsm
pqofXI/iUXGIWDI/e8Qj43ShZB5f7RshVPTeQ3Bf7IeDNDpWjI85l+vyY/8yWmIo
L9G6QW7J22BY/JUva//vgc1yD27s1Czo1V51gvI8YmDgCbUz9jFUyK4wNklwta/x
IEzA+y9mSd0BDKDHnXAVF7LInTdmwVzfBABWwMnR4Edx16l4Xs2xmSFX4VIuxwB8
IOc3wNkdWW24ZOO9rNMeX2M8XtkgQ1WwLPTj970JbY91rBvuV+1f/cnEpFHqmoM+
wUtG5Y/vM8BjbJa/hIEXplsd1LYH41P8ZGdz6yq7HWmaLv+f4NMYu8PMRmhXLAYn
eXi6VB7hX561KFVUrMok6qr8Lz7gTQM7yq5ZpiOqsBbbxXSUDrFK5lh91Fvv5bUS
rNyLiaqXBC5lPDEHL8sOn94ydmUsrbFoHNWCzpoyXQNYByRfoB6ZDCVgY8IKJrt3
CIkJ6r6jDHV4k5wkuLlTfcRVGPBSHIe1dyutaSAPwL3UFF3EJ7VR10Cva4rQxBSD
wRRoz232+ERaSaC7fai6E+5a9IghmeCZ5+AuaxnIoafcGbqvWOTqHms1NYkZ6YtX
JslysMmlLBcsURmZ8zIyu19XaUCfXxNGT3BzcDE+w10oXqFR0K0kUb1WyhlU8V5r
hz22mNfq4aOr9ReNLjPn+cS1absZgg/3lOvBqUSeQ3yCHY4n3qzCu+OjLlIJQQgO
OnWVK72SJwrylTSyE2i084uKlsauY2xwU4btsFgeyuJ5q1LBLz7cEgjvDD2mmmmM
Ft7oQoaTrsnABxkInP+Ec1azAaWd6we5SUaGvWr9n1zN5JX3RweafpPPh6iZ6tOZ
8Y3uZ6Tpr5QD4OcLTFr8rDxznPNPiuFfoZpfwSO1PRqcFT+KZfyBYpaqlwOnkuC9
TAuLH2bRhpm5hoUcglU1i9cAqLlv4u5OFwUIRoL4V4dLclODDpDrHOStYqIrgyJA
yLdmznc+U2WDgYbMzFzdfgoQfCuwaKhp47jYW0FB/+7CYi/MaSfpaZPBEhgcL1kD
T5mSZdQUOO8W7HpriZgFZ7dN17bx8VQ6m+EpyJ4MOcoMTvjkPctPSUMHD3IcBT5+
OqEDHwwAX5FgqbMlCuC5JB5iGaCYvi4G48Dk9DOqDR9A/UJH4Kw68owTshU2s2iv
ZjTcxdYfbrxbg8EXKGqI5h6cSxjgebe8pQI4pXlHCYr8c9HLyGTw6W3F/CAc8IyS
/HL74+NgISr7ETnsJox9+jQVo47sSrPwgYb4pu1S9Qd3C9YWGb3YSnnomPzpdgHJ
jUnmcXsCC7XjpXIpm+kxpzbG+bOdr+H7OwKbbLez1AriWJXO9X+Hu2C0L8WNlRMS
YoP6lduVffRD64Zs1q5SRc7bQdFlpi69xRsORh4VISFU2yOx6ixi6wUzXgRIsXZp
qn6peltaGh+ev+1dP8xiIb/v90KAN0Sy1mymgPP+XHvVcpf07K5YjxYMu3m2RpMe
hjtegJYdbCIgpritKkICiCPBj3RXLzcy0Wn+RIlAvz5/AwEZqrsZVnuSZocvlJdJ
xUwXIIg4vSo8TsYqlPoqQugig5xj3zAcguxQRSbN7f+CxVGma7j228sC8a/S4Vv4
+joRZ4pWhWla4zjKQXoFutl2Vrnst5V/e96+pPK3qomMLomXa3jEeFZvkG2Co2FM
R1sdEhK1APzZHsXIRovjIoyX2mdsdPoVzMwmXl2MSA30biimrAok9pReXVTp3YXw
NaygYtTQ/0Wl/pF3lBGAyTy7gcZZ0eI/qetau6Dz/B2eY9iwcSmsUc01I4GpUrQn
moECflaQ4OAHEA9TTHLPQSDbJVqX2OuCrb8dvRPNcP8ASpuAmbCFPcNOUecqbNoI
iNsQM0qU1+FaGXnO6v8mFLaQFuEjOhuzyPJ6OKKKwUDEWnZuzYhp52V3lj3DPSf+
i7b7q4WHv4r2JJH+jdykI6UJ9iHgWcqmJqQlcHD0MgerCGt9uK0fPj0q67TIWYjW
DHtnlVsEJ/eq6eM0p6VmAWBs3Dvt6v72ZnBvA2j+LYFp8OMdqz6oKgPU8MHtMvGx
9WCUYQrLkXLrfO2wNOG7iSIEKEROCcgCT+xuLPGNiFUtmJR8F7CKkFoZKp5Ik1RI
cc1KgbAInPKP9D/jrHDn//Y9QyGSpa83g8XmoyyFgkN4Txbl/r+ETtSLgaCUWCsX
DbR/LdCSDJXxSjMZ8kHJjrjh0+QIQwrLtT2ZWVaH2Qko/H2RN1+i/kAqmFxItYWK
nCOg9fkylI68YPWONekxA7UYb5/jqkXxmnt5WKoBOfTUkW+Vf97rCAoBWS/hkyLC
jMeOF3tE4dF87HvigTcIvvDx+6od20PkVNywH7gyxKeC+EbzCG2GjHWOBR3U42F1
tWGjPkBz6Xs6cj6j1FNaQo74hAsYMHAEsicG/mZU743/vZWP+K9TDEqV2VepStam
TozWDydtnhA8k8x+Ki5EXgNnq5v8kFNVTsKFeLkjd5Z9pKKRb3BNxXQUTyJAPfkr
UCuY5FD2N7Q0OKKfarU99FD52hPL9MhRwmoLV9xsdAOcb6CV1lnEKaiSmSKxOewT
+gtSJK2FBvhx+LCfG9xiXkU+YEOfT4NBxuXKKqHj4tBs9l8LuqLa1oXepU1KzgAx
Ez2BCYd6oinC8LqPRutI0weL5ogXm8u7Pq0gKNnzjQNBzWULP7k7b22FQdqNbwzb
si9kRcRAeV/9n5aYaRiephr2qHJmLFRjEacGBxXphjzCGqUuKOHUypWB6Dxo4rS4
eIFPZuJJlIckG19jLG5qL6zadJSFhEmY9K3edYYcEt0QkIjoErFp60Oz8+WsPkso
alEXjOVKiPOEWGDNxp69gvEVCnUJESzK34QEkgJLlkWWljJ7KIEMyT8C1AwAB0SU
weoAIgK72fizCiNhKG94qba6UBRTG2Cpfl9qqBEjZBcyAosKXiA2tzMk1jHP9oxI
xuMb8i2mnUoWr5pOcJFZZ3TQ4h0tt7n86pFpJ0qz9GDoCwERG5SbeTl8iUvnnYlk
VuKpVSe/uF/1Uq5SRrNOItuDIwSo1s+gr5V6Nus2v7UvTW3NudqQ19ekXIqal+1F
n9wZnKFiqId6kfnU34edMXBUBvfW5NwlA+pmjW1HEuEn55vrnV8hrfRWplTnSV6m
Su9684ku5Icd+DT21dVDCu+zzS4X4pt3AgLs093uEnNA7u3P7GTjsw9bvSKnhzu4
EcrVguBZSjGT7kGoKZrOwYcogaKOux4+Sugls05VbeIgHL8jPyRVek+sAFbzXhZP
Xg6C/dhSQqF9Pg0mttW8xNYZwxRlxIErRZOo3XNFrFJ4XRLdEuKglA+YGg/XOKdX
KrwWW9RnyLoUE/COfs9qSZ5jB162WkTi9RA8SZwApPRwzUGhQb/re1H+o0R4FEnY
diGtMl43zTTBjAVXd/GLm+FVeGaX8D8Gju1/tklkVD/tmGd1/r2/5nxuDqlWFdTS
bpI3v4dPb9IKYLNKGDQSiiSD33KNBdf2SlfYI9KFUfi3lVo7X7iKT96efS+VPHp+
BTVT4cfZU4sNacBYoSYRm+PtggVGxvtQ3QS/QPc28nqXCW8E9Y9/xR7UMr+TvBKn
ZwRnn+9gysVXwt2FfiyiwpjPWe+dswijHvVhAr42GxwGXiTpqs8cx/9bKBwyDo8V
STzXON7RLBIOK3Tx+lq+JCrXoDov+EfVQIBsWUtUBxKvwG5nYN+zX9tqu50Wkq5W
Nm06brXIwGDLHdRbIO0p01eOlJGdbVDUFMkp2wtSus4D47HwcomeV0T/FiDXrupA
2fr9aKEUgUQbrrPKx51N4IHldLiY7j+HxljWzGfcGg6nTvHhweDD5jNgDB3MEfSz
84kGIXFKLuE1anSOgjuB7hQSWzciOU0fOiipk9pbp29ILvb1LsgvanQbQlZ27JzW
e69mDD7CaZoJQJujdJL9Bu2NfsCIqTWue7lR05jL7tuf7meLr28+2yMPyVEOSyHd
4zMhPP5IcYYbc55bLcKjYwubJ/ooT/G4VTH2QbN2MOyIwIlS7mczTSalFSAXPixx
KdMaZFbmBMx6AZVVnxUBNgcF2oWv1Hqf5zC0k4+FM/4zBAjgFr3SrXH3RpvPKhZx
SBSz6WLeL/UFB7uGTvytEQ5cwF+1VUtY8zfKoQ/0R2/djT0iB+EW94uO6TZPbS3h
nhWdgdueHjz9y/OKcyqFJvXvIru9yVt2xCNdevrzS8/4agAfBm96wKvPLZPr/V/i
SFnBdlr1O1oJKKr+Z954tqWUzHa+RxdCrN4WQF00RyNWTOSKby7Ba+nAkBg5iSsM
jx3yFkdxVL1M92iqwwQ9qX6CalZYYWmz0l+U/jglY4BB93Hq4zwNhhVcJ8WuB6YA
Lil9mMJ28v9wz000vgcVU2eWGk4XfIXpxFeAu2lXAGjIG/9MUu7rudBuxcWR1rnf
Hpnc71AR08prF7w/CLlLWble4lD5gQXzEe0s6kt1waqFGWjxRtUOtmV7L3zIc+Lq
+Qd6LtJzTPKzaGuecNuIVUrHci08mDq4npZkfQzMtKT3lCyXygzoD8pmBVlm8voN
wlwv18PWl1xzhKHdvonh2GStxbOWWgdmAenbd+qNatrwyFEO02Onpjl9QRgYPV2Q
omOF1pcqkeYG/d9Ysb46P40VlA4RZSFOctS0SnwXoLZW0Fep/BOX9vp+kjaLBerQ
3j5U+A7QweGUnOBpbLciMPV/pg8d5kELfBzwoilrjMSWWEzXAoejpXmOJuZQhTxj
axuVjsd8BGqdZfkHhq6l+rPyCXV9lxYLAExylaeJ7dCp/abzTeBbF0xSexf419sk
1noLKr2WpDddiVgj4DGJ2TdNIEPjWz6WAhauNNULLnkiF8r5Lq/UXcVRfZpFLJZJ
djPL+iEHWzG+mt9RvHLPJBzEr0lvncDmhHYqGCJokb1FF+EZkq2nxcJesb8fxUU4
rKR7JUTSjJqFpGPWBnaZ3+8Z1Wvhl2tnT4qIWRF7VaUw1thGYtyjtSptJIprOjAt
ghYopN4yioNz6MAF2DiCrJP+2nF3V8akrjfj85XkIHd8E6dpeL4IcYXG/4jfmQ1o
davOKUNVxRiGXD6dRpfGJPztO19Mq1Hi+3A+DKFcQW638x1NCzCQgzvcLkVVAtfP
rZCaIV2aHrzVrb8qNzUY6NZuAsckZRe2GBWreGo0ftbWsfCauMZQkR16Wo1SMhbF
B+VnGd3LMSCX8+HUxNc+N4WZgiyUmb6xGt+d+HXSJXkhCRxCaEeJsMPUkg/5G7c1
xyQwY1nxZz89q4E8t7MEGeS4JRv8jUPu1VTZzmOnswYqvYnGhPTPHRvO4X+BqGyv
tb0J5u07ljsmjilRon4JatrmF59729hjxtdAEh3DQ5WFxpjlshqD3R+Ejv2CwmiF
zGLEpavE3PMYC2G/DO6tvoGc470+Dl4VEsahknz+HZPuJm4xj5NrZSI62OoDTB0Q
/OxIcpdqMuvyaY5PONJ+NMwSTHOKi1eHZEaSw44j/6LyOnHQo7RAJZRSD3RILmND
j/69tDiHkoxscQXy0fuY9dXhqDYFrYb6zUbUZn0uqFC4o5ovvffibAoXeyB1aM+p
Bf9tW+TWNkE06kAl2E5M6sYq/IoGw/rLKrcHh1NS2yUtWDTV2NSXtv+u9YpCd2nE
/I9AcgxVmWmNRV4qyKCwHEMYP8Gnzh030RCrWMmQN9Ug0Edvm78zbNSWJkk8Y/8u
TIuu0F45+qgvybgj79M8cnALcgVcan7i9NIITXvp9y/PWRybqk5N7gvAxE+UZamQ
qSMQKwFpA37b9gduWQnAIcIVILu6uewdIotgfGVDoXIOMFl92XcP58p6fuuU9wd3
8wIVm2B/l8lNA2TxM4JJZeXUksToLzMctpPEBbcPAJxM/9u+99AcP/tXRzmGqtwF
mDPok4RzA3vom8XGRybqOnW+4UN2UBHrB4Y6cet01kWrvtYFtzL+IlNMPl7239W9
9mDg5bDnXDLQcqs1IqtU6YC+vNE2SYpqqelRFMLsEZCtc2jq/quHzjYuNq+agVrv
usUzGUzFu+jgxI9X/qdaO0sm9AJZ3/8KtgXGp7n+pHhDyx4kqEJQz7yNMsXIH8t3
UuHrGu1jVD0tZNcjn1L8NgdzhkpNxkuZ3y0mIyqG3KxqvqPJ5wZIad2iwUhr76eU
uRpjGF+5xvJVfVl0UNMh+Ek25TTFAzdaaAHQ2qKGFRDrSZ03HfoB9iF58tYoKBol
lXPTa8vcfL7Q2Uk3zTM99EJZ9ZsDEsxVnLlqmLne27ZCpJLQO2HKYveczdiInvZf
L1iuSlLKptAbFOtO3iSP3QzoEzymWQJ++Dfrb5fWHCCS8OcFFB6uK6i9XxizSZ1H
hZaZ7XF8Ive0ltA4A9uGfYv244qpbsZNqOVk6kUwnMKtZUL1pRXaFQVKyx11BV4Z
ynBjzw96WGaS7M72Zai6G4aQ0YCn6luUyEgY1bY97gdP9/daLhO3c0OyyUum4oiZ
hvksYRhaiwUPKenP9L2Y+QY9JEE8Ki0qrbv00e4HcgV3EvoIUMb34BBI1l75XJkp
3kG6hrrPZYfosmjCMtzzAEJmhAlnxtxxqoG50v/U/kMA4QYGuX9MLO2uCCDVLm8V
7vqY+dYS4EAQvYlx6YBm8AErloKLl7fspz5H4AYXeBWJT3BRFmSCWJCBknwG5fC6
lMabNQB4X7Dld1/bsSXUgQsorpKCWq7npIHmF83RJ6Ev3uR8UQ/YUYm44qw/KC/Y
yTCxhfvYRooF1ZiE4pUCBL8rWobLN2hgCe18y9PGQgV5/nkkyTUvwMICsTHYa9Bu
WpL4UrZVuJCWxYC076P4TOqi5b8PUI8AZg4NNTAOwZsXnQRS4ogexB1UOZbWQ9kO
bHdYbSGYQ3mOIi+lA0FnUg7c1I109pZY3C7m7EbC1nHud9t06U/rEw2N+ZY1ZehT
2rR6wv+ArzzNvowIevNmCjA4ZOL+8H7S3V0e2fmYRbRB8bNKairUHkw6WU/2X4Jq
CZI8YFxgfiTrUQDDlNYYITcvLAuGMn/81OWjkJoD209nhsVwXWBRgyCBg1uyi/Lc
omAZChmDznZgt8owq27aQ5E3Pu+47uvfC4b2F03eyQ+zh71oOQ0uUYs0pWMky27A
Sj6xofVuQEuIl3d+Kv7LyVqotxN3+EUaLI6drDkf4NUuLrXBxU307nKCHK8SsoBr
hsUG4xGkpH+oma91bU17lDAKa5529/sGVzZxU8gma83ksNuhIukOIBX6BabaJy40
OOaszwxI2Dz8VSjIn/IrpjzGR11zU0sNoK/WDTR68c13imyRxeFUwuM3PjdD3oAZ
Y1zc3cvR0RpRXj84jzG+jD/7+sQt7VOq8nCYnn6rhcLuCyYO8YSn3LXQIrMWzZsl
SE6rsYZ5Mi8DC+7JNl39UOY9ixW9wEsbti3mrGgASRl8eUu2Sx+mDwt2AxKd7+Mo
DdFbi21XqA5tNmWYqcfCMgVUO6h0QLjgHwAcBrMaIFiQ3ZOGnAGu5TvT9/a50ssc
8vixcNyhlbLHeO1zQQPISZ1ugnLxXsUakqFG3vl4r6rD72hE/cDOGrRFPbtJi7Qc
Q986Gqx58IPGN9e3VT6yk/qbBjXeYCuNIMKQLykjDlvmwm+Bgw5AA5Jet6TqxCcJ
clBK1RQ4cFbXfDJojbQZKUwiHtcIwvcRiEkZjBaloU3ycqfRMq4nMMNwHSjMY4df
G5bWuGSUumbnS9FnTqO58gCvgSFEKa+WlX9SAR9+Ar2xZRPicNx1HU5Ggqx7xkXD
BwELYO+gz0LWpSyqGd09dfqINJd2dQtenjCqUpmNhdkhJzUd4TV2vBDRKF+TapQg
w+SQ8xtqELTjHKpq7Mk9nHkR7wc1pcBDgtRlnLv8GMo1BJ0QMJWjyG8sKGh70ZBd
nBaEgKYMj+m/6FS7ipc5kpb1Og8iKAuM9w+IjpujIoOypuIT+eyg8KfbwYT/Ba99
FG7ZQuS87fqSiT6RrDMy1/xj1NPdH4S7TZjnhJUpoECic9Mt5gcMvs5K/6Un4TKQ
b3/9pZXQUvV86JDbXwmMvcd9BHtiLP54B91rffVmRQHeGYHkI1VDtGrV7TF/jcqC
rC59mUs7aTvm4BFaHn7yNwcxspc/PxmzUME6oUh/8VgoUNKAk3gYbC89/uW0gpL9
1XwMfvYNSFTP5Y6VmTCTEbKi1IDe8O7E+Y/R5EUFxB7uBo8EKz+23cSl5THiDEwc
1HSvVvUnPoUBWy0rPouBCqzEwAhjv0Gp1HHtESOQXL9ZriWxLLVAggKVmk4I2iWa
f4MwbS7cBozgqG6L5caFwRJtCtxOQUOCVbWy+C2LAigDVoG0yo5eIxbgeAmdxBSX
fuVxVud+M5cmeMagaVWTmDasUf43uG/JHOOLKR0b3oddygZn6UMTKa0FOeVJUM4a
NDX3jVeGWUnn9SxnwMv8+91PdHjd4phvO/lvlQg7WeTeiEu7xxcN//yguXs+JLNt
MjphCLTZ6B+4W43fBCzwNAXMPOMiOG9c9QFrP/Cp8/rMFkPR5sd8iTxUY9X7JZ+m
WeG4nfyWZfpwTuNjFjz36RFKxs2yPby08QJ6TPqRBzI4GFUmN7PG1NmfYMbORb/K
Q9QzthplzQMfN0xMxeGukNZLRPB5sqPTCBVrcfcSkspzRGqxAMPhMLlSR69IOM28
vFl2qsZdZ8Z48+2ilVWiafyEArxLa3oG22XXsy+hMTSckDEAJokzulvD98wJV1nF
jvG3U+hsbFhmeoyJBPn/Yuboln4RTeOHg3RcWnBZe73OajXM5aQDDn4GV3Yb3iJc
uAQ3lIgAlQp2B+axCofEHSI+zLQmtrgnotTGswkXTc37KWtS1R5W4TInNGqEj8Z6
wkemr1qhlIPi5SVzJ5UoPaeTU0H1XTrjHMZBiBsX/AyMVtEFLb00X9iDnbrQ2Bkc
1q4M3z1yFDnDBbg2OgfTT5LMkHlgy16/dDgkcYP1WYHtLOAb7tir+lLjvq3FQ0XO
g42sT+1oEBWEYZXNqK/Gz6gLwPJr6yadZ3hDPpXUXsVOI2Vsd+2iiGVKe/gSHBcq
WwCu8pW5iQsIrsyPhb0iwYyRfrzYbLbAuv05hfpx/zbuvE2eiyrantQnL52L0d89
tfI6jpsZ7bnjawpKij4eNmAcSDb3HWMtx95fHDjif2Uu6gM+euQ795TAWM79yFcA
zyUibSTJkE9dRpaKesosia/GINbozjAkhDSiOLI8bj3qx82izZoFR5d3zjJYJuRh
aV2M581cp/vn5ri2MWAVmG4zri4QVMfclBEMyf74o5Ewk+9gqB098tqQ3mGKKRjr
tr2Lq019lyS/kMnAud+8pN74v8dvM4VlczgRWbbhCGMB+wZVA/geMfs3m4rSXk2T
YjS2fYZVXk/GUc2vvFQy+I0yta0FIYPLhYhKcxktnQIaeb3tO5QmxHhSSRO6kDb0
97LiV+HDFOVQph65Qf9lBraNrNJ4xCW1Dut3pvMXyzRfw+mKTtuXHZhTFH5ABU2M
zfLBAv/8u9CIs55c0O+eWz388M4qTq7ZxasdJOSjiSBTGX3KSy6MtugRXcrQ3q/W
tw5VJtTZdCKdV9oVNiorT1emPSOqdE0hlLb5c3iv6fYqv9uwK/an3HFKIlErv9uc
xPnQr0QR0N17Xa8oaUwAHFweH5OOvEsDZz1KGLBLKmvpJAv+w/ddd1eNqhI5xHFx
mZndWJ7mBzx+2/XDKAcU6DUKKFudr09NEBIfIiJXBhBurue08o/UNrYMnd1ELODu
jpY3lLo6qihqK/Umdq4xPMKDoC8j0kx4tR0bkPWpjJ3HzQ7Qs+SLO4SoOOZW+tQB
vJcsee5tIebjkoD981yCi9C3hFMivfMvNHUBbaqsdWx/REm57EVSTY9Pjqy05Hu/
qt8yfh2zfO90jICYhqyvn0ybZRriiDmMCCfwXbdcTLXv+loYplYMZ1rG1XUXzFPT
FsCyAT04AfDu0yTZQDuVz10y2HZ1KjYdrPebsB/Z7gaEmO2cvhA6Hxn/3E9yyS05
RJfpLREnbCsHFok+ZFgNpgPIgw+97Rgx+nMkj5mwpaCfqmK8z8gzdeb/3h3ubyRn
oOJLdidvPwBpIuGBS19ql9arAZhz6tk8BTcfi5/LRKdZ3FalztTmpnjIXp2cdKYm
C3krXWRbdqOW6zjWur+cgFzMOFk/hdtPHFG6cvz0cbymtsF1HZVcpIzVR+luxt7W
d5rUhm0VVooH862PiuXRKFlwoZSGYDusFujz4ofVeRzLkYLxGtcdOdOAP5RkXo1E
K0Od3nRd8aElckMgm9X05mh89X2rLnoiyg3/HTsPM22dCZIJpioDa2gzgwRR5pU0
GaK2TGeiQzHGMMjfBLBppi3cd2lfHWG8uxNLdkO0wJKTbLVtvr03WEysH6yNXbIJ
o2fsrPAt5NdW7mYVF6BIOgqJyONCf5fWy1w8645jRFbDOJcrzQI4mM2LooBVnxwd
MMnvmEgR5ZKEqdz1DJlvlUkZub8IZU5xmr8XW5xpuBf86eau9AmFcqyKCWnMzgpi
TQY+zBPY4r+YaPKquRa/3bc+LGSYuD/nQq2RU0qcH8/29AQxQJc4cu/sXO2zK2//
3MZ0/PrEco83wKNbtrrz8TOVCL3kefAOitmjn28z7OaBqaaEiAZ3QML+o41FA+cr
Ze/14+33xfcHcaIMN/RQpVji4R0Ju9IWYZT21ept4LyxBrxF5xxQW47J8VGR1pHV
CapkqvIsqccLDH9GAJ8E4bWkQoX49kcoRyZ57KvKMWXavAtUI47adS1P5cKwoZDk
XhXu6fnFNh0vm2y6A07rgn/DlKqxxrKq1VMt4bBJM+FWez3sgx0uzzs44l1aA+Da
7rb3bubm/JKyMlu+Naxp4UcxFVUPIDvWixg5G13cEpx6sz5pwM61qvN7HSC8qdTG
1z6rwnLArLXkw/XbbCz/t+w7XMo2qVkdvyMy07o/C6cgGQ4bmBUnCVoaYMSkXUh5
YFhRzDdL3wQ9zp570FnYhxGl/+rwshjf3nP4niWe090EWqqiCWeUHXheuvw6RPhO
rtMTQXaHzcsd3l064sES2wsYNDvouF5QCwRV9xi9wt4jMIP2omEAjrNNCEx2mIO4
JqyD2OxX15k8+b+sfAP54DYxx2moeq40mKswrKX3movyVMVIi/nCK/M/VGTIr5it
CkLMwNRFFPSgtfDctuoYLjTrxgJDshYYOuwJt8BJstyJo/+9wQWSXb4WUn5AlXWP
UUzWLhRKq8ANWjCrtKq2LThbxXHZdnmveCFeSTeq3q3+M29jHWWcpg4RWlWmtbe8
+H+kE9QbMSbzSVHo4WlESvoPJFtt9GALOXaP1unKnw9xl+HRIb4bdStUCueb8tcY
R4muUuzxeufnIC/iDxv2HpMcdlBd2SCbDDtxNuMKki1Ldsw0C+htSFaQz2nv7o3/
deU2BVVQDIT7HjbBDbYyqEcM0g6ElqlWZ3iZLHfrSjkHQ1R8DQyYlfoh5eqEBJv5
GsciAjZ7bvOZEfoFJ7E2D1E0V6q42q/A0TL3wmkiFQE9EqZYdj+vrBzUYjHn4tay
x4p0ebbEdZaWAfRhoT81qNix/oVnhmTyBztTHwH81NBs9oaIVk76wko5CgJdEebm
fE94CeNTrSiI3AsgZorNS5EasnZ0FYrdEi63gcOdgVrvCeosTdckNSaLufV0/SX0
oGe0cB2i7Z4aySimb6lnY9U5HfeNrbGN4AXANqHbU9lW7HDFVqxJX1oav6J8KFPF
YK5lvmObr2E59S1eWxwl91u+DBKnH/MDi9tiXArF6iejuoylfXjGax8o90lknKe2
0gQCyZP51D2rRM1Gulu3++hMjMrc8mnL/YgUJyrYVlGwFs7+lVPVMlTK3VnSfmRl
gUAboB9re2k7dg+/nqckNpXkJWZ+hMY2njlPsmCwTygX2Jb6uBBqSwivwO+UgkmI
hXM3bMEeDu7hM174hBTlOFo3rIIQwO1qcG1vXBfZfdfOnlVt239W43er1bpB0Srx
gsq1zIllUhUtIdrK4KyDtRhALlJLNp377LSxkPQ6fSkRLxrZ0QRNQiRIqDUbLbiJ
siywXJB0mW2qMuOGhrQBDViV/IsSEUvi90pQ9sIyKaam22hfcvxgMLUQRqQynIKi
S8m2v3EOP2Vtc3Uh8rM4fbUb2FVwAS/H0X8vCGc/XMen06EicyXhTlRzimxwc34a
0XHa71kaPLxdYhUQ7+LsmCnpSBBdVDjknaZwWKm/eJ/UptB8wi4a3PWNksMAI9Sb
70eXJy/nRGBUIOk51qCOUP3BxCt30Xch8tclk0rrVTAYdhTDWSaMSdLT1rukGc1i
/JASwRH4ijEiNPNpRrJdOORVG9nGI34e3++DmIBnzo9JOasMvd0QsdOIr9Z+dCxQ
pDqsynIEVYE+D5aT8ch1IWWzxJl8Z8LCZ7zJlGAXvpgUApXpyRBe58qHxpUu41e8
2zE050POCP7VVSTI6vzJwcUaTx8YqgHC75FejjKQSbp+3vkMsParMvX0V5MOWJpj
AqBrpylesnbgJuOEXNmhFQXKIYAGbp1Kc9sdyZq93VUoQYons42m0sGeaJh43o19
FM394RHyAOK1HR80sBW1xOsz8+0p3fssK+1GspRAK2EaaX0z64GdkvhfLCAw/rJv
QhPnDPDsodr7NTyyilVRnvqzPXtYIjUm75PFFVOvhssHb4xtPcWvFVl3+KMKv2Iz
HCYLEvaTJ1YoWWQSohg/FZ1hjan5YDGNhFkfR4Y/J+ctQ9PMAs2ZohkBq6IFNEQf
vJbEE4bvcs9BX5iQDWug92FwSVAdn2D9y5u3YeurF10mpxr+1hkLTh7dXmBp6dti
Y87odpIjqvSHPoeT7u8d7f5FjKGYK/SxILjCByG5GIk8j51RKfkQ448MQGf6IySD
+YByUKhATi6MXbh4yyxdcnUSMUcjIb0QqD8axwTiLv+fA7UaQB5N75Yy7sySKiS2
EaSMdaixbWA2nHynzahwFrDzE+bgUo92vKl32ByCZl/yOcGjNqFQyxwJi95UcdyP
upshnhXc+VtI26HUY8Jj/pHGDg+mZXAbE6lKy63UfmYH//tAS3PRKlg/xxiD7aru
ggbe8WIhnc6KN9RSfxOnvJ5a37t9yOGUtNClChFIJCWsbSt0pdlwqGjDkysTkNQP
Y+cc82yzbTPtpqD7YQPXgIk+kIBIS1gmx0g4TxrQEvXFYHUcszjrY3TohAgzn5MS
v52gYlnfJ+1e3yD8EACECW9GXKNZu9PxrxRY7rhS5EWIMOYn76GGSjTJIQfGzq+i
QcUrSYp+FxvYv3rYmx4jmMd/M3H9lo2sedtWZJOVnVechIZMG9jQfg7ztdcGX1Dz
UDzqC9LaAzVk1W27YeMgy0Mu41Vh3KZiawjHf0GzxwlBQLXJsiHcTfnvHcKHgWbM
gOh0LUmmBjADqz1HHY4sMVZZObVIUz4ybwmiB9uYpBcOqIz0tjRmh6Muglgm50YM
agjHnWdMaT1dQjax5fMijv9xV7rK5xCfpw0PoVXWlszYwG9C0DhdCh7+XDcnvELU
SdgxNKaipBPu/w6qptOBoQnr1OtFtfcHkPUfHKDxb0YElFAfW8mY0snyKmK9hLzW
5iRjIBmbbOvGuQAAWqyS3KhOH2OaNHhq4CS0nUUstRgwBDX09Xn9D/+kZf4ycXFT
vy9Tov5Zr8v8kzk+62ZB1zCHSh6RdzgeBBMJ6zDefuDks2QpZb2PHfBL9F/8Cq7t
+Lat/N58j+l8wzehHrN5551hr3OlenXadQEg99lVt6o/JFb1PodyHymuEfXtxqQd
z/y8V5jrobY1yBXiNItNNocx2c4cLeoQYZy905btY5qnCLVWGUsO4OVKtn0HvmXo
S0xb8fbRiPHiKzaBuea09X53g6zw4PnJOJmnicwCeBEpl7LPo1i8KUmKc49MSfO4
kcAW1Oh105967DfgwDsD9ZQE8ZQewI9zLuMe55z2zBQ6wcm6NuCoZnXn4leIvJkf
G8wOYCgSSjv0YB/XGUaldBB67wY85ZeJLohS3Tf5YPNpCpi757+r0xFe0T+jJYdM
keZE4Tq7I2U50t2c9PuAQ56ALLm94PrZ8YOi2myVo++nYRJuxa62bkCFHE/xSD7X
TpJeJ2IHnu9f3xFrRacV46T4aE0ZWQuhMyZ3/HzwAsnFCAqryN/XBgVLnnC5jty4
jYEsFDzOBLpYtv1BsC777E+YIFfskVMXAp1JG8ooR1uBIhasHIbjzvEQZeRDEIoL
FfPs4JrSkHdZsfvQwb4jYPCFXTgVkx+sckllIRanfmFmdS7YBYC2v+9ndoUwo9yp
VDFHEt/IU/hm0Jkh32nw8ihjD9XxJoez+xoT4lJPCzePjY3rPO+Ph7H6XXwQlrS5
McfgjpB+JH3t5me527Qe8jXms4BRL2Rn3DIWSa2F6SrgePPteOjBw8lRo8kZNPW0
vOU8ClEbIc9bQP4FaeUQSCRxwJbvT2dKyBjwRUiBdSE5nr3iEvzcuUKV5Si4e+zC
ZfPMxupxWxrYvjCJ/mZTtd4tGLeUOwxDPI+kO71HwratoqOEgkM8pe9vw+Mt6913
Ch4scE1eoPFmz/k76bvZLSaul5PAUtTDaVoQyMaPTQHSmMrKPpJd3kV0et5f9Pei
/BoD8SIAEN9/yQk8cWaAJPBiBQu7Wlog6BRwu45Tu+t35HaHMRUHYPJBvAwbIWmN
5AvOKThnoZsKGQdN8LWHitZ1DXu0qWDp1cp2Sz2+bDHIlSVji7FhtOy9eU21y0XN
KCVMt0WcouOTfsXSwp6Dzv4zvM2iT+D5wPIRPNfIONoQqd4q4uZJeaBf3Ou0I5+Q
TojPwSUC4kD/POWiTYI7z+C2u5yXlt5nNvfhHtteTbWurqZcZrTzrEvUp3CVVFRX
1AXnspJpvB7fXWn1HxliuRBUn4GBcnCjqD/BBPCFpMuMqDlY/JtA2I08+JdkJJz7
TNMGx3MM8W7Y29VNiyN4eZJ/XUa5V7ZZHPtatEBOF//G63tJwuNWAIeLfRYlfWHa
OAc5+xyRnIcVNYL1+GnY5GhliNotU9VajFA26jeIo7ysAX+lmBMgggKxZ0qAwAOH
RE3qq57XZ/YAT7rPjgqGmuydBzuZ+BT9jObapAX4UyRHiz262z2SVjUjmstE/G5p
TlzSsEmRvvfaHDSE35xtIAkDvtdDj1mss46e0tnQLtGaUALj3HnpeObhFr68UFfo
bfUAjIxL3xDWM/ZFiIN2Y70r+00y3ApHOQcc+B4vFLSd0J1HWwQgN8uPiuc35Icv
NIMHFitIsfO3PrWiRiMjh9+KdNAVepN34/bF1MAWjPiWQRHUDaP4rLoPMvO3NR9z
9TBr/kK8EcmvrsI4iEgPrg==
`protect END_PROTECTED
