`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
klAhij8fkPjM0Y77i4c30WIJLl6Gh/OcGHFaio5PDYJmpPXupOKpAl9R0z23z5Bd
WswSMACWnpnANj7mBIF2sz8cMAPS6F3xyoN3ysTREPcSbqTmLazKQEwCq9bme/cI
ZADX2mn2I4hXfL8LdSmWefTlCG42RrOTWRiHlLDCtROQyCvimdBp9/4ByWhoDUW9
LnDeih4vZRDKryM+ctW4d4i3KXWHVGRCgIiNbPfeHOff3Jn/gq80tMYZ7w6upNI0
StjEnKywmGHVdDLZ9VNFKMaLM/b/knp3syrmtsauGJD3akDolCxiLjdjKad7VaP4
wiLdTYs4HzgT0c5RJ3Axl6Ve+al7oel18BmeZpOdG7bXVCTZujUvWVnZ3x0ZXNjm
l9Pa20nJnXfiQ0JnbdWuBXV2v5gBu7igifWAPzt9jgUulseFqkexoeEmZVgduHGn
KIZvyUlidmw6WoqywWPOJsSHu/F3m0cx/pXCsSEkLAvLaZSLr56KyVlUIBSQyxAi
JikD04pAMt9nxe7639zhDtt1X6N/8F2FUoqgHf/b4/Z7yCQxcFjk/2qqDGaz/rkm
QmTqH+qn5TJ6KdQFqOhmwbX+Wi0gwLfBoH2VIFbUvJ5X2+E9DyP1QrKYXgVlWv2B
boJBH4cW2+5ALgTYaIfxGA==
`protect END_PROTECTED
