`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lmzfxf/gYxyyzHaS+KW1qTXcav9SLaxEJPiUTez+p7BIswInHyldxlRGSfqKRCkq
ep3B98Wms/g1g0+pu73rHoz8oykxRVUGJud7r9EqXmelnQuqbGXD30BKG6GIxdFK
5Qunxiupt/5w3X/eArAAmkZDp1RP1/bYAywnKmxoeNnqp8h5Vni5ymD+XNtLs29i
kl55udDvwcEK2u9xtxRltQJ60rRh2SYL0TgvrnvuzoanHc0bZrYlOEwK9+X2DzrC
j0UlzImUA7I/5RmmX4nys0xI02lIy3txOJ/Zm8ysxDF6lonj8qWVsPLFG9M27yIK
r0J4MGCCnfcc9h5x6cBEPHj2nZMd5ThTtNw50l+dEnbA1e6d8rWALQuSbvtrYqw+
J5viNKqPOi8uOMsnVk8Vhq1qswhRq2gDTBZmoMIwBWf9hQH8NpW68c/vu0tUj5U2
/zge0fNSetVhBFT9nJP+BFq4jVCVNRxi/kNTNH1legSghoXKJGKgsJqFVeNLDX5l
a/d1Q4OQfVgbgeVaInglnU4k1ios3PRp9KRIqOJ01yIjAYawf8FOfcEYAdSna2AO
jtwNs832k64XjVXQa9llqJq6w2QuWv7wJ/R6NEL7kb+A091Ah8mjxYVvWzztC5H3
4gMgBZqITt1vdfRe3FPlGa9/eYcL2FJ/VfAik9oCi3+lQOtdJeoa7wur9ZyPsrZO
pNxHqNbVPa9eFKIwsQxCIPeI+AHM5z4ao1oXmjzbt25Kzyed9HJce2zsXCOUw+Nb
ePOyUEkQG+9mbxZO3zDun2Rc4nMQ0KiKC8UhqKUFdsUVKjwAeDk8OErMhhCTdzAZ
IikMUqO2bT7k+0XVwLOHIxPTQ/3rsfFhc+8rzqKDerrfCqdaDOR5v7PReJUPu2bC
+I9uXjsH9Z4GGd2ADl1qYkmClQYr4OSr7i20XiLECuqzP/xDvgJtFoMfct4sl0Mq
ZzdKZQyb7LG8eJ5rQ/uhmCNuw6jod73nUJKKKE/zlB2NPszZ7pLQKbmudLs9OAEH
By2RgBxM7X0kjhAf/Ip1aI+l1Cv7wf09lt22czz7rXhtCeAKCZ8OWXf4AI990WyU
xfCremikVfJbbBbZYUsZjaMyuuizNMrBKPOhGALMWhD9J2CIgPq5jLSq3wJo1rKC
hMBTe2EBSoXn8jYxfyk+k58i/NK//P0z/BsOiN9T9vPQCQTKeAm8tzaFA93T9ykA
dKlsEK1KurS6qcE6gnxTqJCUtKbf914uTePU4NgD5UHirSnpVy+rH5BV1IC+MrH1
6iEm6QVQX5SeLhey0XguYe0iDClDDkUKjZvaEF1FQyOJKd8r3QP9adAj7S613cBq
dNrpqKTGf/ooigvW9SZcs2W8q334C4GaeLVF/W4ogk6/ONB/gn4j0MDxdAMCO7I6
ZXM+w9Uezj2JRQ6JQZhTsKwjs9x5rHOuy3bZTo2vTEbLT4+Pp5G+2uYbDDyFTtZo
TKcBdWUDK6scq68zypXojEPM7emTuBn/S3i4WKMwyM39bGeFkZ7tgW34uV1yIPBX
bIfKM0LcEDp7wbAJzEVe02qr39Msg3TtJgQtLbM0ib5LQcalbBS9vw5nxXiM23eJ
iBaigF8lyVZuIAD0duIKNCWqg/ztXasXf/n2XKIl2Xi68r63+9ck0Z9O5Yz2sb3+
YbqwKCMgm4p6iJdF/ntnvKaGnpBo6YpMBPaP2mDkjudXqa5OCd3y7LWGvNGPzXNd
e6eQJEyu3FrzxArKsqMAgltXIlmXE7bCk7JCePzPhq7c8yfHzsnXYJgjcMfAP/sd
rC/0G22jW+oH45rRxQQWPr6fRgd7lydlBd5UUkGZ5Xba3ZQKvFTcvTA8osFk9+ab
fdoCIeve3clCK41sF9TZBM5CYtQ9Lu2Sv/riOcqgQ3Lge+nxyXO1VebSR+cw70tx
Ok1R0R+DfZ+RdqZKlKqsEmDTnICG3RO0Bfd5cE557vQncMnUcjg0Ov5PZww8OwAG
pJOoaCfgUFjIlwesDJEGjX4nR3fGOAvDiIlYtODyGxlgKxvBmUaPczlUslfLV2Hv
+tJZJwewDi4G+Zt53fAnyiNFaGzQbdu75CQFAFK9L3DUUaeXDS4o8x4/sCamaxe9
GLgz09bIN9mraFe7mohwAI1t4kJvnRNoTPrhpmoaKNbiiNiFf4rtNMRCOOUgoBut
eJoeM50zjtiToGTUAhsKEVMjwInIWVNhQ5G/dmOOUxirTUi5jDbuPBJ9EDEzRHf6
WF1L5S0/4VwpBZ0rQ5njqA==
`protect END_PROTECTED
