`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XVv/TuQcjYAoPaWmmkeDdEfz6cPRgaBgdO5wNMBhjZuLeT/WKFueA6rH67wLvpBc
lwdjfD2hQ0lS7uWoPPK6oo/207Q0dwkTtpVRHQy3PknvxEc6dmKvV4YBRjcRIY6F
qDtXN+VQwX5TLJ+C72DEBJNKc94IJZocANdL9mf0Vi9v9e8ccJRjFjOAHHGnU9B7
XVIqybGqzaWqxggQhR38Pg7QIFYvXIaruPBlyZbP91wWSJiSu44ap2mvkb5AjrFX
oPZ5qIA63JE5vdsT6iyEV9DAq4sjCGJp+yxpHTZfnY8/QiYQ673U7TfcoP5xOQ3g
AzL/i7wrRrX/Na9Qjp7mK1292ynYLrqapPsH1HMuNOnsShjOlrxySclKaEBLeCXS
orDdoW2Ii94KdSXIJyDtLm5BUDH4Cfx43c8FLCzVKISDPSLsXrvN/3Ubp6hmwjU+
MvVaje7Sj39Of1bzPQbBDL0qfaoIU8O0ktfPrOIwvbUt0dP95MaBOXfDS2dXgF8o
prCoDMCz0ivNk1i3n+nQ8jJ0D6N/eQ3JN2OR5tGDo2kkqs3lgLSBmlds1+sexqdF
xt5gyy3e34wbx2aPEXWMiht1emlrkWIJSyI5JWB3IVD0r9HOZbXr+xV0eSqZRQQo
rFcVIRsiLLo4PpbtsLOjkYrPgHkdV1thaFbc+QlHpcrx9PJh13AqNUJmyVTGnLRw
GiSc2yd1gZzWjjTGNWvtygdldeKoXMttSWwuqnQQ2/dE5SmEBdUnaTlFy2emH5/T
+mcMyb/CapeNXyanEebQu/LAayA1qgblDm2TRrM0edtnBd7WQyT6GW9R6VFrvmrm
na0OGqPGm4Ftrx9sg4WvktCzUvPtXue2SS9qPLKoXZDIG2nQTcY41+y8MKy3aul5
0BqUXQKp11Vy1o6Lm8FMXDDhiDyG1QKBRIrDdeOI6jNXPNkV36AXOTlrM3Uw575O
ZWYQR5KvAyrlTAicmHnmRukWB3SSPELIkOyH/kRyEX4xQwTBuGYdzEcajaYDluGG
euzzLH4Co3rcHPG1UL78ODL5BWEfqGZ3tKyDjF6FnSuP1tMk04lKwjTlGIeRA8r9
grG1haPLS7FbD21Pym/FWbvxOKvLtFYx9NB3QsjM6NfU1fzwOMyWKmSxJ0cK8xtv
sou1U5xFreznxl4ZSr6sRx4tI1lmMZX56sTgEmK41GMAxwFSoueySVh1x7j17zPL
I7G40IXxtmDMdnMIGnZPR/xJs/BFchTa6nXdhZkQO2I=
`protect END_PROTECTED
