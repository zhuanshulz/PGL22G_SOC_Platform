`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9nTaqHzDL7Vnlt2ygUdFyqvVMs6JymN6WyOpKkL6nDp7f6MT2QvlADVwzQA+DDyL
eCmTRCZwgHwpQH5clhvExWzcmvQYYUTWSQtGLWg3koJ2/mDCaBvdv/FnbGRCCBnu
vyWjl1q9GS7UoYEKOGo5/FYbhEyJHXCuHNMwruPXyLVN/zNtafTHUqkuVIMRP9YF
M53jKDpzQqM7nwJ1c2MNZqXHgdMSFROEZ7tCw19v0q+r+c0HFnpK0nQRZ8WtRiqN
lGIHTAfgZ8JIjqwKmXQ34Xj5rVcx2hBFJWMF7c4mG/luDLx0yEKBL1OS4QSOTPvm
pIc285YceW8bB2bbNlWBf1RJ/F2jPMP1ESYR54gvaMc2svCPYKHZxkVn83AVPTun
UNsaTuRb0WhBR++V33ECyAcMs6Dvz72VQho/X/d+6/IQ7L4v8C60ifWV3tH84eH/
RIjaCG5dimPQt2/hy638/JCpQrlZyIeK0TL0ieGkR8nQlxz4oQDOlPwcEyqwPL/C
`protect END_PROTECTED
