`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+H0kb6rfsUO3yMQg6Yfn2O9rhu8IsLcZL7xoFOy3toe8q4NWNe3wsqgwDgxtJayQ
Oc5k5ZzdA2A0itJDRVlhIeDVtTRtwofSD43+ks85q6swrwvKkD8Fy+BRLmvj5hYd
5oewtzLpbT3ikP+6vh4x/neuTWmVFa57xjc/BiDuGM6YzhkM7UQc9KIbVj5SSmqw
romaVnoMpxuVoFy+1UnzAKcovz2l3W70dK1CY2luMSDMVW4iiVStX1k4dnujS0cS
lFaICB+zqfBgiZmfe3TvC1nOxIg3fo2OS1hL6LdX90giuDMOB2Fi6H+QO00pcQsw
Cyqvl0FmQIXG7lFOttJ51pi3PVVf3uLlmdNUJkTroZqDReH4k9v2FkQKjNaYiRLx
w3spA3BQlL23D+PesU+Kr1s6JPh08Fcczu7aVAL1WrDlwa12LoLF/QpGO3e5a3UA
BLNMfo6Z7SK6FYussd46iZDIc7hTxHv5cbA3z46G9kblhiGfoViL1GK2ry5l3Gw8
k1JELBIhsKx8jdleKMDW9oCwKABT26Pfhe8Geh+3ddB1ef/0pIcQ2keZfuK9gNVs
`protect END_PROTECTED
