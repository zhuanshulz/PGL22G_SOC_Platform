`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vbdGepcUuXbIpwJMEbVMewf5doTQjRFBbCbRMTvLBq48ArMMNFX7LZVggeZYQXQc
VR8Ynx3FGzf+tm4so6BZv3AC+U7FEtj1qTVBHfCXtuCViqBYBq89EphF0drhDJxR
i3Z6Yb2WwgXJh5zrCwXcofyscSDQqzT5FLOQh1VY0wXebhoz2VO0YdH6W/L+uxbw
3sQEDn2rN7BxG6LBJMLcJiQtiP/uJBfrBYdGhLd0/99ZF7g5zRE1inrNQh/4xePb
3ZLwgS5Z02A9dElyLDd+IoGtvtA7dmcvLaPFVv083w1cymOGrWakEN1BTo7gl59K
hAmbyG86Zn8DLGY3q6//n3MD3ZQXPHb19OuKYPwKLBwXGu13eguxCOjhnRVETUuA
Xu+0niMpig7A9YRY60K+alzzFy/tU82NGIZ1Pk8VBbygVB9oZfjvGqWIjTlyXHvC
J81wJVo+Y+TbURpqnwF4EM0DqAQMmtYhyY2VvoD3Wd3O5pIkHtb1qw1KnLdPPrMg
rQD+XpJ4V85jjw+tEB9AfTaH6hjrFyUbGU238/lTeXn9u4xI0W6VmE+zLPqqxL64
CpU/7LJxr8/I9IVZ2VwqDXgsNWOkyNxCl5H5tgqCMGQ5tQNdbf1D6qY2zQ1SbQxo
8/YJ5g4KeY/qnzWzLQOuLDcOLMgkpdManMmyD7h0z1i4nsyTDNy2EFpFow3R11on
OLkoVpvgoAHaa5Rm/Rfn+3REAFQd412vujDcj+AFv6TxP+XbH0xmRcwpOzxDh4wA
bEG0du/+Vy1M74bJQhOZN5E3/gxT32pXKYha3rcqiCDQBz1eqOPEXk6/vTKy5sue
anqR0Wrcd8UXE8UiWMEiV+2w2lRxAwJY6dnoy8tIDL0dwBOXwRGW9v8Ce2sDgbeo
Tq0OqmGJMe5q7ZHarr/gcm5p/Ptgbwm9fW3C30r6HirZOtgM3K/5pfw9GaWEwxmk
KIxbzTUecXZjDsHU/hj+UxWy3qAnbSlvH8Rw+imbGMvjhy01QcB1gpWPRJgDEkvp
Eo8iKI+hk+W+Szg5yTxCA0/5Hl81VeJS+A6WZwElVa2gQ3rkACdArLlywiNb6kGj
NvZdvWA309ESPydzNvospqinMtoC/RMzsFNhIvj0cwleBqTt4RtnExjQTuuTsCz9
PuaZjzjbmNbvPnkNuDmhLg==
`protect END_PROTECTED
