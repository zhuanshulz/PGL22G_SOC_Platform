`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xIbKNlNZuvMLH4x4CT4R+OFWxlarDLDxv0tVv260MeizuOad9r5t0CfCLlH/psW2
OwAYXNdsd6e9a2jPrWvpl9XE2G08OH6+rmzW4PgWcBOAsd51cGkUVZyq4avBp+8r
rmmXRSPWlDpDK6vYWGug2IHl/RKuHUZpXO/uPTajd8t1y1h5BCOEaqbalczpd5R+
Y8VWEVyCPrpgkIpw+mKaTKKhydLZcwMdmrJrV3pQ0hP+brMGGoC1Q4dW4bhu4ypU
AhsjWDMa04WDter6csh0qlak6l6S2Gr/uLOvrpgrfFfuPGDgCqodWU6K/BnOtqGE
uRpdxwbG7CH02tPuOVxzIkcyym18AFRAMHgsnAswYj9JEfTLghc8cN+2mvgo+cmn
/QR6c7ZYAmhTSL7YwCNG7+Q3c7vdLNaffNYCt3fE82JmtbNtBQ9jvgLx/2YOIvqQ
eKXmfNBNY8RC6wS7XEl3nvGEisGVytAkokTuMjVncgOTD+iYAfdMolWxy+zmangz
bK8sSTo1c6gJIjZu57GUNQxC8S/CQDSge9pxXv76jIl/zgqgJewDnNLgryd9KMZf
ywdRUhrmUGTdbtZJHL+LrrrU8YEMX+3IKkMhnJTlBw+L+i9iDWIW6szhHXmWI38K
0H/MPeEYrZje5+PBjDak3LDuTe9GcQwmi5hfmvRxYB4ZoCGdBct2qILZGqKZjN7V
N8U/uOMPO/fc3cK9z4spvaOsFfOaidj0ZAcL+cMFS7sH5lPVHhYsSw9Td+UGu92t
5QfG6Uq35/Xc399XLNmdpFKGSya3HXwu3KxthL2rZftdYdRyBj0+OKbyJfle84PZ
fWQ0Us007s/Kbg0S0zeZFI2PxW94Je0qdrjxF1JuR5svdiVygTsnztUjsbIknRWm
EIGaq5Jdd8MRGvOmpUrlDW5V6T+xNCvNHepTUbUINVv+tA5pAS5lfLfPBuALWhPR
FXbVtqjrFvFPZSvFifFAl3UoLH5TkMW0EsjgwU2woW8=
`protect END_PROTECTED
