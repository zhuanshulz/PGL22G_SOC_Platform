`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PVq9gKSrWdBbVAfDTSdE7fHZVRxXYYMFtM04OZ3CtPjddjPJxGdBkJg5wzfUayT/
p6aUQQGTc4e6H6WKAKXVUFAAKzb85soScYULk8j3Bo92Vu0frR61Qn/0AwFT7nV5
Ng1v1sCts7aVaiwNBWi8G80fXG2eeKfwXm7wxn0chdqa/DvnpplcczUhYEsbcMx5
PZWwold+dVFFzZyvhDMrMCXCC9qbqrJKpW4TZjgE01bP/bGigN8AXjqDfmFF6VZ/
UPifJssZIJDyh+JBrW/As2etV0p18LQ8ty1Xn5LHib1JK+5dpnI36nd2y28GIyZx
MFgRUf0fQerBtYwnBvfoIoZoaXWw1FJtxGF+bB22NLrxw1WqAL7zXL/0jlWGljHB
ZuyeFFYu6MXf0c4/hfdfb116OzFVYP7OIZwag/0AwLViC/UAv3EQh/YfFWWxksrN
K1SKw4Is7u91QdB7TiaopY2tywjQmoNZj867M7KQIgD1LLjc4Xz6hOizVz7VZGNi
I2C5wJPhahs72PVysZo7M8Yw8NmB5gVPW4nbEEWPCeU+9hxKQqCbep5//eIfvtYi
GsMX2ueTMjG0Nr+yzNfQJ9Dp9hjQtFHi4lhdKsgb3F4WmityEXTP2t1TScS3d5dW
o96l85IFfKz8pmJkhnZ6g5js46zz+PPNeerbNKYP16UThN9zRAJVK6shrO2eAoKD
ypEyx8Oq+B02iyohofy+12UXe5IQKvYJBJk3l1qeg/Lvha+l6Ej+ubXudaz19+5j
0sOr9W1MlVU7/dP3ex+0MsIJB7+LuNM+R7+b+QBG8n6IN4b2G2b2CVzaywqATNtD
aIA3o2S3lZwPKpyGJDaHWazuy4ZwNKTATGTVlYzuuFhRwztOfIfAwp1uwsvdIYIo
`protect END_PROTECTED
