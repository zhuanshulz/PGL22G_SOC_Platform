`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xNzgwKF0w/5MjCK95HosPIfcxrprBwTlCDs0nKN+tQs92sB+hC6UeRbBIB5X3WzI
ztxWM1nbIeup4/PvIsQrqrMu9zgr7tcPiV8UBKoe0sdrmVAgh9ztPxy//eODvO0H
uiLTPBpLnXcawVlbwF+YRSZvzGVJ31CBPoYl+IOApp/kzn0Ld95+T/ycr+lPLyAL
77TclXNeXmwxw/iFugFPEsvwXUVRtOoePppI+GMDfWUTh4OnlQam3RP5CwB2BpKO
zgK7HHkMxGcUkBKqXsTJT/6Rz94Z3Mn63PL+4+KsRlosbpUNJQy0C6gc+bZD9pun
WO17v/bAQumws/f+5QXOnzLawcEuVBSMpt2GAUpLOP6NgI6dZsEwYJs50aqu7lrT
PUytf/kFz6X+etcuq1XO9sHoJArphIvRY3VWIu3luuE2NkIMJG5OTRFeX14g2UBj
6QNOOmQutM4RZtkVZjeQRipA2yQ0a+eAoZ+G9ayUSOsVuutQzQWb9JuH+lUf0/Og
ZYdFcOseU+2aSnAB0Pu7Mk7dBiWLQXoW6ogZQINkXatlrJPNUMNMiYh2jLPF5x8X
ppSrlzv2+hu7te051XM+n1U0sXedEcPCLC2rN8wOS6dRS/Ogjgjm6rvB4uGIcABl
qv5yPWbOixxcW/EYBvrN91wK8lxQDIOxKWuOByBIaEYpsTvHcEWMOIT6fulPZRKT
eZeSArHFPrbfnrFNCTdYHg==
`protect END_PROTECTED
