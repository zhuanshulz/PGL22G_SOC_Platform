`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bHMsKknON2jHgHBd21cB29d2/y3fiTpl5E4cBUYtNChgyA62DYn+X9JyLkBBvUJB
pPYECaEGvcXXg3ZxxP/fHVnTeqrIlVb/He0N+TRpYt29RsvOQJOJMpQGJytPaAAA
P1jHHglncGrrk+SFMdg6pAnO6YTY4xf6m6vtqTvrWapHGZwcZlPooU6j0u1b7oc6
rTkn9EEaKqJINlQuF1dv9Hr2gboIEo4sfSmJtWiGMAlKV0fEOTgmuxAO/NuGSOhr
0s+xFxz/fOHgwrOe7fYbWXXrvLHL17sQ7euGDLZ7jGdrMvVn8XjbAHQjJWYhOVaY
Yztn3uwLym/ZRD8KUG7hWIkw+Gu6I5qUoTp/HB8hN3REs+HALna7gUv9inyKjzmE
A3pkraulj6dAym1vj6Ab8DvB2haXkourrf8srkmt4rV2P92OIBqfJXTINYJ4Qali
pNu7pAOQ+PqULNnhobRkwAQsUsDNk929q9hZdPvbNMn/2fsmei5wWiSlAINKmywz
53B2ksDeBfPd6GeYmCKhNYKVIxwAYtrD1GOOLG27gjLxeMIVw1167vzeNjsqSuoZ
V2/T28084XiZvEw1ZblDRCS1LML37YycN+rt5HUeeFUYH05IBRgutUUBZ1kWTh91
QyXGJz3Vm/0hVIJrNt8Cq09pkL03aRXcHIDkponvpu3DeFLgdNGLrTgDPsxo5emk
wWD8dcVotkQXKWzFTlUFy93rAMjMPf/5iUcMWiZJHFFs6CXW4YmHHVnBg/IMTDqL
VKve5uUhb4M8Pqd7Cy3i640SE3M/T0o7gwRaQRA+G+o5DrBzg/RIYTVuo+rWsHgx
yMON5z7BnRSMFWaxgL84JJGTc6cjcUzkHCk2/Nm1oHTLv7fE/S74WRJdenkMnAWf
tsyvtMDPDNCTzIDH7RtoYGWYkqX1cSkdZKUjgZWD0wXpU4i3OZX6V+FZT47f3ue3
q/7x4hWslsEy8BLlgsWk/ySFV/fVaKO/4Hnwd41+SVUfeX4yLt1gS2kjzTCRNl5h
`protect END_PROTECTED
