`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7Qu6Y90nrR0tGm95pmOFJCRSF9IJ34J/3kQQoTjPysSxI0eyv8y5DPTXS+LpX0fB
BBNeAC/pH2M86WfDqqVSD7UgKoJh6hSQCued7LXS90PPbPY5CArVYMD6HIq5ia/s
UG4lugXuUaFeUktiphC9Ur0NLzgeIrUYpVTQL8tu4l2adDpb1ee3hGsBEffNDRyx
+34NmMN7xGUp0TzfX86lDBvJmTZZ3XoTblyV+tMwlSgYAm119EgHXy0LXuwLSSLh
3CNVM5M7eWAeaF4Qd0AQjFgFuELceyGzGqOpQGeSrsfLPy7aZwAqVjqSX5nk5Cte
oTRehDQGo88FrlEvQ7CfRMxv5rRxJsmuY/yNvWjXeSSdV+dcOnjOvKZVyauGUUHT
FwHKINipcamQQqRH87OJg8dTI7Ybv7H1QLdaqwWe6UX1mMwBkWYBbawNfJH10vdG
VNHfaDsxZcUObrsWW1pvati4zZAR87YJBoXB93ZzQJHW7qoygiGsxsKnNyFM+lVY
/Fvny4oGg10EcXNURusLBhQWBmlnFCf5JgAj11lvwWN+c6lurLlqI/WZJOoC3ahI
kaP6/MN8VBO6/cpBEaxlmG8q6bkmSM9m5zaKsn8reFAJ7jninaRVey+J7SM2kt1F
bd5Eu13LRl/ITqK9yVpthAHfxe1j9Hb1aUZD2lOlcFL6VQn9arZWU+zN6eQ5r8n6
SD2PeNdJlFtjhQ8IN8Rd6YAw5xWCwz9AZhhTjp0WKWSjSns6+hcuZtgrpf8cbGOH
A/opW9EylxAGEcTCS5ljJVQnGj6xqe8exkw0GL33Cc4ZNkhxnCoVvU3HcH7nGi2k
Msdvwz2FO5jtjReUXROZQ4iY4V38fP+i759NTKeR6A1PU5Ib0bsK4GXZsWXtpugw
IEjZl8Ky+UEW44LgOgY3ktKxTAfsLUEIC/ef8q/u5A+zxHwK6uAxFQJ4POWQGnuq
QZUYeQQaqivMvHSyRr/DWIGdfam+jtyA90e1F3xktDH5xZagUNqRlj7FpSrDNqdI
HnBSIPA2nH/DM6RtmNHnrMFMusZ+Fh6gUav4x8PXuOcVU4UFcNpn7zskFBJIQwIZ
AjQ8aGYWqpuri407+sDf1kMhiyXcETaRvaYfFk5gixVRRVwWhcptvyihLp6H/oLp
k0qM4dv12vBl2Ooz5hu/QZak8gLcf1ssFALg1Xkyn3VWbDEPyUgDm7CQUcvlcgYm
tzYaEQrtpvpWDJFOzlstT5/giF2JvoRSknWgeBnAP8+22ycVC3bTkOsds9rrCfm6
1TWEpZi+gTNAcO3XdTYHuki9plYDCJ6o6Ees3sF/RGd97REN3fXSoWq8bWjBtxqa
UJ2JUUlmG6FNi2uODVTUqAbMGyGa6NS8Fs4k1cExTJlHc2bSqYtXeDAttODtrPd0
JafkkZsMORDZa+lVNplRnylwA5/RN2b3QYB4qLFbD3J5geJsxq9ZWmgnSsA2GKDQ
3fALYMQgW+VJ5iQ/4ifBRE11OU24dib+47SHbZ9O8IjVHW8WfIyfQcCTUnO/rkxK
BBrnkIus6OcHu/ZOZVVReqwbA5p7b0Hr2vcDOYT88LTKoYg4QUw7aiJWg/EBk5Y3
WRTfvnJXJCwLmwx1Mtmblu8OLaJTEeVJeehd5rw3mXhn9acwEJV1+34H6KRjTP4N
uqSmQ2aWmWtaiO2v0Ju5v865RJ/bMKQU4AJHlq3pfxPEW1ZIvFxI1I6lJopcXfY9
x7s5K7FI4jVIpywYE7McwCB8JBV0oQS3FaW0YB6k91JkpE7ZD/Cc/eukSuuMzAor
8iyOe9jC2lety0O10DPrskaJ/H1DslSr6jHP+0p9MmK3icYRdZNP5qW11x2vXkAW
xOx5jLV8awE8U5u8CA9tQSq5U3RlcrtvobMMUm2anfvimYT5xF742JZYneTZGkqS
fJ8eYWHCg1W6L4tPt54CW65uzMt/yyrnJYcgSPwsPZcsK2TLOsUkFt+qHOUAj1W2
dJmPWyxL8satFM57ninW6YBO7GLmeRfizZlv6EBo83pNMtCyuyINBpiK0f0FJZYX
SdSmJTOmSVVe8L2lwCfAaaGtMT/FMsQSFeLkZZ0GINlSB8+Hi5i9OxkUGn+awbww
KYXrnkcjqzsppxnIaomESJasI1gBo5DdFfXksbk6+TSjN82RjAd55C7id/4U4uHo
SDdgoNaRr1j1FSSOb1dnWqBJGRf9hrwyxgUWSB5Fm6XQRPcB59wFXWJusEa1HUve
Q/EmiCWmSIMxm+s2DVoKIrz+oTpXciOoShLBfE1L9j2l0yGlyYiitBXhuhKs8b7v
qtzcSp2E+CCiWQr2TBPuDVR4FUhZhcncbDMTjQNpvVk8pXjWZWvUKycJoAUZVOFF
Ud7ZNiwHF0MZolZzu9J5LbTvTm2PzmU6hW5V85ftI2JY4C200FgwgCe+fZ7VqQww
i+nkxjTSO3GJ7iczlLADKsGtBrNsinmEpkxHQQHRMsLDRFOqh/cFDPapVdml9ui5
bYgi4Qx84FAxjMvPM3syiskm17/ssXo/c/yuYPR4aDFA9skEtqfK5EKRGFERAY+m
oj+e4FzM+1tkcZIADi4a1xfhnSZzPny9ZxMKwFUYUjraqrvXNGUYvRpIylEEoyP1
UITk4Cdcmqj3SnlSUVuudShA90Kp3g4276dTl53bTQl2+Uxp6ocQYxbtJ+dLbjCq
e/+bPNIdRHOKtCGM1fnABktWOVvlEkbaDqcqUibBo2NVaHgigCq9R2CVZhRmivp+
WpJ2W4n2raOuH2dopPsEiKvgguxRhmPqWT8sw7PWerld/rdfqyjjFNjM9mfXQapf
uUaQ0VYlmFYpG2CmBhvA1iWo7E1kk9QE4gE7ILyYgZXpV7s6sAZn5HXwHUlRdBSx
S35hUSgWhxr+kqwTV7IxMQHl0x+j7IZUD1TTVaB5532Cx7Rto8ZNvVYcaGEx31+8
EPbbxRQgOYLoyhTvZs9ihA9Bl86XLhT9EAIQKTrjpyXdSxSgWr3cHY94jWc9Acbb
4ya5WrLJ6LLtIJqKIwTc88yxLNc3VUl7aYmH7mDj4k+Ml3guu9JLpyxRJlj84xB0
vmuMc3QlXqEA/kRnyKSpVqPK9Bhtx8l6RMrtE37O9UWG5xzf3oiDmHqKZvazE2A2
M3salYI/dQwgca2HTo6DbJ60rradvDUcBSV6IZOhrPKVgDDciS+9FXrLZLRvILwb
KLn6nUK/AnyJhOkLERctTldXOwycXe/uQW8mjuNJhJupsVTR+UA7Ep2ymJNnHpAr
Q10gHZBTlYQ97nULvfMtI4AJZ5RHQZur1owg1TM7dIR5DrhOSe7QsNp5V3QFxwGK
GJ3Ac1Jq28XNkWm1yTTWqvJrqRDxWXHcG0n7urVkGGozoigUmvX5pr4W1edu1Zfr
Y7/cdVbxtHK6mm6YQdqhiCm1fRAOGGTI6d0mO0B5cFiAkLrkNspLk1y+Tt71QuFr
SSwpuiZNvymLul2tlTu1NbUJsRsFXLiMUcNBOhluIGJBKLVaQDzuz4tbqIlH6cFs
ipC7ZVVL3NjRJN88xje9uotzzlH55oSKjaywLvvc7Lf5voUJ0WtS9bdYKkuTM+sF
zxNk7/3nbcDS47NRRfvPbKPTySFsgv8GnKj3GjeeZcxmsH7toIate7RIGcxuiRct
EQFE6JA05dTIfNgIBQ4Qmuw68jCRvVhQE5h+2eN+MUxfjENUTgChPHQYPr7NvRw/
f0x34gtnrN4eySljJUD/nc/6MmZvzmumCUffVaRBZGpFpvrJ0nIwUO8xc5K6Cnj4
Y7FBhRKfoqXBUTTRVNc5LBo0uxomXk+3Q96tByxKkAkZ9Dh3XAwiVbDKeRzfe5ms
hkAneNvF5Gr/LLXM0MzF5d40jOFGgrsw/tXo6uVPRgq/ns0qWcDYvMyJ/eQ9NlyJ
CwcPtw5trRmDwpW1HdV+iviNXn8NmplY4Yjs+jU3qSjxJrdAoMY/fTjTluLb2kxy
Um6vdXrip2cZSKe6s5dz2T9WEObyIEBv8VhHAcX8dpU9TY+wczlTEMmNiZ1WFZb7
dtZstRROYpR+O9tNQySy1swz9hWQ1HlBtvPb1wCU0iKRcl6NawoQSAop7qTiLuuV
kczgHAzcvxAbCFI/5JkSXzmGrP5zF/iUBj5ForcboWl7KLkyNar/pg1H9+RYzWWk
jWkFYuKh+egxinCG6Iu5bXhVhewJynJ6ugiG9jRvCBJHvliFo+seNhSyhs9DK2OI
TIhLWAzz2FGQ2wmQLMtUhm8Q7i1wGZ9OfdshFIj0zgUAe4N/b1oJujCxzEaRyBVj
n4zS9IbrPKT247yUC/HUJAoPLFR9yn/oj+rXeV4UzJdiD1G0T4uNX+8YOclorp1M
kPhSONaSIE1VEbCQC62HdjTgxVFG+3Aq/pvoj7go7yNm2CAFBnByY4V6Hurbad03
6qQB5BSYbqcd2GtLp42dkna2OjtFPl0i8PECmGX+/sGu0glxKFRlDVG/eshjrTNK
9mbKUNUQd+CAunnVtyaSJZkThkowgP6D17Dg0B9VIOfvJ4PcoyMFeUYKB45jOA8P
EIN4XdEK68xeMOFdecc/mk1csBMdO82DV9R+rzbo+Xhc/fRMF3UAQtMrH7glxDmk
DqmVgvTU2qsgW5u73O14Hf6A4pyuJxBDBrBikfucri8IpSm1SxJERppALy3tJ0Sh
EsMiIZXgv/zcpS3Tfo3MVMyqQmO8LwaAox87QkrEjCcPKjyG007R+tLzVbemj6GW
+4fbbsbT4/IFrHHVcML5IsWPg4WuoGzrAUavQcl2xqo2wpNkY6DKO5y9CupG51PT
Mac4I0a3XDaIHCNIZx/d+aS3zCeGqpbRZzwIsWAB9LPS7JP4KuF3m+lo4IkG7sj7
3hog/hFk5IzXRJDht7qxcOKcBgXg7vkkf8+Sn68svf5ngnOzruU8g9KN6ktkovn8
DySebjzigYyGPOTxNfezR0Ev6FxCgQKML2+Okp14DHLos0fmj20DjwC33xwpVmE9
7git+XMEVUiqPgwsNMEwunXDXGAcEPRdIQaFtfYT4htJ4OFGE16kgwfJjcJaYqhW
7sVr+IqheILALPwbCbGSL3hijVbwFb1LpRAWWVvygcbmhCLsDzCtUE3n7PE9C41C
S0lOnXo5HfxeuNRTT27WUI1X+QzQX/SDrfoqk9xF30eyiQQ///06pe9otmjBi9je
HlnLPECYj3Fr86Aqk+tre3j6Hmz1u7/pykaBHFX/iYIDr9e87u5CAxboqZbagyA5
9u5M7DOWJ8lJGm6Ksa8LplvifU0JxcSM64IrkauQD5sXOCGOJzjH+dQpEH5zY46S
o14H87ZTKHdSgpIbqPSwjGgIjUMYXlowFEN4ynA+L28yEGtsjyL3gwx1Hf0wrgw8
S6eORy3EpAkzg6adXh/DX3QElKbDce6vHC2pXsxbT1hiVPivSnHgqwxPh0hJJzkE
XCjVSRgBzAwuJzB6mPP/SEGShs1xljNNnWxYhxsUHHW4yNPgTfKL0CLWbY8WAVEy
4PP3g39vVYDsUdHCjqfc9nAEB9L+IGf34Kc3OzvEmqFpidhRb9DiWoPOR9I1cCAI
Cr8ZqNzKjlVvKcH0n/syy6hgbYCz7CUlX5aQyunMaQsf1fsxKjzo0shDa5yKIBm9
2+AS46bnSrxdxRXPQblpmXLdv6XC7OwzSCjpavndnRmbSjbXylNI8JAgMlr9K+eX
iG9Ve//SXwl0zQjHnQHplJbHg4usE+rNNztOsTVc2Kcu5xo7crnBsCDuVK4tyn7A
y0pOm7mCF4Q/jF8bYnpAIIWGacF/l/3k9txv6OMe76Xb/sKF8KaagSreqgZcEvK/
7tTiOK5Crqu/VaW1F2OSls+SEryDzUbbJg8+QEhNVKdAwlBq7NCHfp6hDtD9qqVJ
nFiYrxYG00cInxL+v9dnC2SszZfS24OEIi12IHKvdZ5XQrnH6Zr8mGjQ4MZ/K+vm
tG2xe/U5qi4j6dAMK3gTN/yJ/N2lA2Tf+yH1HXqLt0D+yKYmJPlWn8q/FjXYXIcB
zrb+ON8VgmEpWLGVSFrRf+mAVb0SehJ6SOIggYlIwbrdUbB7jlfdSF34HW2ijnSX
EKyBTJkRmDID30kvUwm7sMg6EbvVf28KOAmi5nFT4TyLpCcUksWTAdB0h/YZDACS
PGFuqGYDNj1xrBBl+8+0eW9exHuSjgbPrSQiIHrRNBCkDcfaPvER7GY4V3sFyNWe
gdOTtxIfVT+sjY9Yo+Rm0QgSgGj5+MkBNOv2DnjOb1gUBjyDcvEd2D0khQD8ikcg
ZITwv8VoC/GZ6LJnrFloPwdBJqrlQpHXwDpGr7f8UW1kFqvzll9LNmoT58DadTgo
zx9kSEemcbOmIWa48fOARLRT6zTX0/9Sn2n3uXQed3iAtkaTorXmDvy3DHm9ZSH5
nJHUwuZgI5v/xNCXPQMwH25pFvSpDy5Yq/N38gzsBIL5syWMvitTttHXMToVarye
OfizKCBpJYFVzdfop1MSnWG2KJaCgwB7DG3BLbqUTrrbYlmgeO9xx0fFlqI/qNAk
OZBD7l5lCDjPWStfmaLLFHtSheNYWuw85cSETvCR91LT28UUS9+CasCKD0G1u39f
R6sWs5u/tbBjRwj/a0uDL6X1raZcKo7CnmiTGe/+y/Up0Kr7rPV10mRS0o9DsKFj
lJw2+y7Ul+vQSrEP+GSR1IsUUtj5knrdluQQhUdlFrt0b2leAg5hfLmI9luVS5WP
oSYr/9PpeU8EENUkV4KA0EHmgOyyk4nuIjugB7JUe4MpyqAZ7JkCD+B9vRJhzxso
fng5iogSReN9KWBPySoii98PLEmgWW4me691JgnB5UxeFIacJsNgkv6S4hUvE2xg
g2B5N5t1d3agLmEQIiFZBUjWxiMBYz/m+SpwfcnDM+OyzPXPW0XIeiWrAFSjDupW
ku7XgtzcHCIFYlg3afoQlzCs8BN4WNzqVOaCztmdqnRFBTWtiLVZu/exmjdMrIzp
rKomzp67rO8N7qx1g4zC3Fon4TWH2WUqiVI3sM04fBArrtx+tNvQVMqGn136eR3H
ALus8IbvBpAxJD1SIcUD0M561t45Aj0QrkFt03r/DlxGLJXVKxFUQCL5bmjQFLws
7jMf2FB8DzfA2o74Fb0bB8SBCdrVySeqcCVVlyM1H4OZ6LeBWe3/Ex8aHz5nw8xl
rsKe09zJPtSynz4gEnsH+nRhd26wMpZa5hMthTQW79ujRHDFyVsWB8BqosZj5ZNS
4Iz7yZKiYpyPQDNypNLbQTugt9S76WFQEc0Ju3YuGXGgL2deKWLZiumG1fAshHXY
iKEKJU2Zqp/TDdGEvapWXMdLC2Vb22ujq8klBtVWU0uGp/B5LA9mqQFZOvsK0IUk
p1bqKJQo7VHS5KkWJnwPzXcKLAbW4bIBU2H4NXB6nJsev4TljUvyfe+cbLSxtkGb
jRYu9zsKhtm9HL83NBxqS3JQc+u8I5X0vNlcLGWDROav897M5UmZRSmd1v4DMq2n
K1wFg8IjXquI8XTqnCdPqSBbV7L+vLIm2XSb/4Mq5fodwFJoqKEAd3QSdvZ8LWS4
lW6Kl7uetbREA5JQ5KTMlREZtLI6zBrByOfu6mTuxZ/+WXFIDzkZAC27mIUzh20I
w+LugJk7ML6idJqpTr54bu3fPlS0mhDmey1iwrM/LUWbtywyUHcLDgw6CouErN65
B2+3+q8Z1W9V3aPtDW0T+fwFjOvd1VbLduPPPz9ADIl6M6GSv5BSRUiybif32ymQ
DjiBr0XJn5y9AIPl+Xk/ge+S8aqYCSkrXgVMGYcOZ9XI3abVfwpeD/wCwCHszaCT
CKqLiRT35n6LgJXQSbq5I9ZtQi0+iabNUhS77rZI+Q3NG5dS5fNjC5R8gOEPAJF+
7KCNdBoOGtR4LBf44V5JMUaue9a71yOwNfbabtQMriqDcED2sn+4y384WpxhxKMV
ZVguze6rK1MCzUS0HOgdHCeUw4wXQFUOH9ghQATLZFzdGSkheYPyTljuWPthzEoo
CINC72ns6+sr03+hnlWya862Bnbih5WsMCeE7EcnnIsHv8F8zBvHcj8kyDELI1x2
THdYarqaSdCcsKzoOqK8Omb9tbh2HV3TqWGYxSxMpruJW2qIBT/iAwKex0TorSAx
c4sqQ+Rl0zKQI1yPqDsa1hg8rFKklrQUKFLLawyUewOBvnekUdzchp+2n1i7/57k
0iBQuihJ9o9zlNPjg2AsrKYon/yxaoDBdj8N6a6KTgS5PWXPHNHdoBUuBfnVwTf6
FqRNOwPjZp2bl9blLDiNcacdNurBomUTDaUtAquEAD8oOIUAMXMfQmZ1IihD5W5B
HCC7pu3RDTRY/FrxV3JdqXQ3TQrzuyc9wWtGf7RyHpRA2X3n/+CKGy3eZIgB2SGR
Cgd/5YnDpUCx61mUSzmNhouoPRwv5pxOQK3kaoI/mv4POQ1bB+PAXu8FDsvyr+5m
XdCAQsC6Ch3Dh76C1dvwYYuBk9Mb8QsNP5/MubqVEDHzOK8kazvQ75htCOj4aq2S
TGHJVIffR8CnpBfsCE3nkNEEb/F7QIDaHz8NgekvcPkvg2tJvX1wzMEHeZOOk8p/
duTykGa3aeNSMbA2xUbPFmzOnS/VpGymW7pMppXQVFD9C69Hnhu1/IpZUfZWUngX
yBluNfO3dGqovy9G93BzaWOI2OqbSO73JjjLfcS3ohQNIjDz3nLvnzLYK/ows42T
SRMh2Cz9HGlejBQFCa7dj3PeBl2rpJTgWKsW5miMJwTG9xy2b2R4n3qinfsXMms+
WQsgdbeof9xcHVTP90JYHtxnrOdOJDMX9BOSndyklwk6XpxaGqLkybgFtJtLRbSd
NG4MglrzKKcCVT+8a/BJZZZxh/Z1x/MngiRrcJpNxcUTSvwrAOgfFo0uwLvaq30z
XE0Y1i+v4L1SOQmseP1bmM23EujRYdgUx9EQymvkAiNP7p2ar832EOnoqMNG3++s
jwZD67SJQ6XBBGQaBiblViTjoOCaUGLaiqG1K5MZJo17At0qRtFwF5+DNQYXRYxy
VcwU2KdETwuJqluqIUcc94hrYyTbDRbeyR8P1/mxzWXDSLR7TS9OMAuuwMIDeH3m
c9QMlFZGrVmn//tu5S3voV++y3dh3Me8FhJLiBKRScc426TiJTnp07+lXbDrQhiQ
EqbH5oF8B7246QCHciuGJzEVXnx4l2Ee7yFy8FJyC3naIOEXWaDTQteeO+IeSYzn
PdZxQuy3sVO+icZqkxP6SF0cj/56LS8akCJBYEtH/aDlTGtBdIvBE3Iot9Lk5/wA
w2+Eqy2bhkUZA6GybPB9/mYhr3b4uGWdGLq8CooEljpbOUfZ0vakuyespphafN4p
occSTW7PaW35CniUmm2fZfTAz6XGVAkyQWFl+2YGrEwW9FZunOcYafB7M7KoPCWY
h4j2yffTIeK1i90XklJ8VvzHMlkdxioVIiqRgbg0+yEzzRpT6x8GH4EaOXXmvCLl
843AzLSodhqwQhTIri3of1mTOSg8GN7sdlSAYjebLZ/fZtDKLqHlEBOTnWGSQjZI
WF2P/XA1aqL8a26n74eV3KOAHNpF0gVRH4XeiEqICFR4xxqgsgvccw2GGSjTKBV9
hvWXcR+MDOMnl3g95epXpG0IpI/7SdWCofwr0C1eMLUoUuSpaXqfoYPcYypznZ0X
uUX6RW+80vlZrJ/9zjtBEnRuL/Iqh2QBkI7KEDPcXRkkV/fxO+So2SWuJrqTNOmh
fSAJD7SJJs9IKeYf0RdwqU4lR1uJRmIxFac6Wqwkvky7z8uh7/7M+n5/WwyhPuTo
67YGpFz4s+Mpr8O6mZbcK9waRHSP9gkYMoonkQn7VzA0BX/6wP3d9sIPHjtdSYZf
NpO+K1vKe9+PwSSKPBdaJZrs1YP4ARyXtcu9GGSLGWXcp9fxVtJWUwOOYuyWo0jz
dYdpkOz9YmHU8cVJK5jSIh9pl9nuMworQaKT7vxbvZAU84C06O5S2hJ1YtD5nmhh
XLbKgAbnApCGn4N/9qDkSybYDMmHP6BCC1XG2ynNSLeVROOj3joVKNdjyoQ3+T7D
bS8r779rHUeBj/bMuBG1Y2kEAOOyCddjGdRV02RQEsX8hByo8MYiDlKl8klhx7wz
8LcBipOxTVLFlWFhibwQxecfq3TNhVT4xy3+8lHpJ7Yhise+9zO/7V1WfDkxatHU
hc2gPCNkRLtv0EOWRj+Snc5cMYUXpdTUQuy7Ee7LImelp1mhc3Rh1J+MwhUkYhOe
eDn+vtUdku2I0w1zbOqQrXx1hM3rEgykUHK+YBwmpOaNFMNzp9qrUkTef8S/TK9B
aF+epfe1wV6xz2K7X9ZieRZHERtMAYkdxy4ys+L4Ajd1iMDkfsrSprJhb1opp7QI
nmGqLqdjsGLRaZit3keorLclI7L8vOswUiJsGc+XwR4dvKMt2XdQV6ga3rS1TbrR
0C22ISmAhE2qdArK2tTwnkR4CfAuRTvGNUFmyjhjlE5fBvSXikpnodNtKQSQIefd
yDJjo9kFSP8PS6qxRppBG1c9URCmTNS4vqz8ZSmFtSO6dwfhHZ+ZaUZTxI6YIFJr
NPAFiaRQPNQCAqMc4mMQflVF0IghmXbFzpHlFnWU7/vfyN22ooVnkTL/p1dMb5VN
dGPZ/X7LjafzMkkBbge6mILUrv+OaNIrC8b9BdF89Zc751s3LGECXEgXeYIzyta+
8CkBj6eO3fZ1uHKT3mliBwdT2Np0jyBTMGaqrNLI5VPQsO8lVLneGjpTudgEd1hp
VAnAB3e12qaJp1zCJN5SuPwVQntQbO05Z8pZw/d/dr+kSTk/xutnLVmGP1mbANg+
phR5IlddzJikqyEZK/38/xFBYt9G3QPVeeOPuoCm3/j6rFLMHQpJ+0qc5M8SsunN
6XB5YWTuwt0WijAYOJ3hUhqPngGbqPWSljsX2vckG7WXg+4ZXu1Yzd6mAP51TlfE
OOUdJgVJ0UYhbRZok+0b5Q5mh0wcc4njnuyjp5JY08VkTYSCd0hlvWSioQYi8jiT
X4zc/2SDMHXGj1Oxf1eYgiVRSTI1f3iiiYMZfyZ5QvfsZdo1r2Ab6wgO/1n8DHqq
No/Z7ykVDsB+2uOxc4/R7Z1d0M1FQN1xLxCOA/RHZfrpguy4gmFcULZfzuPOUJEi
+5ikgjd93SDilZb6A4aPhyooGtSxC1b+g/sYUYxc0QgYMV8TgdPAE44OaoeEq5ai
HTBAEbAHIozfe6YJba4qPQhcFd5hiFcgJJKH2ZO7Bi3Q5WpKWbNdbV+jv3DwR6b2
Ivei/eNn96CQGyaDi7IWY8dNvz9ueUW39NWPgSd4v7NJRKKPetMyBWnbgvcQabL0
pLv4HOQkribXZnNK4pCxWWqx7vEGphPGFzYA/SL88GKQCCqFHMjR8grLRNBFXCHO
z1OwcSjUrnqsVYStJTlaVa7UePeWgQo6fS72T6MC8c07Wys0wldpvTu2YrQSWjda
AlCs7eSU9LTpxXnHNJeG5EEZrh3aGBY0bYWOkqg7H59HVxtwtfupEH/HJNBHObMQ
atCOvPEeoNaTrpaHLXTJZF+ojQhnbfWhLxCACEcS+UvcGQtctFGXRqAIYah3HCyD
FvRwfaVPFhLXkEy+hUkjyLpAjDobCxVAgyZY8FNdyc3nvRZBoEUwRqFa8gRjbsN5
cjdacw8Jg3gCpBVHfsLAhaCWVErMvdeqmX8vhqChvgjnX9fmhlqgWS+3E9PUvQmj
RqUfCTJNx7EcV5gofkh2rGImFT7RQ19pRvsvGnwntJ8wybmgcq1BU9VbrbOOPShD
myftzLyVAAQcU9JQMoLkD2YvNlk7pXl5qSSCT2+pAyAhbRvMjMQeg4eMkCxDTg/E
37e0//JZ7p7OLdUM2ThU0R+7hLYZuIMkP92kZHVJdP+iwaE9Oi2M7qVIsA6SrdGg
A6Ujan4uKyHJUQyr0PDCjM7Hu8SvG5Vze6Kbi2D6A/YD/2l0uevYidIZmEBVuyIs
ixroNu7TTEiflnMwKJxWCXLOcrYnK4ipbYVy7cZCezdn1TLWiSONcE6ZHWZV2pME
YR92X04GvMRuI4PM9sOwWt3dNTjLkfQqFcqhoswf0tsNtBfH0tp7H+svc0ODdQzt
zqmvWx/OUHXOKv7uxoM66sKttVPpsXO69HJdpEyzUrZzPmzixdDPy2Pq+PwtiHA7
As//gFQYOf9lvwg7JMzo2TuQjJAZ+0lBkRZgA7OIY/RlmvtXNlbwL/uLTizrRq55
65J6zqWkkCD1YYjoIbCyIrkFvZLUyBagK+uc04iPau12wd3oAwKIC/A5I6X937+T
x2NTzre3nB56ZK6E1TE39UgKVTmjdzOBbHIAkyJTT2dWK40veF1PI68/xzKYY72A
fGgvEMwkAOPnjCTdBmwwmvnClpbQVRFNZtkchlV5zYIdqnPC0q0cFC6pF+D1z0yc
cVcRyfKLUuzyXZxodEKpsN/bbEX+ZYg6Y56sl+DfONvMDR55qswbrUebghtbVEZP
ApEDzZsf9HeYFUjGPI6N4mQPRHLfkb3ZgcIepdIEm+kRtpMgy+rpaYC9ixGkjjFX
eI34V76ckSokGdTRo9lECnyi991B6uvG9SCN5wK/qiZMAqLUIIjkTUAzlJcAGWL2
0Ui7Et9Ohnc7tKEqmQr4tKQSeYkOdFh7+QaNqgNHshk/1jdDeg4bbzlxof+cMFdL
P9wVxmbovb5sizE5InOSXpRDhFr02vy8AhFMzbrvTYZvGOsNuj9A/lXXrE5aLfnR
Z+rCqGz0TXDlP4paIlgGql/tx4QsPHTWQpdFHezFCdmsa9WKNB12j+mzYvKFAwYe
O60aHLPkT0c9sgw4R6QfxCNcNm/5rRTuvZcbDGo4PZYM6N8ScRMj+7epyu6SLtLw
qisqEIlaJvmT/chfDs/GrnDK2AEnYwttsUb5/+PPfh6/hcN5Jm5EYslklVvUgLSu
wWrYkpLisqNwzRZnGcjfHaO4gc5fyxHo/XLofX7+AIsSNVGA8YDBOPUNePL2IgHy
Bu3xCg5DsbQnu0Qkc+io4DhUYL/t09Mn9h6yER12VkzpXXp5TytDYXYNTi+P4CnF
Y5d41mz8K21pf4NIrJNCzVlNoms3TLdHxWMqECOEIZkzb6sEENAULWcL1Cx5s4cJ
ORC6+wropEBtYaUE/txMmpeUAilVQm0D0E4SUHrIuFq7fi17p8NrcTKFYEH6tYgp
2lBLcuv8pIO0tKvMW2sHyVa0qtkuBXbWVweTQfsNPe+x8HXfU8Lop1Z8nrOZHzaY
kuHvOIowHzDNCaIE0neKXoU8fbhPbCNqoHSP32wnDM/hdNf7ZhjmKsPAKksJkK+E
iwvFH9hL8LMWhrCO6DZHELjtYaxLVzXslNWADHlwEr8DsSUo7lP7eIxvieaExgqb
W9KlplhbEhNPhsZ5qUdLKI4HADZQDusPVD3g6iBNgPUGFUeV+a7wKONTtojrQ98M
2Uh6RIuqamppZ6LT8uc9QD+r4Lnl7N8zNQuIz4NK+licGAQnrubtO5OxdY0GAqv9
f1JMgQ15tm2/mWtTGsTsjrIBtlBzcAYnEINKw0HDIhNJEv8+LstjwlL071zHm99g
GLQzEIlzAS3CYxu4qncl8YYR77eTkOp1oTiOPLLlf2L1+DC/gFSKIvijBOrQnJjV
TdIuVY91ZgZ7FA6NAJn9axihk4tt7jYtVFKJylVdmALq5TUDhHjqhI+rwz7DXpWl
zT/8YBpyTM2DnZMObxoFsXOBOt71PWznIcjD52emZ0pGj6gabRJOvGBRmM4LQJ9A
aj9rnHoeRLuGjHA3Sqlp3+pgU2Kf2r+/IA4JGiTHKhTpQBFSadw3EWQ7Btm+AP4x
znDcKNwbBLCKg4Qb6tpSbKPiUXdQekVBLOw2n958YJianJu+tRc1sWKqyxnwHbiA
6X2hC5X6aIBiM+RyTQV12wt4HzZS8/eVhLTvb9+ineyPzjSGrD4RPB7cv8hII8U7
WiNrsoo73sPrYbRBVNLwl7Ad1mYEVgORgvc6fyDhzoa3yYDrcLR6soTPkuqXi1tj
5yPW4vxCoanDZMegZzCgXX1unCDHfjPNq7i0XhR1uiZeRg0Fg6mLWCfIVVjJrb0o
VBb7tXSZ0SS1MR7EZrhcWqAdJ/wam2Mo+bAE2FZknq2VPCzJ4C2tFkkFKCKN7EQ+
qZ+cEAQ5tPhkIl90W8fOecwbjjqcnYNw3mPyX2hy4JhOedCWEciLJYrf2yyOqXhW
oZ4A7BJoKibfcRzTUqkdPjEfz7CB/VV4GfTg7BCNoX1d2tk2QJSa1fFIAllLM8KZ
Gr/q67bWgkvVZ4+0U0yjk3rMrx7GlksJA57SzQUGBrXGVogDt8wBj1v7tHdQ4Hy2
KmkST/Dm9M5XjmHEBJxJawtZ1JMXwipPmKRMKJHHLjefBvBZHhR6xmhkMvHg/Y+p
jC667hEshKuDlg+JsJtbFkk2s7h8wvsH9LApzNwDWqfu+JnJia+U+at6UQg/lDYX
dulEByCochJ86Tc1C2AOq8o8Myh03zqNHO4zdiuP/hbkgKHluT/mTQvVNdAVyMt+
LuNPnDPLvuZKqDiVXxV8jCrrSWXoBku7Yir76Gx2MWrr9BnC4WkC+6h9OEHWGQb0
7pYkU4TiLCI9b19bqjoDw3q3G71unmZP6W8LFaUUcAUSAR2IFVld7D/uXq/SkpHJ
93j4L1A/im9M0POxMBclqR3T4Z6uieeHMk2/vQyZpUDQADe6iBSpTuxyNzo+Noz6
BPoNbuk9gtc9RvNVUTtwI8VrtcOwyB4KQxMyrCfNfU8ll8ycMadrWr56g6S+c1yr
PgQmQSVhkBLnt2NeaZ9d5zZEb0Q4LFAVo/oH/jEcxOMoF3R6DOWnZo9wmYjUB4Yc
2uELX18/rtKxiDJrim4VsEWF+NVnCQphxwHyjS2UVZNV0BueuJ6uoZqZfgILOFcV
0tmulVbSv7lOeK8tcav6WUCPFurpmH6Nh6DkpOTFT3GKmmtWK8LbCvppH+3RcLxp
p92J+pLRXz0ZiF6EaO8btNpnngJA4taU7E/Nr2cxJtB43xHVrGBFB5y722cU1uap
azTI4mIQa2jxBYjXhNC/RXpARIdNMjxowdyBJfSxEJPMXH3vHkaZ7aQQFw8jcVQJ
8878LWBRzr9Tlnyh+UhUfHXsenDZ6T6ESgqtD21hI1xo+91HyxWPI6THX2P0/NhJ
/rflEpMIh2wT4WsIEUrqM1mU5aWKnL+WcdrM34oPUPhKMBqjCdjXs7htGu+aBTaC
jGIkNuNWSJTguCrl/yVdVxdCI27upnWJ8dLCPY8tqf0xnGv4UyJ6YWTTg+eus+ps
jVVqXGfm/BBTWPriEqV1brZX3T0Iicy8FOsSjqpOcSzu92Pc9nS9qGRHNYfrR7Lr
Nvlt6BFCKgkYMEVJMvsydJe5VzVxbZAwcTfR87kd+u0gGQH1cMDW04KqxR1ksVOk
k9Acl9y20nrV1jTduns4SfSK/UMcSx5DL5DHKitk4PUQiWcJFl3NoxmeeVTWf/xA
kXWR53+ffstRvIEVrFJDH7Pe9Ztia/EehDNgfZEkbMm0hPO4vH0ngGrYoof0Tb/c
oNr9qyIZjyKGePlNEwptbtpff/yiFoEp/WcgbrpgH0Zk4pKxyKllHLOCRQRFwThO
hs1lJe30zg9BsxsCPS09Yl30VVt8MdR/J7U17kckBvP244+pvivfogBX59xpvTpN
hYH31DOe41IIM+oCqr8r7KmtbewC2wC2PT1JNPn0IBeBd/nMLrImrQJYaQQxu98S
TpSdAvslMvI/zwPVY0bdYq0fdMiOFWga6xjO5Olhu9JrtlL6Dev5diAt/lBwiM3d
L7IJdmQvCOh5P+ZuZg5jkWEKcDy2qPyS454sMpuofmEFJoKlb09FCxWeFIsB1iPj
kaVquULytlPyTLwPBsSXxS1XMMOsoqbueEr4MIvqWrLKQj7NxTVfZaG/4AaxDbo5
r6d3tMVKQr6Sld49v7xg2vXLpAP4tH6JJrwh5WBRSzspFON0djUWEhuwqPQ8G3BT
gTB8VfAko67Zh+wPyhiVO8iCIGVuAzsDmptiVPZQ5KgZLhVdlmgrf0VgevVv1MiB
syBFw82fclWHY8TY9hG6ng4z5AIE6/K72kxDUdmuIwxjEHqImsXrjwW/ZqZZZwdq
0sokHHUoSPv1lFqJ/o/0bH8ZheLyKV7Sfw1hOgINRz/G2lXfCTHO9FsG6264+AJw
kI5LXqVNCGXJBeVo2SiZBpMDYiTVQ/+D2/uqEqQrgqRr6yUs6EKnVIt9m0oNh4Qu
Q2TW/KJUdUVuLRRwi+LkLN9J6sFfjKFPGWOhL7nBvA+Obthl6vd00Bx6RJy9UTlY
p9m77VikW16s3sgo0m7cjkgKecnOhggTqLsFRPGb5hujtAXunc6z/Ddk+jba8PUs
9dsOI8h6BHCaOKG/vbk1bmVZznJcMgsk6Yqqt27oGlykm5nqzWkkAEMlGL/xrMSt
HvQoTvPUAttdjs/ZThVJv6JT/PVnrBV0aYAJKy5tV/soZmscndLmWRiY1rp4tljs
EkpjhCREKuKza+5hlMoMv8HYOL3qlWI235W3x6SxCgnTG2yJhUx2Rj9cAQK9Mgo4
bgFuDTI/zG1ai0TTenDDXthBVM4dn70vm8ZsW9TUV1kfwxD/cqWg2xZ6krV8HXgZ
l5e18w1FJt+trcym2LL2mH3n5JuFh5wVqdn1RsG1JuaSOJNqsqa4pmF+EbNHwwVU
K+8ewKDqTsKNA0LCvKoDve3cZyByBs2IQYpmDtBdZvhpZajCxq0zbsebTyTDu/de
cHqRn1yPaSLKIn3h4w2SfLD9HPEHks0CLo9c9mthIkI6Gwcx7T9UKX6Td3J2xrtF
htgCH1YxEBtXmN+dc88QSUBaN/rFAeM61RjUj3ypqCXOEQQ94KiBWaLxEXiMnIWq
in1r8tnoGwvoUVsSAhuVLDx71G7BiQoxzqRx0m8f4dUxlnouESoT8cmVVSgj9et0
2p1gWIjSUZnl5ygvwEutNGmGFQC1Vh6UJHLi7/VTONl7sttUNIsq9G6V13MELZqt
UW6+AIMP4Tumom+kf7B6p/Q8LfvugDtx1H6ZfxAON3Um/hvhUdID2t4q0mpm10e+
UDZqaX/xBGA9SbWuzr2RzY0i8/H6PqoYdBLfgjiK23JBgsd3pkp3yTmTtCmvQecI
1i1cxgolIewRx7yhLxX7iulkmXAEPNvxrgjwY3dvQPul8ozLGgWtmW88F54xuqtl
0nX6G9Y6By/Fl+Mqq9DFp0PqjznHVmOALUBitROZ5vd/tpoRSl8bl8/NU1lrdbYQ
c4USANiPL5kcyITaNaf+AtQyDcRm2aW1Gn1xqD7WzjIimCCSdnAEyA4qYZh4OMd5
FWwPn9QOCzKxmHeGSelTlguy+x9/rkhXhhc6wewoVqddbx/qIP4V69WfKA1C7ezb
TvDKxpXsW3ziC7KA/ior5lh3f4GymEQBnHL0BRmNygAFS8xTB7huj+T866uZyXp9
hh52sPaucG9V8oE2Qme77hNWKWnMRKzFlPgkWgd3UtgBu6eJnv0XWLfTfdJOPjuO
6JXx6ZkRT80999cqCrj1THIFpiYGXeIes4hpRq5BQaZkzbsmZD686O9BQJ+BPKEY
sdu/1p5wPmI2I+dSHxbMF16yQYiNe/fiYvPlVAskUbCeQByd7/Givg+IBPQhEIyZ
Bl2jzzFpGp4w/Wd3LC73z5HjnrXUxRItepo5VnufssilQPqqUNug3FG/QA1XIGMi
OLMjG0OzW4Blpvllnd86J7txE6wsKIAdrpUqQv0/iNz/3r6NgFZxPwMrdr8glW5U
CHvBgkHg30wa5v558L0QyNzvyqrIX2NpeinpFY4mQfrtxCKWIRczoDyF7T4k+XSg
SQVDS+M8AV/NqIvN5lGyA9mTjTvl9me0O8FVynl+WWBr8cafRqkilK8/+n0zQpLP
/upoGo6QwljzNGXIWd1wGERxJZUki6tz6E9157nu4rVY5THVY0AbnPirzg1NkRBk
JrYqwBPNFIPd5HT1TUVX/9p+rr0JlsM02AK5nxUKxpCR2nRkV0bIsi2VhItFSF9G
fS+Er+6LJj2p8QRT44sBYaCZoDmO2Ph21HshzfNeDiSkTk74nw/icXEgBmM4DPBn
KtLCv0k3RWxzSIz9Yw5lgHH56mqz8rbT0XGBh4URzNsRyBgmacRig+dwq8F/8wGj
NbrFBMLQ1b7gsVbT7PlXk+kwPs28l/Z8iHOF5zc8awnN8JV+D7dLoazhLg4yNpOU
A+G199lcBIvMddaNld8DvUPd2NWiJR8kHWkeIKsNgJbSvJIA0Lh1ixI8V9sAIvn5
Iy48L5Yq0TOMFcpo4FzKnX5/M/7AdUbgZpdYceFu9vV00xOqFvaZrkNJu1RNpuhH
47ff55ZXpNnCGvlqHl9HULEJukmV3aBkXejm+599ojH6FKlSRGtazlIRbBKsA+ai
3JHJnqETXxOLfy9A1LeK5iwuNxv9MRvfwd+HRGO6D9SJFoHUd+Sb8uHYxV7THRRT
8k4RtrMMK/4/GUbD6y2+Uo4+aPP74sPO1rW2CV1XVVVy1m1dr68sLOmeEcLUwNQV
Sw2hre23zkhJI5343gJ8N3szMNlI0cnnMuw6niVzDEdlfeYq3xR0MbIKHP5DzIfo
9a8EiInvbx453GHDfJWn3Pz/OPi/S8539sjbUJPbs5J2YI7Fc4MmPraYbzidBliE
7sAizOZSw3UWGHgjKg7WVSdJeahP38rFI7mvAUwYWiuw5WXPtOJMywjW0+pSGdbv
QswRrbq4N+LFYF87PvId0GrZC3APKmeqajL1GHoeXiB1wWtWpqsFlqi+PX63oRyt
wrJXKEBh5pJPnotN/Yu3LbEulpiUrQqbAQaTv3sQombuftkRkms4cV0l5Qj9RHjG
X+zgtzPHgiIe+WpyX2t0QrPfFOgr01CSi8b41W7rUZRlCsPCAKY/VOdBU50kHo0Q
PJpEG4eU2ffdfKVdUs2amZC3VE4uR3aSMcXzMSO3clfsohDDmFCEIBXfsVWeleW0
cRTn9KYwzMdA+eNZFdqvstYEnZv0J36eB1obBE2DdCSxSf44igOQ0Zy9BAvxSInJ
AxBRXT9WLwAseEwwtSfgxgnsh6KhLAhmLaKmzu1jNEG8Gc63kdlJ+/O+P/pj9Uw0
oi9Vf0W+G7HGMw2uWLgq6VUwS0H5jp/5PqNdZMKIU6MR3ClrCF+/JOD20HMNa7/4
fEVq00J2vKzfTkDfxT/vld17A3HSklzZEOnhPlBaTEpIWVwrYVbGOXpY6qPstqI5
gf6xDYkZB3d7DMcGm54KayZ4jHbCc4uQX7TAAJ09iwbWE7j4eacMnI3fX8a6/oV3
gkMSfl6tVExfWKn4pgvB/OrHspvPo5Ik8tSCyUDTjcOrN2dnSiwtlvRBKfHkpA23
VrkXsRRx38vErj76STpQI4glhzKPBBXEON8t9UckHPj/aG1/ddcevYAqb7mBN13l
CzQ8s1lM0mL9dumNOMnPmz2wSqxe4ZF1Ffgf4T2XX0F6tQKBq3Q1p6ydgcs4hZ7B
F7N98skqAqWyXe3WXw3hXqf4ChO/3kLSfgrZyUgGgeTm/cSYW/+KKHW03q5fqGC4
3F6Abz/sxA3eJuPLKShHaXfSYHp0m2GxA5/zU1GKwj8ipqJv3AdxFbHRLaihubpS
XLuBUgqrOCvIDcpBbaC+CKBmTvSQGzUf+7fpKj7iSCsgRq39N5Qs5xTKyl3gVAQZ
UhXeKEzj0x/+CVWAs2Js+qfYQtL6jMBoK9+W1DdY05nmuKF777mWn4PghcHGC7e7
0zpztIjg47ECaH56K1OoXZPgqYBi6PyquddI3ddRoWLjbRnp9fIVLIAlsQaI3pZH
cybWjy/RZAqLYcmw/HNpj7OIfMCLtYR9PcU6gwZNRarIUnnleC+0C55cUgtds3M6
ktorKjFEpqJD/k6OOTMl8o83EzafjO3JJCOd83imnUWJfgRSjo9NXzMHH+UcPFNK
4aCA1vrjjZWmmV2jXZ9CwbnT7yql9TIhhbUNDPQbTwlKhVU7CSaDHPysGgZVfnAU
jqssAetS2/Rxjcd5CukF97EF4c2DUOe819JRHLht+WCuxcha2LMqG7EYEkAW4PfP
a7D5PXMuOsUPjdCxS+zjJXnJXwil7ShaZYO0MXbGqLUNCJEFtric2x9jtzo4ESUg
fj4uG+do3E/kT6Mwx8NMt4KWiFoEkullHBSOkRimlkHOUMsWnoRjcOTSRdbHirl+
rDszuGgjvaZ+5pToa77FtwrtKvlILfmNmgwJ0URJw5u6rj0RdxTEDYdDoF/Kd7Vo
+4wofGbX5MJ5tldimjEap893hAKQLy4I5RzBvYyuLjIEBHWOYOlLaFHCRHKVzn0L
RPk0AQXpDSV4Qw6Hm2AirmryhjehSYGuWD9hn0DCrxDhATi0VSxyrPfQfbV3gXad
/0w5rS73B8YfH3EkzTif2rTjPw1Y5OYTpmMIaD0SmRgnG2ATkRnmsmYmVLD3Vu5v
zPHAj77+XonhmZ7vDvD9fStU11kbPpfhtbzOU8IREzP25cVMj6ES771jvbeCSuZ2
bIwSz7646FmyC8xsIBLzji3XJ9g9nBlePbF2Vbo6glOXSsS7hM4cS3U74C3aApV0
7GN+0nC02MtFXD/wESBmf2hsuTEL19cFjqagcNrXGtHkSiO9i3TNnSLfk7Lm13Ab
o1yxw/qqLysWC1st920na+IpEpMR7+NefUoPHlEKf4o7k6DceUmDVjDKqr1i8XEH
RKR+J8kVtuEGpFP8Wn4SuzpXNRlmTpYyhvaGgyzUFtrZ+VpcDsmmqvY2t9CDZ9FD
sjtTLU8ts7bK5QKor2dE67SREHJQjwzxhZ6823PTomqU1taI9F3E6DMtIJDDEDt6
ri8KuwkzUeFBgdz0V2XWA/0JyA+YMcwI3Jiao5ivBYzlIbviGaRHjZAjMdvyeiin
Q635DAz61hr4NVzClUzQd3I48NCk/YcHoAq2vU91w+8KdWxuPmQVTQ/ByyRpC0Xv
EIemXdEkGqlk9iXQhgAzS+1WSMH0splu2gHIsHB2DWjI5gMkk27yjUMWQTjjQUpj
i9DoRJXYsEh6i/e/eqyZrbsDbxt7NEh+MnIx+maA/l1MUKC1kFEDBXEEGFocpwn6
bivTBTmhBWORzfYSIZ9hJaaPLgjpoblRqTVxJvfcraHAoP3cN734AhMFJNpHVNDL
D/H/imn+XzBR0q65O4fZ9LvbOU6k2KkWRYAdzRJ0dV8C6wwYvFXFd7AWr4czW7aL
tRvfVUPEaAC9BN9fx/jRall+VFYvomaT3qq4mv7IIaq8fDHQs84mu/CwWNzzCJqN
rHBz6+FsJTjuFVa1bZoMPkW7r8nyYaT0zz9QZlPI9wx2J2ulnq8bQ8aoQJtSd7ip
DNy0DJMoNZrgnnOZi2scA1mK0FbYjYZShDcjYB6Jnd99hvJ+XfU1ZtS56YSLp/Yk
LO/zpRDGKlRdZOSAmRGlLGxx6qdpNKoQ8AY37yXPDHP9R/ar7ZRJ4JtjNVyGVLm7
NJnSPQkIO1AGMoPqMasSIc1/Yb8CwDtGzuWXOWN3xbu2sfd+fhYONHklgSpFmKB7
sx+3HdsiQP7fbiOLODY3DPM8s2hSUe5IlNGCcO8Kf6lYmhTqJeFkRJcHAo+BY2nK
2TlNzCJ0RdMnmCCaP/TnY5TIQPWBpjVL+ikZ/ydGKlirn1b8lC0oB6FRmxIV4cck
jkQuURGVERfHz5U5feHWHq8jzHq8hK/lIey2XyaSfnyqTd1fdBAw9gFZRG7r1PkV
KXwz/D7gz/+uL3ygajpIIWns9ncSnn2WgzPCBLaLENhC+k86lxv4Sdbh/IWDNQHp
YNdtJi54NZkI0u9l6hrPZZFDTUIEyqTTwDO3coy/jjKtUHrTbxhZImCTpiGcO9y1
SKnIiPN3gy0YyxLeR/h8VGxcdUZdGlDzno9kdRaSn3NTXOP6q+B5c2v3ZJZv5qQB
AFeYCb9xvhSBybnPMquHtNAYPEYcKhOgbJFe6dPcBnLsmwWTiwB1Mbg/0iu090BD
jteHScNTfUjIOVV8GgBTpIUDVZrUB+lUKltP1bKyoPRFvSVODc1yaiJURz7GUzrV
tv8JgZwwkypkBDOKRFJI/TNuGI/xPhACVecZlpNR+2XKJsKwqrLH1LaZemwkPgNO
ebXGfFWnA4JAi8/bEPsLIh0z7tpv2Jiazae6UAaatO1EWMC2096IrPOv/ODHTRyn
rDbcAomubFnahpg4YI51zjZ92o6KnzlSrssOD9s8N1R+2QfDfmYbwoe8FCYp7YZe
D8ba/+JCtHVpNe5I+lsFIW8ufdh03I40L9FjIseYzJa0PjgJAUL7gN7IvAd0RLGc
RfYnianbl3AbPcxZYXTyKP3C3FWvQIqRhru0KLKuYydc6XDMr9EDnfjaHpzd0UMr
uXDYMkjcO7N5birIucrJg0shTvPzw8FK2gphDkGYIjb7xORX5IzzmwZgJstdOe1t
nIim309eA63UeU2ML58XbRwujuPWX7QOqqRXrDqqu/b631sGsTQPagsi64ConKEi
MK8p3XDx4y4rv6dw3x+nMA9LmH+kpYvpBsqsTq+IaBzmsRrX+33TD3LpWNLXPTl3
2N1RQylFXuC+gc30RG+XE3UkTJ7fmzo36AcA7BNFr5wdapfZ28Y1Ujbon8BA06Oe
KnnwHhXZhXER9MMePC3eDQv4CoU5TH9tH74qpu72YI3c+OItU/C7oam8Mc6ZM0/w
5B6r6D0KAKoSRIooOglaqeva2xCpL3T6eWLmV6BlCCxQeog8OI1/0itAD3Jfcquw
lTXmg8Hgp7NoRwYQ/iRKE52Atl6q6giEqL++WoCH8XWE71mcgCZvUeP5gF261/lH
qbOyCyHXZrL3BDLEJKBLqulh9XkM+Noh7Xsw8SbC9N5qTyzsn6cPZQ3cXYYlcsHl
Av+6fO2NqFZGOJKSFmYjqcrd6GJEX0+/GBhuRpC4+mpKWO6dXbNP6hvj63PymoRx
tUzVO2Ek3s/py6rWKTiuSUXTBPxM3gOJuhbK3KmmU30j1DKA3xI4Wac9yPEqWY6H
BIzDI9cINnl+DHoMZbmCc8LJ7SHb/XWd3DagfEndDf90mxavl2DlT5Myd9eyihAr
6lp5xeYMvti0yNUVS6DuEFr2Tv2C6yOFVRzVS2vvzd3y3EtJZ0oG5uUzd5dkngsM
lNo2gPKKZkAvqPHfKWgH/5A0ESmMtERB0Hjn6urvmLyZvGpiQRXdyyIhQFxAequF
F5lEx/8cEi2vmiWY8XIyXYFCIaQMOZSKjJ7zpZj4+BO3Cgip6/odry0yDE7UoFpl
5TAxakJzBDAI/F5zHUt6mLq9F5KzSm3Pt+1eRZZ7N5v9jPepWog9KnKG/+hMoMKX
fqZZaHbgCPTUE/UULUlfiwWgy7IebrA4fLbBKkrvdKvHJj6flM5MIZSol9KP+d09
gIGiEmUH/k4eH2/nQdAqoiCsjO4rob2I7EikWnqsyCuFpOM/hW1qq+PLuJxNULS/
4Jxs/LfJv0q/P/Ad/Acc3gXdLnM3kRAHzB+tqNjbhlS8NJPPJ00sD3eRJCF3Nu82
hn5ZjTlQlOKjEtk8itEJKzRbIOG4uvkqSRsRPJZ/dMpFv56Vij9M0KU1zltgdaK2
JzZ+sZ2yzMSc+z8BOlwVjmKzFNImyl8aTAyf5ltxvKTYMIPQLVNOh69cXF8e08KY
DGbB980XAoQdG/Fi8JJcQhZuVgCNmSKc33rOKYo86lljkiOcleENJ/kgkR06eVv2
PE+18DS0ed7JXcidIzngAiWXxru/xVPufmY9Q84illlxCXlQc8bFiQ83O3OE/SWg
zj0y1Osb9ZWgrn25kW6WHy5dZBUWaRJuT75jjS/kvaZsdWHABPVR8IM/RzARrmO3
5WAeOXtghHS8fi0iyjMkw33fguggfqUFm/LjiS1QGQRntnNHBkWQ+tSdJTjU9xX2
+JpEa7F4inMkAI5EYt8bxg1AfTtyP+vdOY0nSVrnmcxMnEuXEQkL/35cjY2cdld9
EVLirXXOC3a64i6o2q7RR20O940IiAUXFxjHEaslFkxFo18UBb6RewS7e0kL1iEd
imiSXrDgwWPxhNPzdHiD3+9ry/USX97tJd7aAgy/snq081/K3Qh1F0oweYuFWBZc
jhnIXXGpYGXnrELk2HuGira6HnFQDGqioY85z5oRcFIAhFaLlupg4KSOnmqHf6zE
6ftydlu+8JgIi0LGdzjlgojIltRndOjEqizmnoz+0Y+sVKF28TXpHvC/X8XeF6i8
Ma1odSQ8zWRvlsVQy835CzAGMax39enRd/upeaZmu6AmLl7kuyiDpI9/iHthcPZv
wH8MXWqfrb1kQ7st1GvGx0EAJ0EFR195j8/88ti9vxUPUXwFFGfc8rRRVsibNL5c
k6Yijz72ul8sEm14+dze/JcIueaugyGnHcwHgMKDOUq2L8GJfv61qjZfAavZb8HU
+NgG7SE7lVW92W37PmwyuVpIQypi0n/HcMSCvFhLMwmk905l0q5835tGxBjKKkIY
P2oDcAlfYHKMKV3oCCy2g3hAUvCYh1qCreGe/RRgJP0zzRX2P6g3PK7pX+xncrxL
OrsEiQgv1NFpkfOznCE4UtnoqxgvwmH6HJmebbALq9LMD94CTpbKjo6pxnYJPOtQ
lQ/jkrnuUq/IoeZcFRBdNTkVyziWryx0biPvaA9J66AOGgwQU9QIEy85smWc/xyG
3cVbNXzcw8ihoDPfEh17yB5rknVAAWBWwjJxVQbKiYqqrHYvKj0EqjMlxKRM3hQw
3GS5BGkDSCTAVrHLZbCugwtqEm8dptkK42vd1yKSNGYiCqOGoTXEqhnWhltvltW4
jaxYCmN1k3b9XXgj/ueCtOaI7YO0NCuwXZgCGw8n3Foa/Emgd3+L1hr6h8b5TgLa
gUvJPcsmUq74PhxL6W7iXcFKot7CNn6uSfcLLTwmvq7em23vWSCSdAhyYjUpfQ53
2jhwHTVrg3eeJu6zLpB1NgUdN6NsL68VRH+ageA/iFZJda5F9XwmQGq9mGR5uA8y
RXjO/3DlQm2JqdUOWZVvV6Y2MJdzBFYpZRdy/SSC0LV5kMfo/SOfinzuu9xo6MKl
B0+AECuqSgqOlnq6KhqDawNBRf0bguat/TvvCiq1vlix2Wq2S7+CaKfT8jWEzZU3
sSCifftCALsT7D4gqNQmgZiGv7Zxf2iabhsBpwfyBpgoakoi7zIAjAZAq62hhTQY
zoXoEttMfPdfaQeGTtob0kT743XGgzxJne99Flf7WRVWOcQC3sO9Fp9aRK1SxHpr
XQzBcSY7dsZKVlp/uBshkzzEmnuAAwuQ+5H2gyJ4xZOvoLBzDriMYgU6OjHhzInb
EzXrry99LLLd9QgkCOlALGdikP/RUPPy/WpyEYiEBpwY+b+d5VMD5/q5RS01Y7lq
DeLdy+tgFh09kVbU3mculb+7xwtNFaqLpuwZ0oki9oQ7K9ZQbbmASoGNO0XuKktr
RPbQnx827OQ5oiejlgMjf0oLfdkrfi2PsUkfajmizqfj6av57KjF7h6x1EziGRB6
PCc+hTn0BgNCT4bhw9PCibUnIESXuhawntyNgBXQDp2f8ft64ueWw0dyAtHozRTR
VMVX4N6Vx8QmZteipUPUqIWSJyKilYu5JDM0x220MvnWPmQ5Fca4Sr3FoXdRSxMF
VVhJNqCzoDpgCJWUzVSbF9ejHnYlTT1wbdZmix6qde+K3fgw3ohpTSlBM8vZ/nQd
zsZGtJ87AtyNbdX97thc0YJKO6L9Xn0AaaSI65lWRLPQq5vX/12a+OmWR0qNAEYg
XZBtZxsDae2KvYdGZCITVV7OgzZsZWR+YIXfnzin7DzctY9C5cIu20aFkv+hsiq0
v40yGs2z+C3rOTK1hKP5+iJ/Kci35UcBmjqqgBcI09suobBg0mQ+Ov0MExaI/K9t
iJZuwQ3wEbQQ7xJ/6pBGGvtlaEtitLOWDK9XMW4AWatZgrlp7Ge4fwWrOFDbclPP
bIn57Nv1wZqssIsmwzsR5lI4AXoaD8RTKEo4LsUOUA3H1KqyDVqHQcFwXy9+QjVs
/fseFpKfSy7b30uwwXY+v9rgs4H7TpkhpjinyKZD2NWYVjrvp2KDC90m5/EdlEp3
T/zMjskuoaXiTTcVBEGhsb6zybQqDT7IClr1xju8RjExIxeinQtDy1JpdX9aPRy2
cOvWWb0DM1scyx5nqZO3kdqwJsudBJ28r3xnrrAGmvtBEzaWfMOS7dsrLQf6Qdof
hIrPhRHQbn6NZL7ieg8GbXvRy51FWU7JjgCCOyADJbs2j3F0NWWyUHt4guh7WLrZ
h+I7Pd0JEKye9CL8EJL0MfyllXOkNLWBXZYw2+QQZowV/4usNE7wPBIjSHHAN0rL
Rae6GZcjDtcVrNIjQf4EMtsvUUWU21sc9lbzqdm5E6ai1oJPCl65i/b3TQqnDv9f
olGDw5x5QM57gLPT3Dcj/ZpPdscFIzt6z1Nod7N6bMRBpG5QBFHvnmfwJ1/9FGYk
7seMWz6o6NPGyczliReCuwfUgo1GldVY+jiIplIb1KftGn4EE0DAriV+3E94Bn5L
r+Az4p/b3qNIK5tOVzC9EyQNBwMwefZ0nDgCwqtJ2pcbXC2kyhFP/9mTTjbaQGzj
KRQq/DEuCWrQBXGyzbPEXPkLD5+tv1FcCzeL4Drxe2oOZzdD8TsZOztlszazQbcJ
RcOo4dJFQZ5vlta9zEsr0T1B0kmXNeTuRD+fxDmWGmlxSUf4yvH6CFRQJxIkXkNH
Eut3k/geV/7dP2/ilbGoTr7japakKYwffqo33ez+5r+Fh0OdJPJb1xeV5pDEOWZZ
oNtpBkFsoUU2T+XvhioVrKnJjPUe0dDAYAfFO6wZM8xj94f3g6rG6PQrD+l/LeEG
R8Ara25ID86wEdAQSQNa5w0pBaVjQM8/mTWzjFSIytUlxFvn9xp6ltS1cANgDAFs
M8It+v3EuO5PEmj+VHx3S53IZ/Ew53j7sSfhRaH5QKpLtK3BfURYKc9nYj1pGFvP
Gn2XMBpp80l4yTPJ8LvPfCGjsoB3h5A4YAlhYzRHVLOxJFtFMoh+fBpiiaVVXCFx
G9ucKNlA38uyJ4jsAOYKRSulnjXWtuwkNDCRFjWySmwNKlb87Je+Nt5izruOUwZP
Vl0dxuHSQfHTXnZqFgisfpOt4wQJEn+XHUNIwt5Sh9Q8v/KzSSj1lV4VE2tkEniQ
iyLYGaJrGjUz8cjABXpHKUzLVb+OGqy7S6VYRHZWDcIASHUg1nWu4yJPa9pfob7+
136AKFiUqi6z/eIJdqpXDMcD1LsRJhXpY+XNLazaNPhbZD4KXfX1VL+Al5q5NJ48
V7E+rk8w0v5QE/MdvyuO/GvGrZ8OeK/DSJqz1jqqQqDQvo5K7OvTMBSnsO8kEyg/
LG75rDwCoCI0oD6Cbps9WcfF6qVXx0/hMATccBAkXirBQ5ad4g6Q48VIWTyCg3pJ
sUzrPb/ezAmB06s9I7Xp+cgWa6FRj6KBoArKPSTiVnVKp1B7PdKPOX04UNLQsxRI
56uGxGAHx0cBcREgUX6gEPPqpf9lfz0WVGL+iRaQI809lAUO1O9wagL9SBO1QWiK
UrVDatB7bvXd0A3hd+81nA9g+QYES6bYmNQPeGpItVwCKtCe6CLv97a1S0XLZ8T1
/vCzl20m1nD21wgF5ajlP7DnPkYWOOwpv0UZlR/FyQf+7id7kn8Byj21UqPfRfoB
+6fQUV9ef5E9TJjyp5oD+C+jXZYyWaUAX8fxGsASVCT5krBOtgWiyb0ssvSOrq5Z
VsmEsNU/ltVMFA0PWXt68zVemm97EFjoe4ZoeZuXLI17g8SnDz+nB7fFAFq89zGa
YszUKwChJInjcqHgUvBJRQ6FVi/gBbwtX1bc+pFakIHjvj2WqRugkHlL9X0+VbqY
nP+h/WTuVfwDHarVx36QmDYUsDAhKLDdBPdOgxAegaUTBzibQMdfzbKFBfWfOQ1j
/UOfw1OYefp9DYS50gAaFTPs3Wr7KI0PkjQLF0i16aIlKpWdcQybcd5+yd/OyP8V
qGioFoyWz6Bfm9lDc1J70g1LvcrWoLjP0pQYbLNlPGKV3+XT5/s4dnraR2r6dZ6J
iGZXa76XeYCyFGxPhafaqL2oPXQt0vZY3YqCMI9r69DOabhGEGfm9Lk2E9/HX/4y
fLtmcNDAG3W+QbRfOINRObpf51ho668HRS1FE1kdf6GjeL+4u8p5sNmgGBni8Rzg
L8WgWR5AKHQ06hjg1jfYkV2599lQlR6dzInkSeyqKjrxV0cGWlM3NxTMK7lihZ4x
BQ504HMtZ13+rly4Gdx0F/gQjGtn760+oSKQV9WY0wkrpnzsWUvwbgh8ZdG1tHcn
0LpSNnXZhQGfbIbvAAU5aNKBOJbJFr8yPP3WzJMPlkyAeb9b+uPpF5+jv7pmzyC3
kGNKTvneWRESjQC3gd4ybaOmQ1tHh4SogGz2BzDh/mz05Sxh3MVJi6UNYdW7d7wL
ekukHEioLvmIEVpXE4NGdQSt7gjSkDVsXvCvkh2xhFVrVv1Extg5tWYsmIpIXBBO
yIgkEddCl32sbjS1v1JNMOZVWJjc8XnQsEeF00IYuF2k43P8Keyg6KcNHe9B+gXp
AwF+N1lgE73ymnhcCOoSkABKJv5TKW4PFNQqtF7JXopAA70qNwDbpz/A4eEEo/iL
orFi8CnkiI+v/ggZDhrSqiUKPOBr9jIXeWDB8+XXlYFmv6ym3dEHfAdhQo2AIyRr
rtvk+26I4taNk2fPiRleEOtbEU4Pgv8BwNNkoiRhSmcf/u1DBAX0k88EzFPxjkhq
OnojO0alQJTPufw6ALsQkgwWxrNVB1aDnSrPz/2SPf//M8RgYQpR5gdiY8mWsntE
Rq6btVrCI3iSEIii0ZbFYrkLdqAjEvMheUZcTpy6XXw5/QI61eZJ/SxIklCc4CUa
qh4k6bs6ZNjx83h/nKmWrmhlILHurJ3JGuMvEgviEbeLZkjwsi7ESOwqJWmbFbX1
sqVkw2VZUSwqQwJRzHYh+8GlUTGGM7FhiZnjP0888AbySf7LE9IcTJ+P49zKCnYW
cqt9TtH7WtMi4sWYRRNw6+TYOI5SplRDdxxQ7g3cKyaGIlWNIgN+LyyyybqhzWGk
zr1D3EOfGGLwTVChSo7gW4AhM42W1WVEpYZ5Yeedzv/w5M2ex6iOEvv9JZ7UiKZr
ia66vGwHtVve/CIaPgxyUZCtkW1pQUE8CJ/oMn45oG8XaP+tABRKQi+Apol1J5IH
z3OmI71jxxsYwf2dTu0T8ePm73v/5r7sypzTkteegnRInTQvfNAUAWRaiQ3DfmX7
7DU2N0J7OVJ6+HqVaragX2YrgckoFlojy+sIuy4fWg1rTtU4SkTODyjU2haUvT4u
TeSD29DzP/+2zoeKWCBeOhRcxEYBLT5wKT8osLmvsm4w7RAV15IX5ytWKAFVwGGd
j3gOqt8xcvm0dDIp2Ji1UUDBYk2Og/Rx/X4JYQyhiOHMBQMkl60jvkHWRkkE0RoP
RVh3KDowEZl5feX1QcSLw3Oddp7TR4aHzjq7DctLNfZ7Aoz33Dmiff3keEfYAkWS
nzkxCt+ItlLprwoccZwCQAH8+rPVNVyHgddMC/+xQSEpkk+KeZijWwrqvoZv0oYE
hya0f9oMPn222ZWPv97c7pVa2FfJC3EGWhVLcT54Q22V+muj4j1dOaG2IwF5QiV1
7Y19NGTzTDfVIAZeRJhUrFNgr6m2SRx5JdUFioMW7Ko3N8KQGr0d7o33WMjjwDPS
UkXoAw359znhCMaPxovPB1FTj64gMe/395az/lmZdJ4edSBzbWmW2/CD04QXntNp
DOY+aSALDzV2TWcGfqybMriXsBWSaG1WEJCO4BY8VXbRe7lpcfgx1iXc2kWMeRgf
EIK1OTWk4jKWSqiY7EF3xvUUml2VAR5fsj1pUhu/4ktPZqlwIl7STPu2Ow5EsA8B
ZU9R7lSOxGqqA++Mz2Tzx6L53UwiCG8J/HqfdcVwMSBJd7SJ//BfxUhw/VguC2P4
pglPSkx+lz0X2k+Uks7jQn6basaIUlOqewWgltXd916KFNiscQg/oVF0M9ToGpsk
YdR+HlnbQL0pQWiB0N7Dw/VFIFBJwGxUupgMiFN6b6E2+i3OKdwAy1zM6gRUq4yD
Bzb+L1DKOvwgj/mP9AB1rESJNcb1m3xqZEY788Gv5XsX1OF0wyMKk6+BLwgZK6Ou
MCy5Dd6yDaYHnMdSJ/Spa7PM1Cevk5H+r4Oh92U++W0yvw5CS7K0FpqQK3r6Edju
pG02n4A2TWeRdYgNCjI8pt3eW9z+I1SnU5eQLuzTS3Avt6hczMFQGyS6lBD49cDh
az60GrgEBM9SHtmUUJwUHk1b+ZiWHO/XtovCrWpzEPudkBgwpcbxL0PmbrZvdBdd
qN6keYfOy4tlHHmDLFDf1vywTUTuWOwYZ/1jxb/Jb8HvAu30I2rl8UxNgZeP1ng6
3BjPAgt7RXo8RKu6HFxphZJliQY+rH7lkaD72PzufrtkEYRPgXusIDfiH9lfGdQX
rajmaYtKoRc7nw+LaJ9NtlRjCf4DpBidBWSljsfMgopS+/fLQ8Y8daJ4hl+4phdb
oDJ7uTjglQ08aomDVMblEo01zFJp1K89HHcFXS0sNnFg0hFGtLU9FRSWk4UNJnLL
h9E3TIajFLQ6H1lBp4haZyoC5JoQug3E6RVhdHdcnt9Y3/UfZoJbS9FUqXJFqr4P
ROCu12ZYTiGZAcJzLPVEtbWqsY7QZVsM1F541Yl7tTOJSzclTRXxOO4YRGz9RONX
sBQtaH1lWQUb8z21tMB2susmTfA7cnzwh2nXewMaAsK9UAqdgVWdx0/PgEXNHG5d
E8XyDAqMcFl/z4SYWZMTnHq2nx3oN/o0TWZekmRRwJlqp5iUPOB2IAyNz5At0BqI
p4/Dnl4ylW78vZ/O+esiNO4bKxV6czEDTeUDV9jvjElFNHYNn4d4+p5WVoTS+LrV
2iOMV5EdEu3qfhIWxC39SjHwW7ykbL2j1mQGJDZacGwt2Mjm4M+62WYg+22yv/JH
TBrBG2ieeFbJFdI92QuN6DprxzHBQGc2sOIjtFzLMTgp8gYlM/galzrIZ5an1r/E
CTdPl/4qV05NQcfKIiXUlkce3cmvN/cSyif8bPgClpxuPd/+T385ByXxno7e+md3
RajqEPXrUDFS9lrQa8XQBFB7H1B5/lhOtXuCj99cpXfIyQxUW8sM7aMV3A6Whl37
XSJ8OKRAi73oIAiUmf8/dFFcUsdaivNnX1Jp8oH19rhBM/1/N4soAlhbz5nMxhvz
s7t2P8gAK+LK3jAtdn94jkInUC6oq4PYZ4gBF5tHAr1HHCZzw9jHVqTsOZ1Z0pSG
555Vw1IgGw2f2VpubeYsxSpdF7RXKIeJgGLQFf72FQ7V9havqrlRm2d59XjhAdgI
I5Z14XT65J9S++le2eh/w6w/Yn8JIq1yNPAEalXULErMDSjhRGIDb52wync546KR
lvY+ORVWOJ47mWw3WQLN3oWwRSsQwUyLUwJsc5MYOxjIkqLZAdunfubRiXINqvRy
ucJA4ia7kAnigL3mDlCfbQw1X+kkvP5r1PE2TifZh0DC+2Tlmkm8rlK2qIUv4xRU
Py3gds4y5yzlvO/BPAHc1HutKyVzWDWVtfB5cdjOeT6k4s+ebr/Q04RnvS8pdogo
eHLMhmpwe+9i+gHLFOhRiFuSsIuWETA6/3i3LVsWXjtMeRvpdO8ghuK7xQXiajKN
MMBWgWG/wGfOmjNkhUywG3mOtndRa5ZkaYi2cDeskqnVr/XpL72GzvDBwynof/mp
csvSOQs5z6gVDrz4CuGWcNkFZIH8hLoOj/QTYOSHXry54sJdSI5bflQA1Lv0B8SI
ybIsjDkBx0jk46k8FGWXmZdDhPWu8a7IoqW2gXfDdWG3erQOQZ1ssODLugpfBX0n
Tlt0QnVj9EHc8Gz0Gr6umgVNB9gtc9MjHm2L88GiWB9w32vckaWuLM0faUAATUUi
SvF1m42wMp6MxCGfxXK4lcKE+GxNtTr5fR/hUOmKN5bCt8A/bpjJvzJq6O8og4mB
FHqYA6LI1XNdSgvZk1YlwDf/hxkCBbYy7XN1+bGlSD2vk061Zmsm+PBgsXv1C4Nr
RJ2ZkbwXaDdAilUHuujr+nsMkf56OpcojzvzO9hctVNS6mx9tzwPsVi6fEAMIcRM
2nG7s9rHPV8X8FHacAAQpeYE7VLz0DQtW7iKoWTaFu6oZNBHRKV0aZtfUg+v7onx
XBA7HVgREwRcjgAtzjBGMsZ9LNOSX8x8l4pyjuXyC1x0UCRH8RieSq/bYaZBI3b4
frt6XTaJ2j1hxNdSztb6q26kXA1ODH1KZ5cVLGiOZjMaxmZMc84CwzcN03OFQLqy
QCiT9JtwnRW44w4atvCMFJbxNTs1OqLuQzO9FTgbeSPNeeG5/LMB8j78ax8Tcgvj
/m2chGiwocYlBYbcPvHSZdJVlgYz5Uv32GZOPbZTCcEBFD0W4GCQBM7v+y71dale
lq7fGLyp2gpDyhbACs/mRxX+ewET3q0ohS+CWXslXtBdHFgH2SJW2VaKuWwLxjyd
svX5+VgGrKKh0z2ezM4TFJypQAMikqNuiF5++w+S1uS2Zv/eQBp+0K1b5fjdEJyH
wnHNLn3Zd6jxTIZ9GwQrWjSARqwrnV2rGqLrISC8y5voanM7DKLqJ4MtAXpPBYto
C9yOqajsPEN8Pn0IWUG0tdjeoeCFJ73xRGzo7BSice9rGth3qlQucbodr0RfsAFb
0iEICchOYs0l72nCh0kRnAF+JEp7JxABuwFZ+o9GJHYnsCx5AQGE1rxYDU8+sdB2
bjlOL5QZl0J9EdUObdnc53rVKYN3XYckOiNFriHQeVAcL1z6/m60k747cbYRrZSX
Rkw4/kV8Yp7Xfve+cSNuO8rPS0XIhjqWOGgE/eN/GICJaauSFC6/njzPiqKCXkBx
vuIKLuWmMS38kH2S3RUtDljlTQwuuiok0qiBwiW3EHi/WU3860mkxMI3ZGyfhRUr
eRc5x7jlv2laBKIkI4C8zYDOSLQLxeYlhIN0p2m6uYsj2PADP4JhD0xHElpGW/Vw
t4Tpjjy1o4S96gkLOhLIkbxBaeoRcFjjEq+wv1+d37lZdUlBmkdrYjZqURCfX/WF
mgrhzc7DeYFG+OX7N4Eju3ylU1SsVbqmFUgrw4DhjL84BX+NZFWcBZ8AzoFD5hNL
JfOwNO5IEbcCfIGRT3a9ktovwM3Ilk/Dlf5mkcvzIbcNFdJUOQO1jbNNDdMuiL5d
YH4CfrlKJBXx2t4eKawPx+yMaGSZ46d1RuJs/sVixwiefbWb3xaLBd5iCP9t03Kz
jJ5vc7opEN5+iEci+WzkfraL//wnUpcyK1M0JiMocBeVrIjNSaKush5VH+xBRGe5
R7xmJtIgmCILY4IwhuLiedqnzE7PJiflmtmhOHDlO1U0XG3v+IOk4WDPHAmTxXJs
/Ta2FKkRJtFb77hljeSn3B2N8aQMxMJ1VmjkVBOc99hOaZbsHz3Pi/SbtrSWr9qL
BOPo08RyWbACxY4mTNGGPD+xtnZ8cakCAw4ZIOzKSpMYtb+k4OXVY09ECOCyCUkR
cx1Z29rYvNIrc7wJ5axjn6o/OQvCIfaK8qLNdJNkX7aOkjIiSPTKqkyWxQu26mwK
gv1QNIJ+dY+EpWnoqgbxomipJQ37ONqUbfMf4+UG5jJVvjdLdPAWI5ltVCuga1WJ
H+GMLGn7+Tc8KF3NuwdQLvR363NUrWWVcs9eztv5bAHtklS9DLckfw+AungBuCBa
qFqcGgMvdHo3V0pjoxaphgr4V+bf8WsdXGqe9qUIM6BR9o6AXtpY0c4vJzDYXQf8
jr2sfJjCFcNk7mrlB2zj2RkycOAwDn5hFbTVwg5kz5QfexA53R5Xzv85Eg9nYKN9
/VuKBBc782vdVGmYwYogwQ04kApcWnAEbBLM9IZPfUNT9QZg642jP1ahjPFIVTT2
N6pGeOUQmFaoLYEnFjbut5otmvi/4ZharZMoMumaSLJmA4p6UgSPcjrSyE36czhw
tY1IHEw6tpGKXGEcqDRoTBUOYjWN5dv6NuuaCN3g5nMYffvhDLkUHWK7BTMJwBIJ
kZMKHmuFsYhgvYDDUPmTL7QCVLvuUfKJKEKij1P1IYKx83bw+XgdmlGm9tbMON2C
57DtG+pYNLTnUgLwcnQ+WPiCEFvzqadm3a63sCFHIFYg2d9uk/oFbpHLd3vlEEuX
YwwJDlqjyYc5/rNe8+v7ybo/Ue+LJMO0kqAAQ+3GfFBB1tU+iLmJmbooWVLYETPI
AUnY9ienpbZN4v+pPkwcDLc9H/uXxdFHRXNCYuJNaIyGtqVDgOtYGR3XVgnbSFFV
Qf56nfzIktkZi+olyOXClyDkdMDBfrM7rs1F8X0jSz/QVGdVNPjh5h4M0CKBPoYj
CqW3u68kT5QBbLDu1BwMGcocwI1pz9kAFuE5+xxOHUkoZovNLup7lIRJnynq3lLo
R/HzTC2bLEh+rn1YfBxn+QU4GnZmfCNGT1mo9iWv52VSXytztp+OM+T3DnU2oy78
BLGnC/QOz+cdcMnQg9m274T1KrBd3DjGudVlEBKlqV8/IQMDB2rcpOPUSiuoSHXP
1j//bFHi0/uzJS12ylc4fLKO69Vg/sl1VaLlzUyV9sr+nRzySWDXMQgAZM9pbtMl
H90M8Rj1pmkKzFHJcig3paIiaVX7npaWjtl34SpsK8Ibqccobw8FXrd7yma+KyPS
SFui74CpF99+C1VOwodIaDACscXMdrHwcAVXm+WFBTpa88woGe7smwZ7iRzH8mKe
CKcnx/4cdWI7oZcTDnla+4DBHW2rmS6gQzrCD5DyreGAMYGd9aw4hAEm55inb0AC
ErBg4Clirj8T+XpCunNb/6kwQlmht/fGgUN/4eMufFVW6S1X9qy9EnXY3k1ESNTv
zk1LkJ9VCFlmx/cdKuaRSCf9avLvIE+y/nVCM6bAWS1JA1Jxh6vxdyS04d+sfwv4
WTzca38pnKfp8hS2IomY9Qv+EXzhshX5fUSEasyraFnjh4cW0igYHDn+2tZRixEX
64OUBOk1sAZZx479rkj56Cx6tmBm6a2YM5c9Cv8b8U7C6DIRbPnQzleT+BPTG5qX
YoMzHA+ssZ//em7ZTVtT7fPafvkNXQnGO36y4Vm0RonUXmRy4Yc1akJ2L06xe48G
2WXCGU0qPTUA32DiSfX9AFg9/sJEEsnYaQYuqzwJHczwmoGpVLBhgNy4F+KlfixD
0hGg3IQLIaNfJ5DMf9EfGSwvV4lw25mhQ6O6QJVCRQjzV3RHYcCBIMjnaN96Vmuj
sToYSUOoge1JFvmSBemzzo1eZa9PZD45vY7/7OHTt3YY5nEsk36gmUJmRw6qM5Q0
lgA0C1ltf4Pg4Uqcv8G7OukChXJopDBL6v4Qdw85wqOKgGYK6EoA51qsESWSfxL+
LhAoh5iEIsrKh5hRr6rI+NHyi9OSHCfQ+thnNa733G38qBA2DxrKUenGf893YifP
u2tCgF9gHQUgMu30DEgiCG1FlbHIcsNhpc8pObGdQnkDcX+U9eKV2AGEprQajPxe
nsbFRNjFefd5qmSZ1FJCHKj8wVzDdh1Ct7u785jPpwjEaJWWgY6GrShZ4fjLc8Vh
bP/JlKPHN578xaPDXF+JuvHfJyToxtXctVxOo7MDm+m4eW1nTG3OTMrqWtSf7Nwv
SYIKfTcRF3R8p13jtPsZXLtB0D9fylmlcDGUWmoWqadSP3iN3ZlNBlEvtK2/mIWn
o2ebtwnE+vr6BjZ4cupnLC1oh4uHL0sFpnAjJovaLHqr8DN2oJT6zgNjBpZTJ+XQ
pc0CGnSOegFfeKSoRSdw5FYTGo7/qMjmyCB0KBXiksw+Ep3nEOoqbkt1UGVFs2nd
77/WYgdcIf562DgkIlHFWg3RFx+20dpm+id9a3vk4/uHSH8XfR+sDHZTMGVDfTvQ
OM4tAhmCbizs/MtnXJafjm+K1wnLl2xfkVgGXc6r1a/7gKD5DIIBEDlTKip30GUz
uXJLjPHbiluabUKu0mRIaQRjLwoY0Otw8o/CoR3eeU6KSBdRAAdjswUWqbMQ1IvE
4NhxMFXlUx5jOVB5ERFSnE7XgY/XcDq7MHXKP3oM+RW+fHiiWuGrv7cq1uWOLArm
3Y90CxZotLh/Ofu5EGs7rn5Dl6d12RoxsPHw4BmUX3giZOWwsgrOXozcM2I34c2/
wdHM8wqsRlmyuqdkUo/I1OUSqrt4ME7vYk5v9nc4yBM0DOCQxNPOfOLMxWEROq69
VQL9F24SoGtSVjI6dAQ4aOtTfVckS1OompRnlsvGZFoLAYqxBGdUxUnvbivw7ABl
JL0RU/blS4HnroCvB6HfDjucXnuJ8VvG84vaNtACLIg42liQfxmwhnRl7evRh5pD
zGEgmgT4lmVZMX21IPz17jxn2YeRlYE+YHEDdYBU3FfD18YcCwM0Y8OH4QvJlOAv
nY4tf8/aRqp5vMFGdGBJYi6ExDT6Rgdy3go0oKCcsu8ABERvnQ+zRUYI7qW5PwLU
mzmDYSqSoiR9Z0cOBnwu05jSFazMiPpbckJF1eb2I39imJMFu9sq5sGczJAU/2zt
d76DoXk9dn1J6ej1hhpaGhu/5X/PIU7bsdKhFQf5tZyJyBYHFOtDDcKgFmvBClJk
hj408AZxQ8bd1/yeg0jpuOrfMHaw17sG41EquGhRlwTA+Ii0aZ1/Mu4AQoPezkb+
vMEIMl3lKjpgEIIoEn9v3uIWf62V1aqDSFxCA4LlzsyN5p2nm3D7vJXbR15Gdjrp
i/rKyP2G34bna/6fLxdG+WWG/SGFpz2+eVMkm/Be77Nj/NDOPk60FT72Uq1Apiup
CSuw6Arg5KgIdcWnmt2WSqCvAQxq7zHDpFroxLrGXIeRbBV1wDVncE3QnKl/yghE
hnB/PPVwiG2mT6oFJ5hdQLmxaI0rOafGaiOkw3J1r0TfgjVsI8Qt3fUhrukxc7T/
46I0/PIHelIq93pRDpEIIq/8fQ1f5km9UrMeiuLzGe2BEx0eBlOS6KlOFunoE8P7
l5q0/fMs6FYE6qlxdDojTzHcxhqUKzbPbRvr1mipR7b219+d6pkllRKesqp402Zb
2geAzJpqfbVEjvd6XOIXBHWTrBAM6YNqSYJGAj7VmLida9o2HOJPjzYzhia7/u8R
siYYDODwXOj2babW3iswT9wqLuK+pK0HZq0/pIF4+eNlMrUSk6L9zwQT+OJDSS9H
hOJnHiZDZKHFxQWNnQr2rNfMKGsayQt/bvSe/Db5PyDpGpTBC/wHrp3QXSTUWSDa
bFuVUE0wyi+qfnkuOXJJitv6fu9OMbizkzT8RLNfX33FyUPfqy//oIVHeqZzxQuU
AocTjcmQTDPgwOfuZ7EXj1X1LxDEjJmSsTSnW0FmCUUKv12JL7uf7HWERwaBgz/w
h+UMFm1680FsQd5/hSH1jSfK55CCKygK62fmfROBv5u0lvzRcm3wYagC9/xpSd7k
/iZYb8R/yI5aTRx2vTx7pT+nKkH9Fj/jfhobq1n+2hlufrWxN3zU0BU3Ot9WFo7l
sLKe9shunEny27D6ZesO4i1/3ppWMXbhX1fRZ2RO27xxu2dFqV4rWG8bGYoU78t+
BuG2X2Yz+pkSn3CVt9eMA8UD2V7TE3GxPLZD87IsHy0R8D0Mm4LTEEnw/OimnCmM
84WU4vVj8x+VpOAXux4dhR9nKH4fNNlX1u0Yh4hK/yuOFMaP7UdjPeR+HmM1bTGz
oFA6WlZmODBsUzlfL4MHZgDDziRGmtqDwa2l1BDLtV3mwcatle9i7GvVOr+xGlGd
+aPv5ur4L7zy/rY6OZhpDvNJesR8drUGD+R5lyPux4JRY2raS41ZmD8OY1EjtcYQ
cW9VAB+mgUZQuX0hT7yh8xcuo29PvZJQG6n9gtN1KxG8pB3qEUo96p0JKxBsp4Wl
4tQmsf+wmntyTg3rKjhupy0EEER6o85qsL0tzxBqjssMMvbBeZ7puH138cDJ9AFr
EQVTgOa568OvJ0Mu8sbXeixXrdxb+OXPSrXB3c2Z3P5Dw1gPdOPmPJVdQpfsD7XF
myklNT88VA9iunuEBlCmrn/F2QYpw5nrUbfH883Wi3byK4Y/3xBEzRqb2fnkjw3Y
hUryFGmz/f8t/H+QTU518rQJ8kJ2GVvOfAH1zTiqYF+imJ0FWSbbHnFX3eEH4SX5
Ju/0Rv54hvXMesX/3DzCgObSBAAQ9MsRfQKDJJ9YGa9ddvhpVWct8zKewq+cRWjG
Jhpld3nJAFFegC+IhwvE0F5G52F9jyb/E6Kkou80clcoq/tV216O500eNJo8OX6V
y/H4xUEhJfHu618JSUk7gJyCWwZEJmG9QK7dK7R5ecDXx39udYBzuNUV38SVc37Z
uaDL1otTSsBqID5E2tekS35PRUuzITRvuOsEOhbXUD019FPQun/m/rBRNKBD+09I
0Gkr6+buqAo1LbMrpKztPXWAuQjNzjKyxPV4/t7KMKdTeP2JP7rDmhUPRM/wUDXW
hVK+cs/R5q9mjjvtxDcmu4KsDu9kbfA0sHFBlFNLMddG/ysucbxb6szKkRspPSkH
cZfIpK7RqGB7acZMKvWxAAB0MClpB4D3cw+DrswBW4C+OO+mAa8koVrWw0wMGIFZ
EYT3A8yP9ctVF5TPbtrLcDMm8K9MXsy85WTUk6Y4Crg5id3HvnyENKEms6/YAXgz
TX/A5ckvyQiQyQFh4TndtzFkZsPERmBT1oB3jUen/MV9/a8L/WseGGagzYlvux5X
h0p2CokKlo6wISUeIWgNV/bAGBuZjYOSyhIau53n5ixC5MHnPOJvl6u4V7Yb73iL
2HjFU+zT1AaV3ysq0zK1YeV58jCpju3AfTDPCaGMCBmcQ216CKyaH4f4Kax539w7
WxYdvAUf+AgdZgxUqpN9aSR9OMRKn7RaRKyaPfe+3PV5lPMCc5xEPpwlV3+vd3B0
5ro4b6BEXw2cfF3dnyX/thBh42wZXwQm2leBGUt6BRNK3NJDlsJUZ6SGGyf260NU
s+Sz7/vRRRt1YSCl89VCKOKOYwrEpeuDbGQJQvN4s6m0Uhp/m1zJKKkLrcUjIPb2
PoujFvaQXZ5cVvjod0vV6aorkn0bkWoeRwWm0E/0eSzm0qCClPSbhqw4OfscVqAo
dAjsR2jNBSNuXw+XR57sZQ9epRADwpw7kGqb6PZ+GSS+EwMHCU6D4xgGYhz8vRjv
EPb8FCCJAikuY7fDe4a9/g1uh95kPlqENrv+07rco66ql00BOaOLy8IuELGaq1ME
x9SdLx2b++NSLRia0LqDIuMMfhQ0XiU1GFBEg6fmrMR4CnbgjP5nrsQSqIqjU2Wq
/6X3ocY2E2vE+1v1hLQY0JjRoWlmsqA2CM0k2P4xpVhf71thIdYyu3DysPt6KQ9/
BeaOIFObFKW6g6adjbVwMA4hHE5AyFMSJoUSp+0Kdjfuu+t6K5K3cE2tZmefGseQ
BWexgHuISqz5fFUwmHx2gsWqzcqZgJPU+eMSAaI/8pVoeLtlsoSWlHB1Jqm8J13g
l5gQFLO7hpz8Bqh4efJmdVlm7cK87iu2KQ09Yf1afZxZpl2++QOHaoflJwAQ9OLm
+lhwhv+JeH8nV57G7CbhrCMXzDIdJGtX5NAewS1mmVvJ1WhD26CcoOTk6oZmzZUa
cdhWK7Q1LimyP22h6aiO9QiKi2VoVf35MXZnJwlh2KRwGwN+uwF+Kb+55I3isPac
V35L5PuVq+IeFPIuHdSb3bJUkOPzkke4FcbTOlHphBnAs5fCaxVHiaFc85IfAbXn
+Gbik1kuAKGIs7UIlDC4d0ajIK2zJEm4xXmqq2ivBbPFmJPo+9jtsBhD4tSzg8Pf
p5VnG+MATMbicAwKFv4T+1xRKNRlirOw4pBVQuBtIrNwavNn+dVblorjaEam+dCU
7Mg9nqD1kwC2heAS+/OwVcJI4pofxOqgLxFoWu9kUiRZYkOLBAV2wAc6LvIeJ2c2
c5O7MtQzpn03a4Q3qppSBaNivbJk+FB29e2BSfmuy9sQPBK/ub5hV5oToYuORI6E
+ET+GNwXZJ8la2GqFMZ67EWKOE4IJSg7ESuU5q3dZJOOxOc7YN657Y0M0XTxxBa8
BkbYmehzrQR5c+7x3/RbCQDYWoF9eLOXfFwEyQxTcEK9yKIDGtySNoEuX5KYPpc+
9kF1qnNuh7QEYGsjh7BytE4306Bqrpmjg7OZKRQJQWgYqRu63XA1fzw7frCMg6j7
HHcENadTslRMP+g/KQLYeHKhqfzoLukHDzW9UFtdOymQmCuQZMiFZav7BQASe4vG
7mEeVWXZCE3rLwYfO5n6FwjxfOiPa2++GP9oif46thEW1J+jWimlzhQmbihl96Lz
l3ZpJ12snTdFTRJToYBir+J9n462gf03aCBkKyGvW7fCmAAWpwaJJGUw//uonENs
IRL2n2DcYCGFXgsIfeqPix9n1+jpwt7UYNEJPqY+240rjvyA5PWO/053w5N4uazP
CXyvww+dFh57AN3MauNeHWw5115+ANLEQh7R14dJI8Ac9PHOm4pkGT39TocX6OJZ
2hYB2HhHFqBINZC6R7rM+CIfiN+mA/9uVnji0CIghIlDIu2dhypQmn0mCAPTOJRu
5kj8B8vnm4Y38g1CYCwJkXprzxzSs0nHG+KmfBxWMfZrvbigyOiB22F0byc8xcyu
qz7aDCJ4x1NgXY+j9OcqmdhQKXivKi62F/hN5ILNnmYVt21JQGmOvFg18bPinS+8
uIIKo5/R1CEcAHMAOzzvX7f/F7MoayjgwxFJ7ePMFqjJLIc7fkpzpb+ASt4v4WAB
05CfeIKEnu1GgfiZAW8ZJfhijrDkMLrEEClgkk5QEsOIgzUTU+FBzYSJdF6VTu7u
vgiDiGMa+lm+GDY2+QggjtEMC6chQASzh7sJ7heL1ernF6/P/2FN6c2C15y24RAf
PmyQtFEGqrnEj+xUMNOz/dOFtd7f6zx7vDFWxrJ+ymi1xNIx3Id0F5qs6+jvpuR6
6M9nw0yOgfU2rKrlzmvCU8kBHOG0CjV37WVv8n5B71QqO7prX8You+NCcVt0el6f
JZXRX57r+SgUeW4T2j5EHWR/HCvi/uGvOrFfVoIJoHkjJYae2LfA6OpcBbNCleFf
8dbGkg0K6YqZR9+u6q6wpeXexXCU3bHshPPidLXTqw5RUz09aCoFl1a4L+jKgFBE
mt+GwogpT2xeKsQNuViCXJK7VE+v4fDrIa1akOYsuPpE22iF/bCkkvl6Qho4Etws
TknS1T6aiw6DTXGw/Mw1dDMrvhpW6juvOKPvPwizxiO7v4vyqQo3vqsRpa6ZJm1b
nJhL23WK0Y4KsWePGA5HZmCMfzWvRou2TCnvlQ8TRArQl/+ZQ+csMr/JsrEFU3es
ccx4VLstnvS60WzMSA1b8Wr18RV+1hs2xiWpL11E7pzCTAGMPdW4GUc+bKbDrmM/
kv753/u584tst+H14mGDuJVhNmN2/jPVmoDAG3Cs8JHD5dGhrKsdaE93rhrJLQD6
mXVZ7avWwYCoSFWjfyJ/AjP0V3MDyx2wEY2sp0LKcGpZDuHxe0+uTKCKb8NNhqSs
QGC9/8NTapyioXmkQ6cHnxIKZgtNjmSqngqoVZ6/FKpPBA1lYAfBs+SwQLr7EuEe
DoTFLAyA8diyn0f87GwnDv0IOaAdEghy642dNKnpHnZF+YZLTcLlsWh5Q79UqBFI
U2DXh6YNymJeUL22vA16S2HBUKBnsZT+XoE63fOiP2/8BYojcJqUmxcPzAw26tsr
5+acnYLHgAJ2pENvF9ESniCBYvOGXrGKl8XouDcVNExbf+SicwvjC7NqRDDe1lTW
bIf3T8ZXYnkmHzT26nm2Im4waswHCu96dhmVuxFgzq5eWlv/GvkYIXt2OtSw9ZKP
6G0xZEUZpiHYXUBqm4jVWk7s4FTBUdyuXiIFvr58pmQOvroS7i+dcE8zb0+6GChA
mj7IGcnABDFyEQMx+SoBB2KC05ymxbs0+8mHrdEsmPatJLLVlXbrycdX57JT3CvI
4/TyJPn2OburcsYuxu+bp4xb+MIvHgy1tP6euoGiLWeU+DIlV4lDFid276Wcoidq
YoK/eiJSzKJ0w8zPGifhs1khx5r6mP5P6nUAcXX0v0dZfNuvntmf45qpQ7WuXe4u
8/Zg/5TcpZp2mInfkyEwCmLRJnR0YukQcyB5x87H9tx1oZFDAR5ZVKkh195mrnkx
6J1oySEikP8znSzJU+qY5fwT+f4ZWGZcPSSNKAR2rv2boHUzYWUU9a71nyf7Qj34
NgQVKDOUFUYx9nfqcHjM0vskvWASrmbZ0YghJgohcVjBblhwlqbpMZIed9V3JozO
lBCIbvkMuN34NaQUg0+Pp4mO2hlahSoUQ+iM0J66LB5vDKheTyGEJZqoACdAo7jM
YoGek8n0fjqzXmTQzY3GxmUQBbME0O13zDoiwMUOk+FprQOsWuCVGOjiQXLVIcBg
zAR9JjkX0nycpWuPRwEp8jzCR7PDFHlK9X+cLV3qNQxijnNpVKcbyUXbUlKOrXIB
0jvk9+h6fJJsrXjuUgIJ1GeA6hN2hUeyiZmFTuiMnzYyHFD6x8NbRc/cwnpUzYRK
V2/hppEZ0Cb+z5Du0+y6KR56AoXQw6GWBiUm3n0SYzSJxF5H30kfMopq4w42V7dy
aafK/cFXhnRVBeJHwZ7lbK7npbLOpagdJyARlnYZU7jgQD6XoNWcsJobp/DyHY3D
B1PZuAUPNcf8rPjL79m4fZ/LLyFTEk7Q17g3y1xmek1FryO+3IHiriaGShmJQCam
RKIUwAP5o6yMVRp3cHNR30Io6tCe27BOA/ihMQsybSjTthYxo29byBFZb4Xmgei8
e6+QOBQWYpwpfJZtBB21RCPM2FKUpiWLASvty7LTq/KfaKZeO97YILky6Jysgf09
mcCRthz39wUrQgHz2XVlwkZhgvDKKLjdO/DIQE3Vp4wVOPV/VSoU4+uSisqmaoVK
b2pS51YrwiIDX6w5C4b5RQWMzj1NaISPGgaySp0iU8LaMnVjqz0gED6yrSeke4E9
CoLUJG1Z/rDDQ0N3gD1rb2cmjnmlTx55NSMrlawGWTHvAoNX9W/gYGRqxNFSca/D
bTsTuOdaqE5amnD3YJt6Smly0DqJPGSKvHZuzukGPXgoQkm72rH/A+qlMb0PKrox
Xg8zyQ1fBKqFwILrTyz3hcNZn1B+/Nmt3YmgZn/NSyePeS0WHU+NOTEWmLVNnobD
dbtBhd3o4FdeVa6oZmt0kY9L9j73CBLCY3B0dr/SPdrsIvOUM73bWun3BT700+SD
Tfk+Z0E1WUjpUFuj4lGlewCkPEFWRnEKLkf8ycyVyigh3JthF5Ci68SMlrY+kWox
kNLCG9Kz7iCvxsN16HqPcFcdx/uaub5WyujskFzm9rGVKjQdReo/HpJ828B03zQl
2qZlXzzk5XV5ZPjODdMcABpA/K5iS2Ut0Eh/E6g7DQtIbmGGc5cUGFECh7auIirk
abkRqgvUqE1hitPcHttwaJm5RmeavtyjhpRjR8tRXceW95BpYiTv1hkDB8y1Jwzp
qA8bm9ZURmgbyfxEoDEf9wDHmwql7C9wzK7/4hHn2X+RMCI09QCOLz6zSRkSRbx3
EURWReuySJQqqW3OwvXvAoYQHXquRvYEIDH8AjGy4AZd/pO/0uMqyayrgXQtF8pg
73UFOtb0Go7va1tYiaJfpxbyo1IYIoWSvmXCq6bL76TfdSFO+AXsMFgNfiEiGolh
0bk4jEVQrBDnsMXF8w90FE4pZaW4Qya2h2/cTFqIaaMcBgvMhpyA0mb5MlKIU1E4
/pSCeOtlL6USVxMxLZjdnOalIOThPdBhJbSQwS/l+si//JLFDSZMGbaIbFxo6V9g
2tyDjPYHyPnWDlh+4AUO6ArG1UCaIG6qQHopGqHDJNvNRzpF3t+LpFmGW0qA1E//
A/7Bx8MZ/Twncmq6/IO8Qv1ri5MQuRHMereHgWPkEsX1YcTiy5f46Ikfh5Ku/EJ0
h+uoSAE3yAL/mUD+sy+LdizNngklrhaVBYgpBwF1vNvrXr+5o510Cej3gfvJ5Pkl
oOuRPx5VGLiqQwhuxjLP8nQ3p7nCbGa4Xa+Khviwq8S/kaMpchgFrM1OJlGkwRs+
AZ6qg7NXWUThAcY/DspigdiQXyeUXISZe+JeQYcFQUSHAYBXnksWeMQusHsYCsMo
Csc9gbjzoLBcP9DhS9QunBz3dHGnSLJqvc2dvov1R0AoqIaFVQzkNt1quCBlPUQS
Oqaj3LVW2yi/YPBdZmoyGYoT+MGmZjWAL5FrIGuoxJNFFS97V5qresjTofnIlINy
OO8NxnqzEQZghjk0WtKQ1HCIxJWEtOpTKhObHaZv3eZEeG4SVPQMVC5lD09KyPkL
uyMXFY4+r7DYdjsV8tpu3eJL7Pw1q5Vzdcf9eB/RmDumJ+ar0ZC5X3FI6KprL2+b
lJCjXL0qZuJWEm0nm2dRrWA6WUpiyq61HRs/d5I/MMDHGg0tvOsld4OfJcNgDSf6
znoGqLyAymWaCZ5GNNeY+6VWLJ4G8By2wwimSQ/j2x4kHa9IpLPEPmEVaR6pQqkk
vbkZJ48enOSkZv5/y7EaIBkMwVx9/Uq557+H9X10RRZbQvUr8TI+KNUmpxhFOFme
lEz6oQFWT8zLv/48sta4XFvWQx5p4qs1w5NuLolZ56p99dVocjlxi7tEby/mdHDa
knzUwFe1ndoQjtVwMBbx+D1zwQZ9eMZSfWWH8KJdq+Uv+pGqvnlebR6iun4i4hin
11vOxMY1LsW1361WItbGER7sETJq85h29pK+9CghhxUV9+/5EBZbaVjcNKVNQOlb
Xv/iU1edJyd8NivsltjaQSSFbIRbz11rq0Amwci5jDRit2c6CPHPjbWd1dL3M/2m
V+SgTZA+cCs/jwSTbpWcV3sJfviUFaMvOKi33t8l2Hk6b/l737CIMKN9CO+M+wdu
qpS8rsOfUo7WmwEVRlGIuECp9PaxecI/Zaz3EnngSJg+RlG7JlUKK3DwuEmamn6Z
G4siRXx/6A2VtLjKXXnZ8Syo+v3giBkYaWmI1jcxDG7l03ShKHDz2uKSem+aLrKu
Z2VXocxr2v6XpyircB/MZbXt45h7SVvw4gpHPXB8Ti5GdP0JFD8KCcrUqufQk5bA
SQaMnA0FSPV/WRs8VmDtYwckcUwVI2dR8tQ8FR9Ywp9yzD+NTcDrPt627liY8Yr0
1jUt4TPwpiWJk8T76Y+cCzrog6kfwVowvsvInqGNyKC0GVWHLb2pJhjoBPgg7nVM
FcV7HvFdY73B0jWtRoD6nKT205ZtCeq5Ys6slwBFpY72UZgbQ9Xd4MOTWkFO/x1b
+nUkLiVs7OR52uzptSd58AHiJPlWJXsXV8MYQEMqekuiCj19Y1rcjtGPTHJC6wMm
GvVi0B9azig6PvvnLQKk8R+LoC7teYnLq+UoInVHbkhnut1cA6kNr93pRdD4zcw8
HqjKukRreLAfLvL8lTuD8/YPZLHmOFTxmR7Hl50csKcP9acHRwnHMbXz7qkESQ3H
/iIXCqfBTsM77YW016gzJ0aHP57xhdZ6+oa94n7HMzWMXyFS10mwCC52VzZ5Un5y
VXChaQXJ/IfHPZ6D41wybPlu5kHlw4lgOiNEtqnsKFSX584hhWj7mykVlZqU1Gqe
kjLiQIzSKr+RALaT6006tFmd3Kd8nvdyyG25m2gC+eQQi4VlWqwTLX1dMNVjZFz9
OnJyxOrY2EgN0J5ny8xms45ZHXZ0M2Z/viTGb/gXP1R6uhwivZcqHZdAQjoAPuEQ
8cY6/Z8KxhFdxZgzxV4MHhd32T0Mx+G3myF4bVCJ4DkriYnbBO5THqnJ0fQzJFeX
6vySTi10pmTqkcN4mGWYdjQ+jPSwM8In18uE9/56VJm0vS7Xin1aE5GuLgauXcWn
kK9/IHx5Cv0FYpxvxXthFNmSavWqhl2IG9qh9kWBmtp5NUFlN4LWwIPwW+pu22/Y
IGy81Aa91Uiw0xJLYsnNpd9RhnFbJzJP44aUSDumfJNBqvSq4QbmMS83jq2FQEBa
HufUwgTK0P5zd0EQrH3aAmA1PXRG/OQ8gHsQ9sWgvcenvzlzZREhhEEAt5od4rLS
TMCwwf7UKqtlZpU/WTiSlf8kXsiKR778vCsSmGRMq/0WeuT20SmTRM73NULNa9rb
o5gWFwLxzPJnBNmGDeDWH/NsH7yn//zJI3QARTvz5S3uWwmJjlzIw3VuDlvgtsnR
IXzFnqK9HbrsNXB9zqJlZ5JACyI/fMihs+3N0WzSjIb0L4DP77WKkVDQKZXW8V7V
aTdOiI0vFuwMQy7hNoatHQLksw6EcEh/2K00Soncts/Rl9VNEUkKGtP56SD+X/E4
IPgDvT24fjukqBQU4s/UAQIe4wZKu4sM3XYHLjYJytXWfncOuOFnv28DxP46jNLU
t6F+sktfntQr6GCyXquVaLzK9bD32QD8Xv4uBIVizt4K76+cVaXQJe4Wgcyjc5w+
F3eHbSOC+n1y2+KMuhB19tNC2jpEshYPtab3WXA0PKfNCalb8HWR3Sb8DmUMDkST
5gXQBOMqGh/pvKXhSQCrZ0/QsF5Q43H1FZQdnelPw4l1d+TkMWcb4Ok1v0HDKka4
zQ5gX886n2bKMRpUhmQhs+eOirzpK4WV+2MLjvtFFSc85dozyDifDV/D0Yzc2JCs
Yl0SK2FD1btkkVSKDRhACDROvUNlGGSafv5ereB9eFExsf/Ec+hUkhlNG0abHHL3
ZYHzLezotW1FKZnrhn6t/23xleNle/tOX2CG5s89K3wKh/2rdHeCxW1DtPGV+azQ
otf5WXiY5ZT709Rj14Hh/QRTzW4KgRReKy1K2p8TE+TZ7bBlSRvuWvCVUNCXP0UH
dQsQPnXkcRFxudHLxVGLGrps4lGQh9bTfi1tk0bVc11gjRDZWFdzk7zMf6EP3xcL
YCONy7Mb6OGXjJw/FadADeq0sa4co4H7a5/cVyWPcvy0rc2RaO/tWoLjLxLgX83O
mltKZv8Qcs3Kv+Rro/y6WmcOWt31dLVAjxhuqf0BBe5IAlDB/RTjj1cYHneDhBbd
doOLNaJern/JOCfyD7sKAFHanB9L7GdhIlE2xjLpjb2yaQBbX5P9aB82JKCJ8V49
mp0UwCK/i0aYr05CM3LXIpcKezG+qvkCg/qAlaGeFowloYyos8NSvmW8Py8X7zS8
CP/xSowh9Mh+k1kJPXcKJmKKQTvL68TLyhfsgqOcM8f0LWgfnffb4IqHSzL2RwZi
L++aYfrZp11FZBvwd2DEvFGhH+GWnSdC3KxkWx9kMrpaJKGLYb8PZH8GRBy15FXP
qz6tUIgP+ETt6DSV72ws9PIDDTayw3d/FkVzfL8J19Lk/ptlLaASHR9Vom9gZC/9
7MUB36IbBJsoA1UMYORVKh5G/imRB3rWxk/WcdMor5xsaE4viB2/lxpa/EWCRmub
hJmINVo3xbPQ16lAfd8p1KVdGo+Mbd5Shx05Hon9Y79jtskrAq/LpJA0dLiGtwsD
fUUhJ+Iv3kWQZNt+EhV9EutPWGxFkmlVQz7XgsVWvfs4BI57pvMpd7+6NOyCpyCe
x0liWi51vfYxl0rmgCf0jPMpaeJiolgta0Cf9NmI5BuUaNYjT7whXGvzI6JtKyJe
/pXtdWA9Lo9nAKNCklpoMW+VRZLiute/Td/ZlYP5uKJb+qcqCeEfQBf9aRZgAKI7
xIPidOhr2n+n0rU7U6+AkGCY0Oi5eNmUVqjC9AKZfXi7gTkwVNMYezvKqf1z/qYI
IoEW/Jm6iaSknI1TR2DPxDaCG5q2cQu8ZAA/hXvp4BOoSwFsuKLZbd9h6g+W1Yxi
k1ULBIROntIGXQRiiFlYTTd2jF4ev6Hd3VOJWs2fPoysNzJyj755khgzbWNbUMmz
adkxGTgbuzhRN5dQqqZUQDDhgr+sUgJuSCSBSfgGOFl9XOQKPxJR+hjpYYWQ+mfJ
ev/enESAiLYVqDhHO7QhpRBTeqa4Og7u+7F8V2nAaRZdRzRrPxkBWebJgMEi5FtH
F6Dkh55yaNf9O1niDs0rP+KrMQtVjboOY4OIMMmNbrAIr49UgNIpqeHpIpMaljh6
VuhctQDrpzFH1edpycJwF3rf8AoccYFUux0OXGPAx/ZvX5T/TeSAeYhJV1ZXrLQK
Xkwosa+01qeaagsiaAZRy7Us/MgAwSLsS6phxtlCDD5Cmk9S/edpWEjSafK9Llbb
OgCscEWbSxU2XI8RBZw1VJf/Dnbjh8ir1qooDUSpl6ixYZ7DfrqX6m5hH331biZS
lpK1y27OO1IrDmj5sE7bMW3ewFqrqUBz20ci1OqJt4YX1KRQuMIEZ3NRL7K/pCr1
BOvTvaB2auN1YE3c6LQgLFtcpRRhvtx3sZfTgeCxY256MmpTQUV0d8cBwCWt9nuz
9Jazzyy007CSbyT+J2kmuAgS9kwV1ag0LFtc/GoTrfLgymQQRv9QTuTlDRR4iFB9
5w8JOZkKUh430okSvp/mdNznhW5N76jKMGvsU94QWbcEpJEuUsQ1DHArHZgL3bsy
0i6yZzSBtv+5QMwC0Wggi78OQSohVMCeX+0oKnBzt2APw+og4n9U2MTDjgQ/BPnx
ZIca/lG9XnxGM8+H4IiOrIT/Fm2JMyxET2/ZvXQIAX8DbHL2kJT/OBdDu51dD4kC
wEp0P7t4ij+wcU8i/VY520qAf+r1AnluJ4ro+JXpWHllAjxKQB7Yng4Kztyyrcnk
C4Sb0ioEiijiOoJgMwtlEFO7cA+Krf+yNHPQDgKidBJy+7R7nTUwnX3TDjwTe2s3
Af37nNEj9swk8Yqrt9o/w5b4DleQqG4JfcSD3AEyL8WYylLvrhWkm6PVTk7FxffU
m/XiL2aD6zyehTw+RF3KigDcLpwYK48AjlYhA43J2ob4ykSu27DGKky6fFSuytl9
8pLoJel0A03EmB9NSuc5mrZgmXqJdmCmJPFhtIKJ6kWk1kZTT0z+WSf/U5sPBRpQ
+D5TsIgEQzm7aMecZLmBCaRn8XoQ5ku16agaSWO5Y6Xb8rFr9Qqj93JeBFIFwD1v
AzCLHW0duxTKU3sRhuXJQlwPMlHOkPb860kPfGm71RAlhKVnzc2UcTFrWY3Iie61
zF9NBfauj7KN9NvhhJKICIiYA66RzFPbFKCzDFzT8RmizYjhuFt3/Vdbnmj7fV3y
WM7ui92NM9FCiAEmaMOYoWlC2wzqaNrc5mJT9dCby5klEJ/2FtUZfvXcXYM/OY+9
IH9OUUclqUmIx4WoNQRxpIFNYUVcIbuxorzELD5fiKWZyONup6JrYA/WjTzjmTV4
5S9mOw2zQqAXrkMyel1cMt42gU9rJbCOtjAObTLYgCE92zbWLWFDIo+OlKKjBk71
sdGS0dEhS195ocEqk7wNw+jcnC+MJKh2HLkKyk/PLpuA3che6Oz2UuKMejR+4Rwd
Nt3VEfbI8QsPvLDmP2r4WetNci9DXFo/tXv/r7vyslkcjTQcPaLf9rMsPeTot49P
ShLDHN/6Ke7iSwexvzJsrQFmfprjLheEXyb/4Lk8CBXwK7LYZfPxkbq7Y3Mo3spI
7LytCicKecbc/fDBC92eBkxQ0V3DrTTMUGhIrg0K3Z8KeDT5v1SzzLK5Hp28N1Ev
0LSRljFu7kGihCk7gN4zf8o3hNzXUwXaLEhOUlxW9Niyo4PS+nHNbgITALqEkk9H
zy26WUtiini/ClytEE3DZmo7obyWkvKanXyjQPnckiDGdYWw10ze5RSCjCBr2Mbi
vsg7ge+hcwZXaFSKW3FM8UtizqUxmalX2EXmHTTcsxLxsZ5Be7X7h+PWCDeSL6rB
cr8bZg4e4fq3+/jNgvFoI9BaYLvtaWEEccXU6iZuY8VMPMigp8QJt082GCpUFsZm
clKXcBDiEuoFkVVxf/hDQ5+04nl2SCfk+yz2jrf8dZMYBxsWQ5Hd5sMlBys5vVbY
TEPVmDQ+fpehrs/a3ZC1FCpQ/lN6f/HN3peWHOx31Dx2Nu8PjXHGvoDQJiHFZlxd
FBygASkM6HN1z9sUrrd7nGW6sPNBBpYQrBCn+ja1uJlQe5Az6pMBVoDx7UiO+9pu
4DVI41UJ/iRMWR9szjVIjKp4pcd/y007Yy+P4mIwJ96rHeHlvPYfvRKmJx5w8FiX
nxTGHYIuOUEyqrZY15Q8frM9I1ySgFFLilMyGpi4h9dcOHzzYIycNtMmNxyvWEci
c3gqLGjR0Ms248S7ycZJ/M4Pey4RoY2t3u7Eswfzs4HHeMheFrcLtkDyuUlJik9Q
d9lWb+6WnDKyYDqaPEnxolkk8PkGAyEPhsNKxMHd12YBlYfJOhg9bVNPLnmuDZbe
RbA0iKiYjPKCeOvBti8uiOSv2tuhPm6Lb4pDB0LIYkfRp00DzNHzpbVObUTy7WPv
tnfJO7770NSKjYRGDQ5le/5j3ZwvM2q0T+rtCR7QtEygIeBsNaJuD4alZvbjaj2E
rYhVn/AB4zqAFURKVNMQG6z9AT7Fr9g9RiW+jmkVZhZ6PC8lybxc+MuDWyi7wB/l
IzIslFwxm4iMdMfwRXYCVOi4Mc+7lPqa+Qt7ewka8zksQsTreL+UHyhKFSP6mkjW
ZPrXE3+j1gV2+G/xf8btOYfEvjkGDcgo+W2YpZLNGC3VFEAR3rAi6+Dd3ECmCgFX
e53vYIH0wUD4LpYrRXDXmz2lgeaewE3C3xnsPaGIZiQRUEderf47r08naVeQmWBM
XcevA/Io/+3sEaN9+Gc0yaSON0kzTR6I/6BzW6GeZk3hWfxFRfTTdqakPzLpeUiY
8IYHXTQLJoNoYCxv1GgMYksZV+L0ElL3gQoYidccA+9bQ3Mkl1GwDahR7z78HKMN
Zdko1IQUXOM8OhXszvkm9Bm5hLC+LE99H7HsvR4xJN9OGom84urWoDBz3GIYHPBQ
nD1qJiNfX+44vGWpFFLWXaV5e5/B1VsuoN59BQGMY/qq3jsrFHELP+jeNX9q7SjL
hkFD7uO0LvTptFrOpLNyd0EEU+Xwvc8kT/fNziH3UiXDoWm3tvAKkRDBbIsHBbT7
Dlxxv+clHzz8dIvMEHAxqwg335qKn6X0gMnWtzUrp4agKJK2cLhbsXuoy4jnadkm
mavALthAyMQUsATQ1fCNbjVeW1AbXdmiAE0GiR3ehBK+8Yyt26qcCcoBAvrPgIuD
bkhUTZU3DLj1BsKK1sjZuNJymQegje4XuVD959Q+38aunSR2Po/zkFYOCPDTc0n+
TbQjvO7e0dr1o+IWK9CYxzHBI61fzWm7Dd9Rqz0GMLQhbwf0NZ88X9A1bwgPHiwR
/4HFjEMBwXj3Y5IWan6R+vwGC73VcUHsazh/qw5BYJ3tWw8B0Y7BN9G0l9XuDaDP
9dog08ASa2PBoCzPRgKgZ+RTNXTHi6UAqsrGsfH0x8ba1aPyQbcfMYR4LfTb28O8
P0mVDYpTgSjN/glmqWssfiJln+W59SQ5Ft797qQ5Q5Eat6GokR9IK9NEHQgZltiP
qpSFOyPMaVD1XP3UJVo1m1mgVQ04VLZSipSkMUkgcWFVlOJl9auB6mRQOh2aXy6B
d9LxTRRwXsHSL2rL+ZI9ZIPn4X9Gvp0MtDXwRIYf8rj5LBZ3kogJyXR55luwUUyR
I0axFGh0DU1G9CnxqxPUuLU7g1jhrFAGrKyha4GjkHn8Vu0gNiSynG0XEFWpe5EB
gSBieaAXG/KRsNO5/+HzpUNozVwfHz7mabBPDNJKvzl8mvPFFyZ+kWOo5syoyTUX
gJJVo+Ba5DWphoJkxx/eGiobJ87XV8A7ZvvRlxSqTAmBWh4nDLCs3Dg3rlCAoX0L
RrECuOsq8anOkr+KEfRlcy167R+YSbIqamljlk4XxJzErpNN3ybHFatBqDHqnQpF
XsCU5b9h9dLkYl+nAnoVmXYNAbEWfBqr2hXoKGYkeWZwUGDt8pnBfQLNxuI58sJs
oJjA6tF7mNtlGCi2PcT7T1TG02E8oTWG7GxgJuDt8hSLKM14hVaff/f1js6qMB2r
UcwR4/tFzAFFNl0n6lho1I+Y7L4Tv6jzoxfNTLFGm6sCLcueNhzYBNNpd4Mep/6s
dg6ZjZDC/0e0whJkJlh6nNdrQJqiLJKP5hnhKUhLVrW1b3NKczx52Dmv53Gr8Gh5
Sv5rWMBmbec6IpCxG7+6cIvthth5XvYQVvMIyRjcqSTetdLc+NavjD16W0I+uDim
b8BScg2LT0E+x4PX3PBEH1g0ZNOPMKmeSGuUvSgYuU2uu8aVYySY/UFnqwIu2Pwz
978P2jZIccs6/YERUO7x+Q+W+UTU3tvKdDcaCjv5kxrwm58qNBfaiT0HEB5yf2cQ
ynirIxpDdxP0uLlQpCF7yE4i9EonqVWqUMr7bt3r2jvQRrw5mxuhOllLqVsrZzyq
kMF0CgLXaewrJ2HGtPNB/YSpJHvnQmzFuwNMq97Q3DHFSMJBW8OcVAzSLeJhdHen
PKN0MkCW94imorVks4oz6N+NIbJ/k/vWt96UZ1/svM/3kAq8KUT80xMfzdOT2gSp
YGvuptxUPurSbPZ8iqKcOUuiL0A38IcYHjT936gJej5RJ6cuKL1WR3mZYUk0Hraw
VaqTgIh1sCKiIcGfBmRHh3H9Byk3YJDlFVvMYoHwQuH7TosBk7JUpSMCdlF/1iPH
OvycIGP3+JH+RDxPl17LWR158J+W7+i7ImOyFy0VNYNO3ki2DnRneyBsUt2nZREX
twDvmJCIKa+1wpsANfM6MB9rNdnbaMKwRvxQIjqhZXkZdwf5zHAAtnQq+KFg30Hh
5X+4CJ4I72a2XV0LYrkVWYt/wEDMbj/WEevcEfY52LjMqtmp/yaSK5suWEHDcUgP
xzQMVqIAF/AzlkF1CvcZaoWd20Hiygkgb2L2rjEvjHJtdxGuEDD0nUg2Dw9kyOI8
cX7XqrrAutagvDBUG587yNMJVmP8zfvGI60YlWH1hV3KTlP+CXxU1YbOPeYOCMTF
iKgxvZQ4MgM1D2CUfjK4O93oKHWLXuzwjPWNGIJasQxpqMTPLik6iCcHRZ9XtAch
tDjggSYPDnnGOOOsjIFirkbF+6FSSza8dSLXLGcShXcv2998JJbxZsV1gabYajgG
8CgRHwTrq1WThenCBqIoMtttgGyvhvBfovn5LtAOFWh78Et6ncCjF8/uUjIvslFn
qv1Kymz19M1mhedmB8y9DuPQZK1wZz/2oXdEPr7Smgmlx7HEF2qbr2t71fsic3K9
AjNKHAAL4W5BTnsFJeIMKc6Gsw0ikWYH9AzMbDkykky5XlnNojt9ypwv5xqZZYNN
MaBSXLURiuNwLQytK8BPd1iQbPbnfL3Ujs8GmM169SdthveY+2GwIKz8Ty9V7IoS
U7ovdrUpbaL6g24KlPjoNZWQ2otAuL6L83fdM6gDPEfTVEBjJnXeipImsSwvcd0U
nlFEw/XOOmmorsiFPAuCtrj+Oq0qm2Ozozwya73JfuvwNCbA0m9EfqGKAj93eYYg
p6H3FWpHUlR2Q5abtsDTNIHuIBu07puSknItZjbLqASbv3zOIq/Fy4QCDSJIDY1M
0u07x4zJgJQsmMT7q/Ymx/4vymGXGNXwpDOiQj4POnRsePJMrw0WLKgHbh0PyPKf
5mLuVb81xM94TTsk0oxVtUsSoD98Ez8kMahOanZQvyWvjh5soaZUiNSMfx1T9sIe
0KF+1AM7lI9WD1HKghuap1Kv94B6lnHKi6jRt+1bmbTN2Rh2UitGY0zA7DADIYmT
Bnozo4lu4MvuhcCTTO+NAi6LS6wAWjA07cWVMgxqKmMbwy4Dvi3PkiI6RWgba/un
ew67vmUIhLwHd7s4W+Bked0QtMmO3LULkjOMxryBNf0xqIyV5RoF4oyFgOoe10Cg
Pbx7sl69QBBzdC4cnh47dwBdiQO+wZ2NY4Wx/+QFayXwK4tu1uNV2TUDhra3oYvW
2Lm6nV97o9I+b5/acCjfTp6JlFfagApHDT/gu8OUpl9TYr9lW9uUKWCBmrcaYqkB
0lv8Fz/+YmpOIrk67SKagcB0E3bUWpbnGGy9l4BRzvzyapA6d54PaP/qwQa0DY5/
bKhOc1IH8L8YgHdFIAA1/5P8AUjCCPhVK+LX10nMzNx9qY1awnEvedtg9DE0VRuG
fnYx3rCDYPuuWUhRLV8lCr3d/PgMy3EErAqWxlYliGSCYlLQozyZWQwDU36wEjMi
4u62LXia9BXAkHo+KisYMtqdaCEvt8xptIJjInF4xEihb+zA661r6VqauWz9d1at
nIB0YZHu3sjgflqp262XtxFnyP/HaEFcEgZisH6pBpJ67MEgr+ZoH2gihZ4ktuol
FcL99YLVCxvJzwEeWrs2vwfVz04swNbPtBmByf5m925L7yMw3HDYWbOFLgh1QFf+
O0bvtLBg2Q7vSTtGxd67oj9iwvJ+zitzun+0ZLE4PPDhBYaSVFbCXJUB3//qHpUg
Pg8Pw6El5QL+ojjHjKuHclnT7TLXkUXSiQzvikW/MOxkTQ4hceApaUiQi1CwqpKQ
xXxKa5SZqXBstKBNXPFwVw/QPlzgMV9QT/bGWIwDG3//N8gj29p6R1imbjCBArE5
IkLc/0G3tAN7USlhyn0P8Urg1QIaGYtKHPAFttj9hOGk1m0vcIjIQg+BdFfBK3Xu
+ab6s84CFhaNudC+hCJmOpmRjL0rGQhdZV/r96VdgALJIjYIUhDnXbuGm7FYtc3U
hITu9FR/T1mYXoQe4n5I06WvGSTr91z4p1H6IlnPqKYT1o2nHyD9cwPkJbPGioeI
1Tx4xtVTccjdy8UNemunndOJ8PCYCnsl8AxN20OGrPwanywuPJ0refKcYOAb3zv+
kEXFVnLCvgWKinvWsdtoXf8ywM/q/+NpLpnfXfKpsSefSo/5wdYybmLjkClUmPeQ
PW4SkTgyg3N/D00TrggOa5HDnqNYGMKPOLYYEaa8aSHNaXWfaPQnRHpFlaw2ebdi
xD/FNmDo6Cf0V0lftqOU8bEvTPfQwhrCfqrUEjEwYoF/rOpiUDdqfakq47EBTQeo
MkCBenAsPYXy9Bz5dQekpmj/Tik12CUNjLxfiO2inYligPioaP9QeCmiCUiEU1Bt
LqIIQJ17I4mAQL3+X3035nUmxBtLWKLkFISA5c3yCmUE6UYPDla8gNgLsrHcrVut
4cdlwSMA/78haxMzBREadhdAkdBiMfiNunuDssa3qD+XQe3KwTPr3LGivV/5WSrj
Ec9ETh7GVcy0a8jGcHeeJikvG/uy24EX2JBNG0IiMiV65IEQqWY9uv0xWK1/KyaN
8PiTmDRNMGbDjIk8RF/6cPyB5k5b6hfuTimiTW0CQQ+fosA1gdPwOkde6zfqdOXD
u9xkLhMKvhYU/rDhkfmFsXSnlhcl0ZhkdyjvXxN7Wd3DQ7zN3R5Fvv20ANM4+2yg
0So7Wk4pTwWRmWK12/e/ccg7konn18dqsJdRIL5l33PGmjq6XgHGdFTUucrHhCz0
jrtTbUTBsy59PNBu8Y3rq0ecue0R3vzSS238mb0e50A8bczKN6v09u7W5jWC62Fb
b2FeyGjk/lOFJnJpMHGJLZYFV2TfuciioA2YmpOsiWtjNgeedbmUAQ5tAnkKPXeK
8FFXsjR1bf0ZVJjmKO1PPrvbU1E3GwnZ8B2mYiMzyi6TJvX6HnkU2dCr+sI6xWS7
SimbwO/IovNoOxkR274OqmnmAnr8wtd+NffyMIBtWLQ8A+jVj62QvJ83Xy1wS+vp
mjplBms+5+aWpwjFNWYJmyr1MtgMeE8f2qRHQG+WCm9PJV56ZQ1bsN8CnMzesv6J
FFUT737jEmhG7SZ+Km9mUFL/BwYTJj2uz6KY0nfHfTBwIUJPv5lS5RdUJoL/W3Jf
6EXmJirBJiceOCB2hNx8zvgP97yENGVVcALI+M8bziEMBxtFG0MQCbx25fV1OV3B
uEsf9XNUjSQA9T/fD1jVtPgsxaxXKFUZaws8dOMLlUdlxE3atHpyKVGXMHOWGXOp
tZIvGEpu5M/XIYyN/CBQdJN3042ieoCiwOok6LhvLo9UU4fSN1K8SKFJju7cf50Q
Cxi3uJa2z3gwp8zs8XqRU1etMG3rrADPIL+3TeEMqwz76doETUEpYtplEXp6eke3
z8teG9LyyiEmVqGV4E+0eVKvNTy3mCZn1r+LHyFRaq119zHfI5sBfcbgXIl6auJ0
oFsOJWsb9cX0Io6OFf+VBO9vgzXY3DP/IRwCQfcYisgySaqbswrbwDZNxkOqpPQe
ohTNF1a8All0MU4MBLnK0GY4q3NvNWPgmjX4OqpswXv/3pp40fCcb8zHTwgwUhMk
/URKP6v+7dyjmzBflG3wKinDNywSOXqIutavEXCMSP6M476Fkxb9MXH3Eo+MqPSF
AfV6fa5I/+D4Pw1Bj4V3UkBXSC2bzjWG0nzGCBXUdKoYjWM26F5uz21F2dCMc4qL
RkU9zDA2TQ1n1G6VQGntH1kfvwp1QBmni4Tq7pdim7G+q+d9oxXhMZ5pDKy/zZ2z
mWlamNySECnANjg4pbbiHc/XTnmYxmh8rFDEmR4OWl1R57BEJT2Uxd/ABPGVgajO
40nzU5UUviuPR2RLLEQ+mLcUQ7XiH7aHwPYzFeyzGw8ZQFyPTTeTC097mPOeZBt/
9LESJuJlsWaxCng1INf21fHuhY3345wYzRnYTdyd3e0LmmWHbjvWocTkWVf8oPT6
6aY3paxH3b77MqWRrnqXnaC3geMfT0tFTcgNw+PGZq9J0YLRJJ0b/1nn4Poj1KTD
tpr74PQ/l3PyoXAAQeuYrAfRoslY1QZQUe3xPU+7lUw1ZM3zed4H0jtyTlvhl9bs
BcHhlkpnpT7XQKcTbOmbktIki5SStCfwNOXm0uL54VgqvRmGn3NgDAHLDjgonlwV
R40dxaKtdnVh8W3u19CETLLxEoYe7B/x//MBBT2vSyePtDs5R2OEmUsPl3ocgLOs
bZ7wIwEb3EkWzNZe/a8jZ9IzzujA3ud5bJ8eHLuQq7yXHmv6t2YoWAoJWe+KTRmD
S/hg9a59ZnFnc0kUOZc0iYpgLnfurhBm5OE29iLwV9vyjDQfSXjaZ+u7HISXNqmb
rnomrN8WjbTITM9fE+zHYpVLK6dpLMApEg3XMWYl9oeJgx8DmspMn/f/yOu17Vk6
QYR9X/BQoAYswzaVJmKkYBXUwLg2gSv+QZXJa9yObac7x8iRoFH+CITW4ijzo1ni
YXXnXSevvVH5oL7eZm3jDdQnQ4A7n+cG2ew/QfgIeDlm3Z7Ga8XTsOC5gYeFv0Oq
qIXgOv9PSwzInx6LBRjvCHUjBcrNGOZXFtPhO/ac1wrs96ygAWMans5M6hKnRjDb
rZ7PHpbIQKxpiotrweA09fd0tIknny7tAQsFsV9e98b24lpIWctT2IMllm5dWKxc
5U8JZYx4fYe0d6lz0+IIuVd/c1SOA86JbGS1JUV5nXWHrYmshvnSPwRx1ax4FY6W
vCND8btK5klN+Vuht/qLPpsV93V7AbXQ4y8jPbwhRQ9zN6iQrgUVzAzvr4mPEV/A
2xbBRg8ePUJwTwNEADiYfFzomvrOJObYwCJVyKjNRkfhjtkHthIw2AYiPz03X2kK
h+pt767R7iavf8XtGmfCXNW6idq32yJK9NSXYBeGGCPQRxFkIdCaxJQeFSoau9Ez
iUsEkKmbBOGY34VWG7UfJBtE9KRp0nRkVIMhHfKwONqKV39OB6Ykw0aDI3gjJzbX
JlPB5iHy7gnZHoASt8nSYcBfziDUFfkifJYsqn+hqHMsWk0CuHFlzZWyz/IeEsVj
JZ8SWgkq/LAoYmpAOGt4eUzVGxJDYSwpLSnQWK0eFbO89TX3QUYq0XSP5UdDFIwz
o3rrdVHTkQX4ZFZUXILL9tjDvpkbnMyOr2brzNGbfMybImKwfu8BzefcwbnB9zf1
bvyqeq4WGVlLT7RAvv6VpzirADm/blfd/bgy8Dc/brFMQpld4Adc7qO5fA3Sx1fE
uz2Myb5I3mqlYEvN9nAxBOwWVL7zh7XVTDobyZZvNEa03XTYTYVwsI6FU0SappFe
3XpN3Aqolj4/nG+imka+rJIXyJu7Q5bphx0yHpief723iH4BjDDdZ/P+zweGuS75
XX8hvwuSI7wjgaNEiepotJbfiCmeoyGen9iZqKi5G2EXKsF1PMYIe1TZjeT22k0G
GyTVfxd5Yf5vIS3va9zo3D2nltbMYFJ+0vJdFeBYvchz/sVD3M0xhJh78tSTgnPe
lnuLqEBwpQz1GfaroCo53KZVyYAmmaeMDpIbeQwatrA9hf1Q6QbhubK26RKrNp3F
5B5LyMGq1Jf6tQjb8EOraw4HsLVMq1S0JDfxmC4GoymZAxFtkr9mEr07WfLNMDns
+IvEUF6e1bFCbfGYIcXOJ1mdtxISoAgk6eVkVPljA4DsIxupL4eJi2STg29xb8st
0WKUj+d48L4RhoIhOz3m3nt7o4lgWdmPHQZFzjk+E73wsJ6d4c8mtBMNzmoAMg2l
73qm6vovkLsJGE6QI+whBidyt2lAR1y2+AvqE/Kwv2rNJj3Rdzif6VdfG2vDQw3K
HmiCSQiCI3gzSlyUOal23uylKMAD8u4UrYJyiVFIB7wLr9nUpgkVQUmTVbAqyT3Z
UjidueDGKSdbotdMzJ6yWaC7PRfJzOLYvsHjAuyWxenuUNPdHrCPVWCNmr6fZhdy
51123sVb9FCailBPsUzS5pbT7//BZufCjlAtiPnVJ43GsqQkgjchuOvQo0OBZ5JK
dRnaFcZYyh3QIBvAYZVKoXzdsF2jNMtdNLFUxahyDpfPZoezgsLwc7NTwVeX07oh
UxDjWkiAgO/4N69Qq/s4YjeqwToOvz9ZXq6yjJRC0Vyktb/xihulSHct5qhpEaDF
skgAiEGG2fbWOwx3FoF7haQ+r/GgACtFRY92CQxYqc8j4YORTS9tjaOVM1dOtYL7
a7DQnDBeoku+5KEERLFy96pHiFWhhgPv7MCy7IFLI6KNJZMtGpNXo7v8JO2bv6Fx
zxnzzwsQjNqZ7Imy40OUizw0VQfv+NHoP23VYb7b4rYklScrIiXVisgElkt5p8kJ
kkFMEbLV2NgcZhq6o1p8wonHKXd5/miSWm3FGmsSNz8UkDehJTKwALRfI4fK/Jk2
a8DR96XvJhTVlz4hkbrGf/QaIQgfLwF5ncpSvpP+4N74yTlmI4bXbK2DEulSgkYw
bLAs/T5wYl3m0laxudkFWTftaL+KpqVjgro7B5VvJ2ZadISE4SHfo6TXrdKG/ZHb
4dNfT6jYql0eAk5GsnhESYBLFmO8ixwYTtRfmTNzWCJEPgvZd5bB1m9LFH2EPO6a
nPiyXk4C49bkwi5r7NWJR8/PhxMovbtr0KhTDNtsgSVN/iiTv2kEN9NjHMNMVcjx
DpZLjr3EGJM9IE+Ab6bHHcIprEXm81mKGRC1wxed3WocvEUecbUli1dIEAr4OorL
CeS+oWtylfr1Fkbq5KXwKG/4t+V0z+rG0A5XgwdqGU3XO1Pbj0NWTNyj/+yVFgU1
IRBN/GEsQjNDvYK/ozM+r6Vne2OK9eBcQRayJ0YjN0xEarBLaG+YSKCiDlJTBNMZ
Uzo6kdwSplCdtnGytlF5VK7fzgA4McGMUFY6YdphXEbRq2dlDy85VhtooG1iwoKR
TI93v4ctWRLoH++1Gm3mG6V9n/vmEnFJGb9bPIP+90fCfcXrrqZtAbN4HVse62tT
1Qe83tTpBQPkCCvolqkjOW0DiEY4fTpa4KLVtVBi5He3S3Q+N91szN/QGUrwJRtk
Mtl8WU4nuol0ghEF4bCkJe3kTuexrpb62CJcN4wxP6lYSAKNGnR66PmMJTkUIYW8
cNoHRwBTvTW9KNA6wFzzzIAqnVDs8wFy1Uajm6dgYoX+q2+JpvjTPXG/ucP9eR05
J+ndDTyceQSP04yRRU+ErZxn0aLvrQeS3vu/XgNMZz1lVMu3cw38NQqNieM+DBAn
HUWpFG2hiDAFW9fKcDnn5KDx0S4vM7Krs6exA/6c5HcFkSaw7HVxsmg05ztTv9cH
zTWiPuxghf9DPRGkO34ypt03yp6bvwXOKtcHyxduYtJvEUgasfhOU80gcCE4TpCt
xQcf4daHtx1eAcxM0VFpNpsYYecv53EdrFd1qQPPOxgQQ2ATqXA9vBd0gpC+7iqy
pPavZEtMIBvVlEYhGTMYmVysGejiBMzJrEgdNdr6eeld1OhHDEhhe3xIHvu1QHcj
kI2mTYOdd0+/iuwSQijvbiVkv/KNikw3JGb/yI2rjSxOVLQkHpufH+npYrMbFP1q
nxWnFW4ThS5u5krqDykhR+lnYMx/bSLIT8xAcX4DdZSMsOmPLGsbgUovlBxiHwvz
q0nToPE6r7vdfjuk+UY6/1mGYgSyksdU10DdJUOxCsGwTUAOdraCpoBPa1e9Pn6y
nM8zdUYBOzATl53dS2xua8GQOe63VFMgxBT2oA+cBo1NrGBaShaA0iFtcA6imQPJ
qIvUoA+FGHVtfNtNL2LtjhcNgOVmm1TRIjvwWwT0RyqmRInpaJz3EHvD6GepJQMF
W0DfCf4ZNCfVhqE/kVgUmix5rfwtOeQTU5jICvE6Td6ElUDzMn1tRO/y3ueLJ9oh
9wQIOdMFbneSAeQYaQYRCejbDPMzo9k+AbTJ6QLoIwbzzG8NsCgPeaX2biflj1ts
2+eVWQGNr5ckIZ5ATeK0NWT68IQ9QC6ZwFyQFPo4xsDNiV/HGeGLAmhQdLv+vPKY
uUqFDySoXUgAP51IdCZLi93pXaApgv9D1tbee472ukSKNo6kVtNit3Q4x0OaRNEj
kXCZwe6/A97JaxbxNX4+/38VVkZ1VjFwPoa1fhaKbUMgrkVbLcH/WuPrmwk8D1KF
TyX2Sc+zTEExXq0Z0qwqtWxyka51u8O8XkcVv5noC2uMPC8rmcXLSpkG2IKAW4Ak
ApCCGE5gVqgdf87g/LNog2AuPnS1SO+J1xGuyujdmxLUpMAxpzdLv8mVXvpyjxGV
VhXCxX+vr+I5av4h9ExPcqB52p/FSwejHaZNr751bfiQv+QGaUoaKlQhnhQvW9ue
3P0LoiWJjzFL8QzjVELr5urNwiGE+HzkV3O5rggli8fKFQvhc9U12w+Wr3P27l+X
EK6Hn8NGnYcWdgg9W2q3s4k1pGN3g8ACE4dpwJhCwbk6rGkyo6dGePGqqlY2Uifq
7ZGw1TiAXGQSyw0XEshicSnq3i463TIE00LSBVR94FCmjsEqOjACMMRMypQfMt6e
PII6WNSbUCrKulsJQIcZuqf6XzKVLqvD8DEdfI0N+SXDF6Y2QykUeUkbL/cPwJMy
NX9AhKPsEdiQIgEfGCdilNqx+OEnCeBnQZ1Erlh4uSufoMOlOfsqxVMYApboqnfL
oKc34KenV6UkU6kayjdhzdBHrQErI4ehy21PilkfnpNEoEJAIvaC1EdjYq+0TU46
5wZ0BCfx5GnyGzdX/+QRukoeUm4Rsx0C1NMLRAzMSTjiolKMyE1g56GUIkkiiA2D
xw8ZYrNoB2zR8o9JA08crVJkg57zaUDhxsmJaAOnrizv3APNKotDh0D1v38h6df1
u6WYc5pwI8s1Zcxh7EH9E2g9Nuf6virEqz/vM8YHucUHoO3u1kuWd/7E/PoZRETD
HQG0S7Dw3FMpx4kzmW4TDM5DfudMimL992bGH8gF2PEGENH5os2cmGn8bVdLIdda
nfUf/wHKOCUUzqbD3o75PYp+1E43swc6BXiER5/7degIQvjt+O/tdqBXsCJHg1mz
0TQkB9zeD2g7Qc+Gs/TsXKoKv3ZwKvYu1NxhC/DEHlobcrkeFxn0RyT2RlmBtBaa
syPWTV0cAxc0ZpVlQnANBWtqL63Zq86jM/iawyGSwIIWcvJljsanRMp5TGk1+R6k
ovpVAJcaWk+DSq+xe5JObQjXIgs6yiUh3AGhmFWH7kzW2Z8OvWk2gNbR8D9QNp/2
4FGG4nPXbtyZDQuZeb3DatFvpi28Ip5vNyfUS5E3F4gpHTha5wutM5qdCaJ5pHFv
qpKeSqtc4bF5z+GZtZPF35WHgrzQO4jxCBZ8FfIv8KXawQzZBdXV16XPexbTiWRR
KSOy1vagkGeqgFsAq2HjhB5/41O06Yp2uDT2JO1G6PK9IO1RiOKYBsU/vO9QRQ+G
4Cba1JAM9LmQI9NRPqruRQcI63gJtMggaawQDhHZo9r9CRefODsJS8EY73bfdsuu
vTl82EQPdbc329IxaJ48Huq9nC7hXDG01AzWAfKXixv8MOGt4JnbDmYW4MUt8PyM
CWAIrgEvJPZMAw5eeH0FJ15FB/ny21hN0SvfLkS8fAtST+6DYMUiliNTaNE49DX2
eFpZ/b2n5mfEE3LoVNMvwtTCJ4HWiEvODLlB6IGLPbr9syghXQQlHjl3+NP8UvM1
w4tJa1UEEjKnLpr6tEN2pKVy1IiZJacjylWy0ckx0UZUp1Ol9U9kMYhBysEuGOnQ
oI/YuPZrw/h21j0+On3dUuDapXQkfZEqajofwl4SB6sbxYNlMQlwrNncPygzhyRj
RpzBkD0XQx+5p11rCFJkwHqoLqxJtvUcB7K1v0n1sDfvlS+noLHOuWQbFyCOTXce
3lVTErHHpOPN0GHy2u7/jLYuEQqblNVU3Y3m9eHjBflmebWWa0aA0bSX2VBOIr8E
ukb2i/jNggDY5ZfWtmnQlX9TZ0/njaEO61ZUQZRE1xulQt0/0GtCIkeiKuzEhMPj
vpw1BPF9R3BmaFFxAODvkKqiXZnlkIDLNLDg81TC2BI5RKhJ9DOYZ6lO/RMR40rL
kjr/6MhVKfSN75jCj/VmN3OuGR0GGgcHlytTYXE0YByA0b0o6PCBVTvLMRVkp1oU
7ilguSCpr6Gv+zzWklTR8dmmELj9ZOV1G5nZL4uXFveHNpj6clf5yasnAHeVYqJ4
dyTrLRnaMlBPATk0YwdtubWDOpK7+3hzISjS2F8g0W/hIsEBaLR6rAA9+9c1A8Ls
SuR1jFiACrP0uxeQQF2wuuvOo8klS7Qtod7eC1C8yLoQGZXC62j+zAUCP2bMlWnX
Y5bqR7bf3VrT15yCQMq6rHUd5ITq5kUfgbQu8lJZPHKV0BlFGMjBm7j7A+Zj2kEG
R6qwxbdsSWQrT9gAJzqMRjhzpP08X5h/knVuilTnkPOZX9Ialbi1RQ7oVoRN3iRP
VDe4vEbxZsSb9D27uWi1OFSwpXa+of9r4y60ttbyJMl7NayOeqxKGJTVZp1JYQ2K
ZTR/BNWep8MPw8V02AHT95DRSYI0oa1NVt1oNuzOAV0elM4/R44OMnoOw93seS35
vLt36t9boymVd+Dqx3eUPfRSYjeXW2t/Yg9cdisO+LN7unCM2yDfOwoOsyEK5X6R
fgvSdJNU7c0sB2q9ktGCJ3/K26V9LQx1gS2N4Un05ErLHkisoho2/v3jDFSabnHe
LIVE3X/7RQzPA/BdLXQqo6dCn7jwwVjCIl3LONCBtoJaspb1QwSJos3dS9ZskJeQ
FaWyF2qdY2qef0lk/hYLN/SrtSSyu3f14LPQm3UAgOylMmyjlPgWR9CsH6uK0AuT
830/ZjBz1Q7z0DvC+Nbp5HqmyLrzN0UrUroTFv984HWBWduc4ZoOMd6Wf5TEHAth
b/ClIch3I3HFmjJMps2K6cdkdjByia0/FZJVoegZPfcW7KOE7az6A7gwGh3mtziw
vOK8l7PAdMBAE9PKlFCePttX69cpKjmGQwMHQ/ojMwHmovorr7FvPtgbrZoymbhl
vq+E7d6NafFiGZpEu7syYdP7mWiMd5+oNv4GeAEVf5eo4HfZ+2PhiS9taB3VZatu
F2vva1DIYFnmHOYuUCq4hHhCLf+miEE9L2TvdaOQgCFiBbJwMuJM4/GMJ9bkUVzW
YtEd6Y3xk1pNYKMcNoVOSXaIHjaadkknGNPAJHeUhxIgD9cTUIW3kXSpJVdYdois
tI5kpMceJE39S9KHyBVBAfYUELPF4wB00ftrdIqU4yNd6Q1tQQEulgnj+bIKWTF4
WGbs00PW38ueqODkMaNUiFsvXDfE48jgN3Bx098MP3HgQBwr+y67v3baMJdbJ7Dy
SgL6EBE0c+L9hAXLc0Blce3UmOfIT9DEiHtI2xxFLb8Tta0zNf1OrOylK6pxKy1I
C4zqcHPQWicdlK7t6LioQi5RlHh3Yombw/pYRlvwQ7H9od7XJFnr3cGJOi4d1lJD
BYI5wuNaGjVkflmZWB0FX0ZUv2bmdxgB4UH5fan5j9T9eeHsdy2dH4ASc0mbF8en
qeVWoqTjHuVaB6D8+vuUKVP7pSyCvgUhiguRTpZI64qRiWYPBcXRr4ejc4QXFH+d
u/DMQcorGZ2gIZUseoHx1B6Q/gtkxuibrdZeMpmi8CYgGfh7/LVto/wYbSy9Tslz
dZ6BmuzCrNiolKvL6ixJ1OCs3wHmK89L/nsZjHs171Bqw/MGjqsP6BS4rcLJw6aH
hb/TgIEw6cQIPg+qZvU7fE9FgztZ4DWB4epQLVsChb36HURYMmJ73FFqy21Ucvoh
e1/ORUjeo9ngXETRLSBA+8/9ggGRbNTa3OCXfazti3GX31DeUkojA6Fk2Xdj2tu5
rR4H2xq2dAm5LmGg+XqZCnLloCCrUi58milA9erxi1znvKdpM6ElatJejwKyatuD
k2MRei9bD52XQ4zlYNXZ5mhV4Z+gPdrA39AcGQo1uvIHWmcV1qBpSUA5FEBfi98A
kx8iGMau1zQK/he9XM6SmotvifIZRKl6vba8f17wwzwaltSZLILWlew0+3aIO0zH
D089GGqeS0Gl1uxtww+/5Gn2yjqZXGs98NosrCqvwefypfdRTq0H3BM2HSQC0heE
EzjDbAGykz9XjemPMU/GkAgZxBqfZ+1nm+cEg5rmRAQ95Yje4Qq8Bz+tCa7H2lAW
TtokwkIodGUZKbhcnLzWmcNKCmmZAoyygzjMhJtjHVHXfqz2OsLomjm0NkHrgdOE
cB/LFffSIdxjf8i7dZm70oLTgnwwZzO5sxZfmr+H6UeHEt67i13JXHAVN8H5qhH9
82hxtQNDMqTxn4o8WzZcUr4tSGw075XELocPuC5cO+8qxUmtDy/FEBGx00YDXIUa
XsThpoExl4TCnwGRAjUD14KZANmO9RwRJpE4w+RXlGOhZJFRAqlsyBmmCoDj8D6y
ELMyJsa0ZkEONT7+CLe+LbUzXDlgMj8zX7XhMqNMwq16rlhSfpk8YhH42nMNr8Vo
mZcI0eEClDy/4zkvvx7dl5LAgPCPzN+i52g2IVhn6yewYWbkRZpaRue6A9W8BbHG
kAcVWonRQll8795NDj6pwGEXBknB/cIfbFqKfiUtB9ZromWhHJ4KPb9x43xsXLM7
b8ZOHFQvMWf/3qJzYdK+GLDy6cqiaLzIipAsrUa+EK/jOUWoJuuy94NyB5ezUcgI
+daaHdeSUyEFhOCF3Qbr3F3S+nqCNu5+2LNDmTxiJum2lmufnCqVMsb/PQAHj5MP
bH14Q///zcVPCTtBoKQA3GXjaFvX89Tr3mzPAi9hMDWki9iBwls2juuNozcJoxlx
5Kb+uhKVi0PvTY8O+a0jaA5w9VEfRFJmtj+p5W9CrkVI35g01w5aO6T6PX+fEhWw
nZ5gujL/lBbsK9eLy13r5PYOKxJxz5z+oUEESAMEoB+wXr05Y/t6a9hdHP29xwdj
1upWn9kUmoFFOCNqWegxPJrbNjzLC2EiLEbQDUIjeq2f/43uHe3pKBfy9Erwg7BZ
e/mMbxASjxAfldbzxrb3PWXQFvQhTIWzja2n09VAP8LiXmoknwJSZBkIysMM/bc4
SYLCpXRZ6MIFhog8qzWLnDxG3+d3IUhT5SlMNUJcDItTrLjq3Hkt/6SswdVt0OF8
NWlzR522PrvKcGV9Jqe/Tf8chUFwPiXhk4FS2jaE+3wqMT/hVWjHnSIyW0VxiinV
dbCOI3B4EnEvivJEyEvorJw/cVCK82275ZyVUV/CXUrUzBzTDjoXEho8cRNoI2Ac
SPwNCf0Wk+XV9m91Pyi4Fxvvgt5R6xf/ntWNV6C64vrg1+xG75XDxflqt+DHQIrj
NWwau4h8JtbEQV9nUaq+iXd/ugkBTnk4gobeL/nBC1rAZ36DLQZzTLqu7V7EKfPG
IRKHuBAKejavMkNU8seSaKJzK8zH0kDEMx3Xj6wBWcbXPH34iHiu2OntqJezoIOq
1rvOmwU2qT4tI4OLfcPAVlg6waRteypkAOowscGRZcMzFXEhXm/EbGt5V4A8t2rL
x891XpXwK1IwkYVJTKXvdZlLXne940VP9Krg1K/obNU2Whk5yjOw4sJGPG+LkfdR
KkfoENQe98K8Y+rkOqUI0fvJupXTbS6ZWrj+KWc7oudTxPVhH1keUbTfdp7dOLIB
bIZXmq/D6WGjONduh+DCrnqSUtIGOyhudiDU9snR/Gbf/hFhg0KGsjOf/pMl7WRG
GpraLbVP40cYdBZFBgM5jl/gGdoZYGYvWH8RtXuEQ9R7GC/usB2HiV5XJISB63E+
Flhd0fvs+ZJtKn63gp06wLex8zK2KDgvO8EUqt6OzqhVJsNiympYyhG3qKWdYIgR
PxA1MRSMlkmj+1omgfW6/VKAt+AJZmnUHJc29mYh7te/00qOLnGD0ImlfVQT8G4Q
m9GCVBedN9QqYmOo026fRvimiGRt4iS0a59BnOEuG3TcEI5bWZfhUeF9dv94crnI
vnuAIVV67gIyazbpO+vihWp3MIwXl0c0OkwG8TPBOZqKMknFs51iZRy2FcKjIgHA
WMF92KI4OLTqLTvHIlFfNuInnoSekLml0h3qeldFihBuXER+9VOPaTjCTNpCWQlJ
efZgQEfM8y/UerSivuxulIeDXkA99WMZ+Hc8cjMiuCLARXt4T1FytQByd1B4gcxS
2BsX51ajflqlPQmkAPDrd3fIMGJFQKHCfhHcKzzu7H5Jr3rggj4Tudk6VCxs0HAA
r7k0saHy4CPorLrx5bp3EfIbWf2T2CnBC2IRij7pwsvMuWYiFrSxSO6ZveixrgWL
6EIR/etFpr/dME02gJpPXaQ7o92qytBLJeXRt8AH7LQkKV1aCYr+i/9ICo5gdXSF
Gzwv9YWIKipqK8RLAsZYkcN1dqDJ39HPnGdEjPuZc6FcjpeJSSBhr87toC6yROBp
/ghD4o/ndVdGWmTGGl+lxTo13hXczGR7MWRwsl/t6FrjuOB5f05wES1B48vw8du9
ITQE+V/WumE+hjhECx5FGqp4Nysp/sVHW5ftmp7u+pkpPVLGuxMkB7oZYwGF8G7r
5EMfKlSJCiAlybX2wl8bX2F4jsYkcRsLv9t/W3cXLx+H7Rdaobpg+N8YPdOOmfPO
u4pFdZ0v+t6vspGLVZE6XMPdJ7Yd3GFPRjWW2MLTFImtUxxRmpYZtrMnHL+oktEd
g6R73BHqH4S0hto17ld38wb+8xgnZ1KthA2qeqyRntTGbyn3Jl3dRYuukb+xlOsc
71ZhqoXw1UwODxnIsAwPhanjYsF60K3AVyGozUMC0w9iWsjaZ1jNE6R5QENDBEUY
NjXuUbS5xlu9nBQ7B6mzb66/F0SEZND3/9OIqO6/VXeB/iof845mfkNNq8l5tcd+
icxHftwgSF/IGzDZimdEAg9eiWGfDVbw7uZMVFHmq3xKh7mQqQV1BvsJikjqwPwL
SUektT+j80GImN4bpTWc0qRsVFKVWRpXUkbzCZ94UH5tyPA7PKBCqBcbkdbbYfJQ
wPiGyrVpFrYivTUmqfgcv7JuAd55uwREArG+37CUPNhBRGDZHvRCpzdawoqJk9S/
eMRJ2s6VSAfs3xH6ObsnSgVL/Ho8U1Npy0rM94CF1Ieo4N/eq5B+D7P/OAMq0dTX
aPNLBheK5x7K1KEucyhQj1LrpaIepxC6hb839IZ39xwrlM4Hr8+jhV8fmeJX7xnp
9m8L3VJOlnTjRLFMVZr2INQCjPjmUd07kWiC4c3Qq2fSk/FIBewHFqdeq+DWy/Ez
FesJBqWe5CNMqYJiGtZJhnOPo3VisNqIac405qBPW3OsubCKBvFmW+MfWDkyZ+yH
d1iFUaupRli/fcG/VfRR6zrONmEXsSk7pQLT++ZcyfRFwDfxqo+PYAgB//BCez3K
AvTEMfp8se+SSnPorCF3g4KHNxtkdf9e4+yYBeZMLStU8n3E2xOla/bAAhUaalxf
Vsqi7gSe9x4i8IuP/gsfzUleAPsrlkuowJzH+lsir/VvdvzIYYnnz+69U/OYGBdi
ZmLL6yrpJaR30pePsXIP08HY5trEuO4/ROuNOHn8PRLcKyp4aT3ldz2Zj8ptXLD8
+DsiExVWnzKUWPk7/9tHTYJlJ4LzT4rtFLrlCh4SSQukKKryXsVIljPAaCx7wuTr
wafsq3PJSKYHxRj4uhkEgX3A2uBap2SePTcTkhFOqrlA9Coul88TN/yKKyWb/jHD
prm4uVtG3TyjpV5G71/cJAAGBUEeh5Al7rGObL2jqg1g68qTDFVRV3GQs2D1jVf5
I9+ihOQIifRb4PSb6BgQaVOOUQCevnuVY57MqkBJiXoZRT4jI/HZpSuVOJcNKLWC
i+4wJnZ+v3jnIF6R2nMmBbS6jatEL/9dxB4m3XnoB+3EXbQAA2qkdNuIWPSRjJq8
MSXMPzP1Ls4BmDvD5t4snujdPve86x6SbbjzCPS6GObOmkFGnl72j9+xi41WX4JI
bzSid44KhXDZzrQJnJkWx/NVqGjPybjaSlF29TECiqY4oyz6yupuNGLlZ/2ee7SJ
0CKoYz/QBdyyzg/gP+zU9T7gAnhGK8IpjnWkaKp8a7vSP3IvIpIs5JME0esx7g3Q
P5Vcen5vTvEnJB3h6I20KCaJ7MDlzZRUaXdBo8+JpQ42gOv8fnog4re4jvwHrprX
x9/Cl0SEgOQ6HkZpVbKBV42ytHFCsMR7Z8t3t08V2PVHVFj7QR6UP7d7L1CxWQ0h
22KbKe+io/HxgHkImC94XgVC18Bl+wqOegUr7KUVvG3KQ/fLOtKFUgCrVNzcLyTW
q6eFH1r8ET5rCDPdLmLUTFZcOJC3TOTMsYG7yuza8CybWSzAMATSRyjGaOvLb6/c
2n/WfJJflm+JkfPQ9gQZ0v3PRMfIhFYsMAHz/i6lDYlX7fpoiUUumz9AMCqawL7f
g3fU8fntF8/sZ5z2eZ/0RLba37Nseu6NOCelzhY26Oz+SzK92SODzJyOsGco90ae
oCLrtyfCkv75QJkSOGL3nT48C2nidgcICVJidZrtTKCZgxrUg+cMvJ35hq201AF0
sDbQWGEEpf36hR8sM2GzwJoeymaOU3ssdCJ88gubRr7nkfGwFZlZn5OfImPNkkG8
+NfSuOFyGto/8Ph86n2AvM+yz2zj6SJiijjvO5kuA0Xk/QczrlSdE5+ZK9dOAerX
6TuCSGEjus48dTg182VJ3pldfRxLJaE273bS1/pGO27HnPqMcYJf9sHGlhyqcQvb
`protect END_PROTECTED
