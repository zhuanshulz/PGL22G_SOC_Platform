`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/v9rxNVZColb/U+KecNRaTnuBsJvU5+YJAPj6m67jKStWg0i2/ze5s5wdOhhhQzY
tZUh5zBEDgYHwOVP0herxCfkrNsZpDqUPJmGpO67S2woSo59oLRwwl+NMkeIk9U3
vBKhY42FogDNoCJFBqZ4tftvTPPpXF/Y2a7fQQxBC1qCLi1vlD4kQUWErm+pg4mv
gSZVzXY250hwS2uhyJ3FkOwN0Af8ngSAzeM2Mdd7O7tD3Z7TCquIWLnDLCHVtlyz
x0NYQY2JggYG2WQULkX7bzvo0iS6zvVTiaUYrGy05UPPZjkzfHf1kSHQlCx4Kfct
LNZOzecu9ULENyhx4HUJaA==
`protect END_PROTECTED
