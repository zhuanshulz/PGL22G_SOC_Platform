`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GhTa6OBffHzfUsasRRpGJyJ6759s63ExToGut0RWjhi/ipri83+I56zNzVmv3TIL
OUDjhHBeu2TxEX6JndRYH9L8tBZTNjOWkmNwiWsWcUrcVhbVacONHqKDtZWhSmhL
hL17VypPBCW3gQCUHxSvvEUolB8HYkL0p3iRuDCS5KOycb2CUlALNnRHBbmdTixN
C672lwHkEvM8vkEQZ25eS4dQnt1JeJ5fwoTWn2gCkVG3g5B6gEKD6bHeVTWiZOKk
D9GGQaEdcRfrjK4qWeJSiaNBfreyZs4q8FftNI+4vJbVnetpUw6GIddTBu56QVs1
hiRjc9Ni2U9bBxciu0aGW8W2Gz4lRpW31u7iVi7L+ec7MTZJVy4uW8ptAKN3sa5Y
kPM0aEeYuslM8jkQRXDgyrj1fArzs9fH4aBwxinik7blHh5vdt4nvRJUT3eCjqMs
8/uwL2YkSARGuloRJ9KCeuOSnl/pzj7DIb3RTEyEBqwo2i1xZnhCMTO5SrFO1XCn
mju/VF8Sf08V0w02CJWiNSrUibaPKCcBxn8TgnT2PMIglbDlfcsBHYX+C8fy+u+X
6ZL9Sd1gGHLlRoB6dQK2tB/ofTnrCHIEWRAxTfLmUKKymRM2ydRllSYCW7B8dadV
l2ppY1TnV84LFYSjCBVt77fb+FNIwJemdZiuwA+4QWM+dZlmD3RRNXXByfSvuJM/
VRM/RgdVZTrOat8yZlMLOuI+X6phioIekh9h0LgK+/MpNMNOYvQnEANcmkQPT66Y
mjCDJtINdonh2qCPD9Druw==
`protect END_PROTECTED
