`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VE7gEZZogexeFFO2+lwB7tSVOt6YPFgC933w7X8xrTtbLb1KovDOdOt5xiapJOte
DD/dfIEbarfZW8RT75OSycfJgipVNw6jXt9b5b+5FAgU4PZpTONpJjsVNCV1dijs
aDZOtm6EHtAAh8KkBCKOHO+NeyRDg21AWzLhoK0tTjEBc/VU3v35cKDCAbgZdxT/
Jw9iyqN+XkhJ0pfvanhb+aDkIRp8fafiUCPOT4JQJoReUJJxgRT1wbK7d7HLQGuc
4ajEPjY20G11TMXWSp4LGjBGUDJlNBjlqr1YOY9qPb/+h60i6ib/g1yB7NLOFKpl
q+HjjAmdDuEZIRVwCzEfV8FQuTuQoiVCEO6DAZL23EYcQ5rKdRVXGC4btAj5rZoi
BRZIj8y+mA5TkIblfYgS6eI3FmcmaiSPxG1svX10tGViZPNhlR1YhR/zd3Oy5cnJ
gAjRItjslQp0WdBfurNbXCH70nXYmbH+ajab6RDFtzcnbqhhtSSntyDh9uRxYZdK
9FkJwKGtsCraGntRV0hHcA==
`protect END_PROTECTED
