`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zhEkeV3efPx72yaHzcFoqayJJ74TM3K3ZzSUIlNG8Iq1cn/YOEebf+jCw/yfOLg7
hjupe2mysaRfo17BWaOKWZJZ9yb7CWP8HWLdN5diluBRTnFox+kI6X1KPT/Zq5HY
me9SQTwjpYrxXZxwwYsmzObLikqWka1s7WyTMQjysymKBD57RGjJ3RW9atOiRGFN
M5l+8/82X3wlHTifneyFEeD1yfswtTO2Fkx3Pu4a4sCMEph05jXtaB0UcZamHj9P
EuFTDtl60TuX5rvAM/yngIAxXG8TLrdoz8WsAPtakg32x+NLwr02AiICd5m6D5la
yowvmwbXjDk9IQiazUiwyu1MAGbV4eoDX0KdSAVOlwXvompfN/IKJ2amq5mEjZZO
ptdVRjg6yVAJuQeKAhPsnmy2H7it83/L9rWU1dY2FiLy44TGIl1JSOtPdUooRe+e
XxqZg+Dpue+7g7VqKgDUWdGAcZqzxff2awn+6+dvf6zYVEC9Jz0LJeR2HOcrLxVT
mhlKftd50MqLAzPyQ0Vyq5fJzstCt5J2/0lQhynqWvQORGTrXJD+pugQsRqeCtLY
AkrliY3Qwm+D37ACHgdrt5gv4V9IqkAWo0FuJ3Y5CvChEpt+lUvECGPUBZq0CFMx
IwoOaogt02svBouzOUEFeOZa043HllkadHO8dXAde7d9BTPD4EfbeypHNmrpUX4t
JoKcsbO0WFu2rwCmXDM22OVQljT9vpUj/mdj8SInSLo45/OSXAgEDpCKuXBqVvws
ziMg0WZIeowH3U1ThRDNJxvPfSMPYZZTDrhUkQf5vWv1wjdEypVPZ0jF3/HAJwbp
S7SNJMBgZhJmeo31LoAY/SPuQFsrr7+DrM+8nvKxrzQAfjZUYmU0OSyWBq0BXY2o
txRZhBJJoCRYJpYn4m3D5tNAfiJYG5RPk8cgtQ09SZWYentKwmKnXhycZ1vLtaVI
QB4iIiEDwGirysZuYJmywDavXDlZaFaDebduLXlv01nnbnUzUG3trwa63ORvVvGE
jtIy08AsIfLmR1zMARdKuue8fASMUKLOoTwKLI2YTOts/dTjLcqEFI9Pd0cR/e69
4RWJq+Og9fqtYc8LVnXLBe+axNQCYjCT7f2VYwpr6MPKcKtDei680WdbzSzDHOWs
RePsvy/9cCunkNBjeKFmR0CuBGWHu9FVNQz7TOzvQ5vtq8fji3mbm7+D7+Bmy7le
A1kXs1rcebGJRnKJrpogKCRzi4P/0XNYGYxC5i3hE/VybgIcbp+2/sdfh064g1KP
YEP0i0xogsWytWVS82E8HZEPCZ9fQO6wq1hQvLbMKVZwEF80erTKOk+tVw82gRSr
5B7TNY2qSeC6LWcWrqa19dwNCrmdMOjtQfT467RxMyDCtCxV4N1oBZc6d9dHj02E
Lvg+TYTUpK6FEYLpwqH1LmpNKIRxg5Na5ok+XDQ02aIJV82TJ9ps+P6IH9Qesz14
GIdRKgb9ugsVxoZzMAcze7iRxAlIbvu+qBKH7J8pf67PSTHFCHU9SZY9A/USLnPa
LSqwMBAFIQuPKadNwCh0YcR23xXTAyFdK7EJaYYGWkBT/TcOSp/61CfNyF9JXLmt
iMRixSX/8JSH7kdjg4QOqDl0E/p/uNsH7PyXWK5RxM2MIW1rCR++xQ/wks0b2/Ow
327vXUhtwQq/TXNlHLJwChIGiF9NCa2V/cbEqExs5lvBGv8DRRXzlwf2i4sFJqwz
+NRAqjVoKO/W5Rm1SV3A7LFRs8skSAYpfMUTHV8AdFYARrOe7O1t1yOCXZcyT6tu
lV/NTDP1b9ASA58jlEQn8YRfYiYPVaXgLeT4qmo3/9wBU6X0d8Z1Iq38SYoNsMBW
rh2efkDfYCkijjgsQSrxe5rj55bEOPMRrUj6aaM9hsUaoz485RW9/dfpgWMyF8UQ
i7T7KPCqS2cYT0bFc//yFFInkgvuhMQNY0mDjMpYBfYdF48CoVug3jYAHWuAVpCz
yOAYRNvkccT9jyxMKPK5B5LXCg4bDd0z6I8J8JIXrvpCkqgEq9ounV0CG6iE4Ler
9yYo2Bkke/Az/aBroENsDKbBvDMdAR6bAAiiGpXO5Gr8tjSjLpTmEz1OMLynVEX/
j9XUSvj6iK//rrtUpMjrEYusPqGwe90aoq4c1BaeUAkoC5p4Ymk60oyX2TDXVin/
O1WvVwhxESKz7pO9r2sDCx0inE4mWHUFr3fEvNdGC1Drkg8As4cyM15I6nV6gUkj
/nRY3v6VdjPqx0I0AZwlH4Rz/9YQN87b7IffuxZM34RhzT7KQsIYEIjOITWn1irj
thIwbuqTQyJwntnKY+AHyTU2pjqHeZajQodRfM4yuBjsPb1z7O6w2w0ymIljtGKy
8+FCj4jlzxjEm4mnqDTTX8SGapDtEXCkLqy4nJH/Ah0p0CRfU5FG8wzmppCv2P1A
BiuiWw6TlreUVeXxK3xLx70LVEJUJPqpoKjTV9Vk574c60UIOUNATISTHSrcWsO+
MAWEWZk4IXD2QM6thqPzFsyl3FID6UXXLSp54O7p2PJP2rdyzqkjHY51RAC44vXI
RqIi//y3o6UQi5dOtSQa9aay+i/BqU3UWhEmJVNut0bG+f1wUcp+x9WVDHWaQgNU
SfEAAr23zVPAifnGqG02i9d7bTTJgayYg3Tj5Slcwxkbu/FJlTZymvxPICUXjqoz
dSnYm6hvJ6FUb+YgEV3Em9wOI3fEGUwBUMmrUPUJ7ezfV7vibq/ebwOIp4rfWq5j
JMxo7kSoAJkqIfUBlw1eQw==
`protect END_PROTECTED
