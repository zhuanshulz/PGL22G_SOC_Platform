`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M6KEzuH0WoYpfsvQhp/FMbfWS/UBrMgYqHCDRRkO4YYP7rGvgpIOIlM7khGcos5g
OTforviFgxxhmaPO2LETIAVx1swMTW5iBmXfXnNia/Xul5xnnaVZK9OfKV5gozZz
0YFYCv2QjL1Yc9RVYwLfeTJmGVwd9ZGTQzuqwyx47K0kglzHzB/VaKJWlsmFBqlC
TjYnnk+jzE4xKW5W13a7AtUtnNCvIqqcyWozgtLreLdJMOMy10+FMYY5J6LN6W8u
+mTSCCOxZtva94c7YFJYW9HhtSdHgBeB7BLR7bjXE9iOZFm0NrokvVunpdkG98tS
GBk8qv89GoefO1tJyVtlS8ebnCbCkSVF9ZXnUXMGGzuwUHx4eNQSebKE0Fn+RTqa
Sk3PSWAVq2XyEBcVozFu1EGYTGvwOwLiD6KZySLvIAB8k7/rleM4eDuBY/smNcao
2XI+RpAF2YJHJJhnuKrSgjPGUZ2GBHCijDZ/6J1gb7hWsquxBdkpQerQwmPfirKQ
V01fNId35GCl7jgZLKlHU3bWbS4XtsiXWfF+VWsXW+gj7D0FnkKSjJn2F3+lh7O3
XW0FuDRbYWzfSsBAq0DxTyk5cOD5lqDiR/NrvhjeMBaWy9qUWH4SGB9vzIbInzgE
DdQLf13nTFlY5Kdh941DBPWnXWrl8tOKE8EP9Yt0XrCfs1KN+6Z/McSWBKtrzZhL
Q3xtprcl9da1Zsgr7p2B+rMLdp8hwPFdb2rV4O2ltHWsBexjQKqwJNzHLsSlSIDk
g6NrJcW/ACQmqaczfehuhgp+v+REORlyCGuSekFzdm5ulqoFCeBIGA42fNr2N4DW
jQ9Kzwlf83V+T+qZfEz56S+tyjNPYIrn9i/8O11zLaLEj3ic3KPy1C4NUeo8ZIMP
Vbno+0wSo7TYiFX2IsgAyIhxHwvOPDU2/Sq+vzQkQ62dvWgFVAT1qzp/wNBSjlYw
bdBbRU3UlAzoNadHA5aAfZXh5T9/LNt/BcjHNg4i2yUZ+LK8N85qa0ilLPvWfHay
QcPCBXLRO2pzTR5qTvKtOMCQOcXWNcXY1cOnR9MREH47QyQUGnaI2k4KeRs/tHYq
dR+8KPmiALueKnjLTivmrnQmzx9dHWBt9sqhHKfevf8QH2e1U5//nOYIXWE6HJpG
iBcYW4yAevCLp8hJ07/SKrp2Lm0PdcutAjWeHfUw+TJEKl0ixuGSu2efiJE3hZ9j
/RgTynD9cLrwZVH0Wh0o6oYq0i798gp0MXC3NKR/3kccSBjQ6tSQCASxdkvCC04/
KiXnNL3dK6m4JqSSCeP9JxBXo82NNHjxVjZZmdvsFIxQeQXMhj2qyjq+tfrI2mJi
tTwTZEf0m/U4CpwNFKXSdtjL8dQgzxVtPlhcAr7OANR480kT5N9i5NctcUE0knJT
y6xkjGP/qrxVTE2cxTzSPh291IbYTc4CAzRhLaCmV2dILENnAG/zNDM5oChLSovX
kMqAgYfIlXwQ20GTI3K8o5M8xWdT4SbuGsnv7IlT2lYLGY1xE0L7OHRZzI0qqMZc
dgP5jZwN7P5ChSPBr51vWc0AprkJDr/xQWxiF4R4NbxyGQcJPWs3f/VkGLTs8sSU
sGMAiruYQHv7bxo/Eb9yVMe6MDjqXAyph675OxlRcj9irzm528Mu0+dTkH54gCMD
NLMfP+g0XueLkWt/a4iLL9pfy7098TCW07RBioHhKKpasOYMa3EoebAsXq3353o5
2GTPgg4pXhYyDc6BBU2ZvFaQh6EKE579kgOoyZ9V5DTxnOlHlP6bOU/1iOR3Je+j
NJBL1Hwm3O9YMz0kqMjMUQ==
`protect END_PROTECTED
