`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OXCyDVLLN7msYLtN3joy7bkRTR7w3QcfACFCZp15udZCP+45Fua67KciBCakijrG
SVJJc3dTvTfCgNBINLMQhROX5RMoahKDPOs+lU00dj13LPsSJgS6UG6+B/UHYhJq
UYz/z4FNi41M0Akj+J0zHn/Koc7FLaYe2yx84oNpJTe07ZJA//2lXnZljLX3L2MR
hP9kov29AVvZwcN81M45aU65zzNcr8rIAd4oC1JjmjLk0dNvoMSCSeYV2BJGatCP
Ooc6OOSjDjBExkedspbTQZGloWpnhKqsWIm2/BMLdpQ21pYCkZR2AD+Qa4aM5aKC
EwPVOGf/4kUi05ks6kU2KeFznYVrLaJ06qCnZ2XqXBFN4YSzDIoSPn7o55i4NnVl
kwlar7l1Y+MHSjQ4/O3r+377gbcvmLOvSSfJVPo4rNHK70IuhT2zlxrDzNVpHjR+
5/NfPi3wMn2nq6l84FkVvciSvACPlDNLhV28pBQnEmB0f71RXo8ByFtwetjIKmWn
o7Igtq1iZ9siiCfoalwDA3Ap2chk83ei2+EYqRzrM49BjtX7uP8JAayYuOgdQdOv
vEXVwSTzQp9F8MLcDAKybZCjjWlsB83Te8gWmZrWjna1uRYv8ZSQM6iUm6TM9K/4
+bF9Ro+EsC0IjW86OqRHg/ldLf36tAJ3ggyFaF/ysph7Ni4+xHhW+RSo61L3Xz05
`protect END_PROTECTED
