`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PyD7yG5HICv1x2R5wTPGBUY8pbQfmg6F2kMKDrqqQODsC5Qgyb125NeGTh9oL/dj
6NPFHGGPgrL5g2LXgqmOu4T35IRk79VmW+McrqTQrq9qw6O9+WM3Em1sODBhNa2h
pfbj9qjqMcnr7KFR7Il2cLe1nttN6Nakt7u0pFXqPhbQhQORrHMR/Ln0isNFroAG
73c3hkJp11UY1pmOMCKrrcSmPZRaoj/HfCWQvK7eLUQFYWk2UfgfFVD3i5Jb/jaY
7c9Hxwm1iknh2BRK+Tu0QA6w4fiE2qKrd2/zYjOWoi6ZT5jy7Fqxn9mIIm+neKhA
CY4+g+5Nm0kY5hwNyg4mJj+BHQg4VrZ8lzIlk6sCPQBzQS/lhl4sf4Z4+cgLz019
JtqiLV4yE3SPbNQ7sd9B3w==
`protect END_PROTECTED
