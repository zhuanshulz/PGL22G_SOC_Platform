`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iPHqQMsVoz40iDUJJeYnBnXYVs/dM+zgTTxeJH6ImhFpGx0wWb3ovyxQfFBzbT2/
dZzU/GvyGOdLQe20M+3lJT2K3/gzaM/GKsTW9JihykilexJLWWOSdGKv7nzO6jvE
2/4cuoM4YlC9Bhcc6f7AAJSf2y320GcBCRG7gWYMEificrMeMTCdVLe3CDgDT4Za
E6b+cu6CVWQslUjcp0mfMvjPpnrZvZaNbOPdlh34LKWohhWCsoMtU7CJ17qnglw4
yCrPx03/C+vuuE0NboWYqZ5d0QfJbtGtEsaw4qN5MqezJPe/X0+3y9iNyfxHvisY
S1b5/x89quktq+4Lj9Ko8PvKpEIAF/9gk3lfwUpuqHNFw5DAhm2qPwBIzFQBVPmt
aknkWGabthSm+rFGby26BwBjbVeApQYaDbJ246IxiNCRnL2u/dVk0b55GQ28ABtm
VRmxjP3gQ7nCqP8ijqWQ2SuOv5VQQVHXNbJmJzrZ9X0sEzajTivI2f10Lt8B1efT
3oMFO72DtZaPPjqKRIcQloLeYi76I1GyA5ZNQS1Lg6Mc1uuyfNXqD3KNMHdTZXHU
dNLFWA3NjMtI70WCOuVRitucHjQjzV1dTqs5hIaAaiqHWMAlgu6DIiW6f8EV7lB5
GVxZemTxpqzKItVviFQnT9gtcx2y/Rqa5dykM2oZsSJehCx1llqbwBugAbM+bbzr
fSyZwQKBRQS9krx8XxoCoF+E0cxoe0I5gVYcuKFBOZ9lkAmEowK5UeFRZzq9AsJm
wC3BXx9M8+BBSap0Zjfvz9RQ8EWI25VldNcBNwPtM8/WipTlXD9+a8+oJHKLUZIv
5wZgtlSSWxVfvmYYykagXbMffe+oTD4teTEroVeXMcMl17TCOxe3HLocCpkhFugq
FAV193mjRHfR4K42IiMZLMMPMH2yEUgV4AV4VyMqYlD+mGmjIkD871MwY2rUgxut
5ajEwE7TrkRK4VKRSlP6xkyohvolD6tjrJmfEzpDN0eJZEbJhXqZ11Aa5m0SzkAp
6tDiqBd9jWe6QssMvot/dmeirceg93iWO+ScVe3xCjKinAKiBKRGyc6JEvFr0fYj
zH+kts79vrGhMhi+wg10n2ocDR6TBP+Hg6LRO1SORCdOi3TIReE+xlz9JWAel6iZ
BUgJPd3S5Mb8hfvWHjld83bKEYNC6Iz/cx8svtWBfLNCchAU3rNnTJfSC9V3Ay+m
vG6W2OAYerqmgfpLljgBY/rMzUCz6QqgxoZ2VCTgT4A=
`protect END_PROTECTED
