`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
STyThIdioBgaIoIar60W1vxZP7IJXAHIitbjNGPMaGs+CdD1eEHJKJKHg6y8c1KE
ccFD8GdLUpRMpg5Qxhf+Y9aDAjJT6DgPK/33vOlU+UbpWwY1NPRvCYA5G1F+3ipR
0pK31kaGUdeN5m0Wf83jchu2/Vnx7wzOEXZZ5B28iT/FXV5cR7er/qaZ1HwKfK3y
mcNuvGuV3aALaHsZy9l/nufpLjhPLeIsmf+HNFP9FtBGC6c5SA4ob/IfXVRy2GZ6
LY6xSjnPvrz3F0axyE+yfMwd5/0zE1hCtlAvA63o4GOfqkIaeI2B8vKzcZ5Jf1nu
vFAwZi1VlzwqzcPFCGLCpMHWwKSjInpLFgtMNmAtfWdVnvQe/6WG6W0FPDgsDYIM
aC8d6ySmcaG9nU6+hMT4jxrxCc6g9JDZtvhY+7KBgjYULh5XHYos2Z01gCYGA6ys
NmH5kGclFE48Vp2SjkJRQw3oNLfQgUkUoxlVKzf77nyc0e0FbzDyCmmEge9U3EHM
OrWxUhJd6lVzWS4x7y0IjTfF5VTdaXgyoFjA1gU7LQ/+T5/YN0+43gYVV6wk/DuX
OyLy07upTmKcmHq16fw03t3plRNiBqTwc1NF1pnqfqsT7907+eemPS1wT9myEl01
fENn0/7n8Tk3B+RqH44omr99wMv9FOSrYJiM6sDZk9chRklHSAQnn/XbOVNKIFrZ
ifC2cJaDlr+Ror2uuOMZeeXb6VHVDwRetWp41fboZH3pkv1bUhpEEZFlHLiLXnDb
4ZgbQIuIShDZ2VDBKyfodTOAkqrU4VP4fbQp+0ISPk8=
`protect END_PROTECTED
