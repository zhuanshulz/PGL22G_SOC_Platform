`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5vgypB0C72c1LHqCRO7WAY4VQ7ac5WJflefxAlJb9iEPGVTWrOuJ0+lCbjuMGkAP
gCtymIRd6JmBxQVU07eIlsNLFN8R+RBuS+ImvVUh1pGaMbwhuzzi44yNl6kaejwi
j8xFzI3slGcQYOJzDnotkVseaIf9uJwTM4YKVEh0UvQLHM0A9Xs5+rCW+3Edr3NU
HfilNotYQ/fvp3AcinRRpFiJgmUPjk5UKRCqESIeOU3FhnhnCbKgzZxCdQ05z1Tv
X0vkQd6SKX+YjAYTm9SVd9npjkLquGkDJ7kt+QukJVC0YyBPWLpstnMbxy+iK+yp
hBgm/pCx+nfsFY2zM5khuQlHJNV0pMwr7cWvYpoYVe9VSquNGAGhf7CRuJi4Zc1B
CzJdjO+PC9dl8Gfs//T8ckBaIKNRu4GQ9HLCP4kQqWBRCS6RjE15V0ZoA6MhsOrF
CehBr+bg10Ha2uB36dFb9v3fioTb7+qCM8gPJPOXRz3idDQUHtAkndNUmvrHoLWx
djKowxfiLEXMNh+TDYN4If+74JyFQdPqlf03nPpq0oPhFK3qoncQg99tVrJdIPTC
z4dEL4Jkz2TDF++c3+q+M5PXImhaS0kMsPtVdJePc/pz0b3ZQWit860Q8j8Wfr4M
GZnbMWa6UbROPrQlp4WzTT8TFSSuQEj6Ext8X6MKvE0g7yz2QycbX0Po1x8KHfns
EeHL5BmBppGRqEX56zJNl7ZasaDTJ8WNx7PwHkQ8460v3+aViCQnjP1giG+BC5lv
bhvyqDiJTWRi37wmxtnfcP32zk6jkpNF/AO/HVDkTus=
`protect END_PROTECTED
