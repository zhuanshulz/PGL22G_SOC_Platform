`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OE43xUxM9PPF5pCdl5DeOIeB/ca9Zj9cxU6NLJe7iLDoGTi6E+iZCOU9ixnia+mp
u8MM7olMjOLiOG/5bX8UUJAbEUM6W5sGobKWDZjCrPHOxIHRDX8snUryRdozyUK/
Oj4pEBaVnjda2FqhaEV2mlmbUXumXC8YCtwxiJY2fRjIxWWVykrXck4tOG0wzhmW
N370/JvPzHO0eQutirw2wR/PQLV24ex4lUg3oKnHlGRdzDyd8ZFz6cQcoQblCXXT
Hwi82TWA+RzwMydXs74KLc3oLLMU4WaWj4YIoVggoles5wSU63S6uSFVteRi68Af
87XUIbMUw687OpyJze+rGKzq6slqKj1phv4+1AwozcAEi/P7plyWpa+FiW8vg9ea
NZKIiP+dAHotNsT6dB1Hqf1/faYz48yUjJpWvpvbHiDmiUpitzNLuJCkKIbcSLI0
jKUGXYGQocTKKerjOcvvKaKmHPaHq/1Fmrg/oCIP95gP4ELD/Vizy8Gfgfk3y1Li
0/lpLIOF1UpgPu+ignJGm96B3oFPMLhVLnxFSnmBihw7TMdJeZm6EWN2o41RawCS
WszlyUmHW4UJ57RxP2u7TL0cGPSTbCBOypQ6cDd4DDOQRAmpnddFH2+5emS7W3Yo
u/W83cAqU02CEO26fe9f/oYm2ptzS+rnLKWkHZ6SUs2iHnHaiLAk8sFLUmX98PFI
OPjl71zh8+jSlHHPqjjgNGVm7OnKlpq2AeLx+MfeCK/9gXwDAE+CNXNMsqwu57xp
/tR/Ebmxp0WlBrubh2IUUVgXN2YieomRa9YT6+NzfLFrwfolbdVxgPdu4CUHrvfh
YylFjYX8QZZe0CI3BAm0KPBFIzG09LCGqGMXff8ktUNS3JFIIx6doR3CjhUQ3Z8A
rbKJORjn3xbbo+jfbYJvf0gABeue3LRoAIuLv4xGbAhIZkN+yF0jZkZzZfEmyW5w
EPo6GGAVqUCcB4qe7hZp0SsPp2SSQoUf0jQHCBvtC+lHDLMRwXb+pxd5+leAa/Gf
65kYfouyFwdLA1KUoQULP7nzPwh3zXw6w7kJkDsI6sNmIzYZDOBNQSGJSMsMTUsE
/A0yneJtiUy/Nln8Il8QVWRotEMN7URc+3Esl58rW2i4boG5YTuXZCUy+9XTbfF0
XZI/kCY0/+FT/pvocOukR7smtuwGGrsEddO+JmM7EUJlOCqV5ostLrkB2OM0qe0W
eKkwiqSzxJIG9QNGJv7Z8w1Pd3rC7m0caFORFpIubLpmuuQAn5JeAu6OTcCiVMk0
T/y2a6RCRZNfAFU053iIbBILo810X2WA6yhDzoOQ9ISh0PkrzFRMzjo04dpyPRYe
tvqIHFLijP1tuRjNDxwE+nyAqsemdkL24T4JYJcPr3x9VKwSccFQ3BGs6V1KxS+n
EMfDnvj8JhL7biGezsbY3bf88kuctRsGHK0PzRWRx6vO2lB0GZly5fH/ySj4BF4o
9TcnmnDvBP69sgopbbnVRgZbFSyPpQbV14JXARDZGXoBg9nDmkuHMPX6YnZFXJXU
uthHOntFJeLEXNT+rf55kcTf9bwfpJdh7T90MdhOnLO2DO/3/kEmn7GbdO0tfNm6
V9jPOOf/Zmc3Ky3mfTAQB//7VjajO7XHTccfA7FqIIyn0SmWJGrlL6VucWHpX5hv
EWb383SvnzZvsicsoSoSqEhCmpoWONsTigEn/HJCLagtLXiFOiN0UR6k+KKVGRmi
JwjEuD2jL3rQx3hB7AX0pTTiO0gUdqg6+FZ3bEfjJO3zBYpfc7Ro2kDFT7plFE0J
iceov2CBtqfkWolh8iquIjNrtBNsJxTup49yyp80vZZtzsG7hMXFIHs5yx/gq/AP
pwc4FQkUzCte8BlFjKT2ssp1J7wEcrMoOvKxZrQpaT6SXV56PBiNoIjoqzPogxhW
ZVGmegt3s2AAWkd71BRrNHUrjIxiuWVLt0CYUUYE4o+/ZAARp7ZUeoUy/G/dGGoe
tMfCD8FFI5OVeopkbBLaeQaLtVUQjqr2JwygoRiN1v8LD6IFYPoiLe/2ZbkeMVds
Evtevge/zCgK/0T8gxn2v92sONf2YGDLFH/P4ToY2N/CdnZDw60MrGqI4ShGOBw0
10AeeElK0whvxdPAeJz6OG8gaGZtDhR4hONN/BP/wJ2rsbBjZ2D6YiiBfNDxDi3p
ammRxidSXIsjVP7U+VHJ3xo1/Efh5NKOV/E94apoMTUHWHGNP4v3yZuVuY3j6x85
mQfZp4PmLDQAY6/WySw4uWD8/XsF/qbyM248CJw7WO82wGeExTVDPXiNllYwbCo2
KSj6JirMglmCgER1ZAcIkXvdKMwkNiWqaQSvZOKByQzOaWWSP2RwVyfgnmORUPU5
kF/mT7TzzqsYTBskzkGazd4dqubQXxBVHizdbO5TwMI1Fevzkmgs8iYfMOOD/XBP
q2x+UZPVJ0ounJXbpm83zzEZ+bSO6QnFqOQ5sixhS2NgmVF5Ll8GfF0Q+gp96Oyn
wP6rZl2DI7pr58Aj5zfIsiw6u82+pSCWj57tR/7qwZGOrw6tjcsVxE3Z6LNl6Val
nm5cT2hdo13TP24yz4xbgJq32Ddf3LDE79/CKqrJpkJLpxHu/KLGgcMTNy8Ts+TA
pFz4KUaY87VS1iAHc55+/wXEw4qdAKKVukQM4jnlSs5EMfzf7xxW6p43SbMoFnAi
W1Vv6zh2nyv5n88BIqrY/9SpVAfK1qbCXFtXflyInYp0O7ky7iAFQpDu+j3Zar/r
h7CqNmoYU0ON6gpqxr8R9ZGQN219IpHui0HpS/bS8oYQ8C3BjGNDf2Wmhvnl68i4
9mNlHbVmiIM/v/pWsrTi2FLX392DpGTStTdL/W9d9X96IWHA70G1gLjEWumARx9/
wQn7Yd2TCHfFOYkRKcZ7sQhBcDOOlS70HBvXzPC8UiqO1tqoHtHG05D44zgMc4VN
/8YQzK6kzEn8Q4DmWK3O1LCNCG8CB1K2YjIvBOZ0wcc8hLKWzX27IMQ0MPid3qjj
dwGAQAZeD3rpk2+5Hr3NTVwWM3i6UpDpn16mr+qCkJM88QgQkxoNc6PAtozj/Lph
6k/yBAPbNN9GFgADmgYDV8zP9Vq8Dcuedp30AUl6QZ+9lvfbFPg1/zNOzeoUkbBs
hjWA+eY2+P3PnHpFYCbP9MGGxb+lhjXT92jol+FeB9QQCdaS2/PCqL5KpVdXE5js
3w5s1lIX2Ep7MLkh5gahsGLT4aCE93J/ndXLqZAwj5k09WSfNL6Oiy1ZR9ue8RZ/
Uh5/p3dydnv132ECCwPG4zP6OKIM6hzevY48JZT7CQ/BqNRFRytCThWAA1eRCd50
AaeX4zvfVsMiyh7U98ynUJ/ORGysk6ZWFZzwUwXHwLXDXCB1fiMboCtYjdS3jelb
iIukEogJgKhaqgTNs/i3Us9DsZ+A2HC4ap3BwWSA3MafbzZstxn0Xgi+2PmL7szY
fpqlQVo+1Nt6Paa7lQoKoPmVXVI5q58hnNVKNP0gJZrGLp+rRVp6BZ0DfjqIOEL7
zbbWqtVDmL1luA7IvY896/D9+QCCij5kRZy7YIeZlumMTgcNKzCpqKM9Rk1OwVHn
du4AIhfW7ji7QfemgA8oSs4LJaTuvrvMEcRXAbChd+eqEkjZjCoNvV0dV4tlMIJj
timvOQT7DTqNNndtLZO1R2g6wP95viNUMmGBmYIhcqOqPaB8wWizPqiUjxRa/HWk
Sxom9hOqXo1NY0FgRNMp/D8peFkO8NFLjqOV9kglgDc52smhY4QEcig6h/nVEJHV
KCBYbjKEttpGA8rlvy6hKLIUtv+16UtvXhYDxHTP1XiINtTp9pCSPKfreDVyRl1C
PAsFZlaU/oxg+9EDkO2a34YYVufoDmz6SpCn6q9DBEBVyORuSu0XgfYa6bPXnXsH
vdLYtJKLSs+WymHt8wUNfjJXUixVPs17XBBBigO36QhGEjJS0ELS7EbxZIbgR/Pi
6rN0MLEJg95wi4Gv5BcHU9YRIKBsDOtu+FZeluW4TF19o0DMQAKtjtqSUsns4wVB
Cu+xIwk/UrHlNwvtCNvs4zFLppyACEfytN8CWSwoPp9ORW4Uk4wCPjg/88CBdqli
8jc22TNRhI/d9qZHqBiSqiHDaMdk8/LK11Plsyab+ByMMfQBhXfcifcT/0vzpkuZ
DtjWevApO708s5357xXTL1cSTYVkoL16gtmPtpog69mB3s7ghEfRek1KQ1d4k3jI
PNRD+zCBTHwSHfmkjREH9zQmmni65nLb5uHlEjb0frQi7PJSCMrWIYyghXEFSi30
cPp/6lniNqm86IOTyKvirf1F9vkzfS6SNEMWo7grQbmsexM1i9NqYBG3wzfOXtUg
SfRYh9a7gnTEl9TZ8ByrbSHPYGcJdmjr7cGKvWkPkx5J32tpca+vgq4aPkMYE39h
SN6xHghA5JZeor/ckP5Qu2yzQAUYHfGYdLbDtYG/eiqHS/h4usEOgm8AgMiUGjbG
GEKr9bqEZ5H2ZKmgRWLtRT22+46PqTEK6LkpllQzUZt9xCnkziy2dHLsPHtC/uj6
zPaP5z+V5sRC5o8Va67hYR9yc76W4c0j2maxqxnwI4Zl4vKatZbAlf2ZMYG7fUeK
L//ISvaN7zYaPfRbYHBr7Dt2B4b5XIfLdDUOKrFEegpEC6gJ/4mZFFW3yMi8mQL2
klB/cSA/w648gAN3xFMh32ZBdAsy8mS6VpG9zDKVkdiZKDOtLrOgptuzq7iBIIB4
gpY5RaCCRWQHVnA9Et9vZkcvx/POYwtCTwfCPFmid9jc2+q3Wjq7XUrZKMFM9cXN
aPOSZJKQTpg66At3OuD9Fm9+nSaP5DOwhahN3n/AKFUFtziK2aYj0YiyeGyF0985
+AT4svsyOxZlsvyBNYj0nTSkXDfosxBpKkR6yLilRioku4t014c5bTmlCBXOLGdT
uhaj8CL+pipe5N851Lvw8pOVI/QfMGQ68KzKHAUD6ZKfXq1UnpLggec4E+IDbFE9
Jr7hj6EHTlFFZab0hiswtcwZ+JHSlJtIL2h9B9OYKjc=
`protect END_PROTECTED
