`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vyi6h4RNSP/Qwo89pI9RQjXFLpH5MVAtUqWrnjkOBPSUiN1SybiODJ2tqf5z7InS
dJt8VmLOLE3hH+Q9PJFuTDxEfv3RTuOFJGXs9uIFOKA1uAbg+ALoO5t7N3D4gpIZ
bbsPMz5MUUnNTsjOFRqrIF8DpMc0YA7k49rWzPMldUy/vTk/fiQPJoNJ5KC8+BTt
Ui89UX1f6Jsmdv9c6V19WtTOXa8Vwj0wjoHQQe3TuPanr6JZwnGrnMsLc/0RoWA/
Omy1dAc6Qp1aCH71zfTwGZE/DT3OrUo9kU4VapNY3JzWFUg3pA1ENOhtKLfb2v0+
Ky+NJOPB9DofZgdMCMb6XGFgZCN0WV3FhEllkioSHk0qIf8dT1pc1H7gY/zkU6p4
kt5hCcfOQ0BsaTHbeQRAoONDuIEtsJhN/ADKMi7RqXwJ6acL0rh7DUfEbB6AbJhP
Duj5BijPK3axI5QTGAoSfvqOjcaOH2URajsItllrwI35ljaJz3Kl8nFHLXIeIPvS
L+SQzPmBRlwMnm8N+3L4AC8NR2KnYQA2Jgrs0x3vNeHV9qFxwzNqAMRZSzKLAmcN
Qs/F7/ug8zYbt/irCYWMtoEewFcNjT7a+IUC0cQ0vWur7/fCcGH4vserheywW+Ml
OsTat5mpL8rG3QumMadPca92gqH78TpVY3XY5XSWSZYsiGK7uw+9+ETH3JUmUM7l
zhb0776piR3u0ucfo8IxBIYmgfivzZrVOTjY5osYMRJbmF94eUJ3EWfHVDVhQMSy
blBRbiUmGOym7PCAvnyBMPRVrbDkCkOm49GfW2k5wnSDBXwqfQDegybNigPvP7ql
0GNEraUcnjwCOYc5zd3NQg==
`protect END_PROTECTED
