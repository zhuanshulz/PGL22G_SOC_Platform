`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KQFPLJCldfCGD2zALAgbQviJb99qeDNPWCa/Y8BN+nTvyajGEoyB2nQem9GwU2Pz
0ifqcmlqyAKIMmbQ81BTxS3wkuNxSNE4fx1ust/hoYfB5Ti4CPn74K+u8akrRgLp
brqWI6dgmG3wWnyvYRk06yZ26+VpAeZoIuTSJcNMXfHd0H5j5L5p4LOcEdfG5t3q
POgR2JX1iSvfK48KwEHkItnDklXKwWQMqrZTTupbY7w45J5D9Yv86kZ30U7GFHzT
pXoFcc0ZyriKcRmaQe1wvG2WiuYdfKHibzODUSR70QYH81FDhifLGe0NXNZY+n+A
sZP8s/C3AqoJIfeFLlEZLgaPTxfREfZDQO/DPvBzp8Fv6t3Im19EOYrVB6wX9pY5
YpzTKAG87rNrBlMhfP+iAP63dhdP2ajG96qH2lly0/wAOBRRgUM8DwHVZim6T8G3
65K/4Xh8D/UTRZv61geDRWV1eA7VweIQxPMEkSivk0BuD+fIvjgciH1d9ooiLhFP
D7F3HYi3MwZ05yTlIfmARMZYdrXApSBdMzYmD6o2etZvXsj3bRh/c9KRH+QwkGT6
LOYHgoCS6I01Bmwx8iXQScUtecvzAihWv8YmPk4kyVSpFaoPFtNN7cB4eMQzZjcV
xFUx/H1bZ68aU7H8iHKbe9iUn56IXzZ0g0A013pkzymhV1iSe/vqBbonPoJ6TsQc
6/8sE3DLHMV+/eS3FCQRz/H01AqxAzjBTWNEhko1A7Z1Ex4sFbLXvXlaGjgmjdFJ
IYur747Ul4AD++oon1Pd2YaK8k8PEOiYvof5vNvDmhyTFGJL7ft2J7sjLyRr+jZm
RCRkxoVyDIOZidKdx475tbHfGuo0wjtV+1gjyci6v3vbgtdFNSPIb86bBU96Zi9X
+l21/fbFCFyHnszBKHPzhP1M0JCi0BIBu+kC2raHoide7n+EkJGKDOlLAkVtkbmH
nS5xX0OFp8DugRKh+HtMtfd9OwxXeR0UHhR1q1wllgZlCbyCz2KZoQrmoWA5tq6c
+6Nu/IuVrlri+3fYMRB/NeuQ1ls/Y/jApZtzjl1QP7rRLm3Kxip36ZQRSOgYfmNz
q8p/e5aWpPV/RJMzN0WNZT0+iqLgUlnozb0w7PC2ie5C+OFs+jqmCa5qLQ9/XhJw
I3og6yVNZRDOh/fRvYipp1y7YvRCLYbvWFMmq+ZN0S/i8/WaGPPbUTrixvxtF/BM
sUP6pPLWhv5kzzKbpf6/LBgyli7rRFgEaRLpTSUDA89SXLuU3NY05ykFiy0lhXGH
CAilNeiajS2apyNhH/g8fbHTGVbM+CVLgc9kKC7kZ8uhKJNjg1XwVsXLIy1D/fWd
J7RXzdkoydHPd58sV7/Rlt9MIW5C7ya+XY1WbZRwWNGu8MSWL6+7GlK7ZASkRM96
SEIdfG/bw+kubEQMePAzPyiVQkdDyuMmv40y+7iAaIIGjM145c88K5Ck22TxP67C
VZryfheMjm2UtPgkmZBZuZP8wmN69xcGm/8wspNiHtFbP5DoudkhuRkqCtA+QlWc
wGw5m5XupCR3h4ShPlRRAprSxtgfXX4lNIpx2d6cMYWkxwYnkC8qOYgojKEFWf6/
T6cF+wXw5dBt1Sk69iTPN7oxQdnk9XL4eE+V8yU7jl2uoAZKaBNdDVTGMXyGDh+O
48FUodxLBdLfTxuuJ8mcaQ4QSLzi2jjn44CtgLgO39UJ+VKVT+xWD3egWD2oAfZ5
HzQDJdafJ1yux42izYMpbx0E7GX2AKQxmaTFMCS5dawWBpXaLWvnMlRbcUIW6FS6
AaEtcVpBB71Lji2o53WzBS13nfCWDt6gsl7BJWPeJufkNAl5VScgALZfKL59bYlX
y0MAm7xV0CMN2UMhRzdhg9mAgW6PQf9n9H8K/cZag+8o8uwmo6adP8XqVuZF3V4K
/diNjkh4uBq1ft8LhYY0N12bzX7SKDAxZ712BYVzFoRS/40HSlx49g05SYWiMl4A
8GgNR61LvOXZAs4K7u5VwGURR2zxPp/j8DweinFt1IMp0rhFLf2XLBrqB09Ktj1x
T7i663xQNyCAppG6emHQeV0Ce0gnCCqjKJ0F2cEuOB8NLR9gtiKvqlWhVwcXKqDw
hM1C/8DMAGI5/v4AaGFikpQi6kQOR02XId6P9l3xTfDGTKu2hOKvm3qs5Uo8Dyqc
GToqRnxgvQio8u8laSkDxGq+w8OcAFJBLE308fCxWfc4xu7WvN1YnDLkRaZH3o75
cuVU+d0nTs+VFE98pbeTmoGDeDq22lI6U97VCGpTKLCRQK8hWH70/wlhwrYGKCAt
7XotwXrKa3baPhM1sO8azMg60YJMdPlWGDscArenLDN3gJUO+lK4Key8IBbaqD6i
KIGPkrI9Kj1OM9jsW957CBOAtUyyaM8UhLATulyy4rgg8zsQpuiQKyeDSsyVyjqK
bL/onkeRqPd1ri6p2BKcReeZjVqJA1JITM++2NwHGXZgb17SjlduKHAxBjjJkdVQ
61NiERO6hLh0jeSk6rLwf/EXWHFEygpXoAkrRy5OhUv0umOp9HvlHOnVrHQXPpXb
KMT2CcS0Qn6uAT1eTdJnw4yakT1N0uWMZiKuggByghBtgK5vHzzmdVYZdX/aH6GC
8qPCYv0mKuSQc0WGsIFfPRQvyextFCsmqs/XLz49nBd6kKCNOmv/kHEE3ZJ0CSW3
UEH2dH8xC01PXYnz/YeTKH4BG6umv1lZWSlblLq+Dw1KF9GC7L38hCKf+C55Oe20
7t4AJOpKnrsVuXu5MHnGWyYVkfLfNKRt7mR2fv11dBNJgGNuR9ctsQkoTyDfhNTu
+6CispMRBcybRxgW/Fuo899Ey3+brFiMzCjBfNkPXhXYhvL4y3xHlWmqASDx2sTB
LcLcyUCMS3056IgflbWcsESFzRY+1nRfQVrfPglGn2iKM5ioo8W8dNxQymyybn9p
jfHF6seHLOg0VcPikken4y61a2SiL06J7rNCRI1yX2xfYWx8r19yiLi/TwTm4d61
HAEudkLk9HwXkkzYnGpp4OqNykrR2v7HmA8XtILMlyl83NNCeR0e4MMS3gJBrG1o
gyM8H8T0CvjvfpIVABv0/86P0gMnecGYJZ1uZOhE+Zq05/J11tOZmxI3FxIJeFhy
sPws7oRrz+IUgBph+Fg3JQ8QD0o4DxYJEMTcjX/4pVCnGRNTvbA8sYDmB9mkdoq2
DzRH1HhVfskczKAc5I1U0ScyIXa85T9TySZbSahoSRikv2zjc1bNJnIGu/9200cj
KNRmK6sJ/s1Mrra70G8RXw==
`protect END_PROTECTED
