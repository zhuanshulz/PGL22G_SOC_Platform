`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TYTO1wMB6/YBmBiKjRcXcdKgX6iVxlhwEGGeY3YKUxMDSib8QC9eEMeKy0fB9MqJ
uy+e6xnenlQMsktazHVya0x3NwCPQ1lyEoPMnZQPWggZQJshG7BO+oROzGn8bhMT
2vnW4XUu9J0QRDb5TqdIcBYlSFiLt+P1zHLmv8rRu961hwgQa7lOZQz3hsDEq3oy
RML7efsJ5fxzsW7QpPzZWO/M3KJlYCs4w32SNdM8VZtPxJlsKDLop97zYYhalJpw
tX2OsLWZJHmdhQb9q6a7kjW7hZ6F+SHm/hf7+15jWsfCqmIFSdKEKzFTeZIGbBgD
odyEeGLIpF3JDM2d9jfB7GQh10gOgNE0eJ/pQ6nBovpmlSK3l6RejCrJv067sbSz
BHFCAgLpJ4szXqopNgqTx2Uo/Op3R3zChoEoRUlLjgrvApPK69aQxOMhryWe3Ti2
mdXJ1P/GzvIiZ14tBbXDoiw+82jD4aoZuigQ84ba5Hm1Mky9qGQf2VyXcKtoUA/q
sN7gNDM7vVf2cUGY4mvIMai30TyA+X8Z0sOAa1zcFxRephMOWe6Xd/AlaEgGUWm2
AYDGNAsORqGN+Uf+AJ4bbD0VCGMSAUDozIJj77BMJqkAMz4n7ncWQ/VJzlO7eCXh
JYZKDbiqWDQROpRbxvijg5JskZiEHD46/AoAP1yhMmYxfJP+IBHYhGazhacLqczU
z6MyjzfMkpVYZCdVvDRoDzj0XW/oo9lVWSDxM023UBUo/mPWS41QOMg2UDAsoS1E
P+F3EFRYqgWBOHwGm5L5ZeEwOAyZib/eek+sW0hIx11iDvXG9zcEZQEDpaSRWguV
OTRWhf84FB6zVB3c2PPgcovS1phJOeK3QMSTVAC/6mTHKPAUFTT1FcfyIq7Fhhoq
OMnfvdSdePe93xYWpSA4CFj2dYl9ZJybBLjOPYeDUl4jTNOGcUF/y/xZTrj3wWxf
nCjOyr+ZRWax5R0lJ3vWrA==
`protect END_PROTECTED
