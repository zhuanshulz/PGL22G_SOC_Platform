`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mE0L8GGt7UIVQrFlCqn4oYws5Z9THfkteluPD2w2RXvoFl24rbGnAtkQNfco+YPw
GvqnaRP1A/5H0t6KotjE5xOoQ3E4ShOVJOWxLCpKhg1zA3oqsSfj65LJsgqgGmfW
kYta/Lg99CBMb/0OTz9pT87nPcmvyxTgBZFXSidwFJawaHBNeKxFzV2uFqf+1nIk
GL12+kMkdZ894+pH1UopYu97zVbtcF4joMCbkJH5/hcfbfAfHTrXuiXbGGX5eVUB
st4qniau9j/cHRUIFXUJWYpud4BS6Bic1T8guBejeTEkix3IYjxxaf7/NzaR9NfS
uxDTINUShi76L6arQ1db1hrRNE3fwNmuyHTdvsZJQztjYagZXtGLC2BKv+wcgsxq
1JHBEhcz7fl7E9FE68fFhT25+ODuSR+pYJRGk9nvqG2GnjIPbkf0h9Nzw/3OTVbn
xzrzfZ8h72UnFvV52PYhdFKbTjhqw5FW8WUEygtV7Vun7wGrAzvri84h0szLD52C
l1FOJUwAjpcgszlgRyxLKxgpyZnC6UriVRZIyaRdWMOksIQQl0bc4tsoEyUdzZxF
zFFLBC79I7Q3eKWiC2cElxjLidKgNO7WCPFrOopytVWKcGD7blmfyINnh4J4sEZe
Wa14fggqL2ErKBY7TfHKhqlRbh7p6t/oSA+fFwDX8NGt01ilgf98DYvs/YQYQ9XS
izIaMx0fdvjEXC1oV3lqdfmOLdgBcVFMaU5R8xmE86MrOANzR0LZmt2H1RHUwylp
HQjh2seIULDuoHGNJopDAIvMY6MZ9NUIkxaW5gGMaN5mRq9/30Z/I0waA8ofzz/F
/DwyXnYX9rsrdOEMQNG4nRgLZe4vTc2w3V+0ngFSAjWVge7mLJY8qScZCnDPFYy/
peTnnfb8qmH9V7CzxKFPKglC5T8AcJmJbG6z9KiUN+3EEz0yKEm3PEOW9qOnXvCv
jw8KLm9r9+pZf0GO0g1SWyWdMBLLVuSEdBN17h7GHmz5qdK2fEdRHrzA/bvNmIGt
raM39p2KurkIMnSG8b0ygSO8tSOJ8y4CV/kbWRbMi2coYI59N115x00rb4nJ9OeP
K0ZC6PagZgm3N+atZ2717A==
`protect END_PROTECTED
