`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pHIeqsYW+1lQUVF6fEc3ImTTY3K+uK8lpm5eWoRK+WUwAO7P5rD8PmAL+n8KpsxD
o92fG03y5P8OPlDhYND8IQ7YOTWSrxndSvfyHFHfEjAGobj/RuIbsimRzTUne/4I
GAo5w/D0Nrywph3L0lZtt6tTYsUQsqjgsdwen4lm8OahZkL2NCU26yGTgEe7shUa
50qjC0tgEiQYD0CsgSg3DKnzGXdj5hNBmN/W6c30jOH7IjoZWa4jREmuXh2pFYdV
1dm8IlC43j8G+81L19Oms/l4pxSHkrhx5HUuic0uADonxjHxQu0+KjJzL4GWxVMS
/zAA4BWeYiNeF0U16nbahLbVJLDUfDW8lwmS2q5dOcsWQ7YTXwcNFZ4C3GUuzQkJ
aVsyeMF2o7YgsKADoCBbzfgbyP+mB68vhTwyFOsVaVOGtvLYWMskLzc78CImRVxy
4XAiecwzeWzsAgnsypxE8cvc5GMORoa+wvMKLEic4fiGR7InTv6Oz8wU5vpgI6Kq
nymeUcjiBduUW3F85rsdTFDaUeu1potJAd08shFJDraAUi434eEhxAEJ0x76XsDa
hxSq9Tspu+4Wp+EmZ1mbCuwszi+v48T5ks7YwccO/5yMVUqIkWL3JPX3ySfpGRou
UjJAugKUYsXF6A2Frv8x8Yn14zyDHNwTdL6QS++6+k82Y9Whpm8cGznDja3j4c6L
nqykIx9cQPoBjZ+TvoLIqP+Sx5lS2ryvpPeYCXT2GxckIXHoWNiiiU7PX/hyan/K
o1pbKLDscf1THRX7ePGy6NKjEP5oTQ27N11ZTGLd2rA2c9h6fNkFMGyWjDV65yr3
C5G/d86l8C76C1wKIM4N+IvE+byKf7YVJ2Pi8P6Q5JEU8uWMcVcKtj0pd27nNN1c
0Lj7etrXUpPapRk8GS99vfUw+b9vOtBkjg3oNWhW6l1mHQkZWAFmniLtcTw578vB
ENGQQ/nH6a6uK2hLcoFBmEOgJtiFXznAbnF/tnEcnD4ICkypjNp69XAKRujlpJwB
GJQWIZZfT7L87LdrTxvyDxbqP/IkDyA0goTaaZn/rGP3wad3tuiJkw8wNljpMJaw
kddYSb2qDiGQUp/KAlZ1Auz5VflvBO4kI+mfKRyBqhzhTh4cM8v+48JHDMqmK9b7
ttbA3vb+h7R8KSgjjE9Ft0hXHJEzDWFOyEe09qo0L6Ospf5g0rhgJAzVl9kSLoFN
2gDBG5gmHJUGuzcPyMJUSlRvChKET6sqDIHF/HdrQC7KRQqRDzG3uyIt4OykbV6p
gjSK6OUzyLt6I0AlzzRwM9ZnR8ykoGNMl1dSJUkaCYxyHH2ZCRN3yPt7N6b883C/
2mRHTpFVLAV95UArMl1UkOBikgVNleKrN19x5n4l2gX3n6DsoKL1R180uQd0uu4j
etb35WolA40akb7nY/lus38FO3dOimL9Nr3uDhqKbk1QVeGDXQHDsvr9bPLJsCux
BN55R6Vih1U8OIU0SMyd5q+xsmAR6b7Mpn9Cn4J/bo/9/OTNjZZP8378TMI5PmjW
P9zwYM5p6aUVEloEgPD5fWMoriBLdGZ7B+BAwFWFNT1mMAjDis8VceTJVYsiM4Bz
QLpSjUURyTRXYUIxgU1ZjxzOy7CpF/7txwh+dBjnssIkAfMJwQG2obxcrIiYs32/
vIp8xM2B2jbRBxHubfLplI6uQAw6c75uJFqDkN2RBrb4reOZefqQqgcQY2482L+q
9T2P/yre+yaE5l9Yk24Lxq8M6qTjI9jE5/Fnf0ExOqb+ZzOdT70Y2WsUJsJV1Q6D
Fdu7IhuAL5PrA60zQGAVVOByzO/xYWjnYgXQwrKLu1D8L/hoCqf4k2nwoqkXDFCU
mBZ0WTu9AOCxJ1KR8qNwIgkxSoDKMXn38ESVtcOE1ycO2SnQC6QBEdCmhun8fucV
Fvwbg2ooyvsLPsWr6bQ9ikr04qd4mgg+Ok8LcPzgMEBfDJWzF3QXQBunUX0UgVSA
6kDqZFNvrQUEJsAkVKiX/VeA//SozmAV4LHtzqyS4c1uQB/XmqEGmA+9BKgWoBW/
uDHeIwyFc+LdRIYWwCpd2SteRGvCgVv/XF+pV+rokvDxIacik5sp4TgVSTJdfIu7
4lDK16mR39eV75ouYL7klgXhHA49FvlZ3hsGE2yjoDBtQ70UdwU5YbGEU1mfSU1T
CAdqXRoOqcYJtz8ONw+X8xWSOR+Sa1eZ0haQ1P0JVmijahs5ChJFQj5qniJ8ScXL
dE88tge45hRmEde3MxDHNEhORf2qzWpgWWUD7H8S4o5IIz9qCXUtXsiaJXLT07fJ
8WLvgElnxZEA2T5mFR0il4XTc1+o+c58xDY8cjvTUOe2wDFwa/qhIGB1Ii+H26dO
w+J//dsJlfF2l3abT36rl4rl28QSm5DP+QZ3mGEQ3dqI6zitno1AA5LpbvuHvG1J
HqZX21az15QZLq45JZmEsBKSPAU48Iahn38kPcTtQB8=
`protect END_PROTECTED
