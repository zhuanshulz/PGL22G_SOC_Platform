`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gjE7RqUzfP1T8Z+GzakPSTwOA93SXxxQxH31NX8d2AwKOrN3ut85WhEJ3jZvEyP2
EkTPoX4dHJtTqeqAFSNTeSmvaiQ4WInsCtw9mcATLA7N5DbNjQmIZWqeWtPLYmL+
TOhOllEJgFkk02Jtui8XS3bsGgW2Yh9Qfg02pvBeFRKqoxl+QngJAlQCgnjZVZt9
FL3N+WN2ac2uSNvw9uVCbf2BKafzmF8z/vhpQ/Yxcq4F4sL4UWrEnFP1+jT2oMKf
fKsWt/PyNhFUKUu7Nno07dtG9yBEWyy2AtKbQ3tPNHmFMtSiIva9t+P3/Jqu+EIJ
KQjviXjQw6OPHe6lihFSmnKjsrSbubyCHvBgcIyv4ckr5OS2DVVEGVoMiCitl62Y
`protect END_PROTECTED
