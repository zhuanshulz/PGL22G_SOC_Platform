`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LmG2x1TlfsY+fZ3Hb23sNgayZZGW3Ph3N3rSkGQhm2VXRSRYnLRpTaMt161tAsyK
cSwBv09LXKs8fyLn3gNvuC6yLnurobnZmX88MEDLILZdIayOgUqIKoTUgfwJsvlL
6tfyKm1YlgrGS3Wh1A+phitCzRc4oE+IuJ68ykM000TZ4HzQCh2W4Ebj5aUC6JJy
U4SuH127fMUVPgZjWlASeUxvoV+prB5Bjx+pAEKz0X/IjgfOYdzMot6i4KioGUUE
h/5Vvtr6c1J9OnUtVwIMfPyHwWguLluClsM08TEYVw+vfCkAudqerqT2ag4HXGmK
x3c8G3b/rGxTf+1RiFA8eQ0TL9pwbRoJriuLbBO6h8rMOaOY0ymdQPgvhAJJ+l6x
IsZFqf7OTqZDhz900esIjmz9PnzMkDlNQgi1eJByYLIKRvZ2rkIV4IsvWbep89GW
6JmT20fGZ6U/BlUGZVHk8W+t+I+TcRUCRdHTHr5B4/vo0wk2g8WZmR7UPYWPwhDI
vUj4QfM47/8LLkRroKbsmUfQIsYVyIDsSYUg3ZS+L3UKdBRlqQbnnwhvQMSEDJU9
PU4zQD2SchpRaKbnZlga5sDpo8gS7rDKwFQtDE6zk0wMQ9DolhsyXNQRuUxLi8YB
zQGM6QsCOE8zKmalXDjT3SybvI+rEAx680ZDJ5nrst7Nk7vQ8DmWxtUelGGBVRss
J/Cu8IQCN+h4X8LeIfqgMbE8saYKgJ42v7PSxevr5JqT3XlAG8aaaqiPRNiGLjMa
iYFzFauCxVOzoEf0QIKmII/uQNd6j8EqDsFV2efKu/K4sUFJGIsy4BpB+9HrH9/+
xXnwoeE/7d1YPgSCTi9BeUxrne56c7XNMssIjoQvMhCnDSqJRxECi5BAGjuDGfM4
bwyyFpiqfNdcEI3EVM4VXME0C5/8NBAHallhVrvV1Cjz7pa5zs0tgm0w84uewugc
YdAuLAbyZFp7vZSSSOg5asnvtxoIsqkHY5CxPIoBat7lu4MG/dzjHthW9Kn1N58F
F7EG6LHCFMFTC1zA8z2/F+nzu90PUKpNEt0q/Aycb6s+GvnsvHnKsEJ2ISMq7ba2
a+Yaju6U/48JIpN8akcBDOdn9Rh+4ZCCUYYpDrdq+mX6Z/A4a45fSOGo0Q0QMRFg
EDgR59zrvRI+OhnkmjGuTlIUO5uI6xBgjETHV+3MfIEIVMly2V9BxCcng2Ys+zNF
iFSbgJk+wy5cGJSq/1tuq7jjNc7h7+CBS63CLv1mxrcnei+jq8IysNWfpzYSmlRy
lBc129lMRVp5ybY1/NytqAsi8eb37fOCJaPaLS0wRx9SO84vU79mikOFL+OXRzhC
A3QQOVC4akAccptM3sKHasF38Rg144VwaZSOx2WuRUUTrPFdNGseR8gaJpiBxpie
qkFfXGQqWHiKdd4/TEwUhLF16KqEmVFiDneDMQKeUDFTDNLSsz+ux76Rg5aaEdeI
j0wvXnelQM9JKROC3Gy2R7GDjNrvkmkkBJbHEeuoucx5S8KvpWet9YtqLa2GSRen
YnIeKXukYOb6bOIJW5J0iClkwdOEuP8v46i8qrocWz/UQ39q2i/WdA/JJ8Tm+y/r
LrzBKiBfwKMvhjZ3mdXZ+aVAvWCGk1BdvGpxvIouOiFGO2/+lUS42t2hpx91DG5u
x9mil8mOOfmO0zW8XYZkY+oJf3l5p3m9D9bz4WMinq+0QTxD75Hx0zfdJv39dnaA
lGPabZrjGNMPUJrR/sZpboQzgg16HFLnem5OU819F11z8eP7jijk4zs6wfsvpxm/
e+LH9cKikggY5Ub6SwhYkDmMPfv1AJwrvb+Rn2Kalsw7KKTctLQuViQqiQh54Tns
g5/UQUA5reS7Rju+2EpzbLGlS1jNuw5ZuKj/Wa9D2RG2emP8j0DU5nWvH7MI+SDO
12hgFLvnkJr3S+R2/2zB99/BjFnkmOq4MiqZ44nKc10cHVz5GZ6j59n0spKXCfXg
oFBjljjs8Of2Mrguf8iZn/jp1P9atl43JKZ4mqwP1zsDJ2QHkTg9pg5WvDHFyoIS
VTthVl13Jf21wWf6PPUtDvdLLXsFwMiXpdsqRi3aG1iPt4w2znZxXOI61sPqc7e5
aNwDmyaGh9UR9nk3oxee2G4pgzBtwEE/IuiXi5ell+CeM5sY6DpuB3fL0ps8kCZo
LZTClJSCAxlzUJeIdbl5d3NJB+bklMNyloYazk7Rt0gtwWHUCd124vRp77QBXFfr
0u9gNje/+GQ4bpANeW12Olqj5YtANLm/Iz9utPImZysbsqjjXoe9yPiX9y4Mafus
9H3VNICTmFhFC9LSjKJUdhEeZ8dco4VV8vj0wUX6RVNAoQ899nJ3oku15mD5q9rK
jvxm3u0bUThdEdUxCtquJq5ZagN5n4nt8xNb/ot4NsepZyzm1nz5/m1roT42lOJW
rOAHi0K4PHaDD1fOIbdyf+5EVkzqnhk/zNhK/w3IlkZzHPzVxQqPzJ1n+oAbee6p
k3fpzXVYNnN3yjpvRTuyDAuLKHhtPIes0xOyA0vJ+olgedIUbRH4DfB1hT10kWHI
RexHR3TqNSeqVtKW6JTQvC4VwNOzGyrWjxvAvQI6cU5TSXeQEX5hS9uc4vX7P4VS
y8FEZlA+51OmxM5NrYFmwhdphe+YhxPFHPuzJuLmqENIfkxmMlVSgMxOBbAsZe8Z
aH7zzGLgwkfGBjikjBW5BNSNQn3+ehIPgRG3hM87eKlzKKvogoBSkJKc6rn/rWPJ
Pv1OfMnL3YsRd4OBo2JZxoGTPwa62B4POZ1aXqtzvpgugjNiwVyA60m49xL5G4lT
UxBBssj+Xy185aNGGrBOSpQdap+wsf4AKrEYBjrOky7exzj4q2YzdfatHXxpVDKW
xbVlH7IFdLG1AJYSMlLwuxnYQPm6oX7+lCIj+rOsWDlo7NNsGR6KoCuG9RiRst0U
c7R4yilkkhMoXZ3/CwqVkENKR3NGVCoIapRboZh1P3HvhwANSH8aE8ttt08jKiGG
dGL01RtmVvs0dBkA6nN4zgA3ICMjY6Jy6NdCug0ZvNAPyjd5Pr+UDsL6yXpQOFY/
CoR1NaXuKvtM0OL9FvGESi+6JKGg+VwwHgONgYHAQCvLFoCg5Z8VkiDN7gg5LuYW
bXFqf/vIbH85U/Fui6FowHwSyvAEubkVrxpwp0jSHbnAF3n8TdlbaMQ7owTx9Y68
RYUPLbCo5ujJwXBo2ZWH5SNUzFvAzcY8nIj79JeAYcpNnA7UNT1Jt9vWJ+IPNxU+
VxmkUa3n/11Vs0zumg/IVtS0AhMrJRE6ON1ghovOs1WT/XKY48Ceofoou7trcpqg
vyCVm/Rk9lzOMIFjGbcoXp2uj60jcQ9g59q9ipT7Xnx0/EZLrkGl6+kGHRzchCit
AuOygSFnrgCUZZHlXFdWSAUmP6kkkkMxc9FJ2zn39tRhzOtQrcaqBH/gHZbpkqob
ipduPzGSISGVFSM79SVxoBctT1p2lxQGh/JGeJIkcRifbs8D83Kw+ur9lLJK9RSt
UyE8DKe1HoW5ShuUPW7+Gco4Ulw52ZWxQkul1kJtJV98B9gQkID2zSGFSelMZtNs
R+aMyREvIQXCcGJEvbQf21YKBPKw4doELbJaCz2vWC+68jtCLewD3WQK5jvsXCWW
yTko3u1J8Ctwfdxyhz41P5FYBLGG5VHOdsMSchx6LChnyfhzeBwjtuqSPxTY1f7+
4/R70+A4h7u1G86naeeRH+ekzlqk4mEhs0tbm77vpRw3xADtNA4K0VNwwWQOGNhg
fffPcgFhO1pSwfWC1asdi6QRuW2LJZUWRIWX/pKEX27muJcW3nZs7P+k1kYNXzQ1
Xqqg1A70P+pUzMk8N8Y6la2EkkyF90tcXEeXNiN/YvF8NMHmBFlr3V6v+ibxCEB/
a+k8eKPAdaDdIYO44ruaWQ1T5cBUTh4ltw3SsB0dA5MuRzz6reYej09Ly28qV1ha
ONxplJ5J8pdXiREZXoeKWEokdiQsklXo4iY+iDyHHfBgUyv+52C8O30kt7Has5Op
5YTZBYywtL/lXag4u/yNPxlHuh96dNS5tBmeNg8Ayh37gCnc0uz4gO49SfJ4FGlc
3nnCBdSUYKaOUvVYlj4W//H0LwGQ1FhoBWVbDB5nZdvRXSuXefNEEObyxCi2Plzh
b+FX3I0o6K7D6IbK5cDUT9kaYEWd+J7P7+saO1wnLe7w+5XBlzz2K7HSyjAOmrFa
IhD5vCFvZ9wj2LXfUzRqlIkPtuVm5X9+3sTAvYC91KGZOgZGyMuXdsycbfVXeYKE
01XVxYU8/2DbpIXw14e0q1OA1SyM/uX2GVQLwQk2qrPco3HMG6LVqjAcL3xt2BYb
UoqbICJ2nVFVp6l4DWarqCxeX82dldqHJuxSkEIMWpSMXtPlcgCZuYIDndPrDMIl
jew+P2dfgZCS99TFngPLuMSSGPhjTPghVsv/xTDSc1nRsNHEwfHTtvEhiCI6Q7dv
JGdne+xLPGRAUYLpoXk/+AtL1Q1sEbIlW6uZDAsdcroYwCAayIZ4mdDeplFgpV8p
Zb7VHvedATGBlkErVuTOz+9t8HZLMl1XFyQBuUeljJ9RdTGgQ1whymaGJUoRX8kP
et4EQpu0/9eZ5H5wxmYWWCOtEPFgyUyvaS9CB8a7RD8YkPhFXXlqO6k5BWc3F581
GV4GpUDozQjCzNu2UV9MxR/LevjvS08K68m3EiKsp/DYVdJgWANGPK4eUzWCKaM+
/HTBtXM/gNsC0ffqk5uWGoTijWZ+u2YZwzjPutUht0Rb5G7LKfkxFj5102ek7cl5
mMeuhFoCKJInQhJ7r0+ka2EqQT8ncFxq8qt7YCTvUbW392by76tw3B8NqrJJbZef
k3TEl4w6k5udrQ9HfwOhKwI5j6wdO4m/wtTIlpWrlR/0CoUkfe30CuuwkdeVIjW5
c/WIoIr6Dl2u19w8WqWG+BCZ/GK69G9KBzL0p45qDoP5SSjMH0xu8u4ETw3LkbHb
GWE9ypE8f7pOQsuVIh+SNSDIQ6Z9/LIMYWYdgbhZmsCfzhje0xqwnFNoQrSq/ijZ
O4YfyIOTBfhuSgZcKhdBYBMpAez/WJ/sjbX1v8lG73jNho7f26exZfwEqND/4Rf0
7QLnr6gKhhD0BpOKQjFZzRdO9BIARSaUFIT8RrWUaGUBTq1x1JreXwE4z5NZiXTA
1UNPbVypBzgt7Y3/sXdJa8O7W/T/5Vw1E3jYlssgG597hf4xHOsuZsj941xopg/x
GrinJ/kIFwrDyjX6/UCHL0vtzSeQbHvSK2F9I+Y1sJmihgQv/XoyjZFHF4IjqQC+
gw8ryeLAkAqt8w7UOKVDlPDXQUxr9h1K1r/G3GJh2+CFimEQ8d0BGf/0F6PjVz82
utTuR2eKRboo26a3vKQohQvfE/A8LeJkbQR3QG4Aao6hxY0Zj4gxb6i2HrwpIVUO
NfDEq/cT9n6vi4Tz+WgwY3PRBNsW47zGVw/2LATrntoXYTk+pmgwM5medwP3TV/d
I2uhIW5rPH2AfcodM4MD9Sm0uiZvj22Q0hV0+hlXc+em+8F45I8OOxx5JLE73ng/
L/jwHSUeOPlrxTSwEoR+N2QJ9+peeioT8ExYEOnBuwojnfMGBTOjNhfmZSeNtQBg
AEpD3fXb2CKHg8mje93LwM87adz32BOZ2AtR8SP8dn4/HCe2G7iYUoB4vjZL4q9+
Yc1U/kk3uPLdtFRcx3j+/q3HcixTrhHpetPDmXLIpF10HJRIuW1g75nvdMjUGHsq
IfvobD0HQ1DyyeBQ7TX1SYW6KFOBd1rbrv+AeioyeUb0ehuYXCkvzW85v2RMIWXk
S3m3thvBBe1yaQueGBUD/H8DprYJKaCwlYPIcUvG454pp9qW3x+AeBPS2ebmusHj
RgcNIDGFHszN9V4fah52LNuzNto2SnfFOBAlQnsfDYmZBn3mOUieFrM0L58/w2RA
w07wHRaLoY8nDjkdm2o9BZEx0maIYJwHrVhCdnQOzyEgbSuj28gyHpKq0Yn0YeNk
YL1yfvpN6TOlBC+JkmWS/fHBOAvrwuVEaqW/eqJaEJJP+l65Lw+6bGPPjQOMFteS
vjp3RWz2ynMg4uK+qSbj5Jf2Jm5WknuujSmyQz+wZ0h1XncT2JwkvfUWrNRUWp7V
paK0dt2sDbbMhZ8xG3DGMQToxquwhKrA684HFHj2tsOK60X0p4e4OikIwRHGV01y
dlJqJftfjbc7MOqERniDqyRaunQWLF0W2H1T85TpE1OE8jymfMfwoUAzSbnw5k1W
CAK5hzOtwNDpbEIOE3OtesDIK8KUyrPZwk6qt8YjaJ8zgMatqaSAu3wnAHfrlYpQ
0X3Tm+B+2Pqko48jh1IxODeqSbp9LfuPLysAH76JFBI9b42p5dSt3wM7NQg/7SJ8
StFvWwfjjLgF5bs9CcdlG+/FoGGl7vwxjMVoRc5EBn4jQwFZejZcy7RNBpQ1fgfR
H5ipL++AiExWS7XpQhqnryh7x9bPpqyVzRFtag5MfFYGdU6YJTOmXHy4VI+zlKGI
yUs4FbJvVAGG07bxaQK/MhSQOANXo4Onzk7dDFNTsmqQdTZmRclHx+/njV1ui4ae
wd5IM9mp371wqoQIWtgiQtJd9Dty3BKgKzL5mqI+Gm5b5+CQZZkX163c0zTphuUx
sXygsDfVslmM+g5JEKPKQeQ+lC2c/em3Q00Q9oL8Ge+tSXs9+lWcHx0ptPR67V6Q
lcgim2htx7iogo/5oomfrt9LLvgZ+yqiQLQEutjsQKu7gfQz3mRWY9u1TPR5x6qh
nhFJw9eXyZxV/vehCieurlA1lYCrtzrcuMZdOALCiGpWV808cIxbgmJ56fBJM5x6
tAYnm9vMFkR1BSVCNXlTt8YtR1a7/HHCWwz6eCppshkGx7Gio9SwXKC6os/+C7Us
VTid9A0nATL5xdpqNa1re1hCUonEGPYDdCuFk4/Lk0zAThWHw2AK8BIoo3lIEBEU
e66mq9smAsgHlP6EBQfKpmctOKYHpjky6zq+UoV8m3YImWeqprpNYVbsOixfDxut
loM2kBOwZwowjU0Z9W3IO312hKabvjo2vVy/6tq/eUCaf3pjtQb4HOhwKHuOw8tF
W6cS5L8x9L0DihEUf17jIKLST1IjUBBYkwdUZPPYTZrIEDh+3qzZCQCneU6KMxMQ
s9K0zr4oiJPTOXTnI3WiTXUO2dkXJkL5FdGj+rVtwUpxIFObJLjDy4E6IdQ1N+o8
+goG2aCEYC9gbzSrWifH3SfFmEpkFe1qPHgnoNeLX3zKq/gJgGYwsKd5RfBsbtDT
uj1hj9glk/PiIDmo3KwqhM3gxILSmUR6zM/dXph8otZdnDlvjtcUTpQjzegOO3Er
cPYdt36KWLcOWqeV+H+ui768AOiZSTtZ6LSs6KuctKQPAqIduFnVCDf7rfua31J2
gcrJGyR35HKbojrnGFqetSeCS3Vrf/RwUeLn3wjFhJeIAmcst2/tLbt68474gua1
ypq+GDNli49xW7IzRBjOsG9ENQz/wZTSNVGIn4BIQ2It2Y3ylMuz+duKKFPWwkOo
qmo3jicErwoReuo2xpzm+1fiU/2RDPnDVQURZZD/a2bnxqnKPnY3Si8aKdc7ITnW
IKVrHfuEobjRU3mmRXcmB3uUDKVnkpIMOgWrl4Nr9HdMKRkg5tBlW73SZceo0Zzx
rPaKlTEwN07cUTix9SvfGagr0Ts4IBBqphT21jc630WXMNrdlRVGpO85kunUR97u
jydaf2D5H3jZNjLGhUIopdWKbp1MfOkXk0BrmLjzV7cnXBp0hLCCGfdX1SDHJvtu
miLVrHEDZvtdfuNESWoZmPz3AdVItNahyOW6pRsy8J3yJW8N0ZkQ4uR4REg/9V4e
/ZSBRVS6uFm1mieC49k6OCCpnsNY1PLMi30XQHa8goB+P9KcMzCHPaaAQd9p/gJN
mKegY4YdV8i/by34f4ibfVWP8324Pgq3HBN+kJS/6Vyam0Y0VnfkugwZmXQzKo8P
kOG9+SlxekkaBvOYGbU1M+Z6AhCdzHotTetvmHnindvDXHU1pzR3QF4sleWE8VON
jM1Yv6yTtA4jAchtN5LgmSdUTBhNbztW6cLmU84+aAP2VfbEa2xrBQXUbNMlO+z4
aZzzH9+FBwMW6WWkAC/wei0Msxx4ZdQI3YWBZtaOQTwaHxIVgJlHc9DJB/j8XtX6
UnbBw/WEPIYeZkjFiijlyOOrzYN7AzD7CtWlL3pfrXDYDuLHkf1Ic9j+o47fFbrn
fD94mDLRxVJicMgg4I6SxbvHssXiKTXQimAXfPPsxtwlNJAqwWSG8qWB5RsszNS9
Oy95xh6YTvvxFz7HgvKsnqUHxJohmrYHrJEjelyM87knjZ6ZdRhNII+7/3+H7eor
9Yl8xsU/hMUOxUD+lvv9lC6fAoQgS5+2ppIoDq93Rl6pSwGZqN5lh34YTNvaTEgO
fL2Cc2dxu5unoKyIoqkuRKznfmMtVdBvy6rjqh1NjhTHiVCjLMGljh4mSPJVOvD3
BBS+h4XELyOu7rtgXVNvDOqHkhoZsmGqWLPe0rMI8a/I4CL5cg1DCdwmSny0IJRa
sBuZER78wDukwIKk3Yi2je0d1tBP8Xu5VVpSU9o0e1aYZXQDmG/Boqk+m4kk2SsN
00LIRGkudozgAS5DquAxNwHqPz+HrhBSqNfDrL/stVf/Y+253PlYKNd3XYDinmBO
LwCVr4dDwwzaASe503lMX7g8IcjsTwAPky+tYTsnn1EXJNKr3koOohTNgm1u9Kyl
QjL35LWFDn17PZ6sTUck4l6DIRo3ExjCc8IHH0Q1xeWX4Z7GkYwrYdg98kwtv9q0
OxvQCYtykg96Fi+uvIiA5nmh9CSTZWf6pqhzPV8sFGcy+vrkSYZ98+WfwSoxgluD
qJ/24Tze3j9A5e/vGlcdOwcnFIRsVPHU0FeIcYqMqs6xsgc5tlIa+amEgCvP7zt/
VsQMxCGH6xoUE9frHJpVDrgyiDWTUfH9EgnuQkeMYjfllG218gN/Cvo7kCXxdkQX
cqB6xasOsubFWNES2ZmTYJQrpUJgxMQnncJyix72pxuxMJtmelZqPin6LTHEskj2
W1srOszwtu/zge2JTrqGsVWMG0p/Kapv0ry6gOZyT9+XfrNNabKur6llP/SXJKFf
A8CdsjGGa84TghGlW07Gqs7pL78qW0z7OcFhjR90pBiCpFTu2FOxcKmCVq+FV4VV
j3nY2JavXTo4Quqtxf6/gBMCTvn5JWxC+NXBP7uk5kx2x2x8NOpdqR+l1HW9xOkA
On1M5+eOUkrBPPKt2eZkFYCYk2excEK5P88I/KEInASm/kQcycWiUYF852MLaHYa
nfXNNkgQuwtb+1iJ7yadqONPhba9CdPZBPN4sAGdxto0teOstdcaGxc+okRWMtsV
gSLBFbV5nwWW8Su63wotRPBS8NU6zg5e5SHTFhntGk6mygjaXqFzQeeQEktCCV12
xrf8rvEr9CK3+ykXrL/3YlkmFHj9ePXeqvJ17jihwGRmWvAXOpAz1MXdfZjvdbJS
as742OLPoVVhSd8hK7/3W2mdlL/AmL9wdp4/jIegaPtz3YAhCv810XxlGwRxv/7V
4WeZszaUQ/nesSd5xzU/OUsf5LZhkKkNfQ7JxpKicZbvx1I/Mq5L9Sh+gU2a27DG
kyr0z7GBlZQv91+KJ7UwMo8EQ3/nXa2Y40MiBtsn3lH+hZYhkwB10xI+5X8tQPkc
Oz62alWCrlzfJ2pDUUmcRX9gw6GqQ16c8oGHdQ8YCozc5coPMyxbzcL2dJpT/EWg
tqHi54JT0DN5BnEVfw66qfShPamYy4cTEn9RGSoK9xNJhK4ROC1pFlQ9Z8NULi+O
wzINxZAO59beOdTaocDBvsY3zoLpmrtTqNCuMGBOGOj6kK8oVRPwKyL+1co55Ve6
x7+h3pjkCW1W4RWm+jnWEbpEaj2Hw9vI+JtWMPqJkyx0ZWa518wUsRI2WL8iSytc
K7ft1YdapLIPCKHSPt3tEO1k10CTV2v9xV9WXt3EPuSzMu3MQLn+DIf/St9FqAP9
hjd3rUZWS6K63tShaYlgOnuDM09bTuCwWhnA7AgXr4TR9zIU4YQjAi748uBjQ81M
yekXBTEuNtsib00rJOYJDlRHMyMWHhjPxneUubRYVVN6THWpuzASGpP6TkpD0D1N
GdGx7rASC9Dxz4TgoahoBgQn6d7rLSArIgfORSFTL79sjBMoBvd8WrzlfKLRDRPL
5cu4uBRdWL923H/Sib2Eveg1uP1VbyQPmhc7JO6nb0sir22ogvHSTY6iWF7Qqy5m
GHbrAHuzzI49GiS4fNawX9CdApYSz2TxseRPYMe6DvCihzBPtIlpHq7Sa7Fc1Stx
64R+tTP5Cvd8+2hjhvOAl1bZEAHOgbGAOBTIsaeIYS8vkRIt7FkU2tImBUpoNywf
XrC4yAMx5tvsu7MTE+JR9ZNNtE/D/epuyDSC2RA+5MoCwIjDiCyNz6xdbpOwsd5P
Ou7cXjbKBdyxtqayOozqrWVu7X45Mqb6Vx9zZViJW739FFfolkDe/GZbxCCBCPy4
PWwDCf0uD9Vf8xoMJAzhYNxJdN6wKm2mca1LKhlEfj0U7jFVLMEmbk1JHaLnEwnq
UMpi5ekhfaBUeaY5AbYOcAor1KkSbF86jxVc3PBySLdXhUtZio+213U2Dw23pf4g
Iyt0l0yXzfIU4C/4fEXVSJx2Yq5s1Lpfmmcl1ATXgWgWaefigGiKm/uVdgxWHjtN
JiWP70dzPjyfd3zTuQGg6cANzDorJdJ80iBtmaWHbcuXuPWJhJWPzitiuSVFNj3L
Uuc8yqJ9Swjjv6eqr+mQyrTYYoQK+rI+mGoTb5PgwdTJ8/IhZ46dkIAErq2wIFX7
yGVhpnx0vTPhrqWeTsBcR/GL/EJyW4tESSxSXkvjKtEd956hzeNZq54RgJfTt5bT
SADDWxeyNLhboM1EUs8kYjRB+iMoYtchpeRXWLQxdX/prhzH1kx574JdsEl137p3
iVR+dxQy1TcheGJIIpveqfHyuFrx5NLKe1SXJKZAWomPA6VKKdPOv5+sbLa6YJaX
WtVA/lxOpcGRHBlzIwWJSxJfeXJrXuepvoSe1cklpVrMluZJfGOBUTr2tIME5OJ9
upOWNtleuDnvijeAh6DVsZjc8NAmVKEZyL0zenBCp1JOGDo9LisrX/WLZ6rVbP4l
cot8bN2kRVC8tTMb5s4iwIUl9wvtB7VbYibXru34cYW5Y1uL1DpaPc8V6UIibmDZ
g7/sIqzDFLCbvTHe+P2OtPb23qoHA3VqVTLQ+H+06hOn1UXrf9tGtUvPPDlWN/Wo
x+3d9gsmVqFGAarscDq29Z2iWKqz79wNbR0sbGKliOnr+NDSgrZfjn7xyRxk4/ae
Dh+B/Uecyol/qmtBhvEoJkQTqvaX0v6XURsYLPY0IYImTcRxySzT5Nj9kBFmmimy
Cl2GktmIIo+nmciW5NhfQVaiIuBRWD/NDiPzQpr6047+WgXtfkOyJ63EuccFozPe
WoFwp9hHB/4zEnD9nG28JaNKf3nqxy1zEe1R2zOHbHFq8RbSdJxRdBlnXvn98Ycj
jXFjDwf1uobJAJFfAVrqAnq/mQ6v+RARnaEc5y/2fuPA3NQE5ShqaiM4KLBQjf7x
wek1/SS+35mYZRwNPYDhaEDj7SFiEC8RE+op3usR5ql4X1G/ErOwkkTGUxunCgEu
7WkCXo2ojGf/Vc3CkuTBZXBeR33ghMgPve8VA0pnGi8ZeGrFkGiuu05ZkR0/kwh2
CMXOGmIvpmUwwfW+riDhyOEjAW9MnGGhZ2IICAbtccxpEOhT+bfLph+WYjzNRe/c
wu/K7xJvftZxGee/DzBvMdVq1a5l3Q2eBauRnYT3ebZxVhAtHIqu5YIc+dzKKgcI
6HCy9beAkroVOPZgV8CJEoaAZ/K9kp0shtwIyOKHzFoWYduxsoKceSe5XfOFo2uY
25/9MYCsOhky/fsbYl1ARptR5Y2Dq4TFYrSk8L5/mwqXBYgG0+JHUShYLwddZX6d
X7q36cgdyujB2sTZ1mhl74Lu3LSbmWL3UqZQ3GAmKs/RsdwEtqP6hD3dfhf05jpC
eMnWlzMX349IF6ZGHJyR6lQaTLskKRjAYLnefWlPs1nTsW+cBYLQ/HjJZvHJROGf
jhkVzye2dNDH4ebwLouIdkbcDrWf01eg26i/VanCUkeWxC0719d4IsumeBPt1kbI
fzpEPRzAHgDTXq9q4NmZb1mY+ZPkvXT+r3B9k+Fo3MhKrL68svytx2vYB+Mtm0WY
jFp9ybmqpzlA5TjTY+RqMJMWU/M6Nc+mPi6MwVsKw19f55RGMLmuS8V1z+Fzr95i
EDXKipdhUfzzHgaAQjocVA==
`protect END_PROTECTED
