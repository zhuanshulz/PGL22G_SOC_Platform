`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8jkyxF2zEeSaW3Vejs6T0Q8JbCuX/iHoud6goNKPFtJ443qQqLFctPfLE3k+4hpe
r6tD15dr5CXEe0QY1GTcZdi33WjUQq7FvV1e0oMxnjyxPYjRdkt1QC11V0yMEnK7
ylotHMg72d24skONcxg6n9IKQ4YzX6YpqxMPxlXzjlFVSYfrTyKvCzIXKHtwExmO
k8h7c9PyvK4onLOj0Pup5pE+n5i/biFebuNZIEKZWHbgVhFdyVx1TFIVEozWDek8
Uvy+55LXRHkO0ftubwxedLpYYP3rl6UKEztG+REtBQroVGYCPHVdiH3tH4qvWggA
cNY9pibtgIDYuq0SCzAs4BlLxS6J6aG1D/4+mortRkscXgDYOYXcXSna2MZwJYJo
tr6JAZexP4ZfSpyTMewaaSKRYkU7/T7xFMsf8vAJZmMj7dzMmh3UfaCqid4X8J9L
UyfQtQz1uWFvap1jkEeM4KJiq5HNlufFgqu6QSNMXh+vmoPhjkMpYNKNfiQobjXN
w+TQKkWjCLqyo99WaE6qO7eMCN2r/EwfiuMo9Ry8NUrwCOf/4MuEVn7OhBAq6eX5
xyAyWKGn0e2k7XbdLxX7cmb8ssK4lHobG3DUi7TzdnmUnVOqu8lnYsihPaL+icSS
+uejGgOzGigwe1yprpf/beLjKJ8bSE4lki2Rg9h2hrdp6n1+KUcsO4mWbNiq59je
YFpC6TmH0r2QGb2do7ypweshwC8FkARvypG3laTEhLL/oSr1D2senH/VCulU84Z8
+7rvCF/VAhlC2RFtiw5qrHu+gQWSk0NBcPfFVv1CpRA62V4v0CDp3kRenW9pv84v
VZHsAUTcZajp7+62KfGKHYelZdKWKLYkrB7/hcBXPRfLobsHmFAq+sO/HbIpsDc2
pOLtVk939ot/6WfVS0i3tXl0CGttjwX9Cj5o1T4RlFKJH2ilVWbbyih6aC5ks0n9
NSpcKyNni1eIaQ6fVSEfX39jAaLhCwsOhg1ClNNyJuCeXktHQNgL3f94x+vxiQqU
DXVEiRlbU3Y+tDVh1VyVf50L2UB5vvnh0IGcftEMiN3Q5R3MXHqCVmy8/m7LXQTB
I/DQo2IFLQtOJV4USf+JZQMSOxhdVG4VwOTjvZ+9XzP9U/4yfbz1gIVb/lqW1g7k
xWReE/FIplvATgCeP5S0YPFs/bRHOItWYeP/b9o7zzaqyJuLbJgoNLfw7ZFCX2T9
lVgtWV9PjX6LltvKh6uG78p6LE84VA8TJMVFg1JL2YcppEe5OAikPNp5fwWAbbsi
8Lnl3559KSKZwH5xJjILZA==
`protect END_PROTECTED
