`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JkOpYsuUDN/UC34SUdudc3cvk262KFWkJiTxJGKDVbnaxuXM8pbuY2dk2+/aj8fo
qirrvuVeyyB08aiDagc9AzbsSf1provi/x7RGHVcoF/19EZGicsxRasgDg90iygG
bWIT064I1WfSouJDn2aUNpV5TTX6RKmANSuks0OqiErI9DnFBUvhM5GmrlXcSu8y
eqFYvN72gHS8oL+E5Dn6qzuiGKNuxEOAGtTsLkKxl7kD2OHXTIi/mxzD8a0oceXa
2GwolTunhvBOtjdqbsORZw==
`protect END_PROTECTED
