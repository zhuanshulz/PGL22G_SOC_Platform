`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E1v/e0Czq/s36Gqix0XDBoaZG4Lda5AKXmcGCGEtfU9KK6rgDXn759uQ18a72NBy
aHKaIa23cvx4P/d9r+Z7zs+pRUqmapGud+idjHCL+T80pKx0h+9y1+Q2N77f3JB5
WtdGJQX1WTNdwg7BrF1fe1WpLvaIDV2X/ThZ+rPpIBQsQ9F25aeJU8AjlbE1s9Qz
0VCKzyrJeqO0V1XMnGebM92cZ99CXWOnOR9UdmXTEdb8lBDqkvhWcEYDbNfYf0Sl
AhXuR/wiOHmOENr7LX8xBwxn4mLhUjNq+RpbLJxyvXlyNW0IMNgvE8DJ6CDIJHWE
Y1vW1RZdlA2wRnDFo8Gfv30yS+cF7FPJA2BZVncacRVCnVfQDvaQYiRN7xHvL/Yv
sFZ2/J6XrEpOXRjtK/CZdNKKO14QVO/g/x4mPJVxbznTNC5dJkaxvsJtFbZ+4Xkj
00VGmELA7hdf6+H1LJ05ZAE6RW/Q/NJJyHRIwHuhyWyB5kf8/6whZigqk9wl+Ugx
ughuy+ZwS7nq22lClbHX82qoan3ppGtn1s2mZ6NMvOBx6TJM/yayqXq6hgcsEUFE
085c6JU9qKiJwGskC2CWRbSpLKgtu05jKRffjMNN/rCyex+ur1PlHC8UrH/NC1Yu
JXAv2KIRiLZnPM3oHhyWIa3Qakghf8xTfA0vxpYkhm+tfGuIWY/oJ7ydbtVPYgNw
5w25Qq0FN/5fAQH1dcvEje75Nr+Uz3UJlMeuZ9ET80t2e7w+mQ2CFCsGJ3tQUnht
ci1/QC9PMDV2IZogfeu0uWIxO9CDQJCoUZoRXj7pZr2OSxYl97PxSpBsQXud+ndN
/EFVx9U1g4sBFCw12p1iUB7KM7aZFoSK6+h+qECwWMqEAtImfMspqMI01wOuM2YX
WZjzBpr64LPdKXZ21DPBlI4caJvQLm50/P1ShqqXAC34VmB13xMyH5a+02l8qeLG
Majhgyw1+q1m6qHxzVxUoNVnZXXwmgcZNAtMD9CLfVUqULlRg8qE01HdIXMVCpYH
M+4NIqCrLLwCCa6t80sP82sJn5NvrOyJt6SaK3u4iE5gePJYm1YWo+YOojw9/usW
EJyiATVNtn/0K2AGtwGoYn/DbAZuj10yQEsxLloOU2HuY2DIHUK9uDkmNEvCkthl
DjghPkZJ2AsfmeYwDTlovCXn2Nf7kozb37hWf060I6+k8NBcLnU5FvE3ZQNc5VBL
QewPG/rQRrzOKH8HBfqMdynG0n2P9xBKiFg4M2Qsp5RKF53+Jh6KjPUcOrZLFz8a
3oB0HFCK65WKqAZHw+IsfAnGrnSRBERSs+J9/T9KNxzowvAez31Sp+ioo1yGCAfM
yc478+xtq/KcJiTEY1q6o0CC8GUaK0NaeYpOG/TEoxZAR68rVoHw/nS0SAeqJMej
oqte+3AUiRnHTW+KkcXIoQZh6Jd9vBDG0kdB9YpqXYewnM2ajEkzWuGceCm4VJYk
jj0UCDjjE2T+rkEfsqWs1MACoXElt4/wQmiybXXsstdTU9MmP2E6CRwoh8RS1eXx
aiVcvlfNW45shkZZlXAnytjKEr7lgHQJgpsnY5srQW5FETfZqcM5jRliFamG81m4
fmHS9oYJV2yBhKYd4J3c4RSAf7iAfgM3ZfGTlrSmV20C6qc7Cmoa7+2T3nx2uYWb
AGhd+BVXoAQBsGyjHXJn3VIKJhpnd/LheQOFPyX+0fV8ZvcRmlOryN7s4vFhCV+E
uKDZq7mdBBQIknbXsGk1TudSv3dtXelUhJufzgL2qX3r/ny/D92I2mesgkavgFN7
23JmiLZpwMG+gY56Cp/rCx34tbnLxATYyvELFoAataEbZVZTMyVzgpMplWLjmm7F
jNcntzt4V+ModxU2gVYpC4CA8KFL/PkA+kq2N0IZ0/tW28yszaG0I5n82xfG9u7B
e9UKg2d11FRh6BbBF6oG8sOWA9S3WH+o07TtThJ2VHvbrGANhb+smKVyckKGqvIu
6x1uJE8y8wOCaFFw4/0WYb5tnJ4tOH8cNwKPU6SfisGfveTuKXVcOBP9uQl1Bh4N
rjkPrxclft2ibrnhkhoKNitZFbUeJIorCL9tPUxJRIwpEEL4b6h/IJ42HVd3k+R0
3vswTqoTetpjmsXyGYdsRWSymPYvMI+RmyUsTSBkISsyaP5e9ydeikDg0tgcrxDv
AsCxrwxPaBjY0pl2jyhrlBEA6XZy7C0FcPGgIGtJlP791SHYLWDXeo+KFwA55fX5
P3DBk2MZNIkrVg5MENBq8imzk+H3jBmz4fNDUUy1zouZDaRUVn8IpVAnt+fVhEdi
iLhVDgXIGGaseASiMfvVzs6iSveY9Of9V9M9vqgmd4kMvlxUnOnXZXptQgXuw4jD
h0kCf5hzBj8FPZI+EH/G3kYk6awEgsyybtrvqJ2HCcV8jQ46GXlQYOJYPkiecbUz
YEUQfdeQN051ICewWLcCGTXz8kYUn8kcv02BN8wRjsYYv8sdlDHPXUN4ll3bNs08
Pcr8OGcRKPSOZEfhXyarm+sxwtML6/ckKYILBN33F8NtLFBKz2yh+R5vhHBYOqX+
6vXXMu6J3cvZDXSyHGzg7XoPuPK5hhHLWG2yQsep8jBdaPHtoh0MMugsA6n571Gp
9pzHjNOlyUWcixNkGl2SzyBW/wN+zZjG8sEZNgDF/S4HV+yBlhJuyZfbDmLrtSxm
tjJK9N7EBta+4ef5yRcOUSfNQCMnRHCG9HfqlHljhttMZKYGD79aN0F15hvuGP63
bJ4RXFln4sEz2bgk4MXfF7m4ni7NHF+tJIyYLE8oUhjnKTY3TImbcrjfCJFwA4DR
A5UXHbeuvC2JyaQqmGYJzg3GUFvfXZOAkM+vUeX8+sKoQt3rhP7O7r+ftMxU0fZK
pkyGffzpIDmB0Fk33BFjs/LypfhKgOd2SpwvB/d3hl/P4mf9IXMhyaBFEFt8N0iU
okPDqTsAX+atzZ7dnZVjr6Z65JjbNME2a7mHSTL4ZPSY+giO1vte+ygwu3yNde/p
502G9ac/78HBDJU4crq1gPWztmH0ZWPmgbh85j4LtHmv4zXijY5XHBpf4pzX6nhd
eKrpC2KcR49/L9EBKg0P2BaCy3DRfYa88yQT5ywq5jopYaHs90BYxlWQKDYUXJd+
W25tLRZfCHazpyFpOfqkDlWPpNTJJrPedEAKCLfHKw1IwHeOZi8bf0U3UoUjc5Z8
hFEsjx5htwzTCchXegVyRaM1P7OGUkcbFG7UzR62KiwpBi5qV6uPCOpqOxUh0DaX
8T8xFWjygl74eNx5ZO1h1hqeg5xBKTaAGY4G4wc9FG2lvlQHC6G+/pFfyDAFw46A
lIMaG4aKZL1h8tcSqV/+dD+59s46vk3jiP40S6psFb+JD8jZCuS/HeSKzCDm5cyZ
e9CRaSoLCgwTyOd0GaS4Lc0M2VbuzYfDQZz34YrWeY/b/C/l26bb61wqvoSva0fI
yXVko55zkHp+qeqanJdpXX6Kch9KXrXWxcekdhp2V/mYGkRuq9WP30bFfiXpJF+X
HoBZ7qVDgKk9SpnUV1sZyyvLb83CWMwjkamEIySZUlAaFMdEhX4gq3Mt/XFbHH2A
Jc1c9rKB/YFl6QN8CGKU6g==
`protect END_PROTECTED
