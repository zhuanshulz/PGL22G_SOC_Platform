`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oc8m6saj3nUadNYjKmdOVEb3nPBwOdx/Z1z+l3Ap8CfVx4YusBRK2vWV2QeIGgHq
orOOvGzjB7Tk0hNGG88sgv46asjA5fg4LjL3BlnzitbIfjoO5WWQICXmJ5CLqgjo
GY9DaQ7mD8lvMHM3D2HjqT03PVI9zR1bzKYyhDaOd/3C4zxf6GfWNDvYNVO7KGJV
lH3AIXK1fcwEonRVrO4RJl91U6m758NqO4ERcbpLf+bgyqphq4I4572W4ptIwTXC
x/CE9HmEYkIqllByPiFlFoSUGCe0DVQd7oXArHiF0kRsSYVa0gb6T2edgA2AerQe
YF/nvrdlwvBOHv74jj3eibCEnY3y+zequiZ0ZxwTybZNDiMp78xmZTOEytNnEWr+
HnnSiKztn49vsxVV1OIhYeTMLqm8rbxz/3vPDA1yvGwvEPQcxRroS+ObilL1J3J2
AO0uhTiHgR7v2d5Vkh0wxWYpf9RArqFyUwciriunCdeXCzQLBx9OQSSc++jkfrgl
BE4gDMwEx6+lG6t3hsKgGTShy8U2kED5c0envpAUKOxpChgdqreFnXCjdrctogtk
UreRWj56IWDQWcjvn9PWekOlCc5c9h8iaNDGBf/hXvq3E544TUAbnVtTPqfezEOw
U8EFUGaVyMCvW+Mm9dxFjmLI9rhevAR8xjXslIsW5MvjkhB2rJjZ2piVNls1kXB3
n2MoHHnyJk4/iTmfC9qVk742rPZC2mqLL5LvqAEBH9O1GmOLdDefwILjUy6K7/Ge
CtuCsYvhLX9ra9V1e4iTX33CU6Jaf9PUkSpvxG7NiCO5T/FLgs5KtX0r1za6y6ak
ba81/CrEIPmh/9lLdvEze1jpvxctXEV1/4a5fq6rIdj0wiJlgRG0Qp40MC1kL4br
VThpVBc+vPwFi6PQ7WwLXtQS9GX77d7kuBqZYo2XC9m8X9Y4hoKxKHYHes7WobIv
Rgo410XBMCIZTRXoKnkq2siJdCuy1kLY4pZDjS4PHaue1dapXqQWAOgk/znmcwzp
sdO61dhQyst/RhMvMrtBrOjDiz95NWOalmM8lkKQvQUse6zBvygx3A7XQFL0SuXZ
mY6rS5JGV4Vc95irTdejzLQf2T0T+YIWe/zVOpW+JTWauVbg5c2GGnbiqTOnfSOt
hlkyRyeHetkWG/lzXVSfziict13ZXVonJmaWTpGbQmcD2Lw+GenGth0DvmWeL4DL
fyFaqZpTa6aiK7Yn630377KTD6fEjq8dKdp1byxIrUHP/kaJ07HAJQfayDsym4W0
WlB5fKXKth9S2e8+uDx5+hbwzW7VPr40nAgFmtKJ+DEzAwgID2moIDDPVVHiGqkF
+jX0YQZG6LQ/K/sL7DSYC/gfEodd3YuHZ3lwPmiATTUtyMFsAWDFizA+wppfUafq
61FosgNC7DYMyGztUmOSVD+zE7Kqev1+MO3B8rUOdWNJJZ+A+HOlMxnTxBj2baom
OgIRQIeKKpnXrcl/o26ejg6400WidamqomSiYjc4qmNl9GDQc0fOMWW6Xt864ayE
Y3Y14tDVnyFinY9jnfW91vmD3604WTzmbjSkLQokqxUiytYd35XW6cHEc5yKx7Nh
prFQri9NTXmUiU4q1HMqP7+HbWDLUo0mQBP6oReQNvqrPvMLl8sso2iEEv42kGxp
uum7czthC9DQh0zW4ZbxB9NFTgm/dPWaHDyawKkARrwP3cDYSTFeNks8IMizguVF
ribpT3nRFQy0Gz71RbgTmuK9posGDrgr+ZLCqLhazuECwJ86ZSkKWL7YjMo+xK97
1awpzXybFW5AQ3hW7/PanIFdWRQVrorTZEujBJKwy/kPkhW9QaPZRYUBWQhC2AEP
BJcHd0BP9Jb6fUgtavI9ScHODsQ4IQvtaBB+T0qNR6xRdPLcAqVSuaEOC7D85GST
fvu70LaGh69TTRu+l0EBvVN87usk32LQLPu1qzhozbqaI1hEpGYN8ei7YD0pNCgz
prCFj1wrEGB6eosXO9FQ2X7mUODBHNtzHjWDpHJbtwUB7tT8v/ZYzhHRNlE3bIVz
fKOw6DtO1QV9LVpbbmZlo4+40va7V0xt3q1uqzP14WWH8XP7LZfu6pCX/dBawnQz
h0tVjfmn+ri9at/ICE36u7MRkMC8hdbix93kVLEIQGjf0M8a0UtiHipnbyCREVX7
Np8Xn+IM60N2gq8f88YnhSEe9G5siUrP5m1MHjC6uH+tJC8xg4kYm0C9yMoASei0
8ZPQ76JDaq4dwjYBNc8CNjIDycjxDYK1OTnJ4fShVKaqLV7r4MsiCwSWddjNrbei
aKWtt2nxLwNEVL06a2KWtCcse2xfghETYYRhcPv2wZQurpzXHKvgozyOqEP8ROC2
/AvrJLpRR9+8ymVV6yFUK/EYnV1aer00uM+0m9kxTyCE2AM5ND2mNYDVMC/LWDu7
K6Oubl4aTUr+2fquMTF8q3IbX09e+BKS/tkN2wMszd8uZIibBEgDNFWPS5AMI/Ls
j2b+KBYxCgI9BLBZAupn1srxI8GJnwybBhtYJg5t2Sv74Xr7ZN2ibVOnBNbmHqXE
fX6rC5j1M7zVbYyGGQaPbGGI3UO5NGhXdoonUIKdzx6F39KhGR3emY86zoWQ/bV8
97QSftKnUaJ00Jh0KT1NOPybPC+49aedSm2apdNsBtbJWq9dbthLne0oF4xeIvBk
HHnQCWtv/hwJ1z4YKyDT0iWujMTQzl7cKcrjBHQTEbrGEP58nasXHVTpRhniCBHW
nyPmfhfBfPOFtbr1uQDo0P5x0ok4eE6u0tmMHbn0Zq0AmicORg0VAg8eHSINJcET
ELL6UgAlY5rBIW2ONiXuGBEFIpM7z7rOz1Z/9q1pvVm+PUINzXuZJFdm7yy9eMcB
YJ7PKFdmM4+UIVaIqMx1MkOFg7jKte69LAWl0Ae0FZ76GuDYLbOsSNomDh6ivVT1
pdpfLrzHyjhtW6R47TiEVlZv9muGfkgkf3Lroy4FoeAig9fqSn1ayu2oM1keRucz
IJMEUiDHFMaf0wMZN5uC61CyqQjpFPiplnbwVqI7/6bb6B7oEOG6KazEYtfZpNIP
JRIddq/0zLAtEm5Z6Jgy77EqY9JIAOukoFkjsSx//K+mogLcvZRh0TmuOmpEtw1l
GhBr7b1lxPuY/srO67sM/Mg78gRAE5SlFQTZPYTsHw1x4c6sTmpcZS4EThnTXel/
YUGW+4hNXEejwOXcrwKTY1HSajiLMGLSNoDifNkBkr6+779sRc1+j2V7xHBWQRXm
lralZEUczpbWkUTvqVqiviqtQ4CGuZJRkjQHccLIXT30122efOgZNl4/V6j9gFsh
Fq07jM5wNdHzRcNi2o28OpTg1f2Oa9/4dkFkXwjNKZT74edQy37Svb7STCfKTR2i
7wpe4irvhOrLPHJj5SLFVKm6GeOHGQYUs0QSbKYN/WVnd4IxtWE9sQBxZeFMst2j
DghatSg5cukyjrRbbV1FCsi9E5ySo4wDbKYTwkYFp7A4RGwno7v72NjehhEi7ZNb
OB+sp9V48NIZgE5N8DqUOvo2ZBIWBakxK0gHCn4a7ulKotvmOhQ5V1pxvPU+Jdbu
dqi++1G6Hqkeomt9roq1PVJC0lm4evKCwvDpQ3+RQkfWJcFTj7KmbiEeQnVRGmP5
lRiApjwhf6ZmA9rKtp3KewiiiVxLCz5v3iJb369rDN5HnURy7lHEROhhM2QIKnVg
6/dnlBszlNXfHQWxTxsBiE8PuPLsZdRGcQlZY4XS1MVA7ohz8gJIyveLA96eZbER
rmD4U2xyhDc3xuXQjX5W+kHgAdvi7tgqct7XLNWKoLtOIM4Vs6oSr77bkLCD8NCO
oLhKW32TFFthjnWo7lG2bWxFiAWOvFLtp9KP+P04dv60xc676VI7mdtH3j+P9Tqd
2ZRta2SbT3eDHReLE+HOLyEDUppzgt2rkcIEeLURQ7nP7CeFpn4UP5MHI5JuLLLj
mxEptarDpqb8stc2m3WG1Twf9F/Ut/YBgU9UKFYIjtCTTX7NX6p9SzEpYWcSrcCi
tNXtkEO3f0c7TGPGseZ1iTkcos2XvMY0sY5EMicJtu+IY1PaOxcOtTB1+i2Fujov
rC4CkwvSPrvVC+i2m369t5vt3DH4m7+S/pWuSqrQ+g/uyfZ4hROAJPhcDYuzm8CM
swkUGYf4tQdZN1x1ZEjGSDlGpVud+o1VsW8mhIMjgyPFTtEJYMuywkIdzAkPdhyF
flD8JIch4P9dqhjJxtLztWtusjckAODrOhwbPQk2XcY+b+o8N0DS8jr4V6An1QWj
ntUebstOaZKj74OJnFZAAQRAb8KhIYtxOMbXpVUKYWOW3CSilpreKNLZTFQ+h3b7
kMPVK/7E6rEPZtAX2euB+43B+HCB5pkeyKecPi5JJ9SpL1r/2im7vAFdTJCpDygW
8rGoIhee0LdWDtUGgZbwbFnxH5VneYzoUcrbm3d4yfYv8DgSJK/MqWiLogo0wr2g
yO5bOzEHrJpbwbuyfo4uC55ymAX3Dvv5tkEYg7AInOIgQVyaCzAdoCXbLf6CBTiY
CFPN4wr4TwDO5on5YOIxf71e77BXp3XnUJWJiQEmYr2Bhcd4e4RiTtXXeHKU1QlC
d3We8R1Dk5KY0EMpY7dIRsU1E4frFZewombe8qdqsEFMMHwtmB4ljeJlEc1ZaBg5
Kum+rYP0cM8IHYXmSeEVxsj8B+ImvMga3oG51kt8ZVs+H0+2jIDTSiUW9V/rzARk
1LZih5JIhcj+ESO7U2hFWXuRyzfSAvX4eNxDfuwa8AH6ZtvxGL4ygjZtiWjSaqar
B48jguhIsqRIlsP26pnyM5/R5BK0jhgNAm9tuepiuWyLIFanTrQ+t/OC4AIoZsud
WTjCAnBM7Vp3lGX78dxnWtXSZRLnuks0NPHy48fj5BRbQbFn/Ca2YGrbUMA68bah
sgwB8z5OXxHdHCMlyjHmgHU4z6+w0uTHZM0Cabbg9pnuSkSfRTHpeHt1I8AV0uDO
PlyFHboqy4VtDBvVvzz8FPMXc8Cw5zMm1hZSG/g5R2Jfckv7ahJrdK0WQmte63Wr
S0wIcB6IuyZtTL8DDGTVE6zaIi9i8QN+dlMm6UVhGAbuEkZWFdwUbcXW4qKfD4nX
m/9Om56FFfWIYAkIAoMaHUrWPEOvp0X2K9PavIeGWAoj0nFBTvJxuPVMofQoMd8l
n02tNEcSGY+9ijIhFILFkn4k0bQATM+jHhnSvLZ/Gc3mwZJMzxpu0itpNV2x54UF
YOhKDXc8linUHLp+mVUTaNfPgZBjy4koiToUiLccwsbcTUcHtVY8Pb3LeVrDlNvJ
ei+54Cv9GPkj0ozRVqe4+8/Xk7q4eT7X0nTkle0L2Zi67InZ3xtBLWY3WSbzZbGu
DwW7r6lOCtKzNUOeh+T6nfqHVgtnYX7sFWODbEJlv9gWNRhpj+6o7mGiZcEmzU0+
VDmv6VYMJviMuQcYXi+4rROUHFKLAQEbOiUJEXPK0VtPi4b+9FFCn3lbkufpD2lX
pKDu1+6NAz+ZbB8heuQ6styAmyZ8l4h4HAG1HYHQVnOfca7QXc3t1XynvJs+gafb
hhZe+Uj5encrdjzHiAi775HGvvWDLGehZ4YiYOu8XtA6hCuhyE7LxMAP8F8NjMze
xXETttZeL5Z4SA/6ul99C3S5WTKr+LPQhAyJ2Cb36UMq70B5T/8uAgEynRJY/S48
OCKJYpGaT8ZBSHqc/khljQ2D2STXGO0aEuRVwKekov1LBcM/NF7ih2j8fXtu7rWm
GklLJySGzbqQ2ij8LHIq4eIDs6fZtOQMR/3lHuW4BU89Y/jzRlnN6VM8ozYxcqyH
G9dgpHJu4qzVl8h62LKt6f34EYbg0KGWy1QZd3fwNaWtudsvt9O+7ULsew7syUdp
9iLXqrlKj+MCVU1rYYUqbdC1UZYESTfKUZfvTMsFh+vR9Wl/7jfM4l8caZ9WXahU
AzvAbg7xzZm3kIy1Q6gY132zbQYmJZ5wwu1bC0ZtNZ1yhiTyjG5KR8a5nka+IdMS
FBaUPyYRKlVX6kc4S5zwx5Kr2He2rkmaTd8XMoc8iYlDg9fSWjRFj/Ce6SsxYzq1
TScjezH1Mj9XssLb2Jv5RuE5W2l7vmyYNGDz9ck/FZNi2w+xEogcOgRX0Ao2Gs3u
qL2Xpwk8JxpHsvBYpfMlV95NDg9X6ZF7iFHwiYeUkLAmDk3JIXIOewUEpgb91eJm
aMbZOC0oIseBqgK8/+fY5tDEbeeDXTpga9A8/Es2rPAh+DPqX8rXKkgqmbbj6rBz
qsQDmlrq9IkaqOXC9w4M3AHdGu7BYZSqO9DD+zgj7NKU+Bmz3yQLjyOt9pcfsP5X
XxsnQ1sH2z83NfmOXSLVA/6W79mb7dPsPdLeEDrBuyXl6dDrqYZpQsU5t4lmOxyL
qqMm47pC+IHmosp43B29182FsDYmSHv4J25etd10X1einF3jxlFwXBMTfrB3cSwX
932RrTR+o9YgpZyE+wUwCvWzhJYdoCK+DedzjBQYm2JGRAb0zjUWdFyWBb9RpEAW
u1p7x3JUPlyW0clrfBJEQKCZV3tJmTdWJJ9db6OI7S40LgEkyOYbsdy6qQsYJZsR
lThkzdJeRC8Y0sYcqNXwlSt+VppqC/6ts8fZjhkSq2yMc7ZvasCIn/3cspDontcD
eHC/CNlR0Eto6WuFUsPtrN9ucA4e4eFFFEwmF9mUX7wnn0BWKcFAGVp6nyzcMG07
FLAurCrVkpvkZFAiKxPSHsQ+3e6oct8W8G9Hm3mLiifyoe05tBtM5JV/OmJRFV8f
kcv6N4QBRVTyce5BuAf2BlJ9NYiFJhbmzmqo5b74pP6v9KCyrR0C7F3e2zaypm8y
bbZCrGZNE7Tx5e5v/VFIFkqSzVi3iIoTiOFL+8fNf1l4V5wgrIRr22v51UHDbqM9
aJcauGvnukDxiDKZzkN37yPwdWptWuVCIjar4CR04TeD9XeZHbm20AdrFsh551K7
UJG9qxy/RYj40bBW9Vl+JnDdIyZpsNlFveWDBfWOktIoMxG9xqXI2dZ3UfXwLnWY
6kNRQP3cS8ySYBPXmxnS/gD2caJwa03yFMsLtzlN7LIvHbp6A3l68rEJpquWBowv
QegxmZ7dW1g3s7tALMe7PEZRfNMcf078hHQQDGgPggZB7ng6C7jXCl5etH3XIpIu
z1CqA1dEXyoeWAO5CNIt9lVN257BgdsRxE+sNnrdjBggJb7x+No3RfncZda93IsL
ZqPngggLk5qZ01Qp5BGpC8vawpcWqtTzAPqSvKOKNxhuyX20BYdPErqyrz/ylOtA
OGiETgznDFsD21dB80qv+60R3WH/8u9wHocOq435x/hhBGB8ABukAmywFn4zNYJd
IOv4obn9+Y9+Wg+fafXXa1AsiYhmGxY8kmMMGEccqm9vQPzXvwV9deCraSOMTxib
W7aWVWoDi5hA8GzVuOZm/1pMFJxERP0BZgL/Lufbc2H3Hch5gGDkG0qngjXn6Y0q
9o14AvaOMwUq3eOhB/vSnDh+CuHcpAtKjjQoDXmgfl36aO7bbNDpffmvt4nyR/Cf
nrYGu3+F9BBuqCJsTh77KAC//zTALm1auTrfH8mKPvd4eIP06y71ZY3zeDir4AJf
3pLJXC61ryynTwCU6zsPPFBHE52/CFp4GdTTYSaEpffDfuwMonwQMz/dRyNBl6j7
Txc7iyISRNVmLkC6BHYTSiR8HNR1mVGv7W9no3APSW40JRFxi6c3tfo9UIFmiosH
xoVvXU0Ryb37riXYmf5eTr24v6VQA5YE4HRbpxCUtKRPRSTwfT7j4bszUFdBxC2U
aYOOisLxO3inxjWgPJmMNRxNEtfn5YuxWTe6wVHKIOJWPKJsAxvtbV949mtjToem
RTr6b8Nc6zv+AvTN16UUR4iH3lv/3f34DVK2Vfl3Yz5BWdnEpTIVTv7xRBk/bEur
4CPhwhJlZ3LeDuoG/H7H2vMPjUp48kEhpo+WnXytOpp7KUeQCatWcV/G2KOzKEg/
Bbcxr5+/WTnh99n2UJND0UCdemLgg6unrOJ34g1afALpk2JsyQx0fVTgl8Hpxc+X
HzRUerGgqRcKff+C79+kvsidYhRaIG/32wT4kXs4wadp3HRNtnNJlI+IP5URZlpX
GNUH5KR0luE8sN5XggqCgnmqYHpn9cV2z7daGZ89Y1ponHVuJiABEBIWgH6GxrmD
yAuf1SR26TI9di8HZjw//V8O0/Y+PJP1v6qqOCpsKtmIIwNNx7kK6qJlwd67MMHX
4Q9zhxVwJmwTrbJUQ1ALCDAI8N0GNOVGB/VMkRG8lOyzx/E+2QK96h7fk4YaRNqX
PeaBTMoSpR+1ev+qqWVpBZm93JImf0fgi5ULLKNSxjjlqn8PougukthI5gBEy8Qm
QXmueHLu23+O0ZuB3qRTIgGM3xYEwdayFc7IJ6fRqWLjuUEkVk/1R6GI3mWKSZzu
hWCnz2vSmzFFgLj8+Jd9ZdgPyXckSZ5zpw8yEtIrGVAl6BuTma40AUziyeaUmd+A
io4gweOx2eN+pUAIZIRbKjOWVdpS6Pg0k8O2QKnTiCtkxE8yA/V9bKq7q/zhyRSb
WJw30Atgupa40WsR3ew72GUWkeMkkQ4zazLssLp/4eeWnw0uGNOhikhrFDXYS+mt
gOdkDM9A1Sc2/TIngRgAiT2jswzsFcJHEhcM1y4BjX9SsOgZFWcyfydbKTj0C4ax
LAEJr+RTqB2SxDbChu93/9Nb3FjVYaKQWjK7pZNO3hc/hXy6xDV9kB8bpb8Tlfc/
kuUMG4X+U5dsBqfmsN+YHvHDmm89s9HXFUGfVMHpPHdU7DQtkf/EWNibzYVaH8M3
dif0DsQCUsRhOCFoUTAaoC7urzG1J7PkTx+fodSSo1kKZ6XTCLoYHtyf6YghrkWm
I+8nUvkL0o4UJj82tnS+RQ3E260cikNLsXsRLb7Q0ZX2W34hbvjbNoowQtNV6FYO
sR9v9218mzIoNIOQdBODqxgG3QIRVrsoYDAfXjvSeY/OrgDbCUmBGJSptc3UQNGX
YdRr6lACiNKLNxEc9j4HJb2D+qGvpOv5/Q4jPQV0NyeC764AzimMIEQUhu8EEwwl
zg81qQp88Ba5KpYyY6VdiTBcgdpEjY37snUKdqsh5G37MzKvHg78dZDaNz3ikV+r
diOXnlFSgVnXh0QJZwZbIJdyPdfA14hmiOywwwd/1g+RKjx6rKcZz1ovywRyA7sX
holzXY3C3grN+lDIzAFmlA1bvubqcD5XINo6cXtE1V0msZ3aLNHpjgxGzDt80Mjn
jqsY64+Qx9oEwq5gnhOYqgC7xR38znVeA1dTlObJBvozCuDn8cQgTLrxqKOqlR6V
xKMSHWgTm7+UwiKQRjk03UkRvUGSdljeDNhauFOqy/IQJ6WYliYTDWdyjS3ALiqM
E+jauNIXkl8gFPuqxpFNihIncYQZJqWDR51hlpxI4nfLOBlw9HPJ2Hq38l33H85X
1BmKFlFXuTETTtt9YYk/MgJCcf13B/WrNOuBsCvthuCrnxd7K1YWivEc7Q3UAV8K
WFyppSy6DnjPu9zws93cp8Zh7qknOj8SAcoF0Tc6YezW4aM5DrhP1UgM/GwLWs8k
Bd36TJV9aeNWUnuruKd9lIr+fC3kpvzzIubY7JKa/yhNUx9yPgMUImQ2YDIYCT3N
gspmHowvjh2W9cP0/u6KgLWP5gaJrsPYNNtFXrerHhmSpR/UBS0pxF3914yMkTdW
MrwPAtadqWozK4olqTO+FL9qeekoI9wapz2g3zF95F6EzRLYcqsLtV9UrhJn7M1n
SvdF8Vcv7VcxdtGU7uLC3hzciCsqjWow8mm7rll8V41AcW2YBrVaJ8YB2Gynajee
GtBCLsZdtzO84fhpwsL9DNVpGARFR3iahpZaQe2qyJ5y2jqa8EKRkvsNgxpEZy8F
PasR68cLUoDHukJSnTORJ6h2SaXtAUDKpxQSBn10pNlVimM7Wg0bjRpi6RvIGdlX
n3yhdfBFliP6GhDpZYGB9ZRFc9bSYkOLR5fc2ztAi8d+bPJ+WT9qPVV+cI+JdUd8
+UjLVq1pF40EzK8D8pmHrNtmT/oM2y3taY+OPuaPgmlEuJdySB+6HOwq8xyhQvjW
BE+F4ApUkKclYhILI26gNlU8740vL/JU/3vd4uIVzscpKqF5/j7ltfckGCbhEIAS
BiEAc432f0ARgggwfRnESCSjapUzQhXhCcauuc8PDOV8zmAF7ZXoUiRZzXZzvOxT
z6t6AXrpTJg0DREh2Ku/AYd2xgNQJemSItKeeUXQKOIVvFplXDnA6+yTf5QjARnx
2CJsfaA3gG8sxGhrWTOdQy73uFhTCP/JiBpHhHdnI5eQ7A68jSJPJv7I3I4eAyqP
OQvuTsXUtNKdrxw4VQKVjNa73Gwp6w8jt075bcLc6zsRnAwbgyt+ZTAhaR3k1MbA
Qn7R8BtgNI/gA3EPeNeqrOF92EsIEvVal2eenNZl4IpTe6dy7j5SBnojtMUxnVLF
tlshHk/ZgCLsdl5dsLEB5GrCqzW8HVEohMWrbhIdjxnV9PKXOBoAtAd/iY4OQ6Pq
U2dYjkbAl7AkZ5cwOzweEK5GGVO0xcxRuktDT6w0IIYOTioHK6emOCYQefAafYbT
LERL9aDo9sES3z4+FCr51CuJ0goc3B0TyKfrXrQLj6hWNTIwmbtSaSBZp/dHWJmq
mBJ6Oli1euklO02/Aux34WrSNyUjPmgJTxVtO0BhNrwzGgnD5Pz/cXOBzhMzsPag
e9b2N9oNeui9IRoZ73C73ie1hWLCKo351KxcTl+rG5hRHrgLMI8TEvTpIOTOTwey
cGE+nnYlYXXXT9p1/foARRI0ZZOKkjuL9JMyz2yQCRQScvnekAHgbBxQcHC2UMtW
dQTOKOADD4dkLSsrkGHp7GzLAJ2xS0xI/WzoLT74j//LEgVaHto4Jj74+U9jH9Cp
aba27cQlSgodcnev9iatUmBtd+IOXYoNPIvWl5Tiu0yRFlccrnfyShJiMyI7SYvX
Qx/zaL7QrMixldd1FC2C03bow7g+2k6KogNu2TkSVGHDVzfrQ8LGxfh1KbjIfpPD
FHqmD1q2k7NL2IXKAe8JgE2kBKUfaTSSoNucsdkGOxN5+3OypvcKL9HzjwZ83wKn
t35JWGRm3XoPxCN5QHKcELpbLz2GrPTa7Du7aGYIO8LE1AFukDGjA2iznVVMWLqR
cJPvpqY4BXHSyE3CRgNeaUzuhdDPZvgMucrVbqnizF8VY4tluHax4aaLjXgxtMgM
azo131QrjwyopEX8+/UvTPNF973VObfaFsLcrmS2aUwmbp/sywiPU17euf85Da4N
rm3XOQI8ryuynQ2KphJK8dRvYj5dzJnfqmiYNe43a30dFnoD92HOHiBN1qtvwKdV
o//R66WgqTVKzCwFpfynCmoPQV1T7LdXscUSpZ7DfJIN1x54PXlFku1/ajc9CEF/
xT25yk1F89DjBC6A5NT01oGDISHxj5wL3xwjhBbwtYRdErqhqxrQbi8js8kFbD7a
CkAnItNUTHctWl1kO728DWVrrJNs4bUjT+2f/H65jdFfNce1as8tdZ6//w8qOmBW
7FB8aqUenSFhfN0TdVL0JWTpnEWngu2+mCvvnJ9zLfUBlpYuBTvkDGfUr0/ThA1G
50gOqgxUlHDYCoZg1FT7DO/FsSaCcfIDzKWIOaLzDY3yfquSBh3HoAEWo46qNsof
qi3JxZh/fEuvLCMazJXdzA7nmfNH3X1FATvlOCrRKyeivZ3cjZUS1xsaO43Qx/kP
BRj9cpIFGWJ32K5Ke0wKjbfa5Mky6Jxo9Q1rBb5DLYOauM5y1TTy5Y9AlhOPdf0W
Rz+gWFf2XvSBnowmJucG0VzUgzH/8xBTccylOXmRVjQqXBln9N9Zri2HR2DFn90O
n4mD28NalEsmPBhQDNJgINp3NBZ8zsgoEud9QastB2uGGmYAnBvIMgIWYQza56lQ
t5h1FY3UDehjkZO4g98vYKKV7iRKlVA/mP9YSDW/uHl3YpSK3vIex4dU2MStbErP
Mov1eASq1wOtWB66hgtkgX3ooTp9Pq0vQKDq7NRFShdvnXub8NyTsT5c4rojfb2Y
K/JG7ofJWLmuTDbJlUJvFmLZ59iLjCzMG+VzNsB473NFVlMVD5tlFnZXpkFtPFIX
WyBG4Acj+3Rr4/lVOGgZI7agoAuDffb8QJLQy6nci1JxhLmNUvI1TMNPhLfNzxhU
l01UmossFkhZtbJj7fS+c7frp/I+H7N8k+REF0ry2QEFcFx03vb+uUr06kXgjRI9
fmn3LOFetJF+bH1GI8bWYS6+tI79dAEhRcxHVVJL2kbwfsJTVV93guqYHIbsUh32
cQQl/VdGhNh5ycKkTZvLuPzazGJPPeb5Mcs9jwVUQJM+oQmIOUDhhBR6FugsHGa/
FnsalMXz9nITJDH6ZAWHauckdtuRL0Qf5bPCDGDbknvD/2dFtAM5CCtF7Ka4QgHF
Eyu52GHx6WcD54pu7QqnMd8vhCaaTmVxG+Bwdaqxvvqn6yW3p27WBq7jCka8Qym8
h9anuAu64rjTJT+dX+CRGSv0bwtLdtN+Bok2krEEvCpQtJqAsBb9vl0ln6WawQAi
KF6NEz6w/KEMnLWdzEWszCMi64Q7YGl2Pfr321DooqnXOxUdfH7w/tjUxDkQuMmz
H/OuJDXwAnQzwoLuOE72waTX58JKJBCUXuK5vrzJ5Q8PGeRQL4sRDqeAd8s4/g2w
K4KGXBLMktWrKUKzcu/iP+GwCa/KIrWQayJQXk4LseuWKgvxE9AyKSqz0xPATFal
51MEal5SczJMPYP0fCmtyQLwp11uB5qkkyZjiPfDX8NYgvmiP9fiWc0vSASHUr/Q
Zh21tIyQ1kDz8apmawgQtWZIk3rgGxo/xHj6Aw/2OW9fxlXIZLDtDilKjJD+mRG/
xDkvfaRa8Ngt5ZLPtn8c5si0znaBotO5urngbKmxHvHmhdKcKg6uS3MUV2WMis/v
KoygvU59hMC1imAnYdvW8+ceNyGc8bWSSlZLs+F8BDxlDQ3ShCX4fQnylkcO5vC7
7Q9BMUhJEGO93ZnbXs4Ck9TtX6GKMQ+7IqCXdqK8jyraSx4n7EornQ2nAHf/Ytu7
zNV6XKrcRWSdAJisKameR+2QI9BWaYpP9UwgveGxGMmMg1AhlXTJFDBShf5+aRTm
ML8KYoUDiTT/aRHApo2s5HCwc9ZMcvhRuv/qDNF+xq2xLtpl/4+V6bfZw7cjNdEU
4P1hSiW+b1JiRP/ZMrLsledxL0R/lk8cf7aeXVPggr/FyRYq7hz6me6f9RuQrFuw
Ip//SYyMP4osRoSXPPru7Kqoq3oZOErup5gTSGX8RaBbpbEQlfgxJBgf3AmhtnyX
am64wfz5SePbJqXERqGx29KJI+gqVv91vrMe5Tvx3OlDWkzRGvMMVe54+brPEqQk
r3iT9LLsauv2a/nyUg2rqZgMINRrNDUw4ZjQ0uvLGc+RmEZrUFEUkcN3J+tAos+N
aRKTZawr/FxxhXPXM9O7K07ahJVX6Zn/51xhsFRAmHHu4S7Aifbwk4sr7qzMergn
dAPqNjMObpXdaoN6qTaIEemRh6ne17rDIYkQQ1wJNp9TuCZU6Wtt0FTMUpaygXQZ
x1HtKTR7/LQ4h1LqqxvNjWU4oXRaoPW2vIHW8AuHcB+3F7r0Kz3xuBlzyw3sTjMg
6gaBsFwvxJJ4krnvUzIFZNc7d1gfoJvDQsg1GNLgfkfkBHiaXkvxRXk4TVjHccz/
1SkzALZb0DS7Kokfa9vzfuUTJpsqNj/Qj1xJUsM+bklhQk3LiJooNZ15kdxedq++
lEFxAneEBIV1kEYg9nUdqxy9Iqv1gkddofmosvaadQFkZblmyfWiXmzRoWtj2DAr
fjKAEvAQbA5T3NL9998tcuoQirU/lozBA+h3eD5WXxCSWp+me37yc43J6lHikIPs
7wvWSMTMZ1n45Ab+zfcn26f4kGUgYMvlx/9lAjtxknwLPS7QT6wRUQmrqbKDcYiB
CFq6+N+xyFBnIF5bnJhc4TGpJBv4zZhjfbtGVvEIKJEFW0Pp0iKlCJseFUAk7hdz
ZuU5nf4H+MveobCv9CIoFAcAZqARSN3zbh4qCuunmwEpeYG/idealNciVTcdJYIF
f0+EwLuZEQMFeUg6EErM5tzckLHrDIQ3Ut6p9OvDuPg6jhBmJNXBkSEXLLV5P3Bk
LOnDGdUImNLNGqyRe723aoXP+TuMp8hMrxOgM8cHqSaZRNTRmEXYDqt6PMuBwQGS
Dxx51bwg5eB9hzkdGr5xgMpkyQ1Ygzw38I6XtP6Mw2BUXbAafxcaNIvGya+wqRKB
tyTlvYQo5ANN9lkQVo2ehYrQcPc4soQreklJyCIAJkMOOVjZTPJY4JJzH5/dtdaQ
SCqGeX2iOXCF9/9cBKXopDwLW4M8ig35TqyDGpsJGURShCZuEYq3gAmAMvD/+GsZ
wQPTrAeA9B4phdoVjsZmGNpPgxozi17DQZT7XVvdbkURP4Nr2x4+vACbg6a9SWAb
ekkiqdWgFiN1ZR/jMuy0/FJQ9KWKYsDksGzGmwT4udCsRPfkIdjXAEeCDxhfUDCy
wYUEfj4L80gKZTC35XkZFiWgUc3ujCefjceVwKEG4IImVjweH52A/E8k1C87IdKz
+h3Ebty/ZQrPJxwl/XUoK1YXGuleAdLWn5FRFb/ijn7+k9Tjr+AFClqeE1dIq2fV
SioNQ3aLroEVR93CoejmQKBfnyG3krOs5gwzJjU+7m7SpoyLQxjeopb8u9UnVzLq
VD8WNkSDXmi5gOBrse5wNHRaJeeI7JtNhCVWrJg3ioc7UQMTpLYsxD5AIf/KiavP
mgmjHN6LZg8GuooWEgYWBdcjVvGvtDhp0vwwOLb0388HtfWcFBGtbpDqILmm5rgb
Ju5lmFYymOCZhtynXqEWf87Gf2YJSA6Pv4nqkPML1QNjjKld83K2/IwpXH3dMCyc
5TaoD15Qf0ho1yZJoivi/DGuIzHUQBdXkZbRUb4xfYLoQPjhUY4/5Sozcqss7K27
eObR99tx8lfC+BAkSr17iL0koZrK9SrpLBiAuEGih0NFhDGKjQ15dKlPwiKH4ADv
S8K459C89TQUY7yAZ7DhkECAe9cIoWFQUqI6QJ6pVWQDNxTPPnKFStb10lTHh4iG
8GsWOsfzNROjIMnivy5hFffN3dd4SdAvQ0d43Eh0iu64vlLrgJcrLhh9pz+UZEBR
TT3mgq/tv92i4kZNuUIPAeU6z68TJVpuUStq3pdXo7qbo8Bwnnv7EBO+g14QJuPY
0SAN4XTU/q/KOE652LQPC8dvH07RLRG8WefA2UHps7+6LeSGyZSVkEJ8jEhxiW/m
uTOqoPVN3LvvSY9VnTwEDEhFVSSbLkbmste5CBCjmKQLdi8eTiZA6szr++dY5Zrb
6W7GhwEKb7tuLd2Crho0QO3Ukk+HSUVkNOoKOR00GrZ9Q6JM904zdOqjhsvlr5lH
WfwZLJo098hudIimKq9N3I+49Ky+aoezq5wI7gyDPXgBOq2e6kJjIm8xdFppTYNV
fl8xQmYgbXY9FsxxNqbebOvQlx+Yih1VhbBtD2YTv3TvuWtxd2IwEoleiK+fFlg4
Mw1q2BtbT922Wtxp+ogfMrYATtsx3AHkmNhM4ns1UVPrXn2Lhd48KAgpUt0zbPou
HZgq0wGn8BEbTS5AgtCVCQTfY3iblPM6LBHB9FFUy5+LbeWFsdMFT6Pau5VBJtY7
tEpJk94rl0jDeEP5/foocVO3oH11HZsJAqHXrw40u6A9BdajeIe73IuzoXrQQZSg
XyFToEPrSpPuHPs2BvnyvmQJLcEyYu4qlQThBR9t8IaKJgAjStD2K/iXllFccGUb
vTF81buoz8nLJNSdZVVFJWnAb6U9jk550vHxBXItSrgDc5EFsiM2IBc+YpMhELeb
TEnreFvRu+w6JeeyaW/7mLhz+ocxGxwIU3OAgy0ZY9q/1KRXZNexJX5qgMh8Q7qD
0O4fhRhCiV1SlvX1xZgJrVjOceZuU+PjS8fzuID1hLdV9PLqFCyM1qxbB7f3kv0a
CujkzqZzPGSOWcIxhmDz+Sd4lT+2Eem1sUxwc2kb7SZOLD8X9pjUmlX/wZx0h2Wt
tT7LEyfXXeKBgz4GCuuot21s/ZLbORHLTv0Uw5CnT6TrX09gZNQ4b0qUXwMYSaud
Ws1WYP7QHBnFKlwdaisaSx62iwZNihZgTAxHhJ5Ii8KKIXe1OP09UToqzQ7S2yQf
3eGRSPCrltT7QV76q7PDO7YboldG68ReJBCB9LNQGQthFEMuG2veUGEfoxegyIB2
FzBM8BFkvnl3g3RGolV3IjZoBGunDKEK+H3AQZZaXBEEzUu0JbW2e2PKfrU4PbW5
+16Q6+1hqwBYv5SQ9NDLEyUppoSgRgo4nJE0mCulfR/MrqLecF9WDVHMpnSGHArJ
SEgZJvllhUhomyiprlrIOa2TQhi0tgUg/sauomdIkyKKshiVE731IylxeVW6Qs0o
Ir5CRtLYWDJvap6eQTifLuBJ1PKke3RMZ/SUqksJpWb5zhdsDyDRSo542Yyk3AeR
c6WW1cyG86L+4r830lPupZHuwrtl494midS0spJvrnbvJKIE5roYj10jUkCpF8NR
HMIbKRBWXpSFsmUPVcV9DhZ4b3pKuQE2lixwA2tn1vcuyloigWlFik0E20P5vi1H
O0Oj7ZP6mD505vSy5NOrvhH6UEWj5gBc3u5I9ouN1xtkV4BkkXQLZdgFFFQ2kL3K
wMkbVa3ZBUa/6Veg5ftyGJUscr4glht7vtMu54BZlXzQrfx46dXieQqNWqzrBVMU
jfGoJKFraffX5ZNHTFobvpl2Gy+bZMeuWeoQKQnVAqhUQ+HpYcO8T6G1BuyKCQyl
3sAknIic73XktF8EgyKvZF3nG9bVox9zxutVid/wD3hrBv5tPDsTDqXmOj6JQxyR
bjKtPs2KgdSfzObYLx2uFU755jlgeeyJqBr5H00MO1nQpcO/tH+r9vsbB4qUJopT
tkvMgPN4vAGDtBhkHblW53kwtvhBBhiBSQsLhzksNdt+1W+wwfh4kYE1iyQrkcDI
7sRM7Pcc6uRbdEJwfgApDF00xWOJnGmpnTYq/0AjGfnC9bWOCTL4ZGE78kawQVzE
AxdwYM7XSygwFvRPndnxBQrY4zFSlXVfIE191LF4whwgIG67QxzSz8TVVwKnSky4
bWeUDPicf4Pue1XCGEaUTFqWsP5THK8YMq3PWF+32qsG5jMb2bxYZm74zEvEP1FJ
8Y8oTa7oDVfB68GMnDOZ5mLWAeFLefR71IrV16W6YWu9wwGb810POs/vAt2oESyZ
zZzQkatGvNwLwGOR1SfBIj+dLBYawsIoi76lKbLc7SLq+VHiOqHhkdUM5MiLL86X
tGrRXC9bKvaebU0shHDxfw2UqkbQYLFAiyhrHDaYcloi+aCWIiKeKeMDcSArVY2y
0WLl/Ehwxp0kt3H0j0YD/xI6nGKj23zlSFjTizSrklEOENhRXWiDO9qqbr0oNXy7
iGPpaeY8uh6zLVJVK3RHuVPpHTM2Y1bqIdzZjpwrl28ihCYLmksWH8HsQwUkHBn3
VVBIBMga93SodK7X3fIh8XEgMuy4GgQu/8iI2DFx9z5ECRqY8kEvXKKuEuCzAQsl
lpPbamOOBLG5u7cdIS2EFC2ChDTEOxVipBoNfnuLo0/Xx82TDD9Nd2YoUvXyBB7z
QuVnWRweCJbyM36DrSTvKTLuouLYDjLwngwdG/JoDT9LoYp+qWyxeSXbCKeGYNEp
w5qHtWKcZtgkjX95qCHm2iY9YhxyHa0UMxoqjH9sv+1LZXaiLJa588MonPEE8bjg
wNtNWlDTk8X9Q5HvUz3xA7+anoqn8xJJbMIYSkhNipq/J/U+H8rpi3rH/19SpfUa
BFa78zbKtojk1MWdM8yqLkeVTJ940LR1qTsW4ziuDvgluW5BRK8Z0E2bLQIhE+ZU
UICaq5mRcihdQJjNA/s/D4VEoUiXWqGvZF5Rf7V9WyzsnJB/5jv3eOuEeTiGnyrv
aLp49UF+NtUv5mir9xvIO7zzNmsctr1mrn+f9hmptwgU6GcA2fZ+0ziW3g2ASMwz
imvOlBKvsD9lIJsevQqRLXpYSO7Uy7PuZxOAjO6G73xYNYf4g12n1uJWDdmunVbL
uicGbQ5LxjEb2bAnFadWSeQUaxSVYU8R6HzPR4HbrexjVIkAPmuyKrwExQVH4yXn
FAKnMSse/+b1oKCfbh7zM9jaI3f9P3VjpHN1qplAo5P3bzJzdWOCsa3SouA9mGsR
3GtbyVf0IksRkXmBtyywNoDhFEbZRU6ClON6hqfejGrBetFaynW+/XvRF3pQ6yRN
/dVhtJtKICyQZgXiwR3hmSPNL2NGe7cROvwjwPUytFXbGPH7pcz3azMyq/kN91lV
jw8GBxVVYk+pSGgDljFJqH5z586J4LyTdJUYS0bcQG6Bad+JXXXNYGkiS3eYQbWT
PFvtUza8s6ccghQss2w1gYzA7yATtTc9Odq67FYxYlqXtzv47VPa0UgP0XcgDPoc
XF8vUwgYKuGBv8IxjufMbqb1fl0Ig4shhXQ30oSqNiyE3gFYudC1NJwdYgfW13te
Jv32I2nt0PjASPaIxnPr4WrPYuBo2/JYml7xPk8nMU2S+xWndg7V9HEQEq1dt8fV
Ux7brr8ZIVqp4ztqqCSOkKiHno/eNr56JUqj3Ea1lp3ybUM01nBX6E1O1MK00T78
96MV/jXsexh8NrNbNSjImkybOTEMYAwS/hmsxeLSFM+k9Ea+KS3TGREF80E4Tg1Q
2a5rZAPVfJpmFE/oDBZaKzpwR4ch867rKW3LjQei6YJdXHJwWRnnzmtsmGAxB9Nf
G6XxCDGNd1wxOWINiuMrMvo93Ku2HLA1Pq6zZQQdpxS6jYVbY13uOKvIUA+o8HhL
aaDC2HXuBZUo38nWjYR+vl39TdsqRRt0mS5qfv/z3B915XvcwVCdFQ0nZOOVxI0X
l0tHa2J0PM8QAO0mZJu5ocg3XUoJ2uKitdQaaHISWmuWY0Ai8kiTzntlCj7K2EEg
tsBx1nxWRdc3bq6GDNqmEIolVcnLdd7BK6rcRZ9KaV7wWhMwT23mcaBp8XVNx3L3
8Ng9oxWhJ3MZyCJ1ToZP+0vGNOHe/6/SEOAJENUjShdR6TCCVLJr/TmLLJ9xls4F
+SM5Klky3PDf1Tqj8PO2LswfaspADDuhrNmKJmE/Gl3lqfaF1LW3h+OZEGrz2QkI
rTVvQC9ekvfsFW8EbktjKMUhGAOAzgqAaFSgLYycMEAoxa3LTGXB9grLrHG3i9lZ
fFRjhwARzX2uea6NOWdYzT0B8Wg5cf0aUsGsHw1MKMCTRLxAPxxuOys5NC6ratiV
TLKKMTqUvm/Q+jstWQBpERK1x3zfpKVpyS0Xlu60KSsjkynEDKW+GYkdX1xhdula
bKM9wR7e/aWkNsWDAGy8NRrCqKC0g67ycQU/cTIWFMxrzGwOHBq5LWvlIAtKLfO5
ABRlm8W7uTIRp8xJObGaSj8i6qOYmwy5J/c/Zw8otPRm0SUpMzYigK8QnJEPCGZa
r+2yZjjTQo41O2lAHganfoDuFhS5htCUpqCZjcziA7cbcj1Z/1zrjtrwoR5AowGa
hP8kn7Jyp5zDnHdvjifG5yBH2UlojEzz2HpGvc5JQ9MipG4BmjtTCRbXabeEiEHi
NNQNa2P9PJae4hNjWE6CiouApfFJJQnqSFW3uMxlvr3hEAIo9Hyyy8hMivy3pgX1
L+ti7tUT5wdY3JylAjPWkQ6MM1vnXcFXJ9x4fkJ8lZnaW4hF5zf+JMblTecHu2hW
MaGUj6SEO7PbtcqEqS3K64PIBOWV9FDYAy6tQE0Xj8mBGzRA8i8wTmHVv32HiBSH
eWThFKQFM0GtSJETcw2GBKI7CBQUTxUnIi2TGORPxrkLLX5g1UImrE1zCYVMNZyI
1n67MoXJE/S/WNMHAHb91A46mwgEU6rt3kDymPSRJmHUDvqkaQlpyjeVoPI3XZg8
KClrPsYzF14CVSpHhmujgEdrbixPw27lDtiBfE3NeiTN0tz4JBqfWB1P15kV97XI
G+H+XxHvirVS3fMSwImY7MIJ1u0r6wMJoYR7iEjVzUSazM4En8qXdcWemI9zZtkT
xP2JZzZ9u8zJ/pB2E8skMkm9xJ0SbI0aD+BVduBXNhntPUMNy3Dn3lie6gmxl9Cx
/wJzhqawVW0xWs9JoHV4saOE5Ve9YzwA1gqcMEfcBuDl5scvsi2ly3V7ElNszHvf
iIM3kHA3nWkYEvSx2d7NfQB/K8Bya8GkWSrLTjeuxG5JJTaA1+7Zp7sgi1SUfMOE
PQdvm0TWQHSYnsEysRQtpdxcCNpQjWUEiY6yrWCFXzin93ztIL0yKzhlUhgAd4Zv
5gaJP0jxNVwtMTLGvQtcfjW73lTxFY2qtWxg2eT2FTXWEU+P3fyaWjH5s/v0+yx3
36S8ClE1WGmcNCnwVHyfZ0VvC85HunPJz8RFyOwz1aOV/euQWrNUIHAzSgKb7UaI
KG3raGWN4ZYZyX6CywGGgh1XECM6PFROlWAxXgq4NVlt+iscIlQSkxR6GqfxboCy
ifcmXtsTvpuxV3ngkoAre6NlaK73MZQYZLeTif0SyOinbO5qkqXQVRU/cz8aPK2f
Rdq85Y6xXPMjE46WipITWL1oTHWk9D62F1P4OhXvJVwQJunySD1LXLTbe1kR8BHb
mm1Q3tFTFhLiDwlE7EfqTInP1TeSkHyWXDe4sgJfyrk4p1KGcXv/C81hT9WWdgLW
R9OPJIyPckkVzD8FEkpHVGtGz9KLDBy0+GFQhv20P+DHcrxmupZubhdf+eIsY3ey
DayPA5JmjVFZTLmWNaKovXwtB4/+X2rlOhgBrFcp2T/gnZZhGg4BPXGKI0kN4YMY
/CY7ZlEHILGieTLiz5Q1wksoC92ziC1JrzeEv1rhcGS15JiONXdBGDQMvvYThcRw
rS1hw0j00S3VQSgyZj9QQf5djGLswrL1Ri0Iwky5TUg8ULf38gRbMP4Ex64a9s6P
NRRQjtaWfJtTw4/TdVmQeRGQ4M8R3NjtkBj5p80wKwMNecnyXKmWyPFd25gtnxVC
YZNOPGJws5zzN8ojLsRX/dA3ymVUOGQkJLpu9W63/JK62xsdCr86qPega4MDBt1E
eWq4d/Dio8d6bfU8pykwWwHcrJIUInn7Eoazq3m33I2lulCMNr+SdELwf2zJ6wFY
GSd+Qe/bf5OCTtqSWRdknpDpZlqh91jg94Csq9nsw0U1NK66bv/kBuxzN0r1s/P3
73LppZ1u0MKe/SRZ0MszlqRi24iKPCy0hVdjXTdZgcCV8mTTo1GsC1W1qv4WDvZ2
08G4gk5zUEpz4Zm7O900HBR642MctJPJAHulwme3AsLchTA1ptPd6rg6OffKJR3p
89gv49cNKoABGX/FLUiJQffq/rBOzExkAwehoqc2X8VucwXzLCiYwXc5b0c2PdFF
WVPY0S8ULqBlNIsi4PDYgfiYgk/nX4oxs2nrRgB8ff0mFQKTBk3y7DSmUiItX/k4
NLH0eDOTg5iHt4P3FcREo8jg0zemaa+JuunYKFUpoQzdgN/ixsRIDKw7B8jmJl9R
ZasYEsSGvf1EoJRGSHkEpeF7p4GF33zAr3bgI8sQRV8djJzGyXh1UthG9hOyMNNU
q4eSgRzU0maimWo/woSNegEK0ldf89ekfLDnQUTUI9zYrvJk60CZZJhy6HV1fQkM
X18VMbEINV0ImOVPFkHK8ix1Vk20vrBvOYypANEQRuF7h60WKUdo8qzl9gH8WdK4
D8iDf44BpxyfLWmMvev6yPn1CFFt/gnnEsrsmiS2zZIPj7qXS05Qgq2NWE7KOdM5
KGZeklksrK4emsM4g2XMSHnUPWfWxI9/wtbFBCJ8jyXxZu9EPscNdWYoqRykK+0A
0xR7abOqphi537Wed11W9y/paZhwPHjTY30A3xIpEfQx8uQT2ZaYfXyUFN+spvZC
sp3fc894oS1nZY1dpNnWuCGiz3GWKpBX62BhaiuVK+U7pneNQWR0YWl/gt4d1YFa
+EUJv7QcSAdAZJ5LSLiH2//r6MfCCU3K3iOcEeTTSfKF7ohDBzN98/4oRpgPcc2j
j/tcsYUocW1URzj0vK4LFVQSF9kNF7xBeV8kJG1tkOS4NnuIrnx2FBb3D093NlNi
J76lm3xYA+BKXU5w3JJSQTWsbfiO8s4LYQjXLDm4fWpqG2jkouwydFPix3zZO3b8
tJHU5TY1aX9LJ8xI5qP8nAAIo8TcqFRqN9BXRWToiZIBJeEkkuTE7Vt+twd8U1Em
MQLDrzIiUDwYFW8lSI62KUfrdEXT04dqpm+2efG9Dw2j8/HnNXJvAo4gMhwNF1Rq
G/OyYcdmFoiK1hJjoIkyBnxciZCCuu73ULOlQc1Fbz5hN9vivsbNwBKRLn3KDmSw
2TnCNYZw/Jf8n58yYV8l2w+LIzU7WssC4cPSk84iCrXwzvnWOCjum6KqSNosehkb
Xi13fz5fgZWXcZeokcxA9GFuN46rE61wfBXo7W7ZV/SOXmIjF2BQ2FCd+okjmnGp
JK/Mmr9N/W0pqh0V1UFeTKYIBw+LIxcB2SrpnhjmTIhqynTiW1TfAVSIKL323fC6
ehvGmJfNTtaNYRnUWM0mmgj2MdjYKdzPh5uAqPrblYbVLwIkKdqzcJm0kJOzsN8+
JmgHgaU0xk8ZVUAFaz5m45xcEJC7n4dgGME5G1JgV8STrP4Tsu2Yi3GpnVTBA0Ce
7ODcVPtaStPLo/W8faj3TMNTFI7a/r/6WBNIZa2bq9QgFir4akFiRMB3QM/dWEgH
8prZir6uCFgul85fmtaKj+cu/AbNzrj/3ZHbxfLEBTR3gPtebAXJGS7/bNzS0B6i
4TBogK2YJAskDEHYgUAOa2FD9sqbjmDj0mCpgRs6qgiFeGhNWX39XZAwc69iPWep
PyAM2lb7OyPAAyLL6wV21u/P39WwLX4bbtAWjv57UiOiSeHvcgSkO5wLjRl2/Cee
ng6ju78+ciDhvlOghu0FhGFRoSAPG+weO++0FUcH+TMhXZ2fR0hNsCaYe5mk1Eip
heYgpRsgH3O/ihiWe86+KYkSfojDRJhp78GN6cwjZy6CbMBSPPPRhhCUIGW2U8CS
2rrlXeBxn8ian005m8NpiVbOeg84TR4mwqAb71ho02lrw4lS1qspnDolUxTNNIZK
iLSj4nBFHQHPlIdGhyQpaOcKyhV0gin1UJQeR6CheNHDAarwrGkvDXILV9/F4M3i
pt9PuBJaoqADFFzz+gbbYR5J73rwco42ClaXOXbELxgAY7ltO4GgatBUOpcFLsnH
mFMLr5sSsm/ampyzfpYF4uT3vzXDjV+YWWI4X5PnsupI99V6U8pk39lK9WxHeWFN
WQ0FK34liDEBJaERlwps4feQjytcoS0AnKLo1LvLaBQaX5a/fAhNrC3M9Ece3d1G
bzawmOAcfCA/ZnzjR59eLimtK2+g8+GfuJHvuqBgTXOZohfnp/niSSFsEkPKxV2x
gaWW6/w0kSuHNIbmUlfZ6yOt4gb8roYzZJo35Bhc3qVbSA6JzaIuLr377HXUJUGT
7QkDSiLMQMJtFvi7viOybqbKoT/L9UkuMkM8+qJCgQTX5saZ/mP0O2uVoxn1c6kL
1qxpTCh67nBLS8gYo49Qf/TtTHyzndKAXX9fTL5JjvIMxVtsQ+68E6RJGU3G0lIF
o6dvBMq2+ZIrznqB/w2pScHMhnU45SD16P3GoYAV2Dh2rPJnz2MOl8VSfloanq3v
Mm188WHUTz8q6eUlY9YIrx0P1PjqWQi47n3rJz+u2zTmYicvs3DeOvDyDBIQ6ELB
HgCKxL0yzWEeZCBlRiOSyAD8WqXBcWHQYVji4QBET9YnAjRCx5shcpG2vJ7aujY9
juYQy2CZ6qt4wn2jBeWJBqs0zjX7zEBBj8t11FdSpBV98PVlMtdDXv9ln6An5alk
id/ZObabgVnGdjRorVRu00q32ebJ2blFKFgGTZAzskji+4ryyje0jTO4m4n2oA5u
+99OYZBFLq1IlwplDObdp8xzNm8J0O9Cz1C8QLZMzmnVuFYUmWkK0JKzVwfhMB3M
+Fz4ZYlau2umRyH6g1F4MaygghbaL08EkfZddaO7pXQSjXY/982KtglnEbxO/PhU
VqhV+4m0DlvcRQmxCduOLEYuY2ZyQE9pdcu0FL2aEAtyOuMBn80747U1dOvPGjBA
kR5ACGWj9L8Llejj04GC+YQqJQ5MWr9FNwrEVsS3u15cenOi9ZDPeCa1jNg4Vcs/
XwZiZSEaNcuw4IflVJSpaHRNp8t0K+U8HfVrSLndoTUAFwZi5d2clR4/YjxqZZR6
7k8/6h0VOWvPLtcD/yE50eBEr6FRSAtXlhtl5KwjGD1W6l1ZURqWOfmqlVrTsyO7
JiwAxjMt/aoTUamZf1cKz4znnzp1Ow44x1FyEcyttnRIJdTjO7lXI9hjL8AC2t3u
Z/Pf0phMxQ4zg7h9Dpd+eKMtraiQ0FaAEUK7NsUUCsdbPzSNVXQUZEt0Sm+/hm0x
Cd2uc4kp/Jd+CvFSagoG8iBDPre/q21KTCzXEPaXgNruiOa1yzajyC8Niw/J8tpY
L3WATko5TdEpnqOzDMH6IO4PjD1IlZU+kBoALHjEhzC7/jzeXA9xeVCTu5sc2Gk7
7jee1Z2m9qK6xAoZ3maxOYwsD+4gbv9bF6Q/h2yuFXvRe/uU+nsy9aUtR82Su59F
ksGC8kz6ea50C3A/SsX6mTkcz8poNxouburIKH2LEO5FLzN/kP0a9pc9mSsoIj0s
iNYf5KLCkhEYcADNJ9/9xGhSCJVn07rbJhanyH1HhT6SBLnBqEeVMRGntnWUZOZ7
6cK66QYMl3jxTKRANUWG1kE6EkdScG+ojtDD9nev0xZesKXJJ5vH7IdfRGWz2Rps
tYXSm7c7ZREAVI0lMTb0dZN7LXBrc24eH9g5w2L2FpedaQaFEp3575biNjVEA3rQ
6zzB9bY2YHKpbuIFJf5LMNLCYpUSSHfa4hkmcQMkmOOu/PgPtiSMbLda7+hw/jAV
b5D1wqY6gGeOorQ9YUkF3JnxDAQT8Eg+j+GllYufysDzHBOb1yAPuxe1FSMnJZqE
tiAe0++othWuIicjzKFL7GYWVd4z1GCmOS6nlGb7zIhB7oup+maAf9F71aSNTJT+
w36c2tsmi8KrTknRUmPm9elhidZCoS4Je/vvRDVISdpmxYZa2T8SzmAqUadrJo1U
uz1do0+vVonxy8uFuj2W6XwdX+gla2VW8R9Gsz6Z3gaiAQPE/Oep/MMV8YHeGYGu
JOk6jCJF39Oh/PpJr4YAc4g9ZK0FYAFnA3wxtPtMcJllisDaXMqFmMJlKGW88/wI
oMzUSRJ5DqOQ5M5ODZ2xIt9v51cAXczjxyS6gUuO4d9BYAH+bPIUYle+6cTiUE90
s5Ouc3r+hdcRPrGGBWSOoOFYGP1/i3lKWXmpfragVZyA+GUBHJTlhkNwCeRGNXlo
JxsI/1q8X8Of3BTo0DMN6zf0l6TQ2YrVUTipWflFgj+O4k94FhJVDG68RiBzcxSH
gKtEGjgUq8QmaPlcX/AFXguiNtljVR5nEBGVrO3vNRzOMpxQuXN0bq/Bz6GxH694
cpuWj2eBCAuR+KxL7dC/n29tAdm/l7em/5/0gFqp1A8+1Rg7uHjFQ5cT/rQA1bJ3
lkN1NKzc0AflZfbmnGjllaliPhOk0y2R4z28Ickf1BwTnKyVW5CGLwOn0owKcYNI
h5Z1zaLLq6EvyzJoQNobe8Sh4QBZiz6Lxb2+zgrWVp4dYeiymHk3KvNV1MRAn616
RWOFfINEtVULA8nKXhA/HyGOmRdh3aRgqcjNmDqDLJnAupJGeJvbRQDo+U2OD58m
8PfDAr3H7je7tOslOKY8F5EVWTkZ/Owo2pIvmd7DPjGcNbBq4A6YdJuRcG8jldjJ
o0sfOs564/tgTfHluxq18ECfyxAOdsUK3ox7FpLhq2JjmncLrkPAQxj55nf+i/+3
SjgjL/hWpdSNG4LBysv3u6GD27J4a6cyZ0SDCpMAc/jmd012iKRWIAD+jznkqP6j
MSaddni+iNaLqMXHi/CcKPOMa1Cwj1XzYiLsH25ClWXb9hp9CgGMLGh8Rh1xNNah
GY0v9MXX1gwPjvkwD78dTsh/4Ot+MdAqGuad6XxN/kazRnzDkkvMh22JlccPQ2Ow
EEK9PeQKjLra7GW2rA9LMPmnBSmqNTTSMv1ebMm5rpIUCyX/1gPw+JbAHeEQHkoa
jO/ZyF3/6MfmFJWwxQidkfFJUteq0pzdysi05gIgthr+1mlafTKUn0GkPG7aNn9G
3DxX7jQDriVNFaNukDzZKL67684mMj4xHTV/pBykIwWxjl+17LRPrWh5aRUkKq/O
dmmeu/Rq5cpoL4v2yussgj7ECxdiMnBMUzR3ibFoHHbmvWjFFrbsoOIu/aEa8vmp
Y6o6jAPyY22CR74UynBQmbkcyPyg9H24Cm+yPFp9JV/h2Fr9qKt6YIKqlZRJGlhc
ySNzPbt0DszV5OSpZY+xzHcP0Xt5Tm7NJwEsDz4mkcjaeuE0PvEw/neisSMLhol3
8VsnJqdWix0pwRglodIxBu1uWwU199bIL9cspKX0uJ/J627t5CzYrehPAoJ3Hi3I
WALwqMq9JGYUoUM3kHPpmTozcTQHKSG1Y/K0pbFKE/DAuC1/psHE+4M1ILsoTLNY
5RFllc/nSDC7bljW0pNX1IF26jzNXSCE78rzecpWsyNt9CIAxWia0t4MlxsE6Cnl
VIlQf+6FjwBxbIEr4o5sP3D59+lFYSSbiA2RuDgQKrgpjSRWo7UsSOXmWN2Q6QvY
fmtkr8UKtCfuqdPFyxCPfNGqlNUTON/A9j36vBDy2RuCrhqcUYAkddnsClNsy/tq
O8etM8DhSDSHzc3lAeCr7GSA1DoTif4oVCPNVy1jJoBgu4M25iRjI0/MDQ24r6F1
mhNoFCzOrEXq6eaU1hq7DL9wmGz2hoSSIIgWIVGxk+AjKRRwysD+L8kgAsBwJZ6V
gWqNUrTcbfFT3+zJvzEGEOwIrM4gjk5FlWRKw9Wx5Yt2JjRd6ycWOFJSFFO9YZyE
BNx9KGhtezMwpnAhIJruYL1El4bEFxybz0ioub4kTec86FsHS2egn76nkCYOrMj9
0qZ3tMWeZPvbx5IdUiec8qD//C8hwbIOqXD4ZCtmnT7H9NURs8QWcLvJRCsqxgGg
DHCSVbGZARcsXXH0r0lGhDXqNHCdj1gq5apdE9UFvGscqslyWQCiCRjqpkpr93MC
9IgUBxqvKeZTToXvySL1v4A+mr/gDREQG+x2YQIr6WBfmJDQU6+6sk0XlMV/+9Eb
DVwlq2pvHDtuKlp62pZ/Z3IjzQtYsHek2cuI4S1oCDj92cIUxd/i+zvV4U+ep9iL
m+pxX84IB9Y9ozI+TIX8TtR1lD+u3vwHkZObXV3rYTxzKSMGx90CUkx5dnyeuHMz
sOlold/ARxTIVkLDTV0XwX7TWfxYpV4xsqT6wRWLRImGMGIxlhs53LFyG2YKLiew
KU3t0jDKkPG3ghlWsH44q53Dq0HcXAyuJTr2691TYu+tG5Dh3Kp84vhscDWA8bXo
FAyv4Oss42g0eGU6r6G6z62nk1IYWIEIITziXGjQCLT5OD1vr/ecA/BTENXd/EcW
HqL6+t7aZGUqULvY3a35rBImcW+gcRnjXnrFFz6KCKXw8n8KVNWX2YABD6lhGnQ9
9+RDCPPZjbUDxTl2xZwUYxvHGggydbwlDsqFIPUUJeAV0Qx/2LkVHPAWz/aMLf+T
Re9o+J0aldIqtR0uB3NKDJXsRPmyNTYvxFtgjIK4rLF4ZD1tYiJ8m6SfdDLxRmiR
VZFBFbW+ivhmXy3zArx+Bvsz+bMSbrsoPBqzM98GTXr1qg6ogOSRThKntn1igsJW
GwrEYJm/1xConefTbil7089Ho2MsMYvjW1fs85nffPLhCEhuK+iF0LTGuHUOzJy9
GDcRbVkwq3yHJ7ZwN1OYU3IGuhMEOkNm2D4x/K7N6GR3HlM8lOkQ441cEva9E0Fh
G9f54qyKqOrTfFQMfvBRs3NXpdT75eRWI2x3T7VppHWRU5PRMi/KpjNWuRNRdrMD
LseYo/nS/nqijNqubcfc6zPmEd7usQb34mnohop6kEpRbWH8il/ZdRZTkIgrujaF
srblGMEK38wIuCGMNwbdDdQ+q2YNpfSXT1r0ZBWBVmmLmiHYr0v69xmhBqoWjTqQ
zUo95GyDyaKXtwTyJ3TM2Qwp/35k/RVSGoiYCReSWha4ypBKr5c3cK2BsoGpYZU3
NurxHvyUlGeRj/JEusDFAGhff+6Uu6lwyGAOaBIuKM7yvy9cgMOvklYtmHKz0B0J
lv4g3mi0TLhDWR1xHOA7LyRPu0CujF9cKr8ocVMNXyORkWXO86mzrDLKq+651f4r
Xqzl3JvHcT5iOQxobJWvyqGFVeUL3+WXDAFDFRwAK/cGH/LYFjAoupUAJW5nPJtu
cPEslC50dyI6QHwu57blsEHvfHrFJTTns5mm3Hc5NxS0PWccgU7E2e5GGpDSvOSP
z/XXiXg8L5KHYrCiEg/+gKMX6Ahgpon67zdu4odh1MpO7JYd+nTT4UjHqIuGGKqK
JB4KOACYp/eXfYsQEylu7hT+QuKO98UDk5iu1kNe1CLMLq6kYnoDHS3uVlitXBWa
uOyaCi074plXmuKjULZuZusqlBJT3/hGG2F8C4nZq0UIyc4ypSP2b1diTCL9P3qF
PZEMI2zwAG3Y7wAHq9GuUlT1vFeOADF1arL/77uvbrz2MvOBCZUk7Vkl0Ao+pzn4
Yf9GXY9ciy3ohiasJmM0fnixKwNsnIXRqnrcORbRiOTKXOKWk7sQ1SXlZ0LZtRf2
L0Wrx/YIM/sdSz8fgnZcY1coq9zLTyutjzxCLIYp7mb3HP4n5lnY/gELxeyTHOvB
erfygZ+QVHy+SfSZdWSfI6Q3HWw9hU1m6tZIoy6JIG5Sa5xzYYAfL6KYXmttzEdd
Sq/GtdfR3qMK3Uhk2xI/zUls/srt7q6cv7DXBhLSKCNjyGPq3slsv8VqS6Nf1hus
Gfl6/CXUYV0zZOSyPBMD6ZX0JTCbsY3G4HCw8G3NMHxVIqzORcQS8dfALxeYw3uc
wVkhbJPlvEqEm1KDyyjHO6HFn2lk+dD8+bqG3OtHZMV3WVbZj71GBKqh2hqctH8n
7A6MV7gnchZ06qKevwRi8yArtUmVu3mM9n5UT4Emb2qUUmz+6ina3aLGjLnvhhx5
6D2i54HiNFcRY2tKdu09NOYKfn7BKZjnydwBUa8ySjb9OSMShx7RAEybjA6cUstl
R6O1BL/F1aSJ+gqfF0X/z4LMZjOhZyFhcfZg925HCcv2/WzmmJ9NsNw/33pWERl6
0Rrq4+cn2HdPAx6lpV6gUWr23ay1FtzUKxkHPOnEJLX0zHqMKP4k5bwDWju9898b
Y7UxFvwCcZ0lgggP2uusDVdU0dkqzipVGT4tZLsBt+2U16knJu4JXOPN+MBkNm+y
379yQG187Y1qIZV5cNOCHoHIp40dz6iBAwHX5zKtOYxYkRcPyh0rErMT7WyaQdWr
XHbEdAY4eFY+7suGtoCVKfuXwX4/CDJgC3GrPtXEr6H3fvkfhnzw6ZHhhQtuS8HU
H6o+b9ywQWZPIC5xCaDzBwxuX/jZXQezXOifeyrvFolz+gSl7Briuj5X2B6Q5KD9
3gDhjDrKicE8A1+OnWZS2sgl6IOSdNAe6NFLpos64FvxBbneX0H8PBeNjTJ0RhBu
XJ3WS+6NJXa/gO+Icy4yBUbDw+Glfj1W3mdjytQsUPb/oj+LW9L+HlLTTrkMHRJ6
w7U4mwiVgMpEyxiXgsWcJ+j9lKQ/hem/NOWcyHjmSpnGnCb5ex8DjyBXDI+rX/Au
CuybVz6pmd4te4egjvVYrOl2hBfKJWDH/SdRnB1nLmwwHc/XLgUjfGJ0H0osO9R+
MNVsAoOLMJENilyzpkGaMoD4jnZfvKEMO7OdKywhX5RQ8SvjGIQuXrNlR6gvfny1
eyOYFgkwLdHQFmZm2CKzwXbEM3CwWr8QNxj5jaHEps2zbClz/B6fuLqbtXtUgshc
kX+DtDPuZVCqwiZtRvJ4U5l8ZiUb16jaZGyjft19jvfSPdWtSmCSug1DO1IcP8ja
UtGHaYKpkI/cGMHYmS48nJ0iRJbBwncs+NXP8w3/P9awpEm/ZAkUB9wgoUn0ryJ5
3OPmMDDa0c744olG38iVYYJXNXBr1L1d/sNweBD3u4iC/466VUzTp/4e/B9VtLUt
zWDQ9c6VHrr+O/9rUo8CdcODvejbRfvhxCVPFH/X6ESLU4p6ThbQ09cnGeBaBCrv
AZB42l2MyDkq+OAtLM6w1rkae+AgdkbvvSwWUCJoXHRK/ZH/dNxe2pMS3NHjdxfw
HeE2KuUMUfg4FRMwNCwiKitPn7QsstJPVdfSDwNQtiMj+Ek+DCoKx5YOCZhBM/WP
+fHo6dvc/tkcT9Xzn2CuIMSpzNQILXUGIR+9MpfhcJq5wp5k9+nnrEcE0twrOvk+
GDW5Rz0JQZBdjSOY1ICxE5syTIHVE1WbiqLQ9HG8RcNVG/HMdgRDTBHPW9bd0msr
oQrldDGn5T9YFgbjrYJzarbYrCWlHz8VEiQR8NQ1b+I1Wsg35iRfr97/DCASv+7+
A5p3LZ67bTDjhUnlWLeOQ37TSZyznnP+r5O2xV7Q3lEY3L04PbEzb1KVOlG4nzmk
jfbuFqZdiQAKaeBgHYLfp4ezEE7WJvJCiXbxWZ7HQIgD2HzgssxR9ienriiZVaWf
3p9iURWL6zOr4QjiKh4rphY+4BblDYQ3LkWJVh3z57xdmXRDadHUXyh9rmVRwxdY
jApA0E5N6N03d7706pXF8Cm0gA3ipmeEDwTJtfWONXLlfBw9If/iVhfvyexju+SR
8FNIgR6woU+K4Ot1AHBGmJZ7x0EzMftR7jR3K445rbz6zPt8troH/aR/Xh1dSLOR
83SHcYks6o39WphZ7yFVlwU8mN6hg01W1e5oqdoJlsraw5Y0iJgJuuPFehQfwiyN
mAL8JBQ+k2exfTan9soZZDKwKTHKE7GgpdohdUX5r3GO+3ccZwpN47Zn5NBUXqVp
QGNxq61LSqOLJDaLVYwQfeDeidDhLW0sTNhGNR5R0ocIfiVoWm8xZyc2S/QwVARS
y4U2gkEWEDS0j7mreCo77iwC7y9YgwkzqejjEhXSuGWPDExIaOX/WR7UKGP38qtf
/kIIaOkfUbjL5YZy4cQYCVLv6iJYbTjytjxadvUsuWesmUuCFLbN7jWoWA++KpTK
RqMeUnL+oabW6zrsb/2AwTgouCPEKa7Rr9xLIjSj0hs3tRmJVuXpEuCVxlOJgG2w
iMMjpC4WRThZ6dt3wGtjW2z3s1FTGfU094KWYT9tk2gTcpl56BKANyuJsJUCSLv2
CabenhwtA0LL/79+6l2lG2J82QOHn36Uaao/y5gi0/DngJ81o1FSxUv8vAQgyrg6
m2OfLWnvM+059MyGS0wzbT/zRH9YNqmEusKYeiN6XhjnvB5tpBzp9LF0n2BzuEVh
WMmPbI+v2PM4/j0w5ApzsEKXPiZw44l2fMplZSjR5JKrBw2cd6LWE3AMPaLMQ3Nz
RcidbEUekwYDrHWn0sFh0u5Wi/vZ1pBjko2fQPljISoXgIxYjQiUw4My9OcM5gvg
wV4VRBm/5r0W54zpQPNHQYerD9I4zbakYEW4uCoO+W1QH7m/0pj8C7ZbrXok9jg5
htSDXYMQpYqKpGFqDE1FlKFkE9sirnHElb5Wj6VFeosFQx+qFx24vI2vqRl5cQCL
U+WEtjrsTVpdhwOMwnPe/ETnMVNRLj2fCuMOU4dnrCE6O0dY2desoGFZ4s6lVYgJ
NFgvIZuVj6D5KjkUARQn9Jh3JVmH/FqNO1FjT/ZtSeoyhAp11R068V5PDI43HLpk
YBUl4RZ07lgiCLNt0/nnAMhDtjJMgNXeaITx7umqX3/AKk2YX+XeLyxSkLUy4zdN
coyBDwzpbcutUyZ8icxAOrMGx6bYn/J6jiu15oBBcI58UzSg3s+pUmGR5AiR9kjK
w69t6sNwRFbBL5OCk1FvYvWeUVoGd3x/cilf/tMeCg31SWe+A5nudr0W6xaNVdTU
Qyw8n3ajig+jnEnyU+2AKouDtMqrUMgyLMKOOECYLH/SplUz8FUWi6ww9+CJ94j+
ch4XSA86uhhuIpBk81dmGTHND6ZdbMxjUBn4mLv2cATBCoMSlkv9dbzVFYs2Ap7Y
drzw4v53Y8hnI9zcReWh/hyg66JRKjY00QndLfOd+nL5oWzKXqsaw0BvT/UmEP+p
YuT043pRECvY3Zolwg8xE907vmvKO63h+1kY9iFY9NmE1p2A9sE3tWz7vr9z+w/H
WogQuJ5YkSA0dd4IVVFv/PhzZaaJC8xO6C42LBnwm+415rhaZpl8+0cUQQJP6/Tt
gIrqrMtf5lgnddyFmF/T+y4MMpPjQIKh31vjpB5gpzCMYOoGC1LUpz12VYnaE9hK
oJ10YzI6GhQi/YwPivEqoaut2wIbAXiBUwvIdUgCft3rEpNRUp3oqk0+0Za/9DUA
ystHr072l4BRixfAwIB6Aw08z8pqqQ5+ghlgCW7ro0JskGaL1AbupK9uZBXIjPRQ
yJ1ibVT74eBl0IJwzpLp2U4BIolUit+rSMLfB2GqbBhjW9hoZaM2htPXh/ZkZY9G
pTpzGHlpyXFHOJtaykIcutA1QmXT8X2mxCdqWSdg5tGYO0vG+dEp0JOBYAkQeIfE
zdpA55GxUgpnuc0V6LXduPgu6bJtXygjZdta9Ch2jkp7rAIha8w28pL5hfmB9nx4
ROgvgVrJE2QK/H2Ia3gK0n1u87jSErk/vd5+cdDkP09J2khwvCwPlFsWdWQNjGND
0bclhzm1IXMbbonAJ9B7OzKwMxIA4DOMlFAyRhnRv1Zuwrju2EhgEQ7Rco6syv0J
Z0d66bgbPD7JDnvO9QDopUcGUn9v1rilBLzaOXdxAapxImy4fEC+SfEnorK/r1/R
9z2U6FnxEzo00ZGQWTxiPSRuEUCvkiwm6nYpm1BQPPCGZy0HMCEn0oMVh35xS8Xy
So4BdrDwEZtFQZ8ar14MI6uwApOKjJrawDLtoOSL4h6pyW+VL8gqGSp1PJHGoEpV
29vwRg4mfCzrV/GYIQQexqeOBp6u7XlIEI/0bG0rvgyrbW470pWUP4p7XkOwYbMZ
+1nCoJj95roCt8D/D197qoFSy5pUDByGpSdfMoveapR3r/vYiD/W8cZKnVZ3XSA2
kxpA9vzn2rIV04ASFmflL8VU8FMliBrLE1GaGEUNvJEMscBztti9MedHYkEWOXjj
opYazkrpjACgNWWz6L3snlpp4JxWTn8yKFIK4LaFjYKX4gUTeE+RMTCt9km+u6la
uRZQpBN55ZlqyBBsgZvmosOj/o4ylOUYza1VpMfZ2fYCcmSxKTWd54C73ArXuxgS
8D/JpBsc8tUN0jwKeV6QFGF3SXQlGG3tok+/kjBawtI8bmUUjlQ9EUFK36TU43+I
2T3v8NGI5nR0ja0CiJL+2xvvLC0/c4J0OshlOjBieB25/3gNjKDZizipGq4mIKxu
NqtIzvFXMd7EOFVz3zYLqR91FO46l1I2b+bnQdg3OJtoVSs39MIEwt0LCR7zLB1u
UEZ54Ff5faxB/rxk9JlDJmIY5iXJGaWiVTDCBh7UHwSdcWoNK6UAH2dHu9SyFggy
roU9BLkDd/Tpi32bQPbVlGv955ZJBBKJ/NhgYH/hqWJ3wITDZHalZufmBTkEM4jP
YRa2IPScK8Onhzs3davLF0BgX49SdTyxM2sVo3Mi2SwRd/3O/14R7itGup/S29/3
OY8ZJnZLfv+sFAiTUpVTo+uZdCOYhi7aDN7TlTKkNS6dV+99ntLnFLHYHVyfwCBs
aiNylQ3PsGYVMFeN2slwp2zhhvjZ3KMmHO8N4FXJF/5mkocFDnxx6CNUW7b+e4ZI
xJV6mV8RbCyZ+s9r5DID5E7VEAiGENTmYXXcQYEMsMklebZwu2mtx0CkPEBtgl/2
+2deeaY+p+uHf14PL8Wadb9moiSybqUR7/Au94IXtcrf7PwTsX6kGmGJGoGPtmq7
sl19JR/mWe/5I3Fu0zK7T1Ng7fZOabhN1nN5OO+fsCh3ZXF/6wCDuxfrdHRREokW
InlNVOyYRaE/FrMDxVJw/+7lB59Qsrh3pnkmk4/OngejnkkD6TwfflNy8D6aagIr
gh81rjMYGukFRDIomtGG9o+W/GLitsObLBopu3yGYTlFMNDgNE1WErgEJk+nqzai
YoSeNBv1dlhFsH9wJLcIQNp4lOTjlLM4hjJ0IckWiaCyT7Q4amHQJ/MnRybSIli/
bPQ4TRMnjyz1VtHUQ7jNSlubDXdcGy8FJvYPiQF7PvbCm6jw667QnsdJuDiV3Aao
A9zxu0LtFe8PyQ/TkxeEinMTWuLC17kKgOAC8wo+31No475O9q65ujD2z1xTIoLn
i8GcqxHB1mnJd71i/oXmGAEqVfhYQOXPt2iX04GMm87US4korTCmHqWIisTKtiBC
traHeQo57eye/bGb4kQ6vv98XbS8ykqWCvdfVYAFcSN0l7AjuiZa/i1FKwT8N559
Hu4Sx4qYP9YcsWGoEb2K1gyT9OnpduyXctcUl7otyQ4KQBDLjlPgEz+xoDZpS7kZ
LFTg7p6usbt2fM8R9Auiqpbb/5MTYfY3yNFGGjPMGp2KXdlTF5nNWuOl0mSBCpJF
L0qcjATGwfR9sBgt69g9y6H8MVznC56++QkGZug/CMbBbApGw9wKlGPCitGcODbu
Cy7N96Bi1JZW2/GC57KhBuVEn1HvkgvIRJri4WvSLchscYMM6/w0rWnA9p9LfJ7w
ixJCAOTTeMto0tTXjA0rmupVcouW3+pwOp7XZ8MFV7MKG/aZwhK6QYaAsX2kSc8H
Leu/FtKQWUJM2El4c1BvL8flLpR3GpOg5VCxZ8MwKrV0AaNjiNZ0MGaXjvzAavKz
y/bNL1R3s9e9TeIrYNaxNHu8o5x//p80t+W5lgVYmklxHCd/ZqNoIxh/Dt6U0s5o
+9IMcj3e/D0VS5BzO3khY+J/lNPtGUW6krXv7drp/gZRB5txSfH+CTePkOiaNb45
XjsuSSuwY37SaDy8vG14s61bjxD6Z/+xJhmsf8S4KF9KxVC5zx+hT91hw6q4Gkv5
JUc1CVKyd6pzoBSfuWavkRE3r8znPS8UZxUmIr8m9VI4lpRFl/2cC+hqnTCc3k7g
t/yBwt0ShYlDvDAMVtlxOUG+vjbmM/NMsjebB5pAMPT3MTtMJzUmc6aRKmTmKx/Z
Smg3P1MrWrbCMKklm+u2uw+nmaTfvbG+aqqtJGkEYlz5nwb15wHF7TqIppMkFBJI
yaIypU6HykyETQZ8gSb26qi2LMeu5qDidf4r1LLHTW3+sYk70tNWMZn85lf6QDuL
QE9fLGd8vmaH9QAZX55KLUQmKuliP1nfm6DzQBBMxUZ3AFhksgcxQRdBbv4gPUD1
grySXn2tQkzC2W7Znk3OEVXH+IKmH/u6T0MZ6hp5jFbhBz3jJ7Fb3rKMLg+Qw8wk
OsXopcBgaY7Uj5IsFtIjIlfkU/8YzZpPtWmUZyB5IlvVtvTtbs2f+cUFnzjTasZi
KNDq4vUpIPYK0EzXKQXq3KLmeWIMmDp619kpPozq/e4VdJ/jnpl0zwtxo/cjr2kJ
NGZk2KRKMsfdMOp+NFCFp3C5p3ukeq8MJtr52xKfw7b0pvqS+gon4F22bJdWjox8
K2yamZT0GeKIRwIRwzBu7yxEqcoeOaZt0QFp364wG36B3+T4IdDeQESXVau/hl54
LlbGgfn6JXMChwrDL6yvIyIqvwzvJLayAD/laCwcU4/mfMKjE5PICFL4nctVq26J
d99LzoaB/fhy/t1riftghNnG/UYIGXbKx4R8qE0H3PUqTcuIqhTMqsyD7nW8DsZh
rH7cwFZPlx/mBKsjKl4YnGvMMeOOH7PKx92zwi75Su5oTewkG3Foekxe0Aey8IBH
u6wSpGqSw1Phk1Xr4dF2fOq4Ys37LmAe8S9ZGPCh6AZBfiZXMUb08c8ic0tbBrnr
MJh9c9bIhHPFv42H71q9ehP85qwGoDX55YFo9zC1Uv+y5ubm5e05yKrXDYQZn9bO
pjQnEfSzNTmDuN5CJQSAk2zPTowj2xAAWp16VYWEwL7U8UqDY3n3ETIozRGylolA
y2TDpQ1vkKfAseHmQBoVTEfOfHokKMGpuzUDCb1lnmEjHgIQU9/eF9kg+8GlvZbY
QhohqJfSwLisvzR9oqMXm0EvFGMTTvwqatGd8kKDDiy2otLiUaFBvRJpjyP0Vap8
+cBy4VgwlvapKUvkK8xTCN+k4+vsbd2N/O07TOF00Lnup6XzCpyUrTKRmFK96Zye
MH24RDQeHJgYyW2YTL6ry/w/6IROztE7khwKpIiuuwhpNMIQyovR5r4GCebXuUHa
Kj/CZ28RmWhWbIp+YhU+iObrVyZvGeajKiEb+8J+ZIbo1TML2ipbvPNrmmRwWG6D
V2/pohywmSb5oUv1cY/fLdyGGjKIeH4z7CeLWPb2OTxUVfUGI5TF6yl5IGORRH6z
gKUTPD/GODL6PEdffa/c/gBM5Cv5QIAzE9KSnSTm/FvW26TtAWWGGSaeMf5cS1Kp
RE2+nd2dYvk3WcGl6PoeADKFVXgbbNRyE5yqr1jFegTnfauz1pRnXJFBXv7LANIg
KpPYASUC6of5reRQfqwfbJ8dlYxoa/yHQG6LS4TPUOOipkScPPhpHwi5WBfdAmZ8
13mhKH2cAdy8smke5iT5wH/Ycl1OXxX+l8nNybcLPHKELhtHgRz62acqTPORdU2S
MloZqKop4ZzV8/koZuAKBQWAxShh5WIlkB4ILSH0U/Q=
`protect END_PROTECTED
