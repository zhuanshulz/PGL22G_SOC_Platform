`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8LJxn87FAzkqfmPkKyi2HQbNgjY8VKlHVOLb6kt0xjpD9OFHLFXMzuFbviCuCH4s
2UuRnXBWDWFxKSkiDeKOq0x/fuq0TLuZjeZZRaU1cHYfSGq8KOkY3CxiSMgR/9Gj
tVEgwTU3qcbbJT+1uGbNaPa51CWD1oclP3iMPsy7eAsgj8O73mlkFQt0uSj1+aqq
EslpvXAJSfUY3S6xwYnbspjAwA5vYezaOSrV+7qtKzKaPMU5EVcqpjRBtHaKLahL
4NYrwdPVVfte+dXy99xKGuqGlv3KbX617irpHPS8MOu++9wi5EqP7YjlquWT6uVg
eI656aYu2NSjzsEqJswQFA==
`protect END_PROTECTED
