`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sJd//Y8fTUxn6okJvD93MoSoqrsNgsdN4Qm5Spl2Q1ZDamPvz1PJsUCSjLqWCU23
BouQEETUgKN/SsQHlhiAWHG9lJIqDLaoIZwE5xqoBw6/KLUoc1ISsH5EEh2TsG1A
FQh7Wd3xfd6arsXGCcgOFFdxUp5HxVrg1R00fr/Htw9fEbKqYeUBcEnJzCv+eGCp
Gf1lS4oXeuSdz9lHaQCrjJHh9zgpoMQ5liBOztVJsic0j/VJiK59JCuc0tP0jOgf
dGYKBQGvRafplojiKwAE1ngRo1uA7Oj/SrMxYTm2VgvDGDaFG+MsnSEploMbt+kE
MmZnAVe7SSrSUvREb1FEj2gJ1bGOfUKLdTl6V3Fn+VtPmen4uC4SHy28rnEhLiVk
8qiPz9FwRVLzvTk2zZTHRawZaJtgYL5L8AxEECKQaDRyikW41e4pvRqWmS3khbDJ
/sBGAsJuBNAcX/IhQK0mgRA74ONLusLf+TVs6ReKsL6qYU+lCYOlg/iec9xM8rR9
fSqVb9J3u1Ccq0Yh+Kz0+8E3VuVRKBJVIs5s7n6AdYvFySGDpqHaIqz0B9hKosf/
ZqvrUiwUEPLFz62Qxy9W67rXx2fyRBvXWB7LrbBXsP01zQlzUheNxLnUvdsbTe6+
W3slvecDj05rfvosQ988xN6AMMEyuWlMUa6s2mCwFUzdFf+zEtBbm/p91jPiEPTu
`protect END_PROTECTED
