`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NrrT66f8M8gvWMWGdKIBy2xG/bFM4n4o9uV4pbs3l9tQxr1rjFLh+B8w09SaciM6
G/ZahF9EC5wkI8n/U+Zcg1tMYgPaQsMycZ4lGs/w5TckEXnNv9mqG8w1ZmQHw/qt
irACakJO3r1MbWtwC1O4QJI5FZwDlPr7RKeJgdXqab3QZvNgvrXVN3jYeAa1mUp8
1rPPbqw7u3Wx3T19WKbS0EYITFjh06vmlCZ5x4q0nSDdgDvWsXB+0tCsjaFdxbpP
Zzp5VxcVz7r4VPnQVufRbMKBF36IdU8jO/JlGjJR27w23fiDP8ZY3hJGy8Qv/hw4
81BdkOXzG195HFbmJXGWeNSWhUOmQJ+5b613iIlKlL5oIf7rD3CQdVCOPXgsLLWs
JLXIkGRtH0bvriXSMM1Z/PCKwH0IkR/Uu9EWONsn1dkBATofICW+dEJro85iX5aE
0D5ZckuAgMiAjvnMauDgIPEkgSBBZzj51h/cXmaRoXFay63yql6kbi1b9MVyPQhL
M3QslKWB1W8r+3ghwBE/oOMs72QX+YluFb24LbH4dx9CgljUqvF+SV2HKqjGCNAf
H1e6SF9uGZBaq8y0iqxZgA==
`protect END_PROTECTED
