`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0sxTjuhTu0d1kYwMVua518kXFmCKe61QxReL+Zmsr19Fr5/57X/zFQ/QGvNGiKAh
Nrv9CRzdZbMPjd3HV6zIJMCd0dK5ZEN6Em9CEHpgKnqDOmK4NiutLdeQ54m605gB
fS+jKdWKpTHbgMj4325vbqrqbgvV4mUujT7O1he+h73f9ahDr4DFS5sZadRQDjbO
LwcxNBEQZ72+tdpWYkAs4RNo//AI8IIjHuUrRQlsBEv3AOXhpkDyNDvGv2sS8pRY
f2hLpmotZJMipBASlCiGZWoWbB8mppITBx7R0i5tKZFC5QeSS9Q2LG07BbDbYQ1b
4ZUU25TOvBBXKBWM1bq5HzPs7WN5w3QCCCjr364MeocUXXB6gXZAm5DxcheKHOtn
TYXn+AUw8JTf2qJkrdq99iz/Mr6JdFIKl0ajbFGmlZqZKymY0M87C9Inpq0sHInB
6cuXXtr6YQPzCIKBU0CYjCZhEztA6RWcQzUanRlrPpH2X0ls4VCEGLlnMn6LI6Oe
oeDn0LF/zC40o9iaffDQoLoxN+JbkNJiOypsVXyMGSP56kjLzToOIWigvziy3Nm6
DLHcb8V9Gc42XK3BTcaBLw==
`protect END_PROTECTED
