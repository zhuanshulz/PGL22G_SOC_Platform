`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YDReK1DSwSB3HxELK0sVWytRct/2YgfmaCxke2GC3KjjFP3wWDBBb33t/stUr3Pq
j6mOn0P/ZIRiShMWdqo6GeMLHAB7wW9y2u/78kuZ7tI2vfKTMxG6JBIQuK7+vSN7
aTOzMbAwLAuiCIR3GV9UrxEqzbhpA7lKPzkq6NBnYK73Ay+Og9xWu79I/P+V09HC
4PGD95BhJrCoyArHNg7NKohkGKBawcPrXS2AZT8oi13iXizO9RRNmh0bHtCgwwKu
csLAkRz0SYK+QxMlC+BY0hdZ1XIrOj3Gs03eo2xT1OyuFK6CDtzoDNGSzYHtT2Ph
qYGK1jFKYl8EVRKjrHt4APYBwu4RaTwZHNmdoC3hE/c7XhiJwIyQ4McqD84ex7IH
Mu+RNRiRcH6LfavbxyXZfIwau0+rAXDuYbrGEqXKoRGRlKRuZPnV9wm3tu4t03tv
971UTKuYrheol02z9Qle8FWj4xB3urUknNBcooHwGNZiOFTekLqz7mcN8FEg8hU3
aLCnAxQmsep6rBr/Oba0iY2Ap4jk3MdFV7jiRa8c8YIuTNMKDtkTew+O2vzEUe5E
BgtMMLhepq4nJ9utgmtaYYeq05+G+o/fQjiJzIif9cvOGU6THMN1/j2jMxrQncmp
9W72NLUwPWJh1pVXL8rLonsOXcuNXIGWkAuBlNlPqNbpsBG8PmMNh7fHCCRnOOQy
lMqkoiaSkHcVcDMCYwGsXHTqgDQU+mkNs9np8iW25oaC5WZVp4hvsVjMrOuUnxjG
b3QTaTXbT1FdT+eAQne+ZjSt5sPEw4PktKuWO3qcCc47uWQG9EQBk5Z618vRsh7T
yY5Cgz8Xb9NKN1W1XNpLHeVHHRTRZSFquJP2L74comIV1+yzsQ4JqFItSPMGSoRC
N5lN0eoghnUvwAcRLL+MyRz9td7gHBNLdjsshp7izQrZ+FdMYOq4FdNw1stzZ9OD
5X7Depj4/ZobKdVWp+4DpTOrTV0qxLTBj6lzo3L/f7JoO/l5XmRYxFOkBSxFv7MB
juln276rhTZGw7eEz2Jp/DYx8ZjS6+NKPRVGnYtqnECEfyFJnSSKjd5PCr2+gCit
pinI457433+uj8HSP83ioJURvlCweVcpgkJHZVwJ+a1Oja+AtDbPr7LYKqHXzEce
o8Pzz0dzUgGnBDCzAeDtIUmnU2AZUt2v7kdBIFzj94xftDWcpBpCnAkXo/gs9swZ
ncUmn2NqgyD5JymK1ROOZqJhp7jeQBPS5fgI5zYc1bZjGnS4sUje1H5ZXl6Ev2+H
j7gOlisZddEq3x9FTo0XmCMLZSgOtmCmvhPfLz8FOd0RH62U/remozME4+12s+qP
mHJnIacB7vRIaFF7HhpkqCOczoJY2TBwAyBrE4Nlq/LFP2EGdpcBA1KQcGuShWOQ
ODES0AMLUZ6rIakeQONnU5etKHbpMByUY8YvWgSRsmiKz/b6oEQsLKRxHSfvyays
q3zwN6WgwfrwFnmaGuxRjqqqKaUknbjqq/bBb/AH52LBOqOOC1hcOdKAhCXSjlmH
iXjX4zYQF7SfEKcoEA5vae27KvnvCebcj0ki2cAlCYhTigfMktO3/T+BXI+HxJ5w
fMJYfel3GiuGNe90+GWdGPjmrPym7Lxw4Qix0nbmRy352/dYkSu8EaaNyeaOKxMb
IsCDkYKIpa/YbX/oRzQ/IjfNPfdWX60Q3+T6sACJiyIjrZYdLqlNRVduungURSnh
gg22ooCI+hQkGcaevO/kpM+c3P/XUopsJess8ubZ7dZvb6i4Q58u/UH942QpcY5m
ogMkl0db7CFR+E7jFYeuQsLKthz1AlGaeuByNCXckk1RfzXTNMEcPaaHSPr13NNL
vjt/WmehfgMbgLl0SjdsX2WAlB0dDRRLqV/LZOOMtlpm8pn8CymhC8+XyzjSae8B
/dXcOK82gRgikCDVJG3jclXn19hGbjHRtJEIVfmaeJbf3bS+ZMB0rrc+aYHGV7+h
pIUhaqqG+qOFAdUaLTFO10gXuWbi37+AMfleDLZCX46HjPm7Bx16nqzt6orrVw+a
GaDARgTuPvxXev3dZtFc7R+kJt7k5KhucfZOUlHVOY/PBW2IOcC8v93KVD+gSfFY
6tgQg23fVUvEVx7+4wFhVhBnTHX2K5nHd+vkXYLaWxGElErkftuM7SfgWztGtx7U
1QShpkE0YdQqCBrtdP+t7j9OOrOTxgtQoJIdPLc3ubTWJQX7pVs8d8/mlzb+TYZ3
DMeiPrSydJjKRixk7gQ91189pUrSzalcstndBGNaX7v+93oaC1SVO0teFUjktXtF
XY3qrWtyv0Ajmi2J49dCMIPFcwPqIr/x4XPXvqU/+hhujL8ZTyaRLqfQsXT228wA
e9OTQd/zaZqcuUK9ZOAlFkWZYRRDM0yWstdce4satK4jT74XXBXbzR1YB9n0r0b1
hWQHb2HZfGYMZtT/EqKP1t8Q1M1H3/lBtM/pEAKIDeYkvpG7CQTvlQ1687SuJQt6
1pAPsYs6Nw/KLtdfOb0G99Iw0OTpubvnb84euUK0AZcELLAnabIBIaX4gzci/3/8
BkEtVmJnzMDtJVVzo3OIvJXP6RzqOHOU3f7JpgisCAP+nzFq5cGxOGvYJN2QLWz4
jJBAo8BwBySWyuzSIKXFjQ==
`protect END_PROTECTED
