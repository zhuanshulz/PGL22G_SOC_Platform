`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G6Y4r5Azdfj2cMRfjpzz1bgcINvRJ8Fl828yIhhc9GtMxX6Ze3zKYQouRXkz3aKE
2yfY4nTbin9nphOxa3R9e68wkkIk7yTLEE/hJ6IV78pBhQxFdugvQPTI0H6RR11v
oq8glDQKTp3v6xgLpXiGtxy+WWtz9epo778kEd4cuNDSCMCXneT0HL1b51eAtOmZ
4Ltn9Q6LkwjFC0E35TQtPKC6mHcop2UGDtjd8rEXtIqekusD39XYk5VYJmwavvYK
b5J5VUHG1xspromQ6QW4KFSnaIkOHQC+a2stJOV9E1YBn7xbCmBvkKi6l6KiNjrb
gPXb799zmiHmLjdwWDMsAP4IR/GeMOSRWPsFMJ7dnHf4OeEyuGPlXfm1pfG9N3nX
27cMsO+ihujWCh1vMsaiqoUyjNa87pnpLI+SyijBpKDa2Xbbj5UfK8LP9FZtb5a2
mMLPtotHBa7iin+AQYWXXEZcTI613FTp1+4EBWoSx1VLtU4RPrvvKmpHFdJZwpQJ
/kWGYWpzr9U0vH8XzTeQnPLNk33Rau+aw6DfqefULV17vusYhHfrbEbjUOCXGijy
XwOm0f1IZCuE3WiSvbx49YNFv1BbpboNJNdrKOFLgWbXQQrVSkOutDbS+XcEtMc0
zSngDmNAe5vSO9hHfnvWEE77B3VPkasobBDXCccC2Q17L6SduZcK0+cKqGpB0V+w
1/X7JA9+y2EekPQW34IH+lSkepKRC+vX0bzVb2xywtvf72nQmgD+UOEwokUCdEDp
QVofkRdsGTBkyskW0OcOxKKASkcqIHcWfku6yQqhbrEnNO6SQqFTjegCL7qkic5E
D4wMqBacuu+xkxPQXGIXDoc5w6HQ+UInk5XFk+3MoKVd9sezliTfE5Gg/GWR0RN0
0SKaMxnfgp39WAlkT33jNV3mb9TEN9rJ9hautzPE6OLwZ2Lp/Q2SYOfCWxWtF0x8
b807fq3+t7Hk8p8X31zHdpHWZp48A/ldKG5X1mEMB8cEkFGaQa03POeQ3B83XmTD
Z18vs06dqt66HVpeGIUJFuvFdSczKrQvp4ksYLimrQp5MaxSyqzML7ptGdWTfY/o
+gvxutStiVV3BHgl23zWdrHP5znDYSWv2I7C41P5pnzIbX7CLEwru3abZsRpLVPO
TmUZFiTsCXIgOMEkEQb/mlItlh7PHxNaItuTJTYc4Y9koms3sKMwcV+U3AxEjI1K
RLDhuYSPZk7pVUnm1gZvu+W8m5nc3FX2BKEmaTZHqM0KBAvRD9MV19Q3Um8oWhSU
Hjl8R4/LD9a66410xng0b6Mbl7XhGOPOevqI7SJvJFfmifa2zs1uQY06uo5pGjjJ
hAL8pHSbkoAt+wa3iOAgBqtDDdtfTDrTy4njjBEUKsMmAn088wEsw6Ad49DDO94Z
gs1di0F6nsSTqAJeFKjkAwWhrHHgdik+eZ02tthVipN/J1TCiFg4GdTNoCNbfsLU
2UPrIYqYaChoM4arSjcSSJggecCS4l5i3IP5WZIj9uNCNXdFkQzyVvwazywdDIRN
RtekntOOD+RrAf3R3BcmyNI38Bq767FyU30pCj0QagA89pxwGv3/KZFwz6Sqlm0d
cIqVGerVCURXiqiXTQLMMlgghdHoyOP++oXQkDwt/2aPjfDbjcuadyRByP+EilX4
fli4S0nBXU8x7fixlrUBEa4Zi0+RVBpT1uqofby9sCz8CImA7iEW3OkHVedB6LU2
OFbZeGbiVeqmdyi6GAYIve98Il8LTmWQONPHoAqsX0y/Nm95iLMrl5HOgL2TJLCk
EfM6/eRCak4iWMJ/mq2b1hV+t8lZhP6Eaxz6wTrt6dQe0Djct2TeCTMSeKK4ZfGD
m1dKngZQHVOxBAGdenf9cHFydZapgVynx0OrG1ZxsG9tXKz8mO2hXpGmeGLZbD4Q
flyhRxnHTL8zBsP1TiTgwanN1Psl9Icq2/krpPW9WY+e6Wz2itJ6UgW6DoLkvy9S
NHKVqe3U7W33cQ/8VrDuHk63ez4wCsRvlZZADOE0ueCxpT679JpeGEhCFKIZGyEt
F1sb8c3DH4PyNKZl5VaUJD5c0dihoHIy9Lbv1242QdcswFSty34eEHv7b6ZvRzaA
XOyhb0h8tHqn3AyPIAVN96aa/ZRvDGOmLXUyUhnlfgnrbUheKceLDRNAWHDVDG/5
J1QRHEB5T5Suuhj3k2UqHXmD2z82/txKARY7ZS4BAz3l9IV5ATYihHQFx942HMhH
Kd+WsslTILAHZiIgVuVm5a89h86uwPd+vlL50BOnFIOtDbvq81VYK+E8K57KgQd/
bBX5dqInt4Jg/26aCxp7KWD3fyJ/IsaHsK0dsARglwYL+zP6Y3H5E93K/4IZoVSY
ircsFTav0rQ9AkknAocq6AoknMb3r578ILCNEibDrsgpsANx+5jIcX5KkbNvt+MK
mPZkLfbBr2Tb1mjKeYgf+qXQtoyLv/6NcD0n04mMwmLoGKeqo0oJcEqz+nbgdemv
ebYk/lEgVTkJSmMW0Szs2UlvCHimG+PC/1V1BhslW5ejtkytNjaVNK8k40rwbWFe
J64Mh55g8JdJcQAbZSoU6khYIjPn7QgBKBsU5GcgMPhM/dlvKNOw9IBCy0FK823n
7+4whpIRC3omHQjyjm0NlIYxxQCHdkOa7GqFVDVhpyoLsCJs/EFapkeh2LjmH5sh
se2j/Y8aArFxmuVZMIRqJWlTYEtytN/wxoRSkdW09y8BWY0OC4AqQ/MqLGscw0W3
3pPnYAyrUtoLTqKJ0emByFCMM31fdf+ImNE8QYw8e0LnJXRmKkQj7Qu6cd5RmIlr
UtiHeDspOs/0P+u7PXfffE1xo4c+NvBmTuG8QTlHYbITE4/8ZjQjvnHK03kEGNoo
kEHg+tu8bCNTpFjWNGLuwymj9lkKWJyAManKW8Mh4/U0obGLboiu1XVskE5+gyf5
Mpa32W+bcunh6dpac0bAcPl0Hbx0Hq0oawB3p3I2p0UATkqwsIqd9QmUnhFkWIE2
Du8X3cMNoIZPo6BlFyXEDQ1iucFnVH3tBcz2AJGJWcS3/H27LXYcXHE6VLZtU55j
EvCSEoJbcXG372jNqiGT8NuNLAFMSFi1sYQ7lYnlZ+WgJvZ1Aa4a4+8F1Cdz8pZ1
dFImI4X/Rr6qhLjP4jKo+YpKPFY4fWEIjThzyhHHddOkZE0T+8YAS+hWF5lqVx78
h2fLpNiY+C7ssWN9/N90+dIHZJTTcqOVuG0GxlIX9MHrZVllwnTY0Xm7D3hY1FcO
w3eQxgF9MSs7hu5T1cNm6wKI5aaNBoxb4I772F+ODGjnDil+wgYwQovmeptS42ni
wqe1G9nSjPdEhXGUdhS4hGTl1cb24HtBlb5KLWWb5nlSwEOan4rgo60D17U8ft8C
/QF693kRka7mvQggdpjdAc2CAyT3NicWdaqOK+mEnn2On+LBdrjKjWrKuUxWt6+i
1O4nakk5tOmL0y0EvT2cAkABWdb78NhxlbUpSaLHrQXMuV7MZgRIHaETw7GtUj4V
1jqNNjF6ODjUx6iAWzTypgQMXZ5KUjfvx8TIOifm2X38OukbM1ESDedrIWlIRG0Q
8+3COmCBiTzI4l2U+qMZQyx9niHyBmKWd5d3tOtnQESs6rzutRq5ukIrQHv+L3ff
n3sJQhP3O/fd0+iWNOQ/LYHt+JGXhls0LHVCuTbZ3lO1GKfcupPxFBkcJQoA3hsb
FhPOZcW1lvXx4f3YBMmnGqSN71vlpPT9nTWYbCyML5K+tha24pXQbnPI/rkakI6y
sZDWaNXCtuzaM3z3xbaadga2iX2b/12k3rL79Zstm6PAYWCPUEOrfV9wzK43AdHS
yix2LGwmw7UH1ueYIwK/uDH5V7AEr5AXo9YPW3GphfK1TU1szNJgYM9n+iYXWnww
ypdnoYhE8vSXPTyymatLYnSN/P6pl2STQiC6bESGSCDNvNX0TBN428j8lW5KCDtm
ZHE0/+u1P91Dkf85MW/MeayteoK91e7Bos+0fCAoKYDtsj0WTDuh/QuCC5Mo4wRM
h+HSXx73mZHwiKcBWLzEM8LQOLxNZe6r0WIIhgHA28aTe/c20uHwPB6GfoEf1/J2
DxKYdstbh8UYBSvNmkpT0xOjYan09nO1x4N3FQt3yMOsj2DQHSoHErgWhskuk1un
1xqSyIWqiZhf1YoCitzfS6wFZp8ihe3BF0wlD1tu+f3kfe0yS98lJN15odIHnlXZ
J8l91SLBzesN95LnkVGA5ZUuutzDYPZXpp5ZPeRCfAHZHDN6FL5Sck3uB9TIe/Xc
J5Oh3rA5RMzy1Y4kF5w4POh8bk+xo+QBRxKcbnF635oBs4DLzAnkymGBDFQDvAHN
qZgobRbSQrECKC488jhl470MrppuygivqZ8G6xMcoU2gMSzG+hQHVBtv3ilMXTi+
LzriGP3Ya525vwNXk6uItx6P/UyO6XgBp9SPrE+1jRUuXP40EUU1OzHUtadqlo5w
AB9cQTpaWCLm1y0YfRwtBYR1g4hpYTLG+MIennylwPfzw13Rp4XEnDSS5Za64Vm1
Rp7Pm3yuY0YIhmocyKQW2pHMbiEywdJgmf9+Vc3kuYI+35cr6MSfW/RQ61doi+jG
lics47WgGs11AN+uuBEpFyQtBCIUpRYTSvllNusrEfHO2uEv6h84WV72j9aDXx5g
B6I2mCxDl3jbiMoFFoKs9VkrpFg+ebDeDk5BNTeiH+Pu75XBMzw3a7CwizbN5fFc
K5zljHXLTPPTETeQLsQPjMDO/KETUulzxr8I0fAEzBpadYUKFQvsISdSAS34Yzbo
hBaymGyQSny1h6oBwp4H+3b+kx2lsJ3wO/8brJsM2z3dHA+e1a0H6RmuTgPYpCli
/2xaSQnvTjcc+rjguM+TeYFVzaib0K8A1cYmARh8u3JW2PyF3K1A8m9YVPurFiY6
SJgvukS4aRvp/KVrvX67BaNrBM3b8tMFB+au1SIHXiVUeS/VKvyWs+dZXgyYIBL8
eRPkqf/gn4SGMxmYkU5EUnfExzbe5ape9MQNP98SL9d34pE9PvhxlpNk3qgbSwRP
ay9KN3HteGEuPDl0KRn9kdITdwjPCY1nCiHnRnSnHA77iavUEZ3FioztkS7pfkg9
hGMtVWkRm46DxdwEkg+/AfZ0nbDWFDO8c6resZ1sNSB1fCSztm7aqEn4kulfzuKA
apC5DDBu/Yh3YEkQOwVqswvqB1eKMiBnwOjyYQZPybiLMdvKVXs/BwTr14QoMuyH
BTR3qmB26CI86+u84yYLZEv67o0L0L30HuEDYi4UItmJhcQqevUU4KVlTT2z+kur
HSGrarO/E/YTeDi2ISemOgXQ0VFhlZ3gMUjG0t7dh3+GwxMaw9SgfZ5dZF/NV+ED
St/fWr2OIDwdYrJnSQoxitTZt40zesQ9tAf2Kx1SpXTaxEGj7Cou1vO7VFLuFd0F
/8ap7blnddKHfPqX7+nEIF+Knof1l/o9DD+bCaZx3gFsungKbg3Eh2b6M3ZxQD9Q
O9irzY1la3yKSuf67jYnBgl7KMsfjV/FtSfL2oO9erEjpSV1JnjcQe7P7tO9YO/V
l5+Z7OjMV3gRhc9+Q/v2iQqeN63X4ifT+TzeyEdpJsmoUElXMNdL6ljKKRg9HyYJ
ac/N1BkTJl+39kzrZXhSCbHQtZZl599lZq0rHQ6UZ9QFYER5JM6+XGNJXbHeY2kY
wda+akuu2QgJ8SxoArkF+zdpuffTbXI12pYuqbEHUCs8i9jEPSyf07DgdCmI3oC5
cVlJP2/ol9BD3/Zlic/GJW0kbUN5/U8iLOP1fOwCmVw1j6RugpcGmyMgTxSyFjUH
Xscp0bZzGQYoTcZBF2zqgqjcHK/j7PkM46Sxq77qX6zEI3YpiWk6Z5VbBMGa8NUp
XrYvqmPCcmwUveOZz7+MBO6rDZSR1tLtRoER5tfnk8x4oW1keUV9n8sEtd1+Hdzp
9UhQkIG4J+np87biTyVWEirdK+stMIEmcNCc5JtVrwSRakxCMU9aWg9t0KArrfP3
4wA+rhjQvDWnQ2LIjAJbTPeutdZ/Z2vYotYWaSmq85rHj5vQGKrGwkBTh3J6GRK5
DyoaRhomly7MwvR8zvnuFrizJW5RxaQWfbrl2lSI0E0/qQY4Xz3cAesMCErXwJkX
BS9IXGLdP+sjz+zhaKI2ysGKfD5PFi/P0DDjTdPkc1UrAorsU/08LD/sNvNfpS3Q
0hz/ZIHbBz0/3pWeO40hntPG2lB/hAiQtOeXCv8mZHOSebca0ls9ZdqTz+nrHar1
hlbdTBN6O1GWocaKbBD9fTxULxU/Bb5oirjV/6iFooe0+WkT5XLoOJ5CjWIGca9o
90bdKLhfAHLVUPrQ+MxHkDU6Y8o4V9ymECKYW0IAFhk8K0g1EzmcaaiE/knPE1kw
GMn6askUN/S9oYQmf1g9GST63IS1txI6JtxjAPLjzwggUxH0t71V3aVTgGQT99M7
5z4zDDIbsaQzbE6Y8KBSoqgzW8etAEoMprO1tytu+3qP4NLaGCg+WAOi8y8Icbbe
y9Gh2zr2OW1MyXt0L/BAPukHj94uoW9bsod4QUZZpwOdLmj0Uv+IFUcFIOkqh1fl
BVqgH2baZLX2bUe0POrpBHQB/Xnoru6p8fBrQeeDF+bt9hi6MAEfEkqS3bcT2a0u
MERweJGWAEsF5GSE9WSDefdL2HlEYhMU5FjfVM/c4fFedsGrJjSA0e1JmCI6lcqB
U+LE/+iE5stxjoR2kR4uA6VIA7LH4JlS7LcKLBXmMHOLGWXNz2iUQWRqOma0k2Kc
UBdIPRMyicZUgw/teKBvEXSKWcatITV/xP/pqUrs9fIZU99ZTS+HeG8QAUfHLdfl
iSeZ3k8IFfcaAP+8TmSA+lG41uvSZ+OKNiGSP7L7xR31Inxq/uOnPng6c3BVvwTO
znbe6PcoGt2KtY/7K9rTjMekU+m2iZOfJOm2Itcdhw36CqdNGY9FEoAVJavYdG41
04fBABOWMhOpNZWv2Xp+GXE6aKx/h9Qdo/+mDcXAb0p0kjx4eaJBld0qNl3Px3Zl
COtvwMTiUzq93mP/ySKtnUyXBc5QX9086Zoniwzbk5/0bu+REQorzjOQ8TEOnL9u
oAfWpuoL7SWPQ19tHn4A0vKFZecLiOg7wFLr7oNdJJ8savEcotMDKZV/dRhz01VG
lbzuW1dwY7moupjn/ADAfAKG8HMo/ITcRb0hr0cwxamwpC/sBbDsb/qEHm+H9z+k
D2h5ldOZChAKkl8VDvbtlGI7srVW6f0XYz2rOADX47KIUJGX+/0mgUC2cqZvIZuH
EIInZ8ybMrH/c/nap9pd8Fko0f+vh+HPEO/CjCOM5DbAhNNH5Q97IaM+K+WLVt4i
wbgrO+XTUr43rRt12Fq+sX8EZdA2VpX68iqFo1Y16sxnnTAtDg86lcsYwHtLZh48
M9jA/QW88PzEJIcitsfRvgbH2XniPjXiV5hhGPnzIdKJhVsP0q51OfmqyJO7cfGY
ayv9UqNDpQ4RIbATLgCL7B79O0/kvQ+Eun/KaY7By2JjB6kcqDRuJTjlGwSuWIim
X8eDkFdIPrto3EIj0YYOwFcAPhVwLrlcgmPz9fXG4uC7KzTYcL2HVplC3wcGKhfm
/J9Qh/0QXszfvzG64BfE47f/+2MsLm5GouCVeM1FVQqDNRY7MbtFEusSEL9AAHKH
wfkovpF0kVQ5bXJgP7K4obscCOvEpHDbKA9EtOxf//cXLeV3z4NreA2x9U+rtJ69
JB9fFOsM70cZVtvVH6gK7JPlmd/uqDfbFvWAMRRO6in8K6L9BlGRtW7lyR3MCnuS
N5ZIXTgn7wQyp03elh+02rVbXgbt3vYIIgasJQUkPb4SFMJknNNpVr9bOe2Jc9I6
uGMvNkYxqHz49ZUGALGHcJ4M2F2AFylHul2NGf4a6qpkPPYzubPaN2srTKLzJcUT
0KKZ5A3oeLXhTYRYKtDBVOgC+1r9KzuOogD3bBHFiXBQdbvjrR9EHbp00z6jTRfx
GAo7OH1qUIjM6lcVppTErM/pY56t7yi65lNU97R0O7CfMB0O/oV5Oq/KBZMFU9Y+
8s7gvrGwridBZpLFqjNfaXXW+/2sCY5knCU2Y9q0Ap4A+h/DHU0HSpt424Fh59nG
xBMyhZP2+luiRz4qIQKJks2SQc+FBd931JPxO9QAt7DD4m7cMwmnwSaWEu2F6bTQ
z4om1y3PUHh5M8pben/B704NLGrs4cmZdnSGcQR32h6XqlkBU2y5lU+QwUg2dFJm
DRQJNklHO1WsaJbkne+qAo9/5ndVbIhm41xR/F3F/AE7xS2pNOMF9D7KrYthGv+v
dyLnJVwU7KJuB132uBFlqNFzJJMjk8yzIoMiZhmVZOsg4i2H9PjGi4U0rWvBQjh6
Qnbl5zw/UUI85ZWeq1JE417yKgHFC3FrkhF6AWe8lwJvZMaApsZNke8Ra37jLutz
yIFVPZLw/4NHCb6wM4F+rhInt5JysJPKfh8l4rDLmZ4Caw7DRXtv6ToiH3zQUau8
/FhZxH2pQPLPS8dmn1h7WsmjgWmQLaMHY6f2vbeSFQB4U5Tl6TIds6F+SB6bglJY
H8ugPWQpftSUhYIg0qLqczTgmbHIVnvqBqWWh+NYZGe54u75Q+jOWa0oYeYZ/FdZ
ntap86n+vTnkuBSVUMfeW/Txi2qZCLbccQiQg6kkfNph2uk8WWdV5bMkdKvzTkLn
fBkZSuNfcGq/kzTeP4H8YrlbA8VUfvLBHUq+V/ByQ2dhXsquqP6fBlT8EZWK8KAF
XIuJyZOkGT+9qV78uWm/VeGdiIL/sBVImscbuVGjr+tV9u62eaSZqSjlHr1J415p
iSckeO+85rdQQJfC1VtzKvvjnn0FB9MeOx5EedYQqK8jcxD/uUDID6lkT1MfcEJv
I4mo9ISOr3dfgOHREpITKIit0r2IeBytZvPmkCkORxR0QI4OGpmejtsUoU3xJ4Tk
E2UXYM9IBgHJC42MgxrM7oQF7v3iCvkvS3fjrYqehYx5BkcI+1ot/9gG9YfyNm17
dJ1jCsXs+097bzJryIcUwqTVSD17tY6dKyf55Pr6+VgP/UbYzW7/NZ0mmJv+NuCZ
Vd3k4Fe5djRSj103RqhjUCe/SBqNnFsfcSm4hIbbml5uPV2ZcPHwGDrj5s0tixkI
rWDcWlhmBXPdm+Gvgtmq89QOLrQQ1gHoZUEharW7QyH4G4xln3zxBAIVzAOap4UD
y/XHjIS+WdazBL7x5jMXLp4jLJIK5d0YvVY/Fgh37Y2nMAf3ZXhJp7K2gCBFDZgO
lp8PUeQcNa20CRKqfh9LGSox13k0m1XP2lN0ryOLA+U9DCGPDh7JbDM5xADas2tp
hRMtwYtljQVE0Q4C8hjE9mcJeZIBy8F0k346MikEoYEGTrGumIQ+2zYr9ZJvTUtt
b2QSMvLk+/4mgJ0NgzRoC0K7lvz9l1wbV7MOR7i9BVhNTxSyM73fNH4CQKrO+xCk
qVK6jhx2WmfXH+36iM5THY85EEwMDTbsJuZB+Y0/TpD1+E8F6NKRpAZB4qKyXKyN
hDwqHexsN4BwpelkLj7mPZnkwrUQr1DytF9UP3QRUFSOCiczEfKchIDT0uTxwiWM
uoEusnX6XGYFCJPWS4ebOdJCctKynx37s0eGwS9GBMimtOc45waUQE4sPyNFsshM
BJj3f1iTKLV3St3yn4HQa+ADxyYn4sTkDRLogTwCIgnTPEAVhdI06WoC07HpyU3I
QZ/YQdUvC4QJ/n/CXh0djN693MJdE5x5F/k5S3vA5C+brk5qjmIpv1JzKQq9TgMu
a8Ytrwp9zMQx8RLtB+CQv2DAgmTUQJ2tCR11OMspDLzR3BToAm/Eez29eiqfO3Ve
2vlQkK6hy2jPfUbkWQvVcJaxVkPvUk/XmMTnzEUAsTHaPR5h1r+YjM9mFD3kFWix
VaeEppxykhDTyWWb5NKjiFIMsKSC5TJqRVHMiINh6DNwCMX17bEVkmyruymb2+jP
PZDxNNuSlkD4odNXiSaXRqg3Mwn3Ui9DWZ0geHa1dQH/d8mU5p1NqpGug+Tb+VkG
AamFK8FMarsf3v1TKXGfNaF4kMyDPwyFfaEPI00QXGg8F+6Yksp9K+JJ+4Pc262e
GNHkTuWy7OcTkySh6yN2xfgaVfwUdnUENpyvp85cuon/S9vB+Ij3catBYWiH1xxX
saT1lBufnZS2ZmHSCxkNDX+weOau/k2oiANPTIsP9QWfvy2+uTZbkWVzhP23HzYO
6/BDHLi4DCTKSj2Z3xKncLKUKGsq5WZ2qKpynMAq1fA0RMsvndU4h6RDFVCc17BO
gQqgBIAXxGxNOcIs+uSPZczLWXzFoDORS1qlKNupqc70OWHIU1YqUtpeazCqJT7+
ZzVsBFY306cc3kSEqnsoVxA/Nx6nJSMIhURP6Syin0c4Qebc32CzfcwLo6jsOm0a
Le/6oZ1EPf+rEoCQa1v85tCB01+e3asDUEhgy5qi2tIcc0YI42Wnp2EkGs5UBodY
7NKWY2EqfxZZ6mmbnleCMju34lgLNSJtiu3JtjEXl4kTcKHAeqz3yzMjsNpsxieg
M4N0xYWmwG5pFJrgPeQSlHjL6TZZz532L3msa1RvuucqUHDxXcI9pr6Ykx9HPYqW
IocYkJjRe911kE1ASt7cqf6LjsH7MBvRKg8cZ9UZ7uEdYbhjpKKFBR0iFMakgSgA
cszEGY+lobUSQsSHbXIg0CddcKk1heGl0JqHOWFBhhyVWJys381S+TWIu1v4o+Yr
QsATgmK+4glDkTvwlgpNBxuw0FThR+A71wpoH/bdfT45nzp7zaIAC+TTtuE17KoS
6d2KzZ0PUlsHdOUkQy/6J/+SIx7JWMmbBYQgwk8zGkYKF4bHlqicALNpWaKDcAWm
tYhprcNt8fveQUp3wvZnTzJKh07elEnBLVQ2pih/QQ2eALjsip97jd5oYrrmR2NU
W4hK+KtJVXpA2PLCUXfvEg7Qpq769qhVOuKsrfg92e4YncP/Qpw8U7CCgMw+l10n
+KIalMPku4PWOXG480TpmGvGSzIg4SVmrrtG4h7e1rNFTI5FqQOc3BUPvFFt3Qch
Msx3vsM2Gf88d0CDg6BPimHhFUwGyFrzznCSC66A1pcRFzupyQ3uz+hlK1eEehrH
yo3bEmjpUj63Hqbivbblsbbd6umptzr441w59VkNAj1UI5kAGbwl/RjJFpbgIcu0
86Ou8ccODvTKN64krKNHH0OhPHXDnIyi6s8skSeva0F4cnGT/Nzck0pWAxDwbCBR
8RdVEhfb7YPwmWG5OOhOCsH6ptf5xyQR7XWhzNFgp/Xym1OSGNRMA8JOHB/8A18A
xy4ia0MvZpx3I44fYBIWKItOYFUsqNa6vx52VS3/2850tWDsPQE5x9YzYZX83NrW
rL1rCqDvqkLvTNx+MTBlW+gEyHrkMc07WpI7NrDfXj9rXdQh8GIEbAntIpPKAgb+
5I8poZ+iOdi1axQhrhqVfJ1GKpB6mgyUBtZc7N+gdpJGfq+bd80P7PefJGqiQpPx
kGRcPIPDQaqVrO7ygSbpPmpqevBoKNlyiY973Ld2JWu+yyiASXbr3tYwDW70++Vm
VtlZP9KvqTDEjz5KlSnRM+Y9vo5Rof5kyIKobQ6c4Se74w59vnX4fn3t3y0JtJV5
GGbyvMaN2DjfRVnUSuHUGIh9SRCFtiYSoVP3evJnsslQVPJDmnFooPCb+nupk61Q
aDq3/KWIlN1q8gJhBQm/i9i6IGaxkiOiMBegO+QFoIklFZ4ruxc4SFApZYrdM0I3
cXOGwYP1OC0QoU8iVzWo5RVpQnaUVjIkpR1CdXLLlbso9j4LwleDQ5byjm+4i8EB
HZ1c7hhENEYhs+7u8qYCMReCRS+w2nvoSjGLyLSSnOVwNbqXY9JLtrkur9UzvBl1
CO2Q9uCm9A3Mk7YG0gRo8yH0MBAflE5gh/9uRzqdRw2jkuZfTf8d+oTZe30W8054
ltIIIj+0CiMK08+CES+gLEYrTDbFUBg6fcvkSptD5NU06R6emeIlIhXdowbgeR2r
6BTT7uoo5hA2M3nrDDWBh3oXrDSd23brzsyydtm+E6l5HR3F4p78f4hex51BhlEV
BlS1O3Xb9yIbOulu4xRWfKAeAV6CpmoNYYbceCYC4k3vbxSwD3NdJoxAlgi8CXJ/
Vu1zeFWmFvIamGkCXt4z1JNy9lzbVSDxR989F1Gng98cIexyiJG/HlZzIALloUSc
68e0SAGQZh/ivV9GTSRYs1nyLn77mnBZZ9rwEhk6MUz/7mYvDHxvrSfmxuvuz4Fd
bccJCuryAnP7MjGnDYBatHGpB9vmwIzgg4fzdWS9QKcGh2o2PTIUUmmQ33bnQelM
SFcoOfFuc+VkQFQkQqakzaJ28y2VfDJLbBp6LczhVQYu37gg1U8IHuR/jMQgLyRp
MoQr08VvgggxqaJlpAo8Vx60/TmaT8KUQcnR8BYQtjMPEvZrtU184xAIlj4PXoMv
jMPZenvcb/4MtWvM8Gdw5gN3cdWr3XNLglpGBDwR9Qk8Jj6+X8DpDLVeFpNedS6b
PmJe+gkkvp5eEg/xRx3dRZ9ucz13vmrH+IS3RXMZwdcK2cM5Hmo/BbjNtCGUvxA9
kZDUrq7sgWkAqm/McQYRZB1zTAT0qfR9aLozMAA+mD97jQBnomfOyL6J5hv+rfb0
A+tgtJaNVnoiGyOA9HsfdvuoimyZdMY3IeS+ql+Jx4yxxn0vPG7bRhMxbfK57Pi9
gDNIpiio1o+0wYGCLYPUUnHmgbaFj01mZtVTM8tibX1p5OAGHoKDO4SpG7jKHf6R
EljtbHn5rj4IoS+HNzivb3Qnst48W66DadC4UlbxTOUkwsN+rK3kf+V8NBN8YUZM
BFjHHeE9cRnsi3kJvyIlUhz86M0Hb+QigD0rGqhLatpME6LlCo5sJZbMh2wJdOJo
DxCM2KOVFs834AwdnSCQF3HRta5FwB0AdlVgvYHkqFniEgTxYOkb2t/yp6XHGgq5
L8agH5hSHxwW9Z19KVnn9PrgswV+6zfNua5K5t3ujnGTcaWySgG9c499O/I/pNeh
wtGodqVPGzUeG+8jioComfCYMlq87qs+U70QwnAQ2o8woNpBKM+vSSZP2vZFof7B
OkT8efHSOugfEQRU2f3fp17vKFh/71qeH0yLk3+u1VwPFU8FQMDCfl3MnLtKMp73
5cwllp67dqdoCz1gUqV62SrASCOZMUV+VpbxGsJTX7WihAbDjXq1TIIY8z5fIS5a
gWg2WzHgzzC42ZQ7RTvA2q92p9wCyPeknzboE+Y6Qud/ZK8mwgrsjB0ubhx6fnZe
tuiWyUqMEHeFLOxoc13OPOrMRN8SIOewHo+MHvmsN9RGhd5uU3B9PkEao5nxeYem
ICbtPxVRlzsePU3fR/UwWOtuFjX4228dNvsOJ07bRgdJr++6DIw9PgSRJosslgwB
wnLqtP8HjtlgC7dr/jNcB4RUCH8qiBEyAzQkly8wCNc7Y/JMV30v6/9UQUE6EOPR
FPHCA72gWaH3sa5PLgGDX2srfsUIOzgTPYNl5mU8ckJONjH+CAqdAkWL6tB9wFSl
OA8Ud3JvZhCj4D92RA8i/IEr1RnI3aDJNc1tT8c5SD5VvKfsRsFF1PFd6MNfOzNT
9Buk/w5n6B8eK2Fqsk0tV/nbEqTo96/59q/KAl2jvuPfYWaDi9EB7fNfqd4/XnrQ
eMn4eRCPYjy8ngirITjTw7EdMGVZHYf0HslWdgpcAS7qQGOp8uqoHgMaNqApfBJJ
ylS2jmxAIf/9nScPovCSX9AGuXillqpZ5ctYMMy7jth/zn1ycobm7seuwpghxMkj
J/eusGrCo2zdGyMSTDXRnX5fyG0CSPjszj6GQ8PH6fhHhnl45M5AlyCpHcsolFt1
6NskxN6Gzk4a6mBA2HlYfM4NfH1kgZlrMl8FRyG8TWBXFZpg6UxPHlOEGwR3mjEl
sBYpY7LSF03BXlSEZfePXlirHSqPQ18FynF/H2ANiaH9Xs6U9tBsKN7pdsLbsH5e
8xWjLoLBk27lo1VWwJBUEMwAu24c0LbpRmaDjt615eLzVSqVZwFUtYEAAojFVr58
fOsMRYh+CHytRkmqM1eWc1OhdFtyjDbkVRZguyjscsgjKePpZpkO/MN3ra7KY20s
V99ej8xzit+MX+Ox+bpvOS8/x9E3wIrUJCAjEXqhU1HRAMkf5lXn7BniBaxvn2TF
JElB6YqjhIwgeVs57rwFYp1TmyUD/XAGn9uhi769+Tz8uMBkt718s28tl1isG0Nc
Jn2G+7J29MeIA/0OZ/LMn6Dc35SsGw/PTZeM0Zrldv4KfuOH7oESBWlSlN+9K9pf
kHAoUQ7sAGs8wnvs28us7jTX9zzBv8gEGYFL/zGzjI8GcQzCFOzLqbUYaUKh9DTj
KU/58y+l+0OZz7U27T/XNDCiG/WJd2ojJM+ptax925CkQ9jN/KwPfwnGOarO9ptf
h4qLgeU1VLvHPwCmz3r2sO8iVBcIf5IVQEJ2ZixQ6w9mYTg7Es12iZ3YlB+zx2ac
eqgYzGMOLcgU67mc2DmSm7yVnzIGCkkl0LTWtUowOEyklAYZoYtWYRwjLZ9BkaUg
YEjQSsixnKuZS4O8plMIgwltJ/mKjuZ9OAWY8vNdqqEbvKysbTu0dg+I+Ea4jtqe
iAkmd2jTeTXc7PEEeIOMYWL8FiuKlDTVHLOfhAZ8vUmh7AHr0EAWjGyR6a32Kqql
2Meymm0v2XGtuI+syojCFY2PgR2G1/TBxfwAPnO8kJJ+axTRZDHjt/iHBGf6440a
f2zgOh4RGMNlMDuK0K431yM/fOa7QEMVkgaj+d1WMSKJX6l1gTar6GtNg0XpYCvf
oIbKZ4gytPw6J+TaEhBiTcdyJHIea+DpTqLZj6VTwP+309TSmIeycOh+XBS5P4Pp
6HxK/1ulvljlH8CYSzpElXvH9JqpU83PchUr2jxnq+VxonM3Am+V77j1hPVSk4vV
IbEhAWSyFWOEdCIgl+QDzjvIN6ReGXcPv5ziVUmDmACqIhMVaByUAkzaSgnbr2tB
hVmiJ+PngK4W4YQiLwirOgx1+xeUcs0tPvKOf9pniecimNkM6FHQgVtv9jXAPTGh
0L+dbWJOJFdZg+dfgBsBrWjbFW08W/xYA0+jHaS07pe6p8TxjjuItTyYedRtnKgz
TlsiI1aRdVxHaj3O/DnuMjrDSFhqF9L4bG6TF1rV1QCMOa4Bb0mG5kWjBIEJs5El
sg1lIS9ntG3tTUNmroLdnoCkXRTbsT2QcN5mal0F1kuQXIYFJ6fg1c+ggjjqRnB3
MsGUhfc0pnp3Qs0AsL4VbUYXIgp9sc0j0+G3ttO9AGoZLBRZ7aYP61+JVWReI9/j
PWDFFydrh9Ffz64O0bbuXs7w1RWPt5gOCaDQpwPuzywwpBzMPZmEl1U2626Xex02
547FH4jbvk+3e9IuScOj/jrqcXcv0MW1biz+QMRmFS95vSqQewsGvTsAtbWzhK1e
3bKDLTd1Yc0FIuS3H+F9Le4SvDMJ1ZOxpLcQu4xElZQ3/TT+Z4BuJOqAS5tFGKkb
voOLbZafRmbcZfe97YYLPP2FoEXszH5imf0jriBJ/9SX0WaVc7UZ+j1+txLqZlcB
/ltieqK4Xi2r3sJDT9qNS/DdZML57hnMEiDGQ/w3OK5T00PmG4OfK1tSI+/dS7CW
JPmFmSotuJNr/r8genkv6TJg9gOJN7mL2mcXQGGtudZ55t5QWk6oVpWfBneTcxsc
BPXejeWcUM03GtdIVLuWQiMvOghsS5jO0yzDvuuqxZNgTw16cMeDGdX3Jqh62LVT
TWuhG0co7e32MB0T4Mn7pQrQjkWVDJNA1oh/dUs1YNaegAxGYPLEMf9VUMOJn05K
GNH5ciXUSlLBcfGZNSbyfOq+FNL66afoMdFQpBXzY9JI0MtPe5cNJqaTyTmCozMM
t4qRM72fAUZnV+/W9xY3vuegO8Yc4/7cVa2pcA0zSkf4X2kIvHhbkz1vDXnQnPIQ
Xa0oO5GV11MySV2S25nUD5BbZOgcxAmFF8vkj4jl/27ZQ6PJO4upilQcKRvXWTtg
v75SCHC0lCgOQ2e6fPaSYq5zicqJ4cwdjjZbOtW7KWzFFtRIqSb409KrFEJ5MwFx
eHb9M+ZodvEYZZjiYsOxjcJ5bH7lzGlm698qIZpnjbjNYIQYS9LbKqgPcTo5g2ed
RSOK0pQhFxDVh3dUba7hsunNnhxM4pDiooSQP6UOkdKhsBy5hWdWNCx2txRpfdVV
p8uKq6M45Y34622MZHEP9ZrdkiP+YgJjJ3ZzIatEZxGC5xPHCsNCdAeWAUzo6qDO
NBtzqnY76aiPPUbTnD6o6JN+fE+nAu0ftUkqpMT/wctF56DtMKgifZQjco7JCSFQ
jS3Zh1m+PQE+bLa7vJB0ah92iSp3nYdo7fYRIQN1MRHKZlbLYSmTLhwZJbe5hLUr
Td8fJ5OIcxUYls3ZTmNsi/12hHilsM/ufmTWF4BbxApmOicGlUXmHD3FqTvLA8P0
gLihIH0dfJhluWZXGPHWWZ02z/vCRf5J/8Tkk2dX/pX3GoG9eXnaNB7VsV6GnrHK
JZ4qPJPyfVeJNCFd5GQGjQ0RBlnK0uKFw9+SFOx6XnJbyz6hFAQVaeIdUx6OqJAy
miUQdAzzHAZqfP70GwiNOmeKt+Q7b45GN3ZNGRynobbNDBNXnOVNoANIV+EyzTix
+GXD9P0FD+PClp8mdiDpeC+xMoQFkWPy4dzuGeIThlLkqYu7lCf7HBtUb8MZ43vq
dHJ1B/YQye8JMZXSrz3+LJj3Trh0oguyHRC7lv7KLxh0OnqPGrvtFM7It376p2NM
RFBd0/1Yrhqk1LXSzYuFE75uN8qw7+Rc0A8R1KsSfBJNSYy8V3nok2ZV041lui1s
IE+cCT5fhNvJqcjnueNbdvj4IK0m06dplU78l3Ir1+RXzn0bYGGnEzyQYPjJf2Fo
AyF4yO3yE4BOAdwu3FF7ABidphGNK0WQZFAgkEHOb8pHPh0WNCe4GHyvdsFrJkvK
CquRDJKBdDPXh69GOYorWOGL8qtrJfT6rcWAFNlWPoxEHP684vpq3W6DaIgxLazl
p40tFrSSXusrVKqNj6vKKbTGS3vtHruM63Ak5bmIGCXV0FaMMGvsunghELCS8iFr
BbAvmESTdWgjIsnZjxd4f/FUqF5z0xUNuIwbiA1BvYfKrTK3AgOP5EfyvH371nCW
27h0Ew0i3T9UjX7Dvax77UQhxl6r3XbkYuPVk/AyArKvh3qHS/d1GGp8/Fy/uzXO
IqElHtwSF4/neEFKCrCATP+fRJV9DTWS2vMdM+NCJ2QSGcDzjV3dti+Iu+kp4rxk
Yw6pE0hNOyDvkWulYuibsZAXOObsUPW3xtvtpKWkVcw/YSUXxT7pRHmsjNJkq5sk
or4PJ+1Muun90UR04IDqzh7CzxG8rcideH3HJEZhzIeNpygmYbd/BmJvDdf6BbCX
W8zTqME6+cScWW/Z9ePlF9N93d3OxUqYkq5Ueh+692qck1RqnsWNRZkC7zxKj0Pt
tDsuzyPsVPvTWVY1nsePIPoh1FiU1CE6bmNOKngcekpjOnB50GYbwb+IuDB9ZGw2
6T4yK02ENTvGWDw4yWm8l/3X6W4HUNkwqReBWruDnzUPjEnJtfHI2f0trhkAxHw4
mnvc8SBBVmVj7oEwPubZpdOYbrW0ROa033CiO9kTcmcnr0GC8kXZ+E169lt+ck5M
wZYW6c8WBMpfgUBapCyxM9UnBI2ab7efRHpy8xAFd0asd3c0DIxTvS4vIHbzXB7t
Czci4REka7i4DMPlwMSfYcJ9qJxK7Ginj65aXMLLos4iOR4AE0EDZ/1UygEkXmzU
OqbX0BFgfh1mVMVMdGCm9OfdKQDM/9cXucKTt7BI6fzKap3OaH51k5oPnNMCP5PD
1F0/pYlTFVVhDnn8r6xtYMlvhjV3UyvGuVQ3CeNEb5YzuZoI7MAP5HpzONVEUmwG
NtWR3fgy3YuYE5sIudoHyX7XFrw4AErNdAUUl0kgst9J3Y0kkllY5h8kJbelbGLI
WTt35OsphxeJvqryDl0AoeMxuhuCHanEBHIuBRKPaJKWswRw43M5mZCqQAZ8Q+d0
npQ8IdpLt2a7+8vwkICsfrtrEfMk4rCCE0FAQYSn0HEJ7Vvemh+wgEZutILxIGFv
OBUCu/Vi01XywsaYxYHX3OTru9H6dtU9mxQMwoewizgyYf53pPG5IaAMsO7x35k3
EvDfj1jL/44Qk+azaJ0cxyf6687w2Z512zaNPeQaa7P+bBfY1M/bWEuEHBgqIqUU
Z1JRCpr5PSnWPhoO+kewyI+ouxVQAzAB52Uws9sgh7GJRB8jRjs5V3fFqzTuHrG2
RhiiIfO1f2pm9hQHitleBhuhmeJvQNSkpEoPHRNhL/5P2P3FYicsvLKLRW1YS0qd
YSwkz0UiKZ0lgPX12LXfinLn3IRlD8g5jOyBB0XbDAoWxB/jCmTv9TjNCSYF1b05
nRIs/9gV3+UX19UlMxi5xOwkVU5F7XI88B9uoWlGpvjorHszmY8J9Vshqs25rhSN
+Xd6O+z2Au494AkMjg2kNZfXre9GoS1K/8ukrF1w3c3lWIhaT/rY7nnr35wRVILg
HdDTqjLsl+1U4cAfk8AhtYx+Sr7vbnimuLTOlM5twoWMX6Pjwu+0VNLEXqfBZE3Q
AgmZ1dUWQPXBud/T44gL9+J8ztpeqcEP4O1Tj2IK4RSKl9iEpb49JwtJyaDhn59B
afnJTqwI3aCjHnt5OYA1WE+JDVZGcjlXmz+Rfbw7pa81m1j/zw1R4xtL8zlQsLC8
Gw589Q5MRsgB4tnempQjobg5/xoosx3f8qBAEsyv+i2tZc0GyiqTgZ8m/EtuDZP3
3cF8QZQmZkMOOo1QzFxdJLww6qAzTw/wKBmrS9WMfPp56UFkxOoPe0uMJ9P2Tewb
zq20kl1daP9m10ZJUvrs2OXwjJbkDJQySJe5jXBJeE9J4ZSdDWKUgdzeFmbgGSKq
ICORrnjMNiGZ8RWtJ3+HyKTBDDJKkNGjHV+XRSgG1vuhD9DvlsHEq2DFQNaMEyB+
1vE+zyhVq2joEJfAFmmgCwjXbZGLvi2vj2Doo/x7z2KXlGUaMI5yK6rLYQrd8aTo
PwhLMH/+zb3ehDm/i2remIobTBhcC2c/wuYISH0rBcRlgZbqvY3bVX9ixaWC6RfN
BZMjIBbaB5i4taifiy5WGSQyzgDv88FgNKozXDMF5L1uGv6UayrI9Lgb+qLP2dQA
cj8UO7KA9/Sn1O5flN0R2Dx721n+EVYqoSPeNRSiOW7Qes93gXD5t0ODa2cZXX0w
34Yg1L+sJ0xJ9Bv7capfUTuiFW+j5QPn/JBIAW79xBs3Ax45UnP/bY51nIsCBBVp
eSufyy5IfgEhvj6dPgSAg0MKx3iU/KStq19hnb6mcB24+6nTD6zGvnKaslnV0G67
cYaZCAwNee78uK50RuhJGcbkiFuIKWB+Os9A3mo0M0yakkqefBy+6Euz6tyIDdfB
MIFrH9u5uX6R34641ZzBS3rKn1pixbdCBk1Zo6/sIJYh8gfI/YUSRx5+xK9ITYjj
0vfg2ToXg+5wZhm5+e1zkRxk8sYAAitHI9D4Up9Vpb0Zr1cOeGWsqzJsgLUX1hyY
waTUBsKJ3IeI46NU3m65rOTuCaAemsvjlB7No1oUossHhBdxpYBmgV5gjbSyYigJ
cKiUAaXSEatSEA28bH9JqzAQMY7J25JwuGpXNKI76U8HGmltJxcbCa5Lio3NmhSj
WLp0u8OMqfyv74O9q9bwYzvJqLgkYVRd9Ay+bsENKayzrwA1wuqcSMrOQ7esr29b
xm1YX4fMCiZ71LLlVSzBSxIzzlC0WhI87Eu/p8waitn9vO/uSps1wx2oLINpZrjO
kStLgCk+lqqCbynYGmVvWFVjJDzM69aBHQOUzARwookmtzAR1Fvd4vhDL1pefzX7
EzA9eU0CvjnZNoovIe6SmlSVKjryk5OM0b4U6M3h7EM19y3R0n0HjaFpZtjH7GRX
VdWsx3/TTubIZPQv5bjzg1iScipLw6FrTx/92SD0MocckbLLBWMrCBpQZyiw585a
Ipukvg64rqSWN7LAv+e9JBaz4sJr+OfTFO0N86G3czAfbm4EBREBbq4nXfN8mxVG
ydWIoo/IM3wta3CqtX96PBY9BNztc5vx6HGQx2Zd6+e2xz5GzuUgbxE/HF6PhASQ
XhH8ko40zQvSJku0fq2V+M78tnEoQXWKn7UZD5CBXMj33Z2v8nXy0BH3TlmbtjBb
hiqKPR76JiSkMjihF0hm3erZq51spwR/OfKuf84ihlTWfbVcqynbtge4CQ6y/pfw
dpLHYCaeZwWZEpqbUIaQHDN6FEkIkPLSaUQlxGUgJNLI9mdsUye9t58gmf/thRuU
88RYCfX9DTjkBPEFKSdHDYkrwGAKDH4f4hTuFuZBD5bopl2b66pGGG08Fm3S+a4T
h+nEQn9xdsdyN5K1qykhP039b+BktihCN+ICjE9z75143mEq1vpztZzjAaOMXEUH
JKEs34jdxlR+U2nsOzUyX7jFYkVp4ehULCWTzeeQgyO+SWNh0oVFnmzaza6RGC6D
5Pg9iZwnVY4s/XaC0VQNjnMldJ2hcPEWW1HO78BenhRQW7HUIpRAn48ODtTMG4WJ
b2AdtrTWii/iytt5VYSaW/vMtJNtoMHkLvjqwsS3HupsQBMgPQV8o0zs5lt2yarX
VSAJCFP5O5XZ/kdV9RPvDVcvwt9gwV1fr6s8r4H7o1dJTqRwD6aJapJiZr6qz/Nb
qTg+O8kvEK7WqfIDX6HQ/YEzY1LMGyD1c1q9R9CYJiOSRbimnuS9GTe6Alwn9DNx
XK2T3JodUrgYAZygH/83sdQ1Kt+Sl3en9VACsj8d+tdwGchDzT1Hk2N8cV+qyg2A
i5/ObcBQh3c4Pa9qfKl3MOg4iEFDVID5OrSr7+dhL4ARYqijcri1rO2g6z8GXY7u
C9f8fZX3ZvNQ8D98WJNonwehJuX3a6L5AqzdKRU+uS9JmoWZ6dotXvW1zT2mfkmQ
wKdVfBD/+nTjoAeq6oUEfCzZl8pE4sCUzLkTwo0M+TeE+e/4x7NndrFcfSqX+utF
XOAG1Xolvvkbqpb1MIV8ENPGNb+vvsHZNSWicxY1NoDjWjd9+X/hU7ajL//4lyZa
BTFU0Yz+r/bZDDoC6PYl92h1KW2T6O1qfuA3fZincCPbAeqEI3nqzaRVHPbwK1VL
K1aIqm21j9VAjNbEdbXrIPT2M45sjIosLp+8MMt2nR12Rwf2zO4R4JLjAnUcSthU
hLq5Rl79qnPmcpyIcCbeM64U0DRGTyvLgX9Lol7MU9xnTtFZJR9NP9UA17BI2xPf
/K7IEKaS3g6bhV9bI/PH1ASYBvxkoHsswMF446yWAKJVw/XA8NMSatXf5VE6S8iR
bqVtJghsAvcjpUK5kj3sfGMETVbmpwxbhQ8eRU4yOFEOYYs99Da2wrYFGfcN+M0D
xUG36NUnBSUCXP3ACSRrhRZfhLXZCCE5RPN9s6TNOLVszQykyTKOASAb90MljC2P
FHORSegJEB8TdN7ubQxDrqD4YP/qYFbErXbR5F8yPA3C9gdZJflbDtH4Ha3BMoIg
VpW+FZwrOMFsXknShKwH/DUwdFs1pzHcr1V1AaK9ah8jaTlZZQ508EvOcQIjUAC6
XXb7wrLIKsYuX6PKCTM93y8+bwsbVZdeZkSoGMXWBOhPi/v+e4xg6wUQY/jOHzY5
O2k1CgqOoiFxUhKtNTxmL7SqVlBwPQ/KAmtF7g/bZPd9UNwfTyZ1o+r2QscCjAyK
P6xWtLqTwwLwyjJgqwMk7n1qMbE5QlLLB8z/J7RJp0lXXULRnv4KChSfzp2TWXYi
NRPxwlBwMq0vJ6D62dx/gtY8EQKyvmwUQGasM3wfal1Ab0SFvaMkslqJ16PSylt4
H42m9BPuYngnqQjvOVsxn+qVS8gqdFVlMIQWckQBjlt2xJXCSV1qF3ZqRiXTwAjN
Dp1N21atxEFSPV1N8o5conOnLbTRiwyo0HJDotQKOvYbYJozExOV3komC+C4U4LL
QucLJdf+nqQEXQHa3g5VAkkL4thRuzIAIHX41tUIYQsRukADarModxbHjCvBC0fk
7qwPBSqOc0TA4QveAJM7XYE0mxhUD6JXJT027PVjHruShuynZDCn6cem8DDxznLZ
nkjUCZDRBI+VqYMDaZv5EpTPk5Nliy/x6T1V4zBXhImDk/Juk/E9Spw4Hf7HK2os
uEdpF33s33Xzn+392OgbVtv5MG+0ui3LkHAcd1qkRNob2iZIVeI6gR4Tnq9KhYo7
Ze1LH0PJkgfIiqKmrli1IZqoiiFlCxcuObxt8Dp+u/F5YxGM9oJBXXrbuqoczDMK
+4WcFnOIwCtH8Fypus87iS5RVdGosmPC1XXFohdo+0YKdlcEPhw3GcBggR780GQ9
5xCq0K6UXx6vpT7Ft72dnSnxZOGPD8/ndsKysHUY3ybth1AqB/+BNcXjmIMTgEQU
LOO9L5NMlHFQIKBRC2teHDZIrhV7aei6yxhMhrZKF61q5pO797EevGpZ8cugs+Q5
Fea1Yt0TQJDjr11x3Rl7bXBoQcU7cyJOtE/btVOaW+MFrW9dWMejWE/a0c/eQ8xp
dsCEo05GywJz3D+j/nkIYazoZpJCWckAlXs4sECo3h8NE0vPmGAHWpJuaLI8oKJx
fuJTTZSQyLYoILHlEWIpF22a6gMHHWsohqHUDowIiEDvNhe8i/h5xXEqDuiYyQ+g
Zm6rZpH6kyJAIlF2zDT/85GVZ2teXKFCyGFPFYYq5hehDfgspNsEjS0mdSZwrNf6
oWeC2tWDUN1Ps7LxYIGL3JRT5ua5onP5JzOt/h3p+V/UgwrL0zfvV96mUv6qff1J
obCyqhT/9CxhsF44nY0/odTrWMth4+EHbZ0RfXwqKOHRtMc5hSnDhb8KAyi5JBPY
L1ZvwUQduZlKNeySFYBxYIzZ86s5QUUeaWVnKktHn1iphk/3lFh/+yBhYuR4bqNb
HJ0MGV3FXMdMNrsMDvQ9wCyYCkZGM5aH0DSmnrZ1jEA+q91zM4+zRmX8Akb2zSfH
ip1bW1f9qWZLRuwuTbb8mjlHRu4byuP3V4eawEvyj2i7Makgcr8wgPCIYn5Mt2ls
ic06FycjbXfmTMrUVJ9tUTuKyBYknfJGod8K0Oa8eZYqyhlMfEy3zP00H8rCPeRA
uxuKe9fd/prJk8JoAlDjwLVHqww6HfeJZp8zb4t4Q8X40JLkAXZ1jPpnFArmTEMB
Cw/zapA0pV/zjflc+2md+OhnEjMUrl+IzGm6RXMWyUk/O2B0xRUsydptKGzzUWDl
s7Xu7ysuQyZ1gw07t5ZbZDfq/OX5t5tFEwwiPkFfxqXILoX6UKsekmj8NtOYcWOl
t2HwOmZXLOUw5CCMCshcUa+9Cx1q2QnRn9O5IVY0LgpvTSH6ty/AW7005D+5Io6k
goN/tH3sA30riZ4TjEYUzBeZrFkdvU7gKvNLPUdYiZPOq3beGXQRtRmYBK43L8ms
UD3RdW/uqhaCdAwB0MccB4FhdzgIAuI9nPji7OSOTJkKjGzUtvH2Tra4wDGvdn+e
MCVFjI8aT3FjVNzbn+yFYnxO0adAaljKxF0JjieZaJ3mZua3gbIehB9io0Abn5aM
a5/Gpw1iO+dVxeaCfjxVbpdG8LhNOrOvEYyZbUhS9xa/xK9qyS0TUzWhQqSwo3UW
m2kzldkWkNiVzLi7TMgthNdLlkmJWJ+07EVtGWxJ9R4js00pcPvp1xdoAr6R8o83
vcQ+YquVEp2uGgVct9bHTjo2IulZqXzh2CDmG7wcFUX5qGDJL6lcM77rf5/RIFPj
C7qVYdoyl8ayNtXQhGOjQBOR4L+1gehtv1eN2TkNtpT3+Fpnyrm7LaJWhjrpSUcv
ZNXFGL2PmDXSrWlk0bVnLaCUVIfpbbG7C+b/wBEvGL7AJ1nLxROrkqNnipdERvPv
sq4nYgDIwxYTu8tjJwIPAizN+y+b6oetPa/nyNnJif7iaOl6DgNjzrhlsjNQBWmR
+JfWYw+s6zrXfQxnq8CyrRizsOhXS460ozxuFUNeCNigzjd130OyZdwMhD0nCdr0
m1OrGMLcjDqpFm/RHyXrNGQWTLe9XCgrwXbeNT0oEPdFldqNtovtevZN0Zc+Nj4i
mJrpT/iFv0rUe9kWz1HUvNyBf39nSsYv4CNnS4KQZOjEFBc9qDTKfZtyXH665Kpn
mD/JQGrKPfS354vQCEqphPgUufL2QHilOdG/yYa4bWWj+L9uxeS+Olka+wp8zZel
IcfTYLYQb6JbxpB5hMka5aq9T2DgI6cCJgJVMV5yRCfuUX49v5vJMp3ZP7tEw7Wc
5r8qMn+fS+xry4XIjfuYMmZd6cWYCu9MN2cia0xTIB+MCf7qU+/26iwc2AyEacSa
godqmwgxq03hwRxE4xeYU3uGwVvn1s4utCUHdoXofSXnkCuFzNcyDCZNTUhKGDZw
sgF17wXsceOWy1+FT5BbLJsrmHvWZ0q02+tw7paA94opu7br1k01s2K963rps533
sEYhb9VlE8AY7gBcOhWcPyYrmN5L5uoFK27UtNl3LBZ3af3hZ6lY9ZlMYY/Q6BAf
BPRHS106oROLV5Vy2lggQprljPazhtFKRLR66df8NkYvGGY7aMNUtUN2OBxg1O+o
U8ZrOn3pTIRRLxTvI856ZJpXcUtQW5Ctj9qdVMiCD+y214mJZ1yxBfQTv5Z8prsS
6VSeeOqB4oplx7DD/oBDiy/zN72SRBT6U2If6G/zcYk/HoY345esPOJiXpjFvDh5
I8OlBjInz2PfPX29z1bSPUsvMz+Kce3/WdiIPBlZmeNEGdmSVMxS4rzYLEWf/lVJ
Cq2K+acXTCTLYOUAr97oxuI/JM03G3lWrjwXmUCDx9rPMwk/56wMNLdyZR37IT4y
7qitfvZaqAx+0LCE3PdnPs0zL6ExlVqLM/KvY258mpkDg3XzokCqM9/EnJHEx9+5
qkCuQ6MaKbqPVhbg3p9xal+9ihEd4OEeIAFjKfhKmWb+B+LsuVsplbRiywVb8h3G
hHkPTBtZdK46pHoYSZXKA3f0+NHCL9LfFQDJuw7uYo4TY9eL7sTIakdTxtyCCz8J
Xw3lFuzPEWOdatZi+NSZ7iHZtDkRlBkVhUKjXd0fZL6Bu6j+1es8AkD2nSsAib4U
Y6GHmpnf8iIe+b8PBzLjj0R/hNCh/1Jdlu8GGb1z4WVvrbMM4bEU7xYCEMArQr68
cFGzJz/TfFKbqoPLLxZdlZZ3qpDiibvGwhdnC1WHOPuwpsA8ZUebgg8FLAA3l487
1YOUurIpQbjq7XL4zyg8F3u+iS+0GvJ4QVeQw9AZVhJlNerFcP2wh4cblPgkhCQK
HTMbrTzjB5vDu0aC8gaJTMcHE09SsvEbkmIyCjqnqujljCNOr18lHmZJs5oi1Kzk
eSEx4XTZzPy1Zq5SnsEIwexqammZOmK4zhq4Axc2B/N49tuyTPBAGjR2eebDskFx
vuhgpydHV6WeEGv+o8VDBl0dDGm9rEXRh/OUwg1SdirYnoeUnh1dTxmhM89Jx31b
t78IWEg30KcYYcK6AOfe+IJH914wcdDL7f0En2zghJATPzeJN/VgszIrerFT7oN/
/2yjdudFY7TV6/8ou4l7HXBUHyC08D2dwpSmXrEMJGmNh2D4RGKJm9fniEh4riLR
LCknZEcTu2ttsGLhSaoL2uE3BQ/j9n0tpOkGvsbLPaOLyXCAdkodYa07YVNJr6OJ
+tPbVWH07GpDXiaBzBsRQqkOI4JT+apRbwoaGJnACBkPOGsTnnPMtdaaLKTgwtVd
V8FrRYXEwry6tHrjJywi8Oww/wj9RYaAC8ODkZAU3DEE8tcyhvtU6fQEC29t7BC8
qwZ77baSXDXXr2qcONRpShqjLuBlJjsME02hUBNy5kgmr1/iLQ/WEkqfr0Q6iSzw
CIHbxaz2gG7h925gmz9SluoPkC609+COFb/CgcunNlIzOaupm6tvsLHH6Vg1F3Zj
fZbhui4MPzP+QCZ4KjgmQn9Z+umebZgWha6gsCO/3cbl275IXNdS5BCoJS0l9ZGG
pxC08sDjLeFAstM7TKhQxtlO0FiRIwN4W50p0yZHcm5FiRBHR4/LJtQ/C4/e2rbb
YSdQ1xI0Vn+ows/b2LOkIoE5y8x658kM2b7481ueoUkCBlXsuup7aM1Yj8piwDsQ
Fk9CjWJVR4rLY+BWu0iNEuPvX6Tumgz9eX2U3cGgLuLFJtzxYVMqkooEvnN7R/rQ
gqoANJjQNQRB9ieFm0la0M8+zX0J4ej5zdhUaxPDths2yBm8h0ri9dNaQADe0NUz
jvwLgKK7ZuLDRITOW3pNqCF+8QdKpxNM66cXasSlGLCLBrNw2FtglUjABKtHo0EX
k5VVMXG0y2//eiHJovC7LP8wYOHa7Qwmli1phVEzTIJuO2Pw8WWVcYa4QrnNts9O
eQcdm9Gnsfh68YvEjPY3coOpIV+R28qlnyXckqZ8w6dxYnOfsNDGqYy6HU9U0lEZ
DVi9XCYF5TErklS806mdu5TDw3UDFmVGSSOLTeA6VMoOL/Kk10uuCoxXOfHzv2nF
9gVqhi9rbeyYGBtmimb3OiSnhSpCWNKHsOThTzKihnjisXL/zSJammfyFdbFEBQX
UJ7lgCw7iQELJh4pnpryiXLVR3eMMcBPunFrASl0gXvo/1I4lh0bbolWFelrm8Rf
H0AXVz0vPL7aJ3m0p/iA5+QC37q1unD3Q3v6IAeXQ8oryPK+8EFpd9jAXPg6nzJO
nUjX5brNGsFWfDAGLBSaKDOpLKdC5IYLDh1ZwuOCI9HkuqeL9WzfleqQoCzFf/I7
BkZVwXz+wn7FQOxnTKzyp78cnsgRo9uRtgPb09RDE1HYVjSv1vA+89MCeTjaCFxF
qSSNTqgJ9ey3OusoSr130q5nR5tRevT3jU8BUUWLfi83b7nigIZa43F4sRsCQ1O+
ORu8iInHRq8hwAG8c0Urj4xcymDmP2P6CJOEsrWdK2DV1Ul+89rLzWMxoLORyx6z
B4NJyQom1MUL4b5tj/4B7WSafsiTkxU7HyHSs/urSTEraSnwsNaxV5Mz39nWgpY2
LILHlRiefvVaxyBEo9gFXLXJz/8Q26fiGcwP5JoPbuTunWYfkm5/jariFXXvZ9dG
NUb+Bd9W09Drml90+1Ifo9mq9imF/IiXpeVNiR12vBfyib010Mnjwe4cQbBKHL04
WNwCp9D/e2WBX4Sw1XPLoRJMJvx2jSID4+zD9cKjGH51UZIhiOOMyhN/w4WntWuH
/ftZEVxhEOgl1aBvJFUzyatqOHFElIDrUwaZ6JeusO1w+yPDFpzzZSjgzNhthrbc
rM7vx9E4NJKcEHVt5Ly1tYWh9KkT7ZLsen3EmicLhoKaoW14UFSz370vK9btqTus
arm26flV15220TSr3KAfGD11BZiayJEe2uHMr5taxIs2P/kbybx3ZRjvNdH/w8X2
a92pSbPjuZwPFnuaBxK/YJuwbGf7gMg1Vm2Ve01/XLI0fjbE+AeRoAMsODVbvZYQ
JuAEe+p++A3op6OA2ocaloTusZJtqfIpWJPjTMzOZyCr5De+M2reAtU02jja0hcJ
k0fn89L8T/5X7rkE/B0qnyP19izmfGvzg1fDEE02z4PRyUMKO4vzzXs275c589YW
oSpxYfd4nvYmXdbm4P50AmRTe6k86DrKu1R9gR9DEy9c6gySvjaPU4AA0XHtVQdD
bLtC+hZjWa7xlhEJLJW4xHeuRIOMlSxN6cflKxA1Dqz1u67hDfLFiYEC5TsT2+qA
HpCd6DLUnQwsRpoXMS4xJRBWNVcW0q9i5XFPbKsVTYmxAwTYCbDrR3Jm5CG9q1Fx
HdN9lpjLdwQAI5Zo8szlQaGeQeoHKz68rLfO+hl2ZDP9A73qiVmi7nQX0kycRAOI
IaL0C5QMVC5t6Q1rgKszURuMQkdDChZPerI00rPsl82i7OVF445Sl77jK5fPYrfj
yOiktcGHrEssl91Of/lLRvOktGj9hbkha+96I8yjw0CtnXamppqLeWS4RiooBeS1
QPePOmpk5XTPRtn7IyUi87AOW9wf2JgyJbuoHBXyZlSFHktqrHAbq09lN2NzTjYx
ULqFl4XPfGPJBliJAAVGXacQyBkLxG9/DQzjLAlTsfHbX3Gu7gLuQzJRyFLB8wlV
co01v+6DAtwDceFjqeKTwnyTJ3w9o+eBvOX6qlhBb3iSP5UaBJm6aHTgnT7GqPOj
xqamODdfYhtYibY4Lo9sEqe97k1+LASVye4Pf1dBRsrwW+UQduLJrXZNoL2U/ad7
F7D2v+xYOD5svuwx7W+hn4opHEy79tedeklBQ6smrPDBE09mwAwQPn2NWRw/bLW/
0xDNbCtgkK0WH9hv2uzEYt0O/KL2T95TM5j7aTSl4hvIEweICCvTgcvWeLDd6QaL
OLZEk7eiwlYLAl2vfaWfsuwjuVpeECn88aafQj3O5VyUk+8aJzwLmCEFtLSuRKI7
P15rAae7hbHDNQ1EXT+jBmKG0ZEm02ZgvudZP+HothxiI9ldjpMgplmAh0Wg/hnY
GYZO2iyEhgN4J0D5HxVggyQB51i5RE4n3Tt6xjE22EwO6HqIGFkBVayT/lvjqoc/
4Ah+SzMAITRvD4ncb2se72csmTjn20Ir3eqgv9CBChQt6HbCh8Uo6bg9LU1C59re
jo5ZOt4oSJ04FfROBemOcVBhlvI7g3XKYSBf6vcM5uBO2drUniYA429EWq82jFs3
yrlCkmscsRE2XjGo5W8dEJzYwpD02aOPadVbdEHh7NLVAxGMsA9CJ+n20Rq6yPm2
jdbaq0KKiOAZmF5JZ8PIIE15j/PDexmCgWZ+Ql8RgBGskVvqCEhK4XmAgQOm5lV4
FJ/g5nZWL45GqfI2609tmcGIWLevksbBxLIlpV+Hu2gdbJh7U4kh4GBWyJaMID9X
kqge2tjKiTbhgVGTkDR4MF4qClN7JZg8y8KhH/VkznojJzSUSk9rzC5N+MZss0o6
9L3dVIsB3tSMvYpjJ4gDan4z2c1f36sUf5QX+nbpGq3k5uGmJhAKMyL2LWNxRvnr
iD2CG+A93zTdBwX+vzx52Kny8SLNKj1pTXeCRKO11FECiVfAfwxYt0ZiTFQxeCBy
s9IUaIBxq5EkDXsopi48Wf0mZ0oAH31On9B0yyJQ1Ue996+nIZEXTW2uSYBphysp
aCjue9RXUqRNcv/ZD88SxPtFPVC4EW9hQLbt8s/Jul42P4KpYbSsKltcn9yUQuuN
1qrAzBbqLBnNrKIMQcurRoKMiRG0OA9QtQ1wk8ytNPaiqLP69KBx7VDmvFNM4tKL
equaw3dfMOO+YAAMWBsSzpl5m+3RyPhl/QB38mY7d9yoReYz/VqrgiTSshZhiYLc
i+zjOI8OAPZIG5LBP1vV6p8J/XrdRGAYl16IEZjdWRveLnJuIq2K17ci1AWHZU31
j35XSRIk7okGNeLxOAFiKSf9v16VefUS1Jc1vw0+NlrDBICNIJO1oVRZj6Mg4FEH
Yb1hmbUJaZJUyqtENUDm8rg8WKoRAfKrWxFpcHnxCl1HMJc12BStQeXFxrUbYWIG
TBqDPIAECguoWsdFe5aYtvUI1bakd/E9u31va5CH5hM0RcGIiDw2m1PNRco9hxEo
YNEo26ffjn0rHjXMKovHgesST9uOS+eDdp58GfWVdZs8CimqyDggKB8YFchJrwaQ
1EcPLGn9NppPJiAWj8atjk93/C51BRH3mN3KEA0EY9yXPBYfr8GEseQe11lPXSqA
GAzk5ENP9Y73V9nMENOXIyHuvM56UGyd1OLFPYHOriys2mKWmN8RicDGCx0LLN0e
2SmsNPiHk29Z8tDtKz2qrWDTxzRIFkH/Xbzic6NBEgPNG2pSGnr7xd8JlQ3N/V2E
MgN/VGUd6lvxoKCkThSik5Babew1cxe3ihCTk5oQGnlBx6/qndScrqM+cbni2kDv
2hkfd1InhW//xdOoALYSdkDAJvVMLKEyvqP7oX/0o3yzku7ROsc3NVaycIatM6PV
wN1FtReVDSYTTCdptWDHX/neSxTn3T4ZZgJ8PECECxuCrgUNV1SWLDQ8eRuD1tgh
udJK0XjD3f5cVw8MpnER3NFUyrvrD/Aw4eMa0S5vThyn8WiUkn2NrINpEX3L+/FT
sIxvGmM+Aob03L++lGp5ASTN+uLwtx/u/8VZzWzNLTTPfH7hJibQpwVumX8Dxegj
w2HN6oeRk6JbGgGP3SVpz7I5Aj9dkKwQ0NvIiyWT5yS5qTsOnm7Kd3vVe9Ui+Dv1
li3UwxgY6/uv8O2TTc4EsmOcRq9WfKH0uIhyjm2I6rRxbqrPni1vbn+uWzrNKKZV
URwrieC8wzk3JjmZICSFZCmvYq+ZmxQUIW0PVzFd+K2l2qwG9deACvlKGCYhssaq
z/eZ1Yn3AkQVXvyfBV+l1MBYtLMUEe62oG0UuIVPwBuUZML5Dhc//L7PB0sfIy0r
1PXk4K6X/o6JQXvE5KaP6N+8bkkIoYJ5oABJxJJkfR2JRubQCoKczLfUnLkokfAj
MHWHVI0s5OyMkmYpt3nprS3ycdILW2MNZf3D7PySjuBHqaxQHtWDurrmnFyWwIjM
rfvPczSzeJ2fzskuhaF+uB0zHGM7LAc1o73go/pTm4h2hTLINJiiuckcJZHnsgwn
dG7xBrlrW0BbJ3AL2RufzqsGiJKxAmc9V6h626v3jypBNCp1IyaE3Tx0pLr2c6CZ
GKUPxcjKHLfY4J43blTB1pBUv3SH+rxP50UqRP2sl0M4llKPWSdGwRNIFMq9A8U/
TDeqKB5WxJzjgNtYaICBu6VelIYr6a/03VDoDNAGapUAJLbQfnSR+Fmo/A6NOYQJ
RuVUgbhZu6fsjxxLsm4IGymamxgWKavRndeB5ePns6wtpBHDPLB4aQ+hn3NIaasu
46jvMdt/ODWmyCnmlGSsriV1mC0V6y2FCbKlI6pY3rEboHTCzmnXUaiHdxRhY5fe
LfcqF49GL/G8YkooZ8SlKgXXW7MpAE8owkDiO23gUrTc9htFoiXVhg7IZbo41ipI
aVfRq+R5PtsZB08Y1LMKIGBzVMN7uSUrfNmJhW3vLaQ428E6uJqWwXJfdxtLArHm
WRC8RsGcEi2J4nqZGMMTH/ceBKeJ/dLj5JRT1Kt3BXUyX2SANErPQVUt5Yyo70Vu
S9XxARboO8NiGfIDVV0x9WwnOzxe07/xfcEVnsqP59AuX1UoNotKePAoqE2gS4bx
MuLqF7C8aEOJ2VqR2uQU3JWDtWambb3VNprUNX/JDLEBH4iIj/7k8B15fhfMxB+7
IeiNd5DyZfz0NvYw1uu0SjQsbsMYXCwsD9rSlynFg53qnPNZKgSMdG7LKejo4zs7
YWMyppgYe/BTfLse0HyOzEkOmYleLsZpJJN+XqtNlwQWTTB1FouukdEN2sxfC7KD
yto+3rIKBAnHwBBtLYE2HFNALWFWTN6qDLJp99Y00/CHqGCeEgd0JhUCTelbKLeP
nNNpjSm110F8PDZNRb+G4LKDnW4VjWTbOKAYUaXkpbmjN+nKAyxUGZhtq2NfAHqx
DhotBDuPpEg1/Zo0HSWB903i4Vt0UUReFibWDg7Q76tSYW0wavFlmQ4flKEzpEOv
d1f+zvf4yG2G8fz/OAN0vNcTAM1wWjsDwgdpZ9NYviy2GreB/fsrn8NzNwh56MCJ
Sgoj1fiyFVIy81VweLy/CV+xlnB6zKYeJm5uhs/qbeIaXUmr7jymrxf5D9IAdnHK
Iz//uN0pGosAke4ch46LAPchUfhNYnvFDfwCKLloekOW95l9WuodwQISYgTxE0Pp
8MF2gtP9qtuALZnpmXjpuJsFfFsL0973C69E8RYJq1lhyVn7tgyshNU6HWJIVB4G
wJv2D+gD5lKa/zla/tliBe9Er3cF97WOgfC0bELTvfpUWd1Tx9zUcMVIPfrUHr9E
67Lc/+ulctRVKqMJ1JsZozgdd53HXYx2MwvRj7whLg9Qns7WGPko7sO362hpGJIS
yMEY6dRw2U8czd11GIPyvyCYrDjTmXdHF5elyo1ix6/qHzX/qYn3ZiIKNR5X/rqy
81qyTUHKSKZgNEir/8yzANsCAr/jDyNCL5YNOe79AN4QhlbN2Slc5Aa3ldOAMbvP
0GRbATyzNbNoSNxXlYj09gYb0TpRrw5QWiPRguu9vafE5OUGiTk+0hIJiOwoC/Tl
RXo4S0eZKZ+M42e3FW4JGc4uKmv7UllwTErX9T0LGogI7l0UYuNebsuCcxRTpKyV
FcAzJZL9bJl8FUrVFxM02jful4rbTkxEW3A+S88uLG+hVMj2RbQyVJMYfLmUFK05
QoRbGV5ZZE+OjWjnvw9XWhP8/EB9yMToXWQj7sDuevt1MgYubur2c4G2rU3oPgWY
o7GfUAmGLx9qck9KKtA1dNvqrDFs7qGYb6QTmcZEJvWHIWucz/6nnjKLyZ6O19I2
6w4fsHzehDW1vttPZlpx5lOfS9Cq9LwdVX7lkxyJKNzLFkDRV1NYvrKlwYq1Oihy
07TsMcR7RTr4kWIInlpiPswsawlQDvGopV5AykIKCpOR00Mpz8lFtCfXb4/D29Pp
M372EcoMyWzU/p4/XSBDJpQs3DLbeauDnkgGUXobYhlS53QuipKjzlybI6SJVhO3
KEOJfSDU+Ghlp1f7pUEmvwY8OSh+JOdyTmKnNb1gxNLTvcmK41SxuK902F4bnamY
ocGv2eNEDl+JVxorsvV1CdXdtd53kOMwYDRlED/Coz9j9b8QPB+zFrA8+MQaBdVY
cyzZcVgGA05MUpOKi8vkZyjweEoGwRqdGJzRWOglYDz6r3BrWM5SbDoewYt5N8Yg
bQwlKabBGpo863xagQv9g6G00EESijpls6VHkgKsdJtH8K3aW0zCkD3FL4SiZWZu
O7Lnr6MYl5g2J1X+O+40uany9y4gVlxCRlPHqx9C1yDtXEo+Xe+XDNtAj1bdrm6b
HelE078O5dy0/UCuiMJDggXFriNXDQUMcGt7SL8xNBVKnR2zx5wlPkUM6Dj1DeQB
gEswnwTuK39XfjZFgi7iJzbkCXho2XkwcKrk9PXP93SNAe/FriYCc1nowi9hwyZa
kmllIAjYDIHjU7vlV7vNgHeRZpgq7nahnNi+Fcjk4XCRE4zWAlIQU1+Q5mSFoofB
QswJF/Os8QZCK4toCytDjMmWdd/BQXRsQMs7s+bZAMgLqvQKHQaHXA9uxkpLur9E
I89OqmCfMzvUJGPbf/lskfXKNCLwEemngt2mdMli/UvG7FRj0MwHkgHZDcL8Jk8x
nRQpoaj7Lyd+30RgpwSnK579BN9LPFHH2kZ3Na3i179neUiD79W53rOR3QeVVprr
NpnSslIwlbqdYu0farFP7C7yGPQSiJRAEa3RPAS6uYmJGDb04F3BV0gFbHqMJRwK
zbsPq+rFc256jEtRl4QLUf5/0tOPcS4g9vheXDV6rKGP66fF+tb99pQSQVMklUhB
ThdEJafomva0voqLhZNH+ySzC2OaDk0LuI3D6itZJb/hZKSYoIreGTW1IISyMy57
1EOn/f7dD5jYgGaGIepKHMFEcSUdtFWd+6MHSBhhCZZcE4SqwyWTccH6K8aHhBTS
I7WC6ThNnQlUD3Y38NAsUKf8y15/K3nPPTyZvrrgNq3lt/eJ75mpQNlPftiKHPhc
SZ6OoEAVNA+2Bva2fWN1Wj2btyJStOaYRSaCOICIG8lJ3dxsYQ7wYjXHYAAy3im9
oQPHJJ7pHXgcfSYgSMrkFwGVsO423hbhSAckhUV/yezEfyY77JwjPeJZ5/ht8XIw
xwJ7iasB/HLDOZcG+EdVbr2eE3LpC8D8G61TYp5YEerUxeICnZBtzYH4j5WgEuNG
Zv/uHomtXR5sa7J4qN6rQKLEDldrLTcZVE6hZvZm7oL3+zvdWnUsfjOH7dBMBJBH
8j/qn6vCoIE9ppYwUJMaDC93MsSvoTM+VvHCSBO/lhj48BKHgKK7Ajloiu7HtLMB
/0DuXi5Ln5I07PwA5ZMCdr9L99HGaEGO8NbjRzAZDpoe6b7WZGPiT9r3dWxJOPhs
vNG9KrG/RSbhlY24BaelzuiZzfAAWS2y3N9J4YwO3Z7Cko110A5IvAHO9j95k2eb
BiLdLHBtnfZPFv7Pe1w9J+BgZYDXl9zFCHD8EuObe4kmWxa606hSBX761fA3PF5j
Yzevo2GJrgavjTrDoo+SkHecOeM6I5CFx4WHWhfF5xqFVNEVnrut9Zd6a9HZpYF+
KnWYeyh2ft7mCrj9I6DXT8J27RQFe7ifd82iTMWCldVwCiRwptDFyoyfNURbKaW8
ddDTVjFkKEeBOvdRCneu3WsezUa8BEBo3pXjL//JN3FAWIMUrazwx3hQcow4r/ID
UOOqVRVqSty/AlcjhUmX4EFmAZqhr9GeNgGt3Lqw94oWBvK2242piJyVnsPAdiZR
7fy2azbOF+2Wt3Lbp0+r73sOVmzMq5Xg4BIJEy67ba8MJmvsgVbhTVVTXyz6v3NS
zznw37tOFwZV/bhrrLwxt/BJYVe2RgMQuQN76czDnfKCaNPZOjL2j2Rvi/Y5iXRb
nbDoiVJh8YFZBg7LM/5//suSY7PobtaceFkFxqqjTPbv22Av46eJBCyxLXsOgJWn
H63kNgCDv4SZK8oaLYt1Pu49TKDdpmKYHLLOJi3WjA4cQ84aM1LBLfoODlJKbni6
/xVulpz6U1oUu8S+5IgApnVHCE4aB1mTyyn+elxl22gzmJYmxmT1G7P0qsvmqN40
yuKJ7blybljRWWGVCV2LyNN4l+FfiM58e9tQ1JO/rXFmjFiMF+CksMatFn6W3VXh
Jt/ULhEv/minn5eP46MbdXoAeEC3QjI7R9kVqfPLXoiJxWZbM4Xlbkj8I0KSSEEO
XXSPOPgGF0KKfLfa7BnXEPLMld2aw57/3GSn2olY2GupW4YuxSI2DSdJMDvFNO0y
M1PzN3xe+onVjyPd5gQoRWi7Jiugk25aNMsJfwyt+P4+zqHoeGHfe57geLCgfUzz
/JSZ718akHj5heA3l3taFkmjGLNJYfF2S/Kda13BPQj2KyowH6zH/y1dLpP3IIDo
FGkkjIYJ0lwrzpuDqk2sbKkID12gc8JveJh2z1MjfWy+Lcd+tNVqhLLIggJOEIDS
6Hja0uqaXzHk8mUBIqHaUPqdCaYp2c14vIxt1M4MkvBAuSbDfBQb4C25l8Wp9sQ0
SYrg6t/tt9PuNlnzGkXSDIgQcXUTbCP3vkhHU1MGVUobM3V3gzt0pc1HflgQXgNl
sJpus97Gm9BSzrkoiP014nnikHn3UvESf6MD/j/VOXQ+m5krA/jX4QGcC/f8VrVR
bYtmkhQL4vpWThx9io4gC1OTw3iU/f9NQIn7mvdw2lv1jCTOPr7+eV9H7jwGeH4H
/Q1vss0Gz5t8vW4n0HWC/ULqxUURvAdIwxa8dH0XPEFrswPrjSA2V42kkjuWoexr
SrbL146oHY9I62uNDgl69oZ3Ypcgb4d25JXMeO30qMexLO1GsTp4b2v3KJvf02Ln
gqZ2AlOX0UEbjgMOUf3iSmiR3juWGe6lFU02LMV8yQfkW0ETajEwwhjAkjimaZlL
VpsHKrQ9AELlBTSrYT7CFRiCrdJsndVjl+HOBA5VGgMsoQAduUQrhtv0Gn7pb2M6
DyQOv0t6TTBE2K8sWvp9BwVgwta7yN/zrENM8r3vZ4UeYdfZsgefjYbtJY78uC+x
RkU03bQ2bvlPUZaK+xUHpG0Po7OdZhKWIV5DtNn6GIs4R6WP3CNjXFZDvMonRI8X
33vpVp9Z5wdz/R3U+8W63BUL6Mf6gay8dSsDicM5reP0ZSuIbFoyb417XjqcTppj
NJ/tT4SODaDdNIPpvzPVWBBoabv9oTxdVxo/AtjF/mJWKdrD24bWSwQ1vaoO6i2A
8hAFZtT68lxGZvbTkIRmAOiipZY/Kx+pWRX7bIDQoYCMe8V/sAYhZW0iNLq8Rofj
x0dBhgugeadQIhG0HmzVgNeUcqxV/roPGbWW5BcBxFUxnNxFnZcs/pfNj5t0mVA5
a3Ugx4ZSQ99vUSZeAM/iXIJvMI5NhOYtfs2Y28TdCMlvpscXk1ljUs6jVmRYv3Nw
TJzW+lmTzSkTAki6xNKnY5dMGFQkhncFYMluYPZNnRgdPQwZV0xmEEXmhS6P028H
R9xrNhl/WzXoZZNfePovqJ4FrERvUJiHktHuxZuq902TGhQ7PAX04EnlQHTQ0ZoO
Us4G312TDf3zFPItBsssS4mXpUO6KbqqUQWMr+CDU9cQO9ujb2+HMT8xfQ9G0Ojz
RKJqKIzvt3skiXPlt272hZ0deibj6tAEvDvXizvBA/8UTlZuS+2P1oY8DksPxNK6
5We50Z5VKXGFRkl6/MprBnh8e6/M4hrb5Q9M6wvRph4ijPqGYTy+eCjuwKd7D0qS
gLXeK4uGOobbh4pSZfaklEd3S7vncsEFhbopEa4a5KiWOHk7bJNmoz15fLzrFcbE
QU3DSc+7qQCL7K2URIU/8NwiZ5Wu+tOzcRA1/Yc0H+pmGplmmbfPv0S/SB/4yyMF
aljTmJsn2GVoxWjJVJ6G0GJ+uNu5EspYqtktCYlACPGMgT+NnC/M9qtPPkyOhOyu
kO+1qxqK5B1oD162uRVTsVWOPa1x0KBpiqI4oGOFmnvxnfpX43AhbQ77GYWfFGQs
AxIfaly8CdXALyd3TNdjOlYWZBVsb93MvF0sEQPbXfmjXhmCR3GjFvVRduulAnTb
h0EXOPxjykmzkktAQ70EH3NxlKZ7YRoyFqJd+z9P1SiwZvF4YW8iTZes+pt/w/o/
zI15cEI1qFUsFEw+tw8hsRzBGh2vBA7qQApxjLWjf79QcfWrAEQ9rvlzCTRCC/6x
nEZcmSYDjc7rXAOZCIBm6ODGP/KEJuu2ZxsewpKH8F/DB7wYMQiGssDPW/V2sMtl
jRbgCYN+9caoK4HDykm8TYcwKKi57yKvLzvzeh+WJ2duv1mkFGlWkNO1ZZzGxuD/
UDFdKLf8d5FFws0DoTx0Xc/iO4XdU3HFOEnIJCct1rUJ7je4S/loQ2VXh73vHzV8
X8trUcgWccI2y/41kbtUmopzcZJ32MjzcKVayDow8Ap8LlyroBAfFjAvqf/n8rCi
dKsLZA7cJSYrpsRGDofPeFJO9aWjY/yas77gYVh+6thH9Obv81+QKXuLGxd/9puR
iOxEwF8mHF/x4SxzXa7Z/IT5BnhqN999OyWs1VtKMuLo5cRljeQ6wDLMMwhsYq2r
YH4QST23Xz5VlsnkuZOkocTw4JmrrPk4mjp5LAX/EhXOF5JcTxErNae0+vCnhCJl
cMKTq79X5qHZvKhjyzfqBtTA26TRN8x0Gvr5r+eX3FMx6A0qalM4vutKOZpzjCHv
ht9saLC1kTclS4RGpJLKzFZg5usqMJu0iOuLS0gie/xHNMq9KweS6izOJ0A4+k4w
w4CrPpwbKFZ/v7uKS7OIkDz6T84yPbFAFM/3uR+VHafFlTzW7FilE7yF/Z4Tbgea
GZ1DyRZYilFIQZ6ptpZWr2c66iIDLmJcCS4s1tSFZLHGMvhLSSPP+q6HndWNkU49
OfP731OzyDdbVBw7SjmPZJad4UT06FVwEK8U2yX9qirfvYlSUslKLxOaHo3rHmug
sQNwFE7TQ5GPrklUkvIYRQdw5sHeGFKoli32W5oI12u/3DuBKTcSuVcOFpkE4+Ui
CRy+3x15yJooFKyHt0D8tgdJTvSqTWWja1xoBtOgOYA7Dr5Eq3c7Ow95OrlLhHYq
cypVCiYkWXsy3iovKemXKsqkB3+wHVGQ12ip7tBgMN9ncPGyBHgZHkokCNgJrxIH
wXDG+QtmzFjS3Vo2G5WGElV6CYtKcG1EkgWJffcP9YpunNM0wViNsuVYHURI/23B
W1lZbbch+60JTIewqAJJqZ4VVLqxhdoB6XXFrZhpXU7frhSpeAoUrSv9rbwQAXTl
rYNCoyAsI60ElyfjRuKXCdrLTby1Ib+52dBkObqi2tygQBTABLA3ecZytg0Hhfp/
ciIKXN2/kbAL68T2YREWO+eB1FkFDUMNYe/uNohI7KhrBuHzALs9MLo5LbFX58+E
GSaUXWFCqkm7855l93JmZVQ84fR4RK/WbtRZHy+hx7hWk6ajvwX84BTWxIUvE4CS
hXP2YIlV3Mwm20ltmxUi2MDUYxem0on9fb7KjvcpxR0hbK5Jov/7Mot+myF4Ayuo
WY/fDXPFf9st3vCokq1uG0gm6dFnjZXMgOcLABndjkkjUo1Zbg4mCWBA6EQrke8K
8gHjjoYsH5unY6foMugL08E9FBYdpaM8jA9TayhkMdV5ISOL0X8ehRQaSsEdPoG7
MDK9qERK1D1YMABV8T2ps7xHSGksLOzMNnePsH0kJq2ZrYxcxiLu7iW2CeFsndb1
y93IpfaYpF7SPNzncPA8MmAuHh01qB6VUJNG8R8MDJsh0+OiMV3bdyMEoWd2BSkI
U4ptVGIXsdUuj7wC0mzYqRr9iyF8g3Op5IQ/qPWTZvabtWZ6OBzxS6tNabXjpqFh
CqHPw4Lp24ysYqyTm8icHafmhgoqbr8hv5m+3w0PpR4jSsi+pRCytJP150OMb41J
qnoWUXtOILOwpigkSShFSih5sgGxgAv+YFSCe7QZzDay6NBacAYt0v/VIZ9LJfbG
+AANR51FPG6unO9DXauOMGHqLQsI3YdrP6DAHgy5n8UUW8mwzsoGcB1jObJbgHwZ
NwCgiRYsf4lGB3rd6mcPTy24WaaH2FzG3bg8o8SSX/8=
`protect END_PROTECTED
