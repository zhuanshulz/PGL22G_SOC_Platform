`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yluGkZD1GG6UmgyHE8/f8TrxnbJuy3Y802l7+7XccosI+H3tKdRFUjlFtmEVI2wh
7MLiPV5ZscENeGXOuZBDrWILOBEgil6S4WzYIayze0m+Vv45L30PCxVAzoUQaIi0
3AtRAmEgxgwnF20bEWq5HJ78MqszqyHXnHGCn7LR5rEQTkwFpiWR60lUYZjMpqpe
ym+2vllRpeGU6YhXQQQzAmUsDCk6J6QocQFEDRaX7yWSoCvhkdwtYckyVT71eO4c
S92dRomfdtaHf+GWz3ONq+1+mCOV494zI8WKL09MY8CTUESq5zOqU37q8JgtYfbY
2mbpqWTVWyJAMkSGMMC8BfYSqqgqZcvU8uUgazrt7UGNH0saCBxPDHj7mj0vkXeE
LyKvWlOCn5yFayvmYY60hj5NTrdKuJ9Uk2j8Uqv8bPFXZN1wbSrN6o+UqRuJOVYj
AwZauor1fExUEONUgFI2Xtv4iE0/efkwGQCZ5cZrC0Cy3MRo4B8z3kh/1TY5PJy5
+487mYl2i8VpuaOiOJebByKhYA5a40xSRpushvSKXBqMpxGLQag98KScG6Som8N6
H2n9eYxwEaWPRvyTwBcyE6IH+GrBQQlK++wWaVJTCoPQg7VO4LM8RdukpC9pFyET
`protect END_PROTECTED
