`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
scBzVY2ZwqsDTpJNcksCyLfWmfT6aK7OX2x4cHMYPP4qy7+J/cUBlOpukKGLrL1U
zkkPGLn4o0scPG8mkaatXVHFepvn21GiDyIcpAZhak21PNPeja2csEmw52L7VTpY
nkzlnVjxEqhG81zpxYoGB+wVySgkOZBX+65OQHNL5nBXzEJgmQ+lK+7ikPMdJNLa
CJHOg9rfusD2rDgtUok3t28Apwfad5N53411rsJGUmgZ//m8EM9l4QZXk61D0KB2
0DME8SItp1aauWa8sfBc+UKgXWaHWm07BAHAfn09huTUaoChiihF6Yt4oU/ACerL
Bt9aiF6q9Me3qrnNWYIPjVciRjpnAuBtZxe81jNIknmBt17oc2mS4agH+lFYQ/O/
B/EYFJHvItlj0J/ZYF9AN1bRhg0p/AB+OzNaPAdI0xP8GBrPXeGkWk2g8BRkpYHt
`protect END_PROTECTED
