`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wmk31piwrGLQ86ZJemnpCT2KB0vK9CSXLHzEMztD64deS07XIw1PxeDgQks257yG
Ma2GSry8l93+5LGBwtr/OOR3tjUQdjjtjFAjcPQt9MghZSBVMK3jVVv0BG/tDGq+
kBs2QxCxOZXCIdEIEFilIxScC+QACxNMDTPWb6hR6k4XfEylceoXqxsXJvv3n4RJ
V+BFpLSryZH4BmJUUlQ9lKH/WYavWikNSqrwCwf4k15xTO4QATsMS1xJ78J2SZ4T
0tMQbGhacvVRmZHuyKOfXiuiaGuc5Xp1hcDSF/f7vLEE8SPlPo8KRIR2vwmors7F
NAJB75zJ98uPVO3CNvgpoRYDTnxOT2YAtuiAaG1x17cuUlaPRIYe3k9XvwZVE4+x
Bx/BklVjoVGB7kTdlty5+ZECIR+x08mEYR+AtpC2HBhqDYyjqOrrkF/ySybu8Bx4
bF0Y4s7F28nq6ZxAHpddEPCyVqmPKj5opureihdDek4onsL7/aMaNq/cyK1xc6Y9
wh5PfB+Oh8NtX6jNq7Q/p9QlgUdazFZJ4jrtxLRxuc1BuBPW0NnAN6eNXJMFxMPN
HaTG2hJohwF20UUbM8JOGNTiRDuLOrH0VJ+GZnO0PCqds4GVLzDCQRc3BKryFoHc
8vN/Ct4cQVPe0/1asiqvUy3G+3S9y7ftWAGt8BdGJfo=
`protect END_PROTECTED
