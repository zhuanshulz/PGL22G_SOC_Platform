`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H2V7BI2VIlt7t7DwZqIIXT3bGmSzDwjHb1ApxYjYo1s3qEI4bERJIv9KWhw8G9Vc
/8W0rnF9TjlH3POKb0TfQjLz8rM+DH4vTyRBcrWBOlwR2s34iC9uk/Lk6CzPpQNX
0iGaNgOvmhSQmzrv/cGP9HbHK+xPKPK5invqBZ0rNxK97D027elp7hCXUjzDXWm2
s4u0oOHG6+0yZgfBp1xsLwDHBkxdXTl4pzFbeWYSf/AohjDlJA3uxZk85QjqBFL+
1hNXi1xVC/HLQW2CdQ8uNE07bFtKT3UTXEDRPvCO+Lk56bCu41Br96voXdYTkkDG
0Cq5XEO+1+TLEZVKS74gjT7yqbXZb/IF9NHl5F4hhXICodIrXGHTWzZNLZz30tBX
Mgu1vs33ocHl2SyWBHZJSHR8cy2WRjCWLO/ubRRfleBw/cTiTP45ukEM7dLnWCbt
TVKz4r908NmKHmT9PhmYf1FbCLEvi8Y6BA398WTd9D0IzCy/n+G7n6bf0Gdy72uu
9Efw1gB0mbeDKcL1sBnC+Tr8llCeX0g2YT25uFuNo9Mhl/RBlKbw1CGFaRaBST1p
5ydAhsxqfl+NpyYqUOje9JyzJmT9qXoVSDA+5nv1cFTqNnsKyW1qZP8xZHevNwfW
/NX/YqzWCtC8jPgOE1puevTa3ohmzsSlk6ERJBjTcMqHA/NHR4Lr/Z7N753a94QG
OR5lWBGKxkg4chD4rlkE2a3dZu+mtEicBxs6Q8mHkv4NGz8XOUPDlwHXytaVEGxy
Qy7mmkmXnQSf4MSoOd4779lwqLWMIEzYShoXvsAU2H12hRHtm2Cyt9kkKMBbPhJY
XB2FKw1KBd7ZwOUr/OKjribMjO3rDi9J4JZhYjrJb4fWQMSR2OaIM9tBBMxZrzQ4
ZFdHWIEMymQLPaDLMCWbtJhfHR2Tvh50JqaKEd0aCOEJBJTUoVB4RmlgnwWQX2TC
0bxC3Tza4tCOCP8YQbErxCYE/ZGrfrBS6vrElzbsVsa+CezuU8x5uk95diRyoTN6
CmBmnUv7kSl2LhkaHPQNJXomRax7hKXgn+GTn82JzFBQIkDilT89Jnbr7SBtyuYp
9HieTcpYu5gxKsSIrm61Vqsv46aQdaYIQITOfXeCG2WpAWgsWnkLfvfU/sO8CveF
XK+i6QRTrtxF1xtEqWmTopE205AGjQSb+hosV/oCJ+qrVkwxWUaWjrvZwUjGslzN
dC0NGAVgr3knOOIY9yIBvVgHoQOuiNrNaxlfuo9keijXArp5J2CuZrYlpPcXfs23
oCR3B2ZCChr3MA6ukfGL/GECUFZUdFjRc9OqeX830DBXsqhT8KJ99/J89Qpz653V
xlgI4UccDKBMtWWcGld9AtZgPq/3BXcHnfl8DkCoMytkDIFwJtFuUUuL1weDMm04
YQPKU3SWs6/jej5xAFBGkA==
`protect END_PROTECTED
