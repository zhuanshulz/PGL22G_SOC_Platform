`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DuXXUZuJWfyMdtlVYQhz82xR/XyoM9xPlU9PZwdY9sOvjkqY1hTZZsjSJ1Js5Uen
81boa8wTnurno7QhP+gJFebXqE5eqjKSWUtEWGIbilak4M2BryYgCSFLT82LwVPc
0bbx3PvrFFOo23V7KdgjU0ho5NbFcR6LNdLDgTDBB6GfSxmT83KO+wZ7oP5UyXB+
rti9688zeQf1akvn1GfdJ+7mf7uUIqwQYHdC/FigGa5Tpqmnhwo0m6J5eBmYraw4
tpHxQaL9dQHCYt4QoJwy7Y/DgJJCT09jhAixXTWckd7ApWKiqdEQNTqQUx96JLGi
T4V/bJPA/nqLrCZrX4nplav2ARGc6Se+L3PEHJ0WLAUlIE1LXINL7yvzdx2GLt4b
G/0RWqog9+T5dKpQrbPyHqpADZ13oANesJbo++c75rIvLwCSvW/imG0wk/UoaSWJ
/4MwO/3xeyoRmMmh9jmDF/EB+ysHAgIbQd07nh5Z/tnO2YpUCMeW+FovbNU9EX4Y
uoJ7uZrjSih+h40RIht/vpklFa25JpIiZ1XwHaIaATMzLbMntloz/NCl+RFKkjA4
lk3RVJDUN9IiGh+zVE3aVHl9YGuX3Sp+LSV087qG07gD+h/FgrvEJPhi6PPKhMwJ
ke7z5rwt7HlWaT8U/ON6jsYPIuoOZXZtG/0BrXKQQwpjJUyFHgg3RKVd3m2cFD1l
5X3Bz8jZeMsOxtyM7/WLWRQd8NjySPOEtGISlFgg3gR7l6thqD7IJ/XWrN1QMCmN
bzj/b7LDgJ/1rA2PMtsCyInQa4G5t//ixbFuxScTpuePq8ITh8bK9EJ0DoHABcbT
TF7npdTYCsFM5ctJgFREzlJFYEHEcIoKU/Afc8zGw9YbfBlCsDWeAFuhG8hKzaaw
jr1vM40cXmfcViwJsf29q9zk0WF4PcbCsNF5xR7fR3rSmZHm135RuP83jh5dfuUo
nvGRWeNWo5kBe/dlk+LgVTg7u4HN2mwlyJgwAjTMbKv0WLftd8622SMtRgUeLv2c
JLiSJv7Sp/IChAoUiId/mIj58yJ9/I3iPtYbF/m7VbKtzUM9qory1o3wZM/JfRHh
Nn43TK1sVLzcM2TQ+c/2nis1GWGKACPuN7fb6aDwhm2er3HnsXjM5xIyBPpOQXGL
ZcuVfLCRaLQxAXBGmPIpL5umbKFTh2sP4BKqgLbKjCn8Yeks9E2EM/El2SAJvRWV
EpOcjFPcHlBfPCYe2vK/kwVEoucybqNtDEy421t2MI1vjZ//FraHKunROtE6t0D/
0fF1/ZAMy+RKpk8CHpZ5/PxEa+0Tamj/K/juF+E6tz+rbkLpiXjhqi+ycYRJyS7x
NRTUSzUz4j45Vlco5en5eg==
`protect END_PROTECTED
