`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0uY+IZgQUYnVK5K9iy1ULRWdB4EIGATBfjwn9RXYJMal/7+q+4ZFsWQwkkbALHLZ
e54K6FE9FBEs86aHH1p0elyhxZCzCpNnXtyiH6ya5LDyLZ9P1W2cjTEdYnOj78Qm
mM1Mm0X2NGZ9bqJrrGJFmjusHUCk1MeGCqHrj72nI7hdna026CEdsTILsCc//2eB
w9BVWPFJ3Jgu9DRL18lhxBkzQJlLD1jw/mBuIXGjNzw2LEAYEwvZnzaXA8JVoRwv
pxlBVpOysVBkDV01ZGmU9wWYcO+x+dbUaJdB1og1CP+JT798iKFpN2R9m7lUgPUN
5Y/c1xp7rEbF5Vw/vyYiVoIXDCERyWSRxZTKict+yUEeVL9/p5mSeF7/Z4RM6NRb
REtKJ/sMmfUpXpI5/t2uxBqc0eeaNZw3ixafyo9MmdtpvgPXozxi0s3zs21MHhAF
ZNDWKCUXa/Wish4D3K+6mYKCben9e8JF1/+WwMK+sZjIuEDSJfOsnojDX5EEDC5E
PHLxZhtg6VY3s7z8iO8W0AD4bf+KKCDOek0hw7wvW0t1UKNxs38eSzd12NVy/i4+
Di91uiRVHHAtLi+v8HaFtnqvPi4RxlQSjbjaYqOjoeli5urnU32FLvJGLvLwQHUp
5jumomn0rZe30xFZqqCc5WPexPuwRKteH1xj5Mv55XB3uV9u180chMBncrEJWLhO
sUZgfrUimSLe5u/7lVa/yrH0drBTmm12S5+y39yOeowcue4NjUkg67AdmRapWx6H
uJ//rKOlAakiCoGlM7TlyynmUkLhBF/fmrJJa0I2Uzbvl/t6/4hgQ81RDPjcUsCB
sWHkMNRYYiLapsDCywnH1al14fhpmCDvBnxKh7RY/GlDw0NwW3kV6ABM7T5ia/ai
NwOgxTpQaKtUE6kpnklej26D7R/K3Oq1Bn4QSCZHBpaOZp1jdxueJLVOojf12RgA
Jsv71SAO7V+zL3ZxRrDDdAPDhVAD3SvhcXtEvUxeUdBQsZC4vfn2DLgqPXtfO9Ua
KlcpmskM3sg2xTBAKt5TpK6Fl6ZdfozAqVNbNB9aZrbSLTzKaV/lvGVgnGs5Z65a
w8JDu5j0AsT0ASPW7BVHWXud35tGL8N2P6cb4VhEym5DY/MxbknVscXSFBXIv/ua
yMF5O33AM/8FVZIxhVCU9P0a+T5qpm2cX9XcMjGmlONxsTwE7H+Gx0VsG/5q3y+6
98D+7UyaDzYo85B8ylt1wUqaLiaOGM5zr0SQRYKnU5PNPKLqpgachtoxDJqQ1jH0
mBnNZPM6iRlqzrOOuStKFZFxytTfnvaToMgn6bCq2ZGzaFlndRteHOnaDfDdMEsD
tTQgP2IPUM2dQOwWlOPmS/Xyly/NBrv/Sjij7wM55GD2abSAz1plTDcnFLtudYE4
KkVULd9+bQsHYLLOGS31MYVcU8xsJb5UfUWBdyu9cqk7BYLCplfRallsJlVTAAC0
D49z+poJXgSchKPjxemFuhLXOxkNs3IQX0Few8uorXYBz99kxHlF2x9KD0rcdfcY
bLh0k1shq77f4BAzv7LoiNrSR16FNzYmQf2p+qi6w2oNV73BmAcwkcgqyy9O2Lub
K3j43+rpmKot5XwV5JlbaDoxF7SozBMUdzi/mcXPLwdPW2F56SlqSyMdb3Uj+Zbe
enRvcpJ9zwmxCJZLI5abhsbYYw3V7qDpxuHSQzJbKz6i5TR9nwF4ndNrfdBRe1Lh
msja6pUzNeXxCM/blAFFeQ6FKjyaodqO5cbo38B9M0YygwCMm7il7Xl+G1Hj+ihu
TfrgY1Q/45Ps2Ntnlg6HSMyzQftIwAcZyp/Ne3Rud2QFbH/OVzRZ0oqQ8qdvb8RN
ZuinRo3mE+q1Ti5bXr4kNoNzNjgvckV5rceO20bd6kA=
`protect END_PROTECTED
