`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mfTZwQFQsPpkrp6URPxs2utHqvrDkT0t9M3fJAI5z9xEmNZAkagvMQzo/30tLC/I
/dYHq765D0c79N4U4xVgztmDmeL/hv5mr3nd58Zp3JQ/bpVakTnIIZIY15EaJhDS
XeNKQ4HiQM/bOtRip5AhG6sAcoqSYtjARUEJpYBoxOeAel25cb112k0yWlxqkyw9
YxPutHylex8zvmO8zlJGM3gY8zd0E39RC/tBaS0WtjwtMbFUR1mdGItpxYRsJ/i6
lcV+e9CgS0bLzfcvLyugjCqJXHFkaqJjNeLwOVIu2/skwyAadR+akniSSwdTNr0C
tGm43KG9lEQHQYk+ShT9XCfShAdoPrpauxY/t7xPOledTPZ/HzXYH4flSFy7NeID
1Ijj5k78VJGVBbtnWXWjSZ/CvrrHnIr6hjYwueno2v+ffQCPr15zR2kEjVsjf9qA
LR/d8lTa3DVlqGz5JCp0PkCopbbxHMAZYYMNy6qa2TjaEZGtNXUSfxiqGSGi5F14
htvra2T66JdpOW1qOztk/h8pFyubrjrfWXHQ9ejXfZ0jyor7mSOXanqPxoZu4SPc
Jh5LZilkYPqlGIv8lBNpAMQrztKJBA8/0VenCoohKrEHohBZDRoBBtMkC8dM61jP
LtSJW3g/EemBMYtXIgoeU3l2mf+s0FknMXmWRrkHqhLpTCuoNrfDinnGvITcxKRh
3Rey0BD0GLeKmhRk1PFFe3/03JhaWWMeKpWpbTww6NikbBT+/ngroqCgbP9FUCvI
80MeWgA5j5Bwn1mbCUohwB48U+ENBGznVVaFlApRv8pIpkw/r8xYCNYDqgaHdGTW
8QS87xHIVSyDU1cCGT9FsqAhIOONY+jiBVHr6htdt1SfktJRx0/ijxMu23nwinsa
liuqiZZtMnZygBye313sl20LlHM5RFFhjuxJ67jzhdCkYW/yLQ1fdK1A7GUKE43V
cQhWdwXLC5clXrC8AdxThBEQ7Soh59UqnhMGyeqd33+v6+EgKHwOlmkdFnlgZvK9
51D/uDCtuWn82ED5y6Y+X58CMlGg9mp4KcpZbrVpck0iHCMLn+TD1ASbnvoFvfat
zACnf2olQxqkpG204FaUD0YqJCOEXFcD7KJHHbVh2MVVajV7uTBaBTksuIpYrp2C
MJ9du7lSppsQfINhctzWtjrUFSPW7bQ3hc+7bsNfOpSRXxs5icRmY8H1La6RAGYp
`protect END_PROTECTED
