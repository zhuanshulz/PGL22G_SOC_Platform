`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+k4LzC2Lq0jpJvAGw8LHaldOXXgp5pkgPzoU9GyP5kseWv78oZPrTFtBjpfO/htG
9zR8GKzxxqLNxH/Rhlty+q3sYgZqgYXi/QpiW/UL8OoZVts71TxRYl+5SS3N5p7S
nF5T6mOiREIoPgREVa+D12ywD9dbVE1yHZp1n3BFPDYQQ9BjS+Yv/tECW8yXRz7c
o4eUl5X7emjTRM8S5fb/KRfYESITr+hQB77RYBGXjBsEsE114m4e83f10GsIrwp6
gANwPgclUqwOnJVvoRcd8G7kWFFGfjocKjVQbvbtSgmzIxetPtrIxEWuSOzzONet
HeRiXpA19UuVhOvJTr847nwtLjkv9i7a0gU8RAz6al6oqMdnAK7k54wOx2qCzERC
`protect END_PROTECTED
