`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S6hjPMTfPotnaWPPLDkNTizcbV0jpmXPnjy7H0K1/c2FwfpBHx8zDvrjjN0orhte
MFqYw5Ovjh0LCtJJAXOE5VQQ5BtC7UjRm50withuhx2sZLkqGYtN1s2ZQmbRQezr
yTLKM4PdfF4B97tGxJDVIQd1ZibOo2clCYM7gtEr15+nnAuRMkRsIz4eHhtihABV
0UX4hiXalJlj0pAQbXAwwwMxgP7LvILFAee1zCGnycwlSILcMVwHl8bldAB9sRQR
klRXC54nPTdn566hr/B8Q4Fw6xEbxOqY9FCvnSKpPAnC0Hv41GOaE+GxKAqBeBub
qRfv4kGWKMuCLFRAR3xPPuL9GeAQYG1DXd5AmEmMqRWRZSzmcbwqFcNZL6IL89Sh
LMC8/k1RY8M3c74IkEcccBFB5MjtuJEmCkSAmF93SYGfse6fkXeKdaSOulF88DfL
QTcE1c4W0XYhV++vGglu1PZdIXNsb+gDj+O1FuQJU+/VYsGDp0hKU38+DuNVadUt
WwmidLjVy9GA6aR1jaEy2ZkX+XN29g4wtMLdPdA0CdzzPlyQuz8noRJtJgxyMLA3
Y0URhaIQ9QR1W76D5mXgq6rgMBq1RCLksR0AicUr/GnFU+saEL/aafnjHNUQQeBr
ID5XwWjRSgQebZ74BSIW2ER9atOeLioRG7cruJVoswn4LQ65H5ifOhaaHnOliREn
uNYkOWIp8VKVHjNrWO0KilygbYWwHZLUqs0Wxm47w9p3NoJ+MuLS9GvT8TR/HRUT
u5/z+m1eiqMbzaNSxosqkR2j0hfmCrekV1XbbOF38wAhRS7WXDKIu5Kczeb9eY2C
4GJOSbOrcDkLubj9qVWGjq8iG8mPuMh9OfbuCem+TvZNYbo3gYf3tFCUJ761wxiR
eOywZ1+iT3xr8dV8x8nmWDEGvwXHiejKlpv9Qcibpqt9YwHM4pO9j9qJZvzBzYmh
Jrx9e8SvN0w3YwFo9gjnJKgwZ5So5CJodQfhxT8StmrQiSjgd0s3Sk64vhnmFjhl
nv48/ZE6LGDjDq9MfD2Btm5XTI+PmGkxZrRnJEFp+BU6qhMCZ7XnoCzqI6dtETPu
Ir1q2tMwO1/OBC+FZblmd8MmhFhKdY57599IkJX00ousVdQpUXvNdQqRShKSUuFx
wXjDjzRawv5sKiqpSBFTVCIV/F0y8CePkyx60jYEGBuLWimV3AYGDrSUKbifqDGp
4kWNEfQnnSFqQckKcsmHi2KrKKvUMkJuf0dMYrH4Ohs=
`protect END_PROTECTED
