`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JwvfanjTBZhADvbYujwRfqaVP3jVs+nS+NyzYv6l9ohXc68KalRBd96LSBBmwGVx
0UsyWljAXV8waKcqKTmP3fD7LklTz7dIsh8XANBl5yL40W1CzlJJp0nUD2zQsapj
6MTVzWP/KxxkaQxi/u5gepXVYylThVw/W6rqw1VOIO4+dETsjsg2LUtfc1PEgaN7
zXzEy+tHjjbcTjEu4xC/DjVOkT6j+oVeUu/a+iWX5HbVAFs4rKUAVePIodgiGXJ+
pv+JN9IrjMTlZBNNM0Q8HH5NbuLRt/tPKBlj2xk8N2Cz/PhdA8HRdq25VZMLQY9G
Y8+cFVB3qYtB6o90rzaL6/vycfb1WdKs5tiOJZ2vC58g0Poz2PNcSl6Y4fX4ZHn3
u/VHHb/7GoGYBeDrGREA3Dy+Vy/Na7BLtucFi8ZxspszEyJMmFdyCJuN+p94tRGQ
4/hCAJR+sT2AVaAPsZxoRTzhjDPWOxH4vAI+JgYnM0nSh2mxmdJ8rKPFhEVf/EC+
`protect END_PROTECTED
