`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xk3v1PSF6ujBs4RWJQC21Gr6gmjkldkmRcZBvuXDlBiiNZgFqotjntt/mYq5d/JO
Tg5rvq6eCScy8enfx1lcWyv0uP0fmDNK1klOd3WgbNNHEl5NH2xwe29NXPJgS1i4
gRp0dV6gEXF1uG0obN7t2GH7JFeesgUQ+AVGFpVic+odEGlrioKz7jw5RZrDpJxx
9xBvfnBUj5yA0SItLTZhun6MegRGz15eaf35LNmtbgCTwvMDy2t5s63/ILIOq4T3
UxBnwnvuTvw97jlCi+CuT7JLQYK++B2Z0elocPhC+Sgxl4Qy9tYV3YzHDVM8ETYH
8qfLd8w778qc8P/MhyW/8S/Rw0aOzf/0u5w4l4xWHmeXpiTwAi8hukTrDjxu1j4V
Z2E9XbOOlm64Uw5UACm5dARq6kTcG4ZMrZ0WlQ2XWGWQAS5DsElVmM4DyshjGE0X
NQb+CEDtChZfwKb/1Fldh+pr9pH8BkF9M57+MXO6CxgBUANnGtTdgIIRneu23ndR
p2YP0Xj6NX25NHR6nngPKluocjHpQTKlkl2VIAbbovWyoapOzdxRZCxTbHYE1fIC
6jy176HqH0QxRPogoLzWMW6C6iRvpkts9dYXjmoQ8XaiiZ4QEnwt1fEtvgF8PEZA
dRhtLzYnAvQrcWTu3SLuZ9iGJezrWOEiIz2IAJdrdTfBL/ZonIWsIT6d5rstrg4q
JcM1xDPx9WuoueKNyqIj5Qp9lAfNZzDJD6Ky6EVB3XIbZcEGDlIyfmycq40/hPfx
A5KkqwuLdwgdJcEGu1gbw0YAdP9ehzBi2mDD/KQgLoUMG6fA/e9Zq3EjkCpFq/Nu
qwVx3u9dSsh4JgKVle0jyQ4SsvYrBerL+nFujZ/ODYebxMaX/r7Zf5LlYcEHVXbg
Nx7c3QVmP7Kpx4LBYgs/KMv0T1kNfR/Mq5E1YXXz2/Vl1zHvYFGI2IMRRFvKDZYD
8wc3P+9VOVkTVER/QizVjHUCo0ISfWCLV6ml6s96g2pd2m0VIaWLEddzHP5sk+l9
AnZac+m2nNf0Pl8CuyP2nHtQRCvyzwFbAMsw0GjtNkpPzkp/ZVOoqxLroRGGWYGC
KGVU6k+SIIXlkax3WkRUulp0ewTVtHhLqc6zreUjQhVAvzERySqC5jbf3BP5rExz
qz0ecZP2FJmp3xa3Y6oY1y//y96Fq/1CU+F4Q8l7JpsB5LlZsnk2kFZnN09O0U0c
djRkpdNtkN9gJlSUyo2UBvwyGkXuqfzV1jlkxZ34S0S1tuiMQKoVEGeogp7cxfPB
4awvtF/HXQTB2gukbi6FOwaptiauMEiwntQuly2q6ld7RAFu0mhKS77QGtKtFKzs
Ff2GoL84EEv+itllv0htgE4swfk9CbRcAQiilVtU2pJ/+xrBKd6er2FQ70ucjTE3
eW1LJaGRy7tcLcKrQJ6XtNyR/h2aJntOs9FBE8a0ZBpQ4vt92xy8upxxCoPUN9tr
jLUs0gIPtcwJFnTAqoVmzLFipXM3yGsm/lZIVqsirdX0utN+wUXlw1J9PUUZlV1e
Ux8qitOaa3/ltDcrHUlc3BIrxgG/jL0Wgzj+14ahgUikNSfF4rQmmQQ3Ip660upV
vNq+c3DhQumpINuJh22xC9ElzW3FJL4jK0o3N4ny9wFokezPR6LAAVjDMulC1Cjt
7QdjJ+5/zNq97bM+1zYCaX1C/AK9MOYv3sdC2p9BZkA=
`protect END_PROTECTED
