`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
81dwf8GxIr4q0S4TR2olTOXENk5V+Yj4ICr4L5W4NBe5HYSgCoef5tLQNY9aV0II
6hVVY9qQ7kaQUWVLmTJS7O4f08kplGRBUOTdgRvs7eGAMXkftkJOVmW8M1DMIOt1
W/l+OhJ/vPaHaWQRPUVvzHk38EHSy7+utFRReXD01BNyfJm/397ulasNs+umbU3c
Ovkx/WtjgLKYadKjKlSOUn6XIqQ+3kvdMulKfUg2sEluBrEL8IcqMT6jVppUvB6z
s/QYwiJOttpUnBl+lz2Ou+KE0fth2KVVvXDaT74clnU4c2ahdIlB9NETcPIOkuAA
PtJ0v4oWjkeaISxTLiHL6y3sLwwWd7LIV3xfCWBNLImBdj9oNxU/WVa0x5XaA9ma
mfAxCEOUuUpeYkeN3CbT9zzZXbJMecMA7UTR2yeLCXQNj+yCBqtxB/e8AEpCqgWz
tJCe7ByMqfRZLOHgzOGTCMHZpHweIesG2RTc+LDN24fP7nGLfciz7PNbLNrLBDVG
ntc7Q46XZF0JJXwSNh5/fWs8zJMp4p9buyOUGjIlsh5XC+mFivNBmwrmLIX5wID8
V2F9RiIaIdkho9x4bb3kKDiq+T61W8sL+MhRhpPNuPVC7BA/C7s1FnQ4G/kiy8cH
dyeq86usk7kAhV0DmrvuqIXv2snnNANalsK9cCTnETCXK8vp09NWo/wzxILSePu+
eTPOHNiuJ5tbSxuyUdrj2BZkqhuAPwG/LXKCMw2nyAZR2kCEYFAxd1xlhoJdhTbQ
+XjF07FzmUX0tA8c78O3J7BcL6+hDrBPXaC31IGkB/rOThrAHShysHmRTYyOEySn
5ZgMGbGG6PCbV26ijCgnDJtEkzuT3TQ15hoOnckrTSgwIxBJaX+LlKy/XWAM6Rmo
d3rEU5n35L6GmDjRHPlXbczpLTKs7kzJLiOvTpvb8HecbFBzXRUxDhkM/DhFUVX6
GDqbHaU+f4VYtfThUo+GcvobOe7Y0lhtDAws4yR1WOiT6QqZ4sad9aGaIGkdiJY0
CjZX1+Wmw6yz+1j5jg/qGvkWiQ0Wk4wTZozVx5ivaz2saZckhWhTW2U/sfCSn0Tf
TzrPWx1uYP4K0nzBJ4KALGdoScoZMhNTBgpH1gv0igx9Eo059FkOgXBev5EGAMxx
M/41K1ExV5cM3a71t9qMt8qxtXT/Ms1w+/o4xz+IoBn//sH01s8Dt3H4RmAKT4SC
YwLJVt4HUHFEhmDm/1Kzj0ZZomyjROFOU+SvqN0B/4NuV/xPO8WYUPzgoEL4kMfV
hkYVbHs5zERmKtyYzlVEvtVYVbZ5hQTmGyicwY20mPq/VxQsgbPXH2J9Rd00VEtE
X86uOlhSoBFqw12ajDFfCqloQg84w1CTpOYsHxbcQvKnHqlUQosl5vbTdSUruFNe
tZUEiNqL4cQpVNrISa5nvDcbeC/slqUfSJXCqR/HEjezO14OzSFVFZahY4RqACOM
jxvZ2JgIMAvEXSpcPsLNJ38wEnm4m/0MYYN3MHNkU/VbZ1cmCujCrEPqmRoNu6ul
1yN2Uyrk8UL8FUiU55sS/2knfLUmlUrFRaCZ8FwcVid/AtJc3F6NZcq+otH9tnoZ
CBM/ltPV/R/k53AteaBCT/w2OV3CaHkSDjIOtHTSQ97G3RMk2ujf0di77H6sBS23
N/pg22MR1KBV8k3NJva3Q6RhiM3sfCBFL5KfLJbUAfkoJzodA/t930nvQklEgfwx
JBLq1+Z2/0LfHh+Jb9YPYYSvvmmfTRAvTCeba/jYJ5CvQvRvo5JKOiXhFk598Q/J
rx0hemjabbdV2TPSAmBM8UG4ZUq3COwipkBV0vuo2obf36huVg9Nmdj0pCnT6ft4
wmDPX+1Nqf7G87ZUO71udZ8OBzgujMO+Yt09uwv3S3NU4NOL5opyHsUr+YxYeS3B
fbjcqGIbFDWC1njJctyhPBF1eAmNI8sYLoOHJboTmcVptRNYJ3VoiEeP7lJ2r4GB
eAXl2lAeOeR5oOMlaQ7tfU0e4laMncnpbk89RX16CEfv6Pn7IiWmJE0VWGrL6Y45
HRk44MpZx4sE9Bnq4xrDlMJYLURx81W0MGPLOMxWegvbj/wRZGk6TL//ylVEQHkR
khEg1v0+KsuSckuZYjNpgzq2k8j6UiL5PZyud1UPNzekbjs7jWB4dVKDnuhlJ+hD
7cdqsOn9SthtkknDcl0BkwlRZFbpBxo0M9A0gbGjQDKStR8GMGLDA+C1RRXg3/mS
I6mdZeF6L+FxfQ6ywGvtCJQ0ijUiPhrdbJvv7/daDa/9dhXpO2bD7U/M++/TwAJu
V/MCaxOdBU9jUPACH6UrXWOWNwLzaWhJfAC0S9mkW2XISsjkOMG4Af7Uf/GQvP+w
04/tXHd1fvtJtrBx2grW8t2PZhwHBdd54Nix0aIb7rCr9+yam9dTEbkRbldF9F9e
f2MdodSe0ivNreZ9jsQmlgmvKt2oErtXJzlRb6JbKYHhkBV3fV2J38ZeDEBWA+1b
UBG6gThNg4+xz1lt1fXAqXRBp/T5ieHKBcvF4GBIGlNK1UoYEVEun8TaZWpOYSuN
7j7cT+S6f657GXKAIKmWpTgz8GSHVT6ANFyT7aOII5eY9tf/CJM7MkcxhqE2CVUL
ZmxI8+Yaq0wnLHzznVgcU+YWgTOnIpnSH2mYXFb9P1DjtKidsTNauHO7ipTWi04m
8femCX5DphgH4YAqj5ZqDaxyQWssFlvict34ID6UC+rvNjaH63GteREI2Uzwo1Au
u/dT9ahc09g1s9GA2d9n0KfI8hYsoa6MqOq1nKPzuH//9vgOsn4yL+Uj/1y5ohdI
8mwEG9wmxCuosuqn4w6jEALMk9SoMiNfrq7JjM3N/7EM7J07sBpXj6f0rYPWv9ph
OPCs3zQZjVNe/XW0ggW0jWD5VL1UPr8vTuuA5WCWz+W2K+jjHCccLmZ8iAjf3AG0
FdD8XPNZQ6gGazskF3P9ARucnaUMZctWQ/LG49nPPLWmHftCKOa5uuLelgd4Nmm9
3bV1ii8sewc1GWTtncYZURYLU0OnSBfklIacExQIKTBVaiYCCxCsfg5eF7WAq6Tg
/o+wQ/6POaNII2h1kccplctZs6Mm32nSKCIBhMfcE1S1TwBd/pquK3N/CDeSDR7m
QTUo0EbyYLa1zReALOyrEA3F20RGOD8+i6c4/nCRlzJ2p3bG+QmtW7pQmDXFgDUp
+96Xkt5veLw5SVg0+jnIjXg7C52yazf7C65uP7G2t3XY9N/zWVUhfNAsO7FPsNn5
6+gKGWuopb1Ks5+Ix/FUmxABENkEJf49cL4yhmNnAzkBiUNdhzVE/eR+xA2u2cfi
2v4oAJR4Yehm+Co09d9M9dglv+cBRPp2H6sHhVJC80QTmDamOXXPtbNzjW1piqq3
bZSg9bmY+7xDExPkRrF0LQtZ8NiZFjC0fH+nak8wxxEE/OuWfboRdWzZFH7BLjkQ
r3qK8f8S3Nscy/Evahw2PBo0Bete3WUQLxkEhowk/uXh1RHSH5FwkZEdGKo5Vssc
RoheHTkuaK8IRbu4mTl48LW3Dwzt+qlUfvdCNW9ejqlYCdwLMlZF4TJms+45aCfP
SvRf2gWgcLqnwXGpcnTHsNnh2psgBfp/i7nGXgJMpb8cMjn/sBrcu/cBLOB6IJ17
ZoLX6rISZC7zfv5ZnNpRAn989Kn2X2srpH7TSlyNp/6fa2WCcCVv4NcJlgcxyW8R
ovHp9EiHojU1JwqetT7vqIRVYyeenPf+zwiBMglsfDu0f7Ay02LGtPxQOUQ8+m1H
wExkMVB3PL3r/tU5hZFGBBE29X7bVy+b19YibSGqHQgwsBgXlQYxf3D4915TkFTv
gcLMZJaQx1veOWA6Yvy33BgFYQMkmHhNNHll57peQaU958n46mLuieLcW52Po1Pn
oMsdhv/crCtv6GDVSlO1yA0QOo5C4YIoIabGpYKIAnSvzc+uLwdfaXfyaz/8vz+6
bEClLb/WoS/wNFLICideghybfPr3d+FlENmY/JPc0Qq3/1uIfC2agDn7fAlTklg6
jF3fxXG+QixWQwTmUC+3X6amdsB8PKR079AVyeI0TEB0791zblFKkNZg/b01bdBH
6ZfYBngWkspmDrWxV19kYqi6G5ZN+CIvbWNdRyFs76+KItY5EOjOzIRq/HHYFVC4
XcVNIaGGuODZx1mRY5DUeWeFTDGBY/WxdHQv99EbnL9Ys77UsLsft3nGeEJdMBui
Cf4KLnsUCCOSOY1AyZ72vIW2dyv0ETnoZQKQSIakYIEtBATSovTypbQhOMPcFuHx
sun3wbz23rE0mMsPydBH66a1uqoGBlv0D7DBdqc3W9vZDfAKPnzAdSFrhky73CSp
uQD3Mk4XPZGhxKCARRUbwvpwhr6yaBXm+g6gMNI0yaML4iISpp/+cJ+IBFi0NGbZ
HjdrqhKUAhV2sZB/HdF+/yq+QaVr/7pL3Kb9vJLQWjZhpsGe/vQbxm9cN+NL9kwl
9X4v2hdiAETZk7V3ykHEsMmJPCXeLyvPkZA21FlnysqlPaC6tD1Rmb9jhVgEKcoV
+JIaj7PxGinypDtcSJjwlKS9ToGc2+DuETRC0dojyK3r7RmYn/fPFV50t2F2Cw7P
wBqUvna4Gk86IxZUDeFTGFEilSqpWgUeMlPsBT6/eFrBZqFybZF4MAHFucR6nhFt
CR3T1dqS5znh1YNy1XSmK+ryEuLAA2y4GxzdNcGBZgilUqJRSLzGHyJous1Z3oGC
N/XShGMFGcYNcW86OeE34mkMLpQlumT8JINsijioVC7G9xCJVeTuUwtkkqkFYDD2
58VBiU4zdD096MxXr8ioeUX63vjDZNHOiRYyexR7WXwf1VrAuwpI8cc+1ty7VWm0
fqjdneHbW2rLZBFh8vpBtFiShJLNX3JLJlA6n49iSUm6vVUgmu2SIOmaUcdfp+cc
v2e8PRv204aXp55z2/TtetmfrAPsMb7v8aXYrnjjwpIDzslsuDslHsyyhtbUS6zG
k28YKvnQMpg7XtsRSYZs6uqnOLnJSQgpTv0jfAXxUcscJudnYJq2OSIjzNrWzF7p
shcf9bSubBc5Sx0p2N8VF6t4hvNt8dhnT3ONG2PwKP48LZcZQWPTs5jP0k5zfjTz
Kl/C4W7ioiUNRxJnI71oQzs+BP7vF/N7r3R4EDH6DB7/LCNCdwYjRvEjbmBIGEca
bj6vRGbIBgALqHG6u/3Rc5ULXaMVUP8Ik4gS4umsStmUw8YKfS72nyiL5LarfULg
0xNZkXowGFqMCGTKoZIaRfr4C+EcRAUopzYtRQiaA/J7GqyFWBAO+NKwqcYWganR
d9M56cnpU0Bx9m3ofCDdYfaiLyBRG2cMTXyTx74RZYzFpzavX5b3W2ht8Trowgm7
AJQLhoaSak9Dvpek9WLO3q938lkbj/SMYNePdvVJ2N3SzhAHarXQtkduJkzvj/sx
WTKosy8AiXtnn7wzgUZ4rzKOKvEyDTke66V5+6WQle7QKHP8tLEYveyVX1zhkDpk
asCYkDD5CRHldMFLiy9hGWliPhbJJbbZ41Jlt93+jQ7v9edfIPi12/U5bunQy/Bm
WfcpbFNAM+oc8Ox1A1xuk9YKtYuYxqeq0dbjQa0zWDTndG4ZWp5Ue/itOID4ENLr
bL9v1IKw4+yTkc1u6OWRTPIWHMof2KvYjV3V3vV/GtlFBZY0gUGtIVum1+K0bItf
RWmU9jJlnzo2VALIIsmVCm0cf2HOl4WBKA1wNDFU0F9G4Gp+ipFhe2dCydkl8Y+J
O7j5GUJmaYcxLivqfXtDXbwpvg+kPbnDJvspFOYE98pRuyo4wbqFVhQFTj6/xwRE
WoCKKpRXCDlWkhyK3+b0la5OpnBX2oUFye/e+B2TycyqSSw9g+/GV1YHR3nI4tso
4ZxDA8f/4DY+iAYhZLTGPCZnVp7JQX1dgWLAuUdGi7FaA32hfWYTQLTchkfvAcmM
3dgvA1obny9yqttyfN9DWsI+N1BzMDldkpHuX7EhcC0I6SjYVHR2e7FYdmE7gavV
V8wr3bmSanlSqhxBz+HqrMZHhndet8yVqyj8pXdg+oRB8issFO7QWxr5ZShFVYK3
iKVvXHpetXs8IntMlvr6FRUVgmMiF+eHudAAg9BFw1U7BXqBucyLzEmVuc/RzYjt
6l2SsCurffFyGQac2lCl7XIBi+XVehkWTeWNopU+NXPRSYF1asE54qKvXqPnZ6wh
tKlf+cnQajO2R0ToglK9AzIoHTsNEnTYDqCo9D5DXnCFaSjqU8bhSPR6KJ17kSjr
rHDL4kwMRoajSVpA1d6wn5D0vUV+8YVp8k7RRBBsWBBLWjU4EEyVBhDSpkGO2cM0
kUczoxEz1aDm3JkBPmRnSIZtQJ/yzzbq5A1iIDm4wwD+Iv6a+TLv8000Ibq1h4cQ
epjWMgSVILdv8VVDoyUkVPBgTNeVCNNZrKATSrZjp3RtUfcnOBHBLVO91k7Y9e4x
3CPZsDCPcRhBHHmgpcVPBW106ZMiNj2VPauknKyL2nVTUxVrzWwKMj/keq3wVr3X
46bULvuhPyzFGM5STSEWJOviYHCyE1vZKMUixJqV6iW2ZQnMS2/kDBs1nEkcqYmS
Vs4rUXH3RFPN2aLp+aqQCfK7kf3NkXILEZ1y9s961z4MvWYf+FyeqM5LB4OLl5oa
IYc5B8BM9m2j8nvobTw4qWtek9NAMDeV+iBMBwHlKX8+990IabB7PGuef/KriFV9
ANM5yj31Ds18snEdiHDA4L56/HSE54wyk8kAOX9D1Ew4hOhjgbDOAR583gPH3Lmf
5nHB3FAVP9Bb4bsn92ljWPXSVSrk2NcLIccTHrxBtDw3DKjZ9afOg5qBSQJv56o0
kc6L+yMfarQsGNdBmt25hHzVbBxPQn52w9uk5LBu3VTbDodC4K5MNRNAaHns6dVO
0VppYpByEc2hMatkLLVj1rgnsfLtqcJ8ay0NXQR75wML97I8lp941K4rcGNjriiT
lL2nzvD/t15tIwcnzCdTqWGHfaCAAWiXam2mbgbHwJwDQ/oN5795WN54S4xFnjqo
kbtrEXgGa9untQh05AftyOCzFxn7bfZxZM/+HP4QdXCDj3IAKH8lGXHN+jbX/cWH
AnoYrltUb7KsY3D70bIQvuWt8WpZGx+54ax6NT1f8kI00jFqP+3TtrdSsMqgDems
oMYmlaYQkl5+ZN99U1cLMTkf8y8ouYFJLe/wVUu45m6hLBzzpRXQfhbizyJVGjY9
3PtrGvs/P8zzEEzhJuU6haL/OvGNreHJnEa5by7+GjWMieibz0zWNfK15gAYvXbY
hOJjtABYOrEapv4x6/GvLZQ05aV9g+5LA8bMOowqUoetTl+zk+OIDPEUOOyCCRNV
yARAndz20iAORUz1R34v3vPsEwRwMoGRtKeQdd2/+GxnOVs9WNhDfmneJCfOXRy7
I6YCrasbD4bkQFdjh3P0JUhbWgboL/GFoza+LYaJiubl0NM94Bl2TASXiL0gbtoU
WMklFePJyxwnLRxpUA63E5im+uSm6bi8xNnxZAb+ut9Mqa4/LnAB8fIrG29+Thc6
oQQb9oUGQQ2SDrV5qKEAXN7vIosMUg74xBL20faKsTu81iP2lvxmGMSbCWvR0QyM
3BZoD/AjovKjbaWKHmlHCw==
`protect END_PROTECTED
