`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kiz5eO4t/RuMw69pdLVfuCvT3Mw8wPG3gFlYKZhYTw8x83T0ZyuF3ThpehqBEULA
W4iaWp70KNuvrZzGtZaF8aa3sTl8DrX/SKQCfRIFXPHNb3TUNZwopCzk0Ck8Fdsc
+vmmHFixDKEH345zJGrZTSWAi5SG/mk2Ui1nXvAA7+BxT+5Q5lhBh+6/Mhsf1Bim
fJdYLeadoZVyh1e3OuAj2NiutTLOhsnQDj08/VtJTq4zKuPEUSCTaQ5WhzDBKn2y
/xK8KLBPXFGp88FgLT3m87eyV+sH2Gjt2b68C8Va62L4Tzr3sYxK9t2z7ltDL+Ip
Qz7yjRN61Lwt+wlw9E64o8mjWOMTKkOdVtpIWuh2Wc+JaJ37SGo3xPYeAYDcOKVF
36AsILFIewZTHPS/jpv/UqIUoiGKYwlxFavg1H0oRYfUUyL+a3jYseqWC3FeKQ7A
J9A+Mmrvw2YbuJk02pAGPD5jG26uYeMlMFK+OTuCplW1lfO3pk1j0iZCf0uWC77A
g8TPCkbe/2byRmWXynS70tyrjCjdqG5WNAOTaDU6zps6gx3dtvDIX/RjP6Wk5/yN
ASMT/9Wt9mCZVJwMU3QNXr+cM7MIG3XrYf2wZSuCXjcJWklEw7SntIY/gC5j28vz
mJcpV/Vrxzs1DZ5yf1MAZJ8WlqWDQmfQQNvD8j09tNIXHs+ujuCc5k3k560JtWeq
flyCSuAN06UYb1gbf4SOGoF6xKko0S+Ad1nTfLapFa39dNtVdx5IMbdFx8dYaLBj
RysujNk/PES4fUDYCkWGVuylUVDDV0KE4crSPzm4yb+sFVWG+JDX9VK8siqtu3Mk
/VcJ6N7fA322UF4M0xREstO/MHbhRytyX7tkJzukL0XG4+IXhaMQalZl0ZYlWJR4
wtDetFOEKn27gq1nQBWNIaZBBkU6EZxsJ5M3wW2IIBNNEjtRVamJ+RqlI0MuMT6Y
SyxKejd9NXojmT39QcbJuvs3xFf2Mt526kOovEwxC9B3lvlmRoqy9Yi2rnfiJxUg
1vLPK5KZUZIOSaaHXFlcWPFL9KgbOvV6RauuzVlRFZr6Wz5r0CwwLgVB0613Z4md
E7xV62TRPB5AMetbBU0tfqkpIJH4fWL3l7WwOZe3TZdv1nAh78cob+N7dx6saQje
3cYqUFrsojIEUfIgq/4QkHJL47aXmRxDLnxvPB2RNR8DRuYdMsXBWdzPD4UIti2R
llb3EgOnfc/nGPN3zuMaacO3m95H6BI1iyyNorGdeyiRZ8+OQQ34PIE14PxB7epD
S/sVPlY6zYU3/cpdBwYlKq3ra4KvtRbKbRSTTRZG/9nr7HzM4btGOGXhQOy48dNP
`protect END_PROTECTED
