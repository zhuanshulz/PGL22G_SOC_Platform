`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o1rlRf63kZmwBNNXlLPWi4BNKMIYCc378eQ0GQjK++1iO/MN09QNtZtA2qlz0znX
cEbJF8HHkiJRFcYrVJJ/I5ZM9UXK05IwJaES/OsgGZ5yaxHlTycHl4chUFtUsakm
6GfAu4amG8LlIyKqw+X6HrH0q0UXgiWJxSO8pocyte0mg+ug+Zq3Zgbv3UByO5wb
keMFgwMqaSiotrgufUVBb4l02qC+b4VFdIoUPxqeG23m2w7DzNn0SByP5E6HIlgz
CAK98/uKiz2enjNNCJCejsUmIonr1fZ+4HzJ2X9S05ttI0YzJQnKRqCI5uV0+7/9
S6Iw0aISZgI8xHeIiSQnQ4fl77qCfNahruxmtfVf43wySQLS6kg5qrPUL8zM13JO
jS9LsQFvI66PuTEICdIJ3XtCMc7dFNJs+WPzOGYu29rl1lmvVX+wkzNfQ3tjH10k
`protect END_PROTECTED
