`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WR8JevhtGO9x8KlgQY8cxGBFTIbYHLkjwKyPBABpoec7IAqm95tqHsGI4UvLShm9
WC4JI+Qs1PHZnB4ZO0C1iSwMplcpeJXDqYm+tKRLGwFQ+Bn2aMSjgol/uTUUpvMW
FOySfKkWKKeA2ygSgvGzP7BDUHRBq0UnYDCD2tKYcHHoX/fTZLhJFqc3J1DD7Tar
nG/tEbyng11t6OwB4GSfxJRGGC4yk/goKEGc3fFN4E45/zl4nAsWyEVQfQqgUFjG
LkGQWgl2yCxJdybMwLZlCaUmv9/EEEAev750Au2u0yNUvimoDy/eIICBIJnopfG7
AlF27qHiQGwooYInvAR+kzzQ/gUnzwdAwvkY8I8KB1ANLL9o2zqj/0xqW1IRwsRz
Fij7eQkxe83TxOGToWMI060O1GFV5vVL3EAeKOEXD1aM04siMyvkC1SQcCCPucNP
xH9F+ftulTZpwmFRjHcELPwrfE3KG9C02T6FJWbI90HIr9b5EfMXnTH9o30IdTDV
yXaE97iIho6YyUjB8WUbDtiZ0zjJUsfuSYFGKeHjvOSDzSaCfu/g9IMAxauZobtv
bldEcUZ/GHo1d89HozeLIMjjLWV+bW8VDe0s818ZbrUD9V76fcqH4Tn8wTWcwfFM
HxIyyq75LwgHRSE2wZu8sJXY1+PNkHSMnNmPaxpSOGyHrMH7iR2HMtuzN2MY19R4
0bDVS3dIxq7J9RZpqdQOa+Ay8IyRPGpKc8qkT+GAOKXWxdjeA4VZoOaWpXf4REBK
x/1ikr1t8LulddqI5fBshjvn2YiGR5+eajXdkyh7UPo4dLYfLeSPZGh9z/ZewVc4
WlxdbEst87SwE7Fae8CBIw/MKt9HDAGdE+I87/9rcrvYA9dG9XkO7G/D9JyOFM7n
/Ie/y01lZ98dDkPSzaABMdmBDbxExbu2/pMNYPYBUCxEEXoMzghrqJ/23TBQcSw5
SA2nJ9oN7fQM0giURWvbtOxqZtNYh4uoHB4/A5ZWz5NIE4JYndl1KZPLGtXT/7LQ
Cw6/MHKYlkSZORp5LRNp5AVx2acdRqeXKHrD1b2+swbyQJQP2jGNSpnLYVinekfF
88/KnIrsTWQG4Lsyn4tZSlydzhwqYTZcSGNkyzdp9YBXD+3fQ8dQKxhOHZehfVmF
51n7ZgzmfkvhNvQUa6ccs0bKWM6IZuzaCqxNmCS6wLhz7BPiL3yFpJIn2zV2lnsd
ItW0XOtFGc5AvnB/SpGJ7oCVweEhird9mDJzwD4qNRCcFVJUDA/i6AHZzTmvaag7
I5DpG481lpwNGWKSXjSR+TWLpsqvT60W6F5u/YKtyx9erYRyAHXUEvqp2qqReLV3
VkrUuN5G98XHgiyvPbNGxt0HIEhr/kQymZlzbuHBogmxoaQiStvpW0aD2XaJciTj
GUPKn7sV4taJ68zgNZMywuF4K3YhiLm1hmDqa7IYQ/re0tDL142dR7LZyUb6Yhc5
q5Fp3FH1aanQsdmk+rLyVN+WTOmbl6hEOIGmUlOvbBO5eSJjPRoIbzYtREJrKSz9
L/K+Rh0vIN0yVV7VwjmNIztiSZ3Jf5imcOdpIywsm/IplblnpYBsD+Ni94hrK9fb
ql8EOfDgigKg4WHECPgBFMdveRz17STE5cNmkj2e8DmivmckO/U8vFJI8D19O+bA
B1+hb47Pic7rsR3WZm/BtbHb977V0Lgr5E3QvfoOtFw=
`protect END_PROTECTED
