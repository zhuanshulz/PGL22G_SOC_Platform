`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wer9KpA1uFOytWS1sf0gYj8DYV+4cB/yNWjJNdmNdINAHAV0MBEIeon2S9pfIppS
oXJTLfqsZIVLpsnDZGlQIRdCMiNamgvChrgp6+e0Jz6aH0iHkTYIPP+s2xqZh0LO
WiISkNsyMwMaQf5e9QZ0xk57hUC7qQzK3K5ieBrvSmS4Gf1qb+Pr2E1s4tqizh0K
zcicajPO3XmTf1mi7q4a5tmwf4UOxAkmzoW2g7Z5jguBiyhTWF/Sp1q2H2kB3H+W
GkSiXo7KEY9FtQIsT7/7dNvQdkmcEWmjtFmNHrnSVm/e6+DDBA19qMSqf5zCZ0Zl
4UTT81p7J7VZjPeadA5Jk72b2RfXKYeePFuuCECB7Wk9mD+amu58DGfsjGqbHDPv
NqGJtIdfxaZS5izxhJVHrlDXRfsh6tnC9Zrl/zAIqrl9E65EHVbgV30LbVeiwU6E
OWT7qDfRjdjMf+9Dhp7l3Ppycmj+U/LSAg6JgpHcVfw5tLYhKxwOn1qe4GwxPV9f
Cps8/UdILyd3qHEUo7OZtDucNrPS12MCDSZ0B6IaYrklu6AdL4yW+39XiH553Usb
USaV9DXMaN3ys4C+qmA7eqhV27kMNUvRH72mUru7xMadant4IYntg7P8Hp/vURNh
Q8wVlLth70gMoY0ekgRpfFovjQS8i1dWgY15DmsUv2Y02cEa8EBIv1znD6XvAtgO
AA42M0Hj0hNDgNO1T+mWXG5rRH9YblJNcNvGjMiJeFu6cpDO16IpAdgyXv8Yo9if
F6xavXc7e+c0G/Q7f3EwT1mTu1DHa2coCFZjDdGAAKpBvEq5MqJN+UJu5eqZ/jqi
xpFWDXH0hDPJpyfMej6gneGWmcIK1oIErYeozaVhAII1wcHZ6+c8V5MVCjUSQ2V8
C0mRNcWycgUIf/33lcATM4gmFb4mn7cQou4vJsbMN8aSKOPeEE63WZbE0m46eIWK
PwAdt9316mwGAqVtcRDBkaEW7jwKc0d6TgeQll3XT1aw8Bpym50RmvHgPjOWwYl3
xfXM2PF2qoxgwJKOYvpBjnZpGTMyPWald/9Xe9vtTUM4v7FplNRClKAHOceeabd8
MDxoBsJYYj/L5HGyO5WxrpvAnMt1nM2N5HomPn0d6O+GcCx6Z0aQDYEMjoScPDc8
IX6nkG0GQ+UM8wkPAw/kGVHHNdBoFGR4spBLOpwGDTbP7wn0v5GtrrC0yk8xP9T0
Ur1qs4FjV0Em0YdD6baTtDHMUKkzrmpxQxnpQonCWDfu48ymFxIrpUoi6PMfwQMC
5GasaEQdy9a+VO94Ji5vLUwZROo41oYIVhNf87K8aC0p+7+rKl1hVHiTv/lQ79S9
YRw5OcPP4oJH9z9CQACH9LizVmud/0llMZp34JshZMz5uZBfcwzdJiYv1tSHqdsh
S1hiGYpQ4WFOpqQAupGd9DmleJhLJ+6My8nyVjRGWtKmuq0+IFLJ3oSBhzx+IGBO
5CbiQPoyLKkx/wZf4LH6DJgtdqobsbNjaHsATzmvvj0pH4P1Wp2lBXOLEhLo2aYw
aUjmkezMa6iusdorsFw8yXedsHF3xb9joKZ1RbK4xms9A+c26NwMCwMh9fhAIOU+
JqKYWENxu2WgCmJ7c6TRLfah+HcyMNHRg2cAmMVPE1ooafHDBFLswEEYFTWdP368
v5h9+1gGZ424iXqJeiN9np87Ky19SilxcLCLJj3Nek5qv0ihRtTpRXQCLlXeUJ4a
j5uqnKJ2W9MkKapE5GJUdAJlSuw/7gY0yhvMCEmrn+Gzn63PvI0ia0WP7QpIauql
00wCIvelucQqnicxymL528iFgmukBkHsjNiQCE29GPx7vh5qCcsw0A/J9sPKFvts
WM0AzS4CD3Tv/2FmGfuW9yZnmyBZSlL5HpmoryAH6d54ansknCOMlKRwQtEpDI/o
Prv+UC6UTqrbdDfXV+zXSd+rhRkumdI9BKw4Uhmrevemlt1MbHHMsmVC/oheIgUc
Kk07AUZ44/98ngpB9MYdnVYGtwJTVnB3tb5LvZzRDPf6PC3/E38dOwmjjvpWAUe8
+WRGodbcuTE8qCJuA9cCmw55CtCCE4+7PtuatzIblax5+WJfimm6GGwMvRqQYoPO
8UpAfIOELoXTJNK78v0aJwZvq0xxsQqSiQjNOopoj8KffepYebTgMg5nQ71hvi/v
8/bF9SLmkJu24EjaI3cBdriRH3oHTfjX5WjmmnRCf+TxdrKh4unFoNuIwiSbNa6c
4WuqqR4+lfxMI5KRqXNThZbKGS7GrWimSEK6a6Bls6Pxf6jE/X9JJ2jFNCAs/q4Z
Xhkn+OdItb9iVgIdkn10zKtM2skbIdJqJ4iLAFRghPqZ8BhG0IBlnfc9VJVZNs0c
kizIovsQ+FMC0hsj13VFme5wAy67uD+I9KHf97CV3jCub3pctDr8o+DQlsZpYauD
wEbsUKn53VFhY4YdcmtwlE5Qmhye6vUONh1Ap1BEfqlElWQoumFU/yG29fZlbLlL
9TFsIKtNgpPE7szD49lqK3kFOrcIANr18SLbT5uYOvDObmGdJuDVQBJvrhK5wMo9
O5W5U1sHljTwaLc4dcdPISKIrZJs+0jBrWYbi20t/Gki3SR3dOqrjxpmOOJNvmyc
jg9/hjZ76nEU9doHOiZmCw5ttKwbYcLDR9mtRF2PhMQzGJA7bv7gzfPZ41hbyxuR
eHV5wNnBk3PbqP/IrswG/uIy+n2pYfvZXpWJg8gjy2XIgUODEMbUo0QY472fG3Xa
Wicx26juKmpLiWQgWufm5qN1gKglKHb1jTR7E8uV0XmWZkfAPRnkZvq7LxsnftoB
mqYbZSpt6JcJr4Zffc8iJF21pr+LeCjXWD0qbybR+s0SqmlKCFPINl+jxUdg5StW
rlNIWhFiN/nh69xB67xSHsFgpSVNWg9HPWA974QU+mN+iJ46cyVx6D+no9uwJ053
D4zcOg6hnq9dXNKuRsD4AjmUdK3bKA3BUDaydCldaeSoyImCvQTcT2idkMzMVDh1
+3MjsA+QPiisfocLIwMeWdQ1e6Gjaa8u9zDWndbK1aqhRA3z9fgRxJediGPQ6LJa
zffYtsCVRw5uIvvNZX1CcZwz0/rl0beNQKnXxO9tdTWxE7WWCuNi32XWscYDc1G4
enpCtJKqrqzezuv5qklcHQTGA4LDfHiyh2l723M2AVd7X34IqYxTowtKCYg4naE4
wVD869D2cF8FuZ0A+T6ZwKKOm5Q3WNPAecrMlR95KF6ud2wltWgE5gMxsfZ+mFw+
fakNJmQX0jPpXnerbS7NFDBJpW9CjEO1xgWmAoKO2+EjE3Vq3/63pZ6jTWat6fxJ
xdtm+50sYhv1aTv3ZD04QKy6Xvlx19UhlbGpJV+oDkCFAEcug2kiBpVTgEoDcqA/
3g8Rxj88Ikc2R5RKwnhsaQS+ztsT1r4BIJTPKIG+PCOBruDtSEYqeysfMsSV3PIy
oPlpdLVBz/rW55dPYTqcDOmR/dtgYtGs/N3OkV3RkGeG+OJ8vnbqCWVJKicaWyU8
6gU+WcaTPJOC7FIbxihMy7Wk7F/DAQGtp1QsG2LBeollKtlo19Ejv2LF9uMaqK2g
vHRXInb5PLhNT6msBT5Q4KJ9V79XAbrphR4Ilf4lqZBBQLFozVaEWPLj+Pa9a9VM
h2uGpwFkcSfvdBXHQ3Uv+BUZ2CDQ0IWzjFbA0DlASEiR04pU74R6eNT01CiZtFqV
4v7Dt1rWp07PJHuO57BHPHo3Y2jv2Ht0I3dQR5ICx0moJXxsyKTeF5G8b7+W1psP
xl12KxBIj9LUCLc2Sydz7yd1uMLKUt+LjGVcq5zWrWnEIELoScPdqWAk4zWGMwAx
AETEPHpCVnP6f6qmEqqCOBArE7PwkIeqGuuu34JvnKMwfVKK0IaggPj3Y13/v2i6
wfSDpC7lF4PV30UqRXShLaUHiK7jjEHr/Ekl8URICJ/bEPHL46M24BMJTjaS6cUs
bRPukmYTBvgtLq4j68fBuR2yLmWLqHS5XNvSDIF/AZQo2wVys/6omR9F1yYGBzTH
RFQfC/6359d5Hn/wJ9kYAlT2O2wQx6VpBaRKNKjgf5pYEKgJJyEs+iC64/cRXHoy
z2bxvps6iFYpPRxTvo1fyqgr0/MMk6ejUkWF6d5aFmc=
`protect END_PROTECTED
