`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jtgfcpDWHSOJ08jTJZWjFtk/BJj/3SHRNLrfhuN7kzCFUOHffO5XHyQYR4oCRe2l
N5XU8LX1wyY+OmdRDEBMgOpzcd5B9WafxGKtZYfXPmQq4sV6LSSTriY3CSVW5JHV
zG94t/RRN6ULLtFsJYsWxSHdfXmZKpqvme8Cer5o3fifeRYuWYiD+mOguxQeHFuL
DlfwVnZFLoGrY142fqphIMiJJ6+GrCYHkIgflqA/J5/5KM153D181/ceMe0by8sL
J72Jq8HggdJLF7hlrqFOxd4IkVkA0UeJGj/SvoUtjR3CIrfAziXK2DaGRX2XVTae
Kz2YgQ6whUPX0V7ZMtwFCBAmsY6qnSQNV6YB9QKPDezGVmpOLfSb9aTDETeGqUpO
IboKPQtN6+VANsAwKPwF6/CqtMRPRSVqE+JAV6OwCOKgHwTdgnUo5tozCr/d3mtu
b9l2phoujebTr4m7SkVcEowKKAH88PnIU79xfKT5gvDpuXVTf9HHBZYKvXv8+bwM
+hB6zbCfpeQiq6Ov44uic3lBwdoqCNbl96ERzKBT0UmXYeQMTJPmj/N1XpomgW5J
6iOpgzMJpokSY+VAwxjrEOTYk43RNpN7CK6CrEiP3onVmkH8UHtpQs7EpIvhDu2Y
NVL6c6K93s+jfX/V0kCbr9P4Cg08uBxkGEPl6SaPUcuDf2SNYiWO5R8nzP7Mq4iX
8VNxEkG2IIWuq4jaRzPDxSSYVBo3DSKZ0N/en4H1GbiSx/diCUJR4MWnPbsaxh7m
YnE/0dEyegOLCNCYg+3B200Kz6lHF7oOgoh2h0w2EwUMZbhouTZTPiCNF950+EWF
9mh2AXRPcr6fWh2WRUUmzkHQAk5mrA2Cfk5hw5F2u40bG/b36/rHWsTRnpikF0Dn
Gr9nGorLsEI9tQW0e60oaWxADOssCKFTlkjfYJfKyhnCe60xmXSOO+dtF0h8vN+/
yEgyBlUxtvM8ibfmr5wZjlkYZ+R1alFrnIq88Bk8mx/qonif7vt54VV77GN6aD+W
fKtX5rx/YDpEnLw8RCrQhi2wsTd302LntS+sDsozdWvxV+NJkpB0SABnuAftFJKL
lvaT6eGz8kqIDIJTRjtq1Zfp9Innaq/8itXrmuXIA6Crj2zsO/jUqWajAMlrUEhp
YOQ+f1yRdd2hijnF0KibSyhNADuVBkP56EH+OGn7EVxSfmNPHoTjxmMAVvKcUMZ0
6tEemgMsktD+ZQ5IKghzx2fiVb4OPrgRO04flm6U13oupPcK/wxzlMpBfrEWkMNM
wNVM6pleVTtA3k9d+wWISxPMgy0FUSa1aEYaG9RPb4Rj/Or7aDASI+1GEVctVJpB
1bZYFwD3YMTV4fyM+3BX47ZYYpcOVWS8socDAiG5EYGnVzavtofdPA0DhWxHeIGD
yFIvChYAsjVD15d9gDprUyyNoyPXtDsyb/lVZvixuYHC4m0+YVUYu2OZVSzrgSf0
9zxtUPuBiYGFzaFvDX5WUV2Jl5f0QEzKiL4WKPIC5TQShpsioYsxWcK9bS7AIZZ6
Bjw/lR+E/wC9TAxcFYTwuWm55F2Vyk+sYSU8Kj+8uyTklM73mdSiXvpdcQkmyQPI
jVV4uXRzYlOUfZNWRqpELM78/B9KO0XUY98JViEo5S0k6ODN95hkozK+b1FUarSv
VgaGnhGwulwIVt8wHhKb5BJw03OYxOUaTlU8Omar3XViYIOX9bybImxzOTC/e9HQ
kRHju/0HuCWMjcIgm/Dy7Ga+4GwT9wra9323N0GA2qKmSFwnNvCSr5Fuqbn+x6iq
AxJTm8q8zVyV4x+gPRixXgcwq00yg+QT9AvtYIZpe2LzDEw3rVC4/nKeIvzwU8SW
j0nlbt24X/bsxv1Uk5wCA2/H0YDuhTHtfQ/o1EYOzkMfe8hFPK8I71n1RRXxlDRI
cvmptsHxZhUypk98sahiEr4pUIMNf+jwqY063sYrvESBZbvr6alPK/Uhpmeqf+9t
tGBeV5RBoKUipktVhXuX47dhEwp1suw0cNo+e2fLCCk9MUyrJuzPPohffn+6ffk5
fWZOr6qwGw5HPyhK6LTQzcIQyWvlhhxLWqAhfD8I/yOaZda7zrHNdLXoGztr5cI0
4n/0lMHFcOV3jaA6Jy5PTH61G/6FRmOThTOlN8PsyVe0vvhHUFWnfGo9gZV9QI4O
nDTIbigSFYYXUOO6rgZi9OCjFT1HHSTvE8mGN1uBSlM9LPbwV2IqQ6Saz1XmrDFa
tSnYPaivpbKCo8BcvaB97Bqi2i6aCD+7I+3f+dPFOaKyKNcAdlX3OPoF0Rt7on0X
dxgL9Z3PJGxN0tBiML5MYbgwQI/XvB67TuWJFvJhIs6XwE+cKg6kl1lGDGflgcCt
DIBIjk73dS9S1bfZg0kQjMzxejPJCRNKbEY+5jiuSSKGheY1I6cV2wBWfGUq3cZ4
GVlO8doPazJ2RkhoZw+SbxWhufIcLw889zDKysSX9Maqx52DJ3e5zviWy7R6vG0K
8uXq3i1u7ZhteLCuYWYD82a7Zs7J+SP6N7wRv6ztokPY9uo5Xv+PmgPUfjkcyd5X
iyVb6nbzig2SRM0ImTr1mEgET/rHLAQd/6qF3LMVGUcdNvsKM6SoxDfwzUu1YHXY
q+sfxWHX8poktkgjF+qYi/nt8NkuwuUW4Jgrf4YtE5+AF4/p/cEiNIp2H0VCy+69
AVzE2wBFmUIDjp/eNyGrw2F89XqNmdiExd9KfSuYhuF9qq6U5UnT6dX3EnKNx+EQ
upl/R4FYL8FOOxKBN9GYu7vHh1UtgnAX2ZpmlW3J4/H53PKMKj8mUp42rbK+Cehw
tkddBHFJuFqW6xpDoSVoRZYVKiR/UXcq2RqxVqvKYDqegO0yJrzLeAkZvh5Z/Z7I
uzWCxW5yi7ju5YRGhFzQvz5vg0Q2XZPdzLI+Z8CR1OrbDwNtMgXIRWglKlv4iu1I
NT9OiddAzLbMrekX12lpiPPj10ojdiu3UNNFNAzgdFcIxP8seeLTqMhm642VglQt
6FAY0Itxxdm0HShjlCV1RiLWkwB8EFDiydT6xKnX54VDz3Wv2Yrt+8HlEgc8K6cP
V3JpGcDX9KwLZg8jQfnoF1311JsNiYe+n2CS+DbAa/59aNXKZJvzoJcYfqk/Zjob
RGmIOXNpkfA4fjnmm8dtkR3aZNsdf4s6mJCSfVPC0ixUpZonYSTPtc44oJLfAMCd
eG18W0EunIQYt/hrn+1wmUb05HT1vzZcXKgBicdcd/fi70a+baE0DKnzNPV9TN/G
gMhp50vGBbp2UwzBYs9zZzGS+SaMIPqJBRo3TtPZHNY0Pw8meNL/XDP7MXh15y6f
4WL5ksnMJsXz8grF5zIVQXYcKKk1+9sP23tamL/UaussdPj3HcJl8sYLy4dYSRHE
1hZMuCZrjfVaJBfknb2wJnXvyF9Gfjd887qHrxrB+PqId9+gJ/Mm27PfIfNmb0QM
rXSwLopYDTPNnSvnQNRWnQqwX7xU95LSISFwgBUQhh1FhjWQ7YpDViKIk8YFQQRh
vNo05SL8J2tG/YuO85QjIyukpYulsmer1KB/ujNyyUu5Qjqb8nJKmbYbBfvW0ac+
GkoI07dJDTt4UzvkZYO49z4kTCVgaYWghcSk+Z+V1rnkCletnXKjqTSj8+ZR991e
OA71qT7nGbDqZbsN3lvssZBZsgm9KjuG8lr/zhaK6e9N8pJggCv5jt5hRPQlAiGz
Lmc3IulgRkBoN8+KQV+XIQPfH1ixQm9nmUkEHuhe4hhPj0644Z3AZ1nRmSusrZqD
6VuWSnc8OJraRDpY7cRDgOV/0DeUXCH1smkOvAuPILRx6AUY1vFf2QRVGBd0s+cJ
/TGLg1acb19fWy/+nfxDzt05fIYgp7AraGmgVITuJOD3TTxjnr9pViUsvyKC3RxF
oba0RxOoqCuitc9GoOuV/m9LTz1u5jEVXk74G+CU9OnZXwwiIQuNxtVBr82rOtd4
xAxuEdIP+gOQULNpuOhDd3uxuTJf4a83dPmVwcd2ogY=
`protect END_PROTECTED
