`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5AIZXFqImP/cZ3cxOo8u4XDK66SbwOKE/Y9pm0mACxF+xeXXQQZ222CLqWM9Py+w
J8ef75MBthMbYlGDq899vu8ep2xzLgz8ghr12GgsPiU8ZQ1pYAID70Bi06gknAZi
+QXE/I5RJg+IZckpVGIbsaiXjX0v4pE3mdf/1NqJP9fgBH3jxvCfcfdY6Rkpz/K0
u8Phachz3BQisXyF+QjKCBQj4xzPv59R85IrJvU8q6iYvrnX03LrBwe/7EPFifiB
aHuoHN/HDru4n1UpFzqeA0qx2aPaD5WnkBPMpZRAjFJ9BV9IOwrDn5YKY2RobTGU
+abNI2jzIbHA7tA5tQpEbrom9H+nDWw4ON7MWZX83+uDZTAJgpuGOCrWpiay13Ti
NfWi0EMTSGuxr77OepDx8jGixNHNDw8IRAz1oZU3g+GqFeEsGelm2Jt4Tg+N4tSG
lksMobq6ZwzSGBEE/yx2tyt8XQ7OfbXLq5hT7CEkeZItvZmASytuVTJwD8BJTD3k
Pa47KeTolVYGtrP9O8KqxLaVbpZRPBPdyh9wFpFqxcnKbfaQ3THLC4JVOErgxvmo
0ZBhWv91aIUAIIWAbLcEatsvy+8iJMEq+Lu8zSDVEeLNCdvszcuJtLVXSD57m6Th
bXW7CeGgBfp3yzG9kfbYmsmA2Oaa9wbORzYqU5Wm96K+dZ9Tq7RH1RESvrpM2B/T
EtV8g0XmQ5x8qQYkbXJLrwWS+/VGbsJQOmp5jHY6OWox+G7R6PRGX0w3akNBrGXc
OVRHVka2NHHEB7H6Ev+zv1z0IwGC3Tf8Hd4mlVUil8jZZ+YawosWpLRi230lhLka
tbCmOZPMjeKEl4cG6bzwfxMGWWmxMLfSuxciHS9JSnhamnROqp17zPuHRcKxE6HS
g6D+UhwswNqr4WlcFgNFxyLrtKFq3E5AoNqE2NXCF9c5FaK9JPOcCJl2OP4H0yjN
jfm3kXpzAo3p4ijX1HF2Srmbs8FlED424DjgUG8lSqeVldzvwJ0p+S9UsttiQnXt
KgVnMozvX4GmgfDqbLFKt9zBPWEVuUfuCLKGrnC6JfGG++WyP7LW9wtDw25uUfO/
1FaUk60JmH03pbasq5aqzk72xghhnxwa4Na7cahrsOwrPw/dG8r2UjUQuhhxRqS7
JkLStud+NJwoK2vYGaFuUmxLc+27l8b1uEsNVHISTM6AmE+MmQfU3nJdvcOArNk2
JETVPSPIswYQzJjlEsHCWkzeCkn+fXtWOjxK57yEzOQhJXe2A5Lo0bXJs86K+HXa
w9OQGRPJtEx7M8xsjMB174rvQJPzqi/dy9DaU3JZha4sFpShylYqvFrjLdApeYm1
oOdpnBsAYKRGG8wXv/MhXTLoibPkq5bB5WFGDC/E4RM0YKhAvz/4iPh6vMwrA/lN
JqP5634l1Uz2ra+j/edXYQjcxMkuNeB8CV696JnwUicCBihVA6pFW+Kl4/Ozcpuu
iUJaRfZJwGwQPCRXU6jkMzYm4ISUkSaDR3CwaZXJqrieYp61AIX2bQvMsjus4NEP
EmVpBMAai32jo/9X5Pelrl/MuDeELzHKmbLP1rRRPpLq6ug3dxY+YCboCxRDzspR
Fc9tzJYDMjDDgwKttcHj58iC6BBB8C0cCkhYiYEcGVVAVWOtNLHLwZrxPIBTkjGE
CZ+3cr2xZm103pOxpjdL9a17DYgh+BoCO6NEB6HkJAYM2bgWPWB1CZjvspnTAHuX
31tlPtEoXLRU5igfm3dkpGIJtSeAQhj3I0UeQCMYzi/wu+ir3FFA/GvIY92ELdK5
I9yaciGrDfdFHQO6gWAg1slEjO8Y0CGYxn0gMQm2yFd25ZAzC4sayNkUBoyXkWeD
c5AGCLf6S/dO4W6CeI7/xSkDVx5Y31/gRKWTP2BYETM/mfrpRaJ9KPkGtdvI47Cz
Uzlj0EMbcXlUAE/xRoz5Nn/sL7Z+DoOhgvZi0p9gO0Fz0KGsPWK9g7KRpFfg9oeB
DZIlZRGNvZY+t4IwU5VozZc1ZRp4J0gVcHXCDl85aaEUmpLo7FkItH0jKepv47u8
0rmqJrwX2Jzd8IoDx+wb53DjVusq5Fr8hB2XJH2pO5rh6UBmEe8y0rTgL80qUi4e
p2xQTp7PTifeehHSzlOPh+ZtysIdRRzlambgvRnewo4a7rT/G7sapzwTimFByXc1
mfYUh21gHuzx3XyQySprB2D/yLQzqVGhbeo3QTqRu8140xbUjb4CuVuKbZJtdB4g
C1wF4nGWYi7KtXBap8cIEJVJfIRhGw3W0Z7WTrGTf3hHY9p1MQ4LIZ8pYR30Hjqv
lvp7N5I+kpcqGbzaUSkXYTb1MSYwPreBd2cUMqt7MB9ANIYUHrJy594Rnwkx0Mv6
dWUfIfWbDcRn8gD0TtPf7w==
`protect END_PROTECTED
