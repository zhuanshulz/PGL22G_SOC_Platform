`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pNeBJd06Gjp8d8Y/j0iaCYdPlxmdwJXdl0Xtyp1SFa5uAg/pW1B/PXVi1BPN+n5D
REWfQyf8D0HV1FLLGsXQSj8duyhfH6Jm/FQ8QeYj0CI3Wwzve06qh3e9ZGEsd0uo
DYZihCqo8vQbsCI3IscHHil26lCaFD2eKLDW2QFdTPJ2OFEcRs9ytBrGxLno+ZaI
5hqkbV8bgz2IUL3OYLT/XnJ1nW8gZ5Gc/ORgRLN4naPyWAip3Ru24mgzt7biJH4W
zmrJySRW0COCa9uG0SgVgX9YMd38e6b+IoS6GPaDcjybsflW6WsnhJydt9CuSXcD
kvIQ8E1ha6AUcTRPqme9RFnxE/7KN57nEDvS/ULX8wFPAsE4jUsx1zIaqmovjoph
+pZuRD96QRMZp7mLGTM85KJXIXCdJlnBniH6mffdx+fR1KIxYMy9R4Low0kn68CT
V8BWH5hZNLEXd+l8AxxqjDNZmB82JIy+ddmflYjhy7ui5eR3wQHuJEdtJumCRtWj
62ezrQIuWVrnmD7qJSr6xB/RxTnkHzwfZ/IbMHsrwS1sjItp5Wn5g66s7FTyz1cQ
cb/0xaJmc5Zhi421GjLaXl8hwPIRsF1FN9X0axzmN8LoUDJ1rXkcRzk/roZSHvfH
sXsz/THc7TSLOChttdZB5KIJoD5WBlXjve7HsCcpAzO9mdhXiCEOSIRU2DFNeUPf
7eYykoX9Fs+Di4DzIiKNqdODAz7bI2IDzcCD93x7xK1H2YPGKR1sjMfhZdQyMc+P
Aomu+l/Hv1+yePh3WpCyBoZ38RvbDTlhGs6gOws/3hX+mS6wp1wWPbyEzktXdU5y
C3etUtVKZ6lgis5IkYPI8k7MvvoOsiEFgMOBl61EgDIcfR/8IlcNI4gzRQj8mJPh
2xrUJeZ938A3iuzzbKTWnFukLqpJ+1mMmyuLw5IhpXWol2LWQ+GMeZoGvfUDF2dU
rTRupmprj9YyUo2/JB1OFzRTJk78ZaBXjvd0g79SYlKRAQLelaGaguIi3YjCf42m
sOj2QIoY4eBPA4evkd0X9R7yTaAWJ74gkLzwCHJ/QWu5R/VxhaNrACTOKKBVbKlu
jUeLNbON6TWGidzUoiEuNb1Vw6S4b+BeUoESrEGh4EHJHyGa6w0qcsmo7mE8SPzq
NIyDU2uCelgmsy+GF/IlVDsNuL3WrDvblOB+c68WjsfAufS6yivV+oMKRBvyX3fB
kUAezRwI3Nz96UC8psMPONAUgWn6wGbr5cc4MdftIR71y26k+p++7Fyxur02a7G5
TfKRcCiSct3fHnFoyWjz/+LGuZWIHu6VptufpBx0RQnraY9wlgP4ovGziMG2Lwkj
SLJSEWnm+DoSuq0Rk5aHBnNwaIcfmVjWoC4BWWJRqXJjll121dAjuzJlRUhBmdMG
5AcEDVU/JrsvYsNH12ZcyU7uWbQiRQo30GelclSK2cyGL59+Wf6UpX+gzW56EX1v
AWnreC4ms17Mvoyx3GrNxwBbeYyPaluDN7C9+Zrm+PXDeh8wkCVpW4nPEcP89FfM
NWFATU4u1VFlTKlI5XpHiYOKdEVKJksqVRuttuphvKm3D7T+Av7U7NUCcHwavuZt
a+xdwxEImwP00XigpREzEgzKdCUztzsGdZGdNmcpb9vahic0jLZeaCGSWY89hFoW
I7nt0jdPYXS6aY/r7F0BhpasDdphx2LCWTaOGqU9ZdT73JQSbqC2uRWF9mJnv1iP
BdgOZa+2JDGQj+2u66Kmm/nIpWCtqhzyUVnw0UyE1JGIscZ/tIA3PbYb9bfFBlfq
7mGcmIgk0xUa9lhvXrTWJs4InwefWhuR+HE19rdQ0C4aV5Li+B4agFk73/iImOLA
gLGLHt/ITnUxn0Je9rhrjVEhdTDku/ObHIZS+z778HJDz5LRIvwRfWeIVvWqrtA/
w2TDaC9j7rbJRe27aG6vhkaiYwj/qTL56jrj+IAinvGMhCtlWAO7spSQKoX938ja
twjOUVAqv9HL7IYQZuQLKxQV/UB/s3lJ4O6gHBot3dtYzFJhlhEu4eLdWpGPAxNY
hGvd6DkoKLmPafGQ57Kg+RFLHYgIPbknj8K7Ue6P9k/NwwuS6sc3zVz/+YVSlS6A
OMikCJ/0scmSLwoqPk3TdQ7cpV+EStIRgGS5fFIrOYXVxT6O8REBOikW/qgFquVi
jmcQXfGkgIJlvQr9H7dw5k4rWe0qn6WmQVqgg2nyiKPiJUyfpQ2GocVezZy+BgT5
F4pxmcvpLscYyQDXeizL+NRdzneflwgYXZlkXMwBXXRatl6cHbXRl+tcf8IRnRLS
fmZIxv4D2iCuaTKoYV/kmjhaPnLkQbgjZMNb2jShsSc=
`protect END_PROTECTED
