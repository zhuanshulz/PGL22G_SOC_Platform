`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RESQi1uw+sMqkcQV7NGhVfXLvXoNrmh2Q1M2UZ3kRm6ZiMFnifFFVyrA15p9VY0Q
tBmHE8V0NU0K9qcUTc0TzNgJ3basoJ1Esxo7w5OenHiih2iWMpCsao6HGnWkEDWG
hlHQKl2nHpHSpfU/A0wLdXCaQOV4ers3h/5iYWt1DIKa6Fz1+Z4fw2GUvNSq5OCY
2FpHyoKlvnRRhm6RRzMH6N6R+Vuw9MxE1TQfaXTKLAnsXDyxVWwUJDVpE9crLxGG
Wpy0MVsC1BC/R9B4sOVRD2lJ96jZdkCEy8XSBUDRkrt1paTVXeExOs9CR2MGfVf9
PYFHwbVegrmfqN9Ea33G5vn8cO/ugkDy5P3dPFYVEtm/si//Bd38lxGZ31kqlIlD
mO0qKDz5EwitcpOYVnfDJl0ory/wcm0tq8TeG/fdLF73TesfvYZyO0Km/X2qoBAv
WLYvFOeVmjwnnb368vqbf/2liY/DKOVAH8Ji1oKqL40vxzxENczOgCVU4rb0cGo8
cGjDdJiTdNEdbAWHyDVvxGDg/RhjTPbtTWz4+pCjoZ5Z1lgplkX4olt9/X2eTnkP
08NpT+vf0SYGaJIHfHXofdgU+f7zT7u+cHy6r3aWdI5fGbeDxoYFBmVIhpgCjH2T
QYVWGV17ORt46I9Y9eThBtUU51M7IjngAHzLqhsEjbp1m/qvzaRDmDjD6rqMQubY
`protect END_PROTECTED
