`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q+MUHkQiReKRot6B5+BmGNpWY99cTE9Ix8kR66sCsEOCP85ifNgPXTXRgtumOFtB
GEKHMrM7GBjHcWao/pdaUoqD0uHwW+ypKJllS+zR8ARQtiNBIaVoripdTcBuiA6R
9aBv4s+Toiqfh69AeANCYN5UFTY6mEv3uZt9bRjhzYd1isdMnESc3seMmTntfRN4
E+eHBk/enZ/OGEx6wItmEbnXF/ap9Pd7eBSvkdTl8mt0hpIAuYMb7EsjitUjLJMM
MKfXC4knDwuoZmpJgwmSaNf+7UxyvzBguIn+HifY/0+HMQCcJ/ZbnVn8UCeQqzk4
r/TzHN4LyQIs5QcsDNTN2ruiPthgaeg394YQ/tdEA6ECsam0ZgYXtoq5iEryo2Bw
Ut/pZmXLQDG0Taui1eY7UM26TGzGte/j5BQozLNEiFxSDZJQoPiPlDn92Eo57DYC
ATJKSIVUSvwebBaEy1z7Hjve2dXRP3/IC+U8MRRe058qhBBQxZjYQuFc/bjAVoqp
KVhiGry8Fl2tnqFt5AC6b2Vfyg98fgoTy1xguluAEjsiDr5JnfgOwfge5HXVh07x
Mqm/irlLjMneZ3Nm3Q4iETKRk5n1AZvciCZAcOXpcj4oCMeLaoGLoqjWmBCHwNe7
EHC9WZFqXN/AC0nIY4P7klN5t6a3+KhMvDVF/rtDBiwxZ6S7YsqOmme6ZR4ULLhY
ySiqp5apRABa8FftfOXJBD3SX96ShuDrBpS+Wch8vsWRXYY5mpLYxKa6jPClfg7B
Ax42xqAaqLK3upjDMwncBaxV9TKOzEMSf7S8bg8DbTguC5oWOvEllpajUYALa3TP
N24z/UYVwdF4ABzsZoKboQiu6hJ2RdfNV/hk9bywOLkY2AE7Jve69AOMoBGVWcw6
56Tf7FsMQl0NhxLgkJmn6lwcJK3GP/SiOUVYre/hqurUdgaCu4JVaOWjtqtFp6zu
v8g4Jyv/QLOVZaz6ixWlr41WI6bTypBVfNRb4Aq9wfgr1a+N8ndmvdKhrMyViEE5
cuOySZa2BU62zACWensABMk46NWtGw3JMyl36R1oTK/f9lfvURVR6m4cqas1PlN3
RzxDEG+jt0eQdRjxlzALtKZCtpKpg3DKWbmU/r9aX4WYvapEC9S1fTKoWJmVtNAJ
alB4G7XdJmRv3Ohh6qFiBwzaY1pyI4JuJ8GNBDzigSOeP6u/edX2e8SWSVElGS5m
KK2MfAq0y9taBTyTXpk1cfGV5KfzZa8409c1lehSJC5llLGSyagib7lmeEq9ggWj
Z/JMgAq/SQrctvE5mYfUDZqszi0sMcSod2grQXKIgNgKXReU5KyE5nNVrpfokfM2
5oYOtgyqbAt0Af1tIaWCMig/GzDJwCLPGEFbTKY1lGaDcQ5P3B27DfEUhv2UazA3
5SIhf0qEzDKjIzI0lZbZ4aNOJ9pVfUkDF4ZnkVOtWtjy0RZMVn1ycyzzqb2cm77V
lNwHeBBTbvvv6J1acHrV+vCEtaJ+kiFNxP+xc9zE4TG/MrumN1+6d4ZZ+I094HMq
6+8HlZXbxgMA8JmZneb5z7TLkeGdBpKp0JS1NCyC/HqJs2BSYSRGJpcGdpB7TSZ2
35JnYlkFb7GA9KPPf/hJGclmOfaHU6qPp1XK7dt9T7Kof70kaq3J0F5yeUQpvNKn
uA1bH4mFitTPz0wbs3o8c/vOY/K2qukuobOAZJY1rYpBlXTmLUPzuWFaGEeBIkUm
dmbY4EH9dJnBuhWu1yKZjmBihXyW41Kx09MrXQr2zhmieiVPyqTAgTkM0ix+CoP9
x9a5592MStMIW08fuBk8Emdob84XUazqgpHr4+fIbSlk86ByIA342vaF9bRDMuJ7
V16qOxxZd78owlce4BZdVPWSnd71IuPBqg+1Ktyu2vDe0jWYaXwURfyEz6fgezGN
1T3nhg/2WxTnB4C9yTE8t8JooCaAL5Z4nVvvMDpD1wMwh1aFP+aNIFCR8lorAI5Z
2y1P3ihlAASIYjugmuCw4p/bD6CZFk3FhrE4QN8Ookcdf8+n1HdFajrUAOH5P8pS
vrVmKZa70TdYW3QuVVi0uloBqQNNNNvJEY0+VoAFt6LH9DP8X/B/axUv1M5K1n8M
Tg97sJPFTtxWUirjmU3DneMmYvl0sByTZ63iWx3R+wgxXxbRH64B2wUt2ULaEHCt
5rOKiuDC0ODNiDUOYPsailqVbhkQj85X4yuDKxP29EOhdZAzr+dVqNrK2OOr5YQ2
epgnsR5oJIZpNBEbfCcr3D3LyAMe6Qjtj3hsiOF9DCR9v9aKWLUlhXcoJBjBBt7C
DwnGpzMqOnfEQ22da0n/kEBmLqRkbiO7uF0o2pEytsWTvik0n6sVlIBzfHxMuqFj
zG5ADofpgjtWw+dIcfIfNvrOEzu1PGrLOAjoxR06ffg1Dxu9PgZiYg/BxfKQiv1i
39570pTLo2p8zDlMTyTeuCqKgE6tLGigHIPs23mZz3QcAKe36zFKZ9NSm+0JYTlD
QzlCPDDJEHDravIQqvOrlNHNwnXl1v+q2rCDAqeYvH7YSo88CJjzrVyChryjhMgR
XD8ef52nYDW5bWKWNizTUi1V049mXWWNVDG6OLNHYEzZ4w0oO8Z32btFjPw5okC2
vSTx4WexZ/gNBGda4AU27YM+qNy+bUTcraO9+5ts+rPiXCR7G1IusGD9Lzd1zv18
Udg6HVJqM3y9DlLdiF+AmOGV2bvz+Ibohbyyj4j2Om3eHT0/CSD0j6yU4Kud0lQf
kljdMCg/TLJwfDE1n95DWciGAQOdt8Gmem1sBFCahKhKRAbDhxCuiYTmp653Ayxj
kDatItVLOr/5GUuOWL5Jl4OgJMb9o+6FrW3hN6dFw4VYMG9bRVC1N9eKI4kQDBUI
tGyPaW9YYQGkCEt7ZUKshQvk18ZcRolhv4OJceRXNSdRUsL981hEvmTLKIA7sBJl
Uk4rpi+EmRJaJbo19OrJ2tU4GftFUtLlhSLw8rISSLoa3hu+rSIrmAi27dX9nbp9
qAP4nhmckCeQuKYD5yeEmKiB+5+Zf1+hpE1vap5OVIgAAaq8rf0GPr+DCF3scbwl
MSyHeSkWFooP7uQDOSNSMIHMTRVmFWhVg39JVSpi8YxEBtiRMaUuScC97+2thXJJ
EY9zk8C5C8O28Vtv3w3TWXM2nIrghZNLrV0MEGBc7Fy6KMLS2dCrvuS4JS0pa0+i
aEoFdyjW7K8Iv69o61FA6mOqBkd4Q941UOmzXISiGtpcP2CfXfAEcNr8avotJgPs
eJBXwnyYAYKrIZj8X4FC2DxE9CUdBfOnCGN1bsGqdOY5x6RMfWhqoUu8WNYtql0s
N8ZZullBs6C/F2vcDz2hDUzd1A/qsAkYwX1D7u10Fym5+x78Hj6QLjVLxA7EZmgc
paXlh3rejgG14Sut8KDFi8PeD2bzFvFaI9YQDL24HAbcBcuGhrFaSS3/byGLujTL
RQHVrnI4Qk303L4wK+xg6+16t3R3EmQzUan3fqEq3HX8oZ2jps0JInqpbczf9hNS
L0WLCFEFJ1RKL3tmbr5/LG5aS+LhVhJQKypl1N2RQKThJqxOvkmJ1DUA0knPskbs
1dGgvNhuFrqVXeufzy9usOnmbq1+nNYJnGR9k3gjcMXTDmZNYoVU8kPEl+b2cU68
uX99mAWO3YdFSX6INL29roeOJQB4rI92GS9rPwLmoUwLGY1t5XBcZ+lE995XSPX2
RE80BUDJ1K+T8cajFTqPyxk3tfCBtxfwsGuLoqttcl5gG1+PV06RdEoqHXp7TTeb
kWhu1f4dB/YgqNAcv/K1aFaItb/tkd9QsoYq1abKRbIdQscT8YfLN2+C7LXY0etr
/DFtdjzL+5xDAiry1I0XDrdh4yHvpJwxbJTd1eVUdTIp9tadThWDAMD0xp7SuoTU
Md1py7vl5ZxhoZHRc7DFxEse1Whv/F8lXJKMqhf1Qtf5bQiehDumfXXEEPfe1dL7
kZkAjFllrx/INajq8wDcQit/VcKu60EBOzxz3hHOCDyUg33ZEof3pmGsxI/JnUF5
YkgNLXbVb3sZ4WVKWk28gesl35N+G1VadO0quPyz6D1SF0Dye64jvbxye7S3Acgg
N+sFLo1eUey0KJKZi58pyzizY0luIDbKmSPKRPe6tsOFiRmVuf8TX3p2k8xI/xPq
cx5A6GYje8zXYzVkQeUTrUUxEA+gWtNnh9KycZH1qKfRvIt+KVP77rJY3v4JC+TV
9uyoC6CCOGktvNPQ4/7fXzoQ3kHpFrs4NRXgTiUCK6KBN160xSrjXcO2iH5P4yrM
mMNff2tiNsYuns9q0vjC+akM2qprpSebPuOkOYVMvX7ONzqcGw8hDWCwW+nbECm7
/eJFqATjVbLTNnU3YV3BePKDGvOzILuuivz8TFv12sZnmIaIp9m/Y8ZNmJYAKZh9
sEfti2PeBL5r3hPD9vJ3S/WFlvU6KKYfc108NnYuBga2rgQa+2iEvlZQXtUyhUJH
cKmt7VyiZy4+ULx/1tvQje9/RwNjbgaTr/lTI7bWe+ctdGUJoL4ZzXZ9/dKD7mlx
aBa2I11Rya4M7zYGGmzmSqZh6OWQHydRSv8idKHky2ee1mh4gETQN25QlCrHuPFB
jO2kIU46Et3Apug6xAxOeSuQ/8yzFZ8hz/W+SogmXYkKCoJK16PGrbyEDGHTowtc
xsFBczKz+MMVBw6hLGgpRexj6z53AYAdIKC+XJR5uE5owMOyF2eoYcD/mhAL2omd
kntyrAHVGxq3B6YQgc2kk3rcE6wyro5rErO+EfsFhUKJwOJZWWj6ovtnwy8hooNQ
X1nslMG+FiBAlkDbMRtjehsflBBJA/ZwSzh+hpiJ3iwhnwJdvXuCnyrYluuEF5iR
qln7U1CmE+IVCDOe61EmrhhDzoeO5BSyxTqHJM0x3Vngs/zwsBueK3oeyon+f4Yu
ErBT8i72xKnS9Fapoy6MK6vwsrfAmgJfGaqPQVby3+4yrjSLYhZKG3K3IwQ8VGbi
MlqDr6JpUHN/2s4h38UMpK9ltRNMgu+xKEsgVuzj6qSBSzKBbZ3C8txYSFHUqqB6
U9raxArjvedz+2l0SyNCI4Ghj0qAO+bDt/isnAz27rJBV8YdrkbjnegdkWLfA/Ea
BVwKdjdeuKBwIclegQeaxdJNJjB5ENzkVGuVWqka3JRY/Z7Zoq928d5Kh3zkGD7E
ak9bdHRfvz8DI39Ji0bS9PbZnsASFfMC5Z1iFkhWH8uuz8XZojBkKH/jX4ZrA7V3
2B5nuX45/Fym56yEASGaF2RfYMFm+6yRaDbBt54M6PtdT/elNR4T4SZnAmJmkFrj
XPlQQwMmXqbZbqlqRYl0iCp317GlvgKvqWfBomWaD0P+wPONk1sCyVP1i4kH7TfW
LOrGN08dC6lyYJHZAZj0Pyh8LAmpDN88p/PdTgZ95g85iMyh4jqIYGsw59Fyn+zn
CQFSClHeAFhRzw+yPtFpsdqXM+lKb+MaW+vsRL4Nta9lvqnPPKCe/IF7HtXCstRh
TuxunUl6AENFQi8Y4HBugfVFtfghGi5Fkru3ZO8bCG3mjaeXQdG2yn01HIg3N1ea
PCxchz+hu1GdRkHnE54jmqjxgmGKTNjRv2d61h7qFsPxgJEXekN4Z/JnbQI7ZcYx
ebUVnCSIvPpmK8iRP93lTgzKCuDcwU1bzoKaauItumK/vMV/cmcNaRrNUxTe0Rc4
mTwj3aIoh/btx9ItZwdWIc5puZr51Fb3U0TtaG0JBu4eT8Vw76CW2WEA3cKM1/4r
3aHBhvN9o3gsh5FxYb52xH/OP/CnF6sNSgo2BY5mOAk+vSSegqXv3bmIskiC4Bkv
LwFK9DUSBwYam3UJYj0G7cQmYKTiRCscF7OWTJoI7jq73g7AYmuNMxbBB9LlR+Go
7a3ZzWNLHZbDT6/ornwsC4bZfRO8gzykX3TZOe5+X7GLgeYIThgE4WM7xMCz/PQc
Wr+zUdBIlZzUqG7BZzMHu7s/WKTqoOh4m6DoUKF6QZZpo/XX10BLFNzOJTzyZmKR
Q80I3WmfCmZorPk8U4AK26aSWqVu75mFBmutBjEwLBakgzqcWimDBy6NXy/rYbhn
q3VW1xftf221oB0xrGinU6mVcnuFabyDX3V3xJFHqQMwG/W5SXcOS/Hzj5oa4Azd
+R24AjM4UrD4R9BJ/fN0cAMRc3F6+ubXnWWCM5/YEglSyd9CRXLyLdGU2zcz6Xfg
R46sT+86k0dhvEyfoAn1hVvQsrWAh8v7HxQxZ9onU7hCsx/bursVVmuPwYvahHwa
UcKbDdzv+2jgmUii2Nw033CFk4rq2DVkDpGQFY553FHAlBbFMLfBKCVNk2rIlpst
tGOyp81fRKpPrcVDoP9YO9iBRYlqb4wgsbg51c6y1bPeqnmCfc+D5e/7dYq4MXdp
FS0813SUpVxhQnjnMdzloUIjQ7O5c447MeGmdR7aV+NVCoYe1WwiIkA/3lP70HSm
3guRp8LrXhNpxZ9zCMru93TXv8Iem9xrlwYYpvJQBI2zUT5t254d5GSw1Z6KPLsg
uzyrE1rLpF6CHIp5a6e463K3EWXxpJOWoTOg/3jX/nIWqOGwQdlGIqCXTAYGc7jB
ME94mLuziVE2bUnhtMNLT3YzWWfQsKw7yZHg5V/5GlIdC1TeXxg2Xx58OcadEJFD
dunt6o/Wz8pyGx8+RgeBYQeEIN16dw3/p+n2DwBXKlfxvg1JJhjXnucZ4iPA9Fih
VEMNYRowA2SeFhAOP4LIXYt/xvQeg6vlI9QDTS8HTfC1QOuWX8qD2WrmWL1gMkXu
s/OKjGQH3ddPIqXGr8mYSLgJ5BiC5WVQEHAPv+2HawWCMqxeRxSdKlvDlDoHwvHj
TQQ4eiaq1fYNUaBT8Ia4memazCKCnVhj//7SY5NLR8AM7LdOjvXpfFV0BwIOLR6n
F5lYG4VT//DwDM4L630ItI/5YRiK6mvLir/rRbvrwNRs3YTaGdt67zmq8p1hNkqD
QcNddnlYJPaI/EqhHKAz5dOrGL3sOYkwjkYiBfKU8+X/3oRu6ExLCv5A1tmXiZdS
alGmujXB0c2cic+Mqfn4r8PAcAmMYVRIPd1o/JSIlURJSFyYbepmChDxl5DGy6OQ
Vyp8XlbR5ffagsezXcbjbB9PpNsWAbFodBwBreslzCydFnzyANGFSNuOh5cquPjo
QdkDSsiv98ECA8QHlgj4OzdyJy2tfpoTqEGWZzsSypcdXDlNl7fvVx8YByYU1tRc
QjNtI3u9saeIfPwPOftMDEkpClQydYI8BHoO0n+noHX3EUbV/VA4V+TGnKuqWNYa
RsXUccX5KLf86bZGtrpNwAN15/SakVF39FAs5+iQ7aZY28INXIp/3ojFN1owU9Jz
LQe0g8iW0y9bY2yhsfCOipwIjSW+FlRlO9CcFwBO9wH3uvzLyjFNICC1fa4I7NL7
9OkyeIS5sc1zxv+fjm+UKVOs9+mb/j0Y3AzSFOERX/78Z30FwHubCh3BYeShSyOJ
uiK1M/4abrH1JR81fNjXtZJpEhNFbzM60L25UNcBAW2KByCEh2bkjppkV4Bx5ZDs
/FvyVyvX9PputgjQ6OnAfQVRkh3zHxbgwsmgAKRGxCyEzfrpcJscAXviqJL+aVBo
rFpmWPXWBL7690wP7iA50G09ELVFXgdgee3a0jKf9C9If/ey8Ev1DCxJ97iZZk7Q
wxHzn02KAHPfqTYHCmtMZhTQuiWWywRBHTaZJQj6c7cT33dv669LkycEa+E9mp23
6iXr5h8SGJyXc7P/mGs+ineaLmHkAgayq4Ba5hCSWyWKdbAE8JJVm0fZbnqe8NWc
GkdmqyH3QCLQ8ugHv2YEzwsxFEIb89wn7U+dVzJ1Rp4OkLdpONoadWIFkyY+m+EC
Svaaw5MhBvGE8BaKmtYsga/H/yYxC/rGIA4StI40zQ0NMz4Vql6R+GVY+bOsYvUP
oxeqkccBBoDs4fhlHoIo3ggp9VsqBQxr2Ifvt/U/cgb6at3kakMYCInN+O60Ijk8
jz9hSoVr6CN/MAwOfD7/U6M7kqhnn+sEvIvV9ZrrDgxvQjn7qB1VKeQearJjuN8C
OqyoUVmfxiRm+e9QGpn9xgZg8NU/RUmNUnWJ3Zh9GLfSE4Z0Tmo4oISqH0GbSQKF
m1CGj0ZAQLeb4ihX7Kob5Fp9uZA0KKZlh9+wnryRKY1f6u9AtENEyWEkthCTCNjM
/F+l2uJoLqtKdWbrT0/r+QCcuWoLeGGAvb/pZ1WzZDz5XzqX6y92x5dNdRqa2L7x
pd74a/sTH77qIAWkDl0cs57Ao8jlgBoSxaSAp5nNb8FKcR0YkKhZeTB3VyKDv2uy
QPXKNPW+fU6xB8iOsN5QdQ6/P6MqfSWVn2lge0VF8Aw0izN4oz61wGHAM4j10JFT
jYkDTHnM6cUYjP7RG4TEJcCwNd/hZZP1eHFKko8dJfeU514TC9TYtORYI/UKxhr0
NTxQp7NsX03D4wjXL3bHy4AfO+C/VZ7zU1TSQSFfM3UFjzu/OMDeWvRGO3YJtzkc
s6XOXJjcgrpH9hIhRIjstCGZ3/8E1Tyu9HHBoBZNZN03YZv1iE+HDgqTwLyuYIsb
4Z/tvyzcrEZMficHsFLfhr2ESs6AypDa/vJ70dKOrog2Vtn1y+W7Zi3UNHlJ3GKu
YqLmiDNQi82/mcONjH+WDk37e+v1xIB1U0/M7Nchu6PlbjDdng7o8GVsisqJS69w
Ka6x1Sx7LB5Pg6Sx9oL8Oc7OHLRlSBndwK8L1pGHKIFhShYEFIIyRBXWgfX+T1df
Z0Mwf+0rrpafbz8or8psNoQtggXvYLcHP6vrspvVFIqhDyoC/r8F2uMFo51lsS0q
hVxzaw/6iScT5Ui03rRgs3/7TjEOSPkrjFWW15L5+hCtyfdIaDjhu5ZVA7hhjfK7
1uKE6ck+jpOt6mljmq9lGOzakE16Y2M0wHpWQwF4bKLg/D600k6alWn+soUn2LmP
XIfiBje7k0xAAhUxVJSIYb23X1H4Hr/Yk3wn6lmKEF59xGMArdhAXUyfxE0pBKpg
ozUhMXfaZmIUir6hgRFWF2WvVfF6OJnkGAYqAnUe6yMBHqn0li22uN6dX8Cj1awa
C1i2MXa9gDKBAUVV+S9OWiY3EIEvb+ygi7NWJYWXXedPJpRvVVn0rEN1Gq1VU27/
9cUNg8FoZyfpmS2givCxULitU0QsJmNyzxkDJ1m3JSxaSJUlLVwuWZjfxBkpqbbE
VSPz/F9t6jTOvrDf2OBfkKKRXYWMmf5aTif3PFkXWnJsXeDihqTSXDpJvxcffRTd
ERZaKC7PaUXuM2N7Ocr1FlJIqWc47ho/665kzmHTwUf8S5TuZ3kfikr1rW4sdxwF
rn7Ky8DQ8CJUhVvZSZP7HrICK7NbsC80wiU+BW0p5X2m2Q2EQXmjxcl8ZuwGS3sv
0RN9q1DwTxsWb0WJfkrHhs2VJj6iD49d2jTlsn/OmYdhB2xz2AJsYlhajY7Z2jv5
qQZ3l3ECQlVWjWsu99wCLXfpbMXsq3OhQdjpWxqWhVZVcAN8po4nDs+CVIA7tyOX
I9SGOTDb0DLf40hanF0IdiCitrzDuJi0Bk5zhShIO+i3yv2jiJ2qGXJoFnC6dLhI
dfvOg5D4Xh3I+ahd/BwblL9x7ttuQkTp86saxUkmogTz+a+Ik+J5nQXxdjGpXMv7
95g1pV/IfeEt5FzVO6anQtP0/WHBk8yMjcgkqlSzVr1Cluhke0bQyN5h08GeNkjv
z/yEbDYwLLLidjVvnGOlBr4jnjGvVcf8zUGHeqRtjFw91b/2I5kSBLkUx6Fgb67l
gOh0XgbWgjjkleFAblz9yGz13224kMoX9Bgi0atlh+CMt8odrVO8F99Piy9zGH1k
JINyXYuak7yKSfIjvz0leh28rrNDWD7/OUXX88M3A0J5jHyLCABOaPuehhJy58uN
2D2IgIvnB51zbwqwgqtzFGVBWCmToNw/F/M8fQ+XB7c68i9LydUxc+sgWM6Dti/C
NQTiXXUrsuywe4qS+slt+wk8FoTLg7/nNkGAXoFDS6S4fFba+7LzSehLLw1KGM4u
rGpEpvGLppaIsI/DYGLN0B/O1Lftdnt2LwmJpOOEYZtF7vZ9les2FSYpJjq6Q2+X
LP3RSv0J2RYgSAksTFlrz6OW5hf2sBRXgRem4Rdzvmc2OgEkEWUDOmJjsKhXhS2K
EzjzKlTiHzD5wISSznhE7iI1u6rRMpXXv77PdGo6yAaMh2iGrm+xZYctOfbFhQu/
0ObaNK2Syp0ld87u5QVI3l++75wXrw9Wrqqp1xKpyX+UMEdWaKWQ2+06GvvTjkdt
676z6XpnMLWGR1MQh0xPLVD9fIL6uI0hslZJj+sWhW8T9PkUImCDhKjJaNSN2f/V
JchGsVKE6a9GkS/zLU56rURw6e23b/8j9sasn7BrGgOOPcISVgNcRiOAn3MK3Z3K
9Q3IndIjGwY4N0D3jvLPsIQmT5lNH82JWYt4sbHO8XCkNLlJU00Mj7Pq7/LgYx6B
fcgfWa1aahbcvcs0rEmipTqlvcDtMlmrbYcMn+KZqJGGZKTIGUlBIPA+Vq1YhABU
r4SmkQUGTBI8IbM/fFj7Nxh0lCUHUwJFzm3AqeaKhIdP+c7I0/JJ4JUEnhZO03LI
Tex8Zv0wxAQgRjt2iClenxdviervcFdAew13XxcJwOcA4j098PmELifHl4wS6bTZ
+Poynb6x6WYxVUPlOvzUidQlQr71ZM3xqGXaxfLUTbpuC9KQZVTafcctKvsmcnEN
5aWK2mYZukDux0vZ8l39Y4msvBXcu7qG1c5ylvHIsvXxz0K/+z+Esoj2rkdaZ0j+
DTma/Lbzm0Bh1GHTR2ePkSeqi3xbhyDNujHqvU0ZJXSqLVW1gHIdraPgSeb/ECEi
O+FtcTFVdMepWvT6s+BGCUE1avMI4HuMyPFQFY4P05lhxNbCkntM1E/Ga8VfTiuc
4FBaLmg/suhyq4lcyG5PoaYWNngAv5qiIXnsOTgtEotAg3Pc74MUUlKIe/cbzy9A
nbzmW33CQswr8dCMAy842qjYQLBpen+mKCZ3g1TjdfokB/faymfCuU1FAWRea+jn
Uq1sfHI4BnkfhlCRsZoHYs/h+BVAg3sAcCl5AZ40GWgOKdGlwsPdbALJH/Dg+ytd
exijkj9FQGm9+A28zbaFGan3XwFeXt4BT7yQ+xd3X/3nOdkVKQfFWodyBZlSxdKW
aOhFB6LRBeUqmGlbKzQlJ6ho3utRw/rbNYIDdmDdSp48wioB2ko4yRqIJIm+tlhx
3FEaZVhAXmJDXKhl/gg4MVEO4N8VvjWUIHLSvIPvnZYsAXrnvVkWsd2QmJzJG94C
a91p5hCnvxCE9Ce/oLvuan9LrCRklyBuaEQPIuT7HrzB4KeBmDiqJZzuNQ7xW/ds
Urp6Xu75nQfyWyKdeFeYhOyWuNLVWtRvNlBwmwhl2EFPrTmtNw7wz8jUZvpT/008
8B7WZ2JkrPHIrEecyHIpVfsbYd9VIU8gGowdfLmqbyqb48oj1ICogbMrq21l3ChL
SesuCnEGd9q8lSZcHIaOQa4EU+Aexe8nkj68v/XdxrLN2JqQrVR7AtCKlOZ7k/hY
CtCTizh8EFdp14s07ib73LblDLvKV2WgXPXIYXPQSiQN1tqQHtshbG9iFImjZ4xt
ag/p/U2AuzR3TFkdqwTAJEhrEYQdkQwbwmVIJHxPZD+pH0+zwNpq/OGAl8LQHqus
W1Yle2xIjLiI2QgwTioom+oWQNzSi24sFA2gw3rUuU5CvtIpNrpL6dWuh49daIi9
2j6p5cInEqEcY2HgfDEVg0HjMZrQ8Jln3t+R3GqpKwVFbYSeNwSqI5YbfZs6syeA
x258uzmozN0f/vyAWQvGBir8UhszWSnMkPXQm4UozQiVru7uBqe3Uunw++lIOqFF
Zdg1bGDKxuERECH0DM8qGzw/J62Sy0KUnA7UkY6kqYNMWlR/wNvaa2h0MCeBYAeJ
T+WuABDTP4hupugBHrZJfr0O2A0MDL4dYwKu/E3heKVQNdnZG+irNnxefqmtQGaE
RV4fuxHdwTBl+QHDhX2p7hhQ0berHz/LnBqc2lKcY8M5u4hypV5JNHU3tvnda8Fy
ih1Y0G43WqXeDwNIf3ugfYDyx4o/5c2+5M+4ylus9TVxXBEdfuVkVrt2EwZaNvzh
6ephs6188bPxFHZ5DuNOENIruyl29O8yBiX5Dc8aZu+SogQWRFNW5kh1EFe2nO7R
BjfRgXxB2/4AM9Lg6DZsnq31viTJyrzrbjaJEy4gdM1mCU98ScIBXcxwjnMDNRdr
PwDZkB6MWVwWI19+DQ67vybHtBAD0ZS1/oNuiPWZJNXTVEz+4VrU9u2MFoQkSimb
w0zTLyV2KstE6cdQRgUrowo/PeKE+pmYKYGxxfwSMZbpYfs+61aBHlHrjbxMng70
6jCQr2cGCl603ScyWBN92ckZ8XKVmBr3BE1VxWAXV9drXQuR9tFKMap6imVX2Bzv
TG8MqQkTvIeMa4nTkAQLHV/ZhxDpwAyMlXOuxbLaohUeuYojIpfVJIFkgJAhM1PC
EstZwtagJ+jXqJHmjO2VPis4DHJEbmLAzjFGmtF8RlvYuvYq+/t/07VTBuWhVqs3
s0QvI6ZnzTeIGpWu7obUZs1Bx8SXdn85ibgbilUjCAsWtua5iL6UNcmfvkjhdI+4
nGkVV/BU80DAckfm0grCl4JZYUCtIjX0hxlA3i1qiczN0g3z9xgIplul3z8k5vff
tJrEnrbwDDJ5UhbvV8a/SzvzP19+3IdYwaWh326bXtRXg06AtLtkn7/LYFjFIJb/
rgJoWEiteOR3CwqAfcWPfsvnqNsrqMnmN60VnjLgK1QTDTtjKlnf5gwlpgJiixMa
uTYzZflSL31NI5Pro1dIuG4K6OGgVhlskZKqNXcfU1UvyM1FOOxKiJLkXDFgEu0x
FwvBkmBoDsfccFZwS/+AFm+tq33m8Kg+9IYoUIVsAU6usJ9tNyvOgwpxEqvGF38w
YBIvLKa3Z7jQQ+/z5aiUEADtyEbW7ScQtwdeJhi6aaCWS/dsShRlH0LQ/zFUX/wA
Pari6vqMvhaqjwwfAF7vl0Z5kvHdLJbPm4vEWjKyYIkuLUD56C/Z8M8mCrJykKUC
DlQsuryLr8C8o1qDk2H4aX3ee5BuMlBAuwfyTfPEkBXAfWzn4+bGv6FzpGghbIRE
wl/HRHEtSyuXhGiVl2SjRb/0HFTY9qy8vULl+uJbwQoUDvDQf31FG5xMJw5NLQLH
ueEViAszDSM7CNk6Cq5LTVNdE0dx4qZ7GpP3/gTG2lfbfSokML/wPhd5KoQxW6cW
be26DJpVfsnpB20KKmQHOzraSugwL9CJtZUbBee0TyAFBNkFvxQ1FGSojAJrc5iO
5LznaolECfzGtZloR1xwv54QK7BTqoHEI1PGj9s3pZTSJwG4RTG/J2IT+BSO4Hj4
DtZBjco6U4cnQTLss/RrcwZuvk2L5f5K70oN7DdYoWO1fcAW/rsbWpjiuKGqHMdv
AWtkxtHVSbq4MRc5aczCGppubVuKXSH6LjDeSvtMEve3HjtjX7VFjVNnEf0zRgVA
y2HGzvjgTfb9cgSzwgH5EaZ7N5pKuH6TZbGrb4xA2FqPbfInePXx0CshfZd59/yE
9FOtwM+t3wS379r6gJ8xazeRPJ47uIGP+34e1Q7hXTrd4BAkwvBWNhBGyb9aNnlE
ikXXjj7BeXytfM9mjG9W4OU+tOHfTO/ZrvN98AZDfgj/T8jK7j8vYUwG7WQbAiyw
FffVk1aeu9jmUMYzK4X5zFKUM3S5lP5SXUIWaSjLcG3z8ZMTgOXpFesbKJhWP1zv
X7whinlPgMsRhD3Bvms13IQXMsuY5IHfPXA2ro00KRtUlqTsKBjeJODF3Rd0YAOe
h62dFjrxGAwM9V8XlOD6BjeCcvwNJLnstjhaWopSwLTxXJRBaJDEsK50cZNvuHvx
Y9iQ/YBUxbGj8HU7Qzntk3/3ZvEYxQn1iUVIuLn3y6RvLc4aRH/9pN06QGUTzhvF
QfCb5w8YnRn1hkOxYRNSLhzmK3LgfjyKRUe5U+G4YyW+XT7/QX9uHrfakYpLaPTd
2jrIJQdGmPdHVVsaM4j5+mxbaePT/IisYne914G7WZkBTed5g4Ph7ACFlPfVtgD8
/3gNu1xn0BThKDCKBqE2HLW0BsrEkCv0otVkSUUkoddNu53AKsLr9Op3pTH6klIh
4Qz9A2DQCEJ7JRf8RUsuLFzqT5V0bfVzp/rdvmho0Zzmpj/r+otML6KHAYF7/kNP
jRSH32lGBYLNAWn02osu/KY70GZufbg3gilnWDv3YGslu7fm0ybPRzm6PHl9Rt7B
ERpgPxan184LsbXFgrmXqPGI0xP1Q1WgLuVGYu7Fjfk2chxXkpvfj4+m0JwR+9Wx
g+YKVL25al5Qj/rGNCR3hAnnR3Uty6uCXdU3A9B8LeCVI7aqzFbT0jnqStAc9X+5
NWme6tc0MaCfouX4lejHRmqzQuD3/ne9+0rkV0CuLIZQv05y9tBNggKo2IPqFeGn
JgHHUC3sdpGI1LalVFgBPAbMEcyc18l2Pn+3letrlqO1U1hbqPd7YR61RtZ1AVMc
DZYbECRm6g0ha3URRXHmXyN5nuBapmMWCs93nQEax4ltw5gAv1fYK9cwUGkxALQW
sXXlF4VO21NS8o5hWXwrHuUBGOQZyafDiEt96bPdK7naxc3TqTs+Ct218inl+tyW
1ShcYRzmHlrSn96W/kHrrShDJuqcuRHBz/4JtIZN5URoJk/R/7jX5yH82Tx1nb8I
WhT96bnB6ruQ55iIhSNanzhAWiV0AwpIyhlz8GgbXzR2uM6FdifrtJQAKBHr8jLg
xE0n3xe1+qs+XZpTAJxh3dKCK8QY3+fNWwE2do6t8+hnpCoiH8kro+qmcCKg/Anl
ORKeGH5M723pqp7XEPZTHjC2051F1ObLo9ukdaHMFfvXdi4QNEH2JSUXkg0lU6bf
cS7QYRqfYlL00Nq1kSGwNjk48vd4WRPOSdRtA6aDv+SmLDc+2XKk9/yQuDkdtlBv
tE2LuMb1dVdVWH5VjARSMdjt24HC8o+Ut5lrWPCHt0k=
`protect END_PROTECTED
