`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VUl2GGFAJYetLxD5z0++sTuIRY++CNzMS/cU+jDp4sLQZj7IGVSGXp+1914QeOAk
Hq2M2LqdY97IrSZvbt9nrvSEZEFiNZiumOzkh+JjMI3eErbB3B0PBKaHaZzBIPuM
mV5dYvaLAuksTObDVT0ONaBqB+iE9KrozEpiqjkeV7hP7JDwwUs4OaLWzWzLT3+C
FdwBugtQZNVkpT0RUUAVvyrmltZcNS6ctTlzkFJ1EZYjayf9XoQWXPlvyWQNGlsx
/MsWOfHLKxzDlQAOLHLCQlcgGG89HJO9mBm22r5meOIaPHJmzPslIMJDF1wYRKNP
O1HsjpSiYJnConwdukwX9ALaE2E5g+x6IBVRivSdju5uBwFc7Y4ztDuEQmEbLw36
T+Ewf0mHigSdmBdlPnwyTw99SbfY+VncYs5GFURP2v65Y0JCEm958axKB1MwfVyI
3c1EHu5CEbFf+4m3oMW3O1TEyj9rxZx6cwynVqDj0nD3ZXbQEHD37iD3kZUhdyTJ
uW2mHtzmi0gRxjnaQENYvM++MX2l9dCJUNwBksZfgI7+CrGWpXQg1DDnkVjl4/cc
jgPHMgmiWDm9wdu8ahl9jaO/AQZ4jejwR4M76EXXZ1EzXqoUelS4OsHxmGJyc23q
dWUU7YsYIc8Tg9UEpmVACkj5hqDYYyc0JDxRTwe5VJY=
`protect END_PROTECTED
