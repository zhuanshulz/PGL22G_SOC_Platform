`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1TFt9lCYAZ8+ybMCpkvUkbuoUUlQTtdC3pruBXNea9CxL72w9NoV+wNaJsdjCTPK
u1FtRvAbVr5etsmILxNPxFtzV3bcExdo/PcIOQJm2AlweZfWY7KcEDBKLO5dTCdh
0fIAKOPIweJGPm+A6bRV0KqDJw6ttAO3VPpOd6kzGLr3xOmNymB9VUqMOkYN9dvo
2t3WyfymKlqO/a4ZXQTcau3gkbx5+4+HDIVA2mi9QCmCSpRFKcPaAJwCzGRC3YpB
EPk4AVFvqfiQRdOrrCOE4cF6FfBVmDHOcyyXEkkRO7wl1mLuY266hSNiZ3w7uleB
p6geJ6tbYiuu7Ug0PiVjVduckY/RW1YCMIPOotIFqwTNBAuIRHl/oQTocYbfB93G
wFT7LcPZOetvkLeuKWQfA/OPZQPSumysZFuCxOaL+znHPRA6jk6oYZjNOdAiNlj0
KC5iCCTgtZiWPMDAep77SsEx13X8R5w6cBT2FEOoJwnsm/YXcf3gqYmkNTBXy5Dr
/Px7DSOwzPogbCW0GiW38aYCLNWD0nWOHXxkMCS9fyvEUTrYk5wSmM7lQrz1k53W
5Kxmibjgr6lwoj6ZC0eAhVZwWFFrq0YvoHqUI00bw7WuBarvZyVHI7TSMXYaO82T
4qis9gkKJaeZ0KDQCJoFUeAatFFglIZEayzwTwJ1oFPYmP/JyxaDXkgYl0yNdbie
U9nX6UIFGpploLLle6GIaOh12igqnqLui2JuQxWZaafpJ6rcZWSoiFjUJcxr9ReA
tiuzl84Yz9TKlv0PWAcey4tSdUe3TGKbZiJxU2raU86KDjG2tbPx0c2bE6l4tkav
yJpgyDnGE09SaD9Z2emoCN+9CfLxFTTr7prmG7QLVYQHjgOPQSUm0lzImPAXstEs
ZdpM4OLey4xLsoituyuKJSlBVUI5Q/wWwp1Gc7j4AFj3MJ8eUGu7JIr5OocWLPnn
Mlmd8+1Vap5zHpnWMMzO/8Yot5GzMTr/nAoa1Wx9mr9ZguuZffLi/wWDJKijqFTK
gULRDua77zKc+1MutKMHqpOi2xoknfKVkkwp+ikzKKK9h1E+YxGRhOb93WkYQMMb
tzJWxF6YTXVP+iUkSYVSx3rtqtK2eLfnSsluefHIDGbf2UQFmKsCpNqhDJhpvplH
cw0S3CkxeDZZnUoPOck+XvjnUOV0R0NmmXQsHHhg6ZC8zpcJZ4s+UkArHQpcALOR
XOP7CKUdNSdS/hoft9oIux6DbMZLCK4XS5Pxf1pmWm4t1KHfeyivE/Og1tyq/PZo
ssmlyMgCxJuPfEyjCq7WfsSvR9CpWICUmR2SulmbVLEpjtEOBdvqT5F8ks9HikoE
3OwWC9642sAvLKbe77U9vkl1FBMj2nKPkgeDl9Aectf07qMUKmx6h1HmANrROcpN
MoFsnDRhQ16VNOY5i7OB7/hMScqYIS7sYsLRwKfPvfom0odia2JGaCI0fHVDoMHW
uLZdN9eNetoYcisDc8Hv7hz1Q9Ei7Rn5D1atL4u4l+WtJuy2zy1SdEq35LOFxVkb
xO8WqGin3dNtdnkSn2lrVO5B1J2JkqRlyj7p4DQIXJ/EHhPMe0ztTB2+ogcHhuc6
4hR3VgSfH2/Vy1CRzGjBQPzFqC6EIogRokT+O0d0ghhkbUlm+EvBhtPNg/2zoMcM
maBnaiKgndB9B7KD1b/S9KsQZssH2v/peqhRwdaCJpygyVgRHlmh6rBZAjDZ+QqF
EeATz6AjWfVGNRvvLby67fwZ/GrGod+We8dzNjDQwpU9eAcpVXGiAMrKe7RXBfnB
djMxuJIXkEgVMN3BksjQ1gc8Ib93Bm1KInFx0abl+It7aBmZHIhIuRsM3hmArv81
sm8n+m2Z0e+nzsvqeVS4X2isbuaI+2xJ4bgmmL45T1u4cKbSKjSECMd32v8ao0gp
/lD6x9eCY2MnHG9K6r2s+b+iFwRT8ClSK4paENPONHx0CJ84sabpmGmkYWin6Q7A
3tH++CvCQX3dvaUwN5I1Fp6U6KVjF+3lbholNoyg0qXDIdYbGPE7RsI1+3cdTI9v
Ma+xZpPtx8ZGRkYWdajT2HbXF/4VEOCGVOLHODaBhCPIamLPNu0r2yZenKc6vwBP
6E+1wkVCbPYMAi9jwQosCBk2/Tfym5WlDZoLDHe+fWkLvwhSqRF1q8f34AScFoyT
NpWJaX4uRBdOLdNrbwWbUd1sYBDZw1MPJmL2P5ljItWkbO+hjjRr3H79HEWDLRYV
ZlVDPSiGIR3o7VoRZjTHhcCGmFewFeXfYeo7NopdLPr4h3r3WQ+I1oL4KyFt+Nwf
Nt0UXxQh1SGyHjJa+l0K/8Qn+NCOcXAMEzFLWPy5kwQIMThcWrp8YZP3h5+JhK0x
1MWwn3Sgfzk0gx/fZws0iralhTra8HSjWZ7X4mfW73PCPgfkt8JPLx5BBtNZ9DgO
GY9avyIxoJvgC05HHZao9nADWah8Kf5k+66dDabMDwRuWZav02MdYzygxPRYKYd9
EsFGSIGgaxa0eKY3l/e0FulfiRY1GXYTdTr06pehITPCk6n8zVEQyBp4VSDOJG6N
lJ2ycZMPEArEvnHeFRLW8k+PIYvdYFFTJyBqhDPeXnXMRXl+Cb9KEg9q88SigXOX
3en+LM6jFDp1CAhxB3gGRWE1H6y2hddaoNyxV+NCvAnTtl/t1913CGoeNyXfivt4
sy1FBHhWsDkG1EmDmU96jo1yFRbzlBEKY6UL0guRiQt4TJiYTSaGj6ogGd3bTy4K
Xn8p3v5e9Izr/sch4sVf0XM+Rdcb0ODHviIJYZlUeL5+jfj4BRTMH8bFt4Fv+dZZ
mmvoz3+zD1N11whQxBD5z3AwaFMD4N3TRySY5pv2Yg/kMZNBBfjsbzBJMhlXapAA
xyumzHmXgo5Fr/nRSYU9ygse1p1ugRLig+QK5V9Q9ZxF5JERVldFP7O+Rsc9mzHc
gbpB5KI9+FhNwAhH4Th4PwRHoC7dxbshpKncuXQ5SaR/YDO4BGZBTj1GSSOJvsxX
snzQv0edaper9XHueGea+DnmHnhya40GyBwA6SzreNktSAPRDbhcta5q2TJ29Qa/
mw2SmMyvhu3iSjezUrIbtO8u1Xj7vaRnAFyCaDqh9jNoS8T1vQROu1/FG9gToOB/
PeowGuVy7JMKGg2sUDpUrcWDyoZzPqnDMdrNIBiXH5dFPUi84V5NP2cZsRvxr4Lg
05ROqYbL99X0fJ3NM2DDhgdI/xfw5htaBNzMWzITxu8BdhgAuU0uMFIgZJrvKVLn
S/a4X28pJW+mag0L3BSlRh2e2f/RxYNeQs8kDz9RK45ZgL4yzv3WVNc/OkINaS4K
EdwlMn3xyXYpvq90Tk+91UBXtEcyiNW19DLBr02RiefV0CjeCWFsdkUeuSNWHYWX
DCd9wcx22zMJNUgmNKA3x6yQVXJL6t+yNP+lBFjNnCT0sSvQVy/yQzN4FKbu5oW9
oAqZQH32/x+QuUSxUfZ2kJBUOD0zfNbDkbCLJygRJN0XPQznYET6GOIWNc2cWWze
V19WmMyLaomLA0Hu+G+hTYtfcr3SAFvLfxFspMj19R7H3XgejoyWCtWFUuFSF9cA
d/ThaTF9eKwJxl3f2gKfUgzjCQYUsua1y8DCB/6iaUtm5DrYlrU1XoKBJ1l97p1U
HOM+RsDgmbt25QjL1rz/rL9BbCWKpNMi9uvyPjDH5fwnoVh8cxBL7KjNTUQelPRG
RAcaOE5qH9BQvuTW4BSB5PkBwrv1IN7C2Z9pyjF0f437sCSgvFwXViq2Q5RS5WAl
vD9QPGfhWxzdKZNVe8bxHh1hGyxMsBKgyzWZY+eOsqtb9RSz473wNtoATjXBLRhV
c0gjaIqFTo8vBeGGs30J+1fJ7jqCOR+LoAjzYgHmXwj6lksK5mo//qNVPUcI/ijI
g3AW5TPv/GvNRsiwDD6d+byKDCMEOBOD4mnS0TluWEh+V6sdGsZ0gZwveiQf+aNG
AM95Njt7xhVPzlF/hX6Vcrov8hJNqz9kBJmb9zAIYXb0yqqoI0JZRxtHcqILSOvE
59KtUqQqKHASZZTgnKbrgxXFac9QpMA4lkGA9IhDJOqH3LwPZOtJTDQSw4Juyblv
3qk4NKmr6bE/SxzfAayK177wcD0igJAU4JWMToHSXzWNRJ6yOKccpr/OnfB6Hn8Q
tHTKBQETS3f9dgShIYpt8ayX9WR/QyJaW3rRz2pAgOT3R5mgao4r0w92q7Ykmu/j
s6onInn48kk7lXjYG5P3rQ4X2fZ/Y9f3UYLD766+BCd9LXASnonxls8QzdheqAdO
25UW+yrxwELbYnxldozTQ2yaPpwa76PD/0NYPiiMWElwIfH6lFc2tahJVMBSbvUM
xDXjAeQksg2G9TF3Bm1NXwOP7HKZq70VdGvk/5Z66wrjn36Qcw2lN2F+nseNBja7
39CpyOT2uqfX6FlrnAr5bPL4WrfvIY+xyxRyIMvrqVIGOS3jcHdMu/agdJFF+Wkl
GzPXA+ICDxWe73f8ZFu98k+gByb/37unSHv8wniN4GtFQgEPmmxC8Lg3F7VtSteB
7Rbdy8/XOjGDdOvfRisYN0l7/fSFPvHN3s/aGQSKaiLh6d+MU/ec/X/VwhpGICP2
euGTlgB294a3y5STeoAKuEdAFC86Vs9iLyk+0jWnGUc10Z3gnHrgXqUUeG6KQeV3
uKoaTjeze8/QX5I4zvkRi883h1W89Z9jUXgw7Ky2N06CBy6ZVBkIDHm/fE/+29NB
YM3foAXNNmAHGp9ZGKcoYrBX15dsAtfrk0YLCOII43As4AIG3Z1fCXx6m2Wt8iVw
TB9xbnZXgK30kOdHVLGqkf+RUaT2OgqMllOsR+i0/eI/k/F8wVb7p2cJNC6kyspU
xMHKSziIeiBVlZMbYvaIgjE0MExN8Mds0KiQg44raQ02mukQDcMVTJpZZrjrX2y/
3AD2fV/AjB4ytOHcM8Vg4ust3hBFoTwQXUlpVqxYX8qBfLs0jhEzfPkiX5ylP075
+asV0hSYxzIH6m2FC+S7uUnTLMdARTwAMki0F+fehhhl2BTq+Ks7suFaF8+Oq8RI
e2EfxXEjRyhNYhBbGJFBRPJpBjN0McYY8s82oDxYlxZpivON2BMm6icct+43741I
Oz0t0bVfsoQMAcdxDxSSbMNZxp9bgvzYp7k9FhVF2iAGhVvcLIH30d00e34qDEVa
3Ua0ufeJ8r7QeIDH2S8NS3JVgcOcuLDd3pAZKivfs9AFtN7Ocg+QSfS5DvaG7bVe
U5Qn5/+zk6eVEzL1hXChJzWTvwJ3kaeLXmupPkUwjdFiAuYw4KhF3stSm90ihclU
fLI/NLUilsZYfG1txvURxcY6JdgAoRnZawpeaFuoXbU48PT4nrF9X7Z2O0qt3nxT
Ik+N8v7ARuiuKZnB6RA7SARrQqeDc1n7lwLlpL8GwULpNCfMq2TMwAqi8ZN4p4T0
5R/gxbOb5nKdlz2gLoMeHugJ683TgqE18RV3yma1mZCutansjAVW8zNbOtFa8Zs5
2PzLyU5mnrJuFn/2L+QdpQCIKJas6I1Y22DbHC0kMZ5f3h9iPzNdlgSeo1Bs4n2F
xjid0zL/5AlEMi32qQzme9ZThYNdOThrS8QDXdYBHtnOZ/GGLA2M5M6zRURJL/3i
9L+o7OvHwIu/hM7fG6SV9GKCjIV8T8RCrc9ih61EXAWp+HC99lK/3Jn+KeRuzPHD
ZPhxog5vCtTTSwgVZQHEESrIfglzVe3O0t2lAXLBvRH+uYFHSYitMABMBBYlFYNF
bfMlbTBgrMn9fnaHOXlIE3pL65G6jy5XhfbqdCngL1AEn9dSDVd3aWs7GR4rw+sy
S7MtcXWeqOEpG5+7zCpN6bGWB45UxrQgSctUTbUoddHTfNStjcRRVcjUf6zUK9G+
XeHZqtBHmOa4lzsrr5AXRQkO3fZVe4ljNWISBDEqjhM=
`protect END_PROTECTED
