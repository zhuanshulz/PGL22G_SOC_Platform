`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fHlSXASsxvIqCNIjFaGARn0YiTs1ouqq2QVOSuTqa4WB0H2XB01E1SSE+sF/rFRy
K8VVOyeBoV7SWs05LBFwFVgnnjRBO020D8ipKL1TWGuNZwnqbxm+kI1RtkIqDr6Q
NyyFJTeGIciv5nPJNDOMe1gnpezicng+gA7eXb07A7Pgu83vUUmLQv5DLH03f5Qp
723oLInIieRrbzdGiu+HhS5cagay+nXZ9oWLWTxirdhAGVTb5UqH+Edk9JfRO/sy
ssFMFh5Mf98qEAGl8Iuorl1aekshd4Lp0Or00GJ37TEHpdZGcRWsF2UT+JNfGz4Y
g6eVWmxZkDxBXbhrgINjwHDmHvYnz4M1Wc8YGWwlTCQ98FtQKBRpGSov/QBgLZrt
72SdGoOZVqg0ISl9s6btaOzFsDiRRGTeyEc2PjUh/yIA0C9MJ7rD6eGeg8s+zPbO
5dYSx+6/5GPbhJETUbn9D6Vpcl1V8R15dHBJycG3zRDoG4E/rqkQE2hzPJxq1BXN
PiOiepyMxDKIzDezVSVs6Je444pXwOKadkjwgIR4qKB1yHh5m10WjIf+Kj9j1+3W
/CnvME/PxbYQQeM3QF+jKpkBlRUt0HZQFZHrbjOaU9ZxltactXVF0cBXBj5/eFWs
OT53ee2fe4tbVPuT+vlj+Y6EoApjh+b2gntmUsFkYiCWvHBpHT9Qo314ovHdnGy4
ptYkxkuzIuF7BtF5YHglP7YnpjeMUYOpNuahJBzkx/tPhhd5YoHqKsjfUWNYtkDU
ULDgeoDfYuU7kCUDyK8eulMw4kGu4jY8U3EpNs+rxF7/7UOHXmqWy6LUjTbNuYfy
CkrSxQPjbgXS777w+/6kxFh+XsOpalPfIrafb5Du4nrLSi9hFd+JjUg70ZiQ1jsS
UQpUkZPJyycUr3ddfNA2cJgUc4Y6g2tvgUnj4wCM9KQpN94mRbYdfMSovA85sqxv
eMmCEkhLu8LgNhQlUYurkGzxGaX3UUzwGjZc1bE+GdF78g4IghjWUTuRgK5E281q
`protect END_PROTECTED
