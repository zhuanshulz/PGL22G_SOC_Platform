`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pgHcfXOWXjpFmL9j1C6sr7setue8zoUQ1MAntQJ7Pipc2gKyCGxQLPwuJpjc4JN6
V1o8PmyNR7tKsdlQbDes8A61vHI4g4LwMqtCOM6wvd0l7Yi88HRTEbCyG7hDZTKG
zvrckLCU4mZFEC2RlVh/6OF91x/5DeCdUGVwlrNR/PtJcZHaq0TWmrFstw+Ro+97
+HbdJbbXuZHzaSvSosajg5qN/AQH89W2wS20AJIAn32p+IcdRtHi3W1qW5ZUn28w
n1YnFHUQNe0Bt6vdojSWBdZ2woHEkiNHWMURWa47bv1aTKx885FzC5w1y4U31KlM
VJRyxc1NaLZzuE7BERAis7Z+GjP/uxQWeBt/uhBB2xbwh4loucsYhI4RmB4HxONj
9te3CabwYS86jxb6eVbZCNe/XAy8c23/dm7G9x63BCxYyZfcYZKBwY7nzc5RW5/V
UTqbWzmu32ZoT/lfKq/nUfKeQAiETA9J4tE4tlT5Pum7Jj8z6I82OpEppko0a5+T
1qwDEd+PY3e/LayfImUbmSaYSuMHDkgZq0OnOGYTRomx8e7UanQ8LuvPYKeJs2b9
V+8Ap3f7pWo4cF58CSQRqw8Ns5bLhb0Ob4Oh/iosOf31/4xa3cJ9q5jkAefln6Fw
4H5XF6OL375yDjgwb24GGmdMYqLhqPb0EMDGDylVIjfm18LZhs8as9PlxaOOxMes
6JmrA5n7BT79qFYRwXmnXWMjqmRzem+D/envzS+t5mXttpwfsiS595T5vgW/S+TA
HQ+JkZDnDck0Qki76L+Wa8gK1fCStB8/4lz286c/bdhmYHyxHTncx/Ra6+MX4NRM
FWwuZIF19EL87G8u/MsDwcgI4/3rutrczXDJyD7fvDTOphNDMHIgs6hju5PKpTb6
/tKphkpL3/cVX9EQ3A988VTgujSw1WEoRUK4Bs6cc74+g0y73eXDT9YdOP83JnC2
`protect END_PROTECTED
