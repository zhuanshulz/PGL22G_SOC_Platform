`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3motLcCnHV3iU46XNfrrczF0sebkQPnNEjlIc1/eb0y7HZd78H+QxcL1EaJKuK4t
hnLl2wQsamsb77UN7NplQuTAkOSitT4e7wRwOhGYCEVzzqWogPgaViLmJhvqsg+W
4UDcKIF5UQzg1nPdcJF1JkIezv3XtGLufRT20/5R/m2hV4EqGn1RzIU2DTbTYp90
q2ytNufGBuu7kRmvv79lbN23wdsuxY6SX14OpGjA+c8Xg9YNdzyUCBmH2epYupRk
b0nNITJGsX7W6FqQEgHY03K83faud6DvRpiQSt7kzc/2GfGR08tLWYyDlV28Arav
tO55ps3GuMfk6tbxDdhCvN8ndg6xr53deYXla1QLHeippCIyhPxQSo0zqtBJWnrL
Y7bOdB+ILJ5coCeGh/JDIc4i60nXOZrKQhA7p4N0YCTdl0VCUm2KQUB6jvU2OPmB
jqhFKWhbZBoQ+AEbMIG2m+XSJo+1dK680tFu1WrHKiG1fbgxgA8mbO1qL637XvhH
3GmfB0ZF+JKV/mVCf0W5c/QWidEzLvufloUtO79KXCDeWED15/OpE00Ols9KSxel
nBtWBYZWBb6ORJfZDqjujJHzkcIwiX6T4vpYwu8jxMF0IgxrbbdwO9zv33B+FSB/
6Re1yrGZ5o3kOUbMvEdh8yokYZvWQJXiQdxEwSAMsE0r2DEq0z3ahgYyNxE9yO0S
gMADPnQnbuLvGmXk8My/qOdwWzKqwTnBxLEFZpuwPQAN3IsY6P/5IsNOwW6519uM
NrqbcaSKNLXqqv03RGh2I6b9NUz/RICvA9eyoffa3DBqifOlj6MYhicX5SREbikS
WpBSHXj6yWD7td+3EuyHf2dxLVwRCim2H01OMHVWMNQBKtrwaTmHhg0/o0rACbP8
IxRWxyXnw/vjE0ac6rN1LEX7ad/73NqtTkq5tCBHJJDxb6WLcqMWfzGhuvH0lwTo
VqAxjLXjHDWcP6eN9tVLIFgOuVSsElae77u8Yzujbj1LlceWlVXcr7jFvO5Mqsxz
YRz8UtSTdaq4ywiMJYG6hq/zjKwp9fT4uOlleQ5FuCvFo1l1tosI7yIzOkYZhlNp
dJTcYyKUJlmklSfczGLzkY5G9lF/6kH2vzw6E49AX9GzsGHuNLPDQGBAajqVkPrB
nNVQ+pUSIrsc7jM75RqqtEsz8umy8o1lydBlTqWR+3PnS+3gwfp/pqJH89NG8T1K
KSOHSlWNTNQ8SAT0+lmZBcvNn3MImVeCtrmgolyHqOobbjHFScoRL+WXjsBH7eQH
RXQ9Q9BZvb6MJNiT3lEqlChbxWIvA55i682QT9dcIBX76XcVvi3Hg5Bd2/3GDirH
7ECH57Zd1QNbdAt2YXYHAebNkafu/+4jBxn11iXDOseuNV2dcQDWIOhxNRnaCiBu
222TT2ve2/92G15TpehwSpsB23v60xOTJI8QYP6dQ+uz55IjiqQrtXQi8fUXmo8D
0d5db7UDQvIWtom56hi+0VNV9FGJPqixV8ILx5OtQPaxpzHs3lX6/rb4OvaONyV+
5cwhEtf85nnw8VBnEduA2bIO9cIQ2ubKbzeu+//UKk+WQJpezCmZiiRkyIEMowgF
OEnizKPNva0XFBUdcN09OZTaNgsuut43lsC2xH/MrqOBW2FrLPFlrMvaN0RIHBZM
WLoc88/QEQWiG+5YpvCRodm7HpRvl1yTmR/TEWlbo2KmEerlS6GZec/aFPMr1w0D
+TEAbcFtAqkrdhWTQNpJ928KZu+Ofecuv2xzmihAb18f6ypdB59U3JAT4OJWkvOU
hUDh9qn1dCDWfVPSejlOh7sF92HJps3vv0M8pb1lmfxMl6ABKrKd/H71fgpRsQTB
RjOFM28lrfbhFD27S77ORki0JcZPaC381QHS23pxjWY/yDMRf/TMDKOgmt0c3TAN
lDkSJAIKpS5ri6bsNdT7bb4IPn6G0f9OvN4nW92xbaH5eX4sp4jCdnzkEYe2Um92
2NvYXZNdz2Y0Pjwqvs0lRalr6aaeGM+2Q/uKArUSE7UbY5E1g2eb9zmDaCLx0KzS
qUjfzWtomDgADGO0yiCR2HIbXFicV6YjVTLVYQtdRFBlIeOxOvUmhja33pMo0xu/
rLt1ewGIQe9m89Qiq4uaGBqXzTZRiVSWUc92s+HkDOcaJTxXXqJLP6Unou7olMqh
fA6oMeo3MIws1VwfJruZOreaciYDrkjtVjuzxHCVXTs/Ms610krtsj0EPbuwxwgc
XQa1S/w7EwZuhXR3h3OK/mF4Ew8Wmt2tAcp60Yt+u9piOpk393J/yraMeb9rtBSn
wOEjRTsaja/7rd3E7aJ/gTp8nlUNOhSZxQzjzAkgSo8eFQ52JotAX8UHbOSHa/Eg
MMPM/s1EkLLtxnAO8LDZ+5ZP70dA08OvyE7bEuUV5nbwd0g+UJW6LG30lSdPfzDJ
vE8CYNXXW1G6TvUDsOYdPWTPQzAgXHYLc/um4MrEEILN2ODFF+KRbJeBPLc+hztb
UF3LjETuBN12tv26MKFKde3JZIiXIav4LDU7SSFNmFobmsVHkK1Nc1VQVnZjoF1O
WvsQlrEXb10c+q7+9wYeLPrQ5JB0RhgP7tOZljftLfc0aSw87GGlupyZgivy9/sh
cKOGtGLDVDeQnuOEiuUpy2yzablIpGblJFWMjkwJ771qBHt0mdXNJYkvtMBYg8t3
iFSMHrr084+3/lJQG9/zUcDeX1cwFQKQNqFFEuoCqDnbAi7Q/mX1sOt/BZ3sYq8i
ANPh4kn55slGeyZ5LAvltw==
`protect END_PROTECTED
