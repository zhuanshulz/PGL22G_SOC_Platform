`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L32yVWasrqPSOHnkY8sezLpxi+vvWGrbxxxPwOgeRROjyyLJcGJqFgsoyoFJ1kdQ
NpX81UBhoKNEsPxnbFqvtBtjz3i33Ab6UHbZ5ftih/27roJ6UiPNIZqEQuRVFdE5
KtjS7nUJ3WmTf1bQSfmc5mJSd4pp+XPRz6y2g9I0jFDYRwztuJqb763Z4O9IBFoq
aquxjtObf3AN7hnehLqqkO1GIAL7SmRGNkgiihmyEGDUHz5x80RpfB+YRqJmxtwN
s5e8P/sSRxAt5DkxiNN2Aqk/sb+6WB1DxqFRgSEuut0N4UTQHdlP6SNHTBZk561E
YzvOJduaoBH/YLBW7+FSdSnlvq7qw0rXW9QXuxxMCvtbvqlM3l09mA2/zA6mCng8
ZgYrb3oEaznIt04cFKFVLGHWlMNo8nsz15/XowtJ/IYPFd9YzUucm8cpc7lpEz2F
nAyzVb6yQJKNsRI7QFePKS10kMPEZ41OR22nn8OyifVGyHAyvs1aMbGUljrM+dMK
a7n4S6U5TKWwmct9VsEJKXFGmrvcgtzcW95N1rQ9oaW6InqvxHC5FRbSgBS/6nrV
9PGOIVMoCyW0Leb7Q5YuM8e9R9KWuGF0u0LGRN1PRS/wn7hAobU/GAiBSup3HRdg
/y8uUCpCty8RpjgtsTuMaLsoM8lUOOLpsk7zTKPdWfd2QURwmpK+x0j7rAYi1Pd6
bVt2BbF/EOb6EGNzFqIj1OQa1vnE4K4xGv7d6DcoX5JiNf7S9cYjS5xq+uC1p0/1
+r75Wc78fLJSUy+wojskzXDIPk8Mkvzs/PC2w89HyNZX3obBB5pOFo/Nnk2RBfL9
3GrGHcSZhAFChyOYiE/f+p85GXjATLdHvNe+5EqFVGFvaufJjvBvsv2vcXlRV3e6
x0arGityhI14382L5+haSB0KkeJ7mcRMeiVLmnu+USWtmOamAekqd+pyyphp851y
Lgfh2/8cI1/xizjhRs84EBWk9WmK6FcoclcsDuXFwxmY3nFebP3Fa+2fPfqLugu9
r+7XDm5oMa7qh5hE9GiL3Y0arh9Vk7DGmYgFcsPNEnNhq8VnVkit0mEWftEDjSPO
6UQU6twtMqrukdUjVJq/yZ8GABebDiQtjhnwBzYSa7ugZBmwR9xOg/suRjEb4n+0
Zmtk38bdg45/wyaaBvElBSSCG7Hy3iN5sG3nfT1fIPFeMpFrqSH5YQ0igmSYJDkr
SAI1q87haYmEN6aJzbocUklSaQzfuxZ2kLCTZOgPzifY6Gp/MKVb6bw/ni9RhZqf
DtJpPOmX+m+7N2tJv2/bHMr3ZPhzf8G/JK25HUOAJbS5FisN0XwPNjTTTwGn6gh5
hCgtM7jnsR14lZruLieZx3zqjJLjy4JVoWXwrRRgeYItsVTJNBa4qsuourXLtp7J
QwCRi7IbOj4g/VM+1DipT093ykZK7Lju2cH9GESLlc5UPAvw4kaAr9Xnsu+5hjOQ
19cUPaObjnMFKEwpevVPEHgqsJ4f/Kit2iqb/MOcgTF7FMoJap+aZWHnkUAUSm1b
ELF58HYLDAL/LDbyrFVxFNHBKzO37mK88d/Wn9DNcoKrmQpVk531viPkwSYDpFhy
MUbe18hU5YgF4ijq9SWNA+uH5ZoCkgM5w448Y7FTKKKj5++f1xCvUmXbhkT2sQVv
+qBc1i3ml2Yed42wpzGO2ObanQAttCNzMqUhdCK7KbPmYpVV65wjURg5sCuPQPOL
Tw9oqY8XmwFSk2tNccWZLk4Vo0zXhc3fWKYDiP3BeFEvthSzKlNlvgWn7x26Kkzp
Dj7IzE5n+CqVoNVviyqVwtGp7mFLLOHTgsJvASFfLlKlcesejVRocLAZBX5YO9e/
181pBJcdHliAPpDxrFNWjDl5zrvrtBwOBkRsBz+FvT8J4aqFFZV48J9wO23DA/lU
ir8mmMh0WaCzvCUqAbkWaW7gQ/TaHsGwHoXDSIw43ieUgri+7eyHiYAb3NzNg+8o
M1EQNWaogVp/uwp90y67LOxB/slWCz3NPuVUHaFp9/JgMWydNQV4QfnXiz51YcN7
MEGzmeXbfGbJSvScthH4lm2KJ3IXRPRtGC+QeYPpblxW3OP7f/+zRU0zQB5KIJWd
GmiSLSO9ArxSJfWu1YNieAdk6au/10Gl09DzaUczERVDsfNnkrP7ho52lyFrOJUv
tJrjV+we+VtSCeikN3TTOirL2Xk7pkcn1O3Tg2VJLRH+Ss1q9ocr5WZEmeWeuXll
VQrp5Ki6QqyQsAYteeOt0QAHssNWXi9W2h4+ErAWmXXKimaif8A3diXbdbh86uch
aYmCgdKiySKLU+yw3GhX2F8bLaMUn5Nwml1pKWssbEf/qiJ4XcjYDXne1xA9nH9F
x7Uy9U5A1+OlsOyrcfsVxPSLykAb8xEHovHEtTuQ6unns6A312DHVbTl/iobZPs0
ndzx7inwQCiG+VXm55QSpRGiw3JKZrRsgtOabPVLxIWtJo0DFL5RjWueLgInCGsG
eYOXDcFBJZRwChR5Go9dKmK4cTwqWH1Ag0eSrZ1/knA6QZbBr3ExJ66eajGNzpvO
+ibXzgDPhmoJIKoP4/M1pszBxncuhM4KS7vWZgwg8NQuXz+B/UIvdTEBV0HZSLNG
HAjTSqZBrC2Ekjp7LsR82gF2S+ML6FaIKIE4lPMn0Pgg10h+GsXVAMFzL3Lq3LwS
cQ9pOwSNoB6jViaKl7pTZlXAlR5HSeYt7w/zt/NHtZtqydsjDCEQ5YfR8OEEL1VE
jXS8HLQweZpwfvYz/gJe0OSfDHUZSwYd0XiHv1e+F8kmedlOh46kNzc/mSCBW5pk
tp9pbnYx/eqmjSKTIJa6acFCcocKLhWuF1wPZN8eTXJzHyiwC6hgeitM9zOC+as2
Ya8rDqpA8MGg0XLrGYMjw5YZvoB+aaKtXEpEQYyQN0IXN5dSRyudnlPg8s/EOa5+
679jzvD7FKsmb/Kb8e16qJgxPowpvBXR4h0/dlGTRduXuF4tnjDG20O9PmLhhBgr
1fz/Rb5yINfTRZog/yDU1h9T5H2DvVF89c0oxHlGRC8oXlF7HZLCIyCGGHBggc74
jVicRdyw1NRQ5k0ypGL+aMLo5yrUrLIMisjsqQS8YrO8DEfbm4bMEKjSLF4rla/m
WHsYaqIpkfFN9vkfLS0TtBXksiOVz9iQDYCaxk6xYeanqPZ3HiA0eNxgSDkSmfLu
N6XJDK4NZqrmM1pvddYbFWb+QJ40/AXH52Nx20Nnd6GlzsjxBKUWcBFRyC8fWO+j
yOZlDoCP0uUa+uOGiNvYFGAkbA14XLxY87mUci3uj/qjDHap+5wH0s53SQ9SAb3C
YO6ke/r9shH+Febw7FFYV4n1LyldxjzmnwyHy7VBGnzFXsYtBgDvWYy/U2ckTEAx
FLbpey9rpYLspmAWMuKMCLJHsr9PrhgPrgmpxaPMyMtxVFkRp8Sqv4nmFEm8BCmW
U82VZa+E6gwHV1kv+KT1PaoU8+Z7rHWXsy6qRHFJFB1zMUp/RlppDtOI6tPnKsXR
oUY8GU6DAcBWZv/AOqN2/KsqTitVe643mgvERCW2ipp1MA24UXjrcnauerKlrCTd
4O/UhVx31xwCo7FHEeCZ+L2UggVfM1EhxQ+238HDNkZdFkoRovC92BVPLPBDjiO0
y9Q6MST48rMGDSndTlVTGXm7V7RFrjE0FlWkUnAnwCY/nr9E+HgqqAKlJfEhFsuC
OmryrMcNXmLdmsxfxFseJ1gM4F6mFJDs9tkw+66PTW+n9O6uiSSVzOrDKbWoxsrq
eFsIf4jwoKXDvHTqSyTlxWpIHFhtyV3yTi4zgLlE4/vTnE7dHw+ChTyuI7X3hLKU
tB0MY/45OzXbNvUuY22Fa3f8ETdnia7tJ5J3z1lUjDqO7u6w5d3xTYoTXR9tq9to
PvH+MPDIj1WeuI9ZmE2EGuUly7PfbRUBj7iDU+VlxK9KmsoTjlfZGm2BcnoBttO2
S1BBwvuY8SnZfTIUEkN8av6bdbzT7bRqGlKsXXhhyIoySM2uekA1gzJ6OeCz/UBS
JHurVmsv/qFeLdMKqgce6kOX2pFrdkIW7L1D6Q3RytoSGhZm2pJzag5anSFMgz7v
REXGTqDxQlcqJQ7qM6LbSCzwdjLs0q5/OAlsvPCRJIBWkwaZ7HgMOKibYvOdpaq/
rdetz5KwV7BVr2z4gmbYyR2KiEoqBhzQRlxK6FO7q2PoczXU6en0d7TXtxWvg6JR
2V26/KdCXfXDpt82kOvfRnLk+qzFjBE2gArjZy2NTSocnysdiINqaMnclkuf8UVN
UeksbRSIqwrZxX2it1w7bb9om7XbHKtbtFE27zp093MiN6QBbCCM/W9TsJIp3FoK
JvdGYl+6PyPcxRZ3Dw+gfurYg43uFevP3gijz3TzMqzOyAQ6izI4M/7yLEwGhzeh
yeLpQbSsSObLH1oS0T7t2BpbIbWxik48L+cmCsrXc6IOoclR6z8TwS8P9gXDogT3
yIuV46NCFsD3nPpFIAb57AXimjojhJuZcHMQ5BooUBBBtGNmPibnwzoB8WrKQ8RB
utTpEgX5oMgKRuAdX1dY4Zg6vCg53nZ4x1R3Us3/jm+xVZEEvvYOBFTmUokBoK11
U9/g6enM78r/8hGNZ2P/Ieeh7RF12agfeWXAGrenVkdPg2koowsoKpLEe5FpwR1l
I8D+4xAax+Qw8KeIMKAUvBYUHvTIbwEnUymsLq7zShUkp5oOCrS0Q1PAN+GkNC+2
9LYJ6wPFyaud+cH53SHWWLz+9n9Yj4eYx/i3bAFzkDD/vW9MnKA6NqfwBrpJuNMO
Tv/TW5wAFv0tvXDSsFT3DgGzcfdT9FvdzozLfxrv0Hb36PaLP2U1crb0sJDeQ/ke
8n18WJAXpnFB2UEp/bBn3oW9/Jp66DWuIBe/laAa4r1Qfd2FPdoYDKzeHNKzkTBE
l0g73199u8sXv+LlDjgcNZojNJP3PTzciZbL1cuAEL11VIbed4Hg+NkJF81e2pLB
3+pQJUgt2OwyzuDJFMP8tSgD7ozrhH3MgV0CH/YP20r/A2e+v8msdxO0LBCCgFW+
SrdfflH7WdpwVQ8leYJ+dqEdmClWb1fFAgywxKiJROmnN5rZs3Tb02JxT34Lyj4l
SJv76HDAqmG4OPKwKR6vBc6AjY1fWrwocnnfxa93b4ZNUfZdPYgBC08sOHAJ8JQ8
/iibZKK1CzAniMICUjVz6EL3Vvh8RTBS6KsD5nOJ8lOForSydoIvHctCqi1neSkg
jkHuo0KcjagUKUEr6fh2Tc3xPRD8jSZz7WOfE7SAKWyC8XnOMBgrmfqtIMetDXi+
Lt058r3psqjiPdU67SJbcaYIIz3Z8R6Mqk/HgoPeA8NLurljU6YC5gn81j8bSSIO
wUuKqpakpVFZhI14Bksp6vjijxeRf2WFsvqNFq7/Z3YPxmXK4QaJ6d8vkK9KwnTJ
6SnL3QuzBU3Se47Jv2J3lJiRZiqlqrbraTsYGaZoF2rDvt9wHKObcw+B3HWEOTlT
bp/OhqnWtEQpakFYeP/xfLI63aAVQM/Jugz5/yPwcd6AEBHz3pww1nudK1rUX19l
RH9d9lLIFy+cjG6If00YwRYsZooJ1sqL+Ir8U0QKWKcg826jSUY+DVW7eNoIHr1g
LyipUqQo/4b6APMbX+B72Uu6GHnLbu1NgUsNa4/+Amsez1iK2AWOOhY+d1E9w4s0
h954r9RkbjRotxlIFZUflZNzoqgqWqA+wHIGvXMNbs1hI3CJq2nnb0DzdBjiZbXj
kEu9hf8hsLX1nmPK+h7GAVKe5/nLTL7/WuQC35mVNzREeSfbMoYC+PsLpApHw7hc
zlzHmYAyCse8kMuvi5KwU16TRk6OM9tDbO4+A649nWyU+oUPtAWf8u1KFK42R7Ot
x1rF9pabip+CpbP7d0FAdToz6IfK4csDTK3tUJKsIcz9rIDCmEvWA8LT6b/3GBpc
C8/PU/lYoLfO0vRv+8JspFdBvaS1GMbMu4DB4ZlecgAriWJFMy+e0r4cVN8EymH9
7Ecy4YWh8pX1G1G3pssbFubxhosJ8HsbCWaTpUcIU0eeX15TcvriTev9YYayzL0f
BXg4kFepswZZE6tAnlzrPBLrQC8DP1Wf1b290gyaTXu2hxv1mNOU3ZIub4WBZsge
D/WrOAGvHKURDOY83LjCVwwE0Rl4kg/OqTTvB16w/NhoLPMnj/vgLMERklhGq1Sw
o93rgp6l21+rnG+YOSfew8/fLxHjheZJn6bFOwWE614x9NUxKC/5mO5EaYAJQmt+
AekDVosxW4jGDl4xi2zYMWeT08yyXxoGOMY4bJlMJLgZD12Vx/jb4+HMyBTH/XXl
hRwi1bzkzs+7EH/gwsI5Fw+hvkI8vY+Nys49dlX16XzaIrj0DnvDB9JdWtelwTcy
kKD4GSagObikgnS5qF2FpUdgdwYED+UKFwsCjhUHs1mV3JODS0UZi0zhWBMeMZjV
oNuD7TUIM+12GpnXfXVszvH0o5cyfT/6NwwQ/Avo9Us/4D/7ECrb/K8P5ZWutkcN
qBtvAloXoTOeJB2qOTAAktc8BNbusyZSkzwIasky9tey8suQU/lh0cqjP8bwBthx
9mTIGlAEv/XKYgxOmkJNyH3nH3nBl/fV3tL918qGVkZGwqDrl0tvNNDCMyoaOrie
XrLBAwyLZE5StAecmGQ2Wu2s46/jH+s50V1mrVQGkyzegz//zZqdN5FTUw/iclu7
4fCXJNgBlLP/ekHweWyGoeaM8yvPaeiVYaDLec+xp7ewtYEIz75XCO12oAepHFyL
GdWc2ermVu1Sz43tWxg84uFiQokGvxlfiT3ngmcL2AMpnQBVuxKCYAeMW4uNFPp0
iLIO+ElFDyb77g6GsC7nUblr5Z1Q89t3m/75cmK3HM8sBaRO8PIVCwNHRtIMWbQU
6MuZcXCr4pQh2BZM8LCKYqxtsfMSwS8RXFDGFu+NucsNlVysLlCWfZ5H/OJynUii
sUmbuj7K4A1xjV07vOBIk9aeDjkj+ksNCae50rTKXSR013x21UzH9+79MleeWWfY
xD27RXu9Lcjaa8OWQ499yMA1oI97jusaJHjSGvB9dNMctjo4xddgWp2Yx5uiDVEa
mq6e6rtkQ9n/wzUh6J+LHfqpgferoQJLEjjFpRq+nFUEyP5uPfVroObbaRykdSqF
YyTICzxO1djef3T2pueWknJKYKilH60P+upVV+csbWgJLnBnfXyyX74tAJI0iwth
yEOkVCY3PFTfAwnaTGroKqB9Ik9P//1EZGV7PmHCyHj7g6U8L7yvcGalUZNoSGfu
7E/mXpJXEY4E61nIBqGjyZSKuBTwtTsUizOeFjCiBxF3whpxMWnAkh19Qd1tsfMZ
GqhONCavha0yaNlE0c9/msi/K2jYTRuWH3Jto2q8MDI6Qbx+wn0JetRyIrIwLm0i
Ast30lRlsBo0/Pu/nMiCudVHVxZBpptaW4QjTMDcpEy8ACj3V1+tjbEbDrqyGLe/
Lb6C79nVrP/yBmYEn6D3JXXqcUi9OHrHmS3XO8OopxJBQxduiChdPaivgzEdY3Ek
09FfyN0Ng7ZTCTApCyq8BPdUMBHiLP5izfmShsgbVdyt3Lhqk92gEM80gLAZmzfR
+IJ2e1yfav7Qq6r+GVvotHShi+E5zami5o5xg0+36F6TS2++SlpWgoRopzHqvQNy
9WKebwvzB2nC2Ohpm1BMZMHgWhqyOpEGE4+o/A+LCfoFRl9mtnxIaMFYHRknZjk+
gG/uxY/FeO0muE5iaarWhgFLlJV+BpKm/ziWabjeDF4G7kMgVcx1Kb5CuWIylIr5
Aomv5mLeo//gMShzAjz1gvR9KJh5301K6En7zcQyxgOWFBb4UH5OHki1BIrcIpzZ
M3RotF0aCptvLL4DE2UqEPkG37Z3540yx6VAe+XAyA6dapgcpn9qmrocf4HQsdqc
tWb1WlSJ+GRj2FoIBOMjogSYhALwng54QAM8cT21GpzD+9LC6Xjb7UsU0rAb5yhO
GCVsAQBLX346Q5OilDepNJsRKyT+1RTa0RNTPjRKdZtEew9iT1kyeyQFfbP6lGa7
QEJs8gFFeVYO+c7XsQBhNIsHaGkEt3192VRkrNNEVJfjHFGE8jGzrFgtGHGaDB9Y
+3iep3l28Y/WvH6R27PgbHOWJoqLpgxQ8xuXzRnyJY2k2w7GuX55Yire2JAYR820
6AtDS0VtU3CnnmD9l1Guxx0tmD5FQBed5N/lke5Navd3sIXz0HGufc9dLC5zHwZa
VR45ke4ADZa08J3W8WW6B6uY5jq+5ohxmXueae7eP9ry1Jqhouv5XnyVf08pEAPl
JW1doOh/GNF6BcT4ib+LIx9ebv1SjihsL5nufM1WSGgSXo11A7Ez5+RxMX7reOAb
teOwnTU4aexrLiaBrHQBAlXK9HuCWU95F8zsgrRDzVzUzueTomCYAOG1T61w/29g
7KqROzc/3paFOtn0aeWWCpsuG6XOcEdm8BuflbHbAFlvK18WUM3y6KJKcUo+WA5+
JfSj6PqNFOq906zLdEc/kMDbJxE6t6I0X6jEdRrsw1oYRk3cIZiHDzSo4dwd+MvC
gxwO01Gv4gZRbXO1EdtnMREQ3oM9lBaIH82YC+9OFQk0NXxGnk5R9DEGBT6jRIUk
gyRYAAZxkXoXQAEbqq+KJA5z0sJ0l50HLkj1ZITLhOayyHkFWmhkhp7zi4uApaK2
hbvaSMnEwmws8EsOkKzS4x6hM2frnJp0c2o4c7ddAtCJhnIxRpbNbF+i9ucLrl39
yQKoo9ARyA4g0yQAC+dSYceAJKDOvILCjTG0v7oWfp48Q/EjpdVz4RzFpfw7MsCY
8kaqr9+kGMuNVzCXE+Gib1fX+uDPzRwHmeWEUE2otPkEtqQAsPOI0lCZgfRUtS0m
gMneKJFR2AJCVglfOU6NG3FH+uHhD0QCxa7jWCXsiiq+XAzyAgkLy/AOojbdXdnV
yI9lVA1faC2Gv4v8LMzbr0e7tPgfMdkpvcBXi3ZB2Ty6evu0wdCfvBjHrCQvQpeV
6DrZjBWv1gCrBfkuYZF1K4EG0GNMX0Wc9zJCXTbL8BfhEk7a2AQo/DJaDgQnTT/x
8YJGrjUPtc7hEEiqnewIxksCCQ7sbTmxF1ff92r97VOAMyF7uSsMz7LirUV92sHc
aKrG2ltFvrb1rnJUAKOh9nJkzYEO2y+6Nbiq33mWgAmpOH2jAw1rO09/Mj/GQFMm
0vx88+tCra9/IH2P9mNbE9iEnLvDGRMgeGuS/m9UGe4D3cFg13mhIkqhP4GLzZhK
g3L6MBK4L7dE/tS6ppTGmBYtobx6EibQ6VqFQKY2u/0zBYG28XjilkcHJN91i3EG
0zENzPO3bAkFhWaUHdonqRrjTm4/Oe+3oldg9JARjK5StdUhBxV4mLVcvHwwDn0J
wWp9KJTExdfdADrtSsxxZObIJuPCPnGb/9M/nlCRxT2DCUy6dZ+HzTrJncAhYKvq
ed2qLP0rO+vLLE/ityCFUzSmVKDKnfa/H4C3ooU+47oySekTvLdIXPndQbSVH5TO
x94pEeeXPacFG83+LrEjdHqcD8ungTZQPWPfGsMngwPwGNFTLICzz1zjUf5KhOf+
udVcI9GO16taH4Y03z0UhHEsn/8bobLvDGYJrQpD75Zirg2k1/vdkTgBiye16MAa
lGkZF6LJs6nUPYAjZmdxa01wwWRj5ZR8VRKyjUIy8k5VVeH8tFCQZafMAQK8J1L6
MUs6Xx4EkcV2BHvDtPi0iwTMP/r+jPCj/dnhSu8ylJANkib6o4MKYgeZtRGeYYGU
sEpVDdm5NM5VTH61Kz0jQO2Ir3vaJtn99GvFf798cR3K8RWvBnpnB1J3JU7lL/am
QrpFEEQo7mInpMLQWkafRc0U0OaL6ZPz1Jc6KjAE9lzfSIebuInO6IvekBce/Ggj
sdJ4ANbCPzT+IlgErDGuZBXnkVs9uudlnrQY+uar5tOwlAliVrSivyxKp6anVUMf
M1eVX2cJSpCfrhvn6I4u9bJXJSSJElLsEFLVDCKzmfhxXft1Z8en9yNUrLLc4prl
wo+65/99g47eO+QLSkiUaHker5QwN9NpCELHz5Y4PUf67gddiY3ms/weBNrLH632
kzGxgAtv4UpAOwaCwcCp7PU8bCFxZGRTpBReopJIVca3r25rTI8HcEIc06O+p8li
DxcsEyPbX0PBxiyCSe/2UnYnPK5dAwulapUWJ+y42bAoKTbVeHDKywvkBymcQB+k
oM/8SlEbmHs4aB13B/AoRBDF6ZalwVulge6XIgcrNB3IoS1CDFf/AIOiezEW12l7
/o+TccDOAdzlmg4vaj2gupuSMz64EgaVgtPv3UVXRNmRfs6TLD493wie1cvbRI6H
YPC30ImfX1Ss+iPfuRjjr+bvxVw91miPr3PZq7EFexxXxC5ExFvyafvgb34tSdfN
Lz2o73jueo6Qy5mCwC5fpcsncqUELQ0/NyQ8sEbEbHe0U/4m5Io/MjQWJuUvhdsA
u8WStG9vkFYQQMlT8oYoylLib75JZQch1UlhcQOFf63Re2znjYk07Q6TbHbRTosf
AWK6wtuv527CRMtXqomQpEkEo57joBqiMUCqi0Y5hbjXPoJcD55Vg466GL3FjzM5
v3q35ZaYwhSBJWZIAI73RnYbUTaNVyiGxlTHwQd+BGQDo7ZsXxFvkDbESYA7h4cx
SWsvygejvgZCvqP1iPMKAEJImjbuSg9rvk1EE7IrkIKecz/b8iDDl2ZkfC6XFDQt
5qKMVq87e1SWRuuuNrRdVClYRWhrUNFq3awv7JclY0NyCySCXu4Yh28skMFEQPly
pKE//ixQl1GMMhffj5BVelu9xEQj1M4mvym/lE8xVrgpHtz8Dx3lWc+DdnoevJ4T
rUbPprsv0Xm+gj59k4B78k5KKw5sGY/U5M2W72qDR+5ypBEac27xjMsBvtA+RV0R
H4jHuyH4H/RJu5uvkH9nSIg7i8oVuoWyYeHBcMtNWCAGGLPb2s5E//mqdW+MIMPh
OZ7mmDZcOjJKpN1rFsjFl1ofm57Z4Zw3QYjWBGwO1GuuTVpaNQPnj/lMhBk5LeD+
OWSXT4lfqZlmZXdUGzWp/HaYBbwJnj8HFdtieH1A/FhrT/83TOftoxcbV3qE18/G
PnBpzNaxAHovIooL5TA/GWFchMrJzv2O4hTof6dnXcyeiptkKgcHFxY3UAEW/7ik
D5V36LnafmO6kOnbJZeKJOa8Yuhausu55lHGqaEB84LFgBfeOPWlzhKL8c6HmFvb
cTfnYrIZeOU292JoW1DiFiKz1wzzOUZgXPdKsiTS9n2+oQD+7g8lRzi11I+P1mac
hjnjP8+MZ4T57vErleCFnLh2E94Qcc5TPD5cj6r1bSMxtrywJw7vNhNtfS2FYdZk
leQ6Oz1KkWHG6qJIhnoXr1blGJnuQndOm8McmBbeiRfGrzsWPvxSsGpUgIZRk/CJ
QD78Gt2pBdW3hTV1YWq5AJD2dVAYOVSY53nWlxBWjBCFoVyf4ZID8pDt9qNRXJjT
sc0RW2xLCjK+EkuQVo0EJV/8YNP4XT6izZIW9M4x+VzHvEAkbPvPExOAO4ommZCD
j/xNFdiU121mbfOaiZHcFW0cA4KCRFMAO9Bcz720oJYqfX8e3pca4MLH3HYonWln
U3K5eTGF65sz3TRbKAlLHQ1fn2xrbhZJbw94xVELdyppcb3HCJ2giHLhl7jpqxnT
CRsxdAzuQlvD7xXin2Rn28yihPcWj59KrpR7FK9iRach5Fpf4cjk5GjyqjanZmr2
3ksprfqUS2MLYx1ADt3K2ocOPO/xlS5r7xO2liNtakXXsSZH1Z4ROdvTPyYMZT3M
41N79VR77iCqZWrrxRCGiu3jQDTvq9f2igyl6k+m2BPfD5HmDjVywIBfWxG4u6mj
wrbVdIXE5gk6HWVueDseE/2MfkB8briJnWW0MlrxuupOP20mqwfUI/fbl714osEt
riFexBP1suZW7u/gUS6k+tjwxO97dDzgYpKqV+UQCELXIYV0YRdUQpWJ4M8N4S3Y
brIkG7mI2X1lL1fXdZBSkoI58XVChTnbLLmlUK2lw53qhUD+pZM1WJJKrwDRZ/DX
xbeo2vekUpsoKGflfAFlfb1u0dAhFKPvLRpkJLYJtzwASMfWZD56gJ9LyaFQAHhp
spQHlNvTJpjVqFeOIroU6gRgmTEO2mCNCJXogqs92u5LCyolPah2ZEwa4ZiKCiEB
DyV5T1bhnLNYqCEOPqr4FVIZWRYcZwkln+8xi0J8bMTHG+sCsdzN4SMiSaK2/cvs
WquvqejxtB2qh0hQF0lthLFQmz7WST1Q9qaXCA9CzvOTf7K9TjAjTMIA96uia5Co
ImjgiOjlzKx6Xv4GTejnFJGDe+zgf7lHHO+ibaUqqg9QgDh4/VGz6havyXyA9CHo
sIle+veLpywTf/NhYdWbcHCOtx2JSNhlqYa7holMoUSMIn7orCZmQfYJJ1TTVKN5
hWvmoHcjLcuWARSAmICd2KEN17otatBiORnsSr8EKKIToDXCm1o5noXjPkTIhXQA
+1G62PcN2raYicLgt/B1lQ5q7CwCCdQoj3HazElaM/zgg2LnjMY63U0M/irMU1Pn
gqL7cMVD7Sb68+NxKbnC7lym6c80zeAmQvMUhsAy/DjhjGlEg1dwmiYENH6WvmDI
`protect END_PROTECTED
