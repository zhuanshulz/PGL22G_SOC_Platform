`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0FNhzziSF4z/R3X7MyHv35uOJMLnzTw8Uxl+q/4EickaM2lZ5ueFqTdqjZtYfvst
JZIwn/i7WF5plriatLLKGvvQEGewYzVWIPkN6EHlTJ5BjwS/SMoynWfcEnCDsczw
6HHTPkuzK9dQ4+HH3qsWDWtsRo3VqnSuKZ63+iTnZWUj+FJ1wCn0ASuqv/lMUxys
3ky2NlDQkxgMdjuQYPTXcuF7bC546SyZqNp7BRMXyNdMlqQhFxyAnacWDtLRnVn8
sE8md9UayIhhJIa0u80SHEaZCp9klWeexWUe+1M9v6R9CTbb+T4QiWAXplathvY3
Q4wZf9bXVrW8uhRdNKcdGdEXhe9iLJM0uaUAPNRXXYyZIOQIivDJ55yHi8OONcvw
Jf+VSb8sMupWk5xM6nA5jM1Yu2cqtJUkuPg2FzWtMMGu9L2FX7+gv9nacRSuLFDK
Io43INfaOu3K0xC7+WX6ROMiQx8j05Csc1iwkGtemqkVoQg672Qq3Gsu071p0kRU
0Hey+IrglVR0C9pHEBuF40WUzn2HYW8h/9s6p4Dy1sw9DgRUK+1eDhI2PuCNW16u
2DliTugvQTPKdvlJH3j3lxq4GkcmvpypiTp06dtHN7vhnTX2Zk3iEbwtflhc0zT3
yYyvkn3mqZrLHY2Qc4/PZNCNsLT/O+HsafQ8hcqhUZEYD0KSNR1Ss757Nrtj+2y3
GNRgC76gMLekdnDfjJyRczaMVRRCBoC04Xf3+ONoJhkA1YBmlrhxrj4H6z8C6Va4
QA6eTtH5CzIN0cgU5Eaju+sW3hR3npWG5HOo9/+CLaep9eUe3IRluY2c2FW16Qff
z9ZWpLytsagBMbRCq8Cj7LAoKTJsXooCPlATGwXtXQi2tREVTpjJ4mbVD8rFTAbq
NgOFocQLDvSWkk7LTKIQlgx98Tp9t6ZJ9IkqwGr7D09h7aaKtNXcp1zrTPjAJ1df
rx3CKXevgj3G/ZBBLp/9T29b8EWHbsHhSahG8rplH36Qv4FfMsS4DHjEMvQWROuR
IqQ7jnVhuVhWRk5pDrE8fjIatyLdLsoi0iPcUrbmUxOZOCoHzfOz1iYtvH96mAlQ
D6BlUXMqTh1tBEc5lU8MBhI/td0JucXI2KriDwHIEkyPHw3jCMNg6zJMvCPkrUJt
URb8n0nPJe9fly9BM/x22KOsEgu9nHpEi7uS/0ZUE3wcEK5oQ6hM6+mbQzfZyzta
hKrDaCkCNNIhxyFrjCzWxV08FfUAzrbq78sRk6XaaiPFpm0YPQs6EKR4r6x7IDh3
VfIHpckWzG02FcWM+L7vw4BsxUBYcUPPxVCK6yevIrxX5U0+QIzLI7tA5/gj8psQ
V5uIn/bUt/WNM1ccrYbbuGcUn9H3pPtI1Fju7NPxQsB1bHM24AtJkrL4OysNNEeb
uv/uWSjnIb4mKjS3JOoyjURv3LjZmxCneJGtAqqxN/eX37PG3A3rXCsESb8tCiRL
tHYLWFAUYemIRTeqoz1CXr5G6CpNSKvgeiFIRO/m6B7dx2GziDW9Xs/OEMLH+agA
lCmdNw3cqCCsi0H122Rxyu6BObeV/9raa3wcTv+yYydfi9A9oh6q+dhUXgmCxRe/
BZ8TYQlHFVsblCVMX982Hc65ODFHFLSsm+c/92XTQRD1i8oOuT+sCcCsuu4bAbzD
ifopsFdbRWuBcVZpnn71EeaSDucJfUOmb5Ox/P4xoW9QygaTDqnrPnkSmgw+8Bo5
U7zY27shNpYYBURu4jCYrBNTmoeHm5V/lTUbR2RVTJDVmLsF44XNp6KiWycNppab
FG9PcGAAq0Q/ZaYfqLcV8pOmqp9DnOBaPCOtvjltKDjEB1yHmMtQyP4LsVrpadJK
amdtfXzj9u/zYfzxbJwPEwzSSwzPWZgePx2y/w4l+noD7br9dREFQ+64dpGM10OL
huXEyFkoqQs7i9LzMAG303O7f92G86IKETUna40sybkzDbsfQEnANe9Bt545KOWf
r68MIx8bhvVhu1vza8fQz85CEV9aI2QVvdEx6RRVnwbPSDWXauXuyt71rVIv/lPH
pexYiIqWZ1ED4HUKl4IFG5RX36+BLPBPWohM7YC7Tz2TECvsuG+jA4ADFJqURr+i
gpg6hpAG/fUpazMyFnInUSd2TxZjCKFX4Llj1CbBjNxofPJTKRhl+8XrLsEpO8VC
6GnB+kttJyBu+vM/Y8wATKMOy7WrPlTXFHAqKBCDGzAAIE4HG0yANUNzl7eAD4rl
IDVLmrI9NU0wnz1DxmfZ6bzq7qxhul/mkW/vVfnUOuZ6B7ycFaGi5dYuhz3sH1Cw
qHeIyMf+qqdYqZyyeze5PZeBgfjL7zadsL4ElmCsSSvCzjt/VOjKgvjI1MmVCKRq
dKtlOl4Zrco5W1IMvnXYqsVDEJCqLer22URGiY+dL1Bbzv13clwYpzk6xl/roraI
GHcSFnBcwBTE6ZejgZDaX0KJzJ5Ls1mD3xzyd4NWc8Qp5jxCbEiWPWdY90MwwUXi
K3CEuuIdw7TUQesKQvHtDw3YLnwhW2aDPfgWFCwTR2bvf2WFHQSddrT1v/m6VSKI
`protect END_PROTECTED
