`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
djF/orXruHSRw/xp03UA1HPnHq2lEU5D4ORJE0Uai6OUpbarBRhCJjEc/FhqJ6L3
Z+tXFHWDHSJHrudhS0QZF33P7pkdHlXwx8Jyr9p77qcClrl45z69kJcFBJLLr7Q+
IPXTgnZDsZsGhzTpYZWblJrjWc+TJ8wWi9IO0Mpj9f6mwQyr5GAcVgTKnjg0N10j
HrXTE3pJQurivtqzKM+Dm7xcHOhGw5aDssh6wxmDMetfJFRIXTOyTR24/kY+wqmB
LKTEa85WI2lF1XXE7/Zd3y1o7B4PE+u60NmamWHShxwuVquhzPQ0IaaNi/Sgra8v
hw8OJgseDXBZ7EgXawJknx4eO72wARK9ik+5NKdxa4Z10wWSdcHMlB84aq6xqKwb
7dnGXCnS00ABeeZCFK5vJlJpaacTQtSACnqopnM7g5uMuhqxYyKR8+ULnrWzHRfp
I4fSISMW6inIio051o0zPtQUEZPycNzqipI4Dp+RYRA9oIeWO6TbFya9O3FVrPvn
Ork+n1eKMEDGH4vMzZH5+sHfp0HwavdFAQr2NXCSRlMKfFXRjxssMqUo+Ak/6hgu
KHeuP4Y5m+j1CE+BZx+QePhkxJ5O5aOArHGg1oylwq1n8kSoDF42o+1APWe/3uqd
`protect END_PROTECTED
