`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CiXdJN92FoBVFDTl3kwLpbCUPoU2NnCVzR+f2NmyODGvdu5xI2/kriCPypv5rFdw
GMkbgsyayJ7ALtrE/1vXm4fp1QHNyVvXZvI4Gv6UkcRjDuppN2ovlvB/mpBgWktb
SiISn9/UEWWKHJaYOwa4dzWpYlwqlNPnKt/V/VzLyqaJqsO8G/hLNpWbiStIpjF3
wutS2dd68mAVf8WlbI0m23lDNiXTk0AYGddpm+wd3s9lPjs9dO7ImSdBNP63eHQI
/L2WgObyhQyXP09n0F//Fujt2xPMJvzwlHsf0tVUx4HDcJ8i+Nnreq6PrY1ToJyV
YZwE618NBYQDqP4btfMoJm8XsHW1OozU+CRv2JRE/w1EV3rDH2KpUmlk82eBk7Dl
cIv/v8BbUUrEPxdD//essB2cYoQQSl3E1T7cFjbIMosHjtigeFt2UakorjUGtmxR
19c8GoLbTWSxiHTNbzrYFW9+hQankiwvkkX8YtEt2QvgPTI67rphZGcr3ZkhsedY
U2TPrRefy5H5BV5L+Bs3RpCTOiIruTauihe+n6ng4EquE1u67L4AcpjGVJ9SA9Cn
fMOwJb91WjFkNh/Ee+KkmlQnmCr/fZQKURjzBDApsFIuYOQ3drXY/5t772Eb9QtT
wVQff17VubpiISZCoRVLQNYfm7E9FblTme1Ausg5FuSuigj/tMlmxyv1ZTt4h1IJ
Enrf61xxVXp8dDxTfwCU2FtpdhStE2/Tdr0W+89O6N9597G0q20GJtQc0es/t/id
iUG7rBWxo5hdOVsf+SEnlqBEI4tLF8yNHGmRXWv4R5/8rxVt9DUkLPr9nUPPjnEg
AOCjr+Vpv798VbbeghFXyq5KN6ca+ohYDO8Wnpm/1cIFrzhmDU1y38J6o24LHZLy
AE4cAgbKJ0Di4+knawRR6k9hXcSBdmE8PMUGQq0oZwM6x05sKuE1v+akh+P3ZUip
FzpLSsdF1l+yNT2B7sHWVtOIW4IlJagVt/slND2DiVnDit8EC8PyzcC8ruEHqmT8
QANkYW/2Wuu1v55zZKr3yU0vSvQB/I5iQmjGHSw18JGGYEuwPDOtLkfPu6w93ZLU
oZ3t/w3lSAeogKUX9Ur7iQr8U897bMvcCalsmke/hAvEjLYGGrSTVZuPyUnrr3li
+ixUgz5r5yJvXQ4702oqoGRBMATrxCp7zqaeFBWnQ+foBaCq8WGyBBOcl/yOmiak
SCtRaJuLMH4BZrk19K+FBXczdEBDBP1SujipAOxdb9Ryn30dYjbi8YSN61OJ7gcs
kf+01GkfF9q+7BO3/ezQoSH5w5CXl4K2TFZ0PbQCAEbNU0sXu0rzKEiFdpBAm0hv
36EHmt0k5KbHAvgPhZmESw==
`protect END_PROTECTED
