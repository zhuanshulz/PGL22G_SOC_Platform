`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iqCnsIVXc3KhZkDoc1Qzm+lACRiOnCgXZKEU8OOvM0DwCjMcpLu5bau46zZxnLP8
uuzEOgwW8LBgYol67wI46axAgLoZ0B/MR6pXsKxas25q+8fSNnCuPcmN1o61AQQ8
S8PUw+N3uVP8DFuIHYilfGuun2+g2hAFKEdf+Hka7v7l/eHhA4Tk+nIhOubaxcga
yxguvFmfXPE+hYiJ95XeFjEOpXdE13BL+KvfW9wBw5uKbcdjas8cg0uTLCI1vbox
x9LgBBRK8ihTWsEyRtX1v782/2JJbqA1S3DyEy0ey8sWrRDwXVY0UZQe2F/83ARg
E1lOsJlENkw+A+Ln66EwhnRugsgp8H2PLvwYGPSSQj22MmPjMxczs0zDK4vRdS+y
TZeBLelBVSVZ1tqt68OnY3Xzu7x925zKgFTLzKcVkFPzamucTvuMoPMrnK/lfu3t
M9a67BylERBA2vihFfYXaZEM/3EQjsQATN8Nuy9vpGTd6PDe8NhABs/idVuvLnY1
jB/WGmhQjKJhsCi5V5RqLyvQR116PYrz7MvNqUFlg3qVljpxWDXMg+v3JBv/a7hq
yMGRaqCDmcEV8gAf5zw5upHsVMClPopVxrhgW1zAQjiWMUU61FNXqSDte/z6Mua7
CrlOhkSwMEyQjEHnQQmQMOKVf54GJ9VuDWD4ap2JBsuB2eMuoCxStLg56OkVckEn
/PvOEa1sdoo6XAGNs/CC6VzL0OfhXoMUA9nCLeAm+X3SDrSExfmxJ2n/0AbDPAPl
Gwr/RkueyQNw6gT4spE+wBpq6qwBEtguWY2GuC5lK7sa1VdcsHdN3GR5LBS9m/y9
PqENEksyhG/AnFCcwshRKwzFfF7u4dvowfDiYeT+Tb4/5rgyQU7RKsXSUWWpsqnA
PbSfDzgG1oS9LzvSy6UboA6GJa1WvyxxTWOmHr8WQLBVITwmL28eCviLCUnh3f+K
29KYI1vqN81t/NoeISPHTeaQyqXqcxO4qVnVmA2LBwjEM0WYE9IcYlaL377Lsdw/
Y4+OKVRhCsZt15uU3IRVmeIaDA7jBHZZFc3l1t6b/GJrdw9KNTUUwPufWrdSDRWD
sLtICLicV/ngtVK0T5LARkOFMsotn1fOurc66tIvB9U86bB7ddyaris3EMhIKvik
JWWm1CsLsHbFWKLUJaBP0OUlsMETx649VhL9wzCQe59ekNf3mAgOga1rLqHpD7hv
cH2K2/RqmwPmV7gEyeG+xj/h9Y/XS6DkwUOEY3z0tpEhsMQgfZyc/ssqXAKYxCQ9
Lbl1/TIz5uQBG7lX2FZJr/pdHh+V1xKdVDeu3vaMrMg9hpaATsFBzra/qvWUgpTX
LJ/GovsH3nXKVle/uEjqHpdaG5Zxt0U+N7tHuAYm4okR4DrmPc2UgSG5/FoEK95k
CcXV4le8Kh9AltQVz47IgG8PtPtBsKhwnscWk5xAhJnKa04iNC10N0QX/nG+EpNI
qLvUKXJgMIkEKqIBVJr9LQCWyaZQn5UWGWUYCwANN+0RY69FSemF+f42GXjjK1/r
QQFcGRRw7d8Ls3FoZhxJfm7g90UG7YlmCctPpiVsvqn78JgCuPGlSHMJBNwHl1s6
NT5h7KWFLHEmVVmTp2gF1eBtpOSIfgi5XMBUAHgete7hQzyfB4BKnKoqeLB9V+7C
FY/KGb3rGDa+qZ6O6o3qDKUkPcI17kPokmrd9BR4TvgA8vfHJEGmB4bVaByVO/fr
aojTRUAJtkvZddbq5hhaqHnPoKgKubLyofet9QR6uqqPYGjXslE50vCiMu13RCSR
Jt1Li9aPyVg5FEKQKCXhx16z2WMrc6JVWkkMucn9oNvRSQprGe3SuX3/DSQ97lES
oavt27j21SL5RT7IFTJMa0A9kBYm9VsVR2Jmon88uf2gUsbsWP929wpM93P6Iw2o
EQenVLnedLXZPxvJC2qaNcQzpw0/eamMBHTT1V1xn4N5PBhYyewlJ/IaSbbUQLu9
GwbrUy/rQfvswB6rg3exd2L7h1MricOfI2fqawMjLJVwi2jtAkOJ9HNs2qOEuoOv
LTeLIr7780f1N3SruMSjDbMTicKl7xGw5FHHj3vKCd9yM40/EwbYcSG1oebQpgwN
++uefQKgAznCmWqJMCHsn8077xmnKcbiP5na7KP8gelzEx4slDKYD6q6YUG0jOva
kwKY45gClXkLiWyqcoI0tpMWMuFVp2CuvhAWHpqANarRtvqrRKvn/pAYpESOkAKh
b9f+OxXvGAtlFJgEYayCR8gcuShnNb+SXw7vqVEw/vLNysg+adQa0gy1+9zmhUSM
0YI+cWkTIoaedPiDXGoT0V25CxqmnGO+7CCkxZvHRTACPiy4/Z7WH++bELFva84R
ES5USlyOyKdvXPotA1IqIiYxnGGYuwpmJwOBJKuJ1mtKn3x+iPWfnni8yRhvTYXE
Ea1i3byyjeIPkMIvGQn8wuCEoo+FAeqZ8hvh+RDmujE4JSxFAl5d5koC5p0nS6BQ
iTJYce0DOyX7RYyNpMCQE25GxKGuHbqHOhkGa1OrxWQ4PZ2wDzqwFyTpiBVn7jxX
7Hi8MqsB/EZ6L8VTVU7jREIYUjw8nJzq09qKk5ksJddPzVj/2lD7Z9s9Y8wfnuyS
+Kink0BjVMh6XZbrQiv5QJEDkxA1gCI6KEZnf8QXKk0CQmARTreA2KDDy1w3jl/J
8FfH8tM87f+DLxqjhi/6cB9GLIdUtWIgYhRDFWG8i24b+HGJ5dSb13Ko3IVnqUeF
ALZEW41T5OTgj2r+V8OI44ATiExSo4eJO4xPnndNMxlG1xQuAA5SGK5y35qo6Zkv
375l6GMKb6IB7pIEm5zgdhfrwn/sGaQKcDG2FcghOjUJAChI9uAwURlzLaKNjo1G
qKT6+NbxEKtlnDE7PRcbJva8Tr0NPrBDCnhPD9dmZtB8F2QI6RznrI2oHYRKA+ZD
Ax0RXSVJbUnlS4IoJNMKrTGkEkslS+Akbh+C3zRycaNzmHFERfdNp1tV5sWIcvBq
+5853HmPdIK3+7LaUDkgQRvOoLzaS4J0PCYjy3RrendK3MIUiTBgh0zIPlXKi7rd
ew9zvVdYx49eprKcbiWJfeXhi8crNNeSteTCjwjcdPLi6G3ujP9j8G60pdoIY4rL
PDM3A/XlUoykF3+h7Odkdq1N3InoHNqwQpCYCv88Pm10A728lrZ7n6EC5xzxJDDU
cjpoh/O8hM4LlaVt/sVLBE4TN4bam+ZsJfreP8NCwrg4s72H07T95lSveribCAg2
V66+FkTrS9ZU4os4kO09AII3KrWnUTKn00lMW1aPpO7jWlsHM5dvxz4UzGynCYyX
F5Y5hOY0LFNU/+hmOsgjmpmW5YJIQmB7T9zXJ0whGBWWruaDLCLPPqJ0Dw10kaVg
CGiVIZDmwkyJhYma0YRlttJ7SS1E2RFIkj78+iv3TRNUcXbpgMMqf3aKwF0ZhynR
7YOzz7gncTa52T43smZeN0Ie7lyJXyBHeTjTuS93GOBkqpdktEfYdkH38rBtc8WS
Moa4ZsuIQlSGyCuGVg60PI/fHdjBim2d2VX6NZ17TeqRUKZbSf/wOqGTkEHB1aKe
ktF8ugi2/7hL7FgDi3+9DL+908qcCuxcacWn89L4hn53U6rUKYgTlPqAoRaqnNyS
wKjgwoze3nBCs+bBvQGObgKsrMt6KW+FQGqpcR8lqQ2to8HcWMslDY8fcq38+Yiw
uWVftfAD7+/0bjQ0UO1EPzLdwmG5pr8uxmu1O6bpKxbGclLYDeHw1jMFFgcfA+x8
73hgtrVR/PKjouEJSxlq9kXsvC/U43ehR+Uoc6/1L2nXlYVi++q/4xK9mgqknz73
GLYuzCl0CQJSLk1PFQ47LpUcI8oBhGKNo3SyxJjp5lqNhpQ9su5aUhrQeAn9spgJ
40uOfYd54wQoLerNLGzfeT3ywqybev2Sxh2tU84Bd5tO+9Mn3wFJZWlDUlcVan/G
oAznw4/+AOPaKI46lO+g1dXDhkqt0eyUkEGlwZlQYj6RHWANEFEGjljLar+5bi0p
D+/4haG8jMy+nLC7M9xS51QIZKTZSGAOusXmDISUnaEkCyH4HYM/vNEbuvxfuq8v
dTi9Ca7i016b2RPLlDizvIFvF3toPxktbLqnyrDLi4PGPtS5GKg9L5BYVb4OV05i
5aKwEUDncvondnY2ECBbJ40jNJVAYKY5XtUW0Dr3g92MsjBTqHJdSgj6p/2S3Gqg
I0H+yeWt4JHKzqUAvvJlVOZ+iTg1KlToTDnJnSkPYmhEd002ziI3wS2vzIDJyT/e
1sETaOXQs/knDL279nLfaoUfy9w6BAr+sWOhI5DV/H1hCVhBduUXCSrwButMnBsp
S7+b1hm628YcIb75oloC5lNCKL9SZ/z10OuenDcK5tzogTeWp4caho7iKyNDkO+d
2ljr1iNvaVBCm+yM8HdQHwe8qNMWj0U+pHWun21+1tl3qLY8Vk5TVvY37Tzn/doy
vxjqSwii4zE7gm70qv7sZ8bBUejdR9RvvfF1eJrv3aTW4mHCEdgfYsJ0IpuTEW3Y
4iizVlaV4B2IgHeJ9gVWr7oN4tJhzybv6K3CXXn6zetqVpQ8NkqimSo9sAAFHRfY
Um7Lo3l2fhtRjwjqfw9AqGiAQJhpmU531RDwA+rEeIop451HcVbXoQpB3QUSk2kL
o4Sgzp0LBpYOlwFRbk8i8jsDGMR2FeL682Nl2GCebssEs8+gimaucSx41LxB4iLC
0/IsdtOkt5RdQI2QtAbj0N1fzPIlb8IF/xphkw7Br3WzL1oEdxlBcmLsKClL+LW9
K/8vp8A+E/biP2Bs/1biel3lj7OTS+5KcqFXSmrENJqmHQ550ZhxYBLlMB0jCJO9
v5U78dnF5Es95/sAQPZ/aDf/LKX8Xjzlf7n7jsahruAss3WeUNm0zeF2WTv+CRne
A94UoufR/QBrgk1UOhnH/dQpeEv3V2C2pia4sg4PVP/wYf4lOGhb6GfVCnUOdDzJ
Gtp4zDsj2HVrRY/wlC4mbA0EH8tlwD49O8HoJ5i/+vo+dx/b+K64R/htfFr2/9iT
27gFq8QZkK3iXms3QHuoaJMzUFBQiSPUJS3HmH4A2FxEx6o+uAaTkakLKYpsVtL0
2sfZ1nrsALPOpZvMoTY2gbaA3nF86bUYeu5yF3cLxdlljCx9e5wmt7dSK35m1PCK
iQzR28XMaUsP51fBzKR36s0H1/ixyytRMHlqATyLtQjOhs/vZQRhoMBHeJsd2Z27
RuNGpuVQT5KD6OtT2FuylCJMYhJ7Vwic6Q+iC3O6thVazh0oLqUkudccwc8Mm6Vo
FoFz7IyCdpZ2EqJ/k6LKF5Cm7UnLxqTAtkz4ix9V8t12FqlP7vlFvpexVQVowS0c
0J7rPr6gtf8XWO4pAkBayXEgReSLOKIkKh4ZzAIr3vU1q8MqZWeiFdT13TSDCmV1
E42+IbPwtXwWMj9fXtQh+sqayQA/pc+ma2r43d4FdDxD/N+AtZl5etW1CawnJUCo
dd+p2ioWFfY084za2Pfn7HiGuIBwK5NXHaCt4IYkYnBYCCllbzQplMUPlVXGBsfx
7Rt2OCTq06Rpb6Kq3Y0NW9Q05U+s5Sw6X03b89bYDC3bSyVgO0Cqe1oSVR0+FYJh
9clsIUOKFZjBIG/FDFoO3vIK+0tjNmjWPJnRAEqi3RN4DtA/sU+xSv/2m1VAqJnV
LFuPS1tPnsT4S9121MksFfUDKNrwTJzDj3q27RtvGvc2lKExhV27QmeDyt4aGS7I
6pUsGuDOFhu1cpKaE7GIxr3UNTeQiJK62dA5yhn+8FAEA/X1jgkrY6jeWkqCkkX/
JTnWKGmX8yMhqKU5g6XZ3JhRkXSd47CmMNiQWs63PeEkA9KMxcLDBIJ8/07+CjX2
+Z6Tk1MapPNt6GvLR28gNSMX19nPiKU6kDLsBSfV99m2Uuq8LZJ1f6RorP0mIcTt
W8EnqyI2eug3eZHNY+6g656nShXcdNFHM6oznDSpvQretO0O0iVAcwGpN9XOBsW6
sF/Hl3zXl35MeUwBvdIGgF+pkKeWylnvIolGQGsUs3OcESM4o2zwqEsX0wRX9635
YQCdBCzpSIzCuwPchnwCY5VZG0s/c9BHjfnVXynuHmqP/NsEJ0+XOULdWUNwe3Y4
x8SuO7ULNsvom9dF8wjGQeDTiRugM64QEhaVqU1NQuKkWNxFpfNQUfcXCKseojRm
Biphju1WXXL1fhDcEV7AC3mZu4fPMxDt6F72rtDFTsIWYotr9OutLuGj+/W/nzcf
HROmYsBbIOtNlUGl6WfuXlAZ3SD9xecgCXje+9bAS28dumAA9Ec9HkRV5rC/Om1Q
tpli4HwSrIHBU+nGz7gvEvtebQFrCpta18F+pVmsUlgF9TJ44a3CJ/ffSI8ftMha
NTFXEiOcZlrT54PZ93tbuxg+jTpWuWn53U2KKauXzaxqTlhQbK+i+9lxvyek41es
u8RyKac3LSN03OjULivuhR8ONJgcSlIRCRE/+TlmVoeCJ7c+A6CkDWB5IX1I9w1f
GKeiHy0VW4YjNcI9qCWL7sWAtLh4a/IW4IzBiW5f4Gz0CY0IZA/De+AIbYHlw5Yc
rKYgTKfeZjjrb6RrWLhlJlpN/zPUtwaUjtFnM686AHXqV3blorAp1jAmkCPasmdT
S4NWsWIaqd3qP6GREodU7mnceDNmxVVOYraFOGJ/UCi/7aWdS+30SudSyJCWdeV7
4BrtnOJPPat2tN4055/c4ultZ+JJgmFUDkOZ58teIm5t37WrCX6DoSrxX713AzcC
MIt7EBT2Rub5CEvLtXOremIRSrVi3VUGtirSnBt2SYJRS6YQahyjUoslyxEASX5b
aB7mYYSt0Fqk3ulS6SmFzVOG8cUlzJ5RFTkPjMm7qVLGWTYLtzqZa/cuA3orlCiG
P4D7b3lDVY577gg+RAEPnO4KyxaP8LhIn1LK+OQyQUS+Ue9NxLKxqEPrwY2Y/hTI
vGf/LalMQvvXoCllyuZcxNg6bxaT+jgN3pE4ctyMneqsKTiPmHyor6G+wMHuHizT
I0NIJw9PoFGt7ljgK3P3y4u5iQXg+yDyWqFukRZcOrJD9tr0kGs0PRSVY4HHDsdY
bYN8HsgAacgNT/65DVzECNgJdsIUbl9cYURm+aF4ZpOIknyFVfdcD24OLhWjGctB
t0n+1SSLSgiH9u1nJVlGPTHRYk0jX85i+65qGCwn8piykihUmJJLpwp23YzzqYr7
ohj8H8mluYVmZ3AnqvXi/ajdCvgRqWX6x4cf40vgs6x3Ia7JWjfE2UD6JbFtesHx
aIX0TIBCUCpLsuXF+eiHfJ7PrcCALg4tK9/jO0rbF2wREzxFbFSnYcpczGmR2z9j
AJRM9fngFQ9Y+K0woLzXE30O6qvM6sJNNXyKJJFkwInf3Ih2PCGQ6tHnYbF34bDZ
HRJsqSy82KlW+5VdqWDhn3Bc5rrjhlUsyJ2OIwOU9Lip6gB4HOMLMyN17UHu9IZR
Vq8m5XOwQW1DKmAaGO6Jk22/HbzkvMtw1FM1TWumyYmp8wtdX1QmC9+VEYeuWksa
YZrkWS7ScCWmUP/MAXBme5BCD0D7mN/3hEr/dij2zsj3jXOdeLiCQolB2mxkztM+
ZXKGFEtqEixQDxslSNhe3+dAqw/FBxfmUA60hxYTez2n+Abp/XS/0JQVeR3zThVk
eDuu40X1wyzosgFSS1koEI1w4W2gUyvJ7AstXLNWptqfvgY3NG3X4vhG+eoM4PLS
ypl8TPedi6QUJmNsWXSMWfBBQcZdvaP/vxO6RztFqP/qb7ZPA6AMYOAVBY7GpqiK
gfLK+1IrtLmq91n6DxdinsJ58xHcZjZGmOcv5o4fKQAKVm6rb3DHXqXX2ky8ViCc
7WdVDH9EXqZ2+UQ8kZcU8VOSlqY3hMz0x98XFBSkWa/PLeFwYHLbNYQYXbiE20VQ
Is0/PJW3e5me42GsFHYkV5JEpxLCqilJGitcT/Mvq9pdBcSacqUcyTyXdovtkUZx
J2D91ilG6PkBKKtLE6U0ZeryRqDWxJRIrvPmC/X08vtBEN+hGKYaZrlYbrf2Fjwy
CywlL9IfBBWFY7S/CzszjzKZiJ4KqKV2wkXBv4HBX7B1DYSnGoKZaZvflmVv6mR8
9L33JdkP2BhZA/YJlKFCs9miXzRlV3F43Ubp37fuZg7gxZBzA0sCPxUE7w1IA7nt
wb89Zp9RMbfH2PhmxXl1EhOOKVXicuTGg11yaknvBerMzYOOuSxtT36YW6vmB3+Y
O4sypfoNb4I+asLytffpMLPPh1yJwehmmyBP8TqTfgdWAOFGE/FpreVjo6GtGoaH
tZAkpYqdSGMfiNChlntkKCH6+wtPrGPjqBLxWyvLltLZhQ3Vi4tqYtEiupwCPtcy
ydM9VsWWbhfFq+vIwP49ehwt2usQllt8YXZ0dRdisYF7Cx9y/8Qu83jxXEtKOL2P
08p+cOcikX2nI/9zKM5SzfAXKpIYpCkPlID5N4f7Wu2dJ4ZiJnR0Ka8m4lG2zGjg
xJ98+5ffgXTbXO8mkx5rRE7vl2CvmrgQ5PdvmAvqCBUmD5BJQTYOfK1lCE2fVRBj
S8DT9NNau5S88Why3F5kPeyb80T94nNZD2aG35kCbOL8kvoC4JY8AGR0u9R3L6IT
mu060PlMwfbI9uUy918x8PmPL59/Idz/Ufie9OjSOmKV9I5D4vPLozXwhG8OFJSE
DMB93rB4yxkpyMpnt59ZnydSuz92Uh0LGLBjQtQk/CuuO6EPPl+rqQtAmbAy2TUT
1SqvN4YDm0ZmJlA94bi71DUSg+O6IgzANrQlbXeDh6ORaGtpjhvzhs0duVEBOzR+
Z+C+k1wGAzzSVIcQjRINR+XNethyxVaEEdBKicSToyNimu1/T+Fylg/qChmpLYxK
FKggyMKttT9Waf/F0c+q/DoA3NWBtGzyB6NmJnRMvwHzpOIUqbZIzhf4NZaVmf6L
3KYmjT0stczmLUy/GgbWG6F1MLyx9fOxNfCQmbzS7RcK6e4qlmFa5BuX4Hj+nnst
GwRQE9mLHNIaKo+2HUMVwlpC8MSVXnr+OqmR8sc84SXFDhXkSpXVyfxa1FVmoRog
RFTTWmpyZwEjD0QiRSXSbz24IeW4lWpG5GeVHCihu9L4oTvYYlCP8vOOOp+4yAIE
tNI20FEPmya87oWYlCS6P2O3+GZzkHh7OV1DIFAPVvV+vFFYRAFlvRRa9/pterrB
Do/7kkilcqVZYtfZdl+hJOtiqwaqkGIdLgst+tetazHUCunbEbOoiPXs+aGZGmnx
avSHMdVcVvVzUO8ZOCgpzWr5XYqQqiQJ5v8S5ZN1nyQIdtMsqKgADyAl6sI2DAWI
JkmFf0g0amJzZcnnLRE1X+/aLPvgRhcjXndfenSFsm6Vk+RnZVcg4mB3DRrD9Tez
+zEWRcGFuoTwC94zoOTqSNRSJuiZJp4miwg7xEtX2vrtB+meHPdipy1Z+LoieIYp
ubRoiL1dsBwpT43rK0PlgBu1vBP27yW+U9ZfxLQ3qJYA3WIyNfmisYk7mSWJ7acb
wJ9kv71E1ndFthtPqf+MMsZKVnjFTEJQvwd6UiToU2kGnaMbXVH3wfPp9TkAYWtN
eOwN3bl8KTux+0lAfEDIaOKySLH+LUrNnEc5zU2L1rQkSkw4BOC/xpzGeFHwDHDb
cxbeB3dyMODGV+Nhueta4fDaWNGKpFjsNkEVRH9rytxY4jDYAfl9ODP8kNpUMiV8
30vk1q/tuy7Mjm5O8mOcG7ZRYp9Ygs+7Ct5x3qIfie/x2EXV4bjeoQLNpgAs4tF3
eYwEyycThkTYfGMeKTyI+Dg9jy5c92q3Hj7/xMO+1nL7ng295IPta9XyEXpp3XKf
qLtzX3NixpnOtKX5mdK01WTtOnFQonSmrAEVs423vnTqdW8UEXiP2JJ10XAXBIol
wRq9N84T5AgYzmVA/pC0MyDKohD0xN8m1Ghdncpv1/myLw3ELQ3BXjA+tRhrZgUk
9qjfqWedrJKwRC+h/dV78HQn97n5aL5/ewtaB9z2dxJ8aXidYiHTxmmLq+PlcISt
VuF5refnwMsBsthmOcP3MP/4f4CZF2SHTE9od4W5NCA+jQLdr8dni54w9oIIO0oG
K8jkqOZ1klksMcOxpjub4AHuqo1P+4hdbgJDYeu5FFLC4htnKb6Bn6P6jm/VzakR
FAKAB3aAcmGniP0mcEJlCOCyOiWYXuypfMkGy3eFn+oHGtZ1Rc6+cTU6TsE8yKHO
DSjC7wcOMJp1USS0TNUxB74MfZqj2WpY+utyaM6CaSDfAyr7O0ZH4rc2XrIWzHy/
1Gpd1xfgZYE2MnYd5hXOAxsjL6jtgzCQ0TVWyMEJfK7SCbtyPEz2/5mR3saTL76s
LNoYmgBiK2w/fIshPMLHtXij9tL+I/g6dcW/7X+3GPq6uLxR1G1TGGH0VW4KtFoy
DctZ/OUlUqzatn9KHKPiKPfIvz9YVpURuAFxuS5Mdij6csrWFMkvUOKtMTz/55kh
3xw4hNxvtrOEq3onR2afQkzM+7ZRV7raIrnmjMIlaj9D1MWlutLYWQWrO6AhK+ag
PUw2hKKgyCoMkFUlPXyKzP4sztM+9l/70WMUGxPnG66ob3I3groDm1BMEnqBRBjt
AHZ5+zxDM59TfvUkX8vkDyyYjp4cxiGUgbk8zVPWR4XTLOA+ao4U37zYkE/NL0/x
misM8lpisqSRZA+NmvjjUuejXlifv+txilVBC0voCB/f4s80G5KZokwyLDZ2W2YX
hYFgeLwh4gqyh4OFKrzZ+G9bDM60SiekXLqNHXhsK1rr26fRMi0SjuKU1to6lOC5
2q803mS1W6X6wdH3DqwNor67pBfArih7EoG/8Ksz5X9WznO9CLI2aJRnCX6gbEBo
rqEm9vW7Ys/f7zpnLTir759/d8tQPSY8iRWLsYrqtaJEJJRBBCEBbi8mklmDJwnx
kgBA2bYfgyOtbXjaIyiYmg==
`protect END_PROTECTED
