`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9JLFXygGMmUfI1N/PuzMKaxPJOUzXpsVodYanv7mu9oz5amNKFzAcNAbQpvTKmFg
oVTdsOD93kv4Tx+YSmPs+wmN9RzSuLxUROLvWznwoZS252PEDanXhpQ8Ro20Uhwq
aPtX1bgEcTfk/1AgqxxqxA8o87Skcmg7DDci9QwV9B+C1o/gbkLmu6z7DcOB/i3Z
ZjifursvNL5S74Z/AfJ8OFqLPRNQPGRDE6HU+B65bvnUhD26D5AQ3ZIAx/TcRdRc
+Dw+Ko6F6JAWYnTJk2JmvhpFbM5CBxsUX+m0CLYuqDHkX4m1Hp8EsKjiLKlg4JdD
1+yD86JcTS03H26nYxZjmsDprO3j1sAr37uf3gV8fulHY5bsg8BlVD2BIoPyLN8G
Q0YvPP2aoDqjlOl1kHuYvuspvR9NUeGtPgWiNaEp167xPS+YzF2AiyV3OcRzlcXi
OVv4nRavQ10KVAfosW7uddSU3ByKtpd4PzDgTbDb9gR8nH4Er0v7yY7+H92HInfq
k1j6kH94inGxjgRPfC7fL5YiMI4Xs5Ew/MPI6s9IdBI2YADlz7sUkCbP0bzOc70H
XBKciM4obm0+4QrycaAe5JJLWn/lYPaigiFiLAD514B3vUF8EKWAYY0xuYGvrwqF
ixL57j9o7/MaFabRJu9a3vc6Pbva9I4rYaw9+krxC42oo02hsL/5z4hLauHujlhT
CUEq5iEkvD+kV9Vzp4Q4pP8haysL3ywPSV/pJYuykTdq1U8v5D2NO2kdmJG0azxj
BITOtevgCaMtWA49uJd/gYTgkbWpd0yKdLPoQ7QJ3uzGxm4foVzd1RZclL9mccCh
ISqMmvlj7ZTpT8gl/hSxm/mL1QJutoqQBNp+tQNghxHxjIluq4a03Hncjm2bpFat
wh2AQRq8Vh8cfzpPbtnmIeaZFYUCd9Ai6OiMG9DD1zTW3AygcSwB7VPJKKFos5QY
zL2Sm7x6KTM4+NRezzWgSe1AhtU+vnlukWbib/kh24K/jsRrO/7oyzLP6jw6LVmg
5W5wgkJmaZZNso1DVsK9CrGgYscTU2nSTslzOrBJX4BF39fG/OovMeT9tTuNi6cc
1uXBQz3skVobFFwn08fhNd72aMVOwvqYymGkrsz03hpVaU7rfPK55zR2rWvcKO7B
qfU3lgmCSGijA0eWIwhMOzWsXKLY67tWhUwA66jVmbr0ajRRQWouPmQe0IUP0Z5n
yE+zO63pV5aAgQq4hhQRwSN7X7u/XK2kPVVNb4JHhBugDw3+ZGEhQ69IQ3KBVBbS
qUY+mTOB0BT62wlC3B27q5lc8n4bMj3DAvH7WHm2pGdHiFxQyzcynkUOwAqVxYb3
aKfeJpCOt1RAputy3qf2IjerP3lYladFTSNN8bl530V2hWYHa9yMQvIBmmiiNcSD
PZHR35aBG5T2MCSiA37fL8JO/+OmT748vSGUaddWzUx9XY+y+vOZYfj2SkjigAT3
wS2rh50YcfpMGYX9Rt+Rl3ltYKEe0O0JHyLEUNSCCqqIqBWoVRzNXL3+mz3wHb8t
lk5S6VaV3fIlFS6q1SqcZXw0z7s0Ucf/sVEdkTO85TD2l9yKldt6h04LMHlH5CwH
jwEQsKMpXkQVkhb5Hn62ZSsid8liI/touQLUjCTYKEb1XWTLkeYJlsNVByDYv0wI
tx+t2/Wetp/DSXMCgKeTG+tAz8THHsAtzA9eOJsNLFvAn9MbhNSmZdOjE4jvNjlS
JOWgzJBAlBeN7RBsa05yolUV7MQLu0poQijSBTjvS2s7bz3kB4lu3V/95SDnhagG
NIXNBeeW8Xp/JlabJo2LP3NOuND+gIXw42O6A94F9R59Q+/0/dB4Z2Z1QIu9E4h3
mXu3UDygkdqYD1RsMjpeIekeZwpIRWk+2DFemB3Rm2mWHBA0Frz1bZj7QXG4ZmIr
5sROTnHhzFa6kEt3VxuimaDVvuJinHh3SsJTbHTXKQPq44lX0VLdIa3YhBfPP90J
WQO7MeTiyD7qxEAi7YpOQXTD3DvW+2xARkzr8DU0GZIm2onuFvR6n53mD4hXhkTG
+969gh3H/XXVKnoMal2US4/sbsAv5JW9LldNQoiGQhfXmPkgsSK/uVh5V97p7fCa
4R56moq+5tpas4xbbT2ULtZE/a6pgjboVKenQjenNF0KOLNtWKV9kiq2OdwQx/sd
tgOcrpxAvwgkpfd9V/wJy/zysS2yrPUKESzfH69Aqjb2iKsuM/Ysv+OQfhwffetR
jqKEXtdIC+7eVcz3Odvg3M3hVXyjdLSfwF71ekWIWv96PmgjP8vhzXZDAPRol6Ip
NE7uOCsG0zxpY1kjphcKINejBh8VptEH2csQFbmfqAe94yMVrGShhUX0JlwJT2ro
rY8+NQmFn3cHoNvtooQKdFlHgFav30lGFt/JUXFrcQPG9E/aGvMdyVMYdXEWZSWF
7mts3/4TuEJQyWasnX0RETlSF5yn5BvJ/4+RyPGQE7Tu7pF0lJ7c5ATMEfBYIHVK
qxVN7RifS8oMuLehuuJNwSQy/o5cuu33UFXbeuE3mH0c85OYKhiedRiZ5FYlN9gx
Dxi4o2H5mYgQeBQRa29lM6izRsD5Lk7f/tuTAroH/WKHoFuNZ14tPcBVzvXyUXhH
ZT9Ec5XFTnyrgl0icRKKa/El+6ehIRyPCiCQc1j769yqCCV2PF2ztdlEjuacRgaK
Q1vDQ6YBlaexRCGBlAecS+yheBpzPmF0BcrmeJlTqOZnB6P2wNOWKWyEgY2pwoz+
kNvnaUEJxD12YRSh/0DRV1QCodydRA7BLMAFQvd9hK4U3z9bcGB0DVGNN+K8iOMg
y2+X8R/oeHlv1QobMX9yihRZPlYDeOtw1D78126/o1pDyRAU+BPcyxsh2HErgs6U
hcz2XtJ7JTSRXwiHXG2b9FkXWf4D7M4khfT016460QAbWjzHsEpQLMf7tl/7mzeM
m297Z84xnyQtsIZWg7ppclK5Kv8eom+j2OX+OF4NkrIQzxDahUtMw4WTZAoPgoB9
xBO7bgypMu1+533GUCswiFLi+I7WYLuWj5Gm8OJcs4iMtgKfuq7cLGzJxhoMZx9O
2yxN13JCx13Jay4ob1vF3nyw1yAX4/ADJK+1/DKxHhMyi6JCqTO0CshWchz7xavS
PLQ1F48DfCgnXZEHVaCI2wj9944yYfEpbFxPG6+vLGZVFrAUNidKYDSga0l/fBzA
0nHHeTuccMKTPpvLXVYYaDpV8c7k1JMvwSb3XCiE7esWrRc8J24ywVVL6ySkysd5
dyqetZas2qEPLxT4ricOQ2Hlkwf7Ee6Z3hMYkEVCs3K+qImncFlDTU9AVjKcDIbQ
7O1O/ATEXblcdnyFcn+WP1ov9Md5zYj2nKGmqDHYWQnpA4+FhX6VgDktUWYou8aN
JQnnav8d/p+qu7zjiyD3M0fgL0kNfLHEONh+XDckm0x/nPZDCT+JhGbB0d/uv0JU
0QVY+AEsf1s2BeJ4m59WzSmBJD/lq9eFZAkfCohRaiVadveDIfiAt95LCZSeTGKC
pprS2HpVtc2lCe4HxiC8Inzk/09DevSID93doyKkn5QySk2ENDT5SFzponxX4pxL
1UbG5+mpoO4tKbM7wFhwo2EFVmAhntgg/7qFd/yxyCKEAk/XcdlGbFXawwOty8xZ
sPTAbHY+IjQmsyjUXoRuOxTpTqfRyDkgtOFAmHhch7v+FuCXRSWz3gZn/wMPL/Hw
U5NkKtYkJHy/rMa62w78zWjtZhh6pDIJvnbEoiItFv1SoR2+gUTHOXvCUpd1ZVu0
T8YlYngKLmInPl9WEXD2bCgXHAFD4cb483DkyWNQKry+FsRpmDl5hBVFvsQq6LWD
plrOnYc3YYIuNZyzpn3aq4Xxzaqt1J2S+E6an4G8mRHf+33DHMUvmbGb8B8j0XdO
3anye06PtYmVNpSkTMhSRbjUjKQgyILBt4aURH4WXRELdY2j2P95clgAGACWBKDZ
loan4qCs0y8RGuLZOo8Y4/tfhgXTcGPaJYxD5rgSkbibZir/AcUoxpNmLLB/wpCF
Q1T6mUwBiyoz3znxixSfe4jD2eo3ionsjv12RWa9m//rrXzevqBMVPetf18JFW24
586q9Nfjeqcpe9gyrEN6y+FeVywxxi+l2WTSRJZh996G1m2LFhYMNpwAs9WIDcnW
0r4lQDipT/rbJvIgcViIDkGidnctuSdQk3fhmQrN5I9CVYGM6wPog0Lj3PV6iXa1
pozryhUQSfJTcZEwyFb7ph/2Zu3NbqHLgM82GwVsFEsLEGm9NZYOtUVYupkKLas4
3J3oJ6QwklKCsX38CoQxqDpGB25ZOxN3WUEb6XpSKxrQX27yHa7ku/7gbDFchn11
jxT46Ev06J0kcykw6P+6YYSLf2aUt6EYM/No5q8sRgQsYsW1zIFzy38gk+Wt+Xvd
/qIgdEkf/XrsamkS0gle0YtVT7yhXpgFcu40V5gcDExyRi6tu/xITFN58i5Jo0VO
RPZPDQfwPDpmcCPUxpNcMfz2KghDODJb5oXlHm28wNUr0qm4ZGbiwKrSDqgFC1oj
/vDh41WKNxutwZh5nuUCxtmdsxrzLU21Mv5RMHvlltj4Ux1crdrDDu1OzufvQSvD
FWozPr0SIxXOkrne8m2lyFXL0J2XT/njw54KNNs0qKgDsHlCMo10OVGtglnWwlha
GLD/r4nOz+AlrEjNS4CX6O82JlXrTWvPP24wtzYiNz2ZeX6aP0wcwAhIfHq8NnHp
wr0YD2/jSlHOkt2X76L9Imw/VBBtZX/LeA73WTFWGS3O0tCE+n/oyx3SJNiZZra/
AbrWtyEbYTErGsrtxjKLgI7lSQT+EVSsRT8RYRracgWbiVdd8Eg/GO6xNgIDVS3X
YH5dQQRXjVW8F54m1oFsIVRU09b//GWHQB7j6SFInMpzL7hBWcUzti9VDIfY9A3N
Ns61vaocc5XaC2i/btQ5tyUczmz+ReYRhTa+z+CAF33ExGrgQl/QHD6fYv/PLOFJ
+EPscUTBboVwtPRu8RxaOa32Ug2USTAmhkiPkZrFSnqz4jpxSVunigUiDNTSPocl
IzZYP4FEUe/1B0Lbt3hRw71T9oVmZwYAStpulu8rMmqfXc3F7dOcUYGRHZXyOFkP
y0YkZqkWHQpZkbEN2mdOq8c4LaIPLJvDUXsmn2yfeIUlP5AoLQ1VyZvIUtE4x7GZ
7S8ODjpKhFjMoj1kphUzfHSEVqVO9sufrukezWdi6MlElLtvCVJGJ+tMqcwO9Lgz
T27CcnTPk4Dwm3K/HGx6d0AvVcQzp/oaY1Pf3UHV3FsCNZ9oRnwBgKLOnlbELS+M
nvSfNIwzgCwA+Z9MOFRedxMLnO3g1QyoeV/aPvBnE2eW96POJ0MURKWgRj8fzuM+
rIlabZi+1XkoTGC+Os5LZUDBchks9Npz+IW46ni44BSNQI9aOZxHv8KqWF+GFGLP
hcuMREPjUOIh5SofB7UIVzH9WzVgu1nr/I1U4thSusYVQ1MJn2PK/CSZ6IBnUO+Q
Z4zTxWI93sIdiLVHOUGmmWbn9XMU0Z7Qemeiyb4pSVM5xipGjXLr2qFe66bpveTf
wDBbZ7noG7D2/80IL5tC4z9uJ7H0MRs92MSnZc0ND3g0SIde+IesyMhA3z5bglLb
FeVLfpVl2QjVk+9LAkW3AQDW+mM0A13BOFOcn4cOB3Bz+7Kei7FX9IgUHegyb2K7
056Z2FdNp9gPgtQkF7/Bl+JkKojiYrJ2qY7PAFSyLSMCj2CvnpEQjt5OHvWNT9JN
29Zb11NJKirIKIJdM7A3ny5EToklavR0YZ7jch2Gz7gQ0AhT7zbv7/kTlHvGpmSG
z5cUKG4BESSvKR7RVlBwu0eiYJhF8c6YFV60t1Cl/JBMUWCxJyCsxCaOH7NfJi3u
MZ+yeoyBteEXUgQWdfR+o91iRsRvC4zH1wOTQiSrsQGU2JiLOWYmrNg9845olzxg
ou9jXiOLpCBspykepF/ssPKwbE+KpMYVPFFDRVBpc45di2yI1Elk8POG8+2pGyy+
CRK7Z9D3Kgtd+RrIQQI6zXrzjKO+DG/avGXF+P4WHvqferTBdpEKO5eOvdV6SHNe
VGohGg20yGCUDvmV2sg3W2QnzWXU0S++N+NxgZbQvhAJGlBAZLb5u3Y4jQxTp+pi
qakJedP3A1m+er/BenZPZbe5IbjNtjfBTtMSpwXVPa1U2S65/gLXJzn5ZWuIV1kf
QSBhWNyXL6rGaoqtxiZISThYHJLbzfCm7Oh0DMAFrQvsEa1CagIgXz3G4Nug0Sjy
q+d8CsJ9fVh5SXoJqDcxSkfv5czoHOlCdb9J/8lY/OBy4KcOj7X/oKqenRQ1XVrI
kS7HdlrliliJARvDLWppOO+FxYcSH3Bh5V+CO2vBev6Vrv4ff0OX4xxQV7e4zMit
M5jzrlj4hWzhngyutEqESE/8hJLs9oxz7ywSMyMUasu9IJd/siFvp5/ICrCCw86i
M4T64RzuPIZaEnKoJKowuI3UgxHurYrOd7WmBSivfWDZM9+t1UhkghPZ3QgefMKI
U+RzPqXWrzcML4+kp5w4ztM6NEG3MhnXgAJl+u4+S99VXLNSUxWF6QnADBisBRqQ
H6Eu16dH+FagXZdG3hY2GnCe3htm2WLzak3NdVGJFlU8ULOR1e8MHFn+eHv49chn
XWrG+UySSeyPClk4q6N3iQP4b6PTZDhsGqnnb23ioDWC4R+S5dXXQGFZYpGWbvVY
CEWR+vNUShZEdFWNOQ25fm4U2RL1eJHzu/6YBKnhWHTNVq1NSpD0s4K/GnMenody
0rXC1y1cfDQut3z7qVpmvvIL4ko8kDt1Q730SQBWekbIJU5JygGPjj6xFM8PgyPq
PRgAmHj3lGGUEN9fMAE8xWvotQbxRwxQQNEzvRCVZfj+eMfQjqlXEf2XY286rWss
H3+327yafPGrF8P2OkpK62jq8HGNXOoDWSgUH4vJ1Pvgo4jXoqHgo79XsnlD8+rJ
ZLxV7s0CFPU7nUkO2mcwJpki6N4aTixApQJXt/VI9t7yvvJEL6UKTyUCyYHY9p/H
D/rsgSNf1xSG391agDeQMNqPin5vwSY82dPZuw2PSXaM+HnC0Kty6FN3cBCc9Xbf
SkxlJSKhVs77VoSxJPA5WRykPkdtzfk/oRo5E5DTEsiKZyV4qijrNlwAe1fCTRYK
PtGuOo/6zk/louVl/hbR7oWvssD8kko3LrQK+LP8Ahs8NJGDuJendG3tAG30oa2W
bN5KH0zIsEvPCY/zz6TmUzE2ujucCATXmTKxmIvke/wcoIIUmfix9TwiYI66RKYz
/Aj4QSv9WVgiLrJi4sfjnpVIbUZ0skdoedqpD7/ljAUh6il9dGkeetC0oehokkFT
AGcEU6dXfBwYWJZW2vdrDuXOHktDUpi/H45fscKmGJvWU3PvSnvnMssAX0tAlpbR
446sn32mYO9DyIdqxwTfu8dlbJ9txD9tQPh1oQbLuOjLboJFeTv5k/m1c2x9q4Bc
a9NZaW8Hb+0jeWAQOJWXXoRqcl+iOeDtCa+9QSG+tN2K3EdjQJ8Vdyhnwtu99/GK
/TODI9mNRADzk/YWiRwAZ4ZmvbXtK6U59aHayzaV5ZuQHKH/B175zKLRTZ7U+IAZ
OCOgbinKdrCwiigrqCFZX7R0z9flZlNSAXuEdHieZGbfVdWsyXrNWKz2sVMI3/EI
V1nexyRnkyx07/Ej7hwYqcjJQrU5s5CVbR3pA5pL/xHTvS26mF6ohFDVqyFljhqb
rxl4N9sTWN8nxiTB7809HjU6a+0jzAuBLRnAoeJ1Z3Lq/9spzM5vALG6D1cklkCj
BgeHXOG0/PjZBC1p/TDIw1nLqg0Gcruur+AX4XOfS9E0uW6n67ElPVA7EDBZAxPx
1XeZOJrFSCsUocXNLoMbeTWrpA327Sm1mhtzwW0zTY6i/T/xzl4R86DR2BnlXm6D
OIQG3tf3MzAMvUHfnDhIRlq9o/2lmDlx4GZd/oy98KIe7RKg4ydckFyM5s6WfQZA
t/XCbj0tXdKn/norCdfX1dyZFKW+2lnmekLk9spKUIV+qhNTDcwnokH5u+HXqGfJ
RcEmhMd5a1ZO8ZW2Ev9mdt3K2Gv2o19CHERX1PiiDP9Hiu6qxhqljr+7cQf8myJ7
fBa7Cgg3Uh5ZbghyL5Lfpq6HEUnREOtTuRa6UrzmmXbhFQ2zlL468YMtXUxfdNoE
gs5W8Ild0X9t4UyE1Y8oblh1bcS+HdfOPpt67sU/oQXvLq0zUDXivD4ItDn1xRXq
2qdEKPooV0ovNaVDL+tQqSoJXFv8nv9ftXNBJXzeJphyfQ2mugJTgyucSNTWYPme
sU9VlBdpOsEcHcjXTyPHVZBqBzpkVjhknQV4IClfgAo3QvSXzMMZX/f/iqsCyNJp
seGW6B/18/71sLr9oeHHE6FjRqcHvZDe+sWVy2TBJbwrzmW4/vIJAoQFyvLc9cMn
8fZ+fzhKkKucxTOxFzaeWto8sBVATgt4valiRhhN0hdTBNXH0n08pjguinAoNzu1
FK5qpFfsx1IPG3BkqiuTWoC0LYEPQwxDmef1MzxvfVbFKiwkaD6STK+cjZLm7C74
qiZY+V9R2VtaRvrbi6ag+7tEgsnyYPDoubiyfF6pJv0oOXP7smb13DtH2Ulzdvt3
Sa2kaY2tl7wxqj8rw1V3NjERyaLn3KPEPc3KoLpfailrspdH+yz64FPFX8RxOLN3
mHz7goZ72Oms/4HCGv/sHJXGnXgms2fNqNo1xWUps3OrY2RyKUz4oEMhmWF+SSYS
VCZeZ+jAqF+MWTFdPOPxjGMN/4y1ML3BLl23E2Ctxn8zQvN1tCN9py+tfDPqqx1r
/6upCc0B3XZXY2uo8/9ePvivTH7jgw4nAnGKh2JKbj+QVAXo623vavXAaclWATe9
ZW05A/wKOyp65hLJG5nNzOG+5d32MYy371AmvNRwbsSHQrEN8zqxMfa6Von+t3DU
vn1DZPH8F7v65VxJFhq8wtpv8E0trDsWvdlxx1erc1FjKGo2TRZnFvF/5PgkN9T8
5nzgKwkRyiEkhxZLAjpL7KLeyct9wAnZuuPosw94eZQ7unNCZAuo7ccMfMCC/CS1
F2a2hSD5e5UQWi5viFCQeGTvkR1tUbjH3cr/M1uN9lkaRD0spIXrsAP9quR94C+J
5DQydkF+4qdYWC5HnNC6+6Ug0MZ5RhfoZzILISsEJGb9dRQIUOykG6tFJN2DNNll
du2FOdXeuX6AB0gCvBhs/0BBqxUhuuFDBhBK0G1xOD5gp0gdTnGhJ9Dn50rp8Ffo
Z9yn9CFm8z55lK9bvBX8RjFrmcqsptzLCsWRfh99qV+Hh0ATwXmRX5eYycDDode+
ewEYAlu67z80mUuqsJazBCwFAfmjfQLbzSyNpPvwHyVgOqHrMA0R7qJoZ1UEMxsy
rd07Iv6ut+lQt7P8Aeh7ICLRu/dMmEd3MWVlLzIxhlRjGyHmxZfUbWPtNIsEBrjT
NiwYy6IZMCT87BPVsgxCyC/JD8lvQWN+nBGomgC+ln8B6YWYOlAZkk/V3YSoE0ME
FgJpQumOYN93hFEBiPNOGqc1tDprsmtSD/S5Zdti3ctIX2GY3qr9ppnnCA2P8A1i
6FOPF/IB/H+PiuRSiNCiw1dF9VGiZyX4NWEQRYflxRM2QVnMX5sfEbNmKnH6n/dU
Q+unCEWyH6xHRp9bZzA/V9GzCU+GJuevKI4LNmgCrZmkv1flTGkimRVioU6mawsG
llsfqiU59b3bTcXappPpOu62Oa0WTPvapHzGFpe9cQ/+Sjb7JAjD+XOzkY4ICDm6
rCkJXBH3ma0/QmVInbohcVeqsoaMwCs+YAOPC16BvjVj554TdlQEoCfU6ROomCla
CynqeBNTwAshn7qf/zq7oqrFSNhfN5ujwVLcISJY+X3M8h1j8prb0OUKN3S77nye
MA/vVdT1E1plVKmOcTQ9HPVulKkQjU+M9JpVZB5FZ0Z/0ijus2yQdJqP1EBYhq6y
ZAIH+xFMv+kBpOojj0Myk25FSh04D0eOQhcd9HcOfqWolJ8HFtgIKzmGFPqJTKqK
umdIxDF68yj2q8h9cYnrGGR2zqsdrmz+Ik1DeZms7ZxV3xFoNNt52rpslQcvBdQk
yyL0Yg027bewS7hTQIvEBL+gzjPkLPXE1xMcn34t/i9Ax48+hvgV2/5nVYmjlyfC
cddZZRlcRtOOSnQxQkdrQeLseSF2qXarOGgV33uY6D5+SrFvGT9T9r/Teo4/Uohp
ZqfDKtdxwteuyZq3Uibnav3wqA04uett7OZHux/alLGgQxVSe8Ga+mpaReY9nJeH
+Zv44kf6x7XQeqy7bjzBNPrv1ae+o+bbqB9mWk4DpOzsDpta+cdqwl+PXeWEKUAr
KIC80nYvPxrYj3XXrzBWO5Jz8SQgtCK6GBF6MUR2qQrm0+QSq96+ARA+EFhSD0Qy
KWRwOeUtWv+2e2/HnysfWnBT31SZynDuCLaFwmqgaMqp+eMo7R7BEqYtBVUUF7M0
dZERTBVm/7/R69JK7XQFrS6ihK5YQ5A10d9Qs6Z2g7Gv0RED5Cs6DhXyB1WbJTLL
+tRtaBLoFFqZWwPLGUtEfq3icWX6uK2sR61dfZQuew87pGs9oTK2drrjAeSd1ewN
jT3O+8ONwbpwHoPZdA6eUkHru3yBW7a5ixeC2zVUC0tKYnGZ4Z5vmE2JM9Pyc2m+
PRlf/LYLLqgCWYq3a8Y7VwtPam6nf7oepnlR/Q7jt43z1sSOeTe/uX2awYmNY1vy
dpzmRK/9smzmTw3X21Q98Hc/4+LKASg1bWg7DhHtbey7qHG2SLWyrFIJ29pJtVNl
aScnGqUUsQI7oc/b1UGvBanhMGbPrADy7pnFXdT5FIsacbVejxJRjvSPE+T3bi8X
Ersf7+inQqeiJYuCbMIqAS3ewnyWWoMqXl+IlLobLF5djZZjPjO9dU1Kp9W/faA4
TzhJ+KSib4PSs66SV+6ef2mpGSHAXucPmLpTWQ7I6PU6sSfUC+27PTv4GQGX3WBI
4C33qXgUNbyJc4j1lS7SuLuK6GiDgONVMK1npEHiyHdRvStj+d7EsvRC/82A36e+
YwrPVSwsmcWXjrjOLiASl2OZFSVYqtLLLcRz1I7Rr7z/4yrTdYoVCQtke4nXIfdL
Tuj1qW/t/LW6laXB07IOQz6CWWWrciMKZdEMbwR/WXYG5AtGzRSR6U5JTcxpM8I+
+MKJYwX0dAOaIVrNrZOX0qnmgRCpMbtIWZcScArfOdKaAphd3arvj6tGVhjDFaQn
DOLZFGNkqL4a7/AxRUuMcHHOmkR0lZLCKXjAz4EMpLu3dW/TEVrshjCCEGuY/CJX
1vWWSKoioODPIDW8pruNZS9Iurv5zx1GF/1R68XjcfbnzEAH7bhwFzKHiKCqhzfa
X0nE/HzUa6jxnJjHpZBeChjyxVeDPsjR0tr6c2oIMs0NUIdYgrZRgViIlkDL26m9
Tzoy2MjgsWTQekjHVvM6mqareTcbniHStqtgKOjy7Cn6sRY3pZRqhi4M1bJtJDim
lraQQsL+Ymk4C8y4xExDeInrH14ssSJTHavqPK5ury3DmVJPIzJ5Hyk6zkcmRsYt
yNZ3EjSqeCeIDXdDAZsN9l7rWyVQjXgFueAZCTbthk65dK4YZYXAbDEgq0JY7zTR
OJnYudiYXgFIuv9NmVHR0AoNJwzbSoGqUFQvjc8czpf0yPLXb4ZFhWkz0zJK/7mH
jmgpzx2fG2HMtWCZhUYymQ6MkVNQxSL8XozF55oHMFXZvvPW9XuGwNDAkzerKLyT
44lfd8zjFhGNVpfpvfMJfjziIOyckEBchMdvM5hxYRatrzaTVSW1JZ2UQi44HO8J
hO2mAfSnkft4CXKMOlV2o+1+ncBFzyPnqPH+7xYc+z4ZcQBgePtfWR92XIhhd/KR
qviTvferJo3/qmIQEB5/H0tCL4cHrjvMUAA+wDSDaCWlDo+ocl1He/1lgkt59xyk
TVCXWME2Cf2rz5FEY1wbKuOtvMyaQ2eaa2mvENdHxGR8l3nTNP+UrzBxg1LTYkOu
a9c8oVgyfromYGXvJSFOjj5FTD2/JVriPd0x2tV6eB+VuTn+o/C5pw0bzgfU6ecx
RkKz48tnad3fHZlHh9W+DQvGgsMPiqbK/hY5If/xB5WCcr1GOnJ61D5M+bGg1oQW
DCFvt5bB1irhQEk4haDhY4WCFz4iCs4clcKWZ5UmyTJ8Ri3qh8vP/9K1BQbwGDQV
/HooWlV0PYKU7IisApMjdzKkxZXF9qEu0kycOC3qsd18vgkOxRvaCgYdE0jG5tRD
40kUxq0uEAGKBUs28FXtQ1tR9CqxrCQGxRyctXXk1oSrOhgcMnEdPteZS21iix32
1YfoC58hZvQRIwd3OZBnmw==
`protect END_PROTECTED
