`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DDKNRDzOOlBTYGTBCnFm9JWjI7XoLWUOlYu3ndQEb1azFjknMAZmg+uaaSxbcWCH
I3/ngSc/wkDRceeAwEmrPFU+oBl5B5lPj0EPDBrZekNnkubCycPpUNr1DPE59ekr
z7c8a9Av+4G2/80j9IfeTjZlWcg4cSlvMDPHx/7SVmORdyDuLOm4c4k7wAATodcH
Q8KgXZ7d0oODDFfjNrm+Xc2Lfyqll5e8j+yTaj5UdIVP7yFYeZL01DO65W0c7Fe9
SEV6hMOQSdAZ+n+Q4NulqQbBgRr+qbBMwKnYYY/UcHMbmzwGvRaDoV0Cht/aHbUY
2hAIB42/i7wjyOyrmjo9n8o587Pn3TjYggHeTzrgO2tpGeRx7pBga2pkTsKu6GYu
JX2u27JCE/w6Zn/LIDNdgbSzwWboUYSQql52jLdTBn0miN3UYrmoNint5RKDd0Qc
WHn8zTFDZieJHyIqtg5AsK7F+VZ53WghblXNUdWlg9dfSriyYKU8V6IdQF6sU+TI
4XnuhtTmKW7HdWqrUozOxMKR3RpkCuRU+tVJ6jX0L0fI3Ygrx74vIfsquZiaeSIi
Txx4B5H0KjOsoB6WfzUCa0ZSEStdMV/8V/fCyof1jJJoHf7+2N6rN7ReC4APBuTx
8fKoKvlwmn5DaZ+3ygNhtWx1ZznSte07DYsV1Ynk58bYkcfH30WITpoPDnTeWgZJ
yx6M7xE+RWSyUmEqSdTgT2PnVlxlgB2GE1wEmqABRfSGubokMtwQ9Zx0vfXyOwoE
l4A2apXzunAEwvwM9rrxLGflsDOtyJ5JC3Byq7KwrCfda4GVos3Kg0Onn6Fchh6X
6bQGh2yFegr0uXcY20tqpjVUK+UVClFXZN9xXG6ZTlwEIU8RSXFFn53mIA6zQXfj
LwfiArUEZ+dWCj3GkKYBs25aHODVRQT7FBBBFRLZAs7lH5wqVtnhLWyYA8W8C+Qv
JMZlfMZkFXHwIwnlh1zMxkeqpaxtHYEZ/bu3ALQVHTxny6wzERogc989E1/twKFr
6LT8fhKhqhNhpVTi/gpWYAmcKLmIGLKYhd26swDoG6bqUcLZqH8taL/2LwwQSHRu
nTyg8U+sRS+hzQFJrDAkhqOtwOjs+Dq7nuhVxjVR7zV8d+Tt13pPvLJxO6PPggI+
mUPmyw3V6y3mo6Xuh8YxAt+amP+te9k8vzDxD+Wt0qX+5THS5OdglQwR4yV3rtG6
/k+254RxKoRzhhNzjAIzDB/1/Fcev1FgOmVzRDBGd/L2wsB7DZlQ1JilIUzFdYOK
9wUbJog3iKqXTAaCL6LnchYINl/51XgrHHskDIBrfI+zfgotnnLcx2HwXm+iSQuK
/ex1PJjp6CVquXXGd0FYF0It79Ju0LSoVw1zgUnnZ1pPNQWAEs229PsvUViXEynG
J82Pgx9vEKRFtvR+73sZCWN1R44P904bwXpzzSFZCeL5kblaCMlIy5jn7j8woTLc
rFkD+xa8fcAYQGBos8Lc1jqkDVBaXGAdpZBJWvE3x+jEnuQMzVwBogt1x3aSlQf1
egOs3sZBn4l73QkypNRVBfbGnsFX9+O3OGD7CoPTYA035gFj4Dt8nF/iIVl97Qh2
xbiaC5l6nDe+/45vKY/aTz9EoXXrnf3SxIiLET86+gaMoNC1UGH0VpsF7Cpd7fii
lmz2ZHMZzZIwHupD8nPoWUMASaMSbOKdfhpWqT3lfBby/oVZf+3ptiTILxYeG3GH
qeidt0FpA9PLowZD3pOp0yXZNkABs/4I2Fr8DUGhu4po4wXUnItrOv6KMdLQTmuf
62itAbzOhAb+nbhIsFw0m7ZZyi4IMHWL2kV6jJMYTPamqOhpVpIk5MuwJfFIO4/t
Fi1EFfAgLpfeTR8N2eQ+49vwUBkGMNV8+DkVO8heNyjezAwFKpVE12bDNOSbdlGc
8jcyBaXfu//OY36U3Zor81bJScO6tpVhjxPcI3R/O6DtHZfJABTG5X732wLfJp2x
lyI8OM5dwa41nhRzm3zApr1EBPjIq0SDT4l5yk8l1D6w3aXGPramfT0topL7C2EH
zoSW0q2RtL1oHoNQpv6FZYSdh9QPNwtaEjKO4LsEU8qxt5jzdTuygJqmbBnvsDR2
WQ3ZyvLUzW6X1rRIvO102r+bd1p9/P+J9ezoxPLaH/BEG2CuuRBRms+LCbWkVqJF
WMnWYvYs8YmvyAaoMG+PgH93i7rj9Gm1Lyc0UaLYC4wcsytFb1fuURnO6nza12Nl
du5vM3AztGeq03NPi2INRr89R+wRNOb5fhfTRXPSEcAlJexwTomV+ke+tfQL7P3m
OBBVjMK55nKzFXLl4GRySOMYUvclFDULpIyPletMpynG9DFbD3Jjfv54q5qjl6Ov
kuzFPwdNaKMXqUpYH0PwG5s59lo9O4dQ1hmLCi9hvMMmLLiXo8Nh9sUDFyCZ45Ko
691ZNBpThimPB7+NS+y5qo+zki1EUkg22yvcy31NavbtGFzRlKn1VeTXdKYqukjU
MkWD4ztn58ieUD4dxSTBzT60uAlsUbMPwjOKaYgIMidRzwAp8vgUf819vwFTP7Jl
n3EQkGhI+KKzIxjjhOJoXtN2mfk/3SFhdsIHHqZ3Cx2kiIvEZdrH/l65/XyL3vPm
Eas+pEvF1T5kFw+sbNWhKw==
`protect END_PROTECTED
