`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X1Du+941aGgP/BqqFdjmZzMQc9D25nEDXJqs0hb6cTg2iaNM6qc9/hBwKpMHsb6Q
ToTAZ/p0IxTUcQDNZM5lxeElMqrTYNuRUXmSpsimseJnVAv5cSHjEjvtsJvVwLNP
vTM2XO/nlQGyjdcmXLeT3o8xlftXnGeJRt9L2DGglMi1qbtHqRbXFBFoTDl57HnU
l+6R0f5Azfzh/+uLqw4UsScbhLX8g7MFjdUhdOsjgRWX00pDJnoSUvy7Q1pjybLJ
XkP+uN2n55ybIagOq67gl1UNLfdm1TugPa5MDq64NvqsUyvqSqhDoAHJnodcd4G8
YcPN4VqCGYr2EpRH7eJOdnQrwYdpM//+pc8yw0mP5k9Wsznhd7KceAWvE0/Tkkgu
LY5ANOKGxH2go5MEwLtDCra9YwfyJXIT4Ni7iOVeLSHNvr/6m5nbDbcQ01E+OJdz
aVNdy1TDFpk+DuXbRJc8vC1jR609JUKRYzDXfssNj/yTSJJ8gZ4oZCU9+nIWYn3F
mZHVIJ7eXijxYIcEM6jMQgh/TeML7IkcmEITs4+dObaNSJ8dqxCPzj71/VbhD4B9
H3ORHh5wvVcw3muzs4/66dwMe87nWIBJ3LhF5Xa0nYj6otnt3YQnUXNGa+dE9mjk
4NtnuyhrpeouxxIiFQOdTEzkp0/PZl0K/IJUcFEbn4Iva2Nqf0535kKmsiZZ6pW8
jrPIQqHscl7hADp3epoetzYuzvbdnGDIeWnwy97uqS+s3Cp0iMehNxO+/26usrzQ
ojpo7p2dLrkMN45ZaeGcmRjUjDtZ22aWHGDLtHn6uuCop4wZfJ35VPKTTaZE1oNo
6wLozO6DgeZ6kzvvGmFRJMkz5SgqamEy3B3O88R8yJwE7itNkqDg6/aX9C75PY6w
HYPn3zTgH2q2VbTLw9M3ZKMho/SZxhoQzqLPuusJUIzGd14zyNL8GU/P+8dZj5dC
RumH50AKo8/dwBDLz/A1cKZOotAkQLdd9J6XYiPrNmc+BSAMyQhVCIhXbQOjHrVX
xzFhPZn1s+tNL1ROy1jdvZF5ImKPXYmJ8R0oWEimmidX05YX0U4vOBlJVs1Im6iY
IYl+t9hpdsPprlZcoTOOiaf1epWx43WOGIN3bXNgr8QwXJggQziH6+p5+3RSOdCG
aEjxnnETzzipTCaYOzDny1DcNXsXgueW2Fpdzyww+7QzkvvuiNaRrTVX/i4Labi0
q9BgJZ7LiJbCFhkAAmjvU6A5/2udcIFZalhm0sxczrk+mupBmHJ8Iv7MxxyzdSzZ
ZOo+R1OVfgrb9GYMk976Q6/47CnKyGePg4eFOLmbnb1NN29c8SwSPDZUMblL3L+k
W4mB0Il+wbElDx9YhyNArzu9qPbADCEM0ZtRu+R+mG6hRgL74ehSTok3EkTYYMQI
eJefkIXj1jbIQDscnRAYBX5X3BGQ25j1Oic+MZH2GtmvuEnt9rV3jqdFWPFwsAMT
oGS8KkRADxGXLzIY00H+k5+kXz2h5E/+bM9y8Sd5lSB7My7zA7Mq3tX3ImnwFtGj
hP3G1/ZlWtHHMbkN/AehSCqghlq0JSsHgCd7PS0cHqIeqNOpnZGyj+HRAqro7JXG
07fPt2CSFp5njoMLKC6S+tKQn9QJtSnw2UTGNRy57iySqbNTxNTO9Suub2LyUSGN
Q2DOjfdInchTdT3KaLOfSXqDHF7j42YLcsbTBlIH/BoGHpuuugWeZ2f57vmJGDYe
OJXnXfuV+iMxQhbDgB0YxPtYRy9ERGWCX5mbTMgBqvaMd7GSPfUgYeZp8+E3qNhN
iFZbkwK2GKQT7/OZC8J9TPeeA874/cyWDwQZrvMSxuJhxR+crpHfybrSBXOCQ/gT
Q6GULz/RoSD42rUEKdiZQI4yqMJ5qfN5RaxbDIsh8/0dI50q5r3RSQMlkzWBImna
JVp4fqIUP68oBElH/bsTzTX1UHcjDBbgssvCw+9oRczsw5o3ee/x0PJUr5sue3F0
SYW3DOu7GNmXBCGgr9aRk6rBabXlOTPm2bUiwSIGw8BaxtZm/zwHg9UIpt1aIceY
kMZMQNMqovSRc/tyJWE6jCO58sJ4L6S6eM/Fx/PrNpRBHfX5XYNK0ZAvWZAjzayF
wQnfPScvIC21Satil89MN9UF2Mksxi3SHDLZed+auGVG6iCZSi3+gIvOmh3Rxszf
i7Sv3sjG89tMnHen70JywcfbYzC7dylLbB+gR6FZxDGeFmt1PnuJzxujKJllm+X0
OAo2mAjqFLFmcyfmgShipWvA+LPan36okrpUdWd7dJSMuK8nKSxY2BCD9bfM384c
k9v4CN0l12BKrbYcEEuJXkBj4nAvrvR3dA4/svHoZIbhyCi1Ax20UwwRASnwiVyW
iTzSRdJhd7g2fruGXmwTRXEPhGYyFqeqH77JWcDKe+9Nn6uN4WTORhsw/58UoXgE
/UM6FJST8QEETzo98soo7U6wegFb6+SwSE5QApOe0vSBM0MYRCQBF1fgnzcxomkv
xv9ZvQjmR2JRI1uSnre55brBuVUj5lodvnUKf1OFBgT1lr0WNLwMAlmYPp2xVgVQ
si2tDV3j0q1M0Xgb0frxOYgH4LlrscIPhpQgcYZPK3qTXFn5jJGxV1zRKOj5SFJH
R/XVZz6JbZ66Rw3IbxwNYg==
`protect END_PROTECTED
