`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x/PziNrxtd+qjl3DrCrLqfzrH8GMp5W8kprWuWm2SKiGMn+XUHChq5zB8TC0lGfa
ln9HLMgn4hqMJKmdqgi6GBT/OknZUOi/s1mzw/BQpqvjekFosuhS4f/lloisMHiC
PO7mZ6MvMZrMn5ZmnRcsN/DJM9mWS0qwwwoKdSbafZANO8rml42zVYb9QMI1It1N
0tbloc0Lb4RRNP2Gs1BD/bS1TZUCEE5j/5a/dpWoaEbJRaEOoO8jNBuponiUUnc+
XdVTQgLir0+RuHkyxn5NUvZoXYUPbqALxx+CtYVdm3gK13XHKFsk33DiNNQ5IrGA
P4K2nvprQ3ueO6A2NO8IXfojdxRHihtvUM5voSCvsuxs3r8su73ZnZqTM9/Zoylw
oGTMMurwLOOkKsTMBPjj+K3YB7kcYQuBbZG7LZ6svhch1t7fsDe9GrTZksQceWGe
gUuFFdPT37H53iEzw1+/wiSfxN95QWO56ljHYa4Ih12TeMUiVLWkEu0FxT+apngQ
FsQMSNV/WTwD6/gdGXI6H4/7JI3+NLUMhfi5GYQekFoprb1DijJjLXR+tBc9DTWk
/MJK6O22PYSd9zvmL0Y9bjJkZJTdcFo5ImffrnU5jqNWDj03F2ExCPwpP6FmZMup
3cdeKqTyC0c5aX7k0A43Fvv90BILp6uR+OxrgCxGleMwO77Y1RuKvUCjKCvWlNBl
Q5AhFQ0kvsl4ruGxDI4B2RSoMOkB1SrBv75RDivRK0pZciDmBoPa8zwkGgdIQBUG
/isTeH63RLO1oEkrXkAuRMx+pFCIw1g9k+d7/FkuLtNAE6NdCovCKzkKwIssPv4b
FaGrQmWu7TEAZJDntljwaR7rFhofYKTxZ/4QRQDft6BDt+fmIVjT4r0PMYgXXHEQ
l+YntjVogVfG6Sli4O2bDSqeCCuZe6OyGsesP/teVTiESVGJRJxDxCQiMH/21HmX
3X+Id9onXaq1cOJYTHy6sxChliCADMiP2X/nuZ3rMPr6zW3b0TFTZBjtoDStjLzw
VWuEcm9Vom1c5MuAV/rFI6hqt3HIDI62bFWLZcNn2QGQZCha3eQZqxg0b/7GMTWQ
XZe7s5ckEOkdqR+2TrV75ZZSzLa4BdHt3IPi7AHtNSNCv0X5/sYB27RHJrOj6vke
L4lhjbeXQQpshmngGleBJHl9gi+WO0/vAGlPOs1rfx2Z4qsBCWVvDxOVhhsRK4c1
prGWD6bAjkqjuUg/n5V25YdLY9LOtKqlysr5EYPlyEs62tUyWYQsVCoxH8a2IrP1
3i5cq0yY4Iaa2YxJ9jn6kI8pqIF2u6gWXc2m6ajYlWZtlwJRt/orK1SSVx8Te6bj
Vjmue1tpLrWs1QLGHf9QjcC+ptDuiZxtvII2ygmrxpx7zp0jLBE/ddFk3VHxOtNN
QzIil75br+GxGSskPDSAE46I5JCCJsxuhkviOJHtQC6SM98NztGmUh10Og9Va3t1
fei2ui0R/EkjFDml9jAV0zLqO5PHQOvfXT8Y3LYuqae/ih+ex1Ocn1aIX4+LU5dQ
gC5aaUaBEfy6uTJwrbRBqwDFOhu2dcJssrBIgOvmwaNUulyLM4KJxp8o75/dUu8M
YzrpVbvOHKSgSF5kKdCk9g5gAmiEpdsd1uZTKBno4HrWMrWosZTwqeGNFBZjenvq
3ZShJTjNf0TlXmYSeRyVKD0rLqBvgf3E4daO8wNSPtFc3rKdzNRPxjxuwcLlTEOw
MFj3hYFgc9ZFSxCXh+jImVAKidiSWlUvcdNfw9o0uHvoo20VT/p6uQL4hIraQmvg
aTfgY00L/1biURBwvoqBawSjhDRbwiXieVSF8bSawJHe1HBCXkbCFmZCf+GKOtJ0
LXBcCaC6pO+kuxx1zSBocwToi4YQB4Z3/hnQY+xGU5zejziAk69fap4DsCzaJ8iF
tJJTWmOUw1j7G1yEaLQ+UVHbHJFiw39Swa0PilHHY6LZn6V48gfRUziM9TKnpkbb
5W/h1uMOFVsMaXucyRQTkbUGcmvQdt6SdSUmRBynZGwHst+C4cZjX7WUseDpl2LP
hXl3tfkt3mFMzoTgrabFhYGYdPqCnckBKiPra6PgDFuRK39oWICJc0dQiRH2nd8Z
oWRZL9HkV73Af03wb0uVHQhgkWXU78gj4EzTo3fQLm055elLa4x06Mt8jw1c8FRz
vJSl+qKNGgF1faAQb4zX4NPEn46LQjJDOdbzKmbSf6VCDisAjsinVyYmdo5ixUX3
oqNm3qQ+5bxYuhW54fSHW4TC/3RYKnAS01u8hQQRRS6cKa1PdXlrTz4jV1BGhrax
6ZoiC/nloCdpVGXiR87EAasewY2KVVTxaSuBlDuLUtv4pkSAqXCs59CjlHd0GoVF
G+VtggznblzM3nULId9eRd3mcPaJX5seTOvhPxPSc0UZE4SjT38ZzVHtXN/2EfdM
Kx1S6Ac+ICqJuZ5NzefubGUoYqjyKAJOxtNbx3UEroiD1kyhbzVAAAdp8ojqRf/N
TQvVnrI8sLd1Z+4Y9Claf8M0v5ZLbeJ/s9G3f3mi0I7nkTv8p5qeM6NaE1Gv97r/
wT/dm+ZQ0aGJfy3oIBeVFAAqtKHHgb6gbdQLsEfbf2Mc1PKMWKM/vzM0jdeOD1fQ
cbGq6HqUDvW/W0QySPu1xkWbTclk+jKhIWTUGnzot6CdokKRH/Il8sSZnlOolR+n
V90m9NbC5xrkSFYvUkDK6Re9ihnMCfCShvgr+638obqVaKzx7lVQvruXDAuug9HG
4xVSbJMplOLYwMaQroBckqXl9wCDNI9kJ6Ef2x/1fpJ+BsX0ak0mtBLyUmLlFVvi
dSkfXoDRKq4h/kNDWwSKLJGhAxAzjWfieoNR6gDEdWSfwbAwU5uO2sUqEfJ98HsE
7L5JH63lYgfhnzot3EjKnNyhjGGyZDcSMXsbd5Hq1d9wjDeOGBRJuF2bhlw9e7Zt
1vdWiPLofzZuLBMaMuBuwBovvzaVjE7UnTv6nqVfYUTihzJPtlyfBxDT9DxA7rmK
ZSzS0eMtVGR33X43wMS/jmrDhO7YDoiDQ765sIJDuZG2ukupAyljIMzZoAyBKZ93
4b1lJx2951FAo81UpvogvvkYe4suC7qFhhH8gE6z+eehTHnhNG7Pcd2xumCCLbGC
NtKhnBrju8jcxb9sT0GFEyVArAuOckU8eqt01/ZQ/IqdbP4f/8UCvsxrkon9aB0m
53LONl2qLF3y3YgCQ1nNcMpUYR2kEVoolXvwnCJ2Dlurx36MBJ0dROgG7lP146Jp
7io5xgMB/cbsoOyOOa54Ak/kQeFTyCLEGs+5ayavNhzQKuk0KpCmKTKJ8EbOJVKr
z4wIKKulQYK/buydsMlNyZKoylOm0/2iev7f2MKx0NC2pWXOebrWAAsX/jqNOQH+
e6D9YTaJ08IUcOeTX75Y5JI8yijtHhbiKyeI5yp3hs4h2Etcrm0TZyYsbN9xtb99
jQz1u5EmDZZUG/l2BYYLc+0dj6NN/ONO/i6MvRGGxYds3FF8L6YXq54o44lScxb+
DBLHP9EH2bTGRebHhMyunVgW7IbtYMjcSo0hsGGcK4XTVjl6GVxZjnWJuYw8MNQl
VebPzQXeS0pYzMCL5EyCWRAAzRhFvORo2I4NsScTfiYPMaS1TZVUR0XA4+pawA8r
LU3M/1FVJ+BvIhk8UI26Xg==
`protect END_PROTECTED
