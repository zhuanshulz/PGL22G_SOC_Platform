`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zdn5VmmKKA43VRDOLwZ2PtY9dMSi7yQ8s90p9cFWR3nBh1rFtq/QdkDaq1Y5k00e
RFHZl7YLAPZmPezGSU2t6Yly0eI0yNZSTWdHpmz/Y5tdOLyy5I4lMHiNNNAFU529
/tyRyAeKwX3okjw2jssXZY75OljaH80duZIhbISwr76kuB55tbTR5AWx8/STTRbq
baAuWFaN7gtLPh2N6+Do3kLzDgUOtgqAemEHHrJxDXZQhatSrVctCP7rhWPtu7rH
P2UubqXovu4xNDnDPG6pYuyyYCNJ74U8tRZIRlgDxPpKtwyYX3Q2e8CT+OUN8kfb
ERo/RnbxO8+hWOogKzb00H7dsBl3GeaWVziuBcc63G2f0h/eGVA9ugHyfr+UqanE
kkzDUYTmT+rDH2YEix2rGp3ZsEFkwvMvHzlc2yJBnKZQ7+6EZgqnBv62dPfqkIw/
75bSTIOdaoDdUli3OGJtsoWKMqiIXh63IwR89x0b1plhDln1MeS9aRUnbyI1oDHJ
wr8YfhzUoHoitgqtbmPyCnxH1oSUZ6OOU7LWKwn+TUgCLRuErefqTJH2ReqDHFhl
IbIgqtm2jqHFZ9W1EVcAbZbjDLyRbaqewTul+bW96ip4ES7X63wOBSYnZmpIU0s4
`protect END_PROTECTED
