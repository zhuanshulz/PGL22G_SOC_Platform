`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jaRZkXQ0uGS5h+DDv5Mw7WRJcWMlMZ+mptdpYbTwPaOI2pkJTWjMG70Y3G3nTimm
wwN2o60RgXl/mFghl/YReYo2KuLSlSH3+okzdh8XvVXzpzqcnjdOo414a6U/MpvI
ogsohRoMbxJNkztsDN0TaOrcxV2RyvVUd8zqHb8pD/t12zrQZ+3RS/SsdyMVN2hS
g0w00GgVy3HyXsqQeoWGD+zxG94UXqoMIu1Nf1Jo1HztS/gFiK8clhzqrXYuIEgz
6NT/IE4D/2h6FhvUjfwlcOwOISUU1x0J9EOJi9LLTRz82uG9xvWUl1tQZPFMQ+44
lbp4G2/Vna5XUO4tvhs1C5S4kXrU76p9BbObVQ5M9tkITgqRdDhCZfmd8KcJYRfD
E+mB8u4g8xbrlYwAh1oMbDZ3V/OaftHDXa0y0SJjHMiZseRTBdwe9EwX81xkLCmB
22+g6C1zlXRRQ9m4jFgyvfhDfYLzUFiTq1rRyM/InAab476GIV9zoiDIAbNj6Vsu
+he9ll78ExSfau7MjzvYPXjpDK5dcdXFDctIj1ZZLxBZwGSvJrBBenSgLBq9AtCl
oZ4hXi6RNt0MHHH4JWYYVSHl0rzj6Xygaw2fWfX4u3wSIKRCzEMHc17FORc4bj1P
0NEzCkqbidYMlBBza540HiU01SSObvharMjnW4mhLTkrO8WZTYgyQNWX4DWvLtb+
c2O2dJOlCVFXwFyWMqlJVyWWNhzB9HGm0xZ9BGqTC8BGbYuyBhYMueRPmd+lndSM
tHvZwv1cRiYq4dIaOxkThXc+jdOxQvfjNfDNawH5hGDeApI6ZrFGb2wYWg9cOiBQ
5S21Sj2F0M7txh0uUkSHeSroRUgh4kiiTtWKTwFrmjhP/1Eo/BrYvHpnk0u/r2ZZ
UkF0mIgeUkaasE5wJQnCaaJmrhBAi1q1ggt5exUtLtC91eaX7V76z3lOjCJPw9dC
k0NlZ8LRwXmTcSNp7h0XACBR3sEFS6A8QMB+OMqJ6nWAP4YZ0qo9JZNzSAYK1736
puQO+GzFtqTtpzxb35IANTdYrrqOxSZjav/egFFTk+ntmOo3nm8BhztWU46lNYQA
hqgj0PpnMtXOV+SOvYjBapPz/Yp9uIP2KqX/KFOoDfbdXmezbx7+FAXliIs20ubk
dMDXwSQGPofrkIjVPRza+hJZ7Qh8E2jpPoDmPqxPn1xLDukzzxoVevuenSoV8Hox
K2w9Y8rloESX8bQAIblM8q1DRGFWz2nGPpe16cZq2gZ6UCbYhZRRe9JUdM8ejpNT
WhY81ELFZCg9yNzknaIZbH08WX29ZhKxYqNfMYBLgW2jzz23/70AJQF+YD7oXyUt
grGED+o/vMXtskowvA3JlJL7Ab9uqLZzycQx8psgSDbAChrcChYK8HunfgvvEn2b
0XimoXcXjhCP7SX5A2pIqEfuJm55ylH9MCMjZDQLBYQ5PGCH2Jc27d9IZytzb6wS
bkly2Q9BfesI34tdoh1f607JNSsDVUQngTB1530jhRzuAFmw3t9nqrMAGY/6TwDV
ePm/tDoUcj0hAkz6C5dfZerB/6RJMAWrNzlQDNcS8jI08d8E8htiCL72rbcJ9yHS
b8pblQr+bgr4FJhL+VOvk7JP2JlnBsDNZxHwJHvSLj7Nw2L/BPq7KYE3Px1OU7JN
WifStGbvKMjNecA7XT//pT7d2RZAuP5hrQKHCjlc0o9HrNz+c3ONTUqZXFwzpEdy
U5osA+RWjtRUQFF3CNOxX8nFe9dzP1etY29exAUIYjufuhiI8AjTE6warHwm1mn+
RQdCmY8fGxI3EQ1w0k0Fb4xD7ni9Nd4vLTZEjqKA0mTkGNLVvrEmCa/AGdlP1spu
QKKedUk/IP4gOK1XZOu5mV7vs94ZVkMrwau4bxyQ8fwYnRTlBQudIwaHAiO6JGGT
M4qwWr396NxoEL8jhNLjlDJaX61sQU3GqDVkB70KrPoB6BBRssVRS/LEk36sCQUl
ZyX8FpcDHEJgNkgj8g/H7H7/XXN4MCv+/MmPjo66sFSCmUk2TcgpsHfEeLxo7OPJ
fsYKlHVeZp11gKlF4mufdAvsqlmz7PRsEtg6gY+YaHtfuxWSJRVDxF/v5/Sqk9dp
bZoLvxRWyxDP2+EL9FZvmQf2+Et23fcb+eqkw/EebSvAhH0FT85pUvP6olD0BT0L
/e6SGseYuNn+7Pa4gVuuBPPO/Uysrxp9IoXG/wZSZGlvlF2BPGwT7yQxhdxwV/TL
HXU+xmxQeTRAbCJRfWQiaJEUIdH4X6zoEjCbwxHGbax3ciS+6XdlvMI8VDiwaS2c
oc+hkAE7zJoPdDObVjT/8Zns3pyn+2cuXKJFdAElaIMeiJwm17NAGrgTjClbNAW/
FVzo1koIldclqdXNUv+iVoR2IM+tusNDqx+edJz1/XgAvlUjkFa4xmEn2QFUFZYF
2QZo5D9sD7f7fir8//Kf5gcDWxER1JGQCwhUjk4qcs9iwXIdi6UBhIxKCfTav/GU
31voc8mTCfH83ZRIq4F5NweLqVzIa8VThZBr13y8F9a65PKSRnSP/CyyWw+X2Qzy
yKsJc6kWa6oWmX9CA0Y2UGfm3D3VVsHheCP8kT2PSy8z/0hBgVXhga7agl87D+Rl
8sv5pFQV62poxBcz8ikVQGjtQA3O0t+uZSzhrCvmbIrFAi8stJVb1fzWLlaqJ5wl
Dc4bivKJI/bKgrWScG/5+fbw7KbLTqHGzXEG74Eqgm5pqSHgSYdiP6kj41BcH1bi
kcYoynskFxHycODilJMX+9Vw/yN8flca0FuYZSFZTqvKoXuDXwJ46DEQlRzDRmV7
8+A/kPWr2NLsPFMidZVWlW7NGa1V4WROGujHx2bHz35DCLL4jSTNSL3n1Qg4JkIH
NpqOuIIk5YQU4cUOyA7BXH1vDtUR2Apqi9cIsqPOSPDMZz4qsbHaao0+moqMrcIU
4jivNDaDm1OnzxogHZHeczWJaMfiwDTmgbjV8NHjaJxCaQ3AmjzfsanI8E9D8ccT
4MFuTxjMtULwesGUrdWux92bQBddZ0lkxpI/96ZjM0WOAQfnYNLm48+ieKbL8oQP
XosIB/MUV+V0wo4Wk44Tmu5qzHcrlvNCK6FLEh91jffzH92AtT61tjeZQC+U0XKH
nHuF5o0szf/mgu6y+F03uWmPS3Kh3swlUERX8ksIBmteOYaXPl7/kYJxVit0UZOa
RTA5QyiQ03sc5cJhFm8vPVeAxZftNikjkbUZzxxKhMfWsdmvJoW+TGD1eiSFqJ9a
uMYzyWg222BqcJLENvr2EBP4BADcOZa+XP1y05KLwAzDi/OqGLUhw2ZuMr7ghm/E
lYr86TxFU4fJXTWESfI+uqf8OIb3Vl7rEkZcTgdwbTYGVxWWEXdL8zMqIv+NB3Zg
CC78Q60GFRpCRo9lZ4aTv/E3/1+8HupJvH+4Vc1j27GHIyWlMMuWAW5GsO7Wy7HX
pK6lTsKTAiBjLiFOWjuvanMW3Rvr1/xjx6Z5TBLySIur6Hy+Jpiu2hz72il6/pVt
vJbov6cjwHm55ZlXYRoq0RNuXoVxcvPioMTECJaMxngsWhj3FXRseHyfMnRpOd/X
Da64SHRgalCW8Z+Kk21ScUAejnxnDjwPkskvZGTjP4CcDsq8fuBV4KyqmAfr3pTI
gjXT7BV/zYmVHiPTOWRsQGItDcW/ph62UrtaJdQhkW+u/BC3DHVBIN9+PSy2vIb/
qeJud5ZBuoJzO/iOcf3Xt/m9Mf6CFYfDJM41ARMoj1jPp2Je9yIOEL38Uu4Suedy
csL97Wpif3aUXRuVDOl/MtxbObJtqE8g5t5JvG/uzalFbET0fZ3Rs/i16J/ZFZX9
EwJtgoaqvHMKQ/i0ZMpKy9G9HPYWrj9YL1qWK9LTpqawgAB5xt52uD6f9c8eAR2M
Wpi2cQFVpzxU8mpR3MvrI44T/2oXkfcIoow6DUlI/KjoIlrN3WjHDmaG1KeWK6X2
nOiFaxCYszmSudcQaM4wqQ==
`protect END_PROTECTED
