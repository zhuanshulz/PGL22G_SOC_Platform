`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KWZAjp+bxFrTX999dP5V2rWGOs2IsD8T4JuDSnoF71vxpHSM5U+hQvzvROivmRoa
53KBPb7V3fwtaTsMp1h0ImJYY6vCvqMdpAOJYy5hqZ87UbMaOXih2WV4phdF+swI
nBZCqooRd4fxzym3vPDvTu+pBETWL6fDybdTouycxdfEjFYt/bGGpPrXAEDERGgr
y0KbU8Si4dKCJWhirOj86JFcS/7O6spj1mTceTMlr7OxswJIbJx+Y23ZmjZVJ05j
8BEC2w7sI79kWygbfJ2AXxy29bi6GEmkC26LNC5X4UeJDwAWtp4J/fN+GeaBZuO1
1gANyMK9k9coVnc+pBGYxzXWBJI5soboUqP3VG7exsYcpt5t6fZ8EuyRzmlPRPIT
M7EAcqg6f93eEEtYgsjO5X+aq5Fmkow3/kuwA9v9sBMmk3Dv3t1x4TZP9wJDDYP8
Ax0oC+YjexpRdJDC60t+azeEH7YKAN2t0Tc9UFXtgxm928nW6yW7eLr0Ag3Y8fSV
EbIAT5380UL0CkIiT6eeFqwImAAUXj79ZbftRDLeqxrUewyXMpK9IDIQZLgD4r8g
MvGNRGolpKtD+GtEzEVNkpptt2JdQNdM6SP28cGxrDd1SMQvOnSiEvwi9gxLjtyB
Lz5zHu/TsqwxOdzVqc2K50qlCResxHOXBrYtDM9PwDMd9oPQmDF2O9gCPzmcdqsA
/WF5ZlD7hSKvfJWaFl5L9HyPeVcn3Lmuven8dWCVi0tAVS6OIJjXOtyEGxX5YIQs
oCO0Bj4J04FOZUkkrBxZoptGHktGl58W/+U2+HCYwRVmQtarLPLM419nbptnknH2
zs0113eza/6PnRO7iyNkvBuuxfuTFr5nq2Qcma330NCQwXEJuz8dxRQ5z6h2AanT
NU8OwkBf0GJDOieUKKVroXNLnJWMdN93K/gONdS78ZAoCjXvoEBCVvLr4jG0Yx8X
CYdaIHyrO2zLX2R5sBxbQFeMfIag5FUVEw7UrdKly1Rpy5wx1/jctjIovkc6xlJ0
`protect END_PROTECTED
