`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hOysrgtHBEFkumonD7C4jk/lafPEmBDc/8y3efI2/VQD7m0u2bTKX/hiy2CQd6Xi
wUKZU++ve2U5AQXGRkhfMvLf2Z4WSKLuZC2VTzfFGrByI/pGnEObYq7PFjB9RBFb
411zT55nCp9MkI0kD+RoGQ==
`protect END_PROTECTED
