`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4kSW4Ju+sVAAZlE7NgFpyaKDZk4Pnh8vW7qVyz1lPLcMpS8aNcsNSh2BqGEPAv96
73wlME3CuymnXE8hV+ZNBWeripx1Ikk3fJ3RcW3V2CSSzLqQI27V7w5BsOmKz6Ls
beUgOKgJD893ETuThBgKC2rjrimIbnf377S/GOJOccoFNh/jfmxplxQFhFMDeMPQ
Xzr4EXTvQtZ/dz2nOx+Xr+YwMekHqAYbed1IPp2238cVRhKouuSBhT6peZz/Zdyq
2QtZX5Wp/uQUNiMBV5mtxy98tO3vvNmExkpWu3CSjl4Bitp/PlPseLY6CxpE5zFz
DpeHvbruoWWuPn0/U3r9hOfEepmnJ2FZy5Lgb5rVU0rawU4zbZ7x3b/btDNHmypS
NRl0lFwQPmpI1s8uUCxEr8ISr6DkhUdeQWZjFsrpO2hjhtaaNzBRCbnsC6ZWqXVw
rPQq34F90C8wR7qKX5D/M9Xfx/YTybR7dsNuVPinw4I7HmBFXoEXhzZJBNgZCsJr
EnHKLrfOt4FeRrrajDqplYQYORUKkWzCM6RkwCUp/iY7Gvv+YPIGduljGa/gXafP
aG0QXsEVjdNjZzvYhwl+rYvdCUzTbXmp/iKnfs70SsAkC98dHAYGEToDPwk1uE94
pIK/cxypvpTXBpKu/qmM9Ytm/qZgniBdXKc9U6VOU+tCMDOvRRIRlQh5APwD92AE
wUaFoUHOl/ax1ZVxd10gUZaYTXjFwezMslZz7SrUB8+K0lsTmmUaNNkrtAOvL+6G
KN77nXGr6vQJ92sc8Fx9O7X3OBJX/l+0BIfqOu0kUGt9q/nogz411qBLxgibhT5C
kyHdclgUuocV/ZiLgIJdASavw6OHh/Gtb6tmJk/2GVZSapnt5GJQysqk7RZkiDN6
57vsvwLTQKH2qlzWGp/jf6U1h3fEjpTiOqMOUetSxiLCeopuP+Qj4LfL38zaXZpd
dTpVsu5+WN5LF90hqZhNb/m09xH5bNU5Y5AHYE//vp+SjYHkCzgjuc3zZzc+ADcU
4ytnlgUPhliR4zlAUBPa0r7obbpPNqgbSQb65IbnwXQb1+APYh+urVGB5d5GCY53
w0ksz3w4Bo+znW01TDJAdSUZql6PSSkhkKSNw1h0s7ntvmDmqkzenwCrghq3qr/L
XYlJm9a3sfk08G8sZchItk3ugcAef0D0zCaN9wl7QEyPUH+T0ww3Az+m8KJUIBxl
OV12wuBACTD0CtC2hPhMTC7t+v9c6jRLOldyhtVoQbjbyy9Yjbj6udGnaYebcS2U
VXfoXij2ilRjDb09Slt8hKIRuUFYysszVcXu6k4YAR7sjxZ0hXss1Yo9YGnJFT4O
q3ioAKz7O5uzrOnw/Q2swxI0ogGmVGMtoKY0bKi+gJAaF7WgrA4eCm4Ij3Qx4Ok6
LxVdv0bA11oP0R/JlPCQZ9bMQ/NWUhecIcU7L4t2YCaCVg+oHEAyowqB7aT83Gcu
y3eCEX8lvcAIrL6AEwuyPIxfA9QAMwXMjaOh3Z0BWb027KblXUYQJ+QYY86hFuvr
ZCxjjDbyYdZrgFNQajTJLS1Lxt3ibI1NA+izdElZj3PsnHArBFr1FtK8yeoZDPl5
/Ij4xLEQCYS2EomCqOrBB6H6Xq4OR4/DZrg/lFzrM/zDRpDt0QAkTF/LHxHktfYO
mmpXyq3Y/xMF9xoFMoTP3iPHRZINCVaxhe9p5DlVfSPA2qK1WBiqvqPb7xDy+ver
S076hG6mmhbI08FCYXXMmDcXuD9Zd5tdhY+llAWG8brkW39dmKE99+xfZ86D1k/V
aje9uWE5KPw/fdQoW1kO4bV5OWLV6Yc1/PGRBKk+vG3TaST3B2EISv9Ecxi4jsjr
Y7SjUh9hSwfDGvfY1/LhASzkoKWCOHVd8nD9Aj9bRqTz5VI6An8/NWO8UFt292Yk
P9fRR3zegEbjoEX4ImeCwHGBi5nSTQTvYCx7HW4iQXwX0JZ0YiBq5DKWRyi4PKHE
pruRe11U7L4BZQSnY0YEhj5yuNdKNUpvehqoUpNCbv803egdGlsh7wxiSyysO5SO
Qhg6TLGxnp4OSVwFr/SRsvbYU3xxH54oWvuNvObbIs39diwa0aaaIruKv+Hdacs7
I86ZWYi4dQR/TRI1wxi/fpu6jGi5sOCpFXJ1SePAQm1mvMwNvnanRDZ4ZhzLagfu
q2sSSPxpYQdklUJMcRfhW8xgFKszkCIShasfN2G0NHoF0pKLXv4QjJZPfzAFmT/f
ITAw5RZLJc/8R77n8DPr3xDbvIW7osiK9kFE75VI6HEMHcI+Odug26nLFdE/2E2q
NHB/LbCmbcSD1Shjvei6OWqX++sHneeLVJxBBdkYu+7AERm5tlvVwIJJPim3RJZr
S5d8yc08ccXqnG2Ig1r/pDWcIdPkGt0qTUcdzBUq/0NvmrVoI5y89DuqOCFOLAZz
OAPVSob8p7N9KoZp0B2WYpjkCYC4+2VUkgvK0LpkXg7co7ZpuNTC7+slpS8Eq56P
kM7Hw//yWaKTumRrtWKlCdTn61djjt0aK+fejyT76SS1yn0UH5ZKo/goDDjBpobm
+l+bt3cvgK/9g5kgys+WkmuYulxpoknX+1I838kbIpDbO7ElrfCMIpUcpsCq6S+Y
+x+aIrSblDfZdXxkfQgo54g2pRoiLluaVTEXWaoCAasQ5jMdHdwBXODKHMkxXPQA
uQv10KuWD6Po0Boj4YsCVShHdHcioG7AwMGFRrhr2pCkBPiKhMCshY5RgV/Uslc/
UMDTQMPVp3LcSn+m37RI0ZByYQAfkgCesF9tmIWyD5ITNsUEnyoPk+VFoQGyQGyF
SCPHVka0qin8DNp3yG+PpZSQ4gU4Ygn28qTCW1PwdeGgdd4itwGXqM2SdkoHRNHh
7hKzTOD2lMVXTnZCwNAXznBIlTTTaCrgtVTmWKc+bRuWHLkW1spLs4plw6qoys6w
d9CsVkpWfXyRU5JTp04JTiuFxpklae6oKdYVSVUYqY/SF4t6m983CCoGzSGFx2Gp
T0MPGKTHoaCF/MHHVogeQn9UOdyOUxVYfBZUAM1gZIDG0QjcolIzpQqxVJPFvvwN
TcOLl7quR3+YOuM9sjqcwlr64LjjngDk4M3LMqXo5i7JJOwa9pb6+cbaVqxNrvsl
7FHD0RsrDnaByIR5P14a6HgH/P1g0rLPHn2adDEam5S46oBUs4VSkTNISW1jcson
y7lLawHUqBd8joUEMkQ0nqEtIFcFVswEQhhqzG8t3ep1qXN87lPK17/e1Y/IBTPd
14K3O2KMjCiuBhcydfHm6fwyrvVTYyWHRrwnN+ie8gkGofVo1G+RnLocTxdzCEr0
K8fxid4UPIfZ7rSft8MBPYoo5mdpTnqfnEE8M/Xpka7htwY6F29BfP1LzJqnZuKY
Dc9YNSJIt8goarCE7y9SQUql1khK3vtzwDWqXjyxZT4ZIEZY4F9Q89hqD7zW/LJf
gF7y1M5xvcW6PBCE+AS5sGjlp97+167Kn8tJ8rVh/ZlGP12JIIN1Ly7g4uuGsSTx
iVdpOjzsC+n5yeBoEAzkPgpACUyNpwHkqTaD6NAR7kgOI98gSt7K0bGGxejMzCNY
s24238qTS/hVaL9ZoWPXMQUOQta2EGuztpIu+I/748UHlJkh2nefQoxIMgvin50g
hCi4vwO/Q0thBlMH32iFtYbaZbsfQGBmjwyxZDQfUvVehbCnJoaNkm5vFwh7QRS4
4OWZIU4HHcQXlFo7KB8bYsnB3rVu/ZoxNErhHH1IO3jgKvE06udHN9u/hUhHanbU
6amxgvFAdynQcW1uF20LjkQqcRAY/5jGaEPwZmyXz0JujGIQKy8jgML2waCuQ4dG
JDN6tfiOFp9X1D5J6o/hSM7tBvR7ugvUt5bfVsJQhQcchZ+Dyg7zpAP1yaqUw9Za
BJGf6G3bjmayPwAv9A1TR+AXP5lqGifJkxcjHSb10dpmm2ADY98nxo+J9OAglvxj
j13t4cSv8Dw7yHJcGYHh/yp94196hw4k1TUFg874MwGeE7Gc3jJVV3hJgbETkHAt
8gVj+0T0HU/qLX2vlLbp/+h20mq3VTDx8mOwtfjpK36fWxnZNb2cRXJQjP809kb9
Kb34hn/H7O52qEP7ViAtLqaq7QMle2KpVKm/SgxvqUThxgQoMeuUMfKCk7kR7V5H
OMyHXPVX5/rN56odVrYWW6gFuFnjzUZZU9a0QAu8chJob0amF7kILClOESnMBcxB
vkcsVCDpWjo6VZMhTyDxQcZRs/Y5D1qbtNEd4UBwRRG2rvbCve3dlF155IPfQiIN
A7BPu5CFsjkNOjjRqMf4lwKnhIq+lgG20FFBRB4okY6wGfAoKNI+NYe/vJGQ7Anv
zOSHNmyvNFpS/uT0Zy6CPJjPkNUeWeYoyEkQGpAx2qTtnlg5C1Dm1W1CczbrUkVp
MTm4vexVHLG7iPn17f4KH/h1k5iI9sVc8DUjExzOAEpNb7SFwZWzHaaNUn78GGhL
/NxKAcy0HEVK0oSjXMYY85XfDeCqeKEAv+v8Ml2yMM49lNoqlmbY2SLF/tvvjso0
5HNeO9KWMZL80xUr5ALW24Dmg4BonmYa5IZdlxOZiWvAcnBV8WGuvpgI5Sla2sxj
zBS8tb+SDIZ5WE4+f4K9dm6NfH2l+0UDebtioDbNutopJhikN+kptGyghG/TAnZr
rxyF4CgKknFIM0r2TtxG9vXb9WCXl6cHvLeX7A598+41ATsgzKVdWCXJzvriRzFt
CiftBoX1kRK7n5Ih0P5sV/oYkeSUN+XRM9lPnPGf0Q3/Zrkcu3dvSi6ovdT+d+/k
GneKsvGv+Hnu872XjXLBCtE5luxzVYDwxEWvzTzaaFz5GdvDVvLfVR6bAu/DkbZ0
I7Fu63HCfb8ngxq8zE2fT+2Q7NN0e+Lg1TH83LBg2M6MX+3/XdKZgqX5xNFLjLTb
xy8xbtZvVrxTks0I//LuKye2aQQcD3kFYnRT2pkuiKrhGTQdby7zgRLOERJDEtO9
dixY8SANY/Vm0qXHO0U4yp1KzoC4p7+Ql84i999wVMw0B2hN8NrAWCSu9mJbyzSk
55K+cQGmTPOzpUOtmMlZqAcY72XHPwZvHrHgL0WUuZ1krRolIceoD7YJnSnFYqqs
zz9NOLg+YacU3moyfBvjoXE8XVVwCtg7/TR9RQCvyqQpDyh5yCgiFJBBGrMNY05R
YT8mO7tpRyO2mNfEztDU7CVFV9VcR659zzbm93o4Rj9sY3bUxIs6uprbKOPvZ/st
CtG2hUgmGg5XmPL44l+24ajDPV6QnCAE1MfdnfvjXJykcK045RXcoX9QhjROsosR
2gFFX+xjN6uPRLGbbmcW/ybIYa5vqxa+rtFqR9Dix0Yx3C3krSI+tCb5zABy/jdM
HJroaufVy5s5BIPgSmZZVLtjk7/PT3eJQBWbM8ZXHx4YKHr8aJ7oBjCE8vK7zsbD
43qY3PHKwqNTcST2j6fx43sZD1pURSAK690EJgO6Xkc+EM9Yw3tMkHv19hO4JTsO
ex/UgYkS0fmUQjKUAVenAhBOey313G4+85csGeKHRwFTc7czauNdU2vQceVPccf+
IS1GB8pt6f5E6SZqNbUiMS8SVrEd/IsrqDdjWLWIgnepLNMluAayXzscRWvmAURV
5PWnV7yCJc99FQzB/iAciNZpUrBzBcmtJ1st1H4YHWWOBQkiUtP4iQyaEbQ23wlf
MwDvRjNtpGy47EshTO4UpVc78UevvDc/wiyzk2fyVN1xyQZF6Ls5nc29B6v+uPcT
n13U8xx/9nJIL3xir92/Nl75TnVBtI9TUuztatghfO4gmfD0u6NPOszRwnWAuKB8
0vejcJ8mAAlHAWCC9XAYdhb8vy/aCDRMh+gLhzfjpH1mamgt3dNY2TEq2iHocncn
TvJomNe4u0O1sf62Wn14n05bmyvMIDGE2FxHBYzN+xPWuSmhrnYhuxOCJ6dQ741i
eWN7cWEuzGDMp99mnlbSI6V9VKlwwwO10ciF47VMvgDm2wWDQ3rcbmEZ85JUM8vs
VXg530KkgTvLt+0VCLHHtbOcwupURd3o3hKkNyAuw70S44QspDBqHMVRWosiTH/V
M1mHdReIMTRK6kv2tHSYilX0rUtXD3qfV25atJe9jqg9GAr7AHsFi8oi+J23cIs2
0z414SKYYFqCwKDhkC4N+iSFZ9uTH8t+LFky+nV5OfaDKg0AJsimz2NIRMB6d5bl
MtOem0YhXUxU7OQaGL32cnvHJKmMcI4asnessgcddmJrcURUoT2ThaLZvSUr5/L4
f0BCujaDH+y0i3dMjI5VXSX0ZmJsLesv8qCe3f/326w5x1IuP/+KqpNL9BDSx1z1
r6R5Jzd4pnRDKQvB3jy7P5XgDHkthGawui3emJhHfrKIU2fh3vN48a5xd69KIok7
f7tyUuo6aE+OEjZhnWd/hUw3ppe8pyUSqzLx98oaYHMaXK3PPVIxBT8F8A4uvbd8
RCkRTrBjoHqqTZktuSLPjISrXTKpSXp9m2Kq1oUTzP7UMarvjqDzTx4Qll3+97Sn
Md+gxzqP+GgoOqe1rx43ThQA0Hj3qTwMfgHQK1RAUwjY/FMW45WFLDgLZnc8nbbn
70B4Im1PVcvH3yPJD4FbA0AJchLj3C3cf84mc+S+v2+aKafNxhssEiRt0FK7EVYF
RDFzBlzS1KLvwJcyVWArf45Ju4IOvo+iViOo0rcEo0iJmD4L+fnjamf/kpI/Qy6X
f8+ius7zuJaKlGsFYif44r8+p9KyyFoGyYdgn12WMriNe9esiu5q9hYC3MDmRRZ3
aHcvDJSediQXSQeGgQRyWUjFnxzh9Yu/y5KYHSKrA8CDzKCd1TG15cXxph4YJxLj
5/3uysWiKRK9CreXkM6CAgQOiynxNoLX91nNi+b9rSBZiZwM+kExmPirA5UZCVok
LBckqh8Dddwxp1k+0/SyvaRccqn7h3aarqoExS3RthndfN4kJ8iVDkUWM13Lw/Ij
ua50bzvUwuC4Kz5NvrlIkOWu2gd1DNTQSMHBh2IrdRJZXNmngN2Fa0hWlL1scnSr
w/NfGy2bmnea0Z31WfFVN1yCwuZG+j/kqv4xt06Yd/0YeXUPpy25j45voVpdJU+c
Ogwh2k81DuR9WWZ9TtiKpFMxYkMuBNJ49Almbn7cUkrK5mk06gFu4IIio4fB2dsm
WOaB/9EoVPK7RWEulgURDhrq/+CJXDbjJ+c6PrQpxQLn9c7V2OdWk38jdtkN1zvE
xUJ2N3VctFyjleomgBZ29FSmLMOxS75oVY9muK6chIfTplDR9CP90WA5AzFzW06E
KMTNHlBeeZgiZY1FfTQTeYPbjKmGyJGKmszb+B76ksT4AyE8c1Nxti/P4IBOqQqP
Zx0FBiYmfdppOBUYE5nOk9/vTFTKef7ckmk7sY8P1KkjhnmX1yvsYJ6Z9ce3LG8O
Ng03dgLQRGQWu2o2tUREjBJEKokjkRJzBPcdTL3WwnLhzNh9uM4ty1hYej1qeIdA
AzoUCLhreU5eICRG8Xp+/v8f11XhfXzznnZzGUBJh4q6+MogYY0/SkGwsE2LOzAS
bwCs8zjaZwXOeriDtNzPzpODuUInigIfq0QRdU1Kcx20udBC1SJ3TNruJXjOtjfQ
nXLK6lXxE8VZ5PSSYowvMiWZrvISCe2IAnDBdlHOonHgeav0iQi5Fc67wDIRVR1J
931yoW46ztVK1OAkITWafjXWsYAbBv4QBy/NXeRTs0w6z8lbE+ZSScBdypXSeFEL
lYPK01uEVRi1F5KlNCahKzA0O0r6jvNGsROroPVVOZFz9slbDf87qVRTzyqGuVU2
u5kuAhKb0lAao4+r5AugM4OH/4Mz1Jg9pehPib2u5yPb+aF4+n9ejJraZh+9Ih0y
QY9qLJnDMbCArX8N/DyXYCZMLCY96Wi8ifXSQyacrQTiWXVThbMCYThyfRCyozF7
RCbiQ5H6wdv47FmjP5QjG5uvWYaI8kr7NjgsWt8VMxJZL/EfAFmiiAwF8tWm6h3Y
q5rm+VG5Q5zkVG/ubIYT11+dAROom3Kv+vBwxGpXPXBQ6Vr9gDu3/LdjZ2sgTRdy
Zn3QwMr3PXK0eD5wjXWSVv4dxd4mbd9Dlj3JDyQ7kUFjCmlqbueP/guH/aGEdNmE
VOsHNUNO4zu5tueH06dhFHMLQP1nn/fsZSGW9L7X4su3cSt3wsU9B5cAX8CmJZIr
r72Db3020diIb8BD0YZnCcJ9gipwS1QBqH692OwKCVK+HExymTvIk+v6aKhJB6s6
CYWcH6/FngvMbguxh4PFMhA9XyAo324BSew8Wh9YF4b6i81NuW8yJ/e7v+aUm4Sj
rOAZgTi+1ZbpahNpWLUYNloN4PyXeszABxae+fujiJ2IQpAsos/ErkIK3S62Z9tP
KwTWNpITiUuBZGb9AL7AcKFQX9lFhh2VcZHM0j/dgqsE2aO7QlM5YwArb73/Zoth
2k5/tcEUtQ+qJjtZT94VdpgdJ5d3z7BXSYSv4CP/awn0MXJmI/uWBnJwOIckGLSS
1thP8+/wTljvickavvuzAzlquvxQCXAjraIY3Wl8KVm8ig1R5aHlclrSXzvx+vFH
f+8ft0MrSuJBpGH5eoWStXKfiZgKckDKdgiouB0M02OHivnODw5ySNrs5v3d7mJu
QNtjCAgdBcKAsuDbNauq8bS1/Eyad/jeOmLv5/furfjEeeFZsyW+E61NaplxbJfT
XtSMtBaMEo3ub1eN3TW8IwIInfHRoVZgrGFCvmCcmjnvvmJpcW18C0JVHTFT7xzd
0BdMUtNZh2RJcoxhMePHWT0F79JD+1pjc4Jnhx8WLQPEbqEm89RguozbLlDAjE70
e6l/+a36WN+EpzEl2c880s4iXKfHtzVS+C1/6pORn1rHX7Q0LUvi8yGvP26LnDGT
53d4gcGJrNxkN65MwribXy3lgjSWPyoMIYNVNrCn500W6zziVyr0JuH9jNjFdfJi
WEREi1aG8yNypXbiou6Ld6g3YLC+VcxWAePnQZE5xMKIrrCnAhQhJjCqmMCaspyn
294uScVrv61h/vewphybLWZg1tTg/x/tYIovgQwLkudzPFOHGr5MLzL38Skrax4m
UhxP/ETyQ2jNHPz+DSzNSKjwLK3KwBCEE+/vNxIw58gPxYhkRAYTk09nxOhSlVGc
hEDGJ2aRP4EXfVwhhqg1ZCL/ljjkFEcznZvDBH9SNiMOtb7fRm1SRMxsCAJAt+zo
hM3r/zJmFHpeAdm98+77JoZQ3nncCzMbhzDNGTl4X12gCMmRKA3Z0e5+i8QnM1Q2
ngKgiaKM3s/u1uYMQPznwj8M08u/qyZ3dMPS6tn9kyBXIudGw3DS5u8VHuz8tH1F
F6taY9wtCkkOgCtfuOC6uuBM0HfKGoIDmN9Wl4Oq7+8ngyxjzq9EqFySil/Gj9l5
yxmU6GOygT1lykcpnadDE5+0WaIDLYSrFFJR+DmUdd4T4YM8NXkLZjuLJNlo5nQh
bfjAKvlmayOyL3NhqNX84R3IqB/Nt9BKd4sCncsOPRkTHWTryJJ47eWIKsPJBGjY
CPbActx66AR7LGYUilIuwLg7qBFbtT+juzchTCLYiyN29y1D2N0gpEdl0dK9mfe9
Qi0oakmqgpUux4MAA2DpUOhq1+DeG2nZsFrq4YDyXgHn3YUQfcTd4o+kjjDKg4HG
VXCWvSQTlN/lqzE/bdS2WzIeAlQBdhlbl4t1bIng+NhywswOFhu/e0BddFmHKxem
hZqAktpeT3Z5UcIKo8h3yziLDNASCcPNp/PUTSc4iXoyrSAXAn2+h4V8Rgdcncfv
/3r6PPGp/LZutZF4JBRW8l8qEI2TRk0883fNlRwVJrnnRQKZcu5F2yXJoC1UgjEt
H+kuoUFQHrauhW1v/1FQ6ZLSVGW7GwDgF//MN8mYIUHAdhbIypi1xNu/TJ/YwMyG
QgS2t5JXbcRB9QZiAJR3Lce/MkQfULG5cZP03UJfwL3s6VOvwvBnzrRa9MQ5Aouj
N6EtErBkmP7Q0m4C6gQeddXZOSnW9t0SND1SMdBfa7JUSmVMigkxxBgQho8SjXAa
3t91vYyVBTBL1dh6uqkC9FesdzS/7dz4za7dKcTGshWfPFLD0cXQaVYRzj5MIQkU
WZJttDlOoEh3ek9E9VP673O+Am5/VFsguPKzoeqzVuq8Sqirp8GjF0wfLygkP6J4
v9vQIkgPa2jIvfnHSwG102iZlHdT53jmf8JuONIaHICAqS0pU+RL3aEknCcrENL7
dOxgXZcjfblqCgTYwPPNHJ375JiE3IzN09XSrw3o/vhv3cDvtxguMYmauZE/eUO5
1wFqEPy6JtjaTimbwYVz1Np3HWUcFJ7lkiFAErbdjLzKHXoXVcoppBaAo2/oxoK4
MNt87047R+Wy4c7uOQJtjoeoFzPWs05wl74eitTltOKfLe4gL/xCyyPl4u8/Uyw3
+t3q6Y2AC/p1mutcK3sGZLPVtsoX/1caxtfYehcoiNR5v7j06QHMts/cIqFNTEu5
F8cpofXGP62MtT0KU+AxlydUXGQjgHY/fScwBp5J2Wp7fx+xTD9W9vbUZAhXhCtE
b8Jem+c2BHqn9PYG17pbdVUdtzHe1JnneYz1smyyzxzua6ZyBDq7WyXZk8spKwU4
HGnPcXkvS2+SbZpcY3cuuJ72f9B59rkM5z5IRiY9Wr3MnIFlBBQPZ2wCi/o/w3UP
xFTaKfcpnozqhDitgSPrJHKv/RyoVCGlKCOLYX2B0ihHksofZfR6KmTXWLJZZxtp
B0w8ER39FkTiJxnIGT48wRRjmvG/StLFg4KSpS4i0QuvE8wMH29oFYC47JJaSWz+
tQ5W3GujG/JMVAeXz3mLfN6a5A6ktpMNqeWXdXVKdCoifr/JuA9WBqbzRI6DRqpD
atUYVNPl4Yro9Hgab8oj+mHNAPOgwFGK5DRb9SZ2KzfxbYv979UzCCxVwD9dV5bo
TjEso31QYUb0w8kXGKwVf4cezL8gGOhw9hk+SRADx2vxnwTzFe+4oa27b5fFH9DA
ws3SgQKdmXhVaOWuO5EogRpvQqDFo2PzuLKckPb8MTeqpo7tE8y/ZUW7Hb8g6SDL
1s8K+U6USwcr7IVOupODaQZRwkXdJftyrzRlwbpfXczqCqQ2GOOLU95dFS0GzOmG
HmUAzzx1o4yhtZAH1YZREn8wuX7Jz1bh/rRWtg6vWIfurUUM8Skw7AQ7fh+ojSq3
Jr0nLIIr434h8kVp4czLoGR3SYL29+R046WzeXCVyz/pe1197SK78SBp5792eQvu
sYh6da+nl0LfadbzydKMT14ohXqZg0gfr/knbo0kBjcrLTkqqMmOzAJ9NzscxbvP
LFSkXRPe89yq1L7nZA6uld8sq57ibzr7KTPl9qJuTG0ssfEa8oBqYNgIG5xhdsFC
A7lpffsOq22ezCBvlayLHfJR0jA+45W1NxmfvAPSaHzalJfgZZ5XFBkxDgxiADAW
xmRrI2BxxY2JZyFpRaUjz4F+vaLx1pQG+w69D38BMwyVgQ6zFPWmwmY/rd4BDCx3
+uGJY0O2MDAgtHOd7THvKWBDN2kVdnXAMKQ6BdD+yUodD3QofdckMSNWiIHjoaxP
VbpVvay1Suzr7ywVVE+9/2Y+5ldStdPzhsYy4kWnntEQShoi7CQmW3hW1qQgTRkh
H4P8cl7WQXYyQdFbcHxNn2TtbHiYxM76VuqIMfECq7p3h7t/MqCoFNFOjTtetO3z
TZAnhxCie04ELk8kfuAk+Nnbr/YdXi0pbBVae5YU5DnAMZIH5nTqmRLya+L5uwx/
ATSN0SfUsof2fQ+PTEdkjpQjYQHKun4HaEbiZajT25KUSJTgEIy52ubPusvO5+4V
cdmHbfEnjufOsa5P3LwpRy062OJxLfwRBSoEyoArCioCQg1JY1Ix2ck293z1rQSc
YjMjI2AMSa4tZpD8Hki6dRGq0VNmNU9v1ufIhKbHA8GAJmJnRbOxUB9FoUwu9qoz
ajT0rpZ0Y28jt9aPR/joSyjZy8Opoq5CE/OFWaq8xHyJWXolzC7EhbseEGYO3Gx6
vI5Rxi3Y253U0mqTxq02ZNkjGhFAwLB3R6QlZhMdygs8mrfbLj9fBnaHPhpqpShq
zekz3NNhQHPhZO6MblaBSQy/eCS1ykMy21VPEWCSihQxs+gDcIpQk4A9392TFSWx
2bVffcwa43PoN5Z63DL/bjmqZgXjsfKiA/9OCw5PK78usMy/EQakRqvuW7hhYwja
SdCA9OprRDOMDhRmHPxLPPmJPijJ4FFgX2qJAmjS3YAVw9PAAe2TvLzNFapywE4Y
Jh/wDd0HnXJIcXOGT5P5t6XDwSj8XXsx8NrRI+cYmKreuPJDbT3bfO2C8HNHre+I
I7dZxEyafMbwoZjvOmsSGpCIr1Z2lu1fvw345CkroLwGKqgzTWxIP3m7oP1UMCJA
OnAiYyjqdn3mnubkkwFCIqLXREM22lwsJyZas21hOD4ikmEierLAJeUDe3o2RQa/
KUGmhyMXia/jsj1G0VUcXnr42WU1FlzVly8+QxrIbZvRA0gOsJJ2aC8Ugbqpm5Nz
OdR4+zh406DVeXclzYA1O53LTed37lOYEhYurMiaXxV0vrvlcveXsdHcBMw5KBlR
u9JJcj3N1rMsoGICbr8x8R6Vasjg3yar9tN2/eult2RW8ySGzZ8KmHeUITt6UqQU
/AGneCTObfJcX4NlOJHsSN1UjycYu581Ob61k0ktUpZ6fSysBrL8ESJDpiDTOIDe
ZJ4hbmtzaNTPDBZiRu6ftjJ55XTCuySFvUQbUa23Z9N8BdCTqlsR4XjyL+Okym/H
eoUCjBK0rFP+qSHod1JlcIo0RTPTWEFXvTrvFe8seJhppqlVoWXfVf11GttRhaRH
HCMXeXnv/Ni0oA2yB8roM/BPKzMvIM81tunulhCGtLJOV/X3pGH2U57b95PjgnNh
et4fRN3Fr06M8eNiyHdpgivi4AzIMaw3sNOr0Hq1XQJ0gFQClGWXHEmL1HbGc/lO
cMFcYersCehx0RSqIpKy3Bpj1s7/HqllXX/u1vyi85/5Lw/7N3CxkIIpH7WotALt
rO7KHGbreH4Pi5ElnrUm73hnVDaQ0FWLIR/2twwnGLjFBf3/FAUMzcixxNMKqFPU
aCt3gqf0dv3Tf0GKteMRl0kPkAEG0nXZWRtxqpcKukiR/+4HutyuQWrBjjVKRcPF
gcsP+iUvmH4wZp0Yof8pbHXIHubdkzoMZxJpAmCWHrXxAWzpi/4WGccYgcurMjTT
mmLEXODxzbr1EQ4JRtDfyFjSkFgERMNLWEIRJ/G/3kvSx1ZOUdxxkBG0HWcoCIlX
Zrq/TtfmjC27T4Qu79/YCq40pjmGpNZYAy42EScNWkWUh4GXWakun/2t2EAqac8t
N9aFmGsYdxVRb0R/m1LyQy/dMTHrE2haE/29ukp/jYqt0/VXRpCv8X6oWi0YvYUh
ItU2OfOGEfH8DPQz0uhulgUezV+oayw+TFI6T/jHzh/kVg9AylajdwIb2CIX6Xxi
+GD5VTxF9dvc8ksbo6IflLWrshZtVpVB7AGRTlLrR3GowNdyjJrtrZYCeJo+TKE8
cEYiX/D2BHu2wNd+fLSqCv/AKY0zbp/ssBvVbYyzoKqn9z2LbtNWKAXvg6JRW51a
ih3hdtZ+Egj5AFKspLaqMJbPPElnNZjrUM1LF/T4LkJ8QvXvJ/HHFB/L89jiq36f
s2w5laLoXjvtPaquLzKD+85isKXKfl3J3FxD91HF7gYkP53SKa9gN61uFAIY0BWt
DsoQchZLKwLN/AqRuu8O/srvE5OGe4G63Iqu/nyHsaRVZpgpDtehrYJS9z/Pz3Xz
pzGaU6RRpACVRo/yIqA2RucR+P17a+DosaxEgXdlAuhoAoWiRRYxdmIt5LhvHXa3
SnFl702sAFEYYy+WV3qRsN78jbd27rL102yPceCQxCMTkHdrqOTcDpG+yZXNGwv1
a4ekTc210mHVsbFrAL2cmI/MUTToTGUrx4gcp18Nru6FZmD+7m/t6qhRrn6pxnps
d5mWkV+u765MDH1Xh8ulLNhlYz7FhMxXWN7a0CCPHZA828CM5biR5cQAG05A3Apn
EZSwYcAbvPQuSEEx/4UkYOgrtAHsz3nDO0XEh1KRYhMB6WJVgR8U+2ollmqhYekh
TKsw5ZFZnFqL1T7Ss+eNCuJFV4adcw+On/SjuTsEPL02p9DXAnMUJweN7WR8ul5G
r3V63XBM/XO1ZM2EEBDJ4ZenZmJahlxq9G88bq/vcVoeqn3PAXdYC/Wn6/ji9UoR
SQVcVW7qsWWaOxoDbSrZo+hmjVgD/kGpc6tF5kJlaOrtbGd/G511JfCiXP2EWoZD
0/nH9TTyhPi13Yn6nn87uWSpdfeh5O5OseJtYYp/xwAR+fJ2GcAC2/I7J5wA9O43
VG8rkuaJhAIsgLAqoS20elt/0Vh5yk1+pMZ72qdHV8smgRdpbCnP2KSU5726CEN2
Cg+9DO+dTJ/0pMXwM97nM+G4HcMTP02zqyX0AeQqnaLdV+1lzv6hYM/WxbIBkI8Q
qtrS6EARr1C+L+I+OmFhly7BfzHFy47ilLQ8e7ps9F390IL8yn8cOB7FMeBjjVtY
4iTxa5jrVuKU3Y4QgiUrAXDFMqvK5WkjGvuh57RzTlMxLrJcRDuxw0AGm+2EgS2V
EPLX297pBGEIE4iqyYU25xe15mIVvCCL3Pd9DeZmZuIZhpOo84Wx8WhPGO+i8NUd
q5TIc3Du3GOL/ZFIoyEIjS4ZTwJZcl3OHC88BL56f9cOf/vLpqODyJHpewvc3YOG
7etgwzcPQirIRWU9O8X2wx4oNIJgg8vm2AwH9va1x0ka7eZG4blOXmyWToy9WeMj
Z+mAFntg7XRp5omSNjHkVR7Wbfm24ItJbh79PeFffhXluGaDQAlmXR5Jl3fAusuH
zUcEXe9fDAxkzTDxWvYxhn9CBZXsGRW8dN7/ZGpMMo/yejxQ9LilTwN22o8QPg9o
rZYNAn0CpKNXzEPnNBG67LM8z/FhrsLho/UlHQz6q6T2YKRqZD6DeThdmdeQOoVu
48rrJTUjsy1BnGNjrb5poNJWEryQtTqExMwB9jKYCqm2FVvX3JMP1F6o2inLiI59
MNRbkPOnV1et1iWKbau2yV8vovhuUp135h4P/pcG5PeUEg+rd4EpCERXTkoTNYty
O5JzDYOSsFZ+IVVYlF5WfAGbU7LqJL9O/wyRH6yr0XW1a5GB5dFQ4p3ELKtJryy+
Wmd7RXJpPonJ61t6dgcTIKxYuz7IILrJsNBLP/rMqfUBb3hP9mhmvzBL8dczNKvs
l0SAXUPlWd5/HUAhoTPZF/KI60UM5pItRfqyvKdr2X9nwqz12qt1c5eg5ZExBEIf
EJI8oLLKuRaDkAn4HPymNYVv5MORyMEDVRXT/xzq01J6ixAPIrhBaSTkqkNMt+re
VjE+OlWn3CJg3My1BP4vyza7RrZsvi67lWJfVWBZqB/6DiPGhOUlDehv4gMQyqUd
fzTbX2z/aiqnZRBq7OoQI54qDdzhof9gAIN+saAKRG80fpDVNiW0e1fJQkpXQi3Q
/2cAbab3ta0cyENAshumtRJ6BkVHXMI/3HP2DmPHmBzgVYU5a68dEMhat/qiI2UA
g8MoZ99Xxy4MH914YVFJSdfT9ROIyJ/ak0u+t+E4P2P4TLlB1bqAhcerBnnZbx61
UaPlFahlu7g6+xpgz9gVdt8nMhdvN7ay6eelsoBQKVtOUTqtfYtYtT0eDlohZ3OK
LUrfg9P87cWWqehsLZOq/vkB+qyqdTGg/Knvxm2Xtrh6KBJPYp3sifQ7GGR/OitN
VgaqeZ+WZmxMHcc6LBWMj0/fKYIS6ALi8hg4RiGwXV/dc5hvnovIW4A1iEnxjoUv
kKCclos8Nv6msEgQEL57/RkkIC5tH/ECckvTHkfB0JVvSJwbeQTw8ZC01sQacXo0
/c2u8I2TKIwZlADwMeWNCNooPRtCy/H9JuRA5xFzfWSs0R+WvMYav7AWckMvqNj4
0Wrxeyc98k5yJBTntPlnQ/BWGXxe3Bmimn4/KuAVHQeajQux/QgSg8XJsOF7MNtG
RGOIguaQEmIYHfvIXnkGxVyDR4xxLurkFXNnqK/4WitZJ590vhoZ+shI6XO9onR2
63mpprXSMNV4aQ8s/2yMgN/lUv0Kwx7TjHUDWxVjhbcuPoHWte9/Fvd80bLFouTs
Kbk/YAtSQKvYQy3TCNLg0ZLY1wrhzOGn1Oqu9aVBOk7i7CLy12yL3pAJirqnZyTK
+aMdbDG13fP6MiVEf39TlAye4ZaFXfxH7BWlTEBVk3qUFBX8wkGMhMp9ndtVzs2z
9YK5178VxIvWL/zcWaTwJhqAjzSxTeDbi9VBwyOmIG8uwPTw6ZIRTwdmqGXfiRIP
NRikU5cV+nLHdQ4G77S5+XyXvPeHLRdOx4DqmQvjtdAMlWTGogXZXOJCx1YJLrXS
2Sl6KBKUOlt3A58h8wZTcsxNnuOK8w0+4YJvnix0udOoQ9I7bUhYwPVE22R+ofdI
UAVbDWLg5Oefi2MlGqa7n+IWXQLkF+bQjdWFbJ9ezjA4H444T1oY5114BYeOq2Om
aHkU/IM7zeybyxNc2hxOlzesMbHTbZCu6bWyA8C4KYZmkaVx413hm5owcBlk3Q6m
+82V7AJ6+N7JzmYTGW95UpbI2zUsZ/xmOcWDySOIu6HJZtkR8eMcxRvrbmcUJMck
zfFKEGfUalN4GP6VKeqLD6H0l9+ZDBkMzpuoOkfSlIXMICoY3v9v3oNV4XksYiKL
vUcqnLSL29HNjG6QhLivNIV+8qB8GuoKfKDnjB2F6ijnLZ+r0yoZHybkPoUCxnx6
zGk47AUjE2ebHLrPabJNh1EnWrEWkgox5u0amew2Vv37xLacHIS9HzWQP9IfIRt8
wP9k+4gAwQi/lvkiVeklKKCKV5suQRd32RjxGAQNUKrAhGsni8LkvYOzcYyR86wO
oqKFnIWAO9WQqmeez4w0GD50ZWMD9HW5G/2PD100wc+Cm6z8loCWZRCj5Udthu9I
UndPQnHaRG4Oed2GAm5oIQT0pOuZfVyuDE8LjLcg7eNiHu37zfyoNJ6v6NXzDEbA
KKPR/Z4t2tOR2cxe/GH6RF18cwcr/YwaZFF7I5549mfDpqhayx/SikA2WE0Ft3yu
zza7lmPQnc7H37wFHUbtefTfZSiwCBRdPgh1l/Mk5Qz7FTwUeVWAru/PsNQxd3N2
tpBjrqlduxXXdX3rqDkhssRgt+s1G4WdvMa1ANSaDkaRma4VBEaBznfxXmls3T2r
eyBWxFUA6hX2FY3Va7LsYTA5kaTCl8qJgGWp62HgcoVJr9oT1cXiHyY2M1155hfI
xF+rAg/lzoKPEu5H0HZd7BjTkK43BJtvP6Pv3sSmc5H9FIdQ4YcYnC+QREvOc6be
Wl2cRAUrYgkxCPY2/3ZyJbP21lwSf0xmZuxj4MaaDSJTm+3Gq66EwCRfvg7sfQl2
nCtMD9o193k5/zgfRR7iMFfzW/9A0J416Z4rS/CtG7m5QhslnNioFzPBeNQ9x6Lu
pbxC5ezEYLS6k4yNaFInxiHsnLEpsuitx0n7mrhLLyaUSiZ9KZH6hRD3GgMsFrP4
C9ZEu0uDlZPPdrUtQpX+PtuqWtMQgz0Z6vOnJKWXhokhZjdPXVk6l1FCQUQc7Am0
rqUrILWs3vItUQjcbaYA1JonUp4THKntovVfFa2gD9gMHS0pN6vRgevHpbZCYLlF
WCjmbvRbJCJoz36ruieQc8ZAvgELaYj8e+elmNvOO8JaUYNvQhz+Q4wWuBmCoPBR
OZ+LJUH2NlMY7auuRIJCkX6NWBjMF9GidSjgWZ8rNO7nDxgUrsBLkadjkNRs2kE9
+9bxqvqA6++VINrfIsRvPePo+de4nCQ5iOnHMXraJa9sHGwPKzpZlXlG2pk6lr/W
/XQfxX/sjZ4Tx9m3IvrPYMevL2NpKbrAw/lIIOzE2y2MAx4BC3lfyzcMgeJxCWDp
Id/+hnflNe88DZ3NddOcuZM3re9WN5n5W+2Weu/HxGBbQyKXdi4XuMqBdf1KjygY
m+zKAcxGTQ65S9dnbmPTP/GRM4TUHCoaJzsyVKnpItAcaH7n9Ni8J1oTsiQ/LUl4
o0T8A3YSrUz2D4/XdlcJTM9UF7Sd7PON3aD+ibHpC2l9qpQaZTnyqJXcYob9fhOI
bWxxZtWelEwIYWgaK1xFLaaN0i683KV6EBGBI283v7I9SCSFrjnICFsqXxrUY+97
5RCgpCseDXcwdG7cQxceYInWZMjzyMDKZIFaQE2AwxCsjdePusBTrgW/S/HVOYzI
xkPv/z+BXm5MEwNtD0jcLKfRcepiyuw7Qb0lystBlZg4X7pSFrG/gXScIXZw0GI0
WAyEcBkk3nz/2Ai/9X278hNf2JuQ9Wx01uqbiYpWCu27K6CA3vpUFRRMzEUJypk5
vaSzvMWTPOofZgzSkMagfgLDh38QvUiLYe5qzsVNIOX+TA+RShOI3mGCQc7TIA5D
u025keM5qpX+WP3kI7NpePWc83fpBR5VPSyn7oyIfqTWkW4UVWxMV5qBpSk5SE76
R3zjPwS0+8EZmGVcozfzlsGoLOWF3li8oayoAtGZTWoihAE8EakbJWcHijE3HgFi
XzSnCGFdV4fZc/mq6mwN+/ZFPFwZzwfLPluUvTsXjHknb8EA2jCazogJbPJ1xtKY
U2vBwXlzXPvyrRbt8XyMcb4zL3+hn6S4bXXlq71OcMJt3tOusnTxCGnFfUClzUsb
3EQvsrACD/jiipT8dJaBkYWIa87ktBOpbH52OU8kmLBD6b2ZN9VivlndMd+mqNs+
MRjX9Ryvws2knNoY7Rd+cj7Tx7LG6g4Mck1BYf6ALOS4VOiZDJe0YLrWRlUCgF7w
9lF+Z2izhRLcvp2NSjKFklEvySAxkRM4vhLawqRuc15NF/zqzRAwue5tepaZ71sO
X80NdRliDqIsJBtGShwnswFs3mufKwuYnc4ZSNOWSR2iso7yTsKu5KPsXMMCpaFS
U1zwyB7jsacvKbfkKoFnGpN3YqRyKtmEiJOKlxwYkRMZNeBsEHwd+ybIbbM9iJL0
6zegOsQyMbEF/GhgFFu0wmeZWSqOWjHoKkqU7s6to94H7nIq5ibzyxbYThMnGlSl
8DlZ5g24iAhts+PEzg0LhAukLgVSkDN3uDTULqFk3nQuPEdP4Q0faeNWCnvHlcZs
UQro796F+pk5FWZaGvyCUIrbBVLnCrh13LcbJqBoPGlW/hpn8Inn1fkExtgghfJs
/eyt3QqGre6zoENzdtDrYL9adZtUu0rjcuoS2FUAlyxbMw83SsUY9S5JmBA/Jyhx
uaxaJQtnEJASUN1JMfQa0yj/IDMFS773HymL7NQV4QbwxwS6ut0kvr7wBwpseCID
3rgAVc3TuU2WNUjYx50sacCwZwRkZ67zFOnoAjUejUGSfbztKKNQ3whn8W3AcO7g
JbkoS5dUr6wdwy1vDMXkwc9jVA73LdQSwmZNOaDIzcevW9hxxu+/4SsVagQOrmDz
jYS2tjvEYMbu+pCAOgqe8eXtxt19pQZcKyzHxGfxSMeueJnBEx1EqK6j1/R8LYs3
yO46bk4piNv0T9rBefDtXUaFSxRgQ82vlPTUKEPL+xylSJrOr+/3jCgXF65nGTBq
miB1I2fDnp8ARTHVn8xR+PgtiE+laSqzjRzCePOdjTdcwivj6p2FxRalFwaYaLkQ
0aYkhg7xX+I6C4GhmjOr/B7yJXGb/qdwoZfUctj2+vD3AHvjuRj483hLjCE5F78/
LfdMRnc27IVSlZeZ0ehz2fes/8UomWl31Lex6qNusHSZt6WrbrjCMgWk+P8ZR1e+
2cRFVnEtcHZJrm34RotEoH8+Zti2jw68cZOxYTKQ4ibg/yU99q9M0YNO+ZtDNfdG
N7KIhtvKlnfSUod8sDEUdWfDxve1IGu+/ZPpCqhotuccb348hrRi7tYqQAHgqnda
o2skxfVS1zsvePsZqXavZJlhctR4p/xZnG/spQoJ7AMLDMsExsnTcHWboBMQBFoQ
m2Q3YwfphGgfmZlQZgRl6AYuECPWPJHxXewbmB2adweo7fz9SOd0/1ZW/BQjewhi
FbzIEX8khtHTpf5zeP0OlWuk5+nQKuX9Vm1Xm0R55Kv483ptBrI20UaXPRuRwERo
HxwaNJAXVMEDvOIDFSfSzuO50KdNjoagn48ZDcay49CT2QGQge5JAOknfFTcq+Ty
WotU8LPK1n75mrv6YjQbwD7OdvL28tbC0RCTGYYK7IgR6gn5d/C5MnS49qh8bjPA
Cp045ao+yrD9Ua4hUGRICE1lQfExkapTVHqzKLbTEmjlIC8YI6iivZoCNb8ha5NL
tRdSYQ9BGpQ71HquRKGpySYVZ1GlhNnxPIDD9Bg4ssOIJ+0uh3iEGfJPSiTixpkk
J57bKDXrlkU3VmlW1L5x/cKxYdqRiu7BlRaxljl+Z+RvEM3mYzE6sGc7D56eXCTR
DP1go2KcIp4yQ6q0hCFd7WfAijXVHs/2xScGlOTeMrwyyUAHceibagGY3kjm5Oyl
bXav741KEX8koBlZ8btqci1QC58lHHKInzNA0pTFeG7Jv8tFwmiykmx4LdYSbJkb
k8BVvVND57QDYRpFgSwSaLA66CrkyMS47tzu7LM9nDIzx0/FAUtgtBdHwQQ3Ym7F
QE/rR5emLzZl8/w+QAFvlv3CZSR0NAxXlvCs9jO2y0eObWjL5UkkVkvav1Q5pM5u
pPF2w7eL954lHfqanMHZn2kBH8lMMILlN3zhuT6deV4Ad+cvaXFzmehdXN8hC7Ld
II0EvwDv/Wha3kq7jXy6A+nUJnxLWgi1doThXqkji5yYWVKk7aRgz6amQvrrrLtf
tJrjc/up7yG7kED9PGwYMh7x7YK2zJdcLnN7c4BR2CW4hHxtDUfjCgcl2A6qZ1VK
sDHDC28efVwfN98SPLDvnPc7kCu2WusIEJDtHu7y/bNzTJzRozgRGjRTArcH285f
yRgHFD4BwFtaw8xq6VmpRmT4r/6vX/rpvT/5gar8FLnyDvjP9c5uJr3pFx9dCBpN
pkmuzWA3+1ohmVtbnfrODZ0CzROznV7nxnExdZ5vCI3LU+eaJ0/LaD64+3xzXmTd
8/KhbFKLDMYR/GhvDF01e5Tvo8hM543KdMNdlFGh0MKP7+mK6m1rkrdSMO5Fb9av
I9hiaPA6Zs0zZMdwsLX4pBFN0DRh/n33M1KLk864Q7BkFrLNQNqqbnKiYtqWvK3P
NV9nb6WHDTnIZLfB0aUn32YtNsFOS/yU9PJyZO7ej07XeV8ROiiSLoitW0eghn9K
UjN03ocQpuKHRV46YjNxxiEEDyfBhHbIojGMbhja+2f5ZIi8CEMD9hKbbRftxt2G
hxoQiMIon9a8fHl8y9gwyHlQ//2shcerncnUq5n4MaKCMkuyTrgV2WXqJ65lfHHj
ytUIjl9YztVW2417VTmLcAMs3bMtaQ1lO/FN2/+Im+DuIgD72nKytoOfdlg7FfTJ
JIHv45ZpgkAy+cRe4o8/eo/OLos3Mhcc6B7e9qF9EjVuYFUO9zywD2a0g5lBkXcr
/d9yBkHIuQnNJm+h4Aw2FBuvRYFtJFfIyipZIkkLn6g1+rHYmPdHHjJ9kT1bWLhY
PmLhzmDiY3lkYOx/TM89zBXCK3kQ3YsuY4xsPeT/thHB/Si7x2djo87Ed1ybvwOU
OvHlzQ8aAL9KRpLJwmWGyYixCNc4UJBb2ZRtlpuzplPq0v50WNtjK1abPWO/cAAa
6i448pZ9QgUXyBNz7xdW2nFgcAZtrZyvdO8sarJAZWnt51b8jnwvMeL4rB+SQFfq
Rukefu4t/UfLExqfioSQpd9s1qxA2O5jio/hggkec9pIoIRmUEja8kYJz5TWC0tH
9Bsb/fO88kvvhJ0Mivher7njj+0aH0rBA+sMMRnzmCLK4PUgENQzIKC/SHUXygL6
tgn7la49kcb3MjkmM57rhbB/kO5wJzw0qT52LjGkjZ2qEkFZkgIjqcxPRJjbUQ1X
T9GoAeNa/MIYj39/bYW6IPh6OWPejq0X4zRbsHHqU1DjNERpBj+5GXzJg3wIW+mG
c+L8TiUp6DqAJtfAlPy2DidlrmfDRnFyVy+9L1Kq4oRSd1N2BdGhEylZjvcs5oBA
Il5Np4VOxGR8rOAxV6j02MTfqmjWB86Fk/lysoTwKNLDxVNGmF8uo/G1t5+famDS
J0l5vBY8ipa4GM7XqiBZQRrRCDufHEjQgm6kxcZxYTr2MSpS/lHXVE64fOgVhiVa
GWNpD4S7F6nP2uIsxSqNXwY9AxOzdltEzKLT88qUGNiPtENnCCRapHpU6aXx13PX
w7P5H7tv81l1sBp6mZ6Y3Nr+ryXi0xv5o0GLzYL23L147pECtRnlFaefkO2wREVb
r4zwgzlF0+AAZyZDMfzSrN0v+SoLwxeUmbeZgTyHhZPiUeWn2vsLTlPEMcAv9Rd2
j/HQ9KC8dyn5X37p1mUb60d1bWWQacKEy6kzgheRc1y5IOSn56nVDMT1RwOwmTfe
+oRlXuW4soASdASw1dbVTWL7IyF1OX76a16iS7Vy9yhhvqGEFChQsFWllfDbs4Tg
/hptWDftC4C0/4Yceo5Z+tIN757Gx6D7aWcYlbnRof9UiEV0pSBWkCUv59S7Hesb
qL6uWwVoicF2X/kknIiphbQkk0EM1DMaSzrSDHzZ8v6Bz98d3OK7vGGsEdh7th5f
x3OAbUjiVgLiW1LiNBZi5VY9mCXaEgGKLn3gXtdPwWBtzePHHuno07PbLI8wDV56
w354oLqkecFFXYoO2Suc0OwbkUe2aWQuZOClSBLU5y4lHjYR2XW4kgSMmo+KUKvw
QQUM3fQIu6AeBU6QlqEg/hUhU7AQZgSzp96nXNd7OgpTP9xHzhX1RP2oFm1CMto9
Ahm9Va2zMn9RPHRyCFKSF5In57dmMQDkK0nT63r1mPOvq6Y+rwY++XlgtiMZ5hc5
GhgsGRLw/helm4rvyIoCnXGki8/0IQ78+kaeY3kQ7AHeImmGfzhn/2erCVYwQfjP
ydfbQ44C5L8tXeU5TBrz6JTN+gPIxmlshc2MPjSTuU0nCS2c3deFWaz5J7eeKPG4
GElw0nDJdDdzEySPBqATT2OvLrAuNWPssmAS8XOWwLEe/Y6mNyw3gUKE9GQNK8wM
leLiNxpv8BDvoVtlbt/fFrEePq0/bgmVgBWd4NR04ur8Z3BNwT+iOiD72a7PoaNl
8FUd2Eah1lLlVgSpb92mjT7n5uRANEN/RNffQ5S1HOGbKkDhoC5q6MOpg4sr2rzC
PGpfj9htwpvDO+tnk+lLXpPzvgTORL03ftY7Y50QcqoXOYytOUFMCI0M3/oOa90Q
no5tfBhYVq5Bf5v943zfRjnwvOZB4e4jw9LDMUFAZvuB4NjfVpFCtHBylNYe2ENf
vId6k2EsES11OZAmTvppC47EsfgVhsqW7BVvAvkOZo3p4qIUTgXOtwZuW6qG07yJ
UPcdKn1G8zr9vaTbmOAaKnekZ+LheYd0RytoPPgISB2IYMfUEnCAiFONDwdayQci
xCUm5+7caJ/DfUwCwoKP+jpiyOl10Sxf98f5+cYIF3a0xMsp2nlDOWF9Cpx570/P
4x6yFdRv5oRBS/GQVP4EfbDaNvA97GXhtHS9GjDJqo6FpmbhsuPmHABsKXLnaRRs
h/70kv2KWAzf1a4+vGOZUIpWFpGLY1Tbj5Jug0+OOrFftQoCBqo3inJAOFP1XQR5
sS0tECXpIZGb4iLeWk0CgYhKSFzlSlS6LOPG/wcgoIiEa0S5UN8g2bK66BgnFjYK
8PEtt/PMuTVImvXj5CRTitjSr+0BPM6ADyrWcshTu/BBCY5uBB7KX3/LPSxnJsPc
ACmm0SWCZt4SnqW5z0kxel3p34huEcI3VlGJzLi8YTk3yzgBqW7ZVRJVGvZWXLoQ
4wT/LLTJ/6nrzdtfb/1XPmrZ+y9q+1Q4GLhAPLHD57+MTvqZeIex9tq8uc/n0T6k
41+5Z4fsEO8gKJxk28qO3C8VRb+Fo0pzRDJuULee3QsAxCIGPrKX74zf9dS9sTlU
rhjjQDobVLLPI3H2vQ0cc3ZlcEm+qa3wXu9kjdkyeYvSLHsC9DD/zql7PUEq6EYH
aAm+5D5v4VrhBckYUWi74yoNsVnz+h53/w/HSNVjyrfbhiz2y/UBDi9xZXYnbx0E
k3x0jj/2iEzvoppfx7/HV2s0GW/KuSZTs7152GOTP8DbldBPgSBKfw3UX14Afwn/
n+AW/mRLHLtD6YvJeutslwTkumXYyxtlHXS06YfJ6EHEtoJeFKkj3fumWTeOT3B3
0clzSORuBhq54RAsvg+evx31vo29lGXf56kKiMR9yFi9DJoxMwBUJm648R3+M4AF
SDjopxDljVQlEq7OUSJ/02KUKPFHCPC3vRkVtPzS2e6ixqRSmKjxL2hF1t4nZdys
HZLC68JakBpCrQhYI80cvJ9r1knHljt9O86g62z6c9RE+Dm6kzQjKtc/cxccDUQB
/T/iqghWJ7JRCoOxscxhvtZNzGJB3VLElLAZNSz+T52vroP6MmE+UnTWmbPDN3Rl
mGRjhT1ruPOJdvNgAsGaBXxYrkCMoqrTb92Kp/ERS2FB9CQeBL522CVtPH+JyJU1
U3j4CWGa8D2gNWJWHszrGssl7eIc0YKdKnnvMCurzjDQ1EFOG1kynZCg4859uz1P
Yeho0r7iFZn2Ue3+VroOKYamTiBz0UcUnhTfKmDcLQkOfCZYnzkq6KyalxeyNMvz
Vn+nRmQiupfHUurUj1Mv4SUn32QXWPRJTlWwD/1hOMz+I3dHMt9nux3PV4Hh9U7t
RBv5YP4BMCzI51FNKuvPrJtRgc68IjwKVb861D4+JlnSO55Lz4sa2chN7y5s+qI7
mHrN4cbVZ8BRT3IzhPSobg1F5HxBqB9KHP17XtUZT1uf6tj+4S+yeoTxo4H4O7wS
QVNyuioC1HHHoeDM2sG1ztdqdhdI0ten8Pf/LTDPVvcgIBAcaJ8ARC/5L/YMlKgT
tpcp8hwX6MRSqVooR+LUKnQpfEF3QOM+nxnkTiJsawAUrxw+i2ReXxH3/IZfs2mw
y8GC+EO2HD/7vfbm7/B+bOk9O6ZlpfuOPa0wbgb6fS8k6M2pW691j4GqCl+A1w+w
Tzo5EVkt4GJyWt6cXM8SYWIaVpBI9coqhwsRviApWvaXOAkNO3lLnO3yvWArIibR
fl6PpRklPCF6Jn4dRRjCPARXfNH6YfcN98iERD7SmMWeZn3AAfkwyS0DF+Esg6ra
ELnijoCn/MGmBL+R0bNQsGcve3mAZIpRbUPHOgqxLdWFRVmD0Rn6j57+zaSaCSla
l6ldmVTf63QtWU4HtTkhPsRKIr88tcE3elCZb77+E8GS5yqQ7L7Cja7RZO+kMtt6
rx9UtRmEYmiAm+cukKT3o1t6gpZPv9reth/Im8nWmzOtYRg+/0lG0BRhPgckNGD+
z24X8hFOtLsa8XXwf5dmPpZHSFXys2fMwrPDRnCw6pv53+jLla9SQ7R2MlWXwVUF
8tuAUc7f/Nt4Vgu6mK8yMMHmXL5PJrtkQqDwnCWh82akC8UxDxIqAsi281fjNuDj
6DLPMLRMkjbLNeOoWNAp+oSEtebUUK6bLDztcM2t22gSJKay0Bv9JjYTH66HSXHy
AHjGMY7IAWITny1jQ3dGy4drvAKLOg7mK5NAfCA1VTdjt6SPyiMhphF4E0zmFSbm
yh22LM8QyrZtwFTBAM+pQ+hl9BHJ/36x5gbVTi2DFCAc2HaFpnTcXdq0CFmY9GWU
mf4NJA6IexpvLUmsyuKSLiU/1OGJwBfRUooPThhFCL7DwranfRaBkOQchTQJNkdb
PL4fo/krJPheUGhwxIJqu0f1lhH4q2czmCIAhS23sjJPpb9g/h4qGEZrQYCmaTyD
E4Qs3W34WzF5qXJkQtBms4baqhMbJehNw+lDOP+U1h+VUN/8vi//w1d6SW9d9LA4
++z9vM2oxm1JnRl9Oej8lZn4WexbXy+tNPVNvYCep0Qiurok9oOBtcikVqnxHIyF
cKSFuPuoGu4wtVfUSGE+/+1hXyN8tOfGASAxPHc8PL73awTbWCN0zoxzdptHhgnQ
PymXhC5kL6p6ttoRMyNyza7wERmvnvj66sdJiDlc79HG+vaVl7rMBaxOIpeN9uPD
kj/3bpe5i8mrjQa7gSno1GgKrFWbZO5mxZf0+AtNY7nSX5+k8fO/P7dvyIHfCZHr
JOFUUapYw3k+zl2GcB39rKXJLdnVouH5IUske2wZAyhFXNN89ESlqxKgalUIRI5q
ec2gqRNkr0QqO9AI1uS5RVbdQqmX6twC9wxGdOWq/aLFxJ3y3jTaPhNVgPu/4afz
po2pEgXcprHF0lNb4M8bpkGP1hwRiDoImrHu+EHug+ruDo+BhfkOdKvGpah+GplK
4V5YAXjR4Jny13xr9ghhUJeRKrjC9jLGhQeicJG/9RX7DcMgoAz/WzV4vmJHx1AS
KO3QVBke847B9X54bdoqzE0phTGdJ1LXpPggu/TJXFH/Imm3PXqeqmwfD3eFfeaH
3lpc2G61mFbhX/6C1zFK+o1QGsC66zS4drOi04NFl/yA7EX+hYHV0Z7BdlWW9nPi
YenGkL6cI2Xjy05/THGfuT1I8Ve+Ohpir6DYE2o/CR4kv3o64/bhHanSzGjEJ5MZ
ETgzAE4T2oJupQsPUiGJoWRLpQWRIcTQ/Gu0/azajn/jeeG2XgxJHs01dS6bIfof
YMSiG8lRwI1dCrslOb2Ey38jdFmo5ceX9lUJUBi2oNNZgbcq6JPfV8c4M/1x7BXC
e7IaJZGSWNP48w4Tk3nwX+NUejz2SUZ2tq4DQD9EPXzXwoWsb+GzY7Rue/t2VC90
A4zpxqMCYRUlXdVfQJcpNGVvf9ehsEUur3Wk5a+NR9kEgGe5VGTeKZu9rGQbte5P
3SlHw85AVDQXXwbraPZWcUZydE6BwJud93CPrTLbs4A/EaOERf12SU8mX3PBVh1l
GcWZQrNFDOwwtmB9LtTJzcN9edwnZz+q5dM2XaBBCWJi5xaLVz40w9xOkMqePr6w
ySZvwZYw5Oe3S9eUZikIkF6wLXi5yPwLTJ9rX32e3F+1e6vgsZGXdJdlCtD5d4f3
UnltQan+Cu8FHrc3mmazrYLEa55cVP+new9F4FFpxbp7ulY1aITEBnqMXUAy64qu
zYT9l8Lfe/wZn/dQKo0HepBZJRvd8yMTWZ/ANGhEnTDsGeJr7FKp0+rpiiYU2BaI
2D7ZHnPyrL12lMxFTu7008dE+VyqmgsAqCI+ffTB+NmZeLcU3rBQr9P4XYXKEbtS
Uj5wbB1h5fSvNA1Ai4A/4u7p+fYaGsKlYJbZ+acNhs/3kt5waNxYykHLw6TXnT3f
DTInOHIk9UXFVxY7h7uHzoIRbInib0uItZiuBMJAYmpHvHUYkxukausiBzWlY5Wj
CP3ezXi2aRy2KRB3waPWyYLnAV+6TBKpuxWLyhQ20xv/4JZEwQVz9889isqzaiRD
ZKhTekl/wm2r2cQGvnNtvLPbHWztENToSXEezYT3/kERB+74r7vkoRDcea8skJ5C
PmwVdY3L/SBNahd+uzX2MtOCvCRPnf5ydlINJtsTBuQIamhnXGWgLIM4BQKmvokN
gOvmWi8cz/s+NeVPu8hQo52u3efuUi3D0ZFnR+rB6owKNCI0Bzo5VwArC3b4o/Zz
3QYkiGwkGYMsuglFSQqhatrnJzgd///QvnlffTZbGsuhQVor1DKt26J1Uc+HUgd3
Zuin/yIJ1Ys6mMKVxr70+FRMAJ1s9ZFNcwJjh3vg/T9ANy0OHAG5D8k0M8xAUax2
U0fdHQFZeiB/YSxJVcTxfTvvNgOmQn5ywp0/JK/2sh+SLPSYA5sLKzf1DIDcvnzk
WY1CU37ivvUl3EZ5/v75c1wrOUdWhzEuskGq7JAruEXnA677XsWdKwVuVVGKDH0R
Nb6v4r6bWg+dQa+jDzs5NW7o6uGgBEsAVL0rFLkpCOc6mhGJcm80aZ4BACGUgwR9
XCqE/gXejIpYH9Garfc4DmEDuxqv0HRCvn2j+FyTC8hhjIqjwbfYiZFM6M+xbqNm
iXmd+3PADz+b027QAzymYSURtfVkj2EdY5iLgBeZ6xuamjRxEuL9YTZo+jEx/Iua
0F8JugzDKloJy26bhf/k9IDHMBXdkBJTeqmcjAVipusCoZvBGY4G2ZjNeEDE1UuR
+LUraexcxX6UlRoRnyQSMnoMN1/a/p7BUDza+FrFACrKAol+BxyvcJc1uhDw3qV3
i0EGQm067szWXo+XtQqnekgA4lCwjZ6wzyCJtoSWCMyB1VmlGtKppstd2XnE/Jar
TaAJYWiGfNLRJe3OKfPIeYYW1OQr1OOwpt6RZKFVkogXYocP243qCTuSLwLlkDFW
pWqoXo8/1rsm6cU4EbelHsPXMQB5dRCUD1ySn5pA9ZFqyBjD3YBuG4l/CuJnlmQk
JjrmrXaKi+TL4bu8n8nw1LKHAHaEvRDpreGXMBidaj0R3xYJsYW8FdUjzrGvUdKl
nDGf3EAHkEdSQt5uB44Bpa6jdCTq1M00x/nJzy2HW8HX0WXIzrleH7IIk4+bWWkw
s1twMatTNcom5tLLjkURsW3PIC5yq8vBlzUSS4qdAhOh1CuqWgmxE7xsjRGmUu2F
kwmsv+j+YcVl7oM5wuv2SY7xZ5G2Et3prH2xxuhFe3Tw5yF5R4gsu/kElcwHXJ10
2cFKZTcbnWIF+obOFcptJfV3YHxJV9SfhZXbAVTdcavfjhmXnmhnZ8TTzrPHefgH
IPFa0F8tuQHRlKaQhVpAN31/FbP6EhLARTK2AJkES2qPH9xyJ4vgokm59sWxRKFh
ZB62nl8CPP1EJ6qTJrcfu5U30AMOqh6zrqac41XhzQLtf0Dq7yjPzyi1KxlP1SsN
+fUKAEZR1rzFt9RCumJHx7DuKRpajRfwES1Y1WDnPTDuJ4gm4Sto9KUn3MDlAKfM
HPoZI0AZKALXSVZPKk5mZmZjAA8K/UFtQphi5LgLARs6ocgb6KZWizKimn2SYSpI
q3VkFTNZ5ryDIWYb4Vtg3ipoHv6DZBTu92mNt4RB7fkNiAX+9W2QCsdAKxzrgmSf
+2jpp07he5XCt/9GairGe9sebg5AV7Qfdn7W3RrtFRnRjVSVRcsMX7mbywNUQOkp
K60OCcFsVpDAC3c4cgvNYZqUnL/sVVo182a3MCpGJINPaq+JQC4Tyx7m/7I0KNZB
fKB33dCq4ZXcGOsPW/jmOjWD4kwWe4k63Rxjz5AlyudYuOJHAnjK1RckwsYPkSbK
JhAW2+EA1aocdAtSUqPSJoNLBSMygQZQjA48faS2g9TzHgLwFot2x9WPLsSTVFib
snmRRzwB6XXzITX0zu/bbxp6AWIJh+6GucVS9Rd92PlDKILOJs4vN6xYhvN7OKX7
LHOVuFx9a+GOCN0IaqvtdnyEgSn0I7WFSExKgfhFJPRuD0HQqUPjVdtXMbKBkocD
/7sgKBaWVYBaQXHHokPXEtlfdT4XV9gUCyoQ7/U/5X8SvQSP7LgU3aVbIboGfsME
DvSdQ6zAt6Tu2ooJaGCNJxTorwT9HNZe6Fpfc9taH8sxGoe4vD+tlBtWT6vydUAc
Bw//+wocWnukoowJwEayZh0KSeEL1dLKn5y2pHvP/qxjz2fHxp7GrTDouHUIpHPZ
wMUVcMuUE5qbjCtE5BstO3lRw/GG6+0jJpkJk5duoS8ZaMZI4SjU2g5mj2iuZtR9
pZ6K5HBH7mpwzGCpjxM13VEjvlQJXZOpisX+/zCcYcTvQpMcY/3skkqkVloGHbRi
Sezwuq2je1V1254GsoiFoaclf4/cL0kcOeN4PkGAFJ0rWL6jqqGOev2Yk4GtnNdO
arDfHT+LfRbN+AlneKHczMsOQVjgZCBCj2vHe8oQ3NANBgrb51oSrfxlpoxKfnEk
RnGI8qhYoePdIPlwxz8IkvC5XwaueZ+0vRFare51En2eERNeMNbw5xC/Ivegu4x7
R35hxr4UHqdKUMUnq6zZQAUZItmEbjPtrIBM4L7/FuKoBHj7gcJkDBV0A0NwlFZJ
RIyNuvePpDvQjAeoz5lnZS3Vkje7AYMqMPPYJMCcWKIldtbfcVk0R88osxc3SG1q
YN8QHxfdxTYLt4HBnLWle7v943hSir+0oJ60AgCRhXSOiHtQxbqI3LRe9/d57wMW
yain5zmqa1tF2K/8iKoAyFl3zx2lIZDZauaXCNtuMpn847ldgUfACI/GxPOz2jqU
ho/Rzv+/OGFWckP6Z4h0DxVKBihNoOsZlpS1GVjixDHg9ZSlcLcKNFrq0oxNWdJS
23KM1ETibzMxEUeJcTQuU6Axw+N2vxozNK+e6smD4WvtdA38kWJp82quQ/XEtDHB
3TOm7/KBHuJXys5s90r8ii+O+HrvFAXKkoHD4E9uPTwhvXdlp45uLH7lKzesoeqX
4pdXh/kmkloIV4rg0w7vAtiocuD0lvxxdE6D4HrHtmmTMhXu7u/IcrubunqwXiSS
Wo7fdzRcC7zVfSyMRfbU1OyIHVZM6Ehnxg7UreqlxpukGy6b+QgEw85P+PcvHxSK
qOsScOsx/O3cmVGq/oHSMsG01lhptNnSWkfQCVsDWM+T5QjklJE2MrFHKsdBjJFH
FwlahkuLCH7CS36kcNGXgyE7EGLUzNruSIyo+d8zwHW6dZYaGJEruEpkp3mm8gGT
P5i8MDtJFhkJoe3cj/8ipoJbN2PY4M/1cULLP5JFzFJ35wU55HtgykivUI5gzbm0
bXOY2qA8wmsCyF1Hm1xD/CWfcHgCQSrETeEpfg/oNUFDD05+LM2op0tXivMCZ0Vc
HKuA4z5b4JUTKa3wGBD60SqVSY6iY24zAFKX39J5YSNtz8Bl8GeLeDpja+2JW7AG
SBq7a97R57oZNVFOcErqgkKLK9JwA/2wP26teGtLWPpY1zraIoy2bHf2E1HukIzo
ssoiG7/MC/iG+L+HO7QwA61T7NDDP7VsE1creki8FOMFtREItGQnjDALP0Ir2OzT
ilmvrXUouA9U+pHwHHuY12Z4JrynOTkKw0MIGwUDmBfd6tZqvzpyKr7X7vyEHr/M
YEMY5eY+kkVF/uFp5yskZpkxKsryKuN0IdsRJPwH9nzPhyw4qvagSvweIprVzUD2
476HCW7uuHlbZpo7byM2/2e4omC9WhX0B1H0KiC61ri3j1lxRvcsL8JykK1mj+X2
OpDKyiHM6ViGvk0c8zuaUAyf1xYrQDjM/iUVwKPj6Y/3G5G7BiYAKd9a1el+gJ89
3NBJcZWbtwIpMUkyyUIL+NLKKF3IwyNY/aKaSoEzEb+xDqc8qeeYuW3TIyRKn2Ii
EMUgdorvzMBddi0Sd05mXOKLkIPzq/zYwgfVveIG35f/2x052LxdZXZTQjnqNwvj
AczdigTruRE/lOkn12W+H4pDLtvsXYQAe7lzmAy0h1LmyYO6tT+j50WdU6RuMoa5
Xbs8wIb+NakSb0Q4y+rP+wZiaEMITk5oa+HxVDmPkqvhKpVZxbk9XcAl34OxTYME
XAdWbF4gY4q3ZGhFUVKVHemiAfo+rvJLSEG5QXvb2/WaPCRifGZjn826o4OX+Mr3
LklyBaqA5ovxYy4ZQIK289br4tMlGxWFajN15/GlMlaohZQ7dq0i6pTcPzN2dUEo
wYaS1U2W9xGc3CANUmDn3U0IsslEG4pqCW6g3hrHFibAMpBmh4rkpMnBKFyy1WVN
fUuaRy/2sQo/9+MP2RqQlFMb4gxYiefrCgOIhQKo+P7i8UKXRXSVnVxdV16lhIsQ
UNsUk+C3+TnLEhoNFbuhFejoxJ2zTy4d0Re9ofqyeT/H0BGGsdMxv6j7JtuZXGB/
IqFFcoD4qYV/4v4mbvY2xTziXhun022ntTt01endY3sGh1XVqztjACLer8YmTEbO
I9YWzrKWAti4lHB2bZMfcsWNAAOJK2uRqgnPO2PzlcryQEv8usuFRmUR9JdaXc1p
KtIjKd/ICDPSb8jGlAPdIyjFWJ0t+oO9xOJLl6BFNsLRJJ8Y2VJrngOr35zXT6ad
BzVUcJeySPjY6RGPNpvEKeM/r1nD3kUDPIEf2nAjPxECMJL/U0/4Uq1e1tjN7Rqc
12o1Rp8mb7jK1KMVvu84uQBV5uFzAewpNYie6DUhJyzDJBY6/XQWWpgscLCvJm65
XuX/WKAsaS7pjaAd1/mqi2Lag7bwO9xiuTN9GQsnA8I6byp7ccIBXPEOjO+vwdXq
AKq9hOT6Sc7QksEX5+5HaBNdVyPoWBY5cEhyCgXzeqxl5JLvSItJvbBIRQZejN7j
OKkTzfjtQOuoSzCo6qOD19wSr7P+bqaE5Fr/jcHiejTr46J3Ss8hqcUJ/58gcqMx
I/Se9JF+jEmZR7GE2fXAr0uumGKFYpruTIWk1xrIR2tHuI4bziNYw60BFgZOzPpX
KIdhLjftXgtPIwcDecic13IaaGcstIyjWEuE4SVXnq36bVQG1nw1hMXCydbkWIKE
5BidpeOT0R2UjQfoHXy4xR+nRunX305H7nRlHUmDqOkVrErfbCxstpvQi1cRr495
y+oJ2EV852ldMRjFPE8bpekZXq9WYc5d4Tt4eRXVs2uK6j9WOBFm6e/Z3ENZcPVE
u2TpIhB/RGkHTtINQrl5rnYAv80zZYidgMYYsxrb9/lue2Yx1ngdrj+7ld/STlyn
fsBqDssf3od46TDqKsuSMixfHXdxZ90ErWNGvzHogsQvFHeyIg2+6sAIPd6FJv4S
mbHRNlePWPLjwAghcfRxEDXfzNTL2Zk7pYcIA1ntpihQzOMxrlB6cG++/7Y/VeMk
plfSW/UOtPFVQJ6XFx1/Vh5RPohJEOqLmn9d0TKyA2aClW62ONtar8qVdW4rY8G9
zxMevt1UJfji22g01yk5FgFRLtuAvC7zlp665VczJIqQ8OqsnnGTLN07cIt+S12E
`protect END_PROTECTED
