`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QTeTn6B2ZOMye36GvHdcCXDZwX/D4iPFZGNQ9zYZ8b/5I6gABTJgcUB4VKQo8brs
Whbq6glzeq6V1+z2jE4BZdIiSPq009smMzchw9/m/gArFqWkAVoNRJ6w3YOxbY8A
C8tme6v4dNMmRshKLi17ZYdQ6NS0n1E7nqnAJER0QBdflXAd+KFUoYnShSkOjsA0
XeHa4A57k13RrijmrnlRhB7wdYLjfQBO5r7m/8JgFvkxa5dR9a6JnVe5re3yIPlI
z3ctpflb+X2MSKfb4hYciICrv59uGQOBg5pTPbGolaYVAKWCQpoWoTVE/MXdmpku
1I4kIZ6mB1ws1xIQ8KnuKhtoAfT+3RCN2+DTM69lJ5ckhrbSbEG9ZoKBGrJMunTb
qJxrUHMJnY9nRKU76FVm/Mwb2Gn8ybCiEu4+dd4n59Yy6d2lWiOFqr3M/381+wEZ
EWhWNVmlxYRaMrFs/hUUqpV18vmzStD/XzpmalvZPLS0tdZJPuHlHplpKFW5kIK/
s/NXwCPn2OIa38Q44HDDz+OYg/feBNtodSr+j0GQdC2ytdnEwGN6lceiZHkLpkmz
1odZIq4dk4bYFyHDYEGhUr2ZqYnT3JJKjeqIFSRu5SE6WuQSSQO38493WeZzoLad
4JfTD9ypffJpHzUB3HfMsZky8zL60i/AqD+rz4He0hp84gV6KR+TSmJ8PzjpYtBE
MTkOH8R7Z5rUcD1glE8NshIfNDxsT4OgPjcwSLzbrMNzcnihLFgXF0VZJ7tKC31k
pfYlMUCL6su/Ck1JB9kZtk5EY1fRMOIekP5Hu6qhSMQUr/Psn9IqX2FXzH1r8doK
u1ij9KviGxrviiPE10wa/hoyPLOp07qpNmmr4RycZpu8VLNM9t+pt1QJCYrRrNhU
7thihAArmJrSlk4fjZJUubn0PEv+3jvq2gep5IvDDjzmRyLrekKjlSepctP8A5NF
uqt2RyXgCVkj6FWIJ7yRBmETfN6p5TH5cSNdlTKkBgRQpuz3jf43ol0xSh2m/F3/
kWLleg4kMr/ZvpYsozyNg+TPuXqA9OuC0sZ2lFsBOipASl3rYf/fF4qU8SsSkcu9
/609AX71QS53UbXw0lTxx25tEbtciEbPnq6VYtutOJMXSCNeB15ByAvqOmzE7wb5
LdEwhcchdv4N3Lt2NK+qWN5SzOLOAp0qII0jE1ONryyx4yNSTtXFMAxF6KMvFnhm
Xrw30K7/n0Y4bndUHRNnDTwYNST46HtogiP5hGoulYglx2hZ9zx0cJNBASxyzSbK
+s3gj3kvo/NmO0lcZ6pvqw==
`protect END_PROTECTED
