`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mglAv5+NJKEpS0JNfWYugtaM8gJY8fCPBRqX2jpcxJTf/mneMwlaJGujPagZSguS
dKLsnaVU7qpHUcfdpIt0JNOE53q1SqlQ5WwTEMwDm2HZuXc6tNwg6DXoDhLXYfwI
wwDqxUGOCGo3LmpftJmi73LTrlGddNM44jw+8RBkSACAyUYmUVCTMuLZrjNNuwDw
pZ6zuXilXwzJ02CfW3rrBJd67iFSqE+k5U+wo8xjmNQcnabTb3ol5zHWNSJd+Lg1
uey+yc5gwei5r1wsltwdTIH+IRh171RfoPIpak/q1/k+3YCsdYSE8O0nLHIwWT/P
ewcyYsxOh85dturg4M/SLdzkDAaR11288VbfL9pfAWAWxazBwBY2A0wY50JcV96T
hu2CVPuFt07p2xha9+Nhp0Uvq4vxOmtI6kJI+3CogAG6SBIGQ3bcFtrlgsQArz0R
fR9r6oW6pxa93qbw84Z3b4HLsmlrKPXTXyu+JWOoEiAZf64TyI/VbxK3pSOf+sR/
8e5ThSkgF8lkVI0sDg/ljbuk4Lshi04Mhq2VGLKX/h4TiLdMWibzwfEo5UbuZeef
ExcTgZQBHSzQiLsDprFdyd80m4PAjUXeb7bCwAgoZrwye+WLhtDohQ5qrQXLKepi
OPLTIvOr+PIgqWdsyGnAsaLMIVYgyWeed2eQpsE9DtWEA6onxhxf7Qw4ZkD8T+i8
IJQ6zGWET1lfmHMqj5y8GP+Ja21EB2zMlK4MLCt7oNmJudqdFE8rWo0uIbHyOUGF
xkqTbyjlkQA7De792PbkKKATMnw/OZmBUqOeTNA4vCf8H2+k71aJ30w6ZccN2sJF
5fU/B0/pbGGBeOO+o553du+wGtvB8Eo0BY7Eaep1SuH7KbOo5pDBV2Fkzb1ESqzC
fcWU/0vpA0Afy2QzoQIRpCYsEsT+HI/cYNbm+uhXjvgRT0SESy+Ik9lK2MUXDZcn
wwTU4bSKtgh4XGzMP+RAvTSKS+977mroSRHFPxymoTKt4bLsb/o3ka5doHhwcg8Y
uy24MistCkEvQd0yzYle+M4n/FUEnH7dbX5gxGbOvGuPzwowXPgpc8yq2xVAiL0f
dC4pzAYRPkOiNXpI8xNLWwnqdJRFSXabsq3jhcObQ3rqd+4iRSE9pjQcIjmMDYxe
6AH+x24qIHc8Vdnpw8LBUY4UjpIwxWxHYvk5JNw9RXr+TIaQbknDTYXpLR1hUlll
iJn0vq7Bsit6v2/xlLnP3GxxTO+B74ljkKxYIO6SLJkGhbjH5GJRc/DRZP4tVfpz
uSjs8JHho7NCwB3HR7ymibx/0dJiLuXddYp2Dp2WT5HKDlkUlHi2rYiKgLYV+DrT
KQ1f7p9F9ODzAaKvN8e7PkHwp2csEBgsS15eO10ZF9KVgHlpyyXyfE9kAPuYJqzy
aWGEHfAD9t193MxLBkoNU4bCF3V1UXUxXCvmcNSnqKby3m4oNabHrDZClNdkkx7I
RtoeX7P0q8h+vJj/zsxWj6yzZfQcOvSDQkKVwcFPIfCBDg2rgRFMxorG+sB1h43g
+emGFrEoTM6H8Mq1Nzge2sAIeEI3L88lrVTiWq958SkellWIml0b1xAUz42Ojobj
QENErw0gjV6q/AcWgCqFNB1pE1358Rm5CPHod9DxvfRMeF1XwZEqM/n+l4Hop2mF
UTKcN54x2Vv/52xYhFTHs2qV8qDBjUqwzaRACMBYucPk3g1eqSrZeQE2EVThUTSz
1O9YdpeYI29Lt3R4iTsOWIFmeAh1CYJoOd6hp+hZKUFdcJ9GnsYKyq7VBG3ULbdc
SELUj/DSUv4jWAj4kec6GryB3Wul8c7Q3GKphI+y8b9+/A+cODqSYJcsjyNBiZ6e
rBwk+w76iDsjH7Y3rWXJY6bpjple0n68Ha41h8GSNZ7oYWnm1o/f4tSqe/yDION7
370+w6hWb30LHHcz7984hV+CvIOzKNGVocy1jmQi4RfynzCDj7RdtGM40xUk1bIc
NGiXEtr5BffoQgXjZ3EVFVjRBKo6e1myIh8RWQyHPE/FB9JodZd0QUr8Av2pluXR
mj3wwSJFBMXkcTJaa8+6QAdV9uxaAogIwIigW7Elz43l5OhtnKCIOmz3ybmIpXGr
Jp3oTrLzQfBx//HphuuSksswQ7uGAly+Xx1KYJvueSWMcQmc/J0Qggq7AwCf7JCV
xzMU++KJuI2vyennxZxTzPc4PpcMJD+vJtfAvu9ykKKH+i/DFML5baYlX2kRzQAh
UDTQeecyLiNGrvxz4dURWuOg6zbiEvHGj211EMqUERae3QXScQ+eJQkE/0STatyn
0tYiYf9FBAkqon399MLMlRx1/rJQJEA3Ekg39uM2BBnL30VTsSnln9XC88A1fETa
Y1bsJH6AnBZ28m1RRdIYuPIgJRTe/Fx1+S6CquE6P1GLT569oK1Sutfz0sJIrrIL
BZ3yAxn4DbM1P1P0fvuvdSPTH7J+xGNGs3SnMJvgKUF3a4z7KGpPZyhc1Erqiohl
WR+jhFEK63cLdnL+wRj81tstJfTQjvnNoUenf6TBK1yoGb3ttITFoh3aTEPdM2Rn
ZrN43k2HufjzgdjcMh0H2cd5aMQ2Xsi3wQ7559OmdjRBt91NKXM3RxHVf+NiCZqR
0a4V3gxofAWqmCzW/IUEeakFHqtzDOYp4T+SA93OqlJpHfUYmpf+HaWRci19Wcob
uhXXux+A65gELjLVIyqN8VCfhCanymS512pEf+w7TEHfjbA6dxjW6UNqo/jIiVwj
PmkFODMWFnxVydnNdhYZS8TWpBeW+7QQmDMspQDiebtvbogLGVYmpQ6RtWut61tM
2rg4cBeKxCsSU/8rBjMclEFJkuyxBw1UDHzSRPrVGgoIyWItTjsFl26t9L5//7NS
o3pT0j41EeS8Erf6m9gfUSbf/pXHP3buMXpL4fFAd0G6z2+NJhohYTJzO8r0RH8E
zFMCgLXrJjupFmdLsc0rfuAFCm7YSHa54msNLuOsVwLJgIIaUtk3PugObuJjK6n0
U5T5rlFNX7NVNOsZaWPLs3OyfKIVvEMjvFLRI0bGhzidCes57ZdFuoHpdQvpXNl6
KI4ioeCCZmLCU57GV+d5tS0Te2yPOHhPGCrgxAAMREE0tut3y2zSfClI2/cdXp3L
2LvDuWeMbANuuLulK/YyntIMtjTyMG3Vl91BKZihQlVdaA4YwJjLBqMXnYu3kYfh
1srNkh76gcPfZqtERe05zbBFQ20ZA/yjkUxw+LpkTzR42+Pc8foj2JuUS+R0CgtN
RIkTddKMuiNI988JOHwGgxMg9ACb4OG87IjeG/a9qxJ/2LGQlccfTjrB5v0DQrB+
MsGke94qSBuH//cPwZM8O1UehZlPfd76r9W2QJNq33a6uTLcQ127rzMvrGhVGZtZ
2QconlZOAARmcD/jDViG5DrMBe+uU1XiMf/KSbWU+8y+qU9/CQWJWXAC16IeZC00
mM9MUigGAt35bZzz/oKLTlVd75rhDPfZhuaO20fPr8zb2JF0Lew6zdiFUKaTo+sf
7tRNQiy1Z92Or+/N0CjJYyUam8qY5wFB7J5PeMT3cwTk3M9pbBAnKuvqemPXCpS7
yQ/8VNeUxAEfndeWOm5R2DiaO64QUGMrLc7hz9ikqlPIxxNYJbFKImIcOFELcumu
ly4RaQ7UNovhhAcrO2F/58SwSU65pyfhNcvRVIDzLhsxbowfVSTW7B0yX6TZaPXU
4NVNruz7emqQ6acOrvnQuetyZGSUd+w59SYppvXGxyrBr2xwHbphwXC7sqeJAkkt
hK1fpQt2l13uVYYeeVy6/YypG32jAvFoFRk/pUeP3eSE9X/HCKRWZ2CwbGM9smZc
Ab1rsPLqfL12QsidwfobDOH8ZxszPLy3h66UJ1N0V51rcdUl3GVdkfFqMb1+wYhV
KmwTB7ew45B2BYnr8RVII8wroCsqRiT+rKMMMLAq9VkSt2sFDAsTbNov5ANv3iZ+
0MB0XyOmtO8WRGTrCJgkebO2CX9h+1hFB6rW2oy9bEY7eoSXzCFfw9QmMMPJJLOy
XDWQu8bKe0FHrE1NDKX4f+7bRnGk1dB6xSBaRZRtqWQiADUPbac+WUuWLXE9bVLr
pXR0GmxRl4Oa36B7WpI67wp/zbH/LSiSk99cbGNEdbtBF63TMAm0otOEUgki3awx
USyg6BAgF+7eGYIX5u1X1rqVSLAK/2g8ezfV1a53361tvS/5PY3h7Iel6epu5m16
ZijQF3PLVWmUq1kxilRBnXrms95bL+KrLFXuSbWVGEmWG36pHlasRpmVio931TRN
tkuH2DVRSTD7sPNfe0mvEv64AGrC8VzYXrQgdDP02D5/BZKu6DSJIKYbR6bs/f+2
1br3d1jrBuiV2lJXBUJZ+Bj/m+WsESOuJV5lZzbVLzJhRwVkkL8PHhlNcy6g8w5J
RFgXfF3+MKbURjlQBQXoP1vF9xhLEKVgAOdmFMpWWKhmJw9dtQ/B9nTQBGqEpzH2
mCf8sqvfUDJBj9w13vB5EQGEgMK1s3k/4MgvPwawWeCv0tUxF6OicAQ49yTpgoe2
T7xEJKaOv0s+R5knjV+tIGfuvfY2Nedd+96ZOnDVeDHXBmW5oSl+e+tWowu9Vm0R
iGffjZdmIzKF/mTKGtZFy5Via5egWJRMpeUufhoxMMKVHhZuQMsn1aLlJQ5OODlC
iSg4dQE49dtSQK0z5FRqNVKCWc4QUbpiMe45/ce1wBQDCuACGFF7mEjMmdsnW026
NK/rvDSbEWyyQlc7IZXuONu61zje0ed4N9SQUMz4D0DGHTFdMCUGXSbQD72bL3E5
zJLLoHhxV60fv4xppTi6swdoj7Fld/LjSsBnh8bHRksqCnUJOroh4BMItXwMe2sB
LCC/T8vrSAFBjyP/EAmGrJ48C8bdgCGL7xUKYD/1jfr88UhqRPJe/ZB4m3/3GqkK
Em5GGTFF/AdDqkx5hZfAGQNx06zx2FZ1imNhu0CGHKZKudCoasWiWIHChtzE4DRd
G5gaDo/9c7Ax/+ZsrwZvSghLOXCQIHZE6bDlX9e6bbGxhz13PIgTLPS0HLUPi/Lt
pdJ4raGFYpxXrw+zitH3Igq/8X3njTByUfNnnNdEfUyQ1sAjaz46pNnyJemxwPDd
rz4msgtYOC9EsOdIVRSyqCgGeuWtOuD/oMfH9LLd/0L/B67AvC5/LXhlo5sq6tV2
GlZwl6wUW/AePcmGaq5ludqyGNhOs8xYqwzpY8v7zEcBrG4JAy2U6pOpwB1V3H9T
y5C414GIv5hFV1Kyp2sgxK3G2grnStNmSpKZG1ypZzhcHuEoHflCm/G8c9xq2oA1
JUbnqTka/W6FLQAWb88fcU0syaIUtjRamShU9oqgfr5XtEYVaj99pTLVbnDoFJm7
kyEOy7Mi4Q8P59mFQFXslFHr+8UAdm20Q5qBp7cAp+N6rqozspYQ1aLT80V6yCdu
7UKjnQ+vw2TGnMM0R6ZOT7fNPwFesaKbK3Y123jUPkK9BAsPtgEhQFMrY0wVwQx+
Yts7wtIP7dtPL+iEU4lDAepcc/4iFPx4N1Cy4RlSnO564Hgl5skHeppV6Mhm7Bl4
aUV0IjwjiwSDh4uwYDGHbZ/9EdgIuf+kymMEo3xSvXk5Q5qELYu1d36J645n1c7e
WGmUZ5+IMLFqBUoouxyR4FG1N9edMQ0dQSrlI/FjjrMPS23sieKS/tc/fxzgcriR
W3zh1VwgfX3YYS2JVDmJ9S8u/m2nnLwkDdk2tk9cpVu5eP4d0Hcz4g+CU5eao8/T
HJUImPyrJeIEGEpG+918tnBIDYRT3aZQiV42P+le6LZPli5JIBKH0w370Fa4RXLu
s5W30FWQHVYHf4LX+fjY4GQwsMC5QXPH4f3fjbVTqe8keJju0kaq5oBFBqeS/+5m
rhnFnY/qeygmr+tV5teX8q0lP1ghbXtNQi8ZPSHML/JvYyQRxFF9wV3V7/G20usF
Tuzy2ypdP6M1hWvjvZtbFOvAn4d+GdAH6ozalwQA0skv2KLofanZprev7m5ebJHE
MN8m+I7DQkMJ8PA1KyVSWYWcXowwI1hfTsb3o9rFF0t9UWRv37RpOGrPqMu0QXJF
fPuMfVJjcqDFDHMEPOCamplBLPHrTn52LP7R2EbET3yUT3u2IhfCWY+B0CzE7AAq
o0mvjVJ5ZbYQAISwFTcjNjK9fXAmNs7KjcOQlZIqzFxV1gdzxmHLg3Vs3YIpdiwx
F1zigC6ISZIOYx0rQvcsSOnV5Qshj9+OO1rNkj2r2irLG7D3PEsamiWbissuZ/Ic
gu9Gdjft5lUkqLPqUXzRyforJ2UWHuabO4OcAFYFFEQr8ZTV7TrmTm80+3B80ZGh
o+Ll92KdbUWVFw5SfWyuo4Hmj0PbzLO4uby4Z9aw2iRX8eaHMrsTQi8ybr40AfuT
PCJilc0n+FvK3OvtFyobPW4f5nwoebsdwyWRxWvkAqzigY4ehs69Y+OIfn1Jo7uq
EXQb2Yz+Um60BQwk9/vBT+ND+rqmbaOksnsocU8dZlYOn5PugLQFB7WjBW8WMx9C
DgXsfShpZkgQvASIZNgFUPkxYwNuI1jdfbsp9CLRw4k497BTSbv5P4zN/TxCe7zd
YWv+ndZikf1sG0QEy3heVy7y7KrAyLSyYYHsqSYKjLIodbzH4CGneH2/+F4rPO4u
4JI/c2tfsGlwvYbuiaI7P1irjX4AlJj7DQJHhIygJGB0lIOGig/wTZJvxIemlCly
VsAWl7oG2/+ye3gbUV8Cx2dK19zJAXSzUufp3jmM7EwO8wiE+I4sMM8+NyKC62Mz
+Pgv5ipqBP0VTWp6vAsfI+7lTg/JiONlsjmiv/JiKi1HFMic+KQWIiKoIZsD4tii
8D+zad9xIoj7e8uMTK4QAsua4/BwE5bk10T5WgGJb23GQjljx/I8OK8MqBXeVi7F
VzZU7qZIctkxK6mvniEPz4J4uRaopx7HK+Opg8U/5oITTzbq4TemGgkSTGxArSYc
R3+vcH270l8X0TtZgqIb5ok5cS007TIzA/aLdP0QSQd9wqXjRlKX1/OMURXWO08F
/BGQxyvSWjvKfOUmp7IgnwFXgoLFIylQHp2pJEBhMlBs7bM/b+mYAVvNGT/fpN8t
sa/fy4Y3f5xWBpnAYvhb+5lHmc8bkJT9x+qrnAiFpsvlD5s8Dd3ZTSHJkRsQfJAo
9cvAwdK9LiFa4nVbqPE/WctxlLutatCVpXdb3UXwq/Ng0t7ng0Ibuur5CibFszel
rDxQPeb2W/0GiSIY1Y3r0wYFsaMrePIy4RgBesFXrISbjWDcNuC7kz4mlaRr7S0P
3Ha0FBqGKpR4Js+rlNE3x60eFLLkFH3s0sCCNCZcN7+P5gtfmk5yLVeJlm7qqob7
hiX+BL0QYOmX2k4HpiwEm9DDM67ux1X0G1oizE0rgAncsO9nBNouZUh9hJoaxXP3
vJeETahOg6WoGcSMhvvBnpH1TRFZeM41ItmAtHiqXhAmS1f24B1ppIbb5coIYxOG
ssOVNFNGpndvG13/7ZPxLVwFkTu0vDRhd5BYNJa3mLuY8QHY/1V47tMP6pMy3Qbj
WbwJgrNZnOvQl/p0FOKS964RwR5DJ02UcKBSbbPxwt2r0eBo1lUDy119TmvSKW5q
DBUZX0SZ/TA2sYYgkV4oqfX58BLHy2SnJgJSmGQHXiFZYezjuGpUaFAx0STp2MmX
IjfRNH6peYputRFy+0MJUMn0uGps3Llp03NPktK4AYKQe9h1NaJ8eK7czSU1cNJF
S6TwjEyE+CFoeWpTb5IaCLqITnlcf9pGsoYQu6uA8XBmLv2yW0P8Ot9RPVjYkbCX
BgKko7chPFQoBPgl4QWHmoQfQUT7yjFxaprmMRWbnhr9CW+g5eyShIn/IrJT1bRP
Ey9YACjvB5PGCFfQejNEsNAZpFS5WenwGTM2Nt2T2XAF1nwgmdO6wz2hYcU/do6h
EYAN6Ar3wulXvD4u+kLD+U+XJeua9zaNXw7RPhH3ptSXmOAQQyetWmsjEdo4suZj
stmEyDFlJO907J5NoSSjBxue7xVrXI2fL7qBXn9XqsMik6AbLPV0rlr0t4b/8Giw
5Tvfhcsle/mWvkyDL8/7R748XmeSrJlFQcBi21NyiWF2BIkz8/h/JtE+Cp/uO7ts
ua0OLNvrj+TLYwRKESvvLAlNxfKuHPjk2lEXH04OaX8XT2rYc6NdhRzT0ZLMT7Id
QlqDTC98HItEU39Nhqv0yKz7IkbuzmjP5ZwR3YvaFyn9xYoRMmm+8TaPrv1E3k/2
8dKgcnVUkUmM3w9gTJqI3a4n+GcvaLA80dBG/Kde91YimNMABvStUeMX/tyyCf5V
nj97rM3mk5tGkKr1FKa/TncbY5ooFqB3uNFawe+WKrPCY8LDLar8DUeD5DSnlWOT
abFXnAe+2SbIrEfllV1xGcjt9ZGfYRJyZ89kmeAZKtoGUnQ86YLRnUjGSM+wC/aJ
0fmsTSlg8ZjCFgAIDPLJgqQ0u20n/bASrZJocjyOmY3G42zcdKxrGsJfqsWVN8mO
EdZYEizGKOR7ThT0icwzq0FVf7/ltz0wzZp4U0TACcRlEA7VYmFh0rMoh+o1ESCu
+cA7Z01xwlMEVjuCn3GussLEw5iZsC7awuHlaz2EyPSzhWFHMb6ylYtIkwLwk/jj
9X6NQ6MjwcnWjgMNdtgBICMlCQPcvGRqI6uXUtK/ilYUs/8NU9I1MDFIEv3MY4Dy
87Fue+yc2dv7Cso5wEwO+7vL1wYYZmBk4KPp9NkVKP0x+n2UHA0VBwz2ycgezcjD
/jLcQg2pq/nTq1Kn++sJSKdGQ5AaVYO48GilMohUFZ9ZIxAWH3dSsjFg2qvJRo1m
hfQCwnly8+Dl9KKhUEUEk+fl2SooWGSc5cpK7Ef+Vn/2KK51qmfMMoKP4NsbnJs+
+2fTg9rsLakAqb9LAdWm/mBdsVpZ+mlSbyGvL/t1ieXZunyrJaGGWt1i3tTQReCi
AbA6+2IloMdvMmO24sO5hzYP05ZhdGkBpfR+NgPhys1TooxXZ0bJt5ReYBNng+rk
Rtb7O8VYDGd5muZ7yfS3do7zL/Eh88uRq1ycmOaBtlghDtKBv5byLp6G6dOwBAEi
HpBFqWz+7spTl1InICEdPMVS93Kmtq6uNUyJ+IYjjyo1QyL72aZTZff0i4c/ftVH
6qPDD+r5OHrQ3jHM8zruObMgaC9IWaMO2oYeppLCdo6/QhK4fKXV2jDKgEsTtxxr
rX9CPxIhqHvY7Ob0cD6YH85v9fEh9xNi5Y6z4Ov+nA6NYptOblSO8uyIZ2nnvwvx
pRBP+7wQgmW5sj5suxzrEPYjTmmUb3L5X2c6fZ6cv0n0vhFifqRPKzIwl40o8afX
9AIAmVQ0dVn22S3YbIrWGvO5/CWnB3yG61EhK3vHqFPyCoz4uxzhm2SxBJZahmVt
cyIooxhLW+7x+p7w7myiCeh0sK9Va4Ksp/DiweBiVlAD5VlcRnvrOsKSx7PZH9W/
25QGuGniXYygdB0eCTX/kgJEIcQ0ydBaAWZl10/zmNdQKzrzChj6mQ1DanSbl3g9
4ZhhptoyQ0Am3JX5ftqhJihFvNKhOQpEqTwzSmfaGCtAR1sx/R+lDDFCcLpyQj1T
pbCO1CL5W7JiirY5ToNUsn1YR75x3wxzt4DD3EXAwQGmbos8UfCVyImVkeoKFDY+
quZ1uhVEpVpBRnVfDS49BRGGZsYb+0Fyc7j/KHPPWJrTf/v//vwYY8ykEHyZyZVV
y4EC2H3QAinQxzSnFimtjuESL+2c7weRiBBiU5CpOwX0pZHRN28EUtUNjHSZMwfh
fEF6YwykJPqvX2foOh8f9Ilc50TS4gQywComLCeHUXmqBtsUOU0j6wIcblYKM8Wt
0g2c0gqJXHA6CHmk9/OT9XssoPZ8MXKjkyB15D/x+K61N6d/8lbZJxZeM7OUq2Ns
T0mDTXKVkRqphsFbSY8HQ55m5OVDl1zJ45i3OG2+pzowUZLb9TmxBU5Uzl/JaD+0
3+aJ34tMAtjxJ9yxi94L5fhzKsEgPKbhDm9Rqk9TZeDQi5sZS1TCWiT4Eeb5GlHl
LuxPTCTk0UrWHf8ODgT6Isvs89lp9A2ezeZsiZoXHT2D9MaohjeOzA4iquiUBLCX
b8IwW5mzKsPECkZD9MC8ylbAdAX5NmViAiz5VUngYcsUnwcS+0ImcEjy9m6Tmq2F
ChhBIluEfBz1L6g08Qduev5TzEotCLIHIn5fjR1bn44cvDme2yvSFwDbZ5/U6oiu
rdTtYHdRSQuX1rkReGScq/COpgheFV4MCUfYJD6JGyeC4ePnKR+9htf76KvY4zEI
rQABi3Qce87D4UsW/rD7aVD7CpyT42MOl3ASsN/mE+0gJRjwqxGJRk4RFX9nfo2I
XwqAJO0fXHyV+SJm3hldB3YF3ubRrX7RFCq+X0Zv80825y4b+fsVTOPJ+uyZoPwP
KohNhXoYBGcTdo86p+Jym3bNZq9nvFRkZYULz53rz3/lI21pLV9uRbKlvz9bGjBq
vB5uAD4TSHgswuZvDgY5XlkjkggIbE9OCNfqUU62J0fq4nZfJ2k6ayRQGEscj76g
qRxhD1JtW4rn1LdHdOqWvFarjZNHNu1ko6V//Fd/5c53gCxEqBkXxy0aUVXqgC4r
KVn57DF8+UlWPYKCo6SPvwwI6M5O9zFBiHPGtniQdkR7nNw4vpfdpvF6sd1Y0zjT
s3tWtvcHuAU74ViIYYoLmdlDsxxEut2DZExgSHpvGe5y4UrifSx2RVNkto72w6m9
vjW34zTxUR2/Ptr2CxQHIcBAow4Zt9zlec9gjVjqvM3P1gacuvV15Igc1ymRGv6a
sZZiLX7ZSMPxxOo/tasTZJn7NmPBTsByVUShAM4TT1HbE5ixNB9HgSD9d6ivPwf4
fAfaKZoAanGBGOCFsmjgefyWM3HKB8M8ABpt5owtaqsum+4Xmtqb2MmUXHDEutol
+5qqV1fhT4XGmnN/z1LD+HY3ZQaDNfB04vqdy47zGYKgNlxMgo27Y97yrfFh2/P2
PVi3oimW/8nPxmoiripl+hDv291mUsgS/evJAEy9nfsihXyAiDBtJCOEzUYxqxSA
KAFW7E2RdvFpPbjdffkGVAToRCKbwBxqwTvlG00byjlu9hQROuFhVPGg0deGNxfP
4lVRL6zn1736D1b9CK748DpD4xQkuy+IQMIASdBLfsGJSE7FAo162j/3WaRk1nUU
LBOrYkjl3XXL6EPC4M3Q7Q5OvZ2SjJou928dnTOQjaOywgh4MmI+ayRr0uwKBLqq
gFa4NTY0zZSFFsGMKz9LU2xqlEri+iG9w+XtvJsS4ZKpQ9jVBl2QD2T8U7nc1fJf
+ttUuAWyZM6V8byeIC+ly94Mvv1HVkKO5ExEITdK1JIIeOLJF4Sn6m5ikXgDtuz2
DQo8b8uSSo7WQ0az9nbVMcofETvkEBm2D1g97a7zsn7etARMfJdnnKm4LXOd4Xgz
RlM7IwRS4tG+/f+a4mB6I8wyKcVsy/Zon78k1zx6g4rqI18HOD5cQmHyo+hrlqUK
inyy066hVn/EnUvaZOsAY8ctQ6UQ8pwOgar4qVlCbkz+drZp4O4UadVh+BmPsKdi
uk8+gSj1tPepvJD/6+DE/s92oK1pUgNpRSv9EFhtLNIHLEI7VsJ+/420YaNCsBKO
LK7gLtQpwBuXPi2gQOZnkDHQNwyJXIsOChobflVV0uw5VBfh/Smzc1Z5zHX9BMxL
ednXcDblxCB3KIfZKWl2wqLUUQSJgrHi9grmRLtQaFZq51ekr7/NworFNInyRTdN
aG9+YCOT7tpv3Lki656yH4MVsFqMme/kZdx6I/XzYGVWP9rOn4gL1gNA1j2DQfFT
2f5KLHoL8oYGz7wVNpsmREUci6ufY/GWuJWdrfFs3F5g8PnOK4PlZtHveK+0xGS5
3hJGCf9CbkDJueN5A3uB8SsotYep5JTNxpcvDSmEJmRiVPXBt1tElEOwrGN4uQNt
Pntmkv/CzC9y+4WjegQNiag6/mAKlzUle2C/DMHVPSH2ZYQ7TCIoEre8wWuXqfsb
GBZdgSa1B6rRoJ+eSqJi77CaPtaom/Q3akttun2cgKo=
`protect END_PROTECTED
