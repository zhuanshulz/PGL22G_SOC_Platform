`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gk3CX6YNR269Sr0teqHC07mF8mPjJOg+WYYk5X761CRBZOtoqU1IxROgXsmHta5w
VAR6DbeC+oHkwJG/cSFYzaOKSrhhdxPxjQO3NSw8SSTrGdWygaNiZ+n3ZcCfn6AL
ZNk/eIwbv2tLcmpMSYo24E2VsNn1LFai4EQmf4v9Mu4w0i+JuCf36fxUmITG3yEh
mm/LN00tAy0Zc6CT0sHX25keg66x91V1PvKrQg/eNuXGnRwAEk9Sz3It98xpuCiK
sZjFP9/rGK1QtwqC3VqMRHkN4RK12LNTIbHx4YO5/z+Acw3cSPkLaAhDqdeeNhPj
y4N2K2dlP+BXhXT2pqihPpRjc5+iIIAlGlPp1lM3zGSrxks0W4KHCyCeerQFN78j
95t3hlKzgVC+TohXZ9rt5fL26bANzYhFfcr5wH02EuOInMmg2XH1bk4K3FC0O0mY
tg0qv7bJZkOVVgXreCEo3BcO8YEUFE414MFLsp0s1Kiu0TgM2m+75kNFG4WznOqI
2LwmAU/n5DE9b4npTC7SXJv8jmE39N5TAvrQmEFJqBEXVQXOk50crBHYldOy+GD9
hb/MaoJW7mUA06SQQpBX9BScBPL4OI/fHyDAsViy5pJUN+13QeOPU24+vMPMnWjM
OJYiWRe+vgv/0W3YPLlUeOSrm7oLDkUN8BNWE066huDa4ZbyPJPbFAe5J7kJ1vYG
pSuvp7edzBLKsy0/5E0Ymd5HRtKyHBPePgezladM7Y9aXTberthqWw1wdkxTzbJH
MuuPFJP1gCYW/A2ag5Fw8aSLK1YUCO/A6TdNYWH9ANyky8EIcE95VGVOYuVHqJ2V
l7QzjiHC3NvU8mYx8npwVGSAbfYp1h0it0IoOjvkdbufg/5gnbagbJHeZSmavm6n
O5Y8MkPDUsR54YK20K5kOJntDSO0ATFVeOwPO7cXQVizUsZR4mAYCAdpASPbyvCu
Z5MSb0xdw6XWUcxSPumCORHU3bWvgZCwaU1uLERMgdZf4jP/kbaw0BmTfp6IieUG
qD5WQphIxJFZGtnSFTndBs9Cu1xzFM+gGtolLnWFKGriq4RSiNiue7AEHMsHes4s
aOL4sWFxWyFrrTSnZ+6TF/s3Em8tBu3U9ogX7fMXrD+aZkwkbZht59HAtF2nSmfQ
UXxQ2E3xaXW63UmyzpeoD8/BvMOgqUYFjkx8pV2i1+bGs/7+Qxd0qb5BODtHNm4Y
jkhejGLFXDdRfmV9H7WAY5ihhpzSApxLJngDj0sE4NteNh7fr9wTUTFZjwBmMf61
qgmK7V93Al/FSndXQNbv8AYkI9tJ3/lAcPNQw4h4XBOd4XND9WyG9kFD/m1bAEha
WU73OPGhlbV7YTg3DYuteQD/HUfwmyM6iqnElPkPTzFvu08xTmLpko63vx/nip+K
BNyuurymqweQEj58mg0/bfdytz7KAGd9teyS15DwiTsehxHQkX0Vwy5InEM62LO1
6gNXdk4i/6NkowvDVChkuk8Mt5JTLd4Mne+ZA/jD4A8CqS1+DV7+azIxKmLEERbZ
TOpeUORf2CunkHF7sUjkWk4+IZuPlvrjeHq31j7rnLfK3XZpLqVJrGdW8tGyfcxs
FGfZOKPnoWIzDPBbMibRrzyV4a36hcijZzkL1EpPafFFAeAjm9Bin+f79TCz1Ex6
UEOt7O/tBHxaffLkgyQ80hjc3Sg6ouNVhb4WMGQN1OLfpMTV5MqftVJeONxV72Za
q15+RWkE3B9aF+LIZMus6VDBXZmWxp8px5jI0wdYKz+y5wgFpGO2xwWDeF1DiO62
2AGW3zrxJ48Lr6qX10cSP/3HOHoFVCfQN7JGAO2x3e6h2/b2XD/PfG3uYh3Cj8QU
Cy9ZRiPtCLqSwLQ8mbBw8LKhUoMEDACvKedENqeWMChPtmrQAQRRT/tmoxCDwbdN
2vseG8iFnKryl71hz0EIW8kKG21iaB4aVf0B7g9Ed1r5ru4pU4ZktbHkr7tFXzUZ
p2eSQF6NDs5dO7Q5U8dHuPXb3H4KS85bPFy/M0TMvUZjp47Ggz2CVEh4hJB/jAmY
hs5dO33btcbcCfYi8dBhCd9CJAa00ePDjbIxboK3dwxEy6AXgGbYJlCAWkWU+AKw
7FZwQXlPfE7W9NcXeOCjP5mP/X9JJ5CdtN/jAOw8umwC4nzacy19pBTBwfY/Y91A
6u8qVd7/I/QkWO7dF9QrcbCMkMFk/eP0u5YhUa7YmUaEtkGd3jI4Q5vELbmr/hYJ
Ulb6hroLOtJN/RgOwmgaFMCh7uONA+/FX94+rvbZZQxTpX3B1LSMgJZeeUhIvZ3c
JqSN0MQhO1tY85+ty3mftqKG4B2lbB8SCafwT1+sJNtiWdUvq5RLKy64hYRFNb6s
PzDiH1NqUXcMFwDxPX9n0tmymeWjXIGQ8vw+JOUjlZoBQLKV41P8km8o/OLiHP2q
piTaxPeJHdT5kAWbZqwWMD5L+O/rzhky9peLDAB2aM1p+61lxnD+/yH3PH8CX0DZ
lJvZpbUcrUy4bH3imIkB5ZBhiI7tpKBPctkvcdAs6IUE4eehVmFmwV13pwnFDGZ4
q1YYWMMoGckg94/y7HktR1T7pISfpafq8Y5Pq+j6fdlkikIIY1QQJLTrEupsJJ0J
8MUsBMbeXbujgYsHSwiYoueSPYKfvj7pIhMbYtELBDqkaDhn7I5UT5OjLr1NPQc6
XR1ANuQyxfWdDddmXRJy3NU/CJ+O9swBYSOYPocCwb1nCggcnR3oM4Et/lQJ/42n
8pnJZ8DTzmqqhc5Sm+Ow2s9RXccKkg0o/TgJ8z7YSU1ybXSBQmnw5mXP544euVI1
JqBTfvXxAiPt7r11+NR1xa6skzz3kxjQ/cylj6FEBYeFv9bdHaomjpxVGu/l1zOE
cbxfLfbREWKTV0P1ahjs7yMyjEUqyRjUt9TmTIuujIPKfVug5k2tbhccGXp81ujP
qP6yUaGTjmbKiVNZc4camZMkCzmlVdRknTvKWCTnweuBMNlTa2seDZ8kAQ5QpOyb
b65i2kyTC4UKfaJzpFbRkMWBFQO7kbxrLHqQWMxQ1Zus9whXO8865s0uLvD12Oq9
FzVhxrZpquiKOdNXbJyVOV7Y6Fm/sUjU9zI/Sb8IOk/IaN0G7LJ7knUD9gvMynxD
BKIzWvPEVqqwXt6Uwyvh1QpUqNt5e0VWoknPQxt5W8cEWQ+q8xdRQz0VAweVc8NG
2Qf7eSdnUMOV01/KZMl69X58DR0hLJcl3+HDx3+9/SEZ2VfjfZfElQ7m4u0RiR9K
dHIDHk/KWb1JVajRD+qej4ZFRx/5nIR6GxcskjWcscthgssoZR8Cid/kciLIphXo
s2dGMnCkYomjZETlLQ/UWv+iuzII7Mtm3SQHb4L2PVdQWHO2kfWMoLExRA4JlIT2
mUKmZv1Ig+2BfdcMZMm/DFNYwctP9+2ba17QyRb3KIXNQqfiHE5QxtAl8Qj+h69i
Tg2IOwaPR2+xDHnODE7tI9HE872t/dCMycIynCUKXuOLCB/83z+8Dalv0LUul0Oj
LgYgfOlVt1WAyfF33PLr962C7bOcj3DPyiVKaCPbJdIsnk3Yq8L8fHsIFmjHHinF
hNsFv+nrJxZNJFnim9cPOU6T5TkdPoA1Nlu3fbCF21Z+oNTrS/NZ4MCxvL3r1gYM
//SqqCTOIgy10/6hQZ0liLIoOFNgfAngiDWB666fK+UPZ2Ch1W+8xC1eTRkbuTQc
ZtMJ65xIau4aqUGNen/lJxCUktFWQB/B2x6OWY1sTL5URFpFuGEC2NkLtBMAkkgF
L+gyDmp8BKLLplm4h7RoOWE+1vB/3CvbtCxME3q/frOycuDbkHORO2WeCZfQYgYu
qgEaaByXdZ8QkPBzwRjYVpO17VC84vY3IUf5MbFEo2W2Kf4itmxfBRJVbsATPHm5
9HxZkoggmB9JKR1l7Nrijyf91m6d097ClrKVa4jjlArg9ZPEfyBq5SLAypi0TqFp
d26JJxdm6B9IQefVmyTUnEQuI65Weq9uwsglGOflBnz0/1qVaSbCGh1NQRLQ84Rm
rcDGWxvrezHtw6QqJK2vjNu6tKWIJlYBOs/rEGLhIX9GV+c9ZufwUMxbJyD0AifG
K3ReEnMovy8LuDH3EQ/6AFb/jYGC+TVY68hIuCwDE4D+lj15Sidm1ZlhTpKQMpLa
p/Ycn9O9gZv8ywzziRBFx19ci1djgzzXPGp2Uy+B1mlnLkB3Cnld/rAXq456tztu
aGYy+QeYXYN7KkLEk4IsE0BQhyIqjLtWRf16vWzkd7h73eZ6jcjC+xca84exR0XS
qgJzeT4qrDyTGeWdOz7uQnNaoxxfF3YTuNwVOJ2UHqBEQPvYHcxK6vyzYb7e1nrs
aV9dPkxfYz8FTeCxGR1ZWyML5I03FnY//dd8hGi8Qc6JPbrJwYeRy6W1TkbT7/iv
uhn7Jlym+BWdpmxECfQLoMiRKMw8XlOBzLXIhkQa6C5rsKiK+KTfG6x7Piyrj1EK
rrDKqT87zfdmYTpTvc6EhIM5Ec80JSk06GFJinKCYpfuvkcDctUTwd0XaKNn3pml
e4eJVC+L/qXUUnQ5Ys8rxR/xNytzR8SS0vER2BjyV1a1v0Abe0MMb8myASwu29lp
5HdeHG6PnjO+VNV52MjwB6aQRCk689Jquf33UVq/iPj5wTD87ROpqOD0rt+MEYGm
3Jibd4oPofsnKDh5HQDVDdFeVka+UXYScjEL6FDiVXEP3hvjqIYbpiT0qGtT8XQB
eQ63tARRmcuqLjiPlQeGB2I6twVlJYSqPWboMaS3F8j1O+nExxoV7P6WQDU+M2wP
L/jzYSQpXK/dhMX6rmjb3zJzHtlUQ30VYNuaKGiOdeXi/9/pwyE0OkStBVYbH2KC
zb5dDt/Hp2ugpcYPMQYdz+WMyV5GtI4Xp8TEkSFvmhtu9+JrwVJcX2CjlgR9fa5B
XZUdI6e/LzLYynjUFXziMgXNh0g1iwXkmw89olHjkm827LC/FwQj1+0oCWr2oACF
+toroccZRhsMGfCGEgYxvnuOZNeu6GlPpNyCfIr+VHJH4+BR93sg+TyIc2zT8jiG
P3F1t6IFZ5CZOQHI+wts3m+27xL4zGKgc8PXIarPAxEHhhFUJ98dUGKVfMHkCian
KdzpYJT/jcgTcTKmyaxIspsgW1//2Ft1BkPlKK5HunNBrXDumuzsj6qtWZy8pcCT
EX7FrQfEvfN45M4WGcas4yKCS56MckzaaScDpMJqconO9k7WW+h8fGigDCDGNZ5T
z3T48mt8W4OeDwn3sPMtou6nKffEVqlexEfDmUTeR9IlMJ47FhxLLMmub3WmA+dE
CxgkKsQc3t95PT02X7YmaqDwDv562ZI24alnM6F/fd/0vDgeR4F+1Uh6ww719E7E
HQ/mvGb+bJOls0KXeQFCWCfJgULTvjp9rAndQ/x/FiWnhonh4S7HL/ovdClPGGzr
Au5nPleMFAzHRFGn6JJ6L96yVQJ8ep2TN98KiIFJcxKNEZyLI2ePnd+hZfB1+zBM
jmCb8b6pAq1yPmL2ykB2i5phIsFv0wCHk7ou85s3Rt+b3x8ULtXt/awUimLDyMpK
KLpG2eXTVTLP1OispoxciFtdSI+RM1OvVqeetDZSx5Pg1PjD0AwjJaISd3qWYiX0
CdLoxvpmkX+J4hILTOvnxzDL7c4KlJkje6Kmif3z4NjNIkrGMUA6PZelDaefsRce
n88mfjhyQyufXMq1rx71OHRxgqqavY45dB9bkpOM5vustmEfSgoiVvw+ylSjaiuJ
MoT/APCZkZEpOD6/wBOMsH+Q3UFfAB3Dd6Jjf5F/T4xA+l0FCUnsCvp/CaMBtOzI
rw0ABzI+lleYC0AyLcMNLXhbYtNvOxg2Fe0W78Y4K/faaBrBMyJR+FIlbDtaUdJq
YtsQTY16cysKONhd8rFy3pnOBSOGyfUII1NPwlKL1cpa6odaW3cfRi21p+90pv08
UdXgj5qH4IhQow7/XOk5Xv9drCxuaOKOuXEPHG8WC+MJlYh+VafyUYsp9Ju5sw0Y
j6jViBbuiOBNCPQNBHe41l5FTKV2Oytj/fUYrZ47su+FlACElP3GM9qIuUha0maN
96zQ50LCoG51oEUZ6v9RpwsxuFU9Fe1WO5TKRlHhhp0ZmskRzvC1BNml6uucpFjm
XBSPn204+xxD+aibzXms4kAFwodNLvEoufQ8JmSXme7vLJ7TImXZE2/s52Bw2eUu
qwvR7l2l60lErdcmvY/EDZ+J8UL+mMvt23QV/P6UHA7TzxXJM9QElIrDk22le3Lc
Vq94s0pgiNEN6KbTZd73rXZiyajobiojWGzzgPjT/KBOgK1av8pjWJiWRem0xrde
L3YBjKSfPbGyYJbp7nXe0ISCQ/UlxkxRmXggDnj3oGumemFXC1fw2VrwWGrZOtRe
sMBBoUR5OMW9FaX8ga5C3dobGVlRtofNGtHn5mHJJpW8C1i3Y+SLBYADV7mMYQWN
49mI94c8ozlFHB55Y+jBoXK+bh/pCVLgdM/UiYrxrZSZjUdze04b7g5n4PQrO6p/
EYfroC13V5t/PKUKzJLGw1+zJ2e1eRcjPtY6pSr4pwJT3rXFyxQdY8tvpoKKxVl2
p0hBU4YXK7/ivEGB4RVnheLcCZqmTl6C0KZj/pxWbWee1hCfE7eavfam/egpUNHF
R8YDITrz7OCcvV8QS5o/RRaXTj/cXPqPmdYfcUHMKMttNA+Ql0qnl1xPWCJhCQzj
fBOV+4keTU7VhYeoRuTURsCFaPJE+BNfOIlsODJtLjWXQyjZsGNcqbNJZ0dL8RJv
PLcWqYPElD46evDYWOCC5ZsNO/p6ouucR8KKkRazO2javMRsD8MA7nn7rGL8JcWA
56jtts/3AIYBXo/CGz/N/jo55ymyawAtLfLv/VoDi8H9KpTktvmahwMTWHtTCLKX
JzE55dgbtjSpjA+XxIvCV1eMa+CsgFVi4pxp110o6v3e8RyAcmSXqKv4L92oCWYG
jByrcD2lh+rd3C9hQRMVSVyQuLFmkHAvU1JBhQicO+qVcnFRWsRGhZwMDyYR03IH
DfqoSQDvHPQqWtiPwt7U8bT4luRwXCb0f1LXgIU3wTkY2vecQmvLG1Ot1xQ9UGn8
79qFEmGjmWMwxeqmhe4ARoSMjaFV4ktE1ddg59GMD8A8ua5eMPNol6R+hTH62LXJ
1WSwXtjYtldbNPBE+ZuYsOLDNvz5dJ8tcR112H/rtoRwF4SYEIoqVXJRY7tgGD9+
0EAoWYM28MnUDQuk+5qe3fYqkEDtxS5JyBzEbdm5LVa41HYAkG/mrrz2WNJ2Cyyb
gToEXNRe1JsPk60ONMsqUaxRblSP3VzSPdPP8f5cYIzV6KU7cnvIaPI1NCcwe7BO
Q5OHWB/F33hxI/AoXS1K+6NCWHJX34qJHZjsypOQTh2G3tvriQ5+4Iyjzj5eFGBm
mC6IVLJkOUUyRN57hWWntrh3kyO/WpGNQmgCiqUHrIzN3GymOrmsbKyFqfThv7og
vtesQodG/pUAGWS2sHZ3frTIxlfjnKQuV4N9IgNQBu9UlpGaYKUqTs3uHYunUZOz
l2ujT8l6ftbZjcatJjCZNkzOaEC1YOTMSxKC7yX+e5oaLu+qXLR7V/e5AAAr7+RS
ggmGCIwD7T/0DxyqfysxmblbFeZXIrdzFN1Fh9Ho/pCo4isKwJngm98SeJMt6DQY
WRDQuRzh5sei8hnymWiF5Ds5nX0iIeDCTX9nRqQfKcq5ul3VCaMqcjklQ2+Q5tX2
ofcj6rCEkOJCCVDsrJ5Q7St2y5WA/BmuqoGAZ3bfYLoT4m95QOz+dTJWmJ4pXZYv
en8RtVtAdua5mXIEWk95UmqzCDzi3aoj3ho1bJH5LLtgpUg88ZuMHn8CB30cveU4
IiqKR49wLW88JQYA5O5pXBhB6Qde9yV27E7kGQgV4Bxfkdn5khaX4sa7YUmZto+v
aSy5Ys9+e6o++0cQeITLZnL7CdYM2N187OiR0UQEsmJJn4BPD4pXyryB5EHUExDc
MTGlV1cM6vR7E5Fz+XSB2HosVwkE1OGDuHEqVQFYKTntYNg/ziTdX4ZHTNwQyEhX
yRj1Av6UP7z25pftk2d/EuJEorPwXl68E0cqauQdeKhXJ0/y3wBljKVyS+YxSqsY
Vhac0ulwou/bdBINqo/qh7i25jYJpbOI36GJBsVhu64mEpq8T3aCJVWveILPz0lQ
4+BkSaeDQMJJmjJsS6iDx93vZ5DmocWukW5lVO7rkTyFPaEbPFojIqcT2UDwBmT4
P0DTrUKCCxpZacrkPh1m73ohR6zJZdRnbCcdO1V2bqD8S4YinNATLHHl6rqlRAPk
UQBlTeGs5QarqfUDlSCXDQcMYsYlKMoNS3L48//Mjbui38dSty9Ixrbk3p2DxFQ0
qnOPdiQOGPuHh4oqtY3ZbFRIxop4OcW5/ytKPFYCGq1li3xm1N09OgF9MCPjbiYv
gPK1JV8pIxwXPGjOEwLVtIizRbP69ZJhIZlyewqcouanhFj/Veeo2L1mpsIfZX1l
BIHaRhGdghM8dqjRelD0B1urqpIFzPx/wbnx8sM5+FI9ZJt5sa+E3aHrSTYw1vaP
pdxcbidmy7jJhHcy3dqR6lwjxtR5qtlaMBUuXmR/OKGfyEUD6t5scafJ8vx+sbOu
EtA+uOM7jiQ3Bt/lRW+hZcMCAA4qbFOEiuhg+T0u0HEthusbFLkl29wc8eIkBhhV
2QnXZUsw61t9GCkYlwg2NMS1uKoHaUlT8TWtDKKK0soW4XMHPssk8Yh+MKbl9CFK
ZsxrqYG+QuWzkmMjZal3+aeJwcbv6Mb4j2RKqyR7TVMDO/EI8jY1UBlemdKloiwI
nK3YiLyXlhP8xOpsBIOBMvDA3qQn6URSpxf2k/RwWkrI8ARK3oEDaRnjjWtrLPg2
GDwWHKH+P7sFOFUgWg2rRkl0qtzF+w00g1+/D9KejkDAn8XEXo0134OQYCNMKx53
wIaIB2vBgzRuidBUz85vwgpaR12nxWh0czqm/dJi2+dAfllWqnBe4hQo8+IqDMgZ
bsxC+kFoPurGXsyoivEddE8y52nFaA/cgCgRF3gigeHWp00IU9BCbHD6hsgyr/Jk
DvB0OAlC+a6/d1NBmv0k3whvr/OZWyIq4WYxjOuV6u4/JIz7sCmoZQqk4DnucwUA
jE+RDzfefZ2MLAxL1pz8axoS2G3bJNAL97/rBJZHwlsAXGGM/AVzdDOGoHWlce6Q
dxtBiFbImX5EbTorO42XElz70iBhM90JXCwSbb+2gOoPjwG3cTHdBwCadR1nIoKk
H8wTzNernRkv0narwii7dqCVnqfKIwXw/V25Q3Y2Bl1XkmGSBQtu995ADxg+Ls61
HW/UAINJp0zMj0tA3NP/0DKun0aeKrdRJee/3P5/BfV10bh1yjN++1aVzS6sIA+G
BFwTz8LoLd1ZDtypLeUqm84IqsSc0DMVDOZSQuSf3SFynkD1KHDbRfTCEPz6AtrI
HcVY6prgDEP5cf15kgvwvuhT5xFi79BNZQL2NTjC2W0el2SB3oxbC2O23O7+vU7K
a78Ueb3JuNRZKqvRuewXJqHEEj6vmA2rB1TlebinT4fhPePkzSNJMNH/n9Pc/b+d
LXaZ78nO0nqR6cHgQvW9VuqQBxLUFofonms22GMA/kH72flBtIY5aWtDN2wV7edi
xIzd41X5HD4rV5yGzB7axrH4PrFj+i/CXWaFuaz0GddHwbjKqgO1i3qVkhjwZ/6w
al2BYlY/UbKiGQodnbUSI40XwZmZDmf6opz6fWxAL2V41kvng4aAi3YQFBfjrPkm
cJQ5lonSRgCsPTDi7mBagzGM+GZv9EKdtfPfu8lkD9g4CQRvSTEYVL4q7okEM9B3
cqtslAlu+D5Aw+WW1GAM34NCiauPBYI2gENva0atQ9KeWTpVpmg3YjiWiZyjIqLM
z75iddUXcquuRjmIP+OHPB0thmynmPt3RlKIezGdvFnJp1vMw0SLlqTREl8800Ek
M+BXq1vtE0X2erQkTtSRF9ZON4VGseFFBDYJFWppTjdm3URBl9hV+lMLahNieGUz
bNoY/MdAeIR7myGFUaGhIqf5wAyGKZHZ4P8AYFM/bOoNXU+JZe9olQ1GEx4Na3G6
VfBoLgHPqnMT5fCoa0jB+0najvvKLoiIpNo+144BVJ3hgvSanmx8XKAIFJVoUo8Y
pjR7eLG7LZQcjegl9F0lPmEzvouyHZQTAiPazGUojpWkaIW+YGtVSJ5hAPiCio+q
JCcmaDlRozeVursRWFcQ0slEzkqub1S47dl6TtOHDf0QLs2oRbuGo0irJwplqZaK
b1GxsI8DPp9btvaxZxzd6mNzfc+YJwKYHHgd5uvpWKW3ZHQrjc68aglCBsAPCV64
URnCyn0AcQ3s8aMMFCm/SzO8jNj1L7Z+u/dhfyknDt0zAuvFk8WlgnPlix1SN+be
`protect END_PROTECTED
