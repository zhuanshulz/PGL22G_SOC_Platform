`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LnuvuyE2ZBkGtmdAhM1sheDUZraslYaC7+NvgWj9lWAHck7FcqAEkW1z2omgW4Zj
TX6BzY95odHYw10Lrqo4qAj/1jIVcwZWAWhGt3JfPCqkHWOHZqI+rutHqJ25T42C
VLAVa5C4eXnzP2XkefuUxHWGZUXhqybYqw5Mo8dADIQrbqyXtvPESiFxPUmFJw4E
9Y6zSNmgI3dPl8suuNcOc235ArUqpqYLkK99yjMg26XOC+cCkDYWLRTfpU0A0p2o
6/4rSrFKKjlL6jGt4i/o6Ma3Uv7QxXMZrVhaEJgNRJVji4+Qde+DmchirQqzy/Oj
xoh1mYQX0YjHwtcadrskZvKSx3GepKQmm6zqlDRKQs08qd7zq+7dG4CgDe4v3H03
jJEbhDetLDrNHzHwnEbqZNgs5lsHwgMePKAOj+zC/mg5b8ir9ZHDZKUwi2d1TYdU
f+PprOAf6Lu30OKsjBttWFNHyEpk2mGdg13N2NKtwVdZzAeu/cckU6oA/bNUKowz
8O9qWxcpOAAUf1WjVKfxI+RNqfkA04ji114oYSIfKpB+MIkNIDsSBrqsD/tPhqCy
adfHK9eSs9f259Pm8qG12tlTEBYDdEsdPHaRpM9s9yHRhLj80XxBA2xFzGOQpGhO
Zpc2Gu9re9ZCiCuxm75x5nttxWJ9TDkwpLzDIfbiLTA7iwoXIPzWqQIOzIpRKlja
oCkoVHUOy9131HL/TgNom9+BpJZ93qem5c1KKiloxeNPXAmeCQtbzjuexB6IldAi
t7lRgx2ImVFeV0vePJGndCOh9hvcBbYjc+Cr+eESINuSn17qm7aHFHf19/lmCegg
ST3EnlEQ3p5dRUkyfA30XnfhsrS6syEf4/M8EyFwVi73rieJoI4xVBWSsOw1yZ0H
P8mOOwijsMlgN6RHAovJOIsy+QT7R4OiqWcO6+ZA7FkZR+iVx5aTre9FkzZuUoOk
RjO1q12kG1ObWT9zL84B8Rgw/ulDBUvnxVtYPsIQq2+R9wuSRJfta1JMbmQYOsyP
mGHAc9bsyQ8A1XqkRIbp4kCYEbzAsMVpRb1ER9IkVg3WBInJJ04sOOMdrnHkK6vo
c8a2SV8ury8IY+vW7jA6sq+lqeU5lL6Q9N8CZo1fCXdNj63s7tuQUavJrJ3m6c7i
pj0E5hnnCQn6qgQDvGUhZK18tA+vKPoefDPVrmrtJ4VLuxeh3HKsrPUKpV9Z5Zfj
aWlmJwjTO0lDIBtZa+88dicBzmy0ZsN0v4T4JQFWy1qsb5UjnkR8zM/xQ+HPY/L3
n404Zpa4k6/A1Ody6N78AhPI7tQDPT9MSY4z7PIROW5pHqnQZ+GvUNF/+J+QA54f
H03gCS8dbaJv38iYmSgkuKj9Rfk32yF3VVhC9iWyoX4pJyEwawwcVFqvENT+r/fU
f8S10vstM1xhySYIJdv8HNXEJMuh9QWRT4dRYYiezf90MSgxz0oqbIufZj/Yuvzm
RPSYzoTMpst/e0jinLm3Nio7RCwcLyNuniOcgxDvP5bh/NCKOHNmKjtTQnfvMeD+
Pp/yyFPCXqiiUXmne5x5RZnTJcbdcsSX5B/09EOx4bqWYfbzuNsvY5lzHM7aev4l
vAwYvDmOZQSyXo4pZBZRxBCzXX0viYVyZUsDbrifiv/uv76YpbjQNJBayAXQZmHT
pfR0/yPg808cyzjtNGPDG42bfjoRzfcYVkGWUUZ78p6Aso5VF8BHquoXtwNNiNqx
ye/XjhjoVX1nugO8tFntoWKetlNkXG8QIAw538TngmTHyCbqe1UnCoanyfZHDnqz
KbC9w/o4Q35w9J/xvyNeNw8DiO7hcpU81c9tcV4pzbXCkngxRwgHxKA8ehLATGpS
`protect END_PROTECTED
