`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FgseM+5w1NfOpE41hXlhd6zADMw3u026eZjhNYaqapFyyZBsIEIZI6BhUJM89LsH
3F88xjkURRq/GR5L9RTNSQfShTzaPnQroPeqE7xRgRmqgvoNzlAVNBBK2TUGCkAm
Rp9pKVEXublEx9gsXyw4tLBI9C44vIie51W2cczZ+sWqvYDi5vPYhTdFeZQTkmyO
5kUbDGGUFqrs+mFf7/nOym/u1pBpaATT4GTNxrWx/U2WafAaX/HtPc5LfdggFudL
WI2ycz+b0gTn2+ed4Vlutw==
`protect END_PROTECTED
