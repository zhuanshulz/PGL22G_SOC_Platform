`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iYTdCjBZfB7bYIC6Yyy7nrDOrjRqlI8l8W/gcaWsE2FjJcN3eYQ7aEEdmxXT21XR
TUJ37BzF3JIofjUF4mGE5nS9TeDAbUuh4TTyXhBLqttRvOYxqpsq1JQA9r7abUmT
41gKch2p6Fidn1SoF9kDTZyyziWjNGg/bTgNznAag45M8ylK3AJ/mSSJaZOZ0n1r
J4/rscOOwg6QQ9uoaI/NAd6vtyVieBr2wK13m0qVMnG9nGTEUFieCRhopmlI8AKe
gZsPvXyKRUU+y4Nd+OV7phWYjf1AWN5R7dOIeaqCFaH2P/oj2507BCZqk85W1kg1
Mn1JVFOfLgtRRNsU2UKtmq6197nQBkdNI+eWx7/4o46vNJErPbiAoPgh8uv1FtMC
ou/5h/bU+Znf2DHAG+d7AmH47EUXP8zU+1FZ+Al+u1RxC4trLQLNB8J4+y5oRgPC
wIXU8yK1DHAtm06l4+Arqg7usMipfq2BR3aS6mcYZjhtKpDY0bjWpiEeUphdCAVl
izmC7MP+10PRaXFoPKzIwDdY/EOGF0Ncvc/GtuvPGXYXuInCrkElDE4t3FVvU2tB
RYt+FLRaWRaaIRUhJHTzaRqylvVJXWziz4Kwd7qYaH125rlHSPxGMBNBTw/Rmq9s
cqk5z4JI1CM71EpGrfJ5SqrWAlV7JWAjHf2ekLzn/gLcYRL4xUXb71E/4QEJ5gt+
Icy/2Fzxp/MY0c19JoTpVdnW50wCBBs7bksUwGqFjWBgAuc7UtR4B6xfvFuAZNdF
+NiXmK807/5/ZsRPkLIATeEh55sRDNwUDnhHOHlVAw6cxmxNf2NyWTFpKDXr4oJh
EHXARXtHvBnG+/H3YHMm3HMJlKI5Pa8N3+BQGmrKiNEvqKzsTgxTeTgMZJfjRcLY
8iWaYjjZa+p1P7nwfbAlrNZaa3846QgD+1LxKFhu1K14mXEeiiYc7ILVKUIRiR+y
DtlrjugowvXBvzUR/AGbsOPEc5P9+tgVCFg7cRHxVa4zcQtylBFyPbqqY3zTMwzl
CfqJemkmB2g1uGO/Pu4OHA==
`protect END_PROTECTED
