`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vzLbbkYHTJHXWDCM7sLhOHO9KDugL7GQMmtqyt7NCA92++9rVl2v/tqQfuxux+OK
EJqi6TwZkqqxJvw5kRefvjckp8dTagRmGumhNSMeehT66PXOLCV0wZztDLTYZ7gf
xIuT6MXYR/9Q5DTqajOhMe7JoYQPkwQ6Qy+ZOu8sU7y4Q3PJsQgRQ9lOtQJWZ9AZ
f10sZgoN2MyXbKNJGcbxiQPn+OBdNM+8+qEEvNdKaKMa4+fBdnZmnFQHuTYjq2ZU
AZ7YEZ+xc7f89Qbjlvt3EeHEQkirZey2u+zMkuGP7HRshRc1TV94EY2bzHBcb+IJ
yWunU3pgMuYS7HRF6aFZErsAS9Rx5w0t1ki072SdL20aqAzReuZ+Wt1EXjOTRco4
kSu8Q9yzkVc3UdsOCdgW3kUqh2N9Ri0jNUUn5mSmnHUiU/PunCIlfeZRQHTFZi4z
3S5zMyP+vHexMdhgbF+fIIu49W1e0kNBbKWfjnCV/F9AhPvDXOAsxEdy0+JR6hHb
h1tNPP1IwGSOPn/QNAvEM/OCS56HykdaTBQxfja4AJX32YLGTL535w8bJELChiYM
EkQ3TATxtdwVUa3IjQettyYyi/8z5FZa/yoiFVExX7HdY8IB22tEdgQJp1fbIRx0
GkfFzU5/Jgu8hb0OGI1vfQ==
`protect END_PROTECTED
