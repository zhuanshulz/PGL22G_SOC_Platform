`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5PlfmYJaAAf2Qj+Y26bSek+E9uunTsLpyTjTe5MBtPL9v/sCt/tsxk9b4xQ3SMoo
XZ19iFZji1EEZlUT46obE+UwCTAqceSHRORbA2tx6H02MmHANC0FjbCi+U57fgPg
MX9bmu6la+8gfEIBLAS+2IoPsIdHkB6LKpdr+DpFJtCQcuWW2LrFPA5yDhRNonmZ
0CvU36ZtE/b3Nx2vQ/FUcq6xpwXe6dopYpD1EMUXQYvLJP+l8+0gykAzPKgm1wRi
9ElK5fMqUL31qZ0BQy0DbwdDNq/eDLBD9gJFzEBl8gm+78J6+aoZ9iU1VWJtq9KW
OpZhJI96r+TbSPsFmtKb6GXnK4BfZBPG4gePQauwx4+VOf+Vm8DLEoV4Q/x5l3Zd
QdNUutnj92TiX5s/Ci1UzLmQx1afbBYjW7kSAffElXqMXfMXcmd8j6vkXRzCcWWN
U6vIzxj6LdeQ3BlT7T2npjDQxbLEzAFL2ASVH+Ap2NJG9HAeEMMbU5e5CfyS4qMu
//ZSYuIaZ/xWjgoyAEpSkApTQ/vZ/jJ3DYDY9qvKWqZAK9OlMVHrfM7RIKxR9ePJ
3cWVu2zwPNIpnOElJ2vVpw==
`protect END_PROTECTED
