`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1DPa4RXmP5jYeqWXhta1Qrbwk6kvNFPXlRMN8VCLKNBFfWID1GDOCN9gEeMNiFKC
S1w63rbJb9p7xg6a2bcM16k1F9UPmnmjLoR/MMdoaTC46O2tL0dt8x3oBfeFfbeA
wregmjZACJDGc8/QPsPCF2PFzAmA2NtSW4KJS8+KwdLS2WnfZW2fYtS94TgBl/B3
mmuXCWpgCHo1qMoZG54ezGBHjnIMID3p1OSydH6Z1JcX7lk+c3ADolLtdpmXZl91
Id9l1jPAaZdYBblPdkag6stmCiMtPsr/66ZtPY5XL6SwPmKeZ1h8lZvPl5A+Ew5g
lpjE504ZjaPiEoledpLc1nWXVmhj2xn6YDTqMrMKi1T3p3qVl5mx/bTfOFW1CLBt
/QpntBzvcmOu7S2joiS8o/3CZ675Z29BnFusGbeMONeKnGG6oO4bmnMogA887X8y
c+hPYNQKoMYUkDdLSz71nxfnH3Isujiz5xCeNe+XM2BR0MVGQgVjUMU6Xbqf8D9f
00iKnLs2mE515wNG+53illHGOTFo+v1JHzdpWK8umSktyVPh5n6AWTUA4sgOkozi
FN+LVW5UfBEnNBcBOtHFoICajh8L5djJPsKDxVICv8RErEJk+wsRJWtH48D4DNcY
ayVKZcOg63Of4QDSJNDHmloA569wlcFGlz0/eYEb+iUr+Jfs6V5gIfYeqSD/4fDK
D8hRMK6N0mB6A0pGM0X95w==
`protect END_PROTECTED
