`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3NCTkmbYGNsp0zLLZwMvu6BQ+KGd3jR4Qmq0nnrSEGHRrtGqIRAEnuzqs09swZ4N
FZHKHa5rCdC+N/nnxiYcjdbXMN+mmgtH6TBPTWggZoYnrnSGGrJ+9Epww3/zYuZS
J1cSmYqC39QJ1W7VEBq25VFlyPakPfCHiY4EzbCWy5UVhu9hY76Pjk8S5J9ny7kM
jRPedFDgTC+KJmyGsjJ2VRQAN0T5heIcnF7QZCti2HFe6KyfBYTiSN5aIw7m3K7s
pKOhqWVTAv7I+isj1HCsk1hbuYbskoNNNkSqehz2a5ZQTxemJvWLChBh9ZDDZNUs
13gmwAd0RVRfvO/SvCFv3uS7D8UIp7+90hs9QjIHQegJN7Y4zsC5JCIh92d+N0pU
Um3uPKLA25fIqTOpMcQrK26WTaK0+u2Us7XfSal1sozC6IxlusHjw0ehmrLlfB9n
hioCzfTvcCrwC6w5bCtiYZrg09m8klRcNWiwB7/RTmlHHn+ncLYeH0+drjOsOM/q
o9KOgwwNvczUvWyor5rbVynov9hhQ/7ZXSUlMAs+UYSusbELkktIeNEds5AlcWOS
98Ib77uj8DI6mqN0c8pmgRMBp+cCbYnTLHqaXJH49BLLHyNuDcWxpc6p9JdmcxwS
5btbVvRH9mWk79ktdoaHv/Qo3OLfeLIF/bQYjwkJbp54OmML9imX8IvQqSk/4MSR
B76md1cwxlHE3wcYKi2K4UCTzmT/u529UUywn0xNoNmu3Qre1vysuh0W/EMfU6Gy
mLYJQQJTwCB6nZv3TT9bFJ0BrI0W9jJFyp7H//Jh6dTQQ48ejql+3M/GB2xBOhnF
do6ELt2NKrXdeKPpWJLpHMKfl4XtGFH7PHu0jvZPJ4+B3bufu3Ifg9slP6CIHKKF
Quz+US6rbL/ZTUnJSX2bxvbCZcpSX/hVkUjaLXc+H/wMDhOLtf+Zr8L1jb1GNCQU
IsJn0fah7ioqOq5zMxQ2yyAjd2AY6fZHGx6zx0HkoEaxdBvOOg9tH5ZWZQrT4r8h
9RTM16qbQ+BWtDC3emdJpWWJRzAde/k7d8NGDTXZl+z8S2JAdJKZl6zSLhO5A761
+2oHrTpaBbWSQvDVheJXvlKe755HnekHBos33wmsb0144nEllWZ8TUfSqRwGj9xh
RUJUc5Ak26em1za6SAqZcSp1a6ED1K51tWeHJbTe8ZoiR59Io8ilj2jak48lEyUH
LjMX04mcZyfex5WvTxR3YSa1M7e+yBDlo1pBPmO+3tfp8j+4yjJx6wjjj5alc2/x
iW7J00e+tG1diKB8qb77Qp6KZ48rGtYLIwvJQeUJK9kJkx7aKAGfK/DKmvnHrbpf
A/bohPAj+q7GTUQWJ0OU3Ewxyqmz02iR5kMP7IQxJagxBQ920x5ZoVX5+hMAJS+U
Mis5fOa4j01FJIqDKD+RkDcCIUwNoGJX081VntLaNpg+WFcZPhg1MGY1iuy7bRGd
ZF92C7H09k68MKyjJpPBfjGmJNpTqEqGnBun6i7JaJtQLv39KvBPM8NyUKwlu18g
jfROHxOt4pfggRVfPZ1+uLO/hEC691z23QuamPVsy1Q5GDQu2qUmv/WY/YGMiSLo
Aw71ltlErvfrSLx9/Fi1qnMW1OZb4masbRrnCeZR0+Rm/Pnqmb2IaDiaj+Tk89BH
kG39bpIB6X9EQGfQPIwWkJEk+MIRX+SNrv9UKVcCmpJIkGXd5QMfl04wztQeV+it
/hSZ8ZinLny0UA1dF2y1lUzwOMV15pHwlGfEFmN0Ffv/gTv+JSh4hqQGPuVr3hsO
XJcbdmo6yQs4uKwAF9BwD7ptCheLBRqK2YAkVm/ixtGOfo0saJgB56W3ufzJf0yy
DKneNxLUGpR5eJuAqeWj7RsCfwy6MN0W3tpLlf/wZsExzh40uJtVZH+TQYpw0/t2
Le/rLtNhZICEVP5x/yDC3aMY/vt6raYhQFgPPoXVMCtFyMLJsaNnv6JvRWyo7wra
NLsR5NnrritUp90GI/RWSmFGAF3dETZYz/9env7TLTlzNUZCPtt5FAwFA+bWudWd
4BaunXuP+UIMY4sJxFwJ7XfnbjUyA0bgI35LtYhPdPn4am4ph5l/PRdANl8AgPES
C+VTs0o+YqDQcY7bCmK6zfkTNXIZwVs4t/k+bwJpm3v27vRx9V/UrI0TkrzbTxFC
m5VUigfh6LFP9SFcbYqjFk/P+qSwHqVO00lNIsQSr5EwPe0mpsUIgkHelBHtGlSb
C7A8UK2afXESZf1qDC+ZWJ+L1lAWaelpG6MRXY9SC11Mt0YGk54Ei8mhDIPY3A5H
EfplOe8mYJHzvBSHBwAXq1+PL4w5yI8hIAOCTUBRuc0ZBdilHSToKYF+KaXluTjG
pBObAnUvPauXL1WssRR1+xazThp4V7aGmthm95uteZXJqkox2ggdFGUtEA3Rrxjd
aGfFZjpCbtzE4wddyGFviicY6Jo7fhuJnr0TH72MmK7u0UkbUO7Td1ASP7eKrANq
l0gz3bhh2/P/MIt+g+7O/o6WuCH97lNpvqiD6bu8yYaUNejed3GyPTDbIFI9t+Ej
e9RjQklRPc0Zkr/O1Sa7Epi1sXH37j9zTc56Zt8Mu9M1gTdDxPJl27ya2segHJBt
dttmDarCEiD5u3CqBISIsA2tGPhjYuA0cV/QMTco0mLhAen8fE9SlYuu8F0FUMw+
F9JfFJCAcF61IUJmUHYehESAexcQ9TEkHIS5eSV/RNKPgu6Bz444ura4esF6PT0w
TApF5lq9Htdx51Bx7ldfb+5hpu48PO8+29P/tQP6wMBS3K83tNkMjEoJruE5cky+
tJi35srQ0vqNi8DYI+xRiExmzSXAkQOMD+xhn+nA5faArR2t6N/Dd/EsyziQiBoi
qED7lI/4SOQGI1qWH1IB5MU656Qf8LGVoSiOvGhFhuen7hVsi//jsKtNfGb4r1UV
MAUHnOB3dcdds66Ijga09SfdC2Dcumz32EZNhYheZchJZSdW34Uu8/F6YaI/j6Kw
slkT9h6tTn4ekIuGANUrl6wIZEbxUn8gAdgseqnnstVWcoduMXMNcpD7fFQfaByw
AK4hAbfK8YWt0Uf1GLIuEI6x+5CTyYZoo87YCxA6vqmD4qT01oUpTyW1rJmf1A9Y
t8XHnOyaNyxg0Oq55RN5jfwF3f+Quc3GQzl4jLSCu+sCkKHI7gyCiaq7XsjPkjKn
Ao2BlapPhxDu9bowL4muQxwTojavzxb9bftoYKfNiBGoh5IkbanhwDFKrdUFAq2p
bkOxXiXhFe5LYGzH26IkxhsYmqB24hceceJAbs/KlHubKbXUHE4RTWzHWL/ffsW+
Fp8XE1hFO3SFDWXyYIGkcJMGUH+qMTxqg+yY8JbBvtRILY9QYlgQkS6q+Naqmc+y
BwNTiwu4siSLWvESyxoWQb0co2Rqo8eCaPhqNcTzMUY3lfVJqinTS0p4Hq8yHDl3
5X98A9WO0EjwRSJWsIXetk3jye4xSeOfcgp+VHA5TN3IYz8w9N8Ta3AFnBqCLHkW
pGEQQx8XPCjtIn4d++v9Xk9G/jXqD+wCTJ3M3MzWYJwvGyl5HX7dDwSjZnfdghxY
cbcfK2CqFRVvGGZWSCP713JKHJ+9qM7PwkjfhfyWGldHl+hwDk6WG4oayZRPwySc
XlxoVyNQTTgyQJx2Xj3EscF4289yI4WB7rsY5IVk+Id2z/U2frxX4GKsRe6YKLJk
J3L2nMronodufF2gAGeB7e0gE/ccJhYl+Z1+Z9laTOUFF+1n5AXvuC709nJJQc3e
ViRE9D7k3rtvNhDJDmSRJwJVLOT1WCaxwYuVq1gBipf0etFWBkpwq3DuB79noybd
rZy3zMAXwvO+lQ+gUqTXotO/oIWKKQ/3qQ7ZXD3xdP5z9yeI4NAjukdc0uCsEdLR
rbf8hksGnAFB2cOjmRceZM8vkrw0ncaavv0aYPTUc/vmN71Oigm+oJdr1wx7q69M
ZgFaXOVP1DbPOOheqztfKex/BznPpG/gkRD6MR0T3Iag8gvlWtzdBsYyyQHXYZZq
eGi6JQNYtph28AB2dd2WVUhlVEBoewYWGSdM4RqgA07YK/4qSU11HIEdC+3cx169
UbKis6r2kjPK1d98uxyVKvFxDfvf/sfTxQog9dbY18kO21QrBdCAyVyzCxv5/TTR
rnHRt0SxVrOKGEkFxyYzqG7giXyn1aDNu6YARCpWYRJg7Ct0LwuUxPAD/QkYWQwc
W7I35KE19DQVmuv1iFKWf59thb/SxeN5MVx12OMaI3zxQceyPwJjdWl4zBPTQciJ
VffdxltYX2alMZ1rc0pFOtVD43uir9e18WO5ri/EbMYdSUMC8H/wcIX+Kgsf1APM
C9JKQUJ4DldsOyMhQvTS2ovY5VWG87qnRboj7wIFeW7du1X9BKFVlTojKYjW1xxc
jMwvG2IvH7W5RWuv8A6rpnClNuOrxvWJgA4oPcNfWlsqzdN9tru28ScGV4WWrJUF
mj7sO2Xv5XSCv0iJkitojcU5N/Lk98L4dfIheRAVA9xhSovL3rIJ02zHK9DZMg8u
QOo4G/y01B41KF4KW3/OUrjHO95wG3yvCx8awVATxwFkuPbLvZytNPmn2KAuK6QQ
/SJSq7DZS6LXSNeHuKlzm55svkUUwWnO8M5eOCdJ1b9ad4QWFliimlwuk4j0QP76
qH4pY/owXiXyT8XH3p/L/3hvlW2/uv0tyF9hcrXoJjCKyqGif0tyQpo2DIq11FJ1
QNWp7PvFj1vuAkkgyJdAX941/Wr6IDP4ZYx8O7OQ6O6Oc1vbP4sYqQu9GIbQ24U3
l8woya34/r0x/c3JWTqnZcn2Q307yPyWc/CjnZ36Kz0i7bEnQ6OylGHS0SQJ6EQ9
j6EyJW1Xu/BzwaGeWfg4lkxCwYLJts8XgxPZkqRl//OaBToklcIW4+95XrdC/bZx
RbDFnIrI7ubWPFx8d/CWYkeD8PY7JWCRBVKS6Cw/DGUTNKZCmYF79HHDNvNvkmZI
DSoh/uBPntj6W/Ab83enn+Yul/hgev1/AX4D6zwVUbzZjEUA10chnr35Jy48IbM/
`protect END_PROTECTED
