`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v9fKBa2/VGh41ngIZwtg3IfUC/wjjOQGzzLK0u15QxZJeOzFrA03pLtl/A7t+LVx
qg1OXTMhlty8CTj3jFWBRyELc66rA04BhsvQ+ZbDd3StoFRdysuE8NE/jDNo/Pka
CJLE/6wrBsvLUYg4UTINbTeGiea6CQ2hl0tHFCSaXkE3c7gRRjGMDZlb58AbrRBd
uUdHMpidUFs9FasPGoIy/YJPTfM8Cldb9SdIuh5tdrvjxbo8Jduy3vaT1OinzLno
J1VC4PYfS1aDXpOceR47J8lbvMW13mjeBUAFohQrByFEYenpRXYEBCxRa68EcQFg
YWA+kuxyaYloDzs+WByboZ291XVZngRFwqkFEzoD6BcU82FNxQRMh7/e8CpzlqDi
6zpFUHovBaah/AddXQzg+fl8ZzP6XMlCdnbdlUNOWdEURPrSKUvSAUjCxXFZMLXy
cbiyFIdj6VPJUmbmCbzyUXgZEXDfIJRedBHPzFdsKiQzKtMMaDx3COzJOU+D0x2N
0XyC7ko9b+BHi7y3qRNiS7VdVtAIV7lBsv837RazaOSI3GZdYlZdcoTJSXyVn2L/
yxb6Q2lOi91mZ9b3WBBZbCQpyHBlNyQA7XTjKvowZIrtxsGr8/8EJbEiI83lRdUd
k1XojgDLTQgosbIvHblB8o6d1l0JTlV2DuPOz0z0BJGZDW0CBgNi5de4YJ2rJ1bd
FMUNuXMqZMxDPS5pph3UkU2ei4ZcGchTHmB2gBG/0/aNT97HqRCwlKilGb9zA9rC
nl5qBqI/7Pw4fjQ+A245jhSXOdYkn87mjSbdvFD6rFCIlJMY1OGYSZubgkrJbAKF
2IV61F19/hwEO1hqTisFYIA1XV4Tc2+ZT5zG4AzIOIyTu6o8uIZbWb4nRyWybzLL
XQTljqQYfzaht/S+4rGBiKm3uzs0wDuW+KVeKN2YUfblRWOa1hQ0SUu1J5Pq3GRl
WGLyjJfvUESTUiOuRiBA7hDlbXKze0kpQyYYujX28+5KTJdLTMgpbGVycKZswgOe
YbleIw1RODgGS1CuGT5bbIuFmUsY+Y1OGg5kKqc1iWutwuLXq4liHmNVRDsRgJiq
Y8DPTz+Kv+QXcQloOxekKGTXC79YVDvpxPBAENwKxwkbq06Mf3pxAPlkB1pwY07/
BRSahY6YsadqPOF1KUpSMWQYCmMosW2wsPOCwdkICRPC4DzDsFMKlrPann9LVb58
7ECm/oUqS8bKVolUlvkTiICGUU3KvyDaMrE/xlTxyQJ2VX9fxYmks4h9/QC/2gwp
sh+1MCITk+PyS2iAmkCwWcVHzR9B5qm1Djwqvd8ZZIvWE/YEd6tzeH0SRTmZzIrn
Dn2/YeCTv7/Uip3mqx8ywXiZexIPgN9HRY+2bcseKQfeqpTwmuXeVPf+cxINaXMu
CV8E1Pxpwt1qY5taesxaRJj8ApT3GVTAQSxHy8dfeybounZCsM8x2CL+BzKr8aOJ
oqqnJ06RSo1kmJ9b3zWJtzYJ7mjKfQdYO8BUtRpiBeFVl8ADEIGZSOzbQspqFf7K
q0PulhbuU9JEPLeYYYMY7DaUY28i7o+8Hr5WQPiPO5dkHQLj7bbWdOzcuS/XqqFs
+LNanOm8ucLr48OLCWNz7TW09yPNQkECcTi0bEJJmEB07aMhAzX6NqnNOTakouwJ
JY6to63g3szITHGmSQgAL63kJ/DMYdIX4KUzShbl/7/p4yH9tOgONkJZaAagkeIH
PCOkrX034A2FbmFU1GtsShLhrryls3Mw0qgKP3W8MJvZ/6r2XneT1XABLRrV7bLr
KOTmz/bqh2Y66iA7KlbdgiqAXoVeEq6W6A7vQ+rvkgWhrlI/9hsBcpiCPaW6OVCT
gcE+CXrCaNb79lZoRiJHnIE/PZQ82VHR4mkQcpTMLEWkLfsLdmpA/vdYTkpTuH3K
rjICqfnVckH7gzaPwZssW5hh9PZf2a25yWOIwjRKKOO5PIxAjDOonwdqhtYkZ5+3
qGhoFtEyrSQrZYTUOe70ZSfPOkIdWNniiY+9IZmiiR64xxKgTVYMrpIZ5adghYj0
65cxeAUBT6RllvmeLLXO0M47UGXejlQg+nXcjsA9lcyJcSw1E7fAFZwj8F2QQnHk
7OXDlDNJKJy6VvYFfHKUrWKPaxxrj+t0VgKMwzvOHIfz0+n/UZKG1dpqWWE7enwq
Bmlu56gf6/AhLdVjVNTDdlXiRPGdCogkeLD0U2ZBFaWI11BT8NzB43HfJzvDy7Wf
GVmlf2o8xUgRaLj/Kvckou0x6aMlF5Rk0n75MEMW8ZrC9s9EwzCYOQw1IGzhi4go
17SxSxJfnHwQopnRVuGD9lsoWhnxQn6L6iJuxxM9U4qhHW40GTDgmwWPkT4Z8lwX
6kOrRbw9KPbYNW/jOzEqUUZmDEGjD0gIgZbV2EkizOT8PQrINp9cPHp4JlhJ+ZUF
DFzySMv+oVptNhcEmpEekMsvebNgd24S0ewH7UcqM7jYmwerUptMhickzBquwWoi
X+bkWY03Vhfb2vY0IBM3QRrI0atXVR39WUcatITZ9mtPurhKc/BYbkSAo4cGA5cb
jgeGsg2D+7aAUA+e9ibP/wtiQc1QC3wU8OKLU10/oE9RmjtqJgGWnDR+9QEfYN5V
8OLqPovn+EP4lcDwXHFWUKukS6bGXrpzseMtylYIIp4bvUG2VZE0hwMksXJbpB7Z
85FTYWDO9p54G+87xFMy2zkRbJBDdzdyVZdUhrcDz6AOamkRZFCzqU9xoXRRiQyh
IzrBZM8SJx+ccjqdKnpEixYgFWayBEo8mXinOak4P6g7G6z1WmTxH7RC/Et2Rzzb
cnosLotaC8KjDVv44T3oCth3NwJiEmFU08EZ4nPfSoMI2KshYzx1s94cy4e1CeJ0
aNVNG2OMytXn8zXySeBWDfkoAb6mxyKL93ML2WsgRLIu272Z51+BKHJawE1QzXAB
kCk7T9rz0d7JRR5SxKM2YhgTjo1tVH5fVHSKsQ1Hf8UGauJw/KXpf3yOHuBK942J
ckToh8m3/tWyuRVfCF8G9sYot4qUV0pd+Tb/gW9BqU5kx0uxo6a5iihLfBL30tuy
rwpbXV4iadIrVBbLvyW2g7nQCCeYnb8ISgmdAKDtXKQlrzBwwArD3pqDuB4w4+im
Veh/bCKk83k8bnzC77irk0g7VL+L8eDHE3NCJLeBZ4uDl5N8fywYQTj2vQ4wyjsu
NsqiNOZ4bI5aw8Gi6sE0WvbJ0EJGyJlif6k+MCFO9CZO/74EoZ7wtbWbKuyBkeTR
Y9Xpmrm4XkqQgIJAlybhESjyo+5umREiEZ5zwLIwB2vk0Qt5qAn1kojqnG8af7j3
G8wmhxmtazAKaeV35dsbBzvEALDbyqw9xukK4eikGNxLXMj6LQS5F+BXpjXdhiU8
0RQZvzmjUEpVbl4ZtT5u1RrKkxoLQg2y+fjCTFNjbJTG5NqErE31Pjh5ozmhyIoG
NoRHacPmwL0ZT0rU1etLck5VLg/zKZ8masmYIqAyfwAU6myrZFM9JKaCGcESyKNg
D4mGf+6lVq5UAvEIU6gTSg==
`protect END_PROTECTED
