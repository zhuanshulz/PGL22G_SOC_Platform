`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JHw+71umpTkm3JV04ZwsD4p5cFtipYljayLwHeiBWb2MxvPULEJQ7qKxfzYT/DdB
aEYnGVqmQwOc2GhUK8Cc406+syaUzz5cvAV50tC2fL5z+U5N9jyr8C43/2QVExFf
ldQkvXLaVBAQIvLlXKqmFrywkFixzhDoEFMpq6WZNgKe8rkf3BuOJ573+uOBR0Ji
mFXFdq52o0OUgWyIUHBU1q2oBrAgyESne3RPSoM2GaGBxN59HrxKmiNaQ9i8QRr3
ZtHB9RdVfv3bm99zTedS7fUpOWfUKjuieTIPjgxjc1mKLExcxgIiH3/cUg4vGbyI
zWdibJmPJjOoXatPvikiuAqLzthD54D89dE8bMIiJ3cZbFtdnwaARatX7hrAMvOD
nJaUlb7/z2VkoE9qZ9JX/zyIJdaV6PQxkABH/f5d3xioiBxFkm/20j5z6qVMZOkR
EmD5E/iLWQ+IrJVfFemT9JiAtip1SKQ2E0uHuevzBF4jrKGyB2XdTE+HOC2pTKs3
EGpcqU4h4C0WZXSc1PpFiKn9UaDMOvznSHl9YdNYgSReAfgaxx+PUCzwMqtiztAa
NarCiwiDL6svsGbmkqkTt2FI+zj8HMtWncXiy5LT/aNuWgYfCtpC7U7BF38YMSCP
FOE1sCxapnP7Al7q1BXFyepxlkEuLOWKKJdOF+3YarNk+Qgu7QXOQvZUL99H2/1a
rHg6NYVTTWrpc5cP+Hp1qGjbe/N0QEYoRxp0OPr8K8wUoYp89Ek/jXlLI7WtwK2r
qYvj8R80lmX1Rh9yb7dC3gT29weZvLmpZVT37ITIguzCbMP9pj9kmUHX4M/4iGPD
UG4bOiFpa+ZPKwoljdJprtZ4JQb49GbCi7lRoc8qUVYmivVtYsgc/fdrp3XMlxx6
`protect END_PROTECTED
