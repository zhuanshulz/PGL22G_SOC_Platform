`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AsrVhJNLlccTJLeRrMCwwM66E74LTO6jXPX8WBA2Q9f4ebo/FkJvWaZjMLxM4C0f
WTaZ0nr4Xk5wX960wCIj+AH4KG8BIhy8lO2+nESctqDE8/CKEEeLWyaFCi6OOjUz
vgvh2StqdV2bTOs0mqoNh26bXzwJbVPwfMtuPvA5TAWgWMT/NtOI/ofprVFHd8S1
aGkzTQYQDhlp77n4JGDhlN8/J+4ZDS/w4OkwWglbrxGlXoemOdUfKqf/KZAGE+dZ
z5Z1Bsj+331UuSef0x23ZhaD0Thav2R3v0c6gC5HY48862ntqbd+rEeFGcTqfKc7
bqZhWNdALLd2chpjghEkbHf/j2zywwzrcdZ1AidbsFZweoj1occP+J+lxW2j/qPv
7xwuqgPlUxa9HNu8bu1ad5pbOXrvC0w06jE0lpZ8SKe06f4rdKkf7/GvNKYlL+2r
u7ErtCmDZVO575XwY/5RQm7m0sg3BQb4iQ9x2chftwj7ezrrJHF5K4414C3L7fM6
NRovvP4ktvmCjjvkxhR7WdHdgirGHF3kdC/txrSlOgZZ+gdhuXRNqbwz1vi33oSj
O1Nb9ZKHx3K/CUYsWHDwf2RO9l0JHD5Pzl4C9sKLiZH/0/fipNC9+uvxsyawsHfw
+A55WklnEuK/sncJQEsfJS9nYzagqTrHCeg8P6DKKCYdc5MkQLFWBBwFwcuExOcQ
zr1vNnmpPr2Ah4zVlDne85txlVqTMT3kgV32rqdcyk6apafvlsDFefYUcmSnkv8T
XNtyJSnGwZAr0xxxGhvC/03DdC3QifKIl7VFEx4DRf1MnoMPqSsuLMtu2sZRR2vS
p66JpfwZDP+cvgEvn2qRW3n7aOBg6V0kyCStNAYc2+uMCYqE3tX+wIfY/eL/xqWm
vaLRWmjVdbADqevjXn4beGt/sure3BbYsvPGdesyfYqyvguIhnBh79n6/cMFb9Mh
Qe6Q8K8BQbJVtn5AWn2kjaD+vdTqdjAThFnNvOE3kegTBzDStI/t22Nc8g2wjnuS
cK8oGO7V7jGleIBPvNZjJYDSZ62idk3hRVlR+Q02JxPAa/xchaq84K8v+r7kSBV+
OAT7HeEWZOqH1VfgriX251Kf+ShUIWC8GMrx7EGIiNJkK/L1E/mFLZPAvmLe6LMJ
rtOY1WZ1QA2DxblBOKXQIg8BiIXZvg1vZPw9SPa6j/xwyz1DJxaX3/AogweR4J7i
ycyxq9gk5Suia5aw5tNyUGvC7J6tiyzSCWdc5MdggVndKfKTHVUARMovYRg6EUUK
x5GMBedpZZJpk77ZRvwZoGbsTXEUuadqxWl9O+2Piz88H2DjBKW7VABcyR034X4l
qMy71T7fxz+lfMbxfvB7Vxph0B23S5Q9SX5BcN4ZnzzRPEB1zQX3kXZgk+1lIYfa
KbNcToMGKr7vbQ64Evo9GAjoDAwK3MGVOxdlua7wd2eA4N8GTbpRA7EfdhRhrtBw
aYbil4+A5Ka43xAE8+0qen0AYNH1etAy5trf647R9fWzkLHK/WyadK7PD6tXOtsJ
kZubxeAsU4dOn8g2F3GU8GVNPnFZtunAnbTqRRUSDgvfrVFoO/ZtjjVY8tmm/dVs
CLaCy30MOnl0Ssqe+DEWEQDyTrWJ7tnxeOF/CW8ezDsTKNbRDdoCdSvH+tckEG05
5Ko9nKrEViQS4j5tGrOjYNtDX/iaYTuYZbLrR9aff9rUc3bf3tiIsH/7TuUZ3g7b
eullBNOvZISirN80ZPuk2dRiONKu0m0pwdXHS64z9EeRdeMDHoykyG/aChbtA00D
EyQTovEXnSwE1kGCMsUv/PxGuBBuYZ2OiHUHiZSkXgpSuwKiLgHIYYcahrdIccB/
TfkYkQGmNtWEbdTnTY7dywzHtufdRTa7w354c85UmUyPEBNQcNjusi5kGc3r1JGS
c9FmFdDJnIvKtV1MO5qwjJbAlLbbQpnguYVsP/wONdkeDbnndTLGp1033c6fSgLB
V3mixclhi8BhqHDY5GW6r/24PVfXIhiwIJqCXEA9LBtib16Sujb1u4eitopAcLbb
whlAj9g8ea2gZhOHNGXalmn7uhfRgrpiaxI0uC+Zb1uN4DL8/An1y9uc79enforx
NFDwMId5EjvIg9ae/CZ+0PaWpkE+rXmK0dSaO1V8SvuyvgnBPXUObiuXGhEzghBF
3Vdo62vv9X9D8S8nZGzjmw0EohIPfu3fAzysORDZ9tthKd7Of9eTt8UoPJY0xx9o
Wq+3BmbV8rh3P9sV1WpdrnM6JEDbGmdy85WfiYyuhIGdDp7ZGdfvsVb4A/iIICC+
5+lsErKLhE7HcD+21y8s7oAGTBCIlUECxfG0k2+rN9hj500Y61AjDAljbcNdk3yQ
wEtvraIVcb1LlsY2nkN8VnmCzJc5ybWLUz0Lqkkl97IbJ7Oesy6ezchpdtjXaCYz
WYkId9E6u0f/fcDCOWzl6D3fQOG8auSg4Y6KgEAzDNFG34CYlnrzISaxp5cpRBxx
891dSOMKxiRIIb6oNhCUDJR5VN0BSMvNf1gpS7RItAMeO2icq7i5ISu9+J7D5Nec
GGGWNL70R4dBT8c4A8YIxp2vOZYEEfz//HpQPZBCYI+RTlcYEjmiL25keRvKiXvk
wXoP8NjATUrTWU9NyMGfrFn1iHv9sdm2664P6nTgULqtJ2DOxUSs5mSYsl88CMXA
0Nhpa53rZXAj68d+kutfRit1MXS3qg+tlZvID9qm0YoIofN37MBzq0SfQpCRXik8
BUAtQqd0uDxbAlzrPcTGhlEMO1X1dpWaxOCrSatHHZpBEPWjmBs+geQe4CDWAYeF
WI+OdwZHwXQijUAAPm+Kqaosgks2lEPTTYINRxPfXSlxCdb7oZC/SHSkNsBJ2uIm
z8lGyXEbrloys0RGwBGMACQBc1IJXcghtH0lUd0M1J43OXCeLzX/Kt9Dq9Jb+ptM
0Myat/qhB4Xm++aP1GOjVxafXzv+FeKWy41SIznccdkJacTp1CgGJ02lhPOxU6si
xLBX3Z5TKBRYprx4NW3PEV+DrXuUxdf5DcU3S6HM83T897vhVIddcCdFzdLx4ZNY
niMDP2DTsG1EScHAgbk/cFYEkRE+Cc58nxUtBHIu4FcGQlphtayPGt9fHmNcW1ep
ZIiXEDwgIS0kS+OS0TuBzQ1bEabN+jY4OxKryqzqXf15wQ8Q99eaLBYHGyX8RsIy
uiPfGV2i8IYfX0GYdtLY9j0YoXAEj+IuAjv/1i73+mYgBeWPYs6jTrr3XH2nk0Id
sf1aMKug3ktSbM2F/mNRABAstw7MGCuqsJtgI0AvAN+qk/PZ4fuqpZ0ln6tw9flp
jem5WtmX10e2nNcMGcYyzWakAUwuKtgt1cA1Z6BlFgi5tOuhSikubXP6f4RqXKVv
flGwN5TlrnANgUFWOX3QyqYPIjCA3KwDMLg+eSydiKtqZ8qRoGiGi7MESdMijSoQ
zio3yb51Rp4qFo+FUlwqj3uk++Mk6/FG/LNvQ83Ez+wAnuaGe/4b57QfqEuk5Ku1
HycKzpYZF9QG9R5SGE4E8za6DcfT9ozdxX34eqJdoeHa7ubh6LbZK57K5F+Tc49F
OTAwRUXCE2/Bws1abDgbZIysHsDfP/eiA1OVKWCz2rynzzNYUA/st6GqQ1SFSbP5
EG+WmDQziga8WeaNxAckhDvGN9yCd8G7KuFxg1CUsQaVZlP/Soxk6Jj+fxIMzFpU
YSZfRVip4DwIkzJuyLDC6FzLIkTeaI7rtdYbaKJz1QQtwNs3sDwspDNAkaKo84G3
YcQ7mIYSPbciw5l0HmnTRDZh0Mjo6jN5TDX5VUButlSj8/V/Nbfe5FSDlHCp3rm5
zJWXFEjFB+Guoe1fDSs59JNG3tEzVBbLFfy8PO3BcsX+um9tJoxFpGzoZTDXG7rL
1tDwnaJGslMQpK0qV1JNGfajn6I/C+v+aTWbtupqeWu0bfMByEFYPP7TKiv/Ove0
1vh0YUFJMqpW3hDeBtcuAKRQwnqGc6XDdotXByWRPxyzNogaKV0KErB4l/lbHWhZ
riNYJ0E6Zp47ubglBdUbd8cZQDy6rQ25q9hWO4PilOGvVFsKeDXEBGgj7rwSEr+7
qUfgV3xHPZi8Fd6kR0zR0GXeKlp6y/CiArSANs+77CEVI+wr7a/j3koSTBeiO/8F
p8vkJ5BCKM/mDLPto8rLQo9sAWJed2Jyo5orf2RELpDWpIQsgUvMyurYm5WmJ+fb
0aIeRnBFoOqbBJnvGQT3WRMX0VtWsNh1EqzR89uaku5vcOQ2dr67SeBdDod7NfqY
MiPmnPSvUlN+8XDMdnhtlG6aAt5cft+we0jKKHjJefGoOIAALFC9/v5hrcLF0Gq/
bajOIRgeFXymFLM7Ld5l5u5tToRMdRl3mtZO47Q1Udt4dpy9eHnukOYUKZv1hlAq
Fuc09egwkNvafOD3kdVJSAmCrtoQLK4yQ5qoOn5ymmjh51e5/5fbQRHD6ELWl2vw
yGI7fMQgpk+xZNHCjABfPDalpTPcczEa485GNFLf3CdXPk7N1jvAnFH9GNXyHEub
zCzRM5L5qIx2t6hV/2LYFViHxY3uzDgM3A6x/x3ufJZ/3bNW8y4tbjDxVFTrIVse
zNEKnnwuMKdkdcraR/a0n73ozo3gwEGWrFUNaBdsryPXXF5Zq/oO96hPdbRv+OVe
yLODVvappDUXeZfN34mbB4Jbv8xEMrKHNiT3GO0XDktTyd8kWXwOE/xSf2oAvvxg
3P9e2KrKcHL2EkBhyZzBIsBHwBcDcQ8+EINyKoRbKpsjFfGfIW7yofiz0nuYq8xb
A7fFrgVLCCHh1YpntLDTrEWNgnaCS1tuAICnpcI26+MQ7Y1j02Fh1XMSsrz6cNKk
hzXKb+gkHBeR8/NRyLmbQtu32LdelFtZVR0ngxPYNi3sX883subW54FjjeMQRzBA
mZdUhD9q316+dPIpGo0ivdFKUI+5iyuh1/lCxVuM+1yLSG8eRbBVUJttsoOHIckP
vQdbo3MQNYzEhBJJ43ut2YGZCPZWaMBd4C1H8LfaF6ZVJcZCw+OZsW4VTEP4RBko
dwdcKHLxKlBb+zsO7qUTmo0YKl1pMMK9vo9Jtd7ljlGolExdZYqC0dTZpX7MuR8P
4VWqBL6KGYB+6WJC5G3VSRuvSe9yMCKFVu/KTT+AfJDbYs6riVstPBxEgSTfHKLL
g+V/FX7nkSSm6nDUgcX0ELomQiGGvEbesYTDlfYq6i7QaAtnL+/aub8CPDJKC62k
SGhkOsheakvWZRVcu+201JS9Uic0B9nfvR/MZdPqpH+JYjg5drxQQoOXH7n/o9WU
llNBHi3PwqVrCBXji6BmJ8c8KRw0N2bXiFD+WqcMy1kEf/yZc4X8IIUSfHuvCmf9
zZA1BmfPUEB7CqC1RB+ztDkNKMwqAwVUdsQh8blA1apkMjnUhh+jesTD806tXq8Z
FsWZ6soC1zGbb1/kfR0xWnPlrVKufemPnfkETgm1PsN7o52F4zt0M0oXT9oOvcXR
3z4TVU9nYJJjbo5CQYg9X2bc687MZnm3u6HuKNncaaF5FfsBr9E6ExnDfgAWPCJQ
Pv1rKNe15HVUWxJzTsqbqYPp9Q9Iu3vSjfnpAbnz+twjeqNA9kuWKfaXaL7c1Z4c
vHU/SAVZcNYUCyqWSjSZK9ef/7dha/aYknfX2tFa4wEiWQIvaGme7x6nbMdui7sd
oSlFrP49dumVCcN10aXR0Vf4cawLERpwh2J9jtzaJ86a5EUpi9ZfPqFglW1aEZaE
/tl7k7yLCiCD3RaFqcbLJBAqBWXIulpJrl1uoRR2VIG4Wh065JIPU3G+fa4oklfX
rho8U7Wc5WNpzia0bA1Fz5lickORv8mmNf3xEYndCgf4Ouo2+lFLSce3WlrAHA7W
XLCFs9aq9LlckmZLz0wUl1hN8M8JT0vVQDiYQOOYAXGkHrFTggGaKAYpSXocGM0N
HoQuHjRQSFS0TaziuB4TG540SEJAg9mnEZ9W5W3DfaA5Md29HAARfr5XJn1uKJxk
82q4KugHOrS8x1/FYHGNihmcCNPEHyQXN77LF99DPwoxW5NXfUYpcl1jnPggAVhk
PNNunmp+9yYOdFtegrv8NLGNbC9VKDru1mzn6/QCIxGEs3Q389t+VLDNO+9Ee1tk
rEWjhv4ougScyWaprfYHYllhdJZ9xbZ2eep77HN7xn/g56kD/8sN1bA6UuMGXkw3
6f0lT4j83QHZB2eW98FiZmQh3Q1/FA55KyxouGXQf+CxQz2GubMHRTJrwx4oRLhq
RJXGdkvtCxIqIZALyhxWf7ZUVzqj4ueQVajWJl9umL757tVzRO9KiprJItGEFE58
hxOtL+w9C7VUMPPjx7J+RYGL3AeerwlhVNo658Ob0HrqLOLpmbnfmMEIlT9Slw7X
UreG4k2OuFMA9/U1n7n0Zhs4br3oDvcIA2p1hNrGUIv7Y2a/egGNvhT/AEz3lrOi
xZUZWV8XVCfUhdGOoLicSrtdNtZnnydkytMfXsAfAQfrk9/VQZk9+9I37/ZEA/ba
Vh/P+DoKaH7sL6D6lp08gPUjz4B023QlFVyXTVQAKuokIZGq6Q0UqlzVqlZZg/cL
e3hrC7/DrJ+TKG8NoGSVT2m7GZ+6J3guz3ukOeLo4lH232QbJkocOSYj6rxynOb1
BV4VPatEwwUMTkH/iWbGxFA2H/odpLUkle11YveIzW42oZcjZvJGndA/7YGx04hw
TMaMSz6USok9B9+kAJONOgzOpSWwsB2kCveu2cVF8mcHhzKWFovsCBjrr2fRUezb
PN/nBkwHCcJ9mpOF/RKPm/mqQaulqcrz+r9qzh/YLaN1NLuHYttR2FhmYoP86+iv
Y0tdWSZCLHiWmQbQVkQXYk2ihfuh8wLbNRvifmbfAZh7hK2dUTCo5O9JkU5TXxGx
5CRs9xyMBNaPe6+VHfQ+baBTIdxBosngefRHQdn78q9QCmycX0tvza/AOI9FlRxV
+s/zZWWjUCkJijOilCkvaFCC4ZRfZD8onWneWgPqOahbo0x+2qhqfLWJzc3K0rv7
oNvRGv1QDvcqVHc54lajnLHrXUwqhe7MLdxNmpIeTVt6caJQb6dVUo4bxnulKLwQ
OZviC0PHtiOEwyGSkVXBHjJXi5TTC4A5VuNZvxprGAzgqJQdJpRS70BssTmPwGBF
+QEa2dEhMVS2oX1ldJGVUaoFfgsdAJbWakbtAlZEwzZdVEDaXzNH7N7e7Pj1iIdD
ynGmiX2E1w2VHPBREDMiUCA3hgYKZ1hVhwZytUvcl9gc56BKKqGB9K5UaoRTSB3S
jQYJIRfV7TwasZjgKtwN42d5Ohlq83PpNh9exXPNleokkh0t1+aw9oL29PuHg1PX
F573xaPAf3Z0A+2WXwaHdGv+zKm5D0YeciHlVAVe/iamZvngKMHvsowtPj9QRTbt
X4x/gytErp6ieOm/UM5BfkpcQjjSbH81+i3Ma8wqLVRssQNgF5fIoTcZzR1Ap/fo
WOle3aaKqKOzrl8vTXVOBGvnaQ6g9D7epfMnHh9laaZlTsQLlNCwBZbpSZzToJzC
DqawPvjejxBoC17yM3C/HQbRHi6I2KCQn4mGilomh5+gY95wR7TSmk7PZ3FwI2Jo
ldGOlQD5Zbzg3jHZQrOrlOvMMjtui4F8eCxNONWeHUSEHi4ou9kvUwkLjELbtNzp
JyJ/iHRzxBAPKf+9/rCF9CtNOfth1xZyBu3i4c1eJLuoPZ7/t5AU0IV/mhuXllRU
OJsJwJJZHXf30CtUj7iJmjDj98JK4cpkT8T6HFx2pnA=
`protect END_PROTECTED
