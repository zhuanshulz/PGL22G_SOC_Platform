`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9HftP5MesHbHc88nhW7lL0wg49H4JSgDpzG/vkP4k1j5VyreBRh+JGG8hPlI0BwA
xXKHHzvGnOAA+4umfXUY6/juYS0M2BRdZxax+ulwxoGkxUprqavCByyaliMqiOxb
GEF4hPM26ead3FrGYEWsTyz+bsaGO/heApdArSuqoM+prUD9N5wq1hXdIS1UPExN
7nREbNW62q1V1lb8TUcueg1/+oBpJuEQOtUdo7OZJmz8+c8Ij2EYRcKSQaHLwffU
5qz1m3/Z3p1AK3kssyCFTeUxuBNRTS1O1bKP4Ajk+G2sUBXrZWXFbXtOLqBXh2GB
m0RpZHSJcgQIAFWsLI5U6Q==
`protect END_PROTECTED
