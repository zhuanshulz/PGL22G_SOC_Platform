`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IE8jsjQ6OU2vLYL9i63y0VWTD3m4AzTPPJxwyCIjocAOY3tNAFPzXZHwJ81KCgE0
r+Pde1I8UNeFjYRlnU6/+7cqpLq6YRQylUinYuuwG+Qs/uhsxcAAcSTccWFHwaVG
pewqMjvxbhS6lIEoQ+t2lKHdlSh6CZF5wOjmnnFPIUAIxA6a4vfKJ3kVHWsZyP29
j3dHycrPB8bkmNi1KtFOohmWA/MMFwkPUZpya0t/TLwYR+V5N8rBthNHsIv8K13u
MEzmfV1QUzIZWgGHp7p95R3vPLU0xl0lKegbrPx37eNbeHl6Yfalh/4A5jKm/2+M
kX+i7gJAHRU/06ItZteqhBFBPIu7GHDOn1TsyMuCfVgfSa7J14U2Q7VM1K4RN1wq
mUyp5S2z9PAqOL59sYk6ygFfVNcSOvT7I3Y7SEGBsmfFPt4j6GoHvzX2Bu1pi2m+
/Q7IrtAff23yW8FpcqaTetKIkDBdW1ViLK1740uLG4AbWKjNZ+oQeQH2Tmx6OJdT
xgDkgGqrtr0uj29w9BQbWBpq36OwRXS8yBWYGJbjWijtinUGyD5p5W/Qx56p7v4q
9pDdb14HC1XZC+kPxHfr2SnuVsn8K+gUXlH+B1upkQAc7fX2SeaUFWsPyBiSbvFy
LJHWNuoB1JcIpTJcKb+sNutc9UR1yCSMjhwSPUddwlV9+W5+iOLNW+qOxagSj3Z/
`protect END_PROTECTED
