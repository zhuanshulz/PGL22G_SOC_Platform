`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GSK6xzr5OrpAQe2HBQxoFpyurOG59xfAwlj6U4oqjQqXZ7NCeuI7QOvteVrDjqdC
3TNlqOW/X/A+ZAgnOKCGxh357U82i7U3GDAsQOpOkGq/JneKWKg12T1m067imOSn
D2jKOsryC0LuMdEdsEiAl0fWfFIjSPL+ztOT3WX81XsU6oudnl8vlfwMhh0QuDh3
hCdW9VCw96mRflJBb2QX3uxf11cJWMqh7ba73ySpQ3m0/LP6juiTCLCFqOUCwqhO
WznCWTH1R3qpd3VxM9KeHdCIsohx7muMokzJGi+xL/mGJJtlxXu9GsbNeD6AhIvX
p2KwfxPuB93pe9UnPYm4xOyFPt2nNomASfzCwS1bFmcjCIaRn1p8JirxK9YfBajo
aYeiKcuv/gaV157UgbXlOg==
`protect END_PROTECTED
