`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Anew2h4yk3KUJT7GfBAPHFnBpDjKsVxoRJ9PGrxiW5oWnHgwuU9cV/qR0/t1ztrk
FjqKWsqb7ijdQr3ZwjqPL6gTJ8P411oBrlXQdWkIxkCJ9kngBqcXEUQjmB/1dgmR
4UrQxe2/ECctwWQg+VLe1oTseUXZpu4X6Lld8+UxpJ8N/afLhnFB/G8CwX9IQEXa
NysXsCWC9eS6W0n7WZvAeeXDXUEGCoogO/eQbpbOVn8k/AC25dix0/ThLDmKBDiz
ckz1nf72uV40TGHM04WduXkgR1zCOQuCY4hTsGQJORi2h84QlOKbstpNzK3/2ani
nmbOFejKTbYlWVbA0wG4AWcDkysK9DaVGCDEhur2F6e4NAipBcRv9b99Wc9FRDQu
28g9yAMgLeA+ZMlXz2VWqrYJwt+AzMV8saTrCJ02fVSSq5vleOWBv/uUOLIgWRH8
MgTO07oHcktEahyk0D3SOG72CcR9YxTAgqoCoLyY7GPLayyGjYrZ/ax63+OrlVn2
ucBsoPm3vm/23YJs2fWnCCU3xaR4j1OZDkEONF1djNszEE9y5lr5yWaKLhngR34M
bABYkackqMG7n7a0T4GfGuWCCi4k+TXVPP/ATce7Yqze+yucrHrpB2lTQfxi/qnU
P1pkhwehWFEL2scpcNab+c1wp8Hoq/Jjf1NUTunO5x9ttdZFQ8eNHQKUGmcQzCzd
o2U4rYDqD8qntsF/4wvsEyd8ouqnSLlIIfUdCpWo3+eH8JWd0B3T+A2JbfyA4S35
hg7qb7WZTQmGB5ococJEf9Oiq7WuEL0+xEPedxJKIhK035AeNKtp4/Ygdqdyy+Fd
38sMYXgxO7Lo25Syy0l7NQspHChrDsGEXq5oJrTwaeXaVl4cJnsFgAnhmcJzcqZW
kZm0kwNddTeiYWUMEEwwo+fTwFwC+WKO/hKOyXikcpqv1OvwWpZB3GeeAO1MX+Cj
1/AzqN18gm2XwRiBYE8VB8bHMdZunutajtQ5ya1BALDdKy9sBV0MNK+gQxl6PTfQ
9KUQcvPFtfyAbgmC05dMaK3EHdbVvZf6WpXv95I9V12qpXi+VePKBDjYfhzf7cpV
OqpmcBmjdLrcRnREvdsXfqRJp41iujhGhqfPEKYPDNroRaPiX5H8wz/XFkkOa9Yj
AG1jRnVNkENKhc/bXo5t4svCwwP1ZJEGvT4pyQtYwJr7E0rEZj3WgGWbUNywXQo8
SbGAV3YnRi6lQQvnGdBKxhm8rBfSK3mtBpbN2SQjLghdVYZi8HUDfrOpC3DfSnHZ
x9hwp69T9skKry/7ffOtBs0rfIixfZFqk3lRXfg+sR+Oo66WeV1Q5EynzpTb0v3w
12uH48n/lE2wHG5i5mBQOa71F5bMVGE3ncdtcUBm9tPsgvVz/pMplw4oRLLIFAEP
GOyaErSY2RT+NkpOuPxQ0g6+cVo3UxNyBjulYmEibi+KAQAKrm1Mf7q5I/tLEjn2
XnAIumiCOMZrxwsFqfgzqmuNJlwVWN5UKFamdABZ0g4RNkJbg5Vo6uOMOOY0Pm2U
k2otJDuEyMdMXqwk+mq3E6+0QBFfuDF/Dz6RWLzzJJUktChq89CkT+rWLhScMR34
AOE+pVHmddsbN1hMXJmlRNKIAvXegQVCpwY1Wf2OEnVCK86tZtuTq9Uv0s89RBxh
dV+7SAB9elb6CNsaMWevQ7A4BremsWxz25c4Z5oALNOzRMUlYGMgM27VVFm6tn4F
CUSZssTXiONnH0NsY3oQCacZBQoDVjQdoKV8juUy615dtCgV6rG7XU9EHty2MN+X
qQk96aMjoP/1q+bop3MHgBZncZeXduLriWiXKlWwTZ03OLImZPA1st5gTGo/r6jW
lO3NgQwbwW+QLuj6arK6uFPEh+2LHusWeB7xnCqb3e978h2Hti5dX+HsrA4SsqnE
mgdINmc4ZFmMu6JflmaiI8koUDRFWL0xQGz+81EyJ5K3xiLYYhNur/PEFUzPBE6L
f969MtfjdeR7qCWg5b9OlGPRAlh1V/p+53KswHdCud87L0/V91c2gfr9oYyE58sN
hX9xqZw3Cfzh93dSUWVfezHgTDz3j4pYGHpmVDhWo1M/L1LRxsOC8LobFlX8XDij
W63JmLH2pXttp4TVzeCWKkJMtYsROutrb9PlBI9Brc3y7Ex/ETN9NP4W1hA2iwOt
vL2D5UvDnF9NuLnR1aTekHiKQSYwCn58eFxPKcXNDXxhf9+Jdj96eXiFVVdu9W5F
YnLn/1xDCLAUzq2XPBvoxzTKnfAyvLSxYqnpC5MqYvjQWECnG29vPb76GviWSrvJ
Xe9RR/8fpbLhfz6K9FSfsWWu4YIE5/J6O4SbdrCZSHrn3xr75IF4Ymw/hYJP9+dl
MR78WXj1K99q2TVth1GRojh2Y+I3snw+e5hiRZ8yEAR8oW8mZDYMPlFpAKB5u2Im
gB0t8nAgXR5TTb/rvzP5kCyZpBfO+IgezFw/6N7gFbjzfeqOauHTRAfz0XcO161I
7qwUDBOZkWB06Ws0iWpH/2fjMwGVN4kPXqQJIifKskbdM9mCiZWzDxj6uUicuAE6
NfbyzJkyzixas242r6NcZ1t4+wRQctu9lzD7RiqWNFyvVrqdwtwaNLy6ITGn/raz
`protect END_PROTECTED
