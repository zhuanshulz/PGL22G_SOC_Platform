`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V/eilW+YwdwHe8E0CoXf7FMrpbTi2NyuEx3MYm1SRjp/v+up7z0vftQSKohtOqGc
4Sh2K6Q9Eod9zxvuNRnNizaaVtFjaZsP7/lDGE09fbvzmIo6Uyjpg6a+uIQkM3Uq
yT7ClT/ymmTRQUj1uZpZ6Vn9X+l1GKYLDCUYXgXrsD+iXdJwby8f7AD5tgw0ZIOQ
hJJ5ICW7etqUJTjyDUJo+y0RFMRQo67X0vMq0/th9if1FVyKWTmv/PV59JzOhreM
Olei1LMdO33qlE8hdwlDby2yvTCLk3Q/Cn+1Yz7yF1fEbckMLsnaLNvQotBw4Ebk
X6Yia14vz/1DaS7bRQ+omDlWrKeivQeaWHdV5qAngBM5LAgrlItA12DlALu7QpBg
hTfyUt1SDrmDwt8wzDBjTfT8iS0mk1XJPOyQZiZoUHbiMPmJShnoLmQir2o3gCqg
w0SSXbFZkfD13bKU1ygGTgXPUm/P2wrNdTgHf8K0BOR5ffErBvmyObjoNlbsYx9c
c0QnRynWmE1h6WOOBmnkGaED31hf27qIhsWDgcqbl9yDykwnmPplMejKO1O2ZgmW
nEmcuzKbpWqlWZo8jnt0tbOuPVwiP/13j47eDLqT8uL9BGBjUqfhSaz9wcK/Th0e
ivobGc5X2AiclvJJmPFcBHdUbzT7IgyGKbt00+QcQNPRT6CnR0sREYa9L5SxDSoh
3uq5JFCrk0137+3Km6pKpXtnDwTiU3Hws1lRIgQqtrqOwBMBF+ZL4rlwcK0uiuT0
B5A7bGZiAMu5sdiDUQTwtZX4YT0K3Com3cdnUlySraTVw61UF5X5WruB9isw9UpU
4zIEjETJr2BRqvqyNE7tukL6iiy244Sa03frilSv0I6A7WJKSLGj3lVfNJSt6PFZ
yIp2rF7T6EvklxOjsMGGmUEC1Ay2kj/KCgdvmeDYXVmumdxnviwGOnGqUB+7M30I
pmBsRws5jQC4oigPu2kx/l3k0rGSIQo5+UwrTe4cy1PWFo/kHlm/jA2be7KL6O77
RL4KAZw7iE2lHI3XiaK8WfD5Z88H/b/+uu9POyFnd7V5nuH79+Oi7bbooZoFP8j7
RkE2JXhkZxdfmNbNDCMkRoRPzrEQSYaMg4R8G0zSEL8yCcFE36orWCSgdWMMCc0a
ZQ+vzAt6KszbDp+tTs1L78opwmRjIWnOW+72bQBFcnBY/4gvROd/kEHRqthSerhK
U7w95q6c5Aswge0PyejeOVHrKQTGNeyvIFDhQp91bKHchToxNTU/KNXs746TyJFJ
qqG1TC+lVm7LUNYQZYAhePe+Oweyp4vMvpEBhanvVc8W+MXn1zLh4n9kxSDdjuci
1iQla86Jwr0m7/HnCrXutEIuAXK3G7J8UyV6cwrcSaT405Ul/pKrBCTw50P4BtXa
yspbNdqgarRoF6YA9f0uoZqnLeNfSrLMAml7+Au4JAECORIePWfFjj2FcI7Oxfs5
nXoVO+5rErFpQGVOu+tkGPEAsXKjzvj9cKibiUhEFR88zlbL3TqfOLp994LXTP5s
u5ChkaGxwcIhHJlGdGhjiEb6ILeKkwtTMDb6wZtSsYf3ZnlGlYnzfR2DXRx37mfh
/lpSLry4WtwgUlAopAXmcECD+vARv5SMgNoOmmUI6p+yxxFtS+XdnDDVXpPMagL8
9P4aLbNEXemDo8+sM5Yb2/HWjQZmDglzrwK0TmKIz3X8E4N5gSzzh7zM7b2dy40a
HkHZ64hSKqrX0+7jefRbvKH5Slkt6qERsjzMoynQ/h733PlGGfS0LoStIk0Hhj5Z
Hx1/31qFJqZL/MI3qFmV2veG8+0mrTqr+P2t/8JXg6SXid5rdv6pqZHmGzVGJXWA
w+9z2xcAQTC/fOmfJop8nK8cdxXMtipzS25qc7+5Ge+JcCIQakS/kO+YrpBljkdc
G+Q5qCKGPZQVteIckgif1UaadoFBZH1vlip8N6LfCLKUk/unpLJgEKvWGdDqqn+Q
J9od+jGAQtFmN6eyPFJObNl/nZqF7pJHTJ/6UvOL5HsanC5fCDIz3iBkKYQ9OpGn
yPcX1r1wcVmJMi67lyYKaDNPIV8Q8w8K/t7+WYw0QiK+Iy4c4p6gcPltBQ+K3IHS
2ohHkIH9/LkEN2BxdBmodrUnMEJxBbBUJEkfRzVkvQ164kmRjPUXvw4rNzi37cZA
F7KUHnCt+EmRSZ748qNTeyja/Gxi6xZ5ar2NFv4+qkgHv2PZncvW9+QMvidtTPzW
WziG1tgj/7SxvHoHP3snJDz0+f9M7S/ZZITVopBikeD/lkcIvpqBFQQz7d+5vP4J
5zSo/U7NtT9gCertRsBh0ubb+9sDXfOo0uOVlVXWCz+Q8UjnhGSdjU0y8sRcQ6pF
sMwFUDB4J5JcQ+yjd+85r7BD9B6WutTmu4cjBr1YEhV7A1dotFNHvc5e0tj/VfVL
t/QIZazA6EtahdCxMNcIXZPUP3qNi+WwRKw7d8T9ok6tIGcUyZYl46l3kVf/MWRb
MrHdQciFFAouSdljK2FfXnIiPOCGSmyBI5UXn3evjU2Ds8R9+tP8I0xOMAqSKUvV
hckWQFViKKYGiYQ40vyxADfmVL7I9Wjk9XWZEFaPN2ELqogvmsSy/4hE/2jlYBB9
4BJoIRyqA7PxjY4yeoiVdqkzjNIGIRuhBeWhuTeydV2PQAhGFDXQbqIVtvRvTsVO
Pq+U4jYSIWFZQf3DByyPzCbh0gcavtzXcGe9/E1NFSDonkq5oKEozVk35DBAqo+1
EACGyvqJhCf6I27BdhlfXQS/qEXrGX5Ibz+AyfMZocGrN4BRl/gZYTyytc62fl4i
+Iy/PXGY8aYh5ME5oOpXrikpf+fOJlZPazy1eKwdrbQzgvHke2uuxWy3Vw672qat
Lre7p8+I4eauu82N6rIeeDyBgm0NbszYCMpl6CpOIGm0Hsxlhm8yrOX7udUCXeaU
mjACnw2+l0SzTs0ZLri5AUQKCUdnIX937jQ4m88QV+r3foQNOeWsYAfEqtY+urK4
pLODKKLP2eD64NMUp5raSnRtAU9w6sXT+qjWROfNSnZUOH+MRAxT/x3Vei4iCnJE
YxzOQn97rkkvsdkYstzhk2Kxo2DzFlcKYRku7UwsHm07aHmKUSPs0r6+Sd9iMvdd
aqwnIhaWDI5RrAfVjezVmDM2k+8g7cowfp08vqtYTc19pXwuxddV+0+NRDH/Uu2T
h3F+qiupd6AQnh8WSqM/lP69s6WYOCG9+M7QuThp2QNfdON+EtlabNKkCfPSo/ij
6zneGZOsvho3sn9uRh4MSKk/W3OeXyGqbCV5xu0eVJsiGDy+voQpMDDtX+PBAKXd
sTxlCoGfoplHeIHMuQTlbfXP0d/XpSpk0PTTjZ4XVVJbbZtWSGpU8OFZ8sgqjJ+/
hetXeYrWez73tLWZ73b1Qe5lIz0JIHDb2rXGLB6zsbovIeRuc08eIv+b2XJ0KMsW
GRn9PeVjuyBXRiO2gAK48Pho7s7fG8PcyxfEYKxPW4il0+oPQ7RJ8cLycgAKNcBA
SpEDQ3FFxntL1/8yebyssq8v0KNE/MGoAEnSVvGYJdqWdE3n5A376viw1PqaMEGN
5v4NJTRVF8RunTXMCfXfmYvPyZ7YyCEEadK70yFemgqy41Vq5LQW4mlOFccN+JMF
Ku5b7q+93rXa/Nce/vgMk6UIU1BbyRhs0nC9ouD5srumMIax2ad0ikyBcL6vd7BX
twn/Hkt3ZC727jv0Udnd44ukzrMWnWvsNNfXj5YUIAgQ5TGkhxkiXEwj7UN7cctj
uAX5jxPgRbtoXp/BMnuDaYwCPCCu/jK35EuLTHPlkaa2hfQaEdmeqrxnErcvSF16
WriPjyvnhYeVu9xJXCR3lfOTJiIWoXfQD4Hv91m/HaphxEL8M1VW0xSDe/cj+hyS
H95vStd8O8JVkHh/IuV1aEpMNjdAMxw/8fs7eXmO00nXqqm36FuWsQAMrXn+o6QP
9JqQMplF74SRJNcZE83pxFKlzsz2m3AQO5+8pjUpuibguxubG8j3QZtd022UoLuD
od9Hf3wKrM+d+ZXjKL9/Zmm6bgkgiOq2FZBFp2ibqBacxH+ldI8GzNfx7AXMVJws
aA6lk8ZcF2NiB8exUTarS5cf2+mkR1t9e6ASa6ihVK9CGk5DFrf6JwDYoZ/GuX0D
aWqn6K5cC+cg1JTN8PnJA6hxRYgwO8q/my6EoiPrDiyVApCj3vgHIpjb5ST9kXBW
b8dDX6fJPcGDYTANwqAObCvewYPCSTsF9GFee4XQayz57cDL1wFHYYWYbzi+yQE/
XWfK/Jl3Ha97WD22chvYB9eUa0+xRC6AJZID7PZAdbsxYOELwRwe9xtGjZUbeG10
VCfWYdeLoh1NMljoIjlvZ9e7GmgQr491bcbCCLph3q71k5QKlFnw0c1Nz0QUuV8O
n5tI8tpvIW7k70FMjO6fBkSJ+x79zSkTr/iR09Fjlxf7dBPANLju+7RcA/fS12VL
sTChHfP6cQng2FjYEsiHizAxcUYur/dPuBY0ydejXoic2jGpaBp15kAEuBVq80Rb
nROuvmatLxSlXycdOYV+SkZ0m3cxmhgRGrI5zoOa/6dbeb21xRi7RYUrNjSPx9Ki
fO0EWo22UX9XdHWEI+p/rTb61UXiktYzad71gxoOeC7CMqGEFsK/vRewpwfa57Dc
NWEbfWAXbZRGaeJBSHr0VfNLF2mR3ENsnepaVeHunhh8/d0KlteQ8INRKNEE5ji1
3E49bGT+8HsEW3YCudzFPOQX+d0A2LyvShZvgIV1XVN9AsMCCM3dPDh15nrdmEmM
JDa2FBlPPHvFAAD934hQPF/Pnfsu1Pl9IiMzKiZja9vTKUz18Qfe/n9+fWByPWFm
aegrnJYc5KIbtiZlByg/eFz0A5HJmTcQvGSlMemaNHh5/qfgVdQPA59tKYNhh9xe
5/Ml6aLd3vLhWhGQ0+P4QX/w4cQY4rY11AAwow2bcG1YfDbg3QOcc3rMOCMNN/lD
A+aCoCVyTEU2rx5xJgYp9xnOefPzMIyTpEhf7RxkLsi3otKwOHe9J/nhv7QwDHPa
BJ1JM3s8n20ArRyVEsC6iSrGTR0qAQQLMj8XX1qPR2ZJJJWHZ1qlBXOIef6OyFEI
eYnvLfbBjpbAVA48V8LuLAQosu8vfoDJDXS4pAox3jvG5i5ZjSFNhuuQuRVV6/Hl
0mreQuk8qmLi0cCV0nLn4Y/PmS3PrdxrMkPVIXWvlgCm6o7ZmY6hAw6XuHN4e/+H
ZL9McdOl7rN52DMxeyWM3aae+YsZHRsjRBaQ40kX0ziYo3FbGEpTuiGt80RzL+vo
azr8NGTNacSDwJEt+GvRAL0BZtgUV2eqwf/AYacSENEGru8jKpkSs33Tfglv4UCm
enescJvuluHzLOTLp015jUsNAtqZcIzYwXSaHrfUQLD+knxUuMlJd21MfF2BDwN3
Q54AdBeh0KOqX/5rdjfluC3wneg727BI0ezUPkki6c0eCn1JzZTNNj74cDwtgNbR
VdTuxeHWMdu5jF22c1UHCPYvVPY67qnEHaS5LwAjOLHVkoNoW0v8hs3BcAlRw0bD
ct5Atiy7jCUTPo09MI85VRQh23XnFY3DhcsPrHwb+SRpim8l7hJuqSOUbRAjU2C+
YPwUBdPXMfV3Qc0fcK6L39K04VE4Oj9CWSUbGsI3AApqOtkH06Dwadif8mB49xko
HRS9KpMOpJ0sZfDUCzFgMtzXUqTVBSR0rjFsEQWMnGWJxqwKVxxxfN+Kf4R92Ly4
w117/HVKIRqpYUm21hz5Wd8YN6OeMjQ+kVdosEJrHZSTRsQEdxqwlVKNhbkQXaSn
PHl0iaiVJBkncGxZASnNVgb0shQx+5StpPu93e/zTW1tsiiIyT8GqjnVjUqMH10K
e/7TxlgFuG5LIwkFPU+l25Sp2oV5IZUfFjgElBZWmuwLSe+S0PPXVeW7w2IBza1J
yAg6GvDUa14GIcMO36NcTbBdwIxhNho6Nvn1p8txp38vwZOoqEIQnUnAiF5A1AvI
dv4daCGLJeCMcHMa9+rcXFUfv/kQhPCgMBbYG0utrV6ZVCuuqNPS5TCIdbC+yAJJ
RNo0VNs65K42QCudeTtmEO2xIyfPMIvKAE1YGWGifVmvHej7HU/GxFeu3LoxXY/1
ppw42FOzd3FUQU9TQdnOeB6gz7ctSQkz9CBDloGDn6n+tbe1bf7FlzuqK9MxPRgL
XVmVIgLMhtKHg6n5YajA514tfldzJ/zXsoJy1dKByg4TbX+CusTKXmqFe84nVqi+
Y27yhICoXpbflTPdhBaBw/4BbWs3Kdmj/TN6DJ14L4YNoRf7fSeCede32J08o6MF
GOd2oFwUNJ7CEEhe/a1C4UUc4KoKe158wKhGyS0RrS83fxPjxN87h4uR2NNtXrAR
+bGBmqID6d4jjLX0JALyXaE7A7hw/L1NTz1ZLcbV+qrgZrtQ0khT5Jyarn9yq/Ur
WhtklCKAP0ihHBVPcgmM5Oa0HRJDuR3ISecYTHsI68eINsoxti/VR4DkoeBgmTOo
wNG1cVrzgEQl9v57TkRVqW4V9tNPN0MxP0yJ3avhmA2ZZMbOqE/v0vIp2/hFSWD0
hL1440BAFRfMi4tabQFidEM4k0ELXaY4NkXP/J103vjEsR0wImsGIEa+wWznmRMD
3U7QtHHgEgZSLTtmGuzYRlxGFdJxF6cvXq7OTzug+bD/7w2fYbhrBSKVR3AEej63
pzQta425kb1aauf9cESsdZhEPu/LvROQ7xGep/EaQK3J1P5JJ2j4LM2hJ0VohoxE
h4o2tRQye76g7C0e5/Evh+ci0RHJ4pMlnWpLFYRf+VWeGAvAJJzyNlTzEUvLH5eK
t0nkYEHi9h0fczIidWcojfVbDffLSy5aEWlZnSQGPbCRWte8OwL7JoM0GSBApGsH
aSGFmCID/LgGEGI89Sif3zAECxgEJY3JZ+sDaOeggoy+u01+Rdlg8py+HSWZ8Q65
fSDCnG2rJt78uJ/TVlNeRJGBHBUNTDsrEB3YjwUOVyEaVwWihcA5NxmRbamKSqck
rCNmOEaOiWHDTeuy2PdT84JTv6HBzvUNhL4n819c7xsCNd4DJd0OpS1s1VwnGsJ6
OA7TZ3pcZDrY1gAEiCNE7493DnRTo8maFA/TZwMBZBDsVdI8XNNJHdTWm0EE18bo
bxeQj62ey5e30vvUGsUwC2QSuX9i6WImGQIIFeBbRIp4XdVB7U0MO0mTk+eDWqKe
zXXTYw6HpAgpk0QyHEXXCyD2kqhRcvdhs8dbMuXyOWBekxhBHmyzg9249GkSyio5
Ce6otjgnwF8rM2kwZ/LK/AC1lF9vZBp+QarmuWEpVdFxud3YH2hVdIEMHGk9Nk1f
Fkma9Alot0TIKbuogUiovDjXMf2Tncc38SoWLnAsxcrQSJDggUwLHJU4wHjkGcIK
XpX4oeDegmLIq1Cj3DrxvGk3NcSl2mrTKK+//eRYmipK1XlLCCyjgvzGILNR3yOu
PWS3I/bATHqEQrha14/vnEB7A7t86ZkdrJPOHRjBkgbSi7scf5rSHRlubFgFNErA
LPK0iOexMaEynq0+FRFLZcSsGcv7x4sh+oxS6jf/FyIxUjWaDKs9/A/HEfv5df/7
OQiyzVtOwAhuxjU7KoCvp/E9RAZ+1Zr9tdN6IuS9cUSwaS6Ew+Co32c/NCFY50Rm
N6K8pJ/qxlR5FerAZIt3iU1V5kkJ8eCskTKp+qUhllUdOmUswUBAdvUUWh1NnmhZ
BggG3MwGlPat1yPsL+jfoCcWKQxI6D+gHmZouC6wBJiiwPHcKjXcLPFEhRJbjaVt
VJTl1PbEh/7kqQhcx1pWcrTq0+/w0QfJG4c7ZdZ83iO2t8BUffeQB/tIlRQM/o0/
fYDU50kIXcUNhzvICqteHenNpSY+jszWiMDulytfw0RZN7ww34q6O3urkYDCklf6
I5YleTN+KZbWsM2bEMYKNWhAQWwL3mOuQoxbbuMZo2ttP0PscYVUuxgMlUtpW0KO
W+ZQhaT0q4J/dj4ApzPeyqrUbM/EXub9vALgyerkko4lQ8IiQRKock8bnIAOxbVp
4jMB+krCDLzdqqh2BcxQPygOHws+2mLTKz0ikqFbvMD9QrD7N352Jic0rt1qxRsd
dXq++2jnlrS4wa8CQgMWU6SALIoIP7Ma5E6kGOCwpOC6kdiugsDiF0KpwL0pCFAr
D9suHIMS4aKtlXUU8+wufWdAk4IgE/gI3KyWfggko9mfVACBIK/rVGuqMKDafJmy
OYi3enegAhg6jDa0taWS+ACjpcDdZfoIDYQDNW6LL1IShdym0HqcZtlxAwecIdSZ
0wbm4i+4w/2wjbk0HDUWXLqsZyczbq0FU+chWFjYtEjNsqLEDixoVivqTcKJJKct
8GRyXsIcxpBGX+lVsgKDAg1sW8WvpouogyklVPI+BuCv/LTAk8UGsG7lIVk28lqW
Ug18802KVj5+z/xSXKJBCElRXrSstaF5IPkiDR7HdRJKPEL4EI/GVpQ12S7IaeIh
1hxBFrDQUDeIan+LTNnQ06lGlp+V75exhygLjPO6CEQKDLIYxOCLjOr6/T6jtyu4
kIQdMJCkLKvyEYz9OIk2P6JTrXi/TtI9ai1PukGQvsjqYi4Vc6+6QrhGhKv0I9e4
KIKH71LOFoDWtWkh5pH0BlVfEZED1+yVMnYGlDkFP5lblb8rUbVQd+tAFUQHUoA8
l6EIX5s4f69Ja6wcBaKAdLO4mF0RmINAw+gX6AfaLZHkSfcLxQit5/jH+uch9c5W
Ozc95jpYHT6MQWsEiRWQYnrQ26qFfXIUZArebNTF/up2NktaYjjUiUOTb1DGOrqB
ojb0I7Eo/QqVwnvvDGyhQVCLPg6DpmQl4SvPOfesp4CMZ0GUddFxgkfgOmd3UXBv
W3TAUp4JIeBEdyQqDE3XywquH/dR7fNrOlNcmTFl9an8yHNEtKFVzxrjm5N4bTz3
eSs3nKy0VusmfHJcNbqr/o92xZuyamZjiTQknFljvryZZ+jsZTH8JjOzEOo9KHlK
x7kEQAN+StqkTFjIrHG/yxDulWREWscQ5sHxTmCeuHmYPhuuHeNPvBlrc+KfvO57
qY8n5HEICTCN7vtIKLTdaofZaUjsygn789EHuhY6rfXsAsyaAyNu9iiMiGLg29cJ
4z/NglPAh6bPqmG3tYGo1YjiZRsbpNY2DwrA050eay2Htd3mFVw9Pc03GAFuLRIl
6baFawzwHp9KjuJtMaEBnoLO9htIgmTGEtN4Qlh4/TLPD5E4cSTpATK6cZLRI792
Kf8QHABKrVmcIQ3JxLodQmZHBpT/CnJ8xeuoGVHv95dO2c7+ssg5kXX8oGQK3nfv
mUvrvRZp8vC6N6v7OsqmFRmeUkKCTAVXvSVKgwhiDtmW14qHmGqpUfSWNukHEsrL
MfMsO4ODPm5ueOaguSc5U7UM0PWjBf46bHLCvRZ7SSi7FD7OFzThslSBdbkXIoJX
L2g7mh78S7qWicRokEFMwc2Wl5+/BmHsBJyP7yCpliS6mIIDrHdYb/6GM8yl3nRK
zQs8oKVK5dFooRs3Ij4tPdP2dgXBRGaytFN38ayu5XAsbwaVQ9RwbnrH3Smg0yEs
is4zeuWLpACdsMOPA6l1ygHoGPowgliPLXNLDLHsZoaU518QBeXa/17+LMNs+uxt
jYV3dZkyWdENl8LBNGJuA5DXFO6HrvGcKBzxsXnXZkVYo6BjtfK4QT0he9xSfJWi
QpNc1XosejXgPcm4Xm530rk0whoTG3z7q6aCPYvrNRbAoRIW91xWrhdbFATH3oBx
oKZHTihbU4xvjNmXRu13e6nOTfZMMCMmqERg4yGOcUTttW+VjNUIM7dHCWUkvX+q
iZRFhCdtONnRQftVo2kaEksptTUyu9fanKTPiadRILGEsSP4pPOsj6jjJy5nNojp
cCi9iLZPiFLu0opjm/Gaxp/UCv2h4OrawUs3NYx0mLPpHPwTGBfnlRSTIEcH7PzI
iM4O12tDR+wfvKM3Umi8eNg5TyAUG0ru7YwNJRblFWtbBSJ3sC3RQucCHxnHMGyI
Db3GbusEWbuYSyo6UqX6zKZTPY4I3LaAKQR27YlGrEwXOuthWCw7Rz1wi/cxFVcZ
uK0S2ytF2wP2ePr/B2H2UXUetQKeDHm1FvLhT6OYMF9Az7FMSvkrNxEYrsR7Iv9C
PqTVr60TRC2cuQ6jqUkMwORVeuqcgMOKavuiAo3q9pIw9cr/qQ4/RDyIs44kNAWZ
7he/cRhS1PKkY53Zq7fuRW25a6VksgtJoqhGq0l55E1GSQ/B0QUNzggL5rox45Zo
VZnFLWJoSjBTFWTJFc881aVqtItSfhImR/yhjxm2MtP6vYIbUDFgPlIJBgIuOSQm
WgD+o3sQYdrbY8s9wXSDQxIO30lfFk0w/lYCLwHa9XJGr2VoJynJWAS1L12r/Acj
XAI3jVf4tbkUYz/FJo2RuHRZSclPL/Th0lgCWx9Zfba/Ojl/lRzVOVPlX7GA2oEA
PH3Sb/9BXTxWMkuW66l7+bX1VlM1QUCMhmpMkyJr0xrxQLUWEFjftycQNXwzeEC1
OTjCOCjz4Gar0N8Y1DmTQQhsg/H9PZtISwEi3M8YhvyHAF4LTurOuU7KpAlBGAbA
yU0/jR+ZZtruTldd09kmXExvNdqIBr5w6+K0Na5CEumg4uYKtlzebFDabAH1RczU
UdG1FbEwyxefzgg7GqwaLqOkz0xusauX59aLPaZY9BUZlPwPiI53MKM5zkTEBVtc
49LwSP2Vh7WU6nr6fuRoFS+0jIShCQYbHmBZYtXh5jTt/xc6oEen/8XWQ9KzbvGx
fZr2XUj08PrNeRHC0QLDkVtKiRok7LWIuxbHytV/4iEb7fvox8WXYYA/eOf/nw0u
rMOoFhG0T2jbaZhEbwCA110H8D9yfEweEDa79uH/fi71hXFEVMcjZgKDsStLFir5
BNs9J97kaSXZ3y2dxb1Vv+oIf0XcW/evJhZH1nw3wDKHAYSMY1bSR03S2lJIlQVN
7XVSnB62dcRh/3bOVgHPKNsYgrOq+maXOoDOx1dESAm3ihMZxQZT+5WQ4KydCCub
6h+nsKAqm3gE5HuXPUgf6OxU0Bcwd+p0Te/K14ICAp6x0pJV6riJZTcK4FWNrkaf
GL22Gf8mmC0cixLsPJcZT7xr6bVuMVo4ZcLT895ZIuplDk2keYuw3bvfz64kwRBO
puJzS2CEhBBewSZcofo+hDYfKIr/4jBTeATjrYBD6y31N7mo29jfA3D1pNOQ1kFx
GiRX3JQmEcCRYFWRsFD2496bkzJFVN7ITApMjjkYMVrkcKu0pGQNyNPzWmbkllIU
9cvDD+zrq4Eme1ZM55NDyQRfcOfymVpSZgTZ4AlMtiUOobbvnp39X5bzSlLmTxK8
pCMWxEGj2umH1jmgncXqC7MGb9rtKcjGPJg3KGRyJf6+QQ/2R081XG2odsb87p3H
HI4GRuWmGUSfIM6fXRiSXuM5/UP2NA/wx+y5c7EGCNnAw4p9YpQyCjhJVSXTb6Mg
isvTVMFSDZonTAGRQfJTG9MWn1fdQP3hgK7dyM5PW4k8SHz/d/XdFiOd/r9OApVO
CS/AMqFj70Lk6w4jL8O2v8Rud7j0zini2TCq8cBaZghDrZwQiqcO+ooeWFVMz7J6
Fmldlart6APCqskQFQr9hdqY/1XewpOekF8F5OM/H+FPVejLu/Acd0NoBXOgzirm
E1bzZi9OUsw+TXlJol8knGjqdaUtngNsMSOKaRTbsAbsRz/RqHGAcW4U0SZPFv7s
GQ9VfrzFrtJPQY07tWXOszdVpcy2GW1cU7mh/yH4QTyDiSKLJ7Cta/9XFBwra8B8
wDdXlAXzWV/cu8F8O0KuFDEj0V0wTOvvWKi/x965bzXROdDKu7+7DRE9lgOUB6L5
0h4iPQPRORklnvmr9lE6/1fKm8ek+dNvV3/ZZmhbnsJPgEJLBDot7WnKz9HpkFBZ
ZZcWuFwK2pUt8lQJaY5lt6mRr0Qj4O/Kkv63mwTs1ew94AfS+ilI2MXnFc29DlBE
kn3BwJUdziotFYTUhKiDMdf3WSIxgV30jDmZHG7vcab6CnMGmjtfQ+dfOVCG/4K8
fv1Lxyne80bCwOxmHutvKzItoTBCoaZDMuQIbxk5ElosWdhZXUZl0vEvQk/tj+aT
Un0orVQHMy3/BxQxC/cJjOQaZVS3szlgPk5i9mWa24q2bWpYxBO6VYREPGuaBuUe
pJiYTdx2wtw8fNrMsbNV5Vr2SSlN7Q+NkFMkf857bi4mR902fY3wqAtGTxRamQGi
CadV8/Kke7zX+6NVcz9K7ui9whwYSaHRHguGurji3lQpc6r+UvpubpNLIEnyvRfW
jjHOJU6y3fbPQ0H3KMwxA3xXO+xcl+OHLq/2Sw2MueE/vFcH5gbTCcC4bvv4fB7c
4OJ3NirheDoJg1kPX2SR1ROswCciNikSLCusetmNCz21SZsgwp1XYnQfxhJAbdaC
xgvZwNfsHW9VDa8wM6WGXA==
`protect END_PROTECTED
