`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fzu9siCvlfxP1T0xRdf+IX05JYNOEIiz426vFDFVdE2IUJc/qPwpokPlbp46feNB
wn9n5M1G0DoMKjtI+ENfuhQdst+hVgkOccP+fyfgEI+E3n51tQMZFeuQKucwrRFv
x2efj17FXYmmlJkU+f5s4nLIa7CGhuHnsaYPoAub/HPTO4VQ0LuaKDt8ceEwPyOV
Q9BnbleJkKipSAbXFkB7YiNCys09rUvayyQwDtIn6EsyAdJUNXu1S1OPlAR/Jcy2
/eZw/q2WoPClCwiuSjrOTutsGFyu88OD7Y65cs8QODOI0Iua7sKC9IfbMmIHDVxK
x3/loLvwef359IZaa0OTQU2cah0khqEUm/Urffs3QbVIz4/h/dzi7uXPJKopSHHV
yoUEKVxEMFLJ6tZQt1764hRjugzOZwtYlUBiOWnsjfYlqng8KXZUywY2XJJ7lo3F
`protect END_PROTECTED
