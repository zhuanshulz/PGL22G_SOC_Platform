`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xC1QffIcOVIe45aG6rdiCITef35jNR4NOhG4IEMB6EVAH5rvL1uQnGz8FyKnI1Bz
rpYSIqnDg1Twdhca7kxYmoX5V8UDJ5O3HeMj2H4S4Y3ReAXk+Aq0QLySLGi9NfYo
oig8/lFRQ8015oT8JgyMWJeJHf2KAhAoqLSmcPnQqAswDVHYXyYtJeSNN9Bl6Lfs
DjGytOTM86u/Fd+awHDb6PsjDIJs8W6OEtXLaIFDpVdyudx60Oee0siT+EElaiXk
zlpKyaUZg5vp83rIsO4DayFoo6ZIIWuddbR1dIwYSxiez4KpYTvOkHSSCotOCX/B
aXlxCdDEk9JPJxdX4U9dq0TTFRC2XPw5lJ23U7oouwPbPTGS57+9AhKPfCe4/YQ2
e9v6rT/yuwL4tLBnoYnYxuyVAhoHifCyLy1x+wEFdueMJ7sePvlVb5wXCYK5Ovfn
AtpsP9eW5fSkRz2iePbpVbToQzRJhuE38xCdlMjY27q0xov6LVvyc41SE96W5pOS
fTW2yk3890cgypfAVrhy9YYGr+jBtoPzecIARLZkfKi0GeuB+5xxdRmwSXLwCMVI
yS2hi944o6wkD0WhrztOjheKsZsE0XPjgqCkR3cCyxyejVHhrnmQa+JrAG1BVfWf
UAQ/OYec7xI6USQE5PMsKllqGr10Tuw/qFZYtcKF/AUYmM2a4tsZD7/KDHUTSMoB
LF72jMROJ0jNE+zfXJuI42Dftf5/EW7HIYlle0P+BVjia1hDri/XH9tuVRuCurmX
bEJ1m1b6gm0ZnWs5XVLCFCVDdpa7GxT47JCsc/2DNOI8EgARRRzAfgcnwGkVlvTc
KWuPNWodHS/6D34ycymmeZnx44P9JZY7pbpzKse6k4Wgu7eD0Iq6J8uQgKs1ttWn
JuygZRiYqTF3k5aRfiqLMgD2/3pyIQxcxiAHaN66Wox75MuGUhIZ7+QKncqdseFi
a+ctzRcLub8pMi42sHVJ4vMVhQReQGKWGPYW3+vXztJzp2CI8yx0IRBP9Rj4uLNv
S1sApQfjoN1AxWVY315Oxc9jQktwJD2FgsthqePSVjeNaE+zezvJx3Lyqk9tubwM
pPfp8zXwl7uvbX6gByFbGWjQ02r5mvbcd/AV50xFSsvfmasbLgb0rAvpTMDvfUHs
Q4iex/iqGrk7UeYWQ+JIQtja4OrfWDZcH4JWrBe/kTB4d8AIDfkgzBh9I/LLYOk4
G8esmUqzgro0MGQsuTf7W/j8wD6GuWvVF2FjLabozCSdvsMKL33WfLTEAw6GVTTw
hNzsHJ9V+yo3EILlRWiczg02u3SpsA6+frYFjDIObFrZCpNG0qvugv5ZeLyOYqCh
ukySu7njK2QovNee6DnSeDF+uiq9vfpsHFiXA2dwOPZZ+ZRId4lKkkEvUvP/53VM
6PorNXpPnSz3UIbaB9iYYZ0JGBQzOePxML3XjYnsTDX/MU6MiW04Og4yBiIK82HW
KChrubQFLYPmpPWo/vgpmirvhAP2ODQBHUvQ/5iH2G6FkRTqlyIhZpwQy4VU2fbc
hEVgQM3fKZ8aGMAACf5OqpkjCT+6gdNa+Sqbr/h4JpBNAlHocMqt5smEApjAo4tj
s/xmzZjk+r55Oi7VK7GvXq9aCv9hxsTI2HiRz0gXG4jknJotIGzWmm6xL178C0Ad
aNWJYpi+m7cbg6lWT0pO9GS+rcMxvspDRBWDrKZp58xrYy6crcupEGo3v5huBJor
q4vzMFAN7wURT+rzLHOrYPx+Ar186ZiLbpV6jo/bqQI=
`protect END_PROTECTED
