`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
buJQ0v74G8/6BbNspXYInxNbcJTMyHL2WWwlbSDTKy34YMhELkc7aqX96Vra0q+e
/mQqBVjhDtwLOC7+HcFVsrT93tb+hpj7vZ+oOhJeSyyRmry5eXZPj23X+/UYqTSK
gUZi2S2TlyC4L/c5xBly28lF/RUXbG3ATyVHiWamQCefv3temxMrBu6HF0v9+wqw
BqsgYbt74JnjERIO3vwqJMpL47owfttTGakcE1KHZV0AS9xtTMffXc7X6N/uv/fu
zBpXp2sZc2f/uHNpYkCJ9GGqAX5DzB0aH47EhyWx1dGuc8wnwGTaCQh+YfhyCqF4
NocUz1GsozC8C4vUHk9LitYn4uFepBj4zKKvHL834cgu3lEWIbTYGdrvbhJDKQxj
CvOTQpKLHUPCbXVbNTpHC6GAQf9QQ0gequhKmfcC81kbt9SP03EEIwWhAXIWEswZ
YmP/WIf5ufq0lY8Eo+n5AM7oZC9Vv1CJMuo9SNSlNRZIm0Wgr4UsfTwHUXxCOtaN
yhS1tZQHBVzYwNE7ElFuMdku6fbXdOvAxD4EYa0RjGcVCxK8kFdNiYep6Y3pFtEp
RRc0hRkqWnWJgrLEpamTiH2auhngLCY6iwgNwos6BtpJ2Aos4cyVJo+M/Mrhbtwc
rkIdz3u23dkSFKgveTBH7G5F/ZDDtugzdvrY07cllBHIJEZgG0Gg7cruSSRCfH3H
afOin7K5lA6xbwXmPfDHc+FIftWh43c3c5Ck8STDZaAn1ToRewDhXpfMMjPxi62y
u1yUqblrR4NYbVd1ZSNKmbWmlpsRtp05AmTq89UOQo7seuVwXJ2jdjWivmQtx+YV
2bSOds7vSqXfBZGxx0pPR5sJIvclinnt1wKF5Hw+/QDHAR1XcRedHyA3TM8QB4NB
KlqaKDlUkKvvnE+JOzSZYJXINVnng37ae9dh+URt+XUe0O855zDEJn6UOZaOxvqZ
sC8+vX/9DsjVZ+7ed1SccocEFsLY9sMWmDvx8HRgc0WV5uwxKppjKildub3S88Fm
8Pmljudi3w2nhRl1E3dSj/2vpCc1Lb7G9plNJR14smNzJlVnnQOjJg08KF1Pg13V
5icQg6HKbjJu/Kdr/3ORT0L2Q4DGQSzgN1i1AZjBG0V4NaTy4HaNKEMWjJZ1pP6I
g+Ltqi3a3zUz2gMeAT3bYsFQ60LT21Y+IK4o8miZ3gGIekqV1rzSbkqib9jNX4Ok
HGihNSBFcIWvFSjLts8/GUrl/+La77YLGpwuw0yzjQIkatkuTIdlUtkKJ/W5Xfaq
PEzkpRUOegojjZJxOPjxh4LIPgJV3IZBhBsbFu37Hsrz9/pv2k1XkV02zqGGlcEn
OLivM/33VSkh3LpVcOEK6pZlJkdREErq4HgxSXcmYgEGHNKQk+shXS6ApoYJQrYZ
j5tIvWAfyBchuNcbHHaSrgXRkDSZ6SP+W6PwoasoLlwOcU6qbdqWxDETbS2RT62W
MyVZoITT+KKF2S63jufZ9dJmzvcMdyxndD/wfWnO1IaZ2CXxhj1avwfM0L8zcmYF
txYbHtl5JOpUU9atYDe85XtrWD3lycgdCu+3YgEoQxFEABj1/KLw+/Qk4+mf9png
iGZ74gz3v+oMPrTvckA+j+ZBDWvlVhVwLA3Us6cPI7ximK936CTpnVsdIPpVN6cK
tc6Kgk/cWqbX9FzwxKxRYjNPUfjvG2463Jo+nEPBOY9YqK11NyzwHt4R+W0aGFg3
KzN41ZQxVeauam2OS6ITavtIxRKettfzvxfBwh/ZAuBFRMPNauCqLpqgJ0k8aynY
5KTzp0LzZjw64fzOnlJWDmFfXpV1h8+jCdxoBZuDGNp3CBY+SgmGTulNklGYJyn6
xbae7KnC8dEFzmDYlv5/viP5bCR1nSFXEvA2dxYOnp/OI582C4YMx2EEJHrLo1Tw
FpD0AKiVuZks7gu2iH//J0hvLBIdukHh4Zl2vPfTLV2ESE+fBFWaL4oBImgpPTg5
pkOFoiF4fb4LKZN07soD9DwwP6X9wf9Tv1cZWzgZANsnpinegqsO9chJENXV55s5
JGXkUIRY0NwXrXmbtgUEDW89/90Al77AT1lo94DBAcJDwsgCYxmEeUdfy3yOBIza
iFG+CAbl5EmYn85OVuBBQLx0b+Y1fW1cakN8eHpRMqTRj5kWG0ELjdwwsfG8TM5i
+SiiMRvFruicHB41IUFmNG9K5YLHmHHp915H7ApVPCvqka+yPlZ9DL6td9ErQHo1
1zLOGRQS6A46hh5pYbOjGD3dtP0yiDZLp1qTZis5uBMbLlu19CmZQpKCSC5THiWa
unPLeprFRfcE+dgNYclNUOgkkEI8h4RxxlImQnQRuFT2QH4SV9okPkOxvO2EKkqg
PG7vHbtIKUmni4GnI8Y1YDRL7+ErzXXiDryZH5/OYh+BRYed/a1+A04Nm+iuiRiF
Oegqv+SAqSD0la9/SOlPsp/ix1oTqpuYg+QKM98uuyfyLKhuggnLeFqJDqQUtFrq
5+Nzudup6WquZgJ4aKF6qsLfkwYZts5LSwEH4OpXwNbtm3KRvz1DTYWO0vCOjGPe
egIf5PnP2HiuMhlmu1Xb23UPwpGtEDeidMF7w8cxhSBB3UhfhsAGNaAWXk0EFbU2
ou0ZJWJ8UUV++kofXjSlu4ezRbXCn/t8X9r4NR9+yH+WL7ATCh+o02yDd4Pq1tUw
4DWz1rAsUY8dwkf4d0U60rxrnT2AkvY+4HR0hQzFROf+zkXeJ3vtcykufSEWv4Zz
TqBSgeMpcPrE/kZ7ik1OulMiyzH91AFcdisTBcr1jSIUUDUp0xkDLAW/Bh4njjIP
dYIuzCvyhe5IvWRlbxqlXP6g3HoiJc0xURQ8DJtkodTIAkbsyT2NWrUT9+Fs/AEt
JbM5H18B5/XAny8g4begm00TCAjfZl5k0k/Xy0ZdmWYjS/lc5hR/or8j58mVAG2q
aAgct0aPW0/b5bQVyvRHw+Cff8Eed4DwGfCBAEWMl+EEv9jiImryZcYFC3hV77c3
XmBTZq4fZ9gNph1jHagYvsd0qLkPbBr9Lyh18svAOHFE1/sxYRrxiWaJSK+SEENn
matK2jS3S+XzvmSlUxRFwEifqEYo6vNvWWawBwkUYeU3xUo17nf0LAZIcWjiWayf
p6XiPhzJaBTDPRTxFbh9DISlq5OLvXf6Aj/s5ACehO0xO0hAVS6EpUxXQqO+yjqL
yU5pgrmW8eMHHq85FXHz5Ld3zwCk7YHQr/eNvU9M5mFtbrBE/akeDkeagaGwhnjZ
M+jq4VtQ3RgWOAgpDoK8W3yxKoNGltx8ZaPmZXeF0IUyDRdAuj++EyO7b2Avpr2V
CijnR+4MOn57LFnsB+fjjnprgvNea0qGAmGAc6i5bSW1+qod1E2K7DwAr5/moR4I
+8fqkmpl2Rw2C99KuN0DVHxuhtQ5DpmaRgFMk3h+zj3wNedm9z9ZYFOKW0yxywLb
wi+UZwNWvOP4+OsxO4mtrVdOVJb+Mdd8ry/f1R2AF7dXso8luhzK/su4iK+7MWqz
voi3en+HATTFZ86G9e09FP5MAhxyUbUqwdGql9DIGbrJJXYgJFQPF1j7eUEADh3R
oz7pZOlmifGUgBQHe5deoFKMaG/JzInq0BWpUBazLWQnCmWKiAi5cleaiMxdXuTz
+7iU/g0euYKXthBhkIJEQk8u2JmfkDCikur2EfrS2MS8CvKdVqL1NUGWXNkdGUB4
VcSxS/s5QvFOOLuMXjgcQXQ6eUKseBnfhFKx/V2IKPQsqmb5p3pfpDonG5kwZae/
4UB45BOb9zRxvyaOJ3g7KGrFGTt4A26OXzZCz9ihyHD9EKi9cMT12F3dw60ddUnl
4k69Zq9hwxrS7EtHOTxP/odnaFFiw2WBIaPUTOGtxGAQdX8L5h0CkLUGtenZ2Vv7
cSkX8H8iCCWi34+t/OmxgUh3s606JdrSG4Yp6Bl7TaazR+fw4+UIlsBYR3b5lsWK
nh8eL5BUPR6iUe/gGUF9CqzAuuCzjjJHZnGfJtyTBVwapQ7aw5cWgOgy8SXdMNpx
BtWXrS4buJuzf+GqG6bNCcgNn2F/ActlHPIhgeC5L3ChG3hSxAzH0c5SJd3v5Rft
`protect END_PROTECTED
