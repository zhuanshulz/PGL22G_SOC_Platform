`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0bqjGc5cO5hyzX2Lt7tLMFEKj8OPcrwcycDKXNjkIDXJDGm0xbW9pPwwKLrJw4hS
5vDigPG3akaCsV05t1TB2C9lRdb7aihLErMDRGB1HHV/8TT8RwTwv0NGrSHAf+z6
iJgX1QZGGYt3cmtDrpQbzM4pAoBINUgJeAkOlgKapl4JfTUY7ysVZHeARJHvrW0U
zath/xeMAbeKNwlOz7Ql2XN9qb7WURm8W6/Ms0C5VwJB/1Hhg1OnwJ6Go1teABFa
wHTtnS644vNxPkQeJBYSZI9lqZ2EgCsHfYuFTvtDmO+MgIrCvm+cZHxr75/Ruzkh
NhK1Rg4qsgzWh/9ZtMsejK8Z8sL+BBpqX6VVIw6Zsx9/sJZFBUtrg12KIUL9+SXL
yJskTCx8A2uKcx3UKYt80JQqUn8MqyA/eULpXid2mRzjESyPTscExKl0xKfo/gbx
pa+oaHz81osMscgt2iFoeLjbqslKZS2cfb6pj2s9vPRI762nKsM9tn7VltKaoT9n
773EW0ruKFp/wQvFfTqaX5NKsxnm7d400fr9qMZMoXIz4duQvruEcQIr2HYgiZ5I
W0O/nmRsu3QNsBMoF4+oyD2c80vQYe4A5shD/Gq8BprTrBj58QFCe95wcByJ3OFw
`protect END_PROTECTED
