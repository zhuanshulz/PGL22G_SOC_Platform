library verilog;
use verilog.vl_types.all;
entity INT_LUTMUX4_UDP is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end INT_LUTMUX4_UDP;
