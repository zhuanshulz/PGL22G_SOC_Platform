`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rfddt7+zS+MXgSeTmjqREEtjrDxGw750qKrUmG2TGq+UVjFwFBMmaZWBUXoNAQL1
GYWtZvcWA9/Nso+odJ4zL6sFsP6UkL4I/f9HiPW4GYykGr8zFSrYFWR/V8RQc8X/
GokK3MmY3LdU1V95sHKAXUrZEY0jH6ATrxUXthmGYlW7WBNUYpJBVbMObjTXVCpj
5ekwuhQv5N156Kok/Ui3r8nD6fSEeKG3IDRS33YCfRjtmfcUD2ZzvtNifZe88PzT
DZGEZAadghPRil5ZC0c07p/47X0iyW7n9ICncxXiOsKjVEx8mrmcyoZVjG//aZJd
bDWIBuOs7bgrGrP5lj12v5akOBotjkcEBW4IsI0s2Gieptlvhsnh9tTKeg34FUPI
CDixkno9ClRowWvZLSKGMBy+5poFz/kdVJSZAiIcjpG4KocE3YVOht42qYiJxR34
DkcakqoCUI77XEB4/AwsB37I2sT3M5w0pWtxjqCtxFauCEHdPH24I81VRCIn5R1U
lRguP0kDwA4OtLCYwJ7Ov6Czf105NzoGk7ct/TakYY4N43mM/BAObvdKF88a2fgR
UTFQg21bRKeMxs96OyfFbNkSLUQWIkdx85ybh77T7VEkW3xWjC9JNn32j0Nif/UB
clH3E0ji+u0+4Ib/usHrhHaR9JMPCdVEC97Ce4b2ZYHYE2uFhjwQdWO02qCyzCkn
azLNsRvgOhSUpWK2TF8KIt4IzlRJBZhDxevQk9+l+EmAy3b/N45dkGWxMkJM6irI
V67E7w8gHC5twrSQhedrBrgcGGdSALsG5751Iaf3cqe7ORPs79rmx7eqyIBb6ral
tG1EE6oZ2ghzrwU5gWlOO+vWnRzr2zz63sNk5spxzUBB1QiguIoh/aBNKZDNFQhp
+Do9iNmOe7WriWfUG9IlIjOG+DcOY+Oc2sfGXl9EJQe8Kw3MZkYv2Y3Npe4Irulj
7IBNkm2ZL8hLeYS3bhsWmwL8x0whoStvVk6s3E41pPHa9FKUpBq3CkVcjcwKdEpO
rnaKIoPXdcG7AY/qPUjk0ZcpARSiBm5+SPozGKS0zWJOLcOSrSdO6R3JVW0SnNl2
Tv8PrPetajPPxVGGu1h6peGiWWWQK2sHZgvQ334+FDUtCmmmPxodrythuyxfzV7l
Y/EC8u/oMBlWBLxRmcQNX9bdsNVwZhxPBB9/RjVJ/oVsJF1tGtv80RCg609Y3mKP
KI3uAP47kfiqlv0GHfh1FM/ak7fjP2BTAiMFilVQxY072TZQp/rlzvaOBJUKNt16
ddh4lcULSQuefZIk/JQGPG7CjQjvNf/oUtu9Lj7ivX1pnXcJCpD+osIKHOUCI5sd
iLrXLzLmunoqGfP6LXe9fZ2mSmncvgpHQm8N/zspHtRjWTvChvbo/8UnceGLBXS1
tA9XJvFxPoXLP5nWWTxYPKfBrY+Jghhmnpkp3gQ49Mw001bpjTQVHQXe2rFcnkQo
TmStEqgpgPIDj9wajSW7u9fcqH5A8N8IiRiCHLX405F08P76pvaH0kwC+GGXkG5g
sPitiwkHm6O3bhNseeatkNA6NpKBqH9MiCOa1XD+IOzvCxSPECf7oGnO9QY/L5Y5
q8ozuYKbO6qZ8DSEzWpKCw+X5HsGOEov7otr+HHnpwHzOJTUAxKVv6bkjtb4qk91
v0EqH2DYVPv+X5keMt6M86oyNs6oYKMyFu0jjPqVQbCKy5ZsJhLcLui45Pglt6dW
H1qqq3N7GjP0+El3lHaqjg0bJUc1OLUQL1b1Ni6v0n3cDO7vaimrauqtbo6uFt8Y
fy6m2xzLmsXdxu/bZotq1Aw+6X1yuGy2kscR2fNXeJI71owdkwJlUGfB4pwkt+Dd
//gCFlWd8nHCkupNjLuu4rSv7066J+RL4VfTkLyEjlkZK4HufkTCjfHQxR6WtsYB
7aQvaEl9i7N8Et9utrDNmCjH+N9frfPXP29qEBwTFvadHOren0ZHs6Z6O4KGREzH
AlqwhxuWhhgYbYglKyL+hPvVkqz749dZS4T8lnZGv8+MtgEh3ZDOwaqIopeQwBiU
hHPm3YFRCOdf4iepXHP7MAL0UgBmVgVDbR+uHbRYyAQoVHRFiUuWqfOdAjQXNy/h
psU7zhiz8qOnHtfcR1rgcOLkxIK+xbrseS2e+Ofw6LccJBgSX7OmNqLimy5y3AFM
1vu4qT7YEI+Fi/69ryE4j2JaAgiaH3aDxk5zql7vSOjt1+H5FPKYR2mijZ1F2nQW
tm6CJaXXeDR19c4QhKLjJdh23NB7R0AikrUwv5IARSsDtm2dP5iqpnXl/gylNYBh
TAe67C8NkA6zcLinr179WJVvnl76DF26bfS8BkCgFRPPx6+nIaiHGT4WZulhp0Gf
/BbPS2v5V3wwiRRUtzT39QSQaCb77ePvIo2WvdAIOQS2tGze9lBL9hDpn33aKALp
GS9SKcSBWQtHvdVhkGnZgPntamdgRsyzbMz9yaVtVnmjYjbHwIEQ7khJDR5BHJE/
LJAsJihYeqX0/vaz7HCUWpetxyoHkE/Ev7cdb4B39JdQ82D2+VZB0DWVP07GSI02
7sGaOe91kT+tA8SOD5c07O9SgwJSTAlp6anzYYJqDf1yUz53lI1vq8oLd+TBfONa
QI19GerdfIf0uU4A8mp63oFPjiwA/++5QZUB3Bc4glBSvn/hLsIql8ZJHqNkdHIM
HLZl9Pmw7b88o0RJ5PswvdYezklioRsOG6Jz51NrKz0Y/NeCBx9mJKkv8LlPL87g
OdudfibQItR4Ysk/xVy2ZFmgsnSczU6zLV5N1BDhWkqowqN7zJHOl12kBq1y/Kc5
fYd2xcY86d8GR1InteSTA7pxtpZbEvIwdcmOmVANsN3sJOLODwB6LPyikmwKIvr6
Y35A7UjXfN1LcGWkRZ38nnVf+aFz2p21M0DmVS7yuYYT4xLm2WCvdRyuq7d66nfz
xL4FuL3TWAfsYIRn4l8t9LRD73wASMxM6ZRotj/ztm/ou/7qluXt8x5lfkOe9ctk
khIEuNYRSCl8yuTS/dAjyd38xYXzuR089VFIQmMHJIy9SgJ7nmWQuJpMycxyAe8+
s8Sjw5UAxDOGsNeVic0rY/eiqTuCeEtygnk0t4h5TrPP/B38+OHRJilDVsRUaJUh
5qIqGhhRuo5yZ8eELLQRiIEnsRVpULeGo3wUCAhRa/bzfTfaBHBlcyvm28H9buNa
XlTxntgbOunE5KswBZr3GjfEwfPLVaWjsuDRKtZOJcRLTA5eJgkwK1lrUIqeVR+7
4A0j0TpmGxyfcfTvVcBFeIJEyx+3l5Ep6aejYuPxe5+LExqL9bwPQcImvPRpz0YA
e/8MG7boxVNssfn4pDc/vamRn0Gf+8Ll0kk4WWuWGqyA8hF5PBzsGc5umbwsTCfQ
/G2B94M3yIgJlgI+4h+oaYIsLaaPpfDhqR7yCTfomPK2XUGRGw9b5/TQh+g37u+p
WEXDxkw7SapnToGHJuERJDXJREMO20YJgBVdSjlNrgYiVr17NTZQ3bDenjtN3Ezd
Dwej07Wv409MZiAbaxOOEGcfhGDSSIK+0mPLmeFg95aytbd74ttcnjbwaedYRF6J
zsm4DYgNCo8D7OrUsjrdUXHf1Gi4eyRhLHOnwQioiVXuhhtZrMsej24QmgZGK3+g
zJe5OqZUoCU9uX+ZLUlVK3Ugt8IoNV2qHY2VNlNwErGUIBp5sudayUDm0oeCY0Vj
adBXyonyxod5vaDj9+NkEYbyN1XCClMaXh74UTG2b01vzcODf3uHHnSEEcKJ76UW
zJUztL6YNCL97suS2+J71AE99i6vNC+DvBq9DdW4fmLzbET7LI2EjcIE6CHE6uV7
Fa4oKLG2959BUMvUyvxyGwozTye44+KVGSK6upFjr1D5fZp7oIlbyBlqpRFQFahc
L5xdH0zWrEYMzi7mOzLcyN2G9wlsu179TXh9cuudvgYrPYMQeFX1lmQ/3VLpCHdl
hwCWhU0TkJmFHGoAq52ys+N+uZFsabmM/3TGmRwW6nAsNNyU4noXqE4Ugz6Rgohk
Y0pQynNeDoqgPaw8s3Lcow==
`protect END_PROTECTED
