`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UOsrFWlqxpZldHdtpHdBJiinEPqzUGCz8ZCvbJNrnleqJzdzqZty9HwkqoTbTss7
j0mApyTvDLncV4qUtw1G3Rqvj24NZYOTXzieebk0JUhvda3l4y8FJuxDmCazRh5j
VPKVZCJ7Lk6F3zsGxCj5hhBxECfCc9dk5aMmXjwTGeaaDql+/JsRiwWD949GHoY6
hxKz2PNrmqlRpMa+2khyQZS7tv9nIDspeX/BF6DTLqR47FlA4cLQZvLx6OitDvcn
KLpmI3KBiQmK9nvvByUisqJyWqm97TPcYCkJfEobZ2HH5gYhNydPFbTqBA0YurdP
dVYJvu6GtV6zaRI9ISnftchkFjjW/oSJrP75D23tGb9bjftdBagVtwog4Vh6FUTn
yNrjRHP/E8h4H/4OVnRm43O4sQkHbmS7V0l0DOPM0U26uHiseDCUl3dwjA3VrVqh
cmymvNnSozKuQ63fq1HP2ZFrD1PESR+GZxCmDqGVkNc=
`protect END_PROTECTED
