`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j4rVxC8el8t27VhKWZ7xB3xVa8XIH+rCxp/kcNR2Lg+EUoav0TU4tslw8O9Kx8ys
5WvA2/HuKyhh5m11Hj2GZctO30UcVl7n67l1egzQ4CxG8oIbe+WUKQl7heK3fYfQ
ZldPj6HXcH2u4cSl0xNJrbk1GZ/dK9jwoqPVMgP8sBSaEVo1esByv2KcFl/RZvgh
Ljszes2/RxU4dgsBP0+K0yRX7ltVJ5V9eW51pp8IOVMT5DHGVg98j4iqX/4Kyc30
rDR/62wLx9VOc/HbJmG9Icc3e58Sr42AfT7RsWRaRVk1OugcT8UK6LwJYh/wbUO+
ZLeslgs47YRXJF7UjFrP+AFRR1pzmCqY+MTTbo8zsffGivEl1UcXurgiX8QxvY/n
+fI4KdeSX1qn3RqHN9UIJ+4LgLOyyVRMbTrH0BoSDFisS1rDdbRUpkaNYU/jw5R+
XgbTcSgD2SpBgwvXOGYFtT30jT7pFjJxLJ4Syq3OOKuI7x7BOoafpWa1aZkghk55
jIlWzXHpb4/4nM8Oh4lTsCF0DBaG08hZFmW/FZjeuXM+3aCwKwhwu2NG1ljVDtHk
ImEhPbPxPJCtnRkqhcdPEkP02Gj54RbHXCdPqjcq8Evp9A04WgVE72WFfPSnWPoJ
/SD4wiZF2vwmu0aRejPx7lBN69HcWxRrGBDwZRNZhM7wOvlPXKVZKRFS6XdV05D4
e433uPgelNckElajMXeomHowMy+c1VzHYxpcfUf8Y2kwQSi2v3Zs5jXxgIPxkfLy
mDzmwvL2uiocJUlz0XtK+Q38M86CaAJKiZ+fu95XEa8sW/i6QVa5mmcFcQGo2dQJ
ajoyJc4UeUQZ7enM/eiGpxujXm5LoqrBPafE7Ppt39lPsZgaK05D3TdA922cQXWI
wj9eSKnHAV06ymPQ0XidFg==
`protect END_PROTECTED
