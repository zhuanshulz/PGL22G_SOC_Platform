`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+FS7SkMpXcNpTG4cCmA+buPyECxXrGLf+VPM1lzCCjUuvyH/Dva70wZMRPdyBcEU
V/3cmy8IoVKXWSbP5SPlsWG7jKl8WRcSmlt9/hIJPA9zyvfWQkQPqulrpbCFQgQh
po05pusi+Nc/M41X/IjisZxLMdfsdK8LMWF8+eCUx6oYdGqw78PXPOhm5uZ268S9
5vZ2H4EA+WTY2cBn5x5prNXoAbbOfwTbDI36fh7eSwmUf1OjWJn5zR+tbTR+mUKU
tGLLRmtAobfQAvxw343Xwj21RAMjifp35SLsCtGMsKwAwN/KrU62C8WbZIiRZ8O/
azzFuIz12L9IIsVetEEwxur+mkktvI1mgtzJ2RcV8EJTVd1r2xL0c4u9FtsSsGWz
C60JbNtbkq9QNUeXDrw4Notp0ZcJM3049SW1Sc+DHp6gNkP36Bxjae8VqGsdda0F
arNHTR+9ysKgSLQ1W7YXxp/PQQG90UUxWDlVG3lewsbXQ4hojbfEiPQROcjhZUR2
HW3EZaaPgGV7n2nYcYUa/7gduFi7el1YlbVo9hQTxu7fl54Y2+m2ut9aZZ7XFBu2
sDOEgCEDTgWx8cLanYFgLkLQwScLXiYSOAM3pNBXdmA+PKLKpkr0rnBN/yT+ZCNN
s1p/gpFPk6XAOWpjilrZz6EreiayERXLy2hAlG9HiSFZAgDjiO3/6OUV6RNTOGj8
siH7AVq0C+rlB+673lBE02K6V5Vdq5gb3QYBf8z36sMdvg5gJtKSAZWECaZDj+I4
HlXlTCgUJvsVp8RyTMvHYkr5pf6jgJDs4E8Ns0LiVbCwBSFoi/zIFva7AGA889SN
TX/SCHgJN8Nmn3cLtN01rDD3cOTbkuaGtLWwrP7FAZBmlx9DNOzXrlyVoLhDJQ3R
sm+RMYt4OZnDT5BSTLopoGMnTP7o95T3sjM4jgUZOMTRqCyZgaPRh5wu1366/yLf
aydo6uew1NSuu6UNStNc/aFtKZrlifvL+CiicLu8o4V1mnMJwMnco5DKtXK/Ag79
nJJIOLOaYzTDM162mbuu94cqI8adzUt/bF74TKFvS6Wh6m0vXEVVUE+Xaw6yjJy1
pTZP77SPn+jVViFUtn9s7oPPK9Bpe7nkkG6ltyX65NZuQwAlgfcQ6zG1ouh243Vh
yQxac5THfqROJZmN+jiC2wnUMzXWp+U7PFukkilQOasR6TB1YNl896ZBNqtyICR9
rKrDIpcZ8MZbvBjOsV0Zn6gfzB492o93Sc7bddUCFhdLLz5RCyiBiiGjfsNTe9n+
/YQtWPtKR5hvlUXsxhKOvK/HNo+ZEknQna9XVhNc1CWUhrVhiOecXSJIPARcGc8v
jiA7a7ts7Mb3HY17/St4q2Z3vYuDmXnsu0rj+Vx/znRmHUXtvJIOg8+3tuUVHKI9
qnbaGHxToixjULoC6fODlMPEewNhyEVfwo+VhT6NLRlRIX6G4nno+J3kqMADsnwu
`protect END_PROTECTED
