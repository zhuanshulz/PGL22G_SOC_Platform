`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zVAB66T2saB4L0Cnm24M/9FllT5UYQ56X83bx1REusG1ZOkUci40k7h3FEIP9lya
qmLY25nPTLPML4WKtTHoc4Eq40O9xAqR0SzwV1x4YLwwbpOl3jS0WCTKE+9ENQhv
BV+v2R+d/EfjiNWvzVyJxxVXXyRLmCmimqQ1TCGVNOX83Ew7vfu0oOGVvDAFlpwq
qmqDuMkcwAS87Aj7IlOMDRCZ7OcRG+iTo3BFg3dYLi6E0kW8dmhS68jCBlrbaOHE
T/yERfwBMc58I8RnFQYGsKHMGOIBvPcKhlB2R3VSN4n3EA63edvwEf0dNn6ZV8Kg
ZLICkIiuxPh92PW/QjkMlUZi8eZPPG5Jdo4sn2lsiupWmCMzj0z8fRpGHizgLtO1
wvL2GZbrFpPtIrxaUo3rh3RR9nE7W10ZQXKPkVpBGcuSg2283k/HZfVYF2RhdK6C
+96lxox5tfuh2WNXYRT2XSapGkq6BTYxl9VmDE6S0YyWirw3nJxLR5dehOz2X+Tg
+hDLnY/tDGSACr5HUFrEkAf/r5e8VhugBjKiZRGi5D0yT87k1ZZh6I5DM8atui71
2oGdQvd96PcC/VbO6Jgh+ew3a9urhjdsc3rZa5QySqn134SUh9DQPNV3fD/0Pfxp
RtANzvk0tzZWbHrgdu8YdrYXej6vB++DPTZLLNLayq6QPxONStb1MbdtdQ/HH8qm
BBti08EmLCYAYDJRibZ5fZUkDGDmBM9aTXJjbcDD0G91RM1YKhocnlu32nAugKnM
6dE8X+iQszLSnANtMU29fAOQ9D3Bf6+inUQfNc2WmThlD9X/1LxcpCyJgumwPgJo
arksRVgZ9vLWb6+cLOvbWQOdj9Zt7PTW8A6zAQNBrs8Iir/Jok8SxV4ullfEAepI
gu/vyK4uf+fsWT9GoGygAtgNkWFXfiH5KbJ9bPsjVuKqB28pQdeKZzV1Zs6qZ7oF
Rddk1DZDfRMQHbFw0HLhYbH77AnFUN/TRLe/9Zw6tpGim5xFbTPNT/OxiYPfV/ZG
gy3UJbvj9EVloO++I5DzaZqOZebcLPge/i0h5oocqTGRJb4q4cXr9QVVy7ksPhOj
giYN+qyFltomrJyid/FgRa9yxIOrTUmW8Dzvmxss8UmQL205qu+SMMMjIIdfcabD
/1bEfmLEcBXRyJVtQ4pgQ6gDfaA0WqvoslBxj36y4lJeutXgYaXXATtum4awMttQ
V6ZU6g1YUJvw8rEw9bBoOThKrOvXGb0KtCUHIeCE1xjRGRJVK33RCIdePoAvXv3v
m5teHPOMT802U5EOpDDUEB8oBAdKSmhFonFw1hpqXso3V/MYjzpD2meJ9ubme3Fn
ZpHFB9qfE3vHm397JEepNXGpMeUcrFUPkIU+JVgyNVeGjQfEPQ9ZP9lV1WxQ0de6
6+e49D85VejM9xepW7ZVhUvYkdtgwHEf+QD2eQUdOASb9u+hE6l66PNftFEH9i4r
EGZSwyX8tfhrKB4GmSlgjIokEtZgGNGjlRZd0RAsppUQ7kpv9VctbAMnoeqf1NvV
yyjQBpIDaWeEjhu/FfVkkVbkpv32Ayq1SxtdV66x/2auPQGKEz5nPsftgadHGeB0
8hJqTkIzkPQad45/B/+IzP3rmE1bTGksAgrbKF9c2d9wwd7LR1+rocdR7Nq7P6i8
efBl77tDmzoXPnhHr5rvb3AvdsZny05NAl1nfSCtNPDAGs3yYpAQgsrJRkJX4BHD
`protect END_PROTECTED
