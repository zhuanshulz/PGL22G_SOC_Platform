`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/FxzxwJt52U9/4tpJOz56l3xbZCUybu1rr6R5JmZiKIVMJsHvo3dPY/GQJZbkHZK
4At4DXNRsjfN64c7ccYniTEA1nNFjfJfk7YFIr/knFIMkghuDCxBqNqgLjKpSimB
Phg7CsIPl4eF5xbbG/h1Tvi+vMSN+JySMf3NiDw2b4F2rZCbkQHumPTwEgcjaKg1
P4GpUiEtJiLoOWsgJjLsT0J1eqRomv7whHrqeKtakfr3OzI99hIwTg2qsGWx6+jB
/AzzcZn/7tEmYybFSDZjnGCxPw0nzfvGuFu6rF81Jn1uCOHKYkzOP33xNk5qH1M/
+wdnGXuwYMLT2d1lFcMJAoLUwaPBGkMkB9sXV2fNiD6sqJWpmH88XX8tAlQJy74M
CULTwCCVwOOKTgAMKs1cPlARz2DtzmmNKdtmdHsS51o8dYY/22iW6uuhThL/pErn
pBMfFh5mZaFqxiKTWrlk6FBscyc9VoGYytVMuKX83ySwWEBbjJ8Q7gWnHd0BzeI2
`protect END_PROTECTED
