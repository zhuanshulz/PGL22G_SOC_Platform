`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9HbggrCuxhXEkb8VC3UcLMg2ZBcycVC/z9pfBbUft01VoTw4SmhJ03+86Gq2Sonq
+JjuAwIgzKkXE7hWC5gb4Z91eFB3CEJh0BGTastmHc0OqmmGwaZjoy33cM1bOkd9
xXynjDD4Hf+51ItKWMX2C0/EzQxc6eCQt7kv8ApDHgBoAbq7FPbILorSY/mcy/QH
zUgU8ktxS1VjnEMLhUqzMr937qGRzhY5NGOkeFaV2EzQdejcAfuxb+u2IPgG5Yge
s0Ll9aLtlW9VvGG+i4AiDZxM6OU7sHHqSBTXzCyiDHBuYuZzftSo25Na1y0HaeqS
fqsSntOJobstbv6H1OdYkWsNKaw+Kn8D1AggQbkI1uF8R0nHGn6/LpEIrGMK9hTJ
sew8YOsp40ZhYfz+DDaXVGdQU4+8H9EiTKScMeHfWXBd30UsuIMdMwYq00vFDKWM
Fenf904xpiVBG19Q8RtbEIloB0FHcCeUEUC8o7con9iZxKFwDKLU4NgQUgYBZ/B9
c+dA0ZfUMnOrVzfOilDMTkmlCiSNhxE2zwvvx2Hd40pFqzsJi6kQ3Gx8qHVw5gKP
`protect END_PROTECTED
