`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q50efLITpZRJibWArn5UxpPqXSQo6BeRodBb1ylSqQb53S1fi+lANZEOadnfVXU2
CMUzLO64pG4fOcd6h0hT1LpFNX6RCmsURBr6qssmgoqRfZ6gXpLV5ugld+i0ujvo
LZU+f1qVeKc9PycBXdd7Ov8XZKmRXCxAJmwe+NA5yMBYCbU8dUYJmb1slhlh3wGc
QmmylpaHB/aNmqPL4d5tAMKbprT4RIzK5WafyVdYUVN8atVuadR6ufb65rweEyPL
x3oNwQ0thtzYuFumyJn3eIhr8hFQEObDV4gM//jEp9MUFIM7z5e+epOibuqLLTZz
bsj6sFuaZrVld3FJhOZXzBYAcd0X6sPbvW9y7GA9kwwDpnfWApBOIb/+tGMJQhWX
ciOddEH7Zw6khbFwIlkRanPivD/sT8OmN6ATEJOYcY9A0DslvGaVDeGsjsoKKvKH
zP4+OUEFjK7+6DTJDFVpaXrqtO43YW5jCNZQuq4WmvFH4Ydx/eAljc+zK2/p8rhi
0lDYcfywqbzZX6fZI5invP6dtfu00XBuLgj/Fay1JdyxuPQlqpOVdRZCb4UshaAR
BCbm5ZjLinODP5tIXJY1jo7k4FJxvbXqkFj6sRcAJE+202/bk5zMhlx+32mFwn/x
kWk8xZRdCyd7D4Eku3ID9/etLJGMZz6Qrty5z/PI7rI3kSU2Be4I135VHRZAHe7o
3txx+mgzId/OKmpV7cR4GX1/auHuNChFGuihTiRzBYRHbXlcxYK5cwN9/mYO5Pwv
uOhNvTzRvtsxhHqyd1Upeg==
`protect END_PROTECTED
