`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/NuqKY78m3bktt0b2IB05AD9fo8Dol6U/fIe5P+SbTLtNPeSiAOwdEGbqIZOZ+ee
hrQ+/8bJrfnnqLIS5klNRiRik7gNgONjbkf4nPEiLNGDe9n1FV1sGk3nktdIkbl8
fNP1B9gl5ZksGOT/XhIBTMPClfj+/G8dl1Ba+TJVYS36ADuiYjGtuIRpPO+kte6u
dB2KHDU38jNYLL0Kx4DWiLrZWE+IFr10e06VtedwGN5me9yFrb4HgObt/iQ5Wy7T
ka7SAqmj4L+5YTql4JnHaaEmsCOfy577XmZ6KaTg8WvdGdihDYsFEwajGHWUOUzH
m2biDam4vWD4c40vXLhDhF1j9s8039mKCy9T+kT6LIpq4faTXZfR1IdAxQ4JTj8x
uGgNzc+S8H9ePQVbzPIo1u4cMKbk7xz1E/bHaO8anpk=
`protect END_PROTECTED
