`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yeNvRXTmYr332dGQ3fMIPaqveR4G3Q1yK+ecB3x7y2KwgP9OFi9IvDpdhnREEc2d
G4rfRpQGhkwFMU3a6Y/PW1+3+ypUq5iDdiKkYOtvdLHibegIXo0VtnYsmzUorSe+
XjF4JQKk1DqzdaIdS7cBfoRfs0nMaiHX0Gic8Fz4JHJXKNtVmsa8tDr/XuRie/G0
Wp5tP7UK+iS74jU+rPxZNB754ksdZmgNTYRM+L31fmMHKNdJt3bjiXPUwVWUAAlW
aUbVXCGQ4FqMh1Sai99Kp2Gx9HE8oeKIy+8Jads6LuAOVUvxpKCXW9izRnyefPs9
p01tE9Cvl0UHMBYEp5U7pnTgVo1nC0MTqAOEgbV/b1+RvDzrJyIBts09GInZDune
5RWowzdgoQH0s88Khc2LKjzoMpNXYmcoQOP+KfIEJKuuwXndsK/dtNX5WfLtqsC7
gf76qPpt/i2c8y2YhtU9IUVnQMNzrqH83jMGHt2uO3fir0U3VIsY61iBPymf+qoO
U8/+6VRHRnEKQ2ik8FvLv/uUtVdl3hTXkv6W1GqDTESNIbRS4BoRUImOf50Pph+Y
RE+ECfjOWgMwE8B09OCpn+vJqxvttzz6QYKXXdWMDr10VCUTudmZ32EYCc/0u9oq
`protect END_PROTECTED
