`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HdvQhK5ObkGga8NEWoeKF5rqpQPVnkH7857H74RKH7PJpWIOKVgXGqxsRXIai47t
8RImcdl/PDfQrjTgLwrFqGDPac0W9ibnEefMWngE4QXBOPdK8K4En7Drne0um8LF
TKWCXWRMPXeKsvLRQ4zdfEBOQMmf/moMCALQ+EXrNWtwD5eqYKcQ/bNrm1YbJTYG
J1MfLiE5tSjZI0nEii8Yl86dUcveqM7iTH8dWrexJUfGmc+SIT7/YxJRDmE8gbSV
3o1vFdwLKuM8v5RIOd/0tfUq1NKeaVLHJlVTmpvU4XeTbkR1YMMZX7gyH2tklOPa
xXsFXYU8ddEaCiUpgiJccztkosTg3uCVP3rEk5y4uqwAAaexfsxLaSg07wPYd20I
nxTsgRcc02N54Dr+K6RLClHxAgtLtvhuEl/yR0TJs+/lG5Kmxo5gr3h1dLKm3Qf9
54WVfqmtof0wLNkqtu8vkQ==
`protect END_PROTECTED
