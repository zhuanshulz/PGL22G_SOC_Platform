`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2W4bc6EGH6ddtpqCTDez/tQy5HtziwxUGuYSmexHCY16Z52BJPXg2OLDin5x12lg
wg7Hoo/Nyx3zmbgzq6st9JkikwSNtFlrHZZ2/41M7IUY4L1xB3Kh3S49vVE3ahXZ
gkaj+ErhvesbBy53/wUvcBg9PVsKbxzyefleh27wmvJDuJocuYxn0fQQwnRrp4/O
X580GZzSjxTSlunSRE8ZOMOE/ig/MnI0YSz7v3P6bFYy+s2rQA5fvYGLwxtIGvkQ
zpr8IAY5S/gGsJL0FM73evzkyNOYIEwhmRS3uVP43b8S5q19YrGL7lF7+3Tqz14K
AO4/RAKn09ez7343vNq0mN8dFG1msFXJB3bAwg8HQqyzULt+Zu7J2+q6zswpV9s9
7th2Wnz2HeSqg5dkaAxNd8yKtusu3K1LQdO80MQ5O6uH4xqhgMtBk43lvsFOXfxc
9RBLeQSfM3pZk0EdIrGeM5wxaaOVVDrlzAyzLTYfS/qMGS/RZY+soGhiK0Swphic
eaCDyF0V5AclpZWt8W6+4C4a+mESDRMCcgJR6Zp/qiNmUfByzTIVjrggtu2cRhfV
NK0daILL01lbPNWTvsDfcv+oPq8/+3LxOyOBra5WJcWDBuw1LuD9v11Xjsuc64be
yk10z03ZGIut1Y1pHlIybrxvI+Od4dw7N0lMX3y/U28XCtu+11zEtEtPiWcyUVrp
ThF2oEyCb2RWiB1MySuk4R5e3v1VzaenaO0MqFxJyR3Jq1+SgA6+K3auadQElFT2
pZHSIXkDkdm7ZXGLGXjY51LabdAiC8snJXgL71RlZvg/ctASPMhZhQLFq10+ZzNT
4Ybiemrp0mdh27J7W7C+qYUkR3cHHBtlORgbf/A9I4a5NCziqIKjPly93+ZxgS8Z
sDlhjP6ImjOLOE5oxDGKdViXAZYxWoNqBFnM5ozXFweeX+Ix7xinEB2mwax/VQcl
nMxz1rXmv8zFtPNsu1DZJ1iiZkG4YIw0SvSoXYUNvA+qZaZtmnxiQy+cspYT2fgB
18x+pBBFwS5DtcbBX7q9VeB7XNC8kBLjwBf7oxBrmiNENQYZX67+H4p0qhmT4iZF
P+E67FIz9H03eWXWZafL/DIkyT0knUaYI1JXvCa1/7XB3xh2CJwzMHjm3KulxHnx
4P7leQMu/zgMym25dz7YmcWOW4fwBEZXZpD+aEAWZ7GG/m10mOwEN9X+tMxUbkn+
JVd2kDsEMNaXWWuN1D2r2luY4Ol0D5LFhLWHUtdgJS0QRcgO5/y1gGbBkCaZwKVY
5QTttrMvWhA+De2SXrqMz7j5NAhBO0y7vreCnoq4EIIVXeLwRRO4T3Xonl4LOCN8
CsbNX+7jsc1451HY0cwYydz4asGDDXxyfXI7+qX/pdeNKZTy+oV2CAklYnpZSvhX
s7/3etdNiEZPfeBABY49pNGPaD4ZJq99mOOUthOKRBAwmHla/PT9dGKAJRkxccNX
Jp89xLcK5zk6wCOuEsMd7EJZH+IUvklFFeNkUoXuqOtOojiWA8lbyOVKNliI1426
CTd34fTYkt5cvPwoNuH3DjkC3sIfgtm5w6sWRIAnEtwHxAcqyPMngQIrx7giOoba
DyzS38I15PXBOuY+skU9z2pKIcGNZM43jdckwV8nbnpufMVgkPPE+9FUHGUD0GcW
qq9xXPGLpJ9ocWdDysQDMORTqJ5LoP16N/OopIUQi+ShLE+2ww6dguT/REPDJcru
xnKApuycRKlxyAIl3vk2fbESIQxVEEaL2C236uI0Dtx82ze1H3Lg3VbwS0UNtMi3
qwxNDREjuYn8wjfl21+wAwFVYVfSjwqfjJJx7fbyLrzuafeMAHaK89iQ8NOgWldz
gkYvbQXOOy2PW5kwlWvSB5cCozmo+moQbVUAHu0tOEk=
`protect END_PROTECTED
