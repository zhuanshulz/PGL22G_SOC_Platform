`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z6rFV7M+Y5cGlluuI7XJlraDYVj524oxYAHLZyH+Mp2yQw5d42wqyreVawCIz9aI
+lW4OU6APXRWD6uluGwUcd13O6URLhqV5WXZRPljchCpc9/koyvnQPOokEP4zyIN
EwD/Tz+DtutwAhajgk/mHxUkZtxaTRhpLVvTNFihE4HIPFwIyQMLhyoBTOiDiGm/
xg8TmxWVGoU35EYDQzqVHkQfhH9byqQ2JDSFP6l1r87a1OOwSA9dxi6qOJ2NktnB
vPCkyEvpj5aK+hfP/Rb9hhOgA+IYR63ayvrSDptiiXwF9Q3c5jz3FyPTT9Hnd+Up
fydpGcvyrvwnWyo/gKL56oxGU41jWApYeS3ViT0TEEgf0C+4b7stc92zYhpwsBX8
tU/5P88Af9bTSUDv9BMUbD4zsEuP+C6kg6ki8WpTx6us3QxKYRDic2tzOLupL98m
Fbwh0rln4hqbcs6Ixo9jr6d5LH15Os1rn4FCKr3+hcaWWBrbLQXtS6TBiM28zbif
BYIalZ/AVEAsG7qMDnXetoZiyQLAL2BfA4yd56ukrBkLSHoyUoM+vTRR/hLwB737
YuVoamVvLO8M1ssOOzLnwZnZcwdXrripHb32oqs8udo4wjtnM1dqpAEITE4fXaPO
+zciVFzbOt7zQHjmKe7X2FrExWMT8ve+9QR3ITbc5EqaXIPIRNE2FS5DfHChWHje
v7RJ9WEdXECfjNma9DoIOBNNc5qTOK9qaP61QrJ7oE3Ii/cWmO4fGHk2x4ktNyDb
`protect END_PROTECTED
