`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CZGCEJgJC20p66aboRepvXyAZXB1kEQKsXivx4nVn1jOK2UbSdfLrMYAhjbhNtKs
Iu2jEU18UmgG/Y+dVgHs8QwpitzjUVoCCMIaXEIfAMpq7Co1kDRGbq/ui8X42M8b
tLpAvDbZXtvva9BoroJQn4lyT63y/g1s6x0QpmIRNkztfmCv2P93LAjzMbBTuuPl
2gaDNm89H4mwd4IyiylMdHwVuy77BdyAmZmARWnmslgQmDJ+Ahk6rMpFHNUJ76F4
t5meBt6p/ToiSUZbQv2GD5ResMRvK79n5yhPWlLt0G5FgCPasEjNlQT189WLmFsF
XIvysVlvNa7KdwjuZuyUVeNGSFOPeZmsWUW3yRTP340VfVVj2VGpvtS2aNURpv62
50rwEh74uTfS+1iDlKSuENJz0viaw66GLm+C/dtwAoDJR7GVmA0PkOWtBmwSRHL9
ulbNE+54lair4bJKn/wtLoi7At2JijyzOs7znpJz9zSraLW7S2cFY9aExi4K0bgC
7urZPcritlHi1MPzgMM2Ye5BeIfGiMSkvfuPJyjAICKqIv8jGbeWX9cGYo01wUT2
/Fc1mP/F100VBlv0vWuYh+DJoAlIZLk0GmTCkg0da2nGuazah0LCSecpAtI1lBW4
ZlxC2K0Wo5VIQh+AFi8Te5vLLWLci8Rw96duEvA8U0Bctuuq8fL4ZKnZIBNa5NH9
EyVJyaqhqu2rEPZ5ITAFwg==
`protect END_PROTECTED
