`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hH6g22Hegz6EKA3SNQlCKqmDFa/rugonOxjDRyMs7SQ8PkceGt4OD3A43kXO1pji
CP3s1H2t041QrKer7+Q8TORuCSEbgHwSP0UsVxHj5ZTpwcbdcb5ODjiv5lfCm22a
Omne5Y3+78HhNPT2/IvKzpfJWEOlenwYbU3RugLBRfIHReX5w0ZyB4nEDNw2SOIy
FZGwfC2q42w9X20D+He/ch9aIoruQZUNsSRBLfhakWRTYM79to+90aMiOTpSMxtr
A4YciNtiMClQwncoaqucaWBZF9YWgEMo5gdRUdTDD696sJDoJKTGA77jSmG4IDM3
YbqSFTRp3dEZMiwixi4Ak8r9717bnbYYsaf4eudmVSa32FUeEceau/QeoMOTe/Hu
X/RV4Em8Vqes9+J0TwGXf74dPLEBsrxhDZMXJmnq/XjZNUSDXKLMnoun1dSJHgji
Ob79rtLuL/+tpHC+UJ+elEEuchkW/kvkeTE0GangmQIB8yDKu29GhwMWpGcomAEV
d8E1eYCpyscCNapVln8v0643Nn6TimNf48SoKdIXbAE=
`protect END_PROTECTED
