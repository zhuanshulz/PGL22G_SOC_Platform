`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aJF375OcX73Pcon3TTBzZLu/18fCbpK2GmC1YI9a2G6fPlpiNkmdxLa3ljq/Wx2i
8OEbwcFULMk3meeGvMbsxCPkCHwijD+CXQBFPem6GisGD53htNc/Ue9oVCpGUl0H
0hcAMSNjlm7ooRrgJctVbYgEJvyThUF8B3p7ILQEJeYN5AWa39MLoATmp96NAJEC
1dqf6Grd3d/oWnmxoT8WzSCFsSccJ2pshKoDW3RnfUBQykD7C0JdSpmgGNYSw3AD
bdY16S7xdmjCWpWcfYmXC2zTaE/Dmi8yBoPEkLLDOBymIfET8EY9p/2rPgROOT8y
cYTKWCkTLyAKL9goCvz6MXAmAcMrCGH1ilzeU3hY91N3hcCtzkK6ur6ZaPlbO2uc
dLWBfchVIaiKaUQTr7FidrtuF5wzZ4zBGDaJ5dkcVkSvyN4A+AAkUUsIYTmj2tHU
lAgJSgMdD0vcPX0bFDHXrBYlHB9xXNgZFh7awQd/guXBzhNhce7bZKWKvIhxjCsv
LL9J3sddtdNyblb3lwYZkamfKcztwSzrIBREeiaYfX6E8xq0jM2jkh8LgjjnlcRV
evOL9RqMpbYVHHwc93nCqPbZFkeJ24ZRId1FRwwCMSMV0G/6y9X3gB+Beh3NoalO
gHKhlZ8RXT4Ne1ilOuZazXo1BdXA4Cing/Lr1Hd02C9iHaBm2XOPhzxJa1MqSAfS
ts2589gEI+NyMPTgsZ56tkbfO8FQ6U2xpdSfoQJGXwNxwO2JuDxul4rYYy/fhgNh
MCajWUoajXgW87eMRYSXwFOzjxahoPaAYOG66gdIZ8PHGQveTwCw8zMfQZJczDAr
gH+EvjNeFExPpvkcHZ3PyII+USYMlCpOFg0fNizGYEDKhc9LiVIlLGdqQUbir2Kp
AcMnJvijiczN2cw/bdGGNfzfLauj/w83AsqAQm5uUSAXA2fHxGU8c6jkbZ35mzLU
nGT9uu3U/4T1dTLVYVN7vn+JsGGaJHK6oMyzxsbhaRI=
`protect END_PROTECTED
