`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XN/T+cMxiDqq9MTUK7s6TPZPDSO8+ixulXFSgZxa8+tgIjMVFKoE0WvHPt7YJdnS
xQMJR/OVkyA9n2sihLcpzz31nkeWS1/sOMKR41IDzYcAdNm9a6kmaYsEiSrPU1qg
LUDR9ZOuYNwV2TTeukc7DCMJsVy8fjQuFjO+blOjNVeanhDuD3w4/M8P2xyJFxAq
zvICUZRIRo6ltb/TLpV0lbtaiCnt4muv8iVXbRC/ShzjbygxqSQl+TU0Uu+oyk+B
VfIqjU8K2RBfOL/cgdl680XXncm2BJsjlvAE5yl3RFPyDMslutpqEQT/z6vqIlxv
PflwsP86jPTVq8ISYxdSw0BM7OrxmuEpcjEaH7Ex+IrQ2sUW3k2oMzI/zg1dRb3q
zgbeK8C1vphZcrLCvTNPzIVgA4YEJHsYiji1BPv33EtXL2tYUK2NGB+IEtO37sBP
eZbwzH2cfrPJ+ERKOZeBxxSWjk2jR7+xFEmcTvncm+rAAwe0wcvUqclfRvGexFv3
eMfxQASv0SQ9FwV/5ZEwVAr5Qx0HGMgwLzlrrFS5L4YM+UFWtYzOduwVOc8wP0w4
JFf3OldVRI49N56de/mUSNzfe1NcDE81xNaDkb9IAGZw94Dzxv5OKweGgKxcOWw1
6rz6CdR2DPn6AVe1MCgFDOec3zdkZ7t4ItWFWUgMCMkgwRmoz+kMnF1UKTHVE/wK
HcCRQAvmYiqOdyMyVcCSmJpMD1F9Xp9Tb3vP56JihDaYZf7XAEGWtc1mtsi/6vE+
88kCnTXrFaUUlXKYUVFIISNquEOsF8ci4TewJtFfvat4XTCR/wqspKC9WJW3PaZN
7Uo5DZm7Dt9qjle6x+5hwDhlU2ExcKBGdSjEyK8FnAEi+vACVeGlTXvWu1javP1I
xJLxz2Oity9hFRS0ErNLyRf5JchUIbPsH6SNbwmFrcRBBobLBAoXL6onYcRS4KrG
xcU4WHDAnjYV767sjh5weCB92KhK46VTRlXvSIKJ0vuEWIx7idF6zIUcQTHPAIzL
ZlhSesrFrBipXCaYxHr6ebkmJrUp9q3+/m5zTpUtPm4I3ZKWQWHBYO55DnmsvM1a
VH2456974D8HnrpuKm8qEtvsntmNjxNyiK3la/14IWpUhu84MHiLDg74VMsvSm1C
4QKiEzy/gMUrHDTzptmBJGffRXcBt6jrtQK3sJ9yu9aLGh6mQUCDttAftbOkLl6A
eCNsdQCQTekPbaEklqe+pbudhPTIMtXlbBdMAsNQefqW/yrZoUtw7mMVqsS4ws1A
adsI7ssoIu05696EZ+tbV9CScNSZJLEVJHp+LbVK4kYCodQl3aKgtm8Gi+2/fOlj
`protect END_PROTECTED
