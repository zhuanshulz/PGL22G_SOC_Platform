`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PD9c9PYD55s4uHDLcVwfqDHka8GxbVKdvNVB0NyW6rhBeoQdawLNzGZe2eM3slKO
+UFywTKgptKVDYv3i6jpNP0nMgZViVi1x4ynsUMbGZY5NeVPR/EJeZFc54/z7vKe
vT0KK7wl8ZMXqrgfBb3K+ZA2OEvo1jIyilDzxmIJcx8YosOTIUGEHEEqsIF5MO0e
ewiTZvzSRYrn+N9Yu3GMWmh8jnfiO2hOoSn7FZ2y4ruhjWGZc/rw5h3kaRY78UFy
Z99vs6iZZb1eNocFN39pmS2ZVTSyIT6tR38KwEpBI55Iq62+F5BjEuTIkLmwvdKt
6RwTbBnruC5lRg+2bSQlECyhDqy/7Z5pWnukDnaLG1lY3XlWXV0jKlBbxLQ3gISk
d+j1Jev84UrQAx9+FARqncdXu8M4zLglFz/Ayta1O8gPjl50eKnQXebf2d6VJSLJ
mwDrcPt+v8RdFgMWQDIJpOJAEIKeR+HnqQhJu4Po5hUZGojsLA9dZQUqYyxqa5JS
h2Btt/5fL9RfHMS1AX8ETMU4se7nL8T55voUoCTnRodho5JAEfva0mM1kMz24f/X
ozEAJuMEnzJBAKacBvbh+A==
`protect END_PROTECTED
