`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5W69r0Qn2C7eZiz2UK52QzpXqQf5q6h7cxIKqZvu+mLAURQ7vO1InuczV+ZG9vPy
XCaLG6DqDggFu8kStomg/uPH/wxYQXx7EFQPEtJF+OUyuL1ylNs47b3aR05Pbl8k
8PSfOJ1WQ6MFN+wo3VXXuY/S6oRckoTE9hgC8Rz3O8MvF0yVB1NIp1cHpFsGS2YA
UfsfCQk/aaYB/Q1cI8BUGKSF3KaNnxoWW2mcD3Vo9Ix2gP4PJlLrhPhwmLv1Ao+y
DwXS2kmUrAOfAC2eFtY3rmbHWTQTztP045+lVjiyIIuOIaVt34w4pQTYUqxwLbY8
z3NzM5Jz7nenLacVaiFgfHe/J4xqTX8EHiDwDt6vlrbe8Fa2WXVeXB17JqKBU8T5
DtY8DwwBpaA0DvJBiZOateU8j0sKdklkKvYRvbYn62zYkftacRyqKl10Vapfw3s2
1ArzYJDUoWZpo7zK+NDxr+RKvPbBQBRUVNdO6wefeZdjPQZ5IWJD8MRRTfnxJSd/
xMUnOIeiZd1Lbed2XeGcMbynfIhxdkMsmEV5ZqRc3DNwmJs3mfmShTYbJSaUm+ww
Xlo1xhUHrQpGkBYqOf+XD4xueeO3VPqce/stm8OAoHG30QA0Lq1im0QZdFMQTAYs
lRMUBn4IA0vulN5TbVdIJii1FGattdV3rTBTXBYWLLeefygKeRRC8v6IhrwNmwT3
vY+srG23mtZnyAxnHDEOuFqjirIOQuCrthc+Dc34kifvvAw1RYpDpt+31aiTG6OB
o1aOMmPLRvXtAaUyVT2u3SJa2uM9flrPq+tpJOqZUFg704YfOJ/YoxxTbrFHUQ1p
QV9enqOcWJ09bXWNLwZ25KIBB2iVEMCd56zAlqaCJBj1WCZwQndIDDrlktI1MviT
Qf3qhlcUBTNXRN8Ueo8BpX1OQ6+Mnn/hRVRAG9F8J7flbUE0/Xk0hMM5cMeH8OgH
Jx1gQHMWV2fFg7CAZWFXew+a5QIQacU0GX4S2K59hPjtBL8UjqYN4DZ8u9VdWEdZ
Tec82f2ccLJ3R6izY5OrPEDyM/v30lysAWU4I9Crf0xSCs4sDuG0KelHTBtFLCDQ
ef7wBEP+bierievdZQtHoQ6z76UG5bLsHehTYUDQM5Z8xhZhrxfEnJE3QYnJP/cv
JujqGnUiUVOnFJk2lG+Ovne/KyBXHfE1QGPwBF/OEw7ZcaRNGiFgoD2lQD8P+Jug
WKxTvVMRSxzuZmU79iN5/kg6nLvmgkcVy84OvOpc8Z8VJUrVHQGt0hPRmWPa279B
Qi+YWzmlN34LVzzTQbcolZgI++t20L2XgmXK+VJ+bOBRMZlCLd/xmrZYddJ99z88
OhwX+hFeHZY7xIl22KGOW29ePlAm+7t8bBfCq5VRORhyOwCbXje0KqAFcKT9ZIA2
07OrncyQ5fqo9LDscq1vnLSeL3xTclJwYKJJSjSIkw6SvIMDcy9ipTNvLCr636Yy
v2ichzZbX2evj/ktKbHHKbkmjfyRVFFRJbHyXDxorntqioM+WIPOfAwyFfB6s7sv
3U9VlKDLg/TkoPLRh6SOeVEKjjNVNXA4JvOr5cq/3t1A715WqtZ0FHpwuQSaz59i
ieYX2BEaIExHmqMENtKC5GoroboAwdifCRbvBWXzO7ehPcwRJsT5gwVct+6DIbFF
3vsd0LRR25XBVutag51w7k/9GU7Lxt368J4V0aranIbpHj9/vCyP3raD0+QYkO9q
FWZ+X/1elTjKCKcxwYnh+R2sCHoKr9PN5E68/WQZIKmAUva+6d5bmnRKTUi9NhMM
VWTDxwJmzEoFnH3cfSZorjMo8rAHl0MZ84wpxPssuZ/cUW+sbzBiRwbzfalrN/I1
U1csKuxAgN6H4BSV4vcbGlrZyIlc5RccNptf89ec/+nyTNzsddXSjEVw+PU5uUX1
lb5/UAtHO0SnouQT5MSJoYN7Yilqyd99lvA4TlbeTsipcM7v9gpdzVaNC511BrEl
hw30pcBi3G17LG1k90NQLTAVd7nfmWrJP4yVngZ0Dqin7HeKDaYtdDCkLU9ve9dc
69a2JW95jOnBJA6cjPlty1J8cfI69ncylSByBlK4wonTJzgKKcu/J9vSqKWqPH+8
F8mUI31n8PN9IhkU5hstuW8HIuPzOhu3oYJPvnipyf2O6nG/prMz3+ZrsFEsBnoe
LItPLRAbdZD2fms1nkXU+7ueBfN4I5IYVkAdGzeXgmucexhuA1wGBFOcgbohlcMq
oUSqBsjhCvZLuTEf5KWknnDaoX99c5qg0oD4cL/AoXxSAxUFwHmMzkw5FvPjBG7J
hifGKhWzQOep9kanHkxUFIP05QKA3K64oikNDEpl5WheBKp+Xuu+jOO6XpuLoVCx
yc049+4mB2cHKUo4l88sfNJTZZKRTTabIlole97jveKwayCxPiipqDrHy6ABeH3p
+vOMSZUipP6+a7O7tmSA2UcP8XzVj0UTxRwglS+w12BJuN5Onh4G8QpTqya7urpM
A7nc7ooZAPyIznwViZdF/Ljh6GEH1a6zu4Xn1HgGq5zroMu3MpWqSz9BQ2t5f63n
zanwVp3wO8tijKzSoC/NUWd2XMQul3Diii/dP/BHy4ODryxb9df16pQfd1AODOlC
CpTuxgKwt/TdOF7wSAp0/acIu3sBPiAd5fiGuvme/eIKpoYarDOS1e9h3/8xon1t
KOa5xDsRji53GkFbfKeDu/T0QyFsu6AcVvDLXk12g4HMQzTtjtosbk3l2NgTRvHL
vQkKOy7A2hf/C4d1Pp3g6tD7SIiJfCsAEjwJILP0+2P6MpYyDRyFGTF2hnggQ2dn
4wAmJ9s0NVq5T5GKAAXnLimSjWZdi+iuW5eoc64NcHZmXXIuaR8b22NeFgV9bNyY
ozfzp2GWdUYO6qHSFmdLmNY95SkajhEzIzZM3JBPJEc2neJ7SURnLvx2FFqezQ3/
`protect END_PROTECTED
