`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0CvycNNtiKtC09ZGKL+DHph8hwMNEGLkpf5++jE6SFD4MYy4ePWGQOF10/ZDp/IQ
3l6XMykohY/EsyybLJMkkcNuZpOvkI9B9uJ9hiZZ7GGySdYk0Mz7TpYE/n0Qg4Cy
Hb9F7VLzRlYi77/ekLys97P5aL1AwhN4LI9rY18t39lIUGmFws+Xrm+Oq6SXKMw/
RSQyeoJ321kUBb1ko5wG2cJ1zBvEcYTDJvEB5WQ5kdU3i3z9F9Aq9Lm6IpJswez2
jeWaCQV6pvUQKIgLDK/40eaMTU39YXFVMfPLHjYD1Z3UxG9LMqNkSLSeHEt9ZOf+
iPWM1aybfh/79luZmOY8IGDklGJ+lXcH+OBeGSOket9yqKNegnBdyZbCdAqIQA/o
M9YLpO9MV2d2IpWcVi5lBI/dDgGRjOpZLAbMPigd3THBTN3gyZEdNvHMnPBnLOlV
h87tH6Jj45WKzRdSdNQKMRav/fDDoTc8CLlsQ4acgZi9T6LrSnlCCaDN6i7bXWVm
84euLU4MvkdoyY3gJBtFytv7HmKl10hmEWVtS41JDx6Xdv4W55XBJjCg36HcWFQy
GcTSBqavQuF5H6sw1SxZkRKHSzh6+YFyb3kt59u/kXbupVO+yIF/UTVqAfBMs1d1
AbbrTHXYZZfXKrbOHgRSQcqIbcBKH+753k1hmD1HQcQAKg1T7KrzCSBKYZCQ49MY
/XC+tPZJMAz8ZDuwU+MUG0BKI2CCAqMs+eV0V1tVltMgZ7uacVF9Mm8wT/QF3nyO
Cmh3aqNmQBEZkwp4n8FsUz8VKx5YxiUlF+DIwvulm+e44YtI1jNKn9deNMzNsvms
c4y0FHwg1ieUaveUV2/TvWsrh1zrvVr/ULzaRGnWSdWNAVgkb7sWZaasiSIkaRFl
e+ZTf+qxBnYiUMUfVVvU00zrgunAFZPfqQNikB2fM3oEl4zm6ltudSJnaApCGgUb
0FNuShqhL2uZBxf5GMjpJ1Ei16cCoba3+bLEZ8NhhL9o8/uqfZwzcK9rgL8YydEa
EWxjM54llrIrOkt0LCkxC4k4ZRV4tR7NDV+a4eRCbXpWLwIbId7uFFrj7wgs+7Ri
IDSeWXN2ZWGsOLmbNZXj79Nnw9XumGu00XpsCJWrL2oWjTkGN0z/WZytInUr/AS8
XrukRwZAHKZT8WfD9KxRaM8TG3BU0/aLtbHe8menUptani0EyiGRPZi/JkF+9N6r
6Qb5tp6zHGJvFcXv2tIyS1DsoiiOfs0dmQ0yOnWLHXsnmpEyVrtNPRGfjlBN/oR4
SUZuRnYks4+2nKf+BM2mx8Vnzex7KvHVhPBbGR9dccc=
`protect END_PROTECTED
