`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i6imGmcR+uk8CJahDN7/KMiUpRgCjc/Hhqa1KcQPUVxcBn5ViQQGa847Mee3CrjN
zBuWP4BPxhSA5vgDQdik+7ddMSEqt8FgW0a2F4GlC2rDq4HDJ+Seng4FfMBPF7t/
vjveLoDEwNXpRJFLTkRo29pfVpyr3CLk0j/ytqGh3Fjtv2ssLohpFhrALGyujLwh
RPFJUDBGK+PK2DDxL8amrpITZHU0mF8ebhRaIvvphOZp9fOozvtbd3KS+hSUAuad
dNFwU2MbjTRJO/6Pw6Ckaky6kOpWZPm10ihGjtBl0Y73KGxS0hjeAYvHeoWUsKWY
rA/MMNiAEydakYOcJjGIWro3VytVfu27iMl03rMaNXKe2z3h/OUJZDjztoOhxXgE
YhzzjI0rf/zJWWFf4/mlaATn8wD4gwdpDKT+uWO05f0pi4m+eocLbTba5pjqlyEY
Ox7WQF42baqYr2eLcvbAeAfXlqQI7F0M2kuWr57K4c1vjGAfEJ5qfFFb+elb0yo3
UgP2LFr2gwhBDMW+ixIfE20XPrSS7NNbHSZtZ/gfVfRgfFD5zkT6MCHHdMtQ+F3E
7A64YeYZ88S1PB17OEZZBdlFuxo1Kucw+jX9diZAeX5QWt/V2FeupPZl0m4xCuW5
2NoGAcf5fwMfsDJ3A28owt0y9Ds5ZE+Q62EfDV3EvkGLrKfiFaW1WWmpnbbBsxWl
yUPbnQj3rFCyBdbluzILJXvy//nS3wtvrcYQvA4tqmSlQx+6n2bKEH1tptgbW0aI
Cau+QDAhPaq7g5YOwKzfRw==
`protect END_PROTECTED
