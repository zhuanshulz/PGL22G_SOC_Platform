`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wkRWP8A48aly+4fNJ6W2n70EisZf04m26WBeNxVk/M9o5+lQHNTPqJQ59tvroNnL
Xmax9Su03Ktzir/rJYBInuJMNRpZ3GKIfA/WcGvhE5ctWqxY8G6749TDMJmv+/Vc
mI/JbH/5SrfrjAc6IzF1B+3Ji1f71frfVINXTUDDXmBVNiWhD6bZACzvCcsggdNR
qF3CWSTuGl+Xi9wEFpuUblDD4zC65vQNmyY5IlKqKmxiqLtu0e1xOCv50HSU8YOi
72FV/aWe4BewbYokp6JPCyMCa91VlygP7NQ7rKKcUvk3RHGOuZbLGTsXcPd3USQs
Zd7GwUi3jhE4MBXIRkkwMokEnmdKJuo9oyQwNaBXwAH9XjRLhpD5L4vQ7r1wV8TI
h3p32d0FSunYwXBEacErqK1KU1llIoSDNmFYoOxsdlmSZ2pc4GIfgG2zb5gwGBi7
BWxPuOsEN9HkYqFXtgb3FD3yu8/xCQHsxNxXSdq7SxdDJ7JZBYaMT5RKvW8IDlU+
y5u18R2V0/QKw3kMQP+fWeWUTa+LHyXyuSM+YW8BfaxkB9L+3nRMX4qtTig/csfk
8Dw7jX7p2oPcWGjypesT1Sfj1shkwZlMpBw1AXxva5/6BBLAGXR5joJnBubje7hP
xbr/drHp4UbbAKAsyjafrbLfPkOQKVtqGxMRLMVIOZK6Vr/ib3XmOeGKrtdpqb8l
1UEGJ4TVxQeXcKJ+IMoVztogoKFuRQfI0UKUQRXRrec=
`protect END_PROTECTED
