`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eZrgllP5kkFm0gU2XAWWIj759Dhg0/W8tDZ8hPfKVCHR8NY0xaAtavq5BjK58lz/
pH5l7YfD7qoD8CgHUkNUhASpJdRnBqiR0c6JFqn8HZqtIBpdE7O91OEiGCToM7W5
WHCpQfiZMxRUh50mYZ7Lxe9co711tatZ+C/zwqgtNWzoBBsnoysKbWnSS6m9IYNL
yXtyNJTAhmwX83ZCzSDB/WRXk1YEyoZy591KW0aKB4hQvP1dcdZ861IEb8p96Xdd
VKyOLkN8CjVG8JTu0YdLAvKrqPFvUPi36f/FvHuZx95Z4qDei8Lvk8RJZkU/sJkZ
HHJo/IDS6flRhbGPCQvnw30G4e9N8heyKMtirBCFOu3HrvSD4CRdUsCsBzI30eeD
6GRFzRr2Es9K4HjvweNAlzhtw8tcWaabG+dIqtThRvDzQ0OvaPXn9SAYSeuv69Y7
+UINFbaPZko/cQ4109/iniL1zNIslINnUnhm3OmAmwIN0pVKZe9vV8sC7IheGtA2
OJlh65c+HkeYQkNe+SQT6vXVoDslwBM7cRSQIq4v1OF9Qgtn4oMaLFRDaWH/UIlB
5HXsTs9lrzMVXnKBEpXZ8N81MoKu1HmfFgopdojMZKzX+NTio0uES11ZXq9WTRlg
IEEN3jvr/W2XmXjApsvYfx+2z7++KF67D8AKTZn1KqjA+o3f7HVBbCPI1HXjygF7
zQvndQlj7M2TjnMP880uXuhlHsn3qPBbL9dZT5QpfiwSU0/nRGx8FOmHfWtmHbKV
YjhQs9gTv525pk36YpK962s6nJfW2eth/7N4qyW2lvvq/ZILfLxTlbl9+/L7cKjG
khkl6hmVMYf/vlnu+Tk+Rj5BT5gs0vv73P0N98TX9mQZEElXqeuOM1jz6E/l3+Sj
q0n7moI7lGiy1XLrh1SZqH4dEHqFOGgFnzH6IyggnNylPdJlr9miygX1RUjg9Ltm
MMGxwnNSpxgnGv652kNjCmpsKwWsY4M1q7Q8hCzAYiA3yqRVniyt8BInth52gUNT
6qgtQMEPnpnoQnor1Ku64XJ+wG4pJJ4vY44fyFLdLHbYLwQpZUXYMwBxMy8eLEgk
oUgO0gcr1y9rObF2M23eMr9KacRlFEIW28EZJ/MzEglri3KSG3LoFhkF0rlE5fl2
OPOacas2dc0dDhhvpH2MapIM8vzofkUbvxb4K+rkBoNTIAshVmpSip87c13ZSwAW
IcjwHpJDQQSXxLVfFEXHENFPnenu/DAQMKvdtfdjZmZJHP1LnYB8P38kYLYtm+Lk
ZuwKPmMJ0no2gkRwWnC7nHFbk78yW4RuIVLLX9KQMSVKSHaxOsPK4DXbQXLmcxnG
MRhjWiFJ2edAi2zQIVZAiJyFdbAG8Lq3GNTy6apxjE/1GmhWfvKeZIE+fnpTvbbV
tC2J/ls5zMUL4Tol65HP+xxRuH6p7gFtnFBcr9S+07A4owY6jK9v1DLfY1nmvMWb
VZdmLFO2uYj7IAJymPD6JHgzkNUQNcr2ckIo0gdSZyEbVEIima9NQSduukxeVQg5
zwANbAGhXoU0i+6NCYKBIFiGWvWHOubRxhJQmcM63TT30ATD90UqAZ59wOD47yxB
goB2/bBkggVfVhFMHr07Hksxt1+0aD3i3mfq8XHGlsJovcQmUaIdyply/D/VfPut
crvPqRdgHxCyfrn4jbTi33vXI7F7hoqPuY0P9/zVW02dB3z6a4R2qEy4fJmXrVcy
ZHu2Fk/xUelbZR+hASwTXoNvcxx6/BWUsZzHH/cmFtAqnXH79wVHn2Wkx/2eYde9
`protect END_PROTECTED
