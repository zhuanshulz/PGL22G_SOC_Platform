`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
le/lo8xkc4QrX8D1XboPbi3fNQ7G5COfE37WAE84YHnapXnr5TRiLE9EdoMIsNub
EMX9wUcR/S4xAmNKWWtE1U6RtI22ouneN1FCoYqJOd+gp94e1fyzXy05kgWvNxsB
s6KLbQjUmL5jFtfyBfQkfxnXjR4vhLrlVN68mll4qCuLNjYF3C4wSXEbfIw8YIIn
T34Y2tyGh6Y7mLX2Ln8kDhVoHPiHcJTzNWQffRevCe5ra3uJt9VfMxSwCR3TKcY3
1T0thV9BGrWItrXuoEoNJ0vslmV5VBSJ74AxaIbR+K7yUBisz3x/KQ4cX2E3F8r0
A4IkzkU1TOcYybg5cSn5myxU8596rcvv8fOFGEueS8y0lRC/+mIftrnlLADN9/7C
hStDtUqt03hU6LuYqr4fKn/tOAmQpbXg724YJ/NdFfs3OWahTp5L/KPsG0b9f5MH
hFkfK1Th5Irgqg5Cqq07d7L4mGtRaiJYEqbnA7oX6wXnWCLULOhbXUaE3x3qRKJj
u7SdBrJwMBX4tjmrPvBNQ/rG73k8n/WstF3TNELifbna9YP06C8za5ORscN2BQ05
JB+RJCDs6aFQIoUhcIoJKjCl6fdD0DS6wrk1x3mireaVfRZ2VGIFausIGNZV9Acn
VPa/KgNhxFkSxusNLTtXXDGHvON3u4S1Wcpy7XXlxQIzRy8TG18lfBVNahpa3vQp
ZkrUDBkPj3EioS9ItW2S0sHD/MEwikwabxs8qKFMmP8RW1+EE+BhvRTDTamyqXQb
PgV0gCSz5r4L1yDlK8y2ZvVVnBKU8cvx4tO5i4CXiBUmkbfuIENNhWvCcwz6Z46M
NV+15iCoyJ+2x1pmM2exWnM9MmWPs07AwMqll3fZuIbSepbpJtIelR7dexs5ddBs
uLe3kn93XoZ/JpCj90kGjCpP0UgUjh9q4VwUa1XXVTGDSgyFBAROT/abmwyc0IJf
tPoya+Xv4+cyAB/TjbgdcrBKhUcwPmwj7krqCCYjGuQX7KLpWaoH0Tqty4MWr0CH
/BTEYjCtafHpvX9Hr9WPAp3DWXDjUfxPw80jcXxEg5L/qwWA3RNJgZ6NRl3WRJ52
mVEfe270ZrasmhCqeFlSyw/tqEWY/nvAakpsz61TdZhsRAZDT8QK6p14etcZKtuw
FBSk8db2BOKAEftKorH7Sc3i80Ciex0vm8wfkdEZfFrKo+YjP3kLOTimNamacMMb
YoiFEZ2y+M79ZOoCK+LP5X9myfHmCBE1I2JI4mx83qpwzoZk/PYs7o16H07C9bNy
Rp15jla3Ei4iWDU2bzouY46MuI0olh1DuT/8AHgLJvRyeS58Wc8WDYLi8SLwYv2z
wgptHV1Dav5p+Z9A8iP4gfuswHvYOnbLj2ZD9nmzxCLCthqWrBff0iRx8SNhoDNo
86ZYFhVpqnS0cJbc3PAnO99UZSaO0oK4aFBS20u69K4tnaATrMZQLwSF+xKvpk35
PgQ/S7mMclFWc7XMe3M03FbZWuV5CphOXi4tVfSZICcQQ/vr7Nhr8Qgjl/lE8zur
jcLxGpbb7h8J8S0TyQCYmuCczLbLZuYxzeeHXV+kIkRtWbs6tfzTkNcwRnggoy/Z
XBU8E1LrgJt6mpforV3EzUAipgz4pdaQZvWlSq0HfSWDMiUNwmvB82MBsQwM3J4j
IQ1zOOzgvTJTsPBNrf+VvJV6uEbsOr748EIb44QLjmLiFGozf2aYb9N2EyKr9Aa7
JL7N7UmUmGFmYG4ewgZbuSxIkUHuo19wwh6m0f2wPrVDS0p3eD2cMCU2Ws4Qk/LP
DPYQQ7Mmq+NI2NVkhHkCnbONWEh7M/WdeZOWxB8F5MMLycFOe30zxhXpL9hmFRNh
fjpYxoRIZEjRnid9vkwqDDR8LAvsVMibsVzEHD9tL9L7WiJEbOejfuiPo3+nTHAX
pEHjWP9p+PZcafbrwWxKBf99d73FygmSXb81bDNdvYr6dolAKGtfDnvkjBPD00EM
XspRzpQSi7hgd3uSraAHkpUg7LLDFkNDazGTQntcOVUzkRyh6Jf5DOcIR+wa0uV0
Jg3J0SfJ6NuNMJEeb+T33eOK3D2iwSwMlS1Gx77w0oDD6KI61LY5twrGrCpgDQtd
eqZ4rHj8IYbcu5v8hO6WeECuTdaF+fduZBOoabKmhRhw2w2OMWaWF9VbXvwR6xWF
e56axpDGm97vVtY4kcCq3egVQDMR5TaMxUm/j3UEwPw436vzpQYyOXbMUrpQJJha
/HBV4z3xXQbiYGAzbIuLkxEVLjWxWCg6ea1p0AQNHWdHZUSVl8nGw9Gfa+zB0l1D
GLiOZL7wg616b/ZeoUQ8NEKfFEMrIDbSNXA/J3rvVKYJ3OLBihG7RSRCjbvQU+2l
8lFCS909WGWl0SdZZ/kKipnxnDsvncgOGSE7OJdMQPeev4xBpUr91ceKVhCb5yFO
cV/1UZ87f5p0veUtRExfYEL+noRCQ5qdoV777YT42QLkljAbPlp7WLf6ZO+tQoew
ev8wjJF/MEwOQXlq8nqigNMLNShh/UdpZxhkgaKjT86l+VaLaHVS/pp0CvEq5QTx
0wSmxEQncV4MLgJCSTyGE/JAsuNL2FUmYu4d/SoDfL3Ec4crzRhXNZx2Jkzn1Ts+
b+M/Lm5rrAZAlIEq20U88q3Hdttu9SZ3uZ7J5y/PJ1DeR6mSeB4UdXMwcrF0oWCv
UQtH6wv0/FFwYOwH4pvR7bW4f9YnjBh4GWqOb6aTuOG8w6ZOl3tLwXPB9bGA3tKi
nh0z/JTyJO/aKqx08qiReTAHLONIFCbOCSLB7imxU9GEUJcnv0D0Fknd6Y30d8nZ
s6NuktdVa7R7exoOsUFeaiTO1S6fAnYgW8MX/I4y7yqByMMuiKp0HGtc0dW0Q3EA
in983VPXECKZW4ufQNeG8kkfGNjqqY4GRmXwtCZhz2pOkON7127BzJhwTn1mAnov
0Xn49tamFDvPCzN583TeaIuVmzmZxLi+OJ6845cyOkhYzNbYDRyPJD6rrEDmne1l
oOOgqr7r0ZL2vMZuD4NceVI32FZnaOx9yn3xoEsF9nTGnNm+hnel5Y080t10cn1H
joCGcCB5LnAs5v8ACbsrT71z8NSLvM521xjUFIe/Vaom3zwn7SoZk6x3SlVc0w4g
fw1aOlnFQNfOdcN1/ag9dOMT3UfRsM8vD6h5nTQljqVg911FE5qyuDfTEqRz6MA+
TslXfm/B1CpnqEqJQAzLCa5mwEwyl2TSDOPQgWYPfltsPWmQEFohui/kVxq41Y2V
JoaVA5MqsxcFT2WlSKGu7zfEyqhnlCgk077dC7stZLklRsrGs6VWnbttyqFgK3uc
3AbGX2mzsj2yYmsVK4ZAoPI41Oxgg8smJhUlpBmbD+MhUPjO8wbWfpq4VPDT85sG
W8sr3RarpvhFogWVTDlnbBpno5LFzXGbWeqDzfzH4tVLWnIelDKQ8clmTp+s1Meg
TcMnEE5DUSJ0XYXUIQoGsMHzHdxkhe1KmyMyzDxJGEp4oTl3k6Rplarg0JNv5EiO
awkBctxfo5V6JIric0txjWIFvPEv+zDZwr4y9Az4FWJaMummXPIGKO2SL4XHUWfW
BRdBZwC0DsPV6EPTSuAc+ZG/L76nk0CjkShmdaE18WbklgAA3X74fRjZH9eUPSBi
J0GKfIJeJa5n8P0vUtym7DO5C3ZE2eTkBMLdJpfghmRy9zrlG3qrOy7Gbzv1oRoR
ENdRFkTk926ZzVC1E2ZXorNZOsA9dzESdYJaVmOBL/hnEnVUY2Ycy8FM1tftSte7
PZBqncqClZxcZQprPDuS4cpgjTQ5kuU0Md3lkUydbyThC8HO32/6ssp+gk4KFcLR
yJlNM78bn5hbmy7F824SfVLMyk+5WjP8SE1I88JjwlTmAzDEQlni59zGviLeZ5nf
uQly9oVwhV7W1ayDzXqqGSsf11owP3gxOKGNZv0NqlMv2E2E5bP1u+/TF8t6WH+3
AzN2EhNbm/OqUcEjZ9qwkpi0Kl1wHCyhjbJCYD8dZuaBmbgWGMtywHSL774WCgFm
cu7ni440FKq913iLw8O0NqHulYPPHxUdKaP1a2HdLWgUeU9s7N4NCMnkamPL1Arc
QNXcHHCWaefN1tdK0nU2xo+g7+oE4Dz5xA9C30sB1362sai7/mFvTEkupC3H04SL
PyYmo58k99qSE/cBRDvH0U9ObdnLtPb+SW5eeJ9P8SgeeKfPfdJPh7DnqYIQIgmb
UkYPzpdCvXDZb2/6jAkZ4yOyIHHyORLo8YCiF540TLRoo1BF//uSsd0hyj4EL87z
2jnEuvgvIeHsPD5P64/cjtzYY2HCw0byYyw7U8bT5g9nFpCN63kr8zWJaxK9eJeP
toIo27nl1iW7bRMC2yLciUPA4WKpofz4ZEh46z9TP56MKRUMSxlqrkrMjgihX5WU
qIKvovQ1chxHqPYaGVRytlVi8xA6K6osm5DCTLVMEyRUkiqE27X+wh5fW3hAzoxo
Mr+J4RkYEsGNYkTuAZnMdJFz/JCrHCLpG9OG5d1dvjqMUxIGLNCYqECufcQFgEHe
nHzSwFcM/k8FXxfCkwUed++wY/4V4oHKM1v6naq3Kwy9YWMlU2alEGtGU88/bHlo
yCFgJ39jofKNyZfBTslxIf3yJt/0QsblPD/4w/Q0aN4UnWSxp8SewF3az71LuZ7S
d3iZIjufjyUkzYcVdn2x2hflu3w8DV5SaQQ4Z0RPugmW1eAV/v3xvwGUqp9omhAz
Jghrj14zVULqkRrbmgi491oT+RMjJL5udFflzEnuNCw=
`protect END_PROTECTED
