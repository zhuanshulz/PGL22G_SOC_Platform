`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qrqp0d7Vn3d1VNQBOrTk7CdGcusO2Z5/3FuDt4YQeh5o46Yr4EKwjtGj/eDk5PrB
WyHb3eTzl9RIbC/Se2n6n8ToNVu4BIDtgGKaOs6L1VEsE5h67VJiyYFjgXHLvtBd
PJWTF3J5/kgWhrh1F36PXSiWpjfTfWbiX9vF8Mv35D+dyGX7dRLGh3aIJvqEtd+e
L/CQLRtcDiu4vIevVsjUgDEg3qwRo1OFnRopB57ooPiE54ZPERWsXT7bdmrKuwew
D9IgbrnnsoDq3sGHdvn6aFtH4kIlb60XSSNcBeOMTbfaHk352m9WL5qTFYOelqP3
QsrHChizvsUHHoxipg+vyUG8BmJNA+JyiQxVe/JVSqkRqulRJ6l0tte1c5CyKe1B
uG6lLVglR2x79DRZo+YSkiDNxcS0k5pbUUSyCKwDYRyaod6cJV1jOUMBotcc+dFc
k4ffekLyjnphWVsY7dgknmuercMciTObgdMXx8QBdc1BeKHT+LnosFDKKop3i3Wp
6jpj9nLYkmpAAgDne5EBquzXbnX8ZtPGD/s4J5LMDqit0B/AmWAunM2V3LE8nVWi
gBqV3B/5YduwutI3rJ4IrNo2QE3hg1NUvPTpgAzv/teB5jTKNEvkEEocT5nouOWV
ci8uMdcMkxLE03cJMbIKcPa+XARI8I/3L0a2FzyZGrHdiU8tX0VTTYXCYWmSP0QH
mbztXoipB4LS8QhQD64lih/FXUDeUxetIMdR6S2stnuxSUAh/SNmW2EmdNGz3D7Y
y8BLGCCsGcJa1lzXCVCbCRVfqum2hxY6gfJ4ZixBrcewlAzpSN9o0VKmPf5kc7A3
TlveehZT12laalC5cRqhTFtaJydhX6pzSkmqIBmN5o3ov/9NWIiiX4N9fWE3vBut
NrYL6nfXrk1KmnO3qw9FtsmsVAKpg4Df40awPHpTNbOLEyG3kINsSW2FiOr5AMpj
GTSkTOmCJ+UYSXBuoS0c7VQKV2SPlS8TkqdOX1YWqdKqW2JOih/sfXGq8USb0yh6
DYjCXfQTongxCv+IWJamteShO5fMka2GFEvP+6naLmcpW6Nrr5RXLBSS4WsHGkzn
htMpDM1YflcNhzKETtDNtuCGXGcsmsHKXvuuIWbwcc4/qrPqr9Rxl/VRQKRDSvct
zFHodDr5ccFhZT4u5iObYL62yHZJFhU54aWNab+/BQ2jWN5JSDep26Ukh7BrA2V0
wB5W3sUoBjG2hTzpffYm2O+sPf1xeIi2gAHptLU1U2+26CS3rCGc9mkTkP7w6bII
fQ+i0hvaGZaLNOIpqFSZU0ju1cAPes7cCfH0ECY9YOm4/W3b5AO5iU6IWDpBOiKS
g2DCjwWLvU7l67phREvY96QQwFPODTCSJR3cQqNBVKvKT+ojgKVDIt0q2Orzlqbu
L/bov6xy1uPjepz25Nl3RA6NSEVecmIpXNfVE5L0ohWHHQIkleSP2CgCqqs9BT81
ykG1YbKNmyRq0K1WPsZAycvaVDWxCULeC8FxUpfyljEtVZunCOV/Qvodyb+k1gth
WqTJeiKwAn7jGaGkHYeoUXZcb/LKL1xw1fFAnN+C+wmz0YxfpKrrXiSjndvSpuzW
482geuMB381xTjMOYqr67oSeKPq+pbOaHFpnScXYj4/ECDoDsJxk4I8NPpc95zUR
HLOnkVnytFhlVRxnoyeQEqh3N2LndY8fnTpq/GyPWpnEBRjbe75jKa3nMDVyXojD
tSRlzyeRNOUF/ZjmgDBMr+mG5gGXfwbpIdOzBnnRyKBe13XuKgxx4JbkM2vcCrSv
1Rj5xXA/mEwvvNIAAr+7BySgfkFJxPz+wxR73SOfGvmjKSDbjkQ6hbjLudBdyLL1
CysTAjQlw+iN5PpamqDWxIg+qyoNaIeOzSdkCWLWoZuwCjc10fAP0eJtyGWLmBLL
/NW+P+nBhSQ7TJSzQFfm284lASU9wyN4vjkgjT+tPFwAtL6CSbUZcndo3uJBvDHC
aFUlg5xd5sMBATl5CdPwmAbcOnPCwXTQL0jl+670U2xouSVQakZzLlqWBCZf6EUg
ASmqcvmZabag7VDcdS7B1raGOEwyKKRx8IuTQza6Nl29MU9XxJae7AjoON24CAiG
aqNBbcItIeID3CiQE3tIZxDdx6lHKjnRPXYHVDygR5RpUyDHz6QHpWdgPMt5wbty
+YjFP+/nbwpW96MoAqJOd0JFOhS7Ay6nDTiJ2+KDaymHLG8PFxrnZLSbNqKSGD8Z
cr0vNbtJ/ee4YWnJekhQ9bn/fh1VfldQ3faxFMZfmS0Mh5p8+RuWgRlptb0vlPCK
u0ZpvQEq4DSSqDXGZGwXgBRqp9L/EzF1g5WC4N4JLL713cnK9JfA4HBK7VpoVYkK
vZh/DfkO256khkfvJ8/FHsG37ezeN+mwXaYIQloJhClVBqbtZVBz7o/38qkDqtir
31kxpB93GI8i/c0kuG8I+mJgOpXlhw2GKKMO5PzLQa5uAwvcJJnJvtA/Dw7esaoN
HiU1kr07SqLLLPTu4i1+acWvF9q5NBWDE9LYdTK2qDh9rnMsIU5BK9T0Fsgmrq50
Oa4ibeVP9kev1AWYnh7A9M9hG04GUr5mJYLJT5AWgG/2Jt2O/i0ASq9TB2+uYcN/
4gjVxMAybNSyfyq0Qtk4HcDJfRqRRVYmwg833BHVeQMnVeZ08Hf72svpM0eLHSjF
C83G95VqIODenBALWlx3E/TvdKc+dhWUdCS/xUBtjG8RBVE/6aqMqSgwQFrbNZ30
NzdHwdnbFfbGqQ+iZ3QCzAddEGbIMGesu6dSZgpO0pqdH/n1Pv1M6jWyznC0aj+2
iVNP/kvgZiUiizSQYJptry2M+XNJjPqOLIEpHnzylsIDaBcq/cWBjXhn2hxsbHnr
MOAVp7LYeVENSkvh4RRgLJL318x2ZHfq0SwQzJB5OzVnktQaG7kf5Bf0aK65zNgb
88QOBQqPIc4PXawDFLsw4ue0dvdwKmaGjGDbxsQ55w2XF3FZUxfNfd4jU5YcFksC
zCRpcmd0AxWqVE7U2It+t78YHoUZ67BsclsOfOZ5hrXgQDVjE626u3QUPDwiwiA2
xEGznZSZQBOCFmCzG12TduEu/VyqS3oL9raqvi6AUH3h0XLT0SkU3RaStqwciS9b
A9klA1+IBvs/m4gaF9rDtt49s5RM0MOpo5ZocYdQGtlcnILxI/iUwNIUEjeCfgQz
KIjmAbRKKsBUhoLVeTnNoBi1ojkj2llhZ65EdKdt+EGA10DITmRiK3JnNxrY/Vh3
gQpnB9Q4JWHHnThnb303HQ7oynjkG94uW0RkJFBTpRNxcDxEUaavV4NnlLMWhKTP
wXtQc3P2c3A75gdC1mxy/xe2VCBLpbGuaw8bmOiAcReDSQiFW7GVaAyX6mn9vzQr
l9519B4FBh7E7A+Zl4qXFjdiMYGnUdl/ksGdm8oh1AtQH42mD2kgTLjkAa/YjqiK
ufKz5yWxYplBOngjaVXUPwfTn4M3kjweDYdbNQtDFZVeA2MqwzHjU5Lc7borpwv0
93oz6jxcaImART1q2pM1tpO//O3jmsIOk3jFlrjw+GKNef1QbXvK3KJj+MWtsu1g
mFsUwtKTv4npan+etGiXax+JIkJgvUwLgau8R1fKBsVyaEmMUP3WbO7qMxrb8e9v
WSESA/Y0tQUVjBX5ZhH2XinhIQIQPTAitReOjrLjfyOHnxRX803IlmxHWjJsaD2K
dMBCaoFvw/KzPjDshV32im09ilo4Bfbm5kJ5CeBzYtn+r0oiPaJuA3Bpwp0LtuTX
76UtsigmTCsD1VJpvZoAwgTdO9GC9PSIjn8e9VyPhkedBm6b3Ia1ShQ477ysmL1L
joJ3/dSP+Gd7+F1ktfxIFZFQCWcWb96srEwoU39IS1ioJKkS3orbEO5LQoX+Z3Df
8vGJbNUGCKWDWItG/enjQMmZM+dEhgnhfp/sX6cGwRhK4XJlgMQDL6LkzWgQ6ldM
LelRU1I/vIl4PGkUvK9RCTVZkZZcFxec9FJ3gFKz2VTFtjMc62Orm8XZs08qyqwn
Odc4bY/Kt5joFzbGGrptvK41jB1Hmmt/O/Nt4FIkOHL9CxHotJzQSb+hOEzQcUna
hvXymNBOuLtJjVipq8FoBkKVQwViXn7RK0zD0FhQ9n9CcxLJvmGV8o2lLNEhYfRs
B4sRP2R2PxoSA8KvOdnExBVZAjXPqKVbWbp5LZSHh4OsVRGTf0ZN/VSgGf333vfq
fdearljT7iKqQ4ekZEYL6HcGMjnNs1thBzPgaaH7wsyeim0Xj3zWxDNl6cFbibGm
IzU/PmP16dIRprfGKwzNVLL9RXOLZHjVJ4ZYfgDHzeKPqPlpbGOOzTGOzDpTeZLT
qdACH/WLRLr3OekK35ewwhp7XGjiEGw5JNWaNoOFlgo0By1ZhKcc7R/affU2gZTy
pNosHMof882uPN/RaFIxMfpGuT1bT3QpouJeeHdrHWQcxb1CQrtWgOY9X0k321/V
xJIMxl0xm9jpFeDjtnp3ZEu1kqTdKaiZMQVA5BZ1dhYlVG9bja8zkuU/LvJugtl9
eu5jhBaz/0WrGTSvXju95q/HPobPFT3Iy3z2l3L/svQXB7b8uoX6AIFtd7JhUO9/
0tC4bgVDkunu0yzNRRjI4CQq2Xz6ecVB56PqbUgiw7b1ycJ6oQgp6jfFUougX/dl
qoIDIT5hxxHDRTjDx7G7Rn1NaHjQr+z7+AeNYGLb2OWg6BGLF+cNkbCO4WTTQGBH
FEPaFLKj17r4Dk6drqee5i1kw6JC0GFix2Z02Qko11YWpFOjOl1QLTfad7mJMB4T
U03x7IjKR3F1OP+46nupqsQwUQk5/EEyRcr9PuZfMbjwF7KLVKvZhnAXsmLvC9xZ
ISYoKnKexHMMPBC/W8AeJtLUr+bi/qqG8NNJx48QSJ2m1uEI95G011x1gUXxe9Kd
n6cJGWJCR7LM0q3gqTvMd8TBqZjiNkOxg43SJey3/c2qvQ66NPLWqtfBCzZjFbF0
95oZIKlVdt2rr8E7/v0Roe9uRAG/CqeZgLDtEJntQEgy/5lvXIu3uwvg6IDZne2/
4vSjjYyzLtXrh+V8I6M2j8CU9tx9wMBMVU5u8jCWqNXtJRzcbGvzwUytEe2aomEW
n35mpZbJUXLDU5EzJe3zAVquvKARUXZvf7v0HKdFxMqYPChlwctwk7hvGB2QYVLD
ZRMpcEA8MEvTdPleOMRxtqdQxL+Yd+vmredXNz9vq4/8B4yRun7xi2SF0M+AFKUZ
c7QPMG9JWW/s9zld0hA3fxapwoDvTC8tawH6xE+KWHIr3TCclZzlRP5/mbIO6eme
ppXoBpfB+nT90kOyIBegZu1hrwB4LOnL8cfg4Uo9+/ku6UPMio98G3Fv0BjIj9rX
Mqmbr1BdSHCIViLivXlcqA98/KS8mP7gbapo41ItUthDGnrZkEP+HQ3KlfdZu7FE
OkrA6ds+485bT5waVt+s8daJcykXC1LhYnQ6dPeiPoAXsVaaGh32dauX2Q3vivD0
LlvzKhhfnkqhPCArCaOCVdrlfrY/C4qF7BSty3HY06fLko+KMWCU02nB7osjWpcZ
xDeQKliZeM2uf/8b6BhhERTuIVqvoS03yx3PXXjV78kxA1ztt+smW/p1C/ZNG3l3
xUzOe5BVWfL+Eo0Dqh3wiHZ2SJNRxNjv3RuTG2iv26BNSKz8cdHz4x/jkOQYQF1W
I7/4iWRcYxqvX0EV9/5dJ5mDtZOUuIPHWvzK+21axtvnvpRBYNhAdMFMcnbRmoen
P4Rws8fen0FVyZIp5hRE0KMfywXupMAPEM/4v3vUtgMmvpTwpR5rxImJfU4txp9i
saMLyJEEcCoXkNv4Bum9MxGFlUOYRJURp0L03MRuKEs3YSxdr6aAct+DXI8T4xYk
DZZLKhq/m7m+f3hDD6MO5e3l7rie7ONu+Dl2WDCAt6wUaW/nqxRwwXV1JvhJHwFS
BjJZErdy2NNSHiPQbDeXqeeZAOG4zqwokcyjDN56OYCYT8a0JHTJ/50stVh0U9I2
PVtwKOnszXS0J6n2Iqz0HniV93c3UmLtGpQuoBg4zejROOFySYA5OIjbkUA2t8Rd
FoMt8KxCKKOGxQi52CHP4d4xjgLpsPIOdLp/r8emCVGd4vXVVZVfOBpy7aHhrEZa
C/oYjuQKPm8Sbm67R8jlFsEXc+tZGL8NdeE74xoSL50VeThn+/n5ElA1bA86hvdp
P02hjsSkJtusFgDcbUfDDV/y0nvn8dAmIHMKqcQMTn1ku4qbSEyudscKMvqbDK8v
+gICPMwiMToAtY9zEq8Kl4u3W4ScnY3HY5BtPWRECUOD42dISRuhkose7wRul/Vc
oH8N51uZ3PPjEaASnxzHlMaA8KgyWNUyNY/D8etSyKmWWjF8653C56c0Ag4JX9ek
0nqP4JL7DaapPu1yt2T1E7q0FY8oOuhrFux9Bc2Co8MmImIpU/8+HtltGjTeDfjY
bir6qkjMLxaTLH6/o95nGsX4CDLk6DaJwWaOWMhgy+xY3CO+UeGl66aX/rcuBaBz
EneyodUPL0cyi+Rp51PWPccrWNR/2EI1TvL/onlBEjo0y7ksFd5bEt1+wl63whtV
PQpl03uoW6ROYaLo8D3zlvcrN4jB9pbggKGg2GZ12LslWlKcrU3Osmwcbf2TFtoX
UhrCegvY044gm3tI1LcdMGLubbNb0NPL97M4O+KuaeQvNzPT0m8zBWzQCGzF4V9r
y6hTVKAJnQmCggxlAVa1nid5S4fW4GGwc/HTJtmE132yvvQhuiB7hi23ajzSKx49
uF3xNQFkCAYkAXzahsuN0pQOjCqt9zY99G1x7YuzL1Igzc0wIBtAsh9yZ63jNnuH
9nygMOIMNAK9KGlC0WKYquUbXRwDUruXkt5r1W0374qNVWFzsggmAsFgtfJStFQ1
cXVipFnQXPaMZGWNRE5QyGr+b3f/y7i7M1BINVADvvvGyJ8CeVaF15ukSqfBHmb7
zoU79UFQE9bFyZPnojBWPAh6nCqMKF5ZlH4Qu+zQOvVc4g2kxN2nkLvqZS45IjIh
CMi1IkjrVfDfEA6rFGgdbvwlPrhXhEzdX1jTT8+dWjC72IwR1pzunWzfdqdcFJct
QYiKUCgTzguZk5sgt1jgu9LmLXZz8J1mdL7lmLf8E1FYf4pyJUhaIw05f7yD/afS
6kJZtjj8aG35fTaqmuzkSZajk7HepOsprJrM6YUqSEIuNx11Qh9JS4zVVWQUErLY
L6MLp+GiRHkslu+/dkUTJ4Z3KNHDqSF+InfrAXT888PN8meKmi/++XW2fnyM9hX5
jkcsfYcSVjdguNieeecNqqZJKyITR/0jxFiZEA6S72KJW7U3a5OKMSn+Ac9uSOxX
+3U0mKsBY2+pIZlxcfNPAO5W6lJZThSQX3NiXb2m7gRUcP5LBkdAZaKpybYP6Xcq
TdoRaL/AtsxSCPNWjMZWJ8mDYB354l/+yA4n24+zdHnnxZSus+CGXlWXyXdisNMd
yVZ1veG5OcbN66No9fZWKVWZSiAHKVX6ukVQD2ND3dC9H9OAqwwyhzb2zdvli/UK
c4BiLOqwQubI+P7d6j58xdCZSXUlLUhswDa9Bm6Np0JVrfsiokSP2vGSPvcbgkBC
WBce/Wz0oD6gnF31Nqg93C1/nU62Ru9XoU2IC42Nq0bYS/clWO5gtYPRtketwP3D
+9tgzUpVd4D10ZGOTi1ps9qpujMpx6+fLVxwJHGFwAwu6UC7t9aKBYriqYuuX/i8
GB8667VztjWjgKnuOI6tT/SKwbP/TD3fbWrtVeLHkek2ZlxvdfkaKj2cH+2taKZe
/enIWZTAsKcwTQZ0VIAHz/0MQNg7FLtj/DhYfeRzzvPk8Kfy9p7nOAAGbkPkRN0L
FJqlX1mBICeOi2KCTs+ub20lqHUBihNF3kYqvEnxNu++hQG7JRAW+jIJ8it1UAmw
HvIffcRZJS3yBUDRD2kqdJTfpAy6B5iqBZr7mesW7/yCLJ9IFMdcZFnEP2zZm7FV
1sB9fOSLI1BcnBj3Wg9AK28KaAM7Zgw0uxQ6W+k/T+dVVzLhw8pDZRBMEMVq5q9p
jC4lBh7rCjHxi+zYv15aaS72RUa8OVfJNdfYEkAjyO6oqcpokZev5mh8XiF2EWxP
DBOg/FPKVXKvsVlsKTo1/+V9Keq5Vhi77u2SKzfu/dfiOdo+5qpUNjShraFI0JGW
RQNpNSNonsOqYdv/YLGBoR8AUeYkODszvu36ePddBnOzhoxMpM09KIGnk1OFWMsb
w5K/qYzIzjVDIcz5kgim/m9QzEyYqUkS1w56Ee+qIg02Mtib8vk36LqEajSptScX
dgtLOE7Hs+d6MVVCuCuCWbshlV5DivxmugcTa+Rvb0H4H3uZz2ex+gHiVGLHXLEx
eazOrPBXfCBuURJ/Xm1/Pw1/jbx2P45BNTRHv5deeYN+urn1XImf0ynfhCTKPR73
Na2dkGQ5ZN1e1OM/Td0Sv0DfeoDztneijEegOcS/dVJPo9zVHjzzuZWSc6ne8ijs
XSuhKQZdgo9KLCq64YAqrG0pZIzdwL1YO6Xki27nA1m9YNn6kBQDVGXp8SsnXRGp
mV1RJJBnVG0vSmp9d8YWk555zIr1tX/h/Fc27va1CsAXs29RTut+X6CJKPOJ9zzY
O+RoM9Xv/8EUm8NnH2bKncDHsixFtzlzThNMVaRw68FhhBEDNOL1kFajSpyi8Hq7
0ES1e3nOvFbDR3vfEXvUK2KZbiX5vX3IFD1RUI0CM5vAUgqVtOpUmsvT3wX9LI6j
1TIO4oJaBO+V/0CXSSk5PvKlsPzzCiQLlk7jDvlDTcXpcw+I/FbQMEIjMIuXDWXW
hTTxoRqbmX7q/XINolK4FR0lufocpglJsalw60Q9C8oTK/ysjnGaXV+yi5P++ocX
KJhiE40Qd24qWtflsLNbPFJi3jjlgRFY4J3VkJkOIPWeZE+LRzpv66azrQBmiyPg
r1j18CSVITqr2tsKNY8SccQglcuDqevhW5PslEew+oF1ZFT8esYtol/AScr6HCbi
qfEZ+BkBH5CZTburmROADdRjcPLhMRD2MlSUmboc6AU0fBCHPdVctW5gz/WG9TMs
5uvwxGd9/hjTgSwyubIEeSUbSb3SosJLaxu3XcAisz/5Ub0aU7f4CdeYEn46r3u2
88Q4uhpfGy9hx3RMAjPzTSs65shxgtHQoxloWHncUwU58s+Ehl15tUeFL82dADCh
SOAocu0xQokq/QB4rTNNRLCzAUfUUMa7M2qKRP7dI7pskuAxvGfK6il7eWQ1ZMB6
Y0LpGYnzYTeqTz3CARhgVaa1sdc4GvsQ0AMQ+fjcEwIfFP7k7QdxWi6wqbuBJhK2
rguEFjCOW/dTXLuVW5jtcPk3/yXNX0LkQx9ex49lc1bXl2WgvQ3qtUe2JKEvxMRq
+NSs4i0+kBeMykIAZk/lX5HUKl0EeEUphmQoZCRpNF/UyFgsPMe65ZKIfxljYb6s
RCbcAhk4sUznbrrSACAMdKbRkLMGmtqcI/rbrlsDYPQdzOuTHdk5jheHBI1tcpTg
Fx8BM3mOo6hZexE45j4c+mlQfcS6l3iQaPXaLjuqCUyKZElO/z/gcBURkjrT3/kq
xjXfDg/77wPPORwSPtJcGM89DM3XMx9SCk/YCi5t89qARKf/B4x2QNra2zxn6Jo1
/Sf1SMC0YsJcczNCg3iDG+5dAxtE9cU774LwmbfB4CAYGfWBXh5De5c7XppvG2Qy
/D5b7edVsPs3F4Rt9arhVLXO40YQ/Z4NTABIhQxLNDXOBj65IUgOLY9/uBTItvM0
/hO2rJlUE0TOL9CjNKURVxd8Fn226rGqW8bKVmaBOjze9SzDrr6SbYtaroRoI/Q6
EYO6zd2gp62PrI/GQnEIWl8ckkn285AfbW0OfJvJI2jo/4pmaLKATlT6kecsJ3fV
XZ/lrIjxnDH4QgBtwzkS1vYGRFh+TTeJlyk1E1rfZMZD5QdDxL1eHw9bgc6q1MAK
rCf1xNxp95VyybVSjq9SvZirmNyixYAAhGa8bgTzNo/qQY2Plq8Vg38Nx4Jq8Puo
R0EPus89qw4geuqvi3O2iHeDJ6RNH2g6M8fm9JmB/I5E40MM7H9ZXW2XimObjMFO
lCaulvPSpofswGIThsJX41bVMS64ZmrpjT3Csg/UPgRvCJ9czm8zOhCpj+NJ3dW1
luHUM5xWaY6DTfa8Ot8dj7b5oRomKCJEzBoIfkYgTBaaZuMDtQeCaUfcI46gQ4qg
3rq6zU0x4FTFR4ojmU2zQ2NBHweTI8iNCPiLSsAOzPSA5JbJR5OQ7edkr4Rza8RL
BLUnrdgIfzG79ELPqKLsFjJPKad+fUD7uWd6QpSd/plTLVlpTUxdtANt5vCM++jL
GkKbtu/vaAAJSTQCVRXhU1SRXFZh5yH4ipPBuFu9D0Mq/72DPmxDDkEgUKZBTrzW
6SIKoGcZDm5kC9V85+0Fe8/+ne7yz9adkLKWhss8uP7oDPRbusAn4ZbfU6cabriC
6yS8HGcwqfc2JUUnFhgKWTzJ1RdNALDcQMZaYrLH60d9J61/ENGE1CsDlup3RFhx
fotQ1FDxNFL+MhG0bfHHc0TSNXSgPN2R6qZERl+FZh6OLPhJvFCb9PoX27ENPzgU
E3HHoXiDY5FopAJ+okzuJFM9KjIQ/wDLVG1lokiemnDjAKEA8BNfbZQ7Bece1n3M
UADEUXoPNr/EGBWuChU1M7BijXxin/2sIHIsVBDY855hujSVvnP+4h+XFoSBwAnR
gkHETBwQ3K/bvNN37Ls4/9kNIZ+Aw9XMqwqyqAnx2wwgLYsPiqOpeNo2M2nkm2vI
eyRAqlzGHsKk/FSVTxQstIFDBjtz+HSu0T5eXJGATcYaTTzaeHNE5LX7WitoWXak
0a3rC3kae/xfTSqiriVeILlh6tOCf1+a/11K/ANBf/a3MH/ghF9H4IrMemxoUUmA
JKicIGARwqTrAlscNDydwtdVhtt64ck0dhMRzPHFqiz5aZFhPmxVGK9wBop5Zble
dbo9ndPgkEvXj6rMFfrOF8aMwbZZ3EizZ/F1u2dqS6+ZeSFJ96a+zC9UU14V70j4
JcMINutWuMXsk5hBaBIvN/nBLUGeAMcs9Qexv0BnXb7MGP7K2Z2Hl9c39fMIIONO
B+KFH2PNtODNAOjpAwCc+EpGmx1WW+whs93Spn5CBuxCrY7MqxDa92DtA+b5PHuD
1YxlMxBN8rIyhJ2kPsorm+W0qtw6oP88opI98hdNGeuZCP5fLK5O1jDdja5/0JDV
QSaJOq413t9/2rAHXJKnBBRqBNsN962/GMjYIQMm7MFOVaqLQ/IqqfRgsXKjCF53
nPySgCpr7tQCFm+4WEY7RLfn5QtbfzpkVGbiuDk7i2KZbQyzqa7mtMQa8rRRKpvk
/9Pp+X6L/wI2gGHT6qr/hd7U4yBzfkwieJTm/vhPEdu3t+MC84/MliQFkYeMuOJ+
dp9bawndepGadR+/7yPZTJ6FJMKYKSWYLTbK2MvO+sW2XQ7CE++TNP4OSkUdUYXo
4VsmalTmvvi0SadENIzf9Xa2rp3tH75aww9nrn86c3MDa/C1EcfhZ2/f3mQ5w5RM
f0vM+DmRoCw1PE6pBEp9iiUb66XacHb/ZNeVb8cR1eRM6HUQGk6aqONcLWpphiec
0YzO41ODyE5Rnraz1nzwPGYvifP8P72TLRFoMyZBvSWH+vgK3iySYaawPOz4A5ZK
qoHu7C77nRArFSa/OcNvEJ5tmyEUVUhGuzUq0ZDFlVxD9n5Oauuc9Z0EAzkDeRYU
swWiAtLYnIP943C2l8TA04YQ85PieLwKXL31d9XKgaFIltF1g8rZcJ1hOyr9NXFY
MNB6Z3Up4l3dLRMWwRvQohg8alqSRqRXJFBrrmnlqzU2SYWtQvzkGvyJ08DCRJ3A
L8hjQ/L3jTqFJPlxabz44F4Kis1sFI1P5qn2K+20hROCR1Ii43PP+l2Pfpu+IJsM
yTxebTbNEEZrzYBZHCIOZw0J1xmSCFDQODoqyLxiCkX1l9BRtgVzYCIoEuLmUrCY
5YKARcIoIY97GiUtc8LK69noA19fWyyi22Oic53KmT2nII6WMfx6PB3id4niE9vF
JHyWCXxyjdAak2FQCvclYvWUrsvw1o2AXsSsxvdw/gizYw2nP+SCXJLmVuGcwglH
7vReNxHFFSa5zNch7iJuO+AFX5CfQGE9jUnBGIEIu3n3RnFaVk9eCd/L1nq/KeHt
6n5r49dJSUnBjtOvapTX4jxfZwff3ayCXnMRMy4ccsElToCRDM0OmXyJNxueiQ4P
4ttSsZJaFkByX0ZkmVQVc7KYxCYYkPDEXmITG46pFn6epDHY045vkfD/N4YGNQzP
vOcloh5+nXk1+gj4ohMratpFNn6TAkElXWmU0BCXvRbChmNdvsx5EId0582NGtOI
Vrxzbi7muAoO7iS06QW3snHFHMDz8gIgpN6NnvkOCxT74xby3h/qPxbidY6jtzhj
yOcRBBqUWDQu6pQAeDMytnM+iXPbwDE1qNURPfUVbOZ8tiN9F59Phu6XmncyOlK8
TttG0ipyVGJ+BtsiPcyQ/r+nxJ6jQcKTKr/OAqNlJemFZC3q3JCQttV4tRWeDZWc
/xgtHQgLk8lRo6+64DAv+OEcTMjPEaU7bgjo73im43da76IqOnHAqpspRI5Yw0jI
j2OuzUkuXlWV8nxnatfzNo1u/0ZmF0Y3R5dO58wPwys+PUBW+TnlAbagqhILTjdp
uRMn4D4DjIBmZlaD5WZP6I1Uw6uJ1iyNhYPsFSFp75kaewWqTGUYRXBheW3hrk47
IxQYRjBd2530YqVbHoJPYdkMyfsupcbecGHGN7oWQTUI+eIvHc3/4mEDFP6Db6Ss
QiySw5ANV6kUHJ2tR8TOWTJKIbOr1Ln2dJZwPvlmZbBVaRxjdlwdow8CNZLQbGse
0/YOC+Vev12hl/0aOgWdjZDrPBn/VaERKZDvBDrMY49jsuqCLbJI/phGQTuWLu40
boAKAWC/fK3A0LoL+fa+H2huNpjtgc3B440IPL8ST3nFbJWGf2OmYLI2GHQKVpHg
g5rfWjUNatNrSDABx82HdHQd2ZtQMNYwH95UhyQkrsqYnDf7BIn8xbvxK8wBjZCP
zcr/YYvlQmxJGY720qyjjs2zkV8u0Zr5SiJ4FSGrCeW7p3o2anN1XRzubGebLb54
2/6Qp+u8tEqvihWuqrHo/kdtAXAL7F0+jwpjVj6Vi06pULcRb6Mj8waxbgAfEt6Q
V9fMgL/dAp/JfYL6S6baZMoLbhFqndg3IyCGRwrLYf0cXApkz/TLvYhFg5vkrJpJ
I2JcH7pFliN6Iaw/jHIT1idYSHKsrGX/84jFojnKCxVuBTprOQemcorllZLNiG7K
tlJbGnSYE/3OWf2CDuL5et2Nm4z8wW51XSntGiEX3L3uuexCAblW7cm+wCc8kNkq
Sz3LsAtBKvx9ZZRox348FOkiBChTSt0UD+igH79UszIL+BhzeVMksNUqQ43Tpzob
Iyt49N7pymnKuVEliqxwEf/w9i3NWnRykz+QPYUUZDof5lOLp0AkiAU0FohtebvY
7zv3LZ7KWkG1qUxzliAyV6P93CrRiMBneYhbiVgUc8eerhT2q9YnyaAchLM7R+5z
/zTywcKticYpKduKBP8670j4JyYKXbk3oxT2H1vwItDrBzyx+kOPLpzpYweyjFa1
FSWRQfcmSMzP0QwUMIcDkbEIXI6cAHSmm79Ghh8NmFHn8y0Rnlio4nxEyLx4WTBf
oImxAFkcuZhfnoV+UBnsInUUklQDh1m1ptFzfoQGeGPuGiBE3bS82T2wvAOoUnK+
SpKYkA+9OeBa+AyqHCorWJII4ztoe8ZKzqj5vxHsgpelmsOAxgOQlKpOdncWe3Bk
/3mpfoy9bgcd4HfPmT+857+TWPqWjv783CVsgh/WVgm/CnzEs8JCumqmV47lNxtI
Pn4iCiXdmfAMtdtrlMeqlpK3sz8Pm6cmV82Djg3WcjB1LKNh1KmvpZ8ZcVlhgdqh
qZbAzdymAYKMwoVoHz3nY/mvtFF86wkVapr5OTMlkE8fL1cnIDb81XixMBxGyF0e
YOl43G26iR/dvshfr2Khn4Ujo/3mEibeCfqf+MIrl/38r7yhZopPuyufqnFLSgOh
o9jBtuLNRbH8pCieQNYGgtCm/Tf6mfejsrF3ZYqk/ejk/McTi1TFfahJBmnLGwwQ
fP5K0N9URwuJKsJa7qYgcFadylLM51EUzT1X/xAax762Tg9Zg32+hhPeKQ8WWDfC
GY3o83BpLS1srZaz/UNklB8No4IETWJsxDyyWDYpTqZnjQODgCJZJ0zLP1GcIyuU
kDA9M2lHiflYKOsEf6XhI1j4dT6zJN0hyNgZr7KhRU1a8wJBtTQFl1HVz4sML4gR
NcKqwG2eSJc727aYxR5HYp3EMrT9my0RnhBDIPHrTjM+YueVses/ADMNeBW9Pl4B
w+UYB2K+HiWPRY+yylOoUgPV9E8kTSmr7krN5UrDAMfAGn0/DmhEh9hoM3DZkuOR
4yHHyLSCrApcdkDIpR6rfGmuCi55XmNFJ7obFRVjdtey97KOzPs2DTOyHa7UGMz4
W35dQYu/4U6u4T04m6Lf5/2q1o9d092P6bzsf0eoG1PyKVy34KHfA965KrgeIqB6
dzVQZwVYbyKNpuLEH7IS0gEUL6HnahPhCV58KRaUsa1Esn3umM18+ZVVPJkYT4v+
oyfF7HOyw0+bPjqZkriuWpH7q449imrwNptk7YPDStFbpDidZhOi/llJ3/7Qr9QK
ddqvNsz/49BNqBu0BqTqvpdF0dXyJQPRaBygOGLYlqbSt/Aw/k3gStEmoe+qOZ3W
t3y6LKzBO/r6OmHHXH4LZm8FVJkBuCiNXwN/Ut4IwQowGeUgn9GYDU+lEDHcB9v0
sggNwQ2fQsmhmIKIEBWfqynjhsriyOC+pCu9irGq6x7qcV2Ly3ibn4GEVpe6vdhJ
KRhZVZWHf3G/J+7gPRKPnmTG2FgmlAu58/Dzk6kVQAEiWLFiN2TF0aYAEmkXOxvg
DVUTEPPBCLZ7hvNjeTZ2UPGSx9lcf6m+fF0y4H07c/gFC/TxKZ71ZxCnyIcvAALX
ncqaoQTHw460nGJ085/O3EbIeZaLVsaA9TOksTiacBn1jJ74wx/SmFAvJpCDAb0B
1CsAJlmHCXAaStuNk00hivM7iPEikvOHX+kEO7A7RAXSybjP18L+c/+Dy+MXimpy
2aQkUOgQNHWHqtDt12f292m0X2DdaIRBTMbI9vMUNim3EYtsnIymjQhmvpzwSZby
R+b+i3qj9S5Ps2qefQJOEaeZ/an8JqzJeaohnXqAtp0YQyhndgR8LuqJ36Oexoji
o/SVTtivQTzFpUWcb4Ik8MyHQSVMjEZEqyBhUMQ4RCxVczvPuQWnsSz0u0Y73yFV
E+5pH6wp+cysap0saOi+89g/hp6OXJzQdFz6NNEtjnpCCORVybPsUaKQMccSIxCy
LFwY73PP6yZDUI8qrMW0VMMTTZ0xuSC79rkH0h4DJvaVFti7u18YZaBppkA4+G9V
P/NaJuT9P33o/5wjhYYgHDsdQUJUVAGWLHpDnu2qJguvzvpBN0xdgfIX2eVReS8r
JX9fW/mHZ/yxbkpo8rvOhI+mZTk3K5QSfz5n45qpfgv9xnkG7eeuzjlUzgu1DcJP
u/EfYiDdA1D2SYf2odw9hZ2HFWToSSAJTavDOIytx5Z1Z7yV8xE0nqv78y/94Sza
H/m8GddVerkwEB6zlYpdPxZQ6mvizGQIAV2OR80gM0rhUFsrOskp0sBABIj0DAnO
urOiH4uKxG65kEVQy23hoimQWYMufhPnDaLYNTIo3/tTXSpK+XCNz+UDc4aPcmwY
/FT+UYh1wKJ16+c0HK3yrnf+wC3DOtd2C7Ck2hViu0sjIWNxJsOaK20drQ+bQN/4
BPoMc+Zn2eisVVhJyxd+/f8JCwEkWIyC0qrOkSQsFcbF2nGkvv95WcYsLippvvmp
v11/TstP3pyaElnzhjeoU9NSzmTvxmc8L1+WCxGZHsYPoXb8jUjHlnfFm1rf+QWX
62KX3BDskOiJOTjmUatiF+8VXDGDTn3WUtXXUjzdTeLCsHA1HCYtECJDzxs606OZ
FgxhqlZkJbnAI7UWkFWBhh3GnzcUmC1LkeyD1DPqQYXl3zgcJeLKsQOM4dlL8J2/
3vrTolaM9liiU/SNSzfMv9s7H5VilwzV71E5eRy5wHr4k9yv3uTCpOCakqd23Etu
7WweCmqtVy5sjxreMqm2z4CuLJzxvc7upitK44fDw/99WXqThlgqGWZ0rGDZ5Axh
oSGf4kPfy6/LoSu06yCrGRMIcl4FsVdOXmP5pfcbXlghL7buL1EZdcL511XE5Imr
kioLlfbJB4wN8di3GY4cG+FidCmOO838nLu5LXFCGW0e35VCiHiSiLGlaMZ2ImDB
7uhE7+42ryEyZ0/KhXh04a2H+MxkXwDFqoFPJRjmlc3O8Qbo2Q+6+ztembkLhGSk
nI4lcANqUQjVMB6eML3oE+5HooFy9Oz5bamG6Y8EX7WcbTfKFuFk6Rb0IcryyUOQ
G1gZQqCCc3Pmx3IcC9UWGoo3I4rC+Cktq5LIy4M4TruZC6qbfjmy04r+KiXGa6RI
j8YCkSdyE82nnR6CblrVvQRkm4K9gvYKmfEXg1WDwBGEUZPUbw1YpYSuG1LN7g1l
XOpR3G1T0G6dHXFO+Kf1cUAkQdPpwtidcHQAN9bJeV8vvJ/qyei6QTHJkiu33P00
D8c5WZIorHJWpGBSy4Rg904FHO3ZSnsqyyjGpi9agjy1MrfBut1eASSynz7rFxgk
bcjsgouyqoj+CQNHDhIZtrIMBAW/JD44ign10vFUMYDJOEOaKQYgFOe57KdS+gyW
kYBr6jsupVGIAogI3mXa95SEhqbIeyycncvgfeIrcc1Kay5JsYGf19e5ODGIOvmy
h0b14U2PC0NOzpka8j0AFgX/12KLJPMBnGBO70CFZ7nqi9mcHBj5r74zVUD1/jnb
7QkO2SFraDMqGR1tbsa0v1Nv1c5dLf6HhTENmxLHBREUjY8ofT2S4yd8mw/pnZWQ
ZrLILxJ60QyH7LkKZfnjpoF/7Q2ZJteLQmn76cQgF9Ho/YKm231JmlDPKiJh4SfA
oRxQP4mKyL98kLTeRHNp9JWu3w1UaBYQhQbXLmUiFZIqthhxGTIBJY4xhvonltqL
cUHWlJYKb+2GOlO/VXqPoQeK2NJmT6Kjdni5oxc0pWpTuptXgI+CeVm5Is58AnA6
/SigRqODDB9IDoudVKuCUkzEFfvfi1VkYWVM23LGRPPJGZ6apVd7D/leLBZGgzdG
H2mIN5i0x/y4mKvSfKQZoCpa2LV6YU3USssLk9pz47FvLe59FlYmlejwP+TtbnsU
787TM0ABL7wB8tPro8MuG0WeM8BDkrnZhYszBzy4PgMzoUcrVFhtApQDROb9Ahor
khtkfUkXOSNSN3ZmOVRStC4LBCjvLIgDAjW7L8U6zboswHaC1vRDEsh4o/pYl8hM
/+KnlMk9Ampa7iWlOyETMKZNw4absPiWCLuRxqrrf+BwSKETFejHyv0JrPDiJ0JJ
SwCCcmSFWEhyRcRrRImAJEekEArp7GGvKsg+bzrgmc2eaccE5dXW+wwME1aDqR15
VhgebBcP1xJIOGCVvvh6xukyCfdLLgXG4oL/ayyaBsMonB6+vSEctxxkMnvI0IKK
voSfGPKwg17BoCApNsPdbSnxK7k6TpfYFbEyQuQgrwJA13uHiSlg5+60cxvm+86R
D0t2USXOD6Z9K4Ttos7F8ZpgtT0Mk0lsTyQ/eKE6r9HkVg3bzWi1l7Ccfp4gfFUf
x04ug59b0pUNWuy0ryfPcL5Qw+6IsnTzjN19wpflVyl4vFvXOSVZ5ot0LLGtlKMa
`protect END_PROTECTED
