`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vzV/xiHKBs4zsFX9+huhifv/yxj3CFGKwgQMtJAA/QeO9mmCYaHXjkqkx/dj1Cb5
MFCed7L5m//tuxf8RqBm+dyV3t6/ebHiHUeHmV1M8+xFR7VtOhEBlyN/hI4XRK7U
JJeMC6M6bCJACKhUe1MfHnPxggnLpm6vXy5uDrBpPJwJiD79NcGuUyvMcujnfjo5
tF2yq9lCJmW5yMM79H6q7hjrmxsSUfiR81pyykMIzyGClakP6UPKEaIVJbtL938Q
ldPvJHqelsHwrr/F0XZHyKOsLjJrfghGatD/LIzNt3CcWYTbBVpCxVH3cQ/Cji4L
zsgQ8ziVNler8Jo/JwrFC5v/F0sJtIi7OV7fQO5klG2nzY4f/ZHNkOHgzNBgyVM3
qFry0PFGTljRfVs5JtBpzGH318/YUQdgIUjccRqG163YhreZTZZMzsSpviSAth55
rKyzez9u0p7DQY7mLu/MZW7d4ARtgNXYZzwseKewXX568cuHzuJKuBfLT7Otnvuz
Hy70iC70wmfxYIG29KIUjhqVFJZ9RO+LE4EHwkexM1BRpxAuUfHHSgJc9qb5ltHE
knA6L8E5ENrkdyDi5lYd3zMzKuyVBuJRiNE0ZIxv8OchaCxerxICUXHgGsuuwNvj
XgCADimNLf1bcaptgPaTGcXwk3Ga2/QnFR0ofQD/+O7uP3O09VDj+ywVrrLUHiuN
IldAD9jQlPTag0zrVo7qxHIAl/QbgxTR4o2bD+eYD2pthu9tIJDVwyIDQ8+molQZ
5ri9G3p6+qSD4bfseI3PdYrR1o+iT3nRKNktyZCmBHm5Hi0j9/UiBt2TZR5uGNPT
19zdcY4a/YHBFsFm1tmF0W9Fm6Cw7LlGf8xmR0UJ36T6sdoctwZ7sJAhLBTBQMaJ
w90dcQ4ZsjBym+F4wJFALPcKOdpBHYXtVKDJx+FRpeWQW6+nTl8s4cVMgQZXP4qj
4Efal9PXwN07VKn3aNkpIrRzV8FIMqzTqLp8KdHC8OP4/vb9pP+dS5ejFlDfMmoA
z6BjvNBj90bVnrbWLf2FqrLLIY5ytv051Jmg4uGTp2kxKtWd2O3BW1kxqpjA0gBc
ITUn9+D7kJDKTUy8jhzPoByabJcpI1DnCWztltkxvVJYm3jKgd4JQctKwQiT8E8g
U6wPjqMRfpPm7s9g9Qma3ZMk3UCCO4clnCCI38/pGVUqj2quyTNt1rmcAl8pk7ru
5I1J4DBVKubcIlQYWV2Uan8N81EIyoz00hYboPx9jMgmAGijCw8rh/II0QYA9Nzt
Jj0VzSEor7jolrSXUkCbq9+/jiekhaH1+uSwBVMb0DQ72bQ71pM1rrKoMXQ8eFVf
XHJwUd+RlhhSpu0FNd7WkhvbI/L2+Gfvo1/R9iCo1eaGZBsr6kUGT78pWRbRq1bj
0PcIalO0IRH1LYIa/kE0UKjHX5rozDEvoC4VlaR0GRsiS8GdxMcjfIxN6KntnnBK
oGfw+QZ4kLhNeQ2JqVSkxDSXmRl7ah4gVo1H2TPkaQV4VNEVTwBsp5dN+iNbtoDw
8Te2+VXKN332yqwcwBfRTje8ugqYweyPnvQ+hF8IoilvgCJzyDkpv8wivlPN0Pld
fRxBtl78KDCkRfpyGJHKgHhYEc+dwIRHrmCrV93gBbdiG/R8A9hBgC6mYUtRUNmh
ZKsEX72Kc680+CGJe2q3yw/kDFfpYdh7/g+wiSoPw3g+3xfC/VU7ss4XR0G/b0Rw
JBERdbV+/c7XWkk7bsXlNs/Y1LB3dhxBsIup5PSYZWti7c6ImRETZob/Jech9qXG
W2h+3AGZbg+2PiltL66Ld2Tg934TNhdQWwm5avmQjiVg4uVtgYcB79np3WnvHmqn
1PaJIiVJm8LmcSZ5IJwdLlpF2lXgvxr5Z1xNVjy7275SxOu7UTP/qQv2WjndmCu8
3m+BTWzz2wHDLgUJucvnilV0wsivN4CcbkUfHvYUZkSocyX6owAW8TsehsHLEbJf
2X/HQO+DiF8ag1MhEyxioRbKseZCQDt67MyR5YFuVKFbCICN4IyIX2CLBnjVoROq
5yS6Ufa7XvyAPbU4YJ2nUWn4+fwMXdapC2rCVWzkxDJfgrbgXyJIWsNaPBl9bjHD
Z9dFRF6nsyHNoQksqOoo8IcGmqBctG2KRsC8s1c1nqJhRjwLDANZnWsdkTx/c5TA
aG0aEx0Yanvv3sv9JoKEAy7mmB/QxsUBoJy3bT0P4MfF8ZzpzJPfD9J1al1/p9nh
BgOLiD8bcQSPRdfGFht1YT6zV//pBPHTGpjydiwTrtYSaNdN1u0LRblKseJ7F8tt
6GLFOY028hfPSRDyUHyyAJj/cMlvF4cxmmoJsQ6X1ikoM5cBJfSwt7TPvwia3Y71
7Oeu+qiZHwTsseEsuPNgxL5+T7IVayXVMANrsx73QjcCSeeWk31OECcdDtpEdC84
QWR2vPZ5YGRAJJcfZ8FYnV3VO096yqpNEZQ4x60P3nzvov/y1tXFugrjrToR6va5
E4nSisJAlgEz3JV2bsNhEQpqtvE6Bv+AIcim93Is/AjVA2g4rvI1Y9PoP7FLGqar
KqCukknxRqANPsWi8M5Rt/3AXHQ1uu9yr1OqlzJLpy+e9ml13d12SV6gKw+el62x
gG+H4lCk6x4Ez3+8lQIgE2oDTzpfKcLq4Ru5m9S01LDjtNcb1tL2NTnTgkjDNBJ4
OU3rgvM8B/bNwCBBzrCjsTNfLI1GWnAkD8fWnDNgeGdSI2asiJbpUEdB0r+1oEDl
PCYTwFHiks9H2A2mgs9A2EEV/Ck/cojfCaTKCYzQgB/IOkuqenQ/P1M/VWCAmTz5
EhPCZZ3OpATeZ9eLaWGLCGiTS2j6cnCmhgaaRa8o1RPQn0O/RiyDbamxAdXDN3AG
gOorKKPkbtarmkXQeJuVAp5uAVh7aH5WPAq+4lC3lInYOzS47/O+npRvUMp/cXOf
/z9mFIiJaUf2cBJDkWMZt0ouNQj8gda24zuB1gFgxsd2t2Lt6jmryvvXmE7IsL5i
deBpBMWzGKG618m6n4FwOH1YrZvN0I6EG2hXNxHv61+IBC0cqLrnlZWd3geB7ZRs
wcGJ1hdLrAvCLfbetsoBAsWgKp9czWBBVmaYkS8U9yT/LHTe4Zg70wfpVURmE1jk
8dVLSDiqo+qtrCwaAS8TuUd+Jqm8UQzM29kDHULqxNsu/gFGxlsJgQL/kMztpeY4
v4k0iJjrIpDXU/o7toBJkYbbrf+zHeomnioBw1SZfDae/SNlF3KGBi5IUSyg5wSK
tmiiXcTTzilggC3Yph4IU8YS/+zdOwGArDglAflQor1gKp4olezION6dokCBbvyy
kr8d1vaO7jCQyegS6Zf6cbseMqNlwQ6bF1Zuu1NSx0gjGgvjd9xjOnZ3KwxWmJCn
`protect END_PROTECTED
