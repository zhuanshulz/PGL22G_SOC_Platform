`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KYhreHjfQrwvQHKeLHvnF1onYrbKV07NtQFCMp3TY6HNP18cYaraGbmerrP+90cu
zOJL/L+BnUr6f89Ufk9X3J7+uzhF6HADr/BGGt0TvIH6kEEgXd9SaxlptipefNU4
tqzu8j+50NTCVdKIaRwuFhVUcXLbT9an4OE4dgHwFDA4hXvkny446fN/yIdQI2Mr
e7nFSqj6BP/dXfJfWmX+oiSgy6/YerC3cF54AASAYIXKsL+Jse5nLltJZzp2suf9
pE0fpMN6OywQodpG66QuMxBf+CyBaPOAk7lAzymXuqFh0+Jw/9sJZMM+iGwG+hFp
EZiSGvtEoch1HTMRxZcLoLzpmdToBSOMI8J+scx/m9vyW2Glp9gh2X59tYBp9qSf
JiQ2mKMkd29/g61CeCyW60YsjLpHrB14Eg2UoeRHbTEbXepdCemBZrCx3Hfxn8c3
+HkU48fSbEnVVwXHwetz6U0eB29+cLfhzbRkrZeW3OFok3ChyPzkpFh6x5ZOJ7c5
tM5NTYnqK2lkkCH0BgHQJmim3V3k4m9cu9In9SgDzXJwlMSSWNM9kra452/JFKUF
wRM7wbrqWxNuSvOQJcH49HXBwMmn2uHumHEwNzdDl2rfs2EGarhx8iqYxl8uv6Ol
GFMLj+gvGnKWYpiofJpcYWLYv6c7Yb47BsVDzenEO2PogOdEJwGf1mbwPgfI+5rk
ll5krEkBwG1gOmZnfjh/NURhkccQpa2KO9iQbjqt/LdTQaFH9MNE6xBBaul4/6TM
v04OB6+QJdZXz4omzQpjpUjpgzZabxWUxkx3IwtdWzDRxjw/DnMAm57JRbywWY11
BtXeBx1YrmRXOJoMSJ04vTbfj/LmiEQIUqiDkKz7l7JHvRadcUQFwbqo+kK2PyBp
KWKBOiO/ScGZFrr1SEPVhfUGE6ugSrp3FiZ2IatMeFaL2xi0a8ndJUCYjTLrkwDK
8AJmUSKqNsdlc7NhGQ2SPkKPR9vbTHNe/p3q+Fk7BSKhRlYyGG+BAZJJTw6UWVJx
nTu2ARNBfgf0gzATIGltsnZajXPvIKq9xxM8wi38qqg1tj/c61Xv7nLOVYwOXBYO
SpfxqqUMNQ6pcH2Pg+3FyCBE9L7zaMoFnYhGzZWWS271NaBL13ngDy4mitcMoedR
oufVZ/y6FOgvSn11m3YrrKfOIgPUhHQ6LJjJbePEHES20cJoDJPFb/2ZQ9SPeKyl
YHguOaNva7ZRYlPNsfMRaKTHC5SoV1lrN+/sbAeKimpLZSrabzAW2ooy0glLHVrf
uF1ne1eJbDEH+G6qDc9v6gTVhYVjfI64P9XIwg9SaiqTCcU5ZWeysFl5gt/eVdP2
j/64DFOjwEH5KuiNSoRxnfOzzCggxGt3F2B7CZsHHj2ZczqLaOQU1v1sskZgJugT
bNXDQ4tvuiGPDxyHZdI4S/6eu6N4X1lYZou9HBKW6/iRAkp5XBl27clFOSZ9+9dD
PyfGvstRhyAlrJnL+xr46pZ3fLeDgoO0OExhSRyxKNMmAnmQ3QKJ70NtHwNyrv+P
+vN4eo9w/bPG90jMRSmy/EMXEJA8qZQagGHVrPh9Yx0E3WgjzNhKMykPnykXe0tn
5mN2K3RmbGJ4r001aDznHVTeYg0J26xVbWY8YcpKeTE=
`protect END_PROTECTED
