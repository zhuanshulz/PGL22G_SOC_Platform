`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FcEh6X9xBH18ADH2xSiUIwNxa0zU4gEfYUHHfjZX5G2bXbyNOo8PGdNkSlo4boIc
SANcuoYFy1rlMF3CzuzUQI+qJ4uAeW4ich6Ra05cdfpkHQPr5BU3vogcQyiEjT4V
S5kNpRt30IT3H5AF1QJjHLDmY+pZNqL4QySpckp7AD0Z1JkVVU43ECqYiINMcZj6
XqUrghJgdaJvaboP7AUzfI23HMBQHx3OYQ2mvzsDbkYpp7ISmx4+nAywiiCmH2jE
6mjGsdFm6JIZ3brpyI+P7AwV46mkRnvkrMESAF2uaV9uHFuQYXhwQFUr+PmoUh8k
E8ZcLMQt08qeuvjUBPLnuIAv9j+z6l0NUCSoPWCL3WngTmBQPSKu9RUhCBZ+M3x0
uZMhNIUcJogUfGJqbYfKoixVlGnI733tNXz98fO3UV8=
`protect END_PROTECTED
