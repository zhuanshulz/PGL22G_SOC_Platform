`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+pQ9VMgiMko2CgqK7DGxPqzEGQwuc9LBYGRhvwmK6Nppuv+mlQBesNRj3vmcZcB8
yKnZcbq8vyw/BEbaqwhGx8A5/ml9v71P+7Z8dOsKUy3ZHsE+SzANBiFtd6xJPx7r
XS8gIpVLTvARedaARlGPHQr/+myILriKug8UCtMgOsQfPhFlzLHjI9epsawX9CK+
fiN9ihcCQynAgL4ve/3cC573BOqk2K+I/iQRttB3e3ejUqH/F36MQ6Wrv2PwUUCs
vst18eSZfYpmWh5R+Gv+pQfjLXBLq7ka4VsT4D76OC1sW15c+RcMlD45Wqki1BLo
pB0IANJWpu1jBBcMpgdYt3cMncpKoQVdWQln1EHBdQLYYEaapG0znCBkUJa71192
BHmQFk3YoVZysYFz+VW+AH1nPVjXs3pCZmjBcq82mExbkTPBfZPyzjiVHTr9Vl2z
+LCxZyhDqZz91t7kiOjg5CU/CIiGb5HdGPuE0CVRsS394E7T2/WguYr9gNGyZAwG
84vjyvm34FrQKGZ0gh2mkGb98hk1S2AmFxjcBHV/vvyAcgPElrjaae2+5C8O8tnn
O3gr9gn16DSmkuh73rCkuPi0drMT6h0eygePOdNYtQMDz/X4S7HfRl3UVbQmgL2w
/Ym0JgcWb6k8kNK+eUvFVnrvVgfvGP6QWd2u3g5EdEhJHqsuYq8lf0igaVToFQz6
qhcFKliulM2du31caCIqmO5IJs7YVOMnZbcfpI9JOSbRVywbdgMUZzpeQ/ofxrbi
6ImdEY11AzCWonnfWNZUJsduo9Jfu6BE1KnwjKzC3Z8RsBiIsEQNba6i2UfocZo5
qQ8MmNWONxeT4Kn0zwkyKZh7P2MstDYK1GbrbZGrZb33q8Axfz8LPbe7+IxIMUSB
8cTT+59mIoplxcsvhyTochR78cM3V+XjMkYoeQnsWlkX5ZEfJfc8jPXoDhWac8U7
TpJ+Qw2+RhI7HqkFMEraHa6pgAKkJ7/zIxnuEIpUrHx6QzNqnXYdIqGQWrnQr4qb
A+uFJ3aA33sec9N+2jpIxH3D6131w8nEmmiXRlwnFrt1cTzmQ9jU/y8a+e0EH6j7
CygfPJw0t8jbE6aLyNLUNel7uA9AwkQRQWJuDrpYcJ12hSSPcDUq8fpHsLBD5g94
Uj88A9XVzU0gFyXYFHkSiI7sxHvWNBspvLly7AVE7HvTmY44e10fr41UU2l50TM5
iTUqCGVY7FWT8NBej5siDGkPbsozfxnz/6pSiDCMV1WoX6SUXOGq6b87D+iy6330
Ws8NA8NuDLJUiK6KbxJIlhFxFGrZ6wtO3pgS3GBjqNN7UbW2bv3XxacqGueeETZI
kTo6DpClvAjKrQ//7+7s2SbT+rIB/L+uGb88ssIxQag=
`protect END_PROTECTED
