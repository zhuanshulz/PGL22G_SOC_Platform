`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1S460S6qekBd2SzBvUL4YqqrxvlAz7ajSjlerBBSLPj+0WwzDlK7XkD4DcqGTi3L
J7Az5Z+uM6dwhk2tDV29vQ+n+PSArv0l+5xloUvWjj+ot6tvQmKOc1wwmNpz14C1
w2RKXjNVvtHuljp7vFnbnZHqhO1bRiqLt+UGASqOhoVQREHuO9BpBtcVQTnc8jd7
FvnNwagEEEGTpmPQR3fy9/seg8SUSfYmzR9E2He45RXULnDkvSDCur83UNi80pL6
d0e5PhJkO7QFrPcxz87PcJnFvkvgz+38prAY2IjFsixQgi8/hiEmLx/7jUotctBt
4TnDa23E9mRYoVnxiCeBcgJN3xuSrcEO3opU6W9P7UaOQyNUp4nm4nXyS0E9Qf2M
S1HKwkWXy4ovnhJ7FTr3akGGV0tKOILStx+eKKyVumSfH14JM3T845ZwN6iatYB1
8pAFVQcSOzdffRjXUFLoT5TkN5NrBlzdhwMGyO1u7k9k0ILbjyRSdd0ybGJfHe/O
q1Qex/jFsTW2eaKdXDjSjQ==
`protect END_PROTECTED
