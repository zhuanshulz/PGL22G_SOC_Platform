`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r+LyWz6J5zfqQO33pGT9Xt9j87QE6tWLc9y1F44I4/+5QapWaWswxoRDFlRXgIiu
yBhiqz7kLiMMM0QT87//ID5nd+5IxKBPtl8RA4ML+A9DHsOastlS62PPGdRgIv0/
ezVG8N/vAkMQ7LOxVn11lzrZMRI5rn4UNWtwtwZQHqnN0p2Lk2jGN/QHdPZSH3Uy
QIsJq2VKzrchp4mrS0wdjaDRnxPTGkzZ8owiODWea7BqVpP0fC6g7uW03k0KTy4L
BjVRTvQnm+Ds3+JYzd8UfukVegdx4txeLfzcwxgHiaGB3xmc5yfsU2dI2HNJ1Jvk
f5PQUU9RDBB9XWuA4GF7cT+OEQvq8L/2YMdm7VOPEkSwrvn/9kn0weLRvB5jOFNp
//kv74XiYilZC+AzyhNhXd/avG67yj/qpwabKx1dJKP2Svd2ptf7PuubK0UOoqpz
hQFET9It/4M2yw4noQsqxfXNf86zmfJkQLFBYDyUJbfEjrDngMZl7XcMM+xh6oOW
NCpVttY2zVwiyzqo4Sc1AVlCSlKPuoiOnOk+67X+Xuh0HspjeB4a0RoFC9epVzIq
pgyHafHjjJyrx6V3y1YUocNhoktxPk3Gx/U8Y+/L7o+0P2X8En7AMM6HTVMyfhp4
hsWvYQD2w/4Gwdl5f/3delQqS6cRRwGRA6gLnVYHNjZYpbKUs+mIO/XkmSkbinSz
GL963V08FdYH/8mrwJ3JCo0f3afDA5Gtyum6e5+D8smhi6zagHnZ2FzfTbkl093R
UzmJktuUNadzuPVIP0SwWEVp2KWxLVMTHXJnPlrRQ8FBaSysqeOmH7WzCUz9TeQQ
NyvfInG+LfgtcqQapc8FItzg0Hjuh75DWaoaTiclUWGQz4dIDv0LZ7A9DfhWLg4w
xLIGnTGM5FS+SZUH1hcEh4gmg3iwjQxHyzuMW6xNvQUfOcJISXEeSRLvI5LhJiGg
CsaJN++cmI+2D3d8/n/QT47zMQfosEObRPcoF9HyUXUrMWK3hSSOsci03J9ZBuw2
kwUr/6EecqbrHMGA7ky/TPE5x+GMi8+CAfVMKWfDpM0YzqD7kXMDApzWWloROPBV
C3nS4Z8NO8UhuYLzBMHxZukQrY9d7K8PS7IvElAfLb/O+fOy2e/0MdlaR6B3lFWz
g22Qsfn1zz2gltXIi7s7Etg0BSoI4kBk/XG6b/baDttzz7DP60cxHX9AO3MXjKZa
s1cz0Nn6DO0OH4P/gxoBo2NaVoIAYhZHPqhiHwvCpTtqUqzxsJGf++mmgq+la99i
hW43H23DvvLTq3H+5glX2HU8PyOQi0ZofobTsZpK77g+90ZWvADW/7ifQAAE0dIU
7UlwDUc/9QB6MTWt+5SMpyOOImLiqQfwZSK85zScBczSw25whZXqqSU1/SKbVYoD
ixmNUb3dmHgPYTvSkN0GJw==
`protect END_PROTECTED
