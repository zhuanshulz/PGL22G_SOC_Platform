`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e3NPrqJGcsKmvU4otqteW5D8fC85SzMVlWvNEbFt6P8GspvumcCovr0jbAkBk6bU
LgqFmYUnyHPQL6KgRg33Fmt95W5v7iI7TmxMBGkgdrk0gOhbkPq8kQjDQEwLl/Qr
GAAVr+AEXbYN1vWotC91xpOTysAu7G7YRSe/MXU2dFHpoS/DypMoOtHloh15KAB3
h9fgM+IT+QDp3jCIWOktl7LW2nY9SrxZKbltr7cdrCl5SAa1vJzaaK9iHaBgKZWR
KKmnimhb2gDigJ/8XgzOU6vJJDQP0Lbb2qo4XUL8ZM6mFMNDtFbkGB7S4sfCP4hh
evSNbZHTHSid7eKC8LL1Bh2+6SkNgx+Ye+L1KbvtZIl3xE/UqTLG8eLRIBOSa6ZE
V5anZfblH511W0EROiWCd/oRWPalM0fbowFvCHxAWixXK6x31OTy7bKiYUG4IJQt
tAW1gMR2zbmraBNQzyInzxlM1Sdun3oapPhXxb6fxtBoJBu2YdPdxl9Kz6imFeAZ
I4Ss4C43Fe1QIjWNis9iBtnH/mfOKPWM2f284c687o2OKEKx8dVlQYmQK9ALD3i5
F7UVcqDTU1st5ZmkTW7pNUatqqLjiCUlQkK306MsDZj4l5VLGhOMsVpwxUXe+uOX
5wiCNTdXHWBKMDH4ZdJeNQRBCbkDypfYHJhQh08NaxRQNdAiEkp8Q8h5c5urDAxs
C0s3z6flCjVCY0oiXGJLvyQCHqm/PgIpelJjDF8Nl8JK89oQ704IU5Lse2P0pMAO
VVqokZmCD0EO7qtaSOPl+6+TpAxzM19Sv+K9xu/6e5fEZLQsCV8JuTeCgQJ6bWkl
8QXPg9u6VG3dcb16UdEdGLrmk7MLP9nMkgF53YXkrp5gxjcfhZifUepuGlSU5hjX
Y/uyunbn/Bi2mENVdN56lNRHhmEW4KqByJeHWKBNSG+roNe0vi+Dnckv+rMQBEaJ
/ELusNaYYSPAJstDen+t8MxUZEJ2sBz6tuZfpGLes9NtEMtFF0a1PbnhjY8bHlNr
ouV7koL0dYnwGBwSX6r4OmBjw2MMxuXmGQqiwA+8RTH3DiLxKmqcOPzs7NTwUvyu
Twjtle12u58jPUlqFmS7Vhr9Fw+S26iNOjSLD7s/C//TX3ON7eR4wxwNe4zinH4b
dIataOTzW9j3vmpn3q09g6nGqVVyV7Ujd6OKQl9Y39zJGfD11ok2LzJ69MJIYL1h
+2Cf+f0NteF+Nay99tSIcMDKb+gkfjH/dBt+e29ui+E/fPLRdcXuP+XBQFKLsFVC
snIWh1P232T9KFFSMJxsVVNWUvzSkd4erCCESSVIAJYpAGIJzkR+KB+gLj6s3Klc
fAISXDPHqhK8obpNhTcu4BKSg2Hx5AaiGYpAghb3SsGOGGoju+3QuGbPerYr5jq5
c4xHyyMvyUdjzjyC8c6/uXBxFWzXmRSmYZEMROlPn5Y2VVkFCL0J3Ptxla4sl+Ef
vMjDVAO4G4K0fkQcqOzGQIcUeBTJ+vptgmxIOt3eVLh/6OBGNj10MDFuOMHdqDyu
lbMksyv9aA/pV3aPrpz/ThYolrTitdqT0h9LotjYgHeFul10hkwQ8+y4TbWGJx+R
j6C3Axq8PExE7/xdOuC7o+JcLKvTFY6nzBMjbxr08qL3tMWZukTcrseac/O3yO5u
0krltz28tW70e6IisyzM89n1BAX+zP6OZtCzrgaVRA57ZksmsQVSIKeqN7gCbrAq
ROLgK2eBx4RX/FVrt1ssC8b+n0u0O8GWBARDUUX5mUGpriFXln8PAV4/Wg4dTYma
UYw2h0Qz2Cw13q5HScEYztVelPFNZWg6SvE0w2mTrfLRN3430QrtIQg8RTdIfxEm
SpYUmdkQPxPdTEMW4mr/28SaDW8Ww8qBVa2Z+n21o3ZHf6b0km/C0FWP/rp5RqS9
mLLH7Pu6nRyEAjz2sw4H9xYHW747WEm6KvXv4s07jJb8RZqv6PrPi7jKFB7SxTDN
mE+EOtAud4PgTH60JuZXWu3Fp70Dy8fQEyHZV5kvf/Zv1RYLzTEUVf3hF+DKW54y
`protect END_PROTECTED
