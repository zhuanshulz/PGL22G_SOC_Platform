`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tp4OBBdjn7tbnpdgyOO4+xKsfC0oyfWK1UxrbMTyffm+gjq2dbTJgyWpGmvcl8sQ
ric9jtYW0XWi7aRQdINzRqlAkJyihaCkR/yPtL72wiB6p6tPFS8Jki6vH27my+MX
o+rgZNkoTXC3h8amDToRxXTT0z86IeRAGzif9+pptVpU6xv7Lltt3YeGp0Vbd0sQ
vT4630RCOGCkHlqehPXKqnhTmfxrKVTeMFPC3H9UCNh3zuF8cebzCOnxDG3ugEI4
uUIDgLk91Vqx3CRgt3TL4B6CK504B7NvO0IIkIrD+OlcN4tcdoa3Xobq8pBjJ0VC
VHPqwOTQtBmT0V0S5sJv2svEmItzzoiMg9hWvY0NP2E+7Sn4oegA7Otar0UFHMyQ
zLMK/EuEeGlW8gInrPwuaBXyNCBn2thqJM554Juwek9KNCAoumRv87owqJVuWblG
gLqqKn2GXFztVmp5STovvSRo94MRti+v3X/EuoI6ZLeYYfij6pw/LpFthwfxiWYV
S8IKUlk7NFKbqF0q4oOhb/C8jiQX0meloonQRZmgWbPxPQm02ZU0s4etC5hBg5lP
7qTSm1DxbQDnS/TCWoR4jC3tMx/geleuuREmkTOnrzBUgnXjigkyraXETfbb5R/n
sjKwP6UBG4F4YPOKBy3l365IzeS0BQn+AJ2yg7dkMaJAt85Y3Fd5TGYk3BN57hjj
nhrapx09dBuJZymUatQcRbe9uMbcmu0RvK92nqJCl2id28E1XusNrMm8ln6u/iaQ
FFGXXluq+rEKTds1oYPwJLoB2yHwnRjnOWQsSsR8R9g32Puu8RCSofCL7jNXZV/F
cBKfwNVyI5DwVWgP6EBjgJcfG5pPQvjrntAeEY/tVvdac1Ia9/eLd3xgcG87AgkH
NcyU10L3ypVMOmV1clGns2HedGdQWUOKQiknHuTU8d8zcfCdByw3cy9bfS49vH7a
8XEa+NepHLYHKHBR8wW4bOGC0lI+GYVoBqYdzD0tb1rrRWti3noNjB10lpCowgp9
aSaB+gda+fADdr7wS1uFg5jCAIJjpMGAp69eq2rYa4z22XKsu/bqX0ByyYVygGr5
kG/gN9czIVvcvKMFWcPMsSwAwmZjX5v6rMOT2+68CJf3fHTyZX4cehKkBfHcpTHQ
l13d1iHlCumQwRM3FRjt/ntm/tDdhPUnFWqh8Z5aNjCFBul5MqHa5b7OIlooYlCK
n3Uvz1pxIVsQFstfCZYStydvHiPJq7pjEIiXAylzF9SOtJqggQbYTwA9sFP+iFcT
ls2G5vKwfY3kiPsJBEenQS9S/b5Msn9lzg2z5gPeZGEkF4cjoF112Gsfn9V2LpmH
cydhCREKQTmTbGmGUhazmZMKAWA+NzBSiUmLDbcJTEMw9hahw85zr7EYopUesmMc
pQqFG5krqnmogpRkWDIDp9W1S+iorahuZB0gUGMk+QOX2ZTo94JHllLCWsWAQ62a
/v2KDb/EmstROoqyZO33UlpgnoEDtd5ykP2BySTQiSHJP6tT3R2QqiX4et8jJfl7
8ILrvUlUMiqafLt62/LJWCTb6ta1AhITr+taU3kOBRlfp2d61Z2cMxQN9GHQPAFg
02MXLWHwbKilumuLRPN/JKvPBKloUnBCC//QSXLrpDFmzIu9p+eXAEpcEwtdSXXV
wkDkHkj9M8uGRInbstoWVvgK5f3Q7Kb8/HBJ2ytkAa6OqPx4Ftj9EUpcdYZOiicx
L9/P7kcsmPGI+46Nrg0VagQBwhVYoRD7thJunKehBzBu8yr11QPvx0TyfVdYVUo3
n7E7xE2XxHSN6jwKjTzW+NgZYtRgz9RpddXlFWVhl8i6drr8oa7sHfyaM3WyCC8T
0ihLz7zmpn15IkVzcu86p8K9JdcXKfZmcgCIXcZvevkSSNMEIq6ekuJX11Ff0qM6
6FyLMAhxHb2txhrq8ho41DME7dpVM8x1nXbHD9WUJSx+u2xv9IKYw2F+5EkibtOz
uIpVdXDthWqjjSWtxymz1TTKFqSv1bAiRy2UJ+TXvDVdUe3yabPSkytHVl8KoaUi
FmQ73bSnmGcAbKF9P4zk1PGETH4lc7THjgh8zH9ph5wUqn21YGuDW4zTVEj7K5Ke
6Lk7BBk5M4UyZyQXvUuuuc6OXB2eHwItv3Q8GgxuBevCigXSLzQZZJ/vWAeVX18e
hlJexFU6H+Mispjcrh30Ev8hX35i0DZpB4XhGwLLfKGVn6N+OswHPo4ZBLuUG4m4
yEyNoYSvp+t2KISHx+aqkByBXtP1datFA3deRi0k285+EKVono0H/HWVcW5iBjhp
3a++EPFshYlIC/gLuWSVblPmnPM80Amaqu/dW9GGYP2GNjBbvwT7Baoh7Md8wVM4
nP5zIIMvngy/MJkFbQXUewja/PmagA7RXELHgmG53jHRsQ1qORGowC0WYoTy04FD
lW1nEaJ+s/SD8W1uuTVFah2Qjp7EhUnuWEe2W5kNX/vjCx7+AU2HPCbcIjxJnqOz
ed/zeMuzlNFQ3CEswHwLtbiGszw+DZ4mUV25pP/kK+qxJXL/5iLsIMYTKcZGqM6v
jRjHJUeQvClcs08QSWEXTcues6BuCrw1wIvqx77sRv/bmIiD0dODd3c4oinL9J8A
4dP+ltVp6COGPDWVqFZdOf6zBpf3JiG4qRk5z2PD9LFjGq+aDn1J5EU1TLyfjgJB
afvA5YbYG0tSaR/Y78ImmaaK5j0rqt3/n9DjHKWyI+YCmxtth2scW1ocWNs8qu+T
S6ZmMKuxIbMevorttVOOdMspz3erbmhcUVW4RLozeL7GLO45WbMSBgFSL8gMJ2rH
mVXbdoezQleNBiSN6clUI0v5YXznPFDn1zQY5q7dzknzYGalrLxHH/E6IlbSJXbo
P7/eBoRfYmLBQxAv22gmFaPmCGkXLkZ3V+ceH0XKBnJEfqX916fJd5Ol7YOwmp4C
2tSGF3qIOslRyu+v1cLpYCg4y+RnGjtR2+2nd7AXN/M+BzHYQwMIpZd/z7JrMzcU
lMKb11kIUtH0ltGu/yw9fCtCGvSqGfQnNhntDD2PJfQr6UcdwMjsHSmFqBdjGIws
c5MW9neNv0R4lhYo6RQnI/L4xloEvvftcgREqLwcissDl8/SLfisNxSVyd5sBrN1
XKZ7nZ4eCOtH9wcg2JYGbwk+9Jedk3/I57IJtcPx0Xp1ULWjrqyOCALpP1XyCIH4
kJO9b4sBerXt4qdcld6BeHU3EbgaByqFFRmmRqSef1qV58Vwk9XUmgBRgQCyhwRc
1oceXzqszjle6uUsgUDQ4IpovaXnZlQmmEpvh2TyoeUrO/rJ+T3Dlsw86o2asnbI
yBOxIGINTuQB1iQv/IpteGQMOpb2rNsp6RnqtBybAnk8n9875qcdMlgsgWXp7AFo
opW9NRj5NVv90aZIP0q/tXsJr1GVahaBKDl/ywnXqNuiG0NgFZUNGspUJOiGl9k9
qognBhQj3/YrozXhQ82yOnvntx+/M/1dnm2zhH65MBCXP7vzA5c8FEte6eCvCH4D
rwCI46TcpDBEpxAAHZABt4letSW/sxflX376DZBjSynuu1SyOgvHmbl8P5uQxc6r
9YZMaamlWRY0vDdn92ZO7toMSRclyFAGEUBbzJfNJuc=
`protect END_PROTECTED
