`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CXYuT9BVb/G7jd3bIzx84OYXmAfieO07OlIJkT1HcUgu6rHCqgpMs8PfMVdjhznC
ctP72h43DSBC2M2ouiHi9kufYO8aej48OQVLA4u8llvhsu28C8jAmexbXiKmbAAx
QUxUfhocSVvugkn6C//1fw4eeAWgvVptj2s2PVph/KhSW1MDd1eaLxMHGi8aSzzi
MY4pkjbxIEGRlNzZIJHtWroAdKml+d6tzaxOu3FyVcFT2BVoj5FPhSKLHyUfUR14
ymwvCbzf+nRq/FUghSgvf6m+aUgQmjzPR3VYlQr4MPc=
`protect END_PROTECTED
