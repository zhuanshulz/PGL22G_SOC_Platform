`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bVaZs8qbjZts8DT0343XDwP7NIItbRiYpEkPKK50RQlvvCFcx75o6uU91K34J8HC
5JfeRw7ZWfW8PlTbkwekjkbi0MnuWTj0F/bPQ9xQcdt1IMFvj8uebUDdiRQApLSZ
/X5YdjlagAbvqlnN8RNPgWc/GKJYaWMNICebRqMFRyV2yu4M1hEYl0I7QJ0EOdWQ
8GYAyyirg/kYam+NRHb/poUz2tpESkkyZ7rKJW0QmDeTVRqWxcMxTBvLjgsVupan
AaAtKd9I3Z46bWhAor2h/dFEBx8o4wg6DW/Pf0TjZ30X4a5CeBFTtZLRPpiCHBuD
zz28n85Cy35ouo2YtYfDSPD6FYTfSizFy5Kht6NtLEjKl4LHQV0RT9yIixdM3o+K
fMW9HvA9WUYWfsf1rVGyA7lN0UMsNDKVPfvKui8qAt9TCx6MJSrzjpdwjvRaaQbD
jlHQQkRa3MPDavU89Xemh79QEtaxClCl8F+9MIYODVCgRPJwis11q7GQxtO+zNHC
Qozv4UGOZ4cDnhBxQUWR0eAlF43wewMXwVEPT34FHk549rPKOVv7VT5OSUYv5tyO
qZkPi93ggmfvr+vSKaIORQ==
`protect END_PROTECTED
