`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fSr6rNX6RxK0Qio1QUiw+aNSjHbvMUgE9qSt0YqSZAfSlmuN74jIo7KNT/7lhQLX
FjE9F2NSw7a93qzqs4aS2WvZJtNspquwPzKy1+9SDrwJxygUnM5PNkCyxETTjPvC
SOhJv6jwJwCIimwuqtu7Pw5fv921/GQqpgaIa4L9pyOajupXykr1IVHg+Sw2jqm3
Ie1DfiDGvC+wVyI+yQCZXH63uCqRds2FsT/+3nqBi+pixGLKfQQVB2IPZg8LYavD
D7zdq7SORBrF0S/iK0uW6yeWwM/9hvzBAYem3DHXg/wjKF/bPnzDKs6h54FII4hh
EwFS9jnf1xcTnpRcC1ZlYpugxRc8QzpuNymvjxAzn4Oqd1eGH5HyvXJ8keriIT8N
IjjzfvFqh4d0qK/xJrLcx7HR9B1I0L+jWFniMjxrJBe+9S+IVUYngegA2nidzLLn
Av3QkuFgmSzpb1y3C3uDm/p+wLK2pQJgtwqJFNRnm2K1UmJECqbEHI32XC2mSHLv
l9doj9U1H7LJdJ1mgtu1Gh5Qfp3FMI6FbwFjudDNE9el7A7Bw0OGyYIQyDXtAj1L
woOYh5bKzM0bqB9z7LZqbiGD4dalInVfhH+WHqyQIzto+USKjCXHHEP1ihPikwwB
vt/MdvZFxmPFOlN7i5wWmg==
`protect END_PROTECTED
