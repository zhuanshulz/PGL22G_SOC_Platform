`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G/N+/IL1ypRqRM0dQNF1bhVJbOxyrS/lBPZKJWMbTazlgEzzRbw1oAAjaANJXWgc
4W9G87nDLiokJbOSg6J/5u+v3ylSGdnI42ALe19cWuZRIfNzmY0BTHI4RsG9Knxn
VYzJdzX7IXVubcE+iwndJX3FVAX40mup3Ew255C0+FY1dUv9YoLa3JbKcFZSqQQ6
kMIFJAnXDgm/BMgzGzY1k2wvzti0QfD3YbeHRbETebIRWXvgpm0vjr7d2rJt207W
633BSz8GfZFSKv16/C7W5wDg4CQTOB+J2R3/QHldkyoCnJY9Pf/IUmTPQvuPq41D
ybLlqY3lynTdaxk+xiEjyKktkDqTJRC2by2GStloiR7iw3Qgb5WH9eiGAsealt7u
a45z3fwroEK+eZVYMKGCod5ds792IGDOpAXkPBfCYZ/+y+6SthBrsEqIzLGVyLjF
rQvqOiPzaAtXxlMDDY8MIlKhsy5nCbalyG4HACF0QvbCEDX+SkTQynTn+t5SNoxR
hrmRPnj1dtTsEwkY2VoMb7ZSaQiTEvvJtq9VTKPTe+qen0XfV29YQAOY/RFUuhQ9
u/9Ji9UPX6vazLS8AlRUQIJ4oO3jUNlby/aQnvwBO0h2SVIQcCGvuj/e8/ApMK+o
/quvGKfZl1D6s1qgCbIASQcKa4wkg5Ny3JngpWhV96L29E0iC9lszg0BrUDYVzSm
dWX7/a6/rCT+kFmOFwdBlay+JUiOZROTf5UkzgQVbCQly8/vs9i56nso88CAZmsu
V4IvHd+HeIUs6qE7n10WZpQusbtq0SG2IzVJQZFrSZgD/PO3/3FCFkwEmSgyN3zx
kLtooSn7/C6/PnXz4rDgmHi7hmYfkPk5iPWNJ4uNSuAuOi+/a6mbKT7vBRjmORx/
tC42tE3m7O8KJcm6WJK2uUqQSpC9EAFGAGmV8ywq91HiIj04W9nHP8VkbOaa+zZP
Vh/emAJXEniHZq44IcYIiHhoB0Q8JeYaL+f75FPLL9u5NO/48Z7dcVJ4huW2OtFO
GTV6qc0PghQOQwwOXrDn1PZjsMBI6huQBOsUVjJZCOueN1/lNmeG3v1wAmAaun/B
w/KUPs6p1vctnhOi0MSpy0+/Or7WHi2STkXgzhfEJz0ROOLDMo623jBBk+Lj8gDu
gyM3S04znq0deTZ4TqS7zzYziua+qr8k1CDyoWRx5PrMMAO/oLz1w6cBos8ldAEr
pVf5nKuu7Bf2v2BZuskFba1g2GL6R1SAB20oi0g0b9m13sVJA1cHAqKC42ZoGvz4
NgP2QnE6u7zSkjaY7nTRnrCAGbeu0dcwVY8aDogKxvVtW6bO8A4XCeZnS0E79dfd
AYd4hB1cuYRo0VjJCYHmhO5zFRrTL40tAJv0zZgZ4CQ4etMZwuppqdtFvAelJYQ0
QWMC15hWakrjXNDKOTkLkdRIraEUBJSpyn3O5fyL9Kq4sMtOoHOTAw39pBL3qvxq
BxhLBYnZm0xEJIf13Ksz8s1UDHhT4yghmUdPHvA8vdcttd+TwzIsscasgnoLxQnw
wcnswOGNpozW4DNjIORNxqYe+UWco1hgFWMVeI8fAnZ99cJf0BzsULaezv0IkTKn
xDYMsl4Zj/k8q8AQD2C0UHY+KqEn/OShSeMhY5MkxwPhKIx50VSpjzh/iQAXui8j
GMqn4BKTNnvLpc54JOZx9jlAS/Ir+rIRWJRIQCJyScQ965ybm1UeXIa9EDEAbluC
PSILhlzzFxPTeft5l1Ck43U7NryzkNg6jONiLU+FHlwxjRif18MM59zTuEGlu1UR
YnNENdbuOWsdTqU0/vcIqh11BCwS//BwoVhi5z2iYj8FYba3qTXa+FpavDoBbKDn
ZRlxQa363DweHe+6whHiC379XUdVHQuERVwS3i1Ui0ddOeC5GVzWNa4kA6XCmUZL
MWExkgK0lVI/F1NcKAZ5rPKUeyPKzbskC8qJKl59W1wZhgejOJno+kLi0KE0Ojd4
lFmzbZtm7eQEMUt+0GGLlTfBRna+8MCkxYWRutnbMxROTMlFJw+uRLJ/t3Yfwb5H
2pM2YS1IRSlcs0qu4TIQPznSJZPa8CecKB0likZl9AWNdAV/Zo+JLeNbJkK2uu6p
jM85H1MCg7WorXYZPZ7ezMUBpMThyPaYKa3qrh9iUkGOwXBjUrqdDf6wPb1FiUfW
NMBSooqU8ur2rCjG4NGURGK3z3StwunElXiPUZ04UvH2KaOeV8UfMkT4c0GcEla2
hYzmVI8W5rAWq1mV3W2DNgw9fBTCeCznbUfk7WQDn7C+UGqn+RL/7EKXGal0nWD0
uZHdr8TKfQMNBh1n/2Scw6LFrXjyglyDMxVUiBe712F8VXV3RxRNhwG9qfVKFlWC
A9FbGrPhegnNq4ExK52/FFKDIzP0LqO1ZqZ8H0gSXMeHjETp9W7zM/HDtrwQoM4c
a5B/AtLe+08/KqM+LrNOLBUQ4QpIrKd9tM5LldCy7UGnXlUylSDXFqVRg6Qm/WI8
yGqb3GLR64KVbhvbYp2qsguBiZtiyi2g1S2Gbte5b4ADqB8x16LOcprseCkD79Tm
M4lfpMcZ5bVcp1LSUvPl2UmO4Z2wK089GI7sMnoqH+YTZetGBip+ZMnLJlDyiMPS
jWZgKrg4n0pLC8UIivLfsvmKKIob/uFz+yht3JJriz0OTw78F8avSfLZ+bWELhcZ
FXVHbY3g1FPjmY4H2yseBnwNHb+ylzv/rE81tOWj9Z2nyzEF7DrH2m01yhmhYHHK
uIwYNCiqL/Hub8f4GcI4qcoo7j2kRwZT0mOzL9UhhY+nIjtDz7vIv1mdLBtBES0F
NfiP7BisQ+gQUPeV9UKaqhCY5TyDfrnJvzz/GsgfwyDI8WHVTjuUQoskll5Fm2Dj
gyEEyMeAMrQ3g39pc7fwbWbW5/HzDiRL6bQCPqd0lak3C1v1YQ5DdFZDU5IzwX0P
CqQMP55C2EnelUdt6qfRiMK03gRgIHx37rFeAK1J4evT1o3RsBMBAWhi1t3JSgpx
SQ1zXDh6oulabqxa03sWr3omCkzbljvHywlyVZ2wVfUzzCFCppTRPfJzK/b/xjd+
jvsWkcgNhqYlzuN8GJEhsZyaPdcZBnGJZzZBmRSqnLrO7ZyNP1e9qppHh9sNGG/R
rTQiztrZdZ2Pm9hNV3CS7cGSnfSEPRXOOg+hfsvElnRmXCKfxoBKp4ZhSHrkT1o4
q+3xE9xEeM6CSgXPaxsEgKIDsKroKkIWSOgo53AgbDWw4qVOc6Y8WZK2zvrW1eS9
SVruSDgATQlB2XWOkuc2CEuLqc6nhA85On0QC5HPjb+CDs7muxA3jPoRjGwzEEC3
bsiynVt1qeNc0OuhWZQ+ux8JxvxqYD8WZ1uMv6VjSe4OuyvXq7naNT4abiBfa17s
uF46HmjW2Wv2KAr7o/C3xd17GIeyCoIOxFYYcylwacv9tEtH7lFE8bACIs60PkxL
S8wemW+GphOTyGjKz7mfiBaGW+ntAMyUEFgyE5Ldc6zPApFn/oHpVGUXVA4BD+KA
zyOaOcRVr3t+dsvabe/npxPBuBk26+6vsOSbwkDDLHxvU0qYTTxjMX8/p4A9JGk+
xP9XT410RZai4Od+5IyNrw0cxSTeu90JzjboicTgLQndZg1XqfvK0u0K1mP6DIld
nF3/q3PA/gwiXzm46MA+gmaT7McN+aXVd+y9g7A3InbcexR2BsdtdTlCBA6WbnyO
3fOl3nByuUVmd/6Qqv8LkQhiuBojzjo3xd9zpdq+2fURNoFLFKug8RE+RykS+HmK
NSGilN5jzGB/g3i4F9yKcAjUlWdZya5F+/MKYasIBAhqJ9AZh3U+y40jA+q6/h5R
10hxCuF/VYktHbQUxn5dKc3uR+7A8vXQ7dVYKY2Uax3+tMo3IoW7Ajz+UANIwB28
OvAXMkgUhc+KovD3NlL+CeRzSeQQ9sZreXTTM/XwZ+iff7mZb8ZilJmnOZsCzjRY
c5Gjc5P/2b18JGO4Mc16CFhmAo7TkaF4Dhl8F2B23TjQq7wPfOoKvG37nqKn/A/L
l9miA5GwNG8j0gGVPj2/R5Aa5WCr1KQdI5JIEsUU47+qnWyhiFRQwRD/WS4yz8qr
r8ByL2vXIgmcKE/BmsRHNS2Ki89enkga+8KXtb5xhssnGq2Nceo4E3rJj3IW+3YM
+pYPz+tg3DRHaNl3WfMMv6RmNIUC/FxG7wGnTDBQnbBezwGdisrr1f8pVsvERx28
gcf9xqI64Hgg+kM0lamSv1Izy25wNjJ28loPeSav3QtQetE/sqRZg3vDZ7amqBa+
lO6A0to7r/5wbyywYz5VLDwPr/eaWob/qsogGlnlXQwwzCLszr1ZWLJ2vNFeYto0
d8nW5rAR58LIkW0ommd4qHDj23+du79sPrBODuNB6QKuyRZpQ91KrKKByxvMOwnj
nSqJk98u49Z9Bc5OG82zVzbGx0Xh7PZhlKIpX01tn+6F1N8pD2V6GSK/+csxOBrp
QdbuqNJhrqh4bh8NmRf1ILt0cGCsMBrwS335WboE7mmbxbTPfjSWwP+wPEQta3vt
6/fBNQX3YC6QXECij65bpVnyfvaF6JlHGE598P694MWuWhADUYYCSqw31XyLCAbZ
VbGZYoUvMF3PRJyeDtkp/ZagQsCBi6Kze7jCryPQO10=
`protect END_PROTECTED
