`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zbYJWjIKe8CFbDpqvrjLlycI9C7VJG2+HfLbdB8XjAxQIRQwkuSHXACts5udjAOL
LolL6uCZA7l3pwp4zrzflEhu22OWgzF/Lrt2yNFw9uTmsuIx4d0yF64TADjIgM3P
1o+etBFUpSMQJ70RN6klXVe3Cev1urU7VObFPolenLXMRZ6b1pYBDjZ8xzubR44b
lpbu/D0VyjVG3Kd7GbiPa4c4kA6zGsdd1aSlo+t/2vzPLi1WW10Kr+PLAhAfgdH7
OE+cpoxjSy1QMyjvUudZciuGRoUDzmjW8tm61f6dvSBPnunLlr8x+SzZxSPaBABu
R2kQyUIrshFkWbGnfVyelFULj61GYCY9CJuny/v22wm1z6rYPtJS2WLvuKvT2iHR
uevaZeQtki8pW2PyxnJjkL9FKL+xb29UIQWScMCZtE2kn+iy4inpV8xFBl9PJk8I
NQp10V+FoAxPuYHpy6wYeiLA9+1VPLm20SZXhYhY6tcbl0pmsVaee6MPcUVgTdXQ
a6Ra2Fttut3vVBdCrsCA51RkEalbmCmuPjfmiL2zG0sJB6XCNiff2pCqFfr2BMUh
gcx7fiR5cVbK7qheyFiC5bfsJQASUz6muPWg8l76Rx3Xwvr1B0VZ8G6wH2G2Ilk2
GiVAxd3hZL+IooGWTzPOwQo8n9Nik6W172+shLM3czEHQtsxWFPZ5Bw6rvBrildB
a23lDQqTi1BQ9BYcjj0Jpie2f33kvWeU9CjuoX11DEokGDKI2GjvnRPqrHmcooFq
1CpGRF51koalxhxeFvYvGrBte1hwJm/2ZJ6fTAusVxVOBQK/NNernKsrwXnugCHd
gSJsQLPIO2BG7m19mBhm66bHiLbd27jXcGKIRlFlfXZn6uobsBgJ8+UxOflo/274
jr9jxNkthiiO3kgnUKETxgDodJ8/pjjHFFA8aZhetgGl3wlcF6zzJtpZ7+ynzWYb
HeiSkS6ljRUrOKXgRjuCh96a4VAAjfVe2yl1QtC7G1A/tIjBaEeTqO4uan2BIMNb
d31hD7QCFxpb21zgu2+lYDovqqEFK92eUVKlq1xT9TlYfqhe79PEeuMCm5eabcAI
/xTw89pQKmbbZRbEqrjnphWvf3JvBTn/QO5ZPIuLfTLIWnFhpXUOE8uqIqE07YpW
jAHQw/3zr0F7XVTPcDqvE5S36Fw7z8fjoL9lsz0iSL4vP8+TzGqIJ8NmrhZJO1n3
+GYhN6XSp4wMXhfYbNArWjuTZQXQoSjS8ZYYwT1dQ1GgTu1ZtsXALLkWiOO8X3Su
AojZqkxSalLO0j+RJUS0AcZXbIrXs8IpEv19f5xyXQPuls+BK5x7boaLKPeAfW55
JzQSYxNU0YVMM+iAbHtaUYH65E0ZPh+nwf56ecJ+IPTkCv1GZtL7tg6r3RI3kjO+
5Me75NPkD0We5Uufu1KnBwG6o+UN6UilWBoCI+/NPVANBhlVxrWyCQGRrfKgsn2m
631ES27D2EqLF4GFGfu06V/wH+hTCQi9+QF0vagsxAt7DBrvEiJg83IfnnwKz7oO
oOEJFuApPUpUC7tzE96Wm4HqH0KS3k1+qqIwCkjvsDSu/vBBIjpng9cM7oOTZ9Lu
4h71rHmcPfPjLW1O/0nNTdGbCyu6ErhIRJVxo97rZVikslWa7TnK1zdOmVdp0yxV
pkq/mpzjhfofmLFdAiqfmV3qYTeIhifg3eiSz7dNkOT2YLFH2RI1h/AnQxpKnxlx
HMXtMaHNffeNAePxKGvuNUMob1WpQhav+W1v78HamqVvKzSydtxTaPiJj7bqjxNX
dhelzlPc8nD4zF/GtOw0ODtup6EDbzsdYVkivbGoooE9vMna3S8dqfjcKiewgUXK
Aa+lngRihpPpm0USgis1H1WOygA+v4ulvny0EdrORgqKIbitT9Oy+TT/GgcHosxC
NhF5eK7d8YHUjoTCZIqV7uubrY4w8PhPMae6qWRwIjuaJN0/d29H1LwFvXUNDFfQ
aB3BBJlQm1NRJuLahAkbQBvyudliVkPbrZo2xoPtJZMuITCnRRfDfrlHNJUw3ybW
fEkRtMcuJOTKn5vMvSq6XTVsvXOpjJDFFDnEqJynZuDeG2qpNXPmgG9h2MGW4JFQ
hQ0DDQYoOjFfsgd5v0vuhW7Ehp8qQqe2kYdqw2CTY6OGL458Ia1r1DbrZDGvy0Vx
mVW//1hiN2rCsLcAzQaWU3yzAUJO8I3l0EUK32ZoBlyxaczUHsANfwtYQlXbeSK2
CoYuHCJoSzjWnQd7FfmAW8/1CDNhb0v4bW7O6tCAKDhgb6ZKeJ3Da9cSZFejb29L
8n0yyD5/yH9IEqiOUdPdjg4NRTwEylbE6k71EqhFEzV9GBmB1cG6/YxomFtsuta7
nHED7fcn6z4Uw7IDlzCzOETCwgxOswvE106lQw2MTeNlnxYHhoE15iFw3nPKlTHu
fsRwo4cBCAJo3jDXP+9130/3n6EU7b684KqV1+sEiAsSHhuoZMpSKoYf1/qSSKQG
KB485WWMljlRah66GiXCsS2HDJMqlwtRoWpBZs0KeQZvCBmFa1/cvfEgTVisrH4V
QVtUbTIugK5/MPvJnW8ws/h9PDBIR++f+7yiwWu5Fjy6TtwIJF2a6TUfzbhi+crD
evTN1j4LoDVJ9Ebe63dsbuMu/XVOs0q6sOy2BfyxQsvqD6AI3fD9spF5CqnBhv8h
v5CJNvu82xopMZVksLhoFqQGJRTdhmyVLvmq8BNkv91AQRYsncGRLUhSrc7Py//O
RnnowfCWQqKEe+SFYlq9+hpeHpqt6ucYZiZwmPPczxZ9mU7OWw6zSSRel6XE0E7O
1uIb4EJmZv9M62C8cFFY7BSdcBvf4TnFntUEzAttTKvn7rVmTs1KT7iIRJK0HV6p
+F9KN1O34I73szb6Di09hch25KiMIAHBs5VpEaS3PeBCkTSlOSmP/NniQ4QxYy0G
ec1Z4pndKATFakSSbsJClVo6/wTDSXS5bxCByyHuauylYMboF5P/ynNgF3i90o0x
blZrbZVbF3MSXHJf9L0c88uI/hV8BKGxPfZQwAi7VOmZYjXuIQPZDASNr19es/7B
kaRARHw2bbVWXpRvi2zSZs3hLWmwgfdFs9/J8Of+2uVkPlsR6tuqvdniOPrNymxY
uzxhWHndG5CWAqbWmZkpDSLFiqDvFRi4w/N1nk3VkpFCzSqgWeg/dVxR/5IIUHZ5
EgVUUBCXa2KIDkWTRHSXlCRVEWmOjPOHoqUxV6nScC+2wiFjDpctR6JPtosxr2Cu
G79wUPln8jvtfQRkeubIusudZuBFR0lM0FVA/viODL31uuz33xtqmMLOcYq6rBcK
`protect END_PROTECTED
