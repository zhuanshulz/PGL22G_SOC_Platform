`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
of/4gm+Af8MabwnnROF0ppMIfBCymhd3LGNB/KWaLztQNsp5Gt6mOlPw8E/l2sX5
nyCHEg3WMUc++fn0hcSMdSiDi9IwxPUiE+aKmNVrL3ExobSJLHeN+uf7FT9VVeBB
ivFmseIDt8APGrdPVHtn8+Qv6GVhGVRmJknISLFiQTNpAQ+VeLEdrgbjQOll1Jyf
jirbueSx98BiphZnZ2eH/NU1ipb0LIsTOwriX545uRNSXCFFMkW6H4jQ4MhVQHSm
ZYgGLWOBaOYUo4PWsVR4daUqRrC6277kFC6TtiM2pTlAqhF7infDQhRoJX/vNpVX
kKQ9eRgXKcq2jKDTogjYc3EEd2I5jxha5wE2OqirwvdZ7+LCbks1L+QHGFO4bWPC
MQtUmkZmy3NCpYilF1Bj9YZ3RSX7a7rNGatSSnCm593RByFJEx3Hqj4JurDrmZHw
LLkLUq10QXDvrY/yf4kHJXM6yQMRevk9JxN/87IGG4jr06ge5NY+0ncZzXtF60ib
sDDzoYyflV+/gcXZ/o/UMftDXiOXQOhApYspirqmBW/whWI6p8zZPh/t2sIzfkEW
orOd7wNt/Bk0t9pQ2pXZegJ2XGojMhG+oY4TIHJB0FApp052Y3wTIL6sgGWH431C
DItSdzKhK9gY6bIgE6PINilRJoYb+IPxf0rYFDIXbkrYutp2fNF+3KN48YUUCxBZ
pT+BKURixF7Sq543e/CRkaoHVy7rAU/OkD+b3oMAYVZ3E3Vm+j6iRo3eUfWSvJoM
9rio5sLj5ydV3OSo7xi3VbHbSZuARKTz6M1ItvZq90/VT/MJU2xpWvkGQ+dw6gV0
+/ctehYYhrIWDKOc71A/fVTO73+JyWfvwZtA97oY/m0=
`protect END_PROTECTED
