`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m2o7NB9mA/NrrhzX99ObFuVnewTQVmqtpiOjNFj6Dwt9AirKOcJcIporaiQYB1ku
UR1Jp9NpRsuWU19KPr54x4Rs13DoGNSxn5RKPePrxugYmMkwYinRK2l3elEDWUDX
JEdttA9KKT4cvrmmPWiVeovQN29bcJ3U0bijuomHVSzmxquucPn6ZXduTe1FPxNP
mbTYustxVRye6cRIzposZw5R3nI50mbrmKSVuayV59Zc1C/ys3e3NL+dlPUwwvOc
YEharC5NY7zr5YVPLI8KMlIBkISPffOla4oX9HGllRBZnOMSWGxDkHFFjgxHwRzj
U6XyAiLdK6Hrh4L+4yO3KdG+qjdqWHs+Dg0CdF5I43k5rl68nHECW8za4xA3M1/L
0+LiJqWWQQMh2JztzMGjpQ4vThHFnOar4iHssKfXVq5YhXyA/8Q3+RISQc4mrsLJ
4rMDNFqs7RfieN2eXmFwwA01KsBVw0++hkCwkWmJO+XLshwpDazHFy7xuffUBjb8
29ESOmJHEFPL5WHDhBVIdBTSEmWPucy8WVS9qntDwszYrv0ZQtw71tpq8Lkbp0pF
kw3Sp+oELd9mNF9+z57vxGLroRQHjbmrdBx4FwT1AjZ1JelKfNCKn91b7W4X4lkj
uPlg8MjNIowoCchkgWz01bwQU46urVRyqHhGXa1RQxNWCqkhf42AdDp7GGHOFwsu
osimoFrFQbw5BqZL2WALFORe+hAA4QXXq9+rJagfmlSQdrxGhW+1QrymPAGGFOEw
Isi8zH+AwEVWKUjA4OK/3yFFh60TSYjAnlZPQK+/k/gBFewZTQ+BVCivoK7ahu3a
qYYkNTxV1xBgB4/mr3LJV1XbDP7EFUnDVj5pP3Ld5ADXEhGKvZcYCj/es+TPbCHu
jtJHcyGaw7MXkfJ0j926d2d1yuUrYPY3KC8cxtrOishjMEIdtJb6XspO7E0qYxfy
zUgTX5Sq9G8/BldEU0TqiZEee6MUDNoWJsXEB+tXyiLvYcyl4g2cUuEvktas3e+j
F5JYW4y046Fs1xHSPVV2RWdZ6urAsImrMUUHiJCTb5K9EJoGJ1DRLoxXK0p7rKcc
BK6JQVuUMMcHJENL4/eu6g2er/GFYKgh8Su8nTSlhH7zaihgr81vKcKubFfGtvuv
zB63kbvykR2BB7A6i4Kt2/Jv8wM8s/cQhhjrLuLWGHstdUf92EA8JAENBxy3/xj5
bXfe36GfZmiq+21n9LQKqdVXni5TaDbqeTCgBjSTMWDMNCBIIPk76dlwYgQYSyk+
kW7s8lx85f+13b5BIfI/ezWeXfn5zu2XeFKA3AAvTR+N0lRfetthq97FOcu7x7M3
6/P5EV+Rh67YUom3GL+O+4TIVRaPvkjzzq806lkr3/NWWM1SEuq/wyyv+yGs1JsC
NjM9RaZIiNDSfuL7GqvfPQeLP5Qwmz37gOLDHNsOsPIcEm91YUTFpDeUP766quYu
hyNiVsQxuW5nXB2O7Nbw5Q8vKf4wCung8CrovbNrzgDy4o+Y3yOBqhdwNm8rm0Ae
02VHbnL8BXvNzrXtXudC8bOebmUar6JeeeBsi3xiYOmJtf5jB3zuxaX2KKnKFEMP
3KkA+dMms4FpYH/xvmSL9I1LTd83xk+mDPfn+U5NUM8zREj0DTG/J9MDtFAnB8GW
D6LwKBJ0aHfhIchuYMB041IK7vsySe66TGWhm0H59Jk1+Cf/f9bf5+5c6hk2mv1t
Rv4aTaKMXm3n6lCPdkOSCkfZOVBF9GPqZc1m0P6jmmWb5VAScHOPrPQXN0g4urVx
ZG9QG2rlfn/ej7Q+rcKI8NOqRpOiwb2HJenZ/wlfC0V8D/j2kra5S3gZa5X0pcr0
/5WYORAvlGmdT5ldHZb+U1BrA/sSRY/R5gE+aJm3g9vJF8NVHM5bexg6rVkns//B
K3Q/cAMN0Knx95CLV/qT2bjV2Zbt6JMxnQl1KbCiCZQScArMZKmZV9qyBU3/zcW2
8BmSdvS+ZE05tP9Ot9pfh5d8LnpnFacTeceSZH2gT57KmFWLodcvZmuyriXmlVcE
IAa0IoZ172+ttiBpGqixigzRfzBMT1y2oL4ELIuCJlajUNeCrCdbmjFDzkhmRcqB
FSUrPeVr0JMQ35jg1GbyQqkGsyGo+egPSYwDqGby9NrfK9xw9stwq0jvTqLQ9UrH
9WANabbhOucY/Ljaaf+EO0YOTJsCTYWG2qE8wjdIyUoRpQZIHOhr1cehhLSnOT1J
i4IC5svC4jPqzXg5K8qFyli0Y9ezT181C2MiFrRpQA04LhjUYkP3bdzM29Kb5J8L
qJXMomR/EWzF6oUdjUYktX106naJmv39r5kgYnQFI1RWCu70j986xQ0L8AZQ6SCn
jjVCliZCtEXphEh58531vp8V6dYvXNWp0PBEcUJDKVs7zpPD0eCRRwtJDiYnMRJM
Mi36oYke+M1L/4NRAIdNTb8Zq8DGmdmUHhUeP6gma9Z/wFZ/0YIVZ0fcf0glYqWM
aSf+OJ8PZfwsvfs82TupP6fZVpYOVCvXVBZyrqxn9vmuOJM+1zGo8Ty8hxTUTpxp
9Fnqh32GkZbALixhtpCi51TEGbbJe/H7uZ72S0haX6TM/xgBwwNDB4ybbq/HmYD/
k5VYiEpKfpRKm+TieeHoyK5qqpOG4Byo0HVfTa8uVjDkGdGsrda7r+FMYVUqNiby
4/Gld3C0uq0iLef1zYG5OyMLPSH3A/1axIGoBDXjvXG5NGQ+zkbNenbXdOf83HN0
PlXBWn/96tDLpvjcjKgmfKFEXJGmFln8pBlcyt+OB4qC0P8XlPGrvVyn/jO76FNt
voVlIWmHbYgBtw+ls2V2NeZtHwINQfQOt7QVEPo30QSlJwzcwj1Ba6HdHNhlX0WA
llehRMd0O1S0qAroP2eVwo1W6G4sP8lvQ5tV6UqT9Eup4YnR0kfyVZ8b9x87mF7D
DktP3ztaxU8y5TQqhWw81yiSDhfpg5YdEI0yKiZzrc3iNbBcHemFZsZ+WI3uggHv
69R3hNm4sE/zDYtYYapQG861bEaOEDktgGQkHCHwGRpaXgmrquFVbcaOqdlpaRgF
Xej5/JZXVHVpP02IcMBxFdDuUW4sOBecbM74dVssWnoSI3rghgMZZ9OxZmwFhA80
lNBzjblmebP5kxU1v5p81JDoLHRGwLN012oYogw8y4Q5Tt1Tp8mhtwGwoXIDGo9w
OUDT6ojdtSWH0IKOO8KdTU5RMoQvzITefLXj4kZHBWxMv2S657qp0C6wYgPQFssq
xMawu2IRVnC/4pnQ2RCGsUsBgxeNHAAmAfzOvXpZgdDinOBrCun7dSGKkEZFystK
+7k2Ft1Z0BozZckLb8Nam0k/uV23dlJpJuzd3T4g33Z05bQi7Cy4yKNg+mU0zqX6
O+/rPN32CcFg6WH+FzozUKSM9CKWvCGWn938I8IzX6nwzt+bDLE5AI5Tg8OriYYa
jCO+rU4JsNbR87GIvOY0oqI6kMny3cVWC2Q0pJE7ShTCKuGculIyKKsI81s5oJKo
R95kIRFvGYimF2g9meIatZDjbfpeU+k9t7GO4SJpsfybjsybaTHngj+BGGAaHKXs
VhVcRwe0XowbutW3g0ovUYu1s9T1ve0Wi4/KvDRVjWOwLxfDRrUlxUekqWMkTMlS
8Fae0hcUF1kOhZY3KADcESHlhPo+Y6q68lTOhqy4kWujgSkz5d0xOUk9WqoAvR2t
4btBrRjcvSecALomZnUatwhy82k0LnG7HTqglRIJeCO/5ElcYJvH4l37rmFdvOWv
s/Cu6+Ypa5J+Zh4GKw+G0wxHlQSz/pzdTEvUBh4L3K7w2aYjr9fftXLKPvsTE3Jq
iVzBkk/l0Hh+Ya0Y1OP375TLQgx2ZGXRG97cnuE0c+L4vWZ0fGRZIgVPmbgkdw7R
k6mFt9/NnZfrcqOp1fTpR65DbISrtzEv1zbkzul+pAc5G5ysqeFPFX1+rHrssZcD
vtwpRQlYHQKUdPgr9uX4PjNm+OGztX23e26rpR9WotgCG7gBV4w1AqYTYuh/0tdC
3CRfIhMMEJhRJlMtzRzBMHMfWuu29zdtOS0rp+DJMU44JG1G8oOjb0LXWQi+5JvY
g1UhJ48CsBdK5xR82E+QYbJZR0cikqA6fR8yU0FxbmIrSz3tUqD5z6krAOHwqLzZ
d6tcx+PlAU1T1jI1xVmNx5SZVVG4zfnaZEK1B7ivPXcrL+Ax5/ySpTiq95Z0TXoL
uJNQjGbswILYT20d5WPhYc+g4M3GzMARf7+aMBJi7pOsHpwslS98wn4Yvzh+vvhy
eQv6Yjxj+YLU11ZTjHwbylOvyyrFQp/fov/JdMGxvn5kIEeXiZ8CbT9lfAv00wo5
XP0LTUAQcocUFa6HM8T4pGgT7MpL0CMH0yQRU/yTN9Hc9kKJQJnj1S2RzMfF2pze
0EZXJhzL/CAtloyrhcvkeA==
`protect END_PROTECTED
