`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
92L6NNLxhleGtD3S9Q0loQ/zoXx0LMgx4zITTBEPALvXK32stp6PxKhZfo21rorj
pHk3Izb5d2lO+PCSw0Pzob0ZXUP0bFDy3dRI8uvKhunZovS+0rihlsEuldmx+blK
I9228vIv0Bz1SQeJ1qOvEg2PZwq9tfkNthbuO5VctA8qbLrN8ttvnNcn+ENgm9Pk
99iRyn0pksYQf3VpG5rWhkALx+UvNxlo/aW3rUx7VLVYqu4qO1e0+Dc9iS9937Au
d0zUHKiZ/viB9LNAVW8nE7DFctu7gk13n4dqSaI66KzRixB0g4Js1cE0UAU91vTU
pDYoWV3ZPP53G9UIa8S35nFGrW6uuWWLex5B3AJr0eBWrRvZZNWyqahcZ+99v6oz
8cPvxCf6Actz9R+6zVWzSi5ZhHJRl5br+UrtZe+PIxabbjDiP4vTzJDH2v7Jby6v
JIYBCo+5QhU+r0qaLI4TUkFsuQzh+F19vy0SSirH8GtuI7C245F0gJNmJpaZQkO0
IhKqPcSrqO+f5X6wfNq8itUtTlT6UfbalFQ9wAPK2Ju5RHw9QhTJx4kFtJT1RXMv
gW6hsChS6xaA7eIv/auEdBx1ibvg3sEr1VhLKB6j1us7iPl0lfexKCiSjnYdsj83
Ris4aCSMat8oEDapPWbkiEjPAMYy8xJnRQ7qE2w7NIXn1DLLygVrUgWTvCEy0hK5
oE1+x5KHWGLkiLDBbOys5LWIp72mhaTaXl5RLW3DX/MSEp3FXZXe4XgQIkuQohP3
BqkTRdjsfrQ8VoFOwt+u2xtxRTaXE/70SCufQvTGA83dWEMdnENabARuJnd2D0eT
FxLne/V2I0+MMlxYpuQezzFoMUQbK94zMGtW5htN4FNlVl+t5qGxrX2dLLeYLMn4
QMJXIMHMe1kcHQaSoaG6dso5TLCOw8oplyyQp4UymbReG9NrznLmkmOBazrPPvkf
ZzKYk3Y14NaKFOzG6SY4ETeI+fcq6zuX9FT2tNPq1GO9BtQC2amtiQNEWGZW0yIH
2Tun8mjf1mU3YXOZosfvu9L857qrpbFdX4XAD7fFV8erad/KiVmRnCro33ZG4Qt7
p7N7VhupPMI82K8YyvojaysHPeoJ4d0bonMXY81oDKcLNo6fsneP4QNlz9BVJpjE
pKdSXG7tyaVi2PhiYOXxFTvXpamwq96GR/lCBdgKXuvrpg89Rres449PwIQhN+VX
iijIMaPl2VCJZDS2MEWLYXDz4AdM7/QXdzKfURV0jpqSopfnoySQDQihs0xbLtSD
borWZ8XQJGOadXvn/Ddjy17EYQz7ejU/x8HfqIpqLsFSZjga6ptRHT5ZYxKlVEvi
0ybyGWneD7VhlPm9lei/LyifLw8hPOrM7AHiyzCkQDu74j4AGpK4EO4STiP2RrK/
jL77IE5N3vFeBZN9TS3Qlj0aF9ezmbAHV1VwlNniqK0yGMblpSVGJEHvnFg8w0Ov
jsU9BWtCPtPSNWSzG/Uy59TMMuqZeePZ7iAsW8dLI4fcoeNtog4U3CEeZHox/tbv
RyAZvnoDbD13WPEffq6yhrSBvNxv6pXCeBBzJ/kbmhTXIJCSIe156BkggfVn3Dn+
DH/kyQFYmtiqXhgRsVJr23A0iXm12q0ASw3BUeuYhPVuDP+CwuPLrebvs01S+KqZ
SfzZmKNrK7ZRx7NzZ5WPaa9gkSYLnLcWFHnJCrQSWgI=
`protect END_PROTECTED
