`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LsmhJayyKU28rqqk6J2xlC1WmgGA8HnrxrOhzHt6RzyPgFk5bjxpHvfUB+QDvarW
xYcTuGmkAjpBvmbRZ8Sy/f8LHXMV+3caI0vAjH7UiChBEZTd8jnOc4JNWPPaI40w
IFsWwWmxwCgEP01jzo/LZPz0M3c0Rnhocr/MV3NKOHi9RSXLyx1i0RbD2PWyBkwi
lIeS0WdFLB1Jgi4nOmHezqMuN+ult60lh12xqC7G572Uv0MliPwQrxIzVwprOPNu
zu9SOAw+ZjIBUhKdsX4kjEcdbCLmRJPi+WrVvKIAkCdfhOiCkykglSrB3Pds9T8w
pZXAdRc3DJpQMBr6qNwOlT/vYOxwJEftLpZTls5i5hCJgGmPUv3jTRLFXswwipwp
7ogr9h11Qp7cFwRmcUdg2w==
`protect END_PROTECTED
