`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UuAF7s1JuneSSqYiFkfg8DW/WF2wX300mIofNunXMIKCAFGgqq6rK9dRkk0V76Sb
C/wHqLN8wMlniMLaJpEH+2RO6EYgbOCgqEJKjqBW/gyxjD7lLEWildUaJzc5t3Za
CnZPAXRgzR3Fb67RZPjtVkRU5OvLk5KW8WyCixkzBCLlmC6bL0kIHgeI2Fqenn9G
V8JqWMxgytwcQo9Wdut2UwVXYXap38AXSR19wOexRhDfqFzqqXQOV/PJN48tyw45
pinLfuak/6yF7+c7lQy2wFKtXUGSxC5Q4xIb+yu6WXKzN0ZwdI8Z2VXspl5mz8iM
lZuQHwEX2QSN721dpW0JLXjJOIYUYuAWjJFuaCxPJ2tUMKC+OruCAF4Ds7WU/T8A
ZAtz0h7wvih0H7ktjBBNcKMf4AK6V0lsn8Obx55pSRFwYItmjYfO+8gt2LUORn0c
pbqC7ULwRQOoIfc2QRIxe/IQfXTUZT2Fis8lScPpBDv2zoI7K0w8ky7Gh4N0lk1G
5VcSE7DU9oxq7jQDmiwGEtDdnsjmfg6brRlqxnat5C4=
`protect END_PROTECTED
