library verilog;
use verilog.vl_types.all;
entity GTP_HSST is
    generic(
        PCS_CH0_BYPASS_WORD_ALIGN: string  := "FALSE";
        PCS_CH0_BYPASS_DENC: string  := "FALSE";
        PCS_CH0_BYPASS_BONDING: string  := "FALSE";
        PCS_CH0_BYPASS_CTC: string  := "FALSE";
        PCS_CH0_BYPASS_GEAR: string  := "FALSE";
        PCS_CH0_BYPASS_BRIDGE: string  := "FALSE";
        PCS_CH0_DATA_MODE: string  := "X8";
        PCS_CH0_RX_POLARITY_INV: string  := "DELAY";
        PCS_CH0_ALIGN_MODE: string  := "1GB";
        PCS_CH0_SAMP_16B: string  := "X16";
        PCS_CH0_COMMA_REG0: integer := 0;
        PCS_CH0_COMMA_MASK: integer := 0;
        PCS_CH0_CEB_MODE: string  := "10GB";
        PCS_CH0_CTC_MODE: string  := "1SKIP";
        PCS_CH0_A_REG   : integer := 0;
        PCS_CH0_GE_AUTO_EN: string  := "FALSE";
        PCS_CH0_SKIP_REG0: integer := 0;
        PCS_CH0_SKIP_REG1: integer := 0;
        PCS_CH0_SKIP_REG2: integer := 0;
        PCS_CH0_SKIP_REG3: integer := 0;
        PCS_CH0_DEC_DUAL: string  := "FALSE";
        PCS_CH0_SPLIT   : string  := "FALSE";
        PCS_CH0_FIFOFLAG_CTC: string  := "FALSE";
        PCS_CH0_COMMA_DET_MODE: string  := "COMMA_PATTERN";
        PCS_CH0_ERRDETECT_SILENCE: string  := "FALSE";
        PCS_CH0_PMA_RCLK_POLINV: string  := "PMA_RCLK";
        PCS_CH0_PCS_RCLK_SEL: string  := "PMA_RCLK";
        PCS_CH0_MCB_RCLK_POLINV: string  := "MCB_RCLK";
        PCS_CH0_CB_RCLK_SEL: string  := "PMA_RCLK";
        PCS_CH0_AFTER_CTC_RCLK_SEL: string  := "PMA_RCLK";
        PCS_CH0_RCLK_POLINV: string  := "RCLK";
        PCS_CH0_BRIDGE_RCLK_SEL: string  := "PMA_RCLK";
        PCS_CH0_PCS_RCLK_EN: string  := "FALSE";
        PCS_CH0_CB_RCLK_EN: string  := "FALSE";
        PCS_CH0_AFTER_CTC_RCLK_EN: string  := "FALSE";
        PCS_CH0_AFTER_CTC_RCLK_EN_GB: string  := "FALSE";
        PCS_CH0_BRIDGE_RCLK_EN: string  := "FALSE";
        PCS_CH0_PCS_RX_RSTN: string  := "FALSE";
        PCS_CH0_SLAVE   : string  := "MASTER";
        PCS_CH0_PCIE_SLAVE: string  := "MASTER";
        PCS_CH0_PCS_CB_RSTN: string  := "FALSE";
        PCS_CH0_TX_BYPASS_BRIDGE_UINT: string  := "FALSE";
        PCS_CH0_TX_BYPASS_GEAR: string  := "FALSE";
        PCS_CH0_TX_BYPASS_ENC: string  := "FALSE";
        PCS_CH0_TX_BYPASS_BIT_SLIP: string  := "FALSE";
        PCS_CH0_TX_GEAR_SPLIT: string  := "FALSE";
        PCS_CH0_TX_DRIVE_REG_MODE: string  := "NO_CHANGE";
        PCS_CH0_TX_BIT_SLIP_CYCLES: integer := 0;
        PCS_CH0_INT_TX_MASK_0: string  := "FALSE";
        PCS_CH0_INT_TX_MASK_1: string  := "FALSE";
        PCS_CH0_INT_TX_MASK_2: string  := "FALSE";
        PCS_CH0_INT_TX_CLR_0: string  := "FALSE";
        PCS_CH0_INT_TX_CLR_1: string  := "FALSE";
        PCS_CH0_INT_TX_CLR_2: string  := "FALSE";
        PCS_CH0_TX_PMA_TCLK_POLINV: string  := "PMA_TCLK";
        PCS_CH0_TX_PCS_CLK_EN_SEL: string  := "FALSE";
        PCS_CH0_TX_BRIDGE_TCLK_SEL: string  := "PCS_TCLK";
        PCS_CH0_TX_TCLK_POLINV: string  := "TCLK";
        PCS_CH0_TX_PCS_TX_RSTN: string  := "FALSE";
        PCS_CH0_TX_SLAVE: string  := "SLAVE";
        PCS_CH0_TX_BRIDGE_CLK_EN_SEL: string  := "FALSE";
        PCS_CH0_DATA_WIDTH_MODE: string  := "X20";
        PCS_CH0_TX_TCLK2FABRIC_SEL: string  := "FALSE";
        PCS_CH0_TX_OUTZZ: string  := "FALSE";
        PCS_CH0_ENC_DUAL: string  := "FALSE";
        PCS_CH0_TX_BITSLIP_DATA_MODE: string  := "X10";
        PCS_CH0_COMMA_REG1: integer := 0;
        PCS_CH0_RAPID_IMAX: integer := 0;
        PCS_CH0_RAPID_VMIN_1: integer := 0;
        PCS_CH0_RAPID_VMIN_2: integer := 0;
        PCS_CH0_RX_PRBS_MODE: string  := "DISABLE";
        PCS_CH0_RX_ERRCNT_CLR: string  := "FALSE";
        PCS_CH0_TX_PRBS_MODE: string  := "DISABLE";
        PCS_CH0_TX_INSERT_ER: string  := "FALSE";
        PCS_CH0_ENABLE_PRBS_GEN: string  := "FALSE";
        PCS_CH0_ERR_CNT : integer := 0;
        PCS_CH0_DEFAULT_RADDR: integer := 0;
        PCS_CH0_MASTER_CHECK_OFFSET: integer := 0;
        PCS_CH0_DELAY_SET: integer := 0;
        PCS_CH0_SEACH_OFFSET: string  := "20BIT";
        PCS_CH0_CEB_RAPIDLS_MMAX: integer := 0;
        PCS_CH0_CTC_AFULL: integer := 0;
        PCS_CH0_CTC_AEMPTY: integer := 0;
        PCS_CH0_FAR_LOOP: string  := "FALSE";
        PCS_CH0_NEAR_LOOP: string  := "FALSE";
        PCS_CH0_INT_RX_MASK_0: string  := "FALSE";
        PCS_CH0_INT_RX_MASK_1: string  := "FALSE";
        PCS_CH0_INT_RX_MASK_2: string  := "FALSE";
        PCS_CH0_INT_RX_MASK_3: string  := "FALSE";
        PCS_CH0_INT_RX_MASK_4: string  := "FALSE";
        PCS_CH0_INT_RX_MASK_5: string  := "FALSE";
        PCS_CH0_INT_RX_MASK_6: string  := "FALSE";
        PCS_CH0_INT_RX_MASK_7: string  := "FALSE";
        PCS_CH0_INT_RX_CLR_0: string  := "FALSE";
        PCS_CH0_INT_RX_CLR_1: string  := "FALSE";
        PCS_CH0_INT_RX_CLR_2: string  := "FALSE";
        PCS_CH0_INT_RX_CLR_3: string  := "FALSE";
        PCS_CH0_INT_RX_CLR_4: string  := "FALSE";
        PCS_CH0_INT_RX_CLR_5: string  := "FALSE";
        PCS_CH0_INT_RX_CLR_6: string  := "FALSE";
        PCS_CH0_INT_RX_CLR_7: string  := "FALSE";
        PCS_CH1_BYPASS_WORD_ALIGN: string  := "FALSE";
        PCS_CH1_BYPASS_DENC: string  := "FALSE";
        PCS_CH1_BYPASS_BONDING: string  := "FALSE";
        PCS_CH1_BYPASS_CTC: string  := "FALSE";
        PCS_CH1_BYPASS_GEAR: string  := "FALSE";
        PCS_CH1_BYPASS_BRIDGE: string  := "FALSE";
        PCS_CH1_DATA_MODE: string  := "X8";
        PCS_CH1_RX_POLARITY_INV: string  := "DELAY";
        PCS_CH1_ALIGN_MODE: string  := "1GB";
        PCS_CH1_SAMP_16B: string  := "X16";
        PCS_CH1_COMMA_REG0: integer := 0;
        PCS_CH1_COMMA_MASK: integer := 0;
        PCS_CH1_CEB_MODE: string  := "10GB";
        PCS_CH1_CTC_MODE: string  := "1SKIP";
        PCS_CH1_A_REG   : integer := 0;
        PCS_CH1_GE_AUTO_EN: string  := "FALSE";
        PCS_CH1_SKIP_REG0: integer := 0;
        PCS_CH1_SKIP_REG1: integer := 0;
        PCS_CH1_SKIP_REG2: integer := 0;
        PCS_CH1_SKIP_REG3: integer := 0;
        PCS_CH1_DEC_DUAL: string  := "FALSE";
        PCS_CH1_SPLIT   : string  := "FALSE";
        PCS_CH1_FIFOFLAG_CTC: string  := "FALSE";
        PCS_CH1_COMMA_DET_MODE: string  := "COMMA_PATTERN";
        PCS_CH1_ERRDETECT_SILENCE: string  := "FALSE";
        PCS_CH1_PMA_RCLK_POLINV: string  := "PMA_RCLK";
        PCS_CH1_PCS_RCLK_SEL: string  := "PMA_RCLK";
        PCS_CH1_MCB_RCLK_POLINV: string  := "MCB_RCLK";
        PCS_CH1_CB_RCLK_SEL: string  := "PMA_RCLK";
        PCS_CH1_AFTER_CTC_RCLK_SEL: string  := "PMA_RCLK";
        PCS_CH1_RCLK_POLINV: string  := "RCLK";
        PCS_CH1_BRIDGE_RCLK_SEL: string  := "PMA_RCLK";
        PCS_CH1_PCS_RCLK_EN: string  := "FALSE";
        PCS_CH1_CB_RCLK_EN: string  := "FALSE";
        PCS_CH1_AFTER_CTC_RCLK_EN: string  := "FALSE";
        PCS_CH1_AFTER_CTC_RCLK_EN_GB: string  := "FALSE";
        PCS_CH1_BRIDGE_RCLK_EN: string  := "FALSE";
        PCS_CH1_PCS_RX_RSTN: string  := "FALSE";
        PCS_CH1_SLAVE   : string  := "MASTER";
        PCS_CH1_PCIE_SLAVE: string  := "MASTER";
        PCS_CH1_PCS_CB_RSTN: string  := "FALSE";
        PCS_CH1_TX_BYPASS_BRIDGE_UINT: string  := "FALSE";
        PCS_CH1_TX_BYPASS_GEAR: string  := "FALSE";
        PCS_CH1_TX_BYPASS_ENC: string  := "FALSE";
        PCS_CH1_TX_BYPASS_BIT_SLIP: string  := "FALSE";
        PCS_CH1_TX_GEAR_SPLIT: string  := "FALSE";
        PCS_CH1_TX_DRIVE_REG_MODE: string  := "NO_CHANGE";
        PCS_CH1_TX_BIT_SLIP_CYCLES: integer := 0;
        PCS_CH1_INT_TX_MASK_0: string  := "FALSE";
        PCS_CH1_INT_TX_MASK_1: string  := "FALSE";
        PCS_CH1_INT_TX_MASK_2: string  := "FALSE";
        PCS_CH1_INT_TX_CLR_0: string  := "FALSE";
        PCS_CH1_INT_TX_CLR_1: string  := "FALSE";
        PCS_CH1_INT_TX_CLR_2: string  := "FALSE";
        PCS_CH1_TX_PMA_TCLK_POLINV: string  := "PMA_TCLK";
        PCS_CH1_TX_PCS_CLK_EN_SEL: string  := "FALSE";
        PCS_CH1_TX_BRIDGE_TCLK_SEL: string  := "PCS_TCLK";
        PCS_CH1_TX_TCLK_POLINV: string  := "TCLK";
        PCS_CH1_TX_PCS_TX_RSTN: string  := "FALSE";
        PCS_CH1_TX_SLAVE: string  := "SLAVE";
        PCS_CH1_TX_BRIDGE_CLK_EN_SEL: string  := "FALSE";
        PCS_CH1_DATA_WIDTH_MODE: string  := "X20";
        PCS_CH1_TX_TCLK2FABRIC_SEL: string  := "FALSE";
        PCS_CH1_TX_OUTZZ: string  := "FALSE";
        PCS_CH1_ENC_DUAL: string  := "FALSE";
        PCS_CH1_TX_BITSLIP_DATA_MODE: string  := "X10";
        PCS_CH1_COMMA_REG1: integer := 0;
        PCS_CH1_RAPID_IMAX: integer := 0;
        PCS_CH1_RAPID_VMIN_1: integer := 0;
        PCS_CH1_RAPID_VMIN_2: integer := 0;
        PCS_CH1_RX_PRBS_MODE: string  := "DISABLE";
        PCS_CH1_RX_ERRCNT_CLR: string  := "FALSE";
        PCS_CH1_TX_PRBS_MODE: string  := "DISABLE";
        PCS_CH1_TX_INSERT_ER: string  := "FALSE";
        PCS_CH1_ENABLE_PRBS_GEN: string  := "FALSE";
        PCS_CH1_ERR_CNT : integer := 0;
        PCS_CH1_DEFAULT_RADDR: integer := 0;
        PCS_CH1_MASTER_CHECK_OFFSET: integer := 0;
        PCS_CH1_DELAY_SET: integer := 0;
        PCS_CH1_SEACH_OFFSET: string  := "20BIT";
        PCS_CH1_CEB_RAPIDLS_MMAX: integer := 0;
        PCS_CH1_CTC_AFULL: integer := 0;
        PCS_CH1_CTC_AEMPTY: integer := 0;
        PCS_CH1_FAR_LOOP: string  := "FALSE";
        PCS_CH1_NEAR_LOOP: string  := "FALSE";
        PCS_CH1_INT_RX_MASK_0: string  := "FALSE";
        PCS_CH1_INT_RX_MASK_1: string  := "FALSE";
        PCS_CH1_INT_RX_MASK_2: string  := "FALSE";
        PCS_CH1_INT_RX_MASK_3: string  := "FALSE";
        PCS_CH1_INT_RX_MASK_4: string  := "FALSE";
        PCS_CH1_INT_RX_MASK_5: string  := "FALSE";
        PCS_CH1_INT_RX_MASK_6: string  := "FALSE";
        PCS_CH1_INT_RX_MASK_7: string  := "FALSE";
        PCS_CH1_INT_RX_CLR_0: string  := "FALSE";
        PCS_CH1_INT_RX_CLR_1: string  := "FALSE";
        PCS_CH1_INT_RX_CLR_2: string  := "FALSE";
        PCS_CH1_INT_RX_CLR_3: string  := "FALSE";
        PCS_CH1_INT_RX_CLR_4: string  := "FALSE";
        PCS_CH1_INT_RX_CLR_5: string  := "FALSE";
        PCS_CH1_INT_RX_CLR_6: string  := "FALSE";
        PCS_CH1_INT_RX_CLR_7: string  := "FALSE";
        PCS_CH2_BYPASS_WORD_ALIGN: string  := "FALSE";
        PCS_CH2_BYPASS_DENC: string  := "FALSE";
        PCS_CH2_BYPASS_BONDING: string  := "FALSE";
        PCS_CH2_BYPASS_CTC: string  := "FALSE";
        PCS_CH2_BYPASS_GEAR: string  := "FALSE";
        PCS_CH2_BYPASS_BRIDGE: string  := "FALSE";
        PCS_CH2_DATA_MODE: string  := "X8";
        PCS_CH2_RX_POLARITY_INV: string  := "DELAY";
        PCS_CH2_ALIGN_MODE: string  := "1GB";
        PCS_CH2_SAMP_16B: string  := "X16";
        PCS_CH2_COMMA_REG0: integer := 0;
        PCS_CH2_COMMA_MASK: integer := 0;
        PCS_CH2_CEB_MODE: string  := "10GB";
        PCS_CH2_CTC_MODE: string  := "1SKIP";
        PCS_CH2_A_REG   : integer := 0;
        PCS_CH2_GE_AUTO_EN: string  := "FALSE";
        PCS_CH2_SKIP_REG0: integer := 0;
        PCS_CH2_SKIP_REG1: integer := 0;
        PCS_CH2_SKIP_REG2: integer := 0;
        PCS_CH2_SKIP_REG3: integer := 0;
        PCS_CH2_DEC_DUAL: string  := "FALSE";
        PCS_CH2_SPLIT   : string  := "FALSE";
        PCS_CH2_FIFOFLAG_CTC: string  := "FALSE";
        PCS_CH2_COMMA_DET_MODE: string  := "COMMA_PATTERN";
        PCS_CH2_ERRDETECT_SILENCE: string  := "FALSE";
        PCS_CH2_PMA_RCLK_POLINV: string  := "PMA_RCLK";
        PCS_CH2_PCS_RCLK_SEL: string  := "PMA_RCLK";
        PCS_CH2_MCB_RCLK_POLINV: string  := "MCB_RCLK";
        PCS_CH2_CB_RCLK_SEL: string  := "PMA_RCLK";
        PCS_CH2_AFTER_CTC_RCLK_SEL: string  := "PMA_RCLK";
        PCS_CH2_RCLK_POLINV: string  := "RCLK";
        PCS_CH2_BRIDGE_RCLK_SEL: string  := "PMA_RCLK";
        PCS_CH2_PCS_RCLK_EN: string  := "FALSE";
        PCS_CH2_CB_RCLK_EN: string  := "FALSE";
        PCS_CH2_AFTER_CTC_RCLK_EN: string  := "FALSE";
        PCS_CH2_AFTER_CTC_RCLK_EN_GB: string  := "FALSE";
        PCS_CH2_BRIDGE_RCLK_EN: string  := "FALSE";
        PCS_CH2_PCS_RX_RSTN: string  := "FALSE";
        PCS_CH2_SLAVE   : string  := "MASTER";
        PCS_CH2_PCIE_SLAVE: string  := "MASTER";
        PCS_CH2_PCS_CB_RSTN: string  := "FALSE";
        PCS_CH2_TX_BYPASS_BRIDGE_UINT: string  := "FALSE";
        PCS_CH2_TX_BYPASS_GEAR: string  := "FALSE";
        PCS_CH2_TX_BYPASS_ENC: string  := "FALSE";
        PCS_CH2_TX_BYPASS_BIT_SLIP: string  := "FALSE";
        PCS_CH2_TX_GEAR_SPLIT: string  := "FALSE";
        PCS_CH2_TX_DRIVE_REG_MODE: string  := "NO_CHANGE";
        PCS_CH2_TX_BIT_SLIP_CYCLES: integer := 0;
        PCS_CH2_INT_TX_MASK_0: string  := "FALSE";
        PCS_CH2_INT_TX_MASK_1: string  := "FALSE";
        PCS_CH2_INT_TX_MASK_2: string  := "FALSE";
        PCS_CH2_INT_TX_CLR_0: string  := "FALSE";
        PCS_CH2_INT_TX_CLR_1: string  := "FALSE";
        PCS_CH2_INT_TX_CLR_2: string  := "FALSE";
        PCS_CH2_TX_PMA_TCLK_POLINV: string  := "PMA_TCLK";
        PCS_CH2_TX_PCS_CLK_EN_SEL: string  := "FALSE";
        PCS_CH2_TX_BRIDGE_TCLK_SEL: string  := "PCS_TCLK";
        PCS_CH2_TX_TCLK_POLINV: string  := "TCLK";
        PCS_CH2_TX_PCS_TX_RSTN: string  := "FALSE";
        PCS_CH2_TX_SLAVE: string  := "SLAVE";
        PCS_CH2_TX_BRIDGE_CLK_EN_SEL: string  := "FALSE";
        PCS_CH2_DATA_WIDTH_MODE: string  := "X20";
        PCS_CH2_TX_TCLK2FABRIC_SEL: string  := "FALSE";
        PCS_CH2_TX_OUTZZ: string  := "FALSE";
        PCS_CH2_ENC_DUAL: string  := "FALSE";
        PCS_CH2_TX_BITSLIP_DATA_MODE: string  := "X10";
        PCS_CH2_COMMA_REG1: integer := 0;
        PCS_CH2_RAPID_IMAX: integer := 0;
        PCS_CH2_RAPID_VMIN_1: integer := 0;
        PCS_CH2_RAPID_VMIN_2: integer := 0;
        PCS_CH2_RX_PRBS_MODE: string  := "DISABLE";
        PCS_CH2_RX_ERRCNT_CLR: string  := "FALSE";
        PCS_CH2_TX_PRBS_MODE: string  := "DISABLE";
        PCS_CH2_TX_INSERT_ER: string  := "FALSE";
        PCS_CH2_ENABLE_PRBS_GEN: string  := "FALSE";
        PCS_CH2_ERR_CNT : integer := 0;
        PCS_CH2_DEFAULT_RADDR: integer := 0;
        PCS_CH2_MASTER_CHECK_OFFSET: integer := 0;
        PCS_CH2_DELAY_SET: integer := 0;
        PCS_CH2_SEACH_OFFSET: string  := "20BIT";
        PCS_CH2_CEB_RAPIDLS_MMAX: integer := 0;
        PCS_CH2_CTC_AFULL: integer := 0;
        PCS_CH2_CTC_AEMPTY: integer := 0;
        PCS_CH2_FAR_LOOP: string  := "FALSE";
        PCS_CH2_NEAR_LOOP: string  := "FALSE";
        PCS_CH2_INT_RX_MASK_0: string  := "FALSE";
        PCS_CH2_INT_RX_MASK_1: string  := "FALSE";
        PCS_CH2_INT_RX_MASK_2: string  := "FALSE";
        PCS_CH2_INT_RX_MASK_3: string  := "FALSE";
        PCS_CH2_INT_RX_MASK_4: string  := "FALSE";
        PCS_CH2_INT_RX_MASK_5: string  := "FALSE";
        PCS_CH2_INT_RX_MASK_6: string  := "FALSE";
        PCS_CH2_INT_RX_MASK_7: string  := "FALSE";
        PCS_CH2_INT_RX_CLR_0: string  := "FALSE";
        PCS_CH2_INT_RX_CLR_1: string  := "FALSE";
        PCS_CH2_INT_RX_CLR_2: string  := "FALSE";
        PCS_CH2_INT_RX_CLR_3: string  := "FALSE";
        PCS_CH2_INT_RX_CLR_4: string  := "FALSE";
        PCS_CH2_INT_RX_CLR_5: string  := "FALSE";
        PCS_CH2_INT_RX_CLR_6: string  := "FALSE";
        PCS_CH2_INT_RX_CLR_7: string  := "FALSE";
        PCS_CH3_BYPASS_WORD_ALIGN: string  := "FALSE";
        PCS_CH3_BYPASS_DENC: string  := "FALSE";
        PCS_CH3_BYPASS_BONDING: string  := "FALSE";
        PCS_CH3_BYPASS_CTC: string  := "FALSE";
        PCS_CH3_BYPASS_GEAR: string  := "FALSE";
        PCS_CH3_BYPASS_BRIDGE: string  := "FALSE";
        PCS_CH3_DATA_MODE: string  := "X8";
        PCS_CH3_RX_POLARITY_INV: string  := "DELAY";
        PCS_CH3_ALIGN_MODE: string  := "1GB";
        PCS_CH3_SAMP_16B: string  := "X16";
        PCS_CH3_COMMA_REG0: integer := 0;
        PCS_CH3_COMMA_MASK: integer := 0;
        PCS_CH3_CEB_MODE: string  := "10GB";
        PCS_CH3_CTC_MODE: string  := "1SKIP";
        PCS_CH3_A_REG   : integer := 0;
        PCS_CH3_GE_AUTO_EN: string  := "FALSE";
        PCS_CH3_SKIP_REG0: integer := 0;
        PCS_CH3_SKIP_REG1: integer := 0;
        PCS_CH3_SKIP_REG2: integer := 0;
        PCS_CH3_SKIP_REG3: integer := 0;
        PCS_CH3_DEC_DUAL: string  := "FALSE";
        PCS_CH3_SPLIT   : string  := "FALSE";
        PCS_CH3_FIFOFLAG_CTC: string  := "FALSE";
        PCS_CH3_COMMA_DET_MODE: string  := "COMMA_PATTERN";
        PCS_CH3_ERRDETECT_SILENCE: string  := "FALSE";
        PCS_CH3_PMA_RCLK_POLINV: string  := "PMA_RCLK";
        PCS_CH3_PCS_RCLK_SEL: string  := "PMA_RCLK";
        PCS_CH3_MCB_RCLK_POLINV: string  := "MCB_RCLK";
        PCS_CH3_CB_RCLK_SEL: string  := "PMA_RCLK";
        PCS_CH3_AFTER_CTC_RCLK_SEL: string  := "PMA_RCLK";
        PCS_CH3_RCLK_POLINV: string  := "RCLK";
        PCS_CH3_BRIDGE_RCLK_SEL: string  := "PMA_RCLK";
        PCS_CH3_PCS_RCLK_EN: string  := "FALSE";
        PCS_CH3_CB_RCLK_EN: string  := "FALSE";
        PCS_CH3_AFTER_CTC_RCLK_EN: string  := "FALSE";
        PCS_CH3_AFTER_CTC_RCLK_EN_GB: string  := "FALSE";
        PCS_CH3_BRIDGE_RCLK_EN: string  := "FALSE";
        PCS_CH3_PCS_RX_RSTN: string  := "FALSE";
        PCS_CH3_SLAVE   : string  := "MASTER";
        PCS_CH3_PCIE_SLAVE: string  := "MASTER";
        PCS_CH3_PCS_CB_RSTN: string  := "FALSE";
        PCS_CH3_TX_BYPASS_BRIDGE_UINT: string  := "FALSE";
        PCS_CH3_TX_BYPASS_GEAR: string  := "FALSE";
        PCS_CH3_TX_BYPASS_ENC: string  := "FALSE";
        PCS_CH3_TX_BYPASS_BIT_SLIP: string  := "FALSE";
        PCS_CH3_TX_GEAR_SPLIT: string  := "FALSE";
        PCS_CH3_TX_DRIVE_REG_MODE: string  := "NO_CHANGE";
        PCS_CH3_TX_BIT_SLIP_CYCLES: integer := 0;
        PCS_CH3_INT_TX_MASK_0: string  := "FALSE";
        PCS_CH3_INT_TX_MASK_1: string  := "FALSE";
        PCS_CH3_INT_TX_MASK_2: string  := "FALSE";
        PCS_CH3_INT_TX_CLR_0: string  := "FALSE";
        PCS_CH3_INT_TX_CLR_1: string  := "FALSE";
        PCS_CH3_INT_TX_CLR_2: string  := "FALSE";
        PCS_CH3_TX_PMA_TCLK_POLINV: string  := "PMA_TCLK";
        PCS_CH3_TX_PCS_CLK_EN_SEL: string  := "FALSE";
        PCS_CH3_TX_BRIDGE_TCLK_SEL: string  := "PCS_TCLK";
        PCS_CH3_TX_TCLK_POLINV: string  := "TCLK";
        PCS_CH3_TX_PCS_TX_RSTN: string  := "FALSE";
        PCS_CH3_TX_SLAVE: string  := "SLAVE";
        PCS_CH3_TX_BRIDGE_CLK_EN_SEL: string  := "FALSE";
        PCS_CH3_DATA_WIDTH_MODE: string  := "X20";
        PCS_CH3_TX_TCLK2FABRIC_SEL: string  := "FALSE";
        PCS_CH3_TX_OUTZZ: string  := "FALSE";
        PCS_CH3_ENC_DUAL: string  := "FALSE";
        PCS_CH3_TX_BITSLIP_DATA_MODE: string  := "X10";
        PCS_CH3_COMMA_REG1: integer := 0;
        PCS_CH3_RAPID_IMAX: integer := 0;
        PCS_CH3_RAPID_VMIN_1: integer := 0;
        PCS_CH3_RAPID_VMIN_2: integer := 0;
        PCS_CH3_RX_PRBS_MODE: string  := "DISABLE";
        PCS_CH3_RX_ERRCNT_CLR: string  := "FALSE";
        PCS_CH3_TX_PRBS_MODE: string  := "DISABLE";
        PCS_CH3_TX_INSERT_ER: string  := "FALSE";
        PCS_CH3_ENABLE_PRBS_GEN: string  := "FALSE";
        PCS_CH3_ERR_CNT : integer := 0;
        PCS_CH3_DEFAULT_RADDR: integer := 0;
        PCS_CH3_MASTER_CHECK_OFFSET: integer := 0;
        PCS_CH3_DELAY_SET: integer := 0;
        PCS_CH3_SEACH_OFFSET: string  := "20BIT";
        PCS_CH3_CEB_RAPIDLS_MMAX: integer := 0;
        PCS_CH3_CTC_AFULL: integer := 0;
        PCS_CH3_CTC_AEMPTY: integer := 0;
        PCS_CH3_FAR_LOOP: string  := "FALSE";
        PCS_CH3_NEAR_LOOP: string  := "FALSE";
        PCS_CH3_INT_RX_MASK_0: string  := "FALSE";
        PCS_CH3_INT_RX_MASK_1: string  := "FALSE";
        PCS_CH3_INT_RX_MASK_2: string  := "FALSE";
        PCS_CH3_INT_RX_MASK_3: string  := "FALSE";
        PCS_CH3_INT_RX_MASK_4: string  := "FALSE";
        PCS_CH3_INT_RX_MASK_5: string  := "FALSE";
        PCS_CH3_INT_RX_MASK_6: string  := "FALSE";
        PCS_CH3_INT_RX_MASK_7: string  := "FALSE";
        PCS_CH3_INT_RX_CLR_0: string  := "FALSE";
        PCS_CH3_INT_RX_CLR_1: string  := "FALSE";
        PCS_CH3_INT_RX_CLR_2: string  := "FALSE";
        PCS_CH3_INT_RX_CLR_3: string  := "FALSE";
        PCS_CH3_INT_RX_CLR_4: string  := "FALSE";
        PCS_CH3_INT_RX_CLR_5: string  := "FALSE";
        PCS_CH3_INT_RX_CLR_6: string  := "FALSE";
        PCS_CH3_INT_RX_CLR_7: string  := "FALSE";
        PMA_CH0_TXDATA_WIDTH: string  := "8_BIT";
        PMA_CH0_TX_TESTPATTERN: integer := 0;
        PMA_CH0_TESTPATTERN_O_ENABLE: string  := "FALSE";
        PMA_CH0_DISABLE_BSMODE_DRVAMP: string  := "FALSE";
        PMA_CH0_FORCE_BIST_ENABLE: string  := "FALSE";
        PMA_CH0_FORCE_ELECTRICAL_IDLE: string  := "FALSE";
        PMA_CH0_FORCE_RXDCT_ENABLE: string  := "FALSE";
        PMA_CH0_FORCE_EXTLB_ENABLE: string  := "FALSE";
        PMA_CH0_DISABLE_LANE_SYNC: string  := "FALSE";
        PMA_CH0_DISABLE_ELECTRICAL_IDLE: string  := "FALSE";
        PMA_CH0_DISABLE_RXDCT_ENABLE: string  := "FALSE";
        PMA_CH0_DISABLE_EXTLB_ENABLE: string  := "FALSE";
        PMA_CH0_DISABLE_LOW_SPEED_PATH_ENABLE: string  := "FALSE";
        PMA_CH0_FORCE_LANE_ENABLE: string  := "FALSE";
        PMA_CH0_FORCE_LANE_RESETB_DISABLE: string  := "FALSE";
        PMA_CH0_RXDCT_LGBW_ENABLE: string  := "FALSE";
        PMA_CH0_RXDCT_VTH: string  := "MINUS_300MV";
        PMA_CH0_DE_EMPHASIS_ADDITIONAL_CONTROL: string  := "0DB";
        PMA_CH0_DRV_RTERM_CONTROL: string  := "100PCT";
        PMA_CH0_FDRV_AMP_CONTROL: string  := "100PCT";
        PMA_CH0_PREPC_AMP_CONTROL: string  := "100PCT";
        PMA_CH0_PREMC_AMP_CONTROL: string  := "100PCT";
        PMA_CH0_SER_AMP_CONTROL: string  := "100PCT";
        PMA_CH0_PFD_LOOP_RESISTOR_SETTING: integer := 0;
        PMA_CH0_PD_LOOP_RESISTOR_SETTING: integer := 0;
        PMA_CH0_CDR_TEST_OUT_SELECT: string  := "FBCK";
        PMA_CH0_PI_DIV1_BP: string  := "DISABLE";
        PMA_CH0_PI_TEST_FOR_CKI: string  := "FALSE";
        PMA_CH0_PI_CURRENT_SETTING: string  := "100PCT";
        PMA_CH0_PI_FREQUENCY_SETTING: integer := 0;
        PMA_CH0_TEST_OUT_SELECT_FOR_RCK: string  := "FALSE";
        PMA_CH0_TEST_OUT_SELECT_SOURCE: string  := "SLPI1UI";
        PMA_CH0_TEST_DATA_OUT_SELECT_SOURCE: string  := "DO";
        PMA_CH0_TEST_CK_OUT_SELECT_SOURCE: string  := "DATA";
        PMA_CH0_ENABLE_SLIP1UI_MODULE: string  := "DISABLE";
        PMA_CH0_PN_SWAP_ENABLE: string  := "DISABLE";
        PMA_CH0_SIPO_BIT_SETTING: string  := "10_BIT";
        PMA_CH0_OOB_EN  : string  := "DISABLE";
        PMA_CH0_ALOS_EN : string  := "DISABLE";
        PMA_CH0_LFMODE  : string  := "HIGH";
        PMA_CH0_TSO_HS_SEL: string  := "CDR";
        PMA_CH0_LX_SELLC: string  := "RING";
        PMA_CH0_LX_RXPLL_DIVSEL45_FB: integer := 4;
        PMA_CH0_LX_RXPLL_DIVSEL_FB: integer := 2;
        PMA_CH0_LX_RXPLL_DIVSEL_REF: integer := 1;
        PMA_CH0_PICODE  : integer := 0;
        PMA_CH0_RX_REFCK_SEL: integer := 0;
        PMA_CH0_PFDLPEN_REGISTER_CONTROL_ENABLE: string  := "DISABLE";
        PMA_CH0_PFDLPEN_REGISTER_SETTING: string  := "FALSE";
        PMA_CH0_PDLPEN_REGISTER_CONTROL_ENABLE: string  := "DISABLE";
        PMA_CH0_PDLPEN_REGISTER_SETTING: string  := "FALSE";
        PMA_CH0_DIV_CHANGE_ENABLE_DELAY_TIMER: integer := 0;
        PMA_CH0_DIV_CHANGE_ENABLE_SIGNAL_GATING: string  := "FALSE";
        PMA_CH0_CDR_ALIGN_REGISTER_SETTING_VALUE: string  := "FALSE";
        PMA_CH0_FORCE_CDR_ALIGN_ENABLE: string  := "DISABLE";
        PMA_CH0_SELLC_REGISTER_SETTING_VALUE: string  := "FALSE";
        PMA_CH0_SELLC_CONTROL_BY_REGISTER: string  := "FALSE";
        PMA_CH0_REG_PLLI_LDO_VREF_SETTING: string  := "0_9V";
        PMA_CH0_REG_PLLI_LDO_BYPASS_CURRENT: integer := 0;
        PMA_CH0_REG_PLL_HSTEST_ENABLE: string  := "DISABLE";
        PMA_CH0_REG_PLL_ISNK_CURRENT_CONTROL: string  := "5U";
        PMA_CH0_REG_PLL_PFD_LOOP_CP0_CURRENT_SETTING: integer := 0;
        PMA_CH0_REG_PLL_PD_LOOP_PLLGM_SETTING: string  := "100PCT";
        PMA_CH0_REG_PLL_PFD_LOOP_CP1_CURRENT_SETTING: integer := 0;
        PMA_CH0_REG_PLL_CP0_BIAS_CONTROL: string  := "100PCT";
        PMA_CH0_REG_PLL_PD_LOOP_CP0_CURRENT_SETTING: integer := 0;
        PMA_CH0_REG_PLL_CP1_BIAS_CONTROL: string  := "100PCT";
        PMA_CH0_REG_PLL_PD_LOOP_CP1_CURRENT_SETTING: integer := 0;
        PMA_CH0_REG_PLL_CP0_CURRENT_SETTING: string  := "100PCT";
        PMA_CH0_REG_PLL_CP1_CURRENT_SETTING: string  := "100PCT";
        PMA_CH0_REG_PLL_GM1_CURRENT_SETTING: string  := "100PCT";
        PMA_CH0_REG_PLL_LC_BF2_CURRENT_SETTING: string  := "100PCT";
        PMA_CH0_REG_PLL_LC_BF2_CURRENT_SETTING_LOW: string  := "100PCT";
        PMA_CH0_REG_PLL_REG_CUR: string  := "100PCT";
        PMA_CH0_REG_PLL_LCCUR: string  := "DEFAULT";
        PMA_CH0_REG_PLL_LCOBAS: string  := "100PCT";
        PMA_CH0_REG_PLL_FB_CK_TEST_OUT_ENABLE: string  := "DISABLE";
        PMA_CH0_CDR_ALIGN_TIMER: integer := 0;
        PMA_CH0_CALIB_WAIT: integer := 1024;
        PMA_CH0_CALIB_TIMER: integer := 512;
        PMA_CH0_TOT_RANGE: integer := 0;
        PMA_CH0_SUB_RANGE: integer := 0;
        PMA_CH0_OVLP    : integer := 0;
        PMA_CH0_BIST_WAIT: integer := 1024;
        PMA_CH0_BIST_TIMER: integer := 512;
        PMA_CH0_BAND_LB : integer := 0;
        PMA_CH0_BAND_HB : integer := 0;
        PMA_CH0_FREQ_LOCK_ACCURACY: integer := 0;
        PMA_CH0_REG_SET_LC_BAND: integer := 0;
        PMA_CH0_REG_SET_VCODIV: integer := 0;
        PMA_CH0_REGISTER_SET_VCODIV_BAND_ENABLE: string  := "DISABLE";
        PMA_CH0_REG_SET_PLL_LOCK: string  := "FALSE";
        PMA_CH0_REGISTER_SET_PLL_LOCK_ENABLE: string  := "DISABLE";
        PMA_CH0_REG_SET_VCO_HI: string  := "FALSE";
        PMA_CH0_REG_SET_VCO_LO: string  := "FALSE";
        PMA_CH0_REGISTER_SET_VCO_HI_VCO_LO_ENABLE: string  := "DISABLE";
        PMA_CH0_FORCE_LC_PLL_LOOP_EN_H: string  := "DISABLE";
        PMA_CH0_FORCE_LC_PLL_LOOP_EN_L: string  := "DISABLE";
        PMA_CH0_VCO_DIV_CALI_BYPASS: string  := "FALSE";
        PMA_CH0_BIST_EN : string  := "DISABLE";
        PMA_CH0_PLL_LOOP_EN_SETTING_FROM_REGISTER_ENABLE: string  := "DISABLE";
        PMA_CH0_FREQ_DETECT_ENABLE_SOURCE: string  := "DISABLE";
        PMA_CH0_REG_SET_DIVSEL_REF: integer := 0;
        PMA_CH0_REG_SET_DIVSEL45_FB: string  := "FALSE";
        PMA_CH0_REG_SET_DIVSEL_FB: integer := 0;
        PMA_CH0_PLL_LOOP_EN_SETTING: string  := "DISABLE";
        PMA_CH0_REGISTER_SET_TXPLL_DIV_ENABLE: string  := "DISABLE";
        PMA_CH0_FORCE_RXPLL_RESET: string  := "FALSE";
        PMA_CH0_FORCE_RXPLL_ON: string  := "FALSE";
        PMA_CH0_DPCK_DIV2: string  := "FALSE";
        PMA_CH0_LFO_SETTING: integer := 0;
        PMA_CH0_ALOS_COUNTER_CLOCK_SELECTION: string  := "LOCAL";
        PMA_CH0_RX_BIAS_CURRENT_ADJUSTMENT: string  := "100PCT";
        PMA_CH0_OOB_ENTER_DELAY_SETTING: integer := 0;
        PMA_CH0_ALOS_LOW_TO_HIGH_COUNTER_SETTING: integer := 0;
        PMA_CH0_ENABLE_ALOS_RESULT_AUTOMATICALLY_ENABLE_CHANNEL: string  := "DISABLE";
        PMA_CH0_ALOS_EXIT_COUNTER_CLOCK_DIVIDER: integer := 0;
        PMA_CH0_OOB_OSCILATER_FREQUENCY_SETTING: integer := 0;
        PMA_CH0_FORCE_OOB: string  := "FALSE";
        PMA_CH0_OOB_VTH_SET: string  := "27MV";
        PMA_CH0_FORCE_DET_FORCE_ALOS_LOW: string  := "FALSE";
        PMA_CH0_ALOS_THRESHOLD_VOLTAGE: string  := "27MV";
        PMA_CH0_WAKEUP_VCM_RX_COMMON_MODE_VOLTAGE: integer := 0;
        PMA_CH0_REGR_NEGATIVE_HYSTERESIS_SETTING: string  := "100MV";
        PMA_CH0_REGL_POSITIVE_HYSTERESIS_SETTING: string  := "100MV";
        PMA_CH0_REG_EN  : string  := "DISABLE";
        PMA_CH0_REGREF_SEL: string  := "VREF";
        PMA_CH0_DC496   : string  := "39_6MHZ";
        PMA_CH0_EQ2_AC_VAR_SETTING: integer := 0;
        PMA_CH0_EQ2_AC_RES_SETTING: integer := 0;
        PMA_CH0_EQ2_DC_RESTOP_SETTING: integer := 0;
        PMA_CH0_EQ1_DC_RESTOP_SETTING: integer := 50;
        PMA_CH0_EQ1_AC_VAR_SETTING: integer := 0;
        PMA_CH0_EQ2_CURRENT_SETTING: integer := 0;
        PMA_CH0_EQ1_AC_RES_SETTING: integer := 0;
        PMA_CH0_EQ1_CURRENT_SETTING: integer := 0;
        PMA_CH0_RPLUS   : integer := 0;
        PMA_CH0_RMINUS  : integer := 0;
        PMA_CH0_RVALSET : integer := 0;
        PMA_CH0_RTERM   : integer := 0;
        PMA_CH0_DCFB_EN : string  := "DISABLE";
        PMA_CH0_DCCOUP  : string  := "FALSE";
        PMA_CH0_3G      : string  := "FALSE";
        PMA_CH1_TXDATA_WIDTH: string  := "8_BIT";
        PMA_CH1_TX_TESTPATTERN: integer := 0;
        PMA_CH1_TESTPATTERN_O_ENABLE: string  := "FALSE";
        PMA_CH1_DISABLE_BSMODE_DRVAMP: string  := "FALSE";
        PMA_CH1_FORCE_BIST_ENABLE: string  := "FALSE";
        PMA_CH1_FORCE_ELECTRICAL_IDLE: string  := "FALSE";
        PMA_CH1_FORCE_RXDCT_ENABLE: string  := "FALSE";
        PMA_CH1_FORCE_EXTLB_ENABLE: string  := "FALSE";
        PMA_CH1_DISABLE_LANE_SYNC: string  := "FALSE";
        PMA_CH1_DISABLE_ELECTRICAL_IDLE: string  := "FALSE";
        PMA_CH1_DISABLE_RXDCT_ENABLE: string  := "FALSE";
        PMA_CH1_DISABLE_EXTLB_ENABLE: string  := "FALSE";
        PMA_CH1_DISABLE_LOW_SPEED_PATH_ENABLE: string  := "FALSE";
        PMA_CH1_FORCE_LANE_ENABLE: string  := "FALSE";
        PMA_CH1_FORCE_LANE_RESETB_DISABLE: string  := "FALSE";
        PMA_CH1_RXDCT_LGBW_ENABLE: string  := "FALSE";
        PMA_CH1_RXDCT_VTH: string  := "MINUS_300MV";
        PMA_CH1_DE_EMPHASIS_ADDITIONAL_CONTROL: string  := "0DB";
        PMA_CH1_DRV_RTERM_CONTROL: string  := "100PCT";
        PMA_CH1_FDRV_AMP_CONTROL: string  := "100PCT";
        PMA_CH1_PREPC_AMP_CONTROL: string  := "100PCT";
        PMA_CH1_PREMC_AMP_CONTROL: string  := "100PCT";
        PMA_CH1_SER_AMP_CONTROL: string  := "100PCT";
        PMA_CH1_PFD_LOOP_RESISTOR_SETTING: integer := 0;
        PMA_CH1_PD_LOOP_RESISTOR_SETTING: integer := 0;
        PMA_CH1_CDR_TEST_OUT_SELECT: string  := "FBCK";
        PMA_CH1_PI_DIV1_BP: string  := "DISABLE";
        PMA_CH1_PI_TEST_FOR_CKI: string  := "FALSE";
        PMA_CH1_PI_CURRENT_SETTING: string  := "100PCT";
        PMA_CH1_PI_FREQUENCY_SETTING: integer := 0;
        PMA_CH1_TEST_OUT_SELECT_FOR_RCK: string  := "FALSE";
        PMA_CH1_TEST_OUT_SELECT_SOURCE: string  := "SLPI1UI";
        PMA_CH1_TEST_DATA_OUT_SELECT_SOURCE: string  := "DO";
        PMA_CH1_TEST_CK_OUT_SELECT_SOURCE: string  := "DATA";
        PMA_CH1_ENABLE_SLIP1UI_MODULE: string  := "DISABLE";
        PMA_CH1_PN_SWAP_ENABLE: string  := "DISABLE";
        PMA_CH1_SIPO_BIT_SETTING: string  := "10_BIT";
        PMA_CH1_OOB_EN  : string  := "DISABLE";
        PMA_CH1_ALOS_EN : string  := "DISABLE";
        PMA_CH1_LFMODE  : string  := "HIGH";
        PMA_CH1_TSO_HS_SEL: string  := "CDR";
        PMA_CH1_LX_SELLC: string  := "RING";
        PMA_CH1_LX_RXPLL_DIVSEL45_FB: integer := 4;
        PMA_CH1_LX_RXPLL_DIVSEL_FB: integer := 2;
        PMA_CH1_LX_RXPLL_DIVSEL_REF: integer := 1;
        PMA_CH1_PICODE  : integer := 0;
        PMA_CH1_RX_REFCK_SEL: integer := 0;
        PMA_CH1_PFDLPEN_REGISTER_CONTROL_ENABLE: string  := "DISABLE";
        PMA_CH1_PFDLPEN_REGISTER_SETTING: string  := "FALSE";
        PMA_CH1_PDLPEN_REGISTER_CONTROL_ENABLE: string  := "DISABLE";
        PMA_CH1_PDLPEN_REGISTER_SETTING: string  := "FALSE";
        PMA_CH1_DIV_CHANGE_ENABLE_DELAY_TIMER: integer := 0;
        PMA_CH1_DIV_CHANGE_ENABLE_SIGNAL_GATING: string  := "FALSE";
        PMA_CH1_CDR_ALIGN_REGISTER_SETTING_VALUE: string  := "FALSE";
        PMA_CH1_FORCE_CDR_ALIGN_ENABLE: string  := "DISABLE";
        PMA_CH1_SELLC_REGISTER_SETTING_VALUE: string  := "FALSE";
        PMA_CH1_SELLC_CONTROL_BY_REGISTER: string  := "FALSE";
        PMA_CH1_REG_PLLI_LDO_VREF_SETTING: string  := "0_9V";
        PMA_CH1_REG_PLLI_LDO_BYPASS_CURRENT: integer := 0;
        PMA_CH1_REG_PLL_HSTEST_ENABLE: string  := "DISABLE";
        PMA_CH1_REG_PLL_ISNK_CURRENT_CONTROL: string  := "5U";
        PMA_CH1_REG_PLL_PFD_LOOP_CP0_CURRENT_SETTING: integer := 0;
        PMA_CH1_REG_PLL_PD_LOOP_PLLGM_SETTING: string  := "100PCT";
        PMA_CH1_REG_PLL_PFD_LOOP_CP1_CURRENT_SETTING: integer := 0;
        PMA_CH1_REG_PLL_CP0_BIAS_CONTROL: string  := "100PCT";
        PMA_CH1_REG_PLL_PD_LOOP_CP0_CURRENT_SETTING: integer := 0;
        PMA_CH1_REG_PLL_CP1_BIAS_CONTROL: string  := "100PCT";
        PMA_CH1_REG_PLL_PD_LOOP_CP1_CURRENT_SETTING: integer := 0;
        PMA_CH1_REG_PLL_CP0_CURRENT_SETTING: string  := "100PCT";
        PMA_CH1_REG_PLL_CP1_CURRENT_SETTING: string  := "100PCT";
        PMA_CH1_REG_PLL_GM1_CURRENT_SETTING: string  := "100PCT";
        PMA_CH1_REG_PLL_LC_BF2_CURRENT_SETTING: string  := "100PCT";
        PMA_CH1_REG_PLL_LC_BF2_CURRENT_SETTING_LOW: string  := "100PCT";
        PMA_CH1_REG_PLL_REG_CUR: string  := "100PCT";
        PMA_CH1_REG_PLL_LCCUR: string  := "DEFAULT";
        PMA_CH1_REG_PLL_LCOBAS: string  := "100PCT";
        PMA_CH1_REG_PLL_FB_CK_TEST_OUT_ENABLE: string  := "DISABLE";
        PMA_CH1_CDR_ALIGN_TIMER: integer := 0;
        PMA_CH1_CALIB_WAIT: integer := 1024;
        PMA_CH1_CALIB_TIMER: integer := 512;
        PMA_CH1_TOT_RANGE: integer := 0;
        PMA_CH1_SUB_RANGE: integer := 0;
        PMA_CH1_OVLP    : integer := 0;
        PMA_CH1_BIST_WAIT: integer := 1024;
        PMA_CH1_BIST_TIMER: integer := 512;
        PMA_CH1_BAND_LB : integer := 0;
        PMA_CH1_BAND_HB : integer := 0;
        PMA_CH1_FREQ_LOCK_ACCURACY: integer := 0;
        PMA_CH1_REG_SET_LC_BAND: integer := 0;
        PMA_CH1_REG_SET_VCODIV: integer := 0;
        PMA_CH1_REGISTER_SET_VCODIV_BAND_ENABLE: string  := "DISABLE";
        PMA_CH1_REG_SET_PLL_LOCK: string  := "FALSE";
        PMA_CH1_REGISTER_SET_PLL_LOCK_ENABLE: string  := "DISABLE";
        PMA_CH1_REG_SET_VCO_HI: string  := "FALSE";
        PMA_CH1_REG_SET_VCO_LO: string  := "FALSE";
        PMA_CH1_REGISTER_SET_VCO_HI_VCO_LO_ENABLE: string  := "DISABLE";
        PMA_CH1_FORCE_LC_PLL_LOOP_EN_H: string  := "DISABLE";
        PMA_CH1_FORCE_LC_PLL_LOOP_EN_L: string  := "DISABLE";
        PMA_CH1_VCO_DIV_CALI_BYPASS: string  := "FALSE";
        PMA_CH1_BIST_EN : string  := "DISABLE";
        PMA_CH1_PLL_LOOP_EN_SETTING_FROM_REGISTER_ENABLE: string  := "DISABLE";
        PMA_CH1_FREQ_DETECT_ENABLE_SOURCE: string  := "DISABLE";
        PMA_CH1_REG_SET_DIVSEL_REF: integer := 0;
        PMA_CH1_REG_SET_DIVSEL45_FB: string  := "FALSE";
        PMA_CH1_REG_SET_DIVSEL_FB: integer := 0;
        PMA_CH1_PLL_LOOP_EN_SETTING: string  := "DISABLE";
        PMA_CH1_REGISTER_SET_TXPLL_DIV_ENABLE: string  := "DISABLE";
        PMA_CH1_FORCE_RXPLL_RESET: string  := "FALSE";
        PMA_CH1_FORCE_RXPLL_ON: string  := "FALSE";
        PMA_CH1_DPCK_DIV2: string  := "FALSE";
        PMA_CH1_LFO_SETTING: integer := 0;
        PMA_CH1_ALOS_COUNTER_CLOCK_SELECTION: string  := "LOCAL";
        PMA_CH1_RX_BIAS_CURRENT_ADJUSTMENT: string  := "100PCT";
        PMA_CH1_OOB_ENTER_DELAY_SETTING: integer := 0;
        PMA_CH1_ALOS_LOW_TO_HIGH_COUNTER_SETTING: integer := 0;
        PMA_CH1_ENABLE_ALOS_RESULT_AUTOMATICALLY_ENABLE_CHANNEL: string  := "DISABLE";
        PMA_CH1_ALOS_EXIT_COUNTER_CLOCK_DIVIDER: integer := 0;
        PMA_CH1_OOB_OSCILATER_FREQUENCY_SETTING: integer := 0;
        PMA_CH1_FORCE_OOB: string  := "FALSE";
        PMA_CH1_OOB_VTH_SET: string  := "27MV";
        PMA_CH1_FORCE_DET_FORCE_ALOS_LOW: string  := "FALSE";
        PMA_CH1_ALOS_THRESHOLD_VOLTAGE: string  := "27MV";
        PMA_CH1_WAKEUP_VCM_RX_COMMON_MODE_VOLTAGE: integer := 0;
        PMA_CH1_REGR_NEGATIVE_HYSTERESIS_SETTING: string  := "100MV";
        PMA_CH1_REGL_POSITIVE_HYSTERESIS_SETTING: string  := "100MV";
        PMA_CH1_REG_EN  : string  := "DISABLE";
        PMA_CH1_REGREF_SEL: string  := "VREF";
        PMA_CH1_DC496   : string  := "39_6MHZ";
        PMA_CH1_EQ2_AC_VAR_SETTING: integer := 0;
        PMA_CH1_EQ2_AC_RES_SETTING: integer := 0;
        PMA_CH1_EQ2_DC_RESTOP_SETTING: integer := 0;
        PMA_CH1_EQ1_DC_RESTOP_SETTING: integer := 50;
        PMA_CH1_EQ1_AC_VAR_SETTING: integer := 0;
        PMA_CH1_EQ2_CURRENT_SETTING: integer := 0;
        PMA_CH1_EQ1_AC_RES_SETTING: integer := 0;
        PMA_CH1_EQ1_CURRENT_SETTING: integer := 0;
        PMA_CH1_RPLUS   : integer := 0;
        PMA_CH1_RMINUS  : integer := 0;
        PMA_CH1_RVALSET : integer := 0;
        PMA_CH1_RTERM   : integer := 0;
        PMA_CH1_DCFB_EN : string  := "DISABLE";
        PMA_CH1_DCCOUP  : string  := "FALSE";
        PMA_CH1_3G      : string  := "FALSE";
        PMA_CH2_TXDATA_WIDTH: string  := "8_BIT";
        PMA_CH2_TX_TESTPATTERN: integer := 0;
        PMA_CH2_TESTPATTERN_O_ENABLE: string  := "FALSE";
        PMA_CH2_DISABLE_BSMODE_DRVAMP: string  := "FALSE";
        PMA_CH2_FORCE_BIST_ENABLE: string  := "FALSE";
        PMA_CH2_FORCE_ELECTRICAL_IDLE: string  := "FALSE";
        PMA_CH2_FORCE_RXDCT_ENABLE: string  := "FALSE";
        PMA_CH2_FORCE_EXTLB_ENABLE: string  := "FALSE";
        PMA_CH2_DISABLE_LANE_SYNC: string  := "FALSE";
        PMA_CH2_DISABLE_ELECTRICAL_IDLE: string  := "FALSE";
        PMA_CH2_DISABLE_RXDCT_ENABLE: string  := "FALSE";
        PMA_CH2_DISABLE_EXTLB_ENABLE: string  := "FALSE";
        PMA_CH2_DISABLE_LOW_SPEED_PATH_ENABLE: string  := "FALSE";
        PMA_CH2_FORCE_LANE_ENABLE: string  := "FALSE";
        PMA_CH2_FORCE_LANE_RESETB_DISABLE: string  := "FALSE";
        PMA_CH2_RXDCT_LGBW_ENABLE: string  := "FALSE";
        PMA_CH2_RXDCT_VTH: string  := "MINUS_300MV";
        PMA_CH2_DE_EMPHASIS_ADDITIONAL_CONTROL: string  := "0DB";
        PMA_CH2_DRV_RTERM_CONTROL: string  := "100PCT";
        PMA_CH2_FDRV_AMP_CONTROL: string  := "100PCT";
        PMA_CH2_PREPC_AMP_CONTROL: string  := "100PCT";
        PMA_CH2_PREMC_AMP_CONTROL: string  := "100PCT";
        PMA_CH2_SER_AMP_CONTROL: string  := "100PCT";
        PMA_CH2_PFD_LOOP_RESISTOR_SETTING: integer := 0;
        PMA_CH2_PD_LOOP_RESISTOR_SETTING: integer := 0;
        PMA_CH2_CDR_TEST_OUT_SELECT: string  := "FBCK";
        PMA_CH2_PI_DIV1_BP: string  := "DISABLE";
        PMA_CH2_PI_TEST_FOR_CKI: string  := "FALSE";
        PMA_CH2_PI_CURRENT_SETTING: string  := "100PCT";
        PMA_CH2_PI_FREQUENCY_SETTING: integer := 0;
        PMA_CH2_TEST_OUT_SELECT_FOR_RCK: string  := "FALSE";
        PMA_CH2_TEST_OUT_SELECT_SOURCE: string  := "SLPI1UI";
        PMA_CH2_TEST_DATA_OUT_SELECT_SOURCE: string  := "DO";
        PMA_CH2_TEST_CK_OUT_SELECT_SOURCE: string  := "DATA";
        PMA_CH2_ENABLE_SLIP1UI_MODULE: string  := "DISABLE";
        PMA_CH2_PN_SWAP_ENABLE: string  := "DISABLE";
        PMA_CH2_SIPO_BIT_SETTING: string  := "10_BIT";
        PMA_CH2_OOB_EN  : string  := "DISABLE";
        PMA_CH2_ALOS_EN : string  := "DISABLE";
        PMA_CH2_LFMODE  : string  := "HIGH";
        PMA_CH2_TSO_HS_SEL: string  := "CDR";
        PMA_CH2_LX_SELLC: string  := "RING";
        PMA_CH2_LX_RXPLL_DIVSEL45_FB: integer := 4;
        PMA_CH2_LX_RXPLL_DIVSEL_FB: integer := 2;
        PMA_CH2_LX_RXPLL_DIVSEL_REF: integer := 1;
        PMA_CH2_PICODE  : integer := 0;
        PMA_CH2_RX_REFCK_SEL: integer := 0;
        PMA_CH2_PFDLPEN_REGISTER_CONTROL_ENABLE: string  := "DISABLE";
        PMA_CH2_PFDLPEN_REGISTER_SETTING: string  := "FALSE";
        PMA_CH2_PDLPEN_REGISTER_CONTROL_ENABLE: string  := "DISABLE";
        PMA_CH2_PDLPEN_REGISTER_SETTING: string  := "FALSE";
        PMA_CH2_DIV_CHANGE_ENABLE_DELAY_TIMER: integer := 0;
        PMA_CH2_DIV_CHANGE_ENABLE_SIGNAL_GATING: string  := "FALSE";
        PMA_CH2_CDR_ALIGN_REGISTER_SETTING_VALUE: string  := "FALSE";
        PMA_CH2_FORCE_CDR_ALIGN_ENABLE: string  := "DISABLE";
        PMA_CH2_SELLC_REGISTER_SETTING_VALUE: string  := "FALSE";
        PMA_CH2_SELLC_CONTROL_BY_REGISTER: string  := "FALSE";
        PMA_CH2_REG_PLLI_LDO_VREF_SETTING: string  := "0_9V";
        PMA_CH2_REG_PLLI_LDO_BYPASS_CURRENT: integer := 0;
        PMA_CH2_REG_PLL_HSTEST_ENABLE: string  := "DISABLE";
        PMA_CH2_REG_PLL_ISNK_CURRENT_CONTROL: string  := "5U";
        PMA_CH2_REG_PLL_PFD_LOOP_CP0_CURRENT_SETTING: integer := 0;
        PMA_CH2_REG_PLL_PD_LOOP_PLLGM_SETTING: string  := "100PCT";
        PMA_CH2_REG_PLL_PFD_LOOP_CP1_CURRENT_SETTING: integer := 0;
        PMA_CH2_REG_PLL_CP0_BIAS_CONTROL: string  := "100PCT";
        PMA_CH2_REG_PLL_PD_LOOP_CP0_CURRENT_SETTING: integer := 0;
        PMA_CH2_REG_PLL_CP1_BIAS_CONTROL: string  := "100PCT";
        PMA_CH2_REG_PLL_PD_LOOP_CP1_CURRENT_SETTING: integer := 0;
        PMA_CH2_REG_PLL_CP0_CURRENT_SETTING: string  := "100PCT";
        PMA_CH2_REG_PLL_CP1_CURRENT_SETTING: string  := "100PCT";
        PMA_CH2_REG_PLL_GM1_CURRENT_SETTING: string  := "100PCT";
        PMA_CH2_REG_PLL_LC_BF2_CURRENT_SETTING: string  := "100PCT";
        PMA_CH2_REG_PLL_LC_BF2_CURRENT_SETTING_LOW: string  := "100PCT";
        PMA_CH2_REG_PLL_REG_CUR: string  := "100PCT";
        PMA_CH2_REG_PLL_LCCUR: string  := "DEFAULT";
        PMA_CH2_REG_PLL_LCOBAS: string  := "100PCT";
        PMA_CH2_REG_PLL_FB_CK_TEST_OUT_ENABLE: string  := "DISABLE";
        PMA_CH2_CDR_ALIGN_TIMER: integer := 0;
        PMA_CH2_CALIB_WAIT: integer := 1024;
        PMA_CH2_CALIB_TIMER: integer := 512;
        PMA_CH2_TOT_RANGE: integer := 0;
        PMA_CH2_SUB_RANGE: integer := 0;
        PMA_CH2_OVLP    : integer := 0;
        PMA_CH2_BIST_WAIT: integer := 1024;
        PMA_CH2_BIST_TIMER: integer := 512;
        PMA_CH2_BAND_LB : integer := 0;
        PMA_CH2_BAND_HB : integer := 0;
        PMA_CH2_FREQ_LOCK_ACCURACY: integer := 0;
        PMA_CH2_REG_SET_LC_BAND: integer := 0;
        PMA_CH2_REG_SET_VCODIV: integer := 0;
        PMA_CH2_REGISTER_SET_VCODIV_BAND_ENABLE: string  := "DISABLE";
        PMA_CH2_REG_SET_PLL_LOCK: string  := "FALSE";
        PMA_CH2_REGISTER_SET_PLL_LOCK_ENABLE: string  := "DISABLE";
        PMA_CH2_REG_SET_VCO_HI: string  := "FALSE";
        PMA_CH2_REG_SET_VCO_LO: string  := "FALSE";
        PMA_CH2_REGISTER_SET_VCO_HI_VCO_LO_ENABLE: string  := "DISABLE";
        PMA_CH2_FORCE_LC_PLL_LOOP_EN_H: string  := "DISABLE";
        PMA_CH2_FORCE_LC_PLL_LOOP_EN_L: string  := "DISABLE";
        PMA_CH2_VCO_DIV_CALI_BYPASS: string  := "FALSE";
        PMA_CH2_BIST_EN : string  := "DISABLE";
        PMA_CH2_PLL_LOOP_EN_SETTING_FROM_REGISTER_ENABLE: string  := "DISABLE";
        PMA_CH2_FREQ_DETECT_ENABLE_SOURCE: string  := "DISABLE";
        PMA_CH2_REG_SET_DIVSEL_REF: integer := 0;
        PMA_CH2_REG_SET_DIVSEL45_FB: string  := "FALSE";
        PMA_CH2_REG_SET_DIVSEL_FB: integer := 0;
        PMA_CH2_PLL_LOOP_EN_SETTING: string  := "DISABLE";
        PMA_CH2_REGISTER_SET_TXPLL_DIV_ENABLE: string  := "DISABLE";
        PMA_CH2_FORCE_RXPLL_RESET: string  := "FALSE";
        PMA_CH2_FORCE_RXPLL_ON: string  := "FALSE";
        PMA_CH2_DPCK_DIV2: string  := "FALSE";
        PMA_CH2_LFO_SETTING: integer := 0;
        PMA_CH2_ALOS_COUNTER_CLOCK_SELECTION: string  := "LOCAL";
        PMA_CH2_RX_BIAS_CURRENT_ADJUSTMENT: string  := "100PCT";
        PMA_CH2_OOB_ENTER_DELAY_SETTING: integer := 0;
        PMA_CH2_ALOS_LOW_TO_HIGH_COUNTER_SETTING: integer := 0;
        PMA_CH2_ENABLE_ALOS_RESULT_AUTOMATICALLY_ENABLE_CHANNEL: string  := "DISABLE";
        PMA_CH2_ALOS_EXIT_COUNTER_CLOCK_DIVIDER: integer := 0;
        PMA_CH2_OOB_OSCILATER_FREQUENCY_SETTING: integer := 0;
        PMA_CH2_FORCE_OOB: string  := "FALSE";
        PMA_CH2_OOB_VTH_SET: string  := "27MV";
        PMA_CH2_FORCE_DET_FORCE_ALOS_LOW: string  := "FALSE";
        PMA_CH2_ALOS_THRESHOLD_VOLTAGE: string  := "27MV";
        PMA_CH2_WAKEUP_VCM_RX_COMMON_MODE_VOLTAGE: integer := 0;
        PMA_CH2_REGR_NEGATIVE_HYSTERESIS_SETTING: string  := "100MV";
        PMA_CH2_REGL_POSITIVE_HYSTERESIS_SETTING: string  := "100MV";
        PMA_CH2_REG_EN  : string  := "DISABLE";
        PMA_CH2_REGREF_SEL: string  := "VREF";
        PMA_CH2_DC496   : string  := "39_6MHZ";
        PMA_CH2_EQ2_AC_VAR_SETTING: integer := 0;
        PMA_CH2_EQ2_AC_RES_SETTING: integer := 0;
        PMA_CH2_EQ2_DC_RESTOP_SETTING: integer := 0;
        PMA_CH2_EQ1_DC_RESTOP_SETTING: integer := 50;
        PMA_CH2_EQ1_AC_VAR_SETTING: integer := 0;
        PMA_CH2_EQ2_CURRENT_SETTING: integer := 0;
        PMA_CH2_EQ1_AC_RES_SETTING: integer := 0;
        PMA_CH2_EQ1_CURRENT_SETTING: integer := 0;
        PMA_CH2_RPLUS   : integer := 0;
        PMA_CH2_RMINUS  : integer := 0;
        PMA_CH2_RVALSET : integer := 0;
        PMA_CH2_RTERM   : integer := 0;
        PMA_CH2_DCFB_EN : string  := "DISABLE";
        PMA_CH2_DCCOUP  : string  := "FALSE";
        PMA_CH2_3G      : string  := "FALSE";
        PMA_CH3_TXDATA_WIDTH: string  := "8_BIT";
        PMA_CH3_TX_TESTPATTERN: integer := 0;
        PMA_CH3_TESTPATTERN_O_ENABLE: string  := "FALSE";
        PMA_CH3_DISABLE_BSMODE_DRVAMP: string  := "FALSE";
        PMA_CH3_FORCE_BIST_ENABLE: string  := "FALSE";
        PMA_CH3_FORCE_ELECTRICAL_IDLE: string  := "FALSE";
        PMA_CH3_FORCE_RXDCT_ENABLE: string  := "FALSE";
        PMA_CH3_FORCE_EXTLB_ENABLE: string  := "FALSE";
        PMA_CH3_DISABLE_LANE_SYNC: string  := "FALSE";
        PMA_CH3_DISABLE_ELECTRICAL_IDLE: string  := "FALSE";
        PMA_CH3_DISABLE_RXDCT_ENABLE: string  := "FALSE";
        PMA_CH3_DISABLE_EXTLB_ENABLE: string  := "FALSE";
        PMA_CH3_DISABLE_LOW_SPEED_PATH_ENABLE: string  := "FALSE";
        PMA_CH3_FORCE_LANE_ENABLE: string  := "FALSE";
        PMA_CH3_FORCE_LANE_RESETB_DISABLE: string  := "FALSE";
        PMA_CH3_RXDCT_LGBW_ENABLE: string  := "FALSE";
        PMA_CH3_RXDCT_VTH: string  := "MINUS_300MV";
        PMA_CH3_DE_EMPHASIS_ADDITIONAL_CONTROL: string  := "0DB";
        PMA_CH3_DRV_RTERM_CONTROL: string  := "100PCT";
        PMA_CH3_FDRV_AMP_CONTROL: string  := "100PCT";
        PMA_CH3_PREPC_AMP_CONTROL: string  := "100PCT";
        PMA_CH3_PREMC_AMP_CONTROL: string  := "100PCT";
        PMA_CH3_SER_AMP_CONTROL: string  := "100PCT";
        PMA_CH3_PFD_LOOP_RESISTOR_SETTING: integer := 0;
        PMA_CH3_PD_LOOP_RESISTOR_SETTING: integer := 0;
        PMA_CH3_CDR_TEST_OUT_SELECT: string  := "FBCK";
        PMA_CH3_PI_DIV1_BP: string  := "DISABLE";
        PMA_CH3_PI_TEST_FOR_CKI: string  := "FALSE";
        PMA_CH3_PI_CURRENT_SETTING: string  := "100PCT";
        PMA_CH3_PI_FREQUENCY_SETTING: integer := 0;
        PMA_CH3_TEST_OUT_SELECT_FOR_RCK: string  := "FALSE";
        PMA_CH3_TEST_OUT_SELECT_SOURCE: string  := "SLPI1UI";
        PMA_CH3_TEST_DATA_OUT_SELECT_SOURCE: string  := "DO";
        PMA_CH3_TEST_CK_OUT_SELECT_SOURCE: string  := "DATA";
        PMA_CH3_ENABLE_SLIP1UI_MODULE: string  := "DISABLE";
        PMA_CH3_PN_SWAP_ENABLE: string  := "DISABLE";
        PMA_CH3_SIPO_BIT_SETTING: string  := "10_BIT";
        PMA_CH3_OOB_EN  : string  := "DISABLE";
        PMA_CH3_ALOS_EN : string  := "DISABLE";
        PMA_CH3_LFMODE  : string  := "HIGH";
        PMA_CH3_TSO_HS_SEL: string  := "CDR";
        PMA_CH3_LX_SELLC: string  := "RING";
        PMA_CH3_LX_RXPLL_DIVSEL45_FB: integer := 4;
        PMA_CH3_LX_RXPLL_DIVSEL_FB: integer := 2;
        PMA_CH3_LX_RXPLL_DIVSEL_REF: integer := 1;
        PMA_CH3_PICODE  : integer := 0;
        PMA_CH3_RX_REFCK_SEL: integer := 0;
        PMA_CH3_PFDLPEN_REGISTER_CONTROL_ENABLE: string  := "DISABLE";
        PMA_CH3_PFDLPEN_REGISTER_SETTING: string  := "FALSE";
        PMA_CH3_PDLPEN_REGISTER_CONTROL_ENABLE: string  := "DISABLE";
        PMA_CH3_PDLPEN_REGISTER_SETTING: string  := "FALSE";
        PMA_CH3_DIV_CHANGE_ENABLE_DELAY_TIMER: integer := 0;
        PMA_CH3_DIV_CHANGE_ENABLE_SIGNAL_GATING: string  := "FALSE";
        PMA_CH3_CDR_ALIGN_REGISTER_SETTING_VALUE: string  := "FALSE";
        PMA_CH3_FORCE_CDR_ALIGN_ENABLE: string  := "DISABLE";
        PMA_CH3_SELLC_REGISTER_SETTING_VALUE: string  := "FALSE";
        PMA_CH3_SELLC_CONTROL_BY_REGISTER: string  := "FALSE";
        PMA_CH3_REG_PLLI_LDO_VREF_SETTING: string  := "0_9V";
        PMA_CH3_REG_PLLI_LDO_BYPASS_CURRENT: integer := 0;
        PMA_CH3_REG_PLL_HSTEST_ENABLE: string  := "DISABLE";
        PMA_CH3_REG_PLL_ISNK_CURRENT_CONTROL: string  := "5U";
        PMA_CH3_REG_PLL_PFD_LOOP_CP0_CURRENT_SETTING: integer := 0;
        PMA_CH3_REG_PLL_PD_LOOP_PLLGM_SETTING: string  := "100PCT";
        PMA_CH3_REG_PLL_PFD_LOOP_CP1_CURRENT_SETTING: integer := 0;
        PMA_CH3_REG_PLL_CP0_BIAS_CONTROL: string  := "100PCT";
        PMA_CH3_REG_PLL_PD_LOOP_CP0_CURRENT_SETTING: integer := 0;
        PMA_CH3_REG_PLL_CP1_BIAS_CONTROL: string  := "100PCT";
        PMA_CH3_REG_PLL_PD_LOOP_CP1_CURRENT_SETTING: integer := 0;
        PMA_CH3_REG_PLL_CP0_CURRENT_SETTING: string  := "100PCT";
        PMA_CH3_REG_PLL_CP1_CURRENT_SETTING: string  := "100PCT";
        PMA_CH3_REG_PLL_GM1_CURRENT_SETTING: string  := "100PCT";
        PMA_CH3_REG_PLL_LC_BF2_CURRENT_SETTING: string  := "100PCT";
        PMA_CH3_REG_PLL_LC_BF2_CURRENT_SETTING_LOW: string  := "100PCT";
        PMA_CH3_REG_PLL_REG_CUR: string  := "100PCT";
        PMA_CH3_REG_PLL_LCCUR: string  := "DEFAULT";
        PMA_CH3_REG_PLL_LCOBAS: string  := "100PCT";
        PMA_CH3_REG_PLL_FB_CK_TEST_OUT_ENABLE: string  := "DISABLE";
        PMA_CH3_CDR_ALIGN_TIMER: integer := 0;
        PMA_CH3_CALIB_WAIT: integer := 1024;
        PMA_CH3_CALIB_TIMER: integer := 512;
        PMA_CH3_TOT_RANGE: integer := 0;
        PMA_CH3_SUB_RANGE: integer := 0;
        PMA_CH3_OVLP    : integer := 0;
        PMA_CH3_BIST_WAIT: integer := 1024;
        PMA_CH3_BIST_TIMER: integer := 512;
        PMA_CH3_BAND_LB : integer := 0;
        PMA_CH3_BAND_HB : integer := 0;
        PMA_CH3_FREQ_LOCK_ACCURACY: integer := 0;
        PMA_CH3_REG_SET_LC_BAND: integer := 0;
        PMA_CH3_REG_SET_VCODIV: integer := 0;
        PMA_CH3_REGISTER_SET_VCODIV_BAND_ENABLE: string  := "DISABLE";
        PMA_CH3_REG_SET_PLL_LOCK: string  := "FALSE";
        PMA_CH3_REGISTER_SET_PLL_LOCK_ENABLE: string  := "DISABLE";
        PMA_CH3_REG_SET_VCO_HI: string  := "FALSE";
        PMA_CH3_REG_SET_VCO_LO: string  := "FALSE";
        PMA_CH3_REGISTER_SET_VCO_HI_VCO_LO_ENABLE: string  := "DISABLE";
        PMA_CH3_FORCE_LC_PLL_LOOP_EN_H: string  := "DISABLE";
        PMA_CH3_FORCE_LC_PLL_LOOP_EN_L: string  := "DISABLE";
        PMA_CH3_VCO_DIV_CALI_BYPASS: string  := "FALSE";
        PMA_CH3_BIST_EN : string  := "DISABLE";
        PMA_CH3_PLL_LOOP_EN_SETTING_FROM_REGISTER_ENABLE: string  := "DISABLE";
        PMA_CH3_FREQ_DETECT_ENABLE_SOURCE: string  := "DISABLE";
        PMA_CH3_REG_SET_DIVSEL_REF: integer := 0;
        PMA_CH3_REG_SET_DIVSEL45_FB: string  := "FALSE";
        PMA_CH3_REG_SET_DIVSEL_FB: integer := 0;
        PMA_CH3_PLL_LOOP_EN_SETTING: string  := "DISABLE";
        PMA_CH3_REGISTER_SET_TXPLL_DIV_ENABLE: string  := "DISABLE";
        PMA_CH3_FORCE_RXPLL_RESET: string  := "FALSE";
        PMA_CH3_FORCE_RXPLL_ON: string  := "FALSE";
        PMA_CH3_DPCK_DIV2: string  := "FALSE";
        PMA_CH3_LFO_SETTING: integer := 0;
        PMA_CH3_ALOS_COUNTER_CLOCK_SELECTION: string  := "LOCAL";
        PMA_CH3_RX_BIAS_CURRENT_ADJUSTMENT: string  := "100PCT";
        PMA_CH3_OOB_ENTER_DELAY_SETTING: integer := 0;
        PMA_CH3_ALOS_LOW_TO_HIGH_COUNTER_SETTING: integer := 0;
        PMA_CH3_ENABLE_ALOS_RESULT_AUTOMATICALLY_ENABLE_CHANNEL: string  := "DISABLE";
        PMA_CH3_ALOS_EXIT_COUNTER_CLOCK_DIVIDER: integer := 0;
        PMA_CH3_OOB_OSCILATER_FREQUENCY_SETTING: integer := 0;
        PMA_CH3_FORCE_OOB: string  := "FALSE";
        PMA_CH3_OOB_VTH_SET: string  := "27MV";
        PMA_CH3_FORCE_DET_FORCE_ALOS_LOW: string  := "FALSE";
        PMA_CH3_ALOS_THRESHOLD_VOLTAGE: string  := "27MV";
        PMA_CH3_WAKEUP_VCM_RX_COMMON_MODE_VOLTAGE: integer := 0;
        PMA_CH3_REGR_NEGATIVE_HYSTERESIS_SETTING: string  := "100MV";
        PMA_CH3_REGL_POSITIVE_HYSTERESIS_SETTING: string  := "100MV";
        PMA_CH3_REG_EN  : string  := "DISABLE";
        PMA_CH3_REGREF_SEL: string  := "VREF";
        PMA_CH3_DC496   : string  := "39_6MHZ";
        PMA_CH3_EQ2_AC_VAR_SETTING: integer := 0;
        PMA_CH3_EQ2_AC_RES_SETTING: integer := 0;
        PMA_CH3_EQ2_DC_RESTOP_SETTING: integer := 0;
        PMA_CH3_EQ1_DC_RESTOP_SETTING: integer := 50;
        PMA_CH3_EQ1_AC_VAR_SETTING: integer := 0;
        PMA_CH3_EQ2_CURRENT_SETTING: integer := 0;
        PMA_CH3_EQ1_AC_RES_SETTING: integer := 0;
        PMA_CH3_EQ1_CURRENT_SETTING: integer := 0;
        PMA_CH3_RPLUS   : integer := 0;
        PMA_CH3_RMINUS  : integer := 0;
        PMA_CH3_RVALSET : integer := 0;
        PMA_CH3_RTERM   : integer := 0;
        PMA_CH3_DCFB_EN : string  := "DISABLE";
        PMA_CH3_DCCOUP  : string  := "FALSE";
        PMA_CH3_3G      : string  := "FALSE";
        PMA_QUAD_TURN_ON_BANDGAP_AT_AOS_ON: string  := "FALSE";
        PMA_QUAD_TURN_ON_BANDGAP_AT_RX_DETECTION_ON: string  := "FALSE";
        PMA_QUAD_TURN_ON_BANDGAP_AT_BOUNDARY_SCAN_ON: string  := "FALSE";
        PMA_QUAD_CFG_HSST_RSTN: string  := "FALSE";
        PMA_QUAD_SELECT_LANE_TCK_FOR_QUAD_SYNC: string  := "LANE0";
        PMA_QUAD_CK_REN : string  := "DISABLE";
        PMA_QUAD_C1_EN  : string  := "DISABLE";
        PMA_QUAD_C2_EN  : string  := "DISABLE";
        PMA_QUAD_CLK_DIVIDER_SETTING_FROM_25M_TO_200K: integer := 0;
        PMA_QUAD_ACMODE_SCANMODE_EN: string  := "DISABLE";
        PMA_QUAD_REGISTER_ACMODE: string  := "FALSE";
        PMA_QUAD_REGISTER_SCANMODE: string  := "FALSE";
        PMA_QUAD_REFCK2CORE_EN: string  := "DISABLE";
        PMA_QUAD_REG_EN : string  := "DISABLE";
        PMA_QUAD_REGR   : string  := "100MV";
        PMA_QUAD_REGL   : string  := "100MV";
        PMA_QUAD_DPCK_SEL: integer := 0;
        PMA_QUAD_TX_REFCK_SEL: string  := "FALSE";
        PMA_QUAD_REFCK_SRC_SEL: string  := "FALSE";
        PMA_QUAD_RREFCK_PWRUP: string  := "FALSE";
        PMA_QUAD_REFCK_SK_SEL: string  := "BOTH";
        PMA_QUAD_REFCK_DIV2_SEL: string  := "FALSE";
        PMA_QUAD_REFCK_TO_NQ_EN: string  := "DISABLE";
        PMA_QUAD_AUXI_ADJ: string  := "100PCT";
        PMA_QUAD_DC496  : string  := "39_6MHZ";
        PMA_QUAD_REG_FDET_TIMER: integer := 512;
        PMA_QUAD_FREQ_LKO: string  := "10PCT";
        PMA_QUAD_FREQ_LKI: string  := "10PCT";
        PMA_QUAD_CLOCK_SRC_SEL: string  := "LOCAL";
        PMA_QUAD_FRE_DET_EN: string  := "DISABLE";
        PMA_QUAD_TSO_LS_SEL: integer := 0;
        PMA_QUAD_TXPLL_START: string  := "FALSE";
        PMA_QUAD_VCODIV : integer := 0;
        PMA_QUAD_LC_BAND: integer := 0;
        PMA_QUAD_SET_VCO_HI: string  := "FALSE";
        PMA_QUAD_SET_VCO_LO: string  := "FALSE";
        PMA_QUAD_CALIB_FAIL: string  := "FALSE";
        PMA_QUAD_CALIB_DONE: string  := "FALSE";
        PMA_QUAD_BIST_DONE: string  := "FALSE";
        PMA_QUAD_TOTRANGE_FAIL: string  := "FALSE";
        PMA_QUAD_SUBRANGE_FAIL: string  := "FALSE";
        PMA_QUAD_OVLP_FAIL: string  := "FALSE";
        PMA_QUAD_TXPLL_LOCK: string  := "FALSE";
        PMA_QUAD_TXPLL_LOOP_ENABLE: string  := "DISABLE";
        PMA_QUAD_TXPLL_DIVSEL_REF_STA: integer := 0;
        PMA_QUAD_TXPLL_DIVSEL45_FB_STA: string  := "FALSE";
        PMA_QUAD_TXPLL_DIVSEL_FB_STA: integer := 0;
        PMA_QUAD_TXPLL_DIVSEL45_FB: string  := "FALSE";
        PMA_QUAD_TXPLL_DIVSEL_FB: integer := 0;
        PMA_QUAD_TXPLL_DIVSEL_REF: integer := 0;
        PMA_QUAD_REG_DISABLE_HOLDCLK: string  := "DISABLE";
        PMA_QUAD_REG_DISABLE_SYNC: string  := "DISABLE";
        PMA_QUAD_FORCE_OUTPUT_PLL_LOCK: string  := "FALSE";
        PMA_QUAD_REGISTER_SET_SYNCTCK_SEL_ENABLE: string  := "DISABLE";
        PMA_QUAD_REG_SET_SYNCTCK_SEL: string  := "LANE0";
        PMA_QUAD_CK4TEST_OUTPUT_ENABLE: string  := "DISABLE";
        PMA_QUAD_RSTGENBAS: string  := "100PCT";
        PMA_QUAD_LCBUFBAS: string  := "100PCT";
        PMA_QUAD_REGISTER_SET_CPCUR_ENABEL: string  := "DISABLE";
        PMA_QUAD_REG_SET_CPCUR: integer := 0;
        PMA_QUAD_CPBAS  : string  := "100PCT";
        PMA_QUAD_LCOBAS : string  := "100PCT";
        PMA_QUAD_LCCUR  : string  := "DEFAULT";
        PMA_QUAD_ENABLE_REGISTER_SETTING_BAND: string  := "DISABLE";
        PMA_QUAD_CALIB_WAIT: integer := 1024;
        PMA_QUAD_CALIB_TIMER: integer := 512;
        PMA_QUAD_TOT_RANGE: integer := 0;
        PMA_QUAD_SUB_RANGE: integer := 0;
        PMA_QUAD_OVLP   : integer := 0;
        PMA_QUAD_BIST_WAIT: integer := 1024;
        PMA_QUAD_BIST_TIMER: integer := 512;
        PMA_QUAD_BAND_LB: integer := 0;
        PMA_QUAD_BAND_HB: integer := 0;
        PMA_QUAD_FREQ_LOCK_ACCURACY: integer := 0;
        PMA_QUAD_REG_SET_LC_BAND: integer := 0;
        PMA_QUAD_REG_SET_VCODIV: integer := 0;
        PMA_QUAD_REGISTER_SET_VCODIV_BAND_ENABLE: string  := "DISABLE";
        PMA_QUAD_REG_SET_PLL_LOCK: string  := "FALSE";
        PMA_QUAD_REGISTER_SET_PLL_LOCK_ENABLE: string  := "DISABLE";
        PMA_QUAD_REG_SET_VCO_HI: string  := "FALSE";
        PMA_QUAD_REG_SET_VCO_LO: string  := "FALSE";
        PMA_QUAD_REGISTER_SET_VCO_HI_VCO_LO_ENABLE: string  := "DISABLE";
        PMA_QUAD_FORCE_LC_PLL_LOOP_EN_H: string  := "DISABLE";
        PMA_QUAD_FORCE_LC_PLL_LOOP_EN_L: string  := "DISABLE";
        PMA_QUAD_VCO_DIV_CALI_BYPASS: string  := "FALSE";
        PMA_QUAD_BIST_EN: string  := "DISABLE";
        PMA_QUAD_ENABLE_TXPLL_BIST_BLOCK_CLOCKS: string  := "DISABLE";
        PMA_QUAD_LF_TESTBY2: string  := "DISABLE";
        PMA_QUAD_REG_SET_DIVSEL_REF: integer := 0;
        PMA_QUAD_REG_SET_DIVSEL45_FB: string  := "FALSE";
        PMA_QUAD_REG_SET_DIVSEL_FB: integer := 0;
        PMA_QUAD_LF_TEST_EN: string  := "DISABLE";
        PMA_QUAD_REGISTER_SET_TXPLL_DIV_ENABLE: string  := "DISABLE";
        PMA_QUAD_FORCE_TXPLL_RESET: string  := "FALSE";
        PMA_QUAD_FORCE_TXPLL_ON: string  := "FALSE";
        CLK_ALIGNER_RX0 : integer := 0;
        CLK_ALIGNER_RX1 : integer := 0;
        CLK_ALIGNER_RX2 : integer := 0;
        CLK_ALIGNER_RX3 : integer := 0;
        CLK_ALIGNER_TX0 : integer := 0;
        CLK_ALIGNER_TX1 : integer := 0;
        CLK_ALIGNER_TX2 : integer := 0;
        CLK_ALIGNER_TX3 : integer := 0;
        DYN_DLY_EN_RX0  : string  := "FALSE";
        DYN_DLY_EN_RX1  : string  := "FALSE";
        DYN_DLY_EN_RX2  : string  := "FALSE";
        DYN_DLY_EN_RX3  : string  := "FALSE";
        DYN_DLY_EN_TX0  : string  := "FALSE";
        DYN_DLY_EN_TX1  : string  := "FALSE";
        DYN_DLY_EN_TX2  : string  := "FALSE";
        DYN_DLY_EN_TX3  : string  := "FALSE";
        DYN_DLY_SEL_RX0 : string  := "FALSE";
        DYN_DLY_SEL_RX1 : string  := "FALSE";
        DYN_DLY_SEL_RX2 : string  := "FALSE";
        DYN_DLY_SEL_RX3 : string  := "FALSE";
        DYN_DLY_SEL_TX0 : string  := "FALSE";
        DYN_DLY_SEL_TX1 : string  := "FALSE";
        DYN_DLY_SEL_TX2 : string  := "FALSE";
        DYN_DLY_SEL_TX3 : string  := "FALSE";
        CLK_ALIGNER_RSTN_RX: integer := 0;
        CLK_ALIGNER_RSTN_TX: integer := 0;
        LX_BISTLB_EN    : integer := 0;
        LX_ELECIDLE_EN_MSB: integer := 0;
        LX_EXTLB_EN     : integer := 0;
        LX_RXDCT_EN     : integer := 0;
        LX_TX_LFMODE    : integer := 0;
        RX_LANE_POWERUP : integer := 0;
        TX_LANE_POWERUP : integer := 0;
        PLL_RSTN        : string  := "FALSE";
        PLLPOWERDOWN    : string  := "FALSE";
        QUAD_PWRUP      : string  := "FALSE";
        GRSN_DIS        : string  := "FALSE";
        HSST_RSTN       : string  := "FALSE";
        CFG_RSTN        : string  := "FALSE"
    );
    port(
        P_AFTER_CTC_RCLK_EN_COUT: out    vl_logic;
        P_AFTER_CTC_RCLK_EN_GB_COUT: out    vl_logic;
        P_APATTERN_MATCH_LSB_COUT: out    vl_logic;
        P_APATTERN_MATCH_MSB_COUT: out    vl_logic;
        P_APATTERN_SEACHING_PROC_COUT: out    vl_logic;
        P_APATTERN_STATUS_COUT: out    vl_logic;
        P_BRIDGE_RCLK_EN_COUT: out    vl_logic;
        P_BRIDGE_TCLK_EN_COUT: out    vl_logic;
        P_CB_RCLK_EN_COUT: out    vl_logic;
        P_CFG_INT       : out    vl_logic;
        P_CFG_READY     : out    vl_logic;
        P_CTC_RD_FIFO_COUT: out    vl_logic;
        P_L0TXN         : out    vl_logic;
        P_L0TXP         : out    vl_logic;
        P_L1TXN         : out    vl_logic;
        P_L1TXP         : out    vl_logic;
        P_L2TXN         : out    vl_logic;
        P_L2TXP         : out    vl_logic;
        P_L3TXN         : out    vl_logic;
        P_L3TXP         : out    vl_logic;
        P_LX_ALOS_STA_0 : out    vl_logic;
        P_LX_ALOS_STA_1 : out    vl_logic;
        P_LX_ALOS_STA_2 : out    vl_logic;
        P_LX_ALOS_STA_3 : out    vl_logic;
        P_LX_CDR_ALIGN_0: out    vl_logic;
        P_LX_CDR_ALIGN_1: out    vl_logic;
        P_LX_CDR_ALIGN_2: out    vl_logic;
        P_LX_CDR_ALIGN_3: out    vl_logic;
        P_LX_LFO_0      : out    vl_logic;
        P_LX_LFO_1      : out    vl_logic;
        P_LX_LFO_2      : out    vl_logic;
        P_LX_LFO_3      : out    vl_logic;
        P_LX_OOB_STA_0  : out    vl_logic;
        P_LX_OOB_STA_1  : out    vl_logic;
        P_LX_OOB_STA_2  : out    vl_logic;
        P_LX_OOB_STA_3  : out    vl_logic;
        P_LX_RXDCT_DONE_0: out    vl_logic;
        P_LX_RXDCT_DONE_1: out    vl_logic;
        P_LX_RXDCT_DONE_2: out    vl_logic;
        P_LX_RXDCT_DONE_3: out    vl_logic;
        P_LX_RXDCT_OUT_0: out    vl_logic;
        P_LX_RXDCT_OUT_1: out    vl_logic;
        P_LX_RXDCT_OUT_2: out    vl_logic;
        P_LX_RXDCT_OUT_3: out    vl_logic;
        P_PCS_TCLK_EN_COUT: out    vl_logic;
        P_PLL_LOCK      : out    vl_logic;
        P_REFCK2CORE    : out    vl_logic;
        P_REFCK_2NMQ    : out    vl_logic;
        P_REFCK_2NPQ    : out    vl_logic;
        P_REXT          : out    vl_logic;
        P_RFIFO_EN_AFTER_CTC_COUT: out    vl_logic;
        P_RFIFO_EN_AFTER_CTC_GB_COUT: out    vl_logic;
        P_RFIFO_EN_BRIDGE_COUT: out    vl_logic;
        P_RFIFO_EN_CB_COUT: out    vl_logic;
        P_SKIP_ADD_LSB_MCB_COUT: out    vl_logic;
        P_SKIP_ADD_MCB_COUT: out    vl_logic;
        P_SKIP_DEL_LSB_MCB_COUT: out    vl_logic;
        P_SKIP_DEL_MCB_COUT: out    vl_logic;
        P_TFIFO_EN_BRIDGE_COUT: out    vl_logic;
        P_TFIFO_EN_PCS_TX_COUT: out    vl_logic;
        P_TSO_LS_OUT    : out    vl_logic;
        P_AFTER_CTC_RCLK_EN_CIN: in     vl_logic;
        P_AFTER_CTC_RCLK_EN_GB_CIN: in     vl_logic;
        P_APATTERN_MATCH_LSB_CIN: in     vl_logic;
        P_APATTERN_MATCH_MSB_CIN: in     vl_logic;
        P_APATTERN_SEACHING_PROC_CIN: in     vl_logic;
        P_APATTERN_STATUS_CIN: in     vl_logic;
        P_BRIDGE_RCLK_EN_CIN: in     vl_logic;
        P_BRIDGE_TCLK_EN_CIN: in     vl_logic;
        P_CB_RCLK_EN_CIN: in     vl_logic;
        P_CFG_CLK       : in     vl_logic;
        P_CFG_ENABLE    : in     vl_logic;
        P_CFG_RSTN      : in     vl_logic;
        P_CFG_WRITE     : in     vl_logic;
        P_COMPRESSION_MODE: in     vl_logic;
        P_CTC_RD_FIFO_CIN: in     vl_logic;
        P_HSST_RSTN     : in     vl_logic;
        P_L0RXN         : in     vl_logic;
        P_L0RXP         : in     vl_logic;
        P_L1RXN         : in     vl_logic;
        P_L1RXP         : in     vl_logic;
        P_L2RXN         : in     vl_logic;
        P_L2RXP         : in     vl_logic;
        P_L3RXN         : in     vl_logic;
        P_L3RXP         : in     vl_logic;
        P_LANE_SYNC_EN_0: in     vl_logic;
        P_LANE_SYNC_EN_1: in     vl_logic;
        P_LANE_SYNC_EN_2: in     vl_logic;
        P_LANE_SYNC_EN_3: in     vl_logic;
        P_LX_LFD_FRCORE_0: in     vl_logic;
        P_LX_LFD_FRCORE_1: in     vl_logic;
        P_LX_LFD_FRCORE_2: in     vl_logic;
        P_LX_LFD_FRCORE_3: in     vl_logic;
        P_LX_RX_CKDIV_DYNSEL_0: in     vl_logic;
        P_LX_RX_CKDIV_DYNSEL_1: in     vl_logic;
        P_LX_RX_CKDIV_DYNSEL_2: in     vl_logic;
        P_LX_RX_CKDIV_DYNSEL_3: in     vl_logic;
        P_MCB_CLK_FRNQ  : in     vl_logic;
        P_PCS_RX_RSTN_0 : in     vl_logic;
        P_PCS_RX_RSTN_1 : in     vl_logic;
        P_PCS_RX_RSTN_2 : in     vl_logic;
        P_PCS_RX_RSTN_3 : in     vl_logic;
        P_PCS_TCLK_EN_CIN: in     vl_logic;
        P_PCS_TX_RSTN_0 : in     vl_logic;
        P_PCS_TX_RSTN_1 : in     vl_logic;
        P_PCS_TX_RSTN_2 : in     vl_logic;
        P_PCS_TX_RSTN_3 : in     vl_logic;
        P_PLL_BYPASS    : in     vl_logic;
        P_PLL_REF_CLK   : in     vl_logic;
        P_PLL_RESET     : in     vl_logic;
        P_PLL_RSTN      : in     vl_logic;
        P_PLLPOWERDOWN  : in     vl_logic;
        P_QUAD_PWRUP    : in     vl_logic;
        P_REFCK_FRNMQ   : in     vl_logic;
        P_REFCK_FRNPQ   : in     vl_logic;
        P_REFCKN        : in     vl_logic;
        P_REFCKP        : in     vl_logic;
        P_RFIFO_EN_AFTER_CTC_CIN: in     vl_logic;
        P_RFIFO_EN_AFTER_CTC_GB_CIN: in     vl_logic;
        P_RFIFO_EN_BRIDGE_CIN: in     vl_logic;
        P_RFIFO_EN_CB_CIN: in     vl_logic;
        P_RX0_CLK_FR_CORE: in     vl_logic;
        P_RX1_CLK_FR_CORE: in     vl_logic;
        P_RX2_CLK_FR_CORE: in     vl_logic;
        P_RX3_CLK_FR_CORE: in     vl_logic;
        P_RX_PLL_RSTN_0 : in     vl_logic;
        P_RX_PLL_RSTN_1 : in     vl_logic;
        P_RX_PLL_RSTN_2 : in     vl_logic;
        P_RX_PLL_RSTN_3 : in     vl_logic;
        P_RX_PMA_RSTN_0 : in     vl_logic;
        P_RX_PMA_RSTN_1 : in     vl_logic;
        P_RX_PMA_RSTN_2 : in     vl_logic;
        P_RX_PMA_RSTN_3 : in     vl_logic;
        P_RX_REF_CLK_0  : in     vl_logic;
        P_RX_REF_CLK_1  : in     vl_logic;
        P_RX_REF_CLK_2  : in     vl_logic;
        P_RX_REF_CLK_3  : in     vl_logic;
        P_SEL_SYNC_NXQ  : in     vl_logic;
        P_SKIP_ADD_LSB_MCB_CIN: in     vl_logic;
        P_SKIP_ADD_MCB_CIN: in     vl_logic;
        P_SKIP_DEL_LSB_MCB_CIN: in     vl_logic;
        P_SKIP_DEL_MCB_CIN: in     vl_logic;
        P_SYNC_TOGGLE   : in     vl_logic;
        P_TFIFO_EN_BRIDGE_CIN: in     vl_logic;
        P_TFIFO_EN_PCS_TX_CIN: in     vl_logic;
        P_TWOQUAD_SYNC_EN: in     vl_logic;
        P_TX0_CLK_FR_CORE: in     vl_logic;
        P_TX1_CLK_FR_CORE: in     vl_logic;
        P_TX2_CLK_FR_CORE: in     vl_logic;
        P_TX3_CLK_FR_CORE: in     vl_logic;
        P_TX_PMA_RSTN_0 : in     vl_logic;
        P_TX_PMA_RSTN_1 : in     vl_logic;
        P_TX_PMA_RSTN_2 : in     vl_logic;
        P_TX_PMA_RSTN_3 : in     vl_logic;
        P_TXCKDIV_DYNSEL: in     vl_logic;
        P_RDATA_0       : out    vl_logic_vector(46 downto 0);
        P_RDATA_1       : out    vl_logic_vector(46 downto 0);
        P_PCS_LSM_SYNCED: out    vl_logic_vector(3 downto 0);
        P_RDATA_2       : out    vl_logic_vector(46 downto 0);
        P_ALIGN_TX      : out    vl_logic_vector(3 downto 0);
        P_ALIGN_RX      : out    vl_logic_vector(3 downto 0);
        P_RDATA_3       : out    vl_logic_vector(46 downto 0);
        P_CLK2CORE_TX   : out    vl_logic_vector(3 downto 0);
        P_CLK2CORE_RX   : out    vl_logic_vector(3 downto 0);
        P_CFG_RDATA     : out    vl_logic_vector(7 downto 0);
        P_PCS_RX_MCB_STATUS: out    vl_logic_vector(3 downto 0);
        P_CIM_CLK_ALIGNER_TX3: in     vl_logic_vector(7 downto 0);
        P_TX_CKDIV_1    : in     vl_logic_vector(1 downto 0);
        P_LX_DEEMP_CTL_1: in     vl_logic_vector(2 downto 0);
        P_LX_TX_LFMODE  : in     vl_logic_vector(3 downto 0);
        P_LX_AMP_CTL_0  : in     vl_logic_vector(3 downto 0);
        P_LX_RXDCT_EN   : in     vl_logic_vector(3 downto 0);
        P_TX_CKDIV_0    : in     vl_logic_vector(1 downto 0);
        P_LX_RX_CKDIV_3 : in     vl_logic_vector(1 downto 0);
        P_PCS_MCB_EXT_EN: in     vl_logic_vector(3 downto 0);
        P_CIM_CLK_ALIGNER_TX0: in     vl_logic_vector(7 downto 0);
        P_LX_DEEMP_CTL_0: in     vl_logic_vector(2 downto 0);
        P_TDATA_2       : in     vl_logic_vector(43 downto 0);
        P_LX_AMP_CTL_3  : in     vl_logic_vector(3 downto 0);
        P_CIM_CLK_ALIGNER_TX1: in     vl_logic_vector(7 downto 0);
        P_LX_RX_CKDIV_2 : in     vl_logic_vector(1 downto 0);
        P_CEB_ADETECT_EN: in     vl_logic_vector(3 downto 0);
        P_TX_CKDIV_3    : in     vl_logic_vector(1 downto 0);
        P_CIM_CLK_ALIGNER_RX1: in     vl_logic_vector(7 downto 0);
        P_CFG_WDATA     : in     vl_logic_vector(7 downto 0);
        P_TX_LANE_POWERUP: in     vl_logic_vector(3 downto 0);
        P_TDATA_1       : in     vl_logic_vector(43 downto 0);
        P_LX_EXTLB_EN   : in     vl_logic_vector(3 downto 0);
        P_CFG_ADDR      : in     vl_logic_vector(15 downto 0);
        P_CIM_CLK_ALIGNER_RX0: in     vl_logic_vector(7 downto 0);
        P_LX_ELECIDLE_EN_MSB: in     vl_logic_vector(3 downto 0);
        P_PCS_NEAREND_LOOP: in     vl_logic_vector(3 downto 0);
        P_LX_ELECIDLE_EN_0: in     vl_logic_vector(1 downto 0);
        P_LX_ELECIDLE_EN_3: in     vl_logic_vector(1 downto 0);
        P_CIM_CLK_DYN_DLY_SEL_RX: in     vl_logic_vector(3 downto 0);
        P_LX_DEEMP_CTL_3: in     vl_logic_vector(2 downto 0);
        P_LX_ELECIDLE_EN_1: in     vl_logic_vector(1 downto 0);
        P_CIM_CLK_START_ALIGN_TX: in     vl_logic_vector(3 downto 0);
        P_LX_BISTLB_EN  : in     vl_logic_vector(3 downto 0);
        P_TDATA_0       : in     vl_logic_vector(43 downto 0);
        P_CIM_CLK_ALIGNER_RX3: in     vl_logic_vector(7 downto 0);
        P_CIM_CLK_DYN_DLY_SEL_TX: in     vl_logic_vector(3 downto 0);
        P_CIM_CLK_ALIGNER_TX2: in     vl_logic_vector(7 downto 0);
        P_LX_ELECIDLE_EN_2: in     vl_logic_vector(1 downto 0);
        P_RX_LANE_POWERUP: in     vl_logic_vector(3 downto 0);
        P_TX_CKDIV_2    : in     vl_logic_vector(1 downto 0);
        P_PCS_WORD_ALIGN_EN: in     vl_logic_vector(3 downto 0);
        P_LX_AMP_CTL_1  : in     vl_logic_vector(3 downto 0);
        P_CIM_CLK_ALIGNER_RX2: in     vl_logic_vector(7 downto 0);
        P_RX_POLARITY_INVERT: in     vl_logic_vector(3 downto 0);
        P_LX_DEEMP_CTL_2: in     vl_logic_vector(2 downto 0);
        P_LX_AMP_CTL_2  : in     vl_logic_vector(3 downto 0);
        P_LX_RX_CKDIV_1 : in     vl_logic_vector(1 downto 0);
        P_TDATA_3       : in     vl_logic_vector(43 downto 0);
        P_PCS_FAREND_LOOP: in     vl_logic_vector(3 downto 0);
        P_CIM_CLK_START_ALIGN_RX: in     vl_logic_vector(3 downto 0);
        P_LX_RX_CKDIV_0 : in     vl_logic_vector(1 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of PCS_CH0_BYPASS_WORD_ALIGN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_BYPASS_DENC : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_BYPASS_BONDING : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_BYPASS_CTC : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_BYPASS_GEAR : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_BYPASS_BRIDGE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_DATA_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_RX_POLARITY_INV : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_ALIGN_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_SAMP_16B : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_COMMA_REG0 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH0_COMMA_MASK : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH0_CEB_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_CTC_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_A_REG : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH0_GE_AUTO_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_SKIP_REG0 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH0_SKIP_REG1 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH0_SKIP_REG2 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH0_SKIP_REG3 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH0_DEC_DUAL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_SPLIT : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_FIFOFLAG_CTC : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_COMMA_DET_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_ERRDETECT_SILENCE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_PMA_RCLK_POLINV : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_PCS_RCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_MCB_RCLK_POLINV : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_CB_RCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_AFTER_CTC_RCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_RCLK_POLINV : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_BRIDGE_RCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_PCS_RCLK_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_CB_RCLK_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_AFTER_CTC_RCLK_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_AFTER_CTC_RCLK_EN_GB : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_BRIDGE_RCLK_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_PCS_RX_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_SLAVE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_PCIE_SLAVE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_PCS_CB_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_TX_BYPASS_BRIDGE_UINT : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_TX_BYPASS_GEAR : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_TX_BYPASS_ENC : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_TX_BYPASS_BIT_SLIP : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_TX_GEAR_SPLIT : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_TX_DRIVE_REG_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_TX_BIT_SLIP_CYCLES : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH0_INT_TX_MASK_0 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_INT_TX_MASK_1 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_INT_TX_MASK_2 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_INT_TX_CLR_0 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_INT_TX_CLR_1 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_INT_TX_CLR_2 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_TX_PMA_TCLK_POLINV : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_TX_PCS_CLK_EN_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_TX_BRIDGE_TCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_TX_TCLK_POLINV : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_TX_PCS_TX_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_TX_SLAVE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_TX_BRIDGE_CLK_EN_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_DATA_WIDTH_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_TX_TCLK2FABRIC_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_TX_OUTZZ : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_ENC_DUAL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_TX_BITSLIP_DATA_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_COMMA_REG1 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH0_RAPID_IMAX : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH0_RAPID_VMIN_1 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH0_RAPID_VMIN_2 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH0_RX_PRBS_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_RX_ERRCNT_CLR : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_TX_PRBS_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_TX_INSERT_ER : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_ENABLE_PRBS_GEN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_ERR_CNT : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH0_DEFAULT_RADDR : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH0_MASTER_CHECK_OFFSET : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH0_DELAY_SET : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH0_SEACH_OFFSET : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_CEB_RAPIDLS_MMAX : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH0_CTC_AFULL : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH0_CTC_AEMPTY : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH0_FAR_LOOP : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_NEAR_LOOP : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_INT_RX_MASK_0 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_INT_RX_MASK_1 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_INT_RX_MASK_2 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_INT_RX_MASK_3 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_INT_RX_MASK_4 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_INT_RX_MASK_5 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_INT_RX_MASK_6 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_INT_RX_MASK_7 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_INT_RX_CLR_0 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_INT_RX_CLR_1 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_INT_RX_CLR_2 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_INT_RX_CLR_3 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_INT_RX_CLR_4 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_INT_RX_CLR_5 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_INT_RX_CLR_6 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_INT_RX_CLR_7 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_BYPASS_WORD_ALIGN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_BYPASS_DENC : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_BYPASS_BONDING : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_BYPASS_CTC : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_BYPASS_GEAR : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_BYPASS_BRIDGE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_DATA_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_RX_POLARITY_INV : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_ALIGN_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_SAMP_16B : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_COMMA_REG0 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH1_COMMA_MASK : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH1_CEB_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_CTC_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_A_REG : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH1_GE_AUTO_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_SKIP_REG0 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH1_SKIP_REG1 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH1_SKIP_REG2 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH1_SKIP_REG3 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH1_DEC_DUAL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_SPLIT : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_FIFOFLAG_CTC : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_COMMA_DET_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_ERRDETECT_SILENCE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_PMA_RCLK_POLINV : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_PCS_RCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_MCB_RCLK_POLINV : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_CB_RCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_AFTER_CTC_RCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_RCLK_POLINV : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_BRIDGE_RCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_PCS_RCLK_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_CB_RCLK_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_AFTER_CTC_RCLK_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_AFTER_CTC_RCLK_EN_GB : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_BRIDGE_RCLK_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_PCS_RX_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_SLAVE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_PCIE_SLAVE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_PCS_CB_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_TX_BYPASS_BRIDGE_UINT : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_TX_BYPASS_GEAR : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_TX_BYPASS_ENC : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_TX_BYPASS_BIT_SLIP : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_TX_GEAR_SPLIT : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_TX_DRIVE_REG_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_TX_BIT_SLIP_CYCLES : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH1_INT_TX_MASK_0 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_INT_TX_MASK_1 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_INT_TX_MASK_2 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_INT_TX_CLR_0 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_INT_TX_CLR_1 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_INT_TX_CLR_2 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_TX_PMA_TCLK_POLINV : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_TX_PCS_CLK_EN_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_TX_BRIDGE_TCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_TX_TCLK_POLINV : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_TX_PCS_TX_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_TX_SLAVE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_TX_BRIDGE_CLK_EN_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_DATA_WIDTH_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_TX_TCLK2FABRIC_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_TX_OUTZZ : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_ENC_DUAL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_TX_BITSLIP_DATA_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_COMMA_REG1 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH1_RAPID_IMAX : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH1_RAPID_VMIN_1 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH1_RAPID_VMIN_2 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH1_RX_PRBS_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_RX_ERRCNT_CLR : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_TX_PRBS_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_TX_INSERT_ER : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_ENABLE_PRBS_GEN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_ERR_CNT : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH1_DEFAULT_RADDR : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH1_MASTER_CHECK_OFFSET : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH1_DELAY_SET : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH1_SEACH_OFFSET : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_CEB_RAPIDLS_MMAX : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH1_CTC_AFULL : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH1_CTC_AEMPTY : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH1_FAR_LOOP : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_NEAR_LOOP : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_INT_RX_MASK_0 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_INT_RX_MASK_1 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_INT_RX_MASK_2 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_INT_RX_MASK_3 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_INT_RX_MASK_4 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_INT_RX_MASK_5 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_INT_RX_MASK_6 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_INT_RX_MASK_7 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_INT_RX_CLR_0 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_INT_RX_CLR_1 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_INT_RX_CLR_2 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_INT_RX_CLR_3 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_INT_RX_CLR_4 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_INT_RX_CLR_5 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_INT_RX_CLR_6 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_INT_RX_CLR_7 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_BYPASS_WORD_ALIGN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_BYPASS_DENC : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_BYPASS_BONDING : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_BYPASS_CTC : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_BYPASS_GEAR : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_BYPASS_BRIDGE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_DATA_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_RX_POLARITY_INV : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_ALIGN_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_SAMP_16B : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_COMMA_REG0 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH2_COMMA_MASK : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH2_CEB_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_CTC_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_A_REG : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH2_GE_AUTO_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_SKIP_REG0 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH2_SKIP_REG1 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH2_SKIP_REG2 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH2_SKIP_REG3 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH2_DEC_DUAL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_SPLIT : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_FIFOFLAG_CTC : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_COMMA_DET_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_ERRDETECT_SILENCE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_PMA_RCLK_POLINV : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_PCS_RCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_MCB_RCLK_POLINV : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_CB_RCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_AFTER_CTC_RCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_RCLK_POLINV : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_BRIDGE_RCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_PCS_RCLK_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_CB_RCLK_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_AFTER_CTC_RCLK_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_AFTER_CTC_RCLK_EN_GB : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_BRIDGE_RCLK_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_PCS_RX_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_SLAVE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_PCIE_SLAVE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_PCS_CB_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_TX_BYPASS_BRIDGE_UINT : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_TX_BYPASS_GEAR : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_TX_BYPASS_ENC : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_TX_BYPASS_BIT_SLIP : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_TX_GEAR_SPLIT : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_TX_DRIVE_REG_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_TX_BIT_SLIP_CYCLES : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH2_INT_TX_MASK_0 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_INT_TX_MASK_1 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_INT_TX_MASK_2 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_INT_TX_CLR_0 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_INT_TX_CLR_1 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_INT_TX_CLR_2 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_TX_PMA_TCLK_POLINV : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_TX_PCS_CLK_EN_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_TX_BRIDGE_TCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_TX_TCLK_POLINV : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_TX_PCS_TX_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_TX_SLAVE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_TX_BRIDGE_CLK_EN_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_DATA_WIDTH_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_TX_TCLK2FABRIC_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_TX_OUTZZ : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_ENC_DUAL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_TX_BITSLIP_DATA_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_COMMA_REG1 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH2_RAPID_IMAX : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH2_RAPID_VMIN_1 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH2_RAPID_VMIN_2 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH2_RX_PRBS_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_RX_ERRCNT_CLR : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_TX_PRBS_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_TX_INSERT_ER : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_ENABLE_PRBS_GEN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_ERR_CNT : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH2_DEFAULT_RADDR : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH2_MASTER_CHECK_OFFSET : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH2_DELAY_SET : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH2_SEACH_OFFSET : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_CEB_RAPIDLS_MMAX : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH2_CTC_AFULL : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH2_CTC_AEMPTY : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH2_FAR_LOOP : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_NEAR_LOOP : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_INT_RX_MASK_0 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_INT_RX_MASK_1 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_INT_RX_MASK_2 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_INT_RX_MASK_3 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_INT_RX_MASK_4 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_INT_RX_MASK_5 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_INT_RX_MASK_6 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_INT_RX_MASK_7 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_INT_RX_CLR_0 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_INT_RX_CLR_1 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_INT_RX_CLR_2 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_INT_RX_CLR_3 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_INT_RX_CLR_4 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_INT_RX_CLR_5 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_INT_RX_CLR_6 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_INT_RX_CLR_7 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_BYPASS_WORD_ALIGN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_BYPASS_DENC : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_BYPASS_BONDING : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_BYPASS_CTC : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_BYPASS_GEAR : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_BYPASS_BRIDGE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_DATA_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_RX_POLARITY_INV : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_ALIGN_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_SAMP_16B : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_COMMA_REG0 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH3_COMMA_MASK : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH3_CEB_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_CTC_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_A_REG : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH3_GE_AUTO_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_SKIP_REG0 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH3_SKIP_REG1 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH3_SKIP_REG2 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH3_SKIP_REG3 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH3_DEC_DUAL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_SPLIT : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_FIFOFLAG_CTC : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_COMMA_DET_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_ERRDETECT_SILENCE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_PMA_RCLK_POLINV : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_PCS_RCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_MCB_RCLK_POLINV : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_CB_RCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_AFTER_CTC_RCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_RCLK_POLINV : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_BRIDGE_RCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_PCS_RCLK_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_CB_RCLK_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_AFTER_CTC_RCLK_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_AFTER_CTC_RCLK_EN_GB : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_BRIDGE_RCLK_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_PCS_RX_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_SLAVE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_PCIE_SLAVE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_PCS_CB_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_TX_BYPASS_BRIDGE_UINT : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_TX_BYPASS_GEAR : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_TX_BYPASS_ENC : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_TX_BYPASS_BIT_SLIP : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_TX_GEAR_SPLIT : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_TX_DRIVE_REG_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_TX_BIT_SLIP_CYCLES : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH3_INT_TX_MASK_0 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_INT_TX_MASK_1 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_INT_TX_MASK_2 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_INT_TX_CLR_0 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_INT_TX_CLR_1 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_INT_TX_CLR_2 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_TX_PMA_TCLK_POLINV : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_TX_PCS_CLK_EN_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_TX_BRIDGE_TCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_TX_TCLK_POLINV : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_TX_PCS_TX_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_TX_SLAVE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_TX_BRIDGE_CLK_EN_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_DATA_WIDTH_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_TX_TCLK2FABRIC_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_TX_OUTZZ : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_ENC_DUAL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_TX_BITSLIP_DATA_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_COMMA_REG1 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH3_RAPID_IMAX : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH3_RAPID_VMIN_1 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH3_RAPID_VMIN_2 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH3_RX_PRBS_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_RX_ERRCNT_CLR : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_TX_PRBS_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_TX_INSERT_ER : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_ENABLE_PRBS_GEN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_ERR_CNT : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH3_DEFAULT_RADDR : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH3_MASTER_CHECK_OFFSET : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH3_DELAY_SET : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH3_SEACH_OFFSET : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_CEB_RAPIDLS_MMAX : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH3_CTC_AFULL : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH3_CTC_AEMPTY : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH3_FAR_LOOP : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_NEAR_LOOP : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_INT_RX_MASK_0 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_INT_RX_MASK_1 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_INT_RX_MASK_2 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_INT_RX_MASK_3 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_INT_RX_MASK_4 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_INT_RX_MASK_5 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_INT_RX_MASK_6 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_INT_RX_MASK_7 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_INT_RX_CLR_0 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_INT_RX_CLR_1 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_INT_RX_CLR_2 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_INT_RX_CLR_3 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_INT_RX_CLR_4 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_INT_RX_CLR_5 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_INT_RX_CLR_6 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_INT_RX_CLR_7 : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_TXDATA_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_TX_TESTPATTERN : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_TESTPATTERN_O_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_DISABLE_BSMODE_DRVAMP : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_FORCE_BIST_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_FORCE_ELECTRICAL_IDLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_FORCE_RXDCT_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_FORCE_EXTLB_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_DISABLE_LANE_SYNC : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_DISABLE_ELECTRICAL_IDLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_DISABLE_RXDCT_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_DISABLE_EXTLB_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_DISABLE_LOW_SPEED_PATH_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_FORCE_LANE_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_FORCE_LANE_RESETB_DISABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_RXDCT_LGBW_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_RXDCT_VTH : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_DE_EMPHASIS_ADDITIONAL_CONTROL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_DRV_RTERM_CONTROL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_FDRV_AMP_CONTROL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_PREPC_AMP_CONTROL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_PREMC_AMP_CONTROL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_SER_AMP_CONTROL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_PFD_LOOP_RESISTOR_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_PD_LOOP_RESISTOR_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_CDR_TEST_OUT_SELECT : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_PI_DIV1_BP : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_PI_TEST_FOR_CKI : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_PI_CURRENT_SETTING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_PI_FREQUENCY_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_TEST_OUT_SELECT_FOR_RCK : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_TEST_OUT_SELECT_SOURCE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_TEST_DATA_OUT_SELECT_SOURCE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_TEST_CK_OUT_SELECT_SOURCE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_ENABLE_SLIP1UI_MODULE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_PN_SWAP_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_SIPO_BIT_SETTING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_OOB_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_ALOS_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_LFMODE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_TSO_HS_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_LX_SELLC : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_LX_RXPLL_DIVSEL45_FB : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_LX_RXPLL_DIVSEL_FB : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_LX_RXPLL_DIVSEL_REF : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_PICODE : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_RX_REFCK_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_PFDLPEN_REGISTER_CONTROL_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_PFDLPEN_REGISTER_SETTING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_PDLPEN_REGISTER_CONTROL_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_PDLPEN_REGISTER_SETTING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_DIV_CHANGE_ENABLE_DELAY_TIMER : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_DIV_CHANGE_ENABLE_SIGNAL_GATING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_CDR_ALIGN_REGISTER_SETTING_VALUE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_FORCE_CDR_ALIGN_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_SELLC_REGISTER_SETTING_VALUE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_SELLC_CONTROL_BY_REGISTER : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_PLLI_LDO_VREF_SETTING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_PLLI_LDO_BYPASS_CURRENT : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_PLL_HSTEST_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_PLL_ISNK_CURRENT_CONTROL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_PLL_PFD_LOOP_CP0_CURRENT_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_PLL_PD_LOOP_PLLGM_SETTING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_PLL_PFD_LOOP_CP1_CURRENT_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_PLL_CP0_BIAS_CONTROL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_PLL_PD_LOOP_CP0_CURRENT_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_PLL_CP1_BIAS_CONTROL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_PLL_PD_LOOP_CP1_CURRENT_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_PLL_CP0_CURRENT_SETTING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_PLL_CP1_CURRENT_SETTING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_PLL_GM1_CURRENT_SETTING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_PLL_LC_BF2_CURRENT_SETTING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_PLL_LC_BF2_CURRENT_SETTING_LOW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_PLL_REG_CUR : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_PLL_LCCUR : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_PLL_LCOBAS : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_PLL_FB_CK_TEST_OUT_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_CDR_ALIGN_TIMER : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_CALIB_WAIT : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_CALIB_TIMER : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_TOT_RANGE : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_SUB_RANGE : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_OVLP : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_BIST_WAIT : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_BIST_TIMER : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_BAND_LB : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_BAND_HB : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_FREQ_LOCK_ACCURACY : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_SET_LC_BAND : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_SET_VCODIV : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REGISTER_SET_VCODIV_BAND_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_SET_PLL_LOCK : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REGISTER_SET_PLL_LOCK_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_SET_VCO_HI : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_SET_VCO_LO : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REGISTER_SET_VCO_HI_VCO_LO_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_FORCE_LC_PLL_LOOP_EN_H : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_FORCE_LC_PLL_LOOP_EN_L : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_VCO_DIV_CALI_BYPASS : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_BIST_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_PLL_LOOP_EN_SETTING_FROM_REGISTER_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_FREQ_DETECT_ENABLE_SOURCE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_SET_DIVSEL_REF : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_SET_DIVSEL45_FB : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_SET_DIVSEL_FB : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_PLL_LOOP_EN_SETTING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REGISTER_SET_TXPLL_DIV_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_FORCE_RXPLL_RESET : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_FORCE_RXPLL_ON : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_DPCK_DIV2 : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_LFO_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_ALOS_COUNTER_CLOCK_SELECTION : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_RX_BIAS_CURRENT_ADJUSTMENT : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_OOB_ENTER_DELAY_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_ALOS_LOW_TO_HIGH_COUNTER_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_ENABLE_ALOS_RESULT_AUTOMATICALLY_ENABLE_CHANNEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_ALOS_EXIT_COUNTER_CLOCK_DIVIDER : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_OOB_OSCILATER_FREQUENCY_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_FORCE_OOB : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_OOB_VTH_SET : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_FORCE_DET_FORCE_ALOS_LOW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_ALOS_THRESHOLD_VOLTAGE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_WAKEUP_VCM_RX_COMMON_MODE_VOLTAGE : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REGR_NEGATIVE_HYSTERESIS_SETTING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REGL_POSITIVE_HYSTERESIS_SETTING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REGREF_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_DC496 : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_EQ2_AC_VAR_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_EQ2_AC_RES_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_EQ2_DC_RESTOP_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_EQ1_DC_RESTOP_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_EQ1_AC_VAR_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_EQ2_CURRENT_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_EQ1_AC_RES_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_EQ1_CURRENT_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_RPLUS : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_RMINUS : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_RVALSET : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_RTERM : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_DCFB_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_DCCOUP : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_3G : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_TXDATA_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_TX_TESTPATTERN : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_TESTPATTERN_O_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_DISABLE_BSMODE_DRVAMP : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_FORCE_BIST_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_FORCE_ELECTRICAL_IDLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_FORCE_RXDCT_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_FORCE_EXTLB_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_DISABLE_LANE_SYNC : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_DISABLE_ELECTRICAL_IDLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_DISABLE_RXDCT_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_DISABLE_EXTLB_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_DISABLE_LOW_SPEED_PATH_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_FORCE_LANE_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_FORCE_LANE_RESETB_DISABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_RXDCT_LGBW_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_RXDCT_VTH : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_DE_EMPHASIS_ADDITIONAL_CONTROL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_DRV_RTERM_CONTROL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_FDRV_AMP_CONTROL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_PREPC_AMP_CONTROL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_PREMC_AMP_CONTROL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_SER_AMP_CONTROL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_PFD_LOOP_RESISTOR_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_PD_LOOP_RESISTOR_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_CDR_TEST_OUT_SELECT : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_PI_DIV1_BP : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_PI_TEST_FOR_CKI : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_PI_CURRENT_SETTING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_PI_FREQUENCY_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_TEST_OUT_SELECT_FOR_RCK : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_TEST_OUT_SELECT_SOURCE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_TEST_DATA_OUT_SELECT_SOURCE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_TEST_CK_OUT_SELECT_SOURCE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_ENABLE_SLIP1UI_MODULE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_PN_SWAP_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_SIPO_BIT_SETTING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_OOB_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_ALOS_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_LFMODE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_TSO_HS_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_LX_SELLC : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_LX_RXPLL_DIVSEL45_FB : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_LX_RXPLL_DIVSEL_FB : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_LX_RXPLL_DIVSEL_REF : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_PICODE : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_RX_REFCK_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_PFDLPEN_REGISTER_CONTROL_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_PFDLPEN_REGISTER_SETTING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_PDLPEN_REGISTER_CONTROL_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_PDLPEN_REGISTER_SETTING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_DIV_CHANGE_ENABLE_DELAY_TIMER : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_DIV_CHANGE_ENABLE_SIGNAL_GATING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_CDR_ALIGN_REGISTER_SETTING_VALUE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_FORCE_CDR_ALIGN_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_SELLC_REGISTER_SETTING_VALUE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_SELLC_CONTROL_BY_REGISTER : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_PLLI_LDO_VREF_SETTING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_PLLI_LDO_BYPASS_CURRENT : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_PLL_HSTEST_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_PLL_ISNK_CURRENT_CONTROL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_PLL_PFD_LOOP_CP0_CURRENT_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_PLL_PD_LOOP_PLLGM_SETTING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_PLL_PFD_LOOP_CP1_CURRENT_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_PLL_CP0_BIAS_CONTROL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_PLL_PD_LOOP_CP0_CURRENT_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_PLL_CP1_BIAS_CONTROL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_PLL_PD_LOOP_CP1_CURRENT_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_PLL_CP0_CURRENT_SETTING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_PLL_CP1_CURRENT_SETTING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_PLL_GM1_CURRENT_SETTING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_PLL_LC_BF2_CURRENT_SETTING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_PLL_LC_BF2_CURRENT_SETTING_LOW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_PLL_REG_CUR : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_PLL_LCCUR : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_PLL_LCOBAS : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_PLL_FB_CK_TEST_OUT_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_CDR_ALIGN_TIMER : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_CALIB_WAIT : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_CALIB_TIMER : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_TOT_RANGE : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_SUB_RANGE : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_OVLP : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_BIST_WAIT : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_BIST_TIMER : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_BAND_LB : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_BAND_HB : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_FREQ_LOCK_ACCURACY : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_SET_LC_BAND : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_SET_VCODIV : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REGISTER_SET_VCODIV_BAND_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_SET_PLL_LOCK : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REGISTER_SET_PLL_LOCK_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_SET_VCO_HI : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_SET_VCO_LO : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REGISTER_SET_VCO_HI_VCO_LO_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_FORCE_LC_PLL_LOOP_EN_H : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_FORCE_LC_PLL_LOOP_EN_L : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_VCO_DIV_CALI_BYPASS : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_BIST_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_PLL_LOOP_EN_SETTING_FROM_REGISTER_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_FREQ_DETECT_ENABLE_SOURCE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_SET_DIVSEL_REF : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_SET_DIVSEL45_FB : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_SET_DIVSEL_FB : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_PLL_LOOP_EN_SETTING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REGISTER_SET_TXPLL_DIV_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_FORCE_RXPLL_RESET : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_FORCE_RXPLL_ON : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_DPCK_DIV2 : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_LFO_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_ALOS_COUNTER_CLOCK_SELECTION : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_RX_BIAS_CURRENT_ADJUSTMENT : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_OOB_ENTER_DELAY_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_ALOS_LOW_TO_HIGH_COUNTER_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_ENABLE_ALOS_RESULT_AUTOMATICALLY_ENABLE_CHANNEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_ALOS_EXIT_COUNTER_CLOCK_DIVIDER : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_OOB_OSCILATER_FREQUENCY_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_FORCE_OOB : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_OOB_VTH_SET : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_FORCE_DET_FORCE_ALOS_LOW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_ALOS_THRESHOLD_VOLTAGE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_WAKEUP_VCM_RX_COMMON_MODE_VOLTAGE : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REGR_NEGATIVE_HYSTERESIS_SETTING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REGL_POSITIVE_HYSTERESIS_SETTING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REGREF_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_DC496 : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_EQ2_AC_VAR_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_EQ2_AC_RES_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_EQ2_DC_RESTOP_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_EQ1_DC_RESTOP_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_EQ1_AC_VAR_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_EQ2_CURRENT_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_EQ1_AC_RES_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_EQ1_CURRENT_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_RPLUS : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_RMINUS : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_RVALSET : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_RTERM : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_DCFB_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_DCCOUP : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_3G : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_TXDATA_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_TX_TESTPATTERN : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_TESTPATTERN_O_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_DISABLE_BSMODE_DRVAMP : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_FORCE_BIST_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_FORCE_ELECTRICAL_IDLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_FORCE_RXDCT_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_FORCE_EXTLB_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_DISABLE_LANE_SYNC : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_DISABLE_ELECTRICAL_IDLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_DISABLE_RXDCT_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_DISABLE_EXTLB_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_DISABLE_LOW_SPEED_PATH_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_FORCE_LANE_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_FORCE_LANE_RESETB_DISABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_RXDCT_LGBW_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_RXDCT_VTH : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_DE_EMPHASIS_ADDITIONAL_CONTROL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_DRV_RTERM_CONTROL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_FDRV_AMP_CONTROL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_PREPC_AMP_CONTROL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_PREMC_AMP_CONTROL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_SER_AMP_CONTROL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_PFD_LOOP_RESISTOR_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_PD_LOOP_RESISTOR_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_CDR_TEST_OUT_SELECT : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_PI_DIV1_BP : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_PI_TEST_FOR_CKI : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_PI_CURRENT_SETTING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_PI_FREQUENCY_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_TEST_OUT_SELECT_FOR_RCK : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_TEST_OUT_SELECT_SOURCE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_TEST_DATA_OUT_SELECT_SOURCE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_TEST_CK_OUT_SELECT_SOURCE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_ENABLE_SLIP1UI_MODULE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_PN_SWAP_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_SIPO_BIT_SETTING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_OOB_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_ALOS_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_LFMODE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_TSO_HS_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_LX_SELLC : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_LX_RXPLL_DIVSEL45_FB : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_LX_RXPLL_DIVSEL_FB : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_LX_RXPLL_DIVSEL_REF : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_PICODE : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_RX_REFCK_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_PFDLPEN_REGISTER_CONTROL_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_PFDLPEN_REGISTER_SETTING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_PDLPEN_REGISTER_CONTROL_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_PDLPEN_REGISTER_SETTING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_DIV_CHANGE_ENABLE_DELAY_TIMER : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_DIV_CHANGE_ENABLE_SIGNAL_GATING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_CDR_ALIGN_REGISTER_SETTING_VALUE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_FORCE_CDR_ALIGN_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_SELLC_REGISTER_SETTING_VALUE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_SELLC_CONTROL_BY_REGISTER : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_PLLI_LDO_VREF_SETTING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_PLLI_LDO_BYPASS_CURRENT : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_PLL_HSTEST_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_PLL_ISNK_CURRENT_CONTROL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_PLL_PFD_LOOP_CP0_CURRENT_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_PLL_PD_LOOP_PLLGM_SETTING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_PLL_PFD_LOOP_CP1_CURRENT_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_PLL_CP0_BIAS_CONTROL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_PLL_PD_LOOP_CP0_CURRENT_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_PLL_CP1_BIAS_CONTROL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_PLL_PD_LOOP_CP1_CURRENT_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_PLL_CP0_CURRENT_SETTING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_PLL_CP1_CURRENT_SETTING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_PLL_GM1_CURRENT_SETTING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_PLL_LC_BF2_CURRENT_SETTING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_PLL_LC_BF2_CURRENT_SETTING_LOW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_PLL_REG_CUR : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_PLL_LCCUR : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_PLL_LCOBAS : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_PLL_FB_CK_TEST_OUT_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_CDR_ALIGN_TIMER : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_CALIB_WAIT : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_CALIB_TIMER : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_TOT_RANGE : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_SUB_RANGE : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_OVLP : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_BIST_WAIT : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_BIST_TIMER : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_BAND_LB : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_BAND_HB : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_FREQ_LOCK_ACCURACY : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_SET_LC_BAND : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_SET_VCODIV : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REGISTER_SET_VCODIV_BAND_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_SET_PLL_LOCK : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REGISTER_SET_PLL_LOCK_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_SET_VCO_HI : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_SET_VCO_LO : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REGISTER_SET_VCO_HI_VCO_LO_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_FORCE_LC_PLL_LOOP_EN_H : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_FORCE_LC_PLL_LOOP_EN_L : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_VCO_DIV_CALI_BYPASS : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_BIST_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_PLL_LOOP_EN_SETTING_FROM_REGISTER_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_FREQ_DETECT_ENABLE_SOURCE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_SET_DIVSEL_REF : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_SET_DIVSEL45_FB : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_SET_DIVSEL_FB : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_PLL_LOOP_EN_SETTING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REGISTER_SET_TXPLL_DIV_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_FORCE_RXPLL_RESET : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_FORCE_RXPLL_ON : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_DPCK_DIV2 : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_LFO_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_ALOS_COUNTER_CLOCK_SELECTION : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_RX_BIAS_CURRENT_ADJUSTMENT : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_OOB_ENTER_DELAY_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_ALOS_LOW_TO_HIGH_COUNTER_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_ENABLE_ALOS_RESULT_AUTOMATICALLY_ENABLE_CHANNEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_ALOS_EXIT_COUNTER_CLOCK_DIVIDER : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_OOB_OSCILATER_FREQUENCY_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_FORCE_OOB : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_OOB_VTH_SET : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_FORCE_DET_FORCE_ALOS_LOW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_ALOS_THRESHOLD_VOLTAGE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_WAKEUP_VCM_RX_COMMON_MODE_VOLTAGE : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REGR_NEGATIVE_HYSTERESIS_SETTING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REGL_POSITIVE_HYSTERESIS_SETTING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REGREF_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_DC496 : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_EQ2_AC_VAR_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_EQ2_AC_RES_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_EQ2_DC_RESTOP_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_EQ1_DC_RESTOP_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_EQ1_AC_VAR_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_EQ2_CURRENT_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_EQ1_AC_RES_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_EQ1_CURRENT_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_RPLUS : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_RMINUS : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_RVALSET : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_RTERM : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_DCFB_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_DCCOUP : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_3G : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_TXDATA_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_TX_TESTPATTERN : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_TESTPATTERN_O_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_DISABLE_BSMODE_DRVAMP : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_FORCE_BIST_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_FORCE_ELECTRICAL_IDLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_FORCE_RXDCT_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_FORCE_EXTLB_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_DISABLE_LANE_SYNC : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_DISABLE_ELECTRICAL_IDLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_DISABLE_RXDCT_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_DISABLE_EXTLB_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_DISABLE_LOW_SPEED_PATH_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_FORCE_LANE_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_FORCE_LANE_RESETB_DISABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_RXDCT_LGBW_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_RXDCT_VTH : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_DE_EMPHASIS_ADDITIONAL_CONTROL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_DRV_RTERM_CONTROL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_FDRV_AMP_CONTROL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_PREPC_AMP_CONTROL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_PREMC_AMP_CONTROL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_SER_AMP_CONTROL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_PFD_LOOP_RESISTOR_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_PD_LOOP_RESISTOR_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_CDR_TEST_OUT_SELECT : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_PI_DIV1_BP : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_PI_TEST_FOR_CKI : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_PI_CURRENT_SETTING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_PI_FREQUENCY_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_TEST_OUT_SELECT_FOR_RCK : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_TEST_OUT_SELECT_SOURCE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_TEST_DATA_OUT_SELECT_SOURCE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_TEST_CK_OUT_SELECT_SOURCE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_ENABLE_SLIP1UI_MODULE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_PN_SWAP_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_SIPO_BIT_SETTING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_OOB_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_ALOS_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_LFMODE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_TSO_HS_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_LX_SELLC : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_LX_RXPLL_DIVSEL45_FB : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_LX_RXPLL_DIVSEL_FB : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_LX_RXPLL_DIVSEL_REF : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_PICODE : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_RX_REFCK_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_PFDLPEN_REGISTER_CONTROL_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_PFDLPEN_REGISTER_SETTING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_PDLPEN_REGISTER_CONTROL_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_PDLPEN_REGISTER_SETTING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_DIV_CHANGE_ENABLE_DELAY_TIMER : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_DIV_CHANGE_ENABLE_SIGNAL_GATING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_CDR_ALIGN_REGISTER_SETTING_VALUE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_FORCE_CDR_ALIGN_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_SELLC_REGISTER_SETTING_VALUE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_SELLC_CONTROL_BY_REGISTER : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_PLLI_LDO_VREF_SETTING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_PLLI_LDO_BYPASS_CURRENT : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_PLL_HSTEST_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_PLL_ISNK_CURRENT_CONTROL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_PLL_PFD_LOOP_CP0_CURRENT_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_PLL_PD_LOOP_PLLGM_SETTING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_PLL_PFD_LOOP_CP1_CURRENT_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_PLL_CP0_BIAS_CONTROL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_PLL_PD_LOOP_CP0_CURRENT_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_PLL_CP1_BIAS_CONTROL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_PLL_PD_LOOP_CP1_CURRENT_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_PLL_CP0_CURRENT_SETTING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_PLL_CP1_CURRENT_SETTING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_PLL_GM1_CURRENT_SETTING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_PLL_LC_BF2_CURRENT_SETTING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_PLL_LC_BF2_CURRENT_SETTING_LOW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_PLL_REG_CUR : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_PLL_LCCUR : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_PLL_LCOBAS : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_PLL_FB_CK_TEST_OUT_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_CDR_ALIGN_TIMER : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_CALIB_WAIT : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_CALIB_TIMER : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_TOT_RANGE : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_SUB_RANGE : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_OVLP : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_BIST_WAIT : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_BIST_TIMER : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_BAND_LB : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_BAND_HB : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_FREQ_LOCK_ACCURACY : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_SET_LC_BAND : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_SET_VCODIV : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REGISTER_SET_VCODIV_BAND_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_SET_PLL_LOCK : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REGISTER_SET_PLL_LOCK_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_SET_VCO_HI : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_SET_VCO_LO : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REGISTER_SET_VCO_HI_VCO_LO_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_FORCE_LC_PLL_LOOP_EN_H : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_FORCE_LC_PLL_LOOP_EN_L : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_VCO_DIV_CALI_BYPASS : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_BIST_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_PLL_LOOP_EN_SETTING_FROM_REGISTER_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_FREQ_DETECT_ENABLE_SOURCE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_SET_DIVSEL_REF : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_SET_DIVSEL45_FB : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_SET_DIVSEL_FB : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_PLL_LOOP_EN_SETTING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REGISTER_SET_TXPLL_DIV_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_FORCE_RXPLL_RESET : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_FORCE_RXPLL_ON : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_DPCK_DIV2 : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_LFO_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_ALOS_COUNTER_CLOCK_SELECTION : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_RX_BIAS_CURRENT_ADJUSTMENT : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_OOB_ENTER_DELAY_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_ALOS_LOW_TO_HIGH_COUNTER_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_ENABLE_ALOS_RESULT_AUTOMATICALLY_ENABLE_CHANNEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_ALOS_EXIT_COUNTER_CLOCK_DIVIDER : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_OOB_OSCILATER_FREQUENCY_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_FORCE_OOB : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_OOB_VTH_SET : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_FORCE_DET_FORCE_ALOS_LOW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_ALOS_THRESHOLD_VOLTAGE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_WAKEUP_VCM_RX_COMMON_MODE_VOLTAGE : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REGR_NEGATIVE_HYSTERESIS_SETTING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REGL_POSITIVE_HYSTERESIS_SETTING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REGREF_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_DC496 : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_EQ2_AC_VAR_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_EQ2_AC_RES_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_EQ2_DC_RESTOP_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_EQ1_DC_RESTOP_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_EQ1_AC_VAR_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_EQ2_CURRENT_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_EQ1_AC_RES_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_EQ1_CURRENT_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_RPLUS : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_RMINUS : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_RVALSET : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_RTERM : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_DCFB_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_DCCOUP : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_3G : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_TURN_ON_BANDGAP_AT_AOS_ON : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_TURN_ON_BANDGAP_AT_RX_DETECTION_ON : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_TURN_ON_BANDGAP_AT_BOUNDARY_SCAN_ON : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_CFG_HSST_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_SELECT_LANE_TCK_FOR_QUAD_SYNC : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_CK_REN : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_C1_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_C2_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_CLK_DIVIDER_SETTING_FROM_25M_TO_200K : constant is 2;
    attribute mti_svvh_generic_type of PMA_QUAD_ACMODE_SCANMODE_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_REGISTER_ACMODE : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_REGISTER_SCANMODE : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_REFCK2CORE_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_REG_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_REGR : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_REGL : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_DPCK_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_QUAD_TX_REFCK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_REFCK_SRC_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_RREFCK_PWRUP : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_REFCK_SK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_REFCK_DIV2_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_REFCK_TO_NQ_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_AUXI_ADJ : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_DC496 : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_REG_FDET_TIMER : constant is 2;
    attribute mti_svvh_generic_type of PMA_QUAD_FREQ_LKO : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_FREQ_LKI : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_CLOCK_SRC_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_FRE_DET_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_TSO_LS_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_QUAD_TXPLL_START : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_VCODIV : constant is 2;
    attribute mti_svvh_generic_type of PMA_QUAD_LC_BAND : constant is 2;
    attribute mti_svvh_generic_type of PMA_QUAD_SET_VCO_HI : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_SET_VCO_LO : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_CALIB_FAIL : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_CALIB_DONE : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_BIST_DONE : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_TOTRANGE_FAIL : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_SUBRANGE_FAIL : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_OVLP_FAIL : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_TXPLL_LOCK : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_TXPLL_LOOP_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_TXPLL_DIVSEL_REF_STA : constant is 2;
    attribute mti_svvh_generic_type of PMA_QUAD_TXPLL_DIVSEL45_FB_STA : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_TXPLL_DIVSEL_FB_STA : constant is 2;
    attribute mti_svvh_generic_type of PMA_QUAD_TXPLL_DIVSEL45_FB : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_TXPLL_DIVSEL_FB : constant is 2;
    attribute mti_svvh_generic_type of PMA_QUAD_TXPLL_DIVSEL_REF : constant is 2;
    attribute mti_svvh_generic_type of PMA_QUAD_REG_DISABLE_HOLDCLK : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_REG_DISABLE_SYNC : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_FORCE_OUTPUT_PLL_LOCK : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_REGISTER_SET_SYNCTCK_SEL_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_REG_SET_SYNCTCK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_CK4TEST_OUTPUT_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_RSTGENBAS : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_LCBUFBAS : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_REGISTER_SET_CPCUR_ENABEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_REG_SET_CPCUR : constant is 2;
    attribute mti_svvh_generic_type of PMA_QUAD_CPBAS : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_LCOBAS : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_LCCUR : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_ENABLE_REGISTER_SETTING_BAND : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_CALIB_WAIT : constant is 2;
    attribute mti_svvh_generic_type of PMA_QUAD_CALIB_TIMER : constant is 2;
    attribute mti_svvh_generic_type of PMA_QUAD_TOT_RANGE : constant is 2;
    attribute mti_svvh_generic_type of PMA_QUAD_SUB_RANGE : constant is 2;
    attribute mti_svvh_generic_type of PMA_QUAD_OVLP : constant is 2;
    attribute mti_svvh_generic_type of PMA_QUAD_BIST_WAIT : constant is 2;
    attribute mti_svvh_generic_type of PMA_QUAD_BIST_TIMER : constant is 2;
    attribute mti_svvh_generic_type of PMA_QUAD_BAND_LB : constant is 2;
    attribute mti_svvh_generic_type of PMA_QUAD_BAND_HB : constant is 2;
    attribute mti_svvh_generic_type of PMA_QUAD_FREQ_LOCK_ACCURACY : constant is 2;
    attribute mti_svvh_generic_type of PMA_QUAD_REG_SET_LC_BAND : constant is 2;
    attribute mti_svvh_generic_type of PMA_QUAD_REG_SET_VCODIV : constant is 2;
    attribute mti_svvh_generic_type of PMA_QUAD_REGISTER_SET_VCODIV_BAND_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_REG_SET_PLL_LOCK : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_REGISTER_SET_PLL_LOCK_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_REG_SET_VCO_HI : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_REG_SET_VCO_LO : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_REGISTER_SET_VCO_HI_VCO_LO_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_FORCE_LC_PLL_LOOP_EN_H : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_FORCE_LC_PLL_LOOP_EN_L : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_VCO_DIV_CALI_BYPASS : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_BIST_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_ENABLE_TXPLL_BIST_BLOCK_CLOCKS : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_LF_TESTBY2 : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_REG_SET_DIVSEL_REF : constant is 2;
    attribute mti_svvh_generic_type of PMA_QUAD_REG_SET_DIVSEL45_FB : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_REG_SET_DIVSEL_FB : constant is 2;
    attribute mti_svvh_generic_type of PMA_QUAD_LF_TEST_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_REGISTER_SET_TXPLL_DIV_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_FORCE_TXPLL_RESET : constant is 1;
    attribute mti_svvh_generic_type of PMA_QUAD_FORCE_TXPLL_ON : constant is 1;
    attribute mti_svvh_generic_type of CLK_ALIGNER_RX0 : constant is 2;
    attribute mti_svvh_generic_type of CLK_ALIGNER_RX1 : constant is 2;
    attribute mti_svvh_generic_type of CLK_ALIGNER_RX2 : constant is 2;
    attribute mti_svvh_generic_type of CLK_ALIGNER_RX3 : constant is 2;
    attribute mti_svvh_generic_type of CLK_ALIGNER_TX0 : constant is 2;
    attribute mti_svvh_generic_type of CLK_ALIGNER_TX1 : constant is 2;
    attribute mti_svvh_generic_type of CLK_ALIGNER_TX2 : constant is 2;
    attribute mti_svvh_generic_type of CLK_ALIGNER_TX3 : constant is 2;
    attribute mti_svvh_generic_type of DYN_DLY_EN_RX0 : constant is 1;
    attribute mti_svvh_generic_type of DYN_DLY_EN_RX1 : constant is 1;
    attribute mti_svvh_generic_type of DYN_DLY_EN_RX2 : constant is 1;
    attribute mti_svvh_generic_type of DYN_DLY_EN_RX3 : constant is 1;
    attribute mti_svvh_generic_type of DYN_DLY_EN_TX0 : constant is 1;
    attribute mti_svvh_generic_type of DYN_DLY_EN_TX1 : constant is 1;
    attribute mti_svvh_generic_type of DYN_DLY_EN_TX2 : constant is 1;
    attribute mti_svvh_generic_type of DYN_DLY_EN_TX3 : constant is 1;
    attribute mti_svvh_generic_type of DYN_DLY_SEL_RX0 : constant is 1;
    attribute mti_svvh_generic_type of DYN_DLY_SEL_RX1 : constant is 1;
    attribute mti_svvh_generic_type of DYN_DLY_SEL_RX2 : constant is 1;
    attribute mti_svvh_generic_type of DYN_DLY_SEL_RX3 : constant is 1;
    attribute mti_svvh_generic_type of DYN_DLY_SEL_TX0 : constant is 1;
    attribute mti_svvh_generic_type of DYN_DLY_SEL_TX1 : constant is 1;
    attribute mti_svvh_generic_type of DYN_DLY_SEL_TX2 : constant is 1;
    attribute mti_svvh_generic_type of DYN_DLY_SEL_TX3 : constant is 1;
    attribute mti_svvh_generic_type of CLK_ALIGNER_RSTN_RX : constant is 2;
    attribute mti_svvh_generic_type of CLK_ALIGNER_RSTN_TX : constant is 2;
    attribute mti_svvh_generic_type of LX_BISTLB_EN : constant is 2;
    attribute mti_svvh_generic_type of LX_ELECIDLE_EN_MSB : constant is 2;
    attribute mti_svvh_generic_type of LX_EXTLB_EN : constant is 2;
    attribute mti_svvh_generic_type of LX_RXDCT_EN : constant is 2;
    attribute mti_svvh_generic_type of LX_TX_LFMODE : constant is 2;
    attribute mti_svvh_generic_type of RX_LANE_POWERUP : constant is 2;
    attribute mti_svvh_generic_type of TX_LANE_POWERUP : constant is 2;
    attribute mti_svvh_generic_type of PLL_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PLLPOWERDOWN : constant is 1;
    attribute mti_svvh_generic_type of QUAD_PWRUP : constant is 1;
    attribute mti_svvh_generic_type of GRSN_DIS : constant is 1;
    attribute mti_svvh_generic_type of HSST_RSTN : constant is 1;
    attribute mti_svvh_generic_type of CFG_RSTN : constant is 1;
end GTP_HSST;
