`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R07bEjRs0CGYhJECabkGGr0DAlfvCmvg5eDW8GjOtZlL8jssQ4YyZby0CFViYJE6
fiaEjEVjpBshZ9ulD26k9688hyfpbtpMAIJzOhwQo0RtgyjBLeiBD0PdyGlU+pv5
3IwiQyoRaN3Akeg7eJcxriJEyZE4BwKoKjBdxqJ7mpaAzhOGCbSvoCnaJGqViJoA
JvMlHTMgEQMwg5GouYqJmHX6uYJ2ccxNJPcn5wOxOogsrQe/g3DTTQS+roGUT5H8
x+jX9hEOf0PjwED5bMAh6iZla8N+DXjtWg7YA64vWhVGaqXh7ZWpqOcW+Bs7huYx
cLisCoJuokKtUA/p0qx+ObN1hurfCjR0scaKyhS0lTJQ9EjO/FlvHwsVLmY/VKXT
sbxG5OEsNlrr0ECnQkqwWwAGPBOEl68Nl+bZ9JSF0aP81MIpJ3HzQjSBT5Q92X8d
+lUG0j9b6iUD1nS7koBGZV0XsGK2rQak14DoJtcRkvzSf0vZyQjebyeCzhbuy3ue
XLIEnIo+uVBV8c3ewYv7TR7ZOY+qIsq+MYHXP0VukaMeV3byAX7IPo9g8SNiQpeN
b9A1uo5UA6YHO2L/0ZlsyBESZvxkHb9spKQJDXP75OSpW/bkQpcwnrjXv3lFo5jp
OyyqfYONVlXADaj0hepa7QvLoxp6i10N52hmQ/TaeWCsl2oJ53wrbHQEMAzfpf2s
Ll24S9MUcAMrKz93WUhTEUCdkIKn/vIABwmxCNYLHo7rZeNB23GBr4Bnpm967rjS
Ae5ow2eCIxrwIHPTb94d3sgZSSSlSNoU9XiJyLSiLQ1w1rgbEj3enNGGW+iXCaXR
wQ8SvIhCDGGBU1ewojfW/GGsv/oBmyQNk0Hs5HtunlyXGiGuqDscVx1XNiIMcQ9C
OaVUjmJ5v43X9Kmc2LWM8rXcKHBicOg1iSdwMr1+WU7myLgVbuNdOSCcjuFev7Ar
us8KkwoYIkvSEMWktJB5qGThehsrl5qG5vX7Qjpr4h3RDS+BNTa9SOciVQ/PtAtM
m9OYBPo2Oef7Ntt5V4fh+LA1j3LTC42wXHLarkG1FuEJ35tIiSaUZROHGvTIeOhD
Rj/2hf3+sMr3IlkBDKIMlCVZ7LtmCF2hdS+w7RKkELH+5KQ+JV5zHzjxxOHxp0Bq
AJiBqVbSa9+0cQPDnJ2Bo5B71A+3ilzPvFUVYIx/ZZlvFIdixe/1RWxh1Adi3M1T
zYNGY3K7pf+G/tFXSjNSiIuGDMoJHt4ifpmk7boMrDv2NLunB7J8c3f+GWN3mlfd
`protect END_PROTECTED
