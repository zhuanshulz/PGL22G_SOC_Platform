`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k6IyodTQ83guhpidrEzo2r+HdLbkFiEuWI54UdWotQNVvtuv4M3ZmOzTMafuz+gN
YY7Du2lLyf+T/FxCVnf8x3+M1oa+GfWdkeLpwt/R5zY4LZ5cLJteC3gNQttYn5/0
FE/1EGgRjuJpVj8FTio3a7AQLgkMU0auUhP8+u+I+I3TTcbGOlVRMSBXwQ/Q/SfG
Btd8a0Frfdd4vejAD/WBYxi5pNb1771MxZA4miGLOcjFJsW2l0ZmmQ3eAs1bkpTC
WvAFHL+ANK71hcX8KquQglDcrxKeExMXHsX4Zb5LGs5PXoIk7ZK97kCYHX9wWXyz
4RbNb0TwZn4rdIwvqCe1byeeD3X0PIIQ3BXGcZcpwa0=
`protect END_PROTECTED
