`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
64+xXtz1oOv+eXdkp24WxRyiXzJa+P3qR4rmtTJ+nF1qniK1TQ1Z3ALeNZma2jHU
f5xAJYDPOaszhW8R+UA5iqKhIrE5EyG/jae4UHExqNxDSPoUnB8h+vdF4LEMC5FO
pUyLCYwgCyskoWUY93D+ijsBEBdtkRoPcG0VfpYGKsgaKEhrwto2OD1XW9ZcnFv/
rPtJCHoILWDymubneTjwmLQ7KmW5ucovbdQplHu5brnIOefJPPEz2ExqRJS5K2Yk
SAEqLawus0O4g6eYfavw8aYY1RZHM21PUFFykV6woFr5/EP7YhqcnaKdpZS++UT4
rxY6g6faMKR46zIBZ+RaeQypR2AxyE5dNOxhHgiATwVg80xG/U8hsrZ8IykJHgcC
e8nyDUH2BQe1TjN3GgIHmQsF0U1gJ+fDV1vece6iKCvKtYFJcO/g1TY0HynwPbXL
7Df1OFUbmfLP0e0cV/gyhjvYu7MgNRJn5kyT1RVT6KrmQKo9nK/k+HlbzK8spjZc
QP8rjY212JKAZaQzjvqPf9US+jjThCVzZiwSqnxLYnfqwK7GFLix6vb7Z+cqOIy4
V5iZYAEBuZv5XzvIJDnTLXkD2Cwwk6/WzTfxB+l8FhMe94KLdaP3oAc34gViiPci
Ww46MLArciyFfWNtOPzmjyrmy/jvwf68GySHlD9geQ4o7cPwthGqnERn7NeK0ClC
U26OwmTZwBjx1n96hnlE3dbKemfL2BvPtUF/5AJ61HxYgsBKJT8+71KyBqkPswaa
X+PS36ho4nyVvxDqiiY3JXjWOr3ZWNMI+FoudE0edSkjTT+BWDNEPH0Dm/QpIN/o
aP0XRqMwuCYQY3YDgBEXHRkIY5t2BjBbToTGRRoxxQi6RrwWqGvl3yRrTWsipEUS
KWwvXnywcDFf5jEdzIA5kSKUg+6rbg1j2rjaTHFNpYSUiFFbz4ftf4UjSAuYebsZ
TgEuFqdEYl+RJV60Vhv89YVgRt9idXKwKpbEZZarxEYDoaynjuoG7CY/+UotbZQI
SZ8VoEpkWqJaYgmaru45QZvnvm5gktebv2zIZrGJISwaO/Ercxne3elOS122dGVP
zZ47a+dXPNKUY//NAye88HavQMRLhDRA/o1xiYMEUQC4qEMGigoMhzdMoMMGfJvX
ZAyaHeu2BKmbK7pfZSUgEA==
`protect END_PROTECTED
