`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HUfrxihJj/fJ1uxoh31FL8gz8m3vjbFqZwo15orP2b3disoSMk8csGZC56SZxM+S
AJQP/2iYL5Rhsl8ypSMK4scPQqQzFKH77R8KD4CHqILBdJKbE9k1RRAbSTlGlM+x
cAnee4fE3NfkVat50wFkbTaH11YDkX4RUx2uTuofwYQX4CEiaOr2qIrwBfZx2qfs
FInKDc4xkZ5v676b85NqaueGcPDZAdAvzQ1Lvf6ogsLl2yAxoDc+C1ayHxevpBhT
qEKTNKF/lp/hezZaFMV/7piaCvCg537AnGhDcPrndv0=
`protect END_PROTECTED
