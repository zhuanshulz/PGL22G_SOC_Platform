`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DqCWB19gIpX5U9lZsIlLItwqJc0239MnNLCKTlnHr+I92ZxxWTtv5PXbtqa64/0u
bDl436Z5w8GGV4a6ehCivaHnNdE206UY+37I24KJtmz2RYyjpwrPHO5MrR9uM/AJ
pUFOsTweUgvTxSQB03tHqQQLkYBg92AzLDILrzdLtHPuuTNaQx2KQKo9RUwh9zKu
yKAU5jqT8jQ9nyqK8kums44H+nIqosMy3w1o2yChxRWiLxjUrxN16R4KRrUmP83V
ECVM+DiDyVahgzfd91pisA==
`protect END_PROTECTED
