`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3vDf61dZ+KnyiYc1lToOE40RorMDL/PH/PUOF2epCtCWoY1eASHZMsXraggiFedu
oY7hJs1ZTSXuUCGlra6afC5FD+6Z8hdrLzs/kYwoq6BpS11LofsBsTvgBkFMaBuj
Lh1eRIAu3Vf+ptgcvsbWOqKuRC7QvKGdvBDP6fdkolIYt/kohp81qB2b3fN9hOEu
m7GLGzcHQ4cGZwbbi2LcynWhhoD8oEn5Rf1xuhDS6tZ2Zh5VsSv2UUxHQgHTPjEA
7HP6vjdkAVSAD2XeaJo8q4kZV5YrP5gXBbU3ADK0Wp3/fzOQwvdTnh050wKuZVeh
CJr2CwSp3qEgJ3iZEUzU80g2NmBHygvz9sezUyazXqC6aJtVcIq74W2YqlnxaY7a
Hi9ds4md4byK/XV9u8knRaWjCGbZ5Z3bMaxO+wlzRgLgYXovFLmK3/AcCqICyAot
ZgpurnXsyKf2cDCeOSQjau4sjk6UkLvCC6fBMdHpl+Sd99+lQ0ULD8zVctFSBRDP
W1OtZLXuZFcosOutXeO5RcYrqZy7QxVS/ULEGCi39kFgxgB1+Pk0QRhyzkPg2wN8
`protect END_PROTECTED
