`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iRtZS+U0GDdMCBhJ3EQ1ekv71SEdBFJ+fPsOD3gkDDYFmqKb1WJbzqk4K4aoea7k
UTaYiPdILf/dK06O3ahR7tkBYbLNHKIoh0UKBpnG4GeUORieH5aYea2lVsOIqoGS
OilMopiG2M2IUxqjCk1vzrKePU7B3z22/ViB2fkUeMQ4j97HhH9KsLYUxuK5KNzn
C6561dIxelNzlPFlojsfQFtFIB+/jzKCVM+Xu7KbaqtlcDo7O+Pu3XYlEayhILK0
mu0enQaILTtW/6PcvuFLR0wTZyzeG0J9y9d1/P+CL9hx6eM5QkiHICqsqrYH9Tl6
5SjmhxxL6wlot1sEjXe+qUDxT3hIvgngomh4O60dGAsqv91+SKFKzkaOe2Mm6ekj
l3vv3ty6qsZzDRC1q1pbEpuwsj6RTD2ykdINoZf9fi+HgZZn43nR9UZHP3tlNuwW
3e9Ja1CTH5HsOdL5RBmJ9fZO9apcokJPTfV/DvTM4WBqzLmCDT500gpamEiYSILb
l8TFANiMQyefxQBqCto3p0Nc2rpCZayjS81ZcbuY6js7KxGthulfLzQp7GNIExXY
2H+ZjLCiRKwDVQ7Ixw9YI2YD8ggfZjge+aljFF3N6Ypjg9f19GvuBjTXFo4UqKR8
wz0BFZNhKrCOxcNce9E1znVA5UsW8MlhJBU4dvlC2Ac2SBFRKVc5teTw4XPofihQ
Tb2XdT0iHAPyEMi29PyZ/vllrT1SDRhdr0vgS58nM7AsAqtOw1oj0bpJTBCT3n1e
7DAjDPZ+vG99TtWXYZ0wb2/zmbiermhm98yOVDcGkmuuCNQZcnZRCth8K/p8DAj1
bUrxA5uLe2H+hr8BdkADKX0obw3XR6M0I2j8u4GTBs027B4Niye5WU+y1vYIwD5Q
mLdLHSeD+as3WQdvzHv4IXq+A+OWLBW2heTZwheRiESicOXn8JrssHy63fULKhZx
ffxL1TV5v5wKbwqGMl1fzbubjNPKUzNO1/U1UCMQWYWHxTrffFf+R/9V7IAd8I3b
ZPJhwL/uFQ2bqC1r1Xa4+zm0JBaKbVbffcv/QjKANnf2v2auPG4eK8zqwJRv9eVI
2Guf6P7J8tI3NMbTm9hrNicHs4ChZ5bS3eL8paSiasT4RQwdj+crrN+7S0XKvJwJ
p9P+x+N0ucFl8xchNq4A/TKxBIvskaZCanA48fNzj2kFhRMPLymsNS1BPy0hCgFc
QQsYw5SayFOEoBLDwRF5QohuRkgdnLLQ7Zc2z1ioJvfTUv7V3oRGtTfTs8mRqGjj
tqCo7rbPNLdUVhxFhB8e8yvnwjWGedNhG+nzU0902GjklCxYZZAIe2rKPldvU/Jr
Mc+o2N9ZLe9ERXJIHvCh9McVNhffRqADI3SV+HR/dXA/tTv3STZZ1fXi7y+iUaWP
2/k/SYensKUtgBDsiHEt34oF/2i/XmA3ia4mkg4e+Wzf0w44dPaoWLrKWYKy+tIu
sV9RuIiFruDlnQ8K15n0EVANksB8/Iv0xNL7G4lxgaTt6HbCOBLc2ljyMpwmjVo8
6FN8xPahGuv8I2MK2gIQj9pJsDdujpj3hmLIC79Zzz8a8NEom8WpFvfba6YdiVh6
wmZjzdKt2jEVBo2vI+u0CjcpIuafawFvGqybCbr7tXQll9yfW4H39W6ntxv0QF07
x9G690NpstMfnptd8UjY5rbHFqeZ90zyzOkyjZ5OCxN8TJ+o8YyU7UhCsUi4TPdP
32/DOfblkiaMN4lQ5VFtk9IPOgTqIEJXmKi6yx5Y+xsANQ+okh7/gTTqNikbBeJj
GSfLWgXXFnz5tJrZ9PzX/WZB0NNbUTz1mmNqH7aACcyVDKjWxqfr/CUWsUf/EOF7
f2oAFkD2AebbnNEkj0sXIHkRE/URkk1kFS+DARiIi2PYuH/uO04AuR3Qnhkm/kOT
d7izDFJ8S+sEmHP6BigLbK86kJ6KspN0067N33wmetv06UngUcSiblVhLAP6UvUN
kpybfoG+qd3zBSSpeYpe7IuGdFYLzE9LvtCCKccrGYrMihoP4BxZ3lcrg5D6lzFk
TQVgPEMJMsQuP03R9GOk0fOyRa4alZMZpa/BjJhWXApQJF0+LAR4s77tVHqjfLw4
lhC2840kdBAZg+XSh0zBi/p9XZR4cRr8znLXXXKPAO6vQf9i/ltFuyM9aW7WRXT0
yLEtvMYccD5ay9zltiPkohQW8ellTFJH7gYYRWE0nhuffoysCTWgBOX7+CoGKuo3
kYlk8E+br5bBIwrtYuGPZ/3qrfLkynVEJNNDowM75SR+K+vVVRsyDd+tmFacYgUJ
+J5UP2Sjm12VtW6Os7d7vGXOXP/csaoCPoc4cSA1vduxwd36AhHca2QULDawb5XA
PL8Nf3/TKv/yrGRshQO4bA9XRKrE/TYaDSoDy/TieA7rX/lod0hrl+qsW9UrtNbG
0V2+UYCr54er+jgsbuGDn9Uq22czCJQkHvn65pc/MZWKxM2fqIuwk2mHM/OF0dMU
v1Ll6sBE+VT3N0eoQhvNhD8o4j8BkCKgJe6IG9zWosfIhqnPpqJuIsQx+GGQIQ/o
OlrgUD9d0kOg6JYy5UCso7mjMT3l9VAuRA6CkbAY8Xfy4yTduwODpZ5fE68t2M/I
4nqX5RfoTEs8Xt66/en9wORIo2mTOEkaHXr5lAtUa4KcjY8FqdmcHnEFGGtvOqtz
c463/SWOkGwnhgHwego8LzYwa3QscWgMeBZkDh4s6fuLpXKV0ZTcYwAE81jXv8vO
HOxxmt9rztLm7W7c45SYVYlwxlLSvnmIfowda67o5okFmrOiSfmbKbsKrj0MHyte
iMHP8MEO7/3T++YHhP/ero0tGY1edbNp2FGQtAp/bfscKztM5yXT9n4hYTph+aDI
owFPiKPhBSUJEYFEQz0YuuaOXKSIJTY9sIwgjbiW/EUVcAveGiC9L91RCyPAyKEk
5qPWfT6TZHz3zk1yG8miVdMJmsXufqfTAs3k5qb1197yxAbqPwgK3aPPMMTWc3sL
RSWqCKX6VhZv3MrTC6oDDVMpl0GyO+BKJeOG12rWio7Q43SLePClawvs/q8VLyOi
yFPngpAke9jljNzALG8LZTNSVad4rckKGz+279AYEjoAVb8LjiPnVHibXXPlPcW+
1rDj6TLBxWJbwd89+weMfljpNqn5FnTqhIaA2ydMfZRxEfb01uDfWSqbCBcvh2Dl
g82fNv61hvwTU4XJHMnYtn+oExWfhUwyaiyl9WVSBTma6OozNpTltsETg0wsmK/P
6WrKhRHqXZ5RIX4/G76uXDYeZvWA2p8kfGaRhdIxUE5AhVjuA3MCG4+cWEpbyXZ/
l+p78Gzi9hxiYLViPzyPGSPHOJOIsdeg/EV3BrRXQiDfkm1RsvEd+0AXpVcTLZRq
P4Yy1hTRBbqI1hTanEPXuS/KJFolKvBUGwK3mfJ6kzRpigBYjRJyG+ZJgumtdAjs
98qRaMPijQPXfEy7F4Sj25L5qcwqJQJJsEERcq3eV+cBWxgK2TD1TD7aLdNnIk0S
z4283NjtzSNzogmBp65ybGC7BKT7reLbDHz83FobNjUcc2ifJqNOyoai+QKoZZ+T
87xdYng4VSUrACEGyU2foAMM7uEMRo4qo23C4L0b2AJupCwFuJfP0tYxkV9ePock
9zI3IrX/jC6MRP5SaCvk23lQNa2DjQyUaeVHA+S59shD3E0CJPq0BvoykjXQE7mM
HABzgS3tMbXQ5P+G5243M6gmyQH1miBA+hCyTLky274CvEW6O1q4uMFsP1aF8MHs
qlWcxndztV/vizHoJLH4j5ljXRYwo1KdpiCGHbTZmkMr+OB1w3/QAvWEbqXwr+2L
ldhtGRqDg/n6nxo4fvOHwGEZuRoRHu+LaNqEzjqFTMkfxPW7AjL+SMfaeO5ffiKy
Jb8p2m+/Ek8pxXwWa3z9jHb2o4gC3i2Romy7CeGYzLM7SRxWy5k8cG/g3hxog6nP
5y6WtAFwtn8TgkQ7gTheYd4TcuKErVvVxsPmOESQDE+cbpbzWEnwRLjl+1zVRcsu
VH31SnmP/LgPtAbRJx017hcgBA5i2pt/Cm6N1Nvab9DLM6zQuNYF9dUE2gFazK4X
olh3MKry5D1VY5B1wTQlZ97YossJhi0NI/wjMQa4N5yrcZOEgzc0gxjo9612UxX1
cWh6zzzKK9ESWtqX38UVe/3636+hJMixnT/yEmIgA21fdHI36cxNWfACA794zZLd
eBpr+NjA6x74lgKNyu5QPMaYSxI1XnpxtFNPpZMtJUQBlBmXC+vuoHQsYtuHQ1Bc
JFwmT1J9OTClkLc8ik9C0eBPj0m3zcmszVNEjFV/8x1+yLBtGskMIUcRvj4bSz9b
S/MXfu8ksrDf+AHN6a/dmIYyEi7Ppg0BET2nMzMRrrH6OL5/Bg1POYqmcjJpAHm8
jfVjlhKyVcfTGzfqpgujGqpd8yM+83MPNd0ewd/LjqMRcdRhGMwofGVGS/mxEPqz
oy+jFfnFi6JpCDkNnaTPClS6ZSAOnoNRK6YyVXWJUQSaC4j7kFEGlo2AMchEIWK8
QZFTlMM5EsrPqkcMiDrQo0ECBW1dGQyyiIETNgHNCKAaxn94kNO3WsMnn+tcXmbn
+2cEl93/i3XflisO0qWwKGg21t58KCvwXkW76lyc2YQ6g5PINOqMQUULcYWgNbc1
O5w6emP/eMBNVo9rnR15WW3w9Bn/7qLKYn9YepsgeK97mGOCSGQsbXDEBttm9lx4
KFLyWsNF6Q8ykhJKnPSDWJMeh/FZ8Z97EK+HVnDTvzqO3P4iZ3apHd0EuzcLwQtF
vI8ZZXmCzaBjEnfBC+gKKoKC+sbDQU9U7cUGHoSacsRTz14ZbhNbg739RSC3v/CA
txcGBnOb4Ig/dEkttTWv6+IUO5GMUGGD23hB8LMkwpeDGdAgGy4Appy71jAcqcl3
KvCSehL0IoULyPsRSQ877kVnuXzv5k7Xqwsnsqt9aADH7PWpto41Jg3eu0XO9XYV
Y8I6QL73ASPXAGzi23n49BrXvD75pQH9aM29IYb7ZSUtMSztVA8+1WdEPtZRs1KI
nqlqAHh0Zerd6btG94NIUDREd0oPqnt3RATJzGeTPOJPyHCsw3BrHGz/Z7RESLg+
rlET1tZV75i4VVDrjYBOuXYrYsu60iXy4m4FetfIBSLoxCQdvlQW8B6tYrDEMCkW
8KeVyiXDV+kTGxwz6QvQzfzU1L6NAmafhy2HfC64Y4W5TvPPggDL/oiE2zlr6vvZ
jTsVSDdzifmBa0a1js+TYZSiYwRRehd+U7A5VOpZZuUETumWNvCxdnSLmJcPowjY
U7NF3qU5Qkn/4S8Gr08D84dU262ehJrj5FXDzVgl0s4AdiJieO6tXNFQ0Mw1BNgo
jEFt8TOA1N3II75fcaV4g++Us2Gutz8MQrzh8whyk4ss8t8P8kRru2dGGbstL7WQ
X1vlI+mupCxf9h7FvIFevRMRuHqipKC5VfDbMfIIv0BlXi38YZ5dJiJTlyyC7k3t
TeHpNX+u6CbHx7mbuyIDwSAikiGIdRZXip/BIrTqOZGfyWCvraXub4rRC3aJcUUm
gZinCFtGJeV2qXcBxw87ccpGaup0fh+abv19IsfZStvrPOEu0zzTx42W5/0T1BJ+
zg6TD1zNaDoGqTT6hsIkl7OXhztfi/M67tCaML/LkDXcnr+PFjnp2Agaw9JGGo6m
h44YC/FQ/0RW4lXPv069FCaXaWjOaC4xUcDP6Ei9Gg7TQu705+RVUnuNpqbUM0Li
Z1bnomYkkDOv9cfNXAWOao9gRqZ546pEN0O6K9g5YISdnoUmU2ttsxDdWfMGvrg8
kyhO8sgbYlYRGaVaq3qKV2Yle1Pza48BoCrxMpX1t1U0CcQhwSp3Eyehr6m2x6rg
Zz38msdfNA2n2zhB4RN42QQ4Y+WXZNo9FKsQ+gl+5psZ6lm+zcPHhvadlK5w4Q/H
7CrVIGRT9mvVjzGrlz05YCFLrv+vXlHxxYIXfgSNETimjpLCh6CIkt04qSgYzy9E
auMxrzdL9RUCwThKO9252c4jC0AcAZDOGcXHjE1gvQ9d3OCLEUeqWDdGl4QBXEy3
QekqC3lwJ51rOZvaSQvT1kthFxTo0yC+d4sy2y/ech153jMOUdx/laBbLfXyaI1M
dQVXdwKElUqryi9DTIrT9ysNzg2UQKKlSWpdmI0n9Vitug7EiDaEAaXEeTs6NSkW
HLBMldAyOY/m8F7OiWiHTbmrArTodU2dRZA/wMBGHTea5S9uoUo+fNOUofPSkABp
XoaFxdaw0l0bLFH05v9JPjXPpcyBBjhz6fZpPQpIlKYF1rDJfN8Tn7LXM4QJx/eC
K/CKRSKuw2iuTxySXtnCv7XrsWPlxmJNSUQacST3akJkkL4skyFQgq+zeq03wjE4
LEZTcae5l5u3wYSb7C4xkxLbU3ASULnUoKP2sS+lQCbUEPc68p8aZT9AE0jPoLQB
tWnr8dPlljpYCGUdB3IBhwGHqmdZHBi7bkvGhJDcjQNh4Rex+43NfGAqFf7+m6qL
8V2EtSccz1kKQ5c8OVGnjdmUfEW53Y/MWLrKqDJLF/JKxoqbeFEVmkbOzDTuFzlD
f26n9jLvPQ3b6BbmANkLNCjsv4mti0UGQxw0iMax18B/R82e1FLp9oDjXjtSEAfZ
zrI3KyyiLOnu3F41qWL4cneLNWlJnOojc+qsFH7rhm7lCuyrv/oLTf0P00lxCMQ3
xg82Uy5KJkyrCumUsuk3xjw66lEN21TtieWAx0TEo53rrtCHqegTUXva1rJd/Z0x
M6NKZsxR64Q+Z4fLEdMWRn3lqn0ZzYgatAT8/bDPOKC1VkTr5fKloSjIG1kUbSHa
9BdbK9NkkKp8NlThtHZF0gF25+b39DwowOhF8Hs6Dh8h1U1qTSFE+26bQWPJeIjK
aTzt8RZTadQp3d1f8KrObNuQ4NE6TGQSQcdiT3T6BvUdFimX5zCFVoVXc2YTozOL
/n5JbegIISOZ/nxf7R6t26Y4fmklhZkVaMnZ61RhIC/4ubKh4t5IAZ/10wfTYjg0
w+tNZCkKLpPgp9Bbs1VZIZ6Y17yLLmAcANiCNhfz2EZuWycsDiZ1jZ8ZFW6Vvdj5
nrf74O5rJT+4IHQBIUWiQu7HAXSJ3s3XuGd1nE6wPruFd5DDmbrotTenYS2TDNXo
Gig21omKht75UPeXrz0B/G9tRSib+gtNmADRt/Tp5o5NavZtGwd0m8T7iP/hFt6A
GBipnybAqFxFExnTZCF21W3TRJqh+O6HA/ULB7DQ+/2xBqKNZ0yh7i3YbraIPct2
n8kmUtDw97jJxKZY+bGC+cwnkqAjbGWYAjs1Z8Hp4aZHUbddbMspXmFB/E1LjDkQ
JZTP/LSROMztRNpLaHBV/NM5I6ztpo3uoFfda4w/qvIJsVmk22IMEdDJL1Bx+SLi
+1yR2zk5dOQ0Sn7jdJFjRu6+QTbyX2LZdoV1dxYT2Qd67Xu8kyp2R8aZuu2SnFtO
2xqYxDsOJbuvNATT1Rv0BzJTPK3wmr8YKj/4R315tUHoi5SzMm4tCrFx94f+mwzX
q0iDiUttxqeUwdlw6amzRRqpLTxPrBG9fTjuwSjd7Oz/hJIS6r0c9qzALUlKmw55
xQ0TTn8q7utcoXlb2mAhTkViBLD7tY5shbo1XbO7gGpbEInH+cLTzCMUABKBfcL9
Qk0EVGR1CTkmWp3y9oweTtvSpwv+Y3sqYNQGn8xVlxywis94nRHUFaAyn52vik2b
P2v06iUuEI6UzJd7V0q16ZXdPCpVPvZ5OYQ9IdAbEuaEIsyPb+ZXymKhiURo49Lj
xo2T15+z1kfyw/kt7ZahuxM1jw89DMCDG3KukVdVxB6fz5upnWWFcjEWlH90UHMi
clOm6/a4EgDSyXQLHvvk8isLq5cqBO6CyxOlf1LRJ1Ab5lJ2+9QuOYQ9mYn+C5ia
JhdVnKaGB5tYaIaSjRKLAArdM/u1uoqfD9ubqj++XOQE7qjQuOyMkV16sYKkY/Fj
phiTyHeQViE8srt0FQl7nqPJvKYdQFebwihDGVOl7BSU54hyUJHdoRWNh4pcmNnL
lsMGYcpsgHeHg1WKP9AOgGQwsB6QnpAn/CAHnbYKddPjEY2e5JKakJTddmoY8sK/
kWWsE6yf0MNIa+JqAX7tCFU93armFz9Y2NF/i6z2zSqWolOCVTG96pnmRI1I4ayu
mbeyYLWmo0Kg0HSUjNgvDr+cOUUvR1VOA7BndYE5IsNWzdSdECyMTiHOjhA2gmgm
jPKAfg/2OYkpmPKL8nVXkmpDS9dBL/GqldRwm+lbU6mZ7JCX4WeHKx0uNJjgknv3
aZJIfOPg6lYy7ZYDwfXFXF4TrF2x8rxbK41WX+G2LGneGbGLzy9nzHh3naZhVkB9
Ifzn0UHF9HKmblPTCBmehwcPcVA0wc8BXvbMO7wan5B0RTMdd0NTEzXs8MgN28Gd
ngzqOk5Yh3+NFRwa1K+Ystv+D4N+vTZbsqOT1wUEnVfNocWSsaMp7cIQfFpkfWwj
PeK1dan0GCS0A93Vk78mClUksCUgoEtkfxHaK7OVLeBplPdEBoBV6Y/zXLuxGIaz
RVbSKc7+ByPZ2o+7KJPP1YcjeAAI48TO+HumwfgtFul4FJgUS/IN8hvYLUq66jYL
l3Tb7C6CWBBQNNRnuwb4uj9G4MVC64ZRdE4IUSZL//hmcI5XUMF6+ybAX0hx/Qls
M6nYnKLRFmiBhJJaw07t+/gZGKq6QnzoFWNYf3FNGpKVyd6c/Z+C/goaF5a3FP0R
w74uTlKh6NwsRnx/39SGaZlxaqoST7VOaJLXGBS+ralIX6TJObApAjxM35rI2ghh
9BR0uwpP9QbkbFWcjiOwT0VJ4eCumROcXoQHZxFtFaDJMI8gzoDjFGNIlhyDpzvs
q//7JlOYGNb0638LD47WAiRfx51xER8pRTjHPV18VpbkRkxabYLNO9AwQuVH0iqp
720zL+VyEeHb1GbrLYhNl1yMD1GbUVrCdM3yj1Z/FewIvie2tdETcFB52oW+9pfe
lHg1mudV9HPIaYHCPEy7w+cjcv/Q7qtPOAXlz2C0zM++i/XF8p//uYg9V8TZvhaj
dlvNKuSu9cpJ23Uoj6VMd47CCB8F/BsYNRy0PM5K/+OL03yix+xKiq/j8teLKUiy
KI73tn3iMWTEBv06Imt4slUPRzjoQjDZEWlAH6/ASfiCgaHFPO8JCUpK+OqIgLdY
a9oVAKVxn0HJpltbQly/rLWlXiOj//EoqHxAFcVsKl1Uy75ZHw5+z/Ud/K2r6A5g
6ht9zDsjrUfiQRPWIXwDuyY6ZAufUIOarTQsHWatg6JQIEaRG5HkQ/BsGSJSr9Dh
fPE44RTO5hSL8XnEld8wkt9pzvaCu2FDtfj5xxbB4R/DMinOKi+7Cp5MBSif/Cho
Iog5DjvWbowo/HsvuvNGbPmK3lU6qOr1Vfcs/qJC5J4YuvWxQUvmwh1NbZyjUwpo
KeKlZWxhKfHgKkYWQP0sGXp9WIvfa+MfdlaKsPDcx9xgVFVMzCUvIFCvfXB7deUC
QgewqbE8qhV0TVlxfay9g+ovfTH+lFSukgT5cNuqoX2d2LKGMBdlH7WpCKqLF/9p
koXAH+HSNMz5yy8XZt7Y5Scc3ckfBSQjah4RivP8uAhWVtU0PYe+R4cx1Zd1iWNq
K61ePXAPWdei72jeJJJXEID/rfQdEw2ko+L6/DxCDW28mK+8K2B33m0f6dce8vCq
cpGe4CmwJbTk26rxMDKam3hT7Z/1MQoazbxHeHtyxYK0t9v9ReQQcFLnJ57oKeok
FJmvFhl7h/pegTwsmJq2lw8xARK0R87nyfqnEq5sJSxZDFeQLcFMVOAMdZ0ciYey
aX4/cwuP4gbTCjbBG9G9PIqEMIm956nwpef+hKnIqHbH5fGvD4NbPGFMSNSEJbxk
w8+rxrrYs5tZhZdieznjWOcKR8VHTncs8C1iyG5zeqUpjI3tr6KpyN50jnt+oACK
/qqu+uDDBeC2V7UhdEyGOFGJn5+e7vQ0esJtqu2On2K/N2beB9H2Ge58+7w+mcZ2
OHcSW97ov0VzDH9w9Aj3LGJGe06AwqiD5VBGuffK/h912HjbwnrDyolQqnwVDao9
TQ6t0sL69NXk5n6dPpUbiCKr9OKH+7Bxq4kDlPcxnbukCuum4W7OjEb3j5lxoBsN
QbOhfuSsyY2y2A6MuGG/AIAfvJSD/w0KMCkEg+scl9qUX8Q68OfMc82Fu8USCU4L
CeMfC60byuNkTpsHW3pgDod/0aSc527UL+MFmBwVsN+4XpDXRoyES1RLKMsHFqfx
VZ+ZnKWogpk85AxmTjnenI/vYZdNUfUG0P9N3MCm+QFatauHzL6aXb3FoP6mCuby
9npl36lUGXgqPPWmip0u4ncHwJftpYdUPDiqVLn18tczhzJxssiyUAn/JQWkp872
ozp0/mOeWrirWBQfj8ZcAqcDmKjPoSkPSgCQb3DMVKuaU0NbpVsj61r/0tP1rGF6
3JAdy7NPUtgOtUQmsy/djokJftKnMdvoIYCU/X+TsCCNeO7EmC8ODqM92qslumMF
/zICziIw+VoyufKZ37h+B4N+YyWPu5HnyCH0usBCRwM2uM7cHlc8/8bcuex0MA6H
lJLyrPVqrvtoaGSjvdPDbGn/jZeo9kgn4zEE33AcrjSvg9Y1XlPmnxmbpv2/dzhr
Ug75OSptv5Xj9pxD5QHzTE8mwoq36Kx8FJomUf48fFa58muPAil+Xj800Rt0/JSw
EZNYDS3jkBdR7NT+cTvpdxHZ9E87kGf38eHA+KDy6ZBeoLC0ZQKFeYvNLpcP5Ika
XNW0iWj/IxaagtpU9nPLhqNHpRRIcndFt4ABENmT+TcG7DljA8FrWW9m6fE1/4rD
br4yofkmR8L/PtbQipgnl0CbyM9TuDpRwr0q8I8z0XkC46huFq07mSlYSvTZQW2o
Q3uWpEOKnYcaVrk8ht/TcNNRlsLBngh7hfhMlJCU1thTjBuvp1PgsUvGqRpWes1H
LyjFxd0ZSMraaHHEQVAa0ok/7BYeHmcE/dl6qiIYDHGOR0X5DpW4QD1fTVGWj9+j
0c/TUU2BYnFC+mX+8MTNTwJEkEphUYYvkvr/1/HT7bmTr0Lq4ibM7huE5CUa3uXn
VjEaqvZkMSyoXnj1DVa2MQ==
`protect END_PROTECTED
