`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BSvxHa8oqVfWfxtYpvU2d7y2TF7DLWpTRmXDLCszoWbXDvLT5UXM5qKVx95IBhKt
dWjD+W/k0PrzdDSnokxDVdbiF/znrxKJYq3eylzYyv+5EkOvjYKW7m/eawu7qiLI
YJmP9cW3N2PPueQUQOvcu9t1uFUak7+452sL/PxAj/vcKz2W8LedbfEoGqvMjBa6
VvR5Mhcfg7Dszyq423mbGxZocanxgNN/EBY+QrR1HGMsq883jomfU1S51HiqIWAD
rFCSxCpEeT1bMUKSbtZedq/O6Y3PrhXL2NO//N0mVcEJc2Z3carjN+uu2vxaXWFd
9uysZLZU948qlTstmsLBY7kBOdPQfBBCcXJp/47cZFa1zWi5bSjKwTNaZw0u3hqs
w+TY9xD6Wywo9xIRKSvVV9IOY8PEsefuyskqs41+GSyFKErfc1I4h3yDU2i1/T29
UmCQGxuD9Q8MSDdnOMZWG2bg0svGx5gqOYmEmntBri2KqnNP+//OCwNyFqsGklVM
HelMdMG1lcxsj8OK+ij/O/V/BSfZj0/mnJ9vxaT6EorWGh7Hd0R3Y5alhCHZ/e2L
DX8AKqrPNzJi5f0fXNBa/9RFEEUZ5udu3P5KVNqfk12OEtFzgTNNd8VRSCw6O7e2
qm/tiPy2NXHigS244UC4XTk62r8kRVfRa1DBiiRQNy8R5Ev7LjGbE5eStOt4cBF9
FlfoN7+O8SbqziR05AOATxjTkqSS3BUoI8/7raWVr9waEcmFNFeL7PP4W4IE9JSG
amWUUQkopXyDW9rEmqAToRcwYje/vGWZrIQko/sLRz+xbaF6iIRNX69qridBiggR
ocz8EpGyN3Lp78CnDJHjTbN7E91vP9mKbNlpPaBGR6FQ0RkLT9GRbT+GN0GAgzbI
LfZp2bQJrCWRtZuKj0V+C/RboO7FRZDDhMQhQp+ri0S/8+7sKUovvKLyHzCrmsvx
kz8N+iBAK27E9xuek1zGtXdJbJokjj5C0ko7Wfvo92U=
`protect END_PROTECTED
