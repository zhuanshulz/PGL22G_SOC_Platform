`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h3b6I6qVnoCJq0XmTgONuSGZTylIGmwAbExE0RxYB0NIzZ/yR55QtnJHcxheMoeI
jBD0Vm0pJA5FnVODP6mqB3nPiOXzJXoPThiN2gU6gMo2vbzT6QYTVBxukdAzKeDr
CWcX0sQQ42l+CoL3VcHPeJJWtAwB7Pr2bcZbQ36LK3oCo8QbX4pUuR8sb4xDU0uk
m+/GkjO96jWYAatTcXJ9Lhma5Fg8uy0GPwfVAKORN5lyytNqAQC8vp5semHyU8fY
IXmn0ae4YGHjCp+uADmrwOa0HzKzQTyFnkpDJ0DotK9Oo9BIVgV3DlAsK3cFcmcB
8GUu+L7ZH9t83D4aLs0hbTrML2WanDA+IzJfTID9OSknVJXJ8RS+Ia4tAL+x4w9E
tpFKeE306j0Eq3p9Fy+Bmp7p4KLj6T8tIbsQ04+nR2bHH2Xcirgmh390A0wNz3bz
bCJ6BZHNbLUmgTp6BqP3d1iZk55/jHFCg0hxvScU9H36X8iG4OHric1HD5kSk+hD
p1qNNlOQrXbrVdyiXAZHkSG+X+Oc7t/N47I0CNKIs31outZxhD1qv/M1+L1m/HeX
sIMIcNbTDR6ZouD6PPV8ziF0pDGaa3BrUt2Ns2vkgJ6jA2AXUAMVVe43I8UYkaSP
T1FW2js0XpBYxvs+TG9E7C3203Zjc0qu+lS40zVU6BaFo0nwr6pQaVTD671SPg9W
b3Nkjtd6JdymFtjr3l066sCp2z0TwilaAqrSGuMkcIifDACeob8feX3L9fPEdS9+
esojyJCvPHC2LX/+neifH+N9DzDgeLx3YH+luKHWsKFziW131F2MoReW+4nEzGf1
PP0EOgXNDAqmsxOtLaI3DgWPjczvLgod15hqKMt9QzrcNeKfrrfiMqSURdJRCsgN
1aJlMvmoJLvG4VOI2vW7p5ISYJZ/903OQjaNiWBsmHL5VlZwm81SX6lE8/iHP2YE
toKIURPqKWRSM2aEuuq58bIbwbOzQC7RPMGWKNvlpFeUCutL0CGFgwfvR9EnWiY/
LLkmM4J/mGbPia1PhPVfHrspC8gzp0WsJeRfdsNXzAGGjr2hucDsSXS1OS6ghfIw
/CLypZ938N0+CZBlG8BEB+P6exUtFoqW1nLQkMAffZVwrB4gwgjk6xh0YUZzEWlH
Am5qYHUBuT1Of4aGDXsiN+4nwcUXH6ZG5p/8+uyIh8njMpYzZWhwhCU8af1CZGR+
wO3/kLLpASHKR1MwmStrqg==
`protect END_PROTECTED
