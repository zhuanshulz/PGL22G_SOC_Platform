`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hyU8UUCE4EbRlwIePz7FuFh9B1+LouUsoa2STec545x5kKfrQxUWeb5BZyOadoqT
ZSTlYJ7BfFX79B0PWAn85HQJxkeLY0vO6vdrvFGQG8dQnbLoJzXZ7GXjYizOGbRt
yY93HKvBqU2qbexUrXehrce5xrMz0Y86huO1fc6X3iUCy5TJ+IJr6mC/iBLmcm+7
R7hoab5MDSjMRzjrRP5pSIEozQF+oLncXnq0NC4bIu4GPhjMM9mM5OqLwxP6IIP+
anO+wVNrHZ7876LaktW/XoSiv8WKd1pRNX1fhayK9STHe1w8rAiCx1q1IDnHsixz
le13rtgnQOHMvzY+g6fKog==
`protect END_PROTECTED
