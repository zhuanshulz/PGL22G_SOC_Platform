`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nMilpOv1Cou2ImH9Cj2NDCHnSc0PUK49F1tSOSq05q5rYkbXHotT7weM8nUqUJ8u
ZjE5V7LiZZBMyDbIRJmvkN1T312iFOgT7vKvQUh2Z2vdf3nXYuyKp7Mxvlm5gegv
xYpKCN12Kii5pfDTlS1k/U7iXyZuenUeP5xC71cSfZCtU2tdH/OqThKgEQWwYPxI
Yc5jfYhmid6q8jyXatGSW8RfyhFRCHcybfiTTk11mee/XOSjoHdqdScB9zNEjSpw
KGfF+anwOk7PXuhV/qd99IRsnVPjXISk8SwSmqD9tsZD4Pmx2RF43KKslnLXUzgr
+e/HZEzmXQ37B0ZwEb0ktDaUeCet4RM6pXJCgyj3fMKX68tIBwBDJB0HBAC6lPAT
TvNqe1A2EUPribt7fZX1hnkELUH4aHAbaUYsT1lanBrgKiSCApVMrYmS+uW88tjI
YmH32Ivwhy1V0HkDqSHGQ/nxQrQbySlNOsWy1RoPJ6dH/qvJb0WX+1nR3XS5ukMZ
87GmnfAO4H80HHNFo9Acl1PB5gs5L+a2dVOSUp05WwCCKsXoGszlHluGvV62e0oC
6twWqJb3zq2EtPs5wVjKoGyNmba+zKP8/QDKgDQeTS5pIyXxksVi2BMculwtqkHi
CYrio6N0MCDSH+6+Vv6jMNw6fGnMBc/t817/+Xe77sPY6JH1fXCEzCGYL3h0vdNH
J34XWkW7I5RDqNgLPxFVnQGG3Ln4ybv5+4+guYsf3+ZSFva8R9Zol7S22FW0+iiT
RfghFeT6hpKm8s6Wz5DJYxlgL2iaXB4+ZxwVmQ0UEkzFdog7sE7X2lnIacfl8T7F
8ECAPMBpt8DU4EdYpP/z8LYsQ2A/pX8wphBQypeYCn9yw5/ioYBinqjU4wAP4YQ+
eFTwkcSrU4cZVZFm0fhB2Z4hGBRxDkaGdcq2h5rwRD8rUiyJc83DS5AJ+a+gBt5a
QbjxDiPKa2FK6S735djUQtUvNxmIB3UlDxT3Ml6E7XQFgnf4d8/Ep2ZbW3oGo39+
uxhmZvkbdAv97W/VUeBXjlG3/ayuXGxjNBpXh4/o8ZnRw8hzkPtzxR0QQWLkW5jH
bhmARkHEa9DDOFf3pd38RIV1kBt/MSgJaxEZ/Jrxh27mPrWYod8xnb8KkMKUCYQM
vvo53S0+DcUV9si2PNEHTvsy9TZfm1NYQP24Xp5cBDdlu5PpsgPe3dY7pEQOfFwk
KubfnKnU0D+tt1lNBNT3zZAuidiQ64xR1Qh3a4oeIeE6epN0gcdo2IFYdf8INNHf
gUq5LUa327k1kllGIE90j+gbzgYobSMXePugh5C8Kp9WTezqXgqA9nBnx2DwSfTK
ATMycTRFntTQ9dw34xHbj2cJN2fhTHOOieSC893mkiKFdTFxZUeS/vyXaG+/VqL/
gjNDLE2xlMImlGUQ/mkWjLGqxw7KW66UQl4OcJRJzU90IoTbp2ZZDVwUtJ5HoXZZ
k+jeligCcAkZW+vYnYd1imulJ7r5QalQLY6zaV2HNS2thFFmfOz5VsRhXvgHYu/7
ucxYIKHhDbS+OURh7v5IBlctWxacJPnLiKUUAtDZCQKwydiUgfMYWuk3o4g4ht3b
pVw/Gwe9VWQpZmrATsWf8PbvoYlDJ8vjc+KoxXG6geegNou3oJSHNGdTdrcjTc9f
/2hrtgm7FNbTRgKg5prVgZ+2kbrEhOq1AugTEfJdjT3vKPLQJD0YrR07nVcTOtq1
MwiOKNAEk+ZzZ0G7Rr9FW6alRQyRm6pdqgh+B+VYYVv8kdnjKfawNlk20NjrOuL5
2xYBWA9dYpIo6A6bJm4D4nAYNB0uQKlNG8geff8pMknSY73p5KMfsDqb31u9Rbvr
EAiv/myXdjaFc9fOkUCEEcEwXMtQ3nf8BFTfZ8ptcP+f9gSE8dFRNhChOM33u9YK
M7ZGg7myKD2kjqdvPya5D21TfNjR2woAsTAWGBA7GCYVxbdBUUSWC1vAvyTMM+tP
I017BUdzvk3aKS0fdW0Lk4BHPQiv2GnyTQDLqb+sxSM03RsZT8uarr269QsHs69d
30duVWVOgHM8v/FXDmJPOHX7SZainxPyDsHY5/IHa07/tuDFgwf9Seua0RIzjU/V
xQm/1FhHPUa9ogpns2Wl+F0dUQFXNlUkFHYUq2RlUwKK1zZ/+ziaM8d8rg8VbezI
sSot0xP+1eeAkabuPfcJ6QEV+Be3v1jZtW/n8qx93w9dNiqxt+WnAltdn+elM3pB
7EIGIILBnnLPgHrmr6ViJxwbqvknt4pjscdzF7ZknrKvbaV28FLn5SJT34pY7OeG
S0Pa2YfpaYaveYVZTp0YA3oXUimDnluzf5h3tbUVnQVRAc6j2Me46PGsg4Nh09MC
kOWfrPtdoPc3yxYoxF6iwavIBq7QUntInlk9gxBrHxw1giJHDXB2/R3E0EXu3y6A
puCReYIgRRBtSEvcACaw13WmNkZpj3A5ih7VzosivCNZ6PljI+IFgJ40voHglgMX
oCpAn+Q53/hMzJttbWS1UQRJBMHP7a2vAb5W4utenYYDcDnmIhfeK4rpjdfWEP8Y
72tm4ItrC/Q0ZJy8PC5ihhnMNKJlq3Q2QguPxoDHRst9OABwriP08mLCdj1QCEe7
btANOOKYuIw6GhoeFcn/+CPFO8ZuPrcKzCuz1wnM49m+Z5Qz8lW1wxvAmk5W/mBZ
keGoJ3d9BB96V89XrSz4mm65jrTwsuHtE2IkSgWRlHXRtYgKh/T2L5l6OTP4ApYI
MoD02CpC9Gls7lQTHKp8+dLx5XQdgCxM0Dh4AUrkIciCfEs9KNwjVB+qJRKh8boH
oxQq5AKopcTmH2uioIXeDQ1W8d3B+YTq5aPs4fGFXKMw2qcvRl/udgsCcX/okCOa
l0Nxu24rQ19okqvgKGhFhQn2rje3ACVtoRKOLjLtnSXAHlvc49sAjpCjd0OVASFw
jkNHB19JNI83mzEHaE7qHrJ5cliMYSqDg/JBPjGCGD2OfUeNNtbgRWN3R952LgZv
IDGgDsASzf5wmdohewmf4DaKGIjhJ5vl3HheMV5Hhu2W6SYDw393hkdjLw/LrEMV
HOTxBQ4m4/84ITnmlM+BIJgDxYpQp4BY28Udv/EvbJMbg0qW+bRZ0tUSeWW/ZU+V
1QWXYCuXhJ3XA36oYdkelWeeAldsNb92ejoAnR8OQOC2H8CviNa9NjN4IGkyJ4pb
n3mlTEHLRmrgvVOAONwoXYjidiuoYlmyyvDwpm+jjSysYlXWNA/tTTPkfjCovCqu
b+gaEgfk7nx+Jm90T/GXuR/ToPwOcL0Njuv8UrErsLlGyhEsV2KLvjH20ELcQk+l
q3Fbl2AALZ/qnUb1FL4/Zf/+VcbkZNaexgtxLbkfAOp5s46xg6gJ9pImyevROeJy
EMpxUyOBCQBGofKnnQESetZI3b+mc/oEZJmxDCumLTso29S2YfuN7jl+6JSz9/p/
qhVCKXz4KjY3UulVnCGXyFghqOn3neh0OrQCLFEIh/lJruU252aSZfgNCdLbykzu
5cCYpoXAP9Yh5jYYJ7dtmY6PsUvS3Jyh0TTsLMew65qqV9fIGb1ozyLhv+Y957nO
iwSGLFCyB4cfAGEcqUN2pMhSDodYMXSHJEBQ5w5CB97K+DT/q+B9XtwNFXRh29Nj
yAxNsM9pZeS+kPxa9/Kks50ElmIbbxyAo9wDkKIEUO709c7OuI/gnPsa26gKGhL8
6nlXYp+k706uXbMwGF6lQr45hsg0dTkxTNlHIWGlFp52gD4NE0pvv/bTuYeQvE5F
gJ7U+aRnByUpW2DlVlTWh2DMrsrAvcNCNI6RFmXBEwJSDWspDBc9jY+TtyWHUbw2
GUlYsWyCRft29uQGeTpuCbUjsM1eI3oijQNR9iE5Wg7q7XPbYFWubeUT9U9E/5bp
vt/2a/ZPahbZcMQOhw589kSowqe3efNW9fNMXeWIoRwkdVnuttRqLacd08ybCcKg
/fTWYUjqPChZBYkGbtraRkYoIU19b2JGsPqcx/JQykTSfdamg+9WDAE97N5lOEDH
AC5CSoPR4gGJnro1RkiC0e8k7U1dDN+A5NTQQSGvl6Y=
`protect END_PROTECTED
