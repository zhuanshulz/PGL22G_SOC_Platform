`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0CcvDCDal2T31TRMtmpJZ1dZmBAVxQlp1sCpqdGDSsWGBDp6JKtTQxLsKK9gAZMk
YeTQrPY6/w9WKw3ZKaS8PDlkOb0g5hwHs4fA9WuRi3XKTz1cgUbodKkaAyQo8LRx
inqfb4bOChfGAXjviOVNnrJquLxMQD8kThGT32hqz4c0IT5jUbaB5EgPgiOIMLm+
5eBUCyusRqp99fqHf4p+2HOovHsG/al+m6aQuCPHdKM7ItXDvMdyOBAR4KAsrLZa
oiDIYCLcCLd30lqO4kp94Vp6HrbVYgQNzjD1LWlUMGn6M2/JZk59tCG2yAsphSwu
Vo1F+1IUuUsX9SBFq96o0JROfypEWfriZghGjY/GjoXmyXr+/YXwVdKhIyq5tu4l
OybA84+RiBG5OvCJsJtcj66p0pFl6AE4oofRuljXrRuzODeVGu9BgSVGMTHGzLR3
O0k0154X6w0LP7h4j74vpAhGX8YrI3PFSUpZjdRcRJLmyKGSdMXgTLKiBZjl+uYo
tGornELmcl0bWOcQKIwEgtf6ed5IKooj+O3cX27k6kiAJNdlI8coGtdE5G4KBgm8
Msf+E73lUAjl8zcO3CyKsZmmchGAr31+WT8BqrbqI2elp/vZCtiCq3hcZXziRV3Y
If+y/Uoj6M+k3pjWMKWRKHNxTRot09KmpDNg9+v3s+9AB4Zyh/fiThwUWEe4MsvI
q8wwgJ9HsRRieBnScdfxOSlK3+3LE4XH5rTymWlxjtJuWkSYC6kgQ0RHgqh+ObB0
78eMAnwCxQrM7RunrBbB6aAftjFCbjersVk86KpGNIwfdQdABDILjoViZ7uBpZW2
MSJvZliYCmslf+VkfFV8whbAu/tjfO7bxfvakg6ZMpNQMh2/RCTed1aaK1wjPgYd
wSkWEhGVhvHv8/6vKMbx7OCvPff9EPR1btytdxzU8Ez+aJx/mCDwhpqB6/4hjtf1
DMfb8cG8qsA48z5KGKjmJWJQl0qTYkgjcgjdcJfHzeof/cIPFNMCNKddOKpyeHKZ
dl5L6MYbFMVFY15D1hzcd7TrT9V8MukPckH96Y4opDmxA2SWmgicIRMzEK+dKu3M
mg9CUTVBtxSSTdvL70jcjx0W9OPssWuPqUX/tfUK5Vz22x9na/uIMjYGtLPjrz8s
k2AB3PLZEwiiCet0GoPvBysY9yhH9twpibnsXCGC2RvyxEU1YM5LxNL5pEZ3Q/pu
2Ms1XqZI+kVXL7JoE3BO/KJGXtsna+dU7mhji02/lqz3GKwFl0KpKhHyAg+Il+vc
XFxVCob35LJ/oV3sFw8yOpBiPbkeDxpXgokGPihWYJV5Hpu7JkfcygbXcgwCXKT0
ld51crqYwL0KnF0lc0XMZC8kfUEZHrS+Bt0tSgVssO+1YF618BXayvRZaUpKpaV1
nhGhJgHWtzdsaoso7Z/koQ==
`protect END_PROTECTED
