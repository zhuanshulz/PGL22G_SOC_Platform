`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
llJyzR3iZ1CKc2PP4MGgc8D0AUx3JoRbB64IL4bvSA54qVJyewk/vsJoYdnF6dPP
WhyD1svD47UrjB76pEXD6HlHRy2akXq7HKoR4u5y2awEFdYxBMQA9ybIx/1sOCoy
oe6cUg87kIc/mPQar7TO8EJFF7Z2agviWUy1H/2tG746EGpFYHflaCdSfz4FZKS4
zgbuxZMf0oJao1fx04SvXmNGMOokPxKQYdmiebRSDVBacT3m4DnJIn98laDzbqeZ
FZu5b3R7lSkmW06YjT8xdaitK1hEHRur9OTKN85DscYa+t3NjCFuSndhzbx4ES5G
Q3p2LQhlD16Yagqj1DX7h9nkLG5uiUfRLxYXzorKm+cLTjWLoExqdeD9hKap5HZ1
ptHREQyPZrFFg7RfohrvkyTCbix03w05b2v39nLDdvTYkh8YlNbB9KmfCPJFcNjX
ptPmA6ApmXldUzS5JSO4v8+hsLL3pEfV8MF+TiMJZBM5LXwysEgO0VmTdXQPqc43
d4NoO6m4VNMWRVONhWZM2AyB31By5zbG+k+KXiDMzRd5qLJPECxgkV+LegNBkzuJ
Z5y+eQezdTZFuinr19oYCAVXaYNTPqucFdwvghoum3uiK2+sOawR40LQTRu+getO
UmcjaJ+FJANgwtaRcA0Ty0Hn1mm7OwTzevmHv08pGBEpLVZgr8vRXEeky3l3TRi+
+Lv44VYT9EctEYren//ZIfdSXWsCQTfjU1mIHpizl/hsh8ZCW9wmFluyygdQo/YA
91Dy4EFHoIOc/Er2XNGhqgM9d9yVxy/sYTBcBhCOPAjpdJE9N9/x2ey8nl/5NO9O
LLTsURJC7jy1EUaMnTysWkj7zHAvqMAck27ptqS6UDu+Mw8YzLZfxwwKivquf1h5
KLZMXTSJzBE5PvjHgMrOop0psNt7WWo/UzaP8QMUQnT0nNv60UvKO6aL30lt7fma
lnxKPIN+g7xRyDksG3N8V/kYmml8thygGkhTIuG+BWViO2L72CxRr9f2oKYGzKqY
DvLdzXqhVRb3lo7jLFpWSgwrOU0jUrzspDPUe3AmhP0C/IRcfvuUn4m17d6UWQhs
NDarvip7SvvGabSu5fYEiQ==
`protect END_PROTECTED
