`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xqIIm6fVJKt7m/GHQjBd6tD4PMZPb97XBDPawNiqVsQTRFWRfL4ZCHDMLVNEsrYF
DkE+L9br94Gjpzh3PaocSKCR0I1HieIts/qhw0i6uN5B/beJ9IBb3jPEajHcQB3F
REGs0xbebkN6iBasoN7fjrWhWvaOzhqZCP21yifLTFxfh/vcllUysvpsyjOeWvtl
eh+jN2cdNzBzNWjShkaTpCPjPTXgCJY307Ya9HXW/koMkBr3NwLxUxfi/goEWsdh
GabK1XUzCWlOtp+lFvUEcEpQC3OE2Ef2ts6RWpL8+rBjM1nAXD+hde3DAMDw/zm8
8UkiHnEK2UqIXERQjiK6Ak5h7A/VTEKAtZMMM5+wyFprozT6BDLgcho1XV7JxQbx
rvmwt1jcg31fBUODAQgPDo8xU/B6vGSZx4vTXbdautqJyr5sJUuEbxrcpo0vDsM+
fCVqawe5sHNFOTZwBcC+KBbwJT2XNFeycfis1TImP0nCo3f8PLe70yfYFWAFsjYN
tTzOPT52fYnky4juc2JeTDAlhZztzoTMwVPpAROSaySx4TPyEbWV7INiROXB5yk8
I50C4faFeu4tMD4zjf9ywuglTbxOTOtODHdAw/iBj6Lco8+t0NniNQgaWixlcCt0
GCzSHKja7lvjEz3+tUeOoQx41PKRjpMu8ewSP5E0uoqDaZ3GpxL0fPBmeTC0wPzX
XVZ0I1VqCK01r7nht1e5pX83ya4z5tK7ku5AIo5WKus/XH9yXoH8rbdsGm6JW3j2
sSMRnS7u2O9yK60JggZtjkP+TPet8roXa0gIw3WWjkDZYS7dLIzqh3sh5eG/pmlM
`protect END_PROTECTED
