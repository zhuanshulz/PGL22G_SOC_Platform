`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
874qm+3nSrFXF6NsFupFHW8xBom+lhoYT/g3N1CJkZ6VmwlcH28J/OYDxzYjvlzG
wNopnPubuz39Nbpw+eE/tcre4PuQlsTxNiKJZW9mMmNRO5G8rtgBdGD6FADaWlqe
fmqs6ozit2WEEADx6sjtd21+U81CFIToZlWvjVEik45k1gBRfYaan0SgzIcQiJn1
b39UdcUtfCto9KKV2BPkH6YbPI/EaCTf9uLieMS35ZdGO4EiRE0sNJJjkeVkAb7A
jtigLcT9laqS1cQRkVevvegdjNai7Ua6sXOJRlNs4P2ntV9IxXgzU84GMCyq8gwZ
McuaLes5PBU8fHUcMF57MVLvr+8AQ0snnKEDPuJfGM9ncMCYcXJ94XZgaMRK1Im2
4wvYrLWFpRNUpiNdXec9eFxO+Q97IEiKaLFtnwDH30+/P779h0Tpl07vEJXdq022
l6NCOX76vqymMOpqldyRXVqCc28dz/WGZ44zTo+CU0FYoxSI7zXBhgvxTcZNZkxa
HTmsmypFdTsULE8tV2jmgNY12+Bw9aq8wvjMYTsb1QefGk9bBDUChReaxFRP32t0
YoXVoVM5GSFfDNkBkOh9fXaDZmkMlV8lAM8Mc8wtcYDC+ng3lsQ2bV5w0Zm5eqRB
KZryqfZOIoArCrwFZXJQji6a+3/VBq+wyKMa0j8GgCOq65angfbUVM7Mc2hUICkM
Qm2IJSrORqc1TpyeNpe4kSNKlzdieaySu7fkFNivXZQa+KbUQ2PTlM7RmBTWppLn
ZATjujPmhLeN3EDAr0OLhYUuGOoH139Q9aEhY6kJgJftWu1RZ72cDr/WINpileaE
Tu7UQItxIsePTfOHePYPrpHziELy/meur15u8sapBbZnRnr7QPe/vhM0E43Dt3To
R8AqyKJqZK51/Mqe74hkp0OVltpK1Y/Pu3slmdBREQrfCUR5B2K7BiHc0omGVR1S
LAV5eiDtC2rnVAdmbv4d1zdrzeGOtr4TdL3fKjcoUEkN4dKF010+djsBNZExFGCV
6ECou606O04TJoErQ40mKMdp9AO7GLSJZax3YhpZq7ux6uajALw7zCAXfZX4TSPQ
6hdd26cDthnvu+YuU58VX2y2FOAqa75J3vF/f1GRdMdqMhGC9I3BoO8toFDlFlnJ
GrMnXcoaosEittMBGc96Kd5c3WuUcLUyKgcyZQ7cjQ0tjM7t1KZN5syUWv26mqOz
zAiZDpc8FIqBfnkutj415GVH7A89sWlzSP9KGrDHNEoY2dqMBY5JSNaqnrJPooxR
Tf+G5ZfYkc7S0OZljof29vc+s3yHZCHa6ZyRWJjNayW5bzNOC3R861xEra0COWpm
8Eegkbmd724uXSrvPwRRzGgaiorS0DLg49Cumprq7u/0eP6F5h3rk2Z8couqJo0/
/k6cPDd1odYz2YudbCZqjz3+6DKUT41D84mzhn7r0+pqeZhe8dpCocIiZ4rTIfei
z8cov599+RNMxNPUduVVKkp8LzvWzn4K/vUeSSp2DJ55agQcV4HoKShiAVoAU+Qu
PrNof+EXwgup/QZ+Gd/prvxT48tF6ybQLng7+j2JznuLM+AhFPRG3y3gw3hxMSsB
pE05+DKsA1DW+NzjIqAfCosNc++qK1gPD8NYmTPrw6Fy8zpSeSL2nqpDyw4yxC6d
UEw3LN7PLHZiM9f2YrZac756FL+7BC/n+6rclheJV2hAVe0WeOSU5t0KRZBTPInK
YtTb1670enGGKiEIHusEscq3TqcUV8b1j5rVZshjNIAjgZKtGs3W9nLA2je5jbXC
lTzlrZ7qAlS18yLGpIZd1hn2dTqne2Mj6Ktda+lWtmZvo4nfdnEZCvzOavr9kSf0
AiwdhYdqSBXa2KMQPR2e5BCVH0W/G7+DX6khK1fTmPtQGeEpdmwfA8tZUU1vmBFL
0NrDjcgaftcpViT8pUQkeuuMtBojPsJopfi7u983aUMYAhPvtOZNbJ1qI9r8h3a3
Gk8aCJZgQPXFwuvTJiuO6vcl+ESGXFi8xfttqoKV/lxnppp/m/FCNa+Z/bpOS/hZ
kMBc5cq4i8HQ3klDGDmwj+CQoPPIjQ2tm6kyhKRaY7dmDDYvum9qWQFSvWFiqwOa
MVBoMhxlkMlmxOukFnwpQEulxSHmSu1h7OmV/l56wqJq+soPMMD5wWSSexV0Fl+4
dKFVxGrgWJFT36iIF8c/c6ITwNmSQFpX3dbvdVzjm0hN2eogRyJcAztLZHLU6YYm
UHyMxiZPYgOft3mb1XF8NjPBbga4W2ssBPlJZYtpdeWdv5GotRBW+DG/buvl5qwZ
13JI2spAlbu+eH2kaoLZD0uradfJT28qFWaNgfhr4kjR5SlT9BqK72tPtzDZgr4X
TmQMLtdU6OtX/PXqK1Rns+v2JcAvbme6u+HrI17Kt3Bl0SXSw2muLIPObwpgiH8H
OfFmhlcIoqsEh11a8pTk4DzaeYZZTJyBKJPf8GD33cNLCBAtYr6t7rulLf0ettNw
EtRTDL7B0PVxIIenEfY8fdmE3/4xxXYJTF/b28qvm58w1lKO6bLxVB1OW3TynOGv
nWS8NYicr00UcPZSS7VFGe/AyskCurJZQ3sBdB72OSWFMDCPT/w3Pf1gw9lKE+qI
+kEksN1o19YbVRTLX7IkjdceBzPPzmR7vvTLwF383aNeUnWwhaiKqLPi7rknGQOA
elkoglI+j5oFzEvARzxP3rbuNlSUAjKlzvcvD2IoFAtW9SjCZL+MaEqMoqQi8kUU
jlysss0OBE/VJi48zYCKmwrarLHcBtfWIjQYvvYPebLkHUkj4ZET03QQizYQ/14G
ENkBw+lFYJl9wWKLjJ/Hwkma076Rwyz6WjcM5x1kBmgV2O9N0vZc0uQMyeq3U5oN
EwZc6GATRN+5DEyGdbYcdcMjDeo3qAJroLXQFJuJ73TWW1KdwUToiiksr19woZlp
2hDhwJ4yE0I/Wump2GNXpSAehBGYdV698+LQqP9m5SHLymSJsIU2lSUM1f2UdgIp
nAr7u+OpWmhcBzgQzh+T+o36CS/6Y0iVVRTF8kFYkbbcDYHeIKRjfW2T2UqrJcYk
ofOPBuV+sZXRg6G1W1jHI7daJpuZC+zIuEOg1LE0aBSKgQ5yX//A4n6+6kwEjplQ
BRW3gCfuP5oUaou42m3niUuSTci2Fn/O+Fcb05b9czeAPpp+euD4tUrL08MrArwc
ifBBUQ0FbhB4hDG9nXYWSR0ZxcMnqIHcAg5QaBOZjD6BIshh/XNq9MrKmZjsOhB1
0DIopnKRNi52TzL0VzTyqY8bkQAiBaYvpd4bkobYq6TSefolJgiDSiMW3jZ1tYoo
HH0fVud1Gd0BzjfBf/IMksob/+KOYvBw5a0XBrsN4+jSrJpdbXMuRcMEoBQ56PCD
gZ91srGZGNF3WYAbnhLDvMrMHWAlg/2SS1BqmX9C+WwWYm9rs5Hl/qbvbDsP9yH1
w3LRqsUsG9Pb36m9rIlMsDx2NrRJ3cgzi/N835w/cB1NffAuYOCo5sE0K5AOcw/q
eKqCjNQBEw96EyISf0FRvsFkP8u3W/aU9EyeHjqcWFzXztWdeNyC9pqXkvotts60
PxC/bM1LqZONOqnIGE3NXRg/YxJtjqkH6vS6Wio7yH2ODzmghU17EFcFfb5R4mxY
waW/zxPE/c/dVkAppW0MPJrY6zTHWBi363oeENY8dVtyVuvTJCjL7hPvUDRPL9Sc
PnkGPRIveFYM2XLY4k8xpU8nthrnmFdyRRStp2VVGlnUoziW5g/L/8cK5kWX48+u
i/qIK6FCNBYsYTB0JoJ/B6v7vQZPyW+vF1YwMf0Qab9wmrzFbVfrU4CI/LDZC4s6
SKbEp0F04jBZBWI0yQ2WYuDSCxDIyjZM2LV7TBxkNg+Mhppukl14bim20oa71aQO
1JNi9awStDilW/M05+f6HkInE8LYrlR57JUMgKOKOETXK0ali//o1uUt89s7PPBh
dvLvP3YsrlHoMu5m2Ivdy7K3XcAcF4hDFG0jhPVQ2mMtYFQgoBDGx3O2reZmjAVG
RLVd1DRZfmOirxs+7DpksCLZOn6Zc37j8oA50tucevJu6T7c+oHe8HPzKEMvgG6J
SZbIsrfp/oWJ1v+NxHQZLMKpOTboRW7PVrrGrneEmcF+WFJzhx5ygyPS1HvXvezf
/HB9XlzoDgT5qE0sFO/PsO0HQLtN29tskiPk1+GFC8E3UgBw+j/lm8sePjzIZqpn
sKyzGLlZm7VyrHm5RN1tkPNsdyELzEjfOR2hb4OZgEYxRxS4GNGk9d1A4WO62ijd
cjZPSgCZp/KFS29/P9cvZhQuRk/dZoQeNlOUQVsIZrXlD4VsyhvKhps2wlL9D2My
BQK9vrGi08S4/DwqGdNx906XFGbfyJSM8tusLN3pdMfSsT7S2c9VbjC4fCIveZV4
LOfCkOSmHHr1B5mC0Gvq6PGc4WTx8GKWC5iAJKvOy5oOnQ/DPryJbSWjKRVCLFva
eLVOZaYia9WrAh8FGuqLmORUU+Q69QFSAr9+LSPzTK9UdqlXnDH4kwx6fer1FGBn
QwlerRQoag4IyZ0fzRiQg5fSnTekizl1ZOwuJaPHdMR5KKmwdhwa6kjkwosDwUd2
O0s8QbfkXFhR542WNdypslhG4FPGjIWMbw0YeleDUiOxgtQiBmzuMXUFgnnOp+ck
hA4Htew3G4oYgPzd2wSIbWbbhgwUXCZIo9VdjiMTL5+BhFjgvarsRVgCF5McphHZ
C1T06/H5wxBS7m9HdkeWkhIBKWqgIBTNOTdsMVgf2U2hf0i64G29hoV7zHwVenAt
+iok93RpYPXkHmOB7zdG6VYW7tTsQezn781vUJBxN/MJO7Xn3FonRMtbZzKWzGCq
ancTluafAALqxkKBpbQV44WAadhJAcDfwBGl4OhFM1FrDUPXWNs+PUy3AiocFTKP
YQp8UL3RIJKaUihqlOm2dQYc2NOsTyaXn0OGTSKURW32PVf4KEYwMMGDq7bD612o
U0PlB40BtrQ5Bak2LRQ3QmQQOGyzvsnxniDftcNyBFKDHTq8uwfkepxDBMkUiFa8
VEsuT//vd4pQYY/zCuvSR+WJX7x0Hcuo0dSALvJbrElMof/w+tcMNOALvskE38US
E1UY+MQnJHmwrXDvDXMnZfQ3zm+ZFl6KfgJ/u4g6Sg90tjwGuQsje0oKAhTNWG1u
Z4S4ARpWLbJfeHzU7LzFFLJvEjLYTEhThFKvahy5XlhjC2i7BhFVzIjdNypkUkta
r2Ya5eqGcccrfD2mhex1Qh1J/mdJRqB/WvbWrKHVEUe8FgQu5nuDNPLTixnf1SFg
6LEXrXNo1quEVT4xUXr6wbqCwE7gKh0Xgq3gKBMH5tDqI/drPaNTtdk7vqfb7D6Y
zdGuYSAyIklqKCSVOPB7EmMbHubctQNFeH4gJm4EqR/KDtIIrgCcgOseeWgpLOEA
IYqyniN+sIsJkg0bDnyMvceW1IcOXK/0DPsSXKL0DYVaFOHDgELhmEQvKeP6RgMI
wSRxOY6yXLYzToGzuaYtij0Xxj12IaLCUS1eZFqszrkP2kDzYtwq9T2SRUvIfzZp
Bfi9AzC9Z7StKA4I4JJjV2LlRtA6dn9hdkSAYblqyXZ0u5MOrfcnVrw3hQkB3aLu
C+M/w76xK7tE2S/o+ahaDRWvfLhdyT9883hwCVcvQSOKaVBXAjn5u3yaPbdOVA++
Z1Oy8JsBaIOfOXWJBYCX0R5ZkKly0LkXqKgQITB6V6F63HnzDEfNqOYeyb36rr4L
DqW6wnlacr8G79xxqIpofc9mnnyuEkMMjz5hXhLhocOBxg2iEXGVVmPxwPdSyfto
eu0BHbI/qAnXEfHI72C1AZ16sXo42Xn30HlFJmhKdx3+bb7KjVPOOIwtXUE1VVph
EO5H0PaPAbaeriNAPz1V5WIxGebV/dwekblWl3qOxp19pLqSYpFndUhXA32ggoKn
QEGpjnSNBv9N4tLHokOXV+BT8ed0jbtSthhC7aPBmjx5EP3yHAgc17DLvAd1ms1y
ktsX+uvTvDdubd3dPGbjKFmxuD2sDu39Ms0s0SCherS61fjUO7jWnt4WoQpAh6sa
eDUuPY9wbSlmIRHvJ+S0zBY8IEVJlSFDPXp3fH/We/qV/ruZmRkQt0I5grvajVCw
k/3+C7Den+fHvbhceNbDyctVuzVE+RMXneteB1bLkKND7rPBgYiWhKFfLKu09AZW
f58W6BZEIz2Ie92u1IlQ0oSLQf8wLoUYL2QtGYng2Qs7tYX5WzMoC7VnldNi1d+F
u8WopCL1L1//8dj/n1juChbvvshJ3GfQNWWZzXf4psuh4nGaWmG703RTqSyQtJOi
3V4LxIISD1VWXyi/E37Pfj7yJHWeJJyjNlL//w95imVyiS4Ax+pKndOpglR3FB9K
Utt5QbxmRXRg6Nn7d0iZ1CFoZ28Z6FUpztdniXdhDanFS+qjwY8tgpvV728X6yYW
AUdsE/lkWtyaYEhfEcVSg1yCI5ng4xm8XAiy+DVv7RczkRaE+6+uK/QNQnuIcqew
WHapYgAbkpSNmnOOW04oWDsLi8id4DuNY+knZ5mfTrT1g99dELmrwqP6XBHqQ9ur
vTrgI9LrswsowDPDNC0mIn4x+Au5OVyWSIq5GiahPta+ZztjSKFcJqH1h0wQElYn
GlQEOMlwgpBtGiVia2tazE90FZoT9WykgdogbhuBV1SFoG1lW7ZD/l2r3LpIFeJX
fp7YDriZr1itRv8pzB4xNSSjmRUZ/g/vZ9jFd1MLYIZSwqs0QnFboKV9brcsVbxP
BEHxkxIrn6CQFL+evZbtCXIaRd5MZZNKUWG0M5+HjorrziWH5GTjvvfh/pLkPPAQ
qTcQByGFj2iM9qld68JxVszkXfSp4WQRYTKEgIgW58n0tN7jzUu4k/CMczJz2dCn
64ethjr05COFRKhzHF16mWPJMYAiqKkIhW7toU755rCV/d5OptUAKgPpf5Tf4MAM
K6XQwplbbFBL2/stLvAwC/lkTYdg70MX/QT4JpJvAuuU4jjGJLX3f7J1trahUWdu
edTR4TiB65lGbvKAK4WN93A42DPaDMzLWTy8Hg86grOzw3Tm2qBtIttQI4b5sGBn
lNYVWZ4BAZZKdCTl977qzdv9o0ftGcBlTnxaR1tcFQmZhbueUDwxMMAG03/QAvL3
w5shZHEPHTupaQTpthHhDMs++xQExUIH0N5STEHsU6ytRQ/p4ARL/xBesrFriA4h
ZN2vALQ0COBwTcVCtGJ53icNkqYwAcbQmakIMdjYCnLm5ZWlrw92dkRP7lf2jhmv
Af+bJL9b83BGQjaWWOqr1tGIbtdbRIhfqD3szNG1nt6VzGT9bFxgrJG3ZbLzqgVZ
nlu11NQdFem+LrW24X/uPi93b7AOfv4/ec8GObH2NkBNe6rZRBx3gCpV0BzObC4e
VMfmoVSgKyuKXVarqkAOwojOdrCtZ3hcNb7TH2ceV8HKpMJ3jgupJHBRGiOyzk3v
5tflw4dfCeyggAbJ2mctOYE823LRPaFCO6kIcqQKRMsN2I0AOxzqMOl6LmrG4C2S
5DwupWPJup4NZw8XICkvvBQMP3yVu7AMQ6A+PEh55kFhBPPqG5dYZF9EmauPUnEi
gMbluSHmR01ipH6QpD5RIzPtkWQNqkepRZgany+YdQYsz1fYFfl5fLLrs4RS+D42
QPN70TMYG5JJ7pNqMlVNcE+KAxyiKUCQT0ASS2+/GVYd1QM8sl+K7llf5Sk1tnHI
S0op8d4iN9/0wdkHVRVTxHuXPwQNW4z9kuIVw0cmPHhUJF8nl3mr9NbiIc1+q+l9
61IixLr0jDevbefZHIFP13HkgAGaMTedVzBJywA1jATxM0KNhkvySuExrUKJN/D+
h+hO+aQyp5gqhwVYBpk5xPcDRTeRKUe12ZtNDb8hwk3DtigUSjHwJLoucaIFizxo
fuFSPkzQO+LO/NqsM2WnuQnZJNc7iZ+Ly++zXpJ3aiI4CH74tQ/K6GhgW6wofv0E
8BL7kC0vhZ/PA/Lcrbmjq55PRNMGYcMPF5tlk9+M+g6EGgqqgCvkZncq9mXrrDre
IH/tQPrQxXkVnG6+263tXuy4KkQlxH/JDh2Qj3Zy1KtWEOmr8cwW1ywz2h6h7Gfg
DZhXsP74X7Xdut9sVuPPPcuimOnun7UgMdtkUSjGhLpPgQB5dLHUWCAQs/eYw1F+
LWoEPxsRTvzuhUGERzFjNaAC1jciGPGcQ/XdnNL49OLhy3bIWJZ/xO56rZTSwk2Q
VFQdPtB6/FcuMGMCRNeRm3OiqvTNLtZoECxsVvDdLimS8ft8Yq1vDyUp59Hl1S7E
Js86kyOyciCaDJIxNwPxRuDrYsdp1RdPt3HCWyOz2SQTxyZ3DLqc7zmOYwpDPT8y
NmvAi7XwZ5gwO6ijbLCjxwVQa0hCHkncM9YJ+Lo6VlqslnXDYYZ8N+J2m/kcUf5p
racXseIyE9xNASS5zd8Y9tZgtUVmJibJGmHRyyjcDS7HBerATEiVrHkeNQemH1ay
z6Uu5TSBaDCw712GW3o3W1e5PdEeNy7dzsMd4RmnjjtgFO+X6tdU8pK/V8zD2BBQ
VcLR43V1jeoDFy/OSxk4ThYpqbg6BtzQxzi1z/FtckazrGRBWLsZ/pjx6gRbVKcX
jF7DGhow3hKoffUgR3ukNrR9BNOSKafEkx9U0NWV35mbHWyDg9IKe4dzshlP2lnE
FhWGt9y04FO0h3kiQ4sesiZTW0eJz+ZKhQSQNXGDFYm16cLIF+8iG6/t48BssKMr
whSXEGPKPbHdU/7LmNNHrEpm20rR+zHrG02yrhQ5f2DfLxjkK/jUBsghfZRUqj6Q
JEMigXlhHlDyRzFGilNZ0wUA2Xf6sKnio0knRfEhQUVG+PURwWJTnHQh26WNbok7
olr8jpItzFlnEPjwAQU2qVxo0WKhaliGOTAcHkgr5Dps6g1dHWSm9YEmrXoRKmD7
tld/zzyAaYw8sVsihvxxm+gNiZei/3R1nuVQ17nexJR8jYbe8P+epNqW9eNPWFnT
PmFLLDnu/TaWhTo31Ki//Scur0BDxgiBkYGKlYYWPi4QjdDSeqCHhhba2JLKfkWO
YdVEcXh8R9ykrlLz86P7uQIWd7cxGZF3G+MUOJEfJhE/BREc8DCd4bPMIH7LBMxQ
0h/6kWWUiGRtvLzDCR/xtc1FivAb5VkNFEujdYCOaQ2vesEPp3Np8ZGJsyXu8+6W
hAaoDQ1PDCEZYpKOvnvejE3HzaBt9Zd/TWpQI+LVklS99T26Ah6VFksHEbSwJMCE
vLVP5SDlYNg0dtol9HBoixEvoaN/UqRjBI3S5YR8R8BK+dejC1m5lLO+Bsx2yE2b
Ea8ovlAxIkCgW7nkBIsEQafSg8vjnTHZZXPUBpO1yRtptdwoZcPZ9gb/Hz866ZK9
UPoipPAHVFdwEEghd//985f+P/QduG512CvxFD17uSjhcI6+njxbb8TVqEoAZUFE
nJuyo09XjBjbn1JdWa21Fb9swP34Nqa7Y8jPuBqW7MZ+CwwrrdFGWwBTOUkWqT6o
Mq+w8xhZLPVZoN6fiIgDc9UppkaU5ivwSbhLGIcR8raQy0108dnBWHS0orqvur8K
+iQuqrsqss6mVNbtSUtAkV83uz29zXep2F7XPltKR0I0E+xHQ+UqX2g3XFsR6qpp
3E/kRnvWAUuf+UEE1AfBLY77PZw9HhQ9xOdqjKH0XIEoePwYvG8+/ZDR4jN0Uruw
fXvD2rbJfw3fvgO/i4hf/V4fil+0+0fDHuJsmWUAUA7v/5gJ2y7osRrDJ+ZLGBi4
X/AlLT7Cru+TIpWORJwBy9H3L+R+HAKPStlK4BHGvYRK+XBJpzIMkaJdmkvV1RjW
z4npBhxY7Di2o935hBCsaGFssCnsux+jK47yLkZaz/g7Qk+Lfi7O+FNSjQJWrUJ5
we95HL23LhmC983ESdzOW52fkevCSS2/puRic3nMdlU=
`protect END_PROTECTED
