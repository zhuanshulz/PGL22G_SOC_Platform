`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ABowBMg8stSUOrN6bsrd9wjrwOCTArm072hsKa9qNFXsLBb0qjanRJ1ThuVetVCl
vv4EsI/e4lXPdn4FzmgnsRldE87BjNaoO0ORwyClukli/zT78qAlTmImaRFAJueB
Um2DcmaGx8G+0Hxo/yOxTO/sGp3p8elyelOg+fHU8CLa2BIuvirpsHHxvEJbwe8I
GKotu15o5a1BfBKCwlniMTnvS+p8drbDNvXtXudCYDVE3tCpqOzqMHgZNLTcaDxz
8Fy7NS4bGKqwqv8eFRIQEP2HfIeoXIuS8+jBkRXKjSvSTNuVNqbeNhzML3E9P2dC
+D1HqBdllJMyFuY2YPkVr7xn3PoYSuioltKWuiSUP70mZ05VBfNGiDOkg7hciWk/
vWw6rgjmZraVV9xte4d4NbKtYeJ1DSRCGezDRdaQ99me++Q1ep5zRLPeuuXNfKix
hsZ+xVtOc9m83tAC1MoHUuZkHDJlt2EPJ066hH5nd1fQG1qyptWJIJ29jAwO9/hF
8Zn9asfeA5xTnH0j6wKW4MyLp/YsVD0fhtKlR+T8LBf4ravNtkA+bfmbcvGH4BuK
c8Ecr0M3p1tV/QvaQInlOiwVDISm1qwZOPm/Td8uhqfdx+GPk+hWh/wa+i02p2+y
xkELrHZvxLMJ+9qQ0uU4yPnH6moERg/NOPoOzhUZRJxS876ZbbddsPD2MFjMlnlC
60xgahrc4f0VABVyWYeRJaLG7HNpAC8IFUmcSJ0al2WfhDJThT1OxBMMN6O27O1x
Hq1+KTktP0U5dDt1LUEi3gk/gWm9qwrI2IXUHfov1K7Q05LNyRgXhEt7Rs9la4HW
ZNlMehJJpuVGJvx8IWeGE5PLEUuAfUdVl0q9Nj2826Gijc13jWQaLkedhuAI83u5
hlMfPYJhHWM/phCKFA+vAaLaqEn/wtYVBhzMar8WECfIPyM+D6VQyQPTSNu+6qjd
PTY5hcZNLDF4d0phkmUwzRi2yzrp02B+8MuVR1BH7UBj5HoF0kgjzU44/lAlPgzg
U6P3plKbepGdQJbFbuKfGuNgQ8nftg06DxdmcVBiXmHIobiw1BUklUYkZP+GphCw
54QcA3XZPVvVcSb1tjZAwLIyxOPOIKVtXBfz5itZQZ1Yn2YKYtkdC8UEB8O7cgW7
CdF8KN0GmYjnKIK5thj7TD7olLCMRmolaHQ31crvRGeB3Z+Qer965sqIi3T0Rt6G
9IMEhhXZ6tZuiero5BoY+5o/0YeMfW6gzcmEKSXWcJRKRqLJzDsLYDVom0Ll7B5k
XZWNa7ES5cxQlky1bRC2sysmMGzcVqwrr1zthL274QwVRMJaP7HM2atvnBjIHE3n
HyrtTi/tM8izgC46ox57UY1q2BDa0/60We1S+199va418skfr6toD0mRzh4aiYLQ
eFULRGGtk3s+9Ai4aE0KptSPaQaXNVYELdTUv8OExFbCYv4y4jVAdmck9VIxbGNt
rux++/bFH10TKA+zgiT8NF0ZUpRb+iP9dD/D5ZGfyQ/ZIh6CxooA7yAh0mi5QuFD
tSy5KfwxDga0CKRihS50Ilo4A/i/DNEjK9LP76VvyOq3t92f4AtwUq2T/qmfBYeO
X33YGeUF8s95NvlO0VvifzKPt3cQe549xV4YQC0SzBUg7mFJ7RXBzaTBmtGpPgvS
WbShjXDjvlQXtRVSkvZhEOa1Evlp02CemSogUE3gKmjlhKsqg1dXIkOqHwuwnW2K
rOeaCIc0K4myMgEy7AUpNZzIo8qp7WmSSvAoRCNUtexSbVqXTvpClbGDw/077kPt
++H2WrIYh5r28/NShdNMoNF16So3JO68x64E+jJTdP1JyPx9poemYu8xi1WOQ7h5
l+cF1SLYWbUV6765e9rdZw==
`protect END_PROTECTED
