`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cBkNWtM+PAU8ArNfyotfpzzUgDmyBUiBPdcN1jrzdpUbsyvVtakWYaZXqSpOmoQt
Rlk0YrxgglIpca84ZFlTmvTGV1gArhuqtBqQyuZEciYMEcnREngrs/L3uvCQ45Jh
KbWkUxQew7sdzLOIAAni3j/XG1V6vp5nivo6HPMujFqgs0FokSDM49VbLRSg0Lmi
WT0oqom7tHHq6plRSVE/+qR+SrrUiaU0PrweAWlgxNCxsk3drlfUM7gs56XJis5k
DjjS431c5kZPuSuZLtHeRuymvjnzfBD8ah0rkyYuue7JS0fLDHuUlqneQ3OPBnlh
9nHzVoVA1dw5/BLwroS4xYdTQWEZJ16tSXreCuoerBREIBcqyUTEuIMGPWtInlxo
5pj2mivV9wBgNQO97IQGdbBK0AnIjDvYpgibyTn9qEup5Vfw25nXP0QpMiX4AqG6
/xNpCPi66LScdlb0ZfptKCiYC2vCQtBTJFMXA0PERWbVGIpNnm9EvovROTHE/ki6
bVQ3gdWdpNpkXCOpu2SRrWqV+usFSDmbF2L6+x9wITzj7dMqqb3xJWaFIBED4p8b
Ot54qgoxo9r7+rKuzXDoiyDBWa85rGTlkDIb2ZzlhYdaVTShOA7jC0UprNuVZyFI
2ybqi44KiF75eOnnGTbk2XI7GiECEh3B5Ez0Xa7Q7LaTQhf7TSbT7uhmQTuLlh7X
yceDQYMj5e6kB9OawrjDBF5Ed7mFLPxWQ+zyUvH4R907WulD3Nz3kZ4p1IT1/XY9
3h1ztrrEWNg1zX/FcWmNRYBVKy1NVN5jk15UaBGtGzdo0MD2bh0gEPtKqIdKLKdl
KMW/VDsBSbHr2TZYLFjZAf42hTgJNC8mKxXNOFENQU0dr2Vj5r5DLbsHD/+XUnOH
/VIHGzVurVP4PCITX6nxAoBzkQpribH/LfidHz/M+wxQI/vgWirnc81TwZEOveNL
EwHoFUEoDKZnTiS+ja6tGoGAb4UF7xFFgzz44C7cCxELTUoZNjmCGG4FDpFhlIOG
DebE+bfSGkPh1swz3iy2o3Z2RXmWc4hIN35mGOjTCjJFEluZnkp6tUmqJQf6IKtc
O5Q9MXVCUJJjrIR1V4CdiQ==
`protect END_PROTECTED
