`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZyovKjW4FiJCNi7H3q+C4poLtB7oNuW+sSwmLzXQYvfDShzp5a4K2Qk691j3n36T
UJIkxijPYDtYk2oficTae0c1tqZgGLy9Ff7v4JtVL/2fnDTMdm0q/nhVk1o3OCpU
TV//Y0Z/TWYHy2K87kmNOveqJuVOShj5y8d+3Xk5VoCwU6ateU9PgTWBPaigYPMA
VLKkKhqrGicaa0f87kDIMl+Rn8jck/ajX6sikbbanOnACn2c74XJDkfpr6+6Kz88
tZoonGZKe9zZrntVrn+FdXQ4/VHJau/fuMgcflchaFXEYCMXACSc1R7YtXSb14v6
tcEpyVf+oE35gpHeQKvxLO7G1pquarqzyKZ1ARvXOk37+oUU9+/tFTgvanTYlKpD
oGtpBmL8wdvYNg60Zbtfyke+/OM/vgKF5mqjWAtXqBILoSFbMdsrCkPx39iF/7Yw
lOIG93uY3PVJm5JODJN/UK+Xpri4r6zzdh2O5bGcCjOMpVMnyj+4tnBQWTGj8INP
T6oPwcsTV/dGBVSIfa6bdmeopH9XPrwl8PHRVs4OWDvSS6AwlHIzOdWJT8aYovI3
VlF0ppKZSNQ5UHZbLZAXA6EVp515L+FZYZafn4Qe5VjeqQJQxJxEbERMftEpgvEF
AQggLlhmEbFf5vXLtNiTUYIBzLqlEGQPcvG/mY3Ucax4Olx5ivr3FYXzifJDEoUs
KhpXJYoZ0borQtnWbD/HBzVmwiHZ91y+0OLiOYbt7GBkrUL+AslUEDD5vDDCgRG3
+Xyp9nIY/vm6IBGz02MixHWs48+vyTRXI0ZdC+Apji2HhD5+FJnGTZ+btgYp1QNs
A5qiBcYPXoX8IjcHPuuaukCgHCP+GrYDMHC5RogOm995aRuoj9+II+3nWqf+2ox0
+7LE+d2SmkcNPrydxKDFLaENtY4xLC2mYeJQLAvA5oZvp0Pzs/FA5ay7ewc/ZQSc
W3CjrmMTWOpea4rGjAJ09C/AVYMNcuDi3knL9a0dBqavwrkMlqW1Hr8iaTENMM8D
Qw2KUod/knAodznjXDQi9V7ULV5luYW/yyRO3mLZtsdxJ8NeDHDbQPaGIg5FJugw
sk3Z32N1CZn9eEf1wxvNa5ph2O+q8YDrPlYzkTSioo8Evc54RoULNMx/A/cMsQGz
y7ZZAyKES7zsxXutwlUO0mw5TbpVNsubdisAfjLXhMBMiE+h3/Lbow3Bxt4Fwepe
1f/ZOpbORQBlsior0qCUY2XYUHE9e1+LJ7gf9YhqJYYjNgLfRLlpdhTdoF76jVzr
WcTnNIjV9nAmCmroAl9ksHsOAJOLWRXxfKXISqwE53c=
`protect END_PROTECTED
