`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tSe6HAQK42IdSk6PZ5yH7uIeUAPwmGGkR4xJbLAncu3mrCzDn7O7IycnA15twBLN
zdDOOL5SqCarAIAhGlnu1BJttCHg3Tty7Lj9ZmgY2QIpL91qyYSlGpaGq+VWqmR9
wZGXNzKF/KqLhWP6lKaDC/JaGuR7TV1joSymor7xEcaxXV8fPShuLJuF/TYxLLAY
Bqz39B/F7yz6EeQsQ0OqQRc03gdl+F2uv7XGgl1JDMd9a9/3unEL0c0CnSlG0fNK
HDGbc1RY+mG+Oc845Rn/rQ==
`protect END_PROTECTED
