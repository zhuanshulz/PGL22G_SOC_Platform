`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qd/LXwZx1Nxktdu1Jk7lhK03TjswcZaGLbBoeNzgFdVj5QWOlIHf3srbbxM9o534
5gEqmRh5oJ8rCyOg0e0JdocoQb4i5PYvQx1t419CvUIxa73Sv71yfFKWjP5vQrpW
CWMSuS+IL9Nn1tWchj3qWNo4kHlPZqtF4mzBGkBOpk7AeYFD5uIiZbm+DysHTwu4
VPJcTqKSos9i5rfm4SbEqVQAIvhVdhzdIXDHhdc9i/0LIyBiwm+hGS/C62agWDgs
CD3S1iliwih/vGA6LQ2Owa5OPUOnz6VGWN+zOHV9oL8MXtzx3RB+0Ov5BUvdqgRB
xvZl3parknQvVZHmWy3KgDfA8udTaT+yxrqgtUybS0aIjhNWAKoP7cZoFXM2kS2o
sUxk1S9qUAm6mJXJw+kuX1Z4+KZI1VqMy5ai1bTL7PNIJfLY4dIufzYCJInpWx6P
+6ntf5WQ3YTxCzJZs0dTzxS/vkXU9J4UVBGYqLK5oYtiXeNd4aFF2nCnz9kts70V
OMS3d3h0ec7Y09MH33oJfA==
`protect END_PROTECTED
