`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qYjBblz2OWva/4eN4LfkDT1C8lTV7N7rEUBZxxd8fGyGnyeUOTVekjI93g27XDpR
JoAYb+rj6s0XRu4Mf10jqLFJsHsGn+UaDCOtysmyrNwGT+xYW9OsNhvMiQUsT7VE
UmMZsJ7O8H1D4QX7DHqwWRW0EPygeRjPPrgIMuFuv+Zm9GtXSCcdn7rq4Itmu4Rj
6+Kl1E+Erd1FIovB2skfWpyYWZY6G+5lMwAPlDuzDzdf0t4iRld8wICUqPJG907c
FENC39GUPvscUrzluGM/+woKL7shwACi65+hHO0S9KidYuVyX+YSzj7j14rapczW
LwZD38kuMvGYGIPjs2fM7g8GMfXdiOdz6yie8l2iQyHn8WNTldpzpmAzgj32sMg1
BjlAPFlQerQs+Z6TvMouCwclK7YyJAIvH7X2wR5LS5HcuODknq7GzKSno5kMNPdv
hxyFRcdOt/arN3K9NhTTjK2CM8o/WqmO9+rP0g/44Ji49a892PdwZTxsbbRIj8mx
79pzN9FQCqNqj+j6KuvXkSnq+DpTB8khqZYzPrhdbU+WFXLKI6ksDjEisHdnk54r
`protect END_PROTECTED
