`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R17zVfHd9qQ6F+3RqSRrL8I+Fdzgdi2RDufW9OTvaLtqLhxV3WZ7C/kGbr4BsTLM
LWJkrjB7zx6vTNreBLZQVA2Y9FXl/EMDht9cfmqZsklYrHUrxtnthRyCHt93xCkg
3YabDfnrT5ULJPGHFXBLBf7j2a3nN5I11S/cTdyH7KMAc5+00rcUFrba5EHtoHMK
tOLB+GLwkPfnTWREDoKg4/zCfGNNXZfXdbByuV3jYvrIKbAEIN8YtpNLWNNSFwn5
Jf5Ycupxv9Xf1RhIYhiVxQc6pm/gUpJe20Gvth/f8GEGx5uG7CKIsexw8dD4+ib2
8b7W1XR1wuuiv6aZjr9b0KNslTA+rshyxm6vU1a3Cslh3sfABIxKKtX+62/6y25q
eO14HU0ZRg9Plbk/gbHukYg6IcrH+1x6ov6MzUkhSTwXGm/PkYdHyjbh6UiSydw8
+UkVWN6rV6Z6Vi5nlO7lXwXL6ZUXvtCAWV0zS3kuMBvDJzYejRjEtZPKgExJ+nRI
35x9S/VtVxyncI/jJMWRxxAieRsswXZMhl2TMzSyp4AdVCghfd2RhqrMH//x5/PP
qgCfhwfIs+gay7/cZeqE3SA4tykD3mUEC99J60+QlBTs//ihaykkz20k0HJa5XKz
pP6FVw27BKImzsKWDEul2EzyfoeWmQ4AUnfVEWwUMx9fBHNYb7uclgmKH+qYSkqB
YnAItU47GDTG6PoCQhrBj8DrJ7yoaGtGWyrAlZ6VFf6Wb85c8+G9TG+izNVY4kDr
xWEVulM741bP6/V4YLAGh898UOtA45O8hdhBEpiCIOAp00Dad5W6ewVhpnjPNZPX
KTkJ4zHow9T8P4T1NDR+pnHJ36C9Z9DJ8zU1sm5raXUFKBqLg1w4riWQjU/UVY/y
MWLW4AbuAswPfMJo7FXhbWRe5/X95upcSnAlje/1c1kdC4G16rs5xFhL2q39fucx
gZzt23KDjtQnDnlvXlZbRLigQvHc8doNc8g+KNQQrCt1fIk6uw99+dVud72o9U3v
gBr0jyIxQ86M6I9uW/z5Jw==
`protect END_PROTECTED
