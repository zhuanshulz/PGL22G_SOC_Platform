`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hd+Yfx1ZKsZtMVskM4BNb2B2WlXKx+JLesXwALXqqVdimz6znGsO/hfd0hQHMO0p
SHN6VwFNFjKda+kMFyKVFbDBlIl44s2AQsmHfBzFugnW0zlpZMAHNXJ+Q5c1ebuZ
nEzGqlsoFtVmigVJ0+obPUQDKz6y+0jw4Hgg0MRRMgtZg3DLuKdujEVr/qp1yMdK
ZMbMImv7dxYvt9tV8JyIulgAeWaP1CCDd2u5XsD2wjMSifOwai0uBv4wzAtab+nJ
Az6sZ2YWOESDIXida5TwE1EO1FeDNYpOMG8LhprsOiG3iebdlYL1+n/J6Ro7IdBb
3vFUYhFuXFJOtxnSQ86JfxKA/py8B4qOfUL1nAphAmVu05fl+1M4XPWnvxRWjv4B
uZdgUcXDzeWvthyKSEDLOhrJQMc+IQhVIWiPhqqwY7hmGkGpS5iqHYgh/sP5jwdN
C4aNKahbMX9GsYYrNY1IXGxfxkELMPhGrV8oNDS04Cu9Qg8FMkBq2TWVn5OraFWi
Uit3uqSqWCYR1rMUY9SmArQJZfHiGU108lBawt1+AKuk1Hf3waw/7Ur1ESAbYxok
nxGnPFQ4lZolGg5R4dLwUlsHCIMFmJnO+Bf+hW9uSIcpBGFO4lSbHazWUieWdmE3
lOdCAWna+pjlnpHteJJ0e5p7rlFOaMB8f9zm0DiFIteGoOVY+5oFhRjzgPy9IKSG
plkIiF8MvyOVQwcvnAoLT+NPMHW95D6dK7u/LR12wXmQBt9o4mGZWn1IyennL7yc
pTBobIMmt2H2xqG0+BqprhasDzFyVdbANCS6bo7zDAsVrPfLNeq54rXzFcoYHsEE
dVkUfc/ASpLqol7nn7yX32GPf6nKTnH8Fs1jLjSSOzcQekdKiSiKUoOnmO0IyaOb
iVN42SZIdtloMPRFEHLGNlXoyb2AXt2q8NbktwQ1hvMlcxt3r8IigOTSbw1HG1fk
ahXlrkt9hEH2pJfJ2A8xMIEbcNP40w27EgE/PtTHBAVPMoCLSPYZFo/GVvtbddvc
pFGh16flG2Q1JXlDXtkib9g40DWXgTtiA6TogdBTNKGAFUzHYuiDyPitolJZgKuv
zidDzHvc555WD4TPLrBDctGZGDUIIokuLCwrmk3tCMKgTiQ5jshXWfRNfEXiB1s3
2xkUr4RYHN4Hi+S/a04L5DVwID1/HFMBNleIdxDfNpmYjQaOSqxMFKBFkirUYK25
t5JU5vSGcdBYGwWfjtAG4nh+wzUWqhl/FTWoEzph9CJiwuvWk3HmE/i3mRxIn4sf
wj1h/8Ot+cE/V3/QHfaLS/cKPd1Pp4dtgwDprD7zpjHZxZdJdAwHpLJslnVINuGo
SvjqIRcnX9zncg/cncZnsp6FxNw1rLTWIDVjXqciDU9ozUUptzuN/FS1xHJ/5mWZ
7YUwQUuT7s0pM/E3C+PA6CLBmbkAThc1pn1hvtBGfMR34Y8GKoXV7p3GWiHxZ9vI
QGczzaeNtfRsOUQGWwVng/gekKw10IVbRbx7dH3Srlcnu5OBc5/lPHxEpuQzX651
ix2yXUw5HdT6Xy5v6/p75g+pfArUOSipcteWjoThu2hetsR7A5Mfdd3N5RbWr9DT
c/0XUniyoi6oTmVk0YVUTdOy5XshoWcbDbqFDXCHLEypwQQRcOTn6Pcdfe8Yaf9K
/hfr40CHTEaIyyDVXW1LoaCObNLW0jZzJKW16WwRttdjHQaP0No0GVHTqL0eqIsN
nPxCkDdYo803SVPuDU2mdP48Cu1V08JZwFYVLdBTlaRNxn23pGpuubGjcwN/Q0bt
g12OXTCLXgTz5cUSiS6KLchS+MuMre+1yIlOYaewRvyBKGYQLlUOadhog0vprlsD
8N4f2EI3TQDqi8XNlqQvlPrg4mEPIeVu1qb9JywcjHp4U+q4dW0RHeJ6eMtmofdI
1MQmLFkHxhH8NscVHf28pfNTwutg9h4PYAMY5GwGFyTaQ/+aqSquLQuQUJ3JZndd
ehicXRRVUe7+Q0N8nGFKlma01A/GYnZ6sON104EGs5Qc5dutP9A9zZjOx56l4Qe2
zWbxqxH59IS7QEHWajZoqB5UXEmThsUqxxX89fVG1DqsKqvYBw+FlQnQIrpluuBc
w/RmSjo70kC14HYqhTqE/7m6WLldkpqY57Oo+wHMxtBbnkHcNvk0bGkBGv8Pa9x3
YKOcPLhs/bZHAyqYd/QssRlq5yc392Heo6tmeW2Vn2pTPCp1WK8nRpprfqpNg2Dl
MS3vgT9K20wq3rCn12wtCUoVOw0ZuG8MX3Dm5RFXzYP6KFMH7HDWfB7bKwqeXJPe
HBruiwTmOYZPDnRlm7jD8Z+tB+rDGR7r30XT8Q6vCQszayxb38cOq7ZEE2M5pZzb
094gZuFpzTkgkA6/EDhlJ9SNagMYkeCL5icuxMkwJwX8Z4pR3laOEQdS+pU9JQ8N
pSIrciF8awBjiN3z28jq11ixUOS7xvyrBlC9O/TdZNZ/tnnFCYUuTc5j1UC4+BaY
FVnZDVs9wbjYL8PdtP7exfyV31N+oCbmOMBu1jFvEGOIoI8y9ykLOOocWg6kW9jW
SOhhJqZYGwBB9zYzWB4ZsVRnTQdMn3DNVFGch4D04JXpA3Wvvi57DF7fcY0QzEEu
jtGwOaJpzrLEeh/6MqreNZXOfXYtQW8OmAtIeDwBF5wXoadtH5t0oipW+w+15YoW
09t58K9OdtKiW04I5l/vkDHmjOaQpRIoXp0ilOP6tOY4qjkxp3wiD6p9p3PjipEU
UnfmLnviZCefIM2EfRuritBhKguhr41WkVu1A7pp7ByXlLV7NAXD69qYeiJLxCsn
SyO71zrXbumYFyMkRRWLdhi8Yc2AQQP7cLjNF3TjxUwguFlvKjn5qqcwyU1Hq3sP
DT5mDbm81leXsL+HHoTqfriqX7JaaMHC7rwYDSqnrs60BcwxT1iFqhq2h4PTipxO
KpIn5tGT87sB+rNJO9mH0c6fNaTY1C/fzUtJOvxZKCHt4F2SCxhhDeU0QONtge8h
8f/aWq7qdF09nl5ACZ5gdOG7A5V7bfiuEirT89MeBwMptNzBP2iWymSgZ01fUfEK
qKhJu/lwsT1fC98Z7zQAZoMfWv0xOf3DH/F4M5I0KyfSb2xYpr75Kto/QIOLHfeC
FQBCKultq0AgmzMCQcA3AkALaNmz4WQN84GG3I2LMumJSwjFcY/HIdOOLm5MQVXJ
WzJgV87HwN/Hg/DJUeGCw6wglsHOTwsErPJCBP44tpf60PjrXYDK/uC/j68eK6Tw
cX94+q3yuthMeF6NFClIMjkBxOQcHI7UnYDUnmngYM7s+QEBnwzyaH8TU2DRbct6
PPRavVkdVoyK/8ntqPEqicNIAvSHNwZuhA5PgEjijrOKW5MlsyA5awg6Ef06Fukc
ttCdpCLR++udZQsxuI5Q77iZK3QNFeQJ9P98BMGqFmCBM2D5NnOZqsV5svQSZdoc
k+c7Ef1vu9DWyGLgMTyt4esYIpmFik5C2f3GeuzviriZe6NPccw3bJskNKsBDsZd
lmwa+FD4y5a5ynSDwLgLfRHx3/dkO2v8VmrToIu4AZmbgNA89u13xvjQYLVb5zcv
lhaqkF/qJaCSGlcv+wwaXJA6yIR5YYGvcQzqMAR5HD1p4Vm5glENlg7yyy94f1Bp
qsGXQvTGyJ1TC69+US0t8j0I1rFuSinKiYLmdGMl9CGgIrAQPM2lX4yThj4Cyga4
Anh8rVTP2ATklGMGPAMPFkkiTnr3RwhNXK8jhASdp2tYl3TA+lBaNMlnv4SsC0GT
QXv/g2Lq4WNivTeu8b3rWi5afUfd80tsr6gDF4EEprCAuyP1OhAy1ycfXkVWue9p
XijSHJ+TK0l7BgOK8rzQ2C/Vdk4fXwvcruxgO9RfHt795ofJ1e1OyC58vJahJNRG
WpKs4FrXiWBWoSZzVJRO+T4s7k74hmCf5cHEs/6sFHIwxRcofvZ9eqIGhTjuVWgr
cHfZELe2+itjyYaWWEiu9E4hGfC0Bko+bl9Tkw83ycj6D2Er5BONwp2ErViBXGcl
1/8uX6QVhlyT2ctJz2tsbWylnFNTVvUnjLOnzQq4kpAZpQx/bgIkeKtBd39GUCtf
m8lgGSTs1Lxc59mHCxPmOSimt33xWoWxWqTYxfMUV8lLjZA4Lf+2OpAQf4C0QexT
CPOPcvwnKT5jzGdt31MGwLc7Vyy97dsUIKglbRWehdxwleedtyW307E9scSVQkGx
o9O1eG6iytx91oWiNxMXd5ctH67PstimHACwh6pmgOF8qYfb4DbMC/5WcnvWp8tD
vMKsVF1Gggyx47SO0p0tEXp6x5aFLECKRMnjV6wMCG8=
`protect END_PROTECTED
