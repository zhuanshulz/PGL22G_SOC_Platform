`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iY6rC3mACd6Dej3s2pgMOF8gX4Njtb2QTXX/Y5QIE1OhWQRDYdtWLIBWWHEmbhLo
c+9MwT93Qb+xbuZXBPJ5pG6/TGPe7GyveOewnpF0vZt+gzIszTGBkA3ROB5y08rz
EGgRQepkCWqu3SlyYjzfNnzH45zTBl9UuA572n4Dbqj6puz0KWrTalTrBwdbmjYx
CGp9hdwxDF9bRbhJ63y9BzIH11UrA1FjU+dJj8Bv5RQ3hVbMv2RxG4vt28tj5RSM
8hEohcTrnOxXw3qr6N2+q+ixvwU8t3k0C+bQ0ZsNji52d9ZvnTbZ3FITW4lgOVw6
mCkYL0z4jpc6T1GqXhB5k6IuyvXG7SxpMuH0qUNnZCVz6Ej00xz7pCyBKFpWi3T9
x2UUE95qkm25CXBz2ilL+g==
`protect END_PROTECTED
