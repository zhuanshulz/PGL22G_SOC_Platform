`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3x60378MuZF0uK2u7dZ6ytWfjm5E5+tM5JiMwRAEILzMfWX+staEn5Yiq6XDgjj/
HCBOOHbph/2PET1f8vU6P8A5kCo25RI+as4bQ8s3bn9RlefMVZlaf5cHOdYhlGNN
wc686BlY58+88dxlWkyCXDItLSPa7ocgyBzEhTtymjDUfEbdGYdfGM9ot+TnGZDw
53qb/KpS/AJyrylXMW0IA8IskPxH9OxS4Gfy6Dvg0c3ljKom+n/V8uxfVKyNTYO8
sqik6qbApCg/+nx+BcYR2ig/pdn2skyYWnGZ5zxfPs3g8QjcWc7PxJlwdFqm9bSd
ifdqzpUP8w6wB/Y4aGkfbugrqqp68z3td+3zLUnPDEvfQjHZh8DBhjPVhQzqY3a6
76txy3TyZZ91kiN6sNVpDsUyULbCCJBkA4zJo+uQ1A6DVemWcEp1gp9kKjQybjrx
jV6agIlpaqISHbFytRU2uQjDaVExeZacsfqtIkduB3UBPIKidDDBUzEpr39yDq5N
bm74L1nz20hTZR1MYpaAdIuZ6mQrV21Ffo8hhqLe8liAjYUOwy0H4d2nNRiSE07b
KEgMEFEgsi9/hrf2qVkNxXXqSt05UCfm84PdpK/L3uydEgo6svh8Y+lfN29eKpwD
`protect END_PROTECTED
