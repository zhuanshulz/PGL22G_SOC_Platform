`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A2/9VUDmlKHDpcbGLkOZwN0ZmAGOei1rLMJx/aubCqY4u5dXeC19YahT2O+CxPdl
vD99x7f80jwNmOeOTrH9uIL7rWLEkA2jW5VydLw4PJ+ENLkQ/hgUnWmLcCCcG7at
lOJIQknFTPiJBXOThO2QlX5IJDf9R94Az4qeUNUNOI9k4+S4HIwt2/XS54THcb/4
Deq70tFufJPHwuMKR8+oLXxOs0EtcVlJoNu+8DdhPGq4WPGG7aLXZ3AYej2zFOnC
jtHasXuF+VnD4WeNDYCqNtOW3jNDbAbOc6NBfHch2e9eSoLCkWS2F6IyrwP17X4S
q6UmDlyQ6PrjDoAZgl3HTy5s2D8C8E7eCF4Of6aRIp/sFaD4VYZdanFrxCNmO8+C
oTFN5a4DQXHIRnZRyUPQD7TbVQI9ENDHHMqZsS2qZLXqZJ+hFOXc3CAxDew5Jhhf
4FShCGRjHCzzeqgJX8zlqxLCxj9sgPNAW6vNmoFbs1Ui8eq5Fj7U34cu0/Sm/bUe
CYgknu4W3+Je6DjXZsznhEFvNMJNrkPY4KWAdh6flGtMsDyIO8aibg59qRLc3ghm
+klSeeF+UUsjvYAYFsHZR+JFiovl60rvnIRGQTUI2jqTfMIypjc70nTjwZ38vA/a
4YULlh797pKPSTPOviY6EnWBJTCOvSWjt2s2yNjhxlvaWPtWIhtHVOzy7WzDKKXw
dTEiORSfJiju6qWnMxBMFq4WlF6AiuNVD9qWl4k8LAk6cJiAbk9g8wQGyvf/42Cd
9V33es5w7XlzswB+xt5dVI3TfVOWlOeRXTcqZCNoTPfu72IJXahQJ+qUvCz4qcXm
ZCFTw8AJQtChXmRvOD5WRozwgOQyR2b9WxIKdOgczT5tCpJxj1gkkBAv6tJe2aSr
9HpGXXoC9ptQp3nRE76bJvNw7IbaLCuVs8nx9UYJRSGecZLUJIlUjJIg/BGv/R6y
5ijpM1FdKlVolL9PTsaqZzDdI6eAnQRnajoSfmOxaaZwVnRUV39tiZJMIBeV6Q1/
CcUmNoI5V+DjsffHxLEHucQZyh/je5FF1dYg3uAd5d8iZ/sl9Si7yFC2ouHwX1Ha
BHHSSAHlm2mfcJm0nw+ME/7ZqfpRaXA5iVZ6feoMMmGDW6tqANKPoqbpNTp7Jfyg
cs+Gc5jv6Lm3on741CH17P9ZHD7hy1GSCutOWtnx0oYdNbDQnvyHeV/KV6w4owZW
thrSb1X9LS4ZIeKMuwAMAvJmrZL5NSdOKQT22QSBC0c=
`protect END_PROTECTED
