`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F7rh0orX3/+7orvSzA3fYYU+4zsQZYYipcRaIaIhGd7KA64v0ESLOBJKtXrn2jip
QwdZGFZOtAxOWt8T3t95KEX5PgbchxVJEgeDQYxMty3i1PxhGdz8xKBOG7tj+8Fg
2WuSNpBEZgNQgdFBMv6W41atgnGaX9T2xM2aVCVb6wNC8ha24hBSXPo4biuAG8b5
tnMXEBuhBnKlqyVsveX9+hYc+yw0XoezYxa7nePalvy4k1m1HKrT+Lkj524CEUFd
Jf4K1WJ/3WlnTWZGKwMy7AVhwvfb5MtFPB4qCtk7bXa4vzqaas2hdEU1PfUIFIJM
dPD9YZVIF06lalV6+2yrjMzu5oXMp6GotZuE1At08LL1cY4RXFHvQFtL1b+28JCQ
ala8oF75HLSIfQYJIfTeaogPaHgfhppEkLgUK9zL/eYOhgK1bcRuraq+JlRlOct3
q5u1s4VEqmxAPNN3c2zAreiq4GQeFBll4zAJ23Cx9l2qgIbfxbTD3HXPwP7YIot0
je4HgCaYufijSD6Y9Qrtlma6tClwt5AGOcM3AE7UtYKWROWgdliJzf6TUpwPn0bq
0u0vHCR/IiBiTMI2kCEqssoj9jhrR//dZNKyWafUBaRpgenzr0pA+WFVonOk+ECi
t8jbN2YaImYCSROUg3EqKQdS4JhZGyKTVKnkbubKhjU+ZKEZ8LE3wUz0XGeF5CMn
yflDheK1lIMGhKWoKOxUirs3jrf/UUjrCY7biDLma2Rj/wd8MXZjVPyHvBw6WgsD
hiRoWP+Z8r2lUhrpe3kf7++zyysGuc1OuSl0cjfNWE+B3tZy2ACMySdV43cKYijk
8XOs+zi2xva19SWHobzR2k4d06uf5w00EIvGIttSERDztANB61Vt0LXOdQAGJY5Z
CcZSEOLiRvO7SFn2nhKabRjUItB09zJmg37TZ53xColuq/aULWXmbfZ1G2CNjvnm
TP5fK55S9ssvwyCcnGofn2IMdV69/vbsdnNPbJrHoK3c8POMuQKznvoLN49OqGuV
cE3CpzhwjnROgqj+EYSChWXCBa4YNB/rB/HLlaScBxcrJjrFTlU0CT2QSLCTka+4
/d9UWM8HEKQaGCMnjerU/zDG0pCEHKtEEHnffnQXLVfvJo8dJZn5HuBYAz1r/WVN
0pdwbd6rvoDOVH0mMVzM3r9E27QRqrd4XFZjbtdt8+J6qZtuxzze4kdCqNrUf5n4
iIRXCQRgXjNN32h8WWQ74e4nRi9XYH1Q+OmBBfDL29Crg0ePxYAoTbkmApaeLsj3
FE3a/8gBSk2jt9xnG1uTDiPDe8CkLARnQk+EEq5gP+WM+cIiR2Jdg5FuZ4ul4lVE
GFeGEaTvE3ili0UWJk4zNDL/SBsMztxV+e5NZTnZT5nlcT7VSXaUBqlRQWwfp7er
Q15vRzI7SF+zpcypVjGCFgCGnTpefNg1CHXxauvSjjIyLcLMoDz8AeG7fAi/R9xc
Q3tydClBa5t+POZiK2g8K751gstREHVeb9iClqjfr3ig6ZQCgODtGxCAUOOb0+h4
VRuQQweKWdG3pC4K6vRxaPkvME+972l9Bph0BW68jYRStlz2FkRWQzH2Oxj2k0C2
Srp61VsXFx/9nEQ4On4SzMW4TFVUUOkfJ0tFKgcHyHxD+Q0sXxBsGtyPYlNnEd5v
YsmcqpRGdqDrrztJC4ZMBIE0yxtt0BhIRrKNcua2jTovKzulHs2j468Gk8w75p12
IYAOvQDZCXM3CwynMcvseUztogD/+N9ydXGP13ThidOQ8dRljek4F1NmiD6y4Y/7
HoCqXe81YKyjGVGuGgLPx9L4a8/SlPjDyhiT8GGPATOB17evynhTcBMGlTFAnGYR
OmGGSdwi4SwTxCN7mij5YbqPQMyiQWuofWU/ogGSN5lIdwTXrQUngL5PAFDtV/J7
dYSDIDL5+jzzt5cxi/hZhLPrnXQVEa7pJ+NmmBUxi4fRyemdYTkInz4Z2IiEwZ63
zRAlQ8EU83sY6ilXI8K5zNrwtKKMEFmRvan/9TSzndQOGn6HsUm/8GjlxHDLN9nz
jkIt5SFUxe1f6k5tPrH22r4OJaqpkDJXdm/3zM+lHh2hwarWetsfPGltbd5e4HcP
5tWiinQNzP6W7ZdRa13b9vFZe3WKyEqxJQwRhurW5eCFOufYrwzVJTernCbzYPcS
Wm755EU1DFRKsXp+KQUAQDAJsXvfeV5QCz2BP/phaEN3pfWn3qGfebN5taD70lu9
4YwmI1sCGGX35eE+DFVrRuZ8exbBjA+2WZs5uad97itXaj03c+b37ZoS4rZioVhw
TgCFfDRpnQ/vySsqGyU2xfELQMvs0cdCcEhEYES0VSBc65g55FnJBg7N60xMkeI/
oEJevi9sY6cb/M89k+ILVQxK+T/bfUeKNG56LHhKW+LyAjoi8DXkkksqSC5lfQsX
xMqfer6SHbA97WGGlfjlwbsEzvbWA9Gz3bgRd6p/XaOwcD+5rtG+0LDdJa6a3ZZu
8hjFY62OA8vIbQxoOh69yRN7n6OX6seNH4W9luRIgfNijrMmYa/qlrBvRHuEoaqR
Le6JFT+Us9nKlPMJbfFQZxxeQKmMvq8LTcaQv+kr1S47jw8ovDzeRJ5OA2+6j8nP
LHtcu4dz+KhLHTKxobuYGH675XFGmiYqpAMVWNRrWYiNc07tRDnIO/PZZGnhqfl/
yIq4gVIKiGnnHNEfkwGWwv0uIn3WihOBWqnEI6CcP6gx+QCb+QRth8iywF6lzYqi
ZTvudV8gKvxVsAdL/ZkJ6PB895jdPoBTEqp0H0z6JCSaz4HqKX9yw0z13yX0GIQ+
hR6vZ0LanYiz3Del4B00FYLm0B9pALfS0xIO1R3VBqqoKi6QEdIjElyn2ksEegAW
k1kn56SauZV+clRzqQf5ZtvSCxB/IQcYO5aKIceQcYUolD2yEyepnxMdyDO9UN/k
Sr7eoBsKwvDJ0Gt0eZylY3ykfE4dG5dcP6n6Bhn816ywc82JGWhVEb2+8GmnddkP
kIxTEXP7clCSBuuhPyBbkE29rRFJ7SPh0wHW4LLg8DBzGvEBjPfbAq4PcpgwqpGX
+4GVtan1ybfTUWWFc7QEVu2yv7SpXf9yl4nxMut0Nym4bxAlfszI88PpaThhzD+S
9+ak8MTWsUiybrwa77ekbezMm0Gtm4DaKTqQl8gG2DpxsVahGsheaZ9da7i25iOo
xOpUnTaMY5fIYcEQAPe+vLfEK2saMGQK4n9vfUeOxFeOJCA4k+uYgvNcA5CHqPKA
g3Irk3WnPo8vzlug2Nq8PBkk4lTm47JESNGwrt2quI0V8fTjXhPPmOWLIGLVmvY9
ntZx1NMCR5Nd0N5g3Ll9c26MEpVTXA+J5VbDWs4CZjNQlOqJP6g6EZ6zBSc0x9t4
He1L/8k+Z7EFVHvQUSo+H+iXjc+nMWpIYFklqO2zmSiWQRKubdWwtyDGIZlj4o2N
rBoe7SkVLlKbi571Bg6bqRP1Bxmgt0MPZgkmiV9T9nN0hvg9fnnotfz9I8OOAX5r
1AOh14M+wk5j9EN1Lr851c9Ub4ieR71dPrxtCs/Ddwt1iRsKXkM6qsQt1sBrXMqR
jIt2yVSMwqYU53m0owwKT/5DnHOdABwJhKeO6Q9uzjTaTkcTYzX7j/It/PS1tUbt
ZF7rm2ktWqKm5EMAppzXue5iMDylwFIa810eGA8rYn8K3ApvoEhVJ33MMRMcQaZo
9jdwfBRdMwis4DOWmRySwhLqR0wcNTUOTp97NOneqHg4Y85eyYK09tn78ox9ZtcT
cbBrgHvi9GJ/36lavbkseL85Ic4G3aelDTPC9HTHtWkUgEJ8hZjfAFOk43gnigam
aiXcU4MsI55fDvqQXm4po0Z7X4HcGDpEw34/0UXrYF0ckeh/8oC4mH0aOkm6xZPC
3VseaRB7QFdMXl1iYgTlWyPILjwXRkQ8D+vTy1tUf3nFa8/5UeZn7DD8Ik21aZ8g
VFRuyFkKaasbDaeCJ0xJjeQW/Kuf/+1lFYIUqYZDQRXzbYm7EudHxw0LqyJAGyA+
dVDZa4utu9RWW6nWNaaET0b9SKEZPZhFWOxxIHOztrbbL3YmutLHqzTx+vxCpSa+
HzsES0OD4/O6s+IIitjWbvhY5y+hcP2bcAKRwhRnrH0ozDLRyzO9ICLtzH9DmCmQ
z2tAdI9v95slqggTs2EVLIcY0NuQvajvue0VmA7PaWoQ7ZKxLesKn0rmLI67Fktu
wZykbRg1jzNKN6GcbHLsANzwhkmi0OVIm7IrZRIe7j9m7l3BBZf/X/nGuxqkfHB4
ntGfSxdyxBBOGwh/808PqfBZYAvetErxa8mwVLfbM0lFQI93c2qzvaYYs3tkABNk
fVTpqrn9HD6iU2Ayzql7DXdrUBxjFm9QLISbrKJvVXj8Kj+MgOM/EuItd0FSms73
zdPAcjVxhaow4Mfx7SKEQKSXenQE/+OuzEO5BNWnXVWaq/rtsjatdw3MrA+TP39Q
0yn9PFTerOQfWDnrJKc2ex2773uDOpsOWD4pj/rbG+mrEBcIJF5nGUcke0jPsJD+
q++7LfylK/mWLjhwXVV58QpZVbZt468hzD69YJNHZnWSdtr3IzD19T0Y0oFNqb61
hWLYCINBuIW+OBrWRKzrKp/ssWNJBQzFgfl4MfMFmRDsiAZi9ysTBhJesfn6dBE3
MYED3aCK3ZoVllALioJd/X5n1dddDM3VikmMUf5eJXneu4crK9UfFkSXx+JlDc5T
zF4NW6Go6zZIJ3sDSaW3G0BWrOS1nCAnCQ1YBgszCmeB0zbWxy4c5+KUDcclQaRv
KfCESND9gea/8SrDdJjiF3+huhGiHa6muysX+RD9MGfPUE7RoRNvBSgUBhonFFha
jhKHGCFUNFR9IT6+3Gq33UVDoq1ChpbfOXwobqXjC3x5Va3irNlwv4iiFjLV+TO+
iieubQ+Rj8ml46RLrugs4p1Ngh59G3ngt/sKYmsI0/RdvehohhcNrGpl/YIgMhlk
I4zIRB+XvIlBMl5X+eHTbY3LFGeUyzGLqtqWJM6S6GgmgfongX6xR63wwjWdJbUr
UcaRXHuaoYqSEjEt/2Y23l3DRyf3xZYzOx3/eNXq5LfsFps/5v69quxqLNIyks2g
6SG7ttC0W3Y1rIAOkE6fFxlLwSJjuZrfeXl9gCs8iBUpuP1Xs2HcBfaydCRnGTFF
1nGqcIIlfF8mRSDsmF+B4T7MqAHhymZsdW9s+bH1/VxcrU3RKaOGJ+VlJU0976YM
26oJYk+DN7mHUZngeT9JAg7HgzxplPAltJw906IGFJ+fNOqP+HPQv/XYMAC3VBnC
YV0ONIydmQjk7JcD6mF3QGoPUITGIuYq/M+BZyIqdQv8A2Y/F3IwrGJ8Cw1b1Nfk
AN3WeOofrfyBE7cMoNt/R/gAik47997dig15S4njF69+Xn0Jzva5B/Y/MT49mhDV
QZ+GGChp1iReTowFV/EUUdNeuc9tnVi2W5IO1dp+eqT4bQ3efvO/g4nKiRcw565b
kXT81Ahv48CTpd9yLBVUzSfIAl03NfU1EPyxWhZOE2T19Qn1z7w4aj8kgeRmr1QF
BzxayHhIDmHX8DPM6epYRSxXKp/bGxO/S1tt5mCqjKCXUwqiYCrwUo8HVM/PEp0w
kqOmVpBIEXH0YxWGw8iUoNsbVPoykqw8Z2A0qgfMOPHQjGa3camrvB3yJu3yCTU7
IxN0nj2jaef9luem71FSBH+6r9+ngISZ+r5fHVJQQ/FDeQWtOJzajG0WIh7FUBFb
CGlRcTEgJ+Zcao7Ho07rS60DxfGL0DERFNSbCpr8SW2fPbycwXGtnZE1HtA3cMht
0z/TsNzkrBG94npfdt/J6AfIZua8ZLXlIkEA//+InMyd/sn4Lcarwdg6jgxrO4UT
1HX6CiTK+VCFpCSnlsuXb22j9sQg2lhF/64Kcoyxb29ccElpBf+8ulPMUlq3m7RR
NgF1tbz1XlwpkXY5mkSJqf0XMXKlOT90bAEkIjaKsv4vlGxR8kO3lcy+h4Z1lfco
DRDauJlwuBiERz8tWFguIKx8llahWEca87N+jFjExg5gHWwWjbF2w9cxdO3bq4ZI
zt+douYOSLZ36TH0qteMu5Zq0NR8l2Xwj4BTcNxONO5/X5eH2yrb/2L6ZghX0w8I
Ri3P/vztaP4J3wS+NoCBS0bKyRh1K1ezdVoGDMxBZTu377Zpvtl6GTJAw5c/M3Uw
`protect END_PROTECTED
