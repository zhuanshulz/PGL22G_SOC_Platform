`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DDmwcdnCPug9QwPyudtYqYqoJvxO31sc1N5fU6eEcFHhkcUN6OszY5HBTyx1Ji1s
vgoWb7jZJjGceANmvfohZCci4LmeRSwR2apYoRsSeZBTRRol31zr098WmO2PFL7c
VjWO0txtxQ8UawsFZv/sGcHsDEJRtJIXthZON4M4cT9/tIov1BqqpFhPbWZ7VA8/
ZQ308cufemqf7/Dk14dfl3znNf8lIUnOI0tBgh+z9S0sEA9xzOrRGVzY/DvsIC5x
0ptMPB7yxE7LSnXkXXilIFTlUorygsaDpNL93r++JYf2yt7zDRM95jdaFsPWElaE
lBmzBQtU1sXTY0YU6+KGi0ZnyY1aIjihZaeapuQNsysE6M1W6tRTaKn0+91MMuyL
M+/Ftl7RGsVudAPCI0GTJPIMFpvHBhuu+v3irvmnl24Qvdi4tk8d52/uis3BOqO5
TP/93EdbE2w0DhenbKnPCwrBjOUTD2p69yOfClS1e/5GTN2PVflS+fVlfWiu6aia
oDDkwLo4H/VnE7pwH+ueAdlrwXhE1Rk3YAqq2ZPJceVzl8vDNUviwfxzTZYf58DR
rzM5vwgz6iOTvqvgwscERRwhvI0VlloI1u/Ib0hs+qBB2h+noYiIsq7uLjb1/IYz
Kr+8gfY4YkgUxEV3EkRgrHzwP4UVJyDPcP1qf4rKe0AyMdapVnyar69f4S+gdNWg
I4Lw+d9UIfsWSC/CjryEBYgYU8sN21L2jeO3GD3U2jvDiTIquQ7QG2TOz13dPIo1
buknL+EplsVrAdWzjw3cihO4XFMyGXS4rBWh8n07hfHL7Nr8AJwF2uCeZgVfwmmv
DgucwztmcXbWx1GpuEIhXf3SL1Yv0MbjWErdgk9knqrOF9KWrTZoUK9ixWlEMJR2
LSTBPNjBw3KiETvsrjiZDummB91ob1hf8pj+z65pMIKQMCyKNHaMORT7twU4aSLU
QKbSTyD1BN5Wnm5/tqsKL2HnK6yFUEyP+eO+P9KnnGn74gG9JwdbvXW38/CHskk9
PezwDGZcLmy2nPnOjwLJ+5N64UKFl+1WyaiyVL46gQNqHx4kYK6u9eWWMtnfwF3/
1/QXbemAnQAWE4mERF8/6Qye+gsHwz++KPlgBQ4bKuUfJHobKVpd2t9vrL0j10cu
KJ72d8Um+sdRz4qVwp0g4yRIAH6Ml+aSbKsELvrX+EI9xY11E2J83L1W0hwZLXmk
FOdO0bDxAZMPXTvYTPbEwsoO+0mgZiZW8LBBbpJh5eP+Zu3khX7fKza+boLBsaa3
Iv4Zawl/tJeL0pIa6fLJTnomLizaMmEM7I/00t6OR82pgE7/SpwxmS7W/+gjtNYK
g+FzCIs+/FXV4+POn11297cOpcoiYH9gZRGL1JrZ3dCwpntbfq/REoyEln67bPD+
jU/+oxPEPC3KfVtov3Uf3MepkZ8HuQncHal9mwq7bh33EJwKNosAzXUn91McC8zZ
qQVUyD2iIBm3SZjXD2BfZUj7eHihvGH254xbQYavfLbHLt5mAB0hvyuO2E17jDqR
qFjPrvgRAFfKdQ23Qg/1SPUzcCaaa4ax4Zu7TTiJ4QorCV4SqO5uzGDakheaVlpd
6MbO8BzyXkRBQRs8ni9FG878UXxHto5TwOnj6K4OO2Le3GAoBf9Yqj5INYOkb7RN
x5TNALtnxweijg8lYCCYlp0O2lJ3DTSk+7shUuPy0wRy6SFv0iq1Itn2osBsuZZv
L646E5rPsQVcLqICBAcsOpo9UtP/MOShMcqd8Ffpl48KpvZl63IlkfKxRsPG2i7L
ltAZGkAtbEMFPM4jshx6UxNGj21GEXJDugPuuZbdmWp/SdYysdusAvwRJbg+/LN0
YzZa8njnvFxx51IarvdMY8DHq92WhqI+Pncttl2ulwESzQ4jow4TrGMmb9uAbtm5
vaNEYfuQg90ooQtCVnBo98bUASYnIYd3kYqIpmyA8nhP98njl/iZ6he2RUYWHLTY
nSKtyrdtsMtufGkmp3Vbm6t0/CiAdGB/jZXgtksFA8Dw8ZZTk7/3oi9+XJkh4ZhP
VzheSoy7ZUI4CczDxamKOBHogsCzeQW2wLmU60rmtby+UzyFptX+SOBRNoz9fNgD
uthhoEnPe+AysYaR0krROWkluYw5elwUh9Vfyd44Maf0b+wxk2EiQ8TBxgQDMbGW
felZwRyKi/yb8swg1PCrxAwqfCUmUtOXlpUklDWC2mlJ41e3S7f4YL1EAohObQjq
T19eN1ZaiemC5LW41fZkORz6m5w6aKPIHfyeOwpMzEPDjQ0/9c345UpXhnjkIL/L
JeYHocSr+kdSGJY9jiIVpnkXJX/GN76WTp+PW03nieacQNvb+40s7fPZzKCN0LUh
j6V9m0fjaPrcpb+FufCWcZyQSMi5SyQkx/Kt0dVEJa5rdw9YdIN7NGP0UoBLZvHW
Xt3JjbQCT9IhLvwqMPosidgfnzFYbRyr7QNfHPTpUeHg0QMiDDfQNBUwGb6YTWRq
eibrYS1wbRpYrqzDSY4qjl9t1hw4zWM2SkNoDFFdDzMHv9wLvkSEq/GqpGYeqOrz
BsH2SaQgWIWccjtI1bSYR3SFsxCALwfQata9OmN0ISjbDbdI/oMIcI5Rsf+paf6w
yIgr2dUFHTjTJ9L6hlJhCSPR6B+WXjLNM9k28lXAQTObRqihsaJrF3PGwd25VBEc
YgCO0LVUPTf8euSTKyY3aUTwtak48LZonCgrrnTQae8ZpZAKEERMfjlDAzis1kgA
R2xS2nu+Ixuet0AvVGqsHbT5vE0a2Dkm4Xy3Ye+AQ1S5TOe+bn2UDcRsvgY2kh+z
j5P0WQbabpwJXDLdNN9CJv+8YFsdCtC5M803DWJkeVzSRaAPHnlgPT5LFQsJd6Eb
N/mm4jrrHPIuhq13mntF8raiXL2Lk8377IXvbj079zDBkK27J/RAtO8jxI2ZbFwh
pMZ053RGzUrO4vC7TDXgI5G7NRxBPkcws/oCvJHuWF3PTXzD4jHWvb/16ySflhU2
q/5PYKu8oGPgMeUy5Zzef9zOKuuobM+eoKLDbSiUqhAPoiWd9XsnJL1AdcY6L8IO
0Xei58SOKbnT9y+UUpnpbgtakcfoAfwp05sWDotOFcgCe8dLqmSW0xbDW0bRtrWR
bK2IJjwZMwswgPGAN5S3on84rGMZkKIeflGTk8cD0LKBpwr8DkGrWh27BCLnvzeo
oqXDXlh3p9X7OZo6tNumlMkL9FKl59b3U5HxgRgCqnUWJAzejU6lgkoEBoEGhqL9
/xh+fOYvRXI2snA79NTlzMh+svQ4SF+cPLEvHg7j86dSjZtcQLVD9V+4D9SQfxcA
m92NnWJGAWejQr7zHg2Oj0vzgPSLflU9xvaOwCxvxT3dozkHKPBpCByxUSVFKQaa
UspQLHkyD7Npqx8+fOBoDfa/YIFR8avIHS74nxqIuDYUwL98hny2FF+07Rpn8W92
C0CdvfJ1bfJX6S4y8JjzOfiQAWM+/8D2YAjihC99wR8q41l7YnUjUx9vYeSHUdwR
GQV01fs/ggDy3uASY1O/V0apndvSTvJGJGXtvIe1hTwb4OZfw3eurmMfiuHr1xsO
GTnazuveBC4HkjoFHfX8zJhvxQo/0HDZp521KI3Dv5kJhVjy4+uOPr0Stu7NG5iv
ShBXFmWbNe2WzfdwYMPbs7MAk7O3krLct5tHkwkNILSd8OUOmSCmanuAgDTZ4kCa
QdOWcoJskA3U+nTN/EOjWDd2dDuCg4/9vyaL/p7UU5O5hzxo8Gifh9uwHu5qJ2Z7
iivEY2REvAbVwWpmDBuekQoj9clJamrEC5+Wd+bD2Dpmq9UWDumig4LvL2KH+kO1
/SMoE90E/NrRmvzNcaIavlTXQysIZ01Vxji4FV54wrqNwCsoxgAZaf2UBT8uBHPF
lxPfjpvd7X+t6tHIR15EEetvtInA2aWCMnki3/5KnIXeuUKVWzj0DhSIYdyi3Aye
E0U7Yf/uYOugCbbbCPkcuXDlL4vLKjzm5b8ggpnB6ciqOVWxwszjdidcx0j4B/g9
hjxRQemJDCTt9QTRpRmsMTRJQG/+oPIek7ZiLOXPiN3fMxRuemqqmMf5074Cu+Nj
XBVIPnc8o179B1tzdIjS/BDTRiqDjwedcF4EzGKZV1tzO6Q6+ndDcsxEXRbFVaRT
+I789TTLrprurlB2Sqzt3bbhfkoa4R69XrTj+KKq9TTfRclS6ZxeKbF34mPsC3/G
ZMZiYh+0zSPGlCoy8bNTClSLvvdFiAFssSyayxcI+gFN2NC71U1fu/Iz/ChT14D8
SbEnEdWjPIWrRD+B8JTutFXPlCEigNQQ3l9Y4rzOR7wjjd1YWtRxxXsNY2HTwf6q
YY4AzoLMKKA6j/PaAILBIA5UTLEg1Br4LGG7gEsKnTs4+HCy+WLoVTUXQq0hFHpv
qgLZ5fu7o766bOqJphNSPfrSKRSrQS0J1RmkEGEa/G9Fy7cT1LQvTlxaOE4mGM0/
ORTTKZ4qeBHssDYdHwLLbS8gXACnJEL6bPWb3R3d2OEU1jg9er5xlT6mGzyUKmHd
yNH4UPAl8DX/PPDlZHud5KmKOGsqFOUB0D6P+Au6ijk1s0G94JYjREsJaVbogcYX
WwDAn3as7DeXPMHWHM5bRL5nQ7eRR6SijXfmOn8aVE4W/NuaOKTd5ivHf1qZM7yZ
IvYSmZIUnS9uq9C0JEMA2kUktmnUEF6V//abirEU/wSfPU8+CyICN2LqNgxF4XsJ
e3Q/3dLcK9PBZbWPjy6AsAVsaQhk6kYlMVYDSgNBKjRkqZHYeXkBY7ypERdJ1JO3
dch5Kppz9BMeDkHiDQUOG4Is16HLjdlMx7aIqEly0c4YAKoqcVOMjWtFayLELm4q
4qmFEn82Jfv1bUMLHOjFxY9OXfb4v5MU9IDafvBU5cWdjKxURDZIqNCdXt/Pek2L
XiQzDsjgmHdTqC5WzXNoPRx65NOMucPNy5qR67LHYYZhHCZOX4gXUL8H1KNvykaF
U6tMWDBUmGBY4SpwKovl4IIpyb6NiYfsMhsQe8lR+NNZsZ6JEPYnyle74RbCZk4D
tYqrf6KWj+SThkJg2KPIUtTTbNuS2VYVWZeiSX4Gps1LhdIfemRfjCpIZ+k/WC6i
WTQ5Ul2CULDCu2eMb0oNbvtNc1BeppGJt3AK3jlLEDTnA1iJIV4kAw74I9itwx+K
NQSfq2Zxi4krbgdxxAA+4crCmMWQYXWcsY18F+b7D+D0EXI84+XEytTB12y4+L4w
M8O0QQS7SqpYGXz4nWM6+R0HUpg/bKJe5fNNgw/wgMFuClSXqUb4Ld3U6SK/2rr5
NWxb6EtcPyREwFy5IKMapeO2JVAl+uJAJ3uO5/7Z7I5FuPfDsyJC7lC9vxpQBugN
0ciIMGc3632Gr/xULr2hesy+P+Rq5Qoze5b4DEp/PAgnTiC7YRIgWMosBDOW/Pc5
ABiLMb4gU9LWNwEaLAQQpStJirXdfLxxZ8Y5w75mzETVZhFfKF5p5zGhSFFxs36+
nxyQuekZMwoTnMs0sI4vBs2xWUMkR+fKK9Q6s2Loo9Kx7Sw5YiaANamkt0/uZsk6
i5pBLGTs5txhhvXHmqBe+CriS0kd7+t66W2C0ZeqkA6EE+tZEoSCDJeccfmmwho8
uubYWByLdGahWe6Jbw4TP5QrTckz4TSVaeBnDIq99nvLqnFi46beUB1g7hJYIIfL
8lBuG5toKXJB40yEr/+iytyggDOCU4SXSbVlQniZMf++N/ZHpe9KbtKQ6kVk7qRD
WU7d0cooPyFX6m0GHC9QQZ5Xdh/VIKkiwOMU1S8yMieqS8baGPdTsEhwNPfc5AVL
7ZKvM7T7DXGAdgrkbPu3vHUUR4lfe8+XAcw19FJOj2A924UMdXHKn4v38udhpFl5
VaQwtRyzmc5PPjJvzQevXXfpOQNh6u2TfmqlfAEiTbbf5+mdw5a2VFeeof6jk0F/
BrgYLLh5I0rsV21eNv8/nRfix53h5dAglfeNFdhdSmdmH34nq7IXI7VYSrRsDyRF
wCX6deQnuoINBAtdkIynZAHSDX9MhqMVXWCT3b25rF/cucc7eDWA//z0Z+UcBsCr
VAG33LDbSB3n6r3INIoVf1q8K7ejOUssj3cVaAukPbiuXLmZBKihu606KBEd1l5G
wzjXwKw/O2G0hsqVVdA38xN5F0RvLiFNflRJs9Ho9a1YT9p+qfxbPe2opWEYV+tn
it66WzdHVOeaL13N1D7a2kcATZ9CFQyqKtxLqvZxadHscSTDMT2uVwGIXmeJCQvH
L+cZnuDQAQa1sv2oXYlBnzpXH8D7pUCdO2srIPoFRJzYVChp1lPn189WQejZywtV
cVteqstJ9LgyHv91mNNPwud+shQ3RTovyXqkbNPzOvOX4VsN/z0PNkQlaUxTsDZn
3HjENRZ+oKc7ZutYW5l9MLXw7c29jDFdQ3M9oJpC09bMKx/F/8cisg449A0+IiG5
sNHyrv3OJoL14VclUPtwZyARbC777elaTC63w1iyHqSt8P2QM01SjrdJ6zp8eVUo
R1tQJoX5CEIDSGBvFMIggGNZCoPl5GrEymlWYblNUoDl9pqVFmFoiQECj9Pot5Ds
SfyIezO0P6ln40C28c/ssa1I9wPhe9H8Pzjj01lKyfWZPfolPv9uXKPH5SB0QGKX
p6wQMJi8KGD/hHkt1VsM+cg89on3F4zN7+vrW7u8VDzmmyVCiXp87tYWe/8lk+6e
nejFZhvlp2kbZFGgSrx05TdWPy0edHELjFl2bey22Mw4IJclbCqhaOg3c1hZZyCJ
S7Qx8pszJODBAhU4v3ZHisMl0hUa6ZMJPAlIyh/Oc0a7AFPVbmsJwYB6k3UYUA+y
VB+T7d3JI+SpG/UKqxaosF8dMaOK5cV0jtYe2Q0gSMefjdcoMwldxVYR75aDUZ4l
uvOh2B9rwqsGig3DGLa4zevUutb3rv2qSDHud6yR3hGgVcKmCzlBRChKGLsAaoTX
CUSRdl4vWxGFcv4yaSqc0bbPfLht9cpz+mNj8Ujh7QOKpeLCj+sgV2/95bIbCKPU
n3HXFf5Bljx5/a5ewzSUscPznOw0Z6BFDMb2c1ywhzcS8u5TT7pI5f2ZYiNv+XIp
XjpbsjoZzuXQ+vRYWT21zcKY3wvMd+ko4o3LOvg/l1lrbeP1RCu3P7cMo+skwOGN
ICudtlXV2KYerzR3bO4/4vy+QWmvhO2/M7p+aHxNwR9k/Tq1K1oQBedBGuLaz3nj
nzLYwxy3768I1pTGX9n4aPZusP0ngaFDNgsXKKz1aFJy1j/ksnIWmXe2KmcBHfJR
MkO1ig5uOkfPyZIVBk9hwTRB+xoAIS6cQZiB4BbMBqx+P6q/Qgk2uPtx3S7kwtXQ
PorN9uwKfRagWSmLJMYhVct5cm6Oan+xyfQ3yBIZ4ME7pEKsAJuTWyynCn/gt4jS
bppuxRhs9HwtHtfhK4iS1shFsE8Yvu9RmoJfwdHgnSqWi3q8DnUfWvi2ypD75l8A
FzIpCVwJj58lVlFA5bcpe8Ssf8+2ncDH83CZgD4I6t5li9WaFvnQnL7mlzDCDj8m
8Ph04/Xur973bzUl6HDtIdMDOowNHAJJnBemTCS67af8+xFPC3/CajK2D2CNvHQj
m7Ko9lb2CIby+cvgWGYO51HB67PDFIK/Pl1V+jpbe10YO1s2QKO7NkH0vxdqmGHJ
t72l116g9FHp2m+x7SBAzH1bFqRcI6aNWKi9/dfS06BCMu4UN9XRxMZjNiOSmh8z
PqTvw/6bWeMvnce7nTVtZzgPYakTcnSPj97iEjrFaDZZZLeUEHUzckvZ6iQsyGHX
ggSrYB4Wcdjy79t668Ioj75vz4std1ofZ6QrKxEODWx1PBQwJiItfOBasPXtQDrT
0dM95nRNC744GZLnHvICIwu48a2WWt5aQR9XvcqTrDgquqBsDXzKpq0IoBVNcjYF
EepykegVsPR5LRWYN8XTCyJLhJC9Rdg5BkkW/+ya7Pml+l2F6oKl/EnGIiusamVT
9y90kh9UiDwnBYmvE1d4pajg2RLMUmS5JX194PkdAfHzjwMQJU0iEg1IleHGE+2J
gj8IiJPcxsMC3XTRA24laaJK722hDslO2EPBAx74Uzmc+OKsZbvrb+mWTzrMdHlS
CK6/8wbY70RAMbwdqZhPIKloLk0qRHReqTrtKHIZy0LDXMOhnYII4drDKjNKzfd1
AYDFHSyWKNX9T76D+IzhXPkpkWO5kfiDk0nSYy5MxJq5GYLR1sPYC0XVTeBoqPak
xDraJFyG3QZlGiI45k7yP2/nyPIvcroqndexpLmQSWXqO15xSvIxh7pSsjRAJFOx
yGqiMpFMRYFbTG5+kO3SjXRlSsi+lIYidWPI5LHHIzyC5T72fLQr/wK89rrghpo8
850m09UXNUo8tM8jSvoKJIcgh+jjx32Gt85GK8qCmLNVXVVgXhrRhhoD4InpWnLI
BEzyQxMQEAde4+LsLOpjBZqbSE0pi85/fj0qz8u2UkOToTJTufqE0kNnpM5ei+O6
R54JeXsLCKC6ulKkXnumBpVzHFNJN+gt+0yfI8++aNh1+UT8CF1kn4VXC1YNK2KH
9Mxpgf7FViq/icC1g9f+FFHvkXU9UElf5qhefYLHZdWwSZPsPrlXVvIoe3a+gITO
fj9N8IQcr6IyIbq4+nfH7w9vxyJIonLZttUrrTVhWtaSFD+Fzt0j/WcG91no+RoC
5g51CIABfJznC7goev0s8krLOAYxJl4kVc5AMd3ipsE7NRPlrW5HDNv0MCTdEY0d
KmOzA6tF81YnxroeHwAZMVhfHBIzdyc0NsFheNG6Es8ddY6UbkLV25rHHfDdHUQr
4bcomJeK+tuSyLAAAlHtUI5rqPb1YVzFXNy+/ghz/db3Q2Sb4UrJBNP2BnKDKSli
GP6TU7lTiLT7MxbBE61WrHbQ5HXBwiAew6i7sQ3qNJX8PA1MvsjHvz2g3oObI9Vv
3ldx8G0GylUG9h0u9/DRRzk0IW0in9IajxdMLkGS2xScZjxAGAO1NPg0hWlUWCS4
x4NSGxABU1tNZwbiPnMO5zPQAQHbcwux32WXsQp6OiUU8AJgROcpN1iJZEF7GKme
l7729fnY2Rh3TaDJarokOij6XI+l2qUTvU5MJvAwScKDCGYGO6tVlotDFSfiWgMn
ptn/0y1AaiBOFk6MCv1r7SzfpZ2qTfaohzGSMzgC9n4qtkNQFiqx4lFiiG10hDr7
+iM47/lulVyNjsI/3zkEVuXZ585HmWxygnu0RrNigvGcCJcBOPUFBD7bc43YXzmA
6rdl4BoFHiFAQ3/TjqVoS3GxE9Hueb4zBb/G1V5Uc7lrALogrAtWh3c9cGN2PAj3
AytczswUPG6EfGIvz0aV2O9Au7vpjzB2rVQOAG17BEv0SZQcA2ykUa9trFe9pOFf
L5TR0Cxmf2GyaecIDb/nibV0gdrEWpGcZ0PkdFCJh9P4vOoc4i/+jOyVxoAg2gDh
AJoTjpSLn9HySYzq9UqvCnDE6TJ0DRfVUP0IRsOG+YSGRbg/d46Co9wwf0dqEa5q
nNM7LTaG0o0h0fzT7j66HUVpzevypJDBH2ei4MZj+lENsrPwWu0+nyD8VdDajYYW
TXj7y6nrlI7yHzs2l/lfeB1CiRd4ONK2BVzV9JHVBnL82BawetAJCOpQN9T6S1JO
fZQ/7lByudsCvvlQ7Wx6py7+WwOvM6RcqS6QhVDIOYL7GL1g4YrkLnSt/Y+d23k5
GLhYM0EEQUYTS4aItGRUNHa7VthToSVcmY3105hM+CY16+SRG9VxIECSSaUrDbfb
Dr6xVD8PeHcNA+RyDzYDCarKJV/PZ8ugeOu5kvkbnOcPrcOStWAi8sY9Q95uO1A2
FlO1oyjCptFm9fOSnQ6hQPfVHHiH/MO507vmtRomXqN5sK2VcJjCMxthSkTnqBC2
tkolOY1cC3hXvqbZXfWyXfv2pkNDAQUso1+thKqH4HM5AEcUNl7eH1mhsXNC9DJD
cLDhTScq9bNHfvjmyvOlC6da3VpzU9sOlM5u9yf+h1pTfXoxy/BwR2UP8ifc4UOh
BSh6891uQbi5efVYN3t59s+Wdb0Ws7pUdtRTr/K7Bcviw7IDkQLWseTRX1ZRUUHf
rhu45uETSVEUyN90uBr0jRbiGlV3AQlIwFtXiiLTt3+HkFC9VnPpBfvL19Hbr+Ch
4n8ltVICrV8K1vChFmnlIt2Aj0028yD1GEKG+5SpxQ545WGN5L6JE+OMPA/Pa8V5
jjc78AQ73t3aVkrVSeHP/2Qw4NSg0yvBb4+Kp/L0Ulq+xqFUJuEa9ZKqMTSS+txJ
fS5ywMBkRMvnO+lqm91lll9Fx88g0bFYUAT01+cWo/pD4sJkSX/rZAfpIX6MOSCB
lyJPgtl80GAzUMVm7kzWCnbMs9o3V51AF/t2S2N2aTN3eZV/59l7ilvNLP/O2fbl
HYlFKhUd9N0xZajEdpEvIiqHQuMuRnJKwo97F3rKnTFPsOYQv5GuWql6KdvIscvF
WmY/m37tUgcV/aU4TknzBtkJ3g1F6lrD/Kzi15C8UJGdcYR6NIfphOjHiNogTQnO
6QrFcIcbFuxzmSvdDcM82RxS+4fexbce5yibv41UPgRtoNvbSW0XrHHnL/7kfnwn
hB0BO4Z6z0dkKUSQShv4OsQq01Dk2WX4xQdkRIPKVzL6MiZCrqX939OwnwhGystx
ZqInh9QYHT0bqEniY5NVGE1lYZL88Rr5Fpdq/LgRuqJ7vNOyR0rlTnVHLG4JlKAQ
yrrLI2nqFYpRw4E1JUjGQL8sFhcPkRHlt/Wgtia6cR0bx7egMn6hL7Lcux2aKeHx
UGMX9/hTCm2/GeJZMnrwESp4QmxtE16qoy3sJWi1e3lXQjJjatsNFJYfgZVQPxxa
wrOq1Ytm5GyHCmgcnutIiTiYeTRtndhtNdVsnI0GBqgi+JlwgvGg+bhh5vL9lFn0
H5/X4j6Qd5EUBqHy02gfbErRFoH/3A4OYKk76gOKKNPBntAEex+tRbPUwqplrMLQ
/fBoQnHGjcWLB6rs/N3/Dh2S+ZkR7gPnZ0uv0LL8Pe9X3SMkyzoHopeOccSAfOOi
YgxPCQFGWxHdNEhdI+DVZVmw6XtZEG2+OnIQlhtFNBanEjIrSFH7jvB/RvTEe+sQ
azwwZPvzJF/aqm1j/f0wQO0Go3xBDWHR5a6qtfp5ZGBeWe+MLiTzToSli7f4UbmX
8Q94ZARP9ONdqwId5orPxd9RuaRw+PeF8XnuppyslN8+A1diLgeE3EDJ4Bk10sWP
pNOw4csYLuJt3ik/9AJ6JY9QHT4Xxppaa3SFdVeAnY1+/g1bsPCTskRsyFKSSMZz
dlE1a/sFqvnfA3W/YIM3a5WHpW++4luneS75GDURTmLa3qKv8li8FRYHaV0dm14K
Yn9BVkbWbFVVOdGbBQqB1a7MvGTvFUniQanA8pkNfAT7LLSilhGkZobCdK3oc0p1
6ozSNWPFwdYACw+yAWTEUPWRGg50NH6NjHrRKflrCSB1Hb0tCIWrVmKf51tGjuHh
0/KvOOs63+XehkMCbeZ6+neBm/i8NBV66puqKcF+imFp4I8+pgoa2Pckw6YFE9w+
VwDo56pY01gUJv6mo0cz0pTH7fNn1OE1HH36loIkLZPCVvJfgfmNSNRroyJ+h+cG
jRjhxlaCDqMPjyWnwg4Sm0tL0izRRPtS7DIwTcCJX1ZRGAunoUwldAZXMoMOOHZV
7pfZEoP1oAiS7yTRSBNPIKk9F2ExyNrALbsx2MYKXz4cf257EUA3FUgtC/6Osn0R
vyEjkU9e0KQbf8+vLlqR2exrTOWS/OVtOkKmIpV2inXZRFGmRSXIzI91RGG9JVWW
yBVV93zfCxCkYUR5NH5cF1Hd3xA9E9zay7cxLEHHwhKhFMYktwSoOWsJDYRwxRJm
vB7XlSA9skQFHZEV8fwxl7lSpHsfWCFcoKkltqyJhl7PDVvrqHNEvQmmsTD042az
1gpGwY2jmVpoMR7u8NqZyt+iiN1bn4Gk/dgCgLBn01rXuzRCHBEqnt9yOmfVreBe
6sfqY1jOC5IzE2Jnt9jVCyX4lF6AgNiK64kOLuXEfVVAkGxc/GpOj34o9KmpC5AB
gtHaJ1JtZRFW4Jh6SzvsKd3+NTpwTXcM1eUPM6HHvbHsumeY4ok6e0w6KO3XqJmB
UqRWcz0/BGuh5v6+PTY37zn8NEcpEo1ZthqhwHc4nawsHEE1XI05r6ruJtBOqghY
ZkTxORY4tEkmp7Vvv2AFK+FosKz04K5seM/KQAh3c3514+wOhQvQ9W3vrnm1W0Qp
s2aIxDCCbVCnHu9KTcdWc+6+J4G8tF84mClKheliDGBpyJ8BPcZHpPLs8icXyj2K
nd8vA6C2frYGnCWXJpXONWIGOTqVzHcx6gDr/PJR6+zlEkFOgsnXDe4GcFyLnmm5
yDduAziBV6IsQb4vkmr7t/HFg1S3J08c3LMy35Lx9Ui2u9pcqxxg1UjNokymCdIK
KAp5DHFbAxLAo/sXirtbTvp/3VHH+P621fhSll8C94VPTnRZSgvlSO1GiZuNnc5s
JU1gITgGJZQhq3MCHlG6pwmfbMvk6KMaSH14hx4Lto/Weikd780zyyJte6rWTflc
Li853DP8b26bQ4rkJFSIRuAJADvXnAwYeaHKJT8g+bSqajqKPmhwpMXx71nkqtXx
J3rbHO3QxGBl7nJ6nWSNL7f5vqkAo8zjPr7csqfMxkuWvTYYQIV06hErwg7hLzM3
4fHgF5DXwb8+taI11ashGsaJ3cP4szoFoYbR0tg8tTGXUvxyNmAZK5EtOy1eL773
/yvLCEDB0cuivBF7o74+SCpu/rXmFuD5qcUNHKeU6RRUHLNBcwxvZiieWM63/A30
apnaXxE4piDBrtZk7JtpaNPYNzEOH1x2H0Fr/qHsFakU84Q3esZVd5hWsdSOVDNN
CHwE54gBqh6b4rQ6nqkQ+zgTdvJSXOt1PzQoBb8ZeXUdUSvQ5rugbs+eZd6KY9cK
ZY1VvZRtISUrW5VcL//qoO2l3ZURiO/pdSjyYg4dfsUGozW0tTvEOAm2ejK/RL01
XOgBuIh4tY6wkf+KlIRn8yEU1dDfBTJYYLD7zf6vMeW+Su9OhT2kHfMgJ5kG7gJT
Ma2pVv31EsU04h3f/12TsO6E8LAakIrwRWfq1f9Xs+KSvZOvB+6oMW+7OerQFtQa
SqUaj6jk9ujaDgqgxDG7Q72yR9JLJ3vA0lGtOUGSc0uLUWxfy3L+6FHDd8cytu3x
aAruFTP5ATPGzZopWc/+yK61zGeHMunv5t0LAIrGsO2qBNoXi7eFAmORgz0Lnh7X
edNcqWdgQwW7zjF626uqt7RQlAdWk+zOSX3fJ3u2wZj97NbAmr+ifdz7HNOOMElw
eEzW9M9FdZs3U/BdNNhKVrVWDi2qzjmYTnQjxG/sqzgL+qWsmIVN5HDsAJ3QnPdf
7BVwlmK3uwqk2rbX3nYSyCkqsq3e6w7NXPCMXdMh1GIZIJJU6nQgQr/YyDmQEeI1
GVd+FYMWqOSlqzBKlzpmNZXgzn2EpdSUFlDTfHVbaSJ57zpbcId3+uarQs1ngRn9
t1sGxKX5xyOqvzpgBlD5B3MCIZI5ISXIaZ3hraxeMkGMwnBu1/HVsK4cJZpaQ7bk
bjZyGyG4Qbxg3S0k5VxriOYgx6pBbLjbOGR8XpSd3pUswnbVDpDaYGqDkLedGsEL
uJfgbp7yPd7PS558B8kJKwMgIPVaTZEbRtqhDrGJBLzN8qf1aywf0Ly4HdRGPETj
zwjn5qv2xJ2HnkBrucTpUFNnFZDBsQlQ/7DSEw1+Oz61tb1jYMAlUnKzwSPoGMHq
xm1mbDKFD7NDsuSxrKhkow3l0djic9EYZyPMo7tS6b7u2VBwa/9Bvy1xKVmdNnKA
CIE4I81GiVAfb6q5FGPQXQr37FNdViHmx4nGeXVafdfwPOA7awJr5daJBHZCZ4Lg
1nYo7oABX5egcs1ijKOTTDUvXv/BY3ZgUHhsBR2D9hzbD4opizo48rIAQYvLM3R0
33G+4G3dX1aCD+eHSuzxnd+DBWaTZr2KGAH9SQ5Cfm3Q7FPLBl8XHu+6geSkODrB
iQB7R8pNOKpMdoDaP9s1dGyQhLeoSyGHTPCqdeF+E3rZtN9JxaV3PpotnSEYQ2P7
Mlqrci98F82H2Z5S5fncElz89FaX5BrAPD+qgO8PRWoK9KWM8eBezOG1RO83hfXV
TyzTqEN08XeKlESTcMvVfB3ArnBeVkPVvKJuBt/nBQpXZaNugLRm4DlKP1jJqnnF
IWLwjAOIo3KCRiLDXX+OqwZ7pd3U557bowsKIwWUiXSz/tC4qKrUZczY1JDkvIsu
NYBkvF6t1uCAPBJ9Bc0BnT8sh0pcvgC1vJv/+HjSvKp6X6lr/FrcD+iSjhs2KApA
lw+fU9dC8HI1nApZuKgh8AD4bbYVI4B8y7mHjs7ZtmySxiHAFkXiPVbHp8EYtSSF
hYZwR0EJ2nxIGSPFN1vQqUtSA0HhE4lfmpBRRIODvLI3krgnsFMUD41w2Z5vcia2
CXTiXVHtu657asmuzLj84Rvl/lUwh9LPSOxQrZKowFVk2Bne+u39TOLcPar/24dC
fUnu/j3+hnRfhZL/bghG+bhQrnfIQ8u5Mc0hmEbdM8SNxnQoB6zmO04WZjvFn4wp
QK1Qet9FaMw1ck2zZxLomBph/1LU7aVzBBhfso6FrufcbhAGDcA6OM2bhi7O02aC
9uH+t+TXi17Yrg6GLHT0FuFdcHUtaUn0m8Wr4mXFMfLiQpF7MR+mUmEc6zxbNbWV
bpX8p2rD4wGfaKnYIRuORidrEvu49omKoPhgybMn1yl0fIZORdWJ7k7fa9P/TYy9
Nu68r46mtynEKRRNHASrnXSeNGS9ex/5Bd9QgEuCg53PdKne5hoxxaDd38RUDLsY
sKrBYy1V6LQjow01giXiwP2LYk2m+yzKCC7yqeqz46rxgiVO6X7wYR+xqf2bI3zH
ODGqsf+siU2Evo5gJTBRlaOna3/G9kQ46AI2HBIS/8YUhx5ejGvhxAn63M5PhmV4
AZFM76Jxq++QAdEsAc6TYnjkP64j4EczTIeCYvvMo5OLA3wQ7+uluCsKqG6TAgqH
`protect END_PROTECTED
