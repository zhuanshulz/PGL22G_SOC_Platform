`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HA4f9fUhJ2LHM8e2srTU4x0RMnKfKcJYWo09OKAQa31sdCT0noPYBlu+QwVXh13r
kY54Q6ZwqbzyTGNiyqI9eR/cR8s6JZM4SFHzwQnxH99ZrUwVuqRuBVQdubDLFyXm
CejoJbyE3xG7nshzS2u6s3xaimORQTK8DZB6QpFHxb+boMMWNcUym6fKLmQXecW/
LFPGgRl26c/F8ta1yddk6J0dG+KvZbO3rjuQ1U1+70TDpBrf4K4zHCp7TdlQPgBt
NnmwODADTPGjaQJJJ2sG3yD8OUlesa+0WUH/F/N+2kmIFr0uzVszja5NyK0Dz4/B
pBEhlYOV1/gJfAOWt4iYBELzAqZOfXXFdtnx8zfUBE99JZC80VNcX0FKL+iOMv8T
57JEYpFp2s9OBD3AKp9dqFmXNq+Z3JxP5/GtoeWHKv03AB3gUrrCSwr5UZMyw8NJ
mjTd6BuKqneAONiDwM/FSR2Ex9NyQqRv7VsqBE+3undmusT1ORrUuKjjmkQEBcLx
4Nn+p/PfmizPeLc47lmkXcFaCNGkNbGZpAL6KMJpt2Gt+4Cn/V0IFyE6bZ7N5OXF
oecmvadAbYE0wt5ph2AFcMzncMInUdg+q5gnYdeAr1WG4FXp8GbwO21h0d9TfLJ4
+k5CCK5R/jqVP+5O0tXweycWF/w8QRwQezslvy7KwPd/9/oLvHWM0zU9xhumztMV
gNuLUZar4hftVGngagZl9qF/IUQfzt/22yh3iRBsqWgpzKy393AwX6xhid7Tufhm
lfnbq4fP9FgucQBJMwzw2JjZWkQ6/kiaRz2gBjwbIFiaJ6FICI4Su8XpMFwXs6OB
u/J1ihO+bqXnzrv+xw79dpjSaJrI/NjEGBKnZhzf8rGTJYPWBYsI4BPW0fAnDBe4
qAOPU15t1CQc1Hl/QU6EVFtnHtvvFfAfY6eQGsrqWQu4PTyif8xthGXa3taspGxu
+m2GyJA9OMEtiLZT7IiMKYkOy6KPSxYE8nX5k3I9G+Zvr7NsBQabU6B4/uDOCbtF
+GKijwln/yZFAV3ZicTTjqTvsFvQ06ajLARrfbLlTETrUHrczrZvbJY32j/s2LIG
Ftf/FRafQkDeZ0+Z/NQJlsAo8uhNgh9LgY8oFcYInta8WyCxJiho2tb/ssPbnY89
xwsJBDbiVch2oYDOi1qlu/NDqegNP0vmDLzyQA5H8q9SJCUcEvFzhPe8OUcUrnHz
TsSQi9Ix+Y86yzxnIlDHqAFQeeHjolieCtultkMqAWuPQRiJVcHJ/iOG/9EoGlXv
gGE7V6VDWqbg5gLTwq4u3GLGPEh+Nk+fGPrxN+OERTaBZK20hhr5Cc5Xpad/KY87
KrGyjVxQBUCmT5kG9y8Gpm2rDTmLXlmslnqnoSZv6dJR9KgS+JtOFvYk/zvDbhjU
YWuq5mt//aZh3KQJ7Lomg2BrjLeS6snPZ6TBxbVOLhunHMkSNZSmLWMxJlDsgqxH
oWWGWvgZyytUsUSvZmW0y45wwAFkfb3v/5x8ILdrYFNfTaMlzUEE3JbYDpyaKF75
kQotC07raBGgsAdSWWm2iuPeLbbVCz8ta1qNX+luZ6MLCzecBGev4CV1g8FO29f8
6IgqpknNSfW61g+mfuvzPReWIGZTZe9J4AVtv040LeK0abA01X4NDSncIYJ3AjRF
tDbTTiDrmsIoUBKg6eUKDjEKyzLeyM4LfkAu5rlVdNWtO/Qr10dUCapwTkmIvAWJ
JYpsTKYUEcj+jk80/KD2flAjoi6qLJ5cKz4k9agHAC6wCepZRPbUf1wRnke7v/Eo
twMcgo1bBFsIjEdCQ7lPMXiP/zY4VlGu6kBShal6zV9cW2jYkac8rkrDVh+9eD9u
irtRL3fVRv+DeTrLXcS76u1/RkJT5rbfW0GQpTpP3X8hd5KhQBwINtcWedzRMMIp
r3JsPgwH61dSBIYGGVXPxRNxH078LVpNfRaL9hZgbwolFIcAdx/Cu44sdw7lMCPu
ba/fjjfQlTk4Hjg2VaiTmM5ww/UkmdIMk7zwb9GySHfDCuebO5GUhnsIoRtbrb8X
mQRrCGzFALvjiT9AdbfRo/VEQDV64BlvgLFUOTOKBYcjujU7V6PXo2HtkGKW3j2m
vPezF3LhxG0qdDOebPnObRqIVNBnwWvzVGVM6lJwDKfs9wwHPESGK1JcnYNFja2P
rZc81+tUK7uwbrpE0urZ+vzhPLcv7FXrPlnCyVHASDfWXVoZVBTiTwsCeFrFJPHi
8wiaH6PyxBOEXYoRfQYWfCIF9HRq6QFCe/gUAog2DfOZSb4AUEkNIAgD8vA88lyO
fom9I050tYVoMYkPcl7JkY731jGkG4TZcGpIVVAnsWirOtVQNDRVSPUi4DTOqyp7
WC23EK02wK82d+Rl49ZGD15+B1wgFYm3Bje+tuA4hlLDc/4utkzv8iM5nEUDYJDm
Jo+2h/L1INHn5Vwtq1rXxhPY5i0tbw7lbO6NksSUAuzaiQbu1LTVAjD108l//7dX
uLOIi6bmdPR1EKPEWjUxLo96sLKd/TStu2ZJnnViC3KxZq9bE4at5xGItYi+zsEV
Hw8h7kaF+GugvdwrMmVEqoHB5m7GalcwKbO8tBREszqgy0aB6FJ7Dc/7RjIpTXZk
0nsbjLXFk+1tozwCRH6iWNErDV10ltyyD1s0tidGDDrPy6ba2y91tZ0uZF+gwDvB
S9CoNPkd3AdPXmwRbiCSfU4KfNMu+fdzjG98vet12sjwiWkGa+5Oa3MjLteHU5dz
aRbcSJnWA9C0EqA2bXWTHP6t3F/JRR7c6dAi6Tz8MVgR+V0agXehvYIreRkfVYtM
KxrunRrj8I6N3O92hz1aqHo9fkpvoUQZRBxuDQtfcGJnCRBeeyInvDcoi0bwE6Od
pyazDCvKdOE5odhwbuLg0SjAjXpZMFZqMgRbHoJfbi2nPLMou0TCR2OTLHTMyvH1
NKtR+ss4Tpm23FA02CmlYVkX5jJ28rSr+F2F2/sTJLICaBUj+C0aNpp30eg0/MqU
bU/EHxtRLZa1gsc7M5U1Ar4mH1SYYJtOJA5RFtWybQwErE3nhFpW0qMZ8O7c0ksJ
TeIAmSII+8uvZj6OzW6nVFaFX8ESWeWH64wgB9ON86xkMQeVTge+DzSvM00ujvCG
jpWMVfUX/s6Vvjx2a35ptc2AjMcfLlmfrk2nMYVYs0uwyDVB4g0KYzTnzHsxrj5D
u9bUugVT3CKutNu+6mpunucP8LfI919f2Z8vBmjy3osTyrNma/2qPevIzQS2YB6V
Ae7KLFdicgYKGZLjAYUBq/wAj1iUMhML6kl1NKS8YIwkT3ROUcQEgAeD16I1A9wZ
PH4plKaXEKVeFEO/o9cvMOlEUp1bAVqQRi15WQb9ixfdiN5cEK9Sb9bQZyratNJ7
KPQ9933jtdA3stvfXkn69g2PbTWb6vBblngphaY9aMOH4xzCShUBoUVhG8uL40a9
ja5efnAtZJeXoBGT5CqnAdBUhgj4Vqz9FvhbQXxmFSf77l5EAPYfdP06G8ZxQgAa
/GBA8TfAnK8rhoMNndQGn//xpkjaTlaAD16wyQ13ZmrBWFTjTDdhW4y+DueTsb9y
FTTQBfZfJ1xrLGxM2Hd20A+eDnPDEq9D7F93U7eUN3o/d1p94FOgBxZIK3PbUdBp
WCZGusYWT25tcKl5QniHDwqJz7obV9cadyuHSowB9kIWnyRoyyjn5q1QLQpNn8fX
cGq+yXyxx/f1RbGyfKd3K1ctljU94GpKVJiek+3ZZMXfWoxD+ny0RuYNXfFsBuob
jZR5+1aADmWjJEPQWNkyIrR7XrcvjJESs/OLIEnY8ol6B+IDJPFkKQDo/7VYUmRw
muEHg0z4IR81hTthPE0nlXpcfah3tlGhnciR8CQG1PgXgDCPQbrtMN3RgHzAo5c5
RombKIMu6bDxkoQYnkPG/Pnv4Z0ij6nTMAniKWgMdNLlt+fLRdHBLZ+bbuwbzmF9
OKKSVDCTBrRX0mzXhGvuzZZjOSe1RvuRgAl1RTFg7UxYqSh0sBr7af5v2IGwP7g4
z7/ik+rpIDB4WA2fDHrDXsHMXAXp3Xdnzl+52jPjFk833s3U1miqWMtl6mQ00j5W
UuAN3h4PbLI4U6So5E9BpfwGeMNouvKFUpwwmb1cNmhfEyfqL2Hnpyro7x4Ay6lY
9xUXUBN03voCmh7kJTRwKWKFP1NgOohYLz09LofcoGNKFopBOcHQccAyT4sF10AY
JORLPoQ2jUmt2ZsSvPzQnSB2dyUQPMy6MxVH+Ju/jc8bSUpzkd+PdWzXqnN41zIz
PLyD3dRbNGVzn/5kZRihlyji4vD9iUnunYCofZKWQb8W1ukdD1ksHHHfqp+lH8Q8
`protect END_PROTECTED
