`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8FQJfdscaYtBwKFz/FC8W7uVH7BCAxlycAz/3KMGmKhq6AEVfh/xsuWdcca0EdsV
WR+v9dXlFyjsreiXoIYW38qiiVrM4esHWCCv/jcGIfyhm0uGl2+09IZHYufkqZfd
x9ybPoJN5C+1j8SGVCrgBODUYAaDIJ799oAyFqC87ahbtQ3fMWi1rNgPX0cnDv4t
b2+lsWsGxr3RQGm84siVA0aFGsavF9UIEMkU1X8aseg84L3idAo99sGyXShJwMKP
nV+Y/jwSMYSQxAwkiVe4rLSQdrrAO+3LhEmzf05hF4MDopIWIe6fawviNBlpySrk
arPHcCrT7IdC5UmEJStBX687zacuFW0AIDVMwnN0kBodvU/YlK8JOAJw9hpzI9O9
PhiLsAGK/uw0LGtfqET//Ko6HN8daUMNN58UNAfkPmR44eYVvLDFsqmyY5cANAxE
RvghqpaoPmoQRZ8pET+lxfXqPWIMUUUD0HYz6KBYqWlVUWDmFkLaBoqjlHm0s3tf
sqTX6p/KyPbaFBWZjEQPb7SWjG+vFRAeZsvto1s26ypmJciIrgmAB0UVdsFhCGsn
ej248GQ/GHYDZJaFGsl3HHgT7AoADxKjVdliHRS+Ao3KGl4aJXuwoCKqvovuF5Lf
Ch5ziQR3fbBT2chf4b6aB3U97ucNjuFP+0THDQnyDai+SSQF2DqCl19sQelDImp1
+UXRaAJ9EidPwIIK1KL37yt9DcORLUCJd9glSNDHlCc8Z2wPY3lGSSvBahyg/vrr
g3To7/l2wnvdDIZcSWkWxfqkVrVskQv96OOiL4CGvMQOdLTfqsSKh8r8ZQUOCc6l
3r9gDqEfqzL51m8OArfLYW5cgqDFXgSLTR+tv/HalF9gRdOTjvv5w+Vlt2PD2LAj
E+oShrj1hMgR3MvfatEg/bpZhVN7WU/Je6cFoQK+rCo2hCUyeBJdpjOVdV+uHwf6
AHb9KPhHhjvSvtuOL5cnwbZJ/Ok5GxgCDd+yL4jHv/IPU/ExpZJMHMloDY0f+SkQ
g3bWY/QxJmi/KJTX6bS9VQhrJ2oeAfniszyZGOElFXk753WgxCIgeIaW6qD8pa7s
ZvoRaTHFYmHB+pCdQLhW8AZMKpNRuiQ/2+N0NP0zssCEe9vK25xPUE8YV/H3RKkg
+izV7lKZKnLsIwgg8maYsEaClDAevm4XdiCLzCUC+kpFVnFbCx8mP/fhFPiKVzN+
jbMoXCwWTY8SR7R+rmwlbk3mtmT41ivJWc4uPmdvhRbRext9X3ro1H04ttlqo00+
Uwxi4MhqNtpdHpPleGcVchleqUfbfL2U6pB0B8sRAwfpPiiF/BmOzHnUfKaQ/PE8
26KRyppaXxa3RiFxXKrl1kh6FhXw8QFeRgqPwv25NvHaNpZ8mv0Z2GfIs2Hhvs5V
IKvuvGkhqhPLeqK2GQ6gq37OISI6xstVpdtC2/I4/wtGXPsQEcaAOSjbaI09vmdq
RJjPewSByq4EffNabe5oBg3WkAv+4z2Ms7ASNsYnJq/NJr9lFyg1KilAkfCeiQgX
TAihOa336DTopp4w96KoiH+962WfrMrz7u2GwBCN12/1RUesx11TnD0elj4GiTdS
Ho3PMdIKx5fMe6fux2lI+O90NKTCLFob3AHMj4aG4p/5wpsKvXYrVAcq6YVaxyex
9k8Epe/wd/b6B1ChXYpzBvWl6OKtjzdHyiKEJyqNbJzHsgJvOtBm3DvbYhS7Zyll
95OCznMd3FhJ22tz+NnedOXXUVVGFh5AEtvFHNlh6VEwakXbrAhA+3/cV9LGz7B1
iRwfYyiW56qfuVwJ1abidJufk3evwoTkjyr5smiykRH/5SQH8jIXL0tUaVAqT8PI
8FQDm/9kiKD5A3WyJXvGoymQw71bnV3DR1sl2W9vZrMMEjfbcRcYpfkwCVljr4aK
IJUgzgIc7uSeBZcMH13W/oo7ZVQi+kSauFEjjDMhUfOZHfkCNK2/p6oojttd8Gxf
7ozQjVf4x8RZjRskk+VWFqD/uC6L4Bm/PifefdPnLsqwSeOF6OYJNEo2EOc/ZnJX
y4XwmVi18vt1iZErJCq5AArvEo+5TznAA6DDxFIuzX02GzZvhob+KlF1V6TqwA6f
W4YEQd4nn28xS6ON9tWhWr+iZ/0XkdfE5cF6oeDkynFscX34JTY+oHWpGkdjzL9M
85UUr0kIwhgO4K0BMS0qTrHP16rj51BeRXVSEDaVxkwxTm2fALHAx4ZJdEIXzi9J
K7FEdq8zbG7doHmQ9x1h76fPB0cGYpCTTbc+94CtSQxc1KxhkhnlsU98j35TpWXw
XIEilOiD1stY3cY2O9kZEwwYsMa44DAgzcK57HCxYys2750akuNivnUQnoc+uzSs
UbUUW2ZDNJQ4iJXoI3OwDTW74bKvt7JIMKdoeVyUkap5sEcqb19C1w7LokwpC6wr
/QVuse7ENryEYZKT7jvYpqF3hepIGZbpIC0kkS4jCOauUubwNWBnO+TiJ7OUKHq6
JBHTkgCu71+aZpQeKloapE9NFHYxeUnC2/7BxXGxFcdDZrO5rvFU2M/r+HRq/Y/T
cETP99agjiNVRrkJgMyKoNgqPKsozgiB7lhtYsMevYDoyhcV1fvC3YW7x71rI+4w
aKTxofIhNumiGx71JW/0xOcX0NuaOEpQGlemEwKy3PLYAyhYYyxBJVSx+TukkJrx
RknhXWO+HxOXGLmEluXIvad2rFGsVGCSnXMkCFg9FKlq/4Dgo3JX+UI/wOLHB4TC
HwofJB3MjfZzZx3L6QgwvFPB0y3zI/bWG2trNC4kTfIWlR4vi7oB92BX5a+nLQCa
bFPZHKEUKzvsNWUX/l2OWv5JwfqtmytIsVMfYm3mS1lZc8E7Jmo6WIuJHBBWrzkW
1C7C0d7oC2hQO9kzvzKwNTUD+9r0yEs1bxYtJQ0iKKgfJ+sIr05RGofiFVs9Z2R+
VpbVkUxODByooi5GH4Vk3ZoM5UlOz2lmNcic6ZwrwYUG9qfpDZWYFm7nnEPnp3D5
nkFVP5Q0GFMwBrNH6OesyW/SA4/OsevX15Miz1WTouwt4AJkMgrhGwzTk+cvJfba
4ZYfUX25FNvjpY/Q/q/M49jUxXShzO5LgpcBOTP573eKWiEIgHqnL+HRSK8ycQcm
JGBDVysbSYBoUIznn/QaJh4vbmyw5uoMHYShRY5zvTJ6RACRSDggIKUOLEuL+erO
E01UZEYx7h+mD6p+9NjcnuADRGRA4dkbg6bsyfRMeZyl3rikfa/dpr/dA/yTyFFH
OFDhh+BcWiIWXaoI7CBM2+yrZsMHqeCSEhe/Wfwr8UtRTXX+QJiMDYqYFT4peNJo
9pyfPDOb4LTTsIy5AP1HFA==
`protect END_PROTECTED
