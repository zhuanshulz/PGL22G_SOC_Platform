`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nBr087JIFm5HKSTBqM2oB4VGftk11owEISZR4/DaHz7XeBzNA90KFr9Dbnzf/awl
S3lvdDQcr3fusUhZ35Oi9Ew2nf4eETEPdhjjAa9JSQuf0uVFv5sGe59dKO74oxfq
mEiH8pcwpB0UYCGyZLMfof/qsVFTAtUs5ci6fzkU9MVxzTYKPziYXIUIZUEGcMut
zzkCdanGo4OvuHZ2kE4kqO4YutGcxBvaTg4p/iXRukO1Cm/ALR850GID5HkbAVYA
5C8VWhILRsf2CAmLtlHhZVzhVGLajR48AK9c8lIdXwKh5ZBomcassMWv4IQ7R8sf
YhO+Ua49S1j/VtGl/FkRLBPfjpcAWt1aYCwD3Heja3vuKRTCDcC/5p/rGd0mpwhc
xUqxVbU8SBhv3PnP72VrsEUlbrNeNN8MvGBrBEHKqz6WCu3d/qOX/PW5tDSAMBzG
AAQHfcsdj6D6P4cB4cbi/8Up7OFl+UZJ2qRsNlYcCxhIheer5aGmoZviJxvvrM/o
XX37pG7D26pAW7lTL0ZAEGB6s9GpqQVM4Ro+1s2GQqDpsyo7bnIKTpNoRAD01wP4
sbXFmJRjvlZ61ZfaY4COEsh6dzklTCS4ElLAZ6aHKO0ZOe7TMUrm7xomjerTRA9T
XGmnVZJJCTbRql4f+EZmqyswz/WI2sWIyoB5ZRHA1eyE5FWLkRvn0ITh/kmFXR7j
HDXUojbRpmGDZq0yrjEktN5DX/PhId708hsiCvBR4H7R0K9OG26dgXGWy3QL2I6r
FsSCn5mmQMmdIlsi4A/DiKpXpyCk8guNv+MINfl7dIg=
`protect END_PROTECTED
