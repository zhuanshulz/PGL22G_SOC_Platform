`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0rgKz4TOM9NfLBbLThqWx3BkCdiLiXDDL50GLBzqnGTXnmSKbFDSbNDsdFOew/mW
RJzIZGD4wb9+t6tOhXBWGiB1cGcmuelKPGMrses5mPD71y1HTpqngznbbdxKfaCD
6lLt7x9KHLp1s3qb0OJqmw636VFIE+kwvMHfZ4Y9pr8PQeXaltxIp4Etcf4yXlI8
4K/QxayAEiy/8unriQKLkv9P0fE2lOkfiKHxyJpa7YOUyCkRHjOkNMCGuVlaXVWp
gmd2Po3kDldOfT7A2EXYdWL4Mak2BDCayEFHVTT+BiE7NJEX1vnT4Oees4KaKV/6
beczURtqQR9gIzktlY/BXk66dyszEwdeiUrQ3Desih7J4CfwLpcjv952i+v1pJah
cjxr4iHHwAVmY+CU3aMd/DyQ/zSAQxh721MyK4OXuxvFw5gOvfslZ+WAHSsKyoBe
0fMrdt4Az5CDzIJZy3wo6DDY8X3GoEDXjbpDUDI89+NZH2XwHShFRn+xdNEVqcd8
GJtV4QlB0mi1Pa0jJvYOsIjREXRK34czN1O2g13eZiOLy5mSoltN/aX2sydn5iFz
ceO1dE6RzXAYfxdfGZxLsXzBxkJeoqboHdDLxi/NLE3yy6G/FjINNYfJllv78LMR
AsfyAZfN2lM/VQp1OnlyIULAlioeOwifylMBarWEd7DpVTJAv8kUIDWD0PeXL4cb
povpTlTpVumSKLK2Oug4CfigHTEsoJuhiRK+QU/G+2wplBNvDKIatWwGIIdGrr5V
rfhFaDtUcvN2xcTaHoLWdvWOgCKK4J/ezL6veikjN2Sg14O2CrgQfauJr5gtz7Vh
9FAsgNeuJpZdN+DTXU6PEc+KNZ27ql+X0TG12bLZVPqp5eEhCK24BMPa+x2rvQTC
28/rC8iwW9XGTM5LX9P72+vfhh6wH+1ytBeiZfwRnqIOPc4jnG+YjNsweXYeaCsd
cqucbjWjJuXZkhvhh8aWJKupyKusTgTk+S94XMgojMttUaZsWcyLJLNgC3zu9RZl
LztPMT6t9hIJqrItcNLKrjurc85Y+dwXEtkLe0knva5/OeS9rYTnHzkIN40ug7Ek
iPT+oT/gHNOHI65BE/eNkMabJtHJKR3BoX3lsFkBpix3DbiSUi931MtczRPJHIG5
8QTGPKM7Q9m0CmBaZACkkGLDJSbcmjFKzHzIKVNeOSmfE5nDQLiDXFsqkG7MoJ+F
0NkNKrQ1dLn3aA1aE3ZSV7cpgbhXg1GApzHR0fPlmTeJbndgOzC1ZrOSZr17T8Vm
PZQ6hvsyiQ8j/+fDMJsP7hitbuezkFhh7J6cOleutunYQxLjVrISkmjsbjSXr/qs
JC4lvzJePrQcGeZac12BsPPZsCCvzS8PabYxBqtcRrYiWgpFu1U7nejETJyyOj3P
zmVctHJ6RZ/z7m/KGQRYJ5G0TOV741zWC8BE+z4xPpMd40OHxJun6EPDYBI386s6
xTAdpeB1XIbhagx8R18e7rTtEk+mHfPyK20JxjfCekuhIKSWUNZrQpD/bIwLtSWy
ysfPtkDoVqW1YsuXHuBcRAYSdKG3gvf+CLPso0FmBQXfk1KretHF7kPEpSTq8tjy
vza2UbyC0DCPlrqV5BWNr6k498SALlzH1HJ5e2CpvoDMUqqi8KWnXS6hUW3LaNcr
Y3x7ZeQS/4OBS6IY8jdQCFs6JMN20dsViAEMnr8tUJMesD3/inhnTG59ey7FEaVU
XY5LLgu7nWBTXYSgrqn5D4upm9+nURt8hL/EFiEzIycB19o5dP2tYcrvgICpegYU
XGXFw8LemKqrd0fq1eBvBMTiiF+I+lsxAQLf6h9zZkE=
`protect END_PROTECTED
