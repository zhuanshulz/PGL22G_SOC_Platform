`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FaiEAbmKlwj4FgG9nhmIe5RclTz21rsdo4hlJMzZKhU5urA8F+jgHFEm9i0s5Dh1
XN1jzFAHzlDSEUoORaQkKhVoF6e7HYmVyz00buv6ZasE/qf9NRiJXjkZtyBwOKAI
habOQzqHa3eMZIPF+HKY285+yJAi1BcrHQhCmcGOLA4wFqH9vXIeU2HUGxfZWHVu
D7YgiH6Dw1KMOb3PFK3NHcMwmaqnTTax7F/eoEKrZBc3pUkvU0zmynd4J7MkFZmt
OLFKl4TEpRaRR8MLeqZJK5j755tvlUBn3zVo3kqhWqK7dO6OMnT9VFtKr9v9IHBh
+JEhDGm8CowLSO8OEN2rdgcKGjPUoQSQm2fcnaslUmY/QFDP23tnuc4r+QGHSvhO
lWWw59B+BuTdAg4t4/iKfkunHQb1K12hkBXc+tszBeh1Qg/pm0M/Za5Yreh0iazD
q65kzgN6VIjIpakBloEI+VQfJxGtL1qXQ3Z94NCO+JgOUO7Lqx7m8wi8nCCv/M/w
UNk5Zci0RpdjmaECMZmCoM5Ysyb5+drW+9Oq5mZtcFfEdn/0z3+aZNJrCrm2LMih
GJwzECDlUqcA1EzGSdVmVGgj8qUJC3k8tioPzhwWBc9Rl4AOvpEzX1PHvJjflHzA
ftMwWsNXQo+TjmA7ZX5NNA==
`protect END_PROTECTED
