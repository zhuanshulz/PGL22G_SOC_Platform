`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jSdwmPD25sepbvCRAIGQVyXV//Ye9OpTb8DmxoDgcwP1Y90/Hsz00nWbjmMwkJPZ
pkbGn53xaiIFYUZ2ssfqy2HD7zBxs/zJ56uW6jE2D+q4Jz70ydhpLkEshiBXCSWk
7khljb6AbJRz8gzkWcaghH88ub++Na62AzZbcAVg9xuvwbOtvzIMFm0QcQJSK8eH
ac0h0CHu0ZZikw1Js+aMvWgqz2BjdDLxZZblFrhBjWRs14vlNN6QLycJCMDq1x6Q
cU+tGnnZHr7DdAqMJJ1Xn7uIzYcmfihzjd+C18nPbRpDFDLVmUSlSs1bLiwrJjgs
uLxLmVJZZAP0MGe2PsZLF/0ZJQmBvCoQCB2bFo0BCDvmdd2kVroATXPtRuJygv0+
KD06J269qdyzclp6H45FBFUuyGXrvfm59vqN2YBckGuLJ2YrEmOCnGJ3IYlKNo44
N8MEo7NcNFACgg7ljeaw5r/n41Za/vrAcHNvHdJEwqSr+tBYiwMdiiEMnYF2Vjwn
73lZC+aWaiIcM3/b4aGB/vRXZXOYMiGE/5lc93nfoHM4ND6aDxu2Ph+q3bwskYWE
woUlJiovtngfQ1xHlJBlZJH87v+HEJ0YIdHVhqbxQrwn9tJt//i3hBORiNf8/a9D
9abVAbNyneSnHmHolFesIBlsWFmMxlhuiyVTG9MSogFgCiWtgdGRGBIjdiWhZqcm
CwMGL8yPHGUGVTahSTW2iNtPNOgQAbnSIP90Yh43wE+YWd3XGGoB4Z++LLaD9wq7
pGGmoWSlCNNxn39aUpSSbNKqtWJHYjWXTNOLbpKR1zprbUht+417Zs4mv7IitcWx
oX7ErAQ+to/q5FgVjmD3mrW2A6xwztCcAbL4H5OWWgmdn6hXpBu5SKS8U3t4nnBg
GvCPmTcwUnxs+h0/5HOEy3+ujOVrd8sSWYtFwFSleVpW3daNs4UWToQ2k6nQuhLu
FmyouktwhvkHm25Peiu36000CvhXGQRIv44Br7iuWdNeXgLRU70m1f0+wY9N+N1/
pL9lrsDmxheLLIpg/tdvLpIjWQ2r1KBYAoXy/rrOQYS/HLxhkH9Dn6LRxmki5Ofa
frtF1BFOCyuFhwz4sKW6DxtKVbLYlbBT5UIvVRhFomG4gl4ycKZtt7E2BZJ/NybH
Lu4r44UTpoM0Oaf5xipRcw==
`protect END_PROTECTED
