`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JuEIh7dLeLSwImxMb1dNWRLnHVe/Eike+IjsPdGCKw/gnf2KoLH1213SrM5dhu8l
8BXpz79wBgezjgx5EuF2/T6gws81r/h9ucdwTacKXfFxCA5ZUwlVFG/2v6m/LS/u
pwFc+zOnqZmitvkHOrPfGKXwkiKiL+wmgqdF0Zb5vdJvkXmVi/P5fclLRpHWjkB3
MCWifXGMqZbCCpviXBYxKyyOLFbepr1On4ITq0CwRXKAKeT+3S9ulkBhcME/mphS
OxkYfhRiPW9VXYJ2tMCNOh8YCXI2+ed+VVKho/W+2nmLgsJiRTVDhMThbWQ2zRQc
ObZfE4edcLw4R+I1t5Yznxl/nVuqiSoXpSnPnzkfPjsCnjdwkTGLW5P0DwWeNW8H
we0IbYkWozvi37lsBvJbMA==
`protect END_PROTECTED
