`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pf5ZHpTqwVAILUgb93bHssLWhb/IOxKMB0NkJogunGGhkQxldRhzrqim1PAT7y85
1LyutFzR6oQHTOfynl0CNIdiBIRhQzqbC0n5s4D+6sdCrqMzIaM7cn2CMdlYh4YK
TpPimQFUKYiUISiiYIIWFPrWrCzTmYEScsi30JfladLE8L/N53IOpeMvuq7FZpf1
Xnd29wG/Vao/4/7n0E97gG7ZLTGDQbjPShC/ceSOagd3pVChymarqwcmOE9pFHXs
zanZiXATvV5FUigBZmiCc0P596rEyR2oTfwKbQqZpQToQmlBlbk6cLFKOQesbk+B
rzT7d+vdny8JzA/Oqnmjd+j25yR5bTPJ/N60BeM4QWQXwZbPVTjU4X4DWO4nNgrz
6wd/9xi4TmenFN7UC/INQqjhzv2VD9Bp9lVoC3ihBupmJoQUKKwYwVOr/NMcE1qH
8mej48iI2nhQzPabqDcx1HN5uzL+oLy5McFfIPCAPay5R6nDfq42RJ8YvcKs9Tsx
hECRXSqWXtUYTbTXTOyT2IfDqAJq4xuD7BYTq+uZS+bY1d7DCrOqx63+FOH7v+3o
4Y9wps+LmLMi/W3ppaiakNVbCYq5E7RLPctkPmbmK+Uk9Cbx9UcgxxfvKaTlBPik
p6De/mBAgvsow95NxttclxZ0RjrEbofpPLzjDh/mZN3zw8gYN1LjfyrDpLPV/egV
/6YvkcopAbsZAwjPTAE8xQe5vsCMUCaLB7APZjxW6oMSMnQZd3AGAiNdoR6q2YFf
juFxWsRVyzdVes/B3K6q4OE2hAAIBXvkeB0yysmrwSYWvjcz/vyM1aREZ+h1fcUi
WrtxTYx+fxSnH73eLGQ9mKI59jzuibzPtQCWCaNU6NMkmTzPd86oSodiVaRI+9o2
cvwR8XHdC9vxFJMhNPAmGHuDuIPLb1qmIp4eZXmAR0zvx3889NoEFTRfywU7nmNw
JrkXWk1lcuhgQnTReDTX9R0mRnBXdcYqnwIxWkRKclatxLbYtR7CI3MMrZ4+m2tI
oeOkBi3BY0WQ/mSFGGDTo329/+WFU9cFTb+PRLrq1v19tX6L4Ajc+aJ5kr+qeH/z
WRFwpL9MZxBlPE40M5FTqjMe2+NC9dCUmzkeUl/ZKxlTCtT5gE8GMy+RzdP8RT81
lmVi849bKDHncf2xUdAjYIpbe5krUtLK5F/AnrLGblL1F4+hoCVriKUgY/cVt7OZ
1NtJMqY5zZwMgXXWn80tT0uvmXGJM6fpL3ZQpnJ/i2vYWPzOTC23QElmjZBekMAP
aZsXDovrd2c/M9e4qbquGxqhhXhqjWv9I69ankfX2Idk/TVyc35pFJsuBsoQ7NYP
KzBmouILOkbsH54abfgUv1F+lH8Yv1Lw4oKygJt2OnLEatBRY6uAl1n84noZXDsh
2EsafYSa0iv67eYGD798xxDYS3I1znsR8WGEWGqBt17uNGAp1HIiOmLzLI9v3I8x
JfjIVeXvoxz/DucuEivWoFNe3HEFL6s7WY3vtTlctxgc6OcvDGop9il/pIm6RLqZ
lr5ljtWCiz1CiCNewygy6EpUUZuPPK0mpjeP24UcoaYkWcAK33Uyg96PjPEDpSZs
oXFf4FMsK8GHTWA9n98egtztSTVCmVA/FDoqYMUE2GQcX5dJSy4YHfhs8D6HA/qK
n7LTZJ2OHydlDwG8YzPLKya/QA51YOgDOyLL4lYepO7IrZDeUq/ttKt2Q8qo3507
T2IOhdwvbDqzINKWF3WaM8s1tb7SSWI8tFyWMq3Rqi0dVS/yBm0WF5hXwxAx49gH
UyI+HWYkAwxrG8kGGBjIz8c6yW7UPzb2iA7+xyVA1P96rOFH5eVt+ZQ/e5yp5cKz
C9RAWBaNifhi+4eVw0oBfX+zzoAiQobhDgwcPMmAr9f0TxgAArZ7RV+RdFEtjn9G
2JigUUQNA4mdGV8m5ql5Kg2TsDer3c7uSchXrJmYpSEmOxAFl4sMmdSHECskjTD1
REfCQMemaHLrZxTEw/h36OfjdxqbYWhez0pyES0w4kYy9rENI7hVVPARCT83C5zR
Tsl2/9cACOmtWW7pKMadDedq/3FuL1H2uEDaQ6w/h8ADtz6ntZ7j4NOi8B6wNnYH
G47v4buBUETXdNaTVsp8/9nKl4iOJFun2iLpmEJ/55065Q4X80ClgK7BYADne/NS
b45HaWIfFupd6fXqzIZDpFtSsaoqDlfPzf8g942cRJ6VFSrCbiJvZDjpYiVUz8jU
dXEUBvoJDtL7JxFdR10zTfiec/l+swLWUbDNGLeuIB/eBMNWgJy3MCjCfCECRbqz
P6Emw3MDffDFLSuB/5SG5LokRbQ8VPBlK1BTgqISszd98j6RQOS5wL8wCWuJxY3j
XDs1BqYskxbfglhtyPdQP1+IIh432W6c4wLpSp8kbCogwlW5zkAp5pA9j06XkxCO
oCWtlapefTmVsGq+ye4rSQTXzZ4VjISRTwRz/3gQprhNX0Csak6H1KPCn3JlKGz/
Mbngn7TFCwO4zO9+LHTsMBORHbq8qjqpPD9mmlGNFXq+J3GvrTwlUb1PkS6cr9Et
OMDc976CSBo9YsbTFx9+gGvLwU4wF30PuTrw0F9rjQEdz7mzTPnU4Wpioa98HHH9
dIk/cLjonns7IEaC4OS4+BVsEc/2yigBY3wKhGa/yTuxu/f2+W819LBFoNDrNhIs
Pu0O7n0pQyrNhGCFz6lMwMjpd/oVtHVO3NJlYnSpyN5AVm1JofnxnFFe4nHnmYOm
rHtqbnKzXF9v+BjNePeE22cJmN4r9xFSISsE0V1Rd/zB4AkF/WLsvJoY3i+8Df8+
Sy0z971DsZl857XuMwK9p+9Gers4zRrt+oyzmmc3KNDH4dleYUJkwL0BYHvpTvPo
/DK25+unVSNb/LOduXNyX3UQajE8jJr24oBWULY7cJCOrbFVeUyT//E9x2MLzZyw
uNv6mxSBpGf7isPl0B2ENrZ8pxHQWhcS9COt/AFlLKkqaxQy1YGYQSwr8DZxFd3i
ovSv+oT+lPmfWwc6Uii9x5K+umv5O5q5fsmkf63e2R5OgoVT2llGa3a4JGIImOJ7
bCxfDjP4r8ShW1OGZK5n1nJ/BzFlUlWuyAN1GyHnkEpSTu416Xu1V2GupBrO2Gzg
AiZdwn6s0zCfk8EXPtdEb3Yrc42k/8c3tRIxh+N9jOF1D69BQhjckieQPa7m2Bd6
zyUiJrP2JQTYWxF2j05KRgCyx4YGfjxKmrnCWIz/8IcqU6hMStZkJ7XvjC5RJO0v
Tf6c/4wyLkJs9uVPrUkoMQnUEyMj6Jf48kdAlDEJf6C1YwtAsGbaCf2qzpUsktl9
VEJ3tsWrcwNGrwKbP+QQkWbD7YdABs62QKuF1TCKBIaiyl0t4TRwux8UipV0Z1Q2
Zjuis2a/34hJJcFn1o7hAc/eybadHXtixXg6bWMwffXZLijCGNwk3eX/XYeSnAc6
WXR2gDPNbxfTBoH3tjSJeaWaUd7pBPbPjPtztA9v2HydSTpQXPQTfXqGItKva4T4
ymdJvaznDooEK/BOPX52kEqnewSWQx7bpMwMcvoDD+xydkjf/1PsSuZmNhtA50IE
iT7zbizHPC2XmHOxp/WSbjXS8qSlS6/fuQ5/QV686rf3pDtsVPTAJtVhF5UOh82d
nnhYBU2XeDR70x/Siq2rnC7C6VyYpbLdqyWnzCQ/CHRWLA37siA1c8myocLhvFrq
YSMvDe7VYV4jkMU/Po/N02itrhk9NpV8AkYqSfm+TJpsNIpn2xwgpej9/7T4cAOB
E0hgFYNW85aDRemqYZk8hCI8eUFXZ5+tX14gJaHwpZ2meU9r3qFU1x2iY6WFIEZ2
xDI4wLfPKQ7LjRAKcc0O8uBxOBKS+tY3v+IDydA7ptIBKibaEJWikQN3TMg4gYxd
rRCE/1u0ut8x3f3SVFnPw8qR5YKp7tmIN40iB745yZvbR9Wv7LnHDuag5XxdkuhM
LOiF+O5bI9GAguPIBO+prTWPjMHnp8I2gxIFSzfAWl6HUurjzS4oWxmEQYcHd1Ws
ahNB0GKU/0oImeBDQSu6G4uhv/wZXwxqkq5jdAQmPoHdqp/yVNTQhr+ggkr0Ra0K
cH9i0fJRByce8rPoxScsblseQ5oyt/kGRN9rXHhygRIFdx8Ot11vQBUAtavGE6yd
YNhSv2adZVGiM+bUxCI6o+dxaJtK0gx6DZdQxsJBJz4MwyBtTNUGgpUBGT/r2Yx9
I9nqY49GfPBh4/2y4Jqnrjmw/pTl+AghfqPPwhpYDA8bOFg4cWas0xfcgiejQlgY
7mB9gLm7xauCIweFUtki4s4byct6bgIM7d9TTrb6zhWArR00oP1hWr0+B0m0tGpd
JzYYVMM5awi5EnmFMTuxEQmCaFpgF6O4Yn1R+Uy2BXxlqJ4UMCvUXR601cBJ1QbT
ngjCiSqFQznIaD82cqKSDEVSwMfqaTYpRcApe0E/zLs40crvEnFDnUv6ixJi1o7c
1t9ixkZN5cmnEfGtH3xeD394CoHCSmY/JbrprzMQwbQcyKW/gaetG7746H9UTUil
GHg1w8pEArVJlKHnBpKyQT6YAmTF3ES2z5smASlu6ztr5DFE0m5qHrBHv6M6AQP9
C4mhNZQHHR8aN5OjDhYfLHXywkwLyVgz1eUybHR1yiTjNLfGMx/VR9tiVH4wKweX
JE1Ze5xEc1QC4QrWBp+G+6lsoS6sMdHc/p+qdTIpjoGcTxNw1lf7TDTiEr+75m3e
A7i1lnXhJq3XW8DlYFVssaqPiSjvNplhnqgU0933LqsCVpVHWagYwAy3/oqAmJuS
Js00dsW6ldlKyVRK21triW21UyAgTl7eKG8q3bwUoYdv+QNQyY04RCepg+t6ZNLd
rGtluVPsfV6HrBRZ28I0HUJGrazydymLsbPFRek2So4Zu1pw2/BdLrWHuqkqwuh9
4/bhap8OrK+CEzLAgIp4GKWrNMg60JKzrNy26CkDDC+6yVRxz/JxbOrXe7fVOHPg
2SSvEHTyFelzikqcLSSoC1PkvOeTP4bwtgsaW/CCnzqyIacBwgyDRI1hehvqt31z
NptAcQrbKBHb/mdinHRLX8wVA6iwPJ2dDBk16vzdBiWlukR3S466SFoHHpiniG45
M77NO7oKzenHjtyrskGMiTT+ElpEuw8Ey5T2e1/aZLFUbr2ybQdXq++LYh2XhpIO
XGaATiEzwbvhsNseTxccBNpOrnl/2XgzlYbaeh+PsyZQRZw/77cGWXLkUsplvYdT
RFVhoDDfgJ5iCVvME3Uu045rBsBAT9Y5Fi2Pum7vJi18lMEJi7Ozafv2626hUv+s
v/Jz08qzkQocNEKwa8nh3nRrtMWX48RVBtjELf+xCgwAzM5L9Q8MdDKHoNnDashb
BJOC7cu84aBV/yGa3BlmNUp5cekypRUxAu7cGQ+XY0ilTNZdbU3eVgdqj0LOQ3AV
4utNiLuRYoVgq6exrIJkzVXhd6UmMbYGRo+zo8c6zftcVqXd/U5Qu3niE27Bj7Jt
Z4IptDsKHPVam5fuaaCCJT5r/izEYArfTa/evi5+cOOBTlsvIu2dGLMMUXRhpQ6f
i/ll6fkuUWDuBdfXiKsU4WZUObVU4FRFumtESSgHkWIrt3P5961gaFGUzY+P4u3R
pKjOX5zIEJdf5bqeH4G/AxXlu3oHB9wUa7TS2yF17MU17CNJui0AN6oBMnq0/2mm
5YMOzOpEnZNEEhseUvrkWxS3Na8RqC+Vdz0iiVh9DwHjH3kch9+i2wfVVbuNXN73
WrsfpA5RcoEzPE4vtOCX3Awf4GUAdGc1T8TtEv8nRzV7chNRqOBxvur1TOBvv5Pt
Q273ijevyLIpZ06ccdE78aKXJMjvPYEFd1Czy9Y8mtcDZStoP2RcreQGiUQ7zYr6
v494sHZ6sFrfFejGnDrXyYon2J51piVii1P50/BEquvhcdKjw+hVNhLVw12VzYu1
Q05VsXJ3lFd+bohnR2srJ0HKesYvxDRuJATjfkXVgpkNjLOpat9m/rBCA2I3jDmY
dAmwLSU9Ss2oJqMc6mczUOk0rYNmUMlQZObKIdZrTnJ1FeBju4WjIX2hzu96MXqX
anIFWAdxBV3OpQSleyZZjeqPylm3bToPviV8cyHY8q+qbvxo7zaDNpM4wWrMI6si
jHDZwRpRhuiUzCSz49kHU993JSLZUiwPTbfbSUINCYartgbh7GoEZdmVdMmvFUa/
NzfGZ+QZja/+LTy++eayCRjnb1gfR8UV+R0ow8/qkUmRzWfZbexE0stlGmvKeOyi
Gldvgz8Ioeb68yq6tjEKPSAT9z0unMlxplqpMdBQKjg0Bx/CtmDstcF40uOpMwrT
Xjlp4DwVk5sykAX6vVv2m287Ftc2/rrN/wyc7pFSbJH0fbh4/1ySfvcnWAuLrHfV
FiJgEsEAVv1/0GJyxhcz8shobSZx0t1450fQiPQ1OJFcic+IjLuR1CHfL+T1Pake
Iz0znD+Yri8hZAZhx4zdwGF22/JDsIboImR2X/kbWTp/0+tYnIHvu16wTeIRFNpf
platJc53pMZHyrMCbNOCDQToh7rPoerTE0mnAX3vcji/4Vopx5Ie1MlrMZjHCBLy
OaThPSgcBIRWPhJ7B8Z6zoHgbWE2pKS7loVLul7kU0gNiNGNvGffsXGWk9CjhJI6
0ZVZiZLrRiFnaCAIlBFSpefY18RIL8sXWLA9q5dJMyoGuq7EKvMWFCy1ENrcusod
vVSqFIUV01JCCtbgOqUjriexlbHuAcSlO5CBNV2APgn84jNbZBvIup0vZyhfHUKW
QqOtzQga5icPADRgYI0mxpCcNzpil4bLht87ulc3oIXPT1sJjJgdjwIUivchGR+t
C+C8IsfLhSdOAGSaASS1v5fB08sDAc6704EZwjeYxNhutJXHM5q4/7AyVz4ObiNz
27h0YAVc1OU/yeT2m8F2IBxziIkHRmyDNY4/UDq/P0Zntdak3dJDF/0g2BxIYYYs
CoMrkGMowQ2VKgPa98FLskmpkg4d1kq5bIje4L2s4u7xOCMezx8qMYYuaejPZa1H
aUPsdZ45Jf6j/0qNkRjBWQGiGcJJtvGenKYkpHQ+z/Sed3bSkPiXfeJ42tgAJOUS
QP50G5SkIfSHzh6B9kzHAjZERTW4tdl5s/+7dz3gwLb6Oa+ex9qqOqBRquCm0br3
wi/NsiR2XIqeqpdI4inqo9e2uXPmUlPh3uEkyrfQvXRZlbiYXmWRZkqPE1r0EFy8
B9OBryCDq4ZR5akulrYmN7XmREycjpK5B8+hc5I1PneNATk7HaCMeE5jhvU9OHUI
+10N7rsPsIy8n4R1wBQ4ww65y83QaX/WfrSScZRbs1JdMH3OMbU1Va9F6J+XAmkC
zkZffcJkPeZ887R/xYtqmPuQUt07VhCr8Qi5lEzwsDphwBtdML4075dZ1P8iS8DI
52/o7mHdW3TxpNrJOjAKoM5PaOkiDFU7z1YpLBVrK5Q53qgOwhFcTor6jtA3HuZp
8bbjXNVCzpZN9m64lUN3bWZo5NIgOMOlKLnEyl++cSxAFVg62lPteFMlbugjgyrb
kIxPM3ymchlFI8PQshbfr6nY7x2mKIp8/LLLNB9x4dcikRtTDzCJLAS+kwfnYQvS
V98VWif+6OPJN+Itw4X7fSTqXgPbjUmk6LIfra66HoD7Zl9ncUXqQXUfcix/yy67
NPYoX2KHu1Il9GGf+1ibOHYeRpBGwRfrIrc3g2Icmzyr0NsMjx9Ein6tbh7gzeEe
0iDxieKVhNoZBlN7Oz7xLHCZFkZcSj5ZrEQsZzIn+34mK5umxMSw0Kxgm/hFN1vh
/mRR5A3NvHPuDOq5OsIFFQYYJWfxgwXXbNNLi1zaGrYyWUwUXSTZioaYNG/9sT6I
yq62SMQmcGg+rrpQVgQPbDp+l7IeCyRMEwHmfQ2WFtW9PQW5Ri/9+pRqEaw3XTg8
sfDs1W8P9uHCCFCgd3uMRlq6boJfFhFLKd6l2IlgZQ9qEbrJUdr2hECfrVuc6slg
J1Ag/3NAJQZnI+n8jMEYabHP5Ab39TmBxEML5ETWpe3pm9p7RbIgKMtHi9IeG7ug
UqecUKnxq5j01nBd1pbm0V6qAbkF9pgWef5VFYKZQwl3xVULZtQGdl9CvjG1BJD0
7XyvBe+WtkoTKuUKzZBSqUtc5Hmzk4XeCQgUJnC28XvhHmdhS0cTkqWxjnC78h4Q
JdfcwlK0WL9lawf2UrB+xPpF+/0vNv9WWfu4F6i2DgY5U6mBl9skma1zydUnwWAD
Ej60GJaeersfia8i8a8Ecx5nSef1tJn3X4+8/h/oGXYSXdrsm+51g6Ix0WxWhhi5
o7V/6qTts7/kqukA965xgCrhTxrJm6UTI9DWlqDLgpihDCps7YhvYfOi0WjiIeB0
6cBeYNQgbZ8MED+Wmx9W9YQG2ZERmnJV5qrdHEKPFCozI8AovN+jLMrtAQ9KjJV9
sEPLdjqokde/Cy05URifks6CSUiGYYQCcaiOAomV7/mm6PKZ53seVtnLOUyBrh+W
q3J1XgUaBH55OqPUqrWiOdyPd8eAVEt6Ld9CCrZThuiftP84Iw4Vye4Hd6612nao
13plMZWDupmYnXsFWZh8dB7b+I7KFBMYGP9DEaslEH1GsgfnN4vVj6kS9B+wLKmK
ga09AxmJV4iaTn0wMFYQzbpKmqB9dEsc6Q2Unyfj0JM1ULBaPkBo3IncmmJxCnQw
6E8QkTbOEupTLHh7qzteoHqYGnlYww1Fgsqrv5ka1ALuYo5p3cc6rYV7iZImEdCs
1UrOXzNX2N2NQMytryXom0ZgsX7cR15c/k38DYkmSOOivT0DjXFNIPVwX4O209lR
E45Jb7Mn2Qyyq+qtiQjBk0nuB6YPmaVBMT8i7Tek6Mx4v48xcLgA5n8DJDuMPX/N
IXzM9fdi9G6h4ztAjbvXhMlODoxhgHHA+BVJJX6Hk39lWz1rbE8Phr1HFx3lnvGn
BwoJhrg7QhgFNnFRva5C05qywf8/HSOZT/EkVDavDEBq6VTKpo2wE+65G+5yNAu0
bKTKpLYcMVKUaPfqCTzyfx481wlnkD6OWsvxLPqzA3pRDpLOkJCbzVcII3fRj+LS
+0/XtWu8185X6pVob7VhC7f4PQ+fncfFd4rY/YLINSF6H1Qdt5DdVlhqtengbxNa
9QhHj4Rt6lO/pJgssFBNqXSuWgaeiscwizq2VZ8oWMOL3xo0sS6KiXet5H46luQa
YA94+dEPmvgBGznXcyKhE9vWCMtl5Nb3KX3hHJN7zkDiVwKsvk6KBRvOBnnROKcm
9K7X+vsXRKjCjw42uUI/Ka5sHh3ER+YLPE6dBN5UqHsvnX49x4QRA4jdmISHGnhw
SoZEEUD2HdAlbCjE10iMlH8Tj4CsguE2C25X07BP6vjF/qRALbUbOlZYr2v7m44j
2H0HjKbRvGhKxFYNPk/ad2TV6ton7TYX8YQCktHJMXukPBbUhjeRyG+35MygYG6Y
i9ExuqmNU+V8M2PCE8n2oDeHHdw+vgVGfduvMjk8paqvqmiyzHUeX7OGRlyOk83Y
atS4y6/JZ4lBin/OUKGJV2zr9455QtQZBDCc7LmX/vHqH26qwKItMqGvl5bSSSFr
kuolM3MVzAz8fdjqLqts2jf12YC16Ozl7kY6p+7g/MjpeKYboqQslaUnBmxtIfcM
p5pTtEOrFOnMYTBBZ9f7X5aBXs6MErS8aXbMneun1qEQ+IARnco/cFoFVAlP8tBU
6tSge1Nk0hTpgXUWrOkwLr9ekit9R+ERzuJBiSzy+vjufiMm/tSMOMItDgOYGCuI
1b9I8BKbup9xQ6acC1fSdRocvIyXb2AdJSfen/kviqkYeBINIIBWY3H0hqYcTJHk
UG5+K7bzImrRLnkc49T/Cr8Q4iMTTWNETqKNODm/tkNkAnV/Zms21no+dGvQF0XO
wSyqFmHlhwNdUj8XzcL9wsj0zvlzmBvGD8YAJUaKZi/WofwYANcQN3wij/mSyYSg
KCGZ8dvDQA3Md28WYqbB1Jkpj6czQSi4XadO9UapsH0wOeJ7VylYhnn0W9qxkiXI
eE4TbMScLTwt4KPqDK4wefTL6kRZfBlxQoSgOUp5pe6JuxMvBMjKlVVEK+jEHsLj
QX3VB6l7JCBO+bKacb5RFhWTBNsPDnH4iSg8+/l4kVMHR63XKph2+Tray5g+ySSm
x++ZDyjara4OfZIm5Gx7C09wl+4UXLMCJvSa+6HuaitLEF1r7gFt7WE1BDmaGPlT
SmY2SPlPYVeSHoMyb9y3JYZAP+Xn/okEJC45mDqGkydUoGodgRwWhhzudABnLTUO
hgqKo+ZWIPAtEsk2+LRTqGHPiyLHORfcbxpX901jdByAWwUSJl6tEKarDugHOS6/
Ii1kgfwZIxjG/4DK9DgfIgD1M8QKhw8eGU7NDIAfvwFcFaPWkTIMM+7YjXBsrkwa
sac3pF0a4UPDEYE4VdkyVwl3ZHNyNJTgP0gSbs7wZhhs1r3Or1M8gUuZc/tJbzxT
WVEZleaaAH3zwWgv/TdWb5aUCWM24ik572INRPYCv6mVKUuo67tvKL4IPvCPsqkQ
/PiyT/YelpOCU+D8lACSbLf6Nm3Qetqhgu7Rm/3/Ea4qoDtZszrxvXM0VGo9Osyg
Y+Vk4fvMGr9T2wk12Jhzd2PHBxjqL7SBAbUUUBY0a4sfbyZKVsu4K0LiXUN44ZCs
U4zynyB5Cfa1XZ9LJ9LuqUxBG/ppbjDp8oM6MgKsh7ubEEfS9dpuAOVCxWH2sAXC
YQqQH+SXazWerOtXwvd/XYzX1XCtVRWtrGMtLl5PgeoxTXw1SmwTO7KtMTF0pfa7
Pag5g90zjUYUll0gAcnunpAFY5S59h0GiM/LrwtXathBk5eWW6RDYW1krS/8nbuF
YBysWuLp/cut0VCU1UsLYNjoN7YR9clh8KxwCqLo42dub42SiiGVTB+QhaMxSiHV
`protect END_PROTECTED
