`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MdEAdAV3uutT944GSw2f+P2nSmxJ0d9A37AZZqJIkTyZ7htT1XX7A5p9wRJnwIvD
Vo0ydwsRqEFJj84O8GmKowwWMeTw99diicAERUSJZKMPYi7krXSA6tfOMzXFf6en
ehaxw93v/NGmB8CsErvHEtz9NJIUcw9BX/TKdJRxncORzG3u/ITwCfk8ezkv3BMQ
ZPCSmbT4E7H4K4bRNEt7TdXkmCdSnaPKOMfM/iodEREUuo3oVJFy70gmDROGokOD
IErt/+VxiVx+U6O8O2dqWhqxUQXepcxFSq2hiabP9KatNyH7Kx5jcjJspzPoOno5
2XQi5qP5hlK/uf4YNkm3Ub4WCSmvMrKnmFZUx1OjllhDZ57e+sOlwVMG0QIE8qma
84Aqhd4x/Y7jPbeo1CzTTGg2H+g4LdaTNW8vYYDI+b+ntLD2+5KulJfuJ3KBieM+
SbJeaUCAhA1CyKKWWtJZEK2LIFT9rmCyWv39dyh1ZhAd1yR1lc7XLiZ+st+4j5BR
Py3xAW5IPPIBSW6sZwAQQoPbN4eEAvuKDcLStq93YzWOgzNzyo0/RB0hRM3VKEAQ
/e9GdgiA972S43bCY4PpfzQuesYhJDYX6V3nfWaWWHEc7M56JOiykI4oe/hd80Bn
RzjhQUYXXXWzVb7m7XF0fxsCTEolG3QpbmQFsTRVuIEe+Cw0wnbiPZcDChCniK5V
v4BQNKtgasprzzhyD3Fxfg==
`protect END_PROTECTED
