`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PgAdxG2EmnzM4ULgt47x3nGNVMEK+CUIX/UU71hwDuDv+1BCHKVW4ZFsKD2195ID
gjQNYxcKttEyaI9m7DVLWLrKXZtgN4fmh7GrMlMOpWBk/nSMBh/UEplWqk1gl3xK
Fnbo5CimxV/NZhD3uudz+NNNuYl/HacPdeor203Vf1c5wSpuPnlA+ymjyI99NZaH
0fEL3TV4M4FAqDQMgfjFz0OjHuMpTQqxC0YAg5Pk+D70ACQH33Oo2W8L5zoWBZay
SnoT7Rn6jm0Af2oRmmA5eTfhw9KTMbK5XBtYJIMSE0M7g/jx/O7tXNjx8+psIZQu
BUGVnaIiE9BWhTq/Gh61PrKUM2Xqc1tcoXtcQXcXGqNMdC1nubhtTfiATU70JxGs
sGY54UzSoxh5JVRVZ16YVFZNfwAgWkDSQlw4lufJ7TiQpOKGXl5NgFy/da08J/kb
Pzo0n+UGYCbvXSqLT68aOuGjWxgO53pj24ANFUaR8QdmXQo+1FgaI0otJoHLHnJA
vdN9Ibc0XkWc67nIolU86temyOEAr+r35bRw6m7fLcjvPi8Hk2TpMDwHTeKbT9nv
GnCfIa1S7EZBlRRhCa/+/BufPigy6Sjv07YI8ZlRgfBv3hnykE6wDsotaq3dk6tv
eGba0K+7UFgtQjODDEyGuy7+b1FxIvIyWqfPI9fpKD1lMC0xHXavFFP3rmEpiHW9
RqA1Dbo9FTJPjb7sakU/cLe63clhPz2VWLKS0cNxtmw=
`protect END_PROTECTED
