`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nVdrSe3i8sP6gPZZUjjamGzFwn+AqrwUJ1pul95HE7MqVbNGnrGHO+nxmDGmAn/C
5MrdlLVYGdtIxtRsDYmRjitJXBtd6dMw/QsMu7ZE/Pt/nXtDUQFC3ze5egdwF3aC
YWqEaFEyMVYj2YevGzhJLhxxjr+GoCCe34wmOlmhkJIaBHMOmm/Q/yKp6tM1D7pY
4QkvEWijfCD9OIzhawS3G3TQ/k9od2AwMsApol+pmR5OZDUIkuSuISlkhUIKTw2F
/ux5dqO1++w+FI+XvmuO3luzauCNyO/Z7JzBhOtrExnjatNWvF6kAVNz3Z4L8ab1
H0J7EzZCg/1HjYFcLGTK3S6SnsxV/Urka4hw/Od+M4bDQG4rsvprsxT+mROwuINR
DfE9NsSPrzZS/1abGZ72iBwgSHmxaWk3NLcwJ8RztvtyadlNMAs+rr66V0FU+7Iq
/ZJ6CFiZR8gQSBZPa/2RKMGjR45LG4fNyQVGBeosYJhAVnp4gazq8irxf4wHBIaz
8hAQxpB3c/Wg4ayB7fiC8uIp2RtWCaN1fGLnz92WMcF2cuNY1B7FqPj2CLjpiT6c
KgGsmRkS3T8FdGjfF0+X8rhiBMezzmtRoTBpGPfja/yPWzwEtUUPA+UljSbBX5QO
tX9eJN0otxhYgQcQce+3achlJ9ex3gDyOEvSwvUOQudmOP7h+6GXPjyWPuECs3tF
E2U46YcPlQQ7Hm4kkepLkVdcBM05xwkSXFx9wba4iptCibq0iI5AwpRi/mggaLVV
+65K743rkC8bnBae8gETbZvgdsybychJijOw+DJ5sdzApsdG1yfGn9C3Yj5r07qQ
pIv5zCs+wSHYEVs9G7FWmSR2cvJJMw4nxk1h4dvDw4kk7oDxbqkUIv/X7G27LG38
Qq/mGHg3P6JjYNazqZrZ4DMHPN0ne0at1bqSayz1Rw9zAarTQF4ns2SfitQRSCet
gJEfXg2R4o2Ki2W+A63H/34mK+Edr8aorRueGtZn7KWQL3T3+MSbeIv3Ecn1CZIG
j8zl480x+GaYv2cuQKek+tPIxewJVzpcL1yOSQkrx1MWUba3C9c0pRq03sNZEox9
VFCy3cIVmFhL+C2VBlY76GnpRaidKwrwkhUi+RrVDUVv7BXzN3+L1P4X7/hpc2nV
tyTOpW4RUD+I27ZQ+no6dngdJNzxuABaAEhvAWxXh3gbbdMTQaCL7Lxefm5GRWk1
lT5E/lcY4QXAYKjO5Vz6DCbp12isGoIWTfzbwBvk0nRTKrVKJY0yGIZYLWB5+fJs
3tRh4AY9TGuRumnSmBaNS49Zlnxx6nwlN6V2A51M55JHcQn5Pf3S7fdQysgFqK8Q
Kq1aVgCa8ZadUB1XO2medpSUF/fheWgRV7OCERSLXQbv0GhlGJy04llQHGi4jn6F
d+0JpKijtnivRNTiaQ5bAjDSVWWLqahg5BzE4MCJyQfIuQWVzD2km7kmgK9yKwO4
CPKkz+YsOiZvQC+pqqK/EyHPgKKmT1BGnNWRj/rtmNJqztxGBX3N0du4w0YxWQti
8kzSG2S0H4wA8tpyccaAwQ90dUWii0UBSIbgBgS0bfEBUnH5nZ1Gk/I9dIFSBgJU
wnQtbi4SwnToLOjyjfQRzy7MfTwNz0X9C9goJ4ePfKWr+vcDH47sYR8uH21Cmg73
XfozC+8EuHYjSe9BOSvAoEq8nwlKKuPAZjkoiobf4hx/mpYBOsz9bT0FI90deVR7
bqYKAlhNxGAKSO5btUSWuB1JrfF2TToDbzyv3U3J3TdHC1FXMCjuGOgFZ8vTcL5R
33TCQ/6ypmspMK1rsh6dg8hxMY20R+210fWz1MPUj5KCMjlzRP2bjkB9sGH61AHb
dy6cRdUEBZdTsK0SAlKkxhY/OuYrTEY2ID0MebaGye9H+bQmqGSwHszUx4MyIkea
h2G/bxWYZSipiFmSNKIZSGj7XpA8GHfTXAiRHAucelNYeTbQYY3Hp0a2h/S1d509
ws190YRRJ379dO06n8/ozLFe8ad3c+K5lbMbX1h1EI4/5eQzqVcOKY4RF1VYesYd
AF3utU4QdHUHuNmNVRDQW1FHym5ySrFZswqfMNvB5EE/POCpB+Mm3HKCcuuAUwG4
XI47tsDqXWxDiSRRhM5pNbEv+X7CSbXMkyS2qBmhfD4XqBdY9QI3+wGaENDhQ7TQ
rUSseKwYLqcdW+jp9516RCeDWWRrOxsPZ0AQwxwNvtdbIOwTk5idDPw4X0Xm3RE/
eLQOymmqOgTEVKZdtvgHdSb8DCdmWaV/lzhijz9CXzMnnUvaRZiuOAc13CMdnGlS
pBz707SR2wgkjuIRfeBssnqaz0Nk7R4+GTsvVEb/qkcsPuykLe/2kcKf+boFgnyb
2Gjy0fRQlEy/WBIesYmxlKh/htvwF2YlZ6eCzTVhZjzM8LSOR9X0XocXxhMO15I7
w4o+C9SFokD5H58MY7U9ksao8PiD+c6M+tDp2PI4dUqfdf6r76aQfO/wLULcHtus
bSEvQmATGqflJGKvvwznrhnrzKx6ZTYf55xU0q91g59clgLwHESJPb8gkElZdN5J
o2Zu+UobPMdN3RGkgBCra2yYBz9zZBIj1LPNOQ9eJSw34JRfzHiWowg6eWkxEb9O
C7y2d2pcoWVFQOwIOT+ZRWksRvVcQ1eMzBRwb8bFu4oYQpx3kOVEeNmAKmVu+6HH
ahhEragTnVipmDZpnYUDO/k1dn0E1UXrk6YZm3xTg2Ev76glaO6An+U5bOjoE59X
h32mruG8dSquG3Y8Tlr1r39dYjDzqRKPTgztCb7lVynz4bCpEvSuGTM87BUXqq4L
f4zUUkU5/nlZio9SfP5Jd9FSbTz71+ChIjSNqf7MXpJcTlI2GJetYkW71ipL17Dg
nb9cutH4PlQQPbrrz48JED/rg84e/8iRyYT0rDOkT7RbkvIw+4mq45r81vXxiu9Z
dgV6dTkwTGIbyJUVt2MtgB4ooKUau3WY74XNaFzZ1im3v5DxafVszuEwuhTd67SB
WnBXMzZUD1rNjGcCK+7hilniHdx4gcJo3O6XQjm7gFYfPbwG92RsvnOQKk5pPeX0
us0CBmXTFxDkiTn2hDrnSm/I/YwtzDhLm2+8Wcc29v9ZIvWdx5UyzuPyLatYgEWz
ac5J79rlFkxR/BwAlwekt9yGHJI0emsxZh//DdV76xGUuMiEhseQoRMx5EmTk7RK
ZxqdSjYIK0GycpXrpF5VjDxBJUiWSAUwOkhz3gcFBA9JKd9hQD24jtXAiIMEygQz
ZliSz0yCFSESKOC+8Xtpovs/8rOc5ZU1ctbqdsIQzQEuqqPbnfaB78PAaV0XSWYp
AcK65/PfvD8tKuSnbv+LBbIOX37sDA9HmbmTxo11IF830G8oCXsLMDWqy8oVgCJE
lSypNyZT7SBuCy3Rs8iO+l7Nd+pzcaSMn/ZDmF+YjLUQTt99GWJigssE+Ntg4MJb
B/ljkiO8SAHsTDUkHtpGnLHkxMDfx6O/09Trc30X1GAVDn84UsRCKhqpbnIhvMG0
OIaAWrybqQA7BFw2Zuk0QFQ0rLDDCr/AehSA2AVOKzFKLG3hz2zOKxBQmp/rfsdu
FJl2aszF+O47QDm2Ps/e0mmBNT0YH2yBaq+Y0eKWAzCNBATHBMnpqABOhLDfmUVX
nJqZH0Z9vBbSBjVBT3bGWyOmGGvoqOtzSeZGE1lN2CPST+hrVhKvvs0raOfhy0/7
fKhBHwtzjJjzNsmgZtLJuReeZpfosEllZI5AqPRHYvbQVcfhhTJvNJwGvpwIo7EW
dLDJ+YQVGK1DN/QNuo2e3CEYAPHSVDocDC1WtZO4B5jkz+ui5O7iyn8Owmr4+RLx
edtEduoBxXU/829uDn+G07qfgy9r67Gl3d4lsqPL6kcvM2Xf88EmytYKZOY6q0dJ
2YXIwuClBdEZdGjYT40b3yFoAmaKw8etrh/Il3fR4+2nb/bnCZ9SlwGI0sLnN91C
vY84JR0hJarSoHp89gVMcBE6mnIKGL09nzNJybWxXdeDigXwnW+UFKHSTM6Dopw/
YdhST61/sn2+iWmfh/k5/LYerRP6tkhrfheTpLl28KKX/h9ruioy1bEEogvlMSnT
H7WuNur0C3V0AMpP30UHjxSYstGLZVAkd7Wp2JLmefL5JN/CW8DZwlSCr6hLaSDX
g3GUBVtbLXOpbL5Fr2ECSK9ZyxYlYwkZdb8dYpKL2+cP63MTLNU57orcjMXBgUif
ezg+9TK0iVCRBhl6MGQrzn2kzda21lxBu50i4VEC65h03ZDyd2LLq7IU+7teNG0I
5Vc/kZD9rTlFcVp0mKVimB/ehneh+vvFUeMQJft30WDFBb/r8qjgBCv2toEpiaFf
8QprUVgG2H5Fm3D/ZpXNvU3H1GX0E957AN0E/XktQF//z3yAaOMK4P+VZCnjwb8M
p1TuYUfavL88qVkpxZRrN9cEq4v2L9RO4G9n3fdUBOxC9nm/rckZ9jXuooHyk/ki
ghM8mDrfTDrPges8WqDjuPeJgWXewadT56e2ZSoSecaLk0Rb/9SVzcPcUCkPFAFx
xa/Yxxsx2gvWvs0ueLDbuxNtoVsehkpTa9n5CeLvK/rfLI2LFcvqYONe4wUC8Ezf
9dNOl6kg8qvjFimvjW+d5ml+UdYmxGbQnU2l3tAms/11naHSlPOQ5W/PLG1+N/ew
+eB7IzwXGWdNOF4ogEdQp/ZrwC1Bixe9+w/ooNDT7ib4bFL1FlgvcCRVK2lnmuoN
LTQYRoeNJG8cK2Rv5Voqwg7ku/EsDfMHbud1V6Bie9h5jnRs2S8/GTK2MP10M4xF
4zzXYDjHOwOK18va055jii+4H/KerebC8EQa/rGfdOseipbWyXemqgEtR23jTdAr
CmUIDlqLBWpqALF4J7D4ZlAp+lPGU1sGOA1HaBIvx+DvywE3hyNSYdbnXTI2lYdp
4JvBD4rNwHeQ/JqQ6V5h6ikK2cv15NFIfehED7I0m8KLxWWlbMZnH32wUwQKsyfa
WFK+OkKHL6M2MtOudsS0qIl1JP8e/YJwej38no5P6lsulcO0MGMXuumuASAxE0sH
LuV0PcF2Y+uaZhEwNSK2IzpHMM/rq+b1w4zm0WWaPh51Txhd2ha7DS9SA9tZbQt5
FPNmTAd/vL3KgZSMjk3fZdh69/3ul65DbA4PVf/fxnTZmkQE/y7dUgTHf2JG9TdO
XoPXVszdP7/WNIUrP6JfJBtvq3VVpFUwQicxdoe+sIza+iVlnobzDvCa9Ezn4pCU
U9207rcW6x5T2i4zI4B2ibx1SPW4eeVN4PSFq583r+ASp8KW6ZBUGns8+7F49G8y
6NvwkNyeiDlqky1AtMFPZdOOKKFpXG2QOwgWS6T5+Sec0Mayb7r+CxRddxabtldB
07tuWPfiwbMydxuxBGEcifhHao6dSCFaAkiQmXUGk1oVUxsIO4L9Gofl/RV4bcRL
CmedGhNUU2tJDxFB08Wr/XQccMfTjJHjZ1M5Qg12w19XlRnZ0WgZPckh9NFBO0A+
LUHpIgUbjLgsFyz0pOigNObf5D2FVzWXcdck0+/vp8StQg6R6tJM8nM7T33PzVUa
FhCNAZ0+xq1AaTUKiMiARGHOm964WpUr4qhgI3BW9ZWA2Y7LFHGg2XKhzkY8ePns
J0lsFh6zkb7aKZ9ymIteLc+KtNCRPmm7dj2GDfiSN6yTSyA1LH6S5QCyA/Ub6WxS
fBQnkf6zhmY5vzIPckpNrEjh2LP4GdC4KuldTjtQgEHyJnGzIkhLZRBqDR7qKPA2
nq+ohlfnTHGiJg6OZx51c2GQ4mOGctUdxD5PS9FtgSOyUyFZBRl+onpTj3rxx/5y
PH2BYaDvQAh/EWo0oJ2M8l915b7ZRriPrVKXq4jMp0NL87AqOzOXzORbi8Pl2AVl
KwaaUVl23hv6BVxfIzLVVLVe6oJPxuz8ZOtu5LVK3cYQnBQjiZwufa7FClwDBdfD
7WnotlHJKZGzYcp9Athd5qYnoAG6SDcR4YekEdaHP1r6il5nKNIsQTOJNIAaviTE
8yzyYZy8SlLnsnuw9jBeRbPLe20LtG2oNQtGvPofFTYuyjF9eAzLV2AMBuAC0kfe
JFrPiEOIx9kU+iWTTGfdEDGCsiCEEVDNBc69A4sj2vE1JEI2AQcEsCHyE7hHS8VU
YSrxNjHBVLUwW7Jkkjss2RIigoXA+joxrzXSbqiZZ4xu26oN0t1v25KogPALRQeH
dceC8TEvHHdW66AM2zilRymW9OU3XzuwqvKGZpkLOn4m9QWdrPrYigcAJ0/mXNvM
c+ryRSm5KvV0OAWIZEExspuk0whIshKQhOAWL5Q3cMYctKqjIHAX2dsoPUWJC7f9
jPI89id3RB0CSZCXharbC0lZEPuB8E3XkFZk4u9YDF5rjqr9jUdzeO2UD0YnOsv3
/1R6PPOFtbN3fDggfWQ8JXgISl6TQNomOqOXhJQZgajJGlTQ9980dDKSM6zJ/WV9
bExvC3i338CfeSxnL0NtSd2HmFW2ecLK/bkV4EYTDeVijb9h5IR6D3duA9D+JmN/
/caOsZveVsSgDf8FPK9IjGvqlSzXt534BXvZnwVUXnIa3vK4R7mlUoKDaGqYAukO
V0+ofALn3NFXzEppmX68dzLtxGcggvVRwL+SZ6EOuImgL/qqQM75TqHtYoGpoMh8
LKqbEJFRwVPMA7L6eQHqgRuE+gYOLBTKxGVS8DKvxLMCNdKKYVNfwiB/2hm7CHdO
4UT1yerxFXgrNAPZpzgJAWnjM28cpSyACk+RtRs3+3RaVXY+2FAwFIRPxEwI0mc6
uiyBIcI9yez885NLTiB9OU5ONUTmz8UWzUCpkJkUZDCyIaffN79epz8IJ0yqHqc8
oZjc9qyUjg+OJ3SQlwy0CVzv7bH9HkhlQbTIg1Dd2u2EILqSo9O2ibUL0mV+AtTi
fA332/6lreWOiS58HZuIpd2loFObnsvPM1bJ5KVWJmZrtIOlvvlVWCverTw7U4ZD
ktCUPzggZdtT4kuAEVnmfAv2DbR69Uc+1UdqakMPIxOcGGpa0f4wfh0Ah0hmUTWx
I+ijcuOqoGPcaSSJ9rS7/HCsaH/il3MPpNU5Wt7H7tPnlsNEqGUAwiXcsZJ2R8tp
r0AFuxFN0nlgTjlK7OS4T9UOMS6mAQ8gEea0Kp9S6//L3n18eMkQrj1/OIASLweX
FjPz+dlkup8nS7zTgG9glRoHvi7AGzOp5wUgfqu7vi0Gvghi0TfJzajsdP/nHjYh
t76f94beXVfMMFSOARBvUqyqSo4oe1iWYx01oPETVFQChq+sc3Q8SHi3s+/27GAB
khui8fk8cWw3fn4DRN3VTHYcViRXdy2hCKkmjlEoxcP8JBGVLukYcvgdndn9DpbA
niniCnhc5rMH2p0YyoSH9+K/llgYC9OKE7x39HvqBHaXtOsd32KsQtrtUD/HeCEx
lD5LUV8NiGsbuONbJSVavlyXxB54Ovf2ZdzqcvYnwQvU0o+sL+0UDPrIbV8SBDfh
EGaV3PPKnEvYrrE2sDfcv4wv7nszBHkUpMkacsgzwuGt+owGSVJB9DE/PVmj0yHT
AYv3qWYrbsAQ1SoFcxIIWxc5cdGBPVjt6H6BQZePq9UCOdf87Pyy4lf5Ef8x+Pmh
GgJqp56fgyWx9aL3em2XonohV9J4Ird/A7YApbCYWqK5exdbLZ42H2Tgd1vdqBqi
+dcZOAAU6qW2HdNYCMGjDhKFPjA1s9oDHP/5sodoTd/roF6yeWRyu7dFyklBp5IX
YLyPGg7SDpzi/YFU8/tdw0anQ3hJGNKiKYp1lBFrZNvnNyyTbEvcFF4SpBNoDvE1
3S6VurGRDJNopG+SwLn5HnnoVCaHkDSeI0ZFPpW4I8XsyzEQNhqt9rn6CkMpojGB
76D6Z55zn+CnBTIwlDync7VsVeIjDRahEjdCBRQr6TooATC7LGHqrd4mT2Yjfm0u
ywldmFubTMrNKi0/hSJm153w4mGo8SPwOc2TVTgd5u9iGpK+3WPcfGO+WUcs4NLi
5ih6HjvFmoPztWxKptEwo8Te7cj4zTAG/HyhiNmaJ+Oq950ZkkTpRpfKr34d75Nv
VPl+ThYTTjk5aYl9b13/4L0kj/HX6XB//Lft3Q9ApAUwyjSaWWxNFlWH3yRkZqZG
K7Aph/NItOwK2SUemcdR39+Z1f2cgq/Txq4/12FnuplBuEEdbhh0s3ag4zlR1X4a
juqjwzTdYJb+keAZHuOUbbHKOiCTtWC6UA2bcqbGI/5m7XaJWwEGZ4q56MPu77v3
bg/RZAGFvafWest57VYJrsTDpy8IFVLJvye/ZY1N6xHsf5kmEwilzlTJAV0/EEvY
/qpF1JrpU5+J+YekEgoJzsJRtDlGtZWTqqqijSgHHN5xcxzARXnvrRghGwrq1BgD
clGEL46KE4e8V63SVSb0xjleepc6QvdhiBF5Vxw6XBfnwF2gz5vsNOVZfHHdMVad
GAy/ntF7eD+nPjvh7rRXGICagXpXMy9El+6lSjVhS6HhxoTsqf8vK6ztSx7TzHyp
cJwFAj0u/3x5zNgfIJg+yrtCv4IRQfRLMjRHH9vfUpknXXitmIcElr+/6P7UlyW2
ez4TMqF6q/5yhTfojkw0tglJKfDmPDtG1VafnXcAtqGPRrKnvPsLpVFfm/S1sFEe
P+ELEEdpDSmFraDBNVynopnwESVpjNjPeiW0sIAyaGNIVvyCYKUQdnqz2lAUBQbY
7KxnKG8xSMCAlUdBsMVTRnwoSgx7xV+P7bUx1HhOESQNl61k5u+MPdbFqY2mwflq
r9Cn5MPwajko1nhYPnTkyexPbwbfmLofgm6OA8WuQccRDr61/zfX//7Mpm6gAVxM
2w0fApF60Df1iojW3ocy5xQ8QuNVuQEvXwCmI56KJ9jgxQ05p07iysJuaDLWTipq
QviqZ1Ggwt21JP1XEnTO8DsW+PcrCYOOrZuGJ2dUq9GYBWXMHIs2yScKarG8FCOM
7BRfU0+iham4UfUPMVtfYZ8nrwuHs0RD9pUHio1cG3IVBwrtie/KTC6evyCQzXmn
wg2NEBnoU+lujYZLVILsB7SGGthxbjUHxaz072rZ2nE9OBSWeqGpU+vO3E5/tNNJ
Dqd3UclRzG/fnouC2lMphIuGw+YHTCk+sGPJANNVpLuEX1QKzkLreI1HAKpeZpX6
1fNeAxwLz16733fR1TlpN87DnPc/iy55IA66Zpg8/RvV22KUXkifAwja8Yu6f1ns
4/Sl8EHHiVEO1Stqb5x//fLAJkjG5NdcE40SUv8dG2mWW1mJjEDuaknXclAWqA/F
hP/D2RMjrPfMRzm1+2jbE4fEqjcZp6FWyYjaAvOtQbmlK0re9C1szVELySEr4OAg
MCXFWhzoAZZF+AjVXUxnQ++LqFnwgA++5FCaiiF8qNMMWLYOgZOpOyrRlvV6pOQB
ClOztAhc1ld8GeZd7xTACQe+ZUclgUPp5qx9AEvRcowhod0jSY8a/vzYHDf5pJ+a
cXpWevgLDbhOtYW6Jqz38RuuOj8nZacUpNB2m2b+Ck6a5/RzQuSyKXjRNQSO61+v
h9HtosAwe+AbmT/EDUgQgULiJHDyKkZO89G2OVsVJclTZoJyJeo79nYJNCkAibXY
n7pDV7ycRbL9OC1qBckrRATgH9CGuVcVCn2nexeVR669NT1zQsy3blM6Gd+j7OyT
JOgJdFuLf+dUvsf99jELhi8LJUFMFz3X1vIjemg4ZauvfJZlLBmVpodOd4wG7y1Y
6d//XvhwEgH69Eb7ShQYGj1cHj/cOLTG6ZBUJZRg6vOkXCWnV1ySPc8LZafqQigc
dLLtoJNBjQ5qztsh+JNBsYdAT7YilPaN4J8C6qfoigsj71pQTWjsNGJ01QJbVbAj
x6kHN37w1R19n5LRpA9cHyWLR1HsRr+dVKjne4fUrjLLUbXsNnXgsVIS/TSvJoRv
REGuLJImKxfRA6DgONpGGUM5kWe0aUfbspFu2Vtcf69xPkpsFZaufYHpKNfLRMQ7
eHbYQv8xgfHSpM1CCfA7eUzegukOs9inbQPW5f/QGKLMurUAqQUa+8Rl1mGuqwNv
S6EbFj+m8+oqQlwB7HWdMnkOTFTczbp8dbIWmXseUuW/+PiESb/Z/aDkK8Sy0J8X
AcoYwsybBCTBQWu/bBcj5B6c3EQN45LPyw/suWcMOpqSlcFP6qHIFRChWoxkaG77
0Qh+ch6/kLzgjFC/nmYP4xUlcTvLlfvjaT8VQlzOq3rUDacVm7AGdRInKJFaofTx
rt/WOZTSxyAeUt7kSpSE9dLU5ezjSKzlpx6bzXahxIH1TU2HWWv5iDGhEruazGM9
EqrdTr4M4dS4/qMOxY0xURHUu29vuV1NMidRTSUmaTYk2pxH/dtiTewji/yZmybO
DPv0Unz73JK5f0rLo7W83afQGUC3RSaF77Q5bZV78Buh7KsQtjyuygFSZXPihYUY
L79aWQGETbfovWxxMiM96PDLPHT6N/kGpb5F+wm1NSHw6u7QOLNnJWVZOm3B2r9X
WAXaMddgCpGb9rhn8syaPeOrZMC0yZvI81Y4Vh6JtzIQjN/iBJI06mPY4o4cs3+u
gCwwrWPFiJxDehWL+Y8BFLeYWwuQIrDBrBdRNb9CjKrXfu59XKlx0dBjU4FhNJaG
2LmbZh+Hsw8J+rnv9S3zuouVO88DrfPJoqFaSPsMwCxABZnbU4Ss/G9mOj/lv8zO
7eN/a2KwdwtaGac5Qt/Y+vksRZXrQE7zyo/UbU8Ba3lx/gDmNbsVXtfaqD4vtNKg
afbV0/thOy+JncETyi5sq2LXXUsntB+y0W8qhFItjmYvWjN1s7u5rEDgtk/glE4G
j0FPjlnS1ahGQcpq95OzmVV9MyWTMJoDzQEWfNV6bxufH7yfnSHgQYfqDAokWESh
C7FUS3ir/K5ZLfolh2uamhOBBIuOvoApJY0Guy5SXxH84xgXfExbykee/ZwARK/m
QOCHeccxMzRV9Rhqq6mWL41ppMx9H9CipfR8EmHPvZGWFW7/0i3KTKqBuWEfLKW4
Mst1SEcR+Q5Z4NFPo60Vw0yeQ+ONJFm9fMv8XfMSHuEsjzqXOH3pn4Qu7llCwA0H
2DjbsvDY9POkMC7Eo8+w2xnsthHtm2h9GyCKQOFJnnxf0nSWfS7C9OhT9lW/9liM
0nRo5adzSNquXLlzGqUb2OxHNAnC/Au1sBy7mruJySC3Cd7BkPK7CFGSIyBm0+Od
4sI54+RiyeYi733OA+4TWF4cYPKixjQ0UDuYvfxmm0RNmiyMm2ZML6eZ6cke2baP
SKucgD/efRcInD67tWD6NmsIXxJuxkux1218htr65RtKeXWpgyLicU51fvOQbuFF
oQq3bD9Y2uETeU5NJ3v3AZ2N0LPigbh26rmwGaOpIXDWrGtNR5f8Ux7zp2WjM9CF
zITkPfxS58VkOOHi1rMdQiXHJm14/rg9kjrwdi6rqq+Hp9gjIEihynq7QbeDtzzE
xqinNyjtvRSA0FItzgRdOy7XDzGx9sRSjJGmjbv38UV64xvwXbm1PCoSqEaHZseO
W9jxLcrtad0aywVxRj59wEKOE+3XQ9gosN7VpE++4kTDNbebB1ScAr3ViR4TLSXP
b6eTW7XaBETDFcOLu4mTl/SdwYxXSXgjkfgvi4UwhQRePQv683SDodGiK2uL2jTu
r/wXTbMLqSjmew3aYktKL47FfopeYNiMbQBb8p4Yeu+CsthULpYLMd1QmKTks/oT
miD8htt+uA0PoRkWaD3fAFJXOfRxEnKgYHQ+4W2R6H8LFEHleLsHyhrq13aRBdpY
imoRQrDe6t690UroHAZHMnvW5Nz94Tm3G79b6iqlr2m/WLWMSk34VRMbbxXhQXG/
N0yrWmOKWZsXq7v8IzQKvTskkOYOv/b+errQ3CsO06fn3sOPG0E6T64Lp7W7yZlb
Zd95E3EtrebhJI5+ujDd/VJM/aRtLmTf/NEVFuE3Tsb2r3eomt63VU734I6QgvFX
Gt4vw6vpwo6PnkmUf9EZLIYr8newkv4P2SUPFJhiiM+doiKjyF31S0uxViNtDiKz
kmPf9Zh4a9wPKYSeGA90CMigLs8hsF4znZoTxNVJgqQN//OJcLGV//AbntA2ti/Q
2TG/cqt29zqKqUS3H2nEHFZtkf/ZQucHEGXsvHwMtrhIuD58zK+CwJHSFthjwChm
U5vRxbPexnW3mg8iwHkUevlshxk2/+WNqyU3FwxXiNF90qiVE27hL7SjRUg8ngWY
iq1tfmGHElCaxoUO9N8Ph4bKvfXwe04lhBpcYFF3OFcycV4mr8SM9i4IovjbQeew
rKzxC08D7KXGh1ewXOas4GABUs+JX2jNKI0/TFCVQ7rlpdQIlnpnz8YMI4RzcJoZ
pK9li1m5jmWiPStcAC0u2GuNo4LrPZvHIQ8Eglsspua/xkc1m9iz3cGhqjekTPla
6yajUAc6zbG5sPufY96VrJtKnV9Tagau0aijQr/mD8hzIGC023Na63y9gBgCFh24
CNgF9j0+5z8ME3vJ3OJH650yB72ojSEjbOAoaKbt5pmELFsBOhe/nZ2+vQNrOa5y
g5Yj13pXASwTTrsfuMDXJnS7apcnV35/uzGVEFRWZGtJbC3cOsJLn3eyhAZV6VCo
SwRHJ3AZbTJkAGW6XpsLH9mYZcVcbgBI41hhJcQam1TfcueBjCc/5Sa8o+6KBcJI
BHWVHF8RCI2ScM6svIGst5iX2YTDLLGUBka824a+598aDQLASA+h+x2NX3+0bj3A
85jWFBJVX14C7j3DoCS2U5ucNy9VIya2d4xJr/4AkSmMEEvU9hrybmCHDz93VuXV
OuYWkSbkWQN+Z/CMgQo4xS1L/Q6WxJVfi0IOmvaZ0SHoXx7yTTtUO5icWsYpJzgg
4M0yBYGDV9Pf2XuqLryDcrJh3B91jZhhTZA06axo6wFrR4n5ZaMeju4dzw9ifohe
VIvYT9JeBwD4pXzvj33xHTYKFZ1ifRA6NzVTvXkCv/h5CE56we9Meg01/CE6t3/D
4EEoPvMS6rpTcpQUleb6PHjU9Mj4Pk0E28nize7auwkx3YEMMpkypFtVNB8EVKdI
Ulf/NYv1T+ku8CeEMYXiCCi9k9n25jn93EXsPA375S3a0vW8JT7h10dg6PT3jy4r
e3hc/ZOP9xHx3UOzWVkLG4En8TckttZcHfFxcBIQKKUNTdlfIiEHCjXpyGdrYfYo
nHVPNzxwreobB5zjKSpNO3yEVzJIlrclObfBl7gIQB+7opr+m1O1TMwwoi6hDdRl
gNzH1b9nS15wDu7ss1HXuRaVSey1o+iLAveu1EiPlyte176DBhVWveRts4ti31Ec
4k3QpQlM4iSPVjh9g6tBm5LlvpNxd3pDw5RJlak63GAjkQiEPwVmqxUmJ8bfRsci
Ue+SYsESJRl3a3W4Xs7DQ6Lei4av/pr8Wi4idPOi479m1PI7QUmEMKtKnAfx43rt
+dwvP0jdR4x67iP5HWW8jLuN8hjOnoijG9WiGtv8vVQrHdshae8kSznKT9buPB1O
RxpE98faP9ZzmQZmxEyFoh5K86BWGWQ0W1s6sBWdRWKiSWACl0BUOzg/x7Pz5zgP
z2IdZ7fOg9hfXp3+PQ9PXw0EvYOeHXJc3Lpy8gGPbFmSHgYe7wVgHb5sFY4cDAP4
g7ZCGibSfwQXCTNPq4p9kHD7y8vCeWOBv0Nzntv1WoLsXg2B3FpOpLCT+iI7F/9n
ug83trZMdgFt1IONUvkGVCQYNfY3AoUQYsAWPwsn89gsiUdlFhF0SqSoV+o3s6TJ
fQUu3KMsVegWkzTBb2lOn8ejBjK4LvAwJ5BeD2nt+kz6OUHi5nuY8jbtmN46fEaj
cs7dVq01ICpyp03wldcu9cyNPf/+EJBmCHHI652wksk0WsriRO9C2JGjiccDsZv6
cQYWqnPJrD8gerDo7jUuuJeUcIVZCi1Op01bwYdz6EtEowqWXGnavR8UCbfhCKu0
jsbiSQQoqxFy+qJZiJUlBB5xNCwS7Qf8ul7Sn9YK070BXl8xZmifud78tGduLZNL
CS4GP4gghKxaYE6qukOdpzJC0KVhcRBC9/naGFf/tRHvwl3jtwWFedlxrTwPjo17
9BN5GifD4tweaAKm1QJchj0nqf9tHsJzHIPtMbvYTwOhsE05UB4Qm1pX+IY9Azi3
UFrOUW3LallXFKUUP+9JcIidHmaU8xII3Ip0kGLbNbNN/iEf7CQuKg1JQITtnrDO
J0AD/KJmBwuO9aHnUIUUZk0x6lLFkxHW7M8N8xF667llnkZVPGO68VZg9pv6y59e
qaY3i8wCrsaRUyqmeKPtQiCxEbg5rCCR97Zlvy7pS9yCxxlVr1Zeb4WxqZnBAiRQ
SYG5QTRd0IudoaWG2FADM5XKh8Jz5/mqMxI0n0SSIgsef/3Rb/fMs3+9seb4c6wq
k60tvHUorNV08vM8eHUDPq6KC4AUQIwvAVAqu+z7aAJAeRpHMEZv+9/fb2eaKDFU
NAC5clODqFGpow6umyr76h00uJsmCV+E53DagZWhGmHCLTxUUdzL8BfEMyWoQU9S
tmEBJGiIIymX8shwsMXEqcec8q9k36oT4rIonI3P+DAAk1i7e7g141z2HC/eKCRO
hALSciFzBCqpa6kJXlZ4SKmv8fkGKT+Q1bhKMk/Gjv1DQvU2+eZkxwevkkC5M5n3
UrSF/PrX9KT8Nrpz6iEltVBib7+XaF42HOF/DcU7T3JQSdKShobpKBHMCWvttXcl
E9glx+rd/FZMShnLKzZVE9O4qHVVJ0y3aLnK/KrVsZzrxcVok7wIUkejz22CF5N1
tWxqOLsAYXGeXIBGgb5wEC/xS3NUyleJwnvFVo0tTHw8KOFNMH8duTuFHKCaDsOM
epw117X1GEe7x9S2DCFe50ZkB3xzsmNuFmJhniYUvaO/d1dJOcPuw9fV3b/LtPeo
RfCPxDeKuCCbL/uLDCWuie3OC15QvAMshcsTXiOaM36qFqCeAJiGV1VwEWLgyJc6
w7uBi8dF5Lw/qaLt2VKep1U7VKzw/cTEaDzkpY+t71Mj52Sa1i9+W1/zscqqXwXk
3QDXBy9rqsnle7pNrq54u1QM8CN6idPmqsUgh7BKSGRSQIkYV6i8ojsTAPUKktJZ
fCjZboYe2Lecqoik/0ooi1A3Y21MwjjK26c0j7bs7lnOGZ0R9Diy0Aup+xAWrAun
+kFVdx0yU/zKDar2VIlRzqtXAEFxwS/oxvwbA0uqbm9rSE9g7rNmJ5WpUGF3GG6g
BQYoUaupKRRFPwsXk43Fa6kBh4ftAtHkhFMbtClZ4ek4UhRX6MDTqQv+IAqdD7/9
vnU0uNk+e/8NfCnWU0SpgpACvC6pCUZnG00D/edlpx7BccQVJk81EPfhMDXi2K2w
4PzGwJZfVsVyUF1bDEWxRR1VcDTdH9V2IFeLu0xxu8Iqy9T8JsSRUwZiDTHz9pKv
NjTUD/dXI0FFlVkw3TrNgTEZDnmWNgIBCJOdr16w3vnKDYVLfGidVkpAI2URRpFv
Bn/ivKYQVpU8FuIHA5ehK5lUeaQhSExT05VMIzWHmEuKGzcfupTID686UWpAFn2y
BhJXDhGvUQIkV0zwUHRusJTgIxxUiRyeP5TG/X+Y2cDW+gJjXHna7vB9qDZvSax8
rzjn6mdrIFlO0u62yUFfRC00GHV2trkNPGVy6ILZf7riDAgDRNnaGaNGzqD9hQWb
zlqIKJRyudBjWqPord5Gy5xcHKNRAaIDuxOd1OeY2Br5ZXRK05Y04sHkF+ChiSFq
cow8ATftNCc0l7vwgsNKP/UTLm6BJzP6dsaVclKTSSEtX9IgWzrCX0sQEFjOCqE4
Rj8Lxu+cb0RtueFltawTQA9Ex2Jw39wdH/vtw7GCcS07vhyRa3AmAvsUZeQFEkUh
jcXKVJBFvI/Xc4qT3IC2Ij24eidiwYYm2+N5pHHFqkgbM1PkqEGFRMU+tvzk7peV
cUqXJmUcmD3OyG6PetO1LX8CX/raHC+65E8cSoitzJnT1/XFnf0vDpNpzhpVmG25
H12pwKxMiZMupm6CR7oIqIg67FyrHB7MvxS3VMrDmxWIQvPBMvYWv4Sk1hqvBX+3
jmhtL52+9BKeBKT3ooIdMFO+4CH3SJ0+acSsfRD7Q9+HwscQ3qajdem2foNsEBUw
sgIB1z2J6AfTG3kuUscwmeLdn6FveH5OxsamR7uOoYgHkufPuP6+EELo8hhNZ98N
m29EBXrqRHVLD26PfmU49t3AHIdGgnoA9YAXCir/qnUhH5LYDPPuymJMoE9tb/bt
9CHWGaA48CRzCPz0oocd8e6ZuSNyE+z+AwwFhYBh3Y/CVYPw/dxdH+WpHckjuWCR
disIOC8556s4YyrZreMc2WHSAOm2fjrqu1koe+SDxase/TWx+9IOQW09ic0c0RHT
UjybKV+wnIILjcUpsPTxgsQ3nUk3YL6Fv2TK7TGinF/VyPL+SGez10LxyF8t85u8
P2y/6MZaSejguunZIKpNzmqaZn2lV/duQ4cdqdx+iHWmcNlosFM0xOHHwN+cdHSm
WVmCOSN5B3RuZLB+W/GLQ/CKSbAGb7qMJUzxGZdN2KTAbij5GOi+1Zo1XlHm7L6e
E5R7PQvk40tb121BFOOV3QY/036jneWUcvoVpUnjlE82q3aKG2BgAm0MuJxfjUwj
AxZPyzcq3SirA7bFuufEE45bnJ8pxXOpVot+rSOBR8emYziNsoBDoJO/xIgJdBAQ
biB2NLDAAN+ia8fcZNBCJB4KvN8bg3cJ7Ew3z1r28MZi1aRUi0ovC75gzSv11dlx
kG8ABb9QY/0vSYuJAuCPxxIKFNEYuT34fnfepI+R2ImDUH104NTLS6GzgJhxJkdB
2Cs4rUdjROZEPm64/93ZNEvY/QRBnKU0ZTJORsp0CjLpY5/y0XbGvl3rnT8iM7wo
IObtSCX7Jq0bxASJJj+Uk2g6tlBkuz2ukYs66K7TpEmkAchwPQpI3aDdB49XgkEi
aXb9aJseFZmK3OiJ5y902oxDyNTQ5JjzvWWh5jVi9hqw7Uq2KQ7+P3pvNZ6m7yMf
DyA+tJaA2sNZ3XbdPZXgfeHI+APUFoeBcz4XpW0wkAwq/QO2WA/hAV/wAFnERybc
MWlWyEm4/OhJR7YTOFDqYiW5OO/d1Y5M50gMckNE/Mu/ocpeu+PmI4Ga/sj8m6Ac
oGRM3mf6Ms+ui9AttnGWQOBs5sKqkrJ2ZOLo3n858Kcq1MYgTV8ZMdpmO2Ut3u5a
QRVzu80RtbwI/hHgXzLoPmCEXkmEQSrr+6b9hit0rn7dgCo/hSTvNQh053vD2gfi
HSwwJ379EacTtU9FJWmzLEeEPFDGbnBmRGuLurUEypk8QgApbZ6PUIi3BDQR8K4Q
hmf++xY6Qs+yeDbSW2usFYR8Elzp2kMWQMT4kctiBe3HclYaxqRqi1tNTaGkvp9m
YS3A3qhCQPO/nmsw7bsiqfAoUvxhWyyGSvYeRhEqZuEHg2EXI6+aHJHPdGOpBp3W
OmlwAG353tVXvmdpm/UwmyVDXKRukoki4cawsVkuJRABRdWOfM+VOYwe88Wd9/Ii
iw5aw59XkjFlpgIaEMuvmrhgAXgKL+MNFddTyHmK0SZCxlMiNmYI6wkHdMto7SvZ
TwGc9yDyOfhGlYfIP1xJdxQz+0cqOB4G0SHFQhYvGTsOybP0vI1W/1wBYCTfdrB3
ITRweIzZvbBM4uXhWQv59Qg5L5PsmfB2lcB5TxGDuJbX26ObeVRsj5bDvEfugvNh
bdHYzB1BXFKFZ+FIQC4JfVSLA8lYENQGVQJQizY1mNrwMi00gBRBT218BID6nCvD
/c1hoZEwHnRn8SQBdvIlxM4qwC3KFpYWj/Ec6QxBf6lo7ROCnFz8681LvgFh5rl5
kLQXmlw/TyZkITmQHmz4RJtiSJ+77220OoU1h3DmJYJAusPYs1xc2fJ3QTpjE7+q
s/gQ3wZr3Z6Pfa1VpWsqqSxohyxrJPjMqJNPN+spsZWS8MF7YLlxXP24HJ4IoE9b
IV+ceictO5xd5u/cgN2LGNokrsPDCYQhni5vnb605OYcmtJ2QbCs/k7Adwl6mwij
CYb4oOafehfZIOZcmOwS5R8jJBXZGsE6If2ZBxJRomqQ7/zS5vQjoifgHWSh1lWA
TY9PT39Kq3V+QIwHTI4wgD5mRd56RjDXTyFNIPw2onzlc6x5IW8thpfNFaHMhlep
MOIvyrEryMYQ8hfMAlczZWowjOiSJBEiabyNSeYpHRCx40VBUYQGGrzoN00PvscJ
EAaRprUqST8ZrplHVDoV3ld/z0sapa6RJobuPnqfjlXgY3w6ryArpUZk4lzb4bBg
TlqQTK3KDv+JaRnbekVgJz/RzImU72IsdmFm0s3RurNHT1HdtkE9bRM95+Rmwy4n
L71pHDtLE3Odskfo3x+Zx/DwP48O+OZE5Ei2gqPGpuF5iwYsOl7qTSN1MY/lBjbf
7NnH/RKyPrV/vJHI0/FM1JnlGYHX7GecQUN7DhIGRwLcHewMgoLywigoNcVe6y46
+oWzxFqPk+NdDjmxaAW2gGvO2EjvngumotY4hwrpNHtKnelWNkYHUFq3rgeAFDuK
miMNs3tiMRZt4o7gUYs+ffKEkfaJeizZVzTT/B5BoIe00UcmlX9kfZatvaPjcC1N
ZoxVCSzWcgSzsiyGDNOjHv5LRZ5UmjBP1NaCyaTF54CM6gPcCoisbalsHSsjIokf
7Fslhwi6GtD38xrAJzLzSP9ssWAyzCCQ8XwF2A/oyvrCZT2FvZl07W18kyy8wS7M
QTSPFUscR972VXjRFVVoVRrh58wjczVLK+ZjqnbyCSTGpWf9iO7DH+3RN2qrBlaG
kcCKN67jknUpnaQLaxum2jRwhqJvQR2/L6CbkERxxtJIfNyduhDJeqNG0tl/BP8h
uNJJlCRFm6FgPyDFuLmZZF5nqrcRVBYtZm+G/lKW8ZT4XK90uJw+0xNgXTOd6e6l
f72U2oz6+Cilhuhiw9L9oArD9YP3isFdYENSYEEGj8OeHvC9IdoSseP0sAGsEMsc
mXL504wNS3NeQdsGG1J/f+q9PfaG1qAmqO2HQkW+4895DR7g6FXf5dPH8Rbu9Ns2
45qZVhUodEIHe+9qfBDkxwf1RSjGxLcjlEAQMUGGVZi4m24zW1uGXtmvKV5L/4Tm
d6YAKBMQzaLKJpzaY6YusQLJ5+cePmyuqghQGycAqOrvN+HltEgrcsJ+7QF1yn3I
3yx4gWjZ+qFobf7aeTdjoR6wr8EbD1JnSOej3rU7SG2UPEIP2htMbdG81m8wesyo
/aL87LUXJLbvl1WRvKUquY78DCYedY1pvs/r8MT8b/b/fzHWl4Op3G5fT124O3af
hxf8YRwuvXAgzsDTWHUNdrfhFgkR/BeDrq9DJJpeSnjsiEHqqRH5g/e7mD3LpGXw
Boc8pNalORleKkvsKFJC2/hcJuInQ2IPLGyH1blxWlx5eAFKz/bDRjL+8YeaY6ud
WN7tytt+LP6Qy4kedkOwusjMJCO5R749gaRQie11g0dAJmgeL5KK1TaZ6ouRG7Xs
cI5WiUZA4FESzIuphnX65aPQqdnJsPHcWieKKiH5kROEsdP4svYZRF7ms/iRkXRB
poAfu6H9IgZaKM3LoEEKl9MMDP1HNuyz+m0nYK4YCphCz/dcvnXfVtJspua7HDnb
ts3gYMMMZL0CKwv45BbEoS0+TFx1kNl+mpC4FMUw4L9kt94BtFLWLNgCyPUJRgXS
FJ5Tz257WhFxk1O7NgY2y7Ac8751kAUSLel7jdmnonyQoPNvYjVHl7H84hRR0L5J
LwmTDkR76igHu88sR0EWt9/t4v1gV6XyHxJtSqvqjrDyACIbJBduiRrLyIZtdAfv
4qjGI+0BPmKNYbyJAcgBn7RKgxvyzlx5qsnYjDFhoSb+IIz2EbYKwoUeahTyyk17
b+xtA6KC0y01iyL7yy+syrxQL5gPOPgJZ04+InA965RtsMNJrddzLLnPJIkLkk1U
4o8O1WB3NR3PMPhyNR0iY3C4R4ITUOAKGyo0/oRG+oJQFZ3PBtYlRodFHplbVZU3
09e8950L3HECL4GCRVtGJz9ayPOVs2bEvtjeiryk9OW673PZrejsiZ/s3HvlrKQ1
kKR7TuIhVkpgZ7ETrenmN3DQTXvMES42sFwhWTmhMSIPWRs6ad8JTHBwyOFC8jAY
otHwvFCinm90AcV07WyIIity/FBiggQAV/HfEHXKfgFcF+9UHj2kzRJMzwZTvDAl
Ba1x67Ub4do1jBK9PQyU1sAG39UbQ0Z0cXY0o9MO6mnq0NK9BqBOY2fjU6EFcjEb
YhdrpffyN0CMRveFiV9wjrEqRGCKiKzCMcjdHgvkFjK2Q30K7TJ/xYGWSoZpNNG2
PJlsrDkLjS7jL/UFM3ezIM9C4Zzy8qRqEjZUsEtjsW1+Sg/md4o0jfDnL/WJRArQ
TbiccVKBOBaNSLZ+aV8E036BdlIECbeUeiNjWt1N3O10vglXGO6omaq6wZMd4/LH
NVL953INIG/tln0t+LJhQFQAJwumT/+PKqSTDt2KQMZ578rKMQLEfH1u1si2NY0f
UvAbhzSUKlVN8a13uz/yaOY+aSIqhjST09Y4PlJcBC7cebI61QVQS47qFlNHO/QY
+EpQgvqf/KIbHuFtf+BSUgjfQL8RQpXKLxgNofVfrHsWeFVf5W37N2A3wCCtJOcH
ONpQYIUVbVe4JWZRbVNFBm/VjaDgI9BWHFBbAtGHqATUUgaIgJdPJEN3W59NdRI0
sfKvf/En3SQNrBetnxgUwMFgbpmOSt1V4AbEraozRaWvSZCB5YlGK7OUWIAe2Y9g
y5n6EQps6t8YEIi6uO5qezdTVM2KmowiK5+0eKqSbXaz3yrys1h+45OUA8KJeyHJ
wqfRx1adxwAATCxw9KmsaMmEsJidvQ/w4Pg7vgIVfKB9YSBKYAoc0/cczB/v3sMg
zoFWiOHDJ7XjiB8f2bRxhasz+yqgF0iwfU0GaFKD+kArkrWZS8RJsxa2k6yqzKZF
4RkaxDAyfOh1WXeXOpHTBovq5cRTKcRXfd7xA6KS+V11k74bin3fta5gaMu8EeSU
rEFh9cSpJ/IFttCGanc0Pw3tXHZaRWTVeSXKjmAc5U6miuguG2v7g9mjxcN/dO2K
5zCOU2Zs9Lwv2vzWvGRKYeIR+a94i2e3JSVjDSQZC5SQlUQ5v3Ab3UguAbWm0+as
PYJLzITLJ7LoXiuY19y6QlyPERTSiP4w/qv+o3hNuwzTS2zSniqiFlrCYohdQt06
qW4Fn6QWVWmN5IABcffmwcAdh5CGiZ3N88q0+j/PMY+HF5L6OTReu2XqeDFEaMm/
gmDstAtMky6CmPerDGLpMqLGxhhhyWCfGn4fIHyp4B5ZCGTsFmZMjqK/tLsm8YEJ
NPJxRCyEykQ4kW+Q5UpJedK5hu9MgH9FN/LC8pL29WHjgaZINH/rLBrm+HnNEN8k
IWG8+No7c/jLcLtNDbetxmVRsm8qdpqQ7gIBt5/ANITq+LikwY7I1B7H91XGXyEa
+UCfynXFH1DYmVCTyu/igTdhv/4Wb1gV6rrBI2mNLxxozIr4QpZN8xHDGLfHSV5U
iwRPJGzaurG5SWsxHgXaUjF32PYUJYOJwpULVq4dQZdYlE/5Azruu+aiUx7d5xPy
LHd2tk+b+9V3FI9QDn1atwExBH7RGugFbV4kY5xZbmhikskwHVCoTIpE6it+daJS
MbeCvOzEX2gA+SfgNYLeC/q8tDpbUGC9nqZD9JaZ+g2RmvR6G1Ne2tvFhA/usMXL
7l+VSA0+5DomRkHaSLsoIr/tZoqARnBLrhdFFh/lQG6ktODP73Yd6xVZVIAvaJVh
iTFYQrNO2iEPsuhrXTPzMX75QBijECpTkR1Eku8oFVrv1AB8G0aTnDUT+MYym1v5
UfCnJFS4qfqBL9RF4ItrEpwzwPkqAF5mRdCetczdGh7F1ZkZYRKWL6PO34Gxfb/U
KZhskyyKZmFHBS/0skb+NxkYXLaUIq9Hqygd+ztbaLg6oKa46JLpRVSBeLyZ1Zmr
GvXUsSgDZ8Rt3VNm9Qiil/QsQTu8Q+TXFKgLQtiVIsXQjrjEcdF8klfXDoc1BGxK
/0BsEil4T+t5yU0jsg/otoLW5VZQ2FMqmozLLwjJnFA0sEnV9MJaPqikwUXsxJ1m
7uU9hsE9dbyaxSQBnBitkb3iM4EJj1WXfSC/qs9iZTwSFCqzmzfcanKECLUxMRXD
vhPfqiF+35OwLISYw/EV+TKxOBSWaJi/njdycyxsI5JIxeD4v382oATb0pCKzJp4
JVL1RsDJ7d1pMs61H1muFEkcTR4i+vR78H1BTHlZH6AkKy0DCaUh2X5zA8lB4VTK
QWabPvtPrn/65c8MTENFvlNJJk1zFu67T8q0zmw2lLW2FA/Ruw0VDnI7MGxjHHe8
+LeUPGE5BA0Gg4Q1j9SqiPpirYrKfUptd9MtYpuOJr/b43uj9X7rouyrtjH52Ry8
kmnebqBkaacG1qA/CzgXc/5j+iFo6BcI/GfSQTFrftP0WrYfMGUDsSL5cnbMo6Lq
R6Vra8h+bbpWeVVXdNugN7tVxt5cEGCANGQWLcnggXoUSo5qnO3J+AKTns5Fws9f
o9ZW+rmupqtGeBk1my8WTVKiXpRP8K7qfKVX+sWL7n4ZQH1LMin3UTglgnU2c/O+
G6ux2eCrpTKEHWDtwirHAARbjpOEb1MF7zE3++8PwvIne1oaTot3sRwz48SFATDL
tfXOPMMWQJvf/x8YKPqci5G2BaIdzk1WQ3Bf67HAyFWSIgPS/ZJlaPpAdPtZqqki
XGs9yOROVUDK7/hfFafi/MSaBGfkPGqyEOgKoLp5eaBVvAgtk56/CMTy3Shy/nCM
VEx7IPwL8rqhj5bO0/M+6rRgfmC31vJDne8D32455rAgWFrYc/D0nF1Noway5Tjh
YBSDkTpiTmhCXczX7ppI7JbdnG+A4FUlqR/nY4q+eWJiYjrOFjzVTCUAmuOH8ixq
JcpA1R0wPkaRwDHHwlUgnfNZkF2CVS5UbRkTz9VtMaIRfEryy8pjc958osaVHG7w
sn24FXZEnSWxpcvaVGN0Sf38Em636Nb627X5kItxDq4svMr/qNH6wd+8Xsh6KFdU
F4ekAr8gtRgnqsg1w69X3f6oOb1LNmcPXGVxNzzedC+JhomRPMgH++z5KSt4GvIa
vJs8cpABLNvS6XxdfW3kiVvaRzhL7CfSf1erODoAQRzXSIdeoFBiuBX+FE/HSN/9
/Qn1gLgTYHhPCEIAQ6lNAAu1RAclG8opyOFIPdWEd4zCUK79TTss7mNVhjt6Hkgk
iHMh4n5dJOLpflTSh7QmyGKr9X9H6Cgoe8uEvwt1kBuM9b161/c9xjFG/H2FfU/p
CvyagFGXbjrkoSF+FsDpFxKKHh2jMHKabWYjns7JXYl8E0hPDGzE+HmzIBxzKQsF
W5Bd10SKUmVEr8AUiESt6MtouOiqt/eNMqU6o2n90AfJTNwwXznJGqQaC38VnkiM
1SATq25u1tuB0zUMLU7NROmsjEeYId7FM2tSHgU5vRlgh93yFmmSds0h1pw5m2pN
Qm4qBdd8Oc4IMibf6N+4s9+57GIH5hCrhwbnAr8Tbf9CNbKbRh+9pL0ZGsOlJ36W
0VUOb+NXrVTWm83oOq5lstQIrMB2i+fjj7qcaMq8QoLY+Yfwana1xOSv5XfetYk7
ZHU8uwrXIvF7ZjPPH/9ZcUv6lP84wvnk2Dm0HrFuMm1XkkCAd3CBC09FBbZGpVyd
E5Jiz7L0vhG1mxiO287RfuvkORGY9PtByC1iUw5uP4h0wR+c5d/80Jj4bwbO0+M6
z47k48Nw7bNfFDXdkwkDKn7osvDxfF3HO98OXqwRr+k2xVesEbD6F7rOpPuZjnGk
NlIPJOCjp+BPQl/ZL2eQYvTGvckjETVKNPo4g3JDWW1qVclHvJxr6vaJziu6GVn6
l8YoQdaFLkL84IVh/vS/jH52cNYrZxnSE4Ik7rgkDOGDMjCmp306bNga4vEo1N2z
/vl3guyxIiFRSyjKu+LACIqzxH0F5KmBQ0ck17/BeKS3ilNnWvV+kPvdzJ6FADkg
OARXAfBOcA5A3VluUxjCFxRoSD6+B80UE3f79VVNi7KLA/PeCKtCl3CB7Kn0ZRJK
ewhYOTCdExGjZFVrdn4M+4qw837na2V4eRrCW7X0aIibmPo1xW10yhjaoRcQwnKH
lY6HcieTZSpeE+IZpvg44gudYWNoJgwv/P4jXeBXaQiVnBVR4kk7bCY1z+GcddVi
Falnty3zuMjFXcjOuGm1PiKJr+v37HNSmHNdTdlUkVnkKaQhWxA0fqmpoCOb97gX
GnOk79E1SfT0F2fSrkb48tGhADfy5lRt0vwZsbPzFvsn1IeFW0mySUKjggF13jDL
E/RrnDRhPnLGJwiidVIWpI6HJixvL/ulflAyvWR1dYdp0aSE32Ng/cqQFXswSC6/
D/JVqzSjKChFYI/xYcJOsG9ynEb69rlcF8iRG9FK0knZN54bfg6GKSVAH4GNZ7Ru
n2PEiPzTpcGCMixt3/QgAmccIDfzZGWVefNbxW0cinzfQp1qMKYdQVz1z05Mr7z4
Ma8o8aMCdY6ZPGZppvglfKobeHDdniLUS+6Fh/lssikN+YkB6+rsgsuZL0b8Fjwv
lD5qK+N19AxjrDsXDbGI+6EuJM9/u/fUa5hjXdsbP74tITB8ww+J71K8WEGfYC/W
Pgxm3H/Mmtihakfo1EkXtucX+D6SoBz3JP6/U8OSHSPeouwxSoDGFGcyNn9xO3kT
7GbTnx3NR0Kn4q50K0sLKI5DpKv+tQC902U+16wJNuKjEinDKguhd4169kkEkw4i
HqLesF2AZfnk/kWcJD/L2f0PNOqxuUZJXg8N8fEvMwjcTlpFw0vsfj+aesHbd/rB
bsXU9CyUKkorLtrI6t5ABOVbwpaddVEyYV2N+cHWYDwRHpxerO5/427MWVkT1zzx
kIR50+g0Vuii+otLbBeAKfCsEdypG00K1Zd0Jh7vMkhEH8S7tyxHVnmaUdeCqt2q
VmwGEDoMk8NYlFAvLr6KuwOfAyv5PmE1FuTgknasoOINxfS3joYIIQmuTwvUpjDr
RAgO/9PQRQwAC5KOmzs3b4OIg0TSCcsTbOhkbQrDpj6fAq8/lGQjCuuQTFGilYLp
S+4xU16M5xY4iLA9Y1MlqgH5diGbt5e/PzQTMydovE2XHpXwFlAkbd9pYXE6BKF0
KhlSHqNpfKJg8PrzaBOxpVEavQm3xNTysamfiuJmMsGTjaAPHXIV4zx4xFBJeVec
TRwxsN7x4U5v853YAK2DBUx+J1itwfUokTFw4MJWJMz4Ef9EZYVWH1VRrl1BDouC
GMgvcdBkLe0wLilkEsN7KkAlxfxahzHt0QqeCWIXNWF7r6zTIjcfTAV92qBjPE7P
eLoKILqahXg3vyuLmEP3ajdlR4q2EZ7VFB3KdS+MyoGtG4vvMzmNJktjodmb4jp3
26c9U3JGkIKsjhwL198BCS92dyJenYcXzs+JSD/Qd7rZhg18uvd1d9dWVarFwQYK
LRizNU21fchbg361OLS5yxiaWKEWtSqkyYm7PfVeUs7ZYIJfRo2YqMjuTol3yP8i
oCwno24hlaMDRDql1hiMa5oJNmOO9QyWK0i4CeH8nnfqU8RacTEHTXP7KJxmd00j
afV7svkMGQO+5J4i8RhnSa0FKzfPC9w/+pKCiZ+KbNpiW2Oz79JtVcC/1pRZpRhu
Q4VXWbJr5WOpXYvw3WY2oJ5EPlsGiQwO06YMWbNCNhAQnsCTAZjwSY25+gfpWnjx
kLxvkbTuD2j4MQ4JVlU6ovdXKDKMMoFTgx6Pz70w0cHM6bYE69kVm7Cfoq5LrVJX
nwFT73Me1s+rgf8HZEX4aMkx/iuasZAPV+TjceNHAlmM/okFwRuvY4zCXc1xpZkf
0KPNiYjYtqMTGNYembSngvpyxH92c8+uEgn+RgHU1vxxdKTG79tFu7YX3I4k4tk+
4lJ3NWjMU1umKmSFbKjxqu0UjHMD2/vQ4mcZmeS36rjjPA+5WO/QHq1+bdODZYpf
qK0vmNH/RR/QDtRgmuM+guWZEYYVYugdU/PhvtmwTAMEcyR1P/fkG+de+fobTcl1
4/Q5FczFRVhjlTwfXAq+As8YcLtsUvd4on22oPtkASahEm4rN9wCZ7GZyFev31IU
7DSz10cmdU6Ka8jfEvKJTktixqYIulGHbuVYm3OvZaLcbjukYWPOZzv0TC8vk+Fv
bkN1LSh60izyCVcinahSgOsylXiUntJpk1qCJ0orh/dvHjr05nJLKsV/jp/NQOj4
fUFSgEjrHubzPgQf8OxG423qddwh26uYggF6de6WsN1dB9Fjw3EBaz+JDk2mvLeD
BuCUVsMGodBV9uuDG64+6F1q0jvNE+W7lsWmd715kASi+HDpDlVFG5lbUhh2n7Bd
4gWx21YxwvGp62Z6N4WS2orvO6yKL+mOHX0wLQSlME0y9H4KrYhWK1VaAksDGDyp
HKF3S/Ig2anktrkzDI+7VdJivGAu75RL6CTd0imVY2oP35s7UJr2sH+vLYyupyD7
ifqprE8thR2psjvaaEgpYoubkxpB0KbNR4ETovEZBVns8GNYuHkDJd27O4Y+Vxnq
f2cKUJyQnaL6Pys3puv/4l7vzhrUwe64jHfuFUpgZth1WpmRQsW6Kt3Lz+vg0cQu
kgFuMzjpzB7M+CPfoKUj/mT8ymhZMwF8c/kScnC14jRaaWcmAaYGNEZzoluApAtx
cr5kE5GmJWonlmVLVIN9Ib8d8XOe7nwbiLHVlToT1QKF9R/s98LgOpB3JDPqNnCD
oVZd9BPUAp7biufMZVBam+IVQLtCggvAUuhlUc6kbuToaJPsBnfO7YBwkXO+IR7g
5fMcusYczhpwgBmt73tRaJtW+OU5UeshFdstHGCindcFKeWQUWmKn7zD2vTkDtLr
owt8Ky4iOjILiWe7FJoMHZo0rUQrE2gBSkFvfymhoMoaGTnbV0QDxPaV5OTYpkAo
Zx6e4lf9D+nSxV07EjpLSin0UiDGD5fam4GOCCAroLh+hU4Fj7Gj2WTeIRBi1gP1
1W06IHWCB+Hq04j1u6ES7CQ7F3FZcGFWE1NhUGuN+6NVOeknU+j151VkWxQuAw25
QWR6Pkg8mam/RxvhgoeTBvZPq8av7274u0ZikZDWLFu0lYRowC+WUlx+f1UgPxIh
HLsS0OcttPXsaCdJRrnlpPJO/hzkx9TOzEDtiJKF9XXNz8fdYbYQ0dxEo7u8VOwh
jLsZJMsDYi4Zx9KyMjLmYAiZF7utRf+/+m0cLjNKu+Wk6Hmh3qivl41TQieEs0Sd
X+uJYRqgmLpygkllvxQRkaPbnb70dtAnesIza2h1A6BUcOrKAcp9eZR2krCql3Qn
RxCkJFPD74JhnmlzfCnJ/Ly+nKc7h1OrxdNCpW2MhGlApqw2jQXYYnquvHlvss/W
8x068pNmvO8v3boeeT+lKq8/mDtniM5By6iILRQMwFT77XTv4IKUq8Ne7wEPhuZg
xuWwPR3leQp1A92+aA4LeYGNx0vMpcIveAUXc3fLmjWbQHb243QYeLvE7zr/qxpG
A0NfueMsgzStPy65/d5v8APlp/0aH46wOdFl2yjKgWRpV7i35sjA+xIZXQErMWAU
dFgvNVs3CBtVmgYsmIg9V5r/tHgLW9yKRnwFxl6rmZA7mZLYmxvFjbcWp/qm5LJO
foZR/t5N7HzLf0Z3qoEyQ2bkpMlsCrJptIgQvv8fS8K7BnSay4tbO9EXOFJDgvX8
s7t83CVzsJtWaXHfxeb+7OnOnmbykql5MK3B0cd4Dz8uq5nl5jsupT4nghcnTXY7
Yamo3IuHUbCaas1DH6Sf5J1pq+tt+dBTjNR4WyEK6SWKWpfpr/oveo+GB600VTpJ
LSjm2wQLXpT8qPNbwy1AYRcC45iyKq7QvwiHyEh/HpGd01YNWWgeoCTGWEBpAq1l
O4zZmOZy6WKrAHa3Y6IKhqgoFrF5X803KU+X+O8LxycSiLf+HfaKh6G67m1irOYM
FS7oeRkFW6dNlbMbP7JG8fxov8f1qkLf3mvGvYuEqPJwdspbjIQrvUG5o+kKctJo
S/vOPb2kSiALKuDIOhpWLgUWsmcnd1kOqce43Nj7nG3uXBPbHKSy+m/zd46UKnkI
PajrlZ9ox0v5sj6Fw2ZRbSqDU2+vkd02VAudjEjd+rTjOXGnC9VOcoi4dNh1jlyE
yrK1Q11CPFOATgJvoTS9mJifNuxNh1OuRqIKL4dDGa6TsaxOMtczj2C7fEcMAdI8
dQku8p+Zd9BxH0lvAs5EauG8Gn8UTpvlwoJZcvoz8wlYmlU6xLYDeLkMT3uTgTih
Wloawc6jfp+/yd6h11QQkOYEq9mK+cAi0Doa5JaeqCXXsyvdNmY1fe3sZqEG3tG9
rwnCmu9LA7V/FaVllZKDlFOsutYKSDWnyyga9d1Z1z791/8Bdf5IwJD3ojk26DUI
fFb03QPF7Wza1WR881H2yyAjUpT7tq6PSxHbzENtgn3vH3hpMLsEugsjHOXVstSj
CZSJERDcTjA74yEAcNX1PiLqRzKs+ZpAwmLYABZQtH0Aqh/GkXnT6WcB1L+i308L
IqkjG9QrbZStPWcQQ7Brt5HALHktCV5XrJlDCwUQn4ndyZnNANuirbdkzyTJ1KhL
BUn3XAT58UqYIN6zY6BhLWoYsor3rrECMXvLppkNqdbrLR7ozJaqTwqKLNMW3Uuz
eTPZE0ChG2C2NPdfPiiJSqiTTduSJ7xLvMA73NwDBYJd5Yjk0PsnSYw8e/I86OfT
pIme0TTdlTOQVy9V9t3N3fL6fQ+m9g33dOgcslZUKQg3a4jwjLv2vrP7UCVfIB+h
3AB+PvdEIpWzYZEqCQB+99HTinuTaLXQ62SsgxRFnSoy6mTR6ZdqltNBZIIT1Qvx
qAhIhglGD1mSbkvC6r01kCF/kk86bW7O+z+Mh1TVzjjAYf8xyZEwlvpYQvlJbuVd
AlQ0YcNy8A8RaBN4habV5RRvbbV1dJbDajQD0zi0AWU6KQyEOXKJRlWrywlv/pd3
HjSFV0SJdCLBhQ98TcbNswGeEcpu2Abws32f5VtH8lxO9I28T4k2gk3NeWzqGzML
sy+eUzB/qXI0Nc45uF5It7vikFLLoZcWsRC2/k4W9tw1YULGEKNZmHev/6u+uXso
6fffPWpvx6WdB9z2IAKalL85xW1AcwD4NZKHsbV50crfUhL/ngsAg5wjrROlasbk
jqz6v1+cOs/4O8ZEIhjBk8YvKeG5krqH1V4HpQGhF385HP8iD/qMGIbQo0eIHwh2
Ki1l/SC31YVjx/CUcArTCi3rKyh7ffMQVFWTJC/PGWosw1Kbs8+m9Z+5jj2bzY+U
06AEAcAifQ39kkrQZQ0JEewtc/g3QO3lUFfcFMNj8TiNkS1VCYGffgy5N+DmQVS/
B1ZgLErq1FBAP5zuOVW3FvJzh6ZTsH0LKe97gBpIOjJCUbJepJRsWypAaBaWxnIZ
AHaQ6Y+mloA2UmvO4JISmq1te8Wsre1JWOk1su+v+GYoemdx6z6xBjWI0Lgl6XAu
kCaZLIDNBo9gDteqo8ZnrcpRiFoPpp5yBgLxHJfv0Eq9Fmjxnx0QHnpu05+WK/Zn
SF8RD05mAiDSs5JfNCzEKWhbPuRR+HHXey9p5Je07TvGek3S6d9XGqshAKwV6S5D
v9cYv8J9vz4b9aZLrM8myqeg70mU6w0PIDm+ErCZoC29cQ/ovL6LwTsWPWbDqyNh
4OcvcefWuoyQEBn3ConD+rmK68kztCd7tF61QR/Ms23LiA6WDohJJHW5im+x3428
rLXu2HYN9YJzM11wm9qS8S6er7u7yzSxEtFXDZsf7+9YDblO+Op44BP+PUFT6K/s
YteZjWXSZ6sxfdv9J6JueZuIOL55C5L/cot+p8HkAkusCI892IZPP0pu5CGZ1GO2
k2l+B9I9J7FKeGkvvnYoyyOCsNmZfRCz6QOk8EJ4dxjkKBDN5f6Fol/uKnid9six
5yy3yTzY6IUt3uc36GyxvGC6B96YeA+CgqmXzZvChPxZ09qdiqDzBE5JnHolxWza
PXURZ2QpDmkqIxBRloa+v3yCHTAQYF56Bzr7AMkJ9GCpqEvM8d1JQg1YNQrV/qC3
13rqAWmpv7ouINeTvFlLJOvYNu42nJe7HkRFOsFWvEBX0NKl3tVA59TOfL+s9N2R
AlLvAYDJu0s+w9lUcAKdGknAPTqPlV2Fz/gH1M1oIlbTmty7gQfBUwmqtrx51Tyg
TIsKLLbg7s2IyZ/FGB3WCFzZAry0n44msBE5tM+F2zLJRh5VPdVl94e30SKon7OG
z8I21ReiqTGh9fIGehD+2W19t6Si4UKJC5usmY8ob5yH3X589ipcvagY4pM46dI9
gbpeEqHzPdHDjEVZqcZSunqmyr6GqDD1CCeV9kcGLaJqUNloWKZ3Ts6OfSVF99su
8k8rmXTyRejcG5JXGlzNmG0rGPs1tLeSFvHfSaETuF7zyVtDUfjdhRhCu+mpiKJ9
ATCKn4y0GLFiUDebbsU2/7XBfFk4T/YogBRr0vUFXaganw1LJE6hb5sYAYR36M7w
zE6LiOhnczp2jKezGkfYMqT9ZdRtjzz/W/f8rD58XrPm3jUUhOeUOofXCQ31I4b+
tAdFExYsQLAIfWt5PVR7DWpwdwrOn+jdO0wzineCf/v9y3OVqCAr951m+SqD7QRK
Y+QqS8S/mj7HVkQZ7qYqcLF4miemk+if8lxQ69XIi2kKFjWbdmjXcTKsZe03Y9Kf
PBy8/v3JCEF5eygvEfxivrhfuP1IQHnHe6BoKcdF51C0sY6WbmkhefsexNepdT/B
L2XznLQDcfTt8scV/CBe9eX7oSluQ/ZAGSj3DAHBBa24RzjpzTwyw4zfnulqkdYf
BBl85F45M3pOYd7Z0u35ij6WMfmUwUwnmlh1/1e8FOe1OFdTM9MOQnrEu49hDMiM
K2q/2LMT6pC895Fdj+fEVSA+lWBo6JFFQzaeDl8QsYtT28zz1JvEaoDVObVEDLeR
gIgv/pfKPwLOeD1ZlmwnKY5xJqS2Cy1zcfayNzKzTR4D7mpOPnIfJ/AJqSze2371
8uXEWwJzsfDmZ4gln0RjOVTPj6WS3AVuee8vIigeA0Sk4ZgPV0slTexhj+QHqSDd
j0jaakqIzHdBxgKUs/+OZwUlTApDUn62TV+8dccrLqO65dCvZX6OnTKFJWXEbeqe
aCzdWXfTd6bJmrTt0wNgj5kJeKXW9n1UxL9Tu2i+nzc+e/RJqhxGRH5UamJlk/7p
7N2y6PiVC6/qRKa3DMmWChlQShfusDjMb3XptjJnQuDxwxPYXLSS5opJejTz5Al3
JYCRPda+CXpSYONQJRoPc2Xh9ufv7NyMaVAadGk0rEriymEHPk1bq01N/zomFzRS
JJdRs3p4H6ZSuObYdfkNQ9sw3WFhoETyZgkrZDSKERvlRZczOqJOIFWCYGggusEo
Qdmd1v9S/RmTMhoTvYKuthVInMKK4XOXMLHbCds0T7QDr9inIcAikfjJVko4w3Ak
A2K3SK+pDHvZwIvKHthsdOicQTseipzh+hIa+QTR8csnT2ZIeUUxuaWHlvWM6jHW
xqQIbzFO9PcTLIGkBBYcA5JcAi2pMramCAZJBKcestgMQJTVrOPoYD0nZ9Y1fhwX
7ld9MThXi3I1Lo/s/8F6IRi3iIifSCREh72bnPkGI5S5sJV6dM1qmaQ6PSDNT5wx
8STf+V5jn2Hx2qVWqWSaNKu4Tf7zynA1Ya/gglSm0Ka855BuREbfAc+R4Eqli1Nu
Czbi+Vb8ofj1/nflPppqzhKelBPRhq2nchlRNMfw9vgmM/OSJMnrIq9P5AuofJba
raPpwcplhqFm6DxQfKunQlzPy8Q/GtpdNh8UEHMFS4InccxOEAKjovGSM9RyNdTc
wUywlkoTC7mVYLzfkZkBrkInMtVMZnqxQV5LAaTQLnwrq2QMAlrOOMbInWPszSgz
k1T+d1DSI1HUuVVvq6eyw2+lmNunfPFBTGQqCgvovuwJu6akEfqmZDGN+hknwJHu
qJ9NW5CW3h/l7dlsa6jmp64Gqkn+hDDvDWgcTD/PQaaou9cVcIgAr9f4jiBBcUaA
HoPmYEgtYvkjixvJns0P+pW+Ns4Ae6+1mgv0AfxXONRK1DZATj72bBGM86TTDCtB
v+wh7hYqWMKhTl4+Wi6jnLt8rKB4lxU/JlI5WqJ1VMhplx3TtAeckj7+Uxm+7dWk
7epu8GObPYO61HturZ+A4SQ87m/TGplB7wM6JQgOTaMo7tsG8WlIbjE9KCyyy5P7
wYS/7u8mSEtAToWPhxLIRpli8NBRgf5iOEyNwEggAgMus3G2bG7jYIxVmbgD1VKb
kidCz2xJr4NT3/b7oeTCgXS1HrAxvYGvYPEKCmdnuocyOnqLUUAroGNbqw1JVuRY
tMN8m3CgxXkxsCt1siNruxbp78xBtb0d8L+GnyfulkvYkSD/FmtrRHhiI/weSpZ2
pK3QBbNCoeZB2116Zx6RJcu0QNHqeqFvDPwgsWgsu4xOYFk01JPDcJdT4sLLvg0+
v1wCCPneqqwm8uPEnQ1sJuX0GcVObtbeQuekCocP4XHHB1xZrxixYmGJDmiwXaNB
/ubO4cR3/KssUk8G5wZ9RnpCTvlXEooXb9P/+fAgCXeHOp0PzVrTQZN7Ccx+s33Y
tVsVcyRYGjWaxMHZuhJRON2WxEmvVToEXMP2OcPcrxFhRE4PKpWBkt9tO7t9qyoG
UqdlJkRCFurcDoSiLrPeRFfHM9h4cmvyi4xX3lkiaJpL2wKKnuEkw0oNjU5hSUBC
/z/yAmkFn1x95byo4KvXR+rp9+BV194xr1Wu94lvabr7kMHb3HmVg7uNfr2C2jYs
07hoPNgNzxSD1Xju2IuGWsT0EM0DYjEUwRPj01TJPS3LRd0goyng/Dr9waciM3tl
lIsAUbfpNTAFS2aWfhisZ5AnBjN4EVpOKXaGCnmoKgkcDrFr/jpt8KC+OduRJUuZ
VCXnw7EBEMSlpwuh2R7/QgdCvPzg7wzlllI+4QtRxmmq80x4xbUKxW9esyDGnGzs
Um/IBeqqhridpjTJnECRsrnfRAabSs9shSPGk0A4Xmqfgn6AkTejWv1YshKMyCS4
DmMvPlbSdm2tB7ZIa2BFoExIkBpUriHOYphvVLGFF1p7LpzNNhfJ0tO7xh7XzMbA
OYe3MBy7SH1yijv2b2Q4h1tmis4T1lOZWSVTFoY8T4WRyRBtAZTjeAsXS1ohyw3F
SxraIo7hzWprtRcA+4dj36+7Bynkp8LQU+/hDyAiLavF4L/NnAXTfI9+pbo/XLs8
3nWOfbLA9k/7VvN4kaoee8eAEFpmPq03rdPCw5TpmkKcWVN0bCVxgQuFHn/ObQAy
CkwCUwPHo6fAtOVpycKd2TGBZtCiPJUj57e71C94ByQkJW5NI7O9XZKIJwAIhuKs
1wasj9DddLecSBZDg1MlHE67mIGkLeyRfFiMknIAfVG5tXOcFQhRvVT7G4UGJA7P
vuqzISVnvD6a57MvnWL7MfSRoF2P3PfZWxNravYvvqFObyAWZT+6njSnKl6XuxHL
Fe1IhQxWu/Vcms9KxlJiwTZZEofdbraPMA5KqXURrGuqF9cBLC7JhTDgEGMSGbQ0
+M/jgiA3cAG91dCeWBAsqJsS1oEv7w8qLkxSgnoUSswqFpo4sOPT2Y71GKEGZpQY
vMFI5R2lLidM6B6o0bO/NQH6526uYfTEh5i9Ojc3u5Dnkyc8HB+HO7C5NY5nR2OZ
NjupbUl5mBpRT6so06uVGpwQqWzKUmDIwChSHXllstzYqUZL3prfQssfiGwGxN5a
UPoGgeM3WthueaJUbZmhPQHmk7tCCK7QNIRxIDgddwrcWOvJX6Rjn2khQAUIBHtj
ntXhVp3BT+JyLK7OhkGLI2gs8HBrdJnEk9VgwygfJlEjay6AlKLbb2u+7jA15Is8
Ci2d2zrNd9aVhh/psrOxeqhUc9Q99evNblpz7gZAqttxkqFZPD4Ee9J25f8u3t3R
MJEuEPpP14xURuHWDPAmpZ0YTT34xEtxOi8DlOGzMBfRvANpSeqkZnBGSUpqb5Pw
8PknK6H67TmFoZBzOuqIhEESHrBjMn77TAcuYtaNfzMcb9VECqq+vBanciyoIYqe
Q+mvL4Uw6er+KO2sIufM4fsElf9y/H4luxfoHSa2JaAzj3WMbY1aQt+7rAEJbHAz
xK9OEHbIhlkZA2C4W/hzRdlagOHciF8F1GVk1oOt6/CG9ZISoObITuvrSA9XoLGv
luHj5+0pWdbj4dUE/RX/NfpRfnINprWa0KoNVzOsTzEb6+HHBecUgTjvenYSzy/J
sczYvn6LiJgsjQI1byaY16wEPB/hL/4cjbxQHcSwpKkRA17hkU0aTmXPYpeIyhuz
qrJHh88jb2SkykaJb9XR3ddtOMLiukRstt+61JZnBcIeo86y96dCEho6xLUCJ1+5
c+ivt3nz2Ufe0hKhqj0J1X+GVL+mhBoJpv7u7hLblM454uVAy9f+yUYGlsbpcrH8
I+w2pGzUTk7fj/BM9my0ZEFo/vchCiqN0ZGNUU9nyC2Ktk1i8248rrOfoyblPPN6
iORG4ps0WdewGpBKjOzLDLsHIgtJhmxyW6y7HBnb93PIRN+9qrLTcNd1Llq+lC7q
hMuJ391/eUOwYLRexxMAjHySDCmD8PAavSrVvPSMrs44yH8rrWiqot4iBgL3/7Ws
Nppt9RKOjOgewSArCDObX413WGsP6Jb7lxefZHj1c7xfqGQ1MyghT1fVXQqDjfOT
XFNeas8++RI1YwpsWs/F6ehnl/Yq55pdcxSjFLcYGci9i/X0gghGZAfSNSVC2usg
sDg9ro8xvU0Jg6G0KOOFAAQ7qGe3V9C7FPwzQJ0RlBjSN6E9tlupTuliyK3od7u0
3fw30jnpajT3yUYj5CrbN0IjF2+vdLVNoTlEijOPYWpk1JRPJyPxlxgB8Rvf/HeZ
ChD5LWJVN0rswagSGKt00pW9SdGfbYG17/EUlht/FnXe6RIpsnTP2v6vKpaL92iJ
73niFPjdLtjXEILbSpEO/rx42kzUEuiklT9bYzcSNG30QeImVBwWt/8ft6be6nFz
R4qfkuYTxaeTXcH+NlnIfWl+0IC70Q18zeYaxFCiprNcBgMJzlCwvFPQqDyc14dY
SgDOhd98Swq3jD2AnhDPeuzXR4CJiQ13kJJAFxPpy2mpvuvFiiqbehETSt2rmWur
i/mlib3vPW3fsVaf6frSJyPigomiJgyupD9UPfIZZipPytHu/yrSG37AJYB5ZHkU
dXgze8pwPwButz5SJjIVEL2+f80LZhrBtb9/NAqjoDedM3tGwUZXuDLfRGeXhFFd
uS8yk1gkTDCQG0Zt8kxUUKETqS1zczqHmaQ4qUUYpdjWpWGhJUM3gT7jNfjvNyT4
cpMgH+Uv+dOTi5kJ6fnbq6eRkc1fJZTexk+9Incjk1EXS+5WSu+1vznI2G7GhW6J
DJK/SGauPgmWJWMJxvVPQq3gxg159HXzenSdrIA+XSy/bV9vzzPtopDWaUZM7zrq
kbgutvMklEoOwayRvJVM6BxFcig4qvW7fSK8sWC1GXRP81JuzPjLbaEzOY+JE4np
o8L6VXAebJLqyOGa7w3SoTHgA2Y8hqWzwSdYryE5a0ECdqC+2tWwhAqBrhpiQlBO
vKD4oOMYaJ6cxLyQpsu80SfE8xre70A1vAZvFm82XWKHYEpYgbtqrcToEgGnWYrU
pWxTQwuJcT/Y/EcUXOEzJXRFAMn4ciokhUaD8ZkLQnHRAsIv+pmP/fRgn2a7fK+D
/0Ch7iOtAWd4otMjpvjTsHG4dvXpGkXpPv9kmQGJp9WM9HeOHjaIHHLzZGcHDwu7
g0yLmspGfggLLD0BkE6JctxWs2RmNhYkr6uSwlHAcxGSkGoNfcNwNTuj5X+2M790
9bjZIVa/NWXFAiC/fgMqubj7gDBppXwz1eG9Tve+l23lDh1wsT5yEnYjchQJ9XsQ
APnfPZYuKP4eXtqLmoD14jvjhKIAmEubM4+SnafR74bktr6uM5H0rR4F+4CMr2mQ
U28mCVx2pz74CVzNWCzgRHNIS/bs/OkuAO7TxWbv7exK6YwsHuITeu7hw10+AkzT
qcE1lY4d+B8s1rv0Ruec6S7vB9gLOpbzKnpglL6yR2V+w1Ies0WzC9bNA6M6x3jr
cvcZCpNYEhllbHho9LkbzISD3l9zRrPjo4cidqU0dSUUS9vPCggj/zCYuHkxiWpO
Likt6e1D8K1nemNB+sAtRwPX4OSrz5Qe2/qcU1Jum4Y0w6lAT8XRhOAzMsOL+3/b
3EAi9yGFEdZ1fawc+p1sY/pRGTpoxwNhBGOuVdrgm1BgihU4HWmeSbG/1W5U1K2p
7HOO2yTOyZIq+IViC8+UixAlAlhc3QFBDVLRP4o9Izk7Ip7gjLRY6mrJPdMuwHUU
Lb/4W7nF1CG4iE1jS0ruv0pAu97yUfNwfAvF39ZIIwffxl0msuSb3Pl7DBQcHYUw
EuFFpdCblTwDogcqdEvVbhEAEEJ5arZuwK6kiAq75kzy/imzJojy/w3zSO9xlkYy
GqZLCHh6EGJAlpINNtNzRBdCltGOy8ewVcQamSTQEG+FeuimEmS0UrARUW4XHuTB
inC8xfXPHJZXQVar2cmipRR+6i0XyBSY79JQyJ/+RgYE775TP1DdI0sOP3BbkH1K
9IRiWsGBWe9leOVp/Isxgpakv8fuac9UKn4unLgB5MlRv5Ra/Vu+bCt7S5ZpYSp2
WSIeMcJeWsVXwrgJu5bS3tN0LtZkUL5VqfRY6LYOD/+zC7mPXRvzYJ8qvgpfyIhv
vcVORva7YR8jCOX1GLv4nUvmdbPWgY5GKhsfW3VcdO2cjfUbRe2EYJjMbuzJ71Og
87Ndu0+oui4jSx+v0EcNpJWToJAfw7hsgYjI1144Q7vOeX6n42j7cJXwaH7S3O41
a4xrqoVSGuIVg1xbslQhyEhkrNqQHt6WcT4yqtMDL2xA+KBoXAzkS4eeqDGGloRi
rXD3yYT/DjfDHKDy/gqlqp/7c/3xF8ey8JRtJ4kOwkO8vOEbPNufI2EdEGTZu7kP
t/xKlYmKdYByOo1aU3CYMacBaYDJzM8kEHMFpznoCtEC/8Ea6egKE2ry4W5KjIF3
RE2c/J8LPogWHTd3B9KLrY8UmlscFaWwWc9njzgwdTGJq6TabCJnttM0iO98RNn1
bO1xKLHmbcO8dyV1IDjiqkqOmZiOoThelsgYJAGQu2LvH9K4CVA7FXmcn2GW9P2i
iXtKHS88go1wXuAiMtucapRrFIVg0WQVc0xhw4T67yVTWrs0gOvZm6RHxSZtDhca
GFeUp+2UXS4S2r8QqsdLDxZhuLdVQ8EHUjeEPTQ++cQ3LH537eik1WURP6V57Prm
4Tam6x/6x1QejgOGHh27jgjLyGphccztcqmzBUA88bRUa+WZxCdDH0k2vS8FXpnD
krjo/tko2YzG1c0bDGkSoP+wEtI+uLYG2m2X0KM0DOOiU91xIQpadp2HZWNE5Guw
4gEbFY+wRawxAqYH/s1BXfts5ZBhtHgn2LAhUPouRwnYtIc9eBcwotu5V1MmT9dF
ZyAVzy3gSGYaTCKIowsZTdxRo43fESqATavRXVtGbrUh2VmW1lGOl6jAqWIESocr
VpcUQIhun9RyD4y2j9Pxluac0LF+GTY6iZfLqodwUVaGNj13DIr4fIo2A2tgBKmT
Ajz8pWmjx8CDEvawqnfW560bZ0+bfp2fK8HuByvN4i5NBA2MSQKERGqOH6peGmq9
fPP9811DCJN31+9W98+Wlu9FUyQRs1CtPiZZjNwUFNnK3P6wdtTPcfPPcnsKo71q
juEzO3CptpUAahPrNUrWpXUcTjA33mnncQHTbjSKKsCV95KyIPggeDcHTDoZ3ewP
ieKXEqu/Dd9a+x5RY1i2K9CCMmluTl/I7SagZfhxzQVeCoTsox+tSVCCuKxCuBUN
ue/marDKxmZAZbEM+XwkEiv2npDB3nhUi3BknYn0SwYSfAYu3Ln2GeRd65KwBFd3
LFBVzlyt3yzZhtjo2VbSh2XiwqWJWgEBhD68ykzc+/Xq7gUG2bnt4H5j9QuwRuy4
eNDzNebyZhU3bQuAG7e7F4V4RJoOvX5qe4coTtD30IUPilDly12AeDe+DkQX23VS
Cre5ZUPwrQRws0pT/+Hj/kK0y6l7F7aqfULNAVgMVoMGs/rcohT24bWpBuLWcouC
/hGsANkGNt9vcvpYppel6rDKLEohRhAYvmHT6ulgqtX80dwEA8SkTS2nxAFQHPat
YbnCzwJzl9UM2nYsNMuIXjLZZVjNCP+T30T82MubY67e4yqwLQ15xYnI/ZCBNwnH
lnQo2l8Unr6bWqT30Ofkyyrc/61oWmf1QwQWxSO3r50HkjAvXvZv9qaJTcqHGQMH
qLZz32YyFCWPJ1+AxGpvMtzALTLhsFd4d2n6iiydg77k1TyO8btUH3UtyDXyeBQf
r4EAiK/AjBuhPjNr7EsRHs0/TGcbET3d9AFHyGvJo+GByVRd6Ss+WgQg0hsH33Mg
ZVTluH3XuNccuGo3nf7AFp3CDEpfdu7vsRb9MKheCjbwdYYeMT8VUfO6dyMaJI0T
1fqEZR2v80epgdmgPUUC1ReWLFh0t5h7552nhCcB25dOrjLnpYx4jV7dID+j3uAf
Q1MrVTpKyahJwhuj+dZ4U/e7L6SbwiWaFvZhBjZ7iz7FU+gcGUEnBWLjzZS8A8MB
fN7B4EvDkwhAjqi5MovXdQpk03JGl5x01b7zWOgLz9+b115TWvcBXzzchS0iAstN
tVzIayOiElZ4vtlp+BtByxiGXiVsQ24gKkdaYPvQF8mVE6eus8KAQOHlikdusDTV
y0WHzVuLHs4+RXlR0szheEK+UtW4w7Osl0taud5bsv10NG7l88ikdufXRZ0U26rc
fM2sRrFliJ098S3cnTEK/zgaOdls9k4Sv/o0nnbYW0caQcFu/zlkFfDOT3wUxbMu
odepUxckYkcuoMeCVpz8WdxHK7Kh0+n44DGJbg2UClGwYRSUTz/1Puckmn7jxY0u
thioJwKHQiZJzP5+YhPubzCbb+bbYAFGOfTlVr5RNr+Q4a/bwOxirzr2pgQiUk6P
bc9i2OvP5pydMxq4/PyBJW5Y+sWVPo6nod3yTPprDocoWlztJMVwCMgZuJWpkBv6
RtkrfX9oLt01m6FOqevkYD9VbzoXVz3O75XZ+ENQlx6PUk6PiX28rF77+pYlSDB7
nbk7IBHyBAl4GV1cM8zXl43GpxhpQGcEjAl9C05br196oBpUJECD699HgkqAFPGX
ZwtoXrclw/P64swdKmJ82WQIIcDBiKrBKu0PcYOtJ3FlNnjPBy096ZwIbrUADyb4
T8WPQfU9Rlch/xazp94OmDjq472Bl+g0tI7vPmZISGoJNKpuMpdgJCTn+Z+XoYGD
prWrhIzLZhpWpqnSXW3kStLm2b63BK2pCFLAJQIEElh2oxrWAih+2CPL4KS2Zh5R
CtxrHH83oGsEWOu39j3ZkK5gz9rc06FaK4JfKREqH4T0+pJWU77mZUcerRuIlxGv
pwkSD3PNizJ8WQAX4XgKQVU7pEvHowWEIN3l5zLanLpOIVYYJuswcPq9433PMEdj
w6JZs8ily61JKlEDJcfVRv9IlMIWHn9dY8e4GyAAPag2HODxnUSxisaaVE2pvrec
rL68q9GIVycWQ46mH0zPBRB5bCDU7iAnXrWlSNwGqvjOLJxz/tRLhKvtsFZ2OHwa
SO1w1dXX/cvamFmxDm1nxzlfkQvKxTSPLFvm+HRMhvw9sJxNXkclj9JoFS3Gbb0f
SXI6qkqBWjci+1PlgAZmuSIumush+6MkPApeOgA8fSjwprNc+1Tlrv5UlMoMokV9
5UeaKyCb4x3YaPFJe5mOPsc7aEr/UhXJ2W6uYWQAPI7riH9tSs+P65LxaWgqEnHg
+iQ1mp5tpWJIlPkjY08VrhJ1zifW+y82MukbVlC7Elnl7Tm1e6l5wOY7Wf2tOKTv
J2zJioxmi4efFi2VFQf435c2xdgY7pxWf7eI2w2/aSw0QUcRu2H6QtX/CwDsanuj
b6jfA7utC5nWkxtGMsKmYdXCXhCzXdaMP8cm3dS2aKovj1skcp0umd8/vmuxO7bD
3rkDn/sdBGP0fFyGFrAeTJtv4jnJjkiQiXcWQdqZhfz2cYFMHpUHNpIn8ffauBvk
Z6lS+rmEjvePW2jNlppQu4tEYB9pjGKXpwGc8MyuvVQGiW93G8/DXQquCihyQEj/
EpQ6L84D1qgkarn3933dKxZ+r8oU+S3lt6gM3azIV3BV3K1PVD1rV1y5BJptuAp1
CiItde7kA9GUcfMZ5zhx5eKHWWSjGYFWB3VT0vKuyQWP4YR0wd7VX+UHmp5eW1Uw
7wSetct+OyOO3/tNkU5IZrSWXx06OMf92fjrxznQjGYjK7UyXu4/DSbEutUzJiWF
rmkdAyaYOESbyMcanwI753rrGngl6OMttTEHmrEwTh3tMqcjMqDaD8VcoXDhTpcU
WzW15ffLZrhUFQCud82U4ZqCKDvPpju7SOxb3fsNL3NktxZe7AI9XQL5Rb5yAs+k
6ySNMEIAbKqWWxA8q1GhnowiWxOqSknI7IZ91Iv9ARVAw/y0Xe6mRTs6RGykptpd
jeH0BNJDHET4tDZSFMU1NFbBh0P5sUNx0EDqF5Bq3Hjs+Iq+Q7JLYAtQuBv88FZl
j8hwN1brKKa8PUEtDtXLnKzJ7bW2OjLf9sx1Wn82E146SEB5WsvXHVc2VtIwIw+T
0mvId4cuAkS+QrVyRqXOXB7/M/sGZad0MPop2FeBSS75+66G7iYxbYZHACMV40Xc
owPTcfAYi5nyCrHSICjpK2mDyXFP9X1WoyhE838r/DHCdtSNN36w8Q2YS/7iM/pZ
vjdGsIba/lekFD/yRiDkf13zgAMKoavs49NP1cQFW2Y4F8cMjQGGvTbDhu2PC3YN
9RXUXXfPslgirIot9dwFj/J+ZumCaeYQ2JresRrxwLi83LvGDp2qzMBniFFnYDVJ
645SlTnrQ1gdfFrQZTM6HDgOS2025nFTJ58GS7Lwoji1NVgPIaea4Yf0P+j4jMxc
e2KnfoPpvNRfOpMOcj3PRojgkLDib0OGgW6rKwdtzUQj59H74t1DSJwUpX8LbmK3
OWE6fnPGXC3GKYpapFkLxWmi0W1BwC6JdasLQSECX1afYDuPiXcpNmoYJYdwcy52
Ow5f5vs2Juu3Ip1ISppgfo/9FKjJxXpw/RJuHgwn6Iw0AGtifafe+w1MI9xlVdYE
k06mnL2J5kSLWeKhe3QsQRW+p0owW4pPbRU2+2yByPb6ViB2+pC6Q2ItjO7QxnpZ
EqUK2tl1c61FKPZmDahwvblMpPJLIfVOQ3+IgrE2YsJePgrWHr+ygIDs6JQM/yW3
YiZRCOtJnIpDdbE0TFAR0U8PQc9j0ch2xUgKgoI12OR7sWk7Y0pDj25jofaKhbWr
OCC6EwTJlRcveIgmbAO27eQ17DcU7tHzePvoE25JwRtu7MJIzoTSES6eFg+DE04r
uMdT2StceBG8bJTR8PbpTXAWbUbOCA8MxRqe6aiXYOtEYoblQIi8xPiL9kjOSPNz
QmhC0wSquVQEt+UYXVX4IFfl83ZYuNFPYT8gPmgDEmFQmol46NkDGvy8Ce6+72E3
Ja7MqhvgKIJL6HiXI9ZnjdqnwHDVxZURFgt8VJKIgnrW7uGlAMX428EdOyloV4Jx
904D/yTR2TtMb53+wZnwlcwGgriNmBRGDaYJLY8LJw03tNa9tBYXdhZC1vuJrOuY
+ao8c1de1cQwVuS9d1aScWOXEGGVH28bKd4S0s4lL/35HEAcoYlIpWIGv8pkcJ8O
5Z4RQe3uWyzS1Rn+IWfNB+FtNia/4wqLC27vYOKqqy8Pld2dfw5h/lrUb8XdUDHK
fr0hzvQLYodRXlnnFXrRYitJYSm9XKYNsIakSYQOTiIKRFOJn3ghez0Gi9Z775V+
E27KGXPY9blyx7CKwHW2eNudaheOPGqUT/aMXTpVYM6K7CROCPms2QfYgOluUORy
YeijGn84yswd/TP/scjODu1cGuN4t3mCKRXtaramhlJU0JfPAb2uB6IMtDSAq2QU
SbbB6NawUqUSr8VHydth8/JX0vZ3KO88M4UQqii8slnwi4a03K14P5sNhr9WiTvI
fVEOJhE2DYCd/lrY5LA18WuD8ceV3Wigfzo/kdPWsxwtv0urzfLs6Y/YEUrOuAGX
zC/WvhufEI5el4W4ZlOP9/9l/068ceUx7vGh7y4sjIOyZtfmyL5ZGRS0HXCm81aG
ClXplnptVKTt6PvK6MIQpCSK3sk1LxPf1Vujcf4i3Xhme5/888WJ6+A1lbB5EKHA
jaKwjhzP9k/1uDEA7lLZ3gDkxxuTuK9WX35dJ6+hHYfIIkYbrGLBfg81U7qsS1sL
JJaCrVqTXK3U9VaygByPcZizYGhX/1v19yTAn4dGSpKMIi31SvXB1bw7hJe+jveM
gp3dn4+nwjWYhiYF1ePImzaRk8ZskwV8HfVtd49VcDmwj2Hbbb3v9Nil23QD7NaO
za3IQ/9XAvULpLlbAQQ14ZrCfRZxIvV3c2zOu0YJLv+w7KRtF/pTLrcGzekwIxRh
fRetw+5BEUFnpPG/dQw1GSTAaZ6s25FugYbTTDfJN7Yg9jm+CFTJvE0fY2lp0k7R
sGCZdQjDF2QmPgPhg8V24QPHHV5f3/vmFG9KCVo5+jd5+DAD+OCC0Gj4m0SL1TpA
cHaxlDXXKk19gGe7aQIhaUZqAXdeTWeYcD9E5tzRzzWIRmPu2ZZkDb1xRbUnbFuz
a1HmYyLCtssQLVDvOC/MMNsgztd9jWHEUaKri7XnaS23X532mYRi86vjtL1UqeJD
FQ0qd0ieScb2S15jMvrhWSbxTzUKs89vB16YmK7gs5XKSgesN+YAda56PoobMPMF
cddzFw6L8oX1EnXfvl4eeDqqOvMZSDWkmD0kYY+OCy83OKllfray1Sz4L6k9of5d
PQ3YAOIgX2CFr4UdE96rJMvxPhWbrIOprhrNWr9DeB3ssNCvTjHQrW20aMo6RN39
+eDHqT+FSFTx/5OBfxxDGnuGqymjgRds6JGinMCqw8Bui/Tf4qQYDUtQkV30FllS
IyDLkWlL6oPZJpy+4F3n+OFfrlj7pGBq7cORx36abhO/nkFAVBTedJ+/z2PClqOk
RjaU287UQhnkPG88VoMt/3818x1wVMXrK7RtlasnbbyxluVoQSMbIQMxLLGJliHe
uB5oRsU1Z4OwtUjxrWriZl4jJnV4lxVOpJlqYaWt4Ipq/HsIU3fz2+ff3OpNMj90
ZXDDDryyVuXu0fBTEgrNPGNxTGVzuvGbWIDdFwykBhjNYp0IS7ce0se864BME+ns
a40M1ij+KdmPOWpbRdL9vOEl2uttOCyP/B03Xfb+A/JVj3NiO/WncMzHcLPy4Vvt
bsQ1nW38FBz1IOcXvRM+lJLkSskNSO0TM5qiy7RzuRuyaXtVqcFp0uGP8a1ppzQc
fwtlfKpUBZWwdHQX4xc4caxXQsSuI+g1+reiCzv6L/dCB3/WebTGy9jshmyf6tFF
h1w31OSEanh1JGww1bkCjIs72SzWyAgtyUavYNnbfLX8lOuDBX8dz2DEdLWA4aOc
uPWt3Hoi4vfsBKm5nzG8G5XcEjDcGTiZKm0Dx2lYAItPw4h3HivvLhSxeb1cRbtl
FudCbhhQAfccGRKO6LbG/Vf4+wrWJSa/rIh6wzk4mYmNOygpxAJh3INsKrFTneRU
SqaucmSyc207qQiBjJcVKYXBUUtdgd1lZPYC3YJy1XNkQDIF/Gyp/B3zt39S5i0j
2hRgbKrm713OMFoW512N7Ktdxwo9HtIqoVhSM9GOgKBAIxNydqTvEU0QjBekkBOW
1pTuu1Rkpmg3zBlcgn+K1pREecObF0EU2zCoTrhRPR/byAihjt8RVcGSeM50EVDu
aV2xr1gFFdXp/4JpoMR2YSEBOWEq+47QOWKlcPV+zliCExk8W3S/4xtDIkX0NkVm
pER21p3DAC90IXcYfAqCrBD7/hLmBNZ073guQNyO39xR8gaMiXVCcUH7/HNKt/Fd
L8OQwwXMTzxp41WvYkj32ZgCQGGJvi5mtoKBeDGldXSMrUPDHvt79fByQvrDHBOV
d5Jx1dpoWAU3xKXqTFOX2nIP+D7dkPAkwkB+7jd19KlPQbBQb58zkw8DkM5nbu9h
T/kgUGnc9hqgFg8KUomrM3ArOQTqp1A+3iiLpYTIMmEGueP4Ti9dwAlv2AmDUb5S
WvYnRmOdpthO9+2MDC9um+U0CbTvjnhstRBhfa3u4eVcrhnj9MAW6k8adOdmOmxj
8UAsWeHnj4S27V59SonVbKYNgAnGnAXk0ygnp7L5V6FgrzDIagxTYzWCK2WQfhj7
dOKgAadjrBE/FbAolt1eHE0E6Opt+P6XhCzrV0CkcZ5Z8BBTIxTdpGe2OTFbQlA+
2FnAn6R5o9Ocgm8vdn9LOGigEo7VTK1mTOj/gn4XqsnLdHj8dbr5D2oiDAV3xbbQ
WluwTmCD+nMY2q+kI4bxiWdqoQSNYFMi/czmAktXmb1KfGHZlUyhN8H0+5gy4k6x
bunNao6+Fk4i9TXDuCaJ1krCpvWT/fCASsl7x90uG+YUm90ZGlJf+8YFmMnouteM
0clqI4Dk2ApW7C3nqa4g2OPCE5kpIbMcMF2MA7Q3TwZu6GCGBV9jhrQaSq4zxP/R
OQ3fkHcUxiZb4af/Rl4niD+k9gLNIhl+T9Vh99dllciDiA9D1BQqMHmrIQpvqPNQ
A1o014vVh0HSvaSTNbglPs/2EHjXYhbffViSFPO1XMDKNURGYZFd2rDD+Wt4Wsi4
OZhUMXGAEz2Bsy2mtOMrEag8ElQ27an3HSYSQIUG1y5zcwTXLM0iyAq17aGUt8Q+
TqSLn0gvyhai+FQuwkNm7cvScQI14m7MC9bEYbNQnQjWre5DT6+V0vHppl8haQf0
5djMWyLY8XXRNtBisCZY4BMA+5CNK53kzXGGMjPsHi74aQzY55uoA07fzSr0Br1f
tlwq9m7aZke7ht3QRM4ySdSu1cUrqmnJqgq4l4JhJc1hDVz0GXsoEauz5bXABqYX
BKyb8eL2gi1LX14sth79WSaaqh2cBUoaC2gqB2Q2Tgqd9asPcgmJxtmr9kuThffR
IS4Wt80r1p3v6StSMt3SzRZRiykIv1wojpp+vwqEhNluj9ZQ0naUqjai0o7nqrSp
FI9kyXujaIJY9ORVQAO8W+LvFalT5kt+ObXLhdeVV9zCeBFmqgZ+qtNI6PnfE+ie
prys9tPP+BkfronRdP0O39n34h+NGH24UAWWBmHMQXcO19KpvnmKjXVAYAJ18UCJ
kKP/z+74QTlHelLRaa5grLvkqLAWK4apg7Snl6OKM3Jk7VIA7WT9venpzxxETK5q
leK6/HNBXA5NJ22FUVARga3Qj+3lcpz+H/LIZpJBtMqOnkrH0l+kPCNXSWUsQFsE
rtRxydvPvS1tiOXWbmG24keN/orhrw2Mhg9V/1m0Z9n5GSSZGIi9TkB+QPn8n9AV
buQO+jkUssrn73+/dlcwgQuqZupb5nvAZ2+52q8FEGFpN63N/WqCXsR62SPEfyTv
ncHU8fHErA5MhHw9EbDUyA1ej5drvAgJ+9aqhSeoe/DcYEfdAkPde1ob2wm/ViRR
GorNZVu8vypN8OT0lWm1gRLKqSroW9WIFNucpogWh+d0d8X2ajN6vU8CIbYUb9d1
WOybY87ZS4bX4z0/dU7pmc6Pxrmy/3e1ORB2Pv8Kcr7WXE2LZAxKifOuj2XbbJqu
5bGihdZD6++1+a0vJdEi5c7VXLmRDnchJEZHWfMIvvsNfkmoav+ar2j7F2R2Gklk
jSTpiDaCKXfPJMPrMk66NZYUEVzB8DguDscNQJMCrMWXUO3A5vg+TH8irpFpTa4h
P8pQ+xjCyLPavtNeWgVawgg+YRttF/YRxbN4517Jls7j2IfN0jUXjngKXaZhGKH+
23ty7G6hV0/xwuAM9mYKlxd0+SYW8ZxboTqdKEKfG0Z58nb5JM8mxh8uVwXABBzH
xJYfdAkncZzTF1VkMNUFQjBoddu1ryhm2sOD42TIh2LrXsuv+23zfPlLDoVK60Sj
lr5SdNDLL31ZbWbfiYJ+P1Z6ROduShizbeC5R9I7LWeFyocBXfz/Hud7oX+O2nvV
h+ZbfIAuPOodYaABaA5a71pueW3Vc+k9GCGLNCPh37bKWf7qpeVuHkcUds2hYlC8
g5BZ5KVM0oZeTQOFScbTtDl6GtVnA78JJG1wRE+PRaxDbLeTDp9xYnQD1eKGwCCR
Fk/mSb3C2+XTF+q4X20WXkd3TQVR53b89ziAOdOHbX8fPffIbPwAheTaCCTYj9Q0
UJDgnDR03E+ngrlo0gJJB08IveYrAwRL1WqXGtkOpyJtYehcTubrvoc34uOgi34D
yl3u2hXD+7zW72xs6ydkEiL2jMuJy5cFTpkWJcQIsbFfYp1fU9KJvBHXL9BzUnG0
E0m7edmBAW8qweU7t7WpJCJDA5q0l+LtLB4VeV53qUws80QKb3YgDuMhfrf1NTuc
74tIeWyZ0BevzRk/P4AU5vjMQTM335dzLp5CfdqSiW3urcq010OV0mXBnVFXAxR2
z2g+ZPhcJsfKezuTIY2Mjkci7PdPaKvC3XEYWkxh5Y1nqCinnuRecElTQ6ShiYON
9uvHFJqtCnQJPqrSOH2yynVHUxpt+EtiUyKEh7hCCdMd4y5tTCvrZwUBzJivt3px
nriTj8a/dKRWOmUqZuCjuvjIYPYmzfCCGe5WO1TJYJh36bs4jDONIRGUJq+wo5/x
CN1SS/Yf9eUUkoTvI0WtlKakx7T4eS2B2CCDpRGTQ68ZyDzzawotg41vqAip1u0p
0MSxT4wR9N+OhvuhD6Qu7wnFVGXe5AcgiJnaHiSQ9Z1znTBuQPK4Cx6SHJXraA18
LYjOCmmh60ULyFsgHHE1KiKUXcCi4D1zeUDD5cLl7UtjbD2nQoWTPXAguFZi4us0
u695PA4LonIQBks5j5tWOqfNdO3nLnDfcQei1QAckYpYkrOGDJdN1MNOYaTVO+XE
xdgRu+JNQI7K2zWfr1kNruH0XN3ZPhPvu1M2zS19VOzNco4BulgPB5pPVSHf7W0S
ZDavnIrr68veomfIYQU3yElDw1Z1Op6wDq7cVOkX9Jen2hGNtWM3Ss2QnqajE7G6
AluCt1aSKFwiS/qK5BB6I3HR/UVbjGSGJ5mM38M4tTBWo/d2mzPje/VkEnfbZDrE
ohWyHZDyxY0lq/I1sTLa2Y8w+hUzwEOFOlYgytHHAjY7mQKQXibwiDDl86EUAwW/
Hh3c8fOWQ3GuSgbdBtxyN3CW6x4dOVSU039JQXwcd8PCwq7slqV1O70+babXIbYb
bJhzIfjxD5UXSidrT6hCtATlRSb+f0Edh4E1aqwa1XaRuRDIp6sSEvrMkYOeBBBQ
f+TQoBjOnlQvIadkfQ1zf51lRifF6GqvmVOxeREmQW0vxZMmsgq0ckLP/xx1LKvS
JNmJtLpQN0NDpASaBAJ9GXGOpGwU+w8sm0AecGkbjN5lQZRGWQSLijMJLHoMCutq
Ov5sr20IOl2SNmupfN4NpOEueHzlJyGF37BxI7G3KGhTvXtKyW7MkOsGEx87C0t6
apwgAKZ73VLZBEYFGchhhwKtuODsGyLh/BfZwYbvuStimGqTpcHHhDKmhFMY/7Vn
kazn5Oexgh+LOTV6Uy5B9c8LQiL3TMxT+/0oOPjgwLk5Z9CJxxzM8crkrs1QSDU8
zpxH1m6khB3uyTGlWjD2/5CfG6bqDfkpsJUYwoZE183TvQtYigps7h9KysCfLENF
KMPIAuZr5/WpEtYcNBB7f7sMpbbNCH9tQeoFMYYY/VOvtdGrapldV2Lm9yxmBg5D
RQ4BzYQU3jxX4MYwebSDPtp4I3MJiXlZNuVs28x6u+KTaZpOK+JvSd616tILsMVM
9oHCk+ciaU5c4coj2wFf1X1gHEGQk+CywqtlcaNQxfoQSZ6zTF82GzTaI1JwJztY
RYrFabgL7ip925i3UnJ7ekLX8PbbpQVrX+Emw8PGrMccTQhmyCsanxlVaBRSaoPf
Pe3QI8nH8UOAr9ObYQ1+cU8ZKoTqPa+ohF2xQV6/+iHzvk2ScgxE+brO+9GQADBB
lniKDKx9ue1ySoi21GWYbZRt7IiSPClpXZcG0+IgNTzMmHJst2UXtGDnGu+6XbqN
ifrM8pkgR2F8hq3U8q8+nCautpuLUluaB1OntQXBvwqx5coEzAOUyF78qK+QWoCn
DfpIKS5qSqXR18HzBIUvOOiwrPJSRxdCIkFvAJ7AWYkNQrgWB5R0XIsMPDyqf6f8
2/mEQMeXqa1YTB8n5xnVRVLiU465i0FOUG5JOprHJBtyISNXBhEfijAW2Ph87QAx
zbQ+MynYF5/zj7lQtHRWP5bTW4rkwxNqyMJd/d71VffFkdCwlkhvXUxw6IKLu0SR
driGA6rqAgu7mzUOYzV/PjgjubqQJ2G/wcusmlHgESz21M3vNpDfUcUthAqhKx1n
946OZgmWV3kOYbGtdbDjl+OJ+OaaWozUqhyiA5MbubZUGN1O+ivvCNyokr6DHQv6
n/iNgoRXRxCbNGFGOiCEQ4A7WyUD+oOZv2R9gmQgUy8ds8T/s3zRR3zvf8NLNyQv
gBM5hsD/C46Q1C+V52icSroQb0f9tD4ouaKwMGrOYQ/+pPzBXVWQEQiRaz1O2GZK
LCt1DRTU5xRZxvbA4k0silatBJVV0H3Gpq8z6IH4JUdsJbWlYX2Kisj7ARNWjmoR
o84yIXB1vcc8V389OXREIeWa/lozInYhHDAphZED2++vXz8PC7wD7yVOrkusKZN0
SOhA3XNr2E2g1zpmgzz5sVDkIKiNVVK1nshTfY4j//4nm76gQfnyibBN17i0Gowx
QTMR9Q908aVGyh2lJuGxifJuK3sgkKYdt8Oyim3+OwUxyPeJmvhz5e3ADdvr6iF9
Kni9NPQEZUx8xcnyXkV9jHtJgd4Lwvcwjq6/IQONyW1cswULy/9VgEVuThZuMEQK
nRgm9hYJTIItnxvAbcpWrEoaWltHLnc3t2I9VAcERrPTil79l43gx2nBRjzEwlVB
2eZ6xEOvmh3WvNnXS6dzT8AeKcpBjQXP8GzOm59OxswFrgdTd2uKCgaoqCDEa8gU
XVsDgfWTD6q2o/2BunwHDb+kGC3JADk396bYGO8edmOhG2G7U6sDFvzz4NBk4GQf
1iOfxOQJCpwn7tFaH4Sf3o6KSwUhgo3/rLo3QXYqVwhWP+6X94nIDK4DUuezD7Dl
JldtwNAsLGXs7jrDk7KpnjXCS7rmBlHaurXicZXcQuY09Jt/fDmG5G4lJzGbBM4O
6wPgfeRZKikBBXcrdgMauN/dH2f+z4H+K5nQrv7Kw3ELPLIhYDskq5K7fZGNsPQ1
P3Dw0pmjp4v4KqvLyhSK8QThA/llL7cdn5x5wJKKQsnpxTbGp5YkTQne0Gsgd0md
dauIzMKFnN3g8isWVqzrvqE2THaN9aSLCl2WKow+zsAaLz8i6SzC3LrtbCQFFsmV
nUAZPbC7lDZXncRpUTj5ypJThlltN5QSmcRxi1DFOOI8EkZO3c81K8Go06tKrynU
JiUrtlCojtMqGFBOD323I1BraH0tzfFgC83nnebc5jTjcTej9Au/7Nh5RWmRkqEl
YvajbMdMnCJNcvVOOyZLOCaD3JmIp5DqUcjHy8Q90IdGpGdATy+b4rnGA1JGdC8N
CFRGgXjjEXp56whO9+u23d/v0EWPS9h1sUWTvkb+MO7MOGTZcSuqkbXPw6QBzZiR
V0bHurH5P66I2e+rXfulbFJhJ5+lsnrRjq7ZmWgK0s+9+TDafOV4qDWd4qmBMR0F
wzmd8c03ZlRosTUbTYTdpz+ZNRPRg0T8KnYmOYS5COhPynNm7hmL4i4XEdDfh8+T
CC+E2JPIdZqFLVas7VmsUhxkixxE7VmM5k3IUmJRPCCX+qgDBLklVLHTH9JGKeh7
wwj1AZ0K3tfCp8xZoULdwOpO8aFr9RSgTOh/QQH3Q06SbmmRb4bwWVIuV3UXzdLL
uuKY7xiZCfk0OXST1m7P5o3Z8Eh63yyMws3nSzkexYcrU2l97vjnrcqazprlMXrT
NgD/adNI0rP3aRpvJp11h/eMiO0ViH6GgKupknvG940AY6aeaeDeDKHz2W8DqVX+
ZBsKfqrqjEX7E1sCLtPRrOHqy0RpU2i1l6ajQlnDHWPULJn0ExdUxNmdAM4ot92P
eufFOMNsSx9y9j5KoUsr+nw1jNVcaC6jzV4Ky1/qtsPpWxDVte8DQzaxrFUWQYyR
yNYEfyy71zd6oAKSqtUj7KZL9XeB2Ggvh8yWTqQMnbNqhqHIdPWt4YI3aGUsg4rs
ZOHiCTNcsdZS36II946sNqSa0FjDDYgSDQOii03r1iXmHqq7SZHQJHFMb+51dCHF
ss8Dy7jZcb4KDFvty+Jor3Kmdo0cSuME22ZuO/Vk2qSY7v5Onw4wRLs8sKjYJ3cQ
0L91k218F+aVAMt9zh82efPuj8V0sRa0JAb9VSV6Ze79nJdGhGNnVCqk9tNrRMVI
LJVcrTkni8JFVtuBIFodVnV+cyZ6YBJoZMu4bHATbIOIFvznDelKRJYFrizPEPvV
eYTt3C5OxIQJw4GKMpp6FTC33P9ffIbp+kRIIw+yIj/PYox/gRZKM5oVXQzWpq3X
AGogPu80OZvXUu57mVdNx5Gh+wPwXzp34MbX4I6cFMKNcReghCvqyQSe/Fjk+9sg
e9RwIw9yaExzCy/IpqXyGoXbxrkf2MjC/3zyRrT23qoxy7rDL2jGtFLyvrAYZ3jc
W1HQu/FC7VZMQQIbW5M74Dy9uBwO7lVahJ1GXUp2+DfEeT3ohYogPge1lClbbm45
5zB2ZnLZpbraapSZHKjtToOAr3E9a4Z7vWPZwB39idw0dQ7MmvgJOx17p3lWiysm
uyGAhWXVQQKVUM8kkXog6zt4oKDUghVNZP/8sgSte+84FW5+qHUr+3UfaXpZWIQA
VKvat2yjXVCVWMPxbJwgi0uA3l+zRlfVmu8kVap4cBRGrTFL25jaFL2MlFOTMLt5
ID8ZFjTQ5kvLYdIqjludJW2C7ZtINQGyQWcCNxsl2m8ZwlFbhHJCf7CfbNK9APim
ny3fPQZAJLhWTniCvtYTe+8cBgB40o+Y5GoW3tkXhh4glQAeEzf1uGMg/KfzGlXb
TopxqO2FRgZJInVVYSLE4f6Szs9f7WYGR4/WXvoWlaYl+T2q6aR5rB+7yo5Qh8q3
djXVebYELFn1fGGNTMHjPD0AoTpJq1+xzAhIqo7cDJPKYmE9+POowyKbwd1OGY++
GF+T8dDM0om0sh8fh4PyOtxJlM6eVC+/BtaRwEeZxfyoPfEk1MTbb+DpAzW3gsUv
d6NGPa9u9Hf0eZN3jembavGAr8A+xcqpwNUxcbQxNFK94BxS8OoQ7S6Evy71V9Qw
eOowJSVnNVY1hdkNSU/O7tffpsSBkUCbhjiNO6C5qBVqh1rRnR0fwzFfwXpm8adz
xu1QIsWXVkanNeHhNFzinKSviLm81lqsziTMb/gZsrQBbsapXr0hqBKKP1QQWD3z
qXsODafSk98NXX4D5yuP6gJLtB3bZt74fHOdLLP0XBxT71HsduPqITOyxRIzDU4a
Zmcwr1XfvERjxpoykAyhXTRLSB14YbqI37O687LTi5K/i+BrgDvyYMsMr66ELRhx
FVZmKfAMKogxgEWHRevVAvRNrPEjStQJrajB286QIGD8hXokT681blMERWDCtchO
10qpLg8w0uoWw2aToBu3ebeB4C/8kWWhoYQWzNj+95lbTDcKxZ5qi9zFZCZaqRbB
6bd26GjVWe3i09iAegXMdc1gKkTJJ477DpAn7WYdJEyFOsCsVBuGTOUM/67kdV5z
KSTkYW5Y4yVj0fLZt7/CrGXw2/5MXY13uHDL54nScF4XdT4stNMyj4Wcs1EBEcIR
JC6eN0iyaihVTVskJJ/nnCIFwwPzp2Usthy2UhI+pveoPicn77y+p/ODRflXoB/3
74JHpKT96OstuvP7jBtceRaOmqxIMkLR9LRUu0jua1jcX1ub/1fmfl3ciWcHlqvr
seyb9icaCE4y7vO9LMm2eIw6nYQmfXkqUTGg657ilVFKSvXDRl1IeFVglPTC30ux
W3kkbCDlelK00FLMU+hnEcsnl+px7ETfbuq54Vn3s1MnZPcrgog6acpmIJxblEZ+
3/NN/nR4dhzgVKea/OTYmfZ0hvWohpgzciGqde2kKcXjjuRHwcSApBxHm5HsGhnD
Idz077RJkxwil+IO7Uiav3snlnUxhwe9/WX6id+mcyvn+cdmYrqlOxmW9Eb++EGy
mVN1yjGc8OHUwbSJZHNDPk7eydyu8FqPX4zvMUfWkJFkgqxFFEMD1QqyCG6AyyPS
t1MSvESKbMo/h8g7ZyInuvIQVPDeJP3HHtt/kjAKLGPW/qbqr6qiTI5A8FJSw1Ao
hlkmltzQsdOXBPRJ9Seti9h3Dmr0XW+TFHwh2sOjJX/2g3l2R6RopbG8dhKoZu4u
RL6jOf76cSrmeyC+d9kuwIbIut5hco3qsOWlYQ8njYMlFd+GOJ8EvZUW53ThuRs3
mKYQZ+zUIXjWUevJOAtKT3S8DMYdtHFJ8LaSF9QRSwlVkzX25WRJ4pCGq1PfOd4X
4z63qTSXK5h/jf5gX1deWoWzLamRD7es4Aw/GOxK1Bnjjx5gyIffSVrbpEKzsdTB
Gpi4fIyN5chLNISlNMy7+mgeHTc1v8efvF23XuF6TnEjpOW7kdWtq0QUS/HFzUVX
GiolDwC60nMGZbv2RlYCCpGrWZdvTe7CXxBe61Ph0jr+xm+rSHdBNfutNlBVFU7E
x5ozreyKAT2keNQLCZiYDFW5qmy1bjXV9wALTwfR3UlpBE6nuHa8WGLWmRQsxt4G
uVdMX01AYtBzqt1/wYnn+Sl/rsW634hzL6EfCWAuu9xgaml5L3DP//OmpGNNmYoJ
k8jgf0DLBhC6O2Wroo9zurfv3sbEY1gfQ1aNY0sC71tJ139Zfk8j1IlhEjoX9V4C
e0DkKzDrrIJK/T6FEZ8HkENS9UOQvU8eBgC+R4XayAPNiOe1yu80+0DVuTZmOBA5
bkDhBdQyxTtXxYFB9pQDHN3l0uqUH5nRHAhjLm+YMUTEEWPNNC/p3nIdfS264QYd
rvNEZwKhF5VisaVmkAJE71iui9pYDJf2MX7S0S56TvDwM4SEjjGzdQ1MV8fI4++3
WMoN8lT6isFR5TF5KDM8Hzsmhq93ut2r7UJg1LQ0i7YHqx+xtLXl7sWbbUpeRluS
tjCETLFE56VBF3tlXQpw/e+O3gc/Oa5ptnc+diyE7HrSWNRMqnn4lpTewWus8mNE
6FZ6X5gcBMSuxAvO8Sq/YtHkuq1Z5TvDpz8Qeym7xUO9cgLmbNM2mdaH2htvv6IW
rqvy1xKSXxIM1whn6CFzwuMf8fbFz3sZWDv/A5NIeOqEnGp38v/n/VvHNJO4w266
HEz809ubmUS8vbQ+trIOekkO06+cTciD3wCXfQnfWwxVoZ+4/YPodSybECKjTm9R
jGOF+6Vr6+Gvd6dAlVATUE2FS6J+vPEV0xIqANngW9DQ9Uj+umt+i/8anpFfmVWQ
Leb0zdzNfJhzgfgCvgHLjy8KS9cI2zQc32hLo7xyapkp4/LQgZuJyaQD0g+7rrCk
zA/FIILuA1n65eu2pVZi763v9aNz+jdUPLFPSqWBTG5wBng3CCKMdQYRqo3jhxDb
NBpsgVCcGihNuE2FHuGXg0Ee2f3F4lvbt/E6AZTGttRPRuovle1Da8RQcAbCKyCT
X9ao1+Ge1RrhMmNANrOOkqDtblBEJJAT//XNR39uLBVS96Y9deXFBf8gJs14t+Nt
jIiw7jFu2a35CmXiksnIjDSMc3v6UsT+BJIdeGuXgTz8i3j7i4RiFv2RuN0OstYx
iIrCZWA2a8/N/JKi2lKu96ifrvJbJAzOUj4X4oYOWTCpe5o9R+FZL9DxzIHLaFRO
L+GIhplcVPyCV5Rj5xaDpPB8zfzgBuyeurt2nR7g9LKuBz70H4JuEkQAEV7hMhu1
xVBurnlxvw3kmdQxhL/DUy5zoIctpcXOaZLEx2StSw8hUDcksNFfQJ96wa/CiSmz
9cVzu0UbPnVsZ0QYd7yhaw0ZIQF8t9GMpA1Ct5r5CCNIuUja3aMedyh66P2x5Oh7
G567RbmzipzdRPuYYahDz2agOmJvDAhl/E9EzhQE0VNLzr51BkSrMTe2YhxN9MOC
9SnzHVauZL7HyRAmcNsuldpjaVqu+wMqarn4c1dVuUnJQZC+6NmP95/Ew28cneG0
SCiKjkIKuiBB+OM+hA3aZq8S0k5jfrcG9ChNAKprdYXI2o+3d7MQGGP4cEhDouUG
WpcLaM3WJIoMTIvcHr3Kb5b317mzAKY2imzF4vMEaWWhBJKN5VicPpoeySUN5v8x
wWdlCua8KS99HxygK1f8ZvNZVIh/TFx6E0Yd4Pt2ER3MF+lb+i1QmaK/0gW8iPlW
Z+inNfkEXxdnRyVtXrXRu36dejQsskMpO4z4vnmUI+4LMCnR8GPwgwnA/C85MAlY
D0x6cl2ef5mCIU+RgMGLgO5AeLgYFCLBMMlLuZxJdJkiHn8UGUypNvLS/W7jtr4M
ChJU/OtJZBuXYpQYTQ4MwVhjdi3+gUHYA05QS11lTGWNEjvs1nD/1RUVxBuhXvV2
32KDjmKhuR0CNWZmz8A1ENULK5KpOz+vWn+bH7UXdQqQScXFjvQi2vwKsvwB/ZS4
DF3AMKCcIHM8yQu4cd+bAeAzBleTtBbiAah+6LpheETivmAXlP6rz0a7x7T448YB
32zdqU3n/6dY0T15zHrPpJftkC06EaWT8An3xrYNcCuGR7AtVacwoODgjd9En97N
5Wwmap74sPN0pq81/zjdkcte67Yj6tpcRRtlYUDuYMXCvE2aoK6dQBllmCl7Blmk
4QNl0EcOr/uySvzfrnZDV7NbKKAuRsRA1Txeo2Jb3bo0WHUL4Ctag1f5aUkc4D7R
j8i4+HZ8dCxzAOQYKNrUwk8uDxLo/GB9AfViVGLOPFFdoqB7ksLjVopN9t0/KnTX
A2sgDa0sfdvq2Sajlsi/CV53yG2ont9UPhrM4SJj3Syu19Qj+sAj+dDi2uOCsFmS
RbaYHqbC+lVdsQvYqq5r3oWZun1/d2Hrwg9xaDYNL45nYX5s7acfUdaXJ6eqpxZH
/kfhFRtb2HbFuTgELNYHXG7mwdOQUGbG6Fl5/eg8sgAPLlMUKbc7ZloH4f91q6q6
c8fwrz/CK7TBiHOPL7tDxrIPcnSk8RKO7BSTjDqzMT7y78RdIp2DsCiaZAYAcQrw
7nSzQ6LYeOaPzJgjA+nzObu3gp40G3I4MvVANjsZxNkUlGI2Vjbi9uIG+WesFnUp
OgaMqOu0JjWEd4edWbWJx1iLwycljRML7SBbwMihBKm2Vrd9ceHu5HbDGaV5uTzE
B+BX/T7PeQgosXOVL+i/zGNZ0Fm93cZZpDdn5hvD+zWVEuxjjBwKJQVFnr0DsEdX
V650vONXMis5zD0dEu/qjm57IO26A8xACDxTMAHWO/bRZ92zZHnwpCATYTlWKDu7
CbblzXUF+1AZI2ic2O72dYvJEpjYJxd+OcsTy6R5QQIl4RwnsYRNebhk2Z8wj/lK
SVDZZ1sWSXWCAP8e8ytzLpx4L2b0B6NhRwFMM0MSAzFukmM5YEr/YH/chqRs+qBl
oVPQNldrfsXkRO5DtNJIR7B+ZrltVC3CtlOQLLYyzAIhTdOszHrrUALAVGSZYtrf
wmbTppjAzB8flUSp8BDdPYqSjfETkzqGCnn50Sl8dDDCvToSSjj55sqCrZ2iCmBY
cxEx4jbHZ4yjQ2j9f6jSVBglutw4kUYKeUGS+yRaY1gGclHfG0gJYzDpkX2KLTSS
4OoKccKKHw2LBMwiYmWGEV7NypDWhPtbrOFIKBFqK60Y558Kb3jU5TAARZMOlN77
jqtDB4Im2jKQcQ/lzhi8BEXkA+tY5zVK1G2rMt7Wm96vCWghQuuFKkbNPLaFG6ev
fguColxzwKF7ME5lLDh4KxBoXJSDFZA/iWI41mjqCh4KxkZ67FF1MXy4Y8gYdOke
oG6/KKm1WI2FbEnNyan9qLi6X+j2q+In3TqeUMu+ktYyCOju+IZKGZovYqqMZvpE
AScPd1sdF+TBvqWbpwzKJUzSajfLc8ntVYPLu3lrXyhjF3GJGRCqBttpmfTVKj2q
YN0KJl6RFHFQ5toizFqNQj4o0nJI9bakAWTEG0kC/FWHXXLQNP1suvTuDaIjp9+f
fMQSD9fuKiCEvtjPkv5WQdfCn1buK0jKD5SWg2TyXihWQEeQ52g4biLvKYLTwkH8
9BldS7XrM3bXDjKf4Gj7UuEJbOyFaTi+uElHGAv92oFZJQOorK7h+W+YmXADR4By
kW22Jufq8QNNhXbhfZnSUUki5u82gV0KkF2IwuTlfXuPgryH63VyCARq+AYi2U48
24zqBDp5qZ0pjpJN0KXN5CI29D/JMogG1oZV+nbUP+qsk9iB9B4spBu34JD/qWH0
WX6DTCMkGdLCiY8Dwekoo6u7EhKrdb+Vme1D0UAyax4v1CcxJVDgMzJICG6cZjXi
YJo22U+i8qa3SNqzx4SBgvXF2JFZG8006ufDqP3H/oZFgBZmYpIWeI4pzPGMg3rt
aqRMcDJTxDPwa/3Suy07chONjh0Wg6M3ix0NZdlg8Kn2IoW4qlYeJ7UI9LTFEeh/
1vvYhQ6nGpwS90C+tfjeuwR0S7DL46u8SCqGmdYna1rYnopajXvSwrEfCDPAzaz2
+lwsFn1N6jTWMVWGhA8h60+IeRsVe4rXqaAchlsvEa6QXBSFVwbYary+hz5LAOTV
06NJ3jG33DH/owbDPCbXo7WJf5pWi5HRLyIuTf3dT3Z6UTD+UzW0NIk7YXPkJv8n
4pCCa2I78k9yTSvCQL2uBkQTLquVpL6ggxSBhaTHz1UaZ+xTmsvjtl/G1B1j2rc2
0uDt+iNOYoq2CaPP9D/AMtVzNKMDzWfzBXvsJRcpHYZPxsMpVMEBJRbkbP6mlLKM
NVbuEz/px/SM2LhRtJ+jDxPCd5FKtRK9OQeRtbmkn0YhosrzK5COM1PVvQwsDaeO
NVN4bmA12otS8CxPIHTuLN6Q5ne6T1aV6M8N2y2uRPX7NtrBSNRZzzTeR4v/kV4m
eeXv0mFsDkRIr3hdLptmEyKqBkWOqxVJ7/ZpaLRPK3MhckS/fp0aQaEMftXX8ES/
BDfE8rB2Ca4wFroePACxk2pzm08SKLF5XTi8lAY963qijvnoSUmPjC1ASTyIXB96
I8ObFxXyoIsBge6KxDOH16SaVrw/72rzH8x28WwBegAsh3OWeAQ961s6LLzUNqtY
lsbL5kPtbS+ivh17pG20QHj9daatBMt3ZO9NMth94tKQICyEmaUGrQKvYtVC83V0
gEAnV5n4YN/6meAlru2RjuHa7LhfLDAHCB+TNtujUPP2jjx+FTZrw3zXXxFux8Xg
zVdJsODK6Nn+LOU80s0F+IkZXjWbMglbCNkvNMzQdZzekcwOonSUnNr/hy3ul4J4
86bfc8aK+rYfl3zhIIKiVxogu5hSBOhiRul4gALj8b1FoxsX+LVloZEs4XlSTnbU
6rXRy1F01qzX/bcuf3gHeQjQcYonM3m1fY8DIAmRlkQNL0Y4ugZy7f1KTzvG02zD
Q+UcjNV5G7LugnLLqPyAIwcKCJehACRNOb0wCjkd+w8sLpP1RummqJoYVWJZ5WE7
E9fi044ud02tVnvmTlJ+tZ42Qb648Z2Es3LzLV4JATuiKuiRJRFEpSL/k/DreLX6
pE1EvaRz/C8v1RHDw1kzYfNjlwftS32UCFJfIFdG/Y3M8tGxCkiiheB4JgQWE8e9
Q59wesntgn/9Av2GkUEbFS89X+1gYbWfRfRmAAD48XlvzO4To1xhTA6Jfr09qIwq
m6okikJeCHaSl54XNIF700y4Uz5fUn7A9mFQaP3hLRs3tRRgxSMCfz5NQcW27/8a
9ibnXKcQ4x9+HXE7Psu4mfb2IPtqyDfVJYQjLRy7fIREOVx+0MPbkdbenn92jy4h
GfrSq+i9KxOMHA0AJqdjNCXfPcJ+Cq753zWCiULS6hGT/73l+ZNiF5KR3FAHRATq
xxm/KYbxV8H3Fzz/Ia7oPYnwesAl/hFfHCFa3jVcFhiNd5QfAhVemvKxF3+CWyqj
oMswIl+w9NK3rMiTH9ogGYcmsR8EfXWYeIONJ4HmnaT4OJWqCe3lSGmI5EWKBWai
28hYiLElLKRJEUOWKdu+YOowud6qNJgCZfXE8MGQSbuUL8CN9MGM4e7iXBZLYEyO
AkD5hHoTaGsjka7SseDQSxIRlLGhmGgOXTq2Jt3xBhXwTmCmfJYPJpAFL3Tjs2Sv
kdkSCziFPQ1mQ41wF5Zs0T2cvHCNo6pZmiH4vGOr3VvXjJLClwKQxY/S0E0hOkdz
jwr0b82+5o7uoA9zOPo6PIFna+ZtVme0kg7NbaF0gAcxGJ3n1UV0oFo8r9eE3DCG
QbtmeKNBOjfImhxGThSZA+ETimj4s1ZzsF411TK4U7NrdXelimL2eN3tq5yG+ODB
SJe9ZGlB4IRTV0RkctfDsI1N2NPnL7lylAJ9aCHyaFAAzE2T6M5+mFWM5aAK6ip5
IVfCmqa5Kruv8THij985ejnb+nkwDOJ9R0AlfbrRkoNMbPA0KVdEab+H4N2kMVFO
0s7CS9ySKybWtCygqKcNuZhxhWyI0XKaieQpp7Sh2opyd2BiYWoKZMaWJp62Pa6I
LdxDGSgD9+unvqN+vhxwnbaV9mJLdYsHIra8Tjf6Kgw2GCGZzF+1CVZf4s4nZ8A8
rByCJ8EUJXdV2O4OZxwASfX3MYtVNFBldlvMUIMSqHkdIRWwVjVBsLQrMV80wTK5
/MNJCs/rwxY9IXPk4tgRs91exXC0V7q5tK4VrtpFGt5hWDGxcHq19LWeb2QSiHsG
0aauIfX7Ip8OMiIBzS0pzaaaJSLstMjN8BzcvKY1a/BVaRz3zP58NKGZAVHDejDa
rVUx5AkU5hnh9cFAx5RybPjeS7J1HJ3Hx13yiIM4raQcX4Dxg7p+XyVv6Fdm+uAc
G9FXa5VhHoe1cxX8QnmtqZJfRvd97OduWf7x1/b0FEu7GgOuVodRMd2R08ALn/BJ
faqIUsYR0mE+F/7EStbnauJx23/jPxx9lfRKALk1RuGguc/mKFMkChbKL1anKJsZ
VHJgwEH+XaRMzH2xoxXAFFaEjCVxKlYvWFmH5QGhp4Eo/ukoSUcaunQyhHJHAtv+
Zj/0C4O6vewhoHNmoIyXoVoiDYiOks9ZlOhSpb2ElRTXD42QSQAbzG7Qxar5pbpv
5FEy6XUDDYFqcnGNzl01YIjtX5nAz/zOws0v+/nXKUTdMa5sryEr7smA/61hg0go
OQN4XfGlDYK/ubzVIN7weB6dVmA2GYfWnZCxxDjf4siu02HQBxIwwPfCyWDWEfdi
+oOXxKHXOf+U5Kbv2hLO3f7ahMARRoNOmXga2Sq3coVg0mA+ob1rlgRoWY6kaqzD
fzWX8KPbyo3XcVslf0Vkme4WyIUJjH7IAVdNqcID8KD+Ybxnor5am7Y/0849KXcg
hmibter0URI6l9w4jaEZS4/NHpe1LuSrcpXDqRrDUmSlE6ZvxNbnP/RC+00a1M2u
k8z1JKsvd62FrUWsJjS1NntiT1fE6uIseSwcBEDw5DjkHN3Q0BAtb85Jev3yo80n
+0Ia/7ojGrEUSAk1gJCnLY0y2CjJTra3D9zVUX0162ZiFDo2LLs1oo9aZnAp0pFU
jmcJUH6xfBYY4vZsOa+dun4SP9g5yH3EmoZC7qahH0N3uuBPy8t0IQgZ6hCuV0Ty
DdUV6CmP/pP1jGKhpMwagqEk5SV93P7hN9e8lNTANZjicYYCQsJhymhDUkcy1k8o
ZY+SBU2Tt4LcQxLLaUAHRJknZpOKfLUVVB77D5q3/YUFtKSF9QVqOCWtjDr15x8e
uwB712kPWOp8gZC5DASLirT9rPnLTYYnQKb0KP/dofYV4lFg+6RgT1cI80m74kNw
peKYSKeEqLfje8UxDtKEPFBtpxGeSn+7cRjwCjtBDaVv7dvcWXT0umSvlNWYapff
8MDMoCm0jvo97QOsUYwYCyfMsdroovz+GEbi+/tXl23crY+Fiwfx9/4d2pvJhGos
B9olYA8MOGsiz0TcIha3ZoTBS/+JeU2FU769NHMF02X+6I0D0BZgmH3JxhFElVgP
4BARlWyy1PSJYY+eOyPulhhjyaxvVqydit79qXNfsrqF5Yl1MGSxCM25ub2liFUG
IUwcVehvT9+a7dWbc6Rh9+FCeXf5y497D31Lp4QmzWCU0hBOXDUyM07yFDOA/o/4
8hDzTdZ3mQ5xS0do8GFYbx066tmPjSyy/IaDIUbtoEr0/hwt+6cFg6NosR9TquBI
NMgynAUcweKsJcjCfY64J2TGA2I2r7bgTObrGTA0NRwZ9+iV1hdTb6Xc+eXJp3oj
6GJFyn6AAe4UkQ7/PPrUiuu7kz+KnhKGgXp0FZDRBHSi47SS9GkHupcZ1Z01HMqT
FN+VuSk9DKN1xuFHR7NsZHGZs8vguUNgucD7isaJbG9ke7/son20JEmoHqYmL+7U
c6FQMJHlrgHg6uGsvb2I5MiV9zpBh8elpBvu4aW+2dXqDXTe2H1STw8oIWdPARet
v0hdxZn1Gv4W6oelvvSkP2j806C3uwg17vbxgkVujBrIdDjODR7W0Ui7+FP38CfB
+Q3r2X4AnQPe/ejjy0XpuP0u9FZ7rlgl8tKwVc/6FBFoncvT+AHN33KQlashSlWJ
pzMzl7XSdMF2TRRsNk2KqyBw0B5G/34NtFyhQOvivv9X/WNTEpu222MREJoGxxp/
YplrreMLoxLvnrW+AbPFzxl42h8yEJu87HGkMW9yMYLGft5jWOZGXUOMf0KWS4Wf
Eo8DvXNu9G96kC9bBvrFR3hWthqZI/WLPvJpJbxRkaX5kp1PgXLTTnP8yioNLEem
+l4p1PYtnBzLBNv5bcxPmE0oa5eNkNTRyq91sKkf8ECxr2ns6CYvVG46o2ByONmI
ueIgxZWSY2C4lHxAoKTOVZiGhKrCSg37nb0GgsNa2ZqSA5WJzlkrawArVnkUPpAo
2CVCgj/ApElHg918l6/PWEO+pe1kC/6STKNNrcHmkT1MWwj55yq2fQc/bRma8knk
quldgsmbzRMqSV1s0mesNSTIWABiqEjumuhY/Fl+tX8feypABjLx4JBX2YO4Rc1J
/JIBNupL1z7TyUq2h/wBwL+hme+td1KHsSI2OQg6sWd8LDv1uu3Cl4WXCCOMEEyD
LVqgY0MfnfUxfdtHUSwyxNhr6iCGcPxcX+tYjhbEcvbUGBZoV5iXNvuGWf5IbhPA
H/B26Dh3b+nBjrr6MCiWPQak8hmP0XlTwDU5c9D6tkrmRJQ05UBVjinrlOdlX3Tt
1hA+oppINB7UDVgmHJHpMRCuymU9RGzCt1BO4/SB8sQ328tPgRFJlLmGu3MxnczD
Qsv8ftqbXE75oG0/Hh1OvbkWus3MeFhv8N2zQaVeo1eq+DNjxq7UTGv1qIkDRuNn
kwLaf/t3s8yIFVSINt3f7CMkZnpcD8dYd0zXPzkUvSSUUwgdLbMen/BlfoMdsTi7
gvLNZcar1AXrt5Fkhz8/0o1NkKr9QxtmZkIza0Pt2bxjyIDtwyTWjgMmzweUT6m/
jzijjF4S4y8tN4bJn4bZFFKFoWMQQa8y9tkab7cA88wj1XqYt0f91IYzHvSfkQLw
wZ2jMxSdOqHmlkohwhwxhyllomC5DukcgsZu7CigA6hIDhC1gnj5vvKblTSrJJwD
7u8ED/1kXthcmmImk3GeqAeprQfIJv7/zKo3v61V09rDpYkMWW3fqGxOX6KvBWe/
W11852QZ6Wf32iQy1kqbCTOqc0CJd6ZMv16cv03aJhdcDuexU9B3b1PGyHvHH1SU
ZOTSL+gqUcBjabeRxgAfL1NY7OTtOgdAjTAwOsMUXkuNfpGwOIKw/xXtA8p8QIWQ
kMiGA87CgLcgXy4ILJKWPlFb1PqQjwHFP1aq9UDot7Aje9n/Xm2EiFtZYRgPdj2s
ez+BfdZ/5FljEpCUVcsEG/CVCn42jMqfsqx1DJk7YL85plAQzH3m86n8jDFOPDO4
D4J6A7L9eQhup8xeiebtCGJtoUh6We+xfFxZfUc1bTXTopjFU8QwGSazsubYzZJp
BwKjd4bU+2w/ylLSGoO60ik0V+sXjl0LMXx9lt5sXmjqRByZEcsE3rpfEnKSR7wS
2u6LdALCXUiEwqG4t5/xThlM00ViOM8H3PjMKe3tzqBkEKgQ9nljaxcrtBEwdcO2
2AfeRhthRZLDp/zZwm1r3gdBePnYJiE7lV7rUTgwHwy9zT4r+AOu0zK5IgFvzeoY
Tcz0PH6wEFQ0KE4rKK8BKnxwHLrILrMbO86SNTy575z0DVRm4helMd8WkObwqwP4
nv9MWWjx/YMLfblNB5yRM3GBdltMDiwOFsyUbPxO8XenRcP7gVM9lGb+HVbCXRBn
Rs1rKr5g79WKnR0ZtWYj09zFeJnXk87LFhs1qdVND5wrv0ffDIwcH+AECsnECxVI
VdgipGPsFrqqhyYVJ2jutt9k0/JffqyH2gRe7aiB46b+W6Ljd8PQQlVEt/iQ9ZCg
ZrTCSVpGNKo/PXaFWKrO1oFhNNkg7tgyRLHbcY90EW4AGG4fy7sUnPHXCEicRQ/F
fvERBKTLdvIrsZyW8wjXHWoRSD/nY7HdsSGkYfllaePiog0FSW7vkvNsHY1fGK5P
9e8uh+9plwZRmy2e9iMlkdAoC7b7ym5ZDbroF1mnA+cIQAOl1B5dUzGzODrzRsp8
/t61dKTjcQuF4p6p+Xt4mxnDQPR3KUVJocP+CVsYSYWvfddbbHCqlRMFhJ+43U6W
kernYYuv+tErA8vU1qrhPXYaWZC4W/ufhpMiOHTuICHXDGbGhoJCB5ENXiZeQU/V
IQX7binpmi2nBeaTCA1+i/jJPMpkNn2jo1Fcc9YJOgho2gJi7hqqDEb/JmxLzdCO
+SHJFDjvWHljYByvMDU0s/RP/QjhsnLMGKKXdakV0fSHgFVAC1eZR18HmS+Fvvic
6juBIGvURawr08Diry8dsfidrvFCobhzfO99MYoP01jK1SAwAHHx4jw1QTN09j28
W6H9RvZw8nYm5pFzHc5h0PKAsZE0+BbsodxmQi8wrrlzCaSjqVmQfEASW/NoQYpq
rffxasDY7W/Sp/MiILxY8OeYsp1fnMItVQElTm7+X3yv7JXzZi9feDL7bS43lweh
aE179pUxOlqt/t70IMWYPjL1Scga+3nGKuHJdAc6VqkXfsftIReQqK6tCVj9D6ex
cM2xGQZMTKwusavikCi75BsvCk83g9j1OiKK3cfOWUeyJi1K8htBhGPGdQCRJm0A
Exyb7wFS82iWj5s/5clkuj4q0DkLP3Nypaf1OGyO+5MNkOIP27m1fN8Ld7lrG+HL
1wM9pPJSyy7JRIKxED2lXJSAFQQw1/JjEeaj4pYe0py2GVxLrs8K1dgvi+9QY0gS
qbaNyM/N4cXz7u6tF4E5jju5wMaz0FvwXjciNWhKjRDRAYtXK7Ck2LBfHv3elpJh
uBZm9ik3TLOwiOxL6euy5veyBeMxJG/dPv7aMmYtAwQfHHUIY/xvqiJdU1L/kL7/
Y+roiIOQSwGGv/AG/+4tnALEhlj7Ggjh868X0EhvJkOqO3E8DjvQI9b+lXVs+bXM
5H/OUWSgD00M3kmV06CwCoiNfnOmhFcAw7q3rJ5ItfeFDSKxAyQM1BqKywV1yQDL
gr9vwSmgA888ZsyDhq7YI+sTnnMk3lC07kEDsF/p9TQNtfOzlC6PYnojd3YUhaKk
oxyKCE142UiDqGox8muzh+lFZbvO7aWl/P10nox9jTTa5ajjwRjTOsi59A4iYVeq
A8ZiKKjemgOheE6sJXqfnUsp5CsXwtwvQID60DVUcJXK5T2IYeldAg70EM9TOY6A
b7sA23Z3HGoXG2CvEi9iLxZeQWxVZ8wcdOHoWl4hjafHh1V37I4Gi3r/3F9mlxFZ
HmAyqaavOswMvRgh8OmM9hWbTC0XjMXsNlkFFNWLnVX2zGliDqSYVC3aUq7PaiWQ
gw91lJeOEEGL+/nJIxP7IUPvVFqtFXb72nhyc5SmNthuYF8lKJsLJigETWNwMbc4
+L2gKoizEKHFrcylJTfhX60F7HaIKBxRLBsaDaaI853OFvfiUbqDtM6n6TczFBqc
HqN1YnV+QcoL4SyhQuBdRVkyQ7eNBvgilaDyNPJFNWP6hSR7WgUZeQLMsuB+reyG
grUPQIrf8W0LdG7lH4tDG47DKhBRdudYR+V5bqmeddSSK/JJ42O8Iyvov4oraHg6
uTFqWk3zVjyt6At84OKLj65pXtWA7CSaDSnMHtv0W0KhAVJYPqLT4lSD4KH1YDIz
Q71aucHU3LAof0zjC1/M3Xe7C7rVABc736TEixx9rj3Ie2rODhsXLYhrSADZAfWH
Yq4v02TBhC2mOmiDgF10dFTROAxC637LAlRZnbMGn6p8CA1grNKWuxxBYS09TUYI
0SJIigrP85Cg1d0dj55FYcZGKEBOgY3jZ+Kf5eLP5WK48XhO0yBVkxWl5as6Kdfn
2GeE292M4qTYm0UC9CQw+K8p7Kg1d306PtpdZtBhlEde6+tLgjwHRhO6ZL8x3AMf
2nt1YiINFi36SCou7Zn6sGXwS7zQglpif/JU9j73VOuFrP5iM5t6d2FDQU2HJerU
hVg+l9t3MrDgdwwZMpMnerO+AyuJOS03l2l7a0qRn+B4HLPw7BOU0aE6cS+Bf6rH
pQVQp3yqj641Su4+/VlBOJA/NgCByOtgLqsc1BdCx5zKm2sx2xv6meywo4bgF6Bn
EbyTaECsbJHsn5Cvn3az7T/+9fECBZ3tGnov9LL7vWfmSArP9rqpH2ah8j1XqvYZ
fC51BICRMeNLDmHhI4MQMVSVtNRAwR0n/NIf0gzRjlxI192okfWVj7AZTU6gN9LZ
TkruLcize8l9Hm9rUVSj75DzHvEjb0qAVEWrOY6oA9zQ7rZyI7awdmq8XG5xQYln
n99XaoKojL0mT61QtSkD9Cu5oTFyMSPuGCnujDBx1Y3CPG00YrHB94ApYu3/DJcO
sYitKab62lRO6aQxtYyITAwKeyuxk9l2+dL5L4iTVBoygN978XCGYPMCeL5/wg+v
W85zfqaBY8vSXspLvFWEI1BInGplgwGmmeHWCo4Wi3XZ87WK+1T2sCGTk29pl1z+
Nr4JzyzMof8IdYv0cKzv2AuaD9hSWSz/JI3uMLye68Fu1mFGE87BWQ/LjDxI/xoY
vx27dMfKexA/f8MKmRnt7dxc+KkctFCNig3nlOr8tOAxeCGmyajItLr/hlyMWVwM
ZSuwSy62VV8EAn2+VpbPNq132ROn0S3of8XTGPvQ09ib1idpRpdplP7cylBjk1BE
AV/elyDDPo1uAX3UHAvvET7tONgaJ4kH/txzTDBZLWGxEjuLF0bolA7kVNofo0ez
DVa2UYtOtS0SBOUvm2XXdyPeHqvMsmVNmOvY+oS0p+cxU3p+BdKivntOSsqBl+jn
v2ZRm9V52cHwGip8NRP7nmkjHthJFSwB7+5guZzn32O7fwUcDIq8ujiCidIt++3u
65er1pD0JVUmzCZDwx/6Uy1tyW0szghKazxkUzG0hI6R1+2AUGUERls4uay6McNo
aWOIenzqy7LAE+4DOEsMIsBLAAB1XX0ihz3BHv+Rt8tbf7NzibVTGyWgC8Ws3LKt
IoD5OToKwzz4Wvae8/Jv8V8brvtu//5Lmj0bxV2BqakfqfH4F82XQyCHT4Rcy1jl
QwUahaySKiCHycD3ZQbNeAZLl6G/c2ze7/Ij01WWufitMAM7/A8907wWMXpwX+PI
LemafJ3M0ZqSlU4I0D5R5VNzdKt5zLt6WBcg2E/PrXpHBytxC20hQ6FGgWYBKUnw
qUxi03b49aElfLn+8fMP0/7NMEa+TLstuI3mbYS4qH4KIPbPFTP4MxWXVbY2o5zt
o+/w06BBNp7Ar4obPPv7kodX+FZyniCMCoWWEJpQulYKoUBrQxfDTuu0e1idfJQt
FT/gUz372Wy768KecOE8LImEJBDnqWdQtzLc70GX6WivDQja9QQ7+Kmm195IMdLg
kNeCXockhqPZPiaftLQu/+FxrW/f+w+t/ZMQOCdeSMtGuO3RdqgESzr5oM9DCnYF
LLyotUrUb3D7+9qGSSP4ypt5g6S5ie/Ew6rslbW6d1xY+0xvyKc5zzeLr3eIkSnM
1b+DPtDKNGCnRF/c323Kiv4vhq/JKZZmN2Xu5hvVWeMDEqIgF64y2GSOEWxUlg2T
FHGrgshz981QIwAGvrJuPtimXPImdGs2nIE573uHmRMIvXW4zbs5ZeE5wd11wnOU
hoB+uHbdgfXzt7TRttS8Qi8iZ54wykKV02/I1Km4Kqzt/KQSCc8xnagSbi9sMVCl
SaxpB7G/5oORMbyeMCjRJH5wPO8zRL+EBtBY1VEgmul1gmnDQrre9ko0j8Cz3caX
mw2xqM7uNWT8tQG2Z1JDbkV+7jJAGz9i28+9cM34wYr+5QeHZy686b0vmatSLpWZ
zyf4IEzNehADeSDPItD6glnFJRWh8z75YJ/m+ArWlMHjPmvmGI0V983yiAYldQSa
z9JzeuEaz4EAEatmNgTHZzKG7GWz6lBoj+McAiDE2qEGCHRc4JHGUAZ5FKU3338v
70exkw8gKy7E35qtbryBtEQbWFlkPNVP/Ik7mg+xDusBI1q0IKy7r/pFagGXLN4E
i18qwpgtsWrh2YkoFFxUe8WtA/zRoMIJE2XZmEGuecYvEsmDNOeNVrrouQfWoJK3
8Ma9si06lx3ijo7oxiHgO5UXzHH4VBzUMDSrawiFRYms3Dr91+oQBHfV3AAdj6kO
4+wrffAqri67PL0JEAU4uh0jshE2Rrqwhe+ObP5HIp/+DtnlYrpPTDNkPaquZu8E
5SuDNqGqIiU098+HjOUIaRQLk0B94L/MgsLhTyrpdv6E+IIrA0CR7IoiES3ELBOZ
PcLD7UE9agwByqk2WEv1yPaEy3CsNDgOoVyeawuuOklMjSIbvtTh1BYVXEXD/V9A
e7p5d3oS35oK8WqB93K3VY66YCe26uZD6/vflnCWvEMxPEPXVezvm94S7oBpCsvn
yrO9UswpOsYBU3D9YyRSqIhECwwBI21sCx9AcFeU5OjVB7MZo8Wf4QAALxQ6nsXq
QtbDXfsmkZyslQjGQF5iRiQ4dzfiZb9KotrJ2E6vJJfBTHP5WLIeT4c9TTg33k0b
D4ypo1oyn+1uRLHht594eq48Nh0o+it5fRX//CQdqXpC9kWqyrgQLe7txuwJpMPF
LTkbUEjWhJidgFwu4gFa/kkqN4tyc9NVw6xWa37hyVPyhI4udZqcfk17BUDECPsl
cBJkebDPZUExyFuLI6bxwP1N52z/ZpI4/C/eUAtBPDv3jDBJ/tGLKPP7DbK61+yS
jRWZvIGTExp8DrNDbGSu4gOJqkMtZCJMp2Sk1V1SKrmV0pyjQhB657P3wNrDTJlt
E4yBjv7r+y99i2RP0VUdeWrruQRxIn6hSGRdtPKZqojeuBCjxzrMDl2PSXIm9Yt5
zgRCowUgy5JaK5zYKm0LdniuBhFGGesPqEqzkEj6q9nScrDjErtdSVmDCkjC9N9G
6sCoRMM+oP3WX3NJ/gl3lNFKHecUe+Eipt06zV2ClvkKQeiPH4D1c0GKNXN8nBGn
SMZC2Q8r4XvImbiA10dLWm+y6HI5b4oVPOVfNcEinxEKM9H4DYNU1kUaUy2Mv6FX
55vMjlr0VHNpDOqz+hgjbo9Di+VYBVVvMu5zNpaYJSojbtekMiqbEKvkByHUOYVv
V6xgIuJJUTxrJFE1O18u4XCtGvBQg34BSQEAaLTNT8mjXKOsVYiAbNRCSWDTDyrP
kQ3/DrCTNkJQO8lPj95EF6ElvHjV5aAf3b7EuF0JF3eYI8tN5X+/uwzpSqluwDia
67RaH3KYuDK3VfK3s8XPRUxQESDQz2DHjMzSLmjAqA7e/fm7Uf3RxrbtT8NeCfuO
wjO3MQvJR/0EU9WHfnTSzDPBc2VkOO6GRf+utx4Ny/gigHoOF0KstRqFSnWKfzdu
oc6SUtVa4LB68Im6/gqtYwGGBmfFkvI82dkY76hn5tTswsk8N+mtFZIC/Tp0tQU5
Qf2cH9ku9RZPh59cDgffyWbQNu67aRUSHDaR6IYCn+PYzPDvuNtrsMXQu1iPaIR7
bQ05Rcb+bCnuqVPlOJth6ro6sb8e22n3lET+fZOwFbNq/AgxcrfZIk85OyVzIPS5
e1cJdhBPOiggsbz1TJ5hde7W1JwrKLKKbhNdeNSJcyipYm/KtlGZvKAbfIHDunRG
0n+QksuxLDs6A+MT5JEA0zw1xvlrCoTNICF2Fbb74vR9E1BmaXfFaD9hGXxS3LhB
qhlwcfUOmms3eBxbsmx1agVVnAYrb5eZZAW6n/e48MifnPpyUvi25xvYtI0uzIZ8
o75vAe6wUy5oYx694YA55htukyyzB+zcjms0djM88MPygL5pf+d1bWP9wRCRd2am
usDnMdCQuXwoKkfCfnmuiB8Syu1FCISiDcFWAyORw0qdischAHhIuiTfZeFWrEDS
IPAsUm7gLBVD6ALeFf423AJDL6BxP0IEPcyTaOuTI0cHTjRzP+mYyfhUyiV1v6cg
ZPABhqjmQxNtLMGqhY3uGLSDKn+tlNyt9ptj3kCRuS6N/qL3DOzpgyPnCY5XfdaZ
qowekz3bMofKq7yapz2d6aR0EdWkcetwpMEvm2HUyRyp1hHi7PO9xkv8PoxbREif
RiODJsA0lqk1WtZhawM0c9r4fbqRzFwgGl2BFcPzceGyj9C9RI2uXm4dT6OoT0XH
j7mfvaQF74SZzaG73/y0iRDPoKoMnLN6D0/kTaPnhA2IKDlWTI7v05AJh8dY6mC5
342TzTPdvVAxZgsmEfxShyw+gunQTcgulGX12Z6fHccVwN7q0GfhF8IUSL06elwh
yR9tlNCANEzxWvH1PSQ10yPgBQJV+ZYUsiP7I7MAJeCUGdTCEuzVnGr93Ctq2ugh
CxbF/Ee/1+V28CKHTkBagEqOcH0yAHLsomW5t//sPC9T1Dw5a3QXswlQ3kJQDOVS
LR/ntaqqj//Hgx7/PhQ9oJWxgGGw+PGAwSQPUAH1gMiZLYMNI3Qs67dTIu5YKTWS
3p4MbkGsFU81QjmfjcpIj0Zal+AmPiym06hlSIOlN/nTutgZr4+Lso1rvgUl6DNa
Aij0D72mJ9d9s6pyZ7XUea/Rm535fUSvBf9jZFp/qpOlFUgCibRzQ4zq2bM2HKQ/
0TPeWtEmHJUVEmfAoP68NdHAvWoo9lXP4aVPjSoLBF22H2eto7xcQzZZLmjnkNMF
Hd6v527p8Vr6Ga+l46juD5ar1prk4yNEV3+4e0peU7MI6NMU/iwtnN7YO4I7tH1p
fcR46BzqBxWdcp4q6PxMoe9j831sSDAvjHFOPeDYVUHm3S4aKeOZt6zmxHqWELWt
PAJ+zGjfs0cI7jrPq8Mzv0u8yZQ+FG31CpYdI23M/lzdvkXogxduDhOJdrPNMYHB
ilMHlD+dmlEhlUPfE4ln94kFz81l5gWn2DpAlWJ5XPqZ/CNO2TdXTXELUGoPG/jk
j08we9Soi1mlKnvjmdW+5CKIt9Q6BDGVqUCCaSviCtreCE/mSSSIDe+0mAwWPua9
jmhJpTS2m23b9wH2XbFx3RblRWRE/YD/FQzyOpDycKyPZH9mpjlD51NjO/IAMq6Z
MidN1bb+QcRAzsA/JMePL5K4XUU1ZhP/IRVwHlJLK4FjStNLFBpngV+1Nr7RHNoK
M88VjHlqA2rMNaXYTkXGFmcz2XdpzZEHr0OEpTu8Iv+OQsou4c2bSWlv3J5UZpzq
RosqAw9/Hatk1CFuYwe/kuydytEvwBR9I8UM8/aQaKiRRqrYm591V6w4HyE7wbpO
mqKdfvvl44eHKejEYzxlb5BaZiOlcEo+bxtsZN3dbt1IgY+pzPAisAEJumHN5oK2
96F/QxGK4VgVPPXFUtwsm6NLmyrGbYRp4/LWAWAE1inMyh+rXu8WFH046YTH2quO
M3PuHH9b9RsyUB+3KBSNBhwK3Jax9wBwjdpbKR4rMh8OTNWnWDnQ9PzznLwNimdb
UWGkGhqLrFnQM5bWdf+UgnPIz3flVAKvO4hpsxfouU0on4TgNsHxmkeOUPAxFFN+
h6tKu3FVLwXgw8U9HoSlzCyTFGES+vxKcXUw8H/cwggpbN0DrFp4NCGq5hmpf1ZV
f2WScszYRhVb6NXpc/nzBMDg0PG/PCTD+JtGhUd76rh9SrdgP6sxFn89NDFQlx9g
2E19JYyVhTgMlGRXvKjdXFovHMVCJ2BSW//KcS2NivbpOlvHrhEdEPH0njlEJkXC
R/DNtZJABhRV2Zs76anluos3XPg0KUB9lmRHpdWUAGKmzQPqDSrKwfbZRnToifq/
scdqXYagzIdZ4SFGgnY2+l97gngbYC76lLPn6U5xqoIEET/KtsoxXUqwiAxc/soa
gxW7Ki99ODwYsJ03qIbd1Za1SBdv2Jx6Xbv2NY3qb75tJ+bGat+jA5na4RsCdbfz
zTti7RHYsD6l8kwx39up9TWQEdVrpNlG5wGlYG2FmS4cEptYDSa7kYyxub+Qeg2w
0uHOqeVmLYYVjbZtOsmOc7mxhRwcMs7n0P5W12BNo4rG0l+FQVDevUCOxX1z9hxm
8ee+pJM6/9btq6B/Lw+RLSVDbodjWlaXMKxpqOoC+I8DFWN9cTOCiDtYYADa4VBL
XkJ4zmynysTJfR0VHLfdj3KtjUitvHuMiyNvbnOjZuYInrIcxgVQVeXTrAU1pfhq
TBNXVkK0cJIVx/+y71Avno/sjBhWajGyY78Mfnc1zYAbsf7aHDjgkia/oMt7yYjN
3RFN10jxliiih9W+LoXLvDLX2ygeokBrrTTNSkRDBycXg65/O2QQkoUCRNbsa7qj
tsytAkU1N6IeyOaO7/yqz9x0TFgoJ5l/sfcvRPj+VsD85S+zHbfW2DEQXCbPrBkG
iEjbOkcNDOGcAzqDBDbZIOem72JT0WM9pPCz96l4N9bqHbjlxCMfvsEJB+boPF5N
71UB9h1uYQq7C2KYM9qZre48vE0JoNkOfrcSj5sCxDowmzTGrtVJrfTj+JpxsoCq
runx+8rY3hkHHoCttFEJiKfsQ0qUIQAL0b7K7d60GbDAn8a1eD/HbcDljUuCEs0l
EHuxwlLeTSozvNGv0+fv8F5DiJAi60/TjEdd10VFA/VRteKMyxDYVZaXVA4C9g7M
vq9mT5oNDr02BAUPEyvC702Zt3eLM7Wk28hson2kgFNc5yvxn3TX8+vrSFNl0gJS
49j/PC+1j5CqNx3f4Ot17YPhDxvQsWcLSuiD0Wn5pfT8mlg37vSoAtRiuhvgbeSV
n7GbOOfg/FTZqmCJf7z6+rWLOFd6TuTdwFrJe2+gc7K/9lfh1cZnmOZTlE3thnWV
ndv3FHbCmBLidLSl8GjMmdL2IfmESZXo1EnKBgG/ibr7VOwFzO+QJKqEdj0eAx7A
LfPuZE0UzO6gUUmQdhuX3ObMuUfkePZHhKz5WI9JD7SkeIimYH9O5Fa23bkKfKRb
V3vBGcZRkfhDBWe1xZakP0NRi7kbgNNt1ZfkEjXs2h69y+nv3IHqiNjQpkjhwHzU
se/laRHGFxEmy4EpWrRyNl57FINXZA1YfG39El7Cijbxdv2LxKQ3XALJh3SLVb5j
3dCnFGrpKEXGceI/ekirwluspnMIg3GgYCZyOvIDMQkf5LnlyzWst6WEgGqDa42Q
bkqsNfOJrloAhbc9FyYM8/32UmzKv8fsTG3FlUAGkaF+ySclrNk+Fo6p7v0zxVPn
uFzh7TrfWO10lwQqIa6NMLRFvNTveHW4zfZhJnHZ7QVMm+3FPITj+ehzIkIKI3ud
LFLYpC5Zr0/yHE+VneY+Y/29zi4Ccf691gggGdiJqfaxpyQawZFnkIik9qSLTNc0
7rMlJ9WSMrdjW7hbjQwxv2uYHfUZw/zMZZiYbehyBTCdQS0vHKhixP2jH7oqOYVE
hMGBbU9p1WDud/VPyVZokNL5j3Ms9owNaJ+RL6jfUjQDtDByZWJwGZ+kb53jMtnc
S3QMxrGoys+cWMoP7aJakniFYrRxKRbMl+5XSQ73RUy2ByQm2VlRNPzClrL3FCBN
pLXq0NLB/CEobiE//YNiHhWKipAYKelZ81NgJU/XBKTWgov0ZBlcDML/1Qk1Veod
yxnuos9YGpdTJavcVHpeWw22XFke2WrnVa2pA4z2ExO/KJ4Cbw2TjfFNPDEpvWMb
NhguNr6nPsX40/LL5dpR7EeI5Ymzsxt+b6Yelmao49rI6dIszHGA76BHcZXknuvi
8TZO+VoEEjEAXxEKdKE/zaVWx43XWbjHy3LE1EIl+J7Z8gLcb6RSRPs3GCGj4EWp
9AH2PSJHxvNY/nhslsAvqwGDd6Mn+8cWkVQDcJJtLWZnUR+gsGc1wRg02kxwc0CN
/ekHFQ1fk3Eaea5meTiC1+5rg+ueol8Idm0Jmt2l73PsQ3BXa0R3zItS5VmRd5vR
+Y9V4qc0kJ+21xLZWWxbrXQgFzVBlgcY++sNK8ZG+svxWEghA+rrow3Ey5Ft0TYT
QRAF6FPn3y8uxFhCxHLg/kPga9+lBWWL2t04ODIi9+eguqAhI9uaksGhiN8+C6kz
NW24rgoclpawTymJj0kJfQGJ05o8uQRN6Bd8DDtmRwPKgUdc+zw6FcShAzE1sCLS
5YyNvTHBNJlFxCnY2VxOZxLI/ieXwevjN4/8czXoiY3+XlsXtxn69NNR2Eei27Ca
40ua0VWp8EcA1qdc4XF4tLMtVh+GPkqnTxNr/ptD4LAieCW/Bz2RFH8jdjWwRPK8
QTSEDUVdqz9neSoWJiXoS/yj/QC9yL4hkd5rw5zdScfmgYM11g35tsZiCloQFnbc
NrHT+GDj9xbTXlseX6XVBoDupmWSRR7dAR3A2nGelFv4iYwNEBxJFyTkHChio2B4
1wgSfka4ftT2d4nn8oGJGja0UIgwWy7W1qVEzF92z/s71Gs42s4RRP+ldOJoxheD
9nEdqfFLweh2h95iAutRxB32iG69VHaZMvsBfFZh1UT8clH76nWN1KV/Lfg/HPLy
rEahIla08IZSVBFmzoqS8SoX+LGYRlFVYTQT5dnrnl0mUrnu4Jnt8NidyClcb6Rb
QSA3SlqCbTTfJJAboqqimNFWLf8L/FdM2zFSzsoKwfEZ7wy0wLf+km5Vz0GYbWP9
D2cQKmI0+2UfCxyrQuQGx25ekRmpPNvk8zrvYeqEUCZSCbsGJCXi9TxJJF3u0z9E
+9RtVTVyeNDcWDRgNIHoRMxU7nIgm1etx+QBqkD8V3PngCUnK7F9+exuyfm0jrIi
CAQeY1cQxan5cDDNL162pvdYpO2JfxL8CDfZb1xY2RWL2xwuh1oZHJJt+T55Cn1c
zQaztSwhmEvc10Dp91Zgcbf/Y0H7Vah3zduVPkief4W+oxA7WsSP63kFpD8JIXtv
juaUGQKHjQQ/lfRFZYQgYhphe7i2xpSmsCoI6lOeM51u7NLWLlEwQXjIXXXvPSOv
bh7n5VRWomzVrw93kkH56+guPyklInwQkJRKZZQPw/reff0Kf39//PSoiMcKcyzg
+/dfcfScDTad+vwjR21NhnVJpjOU6efq/1TaylahLszwinLZ84Lxx7ikvGWaQl/y
DyDWQtckFTktvacElGjHnNMwpe9rlF+EIFtXFg9HcvxS8vSo3eqwiv73iH5FBTWS
IWIu1x3+j1NdynJPV09/nd2KRghfxRo0siNqGaj8oC/4b2Q8N1GhdFOPkDteDo52
6JnLwaa/ZF3j7BoCDsm/nAQ0AMK1wnaPCqO8gL0vayk91r6JJqSJvrIed56n+1CG
HslLE5JBkLzrNwZ02KwOp/5EtxkcUAFYbq3EDP+6JUV9v/IfyOOk+i012535G2Tp
R0xIYvj7W1LYhIhgnTXj/YkNfK689wit3fN7UmVzKD94EVKrohu0IDIqUs6HJljF
JrqLH0Wn9YW6BLgD0yXOrkRTFvAd4w0xsrynnLCwpRnJJcJu9CJQWeAo1RrDI/1y
h3hWxUOf15eojPy3/AmdIgUBY8r5DRIY2rz5kxyHbkkBmcpupO29xLuyvWeR4WhL
rAgmvH28r2iiN9tVQ5tGufGKBteJ6BUZcmHvQz7RSH+oK3oDbrHVICVsXcZoQJOO
ul26W5aDEiemlAC5O69mMrfX4QrNJ1o1p0H9aJAUJrc4IlPi2Gf1SjTc/Nt/Xj8h
7tZhLcGAIB3RChq5oeKxFQo+tSiLBT9aazkso+rJL9pJ+3v2UBqL9rwtQF+3DGPT
1sVrwhjCROK9FClfg0KUPRoqMnSgh25o0gorNVJhz2dS+ZWVIv7lNYoAyPjbiZaT
n/dDN+rxoeqZHR9wBS5K7cXo4BHXLyzTs2Gvdp1dbIRX04VS31awHBgV1tizDiPW
vZyKW4MzIaHnNVwjqhJLsA/ecazSXT4ZaXL7u6f5Edy67vyBjAbf8h4o0EPK5m5M
8jRG17X6iG9nJ68kt4nRojPGhH4ERozRkjlzXcJWIEiIKX3epl0WEC3jN9Hd4XfJ
O8KzHyWz/Er/c1vrE5LFJlXTxv6v7WjCKb8egLC26HWELPUK3KyVBmez+DaFRhoC
gWTk2pfAy82K/PwrjAMhH9PRcKEcEa3fda5yZtY9Wnbj5xcI7m6+d2yqk+KfWFgf
cBXaEK0jC9ZDiOfDlYw0t2WWu9OX/eOhxNvZJAn/Q2ciZA1RrbK002lwLKsFrKS2
pZbuJC464GGKhf1f8AzkoHaK3gh+XNquYkj9Ig3h+iym1SztQk5TV1OXHeGOGOtT
c+dEH7WTnlFqMYqE0dWc1Vu4gRQKddZ0E4LteHQpwQoqUTRDotHgVXSiLsj3QmDF
y8yFHgvSFKcXNr8w7ALb7d5si+jvJKGuMR+6xUZDK1tg4v3n7C6PlArGyLV+ctTb
HDagk08Xf2X1z0qiknfOAsN6TNBHsp3t8IN3ZPLQybI6GqPt00k60hGxh7ZA1zwV
o87e2nQhFS0Gyh0jzgiz3YrE6332SQ9QsB96/927j7ZA5Z6n4LyQnXepIqUDrEsY
nPTj38OIFO9a7cdkE5xx3KmhhEwwEaIVkqDtp1LzCl4RjULoUjBuZzNVXSaAew7+
kqRxvDJSvErOO7NK/4uPou/Jb+N0Jni1iKpBQ4vBmgnD9C01Ll4RpXa88eesG+M6
vEQ5Th6ud2cCs3KSUI53iWZ9S0Hg1zX8b8kolI/NRhJGBpvw43AEDQ8/R6reXu1i
1meMtCSTQ4TqK9PFXE/DZzcqpQo+XkH/t7KdD+fmNi2krzyBW0Kv3vac5GcgbeYB
1DA4XXk7uBoTtmB7Czgv8SC59pbT3WOIDoBjX/3jphKWKr/fUHrN7f8zAtXZ3Yft
NeOU+VpiuLR2IOq7lFDa/B3eUf8WfpA/NPP3cFpchCq0ZDur57z3oTgSVUDegHrO
YowMUtjNZhMnY7VtQKpzwIfsTc8d9s4vwugrW8WXfXtI2swWsQxdfzZrAR3az/uk
a8lpxbgBkkY3F1FhGVRYXw39jiz+JnvH5251nj7p0ame0/yoDGobrkucCsQydUzu
GGYPHFxNgU+wEQFWtpOypTDvw/+8C9ZEViLUIOSIP8tu42WnmFgp5vvs+Fj28DtL
CoPNKUqwzlitb2aIrX9t0zNPI96hq3IQ/vtux+vQO/XdZAI73uEJYlalVaZTnr0o
Iej9nW+NfH1p/I9OeCXX2HTlCQY20g+j+aJMabtyX9wcIhNT6CovyWlJzuFdvhvu
icFuFt8W5XmwNQrJRzQCkZKDjISJSuBKe/m+NBX3ZjmZSEbAWE3o0HNwf4ViuI2e
ecCR3PllYflWjdgTo82CMUjfXVk8DyVWvn9tvcINlSKMBp2++04P9atKR8FrA1az
LIGHkACK/DEnZPnnXRrY/dwoWQlgDDqyhFULNwNcfs3GERf1u+B6UolH1nId7S1D
TlGn3mFl45WF5zkqLgGnOpcYnwJNE7ijAslXJR/WEXIbVrfwGyUA8hjUkd21CCCu
okrEhtty4KpiP4BBsZ5VgJmufm2n5iuXScOP/LbOab5M3bav1LpAZfbvXZr3m/CD
pJFCQSNWPPPxzF0RcG68PQp5OJUQoyNcrX2sRyGUk4M7ZNwX18JKeE78cVRIwr4W
mehZ+Kp5hJBre+VWBjKmOge+ntfhcNINAxl+Cj9MgS8HB2bHqG4Q4WO/XgutSQd5
91Xz0TS112iSkkehFICO4b0UqMCVYdFsyRBQdD1CTZJkQzYYxy5i319FCp3eK2Da
T02hHQk1SfoFCeB1GyzvneA6TjxkbRHXmRKpZx2dJk6KVjyB8vCQOMM5sDx9hIJm
fQrF8AT3Z6Hc2vgUefj63F898zu/lMg1PPXg8gSIEIGpTxBo5JPaGeAJ0ObzP31I
CpV1JczqL+JEClwp4oB80A6Z2ftS62rN4ye3AMAZ9irTVFV/6S1i/mzQDgar44e8
gGH48cH0M446aPpD/PjGr1k4+5wQprSAUtLm+vrE7fDaz/lYkDyfYuutIrBMZH4c
jvVK5kEPylm85St8Ei87LtxFhxftYN6Zw9fV7Ei4+VRO8zmVQGtnwP2TlcvVh/R8
NdcwR/CQzEKYCtRvWiZHKcFHGrkdpCN8QV9sN07pWqEvbwsZhVb6DRl3d7y+s6oY
PB+xIJsGkeEeuR4GdAVOeiGu951FzAsi2sZtVEuUKYUwPVJ9Hu9LUiG2xvzIF415
CEBy80IY/u5zZzIxjlHOkkwET/GvtE77kWaTnaFYgZJwE/eL8fW9T8eQ7cux/TqQ
WGZBrKHjh3joGJF9UUyLeJcUO6R7gdVTf0VzZwImeGRPqNff82r9ogJKJQHee2AH
6cX6oT05lCQ03zVgUI1Aksu2cdQ6HW8FSK2FQlhRt/DyKdqoKMQpZn+xXTp1Gcx9
vUcRPDt+yj1KA1oZhQyiAs6k6oLWgtk7yjFln1vpKQKNZHSp6npq5nuNrkR3doiy
xqfDZZuEq5cV5CI9Ww6bAII7+NsU1cC6qjeFByOt5US3z1taNhhW4h3otSEJwkgS
1H4ctobU8N5O+VAXJmdFGzuVjpY6H7jCkWqiy86b5uMnC7Udx775nqbR5wtf3LNe
fmkPmtERWfUkk6pgmyUO6S0oExYBkgrFlhrz4bBUJ9i3RctD8A3JSwRWFXEmOR3Q
O5PmUrU/2I95KdZevGLTvpXAjkyRHBpK7YIOto8VKEM8HioK80d91lRGkBel0TCB
FmGw7NjFrR/Ly6qMxsnwQyQ+gicPtbUJ4dBU7TUVqOtGTVuuKKvyeQjLL7jxPCr5
VsaqhKBEo4uYl/pIqnnmsmaB2olHaAdY8eNwDfy8zXhGge8/N/rSN1TFNp8tphdy
zdoP7l9zahI8tRHeG4oQuf4MWz+5aaY8sbG+ziCgtIdYKyJgzgIIMhPRII1mRZX3
Cpe9qZpQ2Lz1jQjrECRhucQFm4HJe878rabEQl3H8DCrXVRmy5zNgR7jTWRRy1MU
tP92xDkbFFvvF332+xxVppPOln+cBQJEFnnj+FO3ZTl5DzNTFyMjVpwpMne0/2Oi
pCXKUCkDlLQAlPOVv8O/FuHeCHHxa+jBQ3fRhkXcTh/3af9auJE9vMuxtX0Jnrd6
wQ0+k1y6h6YxkDFOWNyeEHBw9WKHIOU9f5iKvfL8xEEFh/B9WQRAmsjIzaIJD5ly
MzEKqXf6imKJUZtWCJOYtS8Xi7dNUFxpGMf4clCVh49oJWahN1zlCnDUyBkKI35U
coG7So2nNnOwhi3ibDUsc/KGveUnHZ2bVNjlV/x8IHCijp2YdU2/iNq7ylEL6sAS
YACBlSIr/BCOXmuFCzyr1cAP4zwid/li+lQbcy6dcfaADhRQsP3W+ZiSB+IPwFXY
EFhNqwv18Aosq9lASFH4Ei72vGozAWnWdqsGwT8/LwEwJjT+B4VMphJ2R0hCOICk
yt8sZXlMWfiv5pptgnNwNPv8qUCp2wcdMrVXoag7Ij6kKvL/GJEpsMCzNpmuf/yA
R/091f3jcdJVu2ekjf1wztQ9Zrl73xl2dL6+xzQVz5Y1ewjSa+BMOif1NNS4ZH2L
8O9KlpiBSdRlCt/YcRBr7hXumExVHQV2SvLExQokJ28lP1j7ib+VpAeRDEOpD/Md
0XIafy6UOXBr+9hxFSzUTIsgMDTPWZnvVSf1Aj1HePVmkyIXicaoy3ifEUXzhtTy
+Ox9TfpMxjyH8UGGgq2SSlRMRh0Drv27ulADL/1P2JfD3mo6HsIhiJElTBJGf0G4
RASuSVmDZ7Ue1HKcT1K3QjyPIJwCpBSydROOiO8tDUbeYOQcSePtf8mVh4KgpL99
tfUs/KUJpPMwbVXdgviM1+o91vwRH7L6kmeHOnqN/Q09dFUgi1zRtQIlol1tFCwW
2wNsPMrFMPkubgAsiYkC+fXNRwrCU28pq3pt1SAczF9FzqDZ5caJzwYyWjN9pNcw
GohdEVxDKgjHjv2zd8iMEafFVzAndHESac5toDYpli7NVM6bZtlVdQoboPFbLwo7
YHo1ag0yhtlvIdPvF1zDovlZE20ftIkKUTFC5opaz5CAB7QUlzxbG7dpbKAbOc7V
JgJCE7Ei/ap/uqyjfFgZoYh5BQ1EPPEuF5Dmy6KiI8O99v/jqKq7bBG3sYSkE7hS
VA0oVEhHc1MogD8AhxVzY6+ZxTbTqDblCi/LAmbZfJ8Vvrf9KpWdbvVfvNfXcJRw
iHTq0hpDvb/g614JmnSTxDXSXW7WI/4t53Mnoa7J3k8D5vqlply32cjbkK+/pVg3
iGtC8yOu5OaVF9BKStisk/KSLAngcKu8kfeY9HstA6YgmWxbEl/s+H4X28UrphNj
SFOqaQ6QYN5oVfK8oQQfDq9CUMtIkGj5+5yCJ9+WSSklIeYXSJ80q4y7mvetulQc
i92AxvmeBaB44qkOKzt5P4jwTY3XJM/ePJa6nqYnoQM1o6WRPL5NgHPk8H87mzEE
CvGW9SenubISvNW3GnoMcqATLTUmVZHnG3TLdsVmMBaQ9oDh5QtNTtA6EyC20Afq
xPfdvTzQkrvwei+3U3EZBF3jShfN9SRd2aq7U8pSQX+PWPZG+gFbq6bKoWQBnt5z
BtL3iIrs91fyi4/Qr63IvDLtsvRH1m6/tLAyad5h72ld8IzzpmLW3emwoKihGJuQ
IpCIJAdjcfB7ARFY6ZsLMq4vUkPGW7ZAmWQEhfHJ+prSzLNONst8bYW8R+XjJUxa
eDuMAmelmHOCpEbYqI52GjgNESfsQAANKKDMYZtFwZlrzVcky3Gx7etOVoufT1R0
iD2dGs0UcjfIlsFKBsQuSx90e+2CcQRq6MvOKWS84y3ujB/RSy/6cZKAY7DUXHEe
rbIQCYDETALeMzXor9WAXHd73ipLuQotIlZmAAiB7nW5OAKgDtlpNfcqu/LJmGdC
d0+DDl9P4Hf2Xfzwlgnuc6YWXgjgxhAuwv1FaSMshWpzxD2CPHnk+2rtBiJwKWq5
0mUNGSqytJHyGd98A+amPcWhhCVNbI8ZvQ08X8eZyLf79XY3sg1owug8PCtkrUBG
93MmORc5XUPN3Nwi5CI+VoVSnfnS+XL+VQRvoSdAgdOQNSt0Klbb7nXRivvFma4e
VnkfkClL51J8U7iJ1VCG4Zvu4sEzCrbMHOHBlCGewzDWtlXTW28ZsjrdGh+p3rOo
5zBzqQUfNAuFyw0u0wgFM9GsRdjCVP2bDk1JVGh9tOYcL4GgWVzo/lki12qfGK03
+S5zFLs/OGCCe1H1TXhRQFzHRv8fkfw9E7hmCLqH7VAt3NUQ97ekKL+Jlc9lOMbm
NIDEoXCcUEnyPqcIhus6lkkfWsqUo5BvvvcB9ZOjiZWQk8eAYSNrrpWhhbjiHjEO
HRaJYF77inFAuFIIhtjE2QmOXXyYC49plEsCk4+3rMCvzhSRSQSEkAp71T+Yy5yw
I/svg+yKcN7+Yd+Nk9ZLLFVNznR5MU7OG72Z44nGZc02TZhX6qt2tSmJczt0rKtK
KjjBV82uToL6gMP0eDQlP6P72VUWFNrSD6bn+GiFM3c8RAkgsEXAnMMnO+mV04az
6p4c8tmWod4ydSRt8FhlYkokx3LaHRRWto6H1ixvqaX8gJkYc9IWXxu7D781UJv1
S5SsMqBD74APGhzwyeOvA92cSSkb/hOKP4//wzJsDi+MbnPUnU01admTlYss9a5G
LL53lKYIBmsQdi3Q+O3UJWPiKQ/exk1oXUGBfCkq+lPKyzX0OrdLc44Lp1TcuC6v
vs6eJ5C+IRozF2ATY7nT4EJjDB5ccpNKoecEG7yHxCqo9y4rin07X4LCFg5dkG3g
8x+2mGQJYDkfSm3rynJP7Pg7GkS5RJ21hZ8A4I30q+DNYsHU533I6Q+k/AVPXxeU
s2MvktAr25XU32qdobthPzU1Bg/JOmfL+tAulP11iYMm7IaJnnYnmjFtlaEf8okC
2/w0lUamBNd989AZ2ynddKvioGSIL0ABKWKxyELtk1wg8qCYnP1FzknuzybyV4rC
afMVt/MVyKZenCRncVL/iaIx21EhstU5q0gL1Z6zcj0QCzGx49+FbmcjeQWA/2Y4
SNFbTNmrMT4FUnbbm/v5oTCVlvVfO6psRYsm76fcFie+y3cEv5AfdyW5wBKgU5a7
X7aGbIgk9QSEBU3CymcIRQnL9/0X4X8BVCJRoyTUyZGPU5BIuGAxS7vHkeZx3xUw
MHBKPPXONxGwCBvMzVLkWudJZUxGjYsh6pg4YWi21KLPaNKgaot/yobsUIKo5IbF
JUof140TLvgtufr1YC4TOTfYny2i7r1KSsslVj+mi5OBV2zxoy3dXs6u0C47OxTM
QmfpGsAqZyWczAOe3N5xCy3wfuvORv5+n1ftA0p58stis6QQs4qFjzPbDfkc99lh
lRaqto2mMDEiBLug82nt1ih4BsX9UP8a4E6Bp/+fpwHR65dFZcVHkA5sv5gLqhaU
V9aioJ2cXSAiIIBDb0y9HIH1hJIHQ+qMEV+/WwKMt3pf2CseL3QwjcMHkT+YLhOL
MghLQqJvZVBZn2UHdN5mmB7ZG62xjbvW7yQFjdwWpAbGQ/oH6EEiju4tUoip2Nmu
Qtl/YybJ2Fxr2njEF0Igl8zmbnKcPT3xD2dzoRgLdygXOfVkBcgQEuSZbvjWgOOP
hR2VgfdQfbM5sJ6jHdMT0qCSyt5z4T0AEhxvoup7nwn/UOn71g+YfuCli5qtnvm7
iAKQe/TEzzTU0FIGg84WW03K/iexAljAjKbUj2m1KmJhDQaTdTObzXQDQn7kHGNl
0TvYh7V0Oi0aEWS4YIYkGm5Y7bgSGrrXWGFgZOGcwNUnN8L5a/BF+XRAQOEGuYpO
Q0BpI6pH+wA2D/tVRx6ZAFnzZanG901Wz+ol8ToZaldoBwRyuKyQX+o1k64GCSIM
pB1ygOQWBtIag+qHfQYpliuVu7ldU9TU3Rm9hEqoZFLNZO709MEvyMDUjnf/ZJ1b
rPIJin11ZJKOdwcAq+YQXDhAMiTRlByUJ96BVDIuZ0OSU2Y6LJwdhdtMh9veoAcU
rhIfwGNWQOTIZgcYa7OcB/xo/hqegWbsDBYkPCMRvuS3vqWLdKr8/2uNnmo7W15p
e+Wx9fsE0l/vUntbMs4Zf9nN5MagfA8bEMrUsz/uBvnKpnVdBnojBv37tBNBdQS5
GJwPH04KTpli2FHV8dkHycnfcjrcSZUUPg9N1PIHJ2t9BevDn+87FO3NSS//H349
TY2uvi45wXSRrSxmCrDa47cUxBMdbnaR4XmXpU0Bl37COfcpPtDppejqMIIJWNW1
p4C66J3lbB4Mfxp5YxSlywj6XdJiIp4zaKqgPj1wlzk+CGFIkX3lqybhs3u8CPzS
XvizJCqsfLYWsr/unnEqOEpRlMHclBp0vGxZMrfJuFmKc6HSb3CN+PhU9y+KHBrH
7xKKzLZv5Y557im70fRXZRWUo26vzFQJgkJskey/d788owx+jPGW5wcUP1b9OoA8
9PWMTCJxpxp8fIHq58Hc6rkHlCwwWAzjluzaufn0Tk5HLuOhuHiJT30gMF2k8Y5e
n3YRQI94umoPs+nb0NmTDleBtifJjB1VqaUcIKVIAArKmFvGL8c1KxatjvYFCYun
QCWCwoyp8QuG1Lf2RsVHnMadMqMUC2FYrQNVDnP5T5BhwXJr3H6FcYCNo9+INPin
DOCMfpIWmXU4tty1zjPj+wluo18UKIbcsAF3oKElbFHGDDfeSsVj9+LhnY6Wydfr
aWAoE1XLYBhW5aFZ1Yfa85tarLtQry5vGLC2Ym2LHXQq53Ix09jLnhk4DlcbUKsm
ZVnGt/VeYfEbLUffW7EPzDHNt/Ejt1Sfpg7Mug1JXMeFLbH565XrBE0c3+tRn+C2
TasqbBc6emvqVJkIsoLuJu69yc/vGgYHM+8TaKg9U+AgnodQP+Ovt5ga1uCU66hc
8UwcYL22XC/Fk6x7MfmyiL4lDsUdkOX6BTNag3hhTLVih4OqrLgDVggaPlCpfE1y
0v9z2W47vStYC2KyMtBfe5ilB285oVNCsriDdJ66mvm6cU4wPfcqfwuLQhf3cpyW
uROrRRNvNqatGpwV2UKj5A/nAnm+zV8gztRlCu7N+BjFhcm5HGd1A5OxekY5RlhG
GJ06ZATdWISw6I5gpufm0szcudIDxzFurssmEnohU9LtJLPKJ39shlnOB70qhXPD
aY6I/YMtZDAuCIVK0aaPeXkx6AoTCoJLN7hGJVvNrB0PlLZWyCJg4iIPvIm2/ytu
xf2oYY8GpLoAr/MdWnUyzTbfUUlyKH4IJtwZTPR1Y4MJGERM9FgVsPnhdExotVBu
IjCCPDZ44A167ImXz7WctdsToaXTItFr1a20ozPRKq0kpKj35zXfFvc7h31oTDuv
AbTiulzHAongXlvoVzjrxLrImWPENwtMUbRjIeCEEg4+X+j/E2/qOBPR+3biHeDb
ukFxbMaGmYLnlVJhFPCa690Art2QTuIvNtpBMXKfPeit+bF4bObChAdJLZqLcP62
ZB8+4hI1WFCikD7/2xlXUm0kyJnIe2xaCr0bbqeGWtKlNX7/lgLdj+rTWCgNTbg3
WWvMNBxbaNMbFxzi1HgmH3aoH9Fcmi04yFfiZchRp4OkkndLYUEzdpzzgd62BqGz
p1BHE4oCZNMnBKnYSs0GsdcI4+IhKU5PWqXhqjlkqNUnRllzSBmluma6tfs+TXq5
4g2kntWFy4khfg/0KBRUESwtuZyK9bFl7FFzFOba76yuNcnHpDOG/80fhz5BavE3
DM6CqT8IBbRojL0cIG51Dl7fYZtUfHzQtO0GFwTFlJOGTb4AW7tviu1ToZ96Wk/5
esSWc1nIoyS1MNNu/ZRD77WpW7VlSn/aIkKmaxCCB64WdEKA0ylaAT92RU1Vpd7Q
/h45si84SZOYRCSXoM83MsbKa1X6WIOkdtLaPaWSEjfE5OuzsC2ogPqhfN9goSKf
w6ngwvItlbCLLHkNkZD4PQ3hS8XqPnNzKANLtK/3diKSQYtP9xdB+DxncBKR6CmW
Ajd4sY9ws2kCSU6C2Zy3Yp8Bg2pBXCoUsyeHcbltRpffYCqRGaXx4KRbCneTYPUR
VZR3eM58I7tiMlczoTUS287Cx6VFsj5y/xu/bMlboWDqNDge0KMYixO/IuDREACf
cmqk+oxjeUC3C/Wvd2xK7GA8kvig7lfTuSdxLHFC+Te4iJyoDde8dObd99UHiLOn
xYAPcGnB/5hmL8g2jMwYRfI0r9rQe6k54oTcRZcG3Sq9KIdxYjTPvtTR1fpbgFJH
XtzRuZqxvbBg8iWVZtOXA5aGk9W52h/6h6pbihQtVlcPRNLRyvu5LT8JPzZW7uIA
fharhAt9/etfYNRi5U/5uq/jQdkp+EdqAoHqkz+bEqmHqrUyM41D5wOTKppwZFtf
FP+wNUV7KS2VqTseS8KiW03BsSI9lyYvxmrtH0MMotDkMMD90LCsMk7kHNvM3vMm
+e6xaGKhDZzgfxJt/U+HgwRaoqNLKmQQiBpUkz7Anj04mScK9pqv7+bJMtRKz6no
kcDJ2rOu+9mpZU0QdwBj3zYuFfXzhOVa2OBsbhWrNi3GGS7Vq0C40JDM4Xn6d2YF
yFMJozAvF/8qVOVf2oOktfyrX3gKW/uv2GlAJj/I2Nq3g/8zyUKVy74pavfPOaVX
qpfqLQLLA3ySQHYR2vLTfAXA8tF8eXafqF/6hrdyeNTJdZxNPNaU6HgDO4Z+opLG
63JnUrYcnECFH3SrpyDFybDK+yJ3Dz83Mu8KZ+NrXNoXf3mCgu6xpaCBXmc3pYR0
FttJ7WCknOoLf8ETrcK7mWLBBBACUdey2U78OEDO/xaugC1wj7WNy8F6IHFeU/xE
vzw8Zbm4Lj/InBsAVRoyYzxWzGiV3Dgrd0GlY1XXLZ7xPpbUBYQTeHj1GvG8luss
baUL6EhL74P4hwzmYrST73KHWCJkdcYVFN26tWrRnKr+71cK2f+3lAaSLk4UVIN7
4GpHYFAFJqYqV0gDy61rmDlhTxpjeWNPPjB0zTpr0c4g7tI0dL+YP0pao9fEbPxC
f4XfcXTi2uar8tdcuUsWEz0hHwwe8LC5vBbPh6o5/KgEnexzaShjeCkz2qEcXbx0
gmfxwF4c745gqBgeb3Mj/DCdD6tdozeRFGbXyZdpA4UZEoapaIchs+nVQY1o/21m
DEdH37AAe3qv1+WReXlGmN0oOduGMK92IfBjQTxvE3sixdFY1ImBNBTXsjENH5sG
Tc8BGpofda+o3VvnhR36n+iHhS4/oYZ32vZrxtuu2apw1a6MVESfZB0pmIEdT9Sj
SLM/Y7PB1Zs65V6/M/tzPkPNTZTdyz0M8+MlSPDGQF13zEdt7cfmC0ozXxVfoe4a
P7YhZw89totWKdCV3yjnZREVlqtoyTo68naL5oUTcxkEo1c2sx3jB/LjHDHhcSSf
np39qAWXs+f6YlJxQb7GXkBnNzWWUANGAoori70F10n6bfNQVGas0qbLq7bhDuHb
LKYyURpW0bDRVPF25BXcYko7IoS4KUIQnoFmbMg9s+rs9WyMP56YaM8uSCo5XmEK
pZOq8yuEF4eDZg+42ixOv6jNOwO/OnAUQ+ZmXU4r5OB/YfAd88ZyfGeH2Tt5IvwM
K9MASsoAwm0kLMpsvVrMbSglETh60yL4kYywmW2TQQCQMLpIDqiYwGigwTwTFV/6
Cy8I4SHsyfPPS9L9T2usS5lCr0ma1KN4Mm7G57FICU6S1o/Mci1odMdxyGXzfdJ7
gFv0MCFWFL4gdex4rHZJItKDgqHrvq5dy3toQ4dzh/iATtQy8aMdnIGYWdFxSLxH
Wh38nkcY/V788rQVB+hb3YNgFrNGPlP5w9Z+VEtd0vR9CvN+zevzDB+JY0Fa6vUC
Q2R0R+EDHo8ClVEunL+OMgTXsKThuWAK9G1enjYCffofQ/sbuxJhO5blkyPl+Kh/
eSmKdmsUO75FuEcdyRVE/9h2AaJ1GtbZN7kR9GcR0jwzRIi8riyh4HnA6BDaXRSK
dBS4t8n4iJ/eNRyc47g2l3xNc1gEcD4Qxrf3Jg/NDXoQV0VqCC/UJOLoTc0TN7Xm
w7r2FJQTSBohmRXC8+7SuCdqNyrPiu6TvoljBMI9P5mnuwScMvIH7QWgwTX3xAi1
dbIqEEQdnnvyGJOOPH8ZG8aizVYH5WhHSUMt88lEaL3xZjhDeczbrkW/T/fIRo1X
0AryaVVLOGBwTMBXkU1ihOhtJVQ0XvL06iIcEcR92olJanpJnMYyTR6Yuert3cbu
XohGF4guzCD8HYYVeqaHuKgJnMJ4sZ5zbCga0DQ12tKPtSaKq4YmfMFCfkA1hFrx
IpwrP2ru9NkKgzzBIVpLrBCQ6sZXNYOKOxp1CKUOEPAPjaGt2dmEpmP83M1ZMT9s
g0BM20gLTYoNRLYFV6m3nfc3xRvF7FKgiKRquNdpq0/KWgGjYtx5CD5mV3oCSCfS
LhjMHZAxOpKXOr0ImyBfe6hIkkt7AXlHd5M1vcAIO2jFkjLtFnrG3+oXE+3q+opt
3yo3fN/CvUI7aZvNojTDDnAI9wVDFGkikGT5iKMJMax1F/jng0YUCYVnqFiSZcs0
n5I3YojP3pm0CcNQ1hHRXScq79+l1jlQcCykjQ0TQXY+7mwQX0OR8rkw+3bosBK4
FqmPgBYZ3pvWQxR6DAutodcfSiIp6ya1HKu82uamDA8oH8Tua+xq/HvS0NWG3e7u
xjOmZU6MtwPiTiC4qU4DNp01RbXYZy7Fl2CmxKAdpWh842LRmXlGCkQYRiPpPZCH
KJVZzPSUrxtM8zSdMWDfS1RVLTrjdszJ3DFlX/me1qYzptTU6NDe+rPuCFgNLpKG
zIUrQkr+Gmqxq4vKHZM2Z03sR70wIiA+XCrBlHHPZfOfEL/QgseZv3N3TcPCeoaP
Xu4v1FbgmmMs2BQfMuWm5hzgqK+gjFg4h1OPRr42NRslhh7JEvNZ9U9YJOLFZY5v
Wa+jFhKx3O35jdeV5gEwOK2YtsHdSef2fgrCOVeNsrf1y5R9hQ00/WQ4GQY2UDG9
cOeBi4YoiN7AO/+gTij2v6AGJ3QDKoE5oitCpf63FhCFYkDE6Ccv/xZipJNrSwNN
8eV54e8qZMe4nGuKeVkISa5NPQYaEMwAQXt9h4x7iaXxJIXcP+SFbGXxoXWLO0FC
HUuveiTTfj8RFWrXeRFWUKjecZsKawVBCOc2/Lgx7973vv11rYxitDyMdeM3U6p8
pp46q7pq3mf3dSyWZMEd6d+x+Qmz+J0L8Fl0JUwMrn5ij1tAEx0ZptD7J5aVtOSb
B6LIkFe4a6WvpkeJI2DLVbDOpdmgQ7bCXmlvmJdU5JW+YcDH7+mfw4QAnLJClu8L
hbts/3wlLCxyTuX3wXABDd4qwFBX2BoSder2grHG5hYoyfz/RjWPAQex+89kr/9m
6F4xxSHOImHzIu5ViFvxx1Bno5c78njUtPoqz0FQq1by+MLU0c9RyKYbWAWO8DTi
TGewIJThxR9nfccb/GO9WsrRliETVuFg74KaU3rVgHwyTa6ntWgOornV2SdU6mvW
MTGdxCXBeTHMXbo4sPEG9rRe+44NVJ/S9qTYI3bbaEep/D+HlGm4qZ3al0QeVxCJ
OV2G9PA+vVS8m1lYl2bor+HO9YR7xs2Icbby/TIOTlE4ULpVvB1d3xELJGnShH3b
/V9oiRaa7mFTzJHbua6j7s5G7l8qmGE7H0l+7fgrTBDg5qdHGvaAxTkfkNMVu0ZY
fqKwGAzDNcRUcaOMrUbcF+8EGaWL2i5b6mNd9ah33bUwLIvHBqg7hxe9byviJ9mK
NHXMOU6Ub4nmk5F/c+cin1xyeXv+1D2U9ohQNDqvxsXsELb2Cv3+gvaj0dlP/EMR
pQFK9JYrNhYw2+cd9KGm/t11IrrhNykapyCv3UZysnJmVUqd9DPKUzYwSPFHwdCE
lHrvijY4o8KUgBfv+XJSHAyCD31iqjQkIRTALS6EEOijGUyHTymEnpzn+5tQrwrl
vDxW7gvjNdU+NEet6xbYyin2oPYKHoi6dkMBs6ti1fYPxOU05tAMLOul81C/ZJN1
yT1hZdT3WZakzVm6n6U0taoW6RgX2yG0EihZ14RXZXChEaRPi6URgW0hVTcLkZI3
XRm5nD/lPSIhquCUBixlEIJJdlGsdmFa/olZMIEpjsOHtyfxW0pHEUHle+0ITGgS
sGfAzf34n5md1UQGEtuNkxygu4up/Mhj/8NhnFpUe+zEVpgpjhpy1m+aBGGkDriM
auxUdnWpsRcJOqOA+57lj+1HkvHqrG8ieRZbIWS+RlQtKCSihwNYnUdZLGGeoMOo
jcpcjdrR8qJg59tmcKzNg4rjDnzhQZIXD7+LNO2PxO3pF0T7TYNXN6QVTlWRoKEY
fObknha1SpECBzJmphBjoHr+SEzLolTJcy4eqHecyfrzoGDEALbiDd/Cr9Nh8vW3
ob494kdTkNJ65zXP9ucjlkSnU/NzoglUq6m9oceNI+dlfiIgudl8gTBO6lW1oDgC
kCQPOlJvh5CBx+0AhlFKBPS10wehaPSGK5fPkHEJhKVrNqHoNAolDACG8Qr+PcbR
Ki8oQe2rdlq8imB6BPvo6emjw4GVp5yAiUHUz2VpIxTqAdMOZjCaC6kj+3oZgLZW
cfNlfFX+b4obiQaM6ipjn3L7mJR+01dMRQNbo4IBi3Ge8hBCW8KTx0WjPrbJDMry
aV4ehvrmRUfxMle485x8zohxoYn7iTZPQLysVrmYtRGQN9NDI7sD9dqP73NEaL3l
HmLXE4u7Gl4b6g+Etehx1wmlkrvN2quBjynZoi/ioLW5vicT883xEvWmGtLeFUX8
rWsmdb0s2Sy30ZBTFM2QWlzhm46IoCsNBupB0RNnB4/jpISZf5qd0e7aVHmuTMRV
/BWbjo7eiCgyVQWpPXAb6hq9UgtIQRcO3B885eJCCkqizqnlThe+7Qq7gxXv3c6s
3lXRpjHJCbX4hP18bk+Tl6McP8yclwW7JWH5ZS/IuQI4zOJBEJ5h7HyOdpsqtLNO
buiMvbkrfOQzL2rY3SlYrbjhsihWVKlDFCgws4GeWKKc20F91dPVv/rkcURh+r/3
nrDbOU1StfVUkQ5VXn79N+vIWYPCavr7kWNXQphQsJUaO4HWS4nrWYz3lSShxmtj
oxbsx6RJ2vieUDLjctKoPyBqLVCOGFbcd2SQyxhpNtVUrEmXrFSh3rFw+49fNMsI
Eert4DlWeCb7XQhftm2YtUJc4l0CH+KBmvhl8lQOzlzGQZ+PmDMJS96UoCX07Jrw
BQqKfKx+j/XQD1l+fIIr45CA0BODhNi+TKoqgcbjUzqTC6j498mTsPcTgxkaZR5l
NY5h7R6mU5uhFKv/qxQkaeRVo0iLNQfyTMieUsbGxGMtC5I2GviWtwH+jK+QS1q2
tzjQ7Z3W9JeTrw6Z11RdiyWG8Ilnu7E8ZB3NZPxk3VFgz7mokUM1WypddZ+CMz3a
Xn2rVJge56GOnLcw0/nOHhoSzWSw8HjC8CDpy75SFCW/SzC+7US2yDFIHw65RA68
MRqFJgXV/lDgclCKKBGE18JgFqYT5KFXjpeYMU42TGZDnpwIRna0dpgVr3LwgECU
Qc8hcC7Zr+e1VvFaol/7Ogw+8PKM8KerXmb+wR14OqMSu4fO71PBW5VcOurxxykI
6Uvnk0bCXv4Q8upIYtUm0Ya9/eWTkZ1UP/28TGPI+lIIdppi8wXVqFl5qBzluuC7
h0k3m7oLb8PnIz+LKOQqU6DgMTQYin9lex0B/FmkdXJ44vbrqlkY0SSFKp2Xu5eN
Jn0PSKKniNrlbZMgNtMD48wdsAPLKu6IZiUGTk02TfBfRHgAUOsFFdzna3uhAfY5
1JJIFpECeSS8CR66B1dofzVf2Kcjz4y4oH/6r2Hwaca1+R8zhD2SqDOoLlQDx4aK
7BUvU4JsCBDSkk+rufWFfHy5oVtEbe1HImJIGnFgfh2NUGfnF2JZr+0hY7HhcNwd
PcKqp4V2pdoV9w3wM6ntnzjha+WZghFctqx/56vo9HOOfefoFoSiokFGPfZAlMwP
g8Gb/A4rcXCCM/W6SfmKXXA/4nLY+snEUKk+oNas9/8QYPs+eWSIeXQlcN+0KYHY
nvIbj7jmbC0HQVZ+1JVdPpRQ9NBpXujjLZ54sy/i4sz/EnDBMRWIy83J96UkXUVn
ZsfOqZ5JYMgU3+ncUASOAdyfw95ueed0VKXJqcnsqmdjJGn84lwirk9WTOnnTI58
ZXAsWWet6OsMtZ8yfz0WDPjdzOR+2Cgl3gz1oMAdBMCeLX3AwQNhx+Ph+uYrw7TL
V+qKXLtVZNcKMacidChvYJUVkd9umuWPWp/SWe90AmzzeoUnFrxikqMVNeLVHMOp
BPJEzL7gZNo1UyRpoymprrqE49fuJcAxl1SlvmpaR3YdJG7Il9jGOATXSAI7GISJ
XcESZrTrF8Nn0DCCqBjobn8Ggo08P7QDgF+jl51rjbsfTgTQKdgmdjdGlaxOZkEh
Gdt9DBrb4hqRQpDsUkyv1zUW9C9gPq1qKGKwjH/5qE+xK24wAziw4ji8qEqM1sIl
JaC1s4moCLxpioQ6N8DqJPyd+y8CMeM4BhbiQEvSjROHN8fQqRJqBB169frzh2Xy
g2l+Zigfe/bUcfYTAjtbeZAL7v2zJIjPYXMRWxz94MrHffu96/LP6CxcDn6ksjG0
S+lCT/HottbXDbhU8W7mv4LceLoI2yZ8CahcjFxjG3bYZInLoyBwbKdvgtHxm7LG
sqGgN3OoPB6SzdyYIQSORG3NeNo/5j9wByqfmCV7oNY4zb0djftHQPwWFk+fzVtp
mEb/lyL7W/CweT6FLPmMxFwzjS+4N3iD8Nn5SgF83wR+B/HdmBEPU53BFDZhwunw
cCdw0jf4rydAYtzI/HeIUKyAEZxF25jHghOck5LmeomBS/e4iymCGhhJuU6h9Lun
h2vIPZe4RIbQNRMFfmDNeUljascYMvDICNbytUGEOM0bBk9VX7ElJIGMdXvThgHb
aWVEjwvVrBaTPqr4OMn5Z1jz0Lgt+Xwt/KKAKhlB+Ct5KwuZHB4mEPkD/Scs09Ll
aH+T8IeaL3oPLtmE/LiXI+BYyMM+t9hxfQddWKUc22Uh/3oRCXmhYl2ft9p1wRFa
38D9lo4iD2I9kTXGubHTWhKnAglp77pjyDWtk4WeppRGTp9npwTErB0iqBlM3wDR
QIZsdQI0a6hvqTjHOJlMiLttZCczB/GQCZe6z6fIWb1J2GwqHapcQyEdosYgl5RE
P31pzF1rj1MeVE5g4XNXUzB2wG0anxTd0lRbESMOlI971KxdEp66bNZExH4ygB2H
LNISxW6EJ49LtTVy6gMMg14nBufCSPIEOZIRQ0VWaPEN7lgWy/BLx/zVqjIWUmiy
I2+Gb40q/M3WFgwVqkuR2obJ49ChnwCU8wg+uzjJOOmLOjSqTbfL4Z0Tq1612TUY
lj7WT3XJZXh+qiwh3rzWGoVK6ZK+TMnLbM9OoGxcg9Vwinoz+fcjsrR19m0bf3FW
vAqjOxtnXzzkhFfhpRXwCf1HmZ/5Y+13Ups4/Q5xF9x0w2hmZzEe/DpZ3Oglz88y
c2+CTinF/KRgBknxLZALVUQ1xj3SSYzXlymzK5HVuECEkV4ArqwShosuQed44sGb
/aQxr/lOm5HP1FhpboR1Ekb5tlw05Q5Ax0A5PfQgNoQ+Eb5RJKx6nr+bcKyisY1o
UfZZLEV29/fXf6YQG9chTsqJcGYRTiy0cyk/vp0iTVWIyR5hC8OOAxVqwWCsaBWd
D0G++05FjrS6BClyfzxp1E7v+V2G0/3CgZJrZJc1sITxfHsYJYEHluTR3iqOeTPO
aTV0Sg9NoTDMYWf5tUYgt1QeF8p7Z86H/IXqwzooiq/gJQTLKiLtl4Z2UKOwx2om
lFZK4yRyj+1LbPyUATsdL2+iTVgGbHucjTrm1br915O29Zd+8rTH253xaVFluuYB
ZKZu+qe8vVnAzi2ObXxkHdWewBPUE7JP/yvlP3wAblvVeA1b2rYybmQ9J1CLOMte
zmcLH/4K3F+pQ5n3LyHg4rhgR5wUDGXJeQRosyL9COggYj3dHBy0sxExGeB8p29q
IbSa9xmRRJkuHGXtCK3Da6vAhQmYDFS+Dp+8ZPLj5+/AXMUm5YJ8uoD3jOEq2oom
ShctH+mDh4EsMiE4vxCQrkDBI92JeWsOdefgRfFSOR4sBmqZYuruED+GQhijzFVE
pKalmEvmhT4SnXrIJaQWB8bsIDksMPHSj5RhJuZUSZ81SfYKSJ1/fskgD3mfsX9o
2z6bSGLddMP9eaC9DseruoC1TsKOz95Wg3hS6+w2p7Qk6mw1ISLBb0UOLvriuN3f
1M8x8Oz3fMC27UJ7qTQak2aQqFrr6v4mCkeAcy3uC5Ck1nbJxzI/3G7XfHf2AgtL
WCqOAljCOanclygTxzzNbeguTv9up1d6Y5H+Rqbmut5XsILvOxgpFBw3Fwrqj+Zi
n4odzFhUV7Yml8Nol9aPnUBprHSWZZI2kqUoI6zRCE/4kd5clPmErrrWBjqF4JqH
WKIu508n+pJ9oihdPsVPTI6aXW8eYrmVfsoqietJ8+KHdkSTYBMUuJisGkI3l4ZY
DE1o4zSwbzDopFurZamE73Y4RBSQ4lrdkraUhfKmMbI5ZhnYCyy4C3iLRZ7K5Sm1
nLLt5O6HyUEDDMjtPvwoGSJbFuRPNIW/KvEuetE3kS7GehLISWCOcvM+lj7X+udD
Ixtp7Ow8mz1WCcZJtsIDzrUn58JLqXWZk4ahJznH1wAcLkpmI/X6gSpWtvPyaEdw
WtNt7fDgoobIzP8JK3oqBg1ibG9lyh3F2Zli29zzddUgEzPoI4CDbIdbz8RLNCNl
NGPqfrfn41zIQTgzhTgint6d3xQaoGr/RtfmnBCYslikbFOp1SwNYPmOVZR4hWPg
jw7NEr9soqm3IXX4ZV+fWqo2qvzEPFq7faHvjZTCLdK2MfVgikRZ+wDoJaY5MO/f
8J//SDwE4zXolEuI0oiYQmEqwYKGaezUmi/ct7VdSXlKY9UufaGPiYzgM1ZKtLXw
fKYQgkQC39IBBnX+o5nPKS4jOxNnsKqM/+zi2AsQoVd5cMj8vCoD7SyzBH/O8Nwi
StIkVPqupgZovLHyRa8Pj1WsCgnN7bS3zy6rr/3KbvQPynRpqZei2u+k3YUMGCr3
uKIEB2UbxoFUbIXIGynvo/IwA4SEoLBuMsfueskH1yBSy5brWGMu2e9mMQoXWYLK
U+BsCk/iEVX/EWKEFOZ0elgWBkWQg6uFpGTN4WdnVwm/erUdXMrUsPg/8ExIV05v
KpmjZROksnwMxUNnhdp4wSRVS2GJbR0A+IdvrV6LGZAmtyPR/kTkckwU0E1dOdjD
blQ1NZfKPp3BZHT+k8zEpYbpfyg/HZsG6nEErhBgAXIjzD4sAcPpMkH5Aoc3f5T1
S/nvfjzqcM7tEnEA8QdBv5oK48rhAkldOa11xiXOrBVas0wwvSjZgqUJbMnusFpZ
NW0L6FjmqleASjHCmh2YHFQbX+lIeMSlx1OANoXYzxf3+akbcv1Pni/i1lF7d+W3
bUa9rBnNKJRRo2vBRBM4DN72Z/m3Fyyd/fGSEeGmxKpDwj04VN9ETNR2o48WqagU
fzGi1nWULWyVWuvateuLADfLXxuw2DOAqxcS/DA6Ca+/dBff3HgA900mF4FyEcZP
4T9IE9edjtJZZQ4yAQpe+77Abiy8QGsUFjbRzrsknbN2RfIAmegDiht9QFvDuvsK
2b7307AoeJrqQjHuzQ966+neweHPpE8dg+Te60cHziHFP9SwOEa1/+BDKCmaivuj
VLEMYR4U5VM/ixFJ+yzr7j2v71lUkBSFf9rdUZUbKc5G6g1LeukRADku7jKKbujA
bxOM4YD41d1rvOQyT7bMdaNH1nckyvtkKPGJW80Et41VHcyjonnuv9mQV8b8O6xc
MXTMpYHBlZFFnME7dOCrKV2g7eazayJME/Yl3qp5KqzUTsTt44IjETMoOiKUBXQx
MrQGx8AesDdUqD48Wq++qCooX+eEUH1t8VKRXQLtNXNwoDH5++cM2XA2/gAg28/y
DobBHa10ckgMm839kCrhSP6UyUWnyPFWUVdpT+WkKaInVVBalx8Eo7wDLDuWArVO
/CmuM8OTNl6bi9siQWCQK0O/YiIeKhEB1gK7wT68CpO54qPCOq4843O4vbYfmSdY
kgQ4uTrzlmygnGA92Kz10JyJxQ9NOBf97WwV2E4bqc88qqt3L9ni6wJp8Beeccpa
iaijgQvebXgfAYh/fY/kbw0BcNERQTgedPwh9VC2aT/9g7M5axW5wqYW6SQ90KOO
JQ3EkvHFDNZ0N/knwCgUJovvV/oSekTAAnd/Dm5E4twAgjmuQ9psUQa0b0q1yFwi
PVGjnyWP5ZGxgthobtSKRdAK30GjUkKqucAkjmn4aKLfXBLlPT82IC8Jbrxsqhrh
8pQhAlebATahyYiRY/WYRAeSka77Crb30DYnzstA5j2jSB2KyW6dgVIWld3aM0Rx
FrUy2AxKSzHYilac1VUHiPccxbeIVqgAPMjO1xo7JOQckSv3w4bF4suF+Y108SIi
FzYQs3CwHpJyrK7RWzmh1WBJ/d8Edkd31o6CroIt3HddloG3EZdWSmvHsk/cPcrk
c6Ar/lVK2p2htTBqPiNOSnSNyGAgnS7eXoTPSIn85bu+dGe9AwfpWMAIEFBkMMyE
kLRGLNgZEyS5XkSjLfSEhH8pueCvqVPmtFj9ZQUcPW/hA5cVJNL1uY7hb1pi7JQz
ZEApGm/AAPnUR6r05gguIjZ2fqJrDmGOt02k4Bdc9tQC/LI+enSrPG6RWX0SLCvp
VDyFYmABm9AW0elufc36AjxgLvMXsD3vJerVZU0TxiUougjMskTlK8gvm9QuBdac
ZxlnxjMVDfQCtthg15GBFQBcWcvHqQmrt4DkKoINIf3OVqcQHz0cnN6Z968eeVfr
Nxpv6tiDoJUEVSe8NZtNC7Ya6LWSIm9VJexNhwb5EVrpL6skNrmQjp4GFsPxeug3
wMrYLxAO7JNlkNb79/E/QBqich4Y0O/zUURVpHk859UZ8jDPUv1lnmZckvlp7waH
Kk0Y81M4znk/Hp+Xp5FszRxsbsVR+Ji33bKn2Xbl0JK1+JQFns6KJ8p9z2c2V2xP
xAHeayhiArHSBT92avlHtgjhvkxqHy70Y+v6USTcOWjc3+gDC3cf9XlFeQZwYqqy
0pTEw3zIPioj1/mZH/3A0ozyydCXrUqgv95Jc8ovDamG9e9dA21fe8VVtYV1QGVx
9/BmI3ijiBH9Yo+bBCWhTftXGBDQ/RIqjVFtcFDP6LiJU1WxCshuYU+uRTLk0G3U
WKIB48M6tMtwHwqSRLJl6ZtjQR7SVOjDMoE70oZqpjU2O2VlRUaoGdJ9JaJlYO35
iU1EwhdfTtFi0o3APofob8EOq2poVoCjYUBn3CUmMKuqy0Z+GE6U+AX087jGJJo0
rtU2ouKFcH6/nXvruE3HNcjL+tpNq9Ck9lks7/6OXPHtZ6QjjcbYmldOJtecA/V+
TQj7Y1MQq8hKvTko6JbcZ2ZqtRQLsyVGTMidLKfQ3i5IAp4yas8IJ/Q+9yZA1GN5
AKeI+kCM8OyJp8XjhtAQgXTR74/Wi8ZQ6OBsK2lP7DNgYwvq2Iw1zbOkxYDi9JGE
XNiucEwCRZELtN2o8FPVwIcXr4OoKzYUmTjBhEiECUH21dfL80udz+qBfSOLgLxa
EJVK/9mXsSgKz+rwsP4XevruY69WIcrcM73CkDVGjQO2pYMJ67c8cf5jVK+gRH0i
RNrrCASsrp7cbhGA3+Dd6mVUehWL4tQF7XARkbg//dU/Kvb8SThVFdKC4A4N09B+
FCswqK1ffxv0qMxsyJW/0fNEncQIJGWtRXjH1ukg8eu3YbYMfQ8ccTmqpkIpX24a
s3mYKXd/Cu4WeyBH3sjrNeOAXMpcGoFSCZL/BA9Nim7jv3n6qge0uJtXqjXum0Tm
VigkpdQx4Q36J5DGaln8K0uNiLBby/nfVRsNyp5sEdV2eVXVBtdIPGLuZlO7SreI
JuRvtv8ZBeVwmNqiFx1LYtM3mMx7rhhkYhCSPe2acf24myfm6R8KExEvrdw7S4uy
AS/9VDRL6W21CxBHWNR9BUjp0nt6aqNwX/pCI3e2InlGMPox3MHtBqagp0JgCVnL
TI05+Ls61WhpLkNbrZ0A9kBigOfKME14XYCRpTT1LoI8xt4CvhccTETyvFL/wJCd
qLGvy4ci68Boqk/P0ERVh+DiauLCu/1W3ee0lneJWYKNlKFzlli/99OQEFjW8HLZ
xD30XmaYpD0PXK9plW4dgMGxWsrvWr9z9fXQ4bR49YFfijyrjMpWbGPvBOquvTRu
Xmrb3EcNT6KIYXUKJJRtvxW07vLn7ePwddzi/l82p2WuG/rVnm3k8he9jpxVvz8h
dw96iXVSe0cUvYA2vBseFXD8qgm7ioaHHOCOzL1e7Ae6KhwqavgePUzdvy90VCDX
tBdtnyCHgf6S8x/6kIOjyuUF0+Q4CfApvxaKPt+SKeRatzq9x9xmG2DFe6A25h21
xDhh1Hoii25L3o7zonHrYB3N6sDHBB5Gkacs+ymaQLATtU5Df8pM9BExcjllx5ub
nrJmvSjzCj9tupYUDxjq0pre4xxkojmPZJ8HSmdXxISY3/7Ug5NK/cqmSxRXZCnv
W9wWcCRTRrgy+5P5FwYIcO/fFHKy+lAYGG0vpWnntk1febD/502/JGh4RVlxKNBF
V2ef90vRfNTuClulB6KPOGcLX4YbwDkZE4k3WAJ/exfHTgqFkbpz40QoelO8FSw6
INVMc1MZPkIw4rsYYHcnRN3dyuCA4VlAFZ7+7WKyUkCkv+86Y+ToNSPekGYisOb3
DD/NtH5AGM07KPI/T3xtrXqnKffV0ZrfSl/MpmiD+Gwe7Xf/7Nug9sqblLM5wAfQ
6gsnGTLs3aHKepby2W7bJV8XQX0+Rta2hbCuSfPATGbNYQCAUnx4rFOOHjwOSxzr
XULp2vaSdOWrtw0X7Hkm52l+VUwpuHpJJZ3ircZyh9m7DR9llJWSVgy0NZ6F33Da
c9V08z6chXQ/+v0ZraFfH87mYqA/CsOxafILXfbJKkDyJR7cn3bGZGmbKi4fwuB/
RMly7Af9fMajfKw0ON0Xw8uSq/K3XlKkyXd+qbkmS/gI+qvIpU5gQ4YQR1KrQ8kG
y9ipEQFuRO3pg7+MA23dcIt8XseX+2OcPMt+tn9yvr1rwUjSaAkWGsgGIrkLVjnY
x3P7qvGWjT0o7twQVk8QIcjRlp4ssA8/ZMd0YMJIR9D6hbiGaHZr6/gnjY1vjEbC
T0F915ywUQ+++HCo5ez+0GeG1H2r5e9BtmpxfX5sH9J1oJKYmfzmHv4ABovJ7hqs
lZgU4plDbEE6BKFyQEMoNGsIAlgKcZkRT2a3PSc+R2UUxWrKQj7fsQzwXzc6NnBx
ztOgW0v7rWIZ8E3GXiHZ7sSKNhTeBsBbCUidtzp5JjBOlVaCNN6IOURcvOMorwXo
5ZY9sUya6xslfzeEE2S6zfUu5ZseOM2nTQL5ki6p3tzRuJbtwN2XzLHHWh/u9Xsj
tfTkjGZOQj3lk+iqONEC/+jWvWdd5y8zj/o5Y4fdrioown6hcT3J54UCbDjwRga+
2VOpv79Wi6GDnkvnGJHOUnLNRYfSH2FCslieW59fRFILfX6/EMkxtAxf85IEXIwy
ZaVcJb/ZsNdNW30yqKuvosIEaKWt9q/NMDK6MBoT550ybujHUwn24pjQ9LvxVeTy
mQH1EYlq9M4EvmT4iJUGASkSkYpdhPVtTNv/8a/P/CD/VTpGonaaFpgasJpZ6j7x
apjRpbG/JXPk1+CglRrX00yyfgSUzktDG1GZjysz/VkmA1qggRavjQCbewvsP5r/
yubD//rpwkBtKrexFHDrCq6BrCbXhrWouZPQU8LcQ9FF+iCn6ubE3Dr503S6W0oa
714J4rMvt8m8MyC3a5qlayLzeoHMjF28Y7JGC6VTf8E3hbMxGyK3vqTVlNPTIZqb
RgCZNBgGu8JyRbDjtCp0/nFKVNgOknjsL0+ZeE8Yc8idbpCN4EtLP6wwvTWCuNU/
V911Am/akijQ5h7+UVsq8AQ2YlY7zRaRXv7IafDkoZhXsSKFGUltOjiJ5BnnHxBS
82FpceCqDpqfZJbZzgc8svPf9fpW9zBnNB6sm7EHxIJoKsLQx0YoyeU49YhcwB55
rwxYA9vM8AViWbKUam9pssEMntAWzf6DflpHfJX0C2u3rUe6pxI/IC8OPQ90hDID
8K97trwXvDdA4UWukVdngWyL2X70UBbHXGyi8spExPVHPJGjp4gyq4gLlgxUNm0k
onb+DRSSyJYfMLOMKuJ82Jf6OvAzi7P/9KrW9gEsOZywBDLbiBSYVsSeO6iob2yn
iVkUVyobav4uzeEam8kZRW90gMZTNW/djOnjeQqqPQhgy4rju0JJqudXAmkmRGgh
tiDNdxW6+joocAM0WAxmNUCZBNO+cTtg75pl9EbfSrvQNrM4JnBWyPnbr80agoJm
j4BoS1JMqYye1ktXlQhEsT+VdaAFxvjfS5Yd0Mw6+ekBdsrEWxAuPxndXuYM5EX4
IinctZM5lO6A8XgRuyXT+tEkBbqbl2idbqrJxKgdyZCSsbpn/9WMvUn3BdW4afYT
5rW6RXD1bm32cSeL66BvTjW6a53BSKLIXrqkUMkJGCGV4rFjlJMhmA87ZIGIYSqp
clmMyIgZwYuGzrtIyhKR2bdjl7zFkbsmvkNa4Is7Zto9GFtG+BEve3umQ1+hMu1D
idnISbuFo7f6UnnGzN4dTZQo5n9ClfdP1yKYut6/o7erqrjKdOVHrQNu6FTAfROW
IOt5ZSEXy3Z8Sv8i4iSEGaDmLli0x8osj/enc+dHKZSa93c9PHxzRRk8+/H4jQsC
tD60VtETOejJOM87/uuVtzdpRM0jIWVy56EYlX7WoetMl8IQVrDH87cinruyEMic
2FPJ5KB+fkTFeFzQdYUOUXVtHrFrxOO1aEQ0nQUFujnTAv3FK8P5JSRAC2LboucE
chiclnd5tirVSr6yRH6WI2QybE+Tt/nRfUYV5KkoX3BzRQ1+6u/i6byjWj6tU95x
8BQYKwkDaEhgnga+lVNyn33Hl0A5TCVY8TvC4O9SBj+sf7cBXacKDyWZ9VvinBWW
UsFBEeV8iYkxRRC84haWbZBMlMOD1mWROL9lpJH85U8nNDMG8yVFMRUDw9M5L3B0
5weIZwZ7BwPw+lnkDFZv1oa1ResgLpqGuahuPZrmMUj5aNkY+V9bDMOE6R+4ISLx
RkWk0apU5ozJ/8H0EEmYXQsW+Rd7UQ2R3kWvZMNhgLhcgzUDjTJ1BfNFG97DZyjg
uimb0gaU5/3kxhSHbkiodtyADMS1PBYDFRdJUgMkRPQciebmwx4jWNpSujAAbqZD
M3BJfMke7udyEhWok5qe3FFp5tG3SXsVslu8eoZCtg//gNQ2kRhYCJvDI04H1xuE
DxVHSRoMszhvFKRxY7LReSjIoLZIvewXmE9wzUCj5O8J2jidDIhsKiFGyswwmqTm
lJxEfOTBRzoNuqSLRfY4R9Kyna8ZKw/xByWD9zXWay0z0jMNYE8OT/XaWSAPsoGw
wtQzr5PLtaIJ8BwwcPW5EB/atQ0tgy3eoguIBmKDvV5JeoePDTszpvO5Gi9jt37i
A1KXwrL0i2Xi94oQPOBlatKI4nemYM6nQUxDJfe8eUTy3po58q+SnN7kpfW1ynPz
e+O8etKzHCjxtCSXZYodUzayMkK3uKaHfj6vK1YSL4vbviz6uGwLB0+inJy7T4AK
PUHTBBCfZOQdjMPWDA5psJTrUthe+MJphDktH/FkbhQud3jl17bFcAEgwX/sq4Cr
OwzSseiuI5v7ur37FvSVg1Bi8NcMeu2M9XzWXPvlkpYL9JBftgfkLA+52T76euhR
R2jgxIP5+xQZ868JYLhHhKPh4GXp76ZusRYixRXR+yI7nrkSv7lanWaKvXSWXGsf
E65K298x19KJc2P/2zxZjJl0qX5ODnTJRHBdsEPDQJvj7627GZMIUsIpTe2pmuuB
elbR1CBiyKeevQ+7d3xf83LovW50uoL95tC11mvPJtg5Lqt12ZCCqpueVYQ95t6f
1p0sxfh/Lgf5spNWgwjv6/hpRo+OWrIkQbaKaJRRAX96g8fOtT/Ir7ofATY6gZX3
aD8QgPrR5C05N5ZLY/31yCfn2Wo7HPaIIuya/DuixMSmrSENebcbZ/Ai5fdxnRGJ
DI4qzPB92DylRohZME0k33n6sTtxqOrI1qgmR2AfMh8qBZbHZ3jA5EOrzEGmN/Hc
HGQPpLPAM8m+/LMLtsjy/MMjuw5BXUcc5X95HyRpeVxcZJk5GIhfkJQg+dniKpT0
8cDhjHEx8zSHT98yxOu7i6f4WWpeFZyzt/tYqEr2/muNLLP7Cx0uA94xBJ5Cxgdu
1J7x5qxvTYwLu9/oIKQTzA91tC40btIzt3W3zVl1u0p2/uz6EmPfwHX0lMpn/EHN
u0go57dp3xkYX38Pj8/QapvZ7DHt/HwQCC/wWbZGwMAWOeP8Y15x/NjMmPTSRFyN
fKXXuQwAxnPurLNJl6TAACw9OoVC7I84I1vaBN7C3xWksNEtLG3yAy0ZsfgHsOVm
WanTZwkVJilxlI9Hhy5cW+gH6dWLhOzt9m+f2L5/0Glzo1d5Fh4SJwoJcDNZrPlk
kABG06jKI8PMWDQ8rWDIfPPs6fQKCvmo8FexXllZtucQ2bPkZAcsMOSlAeNX4aqp
fstDnBxXN/ez9ntOqEZ4cUUKm5SIh1jvnqfg7X6EGxDeMJmtQFrlUuRiZ8GaZQgu
5Y0BFSbG1uFy3PVJhzGVISI3qG82B/ecm6geXQR3tiS0DqOfCs+Y6QLPe9gWg4Rj
3e/PgZOpa/Vte56W9pavxqDJ39Q+944zn1Z4VrEdag7VQxccROkuVFw9xE6Mczls
JC/dGT83pXhm6Ln4nFubTcmOar3RvEaKEOIAWc3HzO1UkGCpQNEBkf+wIRzugCOI
q64OJRT+0ftbR8VEH+qS25sbcFWItjLPQUvmxd/HhRaXtiTxTV2MlOYiU7J7xPfk
3tC4zkNU1mQU2+CRX3mA8BJoAQ3rAVZVn8ZMIPrNNvGFo3ihtr+bJcgsdwIm8hz8
a6Aw/PyS+Z1bX4ccXcekGn3lekaOPwzHJYh7AXof9wgRvrhiJ99i9qPh+M/rQb2q
r62hYVMwVdXYXAH8Cg/PvdpjImN1k4kMnw1KrStQy7gev44gSo5BiBKn7MqJCHaR
TnJXH7tyagtyQBhAxOvhZzNmIyot+s2YPpnXlGSWhP1KE1sl/S50znBU0X1vANmV
dItLehoV595SsF45GRm9ezLakV17wJuL4Ks7n2JM22nwDMshOQSEYBqKyvH/ZXoU
dRL+acq5jXxPH1nDRKIsxfsbgFr95Uz5nteZ3Q7HKhowRuqgDWQSOVpOhwJEGW7N
M4sq9JAIqAPJq4MeXwBz/2GDaPw39RNUrRqTK5V4TYrp4/cITGFq96iRGtkBHHKl
nv67vyIlkffMyytMxVzjoo0xaqEMWNPy57NnPdm33vuyS6qfcWxd1d174a+TkNth
lDlegr+G/NgypC4VmDO7xCJuWy8p4KF2IXS7L0vpIu6lbXnRlLte4nhrVjS6K65Q
y0pKOCcN4+Rt7khHBlEhppvrTQoAoK/f0SxOvgoKxRo5hmJ3aGWNPArwizKVGcWi
wxWkPkUWTOhYhhe2p1pPnQYuo5qRTf1Xy+LLnQXXBoCP5ng+IgeMZZwyMsbiBntG
ZNRaI/NnWc8380o/gtvvaXzIOt3VRyQAZzOmk0Dl84BIqUquxwBR95acONcSNn79
8Y+naQ1vUYzChLzl6lKnNvLf/1m33umjvLJlTxtJd7T3ousOySJOx2AO/YjszX0Y
FKIXONUme+ASCtwEH7NrxAbODD34vb0mYeZL0yOH67Wwrf+k/D+YOf4nIBIBnDve
cA3NcaEh/PA1raLvHc2LPfl2w6jlBNNAddzLgrYeSjNSCrNUpjw74yuY3+bGOUoH
6Tda5y76BaNWLT3YaHA1xri9UVFiORUjhUA2eWUwDNgAhtMl0PXFwJOa0y9uE5JG
oXDYO/BwS67jN0lR/OrF+4RmbMSkTfaLuR+xOXdPcNlZhOBV3mGi7Obf5mfwtROy
xrYlKJanLi8xj0lk+xEOV2v3IeCJHPUrNmcuHlIIVCZ9qFeb75io2SdlZbT/1DVp
9gySJ4tVcqXZPoDRPwx4+lMYQBXYRCX76z37bHinIr37jLk/w5zrXJ74ZG/XP7/v
kQE2DgWOlvqL64iibpzphZqZzg4RskoITgxSjt0X6/ZWi6kxgqydoFnccCW33cjh
O3N21xa04xlkbQUOvD0QBLEueuMfVq1nRtlzL8uGpXlNLK8Vg6/TQFTDbAqk8jG0
+l5aroec41z2+N2xwSFl3OcyT83m8MUYJ/lZG/InVMz6Y4oayN7PuPoBMoOlZhJr
fj9b9jecuSUkcA/4EyMKuW+aykbccmhDcbXsP8EtBgd75tcDO2XFAAMJZgiu1MFD
YIkBKJIlEOesC256o6ELj3vaPJ77mY6lkiW9neRQdDa4NiHnLS8EL+qRHx5t8spG
oJH3Ld/G+5z7jndYXXVa2FXLK6AFzyEp+zukfn9Vzh3vMVKQ9d6KQveL0qZIRICE
rHvFJzzXlhWCMHEdGPJV5NsBvBE+fzSjPLJh+VL/mnUcCyRqbVW3EwYwGNlYCyHV
RP2ichCggWCDkCOc+NXD9gIq12eBzt4DfB9Ml3kuabYPCgaSb0ayScsiNejTbVYR
An6xQDjbeMnwgqefrGczf0TT2PW5nqsfIAkJ5LEoc3+jmSk3T2LhWfR9zXTQkd+l
EiwOatreV/u7pNOJTSubXQaRzH2+q4NhkiyB7glQJ56uDe3Er6bnWT3nG8ks+9CB
h3eu35AYiHJSWH51hgVCIkxjoEosEuEYrf0YzkzXEx7Ml2uhLWZxDqVMfP+/ggHw
hT7jzd09b1OeJ7OF4hy+QDR0k7h2X2HYFZkIhg50/91/0dktdnKxIFfJUXXvmUEt
4MI6xzEB20gM17NE5mEkFIaVk96qejgINXLMafoLlFtrvIJP6n9GawgG6/sUst/+
bu0xOq+vlnaYLNH5te4u7M22JjoJpXX2vhJ4CxvLG6VlNDDGoK7pqI5s+CIqg2YN
5JLUMcOddhlNq9iBTLSfpslp98lX/a2YMvC4jPKV20jglmxSd3qah1sXXAVGqjqZ
QYEsBoMqPIeVwgveDEIl0d8D9pBBzD9SSFeeLpQHnAyPH8MUIrNXrs8GEzzYJAk0
h+qjWpZps2aqA2kcEMgOMnxLXwger4810YoXaXcfethRVYQ4Qy4B8WUEHM973rk2
0E+Bfo9L0LLX//tGP6dQT3dS15dCgCw+Qeiuyqub5PEikepZDIKjbcM6dbffJRuH
Y8WBolAhph7qTehjfhSH9qq12koxMZhz1e1MV5urpXhR0i1+U8eP3ZdnSZqhNxnX
4yqrJEbVf4Fd2c6zOkBPqta/LNU6MqF5ZJ+i9ub0o0WNnVULctC1FFFEKIM08NHM
58bKAS3rgaATYYilqeK9IDmR59RW1MTX/kmkSv2qOab2Q0s4jC2u5ihCjt7Hs8lJ
60UmzyvbzSi/UbvU/Cmrm25r4lUJ+xZSTtp2r2MKw7CQheAIPCZjwG62V+FuTdBU
FsWIl+wFHt38S/m/DFASXtjrTvEeBCCknFrwvZjueWHS9Bobh/wld2vZSdvfG27B
WxLTk2XBATayY6wqOVwl3vFBi14+2npnEDkO7M6b1345NMNJ5VeYRmksnDlke7TN
PBrSoGyqCR17yTJBlqnMyK5hTuajfYdLcD288ORNnEYc/Y+57WhOwJdadbYOuNqk
VgsMjD7i2pThqa68MLTs6iBJPsDS+dJn+X13ypl/NRFXmAfXqTGEArsQYIcFlIgM
Y/BViB5ALqrcwchsO9LN8d620RF/BaJdydCg72YXtCzu6Ob+dBobCOZvggDCdKou
Ig3RsNT0qabo0Zvroa+W/Au/hz9DqqJu2aFhON09cV+nsvksTg39zoYf8xb20MxW
G+p4BwlVIIYmu+bEU3XVnWrCBFHlb7uadS99UoDJUsANmcbtqUrRVNH4wKzMJvav
6Tc+AJ8tZn2zZ8jNTDdZFgSTXHZjML30KSn45WYv4yPvWojGVvi9fmcpfYOj4Xc/
jElL9dxdJxM0ERrPlSnqq8OEnWrGIbOtCcPITYA26ynMj54AMNXSz1dE96whAhvn
2+zhk08Gk7vujeHA5Z7onvmChjQZbklhcfEfnRc0VyY330xoC51//GNQnVTrIciq
U6sFIfX7YiLbfyqv9t5J3HlVkkMUvHOu/IumVa6tzPf/AJj+vAVFmaL/RnoPoPoH
TIwEItk6tiAeGkYSB8/nh2h5WkkZuWZxO1pS3sTcG98TM8rxIu2tW0qvVMk3e5kr
5McbYLv9JW0MIy3HJOAqhLzVzKKuOdie4dDdjUuYJhUV5O2vBpMsPbg7oW309zWi
qJ7Hk0RnlRDldx7wEd7doDAJEaQ5EAR23lbprZ6vj/+9lbQMM6Zb9H1iWyiuLj9m
8AF5J33nXS3F1A7FN2BjU5vEa0/YP7SHAJF2qDDeuGU7+f5otRI+OzICsrteZyau
IzIHACXcBNQHl65m8fYjx1ZXV1s8vjZQsubcGFjbdNwbyE5F2wvG0KpH+5VpLMH8
ZKFleYepxHabVpFH5KhyOrfZC33x512Vwstkz8TV60Eck3E5MLe+Ntmd85O+paFu
guEM/+DSOr5YKi2K70CGZ2TKd2lTgiuCGvecUTkXefoO+PU/5BGwy9EOINYFXwPg
dSJlwOKtv8rRChk09kDn4MwSF/YPTpdfS8rnPtwDr8uEcKpbWB+BiMklGPg+ZMVD
oM4DKOvWAvvxkUGZ6E3hUiOX7T0jKOC0t2eMB+nyahFJeuoEL8dH6VAP3HahbVgP
YZws+kE25bkMHO4BZGdjaT/Ukm4JvIGyd/ldqdOOMS+Hn/OOumuJ+KZNOvl5H7kM
4ChNMqTby30Wr2qolCS6N2s7XKt1Od/AfBgRIiu2ALkG/2aLcWphaFxiZzWfsNJx
1LA4MA5wuW63UBYbRthp7EtzIU0qxS+4eRTFeLXbZTKQzX0ft7QkaW9E+nBvY7fk
bBEVROMT/RYHyNr2ekT/XAILbiLxtSrbdWoDUgAvw0pir+ygCITxoeytvTmVY85D
f3hZKTBQHDf15HCWN7yP0s2ZNnmjUWIwBAre06TJMhQXwskVb+3MP48VRAucdW9D
59nZpqkPU9ZhJPV4DUv4lIxxzdkDBhW0fAmRQRAxa+oLaHr560zhn6cDjlfiif/t
qXhQ1cyDVAHXSLBoXI17oHleG4A0jPNJFkjw0owKAa+jjR3bO/Jybtt06416a9sI
UvVXUW9t6jVCCBxRATT1SGWBAR+8EaC9SIr8o497PSIq8kjlV/qHVTM5YWBe1reI
TvMDdTP7WxGpWH4KB3Zth2Jr8HNaT9LHhpl2OeW+b/7ilBu4NLH9yozO2dF3iKQ3
daV3SzaGMKjGDFTCIB0sjnAdVUJ47Cu+OXtTTOOGV9kSHMRCg4Z/ODyfyORmskw0
ED84Tgl0ZdA6VdoTnoX/poP+sa7SN64sBZEGZnCj94s7mZ+7VT55hwDEM8xH6JWF
P3S45gUhd2HEOxIF3fTwLFOcqoClzcGCQfNOZ69iyOCNOJoGkGtLYaOVtE2V9q0r
SkZfOxfuKe0JySx75h39J0yUaK7UEuniiBqWDntqZafhaXSi/1UVaPRs1OVXgCAl
8bUcfXfoFEp8KmBpjB7rEvyBQjIinzgosHgehRKUAtnajpVppFEOkMaLG6U8LyWr
I6pUAyBYgOZ9wARlFf33tPlnedJcv42vEYQBIelQTjYyQ8nT7+an/Aq97bHFt56a
C3XK/Lbg8HlIAv6Tebd3w+CX7y8pKkWz4M5ZXvKjZsHu7b3FnlVnpXxPJq1el6r1
Mv2/hBpG8IzooGH8LDFMffc8V1oDhPfnVo8LZDGyBOC1Og/WtHYecoAhfd/YgAvQ
80lhH4mdnlNWfy1AoO4hOr+yKpdSV3y7gvS+PCSGkmUu75w5n/rHX7fmnjkVQbLF
nbjUFdsXJae1+UCbzNOnOJfMQmGgaYaUAU80YoKMyiMlsfRD9V7sQRiB8Hr/yPU5
v0iMBPAJ83+sLrN0ORFQek+0iXnBVJT89gZXGmgpYWWtkN7VOmb+ql7Bd8oKahFt
0jxdIpxKGZtTzjoI1jnzDm0w9GNaWPKIFDZi39bOEuiHRYqL40XvIXj5EW1RnAS3
UBgS21/t427+82o2jhxvmdpRxA5Ubhmb+NIv3mIe9jdMCSd/L8IQ3aSU1yqm2AJI
OCN3M2V348EqFs8HgrzSGrojT8sZ/hXT1n8MGxad9QrqH3BgkLyMm1aunul2OD3H
nENWOuk4qeh2jJpV59hAJnVtLShvZZ2pDbePOGNpzzz383up2K3yFudqKbyprQBF
zyTLU5eV7GHwHbepY6r3JiE2fDR7XwdvDS2mFSBS1VOLyzkrpumBLliCjP6v8IVY
BaCHLLAN3V2XZPrCg533VAltHsU6HlU782m3k9WV9C6OTtxBgbe1s8Iv6NE/3sA4
T4T/ydUwsCQw7JqNDZyHpabBE8o8BZ1giarxYZt0U52mewPzvAIQZJ0lD1VzFZem
ij4IkWzIRVd1nBd2s5WCSise90FtCLoedv9tRyfvlyRp2rhjWng4j7c86QWbknj2
Uvi4Wj19Jc/VhhajsvlYTU8JvyKOU32QMbRGLnTALay1ll/uwRSVIrXu1di1UAFk
D1JXNkrFDogeGrrZ2AFueNvWFMKb0X+BUk2XyhB+qZkuyF7EbZjNzYmEbL1Mqy4J
7bNZoQbfRa3nhZBfUyjLsZM4y2XgMl3yLFG+iZ8IbKVm0w3LHn+Hd0aEz1HrwbEB
myLIym0SahNdpNoNxWGyQsZxTipsMSzEYqwDs2+ea40LdmKwB2eabK+PtC7FSQE1
FGXPa/uokWAGn3HwSroxPzRLhXAWfsFzvmKju9QxsQVFuasekxHkgSW123bk6FuN
fNYzDE+Le6H8ea+4RoL6RRDxiTmrYZsiL0OUnCPrUAMEjPqKU5QdEulBeW6iB7Nh
OWxNzRA/lGECzhcxJyejDuVC++UNbncLT61x5hzqnoFyeAGl5AhMk4wm5ic9dEk/
pwnXJGsWc2KIOLwfGEPAEWJMYG1hrH0dRArGFpSz9wmbjjT/q6T7H/PCAjYhguWF
w/gQnE8QhyOgH8vtf9LSy3hDHAhBQMX5QAasp0nVz7BVJ44U9s6R16b2BF4oTJHH
mkK1A0wEuKlVF3RLtQMTyy4ebfel491FX2WsSmQUxZ+Oo3s6rsauZn1/RpXa/QPb
rvpWewux+fB26tzmamsFYYq6hEf1dFu0EbO3EDJIUfH8u6MuYMIBgmvwfloV6ZFB
S/J0wcRvNU7zmzM14nCHdrjQt9QiHXJkk6wCm6LJXJw5IBe8MZxpLcjbQYZIzb2v
wGCcdRnswpOlT01E+VvLl7mi3+ZVS1K2fQf8ZMR6MeDD8e44J7r/pM01ctRO3YyA
nU36PpFiKMmnQWluDKxcYjLdWE69UKVjj8LrpDoJPdsONdyUrg4sfj6HPKfxX2a+
eKtp4dyRKIkppQceCfP+c+Ozu/jy0GvvFcJXRVl6cQFJ09dwm4y8JuPAjFrJYyBv
CWteNupvulezUD+9Zj9tF8s6X7nhElobFbfcSAYNZwC8lrDlVZNMGcYAU6LsaB47
comlOOBbPWULrLEHA1+Yo9MyviT6/kaqIbzQRVjB+Bw+cIAUa8h/L0e81M6PCOY1
0LiS/NsjyOttjWvRiwpWS/LnHqXaN5rht7Z1ixaCqrLkJATJG8d5Op3SDiZLfzQ3
zaWD3fd5GE6/gOvruJp31zJDxN7v0f9npdOCUtdPt2xTPY0u+oEUcngp5T/VwSLr
yRi0GRppmPU2IHyV1gIY7/LgJq/dElLCE3T7LZz1BH+343ZtfLerB6kJ/P8+nopk
1bZhDiOHSXP0Ypqp54caT9h0Lv6gLUjXqZGAFZoq9eC/uZWRTqBnwl9KJulVhKiF
QbJEf/ls4aIitex57v6JdAqHCMhcTmL66IFJ3Fk3NPF6+nzbo+F4ebm9nUmg/fEk
+XRxHQg+PDFbPvusd2VrzkVOmiDMdPAzV7cgybFpG6HXHSBnwKv0ewYEgP55d8oq
wBZeHgc64AIQgm15uH8egaU8Cgle+V/ovB1Q3kSI0dKF4AMXm78a0oTdGmeX1VfK
dY6ryUWyrXGvAYdhND9tQIyb/1PLn1eBqiCm0i2/4oU9uG0P7ymX2coe/5rFblH7
ROzaYGeOwNLqA6eYPI9rnoIWgYGaHphT+EfSwJ2bh9Gz5pm/GuCdBe9G1LC3Qq9l
2qtJPf4Cu4Y4FH1Hgza5el4FcULK8/GC7n6XYJ5A4NdNoSjSurGq+eZdVAVQ6qcT
73+RcUj2wXwHFIhauXpSAElLoY8+iao11U2e5a4G7sQQeNMOu0UmQGWLq4QSfdP6
8BecBBA/46UrsRp4WBOf3/PSGdrLi1gkmiSS/dXV/mmRCXUjoY0vNRAi91B8+Qdp
CYfZP7x/kcC7JMWreWHSN6zX/0vXG5VveeUEP97MDI6LxMLPbc50UEw+/oVkJlE7
vjDHptkaR/IBP79R448uzXLjfL3tVTxl41YJRN6ZIuTGYk8Adjv+xYjdlq6YhTSe
KS68ndmXveFKfMPU4FKm54X7QvVKES8d55nc/MWRaLquC4PMR7WVhtEa3GpD5Je9
81udTY8csbustpnzh7CDTk25GGvg7ZcMfdOOQtvpdtr+yNziY+LcDXYL45HycqG6
4mMGRvF2tOWZ+8hOgbaebwmGHCnDSv3/QYdJOrR/676br/i79mya35p7R1kov4gB
7ngg6l4WsJTFJB3Rc3wFVHl858xLAVf34RVewJCBUQJVs4VIeihaQQYoJCCuQbvM
x0b+M504laIYRunn3Mv4HtSLhv2CYtn2WwZN9OJZ9BljaRqTp2NOH/bIFW3tW9hO
NQ/jE3v2TfyK4cg3jG9Rm/DGK6pSL1OdmWPtVtR3Zy7vfUVmIgn5F6tftQ2LblZg
2GyB9DeIKWIHMxU8KRJdZhbDLgN1I/guKr2Tdwq+huQhTcyFQ9BxVS0ds+FIoxC6
hwqUCgBAwQmrKJ3L1UuhoJ6uman1tk+SIddMge6ES0qm1CcvBf6zAnbr0fhoX0iQ
PV720pIxcCGrg83dGT1qSr66JaLtZ6KNdBdEFF19F8wYCIEOW75NLuAzjRto/ezL
BFX0lXJHr+mw/JLPuNazPwuhNf78OaIfd7HTl+2JLvmSUifE1RmJjhpBGwR2r1pf
wVNC6ZbsQZfTouEKif+vOp4fj4vb9RNvZhaTkix8WoG0nSJTkdXQc5DTWE/DrwWz
PBEsKN6aXjjqrwdGr5fzOWPpiMZy/o2fM+Po1PNBWSe+KSWG3JsRRTE0l/XQyf8m
jww0whOCrfQA+2rQMc2ptW6LgTaBZLG47YYYiwTGcXS20c68pwdGs8d89gECTAlP
LnjvlFcBhjMuNCVPe4J+Yde3CQM3ugVCwBSUeQ1j2fe/+IX6jKc3tGv2tMhZawzj
Qe39tiTkqPz7mG80e0u/ZX1QAyhCoB9jyj/6hDlsbY9tsjArriecmtGiG88B8GXu
ETBEcMj3PAJwLyYwkNOzqAYjMMkE91661bSLTtxexJIXmyOuyUTKgUAc74b5FYRo
oB8YNIxWPOyGG3oZ4F7zlX7ZGZc+CPfNnZkaP/LxJOqyEKrwAcIVBYCP05ZrEIFc
0HBTyhRpnNc6F+qG/JvtRc74R2XtIIyw0YybFiJ+f5EzYlfLeYd7V6nrOC5z4Vae
VP3ao1wrDa36ol4JsBh8qsyP8onXflHD/547JeS+5AmFqGLmEHDpn9MqWXlUH+Z6
+pexQI517EbdZmteAhWOc3E3P8D7q/b/r5n2jTQ0jIHL08ptvcY9bqVm263QR2M8
2/whbkG90bwd4uCXwVIgidqmcJS+itYW29qqnuvIkNkVPa330gYFMfJImxNgz9PQ
l13vHrJsivwLMVEaT2hd+EawORrG+xVwMRhqvgXEecvV4U5rTy1q94Cnqor6/KdG
lD/vMh/sxq2H2YLd3IcNjhJvEC49WqJHViPYFIKC+OqCZxwJjUkoS7za2lRby5dE
OzFrwnpNSTrr5WXs/Ba0+M22UovoWh7dMMKUIKx0+qmIdtVNNK/Nqmt/j40N4XLQ
v92HXAJPkf9svi/IcPrtEBWM3ICiEy0jhd0h1i9UDNm0uYR3qsw1sSX86FJkndPt
ZD2g3WrElEk2n/BmVD+yoJb5fF2mGBmQEHCyTbarVdCn30iQgtlpFM/EOGIoeMlF
u7DSES81DPZzw6eQmvovvEp0OWk+e4ZQKsrDh5GmD6iOyE7Ub/ojt+6Hbp1G98Gr
tso+Bn33ulzhUMMwVmhqrKV+2Aiqifv2dzIkrZvgZ0fd/bMVywASfxmcsaiV3iaT
/YlQ7SVIk1CCjNfB+uY2zz6nY3i7HG3zi/PpGBVKNpkxg+KB3DnENm0LvQLhIYdY
5H77kgIE0xbhvXce8ZOBWoeBcb0aPzCNgl1Nu9fmplKAu++UHTasH712xxq1pMXI
BtN6ymtIZWKeVH+UFv+9wACQRpmgQmjv3tGxBPw0GoqO0iqqf3ug59OaWiYkLcwJ
TQ/XmxqYZaiw2vEC6pKWdO2pJCxmqJzfoDNX3/ZlBcPSqN28NBt397xlCTIQb5ze
Hy5T8DpQNjJx45Dxp5SpjcESyEkfequL3gKe1JnA3aBUwmaN36LVfY1H7gO6iIVY
7FH41Jhde0h0dPl9MOg9c9t0F/blV0iIm5HGSYHnrkQRF/6kuyD8kCthZq924u8q
LgcIloqU+4t/RcSrqwCA3nNjZQ5CRcKDoEbnsZa3nlJvXaC91RnIj2fqeLG5LCM+
2QgHv5Vgwpq4Ap4bvk8EYooRDOaWOnglCr5g7CNXkM9IGvRleThl9LEL8xpj3f+k
vsQnfDuFZpJTyPVEv4IZhSzqcNEgZHWaLY/Ru713JW3Ok3ObNKE0VwKmIO5efrdr
A2G7VPsCOSBxuRTdDQuElrWY7lrF4ucOJ4+GPUuoObAy/I3z+k2/TBmu3tfK+59j
PHZv1lrGxqPQpVQDzNiRM7adxYVR4FiyX9/TVXvzMIE8o0DqZGhw0spMcHw+DYcE
5kl2atOdrmxWcgQFF7AD07DqFwvj6UnNh1BfS/n7gWXken0RUWDU/yozSaP5rvY7
czcsi8F3Xk+ljdlQBQnwJYGwkGq9OmZZ63d3b7vP2KqC0P9lKOtbccZglFlDTuv4
hE6QJV+W/vZUZgyylFVUeydcrXmJbJAGIp8PEWrE3btgxyA46tZ/0aT+OFGjwO74
AlSN9ohbvV07md4G9MEyOR87NqVfBzNZdRwT60y1+5FinH/YrOD8JihNzSOZkAr6
RXi56m37uamnjZkQHYgOy+nMuLTe6v9T2ueunrEtnNvrqmAqV6hQ/NnuTfp0mRzd
Q+8EkipClcBOVoAvIV12RhF1/ts12wSmfWMsP0Q39a79aaf9hvITZbf51+r7owW+
jY3y5qqeSWQ9/7XbgbcJ0VDp6trIVKmgQ14qTsuE8wesX30T0L2k8hqCuPGMedpo
3pOleZLQ0MlfGzmjaI37xqw25FIRQcseLFhvAjns2wFtNFLgnY8TEWrzIPw8Aljn
TS4v5qHaVD70ckBMAiZ5ba5lDAqEbfzE5TtXEGMqYKTnViz/eW5hr4EuhOnTnqs5
XrrrL8SBm/85GjfkPbHFbwoHuvCoGd/lCLQv7pvFzbTExjq8nWjC30JF+MLUTGdD
ziYlqLHhDyxQGC5e40hoNTXNqAvNjhsCBpo6uQmIabQ+3Jwa7d/9kna3RaabU6Ab
iFaW+mBLCouHNWFD5Boiu3YTfB+gMq1HzngTMdvL0wYj/lflCucN6GEl2rcorRU7
uzvgE/wd5S3JAeEoQdlcBse9pxTxY7e31SHrTdgNWeJEiQYmmEyzcSK2YbsorQ8X
fwNJgFrtzK3BqZpsXeFPj4lZFfLg/QBjEsEyzvi6gci6H3ZYZBLnzuxiqQs5oMC9
KCnEyIiK6C2lBX1irZqEquceigUmnXkFyyD1TijGQamjg10T/f/wA7cXHkx/1Y59
Y7Y4OHcCUcsZhPE3vtVl7+miBq536KgjG8dyPNWE1pOmouRIdmJvrGt/D+pp5aMa
muaTbfh+OhjpFR/jQRc+jpRPtjxfwthW5HPii6qd6d7ZOwP96jJ4RLw2jshV6RpZ
IUpRra1IkfxSY35OQFrWZdK5uGDczUQrVbeJgErZ/OUc7Ly8PrNvw79ftQeQutNE
QFVHo1MabKpb6EpZs1+qwetuONM88CxWqe/ptRKtdJGepz83tydY9DLCaj1Djgys
m7edgwkazpZtiKXgDTwUUQIa4ThsWF6fXUgYhjW1fC6Pm3q6zT+5BFCz4dCH734y
J2/1DZTv88Hbi4xUqmk+qb7nEC7ThbWYXiY/hIDlr3xjtm231MJ+I7kwOyZ88OsZ
m0LouymLIA1AySIQEVm7yjm/qZr8jrJalZx8/WyPxhPWBebk07bItY8Vtgf/1VGs
cSTMKnEODoDO8W8CVoo9LNHV6VHBNNWEikzbRH5qA30O1uMyZYSWKYzCcGl2szqJ
YygtDRcbllLYCAWuFBTJoL20aYhOxIWOgEhq1MbkBSZfMO0ctWGgqT0ATeFGMh9l
RZhzIGzQBIHSdJC9p+raiqXTOvawfe/nhQyh6lmtbNfWul7Qrph+7Rezewcwg6L4
nhO3bjH/j9CJcyiFaN3hUXwEs3Az7FhDLDvaibbIuzN5HbsrDQFMBrXgS2mafl16
JrSpN2iXbrueoMv991IbwaoHUoCmF3wgozowf5V5sHYtGSoD7qdy2v2kdStZ9x6i
V4JzrlnkYjB8r7yRgzZa1qLgsrb750U7lFjF1bEelSCGVIDDIbpGGuurONKUnR48
A4juVlFeQty0VXNY8CmoHME3E/P18auJTNX1va4T+ppPoBjLDF8DKsWie5OFYjB7
x5bCGY7dPMMgfEGvaFnm1TAa8E3KZ2K7A3xheMCpgY9t1ZHIuIF7bkP+w3tBMWJm
Mk6k2uxMOGM7Wgu042jOepEi9CP/kxp2BcLzpY6qpr2usZr50ozZWTZfP8DJ5NMI
FBKdvsHr2XzXIfsda9DnU0YedKM8gMXzL20zR2ey//TmW5AzPqEyuDe/d2Yh0nA7
SwLxM7Bal87lU4ROgzmdbl7qHWzlKb0CiSVCr713muP7rxQ4CcFMtEsQ1eMda5e9
obFGGdZX9CgSdljuUjeRd4r0uMbhL9uMs2nstI/rEEKG2zjnHVBjEIxogKoqle0O
AidEnQ20/scBFQBzkEu7AkvXu3kMDj+k9uLo04sBppC8B5TfGQX07s2x0SH40Al2
0xKSE0M+JX+ThpadsRzM+8k+cLfXcq+3twOUvAGOrLuFOe0uCBtPD471752oaktg
w4NmQIobfgCNNGhxDZn1vnMRGwB7IQko1RKnMWy2Vj4x5Yet+eyFpS/Lh2w321OF
6bj3ZblaMWu6/MsWiZ4GwFEvDgDsKth5lrCCn3eRT6FcwCoD66e3ujTL1FIEAMMc
qselO6+bQR/Ct50gTwQCVx79uuRlgpXIMrjhuO1MIzYTDDxGV0MFnIzfGwdKO8PB
5dXinc5+Kq2DGxOOKXZCvxRvbSgS2ThjAC6HQUhlZBR6PP+GRFPQN0GlUl+v5OGn
iDsc7a9orhpnL/omMEJlRvpqXgMapSluEXFYiH3n8dhtBi/x/qYj82uhPw+ACmTG
Tgi8T3zfzGwGZDtdwaibfRQI0O7FLk+4L1Jc8mO263hrinQwnGpdC6f0RIa2WQfB
pYdZC+kVUvncFaCrHfWESLwRlLclYlyLAUqw8b+aUGZDm0ySn8GKeJxXeFvsvLxn
Ly5zg4bccBscP5wF/mCY0HANIVSmwuVURk7jiHBBDCz9rpj67E47nUSibfOHRZjF
nCZ72bSJ4BzYvLr2YvtcTgnQgn1J2RgC2g1d7YGHbFX99qbTddX+feWbq5eRqJNr
Onf3fosU801Kh2rqUZoGIF6Pjlp81tr4YPgLLerYYyljHliKKG4gbMiqldmiUB1h
D5NLZEzVW2eWIiHJmIqjyB0RufdZ8PhBaneenR3Xx2SCcCn+lEtvvA7hxYDY2aZk
jolg5+pRrukfBb7wS0pZDfrYNWtkslDnt9h4AcV7p1UMt2KzpVQ70fRgwwelMii7
hd5Zv2qGba+6pz4gVzkqEeB8cQ3Z5IXU4WvA9Xlfag5qq44Z94aN75BVtMWJS4co
d1AvIVL3mosf8rUb3GVn6c3UZgKLr5VIYTBV98QjyVrZ6M4nYMkPXY3XvZqfKYMy
wD7Bce6iVnoZewQNUiX6p3ICTdWl3hKYnu3c23ADTJEDm8YgXClMvKHDxBfgFNjd
5IVbiJFpT/LcmfPEkEJl85rHdiRoHQtcMerN7C/B6Z+L30PTxAVjzqS6LDzRaglU
laIHDbWIwrzBuExESNHSb+B5OpUYrNkG7gBm64uWgDEJPmYGSg229Ixhd67pZeaU
JH8f1HpS+KNWp/KvC7oqKC90+yJXkIESkvEe6tKa5GX2Qg6I3VX7ZkUdN65J212B
hDMAUR3t+jUL/e2P5fJVRRxq9XbuBudZWqflV2HFgfGl1BZIAVO+1+52FCqG+EvK
S+NOFzTBYsvL3kG/70RJiqfFY3zmhqSyUB+gWwf/mQ2FEz8wnPbxUhhSgbTQSHVO
hW1KIXn4XZCV/D4ON8LRMg7f5Fukcp4r3fprp5OzP0lrvNdZOEN3QCxAJjDFmVvG
I4k8/ATgYpdCZ1iwlvLMUOZYndw1dA4NksskSXEWfDtESLEciVuPYwZBAKjhJg7l
XAIHhQ4meNfXo4r4fQqT20l9cRMNlXgv6TSXZIrbpfJX3lyQClOwr7q2elRYYKZe
kQCYU6/fefAKIi933qSYdbv6MUI7kxqz0MfVW5erBTHtDzj779ID4zu/QheRSu+n
Qb93zHS72EGukjP1D9ghOsV5jc9nr6IQ3OkOEf46cHEvBOSaiAKuVGthdkHHkHIt
1+UY3OnxqHBIy2mv3v21D8bsGiEqQfnNuRWcNay6pFRUqHPsPf0HzpJtPUMA1Ziy
1ph6QHLEv9CDjhSVnC3DrWlnHOphK72lpfzVfIFsBkffdbpHVvdP/UJ74YBgZQhz
2eyMWbrr71T94E/0TrtDrkjfVaSWRboQq7gQ+qBNCqg9gT1mjmk3tVHtkJWZq6LL
vPb7WtCmWWskU0t2pQaOxnQ1P3VXTfcLFqmm7CDzAY8r/ouXq3dp+xH+qreC1mKH
CIHzHKOFnjHR1hoxp0DX7LC7doWGLAk3sG1NVC5Xnsey3KL9Pg28TN0Wgt6/59Sl
ijdV6ErwqHqnnRwcBvjmBziEqt3odK5/bTZLcTg4XzOz71/ApJZgPZM5xh9MDC3C
Utw5tBa1EJLnLHbeepc/RYt1TUzxegAgGqFA56HjsmBNOdv7mDBAdYQ8gUvwgSrM
0Q4r6FRdFQ9NPU4twkpRY4i4lJS7zZOQlPpCqlsoRnzoG1SOdWc+EQPJKxYkSOp7
6XJlho+XfAvKs737dMdCV+1ynbAZ3rAOuvaMEH0BNiWQI4zimH4n0TRouH5yGY0w
RmMXKMZndY+VubFenopRcBa+k1vYNGaCYqjqn7wul/kNxwr6TnFjE0aY9pFZxpO9
5uLOkoey+NZJc/5RCsLPAxNPEbeKYbAGKZJYK5jK6ykYeaBdFXJ3P7q4YuGP0UVc
/qTiy737zhUF7brU7dfii7GxwKLl9nUViq7lU0NOfXJvLWGS76x/gfJ5DJKkTf+k
puwej1EeYoQs4cCRHr8qWtopqh7/CYtYzHW8tHeQo0UJQW47Qu1i3f4NsN4bpXJX
FbpvUaydMViXMcoX0gKucc0kerCT/AFjuGSsakejSHT36DS3Y5ojItxQF4dGRb3U
5B5rCH8Y+IN/n1wCP47pDkrmZ/MhbICekwmA3QujsTxRqR1XAIrDCwmolOxiigYm
kHYPpX+eNbHYJ8aTCMdlmp4L4E+Y2An00oiCYdlcpQKjsFHhN1f34dHXE8N6B4Qs
A6jJQt90TnC9YJlrvaKYmWZtqDrp7py3ErGb5fptsRITlUAo6XuqY3QRtAPmZrNk
plBh0ToXIe69NSq41G9Aerk+rHBRLQWnzcn9OBZNBtxHo98EW6vtYxfYEHuJIO8p
H9ZYN+6FRwgE7ujtd8CM66rlB+nOzWqi/v6g8IB0vF9AehIr3RIdXn+SGf+C/UjF
1WS60hg5PLuyJXSTSVYzwxqYdqHcFkq4EG/9niil/A0FSUZrVeJZDX63+ja5Ul1X
6jBJ7uKoVIvN875UEC1hxiR4fL0YKKE6WHLHlxXYfVZBLKT9np1/q6GgwJW64EZG
12AOJ/TVEEOXpCMNOolAQYcdDl70VuC8O9boFoMNnAZSbkygpN2gXvoNBC0pGWpS
DhuCrFfOulqrZh9xjvSntgJ/KGsvOI7gubYF56G1b2c+7hZW+Bynw0mbQSBbzEcz
VOxkTyB9snjGZFWAn9gnANOxeMg+QCLiLxGsKGiwSueOntHZBa5Kyocg1z/XHImn
EI7mE2iK+igXi8E2uiGrf8r7SsVLcKKbTQ3AZ4FszU3mmfkDhyHWSXEMVlRtw13E
E3S4y2aXNbNJ1Tl8TGs6McNeVnrC27SZOeD5iGf+9Bj41afXf+W6bNToIBmsav8w
LdOBl0REW7O+gpbBk7BD5nsx6Sy6NvOI6a6FL/ztOGaAtNaJlgpXP7EMQxd+uvkL
xhNyGVgrdTomZL6jyQAObgJqLwR1QCtr71rkCvJGGSH9GdiVNaynGKVpBDE57auu
7ndvSZsLKjRynsGKeN8QK4Xz7BoBoSYeLxqdhdYl8RUwcwO1ca/L4pMkUUZfDG/v
6VcAjqwQW9MIkChRmKpsM3WQLnU53GKJs4M4A48yd5dtaugdDi5LDNhbIsd5Vq2i
5rG9DaOo50Ns2GUfZZO6leffrKvybT/HptybMDlQeTV7X0lqsE5cC/Hx+DuN3xC/
ffJu7Ff8Jjrm3fXinKgq7JaY/X9m44LIY1SIued2O6s2z78qDIvV+qssjbgivE9o
ZeZhUGZTLR45pRzyn0sW/Bj+ddojwpBa4wuh/+2E6emJomQE1Ly/x1UfuuFhloCv
ZuCnouXlHtL9sJOp13NkOg7g7p9fCWU/B6QzLCdwA1CKU0gi1MDEhe2y4RIHZ2gD
ldnq8cDpuM4p6iTL/oydM8WQfP0vCRMgg8Ok/LN9USYElIEmkZ7HpRtLsoQ+9wMn
LaMEb85STJRc2dtQ3o/xMkdrf9umUSQ1PuBZ3YsB0PXflCgegwg60s4bkteeHeXx
OYOH7rGAaW833SSpJ23FhAoAjNYbxp2jEdmGehEpGYqkLbjjwkeUFKXHdFCF6ZpQ
TlBNclNRQxU3fNFamd/Y4ZPaWFrgXmHLkD4EIC33hRUmKoJ4MCUPiRzS0M8r3VwC
OWt0l9gTFWew7BdovlLw2+sNFMiYcjlAkDXyTYPfAMc2p0Ja+cq2IVVFtFxf1dEo
tq9xI8tNCo1GyiKzaOavRFK3YAZabBD/XAqOP2uz8yldcc3sXBjxk5zNf2DjiqmR
iNgfbz+o6Yt+iL12l+YCmRfjJX72KtNtVBgvnNZ2pSnG1xKBls+MxDweNKNGe7f3
gCM9GTXzwnVXLsFtrE+hlQgNHANarBajJ+mX5CJWKXwqY0nTR//V2J6zjW7FI5Qr
iptk5ThOolGCKFcgxeq7MlsudprqLqseeIoIO2N9NxiNj/pIb2+yHCC+WNEjwqNh
IL3WAtF0+IMrNWe3AMk+eqGGbe1/jKS+6rn3X+aru4vclFcr5bFdokd+txs+ScRa
hU/YNADnF9tj2qQLWggE1LEbub6yn2k07xpT6CtXfqrUDtQlrXUcIVS4c4R6KINL
0+i07OkjqtI5JAXFkFnRtinuxuBf3CzJ646WJgP8QjfBOU3w2bdh6p5JVt/j4QSi
waQARLBxNL48mPGF56UGRPJLp6FOV+hpHlOcBEjNNxfHyOcAbJJ7mng9g68QbQAD
Rx0La3MzCxEh72h1vVutLBSwHUhf2ytudCI2oRGD8l7kqOav/wgaqmFrKleW9pDF
JZw92JAsUp5K7n8+c+VWnk9XoeV2BD+62mM9c01lGhIUCDzv+Zcn6ypLqeh5qxra
kgs0+ZerSh0QWemgLRlkwTqbt6KvXp/N5d2E54RYhDjMf9KglZMrE4tATSvUgt7f
GyTUZmSeZEK5yez09nZA0cUFOIhmjQeRSNGH58z9xML+hwe6Ra8z0JR6BU8xCQbH
rEpjGHEtje6jgBuh/nB20UQ0dQ+6T95aroSkvdguGneEqEyqo35XyaprljI0uqwK
IJ3qVqnJFar8XjrJoTeNGVfvkI9y7ePt9h4o4W/1fkAtPI1qDYO9WGOTgTEpFCUv
NJW3nKADwsixuINAOU0Yt2ItL36ngFXoFCz3zk3e09sUHU09NUkSe12f9C5zaUOd
4ocpDgqCMrHGbVgaSNQO1Z1hh2mqp6n2sFfUoJgQ9bC2rsoG0HnzABaytLxmjISj
QTpwvd/enl1E/4/RJ00qTXRMzlRxdNPiBd9/KN5yx/zUDeKLDi21aCMbQNjD6o6B
0R+FBBhElouFxFnfkOTCvJDLf7b9qefuR2h656+9P8+dVKxocm2kpbr5u4OcNfuB
VG78ikpOx6382Wi7sZt0I+tAilLTL2jUARP3jpGC/36yXyB8sTODD3ZUJgmuH908
yiBfZJgX5VjOd1zUX1T0IrnL3CV1XRIxKQAh3hnkeYgBh3hTyxGlXCQr2ImIMAtx
8K25kSlzJvDCRtV5efrgZXekIVY8VkSe+HxTKomD6iqovpA93Jikwnk6D416E4+h
gzoEojQtooXZRb6nY8kCxpENI8LS735yvOnXmi2m9WBpjhdoRx0MBrBCaEmsRrpz
WytsH5fJXodQMpV1idACksz+WsmLVfiWmeVigzM0/dcVFOerMPn+Q+XaKkyUOfGl
4KO2fAB7+k3OWFcnmTPXleCFblsz0UWECdd/+BMdlr+hcDDdtqmDLpHcZMo61KvU
qoNycFaSEwprQQHe/94QP3wk7GlJlzWFLSEK4aXgflmq98FRVgKV71ZI6/WMvnWg
LB+KVLFk2IZumgYHAbe+scw9LN6GyIMVFpOBD74svcn42Sdq5igTUsXbbg07FEN+
zmuLpGgXpgTIEfe4lnRwUSXk2Yv36YW1nr3SgplG2yaC0dc2ZvKapLxAMbA5GN5d
d3CBQBjwyMv+5h1hkdYDmtpS//9eryfMmuP4Ddl5GWV8j/IQ+UVDA1mE64zzM+Rr
YSP3/d/6nGcHHVyEf824+c7y/P9DMSJCfV1xTzMsSSzoSKFTxbSUq+mr2evIT27k
KaMtDBhxfMBiFixcutURzRPNDJzSgBr0964kA9PyBM4JVLPyTAwU6T0ILn/bNa5Q
eREzkS/vvn1ChBfezLur6LyRYzxyQ7sBXR28P3l38vTelYwMtWBp1Td5eQ6EbXpM
WE7on/8rjcrs3G/ToVBzMjFG+NwDGQSdpJnzkEH5fLPOmAo6z8D6Lwpae2fRWOFn
owpws7V20bJplqZrHwoRjB8SftW8SUlbSx8/g2KMvB/ElKWh9n5Q3bcONaTzM0SZ
cq2wxbdgigJeP75UfPy7qtolETr3QcH4+foxAItmqR029hKC1va9bMh1bSG5D1E5
IM6qz3PFTcFDwq57EDZiofntyHr5qKFixzeTkv5ZPSa9jmrRyeVlbH8K7ux6DlZ2
jXia4GVkFWZB6UOYOgU12BTmu5kGeQtsHWPoE6E/Upoq/GLu7lnivqrpOPCqk/xC
cD6efQQop4qSiigWZHDI0fLoeUYPqSC9cXfTFKOSG7y0s1afVDsQ27PBpXByKUcY
1UPaKaBdMb0SaHda2dfCOR+X+ORY55lu4eVEQOrqopc77itAbIO2vButLt/2ALyU
mSPTCwlPaBWPHE3k2PTCLS9fUC60agN3ZLrrOKE6KIF4YkRAy83DJTLXscN7oSIZ
0jvhcVBKrUIXb4GCnex8aO5qX16neASmD++aqc7xG8kRnuOqOUOTxP1997KPY/4+
8gu8mYUu2wQJ/0kySc6xaq0efGrXZrJZTxH3oFJvaXJq5LR2aLWJEsOKNnapXST1
oRBWX/OMNbZesEL/L1ouC05wfOsG97pdbjjNANqK53BpLcbpPhxWvd0GoD+kQvrB
4Gy0lazuALetxpgqNC99wciugwzictrpBAwJI+oCi+nf7kQ1nFtaxcNKMV6KGSJ8
f81f0m63Yha7gHQ8My1ZqSba0SvtCd0GCleJ+0bmIOPCUaKxG4U5CM2YOeSC/eqG
5ykH0Y3gYlOgyENJBi+iC5d5EDv1mcTFC9lxpdy+BITRbtuITmVjFeYk710u3gI7
SsR2+7BfOHeFKAUzP51YGOY8kNIpLu24ZPtqcgRNo/rFOEakrB0LNZ8wqogJh3Xe
WeVGfgJ42c/ryaRJ6eIVlexji6XHBV2KRMUJ0NCqt6so54M5cqRfwU8WsOt/RGXS
W79SvXVSquMIzp/BAt3d7+UUZP4JOxPtsMSc0Ko6aU7AvyGkEq5EcA9wWpuUqbPy
bWwZaSmAmo4m55Lz+ZyWVns60WPgQLAdLH5q/oOXcNXBMyokFu2SL1oXYk/KhVw1
R4JCjDH0MEjVQUkRhFdBOZxKFZxG6ljBOndJXQ2WwHRjUpZKbUxT1Q9HRvffc33G
DZlwwxuthBkV7rSb03ULT8BmcdjDZlIZlfKS6FWTqoADEUNFrv5rCPwVRB7bZJ4c
xW9wuanI9ecY2wKTe+vkAvNRq1TZojX1uoYggW9UsQtfaDDuHgxJZU9/gAP6Yku2
KOBGgxxOC6d/FVlZZ/XzxLD7OLIRUTOvGNZYTkg5XwFFZZd+woOXPAHzwG5Ol12i
fE3bLCI2iWee0XUG25ybuDW/IT6fzXN8QtcRfqrHojT5rQ3hlUcqCIl5htKJ2o3t
nQSz7aYiLNR4uhelNrlPtT68siIairSI7u0mzh4vsWB4n04zlTBagl8tC7HECINd
UHJGnEIrdUHoE4P8xW2oXQIlnp/DzulJQlqdbIwuEu+YIzDiVxoEeajWnOs4ZO+L
7Npu/RpuI/e2UNvO2vbHr6CSGukTDcmZD1IJFCjaBVJCp+wnzgq9uu6OJYb0hF7A
SLYmPlFLKe9UK9Bw/vthLInDzYfQcU7tvjl4vtAJ2Qm9zrHLvtP7AVABgkFhnUoK
xt0cyI2KG77lw60tSdMFYI5T2o+ePqpn76Pnk8+mrkkiOXNkHb0E4laEQd0cCxB1
DlgmSo0wGVgy73ZtBvXUqlo9It8OamFYqe7aEAf3+8j0euh+xZKQ71EQ9brbrxxs
sX+jT+06zrhEJQTgG/IwwIKWzOpB0e/+0eQdmGgzUtyoXLfKd8DShVR1y+/1NxVx
iEd74K821O4J0q0hkZ4pnWCz32k6nqiyV75P2bg8WMm1hfLnSt9ujR9ziXxpnWBt
5rKmlYt1xh+EBTrGuzeELuWuqu6kZSasfaRZ4j6SG6lvdgfDRbGJaMn3dzGVXWy4
/1YyZUypecaVnds9xP1iDSoJzfQkAMJZW/+S/ROPZHqkgl4lB0XzlY4ZNDuvfI9n
kTKibBh9OJsy6fI+hEbT37IvMoC72NjiQqYjCWmRKyZdnqbLl24ImnMU3CPx2l6T
vwA970Q3MrtJEIQaXtGSm7HeMBYE+AarkmfLXF2F6a1RhfoEFJksc1Y3lKigTEoC
eCGFP5A8o5Ps9+k8N+c4uZmmD58T5XEkPVjQY8q43J22KnabK9v+IP9BtTIbYOWU
tb4QLDSoNVRhL/+HtpfuJDpMNdVIpnOHPMLknZp0IqkJrWYSooFtbFv3U5J3mjXH
BEhP6JQmJw52YeuRwFcZBK83arpY1bOEEdrOPumMOsJUfH8JcJD2ESTBY0x5iDz1
gzbDPE3M336s+Jyit77mev//sKk9hvpEKbG28irkPWJJXmkqZM/2QETf1zLLMt/o
MRsXs/EzpbnwzOxk5z5L7OB9C6nG1s+93qyn8Uf5rc4Rv+zz+gD8QPXKT1S/frH2
rky/g0AOyZrQA+8g/FfdSt++wRGfLu5+i84fVMcwWynVIBFTsvN2B31pfVboGxao
kA0sasN12hcDAA+aGnjTwXTC8pAxqwm0RzxeCCxke7XxcBQ+1GuSJKC5T2uZVp2s
qCUdUNao+9Rv3uAtVHaq9r25xIxu6s3W+lNi+ZqGVda1honugauesg4tjAxdY7ch
iwpg4VWldAvaihXb63fuzUNK2vkptPzCh3EL3U1kajcUG23treIxrJOD7d4UsCUs
fQXRvBaq+obO6o/uEpIMbmS6b8TchpzHiP9UkR+Ja/NDRoh1nqCcjhFsYtApDJAZ
k2tXyQ7As0j8TiD62kn91pkq6TiE9iBw2vCLA94wejlf3plEXJ4O/FRVceIwrNJ5
R0FM9qHlczFJGY9mviuYExaNsHiSw32Znv2rtiNK5VqhfLSrllyaFs79zZoB6XrJ
Z0tviyIyML17Z5t8csIfCx7U0nrJieVaPYgT+x94qg5MjlUvRFF1TeIiVDHdpJFb
1vPlo50JuapifMejRF73YBuWqKMA8Sv0kp2btAYYFDDB8xPXBD8vCdjLfNtzZS4N
iYmPouKM0wjCQX712sWfHJmk84N27dqZ9t2fxdK8lAl9/Q6x49jKfBpqHABY7L4/
Tqkv8JLq2c8weItKKNvRGXGfShvsJYldEjzqkpvjykSAr7hNL9IUrc/k6/Hled+7
W1ODxJ/9f1HaOqRiSYLkxpnujVs6L0YInVAsnbTC/L0YhmxTBBHVcy9GTDmfTVjn
sYuLqwf9tGilKf+BYPezMVKGZnKCppP0AdOED7v3+mONhgcbvsq9G+QQHDfG44Na
DW030cQd0ur/4kUj4U9MSgjJyyjawy4OG9xFjR8a5DZEMLhzB1nX5eiu6GdDmJS0
Z/nVJVunV98ePyJkNzxMkuVWCZaubK9xpyR2Y5O0YRnceDYTNKwxA8YBIVfEty8T
kyAVq/9DvpqpEaEAdMWJHfYvEk7hN4r7vMZ2K78II7lCgfwRaNKvuKADElgmMamL
9VWehXpFTBUiy4h5HhzZ4MaYStVdKMj/CO+vVAiLKgvsXpUzFmjtZYOqyxkJXCu7
93uB/BlZ4ISbxVfXXYlAdDyVGQSiPtcddFPg+qEWBzOnwtHy0fqA0hhP2XCATfEJ
u/Kc13atxb27MSBplHrYMQwuIiXIjOqDz4Q2sg5JiBff1nSpT90h4QAVtKROHwbD
5xVSWuvVGpwrR4eQtDemeTpuyB+ExTOi1rAnfXWen0NvrvnVAEEh7btktPQ+se+W
VyXztjNJVZSbNnkKvoY9FrJyeTa0cB5cKYAaD0+GgBIwQcEUvaHl7n0fFVc/2owr
MHxW85tSNqqB45/9WIFeVk4bJ9uCD9xoD4JIoIey0llv3JF1fdzBDGvv8Ke2Uqx+
4J1d6Oocg1QdG+m7PjZzuOSEaxEJLlCe+VP/i8l78oD7DLfdIKpjBP1KEbaj0WpR
1lpT2OWwPyeGwMEkhCiQM8V3JQjKbHDgBZrAZgFNFdK5lmZjZRq+WZXZfOxEBBzZ
8bCXFC0B0gd99WjO/gAxX2aJEHX89pwFzn+CWzXM1XDxT8LvzfJD5wRZc9aroZDs
ZgURG+KbnYC06iWlq1s+vBPfDewzn44OasuVintXuGxV5iR/Prqq4xAa6L8fmP0W
kgcYNoxpE1TSisAgbVTWE8Z5SZDX1nPxvnDQrnV9feFZ2xrrbUZ+AhnRnxeau2oy
ZtYSpPDtYnK3UY9w/TCXh5/bXcC3zx+YzBxVGK+igpcQFtIv7k22gyBePI0SyspE
pMBhYYZ5leH90QIW+wNNmG9fTDSuOQrzvLqfrT5tiQAxZWNHQaEH0tX2COXitr2Y
4/tQ2ilIgn9MhwxVvNYmOmxeXitl5hLmP8nYI5Hog2h8w1iywUOsI6IdE5vPxh8L
EQQbz7PMQp9PbIQiIkMsWy/C0238SQnIwiqzKQKwJbEdZFUHJ9XlNRN2MD7/zRv7
YD6GGaY9Wtkqa+zomCHoaLskRpu6xkwYV8hRBlGQzPCdlA5jzgJJtxwuNTqmY7OD
acfhiR0IUmxS4Qqc3Piwk3scx8fimmhswdh20GyA+u5aYN1uut9Deh6BueeNFkxR
0LCSsa8Q21bcl04c4Er1m+yECSLXkSX5nrSlaN8NSMHbpRn3zDJKoi67UtdTQGkO
vZ3rWnkmywvWpxzjllsb/6JK0pQ8bbkyJ4fBNLqZeowrS498pONruR3FW1WZR5be
BWdrAIRa/cYaFa8j8TAWWcX1+K6fM8swX8Sn/4bTYiWcR+LuUYDGnugTyiOjRUwi
BrkNUVZIBRaU8mzHe2MIczeFrVlJUAj+tsz1V62Cj/VIvpWSPZ7Se300eybAtn5j
zes3myiJawKEnfyyEyXvuVJVZ351gpq3OOgkSr79rcRJVhJ/I3oKB8jQKXuwsqjb
nuwMXRCnqDzLojxEjFB93XDS1GbloqIBEICCAaKJw/ckislAGx/Y31ExkriROUrH
4tL/Mt2T6tA+VFyCeU1GiiHtlSlpHvK6tx49zB5LBUFFYIZiQ0Lgv/wXf1QaMtCZ
+ZLSMz8ExOymUXr75LezrRtLIbf0OAEHrvoKvEGomVgWyU71hySWoxR8MRrpGT+1
I9Jvg/7DEhUMbRrrQu2vEBvsOStq8Y0uA/FS7Ym+VBHV1aT3M36LlU3Mjj/N/PjB
48hBUqDB9Cmh+tdJqDEpy/bmjJS9jMOTtKMdep5fINsx8Jxm0wmBuFR45rkaA2pL
gUqa1eWHksdzci2T8loSZhIZ5Gm9H/gmaResjyRzmGg6daZxJwGqj8LCYJx7/7tQ
oXm99UMPUf8u1g9gquXmh0OfxYuQP8vrIScSNO/dXMDlvlhlf5xXoP5OVZXZ6rwP
5jz3PKfTo+efXh0tVyLpv7+C9rc6ArGSbeEBtD8rJovfVA6mlhEJ02fuT6pMfowb
yRuVGY6qW9JUjuteDf9x22b3uHbthlOGctRFpTte4MUzj7QlVF81vSPaVxdKpnxG
kZLQ/mQUuCd7GGqzdJ4HR517UL12hs+qAHOydiKkgH/FZGDTwlXX5hPSfll4HtFe
cZwGQIw6mn6ThjMyAbOxCLlq/taW8gFpKAHC4X7CnbQHm64OLluYltEGSjTstbeX
HDRvqRhP1ufUVtpcv/7B6Ij3QY0cjgO/U03S1BvTumCXZ20M8SkahBCcAyskLor4
1Oo/zK23mGWR6gWr24qpQIhYiOerp8hOq7MUwdQk6yqzWKBS71eDZiX4svQiz7xA
JS47Qk23xdr7oZCnaIszqv8nNBuYi6VQ/Yekk7IET7j9Q74KPJVDDfmw3Az5Tfiq
SdvbEa1w48e+05gg4j6TNUF4b7YrHgNhspEUg5a+bzgwLL3MwjQfSCcilQv5XBhE
1zmNZDTasSFs41dY4nB6se4Nb+q59aGglP9jqU2+zruUhbS/2eLiu6csyFKZ/e+l
k4eB+IEJlsCjnl9Ly0BttOXAgsPEezpFE9H+hV4PplrsodODeHD2nptDNQl3WMyW
Jy/IPpcV1Xzo/DaLQZv/V3zdgUK2eQgMAbkfq81BHqRB9GSezyL9K1tHgSpLwhia
rX3D+6uERNPYV3/JGF4p9Sdi9TLL8XtAIivdacQxrcNs17KgFuXnIqYDRC/u8C8J
09TnKCWaS4w+qgwh5uurJbwPNxV3ITetAzOPc1OdGSvpqcsuPfJTffTdxKR4qNIL
OEhK/cxNOqvoOojn++fW1hquxGgg/StdryVLjhYX+7CqmfbSyPdraHb6oWGHK0ZM
bZ6PsPcNmRlKLaFPSXfbQ9jYLmD76PIBqjZ50oJSkjymQ+cCAd5ZsEn8Und9RQY2
zVto2mvH6ZkJ8XRDHsYjUzXamzoqWlidtcCMSAmy91bX8UQM6UVbhJ5EwSfY7OnY
GMPnSZNyu8ZdfJe6J+utFEdUwFYpZhNt5RG9lmsziQ+uRPGamQCiPw9mbXULJTG/
VHKBYhVx/RuFKORmfAm944GWPBw6NBepjlyhjQHWoVgMNh6l0X5PhiMN3zW+lix1
r6ULDTVslS6+DHgTZ06CQwZteBRGyCazNphWSeYVPVaVFsW83FF9IXrC66YA4NJ+
AHwm7kRdHMac1H5RGeOlZgIfseUCBqg4UieM0WlMZ2uJElzRU1NisXul3kGPiuY8
QF1TDL2gQsXtI54T9KEEe0pCjuXoQCJuJjWh571PUOTw+jHUjhpMYvfN8DVLzTHO
oSXvYUOhWYKEgBNakRVcJyYnwufRphzg3zbp9lCyND+75umrLC33yEFMZG3tjQEF
cxkvhHopjlE12MBELSJQrMbrV/E/eyhRuDi82M2A98kZMkbm6hKnGVfld4HfPZKR
1foBBbdXh4eY6hz2wyqdOzhFtSXR+u10VRwmBZP19NMjLsg/stSHMNtEesrmZOBu
tfweqkMjkGGC3bHuLX7ghxyPhmAEsHwcGdmzb75XXMmZFEcN+52gI8jHX86Z6D1k
0d0SXeLvZZic3I1Ep/JdmkarBxU05NyCcqgvNnOlUBlczangkIo6ZukDdo6b4YmJ
G1LZTI3/yTqkOO3N4YueUF7HzkT51KRoSEZkcM6R8zzSnN/is3eJtIdJDhGfWIZS
7z9DkpoflhoX3JblPxALT9ie7pwJP3VXKJ1p6XMqSxlH+ZXmtQhbju0eZ5hndBpj
Pka2cFQTL4XpqgqeoykS3Vj+Gtuc3pESD81sn61Ce1hpnuYrMehtUQjLdxDmP/tN
MAuLauqXuZ3HsdkJbHiY2Xk9ZW0adIJruxo69wJnLJBL6qZtvHO619O4gfz5Jgr4
AtIafsTfe84APKb3zkR3jphmbn3Xt75N7TyUQ/Og1PmhoJoqaxyxIHpxnQgMdep2
6+fH8lD8ULJqVtb8Y+Y8xqkAwqe5Fkff3pb1OECFyw00CTbbsiH5Ah7FiqxXkefE
DHoV4olu+P6El+dqkUL3oik8EmfFLzX0AoSRjmBFQgtuuoBasp/SrtftkiJQL1Af
/Gz13Gp+3nsqnzv9Yy9aZPfkSEty1ta0/ZhELpeItVinfygCkGriwGGJNiqqYud5
v6OnHuNzA62QrYUvSIwOwhLN6oj/Uu0QSIh/MANbSYIZsivII6jOoxfYQI1GIjvS
3AhExylrTwKuyHzCaPA5bC3rbxzcY1/yMdWC9GVBYUsUpDxZUsvEIdqC87MULS+H
UytgNXB5Vs87yhvUKKNlXDvFQ+vUFUDenjzaTRsghrqo9u9BdQCl6mnZxddpUIyc
r8y19o5xn831+OfFMTKyNH/fGKm7xIcb4LNOGCV7I76eWuKvGVSIXMf3tY1IpvQy
aCijHo+Om0JIuWGd6e2mB2xqk1IyW2iQWyvwgJfRmEEVC+Mvzyl0bfYse7lIDpPJ
Pwv4oS4x9+kCc9xnX/W9pfjMttjBk7CCKimS7eEfqRlusuPOwzLO989Lh5OLNwDv
+vh+H8jLH1EWS9Z/pp4Sf2bH+eiVQaeNTW0OrN2zGxcp3cnF1Bo2rpJIeNNLRKcV
WdBo/uyh0jqoGLOjfRJlLv+Qaav7W+0npTyscU4qYnHxkTdfxOxPO/NBxJvMvtdR
/6k9UcH91JOCmNhds+ZiR8OrdtQ96MHPCgW2Fuq3JHX157Tpav+OUFz3xf6OSuz+
LOpFuATLtv5dGyGLUnCljg9rtiVHF9Owtmg7wwS7vDuphTpqGEa09VNgOlwa8iix
9J8Q7ylTOD8V6EpyvCAnPkYZ4/8mHILbf3rfefq8R/ARq1wNI8sbIyZM9HIdi1I5
dpu/md01DNscaauySOT7vbMqlcb39yrzYEDwF4hGbdkFniRgkWOPtq7ctDxVq7z8
Lq1o6UtOf+2/liZfYng2164eng8c7Zcz40+pWnX4g+MlTFKGohokxELPPmw9nsVm
tWrRoXh+pPfYu/CyPJUpibMj9ywyGpSRb53EoVnptyh445vSG/oOL7qFbdxBvUdS
ddeQBZh17znl986fgtODJdOQGuhC4D8j+Rh+eV1L+aabgTR35N9Gn06kcZNqL6m9
0DD0h3amu3Le9zBqNUMaeFHoIZgBv57xR7JRVHbMkJ9KE2ZeQjpJF0rh/fHtAGQ8
i5Heb3k+wJu33VM3YgKumy2so+4pGQTX33etdf156xlYuYLfgMp0XtGI9FnRp93w
sY7K0iaefN/FasqnUhky7Kb2U+rrXwGP4OKb+BqhmB6ZcD0UWh5BpCje7KJfa+a4
mNxnQUUbsZ/bdjdNOq3qlUk9y7WzNu4g57YbfcuqZ9/H/AyOgA5znsr0wcRaC420
z7KuR5jgoKzBF/v3yM7OzyxPBz8z5IPAlLw8WRiZ9rWxXvLRr7Pp7nGp6boQeXvp
4olmcnwm4ZmUXMbIOc/uXmVNovrYyc/iU8WMkp7ZFmlvR66tAeun1EFxkKuGh3Ve
dkZTx6u/EgvORoruHorOITecAdUmaibl+g+91B5fnIktgw0Ox8SHqw10iWGqXETm
kiQUkBZBdNoBsye64dc6hxNZbNuUxENzbSJsbMLPzwMP+epgvI3vJK20dSmcwGak
cb0evuLrRS5GGXKNa/092YqTvUNtfnkXIwOtOqIgeMpIZim0t4FeY0meXMPFYx+N
8zep6kuTloEfX+XfOScNBhb7c4UVhMkr2x8BfIEt1o3xIvNjG2hJtV5/z6wDojT0
vZSEuZSi5yLAL7YJhYw17MbBTAAwRBoETDIfyFrXoXVdcIAlfprES8J47TBnr+3T
bBt29opwyeNTSk1D9jwTxaNAB5eiV4iBei9yY/K/GoyPD+Y8qy31HSP+4BBNgVzA
W7EFzGdpuhG28d84afz8HfEW4v+8E551m5fsEbBYgXTXeNDJR2RPKM7EGU4buTY6
GguH00A2dwfz+kzD0WRdJ/7shv6f12WlojeAWY89cuZEaJko3vzd6CeYt3oA6a96
FRhXeAeowjYWhgYOWxqb3yWd9E1pvkYBiDKhKIa647l4agH+pNXqoNU4ajaUhQMW
34iiwtfbyMJ+vvBK1T1Oiwg0AB9lH3SCG0nODIUG2k9domLdBrdkS1jdztnICiYJ
i/biqg1TN02xvXhwOC+yRd2YPC4XupHGq1Px1jFudbuTw9rnZ3zlUrhGp4+XjRDf
0XT9MPQG1KhPkmFJiU5oyW5TCOrJKwURUzNimHPBovndFP3Q/CbxBa4z+TUPfk4U
Pu6G2D1lyNII41+8JEtt1+nBQd4TsSxx3YkMNPGSLzhahGYST980EmZRGw1tt50y
8rjNrRzLaeTrkFxbUzSwzPFiHOfLTaPZaC3sGxrxBZdjl3OAppVdpg8GtUrfxU37
LrfJSVbvCEeN5ZZCZYxl5f7a9BE9X72EB1p9jogmTVZjD72x3MzHIbWurjCyypDm
HvZFRKIJ1IOInKAXy69TqsBnTkpY934mfjfnQaGmOytyiiN+adcneRkuEXkva2um
xYOll0EhpGHb0UGi1HWqXrLIa7Ev2/AeIy6gh6MeqGMNLXkMruCBrHdy9oh0+7Ud
1obWW5aFGefAGZBE4KD98/8jhowhXyeMjZjF5Hpk4x5/AvZALqqaahI+gSfOtEUZ
Zux0Y/krHdZ23fEmi2pqaANlxc6ZYpZBVtW1dEWAaPBqLLEW/0gIlQyxDGFOzZCL
NHJZEyp1NmLYGvuwlBpWIze5jX7xXRoC5ddYwn/CnYSv/Le1IC1BJLNBauhuNuHI
HGGE/uoY0DJZo1O3I7XDpnb8brwYNDuqhaNtpmlNIh4WN6xWn4z5NwJIyqA7GRFl
MezWiYlWAVzQ4XZZUicnPVRvejVNjBzc39U0XLnGXqK70SZe/F2rFSfk4wa7l4iC
nl/UMKTlPCNJRYeCHegsXi/2SOadFZNvDlBN1iXSlvnHQEtg0IbzlrfEcWzB5xpM
tU4TQSVSt0yaGVYB5HlDL3wC4519h/gMXq8QLgkQpXMb8c1/OdkwMPwG02+nTFQh
yQwpv7p9Zu/xuaeOEj41HvN+gYvyFQ1QP0lBLtDo/njx1exMGfWyQBZzQgwKQSpy
3X9ndRWOfZbBWgDbGbHTNqxdS++Xd60g+Rt7mBs2IusA0nWuk3ap7aX/M+rqFPFS
H21F8ARcrLwWVy4LtKHBax4dQb7lxykW/gDKQW1Rgqdbd8uKGXq6tsilV+68Zs/P
cfGLvwFcdhQC00MsRdxr8idsxiPPrHFKhg0TCl7rwdMaa6m2uwaz9LJTzbvAuNvL
0i0lJb0L/m5kYJV3/GuOT2mFX8fxTFKD+ojXUqi30V4n8bi7GCC9Cuwlnc545g0q
T6u6XWOarynCIcGQQ7waauu5qezO7XaUyvj/gRjg8USfJQ7pN8ds20JxEKK8bgqJ
d3XWlI6TkmBxb4pp/yNUdjtxIU6STM4bJ+plW9VLkpvTJBO8Y0u1kjRnt+1N0GYI
y1NVc5qpIYD7xCghnTRu5FuTN0mCINlN4mujN48q/V8M96VgNcKYHjKo2x2HZfUA
WL6Y1x0jeDKToEdthI9j5Bhk74Fyt8eGZHi67y5z+MH6rUK7k2Je572VA5/mxdn1
JKTz0z3oOkgTrF93BGsA6Ew/K6St/8V7p8N0zwcBrJAaDn7VBxMPrZnKlpW6CRf1
5jCgY15yCTVioYYaX9FUWMZ9pxLf9QhJW1lyWySwiTWDLneqTCRbrQPsRh5Frsqp
Hu/rXLUroYBlyfd7icse6GkctQ9yLvdcx4zR3WfV2a8Aa9Y2q877SnxR1w3F6n25
3IdbGMQC8ECb7PfiaMz6F1zdggB+zkrQLStoPOg52vWgI9+7BWiAsJ3n96XsRsiA
eYJw606xxU0YE6sUlBjpwuPxcdDWNfP1a34dlg746Yxa249D+CeXh63/MTE8Csm9
sYdSAA/uWT5HFc1wMFPhBaIxnM51Vvdd317hdHHtIc4O5g+IIiIT8iL1ptDtgqRV
SdiOxbaGRjW7TUWh3eYGBdCV4c3XIPcYA2h+EuT7oJcrKvtWNwVD3adYKB3KyMqn
wm2E9/F2qgKsQyZMnkHmvWQDpSL270KgbBTSVE1+KesvKtvReV4of48re+t/F66H
KQ90C4H4+GWW5Jsg8RyHk+mDdhCyLRFcLTvhkHTlQozRZjlP90zmZwSAmmVYIsVx
D3MZgwJRXHGkW/SUCBEDy2a3WyfVBs2jJrMYwj3j5nB04aGaxkIG6H8t0kmiYIZs
Pq+aCbLIDnT9P9613bQ39xkCokAy7isXs/rQ21d8yXRMmeuWI+ghfW7ewF4AAcao
fmq330+gS7eKxu6CwyQMHh9FZFUXb7PYk+HP/Cq+2w4ciispV0YShKNKFXvAtgM/
7LmmoAWxaFJ3PLYjlUEeOSYIsQXfPzelzHJt/tcZZLW+rJ4+L8MDNQER3icu1r+K
3CZ5K6M6ZjXUybI5sRblfGq0jxBOfVzqbaWyJ38s3rJ3J66rVj1OPs3u3HqH9+h9
suffYZRCnxb+zbgfnAK7/LUNJY59fwrmIdjaygkNrji+Zp3m5PZXpE1kFYXZxsGQ
QtCm8FWFctFH0kZlE/bah1psQ3vducvJGa8EodOIfo6jVuf4XcSCy3011w47XmYy
CsEyeno9sv4Pj7B1gBsR1FhkHxu1V7OV7MQeYiftAxxZWNqD4kiNthQc72J71THk
ddnL6+WLV2bf4dV+PG+PV4ZyLk/o60aE7QYDhUvPzLdpcIqg1/VII6kRZdOXvLtJ
wqmv4v/ZlszPGOS+YXv4HCdawt9rwKxX+ud72iJ9zweaPDHE26eaq8ANW3VLx+fy
X1w6QxKw8JIbxr0lPgZGtbUGE/I4puTk+oBxvMAF4MApbiARtjR7SiY9dE+WNUSs
IMNtufSjqEFM76MRKS3mUZViCT8CjcQ9M10D55iFB4SjkMHogO/0UO2UHUeQ+J54
SGSTfE5w5SoW0n770XoIb8ate9FC+WSQaGqehMKQs16ViS+I00dGzJg0ZjZ33e43
t8APznrHaPjntTHWo+6j6WTWg29pbHIVfK7UU1nGbiaKXkZFpmMIEF8E0zvHo6P5
blRopj5swa7dOm+VQouKEDfhDpPnTh0V+UaZXe+3eIreSp4gYOl9M4JUNEvzk66D
9fvdIEeJ5FJGsTuXd9+cPkbObTYtOShcpYC39AbeiHedLG7Eq5LpLseAXLCS+lR5
+aekw5U2KLeWd2bqjyo33LZ5FWka40w3XauFkeA78pb5yj23Ar+t6icTVslKYvvI
r9w2aHLfUaHHaD6lF1G0VcHYATK0JrnRzAn509Nr/liO3bJhh4wgwAmaOL+RsknC
6A4/UrlmQ4Em2USoVWEASgn4gfbM+eN3SjWiZKgOaQtsagDS1fzzsYGSHnoapBQ1
0kxnT9UjL13jAUjBnm7/ogkSvY9PI7bDnoSvrrzXrLbXqQXbw4ZmDiAcNtj0gBZy
lVjBI5qQJneIAomBVH59WzygGPaP1YUAqzEJZ91IxHeOFiOh2zOv7VaDebVTLk1R
8f+uzhVexI2wc70wVqFg6keu0UZEbE/i1VMPC3+o7fshqvqnhqmWCQ1xVDNURA+l
NfW8Z2KJTJkED2xfzcD2UJYuiP9OOoV+k96XeQtFsXlHQXW4ay0OTzc8qV+/iJE/
3X3qZd48e57QTzp4RXjENJIa8YA3DtDkDV8P27wJTlCr3Pt54hTIzOvK+UsfdDZH
/u+AUtsjLXyBQ08Rh1AYvwehQht+MXPOGUvLAAWYPEZl/orInRmIlq3sx5pwfG3t
/iu53XFLD2pHhvOCSWH0iGy09O01HEFBikv6kXr4QImBMMJiQZpD1kiFsrbuUyP7
l8f1SGK7SYEDy73qzGbTJtqk+3OhB+IEZwJGSiF4zjqazFL6OwgByDI1CYCsPBPo
gXSj5IiO3WChJHOQYdNUmTpUNmkrcgK5tp4qlPKFhneybDbnSGg2dMDi6/po45kD
gHDPHU1ZCvrvvU7+zzvUqtz62lPY2GGnrevFx3t4Q3GSzPchcncefcoTvhtbuDES
aPY1bZ7wq5oKyRFSf/j9ipyJjkEgRoswkFGwkLruI7OuPyqfVZJbUZRj9BPUeAUg
gEieSyi/7ajkCu/7V23Jt92dcIxMFPkzyth02JDPM0h421oNkPRuj1h49+q/7mD7
2xsNGDJeTIIIC4XXxSbgCDmYXin/EBkwQIYxijDVdCfsy6AEP1RxBX/nl7KxRhWi
J6AfscmQcZeEPdndFDM0z3GUyLv3hy4FhmYZhuRYekfpmiztEABi0MBKP7jqUw5p
nKDvwQLUoFHA6zsZnghPQCZiCHd4NyOTqXxbi9tB8bKFzwchQJZUeKwtBwzgScfx
rhHbD13ZeUP2cTDWXKig8lH4Swx/cFeQdEwBIGyzqEcHaaoFTfTElbJIJYfFGQjN
uU+ZueMMcKrEohdfAsQMbdg0JG/6WEMJBjXTBPStXV52wGlvNZiiMILnowdqys5E
sB5azrNJ18awQs0HGjonxttShsc0WtDV9h5Lu5fgqr2IrB+G+1Zt4SVIzBClzgA1
GaRFAf6KjkeKtT1+7NYPyFWvXBmIzxJ/JQlqpPqA2qHDAuePIy/g2XDTC9h9+6Xk
PD3AP+1hK9V8ct8eHQ/5HRWY1LsVtOKSL7cbAZR2oflixxLEZOb3D0HBat51wZDi
5egPVz2uwF93EzEiFsE7xFJLF5LOdBBDCcz9+Ufwl1zo1wFWZZ1c+9qsvfsnP7gT
kAb4SAFXwLw5Ws2fdT+bD3Hkgjq9rgg3CzHuR/EGalehsUEt5P54cTi9Qfe8c+rD
7gRwhPtq7y0b1vQT2LBUPCqKyABO+lLztDNz5t869jc33XSVkdDQA0fJ9WVcGMoo
h3kwvOzrgXBVcPQMLmK4oEThh6i85jdXpGfK3zsh//ztAWZqnx4lGbj537fkT/J1
nkHAw+6+lJeCzDt0R3mEqoLxESvRe+k+DXXdXxVVND6UGHbTo56+jGedGGNWvAB2
BkU0J1mUpzr0Nqwef9fjas/8/RlAbT3pNo1fOQ5aW+QIl1mMvEfSF7Lx/LxQmCmK
ST7LzPyT6XGpO5CA5aR7/aqT//TOE69Vt0imrJK+ngP79OlaBXtYpvkldhwvYw5R
53jdpVYIam/9DIG/2jNO5BMbtaFXxrPBEecbw+EoBxDwX75o3qLR/p0ep3yNRCwb
fMZ31JAvE9Zxawq4NlJNoakzqbFETYT3aeqNs0rp7mGRbK/Ww63Tun6l3oFxXrve
O4GHO7tBOjKvGf7+np5HDLXiyZKry/DwIGeQQqAVSjiExXH/OajiUR7vmbFdjS9/
aT2tcnKvrBumhUYLOezgaHQa+TKj1d6ZEpQSRzvH6Tvkmdy8H6FMPQzkbRr93Q42
RI4OGZ1DYyJ3vbBur02bmNVOKyp+CDdnmDBvaZF81Ow7MxsDmGmUjQyWIsZyk0C2
6XPJicjFaYM+TsxQzM3v1WCl8/GimeLnz0sX4bnVhYrFemDD72jAexMVBxIV1jka
5MW68EWBhWsDLZDv1tGkGWv5fTv1T0kb68LrJJC9pHsWJKgJz7sV6n3U9swmJmUx
nkMYG3KQeAXj/hD0y+BF+bOhYWLg7Ta/zaF94LEwympK86MnfY+IE3XJw7aygPi8
Ic6I4V3xJnlkx+XdNTH2O159H6JKQ5DQoLG7P9ZnKjoXnGLBM9PEgyz5eAfId/Ll
f285PcQmDX2MbgXGyXf/ECWJf6mOYgrj413nw3LU7acifLJmyeUiRTTNjwTy0NRJ
H0Y0kIt23GTlUMgkvFaRdmHmys+KbjALHAhI5Z9lokNvszSFx/p2UlQl4X1s/NO9
pktVIXzcsqPrGHwZmq1XcwwYn6hLpbe5jeBnPPItbw6ek5qp8paObyp2gJDtePwX
/XobNZRa0xswdrKFJincadf0RgMtH/Np7PYomeI1W4CKD5Ebv6rj+ojMvAW7XiZO
AO71BNpmxeqjdHEf6vAF1btHSpcqiLkjainxpIptdiFo+VQZoZX/ZfnqtKWfyycS
ZAogVzNFR9mcAcVqeAj8MkpgtuLY8iGU7OpnZ23JUfupEEzyKTBQbySsl4ubWB78
XebnZJBWSY8Ltjf56hquUUamjR/oR9k10SgR/4dRL5xwdnSs7lLcnhh8mP0hdaWH
PBaVEIxePk3ACpBO1E2wUITXFs6JrfTAFCURTz+u7S6nBNheMt4J2c8H2af542NM
HTOKPtQQW9zxPGtPopXW3LQTyAm26HU2rg2sB3MP8mkZPtkkA6vRWXktwRReUJfD
Gu3d44imNHhACAacs+qlZiVuwFlHw3LmEVcsR/WTpYDAwIXrVQhIDU38GboY/5rK
HJYf0Q2cFCFXBU23Xwpo0wX8FoIlCD4eNBcj4JScvZMqgt6txSn6Cc7xCiFe7Ujy
A2+dxJZOJM6GtBDVsbl7uEnnt3zEj2ymmB8H/uPhWjYXTP+IZH7Keu/OuxZIUo0H
4YLXmDTYfbU9lOyOjVCG88lyOi7XcffuCyDtjr2wUJSObWGmC4d+Cj5QQgXALNhk
ojqCKjZQj12LzYWA8MVudYKl74OBefggkXsWtEhrvjGH5UHIS1XHbwrQ33Clk487
3xw+nO9dl1qgWNgIDOxQ48hW4v4TToWoTKvC1Ezgg5xn7WR7mUSnFvsprOpkk546
1Cdoy8OFsIAitRuFWZpzp+7qaYJ+JV8opP1fGAlxWg1m0pm+18msHySiMiGAN+1o
TOi6RLvyY3O8XZMLcLdedPDEpqEthk5tMk4uRCX4o77VwNwExr7p0948OuPsYb8v
jnv7kDjZTyj36YzL5M3F0Jt8YVCEi7dW4ZQoyVY8f4dIrUU0XDro9CWMtlXQKKj8
rD0/VPjksDywWY1Jx88kaYuU8QKd2vNpJBMYmTBTG9AVGyDAxFqwoXYDShFRZNUD
X8x6iYlzKuHBeCEt5md4VBkczA2vUpQnDtzsise84MibGLbf2n/r/eLqe71Ld7i7
2yKdM1qX7rYpzKOAgyekjtoBC/4Jp0kej1MyVvuiMr0U8EjNaWqgTiyc6BCEZAP8
F/8j/aG0ZVVeKvG4pWDYSiWDbLndezlGPhbSVolNMJ5Zb/peP2jxpKzWi1iV7XoX
+RyZAaETp7SGRHMFmHD1R4b/AflSHOwLzixocRxJFR3WJUGbgHwP1+2qld/VR9Oz
4tEjoEcCa0nKTLNEZT2E5/AlliNJ/2YlWNCcBncFtz+EEwKL9YCttCMqtJAp1i95
A/eIY1S4TUaQyIPZSc3G4HG/GqDzeN2z5Y1EOVOa1csveJ52Zp6ChsMP5NtEt4a8
QGLRfAMTdhtHeW3/uEd5YBYxCOad26ld6vb6V8WNtPmDSFhnmpMlW3c++IAKB/66
KeY70tLSkePWD6ObajcVoBtJ+sLL3tfm2hmM+ziarLE3k9xsH3Am2vuNJBnl9ic+
ZX7PRzlnW+TwjxZjBpPceHZI6dJ2HDcrjs2ZkbQ92CUqWWeeppPobMELUBn9rvGM
C3befKtVdM+DPBOuU9WeXFJIKO/pEUr0KRmeCwLn4IkXVoPo8jnHjuUW1NkGFLJQ
MI8n0cP65hTfGiJ+nygDHTyTOzxZMlOMmleDDV9Yv9Wp1SpzsGw8Vpq06BPAhH2t
MNQqWUnL7rLSa1Dmc57oxPYwCqHPzgf+vyN7eKR1+kL8jME+LEOQSgmfzb9g95FT
hgPOXfVpYmVpoSE81+no3AeUo3dsBs7GLEn0qBVpIEXdRk8n2IIB/RUwAYjUhZTQ
YkOpp4vjqgDg424+MIZxlBkTuJ/nPbvAOautTsb/sKd+lWNjW4pQt6X0K2cOsKEe
bNIf24FRzs7Upsypc+XfGLSxC3I6GeJgaEbX1gAU/nJYtDFPJn55tEzpCHG4tyRV
RLLw4WRweadWTKJ/di4rLwC0iU8/jOVj1y8QnberAnM3ZMR9eC4UCLbDSI/o5Qgk
UAC8jvlSNNSgHGmunc6jCfGmlSY7ccPHEVT2HTOBM8ZFAqKYFpUUoGRtXsoqbQF5
uRwVYOUK/+KXz2UiN2T4UJ2ZKG3Lhw875O6c1rl9vAv/ilrMNOzqH17CGLdfdXJ/
LZLBlAVMZxuqgVA3Mkr9jAE8JuP0JQ+OTVR5eo2kjAYvy/R0vA28VHR7pzBX/Gi7
LAwC39ZZ+qe8we68QWIL9vaeYGw3psNZPU3k9VwrxEn8GaW/CtcFwQvbA/Q7CaXh
fDn+JlnoL7geEoOpzIgavS2c2Zj0JKLAr4cou64AbfG2hQvWgWBHNS4hxn1jK3x+
EfnsuTb1NpG6exImiv8tlZCrCf8aTxwCUkE6nj3bOmwoaoi6/NbdMkXSANtuJ+4p
L9Zuq0Ut67jIjpnAgKTZauJqK5uaFppVT/cuBAFjhCGz7phAZORkNVAK/WUGnki/
w5DzgZ4ZDvy5+C8Qt5jzuVeyreYJy0kFw6N0TznnK0GvJ2t6Bkbnhx3hFxJPX6iD
J43Yn+n6a/fomEhCOET88bNVWqBU0cNKHOPtTz/n02Z/EHbzkHeqcrw27LbIiSeS
z9n+fe/EnhFfrFy206wfm9OdWJsK+3sb4FYR95jHUitRVLl/5/YW9jFiSGbypt9i
0auDkoJROLhUy1NWb/FJZOR9Vt+wkIpF+fe/hu1QhGqSKew+wC9Ew2v+Ssxyn7WQ
Jo2UUIeYOkHKXEzE5IrF1mMbzOLY8kkPlufBiIAy+nzaohlwuG1FmevvL8zWusFI
TAVoliDIREQure0/N2mDQhYjqMQ/vHCY92DgXhHNOJgHFVIyA5dAdWfcN/3PZiuC
FgGF2UJtlE7syrflnxC/8nhD0I+TxwZgVNIwHJ3QUCrhvFapi0fqisg7riOeRqFs
i/OzSFyQl1r0ReZN8dkjhE1GeHtZhqGy3Oe5rQuYFjrv89tkAuxMyjkv9ATzzX+p
Ia8afRpPd4alFJBubzMvyQfe7PD8SQ8WrlvYGALkA3ThKtIOMO4RjikXuoYIgnAf
2W1Uir501jhyIFJOssrsNXutgkMvg7a4pVJrbLQqCE01BHUW+/k7O0hEmlumGDFY
yM5vIq8/AprNT6Ly/42CJIbSbCHm3DkYWEvSzWdOSFasm3LysLHN7UNflHwl23p7
oi5VMnSRQcINI5orh9UmjESqZxgcFcVfkRfhAzJn0ZiU65/hxSG4AGKL88Qnb+JF
o+yjxufy7zlllFlVR4YsoTG9RUqXXW06wyLvhxNjCPOQYhexPig453fkvI6vNr0l
7ojpxGJIdUy5JNqhZFlBLlvcUIbeH82t2CuY3OedNJzzDBIqfjLKdYnBFAIJunZ1
5qChf+z8vcds41AJJv+FBJIz63ZOqN6lWCw0kLiWPe7kZSTWixhDgMTvVa5ZEgH3
WVWmRnPx/ijX2DMsox/knU0vN++rbfxuFA93oq+Yk5+ESaVLzeMDI303OEj4Unii
HES1K+yMIcFAGEb3HiDJb2OEaugYE003NgqumrIr8cnCzWyoJATwkwJUQY44Q4zh
/RpaKGWIex4j+9T8zY+XQ4/8y18Rapg9/Bm+CVmN33fuC94FJJeIfVQg4CbSaF6/
WSxOdqSQ7D8+SzqzMHc9RHIbKU5/Qacl7vlJVkn63W97fhbtTUaj8HVbqJhPug81
ATkIHOMgWooKAiaz7oW4C81C7EZ6JtuzxM9tCvPrEn0MKS4SxUjMCfK3c04oHdCk
oaI6dOxiNByXKTspSqPgx1Fg2B61CLPEfgtiOkYIcTIY1O8WU5XXT0Uc3amF7L/o
+dUj2DeX4jIcLhksQuLAO9Zjs7eyhHyS50Q+dDxm7ViFVa/Ms6LpnPiuEttZ0hVq
ZfwAMOcTttNU5ds+t0feTi35mmzyAv9/EWcpQV5QK5uWPgfy70ozXCJW2CVXSOMK
S+W0cLJSkbFNjqeOiVl5y5R1zcNGvGz3NJNciI2Pl6Hoa5KqCgOtm/i58GQPGN5F
BtukVUZjHGhEQRk4N+wJX2AnqDsqs91T5fb2Z7mt0dUnkobHZuiuCvPdKUhm5nUc
0+fGq4f3z0Z6vR/1T2PjDyW+7noZ3cK5zRvckAshIhnCC2VuT2ZifWQS6CLolDXr
emoUUKfXSU+RhubryIH/7dfQBmuFfEDfPg2QSMN37ct7QKdGLCMfcNytNHWuzRAU
JDJjtYvuUO1rYBtcvUmV4q59UMvZsaDMwU9IYMeu//JOkesmjc5h8dXrOes29QIJ
bCpWjdBL/U3vR3MQSRDzLtMYhKLmv2UCV15Wik1FVFCbqc/xfpinMw+GgwOJItfp
Nc9resd/0a51HGfGV8gLhGUuCA1fplYCL57GXuNpgX8ZLv+Ugeup06ELlpowuX4J
YbPnDmwvRvDq8dXbykdNCBT4iOzooPajatYCRNqnlm5YUOp541oiQgxWPGSzgtgV
r2zI4TUdRbE7d6CFFCwKEV4j2XfbKXPL3Y5is5TK6hr1o3zh4t1AXN5bXLrBFKlP
QSvrjXXIpnNfQbr//Mrjyi8D0kITiHWg1A16fh8yFLAHrqWgDrYDIHzwRvbSY4ow
3BHJygutnjF7lL3UxiohIM9/XTWMz4cFZQTOljzS9DhH/96ELecfcDxWQTr6o+4j
UVNcimQyDeSHRAS5Jo/j5yoNnAzbbxnEvabsgjXyATFh8FIEqHItaw4ol2Cnfw/z
epGQ5PqanXoERwY7mOHGlcGvWZXr01Ml9lMqCEG3i5c24MDUReJKQAH1jfLaqG+Z
3w1B+QQZ8zbSJ9hBKEyJU28XpAecRBCXIT0wRKKU+0sxX9MRwk/kTjAw19//S670
dI3/N95K7+y4jFsvZPJG65W0hh7JhwuMeGO1IQWIZ7HjAYj7cZlFZRQweD724d/+
+t+DxI9EzJxe6u3gpYSomJGnx7IKvROjDcBb1r79MOtYz7S3PPE/DRnVZkU030ft
z9Xc5+gr9DtesSmfa2H+zE+9bvSFJ72O7qjrk95yxhiwzxze6vfGJUoWOx9Yg9er
ZWmxFEIpfSmd9mWjyT8QR0iArbtM0xzbCZHH14C4DEySIPUZwItz6+xsOMZM3d3T
X4gRPy3CGzBmTEd2JiXj5o4Ze6owLZG+FSrXsOnmaot0EWXEfjv98sUkkqCD+Umv
evlMcbOohmIGjLoG1x2J9NNtqes/n1/3XIOyeCXLXPCuBYy3xFgElCrtvt4Xjf/y
oPdnpgZoHcD7oHf/8kjb3lqAidAuSbvyIFc6g3S7nGAk4GSd0LrGMeiA8KQlxo2W
ZkcLfRQwRWZNYni1qrskwcJjdmUgR0zwwa8Q8PKCq/8Nls+WmOTcKN3x1a5hwGDt
E9nlAeomVSKvBnmve5rEFpD8wJi7szXosrsrjHy2gAhPRnpayN18c8LeKYJgyCZU
iVChBynZ6d8UrlKuvTsvGodK6tBEF0k1DagWzor+fMne9AcPyEDFBNE1f1nkaBd+
cu97rMIKsUVOl+oXKXRX6AZXwUBJJ46PPzVTMrc1fSn+Ds1HH3M+2BgpEJcj2L54
6iKLbnuU2fRECRvfIwLam+noYQvFH57sSEGcsiM2vI+wTfHQCW2feIIjovvwUAYN
95C18ZcpXmIXsj2X5QmQXdhGgOjNSYhdR46qxUW7Hd9Vmz1/nB6WdChTLG0FJ5eY
1z+FVb9qNBXhWoU/r5VHT7QSyoZdXQA+32XIBnbUbvEiK1gkOgbgg/+kaRFnkkR4
CdcD78d/gAungv8lzqEvj90bK+3Bkzk0KQEypF9nGIApGGP2xUlIRt39MgOLWlwb
iJKuWu5v33PAE52TMNXdpyFoTA9eeS6yCeHXVi+roeTpomSFyGb64HZ9nRFuCq1S
i0qlVfrGqQGv+ZPGBGSdTDrOf4zyW7UTn0qwD0z8S/Yca+n2TGTfUXTu5tzucyXs
1mi8N7rURNigScl4WK+FA0809OjwX/UIAsvghBo3LH8Wf3uTOD2ztjN5TmEx8npC
NfOBjD92sXoLF2lRIqDZtLD1xrt6gE9vJNPq/qHMpVasD2nhJ7Rzk49M41Dhjvvm
Abs6kD8YdEP8QgoCop5TUaMjfvhkGr5mIGKZ4b5AfIA6IlYKlmBrVJ6nR3SeF/ko
nFZEcS1Jdox1zVphEYx2Hjn5ETXp69cM4ktuM7/Mf3JyZRSwy7XyyezwwqsX5tEx
j+N4JWfD97e8YAguQ4jbKiLPxKPJSc5l+QxkhuKtVo7lKdA/xBsyfT8T5kbHUor9
iJq2XEeYYwwqcqO1hD1i9mnZqftw8OzFgp5+z0ZRjQOXKTREfsh23QxQOi5BHlvS
8lb/u3FMdL5nNP76rxlLrbvQBmBz6wYd7sdkGiS3KYu5Ns9KjSmZDhtDA0fLRzw6
dfg8DJ2nf+bDRMYENBgNFkD6TX8/dHsMPr3+E6JRg96zYzF/rIBJZ/X5qemvazQw
37BYX+nZjU9AId7ivJ5x4Wb3sk7l19te93sDDWuZynyh178CIIt8Nda5r2x4RKPe
0iWziZzhOJmLCxpB3hQbzq/9C9mSIqyknTq83inAfOgXxvtoRQpbCpaco5PkDYlD
+zxCVI+xYjrHi1KebcFIngiLu24qXI9H1wAQGe6StOeSMIqT8ti+pdxVSyjVV7K8
BEP0HFJxkYwvvHKdIMCijKsygWYQDeKn3a9x37ojLKgCz31AePHyEXOhEQXnCrK3
lW83bQqcXVjGRWEu3bLZgkmoZh3qkgz+iOGS+Yq8QVxArhSwAsj/y9imX4Wx0M5H
HUB6N7SF4FxQUXx4/SWgN2+19AMHPj7tMW1Zfl08+gOqUDV+q6a+ouEveDOC8vQJ
7n12czgXuT+u67ZaP9rf4NNbKkGZDP2WWPvhaOWFAMF+H0L+mecMEHJV1TDdp3qK
0S1nmCun2BvjOM9GKMmnjnBvj9TfwUt36Z/BOOcjyhA7GAftNodb/5W2VvCi7aA/
3vM2JjLntleZSlj6/kISNsulJLrnLYCm3DV474qPuo+YbJUgJjwQEPSXXwQta+Et
yqDxIx6oIfGPMuAzZwonIvmwmgf/RrFOKlrRJa+G91c5rA9SC78CT1CPtU219F/Z
CJV1n5SCRZFhsUlNvHyCB46xHnkY9TLIfuxMhvvLM2+rtraBuQRtbbwtzA9e5nfq
9YG3vh8li1GeQFpVjEdkNAB21ZE9mm09uHDIcP/uiCdpiSKD7kkE95yrjt7FnA8c
uFX4eBJF8KL5V6RgaTKhqJRABSqx8aYFDq4azYCjangtKf1jIx/ZYbA8lLhp+s33
j7n6id8+tC0VkXJyIWnQbQFtWeSkH1/j+T5Gx4HVGn6nVgQUchc4Tn9MakYROaHp
fnjsVq9wunSzK8I54NpCZWdrbdPLmvSTC/wxCm7ec/WZ/2iEamIkp9M5Vu/RjgZf
MwHWUsZzJskM1z9qq4e2XCkWn7ab2UOhdwC+KLhygdps+h5opNThAsMjAbPY7+a4
q5MtZMqPY1xhFX5wapYWPJjQwFs0V8Wg25wi+QlFk3tel5DSd6HIHausGYZbpgtA
ecKmTFZFsi+chyAS8decr//Cng+QTK8g9urZHTtb/jPuJzr2dRKGpmLjdrPgrCnx
Bt+qVtwpa8yIa+6iL3joBuQX9mbk3w0nB+k5ZWnHkGG34Hz6m4w9ETmEaT8+fOL4
ppqkJM1tTYbKiU14pjERUDJR9A+L+oadJwG9Y7tVcQBI+Ul7pn6TsQx8n6Ut+XyA
YYHpSeWBPrheet1PQYowyPwQ+AzgkyEb+KNKMB0ay70E/QJsPRM5SEVnMGIMV7hv
yaNDIxKE9yJF0Eq+9HW7f+Xgu5zbYX55Zdag8IOFmYvxDsrvEdb5/MIjXL93cEfe
CU3HnDDIgucXxo35jsssf59+He64AG0YqPBhG4j+5PeUq5Hd/0oo1WT4rU+WOAvX
L/X09ItHu/8+7W7lQE0eTX6VrQqKqTZvpHhDnkjaEmo7jYEAE7nnKnwgtHaTW7yS
KBcVEuChRVpd6ck3NLNU3QRRw/oUGE1LunTctY2MY0J1lY3bxnJ3jyNNEaNgjubB
ZpNf3EHENuMJlLyrt63MoCjdlL2ETjPdLzKMy+uEi2/GkX6Ly1j529s9W/RYrp+R
Ehwn+w9d2aNULMm5YwPBKKe94VIONuVhZC3SJquL+N0WMa/UCvVNJNXu0qPVPZGL
0oHPUNY9qS7O665sS6d2MDTfe+XboWAiluRG/no8k3FGAUOKJoolfjwPykLswEkx
QOWf3CRnpc31u6LiO6TlEIO0GDx3WWaH2X2D1i3Q5sMOUzErjVOvAw2PNzU2I8Sw
kp0b3L8/2ssnJwP721VskHttOTRtqv6ZvK9PICvL+ElZtV/QbyHAd4USLMKD9J2U
uxGqPDvEM+yj1wkQwd6NgBA6zLXeyNYmgl47qmZx0zYI/px3nhiBG8/BaB/VAxJj
siL0dKA8yZoJyH6uhuV8m1Ai8wRpRqDUai2Gv4cQGf3ewcZcZLZqcAII4JzUDca5
j83GFMgwOOgOxzinroTNv4ixt6R4Ak1as8qnmHDtx9USygWJOapafkmv3qrdBSZI
av7Yj4oPbY2SWPred6lZ3WdZr3YF3ftB3ebb4r8Lusag5JFNNd5oyxmCm3n3xSGw
WQ9KPYw5GiVx0ehbZP5ICk5umP9clK3q560woUXaUwM/8IGUbxg6XEuCvXGZYv51
h97pNoIsmRHkNJZEsyjbFw2byF43zfFnuZG/iX0P0edlmoLyUbeSVQMYNBJEy9Iz
Rgt1f5CU2CeLV+2vv/cCjz+ud7w6cyakBzoFpP3fmIECVOvL269ns/BtUAZDNyxV
ovu+tX69L2wpRnZsqsrLPCL8GWNacOUWFH6+ec6CqfP1tRhZ5UaKwNt6dfgd8FWZ
Nrf4HmDkTNK2+zhAy+5B3mJylISIjtGXAT5OuoMnHhf6EILJ20JdJDWoqWzkLFJf
ptXCoiw1r1MbdiGfO0TG1SVZfl86vu0a3FvKSLmGsmkdzVNBJIatuJcPqEX0XdNl
f56W5V37C1kczSfWWzU9ZHq7Bc9pfG9CNzgwk1ehDJV14/UtfH3xMFHRkbKcuBA3
qIbVyxfa3iPFEh3yKSZplHG+I8g1wD3WbDipYUYwZERkASfFLCOAaS4ey6sIXJrV
5MOqBST9RiCim+LRICEQZP4uF4YE+XslXsKPGjnwbVvqzDAl3Q1eOP/9P9IWlWLe
Abj81ADCGjypteCpUtpgmxvNpOMh6+o3Kzp4tzcyIZ5NyHaibZqxE35mGljIqgMi
K0bc6rfNNoJ+7ZXF3D0Qf48vyg6/1unUv/2aUmE1bFAmOORCsey2O21NnB4guUIc
W6w163PhVQOxp8l9iLqcBu/s9zfs5RvSoGIyL21BEFaBFdqHmso/+VI8tcFiSacI
r7Yu6G2/KSNflXoIzrdU5EOSJKK1aNMwWbyVpv1yCzha5Tsww4WepWM8J+BtLNp4
RZge9/U6bdbK9MWDKHSAr1ptkoGfbyhKx8y+nK5XutxLoe/Jm/Hf1WFBJ29OcGhD
xzmK9smOPnVOvqTTjWMtMRXbObMoPclnoGjCQ98hL2L/Y9O8jaBBjgvvDrDGRHS6
jxO4qatrrO89r69chYboWl6Db59k0JuNCbjuZeQfTVMUD7s/RA6+D47XpZWVnJOg
jbacReKLeZqRmSPybD85OMhpwSIZzHhr5ACP6jwNdvgbxS/JS+9BZ0pzHt/CDdGO
yhIxLylA5hLiTMxeD/qudYHjmm46PQirxjcJhkrN6wJh54yNoXT4tedAXaGBqO5+
Ih0bhJReImsXHK4Gk9ey4aZuzDKgXUtk1Eieb9/U3wy36tGpcd3IOHWUFWqY0bO5
157tCYtz6+r31Pnxl9fpfniiBndJyMf3f0W93PS2fOrT/iq86vuGOmzqISP6GSM1
KFj23bmPrVtYRx046mvb4g2+8sfWeaAw3bgEYhKu4f3v0ZuNuXWwj6MXy6nKpoAK
VShll1v43GAYBNbTyB/IXsEsWq5IdpYxdxgbPfpUPtVVaLkqXnbv4F9AmO7se44w
ZhErHB0IpR6iiwFkrPHdQorwjcD60dWMgKvlb7LBJ4hYWKzcXmgY8fVd+zL4ofYt
UoXjA/CytCKbVBOqTXn5cpwIy2EBqBzt/j4UHRyj/x5gr5az3Ynn/HsWqIZaPCBo
HSxbXd9olKdv8gmsQvtFBoAM+bDg/2pt++8lTTlguCF5atZpVVLD7VyKwCWKfGJv
gTXTNg343xNrI1pokTo9GgX/Gthp8yaJu209grXq1D+h7hxX7BIWC8pfe9BRtbF3
gQ6z7qLiuAadBTXBfbxPGoEZzMu06oEPTMSgxDaKvNEggEGush/8gDV3EXOVb/LH
v3Y4IU83Lc6wqfTcofQxHyL+XglP2nk4jy4s1+cZfmfiiaLSn8lwUtZ9KWSDxoca
ycZrCXNuwIr3qoAY6VX6NLi4VVi2OTE195KFFAvgn/IZXSzZIhZWWY/QiWsFxcmj
dTBdsqaD2Af3K41oWBxwb5LDbSekoKOsQ7Rn+RbGkDKGPwfZgDnRqIVAVFGwGNRE
r1W9CylB9ioTiv0r9nki9zpY3GJWXAO5Da1nAmdQxELXXwivgXjfuU2jp+7NlXq+
Tr3vriGzmxKPWiI4DFP/3chyqV5eqYUOpMiQ7cSYznEZbRknULK2sOZ980zWWK4o
6B0+VlNd4e7VcYqZXapdL47D0B4pYchIZrokH7G8eXU2TTlNVI2JhB3nBHmq1t/3
D7QT8yN20WdJP+w6GmRaetrFcxN2BTGIzooIPQTkLOP5o8RDfKULB+9nmLKnOM1d
HbCudqyDUreGKI0uBkoy+/GAs1n1wrcHasQ91geSRqpcTZWCbqXyP+KIMCJT29+P
vCDKvFrev+2qyhc5nUK6VUznsGMC8MUaDNYCO/vJXnfGLOd/8OruoPFPp+CHwMnQ
7qADt0UcX4d9Gkqxms1bJBhvMd8iVANSIKPNZUUn8KpfeDBgUaUIt7HpgL0+4qp4
nHf/t8MJKsxUZDkWES+9JGEJ6hryezyd1i3AVramdxOUx/tzuR2Y2HOvs5ic6dGd
BdYWqR1qUJ/+3Zy4fy0L1NMBEbBrQIc/nc+HkO5QMT8XT7cQraWlI60awSZP8W/p
zZ5ZLmXxX8Tm9TGvbroI9nw2C9y9wrAY8WTTXzHc+9BsunVXI2zLPBQM9AnwYLwY
Y67zRbvk0obr5+fZhIHUGK7IvGCdzA568aBWCs/MHiL5Kk9a4GOS0Cmbfd14qs3K
p48OWHuR1HyOWpRHjtK6BekcZTMPmCnfNA5lwTU85/3CS9rjF0kSzICZMcrGzu1M
OXSZluRtN7PbHWgY5efBTkm4peQcQTODMmOfEAeC7IEKvAX9S5G/h8JdNrTM0IIQ
jNa9dC9KBxF9H6MNyL0JIdrEn2oCbrnOtHyOme9+lik57zaBE5/cqJzv/DGTa2ll
R418N/rHhqKprMndbL97z0tJoU20n6oFLtgBUri8ZPWlLU7b02rqEapmWw8AsLXt
dnaY8ZA8ztK5f9B9sAubQa06fjP1Aop2vueullbn0u3U2rMdUV9bH93rYFCz4G7N
nvuiSyfEPeUZQ4yY7Cb8rOtqqNYWiJgSbO8uumpHz9rZNmmjPOoVtlpninsp51co
/hoO3EeBqRk4q/PQvIH+/EQqRg6by3UmVuXnEuBY5Scnm08fTOUVHBuYBiZ4VPON
pcKaia06QhUGunGY8ewBtlo8VLRFIg8t0HnS7eUnPkoGMKEyAyJRd6qV1cdA+wUq
fTZnCpvHf2HK3wkz9seRFTyYB6WqWzwv9B8q/qSjDYgzCxU89NHqJ7eXNgJtITwM
uf5yffKUdGOgQMm/jCAWViZ3hgbILH4m1Z+t0LYfLfhUA7CaKHl3yv7WHXtHhI5J
bE4vXJlIEbuINml/6qzftCZYf79iBh8ZQcRxJD1cjTYz/K7GgPALP/zA7Gl5JHgE
G2lmpNJVwcGnAQ77EU5mwiGtKtGc5ffgdP/+Ew+8tc3h87QkoZPrAHh5rV4DcFXx
1nD8ZS1AptMJBaezIMisoWkKwhOKtO1vj5yz7O5guPxBZpD45S40v6I0tm+SI+dV
Ag3glZnLyFaJqwuoY/BVKeljyzsh9FeWHttLxX4utwyZP31wzkduO9p53iwLIWpX
/ldp333iC0nOIYiCLYJ52xSU9PVtjIvyhV2+lGUIW6RglryI2KjlvJIyETSQO2kp
i1ssiGV4yuppPRcKy1WEWgyVql1O/8JqlM/E3yq3CChI2RtrVzV/ElyQB+jfLW9A
OgIMw81kBHEQuy+WUKSH/WHeJqZrjo9HN45p3DxFaWFDDtguOj1buI+fgl+NqOl+
u2gBRvo1kAztZB/RWxvc6VH+vtoZXVxhB9OY9w6CRKRw72cxcGPFMoG5HYvU8rT1
Gp605TZ/ofRtz2jTZSj2t8u2EEm8hKUpo0zLQ94kV/7T3Agq+BdqVxwLGi1HKMwU
xXDBN4gWxhqTyQCQJZZx5q94KuSsjnQOvVmxcgDaqbl6RMu3qElk9dhk4g7/YZ1/
UU8iJDg5VRy8NyExvzmmcD1N2ygpSK+sHExjRCdGVFPLNTmVFTaemQmaXbaIDbgV
Eac7hfZq1UcuVsV2i5+rNy0rShwn4RC4It2v3zZWvmxGTxwgG73uKWWxsXz9tQTr
OEkZammtjCU0HU7E8Gf+5t/K5/Wa3CHcWdBOYAsjM3oaI9qcY1iARrddbvjvPIxG
fOvqdhZIcHWn58O/rBouBRHWuvYVjyltHvp5nz9TFa/0G+1qLc7OUEvSxBG6weX6
pbKqjOQ7ismA68xn4cub5nOWZbJJ+UnmHxIhnGbh5WMbuKY3nhB5b3rrLfhFo2Pf
44fH4HOlaZnJurMA0JkEP6NdkGc2kcb5D8BUqvxh+t2hjal2+yLlkS6MSXXEf6Ma
/ogdEDOEadXuhHiEZeinDGpOgFQw0mDsrA8zjzOVXMEF/nS/bYRq+kRm/fj+7a+N
g/Ejq8wMpKbsX6u/NNvNMZx9BanE8poS0xA26i+TPcKThlBMdSo6GwfR4xCKCbRI
iGAEDmcPA/7bHsNaoT6Ssu0I0oZD50hGV2OU6NDhelyceWdC5I2G+AKhrhOkW5Rk
FZL+HbQdSYD5ImX/ONZFpamk9mbM+2a2hZdy0Q/lH/Fns03SWT82j4klH/5KZfgn
OfCAwEgj4UWUD8KTRpvZUsd84oDwCtD7dA1AU+VU7o4BXccoeRWtSLVLP7X8OcUa
UfcyirgSX9F9yJ/U6ldsZxD3ZqpzGOlh4uX0V+Udg95nkPsOPrJ1O5niNNJ82XIG
Z9m1UzgGUOQWz6EGNIG1dPzOs73zLxV87mwq0dNenlNqUzaTFG2kaxgels+fgyUa
4ww4Lgqgycr/I3uivTIa5b4DvRYx4THoLEag4ZgFnGqENdZCulz01fpoKVH1p3pv
urb+KKvNyq1jg6YmHKrVnFKQO3N29nBn6qf0y1Z6jaDPVhEYEEmAzk9A+0HIUQfV
eeoa2I4ETNHvogu55b/moECMZXUxMSJXVmJyAGbWB3sfFRHr0O1GLVDa5mcrKErC
nUA1trhBq5mi61r22vFtJlH3UaXWjWgtnRC5GdDj95j2TLUd4TeDCxyoeFcBopSs
u2+6YNFv4sn1RqzWnSBVGh3tO+cXze84IzEARE7Iy5t7XgOyWrCV6zffhHLaz+Pl
frhbsAL6GcRJBLcRM1CS+wpACd5XWqmdjoHpE/zfEdK/j7002NLcRaANfp0w3SCF
mcsGHo8ezWNQoyPM24R4mYdVm6EYAK7A94MjCPesZkBqzId/mmQLJzIXqKyIgqYY
jTJcjI/mHIvNPyYhctyjUg90yoFmVxWHTZl/r9Q7a2Ol/ou3qLMWsoKEhVu35Num
oBgqtpAicpmhBx959KV5ccxTbAG5VmE6T16vmNHBXVixXWo+AUR3R/ekc+Ynfzdz
Qw3UsBmVPGLqABNUe6P6+apAuYWjWeFJSYstWYPCBPYegOXrw8Jx0Edub7TlJwur
j9J1NaYNb2NMYoAEUoH4Bok2aj0/dMTdrT9FrABU9E1Hl+LMMtVI05xw8p0cdzwc
kUgGscNysf2hOFc5Ct/weKLmOD4Pc+Nu4MUkOXH/7EMFhprdiQCv32L+ZYsW0nPj
sMxfMXhxp8qBYHZKlAd3c8iKudaOoDpkCGY+WxbuN5CRAIv0MoKX+3OVr3jOQU5q
MUzPV+IjYLxvr+egLRKuJCttrYX1DkNi3PJ46uFSypwGoxdk0bgtpnhdMtk+hUBI
zDRSb7BWb79tDkI16SyD+GKsl3S71NIRev2wJIQaxvvVGIknBp+ACxF7j5D/+uZ1
iLmZiF+qkX5ufVy9GU63N2diOoJYp46nx23DEW9Y87lcD0iwtW2lkT6LEkJK6i4z
GhV21bPKWl6+kfxu12R8MuqB9PozSgXYjt5qNp6PNca8xu60QFtUBi7a34Ym2tAd
pBhJOozczh4rdqW650gaQ4TADk/PeuMajuZk6ou4gJGiQuQS5Ov/rwNJuLJ0kCey
FdDna1UGx659qUmeoEMo9D0CYih1a49e7N44s0j/Abu6IomEyq9zqlCym5i/14K9
/azr5eRZMe+306A7uOP+o21GFivsWJo/z84h/HRNagXP40fGHslNTiZIiSeJ6udO
kiNZbx6G3ib0HIuKY6/dxx9o2i5L5zJ5IM0nGPMZ95xtGHlTu0HNTSr+ZB7dvZrx
e5zTMrRD+Dsqo+V3Ns0lGrkzrZ+RiVDW+CsP9AkE8wSmphR2CVj2wYzzl7yhgt/Z
ks/CM1wzSYuRv5VJ0ARzxKxGQsX8hS6jZv34fL3Al7/0NOtmh4ojaJ2ElHYMG61t
Cs6dEeMF14fEWATX0ZObEj8hovCbmSGIQkA3MSUJqaPO0f0KxQ2iTkYaYpeQOKSn
UGfWqaUeICH39UJo0rbFAI417GK/DEIKdPMEA8Rc34BLXcgaEAAxKyix2uMmlv3W
rxZ+kvKrJiU0s9El5Nw4nlG2t/Fwk0R4zt/Ydr1ANNyPiHLIOf3yW7qD1G7631zT
UxhqLzxKxQPoXaTl9UDq/F3fTdnsd2FXt/5OrCvqgfbWgWrvkdD+QAcN23dwJTxH
geM7QS1hPriEO9l9mkYoCKVvqu/Xk+nvtyA69mfG2dn17ZDnCJCnQX5oTr2lgNpB
/xOkfE079slK29Rj9biVSjSQ5r+ZMf7qTnZRY3+juA2S5OY+sab+gm92DzJ4GA5i
JG3GVYXDAO2wfVFkPV6adC8UusVuJLN7r9wfCpYO9UCPkfaZlCr2MunwDS03eulR
zSjzUliJ2xOKLG6XsdAdEOlMzs2URITQ7qETQnBpBvCpHIqfaaIO64Nds0bBY5u4
jrtax+Mc5zbseRwuZKrlKiYIc4Ql86akeBRyxfCRhcRm7icJ3JUWGN6Rpx3mMLcH
rbXCHXhIHWpQt1qnN2OqUHI1YDFNe4R/OaWmL4vfI7DQcos11thiSonntmd9oVeY
tzaB92ciFcE3yCDNdO1EHCU5RSYgK4yTQ1vF7kuTEP4xIT6MItx6KjKjrANwOkNk
UaIs7Lb1uRyjTZ62dxEdfc5sfhle44RmY6WH5OwRJHCpJY7MoH+qrdSQeOS0RY/j
lRKzLSOtzpE64HjXhSpStK+Vtvmo5j3YgJE/oKJRejdPipWkfYWLbAU6boKzDXmU
hEALdem335BbVjaSErHt7bZf1Sg8hWiUX7zyXEQTfw9WPnifuk7hiGzBVLaL1c97
HJ5K6pO+rqlb4Y9Y9fLPrZOqzLtWOZwGreujSCvXEF2VxhMFONBws+kiRwz+nslO
3Ns2Becy7TJ//lqmcCpsy2EKsrIa4f4xElWswUfz3EuMBuItKURnUsUV7LcDWhQ9
LkpplvHwaP/ItoUukQERICkiYZQtzExK6MBKqi7r55oPlniicmQjlGKWilUpr0ca
6DIoCvVEyN+Gt6vnvCUF0zNUJhZB+DXvXA6GB6WBE23i6WzolnhS5lXLeGHMyqhf
UKIFQfbUWg2IgmBnAFW3gkvZVbPkEuED4cNLqQ6My4sES84QFBAexnv3ABVn4aVt
usur+hzHcvotI9Ead1seiq7Ot8ss9QEJRklekgT0lMdsz3SgmSlgDI8bpEjLUGu3
frp1SiCCUR3X4Qd61k8GyzECGZ5ZIXs+Wx4fripbqSx2dTZqEsFRchgrFgIahZcd
Pn9NO3txNobBHqVISpq8hwLY4WMjhPKpSoMTud21eutMTRwvSl/0lJty7QfjGQ13
qeKQG0nG6eKpUS3Ppg5C/f1jpLW1MYD/SA3DPzrhpBRYREKDQnnB2TtUsXrx7ePc
ZEKwc656WeSWevNdnVIxNqzW4rvMCNUQQEoPo7s2Yx8x0ac459r1RbDUiCfXY8JR
nnQrVxdlsgeYkdbMr25DWuR6IeEdpmr7VDJIx5f+uy1DzihXjW01r9yKC5PA3LWs
ermD3i8lZJXFILG0vaCmpH4IpSvtcOpj4eO/8jBt9aaybBcVSbIUQr5vzKsx3OHV
cbyLnTE+1rtAoIMU8HyVs4cnV7C7SlxJ8A00QcOOjEfbKoBoathT2fFFkLwhNsSk
RuVnUV7xqgabqNNm0qAOVXsZBkLHL5uvXJTvuoxWCtAGf2+69fNUDM28iX5DBDyw
4VmF23HMHQpHrJ1P/4zJw8yMkliqSx8oZo8b/ZU+zqpcFZrIQHI/+q833oMQl5lo
NHHa2z+g1gCYA6a2hmdwF9eCaLax9zE26Xyep0EnjgyZcB8CZKZUSsD0XOMxQ6p7
sPF8oYbfRddmclB+aq9oomx2MdoHh3THa18rkcFkbgHegRtFF9jjSIgTPQPiiKkX
7rEWQh1GRx4HfjHWJOXBR4phv7GbOsWs1IFAavLNz8pBw8O/FYMRaJSdfNx2dcKr
5QPQM2f0wodpBRTK2QFLslWO3YpHke6VfCsoxWa/iNgjyulSnqGVE4Y0se+kAcMk
ZFdxxASKiOXtO46pCX7olB85/XOe+AkyYf731BFzVzlUXt8lA/tWqM/kAldmGa9t
LKsijjmlnq3z9wQpwYDJimUCM9rjUVHDwRWBC9c61Exo29Rpo7iUdBqd9+i+byFd
usJoYuOkqaCPCUFHXSvZlebZN043XQDgp2R6wrmQI/Xjr5tzSzOaMoW8OumtZSKw
qA+pg21D6DkNi21K8/2u7QmhBsRYAGhklzuUlCKMf6jtKR5DQWU23v2gDNOpoWMl
p34H0pnqPcDdKtSXRjT3c7/akON4htZneWtIAyJhUxq15pI6eeWpKJXLVjBJ2Fdg
WCs97L9qJvQsthSDtgsnhUOkNyASOUXIW9shERNJmCHjB2E2tUMd46MuTHZhY+o7
uyizAeSMMNin8vw/2y/aEoN3f2ewKHbQV2IvELO3KH/p6OENUZibiuE5eW7dNagA
+2nYPyDKVgnoKiTT3G6NGGqi3FMRAXJJvT77Y6WVihaP81IpcoJ6N0Gv33dliu1u
6KVLvYqbyz/4nqElaDHASfPxip9O0jAlEVr3G+ktfgYHgdKy3HNcibzVR9eLjEPR
USJuk/E+hecdU5mH0nC6Iz/86EFOnKd2JFl+6TZDTr5xPpvmVwnYKK6EyeXSMIPV
7XrEMTjH+8Vh+EYUVkxIbfwVfXtMMEl3+SD7YTm+JCOFXEQvqlbTIp/QJeykRt2w
wSFoktVAfh0Chei4SD25QqOKd+GrAr/xh+oOL9tJX4oWRTHj+ovIHwpAQZMctsoz
cDGZs72xZPz/AAZqryGdHXPSVgdAqIbMCRZV6Y5HBxVw4+RNtOQ+AiRKACWDsgKq
6ym0sO22fJLw/14PSa2r9Jx4NNR5jBgkAYtQTZVULk2nvltzwT5Iy3+SfkPxsNhs
dHWfuYRzBSTxQqhVfw4IkrZidAjBCJQn7x2CJdUZsPGenyoyT2TvUkEFUWZHc4Xm
HndZwdRwjgAOZ/q5WONZDP8DB+SK3OcQlssJvpsn3LEZal7f31aPo5FmfbVrnyRW
TMcrajo9jUyBk6WKYOCNAWCbD7/syxBztM3HpHcVV6DQq0DUZKzZqq0l9LiW9iHP
GuM3ANSs0ysdKIs+aIJG6yq9ys2lEov8I13t5Azqh6UUqRhm46ux9jtOqpTxxjK7
u40zVfgHgPhRYxVSzEmzoriwSPNNl/0tdcWXuGT3bFCnfPu+SV208v9xA/db6wy3
N9YNoTa7mQmCcj8UfXkUyxk+Xr3nTOEllNr9XsNtrH8VStwepOIylVrOsSwUff2J
x2C3p7iELZ4bcAEGAjY8qpL2QlfkD0wIQGqpY225jQMhkM9y2cEwG5WXESab2/r6
nOuF1+nArsYeQRoGBjJUcQ2uP6uJC7rGZpWSxgw/Kkm9JasYbz/EgBZ1CdobvPDq
EksLZM3PLzBITy/v4rZ1P8/FYqhLSdfC2VvSO7Py3MkbTo9fJn9JF+g5XRI2nlDq
CJanoOPVReZKtzgupCmY2NkVE0wh70YqPZIy945wQmjKBADV+WzZXkcdGtNUIhJC
3dLw1Gh4zXJf3Bnd+k8jWhmxHvXKZRzuC1QAqnZbP23/3ApFJ0qNFGIHqJyKlWha
xnRe8Abkuch6Qm87zK6wdnAVBRzZu45S2AoA4PdGAO+lPYBkCcQtJ2K7JsUHiSQz
ZIeZuODsdLKh3+x/twIqmn7hxZ/bRjMh/WhEezB0SF/uoF1MlXPZccGHucuMEMCr
stRm53lTl3toe28cRAorERvVb8RQ06HvMoOzvPk7QFOcUHV5OoKOt+cZrZ5ci3Gz
GQmehTsrRbG3xVWJt1puu4ZgzH5e21xeNbCG1phJptTNnE5XhdXzBiUf8NjKxd9K
H6ER5mxPtGXRJu0VrPv9gZO4iXClR2hgySvXzsXdeXaS/coDz6ATwq3Ev3PmLy84
q5HBRMcBnSZ3oHI/gYklQrnh0bj2Pt4wiAEgvfBd7xTeOFUG29cfiQ30iemQUH0s
tcbDMvy1a5pn3w+QFXncS5agY9ASnI4BMWRbKmCqseGF4jsh3YsnoRsbPeVprSNc
qJHsPrY8QbF6kTgEiz+OpRtIfwGLambKMwNFM6mgEeeqZXYgaOafiDyruuS4yXmv
S/L8XHNjaw/U1gxndnLOCgoj379ELTB0lUELUlUkgS0+xpOhzr+QTxWQpRfEfeAz
JrKhwoAzTbjkPfYWFmABkUg/+Nf7+t+icBX5Z+M71Hg0RI6BeAM1d6S2tfFSWSnT
uJNZ7WasSoXxs2Cy+e/1v8MWVQOjgWVcFQKM7uRcqTtwSCTayZUhM0g1M7bV5JyB
tOpFpUE02IIiKY7i7UTtwWS1gwpzcZUPcqXKAJSuvwaE0WBHnVzNJxveRImquTcQ
+0hmRpOZWJrEC3p2Vn2fq0x3byjJVakqP8ujGsHvb9q1gH0u7gppg/L6eh0S2qRH
9CmA5yQtrS7iEx2RHYPOU3jF5w6J1k8CxXJq0g3HyCRVfLnEsaMV5RD/xhWQLyK0
PCT4gv2nx1HY+qfHfcOgq7fXxItY94i+rPAhBWCTnMZLyyt7pgZ1zZ2gAmZnkP2C
7CwmZ4MpOI51jf2XTLIb4+6icewSIdRFCd8g7WQS0j0XU9nG3O7ucLvjTOPsVpec
b1P90VdUKrwhFrhmca6TnnLeHVWBvVMZgPc0teGkoXzsHNa/bJSYSxMjroUNGMqm
iO7MjVMPeX/2bR/m/IBYQnSaTkOxkb1C53dm/PSMJnBEtu/osN5brEueGP5ju+ue
9tHAZn+nuTWWshs48vZuGQa/NwKLX0ikZwYItCyakc0LRniD9F0eNfD5tExxvbMp
eiy0d/I5PxI1gzALZ47gjVG9du/cj/gCmOF3bGaIUyeh3Zb/CIOdkbki+nFiNekT
h2kGQq7ucn8ax+TXjJOAiHhMrj6s1A6kUsEjnCqWxPFS1Zk/3TPIjqvN1WhrkBtL
8p+PPKT9gSTrYCeKNVF22tpONIrhq+2Ma0PrnZqBjXIT8BhEToU1HCc0qVAMAJat
AeJ5aRDQ+uVeYdRnYiqO40Q33j+2WwwOrtzw1C/I6T6JwdDstkGyDaEY4hyXWnh4
M/wnEoj/6TVgSu0F39drADGOO9cu8lcdb/p5mA7YnH/37VZWficfYhctUWhOMATD
u4JfqLYen4p/tdi732mUHBos8Gw7zhgB6yQLot04bP5flScdFtnH+v9m+7P1KwAl
F3rc3ApChSm8t0Q7yHyMLdHDIv5B/XoOggKt+6MCcuxt47oG8z2IKJ6PfJ7tBzFO
KyGz60Tl4b/LWT2JJrtkXjWGKDmxBoi7ODzlrpIGHDcxGD3MzN5lvc83HMCSU3pD
nwpNHmzjMMA85o5W7F8q0SimojNBH5lySwgBUJGgOMwf8PyzY+E3/khu3Fo4Sr4Z
KdHqRd11y1RTy6Ll2I9u+2e2hcNy8FBWKT29pyTi+67xVqfeq6iwlQT/I4PzQ0d7
f+sRprW5OkRTePKDDWk1x3g5HGklgwwolcOH7Zdh120UE8Kf4aUUCOqj0UTHrIEl
XSOV87Y7v462Bqh53qCpyedcAywA58u1JLNiAU9qlRazXFEvniktgaSWzvD6/lGQ
wTte293LClIY2nBRqoxxpWXgMBKs5CeUn8HGE02kBNgrvWEn/z0v/5L4c4RDK4S8
KUw6nUOE17lOznQlWK8b8Spv8Y0i7wB6ZIGbIPs/FmMrlPfKCdl5yh0fVLEUrH6d
YdK9bsAl1ulDJlT8YeAJb6KQlcOdheMcMbxZH0hcSsCzFeqH6qT47A4uSXfqcA3O
YJxsMzqWNUOhomojzLQDvWarSOlvcROIqIw7Fbt7WhnFkdXeOKtZDDFk5ru84fIC
9BsbadchIY18fQglWl8l2Auc5kW7O3OSnK8jXvRAJn/Yexq8W0ivXxSSZwwusnBL
enRaw3ribOVMdiZC1D/v6f+R9smzrdHjDTTGGhm1taTkStKiPiJadjbQU8T7vXTi
yFAmBoSor3aBU2tAXnkOdZNDQWDxznc/KIPwu02Vd5KpiHPgoHkCY9Tq1hoBd/yy
FlxIL1iyYou/r7hI8D40le+Mhtf0PI32DW6ly0f9vKMReBnXUOTVW1I39D3UBJgG
kSUSWa+YRLfOJu4K76LwTEr4LbJOH2Ah2bJSsf8s6vCeRDzfplyh7/2F0HPjjOeU
S3t8UXQnT4OK7+kdiVsRt8JYBYrS0ubboC3DvnVZSSnAN0LiLBiP5tSLAxc6L5Vi
AXwDpEKtU4MHcp+KYFB4rp+3Mt9qN4hzH/dyt/bdXlHu85JFWZ3pocZRGuAp/XsL
gz/36ybAFPGvkHIme8eqMN1TWlF9hrw6IauOPzo7eYKI8XWwbf2GVsHzimTkpznI
k438VTZmpuEEsLRBIJlknvlTugFcABB9Ep6rJQeXTPLZDftaretNS0vPurei51+p
d4+ZnqjshklXt3YLI3DdVs/u6amOAtJX5z8eGx6ptDPSoBQagAR5/JSwK7AyvV84
2kINcGY1V3xcxaC0uX5VaZHG0UjRsnmzcQRpo5PdWLRE5Ssv20b4cRcWmbf2V30G
HClsQznUIE8+yS4YcJ+MKwNZCCkWqLGoCnYEQT1nUolwMq+9csFhpNCTMzpYyecj
RjRreWiAqv3ZKek0q6yEeAWlgJ55hPflzD3eUDwqlVKsCXT7yCy1ByVmeLNLwGHV
4KJhT+QHkh1XuD4ML8zDMcN1Y+NHujFm1WmT9E7rDEoyY7C47oVIG4WGq+P9oOL4
ZpZ1bJQpk3BN5YdgMDq9PRcK3vpitgKrlCgqItNKsqdhK00gKXxEd9q1+HFDTJ+m
QcAUmipAgySmOBC/Zs+b3BUCZm4bfgfEp9vXyG7vrCV/pyZb3UTy3JLeM3Ht6euQ
iiL6plREupndOl9qPF1BSHL/dkjqfroODOUYD0I94zyTRDQsJ+xNQCc3haejskIu
ATDZzssC+gXgVkqMD3XAV9JE1+nAItc1LS6JvlRXgmwBe5hLv4TuWySAjMPeZoEo
wODGuxcNBqG6tFVWlR9wZC/yMVD4bb5wgv7CugpulxTHE8tE1gum4H0uVQcvq+IX
xZyq9Sly3AanQtwX+bUAPU4bP4T8k3ghM3e4LJ7RJ6UKJgyY29OaVmIf2ZI9DkIM
1HaZsqsvQtuOlONJMVGopVTUReaOgWZbkSFdNpI0Sd+aAzLtQT0Km+YKwS1yrJPz
cz3CEiFrog5/LJX58gRkY+gAb15ilwnfQ7+tv2Nobefp0h3oQG4y3sdVa0CZsvou
RzkXiOOCp+t16fXBWegByj4MYSF5IzuoktfWuAiL9x0Unu+gug4VohpvfJMvTn63
MqfwjQIEBkahQAuDvldxP3Yf5rHvLvr3UkWq2CjHiErwLfOwiEyNXpCkHjmIf3QC
Vz122sK2zw6LvrkswQPTX24LiI3DcGgt2XAZefhzQ3089c6k6wvXFmqGMVqtIt1x
3kSR0I67edn8ib+rDKSB+luG1dQ3jfaGHh7SZlB7LS1DBFRks9YzYhbZKFZ3buG/
Q9u6wqnX09BoH74T+Ig0SQjWMX0pTjrEQqWfljN2pD/7FqlPOY5kUtw/vnhYf1bp
8Md+Pbvbjq3ZQrkwVQdOZj/VK13VXYwgune1p/awe5qcm08rbVJAfBPkeR/1mF8l
swEv0qIIl/NtG5b+tNRpzabaSsE27/+ZdH9aORJXXmtcOiV9pMRoPATwekgTU4Xq
VtgGhixcZV5d8N+pXR7fYvoJmfJEpMhS+tb10uMJQD1zx5uDtwVqKXDu16o4NLsH
DPW5d3inTcTQZFxS7LG21X7HULj53jfqcctW1k0gYX18KzIm8V0h9qsVcYovnuyE
AgdO75IwtmiUgb690FOLPkkmpEcD7FghttTOo1O1GbqU7N26jQBm3pgvRH0yGzsG
megxSrIp/XgjiXHW8Xh9EproYESqSgkc6XG9KN8Y0zrVD12gX6lYKQI2yYizaFVy
/Ogc+tZsGO5coCauIJUtP1g3DPSxDxPR0nPVFUYzPdvp2yvwBlyh38EoQPrxglPm
z4NRKeeOv3M6O5fq+NtX5zf9FLqAyMHUyGUBwwjVT3uSo276MBWCgmzCD1/FDupg
1n2NbLJ1VQE3eh0VSJIuxNpAz1GKK7npg6bYe8TOi8K6WwwyAzek/e9Gdf/NnF5G
DgJwtBf2gMWFc4z6U3Ib0D7+2SkAB9PsMClPDvbXzTD2D/Kn78xU+lFDDf46Ywif
g+Wcrk9gGzYK5h+xwSXX1w/OmN3Ep2uqLV8A6JH1pFMMgA/bdb84bEv9dEImCfYJ
sGPYJUxjGNab2m98m6tJRR/BjvZKI55bkCrVpdvNr0a8HBz6t4mHesnEXzUQInVL
2WroBteOsWWpaaf5QDOPez/rWlKnZ6Acth1eD6o7gOFxwPYR+yuGt5ohOJXayT71
Dr98V+PvnMjdArr0Z3xUBIwawnY0rPBVpYhDkt83NTCKlpYwONVw8onny5/T+C27
jSBYYnwirnQCRhAyklTFYj0M+wCzbA4EWFZpM7nPrSQCvSpIaZE3GWpGyEj5gWBU
/MoY083DntGN+9yS1adlY39QpA4BRUgb7JYkL4zMGEMdHKJi6NehozM/2cWJOBoQ
1kjzZFGAfnZkhRG2pOR+REDi7lJlWto5I6eCgooV4vR5YJTGlnR7Xz1isNeTLXbQ
2jbPbnBqhEdG21rcjTcvWD9G7/86xL7C/7k09IOw/pOJFHwDVH+7jkq61sWkszPF
ufnVS30xwSKRoPD2gPyt2M1oNdVO9JZwFxGHCnuqp3QYgewEAyTBxh3KLi0JT1Cz
RGFDUEoL/B4r2e4PQepyVSUAeZIigz9HSJqF+S4Qpaa0vy1qv+n2jsxXNK1ry4mR
B9CyQfzS0uVm7FE572Tjrg1MX2g/Mtk0hdTi4re7kieL2CW9Alwlp5q7MJ57DTdu
nZHlvdYFdvgXJD3M17TwuHV8BucMaxC8MN4vdPrCzoXxJlEQF2iIgIfzxpTJHrED
lal04Da1M9as/JhJhMNpq0btPx8p2q5TF/EuMiR46GT9DnNZ67WZzItjQyubzB9B
8zWha7U2QtzyTjl9fIC3YNYJLDmqddn++z30TJekXnFnk4/T9S5FZfuRNmfSUEYJ
66/6AWgaAlBlWTvZyGK4J4tTOWQPYGnDzemu77rleleBg5eHn+l5X+rs2mE5IsYE
H3aWdpkOZ4f9FVIJ/AUEg6Oq2JGc2LjKCH08eNkay/RGFQeXDoF+92lOL/HxyqIq
l/Onv52DHOTGkU6Y35ZRfq15o04AhFGYp+xiWrmobW8E1HhzfsnoCEmigKI0YqrZ
8t5U8XTibiJytAcYGfnSvOUfV0Ekf9RhY6VW90xtg9A2rLdzcZ/z3P4tNH0Ku7+g
H0cga8IdHnO05mkKPYxNLEpL/wOTT1yGU/x3p31dcjdrs7V7qOZTYRD/ayXGaQjO
3hUSMooMaCExWh30zsXcf7icbXKcwvc6aBwiIRx1U5uP75RaicTBWPa/eM4df/Yx
6q+RA3HWd5E5Xqgafrt8ygkUlVseX1MJV9/limhFZSiX80SAk7VHq7+WeF/x1+Hz
bLqW8urc4t5Bk4s1S5xTZWV8MbLsqzhdjfhduucsuMujSitl9C9HbrEC4muziXkM
c6ausQmedLb8KlTfs9RHivkEQCNAcwqbu5ZHweHt01BUvLG8tXtriW2K8J7S2Dmr
PRq3CMQus1fERw7qTSwiOjFF3njXd2H+xs46X9EBQ+tafeHdYSBkQ06hv/+F4MzI
uuYHlYiIWjndljBBEnbwQYKdudRLsXhE48qlIaFduG0YW7nX3dY0erXlP9POSGkQ
jDfKvs48L/fdboTlaHthgppijGwYg7yOVb8xJVlSBJMkO2mn7/wwDyv7Wi/guMH3
cv8/pi5XfH49oKcDqxVdIT5WrZ6wTq0FM9r1SkiEGqy9/v79jjLIgoVwiW5dlQrV
MAZvbUXYWGZponntlduh4TBk3l3ofX36nLGxF9O+lX0RB9MBHRCg/BfntwaNjohK
n15IoH4fIS6u6PSkKFP21R8lq8/hZWrhPeiVbsxuX1l8U0TnVHRLUxRKKFIIbTko
jrAWqNDyfbq/EoxQUuQGV8nLPIDTs0C57HTNrzgRRJ8Zzbl4nz/KGiZVU/VbJ8qC
R24Q0lylBPsxhS2B2ko6YUqdkMqtZFYVajP1eJp5X4vnh16sGUY9IpfSg5u47fmx
Gby0wqslO/mQlLOvi7tWgBx9C+I0CoeX7jrlmDQWewoCDXYnHWGDXf3AW0YV8mFR
Yp2/7F9ybVGcXxPwoIQIEGc0yuXpTw2NkDozi5H5Zi2qCrpVKb7DZF6sfnP9hEyp
zWxbV0uYpBIqT31zwk5tSsDt4cLaYD9qYiRnyzVKpdrgZ+BLoRpeJ/oC+MRwRhj4
Uvw0aRh+qNd1g3gVqxuKahsT5PP44GLiCTcxtV9e+FUI3Y4YqzwBDx+WE9gCRrqT
qC4N0BMFZ0KHwZHvjr2Acvb6qfHlwA1543XNhL8ikz7wX46aLOtcLf08vh75mMKu
8bqu3CLig9otuqDzVpOVFR46qCs6yn+GyxFuA45dPhYLDd47839csA0yLxBB/df4
6uzYjEMM9MX0o0pn30a6rifYPMwl8Vo0eeMh4BVK9PmMP3jyANeTgOap/kVOE+tl
JFNrIQ6mU37+kEJmZB6Ertb2K7DpZ5DqUJh6zN0Brs9K91LfZFkU6EyEEuVXPi9n
04MjxoVCOuBIr5A5yeOig4Hbxns/vIiGo3H4f24Ry9UFVo4CujfTqsqVaoeWOdbO
W897KslROjqf92Pt5pd7IxTg9LFkXNmGVc9vVt531PIk7n6XT+xdUGx02Hb0LHCh
uKLg02Okv0dD3vhZY3KeOe5B62jPOFftFe51HG8yACwqPs6k40dCxSPmOiPl3csC
R4dPbJU/07FbieRLQVeDSfq3iFSCm9S/8bl5FJcy3v+Us14hMWJAOm36crV4/XE5
9RmCtIyaIp05UzHPRz3dyLpeukNS+/gkTZ4dbPZwTu5BSS/Nz47CzohAqxmZ+YXt
gY8fhbVypBJEiRRaBzflyC+TJye/VE7phwaAlNxAVRFuekxsli0f7IwBjzfseOLN
O5T8WUgG8bZhhxQa3+GnXcofFLPKEAnaOCHRWy3nXfylNh2wttCBc7YMTe9soIFR
HswZQs2cM8hY4GcMTRJwUqpXMcTXBJLYOGGHQUbTmQ8lF2TC5gB0o+2QLrDOwNbn
M7309Bta06V3EsvVuAYqCAnDKSlaxICQoIHclnDqSbE66fU/2SU0TnwYc8UbDqcP
y6gvITwxB+DDJacbt38tnrh9hpt8mrBQwAighj6w+xsSe17ezfiYF1fa7GBsSIHe
YD6yQxMI+3Q1YkSc4t8zQVAiX/iJiXqSBDKhurlCN0ssZBiW/o4eGS4jYB6X57MW
n4S9SLAWPpu8hRevjF2UBja10H4yfx07ICY7C24yhST+kgYaza3afvnJfHYDK1NF
8lgZ+bIvYdG0agMo6VuK2w02lAiO8fFfi4mzKrZEVOXsP0TmkbcJbhXfs6tBjkAb
N6eXCGOW7A+SRdoquMCrRi6AIn6ACR1q7yB+RAfSh0dz2g+CAGCqDLZleOpG8+Pl
h385vUNGBCeRHo2i2+jxAosDUH6j4j5rs3VXoLbPM+0igbOiOg3vVfYnBhCYWxq4
gSIhDoHYUXmIX28QhFrhcXMAop30d70S43LIeN7reiuVcMB33eCG4HV/7QVbzBLT
sWxam5JX8+7Sor/dTuJV06g+k8Lkos+GonobQj1OEHwGuCPZ4VVfjo1lFScRtYvI
f5TtdCn9kbZF+xFrAK7IUQeKEVU3o09SLTEGgC90k3yPMfj0duL5Lt21yyEa5lan
EFNsbaV57oypshe8rwkiOmh5BUyND+Bmlla3C9mz2pxap4ajop/g1V8AuIeeoqEX
Iwf1X6keSA0PWWQekq1clOCNE7l+vHUfKe8gW0QPdcCPm+ilLsv3iYtPZyRWIQmC
MajmkS3aXmGRccis3THSPmAMKamKHK+Fltcds93mA23+0lJi9t67TDVDPPjfwenc
OUSOLuEnDGcsZYaD0zRqNhqtxsKF4/7/+0QofrHOVOudqMN7CqKDjg8EJJGwzXDX
o+0VABuq4jk+4EZXCu0Rg1wE2fG2HXY2tywp0F8z8SwDh6WcbYpU6s/eKrx35kdC
okxjdeAnDu6Svas6l3YniCmBlr4Zh03R6TFxMXifgF5zLNIslwjgx4Dd9WXZE8xO
gRclRUY6tjSsE/mUPQWVk21CBX+b8LI3/+bB0GTr3mzP2FdRuJRtTVVPrmq5O4YR
NAzE8ed7RmKp4kJb5+f+W9D7XOqAsLqq59Jyqum4hnvWhe3cLrrTG022PRb4NOP/
snnYAyD8v96oMrdtsvnl4k/+Hkymf+R6UHmViZOD1VobJmiDfyxadlcopXWNcu22
gAG2U4p6MiHG81rjSnapKqOlAAcnxYYRqKr+6tf1sOUuBJLL3qSMM03Evk+q0BB8
WeaRxJtwROhSgnJFjJ8IHtu2Ce2x1yRtRfED+NBdjsmmgktxKdr66J7N8l6wm+Y8
+YMQvl/CMMTWtckqApM/8xB/PATyWGV7wL6x2cDAmHdRDg0t3fH0vUCyDmiWMM00
/1bc+TUUc4CL37ykK4kHtLDLCOGgeK4BALrrUSRk4QWpmBsTh0Q9gsk618gDrodn
x+QtwXZ8OwGc5rLE3NcM/hOFcpTqxQVZ4btbhrhRlGNxUjlgJj5xsBSxCdPWhafx
YCvytb6Y6AFcWyJULT1b44lap4Ox7GwcPyUsQ2U3Y9Oovi2qla+v7XyMSZJwYNkp
xVvtgFZG0SgqcggvlmBWZu8mubrkVu8o2BnCCr2FWuhBxYHTYwS/EsGu0sKEbSfY
dFChmBx4ZYXBYfaXjnHcw6aV6hqQ5go+6Vy8kZZ2IKfol6b4ltnds9a1olNtu2OX
UKEQ0RAp8fqVw/P1viSRDOtysD6Z7N11YmmDh+GS+YwS2FwcwYCoGRsgO520C00d
qXediZxA7VOcCDkUrGySGV+KMpUAgAMPybHXwfZAo8vAiGSVL9jP/WiQZsCCHz5K
wb3TzhRep2irUSzk5orXip2tg6ohhhu0DEj64xXqhsw6lyzWRGpoZWjH1rG418FF
tNGU1G1CYqvaUT245W29J/lYhvyzlo0deM6EcMpNaGuOCBRhH96rvmJHZqbfn1yf
IdecDqcMRuVyAoaIMbu72/KM1ktUcC2GgD5yFRIszh95318wx5CmsH4tlj8C1hlX
7HqL+5vHLFQ0IOjjgz6TaTjsQqpZUidMEmvMre/pp29ubneiMIiY7YOleI0JDQOt
pXXssw72NL7NQXNflWwwEmmv6ly1wBx0YUXefZhDBJozEVDCvi/WZ8uIBvwWapQH
JrGUcIWgeA6eSjBrJF4zIugGXz320ewXKoX5OsW61Cr5mCxzhOJ2vmaIswRwfWbC
tPXkl+kvgJ8gRUwV3BQ9jRpsSrKyvA5kSNGC/XYasCWkB5yxABCkoQRJK16WUb/X
jN0Ilweit/PmS9k/C8NwlTFTyHdO4sJr+px3COfnaNrf3QvquIX5GhJVRDEJkxyr
WDA6+GRqE42joOnTOVv5RjhKEip5Jb/fQNHqQzxYOeQxWfYpmEQnzK93xbtrZF2Z
Ohn66Z0u0WnnR6DLJ0BTqpfi1Pg3OWzLUUnHML2MUH50LLaL/0qNjFbpU3ew8y3D
JPM3fJdIYEujGQPCP1tIPJDXQGs118unj6JVXPgjLBBQGMQAbO2xamW/ThrzFs1P
YJmDpw+im8k52OZR4OZALjlWK7+yNqbjh/AOdBP242F2SGy/qeeWGiqnqY86Cn7+
PVJNZTIHzih83XWdNMXQ84f5fwpssMIK6Ll1ZaEDiVR/9vhqa0jScI9eJao5va/R
JoogyQcjNeSgogWIT+Nxv6BUcnHe74PbwzBe8MWnc0J5azjZYTjugvm04Vina82y
KZkuHfN5Eb6tb+2fXNX4atMQb9RnSRTlvEHeAEKNDHye5URrKYPbaOk0ytjXLMPC
ZhhEvXesZEpXe4BcsDL/WmIwSLtPghGaLkqX6ShrxDBnqgqUJT4lKkVVTpTdSmZN
s328YhaFFVp2o+pC1d5JENT5JlJPOQKeBDfWWtjVhwa+UwSyNIvt4rexgyBHJE/a
6bOsAY5w0eez73DibBrHobz9MvAbmxMFUlLhhsm6SxWKzyzr+G8xfNx/L3BG9m82
L4VkoQX3qWikv5a5zxc85vCF0jpc5WuqZaZ2Abe5pu04MnCQPEvWdzM+ocUT0Q86
klqHJ2d9ELJCeQE5IwVaePMd4TPgOWEn1EtLx6r3rBOqLsn2IFWVuR3TmIOuZ7EM
jXBu+7vrP0m10BFAWer017RpooZHHs92Lw+lGkDnK4z21/EN3xqiQOg+Lb4VVyOn
UEvs7/ns8c3/2k7wvNMULMJhwD/xrC9VcsbnG6NdOb6OMcJs1tLoALulessnAY31
kUfT3z9qv0kVjo13FC3U5pGBxx5SwdbNYMMppExM7MszVQXThwwSBXF3qhNLWxBD
x1c95FxkGBgsnZ8Amy0jtinTUYhOSasX6JNw1h9TryWf4mCoCEm7QHrje+j15aNF
I18RD8JIS6e4NLe5rv6BPQEhppjV8W/Q7eFvxe4IKC4TUFR32K5q1v95jQlNQKw+
dzl4znhSd6he64y/IP6ORxzPaGJHvHjk8evgJ1WBMGll0VsuOoaUVBf6MMGMxOzl
EkoZ92Ffjoi2ekWtK7q6z2/jWSYr7aW0YH/TJYReDz6OLsmI2lfFiOOYEW4FuEky
3SYAUtX1xB9ZG+0yrvL1QQ2xnL6wrMN7ngVhYsnVbZH+t/5XzLUXhF8x8NdmhQVH
7kO+XiUFvt7E0ma4VyxjzVAQ01yFUSTzadh5pLNVFK/nn1tRPqMNZ+hHfBcD0sMk
eb3PjFepIklikXo1BVPF4RpzZWJL+4hliOy8BT5vAQOxUltmrflt0/3hEq/qpuNl
TnsEleh4RJI5dJV4CXKZBwIK0JUTLWV2UE6L3NhY+10XtPGsuF/XVG6Otfa2I9lx
Ub8RGFNsnE6Jmuz0nXFWgbVdmPnDaAiY0zkpB2M2Ej5BagtsFxgfn0kodpkZlc1e
fouCuCe+QrMntAZNDjpigK0ZhoV+WFvoXqd6YW0PQn6ftGock2tXG77N0POPX4AX
8EGexTSdcLRJS9kxA6NnpNK1OTjXxPBWcJ4kobdax7mWV6ky9+I3znU2pYoV+/3s
2t/kB8c5P05RMt+klrnePH1O+J68Rdwixn8+cdKGzEoVgfFhyp5Y+KQ5TLlUmxZ/
vECMfMc5P4OA+lzyrlvX5uPWkucSR39eKTXEalqOaZLqWw62u7JWCg16w70WscLb
ehw5orNYb4G5ZiMfmCICa3vWViOKRQhUlGJqll7UcHi8PFyrpj7fFeVlPhC2j0Mt
HRDFi0RxZj2QWy4pqLSnGY07yBtycL3z3uObHN23eqF3aT7taKD9Kr5BW2qqa93M
lyQ7uHtu481NjkBb+Li6iqjwUS9ZwfX8GZ6Ym4H3S6N65zIsqzvpWCRyRsbm8JHt
NLuYpftFI1EE6iR+h0o9nk9vkYTT3yMrIuM6UmgbKZf/2XytxGqHmWt/QDKrLu4e
h61Eym1uGaCYobwMwXsngWV6o7oZ6Vfi7oDrKjrQbG7UkVhCegsnIEUYrW460NEs
zleaYYK3DrEGKpdDyLXWEYBrN2jr+avndhLwNCtzMeMsK4dnUI+udBhPFkgnaTgZ
AnIVbzGaP7XPTMtH7Z3XlLnRDRoxtwl5VLwxd3AwQ9t9j4lzibuWSk/Ew+0kscfy
e0Rp87MfnbS5CaWc6BmjGy+QVX6EfgV33iwx9Z5ju3DdW/fbFa7JY8RJk6/giyQF
r+sG8ybZlFzHoZGLnts31mMW3zd7f14PHdLTBqcU6zOPaiMgr0/7oAyKIrKGzWUR
zFqCd59D3oanfNFvcDaMwjVI080fo5jpNjzJdxbpPaCwaghlQJpHjvSUrOr0BimE
SmQJMgDvspfi8uZbNEzWCbCNLU1Sy0DuC391NwG0byyQM6+WIZ8VY00HGxClpRxj
XLKcCbjl2WrQXk4XTKpI4x6U7II+4v/ump3y79xIrALuBSoF/BqhDeBzqD5yMeYi
yEAhwnz576yrkQrO9OqJDysnEBu1LBKzCiY6C8RT1PIlIWLYJw24DMeYLUCpu+p0
acmKHXOE+KpZ4kOvoLTCVPBm0Xfvv68ENCuQY3/UVmadN+YkSp5uJruRbyPjpF2j
95/j7UfHaLFPpMx7p2DDjRV7ksHeobA0PJkqL8yIhOgmB8sW0Mk8HQ8g6a9A5zlu
LwP+jOeseVMbG4da6GodmZVlFiMpS5hoPniteJRaY6DfXiq4/3yHLgM9Vk5zgpEY
1Wx0PeO9vnqgzh75gqWRZSLg0KSkcPsQyeoiGwSP38pLGdslrpA5hWguYK4B55S2
Kp6zhq/4YEigryCBN8tHJzHyDFr277fiym8mVjhPPaFkrWpZrjHWD630IkNBZL6j
mePfXK9DMdltwnewiZ98XAiY2dtLSzeOewQvW9lC5WM9C+Y+ZDgTt8ipj+BarVe1
B2YC6mKdqnHkQckuErbBDM61TFum94d4UQVbIMJVdZmCJ/bKa6rEv/F9mPJK/Uzl
ONuHMAQJOwhb2fPi7uooWiyinneI1esufzf7NObdrhr+JT3ijeM2v0lO01aTn3Dx
AhIFSlgeTe6EhF0ZZ6hux8iDLLBv658t96RQ5dpPY4arHokJGkLkmkVAETbDtJOO
z0RjuaJK+LnnKYrEOGyDFbBUCV06Ldz3vq/gD4/5Aj/2aPotrY3dgLeOiV9oV6Xt
/X40aJySwvaY65Xu1aIXI1/P/N5ifJGDOpyfD20BJr1Cyoyv6MSwko0ZRQ8708Cp
wdy2FTp6ZJVDGIvwdai4bZB7Ze1tGxgTb8E+hDn0xxCBzNbBsNL7ZCNDelZAE0b/
Yp/tCus3ECRU4HvjURIQ24vmsEW5NSklmCRv4GJuL3rWbMo5lAxLlj+5luwjFWJF
Oe928SAI+ydbkUHOH6vixctVAmerPzUoyPBjFBbBdE3znNSsqQ7L+5ia0zT0FLPu
PUqolWxM/OAKTfzrx+n+d9GGGvrmwJKd4e7ySNJDlkC+pSOe/QD/4xfxOBrY8AnS
Q/OXSt5vEXC5RINF75T1LAHQqZxOy2ZVb26YEj7obFZK3z1Y9rpUnIG+E6Mec+vu
N6KBGNbkEPitL/pmsuCGOAfoKLUIsh/d+qvGTjeh/vzvSIZi6htSk7HLwVpuBHcH
iyo7gBKdfYfIBE1HKLJllhI748qYoOWjbWMHnGU1ogPut9RHjpoDjGVEIRGjJhL2
j4K2j95cj+GjHXJhyoGZ0DwdIpXlTI4ahSzvWrK88pEcDFeWSaevl1s/9lwEP1tg
ocb5XmI88bBmcwjt/LO2Cjv5Z5FGsHiNEr1vRViSA5etjKFLKEwoTUzFem+zqAQX
iV1FVfI/7vnfD65kn6Cangv8d6SV6VfVIxL28fzyxhEgRm+2hhFofLqSO+/cOCTU
uBDfgm+cya4XYy4swpN3uuiYNLXsu6bFpjm2VjG0wDHFMqiCVHYKd/zFHDVHEEL6
k1NjRrgqgZR7vOe3k0RaCKd7T+LPHZ90FJzo1wEnHGtnTH9zqD9kIgXpvgyG6F8h
257W2A87aCw+bLdM1GqooG+loqJPTMGNUdHDEegYAtvOcfqhRlrQ2mpzAuaWEkmL
qW2q+FaZ/Dy0AC3FWED8D3X8X7ROG2c2VIWR/bLH/+mz5JIsUEEjUACQ5KT9+Evg
dzb0EfQu1sYS93aOClRI7VWZBScIaD05A4heioaKZw2kC3ynHRFwzixG5L90pSqE
nLm9i6DgLmC2pXE/XxNZrIqJVLSjPq5MmsoiMDAMiFnKFfnYLUFc8XoV6ORx9dBo
ktA71oJfBKpQAJJQB+fd6RXJLPW5Tz45UqcT9rfG4Dw7FQgmRBsN2gvslvH1qJOg
/B8VOJpXF0ynVcRAc3qOFszpIUDWU6Cgp+US2kolYDCh+Gjy9juDRceVW8Nw6MG5
T9I1Z82QoXP7b3EqN295jkn9bfxsGia7OFKyBfb28/JuKwvHzkGmnD8dMNVMjXZH
YJ+w70/0guQG5FAGM+t1JfJqtkOxOYzDlPH1+an48maDJsghT8ADsl5ZLARMc/Sc
BOTwwFPNW9/5chR6kzbnELLFyw3lNmJYXvbF0djEj/yOrHxE9SHTH9bASgBSpGUN
ahFyW1ECPuh3bFS3dWsyYV6wKn0aD0zSUb49IvB+OzwWf46MqCOj8P1a7uhNUrv6
iLag77PEs0yvCqJIQcUCGef8aoClhTBKb65KW/iQ4pbiFv3exhZZqKVosQSQWTJh
m/yLt2zySsZrcL908vi/GcIrLKUaK+NOfdGs7kSoX+pmR/BygtmoJom7Ifhr8D4v
lN+b5IRfmo17BT5zQyhRuM7DvBifdnvSHG4QdzbqnQlLbIVeNevfoRNNeOATq72r
IQq0IV3z7CMq4aBTKDetjq2ymA6MONdgGyBFYlOtjR9EOL5++YQm+Oz17bI/3er9
ZUk6Y4HYGwbF02riCOoSxVJpYclu2XjMehCCfXYB8aG+Kkepkzw0nRrMK4fm580v
p4HOtqoW3548shloZjoxcyB9WnjEcbCfbs4QWxAH7AU3G2zm51RMV0sbMQB5sH/H
vFb8fvRDIGFLZXYAUP0LIYf/kIJXi9YLTLXSpvJuHiNm9WbYXAiLqHruuHAeJ6Am
a8Vp0ymYZf4FQMTk0k0OrcCgSkuAPq+GwOqHeBfNzukWzYJudmivmoSsef8HzCyU
OYTzgVJXs6X8Woct5MToy/S220LmSIrCPZaO2G1z+s9rqCAfpG3Fo8BMjf+RN4Ci
2z1XsBVf9ty2AUEyPbUnujL+ZHpM7N3q93e9tO7IT5mtu31mwm5uzBMNg0dxGmIp
ty3x036Id4BEFuLoslO8J2wG7M1jGnNLYfntlHJkZxSIl+m7SuNjVpZG9RaH+JuZ
6pILkP7+GzL7EnoKMM6syEwEHSxaVBtaIJpxfK8aTmPV4Wm7HRzmqfpn0JeA7T2V
6CRJZZOOlVQBQfdjgEe3NE2Evp9HU6XV5CQ03798ghE8kwlm2X90KfQo+ecg8R+k
Xadc0cqh+Me7XG0ARhQmPnNf5/sjdwmADhOOzQZDdUVW9WSWKJc8D27MhDMJEfPL
BHG5XiCuxKVWbwPUndEA7JFQ6GQrDF6IHLvUaF6bQethK0XB0nlgR742rL+qEDvz
l+wY6Ot16cKmEUbvymnS+dzby76o++NfRlHbIPV+XM+MpwY2X++lcCpfQYO8KPwC
jJ5Px8TUw/WyIkbQp4Vu4NsOalvwXHUVO1C/dkAE04JuOwTn/kGzknoC75yhaA+F
rqbpi0dLtcnqq2Rzg6Hshhz2iQwjUgu8cgsUFEEyAqz9NFI9YR1jWCpdCNei9QjG
mLBz6KT6MOdoQ7n42JNiqlfBrsl8xiH9p21BNLU6zfILCxLigJYpmibZQV9ahWub
3pw7C47m7o+gdedrjc6pc7XrG0hmMyF7pnqRF25i2x+l2DVcVF40gqS7QC2ia/IH
BNQfCKTI1F8dNNfoo2tKDrLeTdOloxURgOPY3mo75ecSLJh2lFqf324aoPhphx1q
W3C9Il2AnZSzCG10hJqPvNmjDZCqRa0Bw1JjL152/RHttDGmc6Aoei2I9AqdOZS/
fAXkzTJ0nMBS5Ry8GXVGz2pL7xo22gvka33E6f3gQ8lG6d6QD5lPeyIRg+L7+CTd
mTaaeCLgKmHX9eOaTrPLxiZmwEAKt2Gf+qr0ZJAFHDKOjfjinORzmhHJQzNY5rB7
xdiT+80Ug0goNpaNP9gHAxHhHH90bWE3y3KO+Rgg31GjGIF9wZ1bQJqaKXwmpJTs
hIqWNYyA3th4sz4VavaA5kxXLWvcUX0QYJdxkC1zUA20YdvKLb1alIQeSJOMp1bx
n9N2m17gg33cEVkGKWCYE3MifJIK4QEVKEjeVWLbaFdZk7c+Ry8tiUvwznWjvHnB
J3FdJtU+bBSMorWkZIuQmoJCErk4sauFp1k6tA6IP6CjMqXAz00dt79i3w5XPyab
xXXnXL61APFalqkixwT9B+9F1BqTSulrVgspareKhLp4MPH5PEnlaajrfXnEV8jd
ts+9z1eTo+71nNsXwxS8HA4VpEuovPy/872fiZ15BRaJrqQCbDcnXZandejZhd4u
CghuP6cPQ0A1qpCqFrguvD5yPx2RIO/odMmzyOsPEsDXGejtVKG6XIOcqVhAQkbi
ZZfoItgsGq6aJIu556gX3VWrxUyanFZAF4Pl01jnbP8bj+/v3z743F/bbiHLqp28
9JpfpcWZD8b/OM9n+eo4JfqdgEDl4FidVPB22gwHsTIzyfFFUPey6rDAF7rAC/f2
Yzh730h2ij0mikLAo+P8yGxZ3b1XN4iUQjuPY/hm6sxRgcH0rxG4QDoNz5onVXOa
uFtA0EGmXSV4X4GDsI2SoVI7nexylCLR8VpAfdASFegg2MsuG/opV9JHMi21L1Oa
Bpj87X+fzg/jh7dmTnOKnfSAlLKQ5gOpExfrUJi5xt3SK2hmRGj6bTCM+2zF55DX
ZHoWdVSB6lYi5CeusjFOQ3us6sSiMrWJZI0ndQWY4p//0OSo/1ivvo+Rl6pMt+XH
cK8aVKLDTYePaJx3uRv7ss0IvNZQ4UWBr5OC10hqlYKeaDP8qrri0VE9YZxmiZao
y7K4nU443yqYPeA0gCzmjraJ5D9CLOZPlwOnVklUQXTLAgCaUSt+5LV5dduXDZGD
Zd38SZITuliDSIVumHCvTlkLDQPIywcrLU8zbxnkWMiQ9H48MM/WfEIVemX0Qgqc
z8GVbXAhfmQV7C5qaTwNz8QL1xRdOc9LOAZnL071hKNr1BhZ4jwEe/VX7lZ/+Sjo
/uRSTVVrUyp2UdIzpsDVo+BLdAZCGqnGEp8gSp8sc/qYHkqiLmrxLpbdl9vjmV2B
uzDRbaFAV79dWAM/kF8yhFuK6QCEmUE6G2gFohettdZtPIk57+yuVhLeV8v9ThxR
fJ6TW1Q32wd4BXFZ35kpBo3FN9uZFHC/uhV93N8cKxTs3qgCIOVIJ30r0Wmf4HmY
26Ct8UPdvRFtTAVa5cxkV3/fCF2HDorvwPFvNAWD6Fm2C2stAfSN0Y0d88RLl4Q7
F5jc67FJ4nBfP7rCJJyudP+LkOm40S+AnNOHGO3pwwdK675IFVasZAYjo75oMTGf
Gi+yf5e3Lwe0TUCGYW68Ve5zG2wyVGFyCC3MZrZTqNy/EYRPkJgsDzPX0pp32nfR
AXQsCrcQjbYd/t6HLRTJBibdEESJZfYdhX3hTZ3Hj0X9QRRo+9chE2eJaK9aMCW/
kCwc8TDwFlSmXVDfPqKv6KVxduEdFUkWl0vFZtTZm0In6MgX62OP+3EcXdjqGkP6
nucyAnIovPu9BNYqaAFKRnLHvy44C8AKEk3fMpIQJC4nd6WFkuAcwAGDYwebzn1F
XyEUmd64hJfm0TxdNxmcGcm0Y+J4N/YWTYIVhPBg8288pJR3zezcfaNZ0YUQy9yk
wOt7GdGJwFqoaresVbmU33IpJa7t8UQ6tnOXtgbvJNSKT6m5rcA45jTVhCH9klY6
MnKHJOY5bn9r6ywltXPXULVdOSqyRqZGdxDIAeqTIwZFtTHj3+6mRKa8XIzjwBO7
WOFtYZ7fQjdCOq5NrQVewrE4p33DBeVaEa86AWQxbjyJ4rAhukBhUN7KyEP8iyYf
ro8tbupmDS27ibZxDxKGOUIfJ6dO4mkW0uhzmw0fsKVaMiqEJ3ZCUPH3OwAuKAim
WJhk+hdA9lt6vO2uJhAELFWRv1qznq0SdJDj1i3LWpUgzGgABMSOsfI1Ac5lXip+
BDoPP58xnynPRad1Vrv8UsaqyLojhc2WQYzmHdiTTysLgdT/yOxQZqvKmkQQrc82
+PHebjjN3dPyZqExbeIc2GZUVPAQdsGxrNwS5Y9ONDVqIEHqQY/yS4aqEEle10J8
OlwXYi2gIbYFvVOgkrhJXwTigHnNFIrKEXfLeBDjKQtWTNmn9sdmkKYQoHW/3Uqj
gMlysC4vzpWJ69AWMeDa6U0z0QVVWusz7/nsTMC5KUFhHEJJKl0ANNvppWMpU7nW
mxF4AF2NyHi72RyJrPIzNHxsJV7MIccmUCZFKqsFX9++KFuV7Z+xX3EkJKoNt0sO
eTOeqXRZeUDc7uJlnGvCElkadLJ4BPyNgObqU2u9f63UBMXPK9zqhiZI4jcbW/nx
G8G0/Xx0VPPNI8QyrqDIHkG/jDVOoO9fbOvP8rIoxrCc/6H01/7aZy2gaxmhZl51
iKDkuo+KAnRgEuu8uPKUQZy06cHO16RoqtYZDgR3QEtAn+JNcam2sjB6aDW2AlWw
q1c7F0x1+L+FE5F/TazowIOAixq1f5xpKd2g2qRrS4D4D34aED+OiS5UqogxJCAj
0Qj6c7klnfEqC62L4aYS4n+unpKiOFjDtxeNj3WC/nwkn56vUNgNYRXGauuSlUmi
iRdbihOpkuyk+hl6X4+KWfFmawtgm4xUs5kBRHWnBhEst5Iy6t2yqob2fmdwCdCv
o3NUHnOWlWkBj+JpyYuwEEDLg4B9F1ql0e4SR37VK1GiBOHJgJZ0zNNW+/Gj9NfN
DMD+bkJa/tfxd4ebQtBM5vxOvh+TlK844ZBjZCG3d9I7n97sKy9bXS19odakPAUe
b0pzmpq/IEudxkfwR5bTHNMnlSBQ27br6UXj4qTGnxq2iPOKEGlmdhUl5F16bhQx
5NTulPshtGNCfbYx0RTPLKpU/PeO2LZW2t3kpZPATcAbDF6Cg+fxfoPNfQz116iG
rAf64q72ZOKlyTqRfhR+YQx011mecw9rOCjAI6XPYRW7SQy1wiUw/TRqA1THY2Sd
iU6y+5VupM5IVerzCK9S0PLV4XL+2Vu+1w+ZJMX5Ws4NZ/Q7kN90vmElU1fiSeBR
Qn3abVLenaDqJQukuPUYgbgsB3A8orQgeMJ5YFWYl1pd0ib9Lyz+B8dhOEOBARjW
kly+4qBPkw2Kar5YBcxME3ahKzIjzGCUESOYltHK25Hanas6FNG1fwstAgd8IJIH
DrDNLmalpnCpVKayk7EidFYvS1hZouyiyAp85HFXQAhbEy1JYQJFpJIqVINo4d/m
/jJ+Fs8XLW7rNwz93wk/X9YuuGL7AcJIKZLW9fAwwUjYx9CypIoGamP9zv9FMkvN
oWgzjtIdeMRnooORU1zHHGZZLp+ZmwZWC/L4DQ/D9s+kOhm04VGxd0d59FmiHeaH
/a+EZDcNj8aXUc1fdjnqv1q3l4ELqTeebV794Yf9yKoLZnNMR24bPzGQoil8SFLI
X3AhddTumZ6OIZDx12TirfuoaqeWMR497CVYjznRWAqZbWYRCqsy3uPKvqWYsO8F
eromyzKP++24Gijg6naZ7DwBx+yeLHdvkeetEcI17bt8eDnASeHsWCH9QNP+fp4O
9Ofwwyo94jRhbs9M0UH5fnvuR0eSETzaNDwyNU23IHoOo3BIB8C+zcLMqCfGD9X5
kyRcaQNmCEVkrjZmD3VfXmE7J0ObItwAg+GFjkx0ykwu6Y7G8BXflR3Iwdat0De6
y9AfrHW4/1jKzdG1HyCB4p0HqnvgS8WCWoqcQ23du18MCAp9iWq6MmIFPUKi/flL
Ah8xdprYg924kyy5nwsDawcLolltpgnq4uSRrT9Vf4npSeakw6EIXQgWlA4u51Qp
h//8CZhplSlenW4ICv/Ak/tlVAl6fldmTyIKh3O00CH0WppGktThauXbcwR1MMiM
8c9Z3iWOJZI5J160IKjLnSSazyNf5VnPckP3mhlcgdOXMgvdjJHebfaFRhK2bdwI
5ohvTQXPdPrDD6pGMiQoxEwQ4j3gIP9at9iEroUs0xPKtfYXaW7FSebW+mKAWknK
VNWQqnctme2NcGHUXjOacsHYLr07P+SImhvLQ/weX+i46QgcHWKsMCOvJOCzUGEd
MhpqyW7DZQBxKrQ70rrAdxyVJH3rkqT62h3Ugod4ml02E3P0M5AKXkDSBvBZN3qJ
qtZyN4maYlSc2N8F0RMiTQv1m33Y1uSCj0jwIyCBc/Onz0Am+XMv/7ExaL5IrrzT
r58lWXSPn59Lx3LbZOfXarDnnNcH4gQGT0n8vh/CIpMA7h8T1/9Zsy2IX/u/oBoD
ziq9c0wrW8PR0iALfzTpVevWgsra+SYbrJ00032qq9lxxmmk9Xkm1bA/215nr05b
kzBI7RiYOkHtW7HP692q9K35r4GiChBvZeFWcnrIxOoj4/8nloX9pxR+BiWO3lKF
vD5c6kpRA4XEQ/Bliv1Lh0JZHRQv+FRP3Gh0u/MyFeKCpqBsGs291ptC8aRsJk3i
z/K1knEy7YBht3UgK3FkP3FNhuACZQnbh92ArTOT9ZkxsSH5MbZnszuSAhRdef16
gMuBsTjHZIxyL/YnJW6GMr3fapewhIHmZtlYL4Uf8wa8k+KNZ6Gk44A4O0BOXjYk
WoySS8DXIh0MtXsmPsAmOSH4vwtkkZdlZMh5FshO26UQckgIb0jS3jz5xXtriyub
jgf4DetcmT3NHkZXXljhtRcsXqnEiy4V5E/dKqgOtQCDsAqwMeFOX4tZzO9e8iGI
PBgJWZyqbfsqn/r0NlTgb8GpYIMUHeJ06KNIyUsLhkUydquMwIHHLBnUZg1GI2n7
cUlCzzaEKNUF6o9S9CBM0Zy9bXFUDLEFxNSrmskDMlt7wf5Yl8AC1RQ5eyZmLm1v
Ytn0c9hQyqITMGm+esI0eytgCOUiwLkWU/o87IeRQSzIt+NqeI3YdWjlw71F3BFj
GbnjfIWPORGoJeplMAgc/YPUlCLVeBYGqeB1uoqSq4P02+cVK+H/izN/Y8bMP15L
qAakyHPX2D7g///CN35+4/Qeg5fMM7+DQo6n+6xItFtd2xAszdjAwFZLSSQoeaPZ
RycKXbRBZDOFxpi5evzy+/YksF4Dxoj4z63R8ho7bB0tKaHnbrRtAs0DHnFVQc5J
9hIprTwpAfy7jJZMOB25CM4vEOJm3RME452UyXnJVmNx80RhSSSfJguMV94ihXaY
mh5G2s4gL9c2E26vq4MJ0vaFfxRI4gegeC2IiozGdgRqv2kY8RZU+WPaqKFMnqV2
xUet8o4q0KX/6WWuO6sgu9ramIAboVLGQEcScJhckZ8f6Aya2m0YxqF5nAgIa9Pd
PajbDZKG35w+g0VDn+oZY8kg17EL7YjnA1qLRyEdfGroKfZ/Bn2Gn5pjC7INjlZj
mN4nFtQOtikeFeZVaWPAAWYgnx7DH308BwtC9ED1WQncwnbNsV/RPzgP1pMiiU2I
n2/8HQn5Q8lWr6aQVzS8YIJp3Kc8xAsA+zKZvcLBtV4gTArl4h035vgFuy9nkGeZ
U+ATNL428P08ToS8nsq338rm4gfjMhGV6LAW/9zq6TaLEsuoDQhUHeTl9/rrbc/f
F17pVJYHSLW1sCMhi+m6mf1PVW4PfnxtOOLK5X9jS0FPQ1Yp20mirxEoE64tuNve
yoddsSu0l7pxMUlY9URy/Q1KoNHxuOpE/2CdfcKlMCxnj3P7SoLuv6y30smFA6fT
wztks0WCMudm0b5GLLLx7SwG33jvm4CyXBwLQp4KhbOTA0hN0bSLO7RnREu58kJt
tPiL99dX34y4qJmTALmuSG+xP4XIm+DYyeRFUlwn0NFszB4FZDv2JegC2dmSdTHt
oUNJSo1KCgMNf3hByKa/g79wZg3JeXBi1PMlVEaVD2bkT1URmpfQ8bR37zpRs0fr
MsaOQvZzAHLwXmiqbAgBYNwUfKK548/pKbGmYrpdcfsG8Ocn9PcjvBVC1ZpH84Re
RLzXNKt67AiYq+mSu6TrU04nD6Ts7CzlrOl8W5ZDE8Lq+ap9gXFnPGm/KI3WZIC0
QjkWjT3X+MCUtWwzbbVk+Yx9+1C2UlpLt5eaaMA+IUzRGahsN7vitgWow58eT0KN
GkcJuK1nHoKNzH2Q4gH3ViJBUyNRfMNIxVcTILV758dmejzFQX3+cU0EkHu1wuhy
5d61Az1tArlDy/yuQINgk6Mc5w/fbElIGcEI13yKV4zUkzHpCbVl6cA+zkz+kAxo
A4kAUV38GD7ypQGT4RLl74V8TTf5QT7fyEox/KbrBU7epYc2vHrZgN5nN7MJYtSK
qrKt+aKMHEPvjnLuKpEV7zuZKvaJsmHqXsr1EMZwjVmY7VOhOaG26sPnpMUMpHR4
kesFhUuoKCKrFp+EZJf1TBZUYjuuPAgIKUCy9d+uD4Pnw4DXyIv0/k/jhaLOB25O
MOihU33c6Tsj2tUHewdvo76GxVnGFRlquKcPB0ASWWKtLGT+IX6FBwAfCtQyatEK
4Nbyolp0NoreBstKaLsv8UGbB9yb47lih2BtLubLOw2FyTN3sKN06ry3wIF3XceH
IVIjnqlUUaIUacIndK54KNDaWjaXFfGEeRGcRGYap2zA5NCmmwRy5qnYdEbYbtVW
D0L+HmUt4qkjIoK5c8rcKo8v98Glr2BEiFdx6+4MF0u85dNe6/uJoSzGUqsZ+oBv
E5tGS6u3M6snvKr0rvbRkd+bpaFPHLJc202bAVF9kqavvWtLuDi0R1b/G1ikvo0K
LEOIhIz6Ax7OOJ36Y1Czr45EuWv7SicLdlTerDKUGMg4M/XUULaS1xrtXBPe/WnB
v0TiYqGMTdrZs5cp/xXvrJ3imc6vYNm2VEFwox/ygYQgSmpzq0Eu2XF228y+0hI6
YjqEYpU57tM5ThfJxQXs0fGa64eXG1FyCiH2L+T95tWnk6Z7Z3638VrABXw7Aeib
Y0i3UeyaySChElgxN8tyBCMmJ0/euaFgLnro+nSZuwkfaMlO2PP4kyJlGDOZEjyE
GQCfKthJafYYBaD5MPPBZyvK2Qp9Cmnk4DXTk4d/tWGOO74Jv0C5CnQ9KLRxAx1L
pSdaUkevRdRnfsbpWChZDapPd767aLA/nLpih076QyGbUVVuqhSYei6lUAz4xGQM
JQv5FSsgRode/VSJUG6KOsD+3pFshWUxTFyez4E5ciLwY+hRxlFftW+UvBNJp6Uu
++aNxPWqKm1I146fynKanxIYFEUDxuViZUdpBIxlowqXW4HpPgGXUdNXzPw/OY5X
ROVRE2d/DplZ5ZE8Ej2hvJwJW9bFmABJkprNV+xHVAXsDXjlP04x3bQlQgiUqNoQ
PVnmOkOpurOVWcrJsDIvRH8Vr50c5tJytP8Sduk7yg8BGprV7DsQ5HfgMk1jmiiF
dY+lZZtT4NvqA6Yi4ItEIS0m9ujtJsZznt8NA7VKQJpYyTK1mT0d//1BmugZG4Pn
F+7zsY2CR5JJkaRxrsrTFcBWVpC1jWbVceC9VLnws3JHry66fmtcjGoeg0ZtTD2Q
aHjMSoHgCEOaMRyO5pFIBECGnqC9RpAfsIT/vaGF5Oy//h+SqCvuK9wJwcdp8QH6
0Ev1J9FDOqtcgzgVPBpy3vUSBIH3IsorJriw1j71vvYdX7O4Qxs9y7PhZtCD2Lo1
RjPr8LZ3gclrJexCRVktVl70CHRp2eKHwcP76PTPLms6Q1w+wb/9djz4Fy/1Ax3T
FD9wXtoLr5vhsAsED2euAXQDJHsLys5gf57dfHxk251Fp/mZvsxM16wa6owKrUXi
zOnROco2+Q4OnzIeEtaJDcA01aVp7REK1gDEmJGDXntM5MH8A6NDMUFyIoq1ZKh4
PJ5vFzig/p+tO+ygLxYhkGDMxJceab8eXlhuftLtKoA1JkLHc8OaejJxbFhhScA7
vWBnnvokxaubyXli2CcixFxWX4VOxZiattlgyo5kSkiGPVXQ7aA9Bp31rka7bshH
20yP3xaRWQP0qJbu73aZ+wzCa/p1BEHCYRXybInRW7tR/nBWSoVMvY/2elxCk6fx
nc9fA7c6bUWBdKwax7f6SYvSYssZ7weWsio5tdhA70Q/ZjB5j/Vz4R+1+YwNDVSW
FRx7lLbcwWqhMe5Cbh2GJBYiGdVsx+ab12S7QScdYtaBKBdTPrV1sEdCby5Hbjm7
sErYnIMu5b3pTDGgozGurbeNsedQXobZZEPRJPAO+Ldh4wWBaBY5D9SsQoDmaqry
WtSLzI/0oc8ohoUo9IvrcuZxFm3Lomai3i6aDW0YyKkWodeLITdyG+EmfuOCGTcW
4/fe0E1CFzn6M9d4IowNHfeRfLU3M+tGBTr4qMmY61vgsQucDLhg9f1O8kh+IIHI
hTXjR0Bs4MR/ZKVH95UyPKI+dYKwH7NNfUiCjUNZbYxLUSVuwNBFFbz2K0pTGV7B
eX8pmtZYV22iVpuLzLvIMrunbliknBJMKc7UVs+zCqeJlgZAPcszHJWJAalsmbgs
MdmkYAcF77n4PTFowM/HLxBnpRTTNszUC7XdPVHB+7l6jZRnExU3TSdw5SvHlolr
AV6o+3gc0KYrkLOyqkexutIn5W5ivusvpQuUzE2jDa8uMnzpfF+HxlEvjnkWwsPg
G/n1zrcsCY9jMyzYnDeaMN2dkkwHWqOHxhFOKwD3Q2U01998wSmEBb83veTtFYgA
xB6JAknzQ7Uu6LxjO8gcPbsBLoOdVlS5BLSV3xLGYZo2NxzMwsN7Xfn4ZRJdEtCe
ccokS1BKO17vfcJbhL3yPs8v9jbHDJuKFBSEqUenIfSApN5yjSHVxhDGYLjy5vrD
VVaTKu8Dboe1PjaNLXAtqlqFe2YfMgwgcHqNxmDV06san2QoMHMCMFYqJWIdRKEq
ndMvwNRT0HSAYqfeaYQdzS8eKLIYo8ketGmO9M4pouct8lUneYJopAwLPqG0Dh9v
a17ApKSjZn+7GhjCG0TzTsNJ5k+qZg9hOaTsNarwCaLoGsfJM/yX5M0xtQwmml31
wf/YRq0NK8PAH4OcwgXCYmQ7pbvBtSWnVh+ga5Z1tUD5chdZrA4P9vTXzCppzgIU
mQQDmR7gWH29XdzpeMDk4V0XFp7JL1DYNS07ASov1+4pYVdbbFj60D1rejaRnff2
dr7A/b0kgm3IWGt3wNaSWkZdpFFrbhtEHz5YtiG8VIUl/vOQoiw/3odPrglB+D+p
VqQqXut1C7lMLrZG92IMzn+AXPkvAK2IbAfJvUNf+I6dP6r71JEENfcawr4K86b+
7KcCIZ1+VbbwpNyCn7Lc2DjvfXnZf0uD5SpC+iJx4EcUj1s/wYMJLX5MuoHxnMRq
OoqbNaUaJmria4LJ7TAN112puDJeHbSV8TJMJU/6XJgDaOUoNFS7fF1HELOYNkAr
9QoVC/HVdpSeou6s0FrxcAOqhRjbrJHVuT9Ys/VlZgK1m3EEJ6mmQbIYWYcmXrp6
EgtYtiiCZl+Lp/JncGoUw+4qgpwcSxCFDsPXvFmIvnuOmjW6UGOTR5LWj7x1AFVk
Nfr9Eu0k9IMjnU3kKMYCsKRpMp2xcP+3671t2jdy0YXW7CJWuxU9tD0Wjeb6KFdM
RWv3t/xT77dydpDGsNsV6lC8GZNoQV43iKzlAIn+sNxkxRELeKZlwlHhmXKyb/0W
pmuOLIXH0195HaHLa4P+QX0qwoeIhzy9Jy7YWhem/84XlcZXOsuWb+xaZef1Xu19
+s1/yfkDS8k+Z0hVkYmIuGQNzBPMrt8LH4xlWZUJQDnrRQiR2eRR+JWxEwt7JYuI
td+GKSwRiFc5gejZQIxp3QnvjATwX+3xy3fijQIeq3h3S81/LcFn3JST220iSdeF
EDRP2nlxkmoPSXmJgfMLwYB82y8XJKrsaLXFrOEbBSttlp6MJs6688vEns/26pqy
UieGCvDdsu7Rr3UCp9kObfAv/k9TBQpB/SFoRAxEqOT7C2bEg3sE8/eBJ7gXOvDM
DQ3q4uSj8KT6lhYrMSH89lPBq3uxDbFwdXr2zpLUXrNPHWx4UEtiwIE9AqSZmxte
b2V4L988cb1HFBQzACKJRscc5ssFIMQHRFAagLl3liBLXFL4Gl+JPj4NZZ+LJd6c
RNX/PXKusuloA3zlvi3tLsxkHGGGrYtzqBRmi8Bue99hA1QGKAKp2uGFzjyXBHai
+JYRzL0kTqLp/udxxRhlr63mp80wyq5OnvDqRKt5T4k/xvMwQbyA/QLMZ/9ChOr1
YG5g8x9NX22Oxvd6NRhxE1HMgDeAgE2w7qzeFZFxbyUkEC1DHhFrcPTFWXSoJXaw
r3M7lWPvAiSaExuHYhoaOHV4Gq6Mhjfj9i8pwmYX9PRq8OczNor4tJIIdBFMKuL8
yjSINMHX3teBz2z7PStOnkLtLOSdp4SdEjSTC1vKRx116I26npQFHZsHHs8NV5FJ
ETwa+KtZELE+RBdERdQwqNudfbWa2zUZvbXAArmjwdK1+ui075W4pWBxvXPsehSO
tMtgr9qjVtIHL9gWbXRcuE1pNFG7l16uKh4ch32pKVSUfalTxjT+yyP6c+FhmjpP
adZxiXAwpCpotPIarfA8hdXZ1mo9aUBcoR0NkAtFLupFtFxaFHTC1bHHyFlglYh+
MI11T7akDJIiON8iVN3JfWR/ggX6fo3SpBXsjBe1AjxpcUqqSgadmJ619GuKEn7k
mxN8HosHGTqyiHmINd6u+ZUctt0p7TXdYSmWPSb8Uxv8ag6mdHuNMZDdQVfoUayZ
FZjOuYZUFkAaMv0NiR/3lUCsvf87atGeycobmfE5IHipYY8r2Bm6m6WQyPD9YivU
Bnnkj9/zsn/JCXC8q9xB/qWq8w+bZ0TXw6r1TiuBmEV9KX92jXxvPCeXS191/ORE
/sPbr+H1Aarm7tA0kBwoWJ+EeYZGA2Zcj5+u1uzNqiuhovKmJG99Vxzj3QIc6Vh8
7AGE9qQJYeMslJNunUXs6uQ2UygG336P9BPxBdT23mv9l61mP639rohxmwdZKV2Y
yzHkTEc6/+XC1WMo8zJVMsK56NLjOkn+3+RpkUd1I49nl+byNZ0gH9ob9n5ofkiV
pFMBa/5shTEYCV8d0GzH0KVZPa5Bwcx9jM6S5mYGiL64U3bedI+0O9o3Lmwb99Cd
EkyN6kJ7UrDw+xp/U8kG0edTz1ggCWax/LyH1geoSYrzXdin/w60OzqoxRLC+XYg
984cf0rOyoV0K5UKzJhvMRNmWINg/plQaBC0yOIBq57GOqMBpNLDHaDKkcKmAqdG
zeW+MviZ3aw+5v4bHyd+yUUyqmtX43rMiskl8YoopLI6B89XJpgAJpaSSkqKImJg
uN8ge/EjHYXvtBRhTfBKwlD7I+kX7mW1PIywkXPmIBv1SCuUpUnG6zZb1u/QA3Lw
Lj9wdaNEoNUof7fwPK4F5AihQ1VmGLz+1rJVHXUL3Jb934tj34K7jcealwZzWI2S
OsQZ02cu6EPDC+gExrmZllifw3gPaxugXyhQdP7gNA1jTMTIItbSd+KgOHVAsW+V
vuA5kukwMQ8rrn8lGTjUEnMJIAujpHbb+L4KsAJhkkvKYiWCESKNHzuHtHuEg3cL
W0JJLRn2KATKwtNBczZy8QeE5IK7WIZPUyS/rp/ilPbULORhq/Ep0uxf/Tr0FK9A
YTkgEfY2k/0mu2GNbRv9ejM5sQiKqJsS0Z84q+gsm677QdV9mk9ZyVvXyBUsgMRR
5h2SuNnZyPpsEaiu6KPVn/XjeJH33+7+C+g9dWLEIusOjO1H8LTqjB1/ze8S0mvL
hMxD+SUPYwNvO9WVhLaCUzVgqnS0b4lpNFUaMaJetNwzaoJdMxQEOCyg8yBzoQ5+
WO7xIFB0xnHEjrbfSqvnNxi64FHGEPwvMlo25LPup6/I7HLah0MxLP/9ysbmMTF4
r+ti2xacm/wssMqQ1ovnKaPvCKDwxPi/RvgGcqHnHPpK6MVj1rsao7gvcL++67Io
6BGOVnqtuQOz7Fp5vV9RQ87PqSPXb/cY/62/Unkakxg1/d2KFojQOgLQkJjPEP3L
hbCNEFyy+mS3Mt4BlNXcBax4X1eH/30kf07BSdZwJTWywTkvR8m1dxQraHQzZ3Ap
kp1IE+tiyu9VgyjHDSDI4Pd1DlUbTdrI5K2Ml5bEr//A3qYYvi0g1KGgyO5X7XV+
65AJkiaASc3sL4WhY2daWxmKGvNUl4x350fHSDh6gPVoj6L0lp9m1n8lCkqyrlJK
s4m8cdLgzJUh4yD2yv4pqDMdUzOt+jEnlCVayn1de2FnNEfXFzwCBHbIebE4A2cF
YiWM9JWrWu6YmN7Lr+HRxfTcAFLilx75dBW/kSrZaJ5btP1PNaOzEuSIfQfDMTJS
eylG/sfByTgQst1Iy+wTxShvE7UVsRo7jZV5FtbcJis0KAtb2c4q/Y0U+wpqecXt
2PVBx/ZgHeyduU2gz00XYwu+jYb2/0IlXvvSWIPAvwZjMpGv/dJY1UlLjr8S76pv
7qUVycd+vz9w5o/t6TbsRVzwbiTZG/t1VfBzapoJIYFvrdP0Z8bx+9nTmTXXhdQt
rw66J8ewcGUrxdRTs1oDdNdw/OWVxfP9yGDnLveFH4oZoCiok/Izyi9bV5cE5Q6/
pqcTBy6rBWxM/cBjmLphG144ya6K/F4v21O+uxFBw+SBoty0BiotAluqs2PVo8Mw
a84oj/DbAMlZwOSm3mNxGrV1plVWHoOjrqlHzJBxVY3HKq5qOqFSuHujVqPG06BY
PuCGoT4SksmFD8WIVO/3fOpy7p03NggUi8XWEkKJDUx/dc8eafHU57GoWb/ZoQq9
6Yawm/eZfpwzWpS54ruGhGN4TPWjXxBB8WOVGmxISSzZUDEz9c3zRP+3NTV1P5RL
oaJaseKLAA3YnPd2ho3OwqVEUj5xtGWsTSwhpuSkQijOAMwqSO5ntM9w/mIiTeL+
e1xfHm42d4mIxvWVrqa9rNRAg1HOiYmLzCWhJFfKKnV+FNBNWCA1EFjAaSdxenu+
063ENCd5l7BNaacER9l4wINTG+jcJz8rZO9ZCa0VCbz7KBHROBYR/sMzKhx8wc54
5KfDuDDaK63eBx8vZdzgdYQAxBklBEg3WDc1F2jrn6TBwMkbszvVVc7tWhGwmRgf
KnEFcjUcQNehWqYSz+WqCIhDDErvr7Dl7eXapqmV0Ow9h8il+q37j+5WL+lbq4/t
K29KoIElintCgHv0outcrk7zmqk02igEjZE0VQFFYRa2o/wGUKqDJzkVD9V+MdPO
2p/7hgXFRNz3+w3olvluiGNK9yxsPHelpLB6PDHMOQvhJKEfzN6Z+ovQCl6eHFWF
NOVo1fI+jW6pjcrjD9JOxZV7Zf+yF7n+LveLQJswhQyBwez7/q02s9TZsc6GbzJk
w6XAfxo5pPYGsnD6cNgLjA/6l4BgFuxMTswNVK4nwtePWW/GJHtBIPEPz+BzlJZP
diSch0hcm0Lo3Ptk0w9pX/cc6oiccpWN65KyfYlJNZxYqLJSfM95tikTClHvbRjl
343AYu7bElNHN5oQURJDaFLvX0yyamkJbeSdw2QL5lat5aUKjzizU9sAUfy0O55n
88XXjqgbeXo8hCuLvKWoyNFZgCVfVsT/yUijXtstte1L2mSIEsVq9/wIvOCggxyd
ordYPPQkdTEBd+RsnPzLD6WZYrocL7ggkF4zuq8rfw4zw9WrOtvaXkXBT5qFZZ7j
cqVvLTcgfLxCXoF1Gp3yS7f4polQvArKa+c7kJtoNegIA4iHYdOL7z5LByNzLonk
ke6AAu8qy3ctHA8BvzZLO3vlwOyvHGURqbP6X1PwRntkxwgAJ4A29Ug6cVyVVteN
kEKw38bvyCUFFniw2T0c+n8sNWOFamrczqDjH9QyGxmEQUQZ7tZXEGa/DSKEIvwo
zv63SR/n6xzvMskBBRQXB2zYjs6Jg0t1ON60eA8BPb74PNrqzTNljS7M1wpMSUEo
2v4IUNTb9NX3jNBGZCkad4lE825J6nSbx4kkH2n5+32LlFPcNu2GwEOrZraRWI4k
oYAXN3ZLDRuyPvPP1U9wtD3TuuM+MTMqcm3i8kC36xd9b/3/iyNf07vi55RRDPv8
RfAIfG7uPOLqY8i3LXKw7gVnZC1XJAux4NSk4pEk/ZuOJsAutsGicHjfoYN1Y5Nf
8JyrfSFNDFJfDk4E0vaqOh/rw1trQiRtdvEZFBuaGutkVBVcYpeRxQtTLLRRh6P3
eUx7IA1ZjbxI8kPAV5kMSqrCRhLRx96CD87hMIUMLLO383A+YDYKiXvbhj7N43Hn
GpHAFSU6dumv5kBIK1NJp3yw+M4hkCSUREDZTikq6vKBvCzq0gs8eaGX3vtX5rBY
hJzEBh1ZNhL5IuQnhy3QSbgwVP0zfmsN+RlunvWf7rpC0Rbm2XWXU3mhu5wvNavH
zWrHCl0LUaMv6a6Kl8AELaPdBUM+l1+2WoY6jNou2di1d6nZ5+cGWnqWAC/4vT6L
BLTFQ5r0w2ZeOocsPKdUmHjJp+ImWD2tlzn2D/vQLuGQQgKHyGZiVSe2/ITw4YNf
3CVd2FAMzmBKTXHidlsx+TGg1cUb/xAdEgNLjbBCmhVWboLKUo1aBcNP8lW+3Lyx
QtQyxWTz6mhOiGxZyaonI/RBhanLRqTfN62Mj+955a1CasDwDqAvSELs/Mq41tSI
7XVttPQqV6DMtjRqEg/rqOohoQeC4DlTCVswBvYJaxgoA/OQeyhA2TSkXciqeXf6
w75Q9S5YSNVujduq3nqO2tBFtp6JvWOB6TQx5yt0ZjUQP/kJ9n9pPeyd0z7M1gdV
Zwzrpqj9OkZhezEsBgqxVgOFHY7kyXaGUQiz+1691O1pkjQqvEl3+nMDws80Z66L
G+lmHYEVMrez6UrvzvzI64kYmLspzV4ccB3zfEIPtqsSBl3NFnVPUSx9A6kxYy7f
L06sM+3uDDCtsFB/zio1BUp4kw5LR0Jp+ERyUXhcAaBZjfbV/Y0i6tJylevWQN/8
Un/U2PjfmpIsO8FIbyR4H9ENwAyoDF54qerjAvzS5YzxEIpO3i8a71SzWEsgANl+
AT2q8RTze8yaMbr1mim+m7BqjJWVlCd9dm5T470HWogOjN31qUpLdyLLHOOZkT/C
8DJrQj5YuWNUvA3nHg2adrsjlHLhHx1gAldz1K982ih9WOBJP9GMQ1EkxENVzYZ+
A9HVN+KCGQb291FUHcWzvoPviKNjFjOAhI2qBObKvHSj9V3sIswQgnPhtLUgyT+J
CWSfxtJEuEKGbx3nUIQOnf12gGEg9lbZsfIgRnYZ6RyqsDbI8AxAppZAYJK/0zZo
wzygIyT1+uHifJIEzjqNohuffPMYKbunSNGpBqt/11av+96uOxoHS7ky5ObDg1JF
/d4cElfLlVdnLPKyLpjPRFHl4dZpl5Z2+s3j5YTNhYR5n3zMyFb2MythUFGvIoZL
dcAALHPH8mYgRHtUKqC7pknOZBmOQKnoLtOsLBZsk3wZXP+1bPzOudPteUM3AzqH
z/QQlMPXqJqXYAw4ZEFgp4RP6DpY9FMhXEH/m6ceztKQwz81IIGzIXy/4rzN6zoP
MK89syNGLbom/mxnkpAkcCU+4IV+H561KaaJWg0CMtFHPvG1boIjpxphi3BV77bx
QBT41VXm/3JlEzxkXYTXsjhR8Oj+tKLSFgfudaAePpkL05t3NsUcHiDJAW17ev+M
gRu5OYCT/7TOQGaT9JiayqfEb2Vrhp1AgMUzXAKvFsjhJC8bw8DyY1H3KcIcE9x/
NmHwTVPiM/Gx47WnEaMhi3gHkKqnykyHOPswONn6GxdlaWeZN15LXpY6/ez/96/1
AxnqAnABwc8jERYuP9b/Zb+pDg3dzDthHISwx++MHwapUP6ly8dStWODTppbSrRo
f2c3ARuATdj5dFIcRUEog69UTe/w+AAWDbCVuArSw7dEc7WoX+NNDjId/DQnJpbK
lToYlGS6bvtsLDu1apADVMz9Vf7uYjJ5jijb05Tn4+b/bsFIkijYWpbkIhFy8fiY
BlOugnWWOtPoMah30oymf9Zcxr4vmxeXwf+jtp2nArTtA5gnbuk3tp3/ML0WKa8j
sbPy3Skf75xQX5Quy83g7chslJ5+7ZV/MGrxnAjRuzsjoFzA97gFolC3ETJw2Wv2
1dXxOS3FTYm47x4XGtznHk4/UNvciFQV0r9nj7IPZYCgaFVMxQq5Lzhaad0B0vdC
L00nITfAIb2TXWRZyTceYoPRtylA5MDVAXdLtgM1AlOcVnkF0iLvln2QuUioT/Me
HMG2OC8AnOJPt0TYMaBt8tYYqdFzgry+2tzSDUVZxMyWp0GdJj30EdFiThEsyUoZ
yxX50pr6ydbEH3VIv7s+raf9CTuLwDnw0p5/OCEJQlGeEaPb91nUUzYJxNkjbEVj
vLx9vaAg3Y95Mi4VjERLVQMbhsue5yKKK0qT1P+rWpPgKe1HWxUtsj6omYvdhmvO
uuPqCVYbNYyaxl3lX1iXeLoJ0FV2ejjM9l2IzmJEzqEZMwfkT8CQvv8UmQ3kEKGx
yv0gjTWAXBk8QQ5mzGuec9A//k5hy5kSxZ9n33VXPEJcoJEyfpMK4q+lzJLAJTrs
A/Jekp+9zwA+q0+1HeQf4pSbWa5TxF/X80Ks9dmoUIchXSomeupmgYm8GM4uN/wW
P6M92t4L9f4Jn2iK5bZuGhewwt0d+5V6Oo0JgK1N44wwLN1eiOCveVxt6XaA9K81
LGuMB5WREBSAmWpiYSxSJ4rLvNU+5CambDq+TgukNNInE6/78bT5Kk3toHZkpYWb
d0aSgXrze1eA609MeCUL29NAzsoROlJpq2o07p8y5lglZPcwONFihOycFVV2W3FC
/KGcOkN09xD6DFU1RnDSaiCH5xypnGTzdXONvjcSNCjg3Q4X32dtWSztRfyO31SY
m3HQ7TpUyGHGLKskCohjBjwg86q1q3ejCI069T0Dyio//RCUVGZY/WJCBu6youiy
SuiKagvAMwBELwC1RUR/CmHuVPlJuGaVm0fMUp3WxuE/C5qqySUGrN3lVcS5AWbx
04cLk941xGn4F7EbVs3GwWIaMYkGQ5Vmgr4n8J6S81cmsC3woM+Mvus9YS37cr11
SS8FyjLC9Rtz/HAMWl4JFzWrUPj/55Q8DglOSphapKCspbBQM9xHfOLcxwoxVOFb
rQ+L5sBNV92rCn+xQiqrY20wtiyfK8987e+zmvkuo92H+UT9eWQULPPZHzW/cwB4
sBSnbZ2NKGzQNggWjN/NAF0dTnv+8L0t49O0xgzTkaQo0ZCHpc+ol2Ds3ZM8OcM8
PuUr3LCqGE/II9HpotjRKnXJSdsOYljdq9OK1pjrOnEIWXOIVUIKXCniD79mDMdg
zzbF9N5JJGdwIKfQsQHQ0DRcTUz36DzyXArZPPJh4ITbeoM2Y5M8vLiIBc/n6f3O
hJKcIOgLDX9HCuaZAnZRmkxV6EDr/In2mg5R5s21PcRNo2RBuBZb60wuf6v4+ZjX
2epdSN+84aA78ZpPLxjZizyEHogi9ci1UoP2KjDEVBA/DmS60LiKAdqSr9NPgkaZ
hFqiBPt347mprvGVEZEeJnqe+rP5XDZQkFHlkvyII2fX9LtEvEMfn+jGYJI9JIok
6uOggpl5gNUP76er+yUxlVPsz/u+sIhweTck9a0cecfMy219rEnKTvWKYtMoIIGj
xAm7dAPoLnxU/Myf1vZFasoy8cmoyU+YtmyzTzxoQd1H/0G17fnDN890AQsZKf88
Q/Oz+kTJZmyvyNrwK2wUhL8z+Wp+eaUFCzptDSzGm6OYnxT6Bxk2fnLj6gunrMGu
YynNje7ZDs+JwgGYXNVH5hz9XK/xarzAMGWALkqwXCbdXDELy4L9Y7CzM5ryAT2R
fBZDnVUATX9Pl49oUtt6vRsC+x1mA6DByPybVXsTx0sb7Gg4Skm84Jv4RjKCXbXl
QbgI0Njp+57uxf7KsUS/eptoA9KmjPAZD7nCtTXwDdoe9uXKTGgxGNha1JMuqkfN
tR1/lvOqTeCLDcxd6dhSCLNJ0E9BDQ8Ls5TpkvFsZdDt6I0fknpxYl0UTE1xf/gB
6NKhQ2NTtclA0+4xHJKKQvT9lbtJevEMbkWz2/2OxjSKOQIdBZwL21sr3tOCcJlS
GlzYyQfhmBO08CtBOZJbUNBXdp2C/NvoVpK1lJ7ThIFhlXTMqFTWUtAOUqDnrxeS
L+YkTf2/PVIxfukq+nb9d7BE97yj0ywt03j0qojlouVS8X3fOcRUWPuHbzT+dpKu
XQkOMN9BUNcbxp2jP6OPkyi2HoIjzf/bGRsUmBqerNAcrgtbqNzOrafXm/vewgM/
sxRzAuh+Jf+z3OWROoHps/pUT34yHpWNnby1t2MySn3hyiO8G3esPSS0D3mUlR42
ReFp34Mem4hbpCGRTWpIT5AQFO9PdZwC5x6rVi81W5WNtj1jdCGyjgBYPVDJArtJ
e/LxokZIu50rot36LHhcwqpAPnUU54/8HSv+RN6KxBpR61vaTokWCUhe2uLCHIIx
84c+f04CoyHvnl15AWdN+S5tUXZz0HiZ6vZAGpiHqHi/K5KzIGIjj7/H79OTog54
R1sZtV8bXeLwjuwOlALV1PP69wowPB+FfMSZT+kffFmlzD8Piev8vwaTgfmGDwm3
pF+IgxIFRfHGM26iBpYGLoZ8qXDkw8i4W76fh7v8X3GGHml+qvpmpqEXVL4MX4GY
uxFVqKN4uxx2o8tAuh3SC6mBSqi2DP+sDAI1smd9IJiaZJzd77u/7XIqh77ljIe7
FW/DbWH53v4xj8TlLO6wgBhdFlzloD5CdUsFGLc9Cxm8sOpxfwFDKQdDcSfn8Vqp
PU5SAn2SG4gTG8/I+heacwtVj6ofRCmFbKDcDHPjTZP6YmwnumxT+egeVZb0C5Ti
0KR4Kc6xNcuGBhdWgAYrhBFPgNtlsbKWgI/Q36zjviL+gOPy2GHdH9FkB0jaXHiU
L+C9qG3S0rHeluykp5834lOgBmcp2Wy04fxkMabsyva8T2q24sWpKZjpdQId0EQz
Aw6bZl3q/SZ8BM0Z+jQ6FYpGcW55zF2mEGe2ZVbOSwdsUvflvTOc5QJ4BsMNsvEr
kon0wWoqdv/XW4/oxY9odSGNq7HErOjQ30xnQ8fg9qMN6hZVaF+PDmW0pGRLQB2c
j00KVc69yfSCMTPC+zw8B0GNIaV3kd9/3PUuB71ELtde1NjDnHoiHhnjRGcA9ubN
n5X7TrZ71qi55JvTanWFmkh/3JV9wRJ7A/UK9m0ZbAFRviXoe9PKBR7v4KpbQj0k
fQG47bJrI9sEsFj+/F+ZlUuwVjEUh1K3VZvZRbb9zkiFCXcgqg8UoDYgZwLljN24
IzEE7trtwR8VRlKt/WriWE8OEQ8J4pCfvbutSkdvjnJCZNo5uETwm3k7czhH1Dbw
SexBRCmmHMiMz97uRqFBnp/RkKDGvKhrpX2ZJTPPdpZFedLXSiBERwI/C6R6S2jK
ymn2bc2lkyLwGH66uiMfZ8yD3S2Ns2YOHnl8y3DpG9NZqmlJMdbnDzFaCjd2RQ6Y
gixtGlUwlvJ+kvCegFnLKR5BGE3g0UzveI1RioX83D8W2GBLj7nQmIO/5IjNmGlS
GhxVFsUrRfOlrEcU26IRK1O4jIJs0f4ByT9GfjyPLbgxOaueGYWuaF1Jkgw5yLA9
RTsKZwiVkcaeMgb6nV+luZCGRv85USLSju7B7NHh/OMngs7KQNLzOzNIWrEYL7N5
efgGu6QbQPxvak71fO4Zk1TpYlb12rHKDvkZfZDB1PLw7Y3qAIDumOT5+KR+9q47
Z8SpfbjHZF3zNPijm4joVkybXKWTDUz+Mpd/8Fgfq9F5Z3102PURamRLwC8s2frw
nAfZGEB24DXjkT5P/OZ8rclPcWVSPoPWmKKrfreO1jerUGJRyaoO51p7Zj4ZH6U9
s6scg5HeNBJuElviizrF3t8isDZ+UAynYGAWdlsSWLi2j+FAS702bvaqIelmpfdZ
A9sbKnKjpyVADsAJfBwdwufud2HmFvJp+IPKUFW6v3k8MpEvOByQKtwG63rGxMZE
2yEx1fa2MVpeNP8oloLow6w9YAIwJeXj+QuvI32lWiZ8Y6KyHteSBf54ZCxyusw/
unAOMGKSQG++n9eMWcsiA8O1KRC8S+2X29UhnKyWO/sZDcQ8Mst5Fmj5TywKfht1
rTb86ZC9XA+w4fswlfao8GcD0tCiCqUB626bh4NRYWIms6lARkwfddNdNoxaXDlu
lm8D5QCibqCbfQEXPPgHm3YEK5lXH9YDKO3PfsnkxpdnUDlWQpCUWubLrIyO02tO
EfLqNBvEqt/NxKkmdKKVA+LBYE8uZA4EoS6AEyrZzCjkK90Q39pHI8PbtM1GGBir
EPp/dzTo8stUu0N+uyJEo2kDKaPgGT3jlzDLH/5ReeABF08lNHR+H+AvARcu4Ijb
LfwGXgC0k3OYQ9nBFwj3ZVi4pk/Fs2CdDkpIb62hdd9U2CrGauX+pVJKDDmSYozy
j3BK4oApyesJafSdnZjYFilljySAPABu5gkkBG7RrGFVYwKvvOvVmtG3rFfASMz5
7l41ui+mtRS1mkAGL05TSIk2hGnjdkIIq8ssAKskCJ2t7Os4eI+mTHPJxsnUWHIN
62mt7Jk+iUPpYslPK0xYiXATFGhacBdKNaBjs2wjmX3Y4wSXWTbNxAG01xtKk5GQ
uMFpqLuRJod5I8pGm4bAYNsmR9ik7SHyEfxExb2C0u3Xm/eYjahLgcqwTLRrElP/
pGDSu7ejE93Mc3Ptu7JOT1fRCUdmgXCYF09+JQBi9WgTgLZoNUw7Xeh6YADf7txD
xMVJ2c7Lp0Ml1XHhC7hN+jFnOxzbAN+AKjF+VJ3fpiFL2Bru1ws0LJbOnPGNMt1f
F1QPTnEdFBJGSeN6JnQWeZUMuzfCvr5Q1iFx39zmEHZDumaCEZT+gRg7J4vnV36x
tvVMM7nJHWdYaunciu6p56b/LLVnO9dIKwHzHmxDds4ekNIl82e+qFtcC2aa8jRm
ILvjoNWHTtjUVBq/7REDrmD5R8p+lk69aLPpcqSFUWHk5UdhCDBQoxNGMRHpvoWR
7wWYuXRD2RInAp/a8OLmfV2iOZopqfH5f0UrAU2o6EuoKTXLtsNHfwvJtbeMU3PZ
fLKk1K4qIMEBPIcPGR7PfKQ41c0dKGyFyx++ozeicsOrSpPQd2ZP/DrYEX9EErKy
mbOcV0ppyD4lGxKzEZ4z6csS5DUhGT1pSxh9P7LtvnRA9OhfSdMM5tRtwQkH0fMO
TsGyyYuV07u3lBuzY0wc5gr4GafmyBqpb41CYQqef6I4J1bGnlPNeLSiGy5/vf7N
IHya4nD5tZr3cN1VjuHNXF/V+EzpuNBq7TSYonJ+uw1MLE5nizGkRpLfNZHGSVHi
AjWOt73O5QRcEA5QumPQTBV9A/CDwl+XDF9RFHGIsY8s/JiVAASCTJMdvHHQBcGW
pezy6OUE4y4Ljtzj0msyCL/zM13WvXFToz5OFxiqB0+lRS6+vEjVNu71VbixqTxZ
oRJZbAJel0cSzfg+fEnKlcBWpwXxY1r2xROaLTVA6IWPkNASifdhepao19vkRBvc
f8Abp95/0b6IGYqla0Nnh1wB7AO4ZmlqVGzcDePzgFvNHQq4NrDi69MhmJb1EnPY
bQLTz5yI05gbOaeLf9qjSTbqO6Kdn7/ICVuONvI2F2HXyOduK2mN6m3vGn5DBH1v
/rxJRW4eEOBXraOBZ+U3YQth8VzkmyTpFJ4UGUyPhIYi9Z7I1M4lkLsi3Xh7R6b2
zhm3u4VTjPeJF7j+kwI9tJOJSc3SfhMZ256pYeKGMuvUbIRfffxAUcQhCkuOSBfd
/3Tk2UWEoIAFZYPWIka/k1JicjYBbBLU1T+nYXvEu3jm5Ijxjp09Zfdp30Xzuif7
dN5iJfhW7OQusNCsyp7hDopz/Ii79AbGoHdtA7GLUzQTmCmpVxCCBNyexmaEvP+A
r9h9V+NMbS0LQZboa1Svk8pZoVmvGUKeGYsmC6NBDH20iM3kWs1vIpXXb/IvGWlN
9FegoepZ3iXgtRDUjwTo2hON5DnItfxYFctMKV6wnhLYc9b1KOzFIPMAWeait/UI
9k1yhJidygKLuzvGlBPYjIBKvyla8A2DyZ1Uu5U9thBf9oUoIsqj/dpZNa+aaBVe
KepfyYnNWeGcFeWj4Ti3gPMEvfX1kJzB/ps+8/1/2sjtlHBvMEP3StP9dddpBwYz
zspkVHLxTR/uZVL8rl0yYSqmCRxOyMkohKXra1kYlBXTP+XhB3hLcvz2ke2Tntlq
cTltnQIsiWQgB+XTHMrMKRDdtCrNEH7GQMETgb2On/g7MZHjwrkUT936m1mykQvF
xUx31j3sQkQoN//7tg7O5KMB6jyD6/xjz0s6iKfAZexX1Zj0yXm84HJimaqEx1N1
NGEaWDQ6b3lT/njMIeYYV/d6sK6moRu30PYj6tbtaYy5J5de8c03OpOBx5oKAQ/0
Uo4u3Ksm7XXSqzTVgFHjv6y05b9oHni+6RRtWDVPoWXeKX4+o+QZt62aMLXpilN9
Lrjh5BNIFE0cbju7PtRg9LqozjRpSWbcjS12Op8Irv9tsfnbXloetrm8gtPDiuro
+qGTUSpkRt11m7DGM4vTmIgQAnvAWvLFRAheXYyoS1cqgAidgjWh3tMiPWXXg0Ob
okSQMLixiTavjsMDM658upa8Ad77o1jb7xnejg6au00aGA0WXo0Kavd7AfTFV4k9
UwlTCqwXVZl9657BYgo2AsErpJIoS+lbFITgvRFPBNCHAgPKQvE58+cQ1k0oIU+f
JWNX6CtcCjZds3hOByxs486FzhG/eXbbM70f3D02OnBpn64Cak6hfXcnm3Qm1MNl
1NJpzGeHQldMK0yLKdlT+jp/loP1YXwELA/s4LjXJF4N213BA3oPqZtweMhCyamD
hEh28+dQFHKhRErHpReqHmfLftFWj/9M92W30vlm1y8hCBOb2M1kNsWvBsrSGbh8
Gl3Se68kXZj1f5STiX7ZkvW0yCg9KFdLBaltwiOWB/z23jSiAImkHyyimeZC7KA8
AiHqP2QUOSCkItnjerilbNYhgWG17SsfKDORY1QWamP/FaQ6ye/inNE/IY8vV3Gx
488viReMcWxVFbLYHCSLFan8Tj3IChXjKNyPQLPt6bqjVq7Qcgsw3ZtRzghJssqa
zWoHHNQ5nnnktXA0td7nuIHFOEG6GrW2kcouip4gIo29DLAWVsR1albHRni/z87t
NMagFe7UT1EVNCVp/GZuYhIuay4bvyZfAY1csEOkUM6/bDKQPqkRORx+u3BxoItz
28HoOlF2/HDZbNFZ6zUq+V3ptnM/+Eq6h8Lyq5/2Rqr5w5dwSnu8BzRQ6+arm3Hc
QbnKUVYt+H+H+1H/dd3dlnArzDhBDMNRheighJMfM8VGl3htEUfnVvWfGgdXqUNX
60vvkNszUeWvevXGlXsytNUlN1V1KkaCJHrc0rEoYHkPpmej6IDmZsY/iCOaREK+
bYnv1iLGQmEp3hKew6gIKP8s9Ieh3sqnX8tl9XLHkfT4n0zUXxmsvlN3Mp6UIMmF
rs96p7zcF2fxxQIQ4MufQuG5OLx4B9IVSd7qJfUTcLkBF9zU7s6GMw9+E9J+HEOK
OOLsFvwAQ6pQv87RiuURJGFopgiv7C4p8c6ziHJUcPGSM/rGJfmCPwbmdqnwCEaR
Fx3o7avIpBZOkPRbByjMs8aFss/yPzhKSnj2ykdgk6qksC6DTR0xhfEL4wfPjO7D
7icgnOjBnJrOt30+4VInZuN96RpszxxTMaOE0IFFAafMTk4rgXvx7lrOGaFePIz9
U6jP10EuZVtyieFnC03ngjnSevIOnEQeAWw5DMU22FOSfXDu7OoCq9NfaCIFxRZt
tUU/rrMC5dhadOPhahpLk/UfntdetP4YpgACUS03xsLHWDibUA8s3UjNPV2RnCOt
HrtW1BqsQtDTdi6AyZ4rJrPZVJ1+J5I1tknDz8TrMSvBBBgsgRroqsnqJlu1JwV5
db3FNGn8ishQ1AiV1m8M8VSqb6ZWjLUiXYrxtcugeyIfau/4dEQaICyReZvF5OM5
njf5CI3NqBv50lAV26QOvy99BLt9koPQK1berugZ24gq0NeEhSPWhF0EY6D1bHDH
MiapWBkB+9a2k59WaHOh+lwhPM8pPeRG9OUjOHRjvv2M8MAJHO1CxljJ3+6HIWFo
N3tKXqPHu5fcFKheyvWzfj9glX/pmUUTjzmaHkVwC6G2URCw5e7e/jNnl6D1wb02
7HzwrWAEQYzNUEvOAAun0YbbWb2S0Zm/kk/d3KCdQHIUZFnjpKTkGcgNJ+hZXiDY
EF4ZG6/qjwPlJqkiNIpVj6EoJ5rtxgu+9iScn+QpN7neU849iyFVOBuJd1drYvXg
CAU11CUKtZ8WxM8l009d2t1SjAEzMZAscVcTWlDx8bH3n8t85tUIpSYtPp3w9wz5
K2CtRw+aQsAE++JYbubRgQkcBTfKwubn6gVcxw/6NlCMUINs01XUJ8WE8J5aX8t8
anFG8I0tSIapqlZP0K3GMvRrnaEAuSnz0YlPbSEyRGGvrjLIive4g6zaAHsd6/EQ
50Dd/60h1YVtSv0ogUTTrqVmad0wwVEovDnkqejLrC9YA00o1JaAq2GoDPd+B4kQ
`protect END_PROTECTED
