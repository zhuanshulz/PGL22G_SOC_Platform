`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5I/v4uhJbAXdBvQlf34dHgsWvI8qh0hyeMATyHcwGn9zFN3g+uRVUVDo64vVag2g
jLUQfX5RPoAW6G7ObAU6LgE0t2wvGAlatAoscflJ+rudVGIzrbT7ovI79+b48s/d
c/YAXk0mQOhAKKeeGn4ku3ll71x3u/ZrhlZs/SFpw0ez6nhtrCq06gibiV8plT/P
GPfIXRHAjOlMxZo27ifYKBig25Ct6XN0dSw4s1CSp60lOd3z0mtd6i14SK851z5Y
6h+50wzciBeN748GrtTPq6tXaDgmgelTq7B+t8hSTSxoNBsQNpvlocgi4zu7tGe+
14mxu6UirZSxy97/5WDovvcQAusVO/G5wYsN573Q6ytTMJk+TO0CdRiz0Ux7W+26
xQGZ9JPX/7jH81fSc2Ono5TZvoZAW2/2azC8uOFZFNkrsUWFVRNLJmU3+RbxMfjs
A2PvXdCsju7iq11NB4ELkpDCrfVU/nipTt4CBO9IDwblMNQ2lFUFCt9/JtNHd3yX
dKU52DzPQG5EgNQvGbY3wL0siOYpxDTmH8h/kfANO+rE9BfxIPv/F0YrjvXfGlJP
6GtzU2Kf63QF45h+ZV9HuVJn3C6IAKB/c2VQtlph5gqNt1JQ7kgRC+hAUmhArg+X
rmUiRly7kyOgJWqL9yHo9RmZhu+8Dm1Bi02C+F2l/WjPnAZEsMCNTXOaIaKd+PE8
T4TBoxm2fMpTgfgLTGgA2qdvgQ9TP+DF1QgfHFEuksDzUZXIGDriOAxbPMNkpzoZ
bOElvLbskYXfwjjh87saOnIbf9epUGaN1/T+nF+O29bO+aDx/x/Yqz/ug9DAQCHc
iGMXJNvPO+hSbYxinJTXeS0jtUR4bRkmwAvyQVD2VI/w/ZPUc9h3QSmQgdCoW0Mf
Kbc2dxLd6ySq7y08Cntgeij11Imt1Ukc/ch8f2iIe5kgbBgT8ON84gWXndojf2en
IgqBb7/yvZKoZUftBAhhxik3a+j2LJU2IVvcpUN++o8P+0NWE9RCAoHlREW9T1/t
cqy3V7rqyiYduRX2f8tYWubNz157Rc5QGF1+QAQ3YnOeXE2JiRfdFqxoEN8/COXZ
9NWFPbN7IcK/4+NSV7QIE0p57KpGZRQnRlgSjQVqedjccDYKWhSPmpoLGGbEJqh8
QR9JRDC7pT63g4XzrpIzp/orvCxUQeFTSfwa4Gwsskn177W/HFHWzaxbtaHyiIRs
gBljvCSlcCFReIIuCMirDRr3WMeGiiOCRrGU2n8XZUE6EtnP+B6sfHFRvZbXO6Nz
FO3vxD9FgwV42meRK7qv8mQWzJCvso/9wjsKsALb+a4I48jwTBeSnOC7PjT6h6/J
`protect END_PROTECTED
