`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gAVuOQfB5ojalAuZFEUADlCKl7hqogK7b8ojhsvBSyrzkacOFLjf9ccjnW1YOL6j
zr5ZcRiRzEMGmYPuLZjWAHEqQeDm4fkIOvI/0i9B7/ut8XcbFtlGQ0+vCq+lgRX6
HHMGW9Uvs9UbfB2Bqmw73v7lZbJ1ITn9opft8MISzVG0jsVFi3HJyyblH5Z6JTnI
MPlO9HCoHBqncG+0WM75xNlDC3Fj3bYC0GnS/rbS2tGNII2ntOfL6AgNuDHI1LCS
tAYlCxK4p9VDEKeQ47UQ/V+tj94Ez0sCq/H8uHblg5AfzrI8t/3gO5fb5pf1Vsal
nSuLAKnefHnPeUEy5lXSKvgIoUwxH64sJ+HZ2ODgdY3yTGr5TrIbUIGv+d594eqv
mpwMkWjwl9sq5tcoRJeDrqhVEnDcyotUyx0gY/Oo9xJlceF9HTH1Yak9mEhllY5X
LGS6poerszuPR1jTW+cLteee92VyHdlokgiNBBm5FZV1vbvfymospIamCMvIdD/3
GXDRwT9Q0gldhHF3v+UhY0Ey0/bQShWW2p92beCOVSYkKvbEKvmlu5uVZi6T/NYB
2ha5+GE5riwhAjEnZu5z47cpvguIY7bsAiA3R3Oi8jd60ro045fosLDbjDPf3c8k
sKWL7OiVcL+stn2RTSh+tJIzDK+AT3O5N86XF57U72BqnSKobvQBASwCg6sRWS8i
1FrBmZDFAyB7JFHqyw5o8feMkZUZ+hy3HhFzbOT4ol4DToSZ3UgIN9iBSUrlDkKa
nZkmZkScMQtD92N1Pwnyhq/8J4s96xumx/UWYuCXaJJ7nHUKjZK7psrfmsVRVjnK
WrwpJEYF03lT7qDdORxfcUYNdPCuJSjLPK12Ehg+LCa9pubK3vNVWUiLmBk53zlh
gt748usf3VT6+GdM8iRWEBc+KreV9m/OPAHirrk5ecuygA0WCb24kwkvaXU1VIfM
DcJLK5N6SFJrBtbp+Q6bNiRJwdi+SVXK1CA4SdRK5/g8tvg6LeX+Mu/8k57PEXFb
T96Ln1gFFUtLsIDSFwlMErGEuYEJQirtrrpdSBf/k2s3BH5jXwebH3AH1oA/JGZY
0TTGY/2Hj/ii23LrSWI1ua53Nm+Kx7H8siLGeEdaf9HZiqY3OEJfJ/r2Dv0ArTkh
dYR0y7kACMwNX66+g7HL38xNiOdB3spm9zTxk5Opjk7jC1P3CaU/gvHpRmMFf1fN
t9lbbFcKh3pyNyqzlF7RCG/arrZQk/GCyODinSE0cJt2BvI3cMB0/NvVleHxg3x5
pv9UTJUH1uVosKzG1vOlcIsryMPJbIB6kuy68FyXoEokJfYu6zOmHTYvpWw5sACw
`protect END_PROTECTED
