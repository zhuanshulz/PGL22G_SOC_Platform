`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YXm6iaLwiMez+x57CnhPYiRpPOluVwSVIJJNBlmKlI2VuUjZP7URfZ5JYSy7CUW9
tgtKHqFsyXAbaNVZD1XOnt0mipvUMUA0j0YQj9lm8R1oXVRkW4b0NLWC0+aVvFuI
RxgWvmBeUFEwufeScJervca8YpYtplEG34NyjrshuvKdOxHP5YwyBNdox13PTunt
qwNjCYfF90txSBlPHKQD8o5LNr6JBG3DH20JI1MNvnFlOsxE/vxkUTr8R/lHNghv
drLx/iMDksg6Xx7JoffYLg6bR2sTC/gjPjnyWmaTZZlqAS3OGQT6ymNuxPz0vJsV
IUxZP63WfSjWH56GFUt/y+wtSoLUNYpfmmHimw681FEnr1FunC7CUXK9L4STOOC+
9NXhJxeP65mTjCgzQnUr9lecsC88wZsUyoI+kGv1Ba0FT+QovAklOjFkpFCxpK2a
A1Xt5/2+uFqWD+vYqJVc7YSrC0BR1hQnbM9FcbtmRLjTW1cli+JDuMvLX61+JQgG
XVwjmtwpTh5XONYCGvbI0bxeJe8r6M0h3VfKAA0PFr7mIg4TAVXTlx3cD43zdnOx
5rRxT0rmlszg8ZEtvyicuH64Z/zzF0F/++HYapfuuvwLBzJDMazJUXBsodnV74g3
atUt8KJBA9CtWvHVyOCtro7jMn6/xIIVDjLdEKDSLSwPC0iaHwvzN/N+nKBqWsXz
A6VXvfaEdjkWvNjwHLy6eRuH45iQGAwisuWgNsD8BQ0wikyc7mSq797tIeZFmm0o
0S7fJKgRl7sgEswdc6uodvr9GE7M5++vxLwCX2fVmH2J7S8YQ/FCt1knKYljNP4G
gJYxx3nXaEogjxDg0irOzeDM9ehLafe4qrueTg8QxbimMKnjB8lU6VzvDphVwA/0
X5MxYiMygHmoeXtBNFw3Yn3FkyUdmogB7lWInrRxW9rbHQHFiAimZMvxSv6e1n0t
LAr5aUuh80BMEQHlq94YhEdCuhJpHK7IwLPueLY60Wd9n7P9Xxjr93YkYZNdFDQL
j6yo/3sCHZWzjUxCu5gKMB6+f8iXvaDP74f6xM9RZmxKb/xarjfJIm7hiYHit0z9
BmXYdAs42wBCSyTKrYVQEPs7ZvpSPupDVFYWmz9he0ZCo2JILi5BE8YNE02KwnXz
mPrSIopV71z/9LzCXi1enzjuvDrvB2PnkjM5h9OeHE/WHIyyLSy58RSZ+/GrkQNd
oRuLJIffoykyxFHTp+UXovH4B+Tcft0EATg5556TJJhh5CGB3oG4sp5lmVavvkyp
kRD0EHRzPqqZcHGgWYBg2+wajGq05jpBtxrsgklpHlxrsUpcqtyhmfO+fnMTs5Jv
uroR61A8rHJogjPKSvgqOjEI6Xb4Rnwk4zOSOwFllouWoAqTcK05VDAGvjlNdMQ4
L/Yt7z2t+H3dMIpD4vFUIrtlr77BtYh5MNSiOCEp9y+BT8zNWCR/gEfoVTMZz/hm
wFNl1FLqU9xBTt00AbWuVg+gQzeaebayPvnXVUi5Z6xxxDwofw//H18TCJhO9G+F
uqOwA0jjHllGWKVNuXUZagIGAMz9hs+IW5AigUeCBwyRhujFFf9n/cUZt5njZLjh
0rSrxaZmpd+dPyQFR+aR92wEZxdiZpASgdu3mHk8vZs4P0iVH7nLnf+kwUB77m1s
TQXX/NcycJU8Zk5NiwKfMWec32fT0vRJFmqAV9l0BRLVYKFLbWySd/Ev5HclOqS6
tqvi9FBmDoPlCl/axonsCFiPleaHgOl3Sv0QM59ykUGB8uciQs7SO7AWmtrLydeV
n7xFXyoVBure0tU/Xzt3xxE5PGm+qsC+hH3xzgWmzAKGJ0JliqznEOzlDoeSP3hk
882sHc99R6s76c1CwMR+tMpc0BqIAgHdIWTfSHjE2kwSd5Vgip7kklAzGdLYIXrn
0btHO8VaO/eQ00jZLE19OGRD3NAdEpSCpl6P+W0d1ptUljhkomawtqH2VyBufTvH
WWlHpMkOv5Yb0xIAdNBlCljO7yhlGk/zT3BcGXZaZ2xLJpuwXKEcsl/7Ll5bhq5r
UZzBSI3UNauxA8B3XROntoBV/70EDPvp0Ekf7jatNgCVSpBYWS9TTfBm8UfGedxr
KJJAERLEFQ03nMF8SMS5HnSZ4vRwii8fKy79M4RLitaC4Ck1rIgsuSikTNIUZgWq
YEgKg3MTt4NLSJ+Y03a8OYccEH5H+jtSAq6dYMcXG3MHLiP9MrbrXKRPSdIkqelb
zKuWhbu6dQq5VMCFbjzlLm7eSm4cNASwy+D5jTdugpOY9HH5Y6A7+axeOYiClnhk
UXPycFt+DhjVBbEy/6OBqNDkW+UtVmpdNMtwnHLjf5PgoIVJ5yBGUCScmlFl1Kk/
99ty9Ucq19UDQ1Nbq0UaZtrJDWNW4ApPDZbGXyP8sjjA2BpbDeGPHuZhMNqG/Dv3
7hRp/KWuEvmGDgbFkoGbDS6OVgbEwOxbGziWL4hoWTS87MMu63wP9AmCahh+nFi+
pQYTT4VvIC+0tn64lwWdzg==
`protect END_PROTECTED
