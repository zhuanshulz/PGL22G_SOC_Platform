`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4R4Jymn4DEynqFxPtihpK+jTjtE40FaZGGCDLSoM359H3JFX5LyfyRK1/NUBgGaq
VplkfhoO9PohOY6Kfu9TKrQUsH6elX4suUiztc8WkZmai6KiMdFvLmkH3bAZ+C3z
k8GO5NhbMKNWBr7TzxbHaMbB85WWxYCN7WRZgbfaUqQM1qlskYql7K6gTxx+BrCg
1WFXhNjONoW2Piy4zTUPPNcCd3tI4LDcuvhTAEMVBYbRNIDZbdM1+PVpW9txARFF
jbuIJs1fDJcwOKSlhSK5Zy6WE9T+HcSPI9kIvszlSvA/Ka3L1tbq6tUTIXiJl/W4
r7M6b4ujoDRFJ2pMLPubNLc0SEzBldKPayb2Bwmhq/LbjCtq+oHGIKzfzB2zgI3f
06Zf8p0+9R+jfng/YorS7n25/DZSMDdmqEEqgYW3MqRY4YvxSOs3a0xuxER1U/mt
B2D3mBuZQIcWJwSZwloTG8SMhYKA2dl0sFxLb79Keg/605U24gfYKD1mED3l3dPu
myRxLFUdGnpyxk/Mnr9pB8UcstbhQ9J5vEvl879cQ2w6FokRUX8OvbLywR3Fxd7+
1lIGVz1OBrNeQ/NXtQdbUYBE9sJF4vWCTDqrXpzqFNofCT0anq/AVUf2QjDrRZUk
w45cnoLAvpztwdhypgOyXJLzr+kRvWP6sL34mmt1y0YFZSzmPOs8KQ6UK9K8SZTr
cU7U4euF50ANzKxS8PKwnJsCrw2ecuTm5zNawpnaEN/helch22ybv0oTZNTVarb3
R9PHmUBdc91wrzgfYd34WMnAbGwjt5vsFRCw7Vpv6rHA7WjwDy3xSPZBTh65Yohp
nktc14HDR1RMghwhKmpkOcaXJqne8IPyIA+hx5UEbgswDyqAo5eseY+IeGOz7BjY
bqmg6Ns3rnKdbAMmO/Fo0ZbUJTYQzIsgmejlLFMt5tKJ9Yi0RHmXsD3JsgBznmdi
tLpKz9phNfJI6iRGujxsVPmTSwRWtcrKFCafD+8/E4gISRAHfp3cnGospPlcUx0E
DcxE6fSZz27bgI4vzqNAaZORZ3TNEk8WeLZ6bY+ct8ODk5oZ+/T8OTSVyDa70KeQ
YJnT2eutPMTpkUuZ/D+2Fw==
`protect END_PROTECTED
