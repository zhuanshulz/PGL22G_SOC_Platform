`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ei6tPJXu2a3KmEPJaAiBTt0+MdXmcTADMgN7Hq1YnyhRInOEOi9MTj2zb7t9irlC
eqK2nYHwvX1IuW64UWiwIJJt63MJvXoG9LBVtDCiDc2z/Pg8ODCPrIRysGk6qWrc
18kmqhHReaWNF7HjYMUSv84apxkZXQKKwzIU763/yzZgVje6AbIAzfQYYejRKUT5
NH82DLnTMM2DeFRlZitc1oMndAjIw5Gusd8jTOJqcweQIq5vv+Y0W1WxfQJeLoIx
sUFnO1xuO1JmIsAV6yhBBjgpQf9sOcIaahJobv3x7e4+/AVhXmion/oyLU63v/Sb
dR+s2Fpj35/K3cTR9ejbpnxg3S8ln5o5FoawV02PDxARGKxy13QWg/CdFJK+KP/W
v95gRIg0ZCbZebR6LjuYaqyhJYVr20nRGLF1ouqgZIrLf83b5rwHknDqxX8PzCC3
uKSdcVhtpoe/rT3tJsLiFMaxVooB5Y843m7fQaORxO/foJSvjs3AXtDLfmlub5aG
CcCz77cVMXj+KRh50gi7HcwXUFc8b5+VEMdr9X43TNGBuEhdAa0YuR1huOvGJAL9
wUoxwBfAMyBmtVnsMT4GNaf0hfusASqAHiq/sEyRQqSqKCmMr2u/JVrvAMMvh4fA
sIc9Dcux3+AhKjsVYq3IMav6Hq1MNGcimXB/GoywcVkQTf9MK1BfWaSzACUsSkZF
cvyhbjY1lgglcb07oL7EVV9Ih76LkZT90rdeUMK6tKK2qfsC++k1fj1KZAS0Gxxx
Fld+t5qL9TXdAvxsFBCkLpRX0GZoBEC0jpYqMH7xS+BkwoVSSo1DJhTfhzzogoq8
Wn/yv9hZejs8dIdJfMKClIhSjWD16azxo/iINMyXWl64dlKSKr1SO78Hp3YJVJSN
ouq9OdOcwS4RkX2zI9sCjaczAxsR5NqhlWIeSvqHYUTV7oeJDFsccAUrrkay1oFG
+DiG8G4CA2YoC+mNZoF4F6bUoxr3CJooz9Kdrzucoe5BmCLcLNS5ZzgJqug2T1yr
I4DeVxI+BUhc6b4CuFGjExX8zlsuIGUTXVE/Fhmbab+45JJdhxKEbf37ucSLsuAN
jsbeSBfdowNnFGyOhW7fIsNNdcRiFws9R/lceQPGrQF3rfVg0/HLhvOZ5xiK58wi
zdYpO4g2hKutaWcW9fWyokrrGN7x8pPtXt1LnMnuOTpiPvtCMjwJcvMvWdtNihGd
WkJNSYZB3DJp5KE6W2IwEA3zEogMYFLmmn4946Eo43dv6yIATyrSim8pV7M8i5bh
ypLGy0t1MPNuksT8mVEM5vWUacAL6kju+UHEjsDQ0ZnixCawc/9lhfZFynVCcbUd
F/kOSvVZAkypUXDln+68sLzswNsZXmDrzbKGOdizCYCjQq7Q8PBppGCre73mX+e8
4I1c0jKP0FqIknxzy34qT4YYC1+TKQ+kz18hJ9iUTUJ4AFv76vtWlP0nbkRyaT3k
cowdHs9lRF1JIUqOa84V+FdRFrBA237Bh6ihpSgtMXS3Zmg2c6hsCM9gmQafNsGq
aeTYzHvrkm/vlUDmKDhKfQR/qEMO9cspLniHaJw2gT55pHHwQ3ka3N1/0kqBCPma
050FDB4L3a2tVkndzRPcK85zPof0Tu5mK8I7cBlTkTb+bpfn3/VKanmI1KlBUd4/
4HsBqdxaohtG45TvsfUwchwMlXlUKfsiG7sUghWSh53Gd/Jy0VmWtDDM8evmmOlX
rEsjyO1QTH5LqH6X99FADq0buEsVBbkpn236QD5fw2bE+2iM3pMhkFPqh80r30KU
lyNOEAuHmY6oz5xVtV7DgrtgTBXiMnU4q3FJ2HSyhxacn7hSUm/8FeS+5ksiNsOS
pfkfQDZS3Shpgd4b0v/l9QxuRdvpYtCGA4rA0LomrA7htNlTTBsnj/JOUC+Avl28
z9Zpu0mi1Rat2cSxGgjoXuB9ZAkzAT6lB3H4tbWuAQCNrYscnFTtGCvAdfaaeaIb
GeZPq9pT39vf8mptm3jrrETM0fQMC/Ed5GbWnZoenbxbD7NuMaaBnET+JqWIRZbD
grhDOKGnBcSyBWgNk8SJoDNqA2sgfn1OurWpB6k2PjHjDhqfAOdz5rb/lY4x2qc2
keo5oolD7uYsbjSecCSrWfGq030rYN1M/NV+DCBxe6nahvyG+tzTdt3f2zQfi/GZ
KarkVWwJBi2LFRhqQJ7mXh6UtpAsD1KxA09kfsbxfFON5PSK+GCzU0pPoEMQfZd4
Cxz+aXdqlQ6Hx/Dw4c0xfxhKxhq+ogyO7WOiy2j6YWaMsYEFeIAtEyvITQ16K5vX
GiZImLNBelUJy/YSgix6BLNkDyvDITnPRBnXsfPljNSETwhovH24GX3ziR8PllyP
gRm9oOmKlvvrOOLJz8PPjhS8GKLQMgfANqxm8544w9tkpFhT9ddTyGJlWMPNtz2M
wtcN5UHwD/wmMVQQhqb93bGSM3qmxb/cgotSG873q3jngP0RZWBZpnMacr4DKc3W
FcW4mfW68+qmfR+AghGxajTUPAxwuLmPTBIlXlvcxc51FK5oJfPg1xbMk+OQoV6b
lJNf0m+vTdcU1MFJQe5lXbKmncN1By9U57c93FP6i0nZGsDEl7BIOKEDtjw6GnvZ
YE59P9sFlPRNasAXqbVN5FI0K124azvEav2blI/OXFaFRh3jET7KUb4wWVKbSYif
5Uhl+T3GVdxdcK65yIRqgWDpBY+rskFOUT7J8SQ/hnpHAVphtT1BWZnKsWq348te
UT0400KHraULskzYmfcBbg==
`protect END_PROTECTED
