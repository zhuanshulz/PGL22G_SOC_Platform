`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8phA7ng5sulRO5hkz0nvWtTXwDRECSMHf8ZmVHYBPxSGjtKCBgSOy/TEJ3b4nfnu
Ua3qO2HulEilR71FNjHhhl20k/oyN82EvgPfeF65BP3aPLg1tS38UViUMHzOvD2f
pXCj+jhswi6ZWPByxyNUl3f8zGG5m9hXVtTutGJn4pMZ570oyhznsHQbKoFVfCXU
Yy+0wZTX7Wur8aToM8TEiXa5PhvYD/fdONas723l0uYHISImdQaIHVu2UND4xzrC
/6K3q2kYVMQ5RNGq1UQmiT6bg7p4tNTeo76mKKYP5yTdLY/nZoEFioaLO3LTlvAd
8B3Ca9jrvaI7hZfAjOmOemhtLmFhcBOd9mf2IsmtYgfIsEm95458HFZw+JIgdmGy
JQHpFvyvKMP5yfFG86xW+uwUCSAhgrKsepe56XxVPIAOuyBzrAwd1g1DSPa44T2b
eLzFgtm1/tO/w/2p5u+jHI7F2UqJXJBO9gIlxB2XRLPHSUkV/LPrrPb2GtwzmblZ
zZ93aNo5vNStOthO73uKyf/U7x3AHvHLErsLMiCE+MDpFDse20FuwTjF2/8LzLmW
9zlw3MlbZYsn5PKZ4xnpMveRtcJvFTgdps1dMO8V3I5Mxkx4NSow7iv2DvhiH0iX
AJpwucLEpi9ojARcfcjeLtHMAMDZRb0+UWGGkmp6ZZyZ6Kzrrzjw13SM4GhiXlMW
rkUVBbc1UvpO0atuzK4Sq0v3PW9FlIP2XXC3IH+V0JVRMV9GVNtHtLNNCnh7mzs8
ZjOKy16QGK8kxzTF3RWAXeKS0wWTj4J7qujd9eutjiIM50W0GfU4pe2oHXhnBtiF
/fXRQc3OG6cGQFJaVqg0REuflfd3Z6uCCf9sD5LCJJdlblEIVS6IaT8O0EKsyPgq
YqJ3USV85z33Jzo239h2hqH2pHYRsNkchkxo6i1D4DqDTH6JmrH9bG1y5ZDY3W5+
scGTFMMbxVWLDPF/WiF7NweKVLhO8HFADSwk2fx/F1827XOcM/zgsuLaRMx2V81K
mlfGfW+x+qEvAWSrGnAwPuQ2LWGTNt+bYf+W2LPJS3jWyzdPgeMcBNUBW0C+haSk
m1c/W2Nje9ZFVe3Dl4tIomYK8P5f+TwAP2ApcZqcbCfvWhV+eYt+aOtF7P5g3nUm
fAJl3+IBlf31Yd3rSj4hnB0P+9eC74S4/RtDml+E5pCI9g5E8+M71EWucWaNt18q
CxZstHLLjRu1bGw+WQsNv9lvNs9nu4uqm/c5uZNrD9QxMnytgrTq5yLeY4+AWeCO
2SuknOdhz2M+BOYjwa37VSjyOx3STLnGT82d7fES1QghP3oICrADR6W4t1Mk/uer
c/YUHi6cHN6L0bnphrh1Y31JafpL83KSHE9ASjU/qBIcbqbMAn1YTxZriEOvYeA1
X8/KU7Mi1QFufNKgJBYXfEg4r8JL48b2Df/FowwGREmEyOGXJeZ1JmnhOp3s6V8P
BO/3PQT72GEt0t59wWFncPCR6ni+B1odb7+wWJrzuL3PvmkTYCefuvUDDXGzMLmC
00tZkg2NHH5yRxKnj0/CFPuFeA6FYRD69NgVQwb5NH1Px/nriy281mubm7D58Tid
+b0D7vASnhJdgHkWGsiOsZUd+GQaFdLOBM4TKJfJF7d88c5fLaX7eKtALTowA9B7
5XXQPpeS9A0FR1yeR3y6ai9+zHEjs5FT8QBfYm0u/gfYlVf4SsvybvIX4V/UdQRS
v0UinQXF/21PtdRTOaSmngoJ897Yqk7r1Pv15TUupBB6hITMoxJDjFwp4QFPwh6y
rkaKx1mDE4sqNYHedKil2l6Xoi1iPx0PcpHF8yiLgO2Y/RlqgXTU2ZiW1xGGvTgg
aHDGDeQ7wAsf+1lsNaOcVkhHNhVOvtwTWTIyCYu2tEK8g/c3UPNrN4oNprIMVMDc
ytA1YAPdjBY7geA58tZx2a6KlAI8Gn/Zr83u3lPNqkUzFLxcggHeWPfR6vPMsljn
qdmN9yXVR1EfqK0zvnDpxKcBPDLhndHhG4486/J5bcDTk05OlpL4V2MAp9smkF2c
AgQKvBiOngxe3yUWVqW1nkPgmdQ0oMQwLRLdlXHPn0EElWTiIWhd8W/FMMaf3IPK
brbAp+deYnZ77/2cBjU8lto7KyomfkNxw+2wT1Zq0U4F4tFNKLR8s5Zb7TnG7XVX
zsnol39lfAQnShWV+clPYWNV01SgXFS6oUGhmjr8HILRB0YmGVNsQ+AOeCdDUWab
2zi5QXd6dfKrJMU4p9AFV3tqhCSHSBL6QAcGogx/ekl1l8+4X3By9NvIlwfXB+QU
XIca/kSKOZMJOtAkoxeId5yfOuA8Jygi1VRvvWYCzrJ/coi5SypZ409ECbK1ydvu
Z7mXaUnAqwgPaUpY9PZ4U4uKTr3wTaLynpmrRvE0DopOGWYBZYes7mkG4dhdVPVK
7BsbRSTdbmQq6j6pLKIAF1OIGVP5PpQk3NTsyXjWt0eqXd1rMP8lphVVY469ynWa
mwItbq5Ho96kHVXD6Zl15w0SV4oNwjIfW+9yX/HiXcVcpZKq1dyvvvl1RXXgbMfp
5F85+Kgt6ITpZ+28YmIf4ZeonkXfpfWdcV42GXcN6z/f0KSF0Y/juaDCgwZ9GGMo
Jh+cJWBRtESYdBNEUxzJ76mrkJ6bQaLRl1n9rUx3MeFzQkrV5raWJC1RySGwuXrL
fLBbcNhko1PZ2GHwF+XsKhQ1ctEl+9KAi9Z4iYV/mHr7EUAzBSO2jY9/84aPgUf/
vosW+xRAm+w9SNfTywVMb+2toh5AIkdw++43XlVbEAqBYH43BZn2BgYQURmKBBwX
ucuA8EwKXhnD55zEfi9163/3qZy/uQGqJ1FS29FQFbGY5Ep/neH76Erurla4s9Mv
k59Bt44aHJSD0X0wewVec0ZxFQsvYvSzYfcqvIdx4xKbcT2WG2896cqLxRhlcmaQ
Dn7SMhvYksI2M2GXuElSESrEdGt49MryPIUPuUno5eG0fHPwlsQDP/WqgYuNJ3+8
PXQzf7rAyLtdVyEksu4z1GHBg/EiuKE0jDwQpVCi7ZDrfdqyleKUyMdJpj15vCi6
e/mkOyEAO3ZO3C3pvVGcghQETFFbt1N8Bzgzw5yBSozL9TcjGYC3GTShPDsRc38T
Y0M2iD3Z2rPiI4BU2HFjaHJaVSg/00cC+KYm1eD5+xat5Ax3V3pW4lMzpnTTTxO4
DbGoLBz4G6frE6zOxWfeu16fqD2MgWU+tkU1Y/S70f2zuNntovAxxxx14ySXqoi0
cn3vNB0HpAu1mIlBAxKMNzY+qkQyETIEnebZO/pmeV/QhI6ODIZj0rMCHF6KZGnF
F3RDwO5lFSS7MtlqPObZzj/v1lpjfCRpR//ZAASiOKomXGmM262ALNjD5OVVPJBQ
FTyk9K8ktyhlZbm6gfqNVMvapmLqXM+kTi5CdR3t9mPC9g0KwKNwOmqgcUrobduU
WRSletlGfeanWOhTaTrAn6rCPKLg5JdhEPBX/GHnX/6JigMTFCXJnOA/1WDB2Od9
O3Cl8rCI7cahGOTvTb6Zf5vdLWO88K11niJbdX0Cytkzvkwm3VYChn26z/1mJJuy
maaLVX5TKw5IT8Neqpn8OC4416g72ssKqkTCz+QCgWuxlR3IQK/xEJ1jhXYTibPk
oCEvBdX/sJgW7j1+nFC6X8ensKB7zohLQDvFYmnqyDE5YXJv4523Ai2yjziFMkjX
9NM5MivhnY1OnCcAF62yAMHqwR0d8UVFxx6A3pp05GNxdEnUSc+qgWu+O+Wzm1H7
hDoNGn55c0+SFDkIzTRMVwEsgY4IvWqnBZA2H8z7Xn0VD2weYIRORQCvwa5XlYKO
CdXnOg5vsQtTk6yTwTEUzCM569wgakpjtqmp2HxTo32CRzFAf2FfznNQpRHOuJ27
JWpcPyAIohPSvtxpbeQ2/Ki7JWsGrT+LfkpkViOaq7LaUdo/x3YQIcalKENU512h
YRFMbnPIvMbBGq/UN/JwvMYselQwtJAIKRagLAqfwc1eGnvJ2yogFhhONq8tElO1
YVBjxp2DdM2Fkx2U0labzFwi4aCslWKlPop6V8/gmugy8VanQ5kTzbtQ15TnG8Lt
BUG9owBCjKDb11wFjrtSzKK3gx+eglgmYvABQCJm/UnRgDDbjnRvNCVctQbb7kMT
d8lA3PpgA2yBLVrvDcuB3RvtvgRD9WJGhrAKvePZgwrensqg97jFwHdnVC7HNzA4
K3dXwWIyvJM7ZxviUJBruwJAWgA/XVysAed2iPavSIwg3VsiMepAoIE1Qrx3NDS3
DylcpB3uVNel/XifOdwbQKt3cYRKsFtmiCBL3OSpdt9WNN8rebvlAd/ANvZlJbgU
U+B3pTb9T4CIlDM/2j2hlttjZrXFwzwfIaHU/I8IBfB+na8Jf0HD21HIzCee0811
XRrmBeWNscrU/DYz5dtsWBrnO3uQ+6mNVd0P4WHdb0IBXRSYYeuRxq5q2yFYK74l
Rfqq7DeAkY4zdoliBM7l6sljekQmz1e8mZJSUJY4uRo+IvWnKMc0TEf15tehWppa
Kho0X+A7bLbklrUzWq8nkAHKCJy/REva9r4m1/TIBvP4xIlL0EK0EjlxPU92avoJ
OToFOP1WKec2WBixOdES4SDBvxB/IgEh/oL4nar9flDZ5UCzWfirXk0jkgY4MAHh
VBx2bV6Agr14NtR2Y0si74a8Tx2FtVYnwQSJrNgELje9vP+0DwJdzV6xcapZoeOq
EF0Gs/9/dU3l1xltvs3NZDMBNt3scIS3ijENyIEGcYC+zmvmX3NrEjY76oztxVeX
/9iKrKlYFKYmaFG75+QPSHT9EKXJTnvuDRy+ZNFlyhho73tPlDJ5o7SEzoWnpsma
3D2dO6ixH52aRHOLsLsAFH8y1kfXdcNxSFqLmfBMfxQJqEN8sl8SOwZLu7B17XfN
OaIr4cLyF5YwrYwp56uSJYlcejKSoBlFych6ZbSfwbuEbFS2xs2k3Lh4A7g7YPf8
wca4LXSk5PpY/Ctebl7pAqHS7FGBOpux5o3+6O0YVkqaYJdT6q2xUtjXbFxwyubm
FJy7uBKdZp6Y6hts4RiXCcO63vrCHfe8YWzrCAmWSWuYLbdEKXrPOd7PJBtcDgVQ
36GfJDnyXclnBZjibJgU53jXzhRbGTrkV8j/jD0R8WeytzJnsYS+suaoowxkN+uv
Z+knTScazegQXU8dIqG4+t9Ae7dxVUR4mvU6eL3oLGKFdReVkOGvGYRQleHHm+Aq
QcKi9E1uq2hXIYkhaPswSvbWDMpy8COfUA3jJa0YNdLlifrGauaP9/FlZBX9OQCm
gEOI1zyDJZjG0PIhZVjSvTYhKwl6bznsnt86w5JZ/1Gb943qi9+xKHmejgtmSnoX
uXoPM2A514qW+cdzLvQrjpkiRCgBI013vPASbGuwgCHtZu67uNIALsiSD4atfvSj
kWjO9GRHb1DwL7tZVOBNVFcp34gzbP6+qwLSX+fhsoisv9Ril2fKqVg9mrH8oDf6
T1UEODilaOsGOgFgKZUmTbk187yQeuCObjRuar/GAXR0+K6pWQlNjX5GvxPf1ubM
8olVKN5XXLzoHCNdM6AP16ni3qQL4RWJKGyH8feXPiNzHOX2YDLuEB2bZ/mTuJ6L
PkC3eODLUW9pMRSey14apQlV2o4Jdyes4ku3N6zz+hEGS4dYYxCbWEMmzNNcq4kz
Mfs/1KuDHjVXoQ9GwHs8q0AV9EeudVjFjby0u+MBFsuK020rmkiB8AK3zhmm2MI1
TLehDDRJaKU70fvX2P+tE3/jyCB8qJgStMeGq5GOzk/dZKwWtuFvvGOUW8PiyRxG
myaMYzz53ldHkSyFG4zoCxtBiCg1gcjxygOqFFj0uOCnyEOgccaa8H17xigf3+S4
K0Rf8q3syuKtVOsa59DmQoceTlknufFtupdlTJqhv9AtGGuqhS11AAqHabGu2Wo2
PI/KTYIfdxvWTT/ln+vCW1Y2Iw1NLi07B15Le//vA7ShH7kJXYgrmx/P2y+iYYAq
pNexPj6JsrSKeX3gyt1ikbCzXIjLupr4S8nXsJKiN3ZEPDgPg0whAWtedSYa9AjY
Dnag0cN14jagCzbZPQ+yDlRNjQC3u6ueSK9KUZNXAxSXnvympyiMpi8LAuY1AkrG
ZbyrqH41i1hZTkWe8uCwnefvJnacahmVtdzOzNgB36ADccoPCiZx6Hj5+T0lVXHz
mp27KfjsiJjxKLaSWF4iVTjrxtZDSPhfPP67Z2M+kxTlCdKacD/4ufK8WHQCm2vQ
DDNyAlYzlfusYe71r60+ca9YNxKshQYMp2rni4ryCdKEfLPoi5AlhvPeZEdVV2O5
Njqj5kge+OCa5X7MqfLpyaDwf4RmidgTlMsSIy99wQ1zWfijPzubPCrSB0u5OylT
A+YNOEtCj7vGz6cT4ki4lXNF3vVBeyTEAU4n10NR01XS0N1aIjTb7qj1b5C+NfR4
u1nnoEju0AxxceVlgZHfwxSJ0epjHOaWHOGdiEQbO4OpwQhKa/A0qUszASAvlgze
8yH0SodaWydu1VE4khHcE71pH1of7a1A20I5vy4armZDopof6LGdjU+VFufJyHxW
I1hPDSQh+dhdfUpmhe8wwjR0cuxbwcrpRCUce19kcYT5favfRJjk5q9xBinpZS6j
no0SDTF6BzyR79IIERnjG8ZioDakdSSihxFU1FJ2d8961jU5qBK53u/QSjrrpnub
MjDA4a58TU64kgQDBfBinqUniz0p88rIbb7xl/m06S2B0aKdUcQ8J19HeJVBcm72
WwwQH42aouqLHF9p9+9TzrYptnbNMoFujc2o+xAW6tliIldPtjOySCrb2oOOC2ig
rKVpUHusIO08oJAcbEN3G4nMBNg7HYP+jk92gC0LaiECE1Um1BWcUc/B3woSevjO
cu80RfX9mGR2eeJH4pi1eKCR/unv6q114aPSyck1BalNHX/rfs5cobEkFcFk6iys
5/x8LTSCczD3aE4RAgtSJM1yM2H2Y4/TKNqGPkSbiG/RRAkXLwPVTafK+LEw+K9k
06OetFGjsM8NImncqauOhTgvTeh050C7nJqaSg4yu8siMJNZOBOlmQmBdnn9kceJ
cy079i2M8UDsjd9lfQSbz6lt5aAzzoO+PVuerO47hMxRXP5Fab28NDahICM6Xwxj
Bdm7x1LRWYAB/z0MkqoqMYYhWHo4Ucejjive3IRDy2+ATSvjuDzPuq4clt2Ix6KT
rbo3TSEnjkf7kBIccPJoFnFA37OqsUwahyJ4I+ceS8Bi1NY+wgtCa04UEwwqvmH2
TdGJTUy5FFvAQMUEPuAggtIBM2JElZhs/3l2XQ2FDAv++1F61u+/kF802Z87gTBZ
HM1Mp6UpipBr49fbrHFfs4OParh4MiP3juDss3S845aL7BKhuPEdJKKcr/mOsNR9
0SZ6bjnONm4gf+KVnmTTwOWkyvo7vLvqz3U2yYFh9APFf1AQYaQMn2olOSFbgPbP
rgm8cQoXgktXFK4V8BmZJeEqhXPjH0q/sqgDaSsOZnCDWQKJQl+548d18lPcQpNE
N00pcbomFWpgYMcRdX6rMnE6rqdX1TEYkMtkNk6NBZXFuU0fbUYv55W7NTmwRrSZ
B4Fa2gurJNEFjg0xyGMewnGbKMUiJvPK819NsA8vCuJgj0zlT6pKRhLqKUhkMPED
qokSR4KQg9dFkpC2XK4KJDRE8V2RjFRPuYN86sz/VdiKNebaumE9kP4m5nrkgMzA
wgap4cWONvXda35bUlCG13osrh3w6CbPE7eD2MQglzvGlscbbYo012pFgFUAkuNY
I5847Gtc0o8rnxyFRmyypoH9vFHSOIuGK/QPu2X8DYe5eRKt/n05dZoohJimGjCe
DDFgUebLZYWBLa6EEFsnxC5ihR6uTQCusNm/ynacQEI/MRYz7DsLdRV+sxeNXt5F
XsBthJeJGMNTHN3cToNBgy3KLk4wDqeSYspSR4FTRV4Zs4rk47dvzInxztKM8qHR
31+/AE+lGTmV/ebttkbBDnQGApTc45nS3h7pYh3WYqFMk54+7iWjgwjHw+eeOPOv
JBEjHQRyv6xP9/IZU19sVQhFto3ZgQRmd1GYWTD4a5TCj9sdPipZ8ZvBdD8uMfio
CCxa6QZAFJMv0vlR9HaovhwM4Tp9zntDs4CsvT8nsWX9csJ/rTTolo1WcwOMZTo+
AU7EUUZ8SFTAPI8LBviajAOg7V910q7EcoXK6bHvsDdkR5fNRrQscvn17Or3+zky
X4Vv08HT4jQI9B9LFngx2cgHNU+oXjRBtSyIR+T/vZO3aTLYV2lj5hjAHll9kfx2
DtWixyLLVSVNDGaSkFZnkrUl9LUfxP/6pDav6K5LPY3iCdjjBYaWBNx5jbhPRhZR
hZpIs8EGq0/hoImdCpHVu7VW9NJ24fok4n7UeCYi8UI/6XnlWX2WXkWo/nVsCJcI
eD+kPvSvQOIFGH+gT991V+YTrjNR+ewrUOp5y2BpgwtM/UvKLTk99NrxGlspsKep
NMD4HbiyqdVPPFcYtf033biWQPxaDCD4MpCUMl+gzIsiDpCZUR51KllaVoxjKapG
ujXzCek3oY8gDJEGXnVC8i56Vb+WP/grSuAKahJ3tL9xc7Q2gPXJgMgJx32ttmXi
oyAOMOvvm3LwZBcuhxB/2XtUsSgsZ5zGF9Z3RhwCCmQPgTu35A/v+Z33euhcC0ix
zyF8jrxA6yOJ/n19LWN8cprx5e4sgzIiSsFLkTnVDGh6RofcdlGCSzjo9nt8bR+a
1bZeJ6LjEinkHrAp2/bYZSYl99f795NkgsUQWIgkp8sz1xwCWW55LVwWP18+WrKl
ogWUDYtxXcF9BuNkAgISmmPgvkoP9YwHFqsbV9Ocj2ICoDyZ+CgutKiakQ1IgJZ7
Xp0FA+/vKjJ1TMAvvMzYlPPP9g+7Wewqbex1Q5zJbSzpzBPyeZC6CSVdBcNChWia
IaKahyZMbHpBSK+B/iO80Cb43SqX8hdMy1VhHyVwIa6Hs1CpMd1EskRMjMw6bLXR
KqU1tZxE7vMwMUhxSGxxf/gZJnjfUBodkRgOA2GJVhMx2CPa9k1xKmF3eItp+9W5
gnCyGzzSxp1jwxSnWCiX5CX8mzav7BK/H5mw6d05CCnuywMh7jKL+jfCZwo6Wjn1
J5rKdulMTBZ4GDBSRFjDRqKcT/+O6FVro5+mSbJnsez21fQUTx82LYW12StlfWVT
PEo1hlvkTskaTrqbT12V74zMOq6G8CH6nX2FKITNE4vlMPPcfd4+iCHSQNT28UES
+z3jBm36hTGn84oyVU9qHGfwDl2dJTG+wg6+VIWwKLak7BrppuRzAvTKSXUrhZTX
yj9YIHViL1UExI9T3pbMEH5fbZpS460mpAsAs8HnaBo=
`protect END_PROTECTED
