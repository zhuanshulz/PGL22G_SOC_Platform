`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BRBxIK7weOBOFouD0RMZLmBPOmPKKXkUcD1qbMU3J5bBN3XVCRi61cv5dZ1FpKZt
gFvhljERZe+ECkt8n5Frab0HYbQWWf2dXGmxtvtodg4z23NkZZc+0p2gMSH4LA5/
aeC7aqQ+j1xFqhLBveGA+vIlo02jddP6XMD20qIS8lcWzEpgiCAmHZl5jy+96toH
z1sKIeiZf6Td8b1AwmtMiO2ucAAo+Fui4NQmlmch6zs8o0R0mqg6dTRB+Lwvyhln
r4L5qAWwpG+Sx91fzCerz1bqb147f7rqY7RegSqNi2vqa3r0pquylZU/uRplWHSS
s+7+cHBb6GIFDf7Pb3e+p6nLbEmPLN/A++PNRh6c1Pkzl7U7hg9DyLfSsFanFi9z
L74vOd2NnV2U4MAiy+/HIKcNPsxAAAQ6SHvSffK2CBYfxdjNPhhWPykzcArglCUQ
xGe6qYsQGy6ZSflOyiymv57gw6Natzvq9XzvjeqPMBDHRE0jUjKWuGcFLb5RtJNU
6hWtUCe7brgCnn3epprqPnrdzKqGx4lL5serB6w+xhvVoL9kdVoQeG+cFWzP8Nqs
cOUThNnhBAy1im+Tu5DHD0oJo9Muir+P9m9XSHJw9HYaJC8F6rjA3WLrJ6oP0zPA
Jg360qpiUyTvN0IOiQCTPAfKgxa3xT8fn2i+apwMeQ3RV4wT1fMQQiCt4sQmuto4
Zt9VkowtX/0KPeZghJB4wYUTU/ZAaZn+n33MGHpv+jIhdebWce8WZMl1SjTQ9Thq
5OljqPJwvQrTKaRs66/t3K45bw2+Pcpgb6eYvbtHU4CP9onS30Ls1uKd9zl9lb6z
PhM5ypB4yhSrBBYpRDgCJJRo2HsBT20QfGDf0Wpmug+LM1mAkVzVIlYhO+R7h5st
cgqGfEiyWNcEwOwpDcu80PwfZUl01gOCDWGANkWfFmKbQmn//viC8J57uNlWBfmD
tYU9DmwS6x5gka335PkKquNGVCKrs/mHieDECpsRrNNEMRxMFGqXWl/A7lKdvgMS
gqnPci/S3wQJ5JVYfPR1L+MbXxD5XOAKTfN9DzWxvZ//53HQPO4HQAmjWSG1+PKO
pQN4t2hc43X5fgwmirX76LSu4L30ZzbNVxe6p7WhXpJHJDGhCQie6JBtQl6CL70q
0WM/i5uTh+hiFZ4inKzUMDjCOEgoAV6ZN9Qgr7N9R/y8LztyJQrQsmspvMnBV6t6
LqZBdcybQytqKfROUhVtdSwSck81dq9wPbYU8H/S03DHwlS2VzKX2xYX3UyIkMzw
Sp9kK+0Nj9fSNc2JuNarXSi/pEw1UedtrQwKtOQVTYwAaviq1RB+WFEhIPRUAMSo
muFdKGALDwCV9vxjkdaMz4iypRpe9Xh5+d8oYi2TMUiz4diyMZCNXziLf75HvPrt
pyuX6J60tdtZrXt9AJf5k1RCDzmOjBsoeTwmSkImA89wabOTYx8TZx17WyhM+8KJ
CQ810+y0hpplh3wCSOWx4nHwmmBdfrRKbkrNWCLpeENzaEmuFOC94v9Co3BS5u7w
Q5Q+XwAkiKR9aZ+lrM6oWEHtxNdyj7fxlbYvsJffyArWzE5ZfS4tMrF/qWCm84zq
m8Rfi1mBcBR7VIZKlz35klw4m+M2VnHFzO0HMJUbQDV/+eZdQAkDBvjko7g3QQgQ
rkGE29P0xmyyBSZpaQ4SIRyRyTnYNBrtkM97coZQn7xIRv/wpuH8jJ5yYd+yKTc/
pdK988Cz7JCMeEW6Tpe1UQ1Nq4wxN7XwpOTXFrCxxAIkdKqGJNA6ui3qKsgcHCQh
2nG3wykLVl4lgBwWFXNuw24glnbsqRcdmsnHZBJhxgyEneikuBNZ+1Q8PBi6kIeB
LqHZtH2VbR3ZpHaMsIi4pAnjs0rsIXZPXRYBr433txHfNWPZv9A8QcQuRoUUoNn5
jlGo/YkgCkrrR5hKK/XgwiW4JHTGSpM02jlfP/HZmLuzsfJPVhtn8LHVuZ+UjuEu
xWHFzWpmP0g2KBr1U7c9zBY8bfuq+T3wccj9O3IbviO0LM40oKC14rOexoEUxPzu
7x8QczrHUQzL/FgQCIVt4xXLMTjIXEtm1SxFKbZvIyw/qgF82av8/UG5G3LTB0mm
Pyh2BczRHaAOztAOvm59YRewISGWpnC6X6V9i1Qevwy8dnAMSVpjFRYEdTUl11CZ
yNLbi6PamtCkSYCh/4D9f0MwUrTjYQPEwKkm+pBxkcKzPQSYYy0qBwGImyw8Cogy
fZ69AxYGtF7Oit0CN7nSE2FW+cvBZTFmXRcU65+Ohe/rnLLSo4usPvld+6L5tAPA
VtMdn8VwZSelV0m3mUoSGFuENSrd3EMcWs5c8OtR7xYhbXingD/OU9NX0Bi+BaIi
CqGLSb4BF90IOcqCs1fFZHmRLsN9aksCdvCwsf0cVvdOeN/xanNGT1LmYmb1Kblu
L4ecGJjgJoFNjG/g3R7iEBh+CYlIomzz7d7FZUJB4Ku44PjUsk1T+TEFgc0pik/M
lmtTiqWo9nveoFnCgPQBcwbgdGmcNF/thc28DcFecLhuEoMfYBnrA+V9zMDr2C8o
+aK9II4mossGkEbmt6QQWYb7QlCke3MNQYecd8Brum3NXxu22em2xouraJhseI0I
hR2RFYcp3+5Vmz9B5UUvV4KSuRTqxWl73YDOj6fy19vhY/LAS04usAT1qxHN/XMo
WND9ylLA+seWLTswZXnPhNXx0swoctirtIO6CY40ijvxWFGA6Tn99lYUjtUWBIUB
KELkSxDwuYlvdBFOUL4yi94GZ2OQCh8dqCrE4+kZUnebRnSiQoikqc9bo109b1jy
nryrWJpzeMoHlsAwnSIdSe6Rg9x9ALBQLIi0EkEMbbKxNb9Gp4jNaW9f/qnqFbWZ
sVeXnogit22W8RCSphMdZhBBW3twnOGpWq6jH1HrOCmAN6rz1f9rcyv92Eu+oQ17
dT72JsHkgqULfAt61ortGsWJop86WM7EAIY0Mgzk26HltX0A1PPRg3Zd4AT9qUN5
bq1jETHi6yz0iJVUyNZK9JO+7B25rEBaYRoIhToQUTQenz4CetQl532HTvqEWaPK
7LvhtUEtzJIj0if1dejX+4h+FVm3++29yQZEfX2KVL2CiSLiyIiF9lJ6xWZzoRMC
R9VIwwuAGXhE7uXc+LnW9N51rsGcHFsXBZWrS4dKB3WSfsxBr3puE8R6TR5CYiod
QuyV2mptxQGAHMk8wGDA54KwDnhYy8ViRxyakkhFUCNEAMb3d2iw1/g2L97h19UL
xgl0eb/mYEvDruiYbYmkch6QcahTnHBVIRDVjrnnV2cihgGbkCj3UhCvbmImZ6yy
vZU4BXMvfPyGp0bwfSh3QbGVpnjnfAdJVz4Cs/Oy5liF740NkMjp3yhlk4X+9MBs
BbPTEGaOeKq4TrCQo4nracHV9kwrLQpzzf2NtCLXaJf0GOQ7tj33CpPGmdd0HDmG
5huEAH/M+VxyQZI2KiJ/SvauKF2Oj5idza/pKVJ5gC19kSExMJZeADViMzK9776F
uOO6lX8CbpSY7nJ6+eTULV245/TYSLaHop/pTXwLN6sDFHJ+LTO2CUXhnLDJHlDG
KcTT6sZDhipTOgWwu67CIvDtzLrLy/ravrPLR35PvhdBrIMD/NzVGvXfa2H/IAJI
/mqBSlWxxX/tPXznnfXJyBVBdDqc5pUsPmd1peYv1Gdyw2o5Kz3d0hWA2bWRfi9W
7CqVUSC4u05uxOlTtHbxakMTJtYagW8cmJZuTugMFVCpO97Zmf2ZWgR6F1eL2mm7
xyOYfE70HSjg0LwIRmdmB6AjFzGeQUz3M7m5euTdoz+fnkRYprvTvvD58Do0pzNe
oDgxGT0WDGmS9q0edrmO4QbUl8bIvIy9yiq+9zA7HeYwAD1xq+6uPdEhBddSWTAs
9R96Vj8yhmFlNj2yLrVqqsiSryc0pVxUYq8Vw9zM9GyKDxjly3v9kNXvWvNQc6TJ
CcM+Lq+ylb8YKWDx3/xqrT5qBZU+nitSLAPWr6rJuDv4bpGDujYMYAvSTTHUUkRw
vX8tNXtujNGi6TroMUzHSE0DHOhyFIpHPOJFoc1FAkCzI1/RZhhbUChlnKw4Xd3H
a1BbMdIY9j76IPHvJnx5ly0SwNEduONAtbrTuyXBhTdCqfNEPpyb4dUwiA7Y+oZf
LNEt7yhx1rYqn+FOdXVN2Rt3Nmy3/Y/pcZetkBi4qh/LACcMDyRmR604y9T+CWyu
/tEQqKIbXDKifcAh6B4RUHLDYmPJgJgo65XBTpDsOntzseSs7x/8YQAH5tcFlHdi
xS43IDaZ2iSBYGadwF+J8K/03ut4U79Ab2z0OC5/EwcLQ0jRJAp541zxYOKJXS7U
78AWUKJkqI65XUpedRgxPltUjT8MiXi1A8RgdsQdxb9yFdN3ky2s7KpGqcvy0+Zd
ShfE5n2JqohaVrBR4WWTkhkk9KD4hKYnBGxzlfW4Lvkg45x3w9nSSFXgFuN5WGeB
PQXh2rtIFoTTeuTio1LvFjET+FmnvTdAH8DjSuTCnTYzpRr7XoDanBUDitho7z5b
bn89uhvcfdsV3ZiQYQc0Csf1VY7tpqUYAq2lW3LtoMcA6ALkDLG6YSpskv7FjSrd
EOEi//gJVrFah25Vq89O5n1ObqChSrNt/YJBVNOWWuaPCBe7om3AaiomwyovFL//
`protect END_PROTECTED
