`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
efDsMRd9KR8R15i6Emi7NVNQUWp3cU/BOJQhRy65EJnSBaGvPr0L0UhWcAFb8olO
KVSJ1t7m70k779+lERfnjFx6JdCrMsuveZQlZtsB0F/Sx8sozxj4WkI9R9OlaqSC
7jpuIo8Xc4qIbA9ahcxoQ2Qls0i2uXhbRRPAyOA0Xj1EOlEbLPoCkEOotWjJ28vU
Lxw6QBvQm8HXx1XB2W+sUgfKjsCyvDuWT3eNZSkaATLMxuSwmHqiWsMzIBof4PbS
bF5gnTCVD1LeT709gDmfq8iv2BSV4MwI9WQpSjDVWvT/3mQFJBokClvJuzSGhqeA
EzpoAsjUpf9H8eICyBKF11ROAe12vPbV6FeU049yqj/SwzuwesLqnoM3CXGQ9MfZ
rmPWYYjs+bVrDI096heRZVj7d2OwqLw6BGc1XLsZfoCLOFkdWOa8RmhqpVrCkfVH
1tAPezxi0ndc9+r5M+JRLgasFiKDh3GNya0qSeXzus2KGF2a2kCrVhzG1Q6IxCf3
Qk5RI3eCTUSKiOvPSTdD9r1dCNPgNOF2XlnUplCbyLwnkAXRa8RBvDmH+g0bDvWx
/m8/h/M/R443R2uUygn9FtJcj3siMZEmQ/bK7PNyUkRhnB2zaeE+42ZlNIxuW5M2
4YFGOOAa60MICorAwtHb8UVHf2BKvj/T9nczEcKxeDI5eMPxgKN5A0/10kArgiUX
hBM4kyVUV2idA1jCbtsrOWN1I17Y74xxfPkY4+hf9SrpvZWhczeIwAfZhRU0Zc2n
QxZ2qMv9AxUz7PXTBbs9vU6BpkZZdpgjclFaDfFKRU2mQira8XCBIVbchNalk5Rp
7P7+LxLMXMCEJEeXNxtOt9Zh3etz2gPSaNsVh0sUooVbaS7llIR9d3fsoqTySIEf
HdzniLR8g5XHKgEiug/wIH+M8rSbaoG6w27148EdkwZiICLKBH2SqaJt2T2lO/Gt
VSnlH27i+nsbr2pqcT/SSj00jAWHife+eZQeBemVx20ByX5nx4iGeSsDiEaA3phu
6S0jaQkhAa+ZnTkN9vfQSUf0YxzvBPq8CCpaf4Bt0n0I4GDFTu1a+ypmhUbW/o+B
9rn35+Y1lvxKQ2fcvzEeppemtgTZOmiCpk489uwJdgjsarCbbNBk4lv/Vq6QPNg6
uVGY2Uq/tiRIKmALGt9Exb8K0ooAVZERKJVkqDgCnFv69wvkfD/aPahKZOb3ydtY
jrrvYG9l1NQuZy+Ftm17DFsh//92QtccDqx4lUn+BXkbN9R0LpmXeVn57gK+8AOS
RX+tDB/HVUitd7GfG4FpTdfVi9Irdq1i3URVQoNsT2V/kGOtimz6unvsz5nitrcf
DtvWojJysDxavefl42o5YaJRXeifig8ivaGOjrq7skovuC2/ysNpR4Z3RrQy6s2O
KV9DwYzkYUMYFx+5t4IoB7R8fl08q7cNYJxsZaBZinDWmkjSGG7AlwiObK+rfdSf
/bnKAGUhtyz2+tRVJFJz17Mj9rUbljFn/TpdVs1cVU2aFJp/MmuP0fSP1RYI1iue
WkCgVjb3Llh8zO5Rl/nT16Knt8jpdM/RhIg/s6NJA+HRv3rCjHOC/bnn0+xv2u0a
3U8l3UdqK6GukBMFOArDgUgmRRNBE6Hfbmknn13R8pApP68tiu2QVTww1MSj/8b0
NafkRoY2tTTQvFUoJMr/MBzKiqCMqnSLdK4bN+X4ZulZxfg4lyLkcVkZ+7nqNA6X
OoQE14MiDiq9pHpWkWEPj68QBcqBeYuxT1FjbSoAp3KMPUgFsIK8hm/kTsizjP1Q
DkSqfqukymQMI40Cc+krSrZ34fMifJtwnCRutcFOdjSEq0nm5PCyi83R/rs+hXEf
FYK5XxJVgPM0gwx/75vv0Wtbbnpt6G+/ZkaEUtZkAv/TgsLQxDhcH/erxwa9TgHt
hL/4p+0mkMk9hbmIOjki1TKbdlfjEiJYwqy2W23l5REb9O9BVa6Woonoz9u04Gp8
B85abpfkqVurSTp+I9mrhYhhyHUBu+BCqKFOP5xTQwODHjMfJm25o5RxknOfTa9O
e4paBQYbXktKJt3ZYgb73Zhaj8kZqMI/lJn30A/kNjVi/nOMnsyj2mrHWAbiz2Qi
4uD3M2qLiapkP7O08wEkhExjzwY26FIkm4J2ze2RBqQZObDWkL47M9P6vbSHUIUR
Rwo8mNsMGeW6oJIxmPsR9WhagpsNlmz6zjBZVu/0Yo4lJdIhtgRcjCwy7Il1e2OF
0nPtgVbRLPX7aTNkHZdw46Xo9mE0DpPmXUlx4+BLjvxwtDJ/4xYi8cxJMWRmyj/t
ROxRMIe1YG0xb8k465bFgD8yMCCkO1M9BwZ5Wo3AcN+GdzzmBVm2S0smb/YbgB+h
mLFiSlzunt5rVgW2gsh90NIf/F2chqHYB+rrwKR6vj6/ZlN78pL6RkD1F5CY9CNl
IE3hQLD2M43ytCExMnJWfS9eSfVFW9jMh7yO5iQ2/rF0j+QwJPmPApQHcANeZhea
5nBuvPEe0ylfV8+FyqeA0Plr4BsEHnaEH+4hLArblgdmlGPppcJQrxz8PV5T+7xW
pHBTw9vi0c384bSXha7edwrKXoXIIALhJsDtCJdd1quJnV4q9EkDrzdKBDJrpdp4
xEmXva0fxNoCU2X8Rj3lX48hp8vB5tiKTgeMXrjHJzQ4KnaTXIZc+hWfK5MmpW/e
vxJBmBBVPTBAUkYeRPQwEEDauuyO9F8wLtnyhK9kpQkRPY50474UXMvXiFwt+Fig
7ihELNsfk7Ar2N6rXCQ1/+XFkhBzNc+Izx5JS3UzMDi7RaQAPf0Ywiufwfrr/Do1
hGLPXGQVMdMpGLLgMX9gNEeoKV+4HNsBlVrXOYh6xvb/Nej/dt7+W0JZMl50BsO+
DfdePLXimipx6ckl52IthEnscI4y/HnBPe3tyLgJzyMKZcoX2G27/RLryqX98jVB
dVPnghJ7OpwqaXddvSAt3PuRTnU+5QF6nWqcWdoEU6BAJXmqA2Vo5HByqO6nxO8O
St7R/FZ1jQQ8GZONR/olNIJng58rWg2zqjMxfUfJqYYXBagOd5NSZhDeFDLHlrtW
C4ldhU4ri8taMhj9LJgtKSfWZdxBpDWYE9uY1P4NGkuOdAKME3Ll0FbJvoEbU4S2
QFKJdravnymunvHMvlXTzp9TIDujZJUF+Wz4g9AKsKLgcPhew3OIRer+vzdCUlwN
+CxNQQ0azF2J0b3hl2vI/PdpshtVMpHqageWHTJ8aQucwFxQWp25bQVfVs2DnpIJ
VwGX0uqKdgDzag3/4O5yjq63GLlREy0595/eEg/v9MlM7JjS4eFMZOYCRWsZVGZg
JCnMYtDY8FpR8U8a0jCMW7FmTOEFbeDorbWck41INGvDtVa0ivVi3mAPQ4cg8Amp
67rqvfSB20b7juhdfU8BhBOcdXigZeslZ9BVhfevA/pf2GMshIJH6tph+gdjE0m2
nppE+0JQKBCIeyr1x7DRKV/tJrQKMVCrDbEt/nn+2CuZkPU6VOBk6tfXamZ6gJ/J
H/Jgw6jQ3Vh93nlUzyKC/MGUauZVOMnTMWhxOBaw8EwQJLy/YI3PE3N5PfbgaWvs
lM2S0he/rIIc63t3rMspuXIOUMGkL2TrTKb8pH8xGYMYmM9u1Av4/vq8dYtIUy52
nSeIgPcyyAm8VmRVOeMX8cY7bWUtgpn8MBNQ9GOZ/wkF5QGlc+xx5/X+iNNcpR9J
8CaQoJ5w2GX94sxhc1sU/RMjDz44jcGSzcM0QCVxo8ZRD3rUt+TNF4vDci2WIV+k
X9IlBFOM8K8Jdy7WyWUb2e/H+5JTt302GL7KpwC6sucs61n4cO87Wqs3T+IW4xUa
808zzHbTLMGBI7fy/SQELQ8WoMLqpdvq4fF6gWwXjIPoWR3hHiPK3x+lB9tqHbwD
lH3+Qm3/i6dPudXqHTJIjp7WlzD3QUehcuccFLNfyzQr4X5Y33iuaW9YM4hVzyQG
hHe4F38ldRU2chZpTJfCbzOGmmPBLi4FdSoHbHWhNKNqcDP70VzZ+zwaIcR97+RB
sCjmg78P8Anas/DnXSUUhvMxuW0fdpHe0P7Dp1JRNKleLdVZBAwl6EkAmkx3D+0s
BAWkSVOjPSJihoombs5FKm4z4pxu0yV5m3mRMgUoGRrOCKq6gYWQt8T3ZKqc4iS3
ovN4b5zyxmmGivG0NfvokPsz5KxXI4EQCysn2kHPC/6RZu+d0F83P3oZbslk/+Al
ZaVEw5qJZZbboFJPM+kaUgj9u+PLGyxPC3Qa41aMdE6otFtkoxUzyl8dlA2mFKpL
N+kg/sdkuNquHz51emb9AdH6Nj8Csie/HEak69EnpUecvZJJ1RKVc6hqkPT9YInO
4cfvNyj3vMl7/3S1tyWp+Xr7aLqkITNsx4wOqVJGQ0ELGrEXF/9avJOcbXoeySKG
gMkJibr8lCTcKC0qnP2EnqdqVfGyMbZLBeyEk0vLi5kjCbQLS+vyk5xR2odtqvtB
OMdOjZhdyTBiXXUE7k/oiXOHKMQPH5fO+cEWWxbzgbGFzIHuXNic0Sw6h/0WChrU
HbOhbYjMifn0iWeExks3USFyuHrFu+jWSCT9LdiZWCX2fseYw9JwuaVAmROT1YZQ
cFbWFm+BktHmDaGGNd8r85ELSAWHBsqIjSOTkZ36sifW/V3BQHR9qiLjazZYXfws
v4+SbmmucztEegdOxnUnm6ovtfyJyqbUHqATZ4IRLmc6CvbNIg6VYccD/aFJptO6
EmfUIXk7yeowv/nxJtYqHr+OwKFScBJvXpaJPEx2M4EoVcgL07j/W4YunkDxtEQ8
NsGYdp/k5Vd9Zs6JZpxxXpYcNQA/ZaatK4ySwI4ABNOfzs2Gzaxnsh0hLydoS+WQ
sJCpEBXd/Ui561pG8taRLYJ2XIG9UdtjBmdiP4f6dbGgL/4l4d729PK2WkUSBUzs
QOR8hQvE1CrTXpMoXh/CXXpiIKxOqQzloYamBZUSYt9kOi59cq2nMMm0U/iVuibN
usnVIHz98oMQ4XETU7L7tCx0tthlYkIxX2tJ2mIeCfzFfdmOilz3/UwnBJskLcvu
+xnyUXVBtvLpcD/L5VXxRAu+cw3kH6LmEHiLMy/kqJ9yqQjNVMwujao/Conju2fj
wZjEVHiA+NzBZeu71K70OQYM9eJvcJeY7PnjRsHjdkXapJ2dxJ9TgWwKb0ByGkA9
Ixb2n0P93vqZXX/CMNsPlwys7vAAjJiWs+yt7eewYfmEmrbePzxeNeSaZw0Tw6kF
1ZAiMtwqeesL6Tlnd1g8ArdvslUmv1YPLdMBobCCX2m2JLJ7yhpHfV25QNXLC0tR
JmoWwxtGhWGhR9HPmXcgVJyFv6usZPTpFZNLyUu/VYwHqAbKZU/nw4TVTReM3D38
r6VjWO4xwkL777SIm4xzZVErBlRxBFxXtZeCQv4yjiPpdKzku7GLdiTK/IBmceED
Jgt8p/g+0dDzqtdt1+mWFcTH07MsUjN72zRVyPTR2lhpDDFm/NPZ1Sq5cDoeuICk
j/7bJToRy58s7PNAMcH/cQ==
`protect END_PROTECTED
