`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3EMcNlG8cwB2ZIjlFWXejIV3YDTfxyXNwGKgWKKpRCoi3p2q/NzTs+PMMS4h+OKI
17Q+IbynEfjx3ganmvXVYTpcy3QNvPcNVlq00e39mRXhbZMEaopjH+q2oif2lktO
KBDB2jkGa9yEnh3+cbXcXm73amlfVkDSRf6KY8Z3MA3jywh7GW1LGTqTreibZfWb
1Zb26MfCl7tnUshHw2bN6pketg1dWuIzR6c2hD0+QS0bXdZTOfx1kstDPmGKTbQu
lCGHCIipl1WpkXaXnTMabOhvidvB030rthLGG3bgS1gHg+9bEWZDREapQ1mI0uKk
nvMY+m9KRRqbwdf+cA9lTcFSV21GEoWXDPvrHHuKbPluTwvUlS3gYVVAqJCbOfk6
axPMj8GpmZ1676aB4zdaa04S3sKHtci/o8zR5SbxqdjaZ83gYM+iOO8vfKi+muE8
RcRVDNIV9N0A2p1ESwYXpxAnCsxfWAKl0Dda4yRVdoch5WNlP+OoYm/MosFlp1gg
CYFzPXc8jFlIhSXW3a2qBLqoJ6RHMPeabCxb3zM9Jmpv3fE4ZeWSvKa29Hlf1mEv
`protect END_PROTECTED
