`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4xOR+8IOtKIuyHxd2xjtG0yq1k6BcaWCCvmxiWGFPXoXRoA/Thj9DaZDWQvxvdS3
Bjsa9pEu6StNkRDGwhgyoVIJk804jxbSMLjsksj+9scxr5Ualu0ZJkPT2/CUSZBc
lNm9rlmVlJqWC+CqNnAdmmtkOMqGrhfd49W/HOknODzCiOaBchliGZUDkzbBA9aA
P65BIycf6rhIpthHSTXJ1NCmJ6YBTlI4neyd9c7Pk2x2cTMNxSNCvOn7e7AQZ2jX
FBkGfyyMXihybr87OGjEm//3+gZt1pSD4QaHBux6306YgkvMI/aduLPipeqm/t/h
df5AEWUn7JCLfA31dVZApXQ8W0s4WKQlqwlMu9CUm41DGiF22pAYrzV+jKUcVNX8
dCfwH4BJVjXtMRpDvcDU5zl2sNmk4HCk7sdm2gNWL/dRmiXWhA14yPg4AIkwZFL2
aRNCUJjIgoYyf2hJzWxB4h0T+MT90uCTkoAVHgecyYTGtwS9RuWhKMxyvJvXObvr
WmCd5DoQ5b1m9SSGcjiu1B3Hb6g88rYzLxoJQjKXwzpOIBCcUSvS3e+O2+CiRGIZ
vOtg0hwnOXgz9qMqWQS5AM7Idperxlkr75G63i7fn2Ub4WVH5IbLw4Nqct4NwDvU
PoSYNuFt7IXT5FfNFqRgAOqaKiduLBO+JYvnKJ/P9sojvfK4BC9RgmkPFjEykskz
E+/i4z4evWfrR6U3QrNOd5amqxhMhx4KvdtpvNrcBt3RTcFo667AUdXFQ1jCvXan
frTLWxLwXpzgEUHEAZ0wDVjrWjJyL3+pz/djtg8L9iLZ0HMcAGw5VJ5Cphk1WrlR
/lfBfcUz7Qs3gmCfKiZXcn/XFC07qpnJy+KfOm9Zi6t8C8DJsMS9PMxclwn5sdlO
ioQ3NBnRAioxnbL+2RqCn2veqxU1rlwuynaQvvpncNPSsYcUzZ/T9VMi7JVnDH7F
KVc8ZHIYaktd+j2eG69bwTp53dJkpdZ/G0n2doQHgWdm2WnuQenN8pypRsbCvhqF
BQBY4Ua9I0V+PK7FtyavP+qQbuj8wJIIN8vHtrDO4+U3rcFOLSMBWcD0JR4BDS44
NiOIPEN9IAT75wy01bZ16HN/22IB1P4sbqmn3dg46uRtc0LVYGFjQz4ydjK3LKYe
kPPtxte0ys99rhuiG3KR6mklmGrBWHuQ2wlFaLMt/yMYr+eYcDG1jbMbKm6eEZVj
KT305m/HBomXhYyMOXRX6sfIWQ+ma7ftdYJaYD37TtFk9g94WivixZPH8lmrFf8x
Z5sIaGJV4otIcs83lVDoWxgXuZQkDkZ4S3CFxBvb6KZomJMklGTR0N84F5QZ8K9d
btblVD+xaHJpkhXrAPq5Mnu9AQm69e9iNCsoP3WKMi+DYGeYtsSVLaVgmKv8oYyU
OOSz6tbKbfoRU3xwsfg7uHcWxK6TaH1HsKdoFnZMuA8nwgWQ8aD2w2so2XoQFtil
NYyq/JKkegsfG8BmcFO0kVs6r3MfiiDclXhBfUxA7e4j6z595i12FZ48+6gQ4lO/
7/fX7NKu9b3fKDcgZaqYOvbUAOvE3LyeIOBcsqmh/00nJHn6R89WR0bLqKFweS2d
Xkg3EpwS638gtvcUdd1mrOleIGlti/K13qEcvkBAHgSYmf/Kx1oVC0Fd/UMOFIf7
ZBZrqicBNuaBRkmJ9tui2NqCMp9NzD27DzjFN7RsF5iOUy8CzbDgGcJmmod+oqOi
Y6sUbdr8hEc70xFsCH/H6ajNhhe3hg23/qtb00QMgdkjTPi9y++rB4ZSg/WzeUO4
tSxrsDYhUsJJrNVY0jK2EDylTqVpYWgmPDSarvA5Si1kYTpqu89D0ZOtMJa6b8a6
qWDnTbrBy1b/hm6dRiUtIS+/uH/yECl+AhLZtM1sZCVkJ3TRRbxl+L19njXPxZ2s
oPnzkDb9wi5e+ttWUKYy1a+B7fWDWF4MiQhaJMmUi2HdIPO5MdkR90tHDUbGE85M
5F0NQ5HSUI9dF5eDZNI5F6DzWZRDyyg6WeKPfWCtMki0lv5fUHfq1GHPV7JWE9c1
4D5//BKHF1MT5aGihl5SzhTzuGi15++La2VAnOOw6Vi9sVULQHGWDqJe6m4L+3Nq
MsNyswDiNkCloiYyhXZY5NR/X0i+xvnsNZjvujyIuR4tvYny6EinLdf7zyybqwQd
VBWZzbME0tC88st8cHkRkHCK8M+Nr2xKpsPXcnC8R1M3udeaxQUPfL9OJ0aSGOW3
qub9PlWszBBnIjCV9PIWg/ArjqJCTrLasnApArpKMaRilH5F0Nkb2lsXRbOypmyx
Mo3R+EJlBkaMcKW9r9FLd2bMFiLRkzH/jWXCMIomKhr7JB2CwwlzA6pMhX6FeonO
WXIk8fj680zXqCjZHZWeGk0oI3OWJI+7O1Ew68KpVMYihb/sUmYELmJZt/TInSrA
PTObqkpTUPKmxdxkaoduScV7UBJ0puRqnI1I8PTWHTBw1LhH8MLglVsYP03RYPp5
TaG+YEY+ia3bywCqG6gs4JdqhmLbDMmw5P8OoUBPhGLeyxj1rMRzNTMjQwMjVuN3
sC/SGrRXVOlEHSYIJN8SN4Jp7Lv/ThwRaUpwHA8vbo9eICEQvhbTPF6TWvqQPjvS
hq9iNr9HdWmtQ2pYJ4Q5Klrfz24biBONw3gHDzjfZsuWTjPr/5a0tYFe3lXSxi88
lSijAVW3hMtskFmzm5yN6cgK+COA9L+ezZ7SKYJg6ANS6v1OgREnWoFVZESuwk4O
iwj2QOjGIszd2VZWtN2sDBjPejrbeBtoAlsg0l81vdWrr3F5fdAcq8y/V4/tasTb
bv1h96mlEza9q1F/kf9CRAcQGTY9MnSfrQ9vuXw4AxjYsyzH+pevDcqjZjt33b4q
omCPownxkw23aFL9/LN/yPx1I/AAmorEFe8LGGLPLAKgyJw1zb3MMvna9rNAuEK+
GdI/cJkvmKEi5MZckbNWB/0XRSpJZykPFa8QlQ6RV+VEQcfwJCWFHvni9apwZuNx
05eeZsHuXVnYGoGVkS3X2w4n5HjRwkksHdSH3Vslu7+1Gol1zlM3ViB34POs6aJs
3aN6R1zjxU7xaAVgoFGpzmMTjEfhgVgxSbfizwoTFqNmfGnQaJKK2SZ8vpWPNXBy
1HTG6m7W8RbIQ8TPFISuJ/GBkUxA+lckbPMajmLu8tO/gpMQIvhS1ulD3vMi7Qq9
TijyBHh56x/5hy0LwaGIydQkAlFmb6IlSq/J4dA4Zgu1EvrxkBrUGwjQw/7SI/XM
V7LPelOSNk6otnq8ySJO9gka8BuM+sMBcoimJ1HCOeafCsHK1AJiY1wy+jNHnHC2
xbEkwwe2ckvsx36KzUqXhDPB7uJFwKAvQATGnjvpXOiGcR8EWqTGsjqQ5q3BQ34n
0v89iR+n9b3LCPMw/FX9e/qWmELJpJE66bO6pqZ0hjOszExi8ZSMotxLMFyeuGCN
RzOxnpg6E5LVH2TxwEcBuxGcsa2SKTrsnysILK6fGBJ6xYRAaPm779q5JTwKTwu8
+f6LzmFKavhyYk5U3wiqxLTfyo5QfgwTlsmIZYNVwXKORxuc1uCl15wjQEQaNjYF
aP9e33gJdi3ABYvm+yHCePe8T0umQqTD25gD1EzErbnpiiSIIBfykOWjiudRQxU0
h/gdDqu0mjM1M3y9HABCRC5zVgElGoddY4rwTrOE0ho9JReJiw2RuZup4jeBNgJx
hGh2drcAkUfjcJPZc7PDvCeQdns12Hp6awqpBsekk6jM5WxiLtSkJukAHJQxByV9
urm41JK4gUFttUWSRpWP6q0+1++tZKXB3Fy5FXLWvga0PG85RYwD6wBZuFz4+l3R
Bl7us+keOJZi07v0dllR0O3xG2pSkS7zg0AFLEVepOZ8u7xOMl0QS99k42d6ZurH
uhx8O6vpf1FDm/AP+smDvVJ+qk5c3avrydADBiGMlcX7a2uxmjsecK8Yzu1cCqlF
7Of+gOkca90UtaKoEdCyjpmB6iOK/PBVh+mXupPg9o25h0sCrD3lyhgwE60HcLrU
7V98jHv2LDa/0Oavnxm/3wP3ryvvNSQ0nY/lPsme8aLWeQf3FnqztPuqlJpXhBoq
XQMIhAZ2on+x/vg5a6naXX/tYR24y2WBod/eZqeAChdDqzORo/hi1n95DifWJKF4
GQvfp5esZe62a8J9Uv8ZR4Abnbvl6nk7UwepgnpVjL9pvS2TkNh/SzJsvboZs5or
uR8qo1eBv1o19zCJdLtQ1eXQP7nSkd9RFb6ux4Wf28NLWvWRIH+lwl50r/o6RlIW
h75GMtpWYA1VO3mkZ9V3iFHeNJRFQkSj7jpXs4zrUkGB2oKyqYfgwObDs+pnteie
YeSsz4LhFyfFyQ+xBs2QtK37aGyDFrLNVxIXGal0EYaTxAKU05w4Y06JJGTIhcWw
SBA6mUyN9ftgJ5viKbcSySqW9yk6C/r9X4v5B7XL0AwRcMP+XhXVXa4XpszqsfSW
w9Jlpj/Y/muFeqZJpxanj4tB+0qN8r/sOjs2XzN2Xung4OaLxO57kxH6a0eNli+x
YSTX0qixmDHSqDvMEoO54TaRWhURuKdYkpz+fglwKKeBRS0WZYaDyWuOcFdz1BZw
O/OzB1M5Q08KTk7aj2ltf8TGkfamOZImDyEc4ae5qJrhjg9aTAd/IWZq9k+O8xrc
kBpapjS4GSrTHjnqvp5JcegK49iP/h/UdnI988t/E3vPafB3GhdZXQIm+kfwn96R
FX/io8SLbhfiM2wJIZrDTyJ7DvghTMff+siWkB3TSzoSeKjz3ygt2PE5YU7h+sBk
HqdJrL9XGE5Jb2sYxrCEkNcSzdpsTm4pODJ/y3O9smTxGs0HyvvZeLbU/e5qx78h
7lRcco+k54CQXk552bFIrT6exoJduEoNZvaEU/85pzsZzcHWbzfzcWeXrvs3bSul
ImMpCm1dLeIYt0TQIhHUfU3IWLKSB4HG4jghaI03HRIE7R7JpK0w/WxQOwh55ZFx
kbkCLgtromOEJdgfSW3mfqR2jQLenmBGuHSDS+n9IKy6/bHbe6o8abltcKfG0uzT
Gd7aMWg3MssJ/bGkJKPm3p3uDiYA/s9TWCJdaSDFM8YLVTuLlPRMzz7Ah0UZXsdW
5hEqNvAXOcQmI6HAfBszlhOMpdE2xO9hqVP/L4xCAFnDHUCdpqgZ6mcU4nUa+DBZ
V4BJlk43r67LjVFKgv3ThL2JJ8sc9nNgwQ0lsegyoPuCxxpc1CR1HxLvO7JmxPGs
pKLfsXn/lVb3Fe8oACJvf+1NDlOUMN+rAu6kBMjJuj9OHZDjwsGYQUPJr69fI00H
sfuWvyuAtA7b9eKoia9opH/l/n5wH3zO1tqKXjPdNKHRbFNe1edIIexPFR/fYIhk
z37LBon3EfHLpVcF/EaZD4FhKaRcCygIbtX3VlhuIMnQFan7XRLtgcv4aYIFcCLw
VVJiz7645MF09v+BgzIWQedRIsstyJInNFf0EckoQgiGQFoRqvvU7oerB9C4uGCP
hQvIxJ5xAU9QGg8asexBwdvcU7A9aqiVn3uU6gNXG37vCXnQ/jCeWy1VYl50NHnY
Rwp8LkGjN1O6uV5CQjefw8Tek/taguUCddsDWJDa30t3/RXYAiOepAy/yCKfkp3/
x++65ORVTjf6/xDkoT9PPYi8ZBvdn2Q1x25ZJqq6IW0ZFAqR8iI1E8XiO9cnKK6I
fbVJl/N1jkEbW3ntPeouCnecgeLf/ZjOrRu7BFEe8yq5lK5cAHWEvj2jB/gbo696
ZNLcSGAbTiMGR6Bwz7Cw45HBzamnFfXQizkCfAi3Agfb8WdY+6J6NMfDJcUB27ri
w2sM+lTSqRiwPzQOsEy80jT/I28hF3uXptzf1QlQ7K0X0pOgkq8pp467KG/1Y/CW
jgQogcN8IRTTaKlVSdWKvcDnpLc46RcmH9w8lFwcaqVza4qHr95n2XqCZ2fVsffb
H6tAOG3rV9MCczZ8v39ET3n5F3CmIRYdb9iijrxSmqK6RkqDGTRfWRSkBKyhevqT
B6gOGZdb46bw5ncYZqJUUvMPzgRTyhtnxqNYU5OUSi2/RD95eOx3uutPc3yCLkHq
qvZwE+4L3EhNOANvVWEEW5dfBl4tHHiEMWqVfr7FjIfslTmog0wNrVibX9SCaXZh
S/540/quV0FEAVEV0GlqqIKZ1jcS1P00LNm6ODdZ/Sp3o5ulVoOEsxu4EgBazL+2
nBh+vFvvNbqKBXny/ANQdDKSr2e1o6Scuhtnu1cOGAeXG2Z2B0rxa6XZEnCC937D
aWcty8MNtWwyhv1lGK8NYSi6hOioWtIUHThR4vcuZYR7j09H89+2yP/+nIUZddcX
5Sqpvs673O5qYvKynD76RNjAg4tiGSuc79n3gF36j9w4kDKRGzJUq873h/5G0s5P
fHiquvaT7RVUMOJO5C8Kkd4nKPhG+NLdgOukgulbNOzhGKKZv0pL4fZTwFqUCKgP
wBNgWtYodMr3fCqISPFlrD7FBDXcc1zNRGJDKvzLE9ImNo6e1B/wodChX/lIoXti
1+qRUyqCAV2b/TvJ2nWegYzmpcy9w/nMmz9OOmiXBdx6oOf9ieVPP/xpm5z+BlwS
e7LlR/vu3FU/j1tmU4iMDYo/fYtgAdQ6nRTU/COkRU0FB9sra7R/w+nZMi+iRdAu
es/IQrejEu3ZKGupkA9nayIraaXl12JJjw5nnqNXzY+kg52aZClah5QOaoWb7XQF
Ouxom+Xw8gyULUk8nDLX8S4p23H7qksaHUsnOJfddr8C42cgWXSVbzAz/0xzuNyh
GfVXZ3TKk0NplyGwSpHR4lAPolT+G15/9MWVi37IGudoHR4NLfJt6RYqLd6sm0Fw
J/QdFzpcmJi8FY0wxhzBoPwSMdbA7u74jNyfnOYQbNmOBeYX2zYv8SA5vlWW1Ae9
nliBp3EkhOEHPRVhJoWeYTFNN4BSSKsVF6XSKOPTFmTELmY3Hfv0srGBiRxy7GR5
dkt7xagTzp/6qavW3YxKRzDj/DA5WxhH07BtqLlXy8IRjl+HsYADisUlhMl/DPIc
o18mqzC1+68U1fgV+o6CsBLgiN2+lLlmbueZXjdo9XC3ecsYisBfxcjaK9c1zQcG
cvlSLVoEDqM4BVIdY1fVJXDvhJC+Ttc+E4NyklgakVtYQZDK2igQABGYIMf01/vv
O5pd+9xzktQALhaD/4om+Ii1mfCUtgm1p+3XOcLYKjXr3iz9Acg7lmPAPCapdt8x
tCdX1fOqVoa5dBtLSr1jDElQZ5B0HH2ttfCGRgoGTRnBl1VfuRGIfXn77DMd7pUl
d2Q62ljWVS8Wgmz7Y5nw7lmsZhCIW7BS4bhw4/KIePwcDkzF/RkQBkDZrpeIpbq8
WQAaF22nbecHfIRTmOj0pwutZ84INCGbGNI+sIjYRvOYVpTbxiRp8LN4gaXoAZo6
kI5y9Z8dYa/Hoc+4OYBWeq9Ao6i5G/qLe4it1WblqdyH7YgEgtOcxNyYAKKN2LSg
TP2/Yk2miQzs/CYr9Z7DO9YLrCQGWg+iVqh5bj58qKvZYa2r85IKtkGxWUM3Gz9S
+kP5KvJb7qs6FjtFRFy550+bystPIZxZPvThvOsY2NiF8Gswu01dxXzgYbyEI/Eq
LzJKh4ve3u2yDWk/hvWmY8msYdGWm/FpxigwUMyTnYswj3etg5trRS9zVcNPO+G1
dRPtCHaRaZA/FeP188RTCa5IsuLUMzhWP8MH1mzh4BoyTe9E1hcT+HcGSrSv/PfK
Kbtd0NDWNl0dixW+ZJ0J7axCJpPN9cUXOugnsgIMuMM31XbebYrKKJ7jHhGoXEhb
Dh5K8qJlwz+lc9Ov6eZE+uoOHls5MmEpBTlAeRKDgZ4TTR4x7IIs5JwJwBRmn++s
G5S16xsPmKPMuaGklhd5zdGRK+Ap3Z6tA1085UUYVzVYe8/UYxR5nuYB3tY0z/hA
BEZUR6fp9RHuWmyZIHFyzZIn8NRQuU890PaYwPf9WOFKk63BieLb9jfiUjs8Wfpw
o+dlWo4KO+GrYV+mcWFMtk4FC7LzjTZiCklwKxrNZsw4WLu7UG+dq2uFioYFQEsP
YYYgHwPQg/uuK99ZTjwbVzIy2ikkij+3fdmE9mElegyXMrqX31gXNYYCTozKxdfU
KbMFkidguoAme7EmgKC6LWRzW5SCDwF5kh3qrW5myUeaxH7RBSAABshSgSeYN1Do
sS4WFGQVYSUYH8xEsq5p+08gucrvPyqMbq5vbdXpv1zHRDlXrTPPQRlq0Od/WXbS
axnqVt2I+swAZJqKtUr9nqUqQjTY3Y/vhoSeK+YrX2qgOeGZn78gFARiGLlVrntx
nRUEOMSloZ3u8Yevo3PBnCmkvup21cDbK5YA8ySB07agMTk5aeXUo8FOe38++xzk
ifsk30rElxIcFNX7DpuJOqc+5ErHBZVy8O2e85hO5yOhd8eMv9bgD5CVfbbRs4Ev
3ITm4C6R/6HH704Z5AgobqXy4HoauyHWG81Kl+FRInbvQnVAPYnULgNfXlMXWEPt
xCTbrdpq9WISCIgeLuUYcuTUXzDAWs+kbZ+ggCJqZ9wkH6bp++bk+0m6YQ+DNi0V
XME4sfQ6veGatt1SjILenTUN1gAAb0BaFtNiA3e++4dZMO3pdWuTvzgbGYm9efyG
O4qF58z2hl9QCC2tDr8iB10N9/d3BufJxaY2fwRJy6bX0b9oiqHIc5fDsLbIhabA
5K6AsKAwMcNrisYkBh7VWl5JIMk8bLrpDntyzw5JnxRCDNkrzTZJpOq6QVHzTFsU
3GYPOmQuIJSlLKRaWnQCeItH3dP5YFz5eBF+JkMATsIN+nHAm7i/vNrtzrXTLZng
mh3YsTCfv1JeBtzvn98BTlDxS7oOWRpSwo+WFFaIw+G1KXcxMRn5BldCvdpQQ39M
RBEcl2UmJfb2mzazh/1AvITCMLhFO4T+goFnUjkZWWVIDMlssOPv6iqVsezX+QBZ
beJpdbtAnE2JOHkhvizmu2RO+olzSHekRvO8L29XqPkxQO/YUBo02H14PBA2qrLP
nN9R+EgcT+4l+yBkhdoHhAT0WGl7JxUjsiINA8KtX1u8vwYQST37FwjpF5gxMUYB
pOU81H8uDSsdU+SzSvcPZ2X/+SeEG+x2sXD35iWdbGUv9P6DZdtjd22649TMvV+W
mY+Qg+uA8xL1wo2izvsJP7GcZms/SijXAC/HSPsse+0=
`protect END_PROTECTED
