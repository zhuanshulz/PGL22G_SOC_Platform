`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GLOqN0n2tz1cIOL6YdtkUJ7Bvv3P1+cs1CPZW9jte4PCf2Jtja9qPEDN36oUi1UT
aeyLg6kGj5HHeO01CTXbXGKxca1hDM6/tdh/cpyz/xi6AFpz1ZGl+puc103oCX3K
+vV9BOofQlQoT4gU7N+NvFX6DwHgSd7F5Bn/jeMOurNQGyJWK2nWnsRXzM2Mw09J
71tx6PNhnOHE6xrIgkePefkw6F8kyHEoBQg0lOj/EYid7x3B4c9EdIkOB2Q7l/Oh
ilfUQNIl+QCiVNDRe3YXbHFLuVpmUAn1Vq/mUwvEE7+r1NLlBWKC2ZYvP2eeNYrD
7HO49B1K6zO+vnUdiS09KmqwMY9B73OUZPEW/Bv58HAfRTKjxk0a7C4cvYqbLfaR
vnppjXy1cxowEsBQI8dEgg==
`protect END_PROTECTED
