`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LzWrr/lhTFNVV2cjPduODqAfteX/rDCPm89ZO4pOOte4fIKiOBY/eCwukRtpABu3
eaaRZk6N7lqPU6zknSuI7hkK1DriDdsOwKf7M2aeyQle47+jYgWnm6nrDmTFDsXy
v1/+8NJHDL8Ni0ULB6UbTtRKr5RjaxAVimB7/OXd6KB5V9Y8Ij8GUYkFy3c27gVB
+AwkqMBKaOZuWn7TER0KYviUEqq/gkcStWQDi04TYT4lmikThbMQx2f+Ydc5cUE/
qUqh9M0UIfGS8PsgJrEnZTU4ItcXWVtGrvHh6Yb7MPEXZf8V4VY2OdSr4MG6ZaOt
oGx/Cj8gpuzoBOqgEZx8qkBXIoF5dfILxRZAAfk5zekltreZkJpCFljQhGAw7yu0
`protect END_PROTECTED
