`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yz96bBvy5emdKK+8TXvKbkvWNsabQSvzo3irxbjTInMIPT3FZaarFmdTx8qtbsea
QTjKThXiBudwliXnKSCIfU1iFWSS47ZcQcpAkImMZxBO6cWK7hZKJLSKqQ78ZXVO
1rG7i4RCs+SaaOvBz12WMgtF08EnkaanBF93ApseO8KnF2qGunBsevqPdOZlIbUG
fEnRd3Tqn8c9GRzwoJNYXFRIPf1Mu0Q9EbL9DyAvlEtvtO1AQEpEgLAXH5f1NOUZ
gzYUe02/ZPLb3OrFM6Zn36UgwH93cC4c/UYBhe40g5o13RjJBWTw7WbzAyBg0Bir
Lw50pAlvCXyITREERuyq7BPRys/7wkMrWsl07fkOhWJm5aO8G62OFOsnIg9HcVCI
yo/OEKzOtyBJgemQKWKCQ1vJA418roIQLSGvOzTTp4P8/W8ZFYXIf/hSN+haqB57
TgT5AN2ku/lEoUc3kg0WB1+6uh1Q29eOdXfgRr9/zulf3RhzoyLA8Utp5KDZVc2T
a5ewSR5OyCrSBSUDkHRWHsPm6ZOgXku6c+oj4LxQoiGtvzogjX14LeLViPBvLcI6
AvgreQbbC1re60GTVmdeT7eHeVctHfj7GWpHUiU00msKTP4Y/HpCs+SLWpQc7rqv
gPbVubzxZKxzeVOb1ZdEsm2tgcZX2dXch4i7j9TAnQgR2eqDlE/k5ZQRA+KvcQuS
0d4ukZZCNhyCTtnROLqYQY/7Gn/QjXJOejz1jJnDpMJl2C2q3Z3q3pGKaXX4rwfc
QSuqeVtZxdnTmOeKj2EEmq+7gP3iLbvgzp7+wz4I+wPSQu6SCfMZcuPzCew15w0Q
GZuWJSWIjOcimXzbqgvcrtrjbCBRAT3CysawULyXhi7COPstlZIj+7ymcV/9qiFb
NToEPQzJal9Np0xR26MC6TP6xobN1ZSKkFFz3x3x/ngvXwbFigufknO3Xs4NWclj
yS28vuLnvDqVn9JTru9+zZdbhbRdWkHONztI7qIeHg3zE/3qkXw84/2TM70nqNQd
qploO2wCgzjKrEN/VkIVuqwXE0Bk4H+XPUaybDab5cn6zHdWlfEIp3o0wNgZHsv7
J+ePkHKDPFZjpJheGCimP/VXMGLXZqHOG2VO5k+zYXBRq2AU+9RR0qzvCiPZPYe7
3eYGIUimYwKoZ+Bg+3P0VLexRGW9uWSw0dofHZHvTZC/7yMc9WYjR9e9+i6UYJYp
SydqQyyxocDTS8G15r9w11ArLEWmHhPQfyIklJ/U8Mbxc5pu1dC+SCpHx0C51UaN
8+imKHp2YiO8waldbwQzNnQyBOn/x+ySiSDNJg+IfswWcruUQUDJ3M159irx1Jie
laem7VSZ2N1nGj5IdCHlwmdWP7COGPIrO+HoCUAM0CEzv+3bFx7OppeMwRvnBDMu
dzG/q7UyAy4Cmw00M77KeY+/HaPy7qO0lxh/oqLxtA5KkfMc/TWEgFSPaBWj4H9K
+UGF2UtM8+uYLMY6iA9YNpRDpeXbje48kXvL9Y5Ci6Bvj2hz1lG2hs3nkAAAwplc
ajjV03zk5ULK7KXhFs/Xk/vNHWRACiVfLziqaQ/Rub0Ynle5f2Oj5obdcBRaB1t8
evgyKElKhUBQ4COgS+fKKdqrdVHyzEqR0slJGZobwZ3CVGD+OHuafoZzm09L8U09
mDt90qy8SCB7TNyxqCNAPYzkyiiWzMQ9vZ0FR0nTLrsK3QoRZ6gZa445anc/mS0y
RHndAqqTdbpBxB2LZEXTS6r2rL/5aOrFV4Z3O0k2nyD4aIDdmCaiQlKjdtjboqa8
2zeNXSXfjH5W4/7umNYPvzeVSM+QwfdiamZW+vcrb8Gqh37T15kXI0xvc6MCrQuD
ZSLUdC/9lrWu9kfu3T6vsXQEW3mZA3a8IlnjJMlHu60hxxD5yKzUghUmlApwgj5/
rVH1VQWKT6szyqPE3I9af+OH+wnzEWxA5KG3wTEF5XiT2sQEAFYxe4odi8ygB1gd
Y84RUXqN3DdpM0tjw9pTEaBcxvDLEZJNd0bYOkWuDSzYH7bko0BSF+Za8PpdLU0A
OZPC9uqARxmPwxyCqPwG/moCsXLT08mzLgSdMrMsxsj5vLdjY6NOhgWIAnmZuhyw
89p4y0nUWmQCXiGE4LMoIQ5HxK+PeCh42w3yBGMDfAG/tWTlHVLOhnU8YrJQCdiS
Y7Ic5meY7R+tE1lEUNMjS9uz5NUZ5ZUkiadpgPEwCmWmeIIA9HqajatTW9Ve0keJ
r0IQq4oLQfIshpt3YfA59/xIekdc7xcpQb0wNyQP/b+BC3MslgfqKexZsixiIt6I
Eu9bTLmxSVRGob1j32hPMTiRW7XpYY1LyT2WEJU7oZ25adoZs13BZwxT6tlAx01g
TOk8GwNNnxMF+WYcqyLlnTEG07VNAYKfoAvGa+VDFdJON5qg7fefFjHLyXXW2fdf
C3MVZspqNUv6FyLsH+CEsTIPx2rGLbG5NLzfaAJ44CZ4y8w6gKSn5iSd7pBEoL5i
KfbVOncs/ErUhnwa2/IzcunU6IlKRDjxwQ04ueUIn2I5N+eCnLmnBOWM2zQ6nzz3
3WM2zP3WP8JVT39qunM4wbDKDj+7Lu5RMMdzGmRIN5cMBwOMXsEqPyJMOnehSWrf
7yc9WLIEYpPDlo4OqOyCuA9klfaF9XEawH1Oofnaa2lnuScMmwNbr2o8uFeapwWP
ZKonG7/qVlIWRj1XgfSJIHrpVb0nusdPZdSEoURzdKq56DCqbkgtKz3K3bX+WklY
z5+CPSIk6wkuc2ttswDoZ4mJMA8CI+xB9DQmFGGtgzXy1Qasg1TuGitG0JVHP4T1
FGkkzPVxVUP2e2TDWGD2OfzsV++EZrzbA3u7QPAgLUEQcuEV313er03M2JMLePiW
IhyAk5wwYVx/MsNCJ2NcafXP9U5IHDydNfioXjAi+7Wo7KQL47crB6uML7k62AHQ
+p9sQ5iOCGYJ5TztiRoNrdGWv/UPQrENgxc0bVgT1VuWr3vE/2rcp9HLton+06Ie
X2MnTrCsHYav+RjvJGwOLVVI3h3rNSgfPrswi/CsdLCcFX4ii1K9VB4LnE9yiBd0
mdxcmj7/x3YJYe76+w3Dkh7Hnzh/N312vz6cmSuM81IpWS9IBxgHWYkz4UkdRlPy
FCGOV/ULYUIHOMePiUUT8imdolFhGyDp+dTUup7CYRKhWHcHtfgUmeec1cV7ka1h
XEy7FTq0XwOHF3IwEwwibNAZaZS3PpEy2WdyZzmuXo8grjwheO+qNRPGtozrTG4I
mXy47b7YqnIyQh1HTC8BIyGo7XrVlNDftKxE+tp40w7w4Rd9n69GBUn7Bx6IYsrS
`protect END_PROTECTED
