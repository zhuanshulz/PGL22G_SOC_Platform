`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HdmSPL7wZFOO9aUFp6IS+h2O1DZGBWt4b9/QFu46MMsiHfzYlrqcQOfE5O9QP4uO
WbU9iwbxNFby2u66xKVygZugF4GcRxiw87Dc6up7UEZvwW8Ve1glGa70iYV+k45q
6pTM1Fl8/4nYHjQDPzEkrV9xtiM9BLwR1gYbWjsGHyBae/BnEY+aMnsFOPn6BMTM
TEJ1ySnexHiCBZwDpWnv2END3YoqT0Ty8qEUNGcyVHZIyFYRVAcBcFprQCIM777l
ACeoK0sJ56Z5OWpfJ6DvsXhuAtMUgpyckIcVd3+snPrPKU8u04szpGq7uzPv0+4C
3r9lGJ6USIjWNu7BMUJZ+mKrxp/5M4EswhO/UDbWAhWkR1VfD2mcuNnmxOBN58xX
6gQ7y+FX4Plc6I34nl//6twOFJU0/f1v4KsMedRt8d6jKe0ClkShCkB+pCfpSMx7
gn+Q6TDNX7hEMyjGLT2JcJJ38nAV8UKniid5xQ5U4flXJKMDQ5xWbemhc6pFYoWV
+w8OvaAtCBdJGanRui35Apl+/3PP6GG7CfyBE+ypkDbSDAoGAMrNFp297tNQjANe
//E1lQ9+S9BR1b2LC1+7WZgvzoGqQg9NcWjYTidcDinY56Id5OvJA3ePtoaTqJZ6
6PEMynbwoa4ilyZsmKbzseIFcv4RQAd89/BAqmxaI47cIi3FRtglOBjkWV9DAKiA
wxo3iwSKGDC9GiDLWCizEao8eR0+xk29zw05QX04XVC3ZCA+4oiP3aHl7lgzWj1d
sN7PlEmWP+iJ7ozdkY2ECjNTOGmM5IFRblf+V6UhGJU1DsavOnrtcn0MDP1HVAPE
clagfRHg7ywvOyQxncQ/ZIR+GsgqvBbA4SuFqQB2HSXw9qqaVjOEB7qxJXnaYK2o
GkZdY2BKpd7f2iobWEQZUH0PDlRlOtw+srjQFGodEzC63bnR4QJ8TCafqMeE6Dla
KR/rkGIV7PQfgGwZCs+/A0oiOr/TcLOhNoKQjRxLbm2NIRlOVnnQs37uJaEJUi7z
wxSdT8SjT/ZV+n1ua4Sgz9ry5KrZHi2HA70kjwCMRITdTWmE4lDOI/i6iWzI6o3u
rF/ueqgahtPRsrGgMMJrwx72/6LXXN8KYwf5RBSLZK1daDCzOqhdV6RrxI/XDaWJ
s9UZRWn/sqtvyMRq0t/7jQb/S9uxqJTgKuAhKWVFFc/mXlAqGv8zbSiV2Ygw0bhK
Ph6SQEdmQmpkWMXTLRUftsdAPUFVKv0tESIOX90ckxo3mmPHfSxFdZi3ssa6khIO
i0+kJt9Zy1U7OfPkMxB3IYFuk1eai/+UupXVrmQ4Ff1uLGUW5aQl4bwvNYPVamRb
hsSs0lgRzlGAitk0zTG+VjGa6bC1cSW57pizcU4xClNC9tC6yjpCv5MhkK6WWkgR
9Q5ZtKQxZk/fwGpHHGNg9kx9DWAYuNqG7qTLZyLkFdQ/zQUEk7VKfoX3maCz7Nfm
mqBc/3nvsDl5/IlgAfi6wkoXbVsy1VgA4PKT7vQzs4G8jLFfzuxDpKTXuH2+K4Ax
/GT22A4sDcTPM2Rr3h+++/jmgl03Iy9xLWl7hHSrlInNc2Qm5YJ6Ky5OWFG7RQYW
ox8+keGZDQ7N32MNfEPYd/ADJOFyJ4CILy0cjaYG4jFGr2e1fPD0kCB69OssknRt
u/B53sBuLzLKbX1wt6AKEkX9btPEtghySwLL1jI2kuGo5SxC/l+pMmXifnPn7g9l
nXq202jwbahlkftcnG0bSUZfw4iCj3SbzEd8utkK06x8Nw4hPdwQL7010Iof3znB
bKN2+Y7SqnAMfLnnnEvIBKrfPjhXi2xDjZizPhooCOGCFwRBNB1zT9q++hsr68l/
r7bqUfU7Um97gCNDnDGpycJYOD717YS9hef2SZhuBzphFB9mrD0i/hDbVCSA2K1m
Gt4ZomHbZ26xfBHvL/8OPRfGMsUUcAu44mXSKKvmI7jLwF12hZN87Ap+Plh9U8oQ
hjn2AbWklWdcMWWLX6U7nBOk1Dc6W8Vt1m22GmseKDB3lGg8smKZUIoetU5TEbNN
KCVTlxFoLMMjnGTcgGgk0EJncHZYMiBbFTLFngdz25Fi30563jWB0VJ7KrrxfcUR
HnwFfCUTAJEC3ewDohPHEjOXnK3R6YHBcJXX4ZtIHXjuEXtWXJgz3rSGl+7sdWeW
LAir0BQki3ngiNyPHpaqddkff8EHF85Fs5NJZpbPOA4wl81zo1tkkKxpEgftaJPL
u9x3dmzPMGl+MAD1DXtEX+CxZiChXwfdzm8N66EJ8Hyj1cmCw4z1/Ayoy744RuEN
2UECjA5JLX9HjOOH3Ac+gisfJ+fHLWYQu3niXWEMyosKcdURqJJ2GhTvupLCi6Re
XKXFgaCgW8WWz1rQLPqdlH0RjhGeKFMvz8SAhrL5HKD0R7MyaUY1SEuoIqmw4OkF
AgYXU2qK6n2Yhvy7Kg3bc0WHDOvA6Y73ZriTX2JFslUqf/OGyDHRYq7QOyC+RhJB
JOVRmrL4h7vF5LfChKrXeBa9G27qpCerA3SAUXHhs9GIpwzMfmYkkSFFrTM4BPiS
MMRehvFa8m0SUTo+0cZTF+Kj+GsJh//7uMOdwe8MikINFbgxrgiAlBzuaXYkjUME
PROC+Yp9FiGBymzsz+7Ewa1TkfaUo9RZzDiyC5TbGYQ=
`protect END_PROTECTED
