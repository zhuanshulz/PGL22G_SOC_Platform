`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Uob7c1huV2Dat1J0HnKuJWs8CrGLhrMHZZ2tqP9VUPT0sXLzB9B9HG5ebixS9+AD
DGhz+fz/6ola0Fg9A8X1wi/8q65wmZBlRGYk/Jljejk/D70TM9DMTkb2SmWXigrc
51GNffFwLWm8wHdMy2etFsEBGYP8kyv+aeo6OjO5elhll5pBXZ1TLLm+Gi5s0Hxs
agEbAxlBPCd2aZBPMNgGTlJoXRln/qBDyFQurQAc+AChZFKIb7s+LG9gleqwK8hV
qBm8CjteBgIhPY4SxPNyEjpW+gHIs5oZ/ABnTqMkB5MG0Z3nxhx2jMpQLNbOmd1s
BIvQE73Ejw/r0nmyJ/WGrhsSBWCvBX48XiKIkdRy3p9YLWFJWrl5lEmi3W4zsnWc
cTrhlA2AIbsVyLfmiX5P1vkPj5wg41eDrE5pZwuAgtk04IIIiNqEvS5fB4NxofO8
OYDInukoIIr/Cz5rBD2089wfPyZwipJNba6x7B1YblI6sEeMZdaPjNS1lJuLvtZw
aFXaIASAO2Iwvk/kaRikEhaQjXMXNPxoy27tHemamIXEPVd7OHGFwC2AB4kHvDVy
tlwhh6saQw4G7maFjbyqsNEvxq3Dmg8zVaw9/nyEqnsZxskLYzfYeIvB03nsdUHp
llp23auBsZVnXVYNfas3P8ZAXKkAK/r+NH1cNTW5wtl8T2+kgEuZeZJrWHltGvve
4OzacxGPsZxaHBeEh3h1o/ABGp3mHaZNX+McIdPQqi8VjOVHLKp9JOjmYoBW7tST
rxad8KvuQ+EU5A0HTyyW0fwJ9kaXaBqHkzIWUQxOZP6XWmS4cB4swW0i14UhDJbU
`protect END_PROTECTED
