`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b9wQVqnDuUb9vuOUxdoob4cIFLM8teRvIvVCUHoW1T2VljD6SAFpfLhBbWpNpw29
A/Sl2IQXECGJuYjqO/xDIXh14mZ6jDR+nmaVjp45hlCoUzWofZYGVb6bQoONuPpg
y0BOzeJ7WIWrSuOGH2jNropmVGY21+q+yQjDrbBgTzIB/HKIPD2jxH6BFU18tJbp
1Ib9tIvhEVJWBrcJrxnawxdjjSzNoG4RrcEhDR78uV9uQe7nfAZe+7uOY8mHsE0A
p0/bU2ZS32pZKxmvd44doJ/W2d8hqj4ZR8StwkSlswfa56g0cy4/qIz7ZnfX/DVF
RENfBBTEZAWQPk4uCBYBHFcsT2E8DxR6D2o4/tqTnD161JMjDCfBCLD9wSc7OdB5
IT0uJJDOIgE9WkXd+yIyoyQ31U/kg9sudM/Pb2Z9QqjWxb6rZngHTBdhJ7UGlsN9
lKCF2VKtFKOmMILLI2owkV4xppC2eh2HlYlsAxF43k1ZQGY8HFcv/htkAZTsTQYw
9otDqrd3qWUgoKzrNYwzO0aNqlAfgKIxwvf98qj6FBTEYnH+qtiT+GeL0moqZ4zG
`protect END_PROTECTED
