`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NFzCl84uSB8RKoEsanM+gpGZ6dwA6lG0vso2SsOAE+VgULkFUutSj/L9aqsv82ln
yIyTTKKBpDQJ4Nusoa+75SjVmY9L4SySaYhboBNUe6UXnWr/I9XRA0UFEytM8PU0
FUKF67cJ6GALGmYa/HXmpO/j19NnPWPwNUvU1ZOz8PZ/Kj+SHo6E+WrrJJQCjk5n
p65VQ0eZCJPPTQwZbd5NwkUP6wMct25ivd2wSDGuRCOWURvif+M38qLbgOw19End
PQmmGFi74CA9GZkzxyKHZDw5XVtJNqOJYHLm/hvX/v8J1I/cerFos6FujewpfgRg
/K8uCQ8UdzOroIt2H9BXOzp+RYDO1yRqTqJyFQbOQyVUPMkdszha+nvw3JPjW1el
sBEcVOs60CoZJahwba4PFVcUtvkat+hGnpiac4cKrYFtVoKOTIWtc0a9GKbgpjYL
8aDlO4YhFbqSlKJofUGphTvwuMwONfz2X8BEFp2CkV2VbZC3Mch4LERrGmD5xVYd
PzTW7MYp+/OB4y9rPNUDVjscWhD1GWYhhVOfVcWS1ruvYpyTHuNzv1svOCDYUWum
77opO+XE5skbWqk+w6RUUriZFmtGSbPlABlEhA/Vi/nZF3KAgcBqN3LSRCxfZFHq
cX2aUW993AGmIFAkn/jkireGD6WKP+0mbpbddghuw3HnnbkKa3L5nN58u0+9AkaU
iMRmh+DN+blv86aQKI8k8sbt37sI/OS2M7zbKb48j9Mg9am55ckNuxwOZLgYhDSm
B9HTH78yFr18C9xhKJY0HfrEufupAxggdjykYv1WCwGUaq91Z30R5nNcI/KZaqz7
6g5Q8+n/8XizU+ykC2nKhoW9rMX4bnhT8ht5k8fZIfZfIkrDqEk3OY+sTspb1VjI
L+Af/EAtcyfqWGQuQ4cv9wUNfzkcHBuU6CrUgH6l0HdjWBhnEdA+n84Eei21LCCT
eADfWUBWix3wapwHhq7zlP3Zixn4lO1zj/y/V5Bka0Rp2FhWhYwAW/prs3vcQkes
rZSRtSSR8YEaZyj9M5raseMbhmTKbVSYGSN3iaAI/r7aKebF02zM+bq/092LpHlG
Y+ZwJvev6ctTmC9jYID9Ww==
`protect END_PROTECTED
