`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eZmCA7O8W9/exaNcVs82R89sSXjLs9+P6w0DOpInQbeHOYv8sWWAl/bXSxkHwh6U
nyKsNhHWTNab3Ax53LOd5mG1/6KDbXg3eE/JgYzN5MAxjtokhClTymk6phW38tqR
WT7mOTzC+uQ+Eqfj6ipETFRDz6duXV+Psofl88dn/2G+CejMsrCECsXcj8hOIN17
DwgJETmILVrisgTR2mEc5E5B6ijPXcIQVxplR7jLn/JABHhebzwkRcGqTeuIbJoy
KTBo7kBDHqYBiNAJ+eXrTzjPg+R4BCfIObit2iOueDY=
`protect END_PROTECTED
