`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xRogdnYPLUsecJuqNZ/yrX7H97W4sFszHpEv1tRDvw/kkuEc2d6rmYjZoS5TybIS
FP4T2a5RHExeiUdiTygCgFtygtta1ELm/jsfIlr3VS3C39UmzLw/ztOoTYq8OG8G
IoMan99g1ZWv9STCour5GJ3/3q08KwjT+XkzZ0CUfymQi6SEqnqhpzbsxI+Rtk33
FnFxk4n+r1ZT8aGVstr3mRnES17bOSkw6AvvwhS8Pdrk3nlBhD4iB0sGywEH2TFi
GR+KdHEhggkdk0ibvzs4Dj+MwLpk2kH4j/YHA0/fyDkDhoMPgfJuRfYkNAIMKSbQ
dAIkdJa7mCGSatVbLnN10JcbCj6cDjgyi5md9v9sJU6gmsPniMB9YMOcgRy+23eM
vzV1XDeYPBVasUv9mbStYzgBUtHRG3MDrwoU2Pzl0pQOdxfH+e7AybkPguc9z8Yh
0FbUCazL73RTvzrCu781diIuNDKoAmXwqrYSbF6vc6gBZRl/yaldpM5V3aCBmaUE
T6kMxTPX3Lljbt6+53xpGVi5MrhO1J5DaPa5G03H+D2I8vtud8d+PRtZVqXDDcuZ
TPBs4+9+bULJPmdMLl7DxMsTW9rKziiRR0OA0FMXmNbHBYcqPEStYjeH3EN1miz/
vXTRXrNaZHZ0wDiLjMsCOY8afWYBakpEc8j5Bfm4/BKgsPSF1kW6FxuU7hRb+c4T
sbG1b/PC/HnIEhkqCN9d639+b/IgZjD3R+5YG2TrzUf3kkdbz47MqTRQtcKp32xV
f688vtDvYElhztr8r+Wd9XMw+KzFIi7lNx1U7GDaEcmllJPy5hAVvfe3Qk2a6MT3
PRwsrZxVulDyrR+ghMzeqrjByDx3egIxT0HLdKhi3UX3Z7kUE//qBrhOujEvfpUW
8SIzVxrN9pNkwYKVvKrSZPLNQgC6666EFeBFt4dp7BpBCjEnfEmBpffJ3zfyl4c1
+vV8tk02fTeOWsUxLDzjcFkLNVXSteQGZhdmbV9Ju/e0Eqyfld1IWRuHpIajZVqJ
+js5AxJs1hAMo8hiAWt86bSBF/2wMpE6BiqGtWUXIffX9dMheyCh+N4jIMPPBtMk
Z+T5PZ97uSc0+sV38pzSXs1EdcWmxhSmNwOnW9zDfIyjhfdu2vq4zJa21bSU0a8p
ywiLQpI8NLCMQKB+/VjfzppGfbLT4ZiDMblOwJQ53JEIQiStfETTSZHP6LLLTQVw
1q2taVHzg9gh0OkRcT07KLyJwrbA79vr2FvXCDXLdodhzhRgCd55p0CHx7O+Yq8W
W2AJS0fsCgb9OZMgH1ReKtWO6gU7kK94pk26YwGsyNJhGkufpT0TUfyb/R54Ajze
tAPD7SHzwwABP6GtdBjqwzHLcf3MVSGGoMFAnogk7xhpVspKHd4VprEPbNhm4Y7C
a+qG9awczb/SALaFV9fKX/nA3Kzkqx74e3jSFlw8/Oo8tkBCjK0ChgDo+Y7g0MFq
Y1oW+ztcvU+ei8SRBQ6l35wvpO9p1ZYxGDLLUJ6QWZxw7UBJxGXIZHl2vMevagMa
xcf6wSdKY296ZT6NPfgRHMESnPWBxlg0Q2QpyHqju+eSzdw83r3Ujmi6yn8LSE5G
kD5HbWiEj5b02lf+IeGw6x/XCyQRV/Bk00dJtu0plI4QpSv47G02ZF5yV/t/wheP
s2dTpgVhsrZBb8ZHxfGsB3yEQlMtW7JrpDG8lG21LzkIij3mggd/lt7zVSglu+kf
M49Uyjm2uUabgbqrWKtr+9qnFsQmO+uliEzTfP1EAMjyAwiS5ushvQ+5NLtgOOdN
18Z0vWwRfBROowdDH1NQnIaF2xzJB+9nlwVPNpuYXp8TJBLv7NkCSQ4pV6cSeRZ7
4uPx9SqQ9FVosarj4DY+f86Gp3bd1d/k+u1jt/Z2S/IdhmK/Buc/xUpGBJbDr0xN
JPbsAAE9MMByxT79MXiXNXUg4AlkVeVqNBlrmB86wnjX1fQ9cWnOsMIwy1T971Cq
ijIA8ARQPMAw6ZCNLpSZEKU0W5u2EEs+oxi9gB5H3XkwtFnwSY5TXftMvyT1ozyp
cjSwTcQacJodBt1GclybXmVDljAZeXdl1tAJtoHMv4AdlwnQP4JyNcsuOiTENoF1
vWH1PUC5g1cOJM8DkvT1IJv7Rfz8uDHbtzZ088bX6CqPW1uOdw5DMCEPns2x6PhX
SNdsmPKsuASywu0qobW3pAiwPngjGb2nACD1jc1v7RbDE/js6THX8XI0fww0vJgO
EAPntf7RTVI60G1W7ezjPmGHiIbCkXASQasdwnKnoR2gtk056tAXcKUj8ses9cox
I5wpxXlr87C92OSxrX0mQ5Bmv02YNcPwOBZrmTDuwX1qDvjplsejCIcMc6gnZh0F
ZU+85BR+qPd1sy44TCJr9FlaftQnQlAkCMwRERktuo2AlqnLGxvrUTcRkJbpjIyC
6Fec/mfL1RZGJpyhCee5hlxuRBNmDOp46juJrzarf+QqtvKRXIcUYxkVQ6XqSycm
`protect END_PROTECTED
