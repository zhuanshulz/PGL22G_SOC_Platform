`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qnUrR1COsuphf6hb5kQ7QP5lIZ3Vg0fMDoo5cDIwZn4z/gTEM6lx4uUoosTxcZoU
8y/jRXgqvirtMbV+Njwkca95eNxNDJDVpZ/TN1tXpE/TSN89qFd76N9X1+UxFJBK
s5kPatPeylCJFxjkPdZGm6XnIRe2lbqBSVRg/1yGCW5yPNym1rgn13Vq8bo+9QnA
c833loGj+09ydGiGBZUJVhGY3XJeB4KY3poeMmhdr82EfUp5vslMSujN+KUyHnNE
QcNCZeQTNBMV1pUC3TZjCPhDDwObC/Vf4kV4SpCZAokiJZd8y2aSszmK5bP59+Ai
M2vlqM4EMyWpFw9cjaUx5DKPHo3jtN4dSJxaNkR9BSuZlvdBwysP5usm4v1XRfPs
jeDHoKJV9JZ3DB/Ft4oXX/EBv6vHmLAVjjbHF1Ssxmc5ZvpZaVzqrs4572Vfk6cs
pEwPatZYbH+mAonAfKzfIfPDJcjrDI/IYpr4/XeslIMMGDr4NT/KwZijfLXHFjJw
siWqTx7z4aVvk6s1WQayuAsoMnxg3h8s3eaPu/ba53VhnRDI2Nin8pKlshZaUOrY
/72PkA+8UGZjERw4PvOm9VI9f4bs9coxVT9ghFB4FvbwI25GxXZU96Iq1wwDnE8A
LAG0/BaXnKUkszopHm9Sz+HpOG0U9dd6yjfB7O8vav8nbXQJ6qJS2kkt6s3vDj+T
Cl0VzoY7GSjv77FzJ2gAYSLowgnZNjf37IW2ZB7/Hj7ft0rPiQZTWAK2wAC+OoLP
QU8bfvKRWiffQ5Uq/xmZsw==
`protect END_PROTECTED
