`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pFJnOo3KxyT82e9p2cM88IQixqb/3uTtEjPqYcI07RTuyqmBTFufqr6bsJP3pWuV
kimGj68J1a4mJFEY//LOULGB39DNm3io+8Pez1oez4nzuZP+ajnJXolkOcmkLU64
INdKan/NY0ID/qmz4fudhWl07fJFl7Dcb2oymmtWNUqLtTl9lxAQ8a0augzc9Bqf
daORErBwfTSHbXE75GDVTrefrKz+2Z86Ou7WMZnxuavBoJ4TVGzRSMDuoz8CrDy1
xEDSdys6Dv945QaCX15fyy20a788IiQDmVs3t6fT56VSfBZVye9hckqy/GZKvSQ3
Ng2k2q7iu+Rdolv5Q6cKSl9jRz/IDbICvXB0fchZ8Ism2GocBbc9lzzGm7KiulXj
M46mj8HXJGPCuZo9sGx8teIK/GFx37KthYzxWh9kERovq3BJ6gWjIEcBfl35MIKO
`protect END_PROTECTED
