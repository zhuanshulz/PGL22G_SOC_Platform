`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MIsSmCWlR5XC+kjR+DVh9ENrO6CZo7dPzIRNeKQdLoZFqCKTH9waH+ZLEkwUl/5D
lTSTm/SxOk1pAmu/VCU1v/AI1mKnJPtt/EFTOJfmOv6NbG5OYwL8P29j4mpb3IGi
jLodbpDWAt6cmqeEfCGYonpE7WgQwkTH0AdmOqg+fNioItJ2LjtIPbSl0vPfHk2d
r0nzaTdh51eiVQLlf78mObTzo7pUrSz2xLs9eknB5YEjhtqyLoSiVW0bQlsAZ6+D
wf5x0d094q2nXKPjYbTzIf7rQUaLxUsMJqCZ0sTKWPUE+b6OknYbyRWHtuIFwMTj
qZ8zxTghFYdCG4RBAS25STdSD37gsbCQe4y2LfI8EmZn98M4s8IAEblN1vf+dgkK
mZQLD15V+Bhqv2OqjKm1v3yTdws04WhrGuLD+es12/Z+GlOYI0AKSYHSmoEvDWDR
hsY/hi5OGabngSZrh5rxXCzTBnjbN6f1V9rm22y5JqBL6doa4eQaGcjbo0RZHjSk
rz2kIYOQtWKhE7V8ipHKc79nxt6UMtTGbXmMxwbq+LrSKx/s3et/P4QV/ujh6Uf+
z1mTWGw+xaqJvqALiGghPw==
`protect END_PROTECTED
