`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bSBre/t2kUz9JMydZWOzeuvTUZr+00kpSQJx50suvwHqikzMWxFXyAwDngdicWc+
xJoTCuT9gqozN1y+alXSeCAFQzhst0ouMorVUN1ZxE+nHcSDQfGnGwj43JHNQe+p
bn2I2m35fIWXYMyty1MQs+Xx8HXXW97lXl+4Vr4V6pImkuINpIoNyvqzb+Ug9xrk
peYk9O6mAjJPpiZK1W7UBI9Y0FgMB3j6viycBtY7yo8H6vi1rkA9pwIH9nU/J52i
7oStApFa+JtcIotwKNTn9WvyZP4kKgY4xWbvpyj5Pd45tXDldjO9X4VDemXl5eEK
DHNP6rakwyB/NahIJuYs7sYOs6bL4wmYCG8Lsl9vQ/2M2UPv3Uz/4NQ+oQJuT1XO
JqUzYz77eanqhWGNo374k6rZIAYmBRSv63kSYE3idcjcFfaM75HFSnh/NI+NM5Td
KY0VC/c6Tqx55X3jbd2R/MD3wt7Q5ujm6Jt1q56KoXRYrueX8dGmqMZ8w7m782iG
4Y7VaPgao8rDaD8epDFBqAiuUFLNEm2NrCQ2tDRSE3z2gpgi8+Y2nxmTgj3vc2AB
qD1AwLcAspU/LcHfamfEwJmWlnmw0gEaxaodC1Mw8BWK4xxY+VOQU/Zd4Ww3VeRr
aaEv1Lsl6+H3PB60n9oX8dHnHN3n5nGKevqWpGE7OEqqZNLlGiaqIc8Lpi26+EhW
dTBoMW9Nrwct0vt+tOLJI968wEdqY/HbjoUFVzHQicFbBG+vPJPevFAfl5RgmIig
9bwM7E9tDTuj7S3uWBskJrQlOIGUZzh++/eCEbpSR/tdx5b3g/76e+dpyhac1y7I
pR1falOv8DW+ywAqjCGRNBbr2C3uPIoakq0nx2Gy6GXeN0QP3ZIdlWgUlQSUESgH
B8p/8q/YhwtRIGCIMMWEUu4tYUR4HDKwTb7JU5Ek0KM9Xv3ZMNkkYA9eP5LTk3qw
p8Ahx2Bb99FZUFHEtHoGSX96LJnX0R0Wf6uJ2mkyYAJEVA9Na6Q/2SM4oMSvaTkb
1sgHbI/GKKpbkyyj/lniawh05BQOCZqbizZw34m3uhwLIa9+MVlSQL7QgN5iylo8
P8JVHYAMNFsdLfEVbC7GJwyQgQT7+OhjBQrBpz36LydV/cW1Ym4eo3inGpp/wfU+
eCTNVF+w1U795IvoUeAz0GaT3xJKMVt7p5xfsD3qI/mhp8ByBzei5GmUZvK9i7XO
Uy7J+YwM/78Mbyc/3SzzwDW+4vW0A+s3dxxJj9pos+t4Fl/JeyPXl+IC4n+w1p1q
PnFyx16B1r1zIr5N5mQGc0UIFC7qS4WY0xk5k99NjHQLI0sY6bMHXPc7w2QEFSf3
4ZXKuNsBRIpHYkXYNmCjEw==
`protect END_PROTECTED
