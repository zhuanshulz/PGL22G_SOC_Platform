`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IriQ/jD992fKa9nU73uOGm0h/V2nOLSrbLajSGf+1+IPrhWZh/EnlzzhQ6qNyWm+
C64GwRCMCrPSM5o6q55nTgb9j09r0k1pLepNyAdoyzUWdlZrEOFf/LaKsi6hUhSK
ImwoYIQdFtEJCwwyTuE0H0sXCKBHCPgvMmZho3gl38UvWfIWuC7PO+geGG7SSjAC
6axq43VB7Wo5VihbRJBeVn7fC42rojdL3RRHzKqE27S+b5jZFS0e3+JNf2Wbkk0X
lXit6kgfPW+39tdpojJRA9AUn+PZzqAhOngmqX9h4rBsYoLx58oy8y+gSY/a0gaG
gtrlKAVZry+HK1c6KJDjJOwdgzOg4+rAf/fD2y4El1KRs+R2eiLDe7BagpOYvWvD
DD+x48d44WRubdz4SBGj8U5YH/Vf96io1p32sbH4HXxZfuGFGn+WogbwXRk4aEpe
N5jbMbH32y4Dzv33A3pmg8qC6RROb+2a75NZRJ1Cfp5ILuQWrRsgHznhcsLult+X
YCdLU3xHkKJPMhcI7h3r/FH0HVZXu6DP1YRYW2du1cBE0SqbRAoeMrfCQedbTaqj
1yCgl+yg8poxJk72R/2Gqwb8k54nTi+9jh+DeSCYqv56qOxfhw+/EsqFELL8S+Cv
fiWCytW3CX06yG6k/0ZqhxV89n4JcHMRr9r6XffHN4C/VEH+xltsoIEc8cHTTS4v
Iy+NlOPLapgyjYhwXY8qOwBxCq2fp8+pbo88O1tWYF4L39BXn0a2IkXd3APT3e20
Ugmr6HpIkw1iIdstdJtpoWHhvYhHyjU4SH5f76rw3jx59p92+GKiRCYwgRTr7ibb
7KF1UnnpHjpP4SSY8sFY+nJgl+brccMacuE+mQb8uKfV55xizrv/1z4L8HgF6IXm
L2+akEytO84jzm1BgZgaOA==
`protect END_PROTECTED
