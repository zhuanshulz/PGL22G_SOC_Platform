`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j1sXqPfcMg6JBRHuCHYBBmsrVPnPj5LzXokIccAYzJJeVJlliYNq9sTIVANN4ITt
zbyLpNEpBa4wMDfwFYWwNRA6z0OReotxujCdzhQ1UKD0Uh5VSBjv6neQRbNfNGb1
DY6NmCg2GcD3qe/dgJH516l3G0aooanD/aEjGlOP2+TpCTRJUc475ECU2spdop1i
1/OubW3Xdz6Xpg91Smf3FEKc4YDlBe7shzyA3LW0GZuRR83FFYYBRyDLySPlQMrG
9dPjRcEDVkCEURVCmKsfpjVMDHioj2rlMLORP9HFVcaNtaWBhqJ3l/z2pKAkOD1A
fXPAy5LK0z7bjjnt+pzNJYYW2EGJ0TvtM+JqoI4TzwIDO84xje3tBqp9ArrPFSVn
09jAkgFeQDV7mt0bEpc+4DdPj/Kz7mVssOd7qgglr9Vf1ajBEh9/pJafxF2oEvPJ
p77UvKYA5i2Z5bPucQOJO8vSguSNJw/4JdotE65Dy1tRxOnTM892uSLVZA5s2eX9
eaV+0NhQEYt6/jMcENmM8q3H1Hl4Vp1kwpbNyix6b6dZRf/gWPIDVNErGq4zkHce
klVzlXNzEnqvoDeuAl1qcntfMIFRw4y42aJGxIRaXQ8g3Nq9YbeIuyBbfDQhtOSE
VZOgzGybEZnt7+xIefuXUhIjQHru1Ug//QjvR7fRw3YzQryOVvPwiv99vGfiVjhy
y/sHrcv8iC3SKvQwyxluXWvy05xc+bi2AJ1ZYJ45auquURdzI5iQYulxNh9hXw4l
FDSwNdY7eW05Xst3eWa+2I/J2Q2VCsXoOJoX3RfJrQQ73UX6liMMH8u7rUIcuBwc
S/WslNkXg88i1hNidxpZcDhQ2THHq7ak60aoNDlt0K54/S687SD73XISohn3/5ll
wzamHHGimETkt4xE4oVoARydZMPpQMXS0kZ9kwBScxVl5dNrXxqVGWRr2x0XN1mb
kQa83L0cge+gOXWjRAhvFJaVosdb2vdBS/RMd3LmmTrN9NAZt1HF1rDn7ZdjlBX9
5Njh5p8Z8Gn+CpHTc8qElcjcD8OAsnlEtoTbNY7EWpMp5iZOz3G3iYhZHbrE5+2j
n4hA9ARTroxBnnIMKK+7ZCbqTjNv9MIv05l3SDYM4122z6LugLXThqFfAF/HJcLM
uiuugWjjPNQZOGl7eFk9iq7KhKGAjSpV7EPOyKUt0bav+c749ICgiqw7bEAeN1ll
hKzlDKuA1QU5v2OnxVKd5QXkYnM17GDIRZWspkY7mbfzeP/TOWvALcHX7VBsS6ix
Wiy/1bD/ZNYwi13KaFz/1ytwPjs9pGYiqdV6yrUF6XlRKzuLPricxDP2g/nFRfKK
1GsZBPKSETYHlLX/OBbEsRHJEuvKt2xrdM89CvVeM/+w/WvlfuRnjct8A1HmpgzT
Qq1z6KZLotB4D8JpkMFpgA+/9BoNe/TFnbk76og5+wqlJPyxP4yI8fOTU9WmhZG1
EpO2Unr+m2UlIvTp9plhnnToo2SUGuGrjqdhXSzJvh94ilAfAYyJC2IghLH9gJ0D
RDYlkyAz2B3bjZWe1i33dLV0U04D5q64yxfmUlJj7YZ7EDRckSc82l17ZAKrhRtJ
FEnY7w76yjEAi1aSmzhnBgYxtcgpquWehZkp5xqsUoI0huel53k3hT9Z91nrExiP
OOn2JRsmdZJpk7U3As4REXh4MwpxWyW4arhg14UPsnvgUIlDE2RNaPcUctD1QXqU
CqFg30exXRkmjyO0NB2EkCVvdu5UsxzYoXKOJzxVzGpr/EnlVHzgVL0SZ/7nvA26
Ga5cR/l47hIAlaf5m2yA3W8qK9xxr2YKqC5qSSwG3+QL3Y9JBgP+6aGnS1zvn++i
f604EwBoleLmR79NpQbfFCwxHyBZfkUyivwgPvJ4dF9+ojkVRBvyjYDN88+CglBZ
s5oJBRcMBG5n0sNb9Okp4rwfBaanJjg+EQVzorpYhduf4I6kXaBU9x3143RijLUd
p1vq57nObtdLejbnpHGtvYRQnuKn2w+QdZhCou22fn/LrpwoGS8WA1uQ4yxp2kAw
weG3W1S+Ta7MyVXCHxhKJcPVeXwG982dSG2g/AiSPoHlA3zxLrDHadkHQ5DWqecY
eWgjqE/M4uEFuTmBGx+VNmjRYZgwtBfcxLlu+u5hGDbVZyrc+GBML8sEUUGynKkS
jMEs/C6qVuODl9/CvSFMScR0HOOuMQBZGe8cajH50PgDOao/GlPSiQm/nyNBl3ux
jecyjcIQohRwG6Tv4/wIGjdJMD+TRpH47zYIMLdHYLZlvnVf84WSqc9FxWPhXq7Q
HRY5u8UCni2iPNz1QuV0yJjfxXUT0+6ocOJ86Hb1dR8wO6LYsrb2ndq1VhRJXryv
S8/MTqggyUKupWgpdM7XCgY48lVE7nbnFnNGpp4FR8qzI9mi9zZCxPlkGf+/Z3Rq
zTRhDPquA6A4i3ZBjLCFgLAbT8dxgQP20l2TNwcwIhNp6CaQMXIJbPouOpNYq1kN
JZI3C/vvqFz2fGLEXPkinnO2vubMkMkU6knG3kvoBhtTC2w168VspCQ2bV5B3VvC
ECyhpVM97zeRJPjAZ1U56t9mBzoPuDdJ4HrZN5Gz9RlmNBCMF2GMe/pOR0IuD92H
zijwsxTctAtJJMAU4p2mNjME3pfG7Dd/lUK1jVBaFJHmLMPc5QYgDOTQkpPnCJ4i
cFpBkK0Gb955HIOs4XVmgifbsH4eABlBfKMUx4BqIZplQyuXB+UfP02Qnll7CPwe
UdsHAz+wDDkfO39dK61kW345JY0gC/+0OS1GoQTS1g/QOKGaW3gpXxVeWNqItNJG
i4Ls1pJcfu7EYX69QvCPBeqW8P1T8NxV6yjqbOWyrOZHvLgr4x39OUrRQ8Xj3mhm
NjKmMpA0XPMOoPI5BDZJ1X1Tn0Bty9uiZAHOmziaSXwd1/IxFeLMRgU0raxMUvQD
yrrhJtxlcjQcYbKc5KrCT8hNspnRnRuWlyvNJDuuIu8SkjUX5cVFK95MorSk9nPr
7tNTO9IjWtA+CKMJXB/LKxf6nFZuX+CU8NXr209DXN+R9LNmczqcoOXxBkqvizyP
yUiBjT9ireY9UzZsjBJdieKHWpnmNX5GYI2Vt5A9DmGpzsMGozUCCy7lRcE+7B1e
qEPoMz3WkGLlBL9GydqHBZmR7V93En+7VQbpi7jSaW7h+9+zNQ3gz4+IwKeUwjaD
oKsIwYvupThsmGTlTFtr3HOfrUAx3j8alDpjZBlsC+oelWmzLljhdimtBLIlBMfT
ndhchJyPZvYajSW/j1JP/KjC2o7LiZVOH+haKfLZbqQAtBlEyO5HhUh+hKNh5gaK
hhGoQJjBDur/wBsOV2Yqyry8VTAd5R0n8NiqIwvSZWL6KWaY54D5nZDgQVdP6vAz
QOsgBVraXizkRr/tYTemKtbin6U8n6rymq8TfGgnP3a8xRsVNKtekRjxj1ShS/sv
kmMof1nY6cVTr+CIwDgvf+HmrBl29YU2SROkd3llgwDWcwzBv6DZTnB78hW/12KP
kbiKiXZBDlKlGDEjq0KEON3mPXGxq7H6d1xvjM3mdOfI27gLQ43jlyt0a/wEtoN0
ncMGdaFBQpelDkO5pET3E3EQ67dAQw4XJvoH3k0LIG9xsReR1uJ9dh70PuWoxmm5
nNGU8Mg5sGeSBr0GZWD6gYpmq1/F7QowBGXMx8O3bno/bEgL7zB8VKgtbTojNM7b
/DnbrqxH5nkMGXUiHnvj6VX7VHUUzAX5IIBX4SCnvVnKZAkeOUt4vgKakCB/QU1G
QXL/ub3bWBrCfes+m0P3QS2yr+DR/5+KPaCPtD9SocJ3G6vJ2q8YvWb52DjZ6pKt
dwFCTH4mEkYmuAtEjNzxfAxOzZ1A1BK3XmRs/dvDjDPbaXrEQsTCvY32+jJmWwql
bv1UbPaXxhBBMuCLgfGFdnE4kU8/NOUmrqXzOfiVI9ug4kqJ8SLWkmv/9PlQ5pMp
jtuP3diEKJgNPUWK3vKSy9ofXrasiwPPpaDBhzHxiT7r+2RMGYQr3Xss1lau18Sb
EKPgKpewGZyYvrmBKk+zm910aWoFpbQC0KWZbJQGcq92LYxpevTe5W7XGx/EWVqC
B13Qs0grpKtZUo+D9F7GElyNHQ8oBjvO9BMque9jujf2qnOB7NCweiDI+mPbk+nA
uuautzP48s9MIBYuHcfXR9Z5I2e+XE1wqzf0m/uB79ND6aAja3Dv7T4hV3B7XfrF
jN6PvgMLuMtrUrpy3WwqNUuYTBNsV0DlylIZjwo2VrqtKf2hliCVZbNRXcvQI0ZH
P5A/h6JXqMeRIlzd4ojlZ73wASABt+sf3l1phZ76gddNYdbAfVOLU06BjuOVSFzj
GE+/9ZGNbYlAa0axPLLAl+qfdblndyDrupADDTg5tXzKObfL9XMeMWEfLJLYxLso
WSMmdz+3qJbHefVKK2T8B0TygTrgCgH77htZ6vL7bG1sufEHpdGvHI6KdTu2wtRi
mOEeYhCkxJJrenz8do7LW2uIg4C51JjPYWklOBtF1pPVay6EzdtyFwmGml8YWiEV
y+GRSnKWyofDt6aRTxz1U3lqi3kPrMiYgVblURgQ0Nre8YSDspoQqm6aWKkBbQmg
xk/J9TdMuq6f7yhYbAYg10Z3PVYN6DIOMslHHWZx51iAbCby1oAljBy8PxdQeOZ2
SD1wMNpAaSrcTkvxIQ+8AJVnfzNDeDsEt3KDpaZ/pnhMeoxjzX+RunheCoJBr+0X
COXfVCfzzRpM9aPWIfefnUsjRm0AEtuml+v1DQ1h8SStUSOg9cTjHkRRYeEmUxod
KDJ5r3qSj7bYj75bzlBq2dohwsKrt8vbMYl/xQta4ZZnEv2d6oIMwJ4ecwMdgTKU
hjFjiuNJrF9RkmdVRXbiz0QG7AJcjReEs9UxKRpR2/4pjMVSeFM79boIKKD1+ty1
4DSnS37D1ekPs21ftd1DGoTIq1pLt0nEa0jR/7NoI9eXBxCb7K3jsovTL/YFcX8b
yq35Oerc4wG5vsCDvooOFgDEvDwIZGsBxOh3ZCWBZTRBtRa5fzi+3wMzrBPSl/Px
kXmcq5CZJOoXWg9HKa7q0vfqMb4/+RVZ7XD87n+ZHB+gmDraUSRJqBwV6E31gxmU
1yQdAsdola8+HkQRey1b4b1FcQL6vbxj/UK4HKjKUwsYgPdGjayzEItcaXkvnyQm
bCuUo4X5FN5KwQ26I5HFK+oxtYDcjpCl9B9nAZvZBpFga8I8L3cw3dgQf0fyJnjy
ljAXC1ttJbcG5Mu2Ox6dMATY+HMT+6uTVsvfcmfCTv6VvEzSc2EVwSK+slsvvvqS
VukZACmcN6VmkvzyWZu105nJKRqDoVkZ1SaVKgvfhglyWNes+ognNMEkiTJ1j9fQ
3IBqO6EH8g+LV/MMNMZ/jRb49Wpojw5PfHsscrPajHi6CA0TlM9EQsfAmP7xo5Hf
wQAR3pXfgctt7RDVGnrQO8gSEqc6txyrXiBymP3FG3wLpYiqvKz3F1dU06Tnj2h1
55ZeGjaNHF5k5bVFSPucJqEAwLiVjpHClrTReJcgfwrdMchnzkWFJU0VHRxjNS+e
jIp3xfJSBvUa789ffBslq45hJsXYG5mdl1jIgd/iStKwehntuY2YTh/Zsmnqike4
C6he1n/56XwIKz51/hM09q7Rq3WwXb8rb4hO4WmQqsBHr94de2DQof2fkN9PF9KC
/+XhiMTIHbDbOHB69jKQeXAN2juzjoDuqWz/bKBsfgCmxctfGtXVcvMpxuOog6tL
LhmsMm9yx2KtKteSFodprhgJ1ah2dB5J/bbh5CjdnxzYAWuWQ3dRRON46+voQDqT
+e2EHi601IlyFlVhE+gIR2IU0HCfbTQxCJS4Tz0cZy8+/WGC7WiVe2seaZHrx/ne
BGlyBQv6ajKHZUCdFWvliLShQ9ANqsbl/TdYZvRgSdQkXQjyJwCmHYDAlsNQZIp5
DLS2A8fiVmOjmRLOZaaTaot7v6nLBGMsC31GdnvehrTAyCDlFGDK+A76zcCKcClR
4ashIBS2/CFVR88PKDJL5UNqA2F1u9OeqKXfKVRhNeBAqNl7ynMaEto4oVr8lA49
MZj6qezo2JyPshXQ+XXlOz0BBhh9w0VNeDB18pyf1rYXQsDGbHpZD6E6B2F+A1f7
tDB5nPr8m1jOzqGhP+niEEt7TUjKdk7J2X6095u9vDtox2aXNCw3pRexaEA3cZTf
g+IVVhuJjAKVIUyQIT26YnTW8A5cNmOG6s9zVPHO8VYtZJAN+EpNZy4mi2VCy/H4
XmGzSrJyNz5GES/nVjFDxSVkwK2duIsOBXchwSoF1Qp9JqIlsX1XKWPNoirJOS8s
lkQ6Vb1sJWktRaG8djF/nHGEqm0xTKZovTxuWEz7clkwCQgDTRjXNqbpr4mVA83T
e7aoHY058fiAkeTNnGfLahL3UQJkJExpY8jRIQN1WxIWAkwfqOKbwcn6iW02HWU2
+2w/ppq66mzJesESvVqYa1IxJG4cwWu8M5Fkxsj3xD7ZJ2kJM2HMmS7IyuQMLOTM
JaONthQrNYYuReqBvmoj9gwgCXmryE6JvJZsvrsaCgDsbQ8711gBcC+dLqswMa2t
5DE0hbc4RsijZ8jw+P4k8Hy5iVdaeiCEouqkx0EBb32Law76CdjvjenyhTLGZX01
pClvbgvTqkVYEw4B80nPS2jgeJErL+FGFDD/+e03dnwEPoRoNW0Ysv97cwG+gDe9
zCviIrIgFUzTyVNPQLeliQt/PyqPas+r0QMoZXg6v3NblmU64ELiUd6GATy6ay8h
zHhQ/8fTCzWwoABiSnvTpuCHJpkgfUFj5/LqlWu7BLNHUpA2pTrdKgft31ess9X8
ktiGellmA13nv+bO+KiRcThHrrbc4KkytsbRMvBjZjFw6u5wRxe0zp6Wecvu3XFV
jjvHH3B5ymmnO+snXHgQzNf/GVyTwhq1uZ3PHOJvDQcvnwZ2G+MTzv9YaiQc9krE
ttC3KTAQBh2BGXxgKQDzdhxNkTwTwSy1c7DI1dUzT5LKzb/89mwrDsoy5zo413iE
MOS/ZAMJMsvuu8l4fAKDP8gbyWBf7YxueOsp2JdpckQbVJ0fimb0oXKMwK7Bw1zg
rTYyClKDXNIVmSbbi22YVQfJWMP1sEFbN/yX0JbZL0PmnUwl8Kzm2SVQW0c8Xbzi
Tu3Qi0etm3HU1BZg8V6CvvO+WuZeq/HPnkNCxTH+I5bUvG+QU2o5fnVXFSW7sOtm
lxnJxtaVYxPx+bVeNCr04RfnmIO+b6RpikvcFwVWIxz44qdJiCf6foJ5hCKB1KWD
eXKDtCN/hI8n1hvXcmOgkYWSGnX0TbDGkvQ5zMS+LRHj4Dv07bk3BZntOMcbuaZR
f9F/nhnBPUdvbG70YOwAUjLoRBEj3qJT3t+X09jB760syUVo0BttGkFMKNCcBeFR
4FGb1APCBMo77ZDvcV5I0sIJL4RtB5d5ZxaMZhmJNwIy4NBmVw5YkoU731+OOjHZ
RFrxDJXxlqjjZyzQENcfyaoVTGwh0aj6l8/O7hRAMDvZF5KXvqqF+IyRxixA+vUw
tluJeDB7MVuLAsWTJ7mO62+J6Zxf3L/6O7cITuLOUQu+9Khtfc+K1DBXSfcUujGr
DSh4pEIQY/OykTx+dJTG7XAK6QNCoVrdsGZgRKoa7/l1yZzChltml92gBpMO9X+0
MNQgcJa+i54YyIuofJuZdPfzRvr661ZRa9CR3U3c9Xh/bqw5LXH/TfT3DstyOaMx
oZ2hyRBXY8zkQp8p7pE6R5uGqEWvOtXvsTCFrcVwbCNFjWktQOpiuPnh3i1Gw+Ua
xSwzq6TYKvfS8p1ChzMxFECe01j/esqkRJNR+M3pVVzQm5w7rnen7FQG0fAd2pst
NzWWWODOJn1oVrRoBvbqVROpsZUMmKCNQ6fjzrOvfIyT9iOkuwqWsNZ9HfELOxX6
TwMxnLpVITnvuwehfHg1pJT4iYUgNpNPBHE7mV79oUuOttA2mpSFTIbelNNeKtqv
TsTuCFwiNtr8uA8HBQjhQFrSdRvA4fTI8F/LUW3L4zWnNIJZfRAYH5FpJhzxiKE5
sUXU+s2ty8cQsHacXA72xNdUbyTzM9awpL4zxvNOmxP+AS0bydoVqUJsuS4pqO5y
WIuv/jc5CVj9Ks/prekvERHvRFVdEi2mtliS+4OaAwmxgH4G0TAqwMakuOBS/M4X
Ff3HQrXQ2fV3h5/kMF5q14VpPgIPp0dFjy6vHtuatSuxkkKVIPVjazpx5M9ueliu
qKM0846ybCtngf3b36p1cnrRwxNb5C76gjfBbx3JUw7UWr7QdCVckr7fjG/wf3En
Uccrlk2rZmKgBUVc9eP9N0vdaOD28kxbBCvd8l1wiAWrXJaG5NO7vIJL602uHq6y
2PoSnO+N4b10xHlbnIe+21EwuN8vmI9cRzp51jKdi4jV0M6AEF9merXAz1Rir9rU
ynTO78lRNTJuovauy65ig6Kk2RxtNUD/7RVqeSqqPdqeQHd9Ws/T8UnRKT2qzi5S
Bn1dSnQPIlpJG+mJqJFgWr+qDgrwO2fe2MmNuI8L391OWFzLhqC/KDYdT5ldOzql
msIhUrhFJqlZ/JaC27eJ/ClqqVWk0MblvZtmQljUM+9RId6WOpBjG5w8/34/aDvx
Tgh1WGy5D3n3RY1Ix8j4hEpK1Se6K9uBmQ/eCII1lrErgSz0SVy2Tk9kPmmK/Lod
ys/ly3KbOFRKg90oL1hJo+1CvUEprBKwuHvn2VdsCEvHWCU77cDHBDakxVAnze2V
TmWdHtg26AhzM5b1RKyrhqO25VoPKjDUHZ+/ta6e/0sK7pM2dnMv+uMX7ngM0iTH
R5bVEMAJH6OfEJ1XeoigUiyAhPdyiW3ouhq6DWrYcJ1gDbkiy8djf+ASfuqvoeuQ
4MNNI4dJEPXfSTJI/NyGip1xYRDd7DP0FD+p3m4RquYfwvtjp2VD3Cj7uVQsnPgA
uwbv0nMwVfs1QhM8U5yZda+IIeZYs7EDUvNTJBDf5zgOO98uCCO/ms6aItbH9kcj
Xpff+BI2TgszRPxX3yieEwHv1OJf5n5jBk7aaQY6wrNqTcUSeaXxsNSSNU6gwgGs
9yevm5CpFS1G2RDYuMFj6GigVwah8yki7ewm3tUlGWOaME4r5cUOTwiac5AZa0nV
SEthJXAXnPHJKu1mmC/bMoWgl0uBNe62ZoQBypfvORJz2ma33F1pGue28s6gWC9k
77pkQKi0Zh1H3H9tOuPRMfy/6Ueu8yTaYps5/8x2AGdjDBUYBMCT1QYLHi8sE/i3
ASZoc5EBGGUED5JhcdTKrkL8E8GhhfYpYrNLp3bvY8fcb5a3Kwr9c0U9KplOVJxW
wMAuASu1hhc4m2vkyxYpUNujm/cpejoVZBbdtawrbTufElFkpUxPdIK2HdjoJRoJ
JJ4l7D8ISWsBxvRwZiKkKDm+c2VGKnjcciB0sCf2810nRK3knKovfaQb0bT/sp9V
gJFJw8wTAEB0J59TXFHdBm/7FEwruM8NwRAsVDleQSO2/q2LQGOMfB8x12xSycgJ
QrSPo+8a5lh6dRI2zWc+KoCxWZhiK7QARWKTxpXWylXdKBCluL9vt9uPxgFnGbFx
4HFBjQdwx+f0prf+ezJrv7YhUB+FdIYp5h6mTBsg1+M4azPd9ouKuUJz6r5xuLLK
Cp+EmWJBIHuxigFVQGE7BKlYf3pSc6VeqHNLeOgauzTtPxU1feSSE7/bR7fJuO50
xTRzyw/YQueaHix+L4u38kLeLDW/5xPxeuVfnAETRTZl955ZsswEHHKM4zmqyrkc
5Yuxm4CnykTchdtthc+9c0G66/oBObMc/HlcJ7Oi7UETmh8efGFOgUZ3zAoFbLaq
ktNQFYUZT6M/loxK0YErq5qAW/8veT3snDba0RUp8aVj5Wo9ycCC/jhONbyIJxYr
i5kOwWX+ANwkpJg25aocuDDVW0Ktbx8b2Im7hGrbtWF+7ih9iRsES5Q/THBBrpNV
V0of7GJfkCi8yNCj2bYvc+BmbKZm6vdXcxVmtpXgnnacU/+Uc5fZKV3oSqQKfTk+
T9BM873uWuplj/pwsx+fzVdXlArfSfQ9nezoOO2mmu7Tzbo4sDICB39Efst/HgF3
SXGZnz0zgn5mB1McxJcLI9iuYP6qx+nLyN3Ovh3ECDpmegI/gO05YGasK81fG7wL
LMKoOfafy5eniL3sNTp8Ygx/vIK8qdSjvA4RbRogO/uV688s+8tXkeTyqADjxzMg
TPyle+v1lIy1cHamaq0fuc9S7j3igw/Ho+7d2OOPZzUGmRWegGq5Y0c09ixcXMhY
2yVAvVFI3KgUl93RJeMKkP8pM5SCKFdDUj3+kbny+iVwLl9TGhYdbXKBD1At54OM
F0QYhWo2XzyMhhlyavNnDX+A/DsSy4sLLUTfmioZlFriVbSp/9RCMNFMwG48LrLF
yRvP+y0AmBd+sKTb9JFB+FK1xUve8uJCjpcbtl6zvYcdv91h+87+0PePrDVw1nd6
cWYrphf5yeWrikx2nfxWbu7n5QkrWd7qobExUJyeVYwFAtq3F7vx9UaBJwvePYln
c+hB9R1PFNyPIFq8JmnHQzJDraHiO8ZpN8IIy3/5HPFYmephEMZ8XrFQu/u/IBxx
UPaqpm1jEdeAvAl6up0SpsLdlWnfWk70NrBk0ttJSjSnIRKKdr/TnivB6o1eXxmO
/Zl6gIpKA8EBXTDMriBoFIY3WOMcJGRursnexi7NtJXMoG362RZnVhSo9MRdaHxy
Un43t9/CPxijHC18GDFkHaKXGP59eTtUPkANDgEB/w4DQrc2PTiotP+/migLIGVf
U7crLT/9WS8MsMl46t+c57WdIADd+Z6AR5Nr444/57/22R4Xe3PYhjdevtckzlUJ
NboVhzYJp7G/AoTB2/0azoaNJf4k2yB5KqvDpx8pF8Sbl71/2rNOPBUVvzCAbtXy
OoiYiTkcozs/AgbH5VkS3BMJWQ5vEg3Vwhs+KsefjNWSxdBohFpmeRpuvPhfl/F/
0HRnHlJ8c10V7915h6hdbCY7vXRxp239gV4ssr9hbFpBTVpYYOPP1LtaGg2Adpju
`protect END_PROTECTED
