`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
paMVEkNgz6H5pgB409mJrShH0h3tWI7aCM9zkImcJwusw7SX8aAX33n9KH5Dpiz7
D60JMJb+cbdNxzQMyR81uHNnZD/t2nde3qO2efIgx1dS4b9bde/qlRw/SPc6E3Fs
w9crweYjZwx/x6107GQW1xBP24Cr224m9FJpowymnpfuHNdB5HEWZ/NajwByusPv
Nq9l27k5ndiJUGKPGfee2tmaqUSmk2XR723q5S9WZ8vmzfUBn2+pSIfObP2psmCX
D6aw1qIdgphkM7Zb+DuUlN0xUZlpN/GMQejGAfxCkwkr1i4X+8aF0dYwpcw8T0vr
Wj/7FTXcdS5DslRFV++5D/KjWx64Zt4c+aNOPQPMvaqPlGmcPvm8itii6/j1AVcz
eksTwtDtIsUtECRIhfcXNNRogeK0sgOoh80wqKj5zR+jXL9reJr86tHaeoeWtaBe
DICAKhZhc2toRqkZKYcZ+0LYnFKTt2URD7MwK3jAM0uuTebm5RbluhGWFVoDtpah
ivxIlSDO8uPdM/8Ap0lNMlty+HGhmX5Ies9v70prK45cTqu3LPp46GwLXV99yGXZ
axG8AZQI7YzfdSdZ7VpZJyMcRGLzz1lhpPZmxE30Exh+iLBL6s9PGJE/gKT9UwDB
Wnafte/NnjZ26ij/x+vD6J3swkw62j9pgHsvjf/PyRBYrxixl77zaLFhh0pNFiAI
AHXAMw/i773LHg6z3qfM1hxdEHoQbH2aF2U2Z6xVcqmqtLjJHVlbgJ9kViQBHha2
gLf5yAMKDPbCvd63ToHUe20mstoP6jy4JG/cDxNDs1IzLLDC9YhQW0PnP9kb8gCV
XSAduct2aiGIRq4mHO5323R4sa+oY2A77bKonCXJl5cp8+5uHDQZH1trkGWElkWg
tP2aW9hBAm6NlCFTMdHRJy9NvnFoTVEpKB5aIxJ8NFCzUfV09JWCw6MriSgBNpHO
Wvs+GjGMeT1iBDaUQTJ/drKs37WTCjVOHFJ518d4Ei2aGEYqvFlz6uIqmsBl7Xa4
NYFCvu1BzV4V3p9V1EXn/kFWMUhHS0lLuLFr0oURGGO3cJG5ZV2SDiP0f9h4s55M
3OVXRW/Hc+jHII9QAw55pIg0YUxjgIbxpWopC1G+RxTTlyG8zB0J8fNOx3sP2CaQ
ZYsBswtSiEIPcYtZ7ZCpoCa+FJCM1rTSX35R12a4CNvNZ7ri4N4mWNpKgZd3Ns1V
Lgj+QEZDpMwop0tCYQQG06KvR0YZl6cXL9K/YzoAjx3B8Mp9860C9rvnOPpKJWsq
geIOn9yjpEirQ4cOZIMyNTqXCJDT9rE8N/BZjaa9GibEJ8Zfc/K8QLe0OGRsMbXX
V/BIL0/mbAmOtlFbR8ngp5peBE8FdSkmGThgvN5YlzKQg2EX391yREts9UVKvH/Z
9gnvfM20olT+i5KALb4zUVVL69ISaZrjrSr7ft2sk6hhDSnCrrsjMPudq8I2xjUj
nTpT0RHVb/TkoOEp33oLjDfi1owvdqzNJBmp6c02Cuqw9S/mbVJY01C26pRQRGjk
hjEUaFw1U1Qex6OQeYB1PFdVnAMMNxVG29hMbp/5Gn7cKn1DBrF/V1DZZRK2asHc
tk+IBjE4fZoTjK3oHsYLYOIaIMMKTRT7yQJh31Zv2W8LPsUKVivQBAi3pWR8cxLF
Qn6g54xQVKD7vSo4RBlgPFtv+juhChWPbybxdj9BgLVhQYeXmLNoEaw3bEuhNxgB
YTMLR1Bcypp0bJ5iGdO4609pPMacAloK3W1mVO9FkFzUPDBiX1XV/8ZE0/hJts0i
mpz4d/E0M8PEg9NS4Kk++wknV7aPNmx7g9Tl6wcSaSmoswQlNyD0frEaaSdLBMEP
ffPMMd7QgUvgx55uF099NRm41eqRQd3f4vjpa6rNfuZGDtLO/sRUZw7Zg+uGK/AK
uJv+K94PhKO6fC21k0fLsGOAzHj6OW0cT18LG0DdDbx0FI2OQHazC/qm+yJKQ24t
TA5SnENcjdN3A2XTyhsCn9HU0YyFhUsvgsyMdYaR7VGOTZHLuewybHfU6IcSw7vK
8BJspE1LNG/Y/aeNRhagl/pHduTA4IXa+9qnno3d/asUzTJjxo3h1lKTycCzTXK5
TY20Lk5ZZc1QVzEzPHQeOIupOMUR/co54Pz+F/Lo9vw1CTPK4Dwb0jlXiLgHguhk
ywnJpXq7job1LCnIg41gj5f18fgeuwra7HnOL9qkSH+VS28ZtWCs7NSfaZ2Mgozm
51M+bqSAcw7wDSxFfqkNfNrJNo0FJWAsQviJ/fGTSfg6bTda56JePt7Ai9npacYi
aCwn5NUhYRA3S+NiF9ukaKDk+I5oQljIGoNrSp8Y0oM=
`protect END_PROTECTED
