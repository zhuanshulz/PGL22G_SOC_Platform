`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H4IrIeD+SMyTSM8VRQnSTFUtstvGmTdpk3oJ9TqOCZQlPR6G42Fp/5PhskeW5h7g
IhaFMxqAAS3VUETl1iKVDNp8JqsuMSoVFyWXw4HknlSKPWpSJ+nJsxCUF5uDApvK
GkEtz5gosJQhXltHoVNk+fiyYaXdPE6n5G8UCc1s4tbv/X/A/ZxysHcTuXdvBtFM
OcXWRemtohje6CCJiCFSa3kOIROq1CZlFpUsYckumOG19ILseMv1Q3h4V8KFqd/S
r9UgQ4pdPGBuBg1iq/ewLKf/cXww/WSTMxhWpoLUYLH2h4o9aS+ICwNJJxKDmp1A
Ba2XWFetwo2RomoHHB+WLa32n8T69CLXRYaxvcd39028/AUGHlXE07hIKWayHrAh
oTmVwN1djHZKzVpmyweT+FJznczDbjkbj/PkuWoKLbeIcnfm2GtYGQqtP2ZV0aJ7
n8vTLUJAnPykp7ShJkU6hO6dEr+NkR9XYCKTblh73Rj3eK16sQ/QuzN4fF9IYjkq
nYL3YCkLn4pDJQE55NWE4l6rCSUh235IidocTrZuqCrEDGAYDmJtbzkb2N7Lqam+
VYKWTvWsT+enmcW2P7orORNIX/Gvp4zsbB1u/2HM45nTelIndaLYXF7USHVqoorT
47n+0zx7UtZ42eCa4zFrYHqnCW6iJImZ2QMdULuMTDZ29xzeb7+9zkCPbJeppZV7
cNClBqzHgboRyj5pOCLun1hkMxnIatVmEqL28Ko25uHuSaiD0Ik3qXGlHiWVLMjZ
q0GRM8kjOIN4yGOs18KbXlWBNdcp2JL6Te6t5m+6GQFPhp+CSjHDs+ygQE3FaqsB
3UQ6u1eHkIcq7oAcylhp13f0MdxDFArdffpvADWoInT3NEuYQJjuLkUu8ultRxZD
fNXj6fmcBMhu7B0HH56G7loMhYXnOIegGUAjU2hRrZEFeyCerJnd4Bos6YUM7Kzg
S7+ga8/t+pIhNC9u/qg57KqLIRQolDVjS0QNDwwqgaVkD2uaUfxVuz1Tf3uqH8Wo
qX0vqlliXs+Z2Q/03mmI0Y2LgA0Blr+ApAH3MIsZbQjkJ+qbQcuhTVCubbY4zmjn
2L94KVguTsgqzrTIo4sVATf5GwpZVz743/ZZ454HpgoO5FsmnCz63RnFygrX9/SI
ittr4CnUc61QRuJn4K9noSL7fw1HGC2k7RXPSPcC4844EjVZijA+4amPjfCfh6qJ
kRhRS0wQ9FHWjcvrwTEqhV98qZjlBc1IbyPNtt3vqfSapjPz9+fS4jQVE+KmLZ2c
0fEJVd06lb5CGV1X2bua+6VZkpXIvzZyWkcDhL+ztu0=
`protect END_PROTECTED
