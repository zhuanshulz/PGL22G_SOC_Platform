`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lS6EB9n5KhMDkpYU0u+NsBWWsmJQK2pKYZwHJUqs4vfY35Ri3fKW8yYUlL1uzhkD
PIvgxdYhccZ7fcGCoNo803ayt6iEFh4eE9YzU1odMgAZPEBXxqXbdp3r1fQMyrib
a8eeg9mbd9GJYA213JSPMfR6hGadXnf2q5tE8Avd+Bo2RlVVaup11URTeMDgtxia
nrHZ6LPDKgF+SQ5RB04oKEZ8Dlplh8CAYCtrVmKdy9Gm7vsRetriTCmQBIyBW+tN
qUVrvdsdXDXj3NO3G6R5DkWEJzubs+kt5iGgaf+A5IvNURdUHFMuJQlgZnTGOYHN
g1rUaFLncH8jlZ9g7rTnZfSR7h8im8lKuiLwd1w+LmVzpsxHKbOH3xs4/B96ptZM
/CdODvNdS16BzlpNyXuKUBmsLq0v6z2qBbMtPz2P05Owf/wnOXu6xq6w4Ks6Q3md
25WeJVFM3HPaaMAgzBRNr251Mv8BV+fsIQoJVXDyPUd/rGqi1NmV1Vsl3NQZ1ZEi
LNs1jwlKa91ok/3Xw5raXZc2vHtRGlMrDT73ttJ8tSqtN1AtInCZyCXgPpRqNhrK
oiYEmzrwuMHesTZk8v9V4Tzj8fF2aqJdshONj5FwoqKrb5HRa0MFcVbloSeGl6q6
lDY4mU1VEsNk3ffvrlZFG6kjTv0a3FDIEqPl0B5OPKWe7AhtGZ7yWD3UDAoECFb3
cZSzKrotOVaOvJTmsO7+rc2/kQChOpANgBRPKRRCQwdhaC0rQhRr3oTNPzZ2hUlw
arB77cAAcQbatGLqkoM03nhD/Rjm/hhfXWNsNMVXeJ39Wzuw6DQrKMyFYpu8ED0q
cdVwj8h91aDOGlLWoi5irXslMwMd44jWvdA3YVLumuMs0jcbtHBLeem7zNtvFFsC
ENKM3WcAgTJiake+6oAEzdlt9ouv5eOLrsQgf/CYyyglPLAMXCX3XQ4WKkE8+0yA
zmY0e+e63qBoNJaofU7BwP6o/rbEq+7q7aEkw9yomJ2nhj53TkkZ0tcSK0Z3vg/M
tnQJ6B+YFAivOqLlEA/xU/H/DMWgrDy0RMeCybrelcJg87yFZ/13jG/hvIR7pfl/
SnWVQSnZAyquH6ymvgTq/CEX3v7pL74IY02xPqOQF1bGUQAMYlZRUOupsJ/GZFEc
xWXdWpMorTdF8u8ePBOBfQ6d05RrniltSyNFIf64unYKCMAIm1gTogqfJWkBQOfR
G/zZUI3JKqR/4wUppRD4opKesFkt5E5bfuXbP2fd2Rx4QM7x3Swyw/4zZTmgfMOa
7B1lrbXerjKv0fX1n3pFgn7kZiYpaykhjL0RRm6KKh/BkXd1iUW+xeIgfc4NsMXe
CpL4lndy24JqmC9wHi3K7n18nGFoXwQuhCMGkyjJXqZ+5PwOtuym443PtYCFvIgG
BFzqE5O5HWnvElxvmCIShmXvFia7aTes+r5CP0T1Voy60UrhVOZbO30FuLnXfOwL
y0K6+xGzjlT0p4P38SWPhn7eleMQxsxw9JVqROqzfXIjI8vGBWwEyaG+V7TTAtok
X41HXXFGMP5BX+XSntirkYCs5WUkHIlfteW0PMYFLyRyeRotjToY7zVlQuMYiKSS
sQ5nsBQxwVzVHAcV6geZjqzQPqX7kWBL2A+bf8MIS3dPvdppfdKHqEckDH5W8x+Y
zkjxUjuS1bPdehlXgsZpzA==
`protect END_PROTECTED
