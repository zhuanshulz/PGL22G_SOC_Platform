`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Al8B+a33en1yI2Zyy3MOO4JLOebZIb1eCxsM2gcpuAiZwz9v/VE1RG4RFbXXaqPF
Go9p4XGhtMgQ5SLhOy9YFttax72B+fEuHFPYxR8LrdMFF1fNhp7fEELpMNP4p4r3
YSlzu1wYmKFVXfb6pRMQ3SqaUO7K4VQskEQGqGhHZDNAXu5QdDuyDfQquGjrV4+E
rmPkwxrY3bWgeFgB/68nyq64cSP5JVOuwklw3stlMnecGIzEGNKHQx7fm9gdSC86
xkVVfIJr/ZdC9RA25n2KvQ2aavSIUFpgAyEyRiz6P4fT2tulqK2xOViF0RcUxTtB
sz17ERndwEYNb1af8uuhJnxLnpy8NtVb4hDVads97Y295o3/4VCwQPrC9ALgQDRc
oCw1RjbaGTvd0JlPn6jRQoAG1Lbz2biN/3FHDH8m5Bur+xMttZd3XzrhWLMpGfPv
EJRUvc6B5130QMtAPJRh2fBG064v7HQMiPDdnKSPAA2qhSEcWDjNzTT54kxNPpQ1
M/lAV43l+Eobh9Zj6ur1uU5QPvkK/pnxuCsfvft7NI6EUp5sYTaWPLlaGAfDsvAx
o3ueKsR4U620XAiwole2zK0/NW79yjgsx3M+wu0Cj224NFMtATqyFOpg97KpUZjd
3HLiZKeOPrO70wbTRknNimg2gYiVJS3FMtX2z6VIIANzZg9jJi2lLi2MTrPbmYS6
D71m2UcAeKjnZ1+aZO4mjJK00lBERBvbK4R73W+nFYE+8te81CLKecA32ef/q5Sk
zMra68204d9LXS0W991UvT+/bbmBX1IEP1UjXoMIdP5DhqUO8z6rab1v8LaAWnmX
OeLAnbBGhMTt/14jn3EEKPf0K5AF0Z1ND8YR3HfANd7V4QdvZlp3VRRygpwaeJOb
hFjNALenJ/py+kPdZHQZyQ2psZ8kjwIpyMQG7Km0TFUfUP/XY7l6H0P4e2ywTdSM
+hH3ke3C7Y2jRfGP/MLXew5ESElPyuM78sCWIlxhphXVe9mwnACa4ZkHt2bieoyt
7NOq2jD7ZraQEHPJkjcp9BR9S+ubbNFuAUyyCmma7WIfYd74Ij+XksegcHGllSXW
eGVUsLFIX4dMzPwHF833fV8UQ7FuLJ92ZjxRS7zO6hN1YlMVD3yKBFehMQUKKsJp
UGge9TDnAE47KK+O9pr/nJuhO9VX+ElCHDHd8GZ14AwGrfYZze392jU1DUBGtOZM
IWrvOWjXrleXlW9JO7aRw/fVicbHxt+rj4CvL5QLfl6a0TrD7D60ShfI5lDQJdoi
4+YYBWW8ziyyMWWHsgFYWPSGP28YrxXm4czoJA66wGJRnqQDKaH/cr3oDqaHjadv
MWdTiUP1ipqd7NKEzkPSVbGZFqqhKVcLg2vvuLx9i4ESN0E1llBBBGeeLtghbgbl
NyIMqCS//fDtrcYieuxeEvVT5vpkMty6rBi/U+NYIJF6Lo4tgS9Cxm4FRdy1fuY0
36X/6uqeX99WwMhv3d4BefFc7WOp4JFxIWxv6B1TzFcdZpZmCMNV5AasX1bBBy6c
pukvD9Zw4ll8axi260eG4vK/7dL9iLSbkU8EFCrX1cVHT3kOzrfiLm+ekVAmyLRL
xBUn2VoROoSdGiuV6T0cxnQlFOkw9DC08kMkbXHFUxbrKGDkIOBdrzLOcxYFPkLB
XSdCH9qxpTZ3dGK7p/DrFnS8L1Dx3OIzg1gKZBvghc2TlixLAaazLmx+WTOrt4ac
zcjzRdGANdlRM7GQRxG+XV69neMBMgJpQhsNdqdo5+p/YLKKkuqosx5scp/nRr3L
FP67mKYmV+ia65EnZ5+IU50N1uB4DFMIS2EMmgLy3zzeMotr8HYrDztV7AMDVLQd
jnTpseQ/5eK/rDVIzp6pef1JCAJ1h8uo92F2vDbejGvYuid+QM2iii4YMYgf3PGS
ulgyGSRFFnu9z5brmYGCOFFSXScpI/cQ9onODVys37MOIzdJN9P+ddJnYD4evAQM
Zmftz3atNTOJ9G5UpY+izz+7RAw+TvRYF9cf8nKwpeg9cJKROGSPrwt0TxRm0WV8
NM5QJ7u9g3tAQ9NgeI1wo7wXLnKv0dJxq5AgthlFrlBPd/jHaaJvenkfyiB9U5vP
kmwDQAJpnJ4VRj5au7BPCeIXn1ac/wYQ6OWnluWlwIxsnY1uiO9MStHXajRSxN12
bYOx550vP+l5+C7h/FVDb7JT8Xn3yept6ND4popCcJtIM6/dCF13ybhTBnw3Y4v9
oSBNo9dj4l+EiGIIrpnFW4EjSph/HBo+IyRAdNA/pa3sQlYewWgsyvlOt1vt0+Qb
YnawBcFKh53fMk3G1mXcDYNZAhY6jOwoUniMSDWEWUPYT1mcYgtEht07QnN2WsCc
gvLyZc39b1Uf5pVx4KE01jhdrmq0qbGgH2v6Os11PXEB336EvFvva3hn2W0hGJch
ebkylHj3I0eOLo7QexebvGlM5ffufjz67Zwp4tkpkDvinf/2kxpy31EfLBJIBzen
49YodOZBfkIbWRZiZtACP3HfYsd9y3Et9rMgWba6ClePCP5vuXS9irm2c2+ooy44
ukJ2Q9/b+/0m4sKkeR+/8BeKWFAQZKtg9ub2B/rdi8EwCOknn/slpn2Zl3Mq0Gy4
D2oGP9iKJRU+4kGJ3m9YPeAmis/nKhUO9HoQZYCkiq49oyUSS0TnATcWuqToBpmb
0f1BcBzw5trHlhasTb4ZiBVgbly9FA9ijveMzafRAVR8EDEDE5BCC6Xxl9vyw4as
1uYTNJedc4B3EF7DDAKEgKQTtTh0R197IHkCXG8qQhJls6z49f+3+tRljmT2e0p2
Ojknfzc36zlQXA04ezTQGflUlyO5GU2b9Ko+8Bq8nFfsqRcyNHnZdesp3SzhOBfe
jJFqq0vEtBS9wA7tQJabIqCmCZENuPafIgQWH1Hh/2eh9jVt22D78eSn9WdfB1ky
5D9ANmk97Y4QcGcdtvA5PELhkMq1lz8VkCRdKohh5SHsLYidcrrCMA3I3RdmhV8W
vfLu50ym97+7Ll2AZygvrGMAEPHcrY//j3T2NE17t5fPf1GoJS/peufqaiPBUKaF
/vF1Da5ebccJkpSkZzL0ahdYpaTfKcEzuqgi8+74L3l1HLFjgei05MZ31St86GJH
4TDwscQlNYTwuBg3+hhUcgzjDbV1MXgYZW7VPnZ7oi/3azTn/7iR1PoNjPJOLiZd
pD6+j7qKBNJRK+xf8gc4u8gwmucYem9g+YTm0VHvvjaXcusqBrLHUDE12fbjXpSU
m7eWeyeb/i9UyA12UqBOsQVhlgTQFuc0hcKXy9gU0OTG3BxC+/NbrmKmSDwCKa54
2pS3b1u0c2dHqKyu1WZK/QxtB/wVUS5zRYcqq2iDPHpjzYqZJxYNBroWGxDR88fL
Jd1Xo9uzyIMadIO8XaQ/YcBmiM5CfoyA54PQUtZB7dWWGufXdN0FxlsLIYbyKoqj
2Ul2LUVAJHGRe/bDM612TF/XnE8e4JLG5VlWoHkMWYgzMOJRQHG14Ggr1nidTpT5
RosGpsFPqk56lp6LzrqGpPawcKPFYvs3CWm1r8jpFziVzyPN60xZ40W4+zAQBl7W
Hi5RmmJ9bUmP+Ba0oPsaopMLwXnaV2I72KfEuQU5Sb17hBJU+ZMYz3nh8IFnYQQb
AwMSJIIA4ZLAtTgBRwPwh4076Zc0/VkT6PM0AdstlHmNCz6VP/davoj0Jp55HdzH
89WZBmpat/q5DLK6DK7HUMbir5hAPQ19VrN0AT2TWUXJNldvx4mb+53qkftNDIqY
F2MH4rmdKPhtRNf66RI5gieY+B3MuWeoq5fj+33ucPIVKS96Z9SUpSVKwA6KnZZd
`protect END_PROTECTED
