`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dxtAYNw1hit+Ov+GAC/WuaWORocecdSdUHEMGVLcbDbQ8yhTysSQqX5Guuvok7Jr
2mGS/Uw6G5zAu16pDVmHLPdIxLtLt3b6CQo5g/CtyhOyeRqgHS9RG2tSJ6nwEnvd
2AzrnSIfcmDuRka9MHweJbRHu0noCHDKt8t3FuDCbbxmiTbt8LUEebYlrGRIp/Ap
Vm6AdqO1iHn2bckUMYt72SjH39hP5SCmM3xt4mc9AbuxLWwmVnoxxf6T2J/fWOQP
K86ojx6yMPB+Nwkn+FikhRir52PaW3jXZgQCLzmepa+qUL7GUXXtB6aLOocd7nW1
EOQL3Ybxw/YQ81QmkCuBlS9jdMG76UArZHdz81ClW7TbdSjQ2BaNXxhDxAtolcYJ
O2frJqdmeiD+pbojsKv2qF39krS1ChkzDfRy44Ki0DuCEP7YlKnm23gq79vtOMp7
YI1110mRkA3DGNwQceUAN6vGjoav4aN7x1BfHM7GHHE=
`protect END_PROTECTED
