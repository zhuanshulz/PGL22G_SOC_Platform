`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j2RkNG4eVshFZSBzKsL+PXy11hqWTPeTvxjFz2QVlpQwN1KnaVyIjxvHeaAWyWXP
nw9CLcb7MSZx+PRNGrmMzYL2pfGuNuuxctxW1B7w4uZuP6YUkdukIOXRkAi+Ipij
GIx1/RIhhFL2/mugWJsTwG9R7bnx9aWtSnHiz18hrpA+E/WJm9j02hNw0abZ2zvI
M44N5uNzse4d33yni7tNMCS+Bphws2qjkPL4O/KNSK5DeDtyc8PBMSlobAFka3YX
dAOOFGZj/sPlxulC6FZUkwLeKdDSSIBqoNKpUnF9rky52KgETl+/cla6dL/0o7aY
Dk/BV5K1aZX0ho675icp9f8vxPa/SxwMlJwBwHfnv+EqnWPqw72NEFrbE+1gfbSU
f1+gD7wZoLTHNRyVRpa5KgH7LJiPHAHq75dpiFDxgAPr14IpZFZ4Xn8GjFZi9JVp
5Y/pJq+BFwXEPLgKayCweWqDAb7sO9pdAEm6hFk0PMc=
`protect END_PROTECTED
