`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lYcQfbaH6hCBMVV1xwJUXiHrXXlmRPMv6h81uchUd5EqYLZHZxG3Me097bsQMdBF
KxcQjdJ2mUmbb0rzUpYpW89OEn8kju8GyI8VwSOGvh//tjy0SR9t4JM7J3u+1jKi
OXcwl8Jfs6i47cNUZJFWQiCHEjgpQIYvLy9oPHAtMQvwQkcUdAw/VXRIQuInkT0N
421iSTZqldi2MLOULGlFfR/HCuNDeYWKrFxpf9O+bQb3PBeX61SHiE9oP/Axufst
Y6vPlwP5a4PUOJbyusIX1bFHclWidQsvnerQXGdlZxbZx35qkpJauwFCyZwRrXHB
1cNQlm3BSVaOYPss5sz1B6NQrGxnGLUDVCHeDM9m5SKkzLI932c2lvwTuwFDCmtl
4G9p5AMTqj72y5iMyEydVnlLbGdl2kafiuzo8YfaNgqBE31SuCN+zfVVWfUynxdQ
53prR37YR4T/qXRBywrCgjH19Qh2rUPaGO5MWog+3+BCLsazm2qpeBjasYyuhaXB
d4a4E9ePS3o+IhlUn21FFGgKu0FTw099EKoUn6h6B2uHSwKMmQx6cc06V3DQRcFJ
otzly8EdBt5F4ggu3dUgl+KnvmB1WKNTwofGJlK03PCfvzl0DQOpN3RMzr5y6Mjz
DV/eH+xDufH6R13732DThw==
`protect END_PROTECTED
