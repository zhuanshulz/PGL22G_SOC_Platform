`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tt1uwTB3Nu2QpkuHlOG/hEXJuOe3abzGOephZJ+P1daDCao1dTGZc1KO1Sc8cTak
LCumUV62mW/cI75qBQ4IzwuCVouYkESrWsy/Nm4CkYICA7dSOGQM0rE9hClMPZr6
sHhvqw1FdsVx4sOZRVHbWwtOwnL5Aigw85SXCs3+ql4rrbLRtAad1O6K42goGlFO
iOqpNaJwsOirAKUwXbKATsAxAFVjHx3229/qYiQuN8ua9KeXF3bsk/AyJggiM4f+
F/rd7a4CJ/NIXKQbO6OPvNIvAv+BfTo4CelvVYNAj5O1raqGzWAHkTzPAIJYHNRQ
5yx1fZjUYz1OXdWFvsfr9xWt5N5sdPh8vEHs7NKORV9t7Fh39w6Hmc3bINV1lWGC
Z0EMpQybeuULRu9IxMQYZ1m5HNjgfKWmiW9mVi1Rj1YLCrjSUCN/1pQH69W/Ljjl
DrdPyBNM2OfT0kU7b+ffYXMETOAhzcRmUBSQ2G67wniBWlAtzf/VQP3310k4Fmtv
1MnGYKyts2GrGh9dgKXe5+rHzZpJ3DmH2TOixMWNqS9EYfjYlkqr5i9t8vG5JCs5
BnGsWP2OfI/R2C7GPWyCkuVCZOlgvkR1DvLheXxNl102vnCgCWNMZMDb5x0nVgqN
AP7/rbY/tZ95oy01Y9q8RI5vNjsQ9TBtaE7LB+sjH4OrHpboPB4FUNe743+gOnfD
fKVqYwjCB7JdJAs0ZbAkTSKgvGXfP8hvqCqe5ObBjzIA5uQGzlZd5Cf8HIK+LGHF
QS0Lkb85UAgd21+HUaYdIHEhQuR74gTkgkoHakRXgLQaaE5Ru9v8lhbBmmsoj35f
++2aU4tXG5tHZ2tA9oPoj0hzes/s+QOcsy6emm8nrkMOPn3X+VwRxYAe8aWGEw2g
+KS/dYLuY+8n6zBmKOBKzMFd7V2bG+tC3D3UJ6CeKtEnFrRDRfp0PZcwHTAUDNGy
QoBjhbsczIIZVAVrE/Fl9WG6y/7GLXr83Rk3OgEc1MtjvdiiTNqozdy57DjMKQAj
WCiqyE9TLnWA+Deds6JmTxL3z5r35tpqVo1KNmZsQ5fPoDUFJO0vEXpmQ3d86yvL
VmaR1Ufc5mFQbhuBSpNbmfOjF9TKpHAtsH/KUFsuJEkz5AXeOD/7oMYWj0r0KL2u
NjoC7VC7807sXJcWavnJiqb0xEESEySX9/cEvT40vN87/4NeGEI3OIfNf07xTKVA
3Gu4QRk26PjgXRNrejaRMvQmNc+6JQHgdH3HK/E0E4rOLZPbI8W6X8RVJdXwPfXf
popc1ATx62G5X+1HyDsi2q9qTHqvAdkiaNQzRdK4pGV+6ExXPXBsDE3CPR9qAi4O
xfe8CS4Zqkf9PWXp8vZBXD2vYT2iKEpD7HtowFCbcluwyUaLwv9E6LpfaMPbx+M1
2+sbgV92mYX0GCq1I3fvKK4ZTQwiEhE7etDpOdFkT3LQsA4BObZQOvdKpEWcqM5+
/HRR3n/Q770kymjV65JmPyaTMnACBYJd6uahTsqwPZzCHccTYPpfIXx7rvGTA4f9
P732eF8grpDGfyOHDfswv5+qJOMjIfKDLSS7UXBgJtGZlaI+l0QhUqqcF3O4M8Na
ynnhZ6JWXfzRedc1mjKvDSIEIQ57vPh2d7gX+BOC6RA0lHPiFPpVQDCu06OsqiBK
YNhusYBmEn66MkvTLDajV6SVDujQgPHz0d4kv+NqfS8gGlLaQWqLOcUKHUwcZTox
N0WPSPi+f4oxnxQfc5KmSPCizUeGJPGiod/Grbsu1+ybdrRZvNFqfx21xtRPnIUc
mwwJLPOiCA6GY8Jcp1EU0q649OaSe57LXHMFwUII5oyCUdIoGpU09mRTkGTBnkoF
SgsfarlAKqkLSwTRyTZxwWxyPnFRQO/bDXsVrgJWFCeVA6pQlcE2SixrTz1DfdKz
wX1xhCe2zsmd9xxhE/BwiDw2iqrbhhpuvFhfFOl9MBrouIzL5kX0VRQEwqFO8MxP
vfTpLk+stkbZbuzr0Vs+tel+At3X8Cvcu8ufVfJkwk19d2IBwdXG6AhjxnzAjf/B
RxqQ4xrGonXKJ5dzvWZcH+E6qkb6zNYhhqUhz8fxmLM=
`protect END_PROTECTED
