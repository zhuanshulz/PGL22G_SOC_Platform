`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S/N1PK/RBjVM1lSMM4gQ/+RolfQ0k+WgHkbF8R0JpQgIPy6zlVyEQu0RKziq6x4l
x49KZWS6GBWS/C6IzhfRJprKMmr3JIH+3ft/6BAgjSFbVLXAGm86+EIp0NOhrF5b
6PVqENgy8Vd5Im/RH+8bont3GY63WPE2upcmdvpWzoc7J3VN8fvBhRig6rxL1czb
IO+1MJPv1yiSaN3BYL/OJK+mMVUg2LVb+bg0FG4BRI2K7VMzT/0zD6MUNzACuMkA
wtWcQBFHUuhZF4H4agfcwEwMRP6/vBd5+YPxbXEUjbHqvA9XdoP8y6z5W7t9xJIl
xZgf6r+eZpyG7taUlJIKMUbs1TTdonRn3TlboOv1zHYC0W6ovkbfQvI7OyMf+I77
LrT89wIy4SLwNdX9WMYt9kBB5OcMcwPu+QYwWgzSjfy2FhRScFVKo6lNr7mFWRsW
xCRaijtvH/cZkV0RFPqo6U6YeyxeM20jwgwGj2DYLhU9qGO9AjlF3jGY+purYHw9
tLzb46EFFcB6M+n+tjtFN1+ahtVYC566W9OOqUFw/5d12ykAv9lBGtp7IWPYOhuJ
G4gYJV+3nzHJAkNAtY1te4hj2v27XyH6WA5neWvtOpu6xEOwKdZpD+MmufekfQ3Q
C2oGbKZoLL/gTc9cqzCa1/eBXe0VfY303xKHn4Ppe04kmdE1bipigINsl99ve4Ay
Np5rlkPc6bdYzlIAc4uwHLcfye9J4umJabGa4EHaonLU6hwl7N2M7qndse7QYQR6
SzyCVLXpgaAvTJ/WvPcWYQ==
`protect END_PROTECTED
