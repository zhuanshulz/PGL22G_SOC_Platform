`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a+53+q0zocGKkc+unMhaGQaGHrYg/u8/cvjE3gcxSrTu9JLvMmhXEnMTBuRv3YMG
d3MXl1EcxNXREGXJu5gWtXJ4MoINranyELFYLHc7Zcd+9DIpyaKg1ZyHznwwbk6K
+y5kyHurqItHHxu98DP7Lvi5OkqLd++gHJGezrsk36sLXi6wEmqsyNpyga2iAUvD
FRrd6IIZXWp2xfyuUNwNY3hf3sopNwud3CqIvMN9kK8KbAuZASRlWXetF/BsDZF9
oG1fgjo7XZrmNx3I3rQtaysFBEmhFXO1yTC4U5VdutKUFc5p+knN4SelsBfKN5uG
8OjsvacGJDc4XDgzIsiWKL2Db7Lq/031rOFBbAhc0iKZBb65jH1rFDpJByhxafyi
yAUg2CofJf8ij/MJ+DiNlJlICKEXcmhkf7g3aY6r0C4bgq1oQKHJbZyEI1z8T+Oo
PHAy2n0GAonwn5Vk9cDILet1SOaI2sMf0eFs52sUoa8nC5NFUZcI5kCb3Z7BWqmz
DlulU4KTK9QA6c7SL8Ycro1MWe5dGIc0S7jrxVsBkn84FV2H37SmCnmwfoCzC68g
XSD9sAxeRDgnQCjXuOzGcwhoZTYzoKxOdE/NhVQJNqrQs4ytbtWuepA3Vyj4H2MT
s+Y4WJatIEMNAwIlj3nKxk7mw5dXmrlTigHrcwsWJBKtkEGr6y9Y0KDpjYfvasEI
GYVBeR7N/YUcq+BgTeqHtjHiih9o0ZsxxWwBeD1nixNWltBNJac3JUgBmm9PyqiA
AM96LB31Aw14TAc+mU5tM8QKbQiuOOofK5NCGShCXeAd4KuVUVlptQuhrbc4x19v
qJ/m8ubSPzdClljnbO9A+2UUN/uNXY3MayFo95YY5Rg6+HPOPeKWFESS1s+Q1XMQ
b34PLGm4o8IQHcEOiYMs9yi/L5rQvXMU5pL8B3Mdj6YrXo66BcS/WC/PsMMtwHXm
fPS+MscqVYAxGPD0QDbY2S/MAW8e1aInvnWf760jdQ7oZoXIkQ3227SZpGLH+X8J
UGYIGdGW0A9oVsf2BGKAXy8sFt/8anejWhCp+pPxqAZWbjIIpRP8ju9V7tkkErON
bbCPoVd2PqLJu7XhX53DjporElVsOwdWF/fSroiIZP8sXyDEj8yDMar6c5GOnVaV
dYH+eSVe8Cpn+LEkL/+dED1e4fOrQSTjlmzmmFQxLTyL1dZ9qc6R72Nuv0e2pCWY
10L69CQqRsMS+mldMLmlw/CjkGjp3gsY0ypcjgNR7wqStuuRjStXNTzW+QVE8A0o
rUKHd9lkh9g5rVfwEOEX8nTb/IFgwIucunFB56ZeXvu8CteGMuphGuAp6Xv6w1LG
QUidHZqt2zouLmSPW89FoGKhUzMBIJ0SVD3FlwvASj/ZRRkmHVrVFD3JOIoCUIj6
FLSHufHatGD99ydl91mR/3gbz89flGXTP9hmbFabwhiZVylmT9/Hv8Pn8XK1NsUA
jAKs4nB6L8dCwgb9tqqqduwRXK0kOq3RR2f/aeYR8tQKYt6PS4qBlwCWU9YAwhFf
EBgx86v3gUwGot04FwrvVeZcA1+FzEVpxi836CZ1p6LeT31HQqfoaqycF/QktJ1N
qU9jG5SAkAIN7psvRTCECW5Dt0HGAUL/5XztcsM+VcLI+0IFPa4hpiv3yvOoq7Vf
gVHow0+0ZmlaFhWzfDp9Ln4Q3w/pP87wFdtq+jy8TGNqeimZrPo9wQRbDDYtp6LM
AeYYS0zBpKPrdJtrA/eWcaZ/fEIUrNScf8R7/MnSEEy+MR+yVchHfNAbxWKRyAix
xRVXElWj3FmXL/a+Hi9kgz8HGj4z6faoL+Bw59nsuZKxlEqAq3N6PeONr0pCx9lE
9DEE1xuViwXt6kHHO7J0Zxkp/5rKBJ9OTnvth+ThRv2ajAVkNJybpkq0JvoI7ml/
8uEiczq2xVIONbZ7EmqduVrnqwbwt+eqgklzLhCv2dpRthghFNG3iShW+f8dsWI1
4EUWQ3LvHVavKu/xLuN3Nq6uUUVtmiHE9fe6Wg8rLwJURnsdhfMAcDfJVBtEJF0x
yehv0kb8QEGzT+EfwpjzlFd5RbVIqMNiHHE7QdKkwqNWwFvn9DLRlEnFKcrcRBbV
+oI3b73UaGvhbifQkfyKs7+3Bfleep77OfWdyRcVLZ7rFI3P/2mAvolpiVkSPI9u
LCldI8zGWHYZUWtJsgFDG2BPO2Xyfw1g0O0XB2XsCD7c5GU8FzwBfK0knimb5iBQ
YtCNOaBstBQ+RQae+tpA12je1OHnRlcPytyqMJPr+H64cTJ7ylJGU/7hG9qviWTL
lPMZXPzKhLUQZLsPrc/5fdVA3TKUnwotVvwdRyg9pfUSt4weAn2T6RPrUJPD8tOL
4tVodNT4XDjWlx6DNNmuDhkl0snOal9rtHrFewq+FGUEcrCwnHhlAndG+d0yC4jr
gcxg3gX+i/JAmhP8i8uz9dmH/pL2J/8UFen6uOTGSELpkIWf6VjfM7nhkxk8wzUr
OBoEV/kbLxXZmMwXr4q+182Ra7h8xp4JVvm4n5G6AuTctQfR+SGNC0aQ9tg7WRFs
GfLUKLp3/zT3xuhUrBOa+Lp26xb7yCqGUjam9Q3tDpnqoVJG9e/DKaKXp9f+Yf5h
TBkD/G3m/dM6Cec3u8aZ1MuXYa2K46XKEhwIqu/YBXf6CrmGKrLXp+WkeF9YASaC
m6naqw0YXPsASmdJ1GkBfG84lwT5VVMOwuko5Vxl4ebgUX++gR+UIIm5uHMHt4sz
M88+3aiVKQgqgpNq7FTDyCG4LZOSx2kNkywy13zQpt1pgOkz/JiM++Gu2wrAQLcY
i68cUDgY86QoJ8WiE5obL8M6trx+nkvDN/8C5lJNxd8X98w0CTULhPKXyDWOSJou
ukRnPCNmp9CYH3cS6DbYiiqdUro9NKMBpu4sazKW4nvv09q3SKBS6f21b0KpuLXZ
x+IqAxDqgXm/h8mCXu5Jy/wpWOH6O7QHjJ6Ee+mJ1zqZXKgVOBgVebplgmVja2xM
Sp47zH8qiCz7ApQo+be51Vodpd54gIDK4ZH8EFSFOAbJxVKmHbjnpdJ0T667xpyQ
o+R2GGBAXvSj6LEgRo75UVyrt76Gj5kmsiR7Cjc3lDa34pLW/+Nm95Dqy3pOfMoz
F6VcarOK/DEsxlICJsN5utA7AsegZeFOOCq575BuzS3T20cWPHzQMSUhvgW8DYdY
gETInuovfKeFVSQicSxLtClpo0aIcWxGGKEddFy+CvbSiXj3aoI8rrHwSwgnZjrT
eWPiPVjnwnJDCw/4TB3dhE+sx41AUh+hm8W8iTcFEof0q/GyfDStWIqPsunMVzyE
iE7prb/2hOl7R8Vst/JDqHuQwaQaa0c8KN8gIyv1mZkFzu7kl2fNlVyjcePgiEgb
4PyIBrGfld4rt8jvbtjs1FcREPaKoXwgWVuUuZgw/YYQrDIkoekO1JsswEwinzum
L4bnAsjHNn7isuoRd7eQEEtqnWYGc/43SqLP3k24ceTZ41SPwgyom/dBi9/r2yZc
zXMurZt8fuJTU6OrvYqD1ljAyb5Dpu1ki//FdpEV5L17cMq8Pqc3iFHVZtO/leD0
cVgFZ+Gh7JF13GZpp9iAyGm6xwSjaZ5FdLTzfDAi5oJbJCTZQYjc/6ccP4A0cgGz
+N/mGjwWA4bq80AZ0fL6EEMwAoM5O9IjuunrAMEy8UGcls03nLUlhb2YGEqPVO1Q
Du2Dy3uugTgQZmWNW5vgSrIF7CbeHsNQdapIBpu1A+6zF/M3NEzjhBLt0SqVzLOA
vW+9IKND6WrUdhxqX4QWmlCYEIOlJUZkZ5f1k8wFYDolL4SC5QJYbHZLyLXVh8yN
9tU6RkHSJCa54Jy4VtJi2vOL41wVCIj82f4r3gHectIVG8ceg6aNk7+kuZvIKEGh
Tln4E+1XSzshS+40zfczdqDykNZ364v0Ty7REi3wv7lMn2knHjV+5hPTv+0k17KO
ZY3PwBbHCH8w7TzZX9ADJow8A8GPE6H5YGOspKXY+46n19GQ4rtPKxcJrDwElSuA
i906Slzy4NIVDSS4er44B7px8IezR5aP27d3YSWvxFmXxDAz4ZvdfCiOQ9Ig/ZIL
V7GlkwihMk8uPmUkZPfHK/PCKI3GS0shTD3arn+ZPYSWJ2EC87sas7Lu97tU5Tlx
Rt5sfQoq2KrD8Yg2/bkbLN5ealWEmcsVKKnPpMTCsw8jDm6pJGimkjxL8GpfzWgy
Zj2boE/TgtTbG2ce4B6vLDdisbcnFNY0VZ31xtb4EZw1KSOb9w8Bo0j2cWS0HTRs
BtyvrbMeWjsRneDU6mY69TNvJUN5ew7v2jiBnwsp/gnSh3hK0FPc0V2NHCGID3F3
HkPv+V7Rf8kPJyXdHwMoXC04w8z5EcP7GMTcfSnMhQabs5jzXD9Fmh/PgWFGt2Vj
fEDmlhxWnwzAIZZRAYjtEVg6F3JntMSA/lPVKwbqig2m40VZzeZDIZ4Rkjb4t8Kn
1JGSiI058s8j6QLru9c5NgxVqg9Y0+LqSoeKxlCN5h6fcB23RCXH+CmuwDUD2Kw4
wAzRnw+R0nFe2OVZIb6+RYPJONA9Zdm2JmHThLWcTU/b9OCBabQqkaKjHrc7mMAG
eK8EK+NorYgk8F7tYDVKo1KS/U1GrNgH6U3EYA6jBQl9DqleHBSwR0NU5DyQ2WzX
zq+E4EeTocNFRivHFkcC5eZVVrEQyyPmRB+jeZ2L4nnwDLqOcPQsHTiSVnwFgZq/
g/DA6BM6b/AK+DcOErgEsIaY3zInVRamAkNS6g7d6CYgXux77/3/WU9GGkH0pTl7
DfkQMV4v6rr27YMAJzzenPlNgTXW152a7XnSz2qSdEF1/ztXNpOKR3QXXkLq395P
iJuF+2OsihWcimstqnisD7VjAOnaEl9ABq8kTgcbN+BpDYG7GZaJrw2PDN+8uBYO
ZBVlWiLLQZmXOT/QB7cmr2zjyTZ5dnx8up8Hk+BfP65nDW2w2QBQUf0blcAk8rvA
m3GM25wPSTB72i6h4uyfC9BCsC3eIaGADT/CyifZ7pBxJOVmi1ixNlGCXF2TCevG
CQM+mD9WYs33zpfS112sOFWQ/+LZnel07EmOzO75E4dHcK0FCfgj66ZTIHumiws4
1QqwVu8Le811dkYBDi1j3O3uZdZ2BuM2iMgqK03rCh4RfcsYdcWBhBAOKTaQ8E7x
lnGgOEzc+572WPa1Bsw0FRAfne4fVAhea0DNebN2XdZWocRBJngWQLd4sK0DLeo7
Hy6vemr3MGozHqGBhMCol+wIcRxLVQHOn9n0QAAKuqToNOhT9PfrmTycUA8fFjhc
1CMXHtohJeeZZ0kArShiRipFBGn2Cm+4bj9+2eQsEEcy3Nej9rbrZlPd+R7NcxVW
Fa8vh0vcxVTL2M+UGLBI6JEtmI7nWvnbsrdCsrL2q/5Uhj9CshRHsBw0gYTNh0hj
OAEi+CdK/eDGqTKIgs0DmhnluiIjOPtDGqL6zwRjrPNqOQ/fyDf11bYzaqZkKUJl
q9mi2otbhEe++vc/26zW9OZ65KEX+fEs+qrZANiaRAG+brBssVgJrSLaPwwtF/Z+
+/31xrOZRjNYcrba3xZzVSqq9q2fb4Mt3JQfvlbDzzgLqmquP5OXiRg11lXvFciz
hJGrB6+mNaCWFbxlq8z+6TQoGJdrtjw3ALGMd9LQFXLS/pawD4ohS+RhAxmcF03P
UHNRJ7E/l+vgAKHQsRHB5F25mZbi2E2fEC2RkM0BUnmLBEfJg83rzzmIoSqOSoBV
Gx7eajuVgzsTs0rP4IhtN5nwO9DlH145O3VC1CH3atR7LNtpciDIJoL3sWUYdUaQ
oIe9Deypq8uZhagD8EPAVbdMtj2X8002Ajvvi9K62nym2GtKPO4EnRgPXRCl0bFx
HrWrZAnV9qomktp3LxmxGo76q4uQ31SBh6MmFy4mJQHBZvfsCejfZK+2PsanGWG6
e7ZwHGWx2vXae8LlChVDXCOUqzAfpS+RfIQrKpu4acfYuem/Jb8j5xl3DMUqqXZf
UXcd5/Nm2dTmotkLVumZKo+pN2mWYPGA/ocVX7QV2JufFRdWPGf4HOJR341d96aQ
opzuVP71WZdzpxUFm/qziGbzHyLi7jBrqX+HxeDIF7DNg9wl0sg4anJXaYtHp4+V
0QPsEPOSSrgrhDCJHyFQnblM1LDKqzTIeiUTcqILkr89b/qiofjlfVWmFUWXbY98
Xp5teS7t7X7oTG7RrjZ0m5R+s4UzRXhyEFKrRSM/ZzEzdHnaEz2DCHz+xKjlg/ht
opKyzLQyBZuhPY22dUVPuUuikETTXL4MPzOfDy2GvfBuzHSKKCR927HKZST587sy
MG3IqB6bowOeoTfyz/fQQhy8f9CUKO+9N1OMvFddzuRtqdxC/bVeS7goK6wekaAR
XoyhFmnb3Lv/sq5dOV+B3vY5czEP24/KIKZQfU/g1xlTkIjfPFIyxju9sULuW3Do
spqqpWzst17SYzxOQEK/lqS2/G64ecLJZbEbf4DfOQPPsmr3X9FZ4ydHRwAMpqF3
n747h7fkLNDz9f3HK1OnBZRYePs60Y2otSNLNWhNV7QkhINKZM2e25tTuZGDruQw
SEMs0YGNCkD0s7V7w5QGCDr3vocACc5/VeXch3gadJVO9hWBLL/U6nctNpMCHRUV
DouyF/tphrNad1MHVVY8xXwFfmFuC7Rsu9Z9YqAFwg0VOhtKx1Vy+2OCSpkVSmto
gnD4ZAGJGRj1AXPjTYpKrHoFSwedJovK9LF6NQy7Mtv/jaaiy2qC1Lx5tCyQRsSl
Y2a5uV0C9hrMXY9u/fxU44sjQp831Est+H5OGoVKv2Z0GfY9rI4cVOzgwA56tU4s
Qld8x8IAVvHQfzxm5L/2V/u/6Am1kwd8skL0/glsVW/bhXgZYROG/4+UPEZOQMZA
03sYEjcm/luaSP3QJhhKUTHI3gIeT3mi3sgNZ50eR8UR67AGBfn3eDgh+f92Tx6b
sSmUg50WKjcCLS4tmJLeS/VsTJzvDj5oK0yOTh/FTBQVMqwV5sqTy6wmuX1A4jmY
dq6PycP0dbv6R3j2c+xWtN1mox4VK2iMaKy95trqaYBzUCDlNJfRopnk/xJlFOpF
bZctzMfm8BLG/THZYWo5pvJJM7+Zropx5WP8Ihu4YuJunm7qs1v1Tih2TTfd6KRp
DRT+xQmtOZMk0nhdfCHF14Htiof64U8wNE04epeBV3nWKAqlG2Et2ZZnQdpA9T25
IDI2shQB0+WA1dsYyfJWAvspsLm0Ha3sK2gw05Qs6KB5ui9y4gq8p6xKP1ideJ89
//R53JMCTr1Og4ZE0lU8ccBSIamj2jj+xQkpiMnMvGhexlGxz5G+cMHNWaMBbAo0
eI9udzOES51AmjA1XLMffbPI5ODa7Ksl68YUXaXho/Z4OWxpO8egY+OfpsB7LEKN
M4SQJbYZhZBiFUj6krUca2E1TsBFaOqwEBJrm+F9XvJjpHMsu1xBysnJvGOYTODh
yt+h6UoLGIDJ/MUgK/gSKFnosXSh1cY+/CGi1iEhRnoTy/B4wYHlKJ2IsCDa5wJF
Bf9eQw8qNTzSO8a9lgwVJXH2PWjcGuuaPUFlxG8vxRy1VsLvci3aGPoqOh5x3QGR
N6uPItNAoI/rL4dsQQvxN05hGiiSl76dvws5rn3fSFQ2yPzDKTj/BjFziJ+wqVd+
O5TzjZ0TjpC72xGl83DnMWXmlP7MJp5s60Okn8HInoqDg3CnJUs+NYX+2AmGifqB
0gvKjI/4Z3jOb4ECWtbJM8jNcRsZfoIlc3JvNRGa2hMCfr2x2lZpRpnjQD5AixqL
O6qJgO6qOiazaaXlwgZ6aitM9jpKkJquw2om+lzl0apcJ9eMPMWfO2MMfEmLXdC2
iEMlEwMfM1tA69iqm2qGXoX8nlNO+Sylv8NDsjuuL3XL+sFZa+804hJzkpqgNYGx
j9ym64ozbxRxthcpxao/+XQiriUvFV+1aGYQ5vSekQsf9WiOFSD4WrKjjfcKef73
4NzI9N882vz0Kl6L77oAmWbpGgaDJGMQrySNQlB1UbDBznvjwT86n6xIDQcHyxoU
PBFcT2s4s7Qa3uvi+Fi03IxP7sdj6hqPgXjMs3rk0hvOxwTD/9HXR2BvQZNBk/Go
VEuCfbciRRhMy0uHF6zne9q/6e2xCWfWqSyH1/fa75MfqEPI1aBOQV8w8KhxUp5t
XiVRF7auivveYuznxHqCAsVnB4FlJ3PBRm2LbkHPzpXQwtWxLtw5QQ8k0/PkldU0
YeGv/NPPqAeGbTCBxNPOwFhtBz/gs9fqC3wsws+gZmAbkO1c11T30Qz4jeyC+/Hy
GXo2aeOREIUp4tRALHItq+zEsbHvnxS1RPICI4XNC4MSKfRGJNsCBQ2716CSmLrL
+5koUlhuDlNX46h665cAkVtrfbR+6SfYYZc5VZMybTjI0iMGSmBpAVgjXWo/nIwM
89VwebueAwBQk0iZFErAKcaL4Ul+Piv/KBMEwkLsDFLiHKiT8VLjqTZA2EzZAuZG
PEbqCAWTitwNXDfG1sfaB9JgN1D1TcXTyLQWHErcS2YTPpZP+uKyH9YECCosnD7d
CudXA0HHyxi4Ev1lEPFAIXcJXueN85qnlqWsbCAhNl8DthWockyump/aCqCgADlt
Ko4oMRT/WYB5BU4lhzXfEirBLe2+dEz9V3ujPEM97drqcwM24Fa3OAiTUe4sdXlW
xQ3RkeTZtlP65JhrhwGunuywVa9Fvsj4hO1K/+0Zuhw9aEEx1JXLIST4X/d7FmcX
muBNzqZ7wY/c+6nvK9XzSsmiS7dlfo3WOi6xaZTyql0mBnolZ4zaVOuX0siwIKPL
+XMvCUP+QieV4ABzOgZ2xg4HPbHNRcP8V7nmCIQ5BNYZLtLj5I7+qpsR63fyrC84
`protect END_PROTECTED
