`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gUfRfzEPNB95DWdj4oWnJi5i+lGseFzTXqMv5w5IKPOaaBYvY/9IiEFOqelKzS52
NOr01Fyo0Qo9Z+nYpbW30n+9cRiyaaNuouiiBdpy8QO8XsAEtNv0/PEwiNI6jnh+
HMXj40pIFZXJRnqMR/1GP2MfjODLVqBZHybQmqUGsWkXLLpdP9YUoMHcmpxK74AQ
lexg1+m50xw7rCtO+ik37Y4vAlZNQJhm2q0/hGzu24FggIvZYLWVmRaqeQtkaWhk
tS0B7nCPns89oT93JIIfQ9aIGlKhkOP7bNncFYD2QCoTDZgEgwzJDyuwFAlql0s0
yUB7KowLzTgu9sQt0YD53bpjILOM0EeVT30BAdeaH0EZ/td24xp0rXj2gDdk53TV
62qxQuuoCdQNeLnXNRonpvW9qoehaGEngtD9kn5yTy8QGTrM5RqDE4R+BAO1HNS9
HvOYicpC0ZtXe1D6oKC1h7xkZc0dunsgRmLJaWmQEJOxSNUoWhwbUOmMtUob3n/F
GlUWPyfJlOLw0KYxVMC0p9bpZ/noJx0/Y3sAfoq/l7sK2uHFSR8ILGZpwGdVZZYa
tDF+jis3hUdYFzM3CfTdXQStjf8700jhvNVLIh0BxujI/LSrKyy54A1Q6qsNg+qi
8qEPnRnp3xN0rRwe8Qk9davKK9JQR1OMQhdPx61KmxjSGePwfnnR9qI4rKJ1ASdI
oyLzTOxVlZRkI4evxGb/fB8UnI2fr7mfrp4MsMYq/WUS89j0mCVZs2iOMEUT/Yr+
`protect END_PROTECTED
