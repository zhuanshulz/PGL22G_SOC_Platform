`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pSTIPOY8unSBrQj8OFgLyEqjqTtBAUcv49kWVjFUtlzfnYkVEXe/MlVicXRwTgyh
hJvxwXo2a+DrM+iRvKjUChHK5Lg4dBBQKPLY5ykPasvcS0ezrm78Vul+ayoII0Lm
vlhWRGjqnx3dC+dUQI3d4owpqKwiK2sk92qLAlNSTImqTpBGOP0W8fFCgVqa4asw
ohy6Jd4qs5nYPIpuiYJB+TcnsbLzO10pVPXteGXk1iMhamgOVTcWq8nGdyu6at0L
mrP4xf7N4fxN1tVrHbRDrIhMAKi6nnELu9GQbvKEUxQozvyIQsKnSoHHJGlYMC0d
X+0LYGe3U0/hGzviG6oeSPTP7F4MxeYAVuytUC/gZF6W+wyYO0yiF6lFXIoyZtnT
NP8uhveTNXNQbomDcTaviwAjcBqlEj5M4/Q26KWEA6Aphz6/qsxfS4adgpGCkXpV
ulqe1C6+GP0cLwpD9sTCyVBsstHY4xmdEqPJ1OtVmV3voMs+Kbz7OynHlXLup/PD
v80H72rqQ9C3CXXss4e408Qm4HHXLkOHocK/Eem/JfIyEBZsN5vLLpH59sxGsCVl
KiWurhqAtNOwhjJNTNgFLBH9DF9J1rACGDhIsGDQsvyUrBCZJBcUitkCyJizkFxY
CPOlqreNqtAqWz8lhI6Di3wTy+vK0GtO7jGnOU65JJlIeWXxMSRnANL+DMCSP6lE
qeAPJmadJ93KhcBVJaG67sozrlaermTWlDA1gxrCjz0Ggd+CC2UMRMf7Y+fqGB9J
7wJEg/ZYR48yDXPGsYlj6daDlbR59SdzYLwmphw7JnwrD0GQzofeQxrO+j83ff+q
JTD6H4Zkqr8u+JLX5PgaRa7ZvmBDmmmNkLRk729thLJs1u6ctJzbmdlo7ZMtwjZ6
Kxt8176EUHDpsKjU5dk2iAQFD7+cyBNphoLBV3I2JbrVSQc4vC5Ag2KfB4cwcjNW
BNiP0tA+A4iJC2AmxRFAmugN3bl9vyNTmhoeDDq67NmmuWtHvGawmUUw5Bg+YcEE
/sHim5bQ6tXAhVVj27BzVcuB4A0e44DJbtP9u6crbBuNvOEo+i4iXKuNE6C7RzO8
`protect END_PROTECTED
