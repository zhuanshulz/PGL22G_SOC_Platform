`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tDDcNIQ1B6K48xVb7gLKUMK0wJGVq889A8j/G6iHK3jsAcoScU5DLes8YLB3yv4N
wmiBtTiVvLSda8BC4ErrjVduQ/DLjOo62ub2v1Z4jFKCokQAR7VYkRO2a5BUcrrg
X4dx9kNJUV30zdqE5maA9sh2CXipkBBmg8KYQu2GV+IxGFLyYWBjtPfNJ7BfhQ2F
wwempKmmiCnVQ7CXsDbPcmSUEZ44kydJY/qiNtcF9E9+fXgcX9/7qN2qtkh6PSwv
FfsjxOKRO5LRSQrFzB4aQmRbkZ0t1/UEBIl0t95eIvEpg9ZqZWTHkUfelySreIEL
TtXZXRQ2VeOK9GgNUUz8Pyy+Q0bxGJrRADdKfSo/HZ4ziPjSyM7mZlt9K3xhr++e
QuNADS+MxSrF38F8yxzFMOAcu157gnAUi2atUt//LjBQQe5g+eYmJbY0nGRwPj6l
6735wDUpFTZjAz2E/wpPCIwyWZOoW6N0Hgv2TN9K2yTeH8M+lDQbXknm1GixdR4v
cpxCpdL3tark1qwsQLFkQKntlm6cROFBi39GaojAvlARNyOJOHZF9SeMK6sJdUj6
8uPK8n2i90IasDCmqcOYs6x53KzG/u0Tsd9UTg/2wt2MBCM9YDLmBtD3sMlPoM7W
V1Kp/U0i5EKRc5Or4Hin14jFEeZDD25jGiG4aqObCN8UwtRPyjfqwwvser5uHOS9
Run4fSs+IshOKTB9zGWRUoGCYtGM+Y73e5sXu3q0KyxOvu7MLszza3adPVSF9hCV
Plb3S2c1CFK8uM3bS4/esHuQ1XimQ5begPD5FxLPcvqUfEl7Ry1EzRtBOgGoaAj4
buW3dJN+coBRxMvjpZRPPahQZ46MCCfuDDWjuN6YcUMs4scYk4l2sPQc9p4lfbCM
IHmmRQBmwjE8JrcROwQgC7HhydhKI40WEL8K7E/Ng7FO5j4oVIazGoqO8ranG/kg
F3PSogtin6+CSLNeToy122v0AdLM1W7vTbg6rvzMrJX22ky12LCHAiRROS+9f1L1
cK4a6UHXqHJY/AjFEb6xck0GPDTKlRqmM7/7E0Vw6rm41rVf37hHECEVFsfAzGjS
HKAnuUVg9EXOqJfX2ESKuqG1pTEoXuH6jicfZEpvAvjg+rR87FN8LQSgNRaEe4u5
5xU5KQOBapBGGSJgc9AVFA/J9TPkzvtthg4q6K/qE8C7Ju11cHv1BvZxvqHtRtRa
HlOoobWsKpLa3zf30zuum+Ti7GkfJ5wp19kiGWTCJhY9XvgUZ1QgAE+vfCOEcN70
p4uAc1BzO3IhlPKFeMGWS9sJZ2fKYYIf4kwFNFzv/s1IgieeXN+DqxhYHOnZMC7e
JXjoX+vmRRjtDAW7IJKx5NZycB7I1BOoovlbElXIXiBxRx7pD2jl1het998NHDuu
yMgUT3CrQic7g8dk/KATluBuwYCogAg6EzalJpMQcW/gRwtj8jKn9aYJ2FMJeVsL
uhfsimGaLFyCaKJOu7kC51GdHRXlnLTg2vcZb1UmzM/9RWpdQhxRA3pYqjUu+ju7
bFVwxedCTRKvGk92oi8dAsUz4q54Fgx+JtkTvHUBHPtZkLz7zjYBIN8cWzSy3EVx
FGOXMgroiGkEcXysG+rfX/08dHzC/burEw0t8n5qw8X/GuO5WoQkKe0vUl/PTWdP
jBQk+fdGAU63tbd8jmXC7TOQ7OoIIt/qAERMSlIVUHuMMfGq5nm5CYgu+Siy/4y7
oEvpZFGEZpPLzWL8WMvEwsscf5LivyuiyZNskpgzo8QmNZqaN5iBLZU3tb4iX8SQ
3PhCMlc581PVRG48Okeq4E3DVxeijUEV6bHt+X5ufJX8kfEW87LVc35EmslGHiOP
qvT5T/33nut8qQMGtteeRqcxT5RKoveW59TdhUR0dlR53qTLvaS84xOcNkmAWbBf
O3il48YBQC4qfQAKZ6HA/CuXCcq/j6wkPdJENGWQhC4XTeIW5JyzCFX7JCr9IYym
ujr1HCb3ynk0vhedC4Wcdk5VM53thA7EW5bGm3t8yXdqOBnT52hTcPnqTIecbSZ7
nFJdEfi0DNiII0GuqTRf5fZSizggESg06tp864BjQLM/Snau0I15OvgFDNjeoULo
fLavkjuGgn5Eg+3DU1mPpiSNL0hWCi0IgiiRZhEZ4H5ZaKngYvKU+CTqL0rz2jVT
l1LPuIoeWb4ahJBJELp84Q==
`protect END_PROTECTED
