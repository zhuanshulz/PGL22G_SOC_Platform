`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LFkXYTRAnmu258bBkneqQ131rkuUcJTgwdZCVjCnH7bLtYm7jCC9fQcLXzOx/pJo
RtKJRD5/Y7WbzkARbOTraqNWZ+xD8siDbXiPXJYaVH+hj3IepIOACB5oYlwwnJrO
xMtDArlrPNcagqTUWUyzor5qqheJUqbBbJ73f6BZoIXak58l85PYRn26rBg1NvAB
KYqH1sRqwwhkmF1oSdKvl0irpULEgvuZH/M/YZy+jYaJM1ep+ekqffbRCW/R/EY+
xqNSr0d+pRpYKJqOckbYSAuPDzr3/EXw1BWZ4ydidbZrMaaJK9QoIMrTBbLoIn7k
8TaVpfXxDAx9ZSssUvYcSacNGiK8xFggcCpD8CNeTfM5uS0myuPLDRJ5IeAIwbyw
VbUrhrDfil2ERVCg7EVd90E3r9KDy3R6tNLL6gvwKQ2GT6YhGMkIsAUESW3Vp6VD
/V353Rr75Z7Qtkmxql0DknJ8BOghDlh2QOec7s6cNavagqkbAs8QcqlDZsGJwsIC
tcSrJk05ERiu3K9tlAg/R6LusHUeL5F+GPsGraciIA8pyb5qvZsr2SEnklnlr085
poBBygVGK4KkngnBhg0xysX4DbGAaljCP9guWoJn/Ux1f/ljO1SmB0B/JnKx8iK0
5ZTEgkNZLfzLcoB09G+9kL1B5Eg3liwpBAvErHb1rKuD8/DQTDOeCkumi0LNJdDb
ZYlbqxCeZPyF6yDaUTeYY0lLmRFEBSAQ7Be7/RMhtjwjLOROdiVAMZQ/wZYDsKEX
rpC6v4GNEwXJeASDM6ON3XRcsaAzAJs2tK8U4fiI13yPN1z6H0xBAziKwEAyQhmk
zrJSZ9ph01JQwJ+Z6PaDC4QkISKsPXRu7xcbwd00F2IXKA19WVWpz4QKmaJrsu1H
ineiwA+UMMYq/8CrGdiunMVEII1AU/Z6CQfRH5nQj7C0QcKincyHg8tyGCULxdxp
kALOax3O+qPMOUPyANVUeS48XVtksYFkEY7WMX0esnG5Rs5Yix8r3oQskIskUxzl
S2Ytc3Z9AHS/6IiIt4viijgluEryenlbBpAcYTx+E1qmRo03V41sXQRrOkv7DE3R
07r2Ie7Wn6pjM6AI/HIQgDG3yXgWNbmkGbZbIHz5r3X5clYGgj29i8oTobO28TJF
lo0ZrkBiuAD3q2sbwQs8Xac9Kso1NsohD4XYOYuzOvSBBe5KZD2YsB8WDPa6fceD
jBnYFqxPyvAlwyWeQ62htHbTeSQ1tcz1SG1LgMlGJCbwXdtWWsVlJdRY4DLZjdn+
4/7aBt0nwkg+VSm6JaoN/hwb7Q2OKesivA9oRZaX1Xnw84dTa2SgujxHuQeuG4Ho
tFNniZrNJvN+ZR2Zad157qPIKO3jkCC7s1TNsIWIWMbt2zplhjIY92RajNnIqKwo
vE/6dDAz7qihvgtUHOUiwa/6lecSiohm8Wp6AiX18Cu1WtmGPDtsGbvQv8i1Nf/+
oNLttEx3JN7S6NKk/l2wX4vu3CC5tgMA+to3j53y1L2Qn6QznUhDVNNRoc4+0mBV
3APFpeBrG5Lx9K/xJ2PE3rCmNalro2HCrWmo09XpptU63w8N6yM7A+iu1PuV28gD
YGhWkKOAtQQkJ12AYNFsgVoVr8MQfe+BGI4f5be8k2bepu7NnC0JeIZ2TPp76lKo
5GxjCbHjZCTJeEJ+TVeBI6dCFhGOspiWwTmdtpV64yZNvTIGwRVn0lgDHa2sGeks
Exnnr3PUxSm+4jSX2EyowF+tezLJRpMlKOYnAGqPmV+MVm3FzbGBNN+9MARVvhqE
1xymbvytThpReITgx8WR+IWp6W0Ic/RjXLk+5E0Cr0k0Hpyj4tC5/YhWC3LY9rNj
EF8R1lrpo+H6586SxaG1A9brjj2+kqNtT05ENuP0mYiCKr4Th0sOTX2TCSi8VUzB
3A9qG3UwZnmnnVjl8T+4m/iw7PVtEAdq+gQyK8ThpO0mrZs7QYKiSpK2ai+3MS8M
4BwAKXOHBSYyij//PWg4vUXKYAnLUF+kX8PWfiDWIQTGeul8BgagzNdQLYmNZfcJ
d2Tcf9LWjgRhn8laIaMLa/grlXnnny1J9l4aFT0r9tQdC3lL3Trp2YVB2B9xYgdu
vryaiYqlYow51vxte+ucUQZMQhrhprOjYXsCgUmExd9KOXzcFMlZR724Jq/DpFAH
xMKGqCycnkBoVwr7Ph6s70xkFtFtQuPVsiXfcEXzv+ivRjXYxO6yE6AyqxQcOSAs
+m2nlKYSbQPDPD+624+jsqbEg8QruBGBn1fpUmGX6qeitqFE9TegtsSTaNbM1Z8F
njxTo8cn0f7TO0Ng/065yp7KugCDEnKSPDK1xvzJxQH+Qyqf6CdF8xxhqCHcl5yF
j5Z782D/iITsusm1fPqR16tD3DosLYOB3LMzOMscUpckUFfAFiPmQbX9oDp8nrxl
AuyAOKxWHY5KkjocC+SlgcBXthvWhriS+Iuc9YD6WAflgF6wYxlJiWVoJ3+LG+By
pT5V8A6S4sKmYw45l5yd3QUskj4sWr3dtjY7hrzDFDFjNpBqTBEvMjw+KeRZItbm
xhXUps8IZRKdLVofVdM75da3OMCD1w3j0DoZTpzlBHfX4KYMMcbIJaR71bU3qL/t
lHAwiWsT5aorKckWAkcid0FhR1KC0Iu0wP8v9YOoYp7UIo45nWDnLVx2Go3JPMBh
YyEfS3VVYmiui8FthCl4btAS7LBUc3IUCgO/LsnOVPz5sUoqb+wQqi9vOh9vZmbP
jjopbW8uu6YJgIekd9tmtki9ED2s3e47MGTgOcHPSrq6K1JUzfugnca6hkJVY5d5
qshuyoGookXZwc+DUcOPVvriTtJQIf3aK7iSGBQg0/9TuwxwzWzb+gfy5f+JAzpO
9YXdULx1MG7WQ5mtfAoJhFVHawu+GJqWueIQ3iKlW1M19rshfNaB3KqhjTHbjjDw
XA2yiYrxLBzfvQPHtKVhJVFMkYIa1rMddwrD50H/tsDXndfZJEeiIunsG3BQe7k3
llreKcDBfFiQ+8DGY/T8tj60IdrcI3Z2HdMCcevalcpcJuOpHJPg5JEmfOlpzS40
kpJ8G5FLZpPmG/no0t9/27bMtp4tCpjNtqBWGVEIMSdCpa6weBH1lE1cdd5v8S2D
0/ybpx54yunnPMLe+IGqWjXfNb5A+Y0pGKZgea5HHRCJe/dFD3jvhQPbhcKNCF0U
riyTFz7/GgtMnAMsV1eZwr7bQgpK0VuF7A5PluL7FRnwoAU6qauTryI2gFAjrj7D
qKNkGSLMhlb6C1IA55F/h0yN77VENtI7jtOPaYrB6EVIgHTYNYGToAxPfh15Ssco
vI/R0fMKTGf2dp72zioRReLuLHGlvvu3OAzPZuw/pD/cgIfhtECvbLVtvWEED82i
ho+QDxp4Dx1U+Z9noClVZ83A0mCpjIwiBFA5uQQt/SZ8s8Bfl5KITRTwna/jqBQB
220xCis+8QCogRRdZjUXOnhQrHWQnE25hH91NAsny/5122S8bd6CAbjvsPlTt4vy
RR2TzLc5B6LCwRIYkHL0GUL/iDvBJSBWGlpXYsPxEONXIxKDTFBRtOxZ+MikU31s
+il7vpnPQBx7XQV5QTq8ibr2zcjx4bKU1wcgKWfpYyYYPakbDoh4k6bb/1v1TJmw
8f9jh88Hx802INV0DyOPcJCXDu7vbVBjGs0YmIwX9kzLrpHJ5rmA4QpYb5xqxEdA
wQMP0MmuVgbbGN2dPSSxTh0XCBRrXmqwfWqC159gdhHrV+LWBPm2W6bW22ESpb8o
n0FTichu34BHSWftWFoReUDTKTX/U/eOhYOlTWK23WCAzwHDWpfA49hTGkv4T+j9
Q6HP/Zkye21QnttIyXRs7gjhL7jpeec5OQ6oi7N39LaQ0g03POqRHaFn3sAvfWYM
pRwUMmaRDfe12sohOuywrpbQ7TIYNz/AQsGDT1Z4DD7ZL+rovOA8YIQ2Q9BpVLJO
2+gPegTmBXQAt6Gp/WKUjcFMikODS5hAkb55I2IADTfq/yadGOTaD/xV5xKD9yA/
QvKfUH7so1Gl9vOFFK5r+z6+djAHghmDCPa6IYV4YEK7PV0CxNuwvG3YTovIDmSG
bB//ICPyPcq/Sth+E4t84GeuY1//PQ3KBm03VKPpGpo3+7PTTIpnbbsdYgG+yOXx
RJTuD+Lk7MOEZDpXWAR2+qjEtC907McfKnDTw5c2VqOqAamItTYz/2FFM1FNcENu
ux/0Bs5wGQ/Y4sRw2wvYRGl9RkpegkjByLxDiBlulAm2Ko4FQOb+tsSLXT2e9yjs
1DSR31+9NXCObjedsOHMv2gh4CqtON6PWzEb6bbfntEYGW5uTg/q/m3kqMDa2R/7
CfUsqEanz9515JgLnksXn1/oyy2Z3+BJC0W01W4WJ4lmFg6qCy0yDE0IwfMStg8e
1xd3x9PVdzIx93x7aS52Fvb/YKmwStBo2Z1IP9ECxdSg35NhGe3rqE42JVMOW1XX
w+iIwoArIOI8v2WOlxbyYQ7UXAmcdy8GnZngHRgA0kN8VzgvFZd/oL1wir2+5yqS
rYfOl2PAhtqXeyz+HlMjmASv+axJx3QGNZgMgJIkzgH33muorCifa8tmlCxjt8EP
Du4dgqg4NNQyuFgpBunnMJTqvrNnTayF1zDolVl0fFpcbfX9Kb33rCgUM15TRPqD
8OQ+WOl/10LeYqEEe7atqYhXIeYC7RdGQOCDDqNi7AgmHw1XUuXhRYIltcuYMS5z
7sknRcOsPo4vfNkj07bOAqyGOyGbahY6+CjEf+WQ+UEqTyyKJlKPfqhPXZjzVouO
lg4XYQDpz13UmNaodiwEppI3dffHNwY9IH3B0T21y8IDWdTKD+iakJdBAjSGknz3
Au6rrD3q1Zwh8xZr3pDLFh4Emk7VqSIkhOtY616kliJg6+DFsgoWIkOxJl97+pxX
IgDkNlbXDaeahpinNN0DTdgJPmen2RqDyruGrWVRn1MQVaZtRyfDzdXec7SyY/ez
WaWsTJwGOK1rQ2zqQaT+DpVOgs8zonaCiY2tVEI1rVgLazRhTawAlcNpOEwSaHgw
m11nBQxEwqHsi11Pk4lA3g3FTlGFL4JovRh7x9QZ/+OzuixPr/YL+IIi+3HFmhyN
bD4davSjm1p4EtBhBg0oPK8RNrCRxXAHIyRffZs312wgYm8YhoAeCb+pYjfdVBw3
GLLI4yxEqWN25zXGMcuYFiumQ7nUxNyYVkCZyF2cCQ9ORYeZkoJmc3do6z/AV7C5
GXRUif1j5hKuAQG/5Si1QPJJYGz693uzR66Xd13BGjwzsAd2paIbVihcavW4qHzu
RkeSrUSlvZFDOpjo0q9adxEUr7kCXGEmX1p3f3lEC0KXUq9KM8nABqKGvTsiJdEb
ok1Z1pzpD0uycpBjLMBsZWhc/M3L2mkT9EmNLPQrJ9N8gpAFVHq/3xxFSAYCgkg4
JMpOXXBjanNbQasOgESgmB9YRC9q0XN2KDg2g7l2jwZvDVWfkhvJ0iBM0jKsuJYU
iy7mr/qTPxxdV/1opLvc33q/zVx5P7N60XXa0pngc5z7w67sYfXhSmlo7S5oV70f
TD3RdQR02+yh7EEzAFdPq2UeX7feG6X7+JPcpYQ+r0KGdGTNuti8Xer9SJODq6VH
uCISdL0CUBlERbIQnZLUmUyvlT8uUrWA7ht2twheMhnmd45QBvwglMlXM5iqIm/4
CoUf0tjL1vNMKJ/FFgXjWL+mVQ87MmjbkoL8Cvd9na8aNAGx/LEj2rU9zk7lSgno
ETH3IxKolROoN6A/yd05++w9kxxqtbKLkt27lavMqGxi1kZLjSBp48jTF5Tia/QD
4f69ROHYyhTZXe2lO7XvEqk1rubWp6auJZLAZSKqboDn67Sat6ABAsVSTa6Rn4cG
XPUNivQGr8sgxsaMQ7rUXJo1VPmLyTJCoDNzBPVr/WuBrahlEgd9iOEX3UshyZ1D
Vb6SEnJnKEMCGY7xn1S8spKt0u2SaaQ2XzZN0N88246wEUil69qW+hDcz0U+OwxM
QQdWh4ODzMDhrtLhUIIwBU2QafBqf0CPSHqQLuW/y4rgJY3zVRJNNzVU6MGkiVaC
nctiDQwZHgX3rY9tbiasJuUMUu4vSJ8V9D08sxkgkJXVzraCO/VLqRoKaB3XPL17
SxsnfRg7P3Qnd1ydglHENlkcXxMpVYsbn14Fye1nLyo0OtzGyVHU33NzfP0e1OYH
8hTgWcCziZS8Rg/Oh3nqBe19QE7+BD7TLfFccOAZoW8TkktkdyYRfxtILSq6z/0B
8nLCCJO6jPZESbS6cLzE53T49c9g426iXR41Lg0LQJ6yXwpXvScooqCAAJvmJ9ms
d0bRsf7pF2CD+wBRvKe2i60Evo8PF2ymebh5SS3GGyQAhREUImIv3maePWcevYgA
cCuFFJOMB208kzIoTvuqnDUO9nJxjOiAEO/S5cEw5J+YHX/F6anlJIaLzvJaQa/M
yABHKcwZPJFGp7lDXP9iLzQQg09TYDzn541OX3onW4NZU+CPRUrO0L5kewK4mYui
G60og+ow6dZQsxPEJO6Tlc/6IP8a84ZhANjOZumWaSivMz2Wi1e605wzsHGCGQzy
nOUZFiMwF5vKeRZbqhsBArxqdSk2xRmYLC9MW7MMuREyIhK6DKrxX+B3in+V+ICX
ccwhzaO49V8tfrKhBQCAOlY/VuxAaj+h6Y9baGiLErtsCnzuV4TYXYhnzCdTtfYw
cOPCTZx/pYsrNeL9NJm/E5oY+C3mHuFhlblHiro+WaNkDvF6DG5CRvf5Z/vqdNQD
uWWihz0814YhxqV1Cf7HVi4WYljtk+LchepA3S7ujOcSV/yt0os64paupY5tndUr
a4NYFRtbzaxnTyJQV5d6WiL5YziGsxBovm56lqlGEH/I6TnPj1VVH8fpPXWQ1Rti
nxbHwgcvVF0gfmwqiFjPuh6NRakXGYXrSo+aDAl/sE0GCyjXqlkjndDhaQPzkhov
1o0x1nq6XzT/f7/4ele6lA/QynFjV5pA1rYSCu9GFZ3wKMYQHFZYGqmT6z+2V69g
cqqllMmaT1phZQL1iABY9s+wcIqSLjYo7WJpk4RWRWCXSNblr5DRUVsDUzJuyQUA
fsaZacZyHy/pnvZDm2zluNuZLNDcLTqQ16GWOG6XOUlld66k6bRmufp61AxZ72To
Wjn3vtZn+4v4TJoVi5XI9xR/OMdadhIpHQvK5ZgN/VIbJQjjGX1TY7ufK+r3sQEA
WP3PyxfOa3stq2Nj6AHXDS/vcskWGRzS/S3iAkLIooiLDOBDcwn4Wknodt9ugZEf
X5dkwEOI5YacCnlvBiOlCba1SUuwaa9+A3LKVLFUC2MYi8/Eyjfl6LvqUHcWqHlB
NAIHc0/d239JHGnwbAvUnNK2qOOjJ1y92DoOj7Pm7qRfmIVvnI71Ap6Zq/67redW
wTZZrPPJc6/+siEyL9oax62PgKgqFrgfGTRNwIjPfxgCQpubC40X+O9+k0BhGBtG
afBdelSMplSjYkhbS/8e4v/QS0iqqwdUoOH0//QJr3jVscmzDS+WWKKnOIi+FOOd
Q9BL/09cBLcyy8kLZbQw2GwucQcBkrFuVo2u5N8iOfqQFFk7WdHFdBlzShLdUUvz
3cNiQpryhGTk5AiYpwJAPitBEGH9+ByXMTd1hroTohy5wOey50rvAf7t4/PM0LjS
sQpGSZdZDvRVOjGEm+f6Uvln9wl6MpGcmeSSOK015hKDcnyV1ikElOPVPmUi+kpr
c4DCIA3T9/s/c48yzd4KikJwBBE4wskPsa5poHqB2TVW3t9xOH581wr20c6jNX21
Wa/VAndV0KCwIQMmwAF11UjmrNjkuUbfQGVmhUBuJJTUk09Fwx3BGXGYQHFLcYj4
+QegTHw3ojj9Yd8e34DlExglNZaUkUJsUuSnn02B88ApbEQWagieAV9UqPqLCTOo
2LxPv3TfKV1BYtRJURpRtaeUSMc9uWFPz4gxWnMWV3WJOMERBitrIJSIsXrUJJBv
h8F+6mDDfT7NknN0zTQC6HkM/tgUBbqMQtFLneqf2BIlLMiaNHjkUrm+maAH4oUs
JTEhS1o7uuHhcCmzVFA5G0gd0RuppuzCz9oB83fdAbft2VK19C9SjBpdwHi+3j+k
1saisyDS0pdl8NbFpp8CB1rCmObWjqXqPfW12fqhm7sHw4THS4OWqgIQdz4cCf5/
LArlPvC2MJtMbX98FygJLjlry6jae2+01nDTiFEyN87QttFfmu0JycoxMQCQ5f8m
c6tzLOerbF1W/C7SLErNp8i42XfWQFWQVLSLU81+Jo0Zbs+mJRS0gxtO6xxJ6GFC
53RCZO5Hux0EMJZGddDZA7YLEMe7JwFn7mZxvhT67jpwkpilsAEJCXNgzaj+FfzK
JwPHibLgfbRzkhADcm7aRYHCsuH9+Uc9ov6FXt88sokF3THSzpt6RF7f9+lnl6wJ
z/EiIYptsf3Mm32RSwGXnmowGd2yR22ii9Qyce4X2ECKW8NqdSmWgz1h4rZrIFtM
PJWOFdnYn0sgd1un7/1Ni2f3c2LGA+BBU6LCOC6cmfISB5mKMwYMYQboedfLsN1Y
g8T4aHjWtapuUamrJZHb15FFIzNr88WKOQR+LnzwEcoArS5IJd6GjlF6ocINWIjL
7HW6QJANPkz+B5aqIope8QGrEm2fqSy4mgWBo/DnPP57Wv83d1vrBTENrTdLlaD7
HxjbO2BRfKsivk2SVmzmlua4rB3JCoQvaQ9iledhcga4juVvxgpShl9Ijt/h1kBa
J/mLwSphLl0yHGlSHt5OzAirhvXJU8VPodG6MeSnJkAmqV87e1fWpfGlD09Xlh7f
6hppZ7T22Bj3+NeNuOgTnQ6EKOJhJhCBHmGr+Xpsl6G/DZAqlOYyHNYS0vhHKeZZ
JfRZllaf5GUv4RSeS9J+oJnEKn3iv8d31rMa/7OZDxsIVdf4WyCeyp6kNXl4Wsb7
mHk/wGg7iOLqFl8GGkqPSDc6FoJNk/hGQvL9f14mi3j6QPoO6i/1SSDtgeqQpBwA
nqjSw4M11fuGUIsaJFjcMrYc2qOMf0p/6PblcNzJFVoVcJ/DeClCF+6Gvgf8Lmmf
d9k9FXccAmwvS9xlVWDx+jk6DSa0FbOU8sQJx2+oWEM9uShN1EDkYKClUEq+lr+9
mr8Mik78aloEeuBs+h8jaT0tf9/17OBkJv2U3mj/rv8vHfSfe66VPJPFRmhxDfL0
/Hruii3SdDOlropkn6fcB4QzWsRO3FYx1O6KBlf/zzoy9NJmJNsB6OQ2mfU8KwU7
EvnYrAEcAZqPAWdVf9i8V/MmqX5YSppRJFes0ICPqgBGFSEQfTHi83QXMxIzihxb
rI3DD/ENOQ6/BsBruGNTQF11VVC7ym32K/Ct/1q3kt9UUrGfLoAJ7F+navgqu5rv
nzZAQ0PFfc4LyWJ3hWdsroeYj67gWkWrNkiiVf3RfEmrjE2Jn1LZH6fpBWyqePQg
QnwrQx3ug46jJxZoe41qu7A4vNplrLQK7jHcxaMAaYPq7ftQF8KVsPGwig6VUulx
78EiB9neGEGX3eLDAp7gs4ZSXAHpmCoQmn/zwphD+tYyvSFBAEm5d+/0S/Mrxlk/
bVzEo77un1MpJszMGlcyPi+72H/+UtMlLhDHJxE01bJ9JQtN/TxdP5mErDafJDcz
7ipXXknVwqVZAM91Jkm405hc0kVTZkHyevh1rt3eRPcbFXqJAQPYAZJu2oYo4PLY
bUc5exyspH6XGp28ut38ebqQ/bSeF/K90M2rrXEdE+OWM0odQefPXzHIYBYt+fEI
0X650Mr3aAyjHfpN3HMGQwXSNyyCIiRBh3lWNiw8bL3npHnnWglHHIsQY5l3Z66f
cYz9FiRLDya7F07NkmNa75ElXkQXPk5RphWhXSX+ZJycfTN+XIHbXVvp5yeBMEai
dVe8GBL0AqSlPHkj+9F8MQ8FvPzFJTYiquUmjUwxv7vybqEoTReWaeBQ8bQMJKko
5pU7Lq5+Oq2Dhr/RA2FKmlkNjIpPnQx06zBmof3XVlNGYNi9OePAVoFHOVlgj2q/
ZgnRK8fily0F4IZOYmKPlr6xyxRWMFHp6GVFHCertziP7TgV1ri6yL366PRvUw3T
AGkcCpOcp4WN8j4wdon3BAOIfNO7h7kY89/2DAJwTi7Mi76xFC9u8p2NhZkyq7pN
zVbr6IlwGADUTuVQdjdccKkWdKOwyzvaupMHi99kVIDRrT0Rtf49ZFYzq+rSr3BT
+Sm+RZ7lTr6jGblDftadQd078rlTmsCQO9OKzowJpZhjR2Jp+HxI1g3rv9qK2SpW
TW12ai6cnhFdonj7w9pknzYnsWrsXeJDGVRvAfgn8OaFkjdjTXfAy6k6RZ8fT+Ci
DLguHuABlqBmAdgtWq1O+obvphrzi7Fy4HrZcS5jkcuEDAKTxmuJYp8av039ppXI
5Nen6/syxGsHge+nXe5L6i4sEH+tPpyAWmqFKNFs6waoeAEntZEZfbaD8uo/vrb8
+XwAtQ4yyDm6WaWn+aOcS1y/RUh1W/iJSvMVR2UH0Z/w+znT7qUgbhPXtRy5Tljr
YdOsS/d1p+YRUZasDAcq5Ca026+5YcX8awuHb83UOCXj736W9MpE4Xpnk7O6eANv
fds0efL2dfC+/zl8OgxlnFUMjOP6ggSEc74OhN/MsH90pofZUaSH6lw/Yjr2YraW
8m5YIXoJKQzVEl+7S/2eLHDsCkp4enZJ1rOYbSQF/bIYsktmc6CnTF5FABqpVFD6
SLlQffHWIE/hYSsowULMlF5oqzGlk89KfGq9ch+tw8cBhWX3Wj3EIdN9CSVUEOdt
yUvPD6OvyeRg31t7jtV2jRq7DEoNtlGzvHNES4cuyCDOSeyWX8l5pLXgzBww8O9T
VwK+OCEAJLD+nSDMtDi/01rTC4nG3TEKR6fnLSQZjqs/6KBiAjexegql1M6Fxb0+
hNPQV2oKHoHuqUIHMCV5uWJTdlbBOIKOnKGKBETBalYB+exab/B47uNEG4TNC8Um
shUnGsIjGyUKDsgb8TX7Sx7i4hjG8SH3sxoRYhYSm4217FonKyxGqthPLlB1+ZSj
G3KtDPN9b1zYM3CA6NYHLJ1wDhwec9Mpx9U+rB+r1k+z1nm7A/qeaClTprD//EEA
OSNv+umMoZzAOIDIviFFv+AuyVTJ9D9Wdoc/v9OHBNPvjiWxduawXQQF+ohjbbpa
y51seQhCVeNq3XsTpdxhTJJSEQaApBzpyob1og0BurcFEtUJl5JtbRlnlVB0B7VZ
qGWigqWCOkvezzJErPala1ZpdvD6mFPIhoVrMsfjMdnST/QCFfXexLrJ2qnOHwvH
hcNUmsTcT8mwK6bmC4fu1afYVAatswkxNSbaoc8NRcUKisR5JYRhyua/7yjsKHRN
fattOhFR7TrOofWti8es+z11DU4d2V3XrmFDbMlU1gm+z43POB2N4rq5eG8n2rCa
i7thvbAMqDjtY4RmyjUJnQ+TXkL5Ubq4yYyryrVZh9KGLl5q6+k92Zmgcd/Qy35w
EXAm3hDsb0INsddoAxJGprYKakuXi0zByqEc49+yJ7KCnq8vjA3YFiMx0TgXcuWB
GenfBxKQ/o6T8+mF4XuTyA4DcxqyzVCZuXUFWnrzjBCmJ6o6k77W/QMsdVkFJQ9u
O7qLUKJld4qW4Tq8gtDEfmWP8c3fBJBtNIYojxAe6udsuAmGYsb37vmGnJiXvwwl
NjXI71OEAW0Q3fTaXtL6CzBIEHsSOkTHeuID0Zg2SOwFYKhzwMW6Y7orB2VHd199
m/Qr+5INLeJ3lMGpi+iQ2g3khY2L/S9Cevhak1Vue7CQe8FMFb5+Q9KFasBmOtY/
aI4I0mQyCpfOTly9VoeF3lml1r0BYrswTjn0TnO678/55MFsWBhN1hYZVyUMy7q/
mzSJDojPJ0di04EAlHNz1AVJ+v7PpCV2/bfeUpooQUV9clvMe4DKPFfs+gNdyYAI
vkzfpOsvF0EQOTpbfdgHBSKymTNbYpVulkz2PQB3w47niKxtHE4sGzmWpZGFFRcJ
rRka6CmPxjmLpU8G0L2TFDq9cbRCyLsluUAgS+shA6yJAQLKCaGUbp+VBNyucflg
fzrfpeqi1XLWriAJaDK2NqvWdi/6soQN4cslkd3McejGcvqWmLPxIcApZre4NH44
+TpT5Qobyt2EGjA/ibgez47HaWekYRsrfpWoGvQLN28YZnt2hsWQ/07/EGxnqw1B
M6mT0vFW93e3edqDLKr3cYhGXpVBRFdEkjXGl60h8MXEi1hNPND3rrdRbKAhuf84
POR46Cz3UtQ3CYKiKD/lWNrKCh7n1fW9UeQirMY2oBdwecJYwm3+ec4dDgfTcwMF
v0yeT2N4WhwFwnbp8DwwblV1vQ5pjT35Ubx2c0ZWltyq7aDeZuomT4spxul+u6TK
UJj1zptM61J7b8x4Z/p5cW6/dKPiOMPtkTT8M6frT+1F2U9whrRa1ZVyr30wS114
WtnI8pQgeS1JE1fpE8pyHubPuYAg77WptRD4IE5YQGhXiry7rtagvfSi/c1ygfeA
cxwBdEJjwkUdWhkDraOrhsq0cNzaKg/ULuq2FYymdwsAeaaivwqum0FqeWzSw5iR
g7pyWwCyYODW7MP0wXEaeMv6jaNaRXp6KYAOhoQ3POlcIGyxI8L84OCsLaaPyOOM
OSzhhNPZSsYDUB0gmSZGnVdEFE1e6inJ407Ihy55bTILrVRiXjlGQ8FZ5jUTJVnA
LsQCnHWm2fwbjkMeFRswthWubMAwslZ8KI3HgS45klGLpPD4qyKOElKpD9UbtgU6
yJpwdipCKlxAUpidhwsrcDBnmo2r+22HqrJotD9fYbNh7xuRmScypG250kpkYYYY
OhPiikHgJEablRrMYsuXxUw7avSdoOhuWRul0Two6UfL93ktp4lNH5dXbBZ1y9bS
UjmvBrXl+p2zdWRhfwQPSzWT7qb2hc/sv9jPuCy6pFac2o92gLRAfeQLyG4H77CS
H4Idadb+uthZQsJ+VNkV9wrY+5ii4W6UDY4xpAKR8QNZX3Dpu1nP76EVWiEkhJcT
s9Kr0zi1aK5pd+TL3w4fVWhfTLBZC9dPayWARR59zOcBw0z2HMz1zC9Z7AnxelV3
QabhZHQims4em+cStfuD6/htIeZOnDDZvXw9sKF7wMsV5AIYnIFZ5TUcCTPLcId2
+eobqHIk1nSGY3x8c9p1ILuRqbp5eIdZ3lEPvWntB2QWfN2RzkQYyECtqICtVM24
vLOMK5F6b5nlTWHvxofzCiXvReZs0wS5eCFSRkrfiYgjF5ymkrp6V9pnB6lVcXop
1TsBg517MSgiqSNiDLS4nRMjgStU6ZP6tW5+SQzr6N5IATj5uxc6K0PNMDOnqQqo
yYNqcIXW8SO2NjFekX9CE8OdpbZmprqN8pd84H0bvNzz+PwMjOjNhFESIZ88NWyR
kgcTiZRuHln/ApIwqC2e8jFeDb/fCL/0HKzT3TQutC6PM/rDIlZM5TmfPs46EO5S
A8rZeIW2/YjrtRX5ghf/BAA8A5EYM1olOM6qgU2hG95Y1v8PW2J/C+qk2aXRcQg4
usJjapyrGN+9T86Na6sxu5IlV2624ksG9McoeTFEgFA303flxWUbib+gu9Rqd5z1
4ZEiy5/FkROIt1/uhOpcXVGMgUNjbaI/Rl6mDp02chAiP7HzHfsC8CmFJuh7W3eL
+I3/DZv+L5odMR9Jv0nbBX7Xp1vDO0sr0vHBWSck2hgrdx7kVaykOFM+kHMgBmuv
peBQAFLieQz5xPWGEv07OXJnN2EVH0spgo5QOYjM+Imy3Brg3YPujDKrv/qL7Dow
noeuuWaK0DV801rwWfQg6pvT2hX86QJKrjUhfh4hu99pZdznkLMMTLTmkvXvOL4d
79GcmvysvT98Qeka+npENYRL3XHrHvrZMa7lER7XFjfnpTdbpTPER4zp3+KD2M3T
lqLLdrO/Cyx3DE58Ybx3D1OvrwqwVtg/uJbwg+wYVPstGdc378sIVunJTUTEeXha
GiKdzqaPvTAckuGKsgG5Q3HZE9kgz+Bgeq8EAV0iLoU0MfVv4Qs9ggP5trNw/fgh
B0O278zzZ5wE3wfRAmsFt2QGrwa5ozulSSRtQcm0pQQ/9e2NS1yRMDPW9xF+2TWQ
L5kpst56ikqn+QJp6mF62RJohcUSdieklRqRf7pYmRhm21Vi7NmUzhyWAaT2Stv+
87oh3pJfi1LC/sSfTp/p6Q==
`protect END_PROTECTED
