`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ho60b3RoBLTKOnIVmR3Pk3US4a83k6bnF9H8kUt10pF4B4SS98t1JdUbXy9debRE
oX0Nt3X4opd0GPjBcBa6R8KSz7DjHZM6Ns/PumLML7YQ3dzu5hJOA4tuTlLTUPZu
AS4Of9WAc8ba6AcIXl9cAiJs8eNuWmjgIkXlNPROuACkyJDXxsIuuaekG/RqVIOj
Z12A3oE/RjSLLnhYV6qaf4BFS5OaOszVageyG3UcLp+xm5NG6SFcyAdfP2C1gyOn
buDyrnqEJnQptcAmqak10Q==
`protect END_PROTECTED
