`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6/VvFDdxyrH/HpW1AXEUaMIs3qtXePx/01LedIqrIvLcxlH3nuuh1M1hZRyHGSGE
oO9PIEF4ieDbNI3u7kTd1QxgFUq2c1Tp1oQ3lmWGTjypoC9I+255IGZvGAkKFa0f
jFHB5gi2bJ18SRdbsiBbL5kl+m/zoRT6qTJrsLFk7+lMPkDdK3t0WuUip08zo79X
g1FACGRgJJI1L0Fa64GL3at2OfY+EafMT7INPATrHxNBCaCYQiXqMzQLw47XY6Ut
g0MiJovDQtvHyb/bj1jB1JXvW+m3ZXCwvrAlj/HfPMfb6sD19VOPyYOS+inDNuEr
M6yP5ZyzOx4Bd/GljG/CN1uc0/SZuVtyX0hZr6gKHP2taVZXybZd5eM5UsTGe/iK
32Wq7lvhf6zBv9wbvJa1s5Z5fQ81XiT/MhBRBc+L0iM3dZbl84k8PD2otaPd4wkq
xwvuX5zDeIcE1H7b6pe45y1AOpHjU+BAOmaUEdE4DhYXitTrG29ZApjNtNl1agTj
PpLBYlJX8mbVVWZPH/guxC2Sl9GlfHPQ76l1o8ayzjJmn9OJhoN7NGRao1r1Qqws
oRkTBR64FfndnY8vyH9Qt0KJ7CTZLW3Mwdlqh0Hejx8QrU/RT15JVGOOd4LDeu8v
iJPzCsaM8dlj89fvY4lT2rIB6jkPzg9Qt3scVbCb4YF/a45NGLVsMa6efhMZxVVe
TkdNg1iFNyGiTCeuGmK5gLSW7Sh2e16fv4X8xtKPsPOveYyr7wD9QuRwF05CmEm/
NsUpQ5lkw2ZgeKAzRXLAx1RloyuWYeW1ulskkEWYdcAqo3abvUdyzLOg2fkhhHFO
mpF63CjD76qQ1QfDYBI/D1u0L4OuImclTwP+BaaDqxndTo0JRd91/4PipyFEHH6U
eUX+shlDUL0SQaXzwP+4LaDca8znSWePEFLacPx/NFp3AZIPNN0z7ni3h/DB43la
xH/OCZdpcfcuzMor08ys/wVV4L0YdMbtGkc9XtOiolS6UrWzLlLGB/zrmlyfOma8
1BvSMz3elIVA+qcED//tXtwvdBFxyJGf90ixR87JMn4=
`protect END_PROTECTED
