`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r3QUYawl7jHIS8n7/CbLzpqp6boqfZYoyzusHC1CKJO7S9Wxq4chRQPU2DZ+i21z
YOV5wE+yLnEyDG/qTpqh/gW94enIGfnxy/hqcyBoJu48pSYkVzmPyrkksdGt2QFz
66R5BEnX0grQQ2tBGR4EQxe0w+Pqx3/ep47tbPABIztoee9/x6RHTpkPaneOmH4l
YdcyttVECCwnt1b+7DK2kdM8UG9qlgVfFyJDaj1qIRkAtZBZWMOSK6EOurJj1HyR
BVde63wyG7OApGOLkSMYBB/ssL0ZA3NL6DQ6oDvJF14wvx1SOPhfKCIlTONeTNpC
U3WD3PV6gbUhn26niotypQLHEP0JFh9XJnHilupwpKxaKOa2uBsVwHXTN7yEZUVA
SrHp9x875oLJMh4PFzYmJpC4uDKfNpVKdYaTS/o7HDErsgQz8/mF6ahBYepdwbws
nniL8rIwfMdGntGkP4RbGYd7HpPt3NlcmLxAPF8IPssoTvU6W2Af0v2vYJHht84n
nI/s0pmV3RQWczaqidC43S50FtPRuT8kl61jQYHtsnt6YLMRshlkJ/D7QRbgsKBB
kK+JBb4xYcHV/QKdEQqrmzb1wE/LBJk7kIIMzDmsGTuPrz793s/TW24Tna3BiY5J
FH9BHt6QKYzS2JVMmFUeRO131mz3CL/THLzorSew9G4WWPmZpMRnW9VrbFKUpaTP
LZcJgIKT12wfRqDMUdq0/tlj6lcvnZxNzdZC1SkCEc2gK0GL5YVMzkOtG/8pH7Np
apLqe/kWmkeuyou219UUG5HFqi/v2cYB3/xSRljVtt8wkwcDf2dfpKKamdYWiY89
3rrdn34xtNGEnjvn/Swc6rtEfInBu1/T1S7Fgc0Z8mv7tvOkzLtQk/Z2/xV0mWTJ
98pjm1egGNKQt8a+al6Fn9v3ijHFsTNa4ZE3bDZwr8rjcKe+HdoEeg0T78eyYDsp
R8lLhM5LUIFLGXx0Z3fC80D4277M72BX2XG+LLC1FuopYuoZ/tbK1hdRC+AYewOp
piFvwx5bK47+EIKsVBJS1Y94UNs/HaBpnARIqm98DnBVvOZkyrdyFrTkYEFADtfo
oBVaVVAMxo/zvsNqNfB3i4JpFR9TN4dvm16dpj0aAhkv0aAdKGfFfhzaRJgGuSjQ
PmdrDgPqVqn4+QXDXLNuKXKRFmi16uiaILxfgTQ7KHgUh4pZJowBJ3l/TU+nWi+1
aGPGUV+KpP2hhm1054pPCv0VkdbGYn8Il0RhBl3OM6+11nACbysZHiZ6rC/+1fpd
lO9WSmXgu65Ct9h5Q265OPcrs0C/zm20vlB/Mhk67ngKtEG0L75YOnbIa0rQdcFU
t57UnmwMCWSpwCH9onLQ/wqigsijt5lZG6F/v54YAMkzV1F5lwD+8VV1UfeDhrCS
OCTUkXCWwOQUjOAgqrfcGLJbVC0MGrueQXxZNBU1hV5t2daA5n2GX5dIh4FlL85f
ZG0WhOO5VDGJZ4xIGEB+uURmQzixlTRlvsjKJaWnW5/wN/AUPWUBvsXfsLgq/zz/
BLX/KGXtaeGu/yo572PJlnnHgRjKZvg0LZAKLJSsFxcgRR58go7HsIolW4WBKh4v
HIh4TlLNLPQermZczIgLmIbZ9aDMEP4yVtMaIoFVcOWY/QwvNFM90zeRkrUJtztH
I4CQvGfkK2BdLL/Nj5hO20xkN+h+70zlcW56Vnq4U7YyXYauQmuLWcPaWJiQ4NqG
YzGYB1M0mZHjE1S+R7Y7LOsrMOde0STvn5BVQIjPxx6LMMI0DGrLE2SPZwkT4gCE
VR6dXKM4Ly1hyByEqr5N3OcFVrOLgr+CrIwwkKh+Xc9v+MP0Bp5PfVt41rstLnc/
Y8ETUsg3GDa/WKVJA8jVJCkmW4SHhaJv7ESvFqidvUzifDGQRxvCEiaZNY2YWlTW
SoL952HEKzUHfIAx18k6aNWak5uoU654qBisEleQ1k5YpQ8RGNM54A1qHNrQxh7D
dBnxLCu28IVZBcrII/N44aZt+WU4HJHrxewa2EevB0w4u7lcoWdfgWftaH3U+HLB
dO5PNPPRRsXIghIEtrQhLNQPChjBm4gMXt4hD7HmxLzKbp7va7rEjFphFvCRpSvK
PaZtCpYM85WsBeHQ/05xZIA2tKrqhRbt1yKpM8YN8JWwdsYKuqL1wEb+tQ180W+l
U1Z20EDd8xUvHXj7iQJrP4MDnbl4qeIlKJvQPafc4zfZjQ5EdPnXvlboO9fSOczC
rld7AZLW0AFS9r8nEN5wSf53dNa+8GDfv1u5R+qqGH1jocV3bjn+cAzGpVIHIVoQ
HF2Uov6CztWhaIlIBj6cH8ibl835WOW9B3hModVj8vtAhUDoemE+bNMrorYrvrE6
KFRCdZ6avgUKbMJ0mwDK5BgCF0EmvzO+Gtl3gw2xoMNQqqt0tPQmalXpzXeX/URu
0X44sjHcu3BdEOj/wbOgUmOKrnfZ/0DroLvQdDW5v2Kz0BixYxR+ouyw+YAUWJaX
yqsIVmgWyk7wVsfPPBLUw7BUd8Td/2A9xuUElCJ3VefL+eO1iAprqb2f41xTC62v
AfqAzHk0fqjIAGe/cx5FY6mQy0rQHKqIBwQOoB7hPOX5WaffEdJ0kAR/3jww+vox
1gYOkQ+e8XBZbZ8ECPO6PsjGOTI0Bcdi9kyAIa4FqHJQ1qOfMKjVmquFhj4vtrL7
OChDN+D7wrGFtaaNF6BlKPBjF2S255LrV913A/nuJPcuxlkn2BNTWvB+AKdspGO0
x+CL+swd+kFEd1sjIyXcQCO3bzln+71s2xUx8RZdjcNNI3PNgcryKznXn6JSSARI
tpbpsYLKh06Q0XNum0dLg6vZxLeZn/MpZArDVC8JYcDPhlxkuOurMtS6UkgQmN+C
lIfpiqfx92581sqOPJzvKBSYpyWkQaCAFZuQSNP8DakcIRI08et14OjXOZx/Wwg8
29JC8nNkKHXs07MhYXeFQESat+0qo0x7H5mgvbIVT3W9+nzEBrOY+wAMMlypXh7v
k5tZltisNpL1OsnpYcnb+gfdveYdFdEVHP8s3Sg5N2lNhqIA0pBOTQrKOgoaJevC
d7qd5JcWqkySBDeE6Vp5y+XeqGzBoEuOGiy7eq57W+V9wX/5HmO7iY+/cBIzKjSM
rQne+lZJaF2q9312uNhaeDEmiwHfXCFxLZO7RcpEoIjciGv1ftfng5p87+tevepq
9pqlrIjlc4boXsm2t0aCAz/ZE4EbE708KFJRdpRdjjDhkBIsMhratz0BTTrop47I
ryKfy4wu8vMHoPxVbJ7OlBPL+mVVXIP63JUWWfgBWi4YuVR4vr6PmO8UvZ5QZ+dO
n9vVkH8LV+l3+ouvBWKDjXbst/mxxytlBxq2/0HjKUseP5NoRTvcvGt/aelSTcmD
xbBW3HOOd39MVAJ56HRxFUHszncKowVUnf74IDFUZ3FsBv/6tCoUHvR32+klEsNf
pQH5qL2/SZJAMQoRwBWHs4mn/xgRRGKUCvSOb74vF5NOxPPJkP9W7cDtR0XpnR/O
+wOX3187ijlmGSGd/WHaTvemEPGlN04SNPH4nZwdI9ITp+ZLliL3MCmcEtSSccCD
nSlQpK77yDvymaPVXeZBIZPlVT2tmHIbZjlVXhonJ9aHL4sEMgX/yG/JCFEPO4Ez
fvIdnBQT34mQGgAJUjsMqIyyzx9124q6nS2OKX2lMi+0aSR64tIaGzZwlC+awt9I
ruTluYbayg+l0rC3PV2CvyQgTXdeMCmH3P2vjxMrsOGijmCpmvgoA/LfzVXUgYL7
vjTiY0fQ3diQvfj51Sxie2q8tW9GsRWtNwrR2QYuDsHTav6+hDP+x5Sl/iRGx++A
`protect END_PROTECTED
