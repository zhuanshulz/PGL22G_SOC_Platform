`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dfrMqDgYhMr429K4X9R0zB3Wlth9Kh0VAae88BsIORlsQlX3X15+2E532VPzsQF3
zUX5kkPD1FBd2IDqNNqzyajlpBe9t8b0sNvgfGx+xOdshl9436MN++tx6C2G1wGk
XBoKw8WLMb6LooI/bjujRH71SzyDBWxfYaZltxBEUHkNJMrmJAo+zc1R9F0j1xLe
V86KYDpwj7cAolk/PxS31wRe0vQMqfc9Z8gDexTL4T/Sx1BAbF3k0VdyETZV4Wvw
RW/COwvfcTMWvUqmxu71IXXvh4ZZSX4eJvi0FMskIMxo07ztRaHwGt7VN/w+Sky5
q9TXSGBisjX8p/C/TdqBYWiXs8pAQZqEpIT9//YcTCA5304wGCsQkN8+UmfYmocg
yhkSHG+tbCYGN70dYmRnyAQjJZtwfMND8a8iKNadP3ZNjsnf3QQLViu0e2LW5ZgV
tGIuLTLENJ9PHSpWWpRdWuOtN663SvP4pUZoulq1Pp9Qz2NKOGIYZFLloJlrMAqx
bur8xTvtzRSrG9IzsRe85aUnU65o9Zv7crwsDMj353TW4ChyNFb6z5cyK8ODYaZL
i59z7sE0CQjiWmNDRrwDiTBLdYXFwjxoquxH0qskHouobAoMrZHV90AQ7QefYm7C
U8Y1ApM6O78ZFXRc3HiWm5h+W76TzcGCV1uAg3IBTR2liKSe8Ua9wFXo+wsj6g+a
`protect END_PROTECTED
