`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aX/hxnWT6gGarMbK+avPM8wfMnWlScBdMuN7y+Lo5LNX8fFvEC3gHdZVWLz+FwAV
E64Z4PBir96/wE3PRhXFATJ9shK7PwPBSnbFYrM7kSZVugNvG5FIvGy30p+N0btf
MLnNSPkK5wNRmWQsOHZAy0if3Gpy/6cKr2fa3wIHAa9YzCMJUae1f9pUPg6IQChQ
IYGB14/CW9TvSGBVbfQdN79DWASOzi4S6SmuIDIoEq+LJ8uecV/ELrTcKbmI/vhS
3u065AJOIGu0HjYP/XYbK4cljm74CQYX6YAjZQfFqP/yhUNi8zyxb6uJ7FetIWu5
yamGV1hJ3moAKQ5IpEfI7GDMaG+lFa0T0kQMQbeQDqmVs1RoCVdOZVshFx2UiaIE
DJvAZ8KANrDxBqo7+etN5nawybUrsWkDbq4J3tDXUeKAra2gSVTN6yKhsPlyHiUO
LTVRmRnnOAVUwyVqScfmPGMkX3or1BNRCXe324zpX5KyV3v9JAaF/aDWO9qiyEAt
NMaUGup/ALaOOGu0Ore/+DEj9zxoRxvDkt2NdjX0JfumWIs/hvERNm2vPRTC7ZfF
T6OSiKjzb9Wn4dN6/2wJcE8rzB97+PL82KxMsDP/BmNicLJaFGWbT0zcpWtfapRk
Gj+eT57i4rj5OLxeXriJL95bGtUdiPiTwXx21/UgtOWFU54qeFMWGNRcI5y3wGZE
WEFe8O24PRtwUgEA6j1UqjiIVmFrOh3DSGjIpH69ljmv6QVSeHdEn1TCj+5SOjIb
BZ0nNeI/734dYdSUoGThXkUbux8Og4JmbYTcAZbX0cYmsj7atM3cSU37ohr94AX6
jLGseAVz47oBuaNCOK3U1wFPOZ8gKk4DuP3XPlsSDdQExERr9ZV1sMUS9zWHORVO
T6fLYa6aifvqe8NHZZu1LdksSZj7+Ttswvi+9pX65N44jnKAlXiQlcilG8+9ta/a
dZIT9tOH8nxb/QtJ3NisRWAu1sBkYblN7JyYzkrNieq1Qz2t/4kUE9OolZ1Zh81C
bsYbo7zj2Z0/FLm5KtyFa2CpzdBMiD1H2cNd9L886To=
`protect END_PROTECTED
