`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j/ZdZeCwYDkvrcJImbG2C2/DxuPcuocHmESCHlS0fLIfGRhOoWtCM2YJVcdWBh7o
+bw/MoMAigsyfICWyRLBXHlLB4t5jomcPNQhfdskeMEPP0PozVt94AVhA2WUY1V5
h1hV+A4mUf+pQW+f9RPezGwA1Jj97L9JZ7uW0/yPUyrZn2Q8B/yhlz/qq0v4w8bT
DQxrCy/NGCQM3npHxVkZawixiPhtbrWVHLFgc7Ab/4g90uhAMOA2ApQxRsPsGGOV
6HSmQxmdLkDLav5h6dwfcFaINW25TWTTSZD7ODhMoklufVEjXXd5C23rybN9+Yg+
mzGzYMbr7wi5VBEgayhWyhc1Z0UQ6VKObVohJUTQCqF96WFJCS/ceTASOuQTpCGX
b3zI/k6Ukxjm9GDvOVmP1bmk3LcKkW0Wnm449BZX4aXV2O+p51Mzy/uF5rzGvY2A
18fC1VOBqiOMnhcE3o9Z66zGCDIwsSVSDUQitCQ+kcobfwnO0IfDS2UXNY9Wh7mE
z8sca1v2w2I95Tzze5Puj7cGTxJGJ5h8kErF78F9/nk82X8zeAmtJKE5UdROmGs9
nndzQGQh5eoJ2KGCoxQh7xO31KCL8B+jWdOhIvTyLB6g89wBUo/XOlSuTk6m3Se+
fjhgFdrvlbCOuQt0n0OfKy78BurecLx4l7KMvDwMfZoRMGmUrJSwYSTHdGBC6Iqr
LvcKqwG6F6ECtMrNYZ/tTUY2KeMp9NLGnKakMUhpGHfpYqnK7AO8hV0dA87483oZ
88bzxGPEr3lHsWkPHiHwoUDaOqLIbFNi3rclJWgDlo6aoE6NsAxkUqOdxRyWcnZf
Gv7UVWJmRuA4VU5jQff5M7Kq4C3z5KqkoZmFlj5qrUjnNbANDvdEEHqH28JqgS1r
l5Z1lxrg9DsTJEu8Iluv7UawaXNUxFigyNuzK3vbPWmkFcDDqZGtlgMcW86l8uBn
+vCmp6DQ1XaOGQ50oC9zIiq6hHTKFnbYQVil1r3BR6zGXEevO9WtjQKYSelWhm7E
MT47ImODurtfH1SZ8g/lDZ8TUxZN6Qn/xM8FTRpYjdCkYhCCkS9Mul/+j+SzEifq
Ja6Pg9WyDxdYjdVFIg7C/l3QCvvJl5mGM1WzQWwELnJTdH5SlUzifPftUJKpkIKv
BE1XWi0D6ruVVWR1Buz7+pfBXmM6KH/BNU2nL+dXn0JOcspEVRZGmjuAiQzzZxvt
RV1N77pna70km1QFwXCOIHc80ejp1uotQ841PWOmy8TG4RPuVcyKyZaYLA879y2d
YqNUXoycAXvnQbZ5ib83tg==
`protect END_PROTECTED
