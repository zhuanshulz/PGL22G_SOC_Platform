`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FFAVIG8EGT/5CHFqCVRLcbn00gtBMKkpyBBM5jF8JmD6cPzzbVbWXR5ZA9nX1H15
6epVDViZIvH3PhIB/2eIRLV4lWqbtkEZszEFJknFNBLzBpeA7O0jqgpvezKQiuFb
v4vc68Pjzc6ZqZq3pLddjbPYL9HVKxTzjNlGoXJscDLac9ZKj805DKAiAklKA6ZQ
0yGz3sWf46McZMAPURaTL0oU8t5J1dKLrQUN/z6YGOHJ28t0ohdGJEqXW8ALd4sd
JdDFqtA36cO1B7cnSv7umUCKKQus8fFSxjJrlyTyu358ChNd2tnXetN3LlQl5TXr
k1rjtIJRAjbT6tGnBIv18whFEpGEG0RSo0ir6Wr+J4MSttbg3oT13qIBUTIFWBWo
OKBXgFJq+ofZNoxwUnebj7T/oeSAJ+DWwMgqoijpzryVX9abSjAoyFUHXNzIrDKy
oxUZwG9lRpY3+OYReHVUDihN/3KHnCeFj5kJtLm7gjPLkl89WmDIN63sHSQlAYix
AUajy7UyUDfiIapY5VcuqCBGt+iQpgoTABOrffNkQDt181UeDZ8raRL+xiPW2NG9
qHsbX6DyKbsagDTr6XyU6dHydmZUNWJE6dcNy95Sdg/IPEzra3Ap4mvVOamRn2DX
5RX0Zz0SQcQrvFRtyOrXPjgUTNb8x0oMgnWOvryhMocMaoGYk1UfcOo3nkTOQI/C
3G03XrxuRvErWI4Dgab6xvkM4lwPH2MtD869H2kgAjrrJrpNbiQv8m5fR4rpO2xK
nPD5p8l+wpiU/IwCOki8CECT/VCC/roirGCa4QDfVzHqrl//XbebFhxvHApxCZhq
EDR6NVhD4j6VsqoFPs8RLIUw6pKmCp9NAq88tF7Y65nzE2Wv7CDiE4nfLLs3o/wU
+UsRQXnQdhQGQyXZaIk/pyuKjHzM2LAGAP2j47Ze2am6kkex1oJAoERz0R6Tqz77
TjX+Or8qvpZpg37oxzNOpQN8TB23O02AHHNyiBUdYa6Su/tjaTWPiUGMiDahfmet
Tw5O4dMniWvl98XLMJa6K7Vh1GR58Ba9bohuOiSk4QYHfglH4G2cM3hJR8Oh2bKL
8rb3Ta86Y3LaO7948tpzRzEom0r+5rX5Rd/e7C8J87ESMdWkNLIehzT85S8qlub2
t1Obn5QF1cVZzSly/3UDJnEcmDouztRLEOGvfUshKtPLd7rH1G1hJ5JjIDXiQDgn
VJ5eAGrklod3xMwRw14xokXlByiLctc+eaSMYUyG354unIxOULGIPLB5BnWoW3b6
QkSqoVOapu17vTrCZE2fkwrIA+m4BzeB/+PLpHHlNuvbFUPmQPYkHYHJr3rtjylR
/dEOcnusk3kA3of8pfKf9crHyBVbyXZEjzcIZVpTzMSRR+DXxXKe0EhxbV7tiKCP
3mDITV45T9HkpM2N1m68gVhXvHFQp0H5c37Kn434EqErwG3k329JoIQ/SucztqkB
PAGlrFQTJ/4B7DZxVWIgekqJOePX+IkOBbw+QSNvXKFJtSMvPF/DVRwmdsgk2y2J
7dyMlJ40TTpZwkL6CR2k7Z8cJ6NPVpMB/cJNG8gu5pJzMV5vL/INsPaIWR+4FP1y
cpsy9QNHOi8eaS+uF6DiocKE97lDCxULWO+TqYede+lzXkwRrwrrAQZUPeq3lqYi
+MqoEir/VJp3eygbvN2SE5tu139iyle4GfrwPguWQfQFya93gfUGNaDbPzRtTiYV
dbGJi0PC0oaYGX3iHJSEXHkymuU24lz7Qjx5CLU/Zt6CW0yLe78aMkPPlahbcCzh
cnKzd3svmRChJbNW0NAt70NFW3BRx2Vo11/z9tlrCOFBf0Ag5tcgSD6e/PVENI9Z
coEJbBW8A/e9kEZMu210E7NqpOfhXurrwojCV5jCGcgX3mHn7vWQpqg/RlUg0LG9
2NYbjVYIRcYm4IBUJkKy8eSuFsglgSL2ol3FWecuZFOQ0N1tBWFow/0x+s8eVlXt
lUI0RiaU0LmT2xnfa3i8Ko/OJK0G0YbLLMRDORiNqvdL6x11SyjKbL0+ZAy0r0rw
EmEe0jWYl+pyO0wVfI8kr75pHaRFRuSfg1Kgac2zgTor6f5C2lSR73f86dGmf9zx
eJ1AhmuyQhvjzFXH3nKisSiubTy00t3G51VTI8ni8uaMDnMei+sPU3rff09VfdaV
iqbuULBVwF8gc9gXOmOanalAxIt1FvFSd5S7WofzM70VuHJD3MfhcZ6mpDkh37lh
0hKYPFI0+As39fV3rUchWrSsPVNjOexsHTHWFDSi+GUaoutsez4GfGRbP7Ae//zZ
I3dI5+tCAVf+qv1LWTj9BUksnDodWrg1652ZrDODCalYHzSECvNKZlJSjXT994tr
dngIxp625J2nFYaiHr9iKYjjp7P1rxzOiJ7d4zGVi21A9gyVbRpdXvdSkxtImmtO
o+smn35/epjuHyDswWXXod3dk8v9E+ZDakrl/XlP8ygfE0/WBf1664lj/uJqb0Vy
IyKYPsyL0PBQDGyLCGqiC+yM0gmB5+LtOQD5+KHmDCMf4xjc+Jo3TPz3WG5WGGfu
`protect END_PROTECTED
