`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OmZmbcXZOdcaVwliqeUhGnpwvpoExI/JzmqWXFjU4ScFnxn/MZ4YMukjABXD1Hjy
lEQxRQ7TeT22as12u9PaEi0sTUNi0uvDrihj8u08sZE2L+DRhAJHT5JK3Ev0809F
0Htd6rkrVaLmpZUZxojJtAzwIEe1NFd/U5/VU8dMqIc1bX6AKSQn8eQ38n/Vfy+x
7wDZQA611GJaWFw6MaQ8mqVbb0PynNxGGe7p1qXAB5GeF6DNbFVOcXQTFZeqlHt/
/WUvaPVivbTkshPH65rkmsi52CLJCYvNeivsGIoPZITe+dlXteLlvwbThi0kIyrE
71+nu5Bx/IIPuH0dutHugn+LCyaT2qcA5ZMY+PEWz64uRxVC+u00F9rm+Ox45wRC
sPQCnySURL5GI/a0X0md/ZdT0NBiTLCzeTB4+h/sXWvD0MV7hekNJrcfIZ9pFyg9
pVUklsfNDEUxJKold65GVHDULlbVlyLNR2Zl09SIfJRg+zqpODwS9aKtrBZUZmku
c4AlHPHUMAVwCuGgDY+Y7MCMxi10TDR05TkaqedG5e3rTBPEOtZCWeJ3r0txwd7K
y9ZgQYV3VnqPxHx7VxeXw4EnTAwz7qkyjAcpHfiTKc0nCmiAwaC3mGBCsl0Z57yo
PHnXX1hgJelHKvStY1ACV6iG2ew2Ytb2CNMvgH246RAwqMb/vhLMjW3nFq8AAKDR
EapywbxlknUkOrRj0BArcf0vOKe6Hx9DDzbtm7xS5I4mtd6Sl0l0taLmGGj1fRUi
KO7Ziq2t0zpm2Ho7KheWsOdA4HI243wnlftjXAVJmcIWS9zngBiWMQs0lFokV/25
Hdu/r7efEMPBJvWiEJdiAJgqx/iuX/hgAv7mUXjNp/X4atFhmTAzjvGnGNc2lzBd
2wTimJ96aSQqEAWxDwQpmv4bK5wTgLi7+vM4meNKM/cH+tYXYTKtoYhEpqu3O+f9
el5VWaxgbq+vb7yaIlsZoq1O/gIQb0bfyjxP8dcy2GwhcVgu31O10n6/+6mkLcef
NBh7fii0L8koJjsOsANz0uWhd0vcdsUMt8cN1IqLpK3KxXWPn+9AXt+m4ya3tYOo
/9KNFgXrA/mVznVLP+moyDcGjJXZVGqdOHbrI4+iSAfXNdymJHUa46SlDSatAMWM
gA6946zAoF3ixM+h4pH9ggfNrDKSws/UloGZQn0U6wzBcIiCkmf1g03vOJJxLpH2
5XfzjJMV3Sn1FTYleqYudc+UtmDaTVddCTI4+lAMqWJfMXiQIu9rrTjqnfNCjiBb
BiQ8hGeEjMmckoNI5pX4LA==
`protect END_PROTECTED
