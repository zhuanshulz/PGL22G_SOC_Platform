`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vD0NdzTUKMqTkdkEfr/NIaJdhDYWAR0GeEcnQJ79l850ydq57T2/TNySD3+XCesb
/+KoNq7gY/1SRy/TcbJFMubWFUshVS7aRd65LcXGWI6FQwPrtG5n60ZpDcgaNxlN
b2OwMlby/8myBjTwyOvTJJnhE4mdCOWag7MOMF0FhbgTLlF5bKIDh6Cw5mPsLUQZ
64gqtUfrgz3jHuPyle5Zv3je9NZgQtlnz0EgZLmQQmh+e3oH93yXKboPOcdnTaaM
G3zN+x0h+90BURWAKHDsyLVr2dPUSqqJB3NKXr0VCJNGxINgfapIEekOscUdchjx
03OdCDbLd2ogkXhGsl1Lcraii5JE626yjbDallG8kOj70Fx6++y4oNWWNFENFBRV
vxKXomKzmcu+JtHjTdG5UU/saiOr9s2RvRCmXn5CKeQhN8qNZ5XwrR+jslAyEWm0
sRvW1UoUCfFKmy+pm+yl/XUWKGxornwa8yLFDgGigf2GNlKQw8mv+D7WY8MWBGra
6cP/UoQ5obRfPOZfDrtsmdQWO00AfNzFej9z6YzE09z0mqGOTyEMcMoNkc9dzQUY
sMdp0O/5z3bxTp/HbV+NI2FadFy92x62YEfvJpnguSnJKElIHDfKS3BGKW415oID
cmEAjs4lmDWGaF53qHQcyY9vj+nxnqBXuwPdvn12rpnxLAGEzIhA6m97lJZvTaL4
AcCVXozV4bxDqS38k1Kf3OxSYVqu49smp9sOpphrcP/9NvTgxQ17GUp8s/walebD
MBSyp3n8Np6YyNrdGUuJiYMtfvj4lNx+A6G6rR1Y7i5ErhbDSUxEj5WfWHxNjv+B
sm3vlxT7tyZv7/KmSF9EN9iBm3zy6bewl+Bm+hFS7Vla3uQfktn8TDE2s4oqbhyo
s5pXMRCbMSPlBf1mRiU5oAIje9a+fqrmL75mx2r4gX95/FrKof2A30qofgx8SVvJ
HMBJ3KJx9DRlz5JT6Vxk+jTCO61xDqdgHBZyh/s/gb0Vm7LodG8v9vECqy6hlOrR
mz9N9jHgn/BSY8S0VIrE4WpKCC2rSKHUUr7VN4g0K9jjMmvr1x+ENS1NpnupZfqF
AepCK4kCwzHu0ZnT9b601660LEXreHHYGoU2ozAuYvb78cbf1iBP3fOdyVoUODfV
Lnbpw2JIBRKRDE6o95V4ZY0qSkwVTuDMmRSO2ZraGHq7unbIFFYXPiGEBKnrrqZe
K/KqvB9izyx1ZT0nY/uLks1zsYffTkG+4ht+6c81JQmAhyWaDBmhhWSUVhgKAdGj
epBDOSj+MmIKA2kBxfbxVanCecs/7LM3ki6mbqsCzbU=
`protect END_PROTECTED
