`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NV+gFOFh59lhMZaVa0NQ8jLRwcpjnm/gAsNhvCL3i2VuDZ8ZUhAV986C9vvtru5y
TECPpw48BclhuHvFZ9eUyD1eQP3jfM5Bkx+wiRVM4zZwxiUebWla6WPGIhLiFub7
H4lonnWQYh66zn3oHyVB3/fFUzvhBEgUpd2bnHnqomWGkGp90uYM3IcHdlISCmlz
J7/hP+HPYD4+/7GnN5NIqP7rzkTtIsLDhpNx+f0JQhsQ2xWfUBPL5eMsCST9ta26
07MYDqV2SgUh8CIr4VPGvQ==
`protect END_PROTECTED
