`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U/7RU295cErj7aHflj05N0zwC2OJ3iiwwsiIBYjnLMNRLU7uK+A/4DJOnYmnumsy
NkfWyLD43qykYKcpBE1+IlbLp5dVrF3jwj89VXeAKOnZJ+rZ8MxAXTrm0z60vszS
7wn5SgIScg2P/7M8kE41XTQTOelltqMwxg5RhtRlHsVypktTDr+IHZbnpGgUpGN/
46xRxv65sxcHCrEjgUWILT+HuwHXmdrMekBHkWHVUkwdKW9BKbNwWLhpvZT+APWA
NmDxYprrVKtcLkckQYpljENqfcF7vit45CvhPmuKEZY2BwwpLdjLz1E8EKMla4dZ
A3PPTpI1Atc/WEtkDOBlu+2dYbMjl0foSYnjAVsPmMsh2gDec6buhShRAqRL+IhV
+vfF+aFY1l4dByGO38BWQEErheil966wpOPSI1k7QK8sOefI3Q1y+oDMEV9aQDp9
FavgIuC0vtpouSyXBkj8sFW2pWeJmjZLP9sIcTRpkWy3IfwDZbv3uQWIiwAovxXc
p2YqHZblqdREj4nMd62WO/yq17ytJ8a1uZZc3YBh6b4TLXfSJ6Tn0/eDwYY/jXRE
orHMsS02Kg6hyyX6m3ZowouiJ7Mx5wFOA0n7LcLJefsG/WKhYLdq6Cc0kZGC6QYn
`protect END_PROTECTED
