`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/ZIA4xSFIq9Xm9XzG65szfo7kn6e+N4e1xX/TFQnJmLWzEZoHpFEdllmJUETblyG
RLE7WrbyVUjVqJDXmvRTrsRbMuGdoq7m4RcH6rRpTbwUoi2BWhvmCCa4afIhhF84
t6m91RgAEGz0/cHnsMbwtD0ZLHIbo+YjYu8UEKL2tc1iTQQv0P48C+z7f50npStT
7yd/HPkJR0dX19GfZQoLoh6Cewmb91I7Cgi/inQcowc674QVfnxqtepvhV0V4YDF
URlRzyYHrdj20xlqMEEijt8nkUipn9vKAUs9p+uismD+9i3gKspZJrXoZXA+RqrN
I4oFFi31HNCDH3J2w+geSK/1VrFsPWac1SMRwDO/lSuJSdkXpbf4+auac7lz7axd
2/RjcZJaAkwZcfFAaiksp+J2dkfxw9Zh5NbCdfBOdS7cnFYZrJ7KmuNTOvTkv7wW
9I/jlEyTVIfK43MJ0xEdmYGDxyiv5HYjBuoyEWen0KzHaj5xz1jBG7cP0tnwyu4n
bXmAWtZ8ehq5gQTrxFCNwRv1TdeipE3MjfETQHVbUCFPLtENUBAc91X1zC3k9jVi
PPD5jFN9AKWuqG5toMqpfwWTiH7oCGBZUsqYz+7yG2vGiirhSWP+XcgeO4wlVQAK
+yrLzsPjEf3aTzT3oFFr+RPj8P6L+S4fbpBCddmAwhkKec3FkctL2LkMmoRdt6u0
boxMa8CVGeUDuS3mniIYOWP/qyZiq6IN1zS2G+y9rJ6fk5VADFZGv1jkTH26d4xL
706TSjIUhyXwvWnhec1AcJFFCeavvYV/BqKnakNeznDS/CrO+qggUTPGOfYhtXWn
BQXp3x/KMSQ91WOLb6rn8VbqlrMsDMCvE1zrUG0OVCfumo6j7xW+bMPMp4mDZl2e
xWwDnpYtUGaC/CqbYOkl1E0wJLN/U69pUyBx5UntElDlWAVGaPchtKky6v6yy48t
1Fi3JItgzB0cxeuQYHDbHAt0+sASUuj422Z1aRH+p6opqF0hziVPAwJ4vmpKhVMC
LnmGy7cpQHGgftD6JzPZjCjHtpL/UP1Nnu3PlBy0KyOlYaSsoJb93XTnaUGBKckW
7TSxmQEAZDXbtL7juTnzBKDfS9oH1amprH+X1EljbpAPPxvB8e+mkzeipwpH/xUq
Poyq2W4P1ZVI1dAPB91FFe+KfCnWRlf/bM+9l5AtL13enc2kjaHrqCQaEfuf5Mn7
MceRvVm9nqHlxksGup/wyaCRJFxOAvZ/OWzgovK05L8rGVNJZSZ1BNICByTA8xOP
e63bCdi3M02bguwvyIk0VKuYKkc6XVezEI6azIYRKPJr+4cfD9TNXsueCHykl6Yp
fy2sNhORULviHYzYwdNTIvQNhuA68Oq6fYie7oi3dioRxP57/cSlKOpct36aGiUV
DV0rXmCXDFSNG+7zEg78DxauUEi0QtITq2KZXA+5LsXl0UjkU0GJA+vvbkE6SpVP
8aK9ZRpkUZX6GzIO0aeljlNyG7lIskCk0aPt9u6/kngPE7nnYDCToT1+i2rggNb4
/0kPZOymR6yzpJSqtFCDiGAXlISAl/Ae5esHSTmR/ecBl4ZhNgAz1RcmyBpZjSnh
M03jXu7rdLqfYGYnCwf6fUahV5ZjKhEPWy15s1kEGAmtRhxnSXuao6INERgqLq8W
kZMpkNUmn6nHGsH2HHU8sAiCMaRiZ3xILtgp66bwMdPv61Wnm/YPnD5rkXxL32Dh
haWHJj24P7YHNEIAJyfDFFdfNUZvCYkLJwBDgaGs9vYdGEraizKjyuX4GN91+Va6
0rb4gtvuY0cznH4mquQCyv4s+Yj9SglD94eBCG2eFOB4A7VWZyQS+acFgg8lXsVh
aqWDVprUwdj+Bt0DhDkU3vEyzsjULgwt097lY9lrceFbDHPGbm9s7UUR1jxXQ7t4
SnnOyaNmdLWXCfdM+AdJiuuZjQVvBWu3gTb2pv+ftLfE30/Kz11+j/XmEzbeV09p
zqJ/W7E2YEC/6gT5MChwUBAJvYsBzK/DYiNbEVdg9AVm4vKngIOj2Z77DazVfpvm
CiGvX2G9/c/aKLEzmt6uzZzbWbWghll9/IUMdvqg9IuBrPaPBrC9r1O0U6tenmuB
+DJZ5VC/MLKRkbDOkeMG6fmagu8pHQqh7prNM54sOG5VPLUlh0h7VddnHt3iC+LZ
N5LCuJMsEr8rhU4Amv+BYe2z4mGgytqwstZq/SQ2egsyqAYA2gGQCf0tlrXMDaDa
D/N9UDeXSdZgLWYx0Ctk4ilQAFuRZJmmIsC/ICWIKaH81ckqdoF8JbVRzagpg5E4
1mq4tXQoP/QdHG0ENQmVyD6f7Hx1aiM1SVe2qLEP8vtTEg5sgvZotOa4Toz5VuV6
x8v0RckpLit8xhEbUZcF4o+V26L/HUlcjiQcq6HfDzv1/R5Zq7wLLzloC8pJLtxb
aT0XkJMAzBdZhSCMyBZ1KOMuWEFJ/jQ4zYRdEV24WSp7iMHgkJzyNa80UgSA1CCw
L5Y8qvYqnUAEF9jHViFdZh1e7T2fNJyco2WKOXAmiUgqrNJzxGCDbfTwgHWexSBv
pOZhHEDsdzRYtUy5l+6/btXxy84uopoEZqwQT+pdHq/qNTpizaRVRJnRZUZ33DJF
VMFT4VHGPYa2EKnPhlydH5yz35EpJJXcdhtuBR1dG5jQAIdev1sPc/z7WqV7QSG6
RbVDGDTZz3oR+ukddpa7cUzwEEfiiJq6aeyig30sZb8g8SZjLmAX5WnGWv12NpZ6
NwcBX9e9nFlLkf7TbhdPDc1ixRCSzxHEVjb9pd5+FXxZhH5+o3/YMI2IEzCX9dR6
49n0ztBJau/2zc76WIy+mWtPlIhmtP/FvRxOZlIRCu7Zu80cRby+5BlpQMmc6jRl
sDsR/Z9ge5ygphphW3CDofmIuDx2HepoD5PC2McPOyRopz72g0pfBdoDaHMLPQpV
N0yMThHdLbi3f/cLEinyVCcR32Zp7ds68f2o2/p7ENH6VItli+v1WxtMpqtcnp4k
2hdHWdmZ7nD2+127KvIN8S/dZKBasCJsjZe4Za65A2JG6LZSvPA4DWJ08JMYhCnY
5Ku7Cz451fPTlbAevUPeF0MA2urj3s2ebbruoOBoAWfC5mmZ17UklCBJX3FlZpHV
dzE36edC9oia+z5lfEVj+9ain9oSeLxfN/mszdOTvDwnIKxQVcCrj0AaiskzR5L1
rt8vFb8XJE4PBpRri7GqmuyQ42wuPfH4JyLDhdY7H5cp09HLKCEQsKDGi8ZmQg15
n5nGXRB7MNLk7OGgeY5I60t6GYtx+/H27Zdr+FNxdWWJttksNz+CbH73VW7TBlj1
dEcl0VFfgoB03MnWvEscLbQdY5zRneIm9XzsFvH40Y46aoCgjiIfAG0kJaPS8TZy
O0D9Z6aw1PEftJEpBIi2dlNosXq5C/WjjTGYG2JDYmdZyk+d35PtZqJhwOrcw3nE
tPnd9tteteKsK6ecHfUD1nMpTiuLL0aBNF0rJmbgqqmp6tFi6Qb313w4Oewi1l2E
bQtWHcLUYMWJQNBMEcg8KZCf3tfSI32eV+o++ETTfgpNR7ygBxjVzoFoMKJlR+GK
McVWQGZgVmkbhTjKlG5Q9dNCjBde16LtBw/hEH2HatC9AvwICIbQiu03BJgKbbLR
rzOVEX1y6GZNc0pkMLBBLgmhDxBtroo5LY8djLb9S8ysFB+3drTd5hznX9umFsUK
ZOhMFiJx8jm9t8v4QOF2E74QpLZoCPYpnS3OGhJzClT6wLOE5zSCN7YfMk1xPW76
nwNajC4Y1mbITJuOQEURxDSDY4CIakybxdiUtF+5yVBkHQjT6Yp96wD+IfCHKBO6
keVWkbqbfnAKZsD0inCbN/aAus0+XCZPVgU04cuKSfpl5/fqElxPDx28gRcM6S3y
AMQThxSdYktEnpisLrSbLDI0uxaYXOigImDwbmx1mpMcvaMH+l1UvdVuU4NgT/4+
9uPmpD18yHvIgbr2PloWOW1CACQqet3LUmNFE8V0xOwuqMyrdO2cqFZpekIe8teK
a/FnDpMlHemex1vbAznjqJVXGijJtmpdLtDe0leY3QYiQVEmDGlt8Qx2OETAwtZ5
1OZfONNg4/eeiMfar3FgD4fnGIWGyczlquiHXj9SwsnZ+rH4/OXIfoIcy/H1oX70
ShTuRlGt4PTFxeuZnSjRIPEkqBbFl8fEtt7my2x1gtgrcPY5bPHrvum920ZtPHUW
3kQKj9W/BYxBxuri/KW2Pk82KB8xP2UNsXXZPXKtNo8AIGvTFZFe4oN9mTMb510E
786HLzlnUyc9fPe5c9322OiPNDjNA7/ogb1Atj6lRQDNcRLluogCG5P8dErJHECZ
Sr/kL2N359U/uVLmA9+h7+E33pC+/684ghaoVk5yRez6MWLmo52agOR8fsbYKe2n
P/Ac3ujpFk1WgHOcq8Hu5Q9aWj02Eof2QHjHabWf1v+RuW0FwOWUu71ODub3Vjnf
1uf5F8Mne1KO5L9Og7oBNYpYIek9iICsxVWP09rfk5zemPICfN8GcrmX+U87Mgy3
f1oTmuxZdciSzlUi+fFZXew8TNlYwqOqJpjGOVMGZL9A98NzNvPHXyMH6j6Cpihl
hq6ZkGN0DN9lJ7imgfBk5Bf80XKGl6DipGjPw4yYyrNHR26Jhtg1zI4RFGJW8J/I
SArtrTvmS7cbaEZnI5aWglhoUF9MBP3/aTVMUjztkWepUpzXrtNVVz2h8loaWN1Q
oDNBbLltid5MxqoEjT+sDwNCUdSwrEsX1mAszmV1rzsyOMUcgZGSrbI0KpigyXJg
0l8ySCfJRgoSKbOMpty9oMIOMCRC+My1eAPs7sghWAERITgpZAPvYSGbor09sSAl
u0x2wiaXwRZ59O3ab/0AyPT15qzlkDneRlTRtwZomuo8Qz3oG0a+5ez3obwjKfoh
DNYEXSMzo+0MGsXL8N7ZSo/cFbpsogSvb0MpGuazZITAHrFUIWrH0Qrl2/z4OeUl
yKa6NWphtjHlb9dEM5VyPAd8YGtYnk22eKkIXmNVJQYr606mrbi/kvj5y9aJ0iZu
zEI2X+z3XDzaDE3lpBYVpmDXlqz/mWYpZKsZznvYcH3JzXOaYObkV0V7FLlb5cjG
0REqL0w7nYmmgAMadzUt6WBf602eE7JAP8OdaXbZEKtZWMVza+Uf46Bl5qYTIt3U
PYmR/xp3/JtKjT/omtWaHuurZyvz821w6fEEhuo6vVUQ8QIRQ0zUEjkY63iqD8ey
jopGf2pdnEipA8S6TA5Sevk/nSKQfZLVPIqmLn7sGOyapU7nntUN/d9kU2Yg2SlQ
Ngmog0tICF1EavRHurKWMAN5beQeQOrwzWSVg9WXHejg56K+Mf+62vMwZZF+2Hci
p0QIddXgpQz58oZ49/tcsBZyxOB3vyazXGLDP0j6QWSG/PHWxFE0p5bOzO1ZdiwS
uH6TaItr8frcF4lQA4fhiIh3cY7YGysgjG27qK+aFHSy3Z0GHLnh5B+iyWbgmVBN
V53TXf3xhUhgP0IYA6t4bSTa/fSa2NFa3RKZ7JUXVCemRjpgrIEHfw+0hALvaXnv
WA9dBF+iItFIxNDAKi7ZgORSfbi4BlG0S6N4WQN/RnTMHyg1STwbZrPlMNAAI9bs
/Xtd8ca8x9cIRA/NFFEzBxMiMmYHQT/NydWK2D/uD07GQMEVaPROgDn+2xUlpV3c
wRwG6u61gnOLIT+zyIzYUco57FYMJdIaOMjxqCDinWjgtyCqed0XO8jXyVG+zt8W
vj5tEMW/FDNSXWFeBcd5ywUuv3CLweHPsn+OmfBPiTj0yNxF1tIbvgpIjgsxfv43
Q6b2VvtjxBgavLdwICxnX6oBe8I6U7nhelO0YhZpq9rqE1ibhcvl/lwCGFf71VeM
uqd/1bq3K9AXBh2luzHYQYD5+J3E3KMPRsWc0nmBfGLqdhGrDXh6NH1WgRGC1MMm
3SbQk1MwhU9LpS2PeKxrRQbWR/RiMNVt0Ngbbyo8hcxG5Ype4xl21aGICT6BZVfo
sHg7VxNrRphUHivMYLT9+u49kjMvApZHAlBNweIzd+agx3MKTShBq3uO2Ustd0HM
UHV0Tgh+OhUwyXtc1hvbeID6Yn88Mo6fYjMmwaKyX5OZvg6HD1JZWcGbaimX+fOz
wkaar+6tLBlEn8LI8rIr33bMMHj5PDwk/ch7O7XaI0L7hfJKAEvDxw83fBIDQPuC
qkixf7Vnha7KjNErLhbfaXFI5McTtcG5xeMAn1KurVIqjnutehMN4Ap5mc11JLjA
ZFOlFVmFbYXag+ksPabshJqh6/bp0OBL7qLgaeAAorbkjZ7KlC1kieK4xNLwz09z
srM1Qi1dBGoPumthcBrnG8EdDUycUO3N7I9aMmS7iGrw0lIIgwKP2tJidTX1WzIF
+q5d5QEYzu5IGihGcKBRt2ZOxSGSumqbGDUhifD5JRDqKE9btWs2U9kLkYrTZnEH
n8ZWTJ5ES5Tto26UM7Gamh1WSK698K+BqAuoZluzIcYtcdkx6aF8ej0B99kLoAFZ
dDutK/gYu+UZlw8ZMQB32B7T8nb3O26KehlT60L2CzeIo9VHbepIEhUVLcZgGOMp
W9czN1Kd+AC7kvitYWcDUqE7mmNNzl12s5j3uzCqCywQfTZVPgwOHvWkmA+oKVAI
m7zl80QBwqqnFiz9Mp4zmxWAlsj0UqYxRwEOq7s8HPYWtGanEOTMooQ26IMkN+Fj
vngNkohN5ozupIQlMp0D+J5lnLerZuSBbsmSYFmZ9d8/rrNkrF2Q9eIgM+fBbXQ5
/d13V9ab/eo2VpivZsAIXQEnIKoAEs5zcBq/HwS6Fhiu7g+G25sBZsY7d6HORlk5
t/Z2OEmhhUheM5KsG5MByvq2q2XkaWpd+HTDtpyCpsqH5jsrxi2EyuEseUaNVN6x
w5jAaEmMWH2GAx2ZUR3WpfDTS/3zKXt1nwrtDwiMEpoHiD6WCH/cKLvWWTEXF90f
Tp70IOtVbaes01dw2O1lEgk0fbWcUcAnVLA1k/8LgFh8V1TumP3lWf5otdEQW/Hm
/bTSbA6o7AyjTTq0TbSOeNY9G+DNd6SEg3I+NoQEtnMZZ2aTM8zE3t2mANTf1Ssk
4KydPP2N2X10p5YCXCOIdfC/ja7r6R61zuj9FXKnjc5p9jwslcJ+mUQsnI9FbxgS
IIri6fzr+s6oJleGH0LAS/zz8yKsoqVkPHMtEzXVpjEoZpvKnTFDg35pMVSgkvdj
eaCQJjRKPNyIL5L5VjS59PGYNfFXYO9bjjJU8FK3m6fnYkyt0qKQkv5JgfX7QBUi
VE98OmJUqUE/JRIS9o367HloE8j2gO/+PIJbTtVBlkD2V1sFDxxTFiDfkdWC46n2
rkDcbPX/3F3FHkDfsoUg9UfYzdsk1fAiSjfgGWOC781NxpCSyAj19TbPjKxb0k/n
/+U7eJ/CqSjnmxHa4AL/SUaAsFK8KcJZWKIteWjpIZs3W5h30wCEpGykAmhl3tL1
ABFdGVIBscEd3CsaqYBnof4zcCG6zjjDYcebfQaKG8jahSFeDuGMuK2QW8HeR/bu
pLI+zUV9lWLL9d3OjQiV1c7Slc936hRYSh8NE1i82TVlJQEth89Z09FSrMxDxYjq
lZxXyLPIvx5NaS0d8BD216q3LJmeMB3PP2kfeHCxceHyZqeSfS1P4y1NGPP7/RXW
vou1zLi1+VorMcS+VL+St5r1A/3sET7WsM2KMBjA4v6N+1wjQvELY01DtT8Ir60B
8+g2PTLTMxSN8JQdaLUNl+Fknj6ChByX4MAb0mpKmInb6I+IoOWJiTQ7v2100Bet
3+kFQ3pkicnDpu7nlD8dBP53iWO+23Oh00pyzSIvp42sNXFV9kaT6iEl1+bid1Yo
hPqzA65uvAjeOxDaro1bSO/kQGarEvtfTwdcYqDNxuRMEQtfhJdQJvoVxvuUtcQX
b/jzqfV/3o1cqVnysrbBV58KM8o4c5xEEInns30DHL7FrcF8PJxzb4SsIxrwQ/KE
8lRFygFS/7wJWzjkcxZrO+/aD812W8ZOyC3dXk0JdRgf4bQGbidOwflYPJPlXJQY
Sj2Ivktk9L9kZc8IzPF6XcovkeVu7ggTXShflY9cFP88Rn1a/xN/JaU5m+AxWFuE
Oqncm3go5oalVYorKJKCRZJ06Zux4eu94Sq37UKfwZE=
`protect END_PROTECTED
