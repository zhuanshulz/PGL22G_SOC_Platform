`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IiKojtFGgZVxQXJ+vXVROHZv9UmsmBa5N7u5mdrNEe6rv+zibpSsOK5EVUBz7Lsj
KHpJHt0dgeUF9cZYc7IXcB++X4+voslHQlbxquIdKsOkBRWqFzNDh9krvOYY0OF/
JDCQx84cywFOKG7dF78rt+VBRr/14fANM/CRpFL3ZsaR396eh0Lg7BEeR2cJn3fW
MUl5o/FzKPYBcUcK/l5W5npyuX9XgdjU2V9IJI4PMOBjUnKmhTM3UQfJ0JLZ4OPz
fRjfK/lp6kVpp+G+X/3eABikIAlxaDD7HX6GCsUaI9VkTvUbP8M68Kl7farW82J/
uJ6flxaEIluxhWOTn00lKTsooSFOL4RMd/k7e02DolXFlUSIvcNjQAq6NNm2U1P+
e84KMtNQZF1It2h5pzzQC+8jqxOZdH4Ky9owytvr5CfSF/6ydo+OUbmltlkRqmsR
x+w/rhflPYXlU/qK5Yo10cbEyaVa1+WyHJ1Ys1wH+/BaI/TW1tUwMCMZbvm3Kh+A
mrz90cOwqYH07OyJfQbynuOKnk26WV4xO9BJLE6zBy7GiOoqu7hRK18psc7XA0wq
9oaBQImVhjaOJ7sJkIXBxzPG6U4i8NVxxYVwmfcC2fL97YIWZawbK4VZmdc6P5d4
9KQizeXLMttOrEg4n1HzE8r9QaW0q96CofnpG4jlQ7FBQ+CSGenmNkcceTGt+xKZ
e4+UL1STTCRzgaJ/rOj2ROXKfvb6/HIuAgDrFvIZ6Oa1aezYGMX1C3xAg64vaAYp
VrBiZnkbfgl0Fh0usYJhRQcqZGNXlgwufN3S66L27ZyshxckWuv7IYxJw7yVbNUM
+YsPL8hXzaC/izPolmBfd/+kAAdYSncSdZoGHm/gyrgk4FZ0LgEdZt4q5lm1d3S6
51xol6QmiGPcjOO+QrIDt154UkWylvPgF1F7P2Ilr4hoHNt0CqOAk9aSDX6hx4q6
JcWrPClLwkLFCT8V12vy/49l2p2RD40T8GMdy+Dz4zhkoHoS+a9no3mMyMroEOft
aGYJu8QXOt7hSgPFmFgDOW8lIIVmxwNC25Ed0u/KoPk5Rcszh9P8xaYxzqY4/1xA
X6P3gZfxOYjq1jD5YNTS/r3vD4hpqGAaC1u6PdLrNMqmjRlmrLBhzyEzHrC5e7+g
IIDNq96fatMfVmoXxOF0Nf/91neHB4VvmaQwLBI99Hs5YK3p79k17FbLGRFJ9WRa
`protect END_PROTECTED
