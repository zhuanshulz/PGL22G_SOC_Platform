`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HNMPdUSAnGa3UbEY4eSDEZQC4RhJ7zcpgjNvjzOAwcRMf7mEpIJqTtvCcwIS8tLX
KQQTdQorXoDjCI4rtfbbsfVGsn8cjiTGzdh8TJ1i0lApbWyQYE5bw5BPVchOQXHa
2cB9T/BG/wQtrrIrU71Ydqvsnt7nyBoVHm43CrCOGNPOwSGc/19ejXGAhzngaCs+
lrSuwJwdVmrlnFoMMivtXI8H1EkG096RTO77X7ES/PWdm/fpvWeUkNFG3vrvAs1+
wvGDiVJcDLobUUVvSM/AGXFPQqF/xJW8aMo83G/YhO0gzEZL/WGon0bE9GaEX9+W
Ifh66vD1YKgBvqtfMC9dGFXP65e5kXuhsMSDT8GzkMTvsVIeH79AQhcAqxw87qIn
2FwfJq6ouxUHopDAt4nJjBzFyBpW4In+TOCnbOzEpUejxCwMlggEtZsmIIGZhUYE
hUzAy4CDoCrWWcM1UxdFqRdxXHruGo5HivH51XZVtak=
`protect END_PROTECTED
