`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VtaB2ib9syYWYUuWwoeN4/uekwtTbpkIb86/ROea3S9hVeWmvckUhKySVdxgE9m7
mYtMkUAtxyzcE9iBcHPIYXv9xLN3Gmumvsu78EG1C7UoGXs0qzNtjiofVsfLBIxR
VZwo5KRjXLWYeQtMSj2ZQhfHQN/CH4MKf4eWvXqgydVlJJX+N00hbFmZICmBISo0
BzUDyAm4ZZhnIKjdpNd+rTRcAOe7XmmrIAtTxNUBVR0bfmsRmHArAgbMZazB4sXE
yW5CECa0yVDNsvkwRP7Kgc+AWvBP6YSqqHxYXe6CiojukLAXUAeKRXysRhf17V2p
KJ1Yxhp3W2M3GJ72gBt1LPHsBdeL8jUvSNlkERZUXYvYh6OEAO7RIcR01S+n/SOa
o6Gh71F/mb0G5gezTfgt51zmtG05uCXleeGRFVdzJulwNoZsHZ2/Ibl1mxbf7EdN
ZgFJMo74Nmd+ZB3D2PLDEBdnu8PATKyFiVuGWrJQW87V5JpGnPIy90pYU5UvkX3G
FTmBlRac6Y8ODsVaN1aarr3SbAb2zqSAAMuIJflhwkCksDyQLSru56IqL78zcbSp
17xYfc8IK20c6K80KqqdmfEdPpT5q6xtxbO6CbR6nCoqOyIfu9Vml4nJ5nJwSkgO
yQxUlU3Sy9hgzgU4oeyztVefV5pIjkB1Vzx3qXQAGktbczYhVUIe2g34f6wc3rtZ
WNa3g302m0YNScciNvNLCP/s3w0eJLZz8CFdDMtCMVTkG34VjlmzjMJsb/UxmODd
DquqnYdpouTLa/In9OS8Ln5wovlp8m+eu8PqrPR9Gg7PmpdlZAljUcD0LniFY+kv
Xzs7eXVHsmR+1/iLWEwhzahs5U6tCWnwIHAgvUCw9V9qedjPxVrlVUO4kKgatpJp
IE7loCetq7l1xL7PnrxIag==
`protect END_PROTECTED
