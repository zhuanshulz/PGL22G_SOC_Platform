`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MvWgCNXqKgoF+HKA8YLYIk0WvKGwnKgGMgV84HVeKX2D08rB2vj+BXwrJ+yL436G
OsXAb1EpzOhvi26rspeHdcCpNRIr7KHiRkoRGsDqkBgqB1aHpB+o8O0z/53jSZTD
PegnPZ4v/JdqggM7yrWun5Rk4wrJyCYlAK6q3g+ysT885Aat1rJz1y3C0uqB1Do+
1b/4cvUfW5bT2Rdfx2s9jy8UiNrcaXvlFetqvq1fCZKsSxX5E/fqis/NaHA7OLFJ
F5Ky4/UCsEaRnWPTHYAaAr0WzeeNXkYDEe3zVHg5stLWHU9+WjGrYPKcH6LpAWrb
jXr7kEpHudC3h+Ak9Yoinfdctx2bxlnjiBpN+lWdBjnHPglf25FOrI57HIbmLlT1
lPf83oe0QIsWLgG6lSVjM7i4lxjaDW6GgYEbl+9Kg+j35WihM0HwpVmkHMca9O0O
tXKigxqDAJZ7vDYpmT9qyaQ9KHIXnZEux7KekSZ+69mIujRmNCVZMIzWX5vh0m4s
ZfOauc84t5PVmCueqvzagAP3SKlBzu/VFBhmaG/JV4DROCJynhOn/UDPighxSCgq
c0tIDFRqFDskui+Kcwknkfi2QQzLn9ZdjoshTK6fN6cSQbo0Pdytqy8FrmSl+iQq
FD1ndJv+yefHxa3ZeyM1Lg==
`protect END_PROTECTED
