`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A3Soa01sKUdtW83Tw8R+4FKPWraGlljXfHLxqITuPtrWoZKMTzEwTEYsSgo37zcz
2EGEuMvLoBDALP6ychiSenbumt/BwhnPoW4d8tDXF8LL7Y95zeKE3sidpHktplxk
76x5A6wLwqznSBjJ18BCdwm/b2t/iOC2/QmxTObNdcu/5Acl9mx8rF4gGqJNc8OU
8FhwZrserwzL9g6CKhxgTdYcf1xoie/6C+/O4Zp55sXO+PP2f1tXIbyV5gftuDk7
fdeKk0fCfS3U8fTMnvj4xGtLzG4EvJAFkkNwisi0QdSxyydi62wSD4PhEnQVcvXi
V6dvU2kOdBYlKVN2FYtQXChGeFVHgDqT+y3lc+yA8bsjPL3vk/yE/u+FlAptw6Vi
FvW/WLjVm/yVj213wPm77Hc1Zd0P0Ylm1QXehDVsB4ge+mEjcGZZKrY8Tkb5t/6P
IzzFSTTn386rcjmZTgwhc1wS8BLN9ziydWfUloUaC9NtoL+49NJA+0W/M4FWbZVF
zXF6VWVxJil34MV/DG19iXqUCfxA+ZhsoIvHAcP9/DDZzCVJ7jicip1alY0ayk+K
M9xMrqC4xZJCoqbqPpi1DxnI6nt+EGkWg/8qKbMaCJFXy5avxxgw7DTAvTHmzYfA
frZihl2XlPAifCHtrQhMv8tUOMDYmPLcAyVJs58sl+XLknY/eP63YCIoPvbFrAQj
zIA7tFV87vlnRK7xTSRhYEh6WKPJu0e0WpULPN5dUgHfmALl+xn1p1xV/gr6VSX2
8p1uhEwyoKwq17IyG+oSsYV42TMmIRM1zwskAAsEzU1OmQSxsXcSOtkTFxsXHsCI
8SjZipSWJWFIdijLslyrcjbvBAq+jQ4AOU/zlYiqh0GIYiAmgDoABUgCuzfp0ej3
7cGvKvJ+trEcdjSxaONdnY1NzZDFA4xef77uFXbOv5UCVp4EEYhhAHFO9n50mIFm
4ltrASPknOyLLPP2qMmJbPt+ntMaMA9MZDpVUlU8HC2B9aQ2m1B2zdRlqd6joebB
YsyHp6kt5MEInLG8f2gZrT+cgZ6ZTRABMGinzVOSTbMCgAARHQYw41jubmTlzOxt
6g4eo9TVmqpijl8aAZAHiRb9547OWxhbytW5Vv2DhLePpP2w6NGW3IDMDC9v3DZw
YN75iWdVhWM09FGoBj6E+3VloEAglmMdTol9cERTJdfIY2spV3PGakJrU87NzGt5
aUzgcwQeHjCzio2W40wkBYp4hDdlaTCV/dv4IXIJtkZHZlFMmsBlWoNFECr8YdmR
6Hlvk90S3MvXAHbQgo/JE2WCHuRg7ZsqgBzxlCZVSCqDGWPsGIkLrPPUfgvlqinw
gioWiMUJRen32i6DKdrQHCwF2ClONN2uWOfL4Y4qCVkIL76dFMWfhQ0cXFyR8V66
4DTXahcjiP5HGmUk7MWpKMNjO9tcsodX8Mma+aVqJ5YMhUrzJE8LfSUounXjlOoT
DnEpAnaxW5zBgtzmf71bS4dnHBEZI3EaO0FDRbPZnxzxNS3ve0huctQ394qQS6W4
YcP69d6LkDnyLqNrNJ6CaetaeOghreiC8RuXRjTiqzppqTigdxMbM6sW64iSOTYY
qW4b5keqo5t9HcxixytYtcW7kyWY4RV5qykm1piIJV31KQV3NxtcEUHuCOtsFlU9
W3T8UNYVHrFuqKnzNUekS9VuBITTQP5WU61fimxhqr/Yp73PbgnxQJTbFsgI90z6
ynMySHX/vDUy03iTkzmghS83BiWLmsa5zQxzfgxgHvitunzDU9AQ+MsyLTgkS3ua
2/Boy9Q1kVaZHNjrQI7k64rMzzXkTGAF4rn70xOm0xfdFKQfNQBpt4UaQChIC9PQ
cL6w/bzJh+2Co2u44wkxbYYX/5oqHY7lt6n5kcrWyQ7WTxTbfU1rrtmY0ERPJCgx
bY86Hu8pAfeQYO4DrWgTfQ5j3eZbORtYzA2vCVpjZMxpTs23jyuzyVjeei5nRlqt
cVfeiBRWB9rmimQCMUIjxpN0TcsVdaGIhwXODu+6YNG9WlVDwvuQtztWu3dul53V
UfK55kmZWVigpIIpPn9AP1okH7p1qHA8IfLA5Nskp3U0E/DeZYLjPyX9oYY1ZdQn
sVMtPTC1slZOpI8XdTPQhNexLT6ywx21MnBB0oKHxAzN3yhlnnUgKkwrk6u9l49E
NATyz9ZJSbQoxG4zX89WYIA7WltyvSaXoSBat93F00e1VSwW6d0t3W7V+sE4JfYe
VjJviihxFnjth9GEFWlmYhvmUjjsFNEBrCC5e/ADAnpkUrMFHC3//bhPfPpwIH4+
GgaMg0bmyl3lVdQTpBSx//ZY05pE4/X7ivSYGhSpomB7buP2io1WAQqlO5RgkxH/
DRiU31HPPwmiMmknFRhjaeNs2x3TqE8jIGceKCVrCVib0WmZEmjhz1PCkJwQexRf
gscJDUESoItAYOd7Kbpac/e4XQicR0xvZ9nTY4NIO+aKfb5AjH8fH6X4x5PMlSKY
PVPrsf6v5tQQFfnTpBx7wWwmaCaWBdPJA0h3q5EdrlmzuXGyBluN+4eo7Pkd3PJ+
NdzncDPhnmPdHlAMBu213fqiB+LKKA/vcPlISQJ+eJCEGe/UeHdFC2X7TQlGv1O3
fcxZIrRM/Zbe3odZZZDdf/IgPrZs3jcyOOuZHBNAa+h2Se1yxLgJoQkZlJvYAGlq
uhEE0MuwvP6FHt9phfvgnhpgzi/yGHFI/whEYCXwXWmR8BloiI1VW178o//zL7WT
Yw2QeuVZR63uyk2j0gNf1XrItGB5A9uQ/z8Nl8pXa4HCX7oiI0obZAuAt6ZJAoxO
DF8Pm43C3NJKYfhlFLDDBXo0AZliZn3eFThwh446LJ/jS3y2xhVzbQsICHDE8ET5
mQWrWuCn1HMJCB4NwTZnXONcAQgtc+3xHYX6LPIubzWWFj/y8VqpKvYTpJBpJHc0
QxT6kW95z6nYStMzjgGxpoJoFBInG/Z8lb6zpt9FcKiH4m5EuB0rPKiEcuPYLzeq
M9t7WoJujPYmTQW6HDX8uow1XG7gmrDxd/aRX4o1HkVpHaaiYHUP4pkilBcd7URQ
O32MLNpMW1KV2/62J5mPgd5/43L7s7+Q+qfPqOvlkM3jXMdFKRfmjl7QSSWmEva5
iNAByrYnmb7MwPZS51nsP6KLsCXxk7AS1g8j01WKjtwcIicmQ9TJZdcM4Af1q8M2
UWTKHfmv+hXU9sLXzf9V2Wgi+rdKINupKE3VbCjLFQFC0OpCuUrfykM8Jzt3ytpM
HWdGsXijA2IZyy7nlQBpryiJb1pomnOWgQLndtIYf6fyHmqg0yHL0Pt+JwYIiIs2
ln8Y0FhbBBmmDcsKpaIOfavWPdtIHJQXcSjOlsDMyIIqkMF7c8TyLwH4yeGY/fkO
HuYcRMjAJjgFJGSi+75QpNfSW+Mh/P43MZWA0BMU3kR2f57ApWe4RUzakhzm7lM0
RHcEXou+EcN1LsJzNfF25zPjeWYBlnbd+D0tme4GV8Z3vNxvnt4hHp2Ip4bp9RZg
6NXMOVoxXRU93xsNnuJK1UTzBmwQPwqUq4dFbEqk6qqqKC9JQ7/HFuaIzxqpNKu7
fIckyI40PpxSt6Y0taNExWj7yGw9PfowI9pXOENs8uaqBA6nUdds5XKTyZZIzH7M
+X19cAKzJxf3WHY3yWnBTFzO3bE5dFKdBU2OOUJMlfatulQETc8gB0GxjWQ0a1Sp
BX8/J+m3xRZMtrUS9/8e9CHEA65xeeG/P5L7EeIh+8q8fPPd7GSa1E7Sz5AMLegU
jyIKBbRtYKAs8OqQPOLkj8I0O98qasZj7u0i5Nqqn6uKkiEv+9rTHICOGMZR8B/+
flpZ6eKN3+6nUivxW0ZjCmpyrCHQ2oZbAdGImuVsN1nXAxRnPCI8KX6i18aVFl87
1rU7iX9VSGIUszFM3tgR5UzixihYhy+tTMF0IwA1YfnPgGx7FUmMwywXD6jUQyv1
dkgrw9+22cs8v9KynEspKaXF8sih+Ar3VbSPZpQ6/hvqNHpRyfLoZZuw3PXzLt7g
hvxdlYcFNFNhrwccqHy+h4aT3UkNclf2F1biQvHrBpTkJGecLC7vVXgtxfhBGPET
w3WH0wzsPTqMByGtoSS+a05b0Ngrt8muqG0lSt8GbEWOt6zW4CRYZWfTYGHAdxkD
FYn9Bw6Kiyeti/4ZVudGDIWZfqBNiVIf88yjYnv81sB4ANDxN/VeQx899L9LBa8g
zOoc2Dfj/BZ4maiMX2MLu2C4GxxgHEAzw5YrrtI2ul+FXvy/Fe5czaPndwayUorf
jAL47Y8nJ7VatPc3cPKHToPewcMn1P6Ba/8neuMn30/XE/QmHdGSiC8a2oaID2rm
rONTSgAGPvOIIAJh5bo/MScMenAFdw2xV/zZrQ2OxkfbMfBrCjY3PHqWk7nQ4Mp9
GpZ2ZnyP/ok/KlUYlGlHsptPXg32qWj/ylJyJc1SkGqitDMJg7ybzI7LHgU2z6Ye
xKaqVuQo1W/JI8+PpzYMP8KthwNOVxsm/UT0Ea3D0InUxKX44Rnjh5RCrnZumWPW
NA2PjrlchlLXYV1W1on5YYOcLi4RoD5y0diCTbSk8AJetfYwWfF+5Pffth/La8sL
Hc2xbvWmPh9lYO463hr4WkSQ+HPRCUDegij3o3sKtxbWcuOpZ7VN5CJKPVKdjwc0
swOjGDXbiLilfhu/lX6ElJ+n+7EiSJFWeSiyGFVKKaURfqJ7HUlJAAazZ72GiBr8
M+hUzbpNlp4zOog+VAx7grkPORGfgcbY3rm7EIa4YsthDPz8cZaVKNqjOggN0TEy
ciyIfAF7nZu9EPX5OhKpbFae8e0Km74WlRWeBE8pKnxIXapfYQ408zL80CM7nMMW
0bS2qrQxxku73zQm9IGrcKDJKAn+fQOnPlgcrycUyCWOzdTMuwIWvyFY2D1cuDpE
RdKjZ+TFa7I/0eVtFOFS1uBEryOE+erzEqyBIce9YqMndHyHiMidGd52F2svpAEh
lbsPo1iMWpQfMDeid+L1ZLrClCMymAbSQ0M0pXT21ipFm9GOrjTKX4FLDKkzhfq5
8WCcn+McwhezEgspl44PVmw757lAf1CMgPbNvriNUuBRu+/6YswcFfd5C8gi+JbU
XxahyHcxHPFC9OhWU65SElYfClgXBghe9mtK4Hjvvs0Ul06TUUUjZhDenK6QKeUf
+IDaS17jJTflPThL/0gOGTDWVlSWFxCQqxf3HksFaRXtDSGUNI2ATyhEwiehyZle
O16TrjcQ6QcV/W1W5vZ9JGUwgi205B48iacF1yVYJGrYoo4ho3zWMMBeJiomFZFi
b4lQ09hTa0PGhYtXlD2vcmbnzxEuTd9MghxNamggs/TCJwj8BAFNEJUWOhpA3E5M
3qaNet6m9q9AozzOux55hR4q3mLa+vmAvmGd/TUg1lbfBwhQsPKEzILve+wlyIfu
7ztQai6s3mcJ3i6naWk8TE21E9FZh54EmN8TS4B/rsMLd4msBzG7pbhX33nKikxk
+PpgeE9nGXCNxiyWsbCIdHkavXMkte6L7oeF6fswBznplazwSpCMk1STLVzGqk+R
Eg+7lN3I55he7rM73WOUcLh7rPGu1CJYkFXhmms+tmReeWvQOygffropco5PUw0Q
zuPONysYdclGwRRDqJ2eB/+MoSSmU2wK1q6aY0/Mg7UUseGlIeVorC5QVtssVtbO
O9y8io5qddr0bP4kNRx26C5aqgwRhIMX6DOP5zDq64esQJblMGEEQ8JF0kzljDoE
P3FuUKnp4A1XlSPc1ak25Rza/nrzzJeBKtbuZJGM7zTu1HMB8IfL33H88Bhfbcrm
cSdPi9URHqeQajwY4CDdRbcSPRxxTVxlocSrqDFjc45AA/oCrkKB1A70pRB3RUrg
uDlOVfQDYDPdzmYNkYVVI8PXBcj+GkBCYy7c1DufRALwXTJAFfjRs9jMvtx7Z/E4
ksgPn/rCE7+8IGswDAEd+o95vTW3zPqD+Bp6SUO/BbZQ4RhlwC6A6y9N0HydlPou
v+RAppE3DHB6T0tmOC5ZoUfn8LhOx2N0LthmJUiT2Ad5EXRdedVCzK+qhn1ZdNrC
vhSXHvRw3nI78T0iorOXaMD3Wbpp3DYl9cYfYclrztho3RqO1sgsefa6nhzgNqeb
gqW5YsT7ldklPvJgHqbwxqlKdpIcB3Kyf1wR8rizNlg2AZZzN472mJVFSBo/xRHR
WOD6yJgZOebfp+P3F7sr8NB12pecJlOrEK3BFUwyV9lnPAZebE0t/JjwzeoN8h6U
KAuZWT5c6bbNH+LGAR+SUVBry5acHBYJJuA9KjzcC79Z8PYg5JxIZGM+PRPoGTRK
VJIzELFHsFZjAEQkf3C7jT8vDu6ftwMwvzoHI76MS3BtO58dRLkZAfwRsjDrCHUY
nLm+ErKHolvm2XLn9xpO7mZe91f8HyIlyFV3ySYR8vv6w0Qfm1iOe36mZqr0mD/6
LvtuxCHKRU9fVvIxXW52UGc6L9mWnnvrqtdazECpVyqGNxQIF0QqirZxuLgHZrw6
AlN+J7gVF97PSBi634e2Rz6ERB0RfsPzekZDwjyJbuA904SNK7e/sE8D/3BKPEer
9DN3Ruy5yUc1UTVQd5+JCUuuIoq5YnL/UG79mecIQBlWFkBvvBpSVoA6REDwcgUg
JiTEkRY+2mqW33hvYFMRRccvsFjwIb0Q/2n9FVb9G0bLDFYrxoBdv2vq5dskkRpz
QypHyDOLGXXZ3MvXHl2exTqo5nqIraNSDb2QlkUD6hES5ppcaAQfyEc14mDsncof
7N3g2VAsbF10c8uJq6u2tSDRzhjLVyUD+819h63hRFJZmM8buXS0/6LmR1LU5ZUY
cn1g8Aye5GvStPNngQriSk65MGM8onBCP0qgwn42iOHoZQlbk5kvvwj+S83Xccr7
lo7pwZQoKziv+lIP2rVaWrZBYbxwwCZsGxUDQJHah0odsMI/Yu3DzwrLQvsgEVrM
6jBR2iP2JVKT3QR/iA59cox0Fe0byAAmyPC5gPE0zTufKaSwjGvBqDO8RpBDC+Wu
VGQWUfrceT5pxvd3HVnSfRM1wyOictF+QYR9Vp19K/42iZq/4ebcxhRvSnORS6F/
TADB5aeH51hExi1Q67fCQWqahEM3PC45IXJrhItUWFSZkH8uKbxv4djlgtsehzUz
9RnhoKCQpgQziNxUbUX/DBc57rDA3gpww/yqAMWrnxL0UGLBsmAOg6GRGVEEiu7a
nbXKaOTjTSAWPfwhYHZy/Y5orE3MlAo96u5ssAEUztSkX6Jtuz/y7kFxgJNi/Bib
BuucrUkH8lbcuAS4gVtir2kKDbsa+E2kOQALU7q6mqk4XGG4+IpHaL2Ois+NIj6z
l/d3sL3tRnfoX+ANkbZoy3ubEQrV8MlZI4WhuuHhymlIMeHw9aAloEL+FAQbnb8t
vwiE+ctJND+FM5YtQdA3hXGV3mCyYSR9NdgEj9qACwcz/Fz0PAqwfY7gQMtaEBuv
DnCvaYpZR94CZR97iwoXHQejJ4Y8Bgy8/83ZvQ7Br8GqxVSfLhF/67FSj/ZPNLjk
keX905ejOPea7nIkbaoK5MtYVZMrd39zIgbG5LNVbW6Jjgxqqv0FASoYPG/DFUF3
bX9MAlFQ/6ZyTVxcdciejVuTHFEdn52HoWvY+y7w4bOOF9Qao1qN8UWpJJpm0JzA
yEZSh76uYRWfyG2S7cBLm/f/d0iukVT2zzyaU0HMEYfpga3C/cZR1naHYgh1NUOa
QoSEuBLtYdNrhODtn8aE6TnIiUS5uNaXJWn8aHR646bY2BMtl7AiXjTV9z1XiFfW
U7B/mBuGf0eewtDfPRwXsMoqf3uFjRse4xBTphP3mhNJ46J/eTziUWtHkwPoIJEj
Ikq7HsYm2a/d2i2qgtd3gldlEsH3aJ3uf2ELI48NzW3I9SueYi7/wemlxv9y9Z/R
7qiSwyRPMPg0q9hPoQ8lwR6653KqOxFxr9eXjHq7o3G7RrhyLK4k/wZqibKOeOB8
bZyd1PntZAp5Xr8uMTIkhg87AHZvO8uQKe2NAIhJL/cgHffzTG6FdZtVxgs7uDo/
g1OGhxYbe5i0Z/DO9Wa2ScKdB+bRUw4JQMc/HMNx8wq+81FeX0yYasJ9FJ+sQmzD
FEsKqg/BxFdgdjFkEshiJAJvWQJ9S4wNi/PiOVcuHulSxZDssOMQWcVl8AkZb/55
MMHYUwHbo+tQA0gUMqhQzpjK6VJlHljBw3C8BbTlqkYs1YmTsPIwaHJlgimmWWGk
ImrYf17bZvQYpQskmU3R+IWCY494truXdWKpAIQZ049NrIF1OqChVySP3YhazS1H
PalSGKEcYcWUkUOA2ouoqOmBRZB3DqPhbJOBJqweh2kSwlijnF7AasnSfusOyZv+
0TK2qYC7cWSA8iOEfp1F1TfJQo43lLYcej+ZSobxfzR1V6CsItpChe0FNWkbFnRn
flKzGwNP52UZ2AR994R68lGVQF1eo6eVTQ7YmHYb5aVWR4Tm7ydCF5fOPhFEDKpy
gLEFcrc133gP3g4TnyawQJyxQ0W+fkpFCOiS9FVPqJ+ifUxG7Ih+w4Pi1WnDbtk3
dqse5qrff6+dvGk49774MKo4jE0Lw43rpGufqEF6lIuT0/6xNi8frdGBuTCWJyXz
87EHlB1c+X0aIJx+Xy+rs+8QVXuL9fo54DIFdJHoooJbJo+p/Lm2K+6L9J2s876z
aC2vawsvJrxhkc8BWwrWLrqaykuCOsGf6NgRccMIiSZR1+AmSSb2hved1hw4SocN
2LlHxkMObRmn6YRqSiOClrDXOINwgMU33Ku4MfGYAKIn2yDYeZm6NwcbFTRZnDgH
2KKlILzwpOL/NDmzYFxU/M5IDGsFqcLTAM/tVzUtOGLDqWFP7+6W1FBDCjFWywPT
Xhg7Gg7iH17W0/kM2QF5nnXumSUwJK6f+v4vbh3bC2BIIC/RzVv9MlWvuYezcuOh
U1qK/ZOar48Gn1QctwzHXx9pIeJj8LsUCXV2t8fMfEc+4bxISB/VPRpQ1WAbN+rF
0zTyjKx/BsTtkoVAKWc8tqnryyWb2vcupyiWsV1vubHtBA/ZO3JTWbrrWMFC5ISN
VVcyL0JbS6A3t/Nh/rrJzvBlZ7iGzYnQ5o+7tO96X9lnUjR/qHUKq09X0cPuFT8N
pNK4COadmZqKQsGBHswJ6ICsdYCuXy6lGDePtsbVv+PF8Oh2W2A+s14QfpiooGFD
lROnZojW1D1oBbvn5GkOFH+SFJ4WCk/KGx9drlJK0KGnRRm5tv+7tu/NqEwGFWhI
a4Bl9P6Aid5aZYiOhHB3gpq5IF9Y4EQYIinNefHQCY+LF6fQnIXDp/5UWo6VPWQe
mjuPjANPcLNYxDmRMjNOMUPiGydTw7qYd4Ine1qgeBQrnKYyqcNW+qvYKgNwvfsz
Kv1VJ+GlxEYO7hyTiO4xLwgZ0Z7GYFmViRhQpnu1cO+06/uHr8H/MatzyUMeSIfR
AurG8H+EgdFMkBql9/Hfbt7n95vJu5zLANAH1Eu9ZdqDFxIN+3SfiUJ6B+V4gk1S
3AfcQffIaxHLEuQcfaZxMQbnydj+f7S+qZtNxX8fpLQX14deZr8N0/gp4MgphjP+
+lYv/zjN+W0cNVdikinMW9s3+Kl4CMo7HMH6XJmKSBqSTfwzuVj1IzH3LN/M3HX/
zxlq0cTCIw4HEPQT2CDB50MLFIqybLxRdtKpp7IAkZogDJJ+ix0i3ZSeEgKqYDFw
/PvUHL32BP7thwzS+TQ3uZFkvWnSIl7lPNKGdoolJ30gnkqeaGHhVffZz3V/Kwp0
5pfNQ8kmgQiHnxh/6thBtJJ5jN6ZcLCsemIuyP0oSfC/1V+G3bWeSY3zYmQhZh0j
XSVip6nWabsJoLTxUNjHfcYNbGlJLwP9cV4adkvrie/CbEhdfqN/NNGBvv4iARMg
YH/L6+uShL8XqdT7bsUjxbRw5qL0l1WrgyVVwKIQ/MvBK1amx6sN1MkUi/XKYQFW
xkw02pZnCtGprvet0vg5WNSxwoXx2IpyslU2xMcZFJO4mH/ijjVgSfKMDsEKtbxk
TlSdJNQeCwh2n6+7Nz0W93XTZE3xKd/AtHi/BrJEBsIAliaoOiwNlzDJfl9O0TWF
GDDXBqrCD2rod13pBtoOIVutSS+G+q3BOMknEk88kQXBBeNu/Uo8ewT1Ml+nIvtT
9W7i8meifzBjNf7i+ZrPygTfc6r0JhhqXUzxUJPpOS473JT6f9gANi3NU24gBHY4
zgy62rcN8LxodJh5J7ix6w0xa7hXFGrKMMfw3XJS/S8guWTiegEu5xjiPTGkWU1S
hW+Hmi/ybtR9LaM13Cxqb7luDfCHYUgwcVpgEl23wVc1g/2TTT2r+U+IfhO+kHI+
hjh+IrVUu/qE3o04LaCToyO1/1DlJl6aQscKpnEct0UW7kUWCC/Y+Ws0pqegNs71
jvsUCNYbZZSeWYJF+GYzf6MlvxAEOSYMhe/Z/Yh3aNlimusIPswrfv/23sw8nlTm
asihk7JIE9wM2jMbXHbTfjjwvjlEoNRGrdFXRFnl1CgGRwVGC/pUGMhYnUA/PuXq
mHCBQt3UbwmEFhEg4s6f+LfmNHq5kqibyOeWHHYfPIFLTi0o93BWHkOIvapJUOop
HMyzOFciNbAwEbBOiZSt2bwdJxAuGbOqO3itVPS4ajOkCQmf0/Zp4Afhm+/ZeBuU
fO64NGgnioLECBxOU2cgnQWYGT84BrQsq86u9pQ+2oCbswKuN5HwQE7VBlXwBhlJ
66NGOYT3/gA+ox16uW9CHXfkl8M7nryhQU5eWzgsSq+X4YXIomVdcxTDe6LJX2YX
h9fSoc4PkSz53G90oY8l5QM6WzoznRMx6ADFJZwrblqOjNYdCDQ83qRJOvRSnSFk
i4DdVOIHIxQ6HvEDsfXTTagoDzXwUzM8uojmYjZZtuCKUjANeLwrgG1gSYXghhJe
nolC2maQtxJMbxnKUbmktsLydFzahP7tgZc4oepbrlyu+u6+XZsifakZNTMiMFZl
upe3YPMZTiy9y7/HA40iZoOi6PMZlWReGbzr4KbAUXWhvOkmBBz9wOzpjuYV98h2
uaqdmqhWHaQuoMvS3vkLhYOYfNyrrOjdy0T2j4QTYy23MKxuHMxDCu4GcQKQkzNn
dlQZQS0meFDpBtx5T/0Cxx6reeQsHb9es465LKdRGAgLKc3o/r6CMh8cB77AxzYX
pTqSAfueCddXb67nQOu9QT6GcF6lYbak0s/MVXGLgd/PDACHnG+mSpQeXDLnGoJJ
uerZjGpyIX++CcbT2SXEwrViqhP2N6hZO7t4QS6N67VfH8rIwoJz3Mftq/AkYyDM
LgTxe9+ysNCWI8ikOmXIIl0xujs+07Y6pcEMgHazgsktlIuOjJ7STWQaybifczKD
Xnp+Ja+MvEdjOGt44G2VrDq4ty/CtGOQPaPAPbyqtfU+5zqjUfyQCn+djUiI95Mw
VgMsvcerNm97GpFqAoQwZaFZHg8z3cz0GM0/+Wu8tg32CcuMrBMOS+hYrF+ljsyz
902g/zRLskXJTpMljaLa4T3kjw5DMAd2pe7g2t+WQQ4NV9CYAgA+IGdRpbTbJzzC
FbCJq54wjiBCA3zRSklOVWZylQMncAePxRa5wIVAe4RYDxZdEnyg76VGf3oigWGi
rsA/Z8minGh9xc2iSBf4OmwASB+rOyiaa1nq5Q/+xFCVz39rE/aCTghEdH/zhnFu
IVgOS7cQayixh8L5picOg5bMvc4rSQ/oW6SLzej/B4OdRrDzb1gX5+WIbJG2Qp4M
2SEBpAzyea11sPkUlCXRuj5kd2YL7Q8QFcqpMklq5iVoQtFwJXUOOjH2rYq1l9l5
dd8xGbJ3pEblLeGmQNeBbhjmjF+X6Rr4zSSE9rVlHs+2AGUQSIGUJm9gMojuIILI
mGsae0fCVv865dmAw97XYonMVIGHFQAXAyIGkfYmXDDueuLZtLZRh2t6yUC5rlIq
E2PlssLhxnqQSYwSeaWkskswhc/KFFDXHEasYcYbPqPWtrY4wQaY724R+CIlYtgR
N7tH98vWnBUCH04LAXEuT86QPWn13n0Fttelfibv/sR+WmcNt5yPtIReqmuGRKij
YZIWMKkbEyu7p68GFYeiQOD4O3XQSNTuiPjFLG2KER9JX+ZPBo7sFJuf1ahNSsOh
ZWP/OGtT3/82+AnyQC/khRCfQfEBQEAgY8n+FMhQq0yIu92ooICqEzAZNTY5VerV
rl3aXrDGgNrKPiIpyq/wIL7zKi09aXObcgunUXJMhnnzNACqnoU9lham1GwxKuma
BKwknaF8KmQCG6avGy7b5CV9QYWE7ywz/vsRDC9Ij9mBASpaF2786QHmNjscEs11
/N1owz/0UgxXvgDiAo9ka8iT/miVWs60yuF7xqHWDtqHN6S/jlWjgS1Jgpl4iQMt
a8cTcOX3MYXsVB3GS6NMClB2WLGgQMEU3WJqxbVmzdB+lLICtfN85dsltVBfar9k
j7mlSyjfuTdWC9VWgu0Cdo/xyFzdaynNuV7uFer9YZtBEFp79gQLYFGp0+w5xOYW
Ba364Lmm88YMixDqxRGAMJd703m7+m/CXfgYEWE/JNNpTwj19YkdOVaRArRLWkum
fp04JXhopmzVFrTwNKcR51KzS8v0Euis/gkbnyhz/O86yHv/8sLxAUT8pk9rq/eC
+MiRSrMsNE0REv+o3XKozCqKjma4e4f5oXqVh5hdFYD/UvqFpMl9338kgqYlbRfb
HFcseLf+fHN/L4KeqCOcUnJNmmYcdZD00jzmBExIHuUfe2Q9/3hma3DjT2NCM6ns
7KyzwwV9bknxfV/IKqJvWvyba+wXzusSAqBnYA5j6uesSVGwkOsj466/EpiWfMXN
D3pmY51uo1yhJ4Y3sbMIVm7O7U7x+qLYDc+OGlAmph5E29a139lYcfeShisWR7Qa
df2p2WckKLfIVtXl4ctc5cw0WEP5F7DkbccKceZLjlg5WxgsdFWWkO9GzdmtO8cL
jK22SnAptDGdpv7/AgplDo3BTZPCfp3yEq68degmxviR3FoIkskBxRP5XtdARGWU
m70dH717TG54FdGTiL13UgpBwZl1x5dxlZFESHQFuIAyFaW4d6atKZ9/lx0Cc+Ok
PglY4+69MhGH3pbA1mxZbkHHaekqKMb7DL5nB39TTKYir9/9zgSTSDUphwrwD4Ex
fY8WGVX38XIaGKuEZOlW1rNtTCa82Spc3dF9tBmreYARUTWWzyJmZtzknFjWDarl
W0rImbz9IcQ3KAYQqg52kXzZqjIu9gABjl3CaOxD4XD0H008KMc5wHAC8IJfCkbu
WpmRHPD1Y9u13jFKxbU5Rdnh62cPl1ZiHuBnUK/fz26Dv/JxFSpAr/NJmcDde2gq
pUOQL2msB5D9pt+J+jqTCkIbAgxyep3/ro36rjDttnUcYRMZH1J+qiwG2W9VV3Py
AACBl7PE0hH8yEzVS4/l5p1Rz7EomoNgp9m8dA6oLs8UHPK8WsvwqkB9VXLI7gmj
2t+mp0F+2lxa29lX3bR4UW1N1bBR2J6rjKNT5HDtwX5rYhwlzzRpvmlj60+x+9R2
CkM02I/xCgXHh6jtha27H/EoV3wF0XjkE63QKr4Wz0dLIfi6W1u/CBDh0z5Ur/33
CeWJEKN1HuQelsP5+bmLOm5JkKxhhaV22KXDPQ7oTH4v72aB8QdPD+5CrS0B6LTU
6VJaaO6dUwtk+FgdexDDA7s8UyZSsYSA5JovMIv91MLR28qC8maiMy44grUZmB59
A0zaG5Wl2DX13zNjxv2xll3+QEx1ozG4W0T0Ds9gKwZo7OxizROQY/F+3ow6qwFq
6dOPYDsjesOlogOAi9f8B6z5lqCtVpqi6SLWfxPcMWjzN60dZA6OyEUidLZr/F2Z
u/+MRJnfblTTQHI9KUg1j2IoCxLwOXCEs3kK6bl1mMDGWJlUZqabZEqjUwQ3Xs6F
PzC3rXYZH8Exj2MCZWKIdzqTqZh8yjfd6LtXKRzj9zL3t2/3+7lybdEXgSiNvEIx
zlOYA7xGK/cAyI/YTir3zeLw6aI/Ajar2NVGEy2mgtdO+jia6ElyxYIPMBXUeaWB
WBFQKXgV7f1yHp45PBZPytDyR0O6B4150uVzZRLiFP7EmdxDOJWvo21tvoxeivLZ
tDZwje6A5EJmN3VZIqrVJuwrtRUTFLjaeeyKQHMazyVjM2ltxmp99sfACsPIpjWd
lloEWWJ65z1J2bKj0gH3uvwxkL2GDyuQ77B7OCfOSMJwVX+b+8EyCYrCOLw3QDfc
mp8flJf4U70jffGbGTYVZFlP9YB8BonABQ4fJA2IGazh4LA4k89waWtVx5ohj2FW
vrQ4GHBQRhvANq2vGA/hxWZlPm3HRgW9ZpFcFZYuusD5fEQYDcp6PF5yCACMVgXb
y8ttLgqSLs2ke2K5GuPXnGnQyM/a/tM80DTE1sr1Qy/wjw7DmMGSo01l2GnPQhPB
2y0ae48ywj9bfarJ8o+K5CKxsV4y9v5hrfRToSFFVoJ7RuIwhu2iIbXJW8RJUcou
06jRqINdlUNQlaOFO13OOAzOf8F5C3NY4h3ZnRiuiaGxb/9UePrUVLep2D19yLq/
KFEZvR24IYEBjSP0Sl088DkoJTUdKVSe+vEnuExEEuVCKET1avJqSyHRvIRQFyGN
wte04j8eXNDWQZ4Fa1B9IXxmOB21r+j2husFAhnvMT5SEnJkGwx616OU4+GCa6dB
avRn2AoQaE+0+ux1+gZYrtWfSbcRLlH17sHx7h45puYHQ6Wcp+U/epAVGP5YBLNq
PwWScvEn7c/hkpQmg7q6aYdbFHvVVxYNfJWE25TrkqW4FNrGNdhLdkM2ctt5XckS
lC1wy2/QeqZ7FmhHIYiMHup7KT2VyEFXAetEdDDvY5sVdsNMOJVdPOSwO+/ONNoC
1pSddBUREfCwGsK8Igk2vtq8MyJnlrWUUicMkCICBXr0FqX8yYQ04N9vqq7IWN4I
husWTj/C1psXoO/vXErBUaFHqYm/WvEkYoZ7jp7oezowMpJLvFZMAfgaWLV9dFD9
5fSfHO7SObOIxR6pWOZ8cK7u1qDNwvcX0P7K+fDgqOh0UikQlZ4S8JHzOsjEgZqf
mKxUorNRGf7Q/Gx4LbEL+kKu3VKK5/FCICNnTekE70z0UKYlFdfqCz0+Fga4wZa+
9FK6YKsFCprhSQ/eRc42e1cjcVj+NJYRLnPwKOY8/9dgUcYuUHgnZrBCLYuJC6k6
UY9vu5FwTppxtt9ZHKnUbac5RH+P40TmLzkNhe9B1D2ETJeNSlpABU5k/8k9MFEO
7qpLjs3CiVHFZ0NcHAgt1bIIYdAa+pv4YeJW/hKsVBh5QrZCXjOA/9yt1QddYgKD
EhbYLyGtVN7ARnuxjbipXYnhS2a8qyRNUgnZh9TDr54gfpEarQYEczZnVYxYDPuM
S65VsrNl0m/8bumbv8j+h12n/0Y2K+DNvdzmabpM3e7O6iUTJQmLu7wcnLiTx8F1
rubIJbdSw3cz5FCeexKwIYzV7LM83e/wwwRnM10uRu7kQ0+XZ/cf7JC83bi1Y4Db
PMvn11Bsyy/hTaLwZ8BrnU918vSL161o41F4JEOYLbuty2yaJiQm7hbbsLwo0daR
FfJAcQ6O+V853w7WawwBinR8qx0EsnGLH6C8DpsTWZkENvlGBIgGPpzyq9Ltc/Kx
Eep23ftGWKD+bHiB1SPll9CisVj4++FIgBLlArDPteiiqSMEzeKq6/6T7s+PTZfo
SXZ6tniwgsJTlFnBh2XSRXNbY2OpIGSSPtLOe1z+Q9KaOXQlqztW1vY+CA/NW6lU
H+sp0LYLtfgnB531VV/u7oreW/xv8uStVizvxRYN7rik4f6GVbGTSDKCYQ2JpcFx
EWMGGkmnDpVgpYy2Mt3BMohlOC1cJdeRAsoswEWwy4uEVQPlb/GM2l+GDEkVHb1i
l0DHpnnxz3ANEASyb5NGxe5w6pWhFNE1L5dmIJiizXaI9WyuoYnvyw8X3TQFSws2
ZFr6FbFIzFR4OL8c+0C+BqwDfoX0ntue+e40E7YoB96hUOzT6V3/1NXVPcEtEE8q
9fLnsPkj6vkasvKkZAws4ZMHMZpXHICpj0c3B9pVGtqQoYzkyhPbdohxqB+3LbKE
OrU+w54idXYjB/nQPZOH8EisptUDZJ7DauWNUXfM/RE+e6kaWBQ85XMBSAFxDPiC
DL5wdEfLLY2lr6xFwdMb40gsyvmg91JB9FIe49VhjY3s20YSr1CPf9Hb2RhDblfq
w/ZZzvyhAlOnQ5jMwIU96/mZFicLHHTVDsfrYrTGvcGzLelbItwrD2tq1dO9vZvF
ZCZGnqvCaU1n7MRV/oe/yqk4KEtoJzky8VoPyswCzffBZjx8GRStrWZxNU2a9orw
MxEJY1P1HIzX+TkfIiD0wFKLjO39X0j/MrY4Z9bFjZ+pHcromDLxX29nI4B0O4qp
i8tvn/mgWz5v/hgVKGOHfBjndLR+E/zrkuStfXHtOpukKGQQUxq1jSMQwo1BrNRR
QGhEwMeB05flc9SGn/a4BxT9U8ia/dNoex0DjhqCxtWEqw7Sf0rf/mBe+UpqVJtn
gQuFobczUfFG946vPQQV/v9jww0TznZVyXQmlgHwFT6aw0Bjx8/gVYoW73c+BEnQ
5T3YDnqFFCLr4zJeV2FarO7Pr30f/a8oH4Ev/rCbC8lJA1+0GY3ObNI7n6ekB7G1
hyoWKDYnbd96pEIMETKS6oEv1wP1rsf/FB1MsYh6YaLIcHh0b6RR38dymukLr3Xo
aGgUbDeGWYb1QK6NT8CIbSTgGzwHH2YDVtYEbkP4WymVj+qiCs5hO8LhBNzX2kdd
A54Fj7qEE8hwILyC4Lq1C9yTSL/Fsi9a+vc89uZMLtN6xAvIIoKeEUJOJAL/Xk8e
YTJeVbzmw64owCLyuew7OR4g3Q+rgSyxXAa40nKFMUOmo5xno02Nj8+/QTc0W2dy
gj0ugcCkdmFd1bpC3nxF4i7gg4yock6yBVyWPzuDK5NsMWs4UiSse/5Elci9Nt6Q
VGKcvBNay1g/qTTYO+o/89rM8Ey9F1uuAE0CzBXfh6DGAx61LN/4mKIQWQgHoBGQ
mUnLsRiy/gMDVpPMfV2bwVqrWMRMsHDy+eID09yuA0lnIP0Lut2/tBik6PRUSGGA
Y9QsaZ+TWEja3AHGLfTT2ttp3Ffn752fS7/eG+DFJVXqmZyJeo2HQhPJf2AXiETz
X62nSFggrIo6goWLPgIjC6NKxd20xgOpmcVlb2jOWnRHk6pgTF7dgdsd3EGYeUGc
hi4j+GutmpaUVYQJdQ3GCdd29XVH0Zw5qwb7EvB5Lzi0QTFHXdvhIPikNyk22Gdl
QYMqfvc13BYbmCvPCuYHItMTwADFnhR3araYOvTpNUQKAGOm8deZPyri6t1Be+cr
zFaIhhnsseSCPYVEod2iI5Uy0ID+zzHPJkQlJM2As0yrD52S2nMExvQpa+yHgNW7
yUvEMKVGRpjJT6Je3+vnxek4Uz84HQ04bikby3VgAFzPrhEzr98RZXCYHeS6J75g
oJoHweXcih5f9Eqpj8rlwtaFbwn7uEVK+jKyZdqut936P6zO4qJyF09fqlC+k3dO
Uxzn+1oavOl3NJv0R1wndh4aevS+VKKwHjzphMPARjyDD3MPNhDcwf57zvHvFob8
NTmfQJKIn1T/FUJk1tKJeypULBrRNwq4P+aDkfdPPJuNK/O32SgECMwQo2uTvsl6
TW1hMUPuJFk0djnZz5Mejcmrg0Kcs9dmC2DGT/ieHSgf1a+xW23Lyr7XN5+MwIkz
lxptYQgfExwMtipgnRehIv1f2EghSsQ/ZeeRPPsAeyT7RJ+KjR44f5+IdatXEEfx
SSjMp/pbyIucAAuASeZSKH4Rz69nkLhY/XTeSeATVmUN/rXIjTckHsZFqVWhDhL9
TN0Mx10PnF+Y1TwjuqpQHD5/Y+UQW/WSk4Ej4OOk42LfIhfvlmwioOvjBUcuhCCe
KLyYPtceFnJEe+oT97h0Z+nmZ/59vl+bLv4YwacFYDjKA7AMSdJRD6HiauEXCX3h
5LOwP3QuhjBbixi0Bd1ht8MyyHjetRWM9WcxgMchHcbM2ub4Y561xQJ1GYjbf7NZ
RpMxpEJxzaGdBStsNWy0ByaTAw7PFBl7LWUgIgsBX41eOVlsQNFZIDHSFkSS87s4
G9kBrMv8eQjskDoYYsVai57nMRuF1hUquUYXG1FJjlL2raJ5hVVCw/JjoO4jDXOk
iHIFiklXDsTYMM8QujpZ3uk6vcXxqFwHRAUhO5bDZ1m8qb+exQIkwkD9X1kkLYD+
MzxuM2GxVLx5uQ11CNcX52dabhMF4Ji5uklUfmH3DelYbIG3NO91q32TQk0QNmGp
b82zR6Kx4MLnj659HsBisvSKv3PADjx15H/bfOrPJg8/FWRQBp0JPS0vGQQmPdAn
v0Mcme3kymYaB53I/HoYtBa9MfEuGfTTHKyywIkOvE57uuRVmYeUHQn7pc5IfcM4
i8Nad3AX7vv1k3nhFNwHobElTvScSedlyG9CmGxN7OJJt1YICjFa6AsD3wVQ0vrB
AUUS0QjLNpb8OUd2TXab0DaKap073VcG09hxzOghlcrEZlw0qG3nXl/1e2EufxXM
KZ6/s3xsfV4rWrdSpz0sD3yneNMgeqOUY5LxAvImrnirM0ZWJ21r9JnokZ/seeQJ
WxmscHBwWg1BR675EdzDCnBAQGeq0OYUaPRsuGY7UHP7DbkWXgekoTwNCz3vX0mR
dtS9E1xu8zIBBY66RoouRC+hNtCLEKg5xG0gabLoUzwwqDnCY1IDGrzvCqaVytH/
VKLzLbfA3grMsrFf7AhZKxzMdVbRQlB5CAsCOvIWPqbq3vsQtdI360AMGtoThZA5
20JU6dfflozwd7YnaaUCFcmLbmjSthB3XM6vaYOOnYnNkoJaInGVvoYuEMNvIdGH
DDxlo1X/Q7MWjchNZhYbVzxnjZgnfD0cUYvjrLYYNiO+uXMQiUqk9yl2GH3NS1rm
ImbN5RB8mDrB6/2DwLRbkP50AEtGBtZNEtXIGGM+5DxswjpXQ1W4xFKKJZhaJb3j
eGqIC6NpRaUnP0PkG0AqZqEy+4rg5RPXZBp3M+asoZfjHfX4TWYH4recN++s2dfw
ZFvOFfoc/bg+AnDC2l6zT716/UVohHPjiT76XyzZAPGf1fiOhSIRgdYl8swGOXke
wkdKMhd7CyscFcUBnI+lfri/ImQSbD7JPTCR7MRRdzXXuzUUm3WFaCjLaBO6XJfc
nCedYLetliPzeSiekNkc0z9plnu/ti873SwLOHTOf+QxnCjogP0OFgOM1+Bqi3ON
ikhbBRLC17gIDn+NqbZpi/+a6I15JllITizufkOKpnCxAi2HxS0oKiqBy97/72Jf
D9bmZmaMIQ8O5Twk8nEUxomQfTX1aS9+sQprDRGuZtiEgzM/cZL3CFwvgdfjnvFD
b6A/XOKh5fJHSljxYZJVe8ySNrrAwoDt9/qXiG7qj2neulC2sDROfMSU8ilgoGso
GOTDq4oRD95WjtrId1Nm+ItX1ST7LJa4/3pjh82lmfHz0lH65TW7acrYb0G8fiQc
Z5Q2oLXrcwnTToNAXvNEejhcWz6ZGKncChtDE2E0AI66AvCnEVQEo438eBF4ILhN
ElIXCEByHQOJ88YpWpnsFV0TPmOEvJztD2Q2wwOJwCD+8ni/s2BuDyuBgB1H9QUf
TT6FOWbExmtPIEajio5RSonJZzWkfpdLt3yo8ri/BeDhBjnW84ZnuX2Iz/pPDlx1
5y9ZFscJye+3oyZ1EjjpV0qXEuwhLDqzOWXppYiXWBXcNds4YTWyZk7UN5L5rSua
IEoCInyjjHARx6kocBg8tAyFU8DHyUgsJBcWaXFzpo/SezSZ7Z+dXwUVK9eHJMSW
5VRTSvUMsaruQTL+KxZjAGETlVNZGbNqpmyfK/8msUIOYzGshv4JpzH0oTXsuKKc
wJH/PE5gInG/PeXa3tnfeRQ+OsIq4o1fCEnYlFWY4lsOsO6jQb8WZVS26JtBetUr
eMioooaO4x7+iDW8nYQiuQkFOJ5Yl1kVeZDKqlNt873/K3uNgMAtCGkmf2jEADwX
6kwsRyvytRBfDT+U74uWg6cruz4vE9kkEnZac0u689KTffe/9Y8GfMRsoYllbbX5
+KgS/PaP/iV3S1H5oupFKv860WmvHaqAQJ3g4xL1+CMMfVtvbK0tBY0a7RjPWf5E
KF1jLQH5Ml721kctRvG4RWCO/7kQ3i3iZGZxy2figSO7BFeOsagA6yA4HPOmJ1g3
U/2vT6LrauqB8CWfonq5bpRNC0L+oD+j5AoeEcJTrzPe4qy0m+fBywrolSql9Rh5
b56sxMxwUVPJAW4pKIYj1Jk9eSJQjYvzV3A+9PGdsUzUY0rcZshH3aY0QVjz+r0p
Jlphv8hkPeTlqG+brOHLwf7NcaL76wDbau33FoGhj+uGUuCA5YHZz8S/qj5k3cAk
GrOOi9BqCe0F37Q+TPKChv7NtTApjGKJfyj7UB+He/cQ+6mi4QSp37Mv5YN415L/
QYqPTlNwg6X69BBeNM4gg+Y0gCkNTsfMmGGXOzDJ9E9AKSUtp8W2FWeiuLDTi3xf
YEXdth/k1HAAgMwf8UVR89PZmWEVC/65eGKCz9oWvE2oUQd5H0NF3MzCmTITsJd1
T7NO91JWNVyJOqmOVzJPlAJni7QprDQL5SvHZENRyytCwTc6dGGl5n/xDJkrbfaT
Pq72Sp47Nohggk8G9B1PLQyQgPCazW77xawtVJg//Dw8xdUyN1mL9WCDgT2b31gM
OUDMuo/3ZrL53JWrv0MwY3Gkx0xVipSoa/+HYuTWuUvBcMjLVAx5ktDhQ9LjYx82
D8XJdohAQ8OW/61ncchsY1bfjR3XAuy63IHb1jTMPIYVlquLVP4AbP9zMDq33ulx
DDDBc/hrqR92JGlv/YPCBebXslIaAp9LSrUkXni/tp+pRmV6/6X6/Os8XIhreU9U
d10bqAtjk3afc2OgSX6y0dHz8snB1RmBQ35mCI8TrPdkKyq4qDWPDknJORCfqw/+
jSAjSZQ9KdfRfDCLX6wj4lCJ7EIU8coDSaSHDcE45fhI1bUb6D+VYhzh+TIKhI//
KWwOaGC2gZ1GbTiqKLbb+sr8FMNmIJAS78z4KLMm19+hs5Wun+js8pGQxgo9G/+q
KopJ86rsscOm2K0DOzRwIhXVpxQCOrDWAzIOLNYDHVTRWEqK43ocGNztrRiEXK34
JU+0L9/ILdN0deT2iGp4xkK2dIsuE9S+HagynsWVrOBFRhe5qjX8Rl3Gl5leyDbQ
v1JiocfwPxgeDPsu9g5SPZfx4/HQKTMCw7cGVxVBQYzMrz93loPZAO+cugCLGDTg
LI1JQXQGYxQw05I3x+l1KrgkPt/hGZq1oxuW5K3V+XKvjdc4yTHP4rATCYJebm3f
9pVy2vnzFKkdYxwRU+kFwfcLJmfuDI/4BBecS9gO3WgzyiIUsMYhYwkXwe9LLFV6
oyBIw1ET9kKons+ZGn0JtkLDylXc/oRh1OVV+TrCZXFBFonid9l+rtg+nS78LY9Q
cDuxFi7649t1AT5CWqOVh64Xg4udD3XXU7WVvNyc7vGGl4TJ64dj1/ovTEKdah33
kybfCII3vJs17ROfvV4aQKuf0tX+HG8LV4Di8qmuv4hvEEcwTBxSRz/ZhmIpzGl8
SP4l4MrfWaW4ZMckPNfNSU9LKrX3PwIKmastYKXtNHASlxpbqOkbj+SX3RPTsS98
lCviFlEEDOmBfe0+Usz532bCX3gAJYiOKgMyjidkWWtGFWcNpYzWxF4dQiotxLxt
3pjqAKwPjvpgkyrRmGpA5YgTqIBf67RZKXWsNxdquBNro5o5ayKLtd7nrfBV30j6
6pBtz2HvSWj61drCiNwFkWw7A15+xPmtg69X0ZGWXl1SPVlCJzSBLYV6kR+8vvaR
VioiPtIzT3JZQlzZKBee8O29zHQveagRyQphw9g1xylHL8h4CDf71/OVQCV6s7+V
CZLFvvrILrnvfvIIFHPw08lIoVszt8knWtMqGIRqu8zls38EHbd0stFbPymxF2yi
zWuDYkDYvQ5CyQMOt33Di2FwCCTOKdIzMqVZRx2zfIoAkFNumu2naNptwZC2N1SH
0SkjWSdkPN4OPIcZCATTYOIlSr9YcoRRYuot97BpjKD7bTjjfPzotUhFb7TmVJhJ
2kS7Kgc37GDEONW8u4AvxURZD0nvfZxO2/CXU+YMmDFgoW7jzYSeozziyuqSTNJ8
fiVeoKsAq36MWn4zWWZJQ5bXMbdb5+/gOoGSnLJGKO33ku6m/CRsiCAl9gcMh+OH
JBlfX5xeKJqkh6yfZAVcktb/UsSWai+My2y8376a+kYZWWslEmbJw4+OJ1zSIwIc
tuy4egr95he11GnEaqRpjhXG2RV66UQERisRIinvhlx7twBEufkjH1Z4W/G9BTS5
L69aD9mcpmYe7SZXZsZy0YYDA+8+gFs9pwNHmDxN3InUUEVLiZgkthfowNlDTyEz
D0YOtUgq8OiF1eGwnX8yKN7BwbJPzfMoO5X7McA2dqw6DKDN58KViY2oiFyI+poZ
Ak583RRG322NMLbM8qgx7rim2wESneMhwi9j9hCZFfuBDS3BEiwwxIlBmQUN5+Qu
jheOuFwXAGYfLr/2Jn6upYFvGQoA7n36IYoD76vuYt482hye44BF28KgrR3d/tIr
rJVH9Vo+rfVJjyAyPk03frm8nag0rMN3UN0eEGqKilcOpVnbNhKpFAXpNOc4hC0o
7A0zftUCoMUZK+ye4QkyAnkolE9GxNmF0US+nlsTpHKM0hfPgQwN/oJaKDBoW/EF
MEg1F1spmX06d8wpin9ltILnOoJrasJsef1KdB2T+Gby8BE7zST10/QjUEis8J1E
cdSxFWuFcFDsPT1HTdL8EXX4+RxqOPVHoOb3k8OaugaaWrfBYledHTlsoBgeHsvZ
BQujHGKxQ0zagkjcR2C9E/hpOh2eFK+fH4oDZcGHUIqv43iaZioKuxTGuchxm+72
wk/nBGKPtHZ63Fc4fRlxydlh9x6jssOr23+jtAMsQR0zRtu1dT3DEmQ7TjjlcGig
U0goWNBE+rw5fAWtlrGUit3JTEzwNOU71Cad2AsM9CkcprPymKTjTWZyicKk4X3r
gthSuT1lJMAqmKREfLZy29UTY3BlCV5KuUHIq8HNpv+At3zoo8WJ2NaGwWQSFXKz
h+AFyCK54XA/G4RS8Ne+1lp+TsaYUEMM81IcbAkI3WTF4RlM9yZmyBwyJLIYuEwv
RAh97AbVIsMWhYAPoAAAKfbXl2py2A4Xl92k1HRubsRtOpX9z1nhHJVP6mu5nDPw
QHqCCs7TFXXVqvBf4UocM+Ltu1HG8mGUEgurhlqHzxlWd0IbKgZAA7u9b8+fB3HA
NVbJzHLAIuTov5/oAIV7iPDb4jsKJPJHHt/8frUuBkQKoX61mSLwSVObkGEof2Qh
ievUwC9M9R9fNZMTdCicuqUn4l8Zcp+J7+NWZF7FRO3qMpJ2cYcFUWcn8HDid0I9
gHGedHpXOOBHWKYmxKyLQBPzvRWYdQ235Y8Jra47oaSZV+dYz/0y010aRBeQDLAW
wynFhlScRrw1Gk8YdIpq3Fa/gwAbwI4HLqrk5FHfEN1UKfHuj7+rm4F2KIlROm2P
ajoRilnpVlUtw7TJJegLC3VHCGP3iXk12yQVR1+SjERBlhDpdplo6fHUHkYTbndG
yjYbOEG4tXF7lY0cCMOz3a9XgomwrEpBDXWmaie9sRmnOwLixRKu8dvPPbqdDsye
jPHX8YVWljSY12upd6buPI3ttWA3GnG93BDezZ5yHDmMiIYp93dqEjd9JJYle9oW
XKKXyYFXMAS9k2BZ9XJnirHP5K4HA+Dm1CvPXMzP2DbeeANyURO+oGb7WLN7Gtss
5HQfjs/+vh2aHzomXR/XZXaya6IessSNsED7sj22P1kWuvv9nNKo4xJTZaKbdQ3o
eOqROYZAtTEO+GeODWVMSyS4ZsdK4Sa/vxu/exHJOoLR+1fMi7m3oAPjVqoJ+tu0
J3KX7O9qZjixRakd11AE8466raQFdyUJASi7BwqW7KIyGQtGCZu0iQpgNCsH8vv8
GZF/tigr4idhDJJMUQXmzV2YP9Sebj8alGdpmydcPgvLvNVWJc0TMmk4J5inxZlo
XWiSUCZWMpu47BCbTG5bvYfMb8iTdm2XLWwk8FOBowftSE1UdftslndYdFNUR2CO
AqK05qOl3MBQUVle4CrF/RQAopVn98AnvDACHkdgnbNpFUQI9ZU8jg3AkfRgCmBu
DPeLnqjbOsMjl3qEiL7DQY/bIfMZYl+vG9vax9pZKAD/0juFDC4rLQnoVRnfnBxi
0EhpyMEgPtlkzmL8zIh31YpQ9QZKuJXx6Tf/hRkgQy3sncmOnWYbjpd89wCXOYlA
R1CQhuKIfIRKm7FZ5gk929MFfzfygf/fsP/Fs37jB07110ONCsXFYAt8UGbk5WHl
q2UP7QLpWAvzBpd+HVHS3GfzuLIS1SkLnpElf42YrM+lBEqbhLR7hgUJF0v3qCEH
rapqHxJv/pljUbsKvmyQR5GkpzCQDKlh1srmE1K6TPqmDzXDadTjMSHnQ5buC94R
iW5Pzghl3+o6HTVd/a3UjOatbsy6VvwcoocKR9T8RY83kmlp59ehqeo7FBaL4Fji
NVi1eM8qsHCPOh8H65RqJOhRwexbPqcrtj5THqCzCOx0WgJu3xEWHVn33o9/U1Cp
/BcLZG8fcFkH8K1qGP934IY3Nx1zDYYo5FmqqugUcnZNJLAmrVqvBZE5n2eygKUq
WGvrUmlXoUYluYZHnShpcgHRGHcEklroZxIOBBFku/a7NimmnKfhPLJZJLRWzCgC
qT0tdoeYY0tsFn7rVyo/BiBriOt0rnmV1D2I8TiKEX1qE5lYsgC8xO73MLtYnF8s
o0cpvLeMS6oWMUYAFw1OWflAmZuj+Fdygapnt/44kvdQP/+mmGEdbGiqHDklOb+Z
CVy0XAmc6OQU0Z+Et8lk241BGfjbzJuNmL7Rl+ShRlnI8RqlA+6hN02sQugkIL7E
wndjnSFMvyDe4xAH6MOQWWVgaTt2lHEQm7gikZLw9OoOi8JrQyjkpUHfKd1eFggy
WurvJI2VAkE6FA8BVuGIDrCnVUC9W3sEa9o3Jq3Do1S/I/IlM8uSo1FsVpICkxEA
6qUAUu4g2ge3LygUia2GPBJU8oZ2/1jOo6oaCDhsLNwO6OrkkPZj6hQybalH3um/
lDcoNhfqkeVP5khtJfGGx0aCdMSyQAOoOt04El7Net3jHyB/bB7Ia0C56ROyC0YO
AM6dncYzUICFAigyD8hiBqzh/1drlGEmzgalgo/F7F5WW/OY13gYhqyvb4lv+G8z
ZdMwMqt9M5fAp0PM+ukqmXiaCDkVSsRAAKbL2aws7GC0hVC0dxzqaa7HDAdQd7Fh
Kjz4oOZ6tccI01wBHX0TWcb5tPamvfHO0y2pxj3JzJ+HFOVTv8HC5R7aI6kzB/v7
MyY+9AnBkjc5IzQTRNLz50Kw09c7FU+xsG1oAXh+/ucK2KR38hXszj20JvV6i4Ta
x2l7CtDZKyhwQF5+SAbgTY51qx9wHnScWdJhkSdT/D/oJT/SVc9JA5eqDxEglCTm
P3nclZbasC4gKJUaeNsHKquawL5ObxMdJ3sayrKqiVEz5r2EsCZWoLcWbNpveDXe
JygAdY/DCxaut2ETJ3x6q8squHHFJi/oU1V6iyPfSu6fZPUqW6iIfCozmklHiyk5
rng+ymh3OMqn5O41DEHWc56DgkGCROHvlXGh6XqIrSeEWMdQKt38+64egJY+CVBH
a1WwhqxpqOXVaxPvkAh7keOHDj2viXoKIeuNQTyWTSqsGPMTaAwsssJr0jhnGAB3
7M5Cp+dZZkj99nE2YSFVrSTNYb8JCEyuGJFNB/z0N6fn1dw7kNfuvAXbSQheXC4A
rS7q9nn5i8L/q4vimDVb1fTbNAU4QpVSSDjZE4JMpGeBmkY4ymL9Y5vvtJzcjZ7i
DGMARGXwFOkjedDPselOjS34+pACHmQ0n/ZYCGU98teR+4WaDl6tD22sgZbIp/o8
F0Yujx5cijr7u4/+oMZPhqedB5uAhEkMIdlAjFnmG0kkoZmGeoo6RvFZ6DRVs5x8
zE1HEQ2Xp/vr1qRW5nR+rb+QxwA7ZIxND6Yf3FeAeaBMPpAI8i4PgIxoE7uN4yye
v/8jAH9rglreNykPRfu86RcbqXf7iYSC3kZgEk78bGIGYDQFHxjVOgLQS/idfN10
966BRLkNLddl75SLWLVV9S/14GR/WnwIWJnRWVEMhMqSytAgsHkWsciaOjqzsq4u
fD1JaUB3LbY5AR3U9sjK4Rf3k9dSLei2iNwoyCm3r862LC80i6apbIdwBbQ2bmov
1SLT7/uA3yMweNGFvhf0f3X0rwbUU7nDJf8z2MMl5PHzFUL/bbQ43/9qwSEuX0CW
hZnuGazOK2ljwpgSIrZZmLS0Fyv5+igNntMrGTAvUVSstNFba3nWexgJRe9GOqEO
0Uw/MBPBPnRt4dti9vmaZxkWYDImndfK6mjvrATt1gPPdPCU6+VN9wrF6zyUp9s5
6F2RK66I2DROvx8jAAvh38OlqTiUECYPubldHDqEGv/DGfaqIYueBJM6VAE2ZnZm
UaSjG9hddKmKvcL0rwTYTjFwN8OMVejF0cXhIgRrYGI5/sKoO5G77czm6bA8yQSN
X2s9bZaze1SDEQVx5DEQHvJPmt/HIqLgsFr3jqfItr1OMVyHub5D4gkMW3KsYbqg
3RdibnFg43ecQddZGSbzaGABEe7atqIr2NA1wFlFpC2QOKFkBZde2BaCM27jlpAo
/+QFIn2kEQ4zERUKTV+z0IZHbwBQz+eIz2hjvI2CqfM3G8LtdCzYDULqFsFmiKm7
ZT4cShDZwmFzkPAmxh5TmonRaX3jIgQNcnqE2LL7IN25g6PHo9xTxEWWvdWnrzwX
NaM+GL9gPGN/ieSdClEAGClWVYIe/73L5Uv6ZgBxkhubFB1JyBLYtalCK8Zw/NZQ
mBv4RInlT89XMy9e3gB5p13Rwowcr9C6iGBaazmfOlChzidfkbKb5oIDL6/paHio
TicdF+AezRsZAe6G5cIJ0jEAE+156Ei4Vz720Nj7qb0XcP5n0I3OFCF+R5xHQl5X
jCHzDlDQYiPAiF+RwBQOrn+sGt4STDYlw8L7geMAEUVsJGvj1mRmY2S0Tkn9VF4i
7uho+8WFE9SVskmeH/eysCwHLoA4L7E7WZ+Z6srpeLHN9eD4TiAStrRStUctFCBH
A6vbi1X3uzeH6djAljaMV7JEMLAM+8TGMbv7yngy4Jj0a8PV6kp6RVGeSmvs9FMo
XTH28VGU6FCglLZhcz7ZCUBfgz9rqjV7/TwfKCI3WEHtmOFj1wq1UruH6kf573lO
vf/jo0mN1W3+x+A05rGYZ52ujNC/8StdjEqhmFp+nW/HEnb1+oYwmTcMpdSqoW74
Kaf8/mSGGIxrnLp9sG86T+DQ+0TCZM4TsXi2heNbcx7eCkNgxMzMpDnM3ycIDsvL
X3TeFUfgjQhhBI5tX9unFxYnVGaqhL9DQ3oqQtbyu3CxKD/xqp13HLrMRNEGJfWE
8Y2JJf6mP0n/AR7Mc3LF3bCXUuGojAT+0faxIPqRhUtWdfM6jTZh21cY+22Qdwew
RMcWGyXNlt8czShaWcmSlMhEJE7gf8JVg1Phuwrl1Dcsqs8uEYJAY9veQU69rPt6
OhD8s9b2F259pqdRzhG1hGRLj9Mmm/pcMUiaCb8PG3BntWTXtockIhj51E/5mwIF
7oHuNigQvYriKQAMPCcxRTFgTHBfeHZRDqOD36cPJ2leoCVx8IUkWMTv7FCYChAj
+zk4doZgE7mzs6CZcafdEkaUB3+WxD41MNC1L+foRj/KLmKP1YorXeuUZ5DWR4zZ
59+BHM+p0FaMKPuYdmPP1S2G6+zTqn3trELuDXHtDI346diXonu4jgAhDUEajb9S
GK25yxhhbG8AFRRfLz4dw9tvak6XROv+ntBFVnUtmGIp3qu3MjLB3ggutECAXtFc
tJZY6GnlmOhUd+7d67C16kZcUHlxa6Q3xqHujbenyAU4FiN2RQ3KK44dBax6/60D
xrcOH1LxvJmB6EL370tR+dCMwSrK7lEuMxmksKTyQg81WFO2x9U0bbOPL6pK3s7K
TC66WTN6DADFIXz51vuPGwS2TqNnc/qAk9wFsWf1qN2gXhZSmfOnkERD/XKCOpA3
BwuCpvJsFeUKAAauH3tt/+LWHBlWOgCamKuw/D8I6FF0s1LmBTE2jTM5QsKb531I
Vt9zVj39xty3ORNNnzPMP4tj9WloxlU6rasi9KWP/HcVuvoe1g/2KaUDsOx82twc
jAJVrfExLju9TZz1NksktYjsh3MkkAl+hKA3WPaR1Dos9ceCEyKpLheqpaSTLaxa
gdmcjHM8h5SwO6uqaY8/OnfX2CWWHplw0ZmuMYxGTVvGvfyLVXw5rmmlpLqA+j0E
0wwY6mJH6KcjnXl8vCijkAVIw4EHJjoH/XfGBEKGbOXkhYVKIRNABs3KeYQ8Ok4V
zrNVDxC+Zq9rjDn+UNpns4R5YAy+9QtUuloWpljPFiWXwzjxKTFpffhSkdG8CIqM
JKhGjlgHwYHPYdFjsi2xvwH8hO1T4WNFalHME8krpgEQSg4nb/kONQSPPnIEk45l
6AML2OM+qrTeYsVomNT1jQx3+01bVd9ci6AEPCothWWDp3GgwQCIhFeyTczowsHb
acqXBlrh+qWMk215B0WW5uRI+ICvGTHXeR7IFHV/rRfTyF916RcIq49bRhvE38wp
HkIcnkctQArx5pPYvStVpgn4/QmiTlalv4jPoTUMNhOujep3O/7sPfpRPY9ucVXt
KUqCr7Z0BLeCPndedKKQ05N3V/+/A9DkPIh3uJtxChcesTIY0IXipav024m4Qang
uA2XNFoJnFvON03fnrLGLEDMImYurEWxexw/9dy9Z1xXpCFfdE+2C0PEQi7rmmOE
iShQE3XFogkQx1cqaP2rhjoMjBO6GElyJayVUZWw4JBhnYKo7ANDMl5Ca2/hAwfN
vola/6YhgLxNFNXn4OzWjqW2KC+oEjpUhwHhr2uBuCZ70UKce+EPY5Pb5zDim/HI
vhFoyiivL9LT8Jj6LmFe99YVeW/+L07wPoY7RznnuvFqsM2JrWf1GAnl5srG/ram
eZQZQfGebUeIRWYJozbn/BFv3ybo+e/zwGKEIRa2aLEwb7UmeDHSah8ETmarAJvU
AXHYw5Z8RaQby5kmKkI9p83F4qaCzH++VbR15oYyD7mtQnSZDMAif+MpcvxWeXtt
jATaNcgcwPrRDpTkptvnZ/pt1tsQR6ixwlBwfM4eMh7z9S/Cyi9LZTvLennq8ICt
R9bnazwPNmVJYRipQsqm4xYRdlw1T80wvbv0Drkn9DRcq9grZtcBDKpn4YTKvrly
LVFmEvz+MYifXy4AkslkuKtybdNA30zXswXL1MV9SYsAZXHDxBBklKSUn+3eD2RU
muK5xz8ea0fUOpEaTrMfeVHjatFIuYbnLqn75kZHQeijjRA2QS7Ey42VA9M9WlJH
2uP3+Lo6jU9NFEdR3bjyvbvCcWBYIfJXzdTBY23Tn+3wnXZvpmyn1o5IX3w/yVNm
vOAKZR4eknBbcgEBU5P/n83axJvBHlP0f6AHZHap2CCoGOhnRkvsJ6IUaBftT/mR
ODd2jiYR83NKfuykuTFVx4upA+8lb/hNXPxJavwrDKtTLyq+x241wMKv6D0QuSsr
V1pI74hcYlamUtozEZCPbgPr7+bFa02Hxa6RCofvpuH/iKK8QGWm5pl2bGHyyjlJ
ByGhueSTplaDUsJxt7NdAZqf31Y7ood42KMrx3+QddLlahBLPMszXYgeD2IOm10H
qoP/0E4munFmSXCSmGdVxR/UTdTJIep/b7oKKvpfnKoqoMJ/Nn/2J8p+7Nj6Ep9L
glPU2oyeEpnFZUtXh7lsq4aV0Qw/RV5i49sqlGTQ2Wh9Au/APiBkgwDpFQpGZ6AW
dBH1ZrpxSC8PKIcP8yp45DL0WtaYLqNBqSiuSf3r13EuMm+nfXydXp14Xkhy98Hh
r9tm3hozYBpFqCaQ6sG8XjYiOgJzIGcKrHCLk8hljO6/fiDYGJmgFBUHksl+B/JB
n+UVS6eV6Vw/ZOTmyPDy9tDKVmHbzqViUHKCSLk7BzFQLDqa30on86iQ1kqgDOSm
Z4T6EFDI0srvsXtO2fq/fyxWMmNc8c32MxhdDn0u4WSac6Uj746YOwdeSkl1ley+
bmKpSpIyLsiAJ/Qx018i/kPD1RAFdr+H7uF0lAQuWdrecWDAUfRuScoYprnGGauo
5L1AwLIr5O2SWLvRmMwADgOFpiLu5pknh3r1Dt/5kguHGEYjN5cZZ2nv/9EQufgh
v3MDw959jifoxyBqNi1de+N/CLCcExNePXplMjS2JqNLOgp6suPtxkCmIU38KwHj
mbxYzVtV+1owNvfryInwV6SuS9ugLAh+BC0Ogirt0l3ljiR6bErbftCqaVk0kOJE
A2ZCyEmne/GO/MptscaS7TIjQjFeKCwQbqPw+NbQv8AWkHGWLQXE9PxYgDaPDP93
fWrUR6aHcHZ9+qqJqR7Mu0QQNgYHL/4J4QvJM7rOn0GVw9pmqEUgWbRVKfOvHejk
T0sAsRGmxAAxMzECEqGoSlHNGiVQ9zTnOeYaYIumfvuumokO3DPWLVE4Msz/ePK8
Qn8s6aXTndkSSgYwwvSPkwrA+jkQC8vemJCBPuF1XUZvpTH6B7nbK3iXcHt4IXZ0
VAoAiIFgp6wbT14x7qlT6w2+U5kxu4+ZJZ95SVjupnAHHOb3IuPssqOpI4Xv/KjV
7DRIUbO+t449vakf5O+oIsQ2eJADfUUUqOoo9LF1PSj9aidpWqJYPkRGMDArUOe1
t6nMOyEX/5ArpRBNsYyVvxa+mZacKOYkN+AFbkHXZAjBrvf68f+o2J1gv1sQav7E
3SwoeHvN071g2JyslFyX9jHZp7+ITVbiXOH0yHa377THp7e99Zix25ze1Dahy+jO
SdSaptn4jirepo5T9pGDBRSr4zYHme4axHBYK8N3rX9DQzxdWle227J8HUnxkwxE
VEio48YUOxIXQ4jIblJrZ8BB/3ZrvBkT93pSrc6umsXKMe8NwMA44EMdByydyXje
SIM9hT2xK02TPYyT9pyiVVcAxngR4s8CLNkhG6+24kculYNiTBkFbZ/VVzQphBqg
omnavUYXKdYR8DNZPZcKJpF4ca2X9YakE88MBzCbfpfdTNizmjr23agrbwSjJ3Df
lTINe3ljAq2sNESyprvFxXB6YWM90/w87PKcZtOvqwiFSY1FSUNh5xx2JGGX5GLe
97Vo92T7jkgRy1BNuQaMLYvR701VF6WIV3N+S0z+X4tFTGiAFJcHJSrANJuYy9VG
VMN/QvGwqkqIc0qkt1Wcy5No+HddGI7BQK/Yj1olr1MRphu4in4f7NEUxWx9jSxp
U/CjicnMreCcVGmi5COnoNDMjz8YIKcX9MlYVrnJLmWTIUTX4nGUQFZtesfAYsMl
kUGWApJBD5qNP4fJem5qPs5+SPLfDCwZTqFMbB7gLD1f0x7RU01BHjxfVGaJH0K2
ggEZ9/robek7Kd+cMW31Ar5ZSUIE7fkbW4+9BX1sBDFj8ZDVpVQWZEh/9QmMnMfO
S+7nXCo5MEjWgv1SL/SOl+jzRXMz67OB2uhgkIwi9C2IC34npCHafq8qF/Tfe4ox
5L4Ep6m7xIAof+975qEYb+5Za+ZKp58V8gfgiqoXAUWBLL3r0rEt34R1M74ZGRZJ
gr0GeTmtS8T13PqUqPc/sPNIO/ut8u+ZXGulcVZxBltCfm+KWmniXmrncWv4lWTh
NZoov3NWeddNKAvyE2ox7hzRtBwVUcrlm0V2ktTA5WWB7O7kvbh0qLDrKtkk48Z4
iL+8xJzTZMn9Y2xs2UkKgGZqqZ3IO9Dpft0jdLUrnjjgpE+47eW8ZvurqV1Viyae
ZptCBryqlnMgXdoALNSWNlJcPQInoW7UacZ4PE3z8fI7ypPsJN78urz1OJW53U1A
R2c1iDgY0dE6b3xp+5rw1pEryNn39WmrkTHNeOJyMz/Z7FyzSl+6AZNhwXjn/5Rm
K05xW//478cbqjmb2IL/HSAMky+3F6Di/kMNPVCA1m46NgycuDBm2KJzJ3MRtThc
HPa2Yuo7g/h68+RAlg27MhiTwyTQxV1EK7898zgP/O4OxfS1wHY2LZEMKVUHfjnQ
0NhapMeMogfAMItACRnt/NgEbF5zSQfObBLepKC9GXVyg0/61NmZoizuTuRkyHvo
4CHYi/jAJICe4w1HScHybiZJeOHyuSdwFKKE2uhhFNzp58AtsvJgeSle2JrX7Iwu
TxPqQBoJFHK9jNMjrGdoI0W43T2iTOaojZvw7kA8JWfFM1BDi3H13fOPLgOdwhxe
kbkeaUOPgOPq3vzPnvHPmOgyuIhmyXM7wWknfHs0lSR58M07Brge1g3hhlynsJwZ
3JPkBZIeIVIcku7sFERA+LyOl/usYEvRnnBV01Vhklr1zIxheTRWuEFswBh6lhw0
Py1duF19Scuy8AwkU96Pgnq9op1/RkvqhPIuaWs2sKiOjOar7wb6uJa2P1cgMgIs
wDAPLcA7+SGHpjsxYg3EWDwAxa7ySd3kObRtS2xewgb6sk6aT8bOCrX38rTTFACn
Yd9lad0zU0pQh4uMHq449iiRoxHRKpTkVlam7F2jNM6IfCeJLLkHgPxvs7QvkYpp
FDWAYh1gwQIYhIvsSq94ItrPYA0VCrF2TX/k0NujtjWGfh0Wk65qkbzZX0bhpWzg
huini5g6pB+9jVRf/eAZs+0NmYfaUE0oN0k0Ljx6T8NjI/+N27OahdLBxejm9/3p
X7tBUxgwwxrzZGMVNwR4KJeBVlLYvUso0Zc1eJS2P9zacYZ/Hla/2/IiPPMb9hLA
iXa0fxtxUgAwA+hzbASj1l09U8t0hrU/UiEri1NDwXHQJ9bkYHadk4ul/lglVAg7
mIUyZjHi3+q6h7L4cPR0fN/vxzVZsuWzCoEXen9Ur3oIAyUKXC4jp5c9CCbgZGiB
WYHGm62liMMufnm+5ak05U7/+MSa0cXgfQIK3J6QbRf5uMWpOWOf2sAt8zU3rGGk
Sy7KBEVbaRBbc99eNEJmmiy1aF4TkYMBgDobimbSgnEW6KL6cxY8Hg5JDxGMC6c3
LbTZSnPv5P47Qjhwfd5yoFJIotrYyDDUQPamgI/3NP5iCGoxs3N0CH9GI+mJ+ELJ
6yl0ZS+a8P0ljxWTMcIRVUFKycLwgCCwob3lyqGgFcalx587g71syYCUq4NQi/ij
e1iEO+FUPF/tufbBVMQA9KhAofADhTLNzCtJsKB3QGk6xxm4LyKWrjrgkNTxmdej
TtSdaw+MdYMogx2zXzIG9BGkoXDJfaHSkAmzxL+Jp8Rm9TZ3zV0T130TMu4vS/3b
qe9eDNBfyOtrr60H3ISqvyBVao5bn6A0CFG/e2a0EYoY1GUABjrWsd+GCKHxheOz
nSGWBsmd0WobICWWYOMNwDjHYnDftuQcJ02WJbTY1DjTPY4S8BFQFECX8XLRmjc7
F2um2+G8zMnNq5+PPx0kC195K0vTSPYNYCF3lRfLbulPA3K32jj8hNZeJB1vjdhf
mlV3AfzmP/gvsTsXsZXG7gPrKc/56Sf0Xt41n7AfvWf69U7PSU6f0ozQ+HOYffMF
QMCbFVwqXqt3VlT/TRdZIK0peFZgBG61a6FEyyMvAngmFasLT9bZi5vVNVSgMAO8
54bhB43SawFRoaC/K3uByabFhesh2RalZU8PFOhWwoUoKP4ncE9LqOQVQe3z6+Ll
FjJ7nYJT+0XtE2jvZRf7izZZLOUeypJy2pNHpkMyoeREU0PURysmKFTTnsm9B4I1
gvUtQnv070+9qhUdvWjMdNWjP2Pu8WaYg936VjLdVMuez2O67SDqWjulvcAesU4a
WRilFG/8sAGneo5WoFrAKBvE4zgDFDQZme89+yXqxWu3eFeAkt1709fqh1xCvckO
0pMmmaf3qnwEfYyOOLw2RCvy5ucWYZwTUJydQ1jVEtT+LKmis6taHCZaaXOMZIx8
OjaM986PKg52KMursUwMlSaLSIpOoT2oso2fvaeorcLxYNvwCUMMrQHowvyuDODN
UGsyeDW8UlnPSSz7tugW8D2skONcP/5PihG87ZLwz7GQSsOm5VqSgBI3QHSvSLyq
hED1B6lVhPdxbOdXfZ2SMslbQRJvfSdPzQAobMYjg+HxaOBLaJPCEeg1g73GsY3w
KAPWxpIJ/9yTARybuX+c4YPp1Fcx2AxRE997mnxQf2e2Gb4NWWav7Ekk21X9UmuB
7rP3JgccenffF9BBLFQdAYQvcnXvMfSt47X7VlsQQEXjPNYUfk+vaP03SfpCSigN
sdKLG8CXY3TfAUrdMApKT9Gsf/I8LB3Be1FCX5lPscI4/02AOvdVWXDZx+kcnM0M
pZ6sxNsPI74Sz9Gu9mhrwxxh31FUMZBS3pYX53e4Fl3ox80yP1dQol2NUDyX7alA
e1kycATFn0D4oxbsnm9Czuz819JL7N4VP9lL3JjsgrZfkTsHgl7F3vUv45/brYGD
c7iPW5BC0X2DiMJxryJu5qZdoYLe26PY5swYW7ODdTsGXE5lPAPKZZxET0CNNnUF
MJPPzcP9biMNDPVpllS4OD3F+KmHVnepaphcaIWBdWaqQbfPi0l+MnQOm9DQwCsl
+LJkLQrmAxJo1ftOov6fHhFLQArR07uuxndTZjupP1QHRymOgIZcGBgMfHuBQIkj
SljvI/gZk/b0tvkp55jlyM3L8eyZkpe0FEt0ZlcvQ7fQ1Mj8daFbOxabOhDmqjoA
Q1iqpcM5pPbzNCc7/PgSpm3iZIvkpg8hGcA2UTIj9i9x4OT/kGAq11t1OB9w/pa0
oT5v/ybSk6mnLFD4qQefBx3u/VQu2DD9g3H1ttu6bwS/uMUS8pYG2RBRt1Bf28gQ
Y80wqbZ3oFEJkYeYH3Bu0z9BxYQmy45dIYAOg7wUPJ+a9/iVhSl5d3EjSIDvKzP2
3nus7ZeDxm/JVdBj7KXUg/wqzWO0NQH9zaKHQ35CZcJzs39bvXT4oAOxzlUVPHxk
WQrJ1Jt6zIIkJIh9nG6Eju2R0DwVJzsywxc7Y8bn1M8vjhjwB6Qtu5EpmiE6D6qD
rZV6YnkdVXG3RdmU8W/gh1eFVx1u6Id2z2XtfiNED8EUR8ncs3X5+DchLTp70DOp
XiuRVZA+iLU99eQ2kl/8rhAd8QW6Eb3+ZtEGblRb7xtkqUDPw5ub5c92kg54Xzo1
LSvBRVO/WYLmthWOePIn7RodzTUXJ5spu2yBuo6d64CKRnHjqcaC1aw0vRD/L5Qe
bikpgQAyOxJUTCJaMafhDQlHWZ9MnrsgkcD20aGDylxQq07i0dnw6DIttC+odre/
zK9RmPVWU4AytxwBGRMk8UG5YjmlK429k+nJLikGjHLJMx+MPt1DxpVKHwCozv/x
9g+EJzq5+4PND35OZs+cXRyHqw01g6Twz31ukhYI8U9q+zbfbJ0r46agzggF2rHi
z2l49YdsMH6+4jYRcmrn1GGWUgqUz7boc01+iUafGZW9H1zgmd0EjGY9fkjHKUSD
0rX5HdMK4q9Mmk+x7TEgENxDsJ+ZC3tu/QASHrzygSMhCV83rnGsv1RUmDJtTcO8
gZ7UVXrVUZi92DgLCvYpZjBvtR4NAv+61uRunUfMNj7wyG8i6R0FcYapkF9KoRlv
iCSIBH3JOSAyVNK/yCprqxP7uZ2lhe1Xwk6USoHlLP+LVXRsqtB9yaruo+wsZ3SB
ESqOkL33Vw8b2WXD6Wu6r+kxRZd+dT241bqDSNcINC2xZJeVBghawJ+LuGo0o4in
+2bsLeu31fko3O4yc9jaF6bYsLPX8MSdwLbpeI+U3+qD4Oa/qJKCdJW5sTp2D1Op
RqmCsbcw41hcsEWfos4dVzAy8Yu69xJU3toMTCTJMfESavyofiNiunZTLjazfmK+
KtLo3AK5RGJJvZxe0cBPI8a+djgECykZswTZJKpxKcletS8NKPK4mdN/TTValPlG
zq/mpIeS158D2fhXti64YdcIg14VBXIcDt/0se4Ct0J7zdja3hLSBTqORhFBSX3K
YVxZKJICElDCmYkv5puwCyp52uRfUNRlp1fp+Grcocb11ONbyfOTTSX6VWRI38hR
pglGEqlYl2XmIJ9lt5HgrDcWbp6vam4jE+GDZMWY8lcxcfti/+gErDx1N3Q0eiEZ
hhwciFABsxXoKoeovQEkPZMelWjguFhXut/dAZu1KY9KaIjvWrkrdKQFlEvXdsT4
GnP3FUvfTJJxO6ceO9OxCtzfFvt9DqJCbv5IXortvJIbXUg87ZzCMmvaPmvOtrxg
A4I7ggmgzqFs1wcriR38cmRPK+CUHLXtDShnbYiNdC1lOoNkY8M7pB/FFVtpziia
PMd2AGGjwVQXckBoJA6W/x1QMj1eFdDyZ2zFQMGUgdAKP+REKZK5zdh352yNf5Zx
GYHLyU6EMtON8KVLWrBxFx2LZAbr4DKTxSnmko6QtUqyyJYvpAVSjY135UgBVmiC
kNyGrfcNWMxU83fivATazZOGEkB5CsbkT0ty156C8vXcObD8uRpPdR/sjydy2L0v
ZgfE+xW1h321LahuaKHCXg8vGV7r2iqH6OMNzKBEwI7eyVSE988tKXZ9VRyG6K9i
fX8Wg21w8bePus99BJe4+rFK2/mmAmcibIDuzZXvqpLTu7ALWv863ylbjhXvi5w+
z5FCeTnH9wkHa3+FcF+85GpSM3uu8ZphjTyzEGvszwVKr3e7DJj8fNvY+4PlNZBS
rmXJpYgH5IW9+5j9C2KI4RmzCjeLLEuPIore00oqIwYSqE2fuX2UJUhYm5ena0dk
oXFlItyA9Vhh2+6rrgxgqz7A4AHCzU2MqJfGRXB/JPc6c4kXU6+EhyFVkwneyDu8
09/85Lxr5wFfMa5JIRsd6vFrR+BE50n1ubC6VKrgQpnG/tD/tc/7kCG2F9+JOzfA
iGtvdiRZ7bSjgXj+Lfdo2fPxKFakzhlSOFWaZY43Z5EoqHjpJ61AKk39XJDz0RG+
C6yAXmKuT9sNh7MbTc9dngckUnqzg113aZx+RKKrJG0yk3tYZdaepi89DpZdlvsI
6RWcbfuNFKrufFWHWEz/5ltNmjZ1Kvukh9srWw67EY3TXtkamEJ2HxvOFVxyrh1w
l/Ok2OewkdlSUrVYhaocannRThvr8gF55u0oCECn/UGSjB2FNVQBDz4+6U6jbSIg
3Jo8u4ClknJNORvHsAYLmx1VkBpZjPHvwr8MAZje0C/LeH4gYM4h3aCMCqMPeC5k
geaK5FNOh5DEfKtaUDoIDYZTQBFMMjX+O+O0b2pOktZZSY2K8CfhcJSqcldkoIlU
YKp6gI1J9nLSREMvnsYo+DZRoBTJjs7PwoHvhYt1nL+XKo55NLkI7QO9O2/2ouy2
Q2uif+93rlrDebAv8UJ253acer12V/eR5y6jV3IXOBASqAHYtsSJtZapVu7afqEX
h30n0q1vEnsCaNSVLqM96HLJO7iJO4WTbW4AIrbOK1Wtcva9qKVsUNB46YQLOI+d
ZNpu5AFyH8C+1RpNVMSgPcubmSDBKYhG+RNIuTvuidaQ3aPgCjWYL+x/gbURTPCH
BNF7/U8xIYaTHttODZtd/fTlKXXrndrFNM1MLhBjn89VI5+AfkcdjbUFzY51upyf
xbuA8Z+vOlsp1sij/YnvqzOzONuJK1GHh1De3FCq0wlwaC8C6cDXFr1K/Wd9RzBX
yp9YztIf4osCIIedKGRpK/O373VzHLvmmSPhz6NxkBUps67j3g9cR3+WMoV2qdF6
Fc99hr+km9vKPcQTYedn06ISNipKmnel5LQo3GI2f/EHO8LeYRZrT9gK7pZUv/87
dFdT4vyECdaPcjvfyGy9BNWJZUaWgj7/KE2ptf35tq+AYCGdGPprt2QmcuXdF/oo
xksMsxjipbr5qBaJ63vdrbKG7zeO1lio+yWZizEoZ/lYkqti6dk86Nw+LwNkytud
e8WhnSoqoTNmV6eFDwjHIhpKsIBbMozF+rmzNvyS1FVMk93RqNF18ZU+bxwQ2z/F
+v+08n77f71sQCSGgjWu2PA5ZTqYL7XB8UBURrp6WHDxJ3wj74KbAu7h7IjPEA37
/Ltj3Z7zYNM4TlajiMLCdQDU04x3cVEFyT87WVWELHoITynA7ZEAnsRsr3Osrs7u
jlcm052ezEjtJohsslyX8AJSdewyzRnWFrNQX34rKEihCKcuMjWm5lAzq8mCTQth
ooMarnj5iB7hTYdT4c71zFxdpooeKAcL0Vi5YBp7AoT+xR1M5MYId49knRTaxtR1
UBqRfrgTHOvehlrVKepneMk7ljePTMSpiWi59CtyGBOOcS7kui/b5y3C0Pdc6a4G
+DS5dm08PgSECxll7QjQ0fIH8UjcePfI8NrIkgTuPagLyDo6l1L2QRthtACD+kr1
uhMueiw+/M1TBliM5yqNna7AsHa3yjrwATLXFUmXUISDIfkSTKUgU3A3DPiKrlHY
6wAV/yESce/Azzu0Vg2PSoJs0/vOrmpRChQol5IibuP9o2FNT0VPoDg/slXz3Wk8
DbM6bdQc+rotQgEEt1FZWw+to9KGEGJ+ziw0D32ZWgPQU1gRIoyt+jWlWrfpB6x+
SjWfqDouY6Xp+LeyInMKVfeW22PrvRkUwmN6Rq9DT6cXY+OFinpTqRfw/agpSRTX
t+Wb06er/AucOXG/N/7orwJwCunK6lVA8CR5E4nxFhHORsMNE/O0yWAKzpQFH4lC
SQ5YO1wNyNYedj5qaH0o3PHJs7XQOrd520C8TvFaewBkvYbxNx7MMShoTNiS0Tiz
1h0fsue33qA5Rr94BCMXYzunhPgi++yM6yL3H3k3j39Yxdvljwr19MLYKFl6iOXv
Eblc1qzn7/u4y1EGLuW7zEm0u/Pz4VT//GvafS9qu8AnHGQEK9TCF1Y85pGeTXvK
w/ZRTZ/cFGyQ2Pkhh2sU5iXkTiXKAV7h0FlIGPWoZUdz5JBqU62Xy4eYv9wUpNOH
hxDXdZ+M949FrkJKnRJKPXl/BHuPeX1kX7gNDBr5wndvjw3uXpAiluRe6kSYkDGF
uEgmmi6KE7D3VFpMWHiF5JHiMrezsVdMlq48UJVKrL29GsP5uM7+cMUN2Hu2qYe7
LC0XcdchSaeFxTtWzFN/eLH5XCji4fMBs3VPzh39Ai5nfoCEjFpfA09dL2ztTuJu
ZBDndm0Fiman1DH4Amx5MaK2mqpPet4UIQqIbBXvnWlxAvYQDL58lrU+v7OEdkYu
KXUDzzih+E0Tq8stnaXtJEODRIWPvZOuBiphc4G/rAmZRMMXaDWjA2i8NTnG9nUK
ZsorUIiWGI+T9QNhho/ktviE4EKaVGffRmPu7a82vu9NULuWpb7Yl8XN+px6WAWP
LXmcpq9JiyulS2q35rO2g98xdaZPlQTnnasV8Pu2c53bmyzgmQjsr0SNojnCgYlZ
o4ukqW4rI3w/GIV5P12pONcvGvQScqK7zrrwtdOht7mjmZEFXtXvpPabHnKGyGFd
PlpRzuOLL70xEV6CSLrH5b3YwX4TtwTzMZoZbUoRscOzj9TohxT3n1+QlgdcObSV
8MDiSQ1oe2wKz6i23zYVDzwn6mi9z1lrgbOTGluRaFa4+fBbYtDv6aRO52SJDuoC
FTIo4ud5lzt6teM9sLNJhdfWSjr6qQihh0eDI7pHG+bn+vNgnxHzNSQJ84oRaHlW
ySSRbsYKBW8RMupfSiO29HLCr/pWVbEMhvkIH7MH6lSX7GETZ9w+FAEoHc351xse
cfpNLpxXOS3KhiQIBbZCYstfNE6ChCGjbSdKNzJFt/Eb+o2VlMUnDASj7qgR9cZh
Az6lK3W8WZHYlYbdIPpwHaLSMjLIrgRNs58Y/dFwk43pjCvdAh0pcysof28sRdjB
6Tu/IY1g4e8RFP2q/dFm2cWskik1ceEL99z3TbphC6Y/cK4hmzOxnf6K8kBGaDec
PKCzjNY3NxAqiz4A+oPdv/11f/UYhokSTnbQt43+SNkMwC1V1NCT3v2BcPhTa7BE
m3itTkwySI5tGzo540gXdx52LITyuDtIA7MH+hGf4urWPMf87V5Aap2tuH3Jz7+t
WPqzVIJrsHxNSmz7aaucQXtA1cWjEnXy3YkzfD6+AOSxWBXQogVMr7Sq/V3N6+La
2UgL5wuBtYaCrs3xLv7xdsX79frcJUvtN12nyobK9hXqt+ErKcRqGqmcmHLHZkmc
7zua8vLVdFemqSG/R6uWYgNaO7HukSos1sVkPZdMS5rKVLXsQ4I8unwtHBZsBQ/e
5vfn4SY/DFQTun87pq6ieb4+Ir219wImxsmGRnS+njQfOJTEkHvqFXqNq9RX3fI7
LqVyJWsLCwdKOYb+Fc5xraQEadalWg8XeWkn+hfsft40C6k1pWrbPMKIW+LS+I5m
AgjASKOIo+72cKC59T9uaCVn3CJP6tMkQFhJ7RuGBhT5GHT7/JSFcCX9D72T2feZ
RHF1AJ6rMlFQGsPnwrKC/0FC1YsTUswahosEfgoMES6TJwLwUGVWFQqvaFlSKDFv
c7pNqrtgVZPpU4lPtAMsGdlyx1LZQFT+ggs6BuJySS5pMtuagAZ0f24lSaSbZ/K2
OfUakByyQ7w3Fxd53fqU7pqqXE9ZrS+hMejIb5K8QbCDT0aCzBQACwLPFrrYyVWL
0D/Bzt46tG8iIJd1a1NaOabOlY+x8uvGy5CC70NY/NtCiDJQLrEoaJaMg55VgF+7
a6lAHIznCUkvjawbeCTWmynkc7nsKGcjWJQEd3YR09QzfU1I9pWvVx02OSAWxsmL
i+awqxw0JLvylKxQLCt7+YVrJErYiEuwOf79sKcK54g81BDbEGOJE8UxQL9R+4/w
WmDptJtQpG6NiYo+tRs1NFrvn2QPs9ph7k5EU+lmYr5qiczPEmvUinP0zeg6Pg/q
reJaL1xZp1WXaat97/i/VSdCx2+pjU6n8Nf58VUaPc2Tpl1tyec5jofx2rLuam3f
ZlKjKp+Dik8jeY7IqeKE7YG2a2YPbAM1V5IdXVT/nbipGcQMNnPELiA0xTrkfILs
XPJ8hnIx2QBzotNHvqyVuPrTNzrgOIQFS+SiKvD+Ovd19MGlGPHtp454jx4tVW41
EeIDtJwOqVwH4UAxcKlt3y73HQ3PGYV3ggrWVnwgDD4EhXlROUSa74s3n/tVDHej
XhJlooru2v4LYZ9lkDLrcoa6gcUH0dfBK/m2vdj9JfqFuj7+6ulIRcV6dfPNYZUP
+AWHJkBPl3sWa89Ug/mBAnuVWJTuV17+rfovJ3Df2AMm4UYcPScDzlM9MANgSLuI
CO975/MDiHPvL+A+7lbsiL0nHiy8kfV9xuUtztev0I2iiMVAg2OLjq1P7Mi4693h
iW0nQZCEOoektRiNvk2sEIEcQNZLP+Dq69MM1dzteoO+pvE1r0B2G0q0bkcnxxZ0
hVr0amDqz/Xs0YO7khBN7buUP9Ol/Cx2U8bl3mnkFhjoGSg1GvEuA8GHE9B7M1Ys
gDu9bRZQ+Ryg5QERiU7Fn4uE/dZtjYfhiePn7w0XQWuqfSLadV7l3aZHVkf8I/4v
iGXp/gECiKnWHbC3PHO4tc38Y6e8gJ58+PegWdqsY/+f9Ys0a/XqnuBkqQzJXFMq
d//tIK72/2TwArcgrZZ42W1jM6eCFyBRvZY8/GSW1hhhnc9fkvNUKwmOxY7ownpC
Z735sf+DYR9zf1Qn2cl9D36PVVmCh8tyK4dEx0Dna0uQOPl4jBepTcV5L7ntQXDc
CQsIZEDcsE75FWVSR6Afi8WRxdTLXrghO8jmE83SX0ejoqFi7iGqe02t3O2DKi5x
+SgRiFfqpgshSdM15mPVRH3hC+h28ff+SrSVXmiV67WIeUGdRyhoFe422o5bRYgi
UEOMzuXCOUx8o/BlsXVoLv37MpxwdfR3bSJc2A+utlo2eLp6r/VMYbUPP4AS8ad9
98kGiaYEhpfDIzg9BayMdugjPcScstlenk3k9TFHbvxUV5LrgJbu3vXcwLtiKxHi
K/UJKk2Chp4FfxAagaMNiM4ZSSGDnrXVr1ve/hCWm+6jbLZ/WNXvouJGyfX6vNJ2
mzs5KFDbN8lY+4MFlXN0RQ+PeWePFLGo9KHmKp+E+VCC5NpXW3XQ2/iXi7SZuNra
ngFywtt6AXPWVxmWH1fybczgV/6lhbLRyz6gcdH+AEcRmtuG5zKY5DQVpQdgUf40
Q6GVNB5IQQuUekA6B7LZvCLA3cCJ8VwqVCzvUdRH3dPNwRlhzTZ4E4/kTLjRVpB5
nrpk2CVa+XvTQPnIPyRWvQC0orYeXYNlE+FleKnDd+tnOF4WsL8BQ/FzS2W8mWkJ
1vSIWfu4cc+qPa01F/ceKmQAnfxCWyppNPEyQ1KU06Al9i3qh1PJD226DIJwzFYO
dPPo1k3ApVVenS4swUdt4Hzwc1QDxw0GapI/mc+3vx6+GSds/fvpyc3y3WpsJXLQ
d75Z8DkDTIB977g9RtzbxHR9r4ter1owhju1Pnpt0v5laI7cAjAE2LW3BonENRQ0
SNB1kdTK+qy/DBd/oGwE5BO8WCp5EtrzOHL4LH3N30Ey+JvqfKy3v1w1NMhjjINb
zw2aobjCSdQFEbnreP2l6sgrJB63ql6mStEutTCa+Umtw9FhLdDvq5v+YQVov58x
VKzU7t7OYkSfMl+E200xDg9KKfHhiznUfNLiD1veLuC6n+RjE407L4VkBboLsztx
Uvkedvsfxxz2BAxDOxw3xwKABs71HqxqVJx1j8Jm116yXjrZtSg9guSuk5XocLk0
u8afZiY/2r9OnmzvC88gKmFl5fhfMacF/LIp/mYWd0JEigT/FgZhW/t4zYU+TPx8
R6KxxYCvfWNXG9GNUV5HY1Ep2VbXSX9237u3s9YS3crepdjzn69YjO3altPb+TOK
XdcH1lcMOiukbXJQDHBkN1XA35ESeYBFN/GXlB0HfGzt29xLaGoGsJWS2SXO+NMj
aokv80hNKCsYk09jvfbSfhIZEb7tu6A8kHKwwFwKVU5xlI4ryMAAYYqhIyQonXrx
Zu3Y0CkVHksP9GRVsRqIFiqTtlC3vbRMTPw0zuQk/an9Mo6BdgKX4LY/b2K2LLxx
GFPOzsTUSH4z+wdZsQTWC0lgKA4GQhvaH+qwQ1GeipT0VowdzIdSTmijnRSP8HWn
xVpl61v5FkIToFhJu80NoIOwg1rZ/mYJAZlJjJ4KRfFXI+BuPJDA3hYjz2/Z+5XD
QwxBCvNr+jhRSDiEcT/Afvnfau5e7o7Ex0+xbR3H+ULzlG6ElRW3QyGmFvOwUJrf
FUh3dkQok0FCgf5LYql6o6G3pzKQthg8Xw4EVoKiskZggkFdiYpOZH3Hs5XSIv1F
wxr2woDwEsP6dONi5ZHDEV/7PqW8oRpnGY15pYqf53CUItBHI2XMJZWdKW7TSQY/
QeHEOIZsA5/nBYOOV/podmrxy9CslrRnOnAJ4bTO9/N2NQttcBcWK/rMDWRgHPuq
/5M+RzWU9lL5QEMcj73myZ8dlFSoKDTngte29+kJnB3lt6fXzqu0o6T7a54FBh4T
OibU8it/MKYLENv3xvNH2keqJdjAtydrXdbI9Cn5x6+N0gl5+DL5cNvXYDlcSdJE
QygDJrQxqx5SZjtfbbPoitLKaj4jZcZYgqMwkm3Gm44ZBocDdBoSBbaqFcBmruxy
osL9usngL2fxOCsywnzfV5hveZnfnY36hHiQZYkKnKUCHMM4DlHlyuIi4JWSiPI0
Y1KdAjKdlrUBM1vIsFU/TlpOGfxkyh/VBOMN3KzZjqQsuH9MzB77t7kZ/q42Jxtw
QtXkOkMTvpr7c8XHzoDZmwvx7SUD5XAs6ccJplkkJdB9VHQiXPTh35YJb+DF8auZ
jmpNt5LLGPjVeJ0NbHC0afXPQgbTru5m+wV5o8K0NMde/O8AjLsoEQ+Dw5/FOA7l
LTP7DIZmfFbrjD+S2YoFakiV+A8wFRiyuLXslzYQiSpvXW7ohcCMwZevdb7LLi10
pIYzIcqkXABxAdaMmFv0NEb03aCNLrxj8AYtZkiKkcthOcMj71m3608okgUPqVoF
/S9ExThUSGxay1P60Q6EaSUnfefMZ8A++rZr62WChqzkAGstLq2khz3MZXxBdEiz
7aIqqWv+zxPvhdyCdFtFI9o53HGPMznBdmbaaFlpyCOsx093+hnrrzsFbkDD6opy
QgQhMNoRHEXoZMkOk9LcbTJYZ4g0LrAYxleiq1+xsVaJzHlhw6AssDQup6Al5KER
lGaJWcm+ViRqpn90vO5JS+t9wuJgRwx5YQvh/wdOMuXHq6vyBMooDMR4arVBh9J4
vvV4bwCV0XX/N8ICSPCYDUFuclUxKWoVAsRWYnY3678lxqxq0R9XWs5xZ2xvJOcx
Ju6672tiU3weH6vXSqW4y/IweLDyjLK7sib+i7hwB9qZLvGsq2XUhBOmYKgh+ELX
5zp2icZNnxnjBVvZXqj+FF7yshG6qoFozY+ukFT5RIkeY20z5hEOLelCsdASSiGE
aa1BgX0tRJcp7UZHSefDZ0cHzk0DzxHOQwOil8dab2p/SFiqYfNVbS+8k70wZynb
QuhiLYStw5rgduDHHm+DIjSx/DkUpZ4+sZcCFJ/d8R1CR2mlpB0b/KQyB2k6mhld
AoiUNmSgdrEkRLOZRbQdir2koUnhs0Lz6qLSZ7S4sMir/gaEzb1d6PTC9LzpAD0P
ElGDWPG16772c1K6TVgBqCBTjXEot9vaFCq1OnMMW9K5i3ZyuMjIMa99BFevwDSp
7SMEJecTz3iXEkE7+ryBDqve8T6s6K0y3x8+7FkfNFwmck4YSl/joVrtazbXZe2q
lhoyWRtx3md66ErLlvU6HfxKxQ21Fs0jziBHRHbkF+Y0/TwvoLnd80rXnUOo4zkv
zSaQr4Ajw2g3/PTFRp5DSq+gJ9sP2+JJRnrGSP3D6i8Eha+1aTJsVJnKUTDEU8mV
Tg28WHwtS5mPWNIic30zh289espLjKS7Rwiu9F+8REq4JTutl7ElIxsCTBlemttD
UnH861D50GpsCTZJ9EMT45c+Uto17B+A5nRT5AVfwvwHFKVqhxtEgb6Yvoabyul0
k4QZrloZsTM6pSFXlMGanriBNddsXJTyOgt1BdUjwBb7jORcdQKXbnWRtdHE1xUB
YcvcV2SDNQxq4ObAMUewP1SXNgEh2lujbrI+AfmbGuo+vVW/hlixL1JnBbR74OFA
dx1K58DPcH84dsxOQ5ATzFFvZU9hoA/1mVQ+2HLnNBOz5kCmve2Z2aeX12KZP76L
ooi6LoUjTj2lQBHph49hFUc+I87ZFQ+osS9hIFIVf4S34cmFWQ7QLqYYb4yJPGXQ
cz1sda6q810ph5LgRugle4o6QkDoJ7Ia5EUkgEFbnk2QFMgsC13ieuWLDu/BnrL+
esodajyuK53EWo/dr331Pw7MvVrAR/Q8n2g+A9Um/VYuYq80KDFmNoIn2Sn49exL
86wOFEpebW+UhPBWEvdKriQjz/vH3lZIU9bno9wDby+Fi8JFncsE6WLfLZDFwCvr
8VJxGtQDXJjyaJ+IjjlSAVOnFOIucEHi17STKwIbrd1c22MP4xxCKotK7Excjqfw
ILhwset+JFZ19jPZp5a2XhzePy1F+ydWr1mkX5mgNsVI5nwUHc/0hHMu1L47xurH
PcXIoh1WVCNC1ZzoSMKrNNbX5m97I5sS8i76tNArcXI+fj5jT7omKNjIDKajC5kF
yV+shrf1ZUPToAUXOf/7nFu+fFArCO7jO6ilaoL095rBgyV54ocFkaA8aZV47ltI
3315mZT0gFxGZ5ESdP6nOpIe7Gfit/mbpdSdHVeoSCMtC2ugsC8OqEayXuTzc8cs
abp5dIPCu3Os6yyRYniFDOCTR97u1fjhl3LuDekfTucENkunBRTZS0hU+Yx1xeze
Xuqep3Xe5p8Ol8tlAvnauSa4AiUtfND+54GCCpWkajlKZRe5BU2GmW4FZUgrpz5N
R5RBEn5XW5zjlYbiT5bKFBxVxaSeQ9w/3Inq3QL2SEYvzoiX8KnY5fIRYt7CDYy+
ytowruABoAtSuBKunaAHUE+WUKRc9niQ5nrbrBd99BiRz8RXZYrx4j1jf15nNpS5
TDwjE8AVq1QmMkOz/GKpDPFjlPxw+UWeuHC0FcQKZKR85OtWPwLUHh4MChBdMjFY
dM7uCn9ePfhbmWnknT3Xm001IwtIsRB9grp6K+Qv2SLhPgeysNJfjCJHh9S0Ro++
n2SrtArB5fCevF73bbqXjswn6FVaNTbcOBd5NkC1FqzsEwj85/8pAWXCeynIpMtj
aoBmO1UMYdiGEQJrQz9XnMavb5wvZHEBo18/BRUxJ+pPVzS7xc/5fN570GIsTiHu
E4kuhFlQ9UvnlS3lvb/kWMWI4hH+LCwAAI8j7rgCp08pvAf/dqi51yHIQDcHECp4
f6IQ6CHFPvbCs0nefDr/HRL2oHstRiZ4JHCikTyZ0JcNwgMqk6efec52dtC3z33j
dADBe7ui4PTXCJ0VEaQWko/ctQEs+HzNdbgruA38zqapnLSQ0criqVs+CCtoSngA
2qPSQGYXSse19cM3AHcnrqTNAbX3Fx7ms5kLWYXxHIaMUCAa/NXJseqFVwTn8TGF
4WrOpd2POEnA8GuuSB2ebf/1Fp+FKuLz6gab3lNlFoUqkGzSEIKRInLvRwo1r757
EQboIdKmterGnvKLu5gGEc8uPyFt/1W11vlussjMAPREXWZTuk8y70xA+/uB5cmX
zFPePcAFVP8+eVxUgYhSqn1872BCvR6aRgS/8B7hydZ6KnbxiopPhC1bJVZJRg8O
7X+pKM0O1hj4UrvxfclxKF8riP9xLbdVOxFQSbbDk9WRGpIrcSbSj44RabvH3ZK7
h8Mzj4zycqgev7u0kLT3xEipjyl5LFLU8HWRWObJKeL0mJi0i5x8syf4ZXr/bWeR
j1E4Zy6Xj/OFHlU00dlD9gc9WRB4HuGhKB6dPUHIOUBfRfZo7xRwZW4W4DmDOxQq
OqsRpyYI3MxpcsZlN0RbULqaSCI/WbuIsCNim/Z1xTiF7cHJ0CnGEOpae6xWWTeU
VFa3GQ7Y4IzjIQ3fI5ZGyoM7EfQ9B6Sq6dYRsB9aI+p21QXYJXI9Ra/V0uGwNWau
bgQnXw3f6M9DXSIecjjzND94CFDV1SPs/6t8ok+Xm6RnFrqH56bFKjBr6Ie+XoSp
dCX+2xA6Tn0g9g7ce9EccWBzVByM/gWM2YO9UywRQZiNZoWiOo3oK6c7YEsw6Sq1
AnHr9amX0RkZ+8IOMqqryCjPtgUM5MNUKT00uPEDEgZXO7Qvz58KRjkneJrs+KJL
G8aDDLaOYwJ9GeLVsK3GOZBUdrpi3IU7XAYSdz7hqPc3Cfc7UPa6aGK0PoSfE4so
/l3jkmtto+7rFGsx3DngvADcro/zt/rzl3gmP2JPm9dH8XY2nPLdDm1e6ArHt+tJ
T+DR2/PIioL0iZVxKhWutdrlDQ4WjsTJunDqpeG6LKY9vOvah47wh+jAx/nM9dv7
DHAlpvWIdFCqwSMqcRAhxovKlzsuthV5vTMT6PpGDRnn/k2KV9PcTxaMPNWwKSgS
fO1zNQI6pntjQCrUUpGfn14rmuixaQRWw34cLg5kp/7lqQ3EkgNyZ18ZtbmD0JY6
0d88ASLNfwo786K5cx94UeJK4Tnfmnm71d+Yx4mtucY16mt3OtRLDpSVSt7LYJXc
N8YMWvT6ug710fC5VviDbVCqOxxvfFuhzvMX5WFm/BBjvFm6Ic3kWumEEIP3s/Af
jI4K2G/T8DYNaxQIDGpX//faBEWECf17BYX3K1ZLWE4Rab3Usx8mRggBMiA5Jh97
2o/iJXSb2p7SBzEw0louAwzfh8ZgSXnbuSQx9G3vgAiN+UYW6VZW9j4mWJ3Ihqr+
eKT3vEt9fF2MKrX87/+0T8FbcRo90wk/vdtNbb738FnAQSfs5gs6/N3T3NEVsn5U
/no3MaJmtFCz47Va506XkUDZ8BD/6hHfvF9i/ilAOnxrGxI8YWCZcpbgeIWUvaVc
SEjcOi1ACL6e6UhwD1MOjkHxFEZUjZ7hRz+u+GCTbVJJge/ZgqdQwqOreQ566ZBp
2LRGAF8xScYpKBcIzMDM/UtBGsKJuEsgm8bt+xA2G89ZlZOSJX8C8B2zbDcbUgwK
S7qw778ggJz2plcxLrWNk6X4RIYXl5FV7/nXjwlILeHqewhBTCZTZnSbTs8XHxTk
baFWOLahb4Dd7NG8CwSrbJ5YSvXg9wksDy6xtN5Qj8t4NqNFL9Ri/EU/GCpfGfpQ
85nkRc77YT5Lx2wVUISk5xnw2BlXNavoTo1KoBPdTVySTzxJF14LdF00Q8+6HhYw
iygNRVrZBSzAG8GcYXOUtffhxbF3S8pTveRuDq+yXh0qS+VaSRCGNhhw6meownKZ
L8tPUdbnzJKWVaNqz2OnXZHj4dlqbakkrdACd5uVmxUdQbl45zNfvsNFV6SuvvBX
pK5WvcT3yJI+XgcGe5e7oypM8jzcU2x21YxNWbTpgucuS8KuzdRG4ph5q6ZeHB33
J1He2c8SjXtUBqhJERhh2AJBisoecRlsA0vsJ8wTy/OiSq+XZerk4IqRI0DlU/Hw
gEXZnYxbJZRCjyxmbtA7Zj7tZH/zqsZLD5vcUl9RHt4BLuajKSw1yZCWKa60gFX5
G/AdiO3P3d32xS/FBHJ6j6emaPkrK+KbchO+2rx3LUNjFIf/H7paXmS8wtGqV7u/
iEJh2pUyBYxHrtOjT8RqK5eeg6SLhqYjeXxkh4SYbnho8MqR9Sb4CWpcCpPzteFh
pR9yAZOErOxkZQKx/cJ6sN3sf/gbVvGxS2A+Jph6k+PLpgbiooH0n7b1e6+2UjBV
qkF918AnhTohr0e4X0zjUfZ8KD6ne/JEZlVSdRt5AA2jca7m5BFylYgrXgoWVPbT
fQ4+gbRxiblw3cNILupnWHneDZntzIIJDqLAmbi0kMVqEz9a2H7AxFWZVDXi9cLR
g3H1liGhl5QHOuScpXgfstWzM6FLAjaQQeN9nsnld/1ssFRzWnhE8MbhRmP5pt68
1A14FSbfUY7p8N/WJvur7kA7vimuQySiErf3on6ktpgI3QLKOMayN6Xy81tUzs6f
ntl9JqueMR9klE1XP12drMkF7GXZqV3InWRFEuWB5uskIKpCqiehewCWLfgTqcER
hNO2YpJG50OR1mV6hoA0GBeo7wXTcAc8BSk0qigpIk+TYbFR8p/LO+h7bYq0w39c
6rqHNhXsLn4SAsHsws64VZrE83abXqCFtBwwrEPq9eedPigIS4WWG9of2gO0tRaA
iEWJzooQ+5Wz7kCOl1rdbral/RaOln/pKDIW5gTsyCXcdXy9Ic+Yv20J+EBzS9vw
KY2vsuYtLHL7+c+65KOevluiX7fQ/Q7Q0n9a1TtaJLq3k9tKprvSGhqd1RlHmxFu
ZqoGcNjeFOETbmbSA0YdheSZeNbHIMhzShhub46JrAWSsJzXCo/SIVmtQT5yNGdZ
n/p8qz8/V4RWNS2Y78EPEiwTUf+sFmva0rjfglgA2FxI9E8S2PwDDxbTdonH+/Im
rRAih5F4XjQqXbUJ2e9l+ofbSaMVDwQx9yYqe/qU5tyvGqaKoquvjFSlJwsKTHnM
tGyn3Yd+rCcif7ScAhdeO4ZblsDEhn2/96Ohyo/SnfEugn0kR5DVtn8LADgXwUXN
iCdFk8UOO/Ku0TWPSMIfR1f5phfLXo1TRc7mJRzbRMhEUKkR3X62B2UzMGPFcOcp
wd/L3UtFe8QDTN8IpKpvGWXJllf4VIY6ADUsKeESDLph4EVJWBkxY+jICDEaaAUn
HUxaaLNk1OKDPMOj7wZLd7AZo38rvP1Pd0oVHTHs26wgEt78LtdIjEKDDFbPzseV
NJRfd6STMwWo/7/UiyI2lIugLq82qek5PGxbluSJAh8mzXcMw6HNpfQPn2PU7j4E
2jYqFRWx63gD12qG0AHQcKnzlQv5bLAScTTQsPSghfK1nHIxrDJFc7zn4pMHkFBT
6RDD/XOZ/D4sZFkfUnxXD8b6uBf6sCjcFcC5t4VtVDbXw6KUtTP7Ujl2NHrmHrrG
AVM2x1e8VvsTxP3qHAAP/PKoYtK0DtZdHzrf7/Z6KWsT/NL4M/Svn/nZjY3YvsGa
dx0itVInL1iPl4VXknHF/PJ+m2KXvl+8ZpfdrY6nAAgrM7BgWnlfhapg8qJHRhWL
Uuz6Y5mfXOcP2pRllyAaVME/Fi1Z1xmgZr9pzepjybyXXusuZ5uKA/raheQ8OGLN
zVHoA1CDgndEqA2yefVFUUcKqwxXY4M6pJqpGxJMVzKQLSzjyPYj+cD+cITAHB2d
yD/p9012GUg2fTZFSxQ8IuubE4GIQhZ9LtQIykSFBcSWADxcbjUC/OBievpjEx8C
w5uBf1/SLesztv1+ETRfnNDOYZ4d+ZiLrdMqSDGp+nkqT8fthIpTJPS+g1TQyj7E
QyDWN/PvZkm6TAWIxiV79Za7ydLDu7hzGPE9+AERRFMCb2Cz7E+Cx7wqAfE5wvEM
8YNxTxMWkVZWYxfCIXHoUcafzv9H+X5YzTFFguUmhbwztEh30eqvd8PcGkwl472f
f8cgnsg/FsGt4WcOoqs/AhGD4Be5sRQPNSrS+VM6be3t2WqRbkZVTaJbqYwVMAxW
aRuBOsebnbP5nI0Vkh8wZL7ztway1ql9IpjNxlooKcDY/Rw60Tdhx2lUNwcJtMQE
DBO4lsNQhIkEyxwc7A5l0WakagITIRb4GP/O8zaTDhdrcGbrIxUhoIITDvgVmLqr
qLWk/N0dMDd3bDPASfk95QJSU56hM34PT9msh/4sb4JHVHGvHECkfDQnnS43l73E
wwQmQ0MMZkY2J8hicA1NctIOr9egIenXdQv+c1sOKyizgRwvcuZgPUk3h0U/ulOc
FXAHy0vo90vr2IZ7zeKgmgQoZy0Zr1iHjqxMss+tSKavw2yzYZjkV4n18hIffYlt
RfVsxuggqndSvNcPbaAHJUJzhHEq3iOBS2uS9oRwHq4TL9Mv5pFy5tqs81rpspgv
4WSXFiOsx3Fk67Gt3C6NDt3XE5i1AZGHyoDlpw3z069sh40jBLKCzTA4x9oC04CO
XGVh9EKX7CTehE2PQ5KjEMB2q55zQeTx/eheQ6zCi7NahhIDAG2VS/Am/vTLl3wa
FgbO8KzLYza4fR6xxsphWBdAbdy1vT+mKmFYlvvpmhJX6SbZ3Ci2JrhrOdcZdUVG
L4ptpGf+bhYAyKr9kDCH+rQmO4YNn7+8rrZ3BbU3cliOYwdxcW5as1PMxJGKMd1i
Np221/cXMbE71J1PbwhviwmFXBS9vTDi3VUEUhO8v0HfOn352KhYoBFmlFZ9k4h8
1Ui4jr6K/KnWoVVdp0oJOgWMM2gLI9hFcu9ZQCv4GjckTBTa89eqmwQxPuL9fdP/
Jn6xGGebc5YaaMZPcozuLcoZ9oJUaGZ+ofAzIGWBw9K8IbBqvIdYWAxv8g3DoDmu
cPFN1xnsRGv3Zb9mMxzIs0OMES3XdGyelVqn+6QzmDoe2RbOjKulgbve5mwfgc+7
PWI+0+oivY2xM71+ZQGSltJ3pMtMwEJwB97Ed66/Di9VNC9L1pId3QAgh7m6IdeL
cqISSWCdyD+Gmi+1pM43y38mZgWw7z/HDRftM3xvHiPDMRwpjisvgG7ampgRURlU
aprNKkwdV0/CzJeW7drDKfIp+cGAgQ/g11kdDCCwWaYc+BE3VmjySQFbA/7WpCOp
Xv4N9mUsTmbL/KKID3adxOEN7ainBLF7C2i0PW6bYB18Yo2Gt849A5JZcWjIjStf
yFnsFzIkOzMXLAmXrcF/jHKcuKVbtOyBSZxwh2ELZ9dkRmTSVRmABYFXyU+JDPfY
QoHEogA7b4gJXjYs+7wICiDqbzpu5u3J1OohMK599yd3SC4iQtrryd4WBYuykNiL
YoshgLWfnvJp8vStT4Pae8EOFAt/uEHz5c3G/RgfOQt5WE8+TYNPjSgvED3tQVFe
9We23AHiG84c7G5N/hQ6C6QyZNtSUMXpiniAwSOyzLXgO2NqPLZD9wV74IC1e3iX
m625BAzDZS/G+74oV7dXLyWnpvmhguvilCsb4iPZjmmcLWpIHMMjWkxuwoDdsliT
V4cqVkA22GMR6TMLFvDETK6P/aaJECBmM+yjQJvh5zWPlvFlq+69K/JQI0qdaUiq
HAH4nxazY2eB0MmhA8edl99Q+Dwt13kbx8PFz51prVBP1uDCJgnf3mROdeUKn3eO
S+PdceKuAcLjcT6nA5v22tiTnUvD0GVWWEZHula+8ZAoOh/GSL8tvSJCUAH6P5zn
gC1JdUAQq2djgc6lfG+K+2quP6ZlpKqOWMe9q/5OvrnVvOVW472eMg9ZKi8MBkWb
Kek0NBw1cU1saWSHO3nX9zypxgxPEIwC65QfVb1wMp5PAyiiNIJSOHdvtsNsndCD
eZWuvH2oM0YUIb2E9OVyFX61uxnTVGW4XV/707rdO/1gLKxTrhIcCbbbZWQuDBhR
DSTZ1I1K3P+/V64Rt+5mWt1uVMgqAndZ97lxHOPHl0RTdCOkX6l31ZDQFi7sOViS
wsIh1kddl/0tw07LRDOIM0cMAiLM6vZiGGAbSplWttS8bg98Q+kQdazYLz5gMRRd
jUW0rSrcc7sta0MBvJGcdfwC09TW1RfYPQxA82oE7Q+2eik1fhhp4q7S20+RPSch
PPtF40nM17/8LnF7Z4Xki40rUSbFoufy/acmOAIhEDV24+6OW+ucZ1ZQxEZzT5Wn
/gMtmYOclWaTg29yUdxhGQvCsbTMg6ZtkS1IDRNL9gNbMW2GPZFeFdew/DnW5r0k
/IX2HdNf5VTeFG6oc5ff4u0SuYDNMl3NsNj/Ezr9EE0nyPHz2MTlw0F1bwWiqWCr
QNcJdtqdX68n2e6lRNdBhKrInYolskL+0PlgjVdRVBBzdytjGu2D9S8PkSeMApic
25JYbamQT7uo1JWZHyI8RQh9pQuitoAtuusJMqjyGjE/1UKwk7t9rTmNu1GV4SB0
q/WXs7+rEkBFGjMqAv3sl6kuMezqbOPDIy1dvzHDAXbrTyPJswDg067w0g3Wiqj1
q28XNu8lxtGRFXqUauMNZ0ZmjF/SLS91e2IxvY74NYlqrzqPSXBOvIQUx5wgHQw8
5u4ZolYxt6jIOkSBvFxQ4dmNwtI2jb7QUdrBEZPIDcjrJsZbfAVP24RIQk+hkmXu
F5roitwNhiX9Tc576aWq/lGwWX1neXV1X6nIUAK2Bv9+WALD21nS7MoGC10yJgdW
HRoeKU3aVflhIJULS+Z6HqJJEhxEisYlvXe4eQlTfw0pkR7++HG/IPravEQpHUtZ
BlfACwji+eSRjbClQEH2U9+yLBfYk0d7j3JAVaDvyA1lFaaOHZKROTQLJvOBHI3r
KZskS76elvOsgj5b6BWLSMdTtdKAQrMfzjvD5WlzAaj3dtdtgXOLnWE8JVjwpNAs
OG0mR/zSdtQgVGmmZCE7gTzj6RryuLCbYKAUygiWir0xb2OMVdUzWZVsHBH9dCcB
mTEB9qVST8a5HwPDCllhsjt778U7QDUvldLZ+Nb9LstukrdJFAuYsphhJLsn4pfk
nUywjUQ8BDCvbxxoxnF4VoDPWof/FdOvtiCYl1LR6Z5zq2e0JDxe80iqQgOwsIqk
30AMtLpR2edINgJb47ez40aU/l+N+aMwfO06U4tfmeBp7iMbaBmivyLyG4S2koAw
Q5fmI6fixJo2HmOzQU64QWsHwF1VLBc8x8WsJHbRB7yr4hQmNYaqVcRVJeOkuSbN
/7uCUnZKa6uq3aqJ1EUGdo+cw7QdpZA8V82gAXJiFVs28F04bErhzYi4RY6XvvNW
Gp8tNT7a1gwso4LdTjiHpwbQlScpXr5VjtSCW90chIF7DNthHKEd+uhN7YueyDrJ
nAE13aEpdzVnubDKI7m/HsdXgNqcELLMugQnEDBpoTeSlyd0GfabLKmSkrr07frO
W3V6CM2aOClEySbVrjUK46zmW2iFHH8nSJ0drGsMGqWioL+pHUg2WPcUjP6vf+oB
A6fmCEsOIcVWhJ4YpOnGx4hocptlTD9NnYcthXVItqk0HMO0q/GLqGwLrrO5+CCq
7p/4tOr7opTUNi4mgM8LsJcXw4E9DIkPc9bxglsZxLrF2o/AYHbU+ec/ebjqMV3R
RRhk1Su4ye0kx7SJuFRN2MprD/Y7ggfAu+yLbDLEp1KMj0EB+pHAnaiT4whRA04F
UAILElSLt0jRwVVx0iCLCESYQkLSDlw+jFwZUzlc1Vt0ergayy7y400X/bX11nxP
nVPEI8gpKbHRN+2cA+Vy0XocuEv82a472B3hlvGBXaBI9/4CDZh3FNV38alKOhyQ
/a8hlYJ7+D99V55mir41Jnxp+KIk4PRObhhxPsTpm/6J/p08sg57iLWkk9eqKI3k
ZsbuA9OWYLSlNpGl8uhBxpeX2Ci6yS87FKgyVHFRxwhfL1EIee+tXH1h96isNRXU
euP+8HEmxXGyHwzDBqDmigO5VlKS+mGJT/aCmoetLzLA0ufPQKrABYkA7hTQ2IcZ
8ZDBGxoeSXJGw7AcH4eqBv+YYb3O4ITz/gwcKWBEs8S2PHOtYeitCY4IKHw8MB8q
5coKCYvHyWyky+Er38ofI7P6WyGtqnfE+lNLGEofQD+U/1nPpWHe23g1PCVXB4S8
WV5kZb3TGr+wmSb+CBreCXvSp2SWhD7hfKIRnADuLF1nn1AijuNlZtOE9H7ZP4Sy
KKKDf4mQVboP752K2avKhOPxvDCCX5KSEyzil/HcMMdFSwBwjVdtzGqj3AJTaui0
lgrWh3hTqAyDROVt1QG6T1ioe7F8Vxjhg8J747Flkc8+/g0DPoa2z79ifF6gJ/Vj
7SQBO2UNpF4ZNZLVOV8onYhot8FqKYA2BtMsJeLGqWranoj0Ceu/1oH7XzUylASL
qP9CBGedO1gmZawlCHPLGjAmr0Z97u0t1aR1G69kjOYAdjJMcYawp0fQcDwF7Rmu
l4glgJpiMiQepiw69qORPOaOXqMNBvr37NDNydUSW2CA/7HVAW/Eu7/jPRuxy3YS
6CHcz7TRVf59WWilg96qjnr9j11XV+drb7yFk7XECie15PNSAo14et6pWWo6ybtC
VIC5J7WpEoqJ69mMW7EVmybJoTiHHk7gxS4UssB6//enKQCj6HTuJt2p75bQP0rO
6Uy08/0S0v39Ag9AR4DrYSbIChfqqUvYHnxqAfkDz3i1+Ft6PAyws73LtIZHP24X
zdurAa6MbpXDPk8KokD3OcVbTDzDAz1VWAQJZclE8nahJdbh6vzz2UGO9KOM2v17
G6GAMZJHvCaRlvX9zb4OXIXhi8TAOMf4ay5ljymQKnAOsKi516tKvLof6GjLqlSr
EGh1I/TzWCBhGmqEilbcouO02Oqf2g9u1DxwY18zfrKw0IqI+GapBMPb4XWnHcsB
ntwkGwwOhaSGe0l+L0nxdbZTyB9QWc4ZJY4a9nXulJb2giUWxSzspDMyh1PBVmzn
x2D6ObtVPjcRq2vHIobgLoRoT9LR354wCBpdQ6ax95BCx7FE3dPI3SoeI9CvYwWM
giTde1DVAKswJhVc+NSUXVhGiLSYFmr6fKGkIhGJd4BigSoZAj0Ykugy3ch3Fw9p
6w3Qs2sr3zC2FxWyngiHpKnd/2w5vWxB0V/AfJ88csnh0g7zVtPZt+iPacYjUyoW
vkl+XBIylqMRfRHk2qP6rsJMM6OftSP8MnjnfDSWXEBLaVagABKdZ04CW2N69ktK
5gNbbbt+2GG2R27Vaf1Ejjdykg3kWDbVhun4ihsAKFvxmtz5E+xEd7r7NUhoixzN
loR0K7ianxbKlM4yFL2jahk028xrAetFS93Z4BUj4Jh2zJjhUFmPHJV6Tu/Eaglu
wpS/n0OXtBv8oiY4Hoz/xU5hp3UqMzQSJomwavb/81lFUWSFqZRQOq+dorWIJWoD
ps8RDQ/EgE6h6W2iAJdV7wZeW4VhbH4zQCQQfZTmYLKGcNoa2TUOj3DNBkZiPHD3
unxbe7MEPm7Fw6ybCvPLIvy25NGkenBvJ9nrDX1rFceQY4bXPpgNVtD5nYEvTmQ1
zOfqGmYwRjgErFMpSBkxJWw4LhpWfwaZYdSO+WxvPSNaoyimVjVrR4h0mWfhCu0m
NU/Su6tgfCpLT03y+1mLBlBDz/n0C4ClnmBXEom/0GLsHZhtlUlCMhUDBn7UuHbB
CPljz0/ToEsMYCsm6DoYNbIJTMJi76XH56ZDZmyh+/cXzMwncHT1O2RXU+RitdVx
MbS9qlDju2lr3vB7KX4idTjf1lS1P2F48EXIG/O4C7myB6Oeeu5pqMylPDAdsg9g
VHm4iVTZyrqTsrMJcm/yR8+ib8+ao/p1/dvC2e2WN2vZsOd+iNFs6R1orbZYw5y9
EE1dgoUXEeIyNFva6r7i7tzikjuVcboLU51cl56nHx+ZZqbkqpogDwT7vWwQPLq+
FLT5xJkmT8f+x/YMabakvqUsVg8plwhy7c0C+THpLp7P6BBogHZ8gh31QryPuOgz
TDEYAa9tYQ2RkxGKeLgBRtaPHIvt9gWnALkf+oV09hm/i72UJHB34BL5fI9lwANL
NMnoImB0i/Xv72mNGXJav4LMt2nAPYzlqJ9he+DMkt0sUlOxHEmfZ8IDx2ubFCDR
6I1fMwGNydSUVjugU3AlwRJj2Uf7CYLvBTAH2JrTbQI8J2o7dvricjXHPpxvqAMQ
Er3en1X51qyqaoBTLCcRVVTmFqk8uzUFaFqrU4/u5FnoG88qdojzxZpaC5BTOgcS
48cBB9mUZyrsvX3Qh2R81lFp8Ltu6XpOMNpbf6+O8F7v8IayQVQ9ZkZ0Q+nkBdK8
ZEhbGpnFvq8ETkhhdatlOXQRe8iGj6XLN1etp6Hr6Pz3xsEsA1Nkklp7cr2efrEI
y/ybqjbGagkjeUn41cm707uCu1Ju3jEQgxqBPa07qwiyJW0lcKBE0c+wW9f5gOVT
X1y5H46Z1XpBJedXns6tx3ZL/5nvaBC+QH/lMYFJhParhKOtXUJMpgxRkmfR4HLG
4YrU/OIFYzbSc/5F9sdwtvtKj2lzz8UNDPVo/gnO6faMJamtEKBEuuNP0sZNKZTU
5bbnTS2LVOahfNGchfPGRCwNjhoFVQtriaV+v7VhVEucKuyPzCrfKHtfxePLrIs9
KLbxdR/QdPnFYyNDd+9aKEKmUGRu6TP2rZ8WhVi5OG9Ly5K6Th3R+IvrXqC9rbHn
66YOXeL/4hHdVrnVvsHvlty5EVdd+tbFTm7et+N2RdQbeCRl3oGgrj4XH6am0xlB
UdMADJwdQRDbgA6uixARDekWNs8w4xPBUQa1TWrCXhjs57HkEWFSPnFJWbAYv3IC
6MFrVEFysOV+v7eZf4wMecaycJFzzEYQbWC8diMscPbpE0fpiBTEvjYvhka3RjeZ
tBvPfUvT+2812e3ltPY/5vXoB7ptXnJObi5ZRclAd2Ni72TB9XaKVOduUVtbyHtY
BZNU2WmwmIlLBQkdGjbDy6ubXBX83PTQh4zV9K6CE/+NNojB79gVJNs495qIlQLi
m/i6NiDBDxXgPdg+QtvjW5Nk4IfX9QxQ9mJjVJ4n6wdNTgjYnibr9vN+UKneBOsh
ZbhYfO2ZFDBaAdmOPmkWqI0wWXla9o3+CGvjXphudnmEbxpoH0L8elbtg48mu9pd
vobCDK5Ji9KLpSvrF7F9NL7TXq6xCHXi9UQVn+reIJRt1+5Ux1bdLHpFMVbWH0J7
SnYVj2nC9Q0Ivu24bIYUJKZ9Ix97NLFlPyqKQXZDVgUvHUrXoci+0Y+6qjsIMDFY
m7xDbdmZ9uf/4AGI9vZZvXzZXwxjzXgv08Cn200Sk7HdjMTNrpka5gcSTXAv57ip
P8E3B2w3kUQIrxbkOWDjP/6pnz66K9QZKM1/9psE5lHWBkSIS3GrQf6fS4XODalq
hrBGVhfI7lo93pDOXPXRB2HLoD+GWxEccDM+ma/vOC7eShLIvL5osEDwDGOJicHy
TzrZmRi5puWkbEgzHoSyZUq6QMHtCcGq3XsUKEbL7kVGDo8af1q0PKov6uXo57ej
uDFEN8Q2dwwrs5C/yjK/ZSunbmJ061yOfV06ow8JzuUJLorN805L6Ckoq/s0nHaB
dQ94Pfuy2NpxhhAKkXPL04+5Ah9dx1lC9OJm/fNLL01E893Z9Ia5ZLEUvMJtrjnm
C96WyP7D6/0IYz5YjXndmofRvgGGGGHIRMYvH6nq7RvmYaIy1a+Bv0+9c2aJP7RI
zY/EV+5MoPD0oEdz4oXPgDhDCZ8knbAXEddTpJYNGkoNbGDZ5SM2+uWszmx9VYBf
0PfMtm5Y3DcLMIo/jLUXs4EJxYule/zpioIxUwNJyTRhIWhip0DkhNEVReQgun3d
stbgEqXgMf+Rc5KubSATHFihKK7pwmRefOxzBPGwHPDzM2VPZ1AJW0KQpTHntVZx
nAyS8N5OhkD9xHI1MbByduzkF1067IDJ+MhzgBEEsq6bLR7NJ9lkCLhFUSSekp4i
OW5B3mdu3BS2jtdTYxcJN519Zc4WHrQK7pgLipKkxJOnUmts1JIQ0VEUNqSjOqCL
1vCjL+IgXrAlYAjKnSW+bLiJMptwcCiPI1LRUQWN2MTQ9JCbWiQwreowmBVpSNhk
W2u8LyTyGd2p2dziPrkA7XagNxJcgt1dwM/6suMJTTSYduUpNPquM9xFqsoPoC0X
hBqpo1DMxgfxWxUlTo99onUF+R53aLhaMY7hlQDfxQhedXAIn0+4Sp7aFhA6dQFy
Pvfbmx+JLxEtjzLOVUS5nWL2VbZrFlKIi9YUTTr3Ql4yZTSlqjkA+B9jVbG+LquP
Gl7G7inx7WaRYkYRa2h/2hU/BwTL91Phz4fO+06uz076kbvGEn2+fXVtkM4jS10p
b5hLSHYboqGWwxtSHG5aki1x02KC3x/qfVMObbZ8x3AIw/Bgna4HiyTFy1IaG543
IjHoi/6oJVoUDJiXosdzJ0hyhyMzeIVPMJKzcyXo1jXOadOVNhEA3jSRaew2jF6q
+x5DGzUMH8KiO2QJvmqMlTVN+EW3eZblVPi+F2wNQ/YwJQ9FpwWN4x1vaNF0uORX
UGa2jXS2uwUB9mazTYlUQExbctEliTyvGF5eYBcSxI1SdDqxcBP49ZcHDpI4+Xzv
kLrQCh/q/EaWOhkY5bQWN9goNUYUKQNszopyzQNN6KAikCsVv6kEPK5D+mcz4ulg
WGSvOtAz5RgfoYgXIGeJeTx/mhehaCOYLkjeE9E2Y911wf4fjob733nswSNsBInu
TqKPCrwzlTr93Pb10bkv0OH9gORmE/G7X5+k+DXVqRRGMbDWB4DoFcVMM3jHFZxN
d2FY/E4XfCa35u+jDN2RG2MpOnfVy/ULvU1TTW/2+9H2rkmrC4y/OyoNFSjK2U+Y
sk3gNLG1VLdJ2XSue0kIKcuHgTYrEJJYStHodXI4BVtqff2falaN2yvZb+1wB4RT
ovy5EWBHefsMI37HLAtYRILrZB3rXnE0qrGHIPgsoE+xYqbFIPVOs/ARmQMP16MM
qgrFzGJWwqBW8GyHd4ayiaCiG7bfsNkuj8nQ/1WwBZEbxTE+YOLCUKwVtAasdtyt
gun+vSZeFZvchs0cZ4Y89aKj2mPxlTxIyIRg3ironBXkm24XH5rjnJ+mmsA5kfBu
1QbQIswVj8CVLsmE47da0DEON69PdPrDWjsOuto9CGDnglpNatFKN7u7SkxMTsb7
hLwSDCEd5hvYMeMFiem4kffgUopEJ0BTpsOONFqbXD+mU1QyrQdGh5BngmXMVlT4
oNLHcKqz7K1LwZ6lfSMAHj26I3RTOHrTmLZZ7BSWisbBiYWLOSiSXk5BR70AOHJu
GrzJ4mxQRvjJnCeaQCuaPP7asQWTjV60CKPCeQBQSZcTTJl8mIK7LKjlxkQF8CkY
CEhzWZdoflYR9nllIIc6ZFNdHK2drIiL8j2tfuvSFQH2CKLkM/lC3bivbVrz+fqu
o3uTKKApNQprHb7U6ZgJqgXWt4+OU90ZmAa0948FeYPDSaeZqCMZKl68ai0cMQq7
ikkB1w2lGhnyzTD9E1IH+WBcpVQrQpNa9+DrB2O7AjgBPpMBfmsuEDASiINch2Qk
mDrIp+vduo8/aDE7++GTnC2lUyf2VhHXP9HK9KAm70owIYZvwh1pbX+6uuciod2q
NZkFiMp5X7zOaxw+ZeeCyTP0Ajy+Yvg6t9wQ62osAN1d+wW5K+abTu48YYh9o35J
tygaMNCdrCoJSScH4nfh0uzLnj7hpCCjYx9KpnXQf562X02Kqdwr6EtjM6fOcudk
NuY6t8y4mk6F0OGlQ8M03GpX+n0Pc0B1zs9zsWg2qp0BAkLNn8lJ4EBKE2LbWmnc
r3j1GSAg5SnNhFiDTDi02vdZWZsf1lAdMYimBF142zg0cWMvM/v+8uxlvXogIHGw
Zykmq6MP4gWvghl8T7O074bOm4GyCuFjNNSM8JaMu7eMuk1NxxSRlCSFxp+QOB2d
yn7z2Er0dmZ5C6XQHDaChth1De2GNetIE/CjstnGy0Khm6fpG5UPblBHuwLbtJuB
KBtLK455DIRiB+niYvr5EPpREioQ1QoIg9LlKxHxfBFaXTehANiYtT2jMUuz3AI6
dTOdW15u9pVRjmn8r7YmgZHuHYlTuW0n8ktCrt/UJjdoFWVgQGgq42KbNhMsHPeY
ei1ldCM5d4ogxAQ2nP2CS8YbaK8FPgUHk3Pi/+7s+AtE88el0Y6K1ZXMXhX3iH5M
ZmdRqNUFr1J10trg6SsDBgABklgIS8ncvzLyG6FY2tyRikImk+fBCEzhA1EOIj0l
CDEO460hMlb5p6856fFsR23XOBlTFLfOAuB5qqXgI6yF/5364EKx81VMAs2M3D/o
QdY1ulX3vUa3u/h/92VtkOndf8sp79IwcIaraONBsZr2b7dlpfQP4NyjR3lqpO9s
NgDC3VZAcNqSaSy+vxTJ9+VVHkZkuTSc4aK5SZTOknFUDdkJttUcH+1qOCv7Ptet
pX6DcJVL9vG45jdSrGf+IZRvhNNSwAmRboSQ9NYkASamkPOavvf0sD78WJ2gx2ID
FkvRNO33WVR0T3g1piR4MpCqZvuYhTIhSIaUB35EjpQjXlooePqJRwge/tRjNbcF
xn/l1+Bj1hDkesQUxqgPv4i5jeR29AGCmkDSnG7MBygfRIuP6lvFNiBL2BfG01Mb
f+vCHBA8Zr6W+JUkjciX/wjS4MSYmWUjMkgwhStw5h3FAtevc7aW5Mj+yIpGjLO7
KACescjz+oEgoXl6cxf1RQGp9fv2gWh+75U5fdlZw+L0XY4VDV85utyowZ0Lm6KX
XpCUVSEVUmk00ejhPuNPDgh4dOA072XeVPIzkFlO+bBmAbwu7LfRvd/V/IHiVlpV
6NYX+g6HPmo5zIP4K0EWeBbmiGRCrsE4yBxRuD0v+nhYx5vwJ/LxGKtFtsQRj9CG
1RFz+GSo0OI2qsmGFnfS+fwQGcSU0z533BsRpPaHGeKBXUbhrbzRxauNyiojRFSP
g3zl15Zk6BC3V6RUC+BRwqBz823Y0Hb6cVt9WPU8zJng3MlVLlSRZg4RwP2h2Ej4
OnokbuFf2AabWeVkV1XC56h2Yt8fPr8MeEiNvvf2Gtth4A3f180IRmyGDYo0dRKB
9nxHeDYzQjue+qAxvKRunj4kmhuIOak63FhkoVM3BTWjjW3S+Db5t/Uvl59c6NqE
QwwucmZW9TukxNEqZQzpZDws+mDCUzbcdlSgRD/BgJ0wT/kfEk89ne204roVZM5e
N7dWD/llCPEJvOpqjQovqnZCSN8Vtatq2H1V/xgzAacOHtO1VI04b+KqWQLDx26+
zxY/Qc+y7meR3VkgUwTfrqqSsMx1Z5wFt9lBrJIX8vRf7ghSi4JzN6pIlExfM7ge
lAjQBwLDwdIJzO81G4Ejth/40J9jBYaJB535cQJ3GGQwMGJwbaPhRSRqG8UCHKin
frWtqSOyWUFQK4JTJ1gEFvXMOFpYkclqTfq3MY0rAjUox7MObdzVNFLzCzfj/eYI
j0SV3kQA+i44nRCgd8J6IirPV6jKUGqh3zlBDAF8nCtyX8s6iDrsQ/ycgU8KgTpY
s8Pdzj4J4KkJ3PK1yTI5LIDPzymU3Pg7vnbaTptEh8WH8hdJcfIQuBdvhb9R1Uu8
mUAKr/RWldaufW9XDpkZwLDmEciMBg5ZZYBP7lxBmr453B/aEiMjRBKxgcy3PcH3
Qjq73m/gAuilKn97vIQllJgLm7hQpkCTtgouWUNnPzX4IEbNzebZyrbiqpsB4HAU
cau/gFyhISwnjz2mtUEyM9T6QXFX+M8jc+shpPeAfQE89lJ6TShqmhW98zuGCw2w
Hg0979q3KmMYDcV+akbfoiX4XbMi1JgVznN8012oc57229REY1izpjdnpxddEd9C
tH7zv2gcjQNEuHfYF0ASRPL7cQujTzEUqsa/1EOkBCtbvXlU/nbZMuOeOw13Nrt2
ZkrVPEQVypwq3sz+F14PEBQgiLXks9uP3+tZ8tT1+ujBR+xhTE4e14zgniNsyysg
fTuqsXWEeME42Petafgos8ISAmzZCthR/Wy+G6JK9Hxk0a2RshFE3HsRZotHUdXt
3xDijPA9sQtWe9FE+qezcZ7nw9Yklf3YJNrM0qhhCr5Lp7q0X8XdZqcoDtWLLq/y
wcGlZ7ENp0N9AX1wO027+/wgvg5PwD+eXudTG5+S0DeZ0Z6uJG4X64JfzqXzOniD
ItP7ymDfn7p3EHrq7hySyK6bpzQWYmmhByilDk0FCcjUrOmfnacQF7LLH3743RDb
F2GAdUkkeSLa2/z4qIAEuWxHu1GkEiDWSND4x8k7+OHErNn8Z2G/j5/aZxpg9iu+
sGFW5Ze3S6J8cHmqyJC32GGqzz3g48fUIFs3cZO1PDMQ+J9rTGq+QUsjebLs0VdS
1GdJIzhX4jCoqUDT5n4jvjPB9hPkNHBqTzQzP66AxJZFTyOshU4B0qELPoYrD8bs
E+VUnsosoVL7R2Jl64dDc/vLFXmSbRWrbKqr4p+lg7Epnapcnv7Dn8jm2P2Yh6hM
dm6Vz3ysPcEiQN8IMa8EAsuxpPiBFLrnIE9ixV8Lq1n2bKO2c97EOEQITsSO5X7b
bYQCspM3c3rhWHrDtWk0gnL2bFaWTWtxxoWenXgh/8IQwPzwqX0n/4lRfMKOa7UN
sAO0C75dJYVhL5/JgyxY628StSS/PG8XNg2L2r8GA2jHNSeNgA6VSV9GyFDsbCfE
ewW8CI+4GUXSjf1jGsGE37KRPKmIGx1GZHMeA0e1/ZaWcJCyymTcLpSWosrvZ1K8
Tkg9SxJgOAjUcIZQAiRYtlwf+P9sH5uArFoGZdHvWfk6JTGoLXgEuK5E0+OukQDd
T377rykbgRPtDked6K95+GRDD2xODBDTctIUx+7s3POgkrCVn4blNa29Kn5DgRvV
o9uA8TDULtl34GcIXXpODJi8CQMwZhKtL6CL7frIee/SfgtHEdkNSu/Fo22XPcHT
YywJUaXZsgWXyYU9ZJzxvw2lY523ah67oKqTnvwPuCZZhgzSP+eQJ+6u3ry7Cee6
WabY3+p8SBC8SrytWM0lOw33b8QfYmbDwePNwBL8rl23CxMll7Y4K8yS/GI3aozK
jcNisYh9SgrX+PoWVXuKPiZRWAEwXQ3J32yU/ApKMShHkX0NwdhIGRrDGMfKyFlH
VRqUzw7khjHo862195/WClYrr/GcIXZ4uyN+LbIvIsI59NxUyzlAzz2mZzPkaKV5
gfuIiVFe64DdBzrkYQ4qcwY6IPkvy9mNSNE23ZB6V+yQ3ABaNQdsGLnyArdMpqKc
Zi53syXnesNtYQL2qz3JEMYabo6SCb41kvYLvXmJrOz4sKVwvf7Z47lEuHE4vTpL
ZjerJ3J20mQSTcmUhv0Hg6Va1IQI7xndi4c8n5tB1Z1hBi/weGwss6SNp9fkXCYy
tImMYFyARjZabloXNi+9lSI1+XP3ObU2nJkzX8goUWWI2cqDTo5rdPuk7KWcB+m8
5jHIjuMMwHBzF0aOJIuKsCwVn4xB/hRJ+8TW74w27G6Rz3gT02WjtN8BDSr4/QoE
znZGv7Y4D9eJnvmxIXW/Dg3aLND9PYcvod+uBZQ3SWO0hTlpr3epRfFvE7nY8XpD
zZ5PoSIqWmDiLH163r13y8hEBT+Nz22r7oxQ3EUu1jLBdSH7anGsEoXJ5r+E+TVZ
D/uKtufg2ByC1IpkjLSNPhzqc0peYZMiZMvwHa7abwOSb2U2IPJk4pN3huAW7wRg
B0Z2iGvKkm4xxsQqMi1tOIeBI/6QNJE7vR2/vWT21NlHplaMkhhFz3yClKl8DXjn
sspsP9oibEIqu6/1h1boFCHon7+HAotB8AyqpIWJCP0iz0RXJ/aRHOtRGEHq0bi3
Pmsii6TiSALCrxKPNUkdAxL5m91K+k26bzD69bfu6/LsKaD4JfVh2b7wuNj8SPYD
RX9LOI08iUCNxIa2QEYmT77tS66aNAxbAjyel6tSujEH5yoHZyQ+5ZkNB20p9WgE
rrygKGMvyavsAfL1HeDfDJ4bSAhLevQJWW2MZiURWNeM6IDTtcrvZDseaX5eNRAw
HfxdlsLuQBRSgW6bUFQHd+3ddpdfNYzZxsR8EhgC80b/xxpKBCW4TI5Wv8x7uqCG
K1A4YHKuLEUn6MJTY+DfFrTuSOox9owIeO9onPkpCQASqsuCYXKHI4QdkofsRvgG
NDrdFl2XIsK6kg/Sn95/IxPRg/m898FzaLqQn3JZ0nB7KZ6xVEnsgtZP7sd8yBrR
qS+VRqPsjjsu+AXwEfez68QfQvwsPPpbisKlSA0PH7waJmohLSxSCikArEwxUIA8
RHLA4TFAXG8vdCXzoTTyTfVxiRqtUaKa9n4YLnJSoAk4V7FgqqVw25nFGhDYXWnq
Adrahsh4OcVxCjUgOUa4EYA0A76M88Ji0bDMPjMA5/muxlnzC3XM06XYXO6c4Va+
SIYWAXCNGjloI/lylRrIiSxa7EmXoYX5VN+ccBYY04IwY6woenHYhmenq7IyAIgs
ECZwwm76dRcZRkjIIRc/KY7+Rqf3dsIYSN8Mk+xpsx+Xaxnl0yEkZFWQSLH0MOBm
oKnRxc+ZKcvooh4dkEuyx1lZDQm3usAHF8N7C/WKfwP1LXDkd4qQLbpRCCleJ3Lz
Rcg2DeR8TiKvBkladhYudwXCGBsu99n8bUWGOPo3Bw5ERVMNDj4I10ADKYbQZWhN
60hey8PjWoMOibMafToMjlRgGXdpcwOD23aWNwmyrZc8iCwGV5CN+73E2tI15NuT
iuVidhlEyBHaqplT/KIvk0jabefn9BkfU5gDZRkNFm3GFqyGTY52ZriZvdCfGFFU
1WgEAta0Vk56v88o2kYuHN+gMp/+W4qJJ3pohWy1pvI0ax9aj9ddOz+fYHSrFYAL
MotJakx6sYr9bK/jLyl++sizMXfha1W3FBbNV+AbsnImFKgTauzX2KUUv/L9l1+B
0BcLLCeKJrSLLd6ZDJbv08zYp+h7tb8kg1AlHpSnFyclGi7XY8OsNxbIquJOywzj
On9geDYSYIi6sPuU7i257FC/Q6u0YzJFZzy91ju0FZ5iJy9HeFMXYfd2i5tsy9GA
hUfX+MKcxDZITszXnPsmiLPDGqrOFzPimusssbxJrejGMHwrXsv9ep9KwEjSJ+vu
JYAJXHe43WyPX901i9vxxPFLZX/wcikT1qDke9ei0SMSBwYzu03YP4WuWGceDK+f
PeL9B7N2/qMyvZesfUTPvR1E+Rlg2SGBqykVBgPtZyQPUZX0K7ml1I4pk0FsQFqY
ZvzD5iNrL/TN4V2gO6gNvIlRRmBn3GB3dtmRkA7ehfkLEx1XGM+SY5LVzfVBU6KL
aib5JTGgDIB18om0+WS5M4pluYv2Yc4aiuRFDUmaPvbRPZ0RjM4J4iFNTtuMtJzE
aHWxVGJRXvXqlJJN3eUbPP7JgfBRRmG6cEx4gOsFnHSo8Xh2R9rfzDbiwMkET4AA
oD1QrHbA/Ta3AF6kdgB91m8yNT+SMYuyBC/puu89tn2WEylw9qeVf0xo6VFL0odH
Nj0mavxHZNQJI+0VGFgG2TJ9asoocLqkjJac0dDUi0yA4rZz3Jgix/djmXo+KyYs
vxjFQzHMqYF9wayuFmc2l7oYzPI6QyjY7iHVX0gUhgk+6M/YbRL8EqL+TADp4l2s
tJrXxSiagS6voMrLPPmVYsZzzayQjKVXE5Medwgn5MB++a4xnBtoUaYRsN+RbW3E
vrE9IAbrg8Jxb2UXmVZQT+yvd+7jTSko2SLy25fM/xKiIKWiSSxRaG7eBUlOt6BZ
GkkvYc9uVP/AhhjEuv5veA5gnCY53b9Cs7R2UA4sf7cN9CeOhiUOSgx/wiM7bXbJ
mRrMWs3tZ4Hb5WrLgxQWzcbidQl0KICiMprBo+dnqoMIojFQwznSJioFePtmVKEF
nOT81NVViRd14S9KX/l3SNl2UwVUhr6cx5wMGCgU+EmSqEEbj4KUSvqlAV3Y6fOj
fIAen/L6TGCSm5WKyxe8LSMkEo4v8qg72ZjY1eusy4lo1MRrqQadu78+AlCS6Gra
dY0akqNdGL43cOy/e8xY+zB1wv2kAKsHL3jd4E7gEYpgE+6WppO2uTdVAbkAsvq7
/NDFYSyiH33tFzebDj5j8o0VuHl5jIc37Px6xSYtSglJ9EW4uvHwJZLgZGFROuMl
KTNRFPRMhqz/v96tJ0JqdOcoTvQi/aE88/SRl/YmkdZNH3kOEH732Igb/KOAkO5T
DfKkmswnatjJNBg9i0RNf1Wy36848DpuffKzoI5qfLtBmtOdPjPObCgzCfRW4tyO
btmMgbFakcOUhBhOmroonNkB7fUyXFpXhVKJzhDMFTyVPMmS9Uz4CHNQ0gKtL8RO
eN/zrD73UN6mcszTcJuihGB62/As4Y6cXVh6fzhmGDH8nosKyUgRjgms4+S8PGlV
B7Ds6NcRLM6NMWKCNE7l5/oWDyU/T88ysKWxm0SUg4JFCxnFrW9oq2GQID1S32Ub
zqNF7Lcx7o3xg6N/MiWZwqLLiW+fN6avaGv7PK/R8pC0naIhPi0Av5xa084WX6RV
766dKliB7WZSM9XTVhCD+ZIQ//C6ZYrMAsHb0SkOfUNuyKpGUxIkEeSK6OJiHOad
Y0ytSc9mlmCYA0CFA9xhNq0uCWBWLS0RDnTMJj1022yqhrRxfCOxdOlaE2Xp0749
2bMcqrUOUX6vZXVkUP2qyEvSZrzinNUGp09Ct84U2+cdy+yHEUlWsqucBAtsyHyC
nsSxAE3RgBWc5Lffpp5upmJCqIHcTjUUWG1S+03piJL4G9crOvGRvBkRL2Qkee1P
cWfVVVKxud26trF3JqS2s1+nqlTlqqRevMD0e+fVjEEsH1lnl0xPUvVWfDQ7RrKo
ZZhBGQNCtD9pjdK5QER4nB3l41XBZCYv0h+OFRUMSf1ph340WLqeJIZTu+H1ty+d
iuagYQcXqhgsdzPTy2Nlgj4+GM5/gLsSsYoDZC5oYhMbon2xk84Lk16WMIsA+wbq
WjLxWBre/DuNU0/F3ZVyOQ3cS/PyW93UDmjAFq6+rcgen1+rDiHpnmm+JH4aBjn4
5gxt9THfSKQT5zy9BFUglOcDWDFNvBSsbgIhcnutGUlyYXp1vMBzqqVQrUQ4qKox
hNVLGbfeyKfOzxkwskHE/+ViSzgW72p3TWFZ7XEoB868NgQQRxwOKymjJrzFdqLx
VgxQhWAv9gmgu6yxMZ59Lc+HPXIjzYDT7rOcIuM5s5U82B3E3DtyS0PKIDrlGQNk
sSJwixdkz5H6sc1VH6Atxjc1xii3IAHExBnrHVvEJIJI6ABW/sIANwWeMtrBqIHF
maK6qDe7NDUzSKJXQo4VvN/iEWPVre0dUqpIE4TZnGHg97NdanouQ9HlST4p7sI1
z6Orx3rlLee42K1wOFR8P2EICmg6Bb8YpFbig36RqqAYAR81B6BnvN2Lt+2QuVvy
Nc+2L17Rb15b64567xAGzr8DK8X8anAuYPXv1Y4M98b77DEkp8wdaEVRZ2GVk+6c
j4XEROGCwTfw87o0NP+jdNM42DyuNpWqhmpkDweXKNvnfBLtd8SRuDUQ2rIWrWMn
YQaRabmnptBtXdFe6JVqUtbpWFFGj7Snl3/XKv9uzVwgWFzuupjpTAecnMC10cn3
TrAeufuhWEu+FuOAwxJsoP3DMG6wd6OCLt5n1RgyphT/vM8NhpB0AL3oPhjYDUy4
POESVTbD9aAI9pEWUpn7fDdQmijmK/Sfe5Eo+KQ6ood3mJOkBYeD7jfq1ffBrgCu
Z5lu0ENBmcS+3hU1FrIGCVWL0V45gbwqhck1tVFd3KZO6wopXe3wu5gfnVS9SV6K
3f+XD3wfItM1AUmSobJ4X/8hmtY5/vwYV7NB7ZXfNYZI6KCeAgW8pFjq35sL385S
AZ+7ootUmOOSjOh9mdinrPuaXpnh0zjkcrcVLmHHJ8ZGc5yrqOaU0YA7SKVQu3vO
QhyExWah5rFbIG22A6/G4W0ovepdRDfGYuBFUarU++NH0KEWi7j8BCoHtGsH7G2S
5kutU+eBDaKc8LBNYX3uMKksa6S57CkZ44jRMD00TcIjs+fNjSCASkGtVmFDr1i/
grMg+IT4Rh3Pli9ZPfUL0U9w0QdMQJ9fZ47Jp6WbgnblyUMWIIjQytwDd/zwoukv
2xv8GH+gcaQl+PwPDKbANxwos1e9/93NQxwUuJP01rvc0TQZHnJm6g11j+ISMUb5
pGNgWYKRUS5jn8IRQm0oOKB0/XngSM1oXWhtAi9GcQh6z5SI8rGd3DKWTWy+GB2g
Zq5cq03FVYQKYUFvbPcs41dzMnAwsrqcvqFuiAkZdhAwezMC088OoHYpsKdZgT6E
238rDE9T22+bWd6DYSZ0hDNLewFXY2lSd+Te7mhcWST8YPItlAOlvfqtj+ovXQiK
LvvTCdDPoz4uPcT48zqjkuB033WeFNi+9wktn0oskxMP5f+Bnguaz+M1Dk5j1cb/
lFBXUAR6Kmy2s2lsZebIdB5dM7ps+SxkpR4C20lr+/C79AQJEpw1K43XoZUpg7e2
mVjvXiydY2G3gzbAq5ie9rAI/F0ejtfZhpdVgsxIb7yR5kHtqaoJ2vfGvL2933Ys
T76vvliIADn/sKG+LTPpX3So68q+mMSMNL9S4RN/LNr6sJeGVqEjsGo49UoyC8YZ
qWZiQgn8Rz9vFtbpmKkcjrl1cKUiLeO6qDzfF8+5b+MARfPh2mui0ilQRB+uUd9G
YT/EBuQ/4pNJTS1Dj95HG0UqC01RlqvlZAT5rfKQZA6XEN4qYyonCKRb5DEq39E1
uWk46kqNqOmU0EED3GHvcahqLrzYN096MhKvxFFC/kpgZPWQlxMxmFaUuxKJf0Ub
91zO29jNww2EoiZu6lY9/vpj33v49U2QVr7xhrU9dT6lblgbt5Kocu3NksUJMotE
Zg40Y0vvl1kmt2cKRZxphhsR7mVlzJkeTVW0TaQCmuSjQPZgKlF4I1J8TzqA7EnI
IuwujZLozswBiZdDB77x54qXiTuB7mitM+QYE4VCnCoy7oVNzhkviWi6EXkOq3Oc
+fNJOITuNvNHEHZNpIqR9ZEzrxYEKK8k7SqiTLqzBVho20X5b+w+jJLyYVnjnf3R
hP/2fKFnCjQzpQwqmRYfyuixm6R6GMRLVE7mZw+zTM7SC4HthNs27uGqx+5HKWPk
JaHxMJJ4FiZuRFb7ZtP50HCwt1hIUBdnJkDPEKLkovsGOaRwMBM5Eka5CGTjvHLP
vtptZmesyY10McYyrbzk7Rv8QKdMkIZZQS528ApIx8ia8b7kZQwPfh9+M67Txdjj
BBbc7pxZHjM7TjqK9/hiCBvnr5OJ8bdpJIn+M+2204E36U5X7sMnHvF+IhveW1Mz
MkA8fms6Gk/XWLxKoTtEfjKrlghH+GtTr/jqDK8PQTeONSVnGHdcD2jQQQzPh4pA
c6KEKNiThngZDFJ6rrG/sS7N0+Nl4INTyjKaxH4T4vWvSIcGPgYZZ1ouGbGHoiH9
Wsc+7+pLVVlv7cuIhYrpB43NXoTsGYaXa+fs2MgmDis/g5fmbY+enQcuAt8eA7UO
rKbZmxshkJwmcYOJrFokoznFWnHuBmNN0jaqxbydrq9jCOlXA0FtGoIyMz6EJD8U
qtBbTAq3zZng7pnF+0mXnTtnuwDqL2wx/ehsyCO7MpduVL0SCdrWzNdsd5/Z+Dy9
u9iaLpQmow6/m0K5XEYBxDpFteiov6EXDXQbQotRZj9gH/hnHv57WwnVVw/JXm+v
ZiC3SjOfZ1flPXmKStLgIQvhB5ESGZkCj6xObkKd5YplrhaT1pu1OYJyGydNZWaC
S0NlceZpaZgVenfa1nCWktgD22VuRguGTmhdMhXU5NoT7yNBpBLAa5v620OlGOEg
4YEKAwALZcFA3h5WwaKHUryHSXALZinj2OxF4Au9kg/y8E5LnyE8YLCXiqcSJcS8
VbXD5/DppRKZSE3k7SFYHXNw7kY8o8B69KC50Q4gShiZm02lVbqQ7SBUOX71LAgt
+cr8jC4bszMRLoHQ1asY4IvpBrTyz0jXTiNzuNBVJpgi29Ld1ghLQy+GMCeh7o+G
peoLMG4GELr4xDzSeB7s3C6P1DjUEhj/7lBuN3bu/cf9UkCJkM1Ets75bB1cthuo
ggg4AjRUda/tzAcDXH9QNFbFqYZUjjTavh6yIOZhep9kuVyHMAOT5F28a4zXs61g
ylpeq3awxS+QXUgSxsdqhEOmdjW0odI5HnQ/42GPc7yaHJSZWCwVeJ/XPNfJXbaE
uW8/ZF6Ee9PjDjky9O6hAHen7WWUaYQLm0gMJyJx4Siuau5fVCcAhzGedCu0E3T+
XvJ5sb/OqLLsUhWvP/7Q005xFeox9Ii8hDSWnwFxzQDUK6NNgiKvotGyuseuJgTz
h95Q/LJGBSegflMI8Bz1awnFPdCephMGEEOfVtJFghgXMzMzff4B5PNbn9SPQv7B
46IKXtaKfh8R70rPZTarIpEwHLr8VeLSRTcvshVzZsakO4bDXniKOVvsql3AumeJ
XnhxFYH9RxM6v0o3gNP5DkaNYJ0fJ30V+RAJoeviPt0F1ckUR9343F+dyRnmc5ni
WSzkdK3J78TgokqXmagp6H4frN4lyj4O7yJtvHG0BIBBDc+ai/R5bGSQbGTZeS+z
SJhYJ7FS0H7ceL/X0uRkBbxbWRpiAkgk7qjSbO8Z4G9OWznRRCeZQQ4dmYJnGh2M
wGDgr35jDpRVxfYl1/OPxuyaMKo6DgYYcitmkFHmYYgltSsQIe51U78eSjT3EGe6
kENrJfxA8kYpgrVhooOjCteemJgUXr1jenf3GZ3UG3ahHpKc/dyISNZ+KxnN+X+1
yyH0LAqgILvxu8fcpqSoEVsilsgtgLqBF0nEF14t47DkPZV6gU8f/XuqnzzV4K4v
+fdj18kQXebj4/S+ivJg7A93S1KDGgmGau0fk5xE8epLdDdx/yjtN02rCxGT2AQc
/qdAk2AzdljWYhhlUxXqLtsaL5+iXfkbRLI7vb8RLNGSZYQvf9AIkTVDTLeVWFvV
lYSUILRNJyj/QAC1H6sFkvwNJqI7rDlumMf3/QXYvn8F8/Xx1cL6J+7/ox06b0cI
/yGL3+8rKYUhOmHo3f+YkLD4Qcq8LVmOQnp6EEBYv7ZtO7dSH5alZJkyip5OicLz
ocVP8r4XiCBqsvGMlESs9/IMHOTW/srXnpwCvuKKGpMbLLW0/5EAofoigvHnetHu
nz8Dn366QNpgivJV/2irKZ8UGx5ujHVhOygoubX4kY8r9onIsQTRCA0IBkXSFuXz
Id8opTjT6H78gJoYsF5DGwHHtqFiv19VrvGScpqZ0Qn+2HJvqJ+Lmym1ZZ9ud2B5
3qV4uM3rjqCEJcIbIQI6OJRwQJTDuY9bsuFWIBT2AxJMYUX8EgHmLpu4xXrj9gxL
pCPbcZEh85BLKoD9/qbhUna3QNP/+wHBzbQtcHfLvFN7RJbzgTOJeMLPSb0/NVXr
WY5GYafAWoWaPN8+F4zUGTz3CknviHfwmhgW8IRuWNbnm+vVn8RFqsu+Z7NR50Po
r/Uivg0y8To7oQADASJx5O/BPIUYixQSWDe+AQD5yR0dVivkpl712u0C//KHtOBr
8O/+TYcP6XVPt7CylFNcdxdFZYMgoopqN0TkCeUsrsloGPTCJ1QF0hDVDjqWsn5N
mxoP8TYjCrOF5OlI72hUWL+4psLrqSpxrPMU/VLV/MJlKtvDYy9ZxUkrFTpsCb6g
qAfgryW2kWkhZH4cgiKaif6DL/Ewq3pR0T7yU8T16aM3LjTGC59c9RBH85Vp5ToG
7QphePWXZG+O4FSMlmlsc55imk/7UaPp7D0JEf8tyo/ciyLei9Pd28JuthxTVApN
jbaSEM49lgQDFeYtWI//QNV64Zsz08R1BpbXx8rzCLkMVBf9snQpv3ETVzp4o7A5
4mt0SplVr3EHi2sDr+QDaVr7OtntCNmHDBBQhuzqWFs/1nR3q47BRotrQ1py0lN6
gCC1PUDUbpGaLl5fbTO0OqhaL3m4siB91zXxg4OYV9Y3euooThDn012lXFFipSXz
fo956YHkegfuUKhtrV/38wdsSK9apfeS0iJ3M32dQDs1UxduLicCGD6it64Hsgv3
wz4SCi0ir5e6p+Mi0UjAzcZPFxiyukoV66M3QXd3CUZriEZE7nqUelfss9de3L97
kFcqor3JsucuVZ1WV4njmSoLw5gUTMI94vmxcd+WrVGt6BeWuXeYwKjI5TnmN8iB
Udn2R9VpFXOl07tACJbSJtacfY/ldgMfxknLcZ9ElzerknL9lWSWJiz81WqIXeMm
yeXA4B6EMBaxBN8ue3qZJb7+KFJ2wlrqgRMn64zvFHckvHzm045Gptmy0QHVGpWX
oWqf/6swvsldsBBH2ELG+CutOJHctQdU9mp9Hl4UpfI5mP75yF6pMwtqHe/AiAwF
wbWHWpJVPFv/a7pEBl98G4Qy1C2mpVJHg208CFbcbnGUc0Cd8PYMqXmSyl8tP/fZ
uC9Ixv8r2grE+Nb/2VqXBjkVuPOxbrIRsWdtBrRSsDy39Hy13nGGGWnhbHchZmPH
7uMnOaYhFunKFJjR+1KRXCEeeeSFleThT2/ZhdbSxln1NOufCwoSCYsXiquL/F1R
mw5qlSujmXaZJ3JFgF4xGc47PZiHPx7HxzJUH2fX57Jc0fD6rSZ9TgF0ysonhRIA
Cxz+ToNV3NL8wDdaOhvkUvUaiUqD8LylTBG7Yxm/Lae8SXMg6vcWsWrb3X62Q8f9
81bD8MzSdWYlQdgEhD0dTKhc58CnvyKcshO17PgTiOsfFOJ+yYPJlFKkPm94K4DP
BK4CVV5JGOt6Jk1DNKOrL1I0X4qo8IDr2gs1lnMvYbEpIokq6jHBv1Rl3Xm/gtDJ
0McEDspW9PE336l2ocUITSrha0X22QETOq14ikHMv0stqPkvUsP+DDLTSwHF63Ve
+LtVbnawGQ2i6MxdMUznSDy4iYUfKi6RqBb1lA1370Bm0PKxTV1CwnZles0FpXOl
Uo+s2zi+nX35N8rfmPC8dbJ5Qq45EvwT2fK93RKybvZsdPeLlr0HTmNB/OqsCXI8
0bUJF787siHHqXGJ6Bf/EZuzinOd+nbbZXjX3F/lqzer3Df7Mzo5fDvIAHf675kf
xVidkcnZyZQ96VnP+PDA8FO4Tb50/mjF1M/KeJ375iimQCUiwTv9NsHQOj5Ej0YM
c9CI+XXfOge1JmnG46lvYgDs/ajKIweGal0Mikhfdw//o6IuJdrTL7pcwsfZoYFC
YPJMNs5BzqNoox2k3SYUK2zD8y0s1KhQkl1YYuPv1KcxFvWi6Cg95Tz9RHOUgkRB
8fftbmZJyWkl423zoa9PDXvAZ/cwi7lQxuzzIFCXkWAegEyHvZcK20hmZWfyz0RM
S0ySVKVZofCiH0qijlt7Fx6e2sl2PMo2oRlgmbcHtXgwR8asCaLcK3vtc0li65x0
5+19W7/Y6lf8LA1SxSK69TU9+HqrB84XOJ9zywtU1h+6aQ1y4Nku9NuCCzNt6V18
hKmQ7mf+8sBlm5ql5m0A5R9O4g7PPJkSFI/qVff06bIeALdvm60YC23pFQNkEBMq
ET5HqTDHKh8GiXuPmq/PGPq/GwUb+dzv5gnwZA7upR80wwdQ+asil7QKikvjj+gR
VTbrjsWGHk8ItEnaMt2lmcUb7usjLrUgtWzdOR1znnDABCq7Aw66rPD9gjtjiLY+
huK6ftoB1Vw0E7eqgBxDlpEyHZ3tZSeqPvW4WOtaNdG/dPqKVsanXYN+XwbxGtMb
n/ME1lrH47HwByJ3pkstmIMsPMb+VkbWa2wwbZ/QkNfj4MnX7w1onlcmJ6x7cIO1
jMFeslgBNAWXwcH+mEVoDVSeSphfgYUKp/Pi17JIRvcFVkdu3scoA3HW3SfXTwR6
exAvyS3sLYv5SZjFzPCiRXcKA1MeyxxZAFVCdeJJd6pBD8lcaFSXoIr8HNbktCsm
jO4k6SsG/oU+BGCWu7e8rMMVHTDEGEF92qdXlSI+/jsU73vZ2gyX2NBuo8pjQWcO
+72dZCgNf6Edsm39jK4ieifl70ZJEaVSS1to8TRsLgBIXjcCisiiymwKto7UC96v
UWDKThUf05UTFvxBYCsVK3wwjB75z38oeoHzAB6mW05b+G/gkIQHrhpLXP/91rcV
+WXzElFYjI1WXWx64d+VaFxlmG84YrbW4g/nO9UbmK8msrbSCZi89vDyAf6aJAFY
lLcj/do3OI9AMxvyatE5K/JWQrJdUBm1K5t6jHBH5weLByLoVoPDMFs/N3QzQsC3
2JvSNJVStixkCxoXQWPq/HN1RbyHKMCM7Xyj5mbh/TiCiIsK30PZQQCvMLB6f2D2
4Jn+rcOVNjQRfDw8REYYY79Kqa6oQ+hXF7QjzQKSsyHe2bPQ9P4Ek69qYhUynT6A
ST03LsRMNFHYHhfUP7aP2tKKLXeoombYaaG3lZQ/W3fmphNh+25fjmajiJNrwFxo
EC69By++i3Gjz3jFU4QqHCAYxfgARQKZvz+2wRgv6//KrWi6CEPZTjykrRQjzDKz
tXNMQYvOTFsQ5Khvrr4aRY7bgcHO4oMNvmXh5EbxJYJ+rzeN/LdoZbd0MvYZUs3L
YIqH5OSH3A24LV+GbDabpcde8z8D48k+kmCQF38tJFTxeakBTeKWaltXuYpkd1tJ
A5KZ4xxKASFWenJIfEWKAW/7pMG1HEParzRq2TTebsmh/kMK9ybQ8wrWMALi2gfW
RaSQlHbtu2TK+egxEVGdg/E9u5Hdx6Y2NinPNe0lKNaTGlJ1Izqnd/4qrYx6GpN4
i2MGO5cp90uW5Bz9RW20pffmF+8Cx1Y55p5QfS+QvzYvvFb+vn/w001gvdXQDxLa
N7myqxm6xeuEewbn645PZH7SKZa4K+w9c/BAwpPjcF5mz/kwHzNCof9+gq2qJsz8
EX7nAX3lIxQH2H/FWgvYvb2VUB5uiWf8yKWBo9DvR5d0Lix2BI7uMlVcvQF3U7++
95xUx+AbFHxXtjDAlWuOw4Oz4LeuR70+orasPMAWnzAPiROPQhfV/Jahu74KiBoQ
Ao/Iv6xmwgUMpbY9OVGeQNmXggqKjZb2Gn0i10KlFb8C3f7UlpiZ2MqO4cS9tEQ6
u41N62MhD6uiSBdqfEO8HW8Lfr/afoAZeyjpfgu7HrO8tFTw+gjV/bKHa1cbLVB5
/jFLTWkwCdKhzYA5jgyVXYXIK1dPw8tJduH/kBZ8tT7BMZt8wfB67W895oQ+H/3U
hNfF56A52m4v6DEsTxEtbcyc5XK6ZUnYG7MG0dh0M//xlJ1szOV06LpoWlYpxVMt
qItXEc0NM5Q6LmygV5VrZ/sfv5jdCB0r6anG6+6l8NQKsbk+6lmQayWUR21wJeBt
B2UwtIAl1FsFNSWUqvSgBfTt4Ab4fO+h+OZXSJcw5f0gSFs3V98hzRFR76EOUtGq
36fisa9hUXnI1eWYB2Se0cV51uupuVjA8iVesOGtv4fs/uMP1GLv5Hi61LgF6LDP
VpHLr+f9tQ4McEDaJKedN6+E98Tb0FEPrIdK8AZqWEn6pQsfOid1VJMmR70JRaka
bn1un2I6ujXWmGxp1sul/nh8St7Y0oV++EIXmNs+9f5TYf38vvXfcj0oT2Fh0XW7
Z8fZJuosJLfd7s8jyJiinHxTqRvjjWC2/Eabf8KnbFmhkSS6wK7VCnX0/d2ixFyb
G7DVK/tKib5XIiRo//vpKOJSS2sekokTvynmr7Q3fwvRjcscQ1fXVKoLN1Ty37PA
p8rDm6X6HBVS0gTLllqK7WgRQMZyjhw/K71usPYZIoTQXsaP2SPphMUKc2TJ+zIV
ow8fDEt7RkXEYLaVBz1sxvIBzEUAaE1l5vqfO7FCwdefv2eJQviSk3ZY9zi8jjNI
2dzXoNckexwwsiryLxUHq4UWK6F9loNr+sFb/m96j0M/38mHTllAk51gXps5CP29
K+eEFlfZtnhiTtFynBIRIp6COg61EndkOz008p0y0mrTB/MsUsCV94wxSoXPWnKd
r9csnRPNbj09PqOb6VTgStgzLUNWE3ujJtMdlEndhZk5KALC/N6KiXDbaHzQcN8b
vN/UoTXNxQ9QI9tMClmWiBJfCIR7I1Z29PRNjRa3/nszUiQbk4095FRCiYjJdjvN
hu2gCcg992eU3iF1T2PWMl4wb19Opaa9KDu7I9HEvWm07ieRKvPcSjJ0X9A7zLHw
rktFomkRmclZoGU8HnEWzcwebwph3dLeLhtZBENTZEcWD3/njYPqmof++gXABFw4
9rHniKCaC287wtbnf4z1QyE/ue3OfwNG6VLvrtaSXdYNX4zDKusAmHIsaTfsf6uH
m7G/ycxMrYOnBsziEPJAX/NrZabT09kret6FGawl+NLieCmviAQVOJmqZrsiZruA
hBj6vMay2vYJPOWpt9Ko5CobDGDtA0aWJcwfe/iFOcJBnNsrIHlUbA3ahLlzqIel
FEgUbTW0KqM4qOnN4gCfjSnRGhleIWSDa46gMptW7UvNrYUdmuNQ89bF5Lbg8MdO
FhF02zJOj2xsS+4lWcO3rSct15sXB3MSdZjYvtKEweXYmz+uxnmpAEl2v8FBbF2y
AKN4rmM7tl/1WCU4AmAiYvDYc48hcXKgN1GednLMc09JW+xWLDekmdCo70HDy1Xi
hwC/ChR8QwaUE9Ba8fboGv8MOHgls2ANk4vDsTXhhjits3b6+CgDxJOhfTeBSiHC
r1bndOR4ZoZ/JYrQNGNXZupNpbK4SLtplk5LtkMb2z1UQluFWYy5xDRte8Gu1jqd
P+/xW376rnpnvdVFtyKgU3k/CHStSSASY2E2m9/6J90vzQdaXCQpYgrgA4LwULsq
ULqMVXptJNgQ/SbiQhBbXj6iyoHBxljVnhcQUsxw8apCSA6elWQFfaAMlhze24eO
bjPFFl+oCIittoFNTsj/rIeVt6g1Q52CaR0qEfYkKAcXHkztVYQAH/4ZOpzxNwEZ
EIsQdzaJR/IsNDpS/P42mL3x+6AQe0wW7HS1AM1OmEncORS8UOnF05IV2KxpBqvI
uJzgx+9AQhlB4F2q7HpK9Ww301EgYh4T2u/PtXr4uKu5siWeP0laWxbwTHyfOI81
QB6AsNkE8Y2N4/ye1f/TxhYhiIxN6nAKTkZwgVpQO8JqL7SnazjUFd27ZU03Otgv
SGSkMwYdcYAo06NootvpOoB9udSE7FBaB/CzYPhKNm9p6VSHoNJLLxyC5+tnvp3C
2OCxUkyjVLKEmHVi8Wy8rwNJ7F3Xea9wSRrvYsZqVL2OrZRvRFRvzYnQDRHtG4uA
U3Xd3Ime4ECLUoFgZpHljvqn7hIsojsdpWsFxNspobOFdCJ8iBNUniVygz0nKD4C
nnBjJUMRArj/WZ7SSMlIOXGEvLvUh15K2Sjqhhw1uI1mgg4GNmojPzqjJhzsY5I2
wsgySqPy1bqPT+aEWyBZQdzFKHSrvN82iqC5IqQSZeuejGvNDk2NI0kP9LQZasDK
/vqRT2Mjpf/Q2PhHpsOFU/GEqBkKRdjAH7yyyZCiQeKMsDLDejzjlPmr+pVN3NiG
mIYYRWfeMCbNam9FW0cZB30cE3jzQepYVCORMTGQNZFBVJt7SBR3Yw+CKsZ415ir
CqKDc+KlTJd29Ea6OmwmkL12HBcFi3NgGH6M4MDdYs4k910EzwXTg1+VQMZqsKm5
z8fD/DpdEOmzSHYWFg1uoYyLvQNkc81O1fzlnACVrMhg9RrKmSt7X5oDLA85Q+N5
DTjuN56Bhd7U97JUhfeMywUZif9myXx4MrxG3s6ionUwgUe5YWgOgqXUguXL1VP9
i2Y9ICHLePwEBRA/rieaFZ6eO2JqGAEARTuJI0TzbE8byquheOyTbyCbslOT9Fe/
3VKk+lyTf50TY+Yf1EW7FDhUPQCoj0zHe3hGyyKJ+vChJXvWVR0Sa9rlvzkrfvUc
rVAY9M7c4nLj5//1N6NOFCqZPfIlek8JYqJpSWx77hb7ieYnWClpmOuNbaAw+EQZ
MmhVDMZ8Shn1jMJo1nJZ6Hqnlwz2tkPt8zo5igJGxE1xTTDL8p8J2l6u+wFzh29I
dTge9aK+xzcIQoq6o5KuG7sew0dkDdALRjswWXxvSMbPycEOQkw+FWdUG1GPN103
eLYO4K0xCk05JHfgwldgPHodd3/ovMIkep3ZcaXWM1NGbbk1ehP24h8gvq25BBqv
/m09HxsQcmatzHMF+yF+CO/jQYuSfx+Hx79XlDEJPHoN5Qky/zQXAWcrn/Nc2cED
fiMgUDDdkFAXhsrN2VBbfvi4XYaVcRTddqDW4y1s+x0MHwOb4quv5Xb7dulWEeYn
xdq++B75mZ1xCrav7vPVVL/tRLEySoi0zJ7T1ME85gDMMvMVQYwa8MM0L12nUejV
6NfY1iW4vDu3CKAG3Iodm6Q6vxsBqVBRop4CLNkrwQlL8QNlN8HNfwBl8p1TlBA/
NcIa+R4QcZYKu2lkOisdOWOxcGL+YPkjiTMJvT49GmgTL6mBKDbMDz1dWnOZQI5B
EXtXlgG8W/pWm6IFMi+82JTadNS5+4v/wlDYd/3S6w7Ik60/sHYNQDJxms6fSQav
W4ZYK8VoPsy71UDA8HaIOHYMyNMLLVepz1hNhJqV7tvpVLgZGrgLBaS1iVg1AO8e
YQLur32Aa6ScD41QcM8/AvJv/wC0xcPT7SjL0iqdCdMtD51XdTiqNmW6Q6j+BSQo
BfH9QhyYYIEeiCd59HmQDARseQe97YABVV2/mH9unZ3kmFp8CgJZQFrXP4uz/bjk
0DfWO0aG2nn92pQ2lSkRZ2aYZIE7+deLVa/B/czsVNdBYmfTi4zNCfZlzS8DMfJl
B7WLXRHie6dfh9K7rA6dKp6xhEsSIXIoZjK61XIPEIYBQzGyqjDa5i+D5POzqze0
l39e1qrWBFDQyrIVolVcpMSflnSuVROLa8IS6LAfFEYt5kMjaGp3WsIFl/3c0yCJ
q49YxtFFB4Uco9zYX7YuEfyFKbSoeIo6zG5umXZ3EAKofX24jsVpCEA/Y+FlWj3u
Y7gvXdE3lSuI1TtYhaktdKU8sVM/jHW7zk7r9GzknrTYdA+Q0B7YI4VMPoZdtBlh
HiKgmMUoEBinqKkl5P0Q1THONFR+/5kKh66rbBbjWLkJkWLhScNBbbyT1MES7phS
Eld7Y9nrZfoKKknQ8qMnKZQBFKHqybxIUWGcpR/3mWQmcdLIzwfBVyp6USUZxzyR
gh4pfbTZ5PHfzX33DIQZFdUQD/atHd6XO999Gyo6xuZPOjGd68y0u6hcsa1fPwWT
Qpaexedzed2tJbst9DjfE524AOMxftCdL27qu/4zF/8PPm/iSGvwBFQ/zWioGXto
5JVJ3zUql2ckYusmOUyMj1WjYBWevhQdygw3bM8j3cBkLGlmx/NveMKORbP8Mj72
Kf1roIW/tMlBsgJuduKx+VeysUzyeuBF9V6KsI65gTWsbUX2fiJH30DOcW4Ehnnw
yMHMzcqQqzNBct9dL0iEStYtTAS2Yve+0l1fKn75mEJxjnqBYfB922+hVXh3wuJl
FQl1sKYLJsFDAE3sLGs1A0tvp6wJUNM3Qk1N+O4sw8ygghpyBZWYs4WiaRLzir+X
X26lcKreZ93lgKCNLcrKBIs0hQzja2D5RD1AwPr+tGXC5+QT2boAswE3nLV8IN9K
3WzJY21xgaGlIewCUQQcFmy9OYfWVuipmoGZZq6yqlA9reEobxJ2XcFicHi0KwMj
ZoM9Xs5LDkgg6TFFyImusfjnyqtaVfyJzo+nhPK05qEL5CJmwbl+QcZtv89N+6DK
VncACaJsMGlZN9BlNwRUW9hqEMgPDavC26XUn/7mYT9VVI3Jf9p1VY6rC+dUFBuh
cDT+f5/8lhUS1+/K8oeo61zcEnmEeSgG0srMo2VKZkf0B0okT3Rdkoh0FZ4VdTqF
DLvX7RHelC2UPyLGOnGftPnIBaGEQyRBeJl7m799UKH9h8naLptmw6ie1cPR1xiN
TSwkHycjaDjZNltMsit42tX8ZlegolHunMlfI4KE9RUJkVZRz2NOnNm+NvRbamaW
0LeicmoJlSTKX3Me+RN0/AiTKBd7YZaP+5wApUMNprUk4mQhRcVI7xYLN7b+rHYG
8+cXxYZSJDzx26+tfVA4F+JefQ5+r+YeYJQv8Gstr7N7t93S3zgzsZsYDHLtlZ7L
HfyP6nWPHWTsJMmkuUHANhYbscJxEkC0hzbyz14Qw9claxS/OZ4ObcQqgMzZvfJ+
s0P2ROuQS58F48BCvT2DH+9fAfCd4leAgm3r/prnc8DTPmjMitn+1oPugbaKziF3
X3gX3JbZW4saaPXMG757RrTTdTk4a2+t5nRaOV8vi0qR4TfL0Yln3L/uXxmPndNf
RmqULUPVk5LNI8WBw1m5lhgdZD3s7m+D59ef6z8PBVy+lSGelt+pTpySkRR6Z7QD
dL7qOC2AhpNQ+TWZXoxT3c9RV5UwQWdVxDZvXfGvRAVevf1JKcEoYazX1hp1UlUx
NPL8cimK3XlVVRwUmOBf2DETuurjTtQ19YhJ6xUBbM/3J00XXfipn8MrNNC/573U
+XeSjBU1xTX4/t5OU0uV4mdMeOExqLswBhosQiJNviN7JVXfBZfBoRw+CSu8Ptyx
SQsQTLt5l/h5JbtRxnLzVOAuzU3O+18S0QwEFbys5N9sX4wqzD+vgX+SeEPBCvFK
sCGoMf5O4xmfyRYMop4vPlKochJIjXYPodic8R2lJtl3MRXIHDd62EdiYKEx5Ck8
Z/m65E2wpVsAKoyKWTSUWuzJM82B0O2mlitC1MSz7uBA+J+c01Y07LJC0f3vqN8b
3SHJZfkj7ydTMFVtRLYbCBGK+3QZ+uGlB0AA1P7ihfdaN+NcUnCADp/h0kwzHOnC
uIl+exxttiQHiPDXIOtcgOnicVGbXI55M+hNhKIdiWpkVZtA5FXhm46lg21VL52d
kuWK9D+SohghqYhSN5hD6VwYg3WMOYzmbpr2hJfNVrJRkhJithw8rkhHqOosaxf/
XvrjWAsaOVUFNxUn3aR0DgVmgMNi66f2LtGLIJt5BaGarivyljFcec4BayZJ6C99
y2QX3vklasY0x00qr6ncmDTD/+aJ1yZcIgLvGxHYujImQ7ULmq+M9jshhGFNMx8E
Qq11ccZhogyu7eWkFjyCD99kJoCnCZ4hiQvHCB91oY+dY/S2fJ4z2yjjff/sbwEg
G9aKTAaXIBeijqWZ5TED7BRPaRvLS+GDgSMikH7aosyU48kAaRhuqGYLdZS/q2aN
K/UilGqVRiVB4SNY+5ROLgU+4iTEide41nb2/coQTV/TVKDGYa3SJMLgVab0V4ST
2J3sTsWq3ySRLg070KX0QUnrecc7CNzWpQJV7qBG4tFyNF0XLYvNshYUa0QlLvaT
RIwwfu/s886mZohtTbJtc3VkicNmoyHEWx5TTN4A+lNlGLnmST7y7CVyPyfO2AyB
oiSPOlm2YYzeKJr6c2lMZYCLKJMN5XJGif1Sf/PxfD0ziT6UDjpnAZfUqQZav7S/
j9RAFD8T7Wa2ZUQcAbxjDPxXEBK93KrUP+zgvKs6J5KMN8xs7ed92bXtxDa5JnSh
CHkHVqWO4GNHq/hEOTn6WXusmsAWQPIP9xskyW5Yvs1cJc/FZeVZPZQtXpoeoufC
u/NwHSDdIEAUM4DU91SUU5uFuWLM34xZWAa9/XxIPoYtsSMWTwgjat5+tZ2YcImc
cUwzR3p0Ea/1xc21wT3bGFP2dqzb3PYUVmumVmxX/EW865Nz0SnG3tfMy4xRufT0
mVmNtWPS7BzkBWBmbNLIsmQxmyny2PSc1nGHnTy9vZL7fdjCsX8PN3NfTVzS/zDg
zhEMHbM9O+sbfllOaFdbGBdowrMXO0WyhES90ce5U//V2lQ30mnbgkz1ukPHeR6r
srF+m844De1+KPzt6e+mpWNsNbMsmjmP2NxCzpf6nuwnb4a5c5pBd5pVp43l00mT
1yNFYQU5+6zH25G7f6GgskzgWJrRzjDbJl0Wd1uE+GQlz5BJzevaugR807tnLq24
c/ncZyFGBkEWGkB5S7ktjQ5n/yGaAYGYBHFTK2ZzuU2Mfg6rNEPorEiJNUWnJm1p
l9Hsf/oxIdsflSFqUkgp5mEQcyyfRHmBARQYD0o4NyMlRLJsvHy254MFn1xmgBUz
Z3jEUZ0AO2kF0EU5jnG6XOSX4zzYt3RD4VLhEeoV3pJJAXolMeC7pYZ5w7PIziB4
mO2fZwM7r3aA+VNPhZeQW2vTAw7EosiUFNpmPMGP2vfDjG7dZAXI8wynBJmfXNdh
NFciV7PKcdlIujk2fByRbPHUhM2oaBlbBopkD0TPgXcWN78s0V0M8AZ1wMjhsP9k
xuUsTkafrXn43OHJ9PQzCA55faicbl1LLWKJLhnIlUFQPQLwJHuccJNyzSW58xop
sKn6U+Nknz+L2frnuxkMzVzndo42VALfcPe4lVjKb+0UwTOAbay+ITfaVYPGYytA
S3ik1I6efuMGu6/zAGSIeO6hroUxh9ZToqFxs+6GFbKuewQox+pv6pIjZMtiMEdK
8MCAas17cyBsc0MvC6DFwcXqqkocc34/FBIt2oZxAV04v5NgOzmeDMifLGDQ0Lnb
ywX1LOO2suMx4YCbnHndTm3r6NR2cIK3oawptqzclrbJXaI16CzycZubZ6ubIZdk
vsMOlMIUu2Zpp1v47hSceRjR70WGtoPoVtIkX+gNK1qD+zytglWtljkWqiMUfzVF
YN3fsy6ccrBbeE4kK8nR9fBR43SI3Fv0JVd8dYfleqkmERrsOlYsHDW8SAVVjaki
rGn+636M6mO97ztmYB96q7fupVF6gdCjoX613WqhdnfKV07LRnhULCVhTTRXubz4
IWKtrgSGURDcJ9/YNNShYs4ofkZQXTSxP8E1dCvwkT1ZKTNhYl6ODGXMlUGoLWBS
k+yFwB+NtKWCDgFKAlIcMRyQet+IYamzeYtbVQGGNU0Z8AVCZgYvmfJKa5IQvKEX
L26mvH5ejqGxKYByBQVyAiSEKNev3VTuIAKyQGsNlmzwGuuc7tExQu8K/a522nZl
wnycoXgWmsh4/TnNCaicUmQ7PVKoNrnODlvtcTaTEun/+OtP6Rha+ssmUOIuFTR6
oymPc5Yw8hRpdSQZQWWyPozVuKujWhL58PhJGvq3N3EfXY6d6N+My/4Equ3JNjHB
CPzLIa0HZez8b9ZepxUH4IxrhDDdWBrUlBNT3vp5o/LMh3nx6tl80JZBZEmyjjEe
gn4aSwVylWUzS3T8VrclHYTiM2q+PvFaH+/MwYI8Te1tIqN/jXDQURKpJiobq9Ah
xXYDicuopK7w/INQObjhd5VAIzfF6maTecm2rCKJQ34YB8IVo1CzdHPFBORW0tUX
4v5uUDU1nY7ZnCdM0sDbIxsuQ8Tu4poq0RrepL4ykGJPKka7ySJ/5kjenVm+if8P
7884Mig39jJVXNUJE/Fh710flu35nS0ywza8CBnjbw9mHlL+jBDsdcy0LdtzyO6r
MGUsK5P4hty5HmfHuagnpTXkFC7Y131OGX4NyiXysL6qTP06PI0+zaTbJH759vhN
G2hiqj0bywj848zBGmWcOtfZgxN4x7Hz0mfEzDIklwRDcXRpRNxsc+GdqEsOQ4NU
U2wTjbKZVEjGiTYL5zqAdYu3vMG/ja+Dow3FQkLKMA1c7lMQooCVxgb4kBrwy202
dbDMImuygmVi9eOFd4BOtha31XcJPmhASka3DTxL49v7Kb4QXpMuUUXZBWH4Oqta
CdcO57uMS/MHGoREoyFb/79MwHl7vKB45Shav/fdu4KERN6fYXkwmylefBbbPPTW
Sg4gbTOx6IMlnA60AURTtVoqXnicz0NieDm73M9V/dtx3ZeSa9oQxeLI1BLhDHuJ
jOOpbQ2ZnohlOuCTDfVVh60ZM9NyAr2FFB2Up1iePFP/sOXzrDMLmTZ2ftii8UeH
RvVYpXUBicmOGnM2Ny/4G+awDaJ+O881SuUonAOeQTJEKPAv/EJftGDvYJeL1Ab3
jzmzvcVgB7HbxCyawQi+hDFCeIKsjNztTYInznIi2sPsPRGnRkvQKbpjCvrGeQiI
8WvbfzXWmldfUFWzwPW1c+eNleVrFci7rTmaPziCTxxeDiv9XhYmkZPXN+lK+fXi
MMW+GP99418smvcs3VS93HG5I7eX+yWTohrqHZqJKCQZrZT8XjRx+IAtIOQmeEia
oSV6ZcVr881xduy4ZkxSkPKRz1OXoSFcxSLkJCyQq/k5SFuDfUxJVduA5Z3suXa9
WZngZK8WrCyiX9lre6vNNZepqUWM5MAvMtAZm1RuWtCmMiqH/XvLUJbMv+gYN4bI
00P40B8oT21hvGkRWcdhEJo+xbbbCyU5WimRNGtP4iu8e+6ju1gQOwXmRepDZgdZ
TmopE882C2sNaCbpWa7QF2Ho5iUoGwoPTYpSYYowT3XkhT9Hxkw/SSZr/Pqw+W4y
KxyPOMQ+oewSYVybSof7FAVSAhMyGq+e16uZR9biA34GQmdUCrVJTmy4lBX/HAbG
l5rLmILNe/4Lj1rkDx086i9/h7zvYp9avNfWxaxKcX9F23OXRTgnsvYJtLLjO8ke
OnTyJLH5jlDofXufc1SE/wbTho8sPwEC6+US/7IOrkdxnJhVjYFf77FO4FFb1hgT
FnSuGlN8ojmdDETkWWdkfIbV127nIjdvoTru/o/ThiL9ReHmhkGn1/dLmmchxTAV
oNTtWfpGXR2SSQ1O7UMHlT6Ng2Jtc+vvHakXYxeEZMnLeTmkE06KvBYg4HVkK0Ey
Ag+Jd/ujUo0j0sW63ntVj8pvxEQQcLYhl3iYfwJZWWf+KL8NGRmrY+ohbGLF7Jgv
U6CZETuuW0Op3HfWL54Ckr4fC2vT6PALNO/BmXRar6PxsoICN9+1XKaLqrvlB5Cu
hb2pfUlmdxRUVAyJJX3hD9YgXu70s38mH3eQsWwXoMKjdNgqnMlah7wxzyD+x/LT
vaYws0srIU3tVQut0VtUI138TnBywaLi509QI3gfch3B1W+fGSC5hoaMvF1p1bu0
pDFbiWbdDsxAw7JcyB5TV9sYlqRPSJjCSHRAjnx8rWAuHBpN0AFYVeHYHvzCG6nt
uf3nNWI/P/TNgpsimhUDTCBahZiA5ROd+G75fATfB1ZDS9mCmJQreqlLJBFa+GqZ
CA9FfZXkSeSPu7yCuYbmM7Rqfc3KT4f25z6F8Fo5gyGA57DLL4BjRZ+l5A26YUeZ
ko6025srVoYvobVO8j4vBQH2WjgbK0mNjVlWhW+gamHgjSw5Dbu2qrxmgMjQysk+
6O/x5685hE4A9RrclLKGjYToJcmW5Fo7cX4WQJ/lJmwyWmv8PjFCwEcIdYDe5vzo
PmVFWVwi1WuR+/fzhUk06B7k36Ds062Y0+7YUyRo3NpmAqzgMxbOQUxl8UZViPxw
1lpRpzdXyImM9kFOFAhiXPEECRTuKDstV6+fAtzvwPguWfPe4NNyyHr238Xt/UZJ
8dzPLVzu9ZyCRUNrYnCKTvu0jYvf8gEW2bCGKMEprpwiiyNcLGmw4qOErmQNSiqu
D3mMa4g4lkQayNtmV9cWSpkq6Hd2O5N6zmcajD/heeXoIVHcmiXmPBzvkRH4AoKb
+cAHmgYjzG/QBphi6Br5PGOcXL3md0uDO1Cl6Lhp/W96KpsLKF+eCcwcsRotALCP
HOEWJpFazpl2+y5y2stK1mud6eYteKD0TY2RJT6QZCv38mONSOMbVRNM1xFumUDO
4lY2dPn3QJVpeijXhC9oTpSeythsRrMST0FplaA4UOWQ1Dpi3ztq9YrWbLmsHp7B
SJDONhPDTqw1ddtaPl7jn20wAyiyz2iJlbuHY7vT9rnZVsxeZ/QgVdgz98yAPN93
ZEB7wzXzxRYPjBLUAGGc46FVzZF9yDKn7tigM/oTO7KEX33xowhswUuzxkxJALsW
UHJfeFlDZGwRX8BnhIdMuDl38M3vsKdC1cr3cKgQzptlcSwFMPv0xi6nZDUVE1Un
2MbX352as+uj5D4UAOMbTXl/WedGMyegOXLrJacIWqRLtp0GnIWGdxE9Z2z1zrCL
eWIhy/uV4I4Bn4eTE5Kwb7cBZ+XjRwLnavgEQAOR9RbW1zg8t4c0HVhmSKCWof7E
p0UvQ7gycIWVLe8oq6mt7InTg2VjJxGBlXVCQ8db/S1B8oPxVsDpLVbhwA0UHDhw
uiSGTKh4dsjVRhR4qBTsOCrbF2/PWuRJKxCGDefK8IgmegtCxS3Mr46K80WI9c5w
HQB2LIwrouRrAdSNlWQDMHXFH5s8DCQ6EnR2ju/WP+ZyB0pAjKP//6JbAkIzWykj
CyBqzcbuqIBxRoWgmgVF4sHgvRQQNIas0pb6xmBwXA3VJlD/VpHzxV32IemWjZUk
m/fNQnSIj/ypz66QG74jPESaUlci0k7LN06AOYlxK0YfiQwM9/tOhxHTyrqE5Hq8
1OVtwaH+eN5PRn/ON2BjMi4y3HaTtIainZDLM+pWc5MRlUS1SRz0omZ7VixTNHrA
x/lELu0UUygRRNAXjOqibNQtsnaRK9lQlhgX+nNTa7liIc8CvPl7+3rmFwFqf72W
wP5JrMlK3/JYqKvhU5kjUuQC9dqkxaWAYe/KylH1Syjaq86IX3ELkrf+x8Ff6wkd
+HMJg0RP6XfbyqIYqOfvEcaIejLCagw3BkqgcJVctktVFUqM45VCp+fUb6vi7INJ
CTSS+hW0eryK6e6O2b9ZqtueKFqQNKTcV4a/9Fa2NfM=
`protect END_PROTECTED
