`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bTtpVKOCPcLL8Plf1aBy0ZdBcj9XKFRHINCS34l/ZQ2n69gygSziRIYZOSPXCpCj
HLBQuy/MrUM+vmd1cWowq82WlCNzSxZE3Sgnhob8BC8AJ97PDtBzPcQW7NztlyG2
M4cvfnNL5SUejlbi48E5r4fy8C707ziQzUjkwkzo8TdAsNX4mI2FxmOiNpDvVlvY
IpLx1y2e2mT8+gFZO/wepxsWWQ33Hk4daIFjCpQC0Gdu0vNxLNeolmQjC3mKgF/M
bsFLiDqUBwhb0xBPpvzqYGFnR4ssViO8+o+hEBGh83E1jd/E+uDmTKByTDXct3JZ
W3NfrodgSyr3893aH4KYYYWr/7ucq7IXhZK0gU1IMvBVwaHBDDRORQad5HpkraEz
l/JjcxdTwh19SivNZs316+7LEQf8gnqPHbAGK9TvT5EOWOSnP+a+3H/g48AAeiVU
B3oy09t/xzWQjer7blQJzLW/DEiu+crSldGDl9PF+boca/kPZ+M5PBKknO1Qx+nj
`protect END_PROTECTED
