`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wO7tMNfKN7NcM76dkEizlLWFueQR2T5xtbHS2baKWPKR4YrWI6+CFVJb21LfuWSV
Nq4M8UWYLypsvg6qSd+hzuW9DWzv7rBqOZMvrnvZ0y58Xj9VEM/1bQuxRXmw+sLb
uFf3se2xCqk3tC2LJLhO2exrczcGERbsDQvU0PnNog4PZnuzieeapWGPZkMUQ3wx
bkfW9SlLtlZV3z2PPbaLWFM9/TUh61WNoV+K1vE9TKRugDq6k3e5IP2fDaChQPif
JVjQGXaZsawpTDee6PouUfalAV7SSBefwnJSXmPafx294+f6fvurV97+aoR/NH5+
DAldYXOkP53mcO+aF4fHQaOmitzmC6SxVVCQwcAxLTbz17lTSGG5PrEzIT4l2BBR
Ne8iE2FGAlb2iBsEupbhzN6omMdpLLgrymGtKkocTxmH5mJT3WPzHw1EybgGm/N2
XN3BuPuX7K8hOPQ0gY1dMaQ+CkrPkythBrdngvUKUmv2T6dS/KjrxFhud62fxrJp
wpcRRk7QZJHOmDn73h+OuNr4UAuieM9n0cxDr/SHLPwAfrcPh4yIPPlgmbHkxpFT
tEEc4IAXmDpZdfYJkCArag==
`protect END_PROTECTED
