`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KzQZ/mJw25rNoEJcgLhbACW1/8G93sdCFdJXOO0muXhNfkfADWOo1Qxui8E4RKnd
1UR8cct11nGZ9V12YozNF87eBvUBAw3LNARbsM1JYRBJn57Xe11fHHZ7qgD85SCK
Zg4nV7SG+WgnfeO+sY0uKUEC9oNLuyOsw62XVwBbT5+tlF0XeCuyfUOrKo6OlT7u
ZiSZnJ45XoTgPNnymq5v/Jwa00GRz7/FiaVFDhwmJbOFuleIUA5RjZ55dYOajGM7
NXWrIajT2KytAfeydtr5WTrb4IdUEEb5wQywoCJG3PDXjNuNpUEx8UukhsnnRhJp
krP5aZUF6E6VhmFfbvoD8AET9lefkMp8m4jrwwsX+vw3G+KLkp05E/evRs9KF6/B
tpGdSfxIMfcbJVQdmup8Yt6Z3kWwXxribBNZDfU5xPbW45eXGpp9VFDDqxAFOsbc
v1Vq+Y6YCNqrbCIlyG1eLtzRi8uf176+p1gP1SMn0pYAhLjMbyLTcG6HlxhqQ4LJ
4h/HLyozSGJ2Et8e0YtgzVQVHJjQCx//MfjIzc2ICsLU5/CaKfZfUhlfT9XbgZr/
2wjMB8ugwZDDcSrNO8F+4zohev4pcgjPt0y1JEwfxyKj+TdpDZIsM9aG4WQjINjm
C9zOLzMPGufyoIzJ640H2LsAIsaXyRyZSJFnZiK/4CTZMG/sNrES3iwcOa05KgkV
COTsMf6AZWoTgO2Y5PDz90YqYxsO6zxGRf9O9JO8bxn/+fyMgKTvsxDnN5LR3+40
bXNnXhRFgKMj/Rg2jkd6i9ykqfFcIEBcbM1ymcpFeL2Ym0FEYp8HD6unSdPuHKsd
GN7ygxja93DvmdgKtArQBFodHBzc2hRNjKmE7Ak/RKZE+LCiZwJsdgSfzVJr09cs
+AiK173Jh2UiYYoa8uUZfHbzP0xTvY/WLfmNhdPaEj5X9wlhE1nd39PI3Ibgv4Sw
igalA7zq2WO00VSomxPmFEJ9E544LJ2+hOrFyllD6VXSy4MTpZrr8sFkHARWrDfQ
bqpxr2TVK3CsA/qsAX40XoENrSYuADF8mev2ecJ3STKOphq84NEQVLln6ZRc2osW
xsy9qN3A5JNJT3I1ICw+v9yJPQzL5m0nQqxkNqj9gpMc2cCaukVbvFPfkIplyKex
oLMcU+RekRx6TVyCdGdbjO00GSM2+i2cPSVLQo/C9jSDY6bthYqItXsVAeODpfN+
VxSxnALdVkUHb8OPCLZ1k0y2d5sHRHmIq84JAmLPkhAyUVe8qg0+gwKSq5BvjpE3
8wtXtSTePwjzrunb+TmvsmxayTIL+o6QHtR7El2MZEnM8uown1KfN5x810qdyeJU
ZKylZiwy1dofpLbjHBoUCbKjf8NRmpvdpbjMcinnFpqUpSxm9L+f2D13DZzeAE2P
dN/lGdLh2lUloYdwyns9uR1LhaPYKfQyJM/DXmUVnJSel32KY1m+OPDSe3N+zTpa
ZG5j5ba+1cRLkf1MdlAAKNE+Dizp2l+ANEyFZee+YIxZp6b4HduvlW9y9Xig9Zur
NS25PoKTg/vIvdexFl8yeeqWnQLTvpNtNosXrMbDu5ZnrmdbrD9ymcK0QmIsFR3S
YBNey3wQerVDw+aW0T7e195dLTAgpmEH0qvYC85GZKHlgQ0kAh4FBSiyuzHihA+G
EFL30RCUx9uoDYFxjITUNBebw6l03cRrj3/4fmQbGOMiSOUHMNQDcYf/lnBly98C
P1Es4IKlcDold2qBMdUZ/qRBDf6JC0txeKCGTo45wn2qDlqATa1ujL2lEvL745FX
BifkwtOsXSQXCcPgSGIrFtzs7aJw5xPkEtmMpWQUxIYax1ThKrRJjZyivccdUEMf
7HhSDmHcFisU+qmNuAV6V3ts54Sg3KFFS+0RQ+FqnTBrnzYHihF1BXtWvvhBwKFA
B76fMc1rFAIOoNDkVFF1sWNhUtS/Pra4XPzS/CR9mkk0dHKp3Nr4PRBtepTLzndX
HBV+xjvEVmES59J6/0Lb10gMeRcOu/rP04IT+Z07iZJPGacdreb/8uDyyJ4UpvC6
Qk7PYjN4ZTCxmkUljdpyyU2cEDA84PChgOSHC25MIhyyXWSFZda4mJfJHVvr4Wfc
+9TyVtQfX/BaWdkD1EIPMi5iJrfinXbmkaB3PWA0L+18QopGY4a88yHoQmWdnnb2
W9/CMOIK8oeIJJ45K+nVGn0VFMc86ofRWi2KEMoQ6TibOt1c9/N70mPDw7Ll5rNf
QKVc9PG3Lu2ZyPsUzcrXHbWsC3/+UlVeTxwnJG4UfDaUREGauGOU3djmYEGhv0L6
KXKlNi9i7FxxtaEwUZUjuDCpFefekkUj5QuZhOyBoldhnvulHCdYC2rT1HWwb8KO
TG9ej0slD5njH/BNevg4yLRFBS/PAhXy1yOcnHLgv8J3DLvkz+GxghFZbofDt4Ic
/rekV51OMGSKJjftEcgk9V4wEEXYOCZx3FmD4lI6IIkzIJfTRwqr4fzTcJMsq4VB
srkR/vrJ80kDnM/Ws3yqQsYfoAcvb0PV0LhFvoY9IXTwsZnj0WC95K+EPw4ClkL2
S/o7tonyuMpUuACCDtDOdG6VHLC0Q1jHrT1k53TC8crefyNGd6e1JdU/Xc6GM4Mr
mXDbbuU90EejOaDOnM9YBUpoW+I3/lOWrVOxTKLmSog0U3hLF7XGQ4uNkQvgvmeT
kYaLm3W//9eAz+l7kuZaGz+cVYEnwT29OhaD+VEHqdquypS70fjXs1P4x9Q8oFRb
v2MJUdyjfZ+wSqSb4VXtymIeO8Hvym58GBFdPRmS4i+oeMRWcsxoJZRAHUmlEmGq
pXUi4YZjWTpqX7z4Ku7XC0KcJyFZIFLfItkpH0gsIvOxrS9o1siJ53M5hlG2vZm1
Fihzj8UvUUIn2eAaov5O0fbqrCtFzQF5gdNWG5sDP+jmQcON1eZcbFjXWfprR1L+
LeAR+0xiypxXLYEQjhtvrcy0wpAiyJhSt8feynU9mJFr8I980HAVuQLvos01uGP8
Gb7hETBpgLmbe7AknCf/WsT1ae0w0gjiye2l5UFkYzP8O2dnGJFYlCXNO1OeQL86
ilj9m1rTycVk9/1Lf+HvYIykkSd7ztP6YB8KOgRGOiAgBeVuHSoLrFL6DoT8NQ/Y
iVrKN1KlFpgwKYa5+AK8oyw3ZZ9DF01CSbBk8gFbUo+pdTwCfpw3MqCRe3Gikm8E
2rbwA310ZzE6dYOWrOUS5xoIXr4o0dlKC7rwr6RmHGKcPKcptHU1U2U9xHId2g+B
Bq/zgn76eZ8mxW0TTYywfIPmpVTopoMpu4mL+7FrqfH0fkxla8O5spPI11Mcanre
ZSlJi9GAYYDebp7h5osvw5oObsYMsooTpYx8PfOSBW//JnvwG0bsyWshhKgnXaLx
soPPy3erl/xepUOHQ8dagNJM0pIKcSZSllYhzzjmCp1CS/mYr/A894MCVGiXljIq
5oOj4lvrJBi8VjWkZe2VaLMkkfrIQm12vnQ/2aO0BijnZ8eWACr4hGNimAWprx/d
teQKPdg53hQCJSflduPXcuyKiz/bcKuepHzhpx7Tr9eWF9PUqiMjq1Qh5ufTs/BZ
KNFVD+rMh8ohrdGpRYo5AWxlZjFOqA2mkC6U5v3HI38D6hsxKMwBAr1AOhf6+XsY
++x3rvm6oTQ71WVNPmCjOwYnAZFkrAnImd3YvbhqUXoJbT4AQg8G6MKR++3iXxJH
xA7u3OVGRZpQitHkJ1nOzQskzvzwC08KER2PIJ7ej/S60pKZaOvwwdLuVNUdC58M
Vxw75amGKck9cv/fJ2XZs47NcxMK9mcm225zrEUWvvgQXjpzlD1gWhqENOR/Lz3h
1iV/6VN/eEXLqGXXThtSYXv6S5JYpyDXDi4PlAUl5ADOImRx7+IjJTWRnbZNaiHW
wspJd+e83KsWQ8HeXT+KrlbG1lQ35485/PNmp/gLOULP0QI0YRlDec3xr6xrwnBZ
2tsK6rOuNrIvkl4mzx+rEcOlcQGBhjeP6UNDPUS9Igr21MwiKxjUz37LC86E1hkd
MxsaviNeJSSsDbqHjFfsA52jXLT2VVfVnB+wbevAH3nZHADDWnPNTgoZUz1jBU2r
r9g2kg4c66f3mc5eTfiANZecbaD4LbNM3k3c/jYrO3p6tws6X/Ky5yRKryGttEAs
Apnv+n9cCi3xpTdpUO6Pu9UmMbzLecrxIsOteZ7tH2lTbvjXWg/kEsgLYdag0ial
PMCOXgs74toL9Nq74BhNkkBGH833zAE6HaEAZlLrwmZ5GXysfTv+Hm/SQSfBl8/C
qs4H9MTxP2s6NzXjDIUTMzCCZwWxElCENqN/ExLHkCyKieeL9tIOwa9uUhKDoyJn
0NDygbZm56kl605MlfN/nks1Mjqy/wurDIYtfLNGVxIeLr7rzdjZ/Tdm0tMALmkk
XpE/jcTUhQCAs+/XR74/lwCtOqsBcLomaNSy09GcuMEnZnnwasSNwdbrMqCapd8L
7H+57Boy+nFsFCVZcKkhIiB2KCGL32Ne0/pG7m/fTkWD/QBHZ6c0aqlQTdj4x/jJ
bf6e3wmdEeuuKRGdkG1lSNrWFQcwCfkUZl2E7iwOqldfoWienSPvFMoh/bNF+KxL
TfZmldoWdirZmTEHJWJB5PpMmJIGRBdd4SIANDJmaL5WW2VEr3jYWOyKzvP5+QCH
2ri6nk5M0tKejMBxebbKVZ3HbXGTEqMyvnfgXlFnVOXDuga/7eHn2XZdeh+ODBxT
reNikPColpz5JXyZVxld0QVvjbpXRbg3NL5XbrGj0z/FoA3Roha6AdRdvb6VuFiE
OoDPh1YiAyGfQhGl79E7zEJkJvL8GNw7muR9BbzJFtSClMYbTxtA2WB/vxO7Pd9f
dBofRiC9hkpA9RjQ2wYfutyFPVloqamrN1TA9tpq2riogrqex8S+fkmp9PCHGZ3l
FcfGs0nemmNsaD8qoIpAXfGQ+YBwSeYGMGWdzUM73K8SsirgwOt4OD+VvZ917Kc5
lZPkM9udYHmJ1hXtMkeJjrTIPDYnOojFP3FQ782/OA+R/Fr2PBrEHzWEJsm6zk9w
+m9EELXP83rmvTv+x637642fVg7EtwOqF0tyPGdU8Cb/FnC6We4EAVObLmJZP9uR
s1MxwjkThzYy7Dz/J02ggVOUx9d0mAwmgiSqZcASrI3adK1W1n7rd7fAf6Q/86wy
/sOpkJPuR5VjJpZHzolT8FlG1rI1fm77FPKJXRS+8vdQ0H9zS6qzaTsc3okS8ccH
Df9R/DqfMJT6DqwfD6cjQPAsyc4ezg4SpNQNrDseYXB0sTRvJclQXIocZ8tmfHjt
nh2dcbvgdpCiuMu1icOBCb6AC0bCWwuJt5ltsHpgsMhEx5+4DST4g+64Fkxw/9ma
RLQO3iH20S+tjv8RVVtiX6g17BvIRCcHU0a3R3lM73lYJurxEkjzGodL46CPrzG7
8MPMEBocgMPBYGYX28Qo9lmMgebutIgn6sJFZAq2qm1HVUzAvIMWLcXhrP9xoj9H
AL29FhGugtY3uP417cCTAT28aFxJPUs2uBrZCh/dims3S+T5VnX3DRr8jyou2BvH
NLfXlyttISTf7catJPqcJd09FQWik33W4trMesEq5FSDZLW4g9Xea62JNSA60hQ1
9qVV5etWpoex42MS9uRnmESpKR8SEJvfKMn1JnVqLfHzj6xbcOaaa+M7/VIfVBzH
lhnbb+kNx2j9ZbXET9KYj/MSbJvxeyXDrV0y1mDgEG0SYDbpYXxjY92I9UyRwx3X
q/qVn87DckzvqvuMZ4Vwufvnz1lrz3+vWuvG8HVyjFSiagfIOzD61P7IhXDuitHc
pmCxIY3P+Osz26CPsavVrBh/ra4nvOTrDVxjShe+S5cmmHHZTPdE2gNPR3tT2rJb
ABw3AfQHXfytt4UmV6xcrtc7HIjQrx9pn+E7QbJj1m+io4f5QfaASfrJhXi8OUgp
T8vsn+ikANx9z0gbkyFc3DfKUW4T+XCBpf6ZsZxKanCuZk8Zp1hGATFbAhjPSyEp
fwUsrmdINMcTsZZtMbI9fiZ8aFDiZxlr7G2BRa3zPjhi0VMvwfnEJ+QM6kbLYQAE
/v/1otfoM+w1FxI9dMGcDoPRQx84iyiGdUJ9mzK5qvjqATphHFFIUkOc97qRspqH
ngNNjTxCUWRQJ9EtC2+MNiwenJ/Ao3rAcpg+KIX0OiqJqjFhsqjAVWHgR3JyOXiM
W4XgHbR5CD+JCgkEBuOxbfGOWnnQ9pBNYMPqDe3CIz60y5oWGwh3WX/YeniCMOjf
YhKtHrbZeDM7UpzgCsj0kvRWPbKb+RbTY3JAWnxb5J36l46esbWhGB1rGVjuoOhH
0NaiDpUU0zSN920sgFRDZVSvpd6FOsB5Gm41TVc0TPXspid/KUP5ScpKJ1x7cI2e
jPteP59JazSODyyeRPO7CkKEBwCBZbFTk/XKB6rpz0RLE/Pc7A1Y6mjqHz0WY185
hmsVGfqE2D1QnggeCczKEwqaNEmtFFt4HImmAa+flVoNxh6+K45sDxgY37Gz3dtb
57ka0C54COS9zawzwiJ5v0bj9F7eeeQeyOMOy38EGkNdm65qYWlP6/saIapCutn4
nCNwTj9ZdWVoylZU5LqcYhpnT9OF0UQ8QGG7zZr93hHt0/AHw8PaYArGeeEhgjll
+7JtrpRbvaVESFDrpLKbZrpjSzjUFoQrZyeD15opeLF6eU5ZLMRwRZfr6KKiMMJh
4t3dWXzuy9pyHfu7snBgWBqydKcZnhmHtTwOb7NgAFs1V304HJ4Y1q1XcFHGkIaF
vJCUaDBYYeCpxNnenzTIspIqZ1FrBZhl9oQgZQF0hj38ZdR6ZdC0BOPc9ZKoKb6w
akN1NHg2ErAoBO3uI2gY0CSBQzyAdVNznmH1HMTGKP21jF1/SYTcMcbTwiVtI1+u
MeSJJMHn2u7Dq3Apb+a1aRRNh8FNic+D97waJbdidYQ7m7pEmrXUJTmwqqnHAhys
bSk1ByGqS5f4oCE1FoPW75lGAf5n18O69Cwal1uwQmo=
`protect END_PROTECTED
