`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w3kw/oyVfKHGzq+GF5HV6s2XTncmDrjLKfZBBiw0EN33Nmf4UQZgyhhPZdIYYpcf
3kGxFzVsr/vqGkcDNMACKVsOZbV2nBj9g5N0iGswcdryxlqgaTo0AhbfnWVzD0AZ
u+zh1atVejP74XHkL1jOVSEslzZ1JTEKdJ2kEzVp2FwdydQNM6mmLUFtfJXxRI0u
SaikIcf5b+2g81g9RjPdpDmsmkZarxfypSftbWDkf3IoncKmMVtRtP5pm9I9Epzw
LQ29pv4tKXM7PfZ2F97WD8SctkhVGaAroQ4X62fkcbamUONUXHZTozZBUDJXHeet
YfWco+ogTnHbRjSsIC9oHsq1Nb+xgTPsRJZyxtF9hU14L9JQ+XyiRb6BJRPUe6rC
2qvEAfWfpMxDf7+WSAiFvdCDakrL77cJKV1/j6j+AMw/kWK/eyDwEbeiHVqUxnf7
4dlDOIr1+a93bna0x4qg6eFishzNtE8RNrBjScp2VNw1o2uDjSaVdMea4a4erLxg
yMIFhLAifSd8VkrZTxVHhnF2Ntzh7lbetUmRKfx4tGlk3OYfa8HXQ8McRSnHzGmn
6L09EIktxjLRsfk5jlMmEqEsqPtBpyFr86Hb4MoWlvpgm0/F9zjsmFkVJJblRc+V
9ImmLWrLcL9FrUqAPK1FbWqdoHOUV0Yhxvn+Dg2aGn3np34uoXAzdR7GzpdkO0XB
gDUevuREXvXMs8yKZipzknCHoDZ+AIfIK5/UuLZWJLRAxW3Xucc5o2mMS/m06sKJ
kOOAJuvaPpgivGBgcjE/4H3OUCbNJ/7PSWvDypmRFrfcOhBozyVJohCMTOSv49xy
PoJR0IDoTaLHZh3nATVBsUCr7g9simfwIgTcLbJLyeiKW7tXXn5dU05qLNURGLZy
HBzFd4i3jVYHFjAR53GkVzPNyeVenGGIhQe8f+r9sMXjiyZ4rZQ27DZWc3J+5Aim
7dh8pWDHUGOF1+4AyELk8WIJwRlX1QTuZG4I7Qs0r8+g+BJfqr6tWZqcmvPfuWXW
uD6OCD9gfvms0R2Ge1l8X6PCPRZce3y98qNp/ewqEzcM8aANit7dwfifk4giV3Gr
UHBYaZPzhLn32IoRsh4s6VbniuEnuThaf1JdHSmGAjsemLyhEr/8eIvnLq0clT3s
0J5ZhX+OYJEbapmS8iPCnCm6RAmZYnGXS4o9UsRMa605dw0lpbpKaMfK89ERPdV5
/19fuwcli+hZU86BxNUZdfxhZE/VszCSUk3STRiX/5Fl/wRx3i0kS+nbEu9Qg27c
X0am1soHg7I8+/C8DOkBFybFT1vY2iNOrC8JQUC47ppWiqo9OhaP6kLkUYpO+JiW
VE85XHsVQFUdBM7E+ZU09ZGX3KiTi31ci1xIgh3N/WBtRHuuFzKTg/got3h1eYcA
rm8cvzsGiF+umXqq12W4LL67+boKq+yUrQI4pImbPh34mf0/PhDEBuLccmetaKxN
UYVZBat9Am40MN3BN629BRf7IayaH+We+D0tXT9YhpxuRTbunbHuXeSxOK2hw82z
wlV1/LfBWZx8s98zEz+A2qdLHJ0FLIbVCSfilVQGUu8Vxra4N1euBxfYUalguUn2
zRXAgmjuAcWvvH3xJe5gO597LWgNpDNOhsFQP1nFcPU=
`protect END_PROTECTED
