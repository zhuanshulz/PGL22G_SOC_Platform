`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wIzRpLBSFL8mDTsnhLCINukLpDTZl84319qPPMYjb3PjmD9W6m3Clmb9qU0dHD0u
hwwhUEL5N4CDrFBHq+hG+ZYbNmpV6UGgrz5LWdCBtSzImnVN200SZnjatIgeb5J7
y1Mc4TmWQpsKsW9G0ynOo/fpmxNtSn/YZWiihBQ6g4jpSzslh6m6pPtYPUtCY779
47HlFQHKxGsEIBiNJUsMK/UP0Lp99Z9LvyRfoFOKHjOP/G8c7Wpdz201TAlx1n5u
Mfv2qU3Xr8cCO/tPcPySYagYluD1ggSz97FRJkeOdBSULd6WDjJwwSYVusXBfjjZ
wSzF+Kz5WTGXEorycVAUWt1y16WdR8BXk1TdUEId2bkqzviortxzJeoIH20m6wdA
AGiFMuCVvHPJuk25He0mRYQAwAjwpKO27Fboz/Jz4svBVjRrdyhwV0+jq0NSS9hM
sIaKvOemV3sGR1bzVbDhFWQ+XybjbPlc/jmWyOttjEsNYAt92/EXp5JGjjSy1aQ9
VZnbZeOdS3tDZafM6aJzBnGevTd4ECh94t9Hjo2xOZXIq7D0KG30zP6tnW8VeYOa
vcxOyaQcHLpLQ95kvPkCyKcd5xbM4R0FYHB6qs2saCIy/SPB0c8gJz1uEK2dBLDk
vNWT7Ot4c+wnvzmBmVwiFUQPpYJSOqOq0JKqBlwaQIQYByVeWU13dTiFm1Jvs8gQ
oX4grqdDHxZIExZqvlwfsxgiTfbR+yzNAwxcE2Age9k27Xfhz+5s6pEDJLYbegfd
RBW9Fy4xu49QJ/3w/JXWFwEm20ig6hLiYQz+eclVE+YC2gOTGD+MERsyBPaUaBG0
JRYYEctrIxxoh9mrXgPysLMWwbFtxEHzMn+ResENTUpSuuNEB0cWNVAZOAl4ipT0
41LHd3KV2bEocnbAimS2wwPh3+UEvviQjelHUfAXjpE=
`protect END_PROTECTED
