`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ze4Iv1hifJkQffIaX2/fr0+BjnjtvfKnS51jLjVlqP7Z07WRW1xdf9ZjdsOX8UuO
R2O0G/cevGwAoI7OoVnmSf1qY2A7T370jqFertAUXmt+MtHSp0HlOU5EMmPgHGJv
iNlpey8+1cFZw0yA5sCdEBYLoKusAYxeIBQ0Fv+Sybw2Yn2AvZe+7s18fYeSoIhX
Zf10XTwYOjcbeSn80rPi3rABmU1p5jZs5pcxdzD4OVWVkJM8BHqSWIaSlNTiFdil
Xz+AWgoKeu8ERy3ntfkIYulqMy9dwWmRaHncSLrS+IGMiuh77Ci/jixfkE7i9YWi
bg45db/dwpRKVdwIP6rmcTB4KhBKmkfsAa7saQo+AQ5FoSSw3eBMdbimIVzQOv9B
sD0vRP+KHnlolE+Yf3OTsKXbvN9BluST51H0+uBuYkmlThjra9cR37n7Ib6JRQLN
XH7v5t4tfxBR4MKIlewnNef6pLumwZHB7ILtj/0yEqIj7EaEXBDL8h2TWH+0+G32
RkWBll0xqKjPwXKcXX0zVQz+IfZUMTyDTB1b/aNxtuk=
`protect END_PROTECTED
