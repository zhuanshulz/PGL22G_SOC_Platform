`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QXnYjbaLuzulc6ejbwwICTkVYGZJGSg4Gpm4jpxQQUietBZMzJ/g3qmBWjQ5EzMR
E/7kAJSxsuchiO/q0BVMTwhOFqIue2+hZ28rbNjhTUNItb6y6aDbFQG16VxqjtIi
MbxpXEni/Gg5Dne/XyAApLsHmZfvek5M8+6B61EY5rOzzj+/Bk+miFDAJGrIHS/3
k8j8PYcmEpzByEQOrdD+PNo77YPaYrIgpyxF8PImloHhqF+eoCcoll3A6ab3s7OD
mUsZ/R4TPQ9XzegRPPWjP8LpUr1BA5PMrNj2B6WM7BNg0oZgr9O4zlG3yg0iQ8EN
ne8ci/vAQAH7a+t8sYlxoySXfi7rOKyPiZQmv84oIwVBrY/IaC868hLd/XTXSIbc
Cs8iYqeTiavkjEHrCIbW1t1YoOjQjP2C1fkbA9ygm+Ru7je85WS9TE9EpWYhkZAS
wOxLg127njtrESgb1OGQ8dLBPrCG/LTRT+NA6E9gp79chDQSdgeSKAoRCkY34U5c
Hv0oDpgFQQtdV8LI9ME+o2ON29JXefZLjJQMK132tXK3JgyOFdEMvL1eoS5qRz13
laHZ51y9onYujtugE2to0/zPmQZ9TnSNsbPGKldD3uj3A369LbijSsaq5hcdI2dC
ZSc7//f8FZ1ay8mnpUaf6n1QQUzU9XGuDJIImmydfpNw+uGikLQ0cNvi2JhmzWcU
sPjEBW+1vi3JeQIoqNJWYPCW8J4y7UwNw4S5GjhUqCMNQHO/ZZRNdjrD1cyKjnQL
NpVjTsW0JJlGaze3HmWQmPdb4+Z5vx40J40i27sMJxE=
`protect END_PROTECTED
