`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bZGqLLcQ9CyLKT9OlDPXg6k4a7xISVe2eEK/4yXo7311meqqxQMyo1HWLRggqo3f
pAsHKLY5Sk0Efi24Dv4HxySINK5yHnJM6zEFiZrQfv+cUvaFaf63NyIdOz+Cc00G
IGGWEnVYfQkM41Ph18cGZPA9/L/+k+t93eOkKv01vm9OzhEwbxGVHFL/YUtZ4rI3
a7R22Mjw2l7GdwVa49zutMkWvRZVRLp3mH8+jNNDZX/kzhrn8TXFbzAZIycOym/m
3hkO5JOmY3PPDQcSE8ONvEkmX8e+3FeJelerIeH4nZZY5cg3785meWe9M8InKg+V
idbq+upQFF2EC1bshrlv88bpcJwU2vVZRdKwwoDKPXJBlCPk67Pq9whvk+e3UH9M
d+AM50+moninQQyo1FysizU7eBuycI5WOuH6FsDNAuA8N0Y9E56nW6WlTOXzsthK
OXQSKXTPOJpvcVPl8TYcyDbGUj7H91rKcPuMWgijGKDzVBlGlyaqenEMoSnOsIyw
zw0SgNbqZwkxO8g7IaK1OGMeYkYh7zgKUC5uOHP0W168Dx4eMk0AoCE/kpBSmSr6
wkK3GRvTZfO8lniNphIgSxFb1go9PDfQq5TVwuemfr7xOIeDQKgIQ6STvYXVpHp2
QBNwGCizeOrarKQWEcPmbyhdR0l0KwzNmwTWRrlcz/H5L+WGTcZC+J7Wblxavbfi
lpMT8bstPvOh63dHN/MVnGrj1zWpqSVX7ZROKHF5cWIYvTJeueCeuoi+tqWP2tHl
GEBeRQvKYFO4M0F7Fut4OPD1JqUrxLX97+dCEKAHMimClHDNbd1SBzBN65LkklbT
ljnPMv5BW3Y4FWCBfBVgacJlpmAYh27IBtbILCPYxRshPoOl/43Ywqbd2q/a0SyN
3wAElctZ9OA/LIm0xFeys2jA+aXkGvbkpngQRPbf3gmiMqewRePYJ6cDZ4Ra3vJI
w4cATeB414LUCi3/6Sm0JzmGRIAKDeA/JuitGhDK3TvzJscSeGXaB9XtmcFi8bo+
CaEKlV9Eizh6CVdnRNt5zg==
`protect END_PROTECTED
