`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/eNUGXwoi24CI9CFH5aJYZGChQIk2QfuFw3xUyyLW/wrjm+wfQ03K0eP092IcIoC
tVQociBRhnUnCxQN/hbEBN/gGpCGEMDM+khthC3KbXuVM2gY1GOa9fxHj4r3wRYf
eqnIlRRDYzux6+Fmlo4htfEwslzDlLgaC9hLdJvKgFUH28Hiir1FNkHSvShEouDy
8t/XRioFsimR8nlHPnE8O4xnOpXuSTIvH57ydpTu0cRyZmq+mhGbu/kWBecxVkK4
Jlngq5sE6c0pcgYvZ5QfCbANy+yB6HtoCP4yq1xzV1Z8fhjHtaqPMixAxMIJtdFB
DV7tnAO6n9f6RM1yPG+USw7tc7RTDWc6luAHw5RAMrgovJ4c2CsRKxvGaCOQmSBG
Ppiqdt8EHHghD7CRbXrxZR69TIN5OWzjeWI6mxagISXfFne6TwG4c0H8xi30oKG2
YzQPQNUEFQSv+zSIWku46Ql5mcfji+/OBjk8ILhqBMG8E8ptkY4++947nN2gU/74
DQ0AAw1Ec7rmpqN2SRE5ZUXykodoCZ9tINph3Ke3beqSXJzy5bDHLPAo52NB4Od8
6oczu2L69sjssmzNuFhZWpTl2RFDRhKPR3mLitGo5UE4npy39Z3xmsazJd/1R+ju
rW7/y9p91REnc5Qi/Jc0ktbYkaHtjauseCZU60VmOPKSKUDGFCVFZPCN0qqQhLja
/tO8ti1Y22YBZH4SB+KufZKqNKQiU7U10fZgs2l2SV4cUeUWeS9WWoAYT/sCGkRl
NfjWwZ+anfMzI9pj0vI0WVp3PtsPhuszEPSl/cMRCHURcpMlWkUWjgt7CoNfwajo
wLyXMXQ9KWv3tYXC3605mVduwVxxfAPxw7qd2PC5CdQaAOJ08QTXJmAPxOhc81RH
7fVFS2ULeVu9K18OTkJ4rH6d7TyRsFyDWkcKwQNIpjIb5evQhpizbQ8bCDWlRjs7
VMNklYC8Xk1yjUkpLufOZE1eVKwUc24l+lnPF2WT0g71ODWJl/4JP1DKYiZDEPIt
4fLsK6vV/9dBKfyexzrr/korX6pICyhHNStd4J2TKUDSwwYhCKwLF8LHcLu6nwwj
CdzyyJTtbqC7b2DkvBU8DWPK4hE5+utRtsUknaNGTiPWNfIKIcy+k5JhS7ljJk7J
Ags0/Dq37G7yjy83DGuuB/jgYYPuUt+An5UWECyCu5RSSyGzDqEe7VmD/JFIsTBX
gJJK6Bx+WJCb7zjaCEldpcfhN5/R5pPxG9n9E+glorwypUCIgTLz3wyF7xzX5HKP
CqR9fcwERavGudzzMqiqOJyDW/9kYtGm1i9WAMuUlPDCklZBjnNXSQknv9WA/wCe
abOhLG0l1SnxRCElHeD9kPnXKKoIxp6P5LCA2MFCZAmLLUP00TEVFA4ww7M1r50/
NVY1cpq10cBHPXmKpcIwwMzxKS0t2zz9pXTk4+zdamK2Ca4ghIsO4RJtSJcnHFz/
nKrXVg7MVM6UvdSQNgr+V8oGsQJML6suVhkcQeq8gB1eCvjirjkBEnk8Lj/AN2vP
u49T+b2ballFksHQqLcrxdnYNyc4y8Steel/mrjx4VYQNXWkkEyQN2tZ794zMew2
KvVkVU7Cnnc5Hp0dj35fH5NmZyF2MUYkRUbc3gNStjE=
`protect END_PROTECTED
