`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s53lMJaPnmhWhrz5YHWYwwmOnBYwB9oy9q4PesDJaHKHRq/DqzDqR72bh3+Zm/G5
yTcZk3FQr3gybGM0tqZpp8hRpm9t2Te8x2qysxNzXPDn3c1h7NV7oobcc1Cp3p3i
AKJ+yK6EPF600BpZEfsUQ9mLKK/39Q7ciRXdaedLSIINGo1Vo23uiEYESJwkeAVu
zNHy4k45tZ63X3P8gXQH4cTJjWX+5yHkQKidpGPbPxUMl7Da0j8dZhmo1EAhKzf7
Ydcs2zjhAmI5dQP94TBtt4NBnOMJIPSleEyeJzvSdsPDWb7u7zO8CbAfDF0aMYmC
7d5YjEi8gJ1muFZS15GvE2Et6YaqKWMPDBj0huJTzY+TZd7DY5Gp8qNceTbaapz/
h7O4m59WXhtFa4eTOqYJPntU7lp/HmkMra7xO6zIObLSMYBWuStc7S80gez4R6vc
r5gdQEdkj5BbpJf/+vIFNQSP/1EOzPOjlKXKZcV/fIe6ku79QJuxrqMTGlanhZJK
pCDgJJY/LGDxQ/mimGcyWQ9rdjfYvjqxAa76XUBF4jYQibP/H9Dv7x+S03YHojXV
DOe25opnm7BUTxjs9sgNR10pO6ttC91vpQ9mfTQvAk9sBIC3SopBEjJWo0ZHTmVG
LEuhYdinR5JOLV7/3VXFnzTmRIuoGI20WlNiuyh+DtNp6jZiIm21k11+2/ZbQTH8
UeG5sVqLGu+xEbitbeZh/fKW8ugpBUDFy92mAQGFt8P9cHdNPlA9RP39++WydyZi
aAuo8+srkNk8GJgT0l5Nw4sCcdaau3VnwB+rvVYg7VSLkgZ5gcFpBN4dBSW04TLL
tYnEnQNVq9z9jGLnZRTGP1Z13x9UmbUKEvNymwf4z86gji9Bkqnxh22Kdkm54V5b
PXp/0ImA6tq92QgSrHTkbKxVzwSXiH4/gVhRnN2fOhBtb0xHZ/7WfMoIWYtjCESG
yjtnDAeMDVYEM4UF/c43svOze+Ve+S1oN7/HXpo1l5De1Izp3EUPDJbqjgGYEPTv
2RoOdS8auq4aH1Cg9KpMt+OR2BlJD3ha73/cqjZKNOTIQUCYhtKMIrHFJH4cnU+N
OscTp2Pe6YY96bYPJpydc+XGMsZHofN1/j2dJsfRTQXTJMrdBPSrai78MV2JK65j
sa0On6N9vYIViN98ApPmfi76tDbbrq/k8JZsj1SebDx3v/xAMIMehEEIOwGRpPro
fWKfgZdxlgwGaC8rHNoAb6o/Inzy/6Q8DhIvu2laN+EioGTHe2trDo3XfLyjdPMq
b6yfAkXczSHX0aJ3acaS8OASE7o5tK3AMIsqG94bla50FE8xirc3j9y680g8rAux
4unU9VwYfs6RAkIn/RbwqsxqwNbBhc2IHNKkIUJzfLALIEY2XDivbYcWWW88dHEV
hy97+KWq8tfXainB3f4lj6ab9oN6B/tOBs78cmN/++UloUvlk+fgS0kJkcMAPP0N
3ZA83CXtyFQImO9fI37KvgRQVxGimAO880QYVQH+HL/B+E56/nBqZTKbOAu8OSxL
vkSiwpzM2eY4bshOez/+aznXbTfTT5yIFeW/dOGccfEiZeTG5HHN03bORRhcU1g1
mIF9TjD9dRGATiyzXi0RZwNe2SDbrTrcMcu6MmsvdX2EHGGE2qq2ESLf5ZObngnz
GScwAkCQrpOioA4e5R8NSWmdLJfqexUOZouob8NK45uPbgTbImOoAItDGLD/Egxq
dqAHu8/zwGzECrE4loUHg49hMmsS8i9p3DO3+dXqgpXQBYKWuvbTwV0elGok6I4Z
AwaguY3S2GNGfLeFRKnSoBq4Jx5ZROFQk1ol6pCYmo75ilyEJ3yISGzou7laWRsH
oRW3uGHxwAKbFGjnZVGHqWswl9aDkSfaRxQ3cbtD9hk5rUHwXkNTZADV1tGIatTn
7d8PfrcGZtHsxD9sVhbbwzafcqYRgnMe4FGd+z2MT7aVdnwEPY2sCbAVk5WBkbth
t1SVRR+SKga6s6xNbrNU7JdrA7bRdKH+I75ObyRbTeG0fC306Rj9Hvjd89ydhqst
/kVCDoiUjRTujmIaw4H7CmIlVRTtrQIer8rsD5F7poIISX9D46FLmN2Pw9w0JCB/
TVqACJdcWwYCYcZ70pxe23DFCYVVwS+JGi+E1TuKCo2KyXNb2KF/ToPufnpssfEf
n1iblsT+mwTvRu6Q8wYDyBp97Nh+tZI7/d/3f22hr4JML84/gVpH2t275t+rS9WT
8ryMs+2fonPLjOVTU7LCMJdmbPiO0V3rM99V3iuPH6bkvQO1ZbW7NX7OXtAJwv2A
1f5l+grTWAR5BkDk5RmjYRFqG7Q6DKpN+BLibZCMXiz9Bp6LoPpMsSNovrV0r6ZG
9rCYYo9vTuA5q298BsZlsBVrLcOB4u1ggeHU5g26cXEvz7+fPZ2RWpjfG9Z5OIS8
r8KhjaxnTD5+jD+BkYd7M2Bg17zAJHZj5f+oB/XXw7l+SvMdl0EMnRMcOpUzDfTc
y+f6qJq60FPBCyunpvN8cj0KsTKfJe+ZnF7+GTScMRPtL/SuNy4S4/OXDw6q/1wE
Gd4z+Gc/8XZKGaKKZzbQ65j6VgUb2kLUNj0JOCQpmr/T5nDMoiAsAQ+QZTF75uWU
Iqe+cd/6GKNnY2Xp0MLO360ZfhEL53XXIO03hi5qZtF2N8QLaPB0PjexGTJvbwaa
DU3xpVlBalOmGFeQcPlFMk4Vql9txNlT1OEhscXYBMHTgKVWsX703frjYVMkXPzE
VDVHHM2c6oK/qaLr/uitU9U8PJaaAuJML0851j/+Lu1Un/ELujqyCuWxqDMfESaR
NB8pIiqtk1FY2lVixrdRy1udJ1kKah6qpQxW5jntuic1epEJS4Dl+C/fVDW8oqgi
uD8LetPs+idVGd4nY+GikLjhJfWGheKhJf/LkhOwD/9XU+tzOS6J6dvdKDc09UNx
8Rx/AkrhDkjiF4rJom0Iyd1Lzh6mOAd+lFa8iGIk/HG9x5fi3kfPCdKrWdVeUzsy
G/fjqtMTQuPJnVvm3ywDYqkYnwt4AAA8pm3QC/xadjXn1Uaq5tHYrGFI0NVtV/l+
fB5vl9TavyGQrkpp37EGBwJaeK9oTOXvH0AmiS12ZBllERipp6LanCTRSH8CA3g+
Dw8xakBibo9yemcoqNzJAQN7HYjowlBazrFRenDGpV5ZWMODqOcr7Cpy6zNMADL4
hVYz7hGmdONut18zaDVLNlXcqGetNqljef8yXpYNCyRIvp1dpNvMEG3aFIX9cM+f
IGzf/kk342/cCKgifb1vpxwb69IoQcdL5miSzMuFiK9ttzbJ615U75oTzV77EVjl
soO8b+s/odnQ2/19z1oSY+4Ubo1W/BkUQRoMvtXXRAaKp54sEUdeL/RASn0yj1Je
ruwC7jmZo6kQXe4EdATloUnqQ73iCgKy3/NnUAr/h+KQsWGosvKzOTZl+eCzys61
+mDXheI7hKT2ctdylITO1134lCK6G4L6vdg2WHSan1uz16kW+pKV70vFJ+SvjXY+
vMiQJ+O+i+PtmCP5rkTEZ8+UYIIRGiWkUxGU3AvBk8jwKTHWRSI8HzA7fE5ILDln
PWlsrmskYwq5q3cDP79IigDrBQx+UunM/Xb/RqqcaqsQL+VOsexBsYatL9EffkmY
koHLflXZrJL1hJh3oLOHpP9C0zI5AhsvueFiXwEBJvH4AxrgqqBmHD4S3Wgegazs
CZHWZCEkyVXxfNwogjIgZOCv1LA01jSUpuJJQvfw7LhJ7euDKgubi+6fSrO2akTZ
f+MDP12OZVCtJIluKFkNCZYpoPVBzpW3Tfm4ItNaF6ghjRjvVXqKsVpcNvcSx+/H
Qvl1z8J99wxnm9UVIXepnhxpMH9D3LeLG+4RzjmPbbEY20aC6rRz4H8jHyGLhq9f
eBCoZIUFZgiyweCeW5RREN+Euxp5tYvexnPM/E1uePtMm6EWfn0lpUQocBVPwGUk
S29sGLxS4xqTXlinVUuq6W3ZyvKpFpjYy2iKX4YIi2qDxVAb9w1mBiO7qsMXwLFL
RXP/hiGRutEo2ssF+eCoOOS21ANhzNsaiDXcjWI5fKxyeuGRnYGDbarxL33kMt/V
bMy2tFrujKwdrA14qeCMylSYf55fW+tgATM3oyGxIb+bk3o0pbF9k2fknW0V2IkI
20Pkp1BIxWsTa4qWJpHsvK0MAKCN7Um1DZSDwCl2oMCz9NMAlUicrB+zN91S0k7+
OAaF8xI2S7TaLKiWcu7IuX3HlLiZHDQ95UJHrRbN5pmAlIULWW5nqV+RpWfERiRM
wAiudUOmajgooWeu/5oic3DExBE0KfOknLQsFm6dx8Fo4pBrIlJdJnfeGwaHj+C7
heMKyhIB8cU1BW0LmUCcSf3rpNHXtIJpk0N29pQF2dt8GgT3trLrWazMHwty/Z2k
7lpwJHJsAr1S6ZhdJzvQP9BZYCJfE417/3l7YaabGSyEURPjqD//6rVs4QfrG9ax
GZroBDgHQY4qexnPKqotDbYfKt5YP5LLVac6s+Gsfe9trWiEU/Gx5plbT1f3qJIQ
7lnhzyxoIKq7NMBvIaErvTZXkoQAuWhlXoAsTl2D8cQa1va/zn/qj2hrWvP5ope9
TAQwEdZYgZZwK7f31QcvS5rXDpULD8ryQxEQwG0MKej9e4SeXkwg0CpDw8DmOlF0
klri3RzY5C5gRcbhIAVr43DWa/rMOr0YLb2vDeqaAEXSAX/WWxz5G1VtL3AazIFy
YVCLbaKGQctRAd3N/NU3z8MBhu7AywamCZpd3isZ+OnGiVKkBzyOW3263VITK1FL
3Tf3OoE629xBxmTJWfvtNa0/U4CJO11f7NFHXKLfUgJRSzDDamX9E4EbhmVjhAKn
xogPSX4mfJ7XqPSzw7DXkHYzpqrgjgWnG50V9w5LtwljGION69qajht+9K/Z9NBs
F8K9Llq8dGuc/GyW5DQDrQ1ZALTvtFMNi0+jylDN9QCgT9l/ACa6n5apJ6U0P5O8
hslH/yR8OYVIumRezx7nBhqBOaacEuFhwpXsEjqGTOIcjUG3fqfYNCeYYwo9Itzr
JsJi2i3H0pbnPAt4rVBzCfRmeYYk7ceZR9WrzCA/GTKhZONZiUFTF+Kn5u0q7lpg
x7VR+ab5Mwcs+Oj6+Tg1VJs/pHk4PguqUt+SwOh+HmGrirTPxY04IPns6flSUW8h
rbki3ibbnSwx303BxiDz+qiLDrmROTXX+ggyQ5BUZywG3ziShBxr0iBFEvgDUekQ
eNRpRdC5UkDOqW9dh42zeedpk4dH3vRVC8BRh6//mp4E9Cmm4Iz97xfv85jbiKQ9
FtMP+i4TlNC8gb1uvpAVVcA85JJOjP0+KXjoF/inNJt/YfOYpJQmcZ7f6YEcNN+H
IG6KbK3qGG7qTEONRSY8EzN01TW2FpIViGhmARFJipg5Z+dRrJGt0nTj9+eT99DA
U25G/IW09qgLOeBpF54fIP38tWY5zEmZbwM4rT0WF8zaaDn/MAaaaaWh3ZBLJoxY
PNSp6yRpEpMzUtg5R0moeNQ7gJf9QBnsJe894Pqrs1ybEf6lk2oxVbwkfTPqtLmc
DKG0LjCAk2aUN+LLXcbY54hQUNlrA760CCWItjmZjmkID3mqr8NSZ/9ehwtBssl0
wYALeq/BH63EqQSBZ3wRohDPU2cHLQ1zatcJpmTQu2OEVy786G+5xMvjLtt+HJ9/
MVaVg+MZTArZJSeECHp5CTekzNXDsFAITCGQx4n8dX+AmRHhNthj2zICetIbwqpL
K7Xc/xuwTJrGueBsCvloHHYFu4D+VNhghkNMo6qH5o99t/ZAJG1OIKkAb8Ita6LQ
FhbNwqypg9kRuKww6ShHoTQGiwEVfPMvSXwNevmfWeGFgKRyJDbKBsrR16JO3fyM
ohlSoE5nR+46eVoHpw8Fyd3/mPqi6vi7SEEkzTsr3HDjHyeHSWLjXddF3uVNLg4N
bTRsTZVD4jN3AdzTP0lX5mRrqeBELZttLENqISj6moIDPUUthNdgkShyvziIcEes
dBmMzrgNKrfoCAWMZtBPJzWsKJ5O+e1H1SdEzRhwFDyr15uXF5Tuu15naZiehgTD
tVwH3KjGTYYepfV6Sm2PNvbPSS5TZ5WMbbX1lo7ylXBSmWH+OZLsYXgU/OQXbjSN
4uIMrFSmNE5K6Ahq0Q8D5/Gzohxe8q2AnDlrSkW9rJ2vrm9Dw227EdHZv0do/7rG
fkfU1R1VmQpGGu2QZPPO5y4R4RHc6TbPFUWCHMksgNdi6tFhTl2tQPAzNjf9x9A4
T9yn9RSUv/QJ97x6jxbieTfmEDjt0F2YT6CfJKUbTFn+pt+RWP4fFpxWHbunxmbS
NDZWDNpz76une02SDaICruizDwX8JkyXTN4+yueGOPq0MZYh7tP81P3QediJ+Btk
DK+IbnACMx+r9XssoLI9mUZqhEdNpUYMx8blzmhi5Puzu17zpKvEngEf6VYRTLa2
D7s4YCX66D5lv4VoY9skkFpAdR2pinPIXV0eYw0RT+G7C+/9WRIl1FeyKSLpJuA1
JTJiEg/tkeuWYsSBh6iVbZhWXq6eOeoO1ASRAe1VB6c/VL0SVDjsvPP7g0uMWsyO
3s4xw9y7tJe9JpwylQM4Bot69olrOAtRdcNUkZT8eGTsL6bri1WjV/SYXYfLQbEl
BUgycjri9D2THvfw0JL9Grd0IP3g7kr1S9kKnEoXeYh5tMAyGpw1UgcxxtYyWFeG
h3oSp5FgwvqWp3ZiO0W2k1AUvHpY0O+d40hg45i9fQj/Rq01uu15Bix/tnkVVJc7
KywieM4K6ml/Rl22H9qMHC+XFBoFusb4M/N84aHnZNpP1SPBipsA5izEjEfY1o+R
1EBPCQg1eIpT8h1A34CdRdpO3828hrlK5T3tp6GMVNE/HSS/E5mR8omTmWTAKNUJ
rYX4YfE4wViWo2R+fMhv03QUAhTV0oFT3qxKVfJ5UrvUdXSOkqd2cTVhqe9+Iq8E
vpLPEIheAJtQImHIhBeL5ade3A0fK3CrlhXXbZITt9CyTADNhL+7pCIgL9g6k+jd
PcA+0Ptx48x0ZhndBXRhYQFSU5MM/T27xKcRBl3H+Q1gvXRtQNdfvkcPe4Fy+mWL
NsxpOoqqWIFJZ4IfDSRe/QCNycVZ+XBOO7t0WHkNDtvA8YAtK97luS+nSwd9DtPp
lD7rRSLOk+dkEl9NXdEOCSS6Mut5KUtiDHlrg5IEsSk+7UKnKHSji4rtR7NuPwA0
FY+IOEk30RQZkaDTFlrBen+ujdBPH90OWJJUNVspRhb8x/SkCrL0GrfsDdAutkiT
a8PwM/6Wg8pzBpiKWka6BLAj973l+YJzwYx9PImEEZY5RujBgyuhF9z/lygh4KVH
nfeGBOdXNnqtRpdoKiOLqDdxyKTToRcMnQQCwiT1W0YF/JBalFi/bFMrIRp00qJ4
6V7yFxXSuUh5PHHqKWK4S1kPbLjStu/oPoND/mXSRenE/EdGx3GywYSOximgDw57
3yFD6tbRSb4irLMcz2oo35AYaNxkQArPoMdRmt3a56uzK8VyZe1KoeoGDI2kJwRR
+7FQiJeIydOxDKLpoQmtZu9RWcYtzvZmyd703B+9nz2msXP8kbc5lIkUP5aZgxTP
/1kpWfFCmsXNfGIL7xjyjn1o05soh9iv3S3//vD2pAIkPuO5pD6nXNga3oW4Mumz
FBya5h2cnoRKa/IWEpLtcr2GiRMBO+jR0G2Z4eQTMlv9DPka2iH4WgKWvmgqN+vn
QRNt/5y3So1tjJbyd+4vxT7sTMiBYh9DgzC9jDM46cx+6ZmT1mnnvzUhAPwqfy+y
RxqDotilJl3QsYgiHos9FUiS/bjwr8uVHw1B/BWxoeufHIbjGN6vVvhR7+zxxMwB
5AIq/4NeVVb22ORWOuQgOO3tEQWrbDfTCX0zuU6N4C7o5T72E3hxG906Ui2InrTO
leIZUeXE+oS/Kg+WU9cCklTZwylv86/a4K+vm4RllOw7DNPtYDGB406zHWb4/EB1
BPoLd2KujwOBz8aAYNuvOdlUCiE+nu7iheIuYwrfJmALupuPODJjQFTKTx1X58Pv
V9jEwakYOjFHz06KPnsl90xMW4qGfBkKihb28+xRwN1fLTfaECQ5vVVjTOAApD5p
jm7+S9WZcxE/OqYKv1ZxTkJVgTtk69irsLcqIywZK6LzLPb1NEWF2R10FfebOWuP
beH5oHwkxjuhmH8O+GVJZaGxG40LnfoKBnTDh8Hcs3dNIfXUJ4VNkMPm1LjngiZ7
zaH7psbVbexkNdq6bGpCv4bbTezTJViadk7RBRR7l7tZa/jdgEtYQL3irOpcz3fN
SDulrq77agcAz2xyOXzhyiI7FrMbHQtfv0Ycdjya2W3o9KXnbBq0ftxCwQi//FRd
7gRXUvXTHwwqbyucdZQPjrY1zG1gbcDnVXAEcVldattw7JsBOsb8Uv+iJJh9ZPrw
iPSvcmG/7WvJPpL8eYgjEMzJXjgpFz+guprHRYQSeJYu3vWnyYtQEZwjM2tR8Wh5
uwX3WTmA0S+yzjQO6RceQl7D38Mst8f7hDNUec+vUTNv3DedcO4eKnAkh4KO3AXN
SH8TKX+lu358c8MSu9vtRpAV6SQVGlv2aEAebq40wYnuRXEw+UsF9+tPRpWSifhW
orKbXQmneC22IccSUYZ/iKIBhs5S9d01MRRda4pTeS1KE1Pzomvsacgkn+hm49s8
qFFbkevxvEsPN5GfQVXxnY0BbUNFOwHf/vZ5vhs7TTgOXn2k+E+juVtkrnZ0dYUA
t9I5Qv0xvqyRKbOMPqq1l4nsQcGhVZGYQR4jzaSisaEbSIQjp46DBH/cWM7eTyk3
aXotuSeQ+EAxKPyvyatlE89J+rS/UtSsZeEQMWLBVQdCWEsgXvBbEkMBhfYIAce7
7sZnVT2Udjqc89kOi12CfFLO5K+wsaDVro5IZ2EnVVpoObBx0+lBpgBoAT7nlLux
5VEl48vNIe5L0HodxZ2ay2SOgWkh/jhkdR41GHdZUAV/nAjYgO3KpA8mmsLb+UX1
lfJjennX81UbqZ2g28oVuuwiyfd5K0ko2ZaEsjyOYDL4KXrc2zmG/0xYbHXRRWjU
QYEIBIIYL3EyCwHbcEymzzFbJybF41zIueXrdf2NTxZh4uBdQ0cgUkQP9qLy02b6
1PaIOmezH4SkMBZocsl2UuuQbrHlex9gNWZmTO0KVytTAhp7i6dMe8dmsY7zziUV
ySBUQRz7mIYEdsB4OkHJlxFSql0ggDHUZe4F5wCX4A2oawBF68EfM72OK4uHir2t
P8QwlPiiBbsC03nsBqWI8HhwZIJvhjnL5+SPFmV2uuYdJZkPvNC0y8TVsGPp7Hz6
XocFNgEezDLJnSLtZchqbxlw63ZDlLtOTA1DsVXbcsYtKTC0SR6p35EnLHz/5CV/
gLRK07+OvSS+7EYZploya7CjrJpbv4EqLDih8hFX5Mtjrs1/nCdD/TmlHWiB9mN5
i4xV1YQSN29JpGTl5M7z/5sNmrNNhdcc6odTonAEwmugZo2RaPGgW/bMO/peIIhs
R51B4SrgyrteGNwJ6pG/3KheYjNWiDoAXn/0umsSEV+Ur3nYSx2RJ4jxNShUjKR9
NAatS1RvmgqxO4b12Fvf6+zclU2Ubw0G49eprOksFyR48xr1p6nm/a9fZcKqcbfG
O2cNwTh4iPliMMZz/9HpiGhm2WvIq84zl4KSTYOKYKJTaOOQvoBBUne5zMPXANsy
BCkOK47lTqg1cgcwhtgKbhKrQxbpkKV9Vzv/6hpVh5Dj3Q0djmdihLyfElPL9hU+
A+zl6Tx2DHCYFAjc14JCDtK9SC5u2VBOBXa/XF4fNNQG++SWQhcyiHMGj4sydq6N
KQgH/zwEDNEGfmi5iVZAuUxjG+e1ElLDmHnNJkmGF2CJ9+lf/xjG3kipJTeNpx1c
8eLTqjwED8E483BAO4lyKwyiV4k1RRigocN7SLcqQ44KKF+nXaeKJ6gxYKfnN3fE
dCNwIUm35X5L+cEUriYNRL8qume2zryjT/gaIWo8D5sJS9p9LOZQoUwvyeHFPC29
bf8vL44kHdpiWifRgde+1yPkMCUYDLehdaYmJew3zTCm0TeHSsin55fnDKpABjWC
s7RAJOeENBNctO486gsTpeAzRC/2p21TLmivOkivhhUL1aeF/pQu9Z5qOKo3TbjA
h3wS/sHbqf71HOgU1bvz51d/5eWlGHif2/rUW/FQBflGSbL8It2KpvsZeDMUjO4i
VYJvXGcKiHkiA8DxnSpu0dZxUscjC8bkDppFoaepwnkVCbEw/dE73Oe6Ia6ucORT
JEqJBFimD+88xMwYeKSdTce7E/rmJPr+jy4oY5j52Uaz53mm9oZ05zH6Ks6bYHfe
zfq25P4fSIZftL0UXWNkyVTS5SCR782IEa40uBtS5l3Dptst9Wf9wJ/oNdQFEJi6
`protect END_PROTECTED
