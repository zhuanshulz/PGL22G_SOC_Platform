`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rTVJOq7fCZsrh2ZGH3/w6Cf2h8CUXKNwz8z0+k4jR14dadvC0JWHNkVNdHc2BcNg
M8QAPtFBm2UztY+Chtx/3zCRqi+wh7tgqc/2ZsT7CCVfCC3WKXr3KkD75Cjw5iYf
qTcxFpmH59m8Jbp3qcdJdTimc51dI7zU5Lc9OM3n3BMyeXju0aXS7GSZyyhiVXA4
MP4G6banu7lbXARX/bmpNfWZnSofTrazVNNMr+3q0qoE0hzvBb6E7G3RRJ9OmaN5
cAjhMTx9lok1nz8ab+fOXYKMxPHt4+17DL1mB++4K0ISc0ySu7i3kutKA2Fm8FLX
dwTdlr9PSsUlt3ULD4O7GQLx18QeUFqfwhQ0Ld1zVoWM5baTK85QjGfHAunGxDbF
`protect END_PROTECTED
