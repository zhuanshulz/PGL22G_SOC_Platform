`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2iCUvXNG3HfREzcEFDufxUDZs3i/txhGYx/7m/Up1LJBtCF147IX3GJfRGoo+YGu
4pLp71e+pJh9aVbPPWd1pU9wRncUFdCjCpn4W8khSpjxEKk7/C+JpT9k8NE84zl7
Ehq60hlHAToWCtTu+g1cfSQ9bEVmBKsAIN7MB74G5j9LNbQ23gjyX1yo2en2CZWZ
N2FPqT9GvMz1MitAu7KfRPid8msc56j+CPAhCkcC5wF6bZNwJqLeV3ZnEo83x7Hj
cEmuHtgxEjWEkoZRXGN8SaC08IyovvthvN6lImLJJVDKN1nGE54+zsg5E/bSVUyO
4GaFjtpm3HayQX4QjXFXsT5vXpuWb+NmDsWDqpgIofYBPZZ62XengZ6f2NFc5EhI
FVXYd3wro4c9j+NrP/IeiUQrD9y1g59PUQ+QfqF9zv1VPnmyHwiN9b+ugMZknbYR
LK88v3OcIM7EUx6mpAzDW+jGmp26U5RE7FLXA+x6T3bL/TjwdJhrt+35Rm3cBAkl
48VkmiM2A1N16zdqGvZT6ry8W6cj6iFl9Pr2qiEQbxuFiTvJanHFzzzbWVQknniQ
ox1iRd8OXXDLZctQK37huP8EUy1hSU6xkoCUc+I1uEUka9z9XanZC5J4FjS3zRyu
tEyLwPKTIsszNbWefdX9kZPP0EiKcE2L/QGXGfYy2G7KTozJV+W/NKow7KflyBCs
fvdMs+eZ5DPKytq/wPvk6WvZxZH9HQg7L3yp2/FPGnpYuC/f4WPO6DFxhbDtqt2i
ZUoCJxvkFKTGVm55LY5uJIzu7KaNir0UWCu/vZDXMX5dOM2BaisH3Ev5X7mmv1eA
fHy4/FEndmPLRHW/MZkMbRuu5q3t0veH+IF8eRrTW9JDIJf5HEl9CFeGlG0A91Wq
`protect END_PROTECTED
