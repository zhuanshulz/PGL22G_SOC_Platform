`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zBQxW2Kxt7p2P+UN/wczNFVwmbv/O5SbMWHZAMlg33ijIsiQT/w1NpcEvXHDtjXY
zMm+Q4yAJKuhPnC/aNdrrDuER5z7gNKC2CVJghgPXZ1L32OSCVjsUCsVGs/JPl5Z
COCOTJIX1Bqc5MAEj6bZZvlJ+6H+tPujDWLjEsWpUyIBr6JcosqAehI3wodgBaoc
uWFVOxRkiY0QszVTk2uaZI8WmMbnK2MssjEwAjpemnytoiQstXdqTvMvjE/e6Y3c
aM9a2CABl1ICsn92Hd1jMv2Yf0cepDaKzLo532EZtvWVhwF+dloPNS/BbJdcgBvr
ieW8jzR0aAd9baR3LkCN40BQIUqu2Qxgkrk8sKPru+j9NYA1I2gMwJAQ183WOUIo
r0qjfB8MNn+ddVGVNz/Jsil4aC2kGRjvoIh76fitzMo=
`protect END_PROTECTED
