`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0rQnueGI8/JZe+1NyjKMFKq2Pw0SH9ps+y+3T7GRDElp75iLArDuQ3WrsdudjjU3
uZYpl2CC7j5XQg4dtyIY5ZFsLrNzVBtrqnP5bUbcd1E591PyzzqRcakto+NXk3n0
lOGeQ5RVgz7b30YR9J7dsUZTyADL/bfYuvTkCSzOst1Kv27lAZYwUMoLhSnsfQaX
qe3HK9KY3aCBwLtzoscsmRJKAzGU6yFUV3jamQ7/3+CsWRPNFUQVhrqPW8VGLXZO
xlnXWcuvaJDIa2wcXxODYHSNvhrbnnNVdXmcxLYA3NUz4Yfl5kg4ypte6Ekh4Ara
4DSNfosImIMcGoljTuH/ic/Hqpio3UBJIXELyQRi0mdv43oTWV6Cv8tLsK4LEUyh
OCEJdtWlie5goxFAl9EYY31ZoFpj1f7Kof/BUFp/6NSdCKAHoSI6Nou8oiOcwh+9
9NoNbsvTxEVLbFuVF8EcZU719BUxoJ9Lg05fVif2B1HvnNgBqYcOPpmXS1vHi7tw
jtDICGBdor95VQ83oTotX1Noc2fZXHdauk8kDlMv0DvsMBKooOxdZlu86/64ct+c
60NtyjTdx0zhMQKu+LwM6N+ci+sFPHDuknWgqlymlbnaDjGHkdDQDyS4oruUYVEA
K7zyQ2G6LcZ+PFjcczZJVW/9XwpEzeCXPSW+EmalQQWD5KFXrNeyZuYPVf6S8i0M
cYSgybB8c+krnhmNqN5cpBTEG7n76KbNzyiW2YdGj8tbUndtjpP2xy6/HNCp8Mbc
TMjxuyfNhBf118geY9ZqXGeRTBay64kRONFzl0Qlwku0bKf6eOxaKfCBngUI9XzH
4or8uvG7Tx99Wp3xG59yTD9rLIk2+SiYWpKEfMTImbdoC+ZlGqMOw0VplxdexdHs
nnx4LQL94pe6nME6baY8iaYWeIVYwP/GuYe0QQQJAOzCb+Ud8VyVakk78CeGYfcN
1TvcK5tOMXCGKzJNw3zvhwF3uHkvi2hY/3+73OBEdkyZgv0anrw5GfgkTOKKOnNr
ErmYLUWWgHyGs7vMvp+cFZVR40szxzwP5fsjHYLlH/1TUrKk5Fz6SzQLJNIdcIc9
N5Rb2px2lLgHR+PYxMAcLdWbjnCQqJ9vG3ylq5r0wnKFvORVkn6s73lw7hG2gipO
80UH/rEc+RjcXZARZhIwcWR5upbJ/BAWGBA7BWEWUmmsFCBOaDsvDuP5msoLTAg7
xsJa3V+9j8LQuUWixeFwehcKHbXkQEh/RzN2a2DiWNw1fMBa/Mmz370DiYAuiKds
Og/Y54Zd89FWV8I2oxSBFmw8uZHKS/m3CUgL4N+U7eUam0BsWZ5b/XyK1KYw6Xks
SlWnqdgGcR5SftftB1HsjdTp3nJI6Dj/p4L98IOevPAUeRGeMRT4hpHWUyaP7vql
tV2qpDYm0eK860e9ml6q1J8hmF8XPsgnxkGD0P+bVccmtU6MTYEOC2bbutTXrEui
0GWy3KVt9DaC1E0I9WCi4mEiS0kxtoRUeOwuD90gOQTjkktEMhS9p5trysn9GbSC
D8+PFKhH5pGVjUOe2SFuOZaxdYMhqecjZutTEHVMkYAjqlCHex+EEDnqE5sSHy1H
Ahx4dSuLiavknxRHKoZav/EEZb0WSUqBpaOiW8MzM31+3/2e1wDxWOiIMniq1567
O56+Rnd65JofMlK+2Q9kCGtinbZI1ARGJqoKqzL86ojg3h/948UIcpVbZurDFpGY
uwrbrlT5QYI6ac/o1k9BhHXEgmltJR7wmPQyosuJQYxpWAUJ73HtzvT+NMZvHWCx
J8PNli4gm3VheXc/U3fdr/dKUs55eYi41PUPg0/bPEwAJDbOgfTYyxp6so9tuU4f
Pm/i1/qgzeVMUcuYrQPfssU7K6kMAd+/oUj9wkh5oIkrudkDsjICaG3x9NgtaMty
beGBygs56J5l+bwZygSOV1e6WWM2O5jf03ZxULfYQOxoUZtKpX8Cb8a4TBryZAuZ
gJGZ55416DP11VOeG/EJjjywsDnSHOaYOxMYnMX2b49AIIg8nu6106uT9yG5Hxwm
exj1HjqaQzUfKkqamarW11nev9y+pMpdNQa2i2tyDzeFyG4rJ7V77CHbLfz/btNR
/rPS9N12wuxM9VWvqfWUZuX4sHS7bZ+a0HRUWX2xENrQT33KWPTZ9wxGrlIAg8rQ
zpPK9jKRaj/zGKCPS2KJKTaKuOHwwNNMMFijMsEybIAitmrGUlYARcmXMrlfkDTv
0fjcEV4OxLeJZcoMryK4Cf3Afxrld4Iry3+mrorJ4+W4kp32LVpsdATBN/q+RpsA
r1/aoGxT//KSKA6QXTlhLLXk92EwHiJa9JHdMlvRdw5XXBbhX6f26lhX6gRo0IUF
PacJ+cU9Krhrnahmv6yxukKEXbqabfH3SCYu4Yl8+LoMkJA6oqKzErNpQeZ3Lonx
V8Fxc0uHcM6ttk6RnpqDBb+c9bxxWu2Divh+C8RZJdyd08qNwd4UvkoJlGndNBKT
WKZvSU2BNlcV3mXpsIe5KiA1YErFrmBK/p1sdKyZEe+WdZkp+fTlYUfpx3Dz66eb
Pd32QlQ767C2RWWkEqO90qSABYNAyo/+rg7iwr5bP73gAw4jyShbZEeueuq6mX+g
V8VVSNveZnZNHDC9MYqZIp6mrYTeZfaACk+bE/ejaNXBRmiuR4apueqx1On2ZXqr
4DYoCHYBgNh8Z8Aunrjn8SpzONK76ynrbyDFEk6IXTP24zrRq8LEgSpc5eREKeNW
Dovtio5AcPx9YQ7COXab9onmHu1oyIAktMq6yYICo4DGBRC/L2ZFSsM/Fpaz0GUM
SIOMrP7rvYlc/TOD7FI9zRMAqduaKfxMNjGxw9/Ze0Bvvprdf3rHXLa4UIb0zlhV
6M4XvwQwfcqEb+kls5fhnKvayBfcCRE5f5yAbCyJ7abG/xDYMvkVDndz/QPzwgTm
n1UCkwd0UyKar3f5QNtslSIkRBK7ZVoNc9QcmFQtM2C3SDlftJhrpEMZHHXEyY4x
dSeCQPJG+PmyE0erkq3X9x5dTPVlyf5sW1H0VD6zaB9x7GgGZIfUGEjQfj8yu0P0
C1I4SQVAt7OV7rSuzGKs5wohsXn1NeGzWgbJSldCSUw7cxRPh8ezz+xaJ1jKiu2p
trRiYSSwW0CtXr8uudjYxBkwZWeBmGm8BAnZzi5l/+fPrdfTzXQmSh5sEzNAmojD
SDWja/lqMMpRsaUWmiW97ipGLEvpzUTdOWvfDtaj6xjnB2UH/S9bRjFqSf+BzPwR
9HJAf8edY2N0mT9dryEz+dw1o3CujxreY/DPJnzGkzW02KqfybzcT+F5vocq4AIt
m2zRGpJrVoSc+CBnN+LUGpv9VuK4KWyP5kXpoQjczkmMMUeu/Lrw8XFZZlpxk/Q0
cQBty0uETyaWdXPTiZIX0MFdvddT6/53wTkUWQju4VIOFXay43aarQNsq4l1eU8i
ZbrujxIygfZCsamKs+Q2I+Pnb4WGmShlFIcieuZ3ufOPVMQB1YN3Q6DmhoZ1Ztdc
GeKGDoYjSedtpeqZXuFQNALpiWz486LbNt4gxWm9yzTgM+UAcNdv2CYjVOwNfSWf
VPVuGo2geGEccrazd9iGmdCD2hV2PNhgesN/nVY33AEEZqweTVOa5XpDBLr/XjUZ
hVobILyb6VLZyge1+lNiwr7GxYePzCKaB/tbpqh3MqIXBWa6lxK0exngAxV5bfSA
VTPwYDRnogBLLutxNxIPDEcP4YfJycFjkinyJZlGjjhz3RC2mmcLQI+bjuQL8aeX
bYDG2z4pvsIg4lVS2oBSur2YCoWxhS8EvRnQfFsKTx12YfDOs4Lt3EcEcjdCc1CC
u26UA/mrJ2Hp6V/UA1KIueS0vpppdZqmP/qAh7vTo70v51EpgKd+WbxvnwUxOZIk
oRjBRBNKcvnW2Q7aMIhGI/+5mEDRFUM8O6HGT6o7YJgBI/bHfV2rrYicqU8760or
yBVu8h5eCPcObXeENodQwNaP/vroDLlpPqMJgJ47i0xx7q2dyGtfRwQRr8bofpdm
V8UXZQEF5pUUiuHENlKqFSavsp3g0iKkNqM9Rwanti0cEfFukmwf7d1gJMI/zfaB
ZdrYTH9v+tnEZylLh2nuioVcAEdZK3M3JfrzbEJRGZGUizJTvUXSN8S0StkkAzgu
hGOH3+CFvkkMgM68qbJD699BPoKNXNUwb2NxpPzaHwQHCVegAXOcxQGOTMKe8M2I
BTUa01CWr0Ln5tgxM7sx1htGnjxw6K8hAMupVDvsTalQXL5tu8H/TCJrf3kVn4lp
Q7R4g7vKCQfoRo8wdJmGWqO6bCUkmS81BlVU34BvKhbtcG6gqE6txl6zoQgjaqhr
kEknHCxx7hMSTmxA5xlKNUkP6gCqixvRFFnyd3raESaarNfZCfmJmtAFD9VkN41J
6tv5RExuTA+vCa2eBNTleJATI6cp17RD89ksk9RRssPUhXMPrWmk0aLiZEuyM47X
hQB8IqkSyEOWsjuZORW27WTZsByBkBBRjBDJW3dvJvMmWc0CQU9cIbYdVj1GBbEr
qXr3TCI1lneshe41Y4TtPw==
`protect END_PROTECTED
