`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fjod1E//f1Fiv6HpwV40BcdSc1cXRtHHZPwqfhvJ00a1OXY9Vm3aNc/z7ogqbI65
MN0YyA4+Uz5afMVxxYuQDSMJlBU5r1Sp1+GSxI6mu+aBwdz0KRz5QUhgq/kPOLK1
WeqFOlh/2+jSAEwltzI9ZfAzfLixNvu0ugMwg3VrgnvQ6h3ijlruN5Gaf3Uijbrq
ellIhi6NoVcsBOAelFuLzUTiJZV0SpBOlm/7eVgBzXN7oaZXwVi/Ly+UTIm3MojN
KgRDELuD66cZNybEcIuANnOmJWT5MRHrPZ74DX6Gq8VxVsPatcXMXWM3x8bHIDy9
DhqptkHm7JPJjO7AYyZY9gptIFqlBXWXawrF5CZh4o0Xp4b/xk50/wGDw/t3Qv14
kmEQLWgRPewWanczzYURdZcZNMDTHkybr89X6+3ZmuIgbPARWiCRRctwrVNg1FLA
W0Uei3nrDcrlGGM3Hf3+pHVYQ+5hvOP2KushkkDz/jaedvsTaPsQ90aAW+js58CD
rbkwdM/lN6OkGqKCTZ82au1psZWuiAdRvlACDOduE19hWK61f5H+PNpJs7mMoPCq
EzGLGobWCrn6qdGUEUTK8ueJYaCYgeKbnt9eEG8HpNKh/NtluAzIRFMMJ5lybbJI
cx6wwpvYr5x8J3eRIPJd5nTFZLNxzjj1WOpJdC4V6pQ=
`protect END_PROTECTED
