`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BHQacKt2tojv5EpTSE83UEZ8R1q5rg4Qjz5/HRYKtKArKjmCSTmdXhm8ZWX1PZDr
6ROn+mCA5JAsEUtHrF6BGju+8Rg4rYuG5YZBk7JLHaZ7AKMhpfJ/NyRVClDmGsqI
jYJsw9vqHfeLNpCRqcg2gh7fT1SnbO1j2crnUyMyIAGnpgVqMYDwrDQwKnChngnP
Rd9jBW6U6HDkavAimnVG2ORFnp0pT4q1LBeIFdZmPbJqfkpPfav0LCSsphWVMAdl
m5oTqY3gilUxbT/wRu3YTND6SOBS9hb5cLE4CC2XUhRxQxgg9ei/Jms4UamKaS99
I1C9gqBJfmhdCImkXnuJmTcU/0kP3zggplPk9TqkMsurMJZmDRKAFQ+E71ZSr44Y
QLNsXzV9kqoOsCxT7PLy4Yu9dbzArs/9K7gS7DNt/A/U2zh0NutkLVGyKVuEP1nZ
Y40biEY7bQDLTpu2J8CtJt1KPxWiQ7soHdvkWBAqm5FoAXin6m5kYBZNqueeC1Ow
suolrwEMNCrNmqHZKZ++gVbhXQR6bKN3OBoh/XiN7eSZ+Twrr1CR9P5GuE3jY9qm
soO2yzDnIdh3Kmya9P5OHbnjESr8fVDzBPFoeZpV7lnRz9JCSdkTU0lLLyH3Eiin
5v/+n/5WZVMW8k3UAzSRBLI5FfEEN1X7hxNcu1X1Rs4DliPIthD/5/4VIxGVndG9
2mwZ0Dsr0P8eOXi+7snsSh/p0HdRhlf39+F1DSAG+k6YE2oOJ0dAIf/RBMqOPnPo
mCSrAuXgXul9Kb0D+PDQZILwhTpPJpZ4IuDthEHTyU1g4W9zfEbP/uqouQLevwfG
9GNKMK1zGPBVYhqpg5IHh7g5VOj1HAZrtuQkEDlv5Wow5WG0HQLigkwn5kUKFn5h
dj5w0bXCh1jocy8fRGibj1wpcekebpjhVOnlEDjAhH6kXai2eu51P/KzELO5wOAo
Bwsm8FRQ0pKwHfdfndL7/Dgf7+6JMpAnBC3m3eh0VnxjuoJ1mMvHcqkRQotXiCQF
GeIz/qOfBj+we2ZyuP5FsX6YW4wETZAYJIrmixSf5oIoKokTTlnX3bGwds0elJSW
wpc3jNMBZcAb36HxWVAgvjXeN0oVbg/+8UiWy606MepH6K+ReY1of81gptmEFGM6
4j+V12G1kPnEwUMe+Cw39F2SFRBr34GhmbG0IVRfRBYd7CJj4Z0+IwWTsmARj7AX
UVMxjRbhgm5dDoNLSo6NSsvPaNwoPVF2DNJIsQrCkTPumcv7r1InK7VzhOKEglCV
HFpR1jqpU7Wmgskiv5DJnZGZDAizODPoRJN5k6wDxOLG3CgwVqPeji2Xa82lS4sD
cFqI4Ij94KW7sa74I7XAd9XFrrTguQFqX7WZJ+vYokJeb1yc9ySuoGCC6vms6pgi
45MnRsRnPAJ3fDrJrC4tHcw5SZCMhfwROECmvNf7MIgOqZPzRLVHcE0ZXziTKpKk
SZGRpFBR2WlrlqnbEQxg8dO7A93x36jaJlFnnoPPgoLgXe+0IVIOacRuSxhichHZ
heCAnC1T1Tup72s+r3G2yopcTylYGfX5TSr9qtUHmZ+HxKg1mcl+dAm0w451kmPZ
D1gFD1nxi7UcF2qXg/PreOqAoeu83+/GEhAuPEWZLgKdgX9IX5lDPIeUGE1YplAK
k6AWxE4mTsvVgdPJqcVTUek30R+npTINSeIu+PmhGkwwOOE/02ES12x56mEYc9rc
Fej0uFyIW4DZFeqmvjgpo2/4qDalnttaw8a6IlygYvlYBCET2A0eb0msbwdwmP4b
Q3v3fclZ0GQ8iDyxrSkMtjIpOJi/5K09xI8DQ7y8gKYtAU/UxtcUuxSLqpGAjesx
TBywpB2uvMCGJ7EqT0TL+llhrxbdxufOOYYGDex1zO3+6fu02ZTo+4d2Unb/6sEW
97MqhbWvTqTrN6yfhPUuh714i10NGQgXY5lZomFULkt6tD8SJcVJS7Xq2BKsAY0X
9fDIjJsqiXB9mwQiRsxrGW3ykGIrgP8h43UBpyaphkrnUQFYJzEyLkI9A504Ze21
RDyZUsaJI3FdaiJp5xHxa5h3up0xdjW4euuZ4UgMxhV/zQiYYmcpnwacB1XSzhgN
op2+YLq8Ou8CxXdVUGUW607p+K/8Xx/MITKtBeBpqfuWwRKibPtgX+G9NrY87KR+
jIatvjJIN3w6QB6hkuE7ou4T7E7kGwOkWl6QyKlLK9FyHxrsdEbyzQNv4PkZ6bUb
kvrH1MuScPbsiW85l6XQYXrXfJJTmEJNHPaRM2rDjh4UISRTSU97MG5M6UF6Vd6I
ONTL4zqU77LvfPb1xQWDR8SFSGc+V4ECglxkgJyrFn9hFbq7mziYFmXJQcW3QMJ5
shAGLNSQZAFkOZh4scKd4zpZ/jht9ml/8SmM/RbCIpx8w4FJqEI9OjSdxbT7Unx5
sCt8tQTsbJNAC8z+dRCOuHtMzL7oF5H+W3KHe9aUpjpihlZ6YpKZq3tcYmG7rBxa
I9kKmDTRpDTN57EW5KZNoWH0vq5lbomEbdzLeE/Ldjgzi6Mk+zBJ0QrOrvWUq7es
3Muuk39ZvWo2jeyJyWFOMdKV6IIC7IsXBXO//QR3UhGHvJCHEs7BlkA6D4adTWjb
LlL8Hswm+7sV+V+SEQKuuXU5bZ8sfXLWFT48798wqAOSZwiRxmYVFg4tEugQ/IJ1
3jdbb7r1hEPkDgkKxDJtLt/QsZYJwonh4WfHpxLOzTntclS6QqB+DODT65ALI2TA
MaUf7retkFCxSHdPomNa90hJbb9vijFgzBPIUL2os+rR9s9dQX9W2IrS8Y41YtyD
q7FPY6GJWi3dakH7Gxzu7XCxGHE8vZuR/IzGMc7kjPyIRUjLGK9VSdaYAZd9ScDN
CdxFhc92MaVbDeTR5uYUQhvE6zhAAkkv44G33ikg1xXIgrxgdSA7Zf9al46jUA9J
Lk2y7sE5sZzvz5r6mnWRJj741nuJBQqc7xw5yHATo/cUDBi+nlOuXD7LQzrRFA/r
oSwR/VIFUHyxm6JcdwTWp6CkYvfhgqwT3tle66CZqNbmayKKDQ/bmA2c4uTxin8T
Bup6NM+8Y2U9KfEzGp+Q2HeGX/slyhQ4EsC3llbpjqQxBGjRHGzX4n7INm5fkdvE
BeGuENGGlpLCvCv4q+msWcI7N/dy9kUaN23ZhXvaMbLpGRT68TNBbL8/d6x9gOT8
d0QE6mFJeEWka649m01T+Cyna6nKUdCGflol/d2dYsOH5d6VE2HMmC/ZHQXqtS+M
ehwo3VHEb4l3c8R+p/96BA7gpQlmOf2/tHaTxN/4wEv514d+5ZylTp9GV60qPJZ9
FfU8jsXbBC+L+z+XK2k0Ykk1v9CMGaoLjVy4O0lkdqK8JYJm2dwBi3gLJrC++7rt
V0S65It33K26qp+b9xMpyQuwfF94aDooJgSXYscNEazbL/mpsRQ24q+eswUCJhxo
KmL4ABXjbNhEZaoHzWrKbeufjDMmPu+NnsAFoHd4U5I2di3q2Nq4vJGyaC2yc0rQ
IELcyMQHWk+OAWYjtyeIdapAT//rbsXclpnDb6WI8yMZI6OUpckxj7fe3ikDXdn5
ytxZnqTPKgaOuhJ1KBHYWxdgGqLCBIsTjygypSFwQaKzvroZzfiyEbb5wPR/TMX+
u+V1tultTVX9bhc7asBtHRKapxoMc0Q9NjEFvfKVc3GU3OHFbBWDcc0pw8KDx85D
acNKZYtWajTLCr0eT5XzKREUx1O+pWV8hFnQPLGdpxr2yX8tfSlMbEGQ1Qtd5yiV
dVjyLYCFjteULcl/huxQA5fV4gLHpdeYmsF2Q6KrJYoLZxLIQtxpFg3ATKlyRg7O
6wWPwedMbtZzjhd2QcgFFduYY2tfmNxOrK6HfEgVMxR57F8yHp7K4I9ylpDn7Mig
KVZ+2h2QNDH5skkSt4bizElbPY3SSelgszG456ZboprOfa6nLrHA5spMJYFnSgve
jkx/EnNQNAo4GchHHEiONvZgC35M3aNoSgk9Dw0GPcJ3HZioi3ijd5XfFKWCcqpy
2iqQVkLxRHp85Bo3MXxr4xJlu6Uli6XuwwyTY8ip4WDsbz+3QDjh2oULOYoKumLZ
U6y+ltvbg5YnGnsDgrNq7gL8KE5mRw7lKbRR4q5mUvs1PhsGYsN5U5lYjv1I1vvI
SL0X3KMEztoegBWRR3ccsARMBeDRqGf/O2nc7crxtjHV7ovnL6P1zDvBDqoXUTQn
JMfpk6ieDOEEsyT1GAJbFzaNwfG5WkQYKR+MiooI/hy4iKB3n48khpPNro90jpBC
tyJx2S+08pmLwOlu8iem5WVQy26sRPWzuRpeDud+9HPFeRvHEKoL80IkWxJ+hwTa
rTD9WsdjKQi7KbdDH6Y+w3x2Ul+d476IINtPBQAW1SmaVewrzf6OcGgFKqnSod8k
4USD4ciL1dx/z+pm60eZ5/2xDyxlEhC9TKZDT4OYfKN2TygkWmXb0auqkdP8i5s3
t3Z6VbP8jBBPieBK+6cYsKOHRvH7zO8kf6fH/F8Ad9XoqR9u0qLzHgS+Sdvd8Rww
3CgEhCuau+KrR8bBW8jhVGpJMJE7bVZ79BxiEi2iiyn/SmsynLiFFPUbKiasFbiv
fs9tD3zObdGYxAyNq20sm+5TL02CKRoibSVCn484tDlTPNXNZ3eeI00gEUcll/qA
19MDvlTeP3c9AOVsVyWkuQA7GB69B1rkitJu/VmCiJv9bzGRd2xCzDnMI8juDr4K
t6yKwQPrzTM4xqf4m8/V2ngSKoNwI/si83TTX2Y2SKc0x7K/KEiif2QgpyipWq8b
5TeZQfJqY/2sCgLUMZ1s6EAklvm7EZa322zcPC01SeQyGCkriyLHBKXmwqySfA/h
Yr5MFXbb2TWqwk7Cvv8YKZE0SIenpuP8Zq7ixom7ylo5o6u2jBRGj87kUTRhg7oJ
re4xWq1vpVl3ryzvDboxkAcZhZ3miRoT+KMNszxwEfh/1b1Q0dWAkI9bAly3ovD3
jTDFEC5QpKTRTEMfjwofY9J+nCUpJG0iJlJ24Ha3d2V8piwkN1wDENasVbvhYxWt
Y0TYGNQML79jTmahkWllZzcQ+g4SEJEWImpq9eewUy0Odz9TvzqJFKI+JL9Qxjn8
KM0MLA//FfqZINpYXxE1LY8++FFFCVqHoqc1nK5du5rRLuTRKGpEHkeXdsbAtwc+
oiGiavbjmRtCdOiR/To68BJCGXmvT8GyOoBEQQay6cpNi4R3I7SPAhHogg1Vj1NV
2Em/uY6DlcN0V+kgoci7rlXNlu2iLwvhbWi3+w4bL3jdc2xIyEBf48oq0TWBhVno
vgi35EtkPnaW/lqv2oSInvWtECS4DTppZST0JFuuhz3BCKb7wgGsS6uBMZevSnfF
xK8B1xsDbswMNGj4t5jEXdMDVJAcgcNjsabr89W5ES/KvvYPIR/cB4gotZNrM8QZ
pFd/CJYOnh036qtzXs4ldWAjJkTju0n2Qs3t24gM8lYdSmsB6W2oh0HncIT+UVbZ
UF+6N0pie8kaIoNecLmEvXGInVLoTqZtt1mAH0o9/6ajntzAdwL7Al1kr5ZUt0VS
ssWo1YQAfTqp9eWMkuYFBDH6jGFFOIQil8P3HTH55RlN62NU6MlSplYuSAKDAtPr
lOkUAI3wXnmw7s+I0DOxeRPb5tcfqorHjVNzsepKgoZqXE5u9ceiFn1Fbpt256w5
BOgJ8M450mxQYRE+tRl4W92YNJInkaZustRUHp2FM0kTDGCOSpWBMIqJEEUpsaKQ
8uPsww2tG+mGVoUtlfkVFGvYHvFUNfDzL0NZD5D1l+VvW5DU3dnRIhY0lhFqypov
xbG2db70qxMz6FvOmBOQMgFaHVr0qT2cGcIuQ63cuoAp3EWcKFIZ6AJIW9SEtj66
2FvOMv0peec87GGFR0PXgUkyFAmRcLqVDNSVgT5/432y7mfgQjblqMgGQFQdGA1t
trQcgQZpCsG47FPUzYorC443POt0QzuXXBe3g5E5F3vvpOy5cO9zS7l4t19pY87k
2xiho9YaHMQ7vrV83v4WokLzsjUon9Re4qwRjt29s3xnnYRrMg04dHXeVYK4+HQ/
2OyKktQyOwNTxIxqK+UKvfmA0doOvlzE8HP1AJIgXZU=
`protect END_PROTECTED
