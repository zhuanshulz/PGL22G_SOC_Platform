`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sj5pu3B3LBrsUkuuY9rSm9MxyiWFWsZrufWP4v1KeR8XQ4a6FG7zV6YKDgoDmFsm
x7Nqj7vOTJ7+Ayuymqz0pS0aM9EJ8lYUEN6L8hXuVmpHWNW8eTzps4/IfU0tiIcM
7iJi3oVeF+ped/ihEL6ADZXTrH/B/3S/T/jCPLBOUn34w3TNjuKXavAXCQKSeloE
EO3umlIcRZazN66zPuZnI6xX77SCdA5WtFr1u7s+urBOZTTD0Wuh1bKe9w4xrkFK
g6gTg8CoYHKmb9PDalk4xw1Igilx5uAcPusYSNLs9tZjpZNe1lG6EsnleBbOL6mr
g/AQuQdjI4aS8+7c55uysxzf0C+2vosoA207pGfGQBBT1fq/XN3JR9SuQSYJHPmM
nT0G6fqRFUkNvTEgRREhMP0fUh7PD13rl462cSbSG2TIW6LxgGKmMohn4xpVP7Eu
q66KJpdcSEOxUUXLDzPMLY3rrXYO6cCxMmki7zT7FqvsqgWqFJ2+1mkR0xKP2pc2
NolF+WHZhOCvtAwWGxaep9+s4IExqH6dI9Nq6+4w9+uY8ghooRDc9b511rl8gv99
mms1rumfR5gGTEXSBHlFOkSBR3wPHTcSUQbaNmq0iy/QGPLjAFBrcK+OiUInBZT5
E2nGAm6t1m0pIHiqufK7YHaYW7IaIHufBkjGCK1IUqUv7GJaHv19/367B4m+iR1/
t4tKlwKkWCW+e8NRdVO4195zMBR3/M16u5rCys2vtPkqRDj2lAWLe5Zm/yA+wVDu
rHWPJVW+uOshi4V6NvRXRtMq0KxyEf5ZGYCvLrcHANHJyCq7esYBTfmCClW1DA1o
BjVtoDFY8hcmNG3rYFgZIT3xDc9Y4ktTmkT8Vgosvabfxn2zAJpBEUfKfw5SgCMq
nrFrUu1qf3AgTQP1at4YPFNcB7faECBkhKcVGUNahtqD5lfwcqMgdjrs4eA0gFe7
UKJttG9boCFPGGWc9TuNEi+v5rQcdH+swgVzGPMtQQpmTN8Kjl7x3DGCMc3GJ06i
csI1HGoOn/pKq7fSKW70uKng56hav4cVxk0yNeYhOSBOPzJt1CrWkLcyeZHhi+fO
xn9BeCNuB8GScA4Lxh1wNb4XcMwkjaGVDOPEvn6y6IVV2vf3AFEPapCJdlPCY8WV
wZ/eT3yzW6xrES0g9RL+SZPw/CAf6On7+6a/YjxVHbNzQG7f8q0ZR8NhFGyzffBk
8+ENuZkYo1H7/DqOy1X4ZaQ5rDiM0qtyr5WFYtuGew8F1P2/NsYRj/UwN+1yKwHd
hOsb+WcHRSeBvcE0vzhHUCqxSkTn3OvIqvYD8RLdWpjd7sJeM/w/vt+xvu0SJ8wk
o+a7Nrw4lK0QeuEyzUI+c00/0FJBiuQcV/mEgTn6zDBVVkhqkwZWW59FtXWKfWDH
aT7dhTu7j1P5L+Q79qJcbSlHQtXWp1zVgo5afHFG33/Fz5AKJGdsnuEHzfeJRSBi
smrexO0rqgsn62axcmygE6KiQHa7QUsjkDZtd37O+2vPKBcaFvPUzEjhWJOJvZqd
/+yFyBT+HzqpiQGxz72EAEwoBG4EFP6fp01lig9Fk33v39ItYawIKBciH+dTb2FJ
nLK2d7NgGUevRoit6EFLf7vwmEyc4QNnzSQAQWygMbGaQv+wfMLlKFJo12banwET
QiwskQdFGWd2ax6PSyYmYfci+ubGfQba/T7kY2EhmVs0IyGBovrjSKkqozsEAxm2
n6lXGX/ClVMWXNMrOA9OMs2I7PRuuxD6oHTgzoQw8maCdFZS345ZAc0ck/tMXAQp
8WTe65uEHtXPZDs+bwjLWSCN+KVPHkXeoo0UHb0D17JKGtGMOIq0nHu1H2pW9lXs
7POrss/j+uAr2pYVTVbodQ3p0NAMYCcd4z+JAMeQ894uIlEUvlWLVvvWLEGBQwBD
mpDX4SU0LwF1TPG0e71n6LNKaxcHNlc/NyqzZbo497g7IEA8SEuOfO0OLTEPb7rC
5qI/fRIq+7puhTKPM+BUZbN/fRZ5v+5jddq1T1un2pKD2+VQcUsC5XLUlWtu3djo
ljG7ZK0e3noMSBBVZM1kCkqpNFQ7RjMnd8xOSkzkksuEc1Sq+N7CBG/zCCHZkkul
YqKqC5GdF46UnEbPQavXZnt4tMPxw5o6alGPIX2YBL4PAQ9bb0D7QRfdShNxnf2K
bJ3044c65eVLQ0KAnAVMZE/7fUwYp2Jady75/52geey46vMTjjaRAcGdeylWLFEN
2XXqBbG3Kghq/hKRkcJsYPJ/yp64rrQO4KAlqDRw3tDi+Hax/LFdM2N78hsM7w3r
mNxnBfRFwsAgoZF6jk6+8s9PRiDxy75PSXtUnUSM+uHo/R+cojF8zehbkV7nC+iD
c4lB/mmnaGx9gZDY1g/SaGQqV6ELSdCCv4B17z0m2W5W7beR0uTVhv5wCi90njQQ
RoN5pwwcfW0Lg2S0r6Z9MqoCBfhSIe586rAus+MBuNVzRO1rVB9y3GrCj7cFnDht
jpD3iJgHHvpw/bSljHE7YcK1SwLwZZY7BzGAcekeXlxx1A4c+Hqlxe16gKoUaTgQ
Eso7SdlOjJYUcAaSsSniYTuVC08IE70ih7fzhTZcNyXfdP+Qof6tsXdeKPatvLhX
ThoBnBoJeDT4hWZg7HM6bqiefmbrRAxO3nzJJ7pLkNyj9IyhuNk2cdzy6WHrvtc2
kLRCGF3EtgNg+2cfbLN8A3OFqAhyPpQqzh7OB7akZiEZDagA3glc4g3qwLRFiJDu
3mnGRsmMAb6rOxjx3KANj5PJJdNGqnaU86i0Ag/gvVWjTasD9vFjGa36J+tvcrCo
083Nj9H+5sMq1TObQgp9g0ixpiSXq1Iswi6XVqDWboxy6HXO9oGS0k33iT2vUwOS
VWcSfeuwCxRrH06re9O27yA+bGyV8R6l1CL1yrqSu8ZsY/NNnAzRGwjk2GCRLA/u
Zd/hquaDLotx0RnpwQWClsCmAkUudYbydTcKlpnr+ipUb1pKfmqSf1o2/vT08KmS
Y7s7hIiwQ5ZXnHOrAghxqnGlBJUjmF1isv0h9JtA8uJzZqBf5ZCt8zndCtTHi04I
AyjEN9JiD2w7GDoqiO3K/T8Ge9VgiQV1VwxJd71j5ORZdBjT5XAP2Sgrg8+He0Qv
UgRecPu++grOzOEoT9hpjG0G4Myec0INspqfaGkrFz9L+YRDYvDBUIkjx37/xh6h
nf+XfD+b2aQU+YJQlevu21/0G8gs65gfdRvkYWUdTDXvzgm5tkdELfAPI30RXtTS
DU6tU/J6CoArObjhaP4bphj5F9xUrHYTNtRZnF4h/YOyxKzRnYrtUqclRP9Bm/xh
gfVM+dRkoRCV9CVFvmEYHp1/IrbFjSqRb7CRnqN8X70T78agh3mtuPtJ6ouCg5QO
7Y9Oztyv4tXK9P+C5wRIFUC92jinsx0WM7tXrqjKBBMTJu4iyWdJXtyakPtdvxhl
nMfYpsoi54cHy+aqT0tRDcyYgyTKOBqSDOPVbIR48JwXLL3Kp+2Ul9OBTMT4K0aG
WJPSeKpnozO1VlGe8omqje9wt0ctoq2lUvUy50gpvUJorr0AQKiAtzwE3TjQMJ6b
pDNSgQluPV42HHy05gHH0O3rlwBu/u9Cpw4uG3ShiCpJwmY0sfycBM5BMyGVvNp7
cuK/m0lABJ60jRik2RadXvy01HcDLokLTC0TL+Ag5yq6rRUU9EHYlwQfpSNcORMq
9pF3qOLmT3jzkGw0/tqgdnLz86XRHEbKziUe+cux2RHZptyGHeqFFzELVB46N6O+
uceFjcM7wejbxUunSY20u1zngDE/fHNTn6My2qMAGSBUDL4Ae2wyH4fGx/rVV2Qz
4CcH2e9exs/21xlrdamu+k6Wsln5FmpCJt6YbugJC0Dq1AWGiyWvV400wNeFGwS/
fCiLvWglhNNeEoAHUcHJPlCuptj1p+WC6NsxtxDQBMDtzmtDasD5ltLFpM3MD9z6
+VHrhAnMmdYmrUJZXW+WkOAmBl/MHsdBjUcbm9O7KNKNFb86wpJIBOAlNZ1nA+9J
`protect END_PROTECTED
