`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u/Ci537RSgoZDxYlmMfJWWPwOFdPZxH/g3cS2WCRUTHiSzuDR6mxhSo55RIlw/VB
JRlp+Q494n+BVbsIkEXTnvKIyAbn8vaR/Jt5v+Cn5IaN3/oHre0tnLSljXOGeYYr
EeX+7MZJClJI0zuEJ+c7iRnAanMYTcANU34wIbFFV8Udy8cAlF0Mn0BLA7YXpYbs
LnGw69D9TMlbnQ8waPEnQGQdCxR/BeQFesO/c/XGieuEjkLYULPFB0Wgr1Tln/A0
m4PBbu/GB01JlM2AtfmbxAeLuxv23+7RrnvYM2lYmG1E6HpB2VpXIIvohOFQPGQ8
/0XKq6zrh7LnxM1y4tY3ni2+4p9qy3jaXX2dFHrZwoqByh3TgimTP4bnEqR6+/2+
9qIn5Zk5EhRx9Hji0I0IVUWzc2MXD5OPVUApceZvzxnBTctIuJGqVmeyPhzb7zov
3leUj/o7qTN/q8I52ry1wQ8ImE5mq19RMk2Yp/dTmHOygZ1aFlNAXVIePvbkod9J
artTXAH7GtfQ7+NGa0CIkA==
`protect END_PROTECTED
