`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q3QqlbU1zDgjwScjouqOM8Ppn2oOtCEBZqxZXQrWI+rSgATNwRyzQ6meDuUjXl62
piM0LVcFluKkPrLGZQ0ETuKJe9yqqNwy8KwpW71P4P/W17GXaTyrraVFM5gwnkwd
kT23UXlccLPoQ9/ND/HIjK/m7P+hrnkDH5oqEnieykwii8KvJ1ZhSCjoMLULxCUs
KgtN5TtneJdo9wZMd9V3oF8g22K1kBaw7X1+hF90Ev7RdSBeA+fWi8Hu9wlY+mb3
RncQZQspTel1EBTRZpsJPS6yzE6k15YMVVyFjEyK3FXfw6UMkW8OeYeyoIGYgl+v
5Db1njlxA42mClKQR9xeWbi0Msr2PQA+wBx+bxt916hU1JcEJSbgDwBc+EW7dQ81
jthU3RKPdzq6TCz2aXgS3hHsCwZmuVVvrOzcYDRLq2+z+OPhqSgyK7J8h1oO3b8j
`protect END_PROTECTED
