`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
copfD2tNj240TbkzaPTseW+xRtx0wJp3Q9GT0j6Zuq12Ru2i2051CyPb51sXRrae
HkgVn5vzi3ef33gitq/lMZyC9qlFZPLTmQwijOngzcDUrEJ0991lESb9amcHnxP7
21EHRLR0w6oZKkWik3mQ1HSeOnJrq4ZRgEX+3iBuIYJeLa5Zyk0egVHyWTqgdqAf
pJDaccCpsiUH4YUV9LwR+BvDiXXX40W7IRmnfeZYCflAt11HZH5j7acBAf7eDv2r
VoSf07X6sv6wdqfU0Jvf4R6dzNQhJow8a30/uXJoJ6ym1Piq9UV6kvkMIsKeH6sO
kmmKSY2FKfw7CG+KPE9t/CBBInmpzpBNrLS8v/TQDTY+6qDdnDxFi7kyiTZ+N0cl
CyfDoENrluzBQODubpIvjoBs66lpu1W6/N8MIq3sSqe1de3bXEGJxyJYtghcUOMI
Niu4dn8kmCVtZwMcuI/6mI8kNNkwzBCKGu8mgPGGVY1ZZDwNr9Sw2NU3wwYdEz9B
Df/nTxNpy8/DEUgsxWjFS5ZsWU6IMg9+yZ7NI5HfJq6FN73GdN+ghRsOWJl+CLOT
BppmJtIs8o3Sa3Q15PYIqPT46ek8BkPjw6O/6QWumhq9BOCRyQFz3Hc/7RkN7KfV
7ZlMze3Wwcr7MRCwRkwT0XogAkeBi6Rt4SFrjlItUmPMcUPj795ZyG9aAOd7aq+j
aeKKgqPMbcqqK76N6qsmzbTtOgC4Csw8+W0Ilg9de/wYJIaKn1m4oB8oL04iXPYT
+V0X1kjlSK/FNT4ifYRmfosG3N+TAxUutSDp7IgcxwAhnRcGXl4DwKfNQGWuUMPq
tzi7PzTQWKP4VNypAUPmGBvtnamzr+B6OLxFpaPkmXElcZqiI8I3W0SZaRurT6i6
zqn3prKBqvX1yq/HzO/KgeFdhsXMUyppAHJhUPV8jAmm0CVBZKF0iGUTJ+3+9NFg
sBG95g/yC3Buu/Es6Bgt352DJHAgQj37n3913+Q4Fp0Gc/Ct0o+dFcmE48ISDzkT
ocKHqQJB8DjNwuh8Erh7aEqyHAvxxAd06fa4WkH6ZEAk2iujYo6Bcyl+F/BMCQ9I
N+NG91/SH2Qw60rPMAqIwmrg/k3jIjch7Tqj9Pfw1nPcgxCAky5JftkNYgF0eCTm
lj9XX/BYSVCv/TBm0zU5P0DmkZvmVYbSjNch17mbBfUfwoUPiUg1KPetygpToHeA
GCFR7HgLoFzeRp2hvjpRuutQFeKY6r0dpoayRlKpgn8jYLXgGcZ6kvYSYgu14L07
U7Yj02Qtum/azFEk+JrLrx1euoyn3IA4Sbt7HMj6gRDuW/Klm7QrHkQRLVA2x5xK
EfiPSJ9qYLQUkeGm+3Wx4NtzUkeUbvo/lKaLs4moyt1zoQvTr4DEjy7kwL+wGJHu
1k6ixf2lYMbRa+2O3i6VE9loNjObKMht2WC4avSEcReyt+ZEpkqABIZy40X88kEm
1dfNVXYJ4yKsQxcbB7uNzs/SaSIEWjIJ/DCb6C3qN8MrehB0SSOiRfJJuOsrNZSG
KvVF04CeIbik2WtOX9sSEPEtAhmQDpGbfttwEaUHiA5ht3D8JfRq5BH+8AC2d9MF
FklYIc5DeqxxSU8ZyczWZqcxLUhLqH5adJocc98rZVzm8KeLUsPqq1+isnxbzftt
fetXEckXmA1vLngJVtJBJ8abZE53OynQ5f4w3I6KaxLTqu7dSAjFcs673wox8UKc
aeJadJSSJTUi+vkFufMt1kKLQHvjUwLcrOzboR6nBqKvFS525DiamvBP0J13Di6j
TKUhn/T39VGkFEA9Cw+MR0GbVJRobCjYocIFRHucnU0UbiYm3NSs5Y7q3LPaoRH4
ExTLQckDcbtXYD8DaOwo4nmN8qyM0Fw7PLNGYHMt4mZhu8EpDVg0AIfbiT3xdeC0
plmes1mgOZFPUw8SkjdvTPKZTKw002PGOMoK9BX3NTIwAO2Rw4PMvIoVptp4CYw+
VLQWOUkEWorp01xhFHKi1nSVTPb5wXySVacJgF3cG0b1YscIy0jlEF4ncY7klqm+
+MfzF/HvhZLUkq6NdWrxuexG08SZEBzEkwvEF6/q26nmJZlwntILnwZrrSqAFGCH
kt99i0BvRU3dXHm9IopEufCdQ/IeNAAOMLupO6CTjkGn4bARnBogSdUuVNwoQjGh
xZQWmnIx2RmxnnXBP7PwDEc6iYXutC0btjW7u3u//HD/hOTPuCqFH5B6aVQXhFAO
fvODITTNV9vH1+Rc227aur4e4YI5f2k3z9n4Uapy2XzeoZfOG0Rf2D7oufhmEK/d
n/FvskFWJlFS4Yff66mM9NTS/OoGsoM6f7Lbf1q1h7pVdGpLEwwWl/9CNSTbOtIZ
gE5lUYz4z7G7DDozzgtqLH8bKZnpevS49oG8ldLb4HVbbSxE5qJSOelKiM+9eDe2
WGw9hOWMjr9xETdsAyfnwf+CyltAan2MthVIjWv/1+oQrNfoAZk5P4CebcRk+Rp3
UqPsFBxHDtFomrJ4iWKotKt8pCFL/jLLIKNJJlBFKpf3MEXSvltN29XWDDK6/6Ir
6OnYyoxEPTNJTk8Tc+CRnEh2iqbjGytUmaJXfbUbKPzdoJui8/11TTCMWVxGAbmU
KlgOC640jc11bwPcKtnFc2R1u4TcmSdsrMbvWnJOvSB7gA2zOVKMNM4Vzavj5HyV
SRp8SkFEraOjta3GkZg3uCHO1lCwAYw6PEFOIwpXCdiVWhYFM+NxiKPK1ooi8qkg
N0fKDh9F2ltJ+d135qZZJAS9tqbHidf4L1QmKwXLrweG1NgQSRablZsjbwrMm96Z
`protect END_PROTECTED
