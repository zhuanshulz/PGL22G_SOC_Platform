`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MJGNy3VP9+q97yBY8xLnFUePRcjTDLRdRXyR5VTB5AiKNYiEyeCcBcQ7O7GQJad4
/jR+79+TSjM8KvdEiYpKjiFu+vq8Qld4vUJM3svvQKbmfCDRholEVAUMMJoOeaDj
KQ6WpLJdVaNTXkNfL7XP9ZL2PEeoe7ZGAahSVTu1mWaV0vgU6/Uh5Hc5dyrHvJgF
WVoVwHl48tiHVctW0W7kyGNeAKXC4CNoRU5BSkSTDGUNx9hPmPkj52b8AXHMSbR5
1b+MPsH0zQa67tAx64tu/JMjqxZ4dI4WU67rDzYtIcUHmQrOqAwdv4wIDNQPHxBJ
0lic4SjMPlUuWocgNS1+1+XbLk+onugVwRYxE1u3gup1hZ/nD8j/uUI9H/anxVzK
3HGLJM9UwYmJFn4bJPeP+A==
`protect END_PROTECTED
