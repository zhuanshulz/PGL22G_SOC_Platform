`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qma0BtZZV5Dimru/sFR0BtYkEJjLtqNJBzBBCbVFZSGLEOYNLdDwz8jtqJ2JBO7r
TsDNMd/NhKsD96hh1NdhcMszelkp9nXpO2jBB6efR48UfGf5wGSdHDWs7Y2IBupu
NyMv2KRdPA43ati+cXoGIMFjjxWX3wrFoVmwvCPAWcowoQv2oGphBJNdjI4nd1/T
fOp4NZSZgHICXk1duZoqLX+HE1o7UfFlYbvpLmQaMaJpJTm5jclkBocv6h/O199/
n21UbjFIJBnCroLUQbtZKovPB0PXXL+cyP3ZjFCibYs1hMhcW/Q7BfQCwV58iE2J
NjttmSwfu4ZLKYukVbkLmVBNsIzL8s3kKXqbc1l4m+jCDjdjYBJXSlytZXymdR3p
UaFRuyO1/puCmKAXdutKUISfm1jXdERnbJOrSYEf8F9wA3QaXSOMKBmfTUH8Ziah
Sz2bbuS1nDP42eWyFv541bsJknHqQ9AlHU8pZlIVnxtTVB3pJdEuhAYn78JDjJxc
VwRvoNx+Jhb/k2UEIlDYipq45u/wCGBMmeFXeUvtLxAij1+gwmIQJL58LimKZxM4
82TYnFquoR3elaaEs7dE3fkdKaSW49ExriEm+sL+MW5NeRHDfeGsLzwxleDm00IU
EP8YJr7vn2F7ofL1BTD/h+tXdYnTc0PZyZHPEOrMzMnFwV5FW7DlTPpuSdf6gy6S
z3Hp4BG5/Kz8k0ZK3zJUAcQG81RFDCllbLpFi98IrDkOr9vO+CpIfROqYp/ZKMAz
Q6MBUXlAtQJmc4WvgIwg0DSFnt8ZGG240ntiMipbpZhHXZ5AvLx76etbdam3LDID
m36mwIT+MMucenIa1yr1eRYybq+HDbeeFmEzPPejqUyX6totuBAVSuQs41YqvI+7
DvInHKZ4YlwZmthntrVkzi/LlPIDZHIrzN8eSzns32dJjcUm+V8gkQcG2mbk++HA
BThorNxATVRhpOguFqqyNXVCL13A/qCkjatYcXKx+p3UM5WYBIM4MXwfh3DAzK7p
RjVDZa6XgXI4QHx9b9GRZkHJpqtfg8Cv18pDyO3L2HmQnFsHLl9sD0NqnTQhK47/
kzFMJmn0fIsxYO2bvqSzwHTG+CyAe1ZGZvM03Lu8qcUmL0hqKLCCvgVZ8gi41TpA
NVswLcOTgzxq8j67JeRDxi4f0t9iz/AGNdTwCgX5wIPmy0WdHx1Z+MnsMnNS6cAR
cNIUBEtBDIw2Xny9i1jqjGW4QVMhzTTVOzB8Egzew/U=
`protect END_PROTECTED
