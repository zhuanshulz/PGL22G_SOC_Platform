`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SuLtaUB6pPFpl4ac9GKaO45R9PCUbYGgGKqCW36mcrxKDke+n3ydpThFf6VCBFnJ
/2GF7Lke9dgH2uggbpwDiExt8tJzJro71pRcUY+xcQA8Vuk9WVcE1ChaUQQ8x986
NgT8XN8rFXlJmrH7ZxjdCiq8lbEFOhzoV5ZDmmWrBEOdxEBZuyufzL/6M8Mn08ri
h0x94MdOGaKsqDAr3ZVSZMQv/uOIdsZOw2wYSV5GhA6hB2/UKQfrTtRGc8jGXuSJ
xIdfJRQNanU4IETHWS2NYyc2/5E02joTYLjC0liGkcRuUV/kci5/ch2ZdUpdU/gy
JxGUb5ONdJyWymt2DBvdIo/r+HkshIQ8jAq1hcf4xWG3s+cmm9wHhjhI7bxlP8hp
uge5sPYGm9WxrBuImTVNcYTn/REtWEMDXH2CVNcWLW+gcOOTPT6q86s6eQIusctr
Ar3rcc0xPWZnF70xgJNA+xqbBDFmp6JACiJrRSLcnlC8YlHoE8fOQRkK2kcsTtAq
9xW8DDyvjXdQurekacCSpiiXb7VMsFtAQPp83E0e48Cqssm1uPB8uV4kCjlZ4Svx
rBfS8af0v1uiKu5qU/VJnr9crkC+a/0F6OH/6g6NzZTbktBZBNFJr4Q9g2N1QlrU
kgh7oD2lajZehV8ta5rKa0/krt0Q4ZFJjmxA0Ss7GvLqHgdADET3UIcHJHZmZdt9
Pt6aCfD9niY1T10k+lXFYkzyBzV6JfXS/F6yBvj5Mdbh9Bxpxifx0MKkkabpfvP/
NCO+xI4iYfXAnlBHZDrVYP/Yv6F5+e8hCvXcsGoJXtXKH384h/bSGzhUJCM4EAy+
J3aLE7wABE6og4LQ2e0pNcyOUGQ4pwnrVjxW6T9snkMdAJbp9l75NiPTyyz3m9YK
WfoY6TDb7dphhj0VK3hQruIIw4D6DDL0v9RJ5cnk1SMzs72nxyii+nEThBh0UKh3
bZXvof3d3cVmL8XNWZQ4iY7uKSF82TEbwh58e70NG6p/xsBtrrEMGTAkszXTk+X4
JeOQ8gagB0z6lFN7OEMTVJ2GxdERwQOdV4uwb05XAgpgsbtjkorrej2WyUXDQAVg
g0wQuBwtDR6EEd34ZrZsG6TKEpHYWpY9LGZGmFjq5Y3AbE3/cb/i4dVXzsFdrNmx
N+zEH653S3z2tZV+TTvWXC+XWX03ref7rnqnpaPEdsVHVZXJ4q+53Ke/d6MSg1sg
mz0QO1/HWx0ISvPenJbeuwfZ6bY9hfKgSYDQk0UrlrOzFTqZvnEyafdKZdkOCPe1
cdBDfm5dqqzZcG8KWKGJQ01uDFT2Bl0Z7PpdMhSET7Z8hO4q/nCaWRyYrVzCoNF/
3TK3xqsLTNLwf3oa6RsKwdEJ9xsZeBV3zcnE3kO5J2bt2DmMcmcc2INPuc1d/KjU
mGiwGWd3kWLE3jqNTxSnwOHwoIxReJv3659ZKmSizI6Vt2sKBvvgYnBr9M/zXXyM
v/rIxhGq0865k4t6pvRyPXNpA0s7o7BAfy730mugnE5hsT5f/08jVGRJDC1Uihk5
m45IsFQW9Xatvc2xIiUX5ffhAFWQ/PPQp7iZdRbSheqdijyHi2ajw5vis9O71VYe
D+SNEMivC74rlZuz/4/npOqiXv9dfScbBRyRo+6nxlk+TECJ9cWPfGqh2LFkIU5Z
BP9DaSb5oqqRAEnjTSfxjETD8T3osk9S5ISD1ZXI6fkEHCMzq7ULMBcsoWa6eRIW
uLNk57pmVUifslPkjEo9hyWhLiumoMsF/4ptnP461irpU8RencG6MKl3mRIc+LPf
hu1GnGEEGmUcpEyPP81029Lygor0T3eW9OrI9LdFNrwoVk+xqIoXHjYvf03h/sbV
NAQmwm6bJpGLXzVHTBv6Mee9eKcb9hanBnK7GNskcaMO4x5NA5LpNAhirTx8mgJw
4W3HcPNagMtf7p+OzYoHtSlpIe/YmA49jPvvs1TUKzcGkoWS5mieN7Mbo0kjZPI3
Ur8Cmub4J0rTsrOsUfoPVvk0CMIr5cRko/XGJSnyKqcjRv/52wQRfKG29W4CKSPn
CocuG44X5guE1rwXmgnny/Bu9HE02K5Q9rmv76fPZFiafVBGjh1y2Rpo4Dxd1wC5
KP4YeN6/5aJbRaLn4xhaSKe7NK9C5bxFtsoAAlJ1d2tl8j1rDgADtUCp3xW+q6fF
LVgKBITMvGESo7RKm60wSFT+rItxtVgtpWtc8m3yNoOZOJ3n7+6ZiaD6lf7lrhKD
8lhIeYWOlTq/5jFG8jwKgVEftiw73+5n9XiG7yC1Db0CGIkHwHBvv8mCu60jKFuf
mWEuB7Fz/ON0iq6g/DUdn4swxxUfKsdsQrfNy3PtQ0C9TWjPwIUzd75s+2M26DhM
Ui+IYp+PrOXXEas5iZBZg2kl+/xCaLUZH9H08MryOgwcVxdQVRgKihHNLMguB+up
EGzUEE9lPmlvcle/zRp2DST726Vh3gRtzj0ucsMVdN+BbFGcYRlPkLB2CHt209P0
xKd5Orlc23t6+lJy1C+klFy9tIqsuxouBNoanWGOl8hIFIxrhxwfISyyV4s9BZCU
MHRqLWrqD24rXN6/rpYRUIxdiRge4WzNoFGUDR9EIT8AxEYQu/k7EYZ71MwWFrgi
ujpAlFytoLSOvc35C7sZ8IDAZH9gobfHtLQLFqUhapk6t0rkrSuA15ZrMuJiagAd
d8kSeE3thP+0d8F33k5hR2cXdy47g5ZTtEf0O1JK/BiUwiDtLTr8YCtbKRq70kBC
d89TE4skMKypdwT1sNlwbB1bbMlmOJIF3q3qPVJOIJcUk/oIZkQCzaA+VOdRHIjO
XTCfzce2heYNYxW8/kQpdlj1HIFvfJKJ96lXBwm3JCEmLfY34ubwMlfhXgcmhWjx
mRf7N+IcTuMHYbsyLYr+7A+wgKFaw8lKfrgoJwGRzfVLXdL0KLa7ec/6w089haTn
963apRKA9E4mtfqTbyqs1rwFpZrxOjsht1xCt3GqltCnwiB9h6QHUex/XOpKpe3u
XpZV/UHb5FGVvshuKsgptDye3QpGDtSGm3ZRVfbdH29iUdA+LLs9Y5UhIePG5Qmw
4HQQYUa/SrszBO4BVSY5G5SSaM7FlYPD0QJyUTy4Cd53YLn6UET3fUer8O8iAFmj
cN07Cec34Av3WzX0KcRMuZ0dG62OBUcLiycfacremm40Ed2jeJbsTNOgS97FpN+y
7ydro3KrWnXeL6hj9iXOQCFP9GE6pUxIr6ub2juSHkCtTFHLChj6XRL7enHo+gY5
UCIPhgfgzBbsEGCSjx7Q+KdWPbrN5/DaR2eJUWMKFQHTW3XOYHwu245gp7GU0aWc
m2SqRf8bj/9+e9hjdI38e/MVU1isyi2tbr/H7oSTMZCNKwq261PgJ3187Ct+OfW3
KzVg+kMVJHC6GlncE+v3yS0BCg04Ou6R6dXWzbpP2UoITZ1eQa5vUcWgX2gsZ+PB
09YPAyQMPKT3gSmuteKsjTEimU+ohGjzAjji6ICyIMEHaugsNOQ1hD718ZPClsmM
TPX1aRn4PDNaUyGFjPUZAZ17sZZsP4UU1T2Q8MZiccIuKqG2fwCtOcFuBJuRqSBE
a7YBNbGklg0XfzInDzqe5rRi49wxCRhC5lLFvX0hK9iP3+C/+NbdC8TzgIcyHsob
WL4qVCHeu8s3UE3uykqg2XoTABYmNDCWXwN69TaTmg6kPZIy9i2t8JWpVBAgbyl/
t7cemc+ZM1D0A5fOu/AsEuI1x0/brzRcCqeJzOfDPIXKXNL/a/q4lggOQuiXmlz1
wJB2rqime+ozaMqdcnPvxWBJx3UFkD12QscTqbnMwtLEgh+tSckcOcts4MlJMu3J
oTQcij6DZrDlslRNMBqMAvDkqyQTsi6zQ0yxEZYGgP1lnspsVIcPgOywhNanBm0y
vIcYp5lCn/kzgPjUwaMkxGkSLTpF0TaOGHGwqCByFM5le/qe4pebRuA3rNmY6QzJ
duyB5P1eaEijj9Jjw9VUDD8mtj3qo7k9r22CDVDGt9IAaC0yX8Jw1ahuaTKc0ChL
5VO+62qUb8L7JTNXCBEzX/DbqMqkcpQYgrgmBUvEcRONzY0ZKeAbgN+T3fRqhkkD
R95lvtL+SBXg0w1g+pCInewkt/D2i8KulFAcPC+Wsc7h/AMtLnnwsSBAUVsPXq7m
CdD+/+/XKnPKDCLikbkkOM5V9l2iJZnlqv6Einn0OoaZhCE0iDkzuN/K9kGkFF0f
WsG7wWMGAf0uW26Que3ICY1S6SURT5g6ZhGqew3CuOAbrOHLc1W5tOTGhoMmbq9u
9KBQ4KNBTDvnbu1pDckGG2QqgB2jAE8WL5WomCYnT9wujVV8Z50ukGn9BLAos2ST
QQgzK4T6m29Bfwo/5CZ7CMeT9Pt8aIPD2UYzWQQuWgHKzEAH1AeudSuXcDNpm+6f
672vpU14oGViInb7V+qMg5MfkcgMCkwv5hM7zjr23L/CH5Q41Pa9Gym33N+9/t/F
8zn+g9QnrR+BoUqXGU2eFHsiJo0JE5/WKKmD/Sf7A6cpmsDFkmoW0W1+30dZX2c2
BPTowO/9S3JzfEyS1h0nxxeKjxev4YqrbhdkNMllaa3WRvdpQcNm5t93+Uil6gTb
tZ4n8YWfzFKTb1Mp8Zsr/3So2wZ06dftl0dzlc6k/WlJJY+/NLuveqvKUcdYd+09
JC9Mfn43BGHHLcUdjw9dqsg6XUyvU4XTuq6HxM1aMEScx/ooiEymesGJS5JXWKKq
Ie6fQh+ogTOuWN1Y9ASe6BP0Tl3P4X1XlZMi6VGtuKTmafapNFeGCFZ/BNIQAhZJ
jobE1yGOtPh6+MHXEui2vh/lC5iCU3oDF+im/+Aw1c7Crjxff9hJskhG4e4+yS7e
Ihh53CL2rwucRGwszZhNEXCxYbuZkM+cCaHDtKZFVlUrHCjc/2tLdPe0f7nW26tE
tZu5HchHUrMXl9khdqhgTnlYs4jyZlpaCDqQZUSueXI/adVcA2Rkql22W9dTWu/O
GuPf9a0ETfRyHp15CFm3IkVTpaJr56D+FtxYeOG11WrFoLTgnZF9Sjaf/Fxb+6vr
5XLnXRtnU+JCiLX7aSWhGArxnF8QS4Ov1L+5LPiVGYK/iKKIPM660dq30n4vmE0o
Z69EzgzNFpw7aZLP77LyoVKXAEr+YWH8W32RbPrrfdgy1E1/FXBwTwsSnLdUiyxJ
mmCbdDPm4cHDRdyBJ5Qy8heFU+s+zjI+OrR9yfFw8GBRLltPSW7bWnFC0L9VMZ2H
h3S23zt1BYJUKV0inxgO/6S2i7gMhZbVjQlLNbILletHNRIkMDa4RuTu9zzG4C5q
a7YHY6X7pgre9nhFyYOWyd7Ys3+SDH1cSuw37CjF+GF6zxrm+EYzAixO+psf5Vsj
nSnFGGJmUmx6jesxglVS/Cyq3gOrAFTheYsVMnVoErCzXyHHC5eMue0ug4Psi0Ta
sAOj93VAwStbj4TC6yX5bbHjYYBW2+fh/XzburK52lt8z76SoYa2niSkiFXmrR2n
p85Xbw2vVCK7yxagoAGHaPZ8EVgQ+x87N6cJP2Bdb1JQCElpIdEn97lF2ejPbtDB
LfLAvL4euQ7Hz/C8xg0I4wNoR+OdVWdxRmoL7djjpl6xJB2vEg3d5JEeiwOWhV41
ojPHDJY7zunEeSNwRm9d+VcnUQQ1RBCFYlr+loMzmHJPWAa+pzIzUXjdrFKPUvsK
bDe2ABOlZDgWS/obiithiOgdYz1ehaQrk5FS1XKpDiYk8XK0YIAjiSnpgUDThbjg
IbSvYjN4hGqn8HGhy8mu6NTiV3kBc0d5ZU7c3nNtPFaRx8jZOUAQlHh90RewVgdm
9PaIHqklJ4L2FnS3/KLD0wJLdUjpilVViAYiGKkPaph4a79YomHUB2kgZz64YYf5
FcyJFVE0De45pRe/VXvo0loHuxWfj770SHnm76sMTyw5c4dv9yEQOLcYiWrwBp4g
QDttazW/qlP+51WH+ttXFM+OjSPWZ7ngqVCzC4IFYeviNem5bL2NFZfXC9AqX5hJ
9FZBJnxngFzOw4u0IIfedZNgWjf51CEFEJ7q/E05xH31H4LrSaUuUiwrF7PPpyPe
CR9e5QV4k44XTL/Kr4KKdUr9cYVpmVJZrd93FFsGERXXCwx2STO7PK5V9gKlq1Ki
jpSjgQapI+xq8dUgMAdqf1HIB+oNCqyUNvjoKlB9c6ZXHEZ6MNOylylP50dNeqcn
F0eRAZUtOQe4XXEmDV415cFVWf74H4XIGicSuaUhuIPWdHMUSBaP+cwWnQ6tS5f1
TaaDyS45LSge/ASOfryvZSVTeO7RbN0mdbzSsEkNtDkZb9+4L1y9yf7qVFUHRUfs
rClMQOkaJJweV7JyFUCDJY8ltdp8zdhLoLl21jXVO5kYJQAINjJu7etHmv+irGyZ
G1Ss9vJQ0QZSaDP0vZrP2uJh8+0LebiD+Bd2gLUZX4CIXfQJ5a/LwYPJE9lqIlK9
fPR2npRNW1k6w+aGj51Q08pa2a5dAx02kIk58JJKknRIR/diNRHg5aeH+yX1XqcU
5yUKcHd9+w4ET/UVpfxovvcod2QzL25E8dfMTuULzo0LRVLGXGNlbePC3HS5k7PF
/Taq8KKA/DFZP05Nw8GsvX+/KbdAQphYvU7V1FMqhbcsoLf3oNY9a8xbKs6tQqTV
AR22MPi3iIgXVjn6H6E/rdgwI+9n++NE5u00IwR8mY11GYFoKztQGB2/gaNFZUEV
tBahU/ZN6ZWDeO7LQdZsMaIXO4CeYfH02ozbfORhfCs5UTt21pbhO2z+L2IA+dV9
0B/ASzevLcwrA00ha/reCIfh0cgj6Pyz7/VGo9P7h31MUqGPhi58A7PkHkib+tRD
w/XEwF7XbDHQUEHunFt8ez4zg6zUmIFsKDafpaH8Ru8GwZYDlBvXtrov6SPKppD9
0dNRXat3SXSO5/nZIFfMfU7s5rvqGHbIgcFTRxn35Bje9XuXT63DvyBPnFno1FpH
+ndvNqAwKM2zJuRv8Iuls66J6BesrXizIzbzMacUia/B/d1O4QnpSCwRfEIzB5Ca
LNxX94cSTlpDbQz+sNiGDDr3xDRW7cDuMh1y5D/CsDY1G7IX8bDcgw0Cdn5IYbh/
NAxW5tqNljtGPxVzpZV40Kzt9f8LMv4smRwxQqptobULjoXetcbl5tIRXZ25aoCU
RNg+RCp3u9k82XEQsNqXcusPciklip4APRhQSg/0dP2mWqs1mMUuUv1UyWX5kVm8
12xMbSlWFC5/rxBjvUnVp9rEP4/wHYU5nB2zXJPd0vuyi49aUzqzPRl747jLqZQM
+J69+x6kg4KiGpPV24BpTttis7U4xwhoU9DHovsK+2UP6eRF/+nVGzBaO72Jl3/j
x74vwZMvYwUVmzqDbCnz7fpdzk62h7FIcwbfOzlPDYiwjoHFEUjk+m4ReKrhKnzA
9h1EN04tTkpIDNYxLUKSmbxCSp9gH65sRMwUXfcNaMrnFg9nSKMBTJIW0aWhXdty
OscrrKeIycDGHdC4JjwQYYxyF73Mv+Yemw1qmS/Mvgx+/JsbT/g9/O3RElKG6U4G
3rnhgZQLhcam0w5l35wgdxDkA8QjJLwfCL0zBB1gWS0QI3yCUaMBTjLSmegB1w9H
Qk3mYuMJD8DdmP3NkCZF/eIc4FruTULk3Q/1LeX+mV4SlBE4BQTAAlfojdExR8KO
YB/zTVBzCquRSICJTXL7VVXS+0fsumRpWEL8BbNsePLngg5ObekAU/LWfdHZPdTq
JbR6tQIo+q0rxdECXti7rS8+3U6Kw3ymzUf/BGJh8zURrn9LG/79D1pKbOu7Cw38
1oK7zMAPMkZRshGkDvbo6XXv/gkHu/YmZZaQFEspsX0zGKU3HCxj7julk5AcWyWD
kpm1Lx+k4M5TJhYQWhvxDgfO667rTjaBRZPlNlW+juCmOMZCjjmuZ7hSmaakj25a
HCiEL9w0TMhiRbLEP73IO+OXg0h2yGZS0KdNquyflt70pssZMcI+UnzEKJLJ6vHY
U7pKbpGo5VnODrDa2rn2lcQdaHHQSfM5BYtxQbiIW2E6oYjiLfEuVaycKh7LwJyb
ich3shge4q4lwO4Z4tq9NHxg8ANsSacXOmc8bjJ806x+XL4AOlPlQQ5kGf080KZ4
RuDZrX/2RLSJiu2dk4XV0/s1+9K3M9BN8mcyhe+AFlAs2rwB+DaSbw6HWNj2rfAA
wzzBLuCNzYzdOD1z/l73Kkda+9RCz/A/V9GLWwNNdYTfEKHkHtacImh9XZMd8v1g
Uf2JDIOsUTJ49mbhxMiFUyeIyVFxkJzZjfUhWkUqMzmOwuO/r9zvFgxgzm5AC8GS
iefk3hTJXcYPabc3cyGS9JHrI/aLABwM0BZ4sxJVn6L7gNXKAKyHw3NbVVgB1dcw
pkJMBOWUzGLZ3n+zr3pSNtwKTwJuWdjhCHRldKculJ6PRSayeir3WVUnjY6D3Dx0
cKjv2PljjRYrQYzqt/kYbN+r1A9FASUf+sXomwceaCR6aubHaW5tMl4KhKmV83Xf
m39CVhMjg5+5U4CjICcFJw2b/NdEnP3x+hOiLN9FNs54MIYfbjxjXrtOmGxiWJp6
BZSceUhUMyxZYsJVSyRRXfwQwV6v1wKaA322KLtARuqMgNDGXVekZEHrwmhCrnVL
GE2Iiih6SbD5ng1+VcDh/ISmDe38ie8JxJWW5WvPm6L5+Go9/fJr1BqrR9UCTo1H
WogbiOZg7i9XIBVELNv3kdJL7a680r+A8zXbuXXLA9smGcbfBXTQbyaFRzmAoT+E
wcnRZF9J5WaTwZ58CJdv5lRWTmKWXz8U6QE4jbNf+/LRySLQmyqTvqDuB/n6fBJR
0HpUftJ4GSlMv1bhxARqpX7GtpAyDWIi/XdUc11yjHh4rnW6FMj4ZXEj/OygGyTP
gxbQz0NhsZf4aVNZBfUlZZWNbvvC/rN78ZfanvhVyq8eDFdqBwgJU4iptNVk0m0q
vbb98VQxSxG77PodzkANFtEXisaLV5949aP7yZfrwKRpTkqDmYAA8/jlEI7DxijR
jgADvAmNidNz5S5l+szN6pI1dZnh5yNdhwyYDOAszrzt15jvIvSSiLB95XeqN+gC
6mJ5VXQ15Knk0DjbNe5fs171E9OzF/ay7iYrVZESydHzAQbkgCAXSFPv9EKwwV6d
1r5ueimh3R4i0VnKjkqbPgWtwph9EqAmtu4PS9oA3E+0MCa6jQf+Ool3ClKXxN1P
MAHApBzdkIf6TOFuVjuE9GN5UVSRHUyIz2yMePheuX27csBD00S/Q+5E+YGK076y
DH0Ur67+hsKNXaOu1CjYej5FNqAAjomj4UWekBVkBKMoWYMCoxCN9VJ6KB7trF/Y
kDCvwt2zCF0AP/+gqVRSXntmtWF2Cxlc7NzS8KeJyodk0a6esHWQCXfCtrVwmZ2L
72yDLHERuAkGlD4E9Gm6xf+iCbB6MLifav4BCnpXrnhnl1ncc4wM5KGVzuB3fOIP
y4HAsg438bmUG0bNLIU45s2EwWA/t6akxEUSpxl+pnJ7ACVs+xnyfVmsU8AsqvaP
ajFaj+oMAhmDG3z5Jyam93cmP/Qi58CclaHlEmR/kgCCJLWoadSsfEoQeqmcP6Az
PJcR/3vXMI12r5JyTk828ar/+a8okTFkDc+PBqLNzDW4dG186Ynk+QA6oQfpcQFS
VPhO5UdDapJQB2B3lH4zLrYk1JKu2oTanU3eOVQsSkhyQuM7Z0avV36OLAdkiU2H
8SVQoMd/MCyaRwFwPeIc3QkN8Db2381GH8mnLFUaj4JrBm1U3rAAMMSf27MajRcx
Q1x3JxHjNup0nA9mL0+bcz7PDmpi3f5eGVGBAJDlmZJ9r7mqQK1YrgZzVixxU4AV
ADOGvya9ur0RL24G4jTrfBj9d4WRhsnhmT35y+gt35NHNVvNWUTdMnfUCBg5fsjq
I3hHG6z/gfjBVSJ4WojGCMICPlrm4qz6NanYvniq/HXeR5K9onak0otjONc9OQVh
wQKUhZxv8bq8idDZKpbxX/I67tSeKIvrQHIVLuZV9yfp56rWsiqbTX8GEjm0rhLq
haXLvHC50rKwmYVCxh8XzzsM1uWa3oUN1HPa99nSbJzRbxuTg20p2KIgf9bMlHwr
S6hZ6yi6Uk4HbXHmio57c/r1woc6BY+xXf7bRXfTIiIIa2Qct3t4z/R/15opWFPH
UXki178xXa/QZLlsMDkQa7oxEzUbVndE7D5OUiQMXUknVfdf72Yp1K0lTPbAbw7F
A6fLiJBeQS9Z6VD+ebftMg8hKIuknHpX9YdTyD42iZxVz8IoxWQAYNL8FU3AxspS
4ir7xmz2n8/nKAkFL8scXBqtn2Ll/mxxxltRrpPeNEpLX4GalSLTwqE1fzWHe3+m
8XShd6f93RJU65G19Ll9MB84phsLsued2r0avWrXe5jFTACuBNfEVLE2ZI3Kzxou
d02lE410Sz1wH0T/ycaVK//ipXJYVkiXahGcx+j2ptjmSSrFTxOyGwJKQ9dySzQ4
/QdQwSgO7Tbn157Yq5jlFw0zjZkXytP8oPXONmz/4c+n0m5DpXIrv9RrOpY+d7+Y
s47rrxb7tbWCIA+af65r5T3qhVvPwSYwom+5Ico/MdA1K7I7dcUAP9+m2z2RywyD
PpuD1zhKtHOAZZIbUu8N9O1KWX5pg5nxRvLG1jhKaRgx7rR5OTjNp3bl70oaCzjs
Q5S9JUJE5ImsifuYjyfpQ7vQQDCsInQyYCCfNkHcEYSto/pI9x5EG52SIlTpqCOb
EEW59+YRLM30hAJOXVa9vpB/+aCTVQHky/eQ6SO0FPGu/vF386SsZ6IVhUGPIpjh
7GvEla+opBC47jbU5M9SeSSsfcdv+tZhvtfPPJsjeDQTUtcbq680uz//zYTtl7+F
XD4dM+0qYMazuDalp9Z4c7Twlx2iEpBMtJsii6hACHYl7E02BCdbKzC4Svfzcfrv
8C+1hZn+hOOMydkzeb6NRARLF0NSO5PiIEzkx8R7rc1gJw95K/k24qNVJnZ3N+F/
tLYrCwuTpnZC0r4bBSHL7cPaL414IqXaLzQC/QCWV58QTEzE3/xMXeZppCtyNHhI
G0fpDihTE8NHpOIJePLh8SkJl5vc+ynMWcDXiEdP1V1sN7CsTBAAhGDZA/ApXGEl
N/b5iB1CrM3kn1Yhed8oAQ8jv8uCtmGcIjx4T/IUOc8zzg7k2QEeARVfVzdLqTqa
dY7G8VKgP4By5eEYSp7YKJkDI741aXKxxdFJrQKDpH55xY7rq0xDPh49wrDeECTz
kKubCCbMNlXcFaMBoZ++ZLCtIZSmVkCA7oT8IeT/LywII30Yg8VllZjqXfnL+Swl
9r5rbLlQbzgQF3Icn+0tRAzxgOYr6aoFlwxjRYW2yvivP8QqJ2U6MK+lpF8i9reb
uG1QhBpyqHhafzMCqCtGNW17HWUGj+RCUEIFwGlKhXUWOaE06VngIPHAnixYLDKa
gcqzsqTqnC1YDbhjJ/XFu7lLuVkGW9owEJnyxN+Sug45hq3u1ivFAKcOGPrE6Hqe
oWRCjDSIcJ4iO89Fdk/5L7v3bM45l89r3VFo5AByAtYEYfcd1WSHuWN/ambLaVb+
upxBTXU+KLuzz9/9AkiQD31MUKnaAPlGDldtn3Mzh6l2hRbNJ2lAjuu2Eax5kfO5
CM8RaBwuEs1MKR6nKyNX9Ltuo8zZcbOqR/TaMHmQwq4Ybn9gywqTyHW/hkVIxSFq
z766blOQb/vzMFX7fZzV54spP3f8MxnKkdkhKyyUOEAKjxZ6Fj0oqY2SRrWLQO2O
VJD4LHJai3SFdT44oCctmCDIDtyJymRWa6LKbmLctUjN+ZlOONsMObtXCvSdrZ+P
/C+8GXl2rO2mNBwZJ979G6buO6Lv1mYizyoBKS7sNKwoFLheUFJZOZLUtGf2L1Fx
KAtC0fLd8XwjxIbx7o7wgaX6mljtwIWiiLtsxfs/NR7ldrw8mz7ewQ/sIYfw851D
+8pJxuCoDJrm6h/U0FqM0ok20caVSxK+wVS4HLTYwM31Dg23fK7igFKXgfsZC3rJ
gLqB3q8d8pSmbGS+F/wYcfSzjEAoowOGQa1h+xRiL+swg7QoYRuqcjx2Uy973Q8M
IH8IjJcaw9MgEeUgtlde/bWZ5hE0varjSsOtYV0eyM9qW10mmyFGBFCBSzUWlHZd
FhfYu2A4DxIiwLJ8aulCovCsXUNLavBq+fHu9RQVqarPhF+3JB6rPXQQIuI1Uyx2
TqlXAuNpGe/NCFM9gTvjCfseKQmu1kVoiiGPWLli/sOV3wktfLb6NYPbb4qeKTx7
0otByIl25OZNbrQyBmZaLHvbuLLF3YLgx2HUSgDzg+PzGjUTzKGj/oc6iJI7Mvw1
XL9ui+So/L/n460S8dyKF1WDk4roaIF/ZHbTKjQjpRcCBAJ7TX00g4zRks91lpTr
/RdrIPTUGK36yDy6QJluIVSR/ZhaJIlPGB2PYxuR9PxLCwbMti5qf6i1lFXBZTD0
BupuNClS0+zvFLe3YwCUxiQv16ed8JcZ1cxkIJRdXJRPEuSP7EvucnJg+l5ozSqU
O/DwIymbwsJuwWqnmOd+feflScCzApmtCFB8IMsXVX7eikZE98iBjGd0Nmw7D0Fn
SKw61R5qKlZU1NnLRIf0y2ohylt+9rNLxAf78bUSXc+2h0w8xyElZitmJPMWd7Zv
298LLkh5ehO4rRBYk4+QfvIb+/iXQiPItHAZW9oX31oa11jEUSdkCdL+1uyOllfv
e5OkGoaYQeXOAZHBOJLrVFSaFqb/NkQd2f1oDo7a+1WxKI+JkjEMntE4KBY/7hWY
sc49xp2uwuNDatQr5uIAyZGx65xW+JfMljxmk1qu0dtitZH6uqbvcSDZDhcukQ/d
gB5WkOs19a6KDCN2ptL1emVz1lthSqTtPnrqDoae7YiV4Ppg5N529fldZmKRhkK/
TAd+d1SEe9BrD1PvY+GeBPdPiYeNGEkL6MaR26axxYsqVGbG54G3igMgekKA/3kp
OLV0/2vOTfAdCz3NdUT+U2ZMUHRrGhc0d35iKXajjzbBvhc0W/XfKVqu+j0l43Rn
+4A8Wg8byF2Hdh4kH5m+USeVl5wPQb43vA+HXUGAqqjcr2A+HpjV7EccyVEhPSCi
8bBYB3dL3CA9Mc6sj08pKKQRPFouvd+97oJnEGCl+mSjuHXBtTQ4E77CTEEdBuUH
xOTfjDG3inYA4SwOSph11yXXGwudUJI3p2O4hUSzrwmwZ1EQqbygf8ycpWLwJiOf
CAtu/zvineqEnVGFzQzp3bI3z3mDExb6XHBfadTM22RdWInXR5NRunCyb2djCWft
tR3CwsE70UNvKfle+IvF3oOhkxXJ+WyISNBFcfC3ewN+yQPv5087bR6VtxkOFO4C
lm1LTCXjbS5N5+LTLZwH08kWrUFyN4hoSGzrfnPAI+gnZDKLZZwFn6qkAUbWBg9G
7o9X+wzycAnVphDq6msXc+MN4CH8NdpWdySvhlq+clAB5zu8oZmXkq6e9Yv4JQBB
bEvKrub/Wfc1DEv79qg9sLlxvEWn2FREEeM7CtEr6F0n1n5hgUwcaaQCZtmOC+89
RbQAh2wyuPKq5J+zr5vYA4mRJCYd+T7QJzqI3iukaWSshyG8TfE6mEWixpRIrT7W
Q5NfjMIM77cQLMHojlDE8lhR69ScAe01J2D4DyfGwOmCkY/nEIEpGrqNo9CcD+Ar
xlJw1S3q5Fdd1azGM72QmKqRQz61IgR7kvtjA+c1tYI2+OGU9AwZTWhnZoMmHwzR
9GQ5jgkv0/PlpEMT2XyK4Oqt+mF7//U4JQOq1BuIBkl0pqtUmdDwaSRh1BL+sJua
LU9BmlG/8nI0qQUdU013ydE+/l3tlP/q+5CZRFtmJoozjr4pFI75hYyXhP+9I3v8
ArIWXSmZ+t9ySNoRhPBox+ixZQGpDYari3YSQqNSLT2k9GnQyI9ZV0dqceRut4p7
ap2FvRi4ktIHti+ya7i+opsX1r0KbKyqcLr/1YV8KBcnE006ZkJber5ApU6k4f15
mW1ol2GfDS79fSCyy0TjNggof5rmVQ/8ZJnx0qrf+qnUoaM5NskuMTYqBslkLkj/
2QO8dzM4Q3wZYz9CyNrJDV7MauG/35V1MLefpEG+YTTujkhY9PnDyEXbfR/Y5Htb
VQDs/OHZDt8RviKSXZ1VL3x3SrFNMUAJD8WI3tiQd9cUMz7drsqCB7vlQ8pFLENF
EWJ1OX2pg+t3S1jKuSBIIYprNhPi+uho1qEGUXJ5R9LC+j5mNMepOiAlqCB1hhBr
8TYsfBVbsfCjsOnUscsdfKjYqGxi4cGfup0jg8Yl7d85ywiX0qRZZkkyInyYjT8N
evPXqfehGpzdzk5JCc0ThzljieBZMZtWY4KznrqxGJELRsJb6wBlQU5/kTyFK84H
w6vRrbiz/v8lIEOcGmsnsErcYD0ahJLWfZHIGKhDUjs+sJ1T79ibiPNs23IZLZFK
sLxQrAhj4eiTM4T6ZVIF635MtcuogOjT08z51pp/N1d6iOxUxBO2uWx0pf6lsWSf
/DBC88WMewNW1ri9WPdWw7VhEF7bxW7Ixwy3WPJXboq2xp8O8T2LhPZRgxOyLHWC
Y32RMHSp3mLTlgqI1F0qaJ81NCzi6wejiG3wia7e0tu9wYmLBBi+z5vE3BhR3tli
heE5atX8wfKlBDaO4sgzx+k09WUXyuFvQOQebH7bNfhQdCqjWAgfvZJs0bj5i4XT
bhZux0FXzSLfa/K5yht5xi8D89+ExZj98vFwoXKIgyglJfWjiR5qqrpCDFdN4l4V
QblFX4pMf44Y0mqkLRgP993XMBe5e+hVBHUMTDML3uJXF694OMmQGEVaLuFGwev3
sXaWpsMcER15lSJwEAXdByf7QY5Nxjh6w0LJsTHjWMDSVXYh8oNXkW9WKOTJRBaS
oNXuvcyO9EhcWLgokYFwf31phJDT7kcWh539LCAFJ6zhJmE33X4SKPFm1oFit8rv
yzDdnyh4Dbu2Q8jbMuMoytMGTyjoHvObB5NDPZJYbF/RZS1/jvnjIIR9lFjQFVXo
JK6D0RvrHhm3ETeF9a/e3Czj46cMlxAf9hVxEAiMmRoT4Yvk9US5g5cxmfkh5F7a
MLRttShYfFPXCazyNCwLEUAiW8XszWrn8HJG50mUx212esDhufqedNRBlzKwlH1d
D5OrTlnQCM6XZQtajvd5CILfZfooJJNvISCnLtgDResM9hQImLy/uxxDVB8BHFNT
IPCmHB5p2lu/sTuFOlQRkc9Wsz+YiXkis1D6J58DIlBq5jRAYqq6Hdn1iMJpVAIr
C8OOBhZnFgEDamh+F3hHOfJDItrU0B0+SJ0xALlmsUBKmXKtXoaVwJJpXVvBanOj
4AKKIA3qgCwdZUZe4E+iCeEJaq2jGBs7CAcVNMml5ebPKndNasigN7mmZ4ArZeMG
0AViDbWZBKv987v+sT1kOWAKTFh/Lt7/zWhmamm2KrfuiXbVj3Iq0b4qFffL8xqt
M0c5fmzIoRfq8S6Mgvr5cqeJk2B63LvYzGzW0QKW3cCrotK6Gge1p1mxtsMId32u
YtV6x5qyjZQ72vy6IZKLweEvDJzOadltFT8PeB2AQHeuIV5zzjyhlylTgQPNzwbq
6Xmapsbjuh8jq71InGJnrllO+ucaw316iB8Lf2H9EfKx7vOuHHTGp9qqx3EkEYD9
pr5C8OcsKtXlpydfp8QGbAqTtyud90VBwvMqH7XJLdz2Os0WcEqMHeVJuD0tTJXY
zg2v4pxuQfYWiloBCCvj94sTzmQw7sWI4aOgcTlKEj8wAVJrZDwRLqh783ILh3lW
7yQmnRVtIK+xWk9guYBCfwfzH+/Uyq4xA/W81OIPwbvrCj8oUKDwW5B8dVP212p+
bGOj5blrdTkwcYtjKsKFcoN9lP/BND5mclCTCwIZMPgbRijdI83Mu6n3/7ycxmgX
a5ZDu0b2Yr3Kj0vzIYdeZRNBVqCuneJbIKUGMkysMyrpEr0noKFOiCinpHEXUaPo
dMpgNmJVryMhr77DKYpKcOzhS7LilNtjYg3kxTj6dvs+BN6d233ipHzBn+zn7zSF
YNkkahIki8qij9tOjRPmPXUI4v/70dL8d85f94Lt5r90jehmp13+vVX8rU0u8a2+
FXNGHh2NYsNlHw/nB9rl0gMpr5J74dMP8kZgiGA+YLZqW8yAqVTkEoTVbtMB4+Pr
e1sy7cSa6+4EnCodmg4BpGlQ8l52AfX/CBS9VB/pKWlNy9B+YKxHj8PWm2F1vSAL
T7CUyCjAAg76Gj2tdCSY/YVjre3yijASiNpRYazQ7c6l1aYSC/1aWoYp+INB2cDp
O5fhO9QnnzoKMtZg/V3YYXIXfsxVp3XEfztphzzUgrq3FVNNhPZ9ZsCwJhYf+8iZ
lNM7+yaVkYVGxKkbc/Z2JjueNQa/Yo/3GMzs0qKuWFSlDCh9xdYgMUFjXyKjjyXI
WCQFSHqb04KFa0sMn8WUwPU2HP7o8YhMcyR0KjCfI9tc2QUUe7zosX7QFRd7tKTi
ifAGM/PfInTG6CxYG2L5qjKKYSn9RArrq4pHJITtKVrvL6Wx7vXau09BGUFqJoFn
Za0L97Dfff0USQKCxU6vlCupRmq2Ml+tqgZfdxtGEOomRinjdDtkEC3qb9vzOGYk
Xj091z5sKVa+KyG0AtDX1VdanGHKvgl4DVU45X/mtkM53vGi+d2qF9uhUg5kCKrt
83o2/b1uklu2hPdAJ9kTWKQHrrNKI/nd4N8hrehhuGLTRiiFVQKw5NXreHh+pzVg
sDsXhBLPZQi48/nrWRMDBw==
`protect END_PROTECTED
