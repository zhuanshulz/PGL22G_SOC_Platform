`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+ple/bOPOx+l3MDa9+TRMoCy1EyKssriWBJtCpFcjjUyHoNh579S7RxE9HQmuEKq
tgPh9MOqo6Uks81Wa400gl/FUjJnNZEBcrCNOSSbxphGgoSJhoNP8w+LeS2C8bxJ
IjSinSI7BVb4eqhAlBsMGeR7EZFxQAqSslf4Aq0G8bi0YYgRXbOidfXrDap348mF
hxe0qftRoJnkY1SFf3wkFD2RGPAQIwFMY49VulWpYGFQAV+K5BWGndaiNgmSIdxN
wQhSprkWGiNyHpk4VTCSxnfwENzMTf7EEcThzkg2NfrdkW3fba6stzBtO+LVyCav
gMkNwtZVQaGeYQ5/Z9KTirNdd98oodPHmaR8vWYU4YdipdSQbWmdasvejT/zU101
1GnLWwwfq3f9r5Z8FEMBO/XmvsvIIfkuFpPGXrYh+6WBBhyQmEYtvhTC+xIEX4CZ
1s5V3HVqxNPkjUD46UyPQTa1eEurfgtbmkAIDEZsWzlR8Y51bmt9BjLR0RVweh9G
qsNqY0SbExD0IcQ8rmXaoEZSJ3kWBJ75g4qrtC2UH8KWFBFw1xHo/3fjnSBwSJSC
T7Q+50SUFZceVOvg4W1gLZjszMNH4plYQLIumIRZr3FAWTu5jbldEbtGct0KHLRJ
G+RD7bfBd7azxyZUzSLx3FTJ1MpUV2DxrZ5lmsVzPL2GGFUXnrrLNgQYyNSQfYq7
RGWKi8y06HW780wIrcft2bfS8WrKSsQRkFMuXq3cf0tDicedPIDmcedW8H9AZW+j
znkRXVv06Co2KPExgHexUlFQmtei69CLq6/r4Q/7f3dHk4CVvRdVn1Sai2zW1Yyf
Ba+pimimjK7dXptc5MJJC7lZkNaCweffhcZhkwe/XcVARELynD6eUoijXlsfQ5Nd
ObknIsAqAKJwusyy1eFt1JF3Diu+aGLjnQdw7p6297QvgBFZsLBaK86g8Z+9dh7R
DnbAYFy7S9iepLmXxyIjN0mHAcqC5nwbLFZl2HosjqHERpU7EPN6g2U7ZnZ+F+9Q
MhRDw4RCXwlZHAnAtDs+ivfCjh6jEUVScNa6qENK6QLkCFSjj3wrT3n7DqJtH3y/
FvbbPl0c3pCOG+/rI2UOWVyezCT8fIw1qVq99t7kSTwwvPV65Dl2fsBvDbsakHFZ
Po2UWyKF1eMOfQJcdylk9CDQw3A4AYneGHlmjCfHQ9IwtnjZz3jNq13Dy3LjbVDu
OsXI7QrBRsJ5YVpM1I2AljWDI1rMSilZtF+2MtJ0s58IFl3ThAz1OQxWVZlUv2TK
NOUvpjjYQyhirpuJ4Bj58V0sMkWdhb4JlG9AdWo2TtRoyPIKLitbifSgr3Mse8cK
vGZF5YS7TwYzeHsBp41iXinOj+wbL06bh3aZSsQKwTAe7L6+HJWo0P8j29EwNMcn
eDBdr9txwH/QV2swAEZxZgvR21n4HPUey7nAexBGeI6Pv1gC7LxY+LQvq2NcFwFd
DMnQcCAAWYQ1qqAYgLgZ/JPUE0egqBiXrZ4oJuOE8LQ6FcLfUZ+Iow0m35eFTE+H
dlqpr9yJEUvOvzHJBOFLoxMxjy0GsGyBa67u8drGYs1fJUMkQONcc8oYTcyxm5CB
fKxDW+BeZ1sm7WCVDbvW1bZSDBSFXy/N6sMBaXqF4dQ0APBVanyX0lvJWIC2ItfX
j5MYSOcBzlRuhm0ousS6dy2+M4Fnx3WDCODnFIW889VLYJF4WccfRZg4X3BZgA1o
kW1nDjzoimj28aAXUPPaFoWCgav7RdruiKpdgriqQ6PuAyMq+l8+8auGo469fO0A
BIk1CYuzdj4vxxRbrHEpJ/RIE0iakmbS19o6+8IheGgGCs2axq0Wdrluy9ianXjC
cjKlpsi9amlm1Ppi/E6QfXUDMF2ClPLJuBXq04dBnlyr8jvOJwxRimR7+QHPmz0l
sTCOdEpZwDxOE8be857X2XuZuMDO57YgEt0yLttM+WcOYxa1wbWUo7n7f3653Gzh
M1TQuDclCktaPLyxYHg5i0P8iToMii9Zwq90MmJVRVGrH6QO4zex8peBaO3ljef5
HsRfSRMkxxfllhC2ndknqDHjB09PNh1oOlouuFXqBya0LebiFobRCgsAtb8EbIX4
3OqBZjnw1W7oyCkQxux9WkW+i+GeeZ3kR5uVIr1zBZDbfBQTsxMhNpx/rGWpIu49
gmd0sZsb+yfBpCKSAOY9ulzokWvB+vtzHA7e+fxQJjrwb6j30xr/g7VokxPPfudc
tfre+auBgTGeBYkbn/QJdmwPpNf97IG+TfmhpgNaRcgMva82geeleZ0g1bGukjox
vmJKfSwkgNq690fuUtK29EY7wTvcVvZ99EIZX23lsotWCgPT4L0bZP6ih4P4oC6+
EBnArUOJ+COpTLaw4Egy68G4R0tuR7SUOF17l83lzn4j/f2UGzUDdbh0J6g3Ag9l
VlX1TG3P/IQEPwnQ3uJ5vWKeG5XiudmCbRW3Zvaz/Muam1LZ4V712ATHKkpBr+Ti
JXtaUPHreIMC7Iy3chqNMfEHK9FPPlQhA9Ov7VJZSxgGN5glY7swP/7bjz9mLzgE
+auH9tPI2YpIyy7aFwJR2tJwEwWBoiYfA9B566yOj17p7nC4fpSRuulUhsgOnBWK
zUVaEonWIXzZuMB2a37Si0DEaHkMJjTKhYwO7fsG0cD1ZsYxo3wDXM5UBsieQcmz
ws/KT4yA5thMhHyAfCao3sa7WoO1CtqCJvGLWEw5zTtLRtcZGr34alK810MZ2Ph5
AwHKbjsxcPkR3Ai+8Xe0WANSccLmjd3frmg+f71IqtxvjgJdTBYoCFpLjPei+Y1K
qecS6YXP/FaOXdTOFT3HxrMgIcF15BOWBmoZcGv+VXf/tekIMt0Zzij+wo2deM9L
BhW8142bAr9+tE6jdCsguASFlyYmyjFY1fJoWtQpbrxPPc7d3RJp+FXKygRrcf7u
Pmez0AaeK6J/R27AbmCiGbv8A9g2cfm8XbhrpSoyjZNxVOTdj9vnO1tRfN1/LsE3
3Wa28g2oVsumQjnODtay/ggGvWCL6/ZZJzI5kKi84pSUR2B0mWvyMzVicpuCgVex
lJkm0flE1kUlI3TzOOyxc/idjpgrt2j4DVTNvYviaJoWp2Zi4VjknShzKCH7sphF
TJnXvoTLZ/EWu7sr+1INnRSS/zeVayDDl0jsNz4PEOJP7+ykpIOBQshSzqSJiPun
Wr7962wU+TZWUaImDTo5qA5Qcb+IbTzTZHNG4r86vIXDke8PTVlnmfNpkHPRVSPj
b19563wHpInYZizXzne+vrBgb57FKeZiMxV/Ged3CUfzmToJpWHMTJgvM9oGu64d
Tpa/kFRCN8JqqdZx2grPp5Jz64mofpfiCM6xM44C21J/KzDdVDV0d7tqtMrOWrpZ
1IcxVYAY+Y/vpun+4mwvneIfK1pLOa03P89xhOUADr3IntRnk5GCh2dw+ug7pmMq
CFIoYYUtiP4rFNeFPWfmWsPE1WmSkQow7ZAB3LRd94v67aIegGisAePINfReGuVl
jv62EDCvtbaTQgInmK+kbEH+aaN9a1aSHItmLvYVLZeVJxBe36k7RujXyJrDQmZa
RvUymm9OQ6n21fPVTPGMTradu11/igw1PeUgmLaMRV9Aec5eJPJOU8A9m1nsoLlu
LGe/34p23qm6ex6bOEeFmdE9O+pvKg8c/ixt6hRNOw0KQMgYlO8sq9SIorm2kY8x
xkRrcMuabjGbBmb0BtAjnuveWyvfwPo2tTazCUX3ilFyi5QqhlcGbhiWboJJAhgC
JCt1EWJR+sX9EnRMBM/rZp129vaA3QzFeVfLnfcrFjFXJI1TqqypsUSxNIddclLB
0VA6tqYElCHUM4N88d76J9731UVgYmAbD3KtCHuxAlEotcpOKEr0ZOj6IALxRVni
+4QT550CV6C7j7oZJsqiv8dGInX5EdnXoYzDRIewkNhanDN+AInHqwsnFBtgmK5V
Hza9Fyl9gDGVhttGzgxf+hstMfpRayJDlTt7aEiM60zjy1gKCQQkQTkRktegsjDv
R1UXf29Sawx40CnmYMpG6ln2hGD/L6W3d6lQqLXJHdSn4POlmUVXvgae9I2Rahsi
SGzD7GmOqPeHFrwfKizY3rLGyq3ZmLvaAYvBWBFLZAJ3+LfwbXXsVwrTW3y3ponW
3LiPJl1U6Vfk7pV0YgQT7f5LO71YrO4eMok94LdUmla3/GphTKTOt66QTiNgrzqT
bE/vVSS9Sw0ICYRfqGmgPrgUJuCIfX6KD6tB2tgGrpehnrbfDeAWnx4Oa0OIzBAA
f2T1ns8lp1SZuelL7t2dtvPcC2e38Alrop5G1emH4O9Z9opv4O+wg4uXsfoLxde8
UgaEBVnMX5RiXyEnMGoJ9whzSAUz0MQg3uEU4pVv3ItQSEvPMG/nbnOibCyfF6KJ
z/My8XWxzmL4T1UjQi665s1VMLkGt9uSmS0xM57vfyLh4mazKgN0RSipApQfT/Sj
NQUlCTslWdkfK7Rk8cpkTCL34lXN4RYsiJPApUwrKQv1PAhQvqyv9WZDbXewvXkd
7zwgO2aX/uDDygRf9y5XidW2mDhSfxuKDnoPtlATDddnaUcEfbC4liJfE0d7uTOR
urH/QbRcca1H01IVuxpuBrpz984EQ4d+glJxewhsrhZ/zVUxHhA2c+qenTHVky86
VD1V7ptHWP2AUEqWCKzhr85XCiq6WzsN6s8djjh/G+u4BMLQH0aEMvzoCCha+QdP
KFy6dpCE470MDh+iUEDg479JtRLp69jhNyHSjvPnFV29DlUqxMilYcx5kq4y/lOD
b/TFe1SeY5ZzKHhI4AXwofCkwTxUqJ6iKzGMm09VqcISE1rlwkP9nISdPuJzLF/A
tTECTISYDE5ZXMUBUjPJFhMvng9giUmOUXm+3b7D9KJNXxDp5oRRlie2SojVKQfd
n3m72GfB4smimHmgtuoy96RQzODSUBRndCVeINsmhvITgseZwtxWNO5jwZu6uiDg
s49ddNrBSraGTsJhOsjlYK2UO1DIvpvYxRLL8jU5BcHUzjy2fSsDMwaGsAV45dl3
kzQweexgFdpitsNla6mQWrVisTqpdgJUKPn3+oBZ0CVcyfL6Ud5mJnOUxR3S1qfk
45gn0D6R9l5uEosFBDflS9LfB+ZqBquxOcIZpFWr9PfT5serV6XpYyPCi2rXZqQp
226G/oa3rPSKd3SpdVPIzNHqrEUUehHxuy/4N2Ij9PoUMMScMjli6zl2lb15e823
tR3Cx/URvU8qnGdYRBowvMA2QDT3KmjA2TVXe3yZ635OiJnySSInwb16go5n/5vf
KFuQ0CRTJzIARQSvXsLT6VXq60GvHyPhqyMtgmRLYd5UHbsjo37Ompb+m7lsd2FV
QqGux9ewREVPNxAqOBCv/a07U3C4iRpbxGlQhZ8wPlyjzFjiN+pg0a7qVXJWkDaz
6XhG4DeDPYRys95MdfkomS69C52K5Uq18PwNLiG8IUmGx0SemeyTflG5qXFt4Ugz
6NlOVQgMnTRYsH07SwwVTcYULbbzpzY7zZg1dfkbig3GG38W0rqesy9Ow/EWccHn
T0PXheDugOc7rcg/VyohmgziAHjWKwkkD9KDka/CJk1TkMCFMXb6QcJzjEag2b18
IIXew5fBxCzdCnWE3EMJG1ZmIdd1gsr6swu8PEDAE0wP3FWx4Ec7mhrH1XtPk+8A
UT86Ftoj0ZOCY12b0Kk4fUzu/U4BtCqUbEvwvQRJaufP0tRXPtfsArz7pnYL7XGK
e/D3mASIPonmo8VQZNlyyggd+GftF8dbAWFyw01OEEowRAfW3gsGf1Pnh/b+0Jq2
ThGs51mw6ijIxDA0l/BwmRbKdfPYyM+6AD13Ua1Eq5PydeHBIuJcePKc8p0oTA89
gndcP0UWs1+RsPzxGjfXR0U6mmFpdJDnxXseU1D8xPv4+sFHwkzUzv7BOICh7gsB
M9o7WKleEc3k6ETjS8ILXHxzYfFsJGlPdyaQbjMPSCfOD6fyMVrYN1Jr73Y+n6L/
I4ITD/d6Jcvu7siJIqAU26d6WGXfBXuVXiWNiuVPtI/S8IzJ0wg+Z4R3ELg6rLBW
TB8OxJ/tEyKiETP1XJcqMVUexAalBfcEJsVrqbRKpaJkaDOieqcITKg7EfYsZ7fv
p9n49Vaw9rud7o2AvDRwqqPg6/1bLh6so1LOrBrGJOAGxi1zZ9NILf272pWpA7Vu
XXlHjHk8kgPs6RktRWxXLyWW0Wyft+oaUT1FVAsug/RUX4LK53HhzVXmyR81LaZL
TAgFplMjcivYspro1q53JjLLUT3ZeK2PWc/e4za4dXJSgMv5BWeN3HxURSqNQLI2
pcKGNZ1AM8n3d2Ai0ufMOqr3CWE6xT3FEDGhEyuPaksa+1MHtxuTPS3mTEkPMLRO
/gNGzk3YFoZn3XDzwUC1OKmoaSyUFN0M1HNkG5VZ5gnaXlIqynbJFc4keB8YvXCa
kA10PTIwMLCX6EsWXTASzsZGESGkw2XZqq7piXvRXVoqlYfTEh/eTqsc3zErIyeE
4o8RmV44GwoTQ0/fnEgPmc5cTQ0widIWXZ1HW2FrCr9sQZ/sNlcu09OBZvSLef4D
mLky795VlIDIi6HMO4Oou4bHEGWQPYsyfWMdQyydBI0W/xUWxvs06emOzPBkjo2C
MZ/CYPKknWHnbyPOm62DmvkfrSZ/UyLeICa6/N74+R7zUDlYssx4kLul3ZGrzzDX
Xquo2YPDetcSaXBPM1+9SejUUcm0f6mRd3pzwIgsgULLzU2xVqFGTiy8OEfz8eu/
36f/Xb9v5ytpaocOJUZ0XSKKym2PCOdxBghH8ZMqZUFb14nW5maSbZxY+85bEde6
0J3XGx0Ekf/KI2FrjdVhZnU6gcrk2w91zqtCYiSmlqbzdwQZj9gG9ADp4HjTY3mX
4ijBSC8rIxaMBz/BP9SeI/gOs2wGrzSVtVrm/k9iMHu8f7m/rVAcyJRVJHbz/2Jj
nVAEczGLGmdAiaFGodwYXWHW9dc47dqFhggg9xWyqbCmelpIZjPVuBxWBQ294+oY
78hfeYQEkQKzlRIgz5KRZKKCkzn7lzz3nvuNv4kl4ng2ak/jpMn446RvIHeMTeMP
sH016i+msho7XB4OPiyO9vgInipT7UVYWDIKJ4l/bJ6YrltRyXrU42qEHXGFxdai
HKVePOe4XUorI5jofVknO0Ox5SGMO1JbTmIPXoyJuAm50p6RQAKqg0kffF9n7PCt
8IxYOvGAIi00CCV+amwoXLr2yMNtLesItpjztsdS2JO97pXcOZdOQkB0s3dOIB+T
5QtbxFacXwVnSpm7Fb8U4cgvyxoUooGzMVKK21QQrYyNLXYv2Mh9QOTiVB9k6xtD
ny06tOySbbVIMoNlvFS5iulHo1tt2NzgB59c0bmqSFhUWNvq+D6hWrFwa1VQXHLJ
j6hfXpaQq7OW4Kc5fPoWjkErHu+SlGV6rvSluKVspRuDQvmClFMbzZyLAXYUInfG
moU+bz9en1znMK8RhXKT0fB0BJPqll5MWXU9+hAUwn31jTBxtn8Pkb4xF4fjpvfc
R9J6BFCEAHdV4SNCkkdJ3+4ByFvrat29+av4x7LBjgRhEaF9mYC8yl5HRL6TpuhY
yyorgZSqhlK7V1Nalq8rJ9SZaub42JXOHjezBVkWGfrZHWdaLl4nnjN4n67GZ6SB
SN2jZhV8L8yftKj10n5KRLoHJMs2OhSAeeJWSRR0xQCpFZL2nTH8nc8P818Tz4Db
4JjXVlMqLMyWXpxDLMqwuiscZW/7fbcNUjLBl1nl/3Id6iPRSuj4fR14hpWi3apu
7cIvEXpQYlvhU7NNgghOmM5qE7qr3wlDf7K2zy0a4PkIEHT594aspiqW/d3HD58c
+91equ1yg/nOLrStL9u62riUs8zuNNsNKlDCfhR+Twr7Veq622+hNXNdHLy8XvLG
AS4aOLAR2logV5G6zxd0YGY/y65mKmzPjU+zTk49K4tQ+t8zV89g5+lhfNLHtI9d
qoWLdhRwc8Nka9atOfZS8eOnGLp33csEafxG0+DHIqtCVSi4I8fKBGztuTGAKo+B
7cw0abFSDyNBKxEfUgmab/V4eHnou4OgiijFwXDcgQqxPTIq8DZTYA5RqDTuXppK
hPK2WGCWdpKpbzxmsT4fUQ2lEE2hjGYcQEaBVHu3vEAGeSzo9UZ4pJ5oATcswRnr
Lp/UMjJzXgy65ncBtEex/m/foH5Vy9HPHua9xcpSJv49MgerXpC2nokBriTphTJq
BfoK43K0n+AdJL20JsqAnodc8V1REPWtHyf+9EGu20/6kWFWkRQoxcCk4uqp0iI8
5NPSrr7og2gfDA+dA/bydOJo88icKf3XSXg0nfi5pqzTEkBFutng7DkO0op50qzf
rAKsJOcnSTueNJL51IFgrXZXRphePinLuID7V8ENT6yTrEKBkwAgS/Q1nQ5TVuFP
Y+h+wGClbM4oc6N29qpp+u9ZKa+trdfTKwEFV6Mkn3tel92oxnS88uNKENOAR3MI
GK3f8sU1/GINSEN3igH+Jfe2Jb2gSwZQUEybhpQ0JWzK/Ltbdis1RuUftfTjsmzY
ymR8zq7OedMxO4PLxA04yFBHkjQbYk8lak2uiZY95cu/KVt4Os2EAXCRwk4eMaAb
5uQ3S9isr1w2x5Dt2UuNzyAmmtiEby+ZWS0e3f8e6H8t6WG+tU9aN+c840AViD9P
XUwgn/wFOCHjGhXajH+zdIj//TCZ7i8gSOWvmRuw732BRuCjB03fkJn/BnY1tCW8
9NBR8Wax0pIIzXjHRlXyAU6nhXY1Ofo6sOWxPcC6Etp08HPJDzFCDQq8Zp9Q+1Y8
YhfOfuKMT6c1Pv58vR9C8UutavS0yUhp3kDf/8Nq6NNanXqrZSLdwT47NKYElWY/
yPGyYw0WbVFGspIO3QDB/evD0JqScLbm8+ZCHXuG3x0=
`protect END_PROTECTED
