`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J+EtZK6hG5h0AP/CkNcc+TiVe/4vRCz+3TmuHWMNDhRGee2LKBFwrT/ovMUVIwpa
OdzE6L4d3ZVDRSL5tuPmz67JT2KWwUZ1FdBdPpehEme4MFi0kZqABTv6WPXaiAj7
M6YWoqR4hxH3BuyMV3gg+L2iu8lCMEqRk6wOncN+rvwI8gCjtWij4So8vsIes57M
NidgZ8dw2vVXZjW2feMXt5Z1oqV/imvZ5fZ2f8QV5bcJD2SXZwxmU8gD+DpVkcb8
z0b09Mkpt3zktQYEdj/bOt9KhRYPI0rXe9NKxm1CRHnAGeYtVcyXnSpQMdOjbRNV
DqKFOyNYh8+WZDnmPX1wD4AFaoNVgKNK/0e+ATwwEQbc7n1a5+5zWwn4VLjUUsDb
3+BGZWgVJvADw6XALy/APWTJi3KVf7A45CHiBfBilUhVRLjU0A+czGP9YqB1DYBQ
lmDeUXjg23TfhK/CM0tqIoW4/AEihUPK5OAN1vU8zxkWDQiK7qSmjK3AfV1fDdld
+1QtPAW4D/tO/JW3YusrEdNVN5vYOw4J9WWRJSyTNkcQ7BexHS8haMaL7vN67wbb
Ic3Y0YjiiCr6hyEY1q2SWQPOhTngpmhU1xQCcqZsMc3BrxbYorjP7r0PxiBBvbzn
QfvXyeSYyHei4XFEbJFXVP5Os/2/RPxAjRh0qRaBEv3cObtaXwC0g9NiT6GnYZtf
`protect END_PROTECTED
