`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6JaQdyvFgXbj6OK/IkCmUH50EwdRfbWzdbAoKrUZJh45puu4etTxr0kAL1PEEORS
UKe6Fj26aIkPP5yvQtOSQQIBK+kMDineWb44EH73mdwQf9SE2Fvn2t3oZh5aLe5p
5GCkFUPy8o7g+ZLpObFlV1tgNmxgFBFj4lL558sCtQmprQLulTw+cWHOrIA5S6n/
Wgl4aBE6ed765Qu68ub6Q6+4c8BjW2Q0z3gsJWC7FwuXzmQ/Hln0CKnfwG5k1sgt
bXXg63jn17P/uuhek/tEuh2p9iYxEDoTjP1OTwpIj5Cotl0dCHloFwS0iK/OJpi3
mEdv5ydpNPxoJbpZ5u0/dGfHrWS2fojLiE+Newd+p7/baI3jJH1BZwc2fYKbQ8jY
8jAb78gMdi/Hkw/74vq3kOGCd5lCO/jCnalHEgmBA1lTHuqBNUYDaBqrJrPF/abM
GzsZwfS9S218fEvGa8awOl9alhbw6xkGx1Tovj+Eowf0fNEXn5AmcgnMf/hBJFjb
B2mE0d4oPyEuvoNXlhK7WvgXSEYgR6FeYw++HT0X1EoGl4HyGHvyN9KKgmWwXnzL
ubv6XYVuY5PWfAMJbF8EfQ==
`protect END_PROTECTED
