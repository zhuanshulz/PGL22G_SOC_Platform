`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g8FD76JiXcEkypoUbxkMaMK+TLB+HCzZW5V7f6VQSZMMV5tRujojfuNxM4QXDIiX
69Xdfn6di7YDxdPs5gmmG1LYBzy3zG20qLu/Y9eO24ArZ/lSG65JVnjm/YtwhCSa
7v8hX6b1Jji3sWFMiJUH1ZuohnEOJFRnlrN3BaKUXODU55nf2wQrZ10gCaAP2C+o
BE9eEfFJ91mG7t2LZA3oZvrpGErvBaYQrLTlfvCKkSXTE9JVffaHyq+4W0rrFN7Q
mrMr9LbkRdwOxwOaU3K5MNbftiyKZ+XtdgIdbM9HZsIqSmkXV8cGcijPVFtWsgUU
E9m5RXmeAmCTwgGWcnsqAQAQ7K9i6LekiNGgxz+9+KCMJyRBsuCgQEQDsPRmHToS
GJsoROGanVo7bmmtb5cKuZ+ZjEOsULiHdL/HUuuSkksLKC/P9DHCy1bY07jS1m9L
xyHSoE3QkYlq+M3VUZdx2alSwX5jMdwHtOpdSSRhvndViImThdTWsTXMtP1ofaMq
4dDg61cKVXwKgI95qOn0bul3ZAa+yYpBUWMJ/eyC9UvIcVUhTuQJPW0Kn4nIkiMs
/gD81jx0OYGO+YwBi+yxNPoQNpQDruHZOLL6JRlGzqCOGDPgeNSACF1ty1BcTyuK
/akRD+Ln6sW++1nu1IIzA+0JdxpJRYBYDhqJOmI5fGcVs7mb6BUHpF13BghZICsr
yfZBSjssQ/iNB7hhYxD5ciDcSlSW9GWvbizCINgSjQlD4Eh7VSWp6aExPNvSs3Wi
ezWYnvvE6eufrofCze/f234bTO1zn/Ow0O+d4te3sRxsQ+J2wMydQISICn3XW5Ce
hKbtzex751M9o35/zuipZstDvFnR2EYBEy6VYX0IA0RYDLwuvH1zxomzZCZA5UDh
uXyXsH5JiUBy1/WdZbt8vcs3KvwpR0si8052KFz1a8U1sNGcn5OEmolY3ZZdhfhU
4V9h8bGVF+m3B5rDXO9nk6rEE4i4zc+lgeRG4W0TJ3N6puH6M4mj2HfqGKWA3H3D
8zTbu519Ly+JBx8uOEvlMuxcgbI145t1J9Hp9kE2CSASN8Mv56cTs+xMAU2GoFAh
XMmA8HSQWDGDhEfWfTQghW0ziujWRNdcJ/H08wVMUh8BzDtOCFW/vDnkF9A/HVsS
0lDAnfTn8ugjAfozpAySKdB/57tWitI5zrdVPV77fCsf3CIWLMwtBwbRzUn9yMbN
lLaubwZhW+vZMn9f43d5SN3mQCv+n6STCMSZIA+zLqFs1jB/kav7lRYSsGn4uvt+
OUzklCkKGQ2cfyRLDmqg4QE7JdChpMITqed+uwKYPJIc7ZfBysWdZTjDFCvupBTp
3HZQTpC7+vvETFjs+GcjQCS3KsyGFc5YtLNbVmxcktk0cUzTUICM/3Se3n/o/2sy
fFITdKz52oKyTQQuZGtUDPtlllEk1PdljtAyp0hjt1GRA4e75S/s9D9k804F1Bsv
YOx+Qg1LMWGSAzHCXwlwc++mKihXaGlize3FkCHA/TEbH8a5iCV5yCjYhLzc8btC
lG/IHpcR7GaWycjyq5zRmQyuMzAxAob3GnYxLtP8Os50dl7kmbWbwUpt0PSmoLzW
iTeH8I37z+0odMwlQv+0+hrjQgmiYRwZ5niohSGNkYGfE9qkbJ3HIBzAy2HPARwV
YaXO6YLFuDCBjr5XoDkhChMsUXlNazY3WnWigS1NsELqVxue+SL9+vMk77ikCArE
ZcICDCSLgZdvbPLtUGAUa76eEMAuqqkFA6QBmn3Ql4hXBJoXXJIF3+TyBnGkfq/H
zVAHX2xyB6WNWATf6ipfcdDj1afvWEkf1UO9WSCod/gUo+711z2imFTL8NQjDuCy
vjzmRGt5wt0ABr4u/4n06Gypm4QE+65JHCdRBF2AqZT9j1wI0SgPdrwL2xcMv91Q
o1psB9y6ZnZpUKT2RvAI1J9BLBqNpRyQD/lTBIKhZgi5HuL0HlC1ZhQi+qCh1Rf1
u9XYQEe+wirvrFq+U1D14vuE7DJ0g8h011O5Mys8zt4t9NkbpOR/Pw6HmE9w8fxT
2lrGLl62U09ho2m0V8znJJs9SaE0Jq1txHNoy89VvR3Vz2Jlj02bA+ca7q4PtZr4
xPPlRojnm9i8jqektUK8MqWsLE7qFcDAjQEifFPBDA1AQx/AUPZaRnDHlamWZVtV
eDCvjWc2Vaf2qrSe19J3oonMX51NbXsMl7FAyyxPBe6uiQ6Cx8jlYJ/2lC0ECCFt
hvTOJHQs7amUFPfbrg/y36o5xCxk7TNYLOc8xhH3FV6aVUrLzBzdvhAXTLiphflC
4aa1UiPdJqtwN6oXwHyhmLqoQNCXDp5VVsycNkEFC6KIXz4nzxewrvgUjaP7LYQn
jJoNOBhIlvE/SKnGCFWJJutlU8eFuCFaOMRYajJ6dwid7txE5KoUZ1qA1SZT86g+
2gUEFSu4SB1B5B1yFHql/xDc4eND11MGC1/O+Clx0LSaOXwasbRf49Ao5X44Rc9w
OTmPOElb6Gazg2js5+Kag3e7mQISWu1L4st9Ufu/22Q/ddm79nbHQbl5fADUSvx2
1jgJf1q4Y1lcdxToE3NZJXpbOverpznyby7+5B/+n7ibP4OW8XHMAImoTdI7PEjJ
d7REfT3Sb0rYd+0M2igvdwA1WmOzQ2WNFcicBxbboWo2ZfTANz6u1tkTslWto4UT
kC1g6biUSIa/ChN3W7gOUeaYkYtJoWGG7s6Qp26UhIH37LFPuiyZ885wh/ZL6wO+
gGW0fSUYm2wIrSJkuIQUGgYI622E6PyvV6YgS3cBawucm/6kMMZfT1uFaZJA1qv0
jHgqEZmr7wBLfssTMTZTDpsFp+vuHFnLp4C7oZ5Ab5VrLa/yi4YVkMLWrh7TxbNW
ckFG7ImbYjKt++2vIMoRnlMOrYLt1JVYeWt7Ij0Ih3zGKVvgq/ghMjqMlvwP11JV
rp0f/MguQ2UgAldjhA8iXScnHxMzClW9KDVM9h/gxaj09JFyRO8aiS2KxrN9wycc
V5yZJGKpTeazELE8zi5EfzTLEpmCLhJe5/XSIL30TzHXP9guQr43neC4kGt1//n4
HD9A7ggGq6uLB1Td19g+fZ1E47v9Lype8Toh+zPu1G662OkMh7EWxyZKTdZJPxBK
nE1fQbjUEdMExCr2Qwdxgb46wYJYBCcgltLBS4G+dc9Qsj1Kpqth/7wCTL04rZsA
KfwOgDhtGNenayfEYdZguVyJB7LXiKHMFqAmvCxiDCN9QWlAOXxTYHY48OPjcgUK
J4li0dxrsG1sGmGjDVOmUgpBlDeCAquivFSn/wX72VuSNFZ3gdIZbjJOs5kutDIZ
RCl2MrNVgksvbkjTkMerS6yKbc3ZmEMUVQn/T3AedNIWhe4JEWRjPviG8T0+WFwH
OzExdDh+tm3KA9CTUi7LK6upeyTasLbfi4TsbYZAiAQ=
`protect END_PROTECTED
