`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yWLijgONCI993vzEzNNxdfKHWgPQWipZDi73yDlcKSnCNNTASJhNxeCsW3M/11JK
uNadnBQxuYVrFge82nCOfZw0zsEP+2R4dj3yfhyqyNorz0i9rtAIcLFSk5vygZI3
7fN7jDJSe1U2qIv0fdQAUjp+BVkjGJXqzwQxGyjVyTz2WOfeZ10wdzRGiBsf8/v1
LoPsgTTql1uM1UVnopQjWoUzG8Ixro17kXSuLenJD3kwC1UpIahlXCiJPO4Nk1OT
dvIt4fHCUp+OOV5/JjB0521IAbNnsWvkZHlFQwcQpI3tpiprl2aq5CP6NazjNKI5
eFZ0+HcIcuP6sGR3zCjsre9A9h+Uze3HPZmOfC8CpbDp9RpX1FcU64AKdXMGDIRh
Tc4qEkR/ufdKTekmNmkUQQ==
`protect END_PROTECTED
