`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GcwP0f5v9QcOuXA2z8ymR8xgUCyMyTHZD6QNWlgBnzQTKjqvhPdGWaYWhUdt/Nmh
8L6sjv5yVz0Tdtiu5cqwD/ET+pVEhzoSYSzOyUbvu2X7kBIZ0dW7kehg1m/FkGXj
UiL34ZpnaAYTPJr0RjlQM15A/no0kqMX4i7emiA3IRyy7CRM2ipKQygj+FfsRt1z
iyjE+cYSJAFXyF7AOuzFgS3e4022in3CZzWtBW3MD8FiOrKbUMdcJb+/oa6a/8sY
f8vr35d6CZg7HB2hgyxfh4GOmP0bl2mQsV9PaeeUdL0yGV4jRwwhqh2Dgpb/Mz10
W3M5Q9A9WYS4KaNFEv1L74M/fxghgijYSZf0FVOYmuLoemQrNLHSMw0TagVQuPpm
GDXjJzNRj0ef409h24IuQ9zMFm3xmwt65PKhROi/5LqUU/pn2cTH+VPsyzzlUGZN
qxSTsTXh2mAp2z/ECo6/LTiU6kfvVO8MAIbgTcztUJ2u+wcntQJlXIm6KgJWACGT
V40AvPmsVCYYppJ3iNIliYRtqyItK9fHhZ7N7nkzZozAuARaO94JKT+PocD8ANT+
TpCcYqy4Pq90nRdSpNKDvDvVYAyAueegQM9Nyrxs6xraPFtmJswth/rV+de3nCb1
+Gs66T01W/SnpIyWjN1NjJTe3FSbqT1JmlIg4Z8/Pu88zrgWPSdcgW7FtMbo+TQv
VywG7cXGLO6TNZ8DswhIVrNvF72HeEY726wjNR9Rf9KxAWgdupjfhfCOmfc67Ufy
9vO6FA/bE7P0y3YJg2B11wP2PysK3DgezxviqX6KHPXl/IA5/seK8Ajv/VvtHGfA
S8tmr39eSu0Ih0JZJIVQ0wm+hod7BxO3cFn0eDCzqeWiwIDTskntSXdMQFZTh6w8
GcFEvIDeq4Djl5HTENR41/aVhWsgQRv5ORCHUyAunEMlw8Xd3qhIu3TPhPb35UOH
4mgQ0nqGZMMji/Bxx/lJaqZ0+dOP5m3V+pnUhIP6LlvruL4HPUHwzXfK+fexejie
9mY28fxlPg6x65KpL6Lg84ynfuge8Z0Cj0pu4jv8GWEQHUqln7rV9AGUYLeFFk/J
0+DfObZ9MZoCysOUvbVj6j5f+MFfxCH9F11EWWsynNdMv1Kx1IjM8C9IKM2OONBS
HeII6JMDGcHPyP4uz/IQ/c4/b9WlqRiTRd0FTelUYozjSBf5GhCbHiy/KmX9Fuxe
c12Dd9b+KaRg/+G7TXS2KXXDpT1vxj/PGIBIpFmeYHrCw/6EXoyw1/KkMf/hq/Yn
hwIkRknF+GEKmZ43dloDXepmnzmglSsZ/4UaatQTJL2yfbw0Php2HQ9H4ksl2En2
WQ6KEHjtAi0LOw3V8cAhx2weBp5rutUMc9of2svVt9OqOL9qo1dRMiXxfUsS64IB
VoJqTtMhMRdtaRBEjZjHooZ8fjqzoXx0sRH1Banwpp++edLRrkXleZrmR11UXozl
BAm92Q+0giKE7JQp4X23b/EP4xDAycWIM3H1q5c0YSXL6diN93QkSgzORgmGWKlu
5xTy39vYcqhg3PUcGFUdYI880q7hV5X8GuTOgbMg9ioVJ1tksD/nheYmNRr6/DSd
79GlN1MNxyLr3Iqd45NB92rM7UnDKVASlkESSLbmT2yMC/513NApsBmPJ8xuR06j
H/Pl4Ai7ZaktVUfIprlewm6mOXKRnsZS0pKjPteuyc+WqXad+3Pk8J5NVcsRJOIq
Rswp91xXOpLrlnsOLzQ86lCFAESh57usJZyoSXp8QhgZObFAEu27nLWCf29BIdBD
nELt/NUquP0sIAKxrKxLYQR68ZMUVR55De3+PIu/2dAw6J8a72f81DhvO/8T+ras
MzD9D4Y2JA2f7HaBimWrZvVeeeOTjEhQwV4oox9AbutMl1HrMWGZGo6BDFuq++1n
BGEGiMIgbCdb6611wwaoVWly0ukCZyrglbMTozWFtgm43PYYDcUhDNBQc7HMieBW
KSTjZAU3PjFng6nEhHvkSxIZH4NOBMe0qIcd9e82RmMoVOjV1GVn0/EwKQFgOIic
k7Lii7i7n03EL72vYAfFvL08Aczzp+I11mC9pWI3AHFg3ejzOxOgY+7MlAYmZWcq
FYPBXhBnjBP1ofUkqj02rzcSnxa0Th/7il4mHiquFr4Lc73o2/zQbXF9JfUzxVCv
wo7OIc5patFnIDj1MTp7b+Ic6SveKSgH4+idHzjL6Rc0jfxnPtj7aHwkn67S0Ccp
o3CM9VwbWJ3NikV+dZYxT8OFg0rNPnCk98l+4pRpPyBjD3ee5j4K5OpZMN+rDzYv
HiiZMaVOWKSupBnlP9lPp8rY2T0YUbJGp5YovLfr4cyEbs95wFuVwE6cNfOCUSyx
dCMeeYAIB8kBcNluVUI9q57H6BXiN24IdkzEJx4vktSErB4g4yvzoWxsWf8MO42z
WVv8fqeMxRg3gN2wrWU4Bia0Z1hCEZ3qTTe2dR/uUJSxZIgiKRDQeSNcqaIh8ZIk
cJR9CxbcbM5XpOEi1K8Q/eC8JB1BdSMYB5mLHbDoqqOsSEi9UC8HVif/Et5AwMHC
4cpHYuqaDPPchSIGepVMedyI4tG6eNZRS8lKFJi1PFVAeg6pkYBnLgDHnUgURwoz
6T1qeQr/8ebkhejIEpcLL/R7CyD9CzAYsYVkfRmwxI+QrQ/G0wYfI8+83/ICAS5u
/4ukabm6o+ZJKs44KqshfbLeCUSFMY8NbOp33MQOdQKdQCwP1m4J6bLM/OHs1pHS
ByenPsHfHurNmBb3NZl+AXDxBi2qyQKyuvColCRMjbRs9t9p8B7cfNP1CfTSlNX0
0ZONirM8AEFmbebWa/JU3K3q3okJHUU/HYDpR7PJ9sC2Pw2qXw23T65gNXXP4cdm
Z/mUhryp3ghIl79+LdKItaJ0otaXg93p6BojYqF/Dj0uKYTBtAsCTAshL2DJWbjU
qeHQlpK7H74d0m+iI8dytmQ40CKBMHOXsTXnnOitleMC/gh4syDODD/MtZQ9ugEK
prKb8YkOmXW6ZiQoG8nSg0517j670QZZ/2gtLDbCMwhxXSst10ivPGdD7J0F/aaI
7sD2BA5TA2/j93saHx55/3vWfEZC2RSkhce1YqQVNNNDUh/A6g09lgo3JY+YKro9
+6N77OMkFm3vI+x3NqHiUy33Rb1dnnFr00Xv6s2DbjPHA4w0055atupBr+owE7Gh
ZPBd7+fkWXy9ynxDB21CGmFey4jarxSTKvRin0wwe1Bk2Qn7boygq0oraL/SusN0
fu2olDx+XBWO4Pe3dZJFEW2s9O3OsrFlhiRvc9hFSOujRhUKp0NAOqo3Uo+NNHw8
JMrFGK0DbMuF+mZipbZrlTSZYHmp4kyhHeT/AOFW9DSSP9TvpE94dW5hxxr9MfyQ
jHqYZ3yxdYujx+M1VeF75kD2Qz/3m2WYiC4Va30DF04+oemnzi9sF1qxNRzEhIvx
AqiObo3J0Gt/9jwJyCytCLBpK6LAJRxKwabQHYmdEiAaW7FJ4RSaYqvfpj4MAF/0
AzmA7hPt8V6yEtb78478HpveJ6v6FwULrPyNqpfRZP4RQiHGIQag/KQN8MAd+tcw
KpvAzY8aNIYXuCUVNh5mjVi6fVQqC4CvznONONXJ3dd0YJvdva0d+/o0QtLHhlfh
6/i5qf138d3NWeH+hOnVY49FLlDnvEwK1/aC6ah99fg7+aYd0UXlRpX7GS+nHyAr
buPBO000IAHz4DGeFw+TQlG8sNFsX4QDjiUkmOLUzCXT20bhbSva+KtsDQBW89p5
R5gnTORAF8gsjtSNU2R9Ir8pagiUAa8Na99wBbF6+6aKpc1E26rRwacHrNcwNNjy
WL+U3qyiOj4PaD0+lUXkZJ6B1+XTj3P4SdXee6mnlzlFglkUgnhiUL//zRw+VQ0z
DPgmydpeloTgYNtcq1+HQx1TVr6SJ37oI8m8b5i0bui/Jt5PzuKllqQb5KDKR07o
JIjD8bq+dsTt1r3m+uQ6dh40GWBqgg2aysoGp2PPpBQ7WDo8vNNkZxhHre3mYrdW
qjQcdbwNVMg6+aab9taKBnyTABwFtD97qTkeNr5EJ2z3FkQsk0fqffpxedXXEDnS
f3sTvXB48cpfB99d4hwL8ZfoZj1Ci9Qoy+nEQbBa0NEtaImzpazgw4LsWkZgGADQ
IeyTcWI9fBSRXhlHrrNfc1ll3cu5UDDu8w3bnOTYIdliU/9u3Zmy6KXoaaAxzgpR
pUctHlNTnz/bTV25S4T78tBh6Soerc9nubH7MBzZPrOGU672qeTMYkqz5SjBHXk7
+fmFUOk+S9J0BJnBwAHVksNCmomSBeKeQEp/bThKCTtf9Q6gI7JJbWyx95xjksL9
kWOPg7UUXvzRVxU1L3VVASJxsds51A6XOzBg/lzdtwUN+lzyA5s4fzFpH24CRPfq
kLQ1625h5Y3JmP/dLKBn3uO5hg6NV/08c2afrOj59I36nKd7AD+Z83jv0OqDfVhi
rRejpI9eczgGoIzMw/gjF/JdZyrcCenxroNRrS8fUCMzY0lisFQ64U1zXzXtdRk2
nndkSYLLPvDk2ffg2s4ZD53ewlOdDRZFZZxlzrDOPr41GHi+lmc3vUIUGgS8GXln
DU0J7AvI5MEtEF6G1D0MoQzkpNj3XRpvdoLYJN2iTQPXMdQe0zUtjStkBUZaAlbd
Yt8ToyknidlyrI6o+BHrCiuSF9BQAqRobSdfCfJP9ZrVy7JIbK2HSYrCxaohBwek
BGxhEz65JypI7JOmUgv/vVTGd4JQBB9/Zzou8veivzvPBXpoCBEZDe7ZzMOCseZw
dXup8+j/SzjW8qHiWc09S6EidAE3N0sIvMEg3ZfwR1tjIeZ5NOT5ZBqdxAci8EJA
THCCY6+RzKdcS7TfdYdpUsh+LG6ZkPza79wzv6zZyD6sTqPQf5jLo4c2qi4jBkL9
8gxe6VkTrMeNWjZ3yBg8vPO+NkuvDlNGVDJ5sTs3FCChgGTpnNs+L50KImUNjhNB
KjQicZjPTb+dmkcUK3YrQosBBUmhYe2zOhP7CuR6XjOzTp7E7P7rxmy+aaC0uIjh
EBjUdmM6PlQwOfPgxjEcvRRHYgsuC9AxRJ/mxFb/cVVlzav+9MUoXOgim8rz3b0Y
Jh/wWmJjsZdlagOmz1v+LsCdwewbA5d9d0gRl5fZFC58s4efI5OKpp4+Igbbw876
DKIjKs+7KWDgH0Q/QI1HrwKVq8i6eoM2FuIrtUqoaLsY60b8OGJeJiSC6411WiTD
df+YSJiMb7mzSjoUFHS9XNOdt7JHcnfxWyTy+ciyFRUFJIs8h14styVL8ph5UvvM
5woSku+9uusLFa2xiPgE9GMbj1440qhQ4wF33r6xaegYGSebTUaqEA/jEfuJvBta
oyOj5icK6SMEMqRQjJRviUpvs0YBB2F9PDl2F/6f3Ug2U6OOgf9+vsPfckTXM4Cr
eNyPzIXJFMuBt4Zn9q3oHGHe0x7QKnM4IJy24TSBi5Fy4lL/PfknmoPVo9+QnJfW
9G2fyUotCSm3gWfXbtrfhRwTbbby8SjsXgqV0JfXlMyOi/yy9sgKw6Va0/XBK/tz
YYpXi8RHYhAP98h92D4KCeC0QJEg/EFa4FlxKqCcTR3MbkFk3uaNXj5/nYysqc0I
DQFT/PfBF8jeaCmhAQhURNXZ6LF57zCLsrRkLQUIBpLyHRHhalys9M7MbqheDTx4
6bveo+eTASdWY7IkHlQrPK0P11Oc0o8ELeIkQsYO244xsYpStYkVPi83VKoRNNU8
y+jYrUO6RYdOuD4OV83JYCMDYFUTVBbkOQ9v5UhjCiJhIpd+N/PHNtWNVPaMQMsl
INAJfrNuK6az0YlIFNpYnAHQajPuNvgHeXPr4bsy383omyPqcvfM15swnzidTEGb
Ay4STM/5na8hD4uG/dHPDXzbOkBwaUFugkV/Fhv8OYuaR4np+fyd9U6M0b+jxi3F
LVwcnDXT6/jgyadq9akwmsJc6zMN4/azwrpZmXW/FLN2cNncm4Xr10PHIiEl+8wI
snRK6eDc8S1Uu3D7KA14+K61hvn4Fwm25fVOw9siFSVz5EHyrumijyR9zttume6X
uf31br6kYwkZg4jZvil4sR0hnbTFBS2RlRoju+B5zqvGII9+dal5gXEUXRow3SQ1
`protect END_PROTECTED
