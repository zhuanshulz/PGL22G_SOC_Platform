`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
guOnzGHg/HPF17tNPCFWQtXqYRf3ZI6DzBwqeKrwZzfxhpyzw+ECQHoStrmTVRPJ
KQkZ5NqFVIioZ3kbADgpCXmhiNM6XtxZtUDJ9IsO7AYn7rNA+bXLsA2A3+bJyA4y
6PtV2tFMa6ji7hwrQctw/J6bJ4y14iiTkiUU/glN9LEO41Z0N4LvNFEt2UUPtIzh
9ExCxlsOBBgynLSA0ALlvF7yqEGdx4ASwHFxsNVBzMhfw+dI4T1t6wDtK6XczCZk
H8B2lo8m9JsxFnXXsgrfP6Tl31diOIdkwd8SbQdjwns1VjE5wSKWmwhtumBKAO2d
t3rfY4CqylNupK59Qc1zBfxTb0CAp3yBfdyAJZLJKwr3DpyDQys9uVj36fZob/b/
EoMnaUI35T8aVybtbs1HmVYls908hvFRvQpJx6omYZ0X+iox1Zbqi6OmO+ryCVL/
HYYsUE9yINJyn55XESJHFhhB+Kepf/UX4YF9HSVnJ9x3rGHyQTEGStGZYUxel2uU
3Sr+w6U+N6n9thpBg7SlRq6v7un2RUMUCmyYOBw7KxmNf4z7kgvccpUXTrdj2dEe
`protect END_PROTECTED
