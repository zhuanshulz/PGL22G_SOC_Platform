`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eSV5/oO1cCM8xsf0jeVr5T0OXTQ2NZsdenRQq7un2jPYgFnmynHLSkAet5cofAMf
CEa2MgxQG6vvaZS0qmBo7Z2BaaNX1PJdA2Yhq1fsHPsMveAwsctH1858RgGmIW4Q
lnGJbGhXibpsb03jmU3/rvCcc6wUroOJwBZHCsFmqJDoMZn7u5+2QxXni6xKATqz
nh/rn8jPzAjn72SAe57r0vUNh5ldzK0LX62RAY237msJiW/ftzH42a9qLuc6HR45
1L+MoqlNCOmtcCxzdUq4BcH0f4/iOii3t+e71ncyeuUXpyaelEyfccDzWtgHTMGE
w/oUHudghrKwqGS0Qfir4SdZ3iG2CwdoqJ8TU/WgvrRMIuIWjDuAv18KrWKf04sZ
szQLxzeP+iCw15Thh+NRwaxV9rtgHfUt/1xWXmialAImBaPoqR7/4c3HheN641R5
G1X6aSAM96lwC00bZC6ictgn5aJDbVVrFCk0MjdLKGA4RheuaYMjeJGt+pmTFEM4
PT2yO+u89WEEciRp6QW9wg==
`protect END_PROTECTED
