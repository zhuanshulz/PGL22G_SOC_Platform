`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jc91p34u8Jm7L/N69HeHUqNi8TxBQfbwpy/1Xm/Co+2HUI3fQJiGtdB+j6iThkmW
M5hX4DGjzbzsEJgF8VsQFd2mHEvGTX/z8fuNRNn+nT/b11rBtRwzqg1e1lh4n2Mm
ibXxP2jt8+X4yGDJA8JmG5vsX1HNl4C8BrlQ62HU/aMXyLKh8Nd9zQJdKqzh2rE0
PuH22Sh6W2iMlu5ks7d3olOrVmP3V1zdbBW5KGIfRQYujko5miPt1YwxGGMT9/TA
TaCCkKsd/0Bu0pRXZt3NCBIGCtS/btNvKJIlKsJtJAohUmqvs5MaKdFIU1Eg4JuW
bKz/v+35mYAxONHHLEuvRdhJr9XjElgXzNGjKjiXUBY5DxPwZtJVK33qGjIaU/vF
zMDksjdv9P6IU9lwZdRKzPutsKJ0yFIwu13piX1zC8qBxlBLSnCaR0KIMbxPL195
5h6FttuyNt/67o6VKgVHg4JKeXdM2RRpPgSVkOUs4nCEldb0GHEoYOSHEWy9KTQ8
u08SyMClA5RUKWhftyCbYD+GhrQVbCePAChQ2grGbyHvE5eCxvVyEjgh4ZH866+Q
duxRC1DuFbzlOZUouywNu9mkiYXOFhiqsp3/U6o1334IWGgRrYHUCVQu1RS6yZH0
5xDGSCTkIAvt7wlY/2z+0xTm+Z//eIctk4/vy/8C1VIK3Vp0nEDY6J3wn1H7hnBX
rYDvvEUEOlOwjQUrLdmu9ZVExYcqlq2sJ4K2LERYJLg3T6ufXX0ZM0c09HHd9Ngj
y549wlDLtIIoaPlijDuj0pylMxUuPlFAJrwEIHI9FXiUlylKLY30hLbrP9jWpjQB
AWWK72oO7mL54gzH3pLGTeZpa2oLCmzSG2iRmd7FG3RMdZZx7PbvP8guccZXOBXx
+Ea+/bwNWkabg0zV2pPdPrDy+KNU0FwGvjfbKvS8Ci58eDF4k8gidFudU9PPYjuI
/5IqJhg6GuXki2/Hlt2UP7M35lBC0P7B+0MQEyMPBaesH+GfUZFbAmGZ8liV1AG5
cu0fgxEFXg02NsayfVR8aWkfoWj9xyuUv9GIP31UJaDxcGup0vcysizyD3T/HJXE
VA6mp8Y9uH/bRCz3G0PnQlNPmqqadVAqTHaDrvq/pxnDexS4JXnvWYcX8+YV3XQe
RrKd2kaJawaQgJ2S7IFXgvM8m6RV1DPwkoO6Zd/Q17Gg/qlSRjPPPn7BiZsFObPD
XY+wMGwDY+5ymr1e85CQK+a9w8mgI13yh7d5SJEW0zMr2X0UCZOwWwC0Unuh5VdG
eHgh17pl3hXdLQy704SIWVQAN1N4O7JHLRZyv4Ryi9po6V6QmaYM7bMqSUDaewQg
9rMpbP/Oi/Hprg5cnTd5JRWtGnHvf4y+ixJwYQ2XcSPMkaIlQvliv1wBtoZbf69V
+RZMnDmM+cBfKrUxkl0eY+Uo6VjvhPBZ1j+FxF9j5DNGZBFgH4PcZR9wWt2c7Ht0
7OAsKPCbx3l6/WbLq1qMOydfFXH+sKXpnMeIuRLR/4hc3Pl9xO+RVRT7xe8ZLhlu
u9Yb+h6VOd+W57pOOZj3nzJtyYr0wcxANBN3pWlnMitgIgZSY9iyKwLJzU101Evi
hK72y0YHpGh46nDPOb5WapW3o+GlFAlMt2+UbGmDsEcL9etVTozqtvfJX6YFRjtF
9Ec4iBiS8o9Dj/45sXxIIiRCQ0YCZ7Wz0Kujg2XZmv/+vtWcrw0MO090Jbzo6EeP
q3xJxbOHbArOibMGtjzIpghA2R0tfBxs3iM9DkJyPjpfuNH94hsAPwjXMp1Qg8vH
gawQWSrZj8xAKxigaV8zENQVWtDAhb/Jh0joSFQq4wPNoDJA3NfDk6zgBxIoKdKz
R7YQSyNGMgykeRpNFzQts3k9GKJUTiF9fUmT0umSuf3TklYop5wgG/A+3YLsyE7q
sxyWA0htMPN8fQb4VP34+TqLD6uzMvGOcxegZ+S6PYKmpCT3H9eRGgIwqygAK8QU
tHQNZ2MZ0TEVvEPcENZhq1ponSYLlJQNSpSuacu+rxVP3E988BLTgsqntlRtmldr
mNJmhqEr2x1Y4ar2KnEMPEFY5JELhoqbx1COEXaEZyNTBl4L0QBGC34kUOno2epU
YtwKs7wzaD3ZwJD4+SPYdd3LLLPIICHdBJzlOPCx3cxzvKbmxNLxD5DCPAgQYdSq
VVx+enH/FV3wt0jQeqjkHIOR7XQREfCw9HZ1oHjRkIhbREs5Lu/bImzcyfsZP0gx
mac1Wqkax0gjMH4ZflHHJLML6GfX8RD9iRDG6VuIFRzhE9p1ZrpvQBfEpZXWzoRs
jUWT8S4NYVKTtuVsm4S1onYMBAwPwpxMLUw4fSxfhX9xDBtE+qTSt3I+1KDS7vn0
SSXnFrzmYB1NiRYjyNX7NGHuqzLOgyKuH09AEwaU0aHHZtM+8Sa+BES7LH59Q/ur
9jMEboWeQ1M3pguWLC1R/JpfDGoOnwfFkaEcqhS7qRrWNdBn5yQfJczjMG885cZB
H9cdrvJAEXJm9WHGXW/2zg88dqt5dYYQR/QbVIkID8h4QrK979mEYmYMSmSJ/L0S
Icu55OpuSPz3go+AhxdGouV0Dzmdo0T05ye+ztJFbg8GBtfKO6I7mrgMe48e1ojL
FhEzXoGXp1xRct3IQvfPeP7zPh8f5Yq9VznkfFHtsshg3yFgOffERNqKcuZrV2Jc
2UVUM8uWDTKgxRr3NLvNk8UzNhfa2iCK4dAqUbwzz39oB4i20LdnEnqJx0TR1r32
oV2i0Efqgs8wjeV/zaF9gBSQ8+UJHEIM4BXOcyHI17MllG2Lz3w16SlG6Sn8ckm/
gWPg2M7nDUW9CXfCs2w8gh3cSh8IIH1gc0mC2wCeE2OETTbzTcOKmiuxkPvB8uaZ
m2fBqku/CILaa/a+1oy4dOAvMyrHo77+fJLr6MlGDGcsM5cgeG+mwpE4sRHfX8/P
3A0oI9jVac0ZnYVyTNiY9QL/rkb39GJb0diUDMM3D1l1NT7DvP6myq79kczAEhy0
Hqc5WS52UaNHdFc+k0ffD7kJLNY/OVBXrwU+hkIUp9MD41rs3h9/OquJk4M52MJ4
tsEMTQBxYYWhG06Wsg+enw6kTxNyvtGovSXA+zXIkQXUAB6fLO+ebYvKAhfGHwU4
brNXFTukYZcqW4zhZWTcMJ1Dn9yS2DcWqM4FM3M/ryEwfcC0kWDbHQPizUBTho15
x8KH6VfJjZELROXoWpM4/gzjA+iNZGBQxYfpxlGvfeG9I43K9bHkUvXT3lkgTHg5
y1t7pLlc04BctfZzBs65/qHhuHYlqIh/gpuHiE+BvWI=
`protect END_PROTECTED
