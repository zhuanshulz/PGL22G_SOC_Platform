`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IlA/wDtLwOlQwRQujpztUCYHZcavvyM1fy/oTCg93xHfz2RqJ8i95paYUX0mT6j5
QefKnREAUfen6ICw8rt2lZAX3046kmefVmaukezteeqxmefXbmPalfBTWtQ3NmJq
M0mQbDA9Yn1CIWSnATSHyCI3C1vFpQVtw0fFIasy/CRFkyfQW3egsQw8ptI6Clv6
xpgE9dI7LZdgcu2jWE5e1vNvDXjiHDf3QeHzJ0waFd6O1ReTxxhNdOQ7GPnFe+YX
v358pPKGkSXQF0qmFD4Gc9YLeGgDSThyA1RwNhioMKjwpnNo1ui1F3uN9K3ylbIP
aXYIquzoEAQiwADZDF5UfVrVOKtGrtu7zvyxvt2o2uzjsmtujX89f2mjjOiP36OY
eO4E/m5OU76rn5HpfpZPPlYvp8OCV5NeaO/3f2OGzdFx16Ti5C1FiaNU4CplghDQ
COmPo7DM9o1I6nqN55fyxWk3PEtTIqGrm0OqtTLhqLyn3KgvEezsd5eBJlUBbblH
FDz+KyxZc01LWn3yIj1L93jwiDkk/FgJ+8fyzdhjjmGS6RAAndqKTUR1C1GWsP0Y
d9SSaMyxwT6qyTf0u2+dBi1Z8yTgErCvnWavJnSRqKv37IYq0hAOFENNHxBFzQaO
mfG/1XDHcNCouupI8defi741sDXaiBg1BPj48z2PlfmZKmXK3IfNYgRzQOIRqhJ6
zTk1BHf5p/LTOtycdH5YPYrJWJ2cGRQXtoCKGSj7GE7/X5BQaXOq1pV+a6lgQnxx
iDzBsknrLThat3YDyYUurwLdxygGnbYvuZzkX1KJ/z7qNdyQQLFES8/ewMumakq3
1XS83hJrS1zOM3Lth1ieFievbekgQl0YG4tWkBOBPZb1ck2MgCmw+GrNf4zsDZ27
6VmK+LIMCgafqDvHd8+MMYJEok425WVVbtXZEj5hfiZg05CjE/4ussVr0vJuOGNY
Ua2uIcslX2ASmfI/lKUxTfVwFBpmjj/UofygsVU4HmJ8au0xdJyhqnwMTs+gfEqM
gdZrPGhcVIR3Vb/GljeAJFgcUvkVQe46pD8qFwM8S9o7kHUPOOUdcAeDyXdatdWt
jK6nmH77L5Xx90jABiKZhc6omlF7kkDAqQeylzojqKwWJcpdE5B945gqlnjwh3Mk
gE6ve8bPJ4g1J+erqM1VEe/BXLFlAC5+wwRDAHsewIZdyfENGveuxU3a6bVtSGO7
p6cyzOrz+smCA4848VdUCTtIOnh2MtTFsmpONioZzRcdW3VHOl2v9DmPhl1qdBDM
uV/iTXxyMbLaxkRoB3sIJxVnwrQy1whIC6jWZd3MehCyBZsKsHXxnccAkYuIlz7O
+9mOxbLLAnODZtBpusnJhcYfzwlsk7NEE1ioV9zoE0BBEJNO/E064RXauKoXT7jn
Q9jTHsYeADmodF0pvJJyaDp8guc1Z/lRlwzb5eImfZsLN0PPi86mwkX/PFBQb3yM
n+kn0eUAW7In4TCCepOduWaEs1RShopfJP6t+RJA8sFrmSltdEynzCm76qAh3X3M
G1VTPd9/2EnzTURZuzRO75yxFkeBzDPf0cxoZK/lO9kuId/WuIHKXynUVTGESSv3
/NmG1i4RE60BnvdEtHnWAZfhhrT8wxlf8+rtzD4vT8bpgkrmZJmzjV0pYC6yfpM0
dSIag1sv9VGRWqV1Ch2cZlzXAjgmhJO/7DBW1AFtkgcM5HO4TCzOUc/RmSDxivJw
M/pn3FtxeGBnOn1xkGU9lnen02tZMV3CnELc5HbXiPeLjc1WqGO/2Cy/CGUEjpZG
ygZxQvCSjldrHWpmcLm84tTmkCd4AcSN0ZiItgjFSOzveb1rzSFCq8/kcbpDIIp3
v6589Q4Y2oR64d5rBFkzAgFu+snURqgzdmG591B7maIB2OBWVGTkHtbDVpoPpcqu
LbWdyZkdJE+7p5/EviUgmyB4RgpZ8Kxfc8QCwTv72XZqfrWDwOCAWK2TFRsSmXfF
pMNmacYB//wWREWvFLGCKMaUtipczJaeJaH7GPwHoZxCCmDJhUi37wU7yLmFzs2Q
Y2845dwYWS0b2kLSVU4tvxqw9tWja/AqwwmbYh92di6w284wLA3whcHv8EZfnO/p
JIjHxvCFcE79gUIKZ8WmeI8NDT7fUYTGSXQbCcnQ9ded0O5nOPrnGPBbfLpKdbj2
YvdR0M7EJek7SRDpbsivW3eftEuQL4a/8YyYySkzrXPRysPSo7+T1u0YjAtNC0y0
xNhGn3hhk+QuT6WvSdGX3pPpCNwHYI2TQoJJ0BROQDBD21nO2Rg9+PEULUuyXtdH
`protect END_PROTECTED
