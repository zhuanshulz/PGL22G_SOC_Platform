`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q3kDXAUb6vUc3gVhNVyidGIFSj39KZlG0tfpEn/tWJwXltMQtUuHrXO5DTXAmvel
Kns5Fp6GrrqJEcMp8huUerCJIhvB2iBSVCebPcSufbylOknF7o/SX0Urfi7HUObL
5/ORBrZZyL9PXrPWEncuyFukyl2roEqempPiYlCLeV9mi5Kx1UlOtjqQg7yxgZoG
fyE/bE4KuMP7dVSKiHDiGf3NQ/opPpM/1++dkAq6MNv801fnEMdV0px5JVZcCVca
1CSmzDXIPbZC5soPEov8t+ZJR7tVtCmYuoaeXTx9+ZpuzWGy+OfqHKs+J2zcNdOS
Knz3H9KZzQPufj+XFDAQBP3v49ee/P3AV83UFNEzuQL40oNibv4KWAHxFGdDOiTz
kE8GgCh4g/36CTStYLvxLeIQSTUQimuUVkoT56qIfMRXKsk2WKkZqHm/R0fQxjwU
87iTpawnINx2uPGk6XhVw5qpFno/Wqp6tg8HcRBLp1fLTRHpHpqZN/Y83Kf7DDW+
zRHMDUcDnw53WF5RLmHNqXGaAp/lFTKh4bFWG7GUz6g207dEQi+dai3hcR7Bso0W
FJ1IAs8EZ0Yy7UsL6gvDBo7l6BXSLry7rzg0GW8KKWwO0ankn0yJFBeOkYdtv1E3
8tsohyxciZm6rR5DaX/Z4JMma5PgcJY1o45MwQjBMr7bCQ1rJ6Kdbu7kfIU4CYPt
AUCIdoYIPvRojmUUjTf6MLpS7AxsINvmVACliIppkGJdp8hg9sCcrBLBfdRF+zTo
rKX8rhLz2uwcou3s+hC1oydh2oJY8PQzZrqHOP68dLlhnJzKUsvySs/aEAHMoylo
hf5twgUtxxOheqkKjzrc1xKJaN59Fu7KlibV7cg8w28XMD8g8bn5HRhrwHO0Bcs9
Tl+I4Rmz1uxuAK8ZRs3MklII7ItyELaqJWW8y4oREAJUEiIKGFgIU8LUnYfS9f2i
qZmXLV0/2+1cYXjeX5Vckr/Gy1LmF45rMsMjXEUGHKce4HbmjFigBSp//q1NUn6G
pNmGIw1s4iRM8qw43M9FeYUFR1dfXmNsKveI9Tgb1/2AFNib25yv9f0XAzWCgQs5
Wzcflv95fXczUyj8PluQVM8+KCgAaUwoaf6hy1rJnXQ1zJlxmRAJiYbUtIxeJuhc
XDmilsENvT38TqUMdTje5MsOJJy3Llj8yXzLT/R6sSUPO22HBRr/e+S7Y3ERGuXK
e7OAmk13SBP87vJcXrb1aSKdHFaqagRK6vbGPqPJMBCfwTkD09mkwHiXFii4kUc9
OOEgI3NvdMJiBrRFe6t85UWYGNG7jqVOyfi5IIJr8N8uXG3NS73ed9tMDP4V3fP0
6DviolWFwOQ2522iTY1thrzTe4b7ey19vozl2NoRaJe99eCnPNg2CnR1dl0ar5MB
D25aVzS5OM+A95mqoNennRAHwzrp+yap5OMm0Wl795qk4nsPCE5bQIIy0++CSICh
34xx0UdvTy4an/myTjcxuk9NnMWcepS4NgQDlGcLd2IeTPUE42ANwry0CnvjYOS2
ixnDEeFRHk/Lsg5MXYchu0urdUuNYFEyBh+QUoc6e/mwTujtBLGn+QiNfJXHiuec
MdeU5PI/VB1LyYn9WAULqobNadjm9RL2YhOyGsIkrunOlLtwQp/Gv8IbkBrN712d
KGkrarhOy+1x6FkR4z0hQrwo+XV4FYv3b5q2yZ57Ap9wPcDxNXCsPDpMR1M2Kndt
bchb3x4cIrYZ1uxO+dcnJNCBBYmBhpctffoyymbEEToyfWebNSJz773n7yh7q3zk
GB38FC1I7IYqksOXrLTZgg3bWV4XrrcnfZ6Y3RxNrYyJHMofVJYFRLOoPUlmMJ1V
XwCetAe0lD8TMSHRJqSdCdOwXvOFCXOIORwBxyptobqx42N8mYiQh0uhKMjvWqn1
mdgyrZwmmp43RPU/sJ3PPE+m+GVBhxA3ywe5Nt/sFu8AaB81d4pZkzeZnz/LmH0I
rDStbbe/S4CL22Uep8NCirt7bwTyxsxQ6/CJDmVBOcEHyx9aZ+AIAihajJ3LO1B6
3JWDz1guhszria3EIQsZXjPRzlI5FGEVOcYjqolnFzHQ2Eg0VwedZ7Q4U3ndLe8T
sO8NpoPfShMDSRgjv/Ja/hpLDovuUr7DEEvJHWMmyNHa00xRJUm7qwi0G8OAapnv
sQYPMg/pVp9rfU4xfqrbDk1xWfjyjV5gy0ujlcOPnd7icGedOEc3aFZH0QVoVMf/
RVeyhVuO21DZDFyR2rsLgN/DZazC851sQUn6gC9Fii0zeuERckQbfhcKAN61mLuk
3aym3kY/PQq5pWUqvDOVIsYlpjmPsTjKa/wM/SzhWS6MLyd2lkjDsNyts8por7ba
xCEDDHIVJexrrXTE416OFHYBUuA5Qr7hPcSt0A1cORaYMrjBlIricGFbGMLpKVLH
klv11iS5VUBUmttX90//DdfxYMXhZ5bGh8U6bKCCgZ6Fasnpc1cglqjUv9NnF3C9
TxsX709yqwGiCNkidiJ1/PqjjaDrbrFv19QMr4ZOp9zXKCHLqm7/JDqLnLPK2H7h
9XajA5ptB1dhq/eoyjm+IULlOUH3XLp40/IyqsRYDtg0vfLZPFK+eA/QNo9DbGrx
kvtr/NICuemmDQ+8KdS7jpNtafa4EtgP7MYnaxtM1CDFujyD4SavmXQe67THfPx2
0+vB1pcmxKGHqMOCRM347iS8lzMl6UOsGoke+iq8B9SKFsB9YHeWmNah3wZWKKE0
jCInMDdBuW4FzAbUmI+znRvQLNfHYpc8uSX3AbQyDbVidw/xhQrMxmkS/rq8SVLp
vtr9pNqQnw0hBA/FWPwJTuIUPhouLhdDm3SIDQ/tw8GajWe4LvCImvOSW6h+H0T6
xXZIDMWBPJ4Zg4O6mM/xumvMF9g2v50Cf4PFLjKi8rEhJwW3v2dHJkFx0qV79AY5
xN4dnL6FSlfvuxe9a5d4ZBWsQkR1FGGq878rSwJwbupnkRKLK3xMgfk2AoKCVVdm
i+6nZ9MwK5+x0h0iAb6V648FYbC6iVEO/hzeUYaQE3IjFi9+icJs+kNFCp8IzaCw
vebAl3Hg19sGWWLN5MmhlGjCWcWYH2ROokJewytT0c7uXCwbstjRjBw3ObBzTXh3
UZbeXP9Zct8DxIsnBrwFw4eHDlyhaAnR2jWNfCOXBk26cxmgPuLA4sW0os1rsxx/
bgOX9AFJu2hsjmfGxQ1s2Z27Av4rHeuddH5mNeyILIDxRMEcTRvJvsIiV4EVVGAA
7nIW6wCwFAnTOpIVoHVc7ShE/UC/cmuMss4Z+DA5QRqVdfcRPnFDZucsrCQlmQSy
Sjn6ifx1qhIgMav8EiG5jQ2bSpV3nscdBCOzMrjlzzvx6REMgAZqYX7QeCbo97kW
WpjKx0Na6fqDw06ul/ddTQjSO0RLwX46PnwZukCMOnm2q1zFBg+iMVxiy9zqLAor
qcVBVyriO11NHJhehF9JR5rUMapy4cp4q/e2modK7pBsWw9wfiA64RoP+kItlZ8Y
u7wKx5lSyKWQWXVHOdJaHyC/VtHok/AWO1eF79apLAiaw+h+nT0XmFhjV6AztmI1
cmHFSUnUxmt7UL4jQB43iX25re49tyeCVPSp8Mj0P7WlH9AmPUUNA/td13s6fSsk
587YaMRqGk/geOOp6AoPRhfUfkyE3gn9rvKXrakkGd22Nbagp7BKSeP1GDHJmj6p
ZM0uLWkWfGpSba5yw9I/Z0lOGjkIhc9RBL6xzNuKgdkdN9QAV9VOJymZ2VDWtTvx
0K24PjbAXgH2f0Tf8R1xDl0rye8Bt0bZa7POaHv10JK90Q3d+3BE21bAnrPgIZVO
SenG0J97b2dYgbLjbWFZpmJZJQudKh4gDLJt0xX+3JfqFYx7tYvFmQjzXOL3SmH0
C69HYFv8+x4gQlq77zOaN83lrms73+v8EzLSHRHNlsT5N9dLrDWZoKBYODL9OZj1
+2D8jOMAAZ/OpK38pMmKRV9FcOsdwsRKlr9raWXNY2ktnjTax9nQmIcIdZJxX3Rm
natpcjiQ+VPvln4xM6iYKdSrbFbklp4hgzc1w0xV1hXoPcllwi/scg+3WSXa7GBY
SD25xMYdrO+RphHgMWiZ/blLcdWbJ23Ararm6bSTt+GZH3CuEGwnIj1sR+NwK+HK
MsoAL/DdCNACDXqSQgo9AhSPqcZlg9YBs8LYyGt6IriVqzzzGtJ/ccFjstp+b1+r
pQbIT8/YckwIs4jVOy4CI9kOzBKNre4aC2Cj74CV7YE8DmI4mDRz3Uinj4CibJcq
swhvDep+xailzh18RlXk5BgQv5RztyLZdFZ/PR8ciz236L4fliStYf45un2AqgOp
/lkcP/PuJqlLYENZvFHhPkXNsb0zNFOqdhlxG4ato0IiKSXj33BNrt8rI9C+CRzk
SkU9rB6acvw5y9vQHqcaQajbBOW22GZ+6Zh/hsIpj/cOZymTzJAY/GcteiSFTGfF
+GNXdEm5Kd5k2YXHbVqshLPM7iSBa65Eb2PDXIsg2fhW9xw1kZyzXkWeXSQtZiK0
YmNMV3zrMmQIXFaJiQShy67N6ouYy1mcvw3UzDJ9hnYVrvH10ZCMmk39tAxFgEFO
K282EDzrN8VTZLX/Ov59N8nqyGXcaF73SFpnLftzBElBgILabW1dHp7CSaTR5kvM
09DfdIOehwrBEKS8BToRwcQemQgtf2oEs5W2QRT4L+WohMj1VkIHdGfna5wDLuhc
BBM6E5T/LSCdsU72zC+3kcHhCzoKlFkdA2QNTPNmjB48jBNCZ2CUmDKdqnUrJxhN
v6Hq10ewdF74aaagld4tIcMhfXib0xEWjsNiT+ASbYDJaDzsNJtT8nYJwCkKCc8m
VxXAz/gHIoPN09ZDXAXdsS3ng3gIQ95P5oi6QMaZx+YzK5pk7WswBSpcQEJWgb3N
rtE97gsRntE+L48X3bY/cT2ARD8d7P3CibAh9NXKHN8eTWCQyhTV3cIBnUtC6R4S
sCemgC7yHdUH/43ebqUZMSnMZ/qP0fLAiImpTVbXgsdINFJVJ+DqnDNgj2WSIoQe
wAh/N/y0E0eIkoSWkZmOZVn0dA2yvDUWa2ZEbGhRmMi8hUBu/TQSoBGQnJI6kOqH
8H6WOmAV+1wsoQH4V3OE/1b7pnmNNYaRyzHIcPuiNGoDjpoeW1snE0slvAbj4oLl
yqIYdfy6PtjzdWbZHKloBID3drk09wVO+2WCQBViGdo+UAkQBrngbnQU+YvzZN9d
voGdnOCXh9bfLRfXCImMlnLOFsp8ZhvuqOb70GQvc1Uy1E7M5I7WYqFswRMyJtTx
8VFLUTq2hDVRSkEriVG1NlMydRhIVRI37EHZtaCVy27C9QDcYHe/1fKHdxRlM2cT
8Fh5X9/4fhwPwyLBnXd2Seh4yiLaWfksYvPFPlc3abe00/MqAstDvee4n39RYFLI
VdHAdrodxGcSf6Xspmfn1J4XbKHn3FT/6XcGtWEIAExiihjdDIo5vhW8w0QtaZ7Z
3kjDyg7wW8l/WXM8kPKsT4px7mhnTc1gymEEXJg7h4OThzjuepKqhgQibXZA4WbU
w3EZDHygC+NmHydoSSLLvaAAG8L7ncZ+EPLdvUxZDUJwjZNIGWy44TPPRpAXERd2
yaxNQt2yjxpwBTn3S6TZ5NRG+m4B68Qfya4ycpQcIhYp/9qZLAtV+PcPRpFD0MHH
2QV6OmJZADDdS4/3cxWEF7l0AHRSRTh/QDq8bXbY6K2Ytq8dZnmTpjxPVOVsUcBP
JOtm/5T3eXj94kzaMvGgcAn+RUGXs+U/vVDn/81IUVufbXzVnrquRQdLyd1/53ct
WxThCe1xkKHM7fQLSyrqn/S4Neh3GD4Nbt8rppax62p1tpwxLRPjffPhBfRCJvKY
fmHgwkW7cGcwuH+Agv6V+4Zw170nHl4vAgiys1jgtjAsSDnUXQUoDwuVVd0sl0e/
7xtgHtzIY5LhfAnThrzspUFF2B3YV7C2bfbJbmy3huge0Rb8PGo893AFMgvyhK6n
aHK6t24my1x67aeOPBead4Cc90YapZ3tJGa+z/5vOW4n8HterIb60bXgj1tdpFQa
qLyoXlPuNyXrpNbuk92LxwktT5lo/EjmDigcIOzNtSwNEa99pi0V2df3SPJ9Pcs9
k34xAXe3EmEGLhHrw9mscWz3rBmHmykjEwkuTRYM0Vn/ozhPFMsAzieNw2CD94H3
Dzs0mlH6KhMpkLZAEqeCvSb9SlfTUJRcdJnQqlBb7LGJM2FoV5CGYGXSpKdMqPLj
30+qm2WVZAZCKyLtA1yLeF7a+SRDuRP5LBho12KdV0X+RWHYrfhidZvVy7v9TIvz
RlapO70W5yEbcwP2M5VBQmwROhgNmIkZz2tYp35s+KYSwwmGbr4kjHGvONvP0TNL
RYnBOIlxskIjZLReXBU40niYL1RFq4eZ+edouh/5+yWpgl4gzkzFWMjsZ7Rj76ui
MrKhvPG/At4XnH10f6HZO0NWNse4fQIOUHKrnFc/Uow9WWju5Fnn/Adw2/U0KCVF
b6vnxKP/Tkhd5qzCG/XFwFrl/SUS6P9enDECgANo9slCgPgT/Vmc4Hq+tRre+TEc
py8lJ93VK6DffsUazutrViVfaQywyOO7n5EmtJd9dlQN17OzvzCZgPnfEBD+2Lyz
c8+/B9PVxPBEacEysIai9G9gdDmCy9dldcnR5l4CJbm7cWNvU2mYN/s8h8TMv8kJ
Xaf1CBcMezoT8YBou8M3gYNS7T9MCpA/7cgUaPjtn9okJFF1DNCAlKktR+K8BAQ7
Aqqd8bPj4u+Z78mbVS7drU490APnUUfYf6dv0sRihMvl+8O9apbJ8NohDnf70/BM
aHLVAA77ROtZfZOp2j92sx4iPZVGZZHFqm69gddZ/ii9GaxH6fmrKcann6Nx23TS
mVngSpfTziDEA5cHrMuALe6c073kRc5EveLs6bLYUhIvCWqW9FBB0bXXUA1E4KSz
NuUH9/yE7fmi7ntTUhx1161Qd28IMzHeP/3klGzMwrLRvhzOkooOCuTaUIS3nIX8
2Y6ge5KTR7b03D/IeIWSM6JPhRDkMkY0lRoGlMpTsfjo0JCL3NeOPE23vurdFU97
XkpkuJCWVB4VvjvzcmWt3Q/aRHqowhkpK/Zi6pDggJQUrBSQz67Th0W64ekp8EXd
AxioOpYk8D7EEbI4cS0gRwpXjLdWVa/dWBYWzyKb8F4gfL4aoq1FU4m0vTEkqWF3
Za0T0lTQC7ZfSj6tCDPXoWy5LqmeJjI8V/uBImkHnTxf5k63U8nv4ofeH5yJJ2Xf
LHecydAXeGYpN7cS8CuUUg==
`protect END_PROTECTED
