`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7JvonMDisHCPnmFYKnfYcwzHLtXbHUdHML/I6nWZsn5plCeu5PaTJrcEPh9GpIgU
++AMFfGjz0ac8xTblXBE9Q9OdWfTh67qim94vxixHq7cp5zb9So5WOzQ84wldZ2/
idB22QGqAh8H+b07pGqIMYuDgGnM72/fxQD6XzqEj5n6gLm/vASqyWlpDUX6ERYM
E7WNKGonyltC/VJsog4q2eUAYpbcM5/17H4DYQvataQ97Qe5flYZay/oHd3bEwLo
JpkIw7DdpCVjye6UbO0f6WDrgPk9xfaxquT0B3N1EoUIiThGXwhV5JWmagxFrzCX
jhyPHykj1CAp//rOiF+GP1MeHfC7uEbpJe84imsOrpo=
`protect END_PROTECTED
