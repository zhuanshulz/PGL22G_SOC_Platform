`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kJEo/3Qp2l5Ucimph0qzs9vQiFYOlVuorujxJUmzmUjfqaRNgGrV4sV/UvQmZ7BF
CSj1xHqBgQEMgtBtoZPQT/t743CANwMXExcAmRcwq/BtThm0ohcZOnufs33yMyCx
9fqbk+W7Beh6LCJYXgBr7QXXw2mu3sRKt4dT5YBui/1/3XdfqGMBm4G8y1PBDKvD
dp13C6c5rrMoAppHeVsuPjc7YxdQgUntdk3T2LnP80b3DRhf22qbAxICtXpHN5lT
1QnAB9gAaiOvmmWOzrNId7G40Dg3wcxcZOU4SYxr+cDF7n/H65+K6Yul1O7WCJoE
SJQMbRDjXEt4C1rsuqClU0RzRPJ+aUBBCDYG9OTVlkE/PnHKaPEuS+5bN3aeuFQ4
ulQ0spBbJ5as9tj0gb0/3/tYFvW/yCx/WQNPDHplRMhbwmfEZlyiEewiapfhfKe7
APciQnvGf9hYkONuIHzA6bLZtPJRDtc76e5pQ0or2a3CXq0H5UXJZdhoeYrjneJE
NSjug6FXmOrkdWNPZqnfon5/5VMbh8f9JDl6bPYtyQOKCf8w9qMaOn7E0X1Gxl1/
5P5wsxNKUOrsoWTj9hL0/PnwhdI16BgREHLMp4Or4tallEhiCXpfwLhgHDpZygnm
SBVE3QV6HZ+KbQf9658jcp9it4SMlRPaDcui8gcKK0STQFQ7reu355UDkcJ9bWR0
7bJtO/nDS4SbaIaCM0qqz5tFmVb7T1/vuRLJzLxUg16ulr15aKW5X+Ev2WHOir1D
SKy2BPGmqm9DdUaBtGjvUrfpBg9jmg9cr4h7spaVv8NG/eHlaeqm697UloL046zN
64R3kQoL61I1DZ9fhVYQZ0yjrRnxFZ2zkmdqled7Mr21qNbIlXMUXOGc9N9bc6tU
5oyENCc4WZfGkQSiZFe7onfxdWJQDbDyZDDdKQ50jJT3FJvNZcD2mQmOVJW/bisn
joBLax/DES7VzEfeVkhAoruyrRc5Dgsvd/2/QS14J261pc33u1dkmAn+szTOJWd0
ewkHJIgq9rPAiJ5BoUtXLISKzheqD9JITSITKNndH1k3wEA3l/MJwWSN8D+G2rl7
FoB8w/tYnrOAgVZiXxMRn/8hGRZmAGiethKUfM0o3Wz+ZpKnz7RqJAsofqw5E8pB
1VBm2xDSjYbdVVd2es/C/fYrRiKniXlSgb2VKyGnguE0S0rlmQHEWKtqBv1vTWpc
3kBpKj6FN87RnD4Be0G1ccFAAMwT9ls4NwrmccgliePZeWKE1yukRTjpxdR/KcPP
jLu5C2mK027js1dsAx13zy9Opur58OkGiWPC+YHufhEY6miuwc9YXiOUBPqyr2j0
ICgYgfxVZeMS9jZ3liZmn04+PO3f4djAOMmaQ1mUd3jthIyj4AXFj5jcm9aCkffz
AhUlJA0dz/KvJc12Ml7SADLESsrZLo00p0aBOi2/nk2BODaAlHhbY8oCL6idJmaf
2U8WIbzxMF48O9dxQJjgVtMgKsX9tft1aDCKUQy1vSvOM4DOPbPPLbDXvNl3PfAF
wOwCZVV1QINinvvZwHmiyn+1y7klIzLoMb/6Tl/ulo6DzVb8YcfbMRQBquAR518S
xgL9SOodomPBLZEXFOUKwQIF3/lQCpSf3i8+KveGNxqymi//HvBu0Quqn7Ap4M8F
aJ2F8hW1rkG0Jer6tkDbB32guXQYvGf9wvsF+k6WXOtgNwMcjK/ufYKPS/PxZfXx
bntlRw439pG5nsLuZhlCcJ2txhZAQ6PIJe/HNtS0sT2HQ13EBGtvrv9ogdiYkPfN
Oabn7Y+ESBJWMnnG3hM8+E5M3C8JbNi9i06acaZ4EZsQmHm+boOiuigSN9fNRGhY
cyDD7WGHu+D/Epak9fcdwDsUBQrmAJ53gRpCMmTMSD/f3NFkSm8ZlcpOIbd5io2k
ZZnlKUUpW7DcM7agPskqKpWKuFdSy8w1x57ze0gnc3/z659CQNDtDMSLaaTqowiD
33dnQPy0dEv6fRgnwJORep9KTrlKwKba0DHYvlp0hHTeU23rHlJdEd74ifMPQjqb
+FcrwlGv+gewPq6JybibXHLVCpPuVNWEJPY07JRef67+vw2hF56uBYcK86r2V1wW
5Lj8yE1wXAQl78Nl3nR9kePRc6LYL85Ec2VV8qwVyOlhhkN1MUppexSk+403bsUk
PVEbBCI+pkELaWEX+RyOEF3xVfOBTBdnAUFgRu90Ybr6uw9T1zFtFQiF6RFRWzy/
38+mS/xS7OYysOnOd+fadzMTMs4H+l0mHoW8B9GGvEkeBMEt657Mz7Bee6BbHH3w
tqCSN4sPMQSgeHW8QEPX1t87+YdITsTyWs3HdTp1UwRDuIlp98F3H1yumYgEWBvu
JYm/FYQJ8GPUEH7MrfSoL0/NiXHzo/3XIo/YIAz/X7tPJ7Du+OcTQhrJG+VNDi5t
SFlpgiYaqM/+d3LccX6fZ57vetdvUGsyJWIiAgDK2HK83ajYmeLj80hzf0iYIgUO
VDphCS+1520ZENzPKZwogq5eY1IGPppfYk5qSag7IPFda74grayZ+9hoU3W+HyRX
H9NOOufv7gIzgkQVOLTt3LMyzkMfvMqlfLq6EddzyJENygbidMIPfKm36CqsamG8
uEaywmOnZc7FtDAEdDkGPSWlQnjK/ifgjjVJHVSC8ZwQNqbsSIvEUVU/DwaRXaSL
zbLcI8z6FxQ9ydT7gt77O4+U18t70JkBRANKTdSoOp0P60J8Zvw+Iv/1o8e+4Xnc
n5cTGfn91TtCoQNx8ts0AZl8Zw8rZO6EapMeDhxQiSH5WJnZ++7uAsDtO8xWj8uy
CGSTPlSo8GLejSMnDM0vIDaq5xCBNi7H3gKlGASHcLJogF/s/hRoQxQPb5OUTx7s
17GUUbIBHn/W3y5V3ekeSM/1POWhiVDHivF46xyqEDuw0rvZGqasXIuIgHjgeBDy
c9H29L5ElVlohAqotSpIVzjKl1DBkXbb0Tiip/1WWCNo6fvprJqeiWH+ZKQb0lCK
l83meQyV7FYPyo9t5SWo6644Cm/6HTty5wLYxvtzLv++qDZ5JL27wzt3RMPJ9aKD
AEDNhCY0XCPjnAZegbQiPpkrHJVOJGJFWrlL89TWXOcE8zadIRvJvhxCQ5EjbLQH
StdyqEd2qvRY3fWVk3ZiZxv3FXZnIZ8mR1CyQ4LBLy1UdPHR0wexqneFr2CWD4OJ
dXkniB7DyL4F/fQ5cP/wLHwxsU+WXee2Mo4NY/YjuVm6etYMhSEQI9le54ohktgf
rifYJviBFiV8wnJRfOsRWZYZAdzTjpLbEFiM8stIopvViMAMc/XKeAh8d7zyCXr7
RWRqfy8/6BpiyEnpqf7HMhHVbTOH+83IFX7fXC/+Fn6QiRFEFF9AvaEL3A/Y3ff/
4fwq6DWvX+vdqAUlcZfer+RrpiD1xdKXGpY3mnI5xzeULSmrUtvDoQhFLwoWro9L
kqsqCk5HYuCAAF+yNP1xe/+kq/7sXQeMnQcBK2U03Zrr6+lRkrSGvMkY/8drOSm/
cRAkd25T3QjZ2PEsZEkhqtjT4jgCZpK3peIBpu2hxJqdi7ShVHGiXmwzNYWXVIfc
KLjJTV6OjXB25C/pgBj+gcS/4nZKcWoCZjXXkUt18aGYW7FCSucBg/CmqvIGXqhg
n7shltbtQyQ6a2Z9E5l4VESQPJh28EMLOkVrZ2j9DYvE4I8HuHxT9/xjjWF54l1Q
yI+EIeQeavwhPbcCJC/A2DV3lEWla4IzdNxOly4nV9aBvU7hxvW/C8lB2/ql4MUC
UXoTPjiniyQ35wk79XebZ5HBpcFUBVRyOQkkux0Xr+GWCGFdhw+ffq03FF8c3Z7l
ezYujxNcaK6bRV8+4LIN04j8B96K76UZZ/krxbFc3yS1dd6EXaz52ffNPlWB2jzB
tGRl1WT1X7Fq/8UK7DkuIm47VrbvM0mKYzGMMB15+rs4XfG9tv6QMZfPqgmpQ/kP
v/aNCrsoOc7XDijIq4EyP68CMDVKU9snBYzI8cVMlf5vMNuiv6/IE5hcxgZ2hOG7
+6e/62KXK5eE1kTCMz9mhKNzU8UNwUmxdg6faSDxdh8yMQ5mBjd9Fpp+yah+jRVk
DIzJPphbF1YhMy9/SGIzFY0YvRQm9s/gar2JQiWAXEW7ijjHBhTM7ssPtJhs6rwK
5TMDhh8iCJLa7pRJ+jJwlHT2F31NIbt8CJrF23x3EHa4sppOKxwao8XGMiTRls13
LIuYpC7N5je3g+29y/oAOVbbFrHV+S0CGqgNsDCtbuf1M0PNINYCHAIZBTmmVofp
vu8RAdGPgB5B7mqkDFDvcACgiDCPtlxJWJDcZtdTx2UAWfe4esc/9115gYhWj+/U
iFV2xE3h0Z9uyfnY9THu7xW1GqcCWthlFtruRDm4cvlJqTlybySkG5XYy+H7pMSd
Gs2ibwh8byo+agueT+ZpS1aQM00ZG2yiOMDa3SD6Jzp6CGDMJElP0Isvp1MACE7e
s2NlINKGtTK6oX4VQQddz0hg1nsvDYHSJinoF5rrU/Ye2EieAPFjsa94pu8ESl1C
VADnU/0wRhLRePd+yoSC5Zt3JqPacPDUNCTOP30kFdm1Lmms6E5QELJ0Ghs/CLAn
dDs/igK7GaOY985TYRC54i6S5bpwGWy9zcfxDD3ol5wzhVfLOgpBj4r5VUCm/dsZ
IOJmScdbAmrb92HQGAzk88gOIJI35xBkvz1BVWUEcwbjEiRAtno+uSqiHua6fsRZ
afBvTx3l658/vMzTdgWNQHhHNExRxfLp1cLj9UASaSYc8F05Q3BIulKJT15qyID0
zBBJh3XwyWbC3ai0plz3V8kBDXJ7c1oOoHnjwx4zj0+oZsrDG2+FdbegPhtfO6B6
NdSyFSG13vbLffvJT9T7I1D1+W99ekFXV+E3hc0+xIAQHgjSTkkkEq3pzK+U403/
K0ZB23gRRme4x0oRg9O8DoLcu5X8ty+lQH5cylC3+qszvpxbny5/uZGxgvkTF3xi
7QIu4CQNLFLaB9FCDKr6rNiK2JW9ipP55X4bpVdDf5IEoa6SKU0K6BzI9ges6t0G
SjMKKXJqVooOwVyzZLb9u03ppiyjSr9bnbRs6Ar2k0+JM3yiML6fAShqQV4ogtyO
MLlLQRc5DCHq25sUWL3KutXFlk9JjGMKBuewoFIoIT6+CqvVpmKLbqv3D1c5RUd2
2sEhDkP5TDADF7p+jL2Ss2HITHfwL/1bfk0rGB3cbnpra4xr6eOCL1/J2Q7Qjmo5
09pFxVvode3rmI+jhyP/XSPEYYXs7zdy9VOUKv3nePBh3vdhxCXN6d2esIP9Z/XR
yHiQLESBHHA9TWhS3GW29xUBFqfBAXwUqQrWkG603p4VmDWaFGuHvzqs7tqqaDky
JEe+6/hTuTwDeDJJ0W2GTSWA9kfxOjMwhbG4g3+OUCmvV/1zCqVVkW8B4T5MXb3H
WWZETrolW59y0Mx9asH6GLU1gy4zlACT3gXloVYpeGRU+7Qh0PqRgayYNcNUegy9
mvO0SmhcK1GEI5Fji5HQTrnMlSrdEUR8KPFoqvRguBUECtUskNTsBLHO5bPBURwe
1KRDvNgdPUFeBnIMqqalZJW+1vkmoAZJWcaRazvkLMyzDn/rCGC/vyQB0c3VDBFA
XgC2lTlurw7oFqz9u7dnRFoHfl/92Dyil60jmitw0l/qK0Z3hG8Q6eZfEXo5EiMJ
X2j9qJjzvHV7VRK69cOEyx/sgwg/y9hXz7N0OS7v3tj2UIVxQaIM0uR4JjOg8lw+
QzjBIiXH3qwOgHGVNhsitYQ5AHxJRYivmWiMJNTCHjTVPiurWJk0IUSu5fjQjeJq
h3cpGLk7JMG1Y+tsCsgnH4EIdfkS8hv9g40vjqaY6uHbYR+OksHBfcaDoBSslRm/
oJoZuxOPbdiT2PjxPoPWFUcHdAnyWYIaEXQ+k5VerQBPoDqJ+oTwp3Kr6L8GZrQv
OKcOs+YY+p7E5yRE6THT+L4elqn3snT6kgC7iv+BxzGAHFlruFxipF12eMCQKLNf
uWY4qInOva/eeKzessI6oXAGjdrCELHXzArZ2kz9c/cqIPazQfBscGTN2CEhnho2
g/fYfFg/d8uIa+R227Tpw+cArGVst3YyDfNYrvTAk4XXxFIFHngAic2I8hMaA7D+
E6NvqmrUS9mFk8HK920U5TduwG7SDu//DGbZQfbeij9oAdWTqSb6G8ivYWPfBo2n
iFNshbtcahSDMqOds2aq+TquausKaBbi9Gi63n4e1SrzW2CjCG0wGxc8w1a0grzc
DTIOeup50hthfOmw7qrT9b33SRhQBlwXZwW0LIMjaNhdM4ecXUcSqH0oZTXbnOnC
5hY3TtRagUMDGl5R8yF0h7qVMk83FsE/5XrDqcgtxnFxMW2YcNgxZjmwJTBldTLw
h4pSxOKmQH5hYmiASU3s7U/CqUF6kgGf7naVfN95z+aJ58vozbOVqEdUiVuv0J2F
RJYKMHrPQ3dLwiOvSVmCDr/W0okgpdYYrObiOmKCqeoDeLUNVu6waNppVqOTDXrQ
N0PkENW8ckb8YX5v1jnaTHfdUWzIfBq+GvrPXxtgLB9qcsSBd3Xvp5kaU6Gz/LPF
pAkgq2gQTAOfYpyn4lc7/wC0nQwYYld7pp5rXd/pF9HGEd7mHOpD6yct4b9gPGxG
nAgf8dQBXdLXu3WuX97ohD4wzJcCg3msLp8KzFPo+abuABiXw0UJ2Wz/NzV5Lwgr
pcdpNVqt0vs4817fFVOJA3uCK5Hn5uk3g1O/nhK6Rpltoj9GKvFn+lO8MPI9O4WX
feEdZ5914L3wa1vosmbN2+m/hTBAIrJrZHggzv5CjZYf8TVudRdtgTcIAwbbPYPH
ngUp6NYN0LJFXyqvHNfUzKDYp9m9HlYPo+NZ9gulZymp9abMSIXbY0lm1sbUqX6a
2mMFZvnEFqWYoX3RWFNsSfv1x3rSi/iHsxF1MhWIGNg+y3Q+Njgo66UI1Xhd6PG5
9u6KhbLFMtYam8kFlTAelwcWkRTD6NsV8p8T6/QUTRxUgOa7ngm0BVTxpgVNHn2i
OTGpPEaNvdO7pQvzGVheKiv8oZ5O6iZW9+kn8sQMPqGu4655yWAq0MCR2+XAdupV
RB8HYCHOZX6XcVPhf0WnoOrem58UpkeOxcSlYSJeZEd/fRlhXiI6fbtr9KPa+1ZP
9DI1vHLNzTfgw2inFoC13oySgkmj7FZ5Jq/Svx/bRi84Mr4wVlnC1MnkdAMHPETE
BDFIzLQgtLtf1HucnwUCyJEEnqd8cxSi0fn5nOGLeqgFBFjPibNETQJMCEdySqIk
3SrN7cRoiSD1txAw+yiLoXA11ntdMmo2g6TWmDQyNdK2Gyu2WnrA0sKyCtCPpxOn
oy8TT+KdGFs+P9pj6pgzwnPFIDkRSvUMagmG/LUdtF6zR4SNCNukBl7XgMer6rh1
Ucj/nnuqdkm7UveahiI3RGOo1eOIF2YnDREhnYt7hMNBr+bNyymizDKBM01EC/dy
1k+NcctJqeoxfumOP1Tdi8eSwqkxTQ3gqd0FJBTpyF+b3xNm/GSR0dfrwjdkNUgx
s+CnQpz81TlDBVtT5hroOPyPi2rZVKpdrZUDfVYIKMO3JF4sa4+ZIQ57TjDlmdp8
KdnS4I0D4lERwayWXLIhKs8Re9QcbG0koe1vuWHDe8CFOotF59KWpVNX9iV/m2If
GC7tE2iTW8tA7q3dzh6RVgf78IvhsFffYd6RegitzlV3p62JfVhzcrx22FQWCSkQ
Y0uHuyqdEQkvGzCqR3Awe2t1JDIM3D/v3pPgDDT8eBMmwZh8L6HXVrDnMecrNxk0
yAJ1xm5FuQIsfn4IhZFd2q6qbVECWwIPzfNAfzqWZX/VnW8g4iPSTjXMUVm+FFZr
/GQSyQ7bLYP0wqqWFIAHZSHkkrReFJRmKZx1KfCpCuyyKvdNoOWsX9JQnYwTeRNw
+ffBQTdsh8P1R9YExkyZ607liZ8mRD7wUT9OW9Zx/lc0k81cRjzO07gY1SOCNtuJ
UzZlDwflMmSMypuyA/ZOsIQfg5dlD2yENRbQiGliLddqYfIiXcAWraHpAudJI1H8
TZBGfCFMbQXgweP2CzLgCw29t1ddGn3roY2aRaF5/KN9DF6VMgK+OKVr+qgOuKiz
5lSBQUHz0ciD2e9Co2Bv+R6qHCpLsIpNZlSjC1Td9FcJD38kx9COuqRW8uOfu2Kd
JQiReXphY5LhanESAR3F2mwQ1nvcVT9a2E7PPG0bswnBE/wwC/ZgOKLALi4INm6L
kL264gfdp09GqOVtgwOjafWrLnxYfa+PL2H1IbK12utgtleDMMY5laycGG78eoX+
OVfxY1o2w/1yUr5BJaf1GIsv59KeL4/oREUbpdW4jw4iNwB8TIf3W2YOWIZo/Mcb
MlygjDIRrINZhm/MzAgf0mFWyNV+DISTt0Cisae2GZfRP/cJQOCA30trUF0EjLNN
/WjidSD9CNSFvGR/tcbPKOJea3jP12c2j1NBVtUBGjgQ4+5MBKhYd0/e6UEXqbVG
mUgSuFFSRkKh5E5xOwNph/TQLOt0+/mHCafgKm+R9EE41C5hPq27QE2W4Xm3mCPc
tiIDnjSiPzS+BKlpdpOk1ANuywF2Vndkf0GGj6mPkwuzAb3HnRWHe8oWR9dv9Txo
AxJQniLXumCrgLxFudaZITxJReLg3MBlRzcKz4DRTe6CfbAijts6sFainKd1F8uR
x34qejWrkwEC2/sPI92SrrCPgpdQmCw6m+mlB8MrA29FLXAHJ2gtyp269dk6ODy+
2ckk3C7nKYQe1+0C/VCkrBkiJaXw3naVZptXvtbdpJd1vVRl9SpJCPAvX3+RKmsO
NqtRnQdQcuu8+WP9Y/3WHy6XRARMmzdWz3sW7btjY9b8WLgClsrWEiuUZL/TyJns
aLMrFtt/eHcJjXqsRfImpLqv7UK8vTwTkklWXVlAoi7V3imfsV4K3m4SFYFpn7pC
MiNHCK98+4DqJGuZJEA95tYl+SK0ILdGbvOlzdqg5GpfUudBKY6FHoBv7ante+S9
XiQ5xodRoWD3VrerdX7G18aN0qCEROAFz5fjM70EwZCkC9Jrnswu+Dt5/54tAAt5
/k7T6DsvFtnbgz6mqXT6GlZqhi25isBaNAEQW9vtNfPAAJA6IQn0HGFbBrtJxezV
2mMRNdZY+O8KeFDDJv29Bo+sYt2HiD9nGUGP+K1LtzrQj9AviDFurNGaCPGwcW+X
g+1sgLv9f4LFILAIaAwbYETsp1rdyRR9ina66iP4IMxsKuk7vN0BWjPBQjiRtSey
3sDCs7SL/MwwslSq3hqsljhEXKgpW9bVGcBYIiB9Nta/E1NjUxzsrUlBk4ATN6uc
/93l+VG31xzhLwJhhdAbnNMolHrLodHSCuEpGgzUjco5z9idFeU4RQ5U/GNNY7cI
dZY0izWjiJYxt4lrrvjfv2Y4Rk+DUDlyWo8XcibwHtHgTSlijVJ5HXO4pLQ/SUKK
aZd0TdQeaoQDfQfXAqj7KYh9/+dGTlgW5LsfT+h6rqvRgn9cirlUWAjjtUKwHk2I
GmfYjSGAeUuuAvxyLeWVGsZ83UeEauYm/kWNZ7aTHPXs9F1AoGCZj3fj1AOy+nzT
4wEVMgXrmwjmugjvQcHqM4GEk/HsnjJEx3Ifa2W2lVBZarLFR5eTvSJSiewN0vw2
dwCjeyXPNP0+fJWmXp/8F0PCyXBseCLUMV8YAoTP1UozJQzQO5mR0aqycoBoqQac
YtP2usSub1n044BxN9OOS6vRMQRHhAYAnPj3j8R+5WKE8XqQFDbDG7D6U+tpmtZ7
lVwOKgv2ni+oklMj959BQOTabnXbyqMiSl7JUXXHkdZ3D/kyK+DgDy4+yMOBvh1v
YZoJKjzGFGc0RjJcUbmAkXto1zqLaX0soHb8pjCNEkcwkfq6l9JALfCYsaBj/6XS
sfc3cJBgNj7NBmLBZXnMHGL1UYB3WRuiAX25BMFbr0rJrEMKcnPpgje0ivZWB/O5
pOWVsqW0nIQcWnH0BDW0udANycIU+BkHr8sOntZdKCqX0nlaS7UFsYu5r1oPpVBm
0KK+mBMwp5RR2UmuOP6iPpa4UlfX+gzsOOnoE7H5BnnaLILinC2UIoYMKCvKdzuF
/5XqP1om+d39tOrsgHCAi83hr3LuK7QmDcbOFMfMkE29mbU+LogAQV7YtZk1bhCw
W7uyqz9U5XfX6REgvTjKXHClxC7bpfYKes21S6iQupQ1LfufD3DRmwfAhFxhYGJe
CxzKQTc7d+CZgHnQlleCEMfPQpS03HG4dBkizvCxquokQxr/YITCzBNxP+/XVAz/
UjD6883iSKVbw3em/O9GZGxxG38YU+EmyGVCAL2l2/3SDJIcmO1cOHvT/JzIN7kJ
hIhNEjImjILRXRl6gLd/9ZMLQzW24XHxaJMNteNmBIGqn7ypDK1UYwigsp3Jy4B6
dgLXxZ8hnEMF7jmy70hxSaxP06crlUFkLvpudWlS6JE2lXiR3vqC8NLWqkDgap3A
/XyBsYk+6NLPi5HtRetBcEgXrp/2hsBpa4eIkUiIsBceirYwkJVVskd3s2zH47Nc
xg6SUC/0/DGdCmVftvH+YDwwNTVbWvgcm2WVZXhaNh8xVHADAQPgyC37Ri1QTgbm
9Swu6zbuNnp2UK2LUO79ufi2gMN2APKoSDMQB/A5OL0iNQeQOjqZqYLpFrbYieUu
nTH0vZ2Ebuh0TnKkm98ZwQ7/nhRlWd4qbXEDsdwf3xbd4K/9gnaTdEXZBKGnvzdz
4aKZHXZjDkNHpYcIYPU+uCXKyKdhMprDJTKrzMh1HxyMvL0iXvV0UCwFTJqf3Yb0
j+2DtSC54KDk49WAo8x7/4wv3fRbvBDtc4hNL+XbX2Zu+R1siwaxNYJx1aH4gKaH
I8GLQKK0R3an7/xhvpbASYjlsxGEIC18oxNg98A3ivSz2cMiZ9TXSXHMoaX8o52m
tZVu5A17PrMAEBNdMbvqC/D0bNPNJYID2zKoEgVD+IOt7/jUWyquJL3EGRKz9NMf
xqYwAblc8dRZfMFdcFYdVXRcpuCBSz90yBPp7LwpdqD3ZVUsDh/2Y1I2ZsxyU1uO
Z/SoxNxCiARXzgitJzTIqU2ODvhMPUIXloJqBmev0TvobgyBU1iV42WehnmqeExk
yD7ULKYRDWsHDjlXugnjgs1l/wzEShg8C4uaYwkEnP8xB1M6X4FkEVZUqSFS9GvI
0l3ngL22XjH81n35POIxnRa9uhR3Ef+TIPN3SVe3nXvAQcRYcz1ljPS2DIXXum9K
gBddOFOkUUmplMBsRJDKIFm4eFLl8ZIOKHb38rbP0iKemXGVL+nTutPPgKiZbDdM
UStDu57GaTp+TBK20eEidevOJTXJ3hcWJdbwr71UWZsWVxg+pD5Bh+D5/rk5F3gs
/VU8v3plGrn27yQ98jUyy9iYIRO3eJ6dXWyL3zvGIC8Kmv9tWfn3bie9ur4wQK5F
UGnIg3vKH8LI9MbYvFnbNMr17puCfzUxent71U5jgUhKYMLhQu0jEx+EmKdWhxEp
pDiKv4TCRgIZu0duwkzrgR1fX98Abi0nXG1phx32bk0ULWqW/M8ytIiHml+SlhBh
iso3CP+aMM7qFaBYj4HhWthO2wNtvnLDSxTL3eOL99ARMhQhBvAANhXGv0SJSwqF
ChBZk7sUFX3nrTcT/h82BYZFw2qiVoQKs29MeQ5I4C0pDalVRVi0nkC0mUh9Ru4M
+cDhAdiL8Tsi+tiCjfw1zHMfPiY6pnZVcLXQzMqOnAQinMf9hVKU7ffXqi4Zp1BC
bblT0w7B53mGUEIsW4nagD52Uo048pUGDwG0jOIAC2qUPtBIw8BZYynrtwqgsVbo
FPOc1ZshkGtupjV3bwQsrjR6J49Augi0WmjM+nrI1yH0AKxFTHpFv5INggn3ls0Y
NtQSKratoWkaam7/B3kfgQZNsO8qCrVEXKL7pmeCisye7fn3wD1CVidht9suMoqF
y+E75XnHcqL0k7xDWAFHxeFGeW6IguDKRL7MoUqvSY8ijokfAfCisVZNjv1E25AW
AGx2Gg/bRX91Ymv+JCplD8vCmqM4OLSfGkBd6TwPZbNqXIk+RdwWxWm9xnXPCAC1
+3icnkimbGytcF9uWv7MppR3fuQmszQdeLp72WARANrSbKsoTEtyrTq7YUDMzkr8
7vIm4KR+m+3OK0V9Mr91cZWc628KTAl6kVC8qc2GGzaqzfwH47MgGd1dNOhXYWGp
43+pICx9vO0rlx2vcnSw5PjhO7JLS7Lt5cKIco4Fvf0f14vKfpLBN/SALDysckTO
nfed7NtEIgkcPLaNYIJt4OJMR1jaMMUZ1t5vCPRPdtBdopGIYuLWdha5fgqVd7K1
d2YXJKEVklxTY+FaEP5PG8a8cM429F50vtJJtX9A+hjkIdLEwRh2czxfo5vvDtxZ
rN7Bit9H65BaJlbYerbylI/NHDzo6vPBYVHtTlljQ/noPXHDmBZq8To4MZVburPL
WQJy9nWDlUDmvyLT3O7d5rwYO+SgNYDBf7kle5Ck7OKnOYSnglqOZqCCT31QzMwq
HFsBXi3IOM33JqyjdYoeaUVol1FIOgzZFHHRVM+bNQz0J36ENKKbBCsg5ukj5Rko
t+yY5CokO8GrvaEn0qd7S0k7ai5iMe/ImA4BxgkRljXzf50AwmIxKcfEAdGZxUDZ
CgwLkaKV2QDmpDtrYtqVpJEY+bSNa1NxDTMyPfTsBrUF4j314GxbLFJlk1PdXku2
TphgT6CEtUs4C0mIwoUBY2CEVZhwpI7Xctxm19l90gBgJXg8MwDCtg3cyZvyWChW
dWoLaRTATIhz73/lMVvIJBYjvQgfbb+/hsXgEoBML5kkJ+ZtdcNJjr1r1e4IPwuF
E5QrzLjMr8bEquskFGU/ZFiuY/zq1Cg3x5soUlyQPRsQcYAHJK2pW3J7I5/zQWvr
WFyjCZ+/sJU146RoMJStUeC/QdPlQgFThUAEAxa3MjPMAWMRxM7h20k38tWUg/+D
+cEVXNWxkIdIMx168b9qWevDt5Rcu/Xa22AA6nKHapXcjjFT/oZLEf94ozO5mhCv
bZ0v8H7lY2fzO6CZuGu3mAC8nf58seeoKfPYfwGmZyzPShuGLAYwhmnpkuWJRcOp
wI9NcoAOXNd3QEDcm9yHNJyCzL2iq55GHKHFDhZ6QMoHsNOmjYPHTV/28UoQEEBV
ngh9Vck1Dh/AI5rRbBxkOaxCM/PNY/Q5ZE6NTbnyB8YsykA/7COZ0v2xhxiQBLTV
owC5hS7to5EXbADGAbTAhhgC73pWXcKwyMpaQzy2mwmt2yJ2Il7bs7wVXTE3EpMg
bZDXK8Dgp/thNkGw3phJsO18S4gixOKLTDduty1P4tIGnsEfTYB+Qp3hQUc9PV0f
Uv1t9SLg3WRuKP1Qv0B9p7A/NJKwgUG7X58qknrYCmQYL+QRFatB/TMk8PBuASu/
f5UlDZyWlPIZ+7HehEvSO3QnP3Xre6ncmtPmIuY9IHMbT+XtL4qK9gX1d+ODIHZI
f+oCq1fJq6ovwJC+vhK9u5inHHvPR5DbgDLVq+IqooQ4P2jl6s8jyFCj56eixcyL
SGos/Xh0vvcjnTbSA31JWpWCbKSm0xI9bfnCu+XA7lzYn8xrIHhH1DICK5tf9WRk
75QW1OCZgEP5azqPLqfCde4bnlMFYWZlrpe7Z6YqUiptOAJfv9Mb3hKo0mOhPayL
vGHQ0w/A77U8mfVKoVIJ+qNfal9oPMvuL1HBXWjYQoo9ZdOmL0AuYxLylZDrW6uM
qFUu0tXP7/stHmhfDIvHOrTlSZHTSiBwbMYiS1DK7tTDVR9/anmq7vPlac9Y52nX
9HpwmuKALrVBGRgIeJbPx7kaYVYS6nrGBlq3eJczV1rJPhVwRgrVV6JoANyfij9X
J26mB49e0mRkYhRzZueM84g3goz5ig6Xfebt2Q+uS4HXbmOnAOroc9DVoE4qGz4E
786igxuVKX8ruSXWOJSLNj0qV6HV/7OLBbgk8oru8bbmT3Hk8wixrdZ6MW8VoefT
76X06WYtei9bPIKbH7PdMtMhWGjMWYwN9SNY6izyTANsFa+dUuJ6WKXLXsy7lY9n
HI+mfC8qWRdOYMCIjuzLMDTQlvy+6fuor1rEqAwI0eQpg54KpBYc2Kdzg58ZVDlP
2NhL6JtTgbfBsxRSUqE/W/ZpATQpZaT4SFE6MVY9eYhDrLU68nEFUE6sAn3a9jW3
KJkxQMWLCVNL0LAQ+eyMhqhIrGtcgJZa+Ds0X4WkzcPeCJ8cQ0mATTQuhG8YHRm2
FHUHS/gZWqlbpr4Z52Gs4pxdUrEIW6s7MaIZoYxvsbyb5I9KksCer0XAeEQ3VyjE
DEUq/j7MmEJka0fjxrP5RCR1HD2OP+mUkELvxfHBnwc/Gej5Jj+CvRA5DoxtRChW
sxCLu8WaEJZu6SZuzan8d8o9JXnM/BL7EPQl3dEfaoI165l0OhuQxupwDZnRpMIV
Hj8j5TiVwxlmXSRTATfY85Ca9n/ERCnT+aDqD4fn+LIQhIW70DNkjOt1zTYStRVx
Bq5/0xtWFe+hyggXvWzlojxsIbwknaLDl34q8BWdKhJlmHU1fklfiTng7v3Kqqcf
mA4frcVSVquZBpif9uh0YJWASoFxADA10sdXKlEmi/PeAWNPb6ED5mjXylt+c3NO
xYAQ1dOscMbnVJvGyWianeVxFRV2Z+Mnuism+rd4fsnAkVm3uI7NH/372VUqYWt2
MCmeD2rgVSSI6zhLY6Ez+sR2CfhkiWSY0vUiYrT59nN2BJPbuFWwq7NIhnxQTuDa
mCU2q54Mw6mPc026Ru4QuBoq59+Kbvh1y4vs39nmFpT4jyekhadkH8iXhzcMquGP
pZRHZj+3MQFBujturARDA1iMni61mNuNo6HBOXsJRb27spU+UU/kcf0tHFG9CwMH
PWWjwT+hTP37cC/2cTMYQT9wzI9A+z7JPaPnoJdhpJKeoGuREV4bEhk5ZT9RdXya
LXVgK/UZf+lLOBT2Kh79am1yFmyugMIa5u+YCYQl8aLdw/tqQH83nER9Q2RAmF4I
08DC/nnQYw8qZtq0W3IPzWbdVeed9eoDjlOtdjo2hOsX2rq/cMKX0XMBZb1LP+wU
xzmGDgFVKC9TY5NqQXRetJi9IvugMxerRCcdmnBIFTJWA+qkbB8Uxk42l97xPpiY
xafg7ypQEAnJ5SDQ9admbVaI9732N68eKtXcxtxdc372Hs4/q92E8KRnHo4DqcWM
Mh7twKXYDzOqGwSNAxCYN42CHa+7VV6jaT+bs7ADDKtqCFLvDB+wxsuSIDW0F5jO
K6SSsbc/Qs63jn+EEs6ZP2kxXgYMwrDF9z5CLwymHu2Jr78igXkk1gJOOe0KOtNn
0It4wuwhYmNew4a/15B+nwOPsawILia0vmkArvQMXQsyCCECTvt6OJJNO7fDqHnF
WzL1u7SNIbLnk3cR1VN2CTlMMZ1chrObQhYCSU8yisw6FqzfEaaMPe93B/xztQtO
E6PRLv7Tidj/iA9KMZGMcgezmtM0uJzR5NExZUqm6qo8xcgw47+wfZKAVjLXgd2v
rg47+7biW2xrKIauK4h2dKpg28xCPe4Vgh/AWc+4KeHGNDIhtsvomvcE3dRxtvRy
lzDFHx7JGpNvyG0MHg+SOW9TaZdzNMObYs1+vA08YuU02a1HQ78WiqlpUVElRGhy
ue8Ql6BSiyiB053693TIL74am+Gw5gazl1VX0wL07BqiBnvgnBiaNM4FyDZd8gxx
6AOUB202j0yQ0A1vq3/GPrs65NHYmcSBUeM3g+ixwld45JkLxUVTzO6Zxd8rvwM1
mpBMIrQvudTxU4DuVORMZsI4d7PHEjsfHA4drThmd+HpyVGdKLE9sKW2lcfAPNvF
OUyrlqwRvai9mflmXGQ6caVdeAJfmhQzyE3ZhUS3e4ckk02f4i3xJ7mgNW+hKZ9W
wNvhpk2I1649j60aPvmP2RKhWdA/pMg0eVLjFr/q0UzPaKNvfbcS7VDJ9jJScXx6
Z63SWg2foxRCTbR4+0qcAqQK2DHLWUsvy1F4WUTxh6sdxKIfxFFdkPnOWMitvJ1X
0JNSXlFD/lQFCV0h46JzqoqM28N+fyRzbdikQTHW2MeUiH4yvLi3JnfuDCA7q9AB
qlLDE5DSMdFdTJnlDc/r62SzgmYnhcWWmhGi6dp8/S9HxQ1svbobot3IkOq5u6Em
x7k4+4uPhU9nl1nsm5IhLc3b2Hd14gBZe/TcfSsa0jndJDZB2uqlh9y45Dl3MH0B
bhxRH3oq7YX28moAjp1EdxTER4TZoQ/8Fm9Fl1AiNDC3uYyNJcS2L/V+47ze82V4
P1iTveab2NuUHHHIKdEQUVib7GqcoDhmAw/3gDd8otlF8wffGQYwtNrBfgxbjR8p
hBkkyyTR339bBf1g92aqB1B6IO7DH74u2zSxONCrUkVFzm0IcF1iBoqmIFwv8PZ/
Sp4GGaaf71eXUdODviMJ04f0Dia8/rTJrfDqxNVao8L+0sCP4aDqTfamAdwXi7rF
HD7z4cLbIzlaKWvNtB5FXfMzB08PXUngA9VhEG1S6SYGuq4WX7suUOhBLBK1V+8K
yiIfRu7reCsKE0xsHCRRkZ4NHRtbBoldmL0nECxAPnGpRGEWNejej0ikVKCoygg4
9nXCZBMeH7Isx229aaAIXJJK9WSgCkFqiEWSnw5/FsNzGAwVInK7XLfiC7AJ7xK8
rLi3eTZ5rb+cMb4UfKtaGF0oKcUDYWH5BmwV0iyuWe4T+PHI7whsKP0XUy50SnVs
DL9VUDHQhMozI3JwJOmzOwkdyvvEO/kNNdAGiOPRiRXob6tAali7aFkdnp7yjGjS
ekrtP5KFKOp/EHlOppVKr7RkXxy+DAO9QX8i5lfguz8S1yoJjCtN+PP1NSrpM6ej
GKtqYzbCxNxggpgMoTZ4AUO6LXWPGBf/zjpUgMc33qKuHSYCuudzmAARr1Fo9k1j
t0Ks4/AgwvQqcY8/VTb5Q8tGoSbxUaQmEZNL5uNmuOzGwwMSOuuv9NyUImLb1fye
q02IaZxpm0ivUvsqqOqXpZC1V3Zr6PnWQ+1hCvv44l3Qsl2sHxYqSEkUi8HuaUP9
Ay25WwjYQ03kebz2d8Ka0FTZsyBkHg7b6KE24klmJUsvynXoifYaFpnLv0IzK5wa
Mj1ltkM9LYFAnRgJEaLYqUuLJqqR+SWQYdMORPggVsnVICKmWg+aVThi0xb2yUve
dlW0JTiJcNWN89MbriqXy9VtUkxMs8IX1rvCemdbdBv5+rY+m9zR0NSZkqoc6m0i
AuMFaKVoLUOYwb599Qt69khFTMAM62DqnnTOGlsw0SfAoxSt7G5XaoDOIyuRSs/G
nQjBym6yLkRNozbASjOC4dTvviKatmVsO6VmsZZXwIH46GD5kbOq6tmNIJAhadso
IlSAyZDloHvbQnu3H8B81UshZHtUXHwiuCvbGBqATP6OedlB/zQ2T7z3Ktpom0mu
s4CXiT0PFpRwLluwiobWCftK1jMu6r+b6pXerSxnLC9JOpvfoSmC7U5CxMWyV31s
sAu36W41cDMrqdP2BP0WFz6snyMHgSxX+eZa3aG5AvP9Q3kHVPq0/woS0Pfru2EN
e0F6lppDIP8yGsU20c0wagkzWVZI6oOMGGu33ER/v3qp9EM5vYiO+7EOMJxzyyYB
YKo6tVasvxqhn1aAqt0HPIE83/R03NQ7VFBrV312AHX5zdguhdHqDHVJVO3GkC9/
lb/A+kX0v/Wt0moR2dsWHC9Hp+k50eHO5p0cxlXvOMg6f/aemORj8S+cr3BfMqTq
9Z3Vmam3RMyBs5ztdYi4hg3Ec/1gGUnoXBIS1UQFqigocqv/MAGujmCiyxowqiyk
yiJJqjC3PToJv7Q77CmLZL4e4AsiYoMr2nV7+I9ePrFroS8mb1255cnEmjLSa9lO
x0PeTCcyfPkqreWDQmxM+dmwdQ6l9pb+PhMy3YwFjydqPPCaqN0146hG1KwMWNDm
neO8ukdX14tZ8MzbKpCW3Cc46fgUnvSwf7ykVm73UAEIeDGpykq1AeL2vTWXpFQg
n9voX1ooiyqFoTeXZgLUhQ7PPNIZiwAWuc7JccT1yqK1gB6feL2Swvb9zq03X6MU
Ma+ZSgell2g4CuSFGh19wa8K4HFDKc9J6Fclow1aI0zyOefLJ3Cml1FrSnw9lp83
PSivgh4HHQdoiu6+bnd7/mVD//ho9czA5Q3Y9PEJAMH2QXbHFg+NIGmU2+tGfJKp
/kf3v7NAxi/A1rnZx7c9v+7qo6WOfRA7l3djHZvRD0ljfrRSWk8Z+ufNvHb46Jrd
NxVs6bAzUBRsti4lm5zJKPOnxqM9FBeCo6oWt4696Pb3MvKG4dQwXmYjpP7zD9cF
j6bwEF3NZyBWxROhDCpRoU6gQ1vb4fViym3Q7mdyJ6wQfz28KG4mBMzr6utFX7Qj
qFf6utSlULt8sZA6I6NmvdZkVBkkzPeY1q3tMCkex+BpPNtkkaMGZyoksqXfpJzm
hrCWdoJtEPDzmjKVxuyfpy8SqZpXgOc3V1g9x9ro+4gg16QlC9NDfxNlMTNzDxXj
xFIc8tlJAMj9swxAvmE63ZTT3H9JKFsV6DHbLqsSfEL+iwytDPTGewLGRlqzMzy3
AS8zMzxhX/2MTM9s7SsCIOmas4Bzw78llVDxWjBtoXV8+yHRau9T185WjSmAIZE6
RhJ/Gsn4j7AJVyCnq98s5NUA+uo0r4QQXzY+WkeyJhdiLESQN68xhr+rKBKx34xo
xLWA2WLsYsB4lVWsbN6I9YKmTbzMAvUh9NiOcFOx1h2MGtcYBgwEYhbZVsZgMIYU
tHGFl8xPSSv8kuy9iom425paz/vP2+ngskWQg+QuGTMKgv0r9VGNxL4hLxp4ItjY
hgWo/jDWLFxdUekRjl6gD9wXzF7KaLd0KO+Uq9ubcVY1PzpTVptyDFv7Pkj5Yr0A
PnvAmLJtp+z/NcE2Qom2YBzai2SbSR41j3H0KL/0wSgyK8kwLTbozxUQZFLL8AS7
wJFR5c6mOkRoW8qNmwEffHkLsefx6H+82R8Zg3j57ixC+QPyQnPF21YksO2mDLC+
6uHUeuNBaoGxebyY0xC8fxDF3O5XDaK1NOCm1ieZixloygcYwGqbkRgMRrNUm0Fc
nTOc+iloXbxkP22pbqBDnpsXcsS3hvTat5yf66zHeMt7cfUonFt70j6sjxOTEyl6
3tK5d64URuSFaLbd4mUppRZrJdsPEDsa5dLxI2OAI71veLYg16omn3TsoX6EoQI6
M79+TyUrGXmIIm8Tv4acRLOoYyC3Dr2kXs1HLvfWoBDVdQf7Js8zFlshbC8gDFjM
m7bbctPYgygN6NX6IP+w96eSrx8e22h601pv/gc7+e0rwo+w6kcmndrvAzJgf9ra
sBaGUdwleTPD396zMORAyT/cCbbZkTgy4llGa+Xl1NXCkPlmi8BQUvOLsxrjC2Yi
MiFrDxb4iRJB3w/yLZdzQsJmrv+2I38Fc/WYEPDaVnegHP0Lz/suZUyQf+s2geUH
HxjIUFt57rY9W4UzH56N7MXd/HkclOfZuE+KU14n7YFVQgosMpB2Ry8e6+F33aAY
p3t2Sy4PEsGqk1Cw+WzH8FOoUhDjJy/pyW2fzqXfVGk/jPyFENz8/CYyZRaFQppI
qVRz5d/yJHmL0XozxIfdrt1d8Kru5/p4oksCjk/z8kyXJwVc6KdDmT2952PzLfxV
sRkyKlxDcKc4V8+2rcvC5xX/wIYianAdWclm2BccCg/rOYAwnqUi2Uo3ul9jGWpO
FewRSi7ijA9Ic07YVD0NvlyTJAx9pwA7htI9bC68W+IEyOOrKDmEFAOLmhWBXnLK
WftLOVPn3qD5br77qyyRvuHYaXYCkt1DC43BcTS44QgXvqsA18WFLBIjMppYnIs1
VJHFknZRpvMUPZ8vUhlp/Kj9nmCT9yg4zfpIyB1NJjAGeI1fwX5gEN3j3Vaz9wWb
s5wcLMJiVaOO2qcTGBpM9s55eJEqax9ybpu7IyEZuul9bR8wsUtAKw1R1X0JPT5B
g1wvqEaXw8aKhcTUYwVGI5FSCT6EA5dXVKU2Q8yUquJPeP8iFsnrvk7QCw8yzd4j
yxpeV5p0Se0A2lQqvk+0wYqfJFD3zrtkovp2XRNXx2yiG+FMlMZano8FHQS43h99
RiMSMm9Cb6mdWFWsX4Ht4ZXWzJlLhTcTl9n/Y9383oOaAkV/MsfFn8Qu0pXTfthQ
R+/AaoKwqxUtmyzkcg7UGMc7h6mgEJsjSItBa/xt+RylrJquc1JqNI2Fn/8W1rHX
7Yz3439yrnKjFU91EdCuKeY9fV/sXaFUp1QiL1npstOdLrtK033TbZVjg/MPi8c2
YdQliJLQgdUzzv6irHnDs9j8IP26p0j1VU4DYXaq1naiGw/JWB8yb1fpLwE8l8Pf
rX+oMtwuHETL1KCn1uoDevhprx72YBtLTVjB/gy/y+z+75FSB7h5rF2PZ2ZAyDyv
eutmgchuwfPvsn7AlZzfMM7bqCfPEYLfCMTvthK1kzQgVw4ess1KFhU9vqfxvjj2
RPH9KX9g4mX2XrdV1NI86OeQLLNEn6Y95lCTEYL99H5uS9tLJDRjkzGzdC90clYy
X/WVWjbOEGFRCHvbiSe/Q+xHWJbbbRj2tC1UlRKrwZd4pQWOmLWRHHkHlkldbqAF
cGZLp+wEquXWANqmYQUZGenHuogr/sCs0iwe/iXccB0+HYrxH6KWlO0YFfHmif38
OJ17Ji+EswK8s3/Vw/sgpSsaARWSkQNE5+KTQCabUQt9Kql7Wj0T6MSuurMMa6wK
7ByNTzEOljJ6YMTkAqaIQFDA/kmo8qvDeH7T6Pu2+5j1LRVKyh+WD9Ip9zFPhlvO
cCVL8uhRDJAu3RdJRxacYnAecONckBvemRZ2juDA2zUZQ6tb146qmKVHsgIljrls
CLTAkCIS6AxKpdbq1zZS8ZtgSe/P/exSd8im/WkSQvGgB15zR1LA0TMvOR6efSJB
eQLwy9QbWSVhNtAxgurjeSbRd+7mXjZh4TtJ7Fc6lBs2fOdqFvoHbPJqP0C65jxS
yu59Mu7y8eT1ZlVAh8PVWLGj6ejMby3vIin+2pew7y+5uw3xOsGJqyOjlMVxWj2J
YdfxqZySfLK/sUuyx5tWM9qfS8xb1n0e2Iu4hfSNTbh4xq+LDt6iaDAwqICj+nti
uL7NEGHyM7uNXmWz3d+K78gzTYYE3LH60uSFDLz79bF5hKdElNB/zWLbGererYU4
Wt6FVHES/jPxJtdph8U6tfr+aXkYg6JXxqxXdsiC75wbLmdD9qDQTaxpL0XI3jtA
YdlgudqNC8NUfNHr3+lELaBH+XMfp5R6pfQbhE0fvrVjnwVx5a1m2ZTWjgmIL1nP
l4vYruLTOuIngeNYfZhHjyHUm6puv0fwfcWdx77+Cwp7fZqnxWHQdsUvGTNoFykZ
XOWiRfciAILIYc6wDdB3lKBxm/xMUyuk9UyZ6ChcaVaMeAULYHWVKZGxfy1OdqFc
PMA9aCI8B+HVvwNHru+ODZxxft7e+eGdptuwXnv88eobhmCiuUrrVKmNq7I130ih
SR1hMHiH1KwyB7F4xkRhRCjujGDl4N+0ABysLlIxMCl7D1Al+aPpziAmOaXxlXdz
h0UDup2tQnW4ufBcMwRaF4SYPKGCAIsLNhGKPNBI694Y71aK1CrdK2P9+IAqqmXX
KTKLpDkqQ4pw9wQlczZ7RoGuj8387JaowzYWhaKhnJPEnhPdf5J+ILq5LetJuHDM
KKpG/THZ9nXvrED/3MvsNmus6m0m0JglKhHsSS+QeyWmYgBM45LEhmYI0LxDxlKI
8BwI4UCXWeyEb9NV8ID5Gh9NpjdOl16vQ2Ib0En1IBvej9ZKmMIgpt2OCxZ8uYZg
DB8vNy339EZdT8og4WC1AWSDLwK5Px99RFnTFRHKEqYK8S+t4JebLsMl+uMc6M1y
9BnRlVyGh1WZiUCDb6MfYqOWqQ4k/eN+ouKGc90BAm/fGOZ7BmFtFmuCfbWvGqSh
wN1OV6EKzwGTl/iUchsNlpCSvbaF05/gRcUWuyZLbg4UggwXsJtdYvyEWFFJXoyM
rmvZ3eKZ+CTwy9AAUX1Bj2qW2w6huTIl9DAaNekGw+zNpKIUdmL9gBtM3S79bXoW
XgK58SVnTEQhdhmxwWhQzMa3ybzneovYXVi9RsK41JtHk7v3WPhZ8+hHdi4BiGYT
UXpl1g0B5PwfwUZn1fkC9GZ0raR6x95/98vLByXQzSX/NsEpfjdBUGMWKfaUzljF
7kfiUcsqFEx63wGFOuRFR4tLlGtoubub6NBIeeSzFui7JQruugmy/UFUka986hrw
NW0xnGrsZNDE2BynL9kQMwnN73/XdEBGUg1nHKByZh5nBUxVdeTqaSwR8/nJJH2A
//HwZnIgQsH1Rj8n4llgOhvudAjwbEZj9epMnbD27PrnMAK701EsKHraxCrHSV/g
QZNs/WTCI+1ehQmF7lD4v4hUC2aPyWSG9wrYjKAH/dNlySFboC28Jk5tVLys0PIK
BGAMLgSe+PWUL8MUPlkZO1gNCGPp/XT+kT/InGHa08zW0H30rvvoYHCrAgv7sKdj
P2mXvevBFEavD/tW8RSyWG/Z8LMY8lutkqHKdAU4hBvbBCxPNWej0zATHq2mzsS5
h4Yt3QfDv/RehRGv6aNdWgZdIN1btVN+PaS5ThRRs4vEPviRE/QJRST4zcOET+pb
zB7g8tnci2/QXAcOouh0C1aFNJIvFGhOELoJxeYVpJ2MTz32vwt+gt1YvGl39F4v
3E3IO/UTkkVr0vwrjIzaOrRIp2ebmXL/5uVqHOaKiE1OQUIqHO1cvUM6GhzjCFKv
JnLCdzpyoLQEVvtzmE+uFlAWqRC4bWoiwIuDirwNnCotspIpuIBbks7jlea9J+hw
zSChpnYnPCboVwEB7/5cwoK8KrnWbRDBSTVynOt4Ky0b8e36xtHDeGqdHLcfL4at
rsaIcjFyot57YgsZ7j1QSUVwMZgiUx92qAok/WgM7YTIUBPvk+5uKeAvN7Jx68ZG
7Du29529KrbN8p5A30Cu5fk6baWmXj3yfEWZ6DYrwsw4v43FQSQB1Q+eBaVXOph8
X7Pu923lG7aDvVnC3i1MJH7WQN3yCRuIJ8iLS3rWii+jvDUshBlqb2EWFy1nlP9S
lWv/ldLepkooxNHY8rxDn/6/jvabYV/tpkEG8H5lWEX3YtJxeuRygnEqz6vEw57m
cNEP2q0s++BFX/OWYsmik/mCiNaMDdxqdKG/dpP/kLWKrJZh1Jap59Yy1UUKlrgV
Kmcnm1PjlcTGS47yP/GfZkyBVdd1E9YZz9QKgKCLjd8F3jsC0OSnrRi02nyveP/I
tP3PWV5G+t3g+P35CL9DNUNtKbCyLCzhTDM1I+swmnDx5bWc4CDEoc5MBbZD2ImT
J4T+1GKyQUhi5OU+0RzIQgm8+qaPJiMYR8PII/lAWSShPO9B3S4zWBM4rP1Wy2o2
1PfIDalqYx49NhoeOShd8Ye5T2h30c1n7j+evAibayAw9k4msYN7g0ENYNOv8CLu
gOdb6e1xWXoj6nKd44sLViDBiapjidPvP4akpoxuQjz3/uuuFGUHE4zPGAJc+qRX
eumLu2vLs5hz9azmduBz1dxk1q8O1LX0aWutKVgseySkaM76yQSuzufa1QM9ycar
U6sThUseNFX/7Qtp6tYoL/9H3MFtERep+B1wQuyssUPS+VVRyWwl2fg8JqRkAg2j
7OmgekJjVGWUuAkc99mUbeXAM8wyxLBUXS0+/VM2SyGSmxwCsqjznBGfJgdieHTu
PyriACpsMwOIJKsiUkY4zWxLvc1/Y88adKjvT8NOcSXACQK+UZLBeRswekt/uudz
wIUQCvrrxdzxTPezVsU/jhAt912TuMEdrLmpgBJfkhb99PvsPW21GenTfI78UEbH
Yf/7V5A7CqzAFaiaoQinZWMFsiYMgicCSZxlhVsMtE2JwAlGFKpVp+SEII744i9D
5S+9GE14t4Ti01iCrqQN/JvPCYmrBHg0FL/IkJvMOIkEMF0w3NRb3QSdwuEmKD+h
5hOZ8FIQaIg/IND2CerNCtGmZPs5WU7aUzIAFOvFV+Nya2RS0xgMYv+2sAlqssDA
sEW885CGSxBZk3iSxGQ03KkU+xtkpsUec54JGFko7CwvhSl5lsZ9AYQv3DmnUWVV
pvdxoVaWEXgR3sPPLXUzl1oWFMDCjWmHuvnMINDr1xCGzzC8R1MA5oS9ngeiffah
1IAsdjdxM9taXpgGIUyy4AdZ7Loelbffmp45uu+M/SkdZPk+IovIp9WeCaep7UTX
ivq1nmylUKy6As/tPFZijcu0FnzwxZXPXlOw29pxQA6zCFJJvwtlqcFeuNTOi/cS
J1ff81kWCG+U4C9Si0dWdwE1vPDjg9qTxrDCtifkk0KxSeZq0p8Z1StUffQ8ssah
pTwI78RBdLVVCc9kfhAdvqUDOI8eLlqIp+uH0uOXNM0NuiMPdruTFlcImeTQJhO/
NeLL8mj0zeWjBkVwiYGIHrbsCriwxY1kt5R2sonyuaTvzshqgAngGAaJ3cs2/pHU
JfjWyIyc2c8RKrFdgXDj/Tj1+Qn23h1fkMxfA/Uk6b2H6xAWHbGLhqJSl7MDEX8l
K8Gh3Tnd/k7TmPbe9Y1vpZ58T9/jDwCm44NRZOtPgkOxwDcx/DzC/A65iVr/5+0S
IOu9/jVFITqXC07u5Sqdbr5BtD2mBEOE2SPKYdwfGmafIUCNvjy8XWeL+iP76Gs1
f0cV5ed0eqoXckJZL6iWdjxSVWczic+vQwcEqZoELsarNlMVFka3/41gSF+gwQ75
Lew3yljHzjpZvgCLFWTDD7ByL/lRZWM6BjKSiWBFmqoPGM91MIYL21Xn01qtucOa
Xg5w0M5IhRfk6KkVZqkmpR0hv3tk6KLLpb6YE4mg5lZQLezs8ZkMCNz6nmkppB6j
wvGn1mPKrmWWULvSzsX5+qtWOoqpO93HjYLzYWjwARwnAvDxDRvubALAPJQuP2vs
KkBqN5QSNir0ou1sqN7VxE7IZrOOQTQ9f6CP5cqRp6v6BIKD2GXGQ4x/O8u2tHBD
q6JW8cj+Xgc9m134RVhSFCTva6nCQ8a6L0qWBK/li9Qg1yCv1cydAFoqFgrt0tYX
IcoOdoBvms0oQpRGbb9WWch8S4g5aBumqLf4wwx3F88AIxm+sokQHzB7S8l3zhdg
8pOBdgNqECs6ox9/HbtiNScwcYkD7r2u6/9zcjpXM0tlTpvWuif28CFYZa4K7qEJ
+pQZGebEJxs614Ua1AQmwiUPe1Xy0xMP9apwBhSGaB890qIAvdQmHMKb2BnC3i6A
peBb3WpqKb/zD7tOMjhoR+VqH+7zoJoga31tM/j+w06aWVQ4NQNkfxgamQMp+gcl
Iy4D9UvINZfMMKHzwNHoV2aBgvXYGmX1gSLk9ZHTJxW95W9+zIlY8fbVrYaiA7Ju
lq+8kKeiXSCRcwVxwa21W5X39S8KamwfFk0EJIqmd2U05PkyWz+VhpquEmBrcxSo
K35SSCrzPQfg8JaGaIJutm9zBRdycoeDakfT9T8vA8qcgXEcMQzZe6p5IROG2veU
smQ8CydSonpHcwVedd2eDaVLvkUZ8Uoz4R/dLRwHTaqLs+IzpI7pDYyfzb++Mn0m
iLDkDKuhNXG85qYBxfuFxOjSKUwwcYGDjDHsStC92t4d808+gKRp8vqYV8w/SuKJ
Hyx3T0nm0IrbEXI650OFzEBD1Z1E7oGEiOvBkULaMlZ3R5/sMXoGw4HsEkP2acvS
SrtPkj09eewgQYQKssGrZTvyCHPYhs4a7Y578QpxM4TUrp17XZvFqnDL0K4Nuubg
oTV9GLc//5nnP6gGwuo3xeuHp0TyggmlgvrOSWNJq6Qc687JGP0SqGe4n62Tbsg7
LI/wvSVb1LuO6QgsOWq7lbT+hSPjM8KFD1Elb+P2WB/tt/yAb91ZQUP6k9PyK7KM
rFhpEjR69QBI8uO8qBC2i5AxB6PlE1SeWPUW+6wQ/EZ1V8PClegiOqq/bnPmYOF5
qtlxGFHNagID/96XlPLl6A5CZQty0jBrXh0K+ygVu+/oGt3g5rAlajPWlugLx/q1
MWlf7N66u6tofymzyG1GlEo/X0ws8o6RfAcfjHj6USU7HlD505hWsMFyNJylapOZ
bb2BWivGxTQonjqWMKS1lqfsG5Eo5WQNSvVtwDyq6CLgjBbNta5kU5Wd1NrR+tbJ
XlREu/tZCoZ/wgGnURkzfloUi0OK1+1CcyFYoUoiiYG7FOJsiiwtchy6S8lOvZNW
juDwH8kOEDwIajqoiDZBD472r0JuwSHD9UaHdhaFy9hvo3yHm4bIuv/awCxvtu78
Umo4DcIg8iiyrzGfBC2k3kgaP/LG6FSHLBRNrRVZBwMNI4RNtKgVhcM0IXkJGxn7
iIhjHEsd0ELz16YtK7YsGrEOfmtnchZqJYFazwNmFX7iQ+YBsmk+qRdu7FcolSLR
MsiZ6ywReeI5kbM9eKFYtwLXX1E/MpRlzBkwY4KuSklmlk2Wi4lcTGDsov72qGYF
bNWQN3Dmw3rIWUMg09yjV4UOl8cac72c/KRWNZDy3sCKOV20JkecTaLXQqutfvxO
X09c0H8xGnl1HbiXik42Ww==
`protect END_PROTECTED
