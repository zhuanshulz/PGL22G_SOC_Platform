`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YgBdwH0Zn2lgVeXCtNypmTPRB4p3wBUFWYmeBogwbWmWQNHtRf1AdroBXdydFzKU
k9IuAxrae9RdR4IJSDq0ovBLQ33d72Hwa5rbJLGwIiyDISsxz3b0lURCqevvcDPs
sMXPEF012xV1/NC5Q0WmzFLXDZigvbCnswGBfAeyaA6KfDTlpLuEwGy1npsLY7Je
Qw8g05QI/u9D2s4qvf8Q4ejEXRYnx/vWcL5dyVaf1On5h+eorKAwJXpNY0iFEbPh
/e5lb4GXk5WnKEc1dzc34FCXZ7o04M18XQq43WPe7BXj4S7f/f2Rwdhf6+5UFYGC
IqmWeain1cL97Z9zQ44m9A8lcKm7+MB2VKoujA8QMe3XR+mur+NV0Rzw/9YK9C3E
swTEKKtkfFSeArpx1U+9lDur/UleKeRJEP3Rb0k4ENpK0H0v8/AXly5YIc5fTdiA
kiwv5vXL+/IkBUSct1yE8fuCtU/Qt6HEwaRdVweF1qJjXL7Cfmn38gbJCLCC9qJq
Ug7R+Fd49RsSy/Hhe3yOH52uuiBH22w0Z3AFGbtmXgNEyzu1+pR20NnimN3kXLhT
q0fDW+xQbtKLvsthtl1kxWVtadR+D6cc4ssK8xR1WCy/jcJd36FDxlOViTdVAKOk
dH3RrIfU6bSp5KrUYCeoPymAh4RQCT/yyRV2sHJwdFPRImwZkwsc3oYqH+NJUUpU
/trEpLOOWcQfsQdubruphf3O44KIidCROhsunnRXuZmjv8lhk1zEhI8FscOFwuOJ
iKq70aSw78rUmplXUxi/Xe34PD5mN4PUZtegD+jli9VkhtfwPfL7nG7hG8wM+0nX
GwACuA9cqBTWdJlqzqRT9JqVH/UUxMcaIDDdP/FSfM2AUwMWqt2X41apa4B96SkD
N4Ore8aNkLSAMNOYv3EwhXAM4MuSLD8v/DXA9dhqfKg+aKkISaQmssHY8QQ9c7eP
IDfxf3JYwIC8DHr55PArGCvwg/jdcoqfYB5I4ewHcGKA0bQZPEFkPxQvmujYy+WX
DHcymz+h6Q2b9Ih3+eehuMAjrw45lVZP+TWyoUTXfmfz58jjXvn4aq1qoetIrLEl
lVQMToUHL+wvd0KbfP1oDn5OeB+YzB0tu0BVOMb90eSbyqYfdJjPtGOLZGOT75wa
2qoq0nQghK3ne3qnbezExwTEAgLOvW659aXoCbDLxRhSmHfRNI2ABa+QAV0mJ+HL
SJxQt4auNn316yzQS5uX8UbFBIfyPcpZbQlxXW2Hj/x8lmfw80UQW67sKMze4Cvo
60q8GYM/n+Hs0B6f17/uUE3x9mG0TUUevELj5ggZCsdH1e/IbUdePWBNsV9slxFY
2WJDP4QyRDnaEzlLnUtWKaWwhzy17mwUy/957lPlzRHYrD+QspsxBZsI5b+NHsZV
9wNHphCf1pg90XFYRKIoCv/M+iDGWYWUcrlk2kDGoOYcY61mywdEI0EbqG+uo4Tm
U+EK58DR/BozudsJbTGP8lOZbZPMwBOfyu0lJtszBhuWg2CVk4lwl/RFww9SkPHc
rYY9tZF42LhzC0Mbnt2opcjOICYeiU92WKfu0f7MuyOrT0Ah7VhR8Oag5BuURy9x
mbZCBtnYBeRHMtvsR8VeDqV6mSTHSLtuajoUUIhPFEIvnfmx9xUrnklmGnmK3c+L
zpmQYKwjy+7FH/2fMu7f8Iq6jA54lNtMpgY6gDdxpRSLlqZLF9eGnOeqVB0kpH20
iKUi+96nvOYN1Uukc7h4rz5HtOQ+SsfV9oI5+Twq5nDStahH9G2n9REWXAvqszId
nuzDoW7Rtz5RM9EOu1VHP3ZK//2K3HMTuD/7bMWTfb2jYi4TmcnGxE7tXXSnkQOp
bfKhVd64jSKjHdIN82woJkcVURliypjCTZsx0UFKcftOkvV3ut/TtAnEpiATHMFA
uoKuKzBGpqpWqPVBPxOdGa1sBEqYhyrcJk8jyiejA9o3pKy0f0A46iLPcwFUNaAJ
Tr7VwjgsBJxeqpG2CP6pwcg0hKl1728vWLjuLGBtFNJAAabX0Iv/y6b7T4i6s5op
vTrgaykqFMkUHTpAejHX4uob5RoW3/mKxA+Qz95+1ATlZbzkp45fCJHhq0QcPZW8
I70NBL33+OAL8qbLXOPQ0467iTNGs5y6EFSJFBiFercvkwvgkFNsIrbeEY5KT5y4
fmV8V0R2qjfO03ykXib2b8dqfS2MJ12e78RJnNZZpPJ+no/sGpXj/YPxx6px9CWd
c1wguVaOjsiOoQHRunMA3hHXcyb3arWEbxuktcw9e4vQN+UtsF7AEB/UiX7fKmig
nBhwiuujQwsRGzUVcjI7vHJxzt4FiTvmKCrJutMR1IIsqfy10CeY9uKa6lgb9sxo
GSGxo7Lw60Yj0DU2PO8es0elBbYQexa44UkaCN5zI4h9hU4DZWGl+HxBqz3vu6Uo
NbkXZfC+rxDWjgoALJ+ctP77ogUXEtQ4JIZs33/76JJr/P2mS9AZLDQJ5xITaswq
HL+DUUMk5OXLx3yzx5dhTcwomZgN/xywm7Q1ZeDRZ3DteYKwEEsSWw5awQVYf244
h5GJVp4iaqGIUnQSC9hPpHGoY/GKj9DfmLKUl0qPNZYlwCLgnVYCK6w2ZEmRACeE
d119N9Zbjk8PcYZmOeDd9ndAZcwQyRSq4Hhbjzb+XELLeQUHxa57OZrvEVUa3LhA
LVQgxKQSanB42OdkMUwD/T4uBKPgs5J1DsO6p/wYjnP3QOtSbMlsExMnBWQ+Nroc
FSbiSkqNE6Qr8ps6+WoYF9c5BeU468YozYb7f/TAzhRsBnnpPLWJWfyi61J7HAuO
lIg2q5OXKSuCGLWnHEYQGmlrC8QKGe7RQZN7emWXGT5bIt5r8eu6DbiItAI+z4hR
J4BlR5YOSb1O3TXhWz86pE2BU+MvFmhHM9zXTLPgDATBBKUOsMPIPD0YgGuOfr0c
Oj5DHvLSJcuktXIVHDh+0qCDKifB1dyPjhzHTSjQa7ogYMrNKm87FYrLXt5WyLMd
KVDdFh0emEHoJZ/qejv5Vy1F5zHx3lkajgyUqRiKM3VbntyfED3TEY+lyZwRcY7E
xUywBi3eNNkOjiYJ7v5oYEUOYFR5EYttbgMtdgYT0850fhklT9cY7mCHnCq7w7ZD
`protect END_PROTECTED
