`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
11wwz0eZFsvv5vBb9aZ5rAVM1O/fthlzn/BchSV+jtdV0oaZXMwSEKWTFIfdrmsI
/2mvltcX2oEAG+ycx0zVJYgPLcy9bAUtY/NCHMEtCqHFfmFucj76CZM8oQwNj8Vo
2szFue46f1m59G08AhJRI79+Uokvnv2lbPCDS58j+H9/1frltP06W+dIs4mdPiUj
g6quFVcRM8I8oCixLaencj6HBv57C5pIctf8HpMmcWGF0i3jtIWwuD7XKBFHgQrG
6HVYvmqAHtGhitMtX0DAnSnKo4Vvz24ickr6BhShDDpJZbTAMjqE6ujeX2Qng++E
PQSPO7lv9ZdWLXQJDv5m5eZXAnLlP+mJTCuqEU1yICVqec4WmtS9poVKcBm1vEpn
D99eaiWX1opVF/xhNC3LKQ/FieQzTU4LE6B9S5Q5OLUxDN+iaouUuLN2nep8Efmm
y0svYY/N2EffptWMjm7QW3wWEAdYEnfU1OVxGkK7gbBdOUvy+1EIoB5MMkYroCKc
XBPBpTzRsjAj1c94JxVv1l47HBMwdqLJ7PoZc70pOgyYr1eN8YkYDSKyNJItwgMQ
+F3aRTPZPdNbOUF6wgccdZF6I1NIW+wZ3zAdl1YHbgl2/Ecaajm7G94f9R5pyg85
3qK3CgpMFKdmk6idA1t+lLZ3N6+pvfeFJaUnpBfzBj55D3NTHbL0z02xbi3sp0dm
/NUEcSAczALJk45SHnPtfaM8xvpUBtrkFXQqAIBkChHpDKP32Xk2AjPXzx/f7U5t
WCIr8wJx+KX26gxOIoIK/tmwBy4Y+OsRuTdWoJAX3JjLnaeMciD/jNDnEFcyeN8B
eay/AAx8QSObo4y/fzk6cRtcbQHE1U59GgxTlq8BTcvJv+TFR4iZ4QADwtOYCO30
`protect END_PROTECTED
