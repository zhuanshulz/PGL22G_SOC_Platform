`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bGrTwIgaZRLHIatBwUVmLCPNJ++MnWs/fZ52cUo2sLRkWpelST5p9HS5OEFDKyxZ
nF8lCCfXE9MCrOQcb0iC4lwB6SxYyQlNAmxhbnZyx9ams4FvGSeXOcrxr0EK1I5D
f+VgDVpphQWqGfhvN4/E8SipnvUQTeVlNg825pJbElCij4VkvDcI9uhDKVT6N97I
4zlYX8Q3R2C8lwb3Hn9e7Rnk7kRxUT4FXHrpUd9P98OxQdqpQWeEFguBfvQfGUhR
AB3DwU00645WIFbNX26IPI1CVzEBUetnye1skWZ/hwaaroctF1AcbDWlePBZkROJ
IZYv6zoWW6EPxdZBGEoLJcNvfSjaMU9fh7QhLVJTOq/2Wyzbzl24jK5Y8BAOvc19
3W/AqeFazO98S2mfD+E4n4fyrvYwQplczpGzSuMfY8Qn3tE6A+tJi/m/k/rasCMq
Le/EELBHImynmvj6eNloDzedQAbre0DdXLVbcpkFAIQ8ik98/HYm7vf4C4XNrCQu
iNwsKPaW1nLhAeOfTW5XLui7xJ++5yIoh+4+vpbOj2iKb9yYjyKL3EpYlvVOQhDe
EFPy93kuu6zrPGioKquyx9RAu+f2xnXtCm3yINz18y9vGRzcXmVG+QK/zdM1fhu7
wxcY5oHg3zzxpn1RD3ccMx8b6AuYeqFq1KfXPSrRSw9fCpwhzpYdzEm5hEV+DcSY
HvBklTTf9edPJ3Hw8Znfrg+yRJCRs4YiNBOriRzvyoYRPjHB4Mjg2EhwnMAIkMBT
FhoJ3yi/0lxxiYy9r/f9uTKOKCekRjxFOZlm6LyhH1cdRtKlt5VEI1Z1djIeYZiX
ppDlJvCyXGG2N0Ps4oJ2iH9EuEkWOx6gt8q6PKmILJ/tiLSmkVk5YZVgCXBHLRnP
WoaPVgRBXvZ7luFqhGwbqgX93/CMlXWkBMJSa89W7vXVXuM51xniYxol+F7ue0Am
cNzCV9UY5bKuu5T+DH6NzD524RJzgGf+wxRzOV//2ObX8BOWwA5rVu5b69U5yOYJ
krgQYyOpjFI4ufVrS09DHXMcI10Ij2Af2FSvkbtr26GL8rzLDioHGUl64pkUEaqw
0lgvz9AQT6h2LUKZkPHOMZM5T7SuVa+PVg/5tLOENBR9f3m/rmJfoyEyDK/XpOET
SrAQZR8mxcaNG4fYmB5BPoSEIRxTMLB804Yaa+pXuhavIE6MvGFTx2KlP7sjv/Iq
Mja9CrAraPbH98nS34gc6xZ4YzszpPIWlN9fsofIkCfrZw0MMfial0oGBSWCUiKE
xl4Dvm5wCu1JLKS8DXye96EYkOHHJrCwAHKL4Kj3AxiBjhpXphQXRNWYFAOC7VU5
nycvQVq4h5iAZfVLBImz29b7/Wi5Xtgp8oRQlD9Bjx05YEbYUtJAvM0DsUOtxsri
lyiWmzfKrb+mVLcFqkbfE7Gr+0TyVHok37Wp4srcquvwnPHLw5+XU6iLSp4Rn4/B
VOndk9PzVud1a4UdrACi9CvAhViC09be9VbVHlF5D86YBMcK2h7/gCmcar/g8eJ3
/nxuLCkmZxjodykXew4HNn87PZGrDlfUG/ZbnRfQwBXo7sk+VcilkrOtaCnhzNnx
3eAUOtLMIIUwcs+CNTM+acRCUV7ZtDqBHtfKlz09j7fnR8EGV/CyC6sT78nv5RmZ
MkauUKFPkPbbr8jQJr8DAjV0Q7leDwpWR7qh5Ro3ieavRmbJqTyfqe23WKOLjpPf
uH+55PoAMpIC7CKFHiIfxHAN5qLReoeuvI3lxiob0CWDpqhDEtK9ia+tWKuyDm++
n638L6S61eqN4fkOseMC1d/mCTZp+4o44wN8MsCPGGtuunXDC2d3+UKo50wrwlzr
0u0+S8C6WxqmSriajJP+U2qPvCS07882jhu1TfTyD8K20VPlFV922skElifyoaBW
GSDkP9yGo5DGgX2ve/E3XcVLtXGt1ePevf9C14v82da4F1MQCQ8orHMAzE/QtwSK
USNSFITXleR8wC18QSXklwEh4j5BKBolQp97HzE+PeXu0C5tZG2HbEXipWJRC/bs
zL7lDm66V5ffwAOKGjHvfzKOKGC+QP6o9q0ga2pvfLRTrlN0/rpECBsNq4ZHvpKT
IgBTowPzj9BbRb429Ujc7UPy81PjWd3y9NCsZhzX/Zm9u9gEAx1i22Ssy9m/jg98
1eHUFvk8eo/JlsrAR1h/Q5s7FHDYxmjKPtVdEa1K4rBngX+OGqNxiBvWvUreijux
WGa9AL0+cFt/KuCHtYqazA==
`protect END_PROTECTED
