`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9HCgli/95G+tPVCcTL4W5zDt1BRyXqRk+gYN1iLAi8MUdGBt6taICjrpqP9h1Mtp
UuwG9YvL3zSyfCR2l9FwBS5caH7jalNwrUgd2VKoP3u35mcFiuqWqkO//vzFoJl/
igEHYPBaP0ypTRC39McDqxJESucrL3XdM7gyUyPbEuwqlYzg4Rz/elpE/lUJQ68U
q+PWISk78+HA5OjsWS6vRKsRjpjrPIpY7JJC4tdY0bIO+bdzjrZU0Bv5f5vuoPxd
GhSap0EFIZgS53eiSdNqs6hx2+adIQ8RKQQ8Rdjw2Xa9zuho+osueBBoc8Kvqmj2
khxI2otDPHHQX2QjQJmYxNf7eYK3O3kgGBkXOoptcoL8pOAz8/Wu0B+LEi4qi/pc
c959VD7i1DHe6moZAtuooI1uM0zRUDf0WzHXcO/XvthNshAL2h5GUEAX3XeuCZz9
rcwxGOJzvd73loNz3GggM9Q9rNYO4aEsJx5rpskcrpI+Tk5cc7GDXnm6Nr5gOLEQ
qHs5HQCBQScO0yJYupE8xJil02NEQ+t+USMiE1gDJGJL6LMBZUOStD0tYlWDhJWk
1d7R1H/aSBGwi9pEiKdSbs7XsJM2hRhaw1DuFi9c2io/ijbpS8X3MF9DbD1w8Alr
MQOFjkpFH9VVYIcz3lAbraDlbkCf/5S+bQQ7Nz005xYNmkyrnhjq8f25I+x2Myzr
dmShfMET6HA8NpCZ3AHej83rPMk/oQ3iNoJzos5ZiMKxIYyX2VAArPbHa37kMNPm
U8hPfvnrSpocoqfqeNqxK0XZlNs+BfmuBh4DSTjL3z09TbReDfkrsPOflJUOz5Lm
lrT4n3CHqHaRr+ePlwtzoxkuIfg1XRXnl4U82vHro9AIAqFIiLaENFJAt7sR+f55
5idE6bL1ck3nQ5ZCO1aPPZKSKNMSTBPb9TblwdBa6hpoQpN433BV1mHy0PvilyWN
2HM1YXLGtcAy87YtKp8TqdRwzRl2Cn0Gv1Q7aGYFt+ndm3x5JTmGRmudy8p0uXZi
NLsQQ9TqTkMQgxyg8dr8HgY3HBtX76S8zL6N9vqI1BgrLKCfFffhNtd5+Sbd3O2a
ldoFWmq8WPJnsLaNp6M6i+H75oAK1Ss6gt6VxbiRdM9cbLc/72JyIGTyR78qD0ZK
FaNUWup04qa2dfg+gmimM/TbSyIb2CWleTYHOht4C47FekZczkvqd1HT2fmEvGsx
wkfdNG2Lrigv9YwzLjegtOyhrahBwnSefICnn39GANwbe6g2zrFFx2UzmxcSbuNK
5GOXST5KRacc3FVgtD+pKHRQHpNbhrPibQNdVkYm6+E49TngUmQZs2YWlBiogHPA
alSXxZjue9ggfljqJ4hhLf4acS/BxRuV+9ttmv1V36zUjj8g+PqIKFfPBjTPQ0jf
+D6d7+h9M8Dv7acyAm/TM4fesjj5W6NNMpA0p6RrZ1GoBRlK1uNgVye0M7G4NKs1
AzNglPY/yEglT5BEFLX9biylL02eJlHBei9hWlmqsLMpEzRImRUQcDHCNIFZTVXs
O3gByzQrdHKAuiD/ETW8gsjGkJF73Z4RHpfnX9clXoVsD8EJLoyDLQEctdBMDiZP
6h88BKtBqIHevyXzrxTU5w4lJmW9iaxIkFHfnIatDyGYdh3ZEwKJDMFe+4OHbg65
PBDOqPh/npLs1wX+8QKrxs1eOO/zx+dCrlmaAN5VQ0bnvz73preADFHuCn9kLFZK
owqiW31kzLy1G974kKqd5wuapG04TJmrRwdP/+KuAa8UYc7gBlt90Y+BC+F84tc7
9PCk1rYS4CQ5LsSBEw70D62HVckarioqJMdVAQBX5TOWCM40I5zW1h/cdXI/QHle
UZn/bCMhTcMchnYrRVQkjepBZP93Q5CjP83LLC3ZvK1u0ujHyHy6QeWDI+scIwvV
+t6glW+SxUbTH7LATNb4l5mTtourJBdQyDfhXXQFTlDBRkekcSZvuziHuooB5UOm
j/Cn7K4C6WwPCHAPT7Il7cE25Cq83ydst/+56d4SCRgndJh/lbVnO71ofN6W7wgL
I7qojv6Pxat0IyakZyWTPTntkzMpLyeuQXIBPMAHVFvXQJes4FflP1JKhLX0oIAa
VQnw2PMFMP8NWWsP6hh2OJjgO1huUbDj1CPTTVJhaWB0J9KRfbUUCmVF7D4aNrym
ofhHhiD8czSBK6QdUw8+qIcadNseii1BSbiF1+2FKpCOq0hCzo327cyqLPPERWDN
t63v4IITzs7IAI9rvx3oZZ1m1/99UM4ywud1jssKmJieb0bdJaOP6nEhWCyj90qo
4V7WWHBZyWoWTu85IcQpmJDwYjghsnYv8JWmfWtqDBTT/bjC/STZ47C+3sVQAVSG
Xs/FsyogFuC46+ADFbAwBPCYzkTZPb+zmPfJ8eDm1Qh2B/9ouN3kkqDMoqunvITO
HKUH8eSBlSOO+Rg54EvNmxJ/amY26YUQwI0db5wU0hdiRaf7VcUHf2dUcOCIYzyy
ypmbOFqRCJ5+NwrnaNu6kA==
`protect END_PROTECTED
