`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OJPDBcBQtbZTAzyAzA+AA0rKPUjh/rCoS+T563CERD/Xbbkmc56nUVnyeJZMp9qg
inGA8SqTHlASiS4T/u4ZM1uSt/7uXizWb/dF8+KCUqiOSTmuf+QibZe3rrnGYLvd
ZxLW313EmxPqgka7b+5PvmEi1E2vwIoZeZZqI3mX3nJ1eu7Dt3mnY+nqeno8qqlp
1j2BLgJi4U3yLiGI3WCTtY65MHT0uNpU+xoMnMrwmS2LkYpKmwLKw7hACn0C0q/L
okQmUd3J4OOpeKzf071oyTOSmzg4EQRt0Pl/zoEnt0DnHU0248Qne9F4JUOUTzhv
2GZ9nkzNA3AGx7gq3T+k208q00NJg1u7OWQpZYaS5lrasVw4ZcG5G1mqMoiapVBV
saA6rDDViMiUws8fSPI5AWwkQleNJS0FpmLY/iwjXjgAR2Lp6qR+Oix6SLHER17m
a+3wqb7l8heXBSM1cX2QgCbnv5iPEub2eqtyUwr2COkGw/4AfXEK7LbgAvi14QqV
h5TQhl2kIiWCpgbTOx84yY6BtqlGIx25q/YMyYV6UhDdc4kXkTUACaVYMV56LDVg
QOvg/RqBojaOXhJwSyvjSWsFWtzl2lalqjUxngvH79R2T8KLqNUSJk6Bk3AD8XOr
`protect END_PROTECTED
