`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KvUjP3yeqAZkixqZ+nsP+5O0wPg0rW0j52xJyC94Bbpab/Shx2sWByZK5vhhUKbv
wv2Q97+VW9r7BWnF8u9B9MXLBIZZF4HDWG+OG5MrSG9qTPi8AvrChuoA7RmTMQG6
YkkmMqrE2vEmjq1JHR6CXwQLl0L5hGYV2cimdpQGyj5I3Ncm8Wj82q5HiYG9qugU
D3JHfk83tvsRWp3OGGYz1gfxG0GJNt0lgw7duW5Gh+FDRXsz/R2LS68KgdXJFG9F
ZrT82aWfDR1dc+lmnScrMoHXohcBimSwyRfayexzXY25yUJpMo2Cz+J+/n5SEjrO
tyIozfdsKnqHYQWcR9lJqS8deIOQZkE0NNuCko/CGUxeqECcUbJrV3gsZo270X0B
6/MnDdvwP4LVSV9PIUiHOv72h+J1bvYHfRdyM5tmec/CWwNkPkBBHit5qVnRe+2G
GuIhTT1f+Lfv4/ozqTx5iV3UIdYCWxRuOiYOaqQDxjmdZPXOs9hs6r8gY0y3Lyct
HvOZ0vmjJs4CbtIO32kB3Yz6Q6gFCV5mEJwmSJHBBINff3mOhoSHtUVsi1haYvMZ
`protect END_PROTECTED
