library verilog;
use verilog.vl_types.all;
entity V_ONE is
    port(
        Z               : out    vl_logic
    );
end V_ONE;
