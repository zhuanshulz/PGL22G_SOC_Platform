`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dxqf8v5n8QCLBdyZrhLMPZavQ7O0MHvE/7kB8B9VSw7bAv+EXypL68fVbj9Qa8Lb
nR/dSpCAKbP3waDjY9sYq88XscoOhLzNV75Gmm3ULihVsVii5U0ZuNpbcXFBZsEQ
cFZT7VbrOhSL3cprpkgua4Jr7tGCIsuKyb5I6h7Rj4rtQ8E/oAUHdHEBMJnOkOQl
yGvGSaGP4u2xoc96MBXFvqxJ0WUmGjB1u/KcckncqbwpbO/go40mNrG1TjjEwHv5
LiE/tVquE7GtmL70ZpAubQSrSjiBNHrztn8vgtqGOTQbq8sSzspyuTxunkpVd/Yi
Yiy6zsTG7m7r9MvZmvz4W7UGAnTU7pvIXsWupeBi8AgCeTCjKtVtDDBiwfQ76MVT
EPs6dFbsLS3xTROIcoASqn9ICiPDpUjlQNSngAWpeCSBWJVEFv9YdggE5M+w7qFW
qaO+wapHPlR0MF45dsRfQh50/NT6N5aZDfQSfZGqbGZZxCZXgPJCyvdl8MUL7Idt
2GneEIcuOZDHyvmEodRboW2T6JNtCMdAahaHxEIs1Eiw1jXELXi0vgy38Q3afaGc
fiYD4RMxFYOo/6Y8elFWEmKaTpVkak+CYAQ5tv5xqkJyG5ggEB/jBgaStpwHq9ry
cfQlv0jo+rMtUX2LnBR++U/zAmr58dASasrOp7oPooDpAMg8lNI8IKa9FKdrNJee
mQDV1BnA4XKgxdWr4dX09AksDIFd2WUT4VERAaxZroGrislO2W9CRK0OIbYfEbPR
7T5MoBdx10Ecfht59Z1pUappqDPDSPrpRu3QVvENdQByB9kCHfw6AU7zNAVLeUgP
Dr6ofgX93G1EY2C/bPr4xI3954H8Y84L2nMCdjXUKlHNeSSQCc4cdxoAgoRhSKFq
TfgVvtuQBH0svvrjsyCYR+21JvbovETUEPOMB2yIx8lADftP3ciR/tfUjaFZdxOs
CmEZXbRC+3uSH19I7/n4QIWP0fTVukr+sSZmudQMoS40Bl6mKsLIHZuGz4zwk40d
deJBpg9mv82PFmiUBnnveJFSCUJpvs7yff4XC7/BLct6ZeDwXqgalcmadpxCo01P
38A2MZxt7AiwsQQr5q7mJBPGnkjaU1FEVsSfmr3XZvCzqOlS1v0zLonNcXC1H0hd
eJdh+TYC+jk72Yg/wqL3fez7o8Tl58aid4vW04GatVaDCIK9WPrshI62mF8z/WF8
e+3yE0KSoulN3/wxmq7zFftH+POclprou1ptbj+Y5oFie5MZFpiV7zFrgq4niScW
W3oiiQ8ML/jekDAVK7emvv167e1rMP1vpXxTOZ/ZlRoGt6XGEC55zMeG3yyarkob
DOlg8sU6s9d7hlDd9kA6Iqe5MoiffhTU+VLn4GG6gUUTKSgbvY7g570BrCmzttb/
uAmW434fI3lIkiQqT4qHpYGoeUl5GISOEU4CZ2bjxQ3dAHsRtjQ26L9lsi4Ihfqq
34n/iUeDLDHt86gv7ExoEUyXTEN75cTqO30ve9vtGIGZt1Aza5ZWzwOvMgAoPuuB
ocHfKEc+ooVY/qxJwwpO91pg0wV+yNSi8b1oWH5GsQkRJUjWZiLrrCRwMfPGz/iy
tYfxe3Kiqj6Ia7L/OlJql85AGkTlqZmTur838RKV8m52u3QBFdUfMl96VWubRG65
Wv2Rg0hH9PUTc5Bzj3X/oJGT6XYjjfuKj8kn7Z6ZZ9lgORRY7KdxCKMPIJ2ZlvEV
ME1CFNaNAGSNlnCn1oEfPR5qNwbYqIkowMTWtFwYcfU73lKkeWn1rHZix/y5eR8+
AlicEEWuBqr9VQ+B7czinE7wtu3083H+JhJemc8YZlPuiTOPh9TVeoEVlIIsTql3
ET2SYOkgDJ5fi019kLtSnY5zvmHRYJBq9B31+50s07F/9UWQ3m2KpujFbbOEov4G
i+Bk7RtQu4Fhbe5pQunJaFcgHQTxvnvaFEtO+YrZtZmizqrhv0IlKfAqzZZ6/UtJ
rTzjR5B+TLV58s/fkjw0fMI8qQZFoGekG3PR0vwH+5y49iIRivPcp4XS76xJpAUe
N0f+8clcS2yv0s8J6SkMLMOVenzgX1cX347WDNwat2qTduyR+/DNEFH3ceqHUmWT
J/AFaxsm1JvQdJQ7YaKrDkgmEm6DSBUu6pQ9mwYJ+NTHLn5P/tRFGUlD5w8KHh+p
bFgN2QDxiXkP9ZoHKE6icJhl1Hre0lUeUgH3moit3ZRUUS4HyyY5aHKwRn8XL992
zd/Xqzdc8M+uio5QlIoegsKV00zAgnQ5lTJFyOnF6InrYsEJ/Q62WD9IG/sWcUBd
vFmMwkkBFQE3/DvA3q/gbm0jZuEIQBgL4lYJHMSGBwO9j616s4z3mWcVcn0XQH/y
NFnb5iShexcPjLbm/KREEJiGpZADNqya8hgvcqgYAc3fwyIG5yWu3dRe0O2kKU0w
XZ4HebJvwHHeuHNepHJ3rQum/LmrP280jIleO3o5lETsNJkRIZlvai+C9/3/xgrj
EmLVPnJEifXQBjMmRCUe6659n1iaGQt8e/ygwa6H9TGVMPiot0NoBaShXWEHnI1i
ouzDKl7o1IhOjoS2EHoWFHYgdoRnb+6pnogegbIqIMVRK/jDt/tnYypQesUBg30N
y1+74GqrUBqeNfJj1s7n8DHs5v0LIbeuF7yxTGUGBhIYIiGG+ZOW9CKJo1LMGOn6
OzXeg/vZwySFbWyHbYrqkXQ83GplzPykfhrX8VV9NiAbhCQfokPa5aPgsepw8p2y
p/VZiBeCFJAdYu/aWGaeK62bjYGta2Z7vqU/s0Eeuw3jpNHgKLWdotxqj6kZJcYi
nrhQdcTVTVtaI93xxe1zaQR0fQGdoHFxZxqffbI5xbfdk/4GJeAFqGVVsH7Q6All
6+82jlIpXkxbSrB4JdZARDHNHvFIkC+dniu9RDRFctYeJMwuiGDUSXOltxBmkedE
vI/BtYOfzuW1WllDlUbDxvTFB9GjT7W1UDnTKOi6W5vbY7ceI5nOLd4vGYqP2mwY
RIFqBemC96XNzZHvoS5W854/ABiuV2hyZqtG7ev81aECslY/mA3OGWL7EAAcOk/6
mFywE+9cK5wUysgR+SwfPe/FUj5Nfu+4AyK/rx2ofONXQEPv4mgaURl/wrZneUgD
XXkFti5HMdAB5cdt3LdhSUWul2pMeht4veIDXYrlGgQQYjrEqzWCiI/NyyuM31Pw
DNQyMg1Zcx2tAUodmf6hJJCvbdjcfPWprqD0Bs6RzNE2ezgAa8CYzCbIzElduhJj
mPYs4qdtHDsinj3OK+5GXY31bMqdkccLkSSlKpfg/vcc80HN6/cBYbICXwmTYJtT
/uYnddj0WoESGYSLepNnF8Fvs3fiPGeE1K3MPJpIhTpt72GJ5OkrkItAY4nQ65g2
pGhPKqwGhUfDIz8VSDVryCx74c7U03qN9zekP2wYYSOH8FvLVS9REalYX0gQn2gc
a0LGiOWsUGrBVMZS+kA10BhEFnmNR2OtYIOKNyQaUa8IA7DcONEaj6rfS6tNXhyq
54jFQq8ZW9e+AysRPcJonfl38gmodoR3QpJGURYaBEf1BgMXZfs4DTrQsPVAYC8P
XS/I8e08ZEg74pU8heMHOTAJxYE0p6OAhSF/Woubn7BM7I5RYJjPsvavWcVRtXdj
14eVDoJiYv6arp3cFIqnfOBGyBAnllDzBMColA/x4jQbbLHEkPm0ZzgUeEAeWNDU
2jaccx7wAO0PaySa1wYCuA==
`protect END_PROTECTED
