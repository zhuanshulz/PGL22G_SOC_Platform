`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3frgOZsYutH3a9tE3lquEj2j1OGL991uFc3UJ2Eyhw8jevFEuyO/owaOD5gGdJYy
RwXn8QFyr7KLpg5kqXZhNs9EP0lPph8si/QLb7RMAwOZUXvD2Qt2M0qCX3MrV9Ks
Z6yV2TCYrsWfolBnmFwiirVhPHSsF82JWZs1oTq3iyFhay3WzXEEty68cgGQc3cJ
dQwHG5ONmqSBwZjOwBsYFNHxSeeOJ8Rwey6OZEJPIAHafyRAfeTdiJAdcdvjHkiD
qdBGanYKtDfO/Bjgm4X5faPT8fngd9f6t+WyL4GO4fOSr5IPgyQcOPZQ6S4/TIhS
Pbw43UyWwnDOnuPZbZjpN2R+77K6ZEiMLp9m+wr6w8y9hcBlFqGtgiL/zsV1DR30
6EoJKL7sb5JAiwFN34bJAa1ip99LhCzDb3IpqXxhXPqDOzWiDhleoGAUM1kbssPK
zGBdJ4Yt3WvwNSl7RHAkr5l1dLq0tPp0tOzTDG0br++EXC40acLItjzO1M/kQ+aK
klEtc7qSu3HvPq7l1//vt3Bl2gRZJlpHgBUZMlJ1lLDVRq2tDCBeO3djzoImolkV
lk8+6XyZEWlTdBWnrGDRZgsOiqsVK4/GyxFMqaPzbjuJ+wyjG4Vm/hvbWJ2EXnnU
ZLJdy9xrdHSECrqg71Kx08SIqY95Zt89pen6XoW2rf++97p0z4c6W7vOBRDE4qXt
z4YYXvu8Y8APhU4iVV4sL028Rw6aG679taJ24GcjF6MWjn2pkumF1pHQ3GX6JeAL
z5mMCQdEiQ+5wDLZSjLTVlCl2Vbzi/OL8Fnsb+MLhJp7rnGlYCYprcuoczUWtFF7
/Juqw6L52cpgoSzZPqavt1VpgNqGC6asuu8u+fLLBYYC/+GqO/g3Slp1y8nnQlwH
86e0F9smOU+4x1qtcmTs+E9UMJeghsh8ePvg1tRByyOt1SdHFJwkLAHfMi4R1o3O
Zzk1Mxdde4WW7SVNp6+L88gs1N1vLarHAgAr8QM14S8ZwDAkAiLQl4reRovV1zxR
+Da+L/lvD9DGPOXvIyJZjyBCLgn2WTPMM8TWoHooT3j75Bfbn7QWSDWZrXAwJpwx
jjHRyJda7KBGGCZiKvxBCgsQGwJUxL9RjLGJyitlcD81Jv+KMwlUUL7FFkxsqoj6
eLzdSsB/S2FgX5sOSpfUfd2nXnqZLJ6y+wg2s0lJ3ZPnUfFJSjyKXPVHrXV/wstB
nh/eyEt+T3GdhH4rPEbGgbnaJH52ybiMByv1j9y4TkUBzS8L5xi/PWJvs+QkImns
eJUIFRu5EMQMv1obKs+VXaXQaMIdPBNxQToGqFi5qUuCnaGjYqmCcyBa9ylsjQJq
B7bzER29KJH3pkibz2U0rwBUkpbwzvm6HsAIkCD0yLR4UFFc3AVmGOk1sFfsozzS
5LZfBwQcy+i2Ri3NtDvaWeur8LAHqlBQvIN+bKd1Nj55m3KYsG4u9igeQf/QaPwX
LeR+z6qyTmbBtYy4GT1xW3sSe2owEtNftZhel0OqimKZY8VrIehru2ZMDl5Z3htk
fUOKYFEJxPXxM2grXK3INJWIJI+cW8EsR+q1jdWWEPGu4vtsG7dujVJJPPMf1xn+
wLKCVV6FetOxv7VO4O6olfxdYXOEEP4l32gPuy0GB13b0renow+OnDm9Eo7VKPwJ
+FizmIx1LbGOJbiWQHuQ+g3Due7grxse0yM/kak1jAGwtpQbRXkURR7d7rFO4aLh
+SoBsUZWkd3uu1WkFylyrQ6AC11/LRjEeMIUCzEZvhTwjbXcTvuCO/rTbCJMW83o
Nam1fctI8s9JYadCzInJPVw/IaBan9qrNxCw8Dfx1xaMw9W/H7walhxd6gCqQtjA
XmLPxPyY21idi1tFO0n2wAzkkQJmhtfcvbRrKE5NYaHvFiYvz1B4v0VhvKozTSNV
hGBxKu9T2e9zvSkhZC4hEJlCimTp1aFD0QqKf6TyKJPrFnGoknbSKW4jR84WbE94
WP8UzdKdZplmNpY+5qYTscthgBmF62iytVw+5HeKDGESED5MUGr0FmbGt+vIWKU4
tLZTrrz7g78o0NhMw2X5AWqoVZezyqlvwwPHinoSj4PFPn+eZKRnbTI3gcs3jKiq
Ni4j4k4Y6onMAwPnMfbAgdywc1kPhyQ/Cv3+a/lADGnsHei/n5IFLrBn42QBzdX3
VYgo8CLHVfTjE34pcO96BLuHwyFPQzclFGtjlLxq4rjkNGJU+8HMzGX77tlSC3zy
ISSmXNkAYoglx5TlouCQ1DR6L/I9VZR8KIqQVx6P/RwwisgaRXgfXLMvQ6azJM7M
IXH2AHC895nahRZZ0if2YxZGv4cFR7w8PG/4aDfstJCf2LQaVQrex4v1TzItM/Le
d0HrFFevxVVM1Cjwt/VL+ycYn8SlS/NVKoCjgs6hxGM1pVn7jPcU/GQ66EQWC34B
JUl1mCRX4hcEPZjBIUm1XnqO2T8SUuYgI2eUo+yeZ690n/bgRXkxq2MD95nQkxvu
THX+HHwsDXv8Mn+6Thnk2UTCS7YB5B4u6erIUtV+m5YPuXzco+U44WuaocMKGzVJ
5Q7mMUtZf4uO8S/T98wq++jOCGCBxKriWlrPeAejvqAL03uXnO1C6jWijvcGUJz9
kr0d6wkyyUCI2Sn7fSDqOSfiTamBMwYhM3YCc8iXuQ44JKAUNPlHbrumbhDaj784
+yMGTSIa6ur7o/HT5hN8YtjGTIbVGozabOUYHeBJXE4IckA6mh/kqk6hJ1MPHWj+
7Bmc5zOtumzDvUVvi/lr8ZlobtExOMnYWtFP4QXj33cquQmlfTQOCo3gUEebruro
+EOoqhZzu32ux3ggcsvSvus66TLooXeZXjmtm7M4iMlHU64o9rSqpAj+U/CH2K/n
5338NYGZq01Hn5QM2/Cfd+RL3Ik6HjLltZObhxRFgKRKQXU829d9gsZkH/tewmsS
tISy3fwI5Grt5qE5aG1I8tRncaD1XWZrWVoz+YPaMnz3WQ3s8FkeFLFcRmC4N2cG
AkTKTYAe6UbQNG8nEzxyzaj5i2YVZZNczF5/D1usiBM6NoUG8sZkeRSswqTQKoht
vSTv6juJ38XHmopy02Y2oJC8OnJTcLU17f7jQMQ6GA28fT+66ch0paaHogHqOPu3
3DMyIKWiwdixHOYD8HKkZXPw1vYUF7H2uE2e+zCcA5lx9cOQF2qLc0HW6Dcu2Mza
25iaJNXrBHg8YqG1n8GQ4Y0a8g+HToA/yyhtIMIeJ2O7e3ll/eCAbuC+85FTcXn8
IIs+5vcc0VTAhNMCCgDqLsVlKKX8CG6+5YlT+VxDKE0/x+IN4y0RAVh/HAx/pcd5
1ig2uy1h8VjQzuJ470tvmp03sl1ZH1eCXe9Ht9GgAP54dzlN00b2VWbYM5mytBD+
sc+gIfz/u6jIqZdYFhX9xeyYwbDXTsHAV4kXOEjMS0WsU0BYCw2gHiADEr509eb/
50RUq2jEBO827bdddGNlgpmv5Y1UkgBItrRy1RPMPniO6c/ijRX4USb9XCyi91jm
uO2Xq9dzbtkIduXzXXeUuzdDvOIW7KxF4DEiozI1k3fL3mC1dsXdltXLMMdNR90x
zlLsYLdbYaRKyNM55PVdMARSmg2uAVK/W23XQySefSHRqfj14qQcaiwYOMervfdW
WVwgc26i03USIT0DGnnbIu68QnG9BzDNQqxuOHymZVZzKGtS6KZpVm9QW4GhRZd0
/xjsOV5oU/xcmvkQa2wEc0n408Zet6XjjsEeY9KGcZ3HI+tok/aGSxc8VmRRjdtJ
EFA3H/BorTJdXJQGL8DIiMZFKZX0HTwIdqZSFBwhhjOZLoOAqSCPWXI2MMBiJakt
+Rxe4wYmjaEEI1LWXgWLE+z42XLOgHaZh0xcC7aeVIhykHm5Fr3Ez/c9/16tlrif
To5NPbbHrVAFNUh78LcjWmGmULBPkFrpLsSCJY13GgmtZpy2601F49LRZadWk18H
MlL4XjOKLmZCgMBwTtOcInIxjFhBVzhpr6IgcuH/3wIfIKh9d8bBJvBpcHb0yiUd
LczFo/IP04R6/koU7Mt/0xXZcpZE9kVc/9FIDOOdB1WfFg/2IKRFgnU06rxJP5uB
e4LDr4foYKAQS8WCncvJhA==
`protect END_PROTECTED
