`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ps3R6XFYnN0EfkTfzaTiq7hEOcPcYKdLc3J06MNonMWenbeEDz0oWNizBPxogNHY
pP6VcVoMjThwO90ihnfWwKBmyfhgkHIwF1gqqfWiwhk3EaiuwbVt4iZ8TXSoMIh/
yIOldBRD7MikGVb8mXGaEabep8ZQX15+d2LNcBCLrTJT+ZuLzP0nmkBFAfZhQYRF
VoilkKPqg8WJdzeFOtmN51CtxrPrDY54/EAgvCxXxH81WVTA7M1xMq9B7ooUUZQ5
ueFJt/AdfLWflHBsf2sUu/QcBXfYhrbT6uaUOa7kYF444E5kdnPr9j8f/YpRY+4H
5sHtfu1skgxqfcPWcbfawjU+bzGWuOYb3CRNloUA53n6UuQq4272GH1Ylj5q117M
IknVf6zTd9wL/SEcDzWL7U7JdyZGKilNl80BkxdEDKpr41mie30bEurzo7Sa0CbZ
1G8VCISNnh+gW5UXib0rCz+uNuHUU1oiCX22usFUWVrSENHjd/z0nfEq1agsfz9N
WRFOM0szINc+nmGyTxXgKDIph4kW/P2jN94W5U7rl9qmy2TiNg0soS80DXerXDPo
N62yWyVzp+hwKLoVxrNjhgO4jBAsT7RCniQg8ocWu3sL47RpIQi9wukDEzc48HpV
7U0e+1/kdgod7AKXOtHKNLRF0LbjveOBFJMHPyObbtoWqAV+EXL8bFgXKb6HQzLZ
ic/5kUJburj9ZXCWt2WHkpMWw/1LD7I4qa8kUIM5dBPxAbHzacj9OawEs//Bazoz
V5RyPIVibHZSQlfBy9LZDgV5lP4D2+0e5IWqgfGR2HIhz0zmR0OJ/355UW0dqeF/
fSlGrlMgqOkoufIr85SjBD7/MxLt48JX9/+ACsNNCcv4i7qbUUAQTN8BXWRSGjb4
Eag/QEpoeEInd1JLRtGQRG/UeXorKK8EF/GEcMPO6Wbydt188VSZNVU/wP7YNjxM
hoHKkLk2jr/+Me1itESOoHNFehbHsIqP6HdGYR5KusgwmGVoybSt04BVnaBcU2Pm
EzQLN0gq0AygCIvTetCdvRiglBBK6nB8QHL402CpH/syOboAdFFbcbKqR7ivOne1
LB0MpT2UgmUqkb9OVJ5iytg3TU0Ys6LvZxxf5SKb43znC5Q8qfBl+SqZwatBYg0s
H7g8iyaT0JzBHvkFaxfZ+i540O/1e/BQp6ZDHpKCKqMTTEOh0xXdswrs3sR8+k3n
aF2jL89EaozkcgnzICPAJCeDibz5h88Ef7MSgF+mT3ZfXZ0QlOv8l3YyZ6qTKuSt
O1unsermmvwPDls3t3UjJ1uUdhxK2xAdAJgmz56+lmGNYWl/mrBZibkkbIFUMzDK
ntq48BVFWqOVRvo0Ifc3JI4L9QUJM2FFCBeb5+tRQJDEEtznEr2raxqnd3rqMngO
sJdn77CoR4dZOZiir3wGGIl+Rj5CSsti6QMl4kT3FmKjS13JchyJvhtoo0mL/GZQ
XNVLYMQS2fqq2hcfvIsaNkWO0XjqeeIneufnwiOxBc/ll2y5LrD4kPXlJAv7zZ1t
LttkoqA1caBvsF+G+QFNRkiR+Kw1fN/HQUXj9zLi5c0=
`protect END_PROTECTED
