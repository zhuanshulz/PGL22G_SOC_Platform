`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6YrNJrbvQ+gVBFPWKiWmGOWG7tuchImzJkXInja0ymuzXIGE3t1Wl/airohJIwA5
jegjdlnJmmnQ5hNpVhdHcNukdrXSKQhdGum/o4u8MmN3NAg18S1iYQ08Up4oJMSh
qRyB4xmlrMp3tmzr7MpMPkqHnzJX949LcQ+jDKrMhaFEOeid7kzdvyIdoRTKT/QJ
IwHszjCMXKtitR3Pym/GbLTZd8p0emxNohmb3WP+RA42YGn4QVV4dNMnBpbKiXQp
P+HJ7jlnJDe7eCsey7S5oEWQyEox2bVTUjB2rEKBd3xNriXlKDpVH49Q25QPvtlR
vPVDEbZQMP5fwrGCMt7YyJxeQ3Rt3W6x1PppLHbaXkg=
`protect END_PROTECTED
