`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GTCu5aZCUUFHCkpBygSTNDU5c3DIxk4hSiIb1AKfsqrTMbQ9Sh1GSOOfU8yt+4jC
GHChGRnREN8psSk6m2Vxsl0fo+8Nw5/Q1Nvav0rIPBYZtpbiU6eMojdnd8HUvEfh
7u2a7EQxV8cCROaY+Xj64Hoxt5fBgadydw3kSp9vJ29VmfDA8bUr5BpiA6uW5Tt3
UqzllyYsD6RGb7d49gZlk0VqIfD8EssdtQDX9Pg1ja8sT7iGMVTgtFPPataU41X9
QuYzkUsTgc7UbgxyLdSVgk5E/CSRebXN6Wp0lGaX6SRPmUcFmc1i6Y+/hb3Ds19c
Zf7xkwxtm9mq3VfBEcM1D0oFgszW/YGW54BmQ+L1yqwQj+7iAwiXJKcafeCtrYYP
Puc01/Jdx0hMUxxJqEDzB7Gewrv9fORyfzALHTGv7LiPDlx18w2VpTnpGQAuXyrP
4rsP/QnALIODfT3W9ize5nldwQ7+L7Q1F4tWlAk464yfDfjtSRncwaT5KREIvjNY
WE9uxd0QF6yQNq5ITYedKdHTMJg/navKXN5m24hUr130zjxiipQcushAaHyOtsyK
ivqm7AOmMjA9JNMEcKPTqJEtBinkekN5D3zBv9/XMzuHFe+Rr+QZsZf3E98wuDej
XEBCxkXrGkkEoe17tnkoLrRm76buYPapcTuKkkjcsrmA4EyRxzYpz3RgqGqemyoD
FuvT6fM0uOYb0jTAM/S+Td96Er02i5fQMtl5yGJWGxBF5wxzQycNHgAzCyJqY4lQ
H/YztnP7IsSYaxsQq5li9AJJcB9FwuFaZhshvn2IuO62zOITroiCkJgmrEkDoT4L
NP5o2xeQn1/1tyemDgfyXg9GJdTMVORsHk1dp3gjx289M7VIRTaggTviNsapJcca
souMHS8/2W60UHqRw3eoViF2bnAae2KOo/bkZKe0zhbCPn9WEF5Ekd1lsRCgVUmX
6N55TbehHm2DptPTosrFV8JpQ77GQyAqFdYbkYYCC9xpiZO3t9BljMKBrCNj7YCi
1kXThjZeXNTV+xCgi5OrUhAOpYyRU1Hofk/02k7E52fVWN3MQk6uH17PVbBsxit8
6oxQ469t39v9EE6SASRzNK0/081ybGy9qCB4FJJPpu7TuRZ0pvPcSq99L+zM4MNm
dPaQv5iHjznDDMqIHcTsBQBq26Xk7qEoZy5w782ZKjY3kWOYfUZKv2nkgiEbph5M
3/5QMRC8K7lUVUG8pkoItmTadcgVdRkV0B6R7DQLq9wIlFD3HYJ8fQ1kJH3dQTT/
xbpDp5FJ/v38eOfbl95YrAz57VBjOk9hzWnku07gImLbNNjg43yQGAhvDPFCofK/
ZWiDU47BeiEwyQUJiakuRdaM3uIZEVONw0nuAhnz5CroxR1tKrQoVMDb8f+d18XW
jvbK9wreqt78A6PIvNOIKUvAb/fUT7Xpee7NF8xRCDq8aKwCO+3DAQSVWm98zas9
ADHaVjrTjhyON22RCrzf68SmbDdJmIgu9Xz1pa2DfquHSn+IY3pg8WWXwenuV6d+
2LRbXTPrKhVfnpoltI48yF7W3rny1SiX32bDDwIrlWQrMrtG4An6KRDObX3ts5dG
8fUX9VkdspVI9HXYw1PW0lmC9j15reMGDXyqQwWjnbeJsOwMawhMOOZKfDpQ4CK3
KVCs39aJ5NLSqavLnDYvtF9XfG9ownp1iArOxmpAIXNl8Rj97s1w5AZ6I2oJrHx5
8BiuEBVzwdqsJSz62iIe3dynFnAkHikpUWU4Lza0Oi+Qid9kzMPzKQEPAkJecNS6
QceCuAaMhnhdOf887T5ZbIpzVIwZII5Og6hTOf6TJLEmdv4vd6jE+wP5bstAWBKW
34u0DZahtDV2poRtvIzX/UT9OcD2lVwKDPSDSuCvhFgUTGL3F0AMzoUQYxtlXWZs
NIz2zzRjKae4msB/irbhjNtViqz8TRD/mLzhafdDEMjqOI5kqT7odmFWcl4wIx65
wa6wNJo/uW0qy/OKyK3kxgjihPyfCWcgy01iLe4PfSU8vU7yGrj0iOUAtTelufZN
kOmDEO1ikNO/vjJ/uBl0gGDnrnkdTp4I3u5o+sYjMROp+oT6T5fP3Pd07X7xIbgV
ORQUs1luZZbaox7Tbm+EUsj7VQ4z5dYaydudChS8eMOwvLO2fjVFIgTB5MCQZf/Y
TJTClG7DL+LbsCzHLnUpZAABAuAzSUNZ4fFucCyMjpQs4eLXm6/nX2wE+JPZLXHs
z1nfPDrI9VINoy1zI22ovI1bvPaq03J+Tqlw4QCxvgDPyf2FEYFZauEEgXm/p8ww
gD/b5HHEYJgSu3u14zFgib3aEAmMyzOVKn0gK0CWG+Sd3AxGATrdE5n/8nY68rhV
bPMCAJOr/vqML3rbOOq+tBPsm6/A9rIMsWKNPHVhodOwQAXyi8ACj1xrd5hPwo2/
R0MfiwqDCTwux5tEGlJOrtYTwF/Cvj1F7mHKHEjiL8j2vT/kNpTub8UIA9GPHTFD
KRABX2m6RyfeVpJy4opc7ThEGk4QZxQ4oQZgpJM6lhNK6osVrSyOLSfaRLbCHvnG
ddq6HpsDtRwQ4OGPKD/5ZGvRstjQ5mWR3+IPJEizaHNBxFYXf+MXw27e1iIl9LvP
a0Wig3erRt+7eOgJTIDk3n+FOkVvHZ1rAUNghoetlZCPTvzoLGRmXYs54QSTRDqN
ByR1rmv/hSpgm9Kl+qM/PkO+PTxERV4QwsODDF9WC2cGLpNH0GWSCGZSuf3MxGCL
R966yf2QrEE9Debu2z8xvN9xXyxiyio8TbWIAwYkUNNfno3uuo1WlrL/2aCID2UR
VoAM/WJFkLr1Sb7Bj4mmXTk+9qn/voxvDJ2BaQ8h7riam/XNnUFL8RcH9FtvIwPM
D7kipTKuN24/STKzwEkotkqR2qhGib9HzBZoRFbUrX0GmMC27GxONhDVkry/cH/D
sfECju/Z9nk7A6WJuV9noOMGw/1cJH+o9a7T3RIuZGQugOmnl/ZKByv5tUITcQOX
3pNxFiTHqhH3tGTvPtqvnbDTLeHdgRx7eXrIZsHnZAVD1G+WuTYo1q+ixjVHfYej
H15emaijkg/hAji/r6ofWY1ZMcAJ4nA8ITbKkIBAC64arq/tSan5x7GKIefRghPp
dEvYmsUECQwofPw3Lwnwh2UOlQjavyS1o46aoVvtI61UhoGhf8kEE7a3DLJc5iKm
9pTwP3uDmvgxeTIOv1b5iFHuhgCI/NoJmLEUIBzBTamU2zFl2FD93/Wfo6ciA6+S
txLyxDO0qdsjBc2z+vR/tZiPhmYPyIiibf8DwWd9wy5NUbmbTCWuxmAHLvpDxFSN
ZwMGMCbgDBtM6BwTSs5q6ieYsn4xgDPsVPyhsC65Cco/OtqPBHRegsuwY7F2LvL7
5BV/1PxpIKStmESAXd9DMOgW87YFHsmHUfVAF+K6vtTSqXY0h22V3NEHTXBxCTQt
f7t9GRbYkAYhgMME1ryZrPs4imyRfISK9hh3nkfeudZHWDAkKaiBfHB8wmmFOcXG
aQDypkrrvC2Fq2u6xHxyh01NbF8Sogoch6ihc41TCSI4szDhuMGMX4KtTrXR2Zxf
jR7qMTJlQhTX5dvW7SSKeul+muq91STathXdcsi3Q6TYHSvhIGt2zaLEEHOVBFGc
HETJCYSqGE3liGUhvXBFEDNmFzBGPIVUIz16QKj6TbOXLLVBaniPc5sUmEhfrS8v
FlQcBjhWobJpJ4zgwLlHvivORTt9zPrM5HIvaR4a0gkSv5cndo6Ikc0fIltef13F
B5kq9AqtPQ5Wbvj95s9RxU6Ac1cDcM876LeItJBXLBMTCm4FKTJ1nEUxTXM8qyn7
y0auAOmHWgRYbTxcGz5l0g3nehFWoFaMIV2d45Zxpd6d1CBMU6A6nYdYokn03Pfc
jYKOO7bgjBGtSZaCJJKjbj1AjDP3iXWkKdIAIEo2lUpEozNWBoaNV/4mUqai6W0l
c+hscfIZbVrjV1mbm9KvvIXpuTxrrMNrN+N+tYLm6lk6ya60xYO1zjS7alFSCKXB
9F1Uz0JVgLmU+9Df6YICzZ1CaoxoT81E0Y8f7Ze1hlB60xO98kCQBktGXd0yCm0R
0ZHfweubGlxsgB9p+c0a1LsK6J6jTjWSZToUnYfCu8Wyy2XHAvVJI//zTMEYQHRH
lFgVmB9K+lEeQDsVWQkb4Jt5GKNzYpEAihkwhob5ft6rPAYXUxRlRoXEMN0eUSC/
a/Q4JRPSx5k5znBwTrNqy10nfllF9yaQtym4VbDgI5LnNrwNKSyo0G90Hithy6WY
7sLZB4CjcGqTmXoAHcjpogTkkSPQUEdIstseXDC676U7VpYJv1YD3Ok6OnZRG58e
GdOsUq8WNiEVsbsOCyGY3s7G6FgceebYWQZCuIUqnWDoKRTHGQCbJu87zIpe4Ohw
Ai2NdEGX1NTQcGvQi5U1uPtaxp6W6W/RGSyBNzBYPE5c2Sx54EjCQEQQ6dPggxLY
AP3zAcBjlUMfGmlUbx/q/ySUCfaPJoav9DnY3QC0fnKbXOI12JPNGJJSINLJCK70
nN0293H32+WBA3Q8IJ2LUEEgVLSxjJ1MbTFnoT9SpOzpSeELNovPsUW0fAnEl1VT
ScwQ8+Z0cQ0gkPHpQrYgFYPAMrmacy/YICIQk7iOC+YHruHqkdpWi6PX2Df2/nP4
qjsfAwSW8SCuRu2f0ylg7Gk5CC/g1y26kb8s14e0ABmNENlZv+Ij2V9X9BcYhqvm
t5qYup0/SQKgoDeJ9rMaTnKaU0iYMxy5QK6BTnbzaV0bNvpa4l8O3K/sia3/0ZBj
0e1i23qIMFqPH2blA8c/fVGyMQLPg+c/n9h4+G9lmTmyPxMhBwL0gdSEKUQ8hxKD
UoQvWmfdaY7teIVxyJmd/WtAKOPiEZ6wK3gMlYvVGuCAfPdcB1+ySwxMl170D1Ma
HhuFyKnpn9b+A0J87xmjEbmHoio+3kxYBNzxPLrGssjk/VZzDFnmMWymUb4gI947
Z4zNg8vulQNHQP1DNTBICdBJO9u/1UUjKlQasMCCHuwDxvFkOmUT08UJaTEniexw
9U7z+AVC/Oii9Gyni610ershy/2oHlQNaQFTgFNAa7qrbXVEnQ+TguEOdTkdS5lQ
TRReWW3m+LxN24mQCRUlzxmUwuTP9CrHfyPe1o2jGzWuFBg9UP41PJZHiH9Qnu6E
ouaXJNgrZ5e8XXFSHXSSeKNOfruLrGIT9wtx83wEys7FzjLG27Ww8nCqnO7dyJUK
Od/r9Sfq7mwhAFazdGCIwo7M8zRojA0tTp5tiR17yNU+rVS/54YJMR29H/XZ1mnF
Az2TdrIe1uWAOgnK7LROm8teE5kV7wCjP4vUe2XYPoQxR5HhBF1uDudeeuOSrMS6
uBMnwFViQ3rrEo9oVSCv75EJzrWKvt5eeBSlebzSnynRRvmYxx6cCf3SXgLCX7XT
OnWBjzuW5cn66cHum0PnU+YFKNvG7hv0NHBKsHxztb5qHnU7+QrUcWXq491Nx68a
CAjEXaVfmShln4JhUjFShZL83kEtLfdtBI+MhBh6y8EjN7KnEGZ+LQ1R22iFO+vJ
QkLKGUOjfhpAqo64N2pJcDd6Zjl+6Gjsif+ODp/ctPNMihWQeFNIxHhAUF5Nk0NN
FavNtnWEeH+fBd0gYTYvRqXQanhvex7Q6YmDyNQUVxUyj1TdBPXafIXarkjrvPC4
fa3xNQjMJiqDjZF7nYY4z7+NhjOqhgpFMe+Y/qhLBT/d90gPSpAEUyhyGXI1Ok26
uiaiONhx2TKnOqPJkwSaulTIBe5LIyT6kFwRxOnoLnrXpi5VHJsdLJcuBDXj9Cn7
WtyaB05mCRP8QogkQVna+V9fn7FOlFQXtNdCCW0s5zeXVbq1vDMRzSaiuk+CZrxk
9avCBZXAxKd4Yn2OKhSmIGH7iy+I/WmP0NV/zvK2CxmEE51ubE0cl/JYL6AmZxSV
GNHETD3dKQnC9Ve9cvSYsyvz4UvV6o6RbIkkuMequQhcIu025EL+OVlApNdmFvBW
fG734RkoES1/5hjTtl4EDEVqAKhaX9YCguKPRtd08LlmLWBXbjHIncIeWePeu9cX
ETzJxfnIdznW5QxUB2uFXuEdtTlXXEdZ6axX4dJ0NfK7go0XAfSZ6kGm07iDUO+7
ebw9agEdJ6lDjqYwhRNyw115216UrJmHj6o7fiDTA9KVdH6lQXBxR7yAN1r0lqOO
taHSm1caUSYWtxgiRKsqy8RkI4ia5ea8W7z1HRruPhOqMlxmfVZx7Rb833mpWKD5
/skXIozvIbZxbC18QPVjNSjjHhDqEUssLKgRrfJelvVDCeQxb/AhLfQSjklXRya9
0ZI4Gv2PR60LhFcsf4OTSMQwdrUgNWWFqWxbxDLD6p1ciqgK2pyF7aKtXrtnzpgn
kIR4WAlIk7r2CCt4NmywNv8+o4Zoysq/FkD6UPK1YQDk2qOK7QeqDUWMX9obGQOL
EupYm3caS6LpbnESwZBMA5mHdqlallabwwQltE5ytd0Yh8SQ2eOcr7S0N7PQJSdP
DDwRud1c6s+Mc3y1go7FWvb00LgFybdpo9MaWpTD+1EaWaooK9F+rk4rDMPChOZE
GTkiR3YKXAbu+76o6IHQMv9U5l51avy4+W9+6aZDRzf66f7B1pkLi4McRrtpur1m
ZxqNDjznj1VPRpokRQ7ftDTDRm1T/HsiYBM7N6m9v/Ie0VRM9fu3BKn2HY1GRjR6
QoUAlWouVahWhsCXFjB9gBi/1w71GgOCbkXLXChUJMEWd03yTTViSnRywJcBP5q+
APABGfYp3Wx/H6sWsh4ziwui3gZ4N8RmDANZFYY/pgc/VWEx3J9JRj2xhAecflUQ
lI2hSAkWxg9TnaCParrtJ6vRQkH8WXuGc/JhQpHd6hAlMKx+UiH/WgnqGBhS3b7V
QuWXP/ewbKLYG4eAUwvvR8uGUQBFXQDqY2AXnSUKZH/nlw60DOQETlwTLPClGScC
8Wuc21NlpTTWKygzpQjku0qi9C/4V1vk8b4a4IcmavqrWHxlWUTERsu/74NN21nM
qYU6GGVH3FIQyK0/oxgRItqpPnmdLHCH4+ZgcSXrltDYpvUMSjsmuglP6vd5qAwm
9pC6YBuN5m49UUGEcy+avGFQU72G10oW15kIFHd4PUUvuNBVLGR6vZRIFDhcmy5x
wT6vIqQD/6m3G2AdTSSUCfGGoDbsto87Swc67ZZNv71NZAIUbSfV53NpzzVBSnNu
00X+6xZatZVL+G/LjaINouCh/KWXEg/mxcg/kXw082i6Pjum9Z0YoKnXlpAvhluz
l1Dy8cc8vx/U8sBhCKqBPTtSqeNoPX6WtEzC6pvQpMk4Ehg+rWGDKy6lIxOun6QI
7h4J12dr4FPcueb5xg087PMSE1ITsj6GvQPylCdbyG39khADNoprY1swx3YwRONU
5WgXGDGacPQnMY/BayOQ9wUrAHoLR2igaC3R1ppSbfs0c5HMCC+8KmntwYR8QYI2
aOg9JyqXGU0CtfRGQmPoC8sbMd8aH6qRgw2mvSYkGUXdjRPu6FXmSlcbAJm18V1G
lenZKdsuWgS4aXxnrYUtx8btZfjVFim/sTAXhtSngwQ8zAANdKZZNskblgOobsT3
b08E4W4PbCtSkiT9hICUBmWQQpgQY5CKmfH/Qi5e9r7t6gFqWZoBmOohc1JcWgYW
Gxat58EkE2fDa6LSzRPOHEvq3adzgRdxzYNVJAWgzKj+bMoj8FwUPV1UBhKQ8Aj3
MIf9MC+kklMK7J/FzQ9MyzF02+5xsPRZMHDtTS+xv3eSFCo1FVVrVMlpvOAyKReX
A7lccpUoc6CfV3HNlpbrNnGrb2/zS4DhMZ7TQfX594vINlMTyQ2PFX1GjPln70J+
vQZEkgRkw9vIEjwEwUaMXULK9qhBuX0wMXqmp/Pyr85FKNn7x6zte5xkoupN2K3b
vlLZxFp/NKRzzrxP0t5/bV/8VrdsmaKFj2ScrltNd2Z2h+yubNw2apL4/gse302t
o8Ergq0DXOMGHKZ5lhXXfde3kd0hqDk1/9p8/wp51FRUue3zhObGTvOFxP/ifL7l
9D9NCbG/fUskBJeJ0J+0FiPUpcfqp4Em5/gekuboBrPXyT8qIOvBumbfg6Jc3I9l
jwVyHFWW7ZtJWIloNFLmWX3225pkPNLO0XA5LvS+eZBg4TUom1Nt+QWtDvI3trn7
iK3ifftb4ne8NF8nKHc7tI8YYlYBAjSH3xtov/gUnqjWwQTT9PhvNGwQaAj0jr5M
JKIQDn8tDetQEXpNHtSBWt8kRmOh0doJAiiGEBEplCuXN83MOGDwmlj2o206wukK
mbTJQM8G1PGdm8t9g+gBBoYl3zP7bW6PdLkdiT9H5Lil9AlLxGQTb23U0XSIG5ZO
L3BP9K02g35kcfmHN03Cj6xVSPLthiz4sQLI9EO6jP5H9iWrmsx6zi6zaob1uxPP
EvFCd0p8mrRzNVt6TUMYW07ztGCx3zw3qSzG1gdjmvowGossuo6nwL//sTerPZhr
OlgYnfn5mrtpSaDL8RbrNWEDfDZSaNx19ygakcVdnsgjykvk1t1gUJdv/aRFpVEE
MrkzRIDkji0YvO0uI+frzzEYFM4Sib7v0UL9MkEN/kljGqY+3+cIAkQdQfWVV5sf
yEYDLdYhH9TmZL+pB5hgsKBAyDe2kVMKixiKMBTTPe+uAORXcJBcOq2m4hBkHTcd
f4umRpDioIq0DridmEiGzp95R5D3gMYVscxup0wWzpRGlKdiE/s6yiZiXFQt95Jv
r9Rff6mQuCe3miy4EZZe4wHjUkn+OZzIE+OnwOHJxboYerLpucLzWZRuZSt2556p
fI2KKiMx+qoQ7Q2lEyfy/ybzu0qBQ+pp0EACZadOUJkuCE2nAlw1roSvQHCsAvik
iPzeI3wDgmgErVA38bXAgevq3qjz9HTEjFeDdniXhKtt/K1FW9616c/Z181cMmEf
L/kuAiZG+caWgRLDLtwsNzTEJjmO/Pu5TLbyB/BxLbs1udxP6BojJMwgeLNejG9r
IP7wx6HhtyYqB25O5Mq3WoeEDaNpL/kNVZGzwDMAj+kcxn+bIZhefS9fQK79NJnk
Adt1IsAd1bHdlUCRAIabq4wCE2ylAVtQoMf2ZWhheQOPgUXKMzZ6PPHyj6HH/aol
ii9RJ1L1A5/fvXs8v6P6R8y2hrICY/Vdqpsdm5BfKYLU9VVWs6yPmSlu60UdI/7P
h8oD0Q6Llw94VS/Kg64+D+11qs9+ffYTGpJ7FHEpS2J1ow0hWldk1l7SHMuelvqL
IFc+VE9e2cMVdL9IIQDgj2QI6dU7MhqmJy1q1MJ712Y8I5F6YAXHJj0MxWNaIPEx
AC/r3pKxk9zX+Doac70UbJ74di7Dt22OdtaDERy1DCFCVbrAY2mGdEzLwIDI+mXA
v31YGO+dnqxxHiANzosDrwFsNNoaUfx1/pGlB1ob8P1saT1O7x0jtndNbp3g3XDI
kZrhvjAGufKsUrGpa8nwHueQ5NRNmWgGPp0l53lmP79QpqT6D3QSB5rrfrhD5put
N6vDRfIbW2WGHjpg3phoWzL1tdy5QEcrHSHqGtAsEulCOWedUEMICrCAROez/FkM
i4FMcz5t0kFdDxrJcnrWEw==
`protect END_PROTECTED
