`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CLTtxMLhP4ayWCxCYEKp8Pr7t6YcZD9AlWRZkMt2lYI1HTnFVAFSY+IquoQT8iqk
nKmdH0W2bhCdEtFeOO6ZoP1LD+wRqPwb2eVgx+sJ7UkaG1TVI2rjpNSnLLoFan+p
7vCNz5wr+yUqjTLRbE3ieB8Lk/TcNhIlnmD7YkVCnzbSyJOQ4rRuvbCieaHNlOMK
kJ0/wvw5DLJd3t0nfDHXdPx8+hUt/s6PwFN0o5QvuRz4JREgnvkbHBy+EhVJKg8O
1e7G6+NCOkzOgXtk0l/MQmGN04sHZXoZypgUAobP2n8Ao8TnAgAUsgUMb3iLyFrP
B5nMBlfOZ9V5WMpdGeS4CmIwieUQ7filGMnBf/l8qpI=
`protect END_PROTECTED
