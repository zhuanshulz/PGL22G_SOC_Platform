`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nfg86V8w+5Gz5h6bQfG0l/+xtxLiqVehJMxAEryHbEJ+KfhSXaVw02MELv/vaJ2K
T+MdGshQ/A7FgtJUDdDAemMmU3Boev4MMrpsDyrABc01PNx5ZAf7yYq76/nrGbrz
eDncsg67LqNlLdNdM4e1TXzze1SlC/bbgP6do8Xg7gcoiUPO6hzS5hVdNor1rDVW
DQVW6S5R6f7rHHPHgKskFpW90BseSRrYoq3ct1Y5xcxjydlgw2c8abt6Ff6fug/D
kJsswVdI1uadss5nKStso5ycMaMUe6R4JnddKDRH7KXDw//lJ+Q5rnlBy0xX60l3
yeZJLYO9ondBtbx9BvFP6L1VECb7IMArI6IFuI3n47+wNn1vnXqvS3Z9r789X93d
M18UcnjnqpEU/YSh6H2ATNBWapVuoxEXpCsuR95LWxYGD+K73oE3ApEiE2MCHbzL
TUtk8Fb4zTkIqJwVmfhd2umsycK+LpZEIi3OfTx0uHJUj29p/4ecMmbK7VEE/NmL
F1rHmT4uL7xyLBiho4Ls+XUvUeFXnFRoLCxq2Od2wehAyU4goieOx2DDti8t+Mwv
3qr4UU70wOEI3qX608I7XryKkR9xe3hfeiM0TVaZ9if2cmXpW4MfQ1mjM1eWUxHx
C+/kkRdaaFZOx5Qu/BFzB1Yh4aXu4O24ltK989x7l1zxIm67pQ+iVsZf0jbIWfTM
U5DX5iRSjB79YOLC4jZPtCtE2LqXCctUpn9PKsVy83LFmPdPf+12QP4Jn+baCb9v
QG9HZgiplpOAl19MfC8w5SYU72GIkMiNJFJ3IJZsyGz3svUy8G1gCXUU7SwLEkrO
Bf7NcMujoKTsIly2WsoFmu8k5KaHxXpym0XZ+I5K8L/yDdwuH4Q5P6obCuox/sum
Oo6L9CI03C6LX9TPTqchwSfJSIt/5lHjIRvC65jOLX+PNzgMX0PRtMkwo3frr5tg
AlewkFNpO57f/cSJio0yOR33TMbXZ1ADz4El8d+yD727OaQg3TtrUDADuHAep/0m
ry7zBT/mPBuOHNZVAGy1XMkaST7HqZZR3p7BhqoO64MJb+G7Kr4Vw1VLy5LWWmRE
O2o+vX2Z/LSpHa7De+Gxe5FkYL9KL+NEzMmlgVrNNX/mOMAxAkL/Uuu3O2FPRE3u
fz7+q37VNEn/vog6DHDpmLNJhFvfJSVUDPHFZhwmye1a6whpAJvrFyd5HAA8/KW9
wOx4XFbUJpDgQqbI+mwMDKwFU/jmWmZPjT8rrCw0R7DpYRTZDM3aC6UyZn0XqMyU
Y7P7qt9Icq90iYJYgOHdBB6odaP/BsgsNOFmqn3n1Fw0ATpAElcBdKy0MJ0XjlhH
HjbvJmRd9bdrAtY+ubt2uyncG5KtnmWNwrn7F6w/NCMKxMP9Mu/8otRg0M8XtURc
VjS14un6MUPgJFBRmquF56/zeukVHOZyU64Y35b0l7sdvQb41xRp+3BzAbn/E+tn
4GEmxAovGfrprEUkzE8wmVeRayCW7NB9eF8Dqafuq7HkA9faVR5OErSjDRb7QX+j
g7LP1HAGZ23j4halwhPh+0rHwUAFtb/e1LRRNlqMpzg0U+5CCpLj1Q1cgrqa5QKT
CWqx1CkuqrgmKIMjhbIV5qtId2A7FuLb3yxbjOISntKITVRSlDE0sbLCinrWXNDM
O14ZUQqrhEsFGPMKwXaPePfZtZyvlQZaBxkdxjIK1uHfHub2YCJMAdUJnRRscQo5
`protect END_PROTECTED
