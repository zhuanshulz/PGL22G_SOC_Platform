`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zHK57HvE2VRBW1ynlL0KtJZ9R8ZMxTZSudGsRXswZ/NYN+kHBu283S0h0qaccaZO
85JHqx5y8TXxGHY2JF6Uvs2tgFg6UdJhIemxBbcE4fJwerkw4yse+9NijfrQuexz
1QUyHn0qOTan4yY+qvjv+2C+bnU74Sijpzc2Y4o//2JWO+QP2V8H75L2EWDTJc4t
xYh5H2rqb93Ifr16LcyNhgkG0B40tW7i94h2rCypor34osPaY65QBB7AuMo4fipN
2p874Y/JCFsJFJo1r4PSDOgjlfDLmfzMj9qHnohBLvArAUtdSJx8YOw6XRWIqkZQ
uoRF1Ue46p8EIDz918Uqid/LgydhI9nw+CJcJzZE1y0xgXk4t91lP+RVhlA/th+h
/Rde9UjWOZpqh3JFnhf85pk8E/Yob5yCYfC5osPa02nTP+bAVjoYd0IfY7c0y8a6
FeWGxHUbZilRQV8tDxE/vk8dxtDhw/EMUEKH35ootuxNOYK8WchCWe3x0jo61dk5
VZd0wcdliaPHb8iXvri1XCkE3ceqF/U+mQEAf/0SoXFuaL+K/6u1AJ1Ahu0MNsmJ
YSE7oIdRg9fEPz2awiZVKQ484/cBIA9ron8GpFg+6rmSO0F2jROfKGOT/PP74gWf
AOgX7h5m/j3b6PO6Tp06GDOlGxJkmVatFwOQnCoE6hgjpmqfYe1yEzwpeTwpgJV/
lGPN3IRZAzkhyLFjokFBpecd+SdJXfto0EqhR8kgh3t77EazYSez+KeEWkffDA/t
83P5AqXwH7LH8ycshpc8e1QB8TU17s1yYeYofqJ4WAKdKepKARcHhJ0Pt7Jc48kl
RDp4z4e8mSTbNjFhBqF8dhdkkBVWRcLW1InQhKAIgwHp7TxltOjqHG+jNXgOhyRe
/1Cloi5dLizLfm6KcEgBqInYfxbw6QvTNOKf3he8znO4r3lqXiQhdxFC/78OSjaf
xKp8dhiU83z9kGTYiXTRFsNKXow7xquKk5bUFeYOImVWt8+p9D0roZw5+jIVW6KX
+fDw2Pg3+jOeyobGFYx0dRWRl6iI0FQmFBfBBlwsKQXDnUHqk2jW8GR7qIpbB+Rh
mXr/4Aclq170S5F4QJHOzH2xs34HDitObcEiwdrWI/3Yx4ank/Hk01Id0Q2Sjbdq
S+A8kbeJm+Z8YCPZbcSZi3ofcBrLcCbxGu+R40lLoP4YTn9eU9rIhAGd5vRSQ3c3
MKEj6wA+ByjI112eTAMzy5B0myH9/Gt6OK/+WeNZHDwRm9JbZu1DQvi6Ve873hyW
+3RMLzZifo/vEEyUZwPuMSTU1PXi9MuYp3WOcWYbDJSDQAdwjdjoWwFOSwwzvUtA
CmwBVPIg3mU4a4lhmAVuEF9XQBSJdgxCMxQwVaPG+jT9RVwc4nuS63evcZagP/Ta
v+9TnuOwXDIOv5HA/3OtQk+gZO2IQsamvQDK/5yMdNtqUO1jmDrpbMVWi+a2gu7g
xzf7siXq8hTtYMA5Bzjk+RyBf/qRDJdvGdA/IMq/kiC+VBUn2L5mRfdiKKYkV6z2
DJuUulNhP3lHoMt/DHaYgyILwm4XdnYQ5XpSaHVljwO5hOc5FFadaguRZg3wu1FK
ADCkwgwseABvoP7u9w08wXrHCkUSZH73WWj1VTNY4Gs=
`protect END_PROTECTED
