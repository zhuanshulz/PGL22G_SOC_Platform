`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xXfImEIse1oNnEb5KR1swF8D67qUq+dWZrvlw3AfcHyAuCm5jJY2/gyJBTtSjXOA
MkutYslmXR8HNhA1MS+r5XEzmTx5GgPdTHqfsK4FRSVt0iGvb60UHvTTaAtt4wec
FJHJ66PsGSRAOqZSHnY5tnBBaDqehWuSlNsoOo33zNfTsUN7a1cWpHB8iYFaV5vI
J5ebbiuHFWuTwPDl+56RROXQipl48SkQgqkGT2Z0hyKhAIqB5WVlhX9jFBgF2TQg
aLtXZb/j5RTXLKRHYufF38/bMpajlxsraqldlF9t6yVcLhoQWh4jnuCweU1ngsmI
+shSI0+xRlob9O2oShC1WPQvwDJdv0BObaXABxQivq7mFz4wv24FmTd49AfNC//0
lyCEJbuZg/IHyMM+Uh2JMe/q/3jWapm0e1knP+LawoRGTQFPXforFoo2IwHp1dl4
tSgy5MSmzoRBK2Ho7d53LJ6ytOoVEzvbU5aC4uothjA32QShPQ7E8Kq7FUlThdfX
BbtoAw4T10JyMpedVs3KTZIKxU2CbhVsQ5COXbLbO3SNnpFIhM4xHrz5UaAtb6Ti
ArdpuU6CRvRZvI/g5uos+pDWr358G3P3nO+L3UsOOk+nZoMB7Z3XsjaNem0Tt8bS
0Db3Jb2jm8BSHLTj5TxNV+fSa+J78aQMUlmwEICZufJe+zi8DMSLho3orQalF1kl
9q6UPWbhyox7oWWvx8IPMQi9PgYVRZlnz7E8ZosRvB4nqOgX/VtSbtY3xf7Qe/xL
+zEI8z7S+On0oCg6YN3FuunabkpXCE8SA7Y0VvJIcSrJ9GEDJpl53W5bBzkUZ3QL
SSMpkdIlR5gShPtkC8EwSyIJH9pOgOwq+to3WNoc6cbMEI9MPQRKyozfsqb6qF9C
dZU1M8eeWKWtmUopBK78dkvYnSczzN7WXVCyn4iTM4rZHNNbjOm0n6nya2rKdG1Z
6eRc/0ZtOP1v9k+hk388/2ExZByKTQPD1l6gMO1RAG1HHfFWalSl+buhbKCreMMY
pdEd/FF4P94rAQlsPorywwwzP3g9sA7+Iblkz50+Cdb8kWqajTi/EEAIozI1aB7C
0N+odjr1LPti46ILrLmb2Ghbn8DRZWrlisLnycyqp/OjBh5Afl3qLYshBm+oHoFh
13qh4Nk4hi8e/HQMxaXAOx5Ibk/sRLCZdgToVB4sS3Wg8Sx73W0pqMx/+8Z6adpK
irP56B8m0g+0Ts1xAkU07hm7i50iTGHlmYiW2qZO6tMjYdyOLHxqovGliHZXsVRp
wC6tjjjQnj/xybX+3T1DLuGaNsWlPxSjnLGzOOVpohEWW8BNIpwZv2Ye8bKfVH3c
fyLVT5H0/kNkRvEo6t1i8DJzeY9Y3acS54CGNUkM/dxkfLCDGjj0ICAIkoIEg1GP
BftbtZgpyR/lLcLdlMt8XPVIond03ODzjAkLamtyrQdLOcikG+IPC2K8V6tMeHox
qMd70pA/RmmQvLkEzbvTdnZxian27tCS5mGs4j0lbmq9BxdNEa1FSjdlWn6IJd1A
DacRVe1sT6Yp+OJWU/vKEvOrU0/IZymhRictbS/TqjUQV/PCayoO9zE4WUDdDkU1
IxBykkXnEnh3urLuRWgZigfE2QQxQkr/len8rCqMSCvUlNnrQbwOoc1cLC895d9h
F1QXKgPJai4KKyfn3EPG6klXO8mcX9chJtm9FxB6qLRKhBnzsJ4qMma14+0D85n9
lPugvNaXaVV/ePvx5hamlZE2tE39YNXz0FLZZ1vyn9PjsVKsYpTTVx7uUhiR6rK1
fpbTnoFjq58nAjsPvO8oEOVvLcTVI+Ao945nasgRYTxTSa9bSH2nshGeFNyFS2Tg
9Bvp0Pn17o8tPXcG3KRSF6PRsjTx4ku97lgNJM4hL+IAMewx/a18c6VNxCrrxqca
e5iXOzLvFk9BPYcknTyMrq7VDKGXhDQZQjzniCshymX5kd/vorGyT+U54y/KMV13
PcWB5C9KZTQTPwkjOQVnOBbm1DUbdqv7mWrEXB3pLPNf7D/495VEG371C6jhFpmq
KSrPhp+UPnKd0ORMhiTzAo8RNAGm2lBbdxjLmJYNeKd8lD3eq84Mn3/wkj9xL1A6
XVcFQwTWbCnmeiNZtW5YQ3KJI2BzZrHZ0StwrVpNHnXJeZuMBm4DgI8htDAHiUFs
7h7iyPiOPKhkndKbVYGeLYQyIE3DR+c1G6HF9KePN74Kr906pavx34bzJ5S8GLA+
wAyAGIaFwtfEF+sWxQbJUhdRtR98WjDh/UCWvrksrPMuWHgtMs/UlR76KnEr1gCN
YgPdzQ6mUMYKT80Wr/ktl6L9n6cqkId9XgVrNhlmspM2Y7QlYL56eZHlaD7uC8km
8hD4yhcdEwfgerxERffWFWiEBezQwBaAWODNlZZHocJUOZtJ9Z9Mo++h75VfHuDu
OOxALvSJkMPIqsSxNt827KYpjndatSWg0o0gzKAZKAv0GEDi1JVJS8rQnGDqWWgK
q5OusxnWani5d0kn9uaIx/zbT6+nQxCLSiwIszH10F82vqj2LJZXSCEVVzP9s7kd
ij2PP9cv1XWvZkb0012zJOeh12bW8grzUAkwtNm/BWgOPA60SWkoeW17IUvKHiz0
zketvM7t2Y8ozrE2fPw5neuMet7JGd2si5QkY2xnIomp1LmvbxXlqBzDMWdTAYrY
fPlCCL0+BxUzIB+zPG1LIgfr8UV/7GzuvDLemK2UMOVvNP5K6TOsX+LBFvLpIgPI
bDKWxXBpbQlWSeYnRvjcCJzabkHFjJF7FadQXsG++IuOnoYrCAc1k1SfZGaL2l7O
AfNknCWCD8HmwdlAhS9RGumvDi7XA/iaIGv+Oqg2KmLNeL24bKd5ysJeA9F/7Xj+
rDo2rvM+aW3kkjNDfnewyyuaQrKyI0pJ/tGVJIE606giIy0cPIpp66fk/jTMHdfu
3vdBsaaM8hNfrLye6NKXQc0UHO59JDDKsCJ+CDaqZAJvhziI9C9/gSuF+TInAwMS
9TzqvOtQauO1tvhC0oXA4uciq2xpTb7vUDDWAFwOMetxXysP8Q3v5kHF1Sd7JK5h
h6KyDEHJy4e6fQSQXv0koEgEm/29KPFhe9YrTx0t+qdLHCQD1jGr09bI1pubwdlR
pVbgchy5NE/JU9bTw9+vMIe0UEjhe404/oQeJv5vU5BTxgsUuQKVTadzavxkWkcW
gfAC0eZma2vbHzzAIbxC0jGUICp9u8DTLd80cXZf/etfs5x+TnkRXIMUVT8DXpM7
6GV6+cnfU2CZ7LqHB4cnKQ8altjXz//9Q8BlLvkPpzpnOuG6RuHiLkuW8FloLghW
kXwZwD23VMDF4IBcz+OQyNt/bo/fW/amp5VW/+LCRM1JdQGCMZNbFy9+WXizMpCa
t8WsJma7JUk3TSz9wX7iUNgx8mtIdSWsz274n+6hqgqDtiZPUg9qAgHaMpXrqhr4
bBCU1L67kgl2efnWrSN8Gt6ka1WMv6kFIaYKh0V5shSFbjVZY72kJkRsNaq6fLn1
J9BgrnrkHDnGYicWPb+6YcmUwo3yRx+p9Z8M+eRTsBz6imuLX9bOgx+Nk/seRadq
Q4AVSp6CFe6l7PeAIlw+AB1PizfhLUowWBfeILngGQEcN6EEs/G/RmwEnuXM1if1
p/xjh5XiqN+pzO4Y/rpZOZzxrmJn83cjDoIBuoH2+bEhSJ1r/EYBH9S1FB2alsZF
ppZeK8goKtVJJ5KcTg7UTFD+MaEZ+SqfGVu1HuNL69YJV2ZmaEQ9EhwtpqraHteM
6pjEhAe5Np/f4wKKhcKC+sGCWKJtrXobKPXbss6d9kZJBxcRveaAq1bu2KEDQAJL
oHohX3GffGeeyqo+V/f8Ii0mc4NXRtGf0HA2PFPOHwHlyko7J+ljHSMpeRNpymXg
xTDvHA6J+ZyljE4/+oE5VNKd3f+rmhy4TgApw4Q+aBiI8iKKmdOCY9/BgqWtu1N3
bY5B6T6hEqMHll7llDnN4Ox5+GvgQhpYB/ymJVnJSttW8KBEzQh6OvCndgCxnh2i
6xnyjFojW8LW8af4Kwn5Ll4YcPF/m4oxtO0KTfwMIPfIKlzKka6Gy/Yx5SHVa46g
PduGukPskfHjTYhPyOUkTldY86q3jN5BrZ2ul3v5YFlllfLELy/X+918nFX9QR4W
f0xYJJzuuXijFURI41GGiMxsw7R0daGMtq70azKPYue5gssUaNM5bQky2Pggeuy2
eRMY2CjAca2phodV26IrSlx8J/ED7TDVdSL7Y4BWDQ1kAgZMsbrxjzSJV8XvyhuH
ZuyB3TaDHdyHNDtpsk+ZDq1LyKABSzTYTB2tzwX5MUyXKxKkdn7gChALrLaVUnGn
2O3FqAHYiqEQUgnGAuKAVmw5iSugAU2CiAooxxzT9v4QzXxcWTQfmdgKnkx4L+0b
M6tg8gXRVK0ZXCWNXXdycBZVkoJvllQeTB7lq760gFO44LNOPkgRxJX5gxKibQCn
KmaoV6YPbBK5iwxxAIMipms1cJ5zfLnqzGXZ7iycLafk16b2Xut7k9s9nQD/dbli
PCHY8+cDAThPHbBY8JltQ1H3T3EnKncC6CJ0MAsnYuTrlMYdkFWKOMl6QojFl6H7
hH1xr27PDF2zaaK3dF2/Jybq/6RYITDOzAv2HijoP/hjOXBIhPSekt02HPBailWT
+SAzVJSikznqIAuKFIu++wubL9q54UQBKwMaDO8a7e1h+4ziFBOCcw0pu8HkCe38
4sICoMxmBer3OYM6wH/NyePXUzoXF0R4StsjBzJZM/5WvBdS0LoZVW42tj494SHW
CqkHse5c3ECRJxVdeXsRwnhETfczDyx7eTwZZhwleY6tIDYnOdy0U3q3zfkBs6qm
NKWYTth1LLxb2B+71JWxXZwdWgZnuwkWLZdqOExKIchaEc5DOzwfp/klHjdmwt7u
Cy2olzdJpnzQ/Mm90YN9BQImfLmxgDA+8zpumaEi4DrJ1yw3uw71vBolT6RfUirg
`protect END_PROTECTED
