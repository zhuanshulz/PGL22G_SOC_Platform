`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aRgb1RsfPCzVbf4kteNjuWc+AaysCrlNQfQaPoXUKwjopGcy4M8rUHtvxyaa/npH
f9EkGKhDC1F8lhWW0EMBbq7VoX+m1aCz5p8j5mzVyKZmZtzr5QoeaCEGMUoZSVKo
YToYTAZh0z0b+SFcgT08Ndf2iDISGnx6wXFswt5sBKyridi4xzqd9yGe+68LeRzm
XrTZ74xglRj/MLxO/1G2Haw9Oz+EXyrt8MGIAYGJhxVQacNl+0sr8nZlb+Fd2n+2
i+iRPrKpdHqkHyjjI8yiE0Ik6dVNkjBd1j6ACIzQoKo6IX5A73HUwDXJCuO6U68r
d3VDiOijNWMTRD9fe9Yp//v2ZRloIuXAGuokqYfE758VlG8WRdbrAzl9D5IUaFfJ
ObsDW0uF9bxwUdtLNWdUWhVudqvs5eBDCwSbSH7ujYQR6gRDvtvPh2qzcrejIFar
MqcQX24Te1vEy9SB6ifVE/b2b3UyfhcyMs3/74Mn82QIZk+40XgASDMLeXZkUwvK
0xQHdDTriPP2kknzIIcA3HZTnN3LAW2E+yp+Q+Dvnn+rasUhBZaTOttnV4v1c4Uw
5GDitPY8qfQddDDrM6FBmGpRrKzYitPKGcplE75oEbX2AJMQqEwFqRR0TVp+4kgZ
UMZo5uPCrlSQ/GHoi5Q+ByXJURmxJptBgQDzndeHaeseqiqKypkXdmHAo11GDfqo
QeOtgKjqRpXBEMSTiTOQz6NaH4Olvy1pBmjCaJ16EdiCT84wWArN00LMzztW8BfW
jEyncMKLzsz6suiiqZK1ZrrshIU8ZG2HRwkbroV0nw9fOTJnvDLOrle3uqGQE8Qy
zf/u45U641sLRXE/N4vjSOh0Tu8seFzhWfZm3VarZM/rPEfDl/2jjDhS2qICEeD9
VWOy4gamnx22g8z4gr1QNJymsf3C36cuEmcZ7wgqC11JETYsjH74U5/ryYEI7RcP
qqhy9wgHxKFZV9MzJDP5mof+V74I38rzWM0bDi/669baRFkZ5+XBZb5MrRb88CDN
jEVcMs9V9FiYaIVhLezPy4Ukxna2fyQCv1IIb0kfhG7ru7/N/BQh3bVEKZ2K16nj
4sKDXkzi0uAiwOWw0ftR7zHswmgb1KYWSmDJ6u0NJ8AyYvcN+QTRv5N48Dessmre
jpxJJdZfefazlpH13AmaJSIfMpi1yKZLYsox+XzHPPHug7c8ZFNzj/oCeH3CsvzV
pKMTdN8X1dup07yeNaZ2ErR01/DvdWRiw0Etce1UUnTtc1j0Jm/0vSWOSv5GCrBj
eAAv06jXZ0mNG+/rWOs2jROkcX3/+wZZGF1wuTL7MC4YOFC/0ZgLntNkPNyo3vTD
IDp9Nc7z1VGAx8GxsUHWzxmz+YnPtlKACHCmZEEPdsPT02x4e7sfn5iu+hzwoSf7
SazSIUOrCePG2na6Y6HBu05TDdX5FwGPhVgP8ZUTKF1VeCoDBJF4rSdt16tYwtwj
j14Kw5RXmUfNGtxDyQQDbABnrDBlJw0G/9Nf8YOpGsPwQlttG3N5HOCTkj++ORkm
U4fcFM8jA8evLZl/PzQxl2WBNI5Iekf1xixhSRu95liAbgmIpjgf/GMtmfeDF9xL
m4SYPFIAqeSH/KzOtfwkQC3gi4qQFMGEeBGHFyhsQrBqSO08v843rDOPnENYwNv1
iSbZWrpsxS812pFme1Is0HuPnmcJ310lp85NVI+TRR2hWlbaVRy52VRRhmAiHpGB
vFvzUp5cQ/piwVg2qg6Q87b4a3dDig+In6nBCW2a+TS6GqEADk/BrgcES7MNrEbT
O5o+9B5vNN5wvibimPsDaU7AFD2lHcQEp2zudoiPWUzIJ4o5QJQTf7iDT73YtLJN
VCvm33ULhllkQs1xQADyJbNjA/HrfokoUQ6Lvv4kaLMVMBkp2+pD3XOORDe5YH+B
uWoMolYXuc30vVDRt8Cz1K6j9WRLbshB2bqOd9ibJtyEX0aNqNw3XWi2Iyv9Krlk
ysBlMHFFNKTxGnydwk/QWJ2qQsCy67TZIPKb4JdDbKjOC7lnTBk6bACYD253Kh53
Qk1C/yMV7aSxfPSjVjmASLQROtwRN7+L/ri/fgl9QAZPPMlIlCLCXqjyhvoeQMwS
+cbEZeN783fhk8l9dcXI6d37bMOYmYO2SKFflCXIHtTJgw6GYRmjwCGmasUS8d1T
94nXpGYC67D1PpoxfT2MwXaNNeGnvAtF7xth1bChr4wPnDvPivTVwtp5VRzINCeH
dIvDTmaiz47FjQTIXin1ZhkkmWyzhMtocdQ6KXM3ZiS1DLbuYF961Z3IqTEXLM0g
RQ06aHUHMpm8kNU/L8VYm45ZRLA4qdCfL97Hj6I6h8uBGIx5NARvCMUHTXGJ2pxX
D/dCFcDobeHsR57d0I7rOjnfCONZ9p2Odsc/FKr4fQkmjcIhaQwyNc5Rpqb8QJgc
oWdW9SVIBH1diV0xALFh8VlYykH5MybsmCGr++Wxeswz1BdPV752wb671HjzlaKa
DXxs6WIUVHS3YtA+8Sc3Q/3hxL+zmts0QumYEdUes2YYFgGygATvr00I6xEXngsN
PzcgoMerKgEhDj6ab5ozD1mt50cmqYZqJzigReeINrNjKI8vmVJ4ZIdUPqLYKq8U
qrGMw3iiXQF2VGHhhAE+1QiaC/wZRLSL+zA6KE0kQDcpS4BlF5Eo1+7MQCEMFoti
gGbp0J6XHvsBI3WItd4aCDPjUwyi0sMwr3SrkRaEFLXUgKvCnzoaUpOGbKENiXQt
eIti2iE08vc00E3lOw4gtUtH5wc0OJZvsMHBRBJm427i/HgJGX2mznAH0ZK/Mc94
9eRLE//I9FHOTxdI/PXlPsLhPQifKevm1C7hIFpD85SrmQVDM3eNUDVrQiMDOFG0
y22rQ6yoM8Y+NMwU5qm2HjcjrL34hdNhA6PR9zNF47pSDlR4pET65CcCaEJVAFy1
/EHhG+11iq8gadTGCaVws93BdHbPDBFfF8n5n0HxpNDzNd4P4+iMbPr+2DXgXBa3
PcBaoIXJM6xa1V2Pid3gl6ulcZ4+4z8lG2yfgVubSMau8+W7dNfHfbL3lEwR0ryR
uEHI7PtR7X8oZH7Cs0V55OL2lrhm8zAUtwST6YALJOkRzesGb/f063DqjyFxbZlx
M+EcrGtpw9JzmPVf7u3ykXEjm50u6vBMzBsiNhnQzPE157Z7EDkodzN/FZcv/k5G
tKkfy60s7CVmtFdxA8J1cpzTrLnyDOFi/Z+juiNMzNeGnW+G25l07fGJ+6l6K0u9
83LuDGQtqspY/UfHWc8IntN70t3DeONH6mzuml7zF2605gqh0ErHzhi6vNaS80I/
mCUKgW53skMNEkNvWOlNniTYC3gZpGKm/YtED0grfOefvsQYcd4Z12f/eMVkJpWx
HrozExKWaRkKmdnXRbv+eTbybXN93xLXIbStCqiTBeQ3od6zW2YeksTAClYixyY1
OkC+hfaQB4m1e0oKwYwx7Le1KNMBZGe9ot/EwV2q4HpnmrWLwbIyBAkzP8W208z4
pyP9ylEBqktC+RABaBruTIgrso/hVRAl5UB64Yj1WfZp8gRrCMrij/yCINETyl0N
5l/Is5+gaYPEMk1IOpbJtu2KijvdQHSq4KV1NJL+pZ5YUYefednvglMLC0kbwlfk
CNretjkCuD9mEn0e6J9SP35ptgsBt2wmT9vA65MLpJBHujDqQvZ0e+W3UxT0EboM
EteqltAwGVl6fSTdt3HCM6yt+0gpv90kjc/RlK0rGs5f6zPlPkw6s6zS8K9Jjb7e
3lOaFbHPRy82M//TAMK7rUdE7PNPXcOc13lCbJU+kbhPDhEsE+2aa1sEH/xtyiFm
KHUUSvWPCBggtKqAZN7RZKBULSeA92QX0ck7w7BhTRZF2GVTMvkiQoKhdPmi7P+m
1OmBD6NrgcvcccVsohc8NYXKZElDNQFo1pj7xu1Ziglogzqw4KzZRHQ+kjog67a0
Q5DnE/9QVtGZnV2LmZw12I5mgVCUkaEzqi3FOCF64o10Cx6SOwx2P6jbD2KtXiXz
1igEXrzQ+qAEZCAQ5tG0zwZleD0E31CYCbTLxbTFWov55ptMXJBP++LIuPxyh+Yj
Sp0YsIWRhO3DeveBYrMos7ZGHouVDgLNlAIGSaUxb/C/KS/v9l++0/PE7meZJSpV
dyEBnxsoSFf+VgN3KGPxAFe/Ton2jHNQJZURg9Z6ZSdp0FjqUmGZ53udDP8f20YK
rl4N/g9YVG9YAN7gAZOsCddOC8ArPe5ZZ/ESnv2W2RPQtQ+8g8Y0bXvB8PHMaSTS
WOPceDk0wy2VsKO0YZImVy3D1zhuKuYBaA0epq9R4akEUCHE6edYoVK2RqFaEEj9
dzuHt2tnCsgePb6QIRQnOdcDE6L3pNrt4DiVYMW2toHMhWXNzRkgXwkZ5ILneOFA
p0jxBz0pWBRZiuW/C7ajKjwkBvQ5hszakxBdv4FRQGra8bOaUnUNq8FlPtYiNEDm
2ikDY2TE8gPNT0NOxCIFbmRRiu6lOaALHifCT6J5h65LJMkGV4m4fc1jL2AlUhMk
YHLE6o48MP2N1+kYttUmgWAZlgCn6UfMd2Cuf2JdF+fXp9FapGznYlf+80ADrUdj
O0QYqqfwrjxwpZbrxnMNfXRruQDiRASYEB1J1epkIk+/g03TLpTYtFDIs6Z1uA6q
FYGcPuiiOxEya2H/j4g6h7YGyL5YSCZCobFjHBdETf2Rnv00/qUqcYtkUsjc6uXg
Illy78bIOG2EBWUBg2ovlTm/bbhzMO64rf6iAB2ynC+atXfQDTya0Zh43M0t6okn
7vQnriIEVfe1wwjtrzp2zsfs+EJPuc5jFd3o6iBoFId8BEq7j1OsAtvPvZeMWSIC
RO4dF0B0LHS7wE3JcX/3uqaxrcl9zLgD3iiVfia7SKY1OKKQ1ENZboHI//InHVS6
Xe+hgau+ZDDnI+G2AHKMNPRd2r1XHDHtAHNH6ns6zV1tITFp0dWA/JZYV/ZtKnG5
Jo2rfh5p1tkNIgbvXByUdiN7g9dg+1Mz8wdunWewjOhnJ9kSTmMqD3K3AfG+rm9m
LYPHXGI6oNXoAjG0NyEGJNes17C4uhKCaHu8LNixIb4jTSmznLhokVLo6LntaaAH
Aw3cK/iyUPU9fBARtVS0U9Vy+D1o+p/86gzpmwajchY+HXvT1whqcY2R8rETTKOn
X2+K75jRK9R52mgAPLFWZrw6eST6rd84R2c9vussKX0XfQkt9JTJT2Q8IwdNfPjp
ojhmVF38gTw2FuQy1fK1yN+W/Bc3EikIZlDRoYYcXqMvaEEk9JEpCHrTe38x/dCB
nZwNIkC+Mweqh+gitEUYFfvdbftqjsWgwJan3rYS9RjaXn1NzOy04XZNEjHAGAeT
5kamTaK+O0EQaa78WQ/eJLM9+kzhxIbeU9TjBYxpO0EwaE++PL+cqySf0kO4n7zq
ttG2ogA/KJQgk1Am1tYxuU4GbHL75SNGxyZPPLaQB+Js6Rjq5Iq0s/gdsDofHdLw
wa5BuVp7iuZ7pTn1Tp+TJa2F+8h6eiujqlso2+zGcwokvwcuNZSDxq/PIhmMJ5La
bNMXQp7c1ed3kgvxNAW0j9qyHa1i/7v42ZPifEnx+VJrDgbEI6xrcw2GImqYmgVK
Zx/NDu5agT4fLLdetB8V7zwJywN6y2LSqRW81iXAlo0NiMuffU766NfraTbOhZVl
N7AW0jzCnUlJRCaZoX/EsgBuMf+Sm82Xnka2XIexQ5HyVFkY9Mcg9/IsK+KMtoV3
D9QB4D5Ao/EZJVmQEWdFQ0/KaUpAwPo3plqTrTRohh7V3Eh+hNdebqwnxk4RVaym
XRcF910C+lhOfZ7X9DonX83FXaUW1C/WU6fMI7pBh0uE6aF4JDVtaCUsnWQS9hsA
4tRkCxoen4b7UbNLBp8XqttUnOcKYisub9WyRZS8uN8IWseFTA0wMAx98IClSnsU
OtcBneIK+EYkkqx3hBXDnCd7/32JaWXo5l8LsXwfMjuWFDW/5aCJ4DX8MFdP+6zF
wDkbrPGmXu6Iv85K5BasBkOjVOr7zVJLOVYwsuRhtt8gsdhi2dUtTL7aLgI7ZdwS
GMCVIXI8lVO5yc9w0v43LcrjQjdxKpMz8/bmEEFyxofRPkiJ6Bz5oPqXgMt3DOJA
QYAAezsxPVzfcO3oVzm+6fu0SWA/lucjF/jw3OOHxLfV2qXh2QCmMoAKaFpxo1fd
Qujc+HGNFg/DNdXNBZvvykIIdlHU2Aslcp/6lkXNeObzxHAB0ECB94Wj4TUi8MGr
+Sgt+vTgfN2BSHPa3PBkKnLW2DA4u5Dp96OZSA7ghCGjw/FWJLACX+zA6j02wrb1
EvH2KPK+dg9dSEg0sZXiSIUZN0kGXnMfot9bR/7mKzvfP4+Gvg0FwgelFlCsv1hY
8IKMAidHIDXtky4pFYLnv9p0SV1eVvopHED0qQKZi5PubcMlv6c6oV/o5XKCOu2v
wqivG45pkhr3olhM+gH1HjHkrhEwVEZNhAbtjec1urDyP0xuuJDA2Hnv91MxCDgq
FDaGSYWFh4j+tof5E/TBc7mQJtMbLIi8M/JceZ2FjeyfBcyJXzy/cPniA7A/DSbh
QvMqcQMO7pGDrIZK9DW6ke0NGY15EyyaUzKILozhkZnYjEHfcUulq6buyaT4t751
j3ctrVXToRpxnJ8G5XhEBXJQgsO/y05gmduBFj2TapRyr8dj0lya28zTSacW/Mis
EUdUKTd0BEYTyWXCcPOE1FSzgISLnnwx/DzSV6eu4htVSn5icmvdFEedpgR6ncaR
tSp6ClXXtGchuwyPfeuwO98B3OG1/OYpkeGIKmkL3AaSgY2VBfjTV22ZSTLArq7c
mOBWJWs85g5qHIKqzLHB5pT0yfh/CAhIFzIbMOyFpS1mUncN7T01ByXgoQc4a2qT
Y3MAH3hkxnilKBFgyRHZzKtPEYH8K5LlhoZmHx1NKM1BzqYKne9KUnpdAPWPMAvK
TCj+cayRRukz7F0ujdYY7ILqp+fVqDcwo7f8742hDHGqwnNOrqa7VKVYFqXWzqCa
jHD4jq0E9blOjcoTWbaC/3mHhEikSATqmZvJblSfXoBmre1GKdPu4pQOV3zvM6/G
Gvdu0VgWM3ZfgBetgFNmB0CqIYN/nopvXUtuTSF9B1mrePA6BEP4UABQ0wYJEVkV
doha7unYq18fVImcuhfoV1EvX5nrfVUTXfPsbuXp3v2x49KBUV8luruujEHRJ5ue
R+1McnqLqeuCq8mVvAmLaNm+WohATmk/VqEYj5p2IY13X0fO9+qBJox0zw5I7qMz
mK9GUNZ1SbvrPCjwy22ecF3xPuGMxvHHhbloIE/kTMbJPInvQhaZERK/AvqOGZEj
duQawerV90y4yt4vyXtZvUL++/QarHqiuPjz3qpuaOXNl74i+bvskh2p4xXRRo/Q
6vvSxZw8kOa4hPP3pIe5qaCYgr7mKM+t7yhSMuUxymQuOK5dt50fArGUu00zxaLZ
/cbiGXpcs4vsLQ54qBhAPBT+wBiNCpJQfCVDntzHaGWpJF4SWXyq8a+2HgP/jbvi
UsCS1O4esbvNjUbOQ1NiT7nqJbnnM1qbsTzZl4WhZYU0w3i03UZD9t7kYU4/qe/Z
EmX4G51fL4J40D7njAwumIfgYsSARsDX8nv+erlifJ6ehjfQqhMYXYLp9thgZJ/d
vamvh6eaiBp62TBWv0v1G/aML0KFLVX2OQ9L0GWhDrBfZjnS+X6jOxDWLFNo6Cg6
oRKJnf7GtCM0CZ9e1leXO4dkx/f0u7r2VAzsft9SlVRNXvbBHN38uIEizPhOjfHM
0nqjvesGS+LMFtwGTK4yrtspM4/Sj5y4Lnp98uv7AzoMkeiQfwOoufAZ6AgBX0OA
aVY3+HWKQHbSK1LBxSBzci4p97fOY5e+LWTgonrfIzKsMY/EC/UXYFnYqBX7RWY/
tjDRgOD/eCVR6msQ7ZQNwwaR/vkQnyGKq5FBpTZ+ObGhqwa7HAiqyNrtOpQw3mSF
M0n29xoRfKlSlVS3FENLXyamI44574KNwMx0ToMkTujor8rq/xNBTO7CxD2UKzt7
YTqsGffncnNBAVxMUAgkKYGD0fL+9QQJUvY9+S8hiybuwr0ywVeWUMGbG32SG7R+
LoP21ye80lZc+cEtaLbBjXcL7A/0lxBEXCJ9ACQNJCnn7Q/iVL6aODXNHwUdOSm2
FToxVOn1xe3hbKt6yWQfTtplEm9BSblikTfrLz1rDzwchuuUXMZdxeLoEabgXmcu
4yIbhnWXn/XB46qMmU+AhISUMa+g1UlnKzgZe+f5QdWqUZmOZhCWWuIRM6KLMskG
p3WvkkWt/2Vsc+1G4A2j01R662P1LP011SYK2B8lHpGsRnGtHIwsps/1ToSnP7wY
bX3cJd0VFvwTKtyy2u19oNY1RsFR6ngQittzw7OS8GqI7IBkEDsZhhslvQKdV7jV
OvldkPbRogOfM9kNA9+Hj5ymP7Q63eAz2IHX8dmmCB+Uq/IDz2kcdn0DQmscsfCU
0KvA8HZNg7MEAvOkNh4VIbz1PgE1DJnOC06LS5B/B6APfEjIljBr3jIFENEmpxEY
YuVmqwnmmq58io/3T5Gipt8xzaih3zhpuNlcvEkyaZ5xznsiiGd4I9IOkmdFwgxb
PcEun49sbw7ucRzBYLJBZp1U85Xt33XcB5RdQ3egMCiCGKUKljJ7MYfTWNEn5M4E
BLoQrfgDfYqxsE/MnmJj76Bxf2i00s62Q5cAPs7oSoQPt8oquSpifVF+lrdubQS6
DI/IsTDwZFYBbYijXmRANRSvo6q4KBX0iULdXMOsrQmQBmSmTT2dcAGJKoG6TQFS
52q7ShViMwNHN3Wwo0W+9pd6diPw1y1DSnzR8PyT6od99JmktBKkGAtdl3m+zeXq
RQVaVci6S+SHoFfRMBN8OItGnZ23UjWzDucdaMrQPM5yhSqrgq0tGq6NGHhSQi8B
inplFJfleyPJKkO/lLA6v/NbYUECBpyZwDq6fkvtIcw3U9TcKSAHxPVKB7S91jos
N1/5IeTh3eApz9mwuaAHI/HB+zcbbGyHwoC8bcSv3HR3Yd6mRv7dXxD0GfbQXIVw
mCJYh1nUgTgd4BDQqkwuJi52QUTj6FWwAogWrvjBybfbJdoe0ml+0HvPsTWkQgS2
MVO9rD32MObuEGZfamCjnC5+8fZR7LH6EXQrhoqVqs1RK2L4u1+xo4cgpXN1ITFG
s41i08Ubs0X951D6aLmIE5yNysZUq1zIba1zOQQAUFLpGyULlsAByqkUWZ6KqG4O
4Iqft8YJnnpQ5Tm5E4uy6w9qYrGCdiDMWi+QShe/E4TN3CQ0IQNPUtklGvEPUXa4
anSvlxksXpQRNRxc/zzuuWOUjL+Shx8W4cFof2Oow+a0cXpchwxEdm1gJULzIDr8
yCs6GugzgSVjJQZqmAfl5vvMQL//WQ7v2mSmiY4x4VW+v009Kl/mrHUBUoo1RYUh
+MMbewkNRg6vRd917ZHunOzYb9g/nGDSJGPTwOwRRV0FgCrfklpEKakP4FqaBbR4
K96GJ806do8ZVnuJ9RGTkLw1W2ZEWHMxd/t1Mrg1ryhbTYHTxUh4NK8tYs3EeTfn
B+3IP+FewkIdIJZG1rHDVPbHrsLjLoqN32Aq309oP43ye71rzgSBXjyynZE6tn8y
Lt/Hnd0WGA4zxTCOgiSQhdX8D3V1qTW40X1UfLy3Jdn++2h/xz5//0K+jFAhE1RI
ap390qCoOJlfp9J6Qu/A7g362j2VvG7cHO6HBHHuh6np/GRs3MLF9Q7RA2A5t/Op
63Gqq2itX3G14aZjGT/dU8uaY+KPjbiy2gcV7mw9EtjGbvb9gGjVUf+cH+O4vde7
AkzcAm0juBMHLFMqXmsSIta3Xa6hffZCKKezajX70A9z3SXtq7lpDLRGMZiztEIN
KA3dOWEzX1mq0+BGv+AafBfEx3/YkT23iGHRQj2LpUbfERH22kcOzVaiAmrWcmVz
aPTsgs6Mwx7eV8R4Yi5oSZfCogNf+MufdULsL6PEAmJzmGbGxK2jjeymskgHUXnV
NPoJ4tRMLkXV0jUvGAL0WWkBHDXkJoGkciDNfxAFKTatqLww7n5M7UtNZt647ZhR
Ks4I1N9N7/tcfz+ZWVpTQjL2pGOsNK5MI+zAi21Rfc/jifPE+qr7P87ZffStbspS
zeQboiIoBmE7WgYvkYWsLXf6PvYnAD2MC10ejeALSw7lY2KitegqDgqgmNMrnuEq
YXU1CUMpWs6j6XwsgOBRq9TnhZWqCW03GlDfvUBw3KXm7haecIBjclqNaT/ZLrWs
axbcOvWcIu5F5B0o/cQ2SDso9w7UizacGhm3xPuGl0SMDnJjf8Qpt821arpZCtzm
QTulF+KUb+Bx4cSY5YMRESdyPjgId/4yC0gp+FTUAngGhuGoY2OYb/grTHMkoegM
lvvjBJBbauG58/BlDL+F3WeRnNOIMTmktepe5vp5M3K9UuzwGy2ZmIuMuZNR1XtZ
tH+QaSI6CN8udowwFkk/Si1/lI7NgrbHE4cipKgIZADpZLQeGOAUeEDL/7WrCwEy
d3QCj0o+x/drnJJJl/sAmnisbmq2x9V5usBMwL+5XvqVieKf/pDztB+Q1snt4Rpu
eFUfaGtnLAsqhGaSSCxfzu29+ek/knr3vD141nXrUX2N9KtYHIu1JZFRev/q5/PN
evL4xY/zjn6HeL+TkFHjdMsf1uhM+eoxONJtMbXmbq9r/WFP6PbEyDMOoVOym808
s5ewcZ+puQdeRyXctX8dzlnNxsiRTvppljDRa8w1ldqZzDd0akOJNh57XfH+rct8
5G4mZ5gZOSATkBcw1mSH0J6IsJSzUpiNGW3niz+cXvqx4Y+tIRUHvhVW5+sQq5AR
l/QUNZV/mFE8AsHmNw3PV1qLNYSYGyiOdBj6brn0g0AUUELc6Dm4MzNGuakNiduU
Vg/gbtfWpZCuNpqO97BR8sXG/6Pd2OrIDx4l3+B1LvIqmWOQJWDu61Ep7viBdATR
9ptEnvYz+9rz7KNqOJ8GMu8C4R0v/QY+3OviPqD9VF0XWavqXFmqJOTTmfO8ptKx
wxKtOFuhJZo4Vz1J4MOdKKV84m94GJxcMeCE8m3LsY4eEG4oJ9soIRqYKLvtx5Bs
01MLNms9P/WbGy8fLgD92+/CXGkwdLbwB7LIPIY4oBT+AC1djDASFJ7AAyKPWVi7
KaUKBIlY7zXasgYIhnE0LgJpR62Jl6FfMX47obFqMcf9BsxTug9N6da9G9c48j35
FYvsjvg0Ih2/vkaw9FQwqy5mActzMUG4sQM7ZBgKFg2RNP6TpqSTBHB4oh+ZbhuX
CbagodGfynxUtALNXS67dDsuwZNYkyBb56RzvgTaPAHqD0Ln5KQCUg6bkO8A7SK9
Q3U4iOXBNVTSpiANZoFqq2HTddpxQr7hPBAFKR231iIMtP9Ej3G1YL7Hvc27ghBJ
knx/G8GDxd4mP1oiKLQ69cFeK5TA5Vicu7k5SDyPlZMzJ57YBQQbsm04B8KKqREp
KK3mj8yhDX+u4H09K5bgPRI9hcG3Zc16SbTaYVuu+TDjSFjv34uINi/Ti1kUGcTk
TB0H8hpFeXsWehxw+431IqxDng76v6VnZvesF/u4F3dmaX710Rh1hw0Ow0ie0YzY
dwi6nSYhqHM3WHZmCvik9YAjO9YRVz63PHr2Eydiqk0JKI2qDvK2icaSq7O1ygNo
xWQFFhYf6FWfvwMP5yJAmAn++1LfumVTZRzwFWMBHSztvaYm1fGQGgfm927iDBRL
3v1tugsE3Wti1enVr+tYlvXfk682A/Emr29N3WDsRQM654H5UrXm57twKt1nv++X
ZvS3xGYOiZDoYLyDTQMR2YXQT9o+LigVNGNNUOICQUX04XHLmtSEyiLWzwbiziXf
I2vV8RrSJrdLCC0o7QM5CqfiFkeY21Yi6EQocwn4eDRdOSp68H3S+6p+5N799Jfb
sNmh+Ed2n0XK4+fCCMRobV6+ukLd8ORyYs4yxJSDPfVDreF1n9oRWtuQ7AN3aZq6
WWeF5yyFKL1DWCrcw+jxwBUkB+GqiW/DIxz57DM6QpAqQF8ZPvr1YysLjFZxi0+B
hXvsm/ppAnLVnHuAWdYkSDss/RrGslq25DLSQ3srJHY1nPk+HrfIccxPw5HlKD0o
+/lwAWbI8mzfRC5DO42DS+mhtLFf5RXtzO+yFWqRGmbFLa5/pIgnNFKTzy1VP/RV
NHYkXC+oEsfGtjB2JFLoyZ28fhNvRO6+XNxAqBkFI4NG7pnG69WZLNu80OmHoOsx
HMI+NUdsMOIj0/tk4zQy0zojRvku8YuZELvwMqwitTtjXb5GN/vFzaHgnfElzJVC
NmNZ0dzJj7g0QI4QSWo0fEf3+2wvkSOKR72KxehZYEQLebcNtU/eYq81UaTf/Qrr
xbpXDQu8KsE9vIIrYH/hc2TS2BfJRJZA12ugShT0HzNTb5B2j5Kh1qd6YWM+kzuY
Uqphj5/iHOxN9vCjNhsPHopKzBkHh4MY53ioSbAJJlOtmC6GECBo0nsftK8aszal
A6/5cMdD9nN0PiQCf2RvFpz3mTR1yfYtgToC2Yx1VGnFrVjbkEvBqyewRZE4Aigm
Ju/ihwH+lsJ6e9QgazBQThksOmcymmd3o9zzvLTZYAcEM8mOx8n2HABxIYwK0vhw
w0ev7uiqYktdfjsj6Hp9m70mkVubLb+609dBwkswHdL1tOWvSezlUtkQsOq1z94c
TdOOc8P1+aSudnlWvEASGKENo2kYJ/87JP/6Ep33SL6ATZrWqXNg/hcFp5bpXM+O
b0PkFIICYFxjrvEpA/xLtDtrZhI9eZIKPOvzioQWLZg033CjulrO8TVJynf7Dt8l
hrhl9yLS5s20tX07/bsoAUfag9S+D6w4TSCwKolm4DU62n2gntg0evistxB3POtm
dNsMubKdaeyzqyMO7mLkTiqp9DJ/MOM1dSgNqx3yrPoofV/jytlYyIYWQZfhtgEm
bHUY+NKkUMg6jhy5P2inQGR+axK7WtPrqsd1qzPS79rNQNQ0wcWqAzsOzCCGPyOd
2VdT8Oh3tOBfAe2zcPtDyje3LWuoTSPLGnIG23RmcCpOB10Dh82b8l9uMDkewPUL
z4bZfJrw1zHc0K3+erMBliVbDwwTTehO7UhXijKPQoX0xQmq7TKzTS2WmkeW61SR
gabJV9StBWVuTW32DQgDyRHeSRKMUY9se6ZPH0V1O5XNxhqoJU/2umg27QeT5tdB
BIdmC/HwG9qTsCL7qIGtULen6gb7Je9Ap24JLsiA2vY1mT9k6w28TzWgI0+Ehhse
98ai75ovHbN9QSyMiUhjvx1/5DfVZePS3G8PTFRG7/jzB0GeJuvdYpooCSkTxNxu
7H4I9EpWPFoo5Xmuodzr8P1s6V7zpCHMbYU4GhhtIKpoaOJI1J+KTK7OSvn0eqAq
Wokkcolt8yFFcBg/fiUd60ah6u6qYAuLOORRsFzVea19blsNjNLJXBxEpoPVwQk6
sXkGrNIB5/hFY/NNdH3I9hJ/mYgQWSsAglN2k+tpiGSj5B28OkyuNoVH0vTBeZyC
54fxo/jX6Ceh2fU+oVlzCRWRp899XRLHD1rMX+9eJcfOhlScNEES9Dr9IGFX9mEI
k2U5ax41BVnUT5i8WXtfK7Fvqogu/6wHLajbaLS9ynzR32+ScHRmh3yXqynneA+j
m4yLMic6Po0e7vnrXvYdSALVMwPvxUMVqEuk/KqnAwPPfuNlBk4nTLWDaU1FQpCY
8oZexs8G4MVkvBpsfH9A3eS8V9WI42KgZPLUTPvHsxZsK/GN9Wj9nT3Z/y6JR1CR
b1sM+XgpaabPdEVjSWl47kTyhsGjh7/YWzieeWi4H68=
`protect END_PROTECTED
