`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CjSXamHHGfX8jR4R+qVSNl9j63ZLxmRekiTS9e86KYrD9fcDYRepfb5+SdRfjXOw
hLoRUdottTaVrt0NgcMZhFb9inX1IvszeL2koxwd+7XxZ54W+1xRp0OLZcVsuu88
INfl7kKTs9fQk67lqwoO54wN+HCceatV7EWq0SzkkMM2uxvac+yl1308Cz+ZN/Nx
Rj40cfl1R891fkGv7D+bxcaHN1JN9ONQAq5BYrXcaxAZdM5iQ98C9ExDOhH6MDb1
aUwqZYXTRcWJFDi8qOZvXLJKaqqdVqktSVG2F/OYj7uSpreLZ4q725GPjcJMO86b
qZ3cJOQLpM63Ed81MdSE+1eRerlH1SBRsqGpKz9M9rPmJIBHW9gxwe8oTD1SAANf
sM3THMjwr6Q18mSDTsgtFg1yN8yDef9DsIdEarMRSSZZr+ewR6OOjKA7TM/aE0wB
e8J7hpBhq2Zii3EZzCTVt2bvaeGofmgKvzp1WMkVo8nfx1kB9Wg97JcsZo9CXThg
zmv78Kdkh9itaqk4i3eJ7icoS60rgkqnmxMstqvsGK2e6rXXc3e2FKTIE/d8tu1s
X0H7j1Auovs/HfOoAz467sVHD5tUA4DuNTC9mrOdKdpMu/gF5OqtbMs7+r9+oqnv
X7VUMyWYqAjqL37cI/QswfCXrGhha4PRmh1EN2SrkCRzks72Cv5GPzKkxxHVJvo6
D5tFAD5b/xLuLeYBCVsiEMfFNPxO2w5Nah4FAk/lwui7/hnmBf/KVvS2a62oHRta
XZxdM+hRwXLFMSD/Y5PC2A6Ax6Perqsx4zEsz1bILqpcvtlm7VoMMhtOg5rk+igl
O3ld/bjsklELHYGV+BIdWMkD2gvtDGIhKgeIkDiNfgtOd8txlKRjLf7t2wovm5T/
ewj04yBtGaefkpigOGS5LwwLiKP+fz371zZ5V0vy7YmPA+pNxiRSWjsqMFuRbX9A
cfITxTf8HHKhIDmqtkge/lQbmoK0VZG+3W3cll88NmdKbKYoByFGv37i004bthtC
M8PT/o24LSRG0F6bGr/zxwnx58amPntwB17AEwWeGTIyHFAYzpbihh3p23TInsET
0mLTuumW47B/j/L56DIcofNXiLylFzvgOW2H0I3D3YvNoSBkaDjWXzXItRD8zY8x
U3qpJ0TY77v3nfwArWg9doizZx1yWYfOgn/2eapNO2J/63Me2UNSpbsYGRg5UD2d
YImk4lRSgMXjDm+2kRE4SWhm/b4FMvpd1nHJLML5Gi5r4GYcpayhQTA8JskjqYnB
8rd38/yP93C3oAJ36MjzhqOiK8gQToeSV4Z88Iuxeju7XcY54qQdYeZ8IcBUTMZh
wMCf6AK2o1/zD6Op/4/TxcBSn0g7K01M4Vdg3IQCyyC/N4jE7BUKkA9uR3rw2K2X
jFUQWB2HoqgT87irHztBNr5Mdr1F90Kfo/hnK/5hR6pWny/nHzCigNFz5Yd3Ag+y
4tPFlVa4JEkDeupgCPK6JSABhHl2ZdR8SCeEMOoIuZg0nfwmF9ZZ+FS39MytauNO
LzLTZ6Ll9Z3m6FmR2xZgwQ==
`protect END_PROTECTED
