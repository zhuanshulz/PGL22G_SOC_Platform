`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jjfVlhGFngzN6NVP6+GrZK4ll6ySzRD7Fz1nZzCc16okkNamaGCAL3n+TtvlEbiR
Ip+8sTqzOouZZNeAwvDsV6Sk+hNG8ayeZMok0db9b2AiFLiAB135FsSiXNz1sCvX
SGId3ll7rEXt8Fq+Goz7ospt9NmVv/Fn/eeAUrufFbRejxNoiYszdWeLd8Mm6+gm
NRTzXJS/wemxA9QffE5D4O2KLExvjw5x2BJjxYfq9pfKKxgf+DRmwsfuTt424QuS
I+cql5idf0Asj+jnd3vWkRz8vppL8T+dQuwwsfzZnP763cZcd+i+mPAwBz1xBqoh
BRUk6sdOMx92GzPGYtb5KGKjSFP0p6B/TFWa+8nAya7x0z99TNdWbuLRo5z4vCOW
A7KUDwubykEkSna/Pg0ITP9+hNfA2ig4b0JfJUtu51+bKFFtHM4zw26i94h97gBP
LXhwGaaiI5w0dvEy8y+TJAPoLvoMJwNys9PWhbwzMyU8dPJmy2SzKeF37boe9fpM
+K5XMTjA0sVnLVBygc2M1Glf/NZwm845YUmlWrjALtm+29O0bVWoMdl+ZArM9Ugb
wsgG4DODqrsdsrjGXJlsuAVmBKvqU4uxAPr3natMlRUeR2k+FpfYFGSw3Rqj3/od
gyG2QczUpsYLfQ1g53tId2URzvOP78Y5XMjkyOtmkYeIhOP5cC9oxVlDsBD4UPJR
+vO2J1Swq24XrZRSmk+NnYLIBk4LO1iuwa1xc2OLBVUx8HRLs1A2KbGHcbPt5aje
TvIz4PBc9mMamIPBOHWFk9Ssth2OF6bq/BzbXvxCT2PbYxh0A3v7RBydgOqN7+aH
3oOLQz5+kkpXn0sHvvrQnQkXicQ5fbQG5gZKj0LZB3TROEo6970Hzgg7+bSe+Ql6
K6VcKCjckIDqBkMXEDdRb1T+JewbxenQr5j3Epvuo3XCIbY76D8bVOg1xxgaRDu7
HeZWtm778n7mimVarv81mwMhQvH7lI9T1Zx4LaYRUFI=
`protect END_PROTECTED
