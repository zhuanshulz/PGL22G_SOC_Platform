`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
82Mq3Q0NGFKM3qtbcSKV7JoVNarQHD309C70yptr7A/ywpu1BFtbIKs3zIprgxzd
K8Lx6I3su1acIqndxB9FCQ2HEoFLXTsCUhtR6OgwclNwSyDuRJVU8P4MPehciLQF
L2hk7a4l0ZdQf+TkFvRGq392iBtecZi+KrsilwDEKuwc0iB3VYC1BX3uJTQrm9Oi
bat8ZWBA9Sg9MQZMkiiddwEyiXlxweo41UaMYR/wvxqV/48s+pe57bcT0UHo+jFF
qkYjLHtwE4z5uEVNsFn53/F5xY6moV2L4QJ8ug0EJjOjwtJaPDNwUr7+QeKI2WkK
rGGsOE0/bXQDQXij1c3fXhSYcbHIvPrN8KVGcKFWCmiwbWUhaHBFTF/EFiHOMl4b
hbNTmeF9KgDNdopbGZ6b2t5skY/ZFAmD3wNJ2OEGT797J2mQ1l58kTzhRFKgqy7m
XBL4uc67XhrhI8L3wzBwe2kM9Ilq0xbNJRcIDKtHS0so0mgt8tWsaE2ChUn8rRYT
C7Y44/fBAG+mAQV0cb876Qv7di8KQfUTx0p/+F9TZDTaGrulqgc8IxyIvTMo69Cr
fxlKkQCXBLI6LWpQ9rjFkujQl1oOafNLwNO9gx8xtxO04vmlNkStlKtQrjs2v6O2
potCVwRuUUWnDl3b7SDSyGWO9ofckpJDIzNIeROmNtt8x0m6Lxs1/OndIfWp7+2/
QYifJk9oEMlm14UsI0MVTRrOrMCBZ23uDqsHFfT1THBKW/a6XHnnKw+Q9TG1dWD9
DhIm4fArrhZaf706W8SgvkUJE+aD/JTX2Lypqgyox7eTNqJpvRc+IF+0Gj2KtvEM
n0MeXQtNuZ7hRCDxPsmklA9GtRIgV2hevK3QSvesKgSNfBMyN6Q2t84wQjcc+q5u
KkEcmc7MMY1T5Z59YhkC/tUS2r3k7uTV2BewaYWnuutHk5Hab3AoqAqJwTTqZWs4
p6i9D/poGfYpGS5hW1O8r9p7MmZ91Uk3X80n5TEp4J8nKvPaDX7EJaB1BGvfYKwL
Mdf2O18KRma+lrd+2JR4jg+84y7Yle7irP9oFRlNwmh1biijz8Z+1JsOlmZ19F4o
z5UJsKwWp1TRS1cWIEIKRR7KlYL1NK3BtfWgHuivlLJuKwGRpbsvQeAsRIluoxuz
8oKgLzrIUCiU7oSll9F+LLCh28rjQLmtE7do87ZLOBxj6T1LaxT+K1Ff8hpHcIZB
EbzuReyBvtfPghUeGKDc2iZ6DG4A4uLgeZ6c9+sxSqwRj7F9vY9mrEPKHEONrXu2
dXm4JiG8UBc8kRlDiA6L7Zxww3asYjPQSWcWcQO8PABC8KYsaOISWExHQSkAhmF+
++xyZ93nr0JezyQAJMR7IgTPmAIkR3xazW5op07FpZup34wb+DCRUeJwUpSdc4Sg
qRk6VUo/H3eW7SqOghWtWwBXmSDbMP3sbqGZgGSxeodD6MOkRl+s1wKJ2cvFWBBt
X3cYDOIZ+seRzTjJCg2no5Gz38gfr/Dovt6mZaqtynXI22PcalxEwibAq/H6WOZk
rLYJSTLAsnpUhwuBXcrDOpPd+oX6lN7eEX0T0oFkBhLOQoh2AqhdSSRhdrjButOy
6trPhT1ME89recIAYMEFVKBTFXU7v7xst/wQ84+JOliQDIhzQkpDIQRYVYeNtBpl
xwZ5E3twbshwzuMVkvFWhJxP7mbinpCQF+I1iFd01e9Z5WTFM7/6X50UqY+1q16F
lU7JG+Xamsaie2pklHiIdpxjnlabKcgnXmjSIDq31jVnchvjYcMC0XBgwOC0lRl7
X9TW49CfM5Is0g4x0fq0k3EYiD/OP2gTI8eEkiewusjgheCVBhgT6kvn4QHKFyIo
uqm2grUHRMEJqXAxKDYz5qzUqaxKGZqxjqiWcUMCWFlni3QJY7gX/VLBpxGAoL1q
QhcXpTPvA6IiebQqt/PHjq88DiXVOAZBdPD8S5qp8XpPFL+or7IwwJwe45KvFLlT
v9wgIqvJKBbunsy4sUZsz9yak6vn2Xp8I6fYh59DuyHtwgTDSwIJzw4hBdp7nkTH
CljXPnzL9HCd3UD0xFTHCS3CQiQW6yexi7To7Z32ecApQJpEZhRoLs2k+vu7z5GK
zwnv8bW8EwVz/9yEbMyZcs8QZXTeiM8dljNN/vibvWgtyiP0AkVqhbLNy8deJLgD
TKAvxGVruXzoqDIbIMyFQ6stuMYJ+hrUrem4P1KpRZiskZmF8JKOMTXbvarMUyTe
9id9qVdqtyUjeXCxnHVLgEUFN6JEIXXxssb/12Rxl4dpCppnL6Lc39Y54I9mvLtI
T/9c3F3N8lCCn1vD/+x95Y9BeUGz81TQr67zhywwfGkHTgTwL6rulQ5+dD7PdlxR
bhS7uzdRGgFODXQe7bWwaKn2Q/2JnfBaR39oHtrTSgZOW2CLB7tf19iTkqQdnTxq
uuXWBPWMuIe/zQZrmudcHTidobGmm7jFlUXgeEQDNsEEXjg5V6mSLnEoG8JOz5Xt
2Q1WtgHuCWkci/k968UH2A/hIb7WGEQrstCLdc5EFGzUenMq50ehfZpYY7TnAVZr
qmOGJ84AP5uYRp3lR6SGxv6Lx22Vf73/73olGgN6ttUIgaH7WWognwuURajDfX72
/ofczN4tgPPw5dfJuuG7zW+POU6gkPpiS9S8QCdiDLW6lSBs7iaWqCQi2RRHNQTA
VwoCRo3i2pEf7Kukk2Acp3XRH/9UItS+vEMc+TE7TVpbNPEh2gEPqA62IR2wYkI3
vcFPWQhmrltNy/zG708fwQRd7pWDTOaJrzj334XqD6tVKubI/CVeqrLxOBF8aYFf
1Ht0VzbdrVoVdffkLvEzxNatwfnmv2K3InsxOy1Xg5DLQCn/2g0s7yWEs/QOOqDx
U4XsguQ6H0AF+6pw6mVh8r3WMgxYVmo9nJ0VtPW22XHc7Ur3zpMYpRWeBkAuzuzS
6EbSeMrX/puZC0uj1e1loxqP2h0cnKIHwlF/XWoimRyjEHlWgUoGNgW4ZMuhpxvZ
FhVRgp+gzzgf3Jr5GoHvnOBd37N+RXTkOxxLdOGpMFU9pUk3AwW1fD1sHBJaHNyM
9dl1fTtSQkJFI6C0+E3N3ra4Av7doQKJOs/1z7lCzfYDxzk+Ky2UwyaUmOUAIqzy
AZCpvuPSeQaiUrWGwFgTUM/xFkJGnhOmtu+qn1Rxv5Y8nci+9GjPqMh8oxxYBeIn
CiFMcGhHzohKJCQ1RraThA8cfRGe1v8DGF0SXQQV5iCMe8kbNpysfaQlaJ9XlO1T
r1HmEvXhXQSpEESndH7+HemG1rPd13E3/snTn4PZbv8+qJQ4uQ5BCO33JCHyWvIX
V8OTXVOt6VkhUAzG6CvYq5xf+gUKpxhUnThYkIk4VBwuMOLpawTdUM3m4sSAqPod
NA+43M+pRigaSCEKdvOwXWbiMdtp9q5udVxQ2Mjg5NYV8n6qGHy/HqAf55x7Tgfo
NmBp2ZIMFrCauqVFzCEUE2SjhqT/BWwJSNMnIPylESr343y98yswJCu4A+jpMv/D
VhR0c96RsCdB7lOAXK2TDAyzxmxAgWrSL7dLO3OzSKkaArw21wElOQBNYJGrwabk
F5L3Lr9JG0Q4wBBfKKj66oKMAyEJekEpxnLTg/oyDC/ticF0niWS23lVZ2wgtwLG
84RpLrnWVo+2ir55AaLkdGFQTxekKH12INoS+p8QS0c86WfMA9iUXsts3G7kn7L+
0UQHK+pMu3NcCor0QMo1ux1EmSiZyk1ceZgZvTqkEeTJKleZkbzDZ9dNqu9L6ir4
u3o9zxM3oP9H9hMrHAcmLi1yEt5+DSjXHH0sY0cldaQicj/btFqc867LTgmN1juL
FdclPtYNjSIPT2THBfEUD8OChB4ItQVDd3pPOY5uTdm7Kt2kbd4yMg0xg29wmcPi
0711Ks6W00mXyGRqOeTtXJEzYAeag0IFejCnrjcbZCtHcEfErKcNvEfOnhZNr01/
F4azMjpT5ggGHuY5E5Z3nalWi7Tkh00QRL9459Cx3KkmxseBm2Hnt8w9OMLGntwu
JixUuWV7Y1Ug6ZM2BG9v/V6uZ8Ir2UcKyTtQ9S0zQdfKLTD70++5KhERMQNc59Su
ZVasXY/br3mcmgDITdcWtPImSQtt52u1hdQimgV2LCJUE2HKnux6EnhPPOHzGBX4
6E2q6Oa6MDQ+s9QKmwYn8/H+EpuGAEVAwZ/dp4KOmIPBNap2IQitp2e0HbLyawYG
X/MJybvvaeabcJLuDIDtgP6ZKGZO7/BImATopZ9FwxayRadoMd26yc5hVsIlzWB3
Dm69hXRy3BqwlYTRhEcsvm1mVYWVIFZZ78JGo2mEOWptAFqFvW4SGiHJ1safQz0V
M39IOMXjw2rn6/sSM6AcKEADU2WcrIE+Vzip/WUhRM11Cqn6hV2pkuxZFKmYQwZ7
Z57fr/VpOpD3NLhlWS8cs8fpf3gC26+0P/9XthNplKYtIj5zvSUo+wwPxSmC9HEp
pxiRF9rY/8QTiCLr2Xck5rZLzgAxW5F3Ijf6wTQvvfMLu9+87iFQ8fuP+543aqsD
3oRoRWTGZG6v79RZK2v+uQ1nQqwK0hPD60h3fHJ49qkPyRPXm8vgVYQ3tVQmJxCf
Ke6H/yJ6zfq5cs/v2f+iyL5aQVXRNmhP6xCFxmEzxbS6VqTXVgMEe4HnauRxFb+H
6zzOW8NH/XqaoJKtqWT/uGaCHcxpGeIrCQsYZd852xCXDcy2C9bLOPK+LhI8X4JV
lAdm0z4tztDNQyl5e7oWjHLHXyjiZUnv+uTKEKpyKLGAQj3orD/cMVi9IlbI+XUE
7GPg7ZRPd8Pfo2EGtiARhad364Ai3trLzPSbr8vrSy8fcWd+DzEPG0Y56LEIIftq
LPbGfT1kXXH1G1CCvzHjjtDPsUs+c/gGaApRjt7jqxnX0PYLc2SI4o3yq+F4K/uf
XAxRgJ5FLkFoZaaHt3bLJ+Z/VbCK1UTs+wvYoIk7Gheu5R07dcCW7FZisq4C2RPO
K2ZWLSopIKqZWJhqkRNa3A3pA5mR+RSsh+KX/FOGW2AUrerEfhPIm63Gi18Y+8GL
v2oVEx3AvAQ+H/3Wik988hUToctqKq31Cx74P13bhpqs1h4+4we7TdwzcCKkKnWS
xJii0PtUMlGKO5LEiL3IS8j1VC9uCg8HYr0OWopn9INdITCyqMDiACGDEcUeqZXt
3hzKZZm6vzh+aCHJc+48OI6NaT6Ezbs4F10GInS+XTUXJiuW5iANGdCydhdeEyBm
7OpyJ6TiZxgIWT/R5SVkqlYtORL2lzvlToLbCFDUlawWfCbrG9tO87F1jIaHk7F8
83AU3XNCYahnQXO1HKp00NY+IgcgNhhUOVPLqCQ24HQmN0gtTjxBsOomspu/L2KV
jE8Q6hUNCqhgturu0kXaec+fNL2MUS1vXFws3dQoOa+SsZQ4tC7H9Qm405caHDmT
+Z43LDhgSGwwimVvvw9NUwHxmp1+6G8W00ZM9hXo9TW9XCfPFi4HQQoMiL/mA+XK
flBuSlNtx5p7X6FzLEV3k4Wn9SRFEAvly+q9cjhyqrqA/3ZIteLmcF+cYVHWt5rn
LvoI2D5mu/QD1seq6xI4JX2yD8L6I/H5IvvSh6r5oKRfESIJGo5+SPtH+850dpTP
KTbgn6PiLRrBRvfTcS952Zi0TVZbhO3ql077f3CI0ojLjt7QSphDV0ZTDy/jp8yG
mD4PnEykWPNNKOvDZhFRHfi93Rbu74UYtJ57JbS9ZUttH0fRLEwYOzttCBo2jXMq
1DtmO6LGhAwSlK7HKpvnEFMGl2IezHSz0wSBoukxMGcNpNoCFJGGkjzO/kP7GePx
T45MUbmskbjEG5321NWt1UXfaMWYK/25BEhaDhZGtq/XwJUVP15HYt92YL1Wp877
TPN04nh3RSeEZ4A/a8HNq3aIVHkiNukmn/RRSVSpYFhYHotXmfw4wzVxFfkKMJZR
4yLd4NWqdA0OpRBAekd9rjEVQMW8fLBRNdp1N1qI4/+kYFjT4AkeH6Axnirpzf22
ExwT4VsrsnGMsjDkgDkwlnbg7UADa+72hyBHWQ2mp/EI8jyE+d5nXM6T093cc9wX
EQ7LUmkj+c4IHiTV7Epvi//zoB9r+IaoN/lgAQz1eWN3hfHew/SwDixeyYd36qUF
ap+2/Ln4VcGd34a4UTjha7gK61PgfYsGeDwGBDgysqCh39QfwnzmFKDP7vQ0/l/0
q9FNZguOaQ6v0j7BNYnvpP5lSTTiapGb+hhIfA2VZ3PQD4gKR7EfkBrDVSmN4c4z
sRog4yONWM/OI7vQjC+egOvQwifNu8X3J8zW1M5UUg56zppQ9/uD+Ri2n391Aqld
4Tsv0JgXTIWStDPANYLNpaSgcMhK7DsHlBsovf/tw01KRelrdGe4ebR+ZzghRTz3
9WHLVlsVan2pKxEvWe/VG4gV/mwmf3IuANiHW9CuTLLJDLlTX08CJZpVYxpn8kQ/
+9FhfHkDTahj119+YA1mU9Yt5O7Mtmnr5slMZWxdNFJbokeTJuMIy7ux6QJOxD2y
nB5RGyftuwODykidoexaJZIKtWd8vaBgNfU6PtriUsPH3F0NDxUgjEEaQ3N7TTAS
e1vFa2qyQtYsFhFMz6hUeJg+iet5MAk5X3PAS01x99ds+DaFDv4fzkwXSx7hu0UO
IicvEdIxHewJybUbe/iaV7F+Eb7nWHqq88xccv564VTUEfDWTMK/sZjW78P3MZSf
hP9Mgi/UdRMpbzPZJS7SwGgqnl6IoF1tOm3BU/JsvQSsDU43+NOtJDOrTmR4cZQy
yCm4Xf1o/Kox9Qb/29WIoBi/beVovas5kLbDAbk0vhSe/ECHZyRuud/WRk5ylkYf
zGDkt5ssepZrQ2zEGw5IOulEktzs5LYcVUvoaSWiwlHhWcAlAgUn5kko07vPDxKw
vtB2QuZZrsOyTRSoc70tw2+p7R/JiHlKBD1zJVhGQ1zpD0UAjUk0k5C6sbjt1xb/
v1y4qGInQin/+YDez76MVR0fwHljaSGd2ZcQWP2eHjvQLa/eRQdOwR3/VllTeVFo
QUSPGjpxD3IoR/7s2grlcB+JO8iEnb+NkPwYLmtYzyn5U+YA+C6jmI9G2nk9lXgc
h1LF9TRhgFx+vPj306t1ydIlmZEPmidrWTB/f03EoiHzT8WuguCtHXRU3PnUszRm
tW6XZVpMtzPJPRXxD5Zq4+q//EkxXEsFL/Ot6QbUtR4V5gjbY8npNgKW7P74rTv9
mpXXupXA8PpGhWcWXxLlm7uumVj9CFOksSgpelWi/5n5md6cO0VK//2a/tUI2rw5
q/Y6Hxhr/fdwRuqCGAI+qnLokkTfmeJkoEDW870xV6eYl29W6gUe7y0Yx0M8wzKO
Kd5UqyT1y4Yj3YIpXA5H8Y62faryts0WfZ9b+E71p4ob/9BsuqGq7R5vgZsbBHgC
kHZFUL2AZe0yYg/DzGhymBQnOp5fZW9rTaoSKHeYDqJQ20qiXlqkSQhnuHGpQDiW
ewCTytINyx8nJQj+PvdyulYF3QyJE2KZvKiABm86CnXTojzFGytQLymhh01V0t3Q
MjUZAYYmE02Otw1/I23wWDiCqzCf15AhrzZNgJqlVnu8csUOPvkEOr/NWsfnzg9X
2Z+JcMV2bAHCAEZ/CUWzAGwx4tcN/bD1MzyXyRTr1Thjypx4WX6L4MdgEp7p/ZOi
vEaRJrL/yF92zVjVsS8DJWmTM/XaD8rVYfMXUTqnTL0rEbZHUetk9Jy8oRRCxwdi
1DuC2e0sB389CfHygxY1zSVZMBUtO2oLm/P9GzemFHEbjUDm5HGWOFrdf5s8bBn/
eJUk/sq1J78Qxv55I78Lu6Zd5ubyoknlKaruIT1C5JkEvykerHN9FJ3SndiKeJ1p
ZQ3VXt2Iy6Cc5+oNwyVA/PElYki+s/2zeBvFZHVx1tRenCVHEG0SRnvZmSY9l7XT
h54PfR9GUtjD2xvULVoJMzWB7KkCV9kC6lTDysL7A0Jdleg77PvV4jPeGjD/Nti2
871PMcxdlYUhv5b2x8k6jKejqXXF542++6xbVZC4dkenI9EMEXra7dwHRE+Lpa2M
WudXRcO58k01dItxwbKtvitc4NjCL67TBP7hng0UUQmXB9cIJ/F7Omy0YI/3hRVa
FZEnvM5HIjhQBs2WZIEsrobXibgfkDkiyim2kPwdeD+4fcU1XMH02kQYFQoLE0FU
8nUfXMiuTUKXWfLl5c45PQVRjGqaWgQeeHHHFIizuBd7SuIbonEC3NPBULF93ky/
aIbo9f/Mzdyg7ARFVSmRaGn3GIRpatKJFwavCigJpdl9U9ukRXVf06VWnTFW/hjV
8TEyEt7uL2JnhdzT9gzPadlNnj+mb1a83BG3kBIFO/VGgpMB8UKQWxqFlbaNp4Gc
b51SlszGVzC8CtHBV2db1CMMC6DiVut90Ke5sj+T6nGAVf6EBd9gVKHUU02cRPAg
7xmp9k8eNztyNvy4ciy205Kji4ZOaQ/1AoO+IqFhgEl5n5VG+6O9+kVOVfF9SV84
8QS5s6AhGKFv9gIMFnEe8c5eI2Fhg8DgfHkhxFn3QLLYW1dDpeCFLa30X0fxnIsV
yA2aRIKERWMvMGaXAJxo59V4YcZ1j8PnhFR34qztxPlMDFbXWhWu/Fkhr1s8JWh2
QTtG+6KR0fEcUXb1QuUEKIxEwa3AT9qo3tTzs4mXpm8CwLBN4fqgIi4kXEHrWdZ7
Cluv1Yu0eNXjK6i1VMT1nLJYPufU80n7Jqdd747HtRtxjU2mzKaoMNtld8bK9r/Q
twkL4mfiSYUCpLoZ+x3caZSMrHSttxQfK7zyw4itgtAy6YcrlHxZHqqzaCxsQmKS
7i49ErbcDi24V2uc9G4xO99vLOQeL4im97J07ctpwd/iJQ5R72cNkuo5Be2zXvob
juKxmo7hJwiHcdVFPxwIVjCymH4Xqj7bgZl5CCBL8YLFRxYhFi3YcUIV2sldTiby
5siAs5hNE8FI/agOT5R3t+idv5Khw+xvMZ4pb8xRu6CYytVcsN4ahx80/w6tjWt0
P+pealdOoavrCCy7s/K1gmNttavJ2UFEyEi2/WDAuxiFLhUET63+JzMdiWFHwSo1
A3UCJ9ncoxm1TdwdFpP2XVQDvvQr+Jt9MUsomsztB0RPxf4EmzPQP8INznJHA328
53Jp6lZgojdKGSjXikNPn+lg8SQx+6kxLv/uwx+8JaIFXM/QVcMaLpTNQz9O5pHu
kb1KSQwcCfBopmRHjOBS/YYef59S9Oxo8c+GWi1rQ8kpCOV/hO3TNQ1HZO0cdWxL
tOnHmozFYz6/jFtqOAToW62e7NjNl8CrTVvIYx47iInDEkN9eTPqL45I9u8XAfKa
uKMtS44IajNjZ8vydiUotYfjJSLHWCd1DGF3UCj9g1qvYDh1e98SJwx5WjPoNucv
ZawHJdYSuMX5LnvihhpuM4pskSvvP5nBWtPQziiiblq8CsyfvJhHfBm1C+rQMj1B
cfTRBoXfrcy8ypnNfRsgDA96KezkNgMLqWrXRZhFC9mSpnuOQZz462KaRfE5vFir
GKmxJM2snzssR+lEepB5g4onvw9iocem9EH8WEF4cu3OyVj4BFAMMlZCV30ucLEb
sjsWHSAzaK7V/uoGimyCIn2Qjf9rIyEF9YWfIyZTHY1+uuYuJmZrPiOXdTThP48h
F8MNLqac+4rXTP9cQdlRemsuFk1eNWypInFu91fGhsB4iY1EjjBEAxX1D+shBeJU
CvYAPGqrMOfGu5hNS0aZSrD3vvuAxOKGYDMiHbAaKzBl0pOZiaRpwDc+Irg1JkvY
1thESIQx7Z4TVW/09Vm4xH4vCNRB1ADIf+GU+P9Tl11iNgNG1OrPgwgNU1CtEZZm
qxE2VNksoQjOEX3xhTPbd4PtBVoAqV5ggz7uCv3fOiu/f2aPcebj8ccpsiXDT5eQ
wdI8TG7HCtWS97Fb0+gO7jDoS7zSAg+1wIQYg3/PtAA0DyMYs5h1m2tdH/gWYmXT
0icgi+jgOXisAz84aVvsyGS8BY2xehDq4oztGGeIQj3NxOODGhrIfcQpcqGF3ERK
xGFXt5EamkCw6ZwAFQXPcrpP5SDapsXc9VsMoKCJMATDNR3Is3PyDNZT3WeVNHaZ
MaS9QCKzI1roLMGylLoGa+B1IahUH8CFBgeu6qUiXGn3gdzygAhjP4BEcshu/Nt1
l5/fZt5UrAP2gSFJIg1esSd8RpTyjDOvdOmdPXw4Q6r7HW/x71BjDecU2tVy0USk
0zKe4Pe7Q1H2+3XnQNxT1RDvnPQS9TZ/WZOItAWegKEXBSHEY6uFcS6TJF955QSx
+d79/j6abQ8a81XBIe/e50XGamCSJ+4aO/U8IXnDpD+v0UNVLHqnugAgOdr0AfKT
1blEQ5uwQ8tAgIcy+YZrkJICzrFigQAJNLBWCpXOBVGNICBTYuZBtOtWOmdudPJf
lR0x7mbJv8ZRg1FDbqo+/cORnvi0VuWXaMoiHg7Ukp4PZy0Lb+ry8PNmphVnL7V7
UQIgZWa2JmvWdaYSSa2elbPhzcM2lOI9u9d+CZhT9ZqLpwg522L8NZ5OkRpFzMG6
pYp9nbP9JDPsimDj6itCa9VzSO5jAksU4/XbZkpcM1sK8Bl+7XuzgSrrj2jjjVo0
PeJ7dCZeq2DoucSZ2bxyuLFSkuwKaDBWu4MGd/AjzVlIl4c4D4RJPqCLLzztCcDa
RmtCP06okKn9d38zAldDm5cPaZrkwQ8S9qoqAAMXJQU3UV4nDrCf/LGpDE+I6WqL
1bU5JH6yk0AtYJnP0S88IW5h4dwADTs7qEjqtr3PcnJy9JEOT8DyKPeUwD+Aqjb8
AtuCyEwtCb2QPrup3MWS0JO1yFpEnkx7sYRVDcH6tTlizWeHCOGibfA+HUVK59Ry
dCVa+Fou4CoFxrqQg8Yhvha1bDq/pxT0MKA1AurCJOI/Z7fo4ENgRWorK+MaRvdy
jmIhxH7/gize17bNEN547A2TiMbxKhxDrun3Z0xIRGF2s2aepOnruP1DhAWrGbXX
cExyqZohzggvUfpsYdAG+4vAnaE44GCPUO/cnh6zRBiKgdbjqXG3zqUP3sHHmxui
uisio1HRYycOKxyy4/Iklya6TOcxb+nWJwbF84FPBvnpubGGhGrZXvGsSjBvuF/w
JHYmCSqKW7VJ8ZoI6wB0mWw/hNMEf5a9QjO803aVj10udCyHRQh3GjnG9gHPrXtN
kqKpfNUWCarI5NXpJHJdZaKyFn6XhmsHrDKzcnH/5f1eGlLGMFDLUfG4gc+wf187
x+r1gj8RnwSwLNAZUfh+Ck8RLh2eV3ulucxn61oqjouCyBZFyowoRHE56A76YBkI
if4MCcAY4HSqrq/SLQ1lgR8Ycu8X3eJyFKN0TfLdFw3wdwdtjIyY0utzSvFlN/mI
Ftv26ifheWBT8+USpTCviDc+LLF+fgCtyB/5HLgC/suFhZcAAjB1E/iaTD6cq22R
ABFzA0HpdWp2IA4nuabTx4tHP7QQrEOHOkeC58Nj/XsOyyGksNwpJDXZHFsMm0gL
PLvlSMZeXQmrvKuaJFyuHFhBYpoFBVRFrR5aZZakXjfeoGIDlxI+pT8fVHccQhee
AM2j9d7KxY04USmcGELrq9eQOTOwptzWW0Po2JvA5Qp+4lLLNiATOTA0qWwG1QTc
aXdbUcxlTJxCGCNEFidX9Wm7/CpwKi6IUEOZzK8kR8BTn9yq6qGqq6dmZyI6c6Sq
kkjjGjcdGQX8FbOiOARN4OURa9ui+p1Jccir3AIuEjZUqY2Qmf5lGVqgpNie+Udk
2/Nigob9DPoePTr6b016/odD2thPJb8D6wFIEky0RfuJnEW/qCMkgCNQjBa+QM3a
ECOoiNtZNilRtKCbGqjZAHfuG7JCR9+FHL8s69nTtUHwAeJOjl6WIqJ/PEWou+nH
x3EgqdTmF5v2X71cFjk2I9OfuUXnm2WjUrsbZHXmIVk34vVVBWnzNy0ma0VeRnpM
wKqqKqdBqb68T+wwEU1zmE3LWyvvsXiuFyd9YtJWyzH8yWeC0OG3SSDn9kaJYGEs
gwjCu84gtjSwgS2W99VYPF7ygZeYHWDTmMpQ7xv+BSk8NnbcTmBCH+4MI4Kwdvhh
3XfVWrcXxEom1GAyceRzHsaKorkSnpdqwtq0NE5BB8O7kPq9aEqfV1upSRjshJaF
D7/wxMPAw/UALSlFBucP9T0Vz8udHFxmUzRIb+Bwkj0+ZKhy4i2JR0ax1qf/fum5
HXzUgA6JHAi0q2NhzYlFYvrkFRGK/y3ZnM1IwJqEf4nIDDHRRq02D6jzNMm0Xof4
TsjF+X3hqR87Jvq2wLiYsVtawFEpDXhkj/bi3RBPSqArw34t7D/utaaN5lma9soe
9gxxriR/vfqox9NhdNMFtED69QV6LaTBjJP71u+cZD/jrfP95M7xe5QWUULEgv+2
+bLErU4dhkRmNaY5/SN723AeR+6pjrp03v8dZv/eXBLEQ+OtAGaJ/+Xd8whZfyNk
MDnQ4Nc+vyOvxwO3jAP00oQuyrAsroldCVMY2nOxWci9y0gOJMQArar9wEil8Js8
uJQZbQmr3ay5Q1z5AOo3uCkOu9UfbLepCSINcvnXOWqsuuq7BBw6RTQ+oyFD98mz
bN/Ax5Uy26+nl+Rmzw6FZI2HDlfAT63VdFE21xEkh+AatbkKDyke/FRmAaFulx6V
VLkSEEKX27aqYNQ09dF1gr0KJde5r01nnx6TlerTGIW77jgLd/4l5l8Wnfl3bu6d
rJIlY8S/rwT5bptWi4KmFfBTWULPpyd3tsRVGACQNkmXDZXDui3lAmpQ9JrSP+xi
YlokHdl4MjScqwPPTLZ78XLnlonrUKqEMYINlqXlazVfZx8Rhp9IqtSozQvTZx/F
Jzr85XECZlui+nLY/VQdSv7jDkFOxEnojwHh+5qFI3xyx9sodkl3gakF5+f4jtxn
/6PZqSJrhUo+dJOclcN/9vxAoZ7e0/DR5CF1cJXeMvXjBRbcmRPXjcQFjT9e8U5U
7hk49oKiqeBb9RYorvRKBdG5q9jMjguMgAHXc/x1cS2ER+Sd11bwUCbHiT9brdRb
TTiJ6qvfOqtT9AKMbZceHhAUYV1SM0pKU1B8XB2jyrczLwsb59cZl823pK7fZko3
ag9WbgwyIxrpGkwzsaUWbHpgAM6BwipkFv16dqIGT2NvwO7W4xj2mBK2nJ7+uooZ
bIqUAR0hpLgdILR7Y5d3EUSCzdjHJ+WTDvz6hDz5PiQrg6qvQ6xfT5iY55pTKM1h
QiwCarrF97EyUoAETn1voBRbOVZIaNlBMStGq3hEF7nNQA16fLvTnVrgYi0kZQPW
K3rFOs8tG+8WWWSmDKrUhWL4tuERrEo+e0ItgF1UcIld/2yzxqfvvQd0zZwaCEPp
VxPlmXLHui7SSfziR5Bt9r0t6ntIFvheEhS5fIwFR29Z//CjDOlkcnigDVZ/+RUt
hcc96ZuCpFG4wOUKVKIb+uJpHZMysS4Axys0GmgdwP3TWAM8kpXj/WKw9OqiK2NC
qpR8pguOBjMwxZ4tOyc9gaDnSLpEjN9IJUuOaYARmak9h2jJCvjJiwuREs8KjxGH
4McTATAdAMF3CsiaWyIT6xQ9hTPiLlszPQXd8gKAduHuxtz21666Py3JF6S0cHgq
yBebh7EU1w5L+BH4aG5rt7TFMJGpt+2MVvTDFJ0PZUWt/3okR3xra0JDkbnQwT1Y
YVce8ubSSh7uux3bP+lnxKULwii8CO7KeIOjQFkhnTrihu9PLLrCKxjiAL7B1zfT
luLZOecT5EiDDEI5QzFp6OMf3nPt9Gwm27jlBQYY0ADg9BKOcfhY/EEyfYlLKPk0
BeoTs5hkfWOTL7HKTi5gGNmOCYmap+XoqHfG8VetKFl2D1LvP9sbqOCAZa4KJDu3
erb3T9OeAaqT7p8rZRlCKZ2zm0Daz/bp+W0VRhsTzx1Dfa4uNwxRd/X/jiO5iT3/
qHMiQHNRmI2QIJOk+/wRurYEFEdZ3YBahmRs1IK0bOxohP4gY4P7VOHKpY0DZL1S
ayc397HS2N5WLPSUYe1qctXtjF0QPoFvClRbHQVd/luhxZf1UmGbAuEzxS6+gx9D
mqWs4lPgnezN1npSoc+SVkl0L1k92F/PiERTcqnkNU1pHX+iMeFgOdkqWPT467YS
UJaJPHfTKXNJJMVqCrBCYdyxrs2LdhwP6XF0pp/7CxBeSJ618IZ8stFzzbdOfjg1
A5ilnglRMqL6LjPe2ZwitbaiGPmfwOMFIyrOvQG4nBP1ZHmQo375g7IhzHYBwQE+
a7LrRlEojJS07wAsvVcdPDI0w1EKigeXWritbE8VykOYCo71l/P1MYAbaIFwmapR
03TF8ku4u75826+K8squoBXEkQBia8phXBu977XK/r4V/4GcezMub9+KpKafA7th
UZav74P26pOUKjDFPRBe5QzsGxhl+4hahkO8trHh73wUkZlknD6uHGOFouORHYtt
ixJNVxPd6D0UTL3QoCG+y6zgOg4ar6vmVsjOw7JfRq0pJRJJPMm6EpVGF+zEtwDK
oWuNp3TND8te1V29A7R1W5FJsQ/erQ4JSBPLX7zW4SzSqRygsHbhbrRQnobDvy+x
ayh/suecj1J7VUzOweiS1BpDCQo2ca80yvjIwcQrsdau/Vx5hQn9iTW/8c7yAraF
H7GdiOze2fmDe/e9keQMV6KfmgR+OIcPSFYiiABe61sE93cBOBXE+V2y0QEZM5Yr
69gbUiuWwQ18jOsDjzKlX94Rn8P0CeBUaOzIs6kdiS58lr0Mqwl8yKxE5q3vntRR
5iGXmkPyRWVtHt0LWGx0IUW/0AsvapYpiq/29uq//38iBV9kFwjvQy7j0cYyvCHn
ZpkBdIm6/tbWf/xCrtkSBF1E5prpz0oq5LMmKCZ0Hl2OCM9DPy+3IpIFRCnWTYdg
pnpLhvT9IVf56NwjF5y890SZHyxD0zKHN1wiAsy/QdW7Rg2E29rJaQHB2WGRXxFX
oHVx2Kj7KVgELIYxemIQu6/s6IXojKN9vxSTPl6snfd5GVHQnpS2CB7H3aT8krCl
md9uuyK9ZVwBmVJT7swnTqSyCulmdakYqC/ZaOUTqrbcNTYIW1Dy71q5Ni3uELO3
u4stFGUBO6PCD+C+IXmm8gflgUaccJfIbnmzu019mqHwDA1dHxI4m4fyDDUCjgP5
9xoqDXmuJevRf6Vyxr+xPc83viWB7XVBmiQEe+Oym6amVPj8jGKwm4j/ei3YpzU+
s33KcQWCqPMCfJngOAZqWSix/WbClxQg158WqIsoU7UWznCf9DwxMPPdCrOprYWh
5nS5/YA5AyR8D2xZp8kknwGnemRA0vhg5IDsR3vq66aXoAbw0kYWvKuAfKsBGryf
G7LtF3GDFOvAlg548TaRJwiCbjU+32Y0tHYy80VFDbfE+z3Gr/bbmx6fYujFAfUg
FEMtwwHepgHEoIZyQkTKb0R3zB/GQuMd38/pCf2wRZ3jdYyRkCyIbvcwJPpmHSsl
CgjRt/GKDGP0BV8fo7mg5KE5SnQmaIhs8F0hqgm5nWnj6vRUWYN04lV5x5a+X89M
Ayhsu7pfheJD7VrWdChFgCNIbLnNO3NKypZzytAXlTxONLMZLwrJNq/2quOZxe0I
MZw4xlMdiS4uZw1oFzsPk8/Ouk0n/bgt+OQbzNKjaAMEGPJzuhLMM4mM9Np/BB3B
JT8SOhp36xLT/JZUA5WFaWWwV4iRahvhbtZrT06dEtZczPjCIUS55Jn9Ic69184u
JshBO4fTn/B9BArbotCDOnbPOV7YpAzFIel7c7SMtT5s6b6Ba669lE77dhdZgDS9
4MHUZqtgSdU2g9yhHE9VjOAjcvVfA1O7jsh27A6jRvpXd+119xBk+ArTnJ10MTpr
qrrj7spT15NOuEAnU+s60aYhFI0aJs9VQKhdRSRTqMd3KWfF5rCpW6TsLbS331/E
CtsonbMsIPBRes9LbkWc+5iAKkvnL18/1S6FW+yR1F4ywBtJkDSCd/PLcEfWN1tt
aGA4M/DUUXIsCvcHzcgh7Kuh7BZu44Yp8Q+lFRzQcAT6bzbAEtfjQ8rYajzT7bFe
hRxfmph+WlYohZlq+9Cq+GtqLGJamjkn+xYgJX6UX/KYft0CE/Dw2vhiDWRwuXTs
+JaTuoK4ZC0Z/wLEMzI/oLm59jsYrWRdPcVQ3rO6Ekuo3SMEN1IEPIVZZzTKQ6tJ
VMrkqmmFTKl3pSQJAAkPqJlGqKMgKuQtEeSjBk3BNED93nh8n095aB997sNsogE2
zlB6Nau2h6KOXr07Q6+2IZyThPfTK3q91UGStPeRiBH4UUd9Ac963tImoOd7sRUJ
nCun1AKmmXFM1tFD33zIsa7mcVPr7EeXYSiZ8jIKkBF8m8F1nQw+haEw9royD2UD
z2kjuGhF6v+tI/dNNLI3C9T7UpT5H2JUR+NXbOasB1gO3fypJnxOhQAohLANQfur
2ucWnvDIEkT8EOdg2KvGnl+mu0LalriTFODs2bht6UuSOKLMwnpYNDAu/H/7PbMU
kv7K5ZxvP0WgFQgCR+M8AHKXtBl3aL3pIvCh54NEMcio/wluk5i9U82xNdtl2wLH
Od+P4Q253gDO318yLHTaywNInj2/KEo+HhfCSIJ6Vg3W6YcGo6DguLaVrSwzHX5N
WqVTVT8GTW6S2GkNUg1O6+UvmvgWzBEaZnppEA1FuyE8EZR50S4+Dtn/dqS0wAgV
fRxIgln5CZZKxV8ejbKefyhtpNy2+zK0qlPvanQIgiWziVRcEpCuHGhIpIBiAZRZ
HnacLQjKVseyiixaWcoatxb+UTGeSZ/POQLoqoC+W12P/Q0gDoKll4SC1Z7RpLIe
UZSS3fjBBkzmyw1tZsaeuaj8o8+Cfx8NdmCvGtYNG7dGfUSbp3PweC67hCwQujn9
hBDeKWrmCwPQokwNUFTq4+Bo2i5ahZgbl6LPxpOY285XYCuRWvNQVKssZzs1Qu2f
wFV2tckoxL6ajHaZEb3Rag650jkZbgWwuXFd9go460fWTOgZemcIEbQBY24nSwQM
dzZCnvoOdG7Pup6VgU1worWJu3Gi0Ey7QOC4uw+DFC64cvBKm4ptR3WxdyYTXO4G
lonKjsF9Pqpu28VxWKtnTeS6oQfU5ttUiD7bZ373dKps1ZzQ7W2sxrRNgbyz4v5Z
x+fuYvh9z6UtX2s80uD3QCkfZCqs6Lmf6mbJ+9qchrSrRTK9AiPOk3hH1CrP6SFb
ztVv67PGkcPE4X2BLTambnw7GR2ctRp5vS7kfzi9oMXwkDMak47fcqgXuMCc42Tl
4PAh+gUTl4yjgHb4q4DGDvtza9+cgmEoADp5S47j3iKLFTdqhKpAZInICJF1x1ER
uUP0XRQpAHf+8ypBgboF9WbF1cyl8DE67DUsIpO05MQ0aG26mBQtCV2Htm4MG65S
HVYqPBWa5Bchi14b8ibju1PnMnAUTtq4oweLnNpWQ7rSdTM7Xt77Nb5B+Cx4CmZo
cgd7LXVVLKSqKtZCL9kOOYdl8LKHiyWZ8/Guo4pZ6OtFPM6qq1onMHfI2i6Wuj9Y
91/HltpHHNMpqinZ0iyfJ9BmJ5wctOYESlbn/RzNQs9ad1m6iJuLgYfr573D/M78
D80431ABrcxhieLw3JRslL0hmaKLb2GFUjtxMFdFNMSHgeDnbjcAHOcR1kO8/h0i
kPqFnDj2l1pu+Rw80Wgct4k45p5i5BcL1JnZEFnqjtnTgu91goeN0Hh1fI7zkg7B
UxHpMViUunouRtrVbu/P91sbyBP9O+npuGkSoqNh1kTrDIGTIXEWiVUseRqq0vjZ
tbz1N4NMYpbpYzol9dAYcJlrePhcyv4gez++IYcIxErwA7sqCtHCP4x/UmwrpzBq
2slZveVEOha0qCSn8XxcwQ97sngzHf3FG+CRapbAAEKi3KlOmJFft+d9mxYyJD+G
+PJPQBV/9BqozNa273dbU/UWMn69a3G2VXKl2zxyVPK0kKkjT5Ti1ZM5lgSyauDg
d9PS7IY+OTGpf1IVg/WfEJgSwfZekJBH2bK3D+4EABTsKvGCarIygCGy/aFqJpxH
VFTILX6AjeFlXinxBi5lfZvcmLBZLRXzYUm2Y6/ddZeZtWBu/Fas5B+lvlu43ezS
bwceVjpqNF7CeW95c68KuhW3z5nHeHHae++DoU0JsTOMkQ4/yQrB0b0NgCPONAWZ
zNVUMhrPPbdPIOpzT7TuJ4KdWCLS5KlljhzVDuv1CV5XNWyRhDyhk4cFuvWyX+gg
yDZ58OcxzilPxkiCx/QxGTgMWvH0GlBgWwoN1nfZCh+9Wc/vOPmWuFvn5xM2h3aq
V184KNHNVkCndFvJQN5PyVqo1zh2h0H2cDNFo6NaynCSWnwicnqzkecAhf8j+5tJ
CxswpZ6WShGwSjSLjMAmPP2hfneTODyxZZLBbTvf8oLlATEwdnhcGHyuVtAovHeq
slEKtaWgXb/Pgwid2t9UMXedyAh6PsbGySENZ6YUYzlysrcrBUJmXfkXcQwB2Xz+
+EhPrjrsfw3HURaCLZKTzi3jT798HQggNeB2+1Ww1/zZabRpJ6WNkcTOgmFXeiG+
79VNPGMUtQU//oqzeGEvCuoqWZryihoALsUyL3BzJ5yep8A73CD79yiFJ7Nz96Ub
SoFXj+aFxWXBhIQW8al6v8P2gi/bNs9cSzATVTcibVjNjX3uUL7JOm6FJpLQbp0K
mNckiB+r9AAnYWn7FogD0uQ5wbRhhvGMH+BZZwjK5ivW6yGgN06YFHcB+68GE8fy
qLdP6edubH/cOR1PLGOPFzBZ9a4UzylWrqXl/l2H5kV+U5CVm2CHSGrjx4Dk9Bzy
G1o0PxPJMVMRZp6uVDpUvJBPlQu7mb6Pa/2Uu6gSMAhB/dtqS8YQ2oCt/Y8XrK9J
vwunx/o+Br37NatWc3lrSlo2oiRJxQBpXmrxQbdyjMhEhwiKWRcpWCP03b3eBLwu
QkCFDeWF4D6dEF7IfEGCfUJXG/zNb2QdTN8xfy1FNrcU8TWZ605THoYJzxnag6cu
KSv1SVZ9Xd4kLcThg6Kq8oSOo9eFofo2IHLvTd4tzh210wGkN4WlnXGzERiZsDPT
3Rgbm5f0MZyW6wUAmgO0gIhCjVupQHbk/7GZRK9QtwdHQlpB/lxPJ7zudSnng7+N
2G6csd3WbhJZqQgo48jArSYLYXiEX0ZmMDuqslQSNRl0xgYzcYjijKfCW9qux1sN
dIq2ZknxYptQ3nWNO+HgIB5I8t6/oH5IMk8t2il7Zjh5srfqVtfrDYALEdlfQdIm
1med3aznKylzIrWpv6SDLs2Bjpd5pVD9SRypAw9eeb8Vn15OWQtB5HCqUXFj6EVy
gRS1Xy6yHAc+7v6pcEoafnShkfTr4fa1dhR0GtFbMiVzsuyUy6/TAJ548lA+5jiA
qRqaYdMdBO8ikH+7OjWTLLzP59J1cJPD6Po4ia6NLuTzUsMuw0T8DCWLzCFlyEV+
d/uZlVjRBR1j6jGh2Hqiw2d1jnSmMqsg/LjYsT79osbEIGVVokzlNJwXEuIJzlOV
IjvOl99l4bcTM5vhT0ubJfQHtPd56JMZnEEJaTlB5e4mzTYPZDxSQdObVteweu/K
mDxPncoLX0dn6uwLjV2X2oLQXjkF1ZX1Fv8cyHSHpipJdYsWaA4tu3PdAhWD3hnz
e0bSEkOe/y+QZCAa311TNxLkffv/h3qZfkHIeccMZWXVpjEG4CtXWjiF4BcBmAq9
fdz4KK7rjT8F/dJZpCVYI93n6pKa5Y8Hkw7AYazbpJLhpIDoCTHVVpx5qfMFG1cW
oNMd3YbF7XG5fs+xdqSvyaj4uPUxMvD/pdrAhgDhgSSLJtUp3ACvbS77r9grYbG3
0WMwol+loZvN9ik52OiYFAPK6Dwlugjr09X5eyutrKaD9N1HZVKmYrbFCgaw3VtD
gK5vMfXkxPZTkF8opxkllCfMmZwFrZAshsI1DUyyhlExO3tpmKrp6IXaN98I/L81
8lsLbKfBloUtZTyjr6eZdQgpciQWNFTKn+tcnorKoOkZk8c8ZFMXxOPOLvrxW0j0
hmrOGgxpYef1BdewKDlH/4qXkzYODhLUCrMUcU0/uaK6ZctK5uF1yPdol0aQtZng
9VNH++ZKFU3+9p+wFAEwL7Qt5fIeR2G6XKBcsGn5Y2Xc6sFYsTLQphwaF6Z1HgE2
mUJcIfEJq8sY3YV6FqCwS9VBycppXm2q5NAKunxV9FXM2D282yyHddTiecE/aDKa
T2wzrl9dHwOWiqlLabbccAOWT/Yw7IG3+AYnqli53qljAqufcHTHc2pJdUhs5RL3
KBBFhTYN0n1qbERNAWWXSB/7rGqttjVdQ+TETrrE58lP8JXwkG+4M2qwZ6NbZAZS
5+K+KpohdbB9970epUa4NcbKlGY7PeAGOvhhqu5T7pzHrk544Rz3E/dX0eo5ftWC
3lc4+0zO/a38fdCsEl1YXenHr9azjF37wZ7z3+qoLAfeuqxt+WnajVlYYX5viUQE
s0o0ECfPAy81q0g4uDzyMjGpy5wPRxijMs3ASOlEBlJEZBRmqxfok0eR6bgr54l4
spUmo/Qpp15ayIj9XbZr82tFW89DX15uDJD0MdlwJCwfq7FdGwlFAOKsXVB9/4Bz
w2BMlAAdNEm1Kkrz03wh/9IXY+KuYHd3TXpdKfYwk4B73+qh8K54NVfgz9YFKvLt
m6NfqFbGNxjmRLl6TbOD5xzQdFMXV3+G8jPfo7SKvxkuwivYn0uleWoi0U2g11mG
VR26W7tSrEeGSdCY2QuytXXfD9sXPVOkn1HnScIRnDCZXK7YFKmf6JnxPqbEKx45
slQ7yJICk7hoEjxq+PJc7WcYBozcydtWOfaPqAZxn9upDYahhPgxqcReO2VlRiXu
9HI/yl/SOQnwucLcSVz1iPXQvtB+uno5Z6j/+vRoBJsuMrDTs8EP9xoZJzWMX0NO
UWxi0XfAkzId3LOnKlLiQxgU2oXiLCd4ZqDGDhVx8eJgvxKWGUxXFlU+SgRoBccM
X04RniOdt4z78B405yVaf+sW4tGcIxsq/H9vdO1uEQuaCUCOZ6U57lAAuYm0jlkd
OiPz7phekmgjuuyRN7rcOHpN5W4GPPIW/aucGYVUzBdBPf6yX/QRShy9/ge1zfMa
gaPirW5UKgDGsf/6ke0m2+xcn+jayyFUcXZfs3fH2ItxbmpIVLfD1BhYZ8GLslN5
XFOFrxSXM5x/0TD0Frz0hMJTu8FjMxhsAeI3pai2benO4ZCEELzYaw7KpXRxdG0d
z5XEBhjCoyCF2lsKH09PgbPjvksa3jcxVyNoR+R2WILDZijtF6xk9hyjc1TsQyRI
UqVFNYNs36jDvFjtWQVxMlfwS8Nw24VfuWOoMVU5QbqFrzpKhSU4W0V2U2k6t/Zg
jLJW4dn3cLWiHgmnciPhpo64dvEkheBk/5Item7ZkdvfjU5+MOlIc/wO8026VZAC
W+XFjdfrJBHSCWCFMiZ76pLIou0CxaP84sn9fbMoEzo3mlzeddD7j/4fn6TswM8y
8ED8KqOAm9t6HXBx7XFy6Afe7hCgJl3R3zZFCrurraAGEIdkZgSn48msbwuEnKRd
PR8Yf4i+RO9390LuScHpxxdc2eCC9OXOqoW6RGQG76+DSval0VUnhSPAyf3fyQw9
3D2xYRSq1q2v+HHQ44Ela7GqETXmS+M0DR0En21wfcDjVI09nu+wAvjeQVhuOptr
S5LW28uNVYBJcCTcfyLY4akmLkNOu1SMg6UqRvCIgoshcN7KPymmwICHjAEQMLxV
SH/kh8K/1FjOVWBkT13B6aXq6aL1Txu/IK7AwnqfpgpFaYnH5XaN4OOaqfb+gzjR
Ci5k9oh8Nr+pPnXU8175SV8nVORVFzHszNCMP4fb3Z9bvFC2qMrwDFYkV2DQ09Zh
I59K7CJa9gbYffwDotmwVsRPUtr/vP8WJadKPFNXx1Dxp8Pf2+kxTpLLeZJ459j/
yxYtSaTNtNKCKhgAOMaIcyb6jFI8g2P4uW8u/ng9bPo1HHfSq+Gjrj+Kvope5cbN
ukb8Gh9WB1VpMK1gr/uUJlk6dysdnje0hv/yndz6ZfZSJHjjaFKJ4J2FI7ovzzpU
NWKgKJBMVQoybBH3jsDZVuvri7a1y8zFR6wsbWjGYMXjJ+tEjfKpfuGhQtP/s+Wt
Z3WlSWWhaBSYyfUZYFnM9Su7teKZ7j02+VfIamFadvh4eDDe3pO090Lgsy/6u3PR
N+WncoJ3Hv2YNiTpW14MbYjIFYGRP1bKFr9JlNn0EYYM40BgjPMrqdulMiSLk3ib
00AJWhN5n+3VLGd2Dd2dULtJhFtgCHXgsSbtRPdKIlImEmrbY7gxw7qmI4OA15S6
urLCT8+WK9LNGe3Wf0d5n7pD9c/8c/qZ28uyj5QG4oPnqV5q7uH7Vf89TOXj0NC/
Az7MWL9ZblmE4oKgVYb8Ai+pJtTUAwxR7YB+nTQ+OmqPFVTNsoSqUseDEyh7oJVi
NBhyk2YC6L898/mUv5iElHU6t2C2OTzQiREl1ApLunIwGQW8eJ4E1mT+lXrGIQ5l
URlDPVPWNaEK0pOKx+GTvyLhWTx2UlVUQ+p67Hpij8SIpqhR9KbbGW8zJ6SpTmZU
v8KxTD1YexVPyTGtHDe41hUXF2SOm5CTV1s8O3TzbgG8xJpoPrgOuZIfvr/n3owj
iDMgsFXzHu+N7gS3UmzuUls3sbtTNCyAzNQ31nDe01hIrNY1LjxGEx1P+poA9G1I
KNZT0qH5AK2V3mntg8gLctwj9DCYnJNubLiYv1+aNocn5lxkEryto/0g7/+jB7Lj
JE6Mx+q7yOMUtq0PPZL6mBeKA7Jg8RwA6lws8Tod7LN9MSNCDNL/HjGQdJvEQMV0
sTZSI4CtoWziewFemCJAhNbZnbDH6WuqCEv3d7FVPeG5g0UD+Lrd2KTsnKzumcq8
nhAqvJtM/cmFwCeTl3Ne1McSL1rnXyoA23OKNjjFMJOHp2UNqjOrDpV7FQPw9i44
roYHIF5SIUVXqnWottpb5R7lhqY9T5vC8f24QSfAm8T7/P56Dhra5PluWyeHJ0C7
QHSuTTraUVrZyTKpFrFcFx1nS54VVLtceCA2aCvTxX0Dt0YF+sLpbTmr3wZmwxzH
`protect END_PROTECTED
