`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O0Zbmm1zIRYWSVXg5uMlXAiAJ9bBZ5OrK++7behZoYuP93shT5djKYpZUpmoBp5Z
lSTCZN+8OB0zdvaS9EkHUQJpgO1V1hYjFqtViCguDXxZ0933ggM9f3cSpt768gG4
vyA2la3oVAP28t8V+f9WBHp0QukN6rJZRGhO4V3qJ8atuXCqxoSsx0BP/r5cercL
Bkg1WYBtM3RopRdffOdtEuB0GeWBwBJKmFa0pUBylA4wPaI2XfECz0kPsp49d/bt
pQAL+KAgSVpIrndFsaK2o/beau2SsnD+G8aBPO1sw0q9PqcLLQJcEWQpHB0wTEhr
b1qfxYrJ2lvUIcLNAKr/Irzgh650DjW1iVl/EhC56D/SQoMqz3qkUKthayv0FKgo
la33HftqJbqhiZtxS9AxCnFEIUQSV/b28VUZ4L0fp0JLbCqEnDuaA/UmBl7bGPVR
TMjorGwEB7ayF3saJbGrZTbFDtlzPOEkWgtu0HBLtqOhr+c6UAQkediSvxgHkkBi
XtQcjWG9COKxnLVc3Il5QhXrvBD3ZF85nH+UYOkRAXbZJx4O1PWY6TqOwl6+ixwP
hg2ty+srx/eJ5CVIb0btkqKx9Rv+EGw3P0uvQhA65FDNTb5A8K3rF+H47eUdP5Hq
t5WOQmyBBaYlgrtSg7LTRKW8nrPXJW9BJorTkak7F5Sw00OLNvgc0LtcGERRHAUX
L1YmUpOEcRFVyH42CDZlrBKsmazeEXDncsRP+vt/3L4CJ1zLU/hmyO29kSJWAhmq
uvtEKY7m8CwjNo2wB86ybns9ulTYnmUHrPXOSw/iF+6mr9pdy4fzD+3dls+TYWay
3WdUtUH9mB0RankHhWAmMxMhF+ANPZjh74SkUFJi8Zat+Urhud3/A1jlKhGdaNMW
gfvqZHZlPKu0bXSfz7nHTOtyS0yI1kxVvdtWzqjW9c1tB7arvghFzukakbuYjvs6
tm1GN0BP5pCc1x1XDxbvOgdApe0D433tW1Hej3DGjRLTvfnIVuafd9F/NCDXj1if
LjbRlcR9ZAW+k7QTD+oUxYIYxekA9FxwztxU6LVLHFy5oYybWIuHpL0XFTRFAumS
bcrlgfvmnAvhMwanrrHDj+Oi4EnM0vXXHC9p9I7Z8MkfQdyOJrps96jpVW5HNgGL
vIIBMSSVJJxwITLeweL6+ni4U0r22jPnCV/vRQ7R8qaoJZeuJsKjS9xcgG7jTCkY
8LV3mMJIChPugg3oOxf2L1pgDtv2QLE2HRSPpJSshNMRNofAryL3qHjdyBWGCajX
1XzoprJSZOLBq7+5WSeUYBZNd4lGteEmrcWL/grJ6yA=
`protect END_PROTECTED
