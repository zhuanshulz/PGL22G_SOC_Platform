`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J+MIlnuDjod/OFcYBomYhqlHtAdZKCAZaVNZsDsrRYJm7UpV06xxvqDKva0LBCTm
raZz7qCr/gDh+Zg0d16GmmKdlnjQ7juVciMJM+Vuf9u2nv4qELkVUZeqps5nktr9
AGGocoLnJg2dA7WsEF44f6Vz9YaCQPZQCTMSx708iRp8fP2xebgfeu1keQDR0RmH
LMNkMFqAMasqo9SS/K/lMtyU1fTqbamHBIj6V1EkFH119i30rKuVZmDENUC5HyQN
G1agtntdD1W/FD3ns+jaW7pj5cXs3GtxfDXCwAinPdY2RQpysKXnWumJo4OiyeV8
y2xuVyq/puyZi3uOb0oBLBvx5s+46UHeRVvY4aGZpW+qR0w2sD9cksAgKO9z7JI6
rF1/KHQxvQNS1RYna6ya8PRo0+YmTVKXjhrx1fNsILfdQ7LmoC+Xrp1OOl598JIe
tiK1zdpRpN+HlNNkl50e+CfeTMXfi6txk7n5QJKbWeVRQIr/FC86AvaljBPl83dp
hg9k4xXaD5oe99OUC7Z1gCIGqUViX7G+B5yGuOwbkEenk+BxM2ccHN7PQn5GYq07
7c0ioSnFLIudYb+rZiWM6qeiNJPVHCOxs4niMUIBvZe1zq8p3JRlkERsbXv7s7Sh
ea3q6fWOpzp825ZHk/iMSjvlzkEBCy1vISU/QeiVJc481ps+d4eqonz44eCbEPQr
OdTAJeRMzhsbbyRPHPice5m500n0n37RucUS+kNpdrvUmyXkGK9hOlZvb7iEOOUa
h2IlVbKROMnk7P9h3ZpN4mPgUP+wy+Ysoo+LkcoCHVNhPWF949fHZ6Y3uoTN1Tac
L7rrJEYfl17p8ryEY/VO5uhorG67qgSxPAvNOoKoOiJp1rU6QcK/Y2Fj2STIJeil
gOyej4gPlQdP5D1w1SxcR6H3r+xx84KJ5tP+67xuA9Yox8yJI5eVwS3DR8QIS/Fl
jYLkYHYWpd2oHXC+B6nS1DWdsnNnlOaRxAo7KQHzk6OdR3i2Dhe3SFacq9pz9Niz
mfgKtK0xe0TfAkoYxssyqTEbcyQmEneCx3fdg4N0EU7ffXjr4Xi77MhfPoaynmxC
woAXFRuS84JVvyC+46rx0tdoH32SFBndc2MTQii+TEZLdQyAuwHsGpGx0qchAQxU
Qid/8XhSY0hxZvXsSWDow5Rclykd1qbPQBkK6CJy38S5NhT5QO1dSL08nwKJbvHO
RygBjHe5lO3LyO93/4LCF+beuitoX6O3w4Al0cRSicWCgfAgaP7rsIyRTejGgdJi
FiVZKJj0XHd1NIZBWbTjucDvvW5B7aJF3jX2LHSgeajzfZEdsXVrNNOhEtfr2f8i
KyajprRMrVbULhBFvDE1fpLtIirv0NSFYthUksDneQZ4BtuGrCv1UYuAqJd/hJzK
MWiK8+nOUiCxUmEEDWhN1uEv0+jx8FemE/LtdrooBQCiSHxJii3Qk/54uhx1ZKs/
vsj/kM8U97pwPGpIPrsAvB5OyfdnWjJbvJPpQociWPJUzUA9WV+vtsleHsF6LLgu
hH7k2IFBF6j3bxyccVyqBWcObCHRkWg2MIKugmHrydRH+r9R9DlC/mz1kiAs25BQ
Rq+ameTSD9SPloE6r+lvi96YbPE3UU+3c2tGt/F9xhC4vK7zYm4yA/rVJl3/8gQs
b9nDi2joMXvDw5pnsx3+7hzQ0XV5SAQLyhPo3WBi9cE=
`protect END_PROTECTED
