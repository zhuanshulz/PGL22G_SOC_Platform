`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PFHlwMVVk83JtlsBib/hzzM0z84K4VdVBfKbf6E7YVtFmAqz3r0vFdtQdUFHoUyi
uSmnM8qyyvqrJtiQgy1lH4HO8p3GVrBEtcYk/mHoUyeXdf3W/6D4/Tp8r/7xIzvO
DL6WqXxAvT8tTL8ktc2uxOz4zLE1NZNanJcjFDqYsVj2+URjLQ4bNPKF5N/ePCin
EIH/QmCZHC4AJwJ0l0u9vYBOnBKkAGOxTjX6JbVv+3wyLnNWlIc+9RVZcq0rtE/S
sTneJLdwcMos9rfWVScY67v5r0CH3ucHMa23q5OfaMVLANEn+bH6t52S7KlnVt1h
m+5WK8Z/vF/L8V6W60SX9fTKR9oMkOdcZ/hM4D6SvgHBAfFXkwy9G8InIbG4jnIH
CXLccGKVd7nP9kvfl2N0G8E6JtbfMBc7tA65iEkc+Lj8TFm9qQP6I/G546EDCesG
qctIkcb4ZRmEuT6pCe4rQQU8fsP7qTejjRwPIjc44daxlqf66rjqXRP0fRJKIYT+
nwcFgf5LH93bzZs6m6r2yaHnnYdcNq4J9X1viqjbrg8I1vHkU2J7tSbyrASqLoBx
amuP8QEP0an/Ex5Ko/YMCzLeVYGa6d+RC0m7uCtTu01ZxKoKqUcm/beNjNBpmyV5
WYWF2onSO4LkEF+wgYLus3GyXO82x8mrodHRc2QZ6PIHGHWdreAbC5uVwwQxoF+9
dhq1Nj6ve55gotoBfm70j9NbEwqxJNpVkTp1IpYdUp/tC+GNzyYjqqX7tpnOIH0w
c1RM9l5lLLZ8COWoWQkp9Wtn5MJyvOPEWRYnK3XvC2z3wjcpbNFRefqwGzl5lHUY
5FoseKS2fDkrZ3QL4HUG/EUjC5NJRWaIEpQMA93VQq8o5Ts3OW2aFoW7g2PuHTq4
CFrSrcC8Lmilx2MwqTZ4k6/1LJgi4toYN9rexZna4hZgCGP88Lo52ZdF1q2fCiZv
zouR71M/ap580H+1voHSoWdIhhp/Y0n5R/X7iVk+C7b9k32OMF99tRwovbse1gch
GKDwZ/wMdseTaS+tUaBHKdsKSNiocAkNAYJSMhPROtW3kJ8l8Iy9MBqHgyEyMMCX
9isenWllkDTbIBqSc8pa7yT5ho51QDqHOw4MLEI156UKBHGkYNeiApFU+s0iK+Fo
EhmmeZ6Bbp0h9K4NCfUcdQpRC/ME090PSYqiWJF8JDQaAwkFK+ThNO2WpxYwhSg1
eUooqKNFoKvSMM0BLk7BHiFdDvOn2vSqrVMJ9Ih/XyKUkNVkGE9rfO+Vn0nVK+cW
DISatjsBY1LYy5ROsr3bZeDPTsXkyERXzx9vvMm6Tw267JkqIlqHNTTobaljXZSf
CcpsObvobQvTMvMgSUBR5c87qIX+zrruSlQCM9j4ID9efsFKJFMa8v8o8t1viJG2
sAKVuyQzFZcTutylgkWuBy8YMaI26ljEqif/d9apgftEZ0+V6CMExU39w6kSW121
ER6R8NOHT2VCTG9UlirbuJXoKwiru150FzyKoyRPDMAeoNTpZA7Nv0zraRPYKLsL
SFzN+wRAdFXqhhx5TmThBqlVDqxemYqK/zc/giuu1iQ7K4fLss+PhV+nJCFuFjL1
S8+CQfhUt+tBeVM6cz5xqCX2cX4rA+jePDFbg86J3CGJYAMpZSeRHiM2DpOwMVUo
aIYpYS5/5aIpi4F1vxXVQUElsFfRBQrJoKvRmQogSeisiBYmNoafG7PmFA5bgUsN
eQ17pEXA1UqAfl9KbSlnLRAm5UiAUdqqb8F2p3NNGsFnIK8jhCLQRHFXbwNF2vO7
oMMW/K5WeD9zCi4KBshDNeiV5i9bBqBr60fb3SFl/71pR0PftVzN83jwfdWoblvl
U/mGEK8zFr3ImQhGECYQ3uCvJr6K6cyLpEqPLT4VExG9KIy+hJgUwXO8IIU02No+
bseNPBjk+l7bGy0En3CaDuSa7MUTY0rWShKeXG9SfKPyj+Yx0usC7Wp+x0wqLeap
AtjR3A11JlKQGss1TVC/J3vOWqrj9/G8jIEwfT54y/4BwT+oSrWunn3+1KyC0s1l
WFIWGS7wGWaTSZTBuSfiDqote4LnKY+nln9ICcwBpisJfMA36rOqF5qOHlrYOKrb
6LVrBeiRbg55S2zfE+mEgB15FNIlSJQedEybK1MjFXArad2yBz+8QF6zLwAmjaNO
DOF2bOkU0ywfTt74KumwqBeYcm8nNpN7XbmE0sMTlzlNDLZBy583E+LU5IpnEpDi
nJ2JBH0knFzGX1sQNhh497sGwN1/ZtQsFJS6uLJ4oWvaGVNY9M8Ymymllp+xhHRL
GHrmd+a0wytrmcSQGD55SNbxqW7o3SMt56gkWCWXO9NVCt4sEiu9MvSaUITcHgM/
u22sdC6uo9ZfMSiWM2cIgGv74euLyFuLKP9e1i5EOOXNC7ACuj0sLTbi3QxeoZhn
skdWBW2XeM0F60CjQb8dQCqDzwzhz6RoNNuenySg+NrfpHM+/WWciPMu901FbmbY
JU327vhzq8YojOAEPjr09j8tYQ6WtBilaVLyZ4m2NSgERdo0acyeFYhqc1RR4ft5
biLzjdlGWqGlPk5kBitm5DwT33jlIIPWD8waBrWBWxY3CNbEQ4282DLnn6ZTsWPt
4dvJXezOSuLLR5M/BbH8W0cZJUwyj0hYJ1J5Lc05zz+BnCn/ANZkqfOj/o1xzZRo
2dspAu17XIXEFSPHjdPBlZkIIQw3UYraJTFnM3mCjVVSYvwvV08rveTmeVyWaql9
s3VHLH9suus+JSjWHgC/dYTzBO2MeJZR1n480jSgOpoUBbncwbwahjL2Zz+v0gaf
rd4+k8TfKpnBuZGRBhfGIPLJi+icOk4gtwLpR5NCNWA9plzJX0+jBQjVs9DJfjqJ
TDn8usnYneeaRAeJO4ZoVVNk0c7/nApJshQhnnifIXeXueIV/5tREf3j7ffNlJaL
E7OXyEPMUnnGy1PkR7m1ugTzSoP/RAEmk48anQZkYKxJFt79qVqsDyYjccPeeB0u
mcdurqc34wsyLFA+anfX6PgidgFwXbqBllTI+K5lHmYekDxnMTZPgeAdVLvWANGP
0DoIhKGakE7U5o0NzE1dpnIj7m9/jqfxK2ku451JQ0Jwf3Bzx+8Ti79/j9MI9KQ8
LlepsWBbp1meB4gkbTWdfOFHH873MaI4CpJF3x9kmHcDhab5zMUm6owRsHn1WZgQ
`protect END_PROTECTED
