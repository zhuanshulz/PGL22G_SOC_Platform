`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QUJlXyrtQX0ooet0loaXg+CMHw/LMvJ4lRkOcZNlCQeZHb4NeYNAKiaffRqq6RvV
/IMGB47iI6DQoKgK4inKV1IkJ271IupXVSgAVBZRl9xOMwndsRYjKsvoLvbZmfpq
bErVGkm4kee867t2+8eUZNmwYKjRVGtnC7s+Aa08LuFRn7dLNPRd8QNiuFs9aIXj
8WptK6n0bhbeM1d66BxUaF8mNXM7Qi/YkcgmDS/vRdObqTFxSt1wz3FP5N741leM
pBJEA1vey+5JjKg0S4acDrTgm8Hi9ciQiZv1fYolLaLhJwE7+ZlQcxEVTqWXB9tf
KD5tASb8+oi0N6z6aNI4bXpTuwfCcLKe7nUyLEtJ3wFn9izYsmnjwnTgmr4GvHvl
fJMReEgcrcvYbMYtTwnmvdY41c17HfZ1bcZzaz0uONAz6YVT8nmjwTnQ5RRYU30F
DKJf/bBnv04wCeMjoICN4aN02QVsW23UcC5UHoedUn4IJFV5KrtKpKJd1S6vQ4F9
BtFtThSN/xt+fPsRneyyd9AGX7P5qUL4ND7C/KONfNfDbcbzR7OCDz4r49uxQagR
0kcN8Ajn3ROPt8qDv2d/DXVN9aLjTQfibF88prZ5PYKjju2yP+5X5KEc/TSg4MN/
tZQ1WWuYNYK853lLz+DHt+imZRNBJbN6xGw5V4C9u+V+1vF/cYNbBKFj4o9G/mAz
aRKbHqmWj7WU2y4JVbSYjZiJpZCwZQghmFnYyVbiM7zBu0/Fd11VGVJE6xvRofeN
1/9yDGdB8XXWuLGPAB8BuA==
`protect END_PROTECTED
