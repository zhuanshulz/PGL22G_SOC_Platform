`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jdnzx9KApUspgQOnCLaK4DW/Lydy1E/rA5hjl2rROhl8LtiVzSssupBQR7gtpKdQ
M2fwuCPQCiJv9f9GY9T8PSJb8tKBkTXH1bZ0BdSEfg3WUPsqS6xcxZ+ZjuaDiy7c
SXn97teCHfQKl9jhm5YNrv4Xzh0XlTzUK1opTDYuyZOgfSNT9B13NUV6mO1ccUmJ
K+JDLdpVrqn2bhEXI+zM7vAqUerqxPQvWp5DPj2X2sHxLN+kVcRw4ZnIFYU2sbga
v8KNaIe/dAs8cF6+Dt9DfCBzkcQWyuMpru/LwZR853g0jf1KX1D/azK0aR3EeQyd
Tjw/8XCTcdyk9hhXEMAu2tSoVZ6QeNZIbwT/8RtfVQb42loQnG4sqOc85uN3p4d9
3p5ykPZaX9AC/ViF7ouVm0BkDIqF3AXIU3qmNC4+aWpM4syrlltdAqSSqx8CY0xx
CTgnnLqGaPP3L5IqNU+0XsXDuajftM3vGrQQwmXUKLLCbZkZ18GhgWHjb2SQGleR
9poJPew8M7U9q73FWlqhKzFBB7bQ5XgemexB42T8PNmabF5jv5pZevqBFtba+jV+
MhEhPt0RTWHlAU0q26NDf262s8+uTJe7lx4HzelZR275RYODVjBNCuBjQcurwjq8
zKUQi/RfrYzvtNXu4CU4lstISww6VSEVJREChtjQhcynmabuBQM4l+XOP/DMoz53
cLVWhVlG7S4pjcTFaKTetcRKQEZIRgalqFWR/l/xtJS7xp8YBdl3rontKknm6bSU
sEp+Lva6uuL/ZxyPNGEMBOhDLUndy/q8xCgYDf74rdA=
`protect END_PROTECTED
