`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sUlCEK3IJjT1FH6I2Z/AbwXHKS9DZNWIIfAzi24pzR3yfaDfRmLxn5Bfn1rMfcsV
V31cLRo884fmOzgUZgBVParhy2b8HWY1wXoXVmeg/5LN0mxhzqJJicwfrA1AOd7s
08zopLZZGByUp86Zn2kJLrEJIt+/E5ID+7oVdN0mwwcYQuV6J+EcWtpASXhY8fcA
fuhjmpFx59/aWDiJiFxU1TBNYehPyu6vDPwYvykVwbRjvt7Zg4JbA9qH43s2vR0T
kJVBzjBltRd+fGPgk6URy9RFVJ9UB1anPl01d+JuvlT2T2Pov3CQBzCa6+U5W+Lx
ElUTnk0qyOK1nzkpI4gS4P5TwS3rEu0dMoeLSbo5+QG6/C0w2ynOeVnuAJu95IJz
jPGv2Rq5EWKD7F82ZEg058Hx4Z/L/G20lTzbWad3GTRQoVwm5F1xJsI5gCEQnNiv
Z6KMm+mKPt6brIcYlXDPH59EKTJMCikYjJezio8AFNSXl36aEhzTXutrH4RiNjHS
ysaGtGtr2VMKuUEQ7asV9IE9AXDaemKgRu7+8gVh5dDls4D5OPZ+iExwYKZvyabz
KuUdqOfC98y/eVvB7zNZGLtQuUrR4SXuWzwMRs5L7KTBQtv090LBgm1LGElQCaxL
ePO1LzMHj3Js4pyYL1IPR1BH3A8JIi8CoPzX6UYj0eVhkhGUaeFAa+1/VI5lYO5c
qNHlDgIZPJi8rgXWsi22m5xAj69a9I2vE7O9eyKH5ORs2GIPFNnpW77gIhszIPjo
kSJnI03r7erOIrY9xS8tGMHM1pxqLNI35O6QW1fjnhHgX0o+cCdFQ0DcYSnB9o8D
ZgjN0tEeeAb9TFzJwJ3VydCcmQzvk5IqByZVAMt7QX/LK378fj2Y36RHWnLcQA9E
xaMdzb8x8bFJ0WRx441B751MXI7etVkQGR3IrVCchtu1NA+6tQ2nWHbegVUClrCT
YxI0GjNFb5EbM0fCf9HLHHE4zu4U9ctk/c92WAwPqlOmyPK3ARLxD9sYrDAiBFcR
v+MznaAlfLyMhAUY5AFMONlKS+mc3FOmIBWVgIOVg2Ssce69aVkJIYJIgvopmPst
MKmydi9+eHwSmvrA2+b1Z8s+sRCrcyYNNFxFkU5Op13Q15VXejgv6GccTiIS0hJv
`protect END_PROTECTED
