`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O22XICdo85HrgSknLejPmV6isN7wkyyvZiuq/vqY+19pt7HEzcsfDLdbFUcsqCTm
M9EqJViBU5458I0lzlz5rE6Xg2ar12BJRLQLprWpXQxhp0U9AYa06s+LtMOrNDTB
RISO8/J4ptz9AEsfvw4iVzronmKOit/fxx+0J+3r0sEniQp+v8J5OaCyJYcslukC
FgCmihagErL1zG7MaW10EnwYRbB46UZJft/5uHslFUHnJermLoie1aWkHk/jGJ3g
2xPU2NJ+ChuONf/TubZCoMZboi0C7VYwKvdZ+dBetINaOynuDgJBe1jdCYRb4Wbn
AOGLXRPMiztJ2d1mjJuoYXVC4c60Q7Hj/7HWRjFuu48cUfTwARDxKG2+NRgkMEO3
NJDhdgN7hDgm2njBaDZGL+nUAeqdnOqB/dpp9tuJwcg+x7oUiQKAfdeaG3ClMDA7
CrYmaAVNFkpz1ZZwMPsCxbfAAbHSIauyrklgXvOeNKfKW2y2sMVOCsevaXZa+r+r
lDgafRZb4BqVVYCAvTh6j/fLa6tYyRuA/7ZpYiU6FBQOJC5lBMMB8XdlgAwtFFOd
uNF6dWDuKVC7GxdYPfp7ATFBshjCEQ4IgrZF7xhDfbz6Kkes60B5NHySJ315pHzw
sU13TqIJHbm73Nx2mNo/aMfifeqNjTqbY5xxKHte5FYWCrI+4j+wjoctkAWwcEau
u50c+oi61NFx4IxGH/AYBgb9ckb0rBtRoAo/yiiKmFGd9qwzC+haiUk/rD2/mcBG
XOMdqOIJGqI0NFJWQ+1hniRJnsPXBuluh4R2AK8fmHT4FPixW5d3hK1PhD1GWKxq
R0VTEFIy1SFdEZyYepGbNw26ERChZxTEw9sL/yn1+Ee4IQNyLiZexzh6X38cQY+1
Y+1o4C8/u5/wkGcxL2bbWsUkD9wqgbdi4OmHyQwkC6xg2NlugGdLxMIc8JpwndLe
QHxekWQVq2ipVdaOXyYOiDS5CMpxMZvdwyMWCrc6GepKdvOUP+NZhetEXjAKX+6X
i4Oip3gnEfcUSsldg4rKs3SS7Mj0ln6pvAp6CreroZ8n1av4pUdwGyAjAPjnnKsF
HRqjZ04IDcFHghVWAFirtTgxjQ1HR5mpMu0ozrdnugcNLx+UuouDdRGFcUCJ1Ogp
Cnr2bbWLcnysVtq7URwkdHy9fuHh3g+YAAt6TcCoHyIsN/nwbeYWvbFhgCJV35Ri
vRFwUO2yZJc5sjIR3EYZbXRO80Z89eMaJIfZKWe7p3Fvacn96fw+vtBxmyJSgEC6
Mw4xN3EjOhr1vhP930PzuQT+ARsG3juyfgH5TT7HjKcjDMd49kgpyYMkUZ0VAjoK
s8NaocvwRdOlbu3U1h5HQgcPBHmWiv/z4W99pp6qakQybcsGW0elI/4fSchfQlep
8u6HKu/kBeuBPyXEapdUa8Iw+7UYAre3VgM/bswX9jICJC9jyhuldPezvay6Cjxj
tXGH1tWdmEKjVXTyTRr0EA3cf+0oq/1INc0tAKecQNxzGrYlZSxsKj7Li61z6IpN
HJ3miD3tqLPmoB2/R3pWFlh/9DtAkcs6VjrOlhec8rw=
`protect END_PROTECTED
