`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HHqdyTHe+PQl8nKYkIt9wdtr18snD5WtELJbS6Rinml3KepPFwfMGCSZ/0SGwo+C
7xyDi3maEaGJx2jK59wReFEJnFhiV4i5McCZJdRqWtkWtdmaJl4ZX834Mj0Bto22
aHylR2IQebAdAyIJIQuoZPpEE9AkymMblrCvkGc8BnN68C6WFDG8BDg2qLJqimDq
HeISYuARUaEbN4fG7OCWq/Qf8kDozbpAiNryZIG4BJUZX0DH3lp6EWnGBLYjeSEI
mojEWW6qwdYzsEDUnl2K6/c9Ts5zB+HdCdpn7zPpj/YSWHPH/X1Caj6R8z3i5jbM
ueOFSRZpweAZu/4HM674sIFWKubfR12xG8nLkSWcIivWkhKr8i46b+EXcuQ7uEe6
5OTS1gs9fzQkQIlZAiUAN8porSSs2JLOT04rCtKU4a2Pldo7WXVz529L8zIWouz/
QupnWNrlNJGOtYkJhLT+ND/TImz9eJUq5cA/WLJAVa5oA3iHaajhXx387B/VD9Sv
briuTotKLx/p9CIdkNTukhh9S+FTn7+fnOwiThVnqhioCUSKkDH0wiAAer6SQW9D
O/BxMuyjRw2pT4uTvbdGCpyHWyorQCPTQh0yeTTR08f2ABjBvwBxckUy1scL0uox
MBN43VUi7MZqc9stUDa7mKegYNi5+aY2bqYQLMTK76HHLymy/IxGDvIUNGdVtDgf
HY4J8aBsFhYEzO+GsxoPgP+2BRvjEYpVx4YjNs/H794f6deZlgsN2Bm68cerLIhl
4CFPmmdLkJZyUXMD5Li2okV1tv7SwSgciy8C3vVwvmFVyPH/7SY3CNWP6Tu4wph5
OeIOTDqRn7fhegqXzFYBR6R0Nk7KhQB5nXM361xOkP5b8fybHilEj8EbPyErFPTQ
t2mzKdwAD3WbGYRFwTyf+9zuM5gquggODJqHZ37vG7cxjFAzZ/4grSfvCVWYm04O
Ygn3SeKDJd83lmndDMU4BmcgyX3R0omFmZeUL00ni9o6Vrj/vqHUJTdLMt6Sxwk3
3Wivwrp+wIRusYfuNYj1V3mLiNpcZcpwjfgNSVpmH0EYcb7k1fCbkZ1Vc5sBhS9I
lhy+8WYlmstMUl/TolHyTZWeNcv5qzExF/KHt1GtzlkC30TTeVIZYmO7o1q5Hk2x
QeWJZRmwgqNUI1usb2x03AOTI/1EbZ6hAfqS+au/4mO32R/1olZEGuM3eJgL+kNJ
xxOK+n/dmZzJ0rkDtpDYNCvVsz+84I3yYmYuu2PSI6ib6q4YEiMnHt/eZRpk81DI
Njs0Iv78obkX+Eo7FwF24DsmyNGanV4IKKaRkOHOU3aUe01j+rea6kAx+epLExXV
7ksTt2MwtcEIzWESI4h0u9c85pqergqtCTIxpaJVve98XdHP9d4WJvsSEpVJVIks
5u0U4Pz6mqyVwkwy0r3Bx0p12XHY47f0xzg+vdo2KXMuonv516bvHDsgmYoaHf4k
cAh/Fh0hmaixg3A52VPpHg2DRhZySxxOGiEtptpUV47DSWfaXkokJCa0KQO8+ZsA
5cKx8zJKhnkEO/YRsQdlE53Wgi87m8hz4MDB/3kPEAo37fgnbOFPX5ksHV/Wmcqg
ALlOJPXhI80/4GfXDuZdAGg3RqvEE6AQ4siaOlhUiqfXiorNr8napFGKMZBv8Yzy
ikPWyEVWr0Bb2DGtJMOcHI+/0VOxHWGUaHpwwgxdh7x7Se7pOV9Pfp8AFGljoHgi
u5F1QdVHS0HRXeviPUxzou+X9NLimHjJNZ+11jJWBM1qfHwCyZ1wZ4mUxEmfXHY9
D2d3szn53hsAyNpfpYID74yU86YAbkiOKqX5MGVxtUwIrNK06djW0PhRqQNWmF5W
0iVv+Fm15xUHjFrcPHKHRCwVBpYSMwTMOj3rmCGA2ljCeZPQG1u0JxLy8Jlxb3gP
O++Jg5JYg3DYqYVYYCZCpSArj6W2rNDcLBJEkuQ80cZNMG1eJye/mxT8SA6n1STh
h0+7YgOWXdK7/xysOmqeSDEq+m5qMDsMJOjBscjZ5rS2B/u13BDlzD7xFAQnxONN
1w2W1SGRwFMuov9x5jbvOlyOZmXbVOUsHnU2MCG9MC5Wig7cQjYuG5UNw9aC6nJw
gJC7jgNajTseCm6CU4uOrywxoKaazmCNRZBOOrR7KNsVQ35jrzUK/hQvnjbMRebh
uGDdvOrLXBXqWkKtn/c3xZJH9Yo0BKcK4H9szOaGm8Zoo1FNYF960rqxUE4GkcRg
T4ZXxKlkOFBLJ4Ma7DTxAeognXNPIH9d6Bt0VmJRp+NHgVdSf1V+pBHUa6tNG03B
tAw1WMYCmsuhJHcEUxhaQBermYW4B34fPzp7mmueRzGkx4yBhMcgpmFrvJUFxqJU
d9DqKajCNcg6wwEhHMGqHRqgoi+KlEeKqnxu7LrD1XicocM1f9U9PnuMYthojRpH
HIY8bJtL0UeFxjt+nGgjps0FqBg851PytPsEFnzbUzMRVz/oCE7xisYZB0KZTe6I
/B0bUyZA4e5YabHTC1lJwuEpub3J40QGOvhfdCkf7bzTewQ5nlad4m7jO1n3oh8t
JaC2oq3pgGY4ZLTBsm3iVAnVRLNankESEP9B5mDuKdpaC1OPMFPXzT+Rh6l6jSgs
EzV8AZ0jdCU+LWnKg9oEqESr+efej7y8+mIVt3FkR1hf2L59YGlG8GW3T7SMQ+xZ
I9RYTIvFIrzpnFJQURr4G0cAqZ1vWc0F0CUwALB6inEOeYYRuefUKRFcBiTc67eE
VvHEZ/6Qq98WF7/0ZQl7GVc274Z3SQBtug3xwvL8U9TgnemDc/ukqT7FisllG151
Spj6pl3ej/r6WGU2nSroOD+ndY3aBuolFWdF7upQHQQAcerFZbc0uWQdfII248f3
fW79j2soqXpUP1Kr+Z3VL9WMotywxHZDGHl7VhmWiBxWXlVTVfje3RkYZukCnLVC
Q58JKOSpBQEcMhV+XQIdSo7ReJEgs6g5lwJvdY2+V8Fodgw5WV/kj8ZlRIbtrXLv
PA6GE18mjGPaVue7eMzj/xukyzCIfITzgagUEBBJ2dfR2qRcmf1unf6Jtd03X8aj
LtLfhhxahdEN5IPTE2KwJIm3RgZDQS7yrqzjYMW/2OHudos6tmpw6otdbdfHMZTT
dHRAkv7LfTte2mNIo2Js7Ssok19ZabCd/bUSbaFAVKeIlv57YnsBDsOQ1k4UNM1H
aP9n+67kuuVaMwWHyjH9nwqtj1Evi4caBtBwtgIiLCW9YAmAYbVJrQpwLPFKa6Vd
6Hvty36qcVfdx9Z0JGeS+rfzXzW++fXZwNNOut2girknn/lqwIuCKyJB+VNIfQiT
BhHzlhOP+Zy3zFtoWcMTeKyLEtPyoHMWBpGEZPA0gGwVLIUrn6Affla1ED1DuXOK
basmD4AVVlDiu3KHkuCoSDAxXMxBWK3JU2qucPhi9Y3SpYim/2lWn/PruvmtlZ3n
G0ju/fGQL7icyrqrHv1zCrV1/JqOOmohajHRFvnLNZVdPycEswO/HZ2f+8EWP9rl
b96PqTZ/Li0zT7WER2o0vlUzqST+EdJuK20+H3NyrAEkyyn5rAGyAw0AT1k8ZJe4
qBZ1rBCC4zh064deXPtQp7I9vTurwLXzuNP/65VkIs5nOakzDo9rnhwXPb0ri9qx
sDTZ5v4YQaZx9PblKH5Wyc0wS+CzdpMck7CFzK7IXVmf9YMYkQb122+EAKB4Dpe7
JgeEWeVwOG1MpaE+GwppHkBCgiarbzr+bU+Y7IMoXqxw93VRYl5l08kTjQpqhR3r
08MWKM2i6O2atzYn8hk/wch8h6gGRgBG0OkY/z3QDWQSKJAASrDG3I3WPYtfY2XO
+pV2+/lm2WMj/ABSs+V0JgKFyNOWeVGjKFcVpbRkgwwLOLsHyEE0uMkGTY4doyvl
PSce68hsnj6AzYFVbhyb1Juz60Et3vBZW5gD0OmFMe57zHR6RDRyIqPFkZW+5Pa2
SSxwb7/nzzfOxH/YC+f2QS7QB9puHaUGMivpPBMG8aBru4WUr3Vhz70aTfjuGIdz
+I7BeTjWs1TdKdkirGQYzRzmeA7QiO9t7tYuQqx4Un+yjpEi97BLBsKs01U5b0V1
bk865VgqpMwYQg3Qlc7aR87z1xZvgsg4xX+RrFvEg6Pt2G4OAk0eqYsC0J3jZ/C8
1zEHirDjA8so7J3P9Bv3OG/PKCqHq/jVMlz32pUQPI3kz0JtZHgarYseuvFYgL2V
g7gC4Eyho9tzj+ppcAhJvTonFGHb+k+5iskZM5yCUUxuaXlgPCJrNjmZKbvncDp1
xQDx+YGPVOPxe27aamsIhRLnP6eGwO82eleRkhtKQ5ylRmbSL1cJB4dsQbA2MG6N
55jC3xSEJcNdMcC8ZqN44QDIHZF5JW9PWFU8lO//ejk6hTggQmMkf7zyHHpgpVbn
gtLslZW/I92XGtMSZY9wdfvdAEDzYko9YqobAN1Ljz8CNrXLxmrPi/yM++tMUv1B
UCMZ7rmmXTx4OuzcUui574Sthc97sAvS0Cks2h+W36PpBMBxN2+moihSiAz2dbqQ
oBBnNmF3Kbgn8gLQ4SmIfWRMZ+YoEZG0kgl0ug4SWs2KhEO2Oy7a9pVnq2uKWsMS
JyqxQ5GPFpAxoM/ojs3SzPpMMc3uwfSvqW+yn3edZpVOD6n9l2K9Zblx+yHo6WBC
5LRQP4Oaf2NdRlbnhhc4H9u5STd1pUuZUt6Tio3P2C0GXeSxiMrokXs5ba3xIfZp
Gt2T07JTb6Y+ROKAyApKnA0lryFIz0Av1MG7Osl60XUKggQWydY5x/Ct6/zn7sqA
SBm/QU1XGxEv1+/45YidL5lFVTV2wlnAsYmj3HU3kNn44nPNHVGCironk7phRxJc
u7oTC7ODqBhTtL7ydfuPlUD8Ejl2zjfzNH6TI9/fWfq1LQsDRlm9kRGODs5+jQ6u
2A0ZQt27vNwsJt73wLE0uTgw53fW2hhAzGr3kCWb5NqtH8gwdmnq/woSFF0QFKvC
BWKoZLYhJfSca2SHzhEKXZGv8oQypmcUDjRCn+q8nzz+k3vbzDxewjz27HdLXrOj
15IDjVdz3WF1YVngig8VYhuRanMiJGTHWbpVEP4YUhF3eEuc1BNr2oDIOGk3DqPZ
8JfYv8wxYejOk7xg462Fju3dPYJU0aSBBD/WleMohhT1xiBYMQvueLqV6lneVmXC
vZaO50ZRrP85Y7QkwNA4gqGYcsFXexnmhvr4AFF0DID6nOuZP005nE2P98IT/1Dv
GGR7wPo9qEcwbsDFEP26DTWdVgwwvMDb5BokyzjAgLJ8c2/ywG2D6zEiv/LRDg/y
iO0x+yKqEBCcMcD05YXcVwpFlt75141YzdEUoabSK0FJiJILnorRIfiT3pjxMOdz
jNsoe2/pofOADns6/nSLBE//48aak8024z+PlTvbirXMqKzupX8Y0Rpyk9imyilN
1qSVT0Tj4aqlU/S90ppc++ZOgqylL7AKP9yrtQJpFeS+SzWx13HpR1vR4nMeHxSG
SPFQuPRccEflX4ANsP3qeGFnzJEDIM1NpQUCZowg2naG/gPDUQUxd3120lSY1xsc
b9+cMboJlHudnfxdZ5QfGc9UVzEZRK1n3nf1HMH84iEqxVUJJJZYc7csJBbjvEXS
YmgHOeJN97J7KTpA/q2EIVnxN2lRLHVaKT7zwnIEWnv2Rxr0jlcDBs3BNNnVG7IR
2nhJeel3sFK5+kWAKns0JbgrvYyJiKFDe+5Mt3/bBjMRVmRK/Sgx9RxEFGTGfl6+
uGRrry+zceFOARoSUJVhZWzf4VxjWCDkQdhr3qMgbi/keVFa3SpqWwH+AjLSMzUl
2dXBVtsb0J68JZ8qo0q2Yrtm7mdJ3WqEAAkZD1NHWHNp4x5t0+SV7T7TrkXK2egA
uINqdq1bnpAEpKb7TPBUyJkkZNjhhi6wnPBTZ3P55aHa8wYjaoZXn7GrgQCfBIca
L7cxPLtvGWaC5HdFn/Bp9SnqBHvhocu3Unq8p5Yltas+QISn8UNecZZN4yzPlv7x
9pmYX0HSHkYZJrziVciSqOWc81DKwTZHBXgAxwO96aiFt9zXTevD2feeVkftxu16
msNq3FPwKqAnsEMqgF6jc8ynvNy6LWr5iV72lyljJmBHVYjMIskWfWFVhynyRY2y
IezFZlkifz0Zss+DoGDtXjv5lC/qYkhzAbjkCqrNj+bf4casMjIoeaESMHRuR5rT
srLTkW2dfBS7XnKCHfLCLgMf7ntUirTt4o5U87hsi1Yun339hErFlAqOSZCCAWD2
Kx90bTvO1OmR77PNIXr7BR6jjckJwSQPNFw3muY2P1EmngB3XX8EGBffz5Kfw3pS
qX/HHg0fbJRXYPns2wWdHbC3N7rga9EAZK2BJCvSKzx1Ac6CyLjc9EaoS/JbqzCD
Bt0gTdE9Wf1EkcNAhU9bHlwRnLwz1plfttD/rXm3d8Rsxmzt3+2RLuAt8llgkWRL
uXiH8hDZ0dR3oyfbSHGiBnlRhjNRH4ZJ85ow5OKdtEAU/afyEulJd0UiX6Dv9cVa
0VuiSQfUbEZOWrPSR8hjrioiAdGQj9yvtVU69VfqoH/rtSZ8SCwiVa56wu9Kg1f5
xbA5nhkoyOnuwUoYA5M3x9dZyBDWk0Kz5AbrhyAAEne/Myl775T627tOxQYntIRT
F5CVT4gMWGtR6mrVzoj/mTGcaibtbFcQYBUzysF8/fnefIGUaKpUpwlWQHooPrhh
UTOk7Owo0AuFC8UkLCw5/VvSRheKPhHNsD7WkUvNM3b7pBmG/qo/MZVy002Rs2zI
1PZEaw3JXpYfOdntPn03CnrNA2RDrwhp7OImnfJEzO3ThyiTkZ99q4b3NOMNaaOO
XPE5/WzRBx541coIowdqksSKXfqgaNuGRvSr0ErtGlAKPSDlMR3wkSpZNkeeiHOd
8l/bV4d46VNq1AeH/x61bso1JbWMu8q8Dd4/80K18XUOPRaOl3VJB3AzuRLB56Gf
YglWNtWJ94brcWMNvxMpQM0pI8OtgYSDRlwDQCq1T6NL1PUOeCK2YBx+T1tKNZWk
ml6l2rVUeBnLAZ5kFwOGFudtMXZbtsN9LsxzmuSWB1HUhCdp5cIrocxUBZ5LKqjo
AiZq1beVl9ssVHXAOQgEFmCTtssT14YUbNwS42Y5kfIJfLc0RcSd8k5PH2+asI/M
hG+ZZQroLbSv4OfCOoplm/+TJ8H3PUcheVv/FuTGkIEL+P7ygzpqGyDchwjf2VDH
DO0xEMhxpnR/W0Gk+9ct3ucH3+J8CIKGC7q2AXFqdCxOzLvWIzMkNTxEpIILXFR8
b+mBOg+bXOVHgxgyVqEn3kPQnaf/WnEDYEf2W7VOa8Ya9Jpu53uLk2LbwLIS7dTv
s4aIm5QOoVJqf7ql2JI7AhFkq5qu8VhFt2ibv47lTYszJ+7n2NLLvxVEMuHpv8o0
GgfhCXW6usG09yQDN10Bwvrx/zV/uo37dRmoMrLDIKWOLzg+RAtfVsoe4bvKBhgM
1DYmFDjw6xfW7zkK3ewZSnHOd5j2zE+5Q2gEfb1zEiTBHdt9O8Hd1HkjTGm75nbc
01ZidG3R7SpZ9hyeTdN1O+u4cuFH++Qio8X3iEKqemebihQOJEWArbcvX/dW6lT4
04om0mx3g8rJUIYAUGgLqdFYu7/7y3u3y30oHyAOKXcL+Tvho19DkN2utIXWJM16
PTDOrqDDEvWAf8exVate88AA7fLOibCRCti2ksaPh0snHqGmOsH1AVsq6srLy2GB
OjGW/+3dtsJVYBwKylHrxaub6mrVecY7Df3jy/woDiOyvoaPBG7j2fhbtzjHEEEw
Yrr0oDvtt+lZ9V0OSRay2ZtkrxzepTC1zxNu0N8exoeEh3vhjIl+36fx7Tf+kff8
M3SiBJ8hbXElMsgXGBL1NepAWb/QTINlMGx0KATRNO7XsoUNBm9OgFMnGh5aU8nU
Gu25ghItDLlgA1buDX5mz3OF1FMxx9PrdqC+m+KsH8FpLZFm2uTBLvMcoQ4HOlXd
kVWQL01lpjLHQYg1eGL4rfrNuEdE6Zg+WyUFscUie2Hw1OKye/SVBsW+Aon4dNGY
2opINJ9m4ujx+4VMYt5EOhNb5PUwxO7W57s2vR/kDer0r62vlUwTUvQVtVfprhIJ
ftkMKhkAstVwlu+tHO8q+rOxsj0Cly9rP+G2NDtybSnugcUkPVOIix0+W9Gv1bM8
0oM/H0pOtye2aw+XF222M1tGgnba2A08fMo8sSN3vgoW5A4Jr3UwNbF7H61qnk87
DA+/n6HdHWfdiPJE647MvAEpYbpvVJB6Mrjx/3WQlNDj0Tjy59Rf78czwYTblKCW
RVEJbd1oXO84Oj08UggDjmmvAjitdpm5SKSy7eCCr2d4FGbZEnQJsAhFlkgoT/2k
k5D0xYCQlSu+3uWIcRK+mHFNEoUmgTH4VM0+L2cU0+LLsAStEWnKEY2QDqcPZKf0
nPxM2bZM6p4ot4bLpc4OsoNooD5CLs8dDxYiEnPWd78REYygrJFgkigqCQni/3rp
YiJkqc6loGXuckL5z2u1MIkxPb9wbG9Kcc3Nym0dVX2euCSSLISnzmenVhlQri4E
kFCd1U4SCbLbtNXdn+ZfGmWsSp0LQDFO4FxliRUNZXAfGQy8OUE3yn1dCCr7OYpz
wg6uUaDWkc1IgXWemEDiP5GmRbGwt9mPe/+Gz5jpf0IhHjevqJx+/1fWYS/uDpBq
zIYuhx+TCzgDaisqhuDG9ULym5BlE9o36QSXNvHDTLBF5knq7coknlLL1hc3H/gF
M0enzcc6k3PcveY6cglBpn3VLhydvYD9y+NH1O/7ctJcJ+RsABk1my2v+8a2qznk
fDzoazQPpLKP1aQLP1RK9iu0SUHIckTS3U5eO5zhQIYuudeSn2BJ9+0dMNegHrhV
UM/Ujt+9oyd9ylqkTeecBi+hqvUqjXz6fqtoYt5biRC2tLy6c9ayxX0XR5Yjf2uX
p18fW6o72JPzx2+c/bY83ARoxQCGjQyEEKgOJvPBgHyVYVbnhr7VEMw+45VjQb+7
KeqIcSLbWD75R/GQLMJFNEJ1KvYakGgju6lh0nWHoPJpkOASNjE32PQlwrHPR22n
AzIAA3B+2nEgEC1w71w2wngQHtOaVsOvaCgCkTUNA+i2xGS4a/eC0c29xAz6BJQp
i59xn6iSTouVKLHiGwJzORXNUNU02i88Wl3X8kDhgTnCje9tIdZg7Us8OoGj+2N3
BqzFnR6BPnhH+IcaO+bm6Bq0IgUxc5BfWi4o6F4B45sRsN4Vsyy3CEcRqlUdC302
lUXKu1Jt7ljnRvd6Gj6ag9qCE9V9DKMMoF+xpMAg9O80/fof44ostoQH5AMyauE0
wwpZJxX0WP7QSM9pTQzs4SJxzfEB8sZNRjjRjBeqYR2d5DbN7AaiYYYT76mAtVFU
WxUhcNUbvNxcVDNXYuAbT5t24SxASi14wC2BPoc0+XjZ9mkigV7JilianYdP4Nee
lDte7j2jX3rY2wWAW2mPSrBnqGvgsSY5s5iAjuTx4u3BNEhLwbMewA7yPSxZ12yx
QZ9vtXVQQK4EmaXbT0aS0wBpS0VNkcEChoypZZhX218U1lhsP2Fz1rFVYo1thHUQ
JDG/v65Az5Tqe22b2dcIRXoKlxbIk5WHXSqQ0mwUUn+10bg7ZU1whxwQuciZL5sb
+MHvsTURunUwK67QHCzgFsPmnT6KLKQiI+TvSyd61KIRdd0ZOfnhd4q8MaDJQtNJ
lAPDqUmBU2b0BqZzMIZe7B7inbAtdIZH+9YkouWL0ZgFLojs3BksttpDr/wXPA2T
cyxNugnKui77+vv3phhgOHxnVF7p2cFGdpdWOqADFJqS1EjtVnSml/2dxYxXKxcs
zQU1I72FxUQIClUKCAFt4cv6byV2fPMfLDnHjYQzNoWjqIzLhYTnILPARph68Xnu
3n/Bfam2kKn0s4klHXbd45ffHhjHBqlN9bRkVJ4gxDXRPwy/66x/J98DGi7/cuf9
XaQWhcx8wPhPjHbOgRATIjAFM+FUqj+W/15BvVkWlcEeJaMmobv9eUtGOrukXNvK
Q/mHpBAHuoLYiM6SidEFEbgAam0cvDh/LeMDmmG+Z5IlcIY5KTfpMAfUO1gepvEM
tRyJ2w5J6yTxYt0YHd/qo9dZsz0tphdH8PFbsbqFFI80NsiuRqy0+HQ3wawsXf0G
0bp3mks6vAyVYhmhQ34ats/WE1l9ygR1yd/KFxf2C9GBhOEErZdOYWNyt7RY+M9g
TwHZwvvA+3LP+nirmB5OZROW5LJMy27cWnO41XaV5jXE4Y1RDXzKr+YaBj7zvow6
9wQDwn29yJNcZpeeBFzfu35fabrkZWPPt751yK7G5UPiJF4RUief1JVkbkQAPiJ0
7O+Y+Puskb9cA4fowM0xnF2w3530WlTX4RAAaNM37TzAVe2uVlQEUgubMkZx94rQ
LYnclw7xIE8UzMZTvkCXrQyQFMgdBbBKkk1RH079rbeRikICOVFLYzhNVQNuiTYt
vByLE4uYZhEUCRRseEqg/ekSQlpDfjRSzFYCzl6xG0CAefPwnRULtKCPOUIvyhsa
FzY4JS2uqSsrtN/DqIoEtM4SGEFojgFwP4q2+efW8IWX3jIvcjTmh4P1MCAGVw7A
3C20inc0FPkIL+EtWaLHjNGS/gaaZLvTg1jbJePEwAYUMJqIIrOFDi7tvMpQ4g9f
BQMjylCZqTroLq5NPo8m3OFYmKn66KQmxXii4w20TYhI2B7e4TPpiRqtbJ3//qHU
zNvbLJGHoZvxb6ui9HjUow1WoqpJ6Cv9mV7btFFN+nNoUCbbq4cQKKlKkZ5XBdgF
kZHq58guDnuwllmAW/lhl9JA9KahgtpQDPFxSplkluYOyEL/iX5TjQZNwSwO9LqB
lt/RzCYziDrVPiEcfLM9zoxy+0Ta4oGrQJdyfjn++iVJD6rBWU/0qAtUq7PBH8YX
uRhQxlSII3KeIvjZL6wh+TCSkPR9F/J1z4dxzPND9sU7d8BVBhyiOwfrzlMXlJxo
lu/8Sx0iDD/ATtVNFL6ewbtrONLwzsnlgprWT61FalNO/3N35tbyf9DLRpygXKOL
0ptombygu+clBK1HfvrUwU7GwgEkvorLuZjcWFys+r3lZntu+pXoNsqzsALOAiit
351t+mIbLWMwUj8PGlwq1tTgztpPbPSIrBn7NCqF2HAn4TvyMGBVRAkyeimULGBY
muo7iKMMsM4IBNNR6Z+zkBFiSZifrF5mv5WmoQs5UGVhks2OQNJmvS/GQeBIAhzm
x1eBRdjWLd/emnDCEbbszcULNL8mWFeeLUWZm9DNjPzc9aGitUuIK80ER3k53XK1
FKr5todQxCEwPAcJlAW1t3UVlaGfaxG4OGqkPOfh43q1r3e5hcdHpJB/wCB6a8DZ
YpA5E87A9R60sYbRuJTpmVRUN9CrWf63HcKQOVtEHoK+fWfdWODTLYP/1CnezXEY
li3ZaOYNy2AmOAfGrpofpXpnaBN0Cl+0w/gvSua1cwFvCTk3QQ7ac6E7bbLV5iDt
PcW4k8yRnBERT29SS59j+pLxDu6IgvWTMsxj3LhUsHHpcgNErDJ0oYnLjQEiGgu6
ZRQmKu7Oo5BFpH3EyglS7iXEWxCeKkID6pHY0bZO50uRcK2AuiBkdtx0yXzelbox
Oh141m5yCOIw1LXmTSrjeH7jUB08ygQoAmp9qrfm3ib4SBk2sQxWvxYYfHpKY7YN
o+3acVAZjy89aLPZX6MFzhx4QRTz/OQ9hPoOnIRZlpa0ijNpVTpaW+l0eWaGfp86
bFkCRvCLpP7Ei9Wa5qnIzcNODzOTysO94B8Dsr6aBzWNBc7e05NJTANvd34UXHSm
VUwTpsDSAUjAmRX4GtGlLxS91wT76hx/6p68Pdwexlc4xLLeRl5EWMN4SQciBWPg
Uf+YT2F/0DNduDq8edE6b2xU04bSrHPcJtqOVtWmCGlKryTY48f0scj2CVdWkGhc
qoa/pl7+JwDtaVPO9zPf5eYh2IWBgBjdg2gIualt688b0/ht1ESK9Dlqy68cbob6
qDNhzzgdWI4mdm3yCVZFcWKwwb6fQEzYWl5ZlhLh0UDNjrKLyftg9JUPmRGrSSDE
l1pCKBxw4VWqtb6MdXo51t29GGZFjiOIdR9sU4HGuTat6IXX77OBK8ReH7GaY8U+
goN+iJFpUudUFwQ4NoeeSfaEbXVrpwPJQwZND6MBh0hmc2xVkgseMWkOQ5geRsTG
D+a471rjF0tPr51o2ZWdGrN6iFg3yKKDFsz6U2IGQ9NzeXzl0rzUIfT5MQNfqIdO
P1s+OAwIwFKEq1R2ZH/AVJklDfoQI63uYIFnGpv6/NRoE70PudnA11D21F1IHYeS
HuGrAGwkHeAVh+K1k2MT5I1sU2tMp9mFUmcn9D6Dg6w6hjRBUSYi9kXbrMAU/ghq
uynK1npH2nQ/N32VY6DcOQF+x1fqQc95gLWreFJd7Xp4PzZWRoWNLBAV3e5+Rau9
yyEbB3SPpEQB6bobSTrTJySpTglGThwG2uLs9Dmps28cTUcOB1MW2Ih+O92IEJj4
xrW4Bfi5MdpDPHA6Oj3hRNK14/lG43+CETFtHWRO3ooiqDrSbRlGELiwF4c3OfBk
KHkALgVAeNQZZj3vDiyW6bdqspqpuCBPGqyivPdLxiuyFbxnBt0H7xpZaQXOyL2W
+vx/3f7u2z+OXm0I2Xj4O6mvfFnIecEfPgLdAhY3b5BGSqqeMFLCbZXVDXauWH5a
g7BnzOOkfFZdlyc1nGV+5HFp5J4effqfbuUBGqEqJz2Kjsj5nBHSOHUAdKo85/v6
tgbExxf1RUDz/D3oF8pwfuQ9oRonDo1JFCm4bIFqbxTQJME1fmCMK+p0gClLUs19
U7ibNFgy5wyomskcdkypow91K0JEshGNd3n/BqQ+/ixuxx+MxIKUo2r50xRg7HYu
rSXo2gCOw85s/ucF8B2th60XeC8bmxqcs0xs5Dh3SFjXgmdOHbNExi43pI/tfrUi
NEabi8x9m6kw31vGl/Tt42326epQKfegsWEUAwEjfEgLrlTQfzpaoBxSvtkDF31u
EJjWjxfkFVIDkrE8dFDfax2V+OUsjw+f0biEWOn41nSR2eqoTs9tymd6dz9Lj9JG
ILtXpWSdHiaqVPoUlFLC0gk4tIpMjV6oZ1Qn2pd8aD68fo2da+oecH5nBAENs+8f
+Cib1nnNhy7km1ld5wWkAPe7vkMhqVCfZTa06hOUXCusiuTp+mUSE4gn5SbsP8h7
sRGWYGUyvrB/Q3sRb1Qehjx4Tubo4dIEZmf0nRhaVg+gTeHdT1vdHVoZlt38gNGI
W/x9O/xZLGMdNo9d7kS/ds4CuKXqSxr0H1JOI0ih0Nk701D1xvAvqObGL338sBr0
V9rZBuDzpvKccUPQE0FzM41zQUHNCnxRahLNSIkTBSvEjb31d8ay2s+JDChLl2KZ
2xT4ZDrYnnxMSig9G9FXo/W9HudU0Qhzotc9uDmcfky2j1iS78RyHdxoIy3RClr5
XziV2eTT8PcWl0dcCPX7qjoNZSQv7lyzuV8qeCERF/1DCV4lDkXkglmnKehDBFQ5
Q4E7t0H84Fyp22r4sPcvs2z/aKCQAG49dFY39ulB+u3ezELfG0MtURav9+QBNl1j
AXEQxBA0DOZCyHAZl4uShOA08EzI5nKlAS6rGLkUdmLEe+4xUMK1zk9/giSvludo
gFwjvyYdfxsPHi285EfxdBftAExnwjbiF/QAt1mZSgABzLw9KAEbpq1QI5fvbLv1
lkt9QDY2sglHsHBuJx1+bpxSjJA0LHYGTo1IbY4E0mWjZNZhRct9lld78d16m3t1
nKfiGFEioJD/9ThsW0/yhMvkxmtxmAgO86a/rB1u5KYIOAsFWFhPK7q9FZ9vvu5y
DmbnrY1eHJFbU8SXcGamaLuTvJ/vQF+ibp7rlikV84yLZXbF5TSajZnhNwlFKhZY
arHRXzaKYcGaA43+Z8/sIv5FHuoa79CX3W2afQIgFgNuWTvX2NfvI05QwHoEaXaL
24JR0CuBs8E1BeF8K83OuB2qL932oDUmct8w3MiMVsJ1ACkk0HrknYDdiP+KfBU5
D1r89Fgeoks3wrc11GM43ZDzunwz6oAZex5DW3xnStrehhrUPze3EUSluGnhFCYA
Gs3XrXMFXox3usZU2K0vup0T/vo+CtBqi8IvQWkKb2Mc+g/0AauDSDnnfyO3TJsd
+A2qbbbLNYUcC7bbycsjj3XxiQy6VIPUgx/idCthuqSXsdOKsPe/CHCKMEzlIq2k
qr9qWZoKBZXrfx4dEC59ySuJCNCk7wwEkP/F6KnWXCVsEHXuyfixuHek5kFgRbi6
699T22bDuyTAIo717Xtn6jiB4j+mwC0/RbIPZKOa8gEZkFUXh5Z3SMIK3DiNW8TW
d+tHYWesEUcHm1I9B5KwaO9lboEBc1J/1TxOsxjQ554YFHI9OVgszbtZ6oHFO45j
TqOsSFZLyotcYz39g3UD3TukgyWobTrV8RsFXsU6l8ZC/Qgkx1oy9MNSRglAFokZ
KpVDKEBVfigE80gwzMWmvi+baTekFRO0jAAEokESjgWNEWImIA8iuRLN7X+1JrR9
QvgiCWNMqbBkQRAB0bTeBsy2P0iV+AuVQufGpBOesU4=
`protect END_PROTECTED
