`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JIRDTjwziUyDaEvxCXN4SPcIbWTq3Y+bs7+celZ3L5qGFzJ+wQ3jT+eTi4rHiBxD
kdwLMoIX+uKUyQ78KYmYwmD3dCp6BdEusxU27TnEYwvabTTPXqQDTGkvq5XAHtqt
zx5Ezm/QkDbv81nJ4fmGabwTnzvOBF0st4yxbvFsNtQCtTmpbZjRB6gKkIIJuS+8
A4lP8b/Nh1Ll36wujQAx8xB77F70yABE6jt7sIfuSvgS8IJYszO1x9hSuZ/U9ZR7
M502BrLTSCUu9ShqYy989JeuYEFaqQL+jBpPjafPhaVUDuPd7+a5Ml+qwaI0TsPG
ZhFxZaFtKEz9d53qI/NHkg8qYUJdIIctiXjFvdnAtHj5rvbi0JfCuAMHA++PLP1/
s6eP3qvVEfsU20ti6EFDkNvxFjdeTXl6lIXYTYDc4ctnYteCkAlxL5PPeqZYBAXh
TiirtO8ldkO4C46QqtxlWfIvml/yQfU+h6k0+Zg9VOAu+3q9kbz22fRVdIpM6IVA
v/aYrX1JTFZU+i9nhQplJYd82yHhDlB5/mYmoEQ7rrYqExGyUh7Sa3/fLuyrvzDe
QwMHVI+xJTjS39olBfzyYkClGVFfJWW3PR8T6jKslhxNEKDxiaSyYUROp+bdCgm0
2ePKla0ZWWOb7bsa3ApJllmLcGMV02y/nrU0ERR5aR4Qn0dtRetgKt59caPQHgTf
wcCLemADIfB+8TPUqdAc9TWQ7FRNtGCO08ROOY06J7cUvSpcYKGskwCE/szPJZQz
wuj7rQPiICf7kjUZM6b1pkpGyHHNGWqrZOguTYgm5ig6yHGQfrK41043T9tk0CB4
RYpc43uhRU6VsuQPT/JcNsSV5V/Mvu+1Q3HqdmTTDDmGlr04AwSWsFPasq8Kmhcn
VhBOt7GPGQAdV6jMUZQFrWiCcogBpzNqZt6wsOe2870Gi1V5VYLA7erF90c4nF+5
W7JO1Sgo6j0IMdUlqaFmdvVMhoK4MpeS6PwT6edzNa+tjq1QuzGH7L66G7h/glil
5o0TkAvtV2D6nJwTBPf9A7NPV+f4+6gJoVaQJn3a490utnUuxcXWheJ1AplaWQMY
3QIIqinSE14eLIVyYSF4+eiJL8gCIeVYYjfIruJrYZcaLQ+nffedApf8lKb/RWqk
GpFkMTy5Q8ZKQQF4/xSAZ+0l7hen+ylaKzw6EIMFOq6F8TxdZc9vKiMfcgEGA/Bq
a1bx/x7V7TAlwCOfQCNxdWx5PwH1nb0pcGrTF/b39p9PgB9gXUew6juGUBxmgMqq
fGMzOL0tJ88x+9Y9j7Vpn+gMXkJbwL13qN6by8oZRS6Xi5KYejUZ99HpTDxmjlVG
tH8+7kZki5YZRXg+HhMzpbeWaJyBOnJVoU9g7lEXaeXWvzoYqUr+H4m8Xo8ELA2B
COjIXE06R3/KjS+RXLYOBLmCdIXUelKJXRu0Dfua26FdQrjwMKrsVLS6R/lWwDJ7
874/bT+C3s/wEjpI4EDr6hVuSxkvQhYbgHIm9jFVY15Kb9hihc7Ov9Hl9sX2KMvJ
9l678PGz2ZqijgU/ddwrY+hFDt9PL3JTlw8TWrATVlGkYASQDv+L956tRTdZMn+M
E1T1nEFrh3T/4cHGz39oHNcPDEK11fWbjxBsjPCA/DaDxglpYc4wu2Yramjm+4nO
6lI5e7suF9lAEkhVPwS12MibRI9BJwmiYc2QHO4RaiE1yj7tw90BvuDpO/XmzTym
htxgtg0tV6smU5vNY1asKcrnhYnw0jVv+lE0H8WPGXbdAKFM3OvSCmVCLgqrkwOy
PLfqSVEV1bN2zs59MNMr5pTaJ2PvbJATZmHQFy8B3n6zJRtXQkWp5aIUe/XB/c2g
f2OqA4L/HvLuoHh4FpxkSMXKt6S1eNpATc0mGjPoppPdmh81oRdod1qr7gxt2m1z
2chajoZ4HKg2mhjYZJJZU1Mwdiy7ffOEjn2KpZTFGiRF4gSWuNNe4I1MUsl3wZyk
hcKps+YdKonESBLseVUVIlnzjjEuYU27/mbUSJNCFdd7pbX3MZDG3WupJy8ylsmK
NBQAn1MgEQBAX/Od815yJqkYuFRzrlBR2ios8U4vnZ+ml6HdiBCAYRsCLdtNeMyo
hEhIzyyBoKozJfmaxZiUQxxXlpnDK1tOiPXbhKLoIgX0X83zMOonFVEK/taFO6lB
HggX8DKDD8vY08ixMUCr/lWDiS5iLIsJtDbfruSIFMPRPZ19hxJVwRjDyKUCDB5p
C1z4Vzg1QSNvNRsqBO0054oWz6VNXbx/qyj0LKtaG5FlrgkpUtJc53IWYS1+foZp
C/yfgEItl58ruuidMaIBhhsZ4pcZXjIeZzMhq3+y+ytv3MQk9EwyLkbx/y0K5gDf
v83aY0iogOAoNwW22/qFjQ==
`protect END_PROTECTED
