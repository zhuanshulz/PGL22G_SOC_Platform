`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DWLxrqDs0lR2SHYvYT1x0eAipTJQDpBXO2VkGS71yW7Xr9KiitFZYhBxBVoCZio7
TVAH8l5Vz6/n160dsx9rgss2u9O1l0s0hLcMXEKPipeKkDTYA3C7YHo/A2zrqIDz
QbkQfCyrf6d9m8rDKB7w3H6PlZfb2lyWjmPapywkXZcYYUyOGx0pCZ69T/Bs3o8l
HHBJ0B8VRYR7EYKBBJ/Uy5dhNpMxwOrN66Y1ojoUlUGeUrqijsYZDpgPah5CX/yB
KuUTYKfdbTMki8fZDibUxXJbsBVgzqjUEcZrZXWnIjn0MprKgbOvD2gA0fxw1Zjs
qNyutxmj/BOfk5N5cJ3YiHsDwORWfRsAfawiW3r5nQ4=
`protect END_PROTECTED
