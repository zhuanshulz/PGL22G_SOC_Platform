`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WMYD+tTsDPoLhlCexjaFgOGc2kkLnOwMs6dJrzdu6106grzJXMWn4tiyV2EsT4fj
f3JpPLD7V2/k2U9DWOTQN8cpJupv6OxVZeGdE3w9ucoDjQJcSDC9+x6IY3FjWYMU
fYWdR3iNGGmixqX+nyW+kQ1Ah4yiwXFSwwHWG70GLrHgRwezoUvcrmKL4HiEBneh
ggZwJ2dnh/MdpGNY/9ZLtjzGqtpip3VicLrJge9z2cgc6GobRcC/gwtGBX+cyfJu
9ZD6xFORCYPIx3lX37O5L5Ewo93YAT6FVkIYKLDmFPKxMTmw34xpUaQFtnSpgrPv
C/I1XXkDpBD9FYT/5hyQszoeoX04YfFO26dBgmIi6hkDkRq681/QcoRrEsXGE7tR
MitgFAF0tiFYx/7dr6+crsayEgAow42NRpAQKbt27Y2yETQqrjWy0syqUsNr4zPd
BtbLaos9lhJgebSgkQHhjPEhHhnhTEO0aqWqJYM1Fe1Dh+8qKBqeAT+0P2PyY6Y/
YHRQmGByAUQnTZMJqi8pxhwgsiCr+SsWY2a7Q598Ul88svEnY9lniq9lBNLW3+pQ
73i8aOfk4VQ7Skk4RkNPpHIzi7MQx9TTRURdOVU64cwMLKD8iEXRb7MBNOGMvWW9
STPtC4TXApIYImjzRUYg6KGJ+fbDmJ1jlBR3np+3B+5YH6MVz/2tGr3JP/FCi+7e
GJpfEid1hKWQCjMNOafotBiWXmTMUPQ4aYVAh/BQTVfW6L9YOXPcIx6t3e1RrqNo
Qqig4m8yN5kAFgZyUdyQQ0hjAc9nAQfb2bgGxeQ72KWxTYjbsjPj8a9JxiOwYke6
J1p3brVzyktrjpgdE6EbNiPyY9DHbI4FrnL3VnmCct2DevJ8XOfxTJdnsLFf07rR
v84yvf/y3cdpEceZoFDU/Q2Kxx5MF2UyMN0H3miAPxN3/LXo0C8n8FspNRXiRNhr
ddpMEmNDtfDOFX5kFAsBoZQFKBS4V4e/G3wq+Z54PcYwCrSQU8ruijtfdXvvq4lo
scsoCnrJvoWD2FgNux6QYYNYo+kMIPhVcvLqrdOK/t6x6cH8Ar7TppKXR4bA7pNd
NCETrS/xEdacV+TGysnA+X2qk+vPTcABH6FbwAp0XdennQYaOGPAWyBXzQfgwSx/
+LErGlvhGQ5POGGn9m+feVMV5fw3kxJPamvv0av6C3RfyUyPiiJd91wxOkwP069z
RHDbwXaD8PvVa7Q08f6Lzvh3WQdeF+UYdXycLc3a8KhR5Wt7QooA2QFLkeNVpdDm
yUB7DjsETSvrTz3Zm+x8xIg4ugnFm/BYRaIRr1tO9Kw=
`protect END_PROTECTED
