`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AgahxO8MoypihrOl2fEpiUmN0PgjSeBj6jd3r8xwn04SkxQaBeuSOk18A4mW8I8W
X/wC1nnctkkdM62I1y/kUcdw+3N09AlINgSLaPmXrHj3Y7GWvDZ8ZeVulBxQTfAk
uYK/RPCxeNJ4nA1O5rG7L4nLZo11OXHCaULFwkKtkd6hqlsKYgJFrCukXC+BMfVf
WcZruv0FkCWrQ2t2YqcEn7oPXTH7UBynQ53jiTj2LoFuwHsZA2yM4NPhf5tPGSxe
IBTHxcrBwoax4VaXisRabL6qAWcjSJOWi82POtFIrBXBK3kNFwL//W9bf29h7Uzi
NlWFp+OgcC3ElqEVcazWTeAMugK6h53CfZUHlZs2lf2WLIhAwcHs4F2e1ICcInCg
ttQIesfMBmFOEbFwUuaAutyufbnVJkVY0n258cbWS+Cq3/jmegqX0Jau3ZdDtI5B
/Mu6H8kZUxOFmoMiJI09F0lZjCf4h+M4/3jNVKVeGbjgJHPnevkG2Y2YOwtEGMJ9
rUWuhwNVVnyRLXAk9JUbZr8N4DPqrp/evt2+vtI/V8zgBTxXTGEuWduaAOn5BqVK
o+BxeRHTXkgVH/4+3Bp/ab4wodUL3xx2QfxFQR35uP1B9zrTfhw0xCTGtcT+GyZK
PT6IfJzr860ExPS13FNI+WsVERBU8/WpywPTqQ5EZb8GH1GJczahRsYuPCa7ORca
uxYp3p/cwOw1PQFTbPRRGWZc4Ri2bl57En75MFHw/EB7GzB11UzVuVMcU3lSSpjz
UaLTbpP53P/kj+kBWRV3LQ9cNkL6C9bfzVLaEvDMIz9tINCBB9IVC5i8ICWmhsau
`protect END_PROTECTED
