`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4TrJzPj98tFdjhCl9i5WhQHxkDQE/0hjOyIdTT6YyMfvBe1I670hSIPJA5JNS0dI
Suye5Y7frfPWvHc6xGaUF/hha6EH/NpmLHJJoA/LUj8zn4S2FiJexq1Qd/450dQq
OZ1Hz12OvX9q4OCKB9H2LVmgEBdiZB2O06rsa5WXRpRhdKLk1DbTosUCvBTx6Aon
LZNW4ph8zhbFLxJZ1yv3wD4ndz42C3y6dkTBhZ75kRxRVC8L6O7i0uQH+jHXQfto
S96fB3kv74LK802m9MaLqhN5aQJ86gBEHnbKtNOCNx2x6a5GEABjr+hFTq6x62+i
iovxsFuHMSySzRsDuwKnS6XRIiUQWCSIjp/14cFzfgPCw2lK9BDWHslPdBJhhsi1
uFbFqxUYo93Y9qbiZW0QEWWdAHIt1sArDA/OUIeCu4VOap80936NJMRhYIvbIMqm
2vWqozto3x8T5yWV+o59lW0DP0vbJwh7HePkvkOn6noIMPMOqcQtcJf2ls3WN7sy
Q/mqpPvqI8f2uxDbWwTNtSSLyTAMj7lo5UTuwWTDbOgCEip1abSuZumU+UeqFU/f
hbbz1r8ZPhHtDiKJIyKl1tCgwT7NeNu5mNDiInpq+Uno0+CdZ6xIDeAAjA9IicZd
i9zG/7RDzKF3dG6QGs1WiSWNxOcL6yVPG5wSpuNS/0aUdbOPsWLv4PzD49zt1mBm
Nz0kCE9qFUmxUN2BeiVtby92goTg9TqAd7yuGnn4jnsKaWEsi7CfqsgsQVpHdiQk
nBOHOl1DD+QJbPowLdvYF6neLcu5KL2qcb8U7LSvyhcdlgY227ok984wrgtuT51v
ueHY6B96dTmhcoBq68oxfVn3DGSVwu6fmLb9uQTQ2Xg16bDwVHUJBN3RssKaid01
wZQNCf88us0zAHvR/lTof5OLcQpzhtEqXDFJiqmp/5zK5qDed0busNftR9P0qQoE
EZuDqc3kJ4s9fOxMZtZTBWBAdTnH5l7YincuO4Z7XPh5cx4RpBAc2MusxDtLeFSg
w3ADTmcVT+GrGGIZNheXPTNSnzr8WvdctCmcAUfIMQer+OW7A0Ah91ItJlfPoDy3
1xVkJ6BbsLopOiTsudDAfLE11jPBuIc1lDPh97HacvnbCgsmJv9Y1OEeb2cyaHFn
pHozScna4A+3Fr/CDh462uiHMF34J6Ra4oGN+qkyWVxnCy7meTIZraO4Z7ffVcFO
IBp7SOwP4jTAUAJ+9ry2LvIYy4Ahkx/L40/Lul7H2f3iRuTkeIWyETwzIjnKsh/r
maR7zJyWtg/ooFonsVqNWmVuiQLe3OaFrSME7J/DfPmp4a89b1mpQHEMBmlKhvwg
4SGWeJh6opc4cLthtKU6UJiiSjWQ+/Hk/fWZUd8Y/U09GicMmzKQ25GHqOOKF9FH
6iM3njvFysAkbi5KgEGbhvgjvim+gCZTuwvBrcuyzB/R1w9OHHtdxIku1gWzCO/2
gPwJbZsXyFPut/gl8n4swCXUSb4OUEq8WM8/6j9y/Dn2KB0Tj9FiG9OhEYYDTN6z
7OyfjLP2swHDFBWB2fJWYtyWHu8nCtXcx8vDaJqkq/G+dsbZZh2/DO1LKEac/luE
/rfEIAzLalDHXEODPZPzNLkSPQqF0C3eLDfvTUyv1AY7wrTomlFjtms3vzoxBlSO
7H+IgbVIMdieoJ/Ld/aJoZ0Kq/UqCj81hdDhpn7NMPPehtP8t80dDwKb9IHD+KIx
XJ2LfZAOgIanJ1bf4MxMe5xmTJv/+XhmYRLibUbI4e+Vu2loSVusJcI1yn2Biko6
+NUR1y8Bzkd1fgPMtcy1ZksMV9WqYOPrWcCOIzMf89oPXY633T7vpK37nbsF/FYA
ccgA58C2M0FqoBVZVSC4kf+bn30y3cR+iPQGHaWfMHfD5wTC7amtGhhY/MkuHBbc
wQ8NA2A+janlPS0njPtVEw==
`protect END_PROTECTED
