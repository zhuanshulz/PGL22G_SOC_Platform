`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+mDFiJrH8vmkYAIQwzy+voOx0ykCojE8e0pBx8vvsKXiWyspRUwLUqyYjroglC1T
Jhpd7Ca2rVUR7YWCOLODNIZp//Ddfpmvx2pqTgUn89/Cz0bKWJWlAClc1X9hXqdz
mAyu/nYZy6i+9R9QuZFbwPHaJQ1tWEwh26dgXdp6FCYJgVO6+hZy3nUPznZC/SXV
32/f3ER0dMkoYc6X7+2ANANknrBZN69nDHKokD0NOj4T9jkeNllhxpli0GS3Af0D
K3Kc8tuBT6EPX6hpyvfZqmDIhTCd2h8GE+4m8jy4zV4SNbppO+BOA6Ucd++PYlrR
LAA1DRdUYZKYOyHXuhZfDNAUxajVwZL48IaMKMxms6WuJDzmNFKcTxq8wWDb8/vU
Ld824A5LjT90x53njFYJBt8CSbHaC89hTr5n5BvoJ/VN2xIN0pQ/NMPsXbN8ucTh
UBuDt3kPjpO+H8zEFiGc3lMBzN4/KJ7laucFIjVtfElyHou1iNHGQGNJB/ZIsVt4
EWcwCuBMzowxhRlmIAApXLHYkYDez5pCOqnep+KZWCxrrFOxcFCe3dszrllQeU00
3Yw1azoqayjFZuq4MvZpvfnVd7bblYD7ptZ2dRhrSnqMoRicZeRZrnaSnFEM5pHp
l6p5IDQQS2871syuRTH4KF7oTNgVkS2nffUvxldv9SupJgB84nkQPilFfpBgdULw
BIt2qLegdYWiFJQWGMZ4cQ6m5vjgEHsyEqkExNX1O/ln5iQyCBwQmIfbpMmw5T8W
YHm23xMHcMGiSuY9rqIelnbok5x3FdTKy8FFAO0obaaSQ7E98cyr2ZjsdBw75Xai
`protect END_PROTECTED
