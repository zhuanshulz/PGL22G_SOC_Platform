`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VXZj89fIkOzxWxyD+FUsHEtVOkoRScGehYoTFHLZMwrott8i6NG6g5ENQPi4eQ9H
dM/15eM+nIZhJSrhOatHryUpFyT3ynVn2LA1r12or2BlKzpdor1sWUqH1KKryk3r
eRvc2TOndKOlH4jsp/27gfjDQeUj9/fqHzhWfqTEYNBnTzVBYFNZQrU7G0BD0Jzd
repODxD7xYl1v7gsn67qEXqsAX1r9QodwTQgrQo2n6PWiAq46hw59x8++zj17i5X
vaogIZjuVqWhRflALBpN6dxghUpHXaKpETgU5mN1c8DKC25YCHE6G6e6MIIyPHjB
RJECG+BsvKNvNbzeeIQV5R3WyYKhTNuekN3sS0lM9VE98zC4gWwiIEtGmE/WhiOQ
ARh3RASqz2L9S2d0q5Lfewhso/KQzkCUZkAASwFJsmdMtWZOcp70NAcaxeIRFuH5
XUvnAQAuZErECBTxqDW2FbkTisA73Myjo3n6zC/XdPKxbUod+ZqOk3Jq/BQAwrcR
zN39NWKbgtWY9rVx2SUrbO2/QPMMFZnoicxQcjUaTKTm+vnY9KuPk8DAxeMCjTxL
v7GFaxoVLnc1Efsc6M9qy+WLAfwTfdwnQ1Rkxqg9ASJreHOy3p7C2JbWdp++vFgi
qZgVPgYC0z9qrBifEOxBURUlYiLqe3oKIk+TJn1U622+Ew+8u7j3CyvZguajyZPi
ztOTDFqQOzSdAxqNpUralNy9fFrCACm16kSnV78pj3QK49x5CmDVfbgFf/ukGv3a
GyBUbrRoC9s9e0LZit8dxT0LM/a+/wohyQzb95gVWBvbME0Av8g1CiCWPaUTvP++
Qyx2j8NLNH24rceoql9sbLj9Il+ZBNVWTH8XvvpZ6H/NlYDIppRL8Qv3LkWS0+vB
zWzBEskr0fjyYgahHv6ACAVKMlgtTF24duAso6bys6GOVJP+MKMokv+E90IPG1lY
ZIHIELesk8GMf9wdOBAkhmz3tG1tErsbbxpIMmLbFJcBrN+Ztko4TaHMfJDEC5If
nhqy9J3iIDz+CHb8fyRyxO5i5yA4XG8wyn+02KEGeZvlRmbPXOqEyws+vv3Ry4bO
POQCws2Dmg6ssbKxy9O/u5NCdwEcoA5phUCUwrlNmepB86/CW1PeCH8/UMNjUteG
mTAKfTicGqYx+zHkb2q4SVLEFc2imQf8DRr6hSOFIDsMhCAtB6yVcer5cHCCiK6x
IIRO0f0qwUMt3ooZtr4H9Srnxuey0MoT68m9VGCN6QIIRld2MoTfJ5d7MpcWBVmV
8PA1GdLPmJ2GVscWoVpsmIN2BCAcns2nIoyJN0nAFxCp3A/8ENSh02KdFCZ4wjcZ
4gdK+G2o1DlH8c5ihaoB2Kjtw90Jnvlo/bZlz8+F78E=
`protect END_PROTECTED
