`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L41sIChhriDHHRI2z3ndHUYjK2VqO0a2SOFLUeMfpfzkaZlJCSTu+RnyXJXXfhBW
xy5xCsmxQ76ekqUqQ8A9T229K2wXee4N8VDOwJfb1iE36gIwazQymHkUwx/RatNL
AZ5XpHo1zALLF/ZGSPFocoshqi3NMBNurzFhG3HGlS+LBrvH9PYxIdynCVinRW9e
ryCR6Uadkt6RoX7LFFPKKN4EOBkXIBe3LZ6K57QIExLS4D+uySnq+rtuLIG/eoW8
nz9H+04LpMka7BVcKzYJ6/u05zoGUEwnDqdTAXrvhAP0sJ+TbVDLDMpTsAmW6EME
ir6eXHICOyUtgPqAKmXq1NJ0FccLWjgUu4OFgcBZx0uQvapbgeu6fyYE6uCZgqRP
epKNxkqRPtLoVmcsJV9uP0lu9dkIiQORW7YOeCju8gsuCk8AEfIy480cGdL/CWD2
Bq8r2TFlcpqPyEflLuLYBj7cICrV4Tt7jPiGO23DF3+Oxyxm+zwPre6uY5eXnZmo
gJ8fRkC0qPaAHlF/zas1k1osKSgBLl8ktT69Ts+NRp0Vx3CfNwbsjUTYGAapnRNQ
x9ch3vlThrtNiln80RID9A==
`protect END_PROTECTED
