`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4qOSJ3wDnYyq+FxXpnQVHaN5XRqoZa5hKWVunsLfV8ERms0SaruS4arwekIJ+K2X
3aspCyo+DCGVsiTSVXQrN9kakk0rX7R6OjIl2HNLislnEUuy0RstQD54c9cmp9uZ
iN5KFO7zOVVQLz0jh+MgXMO1OeaM0sPkcX+Xfoeql+wSIPA3TpSeaWBTFvX5UIZX
tj9w50m2tIWYZf/0ujZHBWf6gToMKlF5Yz5dWoEgMl9aPPR7aoGClPxHNF+X61jr
Ek2JCH+HvP0W3L/BPQixgmL9eXgrHS/LVSC7s+fnrg+EByNNukVGb7dERQ+ju7ia
KOw99EP+08S/Mh9+G2ElZhgXI3kP8PvgLsPBHFk8RbQU7ca6hD1qchCmPM9365PJ
i8sQ9ls6Fv6374gjOxxnVfHdQisqabZy2sm49tNuk+2+V5tfHwWFLSUkluLw1KUn
zalOSQ79aMNX+vgwuBkYXVajYcdY4otC/YWB8MN80F7xRodtHgmazGB8hyZvUBwj
XdE2qSyxvFLDKFf8nP2mJx/LujOrEusNc5ZW4dULzrs0DM+3R+NUaZOehXKRSsZc
0j7BOxfx1FkWI8nGMe1V8DUHsss1KSORxtwpLs04Hvlxiy1IQyEmut3C7Hik5Ivg
zSWRcvEu50lW6Pjfv1lwL5TA0wGZ3Oi9chVExR7NnFpt2QayGxF6r4Dap/wPD5Ze
G+sqSmbec3LXIoKQqeUJDmhLC7tQZsnnc3yINUafv4D9cdsbl+iYFFirI1kpDocr
aMSbmALW3TLZV9vgdMenXBZN19xpkPgC3PHgxyjjBPYJQhfIG0WlL8HU3xblQXsX
WTZQcPg4mlAM2Pn1pan0pMcKjsemBMedcHn1EH2KCEGe2BT/wtNoHUmdn7Bfh7Qf
P/uDoN+RPFp3kSkTGRjs9S4zLo88zZSuuYGly1rBOJPpuDw+6YQUsTGyquN9TBLD
Td2/v95RNQyI3uoqktgsGda1jaBf6eymMv5zC8Y3VNzNMSzhGwfXbz93/0Ddo7bI
tVWSfF50WR7wlq0TKTPtaA/+6TzlWdV82OzLEtWu6h0Vl3fcrN3uzES/Wa3HZW1f
tUz6Gwn6bxMorBwPdErJou1t0BiLqnfzPerG1jwjlvDhGp0H9rGKBc+N7egsl5b9
GiyfbUqubtBZvBgoP4jEQPmadFJxXBrUn+OlykkLKoYtG/ERLZpiWUYj9YbM12hn
G60iVvgrt8ilWhAy1zZiRmw2kvlhUFYEhFv+ZyGRakwZY/M9a0Kc8nKNxBWguOQ1
RuWhswONYf5zR2QlborJp3KP4G7Gn1peXw4q0ZqpOBh65RJALfwuOwWsUo5DANYb
Jjc5NjAmBun2egemVrfoKcpd7Eo8vqw1PVW2xeiX6+t98se+u/0sseDbD8OLctaq
GKm7O4YuvL07RX0b/WjHqYvAEI8Y/Hg38cgq4/bupK1G8mV6BNQRLGg//G4F5fPK
ifMiBMH9JET+puQm9QWi0bmppdDOGcy/COow7sw6lu3PkIlCMiINlEY2ykp8Z0Q8
eBcYOHTJxXAjkBrHEzVuUri7j+afklGv4KKy7OU5e6mX9vNmCRUPu6bsCs2qUMg6
iHGU+pFPZ+XDTLMIJeTwcv+4GgEbLpSr+81MmL2VmbVSy/FPiUSc/unyhBENZMwI
pDte2pFmkwN9rtv4EepZKlc0pByDB5FVPPfiE2YbeBv8iqeKS8KQzyZrZ8vJyLqO
wwp5xy4abDrtfjfeiCTI6jB8IQuuKYiktOMiflBqS/LhJZGUaIDEHmWAh+gie/ir
tS2nTSbI0wKDLnWfeVcgPNNrOdO2dHmmnhdxmyTQc0y/lejReBjShhodZ9GK6XB1
MAXSAvYDS3GXHrOFGI0Ohp0JpPMrua3HS8/fMW1yonndrmh8UtVsdLCJkfLunkyn
kEKAc9RoCWsns+0dPU75xzpXnLNmrMm11vsPoPv+ZsKrl5rUdB0yQKPEvqCAu6NW
Ypk5keSRN+7geX3rWYmK6IhNbkBWg+gwTahCyBSoX/Eglv2oIbkmfdYalg77cfhI
QhlxrtuLfb80S57oXWD8EE2TTQVCHPqbZlyO3jafySoXduVr3loZSbDlfEJ4/P3h
uIWPyQ2qLWHpEiQN2RnQkMtjUdM3CEV4DEv3nVeuNgFlF1ymrIIJY7uCHviAdNvu
U36RRXExqckG7vLz1ENN59FnMOcYABoGohteUMksMhIRvUQFR6GqcFDBrmPz9ICA
1guXuWKVmvwSa7NVFEngPI64IYg2J3sZgxNUvmYU/WFVu80uMWR2+tg28/8IsQQ4
9WPBoosCkWz0sg62OQ69ghHUHBhPMPIP0cNSo5P3JQsI4E0eRsQHl0zlhq1m6r+e
EQd0WFIEwHbWJw5Danm/vx8hEGf5xhyMroemKNO0FKqgIKEdOv8kqSo99z7Sd2D5
FX5d9f+NMUsQo9UScSK/dcCdn8Tm0dyuCmFIf4EAbDWV92Cml0OBQ7QNKmsd+SSq
fF6tKizliJwAXYNvOeUUqnSLox7ZxDWJhFIRoeE4HrcsvuiYWAlh87L7M5jVhTBo
FUiidev3XT10ICA3ZpVOuO6e2LhaOQqaYdbs4U4LKGhekflI7Gg8xVNp/W6o+RRd
vzIwA1o/wekZz1SYbpzNNpNcuMdhCeU5OCE9ZQ94FYvkyKtZzxRmOwWy6U9TCX9p
D+qIwc4awolDXZgjV22tqc+Jm92myJLsjh23bjNDMoo6i8tcQ+PE7t3D9L1zUkyO
dti+BlY5+7WQjPMS/NKzJZEI8KQglnv93BRxowAvY8smvzy/K6hyMyxylO806Ofp
965PED9sBR6vSenhLGFo4ws5C1Bj6sWdEkyjCv2QCmKf/KePebtMaHEbKlJdb0th
H4Vtjh4CngUO9ZZBIT9KdQC3lAQPDQODaX5bWXJWmGVoYDK0Ju0rAQuxe8Uz2eNq
0HNGsCGF4DVQq3IeqFtrft+cgEE+6XMa98eA3lQZmoQ5dKDXPm60fLpaX3AzDW9s
K2+54lhDrKuC4SRMGXaOQNQlPKuZjM9gmh6VaNbYaPWIyOU/BeKKb6l0/wjQSJyx
8mOCRNmqtRXRyNkPmoZdn0rpjLtHROsuvcGplFCQHfVS6RIHMTWvZLnLsUt4qZ76
ssvb4DyxDX9dEU0qizhBmbfr9r+60cwGT0C9uH1UGVyGMnmN0fL6/qszWCjF8BVo
wRP78APu+xxpc668vdVWVx1AEdckvYi9D9PVE1RawwFUpASvPT/7m1TMpZnRuK5R
1JnoAtad8hHD+2gQdPcfvJNzScJcgNX5672F9G+u5HfYtUhwSQOP24+oVNAgS/7F
FW80cklVpDUj2JDojJc2mV2J/DvpQ0ZAfqrv6hvFAGoo13dshb1kB5A332EGodIo
SpX7aEcnlNCXgdErHnWi9K2imyjDvE1Np4/DvsT2QCqCrGBeavnbmtPk3h5s8tDz
AveU6yabrxvpgvlGM1LfcPEpOCPfFHqIqJ/ZYaz+TMAbqJ+99eCrVAaqBf1slUf5
MZGIJg3mAWXBSFtgFhR7OSBIoCAOzqYkuB733kM/7rx+6T5F425XR8vg8/tswGA0
m27+QX/DERtm3v4fQpk4AHq9qH6wSbpOJVf23FUAqoOJq6tS6tXBeXuI6LcgNGjJ
t9m53MdO5jNaKBeRAqtJhgtssJmx8RA6VhN165Z3XzZk8gBcMaWi2whfhrux2ABX
swD0WI+QN8m31rHaSB5gjis2Cvb7PtUN3loXZ+53pCiVW1HpcJaOioJhTn6dRYU4
vMYh8dsLZR7XE52T7sHzKNEANpK+I79Svrizly4hNCprxopUJtAqxCaqi8EJ0k3L
OCnJJEVN/0uf6W71uLwqALPZc3PR9H/EFCmNfj2UZ7ji1nMKsZVW9AMubnHSX981
WaTUq2KgqTCXBVwIDlkZiiHOAXhv8Grw4Riq2niRoulgvH+bKASeGmrnuJdd5ZDq
PgMRm3j5o+Z4smux21qh9Fu2H7y+31vwZu/rv4fk9VtxMDwQOwipt4NbgpUa9v8N
gPMBulG3mrMDY2vhNDRXLcBSQAIeU+FFqmo0GLGtz+2EZgT4x093ygJCrE5chMnb
3/Mu5OHrgvmKIJryyT2dYOoZF4RVpiowsUfBoA45JMhBFtaDRjbUA/3/2sysoHJn
nUel1NIDmaCAMoaINJRInFaYsTb13F6xETOXRB2tKUcjCXUJEQpI+EQtGNhEHiU4
+GqTWkQLgID50WzkuBCnqEmRpmLzsGgFkCB9HcBi/qhkmlSHpt0Y9amEYyFT8fIK
0kegoIexcbknn0SyEquF6/xRjkL3P8I1bPlCFdnSZdf+tAZdNF4DSUZGke7NOof0
l6ZOiLqDRWoQ1kjHp2jNruocLgSRSaCHmbESqOIGN8le8ckIcUcePSw+4ETrXyDC
ccZl7WZyjpNfyaKvtoQQJWCInTxVeTyW2EKQynyM0QgP0NI3DYmTLwFfLYYshx8R
6tOqpYBJTDfDU3W8wttxxjF0V/GB4bRG6yKmn3ne3JJCmR0TOxDIOo8pzxugETNU
2kxrCN8QW4JM2zvr4EwGe9QcBapdApXF4StBAAdmBwLdbBoeTKn4kpDFbRkXbWPy
elAuRpy9uCX7O1/xg2SUmsWzYfPKKbH6+8y3LCUI7ap9NEjfEZM97ytSJY8wGuEb
CUkKKxHTP2PyPoVmpgGtRMTUbsWFY/gqic4Z17daUfIljy2n3VxL5WIRbgLqHhDB
V+lRXyqARSkpZYZ+BnSYQ5UJUIXIOJrfRyR0rVlP8nnSZD3vO1oNbboSedyo4HXd
e+tVeYbjp+PiYBzOhj/A/BnZwJ/9ajcG+kgGDjkilJ3CK+VANCVMHlVYhg0vjLNj
lvPohhxQFyu7jXCYDXJLrYtqUzzMiI/L4KR2nEIWrxMDXFkUHTIndm1CjmdqPkti
cC5TI26sb3GC4mK7UOT1EdlHKarkmIRZdbZzHgEHtQGMKXfxSZkqERRydagvNRH7
KPeHA+ClG7L7X77YPW/QkxM3dyJ9Bo3g12JD3pvFibD/X8onxtwMTUl62rn74zBO
mpYAZcdldJl6mUx04vQpvnqDyPzcavBxOzRtdCTtm24vVvBMBOoNVfKQACR5sTio
wXkq4/gpvb+jpWib5BP50IlEpXRd4lmj7fYbQRdD3liaAthRB1JLVT7e7ixbIQsu
zlnF8ClsA89/zC4jh1N7Q/PLbOi4JYdrq7tDKOO6p4RI7GSqd9Qrd4QutlA5P4I4
ybiwwdP6E1PrDQWvFdEPlj91QO+qjtGdpdiJLVzUK+0K/sl46ydELd3+MmLGwPO/
Ze5ZBh25u4yJIqPInoC8IrMgHEnIjE75l/HAX6Nr2682R9SaXRhavMBSOEPKFUUY
fQgBdNB6Z8GE6PDxyUwJPZ9fLI9MDptUHXHg6z5+jvGCtCewHnDu9vPieQrq1P7I
Tydl/j1pwFcRlEk3ooiBsnEh4mnuZ+ojz91+JlK7zD6mgR0GKRV/Gtl7D50hB4lz
heBBmFZUbMCEXdAvr42ekXHBQJLjWlesiWq89cWQMifYBH5BZycG2zMITt5MJCVh
KC3biV7eKpJijnUHUOf/rDbvuiRZJg9Cz4fat9DVo0qgwRBBeVaY23Ai3C+4L86o
XnwRPs5N1a/HSt1P4QREkgnVjc2CSICxjRX/DLlHetQGvp18O++Pil7sc0IdrBlB
WT2zCm7FAu3WJOICsQNhJK1mlJToUO78OJFlyFTv+bqFzju2TWTEIBFLVjarn5aH
7zWB7DaWnHr02mFQJzwIKCkoLvTH8YgV5l0xcgXR6dO+UZX7cmH5JLjqB8h3qRXH
AMRC1cDTnSQjzTKDSCIen6BU9tCo7Pjm+a0u7RduCNIrEHrHNEUznRW/Vj5VgXHn
523UAkp9VG1VLY/GuH0St0qK7sB6T9t7u0sz5zhJg9OMeAy0cPW1hxXRmIHB7OwB
xTYtzLApJ1/xrWnpNUIaKkp4oYyfTh2NTxOEXonDizWh/vOOu1m/gRYc8deTJwxD
zDlVQ+yEIjRM6C8FqNApLocmITm/NGi89xlWM5FP7lYtE5tRU/bvDbxaNMcW7qA+
d+UJ8wWkdjfW1KIYhpWfrqfD22i8BveDLuogAjWsBDjfcgim8AeCOAAT5xNXN5u4
vEdok2BR+1mcxSoSBUOGpu9HKTjFLmbQsdSzPxvS70/A7oodfWLhEBhfWCEjnw0U
RvAJzz3kg3Em3H14m7lqpWxHhmOe6CNxrr3mNJb0fGO0VvxVMfEfmdeZVP9+9J84
+LdiYU8vXLRsyD8B14k3Mc4pJrNnb+0P1N5XANGJyctJbUSRuc749zXzjOtrOQ7D
mpVw4j6rm+r97rFcwYHnxsQCZxNg9RHNM2JF4aLkKXIbjCWn269+1qPCYDCzOVX7
qCgfDUsdjm+g9cBPOTah+f227BeJ83eXENSJZLXHqgumYJ9PhogOCtkeZpiyuSfO
wey9UQmXPDEFIPw68KHV1BWvtHJyu1d3CVfNxkZmAS+4wSerjEF8ehm290dOX1hk
OhYJ7ezkVfdwM6Sl+GJAT5Ms2zIKqtOLKzn8SDgHiE2BUHmxrXGBRBXET28pQdLI
PwLVezHExi/VLPXiRkGsjKp1l56uBRX0RptQ5JWL5EcZMxqfMakB8ImeZhUhE1w0
AnNABb9D/5/9vPYPTEXgNyFA4li5dq0SeATRcnIQmT6y9qLXIqi2mD/mapMHnWWc
QsYmRef/x6Ny8KLKGy/QwfMzBCrYRPN07VqgxCkwQE20zM22AqsbtzNTHiKJPq/+
Fp3WFJyiqe4DM5+jP0dHC15Ucs4eS7uQHDnT5Z+RBFd0FpCg/Phlg6Hyq9JOAkIt
tOra82I1C0MAwakOPKda4z3tGobNZBuVi+qNglloTF5lX18/YVnKsJ94RNK2wPM1
gUpub6LlBjByq8+FeneFnJkGu951MDSq+fGy+cND1N6SAxk6VNsFAHEApxqkJcRT
0tw3RGJKKweocEXXDSh3EbmtTS9URVOu+C8BrWlM+AxCinH3z1vWF71uQRulpMS4
zsorzanFnz9suHiRTcxnpa4UjTHUIFH1npouZ6IzEQuN8uWVkY63OgO5t590ttpr
MA3ZBWBBhnWnOE8p6B6uzJFH5yMVu7ioj46FE02/Dg5fpo+qH7wmhmzk0Ol90X0O
d+56HqouIzh94MILMsykNu57Rbuajpalg/qt6zddf7q1ykVLijTk4NTdglF4pWuu
vNQn7TmD6s9n2DKX/NP9MIWCrbom5VhG6hasYtzzRVzEutp6Ekd7iupoJz8byoX0
SX2ybRcrM7L52Zkz3e8zPYMW++mu0nyx3g7mxD44iyXMO1k+FNJlfnwcsnZ81jYe
QiywLCvhi1mAreeNxYG6rCvRtLTrIoxanQWylFA7qfYqT1oSxeBcpExb9548q7Qo
HtAqmPQkpBqOW4bFfGG1pxQqA6DiZ4zO/1t/qDxsve+IbD3xf8WiD5BB13vVOVi3
xr0dv3jhYPLeUaGZvoKg7OhRnn47t91HJglodokoXJdadWn+FCkxEJ1WYDNIc8Fv
c4wUEecNYR66K/BYh/f043hb7ObKZcP/V17m11XAIBsh2rH2/OgaTwmLLlC9N01v
jo6STg7+OhpGwFBDhgq2cp404kdYcVUcIJmaxwuPj99fJjT4unXkdozuVEo7kdpd
334yGrF+odUsOPGwS1kr80gpoQU7ZWSgv04DxxEphLFeX0aENL1YQmfHFEcw/ri/
RQ84yFPuGZ1jCGtvXOogytIj2QpVjgq8+8VRmEs7vFo8XW85eFnbPvwGJj4OEoys
R9uYfT2O8EEBoBNcRjaPqMv/6sEAcBy2YSVYvQPwoY8NNvWbhqz5ScOt5JdyLyn9
9suBaaWLajOgnaDQ9k6O8Mvtaw3eBVV1xQHKCNfRhlQrdEAh0UrVe2YBp/ro/vub
9eStREq2A/11h4JdZBMiEyJSqugyBXgF6uEJnyCLC3hhDDRf+SQXRIzT/hQCv+0C
P7L+KQlgbV3+0g8lHjDKlcYXxmKatn+hvylNLcKZlVeS9m7V2RoPps/eIyemQ8De
mwu9/1PoQH8AhnDk8XAH91ETfGTd2Y20hYB30VlbMg06irJpDTJC1OSNv5TZw5np
N83OMosG9hCvcHw0JUHrnzTMe+vgmtC8Vp4OuDiOvC7KCTLL7SP1wDNM3gWFVeqd
8egIl202ZHFKkCDsZYzSMTb0p8HurBLIbTuihowOguskLJcomHJDq9AXmSm5omWe
qsq/XPIjBu/sYB4cXzRa2atsZixnl3Pb/y8Vml4PfaBEhVnApzFKs3opz1veHePq
uJMciVyGnuNaUYhSeQcs2SeHOLWqyN8WM6/RfEN1VXg9FmgNnpNIPSx0AbEaEgaD
of5RqGAUso1gkDpTictUEzgqp/jEzJb6u5jc1FROT2WKK211CWtetgiTfeA9iqkS
vde/6VpBmoqcObLArNPHL1w4ysy+pcFxzuwYTFFfPqoIbNfO89Gok6jSCLEMIJ6g
5A4VuMDhgwDkn7Iu5+2qX8Zd/BASIl4b0+mm6t1ORqmfxSGft2D0i3r/v0PA0Z6p
6SXwHXLjRJj3fale0N3JXVLqd68/teaA2qFMYd6qn/+jG2yk9KwF0gtJoNXQ20x1
0j+GxDO3CYDDBESm8fCGzyuvb68/kSCn6KXfVXhBAf97Ibq1WN+NzWB4Wbum3QuM
ymp1VCOloFzqRel5PWY9TOBzmivG711kEtmAYaWD/kQieHIbDz/Dc8ahKmVqOoyw
icocnUFbJjWEigHS+mUuLDyPvqWmA6/dJH4shIvtd1d6aRTHeaYainNGe11XQQmi
Tf25mKZ879nBDqRMQBfRZS/RiIE1/lKruSbMcs+64TJtAjvS0yGpHRmbMfp4zPl3
Ia5tvR7j6NOj6BDaRQBPYU4xGVShUUAV+YQx8KC9TnhmQQT5JGujY1SIuxzpjNrY
ikA55qZWylFD7ag9/zyDyVx1OcZN8ltufZKsO4SRTiemGaA/Q4h4NbLX61ib2qKU
niaimv2yuhGVbCsIIm+K72qTQBfKLU1Egs7LEdAGiHRrqdHrjLq9SS+BfY40ylRG
f4FgwqO69dRw7FYPiO3mYdDTR27AQFqWHyNYjGBQ5pPNhZjjKs6QeQrEfmBTnNA/
28CqwJWuKCBBPgQ50Gu30RCBRnOhMse7L3WqjwCzc9wAe24VgW3uTUSZbVrtD4/A
wtcAHw5XyiLPrfCiOTw1p/fOZUVYs1COaW6aySY3kF+gi75w55pJM/37TaD5qjtB
2cvd+tsHX7nds9mRdiBndPkckruLWPxzWE46zQ3AJV4y8iE6lFlgOws0R6KCc9uO
X0ZoF/DQkR+fqTSG67RfD0Ht/p5wZkAU2QUUmiwckEsNSXoqJFJPF3x8Xx5H7flH
Kwv9lvuWSlUqPTPuDlL8BiCsWA7MFCI4xNiAUCtKXbUteAbmWAp9IDU0SjH+imC1
ptwNw6Puv99b0t3wKwNeWuoygxI61TALRSAUJwJ7BnNxXYJS0pbrgMLAkGsruFrI
GFwA8y5afOcFmxhnldtl8nAdVpUe71QZ7wpmIt/r8CRUsqecDxIkQ4uknxOKKpcU
QXNWY51/24U7WDijASwH9x+bTyCyvHkzMXGxuKG9cD/retYCSP7eamG5VCWXo3UI
GT/dM+mYd24XBVGYHu5EYwcoVjBoWoNIV07LgGgCiQlK1LESRsd7Z+YGrzafD0lV
efQHVxWpQwCGqKP6t5f8G9OTdvohLItQWdinyWDQ0ZZA6dtEWRyVezl4EVRFmSDJ
vCzRDFUVLw/DyEmkvcqRKT1YXacoVoc6Az2m4ip8T8XCGA+gLgQQ7ymL+j3uSTkP
lBsC8SicyQyaOFMJxN8hyPoKH1kyTCeXqyX1hN8/ilRI1pM/+uD9sIyc0jjHBPe/
O7tR3IsYEhL5tXb2GHz4UX9vQEyjz1FA2VG7XCh4KpAQowkX8YV5mCDWsFaWYUt1
+m3Kxvy2L266BFw2ZyKsxnX0d6Qc6V7jacstoUPg2486DX6h6c9ra16Kx+BLZIHy
jzCoQladcmBB2qtpuSHvmT2QQOajsRAn/Dy5LR/1jQtHP++t6d1SyzIo0M5lj7Lr
5uGpkNUsBWouqIHSfPo8cJrYi9UEiCadZRQRMF+84J8E+g7+zdUYHxwd8u6+fTzT
LVsc60ZMaPl3ZngO4CxaJn+gYFtV4p4owR6KplEE/1msy0HwPLcWJ62tJ8jqTo7W
kBqJrRRWLDsGdmzfBnloMDXdun0sc/1g/hs+vpAa5DdeYMWTjSmJv2qDPDkBFs/n
jQqLrNZ1LUyJYlJ6xdkyBxV8zyOM1bygfitW/7kpSS6dPzTcMrHB/cvwgDNpIISp
rLti02RgRb4AvmRh1C8C3vVU6pHTvwYj0YkTH7AOo4CIVR+6D/Glz7qmU7ucSSMJ
KBZAItGRKHX6mvwL01yCCCEYUx89zffl57GteFeVEPYzat7dobRa1XpcqFTOiKZ4
2LJ7kpo5ZLNtGm+DwWc4Fte7tFNLMcrv6RgYvacSW8PAazj7lb5vd1DFRLVNDp/1
bUoFblEVFs9o+4MpzrO4OfGwBjCuj410wu05FCBTiQWfdM5kcACPABjrGt02TM7z
MxPhVi5/aweec0htXyfivZxw2KMbfWGNd8SXMWCrF2W4sAY5qSXGcb6+hcofaSxr
icNzbbbKNLRTFyenKGUsJVwgauA9DkSF94bIVLMkt4I3yKM3Su6o53lT550Cuks0
5IUoTNtRm+Itlw0Kwzx128l8zc/wCdjbxDU3Z/qP13YQCGSVZykhj/jfy04sKUGb
pvYXYeMnJzGgfwGcgVvbI4zMTejMREiGRqSEDxrnHncNecwfquTjaWcdEpGYow4z
DbWaJMQenBScuipdR/916uepFBsLXQ/k414HjGn+WLlVvasnX0I4PJPQ+9D9GJ38
cOYRBsKh19XJPDrYsFhIg1hM56Amf5VH0sY8wzSJmg0+MsVgaY+QhJfz37uGv9Vq
0XLgaa87Mo4+k9hlxajN+rUJ6Yh+c4hydOzcoJfo9TXg/i9PRjLJsr2RFxwvz+p8
zEyywSV9+1kyRVppVQBHRyGOYUXy2nkDweqSr56d0tw9zAaJ4e6JP0ZmcTS1q727
SexQ+N2SXhtVYlHy1Z5Lg+v9hObG9O/4wGDVpByx7RPhYA+uBPdoY6kqEvw+WJMl
x1XADRWblYybGRhL4dmMwd81D93P4+8y4eDX47eyXgwo8ij698v7THmOBkUJ9Mo2
dnZ+9qapo5kPQu8ODbgqEBIdh0OJGLj19wMX0xiR3anKLuxLZjAsMrT1t/VK8ew9
XiY1O94n2mj2Cv8Md31HAqU21Do21wSb7L1C+6ZEBB1CVe/FPjFNHJE2JbJhIujg
5KUHS2bk7YDS3TXr4nh/qgj6x26bwfixK1u5sfgigql7mBX4klGMMD7W335hgwur
9znZ6Sm+AieCBW0OHwrJmOiSQ3fhcj7AFbbvH7hZH98Amfkkr0SOIkGPI6SVLUPr
jOTcWsdE6IJoHp23vua5W/Uhgm5gDtD4zcjT6ouYmLr3/Pp3eFuGFPLB1A4zVJ4Y
sQ9AXxl+yQlLQN2m1UFISnaDR7NOci9m239k6H9NWfJsjdWSLakZ8tiA9/28Gxsv
BVxgmm+NiLH2fI6QtJAfJlx3Y95O+dfm9bbB7vTL7GsM1IfbQQkIp2lyMICJe/eZ
z9BUhyjSEKTd6zniWUmMGSRui1z06VhgDnSEtPCuYHdeRTU82ybOEqkZZDAHIytA
/BE0iLMrQUGgN6ekQI0CKIsAyQVHJ0v9WJSX8EVv0GBDuFWlF09Gm+0bUfTZL0+T
9jWy1h2BTkIH3LwPEQifpNpTlSu1LWu8IyYE/SJx9IBXVTkgXcNePY7sLi6Xgswh
DsIGCvIKa6BWbEeGOWVrLDb9gN7DYIy7xXwvTVxPT9uMzq5NXhqElx91LnLIjU/I
kZZVZr9RqmPLhovw/nsy8wLEa3dFSMkvG22PsqtVycSKEPEIQFychSgNp5U8SR4R
RT0ifi8M2CBCxDFhaLR54PxZwjfg/4tNJHIDIP5EfjAEK4zB47OCpL3A+5U5FzEQ
Ac8NcL1VGybcPvr0DtnEgiJd12DK+M73dA/UHyNTSUSLEGXU2r3lJg9OPwBSVQaK
tkRW3whX08d650HoMu6irrSNsCIIpo33wfuv7UcbGHPjeOxsNya/7RUbl4QkU5ln
d07mAr1ihGXTrtJlCGljF/FtBobiGgAYh/RcmDuOsgfIIQ6T7ls2ujNFsXhb5iEE
bCerBMcjAb5rGWkUrrfH53qQTOrMuPGBIicqWlMqc9IWGqxXDuUALLJ+3TJIpEZY
9ifRKqH0UMRF+Q0Wq5rLcva9qTNs0SA+RPGFPuQFFJ3qR2NJibo1N/0jGpgbdm5c
hFguhD/79pG5Qa7RKSp4MUcY/31/zZdPZOStFyhpEMEymI/rdrC68qVHBB/IkjlN
aFmSVBKiJZlymKjkHnhwhnDMNjTNQspSUqYdUPWctB7hxpsDiHm8gfuJRsutQyXG
IeIZmQA2KAdC7atadjvgTvFaflsX0vwruHsrE4y+bs2v6b5EiQER7P3HaNPI5/z3
0f+k7xCw/1hnNpgJYwvpxyubLc1wlgq0jSijzG8wMFGkXWTrEB0kayVFqJDpn83O
357xakJW5I8mamxfu68nr6cnytRLiF9yiHmV9hQ8/yjlrAdFdk/ePpNYNcN2vicb
VgQVG4SOkhePbzCRuxibpxve+ucm2AxfdbgLc7gjbbEycM4FN+xKKZTLMk0lXufM
URUQ5HnJ5WHK8jOgQFgkHiZRCGYUssazeG6TFTrBMGNwFUNFeG1t6j4hPz7R4zZU
7fOiRvh4g8rnvWa8XK+7yxl95/0nzJHYoywVCFcRGLGKKyudK8vCktpULBtUwQZD
FKa/xPfWzCEqGpqDqXWhNTm9SKsjWQf5D+fnFPhbiF55bAsWETlgLYkvXuHcSAgR
SDsH0vqqtt3AwXBvln3eFQmxnZZXn9ME6efPNPSWBTkJ/7DDjtsDEVfNcNhXHgFH
MMuRQ5sLy2vwLYUgW/93vJfk98XQRi0BitEjpRO4vOSDsrGRHZelp5/k6rLzbvbW
UMsy8BGR+duOXGtcCFafFYUZcqgfQBzBXoBFNJaN1VjmJaeKKtgPIBbcPiMkOmtl
ijP22lUTDbKzjt3jf0ghSLs+B9gNJmKQnyVKjN4TgQ2ArpCmfEeJ13Fp1I5JYZJ0
0U7bahIWwpaogCSzwo2HfTMBs6Orgd1PglfV2AVFI4dMrpxHnD6woQsei9aYMHMa
lzKS557p/gMQrdTKcPJesIp4lPTSUlaHVsKLRhfkbFNWP7PScszb4Jl4NeNh0nst
pqgRqKGcJHLC7J5cSbfIJ9atZLq66X/+e8Ny4EWKtF6x3q58hSAbiWW6uUxQ9Tuk
kNhibk8Bi/e/7ZXgLB31TxMxzAijW4wtLOR9VOLP/72xriEoz3Dm64mLyivcewE4
PRCiMG0nYFvYyvr1XjyVo4oQIEoalyhIce0cUmf4QJfi2rSULvfSz7eZPoGXbKEP
OIDTgNFsTHsW2IbeUtYL7kH0AW/JGPUv235iY4Km2nCWm0lrRvlnd8pHY8lPceiT
3Ko/QzBe56O7DdaUqd3G/qSckVdycZPyvHaiy4gXV/8ClSgiND0QP54NcuJkwbAE
QRsSKOaWdEFY9tklt/DtoeMY0eFgJo70Kve9MlObXW/h988qWWHYe4kY9grAqP3P
bZZrOPcLPYSQyGJHRuES3paTRBrcdB8PWVWv7YJmHB7oxQGVFpN9oDmXWDHP88QY
cMTD/Co2sfs1yK5/FQ/eDBKj9YiE2Pj0UBTkSZjNtwjYzRU6aN309Dc0pF3q6NiK
zlW409of1xpSac4pA8E0rgsIoiclaDmkL9kF95uHTz+RSxhHl6ppTdltjy/uMjrF
PnZ0kEbxXct/gq+FKP+20ZSONuv6bvd0+gjtRuOpLOQ/7nFBAq8Zn3jzCDkGyKky
KYFzYflZUPeMsX5TYylnU/HeMLI+WWyjuPbPdIn9c9G37YEbkL5mM6CV58hTrKwS
PgRIxsnsDdasA57G6GVwrk2mFiPP3ZDObx+r5b6WHzEwrlhUHx5tH1/GAqEEMBPy
HVOgmaLr7s1InbNk37YtIv5Iifq31GvCAQKQ4tLxL7KQW2AV8S7wVETY9AtDXJhU
QQSrYgINg9DErD7lVO6OqVB2GZQFpqJc0NGkUfehMB0iSmxBrFQIxTwArSTK4GKq
X/ON8lW6urq+/YeouxNZ+XQYbmUpyc0/DJpk3JTE4Xwb8iFpNDmvLnH/1k4iLMLf
W8s4vwVbl/zPZGtiTR2LyeISw7KQtX1Pv7Bnygf/ITGi1HZgCBlJVsLhcbYjE7ze
SkJMmo3kswe5kDUPJiNjwx5FwAtBPHX2FS3d9ndhJxEhxkxo2h0/3IZxtz6wAukh
7Sf7bSKOH/5AytVmRAzf45es9XO2nzRln3PBbTP2zINkfca2I2BOx89+ZMLGVCOT
PZAAOch/MSCyblWIVpNEgAPp/fpUpIOZ08S19znVfFZ4ez4UxROnO0P0qPbLXAjZ
Set6y/JyWaxhTa+NRjQzibHsreZDdHiaSPiYKRkTYqvIrM9DVjfMkhpSmBwRCoEO
ff4ANUDYRBUhYXAXbaLXx7Uqe1a6O6J1Jp2ORoxpoOomt45wkaVGui2E/jxRrPTD
fe/g1w46b89U2LCwWEHa9aQnlFXfDHbAhMdBgviYdjZN6nHIQpUtsDC/uiPMQPqa
8IhKCBRsAk4lOxPkWPFbA/GZumxWHLiWamPzvWFZ6zCUWWS+e16PGgC/jWpNanQw
9CmK1th8eDCOWOmdKYaO7+9y2S6iFICIs6WyenrNKVVc1kZd7zec3MBsKBwuza/u
s00vUaE5slJYWJ21Z63NxghE4HfOPl7wyqLMJl4HeV/zNOkSsJuUwnavR9myg4bw
Q2BmkXZiVle7FDgjrMfWj4RfiuxpxGKOplXlFv0F+jSvnX084qElKSoIpgwxpfEL
qNReStE8i1JBNiNBiRmuIvFc3IxFxIiRpEEpwIVL0gucdx0cTXPRXQ5i+k77D31n
SmbyS4+Vcl1AP9EfoxXkHV1/zSQ9oIXfY1/rqkXYClRpYB//PZ6gWgVIh8gscvy4
0pKXY0BV4CLKZlNQxEGyZRvmZ8TOxMPOGVMyoAvMGaLFz3ZF9VgRD6mJApvYEKOf
sTmpD178SS9oi/8TKXfcCvAjp1MAUbTSDpdBpPImHC7v06S44tAljCHIsi9ttnUR
r77H39zdvve2zaCFnUOGYYIpArzxaUS3PojeGyECfWtVj7QeHAI88EcZEwVEj5BI
/YX3K79e+WdQykCU7ICVBUV4O7DqRuJ9j1Ls2xG/T1nVASfNF6SCQRfCencJkraQ
ZtnpZA5LuqXNf11uUkcX0iXpV8ZGtskGdjm41omVWuhXdEiBLHvK8Ajoim6kAXHU
HhX4y5wI7pAj2fLG13LXhci0jnsHlde44JJlSR6rFWXXP/igjEIjaNiLs5RgjrJJ
Eb0gx5PRfigQkfDUilbQjgNZIIhToqjPowdXEj4SaFGjH/Cs9OIUmoNbLiTLtVE/
4y4aYOVljJZTwRZE6uisUfQmEOXl83nvM+7K/iLTURC0nMIniL9qe4JpUwXAnLEE
sXg6wisiSdpEqAZJSR1wiR4H2KI6uTDgTajfgbvztxFJ+p943iR44TNDQMDXvp3V
cvbOxqo6KSCKm2WKpynom2iS2kguXl8EhIttXTg02Yfpdz5/mX9K+ozaIX0Gr9v7
Qdlg+pzhlYRPh9+2AZK/IdIFcld1NBfZp0mbTng+sYuJVMhgxgGiAcXjVWlRTTmY
OKILI1okeWrDfbpo8uNKNroF8sAf4b16E5llqceIjn1S/CapSd2LMIDQPrS/NV7U
6ocQ8De/YsleLLY9rvyvW5jVTIhSkKh5jaaX+okTuE2Hh/Rpc7axW9WiwZ+sKz8x
TpFfL3B4z+G9/OdGQb5Hq4oZep0SC/urUPQklrhiwdwVtxVaTcFX0xrY60554EWL
53VSJ30pgsB81uUbYGmCvaeEr6UKdEcueJW05KvssCXM4K7V5SP8qZjW4RrXsmZJ
FNTdovgSSvtnGUjXCF+67NxsIgMQelqyl8IdlHgGZQ3Fjr2HvOikK6NBTgsHBdsl
DstHSKB+RWiWSM9mi7yCi5Y+MRvmxiY5LZ68o+FlrFeq9cP4BmqEaGyT6mMrL7S3
8C0uiwD1gE/0C/Y39XQJzGbKIglLHqegGKr3HSX9zfa9FvaR1eMFd7hXzxd9H3IK
G6MVhBMyo/OWGrPbbv6nAzfnIKGtSni4fX0YT3kF5XdIMRgHYIONyba8/FGoaGuT
mn300G0B3vRVV1iGlGYb1NO9udJq4/kLYi2DJp/3jH9PAkGJNWnTouZRG5XLKGZQ
ZW8F/wRheA2HIMAxxxu3PsjzWkBa+wLeVB0mnfQ7rHkjhG3jqYjRXYfqxOMfHQ6p
lr0dIrnzL/Cb2PlvD+raR3BEatShclHa1LL4cIG3CiBftHjUMENmcA1NWwuO3bgF
42IBwThoKnD21YW2i13rnt53UdFIkn1BRyAg0pwo3kFG6AlTpVflGS8EZjSimXIl
UbfClkpHTu8hOxUq0NsoNsQfiKA/eWCG2LLtvAKUeUIHVf6JrRSSM8QXuXw53GUZ
MPkmGCUXlc7kat7eyUhP8O//dx/lDZhgcaHFUDVntXraNpyj1Oh2D/WU6h1cdhXO
B6JlfBGLPh6qRjQ8g5HcC7cnKyM86LFLzWnfhPo/y2RmkDGl8zTebCwwzasfVIw2
AS1GYVieRQVcBlOHqj0/7k9muzuyK72BBO9l4YkB22EmQ+/rofd+KIpgRJEmfycc
YmhkUdzury9Iqf2p1yheljQHkfy15UYDuI/np8hce4c4SPk75RDVQR80VcSFyGCe
IM1inf9qgI9f2M2l6sfGAAr0xnZRdwdkT18AkQ3/0E1qEkFHwhRzsZew/GpSmwID
Gd0SjxtFrLmDrVVN/b+PjT9v2jj4tA66wt8uGXFtSjNIKzql6/rG0XAz2qWnoM5h
BBltKab5LqB5l/BKfa3hMKtS0TYmFsGYZokqZoU9INVnfIYM4+BQFCiGcWJbIV2i
m+1PChsFADoGjO3XLhEA8bqBLEFsu3bgEcd+F6UKd1k+rPSRMrrIZLWambt8XkjJ
via2SSyX2CqNsEKhP0I8UdVmeSAQ6y2HeuW3h6zDTqTnxl2UzCglNiPKuPw7l/w9
nhmUj7otrdSHP0+yuyI0j2eDkxaGVWmLjkcrg9ZAliOnDFIATSYBRrSqp8x4iqV0
urzk5zWzTfuOqvD0nXh2/iTppZB/fonaBFydzEGtFlIkhxLhkRq1l8vFqWvJuqT+
yzFhNCFNZnUbGkzvu47p1Sc7aOgT+ORCpTNa+IGIvE4HlHLLVopxsTXlDXES6EVn
Cm1xj0bNkRFvAXehkjdh6EMohSvX0PYVXkOPZWDcfFEHbNNcLuw6gEICs7o9jYJT
sdwGYNhlw8d1k3+C30vSZTY+Bg0vwPVQmC/AgLqEugLtm6pha9yXoZUuXpsyEB19
I5g1Z4+klBoSNBikV8W1ULidBwFu34YFc9oDFGva81iB4Hi6Gcu05s7toAehXW2C
ENHaWEnDjUAh3wQiWOdFe0pFoMVhHC2d57IJz21jaGtEoy4YE8DFzdstlDgpc64L
lZKkXfkmmMogwXMY8G45f3DxMP/XryISpnAF7k6nyJ8kR0VKmvyKQRlRdsSOVBUN
iFBTSnsXEmQjTIcx4LynDxx3S5+OgptcRWfJAVj+m7tz4l9hsPQ1TWezhkeT1Ka0
rMCYow0hjjZLV6WfI+vIPx7oGY7RnjqGbT8tExTOngpvTBo08IfzpQI3EgHOPfMu
RJCROM9V8P/TCToGPCxZjvPtIKZ7YPuei5TKtzB+tm8Am0pC8d97ZwzmbivIV3I8
cWP8pyrP83aw9kfm9TMs0Ffgsoetoq+sHww2vOVjyIjlIu9VLdkj4lklRZ5jp8Od
917jQadSoShuoUikJlksb8rAEsIfW+LgLeGoYbw6I59jJNAe/1zOfaFcLNClaWYk
ZmHhmLvdMVtaWqydcujuEGnBBHneeD4Y+P1FGqHhWUcLLDfR4GB3cBJy30NHiySZ
B+t1O3T1iETOs0m7kLPFgyQnw1X30EK+Kmv37IqaW+zm+xnEJrcWz0jGIAaEDYoJ
JzsODQdjiqpeCwVaBQGFA6QPUYSgSiW5vOoqhr3lhofiQEZjBBoGb6vqI2+Hd+2o
f3fAOLYSQOi8KlGxHRmL0v8F/5j5YGZNSyBmKHc8gAZw5w8lN1KthFLNgFRW9KRU
mjj4CbhE09q3KQ2yN5cRGEQ2cXoLViOxHGMmYtyxw0cPmRJpoknUEddKWd6VVfCj
aeu43hRX3cOEib0Ecb0JXfqNizRkZ4rIcKFaLPZdweX7RERUMjyQra6x2ekCZl/G
Qe4b1nhiB7fqGGrX/uZtKPMuQAzRTx8SENI5DjvSbzvIfhApC5fjKe3gMdxv45tW
jAujLSn+BLgfgZU6L3fEr9ds9wyCuSocapC81w9pyIfk7BAE15NzktFwk8Isd1P3
O3LMkgwK+tJvhSCWPcXfPOa3pfmokydLL0/X8twwPnMKIw/xE6mCPjSHn8Q/pagD
G6AxdkPQEd29LA609iKfs7OtO6mhYTX1Wi5FNBH5w9h7Rl9bcQwva82xqK4cumDQ
RW7HWaFQwbtxgLiPWYMEoavfDzRfT+Kzbz/9IA5nwx0LuNrIFANJPXrrG7TET724
A5sVp4ic3OYEUsf3XbtaAsqRb1w+tZJluVs0/LTKxKmChEWzoInIiPJyRMEsCcrF
bsh1w9yDONip4NgW66Aauk0ZTIM3ePFbB14YZEjvQoIq4kRBV8jZvJtYnSt8MWOm
jULuCTPP7vfm6vIaIEE6YTyszr2/HjtZfjdk7Q0NGBZS79ZTgi/U2R79DZuH9bnG
biiaK0azI9KJgWGqLMcYVilv5CbX5o3/Tkrs8g605VFa5MrYFzXNm71Is+1QbGVM
aeHSVVRwPc82C/jxtTVcBzGAcNosge13xAjKFpWK1zAyhofMghFVU2bsylHslMho
UFHRVjx8O3G5Io/LV097ECkc8kcovDCBRjCdqkr6dhrvw6wUr2TT/kKrzhZoO70u
A06Xy+CuoJ3TRo3WWsLz6JG4B+5zlm+LnMnonkLQYGoVqLXSqehPUu7cJMKpIP7g
Z0To//DuilYArHcKqbCRbveHOWSdz4c27c2+1Po2znNeIRzEDljPTIQz199rVa2W
prgrDh+b3o8u8tXC7XMut7odlmmM5BJkTxem3kWWGb3IuqXG9zq+3iCAPqw+72Us
tv6+2bZj/3k99U8KiPjchyoThP6ZVTYVLAt8D8brt7on9Df7yrK10emMHeiatM5E
fzdo1nfi9UaywoGz/aGv6CrQrdGhPWzanV2SLWV8sEK8Q7N59B81JPPDmBS1Md0D
Qihga2O4IF1IpdPyLYok8DzWpA+Z9V5URgYR3ku1DT6A/gmJIN/azA/YTVDdzQ6g
niMWF7mrEsqBND6bIIvBO4lKwzddqnpA4s4sg88w5xH/nioF7dr7YEB8KdsRsiyI
PGEIMfM9l6b6GI9b71G/FFfWgkpDN1X2KfOMmZ3+zvCaBq3q/xj0HQNpAKLFjxCb
afw8MB/YqkCO4s+UC9lbMzEoyPHbX5mxqqcTaiLFpzeVds7JwiNpRYsYYXCHS2yV
DI3O0rTfcFuiAoJ3PaDpkqpB6yOj/Ge1u2Khe9yXHVTyeYnqVGa1Toy9PgQEakaM
Z3+T0Czx6CiFKwTEUVJqqVDrv+u2DI+oUHloK0ABCtgJvKo6D9/rU8aMuVvyBiEf
PfkLnKExSJrylPMFeNe/I4STcEsCrX2bPjXa/u8PhBr50TZLyfx4RZK5VxRGSLq9
lR6U8TJkzQqr/elXcnFWuotbq4lngKwHeuRGHOfP+NiqFALkCzJBouIK3GsHCFh0
ePzPWfpqxaFwK4KnXmdR22wzYV6LaeaOcnG1gR9SBzUCoi2X2YgCSsJ84RGzYfmz
FTVyTtuLr4zzZq7u7N+u/eyQw7Vf6kelntGSxdBxdedXekKMsSsTTe+ymheMduIH
LwQzN4bFt9Pq5xqs8OUJolfNsQmwX0XZuCSZkdDJXAw+dMOjGhaguf8tf0qt/s2c
bUJjtRsz6gtVLEAu5A18vl0BqBu+qfgSTHEIJpAkPRlzWNyyVOnIp0PRCAYOu2Pq
JVRXQpl23KInW1oJ10/Bhzd3pQXMvvp7tidiX7Q0P9Gx5wjm1tzHbFoGWWtLPD7T
DB7fQRUbzhVeXNJcxQGjg9TZfTQJPfjc9qpR9znTloR6MvkKp1iKN1q430nITWi2
PX14ivDaCHkH+JKt/mERD4fc0tqKGg275rVnidfRgVwVmVhmCTaZPEYcfX7c4E7S
qfhSrLKFhZMRqw3y+h77m4BbYC0mRRRyjOmUN6/RSr6VrcHaiKO0H/AVBjjEfPNF
JIK0e7OM4IicHXZ3WghaGJOQyx+vGoLVybxi538UgEdpmE+/QHOsi/EHKRQMBvtN
7+hfxaz4Uqa8jGwsWWZH3+nmbR+TWX1jXyBSB8xw+QmxW29PZr4iJ8LsUC9adiyh
uIutJmL6fw8t3My4nrG6vckE2FDGOZo0bkIzicUI5S0VrfPl4mLnj/yc+kuoVfU7
TrT/fK6umfMzqwzEYaqb1tBS8X30CxwTv2DDFoAl2NUxHvIosYvyz5moDQjK0ren
fcetSKTVlS4hdmsrgJOzESLKMA2D5JEGMHCOkcfh6Luc7WO0Htd6B1+wsh2MXs9J
9FLmk4MjVZEEg2dPt3KNn3yEneNWrna39K9g+36TQYptUdX1sY/u2MSpUbEvo94m
43iY+TVFKEVbykcjzld9EVtlImjdK4P5uSDLBMMF9WAsCeaYzE1Bhl/Fe4mYXxYT
HIYvmuKG51LH2AZNZwGiTz6bzSyo7V3q4oLb/fHwguNhxlvlnFxj80LVUmB9yGHW
z37SYLINGced294NgYlEZAZit1cmPFmLTcUPoDHU2PYT/BmSHae8QYVhfzHX2vTu
RwSgPEFexnfqN5tbj/cdiLY6Gu9nCFE7YbC/bQevNYdgWLYfyoLX60DeKc809/o1
35ukg1TWKsI27viIom08hHQZm6DsQKgQ8qNbvtrT1ngDVkckuw8RBfqacNjCB9tL
nosBDAWMFWM4K18IBVWTuj4KimfoJPVC5clUmn3NmM3Xb+pudXuPffVA8EkWMSAL
u3lUo6gCCqbWaqGIZpDU9b32Qw7fACh/RbIxmcbQaTrY7X8yacuDvzzup4fs/Xxd
fZpw5d/F92hLOrMNEkC8aWFjEDgO0x7SHDWSqdnH9+q1E+HA7ZgphZ2sNNbRBits
iFgvl+5UaRqYmTAKJT73TkjQvlHWi/nI8ayryXFt1wX3b95kox/RXp4OZkngL6x8
iHKPjgG5y2gUiK7iSHhp6mhff0enUhtIRTiafXBPwvSbF2eQLH1sR9pZ+KsDEKJn
4V5kS60fr+tShwlSdMWNGKYonOfSgXEQ3zlCHG+3I8/+CmRaktZodoHO/HpQPbZs
KC2+BJTxEiSeUaQPPZbwvhiZ6G3kooPkT4mRSnCp2lCq6/zv5GkRwcZ/OKaJz0Nj
F9Rn2qw/uPU18Yk3M3LVMQJRctBK3IQW8r4rQBDPEzPsp7Jk6PiRWphs64imAaRw
m51e56nMj+9+6iWbLAeP49gNIZPYAPrT8ORjB9oMbEQkcO+ApCFgX743sLRJSRd0
INHNDH5Wk4bc7SfnRxZAnqyfPDlgJljl878N7g3rmNq3e4JWKi3toyAly+Zfh+L0
xdSfoqPDujQ4ZbQnl9CE+Dsoce2y5zXNAXN2DMoRT3DA++l/w7ctoiEXtqb5af4L
wVFlbR98jojMQMtqyibSo/LaeOhGoIhDcP+1H0p8kjP1GN0K6gD4hHmrm0ufnMn0
tskOKzCR1C3Q+WhCtI0r9xWevJW1A0PCOUCYAlPqwxtd7zkEHyWVSNQSVfDG083f
ogk0JRYx3Hy74H3l1UInidjKEFZxUNdVTu5zA0s8uOYUkvBiD3xILa+1x9hPBFl7
aSR5yIhy0Xejp9eZ3JVLvKB7OeqGjMSGks9vq0BxLTjLZoyvnuUR7v2V/3oZU4Gr
k52v9ehQaS4KdSN/DpxKY2JLYVvt2cmC/1XCj7Sr809Hdzuw+eo3Riu5+Y2PzapI
Q+RClkEhI1q4LrnYD6+anLHvG9UjbYsjovx2MvTWQHs2LNOqFceOaiBh5q8nNi77
fcNLrNoU6C3VQFMIOlpB5H0F/QxXp+AVoC0NNiOkWCAAtk0h1uGJWXY12ZAINqiV
z4Kupe284tVx6Q8AB0dyo6APt40hR1Qj4EcX1qNs0Aw85W1RZEayjPD7ygsGnfGD
ezaMfR56UYqleDW+mhlxAuW/zY7lsivTDnTdDgF9SDNfWm6hJMaDt0K8TM4PP3JY
L4HSh6h/dH+tcnsr6IWcHRqDu1/LMNzV2BlVwGKVY1I92rxNuM1C+/OxsRy68de6
72J6L1XMMq5wc5+XIUaVYbFTJC1g6EK7d1kp4oYwps6qfYHeCnpE8gm+fLoQrjLW
vk76IqoEOyGezAjssJ3LYU14w6yIn0fX33ZDbSseGklcMpj9htNMEq8fcL1q7j4l
CQaY3ABI6Gp8nNgJZauCAU7ONiZlo0f8mR/kK5+5RQOt1bG0ski8vUxPKw/e9FPE
ZW96mOUbXJoJgp5m8UWTQD7RI6yJdjHYj2BiWCejg94DE61VnXM2zQ/jqqXQkSWE
veFC51bDX2dG0L2k1+UYg095LyCkYdP5dPUrVO6P2Phf+nicWHZdM6j+6F0O8y/F
/qNrGw9jNRKg+Pt7KO1l7B8oS/yVym+ZfzqzhQVRdumV8Sne8cGreE0Yjuo49tcy
zH2eQ+YiiQhgDorILktqvnomSbaJ0NDveZdS23Vws6S629BTQUc563h44pwtIG0t
Bat7SsjzQBWxjWYtW0NB+kvN289G5/Lt7TgTLaXmHOaFzp10uIHOtJQgByUlOOc4
`protect END_PROTECTED
