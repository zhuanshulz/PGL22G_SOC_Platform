`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pY92BKi9cdHO60RuGP6kUR9V64JV4sTor06v3tpAZZyZYEAmHTy+dcXvgyFxQMIQ
9jnlKFWHzJtJwOzHCTdEXeFo5cDB/TbeTIOrfPgjQDyUrYwBtfAGGwz4hyNxNXNN
V6cVnCRoXcdE2s1PcWmt3nV3wk/uZA/0oJbABbCAdIfJb72qe+3c/KWpHTy8vZUB
bBw7EIZsgAQ97uVOTFwnAPf1mbx23hGVwED9CZ+LAK6+2Wg/1qKITeJAJ7IfP/53
23A/Lt5OtSkOW4x9P04PjjbJZHYXczXdTNUyKR375WFTx7iK2AQl7Xweo8QHoZdF
X8dUZ/Hjdj4JxGYcPBnV/GLmWEDiYzb6FvStVoUcWSBjy5jmpQUFYNwq2dAmVCEd
k8YyIofCIBgTWapT8U2kcLfhF0Ti5CEB6+ty44L4hur7Svlw6VtcHvNWJs7x7NIw
J4nkDqvzWZQNGAYNfHwQACTSj9LGiRabDUrmJ6FHPkQzB79UPKpmJkzrgYfPFkN4
/eSxkewqgrPEQGLwQIb7lt9reldjhJTqI81+Hblk0wAN13YKaSQ9YmY0h+cTGXNR
6Wy2V0acY6UaWG05yVhoapuWiFP3oGf1CWNaUjrdhRJS0k9E7NRbBcnYMTJlE9Gf
tTR2igo80oIrclqbSG2DDzKUajkn5L658JtcyJYlp65JQfywFGavJifvImyRQmlq
PMznFoEphxzsn+quqB7ElW6sPkDHxmIzSSMj66dJnc4t8KrfpKzLqbzmpeL7Tp19
wpK2ipNPNcj/dD1FA67m5s9Xupqqq9b/Erd9Mawd5mmBXQ/h8gEniEshFa+IQvMD
t+cdNaORS94oyPl1Iap3d3tU3qSQa/sPJ+8UgFWqCRMZIRoYNBOaNeALyVeKL7fh
6HjrmmMSHO5DO8ChKerZgQ==
`protect END_PROTECTED
