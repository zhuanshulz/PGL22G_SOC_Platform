`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xkmABpsX2ysoBFntxrEvMZb61A3SYwVO1EiiOiysD31k+0NMCv7H9U1l95UT0X/I
s6BfCR6AdNbijuxFTlY+XXazRpVEPTuzp7RZ2T6xUVG7URZ7WYnvfORsY05+BcUl
J9s6SOL7tUVBMApWnrMp3I860AgBpyAEzcphIMsCmRmIZy7ujzrOUwhwmd+FxHeM
YspdVyKfdVROEljav1bHgCaJHgPrxUg6U3Mh5emtrhdGPEdVzBP8MElzly0Lk5Er
LsIhrgkcnCoo8uJ6xxbWc4jLIHKfIn+CneDvR+W0+l9gj304FmjjnK473U6eUPL/
bsm++rQfy6lXkEQCi0UqT4ZCvaHwYYTjMWEPQt6sTSUOft9ZwIjcxx0L1evP6KZ4
YrlXFoOfAJ5absRwXukLYpn/Q4qFqGF1QaHcV9osffYTd9Nj3kf83lInVxwc8ySn
Ah0FL0+ySP8lfr/3YNFEnCxARORUV3a0rUu2O8bLRPzTLb+BCi9ZtxWCP0x1Oq20
VJpq9RWh5UWT+d+DHy+7BrbgUBrvUjdj8LwXJ0gvvtc/pob/lkZ9Vn3jCkn69jC6
NbXYg8rMu8tFR20dY47NLdJsxDzmA/z0OfSiIgK9Rl38JN+5qo4QdRptwWTd9IPL
`protect END_PROTECTED
