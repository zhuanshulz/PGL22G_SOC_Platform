`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SQHdkrnQwsjn9NNHAKVurW86/LNQ72ManpS1pkN3PnPoRdoQng3EHiqRMUASzm+P
g7UR4tOE/vclIRqlSZ/HF1fn6a8lfVqI+ritY11oThOiZS919Qq7zvEAfWY1n/Dz
ZPeFVil3gAGG6NYvtnB0sndDM54jv4KU5CBaWoFgN6FqlK78R946ueRbrLkMQC6x
0u0hOGK2YG1VsqV/gqWABVSOEwicUpsBnhJW8CIlXsxI2vvl+U1lI/xoDHJEfvRz
AcqvwwwNc3pJn1Z+t2VFBE+OUQzX/tUvzFQcZLvMCRJR3mz8SlrzWPW02rIT3uCb
bopKs45gXk96IaPjLp6MRUYAaMgSUa5knS86PG/fCrouUdeg8TKmwLPfWa+jHIl7
ZsW4/YwXRsGvaIWrY8PazZy1bpuFTt5/USw4M55jGvjs2t4FUbvIzZSnUVCqbsOB
2SP/cd+MfElA1xhGuYcG4PW67Nl5bmJ99bTMdxQLMxTQGETEwHJmWKLJhysta/OI
Q9kh/yiRJkOKlmcVR8fSxwO7NUuV8TxC0dADXxGHEaD954T4wsXcJ5QZy6eX8Jjw
fw0PeWBBWfU9zKTQUV+wm9yp3ygdOS7CPkuo8zkBs5o9IVo9/oFPxxrux1YnXALX
qrah+0HcBJESlvZOEWSs3VBKcx7JQRCnZ1jEv6O7hksiw9bQCY/1s79JbrhwiG4i
sDA5Zj7RIEL7HRMqI1CHyP8hS7iaQevwWNGvlCwl9dMZR3g8Kx3N/rT5uy5NA3n1
8Td1+jEhkKvG1ui1HSNXn65qU1VppGoeaMs9SoULUsU=
`protect END_PROTECTED
