`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rZPZg2WFAjGoE1MK9FrlYkJB6sSL7T7Yt+vi5UbsKjficKl7BHf90xJTk3pOJaOM
XoP4W8BhlP+9F1CNlWWFqzMTuMhqZgAJ2SriyHgFvEvFwvXbqpRfyGyXt8SaUrYT
EygpPU74cBIUJ7SDc8aMDuUSpARI/kYRRL6wNrcnDmgD9I1x5OZwF/NV7grHhjoQ
AQSqPdxXyH4EFLWLZM5H7LzKOSbiN+JapjBk4dr9H/JH4903mfz8BaOKePmq617w
2N3GVLtR6sU2YyHUKaz5RYfxd9LNgfWnMeXRU2cMzQlf/RoFpVl32IlohZ0QqG5D
3u+on1oLN4N34MORM0dp68QWXvM2++5G88F8jMxjUIP3POYX++Sx+eOoOzGnRpxe
qofmgv0T3Lnfc9nIIjBg8juqvY85qz0ZUhOCgdyOX+PHoZBYup0FT/m6d4zj8+6A
ypNeWSrKX9Kbc2XC5EmhKCIVmqGfomc9csJY6AmIv30/ojHGc7hv2N2K0RsKBChX
g+qx1sxCQ8ui88GUCvLhaDCPSLsBhHZu3NfDGCZ8RozWmrazKMrixAEbH2Pi0zwM
iySaLy5rIHv+ySmeyJq7quCsLo1bbHTOhZGVY/N5O2dpb59p9RKudWih3CEWE8nh
5qYE96Y30aJZgzqbpHnkAIeEV17E8G8NyxAPPdqVCzKJtdBQ+rZktpZAFLgyZhre
4VqBO5aakccMleAqQ08o8GUE9RIMMtM25RCD6JYEYqrgUDUmBuqbRCrBcuyN+mex
TQBPFaEQ65sCwXbFJe/vM9glp/ejn/tFmoiYblqd7CfB2jwAM2ByfxkoB3p5FcQ0
GwYprJZpJ8ts/J5OZ6q967XXAdN4iQcaywr0fROaMOa2gdTGJLxNlIkNoCm0aMak
/KnoguSjOKzTrX/zOBWqbjU6qOREKT2lqsy9Ink0+ok6BhjkvKorNgQ7PuetvRHV
SRDkejkps75lFigt+oi2oslkx+yANBwwfslYfw11M5DMoB+/b9BXpZBjy7vAXY8z
SuzM1op6jgFAD/hCbOYJG1/JzObrIQWnm1ZBthuYyOkR5ag7tohGG2azxjg044K/
+8JW+Gvm4bNFzKahW7EELgZIPOZkCoI8+ioYlKqZLv5Yhst9P3S+GMUC/wV7VRQV
oOOqcN9d3glmo/oaT3KtOn1Z+owwgOuQID8hdci1S6XU/txMSLoReiNdlHX1VSWr
ig5Adj0y8YFD+n+qJ9lG+nf4gQ6bwwQgbq/efzDrQmbm+vpff8Fk0Pc7UKiHVCZQ
WpF01Wf3RzJ8Ipv5uto8tdSye9PgYTmOkJdo7dSUKjfJiqMzXD7r0GbbVK7jZEiI
QNwkEbCCdiHfrfRqhE99h9hHcxqBkFdHKHCS6J1+lJDYMAHkeUwPeVOQdUbnSsow
gnZP7VbepvFshLrtWG3Qg5m3tRyS/ZdPw6wn7E6ZO7eiqKFelA6g/+OgNHzaSUM6
rXMXvo+Fzz/S5tu4XojYKOQ0v35jdop2B4cNX5BE7aZHxgpyuy9rh0Ia/6O+1kmj
mzef8J/dztb4BlQcAXFfuX+6ddIAV5TuMcocWlztxLX/YN73nRrFmPHe3re+mU/R
XWu3NHvKS87qYrBHLsdLvr/mBD6fxJ6YdFTi96Jp1CiT60xDTXzDZEC8ZjEwvzuo
Cdvnny61G3K30H+cyO5mjYjlaLPP84Lu1PN0r2lzgJBgSeh1kZdLdeRLwsw6U7hA
LBPZeegPNc58aN5n/R9ZFDnC3zO40RQhdDmt1LY7j+ZOYtgKUm0TuNIEMhQElEeE
Oqq7aZe9Kpk1gFj0LFOFU9XmE4uZRGhzwF6RKh2W7z98NBs9Nh0WcR3NYD6hjsWY
YjbnHNkQjRyPKJTwJDU6TQqsJTI3ZFrBxq4ljea7EIxoC+huHh6OOpOglKWwAZh8
hmH32I4d1Oa4vuZC1k873fEHJ/8y6L+dUns1TyysbIRD4FMdzf28S8kOxCfRns5V
jNrsVeuCVgdIN3BVrkaPrU3zi/Q9MMwc6/1FLo2sXTAgt9+00G8h3mHmRkDiOgwK
r1HNqgXYm9I6OV5HtUTeh9QTwEE4rR1EIm8WOwuDDp3oRbPUlJRmauYY8PZxI/zM
Cp4MjCIaq3byftk+E6sxWKiJQKy/9flPiRPZ9aI1cVd16ebUKPedYL8M4AjswbOv
9v5wyHflas2bHVxp8uWU4GiYnYfsajVtOFS7AmhOOoI5jqvO2/b3AAnhzNRvDtSm
OZ/6PR2bgvrPv4vNBOOAKt10aABk1GjVhVYtcp3sjBtwasLSpHYVZn8AxsCLBUOT
Tc7vSb4ZFHO06N2Ou5U85yj/i4zhjKH58/hay/sF6CRXUn/YHF9OIMwjTrNVmZRV
VBTity62zxjLB6+uB1LEmI/+2OrtpuCqrxW7BWyxF572nDdiyBX4CO78CGntAiHO
Ceh7rEjWPtpZ2OT0IL/6GlhI5Zthd2HvjwomjETJ0QOAewGreHjLB5yslRFpMylo
/5LJCTBi1thN35dSrT/Gv9yhLp9dVQfZwVd54MefVzve1B6r3RhG3UG90KSq44ko
IHgQZSLQANzcDBCHQK2OSonGj5YmAtkQipO7wn+CehBmv8+IEKDKlueAHAUblTNy
FWfGeXmEXCRZJk4SmPPM15MXOSQJSX27gQ9NZBynihJIJtYKU5aw9qN0tHaTZ4ri
Wa4JUPw0YxE7+lQiignnV1sfomTtPORG9ZFCz1xMLsYXuIcMGj3COd7q8VTxmVT/
gSA3O8nqzZ9t7vQTebXiwMRv7OMouHwY+HfAfI5psdEG23yJ3GngYMZI+q8Otzyg
igBRdbo2szbi5CxfApG8FM/t1vvAQMWsyGYgUqW20h51pwgEvntr+4sXaCEP0lF9
vJfmUemeA4PlsfHcwgCnolaUYn+8uzNR2Z8E19PL06yrngULpKvKHiLesrvxUY9y
Yh694/n5eCKsPH8Rqf6cZ9lnjYt0GKZZHCjkqwErsNKA92GOYWmpC9zcDGClrn6S
IR3xorA7O3fodoPiph+oXb+BbtctG33zFQjuvNvhHThH53W3onhRfUXkz/rseN8n
ej4Zfgy7eQCt6VMae4X6qamLC8jiBHDNNAC38yn8zgcTVJqyDAavVthGJGvA/srZ
p1hx0DOSPkMALlQUVO/J+0/4xmYj5JlthF00+uk7OqVn/jcYFwDjqYSN7aWFOVoI
5rLdAVYxM1PHfNVI4f99Fhfi0H2M5Vrn3yArANpB0r526zN8MIkm2w4K+f4d7FVg
OmpHFSJo/so68Qybf+UPEs7g2QeNE8Nv5w3trujmvWE8WsR6pcE9N7t8coiIGuAu
6QI53hrhMCC+tjxxcRbNVqPK2KUguKceSkKbibiscp1jinFoGl7meIDL/95KMlmd
HcTSz0HSGc+tstDkiuxvkFn4xMnaGCTV4tIkStb2cmllsoCAugWoYQsoH0V9Gcya
vjPGnjR7sPcMeJ7vgYpiVpP6JesRTM4hi60uc28yZTjdY1Huwrr9NpdvVk/Qia4z
jKDsLOB4R1p2Q79hLseg91Nf0l46UzIly9zS+C9qpXS+2OEgepQhU5s3UoBFVd3+
nCiWpHOWuC/PYbkqrZlVcrk5vqXOSUA5w12OUlYBVPoJai26a8V71PISGOIpNUPe
K3FpYialQS79N9v43FxuU7Ej09Wzgh9KqhyIqZ37sJT1vzNAYk6uOJwNNdR/0ilb
hsCNGrAyFEyQUD1I5mlXXclz2fmnyhGKkHFD3ApzFkyORqzODisNvNrFFKTl6yAF
Djg9/Ba03LOmwF3dfbmIDxK0fTxNLnJkqXNaLAZBauy52gMvGPJ4ziB/Tw8WN8a/
6KSg5wa7csaG1ptyREFmo6pIQG1bFIOFzqMsgNxWrWdajyO+8xt8BjfIv3AYxjIQ
PLZ8OmwyZeLzmM7guwmHGL0dKnZrZjkP5kTB5stoxpPc/5liB5Fg7IqGtN8AtFwD
91oGmkUgXxECB0ujgfEUTkbCMJXwDX1AqjYAgtlQOg9emjCxfkFARORKEKOCrCuz
WKDGNn7mIcNox0Vu6QG9ugNxQl2NuC55O+cVM89vrrwj2gXb8hPaFVgS/qVa6c+T
2x4ZyYLe7qrjITLWDKy+/JOZYz+kvV/lM7Uxidalq2g4VY08PO1UVFQD/2AF/oxf
+RR/pDYFE1eBk6hNvQRwk3xTVvUBRJKuTqoBne5nT5lt3Sc9vvE2a1QZUBEmifQX
Dy0cL/u87sG/6tD9yNTNoY8q8n9RJT+WYj8WjCv2a6Z7wCLfEdK337+y2FiMGKsH
crt6QEqYkpFIfhbyLc24DCSkjphNqul95OQGNZd1HmrruxTm0GHwcAqTpNGxS6jL
BK+Xtq71ws2mGisCeWAKlASkZYqbUyor0Oiht5Aormh5RLwDpjcNeNNv61Xay3qc
h9KUnpY3qmNLFCZmkyNTSaj4c8Ly40qdEm+sz2J2/nIrmork+cRgg9W9DH7Cll0H
GgfCsl0f+C4ol1QjFDwe2qTIPsSNgO7DUopizyuK1PjzIWaY89Sf7HvQEj5s2b+A
D2lEKDqfmUpo0mxbcFnqXmHdO3PpHWLKqYtilpUQkrK1t3pjzno44KliCJeW5a5h
q5Ra46whii3MsNlhGKoSpscB7jHEk2TWCqKunK0m8JhjR63dGQYQ2r+Ixx5Tyvpu
n8GUbE5QhaAima1DrcUyQqvHMgah83hZYjb/TLF003xjqrmMB8T6ItTs1GxEpJl9
liOr61vumvr2B+K7iMFEKu2Ty2WdqlXawrPJAmiPsHEnuPY84Eb7nkS9Ozi4AKrv
U5x+TOY9XH1+nI0X+qNnvuf1dL3bgtxxo9U3HvzaCno0Gzo5EEsm0VB6MjL1AFfr
LjvqLf7dt43GrX8nB1JjwRS8nzOF8pSTIbD+XsHRrzx/W25LWFKXihClcVy0miCN
AfKjMYYdCvq6pnYpK5jsz74c8JDhazKQu4aeE4DBvMblVF+Kaydxs7yNUTyRPbEw
DpJPmTquU9qu+tuY1n7hzXAnfF+DphgtNMIg9TpiRAZsfs21+5Wh1XF2AQeB9EZU
vkBalO6vZY6KNyZY2B1v/dctynqg6O4ODPWVaet0j/vWlXefSC++84c0nWGIRXm4
nJT6P885bB+azHnjJ21msNoIabnVOErT2HfIkFXO2npniGnZIKN8D9TaQx2L2+Et
0fsiQYYRevzyJqNh8SEhbscYydCldyDxtLh1HjP7tl564G4BBhKPqGVQ0RgaZLZ2
tUF4L+fyoD/RYESnMHwA1aDAQXR/j3SiXKG5GZA4Gt6vBRxLcb5GG+vmcJZ8d6Xw
XRqOuYRrabHP7OsW6QBqIsC3jACZ4eVPQ1gkx6GsD8pwgV53QisIyqQxj5z1LeZ9
Z0B6DYqrmIEeG7rStdXxwQVMooxgQm7kX9+uERPkGsxbnvLCwXaJ8LWFl+HEjsHu
mihqoJkKapSmchQxAvvAStGrg7ByLmPa8PrS6mBqGUFv7burLTeXFQGMsoNR5zgX
h/QX+If/lOZ/EERJYoXLk2m5jmrW6nxa9lEB3vUdDrC1Z41TdHXUYc1aTwoEYfUC
4SJRRaLtWdd3OVIzVgge8emBKGbmNVKuHZYGK4CmW947VQh95kgmr8dkrhnNqoDL
vMlG9K3N0fIGmUamCErnzuD0tj5JWOcR4e/O2Jo8KGw37UeSR0reFdDaAxBPMAq8
1/qWqrmXzAl0JIcDIcbfB/Rk07pbx/nhw+KbYeBd7Pp3Fur4cVc+mF0OylnBLyAu
elsZlPSWkspayadUfXcqLasYB7qVn+NEEQfJPilXe/XKY/Jni8rYj/6Or/3kYKHg
tzkOV6KcJY/9pN1QHy2XVoY0deJrNF0Ba3XWG6R5C49Jaj3U19lmVOKrEnqbqPDJ
rEGuy6z/q4+MDfefYM9VR30WFZAguf2kjZdSZYJHEzwhZ5x1gD8Yo2umuqmMWAUm
aUMtNKSxCS+uJI4m4NBGriUAie8+OC90liQUw8aBFx86A/6wixh6ZvI3xOhkGaeJ
b40Ajkb7+dh04YGd2ksLsALc7crIFBDXRzyCIj8hcfs6sshSfgmfpwJc6B4UGyge
sg2DV36AqA1VDE6G5J5uJDG2S0LdYTJQBau+gIOFLrXab04aITihke9jskGH7DGw
gLlOVQJdDhBnsUJk2EY6emh+pYXYCZnEc1exISDyGNsmOtExw4Tq2TGAelst0Q9X
fukBzs55RbLMWrsC5HSmgPXob77shwdg+wemSFxNiVhAlKArVogJ/bRkbldmmDkW
v48S7SIChWV/Hy5g9YvgRfmeMAxxsptcznV09Ae0s8SQnFq7anaePhyd+rstBMJe
aXVwtEYWp29lAh2ze4o0NiA5w3eYyn5ekm/01FUUf5U4Y9iJeETeddgQkwIXA3wV
YbSq90uWklmk4ebKy+agnaXYfXfGdpo/EvcG7bhXQawnGNGrDT7yIt18nZQq1lLX
O0Jr/6YH8SEtYQYYHqRfUtxEdoI0k3DvGgXux57vzrWJRogKGFjBKkWz5dWMqAVI
zVCk0AWUZoKLfGm0khU3ePShYsYN+MfExyT1h8gIYSWlMTTF0led7x+50FsxKf1L
NZS1UykFvgeLvKbE6VTquYv0CEQtkK8hkdoewHz9bL3moiJFVUBAr8prCVPqd1aS
k4DJPib7u93ls/JJ85oYEDIhthgCRl4xjJ/l5+8iLIkQyCYo0eFmJa09UbcQnZjI
u5mFLbCaU+k07r4Y1fDvKJlZtiK3fc/A0OdyfUOihE5afQPP4x/4fjjf89f9dFbK
0slA6kcVRxFs3J31YTVMEepgaCsV/8h8DHMlbnIoXssoQ7HwM/OFMAE5zryZFG6J
o5bHHxF9pdhX3mbazVacvJcEUDOeMf9Az6toSykUd+ozibQeNmxHEozQd5MmHd+H
jqrt8HsOTJq8Mb0UkLS9mOyL+S0k2u7A9gEQrFtn4eCCg89tk5jt3IlmCDJAOAM5
sJdr7X3BZ0Ez89nQdpmOimcXSSfgw5Hgeq4iPfKt6vp30pYoROxtqKuYAY1ME/KQ
IavsQ5KbyG0Qu1qXDHkc/1Xza9h4J1tWGv6fnKfnFZqilk1qxnK7DZISlSfylR3R
iOEZVQmFq30ddwqo357qmgT7HRxXCdJ+tagENiuTytv/eL0vRWl9AH9zI3cr0T+G
JiGBVI3/T8M12NsbhQBF+8kp1Z//DixcDvlXcuceN2rtJfE+7kZ3bpCBBqB4FqNS
GYNKTQSUVudD3oFnmHLOEhW5srGbpJZgZ/pXNiZKP0xKFA/PrEz2/1GPGIe7ZGX+
gijzDZcu5K9IL9px/aMH+0FOJQJ7XxWCxMLBo+QOgluDMctP65uNrFD3HEght45u
mtCHZi6Qk/od1MKOqh9MNmUbHsWhsKOf20Ey5dYYz3IrDgBlQMu58qaJAMPGKuTM
RdT/9QexrBGUZMnRQyeTwJLudWv+1qxHNdHXRKH4+SkDY1wW6f9SXteHXgL63m2B
utXC/Ydr4L82tSix17drU+/VH2EeLGlxAsMNIUohh9rdY1yUUZ3uikILLC1YelIe
wj0psuwR2PKQjA3206zIqe7y/4v9AXgpHTUpRju8SPOvtoBCSYm8ebulujsbkyaz
dpqfzDiP1KKnbvq4PNqMTud94yr851Jj/wWobgc0qpPy9eB6RKd5vK1m1k93IQeB
WK0ZgTQ9WdQ/NMXIumAyfyXdmV9f6Ck7H3alQa+Jbi02qnp2p5ql3+QN5jIDNh/e
JRv4tzhVA0TiIgtrrQW2SByJcePlTn81B6WExmHnGyDeDntQnDKw2S6PSR/oMS42
Rc5UIrqnzWTogLRkyR83uGqffpuQuYWB930Xyv4+vibm15kIomyCKy5mvcPGRS0h
DQaqsqlewq4oeDceulWorBi8WtKdA27DXM+KpWFT2Od4FPvP4gi57H3B/eOoLlgI
1zZWfh2k49MtoyhGD+Mv5QKZOfgWv/QKlIAAI5vVCt/KKrgSSmmEGvB3M+jhWmB7
dbNtjDpFbsNEcJ4tMvy+8BuukSfwDh/plncG3aLExpex8Ax2817Uvknpa5jD2Vcu
Hwv8Hu3ufO7SHhjiGxq2lIykOWnEL/T4tkF/Qa+qQFLNyH1L47qIaDdlb1CytRpQ
a4ZLYfuwmwYpdYru96ChoriBVNXV0Y0cRAg+YEXFSChVvgFGjD7JdjoAdhkX/bMT
VxzJXVkmElJ4gScyXh7uhjX+4ZH3vey0ev+V8+e7EMLweH7oze49qMWRlUQ6ggLP
T3iWFILSCILBuVFKndJHiIfth8TeAkbgN4uDZBg9uWEyKtskBRZ5NUZdcW4lzAkx
taeh2t69I7Y9MUdvFoPuLk8kVlwb/TnGiBkTMFK/mk4Uu2vMA8ogU+yI73m/2rec
lV6581IvRlM9WAsoVaFGKcPoV+2ohlD+jOBCqiBiytyBPK3VAj2+171moVNtstuA
L7E0I4i85gp38aayKC2FvBV5PDmif1faQikfIrUGRR6salZX9MtEejSBuIVgVUSN
+GQ+iaIxEARbZY6IpsawxU0Jof9q2mtEsKohGhV5ExS6c+v0CgPYFuZKQk2VU9jh
8g6SEqSjRw2cAMQx35aoaf8kSOmZ+zCDfY31MT5todsWrFKd6tBNMwpoJERjYcdZ
0cWRc2ksJsvopmEC6lPcr4nDH9q1CdHROiyu6V8f1MBqB0NyZx0SNJ/aWNas6gOe
uinWkDBrvDqGilKDQ1Zkf8KCea4H2KjFOOpOZ04e5pUULGla55vQSQFJ36zA2/7D
4+6R0NjuMGAtMVKKfurW04jXaxHJJngfcGzauNVd/mP24crs9YoU0Al2dSowRPbX
xjslL0ooZM7EfW5ocVaL+Y1T4w0uwuayCPcKlu+/P80nuH6gH17e0MYrWBJJsjcX
1z71Q0Vuaiuq2F0zHLkFU4ywQ5n+7e2klquE160GXhbACsTbbNtBygRMKHn4xWN2
YyhoAJsYFtDfDq3uJOGJqBWlqCLyZg+3vc9FaWO2yr3HqsiTyCqy+S4YtWHJyn11
BD1afpvtPsRGboUi8eiCJAmvOTlq26x5LXOyYSrW7d2nzgkf8ZrgTqGSPUeS9wNI
IhnxHnhRp1cvOvOCCeKFgOKdMjFhThG8W/H9OpY3IGVXR8DWPbpq3b34zwe8J4Ol
svtBc0bYNWflzsJxfn4kDueM9B1VuZcLJ7W3LKI6QHI2uvL9MJBYgWzcaIzfGkRm
JzHv2mt9ppq+A1Sh25pRIyyjfP8gC2w1CO9VP3eiiLCRtWH5qkxjR69jh4W7XrIW
UsVjWOl/nAM9FlbHmwaDDsFFjyM9NokIiI+hF8VR+Ouhyuw1EXbQJBCpsfSMdE0s
oQVQrwAgBpkXXRi6cevDujijPkFIpSggylmvz+rY4aPuYO5FuSnprCt+8zPnNSjd
8zoe8avafU+Fbkzj0+/IBy3nLmdrk8ta/1pJhwKWX7Lfr80o9EWRv8UGVpNUDmUp
yl60MniXIpxohno7E8d3Q/XBKqwgipbzeBoP3IR3tIcaiBZzxBSMDjCbkFvg3NVv
sNmAciciuB4h+UWS01PG79RXpiW1CUlQ8IM33lizRfyuqUCgGC15sV9kuO6yD5Fw
ZUPdTH4mzE07sg1SeMizQPpv68dVFzVxJ6pbRjTzM5PdYxFPolY6KdA2gNqkJyfd
9eBTmnfZ+3noPfZIAZPBmxk964fOJ6Gjvz570RB5L3uipp41Owm/Go27lcV9i7Qk
fZiA2uyHQl4GiVwtAkemXULjWLK/Cyz4p2dHmdFMHBMb9cooNMzVm6xA6H8oneSW
2xY9A3qoDNvfTdHawxTbdqgmbgdxn9qvATxeZEZ9HXc8LUo+Dqd4i6Qcpp67CRkM
nJOIYH9GXjvuYD3jWFekaYy8tnA3PzkgpL5svuOsP+eaA/jmYCRfzUxKb6hkRrsi
4VWPkGr/qDVgr/ZzwJr9SAxVA+u8KF6g17ayP5iO0bWAtUThlBJpvp+Q4cKv6Jk0
CUdEUwnXLrA14NwmMJ9R9MISbUKdHF2pXPKXv2hEBcka8gD0n32zHlyWjpeg4cV+
IKf4umYoQX5N/JzzdFH70E7KEtUtz0gWAMXqcR9RvdnHyyXv6mxRkI7kUD5no51d
Zi4o5D2i+MSTzRjJj/zDHKeTXlaQl2rjsVTZjgm1j3197fi04rqFunpiiDIQZKQM
A7TbGONHIo567RG3YoebcRHfgrD1cmqrO0LrTPqiuxqfiqd0VvOHvBszSOAEVzSF
ZFmDv6YWQX2UMznH4CXYL8F0rTN3IZtSv9BjNh4bCj2fJIOOYdw55F3jfg5hYTqi
8efAVRQdD3fKtD06U1h2mo6MEekt1WIECYvQdmWrPXht52gky12aoG/GEi9aZrvx
TNyy9/AGDNo1vGpOpFdgkwWou8VSabzjnF7hCKkMRM/PSjFso9iHOBSvdRAf2o0s
98xzRXaer10J5uGx2DjJXTO0SXBIwaDI4AsahhwGvvIrf8D8YipNFl+SqWNpgwVi
h8qK/3n3m8b1RxZR8GcB7U1CDZy7EVuJIrHPOzkwz57T/O3n6ckpaSM5cv4R/kKL
59aQqmptJiI5TNoLPNXBMiytYgPQS6thrdTrX5mifjqjDd8Ajly2YfmihL7ZSqsI
w0UDj5ZVQGFszUsQmtz0wb+zO3cBjd36vcTJLrUaaIYRsnkO3OoYkxf28YGQpV0Z
9nqOKOEAJ2Ex3O+XTFUwJXLqAJwChgh/CVoTlSouvSesHh68R4pAddORGuEL7Enq
rr2jQMDFzXdLqqUpedRBDyb2s4pmh2P81FNJtTLejAoULsn8YRpKodOBCkFlount
K7G8HfGdHwxyZG/TxrJp/nFZSTv8a1P1NKIdYXcsI8P97grb2UQxHGg2Vd8mie43
XYnfCKOijy7gq9yTQACCO3El43LfUZR1g/RH7ar1omUkoMUJYFk7+Kzm7n1b90Nc
uxPKDzg5dg4uSBZg/k0LoyWAq3GNwejrkeSXEwgX/DijufoRji4hg63H9czjM51e
va6TwTJi14kGM2rC8xeo9aQTIEVIeBk6pEWJpajOVWkK8MW8kSV+tddEb4Rv2OYV
3H9GgI+OGH86uGTWZXLzo/ZB8J04hr4j0TYKr/lSPkgWljhN0Prw/OAOO87vLJVp
W5p720m+UpH6kTztDs75wzIOMx2Y/DbuoMvakZOPKlX5i9zhoUvvXXye5LBT81dv
Zict39lx3WsGKjNaR5g/4gBm54DqYT4ipVrBkRm7CCmXiHh5QR7Rf9okb56RX9Wj
SmdxDvil4I0I3b30aM+CXLMHpiI+zoNr3IT18FoVB3YXWZW+peY+cDZwEabCH/75
M+KOqZHe6aM4k5ZvBu6QDrz/puaVzoGbFMxnBr2Bpd37sbEeP6w9FO2Ca4pmW11M
r3NQLCAkVymhIZMqm+2ZHaX81jHpxUKje5ZprGRnC0WZl42oahty71EsH7Js2M5g
2014CVTH9gvbeny4bnSbHZEgoRW8uLtfTcgJNdZqDMBSGIEFs4ID02c1ydGWYOys
ux0QOIl4FshM0NJM469DqSH8OlzO0V3rRFJYsrQ/YickKv3b8mOzTY0QSX5WXiBA
RRHuuBGtNHdVXWykl4BeKFAOBCXZ/S/Ecifx5TZI1E7ahcaLNy2hDBnCPFy5q7y7
hFGBeeXGymDUuSWKQbdsM2fUcpnwztXBbdaUd3mK/ErjJeGvVSiou+3023hHgj/J
ir1aLYaHAm4hM0W0kYN/yWS+tOzaQYMOPBR5IOYDQUBbh62/sLWACtIwNqd7nYfC
hjG3veElZKjwaRq0qGEA163QgoxPpnKHUaiAFu2LzjkSzQXnzLMxssWH11YtTsnX
LPv9CLxObDnUTGgW/cNQwRsLP/P/Yi043fP4oYkJdhOSkbvJpfgQEMEY/ZMLueLX
A+laMyw/plC+AQSHdZZwkQzIE+2zoPyoE9qPDaWnUqxvJSzCw5L+DYXhvVDW7CgT
L6C5xIB2O4kNGHS8GfhdZ5NwNY02t7/d0C60YBZp2WdHSimkZO8LnL6zoiUTrMUX
M7ZzI0HbNg5CfOJkoWkVxhdWuMLS6K4fWy2qOgxanvpN33QattBwlN8qyYwNGe50
fhRJ8a4AjFZC7HIW/SUu6+7rLqb51Bcj6Qusks1VdNzgRTVdRmW0aTagdbrKV8nM
bTRFgy1amW/pzzKPoFqlnNe8WFLDIfI3UPXU+0fvAhxa/a+ct1ikGEZgH8h4lybO
NN3j9UPE3XlE4t5s7ae6NcwqamBBN6EdttGESLjywYc6VFyj+hVaL5Lt0lmg1Vzp
ir4pH4+tJMq/Lxw3kO0UAMsHppY8Vk+k7OQeHtmKIlxjatctDcIrIV1c4qLXeBfo
P27bDFs5zvOVr9xWYlyXvAOvl2GAViQfeBj7pV1X9BfSN1DHAwjGVGUFwIhYl7o7
x11DLQtkkMiteLgY1TgJhZeHhtrzHWpr+EPIgx6KcfKsgRP7B5ku5/aOWGys2a4k
UzimIoUnHgGj3xgGN8429XscQt9WFbtYQUybllVaxNy0I9XZVOl66Bs0hNLuO/D6
Oma9nsCT1QiC2HMYPI5oxqt7NB+0OD+fkdXyle2lGbnlx1C0bOLndLmChAJEHg3W
Keb3hT5RzMgHmC6hL1D9UUxMlMrei0rwDWVI1QhaMGRH+bJxXT6qaZ3DPhqXZpOu
6jU31ZuiFQssDm9BbNKN4/NiYs9OU6Cimtw3Qio5zCogKvQit3+X0huH8zomSeQR
7Tyk360xYHb2ahMnsz/cp2FGMCP1+xkFAFZaLf3NE0toUlX+grPzxkCuvIZO4aqP
vpkyupc4HE7o7eJjHehCpnfXyUHB764CIefFuE8PosHuOmmLqiVlViizmbKd18g2
jBAC3LB00+bd5EP+xdQUfW68uc7fGUGu9jBY7wEupgnLFlRtWJJix8Wx1zGkxz8u
OGWHfilnzvoJ26nEQYjJkv9MCNgKN2KfhWZy6tfEER73Dwxdlg8ruww9smRFtn3k
mBZlkuSd/3YktmIztGUo3siGoNHNGKKhZs0x5kQYiuKlj4SLgtgg5xQLYRxxl3kv
FlZllpPMijggCICwjfVtD7ohSmaQTYgC/oijlfw/Pd2i/tsptBhEp6CD7c+JwUSa
ii/V/q7VzLTiV3YVmyxU9lvMd1oezh7SPKGbOXoaEkbWVYIIDDV2F2hSdHJFri1b
iJT47kn7riIX2F+CUrTjA6u9MSxz8LesGs1EtIIHIgh7xytFdrbpiiFrlGW4TXxA
a6z/QrFCeodwU9Rk2ms/dn8Bq438o9XOG90m8hHOpNyzLQWaW8OMxe+2TLPNZzzL
iB7xk2hH/3vMabBHDmCNofRyexSyw8GXpSZqi6OYx6njJvRTmFnzmXawBgd8MXGm
42hFbMy1o7WhCD3zVld/Bf4oqzqmGxpmjxiq/uJCVvS5gC0O1G6dNiNSOCEo9C+c
iXBSgJs8y9xXAZU9q5Z1pNBFvIyVNcLwJoUWCKGMe/eQVjWsU5iNpVqIwlUeCOLn
OzrSgLYj/v0RLE+fbKIEUMdKX4i0AdPJtaUg2oYVlNkBQMFaYCEH9pJP6im68IFr
A1c64rTASA7yRX8kC4c4IKku+RYQBP0tYw/4i8WLgtW0QtwY3Go+VKaMPQeatgKg
5T/fxvnHGhfnIbLV57DAFCF+O1MiBbIWxpPfCYhrZepS2tT1rb7rPVl1D64ciioX
xkJhAeejHzrqa65iRtJqi+vs9wfjdoCIkEUz2JAc8jn2LxO8Vmh1p1w19fcvKTHM
6VC6oloU9lDqvQ+q+ZsJlY6xDttUM1ePD3upsmdyqwrgviLmtPiCGgcFMn15mt4e
3hQXKUqc+50BDa8g51yG719RXh9IoaKABW+yBgz9faFZmAEuI6athzGgZe1BKz3E
A13/A9zFde3yiwCJDNhoV3MydRbCtjy9CnPJQzbBXauTC1lNHefyZb4kTpxQvx0s
/ucIQFSYSqTccZ7iFUI1fIFvIWka1GhS66D/vygRNY/u3au1bo5MOrmufYOnDi0Y
vOuEQ9Qx3/bVm+kd4wdwJsi8zxSW61huxVNHAbIq/9/pV55SHSUca+Xd0HnN4OkL
OaccytICNZzzwgG8M+KLhAYRxG73Eto94nztIRjOh+1Ake+8HzE+z++LZApBEVTu
8ldJCjaLCea0DsgRBOoA5r7fCy27bZ3TL75xTeufoooXah25nh4yFle7B48fmlid
s+sQXQiKVavM9tfQ1+cHRKiW42aIigFWKgsi56wXmZPvQPg6sQQFXajcAqiPHQHF
+tGwQtFQJA/GaPCUrCcu0zliaZg3GTOT0aDYxxF66+Ilq3nKU93RnWRKBSW4t9kW
5M1T7JugkMro3oUHgjpGveXIsaJo0J2T/noIIAvcKLEujV8zISwSMj3TGUfvmRQt
FFB8OzNfBh9zGrHF1yiiGvle6PYFka6SjcfCItSdVSmCbpsTC+MBs6KUhh2Oz1Oi
AHOeI890pz3GAJZkvO3cHRGiSu7FF6OXyVyDjgf1+FWSx+kCBK4oquj0E/3aqgN0
NyyrDViGDqOLg5TiT6MfPfTZ8bIIGesAIGXFf6dPRq75IlztK0sQdZlhOFFCRPp6
XSYToPTklcZcu385MhjEQccgiejos05V73VZvUd0cV+RR4gGhg+kEMBqmcQSVTp4
jyUvQPVKguch5DcqUvvvQTHFOsezPmoHC9YHgKLwzc6qn7/DS96r4EO1knlBt/QV
ds91YQaM+N94OfmqJUyLLjyhymK7h7QPuHW/6CmII6PXrUzzUJNTdIFOVSCaDQiP
DI6jKz7fEWhTsDbEZrxtURDDsVLGfP+OhemMNRqz1S1TYx0svJPGqJbxtX22VQkD
cZNxxOwVJePVC1ycmUkp0hOEa3FdVaarE+HRzjwo9yon3Hwaux1QtSR5uyHVIVMj
3h9/HP8gA/ac2OprZ/nitScDnaihBMyiKZVWf19dDulmak7loKXF1HB7hU+kOVGw
YW+5UiYj8xgT64qXqbhNX1AtR2BsOoQkLn140F9sONXQJWW1lgNk0Ms6xBdyTdEG
0NXypZuhswUXiXA2y8l/whhoi0T5TBQKqh/kFN15t+G9aJ+h7IftfpnZ0vwfYWJI
sJIGjqY3hJZRAsfBeYwCUY/L2PBJuyH8jaiITev7Kl9XYc19J4ave3m74AtSpB6W
2foyfo81wnV0SvsA+sit1VhYjr9Po7O6o/lUca+OSCeOU6Blp0Cwl0JLOrbgExtX
fOC+kVMFZ84UoErMI3TVzT625tqssMmFk8Tj1//HsAcyROAm3+PNF7N/HHEriLqV
eQsviyoseLAolvjg4+hJH2ZHyHgXbmCJDfKxxUFucPRo+xTD9Z/TZwILP5L3DzEu
VXXJf5OHm/No74JSGLtgTwhgduaamf7vhGIZ1YxBAFg0SUN5LArB0XqZc7CXtgYD
yQaJsHaYCrBBP/gXsoaI4kBTvuSnVHcS4/9s32XerERnFHQhMkG28impmT6PjtDY
r56306gYCmXJQ5RhsXyCYXZbRrVYA6DSCzZck25RP71cjLy6SmSGczrenvN5OXUY
RfM4tNFhwq7iVYhh9tztheoE7NpJSzNd+7uzm97spbZl8pkzFW0gM6sRqt2TdZ0t
MfM8b1f7DCgouoFUrf1/cNWtU+m3beO6KZmPXOlhz0f3pls6feSF+JpdP6+MvYAb
bRwxT3JD7ZFCwfnSR5CFTQXRHnHzeo9yueGrXpHg1Rx+MqUemarzalBpZ8xDR4SU
EYcJPyhm/syzdyYjsqzfoN1wltcFGKMvdGcsbWnlcQ4GamcuTwjzlmr7Fz/BzuvO
ORcDEbhm0rif2fNF8x+kYZYBkE0PDcASNndnylmWg1XBN+o0RcVMZmwD+iWTCEbc
4HfjI26SGGY1j7JXkUndgUL5/eNtfS7ZjdoktO2+V/cYUwcCQeuuZ8VBqmB4Bt/U
8AfluZoDZvt0etthoZLPIbZ0dypat6Clnc9E/rcsKe27MPYpD+jsZDFH4KMswluj
ycqbsT5kEQaXkbzBkneFbUUqCxUkNsGI6JxSL1LDLGx/G2xbwfprh5G1lm5MhCna
qHcsFLTIqCSkK94jgR949xrzvoWeFA7ZOzmFeTafgfk1yFCSyWJGDFTNz0b6AvHS
YMbVzsXJ0GEIyQWAUBRj1xuj0Oz03YALSiYjZr2yqlw45pYYTfxgNrl8T28sqWsP
xpHlBXgWVLxrjDGfEgTQC8LJdvBsLMuHXjhv3KyvqaQtIbCv23TWOsBp7/2vckzG
GOv8189gXJ+nC1zsSVdxlqE7XfezenmS2qYM/rVKTQ4Fu0jp3yAgi+2mS/5BLt1Z
ac5vPXnSIMYU4XngDgrDUGe4e0ym5NS9U17yDzg3OZCRg5JI/uzv6QM5fLB+dS61
X2/dx1JbatbAeSIGjHCqx8CK+upkQL28HZM3nWHaadRxVzU/lc0LpxX8UrQFqn4e
9i125vojKxcTJsU1SV7umvvCd+R3q6zS9liTf2OhQyp796ApQ4o1LxgSTMYczm95
`protect END_PROTECTED
