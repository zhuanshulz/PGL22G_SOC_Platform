`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q2N5Z0A/YA4DYvz5SSd0DOB9G9Th66DrM413QJBkvNiF01T1/Q9uICybDtxQovg7
SRlXHp93g9glgNSZYIkHuOA6iofzpbLv686wKOq63mUGTJw8Vwo8+usI1EgGhiqP
WFI4PzpsC/Vbp1xdqodWKXHJntEBVPRxiSvWP1UKt/I2OD8beWmf307l8eYR2y0y
A1saGMwCwqAbnzT5vqHsHHHSg1CG68esVkfHOzl+pg4D9CtBCdwTLds/GIf/Lb0n
ak6YWJrELNCk31+qTMQTO384klGh/xkOX6UNPWXajJqLmm0qf2sUM5gGv7zBIfM6
2eM2MU3IMhEfA5J/frjVJ8I9trEOLzzgxqRt6hIFnCzIynecEm6nRrFbHte+/e9J
wC9OIzmI2vj+6KORmXZ0F32ZBR9yc4OdhOmJaQZSPL0DeQQ7HyvoKX8pqZq6ksTv
zLzX1CwsFVBPQdvO6n8Wf0t2MVrGJfJbFLVT+poKtm/ppsKyKix+H6FwaM/LP95N
tcG6GwzhgXmt1wm8dlsAnczTKuVpB0b4MEqO5d5LIG4=
`protect END_PROTECTED
