`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+EbK67dpz7IGpMZi3+AONEw9ozVdnZfBxtdf6SEc3ubKoKxyoXMn7rz0R2woL2RR
JL1V5veJznvo0xsQn47JMSHLpZaH3Zg+qppQ9rp2FHuxYCIzLW4+598mdbJ9Te4Q
iWf4x1XENHxR+JOPy04NJl6+rSqCokw8A63gFexnqdhFPeavWt4utCL7qFjdd/9d
peKzav9jz458MkaehNU3VEaG2uDhEoELvMKlM0nfBZBjN3YfRvAy/baB4zKHWtnl
QKMuYRVK3oPU6xAbn+ke4Ap9VREa+9V6SJERNFCDNZZb8bM8q0I9Ktp59G9Pl/Y7
xBSOBsYQNX8KODPL/j+FBl2Odzi4g3n1H7RAERylvoxBmoXUxCbnlEexyzZbjVd1
zXs7ySCrVhikLpz9bw4mQkXQmSdtkNPNTICP7YCaI+8/0zDPv0Hp6uGBN5SwELas
hTd9u1dGvI49QuH6Wt0DAc62yKb+vO/R4b9kzIauK3hmrLi5SXgSjpyRZES/o9W9
wYOJOKCSwB7Pp4fAgmzl7N9psXMc6vt42L3oGlY9CyfujULIwMF/OULm/pP60+Pr
jbQUqjrtPWlxXQwliHrVuD1oDsIpGrteKqmPApjRGbGFV041UB1K3Ven7ZQtp1mT
EmdfBpZH+Fqk55Ci2boIUc+TH/dMoEJcF3/v2F5XcElha0/FYBMyx8BB+BARZW6Z
6BrKtpBFHKnRJj3Gf9c4S45Ii/Jx0s7EJBRkqRJsZ/It9cwsJhpBfsm1kkooOhP9
IJiouSHO0olX4iG5EZKw7wjznAkWkwG/S8q/7Xu0/V0TO5Du7EMki4mEPWdhFNOu
qwf9Pr17Oj/Qip4VVWyfwb8yFsfBkse5Xc+pSBV3DvFqGd9nM2E2NTcUkbD7Njfh
+ETJKa+468n1zSe2adIqetrERBVYPe/ujassU/Dg/xRYnNSkIo6sYCnaeZFJqP8r
6FJawVHiSJkuGL5PON9B8H9X0Zlds/0XP5mvRr1S7BWXUVXyZStMZ62GmPaFv2BC
YqXd6Khtg09jvWrAAYuYztJNRShT/EK0yl9ifabBcGCVNv6qKSLlsD4C6PPhbibj
cjBhYO6ap6SnyprmjZu/9FdTcv7rk1MxW/j1daYotU8N53YRBu7Qlg9sSo2nvDiA
FjrIho1Azu7OANzD1g5t9b3oLDM2f5jYsH7kEsVZrvPolaU0teAtfjg+vbfqUjab
JxMsT91hPuBQu2xxTEwy5QTt5OJtthXpCIXG4kRsF5Nn8brD45O8iEOSysXmqDvz
YAS4XKBui+eYZGSwIX/AllfqEPnaRPokW8I9dsp8/WWcnqugQDcKGaHWMgL1XSDc
xgAsZyUKe121Ohai4BPaNGf+R3Zy0gmuOonZbjwjoWpnHI1D/OQrJviLo3UaANWs
cCBoFVDzzXifzHb2yh8a1YYtnSUSJGBF1n9TYzoPSXZFFY0Ks9FO7gPRd5cCfJZS
PnNS59xtlqJmhNKY4qSVmWOnufQDBIgvcf1bYSwY5F+Las+076Do8SukNcY7Zg61
Z7UHhqMkttbc81cxi9JcACWKLo33jdNSaczqjDumKuXVnDuBg597i1yJmPzfsTYc
bkF3F6lqmv4fwIUnMSfhGKwQ71xO0j5Q5FadHFYWWrMzwFUDu9yhaDQEQe5aNx+t
1kiQhu8RNbAHFM2a/M+HaDx7dQXmOFIyF7t6Ri5jKuxA2BnUZfpOOf1BkadeLO4r
G+35DFp7iCVuNxvJxFOxsD1/tTgUUSLLcUgQhqpLgt35qsaLocMpFS/xqXevRPJC
Qv3V895PFkVi1PST3VHivQ==
`protect END_PROTECTED
