`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MvR7poLPni1Ij/VuqxFQlZxXFVLCJH7DNwrUEaYVP55zNNq2+wTwyNtotAlbYail
2VhLjBJ8TiR3zrkFM8N07Pgi6chvhnBWD9RecjHlMqUu23cNTjKCtyxYzkQJ0z7y
DCG6KRH+egIpJyxMuijrWuOAfoP87aMpHpcuvDaF3DiSdr4CJCsJ2nF0WfzZb7Cc
ftlhMHzhDiZ2urPWjfIjnnaZR1KBOt87VqMMk8zEc3pYiQJmDxs4EtnODV+hB6kx
MW/tXDGMhotp41FrJFdzUnDw8nYWSq22M+w4XQk+Ja8BrXz+tewolxYWefkKrL3n
4MHYvo0JIWnynPtiGRaxp1jkkLi/XjDiwveVN87nAUix4QebioJaiIpNlu+56Hki
lqnKBHf7a9MAf6pmnfnoGLokhsAPIfkZt4RLI7Rm5cNDuz5e1+GKjsdRDSrWvJsl
lPE2VrR+OSSm3rA67aFAGJGiXgoWdWu4bVC46tpFcTHKOgJ8X6T6xzis9pkRZGsD
tm+MKHxheynaD98Wf9zIhw==
`protect END_PROTECTED
