`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vxRSgYHWZwHzug3m0M4HAwTc7fE0+9ft03cT14h3vU9zMc5iq6AE4++k2qTXAgBp
lLZaZl1VIFA9IjoqzQgKcZbn2hE3bRDyIGtxHiCB/0eeUj2/93bznlxugJoOLZr0
zEppdgzNQ+00VV7EbRXzIN0Z7wDGSxcDi31B0zIL3zi4+P6c7bX2YiktEsHdJ6jV
34qJt706ORxOaYLMPNsVElq7xkZXE9qqiKKAs3EAzsGAmu6sEnhngaipY1Q7PCGK
xh53tQc/7jbdTaCUXbTwe9zaA5jG5ATCOxYd0223hp1ytpoCbW/GqhaubKcVw8kG
F3rzEuRQ058/cHkdap9X0crOPBhtz3ewS5w40Fr72abn4viSwt2DM/EfM3ybmFiU
76VSbfiA/LjFhB8r0QMSG67ajLo9oZtsXtAl4/hbpwh9I8RsMaGabiB2djmeekQ0
ngj4LznMZXvqAEEfRbEIx+LZ5TIBoOQLGefHkvPVLmWBs/dMA2FkVetgfiCsH3/h
uYqBqJveJBdrazsuTpiqymXYnJGvrEyFC6VkajE7PcWrpCnHu814DIAMCxbyO8z/
cEIVPqDHAZTdlx/Wl+N+w7nDKpIhjr14ig6ok7f8LZzsZ2OsEsQ6iXeBnmrU0XZ2
KtKzsiD+rXcAsJjA0m7JQX3cDCx9r4bY9cg+mv6p/VSXu0N1Yvb1M9YIPH+S7N7N
2edaRJbLgm2LStOrIEutXaDOg/G1/zMpNnIx4IYhDGiQrEvIlEfDP8MAUILhld4G
udAiaXx5lgl5fRbht+XB098I4iL9qmV+79jQInqFaYKj0nEsnjBSv1/GnXw9VnSc
wCw1VD+O5mBj4kH9vAM3mDsj+KXyw7PXbtQIga6/Ndz3FygwaXJtFbPhs7iK8Ug4
IklKscEMXY2EDXEJ8Ui78+vT369/swPPtvbZ/3E71R53g1Nz2GNvZ3s3EUVMK1lZ
Dr+DJmfEQctCZ+Wzv2T2lprCFcyURW70ncXMIUu4y4eiiUpRNzjCrCnHsLIGaXrO
p1QhlmyEfDs4X8CdRm3nheGaR/lOVZ8BIO7JqIF5hXvzkK7tuILr/XNzQoILY045
Ba9ehf+P3BQSFGrqi/QjKlJb2BNeX0IkRTfsRZZjE3ktwTJrUHXXV+GklNs1utOF
C16e3g7SiOwjZZZhHyxlgCY+ZBpcEQMjppYoEhssY/Temt8BN4YxYgOu9oKYvoAr
p1jQSX3HN8eKKTXaQ79MskhgAYMom/eH6YritgJWCnu84cOykeUM5VYQ9ri/Y+Qv
bCjLhWYRWJvHMAloq3OqCQ3UG6AVxS8K2HKLCl6rUcFwmAqNTgomq/qk6fJP7DcJ
LUjU/Vh1lrIrzRohCPN0+PU4d5UxwJbXVWDHcWRplgz/erii2UDBUbBv5hDql7i4
iDgkjC8+1XMcoH4gkh4hOLMrPwx7thAUNUN72RToq6cXoCzEv/ThpmihOWfpOv6f
HgqoCMpL59p3AGYdDcJM+vSFzsylYA1220dgpJZ2EQAByt7/7ypPXfOtuRFh8bNR
ol1gCg+l1w1Z9+qXtqPwYVu3czgj/Ch9sUeOrX0DaQhE78AthpSVNumADVUsWwMD
VbqDMJgyBmSPGIBo3dTApajZcIADQiykmKv0bp56NKCTDng+zRYbSiS9gzKiJ9Wj
KqE93V5y+LpAATEqYhe3+wIPhTWcPXnYcJhcCelTlWBUwYSXUFj9bGSvaZo7OHnj
Y9UMbG5EzDd68mNqlM3FQLcpjFYcf0EzpXODXFLhNqMcllqhmtsRsMoF/M5mxI7+
WpzfJgU0O+vH+ZCC6cWUu33anEPhZoVrCFDlBEBGnLlhc2FKXHW6z0aKztKF5ckU
vI/tuD9UrwHuzBe6dEUAZZQT7g2tY7ibfLTsmv42emKXYzH4kSoa+YxGBGo+IgCR
0RhcCkjzkBQBg0KwrGJqPM7zNdljcDjqEMj0PHTRUztrl3VbZH1Aj3gYbAEXdHFa
z7Peg88lhERmNZ6BLdqN7e+Q8Mp2wuLgCa65wU6UVJLH75WjtI0ZA1pmarHbCyFf
J6fdUa5baTxDncvKHhvuYBDPBK5wf913efp3U4YDcbV/8nZChFjWZUdni3OKfSoY
06qLqfLyuipe8qXHBJEH4izqhaox1qlqWL+zts+VeMJC+Y0CWFOxx8OWvdvm6lkf
nzTGrjycysBJlVtDKWgbyZJmXU+tv6hwpiYW/3AgAaYo0eD9GlzbsFt/Z+i6JwLn
LX5kkdwkNCsaDhND6PmXcGFNSMIWKLW5fjt7s1mwoHTol1GRJFbIU4O/9E5RTGW8
CbKTmRs10zQ+/mSTNmnFJe3NsP07WHuC6H8dwxyahyzzp2Tg2SIfQs2X3QqQwe0E
3nntiKuHXQbqxOPfEgNJF4HvzXkndNRMKATB/H1uCnlskXG0App3zcxbhGMeqzW+
urVAOwGuc30kQ6P7pEX9nubwU/KCQUVyVTXlKhEJByQKDisl2dRCMOW60yKzzZrX
aU5uAKit5+3GQa0hm1GXkSD3SL1mXgAGpj8pMkMzfUl4D0SQ+cWi0rGk8c8UWx4w
X5lNcA3aRiQfpwtanDvYplAmWfabSoPBAVtTl/CD8yXRsfqx3LXV/cg8nyQdENPz
nwjIQLaQOSbzwV+dmE4a5LliO4HTYI/jdXrIHt+HxUMCIo6hrNRJnITksEfFE0ZQ
KvZcUtuNsXJhhYhYFIGUWkSjU7UT0mW40UTkqfC/jA2pSAQrfvnKbWByYC2JL0HZ
76Sek/iy8WATVTC408aCSR/zyav4ir7Md4Wy8ELeQiagkBtzqyylzPNUrH6/72z/
p9IWNA4k4SUTZk9ud9edqzfobszfIM2KNpNmpkZLG8pnS7IFtXxf0LifNAxFC7q+
Di8cMA0ZKJIQ13UjrGcthsbOE29vldny3OT07baAmT2ZfYqJxMfy6WT3ViZl3SsJ
X2Roc2LEXy9GB8Nxpcu6PUHtppmUY5C4jLH7SzfgT65MhwvnSdbQjnWHBclzRFc1
DQC4F0HqNDpBpVocp3u51pQwDNgCr37RIidp8NNobXyzCA5j0pj2IH9QIsdr3kjJ
TNWDnxpPzn+4xEzRdTqgdGne+lZQHEJkEX7DzgKoU4O/sHTEIzUDtEllQ1rD9g+A
/ZGXIXdqVhmIYEaMunvfi38IOwsGsxh06J1jHcRgB88jen9a46fbBsx68NoevMup
SNmsDlsvJecB40NA2bC9pvN6fPRsopaSkntobVVaVMm33osUBtuzJPi8oTPdogDW
TMw306imuNzH3D0H5N4BH6ogl6DckkG0FiIlfKYipuGOGx/u2ErQ9Tru8sPLlhV+
`protect END_PROTECTED
