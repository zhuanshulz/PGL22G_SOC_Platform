`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hS0LyU3p4PTrzoirdygTmnHqSArXBb4KmPaa2ZMUKfLQ3qxquQBd4mAjAHSxQaLG
DQJrlIRyD0wzkbH9HXzHvfSjzVJnqw8R/BCFJ0TmIBfctnEYZcGttp5c9AbdhcK4
26hHMYL/QnnFoGfnhfY4N8UaoL2bnDP7r7Gn2vam63grdMeiKcFmDcvhpfr+k7li
rCbtCR9jomA06j1Vf+o8T5nlWHeVgXyoeHm/UdFlDkrFgM/FddnRVDyBw+I5DmCi
z8afBRGg3JEMFmjwkKdb6O+wyMLip406AvzsEfHEdSFB54iF9uiUqiJqXhHNNMew
560/Irl1i/jOybEbTs1PiqXyTWShrtUVnLlLDI3WZobzdiWAxB0oEd1jOUDrfgUU
H1IyFN81icStcKCRFcGkBo+eFOobkOH61toJswCSHjmz2m9Pxbf/+oJ2vCE/agny
4MG7eNVrDliiug0CH3uLSrTMxHE3P7HRAQw9xP1Up8+ckex5JBgJtp+KPiN57WhN
mIWOD3f6CiNSul+pcU+YOFyXtbo2RUTsDR2hm0SINZY=
`protect END_PROTECTED
