`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y+Re4i8R70aywJRyUakvILmwgzWlB1bktzkjYUXcVULoLbMHrzB4oyZbKqSwcCoD
ltZ+nWa9JrS+C9qrSs1dQ9OorBJPTb3i/og9UB2dypme6sX57jOBXTEhIJ1yUF+Z
PJAEHAn4qxRo/f+ldEoGILjChEVrn5Dim2AGJB/m92aacOzTQdsDdHt2pmBo1kNQ
VyDIpToX8HNXnNYq+G1ouK4xZUdshH5J/3yNh4zpb4wozOdwGJ9E+TlTz+/Hitew
hIdgUn0j4bDLQ/h8oA1ZHSPcZd6/G5IBOxFbHArLAv/BRtXAjZpyRsWShR4wfC8D
mveyE3oGmA1kP62mXh5kPlZXJ7ds5LYEX7auoBRaee5sFTAqakTobYtYd87isQmd
0XcnpQ7nZuKuzOPhaweq5ukhKgI8wLetfg0Y6LYoMaO9GoeXbb8GHQA29xZv8/zs
8R1E2QXcAP9QZIY/F8R8dsjMeUWAltQS9t9HpN5vlHgto30A/XFMFfYURYG1+Eja
+y5T3W8PzOEdgHGICgbVN5kE2hzCmJY1I2FC6dQI4S7eiwc+0JSpu7464QzUyuGN
jszbGWH+P8unnO/19OVzq72aTE92exPEA7xIGnyyQmVNdWXfC+dmTY3groDny0qI
rXkyEpmZrlSFXoDfMNS3/0FPwpzzTILTDGUvGXKfQuEtxnsVY1HLMd0+sGaZBALk
C/yadC4T72Zjy15xlWzlLlWtYbHZ9LDcTL8XqkSCNex5fVMnJEARJTdl8A815fbX
aBjmgIFkhA4D9jT/8bYi20lKIC9Hzs0/9xHxi+Dq8pmMCcv/VuE82ehebFObR+x7
e+wvsC3Q67nGO2HXxav9QAukxyUhg9qhySZD5eF+1rYpIojaje2uBvx6wpzaMXCR
PyP3N0lmyg+n6aRy6zHxw/xJlUf58uTG8X4F3X8pX3lNuK3A0HnMNHw23QWKXHSI
i8k7pAkLWMk1CRo6UCneAD8JrCSOGN/X1lp8wpSqZhP8G4/dJOZQRmX8z9cZoP2p
JnnaycCaXCq110qIk/2eQntRNDTrmbTwquZdyRJeMyh3i7EpMs2y0Da/cv8FtPg6
rGkXNgEae4e5atIdjyxaTAqaSsQgLRFMlKalWeLCCvCjjvpKrI42f5L31/moOY5g
hIFpVt1yMYIiplE6HGUiVPGPdvS7lstuyxhAjUn8RhLJj+efQvFdqXr+470FvaC4
AchaWwqX54I1I08dJJQIg7u7MTBNym0pJdi+vSzQzQ2tq2t4rdvM6gi5bc9jx3N+
x2vqezuicfyfEs5ZDprg5htE4hlpnAyzScrtDT18dNxBHLsNBNqbkLkFy+ttxOr9
NzPSYiRcSgJKc8ZnlHhvwDHFMmVQFjBceM2MKxm5SvveOkOV175K3iqP1lODGcLJ
dXdypWt0f0SjOeJKnrSWmezVEyX26q3kPKJ53GTxyRLLvBKsHshGq3QAimj6dUBv
BPjo6TPMogSmA1zk2oDPTwxvvRpdToNeZoU1i0BS228sDpY18lZS58yDE/f2ryuS
gcHbyEWbLdBYk8Fe+GMOd7muaUH4oJXKlxrwZUJ88u2A7FkLArRlBU4nDH1QHcmN
jCXHoTKc5LfXOAg0D0BRs0Iim23mihdD1m/oARGYRsft7YTlLbGl81Q9YTG7K0ze
RZi5KLwhaM2B8Be14uBE/Zvx5Ea4eOkSQTxRbuEFWxg1IO9OlX0NWie09UMIGDZO
7ksAT9/UdCEIJ4CmDFuwWyjp1/iytSfgJ/3JDsGP2oqPIpfS5tp8E1URSzLkvKJo
PD19vJMdsGK96ZDu3Gr6p0j0+5M0gOsGhQ+20fhdkP73WC6wlVkdvpvi0sQmctyT
H/3ie3oWqhzjWSmNhO4+BK0xMvKNizWgJcPDf2/dPbthdIjzuz1uExKvQEaNDIRz
v+ylKXZFejh6VxnmXwODggk8NXwI81pdy0oaPxS085YjqQQJOFjSG4ikJyWvyWph
f11XdtLzCSJxxMJhl8/DalS9EgyPBAObAQRdhFvaVpb83hlw66C5E/yyPWpKW3P0
kRh0DC9MxVf9CxCu87VEBnjpmm5p6rR2s5Gwxi8gDZmvetUvZM/85Ki2VHEWnoN5
lHknCWereohCQ9SrD1bIVwkDZay3KzJV+JS5YcECWP7pOeNiynoqvb7mHodkworE
lW0cik8/Tc+sBwpIFOZnt4ztLt6rLxKjl+8j/fVRrENyYTFCrati6SKa8Zlb2WGC
URNWuSzZdQFTHFtFLBMa2w7VBfXhGUcEzbjdwFadLa2QfRW97D4SKY4c6oNaFLuj
0jS9emnqiw2lMDRoDP9zTZNvzXG7ij7YoIn4lM7NpdbNtI4XK3Sbb2iO7EongVZm
3j29jL18H0zuxYmHDFZk2wc3F2JavCobGL5FbHSzVyUn1dNVtB89siEmTJHvqdyn
njP1qSk/dL8xalNvS5nlJZ2R7sb6bHMlgsLwQAPL3wQFoMbClOW29acZzns72Peq
40vs3P+nQSH4LeIeYTEFo0t0F8OnVYr8hiNZ+A9dK08D3f3MDNW2GEVuAfI4+Wv8
gHQpZbf+3w1ytpzXNBgoP/NbUoCRSs8w8xry5FkuxYa84GP+xvaRunO0IwIx3NBi
y90EcVoqdqywSHNbjg7Gvk6iz6zaQNO6jjQlzOkrZhakKJ2cP7F4U1Qjsrsza+KN
zVJ7PPCAKW7pA78zZOT8UolEd4pVQJCXxNXnlAEIuf3pRmKM+8luIRlimXWpBUN6
Ii7JDdW+UVTXtL28APsQPvvgd+TVEDY0xiclKCDrBUyf0RjbvYxIrgHyA99cswQK
JYZSFyJk14vx2T7VXV4CfhDajWnNYFDfs6ukoIrOsMG/JBlF3cM15TnSzZnh/f6c
ZTUazITvWG72bo3eGPy9/LD6JUo+/HKlge9sP9Ioobti+Bj9uOy0mUhvjlVS6b91
pIMp9cx7iN9bFSMwH+jWMnxIFag2XSG3dTo73qoQHnvYuXSvuEpNGQdqOdLFUlqv
ibkZMZZOJA8fcRdR4FxgSzjdgtE6Ejt9p1LZ0RNp82bjZfvum9gdY4H31McyGMIK
T8sozB0AvLHXLFk84VEsh4qime0zuhZFXsxxUiR4e51tDYV0pRYDABIPpVszq06q
Hxz/2LcWRL7HqPgHvyvbRyK5VxTBMxSSTgLPmQcUbHdR+oc5jOtN9PcJp9wYexIl
kXw3zwEvbkUdVjXPBXBgZf0IESu8I1TaUrCvAjX8845THG+/ba1BMbDmAw4X/CJ9
AQfDW9im1/m9gRjwVLd3ZcF8a7FDr3z3hYRVrx97KofoitNGwv99ijaps5RX4Aw1
gC0xQo2Peoktsqw0142Z69HKkFKu7/NcE2FJHRVKxZMlFRx4xFdLkpCItIqNxvSn
rQxZPY9Px+X7uvsVEwjwKvWui2wZ2Z4j3rplYNqBoHox7tMcsRTRZFSNS1aXCVst
aV7EzEKKFq8lztrioOvAwVvST/RcFeoRzKy8cifGA97TznN9laFErTkOw8JZYSvo
Ghchi5m5FEbi43T+KQKCKYIM65OatgxOUOYgemqHbFI=
`protect END_PROTECTED
