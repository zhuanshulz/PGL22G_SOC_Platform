`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZpzvAvcEf8NEaGOaYw8P9OYcPqm1paBncZ2RWJGgDFHwAv8RNjaNs1eaFIshJpmP
4HhIvcaS1GxjnwNOy4Il8xA28EEOSCbypFLqCpGhWvgF3hQmOAbgffuZrhMxb/3t
96ZCbbCubQW/0jzbnHQpzDYlf4EThkKMJmnuiFsyZopP6q8PdZIDbgBGO7qxU1zj
wNLEbC9yGtd1TI/6U1eYZf0trmG/OvRwO3FzNuk9SaMhj24V3i6mbhTEXrTTS9a1
FjfqzNlqOl6TEypPIbxDbGmKLlqHg0kmWk4ZCP3YourVNnjbz96Dyg1FxaEE4aQX
VVhUPEcoKTFjndJaY909jPmqwsP2dGM1CQgve+WuKpWt4hv5yj+PDCRwZ+/P2CbJ
Fo+51xZBd5sxm3Zz3Iou54sInIjqk3lfWSZc7mXAwm/+4ZK3asARPWLXTwlsWO4z
e6c2HrzLK9+q4FeIABMUro3N0+xFqLqBktGLRi3/+PbX3AJBFnIlBlnZL/KRzLKR
EGzKYORrBkUktiptqpMTH/pxQwZhXNXohWh3DWhov4K+vklfygrUwp1Wq3oix603
Nf50Kf8FKm5fLLfMk+Hjyg==
`protect END_PROTECTED
