`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f/w0ES9S61VyflBaEamU0ICYG0alr37oKGH7zWUaz5ayj7JhqIl2QIO8M98tb+Ch
HZH/mCyn6syHb5uule4GxLamRuPyhBfcysuPPGyW7qb01nPrAln16z09qPxKg1eS
OVG4MBGL2AmeZH6YYAJvi8pktFMaxlyzDHnDtrNVSRShfZYPFgCi+VRQlOLqHAxA
Gfx3WYYzKq55rXmD1vScySWmNaAnr6e8z7bsd5+W5wpCWcOKONxwlGEt6EYR6QHJ
qus+RV51A4Y7f2728IDyprj3T7vY6dAFf+1Nrjjgg0RVpSvaFxCUrwzlLsanDwvQ
CvxXY3cXUu/xL1bGhmzs5a0OkPraw9H95Bl5K7cSqzEZ516c7DRgEQVotPxMlI0H
nVHFYTpdNZjH/MFz1/BZTLn5hey9v/gBRpVornP4NeSvB2AV9ufa15I6yBSNaltB
AIC/5DOPvvIlG/xuggxpe4K1Vb5vl7SVOyzG8hbwjzV2lL8ePfQ+mH2riLSI2jKb
WyyBuOTjYaAMMbdNXPTKukbAx9WnU/SRRFRorkl/FG2AG8l7M5eWbp3tXyKLkCE3
uivVYVwPTiA8behy7pIl0NScv+Ln4JNNscrLZEA5xWkcFvzmkBQMtItaQ+3NKMT9
XZAMkKZuffOsZPZhlUo33z67JOOjsTc44a9jwEToTJHCPXQ9c2mFQGNQpZLqFnea
b39tqf55THK1tDryOT1pjDsP2znie0igKh8nsliBe4oB2g9GUzDZD38F5fmxhRRr
6ATUJP0MA9vpC1RNApJcwR2dTbRdiu0LYwGf+M0pWdGSX4bSxgJboKmEiB5MHzPP
V7zHk8iFxrg+8zadHQCd4M15JNUvGf1rpd6kBaiWPsEUVVBnNyTD9znuGPyewtc0
v3R7h1TN0Re27+v5lUSPyPK7EC7xELsfIkgksx7ZLzxLblrqLralxdmOPqY5h5tM
J7U/WvkkmldAhsNXngiQBvaIKx929Bw2yhDpeLh6oPcDg712L0w9nuNRHMhk9vhr
AtXhmZbsJn88JIIm3tYVG5kvsKSZjIKcic5ZAsFOGTzF0YLm8AcRdGqHVhHA4dEo
Tkp/5dyG1WGsOVc2xuzce4lBYFLDFA6J9OZd2ujQu3KLZEVH9KedcrODJGRG9f1A
m01XcOPwOTMugLQuJb1rtE8l9LBPu/ALBXE7QvtPUXHies2m6QHCGxyRMgMhgKGA
al0cgRiPK5TAAUbjzE6c2dfSZh/cFPFtSpuuHqYONXfFNbh5g86U5dKtddxq94X2
f8bl2qcYnpss6SN+Ov0ZWTiEVlvyef0oElvTrMZuMnnvHWwWM6UOb+z8+gvKPtHK
lehovw/z3cXEJDJ3EBdl6Ff93aPqzA4ghRN5hX+QaisyMHOfQSDppYpb9LDzKDo7
Hq97U++J3pVSLGQebVfRt7IvoGF1Z0gSYTeQhE5+Q/wT0RXfghrUBAzAteHid8Oh
Pan2doXunVS0MxMctaUsTl3+Motx1eynFydg8mqvAN/vjJE/xVvKSJBYaR8m8o+U
07RLYECnpv2iq/P3IEShJV94O5d0lghlfHHyRE4pAKk/8kFISI6C7/ZmhpXsdP9F
IEw81tYg71mO4oFEdykcO3op/t6ERV/4HgZzIU2Wk9ttkZNm7/aLiOxLzFYe3YMB
J5AF/8SCnw38V6XKXCshqDhcwc4a3v0EzofLLqc1ejr4phRm/HontNd/6btnq5as
R0hVgLMrDP+5mk4r1kAfVfIpbvwdyM3r8ZVLl7/SN/J4k0DgcesXMeF/zw4XUdc1
3vcxfF2yYK0txyJ71+A+4rB0om3tXTkUSnu4+CYFETK7JZ48bNYRkSDWf4Z2bJ7t
BQFV+9utA0vHCzPXl9rvOZW+JmBYBsp/fIzoCXJjCFeJpHvJOCU/0/UCqg2xSmjC
dA4h3NKIljX/Bf5vU2NP21G0pKnAqT/yzBPuuIfQa63ydSoPA3lzaDX90WB+B4ra
NW4Csl2dfkyuu29R7rPpehUTpb3gLbcJhPsSOwqZC1tcKfIQdZIpRuCqnNcIdMnK
SfdUbXYGRXeWwfIYyvCsLNX+y7Vel+lw8G/4WNdlb0ik31yoYtfjDA85jkW+rY7/
GVeAmXnyIyN4whaSW65EBSByfSFrIWJHe1E4lAh3cuYIN906NIUhMOBfV0Llcuy5
afXL+FiHAQRm0DwzF8+oRnbXKq7IKFJ7Je7RA4loAkK+mgnxdAfUabNQH5DP6ZwP
Utf1QUJfgpefVRHjb3JRZOShflpm3VkjPthVGv2026qgK6dU3fTeEjHIOlUjNMGO
eC/0OkgOobiHCRouWYJYZzBSFRNGlR5id3vmjqrX4aQkW5axjY4Mmhx9TMtdk+hy
EIoa8OUeMlsGBV0YNVGTFbPfhO1n5g2QhF11B5mBAuPVL9YviCa+tiNvMzDmgxtg
S8g+gaN0FjIThlT4QZuEr7NGEowosah8Y22UupN+uw51J1v9j63yCzarsSI3Mgkr
/5rvlfJoQJxTPE5K8uMNHC/HTAATzIXdf2FqUnzZ2tq9yqSYKOP49N5WxkZHOL4x
rSWJJYTj63SO5DKhcgPcNHgrTu5SsKpSt5OpCJR02hNnCpF0HN7djJrznboqS/ic
s87t4Y0SkbG+mwx/8Z5tcJDslxSvyv4cqxCPM64x230TM/6onWWYA0Kd5411cGUM
pJfPWFH7GnH+plM/TKgHvfva0RWPafv5tgXym8jp3w3w0oovMlrL3Cii29g6f7wI
VoRPtrLLCsmsri+7hYG9X3mRCHGx/WMPYamnWuv6HrBGcUdfxSW/nbiXRtQIJ4Yx
1bTOU3Wk8bOq9orWqcruSGW7M0ZXLZSB0nIXNhPloysiedX87xlhVRGanGYb+j+Q
pNsBEJvusP2Tg9i4LwGOjhMklZedtxm4XEijWH9CGPWzc/D94fxMFUARe8OAZ7/n
FV18eVtx68UqpFjPvTJlUVKhF5EAqXV2Ln5M9BWf480ESwJl8pcLRw6IzgsBAw+k
0MHGxkbsy8sOZNXLHu5aqmo7Lwk2tyYs5SFT/re6d+OETi4LfC+lncIWxZnVbcQn
4+fylBdKYfe3jLjM1f2AMWZbuqW8IiKVVkHUExloR3/W4F4Y2+SxIwQcIkXR9Q9H
6IsgQ/jiBzWNFHRC8JJPrMyzx4Kp79KU7I6sdVL1tobcFyvzZMRUNWkz8gOk5Gg9
x0znqsgMDoJmSKNNzZTISocpJ0lPaPcbkgyi6s5XgOCvyDC+9mtf5VsUTWp1JUY2
e6BD+BFE2sPSpsVFwblaQyUzrJuhlESwZDqEd3oef4yAQQRzBJezLi61JlFB8Sti
OaI3L7N925RJjWcG1iCNpngQEhjPR5Ty7lm3Xne5ZXHCPYArnWistjC7UH8R5vy6
6kqDZZsF85BeHdnLuQtt54HO6wGnH7O+rwyzwMPSEwbS17TPSEkIQEaryekuNiAN
/fETWljV8Uub1gweHZgOCt2ilEfbMsmc8sd8V6oSGooDYyJKwF27yFUhMkduL3hu
MTPX4inGHTc7k5T0BAoZU3kX/QKG0OMtKLDdaIUppIJkUwFxDIltquFbMc/M7Chi
Tbx7E63T0fblU+yf9+tPZoOLSD3rBn/lLlqiQ+ZbpPQEQ/Jo8628NAyjDMvoIZh9
8E9NtTst7ESySlwfWc7H19lyCplehJYsuXk9k3GR8ZfFba4N/mThGeiyTdf/n7fY
oe/O8BGZSweyV4cyOdJs+OmIrIE6JL7Lk6YKTp+i4KCD62eoAeSjny/K8HHOyAdz
9zwBIlgNuWihPVeU+KbIsLDOp0VuUims8YhhNUKgsiim8GtXql4yd98kA5tEnFXm
3FKG/BZDGQ3sxwXOm6iQYmGV2uYlRvlokO9qB62RV7fOECC9JPwshAsowUfNmJ8c
KFmCjq5luR6Mm4S3qRVJI0I0iLumvM5VdyKBhjI+yw+ASmpw56GDDVxpGxzbORZS
1j2V6lYdeGmDO1Fwz97a4sTtly0GL48b2x7vGKqk/f6BkpsrXRZpSHGd1p4kD4Zy
g8x34mOKaCzhf2qb8mnSB0Am9F0MhvqxBJRWChu7C/xomDxx/1r16KvbL3OJgtu3
yBn4k3/1d5wXj4JAV2pZwRxKjMNaXHKN29Egn1glvFVsI5yYg+asXYbh0H8Ue6fO
Z/A38FIAOB6jZnzeDao7jkn9GxRAXkeXbL0iwymdEnimXz4GySvn7DSY+Z0Xpvdf
sYJAl50HccN9+H2zIekKTP+f8oKKZ4yVtDfXWKK7vavbb5CMkuJAzxmEEbjPMfIQ
BK1qxSmX5bf1fJ+SnkKv9yfzmDry6ILujHIOiLfehY8r8BgmfoyRBAxM88M0HTul
lnY67eCrshKE09Hnnuf1YAABGMizoEOqAolIpqOSGEAFOfrIUrsm7Lgfbz7QQyBv
LNesKQJYCaVUzqCqikx34t/03ABd0jQQVIhADuv2zRHh6SSjjtAf1q7JDM8aAf57
BvYWG++y7O0tqoPTomuJyjAv4HxjFBNy2eXwbGvtywjRRG/pSKF6icbfU1/B14VQ
RzLOyLMDGczn+wA/q05B5EzCeX0ZZIT730FsN3cTc0FnDJ9Kzn7WFvU9x09/3gyf
VqcoRc2eSNaKoXwsSltjlK6XTQv/KVnbq0WUgB41mHAU24YGKpl+jNU7Hf3B63g3
UAvjG31rR9FOuxDXztjT5uB45r6qCI/ud+K9psBLcYIHPkyoyba0KntyqsKpI3hf
qxkivufdu887Q1conTN43rHtnefo8Da0aSKXsdVKYMcPyTKImBMbiBSDReAi7243
v4C2XVn70iDSRoJ5odMmYVVOQu5vzD/ket6sKiBpwZmR53R4iPSjDNljbA+s8CMp
EGAiBCCxXuFMFVrxpf6+5CfPs25pgIgHbllwupSK5ztj3ZEYP7DddYH/6/vi/jjK
iygWFjat00xWcXtqb4mFU88iztDv5D0htdNaiD8FJ09gZlMJcijyG8xi4BHsU+3X
rDnwOnfkzaGC4YsgcNxqMYslPM9tR8yeifyZdAoqh+LuDg/bdeR06R1bDO6AXgHX
LYL7T09765JtaQ3rYD8JCd1+r3zeXfiMhDLwFWO55ov/C2XAWe0XrAZjDCL9wY4b
0Q8sjpEDEngH7/JwvdywVYMMrSP2yfMG15EzHcjIqMRMnhyrczO21gzUbMXDcBnb
543LwUQLCLKcqgRloJser1HAyZAkgji+XKvcSvozo+yYkMFpwScbfClHgLNiO5Zv
/wNS2CnYlYJ0WjLi87ijOqLrRMLU9Xv0V+g29ZPE6fh878vPaSRosvBcY7kJD9cK
FtLOhzGuDVQofvWphjdaXtLZ2ILJ1dS5Xz7LUZjo9NARG3OByPZtrzpFWzolODUT
TYyhpT54NMW2IEWZ5kUV5zkt9npRp5sm3MWaai+lJyFaSEZp5ad4mHGhGB8LWfax
CHyUSsxQuli+SeP9dbEo493P4AavySWkQCsYqUQn2PzEGlUVGd0z8q1+6qQ8rj7I
kCCnEfoDvvDOp1ouiEGY33/pqH72o59+Qur14Rf2q7SrC5nJjPqCqjleY1+g73nF
r8N3qLjdSH5phYFbjF0kddRu7lnlo4e8Lvs2RsO3KYw+jz0w5dBxlBCQ97eOL/FY
xqnq6sKqhG1optrlPC/wpt2voNZtf0pfo8zqAN88s0g3CyZBZvh23fCt9n0S1IIP
LoRnIhYeDAaJwVRRPr/mjQ5aF0/YgbcXZw9XTL3tvo0p/mugTWa5U4m2zE0w1Bqd
r8l+qv4vAJK8UXux1pGk9NA2ZhD2CFAZzQ7j+J6iBXWzmoyZcg7BA+FohBjCdjCa
yRemwhERbq63KFCoN0kkbob7CAvVZK5eK86GFM30HwIPiJ0Al01V4r5RXCUM5d2S
L8nlT5obxhtlEngkcG8KKQP59eA9heTLsPJTov5bc95EhKtqIzTV7XG7s7Fh8LER
naO1gURKNKhUWoi2G+9F4X6IyAMGatcwQpBeddDMUyFLDXL+yAr1Y0walG25yRhV
QACwssJNg5bH3hze3wlnRImfwm9H4xptLxsmlL35StaOC2B8SO2nExWTV0VfeluB
KEvL6x80soKPHo+rf+93vwo3iDmm7CeytPFXf8eJDTwi611JuvhlFVpRiPVVBEJQ
DRV17oOR3UXpqd+0hx6EY00u/SHFvdFdnsB0CzuqhztUbdRDGp8gznXf/zGToMMG
gBGVJ+oAFCf0y8YuFGVhWvhJ5t7MD8EnHU2xlsFIvsdOybr/MJMMCM1TUKEInJfI
MMYnp7lW2l0+kgpmcOejHjMojDgCjIEV8OPRvNouZmFaZY19G4CK0+kgy8LSb8Kr
g0TKbwi1glGSGhQCCytXo70UZEm8INyfwRccVR6rjgsmiUgZl1NEM2axnT0myn9l
MAYcPxZB+V6sSz2v0KGOLQtchgG3cHpwy03Hb/61GqpPCtNHk5ttPrua+UvulYyb
pQjSiz6FqXjuD/McEQ47/gFvBk0pCSubMqwiZ5uZzr1qXkETsJp01xWCrOeOSOwW
GthcwJlGqsOyCwjf66aoBeFbUcfgF0EXhump50gP4DN09UsVv74msiPIONE/4sqE
Ai9yvOteNVLLqosq4Xcg6LInx8DdI2vkqCd1900aL27UMESKSbXsQIJKRv+DFiKs
+M7p6j78QO6duS/K7uSZ3ZIJclWOBe7onbw1LjZ6kZVyxHqrJ0iXwEdnSEgrOyvc
0fB5MyC/a6VXklilhV2tqJPuR0NyBS5JP6fGaohcZm5wRjQHTurmPFD81IMm7DtE
Zy0b2rvL0tPslBGcJ/qDMh9IPWW2nn6GZzyX5SOd1ke9rFVGplKMQKruo/kCuYg4
4mZp/8k9UycyxtqGNwpgUFQYHe/RtZl1q+uFan139zhW09SjFADG//C2pT3upgvE
4+ULTjklV0j+p1+c+iiWCoB4g9fEd8DG9SiS/IoZKQgvr7/XgYf2/QwB1X5F/6Kx
UsGXm/l0kEmKGEnqSimz4sddwvrrnahANQtMSuBzOV0FKLLMTwagEA6wu4FHb+bi
+Axh2wKxI9q50kR+pZZJDsaUE8m91/jDT3sxO8uw63WauLwU8WQc/bEgthN0OxG2
cHzNE/Rd4FNmFoAuVNxdA1l71wFnFg44EMs5CNi1Rs0+l5pTnBkijMYa15ASyJ1C
MfgEpuEkqQia4fZcC+Xkp9Chs51HiRKPZAUD4DhyTxEEDtduvbXMpn5mIgGjjXVP
ShbL9PsQpVbzoGErdfoU9A7ofsNF+qdsBHrhwcu4Yz5mOzC7GsTXSdivFtF82QAQ
gqDt6FzC3KjR1b98PxA9YmOLwrCZP1S9CetXtagPd2EgVZqopnbxH4QmDrudOME/
bbNfVZbSH/TzejVTXB3R+SUfrRRq1wKqLIoPEAX924SZoHR2amuloQ+RbeoxSXfq
ceQlv5jZQEIcrrR6alJ6sF1lBiOBNDWXU3wZolLy6lFIlZhlWQ9SOVlVF2nnwvDi
TPK8Lc93LEJkBG9xMai/GmPigPwrEmDKUyYyqLvmkopgf66S7i0uCmZ3Kq2PAcSN
QCS9zsSPSivSGyORWXuV7slY3c+ZA4YbErZdcZkj6qjG73NC5QLvBoJGXODEHJgS
6hcPPBt5oJlHcX9o7Gn2ifGwR2bLJ8VR8p+pRVUPedH6VNktF5UPklVDjmWVLBAK
AXmNEBPVf4MZovRpY014N+THVjHgrc4+KT3vVUkDMM4eidncvIc+dSwwM9rp9PED
HU+KaHb1AIJgs25DoCrJijybWO9GL4THBpoKkKIgMbXxd/UwvomANEJcmZo5U1Cr
y7x0g7RF8/0vZwXhssw0NAb77y+KJDo6+qTrTCqmUgha4r52dngaWGhMxxpQRRus
6HpcikbDYx5uDBSap09od0v/fPXtknEqSkeEHnlpjXyvOHPvv0D2Bq/PYGVS3B3v
iYBwfF1RN+eIBnDHx5XQLu+xb+ls3HYPOvu0Y5Vml/XDudl3hGMO5ewr2Air6cdW
6gwn0jTsQweWf2JiAZMUtyFnGvJogd4jbTDs3i8yfFPf7xd5QL2WZPpFp3KE04ge
jAkWiDJxoomjB1ZalMy9kq1A9f3SWzUlzdsI+6pClJ6+fBHKHOnMJq0PbqhsB14N
wV1SzDlli8knEi3dVhqc28rqJe7x5Poz5m5xelf4QHYuQ6ZFp8UMoJyILlHu2TpY
fmboklIOlPaHmIhyUqcbnHN3yGDYmk6XSbe7l50V2NejESkwBOPhQxlhhWZxnP7V
bN/htKD1SZibkIPy9P4paHyVbFclVdlZAvF2vT434QQSlavQ46GUfq/aCFjHI3/0
y45/V22vhyk9MrL64FWi/yUATDvssiulG364iTUTBPlGv6JQpSsEwCih6VLYigEC
cPd6SgOWdDJZnaSgWZsm2ETQBz9yPMKzSS/K7PUqzxc6+lLyStHW3Non3WKJ4fke
3ek3Z2lGFBBMvsmIrCk9BbHpcVQ860nTgn610fTsfFiXKb22CefgirTCu34KXck0
RZV/55+4lZoeIv9JDacb+GRd2azg+yi/ejMD0hrfQRjmjjqmu8wnl+P90G8re8Ty
wwZSCSY6+AMELRIQoDRI+W6RpnPEZam8UmUMMfzhMRCNqZJ90Cb6VG+BxnKPgmWL
HZQwT29SYPCKOPNhMKmnghKHduzyxQcATZOO1/aiGN8NVyLolGc9wmIOAmPcxTzK
3p23/K0Wh5B3+G+bqUwO1T5385GLIA8Y2vHA6EGJDaDxFiuzPT7JpYn5vhOBkFcy
vUPWchrT1YAKAfEi4PEOaXF1RCci5iQ3Thgod49RdHGhDtEnClm+rLRWZbbFdw7J
VcAzkO6aKi7jz5D/VebfXVe6laTn2Sq3GilLb3m4Xzsxdzv8sD3cjedysisWaD+1
h0PisXEdvbAWFW4A/nHiXcUVJ95d3WQ7s2rp/bda1/hHsPFcrYQb+3uXSexVKGlI
s8JV4aBBHq3G1Y4i7i4BqyM4J/e2wR02LshaH5R6XDD5KEqu4msH2XpE6nXDf5cN
n7q7GcLIuzTa+BkUk8f6l9BT8Wn1hkCh/fbU/F0vqbjbabmOwVo57f5jG5SfM7MJ
OwAHmIsWiR0aWV1MafmL8zxsNDdr4zraVjdN4BNEFwczRvmLmWDx1XsKg2OrLIvM
FfR7hnYdAjebjwZP5wkY+ssN4BqVlyPG716imKmWlYlqch81e7hOYuYlI5ld+0wE
jjuLZ7Rog2pReMgcl1qF9WDswsZrf9tQ07HtbW60TtqhZVJaUbXiSDQjxNuXe8eR
/npMCmYZZpY2UkHFGKgrhbW0xzTwiNrtdAhurPN6M881lzfvIr0oaJXH3J/Pwp8h
nAlIiYPthuInA+xqkTTCywI7BcF7OfxLw1a19jHdLXH1aznaTJ0081YxtCGCk7wy
kNnuM6dE9QDNgITFVC5HOkT4m05eJUy6f96BK+dWbDK0kKasVwn+Dk9TCDnrOS9p
7WWaNeqsPI39Ox45H12fzFcvMPYjMhpzaQ4656kSXSXzDbvgk4wPtf3daQKEyzNV
EBNca1UDHlGqhKm7/JbiD2/64wsWHkdIl77SeB2Kkk9BxU22iHbWYlroS/Z4KCHk
Bcr1RTA0Wo4Ctc1EBcuZ5Jk5osH1aCwvtwCCACf6bQ0ERDya2XWAOahKEZSSfrlT
7bftRjqJ6hXSSa6s6e7PT+9qF1nc1w4RDXqddCSKe8rvMcL8jDbqIqs/l1upKI/A
60fjtKj7+iPVoCO1It2/Oz/YkIJknoRt8/RAejcKCMgT2xT6qCa9tSr0Z0xdSfbR
IrgHrCJzo+5o/hRbt/+FgJiWKlDRP6rvvc2hsUPHDI8Y/GGJKtzZXRvQpUscDlYQ
wRGyWaKVUoUJKSuF00wjoC/gWFMFBSTHZqT3KtvKfX2bHmTAF2Xqu+NwmMtTcthb
dL+kHvydN7ZZRYv3sqzZDbBGD2y4i90cI+vfXcCxXrYitst16iWHoW4Vs/z9azAY
d8tj+kqRbI8gMlnbhaZqPJxiIuy6EbZcgyiaEwJzxAqbGAIGmEi7zD3aLXSoD1yW
CqyTq1dyfv45r+7o7SI8D5TzLXmfqhLPHlvFV+IbdrjvqSk37qVBFflfSpyozXHJ
SBkrflz2LFYD7MaTsYLQCAmHIG4CdpmpiBsqQbpCD2V7OiWRQQt6bNUloXPwLD8e
PqxvF8FVrpP15G5MmGGj3Q1+aMH3VKdoZ99KB1+IgKWztTnecDjC8uX8f3+Pzn0F
ijUrTt8sOoUIRGu8MTt7swVxHuBMjCW7152hvDGbarqvmJLoLczwMzPRqh3zMj8s
lkXFKG/KuwyofR57C3OwhZKuolkT3RkoDemVhh0YOJuONUmBiF/Cb7X7NsR8Wzdm
GXLVg1DruGI/ZdsFO1YFSNR4hs4Hnzs6wnH+RBR0lNQtIlBAMVGy0sRyBO+cAipo
KafxXg7KM8mEqIrg37LdPWfJtgybAkanv+wi+34G73Z6zVnBx0Y5FyQqrGnfczE4
uSbaRZjEx4iuJ4iEmlrU0ET9cZi419CB8N4wM7P68Ad3qaXFUcVIYacAGohhK+iX
L5G1u8rJqQv+0y90vpDeHEEyUWyPdYcx5rcAYwBg8aI=
`protect END_PROTECTED
