`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gj2hlxNm8hrJJ/ih5bRYlK0xCM9pV/wGLN9zK/SMmxIgjGXEOg+A92htflAYXf17
X61icvY+pz6apqH4mZtl+tA4g0rkiwL/d9Dx5YtbIYbA2jTesbOpvl1DZMw73lWL
lW75weB1hq5Fh5YD+szdXs6RrqeC/cXxm8y0EF3sfe2/v2yHZC05jRngxTu8859n
n4JHEGvUuHP4EFWiBiCFgF48f+Yp/xbSEy9Q/ewDlDeyXDohP48ODh7rzBv0i65T
pnPReo3yvhhOS8Uvz1lTETKn6GH27ahY+JJtqaIMx/0HSjopjxOq1ueeAKqP0N82
2TU0qUANBLTknbq8pqolaLpY/KiTY3KZOylik+tl8UOD4kxxlhMPAkgubmaygjaC
qkOm5gIHucC24Qte+MiwA8PTbzxdtikLh4Maqu1JVBAKCuhX9T/XhX9ZNedFa7wJ
kCiTrBIE/Y9KWn02mMGbrGwNWqGeKRGM3tiIqr4h+LPbg2ryD+4uGu9D8IDqY7Kf
r4B4QoVLcrnre5tZ65P26d67HupAgewakaf9ItGeHnk=
`protect END_PROTECTED
