`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gQxxYT+/Gu92pEUw3STnmRZRtq0ByGZ2H7+JTmewX/qQ8skVNjGnNUc4vp/B576I
Pwqvjq/bk99nW5f6u1vcp7JJVn5sMV4vt296DtN5dbCbjhcRYanfTnSTUBhs4Y1a
1AxKhjDwh5Wcl9bMzgxNYSSXNvfcAvJBS0R3UHwpc84F65KiYtNpxBXqsnw2zf5t
0Z6rEy9DDKO6bwcSZpTbt3oLIjYzAFE0HV2KfcxqmIGa1jo3LWHbuDnKx4/pW+HU
20WJlYVMUZ8Wnh9nAFQW10d44DRHuSpLzAOK4f0CTnSGPVTyUubdBCP0DthJOOoA
XjlfBbnGig8RJMY/BPvLwu34fyLhGPDGzy/fQ+Rgi1UCA85N83xh9jyQb5hNLlwl
i9vxbhOZRoNjH1duPjImPSStuiY2tnF+o2In+cYrfYb0wPs8P0G42zCKasy2iqKX
Pmq0qQrrQaUSndRlFbiLn3aoo8TnnwyKSRYESxiXUi30ekL6l+TruoQNNR1ccx+N
KBxOXgrqrCMF+FZh+4LYf4Cpe2/JAx06/lN9s0C/bJ3l242AgOtX2ZBAFUUng0Vr
01h+Bidz8AaKExNSYiiyPIn5byUt1qaKbtE/TIbwC8QlI6kLLsqkJCe5H+2/Nh2M
xFqS7Nr2xHEdrwYp7J2VAGYemAX+AbpR4Q6QSX/CJfAViUFm5L4djtTuyf5ynhEx
YOZvDRbISt8Ejs+HsVdh6xVeLESJB2l53T73ymdrbm7f4n0Ku617QMjar9Ped3Ve
Rsin9rirsd88JsMo4pkb2hfaOKeNkxokyO+m/SnnOY28ffciy0HFGMMr6/nDLKLr
p17rFVWeYignxgSDTYX/4TysPil0XkLW8YjrtJsElC+KlIwXxHgylzTOLkybdttB
LVMi9ED18zQiCTXutZhLFGsPrGTKzzJYKO1tky5CvCVuIYep4uHbxMp8u0rC0cFl
ER4BJ3LxtrM8nmqyTgQgk2JehKpQduq5CkZbE31RPKUBLy6C+SsGvn59jx7S84n5
Xdokz2N4+Ky7pGTNKnm74lV6zIqaozgWLg8Fzix7PCxqCsHBjbGTkWgt8wCcVmbF
g1iVnH2M0pvC7VJ+HFDYtIbg6wUFyN3q335Alk5p5iwhCpXr27ThcJ+MTCl/3UZI
c2oUdQUCgP98XUz7vDNaqe7WaSH7KoEeUqysKckggPu5X0h4FBXOQ2So6mkr/7j4
rj0HEQnUe0LkET0ZGeuygOQOwbLl90joIKlc27owARbRO3G39DFOod3Fgb0H1F4N
IbpjKKO4M9dYzvI/eCCfa7Kh6XLiSqDsccfun0YEYEzedMHeOXZCaj2RImrHUILS
QSFkjUvsfzvmMmlabsl3lquvpYpoVmfMcAR0rorSJ7WFhqc3Tgv5GoVcO0X+IBHC
v0ud96u6RI+2ns985bc4T8NuRYl0owaUm4+utr0C9aIPDy0E+IXwDi6b+DqIRZrN
VOp3DCvNBGmev5Gi9xeY4MFWqfYFFmvHUjdZRnt6SVbEtW7h1AZ1q9nNbV4JgV3I
SInLh6yxsXJcRxMStCGa8VYqr9dZaAKF8SYE6RUaezawvrbmZsjhW3J1wlVai5Cp
951FTpPzvxcWHQrjv+exgLTuW/A/FOR8DVcA6s/uQyQSd65vwoqtGTDhvx6uL1HQ
iAbM3EFR7XxGIWFThomx2IMoC2xoNn6JHw/OLLi08sScQfE95WdX6Mlr0yMzS+1z
qLMTNEFvUMiJ+UhBgZ+ZTMi5baaxHJivP6JtSOEjtjOGcNm2bachJF1BLBLhvc0f
N/GXhg6FZWxbiOoMizAO2aICTwcc9OwD4EbM0gLTiyg21Phk6BnrkzA6Purf2Hpb
XYTQYnq1K7SDw5EaHfRwfRDb+iyfDmZiHuX1yG3EDLA4heqfFD/7MkniDU/ulSvk
vfGyEzHSKi03V02WiQq060pr5AfkaJOYqp+BLZO2MsCGgB+UlOg9X+7Mkj2A1YXi
3EA8sr4Fiie61t333PEH5lFIItZINelfjfNn71FoOY5F3owb6WqQgUo4fPpSdpvw
SlK/W0AZqNjwURGzH6rVASB9supIvwbk6UZn5rm8dBin20IFbUnKjAeh/j38q7nm
Likbc4XzC7w74RKMxh4pdrVNIkbT2n5ZJzZXiysSC+YGsyWROY1+bI7aQkuDlv03
l4t7BTeHDshmSWZbx0+jf3OFkLmiUBO1HdIatX6EihsxTL4iys3rIF2OwATjiEmV
Y3OnxHd80eBd16o4d2nSR8mbZd16XQ1Intd4V9Mjawvn8pE/aBW2kS3V09INyLMQ
7WZg5e6dF3O7LIVIHLmmuRhuIGKd8t2IkL6REBovXTOnEgzeUgSpgfCS1ZstbOZb
rw/1UhiNngtgPABtDiGdO7vXki9RkZsRtnYiUcN7ArZl7NDbFh0L0PqEQwFnHyeM
p2LvXWJSItqkH46P7V4JiwvC4irc/w9G1/b/MGEo0NkzylxaCJr9iTD/RJiTmzzX
QHFNsYTvRHcC8v95huRhYZJoNRGwVtFnCg3Pv6zBLR9dVlDUosnhEEWsOEAnH2P0
mRlZCi/+mdaW4yfiaU897n+lu1KQTz8KFEEl8SHABtw9ZyQDltH+9vcIccH7Yv7R
8Cxf53d4mfbmb/LLlQSqRsIaxxLst3LT0/XR7eZqZrLhOXJvkOFZjzuIYCS/jVcX
c/3om9Y2ygyFOiliaEqMohLjx8ghRKSrh5YdfNfVXaBza0xtBbTMjojBYK2NRMgm
VuOiOfA9wefqip0U3dtuZ2cP/bVdumTuG2VCoZSKXUNdYvAKxcIlvepga8SlI3hQ
NJuuIiaNO9XVvpJCuw0W9Ms1lkwEAZs9l1QQWSmTPOKvgmn1+YMXmyUQb1+fty6L
hrNZbo4CnJLmuNXSzlYe+CD9jT7xjC1fnXav0wuXWe1PBv2UTuYmjlR7W3Hjv/tW
1fAsQLK4PPC+Y380rcWF6OcsL2zPoBW3IA/q5vT3YQWsnfBcJkhwaDhTS/Y9PuAs
EduDOWA9k899crs7uCESwQ3qYFR3fDxjF91lWFPykPa2sOtI7XETeNggenoi1UI1
2ccyn+Zffe+MPMAV8fkv/DZt1V84JVwMKtsbHQfAXwoxfOYrPDUzQ9WjLeaEzrmx
UfyGO9mmMdmbA3Zk6nFoXvDT0F7K/HAnGlBdwIXlScbMvy/nNJ+xaD8As89mzLDD
DP87k8/pV/rwdR73Y2P7wBSUZbdYRHPfunEgyRlF8TqVFj/pdis85peqcOmyDdEG
m3D8ozOh5vgcNdaNOMfj3x7/9RzhizOzpw2Gt8vkzTWrdVeM5GC6ZfX7uTBCsTKQ
5Hvph54s0AQ0QEY9WuX4xUOuMN7mjuiLBQXm5H/esitQzDvV5A/AynS68Jz/G/R5
l0+20MQJF375v4En8ELzRXFFqs/wbZ96GuVzpllS3ccrNyUtRTbkAyO8mwRYgGUW
GTqbapKyRG6tEaf4Oj/N8atCsQXS3SbgM0VZWkpVOupGBpoHzGt82RUfwunOa1qk
L1WUoBO2gmP1eupp0YDjEnFu7yDANpakUjXSs3YdoL9/2HZa8rz5nMIqQhI8izj7
UgTfYntB7hYri5UkjnGQLfeK1nmKctn+dQV7JA1qhssnz9suMGvk56lLA/nQaM1K
WdUoPWxhJfCmjruH9YiCFU0KPUe6QIemVRqkegqYf8VkS6+eb97d1KaBn3iYbz3c
IXhJcpyYxU35obLYpgqhQP25pRCAXB1s7HxAxqXokaw467AQprHjST7dh4qoxYIF
1ZeskbwWGL6hPaZahaq8oCa4hmil26Rji9R8pTMPTZYXiduL09y2/yZyTV8z+DWY
KEHkVKYQIgPanEYkrHGzRYS8P8BgxaGfbAKUvARK88iO9iyNQBHcgF3AHMQa+W04
lvKkcUM3ZG1jtZZg0kUESroHfIm4Ue32rjfk3EOtki/W2JDtCN77EpI9LUueSJPT
yb/0pDBwjf7rO10toTJEnduGUofwhb/ssH5zQAWs2o7ppbl0IOpo+IAwWPRrc4ub
1WyoP+uSqjKloUKpv+o+BmcH3vPHbY371iK4RLdbHZSRh2zJNgPDDClg55u1Jdui
prYBeK0QhTWpdebWi332Pe6w8M9nlssY1r3j2m5lVhcZPybZcsJ5XJ+6hWdV6mcu
dSkQ9f+xZ/mNpMtInre6z6Q5VKd8vVjHpEeFrIDfZsKrtrT/XheJbYMerqBp2Q4i
cUwElRaBUfwg4D+F5EOBAcsc2uGJR0osU9A/JmxO/La7iG/6F9cQMqkoEQx1iCDI
krLbyHhx7MDmJmsLnayj/ua6G+H8Pzbm1dbuT+eDapHn1IkbJwNpgc4a0X2x/Kst
oIZmyFEU4Mty0DNBPb9mjOYSfL8SkOa/KxLEcquekGfAdMzZoj8ytbkjviY+LsOL
CLmE9sg5qVAlTbD5V1DYJ+lI+4MqXnxXtbBr+ljjceSCU+V/CKSin3nygKOBg5NT
ywEpaVzyyuTrJ2DC20PUE98+p4Pc1RD7CpGzt8IcmVfVvSzyYkmth5jnaYh9hnRI
Xn2GXrHW6ZIDqEdJb18oXtGK/B0XoagZJJAlzgZHXY3I9EwAghvZIk2G/AJ3B1qV
zHdRCAiTt1PqyybKBVcVosOpJhCvnfM7ZDQgvi4UKYWyWJouJf/Vt5cRvkKb1RgO
xOkgGYCns0W/0YS7F3kXyJIq28+QroBtim7QCMTDldtZ1ooAE1oKcJAfwEwsMKMz
jwb5RidUjUd4sCZPeo5SlbAXcICepyUYBCe7FIcYlgrufjpjeGJfksi5IQPUya6e
7x/om2PIjDuG0NR30fpcXPZ4T6DNEIGypY6msO0p1YUsHbqG+7pkBGDF1LazwPIl
ni3F0v8kOjYDuPItwTRZB9LaeSucvm21nZ2DBd9kiC+pyf4shJnsccavC3D3dr1+
Um+/8mZY/PepSSisKM1262Rwrz10PqXPNp09rDcnB5clSn9xX7vUW1B5XMQOIp4o
ez9eEwfDao6hEaLrkelV+0xJpT9RLrUmIjjGiDQt1yUCLb8Lre06y5MJtvsmwgxO
sWO3zKh1IgyPG2viTLtmbvHJ2YlQv4tTiVh2ff6wpE/+ADxaAOUiKmRzcOVXfPvE
qrrCmqIgAYbNLqaVPTMFZDWTAHuboob0ttmqGvMBpnjDR9Kh7h71/k/sragF/L5k
YrPXoIv545r4arFfBUbfCHd5uk2wfkVwH5zGYIBkeIuAxWSviruRpTVhemiK3nmi
VABGWv1Z8AOuC0q3ljCEhyt6dygRR4phEHpFaYNp16bKP1Ieb04FGgNEpdsp9w4p
lnQ2r/d8JrdqYqgknt9KglGtKF4GI7k35ZonCDE1D5+u/ZiX5wOtn7viMsauoiTW
c7JcMmDl/M65WvmJQXqorMyM27cbHCbQ0Fek87jgqsyTvtrRsr3LGUe2UwY/nDv1
+m0xLAi8AbXbx4beW9wTlAmQQ3BF5HJ4z7HGZvJyo3m9+DVmgTQU5RvSRnc4xauy
32STSR79XkB02skJyJbuEuQjci6KokojLxtxs5lIdoE6QnuQqpYqK5bgN2mpaoUy
3+exLhKDB4ZtFmYf5fh4lqxKs16bWcwgmscdGkCLXCsJPF6vre/vQJzs8W7dmSCB
ERGWhMWQ8nI2OTHiU+JUqWGz2DkhRAK6+yE2G25ykaklYrn23A2vgMDPrV+iFdvH
ieiRlEVz/JXhwBor1IkyTcMcVi0oKHH0BXGAns2FSLEvLhcs2sTdtL4pN4almfEd
WfEoVQpvLH00uSRX1gPetpaJOYzluLQib/rso5eapFlOd3HwKCAFgUdxz+BVwHnj
EhWo6oqn9V1Ws0iJni5Kc3fHwAv0UeBdB8wKv8QiX8TSHH2E6wrlnZlyhPWZ+sfh
HsyRWfF7DzmAyoDVoxuYr5tSTxfCzxiLGSqJyqKBtWFU9zmRT2EBEGjSMAhuGK0Q
KdPf5m0LuQFWMVkiwtOxh9BYEjZ7KQ7jFi9Be8efp6snn0Slw/+pmcfi2v5fjuYs
Ktb8Lom3Sm7eY55233t4iWjAcvwFtD32t8mMyvIdSe0EYFwD5zm7iml3pul0s2dK
M2Ts7TPtb+ir6HAFKTnErD75R1JIXZ+IyYY/Z9lINAMHAGrG3kkx4TDSJ1d0pOTh
gsXRXVjFUtqqmFNYpNI1TtDI7ThcgO2HTqQWYrBAtbuxPLMOpycRbln1wsfkm7eu
s9IqYHeM3xs3N/C7EIgXmaOs3V8s3poBIxOJDr4PEX9BGLscgsq5Rlzn2J7tNSHL
kz001bHJQVq2kqGkxykVcxBGyZO9JYyCyDOQv8hWWlsFYN757X7nKM5TnjliYAu8
miud4dvir1dtmZ4WAcYRmt+i2mjRMknrzbOOOdfvVImG/91l65nAMG9742/IVGOx
SerQd6z2CLTx7Do51rIPT2oWF7syFJWdV/YtXqFZQvSQco5WG1WOpQ/muvbgB+EZ
odpeKu9fXD+uhAczM+SJ0IY3j4gvf6wp65B8buBBnLodSGnsay5rDAhfsm93wyM6
EnXHmXRAN/xC9mO5gZHqiTioOmftjZo8dr+B+W326TbtedpziPk5kju4+Gzdv1md
3LHM83XOcEpSIv00wR01tbbdflDN0kSobGypZCa+Rk02LN0m5TjWhUhoLT2L1BFB
9UN8u/7piF6WyoG/9vZxxWYwdj7J+ejtOaXpWe4YqU3aDvq87MnwFWYPls4NV0Lv
JhPhYklcRIjRvrRaImJTEnq9Gh9TYkxJqY7HxKgj9Zh0cFJwr5szjIjwSvixLLW+
Q+rUNl4nzMRP6SCCDz0SwSsunVfJUigpCBWkvyDwAHcEX6xYqlWAbXxJwOub1HCj
tNWeGDqm1hFmKst9c2PEXiIYNrO120yHzgp6Vaj7cfDLDubev1kByI2krdcSYLOc
KbIl+ipVxKywL1HFg7muAkC/Jqtb5u20Tu0tnclOaDvlZliHPtJU1Uno4ZhWiU1+
s/YS4FiospQyvR0N48fxdhcidr2dUk8pIpvjb7G6WsdwmZdRjo47XSIQBe4dBMZ1
4LhjZwnaaKxoM6VsgJ2lBgITm3iBXiEOEWlLVJcPH3R+vz+PQqbzdX5sSL689p3M
TMG0CUnwXtTAmSfzXOyPkAD/AGRUCk+hxSZCZZwx6fg5Ulyn3KZ71fRamKOPHP5J
XwH2ELfMQMC3rfvtiCjHyMPlRmxzhoIftkk6d5RceFZrel0F/LT7SYiGteX67NT+
DvWOI1F5dImeuEnj/lwXX9Ktft5O7aHojx01Xz7jqSWSYok6HuqY9zlv8tNl9PPe
r5hKoUlijFnEKvkjFMjUZbkIJgNavYBYz21pfwhwE09NkQpompt56SP/qzxoumd+
IZ6iJVsCuh+3lQzrVLu/dSxfV3v9s1u67GGt+6jOtcjhASf+IOLWLtg7IBza8oQL
3y7MAQ72k2I2HAq4e+K3d2DbRDKNhd9Jr3MqH7lpjPNL78LvFJuB2pQR+a5m7mki
q3LunmVfj+SzPAnMnabW6SZmBX5HDx/TXaMAbdPT31sHdVceqMKmoFjArsdS3SAr
FjnCwBEAqqZ2Yl1pGbjyevzmH22HuQg4R3SGPhfEGhjA7PxM/c+XPYGu7zDihWXL
yulYZpX/+T7979nlOiG72Fhqt8pxBnnoATAU4Kqz1Ayr88XuY1IKHD928Ndicai6
Z+GWzQ9U9eAmFXu3QA89QLxlAC7of4D/SrJI1DAS/NUrGNFog5NWw4DnDWz/puHm
IBRcm0piqOp3D6qZ26Q8DWYo1jbXZpFyK3KxULrokuWiOrq5MybJy7fhI6okHBpY
tBj7l9oSOY9A3lOaC1H8TZKVUU0//BmGXO9mlc2Vy5ycpuRDU5HIsjMx2wV5ErZI
0k6j+Pu1+zrQd/uvs3nBpz5zCJmZ5V4wOpIn0UW7hnp60cArhk7M+bfNkOwE6quq
2ClM2nbYUhISjN6CYR4H5tPp1TOe5qHILnigALUe1EZVHH7Mm/6YiGBFkLgO4qJD
uY2ZmAe5MCrIb1h+GOqyQi7cuz9isQbARzSUsR7xpsP/Xry013w7QaG2wNjLP4aF
YkYNZEyf/JoqLrm3UOMoEIpuB8RU9MMOQ+bACxXjlrO9cPeaDNmz2eyhvMHqGfyO
fuYyPjAE9oei855dXY93sd47+3zDA3eTnoWqzVOx6GwD7RKVearFIuT1EmjEB6Go
vcp0WGFD4lcqkYrlhOIlfMq6EtDB/Xg93hLFYs0OzNyKYPcNZRI0MlLa41keDnb1
zPKZJTETGu93Fqx3G2B3D0v8ULvQh7MJuuvOGBCsJFBhsMjimlZITTHS8HHmP+Cl
zZKqr8wPcVBwk2zp/vBqhX712OeCwt/iDC2c9Q4OyMcFEdGbXBJQR59jfKRTtwH8
njAUulwE4JD1TxTzWnXitsJv+lYuf+1Plsg11qM8aNPQsjNmrBIDz6CvuwuGUgaT
FjtyiieLHYLwRIyLchsIfnIuxSqiArCFAJG8j/eqgI8EazIXoXTHfQ1Th+Q83Zta
Trbf2+MH/362g5mefoIE6oUnNWgIBFs3ZACZtnuC3CWYKlTXMX2GUTjX8wXuNV2t
RVLLcEmJ2zwHqIvBA2zQP65VAZ+Z0dLp1zAXY8E47NNi+3EIAdpc3LmpaHVE6KM9
2n/tP5JHjjBWEVUvNngiqqMHgfwYBO26l7IgulUF2uR0lhrm+l9ZfyiYcrpuuWvG
9Ss4QIgHInAQdsr6cYk2TsvE/1UH2/wQBmqIlcRImHJaFHqDMGuMsXdSg8xx9SA4
fpB+pcFCYQN8e3OPrxsMG0Hypec5Nxy44KAJWYl7IpesiFNVLzGUnXH85CVBjVVv
0P+0ELZ/hV58uqltfYgnQ5jCxQQZlyyAom+Ct9hfWLn7nD+rlrT5WPDphrlSd5Ab
JfCbAV+XGQojh2F6YaEJNpNNRZlri5va3HOdz9XiwvE6E7YAxB8aEvyQmIEbc+1u
DJIFMePUeq5zjbxRoSDwOnZ1vSdOg0bOoqvZocK+YFuj2lQ5nmjGy0Sqi/aOrQ2u
dTHOZi99Ga2AWtk9ONaK+p/E8fBEEKDpILXtmGd4HOd2C68zJsMAoq9Is+M2C5+3
zaCd5+mglmzVhHBpgsU8GxcnYyV6I4/soouxYI+xld+WC5/Is1xPV+ZIuKHxe/CF
NvdrpgPgIGY13AyAxBiip8g77k+JfT/mH6CaBr32kALRbzwdqAapVx4LCtOEaruW
0Uh9f35W+pACR5PhkSN+XiMnA8pFBYokGUdWup5l9SaqbaMKMROAYjgSKdrPGlSn
S2roEc67PCCphOoOHljz4sF3nXh2lKygRiu8pk4MUdTJDsF0uzQ3hRN2VZSqhLVO
ftXhlRQ/aKExqUc/BbttbdPSToX5WKIrSDLutiZxavVTSdsy6TWHAQmAMRH+1Szj
mWQCKP2LEcxt3cI9JyFgHbGk0vmOATxwxlVEnVZOAteMmROY32n9S9l8G2ecDJRL
hC8heQ/8neczCoEUW2EoSDWlD9ib+ZxKUQeNvXhZda3RhPx77s9krpKceOKKRRCU
ewg/bhJCTVCkL+OPBED/Q+rUQ06uwIHwPEPbzwEtAV1rn9+VNhJScB5MFh4CbnOv
KRtlHq8pyMPnyKav8oZGZ3mmH+UmJ+k6ecZGiOFyutVNt2Kq0b5ryJD4x13OaaW6
O04OLS6argDx2/RThy/bskaWtdzZb5KCxgdiHiiFJ77s6WRw8fSB1llUWlB2TILM
QVBnF4/0ZPFoR5GSn3OugOMyA2rT6T9M1xG5PK8tZIEN4f3KnXJe+arEB2/faBkN
02vDLCS3N0q5XaRIQFrhchCO4z00aERcabN1xManR7tBZ/+OnjToioAs60qbaeiT
NToGe2fPHxnk8j1j5+c4L+JQybJjhjcdhpVxZiwVO1g=
`protect END_PROTECTED
