`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HkcmFOJ/VnyYGgwvH7OdtzND9HHxaAICxWqbeWozesxoDLL06O809BnF80lExLoB
QqjNXODFSRIYFb+jV1AU2S1JbqJ31aasyk7UOzcuN34xK7wDjBq9J+c/HHk6yTjX
RiPwT/7Yv0v3SWTUMZ7oTLSGpaq4GkLQwwwfpm6VWs2wcuXIRQf9LGVSWm8HujLU
nJ1Rl9YxgIwaT7bC4tmi+6fhmLW3EAaBPJPpMBf9UgfrK8qzkc+JUJP57g2z5fe4
GldSsNU/gC50hUHkqimgoSSTQWeGPDBPOmYHkPA831d2CO59kMUk+4fDeg2AnjaX
Nv8s2XEoUXSCHowUIaPEurSpCtx76ycWxaSqpd+rtaj6akhtQ1c8X43aJAqJb/Ko
hz69RQlSMcRJTKTZfLzZBeZZIfgksH/C+NUoD0N2wqcq6xQYDlFO3pSvfZcyWHJq
MdNadSAalptErmV3a/bzrkmPtwwr5IL7YZlQCZmSbawYxHpWnwqSz9WRM1ysQ268
iVE0t0I9pnbj9PPZ+6hmge50WZHj6bHB6F2kzAzwlE2RBmNwsIca+1gFOxDIKSZj
a9ob40cKlC5ua75BydRi4wnScQVONAMOZFkeRMyhKbfA+izSQ6p5eqAjBFz0bTzr
SIG2QaBTi5ppbKrfbXWNUPMk0s4j6dGhNcuSyDogoiNmrHQIJLxsinIaO8XoqNrX
A6Cw2jz9lGHaAfymR1Vydl9JWp7LJkFLSCYZ9r23vdWeD/wzYcyBhE7RX81v/6cq
bVV/0ULXtHxKiU1A6ja+Zi3NEkR6x7HOonCtf26rezQa6a8t7E5yYV95ARboT1/1
rjv3pr/syPpZCvBL2EaindLd2vhT1W9ilGtVDLOH9bmPEnUGdS5uJJfTZXPZxV0A
0RA9xL2835O9Dj72fCkwdSsK5UuS/3rl/12krleUDeG8p2M96zTtj1kD7Dd6Zavd
Fw+ygCUILUNii4uzYRxesyP3TP+AsyC+AkviLRfY3CpFCIEFQz6einV5orWZb9u2
tAPCx1lyMzbKUY4ZbU1nybCr+M372A6AMXpJHaXtoxEbsLLnzmielB8GtHUdp8Hk
3RUc4EJ3A3+jqwHZuvKpvw34VEqkFUjliVo45mzZy9pZbPEFMtjSsfTSSEy1yvLt
3mJPWy2Eb12M8OCstIhbjprqYexQCgF8OOY1e13mXdngyXyxQhgmX5ZeiVicvrl8
dgU7SysayVzKUjkPnEHkI/Ax6k1uAxd6vF5sa3C59eyCe502Z6x38coCqIMOo5k2
/3BLK7Bl8cNW1tXRrgT3aj4ZpIzrjfB3KBh2gQFlqWvh9zjcj630t8Exrlf5g0J4
6amuSwXLWuZ0xID63Y30GKopGzh4IIbpjS1pWeMGJDoc04WKPUl+5TX8rbmXfY0N
C5yxKFruplttS5ZBbUCfS1O/hzH/iTbM8tDEvo6hTZvX8ScWNHV3zdoP4Tcm64Rs
vPmoUjQbxQXrkhNplt9k8H3s+jobzo2yRXklGqh1cm+JyKeKTO8TlL1JQgXcXExd
uIuQgj9XlZ7eUDL2wnzG4IY58g5Yc5HyMB78pSQKeXwM7Qgob47pCqns4ieYfvdT
Qd/Qkwjwbw5iQjarffBj9gWfxuP+iX3kL/EM/78+6d+iu1IHsxMM/OxMAIFX22Gs
+9+rVbD6T5eb9yde8bk2irKWFWTn1p7I1z0RFAtAs2RXTZPlCgigjnGkII3Yc/vQ
Y0L5Ki6wGXPWurmeuH3fBBzUa6hTXK4rdTL//C/u0o6imY82xLyxEMm15Flflv1f
saZofEBam6B2sfoOGwlYsGqqjvaFatYZTmXqZsUiIyKDf47RRbCfErTy4GzQGZw3
IDsQ9IhxNrRuchadns8LW0mJshrP7xVtAma3XmC0R742/g5stbyfEqsifZi1tjU3
ivmKyYRvb6sk5loLUjF60PTjVu1TvxqRFbA3GspIwFm0eh3aIXSTSsE8ejrQxvBj
iWh66xulDdcJH01jaueN1dkHOzxaz/hBYnzLKJiHSvRf8MTRJ9xVHzLYLglX1pIh
8/JrM+aFh8BWUNQXqZOE7GCfFb98rNn5DbdnBxv4PPOIK4FujcncCR99CaVm6dyE
jg7EfMOyW5Vkr844Uykd6Qd51gK3dbVtdcRv0YQjiDQ8K4K0vwuq+aL4msumHJdg
YHUMYgGvsrwWjabQgNBj6J0CPjQwmHFrLiC8o4ls5Fgl7OaexuIELLnFB1tde3If
V0z1lM4sxcdKhJNtbZyu2pTMbp6e9X+R812Yd4df2zg6F67WPzPjpjWpLk+h6KOt
0+ery1eaWL18rTDPGIrOPTvqX8PuDLnmcMgYbcHmdViYCgt4TcbcXKhyVUkci3ey
`protect END_PROTECTED
