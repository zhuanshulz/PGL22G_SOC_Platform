`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r2JBiHQa1RCTVRQ/3Z+Ruok1ZJnUaPu4UgSF1q9G+9qb6tOroZo5mU/IR/Yji7p3
9A/gGGBSQpVhmFJCOnWuVzwDFuYc2OJRWqAXkIYMCivsXuBZX3MpOBGsG+N7EHHR
q4GZAR139SaYhy26RiWAmaP+fn8l62mGLnYpgIJSQjh9YnHTz8mveKyByIO+C4RZ
DyoLi6sjKxSoX7h4089wHO4NgO8Npi01s+szVmA8PtEGktHtrbx7luaQBw4F+feV
RLiG3ZarW7AD7rX7AJqN+5JfTO19MCVo069wUwEDwWgL3K6WeUbQbBvuaq5MJ/lY
nv+bZJwvyS2wTd+kNVrDQpX2htSos+J3U4O3y7IR9lY8EgViznjSd+kK+3QVCRea
+m9qhZy8kpVAdmke5Nn1t9jME/GI6YS6RQxRjH0FTt2hOUWu7TcKB5GeVbZ2Brsn
WYfy3jEUOmtZJWlaOdpuyQ==
`protect END_PROTECTED
