`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e1bK9reyUlR1mfLILr+by4cfW4GvwUwPOWQ0JBx1XQNpH+PSjWQxDER7JdCV0a4Y
lSfJOGyn5Z4MGWP1fOIvbsBLOullqTyhNSYxpR74kR1892bsIxa/31o0UCcKi2Yq
Q3ZfBI66ZsYmyzH+3jW+qacNApjbIuFBK7XyMF82Z7/0J+8tdbCgmefwn2/LklkC
2BTWwdW/QzehFjpkRVixYBRerzATrkOSxxOOXsTBf/Sui3acxLKRZ4rhzQDQDLDW
SQv1tRD0awpwlnapvTKs+Vc3+t94iDKdvVcl6lr9p7utkWbc28VYzlF6RGfPlFxT
qth4UT9R3YralATSfHn3SxLe+OrA6t8iNUqpZpmij1Dhi1U8lndO1RuYHBCAJpU6
h2/oceULP3Ajw5lp4fhfb6AcFwJr74o3foeo0xD1dgZJLN1QtuqSGQTMGj62RtCH
Dm4oq75Ur0WKN268gTbpkvRdWVjsicvtoY0Yonqvd7kvZZ8RWZdKf/+tIVwJh8Me
g2XhgPXt7cvLOrUXSHqnM/fP7DUf6mDCfVHWmGTv5fP0pZSpEFmApPTx4ZWnl4JP
8LIcEynISu8pCvDblfvIFoKVYwxqm3bBLrmjprxN9TCpQejTGAYeFrN5cWFNqZWJ
c5WgxzM5OR3itIUZyiQbjwm6roDikPoRx9TcAs03JSvlstmGxnVeEj+caz6mCU3d
z4fqQ/l/dC2xgjoUCKYa6aoeZcxng74f+8058nrijssROI7nGSgmRX0Y0B4996lZ
7Kso5pr1iRmpY444+Xpkep6taR7hCnioxXfESCpWpGCr0nVN+kNd4m12eKiU4AVy
AdS1PBovXKp73xtVZ7zu5GZ0y6xG+q7HDNMLriiNqG6qdGT1wiaGpaBW5xRZGCk6
NgMzyePhW86dLGLdpx31RdZOMkSAnB7BsUlrQIT8QbBSwgzWmnd55b2MHDxIAw/L
rQyUBrYeil4ydNndfva4CFCnKWltmztg2JbVqh39ChIXKZ5GuKQ9Hh21tEnWE0+G
nUVY80/Cvj8ifoRs11sAHIbFTW6XLYh7PGisdYPCze1uFY30JDFzTHpCN0Ul6fly
ZQJmpIBk3JaZV/JTARPZNUHS0PzIIiwzK4aL3oR/LM37Kan5dmIrcVvinVnOZfMa
/LlFU5B36rH5gONoAMHpy5vNBhHeBKhgawB41TDksH04uPiCtOw00E9yXHakTJ+6
EAvwySHbLaucLgTD/mD2jPE9ZwvLOtKk2aVveSel/cuUuDDe+JLi2vO1ZcfzOAC7
Y+T6qKGbJfEPhlU2ClXbfn6lAIDU/mqs0efQXaurTmbfpEdwemueYp2QCCGlmAqw
Mn8cMTp40s5cTklHwlCs5vOxHecM+YbPHSNh4OVI703VUk5i/X5QBEzUR49YaOGs
Tj5/mljWk+0oAqydVLGif7vmIlXJoFORD/zER+Iro3onkJ4yZQua27FX9lq8mRSH
d/wFKWwhehhFGmml+RpxIkSohsgP8o8VkQX/Uo/vStwuLeKgBAtLUO+8yaDus0sT
8ttHUAolWexmMlFcbm19V4ULM4+xziSFnu3WmSFRVAhfGcfioSU3lApK9l0BSd8S
1fn0b9VTJf1rzrHQ0tcqHqCt8IB7tUSb0VaoNlOiY/TPWzYPUj/HB+/nPLh0Gbns
C9idEU7viztMk/e5dzENbixTnge9kVR1bOFVyGh5VpvdG5IaLL0NjNXiVEVS5f9O
mgU28grvFvOtwZ3c02lUJ2wB4ITsjXygiYfvwMeAwjS5BhfAk4gxrmiwJ7oisDtw
HmihSbcIkvScC5tkhLW2GkVO4NTVQIqrCDfpcqx7ITFEGhfE3a3hPF+4UNuT9jO2
S9jvc91hcLDurO4kxghUxAPnbQLILlck0UVKJNpW97GqhKm+OkPZpm6ImiiTpJUD
YeEiRkT/PeSLQHezzGKgzaaHI88z/2DhNo7122XhTzzHYhiUKpU8cgiyelb5gkJf
uYo0Rd/zPDHAVGzkJUAIIOtvfUJo7p23Tiz9TYxMfuKYfEGaFq8Y4qQyCK0tg69o
6Z8X4yKc8H3phdR96VXd7oetzsq6lasCx5b5OdbWTko9ErTJLi0aPgV5Z1QHXPey
DFJCg8+CDVsQZbnpnw3KBtom0ImTzPLi9w8ujWRPc4qgd16iBvrTeJspxn6bHbzQ
QR35dvL55hHyZd8tc0ToN0kRiIxOBbRP2O7ixJcrNtcE9tWkIyY/PxbHXXxsR7H5
Do0Videv5k96WywNwjyCVRGg7+bELq37CZBEQjJbTAd0s+YMx38ZxS8r89moIwMo
qOAk8QBMD2RKeGKlRm2KU4KIHm4BTLom+emS66qHpovuN54bzz+l5SZJqJuRI8g0
TPN6yQ/WBub0z23G0uPsZ+qB+WRLhDvBZOpKCrnIWka0gLdpY19seIcDKIfma1bx
2j4iGkQTLylyvM6WwQeqIpX+rhs/xgqxTzd06wU/SYlDi+jGeyMJsYQ7uTBjjU1C
kg2LhgQ5LGpOUaVmWzJ9SfzgmHFsCykWSAkcyq9W3odmrtAsgKC98dE+pVjUgKj9
esc275gGI/asFaO29/K5S8wAzB6Sz1IxzNsNOMxfJAAfCsOlK8KfrjXO4AosdR3s
R/bDZqUfRIo+X9rzdXNYf8Yo5b0Q4KwJxzNds2f/1irgJGqRE9BXrc5mTI7kt+xZ
pT1WtB8gfLzKyShdpwUFdZK8FVQKdFTsh5XyyJAGjU20kjFNEnn01ZD2ynkuzumn
SfCDuusXc0SOG7Q7gn4s517WzsTc13WmrnTUlq1vebthIVKMurG8cMyFqiOqUjeJ
GqwiRpCTGAqZHEobvzzl660neJOn0UAN4sNKbaXaFaAdubqRzhVJlF8d3qUCxyKQ
/SH1UZ0N1bZLenNNwAhRXLC9a2tjSgwSH2/2NBuGbvimaJbk5FSyRYewDjfQJPop
p77kkcra3ygEVqrcymUIGy60wNjIWirh+Lixyud6mStr0bnLMLAKH85PB7F2U/NZ
Cqr1+t/0tPghqDEbxV+EoKQbbIXkGZVxjD9Ov/AX77QlQT6Sl7hMZ4YwKmdhOUr0
8j/m6JIactEp+DChFciPT8Hcleudnj6Ks9CyKzEQbWlzHD5DPIWNSaIduAdelo57
/XPheh63DtJf8scgxoTSDsnfcM9ogfHXZQEJFY58nC8L4hmMxSs0+0+kvJL19RC1
VtdCbMk4JbMxxjsSBSsTxKdxFuG2NYm0hUo6KWvouVxEHWyC+hjRaSSFDJAWYARm
0YSapx4hLEemtdvpyfvK8IjYDF0q9ozuVUtUF5qTZUagQB5fVtzgScw+fCN++u/J
eJS2hlo6Hyb7rcDOFjnh1KrzWkzoOZcyE823MS9OyD4q6bvDvruC8tmmP1JpjjFH
wTppUrjXB36SzM5bqHchNgk6oJCfHupxfF65heJOclQg5XuSRoTAcBOIHxc2jhDb
bpPgg4n2L3wGXFEulCVNjmQwzGy9HzUySoYw9AjUXsEUgNpNaamRODTgV9r9zwjQ
po9ni6qBbtyfrzAg9GsEJyItBZg0jrUrgj4H/phtBbbzXBoY2PyVJVdXxqZs2xwF
xFOA6n4lcD4GRtcVrVKV85N4QEvv8zfeUw807BEzSNOUETPtA6GakhDB3AOaTlyq
1wWkAFezGATryJ5B8gVN1sx6Kdl720CE/RNmJCMsRVsmYtzk8w7FCmKmofqzX0qO
Baovtj9OnwGXnbvOO7ZKz2mrkRkYuqyTdOXLkrisRutCqQe7fbeO8b/F7hKBWPkJ
1gMp+5Qe2XlPPWaKYzlvc1iSZVMmRXEvNuxjJsKzHEexNo3FR9xYELwraibA6gJi
5MrvLVBeu2SujvppmHDxlb1rkk9Jq2rb1WEIKx8lR+O7qaIbzOIMzQ0iuSeyPJ+j
wyQjJhFKAx15QRCTA7eNkn2bk2l6lWV6lDb7fx6ABpslFPWgQtJaPIBhtYsKCGG6
ZOGsqcIzD3NqxM6eUPmEiqbdIpp7Mtm7zUYEdFW7L/ciBUBaFa/b6KmsZBOuOyFm
Dksn0cbNFuyrYMUQ+137FqL3veqf23GsGUiKasDJG/IqsxmWqHZuHVWgDg8ZmRJ9
S0aQXdonSeydoyHOtrW0/FkUBwVKguLpK0aGdMcp2lgJPu+v9AuhbEEv1ljnO9bd
9Lre4AjSPsnM5XT6RYK5gxCOkQtkFRQZkQ1c/UgX1iopw84bZJV7KdsPKfTxfxXN
6SuFt2yberJi8ip7oNV4o6K3K5BEaDFOr/fv4ibwt4ctbbctNNbplZY5+JfLATJh
F/9QC5zkgitEoF4rTuKkq2dHZCXBGveU3Ibv24JfomIw5n78TOAwAobzkXCSizAk
UzoH2bb9TTpISyCmVG8SEKY6+oVP1WwR4HVQWs9xRckm75qR6KErcWQgpKAaRuwd
TXvl2Vb+/KpNF9f5YOwjS58pNOfqFUL4QidrZ8ohBaLSPuqQNHCUefLzRjPCzRQl
toMFj7/S0bT4kjML8q6Al7KOeRtaQdYyagwrYUcXtz807b4OwRGxtbV+mUqx3UAD
LmriHSgU/Ezf6cNGQhXLV8d09zddtDONWRUlCgkH0ETJRoGE3WgoxozfuR0xqN+w
CaKfC4of83xqLOYoJNfbNysNNLuyj68bcQZM0DujTaYZ8ikosy30SbpVxYLvijjy
YXN6j3Q/Avy7u1RYmS24uTZ1uhajGoEhkfNMMAI2sEnwkGut77G2KFc7n0BDxmos
ZsxmB9FyIBmLa6Zlrh7Um/TK1Y1x/dLWVwNn43UkxI04zn1TYvkDrzxwD4SlG198
3SzScCcu3pMIcdegHCv//osX3sodoSV6NO2qetE6NkX7dMU61gO++FEm6LYjknTJ
mHXC1VSBRV5tmLp1LphHYd0r+VjkDvOs3HmQEnvsTGob5g2Cpq5NvNtpeVh2jzJ1
42yrZPoO5LdhQnFDgWlAUIMLt4GawRYKx2sLsaD8gU4=
`protect END_PROTECTED
