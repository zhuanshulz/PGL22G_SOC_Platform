`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u7vGH4PNOBLTgFMkN4ZZXlFgOFLCb8zIroXuvK9IKTDMaGE5TAvUe4mU6YNE86f5
+zIFSX5jicCMS53+sCEnCYxaRAcmV/s93PVPE0GaHNSsq5sqvUbAsRRWlXxAOwDW
fzofzomu2yw5C5vD6EmY56x1cIrlJy+bbeLemzyUESDAr+BvM+ZAff6Pddpthj4d
14PKpdZdNqRPcXmbDyY4k5+5TlZgKeWGcErafk3Vb8/t2xYUtkOmMhxAiF+HNh0R
mOP0tIEp9bQdxiM817N6tgqNFAgd6xJthJ/LO9DEKlCZ5ai0f0YXvBN6/9aFoKuK
jBQhW2ZGRa7gXnngWzoe6g7UPKy9robSqRV1Mn5x5GctbPikqCMeUY2JFVCi4vRh
Qj6NghTSL4jjTJxw0D3ypCZ/+RS7jpUnsTGEDWt71hKQ22GqD0y7CS/a69r4pUFS
BluDLYKOTF5FUA8ZrhWNrggeArvFgFPwZDAHspF+M5W7JHWO5kLncXp/nHOfIEUW
eyuhkavQG9B9wypycUsAT12Wu+AxQFaAT7hj9umQj89YOMF61O+jb+oY5bOvCX5I
aOVpz83SkoxiDTHHhWxHutKF0QtONGJUBPj8BMZ0C1KMi0fjkUsVI5SFOs+vyD79
QNzxQqhRNbv2u7Uua6+fMfdrDU1ikRueTy7XDHSfKxrNXsY2C7TDVbXUMuYLw7aN
QE91WLTf9x4eKgnvI4S1v3zTu6rcYMVBaGRAtxH6RzMQLxWTPFtO55iyTxOzqwMf
wUq8bUVbn5fb1nyvHV/SngKrfT9omH1nR1xqdpTDMXVNVDP13BndwEWz3ZxtZ+rc
594BlzwuEX1vbhAvZc7lBFu0MTddivt5zrt8isinGkjWdeALuy0K6gDJZPQe4EQx
cHyZ2wITRzUnoHwM9pysrz3SaqBatw+hODFuyKV8qT2Gp12yZu56X5Z/I7kfnRQ9
TjENGY37aov8KLAuUbNtfCaFlJDWe6taqjGWs8/t1pt0MlSf6ZpOSxfCT6ptRB6Y
Mc31xUWwAKrmfUYoZ8eOtqyK+WyIXSzE3gMJ1GGIPtRfoWGKWrhDLz/0hNFaKdsP
pWz2n1tN1NEk2wjVxwMmI5llicSv7EW7SY8bu0VivWd9YmVQyAwE9eNKoPJrPZ/F
O0wTwuGfDtMk9Kmu3qg15IrETQ/1vYnEyieJZuKGqHFOEBcG0mvhJ2Nbi7wdTyKD
ncoWdfV3OICuRvcx/fcYGl8G5RiNGeLWZLF1y9N6lCwR5zf7KNCvXjhc44WN4w5U
dctj0M+DD41SYNV/1ruxR5n8p+XyDjdpqXh6BUqxzYBmGC1ec0M+pG+rgsvlGucm
93R+Wt7v+LAqN3SJ6AKy+0Jo/MfcjLR1Xwz2D0IpsV3vrDihrgxB32CTnGRwSyI/
uqHhiQE63/1t8Y1EjLeHqBKPclGjDoRzwb1+EE5v2QyF2urC4dxT7QhKV6RTb1YR
duxO5IxRfyVq/BrNNgTV1HYb11CCZYDkijjEjuTQUc0uKcjmIwagrx3m06Y6gRcV
ePDyJ+sBRq4XpYGNRPOdvmXMgR+us6l17oWU9QWfwAiHGxYaoga65o9nNaZgKvCv
gTA3Rpc/PZDn6+CWytbDkB4XDWK3w2X2fOvhNXHr0VIAX6piWkwhH0ZfmULjTxhK
HiL7S8OTpx6tRtLsV896HULv5/+9TPaw65qfvfD9sUc3fTAjC9KkiUAH9Ljn6Gy4
no2drmLAZdCgfzvBSHUUPN6FGtdLdHGw66ZQ4ELHl+DorEUJ8WCLkqTLnrf4upPc
keZwauqJ36uc7w8h/6wHt60Wud20jHrrt1hC6K9OZJdLg/MA/5g6FFFfDRmaF9JT
ofLdOeo33bd7mTcaQcL5fD84ihmU6FzzFnnZCvXUFb7Mc/zfw4i/RoHpkDJF9co+
58HEA6uZ/mmlQBK+FDygfZgiMMW0l1TgmxyhGKNqzDPSNrp62Phqp7Vwt9a145Xe
vh7cy1v/jq+2ezW09Wg/wUcCXu/jZ1dXbgOr4HXCspoWfWOdg8r3OMIrusnuG4bN
HRhdgcTKiPY7JmX4QT9sNr7M/tORxIhoP9F/fPTyvqmRfcJyqRN70MKrvTA+zoU1
Mq9QVObnbAbYvIlJx54A8Rq5hdxVPauWZUMgXv2vnCbRX1hUoaGgb7XIEGpDA/I5
wgbCmThK73trZOoe15KosTU1rqurhh2jXCjQq9e4kydIopZ7WwgVcslOL9ozWA5A
23Jdh7Z6WJ6JxhYiWEBqQFijHY090Jcm2/pv8CWvMjHa/d1Lc+8HbdQvYpLHeiBe
8UJsrGaoiM1Pvlh8etITgeJIKXDYAsq5cvZT1UrK9AccjoIn4NRJxG0D5XJMeQEB
f2JgSe+kZt8WaigBdz12rA6w7AjzWrYnYfmxkaPCNX8AoR8HdSC73y1cGS2dGw8i
xBcc0y8O4A3XcUVrOqnTtjRKLLoF9MT7vBQX/1u/TEnySusO+CknfVLfCU9QYFZk
ViQLk81//0LSSEpHzlzVXFYcik9g2oSEvvbYPa1kDfCbBLhQTNjSArDq0wjboA0x
1qT4LJmI8qMUlf8wxkjwHIf/AQCAwlVvv9t5X8FqIpRC/18ZBULOP05KotT3+oyU
raLppMYg1Np1xSij/N3AplSKiKXcPkNMS+x93r9vaekHnAiLdWuY5bilQqVepSCR
Yf/++/j526e3ag1KGCYrXQGGz9aVPXDz2iZEJ4Yr6kjzAk/tJLW1sEnXKcyARLPZ
mOcha+ilbHhE9bv3KsV07umFw5AzI1pdyJzpPLS3c5qNFqb++6lBvVoQ9rL3BbmR
iXHXvnHb8EnA8zgdjp2lXZYD9gWKNimTp50S5x9C2F/FDMoghw4hLvevd+o3PaiF
nzehiI43I/iIA9wC4kDdxiY3ikd4eMGL1RWXpNHDCwzqKlP7DS04hdB4BfF2a5xP
ixihnX4nEs7R3wxjT8oH743v+Sm+37Sv38YX7lC5wRyGko6rRkICSWr8bFyy9tOo
ahdnI+4ue8Ca+CL98SqbbLvMXm+7qvaBU61mJYELokgarrmWGt+gtjJ+Sj/Cg1Oc
eyVysALFCMt8RuP3Yn12htfnmuPuu7zKxdgEVyOWoNybSz3aqILM3crTiZ0Xu9Uy
5G8WtVIAp5YDgV9kK97SoHbXQUd2Bvcf2DhvrNWiwHCoq7CtOc6P2VxGwLY9IePa
GesHTymypBGSL7Adb/aizRS705leMOBRGsiWMHkHrnaS4f404RpG60+2cd6P34qn
fygTwqYsXNTq7jLSt2dAuEk1L0/H/I0uCTtlUa5USUWlcVxSVzSPKFNiTkOgIH+9
gOOtykbZoWbMwjohKQIGshdAaRka3+2/fMyDBMpzBSbXzra0mAq2NNPcV5gBiVT3
hLngysxXhRZcuLBIqd9my9jblgdMdRL6Q/5z8N2ntxQ2uKmcQQ/6fnMktVhS3wOM
us5ShXyd7U22vvPc9wJRFjzkiVg7u0Qn76IbX1rDIIZEdOAdFrJdpOoJgXi1ykJT
TlNol6gU4MyqXe6xfrSxqtqFt+IsMFSVdZzsxCAwmaER2EIjY0YbGnc5h4oiV376
kjaUSiDBcgmUk/5bomcKGQGJBlEK5o8b71wIE3jN+JLu2rbE/hWOqZaDvAFOKJL8
tjzsAFptm4z6QBpB7F5efvBgreRkxduNhBeh3VvNLemtszNzMLHoeFcsziFkOClP
ViNlIqeDz/rgGh9UOdmVWOWFhJJ6dyzja3UlNwj1m1pJQEAqMZTAgz9uGQZsspma
Ud9zoCfGoQYisGJc7enILO/BeujtN6770MG7PSGowtDLJOwJW5N4DvC9DcGtzAWU
awN+v1shwMd3Clf1x4jC89URGnsyUqSVcOLoFulkGpjDHEa+/4RtYV6e4vgrDGTh
kqmfgB0stSzSlkYi6xgstvdlH+Na3uWr1ZAtnLXtp3HqaXaQFcK4R1a0VuDYAdmS
yZWB/DPNpldMPY+tj7a3Dv/XtgpSExmAKCQqHLhsl2px4YHlM17CAnTdm5hwsUmx
UIf63pFrSiDYjMWkg0XE+yPV7Azm+u3Jnz05xHvjDB9Gk5+L72wO/ZP+ARR1bOgp
Rls4kJcxDvgS4Czl6sZEA/aaBsnzEFbFu8L0wRKlITbj28+YDdEWTuhAO+d8W1dl
BmPe5q/Y9hqrOCFt1L+VG4taLFKknTJmrsuGNRW2pNrLajbI67v2wdO/Dcnidho6
UNMKD4FTEX86ifDVS0Hit0NjtKB0AhP+fnUXIv/cCdhN4AzCcUwperCorONJeLu4
D/jMkkL18mC2Gau50bkdFLTYsz168PaSrsrRRgvsY8THWOkyrN4zLf3NVoB46dm2
pWoygOWL1sp+u1QhxEJEpT4YmlyMkyFnbG9lpL4ODZoHIRwGvGeR+agBf+vzZKxN
p9UzQQOUQJEhqb4Hu0jK2k1k56o5q5mY3ISy2OC3BlxId9c2kRo9mbJXN3o7FQFr
ndZddhsdwveBg6PfOfldwQK1ol/16sLUw9P093ulzFFv4a+zL+RvyBFUkmeXcKhA
L0jPMmhy8kVXsrRazmvHCY9shuuGE/fSpG1xJ5JROdTHgMgZnBnw9mKsjiQbNlo6
4CrcEuAVWVzzF/IB4ecG7Qh9kVqZ+Sb0a6MI1DvWDjPklbdLP9VvHYQk/9qNLcp+
UcmvDLwjDCATydRFERMmTP9FH21WDQE9MbQdrklcGtrLXOdVd6DlfIGL7EEKIGMy
ENHhAuypDYfvE/HwaObioUY/QcDH4oV3bbo4IgbXLAYxck44qnfWtMXiKVlv1X5j
HsFkNQSBqdsdMR23BJgyMr7/cFzRyhUu4tMsMU+JaFFHDOnh/Jjdv5jdGQQFvvQh
FwwlGEOM+ZvXAY1CTgwVZkaFuUPnsj9ow4fFK33fRd+ZOaZsmi642daT/0C3cEBP
9Bgn71h9VaqxIYrnTMgsXkmNsqIkF523cPwooD6fDGhVSgKdXgb6SHriYdDHh9MM
GBbwFRu2swOiOqCKdlsaoSKHljvZSyy9Zs3Pu/Vw1+obkVkJOblTnIMS5hJkkgt9
tGPItfV/BjZHeuahXwx5AOxndvCs3fX7AupdKAahffvCfqIGr61568MEmJtcQ+68
avO907b9dYH3Z9T71zOXoLw9SIw81V4Rj0QqMbr+uhCMYgI5K/MRvRfE0TPDOu55
cQNcvWZS/YqFfvxazJ4JieF+GV2eWe3tr8A2g+WKTElsM2NLgUitYKemcg0aTQ48
VSXIyhdkY9olNjzBvPk0TixYNqaVYvTCl9tzUBgcgd2j1DnkfFoseJEa9Ua520zl
jsQi5QeIxF84OFO1nz75g7vFCDmJhoB3QTJVmcaZf82JuLuRWoDUWqbXmcDK+AOh
V5WT6cxd9tF3+7SZak46yJEO5QELSFE3yp3Mt/tk3m7aoXkD1pkcUW0VPEC8Ib4x
r9LVhdyctiYIab3YD390MXX2793Sua4ujNjfZDVK9jQ87rG9sDHu0MIG3K0H9hnP
vd4YfyILOXWVCUHRzqmohIZvcxSqinmdzEr8nnHbJF3/LJv4sgdfV7L4vgULJfFK
RQKY7bmdc1QjPAm/ctiF0x2dDGCSyrahtW82z61i0e/ROnAEdnXLOK8KxITywR+e
xxuWsYM5p9DcxaCpf/EeWhqNzY6fjHUl/X7qm9RPtO/vWAm4nOjiuPkm2OlrhA1U
prKZVURZFIBNtAois24yEg3Jt5RMZ0biRWkss4Cuae7dEWuyC3qUQp5uh7GacNEj
ug+G3fHAUeWOVnj4rNPM9DDWtuhJBG13d53J8YI4b/RaCG9YPIAn84cqQoKAKdk+
jd2Jg0Qy2zcHeMSFS+ydwCCEMz528b919dOCUn67gYQ+SPXUsEWbUG0f4Q2RGrOd
T9T4B7EfNfl8RNqSWsON0T70ydFA6zCzPZkYYLAf4zzALXcA3o3x6e8lgDnvnHs3
z5rgkjGZJSP4cFoTmoeSVxHQUM4PbRev5xqX3Estq87H9XN+a0OkXXvtm0E4tu1n
mtXGIJeQAcRLrrdYnnfrq6qMrjZGlAfBw9Ji6dZA87bWQJt1EprstthKL5TOMtf/
c9a/z6thRR6SjCX2wPc9UQv5w4A1zHfj6P2X8lhLNIxAO3aSVgRKKCsvO6QNRjm0
yG9IBsf+6H8Sba8NcABXYIjQHR7LsvGpqRLKXiJ2or5LbnYtcA0Ja7mGqODhyHbR
ZxujHDBC+s3mRNNnoaiLWQNG2S3kTvs578jNameyxXtc7I2MYjlo8cAtCpmlafcd
P5L4RohKE2bRnqwsYROzH+xRw2+84lNiX5FQwbMQs7lA4YRdB07SF3qDkCHTucWg
2KobvWSkf+7niBtzKTvDx6Eb8XsesqiR6sa4xQBZaXlvtgKF9KsH4jEJtzqZZaj6
xTHrw8dIauvsHvJH+R+EvpbqPNFvSGBnSh3k/VpTglvpc22gykOoUYKs1igBlwGp
OY3mhfQH5Y+RqCH7JOgpF43l71dxe1zyJGF3HfKr2qRKwbxaQ0jxcbFfGyrzF5EB
SjqzaCQCaHhveb9juo7/aBO1treeZmGMDsC4UxGf7YVd4osIbVXnadOL+gudoVd2
7Bb1XBVWKGFn/f6/hM16b2GZbGdnfYvxxRwgn+ot3l/XCydLkZmyANosajjvn+j+
F7d4c9jMlQ3ZHULcWG+wmivCa1zdv0mt64bRCBro13lQIycebuw2uH5AuDs080tC
bSaVRFUPJc/HN1g8WNpM28VDIsLIwIhW3XSmVLkO1i2dhOLKdqx3Yeo6Sd9ofvc3
M3zPztOyd0ergBAUGZOlniOqFUgtGaanx7WAAPBpF6XKNOwxf02elJ1WzjRkKTC7
3lezqMNS+1Mmoy9Np+tx5ZtviKl3rLIB5fPBGslLGseX+Tf1Ss39MJqESlgukrPR
8n3ITAo0zKBfrziISNXGkojq1N1h8g7DtvOrVs+nwcO9lqyLWrb8WyfH2Wx2lTdy
sbqJJwU8fsXqUQ5apz3gUx9UPqpmenGvmQdI6jIUcL0jv7xCvyK/Ge9ld8LkVhp6
VdNecmqHayYfUO5GxXjq6hMuA/oclD1sGNVsEiiiWtquwb2r7WH/BoaKn3BKoOsd
rJoS1cm2se2k2RJmDfuLT36AVzvC8H7cEBCoBUl00AhjVqWo8sEh4XWiWbhs7yul
o8Ld3bmGhgVJ2Dq0SyJxp3Roodp2MsyAYFdtWZR1d8s5qUcCC5tBT3z0Gc6/Mmyf
LKbSs4NblVr0mYGju3tVXOBAXgkyCGw5gyOeJ2muIbN5BktUSnjPQ/XDSpegTCEu
Ecvo5aWMBbtZwHSUcXTNd+9BP9YLFwajFNyLZ8nJHvKpVBhDtUwwcC0MLNzjHsEw
L1k573UM1GmSYDXIsBcd0E+lZ08pvdnx1r4zFgCuTn1qseVJT+P9Svqmjoresvls
eujRJlTd/wXzIxQbiaEzwdIvBlkmlxWhIkw/w9pqlVt8PMZ/cn70mAQpjTLORVgZ
Yfl5EBjaTgwldYjeYJRwbjwHlDbzNkFi0ju0D7cTbRTccRL82GhrPhcgq63pdprn
tnBIu2fo1TCc5j6brRce+UfUrn8kww4FCY/Cjtbk6LHGzMEqJqE9cqZUtOOoxAUy
r4baZF0P7gddWUH4clL7aHTaWx4mQUyu1qNJl9vB0bi/HiG+VMcs730zk1HcIEP5
84PpVgm5q7YnuxjrFdUXrXOzCJIE98zfWxScrSBoaIXmzg5bZqI/IgaQu5F6PujD
Bm3KWSk6ffi58NSblQX4MH4YZ5u/xJM2KAfM5TYpAwPZlsVCjIxgWXimfrGnpWMF
PCXL+I2HB/Gjr2Qes5OZ/hJjLcFrF35vOBKg5Ul8A+ZKE9uged9M6X1L0rgoWvo8
NjZnec3Pk6dpCgNIlsTxbrlqIx01MTn4S2k95KveVRGv26rxBwDFCpzAvh3C2Ypw
VGE8hAqL92JOyUZlmB0Nbk99DYlXNgJd5dIyHI/HJt3r5/uB7XdqotBYY2fiQ3qN
2JEjZZaFScgMvjJ0fqOxpm9c6tW7zsBhbYxsBqsyn2VcKRrCftP4gGaSEtLzBVcf
HviYANXXnc9L8fQ88F1zoAKuAm4eON8wLx4FOgysy3Iq1dQtb3IUUTG8IynArOLI
Yx6aNX7h5jStqgyfrc9wgukshR/W4yjrO4bO2hH8zATaMCoUgR6TZDR8+CkiFjel
AOmROS4tmKwr0jrBszgmtMNELbbhh/0gQ+GoyBEYkZWFQLhb1q63BUJhAYLQD8Ds
RcOX1I+No/QyyEBf9UdjTyUeetTD8P9DEhSSPw7Y8ibPzYkvYx0g2aGRbg5uheFJ
0M1If2mr3CPSLxVxYPw4ovUs/2HN4PRErmhJTRkI1W80y4kbBbXEdhfQpW46AOyL
MT2HWj3WsdiphrBmD4iJQiJThnyjo348aD35zF9jQo69KdNcAkr3xmHtINXVorsY
xuaPUYJ+GdFXpo18wSUbKDTPrViZetL4cdcvXXdXD8HPmhNkDQvNH3JoYunrhCL0
E2vyJHkMORto3pF/xYHON4QYq3oZu1yzZpS6qkLhUoT+H71hnm0DC6f46hZZ51XF
gOi52ujQu5sniNwWklkMvbHXGFzjRlXXVcOuTG5EfCIGwc02w2D1aOoxc6RGoFiE
+kRRt1lH5V6QL9TZZqRIV9eDnEPXVrFM5rc8YCQeTA5Gx2veVfH0L4V9LZw8geoZ
RZU5tPzhsWcqxKE/AChFSBXbfrOWYBj4zoxjLQoznL5cGaYcDrQDmg7fOvMnhMZ6
fXg65q2FnVPQ0/aKHpvicwh9uPWVBOlSbmvzmhWU/Zig6Xao9aoIa8rSrbiAwg17
ruWGjRKizdeGddHtJn1jDh30M7g/JU38kwVKpQ4AzGQoFRM6HTDbRnTng21Ly2a3
shjRxR0Qjnb8g+elFO+/42eVK8XbvuNlRgcuReIqCCddkXn7hOZiKdaKff9yPRC/
2+tBHwKE3VUZ8lj0HLZm4VOsMQ2NYyf5zdgehRhw/DcZPH5VsFKGrKDBOsVsxH7K
/cQsZa04IUEIGjk78v3vARwnQy9GhQ9zKjmdYq3A51Ledx9Bewi7+w7MrxfF/VQ9
VNuYH+f6k8lG1XY6simcXKrDhXwCyw+D3/KMNZtPlvTzYLmuZNjNtZtX003jdYJ+
EvmSO685A8zgjnQPPc9Pw+D4ovdwG+BXXtRgnywNGkKmw3e39xFAJbzZjd4tvN9D
yYRjwZcArcmgocRKjP+AFLQNDJH0gfJxygZS9tNspad8fd39h/tTKyH/UcnUGFgu
MoV4nFSPs+/tVQJnV5AEhc6tF8XOM1NhIqG7DOHQ+cEaIJ41Nx1ccskNlYR7u5kb
CB6N142rPBrdFEpifhek4XhnwBV3/vOXVm7m6KEBCvpr7Didkku1Wnq9hNejb8+q
CVMJa/4r+cd07f+zfcCCxIR3FuQcQepnQZY9QNTUQK/TO1ylO65bwJXQ6oQlsJ89
OKi1pSIs+KGX1MVJIAHXgcKBMuXIGOZXY6Azz6lSV5c0PiJnADkyZLqKCfKnmlr6
VlzsAWdswFkrej2Fk0dZfRLwEfT20//AGCs+MUGKW5HL2/w+0wDpJPYBzO7yjYX9
DNY+0Oz2WotAw5uO1Jyval7xZJkvliNnKE2e6r3Ea7kqDd5YJlbQdFu9DM48ogxg
CRUneX/iWDK64ATI7Q/idX5u5/shz2Oq00rUl/95JAPOkHxx06j4SvQNPZqugF6a
JatJr+hqxrN7DZ+GPwqBkBMsnQP4ZmCmVIKdVRd6hyj0619zEmpxajZGcBckdxsc
NJjZIWeXJpsXd/RTi90Awi/PKPz0s+RKREON4WHphv5eKRPWWQGc+QLRESYkNDlh
3UHy3jgxng/zkjXj9qySk96a3+eO00Dma5bg/YfUxJXjJBzcsaCqPRVuE/oHa/OM
UQnshV/60AHSmq0oLGYmy2lC6qETLE5dSWmWPg2QuRz0cAE2rUMEvgCwH8ALQZn9
B3KAC4L/JOVN4uBOcKQpinn7m4T05gLefL1gt+qjcFYIgxweGAzC1gpnUfSn7vbW
S+4IzHO+BMbSCSgxTLeDAFVxTmNPV5ArwdTV5ZPgmBYr3AJF7XG8QRKBzOXNNBHS
GPkvbogYq/rzfcLsQDDWL/fVaymxeN0qpLItfPmWq9RBXXhj2mFnGovc1s9ZoFct
3pU8d2H/auAcfLU4GLjw0b2LFqfhf7S2m6R0jcmdOu3UXzUGBNqwf47ADcuVPupA
UNQnBpAORtCm0T8oMcIgx0pm+6VPBOJXLBrT0/CVsS1ZaNs3V0XBHnjAh88QQMDM
WA13Gq4koz08UD6apOkjo71578ERILBTxZCi9jVxkCoPK1oOyvB4FUJGZwd7BgAt
QaU8eJR4o8gKfYW+jm0tqMgLQLj08hOm22rXYptr2Mrebu5dZEfUJVtGCGSMC6ax
4DqzJt84cTb5KgSgKXB7GtZpwCNNoBaAS8mo4QxR8fPb/ewcTgoedDj9k019IDip
GCzFf4SofbNN/HMTNyrSGY4IgN52fh0+qi9wSc//rjmf60movjxz75zpqsfJMVQl
l3D52Utf2ROrgY6mJ0b2oFhgl2+otDcSub60MNFo2viRGpT4bUhnTXwGOB5ssRg3
sar9yrS4pdsfjIundUHcbHamiARV62wFbu73eQaR16g2j+RVQWHcew298g2ULhqE
oLntzWswSbwil0BgiUn/+eoXRWg9lHaGf2bZ7x413szjEYr8pT8SJRaIGzw8kM+Q
ZQtvEMauBRSeQgKIlSEaRCa2Q2reA9gJRoMKxXWRlutMXy4s+4h9gx2rqfDytH+D
WTjZf6LouK1axrnHJZUeEguyv+GP3ugEHvsvTyP3hwbqjpH++aeWIV+3DEwVBqtR
S2RphBNFFcy9VI7L3Q3ryCCWlnfpJvgmh1tA2wNqWUN2t8a8iqcAfrmcTIhiizWc
6FhWzfRpmaR185TXBQ7SeWr4cIDzRZGGbraaZmQQ4a8xofNqSXdE1Uf2sC8D81fW
3Piubh1G5quzCU9QymCJT+jSyawIknjFnyaRC4HLxg0I0DgIINmiiAfyYn2xaRna
l+thPZ6QZxFUCEbgM1t4psQnd06MvDLOc7TNnWU+KEn3xU5F+D3yJFf5q0thrXQv
1SCAL3oiWVRR+lPO+7PyfK5/9x3t3KudrYJqAbz6lS95VpWhuyFyFfPDoN9T0Ltz
X0N7AslmlEflyetSVq/McD0F8/sD8Rygc2+T09xjr8ItClAvHI2cYLAWoljwvuWn
Ch4bB7/c8rNXQEjo0UP+Z9b6GtduUD8PVcgARkY7xBGmQDqZ47lW/OD8aFi9N1rp
86C1nWBZKPyYLKVbWIvB1mLnR610x1lBNl2LM3N0nmS3camYkFn8YyPicFZ077Me
5D2P+DmQbYbhBlKUsgHRPU50Bb0h5icSpuHz7miJJCJWGwcbpoxOerLIlwLVBYLL
rmEmTOB/gRTaCdT+rJ/cHaXwvfrMuaL6k09lsvGfUkbKmdi/ZipniOXA055GUFV2
f6CA4AuFFV+N7zgVMgcVGF+cxvA0E+loxVPjZVyt9EKbZTkowa3eKfp0gknjqKuB
0sVaCHfwOcC46QNeMD4OvbcAyPDF7z+gcZYxUajCZ5t3tVF0yveEQQxM6osb05+a
lpVsOOfMtRt7bP4i/Tw9oDMYlsM5MGgZoBBItcvOrPe0c8JiXfIi4uJpdX+HtUUb
PzXyBVHDyTV0aD3VZkB0CPwrR7LEMNyE/H9FSkfuGv5pi2aYzXyByY2xyr4YhiOl
oEkV7Y/IZ/tsEs9/r554mJc6v0iw1ZE/zsWFC/PUTJN/Bc0R2sl0G3QPG30Ma0TJ
gp3oWquG1GQ7qq9vywQIgy1pFcsrM8q1DAXdq9NFO3sNvCk3HlPgc6RtgUgVxxUt
gt8xpKBAeKvb//e1K1v05GvMFXFYHWJedL6efocMuVLSYIalMeVA/LrJpswdr4QM
x0jsefE8/PmJlH0MfxtecpgFo7lxrRlAjSAf6KCFneU8/FNe5JKjl7JIzBMlFxKW
L4BuiC+Ezb91JviByNF/yt9Tgmntd40X5nCaXBKgX5NxuuTFmWyPgCrhuxeibBGw
gl/8tTqb34/onR9ZCKAkcUwTgmY3tZCunDdjChjxPM3GBMr/qASxgfem16VVtg2S
ThN91/BOJCpSA4d2fyXR2QOOF7qOYgpgZiZ7oR4KOps2enkxSBcvRb04aZ+WddfZ
qYZbEWu7Mn0r2UiJV70ytriNzChyHBMCyDYSRT40mSl/3CtBO8EvC2KjH1TqfGHI
RdMsYPVn1Zj4chd4X/xC45+Yxi8NBWsbTfCRSDNtTIXnd/svgOz84jQgXT9Xe5LN
eIXqSP/iGjUfuXD1TK+/82oaKGlxGBkfbcm6/V6XCBTm8aD+ZO/SyQ+DRACT+qn3
eqQLBVZUIk+apIcPwDMpa9D9FC+RcsDuUvAF2b57yaw86Kky0BctfFlxCPtbvT+j
M9DhesGR/Np514GzG51fPd84zLr4XyDxJu6QetKUUl2Why4S554AwbmXougde9SU
+loyQGVPZxxXUl678DnrkMplsxYYUCrnkbnZzdiBFCk/kN7CrWlVddX/151D4Ua1
6/F1QFi2h3MdsXu4EBeIcNYeBWsqi7/cw13Uutwsuw9D1HF0IKpE854X5cPbl/0X
2h2H/9PwDPchnoN6z0oFb2sLlGOcirL4cOPVii7DyRe4c/IcR14hLillSYlxQe9d
R9pdPXjiWC1ZN2l9dW0clcNxIXbQ6TvlUDguenK7WOlD97M+YnX8pabTR2jQFpP0
3K1dXA4d4Isna/VJ062/uQlMyKiCroTXP8dqJQK+2iO+6RzrKnYLMTWZBq2suDWK
V014Um0VUuDzxtWFSfIeziE9UiahLJd0MWb+pKsRYucX7BHFWv/bQhsj9gwle+Fc
vjBFXOIFg2iVwZpGdmLXfSDWuq2AKxCbL9wFnY7F1Z51RBVQ22IyaTP5dF7cmh60
V+dw755LMZpQWsGZ3Dc3bvTcKrQY11HEb9Px75Hd0yTm2XgcqsBq6eXJMD432RoL
0g8L+ZJ1WkXtOYSrgRzAs7w+y18KnH/O1DfKAn4GyBBR6f4eeWgyGgxtq2I9ceQJ
Xp1WUVzB3/0yheFKKli0LF+3CV5peaSES2/SbexFrwr1wXwyxUGrryxWz/LGuVVf
2KtCME/jtLNc2keKprPpapNlZOPknC4D/kof44JXNCHrgRpb7RplObsXsRhwndaA
ikRrQV9lsba7pzVXU+pXqGMph3DXHpFXO0Fttxl2Ihnkzj61o4hcYGDK/t5KizSQ
n1hVsiwgfe8H53kc2NSf8RviTBQO/3tQhCtOU9u2xEAUpnU+8aN0HgiUe7Aih8W/
4zoGUjt4euQ7llZdb7SpyEUnN3fHVdTgLbKtaRZni586jYfpzinCiy3RlhwP3XQY
NToKStFxEXbZ9FqbxZDyEI9FOwdnKNYjq/HHt5nT7np1SYG/eFLfhIDRlKzCpmhS
So700OQ3LUYiAlSgjcmdlfCp3+2nMmKZ4FcYmWOGGHiQR5yrp1nllJOKuoi3cF0B
5aI8+gP0cmOI+KUtrFplbDVJ3gSXfGeqURpYjvVFnMQ8y4XZbm0prY7EOSc/uoJB
hjxhtCldX60pG4kw/NR6sKGrxprmQiBPKSEVVf3W+iOqB/m0UAnG6WrQmEDe6wTH
zzgmrks6gCoyyE51VfrgjZbzhJZLJ0FbKzeLuAfkakdkGF6RHua//ndZRDCPyEQf
MCDDlp4DNkn2F2R923p3JWjc85orF2+EHhfFGVb5EW1aCvp5tMlHM1Uk1/7SQv6K
4WSDdddjQe9FOM3eQkSoZaAz+K28OJCf2tL4np3byecEkYcedRbPdSprldNUsov2
iRCFnItilLLENR1Y0f+SOqLsie9T/cbNYadJdom9pn5rcogIHRS9YRF1hoTkC5dT
ifS9s7r2vwgXGjws/RYzwevjpFLMqLHHFfMEIcebxPB4doFJw4wLD35Xi8cxWmc9
FRUX0fuZ3xZSfmkWjysLlIBIHTnGehDdu6gTO9gf9azYy6SQVU2uEOLfMgEsfa+W
t4vfBHfJFPdk0NWxT3lWRBA5hlXUbLDrDciffyEUdDXWawg1xXE7O7wd40wUldei
jQvf/hv/p4dDsDgxuI6EgJJ+jQAFMLZEb6kSqjnHbRnojd0JgyteUq2JDYJLel1l
EA5VQs9Q0DM4m0hrG788QkYeXkoQ+8jxYeu6+71L7YYTxOagiD7GBknq6QcgjvvG
f0qhyfhFrOLsIFZqI//w5RkxUBmrR40qLad9sivE1/P2jcRdwx5ecg5cG02gXomG
h5JMYnKbUdE8xx5d6Myq+qG1PXNFqnRf7XkLOkt0MCaQ4BsWzymZizjH/haWalpJ
3D8OBZi+oxPLA7uB1xAPQl8ZAzYASNLqbHgSzFe/ZjDFJr7rnVxP97EXvO9QHCSb
vXVXkIPmZpLqnsr/QPnuNmDTu+pKckZI3jYw7k5hdaVoSqT30PRMnx0ENtwOkOV2
chr7GQUuAnTxqB3OgicrIjqyuaKN5MtH9+5MR4e+46oWuN2pkY2xBaTZ1e+1F050
AA2l2SXkz1EoBkND/MMA1QAd8Omkmy3jPcbfY7F4W9IqgBE/IGQ8vydIi2w7RPlx
qkA7ZIF15DYXknJTntJQlKHiUhd/LBNkXkfCeUTTEqs4iEjybVe2hfjEawehFU+7
upnntO8NNP2s+k1XFzgw0OCBraxBv9q4IMLYVyNiDUXC8Vhfg8JQpSjOjuU+Qg1q
wizryFliZhHGzYbSraLxKWaxouxzzvJyXqRwrBlcBaZbSGWsw2LmxkRAAC2ufneo
vNhLBc9Cydp7+xvzzOEE+GVir80E17QTSOw2aDPwYxbtrawdYGDZFXp9iCRLBWRd
ZSanFvtQIM/fgTQihaq5QyfTH1k2k58ZzdHPizTJiD3wm/Fbqj7XgaKJPTBLpYlb
A8T14Zn+ZAg8Qf04MHykHa0a3tCMzElDn6LJc++UZHQzHEvvfg1cgT529bS3f+f6
ffRzlFaw3WXbB4vrqJzdYBKkaypc9rOgfxiuKkYHFfny+XZc+KpGoFtJy8ingo5P
Ik2SCeKTAfl95nj1OtseNc5DFLfePJuMpEyQJdQV3lnrdubpmxaQYsYNujsQJwMB
FiLr9lhY/V9YtIJPmScmNEKo9ZMM1cR0Mh0B7OR4QW8zv3pavCNsAGUeO5I6vLtt
aiB4RCR+ZDJ/BhsXHNMUwn2cUxShENKKDLP0JWMI7H/BChxvFt3JTaQNmccC+8LY
Znn6LKHRcJCQu4EvMX8vkxo/Qz2QCcpqweDdtNtVIDZizKTRfh01X36PcY8vmfkG
9rx80/7CKbVwHxz01Fp5z+0H8oh2gx0+WAAFm0luTM3GGbP8NER+246ADCmhAm2r
3VqjtNp9WVnGTbL+j+zsOI+q5j9k8JCxXR3VzIjHffadPi8Rf43G46HkXWPYZ3pd
KydEcDLVsd+/S9YliXfGhgMGpLAWivICZ5EV5f0ZeAhMUTewXmeMDM5I+0Qgz9bD
J4Zu3fp+RQ4Wo4ILaYt79twxW4GjWoJuru0p1I2eHLA/hA8ZlYmL97bvisInJ8VS
jwkzBXEgiWq9+zV2Gr+fkSzKvRdB5tp4BTA2QEQ0dN6J+lRIXOEYZvA9PHsJo9Kh
yeu9DLe2GRFJW6x6z+JGAqwvlzZVvI5zeqapLvW+873B2NpbqGLHRdLTYYciWp0w
EiceHRAsey39C1BTHkmYlrof6k0Fn4j5cFxGgxhU28A8VInF4fEkxErdmyzi/rRU
5h++9MsFK+TbR+8xi32vmpDX3x5u1O9Nh/XYTnW3G7WLwFmuu+V+cdDM2Fc/nSaH
VZvKKHgH2XvZtJnpQ2qLOzXhlnVycZrIMlJMng1KF89puVNQ3bEB7Kv9kQmxRV3Y
OZMnKkMA2QL9GDR2i6a+LUbf6z1jmUEhBwftWxafVVTul1yadsvjKFTrbhk5Scl8
OI2Z1b/5HazYYQw80rDezzPIS5c3I5Qx7SfE9nkcAYtwT6eNu4DMNcXkcWhnlDod
YYQ9uAiMzVtu/lgRxJfUcv3GZ6ld7tYjV+RZ5koQ8MAVqIMMrw1jaDzeRk/DJrbU
FaVJCpQ9Ac9YEqx0Hx8Kp5/wMulCoZ4GaE3Hu2VXbbgbGEcTZX5gKLiItgl4i9AU
hCF15drZ92AdyMByoC1MPfTVNh/ogXVRUnSOX5X4iAblv9uzoXAeHIIjK3Lp2BSa
vuH1/WJ/JTKkEG3kNkWkgIf+MmHV2dTd1f7ZE8ZSdnMbgQqe6o6CJvueAQ+BiVic
80ZWxYlVRnmFUn/3cYjcDLV4h88DaK2T73eIRXPwCzYCDFRWXeatyQE+na3MmM5A
PHz8q84Ml55XIwg0FWnQk3kGPuYfJczHl4hcbIsLbL6NgjBdT+Mw5q5HzPh+sOqp
M1lzVYiyZpSCFWut5XcGHg==
`protect END_PROTECTED
