`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p6tjK5tNr7hbDX5q1io6K0t3A7JqVeaJzmgXDJtE8Z7zuBSkXboBuh4iyMW+2Hnu
BSwHSZrSgnpSwCvNbLW8ybfoBAtQHc02bEV9Jf6DICMoXpK1i7G/pMgoEUID66W2
14nBJLqMwxpOYuD4nY15fiOtxfnlL9PRXv2t5dsesjdmeH2S2fm/tNKlON892QhK
iZhGMuDSN4EddE9VHngObmxKfLNdsFTJCIhPBrP1VLUhTwnJ1Yo9YvbnNDCtwMxx
5OoAiVZ3+yT98V6yFvWnsw==
`protect END_PROTECTED
