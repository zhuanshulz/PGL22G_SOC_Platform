`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ubX0e0HoWX78xxtF9MMhGhJlQ58xgHParr4xe7jnfycFhP7dG1wD4AC/oBeMwHGd
ELyhAQUHXocLcWS6dsp1w4xr3DSYTdsIE7ZS7+VrT20/rlzJRWP973YEv3Wm3pkQ
gQhi6lkWGbf4oHv0jQ8E8zZqhzX++TqLkaochfb4o9uUXhWR9E+tCUN1urFxjBvj
8QSNuuy0dNm3oK+3GYyi9xyH8+xbauE54G/cnkqWgRKsb3ck/dKY+tMTABA/WpGh
1/vpySaDcajSQ+IKK5AsS/3+2E1r3t2tgXz+diQ2W+Q0KWXuuAMUcbQjcOXIoD19
p1WeXCXVWUnsvd0oQ5eOCfZqyGYpmsJkyAlZm4Ohwm3IsF98LGramDe4IOV6WT66
5lDBpNQD3AlGLXlrPrQULZHMFhUahA0m2HfT8JN++den9qgb+VOe7btPHFUpQCoL
0btxn6BjX99U2qUnV9bbwyEPikerie13jdUqzgeShcuD+fiDDPy2TPo6bdhKKOgL
ttssMZ5o+TBAMnHqaSdWyAYtloJe1A0laVXygSUs4gyx2Tqf/6f1i5eecE2vyH89
zdglQoqJTUnmu+sMCJiLm3plpcp8DxeYSjfUeCjooSq+2XIpmGhRWiUh+C0DNfhp
TKCF90iT9u8ZtIyUzhlJ586Ca4I/8gL2hcyzBouwp/yjcbKJ6ngZuEc3jBgkd2E1
Gs8xVvE4Uiny7JVTimJ5C8gCAzqX4EQ0WtRsfVca0trxCJr2ZWlLgCxbmmNOGRKU
`protect END_PROTECTED
