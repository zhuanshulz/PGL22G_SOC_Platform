`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1mWtDJMJMqO+5aE33HnsKNm4Ap+vqqMI5hhDaN+d7Z6Yvw9rUZmrBN2l1PNKWRRj
wH0nTeXGqT6zSic+Rcr211zpY+2urGqBoLlWva4mj1Ly6ITeB/hte5nbg1hU6kYl
HKH/JKsRHQ1xj0yW2N0ZhgPU2fdRpX0e8+vS0uZEtDt2vf/oixpvE6IldCqZ58cD
BNaIYqtR8tqjqWgpA8lBiwILzQT6pHnUhJilae0bcgjKfHIvVJHrAbok3yCRhodM
pYt7Cr5cxCg2lwb3ALvwQ3ds4vDnqZCmL0yw0zmBGRXDo1bGSY/A2EnNh+9N3hS2
fbUN7mNrM3x8LwFyeKZwbFTwwyaSdlcS8nGNmsS1qGToS6Gij3TEmXVwbS46BMKZ
ML+WgyAvVrOsMoMDkSH19w3lTOPcVtHzYHR6PbWl+exu5PLsCsMEQbOD+Y1qiDSo
YK5/SmC3cTbg0I9R15kIvWFkwOUGKYmHP2IHazPUKDd9NSjpAfeor6Cy9DEWuiVU
M8j+oKFszAsGYVcr/R9j2bwtGTNeYwyWaxzskDoh9Lqo19HYBq++6ooz3cEIWWqc
7MnH2yOz0rSf8iaAP3p/xgxm1xtiY76YeFk6lEEqGlZM2fVOrNNdduhSFBHwjwog
vP9dhe5p4rak4xpnWNbhIPrepHqD5863aUrMjc1UIrXgMzOlYg1C/HCX7X5Uwv35
zt2CUByM32Dp6Uz9w+vFkj2QqNbYuiSS+RXiQrj2YnyzXR2kzdEnWOHKMqAqVezY
oNeDP8Wo4DN26FQsRSeL051X+AHuKmTVxT//ZYKMXONLfFeE/vq0neh0sRpvXj+A
mgeCs8XnJuyTrIBb/XCntQNji2/pCRpLoSXg9P0OUkU=
`protect END_PROTECTED
