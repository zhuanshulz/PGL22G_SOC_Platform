`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7ZoU/wZV+tmXkVZEtmXvZXm7Z4PKq8FtD1rLplkeWVHbaoWBs8SQ/OrZHGQXsdoP
fMarwFwtf9EGuJnlpVSSB6KAp3ZZPakLHLFw4uxWHRqBgE9wDMiZMFiKVgjkiGOn
XeBXv5+Kf1WrpYGvi4Pq768OngKvSSW/vSqcaH0vuTCALdH/G+iXWpLrZWcqynIW
5b2NNGxJxWVoHf5MTijRtlmb6810XV0l5pzV7uUeApZ6A3OkMX3hVYuGwGLgJcI5
ul6I1hMEa4N2Nswt2RbSLb0xFqI51PZNZBobDmrxmp66amkZ6A4kD8YUixx3kxOl
APK7pMMCmK6dwtAM7ON36imQ5kl345wZiT3v0/vhcOCSi45nJxoHz9d0GZmFZb/p
76IESjszE0Qj6AsdWGGXRvdcHi0mieBJ/swjvypnrRB20oHD2aRSnHOz42ef1tzi
AKqX0U6yctNW5d/z/e2QbonUCdj9nGP+60IRFjf6nZvywGlb4cY/8xeHehlvIHrf
sPOYyfy7Pmredj4Qvwqk3BAnIeBHTmzZ8O8GkPWBoE7YpnkT6VgaS5xjDBTcsjPZ
QOIJlJBWOmRoDEDItS3zBLgVPgBgCxvzE4i+ZtAT9xe2LKuM8GUnpLkEBPbUTCn0
DIxZ/aVhFUnU68BjeHcjlVsUY1kEttes/0k9yvWo3YzChq1wOokvVufhzap5igA4
oAvjGQ5TKmFgWi3gQHK3UX0kkehX/97osxxkowrO0IQ0niGE3Hih02bdxbT8u5C8
1SfX+BNfQKVSEULuyO4rnkXY42cyyGN7K4DxBu/sPOdJxBKMIvs2lhWhM/ud6MpB
LSyOQHasIotKVScttKUNOKojJOAQJJIZ/bXjhIBol1iDJrmf0LpkHi/Hcu4vehY6
63bAPlrkK2fuhBmSlY7YiYy/KrxJRMDfa1bJ8XmicRwL95ug3Kn77GfKJzz/m7AB
wk/cgOD1QoBgxUax22Y/VBjh6RHA6xR6+nNtLWKi40jIQnbigltVCc+txhRoscKx
U4t900/MhxTtDsBJRX961ETQW8aAmxZ1u4Wo34SWkzLDz/XKIyjLV93iEwqMWfrk
Vr7M15x+mhnX3nOACxexKtkhw+ZBlPFuX/NuxA5boFh8FELBX/Mgg/aQxOKFiZVr
H5+mjptG9wV464lBPVJE61C/+Js/S+WZxiSYCecBXJmmNuzk34/Vvl2TS7OETxIm
+cm+C1RJdFv6IJEf7TXSpIs1UJ1TYVgZH0fbCHePcA1eNZ85nX0/zdEa0q0T+RQP
Xc8Eej/Qb0By1hiHn0pcppd2TIpHFP4ohqaXswzoklE91Ur+2jYhQoKMLZW7pjyB
qS+1si9b4kEjLT73p4Wn3idKQ0HkRnrEGpxFpCNo4l15uphM/5498Bf+6AXIuDRF
rw02c8qlV+c6jGnoJlyCxPq8psFLuklkiYTsl5uYEFRo/TopyBEP5NHzgotOWRsT
RkRl621ekWrAhVq3bTSsHQp+LjqWpggpyZ/PwORFr0H3tzXiKZmsQAeHk26Seuec
Ym1i19VSkv37EGFDo9hBtS9Z43RiUE6/xI5wtcRYG35Nblr0s+BVg2iTz6WtdLOL
RSGiImzYD33eXx5bK4uVNpjMH3+ODl8MZJjYXja6UjY9FuwLNRvkAJaRbxCFV9wB
Y1JLhG4cb84qG/unD2GVRQsH7FWGVhBDvvilZ4pgxZoluVr3kuprKWCH14ARm6Lf
zRLy/eHF6fR8ST09SekLnOwcr5pnp7Gkcc2Ct0guFpC42uQoNHVgAvAKjFv+MO20
EoFnwUB4xxKm0i8yJDVWdseZq8Vy1Djq5lJGPiK8VXedaawoerldwMoz+r8UMXJ4
XbwuDYUmzjAVmH0YHkqsNR4BR49jcEUNOZcKbVnOadQ1epEeFnayV1nOMPsGROCM
ma52nfukkYdpb0vx/tsUHJhAyAr7n67xgH04eCNsYNZz1Tbd+Qr7SyaI/eUrIHMj
LykDzwtisjbcUXu7IJX66UGkdN3iozR9FMaiG0ZvXrw553S3xQ4EYIZ2AxAIz5F0
JBqQl4Dacon8yA09UMwlBbvy2fGhp2wdDC6hMiSxidyC12xGrUSyw+nB/89p/2zx
obek4pT4wqUzhbwi77SbYnuGZLigPIlfClJuzEtUWipsJYFGge39dzMyRORHZUsh
QMYXgdG3Ibx5NQ4qP8PruYEfoWNfVtW8VRK7H/jmB32gGyKLl3nLDWvGWN3bE4Zu
IIJQeIyeCvbdQXsIckb9zGB5fSwyO7k5o4sIjRYqX3lyXZW84nBfgoh6pXKQNPOA
DvpTbXcUPNMmlHr/CU/JK0XD6kaa7I8non2FIfxJU/tSGZ795xdZnUkPImahq7dL
DXzDh1bnai3/JDlI3U5R7jBWif8OVFmxAOmfy3Ldw2aqAXOSQgiXZZWwBumAOl5v
HiloZTyZycbmyzWf6qIMhOdKUHBbR7C3oCU573fBSyG0IdA0ht0eIBaWH4ffvC9Q
tbx5Qh3wnhGT7wtIRdX1ol0GgICWcnKeWWgQTDsjHmu0lBHq0I//gS8uuklRRbdf
az4i6WEQEpaWmKD9jswqace6+JY+0OBCqpplcItq1d33SOEyKit+TDUisvbO36Uf
ORklXrT9Ed/HXFn/1Pe5bplCfJBRwflvTToGhlZImq2OwNP8cGgPz5ksdqjMt3C8
3MSWGbPaEWcMeoF4wLNnKwgC25RAOW+mSBw79Q1qezWLxhlwWqqLA/pUvPev7CdH
YOSu6ITnEA8FNkbqjv0rOX5Jpz615OaJaz44VSrVjWD3BUa4CvFGALLb+jPo6/Pc
F/arruML5ydKsxQU489RYuVNcThEbo0rOyh88WIp7gXHXBI5huvpO7BsgzC15M4M
i17nWs5LvKy5BBcDTTrXNflkBuiZyIMDQDR/0Kt+YSk/t1lx7kFZHdR2FG1Ydzak
iCEeIxICG5xAvU2S/+KgQ4L0qK3UNsNi65GREchiV2gpbktSt/AmDoDKti2ssWsM
pPZXqvwcmbUtO60J5PGbSvdM4HcoRvAzu1zrEIgPPmfdgOyfcrq+EzJTzCE2QdBX
U9j7TgAJn46p25DENgGVQWKo4s2l1iTWTjpovvqgGjUDD2YGldGbzG9LAS4mzEos
Pr8Fym/NqF8rNUWoriXGrOEtsMUpIIZ4acpJmRzbrhdyN+eLNVJCGuVpNQupiN+h
4VGTqdcT0Rm4VmUGeXPLhACM+LfQcfFfENwQoLo/34L0fX+lqJoo5CvdIlLKqxcm
DGA7cP0mwzd4b3vqX0TeUuxc8Tl6NEsMPU6yow477momF6sOXTHOdujwUO/CSneG
Zlml1S1k7tbAykxiXuKimdmO8Gx5q2csAKFwTc4qlHFsh4yHim0UG3RoDgesf+B4
NEmhbOt7ZUn1/EogTPyRxOubO+SZ6/13hLnU2hi88NHBtO4fgdeb7muhgTML03gE
iUtbNplZVsrhbh3YguO5atRMQm0R/gsinx5WbWgnJUgksihLCASpJ9k5jYJ3TmMR
IKRMQg5sK55XSlx3/LU1UweTlLf2ph5Qu/39UaKgYo9cuMCRSZTH4PvHYeAuUDOr
NCpaNa9oA91FVnVX8raz1sEECJneBOIbLoumeLUF62/W0wT+leVFH6aUX3DeMuYc
ylSaZWGyNfotRFh5DRlRHqenaualdawzbYkPztjdKJrYrfvRcRATvEosOpirxynk
3YYglhc5r1wI1AApw5+8SDz7OnObbQ+4ZP1mca3KPDt6RzNQ9iA4JQ5RDvkIIg+Y
1ggC9eKEwjCfmjlKtHbpDrijCgmd28UwLwt+BkIccCtMTLKOAFjYT1otE25dy++M
mHmOortNtyAWSzjS25v+Upvw4qSQLglc1TsrJEq+J8OsJdQz8BaIe+isjoJGeWor
QrlgQqJhTN0JGaRMixYeh5d7IdQwmXaeHSNJ8S+cg94BQZZz3F9pYh4VryqDcT59
n3OoL1Wkx4uVs/8Q7KrAtuaNNSvndMJ1Uci2HFkRPtMWogayNAB+JM7vY9QZ5ddx
`protect END_PROTECTED
