`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ucwhX2kapYqrYLONU/kHtkeLSy03Zz5+w8Mm+0TUXggAIoQQdiarTzubaNRiVlCZ
eARyKDX5I+i0fAHcHSPH/wzP9v7bR99nDWAUyVhdBH8/QdEwzBjJXc+/69eZoUnA
EV+ik2tMdiB6EnIWQJZxg5KEtRNpNOrdVKmamfZFhmYimPuYcJj+zlBqj4Upf7EQ
HqpbgiNUk11ydp3mMhc+iRHql5WhsQtSQydSI37l+fjom1utfZTr3y0uJshuzYWJ
U13pFKFbg994vCOLKmtmlmdgmUYPRRYWJybCIgL86TN5WTdyAJWhKnTUaKl+AmNf
qKSsKfGbZfZScBLizS5NtqiXdiIdS+8wFNmIY98/DirGTB69vPmhcNSL1yBkvgPT
gXgrv07rvAIr6G+YZLU+M5oeDT1RfbrdLli1kEyQxIj3KQyTbEycyI/L/CiCIKxg
iGJDadHuPkksPwGm/05LaC3+N6xOgHanVeOSF++kgRbbXRtRNiI9dO/xalOlFCW/
zN1vTrJARq/VgEzdrO2HM7gWFQf6esxHRoJEmhVDqJBusqIWsh2z2+aZ2JrsSNmW
92g00o6INkD2sK8qg8GkUWLO75Pk+u3t2/otYyiJzJhF82MsSBT7ODoljsQ4y+XU
s72HTtbnuCpm3OK6YuV6efN0TrMYUUv1uvyk8CkLEn9VG1TICrBf+X9T2Va0cfQP
AHONDwOhAPTh2i35mFSCAlYb53qAvfuBA1018B9IQYaoNSw9D37LEMcM6PVlP2c4
8TMt9VPgDuWPM1qjEbBLcY4xXjDQDpe1cJ31O+gXbgEIEzgbrbqiN9ju2OOFb06s
8dqs43hjH1aaEpfj9XOfQ0wFulO9Llq4rUecvgdBQZX6zOSTAeVYUJg91eoJvYpr
bA1aQxO2HYMUE8TcBt2S5TlaHpfLuaRHhZ7Uk1hLmrT+eQcnBmXtWsc2U+nEM9b2
PP8tNLwMBDcYpkU9ruxdKtswtnNe1t2IjxXoX+TtYpbBsXGlZ7khCKMAn/5pcMgv
ZdjRjwr8cfceo/4ZaoiVpaa5knX1KYKeULtLzvw9g+qDFQ5adVcvaePQV2DRKkiV
eNvVNZus+doTwGOykOSTo37aDt3C/HwVZiIEYeF6KTkQNRNWqAEauBgdCEy6L/WG
vAU6riHOi4zFhlGCFV0K2QbelmDpZHH13KX2pIyCxvJMuZPCqwXWaCPZYVf3sHFw
f4aWO+Z+33cKmHKHG7pCLNf4d/ZKKwpN2U6hrz2ft5+J4RmHaets6+oyVaFESvk2
LfHKqsO3ih2w+7t7F8y2RCOugAZzH67MQSFaJduQty3RB7nib2ftAc2FBjhziUva
Clz4uhxB3CEVgcb/0vyrcvCmxn8zBLTff6c9OyIlXTChVFyrQvJd0EIkivFl4JRr
M3nQkpLNW0jdjjB2qlsX3CdmhH721uWauUcqKECdnXf9Rd+lhsa5UTvRm3XtWqJV
IvitslGzYryG4VkV9kO9Xr896ljbQkaniGWBlejP6SOOpvW32DOwEAJVlSbmbR20
obYdemfukIorPK9vn+a/sARl0CjZ+nmI4ov559CMyeysakITW3EihMpZnRBLXQ+a
YZXCtJ75CUCaaIvoUcas5OWzCPykF9yWywmvPb2K76qIptTgrpwnNYH5xLjOsjHN
N2hnKvpB+KLsQHXbAtXtnlw4nkg1im4aoU25T8JW+464d890uGmtFL+2pc0l76aG
AGf5Jkij1c2kiy//x/JsTz2VpfeHDLzvL3d7OV7+Hk502J4dGQVx7tZ3RPl6GVAU
IsKbXl4bpj88cDNza56M+so6ptzFmXvRUlpXMdnzKpetQ8Ro6OS/rV3K+lONia68
Q2Ysci1mUVVLlwsIx8Z/9UQPZ+9lKhcKJh82KsjPJMEvEiQ/fA8SB8UU5fpMVsKH
AU5V43Ivieo9+yNAyXEJEbWKq7EU9094UKwGlpHv6QLJXdIUWqxp1MQ7khpVeEGf
3S/OOiTyupxgabiZz4UdVB+YQSpkzNHfUDzrByq+9AqRDeMDlvytaD3bFIs6uxm5
PF49q4+ogEddc6fCSZhewDNyLC+9Zh9thocSn6uN+F2zDttfbvzNFzmDmltTMGzA
TQ/iR5bwjzbOrE1F8FV2Og3vNwoYzHeys0s7wmd/4mzbkqeKvqIuieRAV3xpwmeO
oVGjQlmhERJDrFf51+tj/B9bCe1/KekpV8jKaKHidvu3URU76kHd2hkJSPKKGbN8
2m+goTo0jcMzj3RKWNUAzbj6DJL73dbfnGQPxX3/pBcttiJaqLl+YD/ol8Vktpeq
1LkEXgpJ21+/KAx/l/p6Fff/01xRoyNZxddqwFzqZpZyVKLaQ3F2tdmhwLp0VOsO
h+AIqnvD2N85eBmdr13Dv224rdS+zJoxmWckDGFYlqCaTJShg+w1ibTUa2rsifgQ
qWPUUdkaSDGeoN/5rZ1RXmSmA4dIjfoz3KUCGC/3kkiqPFxESIBU4odHjVlFOaCr
3mQYKyYL7aYEKd42PxvZeS85Kg+0+JQ4eovFTgypKSxlj8RzR6llyGwBSBTjX6Xs
rGxekAixq5Ins0r5bYqyK2ZSGwyl6naOOhZurOMRcz4MWHxW1bpgRvNYIx/sjdpZ
2veyuAA48OuQ5f5KuII2yFU4/CjnuvVzcJfWBNV8zmyKd3wv0trBZbTdzzwk0z9I
RnqR9PgcpWFvBFkxWDmthYd3Af3vnY+vnVhLdYrKtg97BeoW1b9Mz4XXTODkDkiM
ic5jupADQw+XP8DeCQuK5SpI1S8XT3jKt6DwtnYcaGCh/G0MHyij4qCW5WoDCQz6
b9GuYDVqrTBx264LuLnMOwHhX8dozJzLCPlpcS5S9igDm+Yz2R49lKXOQ/MXRxPU
WsjUlgO8wptKKgO3t+4Ahz2C1frZLohYMt9YSCp6vt1lAblWpjaAlh2EjkNAGD10
eE4JrmxfipAMzWpl8V8LfiIG6p8We6E9mCfttyOPvFR4s733UdjvTpCDtlONilZT
NKi4SfJIEmjA2YImIKL3DqH3fPocz9PCv3g9so6txwl5bbXeF/V4JOhclAEjK/Cl
ywgkkLTymPv/B8Si2hBvF+PoaF4QWfHpxcU37u/PYGT+U9UaL615AasorLMmp8yA
/32nPreUExrXINKkKPbZoqpZMFm74i4a+ISdbs4kKJx2n3FuMnlMJBs1gDjT7Ed+
ojfP082vpe3NyS0ZUNSxK6IS0PV6i7u/T39I7x6ZQrwEDPwSediGmFGnwLugCBc4
2uZwmXUh17C6+B66ZdKHAommsKwBmj4WWWGI1/DWrzZkGQ9uj/TcvJ9GtTKvpKLe
fYeIDINdJT4ZrStCA9M3kvQ+AbVPDKmeZhWzlhFx8IfU1ZmKZzbp7yl/ZM04E/7W
2Muzp723TPUDsEHm/9z8b/QPQDkLVNudPXuVftl1V743we4o1jxEUA6D8wJ1T1De
kngs+W2VqoFv5Ff3AXaI3MVO3fTIboKPvWu5ZrS7+f4QTZ/flGAmwVlcdt7+/HBf
0v0AyuaExGZy4KrNUVdSGSs1TKQW25D5lC/oNGruiKdjoMNdXKbEv6rUL9CtYIz3
lbE+iFB9jdi4yI4V3qHIY/w2DrpvwBb6uZhj0tVwC2Aek3OEsi0Gt7c7ABHxzfED
e3gsgUuX/7HRCKFootf7d8FTIEnkqWafH5eu0cr6g/c6on6DlY81gVuqLB3d54I4
MI0/CVt5Fluhos5reWoQtBJe9oreZ8SXOiaCwJJEtVkDqdhVfHbilJwoaOW3iJiv
lAx9/fwMEHSbYFl62ceYnczadfUGb4c6BVAfPJzcajWc+S+Y6srIG95/7zfp+Cx/
Dyvv6ZCiGXgmrUHbIbWIkeX3DzGwdYBDeZ+hujKetXRW9SaD+otMfhtbfa9aQ2QA
VNtKfBzpA9tJi7knNQCA0U1z2bPZXrqJC6jHhsvmdMq3v/b1a65tFsSwc3fJCiOr
2Yr7aEhXdzudl71xQ9IVJkogfBukPswq9zBM9ylt+TfBB890Xrrh+GI7hbcaVqp8
mLddxWl13pscKp+h1q6JgH7SjCHYQdNNmoa2ZhHQ89JbmYxeyIlActZk/AzO8jxb
UGVBICQ/KxQdf7nI/ghG73UsTIkvNBhLFmllCBEpTIz/PUSCPh6xskXZJFWArTx3
wSx9O/nj+Jyw63ica8YIdAPkEBGMSAsHyzEt3xFwVS5zCNLogJ3CNBWOwQC7QtAg
GEJIU5DZwmT3NNA3I2LfvPMC6MFw4LoVk+ZPtXoN3xNPQ4AHjf48OqJfu2Usg/LN
55cC5jh9bUndY413dep0v0snupLfJxboGohXs5+WL4DFpevMV01n9DAPJZymhKbO
YRCBheSj+JB82x405sibRgq9tYd1HlVTH3mTu1n3gZEiHHzK6PTufDTkNhAZDDIo
zNnIg7fMeFbyTtDs4ZCWZGk0k14GAaDueOXBT0WfTltl/iy3GkDD1+0t9c7H6OW1
HAtxe1cTPN22NZ46tsHRX+quU+u9IqhtAw6hBkqKBHliSdKIc4lRT4Gc8iczVJap
ic1xLnuhMXq0aUEHNlp2e6vm7BkBv1Cyl3xz8kaiFEvgpwJ/bxm4E6vN5A/XYA5K
GfEN88dwOxgDsYPgikYVJosJ7Ru+iTNVYd8epucKt+NlfEebkyTwYK/vs53rmFvv
QT3LQZq3uvmeCArRR3IOqPadSBvZF3A2iwzhNUz5TICbV0+xX9t9zYfJOWVlC8PY
hG4B/KeZXjXEfL7X1sStyuXVxODZYIU+XimZ+sv/AN5cBOGbSX2Bf0eWVbmJTzXU
1DCHjfaXwuvicbJtkylNOCHrsGb+QQ1zTqNcYwFqmy5caR/GJOTdeN12VGOTji4F
TxMntck1jQC1A2Z/pWUPD6x4Q9ZlMuBT/aWpnG7TmGhP3bEshCDHa1HJJLKb6ljG
SHxR5Qo/IetrTRgrstJT5X1/+k4JToXH8F/gKciNZGLGlv26kZh7j/RThVOtw6gu
1WHVnMMQVZDLKmqfWWe70wAWziCc5jg5vjVeYM7ccUyHq7yGbsaBl5KlrPoBjktq
uC+tEZAq9sNFQbEFz6/OGbI1wS8DH/UWUPKFXf/tA6YYkZzOaMAqgU+Bs1FiY+ig
zhNqFcByyMyg7AD00Hm2XvoUgYVMIZvi3VRaH/0Xo4kFQGwxpsBrGHIe1fe3LvfX
otLMmZKHimc6n/I2oG5/EtBYA/LWdHh4x+2d0aV2s8JNNa707cCPH8T8MkHjFIqV
Y265rvY54twz5UJSy3fyrH9IszXnswSMqHD0Fw2+NzboiNilWyTpuEXsJ+9WNXqu
shSLKnTqHMrFXbpYgURsGDRz2UG/MxnIIuSqwzVH20yzTMLopwCEu2AUebInyTLa
96CGhS+zFGJeqwajYCCn1niC1VNdTQdmtVxX/4vkkVojVWHNTS6xOY1lXgfuJfmH
NBCopyIplF/vue83n0/iq4BriLeelnPj7NyqOGYWEnDSsrQoO+ZsPd5+IltNaYwK
N2eUIi0cxHODkE4mTvRVtB6NaKrVy68tsaZU28mazml3FxlGaU7L70ntkx5kNZtg
9G3FqQ02e7DzmviFRUiL6S5h6WzmJRTOSn6rPpI238+0dJG+aSr8J1qlgs/KMr1b
bJtgim68/tz48tur1weQeZomr4lyAAA9uZmP57YQOw4q7qEJAxHrcfY0WYTwP1xl
K2Okz72nMPmtWPoQ91iTtKcmnKimiPfXuP5DCsV42u8eCDEsd5dwWmQg7Vb8E1ea
kW9PEjWUsN2lE/QpxDa+hLl4BQuQSzhB0VdHqgc4vt1V8pjyB1IXA7aarxafTQsl
B7OwUroHSfIUs1b3q3XlcR0SrpjUfgSh1MKzd3nYA7v6Eka+rmGkmzC/XjXtFrFT
aMDekKHc0ERjiJqtkQySpBzgWhUWPyHH8P/vOXEg8BgZ/sDH5A/BOB15ywjUs2G8
WyRcNFb4orU1TGE+Sn7P4PDJOqVakBPtEF+5j8xc7DkGjmgIOzCafo9syzgx5uXG
4cXW12KN8ORQK2ORzXsrRp+cTYlQTZjM9/XCQeRV0OO/8hZDfRyMzZmT44db5HzC
wb3TsrgGTqgDmjUnUskos0JiTYnhFB7lFVNGwsczFazSEC8BWYFsbEsMXCB1uP4m
vq9mljKUU0e2M1+pT0dlQve6G6mqTzXUK4NxbVu/D1w94aQMSKuF7zNfNiJlFmS3
dh/VlfWtVjaPMlHelS8hY26OKbg3zdDGH0hWT/ZkHdE8iCBcx+tMAQmA1iscs4X7
dvYiy15TITNdn7U+lqHKZ94jn44zcUUTYPP3/+6jkgp8SO4cupCAGvg/5xAEcc31
9kQVH5IOv7UpoLqzL3h1sri8TB2bCO7BTKURxyIvEPS0qaiBPgcNUOhjcIISWeuN
VIWk8/xPE4p5Apj2l/7Pp/Bix04Z6Io2mku9ikHpiz4vZXHbkWM8FEcl1uufHrBf
FKRja4u5QR6P+kmQsaPqZRhkw5W8vnlXgiQ/MnuDegJcurKRkjoVljoHI9FAi62/
20DTV27NyiYTtK8nEngdiifDWhn8umREVtmFLgJvG/Xbml4xpg7WAFY3ONIHqByO
VV1GtqfdKmEXYvPdFkL9Vu+h2jhnG3MlWHwxPjutAs7v+DzT7grCcajNMuxlwI+Y
Da6e8kzsJuABticgc207ulrFiqvG6snxDti9bvr2i1/jkvGMuqnNcOAKndne9L2o
tyijbVkMxDcEFGwjqUqk3monfAmkuOzCRtjGotCBa4Wd/eNSGmUzy1zavi+yxQN9
RpOo+xm0VdwjVOEhQz4naDWIq6TPVp7kHOby456vA7iB4EiQgqoWZiQZyZenXLRF
xEdKbhp+4yyd1vYkeWLWpmdfEtS8cPvRBL0JguRRE2akxW4cYXk70TFPCBWsA/Ny
bq/ruzasuB1Xlq0SuxpM0rnmIKe07d0fNAQw+oPdC6mhfDoTik5kkqW2ID/hLd9h
xKhH8rKX+qjQIW6z0qzMA8XKkIs8NSOjdHkV28S1A17kVaugGeUdEq+p1k6yJ1JE
qZTYWEGPpZ8adx27GlMFazDIt+EISh7ywpmZrreApEEuziIRMLZ2MArH/zQxmkA1
sM9Cc2nP/apflu9RKWUZ7PV1KBzBlirduqha2p2xE4Jo9X8oMShoWB42TSxwt9hi
StwvFzdoRZtXxFIjOekMaEU2BnySM8e6pAHqnigwbNVSs18bw7jek0rX/LVJCpRH
+pHX876VDiWCt4yLbD83ehYK26v4Vj2jx825oeVaiC5vKWNB+FYQADJvzX/2DDmG
sqWzDTG517OOpv1AjNIEIHVrALTJfZskfN3KYSnasx5W4c8TrAaZcU6/vZphLHHZ
XO+EIWfEvcWU20WC1ElQmx1I8zHmajpDykRxlSO9mcf9+fy7kUNGF7SWWC5fTiwm
Ks77PxBuqSjfn+cWVw/nhpXcHvfbQDOZg+fjbzYoli7CK2lK9duSsY+jszb+gBlF
urpbkgqmDwHZu4/b87Rj+kwbQp0OVXA0aqllFQwrizLZZVx1+Wg4dlZc/l7X6zdH
mg/UjnBYc1X7nQNKexfmxNS+gFXDrpZwMUwa+1+EsVme/i7uXFTefgM/vjJk/fJB
lZnys7h3BRVzCX2qa77VmpfKql6jODQ1KRSO+UvLm29WPYmN3FLDmpUeMUMgaFca
3NISpVR5CBsd7eQSxd1zaDqyzQoIBC7yrGVKiIWEYIo1K7DE8yTCtiPWrcAdf6U9
J/67U89+rMfmeqv3yeAbn+/oiqFKwUwKbAuN6GZLOiveZgTggIEkiTDyorMHpSr+
fxfLJznNR/07Rgj5lIcdB3jBC2CH9Noebc1HvHNWNS58xX0m+2GVqaWLhGqaYTsB
c5GU25vjPENaHQFcQlexeLOjb0MMGx0Ud3V90ylMWRLfDv51XKqoGripFji7GJXm
UNAKhx/NUWULH2ZGwIGOj4FaGZPCyZuoHh0hwk5dY6bZ/6UDOssqk+DkocMeHQW0
9HFJkVs0Eex3CRT8tx7HjvAZn7m5TQ0lfkB0eWkCygA1GNnCnMWy/ziP6ah04nWV
tR1i/dZh9R5C87NrXp7QFnmYol9ed66hHMYup1clN0cYmExMnXARvwQnIEP2AWAI
KXFxcOzC9neTDKCQexiVuWbHBG1hQHhp2U+H14dDNhzT6H50jgw8rHt8IP+vJPtT
/7ErvKfdGpl5vWh3yvHwTwg1Jb0duOiph0ahokKAmtrY4hPGv+hSuVvNu2LgwVZB
LLss1LONH/Tv+jDGgXHHaUryyrltvmzdhCJl1qbH/A6abx5EZyNpJsFZeh1QtPIU
8cGG8jFXXKuxpwRgHMVbPu4ybU719iJqUv1wC5THEbwl1qTBXJN8vUMeGaP/E/V0
5mzPMjTrBJ0SWQ2fq6EnlrRSG8PqIzn8akVRqlzIvzTflmL3H2HjotULMCzlZcbd
3Slcho+S3Z1Z5uKGsIR5G6ApLnUswWexfLQjqLBw6wrShwswyB3pqFgSpI+VfGCK
mgPCzl684KDWgW+qVjGeNxPdCmrn7zXD1Xvj+tTWurK5Td/Ule76AMuHEixe+F2R
0HwIn1r9WzaAkyHJ8hwJJBGWVEfu1tgPGnqz6SqNqCasc3iezFiXdYeVgqI8pAbw
L2ftlUjuF+BebL2DTnuANC6PWe+UjX9VZPAYtrUkOAaIvLRVV+YKPmVl70gsIygr
XJ7QdVa5detNLDA7VzJWxy32vof9ASUno3Y3zFGHy0nXSBoIgiXIUSl6KlDzX5Zh
d2LlH4aBOBjb5G+rfTyAcyPU8wM/d8E9NwJfjua79p0n0tKeMH9OVRkI3eDZxt0T
YZdGv1IAIvhe7k/Mx++6f8WcD+eX6HGnX2gwu5kiG9cxPaDhw1ObwX7wbHUaJ3/H
KgOKC3k/htlFN9MTtwHcqbcgf8AwahOyt1h3qvHTsju67/rPrix/aipC5fzWJsjo
x7Qo5VPI9goKAdjwZ8QFrZpjE11R/VJTdbj2YTB/t2c+DvHUXhA1IVver0kpMxq+
GCKYg3OQLAfBg00z6ddrhIImKAZM17UiYsDICR7aLPH/4E3RJzxl7BlwX6gv5/iz
j3ygVrhgUH6Gv3LkiSlubGqM4BKcvdwwtyUr94iD+jp0oVqoL6e1R26ZLTWgnsaL
TnBFcArmqYlxCJdWMxIUZW6HeFAcy0KQ0tmBnkAN8WtlyPnEdvbGLYHIdDU2P8/K
sM6rFKHLECUUsiGULZ801Q+QVbQOAZQRAYVr60m8ORQjDVrz82WjNTTWwAQajBEA
4iHK//C8LG83aVPePdzeS0RpUb4HBCqAcbzjHAo8NzOwE2EwcC03OSzw6QTZrAEw
w7cryHw+VzvRg6L8CKjQtsd3o/NUbAQlJfwn93R4nQdVidQz5IclsN0D+6Y1MYA+
hy0XBIhVm4TS6uKWA7aBPMwzO/cUrW/Gewia1zhnnRO45UZPBWTQVcn8HhyJDBAb
XDBlB7RkiCy0/549i9dzAgSDHt72W4MQHkUZyhiuL73D6uTaij7IdSSbv2ppF0zd
bghtThDnuk+bPyByFlquMWl08fFyd6cxq7WLdXY/+4wS8CQngF+iUrWfGqjHUy3u
BtYdC/1tjveXMKHEM5YExYG5rafn5Dtrw4nuVixL2yEzB+a8apy0iuSakG7bWMtb
D1Y9VHVZGyzJAkm1myx56AgwzUU+RnVRFOBkC4N42t9l/oKv5KcM2Vzp3Y0C2XPr
niwMKnSM0i6qeiRq9Egw28OtqgVfLmA9ro8ITfb6RN46QwtePkb2zrb6uh+TG+oE
72xrRcR2Ggy3cCatNUxhyGEUXLx/+jUJgAXjLvhjHADMHumSzAWVvyXTqrGXK3fP
WZPoflhY5mL57XSvIXskS3s5YH1BYaBm9EOribpnzdzY7XO+NB1pn0+SW9RV25U+
1r3hTb/bUHiocq0U9lf2q3YkfYJNKCEdAZiF9bWb0WGOytZgG3TKDJN+wf6YP45B
MIQBVb1z4/nWEB/IlWN1aLdtJdwbfVeuL2IMLCIwIp0d9WYtqf/BmtqaptLFM/zE
nmreQOtazW0ZBAX+DLIQAQ==
`protect END_PROTECTED
