`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sx6Ad4pszNLRYux3nQRYEBpNvms1XWQ+QaJL+Pa3QtOklIwFR/6ZpBXJ+SRrtvav
k5xIyGaFg9Qy9S2Ump3FWwwui4evjPaXAqMAUL01o6QrPXlMyUNeHSrTZABJ9oIX
wJdTQeCELvFc8MBNWCWdyYEJGANBj36pxXYyvOzggK5Gt02vF31YzDCZCB3L3A62
G/55SkoUQ1zJi9YqpxxoGXSpRN/dZUbHxjcr9vfWmVffpyyKVWHl0jc24mN+cRmw
WWPIsWitDb2e4cuJt7Cr3jtYNgJCdkcvi7qxOSB8WSQ7BvWCbsxKThDKtpMAS8m2
hJx3RqtQFNIfznoSMxTSIDQvEnrSWrU18tHczE1dnYzhAof0KzoeY0pf1bACYeGk
Bkk0eLJjmQusr3ryJWUhOfjLvhhPyaIXBmtPUjM29bPXdLsALT/PBKSA2+79dG1a
OxqGVcfHe1C3+pGhtRL+z9RXS2kGQXTqjsxfHPqkwFM=
`protect END_PROTECTED
