`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FcmcyBn4sAgRYL2OFCV7vMnKwd0KaQ+dYjiMjpHXMvOJAxrXgfDxQKLKgcUxg3TL
walBCBQ/DlJD07cQSg6nc4UB1rNiFEvDUgNCACnDQnU5kdwHg9YXgFFNYTIrAzjQ
LQxPoxeA4jB/NXi7tIX5MOYNr7mb77OjNQXTMPe8iuU3EJGRGtbG/WBa0Cfe0+MB
p92kWRLW0Zd1Gi0UWWcy5trW8PBwRncyp60faZrkREr0VX+VscuvUgfJc5vuyel8
ghNMVfoW+3sSwXgRje30pjib3FjOlhRMXp6O4mjr1KqtIKOrWRexQVg4a+XIx8hb
`protect END_PROTECTED
