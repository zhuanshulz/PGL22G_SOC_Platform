`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z831UruEzYcM3DEbOCnBXtuHPKBhcYWlDQM8OrhK7FCmNQisMZRCEbJ19xJZXKfq
WmaevMXjHFiMk3bORDBKYBuPjHMGXkGlcZBxbE/F1fZ0Z/wuHC4Dukk8PN2Jrbim
ygvNmVQh6YbKIRKw4KlB3pGs0/cq+raViFJwft2jJoyIPgm5eJ+OIoYUpXME79al
SLKj9HlaZ9aauxPTJtj56cipptTiPRJ+zO3RjGS67K9HVkRuhOn64DLwsv5FcDzg
kYnAAcbhmwNusea+5KT4oJdw6AoDrUQcqmgJ1m0T/nyxV0b3v+zgKey3GwB+Limh
Otkz9abPewxLkiK8YJA2dnIY4BH4t18vv6eluFSn8XPDfOBWRFF7jJI1fD3SfWI5
EWpDYqZc9qeuwW0PzT7s6fuh8aVS8D6G6AM7N1caOXbDlCpGlFtDUYsiQAopfSie
zety//9W4d/c2aOwqzcAviwQLFTlPaqMFF8MdjqW+wo9PsIq53ixyO/fo7gGizmi
1YbijjgWfSdEDFfPQjKyC/xppE1C9BEbCi9t25LpFv/A2ZmfdCh/29TNhNbkUVOh
cX4T7YLGask3uy/FXhP2qNyR7kZqFlQfdv3sIMa6hU4YY4MdZmQiVq9r21/2OtDy
wCoKB8vnhQoVdWaUFTB5TX+WI6i4IG1hQd0YA3kChRYlBrOitF/ZJcgqT/5gHAQH
PoHofiT7s599jMfj7g2SIO1QaQfMgueu3nzfZRl7aUdaYuvkqUUHJCH4/UeaYAbR
Ea8inBexqR2c/AS09Mrom9dqKu3GaXsDQIKWrxgFMhZa4/Y895T+5qIEqCGKaxwS
pt3YBpo/iQrMQpME0eG6liE5gpY2okshez6+7fl5PW+gAZRYYKUA+NqElGqRqAwt
FhULUUjjzRA/Gy/PMr67cKZJ7DyqeSLhB59xn52h7vH29j99Dn0rCbBgUYle0W8X
OjUwzFEhYvAOYNX0kzlwYYr7kUdJXbGkhfr0PAZUX9/c2/7MqLy2pgN2cdGPXEQQ
Pxw4/8bMdYUiMPPpDZOM9EL8Eul9jUen3yiNwfwBkzE/0RAi4RwE95U0vAycxn6h
Ncd7oIMoMc+z9h2CrJhW4XQ3+aO3SBz5D0YMwRVcEoV8LQnKhaoJ/u1IGZ0hgf7p
FKRy65ujvz8pWbLw/GsWo5DWtfG3U99ofHgtvqKn2wrnYyggLE1oJo1dbbKyztxM
PYjUyNUgj9CxT6jsLh8otBY5JFnkZoadJ0n4WNKx/fvV2TAuYfmKq1M0TuNxzq+1
DjmWk57tTHeigREfdlBLa3hISUmcc35+M0/MlxSihq3MqV6L9Up8iQcGlSGiy2wb
okW3p1CGHIcdjz+iy2Ct1Uww/0Wf98Qnv3wE7JqwnNNvigSb6Qp5nahWISsIvWtE
mAKISF+1/xi80EsHz6nRislyJqWoBQ1iD3DcbLN+HrwGautEtUJLg3o4ko5CVMC9
Ua2R1ZTqETkh0gIRaTwL5lS138AkjTm0qk0Epi1U6ppnjKxftAU8uM0n8GlbNh98
Y2QguqpTt2z41cV/0ptlmysAKYgZN6RfGvIQbufTnFoVbjcWFQsmaLyBbq+hmOM8
phFOg0HLs1OoH5jeXd7BjrvYrcmzXoR9l/NxNklPf7oslHEF6OdLptVkoI+zpe+R
NxvdL3OcX/xfJS0W012Pm6RUCQFk/tclf8oV8/VtHKMNPtijQP7e33Wfcv1N9u6Y
/U7TxeIxFiNZPYntpqZ3fXJtBNlkPxgyeQZ84Wdy1RWlKWwivG0T3kVEJbkQXPnf
YYTMc+ikboYX0u4vSuDDnAzPxHSylqhtNFx/mM+oWbyyqyv94iqBL9axRE5iEfZf
LknIbh//llPLL+/m5s8dzaPJ+Fm1Rxx7OCd+YIRXeLl/OWLDd7u1FkL/mfCb88q+
Oa1cHIpcks/nnnya0TsOcIH7tczHvLqnP4KRwc8SEZDE3iQd360cpI5Bh0yHESuw
GAcNudTGKQ0rEMQMU8d0FqVC0aIL1YZo/nDOR+4Nt6E93oEqLzjX53KKYVk5QcoF
L0pmgwp7jzXU0WURbQZmfp1EsPbZBKbcWis0HaJHoUj8woBG5rsWLM/jFPdFIWXe
bBSIAVlWlXm58SfwUFsgpVM3H6dkeX8WW62RBd5vJDvOlOwvJtgKhKxz+HDB6sI6
8RVzokuYry0DjrAljGs2+iIWq7WTG4R25U58xjhld0NwDfnFTIJ8R+J93C0LpaoK
t1hSJbqwSphTfhb9pgmdoRaJZXUYSzFnlHXXp3cQBA8Faz7Ld76tQFHxq2GIeu+a
xxwxGK7ECh3r32xaYwzECrt5vRI5DpTfOej3plRxyf+MysrpH4HwWlBxcULzTbLz
6yIJ+QCYk820fV2+F/444GW3GYzjMZXTmcH8jYJMqAM7Vj1NkY2PauNyo5A6INd9
QrTQdrmwU1XcYCm3QyUl6ar6UF+D15dhi4/qGrxfBLlm6fFpdWYQYEQq6I+MgLYH
UM9p1t6H3oWaDkV6aEDVDo5OYMWVuuXaM/27jZ6ZPlFNHAehdCrTq3kWJfcwg3EN
y9WI/SLwddvKGpqXdINSeJiUJk5onquXIb+v9i1A0PLylLHdkPgyVrXahSwLIKkM
TZbsfYbk4R8YENSdApz0OeWiLI7PS5ibc6xd0CjYk86LKeY1e/dgEJ5DGvaRpXjd
7sHBQ88FrqpE2qYLs6PiD98WIdMk9rBL3XlRV1lio59yE0NcqWO9cxcz0QHhAx3P
4MVuVNDjheFawSHLVW/4ixjdkXbF9Kwb90Dt9AEDRUW1jlRYS+tnU9RO+jlo9ibP
pc9e/HECkLNy5WD5M9zrE8TYccLc+AsAV+XyT1eRX5O0vM2EYz17gyWRAdwYWsLU
ComJyoar4H72IHJ2luG/R+f6HPhdRrdMlVSmAfUXIBCjwDghR4P+FbC6ftFhX8Fl
5NxHqWTp2VtCh8vpJVPEtxunxRRWMCGc0ZFmj4acNrEVxRttO8x0O5NjynWPjSfX
Kg3Zw9tbX8dPLsXPuBYwgcHU9TUR5Bl5W+oYEW9DdzcZXTIEEkxZvOTTnRbSjvv8
KLVnbo/2dNniAue0BV8pbXqYh/serv2fusc/YkDEHAcFTiGg3OVahEY3Dl04+Wyl
jajkqiEpIspFTymfzRO4qdxaOhstiNwme5Gm8ZdHQi38z90HIN7IlH+Wfedq0RlJ
5xdUlgS4g//zHv8xAXlWnal2E/gHHFeHcYSLG3xMoUZwtQsqM9RpHKH4ObU74KT+
6Of3VydAESVjDnOFRWnA4Tzo7XlnvWmSvoKIX6461jSJUSz0pF+fLSVMs/l27cWM
kUtXoL/BAhKsySK2iz0BmcE/s/ztcPXm2NOOqeGcnyLpeDdfBG1zywknF9edDkyt
So89fU/0wKH/mCx2RPaiaOYwW7Gtwy1XcTwn8Z+0WYssHK9QyH0B6RzsRikg2EUq
oFch2dZ3h1cXfsrPVJ63UYCn1aRddx/bTB49Y13YYpayeWGI2wVOBQxivRSKg5iQ
tmGH1/1qtnXWWUWKvEEAuRhTQfO+GfGa0LXXvKXZyYjIwhh5jFrXkL/ZntI1RhSs
CcTDwnrPAu1RNFz4XcdNwUAgiM/Ia2EVXAiOcpqUkz6qYvKI15oSdCpFrsPTCA7y
RMA+TyH+u4eC+YptZwTlBItEbPyftGuIZDf2KBF+O+wLHKt3rhesBngF/+0CtAp0
urAZ0GsQ1Zc58YRCo/7UsYEi9MDminbWPtoNFWuJEhJq+dE1ZeM9wWuolDu7rRsO
y21eVaIn9MwUgAhozDToCynJs6n//1HMTAxhcNUWwEZF1uTiRmtpyOi5mGxN5k6S
GkeMGX1ZCZA805a5TeWED+/80UyQfxTTBns8SLDp9iPZjFd/MKSZdPJUFLCC2XnS
cOZpXEQiQuaYd188wQ2AoYL1YM1EuuN4s0vDmzBeiijQ2GdBHX7YT5kkeCvP3hks
PNQ6CvM8KxrKso+AZKcCNO/RBYUEAb7fEOmMFWePZ9YRCLmDKfcksfWR6hpYOxiT
jChuBjQStXFTKiVTALInfMzFfphBsQPjUMepH1w+uVBwXlGH/1K7N9qFfrV9NQtX
`protect END_PROTECTED
