`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z6Het/ejoRqhAAYdxmpvUdUzgmq6hFrD6rj2Ce7td0YiJx2nYB8VFlDGxkWZrj24
4ZjhJmHl9bs7eNRdQb7XO6j1Bdiv6urYaji8N+ReshP3al7nObgkiItE8HK+my7R
jChzzPDVfu3xh/P8z5dLWELBA4noUPXHLqx3GH+6Fb+Nd3vDOIuRJtFDgnM49TZh
/JHtKfvCuF1DH4C8awBNVNNanlbi/NtyAVUp0QjsjVfNDlUmElyfIRrTWwTooHB6
O5V5iKJLxrjQWeSOq81kLH7m8BvpiAuyMVvCxnTSmSEeIbWgkmu/TUckwbzm2Qkb
/3whQ7vucLFGt0UQeXMwX7wDS35Ukq4xkbgWEzsfIKduUwhMnS7rQzuKn40jVK/9
MMHtZauoBbtH6Jolan/0md5zRUoWVqTiA0CIEX4GFTSJ5PWc1No3WUZj9pXhOGRU
I0DWR/OVqwVhQncZM+UGSnXGJsLT0B7RyuCZ5EKKolFCbJaYOCJcgheRZpIa1bnJ
E800D7hXhcu2aV0dWGAi1gny0t+RdfCMsoY0MK0MxiIbkunY9otEo1dWL8Kn8QL+
C5LWHblbsLAjlHw63UDokVYapcIBuvBD803hI5XZcszi2eaem6z79gV/S/oYiUdp
WadoWk8gqJJeAasSxdssXemSprZgNswDIrrJCfooyjNxD8FOPn4laY/koy+XdsSd
w6RwVOTJWFiX2R2MWEzEWZcFANDX/HcYsXCvAk8edxkdFkzAeDVj5Zs+SGyZUjH5
A4z2VFfYy0G71vb8eyoTEb0mzwSB8EOIxxvk1fJCLNqZ/hCYgGutgk8I8njx3OUf
IgHEAUqbts4ETUh4RkUEByZQWdFkXbg7SaOdhWSV6jHrZ+L8g5DS7aFG/Kp0ZbbR
eNCN0xUrbxIVf6cualUpU3PqcZMgQ/eae/W4XEiV27LWqLvJVx3xVOC4szY8hKVS
tJo44dleZCsFH9GWDGBq5NjcijdprNW0kN8EbFmNQ0rD53aaRrVwMfnW1T/MzVzQ
2ioFvbdtaY68Yt4Wz/RxFBbOnPMQJP03iBiCQ2Czh/EzbvFr4cLgJt9tYKxwjqcP
qTGGnXX+RnVjVv1jRzlsn6bFpZ7C3o7gFK69xce3jUr83kxVm7iUUYYqC9LfPXeW
nRreDRkZjaWRnw2r6oWRewGMgADVpwPidw/6awz0rMXozQPvvSwtweLZHITpgodk
r/eZLGVxLMSZmlJ3AE9C38C0xSlBWr+D0YmDDbgDzrLI085/xk6sKMN/4ErtJ9nF
F5hcRTULs8KMnBYVq8BQbONx22wEgy3GvXRchjoam9omTu9ctwrdsRd3Dq8alUkc
oAEzNNw3kkD4ShnHM7LK4K9kv/VfZpCTn3YmVTe/hjSlh9dl1/tgDuI6xaJq/nBD
i4+3uc2ffiFA7Ve8zEZguOXw7mjWY5TnyFq0b6/t4IAyP6EGrB2bSwWKG7z289L3
QlyCNnRd24IvdVbqlBPLEMl/SlskmAiq+4m1N8Q4sPR7ikwFnSbFJ0CmYWDmA4HR
WVKQ0nL2XyZlVkLUYu/Gsv2DqXBbI6JfZt2D8aoPJxNbn5/3DXJ60bNnMrlb9CuP
wU9Tho/Ew1t1+ifecWlvLG+Y/9xQFbtUm8wmY5aUuEKdUlaWQLguWv+PjfrlqpPf
ZI2M+GCDHNxC0eUhbKHdh3F7L76YUH99kerAieFklAe4EEEmpxu6t4ChAwXxHSxz
WGmggOzKD8kDyBNtn2nmxIaoHggFzziroK387aH5KRBy1k4ctQpyqurpknNTNnX8
93zeQoJmxqkrma8Iqwc7uNHmZdFkpzOBbZKu1cXnTRpL4LOU0lqM18sOLFAGvGvI
FvKL55s7WcUVfp5c3qhnJpKelzmhAcvyJ9dLmjvP5QlUdzGRhR5nSM2GXSUIzkxJ
bZQ4ZITHT3ozfpHp/d/6ceJjqd1C9DvM7lL3FV+EwMtxPkxgrTf8dlT3FFjqgxt8
sjXKyG66KPPHnI7k6hZAGNfsLIN84Oj6o9WbCw5ccrZVT7XweuJtwIkrVGdUtFSQ
`protect END_PROTECTED
