`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a0yRkb3o/yNEAPjrvkZ3jMUFRSY8sVFUbV1a5IhTPmw2lnyOUdTTyea8+0418m+7
o49y97VAl4fVw2PRLjl9Zig6ZM/fV+AWQs7vRD8nmxc/jK0vJv906u/RIaiEXJZ0
LJhAS0K2neEJuL1XUzxhKOqcYLz7/J4gnWpwa5PZ7y7Qh99YikrDlJwcTjQUb1Ct
QB5xZAS5A3k8TZ4zUEFMCSI5vnzG0jQpEKg1tOJ7Zhi6jTMpksppPJunfsgWYGCm
y9GFnrewUwYPoRELa0sgaOzp2/LVnlxrJXSCkOqTkJ6YQAsdn8iaZoOKiV54cuJk
z29Wofw91YSr2i3ybvhc4uhJAjnVu7xP8JmwBADCZcLSX/XAV5y6KitQBTbjWZAi
jrQjYEqey64B8B0fVG8KFTbug5DKowai4tijnT0OFHJQ/zUvBerodlN2n3tcySIk
9D76S2z5BsiqtWBtE5n3qk8vi0OqPOWWqQYULRMv4QJ3JiWl0xkAXNjwTmIxKgqy
DSe6Szx97MaqXSJ9dJnUV+aiTIlrb1qI90tjErzTLjJPeHIV8PFXtHsUod3jMqtD
xTGJRx4xdQHU7u4SanDm9Z9CxnIb28SOieGhblS6QHlu+amqgSCbQwurqcP7Znai
w+Seuv5WEWHuZvYET6O4Bz66aCXtiWO3ZjwjydRKZIVCD9uhk0OQPuz4hxQUj9E3
1gc5CmZ+Ak872g3gHfgibMnmLV4Vm0+NqAwfO9JNzD9SS3+iJXgOuaM87jCi5LAz
`protect END_PROTECTED
