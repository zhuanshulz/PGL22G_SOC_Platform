`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u6hfWx/M5zqk5mWkakHeWE8MX4aFBRZfHcU3BvJp1NPjaXqvIKiKWR/udJdcDDxo
ABU+OtACYnJz7P+AGpPoi74F9a2AJxvrjJ564aiXfrocXvv2Sj1ELiC97hd40CG3
BRKRJQIUNwUCrNoAYeKZvVYJEuenrCvY6o5VsBpJoxlz7iUpVbw6z1wgt/y4uXZZ
TN4RB0yXfQ83zf34UYbZr6TEeVWCnS6jWXGQyFWlkWzJOlUUT2efes2eomXHBX2A
lyYNihF+L+BUjPNjPUOHeSFOzgF+UpoyeiwarBnOpguATN4Mhdd8ZB2223jV19gm
4nUCqTZXHfVTwPmHAgQlcfbsJI1LzW7QJbkla7bhtgIsrDclOcBGas4+w4JdUdSr
51VLWKV4eo2ghKRKUDysvoASrYGgwxBCx046NXIpxRDjB+TFaVy9mCJmKwpPZ/45
EcEQC1jaifO5E9TFSjKMictf0i/XH4VG0XnWBWNZDbwtdr6ZhnW1hLCDPyvOhDzz
KINsiVD4vH4nwf7u0U7vlY8QMyfgY4VR2ZuHX+84RNktrP4ettRIn2IF6J4/aRaE
iUOXmT30S3In1VUQsi7IG45CUEESCPbp3f0vspZSu6Ryk0dqXJ7TTIedZHsucBYr
wmhOEwhxtaYudl+ybXHsV0gIf3Qg9GX7psVJ16DjrMQLUUqcFHfcX2R9Q3cCdg8A
eeX6JAgk3PPBNJgMwQ/aEXfb/z32RARdN9XSWdOit+7rxbNnHdBOy22W0BoS232P
rB34Lv8j+0vkGAnDmJEZOEDU5ie/ybXq6X5ix9qg0TyQ+i78yZ0PFj7agjAeZbZt
zklTQxUrG8Kr6G1QG+TiMTlbiofvsegfdg4Jlg+qvL/kXHud5r4HaVE3ktV8Gyr+
KREkIWrQifb5wa8OYvELlI5FO8AktzkjJqGelJR9NGzm7ybTx4r3NNSQHjNUsaIv
2yZYuyTqiLx9Yimit7ux+iPppKLDgc1z2q/4Q01m9Bh8UbKi0MZAVcMaFDdPftoG
zrDBLVk0LcjGIdqgzJNInynu0O+u5B23FdITMalY5u22ZYm5CVEPu7jkibYlrgxW
sMLKlQoQfpCRk63iL7xA/PzcreWwrHC0xXGoWqQv13VEu3kerwZpI5so+TTdFZl4
cyZU9b0ud30KdKHOgULjzDxYRTlpdpaursswihhDkDpnZeE7+57MVBumba0ZNqNW
ZRNFDCccLmaFSWiISjZ+NQUeFMPkFOXj7CsNrxa0jzdq8Q/hhftykFUkNpNrAt8e
qY4BUgGIYHjGh+vsiWaql9oakSz6FIw2+ZVjmLkajNb6idExNOd6o7CJGF/31ceQ
jlLCtOFay434eSuR2HzM3m311/Xi4p67mNd7DjxPDOkI3mwh3CG6SbH5GRkZVvph
fCRng70o2SEMNxrl6lhEIjMxOz65lgOjGQzTqEnHk4AEK/zXBI1+wVRlK2RIrObB
otPf5D83WgqQil6UBqcisALNjqXHUZMTNtofcfCiTJQ4zrQWlaxIclh5UExSzFoO
MMNkJcEkAsar/vLlpS4jpOWZZGfonJWtNxNZ8+nRQAdBg2umSlwuxGzUto6ebvoA
O1M64XP4yyDn69Tk4ncckPHFw+jE3D2D4k5E92/qY8c/4+AMxsSbXoplkPInQio0
rgwCTMdAgYgMJE4aI0/MtlJsWUbVZAzPjyX4rMriMPw5AE0H8nrUSdP8Esj7cm6v
iiYzqPtIxj1we5LU/3kaxzGDJTjvPx/bZfG/ymPjyYSeEhM3I2D2DrIYP9Rku2uI
iIWaojGliQ/MFP89I7lK4Ya87qBW/abab6lQbSZn21X1YDywb+ijjC1Lbc+aHdXM
URE3ng+EMp4v7SDICzkANFiwqAdBiY5mQ0FobI74YCAizFfYC+AqFOAtcDgORWuq
RB3QDjoIScSxflvGRfutDNt7e8veirnvH+MqQWl6r7hJlrbDJd60HQlxdVdMsAYN
QKNosrlCho/UqdcNILwA1YYNYYn2wh5r83fmJr7Q5u3NyxPpgsY2CJO2X0+5ltvp
SwfSDfS4ZJUpzshK9eJFpMrEPpROk79tnPhEByBf6VjR/TopnOLFcF6YeXAXe7JS
J9QUYgjiY0sdC4RKZ1MEcmnBLkypcDDOJh1lIYtU/zCdruK5zH+xnWmEERU//fXP
euItyycmIe3ntWusoB50U8YpG5YIU9hKnzMe0KHrjO1jSma/asGzNRTMtqsIt2Pq
eH3D2RqIQhWZCqep6hrC5PJBqPXOhFYY6KhXJYHoLJxW5YTIWLyhfoNIb2g88hoS
TKUCMKujg43pPa5R+VVvrQ10NmHbISU3dhiViNCszrchYajM+6IWNRehVPFQbL1l
`protect END_PROTECTED
