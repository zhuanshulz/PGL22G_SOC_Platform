`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0KTCZEpx/KafPHJPz6lIU/Or4Ubv1kCmnCk+qZjxmfPoZfRLL7ou06xJShXFosiy
Xw63Zx4Qqxi12kwrbI4l8RaRnefU0SQPeJjdMZvEe/ASxivzBBwup137IuctJabV
RQC5nJfXELtqyVJETUm3+kVorlLj0WXIqJW7eUiV5UBoIjdg0DviogUPeSLiANm4
owgTXalgXvyGjldHf9Y4/VEsSyCpJ93tEBhNf0Tawnw0gERMQAuwhm0wbTaU8nI1
GUZ+hMCrcNoIe7EkD0RyBAeiBBgCdNh9wh2PWokJ6pKhlAsLjozRZHWk4lb48Ixg
hFlm8CUeQtgfDIG+IZngGmqxwGbAPHhP4gdoz1Mf4tW5SZI/IgOktvNEYjcZXIqk
uF/L5wh09JKjWDJHOuJ7DQ2r6BU/YeqPvB8V2B+YGwTeaNHHsUEYtzwo3/VvJmCG
Ts9WkMSwhp53ZML920NCwALVA5QfzVSal6PnU4oxgFe/nfvWK1fzCr++czLG5wut
B3zEGiirlNhSd/gGAzOYt/GBH+hv2J75xobAMfMKizBwfSDaFr2NiLrH8889N7Uk
2HU6QdSnGFFccmy8KMd4KY0szmQ/5usI49A+Kcf3GIFm3NYcW9wGy9g38mg/Acv9
uCESiSOOoqWkvs0jGWGO2DXgGP6yrZmYk7xGZUis2j1YL88x4H9UqDP6Iq8Y1/6K
9UVUrYXrInmCB4eckctf3EYwfonYwWLOWjAjtDBEVvltA830YNd4JbapB4AdbDwx
EwPwT48fem6PIgOtZVELf5mtvusFBUcyhLnL5v7fvgzoECBKyq8OHFh6s8Ob/Pvb
mIVUDV/FgjZrr0yaXoUQN0ntj35sBrCQLKm7044YEaRoB51+wbr/BxqmE2VGBosV
17z9gBJDLKFtReWzYW5p7KZRK9TiDAAoEn50vqRJ4iaAXpeleUxyWJx6WvbzXebk
H3gel0qCGVNN6DQQKzFghil+mKfoV0S18n3G5TxpRnbiP7wMQtTouZ9IiMSM2qwV
TBSztxs/uWaU+/at/zhjPAoN4wq9qt2yTtRkpIF3saYEi8t1uC9nfcOX1sImwCor
gsp4lla8tO1SO4+KtkVqiGItVewCSUfJo8phsE8DfRuSEa2jQt6fqxycdtLwlnfh
GLGKbYrKrXx2BUhBonoC4w==
`protect END_PROTECTED
