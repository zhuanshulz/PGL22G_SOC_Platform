`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6az0p9nMKwN5aDtjjgdbybXZ5CUm5TDbzSSW8YuYXR3MIIuXenCJbuWa9zjNxLjR
oAWnsFj9blolLb3WPl450Azs3w6sQ3AmGy/KCWF+OzZcaODA88sF2aHGiRGM8v01
xIi23i7hQA+OF0HHnPPvVZzd8y+BNjkbjpxN6rngZEOUv5BMUwHu7A3ogPIaht2f
C23LNexvIHliq6kpBAT/BSQfqbVsGi4/xJJD3+cGA49xgP7AJpKLzgEDeGaKyrNY
CmtFbCydI+sWPZZMutnTANJz6gQMaJrf89+BnVBVfFLabHfSlZP51a3hVxN88Qtt
dbHTX2DBUAPqu0FxiIrcGa/klpX8TrBcjt3tunYZSVUloN+z32WDXW+MVR/Qv52a
N/H3xuTPjp3TE+HIk54B8+vu+l3we19+3CXvpYhJi3XoZtER0um43+478LUOr0sC
Hl+i1JFsvTAbrz0ugr42/pbNQLqHy07zBnU8tOmN7gh1ANkZksWZ53xvTdeSqr4j
7k32vystIp/ylTFbI26lRm8UzMJcFS4RlahrV07PGbdF0jP4KC+eNMlf5Jqzhodo
+vpkMSpXgBNvUu8ombEd+w==
`protect END_PROTECTED
