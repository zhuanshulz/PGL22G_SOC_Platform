`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DJ1q1D3oS3WxGi/SqodGaVy/4/F/OfB8bE3W5Cw8Csy6FLrxLE3ownAHt+yyqlai
yEWq5MIA36kwDQlRbEMCMAYvyTLX+i8mk8ZKgUZXu6yJc6c+Wz8QvquxutdfKrKZ
Pm4mZRzWo7XA9omPSmAp+sZESoSlMgCrBgZHJ+ZKBkE5tB8wmfMnjsrEqluLBt95
QTecZZRMmCyLiHqgugsWT44tb3LObLKxjfpg5YubsruZ7pBi5mKaenyBZWeKFt63
ymZF5deNzmLFRhUvFZncGL3zXXs796JQPrMTrZbppIxOFhaQ2QvHwcZQhUr8HOlt
fRnJMQwkUXdyQhMhZIj5dxRKLDjLTz5DdtQL0/ypFdkkIui1C+0LfcAgBbuHqCNA
/f9CDslS6zw2jmvcLT+VQmMJ4cbkYuR29tJrUSLkVAnobOxOCVQX5zOi9XxABgvR
9qhG7obxsDVO+N9lFj75VFkBfBU7v4sYC57ToM9K31cio239bKe3iT5spiAMd9bd
f5hKbfZsC6gWIZSgUuB4S49AxzyqUf3dJ75ZVRmryOPgEaPWthGOyFOQDJskkrxm
LcLdcl0oRLnCef53/+qrmllFD/nrRLHbXxcK5nMj8PwsT4td3yqbyg5obvZLNSnR
h3hmiFgWVqfQXGnPRt3EJsVlPPfXo67yr7ofLARUqR4EMRRK9ztxkJChVbCPtoRj
24weZjyLaRXZQpDbeV+UGjCJSr3IJGBtJ/HRy/AAjAHEmST/gAPw6Sj3v5jxkug0
a/5NPl5Ixgj7EgendUcUsMA5cNKn8RWM/3QD7GHyhoIl1p/G1ouGXHC6BGpkGY3K
`protect END_PROTECTED
