`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5W0N+16FPMxQY4tDfEqDRzzbbUN+S1eYPbnGHDcdBOG1qZMpLy6GjmP85iEW+zj3
VMv3gpglWrx/RYSZBXIHGH29WNQT2Sogr0EmFVHOspPYxrsKWobNcpzx7q8/ZmY+
MIVS8ScdgBz0R1X6sPIaW4hW0GA/NQhk112hb2t77sIlpipN5smOo/5KIAzykTnx
VWHjNSRKAvKYsbJ3JvkLKVRCxD5Rlcn/N867HKyNqkpqCxOd50bo3zbAjXt9KG8f
yNMMBt19hMoHkN/STA3wAIoryv5LxEQtinrKNU68evtfzPgxsySkje0gAYTYT3K0
PiMAXnWcN1L1x/EhW9FhaFp1nwZs/j2xPcCEEF0dF3oQldv8pQWhcHLPL4IxUnCT
rz/ywILv774x8tyk0iuyw4aiac5fEr7pHLGYSHCytQonRW4UbykJ9LVCwuF2x8sy
jHaA88BPECgm7rcmOfWZLFWfoFN9WGKxJ0lDa/BbvYLkEBsiwLaCuKHXcdr+qO1q
JQnxc/1GppwGY5Yod6VTKIM8C8gg7Rt7j+qTH6prhEmEpbn8Ffopy/rAWsPWI3uE
NkLzxl0eViK1HHXIA2hIqh1EwjAdbTn/51NR95dB+6r3uiSJ2AhToNGVa0+phvqw
mAycwTqbP3C66ySrdq0rTle0VGZzmZslG9DBs/Kx7o+yxUCwl3Jg/KBNSR4v9qLr
9UcRtMLwUCk50zmGE2lBJ2t0Bqoet+/OZ1vEvz66sjWUXLKj86b0HFpPFBlBn46+
WhMK9/Y+blYK29wkThHqa7S8zhJrahHlLvnQgmW77mHSo2mlqXzk1UYyjImzYNzC
aPWzUsu648MrNQ5bi/g5BVeIsYE1e3Kd7fidBOSpP2P1j/M+seEZeL8YrtNLSg2/
QTInjmmLnx71Mh9A5dacujbbSIoOfICWov8WPrw2weaKKEpEDmnNaCx7+lPHqB+e
rV5JnUSdKFNj1r5Qlg2RagwEEfP1S92/pZNWKlW+LiBQQ+m+Mkc3y00NiyCUFsH2
DjhCtOE3tiMLpE0hPXhXD2VnaOUnToEmJbzPP1vuHDKdi4IeBkiLvpidqPd7oYOG
vu7aw9GXOvCY5Ahz+T8heOujWGxn2XoeSn9Tto/mfBMWqTYN7CAQuSGmJVojcXf5
KxIsBeB0i7fri6F62BMHgofAJT4img92FuI8LF2aDIxiZJiT8C8fzxN4qlze3+BM
SPOrt7KwgLSS1nbn3W7s0wsOWCFDEhRWiB2jIRbG6FxdUFXEqCvuZrzsABNS5Tca
Gp/V2K3oYpglZlAILdVZlRoGxZIeTRaaI9kNQ2znLfVCuWYikWBtk+jwPMia3sen
e/v1WNAxu6khx+yULSwbWAHV/JAQhNk38F5anOyglxO5q9Dz3zzomLKkbSCrKK24
bfYmpSqrgPcfNL+akqL2T///q51CNSWcrrFC7tmoh9KxJmwqENSP3RGfMmGl5wYs
VYV4ZckFTR7/Q+yZv/EGVbc/Tt8P86C1pakLmZpiLo4JC1GHJMqXu5INz4cmnGfn
H+fnyE0uiYFu15qy2BNJezkMYStpss/4zGZ3ewcK+qVHKlXuQEOLyrZaE5uojBcf
ZjiFy24DBLptQOj4xZBSnyhmnJaAB06vdrb07TaKsO8nUt3I2Ukzg5NYvfLfS+Ub
ocBOkTce6NyYiWV70QH4J8wmsFzmh/H3Min6qNKyioFCdITpRs8Jn9+t69VJIfd1
cY1Nv6ieHjDU15qwhFmGzeOc18jUrLSd/jnCTZDqmzuThCRM259WdCsvRZfFiKiP
yiKGZwVHTdYqwdIbYmiKFaIH6qBAvDSQ8VZKVy6Mmz4IqtJU1C+XRWK7/X8NupVb
JquQ0a1fX4p0csRBuVBruIPZBk5YxM8YKrFm/+3v64/3EQz9cD1iXB+aUGQcLOHn
ch9YEJ9k+kX/lsAfzfQzShJyUWk5+RgVBlglXGjkvbyyEelU3tssXJBmaTLi1Azg
Zu7btmdjxLA8InMkwsB228HwpYDCC/KyZh6my0f+K4q4lLJmEYy9s2Hfq2ig4tf8
hxibmilqkFiG9AwmxSFidzMumDawkL8iTg6oDZw6ZYHQz4rjsdmQi8k3PM69kpIP
fdnSyIeHqKkd73oErQVc0WPVzTSgnDR8RYf+EJqb5Q0klUxZkw7YKnMP2WNJwNbt
PoJGtEE5BShnawDi1PmIM0vR8EhJqBIDktIUP96Ekt15Dk5zpCyXgOOSZzN3ZdI6
QMolDo7MsFTzSfXIpMsUA97NQZvF3SoNjZzf+oGSJgbXyjig5i3YJklzF4P7WQ/3
djXo+0wbILX7f4C9YsS2J8N37PT1D2a6hjpM6B1WdsyQBRTfenoraQKk0CUp9K5g
PsvGqYTVVU31+EloLjwduE/w1B3tS98Y01OLh5/HB58jD81hleB9RVQMVzJ1HXJG
XM7VoxHz/H0ysPjdFszlPMPzIX4Lf9NcFPFvgR5t5CTGOX4B8SgiSjRI/Ympojid
UZIbsl28VdCQDLVYZ295fVfiw8T5zHUkKl4a4BWxRQSjm3X0TlUcONazugoOd6eC
O9qxPvNJQwNRGEdXpRJYEk+9o4TNkEY7U3XCTFaWCyP5wGzidbvRlRYyasYJssxK
CPOTUamA0VZRKv8+qwgt8awCoxhocZoGfFhMC3VWHzYlmlwl7uSRku43j/VqJLdv
5p625xp9IrNIf8DDMI3oh7Y17fr7h4jOJcaNW9BMyFTajSg6WLzS5EQCsPBR4Et8
dl8pvWhvqT97mEtdHOOD7b6loxwl7ViN32Njd/zaMHH3EDk2l74Khy8NoT3uVK8U
lF3im+ydnxd4QIQ1hQhSrfy7BLe0uPl3ZcKA/eFYroZd/OodfCPchX5eEqSFCgiC
lyuF8JQnH+tbxt7RSHEI9XKY+nZ4HfdNnFcNoT7EWCmukwe/FWmfE89liadt7zf+
YDTmuQgT0MDQ+RICDAyPjcCTfdS0fR6Oe66rnp8vJ4JQ2j2UNaCOpPSpvdSMp7NH
vmASpyH56WWpFjPUlRFJmjlsomboWK1rPp8H/Iwp7izrXPo2Xdx9HDjcsITIeaqz
CdDvCLUBPpo5izswP1S0HL7z1OGJuAk1ucIgLyJJvnRpvVw3cMhHowzimNIo7l3y
AIOi8ILSMP6ELVERUslUcoG9hmuxLyT77jLwF8ocQWEwoUvTOxjxoAKt0RxhHD61
/6lyUImoPm05Vg/A5vD/QGbhA4xT1rYGAMDfUsil6a8ThfPNVYr3255Au7o0EFR5
l+7U/i5P1gozNBjMoE6LkbQQMW1uIgCig1MzmMBhHWpsoGKURRAGvsL585N0nbDF
XnUAjodb5b0FrWlMuf7G6nE0FtPUGUEsp3QMqpCNZoF9UMxpqnMFqWfdoozggsUO
CJ1s1WtJFIg3J80lYJcgxbPSHC1Dvkej1GPIg/+IQA2JNrhymYC0KO/+C/jPWVVp
+GZ9atN64p1PP27Ck72p/oSplwLnC3TfX3cKC0pPOBn0upWNnYMQL55S0JFnSdGa
kuuIXA9KqrX/5cCkMm8U7HNPdOIuH1ZXeb4mRNc1aj1Bjc9DVO4UMoBpx0ddYuRi
CpP6H7bYyiwY2KwljAXShu5uxB8SPBg73OKDsc4kZYVFkFWYbFB4Hcj/Ar/1bnNw
nqd4WcJzoUibYCPzxo8VVwlvbyHdHzr7bhYXPR5C8TC9YEPmH9tWM+8LBUt9TdRQ
CDPYeNro996+sq9VefsvZ7YBztsBuebBMf8iG39tD2tbB8cDsyguYQik059GgGtT
O54jB8A3AXCVu6/052w6LOJJCkLcpMX0wLbN1TkCzZr4oW4ot0ls5GCNb/TvTprJ
MMJCDFR+H1BBYSrMsREl6g2XzgAiuSyXDuZBuSzScsbktlrKNJ94naKeL4AdTf/u
ciILXo0zI0nnUjYQE4HHQrKXgRMD7DntlZU6OE5BNpiBPMdTQc9XBEY3bpR/+PKq
sMDl3mXNEyPdKLx3WCnoUo6+5NvaJmr7Geq5IKUwf2HIUlvN287hFbkFRmZItwxv
5jJyGdFYc0jvkE8PUWYwFQvpXiYlrb9TN/CRR3/yC/PUD200BJ9sAIp0JGa7qngV
NzVv1Lb7MnP1OSm92vcgCkZBwPZ09pOdhIyxsex+fUh5rpiXf4R8PDboe/aT877O
qV4oguzJSf3aiXcki24H5q6RBA014hCIeyTBncXOz3uoQcJINzHRSgRBrcmPplpK
S1hPq3Qz9d5vm/ZG/ebitg==
`protect END_PROTECTED
