`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IV0QND/Ndm9wRjODyX8vuzmPi2mquiBEZeyf5VqXbstvyF7T8OQneUhaijAfkiQD
KpS4yV33LQ3oEA6dRlQs5JIw1h2ha5QPuwlWf39OcUbjxU3hS51D3YgPOY9ZfjiU
eQMHIhIyV4uZ8Ct9E6NSLIOvo1/O/BqNthGocv8RZN3auGXdvBihj9GkZGU5R+PG
tl7cJE5eWzFt9yQLqO/Apj5wlc+LsgfOOfLAj2CmfkhmEoSZi1yGMTHqix3GuZ6v
/7ot4NDsmbPppPGs7AQrvsWmhhgsryzUSmVpTjLXlmrqVY4WN2lAWZGbGoMCh2eT
mocfMKXJAKUyRUiZRY3TNHTg3YbzwppdSghEIHRf83BmCvYSu/8H5B42aHrMws6l
PJHZEMk90QxCmtTNEKO0FmRHpC8LC90ZI28ZyW9DmIpqV5J2SoHMEJLJGGe5Bkn8
`protect END_PROTECTED
