`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K2FuJikI2vAIQhoFZbg9qDp9zUl/h/yt5UDsl38JKh1SK91wJIWDX4Tr+rrVcCQj
oAZCUdy7jmjAwNFvSSJ8tlGjhxrSHlIeGHwuagSswZXRSRxu4DTGV/6zwYMSBdhp
pPllWK5CGzNUFk47LURdtRsaxkPrisgtfAeheFkdVHObuPtWS5GpObMRmjZizeYa
NYCJwHddaNMmlOzlBoW3TDvgrD2HaLUU1XlF1fezpY622c8VgIleWqhLp+soWfhc
AOTQ1g7grVZtfwx5VrbYgZ3wiImHfjsCi2gVksKiSSYj4Z/uWlHi0ajfScvHDlcI
cbE4Vd2j0BwhTZpKzPUHToXYw66STQrMKB7kf26A2tk+wkmYXv0eXVs1vE0fT5/x
bCNr6jSno8W6iiZcZzm0+Tc24ZODSbo5E0nKUdefI3d2geuCvE6tV3GWjM0RtfP9
LfH3AUVw59XVwi8xxrOHZVjH4DVMPcn1OdAy3tTxxhv8dekWlCbXbbEsVFLuJKeQ
e1Ykbj3ipRj8AgdKd50iwha0oKKooykyQFGsoI91S8WjUozdr1cucEWYOGwpeAko
UFhHtpnt+B7i0x8PKi2hwQsQ2CGY30gkjEAFYuZjKf743MjvCLw/qLoqlaRUL8BB
+NR8hk4gJV1VvX+nyX9PtHtiYR0eAtAtPxvVuOm5wL29UQCj2eDJUEy2T6XFlqp3
AqO3tsK+U8H2KBTP7YkAMk6HeAa7T8Ei+Dheks1CS1SIGWhvdNWNJHNGjOdhtJ8L
bUG/l5P0k1huxCv/xCno0c15upjZ5T2lZ+EX/GMyFMflsQFHOqxmtG9N+nFWUROX
MaoVO20VSoEiZF+nrNz7rZVjtH+IA0ueHFyGhzUswT67eWAUIzJCLPIkjoxEfXBC
j60McHEInlGydQuftg+g9mN8wV+vVR3dD/jtvo3AQx5/feAiBfox668RL2pMEkqb
AwAZZARiocuWQcW8sy/3Ghjtw7db27tsbrQ+Fd/zkceDRpVsBb8XAvu9eNohWWkj
BiVWmQVb32bWwv8nXrL76g7AL7/1rqqsr+sUzKdAnMk7O4KUgsSYiV2M4tE+3XiA
EZVuxlLwC8Kr0jZsHM7m885R+m8eFY9LRGBM4sr/gZ87L0RxQyo0ptZT+SDEtVME
aLM+dHAUI/8UYJn848u2ziQzU907BLJ/66R4OPHkKdYBeodfMm/OLw8Pk8VwuQfV
4EUw+LDKE6oOPWByCPsFM9ANqaBIsJE8afnp++TQS0zIiJFg0chDPf25Ef8EEBR0
0XxzatrXuYSEwY/pyZvYaJe4DxeXu3nvj2eEzqlkNycorWYY17X4KjUj44PE5iXJ
sUrXyJHOdil0veNwNVelPuMzuecv+2nI56YwDtljoENuDqpaZ74IaGFhq036J5a3
J8du9NVNYVRrvF27XjyaxdYLRD4MBsf0F+PcTDJWso2kPYyBLatf4iW0EONerr2m
lyS2ZUuCPGHnjvQmjDX18cmttQtv/FQ88zJH4bXP7JXxfJ7oIGqY8+ACIiXKj4be
HE9TpIGorfIQvmjU4uUFkwHPNPnMDs3uszAnDh1jIYLhLDkEubgfD690vZOqBC4c
rfxEXfAFyt7Cf3MJm3paKQhzW2vNCIeo3HXWTpm1YBS7aocTcwdN8piC3p/yVItk
1DtIbpayEJuUR/9prgo3cltzHb1yrIbaZF8UCIvqF/z61okXRJlPrkqBmgjCiJAf
vTZK0L2gaxuWGWapse9EvW1FCN31tUnRZIzEVmqn4vFzKNE/141msYA82t+26KuY
bC4WghMbguojIN6teFD+l2nvJk3uxjZ/iEd+2Z1oVSI2MiHEBCBz0SRH8rxb6S0q
TBvEnVg9GrMX65mru3jJPsw+Onk1WUixOEgGQsUpqv5l9T1qNBiYb0Btwt+WnYnv
rRA8NWoR6Uf0FzvptFxvT4zer3GNj71rCdmEVxuVzpFDgC9WgsX8skxoSRfRfVpN
ubCZ4RTMJ2yGehwvmFNrBGhCu4hPnqMUpjAcHzfv7AzIloJlSIN5zVnEaWCfXKJK
ijcFiqQUF1xP9rW7jdYBTYJvZJhAaNaDBLWfwS6HgEBkyeSDpX1yJtO1z1c8MvXL
JblUKPa0qda89QLv3IXkrCZ2rIfnRMDybGvWxaEpePbLYYrZp+6uXPNjxdCdkXHK
9nPzUPsMcCGcU9Sd8PfiGFVMrXTbklqUmc9VDSlXVQTdqO7+sHYt66ebg8eu2LVz
yLS/7bI9kScUj0M5NH4M5MCbSFYq0q5MiRn8/bLZ8QMx9x99wH9X7ApwMC2rFwuJ
7XE5UnjW0q1vyz87KD80qc/fUHDogNeMxrDjdw5W+N6wruq3ypxw/Kx0afkwyDyl
4xKTgqmWevElZVkxMWiihELW+tcg/F2BtJ14BT5onVnHa3k8yePRFDxa9DgTmm2p
ooOmYORIjM9u9teGJ7kNcewgTf2hdGeiV0lAYmrNtwRYmL5jYsM/27fbkNE9ubK5
uxNVrMFHcYYiXfRn1k0ZUZI9IYSMugEw+iHAIMgrHpVquvDG5OiAk6L6VlYm+o3d
QRjAt5aQEjA9uVAx4xm5Wx+OwmTy8xxALsxssbBNWAHYGccNG6OFAW9FViy92nTr
Pl2U6isO3K8Y6l700DEaScMp+eh+3xsT5vRZw1a5lYW7lP+e2bCqRKfrqdjDYiiD
d0Q10tGdJ83YQTpDe1C04Rjw1OeIerxNB57XU2qiuYZbt3B6/nsNaBdqSGO72zaE
xrQm42gxKnPeYrQlkIyE5MqfwfdiYx9xUQmVtD8iAfkySgRT6mNGk61VjlK4mdBw
R6EZW8lT2jBqzEtqhar2o6w6/yxrHtBd56IxBMoiKpTSC4TAYZTx+YWWzCL5p2N7
qw/HXy1m3LUReLV55DNxmxV/1vEIwjR3Bho/68cUeT7e9iqOU3Eq8pfwLRHrM/1z
jL4bW8fOlAXkkEdnRKzAIpVp4IodPnj2OHyES9gj6GpjpUPJUhqsR3WGha666kZm
dWjnyFDSyKq+BfU3hwVDlwF5jhpS31OjP/AM/owfFKfiFwUDUzdYLirHbmCJRhEI
jyp1wBAzIoz0K6lsU9qYSw==
`protect END_PROTECTED
