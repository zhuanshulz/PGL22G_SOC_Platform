`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f29BNlRKMgF68ENLs/IdP4cFznhTN3zfXPD76SqEnfrlFccnV6kQnGCkaj80nmtW
lHKHRJZelbQBqt8nY0ygXFbCNl8cpOm57HCj3JLcgtCE4j3gX9IrdrKvvM624pr6
a5Y/9A9LC0Ti0WB6O2Ce5GHoTPSP4tSgAWJ3lXWTK09P1fdXRGHqYu6Axc439Ou+
wXYouv1jrdDGEu+4I/6P36JDYPxZol8CUEs01l9Ohd9WGvJTtoE0D5s0e+W8jMbs
avLdEKfSgsvI6YWarFVQ0i2Ov7CrUh0ZrLt6fNghP7N0t87yNHhZ8avqzSncxwkT
hkH3XyWFxLIld393UTJfvjNFHz/qDLwatGqapuLcvtM+lvw7Lwc9RhbeukX6uh+u
/QmAn8gVTamRT+lyytPsok+h68M2DHCIdf7Q6cWZ7achZI1koPDLxd12+dXsOFMO
boAVtS1fmriYOyJ1zkzoPapC+PShRVmGUjrJ3BTgGgvfxMkBVz5eAGjJhRe80W1K
QF26v5jjyeTHT/1hMGr1ZOSkrSYYqAeIV1i7/c0JyfkdhxPiKIw10Qrb7vJRz0L2
ZX2o6Jf7j46Osy2hRJmxyxH+xV73PtoJbDSnDyKX/uRHEtQTVSwdEW5YjPKRHnvy
C3uI+YIUbYcuJgBVfkz2x+IoRWixddO6QlRgS7fAnsWmvXPAE9C1tWI8fCrKn50v
dhJhK+l6An+NzgxP5IY0Y8iE6zKk78+tJZVhRKtyX4vKNco4v2kwdQiGgqJ1GENG
6dl8tbxj8PeLBV9j5ZyTzkrTu0RItzJewczj58uNLgTB7bpgDWzBbJodjFGGvEBB
OLnRrHwCWWqpIA+V9Bsr/zA4Kn09nRazH1AApMG57KyZIEMzF8d/BEDh9XUE2fAq
w8sdWjtbh5KjjGKBTAKWAgXOBQ93MRrQuVP3iQdxBjGrFoq/G+ZRf6oDgSgW+QYi
20ZoOQFYprnmHmxQkz2B8PPwLKtddmzi8mLQ8KmwBNg2qyW5mI+cOjk1zbnISBdS
ecsankBSF0Z8JaFU4nTAFr/2NWkG7tnDIH+njKbXz10D4rCg0hTjIwlmhrPtxnBj
t+Ny/Xsy58pUmRTbXzJ40kS1yMTR2Fv9IimRhzU9iDF6vzreARw7mC6ONPbCJ91E
9kAQVXIQ5Jg6RXP2nLOsULDwaOCAZYZDFJXKsPs8x1VCp9Bq29tYeBQ2j9TI4dWH
YRBhXkpKat853qtBHXxYBZu/31d/36CWkpIMaiZqL2tqGSFxG/vWJLdF7lSeLDH8
nJgoAAFbrE+OY0N/KXm53gTFhto/avXn2C7M5uvpRnaxDcbJqxlv8cRJiHSvkmaM
inkN/9Bb9/OWlLKe8s9Bsz+8UKhl1pY61BLv8X6m5b3ZnUlmiXeLILoVBFbgc9jU
QQwFuKqM0w1sJXKVOTPHHOMHejqRGuEuzdbKeqMU5WY8GC4Wgor+wn7jRfSdJwQb
j2gb3dLx3wvxWKsUZgCRK/krLTgip4mTIaJOgSN63BMzfaDBIMONxwgfFyfJddHY
IIQjq+S9Lq6zyRU0tCi+XyvjxSb+7SAPrbm1bz4ILkd4AnfvnlXu7/8hqrECPJkk
2auEeDuQQo+7NFiAqOHXvzXsJ5ZjtaOpk+KfAMwcFWaZC5HL/mXIQAExm6YtRci3
3IP8BT7kJdzr3yH2ym10kLMikVMOlZQqCP4cxY72X3ic759hdgaddxYtBDnZPi4V
Mfe1Y7wK7N/NJJjs6VW2GefM6UgiG0tsxIjTzFbMK6/mVrMfxdE75OVfmoEUi49I
Sl8yXFA/ISRO9zvTcP+NIpFFcqNcl4apEc7g1etGdWNCPdOHui963TPrAAoV0WxA
I+d06vDPnbiiw44HAVP0W2TdESZ8yC4Oyv+ydmLbS9cR8cxYUvPsnSVa+szMeE7b
RkfxeXAiA6r9BqDbU1eOi9D63F9daIWxBj/cb3lSGRqPoze3cFiZyj8sikmRlKSq
MaNcyIebwDaKvn5mrG9NOYX96fh6MJMlQBR3NTevrFHTo703EBgT4P5e3M3fUzIe
y27mS02L7sQ4gL9qvl1YR+2JsYRLgnyjNw+/3Sih3CPJVWLx+njVCG9PZgIkNF9H
anOhNjSfn78Dd2m3XyQMFc+814abmYQ3qkIfLE7TphZnnhY5fATUSjK0zFzeuaMH
ZcumlLDsndTCe0BL+UoWJn+JgT8aoJIN1o8qxwV3tLUGnVzKDm9w+lTU7ja3o5op
H4M+5HHkVNsyhSnXr6MZlSzX3tFBChFwUISrJobPM90n9ZOfELKfkAHmYDT6M0YD
IDEYt0IwHtdKD+ADGI9v3moBwH/dWdadFXyNB2aJtoXkc5fx+tAH8MK/AGuzvnrV
lw0QL+u4Lwc4sTTiZkC6CnRiPCYkpxD5nZZqD2XnTweigK9nty5GYKAnsWL4C5Dj
i8LIFfUqHduonRqlEMECvZC2TbVnPtWcMujMYUpOHGQoFrkK04rG42UVkQrEwZl4
Y736oCi5ovRWbPW4/ioQYiRQ7BU+Mon/rz9DzrqtGLZ5HGpWF+s3NMxC3qaxlUvB
lxFweJUmzfTm6wwzSlxLlqfV8PCRBrXaFw1ZiGdBYdY0P8FtQJDkWeZGwgtm7faR
llauPi8/HpqDe3X/qvebCVH5xFjY6AVLyjC6RKxniKuossEXW3r1TsgHrZKUKvhN
JgcUFICIrGhS1zNhkxv0Im6SIXq+/RttIPDYKbtuJVZG5jES4Ef22hq0PfdSm+un
QyRPrniV5Qh/0OsHzLBcyoOA7FnXEbJTAIO2gvUMRi2tAAYJ4Rz0QbRKYeBUqzco
6Cj0aUyVx6SwWBgcmsru+f8dljPhwIa+oxm0Pd3P/GDtEy/cpNcuhO2GaXicVWGw
UqBC3AZI7i7m5zQ8JSTVNjF8FCw/JUicEo+inh4p5ks0op5zuMtKm+kM+JLJeQja
cVeR9SFGgxICR7g969uzvCGEZjL87ZCNJhmfByyQC7idAhaL1ubIq82wZpuHBayu
k4JdP4mlnOch5CYoKRwbhSJTC8aDn9Vye1KQTSqw+TkOspqQgsTfu+JbBAYKBvJz
QJ393/kUPBH7EcbOC23HPQJr7ciKiP9DtMDkg04lFCwrvRSiPOdcMMGZXnOGBBVi
/hzWefPTXLgCE+fOx8sZ+WkCU117Fnfx3Uq3eLWmD8VSD7KAQdG0ASc1OXFRTfTg
4soBP6BreuyBjD3wgTa+Ga+ty+9lS40dFKzM1JbGvSqqMZgefGbhb9n+Y9JAqSGd
mhAdvDFnqPn3+Bht2vBShahDr0zkLCIMjINAkU9W3BVXx0F9twLVRNWPEHm5VyHz
iA513n+2AqjgQdKN7KG+CbeiB4fO9Yx50WkDfRC6+/hHmxtiO5mKGcgexHDAD/9p
mmKpqT3L10B8+/+lnjlD88sDq4YYaZhlYj2Na2VMHdiywk1m1G6PzxLEsv0Ilpim
x8hP2lpPiO5RiohgEuUIAOgaVVPMuqR5IqlqNyTVNyQM5gnXmrcUoFWbKMQl0zKR
CRVem5Ls/S0rh+tNBhlCJookobFb3xzcBwi+y8La8TKvL+vRtI4rkB2FjLnxs15j
AumgSSiiEK93iY4zHwCFL5hQLkTG0MdP/V83Eh8WTkTGVYWkSMao9w1Mo8roOhiB
03pRIoVoIv5ypl5i7E62Zw==
`protect END_PROTECTED
