`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t8LT0rqoe/AhxXGBLTMsA4kNEFblIXvEZbSLep/NvQEQ9Jmbyi/pj64vY9EgskxH
UZtr0LbyUUgAhXa5n17wHtXXCBiA4Q3hDxlFQ4pp6tMC2MyCACHLGB0Mg1dDkqKi
eJ2gS8Vcjr3SPmRXk3nwXnyto1RNpDdcpO2yzsWHl1ljqW0uNBogvP/9cZC4U6Lg
0kwgp1R4Zh/MBudB4wsGE3VFuR+I8dLVXcKRdGgsxM2OzTcEQ3wwSXfcPzgblAAh
VUtWXegvGw4d9qXpKYxyEfbUuyYi38SvbV4bFpl06qHMx+YbWQJo36KBmJqXcNjV
CPw76ISkRiTOM6ZodxaRJSBG2hdhC1C5b0OlFoLt4N2TJpOMRXwiBev5svWq2sRD
qAc7oq84a4Z+yhw6HCOlCBBRN5ELtyWxZxKIKjb7yghxRCfxgVHOl0qMP6CSmjnN
u05ZH0QHnB709ELJzPw+2JN/JPJlHNtHXHCKSY1hSAjesPcR9p93TZCF389L5c+i
9GanJ/CQrL+AwJ9sbQ8HJ+URoBWvYAceL+fukirTsUSE9RqRmNcnD0DS8Oe2E46O
ACrvCUkuFqw4ELGtgdaswh3+GGjpw54yiajC5u3pw7DMmaJIkJ0ZXRxh2ofPAqr5
Rl4iM5WjjrFf3bX78s2sr4BRiOoOzQ0ZDZ5c3cY4SOKrRxYKo2zm+344BarKWIUp
IG8Z0UMSlCyHV951pmeONWA2xlDFjaifqwWuiu8NUKIgf0BEIzd26Ase5EtjYTq7
1LzTaw4ely70cbLm5N+bdSXe+rfPwKTcSYDrvyagWWFYqrKCjLN5SYOkRQOD9J3m
vJfABzEFC4Rj7plK9xShN3u3xTeF7nDeak4CEHop1BCQ/DDDbjgooeApwGKp3WNW
AP0a13wZiLUtzIVqrMVSkJc48wqZbIynsubjrG1kQHHS5WXiKoiGUNT1LAg9l8XY
xEItDyqg3fGHqIQm9ycLyDNDGQBjGOdF292TQrKicXbaDsXri0SHw9v3BsNGpkKs
fgk2hM0FsnqavpdDhYWMhVL7x+QFQRcMU1chWep218VUctubznnECBLqLDUSXb6X
e7soKHKjHDEOygaahhjfUxbC0MQsOsoDdNkvMgwqss3kr4NydUj507Koby3i2Q+d
ZYnGzDVcDOB80FyLY12tnQ8Nklso4mv0aivaX8zxdDkmA5JVWgXzqfE5BVFhON4q
JCX0YNZ6ZkTm45m1jfFdp1kPb/U1NuAHh0SCAzaaoxB1ptvBqgmfFuvK7ybnKfCl
q702D8Wv9FqJCWfPS52M1j5MPuWQdQL6As1YfKL9xOBRlRhxEQgY55Pp8wAjlvsx
MJUMJ7pSdFvjZaB5zTokGeK4OVcKeVby3cYmTOIbIgBgTyJ3rJN1Y5Vny3htsoDZ
DXlDbXnWoygtA2RsqzMUID4RNHhEJVcUYp7ZEPoxlSRBxpq2tYGDoQ26dBM8oGA+
1mvS/JAWocR42KVf+QKFSmQzAPokg5NR537nKWdRkW8CDw+0P6Z7TAWOSxNzH35N
kgVpXpCI6+nFMgiii7uMNvYcGC+eLxSHoc3c6TKExY9fSIsNDfpRp9Mua2f8Fw4c
FTTv3h5qfGPpby2khA4t3JJIm6hKNj1ZVNk/uL94U5tJE6rLx8UyQgKKN4VFaAfs
m/Uuh/Q5zR9z+i0VnuBLDFnYXf6bznwMx8Oq2YVUJdC0fYVifen57ovJH9N5ad8f
iE1/F0n4Vzlay1C3mMy7x2/nWf+LIwo95AvqxN9iv4Tk+Z7qKJPbp5IZ+uT26fCh
EkC6uwZ9ck1qSlS2obwoN6NB8aYEDUdSlGa83gGvSNqQhMws82II0a3T6lnV4HOn
9rUiK+8LklrnlsljoCMSR+9QwCwA2Wc/TpmGzbx1Zv7CJWWVsmozXlu5hagTvrG9
jHz0/fswWINB3TxG+cwMqSOh/1RbRPS9L4dYtSkTIzY/oMjg2fgaDLDpLJucHFWD
fSpsndKFmvcq34VRmQf2uJPE770bo+m6d2PQgzVgqlXGSEwrSax55penPeNv6DHJ
kTyDwlp1XB+qvAWQsugWve0v9SeOabzGOl9Tc+iZ0Dd8Q+/WSH4au17si1JUtRza
rygLqKk36CMP+mDFCFpKrGFujPTNEU3vHMWVYq+QxAGDnu9v5CMS0JOetrOcQgch
Mq5So2JbRQM8ZuTOXmjEgfbHKFlzamftOg0w7WFYl3U33+G1KUHks8xJAxf6Iz0a
0MHrL6VVDTEoXxcJ5/T1X+rxrg8L4FLmTNLNtsKl9k3C4Jm3JUjPFk8H6MrAj3uU
fyW8Pg9aulaTCMop4X1MgS8bL228rXGu/EhJU/001MqnELRGORo4xURp6fAYivj7
/AFDeez2ajO+eLWOXBPJQjq6kuw0MzKZxrAQ4yxPG56KEKi2rnDydLksB4X7TzVa
NuFQadZ6Mp/kJlhq/kRRj0NWcL/65jHJ/m58+7GapdBQkEsc8xlhiGcf+U2CHzsh
Nz/+ZfK18QxgHd06E5d/7c3b5v4qHtednaFkwYErt+4/XrKvkWvIceK9DhpUjd90
vMiub0M7IhlJFckpoqNq5uuvxGXx9onMRL/nIAPtDAtQ5W2wjXJuovKBA/PHbxA9
8lQ+H+bZ7VnstgBs0j/bTJOYrtjrr7+3JuINCx8r+mssEUxOMrSCtzIGvZvKDu3L
BmdOlsI5xQV/azs36iQnCuwqRIu94yQJsIFWRv7gUh8jZGGJwa6fZ2RyX4aKcJuJ
WiRv7gQGiRJVb3S7bWi0och+aqT7chVGV9hGqo6LInenJf30WjssycE1KjX0I8Sy
/nvyPocrlDnBWUGXqsrieP3ugmg2COsB3maMOX1r+BcHS3Q8wi9MczT05AhcIUo8
8IQMiYHdmCEy3yNJjuXNLMCKCBxx4r6tdiXZsxRfPoF8MLXQpILpShnuBygLEoxj
0lfo6b3ILavyYqwpUrJRTc4rz83oAzN+HQ3hxTEpDGr0rFxE/mz9gNOAo2tQt/wV
u22nKSCuHAp7+08dsZXUGjqti4c2GrM9Xun6srKbWSH5b7k4L4GO9bq0qp1//D1d
eB/YdkpnWsP7YiBD2vAPdil+MC3/TuZ1bkE7LiaiitRqC80FyJsBXsdTEWIqAji6
o7/H7U12zceJLC47TJoOiaD7qg0JJ9lMHcjq36ELzldqc9xnN3NZ8zoE1qCMVmm5
80L38ZCRAjg1fq+kv68uPAOlAlCOATep9q/v242SNKTv0MZhUGV69PcTgnjTCONt
CYYe7ky76yaYaGu5M6lQj4LnnxFbPg0z74JkdvcobsWe+/bj+8eJBsNBJHGtQBwb
ybPq/p51A/QJNpesyrqrs9Rp9EzsQgH/CJO2J4bxfZXo48KVBjV35i9AFZtnLXTN
1KjQ+krjqAFHzxCD/afzWoOlMJpLq/SMKXgrSMlDFcYg/0qdxLOrQm1XRSAx2Qow
VDub/rdWLv0zIt2D04TzdGzpqy1Yl+6V8fN+wqcGOaPtBV6CE6V6OOTS31zHPxUx
fqBodLNspfRpzHp/UkH2Y+I3R/W/hId8asefdBMB2bdVumyuhjEmh9i5oFeCXIil
v5uAFyJ0ve8O664Y2CAI49EU0bOXSI6+BXO+4xtZRa1JysYt9uEMOY1AlmQIWJmz
GnidyeWJ7lKI26O9R0Bqe0nbgVnmuYq7droL0kQnqcJLbqSqiERg0WdlMY8MkOsn
LDTc0uHHDQxCzi/F0DnzY/VFK6kJtdoqjEcnnkJKJ3noq2BMXHn0cHb2uqvXiWN4
T3GwEwxHF7dCDe+MI/CiBVMSWqVltYAG9l6fvfinYnaw2uZ1BoCsNaSCrblCdf5j
SAfoYUa2FaoW4sVbP7A1BVIuaBRsw8t0ApmvY8qBe0W756gTK95fHs2vYiJYEU59
zi7YWkjTLjCno64Ntwi+PdPFA6D7BjqgQ8PIJu8J3Ua5gAA70JdkyrjsXWf7s4j3
/eh41UUoJ+vKAaVDgSsNnuFVDwz9oifMpiE0V09eqoSmBp4MQngZw2sRWVM7icXG
HCIgnuwm2MNOT0SVJdy2q48CwXH2/5eY251skOO8wQ8mKaGZnw2pAJaRKNXHEG5X
gdk6UYQXvNThY1kObcwSs1QOba+GzyzMkbf7r3cnQjfPYdL4hwqxR8/sQOWTFWer
MnluTCB7RC1DWAMugYLPKq+yRgfzh2Qxusb8JgbJylyUz5D1dmPgYYx2xKaA1mlK
lhVcKX5Szf8cLRK82SlT8cQBi4HzvybW57va5l43rnyWaVlGi4fxnxLzCO73TcvR
sm5xTwn+r5fhHjp6nL57Wab9QJU+9MY8WrkVpbj3HnarUp8DEq5DmGA+F5vpJ/8r
pMAO9tReD89BKgcKvhRtusAfn0USTP9zK4PQb7e8XXK9stwGM7JPFzOtG3hGtyo9
qsACaG1qsqizOaXZYmUWZqyj1LtjwJ3SQPju8/lALv7kyYVJH08mwoNBdSJE9LC/
up9mtY3vpFkwjHShsibDciqCbVC9QhH/a2N83Ah/irtYBJzXzugaossLdDU87moT
MFP0QMQhQT1vKWEAvtK2+ZBHU5kuheEPV76APSinEnNX+oGAbVn66svKKpWZQH1B
pThqmx3Y76TGKTnaRbX35eJYYk3DY7DD0ata4GINiYlD/jN13Sfms3VQEe03miOB
6OJ04m5PckY+aA4PypEmg1V+8DcrjPfjD3GWYMiXPZ989AxbALce7W83JGQcs2oV
Ww3hQtaXLHz62yRU6/BNatu2er1LqFzoGA9/DRNrjF9YgOkEQiDO1plho9rATP9U
YXH2SFZRp4GpIEpywyj0FAs3GpeQjN1zx4ncXLohiPNg3PZTLSDzV8/bYCaXz/aA
Qd4RtJKyhF6G++awTa819atnkG9NuaDDlm8ZnBMIzCgkEAz3vMXNyW2KOSzPUiSg
iXCv+hM2EMsVHKD4rBoHD8KZFTFAEJHXBzAPusAMjBTOMctjepJ0umIGzcBQQBxR
pHzg9oa9dUETWqeSNxqK0d/IHN0AFY9IJmAaZvwVG7c=
`protect END_PROTECTED
