`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5JtcNR5/N3NTtECQxGupDqX9hq8Qc9ekN5MtVwllxM4vZuOHEuX8euf1Vv/H6k5R
8RvmGKwdS0ksijXLv8zp2QIoKNiaDZD7IQb3gK54lATcP0aS9kQiyeWxEQpV+VJh
y2g3FdGYn/xQ71bW+0Aop/B3LmvnuXir4XuWNQR2SLNdjq6uuTPMK1zjXYYkNTqA
TZpti5aAYc4vCR/hS/C298NDfutREDl9gIdkwzf8l/AZOUGQTZRzp6fBjUMskoxj
Ux9CdC5Z5FeUYDehgsNU+ZFX7tI2Ar/evjMpkAcwsNSeRsg044Qy/Lxw++4WPiba
K/wNDMRtgwyhQ8zo8CLYb0OEJzKmZtupzjfGqV4M9Kz1jgdCVsWPNdayV6x/O+PH
SNeKA/r+CRbxMHH3wRt0zsH1adMV69zwa3kynQNc/4IaTF48qxitNTa0DQ+fRDne
Ks/0ZjUflfYa97KTA/OBuXoX8XkzOC+I4OycfcPgOB1qQm9QRjqUOR0dI1soBmM4
i80HOQjONQrqfWDN5frUXy7Hr8ybUL5zqDbCDn+Ka4kRdhPu1CHvz3SkDzIY0SIS
awfxnKx81f/PhLlRDz5UxssyIxjHb8y/VoXmNy98PtNsVfNSX0hMMkZxyvCLr0A/
WAQr3dXB9u5+LD9n9e019SszUzvXuR6HPbB03TAb30PNlKaTruYZOsgIqKbswSBn
`protect END_PROTECTED
