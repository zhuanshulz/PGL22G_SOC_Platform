`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R41Oj3ztrBsltURXG8qycik+HUwfuquBHSBWNqm183Iu3FMAMg5lYlE7B0wZts9A
uMDePcJnWrK46O85W4N85WaAHfa+EcRjUUOtzN50A8a+eT4psekP4DZDsET2p2wH
XczcuSmYQt4NL2QvC6ynInv0SOx0Bk5OLeIM9WB1Mc+rg39vFh+pGGeGitPGSOtr
tNDr871hb+FeaGFLUzNppLmwksx2ejM5t9KFy5cePYtUZjt2AaK4rP5JzWOkkBeC
g3tKJdVk3hv+Yyz049Jc/J0fUcG0tTyx8oxNuc7RqEgX7Y0Y2WMY5xHyTFFPwQ6Z
bV/SSgigOMS0IJ/+a8qWJQYOHFcNSwitJEUeI3vQWHgfbV5IRzWXeyQgp9YrnqeZ
SZw+ZRrTcFDhTigKXMFDbGuzY6Bih6ZnYBamolR4nZxyM28/ra9nupSyiXOjAke7
M++RARfPTGLW0P3sq5yqaad5e/CMjNsxM+INM2NZOajP91aG2K3stjsj8xrSyEaP
xN4JM+39YH/KF0pFxpdrd6CYFDyTDfblMA37lV3P+U6F2817b3OSC70X9gILxMlD
/+ce62PfAJ6VDLwL9/Cf39QG5ZTxz/DAXLRYV8gBf0FjdmuD79vFL6G/aPob8PCz
WCbkoE7dF9COW4V0WCY9BMy6scxxrQ8eDmdrpoJCXqoiTODLdoT9v5ieOI7f3/Wg
WuRIUle7zpjf1qVOrQXgHDzQq4OzM94PFa5P9A/pCfCR38k1mOmSUXENS2UMscNE
yycX/4hnseD9qS8+S/gh7PIf2fknuW8MYHch2eRcRMMiy8KTmfiubYY3ur24jcsi
rTYAe1OYq0NLP6xRJwPyDSRPNEa8It6zJswl84YnbCMYfzwopFqBlsYTubrd3LBc
QjyfW7jeb1LWqEt3LY0apKGc++F+RcVTnKeg8mJ/sJwvEFOofJrDB/wHrLEwDSTO
9YR/2ktMXtVVrIYU7TR1dDE5FgKAX7C+N3EWohjEIX6W0g07ePeB3GS3QgkCe2Lv
y64gfLUkSJtehPZibi/yse140wPPF28sLORxAHAl3RTtkA4pq6sMgHoXtWiby+uY
8HM8X2rD1wCk21isNRNT/fKqrq7Uv6Re5ii1LohUhwviBtR+pLHi0gRajX9qf1ID
uggHQmvXyHYT4owOclGgMXyK5qjgweF980oKQF9NEWfSOFzYw5rKEaHY71q5x8Sy
0rC2z3OmoHEpgRUaNQ1wNHLfUV1ygprIUAUV8RJr0hhOK9Ca7myRVbtJOrpcptye
kIbtBRW9hbzcvnVSMotMojWUhSvHPrsAyvBYe6cxVM2wudjdFE6q630oj/41N2Yt
qkDAdpJlv9AaR5GJJiOkyXYTISNdnqReh1WowVpSfMDArUcbEI+jpBMwONnsT2Br
XsS7EJ+xo5WcIj6R851gIHiPQj2WtnvnXm7ulxHqhZtCywPvbeA3JcG20flIwla8
XokhnDRGJHFaMmw1ulUNWnzcT8jpQcTrrpo8GV5ATXXicwAjqzHHDPn+NtxNL6/c
ZJ4Rj6esD/ndr/s/uKXXHRFfMGOKZkleknyvEYJg+yNQXQNz9Gt8gHvqfm5t0WW/
Rk+uphWYrAAcpVMuXlJ7u0VsxsCJXSB7DL8rJ5ZJhf340OyyaaAb+L59F20KdPHU
7gaiavyGsHBj1MxH2HSx2X0ATc4MxMFRZFdvodpYA0NVwE8MzD9yRJEzGJAyR0lZ
Rhv+GAJi0sohTsE55Ii0O+q0P+8hmAVumLlE72caWGJVuY+0ddKVY1Q8wViTrXm4
Ul5pHOEXCfXW9knRgwfcFBrzI6vwd3DtgXWpOFQ8dw/maHEWFC1bh2jyOahA9Poz
pKKT9/7EpbX/DfHLvKyi+5AF53lizoqv0MuIF46yOGi1ganKpfraBtCbHHtPuQqR
hQx0wezvcGcJRBU+1CKyYO/vrb++pbvYfR0k0bdQepre5faEA+ZQ7gQghUONU2Qt
qEH9+Xm9QuO54i3xXrfdUxmUx6d45h+d9Qqf81P3wD9xEqT2tRDnWrSCVvBqZ3Bc
H0a3znCnVioccxpzmGMhw25AcD0x56MbeCSFAgIvylQZ93g9Va4jz4T9u2PEnCgi
cDyLfa5+IND9KNsynzdA+b494bwFqX35pSoTWk53jxVuI8nu9WOifsZvpSJwzT2a
63791n2Qv5z1EbhbJni+c9EHYzCxA4tgX4RvQcbGECVmejXdkOF9qycRdOobKR9r
DJUNSLW3atT9AreORnaLeOGOC60BMQ1MtlC9OD4aq9eusKd3wBWWyZNVWN1T02sX
MwdG2YFH757NS1RgaSwiFo1CdWPd0+ImdqFqRW48GqG4KV5KiLmtvha/MtRX6x9b
rLdMUYnyPNCJhLSIN4aSxtk5rwBlrTIJPoco7U3/x5aHjo1l15WX8Ok9eIbgoET/
L1tkP6G9gfnVjlWMObDV+IpztUzocHtlIrAw9lPS+odKzTETwzUTy56f24wcRdsA
pW8joakRkLzbSytFatH/1OSLtIXxY6z4Ef8iRZyvzg5+b9fKYZZ0iHa2+35wseUH
qgvGXjXHo7YBWq5NW2kHkfNAwPhxyxkjaVJoUER9koZ20mnTz+PtFlHZhPuNNgmR
`protect END_PROTECTED
