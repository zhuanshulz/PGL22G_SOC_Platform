`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+D8x8BG6T6VPjlfyVydjRGI6B1Q1VKnqkppqxFcNRRoAPlqpTwRSVSNdJ9AP4kMG
Crfj4wx+iuCBL00ZTVaKsOSZc7E3cBa84Q1pzI2tzh5Wr7PjHbu7L3Q6Hk/+6ABK
74B+5FLY0ZILccF38XQz3/nfnTQ8DYV/hloH1K8AlvLLjwks5s32X2IS75jRrYVw
X6BV9KvNr1ZJZQlgFwCh854x1OP5VM1YrpW/U6t1hBLRvPXHyPw3tD/6ITsbdvou
wjc3kE4L1Se6QKZj4hil7LpNW2qOQjagz+MhlWxn6w3aaEVsNVZp8IeySrNzP7jI
E9mmz80KGAG7xilUR/CvcQ==
`protect END_PROTECTED
