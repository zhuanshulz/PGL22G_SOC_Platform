`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KY8TCc2qnA25wq+NF4suc6fteAFQ1H+GXaQSLJVDVd6l9S3QNd8TBVVD4mZ8d0lT
tD8rZ8YaZS/pT8fmuI5tj72jGr2sjquv8YjRoM+tVkr00JrJIyMzcI/KeaF8iSWh
hFQv54VghugNUJpObNSCzwEAD0B1f3sxJCywb9TQbsSSTbte5Sm78Q5M2MHA1UKe
XFMy4c4xa+O06NIVHBrHAnhZfGV4+SSvFbq6bK4qBAqGeB7msiDeVJmWS8F2oKKG
lZ8kApNFW3wjPs7GgAPKv8KmkKwC4WpiVBwtBDIe/fSoQ1T/ersoy1ept90/O+US
BPMuoZA5uBZBesLiF0t2qwiZUP9kR1BxWOihtu2c6r1CR0umKWPCSL+gBs9yd+x7
AT/1WG3xWkDUdtFJnG7fB0qwKlqbAAUa+aRumgd9SbQ=
`protect END_PROTECTED
