`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9+Filbaes7xch4+0QoBB/VV9zAi0wluJgTq0a05fKQ+NVI9tl/79OSwwGiexHu/V
FUQgTKurV1g69TyOQwDcQsKb6WH4HCzAH8bBYoa8v02HlwZzAOygYYmrYONssLEy
AFa1+DYuPhEanWgQRN3KUk+wkIJN83qZ4evM0vObTVRKwPex9YAhCBksoDAqBURb
vkIcSfNr2thi7Px+ipbzZoxwq6VnJB3paVD28XzRVxV7xv6kq4/eA/Ratdmme87p
Gv116lq1Qd2y9Um9UxVai+5eJVqMVpa/qfNBmBBjgEhQwVD7sdZeV5GkhHOz+mX5
UI8olGaXTPWO3vV8AkebwyfSa/eLntdsMvp4kjhrLGDMsum3a+RQq9GqlosdtalE
1qRc757t7SLPIWkxur2VPD7xV+Gmvkz//9BUfzuoxzWXGvJdCBVlS9Z7saoL1P4m
58oCzKIPJ0zBaoi9JUNPWUzUVrW/CdU7tnDeh19/+5TFL2D015LR0YtMikhAmXWg
T1+VEsgHJgajprZS5K4BAr0tob+6nMvAwGtiLZH9UtB/J/NifMpJZAXIwCEtX3ra
csm3OkIJS+GP+W2/aHwd5QrfBIeOjvuBBYWu31sja46gPopGSu6bHgGWb0zUpnGf
jl72Mu56r4OfLY5V0ML99gcM0mwacy+Zh+9WemVZ7nlS+38lH9wtMJObUJHjFNGe
`protect END_PROTECTED
