`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g1Lz6Q/BWqD8Z8CN2s2wVTILe8snEGluKDE3jiazhlYEFljL8xH8iqmMReA9/aFl
RRImXebzsUnMLcEyfXXh5EFhvIoXKt9UoQ6Jx3H+a1/I9hCPLQMbh0qp2sT4Pw18
CHFObcIn/Ing6tMv3mM/BAi6gxCy/nosSczhbEE0UrUH7nCxsu9ZhzVjkq7I3vvh
OLPHeOYLn4l/uMtrsZ7/AdJEJeD1UJcRe1IX+UOpVm6rjPByJj/xqV8ueGlQKDqa
5/Cy8Z1L5rNYGuBjsTXvJWQ1MTggLu5UxLrdLslMvBRnwIYag/NhWJ9b3RQbmZJn
oN0PKnsrENeb2CP2eqWjAMxid687U+CXUl5cOcG7QQK+MfHGFE93VQjbYguGWPBK
u253ILylW2TNzZipuw9D1OnrdQUR4/Sx8hFquHY+ZxUiPvftaAH6l+e8H+G/t1rx
Nl+vDxtvdJ+zSMbNpTWqTNfPlLxg8cdy5hL8267TJS7iacF86PiIBAzLTe43Vcn1
Y3fD2dU3iSpoNVHmO7tURpcwUvpPCn4R1IIPFO5OXRw2GamYf1zAPsFg2iVJSp/Y
d2mGzwrYMfdFVpPuxzDocwxl14gn3P+ZsakiXz+AxPsHkZ/ONOEz8FFDrnojaXNe
D/AlKWMUOKuAXtYqztvaaaf9SSH7N9LwaC9ySbkCZVlO0HMIdfsTn8jiIdbPNbhN
a+ISOPy9BSvNCy9vkKBxDUVpbiYZLE11YfqL+KmIllNXPZgtSN48iAMwAB52dWv3
5ufIktzmmSW5e9g2WunKLZVQoikpNgB5KQgpf5MnHS/DxO6XU7nB1koXwD5kwxZz
sRvjD2BtXrSoKW2fxcSHbtwZWog+vEvKUbLIJAFZShMwCxSlG9st/3kluyztzodJ
DIxH2UshXVl9BgoBsmFBWcfoBBelNYv9hE5ppQnnHhHxDaMh+q0F2f92n7BfNLFJ
GOzQu0I5eXtAiqInjAhtfpvbobIB2O5xcMHOo6bI9aM=
`protect END_PROTECTED
