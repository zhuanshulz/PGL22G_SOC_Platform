`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XISJ7os617tdY5P1K9KlKNefDsQOsgKEJFA/zOpdg5DhWnK9RQQ6FRA3NIiqza7+
toSZF0njv+SeEUqi9kc27uNo2iFKj3L6k6QV61Bke6Ue0NVl/L+qy+HOt6l0IJz9
qrwLTEOJKMBuQug8/lc85YENQ5aOaDXwg868282pLu5dDTtAWdx5ntlJ3v2djXps
HUn6qXu3y/8P1dj88WUjCTfoGYF/VmFWS7CwR2jUuCuyCodarGj2oLnLDIKX3Mzf
fHn5rAbfqTW+3K0t6tr2kM1VCei8xqwuFAmGg5UIZt/X/J9DCTZatGvcZe+bNtZ7
RqeaNlTyGvYRWTP9/WyzB/gO8zxzSzS5yEZCwRoigbk48GoHCKkW2E8dbrZ7mROu
XIyqYAeM+Y1LqS+r+nTAgt0d4oB1Il1fkZqiZXusgf1KlVmaqVBooDzfJMiOLdI5
mcAc8YjiOf7FKpE9kKnC9mes9iy+L7T0i8xtfjAeLiON8PDB0xfDFEpe6ty/ECaT
+bHoDzAP/J7iGcTki5QzGg==
`protect END_PROTECTED
