`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2edmuyBu2Nuel21p1QNIlbcSDrMBKrELV6TJOMlp2jCmZrm72dOb0Kt9taOghhzN
rXuti8+506jsX883Sw0i/AEM6wiWfbWhKN3KIMPg7hxuhRrz44OzxAZGtrNDv8Lj
5nC3CbxX3JLo9nmUCyjafVENg/HBbynK98emLkMi/VX7Ilx4R7C2GBkiuBut3Vp6
Dh4h89/kvWFbqN9sKwO/L6V5bA+hv4gD5r97YvAPJgOii7SOa7aHrnZHddar5ww2
V+sdLvBldqzvaXmsw54aLw1arPF8RV3WPapjDasONDvT5zXud2Gcf5DKTmYCxzsW
KWtPmvZZbEkuaYWfBhxo79qyAOocvuE2yTXDQqR2VcGmB+xMa5W6vMgqcXuzpHy9
x7ZvHzysfALktrLnT6bzrDNXETGFrdawZQy4aF2TLszfDJHRdtci/9gMNkW8s6Oc
Y4U7summ3Ol5/pCiNV7s2kZwxv6c564t5nQMnanbdXjI1h+D/8jlqoPdVnqjYFsU
ZkhM2Pq2tzT3pGYdgLhAOkF1AAt7bgPyXErIuS+5aW5Kz16Ax4CHJ/6Eeo6A1ry+
BYOhjXgY5hpNHAXt5ehRJ4E3HfEZXiMTanmp1vEn0lcn6egiIrc+Dt4zdC6RqnUI
MVDPJXf/X0TQQ1XDLgEBFRSnoB9T4Wt+Ty3tGn50uQxT7lB1dt6QQ6zukWiHA2ou
aiYsvP6YcQkeHlIH4MXhIznuKH3Jt/clBsQM1cMmHPebKKWNOISl9cTuIsk4rY/4
VpoKsxKvT3PQvCVnV1rovgpaneBq0MUD5v+Okjb3hYZE/QL65sJip2Q2dDQaHpw8
wJsQmTCO30cynY5a03L3o0vim05nGhDO+XLA5LcidvVwmGk9Kxu5RJBrzTx1VwFO
ni4Xsz21cIvogkFeZaOrMRWOsdXDCfaCEIXH4X1A8RzTKy4Q6CMc8Xi1gQUJf770
zRBqQO5L180eAiazFhkcWuUvWfbU7mIabgLdVkO7ekJi5U0VGjVNtB+6Dg0NK7Dj
2lggxZsnl2f55IWJFd2yY62Z8g00Qx/lt4YtyriBwseA9O9u5Sqfm7Gxbhe+tng6
2axaohMI/vNUfQBcT5r0he7VS7rdFLu40GTBxFWOtvRyqJXY5wMwSfwqDGWggobf
1i0SwHWNp9K4h35/iKIJL1m9XhmDczbB/O4pDTVBfC+yAbBG7DF0lYrhMFMBFqtT
RTLdZ2v2MqbACS3ZrdsbqIENshWeEH8X+KwJweztIwRL1/NPl8r+D57acOhMt1eN
MlTC6RD8nHGnUeORIb6l6fp/m3ec+Gop+5fu0cX6m67ewky88oTJ504GWhbj/GXv
D+43NfVzEKfPus/HdReesp9vJNWnVy7bzReONQId48o5GLbNwjm8aOZf0oT1aT+7
/EpWrEw6OOPLq+XP6zyEW+SOwmZtcTrOeKKzYZZLQLlALRwojkv72PG+ZtCeuBaf
LN0Hk/lScNsHLjQXclJHylSK8iaikLuFFclRwJrcuRr6izAwylluVSAw8eJ5SufR
/UTHzSmf5DlbZBgSl1T/wsKQBwE78kWULX6gJt2z0JjIJoehhd0QaFJaJV5X6VA5
ibO7uIcOZyCDKCRsfr2LJo+V+K4wJQEIv7XTgzz3LpuS7sfC9KJ0RPtFC6Qy48P/
hAh8WngE/8DVv0+nyRoxA0X1cyqvCwTx//lTWgGasMheQ7yXGeUK2SlNWzsmk8LG
981pZVkgHLCRybebQ0d4cQA/yOcW9nPCsn7LgHvaN+7Ij5JykQDBkpO5ZpIbj0Uu
`protect END_PROTECTED
