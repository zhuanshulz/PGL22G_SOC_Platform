`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QIkGYia6MW910PF0XiXnCYFsLBXL4QE9/ANmY/nx42F3rOW7w+jjta1iB7R28HOf
JQqS8ndCJiXAilftQ1ypOGGgqMTV+6w2MzDoOHM/hnRDkMP7V5k/5+lRewHfka6b
VPjgUvDa+pRVoRCbJVH90nRQNO4MQ79ALU6KR08Niu3/SU3qQcryGVm21HvPDCjv
0DdJoiVrbw3YLxTI05E447S73KNBSCFDszIrZitB3AEGVY//bEENIqqP7En+6ufq
Mncpv5zoKJ8jbxYdCW+rERgaXm2FRG/eSvxRL9r2IlT9mjcJs9xKNp19Qsndq+cf
Rt0f8ktLs4M/Mf00Wi4F/aD0iWyZs6RhEsK1WVtaIVbs0mMpgcfxuVG3OSjuQPB6
A5OX4876e2+LyumcHoWe2Th/oiVF9CS+WDe2k+FXIaGY7TALG1oKUisptVmIy8CY
xotxhElcoHoIOOz6csdyw5bTYdyDfFXXpKjWcSgYJ4vAyt5EPYKodfNnzO147nvG
JbCAHOnSSNWn73MLaBWkKN/7xGyOtOF9NeUKeEfyZWLXWhS4AnHcgiBZCVDoH6sv
Ez6Q0gCIR4cFNkczoCLR4quDnRWp1JpzfhDnzt6uPVy+cTzNBP5Mk5jjd5x2WQ3g
ZN0zbjGkJG5dyUuzN6OmW69cKOtcAK1yZJQIKbUddHDJP9bVlUfNK2JvO1rpDWpn
p89LFTSYW0QyE5wXVUA/bSxKMDxRY7DtqEqR/9nA34d+hsWixxY4byFiNOqTcao0
F5aMAoeC9Pge5VJn976FsqeHxyKDxi8hum65GWj7Z11sRwhkekFF2IqE51qQsBUs
`protect END_PROTECTED
