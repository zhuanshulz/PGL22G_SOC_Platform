`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CxKkVJSfpUeAUcWG1p951AOVJ4Cc4CjVjkoIkUNq/sMQ8WUrzlc2gyC0JzhijL50
mc1vgZscY77ZTvSSg6fJwnEcWKy3erkw9P6OXRwEi3IMKV8aNyb3RNl/W/C/Gx1A
c443//0gWnvySrN1qrXxxm4+rgpCCl/SaER6np3nLBEwnmdLGu9G+T9V6AzDQ5EW
f3xV3SStsx+I3GR3gxHMuOl1YY4Zw5ax1l5N9PrI3RDuaP8qw7i9xOBG9B/Zb3ng
Os6LQsxGor+vwPdU6W5iU5R6iPdWsGw7YBpXPg9tFswq2W9ZmBs7Xank04yC5i35
lgizeKniPY1RhD1CrtRHXJAy0KZrjOJoLwhetR/FYpHOccB4yWTa3J+Lz0WKanB1
pUU3D83lqfqCgbkD9+gCOVUUeo1r1qfNSrrWpMAnXbpu2B0F/XwCC5A2tO9GSjI8
Ag1oZGUMbBskSqkVWYs8trKJVoDcyeyf7VgrYbThH69bmZMAEXcC9ajC8FQJQE3r
`protect END_PROTECTED
