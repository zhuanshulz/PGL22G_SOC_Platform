`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
599ujLUUdYWBx3Z+e2ZOHwi9nPSzW1dgH20PYjbFs30g2KG0KDdIJmQTKoeKr17S
jQoJY2/fgjzimhfZNBSPVzxoUMm9HgO6DD9Aktkaz7eeMU9iSzmdpYaE4MF8S6D2
+r5FqDXsxRjf3w5NRP2iN5fm6cDdDL09o572qelv+4w0UpDW+gNG7tzv27ihEH6R
SMsjSWvuRoPlN1PtUGSqiJ1fLgVrI0HqcOjiGll3n/IJa4upk0lFdS7Py96MSsl3
3n8sgNRlhEagad7I1Q0PequDkapArwB8mYGUmRkQxkDg2JcWs7Sxo44slmgCnVSe
cUFDytWN5++R/sSgGHgCEFWeSb0fVxsVJ6xRtjXIAlnqgPxHUBFhSGmMuVruMZZd
+nONp6a9eYMeE5RFcfNLePcHaWzzPyWjfTuPU13pHzbK9+wSSYpqXGgnmBOUUYDQ
PVnVSw5p9qssklnww3IcZVxqwD+ViPAV4T6jzqTWhG6iI3D56TzRmVmXca/Cuy0b
/OYmVHsPMfO2CvmM79tp3xHkkBj5eYYwUv/9ckB8JDDYgHrAg8kUUODyvAsXU5Kk
jcCWOYfNzkiNBPFZe10fl5J4ml+MErgxORNJy1WWHjD3M/8BfXd1hSyzTC8JhFRi
IrvYrRpIS36+a0/rIazMla31GHe7E7wVG3UDU8yPbJ9psCpQer25mJKGff9kDNMm
ZL2idXm/Ev8UyAQtlz30SBYODU2PrMYzGtxn/ykM1SMU+F9j5emqW2SNaeGFjUmU
lq4kjFPfiqlWVFVCFr/ZMxfTrz6SX+NtMmiDKXMfr//KOBYZ0QhAvUDYPsJv0JJ5
MZb434IygUxzJzyaN75kgR6Mzy/huWBBnd2+unMlqkr+RaqJB3xOoM0tfbDSwsEa
mEL7tS42Ci4GOaENC5ZyJ6RsMrHsE5KqvQTX7Z9rq52w8tFyGYMnkGt2aTSobNE6
3MNx63wExBHJVsRjqxRnRLm8QNg3OH/7XXZlf+UzsPCukLHjrxr9ACP/sZdJPu1h
+OdSIu/ujEYe4K6BSbrj9PA3PxsPxKqlVNLkTgaNnP0ireb/q33fo4gLqh5SKuKI
E0g/Ko2GQlrMlyiJUPMBwHXB6ryixlMPm1rCUeyvAOBKbv+EwNKb3zP3P8USgU+p
KSWVfAwVP/MziZ8nQZaDmRbukbLFfqy/Al2lnutKeM74jmiWm4hoVFgvpmaSeOPE
5RM9gE7+pVxQ3BruiLVVKSIGg9LthE6HZ/oE+CvrUdlsjvmMN6p5X11N/SEOneUG
UV1l4jCqoaDxObkQVmPYqh/b586Q5RIBemkKin89I8CaEegbw8+NTIWl+ZrC/dK9
/EsOKxl+EcyMdYx4CqkwE9yK2YT9qKyqm0NsrTCB3yBjdchqPSf5W9ITtPs9Lo2D
1wbdAraWoRm2cs3ETaCOGi7qCeutVhYKgQyqBpGsyDFe62xSJDYUC3RlwEvLR7rV
Ts7/Jo3CBk4B1ynlY0N/s76D+ZJl/o1OnhXPVyZ8WD8vDyDHntzDcYcHYejj548s
EsMdI3zZIE9MWalcUxL2g7/q5ngVLh0I2LqWstsgPQxTCPxVOSSmCQUEcQ5SAWnv
FkYrT/SZMelJyileQyS+BZ2+/YOu76akqoSBJEuTrrPnwq8aoL3GIR4p/8Ecjd4J
HUbztvBtGgttI0P9dnkxqMsT824BNGjxEtnyQTUgjl9+0js1HKypTR5COAarbN0a
b3Z0BIoJ+vw/m6KLa7zPxdf+mK3iq8UoMQ2vMcPUkauoPo8disqxUsFcP/Mhg1OM
4/GRI3Jh1CPSwNydCJZMSnfvgpc6yJfR+4GM5rcpae0ev4PPW3M1VnYLK+nV6ZMm
rKZGpQGVKqoUGuXR264Ok1nCuqz1zO37/gaxHBNxOtkY9X1ErCdo/AVPOy9gnJV0
OiRTPYDe5XWl9+h6qU4OBTb6pDxHvl9ibbkyNdUBCYr7jzbhcfp4H/7d59erIE9M
SVpo/RkTaoRP4eGVQ4cZCdPgIri17DZDSkvozZ5YaUZ2MEmYUPoDve+BHBvfr+Cf
VW9ipMuFBr8zZYo352B3HnVtJwrqoEWFN3IUtsSwaqHLmJJDFLXx3fVFXzN3Ublb
gZt1EAI02ccnBDrKLSy2rnw81PBOwtDtnhd6fwx4H077cEGuPhyJDwk6hxLxNkni
zrv63XAYEyF1qHPhPybZ1KjpJURF3cFsxLO6EvxNou30AgBW1UKOrvkUgv/C+7W7
4nmx8aWdRo4uXdMjfoxT+d25p5JkaMuDkkIYNuNZfYz4CXLyB9RhXqS7vlxt4E7/
9Kdr9guqX8GRvjlzHh2cdiQxyngYWTPVnnTavZcA7OeFL3aIewLPGaBUZC3y9Gkg
8XokskOy9jUKeCfzvHdP2j7RYuXF4F4HuWqmuP8DS+9emzfTHl+2KF2qNYpFuVQu
hyfA9WyIHxkM/2ye+/JvoaJZbSFrU43QfABniBC3P7xJACgAs8SJoB3yeoSLhpnp
KZXXB3RMey4GlUIIFRke+vz7JMlqkGsJ8lpW7UhGDcHeFJ5ZQ2stpD8t3H5uqZoY
o6v/S2uf0vaMrOZYYl1PYAjSS8ryCtRxTASmJ9NRHUmk5iJ87cNqguCUOmt0/mzC
HzTtMftB0krXDnv3QrmLZ6BA/g13rMsCAQC+0jXSxjzdXdyogfcoRmXq84b5qqMO
/oY/KsfRbx29LPLO4SFdgHWFjFt45Ic1u6gIg0ZEigR/u+FxTnCuBHME0uepYo8L
iQoPvMma5r7JguY/xPYo0sI1aRjnI7cysiGQoSmyAFjhONLyTOqhNxaRK9CQMK3S
blzu/wW1KKSQxlyzzUMQTFzCUSVIeDWWlFWFsxw9cSzBB9jdAHpQwjN0CP8bUZdH
c2/w6XYo+hldBJv9KZznbs5ro7hymiJqzQpQgUzzhuR3ZOBGa6U0yHcmk4hDdAT7
XJtGshG3P2kWcvdQnWLS6EMFSdIj6hMs+YRyk54ksy8035XWOK1NicVHyGl1oku0
FNyM3CPkrgE0ZlmqUeLH4M6ZGMws9fwpYXhqom62JU10ITYFTwbX90kVnwyu0qJF
vtW0066Rauet3tEvrOzzwDEyZj3Amq33jbUFXKEQn2cu655bWhPWx7xCuV5YzPEa
QJxs4xav6Lb3ct5nBrvT23jszYI2bnM2/18PEshDZAchiXI8CmZcUMyQX1meDe/z
aV396jhTkP7kdXXwu8LCVhQ0i2rZ7piqZdOn0u8lh2WjvLI2+TNNnK9Ha/0qdeTB
9Y9lRBSz5ngwDBPC0CMhWhSfnvC7U4S7vRXqYuDM8+0jR10lIi60y6KQEwhjiVR0
+A2g5jOcRZ6Ps70sjLbId2h3JiqVKl+8YciBrt6JJFCdDgf9tdZsY9gQnS5ZQPKq
sJz1RwaHYakZJCBrShziLJ7xtEx/zrXqfZIBgGFOgOj7XxwIp8/gt7TVht04YQEP
kzxMyLOZ9hD2xzHr9IdmEsixmx5tb5Jutjd1RS29xUF83d/f4cnKcRdXvxdVdD4K
KsOSMZHDlYpz8Nyxo63Q/oipFeJE/7QJRNfS/h/CPOLugHupxm0Y22VSHglkHlWM
4iLAcJP6XJ7KxByfbJOndfOGAVao35C5O2FXxnoFA+DSOVCmOtvWFB1/2kl4C/Dp
QSPEKQ93LerjqG5BOACqHYHNqQD26zdMJ2x4zlC13bertIiqZYQPkAKYqZJPRXig
KnrCM3k5YGPKyS0Pcf0ohN61eB7NzLzKHzgicemhRAypkEVdJmu4wUlZG8qOfBEG
VggWi5niyKhYsjwh+rMQuDfrpPe34t4B+cKj5f27dkbT7M/fBYCtVNaAAHY737P6
YO3VmxQlMJaiZuSfheMdbLeOcn8ataFp0u8AzC5xKr1WoIqu9fClPz9JJBjjnEh/
1vzm+rnwb/GCEVsxRhL/tcstc8lJh3aI2i6lyLO7gHNn6t4C5YrHLcPoJuwJkZiJ
BzthI2EACPYfAM41B0HHu6Z5rSpuzvqmaOSn/EV1ZYqLDAne8BCJjixp7tv40mIw
jSklfGauALN799uibNn7MTz5hLjm6PK08fUmW0KngbM7wKvf1Uil66nDxnbZP241
eoLEhHy0rMpuIu++ir/Djaqai9sPtF+9BgaXVPzH2Mu1bOiyKXLuipKLUgROnvDE
Rh6wY5MqFi2wla5tRu+lemAx2pBNHSk6fxZgxJ5McXUx6PlM06/RSGlyUMMLdpkm
t2RW9JHCh0xyp2F6vxhG96rvx8NlPC/evdYo7noSD6UJa5cP72092CeGIFTmPxmJ
sSwyWfbRV/ICghpjkuWJW2wzRqk1j2bDoFS1866OQTITeyCFfTaK5g/ApN/FT1j7
9M4YQeFWpVW43NOll0rbw9Q7w/dCoF5PswMyqNAeVaGkVoZExLgnxkZvtqIbVKAa
QxS0if4XYVrnaRTDDZrGh6EChQpMYzbEqXyNT3vg3igwWD3RthCOPzZXyFjmzBJw
DfypvdTXnzLa77eqjbsoRDRsHsBePOdwIcyas6beP8ueqmtmFzZwivhLighbIZz0
MzsrJ1V06dvJjwThiRSD4Cq8Yon3PCoFdUVrByR5o5aWqpjq09j3AmUQFn5lzDRE
lohjKyWln4ika3xNG/VwcKBUmbHTeVPqQ6ZIdMSUGJOeHVjuKj2smc0ZnNNdscZA
`protect END_PROTECTED
