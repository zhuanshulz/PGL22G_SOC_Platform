`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6OhZ7iVutmgs6MwXCs7k4oq6BuFTEMLyXbGNJWKoDHGYZgzqFHNlwEsgczpn1CZN
gajdoA5Qoe9X+OnYjMzJ3nLKxWWu1pRbN6UFUn/Jz4yA05mBuLcR+wAcGp05lQYn
40OpuCLtLwYGOmHSnhyS/fvjoVvE4tSeNx6tr3mEPE+SmsPRdSVEcE2aAPhaNjgt
fjKwhrc5kcnJUjFkbMd+XOT3834d/uc6WijGMUMuAdBENXKPPxe6yTLlEX+M00PB
yTkoW1MukitB97TC6ltPyp4QlfLU0EN5iqje8tiHIcSzxHxE9euFMNtRmwgYM4c+
I7JBsAIMBUv9MwX4q7k+WARRSk14di50ZazebFicNtOJKsgp0mDh7152x+AooNPB
ilSJjc1KeMEiMTmb1nGnYmpO6Pg+T/XZ/b8pvwojh/UfkmjNDj/3jAnSm1MOAdyu
tWMPD64bNeYvvVdHewwZ4MoW3plk9we52o+BtjUKI9it9o252Ae8hz1OnB+Lbg76
tjGC4JyahIrZjUSc2X+YEzOClFyYiXKQxyyJwN7Xa8VZm61ISN10f5wZ46tvpnVd
Aw7f/5RZAkDYFbYCoV7ryBMeZQ+v3oa2t21XKUEVbPsOCfW+MBVQg9O5HfUIYuKt
6oDTOtFeS5uz9ov/YWzYmDkQOWKmuMzqVIqXkOccSMQQ3DZ02fVzHZimtWA15ZVb
Buhr8EtDSciX8hvsY+QRcVA4ZQj0ExFmdfPjJR36zMA=
`protect END_PROTECTED
