`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tz8paSCwOhH+lSlDpIVr7aDz74EHI/KEADHhsc+lb66GJScYcBhhQpZCE/rmIGuT
QEyHEnh2tPm5wsTIgMLlvbJLJIYl5ivRPQcHjNAbqYRzs+tgC+NzlOPRTMCodF73
DNxW7PbWY78KTQJUrqgxx8ueTe93yrBwtdJIWPK3aEQOsJgOCPXg73BKpTI0H6ue
Gu2rrLRW7zHccmh+vqjRNp5tdJcXMAU0WsxM5Pbxq8xBalt3aOfvbDnOF9HMgfqv
P0L+jvZ7YwHaBjgYbFSCnLzqqKtmp4F8pSgFyCzFtSIOZ0ZEWvd1Be7RMIPpzE5V
a4PqGKy8mxBXVrk/CdWSOGgvCQ9Jx+6hWbezI/TQgzs2f0tzuOhcliDEppgMBHV6
VHQmTi3qcIG0Sa/kQdVlaPnUrd8PBvlpCi+cFcNWFo5rSzmWNseX5IZ+5iWcxPor
WVGkAeUKw2fPm2LRACqwXntXz/7iMEVHd2zKQWutbURK2eD2vItQlDRM0LIeNkeb
GdfCTBrRtXH0ryoHoBs/TJVpEl3St9mhGdf3NFGneWcFXnvddP4DXM8yHxkYVzmh
qFvWHw4c5erUHvRQX8HshfjcdNIT7gwMCsNaUzD5adiTKG/fbB3lAoM/wEgl+B3h
mlUE63FFcou3fftcY5pVnGSeu9r3K7nO5jMUQBYDV1MqP8QFGpVweYRpxupjp9Qu
fO+tH0StGxpIjpfh+uAmu72bQJ/enNmQcy2m7yeFThMDyWG06br8eQGzmPUuqJK1
mtNglMjca+5JrgC8aiEDpiLO9hp+/cEMqGU9hI0EWfHijaFt7B2tJ5EKWygOwMCD
p+ua+SZ2WdF4jYXKxu4cbaIDAT4e5bPpyT/zn8WvJvWgHyKCVtd/xPwiEHdoVatV
MkgRkItYwNpzgBNpKYB6Iu9Sr7ozOOlHGnF9H4zBhOb7IKMydCNu+A8syo3vQnhD
aP39fvZ2Db2AB3VVTYjHd8zJRb/YDrMsKTudfn+xdbjnsHfJZCZwl0pnW1eqv6p3
/l89q80+Mo3nEhEBsMvAu2GlnKlLOMBBaYvsjEVYAbUQ/2ZLwPzXrhrLyQomwNK9
nshbeJsXcHrmNb3hFBeKaZHhVFX76cMwlE5sLli4Vzc9BKq76ckFsmVzVdo3Fkr5
iQczi5iWdUAe8Iivzm9COrPctb/dGiIIeOMYdReeMBasNF/nmS3N606K4rsRSgdT
c3gQ/gTAoWn0V/a6K2nfMtE4jbOwNFmtH/LpjSEaLYQfvWfQGCmrUylWZQF6WG/f
6NwIWFVvvebUgE1AfTA/jozyUZiCp/b0AKF9kM/AM9/r4kDEzqUSn2rRGEzRblHK
HEnOWn0oA51+78hPi0zleW0jBc6afJoRLllE2bSbV9Ig7nO8fWcdRKUs0ZE/8fGa
E8zoSqqoPFQsB8jcaDi9kKUKnRn3iPwwIrCewEK6UCmoZe+Sf3BLmDd7SByuDJqk
Qsf7HweclVmatkn9+wMWqCRUtOykdTY7eluZG/2GvlE9hbCYp8ffUKFsvcC/pBEh
skNmPIRmIcoLo336IBUYLaUPtTpYehU7gukkJkypfjh5TqizfVZ6fvqd/ix0pFmL
xxkp7x8RUY1QbC2ZadQKaYOG/QRCiatOJ+E4HKJZNUprlbVlBS6Ah9aE3vR7i56O
D74r2ho+ZGF1MrQ8cSghB0vBM7G/ksVNHZoG0kBbB81PGjDVAJySCAgUKiDcoYdu
NwoaRx5IuOZNj57A4VSVOunnC8Uuxah1Ol00g1yZtbzxtt/BtcnzizjleaZ7/ei3
ix/XYtgN3jQHicrARsf4iJLIq06mD8X9BvTYgHfLYX1uiFCPiSt6nqTOb9rWCd/I
2Q8fXgmDwufEs5owbPoyaM+9J/s3/i7fApM097VWAz4oS3czl4XRwehre9wZGbFs
N/lIWUYnC4DHf5INXiey06tAFwx/KZ71QkS9nT4R9oKMs82QshjX5qFx2hVeIzVv
tRrX4XFFySyi8cu3P5OSbBRGjsvW1ZXgRdi3+33RfdLJOgB9+Z7ut8U1OnyDOPSN
L41vGFP5UyrnVnMOsAKCcDAjDtE3yBg/KmhRTjkDB6e0J4kYLlJVk3kyCPusDPMX
e7IuiFLDaZMfIAV9PrsZsfbopcK+mYXfJymigaF6HhIBdh3QKZjBX3p3cuDMAeXK
prU4dW56he3L7tx9etaqqI0JE6qpmtruVzulMOVpxQTzcB2OJZ/FNA0hIsS7+Gs7
GfPT7gyi5qAa84z4euqu75rd9rrNmuXyhmMaqHQ0xP3rUIArexsTb41tZkmCgPa7
uNBYAATh5vWu3L1LoZiJT/Etq1jfFALv0kbD8GNyqYpz6Hz1ciVWis1D0JfgUzq1
KeYMIY+VTZQNlgxGJbJDe+h5Hiu0XBisGDRGZQOWHOT+tDFH86S9hjiyhe4/qdmn
EvzTdqNVzdv5WKz5+DhnCFimSnXfrY5mIeYsdMi2zvHnD82IUQTdSFuIn65evVQR
ZvNiQIIBEOwtfbxZlWBiOSb5m9BywtFQ6YII0txZhtvgVZJkTIow9Czp32AsX9qY
DmCBzhYwCZlv3EC/iXaK/vzKMSKZNzGMmtv3GhOnh4KkUQyOiRhJlT0ODHS377jA
3Ps8KA46YLkq/4UMe9LeV4RbnLBKjM/QWQdpF5xLuD5/noUwel5DfSmblhUCT7cB
M9HQzYPj+e8H3PP1QDkwthmxPqML91Kz1a0Ms3V64HJsNJnXnU6wnstrlWDo+DoX
M6NuLtCbLaFKpVE0eMzWSWk0T9FLnU/IpgFLrzH5AjWK+8YvN7CChU/960mFa0vc
FGKNyxp+milNv/XQyEIiYzQVl6Bq2uALMhtsbTOPzl1rNvcRR1wWFsTtl2jH8RE5
zXL9lhd7bRK03zKJruJPa4w32+ohm42eLfrBtDac/eewp0eo/6OwFxLDlNhlFgO1
t8WW5g/80dyF/znx3Sz0kyoswjHFRycJcJqiyEG0AGYYt4t8+4B84yG5r6fgJLo+
GWqkGEkJjQpArucfVjt9rmnw+OIwRKfPTDNpGBHoRlFyhAev0uurxug0p1G3DOkC
ME6A1rbAHfa/E4EArAW6BtKCpVY5n6uGgz7gg3/W0fc40HhduJ1IRIU0Pkv0iOpf
z8UMnJKxV//CF9d+qWs80sY2yQYA1TlTfjT2dVPhWJw9WoGZcR0RjFsn6Fq62yqc
btdJMZibpTs+5jCs4n4G3UrU8v+vEvLzYcKyg2yAt8s=
`protect END_PROTECTED
