`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sWSTI1D9zOhxpnGIlCXMD3BepsNuPiAe2NRg7gzoADFL7W0dPEmxwOqMGK9G/bp9
WMDCeNvlNLB7uczNApsDi/DqYxwk/KY7wBiYoDk/cvwQDFE6GLLN4vc1Tx9MWDM3
SdSa3w6L2JnhJkaTwvhrCoa0/XFt+mTDix13Tsq4oPL/oLxCO8pqJIuk7rdwujEW
6X7OFMusWIGmMiQr0DwVlyvrABYbA0jPx6kreempgfN1DUuWi6sVGwbfIPbggf4B
nsyMBzKkxhPLLISQ0tXSGnpXhKyPlpqYkos5CtXnUTndB9m+n1yZ36xEho7Ad1PY
mlanP5sdrHuvuiPGVi1rdMu5OEwXBuoruAJHHKBCBNSGU3+UYSINg8jRgWoXWZR4
fkjcp8QgQpuilvu7tuYJqUfeVdIe4n/+ARpXyzmho7J+pqY24Rr1yJY0JsM8lf0g
a97SPaUj6bGNfT5JRexdEEqRBqA1oDzLqBnBj5JS/0krvLgi+QpJBWsWXkZ8A7k6
gyHBJZpjtGw7gMKIxDXpl8UECYwEYeD2cTD+iWoON2ehWxw1QnglINOl2pWezcpT
inbKAdhTsmEQg0OV3mJtE++2DKP3Fpi574jM6S4YPzZjTeEzQOgf8VH4RKS1brRj
ix2yzptKl1i6DFRBJc+Sfg6agp7q6xQphcX9ttQvAw1EkO79PDWS3I/ebUELyQ/L
5cxPHR0h5infrGsXUQ5xqqD/lEb42beaClc/yBPdke/QVJILRAhN0jQbvr9tu2rb
i9icZI/P3Vt4250PZ27DeHxRrsp90uwPbFs31rKgshgvocrmYLIt5XaMVv5jw3zj
LS1l1VEK9BZFMnIVDkgVwihWvN4PlvkneJiwBCo+Uo+au3Sovp12PXwNo52Rq8Q4
xpSlUKyPfyxYifZSotky0XqZ1DcViz6KBsVS8MObOOVf/n5U+ylayx2BXdb3hpoj
/y7oQHc0M7XkKd+LJiVsjPka9Jf5RXBlZtySGUdVJVukg1ul2LG0+pBtaz8Oj2SL
ZKWu69s3IitcW0hv6+1S5Ha0bU3V+i2VCUS6Ejusqm+n6j1ylEeXaw3LrEBwWp2K
GBKk6tgmceWDrPf56xVEfM4Aac0EsK3Ic4QyaiUpz0GXDdgs16Q1SytPa2Gg+SnL
exs5J8SUzVYztScGRCi7IQMbJPIL4bXUb5BuEvMHmNDI22LeaVVfDTSgIudeUQMI
x0vDfN1rIJqPkTl7l1znty/ipqjcU5MQtHab53Co96FCy3/BOL/OTmCHm2loajif
czoXmia5ceJsAoK6CQWTAx0KXRqyWJNLzqa2sFvvbP9xxXXneN3CIOxY9JucuyXr
Zwwbv8/IA2FIA/vpKDrP9xtG8eUxFwnabzZZHSpLa6KG7AHlng/t70VsnIvt1O89
NiaKsjS9h09Wkh2bDs/PtMOb4m0chng8d7YZHLr1s8W1fQ1WGI98icpXp4JjySJm
OZ0RsNhS+pjwcIUQCClLyXAkCgDRxejhQ/gbfjIY5GjzvBxeQE/zUZyHI6gUqP9o
8eh6BuTLeQMJU/rBZXyUbVa7gliHgP/hicU2tYRjurDr80+veZ5jA9rdp17KRzwW
lUoTR6Qj1sWtXtojSmkcpOYKZKbeufB939unU7YmeCm4cNNDT3fP/hk/3fa1DK3g
kCtyJ5McivQw9tpeUbK+M+wYEJUgct4X4f4NlWpzOWV8+mHSB2xQGsstVkG812lC
RmAlN8JBGwHHYBfo41WeJ9SSrBj5mP7V7gRwoA0tpKv+ZY+jCnH3aXHHOIWiRcDC
y9BzXS02W5fwnHLe4XuEX3XBozzHE0Cc0rLxizafbyLXdAqHExi2CcCPfPjEVqRu
rLw8H6RMW8FpJJI7uLl1cd2J+Z2fr/9C2W9EQjbEXbIrimX3+QjYhytdBwfGk+Ou
ArgbZl8oKoSeNv7GYHQjltdpM/p0CPsDUd9MbNdJWWPD0BpiNfVnoQ/o2T9xuflG
J0qjGS0TP/UgPv/O8UZ1U3pQnThjT6co8Q6JLyTFEGBGEn6YO5E+tlBQMzW4dEVE
8YWb3Rm4MReB2Tu/LQmw32szqDdGB3SJL9/pNU+rizeTgW4Yuyas0v1OnoErqD8W
9iyvhL1gV7+Kn+JaWnBZFOCdq77jUjKQA/TPjiWKH9OOSiwhnroeeyjRlQ7m94IE
3N9l963Edl17gQFoEkgdAofnKP2d+NqM1MlEyd0nakg3rRvrt0rJow8gKaKkBamw
jhkLdbztjjfcj9bcvQF3rN9HUb7b45YSTVvEPBNGI5DjfJH/eqpL6L4dwjP3//ef
f0b3WuXkdzUV/yElFhKo2gFmoLNOwsU0SSfN74Pl/9bnCQpT4mJHc0uR0p2Qd9M3
+ZMh2y0nBcQrA+yWQO+AgQy0ej27pv0FeSo6/I/D/uJkHyT6M+7/uxnME3Oabj5b
UQTprCi9ypsOeU4VVX1z2t6ZjELDCUM6YFb8Jy+CshWYfxia/Juaxamau3gDsONt
AJ1VkOhRZ+9pw3qylkvHRzNT8ppRR+W4eZsCLOoUvQ3dOGs0TyAWUPemxZyjl+si
8+q1YsueIV18YKwW30XhqXw4aN9pd8uXMf5uQHw9EHW35uwm/O95isyiRfwrNQ4E
l1F8T+kWSIMsY2aS41lNemvzhD9H6H24DLlC+GJxh7+w/Eno7BW7iAxlshIb1e5j
xOR4pMwLvJE0amLHDA/XQ3DGCOwXGwTHGksbXE7zMAUOkGaeIC4ASulJh+wRzTNq
3c3Y6fiQ5wp3xX4sRQjMZd5X9qH51vlCASyX2mYULxPn2ifsyoKxDqfc+FUrzcUN
HCdDzUZPyeyZde/H+e16REcpe3ERpJHdKYP2FyFTds2qNAUdVtDgSpVyBFr4kw8N
6mp12RykboHanEUQEKGp9iJsElJFS7I8bExmzIblmfg8PkOjw5DS4q5eNC850zg+
Vbw+IcBqq3BPBG1o9Uq2HD5MSvZ3uSJ0FTZydIDcvNexCBPFlQ/zVFEI3wmFFzzW
vmN6y1gsapFx2L1a2IN/X+x9QIWbe8myUP13Z4bP9fpfspURvy7N5AIB5pWqwxyb
0fSVXhfMDQmUlM0QY0pqp9IXmYfvoPKAwPM+S067SFIolySd6tDGjiUSvhcPHAY7
UOCOGP7Golmb9VNpQY7rBij6QxyHFwDUSiO24rsfH4gNkjmtxvAy4lV56Iokojdh
b+CagqEdmoTdK+oqtV4e/EaIzV3k7FeJFgipFq08jb3cRiI1Ku2X9KLVsOw14Rw8
WbYWWmqpb2JAjli19wuwE08uxls31ImanwGPVDwJCuPkZSNW2nJ/Mne67Az6M5UW
aRxiUlaAvt0gZq5TX5+R+Ruqx+Sm/R2YET9/uSRegtsM32njx1xdGr5TYqC8ou5j
pYaGb+o4m8+4d/I58WvIN2aO/9Hd6mWtgX/qHIHDrEQyfeSsTliezCFMJ1RxU+3Z
rEPME9LYAtjP/UnxHvTiGbAKNp26v+4xjP6sVAYx5PfeBJBNJyCQzsF3qVzmDA90
uiX4/m+hp5q9Pvz3r5ODkTKUy1c8+ZU4lMcqnWlCPiy1p2CYSIwqYfZFVTXzcVwr
Lrt7i86T189Bz3F28kfPOPjsqi7idAs1hkaV86JLbOBtM/VE9zRLWmi+qSvesA2/
a/zUL38CjyYW2o7alq8nQJY6jLzhq3yoSPC6pfSVqaB6tzybqj2svAd9VZmiDIJf
UKUOZV3Cqr1KvvXmOVGaFgj3NTF3umEA1lfTqqpcXFmJJuZwn5iKLs11Kjk+5u/x
oYBNpsCu/jVDiT3Ui0uCD58gbgeMUXWysVkzUTyTQ2pQHWbILMWw62YrWbKdcirN
XP9O+rrR4ptGjBDvjYcOq+Tx5XEhy7ro3vD6g1iHM6aPK4Lspx85486umpY2DIv/
TDPg+GGz5jb/dJMivgKip9WBp0QCwq5+iWNZAxM7+tSPitKKMtwjwOHb9806bNgx
HemVZbeLbXdTfxc/EbiZ7dOpt4TnrAqpXZY7euI30bRpQO0LjFWeH7PaRfsHyQsX
LCc/d8KWxYUYDz8Dcjr+Y73DIEppJH73wfHSVgL4SovsN2/OzQB/uE+oDZkAFoEn
nsHFayE4O976VAceWiaPZJDXn3fCowdl1uLk/xemkB/emrUDmCoWb8Vw4LKD8zts
PugsGPMLrUgJxoZWgl9le8gfcPYXIK9Ui5j0XERJxhphlhwd2vY8/omb86ZOhSan
RvIm4KTKk6jMMk+pyTbPZAMp8VHs8LWvlqAI6pXFfsSRFnTEO52dfcK5xTk43CRs
GdiENdIUZQg3JU9hWsowutGFuH/bH84QT42/77LO2EM0nIOvnp+q7Ellsg0fY7II
ARJZfrhiILvi2690ZnBH7ofZPJPF8K5dSn3InJr3D+tOpYj9U5ydKQthxdHlUOqE
`protect END_PROTECTED
