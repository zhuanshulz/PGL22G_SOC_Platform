`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HZ4d3GDI2iL07521EkR2Kjl5MBlYGZ/SKFknFA9J6dLSLOis3bI4m0EShuFnTymu
wenj5cRFho/Z9SoFWSGFe6yzZg5HVNP932KXsaRovdWvcG4D6Y0/bVJufQGTc0zW
50jFfotrWYvnnncoHszeSuTO8z1WspA9hoM+Ybwtu0LLmWG9u6uXOrIMIeCI78ET
q/eIK5yjEQt8ASN+TTyJrIjrTxgvtIWsf9/ma0+qiMGP7Od7DOnyRelAjgJV01OF
nTVE4ityBie+0utI/p+CetISPzSjWI2DitKbUp4mXeJkFxdMF09kYATfQtxAUHPp
01jD7kdnqCPSuJGjJ+wmPSYWrewtfwRyGIAiJPp4eLIabbNTY5OKuFuUNzNlCMje
VZwUywwyCV76T7AsE45E/cB/cmXKXFrMKPTjzvc1enpTY3UTzSffzeBcPoIrV6ya
T5h8S/BjubA/LMkJe6qVGkhUEslnHWxAhUJnXHg3V/PXkQa/1e/TAo13Vs38Qryr
4dwB5CMBZvFWGKoxz7CqfB4nqAaC+LLBVH0wUVQJm2x6pmiRGdqfXK3nxfFGYgS/
smhUdNzlrPSUgfNTNtP6gsVe6v/RFM88qWfA3+EMt43O5YpfRxzSlsxwbTzLX5y1
RTf4g90Z8eFQ1aoOVjDBMJcABFHR37uoBjWQ62+x68Qsg6YHI9UYqrRH7hVeQNyT
AMAAQSkNGiI0lQrfpP605Yoa/p0rI2qwL+luXD7SyzbnHQY4+hJS7nhtq36kXxVW
nL2UCTTmSAaj/hf1uojtvdQYP2yfVMNlxpSesj2dBXtXmqhDHgc15LhfT8bd5c8I
OiuPjIxU37T2UhuLIUuZX6Q+JwVL+VVsmZnv87tqVK0mm7RgokLrGGlwb3uQrsHH
rfAk503dQf75BPlVylSQ85ZIDDhnQey3Qrs2Sl0BXsHsWExlAdaH6WmKzSLs2nNi
HerECIma3w/Z6HK1qzq9V3npbNXhyZ8OSi0AZqPLKaMRAyfegKCWLJfltR/TuX14
RKTc/HkOfIzvxZ03rM22Ny+njxVoShJSGGkTkN87JLYyiDxWkN6oW+rv3XTccjfm
kU4sOMY7p33+2EpQvW2JNri/hnOS7RtRqQcokrQa5IgBVpBCf8QuZZk8Dnfa/RA0
QsiMvDkr8QH5iPoQfFHDDwHV+U8d7sxdaxWmAIWA0LxhNXPQtoRk9aj/SPbkomas
AndKmh8ZvwSJtwyAymnElv6Gi8da0lJB5Phs4kaWOfyU0In4lAxAxxxpgbMgy8//
bTeLxW5q53O6QhTy6ZSUUw1WOgyg8eVAomrZwjZGZwKJEOhIpVplzSqVl10tL2XX
/WQ+rm7EufQQmJkWD7gXNMgEh5arfo0FMXWN5+1FAcLHZX23E9vNS5Yl44uGfZhD
ZivrJtWuomjy8ukP/3HIfoPO7PGQ0jH6w07G6KXCeaE9xEwqhsGJel76XVRZWufZ
1htIp+eJ6dL1Y5p1CbQ4Trb6QgpjqwJHmQrfYDMtt43WFdTkOiUeLu7Dm+InLdD5
X1rLxjVFSW+kc1cyunsK2gAoUWzpcz39jFBcwwq5oZXZ/5+vWXawdku4nwt/Qf5i
ihqUrZPu91Z9vgRefRPLxZkk0l3bYD8SfEBVFTcgI6ooe1V+elmEJK498BI+AeW/
8cHnOSdoIUePKInE9LhvDFlCenhiXoMXFmrLfCrYOiumGg6O04EHxAxVPVA5URZf
3VvgDtCpXhX1ltZ2xd7L5ukCr4yagM0zGDHcyTKuOw6yOuP1qV/5+Zxnsi3+lnRw
mvBV0nUr/COuohZOyvSR6r1qIlaI0c6edSvQXYIWmVY9wN+fzyHNNkBJ3iEaRWND
ahDUV2unisgrDPFWpP2hrFnwq62oelEfHBvAZnnTQtTiW/Mad+kRGkjWcCaYxlAp
vEiUGJ5el7dLrLALL+c8VE+xFrKqm2eVr6PgB+tpK8LWPNlKuVRGv3XIwqMuvZ0Z
KaoDv/Xr3evnUJQPB6/ttaY94FFSvc3z3sS8/9GlFvFBJ2c8uR0WOxssGoRCRe7z
wPTxDP9ZFRkBDPx9bBVD/lFjEKIkgfKXIfzQrbxabQQA4HdUjqUdudFcLGwYJDww
k0HC/W7KNrkKnRmiKzG0tlovUPfUBVmZJtEy0Q43bh4ntVaa4Rta2Og1SZqDdmTB
oLcROGhnNgUBf+DcmccRndoIarHtgCb8qEpZcZqOKXzTRQi4HlhEU2a8KvVzw0PL
YuiQPVdywCZLvFBMyBHFrXFRZKukQUuQA2+QipiBEppVc7tfRqEXJQmgYdL0MDhY
scHPKrF53QRl4MT/oO9pi2aApMrEpb284Dx2t8xi4lDIgwusAeHfe/YYF1amfEcw
clt9rqgPDuA84CFmbghBxKEvIppp8d03YMMrOcU3Ihv6rxpK3z6X9aBz5bfcH+Ho
S+Tz0uUO1xRj80JYpv44FgQZ/w8pZzjvWr8ykoTwA5pz9goc2lS0P/7YsiBmY/qt
ibg04UrKvaMyil322A+OMncQSJ7iFmD1O7vc4fNOXQf+nRgwzOhYIKpn00BjAuwb
mzYv4ZXZeLGy911rWxI6PRB61pkuGmB7j0t5zBKPdHbd5JN4NmN9Dp/JC1CIOc60
d74G2XEhgIklM8qyCgl/FbRC6iF2bS8y8hJxw0JsqFWeInKvKBSGVqMVhxaYGjRe
2PXzf5Tsl40p4mnOZvRn7OQPyiRWT0S1+hfFIXGtxU9zHdJwwCRA+/Dr1v1L+Cii
eb4UHE+b//Qss1542dYx4D6g3UgWVIxLqnshChvlwKZylii6BVQWky1nmGHfJgul
R+jTSutq/PcE37RBYz0QTgYOYnK8rg+V0QBrb2d5eMu7UdLgdVSC+nmPCvB7WvYY
1GpKFDAURyOccBA6S5wVQA7h+396pvvSVkD7haIyHprkl5vy4qbTr2VsfXbnZdEH
ZjyiM5YSQdlF7ttIGRBDv9LI8a0k5W/xoEZx3DmBq11j2YBNjwdU6nzMx0iWJFQ5
2M0mQYtmhX703p91ugHB5wHGiaj8CK2+0IGnxVekZmW7suJyHSwEYsaVmHzyQNzt
IelN11+J7SteX/QLlkCygR8cIrBlT0+4ZPW/ffrZkoodZG92wJCPWVIu6tdhuXty
rZ9WlyJ98zLWdK5vEjpLXIz+RsnAzH4DhWL6LzIYjQK+1SC0POuaOUqgu+vlpnmX
3WY1ojhoz4G1gye+wcsHAu06dZVl54I72X3OUtbt74hTTS+1gu3qfNwqUU0/0e+0
doPwb42tFJxWJ/+aEO6V8hltSfggA8Je1kcM7GPjSWujRTtkKAuHTA4i43CPMLE4
PoQtDjBgzrfI5l96o5wessWZxEWNcQ6oHX3Z4TGu1LZWSaa6J1tlaYaczou8S0pi
YgI40nZJ6FVnWtCcUxVQ1Ji7YiR2q3pWdvfTG6Vw+hZlvwnbuuNvYN1sRWkZVsHJ
84y8VZvZ2dCh1fvidVhK6liHVdhP2V6ZR6WTgRjOOTQJZLTCT9uvM6dC1bx4EQuq
VuhjqtIQFrxXhZ3d/3vT/9mm5JupFa5DvCEyFvPhrOjHbBsRl/8teWYZ6p5CV5v6
YK3dBc3DPyB6rUvxh0vVbhZkFbnR6aJbwfjmBKBuTX/MPjN/HZ4gqZAH58N4nfsM
y1lAd4Z9jVNgNJkHdIBkNEVR/hpeR/MooArCF6niaaO3xRGvyqJbGd5HZHD8Lao6
Fx+w+DUK/EUap3JIvGzNbWhC5H8OOzCpWe1GYuousuKo1vIEZ9rVjHhNQhQAGdHd
H1jbigH74mgNvOOGCF/FhPFJdYPqAzIlQ6qrIS5mEQ9tB0/rP16Kh9SJ+MrC2p85
D5kFzdcasssN7+BcCcM7UpG4JDCYIKa7dBfc6wS+IInloDZJdDgZ6HwkHuILKtZj
CdAs7bnrdAzgLL+98w1xgQ1D+b0bmieTN+WCSrcuOFNx8qZyXz3UTO1owTtpM+jV
a39zinpx82PBCrwXwgLAMMbNQgmBnuPLfHBkkQe9JIwMQzNBLvLLYoL0XB54dFjc
KKiexVyibVEVWCk6K+fy6L3gXrq69URvMxQRQZusi3cHgWs/FEGqrQpDaB0N5lWT
9BTT7ptuzK1Gp6hA054Ol9bixOQIdafiOMluOgZEYUCzXO8a8sqVQ+gsNIy3Xx5B
Dv258dcJNAioey2pnB6CkkuTi4tXkaJz44AOQHX+c+uo4UNqUYoVt07st0heOJlz
eIwuNnKY5UWpGT+dlQTu609Tg4EUH/Th87fBo7vd0Yc5YYxdNF1l5FT+vm9B5fEZ
cfqhzufMjyol3oTRtmlK8l3QeW+hfBu+hX+yi51QgOYiak/NmOAeti88uLv8cdVk
LKjVM031S1tetwHdTAL1sao6Q80a3l77faK9flgSVRmB+WrPGXRRyvXSnB/6NTAB
6QZTypP21fHm7fRUtCnBOvFUgA2IPlt63swA22PW/k6C2uZEjTBUXqINoTvvaQoN
61pT5mYyNJumRwaDxj1EDSUwdGAD+GmucxQAAKM0EEgZBOacKH9zLcigMArY60rC
3Nqe/eyQN1usfibVwaICzEy3qsU9gbKWFVQkQ7jyBVQx2EXeOt69DatAyoBvBZQa
ZsQQ+tGee9onV2lsMqGbqfl5ZgBA0T3Yy9z1Sc6G80qyqP1RkMN6b2aeA6V2ybJq
uUIwTPzlmqAjrLfVCm71AWC9awp2yUUjkM48XWE1to5bbl4smMPvGYzGN5f4isiL
r/tqjUlu5VvWNEGczpMIAX6869vVAqCyL2+E4jToY4/H/DdMhp4jCZbRjbQ3Vq4R
V1/FLhyz2Rwp8loljeTtHiDuHHrLOEt545e7q7IT/c8jOJ0ENef9o1+vUsj4Lvnm
cdmF62wkq30PIMDKqj4DE67jE4w3DRmsPeWcgdkLhVu6guptod4ZCyOopDYBLd9G
HYhQ/bLSjiJ9zqu4vku0jFeVpuIrIRDWOefSempMyuiFWgrZY02qIwbNevwI2hMJ
750XOm5sRSukZENLPjXB/gQd8aoIo6mWgf1lK8hlTbJOG1JhUNA12q/oLR5MbZAD
9sdIw9w0eXoDp1bR16nYhy+LRS+6qukIuk7tHYmNJB+69+vaWwTbEg0cLPE57Kr3
fzogNuWoUaYIeQupWPItfxyp5PG9rtSb2aVkVHzxHErat12w/KbXf88gFDLu6imk
mzxBq2131KXtLEOIEcOipXMCperOigXrSndoCPGaoTr3talRgg7vHVLwdyzbggRm
C3Iydh4Tvnh9zU2Il+zWPFfNMNKOufP6fvVuYH9bXxoDPMW0jdCbBd+YixthVoyU
PzIaAYPU1YSQdw+dd8MvPq9nYcLJLRUcFsRWMAeFrkYIXV544FtWiFT1ARUdTBNz
ZQoE32CCnZLEorbsHMvSZjW0hcBNtgEcg9FTOhOYJEjY/mUGcTa9y8qKKGlbmLO0
585oFqWbDxfoIN2blZEm4OYWRdn+ToKS/oyIYrrlMf5WJ1LTH/aT3D67e2icTaU0
ygi1GowvQLsb3b32aA6LjfYJYHe4P8s7KCxTHKv2L3JHaF4XkPeUZFuWX8QHVEqK
iVflGNNhqJxPaULuI+K/FWj6Jv0VtpRMSijoHZpEEeKb4fpkfvz9wQhcFFhMCABQ
SCeu4RpMe/f+AS2REZOxdCNZ8xtjKv/Jrjrt/6qZF7KEonSE+Sls7Ioe/BEAm5Y2
RC871l8dycuHL2Q4Flu9XEsHDYSo1g/7o5r1yhEyr9MD6bPh+pYsJyAiKNxUVUjf
Ku6TJtmNr8h1pDmEYfEQoGg1s4XX1ga9XNOE7gdrh+aBqbYoc6R5mzCZcsaNuxJR
SbRn8eHpMGQygUzfrrvcGIM4/dhfwGScXUFHbrjT/r1sHgYJdrYfW8dv+hOGU29Z
8mGCViSCTbHwujXxWNy/UeZjdrWjKN9ee91EyoKJ9WGX0j+49UXS6QGShFG0KB0m
F5BR4s6JUD11QcvUBZGtVj6hEZxhlchxxD+AW+TqZ9Tlyjd7TeQ3l2D/c6R3sFEp
1wW0+wS5xBriPVCObwMiZ9MagFCkgOG321mWIJBqIo+E4Dm+YYFKrCujQAUtfqyG
XM5JknQfl+yXEg5x29qHR/JFRZuB0dW7cUKHXhucYnpv7IEOLgZ9/uj5sJ9wiyBD
YtnYTpp/sqoyHIofM57Kh3HrROhiv8SxqYkfvny65ETrLL3fjSRFaVuDuo+Sr/kc
UbuSgbFki1r/rWjMenYyIE6+poaUVEVLnRyDertQSo0mimfzhWEKL155Ew1YMu8l
UNPJKtaEJ+JEEtBX+UggpRTfeujBaq0FqDgZxbirbhb98uEbfhF9Wt8oQq4sWnAu
DRRfVTYIwxrgN9rUpFIv73c/La6+GBvEp3iPgARrsWQdccFXS+0/xf8E4MD7ocxV
HRqpCA86MbpmOWkfqC3g0hBrcaQpJrk35KnEyDE0ZSGftuwx8elIif8M8E/Q1Gr1
SQ8zBWqShylQeT9y6VDmnsEwrwXqYv233xFBP2N5gK+uQO0+6Pezth/EofjqS+QD
idJ8uoIgeAy8oOH7VyO67k4Ru978hHhASeQYBcjdiDeCT9mFeaacJPCPkvyNSVbK
p+3Eq+p+4Q5K43DxRKtD9CLavniMpTZigSGm+yrmx5o9amclwvAD1I+yO7NGVJA7
Mqk1wzj5WiDot7kovCrSnal1UTvm5SP0a/TkLvsl0OaFNI4esAgbvyH2uQkNseZz
IuTCi1FjGWOqTiVEfRN+5fwTakHLmOwJIJO9PFBNujnCs46DED1ITSHoisotvqCf
YXmgqakr2L/vchJDMlSMfue0xLV9NQncmzFvkhsAjBsjmPcBlCp6ZTDhjPTxpW4v
5/5nPaBl1ooEjznzv+2d/MTlZNtgp3iwi2EAWzaMjH77RZOV9NvNiJD/GLPvhQuj
WrI/PLHhod2scGBVSv/ba89Azj8Ga4hzDdAemZynumuSgTiEqEaBSu/f1ZA+yx2j
nSE2uWyGmtCEZ39gRcu5zRBoW2NjGSPJHCaKzXDr5F4J+ECkF/gspZKkrfH7uWAJ
07Dn7/0QXmZzvcxqnNo9hCi4KNL9BWMrowIyedqQD2sFJg43+Ivp7KqbdNJsTdEt
kGciopsuy2yo7QWOIQaR9y/5/1Kusj0iyQ3QIGFZ22AgN/Kui9oCuFDdPUBucm7a
17XeUsjNpmamVSjOIol9ZUFrJMcydr+7wX5kKRti9/ipmkCeyb+JKbz1Ldd+0w0r
24HwDct68X+ygLPqmHfaZJfRv1Q1mel5m/HvWwVD12nvwO6wtTADxSexWqrcRfP9
17rkVyFoHa3KLxUm5xdtsovhT2aB0Ju6RYCRacZcez8Z34EeIzcKf0+EFk1O38hY
hHb1NCjxQY3SQibINA0ZaNQV22ZgAkcN7f0r0JupHEzxvTst2/u4H9fta9bizY9h
vZ2AbHiXaGwPrICehvy+0RbnaRxE/A6deimYbJhvE1H8rNST2stYCFJZlV9zhsbZ
dUW4gx7/RbNyQ4z3alojDZzXHymy5LsclMW3lLe11o6No0ij2hulK6Z9iM2iSxuS
3SXff3ReFV4uFbctTn5g1ro91eizlBAXWm5hGXqKiIIF+ajtc40mnus+qPQFqOLQ
5CWlOHgcpLtt7041lX7m7kXmV9a77KO+iP6B4MSMUqph4/56bK3TgU4jhyNB5esg
erdZg7SEzScUADOwqaCvELA7+5172HZ5QN+LMoXp+vVijKq9Sh1YcbRr8ChEuX6O
3bmJynTSfPxpAOf7NvmLML3WFFlZmwhhsHTuWffL3XyDXCt6On0BuG7irnDr5jZr
wvLM08b9WBEf4a7hs0zX3QJ8CHOv+WaAQUJ2zVPkcmr9tzcciltGWKMOUFK7AINe
PZpRj17C0gNr9LvbBMjYikeKDL90mqMGpk+fU0C2pVbh05FmSpOgH1EqXLAnlJS9
ghEpKCmEOCPW5Vj2xzCHF5aN6CHIXRSlK6obBNufldxffLxhzD8aK8+xTIge/2j2
OGGrj2thNonXV7ahAncp6iROb0VtqiE9FeXP6BEzvYwBepLUSpdYYF50YKJUJ1wE
EE8Ids3Uqstv68m5tK/6BMITccwPc8aP15/Nj55XMwoBhcafctH0G45S49BMED7U
aIHbiTSjrXK6X/LexaG6Wuk0Aqsfi411+3SYjhuYKnoyf8snpYzUNVDQJD41mJK5
nx2rvAPJ+9U2RaON5beQnVqJKSRyDQgbR8OVHbOhFXYofN9JXVtfYk15mO3ztRTq
FdogJc3YmYASbl8hOcSKFnvqEoNomn62bg1ZcslWErHCLaGUFVRg6uv6NyFLiIAw
rgOUe4CiupTNOueraavewb4q4JD8K/sxN0uEhuVBXl6IbQ3gKX4GJpSbzfsyZhMB
Hgh84JkRA85mH58dHOWSvDiZFGEDy3opGkWtVTU1JtO+Vjk9F1lP3gIugICAo3OZ
ty4XCqc1C19mLTkZgt2tj2zj71RvJh7kvz8QzVnsHTsBl8q0kBKEWeV0XfMyGsKP
K2F98M73VW2u/SKbNt8fuBpSkfQn8iS/0MDYOJkxRujo/XgdYaqHCAIxQf4vwo1k
j7+iijW1t/tDhBrMbwhjolV5+7aegALN1l9HeNP6ofUepytWTQw1tBCp8JDA16/c
bfZKQHjx6AvfHmngw5Ajvhda9EdguBDdWVDUbclDO1N5snc5Sqf6zxgvZrCJzMVT
OMMPlJFdbSshH7yB+uJT97FlpMHtfTw+i/c/i77DxWp3Uvqy3e1PgE+b72bpaF4G
G3ICwU5U1U4Dg1OBV2OcZN9Z6Q9d0bGfWrMXWSrvRiUNEPivmTFYBL4CW8D07rE6
fWzqZ8p7oukWc3sU47IIQS2V3plAChNZhYZ495UTA1CeMe1hX/DIXchhUFTfOm6c
bkbzfeY0h298+P4jkWiVpasaR16HbpwpMvwldpsGgX0a4GEltTLupjWv3x5KdHux
wCppEaYLwZzpL+KCxxidpWBk7vTo8DN3IL2Zr4Usyratw/XNP3WOiA1ivpiUSzK9
JbwS5Kzpz1uc4MLdDfZahkxAaaQgIU3P1gjNUTI7/eTBEteaNElCvLMXFxrdcS+V
9EbaocA8C2dH0+Y4c0XlgZ/qEdLQe753L5ri+/giYgoYN5W8cGUDrWDP3GqUQ0bH
eaVQ1Y9Rf+/FKCP+Q3T8xpBt4sMOqabXB3SxIQcyd7pt97sWtP/oYvkhPzFff0pL
dipeVpftY/VIsmBQAsaHgHdKyw4jsJqETj3sPMcCOY5KNDvBHcAPrzgY0yajqggM
ST7APLGNF15wg2SUB3rCjalsKNW6kcxtbYY/Miwb0TdhyMtIQFxBv39jp4LmZBmc
JVECZcqlFKzGbGS7YOFZ05ddf41Lou5AIkCwJfNJI4wZ2B7jF7RRSy4nJB1v/6Cm
C6ZMnX8EyhmvpcRSPktIS3jAustrBwk01b1rxoxPT2sMMPF+jxJswD3WYsEPCd4K
mKxY0ItQ0SOMhO/H69JS8nRrnmpGYVBNS2aT85GqfKBqMujMHbiqn4Z/KKtHQX+Z
nGqB/bW6A/ik3s/OyqeBfHgSxsO9foBOMAC3IfNUJpykBF51Am6tEkzsJo6XTrwN
3gw7UPh59MlcdNwZBgWVqjW/NsqzZcfzkj4nuIEJ46Qm44NKmvQwjMxtS5D+D9/a
52U4WZK7NuCHApcL808hrQQ1KmjLG+HV4t11eI9437kbONFkjq4AqRIc6yNd+Uc6
m9RRiZyVdzvJEfaN0AF9ztM6HeXm0RYzQWofdqEKqPawTQeWXxJYJjiiU7t7Fkrb
qJXqOP8gnaS4cWGp0KYTceRAMIeOQSLpIEBFqJgv7Xs15zSZe2qCmdE3n4PIiLHI
7WaU3ragEsRvT7EHic2ryZvA8Az7Spd8SAP2oaHRI1k9RCSeAeVTOtXjgbA416aF
VV4shgdZzppXwCKBpC0P4HMczwd8aAtXeDB3Q1J8Q32A+qnozECUM2K+6uPSzOIp
3yknApg9yIYQ4Dh1Vo7f4dEHHhwAN4LIq0eaS+7VXr2d9EtKRWET0S/ivytrw0f8
PFP5Y2xDLMGJ40lfQIq1naJ5xsGoghNdEdONBL2PYWuZ5xZhBBqy30kCRm4SqJVI
47Idfc85UUcYnh79OnI+XmktRq1M/kmwRdBYEAHG4W90dv+Cw9monhpTRTGxaKde
VVyoZ3brbtcmKus7OLSVuA==
`protect END_PROTECTED
