`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UKtsuzSEhkRypSCwIZOXT2pCA+WUi25KTh2ZVJk5aVogBMiTCmbpS7zVW4Kj2wyP
bTddaXms9yYnZqREzKfcv06eurhgJkZwf5ntI001sSgxCYV3rIE1ILAXlOEshjq2
IcM7/3j5y4mqO2YVKs/5dVpZw6fCh6hKEFk9HdgCB1jblzhCGe3mg2cM+5cO/XEL
UjuqqIUwoNEXzXA10EDhh243t2D+44IlombaVvrfZ/XJ+MT/g/ysegvN6GTEv8Xz
`protect END_PROTECTED
