`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gtf29nrGArlF/MqxHovJKZLTGl6F9C8cloSIFQgh7SYWkzOsS0il+x/0eewgbCKG
U0fbmuxtY3sg5Sh6KpYFf2N9dN4nZqppkWRa1P+YANJ7TSz1rzFgk9F0lktcPwVq
OpHsFni9M79VW6QuFflUXj0smvo2u4s2ukPLc340wQEu/tcaZlRuUnuiC/aL8Nsx
8aircHMvtM3wUcNLtvNTu60OlYftV4ua+QAVrXpJsMRR58efWGCZOLfO0gpYBrLC
FXV5VEPWxVSz4MO2KO/SW61z1aCIqCvtCA3//J2vAeu9M2qBnjxJGwLgvubcLYkb
1J+1R66JA1ymzuP+6Sb/Hlo/mDBWJ8cbdysrJZpFXtQa83ru86z6byNDnSNGwgbz
4HHBAugzh0H9SIAt6UAGd3SoUVA5Ctpe1YUsyNZcJckWxr8ENN1FyoANTiDGkrtn
0knDpiAKlsrxuA2EcwDXDeNagyz5n4hCbyLns4pvsdO7uOgitMPBulUR5jmIbHPI
ua4nOPaw5MNkHiy6jv2upY+Lry8U73Zl5mnn/jQ5q8xFp+5CclzdsBlYNI0d2K4W
BjSVWiba5xR3RzdvhfCS6AAHdyvMBJTlzijJvGL92hfnu3mYseOu/b5T/l58rac0
5Qe9xYVPIJXHY59PSs7jY0oK2kWrFJ8HsxVc77M0bwXlM7+hRPN+TmHCTrACLfOx
ipIowrl6l/yyoY2VNm4mbEO+ZDg2Boolla64D/1N++5nCfcpYgNQqkQLZsjhllsG
`protect END_PROTECTED
