`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8FJp8MOfiSTUw1VjjfbBJvRm0NPEsERuI3tD+kMMio85S/iVU4Lu4bv39au3J4Le
Hxp1/hJhN8CEZWaVLxOxxzTAqVcO31L7xSz9aimFlj1b65nxTMTB+OBNkHYbZDes
s7NlcpmOYopayd4lm52PulACnUFLD18mniFTsap/YpvmgXa8/XDBMsX9HrtfU5KG
pcePZ/OwqjgyBNwRBczJBiW4dMw91a46h7+BLqCV0tnrE9QmL3nBSvqfsOCRgUm1
AZn9VCJs9phrqcMg3ys927n9CqOPQQh39Z4Munub6S3PMj7ZhN6DQKX5A8Yq8WAd
wFQbgRJ7UGUAUpfzXWEMvRU0/dt3IkqIr27izXnNWPEq6ywJVg0LGvC+CCl2qkPu
pkcyst2opsAHA8exDDVXZg==
`protect END_PROTECTED
