`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uT9sECf/tLES5Gl71fVn3BrTQhuo+lHME6bdEZjLtUgbYnjERfnJsd4kboTEMyhE
t7lwBCgEfxNyfGx9EceLk5FOQxbpqMaFu4XFRIdI2OB9YQ3KDWB0IcGepEwN0+FC
mAj/RLqLKP4mctbQQDBXk97NkIxx0J6rprDRA18P/375Lf0kVnpTVBGBI50lhB47
i1TsrhDrz/Wl4nw2VeBspLZgvUIeNTr9yTtoAdalFMR0Wgc41tE5NzeMBYhhbC/0
T5BmTI2OBl/I9mEjM8Wm/mmVbf71cxVvz5ZJUWRXcJ4eoLA22ZicJ6h9mguXuWMh
m2t6w29YEBZATj+/9eWKE+EadnzwyKgWIbbv9PH0XCixklJDdP1ZjEjJ7KuMQd1v
yCdV99/DzqCc9WvJcRd77RO7VCqO0rg84eqSYsD9MTBLkhM0QSU3jPy+DDCD3D/s
HYE8kzDW9xW+SZhVeyXbJfQWv4g5QcM3CkKuoGZs2jJfdEHCroMAEbJtax0HePG0
w98JVOXeKPwKYtSzdptFRDrrokiN5qczSCfAGjMTKbs+6/8+BN/QRT/nL6EfmltT
Dty+ac0LLGeM/We97rJhX7LdNsk6om3WySJKXCPCOa5b6Y1gj4tJ6PlIHtmMt9+U
sxhd7iEuJBpdpXErj4nPoYAWyYjeQbyKhVd8Ute+DthhkyqqrZcpUU+rORwtlURA
f0UyDtYawtwYtgNW+DFWG4GVaS+8kqwcJ8Tav8B3LNodbhohSRhF0902vE05c/4Y
Iubb47136td7MIJKqOxnhfO66N9Mzx2ZacJ5dbU1DlfVdstBLmdAA9CxOR+qpop1
2v7dEwSgS+UWmFgKfq9svDIfcyBQGTpwTMIxJBbu5Zungv7kWieIkwj9kAxEf3Dh
Vs89rkmZYRchrOuvxQxYeGMpBLU078rtSwoQYIllhr6gnlifiyBFGzUuac8xPoZe
fh8wUK7N+1w76fN4k+1kXGOA5gD4b3NTIbnlccgaKrNHmFX49KdkTp1uBRBbDSTz
`protect END_PROTECTED
