`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F3F7hR7F3plmsxg7RYbpcfoJtUA7aFVsxoo/HDNSMeOBxPOBHuSuwR2TT6Ax9DBt
wm3+gz8oipE7SLlecu/mwlNLRQlcz1DUTQiTr5DhqHcIOCY5+Y37MKiLAymbfeLx
vP7My/8JxK61Otz6T00dg5AJkYKmsDxOp4+V7Cnw0YoIH9cJe/I+kQ4W4x+HVPdl
RgGrduG+OPRg2vbXK4Hys3GAOctGv+qXeA7KNV15eV20HeVAKq2N5odDtyDkoOV9
7wxHLLP1d30STz3o7hrlrl8GX4F5U2GnhnfXBRoterKCuQJ8sEs8SwWW+PPNrbQi
xfSGwvazliJmKkBq7szAqemC1uVfLVeOxVPaxbXSi4dnx0jWPLGPwsXZ4lzCpDkN
OtQHOaA0gLk0YrG194+t4SQHZDoEteskQKHRRarz1kZKlShOzLQTRgfphj/dwrcu
KGT8hSlb7VtoP1MSnX9VC7HzSCsoR0nXXE/9delTLB/b3bFmv1ctMj4aQPElEWf3
vrAo++ZcM10LPpX/Sb+9ndzr4pjVrVN+l770vf/4JwcKTzvu+ChDWwFAzkZ8nshg
XuHrSrQLQv6J8p227QjDWqTGdrW0PLLhw4EcF2FUkaD8MZClHhYKcsuJ90S5l9O6
7VRIEKb3Ev2+XE/qJgajUIHmtqqBDISpLGT8BwKQitVKq04QAGtda+8iSPZKFrLJ
Xg+u8MsS9XTnR8w+/GoGuQ9HJ9vmnv+WFvT+QPnCl3+4LmQiegRyxmR6s7SgAJOh
TutJ68dEQnWquNNThQcRG4uYXsVwqr2FUmIV8aIJxnOKhzc4G5rKZjLs8qBgRBnh
45UN7684nXlxkLKYq0pp4YNFtWOAiWOmsiynMSh1aBTvHLwyJnXYPknIrNJ3G/Iv
`protect END_PROTECTED
