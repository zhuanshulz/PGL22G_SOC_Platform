`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IotXYEKnGRq3JBa97KAJJyqTZs39ezuZR7P/Dg9gSD2j16SUz10TVX3YgMWr7ed4
O27THQftrxmgb0kJE6JhWT4yrqoZSCbe4pSYpYranf5OmYSR7fLCS8jp9vPzZBc0
ETcEqcDsiU37Z/u7cPISJ8MHRF0xOejkyCzXbN68/QZGfbefBBArKjprIy9U9mPa
hOOQUko3cR3y8cGriDGBpMLzUH+0cwp8jrOOgkQcFd+5WhSv9ue7moVnCmQZrgVU
1uA6HKgx58D/PBFlfKU6vgYDTi71+hWlBOi/vA7UEJuKxh4rVmNn82KrBc5CQpQz
JXmbFRVSViayBQl/SNfL8vcOTe22Ml/nqCE0q80s6lGUqlxV4rkTSYOGNB6XXUZb
G67tFcVBEA51UBdNWmMM2GMs1V+eV7k9NaZgWth78T9PxuAphoaJ2YnCsezNw41s
nxsPjojgwZt/M/RiF3Hw8goGdxnFddVTEqhI0gfqqa2ArAXGNNhLsqJTokLADisq
sGhfD0nKoYkK/8wONFy1EI1J3/HOLbiNVFdRidH6/+lrsQ59kyWIbPLobM/+h9z7
9uicnb+EoCQtDfcG+c8hM1N12A4X3VmpYhrkt1SdLh4qBEo0HZmD3diB5rLvFuLk
zJN9RRMx2J1wwVcv09rhDKOCm4JPTer1W/qLZy3S9oe58Gjyek2c0KRaVA34/g4p
MgJ6YBOJKWUWjmoG3dl5vnHSbR/P/DM/pc6ax3cAVsplHCXmXV5JKwr5WRnKBQoj
0YT4VIUUUQkY+GqB/VfXzdGFJTu6oiTS2GjxXGOv62Lfa6b0ZrAEflEIXqEJI5/S
Fs6NUZSQQV6tJdccBNEqoJYJhwT6SMkS7qgnN9Kqm8vahMzxIRGDmoDFZ0U9lGNb
JKJNel81YVTEwKirNtivaQbGNTdHaHMzxBlmVigRJvc=
`protect END_PROTECTED
