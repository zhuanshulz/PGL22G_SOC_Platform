`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WnrTwuTDT1en8GrIpvIjc3q12y6Mr9d8fKZWKYceaY73Te+cuiGYOLAUkdSu6SA6
3e9uNrWxnK9UzvoBcsoK2E+VG7alt8g5ArX+xjOoJy6Z8hN79uuly73UvYRWS+Qx
CudqfetA0W3YXkSiHj6qfICYjETEVUFnrv39zRR9sOqrKEWETy3u11pT2hNAgQr5
HD7w40PaXaMuAKLAgC8VZVKMjB0BKHkzt/9ZjekG2wuCJSEZqmL8+ggCc9ofmbVq
mAGPZkjq0SLw7sO8JBvD0EN+LmOo3o5acEQr73GbbkxbY25KoyfN2LLNZZZbFRfi
xiSlg78kgSEShfaww04Plv+VBRnMc5mWLcIa5/M1fQ72jyGLABSe7lfNaCZGXNlk
40cfcW3Ad2lDUteugt55igzJcYhgdZgTkXUb5Lrq9eos+qVPrNTHZ47nLG+4boX+
MhJSO+Zzdy7UjYdxihlg7t05HqDysNa8N0fhHY/vbd91g5o2C1geFLnbPjjQWDKC
DHHmXsnYrtpdJR6GLKK5+np3NPiWxFFO8WIQbMCRqYYSS57qeEzQ8IL6e0JdrNnh
kqiEv4P6xn9N86r/FZnKtD6Xa/S7a5cLlgca/bFmUWXVjqgHOXxnBdx7Fi/3Q5PE
cWH0agnMO8eGGl+JYrU2/SSjBvJwK9ILXEE98y6GIQhgbFJJyiKtmAjjy3cDHPFq
0EXX/4DaJjxwPpZnVU4gHq75pBEODzFTgdVY61n7LSqWjp20l65D88us/kVEfiEf
bi2tDShkTHbNGmjb6IkB+VV1ahTPv/QYuCudspHCKhj4+eA19x7yUERb17f8khgF
FN0/gTPH1g4rcz1vKNBZSEUfFhuwofEqaWDIMRXTX67MczjSA45UrcCF3kUdVEph
+OP38O4IFW20X220ceevxEFuWdm2tBJX9aT50wxOuhymKF7V4HGd4sfX7kL5XgTp
ExThZTAYCp/vT12Mt2VKoUxuyx62KUYG1VT2t7GF9e4mtOtNNZMGG4uKyj0OqQc2
TQ8LJktpBku1Taj/wPTsGEGJDTism+2RgJle+Ja5eZxOwnnuAgel/1jmUDnO3c65
XIfBeRDqc4EJMNhuPrU0jArFfDBZTVu+r98SnyjNY/8w9KD13CEkp/RkA+JUFoAN
h7M+lavmhEJIYr0QQPTP7W99JzuR8hbUfbz2B2DloQB2vw5er/5cPQI1Z8QSVD96
jyWD2hBNuLZabxuJl0BUZ/CJhD9Ac6Aj8adf4iOPGYYPX7G2WeO0tm9mKwUPC8T6
Woh9YAceYEV/xcxvtmLNlwYbpyxaEG2b+eOaeuzBcfKxxEqi2VARRdK15A7fGyz9
rcmUkQeAQuvaFBDb0aYXiHx83P1fP/FKwMhHUTgRdWlhfqG+yXinaNLwQRLS1wSb
BpFTnAdrB8TA5+SyjeGYD2NAcYP7JzPzwFZHvMHWIkOV9p3NtNWXGxYkP3PCQj5s
BwZrO7KvOAWE2uwFfooskzb9/5AEdLyFfzd7YEmD6lvKVxyx7is21lhRm3OCzo7f
Boow0ZUz0JZ9rhiQWbPMe8BOPoDK/3EiwcBt6ja4g/68fO5NllYc0eiGpZBfs/h4
AQuMHhTE2DZ0nYXP8wit2iDs/Ur9CLAJRI9cjS/LxL6Sdby6TMpIEu6Kcmh7aXbi
e5eKMh2rUS0/P8g8O8F0RYS1IGqW3NDF9Uer+IX1meS1LSr/H6/yj6i5sDCD+txB
6CRb2K6vTbZPhhhNg7DeGwH9EhW3Dje+4hpPM+eKRimU/6QZmHHvYrNhyOUE6kI/
hChfeMbNBcKB2AJoBaOjpGKE+HdPyC5BB6gDvt+hvfHxtn7o/YH1KGD3ejaqazZw
DTIF/Bs4/qb4ssZgaKIvsu9yBjE4GF2I96XVTc0v1dduJ39YXS4XFLrP1aVUTtf8
/BROv7AsdxYy2XTeQLLlUDRsVMAMlIfg0fq48byn0qrJZH677P7HXWu/9B+4bdKL
gJJbpDz9V9+Cmd/kPKVTw+XMiQ9cx6cpK/EgZ2wwMwFnUpGgCvKzSqbc42/GxOBs
D/k0eafDAO0kVslsvM+qewfgsnpigUnH04MnWfn/fvGSXXrjCBG+PfK39VT9qqQ9
LJF75DbafPj2wazXfkQPC4IRI9DxDku3+6m6o8Oil3N9vLE/PjaEpmXJxvmemX7X
YvWhI6z88KOIfgpKvQU9zgsEAA8g6hlwLLX6K5ZCAisTdnq43Xt2dsuSaJb4zDWg
PSzasa8hfcCGJmZKVddzO4N6BzlFVFFtjjRsBGi6ExG3yWxyooq69zCR90B4Ovx6
L2QZ7IAaroZoZQGOBzuINAvqg4WqJ15U7zYcbgFv93u1y7Wh3w3T8HVYpy2qMjTn
xnlvpyXFEfuzjGZod059Lq8RW7ehHKPr0x/RuA5jZUrtXJogmAVt7QQvM1kTQtm2
svMiC7D1dsV9DVt7G4Q4M9c6o8XL6IcMIpXNU+qXDTIn/ZeF+2RlBBRJhZRmepLU
kHD4XTU77PcLekyOvn82yEartj6jYplOM/5cMyjK5lVG/noVmqkkabcEvRAL7k+Y
zM7HoOhS6ckoS2D5QbJHIk5+byt+vzgmmahpSF5++J2HaKjRiKuoMGEYct0DgG+z
rbBKXnjNbfNgbq+SJWdhM/VQnXRYmCzq8vVzB7ttae4wVJpAvIbVW4jNety2jARd
Ww++pCf0Y9Sek/udlgiOvylYsWfuyCQxLC7AAWAK7tZmDSSp9yflfEyJ6DeD3dmD
55E3CMaKzImGdsbj2DdEw3EJ4/8J96xQRacfZr92v9Onk9OAa2S43F8SqrJXPVlB
Q8aZjoG9ZEimw1ZygF3eeBNAU49nGmKBzMVMHosfv31OGRZawvAcTuKTuW++NNyE
RvNEpuwnWfggU8oJKRbX6636zF/TFpho/z5QCjbxxqypAEwY1lPd5I2xXvelm8RI
vLH3pDYumN85/vWQZgh5MJXRHLgAED0m37W53Vn08BsqaTHMkIx4ijKHJeYXk97m
dSvS6oPqUUQZmKLQdRMdEn8wtEVy9nyZsxfAf+eACWrsbUsBNs2BLRAMRTN5p8y1
0VjtIJM1R0ahfchxasYT4DJEZp+AHeRGjbFvIBqQJyYwescEytHWZZJH0xRb0wey
fMzozdi8X0BkTq3gACtXe4PcsRrOhwfUFtIm7LHi4Fj7NFNM/PdhOooPMbX1o5DD
vqS7nH3DXAShszC5hbOVJ8X3vx29X+cPIHdSMF+lz9A/okUkws7bNqb1GtFBBOOU
i3aEk6fr2I7Pw4JcoU5NV4zbjb5EiQGAkyzINsG+mAiqHYNT9z0+K5NvwODa8pDE
Da6vydC0k1qfykwxo3pPnEyMaFas7ESphwmMJxNnUGAtZgOAkKIRKB2xbNOlboR8
L7D91C9RdaujKVfPZdgnkidrFxqKx6P6lV0T6Z/tYtDrzmuERrnKUlwuhnuq6Drf
3SafSVAYF116ehX7rQhQQx5qirA8RB6vXV4UdXC92fF9Y6q0wSnEOibL9lgLBvg3
fZitKERWWRExf7ed5bnpPUFT1xi5NnogPiogI+gz7Y5Wt0kJ89ZWUCwMYKLV3gI+
662ToiXuQ7eoBMVS6gZfUcubTJbbPcKtisLYmo12tfxS4B4qdq4gSFBG9vulPIzz
Qb7DTwnfsE4Cw36uwVUkG+TjclxzBTmqXiUUCoCHWq07PWJBDwoUKzLA/1cWksqw
9/e4TaX2Pndcboz57bKHH5mj7gVNECz7vbWlKjmyYhExogGTc/5Pom8OLeJYPMMH
aYemm5EP/jLXuU/FEeDrpVaJbJz6jjQXl0qIx4mcogkYLc05up0szivrQWb3S5M0
ZBnbkx3l5bTRF45PMLg2Med9C3MlEhEHEGIRyWlaIQm2Wx7ItFbH4996MN6/Vs2a
KKIeBaeBYGwkfMTFmlY36WMMhme+L9cDFuk0Dsmt3XRGs2AMa1dGy4CcqtzZThYG
2Ce//UA4jjijm5TQv5eh2nieGeoMOPNF/0yCyMLBXw9avfClKVN4xgGpUJN6C1sV
6YoNUN8pQGYRt5RVINcsfOCB53Om1zqF32CYVXpVnYDR+bnSjlaS9cy6ommEb9zZ
/Sj8G7P41GHeiRX6MHoRchdebL5s9wwJ7fEUuvWFqNdo99ub4gqjCOs+fyQcKbhZ
SsOAGMdzaRjt7gEdALYGJIdR+p02MqNJRn34Lsp472S/vF1bglyOwrvYdZ6O1bL0
N5j6Xggu5h0jbJXYfePwcwfoDukqH5Nd4zMfj3uFjFAXZ6T1HweSG+YZV2tZccgi
GzJiyJQTmVXz/ld3BD7H0wcyag/DoBI6o8+HsOAXAveoJ47qtdrhVRZpVKKKxGKE
XJYyMBVwTUnDc189xNdpEnQHyPMagsPaqjn5UxR8/8z6LmM2nkL5p/KXM+08Cscu
SxIPN6bQAtSt3wx4VmJcESSrOQfWXeWhYcgIquRj0X3oxLrbQ/HC6OBS6+Ypst3i
nkfXH0gQxs37+uBwf0UxdxFOHFC23wbQMrE/V/Zf021PmX9POylaq7UNmQzOc145
ZmHQaRMiNvRFXOAMGPjs9P71d+VjVN1/DsjcYC0uzx62JBZ8xAqhzgflPiA06Tyh
L1oYjjhR86HRFlKLj5NKVeu02tNW/+VGpGe0uRXS6E+4ajc6q1TxD4UVNWbkqCtU
JU6GU5QH57NCgNW0ACFOw6lxFd4FDm8e03r4cfAKWU7eSiHAnBAinjt8dOf8rcnb
I5gpJFSDYVfcNT3oarWMcmBj+/vaM8N3ridScvxyK4pVnsNIxZzNkqTWzoaY7Qu+
nTZGauZrRR39qTxEc3chIRigeWuGZtBnjE7iNFOdSXaPzSMXM0oLQiRfpcu/ynGZ
NPZRg+9/MMuP8fWVPGDaiSJbkFDsAHv1zjY9Fpn5dJ2DkaO56/l78nrP2Iqa+Fl9
ZtqqA2ef4guZZnsT/hBqJWY6K8KQErI4febnOfLdwV0vkjPXZRSLHl+pithrNr1d
Fn6lhJ4ZHUcnqoU/Waxyokv3D1gD90NnDWngeZSyvDEu9I41DdFibnrfX7wrmg2X
mPDTA7BuQ+cHxcysi7Mq0E5/6GY8ZvP2rIyq03kWlbQt4eRhnAiLqVp0re4LDMJj
XvN4I1BzwwJvTNQXRQq1fTiilzFw+r1jk1b3RxcyU3bg7C8P0bTNkNSgh7vIQVne
LxemizC9962IFOPSNThwnQXYa+LqPLFrWHH0m1kFi3Dwrvarhy44bjE+y0SnwtQa
D4Ccff2QNlApGXM5p6e5X7vp7dmlqpoYmAxdNXYSatMMzuujuw3Tce8lZ6I+aSvA
0FMl0wMmTtZ9BKb2Ssp4W68h9rj4HjnC9e/9iZjdinPkz/+JBs/cDOkGMn8YxOeg
rXXumALL4rn/tM6w9tdQmClBNB5+S3fV0ZIhomFEpbjxCJ5d6aoLWNzhIlfkSVqc
B83yf+JmO62H5HSDDsJzTvkNkfMWQSCiN+GaI9SPqArm68WOi9KPSxwJHYCQOYI9
81D0AXtpJRlFIFeVXg/1KMZuRIp48yud24ay9XoJzhv4R0DQ9t4rCZuXgCiaBLSq
FDspidk6Dl4mfWdSMZ/4I21lJFLw7fKU6Mu0Lb16b1Q+4Ue9WkJLTnfyDNyEplSD
49jcB+ALRhDdFP0shAn1vDXn+Ur3hA/t3jD84HGnAAqY00Ny1VIWkVRFGfNKgvjW
RFof03KnVkQBtvExKKehAj3LgHEAdnswoqQKp6xwzW1VBGO9PCxClY7EqqBz2bcM
4Q+p5L2YeHglxel8kPVrnuiZvEx+WtLS0iGhUy0meamj8J/Yt+jliwqKMiX9njPp
ChJbdCPw0Fk08cuWcd8N1LB9xEPtvDpyVBaxKjnOshYlBrijeUeYKDT1smnTDUVm
zp3mF/PG1SvxOO+Xh9NFB6nXjZl8MbLCzMvAfFzysBaxtvM9jLm4Wl1977xleZB2
4I9dVi4rnKHEUkwrxOfO3Eo+fBDYOIz+4Amcv9BtS18O5ReswBvi3xoCT/AKMMPR
jfdC6JDO8G4DTuNrBTLiZENoB0124XGDtkRs/UQg6ofQyB6A71KJoJuzgDZMRWBN
aF15XzfLilh5SQcU3lXjtmE7yEsPrB516xC6jOU0IufEzJO80v4gfSFy+BDhnGYn
P7Rad2Rdg/25dWMv6mWQkbkx4wS/3Jba+fXYkO5KNxUjqHJcd5JSBkVt77hMm7TG
wlKAsASbSMRELHW1kLrC3nD6ydZerb8z/qSA1JTprmOHM2jHGX+LUK9AuS7308I3
GzjNe9Z9oZnCXMas++xIdB5bljqiDniUMIG/q1PFP0BOmtqz8K1aldEf6sw4jUp2
ZSp4zX2ZtVwy5eFQu7OzhgfgIcKfzKX48efeVjZsREnvZ58NaYi7lB5q9i4wRi7G
HVC1jBFOwY8aV8DV7ZlpN40oBuX0fFUFZIVF6w9QDdgh/Nd023R+SQxXMGtRmJ1E
DwRlYz87ARUIFlUrHpwHocj1gvcNJPHNx/ZGauQsMhOnkhehvwvPwLBu1i3ltWAi
xLdD1djBzRucBM/8VC8uC7Cy6HT/PZqEZNugUhuxj+mm+ypz4cQQ87THuUpj9JE+
Y/+h2ktB2XVjbCvcnc8KiJsNRawLAfl/hsnDiuLLFWkMOjbt5lFRUtPiAmAzEsdr
KWKWbUL2CzdomWGYTtZq73y1jFJxbjh6xl9cNLrq9A+MnnNO/ECViXQiif1Fs7F6
RE+v7XOVdu6oJKrAwTBdtMcP5O6OGR/jZS6XIHKBbOxaTHBjxXXvpfVQIHbgpbjq
YHQ3jDQouAVwgmX3aqGWUAVoC6AMJB0X/fxDyqI2j+wXSzspk5oLI+A3FNgJ04xF
BQXScqrst47hSFdDZg92QbGkKT5ZPE/9wznoKIqF78K/APtO/FEyMDJ4zdUEJ89t
ibl7o/QVCX/ZJZQK9doD9h61/gAAfgl6ZKunTQVlSeQiS8hSRN2Dvrm919YzD8C/
EQhvzoIgV0kKLHcxW3z+zI14ctXbJV1cvftHih7kzZRTXx4+bVkC5BNWFjSSQ3Uh
vnDzipnV86AUidofihvqWhU7CgVpl+nokvFisXPMI5lCy7yNDL8Nli859pqwA42J
mrZWHB0YAnbyxXBuaZyQ88LiBng97bczYuAiyHs3wY9ShYPGT4a+Vn+9sC/DvQLH
xvgq8aQL6tsmj7bA6cZJd6yxJieT3omazZgPBWdt4VGocVFCuyt6GRxiP/tWtQIK
2AO0ccXDxH0e99hmm/tIFmQeiKwqt4RDarRSC4J598hp6z/mzkDBL6QxL5KvEdGK
8Fb7NaF4eTIGuoO0wIeXsO/rSpITCFxrt92dkEZfLefRnFrw2tGYhlCcpr4Qs3si
aD+2bRQN3l2TNCTULctYh0DZPJtHq2+VJeRGH3IIeRPHS1AxXYDXwVkusG7DqCBr
E5YF5GXWJeelaSzyW/IclIqc2hLW4maUZwkah2XkIAzvBe0HzqrbYbbg8yUb7u4S
M6WPxEQbRqDdGc6Cnul/RJDfwO4yYdgAcbYXUbFF+60HnpE0oxVL8tA30290iund
hk3m06UU6HGjdGDHGwNjVwGap1d6m9In5bxQTQpz67NyDdSaSFT/jbJIvzGTgzxC
dpTyIzmkWEqvrdGmHc0ZJ0OhHRF7eU1oiVl0uJu7144bsFyAXCIexyv/8bYZLzlz
zqZexY+YDQ09RT+JCqezZjj5iwH4tgWNU2ytu4IfQCGbDk6bnlRA7fIWR+GVyp5+
1uF5+kczEokLwD4TXe6e/xLiM8+7DR1Rhbyztvxk2iPP9MqRQcTq6TOXuLJilzHX
xY5/RheI0MlsHmPEAPFhUYEjDRHrEyEbdR4UisRupA3oFukxdn0iGBWmWgXzwXyt
0eIbV2Zgqaq07fwyw3xwLQrFDvFRCe2ZB70xzMBmURCvrYtQdsg3WBN1GG42LDdO
W6NdnP7QuhsHWOuugEH1xpzfu95Ca0Ntn1A82KMAdaEi/WGdh0TNApSI3LRrhBeS
yfvEQouMEs1U688obFWD2uUWfCJSKHTgluU6tA1A9Se1Qp2bYpeoKB5VcidJT5VH
5risy/yfL+lxSB3Do8eQNfp1LEEi2fJQ/dbWD3Uv9vIRMk3/e1bkl7koQOF5EBDy
qTHH4Ufg28ivTsGcZOhg/mx9G2rR9WM4COH+TSv1x+GmwCjup39V4jSVHgnpMeO9
9cy6zmI06rGoQTjzM9G+5GhbukfprXhM4OY5BaWhWQ+NXt2PBltHyKJAiBy01XSs
oo3Z11FpecuD3e6hmMSBb1+3zej4qE4mE9gcV7RyG7ZNG3w1nMUtqtaYwklKBCLj
SKU073nP2BDfIcYv6EPoc0En+pDsvE9HPF/4HTFtY/NsDKbbj64dPoUmo/BfVBlz
vbfM+wRU2CHp4vn79WXW/ke7kgZ+TnaD3csv+09Masc6Q980VrHt74IdBgm/E+vy
7y5iXA/S0ckOkaxkh6l80SA0t/nzDlkuO4DUk69UrasaFwTLgevoVlWOBZv8O/m1
HBwBiZ9J88II58xRBvngj6F0/y3CrFZwJ6NAmenPvC74il5xM2xP6Q0Eryt2VLGP
fn8EZBFhqBf0+5ZrtPuromotU9T5cZwbXXyYE8u0USV25K6ZATXdZhAxG+HAutNw
IpxUXoJ0TrgdPmS4789vVyAOOMiUVzdxBhJN6WhjK1bM7HCSP5w9qDvpgTKBgNSk
JKTdvA/mFPGGOYxmr3RGOF1F+ADsqNMOV9u0zIplGLdaQJ8UX4GmO2sRzf5E3dOl
xwAYYtqsLZJNc4j3sDEfcyFJBIrJWeYwZFew1cSzmnSqEZSEVuCdSeVowQGg9jKC
NRmK1onkk6fGQjLoukERVCPabyZIEQf1u8m7IH5fGGUJ/txgtFkOKhxxt3mjKLqb
AX6fn/eGAE7RPAkwuJ8VAN1+SMm9ZfC/6TaBQclJ++rldmFlzXdrzNGGD+bGSVEE
YxzNPa98xCWKhvGf1mog3kHufSyuGZIV09asluEDF8AW5eLfmElGcuHWF8w0+CBW
v5jocLNq6ZfWPKyfaiTDUfAEEniTnRwKWTbqpimtfnGTfDwLI8c3fgBEeAx5toLR
8E1aEetIGVeM0jIGDesDpn83HrFeXEgD9ffLUyetIk4n+elZoRcGK3NkyiEdvIY/
OsU05OZVlgtodm3NAWqOoRlnsHSbi2hvOkWA1vKSu3cZaX75JsJz4ijRd0Swf3Yy
zZisdCDu+SCgVXYcW0DofMPf92gJ51bql6sgvGTEQobpXBTCzd8O13ZV6I5FTDeZ
ZhlyXQJsr+Li+pUn9fDKBGh8i5Zioo1k4jzH2UveHFmgco3CbFMgtaruDYrTkTTe
ttxi/OeKOkgIxS2aLGS29Hjge2Yh49aM4bJXmw/u77jKStSiTPvKu10flTzKt4tK
Sagjx3KRcxyCwiDGqYpW7CHOojKHBq8/DesDmFZNPan5uYGatMGBMCQipvLspYsZ
F/h1xR7mN+D43sA1LQojGV8wfdlC52aPbWIQv93FOhyp8YkjEljTvGc+yJBL3cve
PrVWZbPA7KQIs+N04TNi16nY/H6V+V7RcXcGrV95k9qGYEm05/kLb7JoeJioSx9V
+IvjzaUYDhOTO5URtlvXMgWHIcZ3zNnwliFUaDa0aY312vt6kxtnYUMZgTyHGxSK
M25+l7uWKVAQXQywmM6opV9Q++eJiyUxhejAol95I5e/m3y6UpyLjrb36ePUUfIw
sy+ZrPyvE/MZtC7mHoPDtrc0CS4JOTBCo0QSDJNjtsTInosgiuhmBBcpISdDLGOd
7fsFNWHb9fTWW5+6i0wb4LfFt2O73ewKwUGmSGiRKFfkgcfCMVZBzgg+ql8xNpsp
rPwbhYhCM8Um6o5Hemd3ND/SPysNyCuxtAtbxPlx4Ns4Kh/T8MpcPzFqnZcNj626
1ZoignawfrgAPwS7TL2YN8OZkapyHwlggOnYLjHWUFvJK4Cxndg9VBmP8fBULEsd
gIKYN+YyC/qyEwgw8Y0HKlAlmeXZV+QGDCkNUwRglnliNI9LmtwJbDlAuwtvLR4S
hCLbAwG7msKY6FqiPWhGoOBmRyvAoiE3PhspoZFaQ8TO8L4J6ng7UU2bpbrTBxBY
01PY+pOuvhqRJA38OgH1jflcdA2xY2ANpLdFuCvHQCddjoPXHj61L+8bEMEehKCt
D5dWKSjI47p7B82kUAtwN2zx6gkKpvuXzFm4kRIkFx1zG9mvnR53moyILMzHrEtC
LMdwubNnd/+whDjrUft1FRi8sRndFzK2XGDbnpzSeeyzV1lJDiid0P35B1/EpXms
qhAxLF0WBeJxaHrzahWDUts5m5MVsmOp8VAKbR5jsl/0dLxVcN46kt9GX4iPkLs/
fcr3x6eOucQnlZ+d65lnrHUJRrJ7P1cBA3m7cfa1c/PYu2ynUUvkIT5NhS8+iJxe
GXHFC1R9O1PQCXHp1JD5XxxCx/jnKgvbA0e4NC+WtQc1Tbt8RTcYXDWbD2jnoEgV
u8YBlmQrM98vgu7P2N5wkJp6VhSOCHUaWwCHsEsLE70HQIeSKgtFPqUDD/s73J7H
x28YxpDNp91lPzhq+MLH0HiwoB5GemxAd409KWan2LMb6LE8eBa4k9UutOGdxl9L
DtnMDrdVriMFFgD+U/lCm+geu61eEIYzHQyMh0ZJZ4Wn8Re2ua8frCt/0sqQxOb2
lXzCY5/Y8j21s+AVX9i8acYbtZwY4OdzsjAm5OlO7fWWneJgk3hEIr+WPf5TNZ6e
u0izq6/PyICte3TbPSRLoqInq9Y96QgChqiZwmpXhgBiIZr9XdIJrUQI/YIM/n44
jD5gtZunKMv0MBrQRbvU0cK5Uxu14GdCLW+X10FgzMegsTrQhf4wyy7QTYoRPixW
ZQ2yLsQkUMm7qkjYCMfOFwe952OqzAw6TAQ+whdavJodY1hrO7u0Yja7SX+36Cv9
1UzoettMSsbV5tiYxZLIYrufXjht+yzpO9BPr8WyWEVm3PEjnZEqVQG/Y/JCcq08
CeCb3ucEhWtCyDw7CjiP/VFnOUP8EL8eWJACRtn5G6kDAka8Q6oSlZL5dXjvAHSG
IIfIb7RwD+pSLGCiR1Xu3EQ0HdxpUCCo7kQ+uelyzq/oPTa5kI1ymVG42VtGkwVp
Hll848MrIKt0tleaMVMsaQZ1gg/i2dtQKEi5IEe0PwHQmmMfD2Apc+W2msnYNHgM
DhupEDsUL9O5HdtOS1Ymh6t2UHkkw4vzJMwP8NRHyHadKdv+v0KvB4d0nkQpGWw6
tZwiTqUdMTZFd5Wc5EZpSYne2iqNeYjHde681CoZJVB0zPtYJJJXgjKww4NTo06P
IJXxAoI9sljYCxtkJLJXNPTzLTmW8zTj39dttvQbfXhAWGBDddUHam/9Ey/XuH1Y
GTCWx+aTlv/lpZgW6NEsuDbpgIzWBLsMe85XQCQG9DGgnO0C4LLDIKhzIog+AB4S
6cGhMMDFBvckP8nNnjb8AJkG2QWW4ijqpbloKDGK183w4WWhvCm/Cklce5nyi6SK
VrUQPXDL91zQJNFNEftM4J3W5SJCgbJLCWWelQwnsXnzIzzdlljYOHnckK5MKna2
ZS82UHMRLi14AX1px4YIl4jrIOBPT2l2jQUjKyIxIggIC6txyJ5y439ZwKiuBSiV
riHWaWzrZBmnKbQeDbb58XkHrZW/lEWtgewUmxiTEn8GgUNeuDVfskoEoScNPqfE
DWVZ4Sx+mORiM9NnLwj1e8Nx3GD3/gKZJqzzLH6eSGF0c+Oitw/3a+Yxts8UopCh
B4YjP9a34cukn9I1rteNF+u8emU3YPijPscbrQb5KlXYHLE4Z7aIPOA7IW69A/Jh
apJwHdNToz+dA3k6nNL0vGsaY1mkhxjaTlNWSDCt4MSmQuq+0Pn7zup+ZcQTDMw8
Z5WC7qPqCJLpruj0+itv/Ae9iltvR+jnWW+gVBnYdGYBtITVUQatsTZnXzexqqfr
PPAEgOO/69w8CXgfFOOCBAOdkPO0nCWCb8rlrygMaIiYdPVaXQBVC9ikFqWMPy9t
+8Oihnez05JBGSHl7Xb34BYCWI5R/pLpqxlI1LOx6BG3dY/fde2I4cIBMGFRiRRG
nSC8i2co5vGGCTVYJJDvVmAxnhiL5yTj4tvrgv2/SB09SpW9r7tDd2Aw14MqqVgj
eTeM0ywt9JdjxmNyfMzc+eOMqfk+hoYuNzH8NpP4AwkzzWJRArP2yx9xQqfyEP5W
eyEiz5R42wFOMOesWLQolp6qFsOO8hKcu7QfQX74lqwGEhEl8QiCVe+t5BzEFNLR
WQE6Fmno95TAugN/JjNjTabo+TQWCjDdqeLy5qJ6Widwv1NRkO5Qs4ygEJXxz9eI
/jT4YRONrjYJ0cOfphqNEgixJ8jlhFIP017HtwffAIAjfGb1mgrx9E12CTnyzlBC
jCnRV0khutG8W4NkLq7tDWymQwcKRMoersRjNmxZUTymn1vFkKQujmmt8zT5NzRU
wEFgDABTFWPgluBIah+l89xrJZtgRGzkZGhIdF7GkguaZMQYp0uEfYMUD0Pgf9gR
D3eEXT+hTJkppT4JQj40yxRyAuvMe8FBs8Ba6n7g6L+IQJqKvYoVkSipj2F/7Nb+
MoZsORs2LfUkIVHo/X7CFAc2uRQulR1w4/jqZbi09uynu81GrhS8nBZqcfPtAFy4
YOy1ziijHx4FrXgHRj1yXq5qmE6ONtZ8OlHqPQWe98qOq+2OLjCeJGrOHe7rKKma
jAL+VGtmffkByahsbRSbw2VC8dMjGbefzGHzYYCw39k4DjdgYETUkUJfF+6kqLa0
jbk2J5UHvVmpsSD5IA2T7t6ZlyM5u2IhltytoDMtE4dRl0KxSOnXv5sOB3HzJwid
6i2252XfQLL733lrqKyDqIYntWsJzChxWvuHHhNn7gZu0MJC1l7Vpp9hCEjq0X9W
feuTewSGZCLuze3F/7VA4WnMdJxVTg7kcUREVqSZI18b5DrQL9/yaznRFlf6y9zQ
ntrymEBPfq5KfbpD9no7bQ/7RxGCPsJoY+ZmYRxv0y8eOOd/ofJ5Uam5YbuEUr7R
ITXfooF6z6shGjm6fqqASF6xH0swxpauCy7OE014cIYRgflq8D/dw0Fe5bE7ahAb
ZrXCeipiMcFup52ZQYlbPRTFjEKw9Ll3HXUN3wNfe36OJtEfCxvtJC4U47ccYW7/
/UmwyvYBeXQBKLtZozik+Kr90DHkKeEttJLFk2erembR+Rjl2W87XyUwOePt9WrD
UjQ54Poz/OZtJs3xrXeFCeFT418wmcd3NhEkOm7uqtjVHIQNLpNaWirZWdHxxB08
RPJixaoGEIv9nkJNBCcde/POPdHFvRGwDkORbbAPItUujD9EiM+McpCTqbvGffDE
4nSnP35lfcLSp71ry2EjYZ+gGvy0C50uS50q++OM61EY8sAH9+LKKtGVJeQPBB88
oiV/OJym5FRCzq463EamzmfxS03Tyrjh1x+f7FLPbEylIUkOAJnPT3Q/IR6Mf+zW
78ILNuWVAY+5hR9eJBcdMukgxYKLr2kjnOWsCTxyxSE3imnIXRikIYyQs1o06jjN
bt859jmg3k5Wm56BeVGDNQmvbmdMM8B0bgqCgyROxULtoMZSYpvk4X6hBGPfVmR1
6u5TYOUFY3FcePkm1vTHmSUlK6c7Iui7NjEBVItmU+GtIPY7m/zY81cbXZ4oDxcW
yTtDIs4QAuGIrmDiKASKzZmm/pBCEu88Ie2Bwxsjc5y9seBZWnj+RjnV5MGi3XzU
ZGXWn49Hy1NHgqSwu6lvlP9wa+augpaWcg+5/yRTfbbQH58q7qucneO8cKiLme2Q
naM/B592BlDcryE2HZ737UVvWlY3h8pcR927JXqIuorOmLfq7WelkTtNlC8cBCpy
tjKynHj07sxkugxnv/WzSFWNFil9CF1oQLUvAZDnelD9pwGTbAagNyRpowamsvst
y0IjyQHzU4lJEncjopwi5KTSX70kKdsLlxrB2ql7NQK70b30A7ySANIfrmQRmRHL
x4yxldMF1utilpFQAvTgfBO0EAlmCb6RbjDaEODPATjaQScCYTPMlXTBROGiatDg
0U3ISHS1QxfxL8+HyWQPx4LiIwdINGu1ABwpbtE0f+3PXWZh0aympSqX2es/Di5r
kggv7vlsQZZFmxoF91DqkhSoT9b5vFIkbry7ayQDK7wYgNuKqUSkS6z2zyc+Pesw
mvztapZMX7A4zJhbNYk0nZy7Fj4C8ADVzwU1Y7Hy3dlxkCeWlcSVzAQh2MhpXyHL
+ZmPcyK+cnUWaH4J+QitFsT2pMOZagOpS6BETT12PdLZJolPqCeGAd05n+bd2aME
dSKr43kQCLbzGVKLO2q+b5B+LOq6s6YIQFlDR6fFNsstGf7hl+rBbFDIBm76jEoQ
Eavpk4jdcV3+pf6qq16dzPM0qcs4E1M0/F3A2uQeAJQabPfAGevC/NP/HAwlYiW1
QJHky3eu5iT+/xOXa6MV/2Me7TPglqmTjU+rqvyV5zOGqy9wwIF6ez/ymu3W6Qbq
7c8iPyhIvoewdDoB5tsabvH2CuBG2RG2SVEngacieXr3neM2Tu+iqUZDNcvyJuIT
lueGRmR/r7NHy6xvMvMUBkMLBt3RxAJHA6hPmwVrcyIXIEJaWlJyht7D6UaGESbY
byWcmhEy2AWm94p6pf5joSfNTtjb7F8ye+GUNXowKyLM7fZqiEp+5k/VGcoNU9em
xDnEbnnV9+7k4crIduNO2mF+lnkaXI/OB3EIkcS2vQsY5wHlBrfsNgiZ5mBwaNAM
vA/ssPUKIg52sPZAGf32TuRIyo1G+qlZeLWTFqG6S7BKG3mcJ/pMQrfbiu7tpjm4
gJebPgd4T49+gIomwXM4o+tt2x4fiuFnZac0hyxolSYdW/+jLKtt5RwZcm5ki8rI
OgiGwhF47vs1Xq1Ba4XMAAVi6mLBebEByGP3H4FuqDwpLl0uxZ7RoD43c7abGG/U
W/ct63seBQ/rppkuBzSzyCyTQlsmbTv3FmjV6xfBE09HyQaLkLlwjXZG6P5iYqb0
1GIcizFQgxisWSYpAMtrqvMWnt5ZVRo37+tcxNyGKDqEUvQOZU5ybj5mQtz3GPQD
4qTyf+knFLux6CqmQ2BR/An+Sa0Qo3onsv/Ey7DZ5ISpuXmHhGbtApE4VelHHw7F
q7HBjfjK78JAmfflMQAuxNtYhixDURL/RM0fx4g7mpXwuWz1VVQGF77UduDnuejM
f66r+SGdKfO80aEeZuB+G6dmXfFu8qGgic0oZiUNyxBGxMnV9dAh9UoeZDAJaHu6
WU+4WUnr5NpoCAaJi8IivKEZxIoyK5CgGyEiYmm1NUS6OdC2+i3M8SvZpqXsOs05
8CLE+zAIRwrpw1/teZFn1eFSeH6FLBmsEnJIO1JG1q6HJU2VoIyprXKDSlbTyASL
DtdvXM0U+0bzoMAYxP9Kyind+zSUlzfSSIMAYLEaXMRzlqcWEndH0uv7Q5KOOB7k
0yG0x0nd+KoU4thwLXtQjgUFcqueaNzSb/m9opC8CR0ODMU5EYGkywOS927ocQ+z
sxaWhPqbDMhxcA2XDW2/QmVRmtoeL8qcGbzL6Dva/vHbN1cem4hme65UZrahdPYR
7iXWOTVrHv5vml5hOKUqbz+AONMYW9ZPpu7xk63dwRI3qQz88t5+SEwzmMQfT3u8
Hhw6TAOOnaEgV2mKgkJuIrrCQSyTPXKvT0uOA36vq2JNIL+mb5YcnXKmFoQ5Iq9W
e9NZMOyzCPk7OXGmQfNqw5y+V/fXnVjmg6+Jxm58jsWQcovmHQTj9MNaiLXMfiSS
9kk1+cKv+2HyG/kLZ6Cq+PgYW0mt8ege7cHZJarPhZUgKvvLPwmHAcwyGYmimcmz
ji30avSjs/AiqVfJeL518LxVlNYvAxO8Wa9PDmfsL0AxXjETj72p8sJlxgrrKJgF
ADvCUDT7hBlzn9qc7xMcfa7QUoHiG9qOlMr2UpDeWVkEi3f5iUDYxhfKNQQuc5Sd
E/3k7NPpHUf4KQnXkRwGY48+0DSQh8RB02NTwd/o/wmSynEtGplP3o+hR54zgOy1
AuscS6nnIOVMriziwwZjK3ipYVc/FnzfmjOQZo4a8PqJZulRW2xJxr2JYr55G//g
yaHSO1SHsRWB9Vayt7qJ5iXk1DRq24iIpigIaedwJJv+6wrPZ5jMKtPgkO43FOdl
Th0MIi7ny3B1OgXQi23At/CDQJlUACyhsdB6BHGUgpSGyXu2GzZVhDOfJbt+mj5m
ZqKfbOMD0OO92xFBT8g43RY8HCQLI3TUgpMdf5TSSIM2RZOlyFiN/tPG+5UTd4R7
WuYvQkQLFkoQyBT+oDtFMD4Okh57C8QYzpoqtYTBgxQ1uyyZl2o2ArmCZLgE8ZKL
ID64DvozMigGPqOu1sp7pF3v2n+XJ8A6tSTDSiGJwZjR2G3f7+HZOil1HxzuE7Vx
SzJXvM/r7DhmIz/971LSvzCu4x7Ru1NnEbk5iZMyTmYOtfTg7PSL9pbGcd9vGj9p
Lzrdc8+xcK5zwSRykBuyf75xIytiUB0f4JyN3EIFPiWSGgedmsZeeset0cO2znkh
M8SpoILteUdY66I38kKzrxDY+lABQBS7YesHu3rf+13gWqv7j2c0tVVDS+qydxrD
TgrPrKDrtIebpUnsCQ6KLrEHWZqujSQaEHzLMRsiWwU7SnliDJAJIN+rJEtUsuiP
UVsBeSCaYxilG6upnr+FnSfsrxBzCoVdaCvpE9n9c3Lf8jTyT0g2cHEjzWtaVDRd
agL3SO2XI4eZIN+FW5IqLPUww77nALGU6dRmGaK6ws7BTNqJByF7DN3YnBQm+vFe
GLtYKOlotSex8bAps5grMkHXg/rYOHEeY62KGqWVQr4655SOVMuic4krHSQ5HLsc
mWG1s9uRiS79ndGN8e6C0Z4Av0/ooowDRTX6K4YOK9EQYjErLcCIq7izS/P+HDbo
0JdxH7CpwEuiGFSfvkldUXpVa/olkWu+PkwUlD+DUbQjnJZQTNs0ctkxzIyjDefl
j2FQUvjtav+MiiWomJl1tOiRYvS1quB/zzhxP/TysLX1tqSjuUuewAiK5gBDW4MQ
M7CIufUwpcSOD5+R/aLQ3EhSr5pAzWVkn/E9YwfNNTJLowq+f14/UEt3t0RfU2Qh
Mdo3blJfKfLzydDH4RIoYwSlofwufOZf7yU14Tic34arnK46d1rJx3s+3rcXAsUX
lZ9r7q6YTaQ8v7yijE7fYAQIhU513NRSLBflUCGVeKItcw27IYbbioi7cKsaFGvl
chAhJWsFd5i4MjUYJ63bT+/7KYD1qPxxO0tZhianLAFgNzxjpJ3XjedUZi14TISJ
1NRRveWw2qt+SHrWIOwqAwfeG2KBID6ad8pUQeAYWDe/mfI+lnuFXQM2/skObaTd
sQkxoMI78f1E+Eia4X5wTmlm8wl7iqqYP8j0WuMmSVCNwUPAGSnSDO+g2QNK3EWM
weJzH7CXgz1r2p+pIrX+jDlZY/dn0zxaWa4vYH6xn1YqYDTIAR0cB0yaxHK+4wdp
ia52oG8CE72SNNptZKa97M3uHE7xEN4KwZKPOZDxjjrAT/TAycYHAoN2zGlVyoMS
fPhI5VB0J6KD0iih8ocDeb4GAKTuhgb2d3ijigVJDsIrbY6lb45peK6LxQt5ejR7
HNiHLIJ9QOalL8h0aqkS7/V1IUenXj25aFIFo18wDSt6oZmmeUEyOlXWZEXgqCEx
bCHnlO5VOYafaX+pLkIdVKUfg7pJwODLjJDdFUAMJsz3OmsG4d+Po4iE72qqoi2h
Y6dyyBVgNHoCbGhsaz6wpAEaUSTZX1HMY1degC3gKqH909tSueGm9dvl8tSIOkL2
knQcZDgkgpot9DWVoFnAUVjjDaFQqIqx25p6UlLo9RBw5+z9Xg+cpqsP0hgAnVTp
2AzcJoYgl5S+uhPdQq4wLcc+Nx2qWCB0cDzjoC/CzvPT70tx9yLzafQ//CgVK2+b
cVRm9SHTO6KcHTA7EpAQBGMFedeuFpBCiiudTpff2XQ7h00VEMnendArYviIjTAN
xd4Snpj98uoFTLOn4rrFoh8r+FGkuYOdsZaYl6DbdgGIXl2C/XQqd7lVV1geu2Yg
P3e9eyEP8LgaD0oUhk4HiX8XtG4aGfcRHBx9NnAqrtcjFwLX9Eb5MDvAsWBqgN92
cffZBjpCVG5lWx9UqCs3dL/6LvvBMH8m54fYRFcpULfAe+CO/uAGmoyzaHnQFKw3
WKshYJAPIldzyQeFqCZ2bE89hvWF9UFsmfXJ9A6ImboCh+tX1OcGI4QlcwhJUYp9
KuBZHWhh4YHybnzmf3IIT6ZAhVvjMXP/74GED6/KZUUxzAAfypRaGU/94T/UT9f9
Nw9eKmSD04juJ+S2N+S1ceh43jmY+AG6NXiKWBuKJBQxupEoZDsq61Ol5eorTe0M
ro9rAkjO7yZoUfI4Hc5nKLQcl1V2LO50omlVXxl5mXu72VLr5moZdKANGz6Jspkp
Lxyo8pmx6EceFBZveWbXI0BrezpikDI10IOhKNJgfbe5aGl22egOXcjLfdnAaE95
PDA7/GCIAXha/Q8wIFaEtksKQ6unWpah7KtIudd23iB9uzR/9ZpIpy5gT+QalbVV
H7blcnQdxh26LCWQZU12yttdSZHYzoFFx3oLKgsCFvYqy/KQELRxDb3aV2bXVwxq
ImH6w6HIbqN2WwFP5ERXJIsOFBFOIavmPGNjy+6mmXJFEZeusnlYIB3WGpff0JgS
iiXv7ZZNjjymlLhK+Wo04hNAeYE0y0uDz8AjwoTF6TI1UEiubuLjeO4wlWemHFwU
JWTpR4OX1+WFy7bgaoLtAtKMUO8vkny0OkPbrBiJDK8BH+TBKKf/XIu2MEf9cxdf
LDKfipgCxIH/9JFJ58gaT4Xrk0zXilqdy17q3ZuI49IiY0VqTYxQsm+bBuyQc3QW
k11XSBnpr+XRmm0CDaTwMHFpa1wDDY7i6SKYHCg0tLGJjQRtxOPmT8X03B7eqv6a
7n2/1Vrz7T9JXVHs+mrBOB4Z6EZI7sPOQL0J6vzEjrjiuq1u66aMe+I/faN2QfIx
0jwLry4c7j2XTPuhFK+cd7lz6fna9B2uqzHTG7J1MPa2P6jcO8NDy0byIx9CjS+o
A0YH5GYnt4KllJXBlnm+W0SVD1HjkY6lOV24/JI90ql5Wyv0gIZEzBKU+KeOEpjZ
Tp4R3O2VA3hnQrMrK0FL/xbTw7WOxn0JAdKumoT9UsaElUviZr+indsfhyEoiLnJ
0IHutVYalVRRUQHmcyM3GNLUV4drPSdL5IZqitY/nd5gHw6CArCmi4w1Qe/uiodF
6aQVO8OMbZaORG9p66Cewte3qGko2IxHajE8M9t8kP8bbPehtgyPismiacGpDSsi
4x8pgwMCB9QcnWx7JvzxrjCiXMy1if+15PYRIbEbdBi0IcJspdQJkBdn05wRVzdL
pnf8+4xdGxM/mQ1ng7qpmu0WaZlMsOnbAs92Ot2QkCiU366lR76EoKESfsXvKHWr
JvhaLP2k13Wrq9Ae6PMys93YnAhRxKWaeqwh+mjDiHNjsh3X9V5p7sX447jEbVRo
eLz7bCfHTlmxH3ecVejUCGSGk/HzUxdwJfhePVLcrAbHu+yGqNyyBxnMmu7YdDLq
PmuRD66R7H8ubp3lCrn0WcP7gIRstt5hYDuthOoz1k9z22CY0hIRT81RCmG0ysEy
jD4n5+uKJCjki6ghk+cxfa6Bq8eUVQodoI3gTpl+qTd4gAG8KWo4UJWyNOXyGxhV
JGtEAkOiNiJZIor/pIF0CciGPykjMi7qCY9sjfFvy0ZAyr7wy9meUWJ7ezyD4zTO
s/kJyRrsK4QOVkJ1X3kMtpWCjRSGaU6fwwDVEmBhNDYfPnn/YwhyFTiMxqpVo1SX
iQsJW0btdskAOu1ka+tgcoXPIgWmBFuSg9VfqnIIaEqjSIA0FcnS1U1x3iqM1Dnq
nANJjflYTY6dPzN9BK+h4ZUkSVy4Pd/eYirvmckF0hEy25fKf8GN13YeyNkirq51
I+IvXfI0uZxYhUNyBBD5JJpzWZ86VxeSvr7WA54x6l81AH2Av8lHzuvTOPkFz/Yk
VBMWutBv91TuUVVQ9T9hNpIzywQTIeMj2f/8TdXk6z1UGH+o1WMfNDTpFQ8YyjRg
Ml72VDfbyMOsljVnCPxw9tnLE0jTiQ+Yq1g7Sli/LEZGkpUH4xq9Dz+zs2InFy2J
Lz9V5Nb9Ehumt8mPqpGQ4QvU+Rk1niV8FaAbPgKZu8AhStQF+cqKw70X7iNeo18y
09k3bTccSLFGpC3DFdwt95zyTzGnWNSmhs8Ua2aUzCgEWCFIyQNoQas0PYsZh/gr
Yu4uAwmM77QrVUe3CupSYmBf38AgM+N/iJtXL5egmB7pGO8XUvOWaBtRAujdotKp
3RJfHD7ZhtJGY3RzrxoD7nyKLP7xdFKngsXx5aB49bTD8cNviMG1z/s/sOfuQPg3
X8Wvft9dNNVKKlWLuj0RVrcK65IK0+FFE6b7kXUcEgo/nCaO+F47yp76/3ZABGKF
uQ5wlHMtvQ0RKn0g+DZ7C3UI1Wf5tGQQwcpnETkXLvUohoXABXHwXls0kVCkZGVW
OXprUIoTjrwMalexUAxWiEZkB5XVHJavNhSUjhxxgTdT7vJMbOdBdrW7qpLFUR2b
rxCAuMBOlu0Ck+3PRZQYmx6JYOWrH+MB4vVRfE4hcGBFUiT3XJNV99I4ZLXJpWtY
jNHeqFbEgb3sypzJrKtky4p0stGGUHR4nAEoyzYj+UdS+vJmiaLOFpU65A2xM9Fy
FiFAMTdF3JIQavDpiYeG5xjjLyQSOMUfh8DRNd0hTawEV5xUfOQd8ZTP83WGVTeH
vEZmaMIaoxDDqU7a7+KysAc8h8NFjNDVjgzvbebn6SONvyX+KD8ONst2h2SNbP3x
/x9mTeN+qHGW3Sqrqm0qw+ZSzwn3mLMPWamCUf5aKUfGPIw53vVfXi6j3LLGctFu
bMgtJP1fAiLwlJeFS0E0kzIRfvREJgj8A4mD8D+e2sne1YzVl3Jw7ykgwrOlbHrd
8DyEM1zzLxli3YFyDBVuKRf2KADpWxvBvkqCbheF54/bbM2CYarf10vdCIZVz2y5
v6QwFTV8DLMwoBjR8q+roJLLy/HePKXLXiM3AT5Y8I7ZUjulPDnZprUE/oMW/Kah
dqakQyI3AA9efzEbJ+Ugzbax7s0Ijsrh8mTeK40zjhMt4DNynjdAjWEwF7SkFpQX
Q/4zq/B+sSMgHqz0XHUoeDewg24h2Gio4ta3sys+IEP473i33XbXtdMyY8CHt7Kn
VCUI5TYGdNjuqPbZ1B5GDRJwBvJ3ojEUXmPUb75c2u+L/TRQSgFm67efR3Stk0ub
v3XGZHUlFQAZ2OSE+xCwttiRBIbnFmu0UCOveyYJCZBcDdS55OaNvfwVZ7t67nQT
9TmJrcv2L2Q+qglJElKznaSBbrgwc21+GfqLR8wijkyq9nz8+L3ftvO862WNIW/g
9ePnDg9flwCvOWPf1Pja6msX78EY1DelbyoTfiniMr7Q3hU/44FdMzk9FvJ8/UHQ
r6CHv9qDc7DNaBAY5Lda0MrlJ6Gy8Ymfqh7ole98XK0Uqoqz2+KSmqG+NlVU+FiC
bDKXtmFIEcIYzst8sMTR2Jci0GkWvdalERlKYsZKTtW1j9ued1weEyNTI7lcXNjP
xavk6vl0V9NZ+DWnwACM6Qaf7EeZY+sdWYRC8x0/AsQ+GoE7PQAEvUV/TF9+8Kh0
MY3skE5UQ9Zn7gTFfIbvWFCqCZ5lZ8YOObn4aBoGzn15CktqCOnX+TPuXUMnTDVm
El+K1nmcXtrCTZsioww003kiiBk4bdTkd/bw5wxzJ99dRnoGj54zvnbcAsYWnJYk
XWREu5KNpVF0wSdIb4cmv38M+q7hRB7fwQX7bDBsavRoqYIwVP9RiYhQeUCKTq0s
rxMlzpcEDBGSCR3hmruZHD1R9uXHTSDv8sXEpVQPzAMqYI7rWAoF6VpBa/4LpqRp
twLuP1MTmo8P4GHbH7ixT7bBmyo/lEse2VEv48GKg7IE5BxjvTPAidpJGOi0w+Kd
71Wu2esP4cE3Kl08/rfTRbm6A/sGYQU7qmV+S8W4yms3uLyX4jc3IhxJpYezAx6o
azSyUBZ1c6G4vmbcE6sL4BRM8HzwIhYmAL46ot7KuoXdBHWEawfyZ9HlB0Qw2GNw
RFoQ85Iafp960qg0BmXCDWSkRNfPST8xMDjJTdGLeuqYRmRrAajjk9lx94H1mHYl
XsVLNuUvpXxhlFgKlasH/ZYdKyx+MOqViSYJ/MmRs5NspQHCABLdk6hYr84zMOJn
YAKFGtmTnJZ/8ne+QscyqAIRILTl1OVYhpoGf+F04osRy5BhzUd8EegqqrFT2trx
qnpeYxKy4Q4uGlX8h9bnhRD8t4NSNxPnEWh7KQIy2T1OPqRVVArRivPT2XYW6mXH
Uqww7nHCCMe3OGA6TIgpJm7W8CPpynXUvVvbZhy+qI7R0DDObqANdsYP8QZdXEtg
Co9U3ydwjHDHsGfBuxjk7acM2jHHgga3ozrobqYL/DU/LlseDOOkxHvgpjHCwsks
c5WtCc6IYgjXUoYQFbJHwRWP3a4Gm3l83ZSLn0XRYJbmi1gWKCDVtdEOp2n80KmH
t1hIBKw/hzHoG9cZwlT/Re6M8GTAEDaZ874xr+t1qBnUldMU8LIPc9mFfZSHtOqK
BDMmH95Xf+hHKOUDUGOUQo49PHF7BZ0Ee3DbpvQf2HAGr+CfSnznXbyf03aIrYG2
cHAjUjofX0SY6QDfNYuDzx4raG+eeTb3xbUgVrYKAfWZcydFOHFwlHXB7FH3hdgn
viXykLGtW+lbaoo+CG1KECN6g7NeOEDjRuu8wKCsi2bYlHRZCzsbsBIbjotSuFv0
GLVK1VBclFpqeuDzV/lKndBFWe2NJME/M0kqlm6xX4BlyoLDcfwqcrLLUguKSRPB
xL1RPuq5yR4u9T0lsXn0vQYV+nadkEWckcQUrOrvU+NFzAmETvMVStSpNxZw7zS6
iEHXSpqxyG6lXSOMdF5obn8bQBpdf8eb/ltcQrE/hrMYdX51tztYMRIVRogtJXUV
8Zs1nDJattAOtdqftQsjivCYHTR/00WXO166UcFiVurS/MxiNTPlp8Ax3BWCIGDE
9JB2A3fCkzoEeRH6fwcGXGklsLTk+uoz1KzfX7Q7qnAoEZ6PU66LoCiieRdutp2V
zDhj2CTN4ft59X5L4woKocbAG6kiGdhyWBduvq1+BrWmTzBG/86kahCijVrKaaTU
irwY9oq2dPg86lsXiQOjlCtwW920F7L1T4BpZ88QeTLZsgzctcw15gslIH0CRShM
kJFgnrrybOsjfiNC88lEO2KJLin4lBJGfNzxqmk77asfgH2dPe/9F+vYxeV1iqCk
Rivd1VERrI6PqHUF9O28JTzOCcG4s2ts7rwDrIV43G5b+4xRf0R8M+iP7AF9U3Q5
2zJj+SvCdVk2SavAyKYd1LuofrRkO3TbtJ4MrVFvVpUEPH9hhgj66BvjvebGN117
AEbp0EFTg/7oV7h2oLVO1iN7lrZIK4HrYfQkqg7fdu3UjZzRiZOMiunB4DLdZGUO
p85R6ZbvJIj+UOEwouo4fuwHv+poJ19bXfLsef4wJ7L4VX4Kw4BPJ+9n0t+1p7j+
Ecll7Fc5ExmN7KGiG8co0BgbtQBE1r+HrDYZ7uMKqkWVjx5UFwtKeYmK/6WyTusl
8v2g/Hy6V71GAVfKq+GZh/dc6GC88vSdV1s3z7eMyzXIxokwjwqwES7AeHtkGrh9
okMAvafCXcYsMYfkZg16J9kEZy/4uqlSIqx2Rmo6ggEVmEcp0hwShDbRpKnYZyfr
2LCm9M2xuovb0Yr0n1T15t3SxHHNDZ3+mwzagEiFNhMp5lbzjNsykLnyDK/j8wuz
DLTiZQD+R7LIO8HEmRZll6Qqrlb/3XBJNUQjGJmB4krQ2T4ek75XQa4NdsmpkVY1
oHIuxeq4PIf/HDlAa/CSLLIhyJtjbTfya7Q61cATkcVNMO7s6LRVWTttcoJdU6KY
E6tBX4sizfHuANZzGzA16+07cTHK9/5pB8sqjpwp5LdwwwQkMNJPvOb9k9St7yIx
bk2/WLC1FPBe5DY6cqM8r+gujMxfrXqOKDOy8+vER+h2qBxujHyJARUdkfH80qIP
Zs9xk7z2emyXWoWrgHha4/mSZHjsX/U/3FC5cxizGXzGbsio3WNkVgauAV+aWtxZ
x4efobyK4+fAsR1PIygLjO0vm+zeC8HxvBr1BOro6Tcgm189kl4tE1opoVAWU1Y/
pwsvOpQBugx8Lyrd+Hq8leIxQ9WT30r1XUQ1qU5tWzEk4dVsliqdjByO+RThyxfv
jvvv7V6rtBbOCWp3tGRQefX+HrakbriznUZc0ESXn3pzZV5H4bDBRzMow6gDlHPz
qK/rMfAB/91n1FwiD4HoJ4CqFTmrR+84qSxpEIngftJM6WA/qhYw7oPoTXKwndlS
sCXc75THZ6dHmKq9XwrZXfrVZO7QLTHoiuSEPYzPkgLRN4bYbUg58oJIDEJTiDwb
TsDeNjuKoleFs4c7AMN7O3rukgeVICJ7eLQWXXD1P4/v9bQcmNl8zW5kDUqGW34M
B+MYUGNp6NB9YXyjAIVlGgx07/QOADj6gMVIYDfDyWpARrp++gN10IcRueJO3KRi
XL1Q4VXamVT3HkL1i0mkrAHrbub4g9iNi6t0I4ztfzQj22tOIn7LdniiVZG8y8In
dR1pJpsQFbB9i/CjtOoVkwQRPZEEnEViBQ8kHgIstb0eySAzwng0yQrPPYobZ8rs
Z9GCym15PDqSjRHf3rS9C1B/HtJOQLIKFGMZLhYfm73HMxy1m/F6uuz/7ewMwKjA
CCVpKbdNeXDiklb2Gmi2EGgoChol1I38AU+DuvOvQKa4tAAWB0fUvpPXCG3i4X/n
2Bm8YIlmD9tvXWyqgIF5msbFyow4x5CWwyoPsnTGnnSnpH66IMYl7FQS1VVESHqn
tdJJ7hSPmhiFBYuEMuag4p04OGnsvdMrqYsNiV6GDhUunon26jiwwBxjT0eILIg5
4uhw6S3LJJ/GMbd8I5u6ZOKytlP1IbWJc0ehWjFConM4y/5c9WNITzB+qpg49O7C
9VF61H+EFpl2AfRHASmCj/Pm1ZNwryh+P7bYkEHweHzTNg/pOnm7a+LhDFhIHboJ
ZSnFY26NQMdZw/w3goxstQFtRB4SXxMSs8jnFuF3mBRsIwlyo0RYbej+agVcgCqp
/7tVi2qD5FBo0XhJ+EGrpJ92PvaFY47faJqbqbYW1YmRDUbGNdu7H/9CzCXhw2zf
+V4bMR418gSK96Dt+btSjvRviO6zuqqJXPSWT0Rkg60tITPm8jKAf28NAlARbVOw
UP+Dx/xKvk4B8MvEIs7FlP4M83/Fl0Y+ps1ZxaW7NRKwlpmxoKM2/XLLrVUJDvfe
gK69XUd2NQFkGhGpkn9bXqYVnKhjOfSMwfg0esv3440LoleKuxn30a3csr5RGYb9
M6mAEVJNFe95jnVoHKA5s1IPyY+L+dFY8Zttvc8prNpchfhabjBWSE9eOcPQ4Xet
qDYFCTerkSZGLKJmizwsOi1r9xEyH9uu0U5JJ/2TTXsSA4qoEytN/6AOWtiAxXdL
QkDLK1n0v3OODSBhFnKV9QYQ6CJmdTP7nUefErFSe1b/NLRG7zTHIESZpur9uBjf
vRsprwUfcQ5ScLjXvWxONreBrADXBH46WAzdB7nelFpRlj+Gud2tcZ1tog5UGlmL
B4BdOGxUJgnx3MICWSTst34+XRsxgJo300NG89+ZLSousJhXIYBTzVviCe7iyHhT
vnbW/EDHKQ+Aie9mP6qUGRFaTnrfryHB4Y4mk/IGlV5ZeLtF9TR/BM3GXlkMXiAY
IJUQZqIFrshv/ahCiLC/lYGzte83syMKRB2VprUPSxCo2TBZKGCEawBQTZBe4TI5
hIeJOtHr1pmNrURCRSllcG4em+qXB4LmJrauMokkzy/lEy5iBT8yvXKZM/0JbEeb
oXMfYJp3k8gchTlh0VDla9ukIXFfQVbevQJXxuktrSFHQUOyCslR/+KBnNc2kIjF
8dT0+/GEUjWJdH4QF+1/kuxSOnVXnO/D09YhJUuImiysvxAW5onRhkHkw5X4TSVO
vhKrBWoogWisGuw+a3yDNdqhBsZILe5XjFTApk1JH3LDByC2FDwMdvyRRILeCAp7
1Ri2fOOeKnlw0rIbH76VaipSeHPgb1KRe+uVjn+52KXJxm3UrcE0OByEjEjN+bF2
CO1opddtFvzG3sVZQjf//0Q53LMMnHX0TNMSVFuPsxU7QHqephceXnavGX7lqvuA
0TLoviWOPk58e4nVhlpFB3dw9wcqwQoMGGD9iPkxVZ20s2PepP27n/fv/x0xVW2v
omJerTiXQ3fhiqCQJVxNnNxxBlcufA4yE37YWB3uWwffCMoIrBiwGJ3opnX2GSFB
AByXaEv5xfh+l480Q9RENqKO4QLRASQoe9DnwkJ8jjGGWr4jrKGX2DzOeqyHpoKS
K9T93c8e0gaUFwUk73tLef7PaPNr9LWEiniffRAsFCL2FjIfDQDO5dv/BFc8z9Ss
Ck8vJczLN/ZzASMZj/caruFe6/apC2ZuAN3EtQ7s6MIt8IuDO5Mrdn5rr3c0DWj8
O+VF5fsi6CtamuIddrHsmRPI5Wjsa51I0yahRqGpBqcZbsCyOP+qg3Dn8YSXjhRV
JnVbNX+wtP0VyBTrrxXil5U10NuIBb/t/IwLvVQNNP2PazXD+GkYWj5l+j+7pBuJ
+WuJMOwnpw7Y6FNwAIW7B+eNels2qYZoF/kzH+06DfHIkbih8Mz8KMtwQL70cPwG
QTzktt3w8Wz545iJzQ01joBqUJ4YL5tOn0gEeGbK3E5h+lLeVH4CqwQtQhHm5S4U
ko0r2TmIOUmza5vmAozJrC1CFMjsUCWn0ngbNWHqlHKj0Pt3i8vj2uQV5q4FRdNK
+CQeEhK8DiiS63zM/utecaObhc3hJXP4VjeLpddrPboaQhrYm7rXemsgVhqZ1jAI
uSRG/edv87XUbMeEZLNLlJJs5akL/q5Lb9vB87MCeB0hiHbscMKAU5jc0slcPuaZ
DxVJdy0MhxFZs7VaJ0scQLTjb5fA+fNoj2yOLS8wfw1JVu0Xzmeg9h1P0E3hlZqs
fylJDjp5Rh3cliMLd7zMETDB5bBy5TzACxMJ2ZriwF3Da8tTLgjuVUTxsnH+etPf
jwDXX9fsrQbkFl6vggyu5Qw9gz6OPHnkvElxH7t0ScN/jwSAP4ScTx6GaX8lD4bf
GJeKp0jjn37GssmqhYncmEVPP14hLUGqFTAcQEa/ioaU4JqLYKfQXliYoEtRiQwt
y1AZ46ZzfFlWZTKoQG61jzV/8GQRkQNwL4x8OVh/BvDggkVk36yxG0cXO/B24+Fc
OJx5DBQzjPdBXMPlYOodWojL6WkaDnsazysddmYcLSUxzCF2mLNhzHltigj4cOOn
zaEymz/Ha+nzCaCvk88uCt2t0umip3nSfruxNtKUHt4z6VkMbOYuJeodNlyg2HES
5HSqeWXBoAuSicIN5t+VnspM0hMEVL8WK6TzbHKGmPCwk8LeoYRchyARfUfPW8uQ
BA1s9MGvcggH8GRRvDaF6pAG6AR9HRjfdVYtdat41ilr22VxS5RccX4EcJ1WPDHz
YsA2dvftKw2G7La1TsXDktdA8XyvNBURRflK7ptHNQa5JhLD6v5YDLqqiObCg4hA
ruMfbAkrK2MHjFMXWDLfDknMS5f76ID5WYJD0vCOZqni6tbwCA92Vfu7JGSEnJL9
lDoAHHUYDZ42D+Kd8JREubqCr5N5QGqhZypor1hTgP6UU0ZJgCYSbCTtW+uQjtSI
1XYNll/fcBcUq1w0R3SJZUgXGN9SqFQ/4kEBHhXjauSBNUzaiLudaENZ9JKk/lO6
2ynmc985Q6TPFhle671I3uMKj4fkeAzMbnwGpbQ/3pWmF3jVgmhr/+8xw4T/IMr3
s5OBeUWZXkvsCEeanlaLswPvhJffmmbe8/p1gAFJf614NPSfq2QFlwsVuQAthh5w
GMTJpXLILCkMVa3oW90Nf0TfqfkTObo9lgMkgKa87KVaPN/eIhXfGM9s3anrUrCM
hCAX7RdzKpBsegYjVkyrktNiqBQnZ/KPWugllzuCjCer2W0+HkzmICgL76dmM129
UIXd0ae6sUYGO0+Z2UlrmgUHUcuLdtesjg4sZmg45T0SR79vKXuH92xeR2fNEd4a
BojU+xfcIU9fda3ca0EpIoH1G5dJnb1SSz9bpRo+KOiLw62ACtU7lBgQZ1S5Qc2a
oPwVeozHtYB4TvkEAix8VCEd7gGLdt+cvDjZ+vISZsPgXT7X+xObDGcNG87pxehp
m3tekQFuET//rDoZN2xuUTx8uBLDJtoHIPJxzkj3BpTADaQMhQ+bT/PdmE+aRvvG
QQ5yZVq+N1M75ieJNIfJiFd76kYEV5Y6WcbT1a8ARufZrnDHNaR8po1ptHtKIJZN
h89Hs+z689P/3DS4WTitgY8IZB5yNAcCws4Oe9VXQz0ce8J55rpkkCqWDAIYqNDZ
ZyJr6Ldy6vNcU1AY6frd4eeS4BPtGop4qkqaL62yDpLSi39X228iFdWpyrWPEWJ9
MKiK4iY2unlK3yrB7tARwucalye61KKif3ITjQ7PSDo1SVhYwf5R5wjOTJO8VBb/
n4uZ8wUsu/Bqq+Mieuw4xlzVjck0QM/p03oaKA15rC39FW4h8Mf7Y6fIDj6hTNDI
bUXljGmZSZNOQie8lWHOp01RMt7HD344G4rzlanbGeFl/1/wLCVmF1UOWNMwAKDQ
7C0E3MJ1gKXGEbhxbgVuWEPX6J3oKSjKO+GgK7/rCwB3lWWT5hXCXP5Gda27BZQJ
YNDzVwfsYQ5W/re6WgxhuuLAobSf3CP26bGLcZpxbbq0H/Ib3Wo3ii2ugaC30s8T
MHJ6CXkJLsjMayDmWd1humJiBuzkLoctOrgzxJefhZaUbUcKBWHs9GUv1X6LeU2w
C1lkrMuYmdjZTqqvA7nZTFwPIRvPjh+lgyKAd8ClbQa+gkPbn7/RX+GJEcqjS7Dj
/A1GMBXZknkWAZ3h3yNLgekszdXHa2W1dUXZp0tgNnflGPoy/XPwJg4b1DlJlPiW
ojmJ5sldt1WmeyB/nyl+ATdg60Otvwf1AvvtpEgKoaTOSLuZI+sK0ReUKT/k319c
LusVVUONcTF/Y30JH2Su+gKVgjybde7bQVTFwaKlp8EP1VVPt1a9TO5Y/uVUX27D
gzKIQgTx9h1XXmXoW0xzbqhmJ1UF+abhDFmZAFFZeDVz6Dt9bO+lru/U0b6swxgQ
Z+ysyN8KiiNi1xu8WwUmG2kJ8NtyLIPBLkK554PT/NnA00iFWhP2VAPgek/BZS6A
cGrV3teKq0ryMj0iG7W+e/zwi51TtqOg6+vOC7Ot2ZiNpy4dCj7LEkLlLkhcljS3
t84cX3vg8pjeMjOHPDC33MmywDsSxl4GV45egkjUC4PjQ6J/JHEqOBiJQUpM6zec
vZbUVh1NBTRZUUnlJ0CijIxvRHAiQPKpXc0MCI8jDS1xhI35CH1+Kk2Nqo1SInDz
J0pDQsiZBmX1VatLMy8MZv1Bioq3Ez70a6VaMDNXgi8OIJYuSLo/dpLRzD5qCg42
k4bGwJYVlIbWHTzo9jFlpNG6B4ecaFhxfAxSmI5mQYR/SxaaMpE8sgZR4LRIpX7B
QwYigbBbCouU9RZtAgURcw9gf8AXU6Fzn/ilkjV2lO/cW82/DAIShzwCbNCxCNt6
dX79IXwNypJKrWfGj1A69G/WrhSVYqs9ud+OYK9dXmh5ydgxOvXXEXZo/u27NG4B
l1jLx8c2+ZDOJWTCDa+cvrWGLs5vwXoB12B/a1Ai+u86G/W+DX3xDALfWH4Iq2c0
gmXrPURP9+Pvqr2siTTHq/PGX90o1rb1EBeMT+JvpQyQKy727vTyJ7sVRcoTSeGv
5k/riE7JqMUb/sm/8che3WkbudTKHG2Q/uqyCpxvVZS38IpjRTKJZR/xWN1hdJQS
xWypwJbPZ0elGjhqi5m6F0RQu1bHTnbZyQL2Ne+IwsZtGUDJJ0nLXz/wpIbg2vN1
ShVraffxn8yrSDC8+pHpHntbmeq6TaEf4PTOQIyzAV55epsjiVFs1vK4+YCsM1jt
7WPtmgMTrefbHDO5srNPtTZjcAceAGwq9ddMFEMV0Ep7TcD2GCz3VALpNp/Ue3PU
tG0trQ+shm4dXnYHH4PEimKKLoA9hkWmEUGDjEBRca1W3YrWDoY5whyx8s3qWtKz
xKXRwK870puQrvTOCe2rZux4S96jqBEOzDzYSUXf71aCHJ2rsHG5TTjeG6EeWqc5
iRGgFManaZL+4SSm79kdIEgz+/FJH3IiHrJTmLE2i2THQMywZ0tE0403zOYZ2Myl
bxynLavoaiAHvmWWzdxo7UDKy4nU3TTAOfToFB83mevAiT35RDiKrYT4DhHU6EDK
K7bM0vpuNfoHq86kz143AbS1xVhWCk2eiipstvl9enoTUzyMeVjcwcysODU92InK
YG6CWBxToxfghYSDfdrKnWJDgTd1xJ2YTl8CabvrBJmxcbb+tILJN7nEd8/VwDJu
a9Tm7L502iTKdpkSkXaB0YBa9afHg52P71ibqQd4K8UIDrcfitV+c2ZdCFRVSE0i
mqLz4D1EW/vUukQSyMEmPa+PpDmcHstMwVeyG0wNzNEMbI2TZhX2BEauh2EJcX9M
gBpfoNFnUTWewubL4u5IgRfAYLiy4LgoJWZLfgiFE/yjGS/NghgcxaLEXMC/ld6N
W1COeaEr+NjCOJKq7IwB0WZpDj8cy+1bUJJzTuRABHx84NLbwa8DsgYynS97WfGY
b5ZS207pKLXaqKrDYxA5mrKcWlM5+6xHzA5i0nvQogxqOzDVbIxlOvemKQOcGnPz
aUwPwMyYknurAtWKKe4CY/u2FtV+/KxI6EShv2P/4kuRNWY4b6jX3ezGEZLNfi1B
uU9JDiIx1CJfuh62iUZuUXdpKjvuM3uzSVORMpN5fHEBgE5lbzpNamcvHDEaLZnW
v7cN6kJWMa+2TJY+EHREvcOtEFx+NRWU16XH/fbeGxZjpqO8jFTQxkIV8FYO4g11
AxVa0I54hHXVks123SD77F9l97os3Lgl8R2JIrz4pju8GCJNrooy5LAWq9ioLyKk
sox1X2NtIThEuL/BBtTj/qKWHGpeloaognlu5gm5beOg1YFMY9YOdX5EPYPZSn8X
mEzWf3Dfycy61RM36dakHtIddbI0qWV4ZKKHgckGzJal7Uz88P2VSxbl2gSvyo2v
LGC7ejvlLGanuPm42r3xEgC2fN1GBgDyCyGUGMjypafzldTU0OfqHrrx3kDJST2K
XKvl4D8EbShYN37kqt+sHD2d86uZ8VuZ/AcId4xuKq6MMHSpnzOQ1lJwNgYy5yN9
vBbtTQtpAFkNjGlj33YmwGwM1VczesiVxqUqUtJyeGmKwGyOVvCQUJzuaS2+gi2i
d+wA/n8JrXxhBdvwnIpfLnxP5kyy++N/+uKrB1K5aNxMzfDy1M+bzcTU54EJPnSL
IZHqP7kuz8HjvSLo7lkl3pK+HI92rXfAkMxRfDeV+uOelx2M8eWzUjurFcvp4t3y
SytuBj7l8mjzZNNd7TEEdZoeB9mLwDEkllOaeZZ71vzpPP6/ehEFhLOXgn6igRX0
KpPqsLJ5epa5HyLmZLgeCEwx/4rp4Erwal8O5wU4I1KtV0V8ss4rLeAM7+4ALHVX
aAxhOmn/aKQc2bkFC5PeUOg4xdbnx1x9EinKO2Ua37TUAdax6cLm7OjFjGB+/upL
7nnxHe5TbdcaY+XEXXqv2fC607cy/65u/OsTyeeziLzCHjOQJN5yjJ5ZKasZRmGS
5sR+x1XdN3mqYEW0OYA8X/OazEG+k/EjRrHCvexLUTza73+7XtayJMjibP0ggwZa
t/69C65H4UuwultUOve982zWt0ixzERnug3P/euU+EqzNtKh1YiVSRKheorSPTb8
eVB/LxEnbTovbPb90ugexrSdmZmQRv3s9AeZ78FMJvmFYCUoAi4TZI6v+BQIt68S
W4twABxsgpJpPvP9ftjBPzMUGNSzEC/IHModIGD74jKAJvQizY5sALXIuV9vg+Tf
7kZBugCzHG6xxkuJyQk7iZ3awHpywKvZuUBAs4nczd2gOcpnUcWHm6+pvEqZxf17
eUZ/YuqEJoUG6KXiNhyeU1JIxzyBaQTBVK3ZT5iS65uhCleVgV4eGdHfoEmTWOMy
x1kfvOs7gIO/J7NLHeJvScFRhLN8PBcgxypf7N3M/gWY2HQGp1wFbSjW6m9wCQIM
h5gdavbtQMvrAvQNaPAffEbCSOzHUa/GNZE5qesCPEAudrov3SzNpHoKhxndl2Tb
DYKV+8pynJFWZHKJvnSDBc+NqrbZmwMGGs8m3yPNQRqHR1Tzb8rlbcGXx75GN6JQ
NQUSuakXiekJqdHW4fHwPjjdLT65nk4G3DK2PRfsdjG2Z7AgbD+NQ7TQMNJnGD5m
W9C6eTPn35UqajejjxY2kUqNC4netJRKMXkEtuClomca7yAUHAgUPSmFNGuWDtpD
K1caXKn47U2ixWG4xG7r2kR7b+CvR5x3dbz/A9JQbkC31Eg4ns4lAJzpUmAIcztE
vT6ciZeKpoP6D20AHjjIVKH1ORF9gH8AMyN7NI4cZMp0KwBB4O5/zRtWK2VmKOCC
oQaB9qZsFtDFJ9PD0Z+xlZYWCd31VcQqe7Ozakc8Ps3vNssaOUjdeHHVjRTvGyuC
/G6mhMF4ohnoPpPRJ5642qY2J+9c3MEhwbMjhQwydQ47AYnZoix9LJUVpix2blAP
195pofzeaMpc3gDKk+JKfXNWeOrR4CEb8TaBUHAS/UvDe+ZsSlP7aV2rOHKRSC5S
`protect END_PROTECTED
