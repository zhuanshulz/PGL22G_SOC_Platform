`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8/6S74yljYWTLkez36HIa4m7o2mcTfQNZ5co737nLWf1DjYsJWOTpSKxhd+gXue6
ec9Cm1kMDaVvlcalyH3ObxGNFHCV6G+ABmp4B2RabYPHqLUGpTt7MiuLk1AJJ7W1
753DNKY+lWCyeAThUoEU4y3gnT/fNbb5JN1GDiFBRWGEFmPH9SDL9T3sQgO+593Z
g5e7FeDM+oMGCfFf0I/nur+pi0zzfZUqldqgUjzsY4DdsGSxV1sg3A2mWEU6n20j
Adul+7vo7ThJjlFIrZul6aG2bw8qDDkJX2CH8GXjmxeTXFSWk1IGs/ShtrXXhNpc
xpqCxM7JiPnMXwIxnsIon1EiRT6Q90E8TNtc4Zv9rT6RRuY1ONnxrKXya/Sk0Hr9
Ksza9qzmVaK82xVN6ulLpNjguIItuhZKOSXEF05nW1GCTTWLuFamkhXyil9DdbKi
06zG+HUxFpTU27Q0v54479DcFtCDpR48YCB4+gxs6QykIxkZOVArnvUYKrixP+c/
hCdHxa1z+XAZlfDl4t5Tywlf+uaXToVLgt8j6m7RzBGE8FGmjDchl9UL1EX7KhW1
agpfFsTuaOuQUNQTWFrPrDQZmKJdArY0aCCoZUKaJWARv6qac0tRssuK/eR9VwxC
ABCNpJidz2Qev7HhHgOL+GJYBT2grwaJEAPsHAV0gNUiCjy2wWPEhX1jjn11DMhY
tXkAFjdH6i/8cdoNUey8JH4uOOPtpb/OzF8FkpQ49Liiph4DOe/rabYZP8dH7PYc
sH/5ecdxWpYceyDYe7wDDPyMxUx0KNEio1DNtayc5BsKnj3fB6IZzzTE0/rB/oNf
4/dDLuHJXXD9ymRaoHsFYrDlwLlteUeC7MRX3u1oNHd7MI7JhE2B+kgKgxHZ0fhl
F8q/EFwGGbW0eyy8NPxADiYiImZXVZtyCuhfuW75cWkApzsSiFTOG/fN0I5biZYE
cuqOkhKp9/wvyASSitEO9sTWa6UD+aG3xRtqvux0MXp8JOZNo066uri8We0dK+tk
FSQbzAF8LXWiI9dVFNE/MlTY69TcXsFUpLfOV5Jny95h0iiNR2tkFOJNUAf7Idnf
P/OR3r7c40wIA54KDSuaTbPX3e76lmOOeUTwwjxC8ohQAoVanEbsbtgnRUIPwRbm
20JzLBcY6mm2ILlzxCk/0761xrHIOCFLR9KTClXaC/nHOi7GQwEbSuTEoDZdMsrZ
kWQ76q7UwGgQtuWh4M6+/UCfUmnVmidcsbxvtQt91vbz6lcF1SnHw2eBZv/uDEeb
zQnX7V7vBkr7lOoJLshZhxMWRZmCnzcep260CYChW8bCpN2hLjXgGwcsaNh7OQMk
a0cUjVRAZWbnI0Gwrh6YoR51v14TJ17UAYfQWK0MZysEKdQr03kmDm4/yrdjNq3D
5bwQi4H/w8IxBIe2WWfJxHeECGcdZykMn7Z9QDBLBhSoytE3UUzdQy3E8ROjr1n9
iOKYpNX4x1MORtaYXLWd1aVMYUSeVJix2X/W+hRg+0M1JPLsI2Cpfy+jj0vJbEZk
NdrZzWV7Z4NJXB4C8KJdtuz2I3zaJprsLZimalx9LZrrMB3uE78ntTNveRWLLgVA
KtJOzpTkqy3zrmoVQalg5Q==
`protect END_PROTECTED
