`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2ujjVpcM3Fqe6M/d8ZZfLJE4yAsANbGHJpbIQ8TtDEF0iIMG4YqMp/R2flKDYKSK
io4bHAozncT4ROyxcyBcEiSzJ2WYmwO4BTvRuUuogpf8zAiSOqEhfUAcdZShfvwR
SJwRjI5pf6ZwSPGOvURPug7R2xtgkrMEOIzbqsF+D3VqGLZFCw6LA/Kg2TLN98je
UkqIf+mz4kv9M9/SC/CxEW8zfKHhtP3D4YQcnSLwWsdcUvlRaYenjh7LZNNMLC/Z
cdgqUagf1vEyh3plbt2/y0scM4rvIPohPomveKd4ks6hCSlMV4gNCydJmZYGQ0UM
Hl9Uujx/hhnRSM8QcYOTaQL/4h9/BFLhAfKAHK4n5LIt0mmg3faWQLrUWyaR+2aa
qqCrJ9360E5sXQxFYGRtSBjHFmVenb5XneMjnDzaurjbHWvl0vdQfablt4sknAj1
WbYgdsv7ztfQZA9Ah0IQV5PHUlbxit+LcoiZUApjnLkwNVsVpQyaTU3JBVuPU5/h
`protect END_PROTECTED
