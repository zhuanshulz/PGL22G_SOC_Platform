`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZuY6gdQ5ztzxYbk4uP1ee4t/W3RhW45s2fkiZ43wYKhKPs82tMUCrqGBeyxTRMd5
vyFBmyQG/usc2YaXoZjV/4/JlCMV1+tNv+Vt8i9zE62D7Z8bhE6AinFo1EDRxrR7
Mcl11t3IgLioYRSGZ1+ssYdA1gzskzlUClF7aMjDxayFGZD87WvWQLoYvAopTS5v
4aBZoJEQBlTAF+7Vpu9vrHM+BoMK2TtwcpSpw0JZ4aF6cuhrM3g5UyxA4vgekMu1
k79wVCdIr3RRHBg0g+a5N6CFyf6JTREH5u2po3zy8/VlcGbhbTwkz2Zw6amMzUg3
rkmtJi9iHKjRYz1DDkO8Wj6jC3LM9GdXYVb10EELG0rGtvAYi9tUo6AXz8Sh3T0P
qxD/enK52azwRJVA8oleGE27v6w3gWuyKW23t+mBKizIAAqPWytroMtuoJm3PTh1
TCKkgh1/P09RbiMwBCGlPVOyrcFhZ0jrfdiAGhdnvOxn1MfUoksCht62KUEwcopz
Iv79JDaWX/FO9OUgWCZx7NoGIYE+CM51Ys87KR400li344PXhW2HmDzVstMnkM9Z
J1K7fXTAmuevtTW42K/iCUuk3a4KKXIqYevcjFlekEAYOQLOZGR3E6879eOu0XH+
uydIBplQM0cKac0bj0x+suOFudxBIivqBrl/o0XCbKwDRP07qThExacd03xi3E2D
w4aQMGPLD6JnCLt2xsWEPEwVzWFUiE2kMkXeYUWouC1SsTq3IO2F4LWc1Uf6Wbjz
NcT8v+BAJDe7QfPHWO6MMRPkVMDRKqgQrdBwqQ+M/Qm5RN8mD4mT0RukPhhC7DUz
5iGo5WQl+bOPa92zgxrjTcKY00ggHrxOkZ7hgk4eG1kHXSlTSW8NDAM7sEOrr/0k
GzRKKBuG4ApynCr4BvL1dvfZkqf0SxwpWHLMWd94JvyXWqdbjryR0HnVLtV0/CXq
mPyC50BMaqwzQpIpneQdpolmrzBYb+Eu9G1QBXhq6U3iOpxQC4woeeEOTAQSj5t0
Wpach3mDjcGSBhuLoeF/i7/sritbQrE6SR3GGENLlEhrsNBZLpren5sguWweEfNg
e2w1ASgG3k+bH+jD9GZAF6TbA4YVph+/fI+XSXDmmmj27ibrWsAsVGByiGuTlHo8
p5Yop+IxsS8atQUh5KBveJPIwlvlWIK7TjXLo2ImPN5yTnLcBsbElbDOOVAcZhfu
4zrKH8ekwpRgzg3s1RBQ3HKDuGaHg8c7ZJAIVpNvwO0P4aLrkBHBELZ55gUYa3hb
x8ifjzu+WrI5BKb9wqzZvvMO+CNTcw2iI2lIXxXTIgZjLwG+JdaHhlO4cW6O/Q4n
cH1i0NJysN7xXe/BSyRS196aAWjt9SZ+kFvLLj1igKhU1aM4QPA1RsVAqbqwghal
ac3CTY/rd/FiU2l+zeEmmVqBEaLHiTNGDh/fmzU17iIA/JlRHrqAWt2CDkRO+GXQ
XP/riPBODx+FOfHLTT+Q/ztnyXBDPBcdzDshXxT/JDLY+hXjKG+MkTl9KRtiM6mX
sZlVrC5Vno1gBP/vyIZEnJrkokgh2c6CMq+5d8xzkFNYd2pUYVX0zVA+SbOrbjFG
BKoJZ6ml9cRBukyUSySgAepPiGlSYi26VZj62Emo1jrLHLUpcx/jo/8uYPh6+zTr
LA89s2ii9W0nnJLXZdvK8hYd/J4pg/f5w3mAWktTPBHXHpEvpCGL7nArJ0tuj6f7
w/z4ruB3ImwfLruKc1TFNKDRrl0wee93PjNRDDvFaih9DI4s4n5gvvNwFaIgTh/M
ygTqVGO9z6LWhowRIG2O5+yhXwNe4qa3E0Xn5r1J8fVhts50kthJenBgCm6REaQM
FNAMVuhJ1qe5wRxCtU88OFt/PWx8CnsmXbr3FUfofq44Z+CM0CHolM7EiT7UlGWI
wjejKIZr26yEcyYQ8gtmsCw9Gf5B+esQFkScRgnpNeJKNmTfqq2hNhn8LjSns0Vd
Al+ju5yP6PEbJU2/H3Uh7OlewERDm4PtalgKXVg+ZKMP7XYFcX+cH95lYYifqFQD
vpHhpy0DF18qm2nGSHCDLjpbjWtPWN2GHJbj45/boulwAKBcvyURBONcS268Y7zn
E6W2IUodirLm/+2JsKCQuuSUuIMmDO7pJnb5S4mcVvNsa2T9hZ9fslrrV/++ZkJN
xA4I7E/xFEvsrlQ7YaQeuwUtb82eetPkGC4cJ4jnyWebwwhaTXw5qLRAQ6iJ00h/
heJVnsL3tkTY/88tM6JlKgR0tlcWhzmfXzbXbTrpt5PAGTeXFuLmdjGQlM7FDxL5
hS3tM7wBiDfXqYVIUNMwx3SGDfAA/3BdE4NyWwTPXLb2BH1dEZZ/fYPkQATB+cF8
fJpbRGSr6KeeJ2ni/n4RWIlWcs6hfcAdjAvPa0hwlLpbbPBPG8IlkBg2bO5wz46w
LbVOT/ueGI++u3sLMgfXb1oAKKx4g+RmKTyis4rsp9qHqxNvBmSSry97QWJ0NaJQ
Z0BRddUZ+RSnsrvTWmMmBCWzD7kgCfkv7Pn2Iy4Ysqun9uePygibLqRtgr7LKuhU
ICNlxWqQ/OJ0uP/bvzszstaL6zljK/Vxm1bLHa3cTdiH9H7ey87WfIZIABgeMBV6
EipYDou3ArOo4rdXMkKrKGndCB8EHjg5MYR65GwTk/e2WavosbNdFEwUCqZVYSbH
LBimw+u0ZtPz4JVwiNAe7k0tFIaowZvg87v4AcE97D3/4ib33O/AYFHRjSPWABp0
3ymZ1vRKQYEb+CatcJCE8yNfM5FfLbgUbQUMldIarTryuil5NYucQblpGLH17w+C
r+hf4GdMZ++rW8Sssbr9uJpKqDMgGHVX4kNW8EXFMPzqzthsfoj+wTukJDU7YpRF
j8qzvPGeBgBLSxmaKtvdrZPZ95ZLYn40rmnzVvrTILp+pjRRlEglEDrxHX5ptURH
lbLJUvlprB89SgmmLPGh7iMDMXvOdX+WJxHIv6i/vxznv/H0SfwNCrFB4oJtg8GZ
uqnZCKFF+b/cID4o/mQWTN7YL9jdcz9c4itZ1u18ItuY1rrq6PB1fNQVxerLv4iv
0RO7mFmTavShpCmga7DDpaxnvk5Q3dLDa6OTQ4BN+pSpF1gg1F5Sq1giyoMg3jNy
eKsr4Q1U2vs4WjW0D+0I4GJ2wKL+3azsM5TAfLatsykcijCjbjag+9X4uL5iO4lL
Tj9FmTc2DV/OsAHkFob1QOgJtFJHyZj6cPPHo05vbnHbgntwCO0qIibIw33HGDTv
5jCrKm9v89JMRrn8YsiUdR8b/YcEmOEASkKaei/p0Eoz5ziDPOFZUHjIoabmg7o8
DzJxYW40Jmuvo+LwKOYuF5lsIp13kCLaLa4PqXE+fhYWCBaMjda4SBuU+UNa1KyS
/B3NjG90xcHWfke7cmCj6MH9VWMYoGbBVTbkKyfcx12L4idnLStDZNpHRTOBPf/f
Hmhh2iWPaXKQR80Dl0yigDgr3B8/l5RcQqdh2Y4BaG00ZqXz0MdFaq67HhgvTeny
3H2MOXTtO+Zn+fnNikGg9MlibccqSKswX5RuDiI8c3AEEeyAl+yP7IOay9A2VwyW
dwaG/jiwHtBwCmR6Ujos4IVodS6B2Owd9OI3NVDRQWkJnVoyW7iBevURfLGAn+Qz
BQYmrVMA33jUrY4pzvUFnHH4m+qXqt38zyJQQp/UhRB6jRfk4zNnI/kW23RMHeWV
E74cerjJ7k7GRO0O5GU2ut0qJmhISqrivO71fK/1Ccl7OGEm0hi9sHt+RW4zZlTr
8uMT9u1qeklpqVkz/aQ9XkOYY/XkuCycv4VmlHML2AEM0TcdbiThRUDb8DXGNAkm
R7OprqbBXxH4X/9SgMA0gIyIlgsgk6+L+dMEelgnhwzyClddH4r3Jqa7aMdv4+/5
KAY9z/2rzYU+o4t8ha/POdWroD9iyJ3irgyfgWpS1kXLLO/BQBOIo34sTgQjjFO8
97kDdtPn2sqUkETQQMUkuwkQZP9dCxGM81UWdU6ingJD+yhM0uBZvqyTfkgbltuA
dgjL1nl8LHrQdH575RTH9iShNdGhPBmH8hzJY6O4B+PXpNHTLAtLzmLY78uStNge
uftwnv9t9HUhbLiq7vZ5P2gOvcZh2MJilH6E76eJ6qdSPGzRFGUXhzYSb1LZZ4Ng
tZ/nXSLIveHez/QTMrjt68PUt118lJCnBE9lUlqX3q2TLeIJ0TAo9rEBEyYe7Jyg
NyuV9ls+fRsqTJe69Vo9uZLtWUhBI1Wdo4IVSFm4sFaKrVF4QO3h6/wJ0V39aewZ
TSUFGt69g7t5hISSA557OPBwQ4V+lB3ln1NFLHKXu0YDD5IFMEIAnBhrS5RPKBy3
bgNACDwATiCe461BxvhKzBD7s9C982dIogFJkhHo5NIwL/BLiBqMzmqZpVVIM2Pz
P03CcuCsYhdcUROXnZf7+BVBtKs2jWdoRvZ1A3JJ7Yn1gp9fazH4icmRFNZ3h1Uk
B757EP3TeGvjsIds/S6307uZf4kFruuCRE4jiNbR4czfPXX3v+e575GD7yiWV6uW
S+j6eD9Wzt4Q1t+PUzIQVPQaHt2Mlk853vuyfcYMdPDPtuDbq54sjZVuli/dn28d
NMJ9bdGRHyrpN5/AaNAzFQJ1+HbtF7Hdy2ve37rmfq+OTObpV/dUhWSnj30dmTKU
QxhPErzdApZbUp+M+jvWLR3kqCl9XsolUuAhBfUMw9FDNh5Gi3eWQioSr6i06IBY
IFeCf+c7dLOTEhkR0z66kILzz7Q6Lfp2z64Yg1poSH7EUoWiqDOF0LcvWHTWFn0A
a182/x4eTXWYdZWbgoMFYALjlw8raT3rGMSHFkyNfKLYb2c5U63PUTpVzAyOKxY0
/B9L6g0QlmyWXDRWj4QhdMVW4UsqO47A9QFEFY6fr3Y+LB12U8dySxT2mPWwceFr
d9gBE5d+2MJaEliasiSvwP43siY0X+shy7OIR+LDRsyv0keut4xEBfzSvYCy9h+y
yWHs048jJWj1sRMvBdKyl7E6g4QWbeN0HJvs2jQWOji2CCHDSzs8jhNxa3BUkgrH
EDKpOqlfP/RG5JPxHETo6r1NIdYEkTqcoi8AiZtitUrc3m8cR26n58yTSTMA097F
RjVS/22ZiFioZGM13FVLs+XiuReGbX7HXs6W5BEVPOrbkwBmXwlo+dzP5BSWrbCk
zuQdpN92l/b7lMDlCqPWr4KjHO7mZuFCI7AeiuUzKAo84s6N73/rS5cKQXH/Tyud
Tfg3HDCTBB2cChgJ6y/TQDQMNt5y39jxKf5UXTVxHf5EJ5l8UR1+PGq6zTTs7wOX
smdUFX9zOCKDSzGrb48tVZGg4UHz+kUf+mSt6n8qQVtQU3GRQSzSOywaORKb4Coj
/or/BdyXu/3NJ9yySG6Pl73Vf6kBH+g2mc8KGPLzckIpW83tR42m/hj53CBl5N6S
c6v0f6PR12/ItTUUBCd/jSYQNxkxy8fA2mOC1Wc/7hAR/urlb83vRnpRom3UIKTL
GAkpqfNvRTsGbYJV28lFJE8fBOpnLnao+JOLm/xwtkqBg9sO/FfSPJD80I4/+3U5
SA7rAfMKmumi3a7u7z0WVGyywcpuDHuZaSp9Xxxylf25jADt+jpXMSJWSvsHyl3x
1DvujtdEw76TLylGxTv5E5Xgk2dcB19b63loWEF8UuP91thpkzaNiHPYtJrKvXvE
ciZiyOCo5SthAoC+C4oqFKwNx0LGawkQ4zkTdFoxTsQKAMYupn5QH2V35R0+RLMG
yg+cdU4fk7wUUSybD9q5IRYYOsAsvigefWNecfHfB77elm5U6aOTJdmJv0k0F9m4
PLZoAtpEZSDH5gJisRBy4Ilwhuu9jZ/XZmI9kQH+jDkTIHqrxOSehmZZYrmzlk6z
VwkrGXtXzifKcglowdOW7kMGcZgWtXL8FmXSnEX6hSFrfy3TSsjzfxUlHuBxnDla
+9GWzF4EDFDwZqA+eotPU28OaHc+p2AOvtU4pmh2xEKl/i0NFM1Zg0e2agYlh3vC
wVukw/wHK/HkB5iM3eaQoFM7j6Qrn7QkZk5gtu8/oH1xIBew8aTNrzh1TwmaR5Hm
vF9LN0e8QaWNZ4WIShUl/xt+Jzp4mm3SmRWG/uqs8LqBEIODecslEAMk0tBViuQQ
`protect END_PROTECTED
