`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1ze4hvHbMQVTRRdm+I35Pj5YfvvsHQOfO8LqBd22W6n7xPo3tafrbT4TjpEE0gs0
s2q3xDjgPowX843M3QPGzTNmhXK8eQf9DIC+tjOhrEchRVMnpHkSHAmIz+DfKGMb
iLsWZahGeQfI8hvR3ggsmNE4tQf5cstRB4iZyKpHQSeAs055/MTj7cDkh7lZpEvd
No9TOa1UUJ4BTp0ylkBk2v4clXtb/1x962HxxP/mnAaTFyb6th3U5f0NmFf2kfYy
jcrgzGmNhCaOBNJrsey1EEBZ+VWHPGckqS9oS0+6Cxx9J0o8yQcJJCKJNxbHqqjI
mMUrIqzCM2bBvlBhxFooxkxw6UideAR8wcVuDr6fQrSn58etQuWROlfADYKOARuP
+KwEu5girZ2GfBZdKkLSgfX5z4fqPiuWtOc6Bxr/z3XeZc4+9264dE4qsQ/8oSMS
45eYSOVI4aoCSO0ju0Fuayh7CgQsxewq44z5hNepcyUjyQLDBfHrJ6uJh7hiJk3K
q0wFifRIELu1bJGh0Aijd1aOWJdzQh3T6DRQYT9iTrYXxK82ftquZegbbukBvuS2
3PklFUTY8d3strnMeFiB2dqBkV3LVCCs0IgD38363ax2Je0yjcCMUdNADO1GO+Nr
3leYGtaJfyqQej7gpF0hBVggFwy8vqlEL8h26EudyxHktQ6VrMO2+PFn8vhdt7Ub
c7Y7N+VU+FpzMPA1d5U75Kzhap8YxgBIFUz1+K9ZouFvHOE/7TqavG7DfIGmnlVF
Q+Xpzot4onx4rgjsuPV2ATvsP0s/EiGo7iSASYWIzPEu0ingkLdxpjnLtIus2TRv
ZCnSNo3V3gH3+3Eg9hh3of2xL3ljR6XH/LhM9R/vVRDT5SFURL2n3cW/fBDDtUhO
Yg39pUFbpIPzdCzeEjWjK2swC+iRVtdlgeh/BmYHu5QSxwHWykRvXD4rfESi1T5p
Y5Z0w1sfrLdTuttlnojKIkJd1QQj4Dbk7R6nFXu1B9wH5a8Pq0ykI0GEQhnWb0LA
Y7mtK+v3qh9ABVr0SA33dWziRtkFjdry5AstYJPPbcCpaeSdKFNbK4QBtiiwVTr4
J+ig4sr9CAqJ14+EPEi+Fvs2E+2EHU4L59zQzsZfZWkJPQbA7P7lgzlXz2lkeUTl
ZtBpJyk57krXiNAfphYOU7dOl4G+FH4VQTadyAIDXO7RHOX4aLkp0Ro7Xorv4JQB
NHsujrhPHIPnR9h1vSXouM82ppDuK7qv1z4DaYBpSKDMh8ZjGfVrZqjGFOeoI4yJ
`protect END_PROTECTED
