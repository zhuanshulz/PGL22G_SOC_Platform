`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZH/jBzoY/AmBaP0XPvtN+DrmQ9eqHcGuBg3Y1PQdWbjNA5yIJCDatvlpIkvS8gQa
Q95Vg2Xbr0TNkC8JbF5mUPTC1vRDVEnvbWU6Nx2NOrRPgDBjNdIVVC9cRifQ5HC5
0cFegnOAFIzUS+uPSMHRN6JAdsxS3grPpY2qk06cp6T20g+gfxRiV4OnjHOzDuxa
qpmJlBX4NQ/pW6wsdjsulgEMZeJMmxAT1MIqjrLrdOvuFaamxlVzpAOQpNGPgv/7
kvCcUA19nuJ9aeeFsni0r0XC5HUd66OQeUF1TGZvfpLHf0K8YEa8d+1vnvn9Wh5k
MnO2yeHSG+pYMuBPbUYOeLi+DH0F8ESIi8kRUKD/ByTYaCvNxibqVH+XTv98mcqG
lYxMT7RoSq0hG8m88YlZbgqKi0cWu1jA9yEKcXcSzV9J4464dFIgS19a7yOH+U3i
PifKCMXP5ikoPCwnePCZGQP+QVGbuDHe1+efXbPfvHz9iceDjsquwfLYABjg1TtN
TQPRxsM1rizn3mRf8YP2/HjEG5DFzwSh8+5/F18xCyz9FHOB4LiC0xwylA2YVMSs
0/XqINAudomZb+AqjQ+BfGl1YNCT0sXvWmPLXUEcy0yaGUB9/eyikmRd9PqE7PID
GsGcKYVb9EyUXF+Ie3KXAVkT+q29cBLYquZKCZgEPM+oTlS0w2N5vOcziEC8wJhR
H2k9Y3EUMp886XTRMfNMg+oZY1HepgIK9KfhGqVd7H0svf9oqq2RmNXa4hEJ48gv
nkvmOioFin3WrQ/kTrFl6vLATAB+pO3dZwaSNh4CH0qbvlWy3DqRfpyNkgPYizfy
/V0DqnM9sTzr5gHZ6Lk6HmH0FN3FGk/SPw3rs/yY5LcItsySjdHsOiCNnwpTt84x
m09NMGAp9t9peNzvIHgd7KHcbSQeNrj/dYvyXFJPxTU=
`protect END_PROTECTED
