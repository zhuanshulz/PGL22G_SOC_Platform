`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PzAw8zvlqZNQlTRIs4CUwjydupmaCApafEsHEDIp2puudz5I5tWYrWpoWcU5G/m1
ySuVP7Q/Uitt7qP5piT+TQz3GEdbuaPaveMJ9tbDumkY74/yqLEFJzxFEpXyaXfK
6kiS/lYGAp9YuL80/haxP4NjVnGY32LAq+K+/JDly4scz2lNA5esQng/JAFePpf+
naDS1WlowazNoExzJEIHNkspGwsH0aR1oWyjjv3PnZKctPj37tpc4A1Pus6IaSsp
sOruxVbeVyVb6Z20b6vsCCzY/UzPj90Tzm9kVEeUuaOzHRAiW4sp4cPHZbBEhIxd
JFBhWq3JERE0yqFDq+HJsoVr0IuCcYhpO9SUd6pKtCmWBdqE/ASR6DVcnl9mRk3j
H3ItrwlTbO3ZBFNqgy174+f6eD25b3KSXS93Js6QzdAGF0+Nsd0iNvG3h2IieT2S
Z2CbHAxq3uRJFGsQfFtigHYoUHs3mODs5x+bq+puOYTeXJXFhkOAq3sVx/vNkVhM
Ohp6mJWCv2/IMOY9+dWkEKTqaSeBmseatbCzu0Vdr5Rfvxr4iECgFjZ1O/3eVyLl
`protect END_PROTECTED
