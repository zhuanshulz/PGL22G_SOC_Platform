`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CODPQv/1Wp71/VYL8g82FATwJG0deAXn6d5SeEcrw5Ov/JneAw7s5kP3Ez2UUSix
7GXPXvAt7Yh0Ezr9Kpg0wR1aobeI3+gHmOf7OuynUfkbseBwqxL7PW3eTo+3+x8K
0DgvLnerybnSuL/FAjN0TLatuvtv9otXRQn+50qrTOOaEUbDG+rNW8ve2yCb9eSl
Fg92P0rI0xuOYH17XH+611PfW/cyfdq034J7Hjbe1vaecP89J0gyfnXc7Pc/2feF
0XnU2BwE2H2hFyaNTJZO7fBScPs83X2hsYgnztL8JJNmQ3wT3AsVpexbU9S3Fgbh
jgMDgYvFNhkZTKDMi8yMWeF3I+g8+TY7j7flTxAvRBp9RaHZNeooJkSoPs076G3h
YGB9NEV2/Zf4Iis/hMut8Q==
`protect END_PROTECTED
