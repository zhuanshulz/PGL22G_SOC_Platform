`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eoah+azLHj8NcEVCS9B7nXF2anOrdIoN240MOYQazJ7p2b3OewQEVJoOGivVvxnI
bbL9huHfY6IPqAdRBKKFibS2tg2+8iHH0+DbPPA7jjH93UEU+HltDWj8HEPqg+Ru
9g/zPdVDh2HUmRuuRFeAvutNTPe/z80kXxaB0ue88sOdDj/wyjtvVHuVdF6LM7Rm
LatXn89QBARchKllcRDYV4XkPHSmxZnrrjjNyCtuZHay+QEHnxh/fT5tAqTApe5r
YO7IaOT0Jc+0BlruyMQB3FuLbN+iFNCRx7NjPjHgvuBKaSVbpXPMVx4ejaRvSHs2
VopcGkofCHul7rzdUK/8WLQrT0LC84DipOVzZyAqSseLVYU+NviJosVd+YIv0D9B
HLsl1Gus0KeDJcwbR8KKd84TBswAwPxPhJ+QR2ghy0Vn5G6c7ZkUWceABZHaJ1tz
253SGbifN/nLGQFeLkT8M8583IfNX1PvTk6SSJCzADUD/Ks3DRplAo69tzOA0Yjl
h0evv3taYnNiDlgO0lWJ52kPygq+FqrJBQ6S5wvJftWYaM8/dUWAxkIEj4mo8Nsq
A+ngq3cVGsGthQ5Vxwt4nLhlk5ffQqxhzFj7WDvvp5iIW+UpIzzrbohKfx5iXrcO
lDhFtpC2d+JUxOsvspPx1/2xT7Vy3xCETc3bQBI7ufRNW2+9R4fC+vRSg4mFWsO/
rBCQfh2bJXUT63jKfbhyXOoXEMUXAkjaTeI4jFgOUC5nOWF6Er+QreWqb6DNJY0Y
u4k5ZWSfenPcuMmvQyzItvcyCJ+pTnfXhPEEp/mItWDH2k0lJCophZ8cYWP2OaJt
Rz+W284m4gduUPwZ+3/VPokqRZI3fhYYTwO8DrxHZPcrrDXBm6y0z2CJgEoJq88h
ALfrL90AHx6DCHbc4eXReXEsVizNFpZfotruCkb4LdnoHYqYcGtRI9WxwNf8Ajmm
dO+c8CaSUcW4Dk93/FDDSw2cs5qY09sOuWbCTzE0VGU3j9UXk0kMKN+cep5w6MFU
Lx897T3IgQsEYZ0ZL+32GMp4MAAUwv+znc2ZRDHcNSdVzumA6Nbrzbmo2IBeFkAa
QBUjAdEN6Rdy5JTBJUGQBTwnYq7VYh2EuNc2/KrZkh5pSsD9sDMsDv9YOdSyKaji
owZM/7UEfMoRg8rGFu+j0JUcUQK4bWDWMRPb1fRkCszmLDY5w6Oy0L6G//itQZJA
S3zdj5WGij5KzPReMnpGMh0432qSEOLpqd897peuNV4cWvsLKEtVGEtF8bkyuHi/
CdCH0nS/QfIuAzcUe+lth1D2iagujaAkPJ1S1P8BjNF8JtxBdP4c2LRl2YxczJ2y
r0KU9iJjZ82Zvfi6o74RQHgAIH9qaxKpQazCW8I4Ik3nQNuPyzeTFIdX9zm6aNlJ
2dv20fIyOGDTZ3c7e7i2jdIT3Jebh2xczlOu4XVCZNOio4XmK8G+EJVU8ZqGB6WX
aQ+8P0jAdCMEi0VvnjUswWsXrC/yW2HOUK4r250Ra6Ww+CI49I8eaeU9GhBvXOvp
U5OO16t2eRDDcFzPJ6p5VrL6pvvjhVgIcMdcjTumm4J935uajCpM5rBKTCxFV/PO
Ngi9HoMzW7Nx1XgAcRcobsmhFciDX+MesseJaFLC4Ll3K0v+iEfHBDxw/XPF97cV
npGBfW+3OEIP+DBGhaeC/4KXU6MWECZUVmIbv0wkSnbgAG0OVgOy3xYTFDw7PAe9
1rBHmnrfPEgaDFUS+tO4xzou1IjN2Oxvp+7CL/iixxtzibkxcQavpI3VTxW54fxE
JHxcuMnWKvdLAflrkxu9dHBKIIHsCGgCdv74CybAWYO2Sr8CHUd7k8DItQaL4q8w
dDB2Lz7tXWL53zz8mMaIhjUJJPL993d6yijfp1Z64FkdpSM8D95nOIzHAP5ykKJR
GiQxblr9doyFsVznNpmt0Zae5v52Jfz60xC6O7ERpoC1qJ8bQXu7GfWvDR9y+B0g
UAPhouGG+0HNjKUoXfQgz/l1TWFW5C2XSm4IH8rHkUUfVG17EpS+L3L55OXGeruQ
pf/4h8C9GD4KCgdDF088LPPxmrxIuijSPFC8+7oUXojw4UxpYHuj1VgHqyvbTv9n
zZp0C0bo6/2xfu0YgKWTMNaUuUd7bqITBeh0MTSLBiK3HWffp12pP0n3q2oZKU/R
+qFRWKiSeOvtcnK6/98RclLoulCvDbZJ2sqmjrwv+pP61nFWKErhxOEnVdt26IjH
gO8RcppuVh4Ti8yaMMc8++hBi8WHXpURjpskqke94pP/2ihseT8/5Lj1QCpNzv/Z
HLfGQj2X7xaU0Q/csrDM0muFaiGjEGt1OpLob+OJHqTF20rsWrsQ4pWRh8UGMkmV
XNPfnpHpVoIdPXo7a2DZOpMXSauPeoYoWrXuGr24/SLvh/tkHHsL+Z0Ab96p1fqM
VSyKVXt5i4iXFm1Nxr/0nSCCkXjHXMmNNJz62CIrWw8lpMZ0FquOPLSpM5MVm8Xy
xqplE38Mj/bDmJBzqM7Garl4WwA7Zit1I8PAxP6MOKxtwD64l2vNG/KIK0idr/7w
Ncrgqn7v0hcSKN9qFakHfyQ/DCRYJYTXud8cc2bAwDs9zB6mtSveQlZBzpgN1QBR
z95By8H74p4xrpw7WSoeDpqYfgl9NcWC8gGpjIYMuM5De+2yIxg8bf3q0+8DFiJR
mdIX7yUxXyImltj+WWkwgNEbKtmDGpPwSFteHSFj8DmSlJqy6Kfsn1EOi/v2nDza
eRfp9sbCaILhgcUlsRHcZbcjYwyptxk4MfIWPyJHwstdG6UL8lEh2LuTPP9Nj9tW
BnJAKHUJ1n/pYmvSVjmuAq/hBfVc3lfwognnybOSNmSWzm7F15aV0oCLkyFBaY5K
7OLIRjFEPg/zpeWwV63Vuw5tdZouAmlLknsdH2Au2XrmnGsnAMMEsuRcJcfW9gH7
2gxzrDf8nCOenKbo30dzz57poy2jhtmqQRw4Xe5RIP8hwDYeXyQCoTHJxb4XicY4
XBbB9CpyamC3uEw6ALJnoWcEaKTfdP9kuoOsAFoDlUtO2phrYu+SA0FpVAeF+6PX
xMHlKqetfzyYojzn5w1IGtP4zgUtCyfYpOoTsWKFLmP5h3aYXHgtQ91tUy1M0jwv
eHryAwar/xy6xNT3z9cFQL3C04RTlrjStedD9sEHqZVPCtunre4QGK5qC13YfBwr
S1dz36+vk7MD0+nHPRW2j6yjivX9xE/BxIeXPU2zOwomHQb+KWNR5p0ARF/7xIh9
L69MvkdpxIqCCg2hYufHfFj+6DaOx8tCSJpchPQwpocQQmQla4GMcewYPgw9Ywis
BiNY7H8hkiFlHjDcmzLiWsSFxEHLlRS6hrQFHMDTlH4DeUeRvcQUxuTodqAMN0nJ
eeutV/h2YOJVhtZtUA/9g8iFSS5f/W6RdzD4ZzQfequ+1L1TiQ/XWq+5iIK1vQle
j7XAbzgtnh33zNwRfMEKrp41MUcnEoDhqDVA0aM+J0W5JVGq9w+ZFjm1qYy7+JK8
Wxd6CF38JgrCuAI3YIHRYpqc62sp43yzzCxa48nWt3IsTbpsRYEWNw211WyzX3/F
hu4eiQFKB80uTz9ITAoU7UxJSSJCkgBWHz/BUfyEYh/n5rm0Jg6cKASTateiZ2wL
9eIdYkGERSNbvdVeewXgVZSW4I3gJxs6sO5NPpaOV8D/4XljoVwFR/2hPidIv1Cn
VvWtUyr/2FNKTI48v7shOoRHCcht7s07f3/yxJJWgUfKC3slH6F8YJYj3S3Y1Xz/
D+c0jbuvVAm5FA3b3cwC/90G84gRpfmSFieASXDMyoFX8m8AOg/VoZZfAhxvdc3F
MkvReWQmFHL4022tzTTw13z0AmIms8HnLLoUgpvc/31pAsjx17QL2lpmY2TpM9Xc
qcFN4aHn0+DC9z3SkCZWLMTrsc/uSU945mVBPTXAnhLRM8F5KOhu+Vksgh9UTBJV
LClXH8tWbi5Cl0VPXDciWK/BR2PbS4edaxVlic8n68/6r1VXimhwY/3uTpiQ2+th
lICseGM9todmm7T7ohRJJoPZ9IHyOR2P4UnHl8gld00j4jofUwd1jTvVRrip1e2D
1jOsYFcR790Dri2FzvDIdwDy3/wcTE21FhKzPa6i+za+wi294/YGubwEi2p8bfaf
f8rwa5FVin8BuRDQWBCjMGug7eXe/d8gBYaqU34rFY643ztZjBDwwEleTTGht6rO
GRKE8CTpHsQBuWYZONQZYQGUg0JSowKbpsYI+omk/MOSm2hdc/ZQ/PNickusRJ4g
oPDvDXP+lI5joPxWq05cZiGA5tIpeEkuW1rMAKXyjfaI5zYU8SJd/dV5oPzgqvVc
k/0wL+NI8krvRjPYcc66fNsf3m7XfLAobphC0DzCtGd1++egb19WS1IzB3xGV1q8
aOeqxSko4+qME1DmEINHQKWB3bLHxvQl7w9RYn3a++YGYAYYWChtxUJqe2xr3yKP
O+mwISxYgDeTbJ/VXm4yHdNW/fZN410BOgw/2wt1tNyftyrbbADuXa4sYvjN7lw4
EPcgUUBen3CUgFRTmbs5+CYfp4ELiRuxXaf1NFNQXS2u9EIVA/+YXheEMRNVKVw/
KNuu/rK0Z6oR1FowNZo8uoz3v5Fs93R5fBNPoXPvjodRa0tU466kVPxNW3w/lZE/
lvTKSZ7FodPQyxamAekrfcqS2w8ukXGr7EYxS4Eih0D0TWLpLA1x3/BvBcwDWDdH
jOdhaEIXjEIvBw9dH3gUdPzTijVYtCtTQgUTaRSe9uKf1tXXv8+ZqdT0z/H6AMHn
NjJPoCjcRZpjGLJyXY6F3Drr/wPQBSt6Sp0Ch89ZWxK0zMzIAhXbMp+TgtMEL3x5
sI47d5CMfa63WaD067vaRq3CjX/qTVt4Beh2HsVeln3kBCWFqqKmFKsaR3ODfuCU
0b2NnobuS9asI/WBpcNITvEC+W7W4EZ7gduTauT9SBhnzTkv4Sat8CbP1Z5Vy75h
I5Z/eLCtWa7NayCclgFHf38wAxy+IJdbZilpf6QAc2IaoU5NMZxq5sOjxT71c7q9
0YG8av/KVnQPnGHkf5Cac3FRF1rbQ3yeh63KTI4j4k7UKOW25hBFl69jJ2gsqW2D
ZlBOdrhzkzkULzYnq49HLqu9l0yjP25pEAYX9NR5HGVSPUObBcDgnU6oGBFSjiY0
sCdyDu5kNe72c1eRYDp3EM3j7NbzbWUjWxk5Y1S2YVkqhBKQ/1sm8DgK9IScfjRQ
ugmKkA+4B46ymGc7GAScokawQZc5xlaXgb7YK3gXuBK3HotTafNWwCF+pG5I5Qd5
cFu6YxDn186wxWaAZTxsoIsPtvwNSKc4hiKEo2mQQcJgQjNhQp/5i7rYtrWSQLmQ
R+iplj4hsJJ3t6TSOcARm7nLwERK7OjA9z0sQaE4GLvLD2010mJseDt3p6ILSr89
lgRAJ92g621LkdO3AZSLsvIv70DRIHwItxH2zkqRJWu2+BUOOX+EIwPnwuymeXV4
iHWoFQGddUDBuE02pGwroLClRGuVwAIh4KMfFyOKEgfH7Q6msd+e6c2E5uz9n5NI
0TpeNW1uuodlYYEfRJHGwgQh78LUj6Hxl1DEJmgEQiuMlgdo767O0GzFT8r18Go0
zQ8WvzWVip0IDuCda2sxtt8tNbicfgf4HJ32izZz0LCw9ajR1HzD04Bcb/3C0j0g
4f4g1H5KoTGX3Ub5eX81B2kC1w35CaoxZv8NMh4gjHKT1YGNvhstgawd49iNqbff
FU6Z8z/FUtqulifNa/AkG/W66rrjIzclyzXoXa215R5yyf4mNg0xAiDo2hmQieNK
qr4i3/AEUssinlMgXl0U5dkrUhTPSE5i4i44rKCuLx1C4iTs1W7yRYE5x7e3Tc6c
k6hEQD0sDvi2R936aRrGgbQITSkQmNlmnax6OB5ODI+tF40XQNEdXbLx8A8SKyQ8
Cqcb/OHk2jqmuHHd+P6mt0vFfipUF818jybEzintca6wlfWKCxCKjmOHsQmGNwhW
cdQEwvcACrm1KjXhJod5u6MQytlHZrj0d6BTo461qywMsssfvQ8PtLpJtCClfUR7
htXlOiiIFHl/+UIHECCargcSBsjP3oM+rRbtPcnvd6q2p3DmXBDFWqEqakfzrFW1
BPl1UIJRMVzbDgT73KUHFecRL/B1M2bawE8bhXqRe8ZGwRvdg8spPCbEQV6asji1
VQZinD+za+a4Ot5SFsz/i4awsgWZXxJ2cgZxwkZY0uezvuppKWSH5ypeOqpp/zDz
yla/Qx0hSRPP/g8oVe8oFyvl5Te3X50ld9hrGQpOfrPwnCVAGDrzH8YfpK25K+Yv
3cYjorj1/0DHoIOU7T0JslVrXi5wMLqrQ6xQcVvj9W5AKBwWJcUxml52QBSk0Em+
r86Fa4laOTJat5uQDXUpBr7SywkD/tSdjyd9S8uS9xKLJvZYn7bi8bdnzxcHtOqQ
HfLTzmzkHngP8hYOwugA62a63inhcoNQHsiwg8io9FDnIsewIRGzUQ/JZKwechJw
ujgAAlqCO4dUVLodKnGGoNYFi6y73Ije2syMKMKAnfZYEiIKWjXsOd9jBl9s/zMP
7b1IWtPlN10rmun7Ol2A7WiLA2qQVMoxfSpzG9PX9gT05zmP3iTNsYVj2daF71Hc
Ptdi5KAt8HAGQXyH2oj8qE/EdtiMR28udUJVPqrij86xDmA5cnww/TK+VAi6O/46
cLNuqRUKgLCZJGHf3rrdvUugoZTnkmti2333mdpyrdFukPtNRc8ado0JJZTN9JDy
fIrgKmiIYYweCVY33K2Rb/ciBMB7ZJByADkOaZstkxlbIojcXoROOdT188UT99QB
eK6TVgFDJ1Q/4IJey7XDt4TIpF3zXXvRWKhDBm/OUTCbVkrG8TGxBDdsc+3yDcfI
bQwrEqe38F+24Ej/CEY4yRs+OJSN/10F28IT0feJLVPD2Ln67M9ZTAQ8r57DGDpw
2FVr3aQ77lo45xUV20g49BUAB9wpgVAKDjsxkB0PsDzb+jnrsKjvpckarnmg6wMb
tXd6AZRSvhf8YDvTyTz7aMgvtyWWRsLkXfYsO89D8JFu/xQddv3BjCBJ/sgCaMTk
ilevKxUrV6e2ic2c4wk/rKnq8nXyHASG4vTWxzE+1MDuwKVh4YXlRxzkN9PLDUZv
1sLDYx1OPRu1ht4GLI/St6Z7Jbudx8wnYyMJPMU06g/O9PKwaouzNWe+yrEJNlhE
T6tTIGGmzgJvYkgGs/nBJ1cwSg8WQm+P4RpJxxGFI+Mpp7afgvR4N2UahNJXhZfu
u2lF1osnAGi/Lr7V1Cc5nz0EpoXESmoPQk3ARBDbr+DgjPfaI4nwnZoYQgGEtkVD
HOKzAJn76x4Gyk6mIeZKOQcIr7E2pBTEVjhMslEI673DUz06xUrIfhVUWaFsXw/s
5PB8geNs68an8i8SgbK9GC0I5RzYYPX3W6NsNasYOtwd2fPgqfzAQpQZXtKthzMQ
ktvCUDs0PiIBVY4yv9XDcy6B2k2nKYbcTSbBWLjWSI4BrVj9qXgp6OYrboRmnoXk
6eeLHfAlFp/yJ3ZEFySMYq/sEFWaSs6H4ePSk5X5N+/snzpQpCendjWyLgkpC1TR
XAdeJqGG20CVNu4TcHT+i16P0w7EsVySEXzK7llT1Nely56z8kRQBJsniS9ohKgc
Oi9gt24RSqL18/kQ3kFhpDLWxpqo9M9r1FIWyvFkfMYc3tQlT2R+TopkcOI8VRBH
HhYHhCiSQHFMlQagD667LQnztiNw9yCvN1D5J7wu821xxskCrUWQxHG+Xm7Pd/Cs
H4jR5++JTp4MeVIjnGetUQ9rJEwtgm1a2Tq5smUCi/ztyeVATLWJtVrxjjUHKs6/
ATyjyv1KKp1k8AhuoZ6mkDnENQ7o8lsI79QfjXa+UI8TJBjoq+9NrxghthvBNXkk
Aiy6zayn7RYlhExIC7zF9fuZkIOwS1QjfkWTV/dfW8ipbnI/WSl6kBftKLBt1Flo
vNMuh6XcpvyoJomAIAClQsdHMM0U7BuAENDg49rNwXKc/KyDYVF/B8G5Y1wt6Elh
AnccQ8K3ltzpcFqX6cXz7aOA/dlL5bqnqetOxSatDae5mmJ4Fy/32/go++orEfyt
pHaLrKkhu9NEY6JBNE3vGUMvTdQJwHHM7UprGQ8/rkZnB1JEF+X0zafo2lqdUS8a
3T+DpwamB5tRkbFQwndk1rNs7tDCvRJHC1snibRnTHgsphAhly/ZmKJkpANntd0I
wDAoWxl+P00+ZrViyzHRD35XWQEz4n4kGnUizb3xyQVqUB+NXCDxdSkhEp+dMVxG
ws4dAaPm1EXAcy6x9ZnR96zz6Y5+SUCacPZPpr+U83vUcy+umK5M8X3brTM2WiLv
jr7Si61QBJ0P0pjvOBNg1sz9RFH34WXzastNGLmFGxIFivkM5csPWvPfsTHAfxzo
boabc3rv3vmJvsYYPrD64bi6hB0ymhFwQmYX2KKbtkA6QOTK/e3fOpfpKFWMXd8C
NLcE2jChlcmQiWY43mmMrTKrIawY6DblDz6s0vAnTAna5CUG5zH/kJi6osWnyG5/
js27jKjK0Js1rBALjbI5eq+kbPbfQVDuowXrm4nsAz/1xQG/WENvKgKsDJovJUFY
eYZGh4C+8J8NKJT718Y3vwqL8AlHvDfu7aa4tG0mKRXd3nTIiOdMu5sP25neBt80
136xBqfaXoebZL3+gjH9wOdp451XyN4a1TGEExg42VerFoX9gf2BM3xEio3y/ZiE
Di7JVPHyErKyQ2uOtopbJS3YiMYdcTEPdaPATGbgJE3xhrMLropt1SA74LwpdRSl
8s23BNrtZHIuY2h8ZK1q2ozkUWHsBbTC5nfnpPsAu+wgPX4MSzj8wdQqPqdjtN16
heHXIdGzTzRzoxKJhLBSFaqS/7GwZDsWNo8GdPj3Ru+8x6SbjxNsltk+vODOJDRu
ZA2bI4ZMtu6RHIOmZDhggoTMy2Cp1mkbKl0WPW28AU3jZxDefOqUKJgojC7fqZ+p
8XsUKMQdLH8ooPyxJLruTyRW0zziSAPyTQKTyMfd8GYpjoo+BTRLTvjLFS2j67FR
fYL+1EI1bfB2jTYZd+5aFS6zUjIRYU6ii7MuT9cHzmJlvJHxQhLQ1ES2Y9ViVJjN
V0L3WepcWAfxVq4KT+JX8O02RmICPjuidSUKbntrk+e3BTAJ29YrFlzDJqIvmUKt
nCAfR0abSRZrWMwpIFv1egCN4OVzd9LvN2q8H3eECWczzuUELrs7P3aIkBi4h07q
66I0eAWuHL9vCa36E6OdRVu6a+1wz3KvqwlUoRwffiZ/AGKcYd6i4KQsS0AZOrBt
8pAOlb3PFJ95V3xG388GTOWoR5UBtoFKv3JUxsDOxGq1HSDxCDIsA/1qBdgyER4R
5YFX/PiBfSVswWxPuJsGPrtLOZP3qClfH0y1Jpoe4OYnx4iH8UsINzG9MxR//hBM
nKoTM4CLUUxCrhJcJBDUYdn/umr/5qTc+AIX18XlXuZlj4wgaEDy6gDJzwDoTiZN
T8vYZ4xwcoi5TZvkvWjxIsEXeevxmCq5s2steEmzRn+XKJ7AGqJnkTfVGHslpmiD
kM2vxF30swhxGR8clihaRty7fjzXd0+xSMIAyqSSXmMv6dvtCPEjyu+RMZhXMbTw
LFKyPjTcUIPEE/28ciA0bQ0VBjlfFsIwVblMfcqXy4AbWWeqSr39QfttLDdoojwa
kkutPLF/PNT5aAKL4q8lQmzko8jPGNJqpwEqmXCKId27ax+wwZ1QQkiJp3/k0rv7
H+0MZlsoh8zSO2kvBVf1r/x5z10N9SFPsCOh3yR88PJnWVdfY1PwV2vGFLADHAxp
fKHHCgckkcFxHCZK0P47oVDc9aeNQA8djIAMx2eMLI7MIEbkXC1MmB9UZ/yWfh2e
k9UJdqaXDJ/5ZYjuijj5ky9Krh+1VS1rpDZAPlB77To/E2Ymx6BCE6TRbgYU4QTt
OA+fE4p192STRxy6W11bbbe7fKCCU9dXvIXZXFDletycuRTQCCnQeyKbNtZPgayn
MGehXNSFxKSGLCYZWq9TxI6C0tnTQjxbSpv5Ujpc19IoD8BeP1X+x+yJhomNatHm
6+0sGo7dOyHHZRb6S7P3J23S4MPQKyc8HHKeQcuoFsNolskOlsv6mS7f6aAIwTIc
uPn985T2fKth2Ker0Op3r8EuGKCB5oSuuYHZo4Yc1QFBHaC+52DzMRkscDRG1sFl
FraJx1uhvEHiW0ig1Ir6yfFXbf+je8KkjKZJv/TGf2kiU2BbRH3QGDT3ILxaaldX
I83ElOYt36kmiNs4jRjasDpJcPrsGj7rs5XohHOXbFcKUscVjKZ059C/V7mjxNsD
GxGitaxdVCu5nu7WbmkIfw0BwpgZ+oUJWB/EttK+uzWJ1PcezlfqPt00fNMr/hMC
BxqTSJXaoo5+ATvTt7VRFho2F1uEJE5CnlfVjhaVftKvfWE06nVYef8oMIrLn0r3
78l0O+UeFd1uoKjkHmxja4Xz38E4WdOmKDf4cZ4cuzkGktg3jgETbXus+gRFpNa7
gWXfftUJhfrAP1U1CEewbrqnWxuuhenP2F6msuVeaUl5Zq5qFV44aQXOeV7fRPdn
hhlff4+3FfL7s1INu1Bl6B9YA0VMDP0v9KvLHhDT7quAdkPUvAdZg5v33i8disMo
usD4AX1dC+H6TaTYjwKRoWuQtQ+tfhI2nnjLMZFDwLMq+OMx3XlnpS+r8ABIW6Yp
X8DrEzV1dF1HZLNosJ+bKIoy4RbM6W2pN0Utt05O5I/0XIQEQgWjnwyRC75hYmmN
QIF3yCAMnGKfEuo890tDP/8d1jCWRN7XhCZ3EtOUmiq58nBsAqn/cVKEYj0/fds6
0YyclO2o/9GLa4kamOjUGV8IsqpldO1aA+Fz2sQkkjDw7x4adB12Vl58c+fT+Mg+
ahS4ZAKzkc4msMdU18YWQ7JtkMi3hxLObK+AM/r0wcyflmfvJij2NKG0DId/87KV
Qw/zh0HoRYjxsPL9+OkkQiVKHsGIUZ/GeFq4qML/cK3SdOvfK2e1ryimlYS+VJzo
wYMLpJk436dnF5vdKOS3gW0UzWirKGh8ymRPfCeYdmbmJZc7qGO8Guis8ku2xjuF
BTzqBlXIW5T6Zfdklfvu+QW0C8beeJGTVyA8jpnVRFeFBIZigXyykoFCV1+21jb/
3Y6yRNZvTA/ofXW8Xkaby9eMjgXhDfuRoUlCD3ALpIeF+LTQIkx/7MpYG2aelTVS
zd2GR0xQ7pIKh9uQSgSMLoZ+J0sU8Ks8Rm99U3Ug4wf6QERHHIs2Yldhdco60F0d
A0jpIUTTB6z938aOg2/v8S4zIz5sqKeky5TOcwPFGYWIG2e4Emmsjvl4rAaUmXPf
ZgI6Frt5DKcSv+GHd1Z06R81Gz/Y9N0JEscCoDOG3zATWPtXETB90wLsZUewUuPg
8jjgtYm/rzpD2Mg/keAlW7LtSxM25bxnlqBy7Ztk4891pF3AcyQTtYjSihFkvAad
1j8EASaPZpIhRE3/qxhkD3MsvoAtnDvHgIHeM1GFrf6XFi7lqtFuM7vmPFrWeyRo
LtSIywHKBS46ogoock00AMmj+COCcVqnm+lFLGLmgLuEm++XQb/hXRx91VxCLc53
nZo1SFaBbNwS4JcW3JWRDhTLH4+mM5XBkhsBebSdO3XQlyGD71GshXeJ/70PNIc5
AX0w4hNwAo+yyoWybYZCH/9GfFJG6M1p1z4F5Dc6DkDL1T8chzEYse2JcVzgtC/5
hC1dZnJaPstY+HG7ydjfYBSrGkuK0NM/rfRA7pI6hy0LPATJiT9cTPPmtsWEDfyd
X/pF6ShJ9K2a4lOCtTXIddJLeBETndsk6ldBM4qiFSdySwvHmfv5Bn7HX07ea4O5
25OgmZ186zM3mdIZ62E/68nq0/sgNtgb00owoQIeSfYTwrs8Z8uenDd+qUBeA9Ed
qKxPLyfTg9/2HKjuX+9J9MjwEQ72w4U8fb9N99rM+x4VleApCzq0Z+qhwLWyVDPb
m5/xhUDcXQOHgOrekWEIFw0GrcrOLJFP60D7ShGxJBh3pST0wGNUmektpqMz5XAH
UYTkwILUUnWokgjuhRVgeVLErucHKKKmWS1I/s66YYan4+5MttDQywL8qH9MPSXO
kbumPNuRQYTaJcZNDZn/YSBk7cPlKFv1UdtcQYT+ggZkCrmjObAnKqh5xKm9IbGH
br/0zM1nFJ9XXsFzPlSqM8KaBAV60B3a93z9o0AH2JHLhJpJOiyVD7cOlN0i2fwt
9GlQGsQyYmZE9FVgDYbqJVnIDsctg7JyKVxTdK8TaSd6iqJvdj8fsqohlcKK5DaK
Qv9RDOjWLTFHMNgxj897MS1Qu991fZERimC3yz1i0Z+MKRBZ9renq1r9ao2CgTJs
lG8gHkh9KJbbS/g6xAbf0MrnMoIAXIFNVGvagFT042awHlUVbm1xMxCESh+X4zo3
SgtlMWQIGZ80J3cxQ2y/1ulrIMV0dheaf4ikCGZnjMm/AwmmkDGWQ++XIzxnBDFA
q/LltOr2eUCAfi7bC3dESZTbmIUiqBPGBnb6oGXbYrbM65fapGr0ZbSpzHn11q/O
HN9JQL+pqEM0htBPI3HzIWhDk8QzYPaZXMG6UcJZHBVjB4q+P/PEDDE6QLxjovhw
btEhXZwOdmzukOobHIYYCDC9EpOvdCtPYR0rzndIrOpTwi4ngOGVdzkKhkty/67k
eNqIswO1pD/xDDoHr7ThY6cbOy4+n5zwXcspkdCrQzi4SzDst0bx4Az9T9t84MbW
g1cSaNLUHnTlfo9bP0ACyy7V19LLWKnkGEY4TwMy9PiAEkds0oYqpW/IuVutIyk5
KkE5N5kn3ugLGC9jECaWStyciDgOlfwqfoZTaWJoZAOlhmudFxwXgy87qoGdOLVZ
0TTkyxBENo58K2+00+k4o9gFto9IbD2L0EJ1VTaXrhMw/zbhqdqvwq5H4IhABJnl
ckhZSz+1DOQualna3+NxM87lqBwAWpkDvD3EUzycI0xrEK+yaV63rvudEirbkw7c
zYXtN6CQAG2+LkAOc1udkcemyNuHINrhIz/Pzkfv+w+oVseSKWis/IjEacrddG4A
5FjytXp0IdX7irzKZSaD/9OqKVDnaTvGF7V6u9D2UQat8CE+wkm3bxrcT8iwsn26
gM55RoLMJfWAtbH0D6jBpfhJ8BmWqtNPhluJVrmgdm4mTz96paEJJejV7xMDP7H5
GphEV3aqe72ktCr61jYEZqkPZ5GW06XdUQCo8bcu+tA=
`protect END_PROTECTED
