`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pJEG7iDyA7SBekoO2/H2BZNEgWNDrZ/KSzCdxi1ANRBvuU6J782fN9Jtlu72Jo9q
N+az4nTWt5wyt/ntJ+MOA/qE6R47CJYE8kYYgjYUbyudngdkeGq1l9GNkqUBwDv1
kau0ZsJWJ7uNNEm7tUT+aFJK3uAQop13rukXNyUM6jpEl31ZDVpA1XgFttS5LN1O
+pWGd8mYw0tCYzthYc0mxrAJhm1Xt8m4JW9OLhuDtqJDwVCqSvqncRauvBSUBJvN
WCljhg30riwpn95WKflXGmd8CQmggjdPx/K5ES4P00lQUKSlQQzdWGnT/gvzQI8j
eLUuxuIxZy0HDq5DhZMr1kBBGPKv5odVB/L8x8ZnSZqB0PHp4wXe01awmoaoNyLb
VYbLJOE1gjFAFQ0Z4uKlyrRvKE19nTDDLXP8grzVZjZe/otS1EoFQTyolhLAnCBs
0F9JKbtxG7DBVm6sTgRqiy0qGCb41LR/TfrxUv6npU+Qo/rUFe3WQLMScPov0jCi
XTvc5p+GF0FlHkEELUjcz6unrDzOP0L/Oua7Y/9ME/oXKLuA+PuuJMeQjy7Wi6yG
MG8SOtapgytb1pmv8IjiEatp9p++8tYYt414r8YadiQ=
`protect END_PROTECTED
