`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KSCCvMcSo5p+/Og0wgRWDCVT7EhWdKyQmvrc3YKEDI3kH7PpTKJ4u1+fsXyX9rd6
BI8gLca3wyYKaqbB5vNFWYjx2I7WDvy7+TtIpc2zhVPVAqQfQA27ByUTfjWLJ8p6
W8N+Kh87sUcjz/siH5JRS9sbzeTTL5zX0R2C1i5OVQILh6wAlOa3imxBM+tb35d1
bwSFC/qqpzleTIBoECBUVvogNWvYpOXmudd6s2Y2NSzSflp+MgagGKNYYEsIGngN
7kQW6QuKU9cH+Dqnrw8RbjGennzjyrke81Bdj0wuygaAFe/I8Zfz21hz0JR83uQw
rXz8I1RI8VXPHSdKSsJvZ8f/uQVzHnsYZn+MHepdrwSVyYpJXenjtZVX7voPlcZR
YcEbzuLjbNjisKHScCzxXUK+2O0U5VNvsmYemr9f823IUUFrJdpj28+VwM0Fs+Pv
ADxN8aDCu1squDwN2zoUGJAwDffidO6n0dtRkAvupO9lA26w4QkiwAAz9CnUzaMP
RJd6BGcAv5SFleuLd2Ioyw6n0oAgeDoJ7ajEq3aW7Qw1NsvAWFz0mOGkcR+6lUt8
gxABea1EL3K+iVwPEmXCR+rTXXnavHZaCKLILs2Bqc7gzcAAcHcpfx/Vn2GKuj6a
2U1NPsEP5vylENwD2tf65qQX0KdElliDgk7m168LrJFh3nNQUKpIAjzg+lyg7hwi
CHcgayvzzyqOBsl/kLScj3JbWDS753Ne6QPb3cB4x9jjLcxZB7MhIuHOncvIEUJa
M0tB88tj/vFvzj49kYdemJ+nBijXSoCvcrDK+uKwWPKa5YqmCXItJCm59FPRejy/
Qmd9KKXpP3cWaztfMFfGQqOWek2+/wMvDqtethajOFg6d3FjOmwBLB9qrjIy0yQv
PI7QFzNtr6OL+pVfhYRFqoGaML6kYLkdTwxz9aQwrKoYxIyE1BnTDN0q+bFrczfQ
CWVoQvxM0tJoqJBrjgJeNlm1Gd/HWkFzcoOwOWoqxe9sT6SI3TYbWL3aPv4vim/R
aiQEzUxpCSuSr+oFIqHSAwyLh6P+XL8UKD9ZxPk1p3ukTyTHqTwuUF6Ci7cdw3T4
ubjKKEX5FM57SorQHu/FVUjH6XglRnfLdGyJa/atdjhd193+vp2winuoEv6Mp4G1
R47aL3p5V8u6h/yF43pD32cNRr0SIdUKgWdTYch932DZeoOBpk28AINh0byDBAdM
6qOmjf07WvXp58xpUDbmoS2HQEUOGNtZXIUkyTbdJCytnW/H8KvRn5Yd6HNDd9CM
Jmg9cPIyDprUmAD/9gTbSVWe/hHVbTWTOqTqRIWqfbBtOkfyrph42EViBTTA8H1r
y6863UfzemBwtd0ZOy56JMfPDoXDZwqRfIBx+LCp96tf4WYN7xivZ7nj0RFAMtnH
9z9f2sPBSGNzIZD9Hxa4sD2d80MieedPt7AtipA/c3zm+ijs3n1wDfC0gVL06yv8
9P518J+t7EC/kzOrqqSixNIqdhNXAnZnxZSvkk1ylNq2RkKxdK/6DjXD2s4K6GBY
vCAn4jNFVRocpWMmc3OoekVYhzST4yi4ZDVcaFMvnaz86teGvnDajGsjYxw5dZyF
gXtlDlKYz1RbnXI+7vROuTpLTH0IW7yEuL6dm/m6jEKd77raBkAoSVIOt4ai6TPm
swToK5Oz4dJzmAtzVtsBrdqZNmQRjrdoMIaSCmw2EPcXi4MqwdkSVy8/7epeSGDp
rad5IuzSMVeQ+cbFUgct/4UTJdASxe51LP+LCjQ3z3RmacgS5TX6869Ysm6/dzmP
WtIgmnw/wg+D6v+NJpXkC9TBRk4eUuAubrgPsH4A/5yIj3Oll+8HK3BsCp5jUfpK
Oy1N5/0kAGvT5ulb2J2AXjWxnvX91yIHIV0/hF0pq/tJRrh+SINzX/pQ1l7hdl4R
3UY57zjbVag8lVyBFkXqIziEd+TrwjXI9NF6H3HA6swQnr06LYLImDhF0ZZcEnHa
RcffjwYVnNGKXTOScZCoqHWQrs2z7JIJIgJomTJKMT++t4Y5T4UcNSP6A4vxJxY9
IldS/1fGNk1NMB+vEq+pPkGaN4dOrh0OTPJdZU/js/Y9gZscNuNARVE3Oiby1ibl
7xCiKIGxjonbNR/1rrLlXve1rnCy6nXbKo17Nd3NFMPAc6RG9UvZZYoUcAVpXlsX
U0iklCFctaOiqS/+UeHEhlj+xMkJPF37Gwp7C/IUQxdXVeQWMSVR4sfbQxFJMYFm
N+avy6KpfVU5T+enX79IrO2R3Ry8WWUGDbU8KNdWqrKHzKRnPhK9/MRQFW2SaS2c
fVdPT+qMRbr+txgTt/1hLMLh+K+G3NefwjYCWJqpmBBMrky1i8jYG8cerCZ5p1TO
Ano7SUhRHfNaTYCO7drgxxMp41AvJWz/WofMovM5CgU=
`protect END_PROTECTED
