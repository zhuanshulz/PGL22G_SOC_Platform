`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FBj/K0mnNRXnsPCcbM1dMRtUg78Yi38DsCk4cWqEjkfmq2ZrtKcuiC8SCEFZU5IE
eNdaZJPYZ3ATbVh/rU5MJIYmGGFQldBJ/94KCrby9ZIcRlxcrBAjBOHt7nJRi61x
MlArgJxCSPN7AygbYYnDFvnwZGj8tLdb1reHJ/K8VQvCba3JVh2S8UfzRSyFoEXX
OSo3Dypec8uulNPjgLTQiDttnoW3URtXfZ+LqLivTxUWEn0vwUgbmn3y7ZLuT5N5
AXFuEPPRa4VX1mNS3kZD4XX9EZNg2ENlRox4A5UGoZxek4Nay8h05XvUO/ugX2AT
mxQaxZFCscNSX8cIqKA+TlyJJY91732525aDpTETeHo7As3v7EisrGHqM5bux2Ws
Rmp44lPhAM6wZt8FfmNuNmws+KxnltS6Kf+5GcJ2RkvjomYlf+CRHMGnOeVLdh4h
ISSjr3mVnYLxMeIzSN0bj4MRzsTY/HPuQcSvDSPWjoOl7/gG4wYdiJyEgsoFr6Az
tquBzk8HCUEGvl+5enxqOL2jxnrerruI9gR8b7Jj5TPVln0xQddMpP6L/fX9pBmd
/8/Sfxo/rjwuRXl0xcYBh2xoYfYWwssw8S/HrplJJNoCnGA6W/Q8bIo/rgpVwI9m
dT9rjfbKZ3RLGw6XQI+iVBunu8CqhhenTkYrf+wSc2mcJUJDMTlUI6qofRH0Uqwc
vISUQKK5DBIVXTD4XIFSFXF3MoNWgNcVv7g8sYefgTouxQZNxB2oZ8GMosJGZ94h
goxqFgPma+Bx2dxR5KLqZWVQsnhoaid8sY1B3ymHQtY=
`protect END_PROTECTED
