`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PPjnCvb2+m6fxfFUmkI+uLTAlH9WbjyN80H1MjEjkxT57+wIjH5nk+MN4dMNc/Ia
+cO1joJJ2XZmG4cuzltVp10qxe+SHWv+JomXi88XyXAdHN4dEfGFatbQWY3WNdUz
XzijM2mU5g2jq9Jt7vT+3zax7jdK86d0lsdTKTSWX3FJG5xodSExZKTi56AOYyt1
qD5uRy8qMyNjNs8x88QvJmz9ACGC+mYPmmtpWrpedJWYXT/oQvnK2GocLaHUMC88
JfVlPqG+NYClLD2b5hMB/r9tyeoioJ2uw72tEP7re18xJLS497Z1y18kvddtZTLU
59ByhnlC3zypVlnVFToAPojHB9nDrCqbdSCEY+9bmoSIfw3IPbMaX6PefzRDd2hH
dQi/0wOLLTkj527Pz2tWOLSCUIM+l5KvUYFVAdxs/sqbNtJmVsrHRFwVrogjAF/F
r42Adknpoa5AJcYaiQ2/WZqEDj/B6HXfDZaHm8O5O7vON9qN+aX6leV1sWcHYPNG
KAEbQ54oCzFC9ZMW+BfjZOMIxVmu2tywvEBVU32/M0u0U8VYSlNXm5NBx9zZQc/p
3KTqiy075OpdoTn8kErb/NNJ8KKFFz/gA7WNdhVcRnwKTx6+8RuHDqQIv5cHDn/W
jJVUPKtekqQvsLrpCO8aOhxwvHgtu4qwtlOsXQP7uYL+XgvzJQ75Oo+RnqhBvoin
pDlBrJF7BKnMXZ2NxGe7h2utVUZHMUsPyR51ybQgn+ImXs1f14jTMbSqTUcRcbpY
zmgCPgDBbVfFmDIdeD7ZcXFt4SUVAySfb7CrOOa1nF3o4vbJ5IqCBv/QTzuA7GP1
1R2Ot4zvjA0ByAoyXGKsPu/pbdC7+DYy+bD+csBuRVgccagX149JKCihfYZpZj3z
n1jIAfi9Y6vasU23u/AJz0Xw2JQeeJ62c1hiuFeJcd4MLI6Azt8bwLLhiV8OS5BJ
48eZQ6usCy9qrpsGdjOtRFQZ9lp3yesbfvU0DfSpRrjW0gLXyi3JppIzOuPmfMrO
JhLPvGjEo87PpgNlyAwR+4WYeI3GiVVi7TB76spd1F48haXX9gRFspG5r1jaEQkp
N9kUGyeJd07OJuvTGwY0PFIB67EFUNnCDdsqJTngKjexvzbkNHioS+NKp3Z1N7Qr
RAXaYYtHgZdgEK4CfYOMQn6MKcrNIl7pHgZxTifkF8GZLwjA7gXvgjzHeRnugusn
U+Q4OSItVrC0W6DTSCLo01m2vQpT8512alo+7kqtQU8/ZVRKfZkt6E1Z0wY45uqF
YkxvjPR8PYaNjZxvHXBa1sIuZ2oSnnHYhM0w8RUtArbgY1bI4KCayqkCmsgI/u55
rvxem5RcwHkIua18oSnHy3EtgEz+0C702R/SJjYZ829O/m75cdUqXtHNYIWhGqBR
DSSiSIdVCwNr0Ibkt4hM+I8f9jJZMjSVDOZmlQOG88azcDkh03HVxQe9YpSIX8y1
fWdlacDO6zPK1TIny1W8WxCB7QFz8Mcu1A8jHW9c2xZ/aR6yMzallZL9sYlG2VQB
PgeqykTVL/rY2+PQ7H56hYgBaZ4gxv1ImpKJ9hBGK2gMWUg3UJm+n70WxUKWar2y
meBlTLcdVgYV1JqoOY/2Qjt8tjOAbYJV/RLksCb6b5t3iRlwGtyN26iAdqNvRXgL
UnjgLtO88IN2d/O1cTGh3w2Cg6F70Lgy+Ls1b8gApQd++m82G6NEUo1ylJA6iXWV
iF2EliJxEy5zhWK+jSTPMq5wuR6/1x6qgaIkbMF9kA6JhpP8wLaGpPme32SHcxQy
cO5NPdo3SOkBhQPUWj7dtj7AZYTWx1rEBH0e1KoBTNA+uzgaa+hO07t85fkormS0
WUZZSy+d1PsOLsGzrRBgdOjbs+lgCJCNdb/qiTURKt1B+mT/Yu/GBAlnUaJhNU6F
aTaS76Z4yJ28NgBNeikzacHXwLMCThIe6HFAV/NkvVMM6rlI/46n06Z26lBcBTl0
1YMXlUxewCaJSAUWWrMPn+scrmz8lY9KKsWQEwkvoVzYWvWdtXZGk9emF/glDTvw
b8dJFAzCyJJlO2RA8k+iLWJuX0shPOOZvoLzaIZOHiDqshWAoWjmPBQKW+St4ory
GYUpHidTtt5HmyXtrlevdaHIz4/SFKWjp0H42zHOfoo8Bwj0QwsbSFaJVlJo3Ixy
7qWimvH3y9XVOgr0KpskQdaTP5VOJZpr1YEpXMHH2mG22l2glQiVMKZvKT1vW54v
Arye/2yykZVwwEHbIW3bIhnRLyk/Fgd3FvKb9suJRag3HJ7MmjVD2eaM/9PwIn/K
+0qvey3I6eK//LzK5dHj3AtGUzjbxosNu6pF6ENTyCnkiyfLnJw791iFnqmwii8G
PVEDQahBdnpDYixRlGJaIB7STFiBWzo4egWy1IXpl3AxZcZf4qUmmT4lHdhJOtt7
O1kC5+vZvKuxIBI+5DP/SEaxKOagvictayxHFtr7JKOwJKcXirVsWjt864Mpuo8Q
5/J8GR4hCistvXJ11fiMhThF3+GUTZU9rjZA/+6dCi6j18Dnb3/ULEeF3hDRzlKq
jfdhxnAH4DaCy6+sVKjKr9O9dFZZcPTbXn33hmCdS2BOlwnucRuXbFgeRX5ShS6o
TG55HXmhzROn/YeeEhY888GcK4ir+o8iJka701++2RQhVP0l5eIwaeM/LkQtE54z
hV9zxKwyLbek1erkLZxgrMIjoZXCnPQY/eJ+j/KUrFF4PSOKALFGfHvT+Sqd35ak
9yT87OAA2UXtvXlPX1SneVT6j7WXdEDSM6frkaP8DRTUBGfP0xLsqOHym3LNfvMj
EPeYCqpg6bY9Hwzq0UCuswJjQbfT/502DeALuaO8WS1ZLBhcOSJEVnx9NlGIO97t
PaR+bfTcGD0WV6ERgei/YwoV+Z87LpK/yHV0oMGtDEQoe60LhrQKY7xENJT2ES4q
`protect END_PROTECTED
