`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yq3BNC5joZmd1VQP3Jr2t57UFFHOo158UwK3vA9eyLBWLNEIovV2ELJeVVbdv7hs
mybq5HLfnVVxyyw+CJMFWoxhD6YEqot35uv6GRpdvJEaCP2/ZsDlIMFhJsHyJwHT
LbFjOWnZlC1+brwIBYMgy2+IVaLO9GXSHKZ/g/8bwEzJP2/V6M/W9aEKb1d9Ch3r
IWvr9qwsYGnZ5V2S8OFbxh03Lr3WPyOK7bzd+LDtk4VP44BVW0hezfp5uEMZ3266
WAyzaDw3QuTzOyfgPsGTozLP/TThZyInbimwc2vQn3nd0VWx2wVIdFW312w2OCyU
TcgxpMwxKcgKqYjBnO7rRrCI2+66FO59sS54yKEMQtgTq/bRvPc0hNHOQKzdSUGp
f9GnTvXyEq2GyhD0KlWikPE8cERZyc5Z/NdwQ4vjLH07Rf3/bhLpgNnMf5VJ7qRT
T4wL3lig9e+cxEaJP0xsTrOFaX1ElLDe3QR7JZCCGRjlg94UpkLVZaui9eJKvL/b
LXJmeDKwWRGEac5pu3NPMOwYF5lhZfzG9fjJViKCEaazPPNP8uVCe9HOTotHSG0W
pP8ybIrna0jStOUpd6SaQQ==
`protect END_PROTECTED
