`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jf3UGejHgK7fxjmZVrz096/ih37TnCCL21LtFPde9pCR27VcJYytwJ0arEAmEsTV
NnXsU8BGLU1a2OWb9J0QV0fXogmT5QYsuQvQWGJaRxKpvOhzIjntV2zW8sM9KJ99
UL0EZmR1KA+9oq2XfTFbZn4cZmiWPmtg/v9ynvdkoc6otLIdTVVMPVz9Yz/8HAvn
zgpmFQ3Qwvw3D80rwto63aiYvfL3yS8qG+BIQFrd0nggsRVJW2mPHj/tjpLkvgIN
Vo8BVtvEwSsPdQMJMHb0H/7D+OXnxFzfjuwEPn17cwn/vU6IxVh7zpOkBUqA2VfP
9E3Mhg771mMGIQtRq4mPs2VTLzoUoqxlsGhHHh1SuvIrFEcH0w/wKZu6vVvRDsZj
qahDP+Xru23JpPVtNdeaaeAL3EcQyQZh3ZHhp/B4g4cRyIAP1dRrT59kIL3dgxpf
zhrsV27Kkd8GcPYVGsgCMUwk6nJjKptzR5zgQtUVwEerN8/3Rge6tG5eKE/JaZTj
0D4fRyB+4vrSFFYFQtTh6g==
`protect END_PROTECTED
