`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vRkO9mqG6lh4VZR/f+/9vK80OLq1hqaMQGi039GqU/Mif8bIJLe32MjDZkXj1uFN
GqciMPV2Jj3FgcCqbBmrIH5k+JVcfKHA5OhH5YnMv+j8FXvrrChq0cJpkzZziDDC
JHS6AGujmVL4B9YE47OE5QOeTo8arkGl9DmKcx5QIHsKGxABAns8rKu8Z3GeohPV
Zmc/TsjQAZoADmUp3zinB/0KHciYzGR7tomPX1xxmIlMqdp0JkHzeJsbSMTD3+vm
X6fazceSI9o05BMu++3Pat+2RcgiRqlDBylGTJGmbX09LuO7wscImP7xhT3sdooR
Rp2boYuezNXCCK7m4e84vrdlOBiBsQQ9iLNxRdpuEbQvsUFp59SY+3dvQMAFSjNh
Ms8N135mSv+jadbDJ4I1FYKuaspZg5Q0Mjt1tyM8F8s=
`protect END_PROTECTED
