`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ul+sxCYMRNMoyrShC/Ji+k2AGzPL0H0cPEwDaUhOx0aZqNkFel5G5KOwWa73+MUO
NXVrZTFIIiFeTQPO7+dx9LAPkq2/c+4z0qsNJN74HG/Ue9EB8gCUft62Q+zzkORo
IrlSG4iKJA8U94ZwbPLXx1skR1eiAkAsgLBG3P8PFG4thabiAsVXTo9MD/HoCRto
8qI6oCGl6+w2XKEEkFz7URFbxTymPNvxlE17YVjcC8hW1yE0OSk4A9uFZFWdqCJR
DoIPnkFf3bNJ4R06l7uD+ufQhnAV0Ehm0JpRTM3cl/GF1C2xhUSpZAbwjvA9zJVx
5ZVPmJPotyVFxunb9dB9vTqDibRiNqTXXA8GAs07310CkwJi1fvbGqdQqk+FJ++E
40qEDu3stn5Pvnzg8sURHQ==
`protect END_PROTECTED
