`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cmWIVO/hSvhV6Nl6MGxJaS+CiU085y03TRanEE0Xv1DudKmK8WDp/CTK3cqrP6Bd
simT5cmbuzU5sB3rDPOSdeF0nljH/c6ynaogCnD2UQW22UQF9NkTGb+/+KcjCcyG
Ja1TM4rZNRvbgS/mSTZwtBTpfAa0BTb/uEXZca3U5HHR/4mKRpu2sNiRBwGBAsTH
3BpEEzehq9Xa2btaFWi8aQq7gaAAbY1q45VeSqH0NjpLp+dXzvKAFjfH3aO3bRqi
bU1bLrLBVk5w/ow6C+dQrojT7nCJBlq/2RGVlf0O6jzInx6/EMn5iHM/rs3rdvWy
PBowJLqLcaP7TWtzhYdBmX2OSLyNtnFOF1KwYnbU+wernLXgvCYKBfQX4hhvNO2S
QX5mzg/17BiF4fMXD8mZ3ggxiCJFDtpmzTLO3UcjyEkmC8Rd3blE3Pezynsn8aZn
rUOvvs+lJP+DUssT8AGPgO85N7dhZMLtAJnymiVWfOikt/qKdaGxOS5eEjU6DGdG
mOsHOtKMfay4n6yXXQK7+Cas6Hgvxr6PeIZGV2fF82WqUUhUBRSmA+lzmL5WZ+/G
HjPw/DhxNeWyTGES16s6Tg==
`protect END_PROTECTED
