`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G028IZW9/8+bl9Ls7wbuRy01FBRISb01JjEZj/dwaypwBWfvNanUt0PLFl+McRDY
DmC23DKx1pTO07i1MuwAZ0xr0zENIz14KRBwh8JsxBl3T3swTfSabnTvw7BFIaxr
R2yEJYZzV1aeuuD/nX8MzvFjht3gOZbbaMwOP+lWfhduiBzrVWEy5OunQcjsizFQ
wb8QAszyD03ZF3EZbLUmsrbQTwKK488Wd8EZb6m2VJFQIH7jUNgRJDX6y9lEZStH
BOnpiEnn22wgsc+f/MJiou8ux66EkbXbwH2zlI9f0qtD/mdI6fY3ffSyxJI9WVEU
AzBIdJiMpEOa7+eBXXkEzifEzowLAtLBwleVWLPh4jdCtotKTlD94mLJocFP9LhF
Esx9M76g6JRxGHe44JlAgL1pCmSerGOnKUmkDRElxxaxCvMR1OpVWJ0Iv3gAyHyv
tiOzK/H7ndkmP6oz4WfJgyDidVgLXHGfS+WQ2rUvXJn1ScG0XU5lrFJVAcYgWRyf
DWDu+3Y68meRG1hAN24H0SuksgsoF3TY+wQ2sE8EDvPNon5iAl6YW4uersmcNjyr
Xlxotj9/x641DOh2hyvm3HQCbzd1L8g3wEJUpVD05sKdW3neOt783W+BHoQvwOoI
0GiVTeRN/gfWNFDS4isbjxaDFIXeDuKXZBFNGToKaZ30WFp8LdNJN4dnoXyeGzNh
YojJciWMucyG0DRblePAdx7WH5yT9A0myQH7NuceidpPnzvzYe30petEW5tZemHQ
8dmVVXFIuzMLTZjoOUsqGcJIZEmzL47o7XmXrLq9vQj9oeBx3umkSCZUl+v0paEk
suN5G1Jv5wCN+crPK+0yTM8sPnSfa/nOCLaj0jNTj5rmiwjl/tHwXWAv3h93SR2y
1xjat9wALr8BN/qEIO2JZbSvHTlMsG+y+sPrf6oq26N2dXqYebDYufNO0gHmpOqD
xh//+spBGrVUIrZLfi0U1HwShFptWTMu/fYApl6gthBeCdUC25gZ2YdGd2YgO9m4
nfWCntuiZScFjbUcoIiQ1GX7ftUm+H7hzwUrqW3zL7K/OTW37igWO0dtpKbmaagE
hL/JEPVp6jTskFsiFlnDLDefgQrpxseIjDOQaJDdpr5zvYgy4l+lnBmRZFcM4ewg
30FzYNEoTIK+oFnquXGlYCxSWDna9lTsU0i/126cHom+mV0HTtemyVDDB44yI/nc
A+a1CWVev16v51t0FnoaO3k+DIdrDdcS1tT6UPRn+ISnT/VCLJxDWqBbWQncmkTC
QTVt/jJM8a+2qarJxXMzKukcEXelnVWJHwUJHhDPso+Np58rb/imzQA+mYB3jsxJ
21r9HyPuu/YSLkWTwDg3QIPpmpS0Y55I2fAf+BQ/ichKYywyFVPqun3TTsjblEBr
ZbBJCNc7xg08RFwR60BP5jZGPbBWKCrjKT8YWxDmdViMJtQwSns5++0g6h8G1tQv
LjUuIN3T53ZX+4WNsno5oqXogYQ/5gmasMxxYNeUjtme3HgESw2uU13QDLd10wJJ
z5KmcIi+fo5MtVx55Ar1honos2Ekqgl65JG8iM64raZjFIfQCL2pmBZqzFsoUREQ
3tMwYvVp+BX00xgxXYKY7gKPr2Vk3J6G0qtGfRuGrayQRJcENGbyw5dBu7dDDdXA
hsIIbXyqf0/bucxsplu9yk/rhmqFARutr2aUZEMF4c60SS+dcdjhbg/h+szBre6V
YNaQNSYd2wSNKhzRoM3ff+CzxNAaHRn/IBS/wVvzwjZZjjh4KrhURLsKySAXLzbo
/6qgJNzADVM9TLiaJv3uCYMtExNY5AeiRScukauRq6K9toFzAGzlsXZ8ce1MMNrD
iK9g8yFnmrs62kijfRDByDeASQJSUILafr8LiUz016u0lou0xqvk2Ecby9pJt3Iy
WuQ4WUZobxYO3sS7BsFuz5vgU5ZCi0TaE7dbq2e05sqLiTQIO/xmcbV+6qEa9AUC
5u6Gm6v/ZWLMy4ebEvTCL+3MAOk6n8F81zIUETGSR3wgOb8iZFCx3RymU0tIzT3K
XvGS2Q6ymxCey2XqP343svZ52WMp7GLgitmnLf02cBjMCbEw5LQEdE1e8lQGNHFh
`protect END_PROTECTED
