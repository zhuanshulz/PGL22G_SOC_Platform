`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0mmjQFdz7uJCQSaQ2L5+VTi8BlBeK2oIm1OK2ch3p2RT55JbgMIjgGo5NgZBEwgi
HRpvNI0/NyeGaYZqbJuZvfnIiXBIrhzRWvCccfbzEKJZ+SdkG5Lr66XAJF3SlSdk
YVBREoX0dFRs2o8q24zV1LNhs5JMORxY8vb6YuDO1zNJ6GHCRD6bYrbNnqpPjXBQ
/HKzaUJao1hY6aFtHo3LGnQ6FkrewXEsmRoNY+3XRqp8dNweOd74MM5YWTYtsjIY
eyB/pvYdbKVqyDvFbTiLdwj6Upn47J88yWCj9QmAMNKxcnXAd7vDlNkUYi3sQnLi
AE9Y39RsJ1KWOw844OFt0wsdLrdFZhrZvlDlvDPm6zj8uMR51BYXUcF93/LObHNu
K9uhMlSPSNnyLvtTl/YhEp2hCQcu/ivxHOLyER+Qdp6WJYe0Y7EGAcHfNizj74u4
Fy6PIooLcnP/dlKexLAatnA+uoYNLBodG6gXjdQo7Rda+ggMVCAzP71cAjYE2h7a
Ze5wK67dzMgcOF3e+FU6U+7WAIHyfpAt/A5zOISNlEUR3gm58jgDruIgFm5K/PUl
SIA4udvJ9Y0oTVhZ4fM3agP37ErluR8XiOSMEsN8mGRCEO/4+79IokdekYXd+YI2
ZobrIu2C4gbooBnUjqJ1eot2otwLS5V83FIvL6SzPyAQlsU66nTc6fTOFRALFHd6
8P+aLrLUtNefmfksarOJarfCCJbCoYg+4b/MrfSH7j3Uo5cHR47Mk+OT6Q56XPyJ
NnmJuIEwNEw2+RzrBycRq/yqEVUm23LM3R3qCvzcYOZ/PT/0kHDdTQPD7MDx/OKA
lkWPHhE9CxrWU7k/lXjGdYAiDho3Tmw4foik5JT2aPfStF2E3gPt6G6IeqsX9/8E
oSWNkcTYhRG5aXNvq4mwiLSrouKtBx8nNVxFj2H3D1sL2XnrvFI1KbB1PLerarPg
Gf4SOWKab/t2FPeD0fyHoUeP9VqokaJ+20hTRpvKwUG7ZXaIw9+Sg2c6QMG/+LYX
nrWWbR0yp2t+w2xfhNXS3BaC5zqX08cN9wEpG45Mp6++EGF9kIxwMJiuPIGjWFjE
lecQNXx1y/9tUCyXXSK//agOFcKRxAgrF6f6yrZW0LmcwP0yIq+r04zox2pTjlKD
TnTtTfOF19YNiJB11p2D/RYc7mqMlslE3vIGQyoKo3rvSZFSffDxDfU8+BeqHU6H
oqyksHFHNahRwEquu7iw8k9GcNprALdVq91/+AR6lLyUnx92TwT3Rz8MdWCUV+6U
jzO2YLcrPpnSAT3emXObVtiWk121eLtl1FS8LBSZ3V/zO6RTlQEtq5RbaiFrOJ/0
`protect END_PROTECTED
