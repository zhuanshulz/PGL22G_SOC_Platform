`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iZYtox8YIRtmSe2IYcv6bmO2Je3QYqBLLy714+ePCBZogG6q/tL8z4edxkPggIj8
+fgLMOpedtQ7oGAbLBAmr0dUw2/ivuOcZmXbpzIrZicM+SpZC8edXLFSaQl5+m05
x5V+6l/zNIL/4n0W19DPRoV96EeYEI574yoz4Ip3fOR8QmCfRcvg0ARK6WhDoiIC
LCJVmSbbAQfEkjZ546pHreOMwcUOHqbT1PT/KHIou/S7l6xxWvf9IiRaAIndPLcl
h7KUdiXxJ354lD8RjK6UUhkDmOy3Lu5i9Cl8gbIwdbjorvMSn2LQ9/mkOuN5VNvX
CKCb/4/NnkDCQXzk5B73pz+BYge/09vxABzCfyrGZIHrx1YvrNvjjo6DmZ81Ah0p
MdcYmUWIHi/WYilJCM9UhoAU3SLJAJC6NVTr8X+0JmoJ1Dee1fCZHWccUX86udKb
l9pbrdMS4IE8V2idjmDwCOl+Y84fDV/ShaCtTNnwoDiknNma9vFU6NmwBCw2MvA9
Ijhy5H2lkbueP6keMcQcvIXIJdkAY+yh7ebwCXRdaurpTqGgDOSQxtGAgPQy450l
JY0Ln51HCT7NDSZr5Fj8uhtVth+83ZTTdI02V5+e6CZk5zULvNnHZARv6c2g7AGn
pD3eAXFoO99Fv72Z/amFgXGTePQOOWYK5I4OQVRDSbBPkOhoyrQ1uVp7A/Jtkfwg
o/IlOStUmpvNDy1P9HP2CVnAldqzGlQ215QO4wGdlLhPkcZmSpcU5UAUu4l5MEyf
x6bGj2yNomCMZahJwFb42J+1Q2vs+Ghc7d31ZhcvRv3znO68T4R5KRa44Q+o2hT1
KaoR1uuOw/p4g6OdGj8a4TiO8wdb3AqHhJ/9jJuK+kvRhaElw2ANxCZlR3GakALL
ul0jmKFI634yIjtKhTB1SbIZOLJYeraaP3/pkGXuRv1WOQMtQv+SxNQbwRD3k93A
PIODRZf2IMEb7M8O1jmy2f0vO6w+ag0DZjV1hxQFUV40GcDGmHdlFae3u4ECPURX
`protect END_PROTECTED
