`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B1g+0e61UIeDuImFdoIsWLGwsM6mKQcL6F5VCFldJqNYih7Vwd1kxw0eN8uFvhXJ
hgiwSCjhTZ3OES99yERghBdRM/ES8/lo50wUnnbretw0URtCn0BO/k2g0WkIbVDW
P3P24doY1pLBbAUF5aWvqZpO4D/oteNfuah+ftIo6+bkd0BYPbWoLY3pZaWu6PKo
+xdQYaZkVMPP5ovkM/21l79pkKOALXH4EhMH7w4uuDQ0AFOVr5Xg5H1Cwa/b7mtE
kRK4tarySyZh8b4k0ZpKOI6+CpRRAEwi/pfnVayKrCOYtCluxQPNu5IfpRTHLQpY
R7NCv3uQmw7mzBhScy27fV11GXzuptSj4LP5KJRYLXt+oWX7f78LdA1QyuFdc/Fo
2uqrmAgcqsqUHx2OMdgDxiML4E4OYt+8qgg5k/L3vp2ID+B0CfvpaJbkdySul8Pu
dKs7Ayv7QHOsqb0LM70Obd7YasB40HJIoYqxvpY/5S3UvIUE7AQXkrepHAoPX2T8
7o1+uIMkpZQZlhaojzPC1XxiHnVbsplOymqyGlNrIp7pZeVsg2mPrpAfd+gQWQ6o
a4F/X1bJ6RHMbZnfqeI7AnMh3CBJUKZ/v+/VM8sii/bk6hNtwaqtHoFe/+9m2Fhl
2lHFA4warqoJPJsMTgS+mVl71Lo10aEXiPD4fVwhQZLIKVdO0h/stQeSV3XO8mCR
fXJ7mGan9blA95DGkS4lMegKi/MxUn7IM/OtMhA/XbMqLHw1FR/THdQnpM3+b+mQ
pYp0I7qzHS71hsHH5ld/FyI+4/So8d0/O8kMHkXVmVQYXZs2TtX/yYbullyw1oma
gQDNna55QWlGOzRwhTOOBcUDsp9+4dy9V54suXJVLJm0qt+asO+xmfwWgqihEc6S
cp/0vy5v5cSSh//E1gDU8ztZ1C1OdncqpuaOLEZbLxGIRK3R+aoAFNVyK2FV6pzt
/2s7aJRouKnf5udfm0ejRnoIgC550MUvhsjHCXmItlZ2kL3sC25EpbdDiOLwvHRj
Wa/6ateqWdfJiU1DQIWfv75KzM3Mc5n8JEwSlnkij4ot7C5dg0aJ11RqYtwwCPtu
lVpWWJBMU04QAsXvDw/40xvOHOo8KjuJUTi2eSJgfPKPfZGzB2rpgczVguD2gTCT
0sNCGLHQ9EcT5A1kTs9zIJsTITOYgs4vKVvalxrZ7Wg+YMlSvgofuRG/nu+IZqZa
4GSwzFX9X04O3w/s5h9xWTdBkbwdRXwPd0onQGQ996lp7VA7O+GIonrUQbTlWzaX
glTEMKdpwyaAzQKgb9c6xi5eCxAT4GDhy3aOB71yP91zVeW750IV0uPL9vWmjX24
bfDT7fi23oPVbuSlepefDX+/7lmKubO1oi33rqTmt7Jb22rgJuz6wT5td9qvtCDN
+Y2vRDxIivvlTWMbk37afNX8K6WK3oM+UIYNGuISR96CfiP8di346Y4I1TqsJUXB
HIslh7rg72iovfzfpGX/C+oJjqjH/LefUHW0mhnwmZqU2FEInmDRLlr+YcZgu1w3
5up/1iXB6r1asp1IodszFj8UiHxEB4qAJCbHdTdeNIom88/MERDqywU9GJ4YQ3Sh
65b3OC9A2ht9lurIB5O8jgTH646aeHDkhzBKWhS5zpdCQHAsre29JtPhu2h1Bbin
1/dY3GMtrmiVvKrTQ5bTcwyG0/UQkJeKBpmSqnx0QZGW+9Z3I1hvhoULas06utoM
PGcJh+Y7KZ4cPE95SY3KtxyuJpMzdrVlfOlbpcBdZtGrFyPXt4+1aOSz7yRs/AXD
r0a1wvBfP7eI3bAWSVF5O5dDZ11iiUhndOc/dEeiyMMxUwV4uINGHhKriQgE+8Le
oU402j3pshV6lTHxHrF4qs2t+ZBMqU17ok5kMYJM4HMFwl6LrOYxNkgT0FR7C9HE
VNKJFLJEm52m7c1JwBFsQcbAfAPtlrhKL1jtS2Xm6I30IAX3uO8F6Rrm/ON216HI
mR7n/EiKYkg5k+VirRDuI4fxDu/v7/ZrdhupFXbOMdcU/KlJwkDwAmBQCnIYIk3O
gvTCE/awFAdt5p8LkNYd9BWFJ2RZ+gzHiE2zmyIahh94G8g2qPTQud+7WMBHuV7y
adBu6ZEoAqlaaMKN/sctrL3aHgIY9h9S25AkrddPIXXiki+1TY+D9jgnR3yae8YF
l4D9u5RN2800iAR3CrrqBjQ7bqfsjjxIdLgKedby4FL/9wFDGvoblZRWGjWSg8s+
V4nVbAghRGyKrzPEs/iqkufdeQiLtjvpSdg5vO1mjJbv357LqSIntXG//hLIgGq2
jaESrj++yeoYiEnqAp3MauUpJSHsbu300HEcH4QIEMLyADQfk5s0aF3+jlv3fvOU
HdaOmcFpsnafpvkAqIlWKw/Wu5iXIv47JdFqL+gVL1raCkO11JkQ6BEI+8SJ1Lbb
vlGqh5lI+qFTcQNJYgmEyAoBnzeIOZiZlW6M1L1hA3VOpXamrhHS834yDab8jmHv
zEH0Xe4NfyFtYRWA5kLXCE3+sVcfEfOhDg5Gk51JJuXhNgKSPTXuXSaHXFSRQ0Y2
LjFlNhGGQthO96ft8qsaetYTjUSAWShOdWQeRWvMh7Qoct+zS1og/btYUuyvzWqV
lykrRRUY4ymen0c/r+HTDYP2kyTbMFRT0Q/X/tZ4ftnRnBCx+nGP5IJnV3bVdiXS
TnMFaLYV04yV4Kg1ehgINS2WwQpxMBbGGLZaJV1FfOiXpEvjkRgFOkgEzOyHel3r
wBiw/ZJL59mTM8tuRcxpGfAn5xlLcM9d2micrcLP9nyugc0w9rWlKrS7rbSczb/T
H8Xcz5zvYpV1j2Wjnhe7jqRkhJMhYdn2vs0RFVXX1odo61hSgJNUCS+1gOthWI/7
PuVnZzP0jQi0epfKZLDQmQN6Kom9FqogAHTonRm9+yThGYutV3557w2b0oQOoEoS
7soNu3ZhE/3MDypdj3fhyHk+Q712SflZXM2eSnJj6QBKFqKqw/vaAnoBUEqImqUg
HKr4H6WsWVUz8NwZ4hRXvD3oi216c8NgqpCXCErdbynHLKc3tS3fMKnB7a4WWHiv
g2QS6qX3FUwdOFvIbkSy4AzWnR3vEJUW5mmErPQV+3kzJsEDvcJyBc5debczNn3B
Q2wyxGSCUvAN11mjL2riVqg7f5UCJioHyk2p0yg+YZAqKTiXtZgfPBB8m5flp3tr
yjj/7mXNK614giamuaihEYovtlpn0WmJ8/pRoZ4r5an2PbElTWMZ6IJZDaKyU9wV
PoAFL4NVOaEVsOgVbcw2oA2Rn9o0bi6Y4VW++LnoT0w=
`protect END_PROTECTED
