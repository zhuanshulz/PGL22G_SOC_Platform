`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EGGrlSnpyDnFkfQyzsoCG155micg05mHgW6xXr1C9h9mLXsnjGNtp7HqJ97CDhpu
mBvMC2icZCM1LP7+4YEYDbnPC/K7L05T0mUw/bXegpUtvV+qX/hNQdRGMgKEj2x/
YPvjEjfhSNzri4GH6/O9hKB5LW4dxJOxpjZhYWGE6b0jM96YT9WQ87H+voVQ6Xum
vLOQCFevIQLUFodSoIP2l8mRDyavs/ggze8lJ+nfwALB6At2woAG2Isd5YUNHyZb
y+wrBwWIp00pMmAHOM7uVcZkhu2TCl4ELyt4stffwxSZXMFJbRjdNgZqjwKhmNzH
lz2yslBf1nAsLweLZv1J7dGSN9eNgucEONPd6hTLPQBsLQntFFn8UCsNGfyo1jwm
FF0Mlmm/QYqG9iZ+npv8+ESaj1utC9e7tblJlZN7xyBVEj/SGzr24t+pHIL77Z6q
qoVFLVmXztTqu5gnhi25KvG4qXy7RKRyM8eI6Lxp2h1P0ja3mhQJmiQI0rt55sBd
MhXogGWrcRuK1aX0D89Jm1nRfcYrZGpItNsNjBxDJzLVU/o6fXIbk9JZGpbU8iLP
EGFd1LJVYDU+Ad1wUoSEt98HIgvrnNsuxYunLBlydG7rLd+5A4vEzTLhjDUyRiV6
hRqLBfT+IIxt+Mwt9a9C0cBDiSFSxXFNDCd97F24FdIfVXwBMa4lmiJIq9h70cfi
sbsh4kLfUDxwea/O3bBiPPpemvssw3Rxm6c5NlV2SE1vyiTQfe+5fXiP0e8us9z/
nh8eLNi8GYbuK3sXeJvz86cVOzFN4IdqpuJ89qmQEBQf6twgHVY4Py6+okuE2fgV
HuWMhgcwSEXTdpFZ5Ss2c8CUXM7wh1DryuQpvAnaAMqOT0ejYcsVfTxOBcuLhDuR
4GXlCviIPQQ4fPONGR63SOTqhlw96XqgKUtA08o5y00OuwjLreDOACIzwblRqg3N
myF/2StNCkVami9MeAjlWzB/MXNfuO8uNKPTVMlS9038iNdleogwB+Z1vFDDdtJM
vUIDW8RkZYuIpXZRVN88MvLITLsUmdnMCkmUH4u1YpTYn9iFHjmFPTK0A7gA5Y2i
u74lnv4kM0/qW8wQXlnEcARwAaoq/NVQMrJ8bYXt6XJMREeEwBDLCcsYAB+dDw1h
eEDxXVsPExq3CTuLjcNCeWNzVHP7aLa5zrgPQalwa5bVxyht08ZHpLj05UmYe53m
4tVnMCB1TZvuJ7b5BCDUApFbldnPn6PzeDgBncxeX/oIg2yl/WhVXJD5RuH8/3ut
dZfas5+JDeHX4lKl/l+u4srVaEgdv+5+/zdkWYzIZ3d7z9MarpKrX4SdCZ+wCuqU
mwZEvoXriH420RkXzMaTE8jFRy17yBC4sdoqkKyscXDetFl9xEUPj3rs+ZRvQae7
44MRhXcJzkjjSgFtjnGpt648Wwi0UTDSwjvoVn1vYCogot/tGd7jtFMoz9dtv3MP
3XmRSAPBw6Sw1gdKqJs0W8XQ2xbLBEEITsMKClfjnjHnz4EBAuOuQT9+wXX1P3mg
aA463z36x/w8ivw7KvoBrYWkqE8iKWBT2elT1lDGtEWtEC9RTBiXLhKCZu+JBgSk
HQ7OQlJps9PW5nA7hw7KPk+6+pMd/taxFJ1WNHgB1bhsi+bgIZ/hjTxV1Ges9Zms
s3wEFB8zpy41X5t0fl4xyzPAIda57igjIR75ig0I3hyyJtUsYieUJ0O81Bu5vBcH
RYT3dJ5L5kJlQUgb3O6YkgNbmAwRp1gLEdWF6QzomDJ7H8IjCWRVzCqTIgxR9kRA
1uYajCwNCzaJ/8nTULkb+VtoMNPP+K1wlj9jeMkBNJ3sbYi50hJRTt66KE/t/7v9
PW9J1s4rvrdX7E+bKJ+Gnoedlw7tuAgziwUGQKaVddpPtKr4ABHIOW61jCexvdZG
hzy0sCWaciPcLYjOoGjzF2048h+4q7jvi37+IyFlrzNGuo9pTkuwCMYtlxKEvR65
KV/bd0jSZhMXZZj+9RjEPyXsoGKFJ4cMEpS1Ke29h0CKzFExNeY8NcZ3WpK/t+74
I5MzEwEJGk1vdapcBh5BXRti190W2hc2SuQuJXPesWk/uuCTJAe9g5uH2aZINPwD
xvZUq36l9p2IF9swH/S+NlDgG/wvf1AnX9aLN8XZwJCQpi7FmbbOWEdQFMUk37MA
F2OS/qc8xETKenqgrI+I+exaD5e3DKhonQPvSBnCwD72OLEAx0zSecNfKnd+7y2P
hArE0OAj3zJvh14OZP9cgGwN8Sult+pohGzYqmtDWq5aBTls5g1Xd71dtPKoXqvO
0YVzRypOIgf3VgxR0G3Cjgq7yMV6pdeWApb8sXXbUpIgxYCGOvisF8eqZhPtwAIF
IehTkoYnaP6lj7Ipx9+bzQC930e+a70rA1iZoJnnyJGe6O41xo/L8I7Cpz7SReLf
Y44bPA7zC/xLyYZYsdaVkHklMUqlQsqHjJ8YOg9B0/lBsR5s5R9Z104HLEJvqNFe
9ldgJTjxYRv1tFBIygzwD2ujV9KcCro5KOQdWAyhLyMlFqF3rGiZWSpYqvLLM6Ra
5GaVW0kWxq6MBM2KmVKev2eI1DQ5krf90Coaxe4OgBvrdyYws0h0R27A0qCR+ZZ0
lrlnGyS516Iw7xtkAAoiXR0QPT9luoK2+BvAam9fwC8AL9iQ9H/eHX7lTM7j1dQc
BOb7i3mNB3BVhz9F4JPIG0BalFDHjMJAmk68l7D+WnJ1W5uo1YRzZY6hBvECBLSg
WqPNt+jXRhOQtwAQvho8irHxzTT2++PGQ8xu7CxqYVKafozxOMlRyroRQMiMdXX7
EIjJCceypEWGdP+kDQVgRq5+Zy5ExzfAUutifRkz89RhPo7ipKmc2jvwqdxEtbOX
ZNNy9z73F9YgqXjA9kArKsPoJd+rhFN4ujFnZrMl65dDgro/MCfM6ydTwWYqlVoY
uwPbLOeFdmEoFS9z2Rvp+7vbqlWRzSm5qUp2AdmkX2ihv0K2/I4V2CKfneAuSM0g
tUa3imNRJvoGatXbY+M5PfohdKPQLdzwcGc6ms4aoCSaYAXAJKYZjF9eDsjrqZ5B
ob6s5h2SE1/Mj6utHz6szhsScIzJx/Qs3EXSr2+eH3tcw8c2Mt0AENW5MImEhRO4
XfKqMftdpLDF1qVDUWt5w8q0JdbdVcSKaMnqFJsCa6Pn6EsRomuHTcrZrPQvZ8ZW
3eslpAtb9ES17J4TgKzqaWGH5KtOCNx5jaPyRPDBg8bbnH1IwCOR7CrgQx8T/VWI
3GkWE7GPVQ25vMaiFWgbgg==
`protect END_PROTECTED
