`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
01RLvPBwpl7A3W7h04inSiiHUQ1YdfWYXScl5Yf8wxn40RbrvGR9hjbchjwAyySS
+vQGX4vAglgfDEpPGie6QnbAhyg2eh0y0v7lLBnZx1JdoJYxDBbhGfJNNwqCQXuo
F9Qg/m11fiiyOQI/TGsfLg/9q5uxKTlr6jPyS8U0SLhwfhXC98yHKEi48E/vEmWm
bYcTypP1vhKBMUWSQXM/R/wYidfHiQ7dbd2nzkNY1g8uSPU11K5icAHJI3wl7084
WocWnI+QnkKrH/F23heJBAJySiXBOhSPWSfIElNo2YRRCkHvgp/Oe5AE2OpNJjdt
Oph/rf17OWV41tRyBqEBGdG76dEkCZEvUVi1eFbJlv/9akjqLVfqZol0QxIk39UG
iDZS5gPAGS5wWuTd2OnNqoQmQ4ZNm1o34cwcUGh7+Mf2cGQU2KPPg4aNZ+A4VWLr
rWApBA8W6bVOmXgFXH98X40oTzyAEvZlfNfgrGDVtv2fMnZ02jQaGMTORw3m14bL
iHFaUG5VPWtesGm0Q8o+KsTAhVPbrV4nuchgCf77wF8y/QbNM7mCEUnag0ZkSIWM
8AT6M+tQUA2VroaYsvokMAwcCWpJ3FrlGe/obkuRfpG+XD8lGSs9rR43j8iE8V2l
RrmmSfWiGobuOlJxkSoyJbYOehw9L4sljSyNQmEZJSPjf3JZ3vl5lA2KDt4exKSy
rnceaDWaFRtfFmWxb1lJKdze+TNZZuo9AIrIJJYeFySvZylAZ9dyhdvlJUZv9fRM
aeobesS1518WPX04RDcFJLuTHhnotTKzwxQQawKJrBLHo5mK6ZnOg1aBH89OWKMe
sYRZLeF7pjjxoXjw4JBOO9cCl0f9p5xBtw/UvNKcBnAi7JU2v3izNxKNlSDSDCVS
xw9kCiRkCmSqCDsbQ5upNt+3IhALOKMpSrxKO/u26fvP5KgG3rZE4HUQOQPF3/ZP
5lOk9iFjSKn2M2ErE/ze338kVatS8h5P/qa15rz52Lid/YuWzBQI6sOoBrHuthvB
qkrMoOFDWUa/NXDwevSghf4Uo4iy5UReycLADlyx31a8u7F+czyn+A+1ephzuYRj
DKgS6hU5QAsHc4lPFjXX+4mpyrRxH69FDaqKTLPkvXHpjiYPpMnH7HGQy9BfCuxK
9nJSQ3WWvgIb5eFAzG7XkA3jd4cH2TmjayW03CYCNdo0HnC/AqhaBpuIdzr0aafL
`protect END_PROTECTED
