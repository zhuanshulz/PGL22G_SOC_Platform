`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dwshOmp/ofUinf6IDVURgAYiZLpxCXFzL9WFmSZaEfL+d6FatdQTbPMedzDxCrtB
FafDR8BWqC00SvMNU3f/Gcz9HObMqBavfRwCxc+45scbJ++wUGZMXsiEu4sQIpuP
2lA/UX/fJcHRspdHoChVdWS+s1eja31u24fvX/iUrGuai7lWJRRz00vb7JC98/gB
npUIQJP9OFYE+qbaS6np4wpZfU/2JSD11itWIx5t2oiCDR6jdYFSw7qcXmWtl7y6
iWDHHunnxC6UUJpnL55MImCPYKi+0cZQe89GzlkVoQKvqaJcZETB6xCAGodsVwJP
NAl19PkDIS0b2vUY4uYv71ZbpiUhStr3zvyKJfc0vduvXgIcScilFutw5rCRegTT
m4nyQjXiH4yLg5aVKCJ/7zzxX9J+DYfOamMSNO7go1Q=
`protect END_PROTECTED
