`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
apc4hsPGXrdG1iu/SpEmJz711UTxnQkmAtRrKVu0muV7zBCd2w1rzO7RAMWIgt3j
2uvFYbJzNYqOl9IGdltKA9V+svo72yeiygpHQy2DbGH7y3wno2uQJeWI9txJ06Mb
JiftACzJJ7hYkGwOcXJwWpnR7xCwUfLO4+PejZpuXUqCz4H1J1r4rZQYcFwyyiu3
fscK08ZWhSeBxPt7YpqF6y/0WS3h898VFuTKoh51BmFK/Kf1MQ+RjrfFa4jW68/R
x+c4xFHCz7A50N/48UDvcnlmYK9dFjm94ZcmJbuP7UDH9q7nu3oxxeJlMR907Kly
oChpCL4kw3RixKNCAAeSUoBQD+Z6MFTMPi6bdR6Lb2STQQJPAkGtzLU2WGQCNnrP
EB2bt/z2cD57WeGkQgwsQXpeudqdh/hbJFN81aAMof76NNyyS3iz7V/UTlpSgQDg
xG9N6M4QAc8opAFjarWB3n9QobHBNoKaZlWurCCrHYDd9Yeq77ZizfpZ/oIvnKAl
udeXWW72J8FRTRIg8D3VjwRBpkiU4giryncB4Vd0o9MPU4kAXrJeCDa0CskfFi6r
hzyeL5CLO64AAuAeLkyuNA/4p3yrcsy+QH+7Uq8ABkPXKac6nhTg6lSTfTyDTZe8
SY+uj3StO6OHGCantzcd1FRCyCdhr55d6cLmiSOQ1CqlFckpu9x18U2U9a840KhZ
kAFe8XM21stFqCf/MYcyjPk/3lOIEBgpXOaLJNUfwQzCMKEsxi9Cto2wiIFpCQMH
GfSjKlYDdYnyUVPpF2qsP+wwPXU+DeYtEzt/ajypR0XcdDmGeho7xW8E/LWl/W9q
Eh9526jm3bfGL/ezAW01wQWsdSnKlGnSxSq+oS51tMgbxmYZP+37JEHDtNQVZA9b
XFUWYiLif30MJ7ZhSsdmtJScnisMdjT5jbcgl02YHAScMjCQ+9GU06Fr22D7DobO
wWNuLCCRFCeCGl5uGoSAwtFKQuTIMeilET+H5yGL31Q11i4LYQava3H9svoq/87s
GUWz3COiNi3UZsxN2J+PFZuMKuB7+rPl644bQfpjrMmTAoIEzY4vY1oeY0oBmchp
PsDBD5VDzTinwdEpeEFOy4r3Ne5TMJ/w+HEL1/SZgAzEeQhiKoSLqh55Mrlwjjv+
jg8PBSteCLojSfBC4TtJvyeOQ8v8TikpsefTFfZHykuX3qEFGN7XgcWwqnin+CS6
vGoXnsIgLPIGyk/glkVB9yYhOup6ZYG95KOqksy1slfTpiBDYV0WxOutJ8rVoD2K
OXJKXS3H4DRMg/rOuoELUOIRssE05VAQy5asNLtpPEaOshC08r+W3JKsHsi7MW2I
HhB/uFDnTze3sgXZK+8far3uQl1gxKiGYFv69B9P8nRYgL+MFL4PWTussq130XVt
fw9sTrdUb5XjpGuYVFM3caEJIhH5kORYEUWGJ57UsLABTQXKs5z6FhH0Ro7xI9al
d28VBSYtKSG105ttyhq9scADwR8lLG1EF8y9+HHl67FSWJZodjzLTu2jRcJ+FiSB
ttyqyONpv0z64kW5mcz1eC1RUCd8dHytA3PyrBspIgjfSeNR9IG0gOF2uvRWqxNr
J6hFedWm7IO2esyF7gNrO5NUrcoTHoRDO2JbAkcMNfVmJtGNXmMeU+ZcAc8YvE22
NwegRa+sSACMCj+nrU1S7sp/FPU1LqNNIYjbdsCB4Z9HkaULi93EFfpU8WAoLKv2
wz/Aj+xwFxDXnI3tOFWZ1uqG0yNC/8Qq0rJGZ/QWe/+Wh6aU+rXqCbj+10JeNr+r
nwa3IQHedsCqrwsIE5AH1agCFw8LQLxE8f/omFW+Y/lPlTpmHfDHJ4N7Ws/+5f7a
7dPBEPkhI857trgOMwkdc7G8QRIM4Melv76OPkK0DvAB1lA8qWKxccXSGNKXlNMI
r0l33Kz2Q9Yno8bdyVh0AfG58+yt5arddWMHKCy3w18LhEMqWOyR9RTBpIuUCVBZ
nytTg5vNA/dwKt0Q7l8B8GtHJY/hY1mGDjbdUuWdQw/oCcL3FqCGkHC31gRGPgOm
DiN2KCMUk750Fyp8AxtYy6Q5NGyBTyRcWElpVBtJLNqBHqm5GFcup3gD36bfv4Ao
s3LKTIBnd67JBWSnQsXt34ofLspsRXYEwAXrsELy1hmI3IDSCPd35qjl453b2Rxm
dmhxczm50C7xM64s7c82R3HnPYXdiQid5XX2VrotUeNdjOELEBh2vIMNNtuUxWKL
o+1BZ8IEysIJno10ACUjQ9rGmvihnF3LXsqCZ1gbCJ4hUNXr4t6ASRWpUno7OZUq
KjNSsjXdT+rh9Kxs3bc1bE0lx3HucG3k5cF+O5awHLpyGrnfFYdPw/LL1W6JQXrb
eTmSbOQZn8SmvU5xTmWPCZDdkzb11hknit5auZFv/LQ6JSrmPFn5it3HfZPO62/S
IE1JEQLwe6CA4MS+UeU70ATUEjwv78qI4dnCo5vJkI0juABpg/PIbT+dO/g+FFC0
i3KqnxocjvbNnPBkONb8NFES8OKaiSuhV/34/Ch78cYtp1iw9lgs1OrfRwCaow14
04v2Zd5JC3taeQY3YfxJ1zM7weLk+kYpLtdveVygn4IMHiZKiye3R34aKbNurKcS
5qSVHViv89fLfG2d8+1H6Oo4KvytqHFb/gIV1q+4cnyYTlQkizKq7qYKhhim4yj2
7sg1kM6YGmVW0bCyfHGK9KxG4uy7mQUkVG4PWEfoyYhrqYfZE54LBzca9UJOE1s1
Ok49fxFXDg8iu0CA7hyofgA4o7m1Ouo8UQR14kH52FVjkRP1eCMdJFvjlp/Hbh1O
ECX9Wsw8UrzLHp6Vmh0KUCCAtDtt0wjttBmS1a9czmwfpiQsPNbVXv6Q6uR7jEs4
Ln/xRgZyn5IjkLEiwQlhUKKZ1HqluS0djUsqdMh2ER0hIQYVn7YW/0aw7vCJsVFm
qH9QIsPp54V1tuhv81B3ZA==
`protect END_PROTECTED
