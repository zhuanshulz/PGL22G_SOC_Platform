`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c67ORO2Jr1l9urWsGdYlCyOsgrlfg+tHCo0XN5OQELIFViMR1VNLLKfZldMhMNAv
MLvv4ZN7/rFQjhIX91IOI7tKhSB3pViU2Ss2oqwJ4CkH7w63n35XtxP/t2TEoO/U
n4Z+yovU9lKCp3nz6md+onhsjql9so3rK5l3NJlWWWNiT6NyDhDb045hu6ITEVka
tTtHfFiwrWE0gXBcjTfWY10k1rD1HEC8FPqL+ZqTVngU3yhITe7X9ARNZ5UNXf+r
L3iT2249JDBkS/rzEnkb1PYmcXEG7IyqG6cHVqI5xxRJxAN9n5lr9/2MPU7NIpuw
Mg8voUbisTRYzdwB5Ww92S2Zoz+izuHw0ToLSkuVGQapG24OEYXVYT4cxfBFiNa4
8ToEQgtYcz6GBg42org3rDT+uGV6Py1Kjb0QWAMsSYFu3xm01uen6xK0ZoRPEwua
rx6/UjHjCmILLQdEhq/nGOW3DhnnR1U8PRhLOIylPVTk9ScTADWYVd0akplrIJr5
xVR17x8VCoLAEoFrhpNqXyvvKpGty/q3/Ql6GYQFUPG0y0ZP95i7X55KtTko/yxy
Liyll/4/JUWgkVe1fqRajAJC7xpk8ztYaEaLGSmAx0cahlgIFm265eNVrKxHCCWm
p30vRrtP74kM7PUbxq5aCB9mRLrjUJb4kXafmMr/nAa+onDgl5+IBYergwX8ydgA
4APDy3kXXyGvfGLXYYJ3JN27i1kcR8bU1Xf6vaaQpxNlK6xvTIjKaOOVgH+X8MbK
4n5JJkLEYq8sMagtgf4sDmA/1GU/eG1BZ9icxRmiFwJLPy8vm7iXUskGcSB3mS8X
wgpXnm1CSzqtAgUrXhHE0l/mAm7CaqMgFKip+RVoq1WwPzMAAsm7Wfn8/USpVdee
1K921EADwIeA/yuaSQV++8Obo55mb3daohU/0TJPJnpyUD9uCp8XVBXUgb+nmBFt
a8K+0RB/no4K2/O6caPNh9QB/BCQr2p/OIy0BlMwYiSE+jOuaMYYvAnqxHIm0FhA
fnqphPmCxE3QclzgkGiHuGcs/l6V8JLqmT13KQR+reC+tyCfXZYKOdBR4UGg+MF+
NXK+82zgUS3h3fuv9oh+ze72G7Q0FPln7XN40A3CfMncDuL5TW34CaYprof4vPqF
dL7N/5V/CZHes/kW3rKks9T+uc7rZauJHNEvyuLQSl8vnTtYzMF9kTiugjD+vFyx
jfd14HgRuEWQB3DNLJGhYQ==
`protect END_PROTECTED
