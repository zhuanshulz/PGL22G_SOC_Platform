`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h/QpJoNr8+mwEPwlCM/HebcREQb9qiz/a6zAXbN1PDUcwdNyZ8WYmmFARDCmaUOT
1p1VHDv4J7YCuSSMoPoecwG7DJ39TnVHI30w1h4cI+MFSoeISj0AHdYyU/qQzGiG
o3Xi/TvX/v9+vR/HqL8rcJgxrTBEwy+G2iSnyFXP0ZhlZ6f1hXCHxiX2ZK/AiCMZ
5nbTjjfBm9xsT22AeXFLeHfL1MJ3/eP9PP3F+I+GMYpg4hwLULeEsKPnTfIYVS/N
WBCop1kYGSgh/lL8Ya2PzzLRJ7GMB5M/EKVmIExejImvH7xdRnfHTo1poxliIsmS
la14l6QAP6GsADPHP5lRwh45zqRinZ98KV6W9SQ6+hj7S+43xP4j2yVe2gu9g3U8
/TfAwYLMISVmhOG9z1/8VtOsKx5TRnWr2LWrpaOqz5/LXmMhK2M01Xw/BnRkvQcr
ddQ8znWYL7c/yM3K5AmXU4gQYVAEy1z23TUs8Ch4gAAiK6Bjw95b24H2Daq/qi8a
Iv5BWj6T1nF9jacnuMO8GZsB7pjyywKVXnOl+ggE53SJ/3QQrGCBSoZQyE0TihR/
oV1wUK9885+VpMgOqssniaTGmUEcHtfrU2VPcKaJbhfV4ixAyD61JNKlxhllH/ru
QBfLJAsbEj0ummdDx6dqOlKuJK+GNW5PkZm8OyPU+tsLFczGBW2sqlTSbqjREepj
emsIRwolCVPLiMRmVnTu8K/3bhAPBKDjVkFf3Gie5bVdJfJPEh/p3UH2qn7hdoVJ
wNNNZoW+MPmmhIvwm0D5k/4phhZ2ckaG5oft+nHe6jM63JspJXZGaewRJPxr1WwE
1xDd6jCAWBGm6OoRjYJFGrOAh8uF1ObgoF6Qz4ba1gU=
`protect END_PROTECTED
