`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0qBRCwPUWjtI6PRZbABbcIYTY/H4cJ5hw+/B9b/eFmQfFyzTiZSyjIxG5Gv0flKV
PSRT/430Dso6CWXKnC8XkuJRcHydtHa6XkoFY5CfreHVpoq2rvbdmMK7rPFR+DYb
RTOhb0JQZZGhik43oKe3GFjQR2l2OQR5WjDx6fYNgzMoul+VG7f5HWfU6DhMyd/H
ksNoHs/WhaIkr1JxgXLk/YFF8YYT0zihlBMSJ5FwcJDpt/CukLieMKV3PVJ37AK4
UlqaydH8bi+zpkbpLEyGKxdjzeHyds7WgYzSMMVWJDtvKqwCb4AZFjgAfvluMGiA
WoQw6yU1oY0vXNR2xLYm6D4UdXmLnulSvghnTx2+e9c0L3wGTSLwmc+rItcN5i1c
H+cW1zqr8ANGREL71GcXlzcOVzWvzcMLWqv51lJ54UfPHRQybs/EEnIJ8rCSSbDq
OIw9KYv5MFrYupx2I4LYsbkeUtDLD1yAukHHKscS6hSB3OrmXvVNqjd+gPGF62Zn
KoDWjOFLmObAsWk1IEP6UzcY2tGoJyLT2cc0ReYSDj1pVjaliV+q6nHZVL+D+cAX
lzNkgQ8s82lFcKSQ0c4b7H8V1nu3aMl570hfFdudQU74IqI38q8DsyD9bBodxcM7
Kj61KvAh1/S2rNTrCkuIHxidawrEV4AqSfsTvar7HAk63Y/YBGFiKwvtDl4EIKWW
Pty9viRYWkDeKt1EC6fdjaqbWZTjVUfhI1cuHqACLl+CnnBSiy7fd2X1pKplCgYf
8OCfHASyl4IjOtJY5fQPOM/HU0GTdylspaRr+8OFpU7fxpG51KKIYRPPypakltIe
kywlNXLPKAVwTpC3buUXAru+DD+AosjJdKRyg5PyBjJ4q6bP6gAPJJoGCPGSp/GX
uHm0O951uqLMZH70gs4jXwA5eYkNLt2DjDTvk7yhEvCqQzwThGAxV4zN73v7gkcG
plv/VZ4382EAVGvd4olOsz35vAtCl/y+NLfHLB6hrRYTliF0v5irZMntA9vprpYe
xMqgd7NvebflChLEHO2XayZ6pzdH8PCJOlipKZ2/WrRr8LTC9b2fYDMvjI4Yvm27
ftnRWO62rL5Ak82GBCpEGwKjFXQHMUov9jBs67g6G3mjKgGpQoyjSHfG1B4CdOdx
M4urC+alRGB4mXbkrRAWKD51KoU0oS4AqGKdFpOuDiABa4rvoe8b8u8iWBfKs1Nc
d0F2J5hqcvmvDMGJQPvenvuBPW2JhIaOb8CueFb9UZuSlA0pZEHJqeu7h58G3SF3
E6m/9nhSjQCpaBKwRbk5AyYkRx05LupMU7TNbCJDfX6rGFpjqPRzeq98Pn8IXi1M
glizltfLeFkCZVqqSfqqQ8z+xi5GuE4S0lO+UTNdwiDnUKSQb2XM8oLljsqrbsza
nMQRX4YSwtGq5ABUi0ZNViwxjI0JUxIVtB5eaxDVrQDonSBoKSnl5O6/Q5IKaJgy
gDeClBH0SUmQJO8k4wY/GdXNe7ai0I0KAn6AzF+Dq9UPjggS9rUO938ZM/e6dkK3
aSqZoK109TP7P8xZL42VJwGgl2lKqghdI39b0VEGEVKrofLivXQZ/y6lvu+RD5W+
72v/VoPMWXnNnbBx7HvUmV2JtscsDFcpVy57cbofTaxEE2QBMjk5nLffQKERtaKj
wQRxKZZ3RtlmAEC1UIAEZ9+qo5/3sw5atYi+251ZObmgnRXG28q4wVz46O39rkd1
uyOQ60EASvbN1Q4AIORUu8flm65+iciVsdzSapoktC3GaU+QqHuv77vL9YPasPKb
+MpedfOYnLtXb4uaGqbr2A==
`protect END_PROTECTED
