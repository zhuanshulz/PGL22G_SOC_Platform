`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
98Pf2XmmTE+gSTcs5Cc9S3FsPcjZA0GAkMLAP7PWkJ+IdFJnQmoAKy9cqOApevG5
xOyHQ1nDYrxfdm5AT58Ku7jrYrwObWQ7JuEAgmMwpgpfpB0emnJZI5bsm3CJEBnB
Nh99Hnwq/i1+hybIUDtaz+Fb7ktcU8+bpazNqg4FESDtzK6HWZFYX3bBz5d+g3dC
CrzCggz5kEx/6RyVUanhWsHPFYcLz1cnimUm7yg+Ioq4nSJ2ogmsf7fGrLhNjC+o
JBTkLJq68RotXMHWstvqmRZRcLl34/uBm+qAiQIvu+1nYDWGtj98QbnEesGhqjsk
JtZAwXmciZzqnTvZBHTkOThsj2mTMDJQj2748wUT4sc1td2mbZTGGK81XATyrkny
zWC9tsJo5CQbRt3wtMGNePQnufVfhTzS08s7SBzqDMz7WR/uww/HNPsOdnEvQxHL
awQ+flEszDuLw7gZ40/xR7/nS/oj9w8XkVP4BFqSY9ZM9i4v9HtXze5zAKIauuVp
pkxDf6Yuy6FXI5yhSQqJTPKVCK+ZAfnDgDqAMKD23oiiE9YiiP8wOGcpfLhDneKT
id4k63aaBco9gdI73Q2y1HIwVUgD0B6Hqe26osJ71KsmRYLbckDbc3QnxmcwZb+P
CZe7uxnt+6UbKrfEYxPFiJ4crknDy17x5ZPKUn8fz5NLD4lKkrJx9Uzfx6ljiA9f
f+iUkOehHtP1LiImdQOdQUOl+Xd4sSI5GuUQMuMiKY3Jq3hz3Dbuh9wliDuUjfwA
/szYXiF5PpJacwF/xEBp409Ztx/sY1P/FtllzTTgA3pcsIjmVvdwdUprcnEyVHzm
1zmirRj9zxUuQ/yeEDRqPu6Ga2yNEVSXMvApG+75YSt9IU+9dBvRMBVANYwU2Ga9
Htn9jyd4daA4kczjO7vhjuIuNq+hEBulUeFQr9X8KPAE+bYTtFA9UoAIkTl+zftx
VP+Kp4irj1T17AdoypcDXZWoQ++uwXB4dJcu1MCGrpX3tjh0FX1UbEBqYVVU8AD7
rQCuDuVNU5EF+r8z+qEPnc8a33uBJ89YBLHqINCT9fDzxlS3AKYbdhq4e5ezQ6J6
VWkmDjUbxXXwQJtW/yKwJXYxdKT9NPl/mbuVrnAN4jl2FXTtgUlCYUO0LqKOuRhz
RG8mUbJ4cO/3svA3TIGbh1TiKH97Fpzj2Umjzd7b1lXoLAxHVYP4576oyMNSk9Ui
MmImljXmCjof7hhmPQxjOHOiqM2bPUBCxdrKYZ88Ob8mo3nHEkfBPu/Uae88d8kV
Ml8jbYdqfpffJGhtehtamLPQ4E9+fGcPUhXebGwcd+CyDLLfEHfDD5NEgtr9tP8w
2c3iePJv7vYF7mxd9eA5+V6e0FjEYLg2VR/hAjbmMZdF6iXzkyDHnvnhHKzsWhj6
6MOCWth8nOs59yw+2e2pWD+v0UIcEjtUkA0AkOoPQ80bLgdWKjswO00uS6TYMn0D
Vu3buk89zc6PN8RRye5LMYce9+wbgmp3GkgDZhgMaW82O6rbgbOV1/1upeV5WxBr
knz2Wy7Xmm2g0P3r0CLgUE95STW3EMKtc9EFVr6mxwQDeVLM20EZVZvlxFUSuPdf
Edep9283NB+LlskWq+eh6uCVhrbmMRxdGGqU14o9M46lHktNFA6+ZxH0ZGTWzLrS
boihJhfpBHLPFRBXEdH7Hr0V8l1BKDXlKR37KDmr/0dr1zjZKI+tuQbR9YNv+7+S
drdGrVuACrc1RRgQrgHCy3EMyf/WjXqAXyupz18Oeoi/prLgB2JXP+snRoYREtlZ
+dQ+AIXv0qvjjQLQEE0mecFs/e2b0kIg4QTpBCNfvO8qUBPuQ2Ivgahrv1ztmXHU
SpW4BTaiVqu38Tqyfb7+c92zkdgZfbLIBpashb1tHc8siLPapczWrX447nzfQiGf
U0xxPdbFvduRIazbq9J6DWquOhZ9Zo50tVA2v1W7nnlyZb7ZnN4+HfFg1ElZrOoB
dK7A1fLW7ur8cE0uPcbCCSFxDxP3y4uYgWYwlHIPh916LhbOYLkH0+Si34BCgScy
jhPi3SGW/cPITJG6V94UrSvcWHp6/yLWwN/EQ23Rg214QXUWfLrMcsSNK0CDyOE6
JHoGKTTxfwnIYJvCH8xR0GUFEBoTypgKulnFq4CZ75MYEoHTkt/Lf1qcmZDCxMvr
R80Oava8hH/nNkeNgMnmGOAB4HCQie5haFpeMomJGdfYqH6U8k+pPPKaE5/Y0Y5J
S1196pCSGiG90/VtxHzdkLLFGG5UfXMa9LdazboCJ5wZM4YrcuuMeLvCS+XHeNRE
DQZx8hKc/FL1gsrJMBi/qGT1ar69+rcyhCELysK1x3ThMapNzZuhuQv/++LX38ch
Yt67MfM4cZdIekKA+lC8it+fzj0/trwv2Z1ViNh/mHJokn+NUIj2ODcDeM2gphrh
d7oVpoCsAKqyg7qYV2GRLHTd4vnco/cS683t88A51gi/VSitrlvjpqqndtalCu5h
U9vZHniqkwbbGKFZYRC69eLVCj0x0DokAwyv8lrB0Z0fvauzKWlOXDKoX0NntMWV
IKlwPtnnjtZo+2p2ocsgb0F5yP74X+SV1Gg6y1k5fVcD4CtsSaTpWmYpYAu2V7zJ
O0tj9MeYflXaCpe1eg9wiebWgc/GaCMzdRdgOrZw6nHdpH2jTTkq4BvpvI1rHUX1
eRwoMQd9BWxKPmtS7Q0JRJ4oCHDyd91PCz6WgonvVdwxaJ0a6a1k9xNmDfDB/HAD
eqVtgLUF/cjv4IbwJnyi4/Fkl6jIcGG+iH79Bcn3sQID1xdnZPmIVx/KIf6KYvia
LTAbbZKSGxxvCIV5vnlacJJNdjdEM68IXLlIHGpJb+3vXkjSKy7dEV7FTjy+PCK7
OuN3GiydeGzWOdeuR990t8+7OSfLptHs8kNfpIyCA+4oxkhmSbX2VA/VORauBJPx
mZ6uvh8uWVvmFVngTk+s0PS2Hh6SQ/tATAJxlywblGHtbdRztl8Rc9ZganIu8FRe
v5iuSmJlrh/caM4nqtANOmPi5sW6JLd6FXV6MMlTQSlBSAr0MFyJdhwQZJaz2PJL
KL4/MNn309Ts3ZG1YG1mOEVPF0TKi6WHwBlmsqBQ3KL3Vl0v1IH7aPtHZ7jBmWFQ
sS/rso2xMr+3Na3ywjw4NZA0KrkcMCp597Nd3hXT/lYozlUqtOxHfrhwpBl+ejet
wOKDPKPrn5wiX4O3ZSM0vSQTZGic8x2ZyT/Z10rPfyopnSo1eFMFpND4FSFAbeVz
b5Af2hCPzlZwJxQO1U1NH8o9HQQ8yEXbcml+iWXG93h2xp6uZqHPQWtmvI/k7qU+
4JUlvLUXlE8Tez9pBrNtQalb+7wrzK4HBKsH07Uo9j7zCCG6zyZVs1XST1kOGlyv
OAVpenoyRWgXDug1fyVZHt6thXgtrer1k1ozFyFHSQfjEBV6+Una96Z/LI6bSYg9
m7YFXMJfwr3TSa+TJr5jsATwcBvL0/K/5d3R7S1ckYYOQHVyM2HI0Bi1VWqSasFa
iLKRz4gqB60jzUnOkjeNVok/OJGfAjHEUpg8rh3MC+OI16R2HUFNQLelgaUtuEYf
bdNfbtSACKJEz1h9cNAp27PUXtfWjxjI1nhfqMw/0TvW5NG8kh7NxKvnjPXFBJB3
FbN9aIo9RCWYLZw9n1UY8/tUX8b8OlRnZ6DJrT9bsSLlsGjv/qeq0iMshqb1jHgY
dLngTQSKLjRn4ks6pKLlVzK9XH9Zo3N7cJ3zLsap6qOHpOIvwujj+4Rmi3I68CL3
G1VkTqkSzbHpQguyca4E0MbQ+xcegrZI8pJyebUboW0QnrKUgs8ygdV0xbtGiOqf
fPPfd4DfvvSueycLOwg0Sy1UtOAKNK+pV3rYij2rPV2uLXlX4iDiV6cXAystMfiP
n9f/xRhmHWaRawnIpwQRv4w1Pi/MKC+S408f27k7hwOF70N9O816FPJ30hfZHx85
ex7yMAv3QD7AryeUZ2yd0wGSsWk5/bxwUE6dGVzS06S/ApoEi700BG7saZ7oh9Es
felPY9GhujUXyPzHqsjOCsKx2YVehLglvx4/uUZeZLyPha2BvCoohznX2uz1lP8y
ddMnZGMISYk7uZuAhT+dzGo75Kjq9oBVD4/DYFNcZ4PFMVIK9UdsDOeV4oOTP54r
MxV0XKEtlxtQrF/Dfxt2PmChS7jPq8l0GnjrE7GtDr7nSNzXzbXlL1HhgEV+pU+x
tXvbWhyppFLcK1QUky8D3b5gdOtyhedSxDXn7VOb32iHWvbf/0k/1ELirsRtgf9z
EotCL+fX/Jgw3yDLGITWiNifX2eitmK5pGaIz6Jq0fi7O/K1V3Y3a9oylZfMkFC7
kgUTLs9RsvDzWy4VZQf4p72YIhN+zMKXdxsQX1N5wdz4WwabGpdNDimvaGD3cCvp
Onh4GLUepaWJWVqRUw2AajoDOxsEh1X1p7FG+4O7XqkNJR7zEBUQ5OZPL6cjavVi
NPVt4Tr7L2PjjE4jm8oqmMGv/RXU/DEEUfXptenVti9DGKh4VrRGxctB7t3I+WB8
3qz5nACuS4OO5hus4MiNbsEcbWyYm+daDlwkVyugOPkaFXnowcmHldNo1rbjH4Nm
84mUJhEsVI7dkymQOg9+aH0zJwd3SCisCd251s8y/2/IvNSW0jSXCAqbgichRqTY
Y81fnEeUs+l4Va/7DTLmvZal270dLaSmiMA4JE79jFIqRFTgN5dm7uvGhxNKtd6v
vSib1FRwcsILuC6QoRx7IffFQO/8mpjMyAdwAmemk6dtrIjTFyLVtxm79d36nOpJ
34FYRTOa4PqP3kPBS6VPDrkhOJs4A3clIUZHcOaKH1UXZcklPu2J9llbQXoKf8wC
DUMzI3EOB+Lxw0MgECPt4Bn8qttqjrqylzh/Rzv0GmjGSYwZaC98GuYBxOvewjO9
8XNUPLPXnLPtPdzuGAFuXiKqc/Je7DGfBBA6cevdd4zpm/facF0iaurCfqRzNEFI
DG8VwyV32oqhG86aSxMM6CZbRRyLvGil/D+z4qK1vDT7UEzkbEi6UYCi3maYdyOk
+sLqI4tQLjXX96t8I75BbkuhIdeEBMHhNB8cea9vX7YEPFUP4tQInBlJxYYiq8hD
mt4pjLzWClu+S7DbFOQbaCSov4qp2Tw0Aa7+ixALVvhC4qGU/F3wIoP0OHfflM7d
NPIQyBsOD5mmVGFG1ES+bsD6OJ0aZRPT9H4PIVnx6WWTSZXzoLrTCtlQMUGQMcZp
pf3CebPHQMCnRHAkG8m7Bptnkz2R8HINK113WOEF+vYLvjNnWnjwbqvQnEdzPXjb
hH9edEbY4/NX7F+aPyyGuUAizg/kGgCK9MkULq737oAGctqy6vjm31rEQ/8DUJuo
pc5VHK3J613ss5V0MIaANAtJe+hbw/yf4ptpWcE11Nc5CEVyqupIM8Jt2dWa+OrE
NkqY7RJDK2y2PZ/NMimS6SwMtCC3s6eX+meUye9S2s+W3x7yj5c9Gy7YJGgpdS3w
kjeQ9z0e6D2g4OSAPZC8+2g1uhYy4n4hcNT0gqlScGqshtZa8HLnOqDmCUVj3MmR
YpAC/vq5qauNxJHVLK4vIvIOua6Gt6XD52gOhbnT3A+tXgrXbygj4sdD2JNtFgOW
SeO+t7tD0EbZGoHLzkTl2W8NHMPs0GBZMDXywsiLAhyzzp4upJAIZsovLfqAdBoE
gxp2PVjDb8fmBlfOJ4WrJjt1/SO+pQJBj42BL4sXwe2apnDklD+T55xT0hiwqV/F
mTmAvp70CdPAMQmBW2BMJDt3Ze8276K6rny+1z6w+Y3gcboo3mDYURYE4znBXsTt
5xGuaFem6jvK6UqYWlg45RPVLhRvUDe1CwXuknElEbBUu+AhHGroGIdk0wHX1tEl
8IkB/3tux1FylhrsCK1MsiwY6LjQgvgLN8m9wxdlmS6JaSnJbPLiA1cn9urCyGj8
BZmxxIZhcOZVyzZ4DMKmrC7nWwnprg6Sxs9pmQHHQD4chuh7Qq+RkZGf+LG36K3r
+D5TNy7arjoTKD6nXJer5/4QugGVm/DuJ1CnLRZIreEikODLi7jzddamioqKMSVN
wTrtgSMH1N0fYYemEGuXgpexlA8hGYNX70BxCRG78UsQblTQp87Zsk5O4tWk1oKF
uRLw5zDVUQVXXSLLJEOVjsY6VCTZWNJT1TPTiDm/pm0t/3HDVd4a8S19gYNZu6NH
CtRYNQvXednAwDlaCwvnQfzmw8y0gpBScRjsV0ccws288lNRx/ELi/KRIecku4JW
sAE+Oe3iWR8Wst695PDHd4M3GBhtqY5QGpQ8qbVCV/fPI1iQNCN7YuwaeBQhpzOr
lhP/QYRFicPcmSpFVi7jLLGncZGDhdEwz/CgY86b9QfRu2PbEkhJRw7MXnygAgFd
LvgT5s+OAXUzwPt5XWn5ugpzAtIzMRrvmCzAlVx/9OROLLedAoZnse+r70FLbioM
MyrfsuWoUgaspMI9gi0kLOEYAFzUGzBxMvi/eSbFcZf6KYQ9/bVnY5RVNwZ4figQ
G0w3EKolbCZOqDd/FDxfhF2u9bAF9CM8i0KTyZjsMEr1TL/xfY113qYt+PqOui1b
aXVLdPDW0pqOmuAMZdfL9ZNbnWRwOGCCAXuMeEJ2eukKuWKOjSlY1rFJ6+/rvv2j
GHouHQfIDDdbeN0KVUCriHqNdtQp5FkOSCigf/FR8EUP02+YfkzWS8fkhXQ6+nQl
nQF4b2waiY3NJDY5ZcdqoOpDy1jDqPttX4w32zxdMRdwbAz22VQmLDEmGV+AfrIG
hQacKlondpob0r6p2bmLQTyOdgu47mML4OVFYzyFOkzk9tkU9NMDEIpFQvVI8zmZ
8J8y1MDqx+z3/YyfOjCVo+S8i3CTbuVz3oGnsfhFUp0JV1CebBw3Ijff1oskR0d0
Yf1gFz7u25/bttEHOu3dXKyg8N9PfI6XgnwR3tB+H7h/DeUGvX+Ds/LDDfxuh9ff
Pz0VZhb5lH30OcYPwd3G74Pdd8ic6/tbYG222ySnt/+5Ue1ab35vpkERHcq5MsKj
rYUEySkcrsq0lNcgya0FOEbcUWh/MNbUunqHK7bN8vXWGmF5ySVoh4Umh+U62BW/
fl8FHE60qsJAPiIa8kxLwvMLLMzHnwuhRbjL4yg3KlvN98DGw8NTno4XRreu+ynP
1JhDw79++g1fdvm5afwF7JtMTkOVN8S/qsgpHOdFa/QMAqoNTCKJ8Ww06sQqIsaT
c6PcmwIgI/OoyPXA+bsqqeurSHcV8UdU6K7x5lW2Rt2HSj+xszTDsnfJfUKt25mr
mtMxJPoyuLO/p7WVyWx9jsXbt1GKcZ5I6s3uBkLkacS6lAYlJgFP5r5MAW/RSept
4WJ9S2ltSzrqVHpMr3jJ4i4nsSPTcw8t/VjzSmtEM1q1qb9LayOEGePU4/mru97b
7xrNjC5uZ3uxlevDLXVIRxStinnAMxeYi6n5LwstHiPupAm/sR5YBy2xPnF+uJyz
MW4PG8HZ6AV77EiWjddpJWbtjfz82q2cP448T9MO4kRK3CaF1eqb8JEcoQ97Wm3K
UVOrqNVefRWA59b68D/e2eUl4KimVpowk4YOwU/5e3bRpPPjXWxC+N+AM2cWZsc+
V6mUJrGdQyU1xFxSCAMhSJDCqiPqY61Wu5ooAkaK86yhY1JM3Qx3bjLrTdGO7b3E
Ezrt7udkZ/+ek7ep4ltJnxXVN3MpYNzDuEOw0mnu9+7PwuSBIB83V5/pA2P9BaCy
gUMMDNnTNlxLTkBRMTVJm1UFvH2ds5LdPAw/As+YKu34pEkoWi4arBVzYXs0vOY7
23Zd1G0d9v3sAW5kaLHkbQbQBXLXC9C92BPB+nfjMMeyfZiIrvKcKi1lM9e1MnKQ
CTWmP4CuX1n6AB1dM12unr+3E6DwrxbKPKneEGPkTuCTYVvPNiKJYHUcN31v4Dq1
YO9b8MKgMs8jLfn3J5JuvOpklTynl1OgoQjTYhNqeE8E1DeySI42hox4hmUF6z7Q
kL6QEz/tIjfU5V2yq/mWZb0GDpDyvUAV6J+d0zGNgvwmZE7P8C3SAySXPDA74jjZ
Rjx8qbFzCCxJYgI4sgOLEPlAjx9r0ubHAv3VFuJgJaG7l484uXMgl2TRBjhx75+T
Ow6mgulPYaFvR7fbzd/rRZyCLG9MKiTLygYdiJ3am/STdcsgow+Hr5VazHe/lD1Z
rst4302YvXDYtQkoFtK1DdBIO813qB3GvANFY9fMc2/Auw6JHcmdV683/y216fNu
FPWM7+82Ae7JTUbs5EViRHfO+ujm6aJcK05C9ofcd2wNqOFzrPkEgY4dMpsJ7uoY
hGHarlKUxNbdEjCM8sy8EbckT2MBSvIEzxjUgErWfYfdpfrAYRRwmxCAOccDS2Xd
lqPCcgGd00eL8sOlJrjfXO0jDzoI7ybPs646uLl+Z6u2HB6ZYhnzEKZdGbqkem+Q
9ohv9do7dXUdAaSOfji0LVgjVBrdSTkWe1Il32twA7Mu24rPGo8Q/xVKFVT/VAzh
d73J1+IwiA87CZ3zZHftOwaoVTnmUq8Tgsgf2BAlNU+1+IqDTSwmBh37KMZ3K8UC
V0k5BEz5PN7++M1i76iUpxpA2TTuGWhBWl+Klrb9onyvwC91nPXpDdUP6ThghPNO
SduZdC2fMOKO219ER9q0JF7DlW/F22ocrxqruGMyca0rsiUs3TWUHBjVIET0d2pl
Ao8xCvUS3FZygmsWspJ9rRU3yp24JjJWqQuvIN1yskx/yzPCTsXQTyO7LkOXFIKd
Y304qEehuJrjP5/Q7nTrL+pPYWpDKGBXIiuFKouSTaXvspZ+12aC0kKqCiYqxI+/
X28YBB5J/1T10WLhR6wZl1116osCOwKphqOZjv9wAima4zkt6UstXfXQuhKxfHnh
/MW9GYsUQf8UkZLgL3N+h1HJF3Rm2tV3anALl/A7HZsgMFhFOXm8c81wLGFy9Wva
cGmQdmj/k+wbvlV3SeD0HAf0RF2EKqDj6Eclf1DHkJDgjZWnzi1G3pjXF3lCD+pB
3vCor2ad//kpZnHrkwKebXVdk+Fo2qeSkd0VPX1y8WPpfcXriCj+bIzJ7NSxI+vG
ZftBUn6sejlYHbJeYmU7dyqBLafWtnRDo04d1Yvg5wWj73J6JJpX9AakjbUGRoO0
/ygQI4IHEsBrGzg6/7ZtVpcYFMd9/xTSY0Krqz2yEqdCbBBR+Zjzw5uadDLOWOut
KHDNWmqocQMrHSOSvU5MngVtOsFaI70JSGlhNP17UonOoVm3zLPuSZz7s1L76mva
k0/FbAIHPYLbxRw9bz4RN052W4B3bnn3NwpIL4xWihL55J9QGKAFZRTfdyubtr0l
9JNaLJYcSGgGKHEAi+ayk1qvvY2xysYihiB9uc9Ed+SSLMx7+CWae8Bdkd0ikqpn
MrGDGiLyUxFvzpz3lJaPI+SYf5mXP+4GX/L2R7KY4pEGZBiFT5Mj3dHtQ7EkqFSE
lOOFMzlkTCKh+lx2X3LIaF+Y2Z3up+vjKQ6y5+M03Pe09SlIsaXhRt0DMfkZZwmo
J+hvhwpF1lmLGKU8IA1jff0PPQNisHBzhCRUvKSJAgOYGqqTdp3tz+KGJU2icgoN
iL3PsSeDbMLc62s24T862zHNUW2l0TUrzxeiutFh5+WswQxEQiUVCoDdI047ko6n
Yfwx6DUByJKwnplMUYOHhY1/gE6JHPv6nO4Ed15z87H526e/MGlprR8zYm9KYMMc
TrdM0H9fT65+NH+DvuqMGh/qcObiMF2Wd8U+GP7ASa814ZhvBxn+siJGOvl0cFoQ
MgiESMBNIxs3iyOxTJGUVOSh9Z79zske9Em2eMae6uaENr2ffixVrmmPyb8UuQMx
tbMLTXaiTBbevvxF2x8gEeDghUNM21n3OKmqNw4zf7h/scvMzDkGd4w5NfqB706b
Cmz4Qbcu+GRRq/DYKvzdGIurRhhVXYSHDaII4W/9a4DBpzHh6+U7XSqDFbF2rgIm
JUsdYnOxMoP72LiGqP+0/mSSzTHvUaRFgTYiz52cPNc7hJ3KcaKqW54APhIqgIYl
t4oIO+XMKRy5IHW9VpVO025NRQhB1yh9gRzcBSFaEXK9DVB78OZY1qG+c7D0gwiD
tF7qOziYfmVBA8KE/klUutvTwNIDQO126hvkSILWQ16onP8RLV6thy9/xrl05iNb
uFfe5UCZnRzhx5E8hwnX+gW6XrYRlB2n4NPLffBgtEUaE/D5RE8pdPfCD9fM9XXT
2Ruttg2ukvog+8eOWEabgpjNZjh/Kkbb0UJRw1QWg8fuxYiZDTB8Fbjm/BnX3EbY
/ACDfectmo9IMeokb39Tz3OiAhirASXXC2vLcGyOu3geJsJ02xSD+87kvW1nL1D3
K/TXPC7LszX+ioyFdexwwbEYaH/ZVSmUnjcnkgQfwesnEsY3U8Qji9hNMg1IOQdN
8YFoo6pjbNWx2kg5BxMwWnEWIH6unrL/MU4He3YZwcN6f4m/fsI7HEBxN7H5KkBk
ZliYwcgSudYiWM5Syh62QnJ/GX+nLgtlS6OFezv1iGgV1Gh/dErbeiciKT1UunjM
r8RVQmep54eKqhnRRPRwJ9K112Pw4aI6RdrLq1D6rrY5wKO5piyn/QiuQDtuitaS
5yDH12AFfbu6rgWfaG/TCjJuwwXnDmAPji7FecwRExM1v+nORR7kSMTqpyXjGRBd
DzzyadxJS8mjonaHoDZ/M0uVI2TrhTjJGs/mztGlFup2/D8Xy5GKE0NsPcJ6DOvi
BizVz4BU10YEk5b88i2EOQSD3r8nogMz6A2wxjNyxTVZTAF97KxdIj15O+vCfFzk
3/9eY0s2jRdR1lgLT/8wiobL1Y7Q/debSsoXWonVWqcFDXbtRyfJJXoRui78Wj27
qbJHrrcqUQ0F0skih+eYWHR3Tgcv4EugDfZAhPeREH2vknbZjQZ+uIyDU6TP8UJi
fZuukNju70IbS9qiiMZxo9kqCPp+rLofTL2FrUy2KdGpDUbD6sxlEPlhx7kx+OqS
UTMH8NQgY3mX0daniHum67aU9jZZq3A7xqRigAqRPQAXEt2YYQL+B/XZuvcONja3
sePuSqceUAZApDz2Iz5zvQg/tEFScv41mAkPYQzS/yOvPohQ01o48VzW9ZTJ2D4E
pXydop8O3g33TEfQ+LpyKPChTzfD+UIa2SSyxTN5ZjGR8HlPEWkvAAjYLDn5KuIK
DcLPT0AehBQHjpXAewU5sylEG6kCAnsF3oSjPGtyIK4s67sdR34VYl7iGS7M2M2C
7706YhSrIv17K7hrROo8QwV7FqGf+sZZHHOcHFO5AfZUXp/3chrbj/Ea4aoKf1gD
3XRytuVRmJbu++I/i1wfo3oZNsHlMhRGu8xfiVwQ9KMcmVsPTZ02wTeaLHXABQsK
VITld/dRVuCJGa176G6Xqn6rLVkfVV7duj4cwThgX57ubnpHrKriVIydD3mpR4Dh
ETFtHKTIKMPAg3oWzPZiooGNXbpFUSRVoFAyupyE2feEVLmtII3dDDHe34mGHmqV
GtHyWVjXjrpa1BImrAPXZ8aPrzLV+e8RyLDOCES2C126bXjmhCKscI4pZTHOM68M
FT21xrVxn1JgApJXGEXq+k05KrpBXmdLom1JjfWEy8bI+GaLorIC4PzWkjop5l8H
E7Fc9bj3AzZLjh+ZYaW1AbbJOsfwiHVaPLUC9J5wKu7jfzMVJfQ4j4wD0yjhh2ah
lWgLhyJ0tR8MmJwW0sNAJZVW9csisAmW7hi10FWhFRxAaMpMXOTawr1C9SxV9Vow
v1uD4L88ogxYQEPLQjPSUvut8qNX6kY+E+nCsWAcMBwY2YmgClYkZgznRF1MBpYN
lptpDasOqkm3vjZY9JzM5+oMfdoTOoo7zHwhjaD4eVeZ4NngveA/W7DZAQsXlWpu
ngDGzrOa5pbag+PUuo7sGkw1ngD3X/IUu/XsI0XXvLWnEe5VDAm/UiyFRTc2fv+C
b4CrRpzf3K7jXsDhqATSs81ZRVeBB3Kl3AXJCcfK3OzPdmxYlZXYv4JQCi+66Q2e
oFIpsUF0fcOZcudHEvhEuv1zs1PL9fMqz95TYw2IxKbrxx/rPu1Z1c9i1pb7yqG4
d9E4ESZCdCRo9Ih2NRv9UvmoxFq7Mf//pAjqxAgwLpt9KLwYXGqvVAXGxVOVFaYg
l+o2CKGWLjtXWIg2F0LNvRSWzkWYP32Xvag86LWQhfONy4DnNbjJK7/WqUCVoS9t
qxazAFNHRFPrrnmAUWTThRyi/kaWJoSFq0gvwyg6OlHti6c+CAXPTSRg19k1Z2VO
w/kc6bN/Ti9ntG5eRogpKhTy6efy05hvFEIEfw5v2yTgk6p4AqQVYowGI8zPfnbb
/Ck2keb9oBBfA1Q7BAsmNmpAqW8updyOLNaEk9i54wurWhVzzYSJ0yH2T1Fp0z08
HO2f9gqlbHb5lJ2CIaPvA+kEii0DXuMAttC7+Q/7E/ix1LQC9NUZpjcQejT22WCX
FqWDA770y2urHF3fJTj/1dLl2MdmuPIwjHnw4I3EXyRqDrdP4kkvbeWKKg92aamk
MgavnnSgDXwPVi6XSZUipkhQygrkZ/tV4Do6M5JWQgbWmjzZyme9Wj2NeCYvMmPn
mJOD8OAGPw02wLdOo9+icrlUppdEOa576nnutCeIQC/7cgajAQBdqykuUDj922dL
2VLQIt3utuhWBPgQIllRDZwaCDd8i/HSTQ/PZIIwhKoBSpPCJ2MwEFpu2Spy7w4K
t7IQgwrRC51AkjBuyDb+eir5WiyrNoUPsLCwmhJ86auRMWKLFDLIVtcH6IgUhuzP
wvHt3bIAF2DWr8NqSJSwGDp8GrTgyFnc/+RNQjo3KcWmzfS/fGapBZ1+SRVwbvTW
Q60F+KF7EOGf6hEuJrlvs9wHVvkeAK5Rs/vTp8/1wgnhFsX18B313gXRBC04rDYe
yGLmG2D0xs2gxd+0Issod1r1prWREna6Qm0uxcQLsrnN3NkF9Vo6HAG1G56N4f+b
2OlrFibicjGq+Fw5mmLOOE3WnvJqa5/vBc9l0xN4LHnW47EpEUAXNXtvHruCvz3r
Thg4ktbahxshCzIV4rJBf7ZJ4RApaHHJf3LeIPUERdT0QHSHl0I8JhRk/ggZ0op/
Td3pT62VeK0rnrnPoFPfldA80BdWzwh/Uroxqt5FJc5b7yd1GTxX9GYVufLd0nV0
Mktgid2dlM30TS3USKj2Oa1ou53s1ZUJMVTkVLvy5w0Hi0BqbXXM1mRJITrLzOs1
xgZWcUf1bOuJfM+XbDiYr4FFZMjVNvJHWKxcfMa3H1KfMm7hRY1bWpBWlHKB4lgK
zrkEo5bGGbu0V+TQ2oXmPmfNdGGDqZCEzTtKl9OXPFW3VfEJShrtLdXl5j9b4gM5
6s74tOPDS3KktjN6DOvxsFN9hYeYU5Q9AVkeptzcS81pHNH1T4TyHHsNqy/hBRPI
91xsHm+dFFcKCcs6YWPHcH31G7i+gn5p8EASj0cr6SZV6rnzigz3PT2ASTPVF/ks
DoLOl0e2gHay70btTaey5OcjV+wrT5JB4VJS4YJg6WKI42IfEidW5Q5IDnzgvuMp
cKbDI15EQEhbILGdLZI1nA6BgPoRz14lD0kVCbjUiogSVZlsK61xPy0Mc2vKlA7g
4bv7y8rJvB3HHDTO5y1ic7srhjgFhJEM0KxJtc/mVUJtKrmZitOF+4C/2AT9snmg
yoGp/h0e3f9hIODJn4dZltvRzEUi+fywDFbT0kP9YeyBCzxSjtg3wQoHGVBdSyQX
FA4O2RdmqhXW2oGOQyBfP1Gxq/DMeoJUccx8xDJrv/wuHw2bDJta2Snoy0nNy4Kl
FswR+2iEfxJqlRi3lXVjRltolj9umF5PnBL/VRAv2Y29VwM626r33n6g/2HkKp0T
8LcA7GxK7tk3ODjVU8azRcKDf+QIFcDPDZhd5rgGTzZXE1DmhT22o0URA1DaC4nn
s81i3tLTKGMP+w5rdrnM0gEh8hwzADRWH19owJ/fCXKwvyFdSosxW7P2TDzvabI1
dyLGWySt3AiGC8WFr5BVDjisgLoJblZ8YBaETT7JaCCC7ny7SaO+iIBkLtcwaB7X
5xtz7ivHgpIF3/P4KZjDEQRrazUCoAJCzMaOMVimKgtiZAfuaBqcqV38F4q/kYva
R2y6N4MSejsSZ2VlH1urCw==
`protect END_PROTECTED
