`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uCUbxa+oK7JQ51Oop+74HzVklQHoTTkQ+4kBGTY5fLiYviROlZ/NV8SmCLI79P4L
C+A205p0hKSwkpYJfowycxg0hXrSucpz2CdYwmT0gnNEdukxyTBg70APaIG6iRh8
8B59iR4DDtd2o7iw9dCIBeGQA2WlFFqXYfUXvOzExQJnkAlGDqN/osLj/YAzcJ5N
uWAzIDlmSj8t55L6vv8kRMm6WfT7dJrjf0vpys1k9/nOQGX0wJptm5UZnCk+ifiE
tMrNT5iLhROntEO4YieIcEG2GEAScvhMF8fquA+WdgP7V1PEgjAkt6nim4iOW8NB
uzVkzYT/+hP7GU79imkw1pf5va4vBDCtx8oQhR0u57WbEzyLpJo1v6eXrODTeCJN
Bo6d53bawZKv1XVXF6CN9dAOevdmaBQAaQb70da9NKYlsEjFwJww+oYPOKidcsUx
KWiVwhQcoEXXT0acxtvPFDKmWN9Qy/0XGA22704TfyIIq0xBiAteUn2OaPE2DhQP
3BXsji8d+Vr5besvkJwo2/j2b3jrCwTa2rY/QnaoJIyeTTHx44ykWZy8xBCS1/08
WevCyNT1B89Z+xxCWCzLuJgb57FOlF04EQWvMpVgWwWRM/8z5YKIcD267/v9GvfS
eSuk9blAnwE3J1ZnjYqGy9JDSCudKBHO7HYIcEFZwa/YwhEH/T3MrTVVIhkjpt+N
OZcuVNIXI18CDyrKcE5f74FYx0HftjfK3Z6Uy3v5pSdtJP+eWm3X/w4l8uvfJbq1
hhAOXleTX9b9OZTV24Ld8KfBg7bnqS0z8n4vjlIpS+23k6HZvg2Wetefnr4G58PO
U1DGCB4V6XKcNfzdgVfJ5imTmi/cQ5oUJ0ZlPSC/i0VjCD8sSIT0Pjx7dCJKxjmV
`protect END_PROTECTED
