`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iqW+h5goM/IIX0BmOPueCIKSIiHhGTwnvGZ8gIb7LoUFTI8RK909uhKfyfrrD7X7
zLqBGu6QZLTEz7q1sKrCNUPPyK4Zvtqj3LSsBu6JImbNAwG9w6LlWukBAL/0nuJW
yW4BTOgRCGLC3qBuxNNPTIq9xvfxIXQ++ljvCyC0yo8dKZQpd6iba4z/KO0g2ba3
wb5+V+LftMGuu5at+aw/ZmUTosr6xFHaPg/ZDT1Cab6SjzwDOpdkTfT34TWzoFtP
IFN3CD3g5QReepcQVJI4+ol5couL/JiEsIHVZeFTqjIpN5nO1c+PYm9zWwoYAsZZ
QDUnnaNzu2KmIqxDyHA1RfmjXsfuu2kyA0akCGnSYeHmHJa4IbJHKCkIW3fwdk+b
b4psG0PVOGKfRK1Ey3uxLAJd3hgJa/LjpGNqGg6fub1UYbmEHs10UsABI2WpA7ZL
yEXNtn2YJ5RBTWgaa3Xc7a9oOUssOqCQl0yM36Ah1aF8VESXhWVKftrAJsMytk2u
pzXDXZ27wT5ta9UrYjTll+xwPNIA/T0BqiWBMwXyYkai9Ji2c2varTcQgl15e3n1
mwzhpDNbG0+sHWzItwNqcwBk5NNwcu9dscX0KBD9nGA5ycCB8ujWxVaR68ljHu3n
hL1mIP6kmR3wkFOPiBMYOesfJ0uWDSkomEG77gdaXc3XMOTYBNmIYVrOXboM84zh
JAz3FOg0/7QaIGpe2l9wc7KPhznX7tT2OKbLP1beYAFtjt+WWjpzHIotq1ma4+B/
HmJ0UsyuNgcY6l3G4QrVOfRGk4T/RFI13bRCU9/UdC8HDbIf91jbkHipcSWglP4u
TrxKOc3aElgd+KTxzC2d6A5PqDdViW808M7EBKtB3fLK/z8c4JPFaIoYxs63fZJt
JiZ3+AfYG7zzy9Q5nTA8auW1vPLQ/2NSpcHdIU0jD9yCDA5lyTNpdSMLnn6W5sZU
yEJugg1/Od8c7z0+xtaikVARrQFas2Z85G7TImntLuFknkwfELFUOd/z1AthKzZp
WBEZnPv49w+KoNmNklIr0tx76dwgZe6maNA8Nmv3SPwjQtyvPAtzVZIwqSLBNc+Z
f95+VO7j3kbKrDLt5ldN4m/pXmJ1Jlcbb+EjfJCGgTTFLqzHytCGZ7FveZLzL4j+
BZiUSK1qxv9hA43AjnIIbpjW6Ypnae9Bb4ivy7xMawqiA1+8CA9tJ/gf42RmXNFk
QR4vDWs/EtvsKpmA6/16ua+Pp0UwTHLT7Z72FKdGPDUZuA21wHCDVNvGIp/beOXA
Qz50o0p2J1/zQx5gdzd99g5gp21kEagOcvZwTLhj688NLIj+/p4+lWBtz1C2fbh2
t7fbTy6WJSfUMT5tpCnjgZlWmO0yQmsGEbmq2f5RPVQbhDoO5WkmQETzWWqSh1Mo
fY87lAoaqL/HyNP+9T7zQA/unNTaXr3UQQLR+FNEtHa4s7+wKpqJPKu+M8ThY+yQ
zTNQj5jzxLhFazrYdjrvySW576wtmbI1SMU1Q52SrFYh+LzdbfZSwMxXgGFVYqvq
G7aliHSR3hLEebay14X3XTEaEWZ+qiKRAtUGKE7O1h9NbI1KoWauErfZ7PduLNbF
HkqUJpJ4y5hI/DHenVnkaKX8TXhDc6g2hE1li18Xf/uKmASZpjTnPl4TNusTKYG4
NdMYIjmOZ/JQ0SRtyvN+Tg+b4T2NBAo6kbnAWgbAXhe4nw4I7+3sxmsd9P/DfjI1
sptV17J1HHg+gaAk9tK20UBvE2d9CLG6FRnvR4TJjVm7lXmJVDGQSQy4BdJg0OPZ
THljJzmcjTSq6y8vJFjgDg==
`protect END_PROTECTED
