`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jVGGus8wD9cV6LFHly51k/RRXn7Eie2olGMl9obSwXOfPLiWX9ECXgfgFd51Sjcq
Ysnaa88mjCYiNjhsbGD/r/+WTuFt+67/yYMfVr26g0pbHqXWClCAuc64qFvP3zQy
io0RVCtTeK9ZwNVobF7jfV1yBSNn8h/VQQ9Bb3yMBxqJOLVJbvf4SEcFNobXPTda
CzYytNCpdXN/rkyqaWh2V64ANCsYdqp7mNgTwGE3Pwns4Hulfcgc6ZFvSFywixzb
kGe1IgoPpQ/eDKatiLOVE2A3IQKiHe0E1criNJmny4am4+KuzEcIOw40rOCIA/1c
nmQGSJQw2dr/j3V96q/BEcSowEhoxpyLhvUxBFjg66s=
`protect END_PROTECTED
