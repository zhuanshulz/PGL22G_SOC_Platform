`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w0GQ5Unuv3XOTULcEMrzV7XQ8hBEAS4FZd+KSGg1iVnUETKbgS1J7z2SBLGCN0z9
nc6GxIm79SDcZ7438DIe7qZk01h5AK1Vo3CbqT4SdvTwLtAFbUOG9Cy9t6cl23IF
3Eq79yto7VEa4ltV5ZpIojk0Z3u+pre23bU4uRSdDZ8HN/rrnizoxN0EQ/siRDgq
tIW5m+MTu2PSz6zZ/lrzutRB8TTkhEPOFmFlWbLcJSGFXhUE2BbSznxELsSElfIo
p79Z1hUt+KS0aBnaRUMiltp9MvSugvLxoyfd3tywhEdnpMk5xKt5XmF3lXlXEv3m
bpV+MCbpBt3Cqf9hmMd8cAUPrph0N8Yd8KIa+2/Urr5bZgsFtFDh0J92JIIpyGGD
xYnNDEww+gyZR0Mh6dhls2i4Mzme45UdIr39Q6ce2kIzteOu809yfyYFEEmj9pqn
y58NCwmmSZpmY09MujkDX0eY68aSH4LcUB9AwOlvw92bt9TycXtG9nswZWpEnb+W
8ezbY9Dp1/nlp2BWVh3k0z4y7gq28S1zWmA7rriSpRBCDqcGfZsUc+ABgMgQuNuh
7ZBfMD9XHd4KoGJVnkrCdtr28mgvl5BbxGF1qtg5Z7twN1F2s/CuG54Cg8OMSKfT
K95Z52Vl3LG+l1/o57PGRVke7FnTy6R8APtA8lvQoSt/MUcFMBuCLqpHnZ6FLTrk
37xSyzVMbV1zEI53ogz4kC6iaBbVgY5teod1vrinhOSVPmxVRFHgzip7h/6fGMB/
9FuqLkpwQYO5tvZX8of6QLWmfFfNNaf9gQS+Rlw9J1a2oZlpgjrcmQXQLqT05Sas
XGA7pggmq9XN5vG9CqBA+/PbghPxDxXhl5Rg1E+6nGWWGy5HAAMSgS7Uml2RzAZC
1wjZPp3Web1Y+vvTc7lrnsmUhmhfNTzQG54jpWhWYNoT280mmErCGJBtFGJGpLf2
r4TZ1GUINh5Tcp0eoei5W3/qGC5OdAzRl/wRk6VZSqWZHPlCD8sOAWQh3aU1NdhQ
LbvvBTf8uO+iSHK4xMuoJ/LOo4lAnE1Y7lpdmcCcnn99iLHN6K3s6VWv7zhmV3id
IqEJozqwZrb/3BkX4QuNjNBFHL+alMSx+uvFhV2eE/Zp8L9zk4HKdH9fGEP3eUgq
h3h/iixthGgcjAnaZ7gKUNSIBVbUjQqcU5IB7GEO2OtQ3A7wCibI9XvOv+wj55kP
sjBEUHWYYWyNVCTg6R0F8fvOROMJKSTbHJe9zTmFcEKMqES6H2dxP8jOk8VscsLE
KWw53DgUQdpXQflgOkf4xz7e9461LzdFK8PBha8KWTF19IZ4dhpRWSyg/7rhXPP3
n4IqHrmmCxR+3XZefJ3rKvG6+mtTIDTSb1b+DexXNJQ9LztOFoUzeflw56jbeaRI
j997BJK88kTOAn+SvAWEjn3o1apj2KcGGujyvUE/q2VzCKLXycShNblJ0VE1n61l
vHQafobMFnebJKMgibcullS2V5M2KSwEQf88A/o8LNCgGD0KkI2Cnfcnnix4Mi9E
Uz+JEWuM2bPeD91tKwet6Nlw9awuXLY1tW0si3hEg85tfz9WhrGoBMbi/RGmrcm1
MgEw8hDYtRDJ6CH9b88sOmX6ygX1byJIj4teANI8gwYGS+AYmPhtdZEV8MgM0MsU
m1P25rsKDvvTUx+xuD1Otra2v07kBPw9AGtovZPZrnmH/hmzZTAmXCgL5GOzujXQ
oX6QHg4QjJYYma/Lg69mTs4vFDpX7UB/KM/pZnhohA2bvj3Y7We2uWX6CvC2fJRk
aFL3G+OqjFDs2eP+BJdJgIZ4vhh9C8rK3/FmiwNiXvUjxKnVlNC/GhSgGwONEZz9
OG6NJQGIZLb3GOJUmNID2vRdjcmqNrFU1pHlQuS++v4=
`protect END_PROTECTED
