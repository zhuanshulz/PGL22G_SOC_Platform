`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+83modDHxqsV43lsSkpIFVdXqnZff62YbxviRwOCr8fn3Q1cZAAPhQdEm1pVsbse
HL/pGI/m+SGhjCIUNeWJFcIvs/Hcqt4tgjRBfTFgYOzweVcPpUElTDR62BLWYOI/
V71i0rDg7o1QG6iFJMqUY8j8pszTqp2ei9QEFHAdzJwUhazv7ytEkNmllk596D0o
zqxU6dfI1MkWQjBC8EaifsBFb5KxS9raeJNpqpW2HaCz5GlGSHvSFwah/KI+uG8T
fyLIK0sjJR5mXev8ZfbdBRj4EvbUK1ELaKFzR0lDxbAQ3+21g5GGPw2Ekj/+pRt0
Bt+wsllFh7P/nXvb3j8MeQnxsRMr2bJMHbGn6bSvRBofcBcixF3vEFYSUz2YAwDe
J1Gg6uLF5PQvENZ2Ac6NV6U1uNUvYYjvubOkdi3H0Xm/Et/dpFkVoEF0Xx05YyrT
GnrrpnVK4bVhYrg+1S5j1DfZlyCVJ28mnTC6mBUelyvNeCon+DO2Vf+IMItW3159
M2R8AIdJQAmCML5TtCc06oSVaYuRS1WnWrLb4UgyVdjckjY0vBv7Z2O+rx3nvn+U
Nagfy3Sml/8iQQsmJLFy7G3YQrh1bwW1fAx9ZgsFKrX8+q1VGjMNHkrXNzE+8EZf
IPfhf4zuwQSswYuMb7Igtz9kx98vEWgtnkGCXX5hMhIsVbPCi0XwRjH97GUYlmnf
9SrvNG51WdpzySzIT+4Roetjp+EaXKgsMQSllxxX6wYHZWCC9V3ylIOtphCsj6Ca
WPmoYOYr+mQKSVaD/2eEz7WYRtJn4gzy+sgj7q8J0pCPAJqROftSf68QLRAVj285
T7aGqKJxoRjCSR8iDWm4D8kgG2IJ0XjV5dURCL6plCHrGAVBAq25CfYgkjorjUAm
0DhGzJqJy5F/hb8gXPynlPzDkbkIEqPnDdYsn8DU2O5Q0hSYYzbwUU94YfNezcs0
6C6DUzM3dhxc1UY2hjstGKvEnr/Zgx5S0vrvJczCecDTi3VhrJfIMu4ot6cWarhC
MTmNTP5CQp6PJeC5+FlpMIVsJxZJH8voIjUuPp+vO+LiWFxbQx8PMs9DUDewL3+G
aoUuVMtHyVZdDQ24b05CDLMb1jLgBxWZgEM3a3KyLZqAC4JcDBtqeIbi+onDND/J
l1BlUtWhhCp+9t/Cdd8k7wRItdOg4Svey5gtQgR9e+a1KvcSVVzeAXf4IqiAz9r+
BQFlwAdZZxX9X1NxKNPnsFgMQ5sOJHAOq6XmJZXw1cqgacV6JBce22LIDQYej1eR
yANuFjoMA4YpKqN8Ault0s+0so20LXdiuwmScH5akfX3uDvBpJJvUObFPXBdxRc0
`protect END_PROTECTED
