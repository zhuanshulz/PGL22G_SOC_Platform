`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
scTsqL5vqDuPNwJNsLeHW0YvEMq2zl2gjr7IVezmA46uHafZneO6ZVp7BIrESOhF
7iKuM6EIJo3b+T8M2Jq43eT08waNhOTSbwiSPHMnQ8/3bqh73oZpBvVVws9rG4Cv
RmbpnNiRachYAuKNP2+sir4rcERaskCmSdVh5wkQI+zegch3s1xYmNcwoNRKw2dO
5expZlYGpDHSUG2FDsUu/07kLVCirhfRjyZIZA9UXZ9V4YMySsQVTI5yvtvW9Itg
glfnDcjs1bN+CT5xu7872J3Wdx2DSNiaqlssIrzsd/HzLXaodHR2KJCN222eqxCx
81UhC/6iARwjo3aMzBT3cNQFOKt9vSI/CrKi+VbbM6MnMr7jZzs7w85fAaUekqCO
o6gR7GZBQda9AnfRxay06H1qhQFqikpm/rWkbahJGipqdyjnOTCNSectW4mCxbiH
Wv3C/JEGjrufpLD/mXY7pb9n6ETmAlA6/bBPJV+gdkMJRpzVS45Njx2gjE/8C0Jx
nWBJvrVaiKiYTiIvWfTPn/GKs9uwOVUcGkk2KWywZ5I6hVDXhtchNePEoZ3cO76p
AlhWj8c1kt1vaVZmxmUAdnKGOnUBahaiGbjgEB/ziAMctxCYVK9+RU8ckR5sLZ/P
KF+EMN8cLUrP7dIvzAtzhp4hnItq6URTQGRqwteeuOimd9caVO3AEZ6gVXiTEKnh
ctUAPdUtNVNGs/9tAgrAT6tUTeyRJ9vadHIFEPQO+8qwWjpoaUrTbk6N3dAZJDor
qmGh0RzvP6q9eOJzaxF8CFYiBcC/kirmH+HUwpiwclXVTu903os/AYB5u864Ra2U
aSADKRjI/ahPxmUgLs8jr/fPf939qVhqLlu7MiCk9dE7HlRCQXc79XZI9narFJHI
BlJu9Uy+aRQWSbcgYKSXkJsZWTa6ybY8J3nXHjDy+OYJP+yItxi2OZ0017yocFCW
ZQNSGCt+neaEGdbI4zpj2ctrMiXLec29oc4r87EGUDZG8hlgCoiGO5VpdhzEUEAd
rVJRJa0vxrvyWv3vgsoZ2yNZqGE1Mp3dHRwipqxVpBI3LRMIlMwodlVtMpOiD73W
mxQi8xLsNgo9gytACMyUeHcCOu5HO9jN+hdfo+QB2xSKAOgXbKnWj31QaUz1wx7u
jAsbs+rum5+Cfgq1fgQ23WnydzlTYT4b+M01zr3JeEyEVq2m2q5tVlo08M0cJtRL
L4fH+ua6H2dBxWRg82FD9ciWSqZ+WmXcq2cmztcMqDAChMdCmJNRPsriE2w9vhYf
w67P7eZJOUyZsqdRRgvtBvr2V9+kqUMj+rNKkX0T6l2AnyJqQi0su7HMszc+Y2RA
yBwl9sf5qtrswo1U5yD/YM2kjdjCSaO8Ze2l6RZUgLCPJXTAsqEcSUXinNSZrp/s
Hvx7KZ6xUJ61DzZwwtrG/mVlUnVoExAfMJ0Lb0HYLXcU2wenO4iH1gudDnZk6mLw
H7Xi+FGbcZuaCf2l4NIF3BiLwex0JAdfkshqN5CJeWivxFaa9WN+jEp554Ni+am1
55RQGrOvh2KBbXNQnNk+J/zpLTdenfNeBG0OQ3IPgDOK8Swndnqm+n+vHwgTIMGJ
k4i/Dl+4Gwcgm4NB5zT4R1MBBS80Js0sBiowSCRwUNA5EB2CCDMajiznA2g6gnjC
99VfBYdzTDgJVEvQNkh185S+iErWi6c5Lb0aYuZSOtfn8g/23/7dBk0OpE4raDxx
KCM2vO+XKog4UvDpSNPmtDHUEzsjiRaEjQp7utTe4vZoso7ixdaI0Ncau5dcyP0O
+xpewZQ184rZIXLD0GbT/04y8oSi67NEBmi/Lvc6LQ4y2I9ADGIdTdgGQVuqZx0j
B0dq3mtYOkvdF0rLbOHVz2BjNF3TLgZQOXOaOV5Nz3cmtLpm/0+aTb+HUiaAcREA
kKFdnoRvCGMUrclsi6eCrvd5PBYkig4kN+R38aMKj3ZzbqoJTHULmZuhOJurDdtj
v0ym3Im5Ebp3q7/bwb0z9VnXuMJwbUmIJQZtbfjoLV5e3JILiAZIpRvaLxVrFBTV
X+/Ku0ZcFez5YDZAKs2JZd41RAgcpHeYzyeY6I98p/Y3sW4cenvnAjfWoNxlaa+V
zSXhTEvvdcNuripGoseAPEy7y6tgjqjhy6x4Xx/7HWXdtRcrRiLpse+p93nVMFxC
M0/MVv2P7qYiLq1i0ZIJfX0WyjgQJsgWtVEyqTXRusXqyYC7RfqYW8xawXArbyU/
TVQPbv7aeOOOOHBqQX/EpZ9306eL8aA25lKr8izIcx9LFqD4WR3emu+4nhqrY5xq
CNwpsaVuknWI2G2Vq0j5vOITpfv9OlMqM8G4GzNOWsW4VF6JWi1sJoo5Rj5e47Xt
DTWkXjmtoM39LWJf9om8LqgL4+h3+Gv8Pma0c2VdhHNQwq1YvF9TxWh+983+9bz2
QR55THYDFEnMIYG+XduGQ9EmqBEepJDVlwc1KP/6UvQMMmVfJBlgSAscYek0/WsL
XdNb8rWaJFGimU3gcshbfHY2Sr0PoJC0uhyvXKrrTUhzHG6iur6c4wvBahPF4Obd
KBv3nf1NgYnzibCDRwSux0Zm4+xgjB2C2SaG0JaM4vrJ+Gc0gxjUwOMFqpfZG2A6
EMKhVAk74X5Ovav354Z9dzOMnXVXx4RW91mAJ4h2ltH/kePNKPaKxaGtBr/AeRp6
eliA3AGSnsRKDtGzC9uVWRTY7fOe/GEqLzHpixZbsomDDOnUfnKR5rxh9C4tJHA4
mnY0NnUzWnYUT3LjLof4PyRbKTzXwZm4y0YUcnzJOWgAMY0AAvg9Gc8JCxTHGzwQ
o6WbTj7C8BTMNvtN/F0MS2mI67j6fCPyt0HQU6lC8kLtAwAw9IcqwKNAN0pRBgyC
ABPJparkp7LeOBvQ6ExfmJB/LktqgY3mes5lxfETaBLq9AeObHRDWOp1UsoHcjtA
kYp1BwJGAIhTWlFqNK7xq5FE+UMnAP2f9hVcJG+hsIUNm64pN56U7PnaTchDl659
XtgHbFjB527q7b1htUBc0XzhSPGVpscwwR2mREQPaACuIWvdHZtaFyVKaaO+sEjk
gWq9/dwIdJ2qyjIX5p/1Tq2vdBGoZ2M3MvdFI5qZFo2DzImmDVKOoH+DYJzwg9CL
k8gZCeEJhC8TYl6jY8hT82pGZTRaNbzXoqeNU+9W9/74uoLXNaoD3/mMlBX9kmt7
gLHXsiw3z0K9sEbbzSAVG/L3Cf4Itn2WqluabLosL8dOmS2IYrs95X/O5iFb0HR4
jPXl/ZCrY1K8U6kpgfDDRwhCaPhNFtTdqWYX5BqZBjDUf6LxM2O4gfHEH4aQyDB+
u5bdJcdlMTUBO686L6ZnYGC+BtFuX5kd5KpKcu7gc+m/j5rpeDAET1m3B4rANGKi
ocS3SD10LqGjjobjyhZMRf6Os8cc0dytW4JRpUDuPJ71/B2gEsuN4yjyRm7qACvw
NiE5KJc/OCDzmxSq/0jUgai/+sLPtDbRL3dgUbXXKI+jIwjkoAStWEY7IBcEEaUd
L/kP0GX334JJGxpUH1mZNGpq/0Vur+AFRxi0081RijCmUVDJ0WwwoCtNZKwHt0CG
m2/WzdA73XlZxrijwwXF9szqKJhTzP3q7ZgwoEiowI4pzRLEXYtw/0zuOFTPM4Rz
DSaXENClVSUmK52YFV3qjrhNRGvrSRsHSaSFjmkMoRScIotKDc6y3mgEGDxqrexg
aWTlT/fQa0/pJHKuf9Oi/3P+Uq+NNQoA6NbSPRK2Lw4laGmM7tPEBvgolFbXnDDM
xHVHdT2qtK+7w1jeuVePGxMIRsMclSv1/JEU9kegdDs+0ZUJe5X3qd5QpDjiTEft
eTfyXkyinciOiD8FcEeJnz3+3UnvLQgfjZDy3xXE+aUdcBlMSfSMV8DXCYPQLbLO
baiQajI6jS/lYYZoFbyW1U/vfSzmv63bvx5uh1SEfvJAns/nua329nQqhD4JeTqZ
gdYCV/YfHalJrMN2KpcPw5LGGn49dmYI84z582sX/lUvjMhzzZW2NM7GomUGhxVN
XVdb/KzJSvRFKvpgLhmWU3nBYotydphRj6dtaX6CoKadcWH23YacX5XTgaGDdo27
DsZhMSnUzfuh/qgSbq5fGOYP4fKdNN2YrqU8zDAUAacJQMtVWXRkDY80ofYkYX8u
J6fE01LEWr6lpBDPRDFEa4k0DlN7lB3o+2QJ0Cm0gzKAoW+8Nsbh/Hnj9NbuEoz0
CEswwAxUzKEpZ0obcEyaTzrkWP21UcpTVxWpehYm9WXa3cXe7wYaapMHPZYYKIuT
CayWz0NpQdVngRdq3fp+5x01xCbkYrQEU5RDCKCz/GvTZWFu5WVwdzKAFeoz+vP/
vfI8hpK5j6FDeDconZczAQAhjZGHoaw5W9m/Eyil2cSv0yCu2YhJSSeycT75kf/L
ak9jdfZmHszRvhqJi6OgoesbG+zu0+wNfl2t7i34Y2gEiHDe9RkUDHUt9c42SoT+
iG1J7VLK02O3KkLpO7qDoFyxRNX4M1R6IyEWLJmpshvsjqLjKctj9CDSBSbiu5XH
FVNZKUqmTIhsogSGxfFOmOfgmRrRPUmOJqhHO+tDMpsDvbv05GkVfjTg5nPeaz+I
hzAd0UQpUpSh0CQzFshbE8I6pDU0une8Wa1Prd5/dTPPtdAPephx8ZhtFlcZ2ZgW
TsrQ/Sw1k31OoTXa5kB9oFTZtctqwZAT2iCwdzgCX5cLSkHh2K+khDHOgYTs/NBR
uY4fwtvMpPPiewCDl++Nf+hwcZk5NtLkl5+74hqkf1M0QHAc+KV5dkv1ELRd1FEU
zA4VBf5vIecKelfy4UUjazraUc48yrrFDUAope6vxT+GmFsCVYo5IKuRw7PDWbAA
InhC3RzSUufY1iN68B2WdKRMBpYNgaOH3r6R4csYO38i+PWtfBFTDxnhLGJ6MCCc
rrGNrOpBUVGRu4Ih+MK5hz8+oLbD92UIkYy5B+dAFs6M7JmLheRncE16T3Q4y54H
l6jsF9d064yc6k+VHuXpM9pL2gNuAVPh+0ko7BQL3p0KWK3YpOmuY5SsmyrRk076
hnL71wwIiXXoYHPsvHzvqRJVB2Fai8b1IBsrvgteA+s7NI6DtHK1qDKCy702Lyk0
y+9uxOkq3hr4VKMTzDnoyJqFI/BFRmz5ZDZQ95PXJQCGIqQYyMQHdLZPUSuUiGTd
GhodxeHoBcMPkUb4FknCHtSh+jWDEM0e7En3FQNS1oP67Wdxv5FdB3NXoq/7tCJH
VliTytZlLNItnZsKOhLlsVDxVthmTiW/L8v+nj0+QCFsfgKd4+rdz/3YlMQ1kavS
j4eAuYSkSzqjZNhycWFJ5VAkF7t91mPc/LB+JHCa1WgkQy8ARX0hP15kmg6fs6jo
dHAqPOFFbh/KaWh9HDmFygHVabrmYmdKNepuMOtWTp7Vvft3Kycr3EMhLFXrOEPj
8zBEi1mPTmocYGKhwHDAv+gvBbbGMHV5Z8g2P4QWtLQ2jajcBKT1zYnTz1zabLmv
rqZIZ/k868MvdsAKTluRTKqXD3x9W3At2hEopSMpSeBiXTGNfb5nnKwnSvmGOGof
qyL6j5t+sc+sC+ifSh4EQFEug9Rs5/1udmETa/coM8286xS1Nxkf/2aoTQ/XMRMk
dznUHM6Kvl1uiTLo9ftdcOaKTmP4WxMDDrnRrpx/jMXtq+RmPLkHsiGNAVeyqM/z
1LTfqTHzh7Rbu6U2Of1GWaBKlj+xGd5B71aU1grUg3vI1zR3jdukLoXw35HAP6Pr
bJlIpZ7Pu93pFf94CY6n1O+DXVH3W9XUXPInyl0V0dI310FBj3I0g1srF3tKpm5/
XoxRXQu7bpW/Ph5OFv6dLMwdOXLxtJAqM57XeoTXaLFyRAPzmzeFQtWyxnEWCPw0
QHyYVL860GONUuOZ91u+Xi2Ul5Kyu/9mQrLe57+HLxCHkhIbbzhhmIwRqyVIbmX8
SXRUQiN2YuvJNOLiVBlKFpGQhQk9QJZcsAnhm46KdaJGDRjmNJOlw74OBK4Fw28h
L1pWXYpsHLEXx8GC/ARuBZVaryPoDVfdhPLklf80TfjBJ6FXC8DPcZaHvEiv63wp
NqiEn1fx12Xez9JFNV7FVCktAZfF6k9Ru+Tx5Nrn+MfeGlfamo+hj6yfEnyR+jN/
NSHXkCX0KSxij9PNwbJfRYeg31GbWOSyUA7MgLn+UgV7JRTQmQMk4sZvPBLWmyWW
YrymmGKtDIpxUY8Qqg6Q6VmGPFkj75Jnxpsy9Fdmrj+cqfGLNTaGOlDg50IZQ9Aw
AMbl3ldg+ikPWc5sp5O33G3mLuGxuJ85AnNdQ9Grn24YJ3Zq40LYJpYBQahjvIfo
gFeAVUxrfWuAUwykq3TYbGeO1tbHFGKg57I817PYxjqAEhrUVhD9jTZDDxFVRKBw
xw6H61Z4annKIwADJYeiDFim6NwF5zMqTVCyppxUbZpVR0dE5JMz53+IDQaZ72sG
/vwEoZPiW3oCTtSpdl476rjxTBmMPQvXpvP1ComNdgxSRFPPmcAAAeu90wsM1k5Z
6fmA5h8qJ+M+MmDFbmSkg3hbzEl1LBspKqAx0kHcPcCoW2b8sLCYCJQlzn35/OX/
LWNVwMA+84gz359u7AyimRVn0QiFCTAM913rV6/yxYbDN0urq2QgccH1N2W8BWlf
ZqGt9woCG34EclH+6QcXoR7SXSW3QLd5YC9MB62olPBsUruTdnu3KfrZAmaXpLyq
ubU4S4OkkWlOjj86ecGqJsdIPpNMShyBAQAbz7N8XnwbYCbw07qMwLf8ZAR/Z8tl
7bkuieNXzU+u9JNkQGxuS14e9HH0GPTtqA0x5dYcALq0huaRLvqykTG+UAGE0P1A
egR5UM9xJBYuBcq9w5OUr3xZAuef45LpU4Sd/IB/oq0sCFr1aR/M/10+q2YNE71y
hmsSJ+S3MlvGfxkJsvfiifQiAbHEo7Pw3KCYF4KqXMR4XxPfBREA3CkctUUCSy+3
I4C6m+ndWFkZ1ocOylUFMSVWvfYCgWHLy3aySZbONOAy4OvXhU7ARMfCG018WaUL
zpszC6IYMuRWk5KzJB3+lMpkHATRFiy6AOZcenkl5uYU6A+GKEcDHpxEg0D8N24B
fKALPd2aBo6AC/KhHTUKh0sfMcPKdKysgkl6DQqis62napterCqE+TAJoalSKSRm
TqTaMSGl6/N3ofQlJUFUCLb0+tLHuEbAyDJ12tDPp4SYrNTrYl+GWn7QHt2DURt5
fn1UddDBS8EMubJAqphWTB4Y7SKgoV35mzyAEGDNM4dcC/o5ioKStHdIPveFN+zi
P3RXcbSUuYdJFtDZOyUmBZupD3Z3dYI+Xn2tj5T0UA5LDQq9VRu+Oo3gcdW1eITc
JLJqCX7WInPOtqnGFkhtJJn1ci93PvwC+fsXEhzQLvbOqBEQyxtyCgMGXkdqHVkl
zUhfkfEI5P2TA9wFuvlR3HQeQ3Bf+qM+rTJu4D35QZzVdTM946gBTWrgJGHE8yn/
7NvMaDcuNrzAC2GDCq5UenxfdQ9owM7uPUyXNCwlhBy+E5iNozxhG50M09kpLu6Q
+ZC4N3pisviYl4FlL7W8Y3sAG3vCOKv0jC8keLnnT8DCkw5J1+NjyYcE9MY0qUnV
zn3P9bXGD7V8QPMpQrtcmRac0SH318KLbap2pvqyuE92k/ffsyq1U3vYLHTgyqxs
O8MOfEbiMVuE3qYxKnGuzyKyrXaTNVhhNnZ+sJDh9+ami/0ccGmGRi8JTjzhE38h
tb6onO33JAGoqqm557xLz3jC3XPCqJZjhYok2lc0PIm1JbsMuaBkrzKGpvYy3UyE
fBIUetfq9giaKKd6PDEVKa1XSj+om4Nw7xkjmXwiqnPA+ZamE2rKLWHjo2U5VZqV
XcSh65q9fvFkla7bR7BlsiS/G8EHKPko7c+4a9pVFtk5q1TA1+7W9AQ10fCq6hlw
1VRR8szxpBxbvSX33HJ0ryyhoxrmkpthAOV5lLIYvd2qPg1pCeIKUxB77vjmfyVR
ecS0IAub507r8n1qcWZg24gAbt0lJX3cq/6zjzuXjFXIr4o14n7MFoMouo7YUqDZ
llviyU1I79NwHKnK3tVmhckxadAHtMjYQV3UMH8OjbGTV/FsZPQtiEu8udYUoxPt
yOsU70hcFCISCDBM5ADRk0v6JuQ9AUeS3zV1urLwGYvyaP6F3E83Ii5P9w80e+sm
/DuwzYAimVNcXCILSYF42YJvJgWltuIHkjZ1pojkH5WswKtTu0RHjaJsvytJw9ed
5G+/3u9OVq4n8ZFUjEQmp+DpXWtTMCd/T+X5o6RBWEDvdPdNGQm3RHL/ybkF3qPO
n/7dzGHP3FCGnCmtEUUNoMYaikzydBd1csN/XioCYB5GQ6mnB7NQ3YsNSCQqrPQP
5oTCW0ex4RAaHjyhim4Z7Y++V3t4KZXMfG6P6bLKP0HszEi2sOuCrrV0cvQyGsg0
62iyfgnFOV4cPJdoU0jkYQEjJL9LbW99M2t+NhXh/FJ7QGl7fIgXZlWX4XVKYxLo
qZfipbw6lX9X7tXln4Lsm/K9qGcAccoxkqQo0pG3UejxzvlA39srJJQey94Y8Rx8
S6ojgtMTfjvMEo+vL1PRg1PKHWr8z8eSDvm0DYPctilOyWnrhX26npwzpQ0W0dol
wDs+01NsAiDaybdZokLBkodw2cfqXEUZhmSnNQQLJRw83fnsX/EgKbC6rd/zMgmY
wY27mnc/RQC/3+CbZjuQbG9pU/tzmEeyaH1Db52haKC9zIXpII7+MqNGwtc3F3tp
yEMkrmm3NuHOehKJmBos7vr6VoXlIITn9JI05tMEvThvPkmHZenDJzJpHyQwMKac
MTHEab6lR2safmaW1oLF0489qQtoUGHJQtpeBezEd8haL0XAu9zZMsX/DqIeAyhq
ZbePViGARHz+YNAjTukYjfhGDtO4MJzLVspzc4ijrR37ZuZtZIoSI56x5nKOQN/q
YgeejY1R9/rBkW1qrU4dyrYg49B48ONfyqIeNSg29z9koOF+kj1GyA6O/Cg+AxN0
PXhIRzzqWJ8Q+Oklly8F3alEQmZ0B+wz2BQApc9G/GJMO+adpgdLn7lv4dLI+1UO
ZlzrzJV5dRsfqZQDaAsBOMS21jghiXGAeGxw09bhiHFpLIwrppEHdx6Qu2nogPFA
vBoHXsa//kJpuiZcv7XuohRK6dyL+nQRUoyB7goZ85wAZxGjQeflxxCTUIC4zzOS
8gvOrrYmXFnxMDFpKFeQHaC1r7IkiTiuOJR4ZdwBmraKUUSZFEde106oqkrEb9mq
CUD2hc8h0mcbcM7gv8G1MMCl9dGSMJHoKCcwVEg5dg+sCS1WOQ3OmPdi4k/GC09O
oBKs7lewr84nete/M/DTGZz6bhWpueUdkP3g29DeL6s2Dsb37Hks4j3WcpASPiTa
EQ7Ev0gnSDq4hS60w3z8O3NPVEs59Ys7nIAGyaG18thAu7tQYG8ZjG2pGlqFEysS
wg1/TVQYmjdYH+s/aeziDKCTfUTTTmYuD6+nJdhD+12VB8spENJGbz6gElsVnivu
XyMPYZuXzErbesgyjoVR5fBKW03tKvdoFICqMF+tbPIMpDey7VJUSm42XNayT3s7
JLpArZ4aRuTooz5iBzeLfMpWyeXA0bOehU2NMTQnd4kjaQn4mDh99CEgQkOD3Y0y
HNsxC0jClBxIbEhUotK/8TdNDw0qB5p2khBIgYLyXnrCQBXQKOpzKf+tbaquOr1V
nq0a8WBMS5vznocKXlXYiOlJFblsRdRbnyt9yWnLGV3xq8E/sRl2af5EIyHEqFV+
Tb5rTQ8QoWf6V9KORU/fQSmqF7ezv9Czv3d08qDEXIwnioES/fVPnEjVTpwwwMzp
toPWVIazhA83p3UtuvAqWzGwnKBPoAULsTyExMp+661KqrOCVArRzmxrIbsggU0k
6UhTBfllWHeh9STUyrNU+e6YIaeyD/KvjLr7T7mC15BoHA7wD4mNdWtQiZxURHBq
/D2jMOx8XsrMweJkXOKJPrZ7IotAYX5oYq0ZVgYm7PtMRVA6O2/5xsILIGURni+w
FguwHJxmRNKeDiGmlSzKabtOFoWBhx9p65YMBzWZxbPI6pM/0ZEBowfJDW1CVqIU
WWPkJx10z8atRIGhX/kRvZOr5oDonOhcreUitD0ayFtvC1q7LtTMuP2+k57BpxMm
8UHvkVvoi10pm/w0wk641bCE1zOZBtXus7gXIFRd+Pgat8Ymx2iIgBWM5q20cgvp
Dqo+1K4tDy1xDKqWt7oC3n626NlDtnJbvz6iwksXYg/MA83uxS/CDvWAh6W8MZN4
UtBvRFehDkqNYgEptl1Fdx26UkxLp+bQ4OS8fDgMp/TECGI1qQ37VWO/6x87GoAq
wnidhs8UYMk3Zn+dWT4VsTuZskBeFX5sGhqSI88GiuogOxI5vHqLrGBZVQfGw2MM
D5vP4NdAFPBspt4DqZ7HqfhCRgNUmVCaJpShJ334+dEZr+c7JD7yZcDadL71psek
luspsRc9YbGwm7HZYoB0BDI5JCRitwfQpjQG4xnWKYzX3BxEFezPoV9VD4vQ2hJ1
GXWEoWbVbuD9+2PVt0Q1kzvfuMOo3ruMOTpLzx/aVNL/dLnuseB6nK+klDllOHVo
DC/M8DpuIbIZsK5rfLhjb3KWrEttyelCrhVAqN6dtPC9utLxM9B/qegZRcUFVDG6
ld/47Zu3KOSW64OT3E1IdkuuLFE0UcvL4+Ji/Ff4Y1xv332J5MY5M/PXROD7Y6Rq
WvYWckW3vX6dg5wmgg1vA7l8YO8pVRUyY9o4tQwDAIjlT/GEpgEkbasmiXXDHW8g
HtirGu9skFbUP+oh9TjSeSgknjk5wPlJLtFjeX2FAFyMkBt/ea7Jkg5O0/rbhUpf
JDEf3s4d6laAWmTeMSKaKvK2fIY8b435fc0CM2Z9E6Z8oN9Nm9yL287QdevXPMe0
kauSlgK/EJMKklK9izMUJDM8iP0KK47S1WtnvsfzKWGVidR4Q1zKo/ZJrvjsqP1r
k/Gg5VO1KIBUp9dFA6EVBUChLCr2gjyYY2uo7qobUCEeQBsFWjWtbOLaysvfNvDI
DJ3R3Bvby+dHnlI+AaRdxU1Mqb8NsWd2vlnXlJkMvmpfyjAM56G5TuDsP3U57E7o
qnUQPC+bao6cHnXsQfgaQUsCizEzNqbHtYF9jeXFI4V3UtUZo8qi8N+u1Yzfpttv
nzpxFvjE95/JwVs2cTh5+KMkxzipOFlJPkg9w106LbdKjBBjCqyWlco301Dshw68
hzTqxsvwgUSH+SP5fKMvnq9gy88m1B/2m7TM1PaQlLvOtWwq8wpNTYZanTNvIr8S
XjxuwnuXFdzXf4agkmKheICaykvXhSjpESZq4w7q4PpvZHUh5Yb9I7YSjG/vRfnX
JH+qwkixqcNxMdk62xz5W7AU/rUSVZhc2o+OcOnYb5f9OeuejKecbV/Wsmn3OoHL
5a6xemSKBC6LAwaiYqp6ZA/3wCwOV7nCEdfcbGizCx6CMLXtz4PXvAALxkTyNmlr
+wrtYfL9pzIuGvFvyKWxmontmyaNX1X0Tii9LXMXw+8XVHf8E+VLYKXgAtQIK1mc
MgHIyPrAFWoe+SwuI7qPEA9tDTIbiBK6Uwr1SwcJ35iSsx4EyFP2JpVsCz3o9QAN
EqUbd5ZwH7zm8qjngwZXHQpzFclmaJsauwDvibiO2otAuKWtNz7U9L7W3ctcrre8
uYiuSP0XrebNQFk6jw6yad+ZqvImUH9H+EXPr3ec/cF9608+y3SbcMwxQGp1nu+p
6zfaVH5e8o1gHd+xmBw41CugaayrAJ9JOzG1Jnq/tVwa5b76zp2OPurqbUnoYt6H
A9Bwp2LfkNzyGJwnZCFAo0i+Shy/QWlSbzp/aPv3sizfmRScAu5MHcy/ZwfOSCna
YV3N0NrwTaUXWjC3W6aApH1M3OL8sbPXtobBhLAZrAiY5WQ/JhSQayvdOfBaYN2U
zSNy6xDTBorP4PFS6QuUyPfclsJgPB75wlLSJ7Vzso/knHKOVj1u34KKSvN0fs4E
oGEMAVrQpPEw7egOz2aKD2iunDnjUEheZKviUJ+bzMq9s+10k7gxtRrjpMlZUr2m
0LemEg5zzq4mxfknDFyaWG3qdqVJiJQDWubZEksVnvBCtTM5AVwj6CrrepOOXYCx
KCrNdWtJZNO4/4T+SCjBLXPVwFgWE0LjAwMwT6zYIIFYSyUgcEt7U0duLJUzX9lt
m90sQYWm9yfe6TT5c86u8oTXgyyukS8kN5XsbU5Rd6Ox0hzc5pKIhxpIVTh1o5yN
inhTmSWvJJd8ki2DSdifzk9JOSxTun/rmA4g0pz20OtAYDWlZWr5byJcEFHQ9gyz
6Quf79I9qEq5vIkrwV6e1gSEinPa9mxA/6QlmTR8v5RBim5XB0EKtR5p2wX0tY+C
Ir51u2+UjPCNXeDYTpCOQ57C56ahy3Nj6IvZezl9GZWmWCcyTaR2Yt//C2LWXsXB
4vKCNvcSZJPqoC7vNkqDvF/r2GqlUY/hSlpq6V18Rm4BPuqq4U2QFHCikVGtoG3E
Wy+oFXoDydo+HTSKR0KXfCDRTvaYgbESIAOkbMo9scjYR7l/xm6U2VAN0pYGLXii
tFdwrEnnh9xvj6PSK9fCjTOjav/plrjhwP2Dv7Hf9itOLPZwh/6Ej1eliMXzCmcu
fyrC3mM22c9KUu3yjJ8seIn1ft3un+ho4wLR19veGcLyfV4+UrB00uyDi1oljsbQ
5xO1IB+b/eXZ0N2bRLRcZpkROqBKHpIbjexrhbKAtm4eMQ4LwPioiFzAsRY8M8kf
pXwGe3OWdwMEUP5QDaAtgwBng2mLiSgBEQ7yLsZ8tGeAVcbjoJ5MmlVMFPezs85x
6QAL7diEMV1Q02qqbvPRiL2odLPRDpineP9V1d/Y3Jf+1GH5p+Ot8PYMLXvI+T0t
TQQZyxrYYc+dz3DZB97/UKtK7f2347GkEBfI58Lb31IqU+s6k15y+3NMObBeGqvd
Q5oXE5WhxCwsKMQd82o7So0JyQFFgmOk8T1CYxTs9S9tHSGEf+EtJitxx+1IPPqJ
B9T8D8vHOvW0+DIJK5IPSvXvkH2PCiXvGq3SDeg7XaS8DNmOYkpk0FRvza8RqQUM
AbFUZH3Bu/6R2Vd7y7z7TFXKUbGe7pgwBc7dz8JMXwaS5LDjnwTCORoZyqGnyi9v
ZL6deNrSm5eqKZzZkPFavnI9WJgvpdBeOAsjugrAtskhMwKjH8Bx1XydROHcK90h
UZnGR3qlXFQXsxBlcEtIy+LZW7WVyXnUiasjnXwMFXSphUvqoVxZRbsNIf32MHDj
b+6Z+ROeOtMpOSrJKI+80P6fuFL1uBr2pjLkcR4Ws4/+3bpGJAAbhSuD4Z5ZS31M
gam7zk8sn0a9TtHRXPO1sXOHBi8mWdNJooe9bPMwOc8Pn2o/IJA9nKAUfhoWy7GF
dZP736bNd/d8wTa+1+9Z3z86NpW2Z7OyRGWfqCFqGngMsnhtnGCkG5Fd0XAXahzM
45OTsulllCp+xxadJL7XbUdySgxxVl4ho5+Ls+O+L7gMozzjtE0LQ2g4u7jqICGT
uCn5ak39CZFYlKTDxuE/0jW/ojHrBtT9ICrZdp2HsC5D+rbQ2+lBMbQGhzT13T1W
qLLvv17dGIq4Ux8w3aoC7iKXMe+J6ZBfDQTsFAhI5LaaL12Krv/bMF320VrPH64J
b7+Pa4trB9lM0a+3+uD09rf3zmFRDr1GMvn9SE/7tAsKH2I5ZkMTVRgFFAcybC4E
ZpbDCvai3xsDi+tPHViDmksVvrX0VWIGba/5oHpQ60d5ZP4YQv7ixSjirKEEcjGs
cx0yUeNv2rhGgQhSWPppW8rupUrlC9sEfgtj9ZXjonpQYAoa0pBbfISZtZOz+Elw
Yl4/zPtM3oA8absS1RfDah1qIKCvlZX335odmqgap+O1Sng2XPJ+e7W/K8SA+XBR
8f9wB0PeX7E+txb+l/DqRTa2Q3jofKc/cf408aZTkyC3pHY5u2VFlaOembjIiy3A
w33Bvb2vlWDBobvtlqrKtq7uBnjiM9Ag3unM58ZIw8G5rKL59JjiSUapjECO0ngr
+A0Z/HNXzeRV7oYcF52yv7B9F7e1X1VClgFgQK4f8o8XuuFsd/hLXp7lMtJWrKnW
336rVqyKAiokNdM8fVBbLkTIgFBJn+Zs2k9dE6DfgKc69MTnqUJZ3APSEfahu/HK
a1zPwTizWYfQUytRwWxJG4IXGLSgVUs5jFFVc7uWCUa9cQbWOsZja6lSZJXMps5J
hB+pEWKTcZwCJE3S+kmqQmRhrNJPNMmhQiW1ipm2dG4YN0GdZTq2eoxd35yBZmxS
c1D8MGAT8Ltto7HutLazoU3j71/s9LLsthlWGZBfUIt0QvKR2XTtMRkKCjqGoeIS
9AVePThCtnc06VTLixL6XyZ/hytP/Z1+8+Q7OqY+C6B5OZSRJWd8kZhFDI2//6lW
nDYfvFOk+X0rGRMFcphz+w2YDKs/tzXizSARDhbwNvvbJcoNoX4bq0FyCPOsRMjC
UVANgQNfyHkX+M7d29gMlVrlPpTeB0nF/jWJRfnlF9akkETvIvTKAahin2lk0ZjB
fMeDC0TmA34fiUfvjCUhRSTAPC7bbZZvKm69wG6R36rlhpK680UaupJ+XI6NT+YE
DcE3lFSuIvAAvLrFDf7VjFjwN1CSuFi7yehTr05gboCtUp9pW2OwF/ribZ4WYGDg
7dBvYT3SSSVusCnsQHMY64D9mgIrV0NvNc47WLY4FSCqUeW+Bjxw9q5/FivdIEuI
vX1lTmzCweOj/W3ZSTh0X7Imi1ODJtUtDjxpPnVb73SNCAovtjWnDIVdEHlqvR5D
JTrIduzR51+/C6blSkgAQt6KvQZAG3DSFRSmDg5IFFb7592sX3B4t/TSG0Ex74zz
ZKA3KtNae1F7AiBQH9Yu0nXqopYt12BBbhN3IBzxUB9AxCZ+Cuh/NycmGim7x2Aa
1c50ySxfKy7miqiAPn8BJXcfexqLEG+PZYGB63/3Rdy0ZFRAwLRDsTSE4x3sAadr
bcxg4nqJjd7u52pQuBhTRMBEBP1QzYJwHc2j8Ca/5BlpOUTyDbQJxAXqRJ8HmZts
/ot/HKFIbfAiCfejT2rZ6b+TV3qgO/hKk5RMQ6btc8V1oInZ00W5hAhVke+rl/E1
AawrdIbklkxRxFufu7gv9fWy6/yTilP+BTXhPlSWYmFL8BedNBLdj7TWEx9qBDow
tqkYXPe/0Ikvvkiu98rpXoqgqQ+7is/dph4RhXCEpl9B2efXZumxCwvGHugPWV0S
jSM6HKgWo39ZJTge9K16+rgTeX6Z6rcwzMY3kiJCNhQdUXo+ymYXx8EkR717WlJd
07QVZxU5oKyzLp7SEUTks/OT2zGO67si1As/hKn6QQtBFDMa+pj2ai2NmFs5DLeh
4QVkPP0nPpwraWtsMQ7qvD3IOlpLSEo7Bwtg3yok5lkQrYc1yV/rrbA9DNa7MTHn
5kwriqjOSCwU3z+/rbg1Lbn7P+ampGE219ze32P7e8IQXWKQcKRj0L9zQxRoZwKJ
UMKeEAeu4k9JRjMBQEJU5ZxtbXs8uAun4pX5fWQSZ74rMmT1e9NZuxmirmymXohg
bzR8+6zF0a5AILhzVVvkMRYrzXXLReruLDEyJUlRYmUrmFZra2q6r2f0DUKUQkeR
8jAaxAFBPO9UZwqqmjAo51BASKfpHpj+C33wQ2NbMk97B/zmgvke6GK/gjOTnwKW
oGJMU++xnrdvnG06R1R8Oym3SiV8byKsB9ufCTsykeYcLFTeu4pbD/YuLnBmWEsz
wDLWQdVlC5pdsuYUiBju555nDeI5TNRoDNaCoWutlOsKPfR8e/IJjjQovMSzM4OO
RVKlnRTNPq1AQGyp9sZcIfJ9yfZbjxWszW+68eNa20+IKXkKhIsKGl7yn3BLMPmy
Ga11Ng25ewDq02mKqYB+VBxK8JnW7QDLm5nfRj8m+DsuWeyJH+b9kn5YIHdaI3Ba
9UBQ2mkw8aMYpPiCUBOsIEk/BXl1J1zP+dc8x++rx2z0K5WrOhFQ/1233wWO+ghk
5xSwXHjOht4M04lR2d7/QFdEPLY4YPo9mKzF8hTYXBQRqM0Q2upbPXQE3nUFSguf
BKMWleq9Hp/O/+mBK7XJ3MERK1UeQ7rX0wDf9FKgm0+ErK2hAXVw0/w1klmulQmZ
grEcWjTyVDIkCKkNH0/y4rbYhTH085cgH8qcXrIQWxuAnJa8B/74aKxyxjIxSXM7
M2fFlAhT+lAZipxSBOu+Igkf5BhLXAXbvNEOp7tkcq9ElIwoqHGMZNdLOz/GPU7o
1rjwnpfMKDaTSJg7hVuOPf3CY70QgBJopxTR055RD0bB+G9uSP9fl9fl/7JAZEBx
pLjjeCf5P5V4zki38DEkvE+sDvS0outXWlqIK8WmR6kDz4ZIIbeoANr1wWJ671QM
YZYfH6z2iU7qZpZQdF8HcaZG6nfVXO0thkRNO0Dkvz0w3foXPX/5jrWpRS+fVcLm
N7x7mKa0rzAB6P2z34VsCEqAdFg+Xk+loYLNmEuFam6a8fUxNNEQsHc8FspmOunL
/ZD8D5pOk1pgT41BWRTTajLc9Nw/sxjxnx7e5urwtY/Vg0PXCT3vvr+KeGt3nhix
37rDyLhP4DXpr94haBhogfhvI/58LJ34Pgy6/oSmcKAdKb8Kvr/NggJWpqFv+xvN
C6rFnqTlPLIWIGy8CyEItzVDtzAY9bXmR5eMEme2G1JzP/Dy7x+Ull6p9uKPWSoc
Q25OHvhT2hqHVwj2BI5Q0kuK5VxjewpHJBx7LPy1JTc9l3l9aBRu/kyXVcJ7fbtf
jaYbtJFR/B3dubLkYKU/wuPWc8ZDfxs4ZhDTq4UdPboENKQmK/9WAKjdSAhZp5jS
kMGvnU85uOqSaznbTX682vl5GMYpJMZTWO2GiVnc7KeeUjr6AMet2CZ9lOiocCqp
FmNkS2fImnPAmH9hxQoEBOi1pJa6YvA5i4B/0/CXiaG76ARYRqNFnFKg9vW149Ct
B4dweoYlKgDHQU4RkqLWHqh+i6SeNmWtI3SUsvZR9dhRSsdwLa8IpFMXRFLGEapJ
gs7eNnw/1n/ammcHgBKmckOTQ2ajYHout8swYO/DgGJRBeYUXMUyxEyEtJRsbBmj
B2MIUlmvZL55hCtWIGYQIz7aAxKwj1h4G3vYCpiob/XVQ2nlHyJTzR1++d7SMa3U
H/7KCNs4xmVd7uCpAwsxKR/0TxX5aJAogUJkHxia4gcTdrMhk1CjwgkJiICHncJF
AZpiESbBJXFc5oyZywhqVT1XV5brQCKncyqp0p3VAAb2zHn8zmGdZV8CV7wVDYNf
RD6Q24WlVGNXILP8Ls5Kg9CFtoTXtEhYsag9GU6lhEaOAJv8yvOfpXm9Jr/tVjww
IXqazVEKWbQl4/HD+z1F7GOnZ4pt/w9Aj4qcHQMKlgdkqFB686UOKl/zuVJFEgc7
dAExDE+4dk8om95DRysU+0c2T/2WrGZckm1RFvisLkcLa/IiyWjGb18dOTnXsD4B
yNl+FY/1RfizEXjldbgPrcitlvVoWify3B6UYB9KWmZlmVWkHhS73kUfRu3tjl4k
HURKnBjO7/mXUu61yed9H43y+/rqWpY2Lx3JAf8kL4tXkWu7Nv5mJFRIszQ/1eyj
rarauzx/Ux0bsL0axApXgEC9fYf4Z9sb5PhIuG2iBVEti4uytKXNlKkevjm2ovUd
bzcxRIbvIqtfILJpE+rL7Pm3i2+UxG9+emY9Jx6Xu6ODQ8Oi+Y2FY9stuL1hwUh9
TMr2gCQcBZ8mmo0HKY/N3AjkOFbeE5rO7CDgr1yGxFoyzL1FKVQyFpWYt0WWQ4Jx
TGJDkC4k+zOs7GgkP0Ujquq3UBlwuCwZFx0jQL4noM7o8GPFP0xq6AQQykimd4vo
XS7Pog4PXveKMBcAZyQD9kHfvfomvidP0+vxgR7JIfhPG7erEeOPbBFEEgJrlu+s
giEdM6hOdhINpStwW63e5vAZ4oohQ6Pfxemh4Fx7cNtpaZjsCp1gh+/B/LORXPTr
b6B6su5FxCLrevvWsOGXiZES+mb8WySV9OP/YDL8JI9gp5I8D2VpYIqPaRKGjF1J
kZLkL7G12iFc7drO8AK2OWWhydrxSFEsEJ3/P21nKflbMuSEiXnq14YBVK7CBm/3
fPFc+ou9F0qvGeHlsQHBJ5ZwyrWvWbYmxDTKBmuHZw55EYW87MXoEEML/JVLt3GJ
gNKx5CB1L3vP7Lt/EYHszlVRV/IP/wz2hcZbxi7AjqFTEdWmEi/1WMh5IBnFf9gL
JKB01IPwEm0IjEIXcJw8uil6QxyXLpGeGl795/V/INg3f09U00kdHwn1QPRtVwNq
+65vzROzMiK5zKccLSVF67BQOaNBnJ4OsBAaZic1NJdGgCxji35mOetbXKfT2XHC
cbpsff35ad1E4ZE0DFcvBoKKNK2N/mVay9wqPF1uEpc9fdoDZi8CIcNvV4xP/dFl
/jQw9WhX9ZHlVYiVBgZR32Iijv9fQrsRxQ1Lx2cd0qmgRaWK/qojuoZx/0a6tudo
bEO8WMLgl99m9Pn2vueK9NBdiYbiXRA4l6mf81i2+5LjoU0+D6xqnlsz01CM9V5c
1dni6VeKARMu0/VSP1xyewAsUXS/JUGmMvRJ5z7NP61XdQ1bvc49DHmCkwsF+LLG
vUAFG6vFTpfZuMYFZ4oqOdnWCOFfMp608CYAouZLASM77UF92KFSYB22axSW4/kw
4Ke/BO5i6PsHGxnP+X8GpGugY/JqzAesDPCOXgVru2pVQkwJttRwR4b1cMDngZKM
vGvS3lxKBw83WQhVzF3C+JvOujmwG7tP3svTR32SbjxjQPx4KBBQRBh7TIZI3UvU
pVm7zbfCoMV5Fxudz9NqyGGQvyA1dK4VDDuBfSo67kq6bqBCPul0QBuDkQR0Za7A
YfVCb2CwHBGoVTi+9c7K1ZfDYqnjq5TE1HNrCqCrt8SgNLhqNAftc/Dy+/sckB44
OSyiENLrryQXtOub+P8NP0GV5CUwdqaOLRpG0MNm3vodtETE6x96FAfNR8lc8sTJ
mU4WaIGP2W5eX0d7rO4xOAMbJXeI+TUuYypUxSfk/G8ybw1dP2O6pt/aXg73c0ic
NYNSPd6GYBZbS/v2H1A2UWY5293pj7DYpDixfex33oNtfES0RPkadlC62aYPjZiV
dAe79cPbdvfhTtYkCsg/lGKHQHF54ZKwx7Ub9f65FbmR8GSGOAP3SgDjs1x2KXVs
1EgSV1sLHYm9ffHzjAcwmED8zG+HrchwWTgVIUnpJJd4HymFNPzn4SeOUmsSrHxg
hiYFn2OSfOe9M/WIg8J9nkPjuasfsxA/QrFGGLjtYLmd482GZShaF/4w2ajN7SqW
JJtROzNIf6D8u1L1n+LEfSZMOTq2JCZzWXNQHsJADgKP8i4LBY7F/xILdXc1aWea
PzqxzG2T7fg0TZc9NQqT67fXHZWS0prQmE6BR1bz2NUo0ycgI0YlNvspoABSvovg
/z2yiCESLYBA3RadNYmSTdgqUS/b+SIfet/Emza69bPt56u6WwRrrYH70xtEy89P
QMLw3UcV9lbkvCyyjXtATMqcL5V2/7Mc94xt7hzp94lOcYE5gENtxFJFZekqExrY
PTE7ogCjUWdHEBfSviQ3YwccRjkMjzM/Ez8FKAfEOlBC10TvmRGLVv1Lvvlchk9p
DC59Nl7w9Ev2BT5NZJh93T7mDr4/MdNjaEuaYMY+U6ycPJErax24tasabwUGUrdL
YgzwJRnllySlxnNBvZmTIA2pffXr9vx8bmghKLXJVek9AMIglkSsX4DeqDdmavv3
eeTBa399r9SSt3XuEReeEzk/UIi3vgmjeo7jmLUORdUgz6h5nhCEGZ30pwBuQU4X
GkLtC9qTM4YKhVELkt37W3LULmKZs6EJaDoA3WCuXdmq13hQ4YyFXki7fSINWpFd
DwDn4tIJwlCw8ckjBICPlMixEdcVjY5PmFyrXWgOKpC7oypXqNtcGq+3mGy1tUN4
b9yWG66NxObpudVem27iKeIDv4dlrFZtIW5d9pgDM8pJqtfwceecc3cX6SaRl/ZK
DfecNI/XirFc+oQxMh9oNoCZSxEyyrey1zqJj+jH3ubdXBpe+AbfqrO2easjdgx6
nkYmIzJhGocoEkqIyznqzpLLgQ96bNDcHUtaJixG5o7/6N2onynN4ln62ASDqY8I
uN9QAGNnlIj0BrFPvHJD2J7qr8sLdMJIS/CngVkgrkRLtSH8oZDfzMbh8P+Nyufb
Jhz8D2FKDCCzMPfZKkLKASjvOcl5u6WD97ot2E9WBwutbWu3ouN+KojQGBVazllH
to70vgnI3nqR+xPism1cKw==
`protect END_PROTECTED
