`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yHgnZuT3TTIfmD9yv0xsRPKThTCj5omCMfY9HlXeD8AxYfw04VzJpWKA8WGF5NCE
0EhNxfxm0cAOnB15DCASDmNYernP0g2CS2cr6tL4p9N+yEI2kyrek3vTTD5OcHn/
1yz7l6l46jP/P0VnpJp0cRKLyjcfDwQNRy6lOBSRmAlCluoO4jNa1ZvXt3I0w+B7
iD7mnW5RTWtDWWzYEUAtyshmq4UqYCU6jNpmz1GW1p9Nfaz+KkPMjVfspUct7Txq
a/pIL/KVeU2NWPDM4KGeDM0+26zIarTQLl1oo+Thekdy2LCUwX6Xf6ttzJ9PC+h7
04h1uGejTMumc5Onzo2RJPYLiHFfHrz0sPtBJ8sxIML7cfmfRbeu9o6/E9hWY0j8
`protect END_PROTECTED
