`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F33RYUulh/R0PukI4c/i3QOqfYogbQ9MRLnM05jHIxJ9Z8cVQxnd/4OekIU0z2Lm
HNcc2sPST10Z6zj1MF4fP7wLCs/O88Xjb2PwcPau2rHRBiVItTzrIeKZ6vRiZIkl
AZf+lXTh7ZX16Lxm6E8Ibq8yE27Nwozx7Ctf0doumxyAWd3IUhz/dUG6hk5PMKxW
8LDI3/b787JgpkqArp/mdDsdT3H2ifMnrWcq7VM2IcygUtYpnydPodGbcgqXMEG4
WfUEsxxnRUy2xSQv45HNFVgntk/DsXMR3X87Jnj27NzMgdo1kBa6sULjq9HULfb1
dNv+q5QhMrjn3IYqJ42fF7uAKoSIj5QCfLm7qNqEM5+/5NxSvWIJodf2SI4vWkoF
N9Ktyg4GPTEmYS8XmdfwA5m9EXuEXJ7g4IAL1cHL69I=
`protect END_PROTECTED
