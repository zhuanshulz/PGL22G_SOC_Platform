`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e74sN1CSEmnvfB65vCI4PCE3I0L/AXR524R/GDsKsL/8gczg8DXjD2tNvKs8vA9R
CWPPn6gs4YHzVU0yhuyiuyM4oSbNIHYaqI2cvJtXsVlvdU8uGB9Nq8ho07MouPCx
p3eWrt+fS2ixmPVpZ20IcsXJbHC2ZCavvDl0vF31ut2maGcYiXIZE9z790ze++Qo
Z1Y+SEHJz9Wko6+mNMOFLnjupzT+8SJTOEF17kNOzdExX+3MSl198b93qM1XE50N
XvHSHhJPoUGykNkIfXl7JpJwnx7E634aAITuSPug8LG5AI6RSpk9ormr65/L/Tqr
V30emgsdnT4suDo0yA2ChhZeAM7HiYGeDPeE/pTzAFCkYqEy4PPiEf4CAiZ1HYqC
03B57pVKNw6rRC5h7gqNAy70q3Ro341gHLvz7vO1Qj8KRzMt3B5ZBs7+cZ8e/4NZ
0iEW38RKyBqe+mZDwzpgKtTzc/OcCmeV1BvCsuBpvyLooZ1E763rrFlrxcjJt4dY
K1Q3Zmfl+BajGagvQEWxjGuR6PrbJ6lD570GLWjDZTNtSwYLimo9j7tEWuLd+Hh/
E3izYZGM+nhDIrjOBOuWWjxCdO51ZCZNAvgePAFggDqFDwNDLKs3sqt4tMUexQoL
Bmk90YEtwfdDSPo19E+ElVlrmiNioSkw6LT8KaL5cmvjCR31WcCqkt+fe1Ne9G99
tLMlX2bzMBcjAU4q+8kJChQQu4Rg5n0rhQyUASOvArY0bdG3LjVNBoPJ2IGKvV+h
Vq+r05A9DBILRKMZ65wMd5/jYkMz5SFLy/d+RwJgsD7oIW3CvedKV7KI7Psq8F1K
Pwwo08bisC79D00uBcPLG0GwyxYiFNh/F1aEr8GeC1eyvXYba+4XsdlqV2NgOPzH
hZvIobG+XHdu0/JCdSdnc3fY39JUSqzkt5LpFzhQk+0NDpSNDi7ammlLZOHAkZrT
0Suv3hRgs0mD2fXm/zmgna3h7Wbtk0XlpPBZDn0FxFRmNd3WvjroQNwnV/5tMxOW
7v6JJwkVhXYo2z6WZRrHl/6H3eGC1+jGCVEw1sjkoOYpLgHhGDL4pv4cxt/kVnRm
XJg9LVxE837pnwd/KENDZGvoZz+V2g8o7PolhB+2R2nI+6S8TuipXCVFKbGUBEAz
aAe43ckPTFCydtpDHCEqesK/+5fkkUzXJUqPTwDb8hjDAVqlzJX1MUsgfIoBJiKy
mQZWYCKZQhzXiI9k4j2V7qGZyZoQw4FvBBZ50YuPOjqpZAyysZreAgHu0pm9GcoU
pw2RWzp89xswtcHqpSw/gZg+g9m7Kk3OvIRFPiiY6hyMzUya7zSFMdOQZNvwJ1O2
Eady74Cv43VHuNtiMLqNQIddhQ7wkg6a8VE5o8UuaZtMi2XihGDwWcJfOQxLrilq
tBOIPJB3MsLmNcfn99qGfudtJAXjfEO7d8MtTdX2tRy+8uaDfNmD7dp5rIXNkCgM
+rrF1jQqv7obPiiX0eBKdVcE7AlMfxETuOJDsg0btayUU60W+0CAeFwAduEYe4N8
4p5KntEQW3QfzN9Slzz3rDrNtSdpZRW5wQwpe5b5470G6u2hdlKdY/yTjaxJ7iOi
8qjeOMAasWRpUax5FS7orOZrsjuVHcV14NYNQB0ZpZml78jbbzsDBOQWF9Qxbt6j
woHukJ+H3+yqIof0QtiPFVk9K1L//9c5Vsp50m/XurFPOPIcBvDHAEUBP6DT680O
hRt8R7jLxjUx96t0caG0nIXvrykY5+lzybpJqdb+tLahwRQr7bglvDCgAcAPokBF
dziZKOCsI3asGwK1Ips2JSIFov5VqeUrJoSTy1Tyw4XgrtHGsBd+tgODXNuUuA4P
wc3t1jAkJTUS0SLo3a+OXlsl6ux9WzlDc9jnZL9fH2miBD6SItRX8nAqY8dW7p/Z
WF3bQKQhQYpUDnhRT30Z4aCvUgmN9qRlqiYBezmKALs/Vmds/TFBCEbJApD2hiZd
DM3sEMStiJyqb1Vs06gVzCNHhCUbrn0WYRAtiq/zZ9BRefFlR8TH7Oz+P+soU0XZ
iWBM4qZJDfGvFFUG5DE2mYm4nTBnVsGnymJvivQfAsoOQiwSPp0UMzsb0zfJV+wF
sj0vZBSzB6fCnHGM2pHAXetPDC+Kk8tkb0Wq2sV+N5+JASxGrTSBvZp7VFNGdr5I
YgplPCQp9XYiwRG84Ra8enEZjbwEkiMaqRVJJZn+k78ftHXvxXQlvCJfwg9EnSDQ
E4TTgDngPSVjbAB18TCkxvgBEkE8telxhL39VfOy3WGmTBr07do6o5NjxHZ+Q3b0
fdesFb09X3G6poJb1/GC94/nAe9M5DcTIGk9kW2HTn9NdrpMPl8RwVq9bCHa1mKz
8mkMmuBSX5j11bBDkRqZAzndJPdDRlZF5CkUtrg5CLoL+RhfqdE1hEyJqpq19lVt
lS0OYUvpYO2gJlphRVPbVs0C71WTiAC+0S0OlJUOb8Ah9xY4Vr/tv8pWF15rFmMz
8PmXHFjidt4vqvuYCE7sLBXQ/HjxWEFoFYvr2/j/K87wzmNMmjZ3bsbI1iOicat+
Pomeh2eQjkK3/Y9F0taIl+uCqwy2c1d0Q8sdxd7vdmNrA6XkEUCDpk4xgKZjgKEb
5deUoA/1VVz5lRvpen7KOxgcEiUjc4lGCHePVIXNByw+3B7B527rqVGBAH9CuMOW
OTyMtZL8h4DqUt56hK8z2Im7O6hFOphv6QOsX87/CK8s82kZoL+Jo+ox5Qe2oq/T
MQxorkvXzSEdOjj0e3jN1g5elwV9yRTnMi3RacjZoj5HFYvrmPKc+hVXKH42GGMJ
38kpuJEWYJTvxwzMQivlxgBH4YZS9P5+99XdIprB8XNBWLpyfSrOuyx1Y90fyo6I
5iVQwBbvMqHFnX7GFLsYO0f9daFcLW1GOlTPRucvp1xRYuOLH9jE5qFCfmpjQ7sF
6BQz+V7qCgBeFWtIZz7bOE3vz0p65DSzyH9j+xfwt4daXmHYdOh9yQQn8CnWiXm2
hSYktkLBVrsfayVcLsJ3IN3TfdOdRQG/U06xLZ22yN2Peyx3xQ4NJY/NcPce0wFi
YblQVNJRxSyP2U19c42JNW2GkuPMF94iIIdKBqRvcfiA16qVTVOB8NLpUmesaR5f
Zf7wa51+Ehc4aH80KZZUu1YOjIbv5sxRaP2PVeRS63EACjaUquPolj7YYif0QKuk
FulqVjZeVQu9wXgjUfhyc6J/4xhB5eLKekf71KH0yT37TlvCRVftIrw2Ra9oibjd
fKeGcT2grEzEcI+TzyS/Di/8yg7Yz6u5FjGEtxYRh/EnIK3zI2vhRLMM8n8yltTE
`protect END_PROTECTED
