`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xc6VVBBwUnHDZbUTggos/F/nJIhBdlWCIkNxRQcOB0Lgc5wLMmvGEsGjDsjURA/3
vtcRBq7n7+iBURGcZqSnA6DaUepQO5JOWMa3wZjxZiCb7qPhhb6DGTvFhBHCQz4w
0wZ06btl7TfE4mES9u1G0tKNx4/sSzHb2XeehY3G1iWsWhd9VbWiujBOZo6EPV2/
Fj+FguzFD/JzBYchwkgDxPMwph7f2pbLQYVhpm8MQVHx+c9OA1DuYUG0M1CGjaBs
d0wvYzS+ELVXAL7MQqyzC8XuOdohd2k6vJaI2R/ezFIbFBFdIiwmJEjLODApOUaP
v6B+AB8evJIQhaf7/G9dp3RJOpl9LnbWw7DRAqOjd9rAgXuv4YzVoRaaxZUJAV5z
4ORHdcl5ZwJxu8uqmS55+fwpsU3C03doYm28EXqTC2g/WlcQRk7lOsSKvNU9ui8a
+ru2tvekfAnQiSNqk+xMCPK8CPnLo4cpBhBF/eeuXmkybxlR/DQuGQwzdNdiGzd+
/awxNWd6y7tzA+zv18jWcthiYl9A5Y2cyDwjMJeBYRNhLbhrlx832u+fIMCYeaer
eCKUP4NPjYvH68Fz11UoBBrC8FLh3BHMHw78gnJTG1IgQrfeQL5wu6v5sxIOniOg
/uYjrKj9QKqrT2uqGGoawm2Miyi5od19ptPL2ADQKiv+O22V0bKVhlFlXjguDjvN
NUZfMhUH23jzq+CfK2OuovaUJcqvhNYE7hRjCal2JfXKIrjb39s/uAED5/ayPTSn
/Y9sBAsz7EW7Ba2YXqzx3ggB1Z64fD3mq/+DRFd1X5Lxv4znVVYwlB35WYPDsU4V
YcPVf+6kY4/IRRHs6q5fWM0S8ExtNSzWiYUkhcGojFwv+rW75ECxpFgnj5krGLfF
lF1SeXc4DTCqJ+pjoSYNr0FglecXYzxX7vyMWpp6d61hMxbMt1jsW5t47Jfxh1ky
qfVlge7rmD3KMsVvOTt+R94QpXadL+0TkSqCM9lKJJ7OxXo3/nsBeJAVnNdjnyzU
dSSlAWCW4TkQu7S2ZfDmO8/PkjxybGTVw2muVmrTngg3GxgaAzgMTG8dDAV4AHpQ
zEHibOuGxW121DVDPRS0ltTIg/mLd977i7kiHUg772IP/yTG7SIkGWyRQEzB4QGd
SXw+C6dDgQjxK8tpntmJfw5wf3XMPjPHaIGxbijG3su3d82CFIm+D4rM7V/T8Szg
y/RJ09+PD0WnOK4BME87H6m3uuy1HAPpn8Fqf+SBw+FhGTjmubi7v9iOMmAal0UJ
`protect END_PROTECTED
