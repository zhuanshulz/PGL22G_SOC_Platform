`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nPW6LveV8RCRQW6k+M+n1zLbuehgYeBhKPsH1Qv+urp7h8fVnGl+H5Yqdpdl6AVT
9FZfdFOTgKfySBx1q0Sn6+Yieyice/a8Ps5gMf22JaHkUzMKCTFCI5pEEGj/9nh7
7hao7EvhS8JNmd2n3vBNP33WUVYOIHvgQ97o4ii2ENw+ca2IUvywSnSgoTI+7HVc
Bp8EGBg6/NIy/PdPjyk2jUWqsrbeMVkMzjvJ5aExpg2dH1BJQxnsKfPLqsxt2O0z
UPA+dNCjHCTK/SqDW5zY2seKnMX/OsJ4hrRKDX2dsasc07WV3u2lkm5YHolO0cpK
VnCsjx1Pjgc2yrlvxNkiygTyzh7GvJ46dGDcku/V5XITwl/AgIb933fY72nIDB/Z
pclaZqzb1tqlBXeHuLwIrJaDLhhGgMBq267Yv2vVyhsRfscJdILpzaEc5nSvKDOs
uysZJJb//aVTq0PC6XRsXjSYJnc+ZYa0zjK2cqOfprf7LkOFKFy4RGXg+UgNgnbY
plQtvJfKh86ZTaSnE539ar4XKdw4em+ux0mBElo/CeRNmxqkdI8Ed3CB81xGFHsx
Jap4nhS8DhfG5hDvaWaNOHLVEpKfUxSbaZKYNGoDSqgU2lxBO50IOiEByt8pgH79
3hzkuON4BjkpDC2XradCc104gir3xty1I7xLkuq7XdWAJA5yXF1nLerMuqRX/rh6
kRMcu1qY5pVynb3BnrDC3yM8QDDi43oLkf8eVU5rRtU6p814KetN1avI/mTpnAb5
7skgzELyt0ffRUlpV/rN/DTFrsuWKfuEasp7jljuLtpVKBiIezjT7q2wz8S2NfG9
v5fWXY5qfkPorFDwv+jnB/jlYqPgGc1mocWNpNbU0mli01MJRWjI6WIMn1c4A0HC
XVeJl/lhQKpr5BDj0BXwf3K9o/X8c7el+BnEvXvB8PlRZG89PqiXcYaRut7Nl8tJ
RU03rnSSXZFAyeWjtomX9rYQWv9/V6aweZuTQ9Lbw3oDWUpebDpiv0pDbMOU1iEm
ETd1HhCa1U43ZCL2oMDEyZWBFwI5JXC3apE/fHkJ10mrQVlWD/Zq4hpXLSDYHJlh
`protect END_PROTECTED
