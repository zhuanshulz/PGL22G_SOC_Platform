`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vjW66W653LV/YPa+ad3U8J/5P/vUFmbuj4nZVMptseWQSNa/91t6hlxTPojBgokc
ZwUzTofW9gbnWf9Up2u4iNB91znIT3zpTGN/4AnhbSOcjk1VeavjbaWMYbX4XGIn
+B7iKnNgAiiAmopMHZRUaSjEUxB4+6j088Edo9C/vvspdyV/iWr7ZeHYfdIgQCZs
TGVcR1d/F7a6Nj6eWiWfEJJesyusaj4CcOKEeAeK26HKhLmZIHO5oJfoIVcbIEEV
cGoJ8ENubqHlsIN8/H3kJgAyBuFspKvSE/W3iNIFxJDhWHUrE7WyJnOZ3TGASLxu
dMpVN8dDr2gwdLJPKbbqOpYDOLxC/dvDK5O2fmUVxKMFK76lYBq1ZmHMIgd8P5op
y57CVGuJ2drP5/Xe/63Ak1dCZRrcg9Wt1iYjDtOYfBc4ce/4313BERXxDOvh3wW3
iUIyAUJJDgPlr2NAgLl+YwJ8jJ/0VIYmoUJf3bz6gHjcNhtJtrQtplvBacSGtlWV
LHwz2q+xNNjww/Drwp4cKYdJ6S+D3V08miSercK8BnauDW3E6DBXxDs16XSVZ/TJ
vLf+0CuWX2Dr325dLZ71R9D51JaFiDb9tdBoPjFLN391H+v109Gu1gutkJ5Kg3Ei
wqP938upJ9Cg0S2PFn7FdJcZAp2y9QVejpTr8PtpG3dYASPByqmD6Z4GQsS8HjV5
KMXv2LQoNt6HJ1jQ5zd8Z11ctTkNPfLJkFWsQ4q14EfRkPxxq5ojoMc7818RbV3R
cKbluloqMdIlSTae0TtPjx9UqJsr+1NALFoUljyULRWFCV9wUmoxPACJPt3Lr27t
jhxDXapMOA/UnXqemS7/SEdoCUz5FTCDsOgWm4iHnhk=
`protect END_PROTECTED
