library verilog;
use verilog.vl_types.all;
entity V_PLL_E2 is
    generic(
        CLKIN_FREQ      : real    := 5.000000e+001;
        PFDEN_EN        : string  := "FALSE";
        PFDEN_APB_EN    : string  := "FALSE";
        LOCK_MODE       : vl_logic := Hi0;
        STATIC_RATIOI   : integer := 1;
        STATIC_RATIO0   : integer := 1;
        STATIC_RATIO1   : integer := 1;
        STATIC_RATIO2   : integer := 1;
        STATIC_RATIO3   : integer := 1;
        STATIC_RATIOF   : integer := 1;
        FRACN_EN        : string  := "FALSE";
        FRACN_DIV       : integer := 0;
        PHASE_APB_EN    : string  := "FALSE";
        STATIC_PHASE0   : integer := 0;
        STATIC_PHASE1   : integer := 0;
        STATIC_PHASE2   : integer := 0;
        STATIC_PHASE3   : integer := 0;
        STATIC_CPHASE0  : integer := 0;
        STATIC_CPHASE1  : integer := 0;
        STATIC_CPHASE2  : integer := 0;
        STATIC_CPHASE3  : integer := 0;
        VCOCLK_BYPASS0  : string  := "FALSE";
        VCOCLK_BYPASS1  : string  := "FALSE";
        VCOCLK_BYPASS2  : string  := "FALSE";
        VCOCLK_BYPASS3  : string  := "FALSE";
        ODIV0_CLKIN_SEL : integer := 0;
        ODIV1_CLKIN_SEL : integer := 0;
        ODIV2_CLKIN_SEL : integer := 0;
        ODIV3_CLKIN_SEL : integer := 0;
        CLKOUT0_SEL     : integer := 0;
        CLKOUT1_SEL     : integer := 0;
        CLKOUT2_SEL     : integer := 0;
        CLKOUT3_SEL     : integer := 0;
        CLKOUT0_SYN_EN  : string  := "TRUE";
        CLKOUT1_SYN_EN  : string  := "TRUE";
        CLKOUT2_SYN_EN  : string  := "TRUE";
        CLKOUT3_SYN_EN  : string  := "TRUE";
        INTERNAL_FB     : string  := "CLKOUT0";
        EXTERNAL_FB     : string  := "DISABLE";
        BANDWIDTH       : string  := "OPTIMIZED";
        STDBY_EN        : string  := "FALSE";
        RST_INNER_EN    : string  := "TRUE";
        RSTODIV_EN      : string  := "TRUE";
        RSTODIV2_EN     : string  := "FALSE";
        RSTODIV3_EN     : string  := "FALSE"
    );
    port(
        CLKOUT          : out    vl_logic;
        CLKOUT0         : out    vl_logic;
        CLKOUT1         : out    vl_logic;
        CLKOUT2         : out    vl_logic;
        CLKOUT3         : out    vl_logic;
        PHASE_SOURCE    : out    vl_logic;
        LOCK            : out    vl_logic;
        CLKI            : in     vl_logic;
        CLKFB           : in     vl_logic;
        PFDEN           : in     vl_logic;
        PHASE_SEL       : in     vl_logic_vector(1 downto 0);
        PHASE_DIR       : in     vl_logic;
        PHASE_STEP_N    : in     vl_logic;
        LOAD_PHASE      : in     vl_logic;
        CPHASE_STEP_N   : in     vl_logic;
        CLKOUT0_SYN     : in     vl_logic;
        CLKOUT1_SYN     : in     vl_logic;
        CLKOUT2_SYN     : in     vl_logic;
        CLKOUT3_SYN     : in     vl_logic;
        STDBY           : in     vl_logic;
        PLL_PWD         : in     vl_logic;
        RST             : in     vl_logic;
        RSTODIV         : in     vl_logic;
        RSTODIV2        : in     vl_logic;
        RSTODIV3        : in     vl_logic;
        APB_CLK         : in     vl_logic;
        APB_RST_N       : in     vl_logic;
        APB_ADDR        : in     vl_logic_vector(4 downto 0);
        APB_SEL         : in     vl_logic;
        APB_EN          : in     vl_logic;
        APB_WRITE       : in     vl_logic;
        APB_WDATA       : in     vl_logic_vector(7 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of CLKIN_FREQ : constant is 2;
    attribute mti_svvh_generic_type of PFDEN_EN : constant is 1;
    attribute mti_svvh_generic_type of PFDEN_APB_EN : constant is 1;
    attribute mti_svvh_generic_type of LOCK_MODE : constant is 1;
    attribute mti_svvh_generic_type of STATIC_RATIOI : constant is 2;
    attribute mti_svvh_generic_type of STATIC_RATIO0 : constant is 2;
    attribute mti_svvh_generic_type of STATIC_RATIO1 : constant is 2;
    attribute mti_svvh_generic_type of STATIC_RATIO2 : constant is 2;
    attribute mti_svvh_generic_type of STATIC_RATIO3 : constant is 2;
    attribute mti_svvh_generic_type of STATIC_RATIOF : constant is 2;
    attribute mti_svvh_generic_type of FRACN_EN : constant is 1;
    attribute mti_svvh_generic_type of FRACN_DIV : constant is 2;
    attribute mti_svvh_generic_type of PHASE_APB_EN : constant is 1;
    attribute mti_svvh_generic_type of STATIC_PHASE0 : constant is 2;
    attribute mti_svvh_generic_type of STATIC_PHASE1 : constant is 2;
    attribute mti_svvh_generic_type of STATIC_PHASE2 : constant is 2;
    attribute mti_svvh_generic_type of STATIC_PHASE3 : constant is 2;
    attribute mti_svvh_generic_type of STATIC_CPHASE0 : constant is 2;
    attribute mti_svvh_generic_type of STATIC_CPHASE1 : constant is 2;
    attribute mti_svvh_generic_type of STATIC_CPHASE2 : constant is 2;
    attribute mti_svvh_generic_type of STATIC_CPHASE3 : constant is 2;
    attribute mti_svvh_generic_type of VCOCLK_BYPASS0 : constant is 1;
    attribute mti_svvh_generic_type of VCOCLK_BYPASS1 : constant is 1;
    attribute mti_svvh_generic_type of VCOCLK_BYPASS2 : constant is 1;
    attribute mti_svvh_generic_type of VCOCLK_BYPASS3 : constant is 1;
    attribute mti_svvh_generic_type of ODIV0_CLKIN_SEL : constant is 2;
    attribute mti_svvh_generic_type of ODIV1_CLKIN_SEL : constant is 2;
    attribute mti_svvh_generic_type of ODIV2_CLKIN_SEL : constant is 2;
    attribute mti_svvh_generic_type of ODIV3_CLKIN_SEL : constant is 2;
    attribute mti_svvh_generic_type of CLKOUT0_SEL : constant is 1;
    attribute mti_svvh_generic_type of CLKOUT1_SEL : constant is 1;
    attribute mti_svvh_generic_type of CLKOUT2_SEL : constant is 1;
    attribute mti_svvh_generic_type of CLKOUT3_SEL : constant is 1;
    attribute mti_svvh_generic_type of CLKOUT0_SYN_EN : constant is 1;
    attribute mti_svvh_generic_type of CLKOUT1_SYN_EN : constant is 1;
    attribute mti_svvh_generic_type of CLKOUT2_SYN_EN : constant is 1;
    attribute mti_svvh_generic_type of CLKOUT3_SYN_EN : constant is 1;
    attribute mti_svvh_generic_type of INTERNAL_FB : constant is 1;
    attribute mti_svvh_generic_type of EXTERNAL_FB : constant is 1;
    attribute mti_svvh_generic_type of BANDWIDTH : constant is 1;
    attribute mti_svvh_generic_type of STDBY_EN : constant is 1;
    attribute mti_svvh_generic_type of RST_INNER_EN : constant is 1;
    attribute mti_svvh_generic_type of RSTODIV_EN : constant is 1;
    attribute mti_svvh_generic_type of RSTODIV2_EN : constant is 1;
    attribute mti_svvh_generic_type of RSTODIV3_EN : constant is 1;
end V_PLL_E2;
