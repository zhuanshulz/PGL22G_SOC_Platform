`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6mMbK8h2pQLNJPuwFkinsfPmsblO78M0a6OCWWa2xB9Pl0EWu+Tw9RLzf7tbvfBU
370eC8lcQhuJqjhV5mOpzQ3N4x92kvvOMBPKBXSOBIrlOzYymY9sVe1GpBx93QMe
fZ9nvs7nj2YKVieCaxGe7qDj2o5KL3S3GGM1os4FgcbWyRPxBp6BuU8udN3Q5djr
B+ebUZAPrvTBnFVxhuOGKVSoAOe3dSJVbUnNyB+HikWlE5/tRmnQqtUhJJ2XEzGK
6tRfQiWe1OuHxDAlvWhLSinFIjzliEbx73f44406UzWPtDJisYwQj/d+I0klK/FC
SnQaRBxUuAaB8o9O9u25bU7yNf9lgSOSIOLIG1Qw65dINFj8oeNrKgALUqz6CBgD
6Qomt+asQpqsDx8Hfd058l7nm8soMq2921IB1r17gRVVXe0bixYeaUXVidrruGSx
sgapjgqqJb6+1p7vh2iCs20ZkUafwSNhSkUO0yQ9Mexs2FXgiKJKqWQwq+Zgs8Gr
D0pZV7GVVBSJV45VV3bvHc/31BWdaGDNG1jEU7NuDv5MwqUclZr8hZUU5SXx28sG
OUtSrdwRGWXNKYn2vPld3nGhKCGTvtmZQi6NovkvwA03/jn+bfUlvDBIMlxAQgbV
O+owWKfmdDk7GXDPSAMS+C6ZBZyiwc8CMsWJJ/cMvcE=
`protect END_PROTECTED
