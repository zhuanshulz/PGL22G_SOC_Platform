`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b6z3+/69fPFhoEmpueF/9MnvTXgGzeu+Eutb/heg6G0R5KS0O88Yoi3GDL2D5gI0
MB+SeMF38NJPEJB4MTwGvZVeFop6ZdoGVb2LNoodMl/lEfWxV/xnBmOR8gWYBkkx
dkYx+07DLLBokFtq5PWzY7f7QFRPMCUoIChKjObO2Vl1z3ZcMZ3qyiMgrHkVQeXL
hWkgp8WIQj5q9/JQGLjJ8e0amTHG36QKj6lSbfJXCHtfubGcAdEmjUV6QQz096dm
rw2WtAILXOqj7eYYcNRFuJXcTCAe41uCRVQl/b2xg8+eXvxJ6zCSIle1UnynA3fC
NtPsWbmdofmFbOUP55Q3E87ELSBvUo0enHFWRprTp/YIGnaSicSxFjQsLF2titxx
dT6KeT3eDYVnAuYHBy22JO2vF2GwgebLuHlq3qIQTYV5bVsamN2wykrLNRduqUlh
ninCDFN1qHNTQgRfBGfXyZlYNHcpwwtEGC+ZBItGARfMX57afBSDMcsqrCCVFxIM
1M2Q+Ftml4H+av3ELJPbdVbE6S4Mwcel9xEGeeqWFzSo4B7KV8EYm0Ml3jhX18J+
nelJstCKAAE0P9oj5a+Dq6bMS3DhbYU8p+QZ1w3wid0rVZewJ/T1uZZmMx/qYiyL
S0JuHLXrFtA3UPsLeOT/SuEtS7YySIuM70FnL7haKBdLetqQLozzfp5S3Kxc/G2n
1KoBHAEdD+RnzGVR6fpif6BkAPeMikWUuJBQmCBKLAhVxeCeDS4uUa2dnE62xJAz
6d+J+lKUybQxzxo6VLhfvaLyQm/22I3JY0xPXtm+oVVV4fEbm6YWA6znz4nryUDq
LheVSf3maZZ7oexiAEJ3qWcnOMwF1PHHz8YPcVo4lfnbhHg6ncGAAumA0dDaYOlm
8uexee7Pi//jxEFoTG7n5wXi90gEC4OahJXcCc+YA5P354G2tsunJ+nQq5fjr0+g
I9ty6e/1oydQvt+MvLouiRLGdGzicYJx0Xv8PSyKeV//Gkju/o1fWmtzW3h5TDCq
VXjbeOActOHO+gFrCl25VRtbWtisOviGGCGmoUZNw/OURf0uvGRfIexsY1OsAAUP
sBSJWQAl3ajpa8B+JszQAeoRxzoi6eetBRf/wJvxcO9vsI/E0Oj1qFFxyXdyykRY
961REJONT+crzy5csxy+WpH0ui6Mg5eGXqZ5+X8sVYYRAkUKdlyZ4qHm1lvylDjF
rDB9BaOxC1+MlDhneYT3dHXtFixdVK1H4KO82HuY6E+tBW5g5M/1YtMyOSn5fvrN
ssnOLnFPa1XzUWNnzO9Dsv6HPmh5wi3LuYIHlNI29L6hsIrWfPQoi2J99r2OwSCm
cFCJw28lCelQZ8BPIMWDE3Vi3kVW5I7ZpZZQO6uBMt3HAvxcJzaZRvK4QA35+OQb
arulCl9iSPCs0ksKlgBW/suuVnLMuV2BWuYuXi6RBrH95Cadr5DC0X2D85fsALEQ
hU+5egeAxnVclSEfAk22uJOObX2rvjkraU+ebojxGqXEv7oE+mgXAtm4L6Yefr2n
W8+nRFK2pbYv+EpDlqOm9zFHt8MB51zjcPnRz0oIGo9P9cz1I8LFM1hC+yN9TXDd
p68rrQbAql5/O+YButENxENPa4pJOTFelpBGRc6ok6i9sQh3D0TnnZKDO9U9WJTY
WRNkAfHS1m58IWVg2wrLXQA7qmbEHId1Gd4KeYSAILYZhrUgQtEppDqmRIFL54Et
HtpfoXS2/EsybFq72bzbxlh0+Vn/HoCUlX0JI0tyNfY1ibJ9ovp7c0sQXQOIZ9ED
`protect END_PROTECTED
