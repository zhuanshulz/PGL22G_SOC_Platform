`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/6h6bzNUV/kdIj0yYUvvujmEMd4RW4HI+h2XSkB4NiWrlHmmUD8ZXrgiBIpZAFN5
f5XxeMmE/F7J6v0YL2BFyjJZSUdu7L0Ztn8F+zsqetJvCihdEe+deP2CHkq3qlgu
Hv6HKrQUNJBLItbxc5E9a8rELGMw+9lgUMf/jYn+CZqMAIVDgFmvphYaA+j5dKki
XVCesGoHP5W+VrnBZaQ4SpUG4hb1qGoTCj6JU1oKgLkF9bd5hm7OUQwSqP4+D0HB
lCG6MIei5FpkqIapguIY+Y20CN4xvfqbg44VYLZzMjAIK7vtNkykoT4QVz9WPzyl
VBRQWySJivJhSSSlE9Y2d9dUk18UdDDom5rbM0niGe+8CfuqemX0FznAgXpfd4Hm
s54vaF+bDSR0YloheM1Jl735COpgLzwYckQkQNOInbo8T11RO9BNgJgsZywtSW7h
B8MSSNM8CWnXnBFGKsvv6yr8sx3VuI+zAky4UzLDU4UvXdKNbRJTG2Q5lqbBJQkg
+IQvI01KCQ6IN3o+86cLnH4E5P7iQafes2Efb3dVzWgxBnGld6eUybL2X2soHIg7
qsR9NNJjR8mGrg1s55JnpRUSTaIVtoZfcXWoeC3hC/wux+BxfY6fsWLqg8mCPu6v
Z3mxT/3dhWJcHX0+BNBrwtCo8gm/AMepVxLTmgY+tElDJgl1bMlEkwfVSyKNAZt8
uBYR2CyikrcXiJVzXST8cfpllhSR8mD8MPXpQJE3k6zivWJPsSOUanOzEzrYSUKz
0mxfO/jyQhN9MV7u5zT34Af856il5gJlrV/xUBawYK2WY/8kdb8se7JyrFa7ypSS
`protect END_PROTECTED
