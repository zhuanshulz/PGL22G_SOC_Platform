`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E8ibJ1xuqpWT/kpZI3qn1Mn3DMY+yxFl0CrtTaRsTdW6UGmDVMShNiwVtL/aHdc2
aF+28G+7OVMxQfg7osBgl05FqTYIQ3YXmQS/v7lk59mPh+nbHBgGv7gzhFZ+8WZE
gDJeY65BdeZHytjOtZF9PBuT6wf96eqco5HxDIYvQrKGjzHIWIesJL3Aki5nD9fg
I3ooldBZ20/TIaIf7HIK+iVAlnxji0QaLWSGovN4XwA2B1hc8I3km73R2TUy99GH
BW3AcQOn9ISVW4Uiy0wN0NYvSK1OUEqSOdtPrjPQa4j9wNSL1gzsXGgJumr4jFRy
sVQYkm0+tPkvXupcwDk/bqDwzKXUjBkg9qC+Rb9TaSf9KaYGlcoUnaCsmc8mDZZX
wFGdYlTcBf7lCLM3+lOIOR17W/YweNazELk2iX5Wta3dA65GOXqYj/rLjGF0oBKs
lBB1yWxie4Lkz5+/Z77T5NUOYnCMvm+5MHqbh/hgDD5FGh5qOCsilNSxbwgHTDw7
sJI7UhXYqMKdzSoh48wMH2flMN+hcVc2D5S2iF6t99QmDbeL3f/Cmfy9CaklkT1+
ZjdDpyYdrLzgjukXLW5XTIePTW5ddGOIebdW5ICrq8QvdqDActJFMnnY1+vQENr3
Jw6eqiDm3fCLK4j4SDY3lh/F4xBxNXUkzqsdN1ro58qK2Pmo83PBat8ec0MTmSzI
p3ihso43JqAbtf6j4j6cIUoEu+BwDUcoEZ7TM8TV0ttghvGn5s0LZyhwMuM57do2
KOp3zNWiNZwgxOElBy7UGkDjYJACw5KpG4Ae9rN+JfjwPXCoYbOTMLd7dUtXnFD3
KyLBlHiu92DTbJRu26xGh+ABc+fzcYYfGDHrhH6aDkAoHAu+UviM5CR6Z/uYQ21Z
Qf6/F34Y+PBrlD2OK/1ztgLUqwneBDWvAvO/dh1UvdENm5CInvSYeK2q8yTEGkET
pqnrj3y0YvDqI116oENNPV4FF4QujymaXEZpQATkF8ErbrIlvLk4sOoKgjAQmAny
GjIemQw+GM4Bk245PAOuFzHT4cFuF68AV07zo+i4f/VuBklKJj1ZzasmRo+74i3o
JlKHrpm77zhnCThiuiOeQ9IwL2STsP0uD04SrEpsDlflZaAdEztB/aq8vCd/k5SU
zHdgoST71Qss0K4vwsClt35YB4TLOS/tuPAfnJLXyTlOB1p7A25sD+fYiOv/sl4m
dIofGTsBdgDWj9pADKxml2zb/iK5Q76YDT5PO8wO7EPC0A18SL10B53NAdy2p5eV
uUiRct+GnSyCWHVR71knQTeCsxgoHrZYxw0ZnbgPps9BxHI7uv0yRsAgkPp9Lrw3
vXAoKySb9oZFjFpYDJS6xBTsLcW4iYn999ihRpS4HsozP3uFw8ZAa39rGgTLx/nl
OS96wz5DMs3dhoLX3ZgcOxrhQnygLzx84MRhH1mH2rARdV7Tgx6xN017k6JDgYKF
Mxbg4sTiSkODLdVlcDsTBetRaqRku35H7Py6daSCTPGTELdcPkCFaCNfNwVwh2zK
f7UtpgULXiFnR1N3s1sjnGI1AZWmWMaWiyepvtJAH5BX72iE0knNYBqq1LVz1YAD
+PBJ6RbEuVFs19lPmTa9BDiGGLztOGcjs2y1Ul/+8FYL1BWadSTUX80QWMpy1gn3
XEdiNVGpbPfIRi7/DIq3V0vRGntlj7hbJpy0HdNSpmY0WcemLnq/AuX8O6UtbSUQ
TPhNv5DX+I+qRbhVKo+tEYBPzJW8JsOJ+ns+HsI9h266EPLDLBLLEs7mPDS+UCI9
JxTP422i8k7ehN8IUyX+1J/56OIkq4B7QrkD2nhR5B8DvPzjic0FbQRBFBHA1HrM
Gd/rQuyA0r3k0Z72wNQ6BHVnBDhVWIQfyYsqqVaBdttsvE1wpDsnwUKWt1K/4zFC
FN3JB6J+1DIAO3qVD1B31pPCiJZjK6VGaOjydkKe/jWnZh4+5JygAAs95Dz9yDuO
JxXmck+YtUpRLbIeqgEpaOlLuOtV4aBp9+dCigsThEPkUvc9/L2oNMnaPAlt9gut
5yXsbbocEHPn+P0OKS3l17r/r0bYLTEIBbvWM+EeNc/01X7krFmojdnLCoMqGH2m
pfcCJLTB+3X4w131qPWeTiYgAs4nQs8CADgk3qZxsXMxdetk0/psta1GCfTpNVuU
kfnwVCP2PNKrIClI79kubqIoORiG+gUkP9NLFUPwQ7Ev91vE/jCfYFu47x+l8Whd
6pX691T64raqW54sGnRMWNbjSA2GmVatc/w0lC2b/XnS5IiVWfjhXMRTm+xL9CJF
xPKX+t+nOfly78clCAwBU0nMpLGsrc8S4J6LTffc7ssP8mOs883DlUUrtIhKcQdU
T/yexYNNjkqODl4xC7aJg/2SJZIob/U1zb/eCdpVjiwamnppyS9yiUI2M9XxMR/u
o4Yk+XByc/u52iI2tPe5ht5AaEdBKe5hzZNymFveD+XMqtbty2ye/pT0YTui0AfC
zvxrQMfXtrXyo224r8LkzyRJb383qjC0OQ39vzG0gbKQ487ZoTd4wTP4sXXnpc47
Po/KjAIBEwZpmBy+WnZLH5+GNJJ3DZM362HHI3QxDlouO9UoImYiXR289ZnaXrMz
C3xsui4PA8Mf741bznR5ZbwR33A8aQ25e8CbO9ygFIyyEnXBkgn0uY+zgZTrpgFM
tHJnl2kEeAP0S9cXMuMLzUeIXtvcHivV+27ZoVmNZRcJb+v+nd0UKhqaChsUATwI
I4OGeyx4a1QEDTi6YYSdR6CgWEtJ6dJVNgKnvQScQY3o1Vxb0x8Z29eDkKHcQ1Wr
ceMMePWpOaRT+AzKgYlgRIXmw/vyxQCeI9TwXBxA7xJnuLPQdAdFYDEr6ALKD1NW
V55f1ONAy6+4X3sj8GRTaLhRgcs6JYeiG+/leOKbPmeiT6NUWKlt5V1MNZp4VB99
uhO1tmATL8N9Eeg/nqmW/0UyfTFJ9G8RBvJ0nuG/r+JTungMnCbKx/3QsJD23dFX
Qx9qDJSbKVUSq97hSjf9VIbG54Ksmg1+khSrhdhmrbYEwhdsmWkAL4yn/lVbXOFP
X9C5b6XciX8/CUA4jkHY4IQLxuRnNy0tbFcBbkuQmKT/9sXN4HhG70wmdo42/NJL
KuVOHY96jGUs5tAvx9EVl2ERr0vtxpDm64XCCuJews0qxwyvflLD+FKi10z42M3Y
xwiDalasT1soOnz8xqBf2rEuoikTnGMnoHnTSYLfy+Ji3jFBBrlS8NN7paG7y8JG
IsRHIU58CeNn7G4jyU5oLy9AbM3y5kTEzacTKXwt7uPH4Za+O8Z48J10F/msZ6OO
EAcpsWUf1i+nugnEaiC0z6bWTZ157CubJAvi1x+4/8bbSP4b6g6wWgElR0olDH2z
6VEodo0WW6tbCEMJQ3IYE2s3ueg5JVJIdiS3M8Y1zttynw32u96EhpFpHjsScqt+
h1dxO+1yiDdza0rPZ4+XYm2PipALrUxTFjQ00+E37/KaPZMlKV145Vgwq4sTmPkY
cSnxUj2cwoRfT/L8CFq6fcvShS1XlonaiVJKSpdn/VjXeOxk7c3L1ISOTUWxhd29
ljvvsg0DtOcirzBK9vVKH96NtauYcFMtOyu6PEW3YhtZPDyPUMCoz++8rGkwO9mb
DE06byLMZla53KPFTrhwEohw9qN2nEKgjbzuy5CF5YtzyxnZX5GYjNiKqYkwcYuw
hPPICS6hb2wpOkbU7ty87gmis8j6dAGDD3QkDBknKVZq6QuwXQ+SkWnMl1adndyd
cscQL+YRRqalHW0G4DlpK9QIMUr2E8K2C+FBNtn/Id8h3FSWTSaFU1ssXORTVfjI
l+nA/4cp5i6bKN03lwpAkBJGi47J2YVkk29pJwBohGqk3JeXybZViWiFc1nhKM0R
lwRgAoZyzAkWzJ4FO8auBxI2XuaKnQ1vJQHmFclJwgZzbsQytML6/PCV1t/j4Hy/
82a1qKlagjKJEvTvzxNUtNbqDjVZSDSLJTNZF0X8eAx0J/z+VnLp1UFpa4QYkhhb
y7PD1VHUT8UGslY6RlLtx0dhknAGsgo+INgPjezbC32iKYHTW2iDVAEVLCsQxcwM
xHYbso9BBozu77HBXxF1lj5GoOkpGNBqedEiJBzbIYthetGfCLOVwEWwy1UaqN4h
/HMk6P5j3CGhIBqlV3nJG2Al5kr694JbXH/Ts8jK8MSw000mO8nNihvQjAwsC7qG
17Ek9XzBlPW8KFEjMh+ATThwyJHNU7fSiXCvcdt2Z7n5DYuv3KO3AMEBh/MOc/dv
WWpgKRnQGGWFA+vbkUlVRhaJYHJyrg0YL1qImv/sIIPlE5O8JkmErEtxXJgVz9TQ
U7Xkrz7QG2nf8wVDsUNnO/LQ1/0mqT/q8YjV8ybP7jwgT+nSg8C1jfeXosN2TEXK
EFhdjp3ncOscnaWoOkbDHzzeWHh2t/rrAb57iXzfh0JOahErlUFkgaGB6DcXseXC
1xvDS3drWwkqpWfywFYSzkAYWpUQ1WrJ+JSAYQHYEFHmdKBe5ff1tno9UBldjGPQ
2ss5f9KVd3e8WFxHelF3JoomaY5GmMIxYA5Nac+ldEeP2KGaDxICL/+lsggbCFLl
bEsftk7I6g0+2rEoZa0vdWlL4CpJvqnGEjkJYdwqBtEiH/ka0Tq4V4LV+EAC3WJH
maODeueZPa4D6W3+URk805GxybvT1lbvrFKpEc01FlJAPO+aEG0iwYMDxawgFFWE
BH+EmcqKraRlPCmnFh8rL7HnYxH0e4BCtXtOep7UhirBNqhzEN4rakSqiXDopASk
tQJT/mQoEt6qcncBJGLado5uuQSTAxoqRsP4bo7cUAAJgAfYgs8CeAYCvsM3dB4D
h2CUAcwVnTY3G8wHR+ZHhC0nMbvsMf2TIO7/WO79YK4rDoFkL4oQ/9haQGhQJ4f8
ENs3glJealhdYCPBFUYZvzPQ74yLlm68pfOu5mUwEZ6D7Wks51BHzWK6Se0EGvaE
HU/b9qaISBPMHzK2D64iHw+q88NPGhmPjVzkfNicBaZZOF0cJ/0SzizHPz/osPOn
4ae8f8eJxo7NBNuXdRXf7EdB21Or8BI7N1EyiJBBKMtYt1Mu6GfB0YDWvazD2CAh
xe1l+1zyXW/cGfBb9RbnxvarTi9pYCV50EfmN9PrSWdxMMxB9l4i8RZwf9/JJ2BR
jOFvz1Mv28xjom11ewfD18DpKMHAtUK1vvEE0uE7C0PbKwQ0eVorPPlWbGnE7tIc
/z9uK4FP3+o3YrCOAynDL2zQhErYRC1pVbOyqRLe3L4oIRZEvVQQzN1oGd/zOJAs
1URq9NaMC1X9wNFOmyywMCVR1PkprIV3vvfjbr9mTJgM9Zrxpuz8YgYY/ssIRp9+
RT3bFbxiWPsPJKjgf2BkeNxYIvuCvuaMN8R6y/lb9rNawaQ+DXwuk1TcS09pAuYc
bboepJUpylmfF1B+CGl6LUtdUR+uMkoM7f7ujQ5pTdy5e1NvEcGLNKyBq80C2rpq
0IAy2KQTRySwtCMMRoq99kRmNNRh5TlPIYjQywiMW49QWkbTmAXP/XS4JuT88G+z
dlcpChth8hEaJ7s/7El/eWcAQm6bwstUXVR0fccteKq3BvB8rYfNEaKXkC1zCX0E
IrN5hsxV7/loQhQB8hbfQ2rXnB8XRmhtycr791Fj+ttjQngN09oGKlDTTd+WWPRd
IajwkOblmwMpC0ls6MaI63Ckfu8mDvhrENlnFIPRxj923M0dK1nibq6RghxoK1fe
y6Ngh/TFFv9xyC7k8E8NW4YNjIeN0RyqoYh8DRLfvCt42l8jRPccE5JT9kRiIDNI
jbjoS0LTYWNhPb4goR7jGbp5szxpDHvqCGtqKrJDjFFqlyVhQFhz2/mwSSKcnYVd
tZ1oZuq6cxUfXplI60Te09lrliV+CMgUgkBQtcsE5x9AjITAjtgcMyB4tEF1+4EG
ODiQ6Rij4hCfg905UDk9RIVLAwL1XvR3D2oiVW50ySiQ9+bYAD2dp9BUI0mK9HEB
7Esm/pkv1EJ/Or5igiyT+gGt84Ony+3VTKr5a/WRRe+PB27nP2PamnN9uD/VNUDU
HGUVkW2ESDWuXlkdNYRYt0E4Zliqz/i1SD1Ur3177MsLU/w/8f0EZ3Imzi2eZWn5
n+oF1w+gjCGOBhPmmPHcO1fcaHRFj8KVNuWyDS+d4W28E7/l7wTP6rNbzjSILi3f
TtFBfBnGuLsDy7scHr4isYcCIBW74RCDRlDgHB/RnVjxyovUW27IivoIgsSeP2TK
poChm83+Q4bZXfx4R66OpN5aluWIp5PFrM/BDMJbRlF2sSONpMtxYtL8S4LTLRfS
vvGPsqYmZwr4KRdA7Mgp8Pv/lg4iUcIZncajrAmRPSQKXt0PKsszwL3dzBa2mfg8
Jlg8bEiHt1kG5uvF8mBaQlOivuDsFym9QrihGSpnQW8HGR6yIWSfUlSperJlSvNA
F5jZv9vrxawvTAeUpEYy9orDelUypN7+GtXj/DFfcRUFQi7oIeQaMn4L1/JStZiB
awcRuZsZZBFFOFvcd0pFBB+NpW1oSZJEas7fMeGCk5DVEFjA7WwoOHUpBV/8JXlK
/Kc3BbXn6rOQ8y8YttCbaI6oEvvBhua0rPsA269+bj4Lv9MV4kxNCiFjNyAaRtTm
x8vjPcXsNkLDaaAMGZkLMX6TCszQmFHJ8wCFuwFoEulSujh/Dl2z98uK6snWkIMC
lNC21w+MjDLfkiBlQhO+e1B1+7R0eNdOnpSxmMraFHhxGKLHhPP6fkSmBXKhrxQA
PC3SHo68YNonz+cTcZo7Maaw6P5/AncXaEPC0HxJpRU/J6TyPwKUENAr2MjyaD2/
RSwqGVpvcweZxtm8ogEXpb9B4Zk0kBYSWlXkhUe36YxSMOpyCR+Wde2/N0rD0Q6l
4gCprLA5d47s+PdMGQEHVHTt/u6znrRLDMHokMBTv8oPVuNJM3X7lrhg8DJ5IPph
uZ138mPK8WiXGvRQ31vkVXJeIj0urrRD0zpYE9EFVhCQq5teSTeD8YDMWU0AwRQO
xWNJo4F/dfhr8muT9pFIQUKzTbZMbF10K0/U/O4JYWL70Ocy7SimDNpR2TdfkabX
iCcrwfaL7i8p8wkchBS+ifRQRHYz4qqbeuKBSm+8rUHddO2owJgfgVLfII185UQZ
F1nX5TAdvwi/ILVSaOhSTVCmFyY4ukaB7HPQDTxUDXqg17uujCIkcgwoMJ3f9ijM
K6zGG083ve30XZob2cOGvOMsPHGPOoZqu6C6c5PZYCbOVZdPuUh46qLp9fJnRWOu
hq2wcu4ijUCnXHpR0rjyQz9ont6Llle+rPFIXDmwUZ0LVyzqMV+JEOpJDUGQpYCg
Nakijd4sP3EcL9+2vnjTu6BigJmgCwC1WHrGd6PPV9zs7/XQQrQq7Mn8ghwVHx+4
6TMzdabK9BI7ofn4rNOoYzQsTXUUoktFLNivo+hECXzrCS4cHDGHWDn+sjhXaHSb
m4rzT6ARReRsS8PI4pyu1wPMOALswxTksm94b5ZXPBlSGjR+QMNFhqcdnvYYnKiK
qYhV8C4kTwP3tBUwKU/ONecJvrAx5Zk/pcylQJHZdAt+p3oRoDhH7jda6ATbJW6S
rFEdmnZu9s1neA7HobUWdTLGhTfThC5sXYQB6CZ6b5EzCvwjQ+N39dOjo00nbm3H
+FmZPhqpEUa84hjs1k7BIOpjzq/rvskrnaeUuXin7DvrGzJ6UtsASC2Z94j/5T3F
4knYKDJ3gttuYNPPtu1JTKxZvGo/B93DwoKAEiSN4VnWpAmS6kfpNpPom6aHzmab
gOau0yy6dzArJ/cUhog31jvOL137qqzDgS5M+48hyZENUVbftpgxehYmFtWqRDQf
P0fz4vmAULavM4+fvtGgD3cV4+8onMJU/a7JGhLQju0aaEDY6skYiOrIrqewIiqZ
t8NHKTiDMmxPVZIC+HSj+g==
`protect END_PROTECTED
