`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3RP7BCfmLqPnttoEgAxuyK71aMlFC+1uqSfjU2eQYLbHhkp7Mn/Sga+gnAucdjI6
Ma6FSfx10BOwI9K6JGftbF69WTxkRSKSGiC9OQpVap3An2nKKRRP1QRY/BnUfztx
WFr8xwtUL7dJe3KkQWUradl9iM1WPdCNKYNbZcNK2s4meSIz98+pkeD55ELUN+QH
Fv2QgVmo8A6CSaA5mYW6o/g31wbE8blhJnBgyxKzZl7BzfZmPBt1pdDZWIyqntoj
P5UZtHKKov8BEDrTL/xTqGuiCVMeXevsS/DuH7c5qxJsiD9r9VPNHEsHaGDfD7pm
VLLlV0wfJhdUydncjDifHA5A1SsSn8FWbVVdgrXiAU8rag03UVVTyZZF6Nqns1oS
hVvNbpcJMTANaFECFyQax1sR74GqCz9R/waHE5Mf9CligqXrVi/aUXFKcN5tbhF2
ELMy98CsMfoCMm1NIfozWcjBov+gC53oo4cR/FceRr2QbpLzQfLvfg7YpGkvMV3H
QGeeebf2syZyzEW/aYHkj8Xk4Y3zOvdrotLPeB/mv3PihzsIWPg0LZePz9YC+xsA
qwOwZdHNlMLQM2C5m6JSJT/n5eIprqLSjW8yOwY5J3wM3nydSuAeaYbxGI/7iZTB
H1HDlnHIiljQt67Cw1T+QY9GX4rJWGvxRkplj1k+ZHY/7cHp7jQ+rdt7qnN99DGs
yJh276UPsmbdYfXUtpIqd/3C1Lh3FOF0alRq5goASmdUQ4SkzBpUUuROycxaVgN/
YNq6G6Iuc+r3kSO9OgOqr4iZRkOwXPncrQ79R55p1PkKLqm3p9ZavxkbKeawMGHh
OPoB7FxQoz8smlWr4xC9rCGf8CxQNvs7vDYEgbZRrwxKRBqQMUIcyN5OyZALOmIT
NruAbhoGMCPdqa7yJIWKN8ZuWs5srX+AnLZCk43XvILpQCt7kzQt+/2AeQmQHQC4
7r9TQRZ/8dGW/ZpfYywqSQ+Wb9w4SqY+Ul1urFmptAJ03Sp3/5IBxLFIFtNvnBlY
cQ73+oZmJaoUJsYu+QFyX7TvV4Bylhn+bRZn1SLKct3PVCzQAU/iwXfPZv/OKZ5H
U7Doi8YvEP3SQ8KaWcvr0FXSS5I9XuByjJl95TfMBoskLkuSmdaY2upQQCkpqWIi
/hxx1usqpNH7y8imCRViA7gmK76YwzVSqQ5OH2XkTovjuFzw9+7oBgDpC5qIIa2W
XpaVcFO3iLUt2WAYGEaL1YOa+5F56LBfoQX8jTQbl3FdJVoLS1eospRmJJeOWQo1
MkdxwwUvgg9UMjDAKyDZR5kXeaBEEIdcKK3Yxbp3IaR2Z7LqO5EKekHVcEJWjVaU
+XBulBA5lCDmeZiGFXPbTVfwVFMz+BifXMRgfinkoPPswkbMNmp6GKobjj3fPkyY
9v9Sn77L2bwTIAYeLNOPjTOcihA4H4GHKIZ9CkStyrhowQPpHSUjzfwdw0O+o481
YvnSTYtTkRQ0L86s/Pkg9KK21zimafadEKZz1v7pknelwqt3m8DL+7heyI/2juC8
hxpfOWEI8o8puyD+hGuSx1yw1MbRIdGm+zJlVEADLQFpJrj001uCiB87MOkz/bVw
jvKjpU+cHdqPLCKYgxTuLxlWl4/muistmZxVHVI6sWUaDhy1xzfhomtpETu/HnuT
lba8VjpZutxwwMKRlGSrFQm07ZciZgFSDFsDGqDWWYQqhb5Y81tA8tm0ostpK53e
EkUadOmJNJ4135gUNwo8+HELhZ77oPNYoVUvKxh0wu09r91YIA16v7RhzfwTiIW0
V8+ozTgmiS7POwvK11bB3e7jpZhKYMueMp3x3s3msA6rlxY0UkeHN6DEW4oq7xlV
KCz5UdZ+jPPg6YRQ7NtICnV/m5lx6eYxIx2nxrjVvfMy4EPgWYsN+0fdGlcAs6Y/
fEfDX9WBLl6vQ9tBLKnwiDfBGZODyCgEQg+Ww6M4stuzmO5YpU7EAiio20U4pgUl
O31Wk0vrKY+31FvDgaYlj9vtURV0j700bht1j9gnVEvfhe5MGmUpAOyEfBl0pcv3
xypU+DM4X49jMmjjsAwNXhiJnuIbLf/K/qG3Uhb9XpNAk/KsNB9gZV+DyLHSZWs6
fT1fWTnDzhLPRuktbdxvFaS1sx3f51qtx3rGNS9r4L9ivhqTON948TY86ZiPBIKv
aPoCmoGUE8rayjYAdi4+8M5+E+3+TXiwArrsGhtx2Rbz69R4MAnLcm4mcwV0gc23
KAip3yd8fnYRCY7eitY1G685u5tydDp23koWHeC6w/ISIhuKqSDPjX7pKtVJpvk+
3EnA8nXG8Qal997KIIMBlfUJ0V5d16mnuBzERvUeGZwxVuOBTmOzxOje3Catcqd0
xkHpsu4gEC6nSCEN6/jSSVRZTpu0aFS169FEvltZ0sDAHTs8xehcgqUV8WxLuueG
3kK0Rq1Hlj3zNegz5Gc5W9idFBgJ9BnpannUxry0Y47NBJdhR2j5P4DS1kQodmK3
YQEOi16A8EP715Py4JHv9Pz2r9ZcjriaVaVLC5TrsIHaAW8f1duNHKLVoUJaBQ9Y
VD+CQmKXKFzM2jX1XG51Q1t5e70ZC/KUuDYfSRTzHTXC/3MOwNIfHsL2bl9AjgtI
4n+1nxtyYvF4SifLSSjJqRExRF1VmHbT7z5Y3iI6KjU8ZBNzmVxdo24JgEkf0kIK
rfYeYMCo8l8H4kt769rc5poJtd4bZ6VYNHkNt4QkIynwW9H09a19j+kdcBu7l0rx
EmXiBTgz1aP7moOJPv3IzPI5WSORvgdG7CQHMWHsyRurwikYoQYZJ+bDsi0tsmRr
97916ByNQbGVM1wtZ8HVloSetPFYpnHk3wQ54XOkdKkTeWkLzCPsv5BIWwDpXiQ3
x6WeSHK6njMsC0Q8/xBxvnPeOcyz2CVCVZzV+wsl/qr4ZCXxvi5BHktY3yu35qwT
Y+N9Xp0+TFcIDnGAlwU0ggQA9XLzSasRPovzgagoudazxjgy/l0JNRN2b+G2ID4X
EtBIFPztA80mF6FFYG6NWUUfCacGuwUP91evC/L7yTmSxXckl4gP0BCxH8uGiH/i
SHw+BsDUUP2zzWXxoUA2uS6/iPbXG8UlMNob1JfoQ23rb0hG7QnsOrOWvN8URGnR
TcMa/zIQxswF+SNJxR7qN+4W2br4LYemXFaa/3NXTQIfDEBCTwd8ow0gbkWWiFJl
nppxPh9W//PUsexGPNCQmb141ejz8GaK8cayOR+Sb+w4YDmZ9PJOovUNrpffnKRp
KZP6nvViGvC8ND9ILPB3/XLAJVF2JRFi02ZEHNVesajSUNeVnmsJcH3g4UqkKPP/
RAZtk5LsXhbl76Ucz6RcnYU2iVEhdz0yq1sB4QXwub735tanA63EygrwZEWRw2UR
W2OmfJClR6i09sbPm35z5LV82YGJBOAoAKMDAQZqWdvoPicwm/0JShAp+LCtO49J
MPCVej9JvrDZ7WlmCLBp7eWz1+i1ZjCmFqjJnL8Vy+ZhSAHJpeSwZvge4dkUvVMG
+xS/Pg+y+zR3iGDSijVtxMVVLTXrHOfm4bCylpfAfS5HpxiX7o1BOykWwDtHlRgQ
mTnxj3TZb/EP8QR0aGCB8mKxC4x2b6RjJwuHez8qFzmUn8fI0JZon9e4sGJKlw2e
sj9mvX0wXh+bjGGrECyJ0KRwz+8vziKHysoM++s0MFeFlFKU/oIIOb67yLIJZ/f0
CnkgdlXJNUuBSQqe0yW1e+WTmRSKW/Arw5fjpYGDr5rrFzmfLwGMmlqp0pWxmPsp
9ZGjhC8IWKkCIt9NKjw3tDjT/qKvT69hrpQRoyrwmNtMMZAfIIRchkCpfTPaiYsD
`protect END_PROTECTED
