`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qhm+/B5ORjn+CAyE7ZMAHZOnKrNDM+BjD56UM2BXTikb/c3FVZFmRAWSVwDbhB5s
Thr1KbFUSiu4Q8tOoEEy0Vc1jRCe2OJ/ziZc6xTk9pwtzpCJUnB5VCNNW3ROH5XH
ue8J2iqznL3hdOQINCVKlIKL1JdwGCdlmQeeFldYEyXTmFDuxEpmgE4UrOSS+mit
aX3+oNIMXo97EwyW7vQ+Cp/kQwPt8cSika0U5kMVMaV/Lk7wxDGKBObiASeJvySH
MG51bBdLISqyhR+mhYk9McWfdqje71K6Ho0nnOxW/Mu/leK5on8tHenP4dot7o/z
zzA8q9lMn1uUEU4xbIQjSN9Xhu3w120CY3ybBmLj/PfpST92msO8WNIEfXKOWr9h
LV+7zJ2SJtq+PE+EglBkrILfPfsJVSjko5YshsEq5WmkQEm44hR2iW/oDsmRpkKu
1mj+5Gxgs0EqSDPLnFLQAoJvXVDKOKiZTmGzthvUSSbJjeh/PXxnUtsuRDXN4Ww1
IaQ2qVgxWGLCb0QiQfpmx6sK6YYPep7CK5jqDCO94kP4rfdxKw5PgcP/Qk4qv7Ds
vRKkHxbXOZON9j43js3NZdGbr4QxX9n5S+NoMEs4HLo5JwdfiEJRKrFze0zTMoWB
YMO198coYLHgB5GDWOQ6z2LcepEglCNcRvts916uqVd/xdg2QrX9FLFQRj6LotX/
OXKjeNnQdQ2Egt0Z2fykUC4zkSnq1JP10aGjitC+yX+VPj/03+tO4tKrxqgX6gLM
KSZSfYYUeMKkahK7RxsU43/4iMfSGm1rAzM+iiOXOwBK0jmFsEiiNKOJMrcMqHWX
ST5f5ZtntnA3Gui3KuLOtX+PFOMfylFcn07QZtOGSzVUgyrnJtWDiH512TbqgZNN
HPe9nrUb/EQx9iY4GFKCqGpqYjUs0KvKtBWbD01DS/qdJh/+gBgJ9f/5V7VLrCjc
tK0SSh1VjkyKBpWLdgjEV16dW/B4GriaGifKo5NHi2vfngqq5WrndJpWLViAYYfx
MZA1TCuWahJlPEh5v6ZkLL+TOK65RTKZR1msql9qDNCN5tFaPbIUJpbg4oT/Ukoh
tglJ8dqmm6zZbmSm3CRLI++Mj+WoQz1Bh12CVTwA0qXts4ulH7PDJg/Nkf8VuWLu
TlOeNiv9yn+KZanzmZ34xM2zD6bBphQmWi01EHd46wwlvrb6oDW+tbo9m+JZbGWk
kf4qB+9A9UbuDGJS/IPomq0I26H/qpJHoVJKxrVxw9Bgt6rog78K6GabGZne0Ptc
VeyWs8HN84SzpqlpD/8csA7GkFTZzsYy0HilHxGfew922x+T1C4KV4mabxOmV2M1
RxFRT111Od3L+qjB8Ti+LFx5iAWJ5OKGEqS6PM3zKU/B/It8Rrk5kqgGay3EEh40
+JefiMFevFDtNsSxPxXp06fECRrc0imRihsNCg98xkomy8baAWaA9c9H3NgnNBjW
MMkJgRr8Rd+A9harM7iXFm5o1BSwQaZjtTCnHrmcHX/Wpo+++uLLppTWTXmHqegq
LX/zmnn/PQPQxZu9RSzjjCzamut2J0m+o55Tqwz1/wsmZCbqYT3Eo931w0IJGGSQ
JLh0c3T51iY0I0hL6+QVWx/4jhy6bWLouP7++2wPvtjMyOw5kYXHKTlszvHoh8Zy
2rj1yES5Uj7B8L3RuR6XiktnrfMXD5N+U5ao396e7M7p/wxsDcvbEAZB+sTzd0uK
pSb2q3WmnmvyINTOfB1cUL4iQP251xPbY00efO8tf3nrXLCa7LruUp/NpoJcZ6t8
2hlcQ8L/OT6pJCsaYvI9lMiR9u+ijWFg26AduI1l6yXbIg8E5/VRbU1BZoT/q7zJ
VhzQLscaPp8+/yCyiZkRGNDMmJamXNcgbnKYRQGam4ei8PSIQVAUvWELup781A7s
LD+xqEfv/8lQwNnniQ3dYsdVgMiKJpPd490qtlcyg+LQ2ubehhHGeWdRiZU0BQoq
PeWFHgyfiy5JzuTFHqMXiAUvWab9B1bOIvWEuDVxsOWU9vPg7m7i/kpi6hqa+3Nb
7YJBCjKRjhIMoWYtuP+5GaLy6WFWA5q78tu4cOZJM63p8kyzYGpI21CkjmqA7B0P
jKMuHdmf3z62rmR+y6Lf3QbfAJVueZBrujfYv1Ezbjy/4CPRo5k8fKe2YE4RJ9LY
`protect END_PROTECTED
