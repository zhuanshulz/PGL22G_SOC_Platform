`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qqnuSNNiNGx0K5yNo80NtQtj8MgkLcjLYBp/TMYX+0kZzAHkVIhvojGvxz3DxfFm
ll8hbT57pVuTem/p3U3ZpmpZqUabVMLGjtzxQGAV1Cb9XAIz0T0u3h+pyyq5/SfW
/8GVkiJTurGKR0r13nyKMXpDvAggvb24+GjuWUM0lw5ID+QorLk6/eED3toq31xR
WRII9crw1SXU1LjkE0xqo9mHv7egMaIMysejVq9KIrfCFjKv4Q99vYSgXNU9XrId
wbV0VjetdK/0Zc1XAsSWaNwNXNFYckP5LzIl423VrmCjJmrdgosuAaq1q6Jz37qM
QynqWXu0oDXwLPatoDfsNGq3TnCTFmsDCYTvEBNZFqGEym7uJ5GldX41anhqzb62
xzIgn92tUhq8I58ULBDKd4tpV3X7rKohpG8z6V4dyB4+8HxxDZYf29Cl2A0PKJYu
As2JyyjKGNkMyeBY6rm5HX9603kKcEUDCWYlO+LQuSowy0ZJ3Wgg/gUju8nbog38
ZqbNRHd3AZmvzjkAdV8Mkw1Prn3+1DQjrdW4RC8yzUcaxtZTu3YIGdDTrfqTvwoK
pgwrpGziJdvF4jAzRHSQ3l8vwP6bYsRdYLeNdzH97wDM6pt5xB3XppiNTWXI0xZ2
dn5qB2t8Aho6mMIGXDiprW7F0q5Ed7gcmGsprn+lYoMqj/Dcfakzr5k8gJYvFg6O
OmkYuWbQ5lA/vbneeSiIDXlH4PwltpDhWKBH5jORDeQc3jh0sYwFM+ZebMcY67Xb
13Vjdjk/zwkYGnu5wo1mrG+7zqPDSJrUzt43Q2ze5Ot76e748ZRNSwCuBWhbzCxZ
Q8k1wZ7MAExEarJCAuC02Ft70l/3YMX81ZU8iCilGgVPmzqcV37PLpSFColXzUUz
bfdpNtuyTUHBD1H02M3xoI/C7BbqgEzwc6wkMNw8QDkHSoJsYggZDKRMcPOjNvyy
6xjnGqEhagEwSjVMG/Aa9Q2ebTRvJT2gaAPA7I+mViqw4Dz0vUgttDU5y5USEl8f
FmFGDRLxyjhiEzWrYu2DU0tOEOuXEN3mhkelLqXkPRXW4Zy5rsRgWLorua/+OI/l
4SaWJ7Bg+7pogPx/yWnQ0mnV0yL1Ck6mkdKg6z0BdA8fRTy/eOnKPl0zTCtGlUEZ
0aivzAK+JLPpwu5qDg9hkh7yjfYQ8twc/RzrKR2nkQOh3pfDosN2drf8odE8icti
Dneg3Q+I6CZrebs58mCIx2XDg6W1beoNPE5OyBYcD0I=
`protect END_PROTECTED
