`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3mFfFm6BwhSrX0F6Z2+19LPkeKMYNcLIbv5stV4bo4mMbz3o6MrdIcecsVBtuSiZ
cocj6Hlzz2BKJ8BT7VbNubfitkhDK3txFrlxPZ133lo0I4e+Mc5m6Tv9Tw/FHCP8
8ZRt2QWksdLOYNqauticna0KvKYNw17IQcBbyPO8qIN74zEklWgHCZj18/Ndhc5E
DXxkQvncQmKyC2UlY5mNd7s3UzYKluSxeJDNQmj8wDkhEttzAuwOIGdvPw+iSESh
qXa8WZMAcxdfuBenAbgMBhAUFaR32+3YjVJkXavJv3YHU84bcmpHL6hsLD4+s+KW
seC6Cjq8pS1FsgPD4e9aT+mtyg4rsYhWfdSiQVmZR5hygIsbOfwdfHgadZu7zgmb
DSqUcbiDXCZ0gSo0K1F1piBx6jpy2bd8neP5peYjH25uipCWYcrFnZAeiMblollu
du5O70oujcOQX3aOjCCU1EtmCv07/DVpPoAbQMxhr2KiKn+h/m03XK5NNuYd30Es
ZIwRBwRB5l0IWs70LNl1OL+WrsPXNJlkam0RTzJ7DIxV0OnAqMeYsdQ9V+6p4bXt
0fPWcl1aUT6wFcfKZ5qovO0doPyrmjK5dfz6lBrktA+GoSn1xAbdncWgG2kMIlRW
c8GVo/Ksn+hlfMVuP3QWQBk4WB4DGHoQlqdFDLgfw4C8QAl2oyY39RDqlPuTzee+
Vy7QGssit9YB8CmpIiDGiO4VbgBgGsDus5wEO2ag7ljBPKVyCaFPbUofXQ+ukmJH
d8tnxFfSs8yG2BXhg+gSRMEkTdrWaFQEyMnzEbBKk/GiNgNBJpaGbzttwJ/EZKho
CiT5G+x2OYQGAQQCP0z/RqYeCfnK3diKfMvD4ePCrihI+jAhbk09tkXdlksiOPvq
`protect END_PROTECTED
