`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3RxW4irTaXGMU0y7x/Ni35elsg3Dw3FYvV27Vw+Z2p+7/RnleNomEbN75crNRg+4
EFwf75cIcR/KK0qyBBcuWFNdm8NiuPuFzZP3JJgveN5BQhzrXj1M1gFmbhopv82s
gNtNSBaSTKcIy7Cy+Y9KwjaboTbAAQzNjoyHBcP0VFYn753zkwgEsaCe17GXmcCA
T1lzKJ3/u9qvq3behWZ715QpjmmG/3TXpHroGzlT/7XM+JRYJBC0XCtK0TEs52a8
zzyNikUS0Cn0JhrQdSH+mBIfrcv7SkFJ1FJ3TWuLa/vUpRK1f/CRtq7K/AtIiwA4
dCzCcuYJ1CDeCuKeX7tPWVVbYKqtcISgiJXyofN1yp3GJUly4VlwqhR0GE6Epy07
G1J5Ocxoes7rTOknN1L+LWXxlGoeWbhfpbXJ8EQN8jCSV/TvKD+4DxqQAqrzM00p
5RwTLKa7cYXibMr0l0l4tu24UIC5Sgl276URy5Oh/UaxPBw2QDK9E1P9UJGetfWE
6AcQEX8PxRcjgOlvqsJOjQ==
`protect END_PROTECTED
