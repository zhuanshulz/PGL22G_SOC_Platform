`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6d20C+5BgJ6F0OQFGN+aTS5W0E7MpJwwjsw/EntjP4LPo67dwsHEAWmjx51Piwht
FYk7CUsx+/bGCzDh1v6bj/FI1KgwKAxW56jgg5M3Ho9kIQRwa6gDMauZx+tGN78A
ehG5RHSdFHEMxtHI7yfKuLxulhqudKjvlvs6mOEOvuFYz7erccYG0R5SpCP9HusW
4j+hHIDveTlwx7V+iilFO/qiG1s31WQ7nM5jblL9V4oO9UK3IB1Go3h9xecMIh8I
fuZFmfyFY/6+AK45FzhwzUoMCeEeHpwnjZRO8FKdFOHYWiZXKZPFfJ7yujAHJR1u
hNgtw8uP4qeuD0olj+EMJSpEvqyEvWAEddCFSZbinGV0uQUmgj4OY4Syguvl9q0O
iv7Hx0wUIi/2Ga3uUwbHjNHkP193peHnD7hhrjg5cOGaYMhErmEzicrHot17xsyJ
GvAiYkB67SJEivbm6qX9UWbu/KlRHD9hqdWFTjJZFwJAOJwVvHdkd4k3B6W+nbGE
L8bdZTMbE9683ESx8LnNmA==
`protect END_PROTECTED
