`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QdCLE6M4q27WkJnJWi8E99O8J0mtZX5FYKfJ6yaIvkDh2I4EZOtdI567fyhJvZFP
5uGnUwKN//YdUX8KJeARI3/saQsomlzp/x2FATn2Edhyt5cfB1uNPDezl9IrA8a2
6QNyaUcl2011+WlGpLg4q71lpT4hjMSeujVyRCguB/qG2/AiGwfZVyYtVfEvpi7j
Xuy5/doHsrlxr5IzQ36R3fYDp/1zneXwHmk854mhw0yhF2WtRX8O55sbRRo3APg8
svVNTKaitejBCyVRe9FEdu66SVYBmpL2W32eMgXhuY2kZYtFTcsg/u6fo8ikPSow
sJWtb6uDS3JLp+htLjuFcc7Q29LAgQEbK1JmCNCq/YhSwA30kFRNBAftjl5wIzTB
QV1bS1lLTEtF0UfPK0Rtip4AP/cy15iAWsJbo28dqhbyrOer4v71nUA+VAUghjyr
lnjSxjWkuTy3Na3P6Ashlw45L/gqvSX9sOh9fkxfaHfpLnk92mrvk5BPVDqeo7Sg
OH9VkZQnb9i7aFo0Q6py4UeTtmh5MTe64zyl4Pocr89JVuTMDKussgzSq2hoFxcw
OTn552fUhWdhuP4WKA0e5fN9zKGDRn+plQhTkK4HBY5fvNjliu6lFcVb7qVsdcnh
kkRYvlYWlauVTLME29VSUCaofu0SM+Fn3ySh4bg25sjiJVzDTIeLQ4DBFlixFTmm
u+0IZk9ghji7ry6bbG2mjqcKVYzkIGLCkc8+OQqgQCM81J8fUWVLP25k35R0i5/T
EPckyOloZ7rNHcF3kpFcavb4UcP2E6NFXsYDk//BavVrvbixWbXqxicYPr1De4Xs
TGzy52dO67545pxG/EjdylSTe6vU6R7wC1QV0PyMNnLoUk+du3FriQ36feirIB0G
`protect END_PROTECTED
