`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7TYgpjzyLOYhm1QKjS6jteF91ZDemkaXA9cAxC5SeKAmz0xMzgapY7YxwoNdb73y
7j7HNGI6KdahzYAq2wKjR4bxNGX71Idj71QKSoQpOHPGCRgTA0tXRbeg3IlKkTYn
LMAa57012mrRUnCv2EHY43VfXmMhKxI5UIyfkylF7P32AXLic17ydi+wziu+iPpG
emQSniIfNUOItApj0hiCDHVpNgWY8Njjsuc6sbPp1ycEnBhZufm6Amc1Rl38XIC/
jDXCS2dwvGXPAv1AuVethEbOkOnLmL8Oh+zutn040sxPjfnxkWsApKtd6TPw0wUq
xUPB6g8Jo+ElOZgoEALwCpXpgHRgsg9KA/hc6I6hPdHDOcLYY6i0/AHiy8J54hOI
Slxuhjy2FRzFs7e1WA/ge4+CY/pWR2rIrfmVlqbDhj+qHpQcDcX1ipDld+NgITib
JiJNrVYar7HkVpWwcoxS46udqNI3dMcf+qgnwTSbv5RbIc2k8rUfXLIUBc3l5gtW
SUfMv7bL6WtilDIfSqYUI9wWA74Kso8QyI83VEri+eCuJ2HW2Cxy9sAYj6yvc2WM
juJPZXuVsmAkluDopsWzQcWO3C+poViKtLxpuqargCA2JG4+QDZjio1XU9pEc5UQ
KjaYolxWT6TOUQEcGm3QPE9C82zv012b3Ddm2QAw45zXc8B9OJ7hRg9WPm/mE9Dv
N90yF2PYKkKxyQR0mS/OtSvshge0vHe7GUNv8yn0lc4eqIybc+B6mRl1R4AE2p0U
3AYiTRh0QEbJVmNKiA/jXuPRimakxZcXwXxJ4rRNIFI=
`protect END_PROTECTED
