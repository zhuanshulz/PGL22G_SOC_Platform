`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pDpjWFJNCaeA02+FrTB7n0DnHI2aAHgAsB1ScDHbCACSW1moNc1C/AZC5xYBiRM3
dxLtWrv5icQez/tiheMgpTJeOxgpzqFXuau2uIqOs188k+U8xglxQmCSo/KZnEPm
730kbDElGSvfanNyaV2QhwpbfTUtzNMvH4FaQpngP3mlJ9193iBky62G4OlHKKGj
IXKBZDvfCFiI39kKFYkMGFAhVWX9MRCInHo5Qp/2E9pDgvKNPWzE44rq6IkpAMn1
MAFY6rs4F1RBTwUtL20kBDz68aFxGBA3DAQF0FjtgcJfKw27Ow17T8lVGyDKA6zI
cXJasMNPctP5py2ITo3QtdJ6DrHR3F6j7yqNaOGEiJFZkn9PdgCGPu5yTrIJo/5M
/c3EkI7l3AXeYuzJfBa7HIKwaC9NI+4/7iuUrNK36oGjHhNqjcwA31BGVbGcTTON
IoazHzb0OiMqi0rewRcQu0wPFc2C7dC+3ewnnCmIFahRXcWacKXXtkBVgSI89L+7
Qxfz9OE7Y7RcU2PqCmD3Lf29STDsJub9VYSR3D0s10Q3g0EtyD8m8MEa7yUblZRH
s4ezexBUoHxWqCK1pqkl8ZTmBNx058nhJ4eJRcU+KhB0ABjhwp3LJkHIwvbvbkd0
m4/2bVdnxFPA4DMNP2Vr7ZAQCmsnmfEzMK8uom/Nrc0hsVPEqCg37+6j95nb0IYH
uu9bjNvUuT95oxJ1o8lxPbMwy4+xTfQk8aI35XSyUNYAOq2Qx2DHGGjymUoVEqli
sfzRTN68lHiVZWK2BovIpuF+UWRiVFuW6Q0vwNkoy6/gn/vImiRFc5duQj76mYj+
VwnVWG/4+791mtOSt/DXElsZhH4dupskKXbmZUBDkY/ZlnAORBtNmkMDqUeR1HWo
cUeD2FB9hg1MmhQ0IHoR3spb23utgFacp38XCrns0A17tUUdmyZ0s9j+g6/OOFMm
o/XPUQeW9GelGAVq8kbjBnbZ14CwRH0xRlb6X6kaLq0LOSBWlV8kKBmD2fHJrAbn
FOzqm2gbTTEIQJAGO/z4NaApuMnFcdeaLZRs9/sxL970/6BNZ7wy9UnRJGFjvA99
0zjcysoWZU1wUMXAyUmMWFYOBIcRm6u3VNBQTfVUVu47Td1dRV+o4PcUgSgRMUag
kK5oEDlIRZnErr3adIdzC2YfdMoGn+M3Kj9yJnZLnp3eqlTGsBRzAdzIUuooJrXz
d9ntrmm03xospJ2kuMTxLECQkz0ZhoN3EAzC2Ef3yJ/sbyLfD4kVso8LLVvPECPG
hwk4mZwYFeDI8UNmNyuEGtCXTxWisCDMRVJ/7xL8sxe+v/vaqOAA09dfrxQFDk+6
9bZ2tGUNjpe30rF+JhgBv/dawY0D674Rx6Ic/dGrR2kdvrXN5Go00HSC5V94Tf3d
4d8VWRAlnwt8es37a10W88xaZjec34pciUL/O2KQoRjzY6cS+gJaaW1Qep7yxUsC
MeezGwisNksu/2Fq8J/GEQ==
`protect END_PROTECTED
