`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
98hgAcYfjeFRn4WJsBhBTCN8Jh5Z67tYLHMOLBMlmjkesbAARV+t7sorYRfmeK0P
udRoFoEB/o8He3eg3fc0n+5b/TqlMzErRHCs4bYsMoTj0GDgK/F0mJdNfemVeHTu
RPy4QGcomTb5c/+PINCrWPlcjaqqQo3Mnbj4fyMkpw0hYAlItWG9xddjVGgakSV7
nj2o1/hNDITIavQo4iwyCBuLEJJ12zPZ0YunS7Xk/WpKhH3akR6bBMckjtUVSns2
F0RpegV8Wq7c3fNlLjhrOpObuB2gUoAm0GHaYWdxwwWltUDYcPC6N1GSGUv5y5Q4
kLnKRe2SrfW8kHbRTRZc31Z7jx7BQA4CG6VdKm5hPehmxJF9KCjdgRZeRUHQuZpj
Kg04rZKM6eUyEdITEyZMGMh7XNAQKNoc8V8miB2bNNNWV1r+R0W2OqnosW/695EZ
GVbEmADy+2BUHAB2HNRuLbFedqLjxX9V/3roKp/E9tHehgxkGTB33RHV7O/7252A
23hFeajXZDaEo7kF4Z72/V1QsoLNzbk0ERkzlDMMpZqHnyN4hXfzyooAmm37VKiY
LnjuW45f77wPSm3mHH/99AYfpCG5OFE2hiBjdWJzqNG0hgM+jTiyaf+Y2em1dKGt
o7fPpkAm2fVXmz3CHMEbl7QukMaWQHmBX4xpiHwSNCVCUznq+hoK6iIhcbgOfUZe
2nPYPi2pKCbc9dxPMimcMrhixImwOwavHSVgcMi5u27Wx2I/N+LReVUxamxkv1AJ
IUOzlRwyvzrw4dIwQQGWdU4YYgyXWkH/aqMCbCARRYxui3qHLr1B6pwSI0iZjAO5
q3JTnLk4E7Ic/idz+o7nPzzeUG2Fbl4RFGSifyE40ett9Jh3zy/0KtHGD5Q8eSMK
itbqP1uzBaNSi0GbKns3OIpwxwUuFmDfGrodR34W9GNjBWJTB3sxU4rWycYaYg2c
K8zfzKmJBYywtZiikOL3RYJUr+GYAoK/67JpJz3Nu0QRzdZwdqC9XUxhkck2Tqgr
+hsPGjcroZkwxqpXBrIzDA==
`protect END_PROTECTED
