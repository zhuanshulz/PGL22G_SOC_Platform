`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IPfyJREf389C8Hxl17ZiGLO2tg8zR8q7o8LIjk86g2/riPxoi8WPlNfa3oa+zkUz
JEENCIT8pcZuXWGbBbfgEP65Imge1jmX0TLQhLUk77M8gxeEuaPlRu/HR3cMjWur
pVlczghyD5d/AZgcxuFzkFm4il+sKdnfQBCpfeteHOQuez5R3Omdk+W6SwbHJYzi
XQ2JiS/Qp/egVJc6BtQtPGh24DvV661XXw6IxHk+DgIcv1eZM3K88okGgx9+ZJ83
j+F9QtMX7Ffj9kGIulYIIHchjInJnUvA4OY9npdeVaEWwvEAA71VNcZrgNFS99th
jfapxlCqi8BimA/DOKjI8BNYtl6AZWBGSRBlUZWonf+L1bkLt1OGRRScihS20UML
PHZCvNIoygcRtVAJObA1e41qDdXk5XXexl9Xlgo4X/7NmfDgAuLda1Iu58uQW9/O
1X3CJOpcmkf2dKMcXUwtcGkriEQTQALRec1zCUeUxtl2thjSbKRdO2Rlj7opcKFY
TH6HcCpWAu3PAgJbH817AV5RNkbyA3Qp5vKtZIL1XSYcSKXwCivbmd2j7GehW/rV
5WmqyXNWcUaKA7GHtN/nDW6Z7eAKlikIiVDzfguEfckyHeBOH8UugUyZDSGzdaoC
j73cWnM06hEF93wLltgbT5kUagwxd8VATpEHhCIzUBddNYaYvmYJ06Q3f++1bCpz
gK64HEh6TX8VZjWm/6IW3H5YcaM+7/hcDWVZDjP4e3EXhsHDGILGc2svMhrNWsrl
C7ebs4i2YphJVKN8fmYDthAsbfTq8Kit/wxt232tVR5/yLPHdsEOWAGpuxpZ/mVF
er8L3nJ4iLL6F6r5AgfGltJsGC5QDH+NIW+VjO0r90tzSH0YY19GXvur9ucJggxC
ToIdQ/4Hyv1Fo2XF/XFh78/Yr+1vqF1scCmscr6W1nlHXkdPEAo2vzzfd0EJXaD6
3g2l4M5fPLFLIpuFsn5GcjUmCGRObMYApptRPTMG+A7/Knlp+JOR+Fwo4VQ5vRLI
rsatn3xmq40JVR/xsAjp++RP/qnK6rmV6tBX0iB6ngS6hjpNWT920k4soBq8Im2A
L36ozbE+jKaHsrvDVM+8XCvxMMnIGOUpWd2OmDh+ltBpFB/m8m5XW2I2vY2q/TZq
O1X2mfN3sdTIGqykFhXVHWzailGgUtZZPquNYTpRTVz/w+fj4fQKkbArV2V4FRGE
UQLx6e1Ww2iVOBxAn4QoRqs75QcvbMBQzEFgOOs3RGGAqvDYvzxfxJqbeTowxYoR
lklK6q9NJPSl46+Z0d+fCVk3NWGwr9e7lEPTJDup6S4nNfexMFxPwfeOi5S9IZTT
xrjzUGPVHlFIbBHpcrjepT0LWCdX2LQ5wb5ygz5QdWfm3WS6FduuOJhVdWn4rMrD
XcH2rYJ/7xrQRZoOjXcudnq0f5QkGKt+BAaw0uBBMVIiaLSB/860hOtjYI1VfAH1
cKKp5fbpZ3dCuOgngre8Jvqdr4UIPooxCOE0b8nao7GGytKKQwJxI0mSGRtwvQE6
nQmM+gSC6M60YWMv5AcfF9TxFfosCrEHUub+JYqttLhJapyX8YYIHMPTTBJUgfLe
Ca2X6IVhH8AkuQ56mU6pJko6iS2W+oy0Ql/nE3mhKQsTFDL4jvxKVKXycbvsYTj8
CVYvWoJK5awTLgGweJgfPqFTEM7oM6ZwtGt1zGaiq/Sl280o0SRXJmNbdK7TwumQ
mpM4DVTLBKW3/rwvvtT1a0O8YjnyPqmug6D4fQjMAmW3Xr2kPaBu8197zNEPpRwl
9wTQhYzaAcR6fOQZa04wAcAqoH56kSYVQpKcVsC5ImrT+TmMiDij3yA9x16fsLFC
z0P1rV5Fsmjlznh++EVrJ8rFAh7AJO9z0MR77TL77kmfpvHf/JNWjM/SlwLu0IJS
lpjj7ko8/zIiDQ3cE8trNjX1VmunB9+sjkRpZwkj8CDOaKjWn3tNU0SYK07md0bA
tcLazsy4aC38GZfDebCmulgGT8SoeG0CxaxoFsp2mNzBmJFCYLDbjbiZSTKyoOnk
3czIYvl0fB2nIT95+1dNJCGoHyLPhBTmSqVVAwZbc5cqvVGJodoYRbWXCszxznyg
+0IVgJsl3CvMMmdvyvNvAa4hbthkyZxW1FCrfRunlT5cYky0iC5PUbExri6Nh3vX
KOPi0q99wKQQ7xTCTATRQunSZFqbaGlxOtZj5saBukNl9LVqPieeyC/GnKxlP4BD
60ZwaJc2d4BH4jFhxEy2Vyb9icZaqhtV/1boimU3IXfzlqO5qYSMvoi8KkDUuUnN
p6b5boD86O72ORbzCmdDUY91ifXJvbyPLe65Mp5Sy/lz/tvVJ/Gn/uU32heuVKQP
osQJ0yL0l/Gq00T7OunArdaY0nu6DnNjDOnqJ/iqqi3/bKF6FtoaNa2UP7eUML7L
IXpNyMura1Ge+2ggHnfS1GBXOg16WyGAYnl4z1GuKDm/A/k4VyYtWkRxZ16CuID9
`protect END_PROTECTED
