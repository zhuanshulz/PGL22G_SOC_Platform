`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
15Stv9RcWCSLvDhsClSV/bK3DNee2WX6AVGnm0q4M0iZ7Ax1HQiKuZuVznnKsT3M
A+D5LnZGU6hFQS4UFiLYEAHmjx95VLjorUwz5EGrtmZS/jpxOdG7P47B3zaY2FdF
Jul2uDO6f2rC0VeKzZdr3PmdBKjUnOviX9mzSYzJajrDgWyb0OwEs4uV/aJMf9KP
Jh2qsXL1q1Bcg419omBmFU6U1z6F/yPkxpTQAh51cLfJIIl6xzQThwOEQSs90BIW
hUIkYV63SaJ5yixq3P/Zf6jPnXEbA1+7IygIEd9X9phzvu5KgsF1PXg9kSLOLxQg
fpm8boHVZs5WPlG/l+5xIPt75Z6pZ86XEKN/1hgT0hZ4zTPLSx3liPf3yF5/wiS0
bLkvUT3WQ+KydtAmijwGeC9DXiZSxLRelkXKXS0MGJ7eImdi85UdBS/47aTlrYIg
5PN3tXq8N+0LxB6oOCoJFkMFFxUcUxDXu3YAvs3aTJ41H7Qi62cfcBrM0+t9s/Uf
u9zXqvnbxoentA/HQJh/1SDMvVfqCxQ3dCyqeMTwlFI7ItdPfhg8RiweJmqm+Q6H
S96Ur9QAFJ4J23kY+huHEW5JlicLcG9qTyLsTs6Io08YViQsKPqEjjpeapz6XUHe
f7I2q+jbfODOH23CIJTsRA==
`protect END_PROTECTED
