`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f1yY8lNkPuE0Hle1iAYHV2DctKPGiCbexpCPsm5skl5n4dZamR0xxDmycIX1ZRXy
yV4UYX8ppNd1PpUbn4fTUqO7QmdOyfY4YyIbUAl29iT01tIGo8rUkKbCPfPrsybf
cMiQwrwOdFy4S7vpm0Sk6dTvkpPT2NNkYoWi23U1pUgzbhRUfvz9+bKkG4K9DlXk
4AwfbXwogTBWQaKFlo0JX+haJQbQSp/qv+Un/WUawdRna3ueCUleEfI1XOgkCB7s
LvIyBkoJ4rZYyEi7PUPVONjfl9PPPrWUCCixrnFF8/WKrKJZLmjHGfqy8rUM6IfB
N/8gbS0DH0kbT10Q7rh4F9dXLaMgXL54eI05k1UxOkscegbBWv9IQihSRAIjxs46
HQUjXcpajdeaqZnt0GSCvQ==
`protect END_PROTECTED
