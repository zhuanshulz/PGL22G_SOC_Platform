`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4LCKaaSD3ITE7btV72bqM3ouqnP9Pd65inYNxHBYuz62xYFj7oXzZ469hyzcSeVf
3CaCeu7JZQl8Yb+dDrwNvpLBuDyFGKepXG6BF5/7DBddo8z+TxcirfL0qeLAndxT
lXDqd05dxjF76DIg9jfl7QYPEIYC8qSCvwlZp9B1p8c4oLNmJu3BzwG/L2poYCp6
oelJiZhtbST5Hh/0qlQBP1z5M+6KRgipu+YGxpBjJQN6qmSAreXk3SaIMvmtr6ts
bBRwtDlvfjvDU0Co8pfKnRWgTa0ZCoKIVKajcx8yGRrV2aVteFy0AFLBmGBNBLFf
o9xlxYLZ760ByFJjDTWpHLWM+EHBFTkNHLuqXrxH7p6XTIJ6ck2m3uDUjxk0mk0o
i0N8kFceYHQ2PBzV1QeLXP5Pi2E/FOg+ePlj1PR7gGOuvJFaGt4pNm+alaROAmmR
CvNuwatissgUROkvLrAEutmWEu21Z+wBH3tNY90m7UxSClkNJvxo9nQSAv6Xz5C8
ClZWv5eOdTqDSFpf/eLTwIHrlYU8RCx8XHMK8x1YHfxN/AaaN0OE4otk0EOr5BMY
3S4CU6Qku0zFxP+7hYBEbZ9wbZOLOTJkuq2RWKpKzvqjpP1zgFi7h262Eimz2FH+
DKrUaD5G6720cDKkI89PmUMM7gM64QKino7o72bUoEZFsb2xZPtUBBKsQ1vkyClX
Qlj2wqSdLCN6j7L869L7mRJtnD5/OIv6yxxdzAaObkXnIXhiUY91wtb1bMaR/URX
`protect END_PROTECTED
