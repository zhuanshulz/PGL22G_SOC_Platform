`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1Hlr7BEDwUF6cxgkfCFvGucNWPDq90YqgkQELr/ZKk6Ym9Yif07lWl+YF2GtWSTu
Ohzx3jpGevxWxq7OTZUcBvBS7SVzXsSnNvOX1ERVFIFQhaXhFmjbV2bOfzoJ9uJO
2ecnb9lFKbdi3LbVXxOoKO1xNnSlL71kWJPYjYFqMp0b477bvhv6TCANRtp1jWTK
mTLlsMVHVTKie7gc0S+pPhcKc93FQzlhX479Ze0KftUk+ngUfccsyGV2VTBxXrX0
06mD70KS1YzpLvi8GHGeT6zjxeyGGMZZeUc+9MB3rn6FXA/a7hANIYAxjKD1vngk
sibMZ7mIFROkJmw45UkCxPMjc/c9/PuVXs+YI+rWcLXGOUZGX3IG4l086se2p+/b
JwAU1MYKm4Mz+QkPJgsdglqfQljCi05xVpHv29cJY9cEemT3quaILFogsDCpAIaI
f+D4zq3IhDA5OXVNT80QJxED1HIMcCptdoxN8qjEVVUpPUtbN+VO3yj8mrMUaU8R
zuca/GsWdNPt4/00oGFognKHADgPN4l6Ch+mfWT8Hc5PHG+eAFSiSDkvJcZC6z5R
lvnAOMkDD429EN0FYp0HF5L33WkeufEXEeT6uGiQICQaIt4v5vwy7BuNzn03Wdbp
UhA3U3EymjEoVw/Xh0G46IoOmKaxag0gndib2ls8+5jJrwliKd5c2/aTfjeWzT+f
3DJi9Ybt2O+s2h5GAIpFE4ABJdk5lhQ2cUlIX53As+HdcQPKvYyZkmbDgcGioO0z
pg9U+xMRY3lFnL4C/5wI/FNDqYl16cMnC0Hj4TVl0omzqVNYfgf1WNpfZ5ZYCcIv
6Bd28SYxiOu8c4qjjRVxNIcnHPKvCDw6fY5/n4ObdzwLIZ6aTpSz1ZKxGRhIThlo
JFvOOf3KRyCb6lBBMHj9ixIlTmzFQ2VHlaUPdwDArv2FQsqtdaCNCoY8Z/Xic2Cz
tKtn1ZQYIOs5MSQ0J8beWl4yNPYJFDZeIS5mHLBzdI8LbLjVZB9jg7HPisIrkjUn
8YZ+ee7rZxI6MviYgbbmSph/Isci2pI74LIW31GvpbTXc+5eX3IPhbr0bUyYwTIw
/H54mKHWFSuDPmBTVQHgUMZroWNS+weXgm1DtD1uBi2wofqWem4NeVMmFeIDt/95
xpdW9AUyyhMHw6xx+0VBSAY9IYIpnfQmlNCVsY1aeVDPXj5dZplF3AWeRrcJFsyY
I4jOvr4lZykYGQSGbtcOFXNVYaJt1qkgs5F6LNbHhQuBnqVTjeYA4BR7+DWJTvl8
I08F8PkKYLX0tZRfaZy9yxieQTSbw8EGMLgNlkm+A/UxH0HZOwTSSuLFRouGNvSf
AJB5aPluf3quiHlzXkvlYgWj8NKl/ndKipdQqe8Uz1NAH3uJbtJkQjB46pAcDTDr
atkDIZn1MjDWFZQzZBzlfxl4HZynylTcatCt5hMGlE/9wJhhH26BF5QNbp9DI6gv
S90eD8g6VMEfz/+Ec23Nwtnq8sKj83nc6nmWUq5e3JcTbHN6+o1RqhTxbLM57e6y
1zexnbgQMxB+dBgqt5rl18W8JI+S43NymDQB1OdyoWoaczPnKURaHWY4Z7iPzeT5
87DK4nPLqppPqcxMAtKwuwn5bhn7i9tsh5lLlspkuelyFGXbQIquxf8uuGmGCJcm
m5fUJ/bcQwYxKtNGPMq/N1hBusSRKVm1UgdD8FQQt1q1e9mdQB1EpFzMUjPO5drM
8qHf8e/mpEjG/evwIiTJUlkZeJwG0gSmJXEZBJrKJYGMYeKb4M9ZvAgA0+MgWc27
PIqU1NN3ckZfeW7dPtpSQVp3J/WctkmeLpE6hxTWrIQewbxNFxD+d6ZgD4hG129u
vzsLl46fnQho25anHt8NTjEHSZ80lIx+ilBW5SUuPVQ7nq7tQb1zmU6XMus4M2zM
NE/nBIdQNjDMqUdGmV/gCExWObueHdnTpb+pjZfIsReofnpq/9wOpinnlMoqgTdI
XjR0OMC7X9J/bD6joZkNThvtKld/3mqCu5JL+4W+sBPx5qEDaJfFYuu6VvGxW6vk
GEaK89Nc/Gg2qhoY22k8WH5flC2YYYWpYUitwwQEidSN2ZFMEoHmZTNhYUCvCL1y
HYpiPgNyWPPGrXoCS6ZlzYkQ/3Q4CfzL/zPT/Kmw/Jw8+OhogXpmCN/HCjZIphSg
ZOBVPf6IhP1X5DiGbo97OkZXUtntpegLr8vuwhqwW6eK+iShOuVOIvhQsEy4TsXE
2kF+zvgKsmEE/9Kp+/ZpnGWLnNiUQmNel0O+UR6/YJ4AuXnn5xfs/7t7aJPF9GlW
nJIKDWtiWXzsmolxaIeTO4niNXhyzgApM6z3I5/aZeCn/KmuIRIldfNuMb+1Kt2V
Yp7XiDbfsxVI1BhLAYqdojbbUKdN5Du08UpWTzNc/tVLa6ViWvgaBYjB28wTytRa
Pzzv6qxnFymdnoC8EjPg3bos+sYIx5524p0znjV9dYLg64FqSXbTUTrTaDXbDsLC
qMOUfvW+Zbnb17sYag+ctHRLCrVLvyGPy+c/BnqupUCIF9p1aZ3FtvGBtAFyTaXr
oJrXnjbrytaDY9MGqfP3enCccVW38MJvTTpCZuZq5/3PiwWAOA7M6hHQurHWutuy
LB/SFziJwAaBVt5FitcVbk+aYcFde2amNtmCfcMYkeKQYrOUZkU+bisg5H2XUkLy
rCpqTxjQbZk0+gIkWJsFLZnOrRymeXTBB74HYhjlZ+X0F7lpwOBUHrrsN2mGhGZd
lLyEZPrFRAGgrsGew8KuSi3T4R5jGGN+YkHwWUpZsk2cA0SiW/x6QkENkO1uuoE/
voAG5tUjipiNF4wdT+zyey6b/eGSf7SDbK9v5woBSAyvHTtWpGkqNrU1I+78PCx8
grI3WMWunjgHwteVPIv1jnD6FUUdn8QZLRO4AbVkacL0ik4bDG8PymQa/SobBLHl
I1wAwOdjoyS1WMDMXf2PXJbOKmzDw77teoUroCrF9R/WqzhUV/WB71nIbHOmQfEp
mH2wJcxiG2aWlRGtB/mTSw3ixtr/r98D9JnpxwjmLdP//1YSHjJn/iUAQZBEN0Oi
cstLTc1E3wQVToHiFal9FFDW9tBTDAaYBmXKnwkFpf/7mIqIYyJMVpufqapSbzij
xz8cBRE2bGKUj/IH402mrp+8icWC+JlzSF6jAEP6/1GLI05FcaBdC22xvoRbLLcH
XKjx/fEEEiAj6hv1yDL4PhjiOvJvv9xKPLrQSdcRqBMDjPLuLs9pm0Rpc7CEDHN4
bNn8c/6PwPM6jujLctQXndCcZxL/Z22Co/+aDZj0eTsb1u7y0Iwb+AsMpckDI+Vc
nqtVwI2ctuQRYeQ0q6bWrh2FgGYASqpT54xVfvawgkPbF4kzE8Q1Eadx1MouXcx1
/89ZmdfmrotGy22qfOQOjDt83bFZCx2vpO5T1jLtPRo4bCOiy7Kv9+XjH1t/SfYu
9MD0Ku6TmJzGilHqH5UoqpDB2Z1rLszY6jtx4l5I5AYvfaNMhoSRXdBTBSUBwO6J
9kKcCFuB5dN0gy/brln14rd/zga4ipWXqipQlhfS9NyClr/kGQcEnwKXWqsVUxmJ
jw8tYSoo8hvvZ8DAdHHGfEmJIXm58xtuRPY1dgOykzZ8mf648tLBIc32zgLxzCQC
AWEy2jkJVyyu+ulLe2kP2RCFifz1mdoXTF72mvFXd9ikiOpjUV1YWEYuvQSAyEeK
zuid8WvmgphVi2q0uUHxeKKCc6IgwLwaBxs8ohxbRiKmXoZfsOfhrEtDXSO8DXe5
t9U+OLnmTeFb6tYDwbCP42iIG2ixGtLqhA/LksvoCwhrIjN99/4BjvFFdzCyOrZz
PEaJp7V7I+w1m0sYJ3lDzOtvUAP6u+oFhF2v7OjNIGObKETPcJudCp5n8w3oWsZ6
vlCUX/I/nigL8tX6BYByPhCrXthq7FKntQWJ3tEldUQcEbsnAlQQT+pY3EGPeNJk
/DPp/5OlO4P1ItXBjB453AAFyavZgx87oYddEhzZQ0aiJgWbQjBQoBEVtXZZbDH4
0iTevggwJnrM1Y1ZpmdKGGTP8IKaJtWZ8wwcFzgDwdv0UJmdx0YqMrkzsm/D8hw1
CAS7s5HTZ0SPUzwH43xtY5Z4WFRbVhaDZWivye93ZbZz4t9oT4jRqxQmzEuEEdrH
GMJMjozAxo1vcBgRRtila9wSHg1eOSEEiKPzLrzb0wGuPq+sUzInzAvMpnYZRgg+
cxNe2w/y32wjsdDQyYXMQPPbfuL2aqff2rxNdxRhDXN7yEYj1Hu6gFRq4NFJK52c
neaeMK7mClKhRUqdTF5f80pAXEBbiTHrJiC9X1slSTDnSPnl+zYYbSUIr92jwkZN
p1zDWa8tTunln/2Q8jjm14tBgL1oEGD5b7aaIrbGYejTDqNYdLgyrTQOCHD+P0fw
OjLhUhkQx5G297ZpUGskh+7mz9uS4FVCMu+MjJl9I1O+8N3u8vXjmBDb3YJswlmw
vUUeYtLSgLEwihulYAwPHdo7diG/PW8mb7QDRxOv2od6LHaVzbYQb4/k84AD0uK7
v1xojUNMsgwdk1xI6TLU+KTvxY+9UDlj8k6T+lJahxPeYsq0aShqR+sKYE5hnPJL
/+qzdeapGByCjmk6c3Xd/zxlI/gBMenKWUWeXJ2/m59nQOyLUx1jpUANB0S047RG
NxShRkABb4tKE60sFJTndrkP2z6IvtXNfRi8smoSpIoRU58+Fs5IYz7aIIQrM3wF
8wNqlExg7STy35MV9kmZTEKIsBEBmT+MAnC1/utnR8SvHMHlybxFifHuatfVw67k
XcZ8/g39Rktu/Scguxqv+THfaZfByZv1o70LAoBbFiBW6FeltBhHyiueD9m0p2te
nVAUaENn13JiyKhM8W03ltROtHoJbO2lbR7nrRb2bQVqmeJUyAjsBVw8L6Ki0yqA
kpea0tgM3q4hHzk16kwAPXThp+8dYpCBzDAd9zNXUWJ0w2tYtqhdq0u9LqgXGPoT
aDmn4OixpKHxBxS1AJzdG3tGReolzyJ4DvZJWHPkU1DjE45X3+rCdZRRVEMJwg1D
WdrbKX3gIKQ8RcsmidPTHBug8uhf3paU4pamDQn72/NP5KgTEbnaj86/goH2YxoO
jX78ty+pPLb3dracjiA266lwFHTLZV1ZFuQ6OT9gcK6hymrJji4RLIZaNxftfvCk
T+VSaOMVYPwUTdJE+2SR3xm0BhesVy/bFR71akfuYTbbHSx49OofFFsRkFVteg/u
vcxGpySoBusqxBuAItkJKhHOFcMD0kAbsOFvX0pMMJPS6SkXx9mHMunW2mAtZow3
lxhikxm7Lm4EnWP0LDDO/vJM+d3icpFrFWzQP8ExH4FWXhLJUYX1NXUj9MzuF1BN
mTUWVkTSSeG6yjx84TuwjxovBQZDvhD1n9MqopdSn1/rprtYuNHsM4u04y4r44qK
3ChpY/w0f4jBZs4pMwTXJ5i1SM0jVJ2LwBx+DR9wuK8yLAlhmIrTA2XksZU8AyTG
h1eNQzYDxGIh3xBH5H0yaJmzJzw7wxN0mOYduHerlO2NGwZb8kYmt06ZyhFbjJEl
G7x/xutW2XhjLCQa4PYoz3O+k0rFsKfs0BpaKxA4Pbbpa0Nn9mxToAAhqvw/tlnT
IAhZUbIH/GYd2mqTESbs1BvKZw6N6Phs+ZtGLhd1ft6dU2uxjF0gUKEtF6ANpDjE
L2vyBYK73X8NJEWb7Lp/ISChVV/5KAhlPFE3FsT3vefsP2rDgsn8JHLYnTNjv/AW
yR6N7zHPRPmc+0caZhdqvIbjgiLTsZqFcO/9nJ3B1e/KbuwRi94z2hpUcS/RVMe7
NKiIjVsZsgtolzDdLpHdDHuY7oi/dVqYKjscEVIUeLsja2iPDRrqVIm5rpfFb2Qw
`protect END_PROTECTED
