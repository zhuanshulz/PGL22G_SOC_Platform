`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
57SBtPVIRMdArgXf1fsJ9waTiCrcb9pqpuxAmSBrCzr9qqnUxsnTwayRO9ux75zl
7cTwadC8rvvx1phEcCioQU8YJDOABPP6XmyGCpNDS7i3Hlw2F8scYQywnWFk9rXQ
UwPG6AYmNRxp/0qJ8CLSt6hu0WtGsABbAmtcvchzbQceZz07VAqGDsuK4UOJAemr
oqvnMY14zoZIu7f3CnQeoJASC1bCgHTIDe4I+4exTQ8zGFgfof8tijK8951d9bQM
jXr9TkZGi8WAe9unbfL9YV+0GitvE0AToD5XKWA9b4LB2TUCUzPDMjMOZmkuAgqO
61NxIqRYHvKy2O+RpNywPeoo/gFI64iI+QHsJvV5dpBo8DIXMSfBaqT+xPQM+t4f
Gxdv1NhyAAyHbu4Z6R7kV2o98xEtz0xzPxdA3XRnUNsnWfbgvaVNBkEJ0mZvGBp/
WllijxM0dZZdtfFELiBfnSlgC+alhi98GHrsNdy5Q5oW3MLZDj4L31/h8ITkEYyl
I7nJ8zV0PQXyOBVqyRrt0g==
`protect END_PROTECTED
