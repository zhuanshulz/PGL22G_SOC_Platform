`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sEgQhaYkKhcbkjqqb7rSNjNvZXvWyYpnTfRHUAnuoJCdIqca62x6DhNEKNVUgs+N
zt6HTSSdaf21H9HNuDhKklnDBOoPhklvrb2yuhZe4DIjwSdNOhRMnLWkF0SFnNd7
7rrnwRsaEptcXEMmXCn0TfJGP48WrNp2oJmAzEDKLu3IPfjL4S861BeutHTwkVHx
0hu7UCfFYnXvxTmwoSzFb3ikrIZxRHMCi860BgHorEmxJkvlr6akGkhCdA7WVOTo
2e02ZzLSljK4IYBokxnQ2rROHwNmD+/YSvmpo7j8wKgaYCpg07EbZkMPNJ0LvJ7C
Wox49Ps0FsNqKP5lXX3Gq3+vuoy1f80dGKOLlUq7Xkdd3nBLqkx4gEV294+hsDd7
5LqopiGFTNNpIZRDV/JhDVa/+wllUGgb8jES3vZn87GmFYbG76jfSesi6WMjI3LN
a3Eb7zgvP8bkX+kHpRIuAIQaoyEfJlZp2j3unMCJgJ6TcYJyklxWi2ceYvfBgf+f
yF1qVn9rPpQIaap9wQw/DhioxukOzsP2BSG1Konr/LFoNNARAFpaxnhGFRV8Ywwh
DPSocagg3iiknhWx72jJv0N3Dd7woj2weIN60kU6QmOwbMiw719EogTT4r2Kl1LC
koHsyHzT/t3CLFaN23exhiegZIVOdgu7sUAom5vTQ1cG8V7yg+mA3COSurfIO5d0
YLDCGGBa1+7gZc+2xJhnWocVGnPedyTHR2/yh0fUvZnal6ukszgTmt+y3RGuZFa3
xDRmTvXdCehekjO4Z6mhILoLPDy+KlWjJpB4qiv0uYlYobShFRU1H3bewrf4Zr/6
3FpDV0b2BfkYT61YA8WVh+5jR9X5NBzhfuQejIM1sCBNVincNOmQTg2hPrmkeGK+
V8LMxPtMBZNgp+UuFLkJ/gG7j9LEA0Y/I3cPD5IGrW2nbmw1CamByAL1jocMCpOq
+9PF7qO3Owwhc76rBEgDGZOr4Wf43FhpJMz5VQp1k7A0nZ/JRBjH/NmY4d5jbUr4
S9YaSFCIkKvuPsSa5lIpM3NDV8rNXMkRcsS/YYVfAzYGAYKes/H1e/BvOEjtf3A0
e80XOQp12HRyD9wLi86YwTQzCkQCTgLNI43EzhAe8H+LQPavO7f5+s6LBn/ivz3Q
nBpY67JDtZvEyZTRqclzh9C+or7MTkNXrSC6gHwkZlsKt0ybFPkTOSyjRUfz4vZF
vPlwv1LqBL993ggE1PQsK8FuUxReLqp4gYI2POoIXRs8sTlxreReh4zvMfVdJXu/
a4uBQqsjVv8/i2G9eJ/eBrX1a/a61lMLIoT+mjJyk2GdAiiEU1jptCGLaeMUrqL1
3EKf9Z4YOAd/XjIpKfwPbELgkturFFt0DWfKd4nja0Yyp4FGNxliZAhir5ArQDrv
iVf+Uj7OI0VOD9VahFhjd4anXdAtTxAk7SYD+GtLv20yxCb/CwCUTcv15jvpY4oZ
mf6mlWtg/pd1RjXlpQDH1PyPo/mvSiaNWDbqzjQeh6f3xeS17t1WRqnHgOcaESKG
87DDFB6BtHzPBzWCfgS7aJ6bWn4+X6gC/rK0/JUTyr/p1OPj5DW48zEIOziq+7Aw
u+7qZGLsRLbbqfrqhrhktU6LNl22LZKeAEbMaOEbplL8qoF8WkM4RaGdJm4BseJX
BzfwoJAEDqbwmnMEZZ6GfAQvnzJncd1NCya6vBiqggfOgKh6UKF+jrD+urhpS+5F
s1y6Khbe/gj4spl6YwpkICkbUJApjOpIfKNIOuC24tlIxkOeOSVBQD4gOSEYfmL4
jhT7Sz4o1ngiAIOzA5WMW1bB4/U0RND8KSVlOSl8mfrOBvfLNvIBwp99+gMwRvMN
0BS8ODmP/jthll3wNzf/yohD74nBR3hJUBT0uxWOxq0zklwkDmmFtWmelg4WYfYq
7ge17k226OasIOFNlB2MpLSSVCKkJ7Df86Kh1+sLLAz1uBbKZNw1xlDeZMFtX0Ix
U2CYheztNe4fWX3IE9/+UKNUTzJitkNL4hPUC+PnX2cNg99gwwQUrWAVHbWbf//c
gBtoE1FEg5xnSjJ/OTr9zOpdig5CshJJCqMPTpFUoA6hqWUglOv5qmVHSbqVj6O7
rcnkVDW3hQ3+5Uh5Az2Pm3BR5sBROvwCCmKRdacak9R3gfLZJ+kS+jGbm07LUstp
haCPJVr+utxxtwFNElchFsL2clkXrTkMmJKxHrtqNOzfTQhbodqFF4XofQYGYAjA
QQ4J6KT4UT0gQPUv+11DDGVUhri29jIGiazJMG1e8z1+wlOwXvT+VibkYgq2ptFe
p0gl+bpMiV6iif4Qk7YPZ045dT+6g0AAqverjLQZ0jrPcFDEIEt4zoytV7KYNk+h
AE1Sk2Pfl2SZn4FeQumUaMpeNbBEDmejDQBE9ODrBAjoJ3GxwCUwI0P9w2rHjf+B
IgCmi071K1VQUtmFzzEH9sbVTbcem42i0KBUL93nTNasjy97KwyYju5mTrwBs8+L
TRVHpuTXfcLkywRA75GS2FHL9BNv96LH0eHia8wpnaQJ0gzEG6qFQPvwjFAwPqjt
EFP9XwR/boipTXV8XVnPhMFvlqvopsiL1nsDAwYT/CordVukA/WtKUXvJUH0Rdqk
DcleB70MbPOxwipv7yxsxXqeaNrnq+NhDP/qWBMJMUoZCFGbrJsNFOn5EE5ID2OG
/kl116GsjiNzvMGvWmUcmWPtqv7YHP6JlwE9iJLiVpxv0DCOdJ/Ye3pgYbolP9gc
dWEiHLQQC0zan72A+DWUlujN9QnrVLnGHTB/7aqDqmqdtRGAIRrUbJ/HnXt7CQP2
caNd6nU7L4AP5rt62woDgll7FWMd7JQKe7J3a71gRK2b4JsIEDGj8nj/WPE/wIa7
VnIj9sEp5smdUuDLzmXujkTRz/9d2o4zRbE2G/WFK2x7qeCsHqvbUM2CRIommgAO
j+MsX2ygLD0Ej9Q7QdZ9U3LjTyK5X1PyH3tT2B28LdzaO09Ez1ex2J5+Fl1kDlRd
UxU1eZ4dqvG6rt+fkeFtXDpZ4eeRqCI+L9iE3n7n5/HHrGe7r0nX8OwYAFI5f9w/
HAaI7soU8dxauc7B1kKYfw==
`protect END_PROTECTED
