`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zgyiBWe7RmugUuMLQMp3ezjcuVHyYeRn0Wip6eo+TckW3Ma/xPyNIuHv+PDtgHQf
b1PWQwAouqOUYNPCRJ3kZV+dmuJstFa+jSVACPk3L6/TZOjS0401lKDqbw5AAKzN
MrKHxPHLJRnGO9DBfBxjTO5c3Z+IvBOR/VAZ7U9lAISd2nSXwWEaCkhuNlyrBlSg
Z9WYxsfxD7nJmm51rgYfn2aLAD7/V71sJiHh7AudJPCF1Y1G3IijQ7DrDWkQ8/Ja
bYykizglofLwdSpAaYL7jWAs4KINnGMf+sSVDMBine7MYwu7sCCKlbUYJsHnThXu
8QBT6ssIIpL69b6rx1ofd2muxP3MEqB52siwsgn97nRbY2RaRV8bpwW8/qmkzj0e
5ttcecAp5g/eClAlg46vMcaTiwvGxYGMki7PJq4TC+iy9QbHusD04nOzk84j+kUu
0Rbo8wMFoCZJCOixbwzaZe1RZmi+4B0Uzu4yEE8jIh5w8g1cmXAGYBuyA4t3hQfl
7dIt1sVnU1aaZq4uTa1I8uxOGjd/2ugIGilm82zylGHnZvHx8FZGS/Fnst2gSpsp
Fx9lMX/TFiKr2T7s2hpRe+rc8SW7OWe00ACxkZulOabwG3/MYiTdRDxdKJ3IBlxP
9Ng649aEdfJSphgB/9AH+i71vAMC3LFxK+3PykvzMKWJl9c3Q+WLU0G7ergLRc0z
5JH1hcwKxFooQcMem9OYjJ4Jx0EIOfO9A94InRiITSuJGro7BfvCS5/Equ+b90bU
zYt0pYUWLNYx1hGdee+3rCHbAzeb1TZuaJ/zs3+qbDTUZFq9qNzQXUGQBh9Wk9T3
61Uu71IOJ0/A+T8Kjkio8VbiI9cAzZy15fHNGtj4omfNF0ijNDlVJtPKPWEfReVS
Nb6ZqxAKiJhBZw2cjMJLDvwSA7aMIRuxH5XU9UNEZ/pN9GjngmBOkpH6obP/R7jN
tuO1GRbamm9ex7RkVAEA7nuB0K3CzHmXp5zkaHsP5KxutfP+vIiYwpjFrplBVzxw
qoFJQbwuSwhB6aA+eznpslMyoXGIuitoOaN7O5J9LB8SG2norKdljH7/qU+kmDDk
YGlQF8tTN2t2DMzAScBLoihXhsxGSob5BlRdj7eFmq3/6XPuRK6WDRCoUxYhIsz7
RURxo+FrcquW1OWtHm83evliH2grHYjh92P2w4ikSgq4zWWSh8Kthhe5YccD27Qh
SnEr+rk84N8NwUcVl1UWpnlgy049Bs4lFfVMxr3VfslTyQaQmcp244Q60p6Vezbk
QDk651tJkH2Px0f2Sj5+Mj1eorV5zEqOP1JibEGDmlRpaqcvqPH7pxCc2WENrLzh
oj//1pYGJVV4k6xrY5T1m8/hZJZlUsdC2fGwoZja6c19oWrLdhHfL54VQZ7Eagsj
u7PkKOLOZo0/61XURoX2rVOPZD2eKIEmkQ+Kcv+uLifVv9+Tbi1rlWu5DJR6YEUS
bp9Dw6pDkFLF4ybgb2UHWl/gDcn2MQ7hYP97MdLEp0dsnmMYDYSXBme8b0kyhLlM
ccoByYDTyWE9Kk9BGxAtYz00icJqu2wcivD28//84VBRJqf2YZHP7B9DwYAoIThq
0nY8nKDn37Q7h5g056YyveVY8XQ7/48jRliXiKGdeSWa5Qht6QhUAClY4IVHDb9D
HqkWOvfn0nSkCnsjjv2c2JO3JlS6HOqSu7T6MD9uRI5oOabPJxHicemf7v01nh3U
jT8TKskAkxI3cnDKD9wkruW5qQtOmmhYtIwV7a9HF69dqNOzwylJMolObbrPO7+l
QPcjJgWim3awz0NX50FxmEfxZTHa3wptUoYS0pO3ghogJsCjYzcFi3BgD6tsDla0
YOH+hAq6VLqmPRsGNnqFLlaII/lMboedOr05u0bcak89jkVW9MmUGeHilS9/aG7u
R1TYV/s2crbaiB2L6wJpS6ndJ91kdjOtl/CKjpBcYHO/rPZ7/Ftzq4pwrx29rGOm
trgyR5fofWPeW16BJDJbwttZbLk1wEqSVA4evn9yElAnjUzT49XF3K3XRoLJIt0A
AKsaH8FUtrnefha1QNV8B5TlqiS3pf4B3+fP7BZbx4xQhh4zQljov+mHoz9nVK4Z
lkgRHFfdQegCRJuQ0Tgvwjyp1gZFhJISgzbRelSMvG80+uWw5vip1bwNEKWgcyL9
751gW/gJFbL/6kAterfd4OV2/6GiCL1fQAPhX7kzhAcWr0ixI1l9oQpn1sPWR5Ez
c/RxsocFEqC6nDKmqA3tjvoYerkUGmKiMmpeh0nzm2Q6Z+p9NN0yiMhQXvYnStLY
ysZQ/IFZpdjxXPdOhQD7xQCz0ZJ7WEcS9XdKqEd3JwW2TZgg/pI7d7IG7uQC0C7C
ecVEdSs6m5UEIN42I+zf79OXccEBba69ZW5o5SB0+5+QInNxA8PZ6zy3agUuEI7S
GZqFSg2wJv4dqu2AHM2y8/rVt2lwsSiahEujftk9F0FuKnNa6JdKAxBcpCETFEgZ
1k3TuOQnozPrdYzUFrabiCw2JfDN/IjBM9d8Lq8wrk7YqbHOElz8o0PomYEINsFA
3XbTvXIw2CcJl24SMR+EpvQisQWl9IyFvm0nZ9879OFsKLOIwZmPqKnWZxPkk0tz
F6tvRq/j0ZpJpBY7mRMoGSH9Eb/QA4vgZkl168YEbhZE0wNNL7eqP46gkdj/8JPd
f+99tzvVI7LnOTjUi/HvNJNK3i79tzH8wA9wJToXcRNX80bySq+f2eyBpV1wsJAE
b2khtkDdkvzZEDezWvpKN96gFqKiMmk86+IMZOxNU5isr8yJTKc8rYZFBsWvE+pL
7pvKmjheWvz/GIOw8CoE4OHiaQwzGRoAHCVNxJzeXWE2Kla3LJzodQgglIrDheLp
KF655jqgXJnYC3LfB5TkYkH3BRRu+kCchydh6fhHrlkxdvRmKp0NVYsjmz0PVxPz
vt7fTdUS55WJcD1ZD1oo1tc69ld+2/KGMqsJs8JkNbd/5Z6gYfqX1x0+6rLDFbzD
yETjnzbNxiApdLdNFDP8B7YK+05sr6BMrZARME+bIWLtjDEIIlbMXqiBuH7BFjnE
7Thf/765v0iygCzFOM1fHg==
`protect END_PROTECTED
