`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vAS7ABOL96nK9ypovGsjiH5nMem8nStvYycgAm76LtxC9xiqb2rRXZifNzrbtPXm
qYM7Y45FwUQlxJJpSYhehOBudZfZev6ZWUhwR7TGeWFlR6Drv3e0nFWe9K5gbhWG
RnbLjOYXGk8nPxsqQ05u5zStc61QnaDJ/QPItXZMA7/lCe7tappqrsTVk35e/iOr
NpNqyy1Rc3jooSjJO0IWkWCVbYqtXq0txcwedFsaLgIBqF058zn4Qu08Bb4yJAaO
X8q4pgGrZC2BqRaZIQIXu97lSVqxUbaI4rp2Z4rmV4pCy7MXQ3yY3rao6FxmoVFD
oYBdM1Vo1rkt8YKBVE0npE4lU6UfLlna6D9jXfB/Mru758Pza4D3TQvE7r/laNWB
5u1ayW0kCQeSCl22Kwr3EwwFMjWr+MOm6a89ACzVWgdiP27//yO2BNsrQWIefP0o
`protect END_PROTECTED
