`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1Y115y5fc0VtpVT0N6BD4N4Ke8RsV1XI9vsMWiRttYjK0+fLMZNzGDY9wzY97hq7
9p0U1IUT2YErB/i5LFPNtN8/8Xc7sRozMuE9aEjoaJogCLXFGkzN2QYPYUSfsfAc
BuHsXJH/Scr8RPOhYf2O4FTk4BxIgi3OniL4MPCMxmfc2yRIPu/9UcyA5T+DbtZp
odZM69ga29HM/s8ejWR3dgnDtcDc/RbtxkssVKrktOMwD+0txbLsb4nmGQMwvEjE
L2PcJFs55IKmtZwUAPbnaVDzws27JURDPhf4d5xnGfKiNIbIyTenGwMGf2xGJM1T
m/GZSdpxlH5yl2J3kRCQVFVMHMIuVdNDK6es8m8/TnZ4ofn1Txgo2N1wkSPFZcg/
U0P9/WW83HL0OGeewbZgYrBnLu5vDNQiR8AMGS5XmA4PlgxygIQwoc+XmxeH+uf5
VXhkbEboB1Jzto5LcPg/aHSqwdcTpmDaX63reNVsYMyFItKp5FWuFo5/1UN6s9PQ
a/5bpp4tTDsmV/RXqkiGQvofg7fjZrpWs7BP6a2KzAqrVNproZhcIhjRFe0Tf3z0
5XcN9atjiIqZPRYjwTJhtGKnckKatZnTLd08itft22s6yzwsy5p91IUAzNvjSah6
jMTnIKbScs+6MeK0hAdPdZoRk1OJVYkBOFUXy2NoFzhKiGB6k3SyawgG5lyGdwr8
DxAQiY+v5YE/r1r9kFoneFflDcuInFvAKOGNrC3+Q2FHCZ/FNHXM4buh1XCV0Vz+
0vjOyCeSePnhRFgBTZUSEgyVxps9TimfvE9wlAg0T25Wpjle64rh8JrE/WGDCVop
ejGKAT2j0DC0nIA/7TAQ6OZi8FTCMtGjNuh102LOlDfa8eGLNXYXG3e1jki6cQDK
MtFF53xNxdoDA2CJ0RndPn4++iVNbf+PyeaAlv0WiJ6eT8fl3IPXPQonCq0idq+Y
uXU6WEOHl2BBd/fdh2Safum8EH8xzkb6xM6V2ysh222Nib+ZyawsA54DYAAh+kz8
oT0lmUKYflbmbi/+JGn3O5+TJ4qDxK0SjzSkRODCE4KFxlpN9V7hZCHXLVyJyFVq
TLkYY5OWwbvQjrVl0YP7Hs854z7bmrqTaUksOTax7NYS8ZdY9/xDJjFXiQCgPiPG
1yjIb3K7GMYtC0IioOBhdcFlwD3QvNxnDXXvI6EnIhacuflrSxU/xR4cL0lRpPqV
RfZUUB3LRCWBWh9KuQt4SFkbwSlCAXurvJShYHwI+56TNfmz/SbpKbMeqlU9WCgC
MajWR/jVIIFvuavkHwaZUginZHLV8SZgVNyH+6bVDCa8Om5MW3dLLgojeafbIC8P
GLXMesTV0z/HhxhjudsR5U2KfmHHuXDMK/97EFgB5Ng3nxcaa/TNq17Yz8zCTJqZ
dS2GgS1+iUnisqmLBjLqlum30JAJY7VruW5Ohy07wMfGq9ZOin6XyFls1CU4ZPdK
YFqxIjQRpqzPjCkKwXmxKRDJUZSLz9QFYxMfGF+SKcGnxLHHexPEhNFgPyOR/UTB
IXOQnUsPecnqL1jQR2Lq+mJyZnjOCYSa9uQBfZrKjNekwCVLQmULak5QjP3/LplE
Wg1bb7VEvfBQShlFNjeKelACFgR6M0hVLhojgeEYzBvZLcoRoM7ATapg2pNT3p2M
zy5I2/BvCEJHp29L/ASUST5uBjugXEotJ9lJy5XJgBtoaB03PGOxonY7qhbgQ7dP
iZ4oYptMIXdBLzcm7MVPAoc1/0TxXfc8dx4tQxPkBcVHEU1GQfCTkD+ibkPNH1SD
cKyjp3FvXmdERETT7RdKElMhgy1KpuzjjDq6Pl85mU+U5+mubeLHhrTNT62cclXW
lf8Qk9aIMgrimzMllYNZvV5tHHTede7f4uQoZebUzWOf2/KGctzzGoYMmRZd14c7
1deuJ02k9zpTVDb4Iw0rER0WDzH8yc1DFr/IVL+GCEqaksMxPFsigiePARKaGH5a
QICp38rxNXW7Sl1fqhPz1s628C/MPf/Rpzmohbm2SbQLSi81TTcy0bX6Z4qGGObP
4kxeUvYNTgikoc0RJWR22mWhDJnLdGtzaJSlZFPTByPJfquljNWOqR9FtKS8EgSC
P6oqXm4hTfMEsXSr/cxXf+FgUVatHo0yR8KPChNsjzKgZHWDWkWjtqJYxkHYYSY6
2o/0S/L2ZeXASIqoEw4SgTMo/HjSDEfGfK46booXLqcLy7Syc1cb6l54P+8bNDn+
ViJ559R4eY/0sxEj+CEU7vMFT8bLhe/SXqOhZn1omu6CdGubEAIxViKGuJMuOH8E
bUUX6qbOzTnuZ4YPsw+21QdmC82lYr5CqV0JuBFq1Ei9whqkYDmXq789LPL56luP
izUy5qfqAEm2nT0z041ny0tPX8NgTCN+3BQ21QsKEr9cnbEhVNAb6Bl2lBjK7KMW
yee6F0rZmVaKrcELYnfOhQhdsPgCMU+b/h1D30YsAP03i1TLQ3WkMIsuko1GtJsM
C8gGzrBxJijTs538so5diFbRE6SoXVHEhkfSo286hrPPX6EaAm9Bgwqvnwhxa/Sg
fwQtiJ+x8uu79yV4jc9wFypCrhlqMZrIw99eX7jUZ5AFoypv0TpQZHxNwnlPnh7e
UbFbs7P++eL4j4zzgulhSHi14AZQDlqHAVyQfzfvHdYW659U7s9/EseSYCbBrP4M
qcu0nH+E1it1jVGxWH+Obik4Cy8CPgPupPVfC+5eyWRqwvQwcT6UK5vpzvQxgDYM
2Xsjdjl5ztMj9keVnqPGmGPUugnq651OZDaLvI4Q+dBPlZzLcvjdazzWzwHKd3Pi
c8TC6UBk7q4rfNF5BV/6Px7M68mUN59eg8NLiwMKZ6ZPW9sG0xXNLbIvhMT3cEFI
t1GHQ4wBNknqG+IQXT5R6kWTou1PlvXfIISrg5O4PSCGHDExTwNUUTuCeCKbc8qx
5kj9c7gSIXqyxWKL+AyyXqG+dMeMEOusrKWJrHn8zsqCQlqHBfhlq2WF2A+gGFzF
WNF7hL+DimaatXSXDue7BafBgvhbWiUiJyVrGCPe16qI7x3Yc/riBDT7ccp/kE0a
FiyYhz96IZQai7WMULYIF3pmvJMYNkfgY12GXxtMXQjmvErnPJK2/1rTIgRelDfM
1TvfEfijWdlmQ+CadIlBdwcSpJu0oyG8iEj4cGWZ3NM1/dn1YtyOz3u4FxI/e27I
aPpbhiMtUTl5H9P0EcgGPPjU7mcAQQUcHAzfNbk8Ei2wx4BZboeXJ83cMIeSPRPu
TzhaIhO6+zJPWRfG8QAz58gagU5kM2hrPB0gELucP4HVIQTfkTMEq7aU2yqOlPxh
WQyd5Vv83XvZbh7RX1OTK92eXcz6PBoRkx5hqal0wt26jAy2j0vqT9rU9nzcd7o9
1OzEc/tFaDzHX9FnaUbUYgUhMpcAEupsBagVE2lTMuHCfb1NcMN7CJSG58UeKiDL
Th1FklTprgxOR3tdhG/pMIncTIEZjQQdexgum9eufVDp2euKTxBfTM5s6BXqFVZ1
`protect END_PROTECTED
