`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PnA4MjAVpypqFDfym6hPcaWeirqA4209kV4kvwV3eO0nhBDVXFdP62WEy8/FpvYq
p6u6yg4ujXD5vnXjd4wkDHATxUIw+b0uTMrtY3wHBqm+6YSgBnyREOTC3Yjcm3qY
aTOVuYjs20rR+A79nQGrYGsogDFRTTfH5u1KLcajBPvhCBikBZtfZM43A0DMdJDd
rhtxZ/p9ecrsmxKLOYvbbmDwOZPRlZpbEF8qmf1GY64TyuoNeHydgPEhqSZa1yNY
mPb+JKR+SpESABfJqbyk1VxXF82S6MU9A3IWYe8ccdQnOTbXssIijGumJqbsc8UL
h11r83rFchvLcB1Vo+4yeA/AF5o9J4khnZk+aLNGUtvRF7OvV1JtU2URDE/TcCo/
`protect END_PROTECTED
