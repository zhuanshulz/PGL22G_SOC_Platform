`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IepVG7MhEHcIDKwa+1j8D2Nfzb+lVm5vReZSSbNjHdjHnxKkUMkshbAudvNhSQAB
Y/55TdPj502KvFvcVvuPvRN2mZ7lhdjoXqRqeNvD3GpmHWi2iIapUkZfIaZZSTf2
KX736+qmok+4mGhQHymHiiU1XkqMFPqp2MaN0dm81oCXt4iSOorFMRoUZacp36vS
Tt/hmPvtCaNN9RdxEUSF2JtSqQK7GYIS22xb0pqx8aqnEmbRvgOYFK4Ht5GkpY+i
tks/n2uHP5qiLcO6fjs6pm19S3lMSda77FzropGsGbW5v+DcHJCqjBJ4iRHTQL8v
XTccNgozlixzokr4vrip/6s9gW79Cy277GaWcJel5jOFlj3egO/xMVHz47/HWIA8
pMJ0ePmxYvJNhc1QfPQvWESi7fOsolD1I8y7svlPWaPeBAoeJ7qHskmzBkevS9HA
1qcCl8kD+sUWIk3rwpMUitd2kIwAvwpaQQaztK2OKimnWUSdbURqrWwyJwvSl+J9
u1VIn2+tg3hpeoxhdEcUl4o48tEob63pkRZIfyZ7HPFfiVhttE1QTePSiaMuIS0d
v2q404gD9Iav6kkpsQlomCqekuQIIB7FzFKvKEvUOUw56OulPxtKYcK1oSNMbJfM
u7tUjp3r80Lypf19HkyKj6L5e1dSdaxpswsvQ8vxhhSf/XJr0qvX7nKDYFrLVyDt
blkKyDppFl/LOFRmCyWIGbGQ2cUGZXm4qNp1VzEr+eZaXMGZMrLaJEabR65tSGHp
J58uSlGCr/e7RhgICaHc256+xqA3YPHa2w7p8mbVjDpwjs1wCsZ03Palq+CIDZBe
kCJn9c3URhfuceX1rR1WvJtHWssZQv/GBBKCKPeR2xkpIB1po+dSTnsEHTS7dzwo
/xYd3pXxexFpXib9WGclQPi50vpZ0Wa0Vsw0mmRJxPhxc+5CsL6gjAxo7zyiZmnA
MlPrAZ0XJJ9Xa5rwzQWAucQFX5Z9MgrEQ3dJIGvmakChIye+AGUOnjQtir5VkvWE
NCpLJMHR2LRenJMQIZMgba3BS0Zw/boKwD5rwT6La7oGtBi+ZOaPNky0g0kXbjoi
lkJsq00w526XqJ8MbZ9DD0gYMwuKX6sTx5N3Pa6Zwa+nQSlR12zLN56bEg3AByRA
KWM+yN03fvckXzP6K6o0JE4UQtiLwHSUyoRuZkkIejT+wR8+cHaF5NQUfoF/97ve
EPJxnajP0QRO8xgstkzLs8QGjnY9o9eKux7r/issL7Kyd0BAh20qSssc/tkUCwer
ajh8vQ1Yiz9jsHLRRABueLY73RvHV1eDbEGxN64JqKJEGCfczQZTCkm+k5cYNkXT
FX9QZuEZaUXRHeKzkm7nuXAEUk+wNJ8zhvqA6zNaHciZb0qvZd8oI+1nfZSMsKsm
CcnG+HPbrPbhLxQe9yr/fztgv0cdj7lYLs1xfCmLazaBvUHxYdl+sMiFjxpXvkRN
Qoq5Svv+u2InSxjisvH5itFiK9aq7+N7w7IffVWAFtEHguzNdXowRfc3LPyR4Gfy
RMme2INev8cpL5b+m5D2VsAq+sRgz4EjPP9cz0nYtg1Tc+qLOBhR4fy9oAhzcpyw
xYG8f0ko53TLds8DncKiLYzeLXyNqeF+Qem80NsBykq/0b8heYO2z6SSzBFCIrHh
c3tm+x/EWJfedvfqcwAMHYGdqMocSU5K80BerM5zHXg3UNMaGJVlbSr6ys5GFTSa
7v+CxbdkIOyKboWUC2jZM2LDclnGMjB3BAqFSjTjeq3tE6WKzbbnGN8tYuL2t62A
GXC6usji6ypb+FhUjjyPb4e6eGI4+TQzuzdVmPMs9NmVGy1w60lSKp1v/TpYHmJ3
oGUvIOe9HG2y6DHxmI785ZuGmNTsiYGrlLo2DWYIrUDRRkcMHJIjb2LUmcIMfo8I
TURdy7ObSBMJbGvt4WaqtiLRli8P/vOe5kiNLvkNjAXfcBIlcf/kqAVhaasdM6Bw
DE6ak29ozciI6ZLoT0skYYvToIWwrIeBVrXE2Pvacd353fSGP57JxPeEv6mtMJJf
zBo1/q2fvBmrlS5opUjDEk3c9iRg7z6e+re3gFnk8nE7sQCtWe/98SYhUv+H3INe
3Pmtarijsgy2grqrTu+cyRxd24xojFAnAiG9V2cMg075PCzqWMe1sHrQB/pavoFe
/EAlYfjfJ2E8J0UvF20/2QKKLirhJk+s0WEb31gHr//V2fnWXyr6Uh21ZOIyDeVb
1fUd5koMRjEFGLnOatK4SiK8L46hAtX36lo1EWHRA88lbdOaqKNb5hdR7LIu5F4Q
Wx+veF3JDS0X2sxG9hasF/gpKDSXiFepcenwNgFO4T/8+wg0FxxggRHdbKp6mXK3
By3FVaiDZVRPALujTe/o34AprzHejLAS9Ezz6cXDMn109Nt+g6Y6CxTNCKqWuYzF
dnz0hjyUQqg4UWJ4XH+jhTT1CxspPVVaR10gKR6KKVJD3Vv4/6J6uf+Lxw0EOh+T
EYiFNJzoywCYAUjBDckOMOmEU+zBcvZ5EZa5biXYC2pzU+yNSbZzzr3ybitmgBSC
Y0hQCyH2jBrt54nedCNun6gJ5gAMoKwDxUuKy1FwWxHK3qvAcmH2go06mZOxtP6Q
Sbey0eMWsoOaeB1nHhWHE2t5bj5SslCSGA8vguT80b3zK3VuNFUEZDXwa/RFcGki
J7N5H4qMr52zzY2gXaL5jooL4pOsWRuk2vPwz2GdAsuirSa2qvVWnWvhUeVfRJSN
ngAlJ+fGtBVMvzy55S8+dvIW5U/nC2H6DddphisH/TiGHTDod6MkAdJ494/e/TMh
wqhQGNsoTVs3mLrinGpUldrTdOroFPM4X/PrhOGiFHxbQfD6MvS9tr7Va96nqYbK
ehNrr9/2+bcVzGjXUDMqnjjfjHrjWrgb6yZY5m/VuFG4kngUec5PLoa3o5MBIbmg
ABbv18X6W7rwFLsjLQNwPQR32v7EPGYvN8XTQmD5dCHKPD9oGFJq2jpxQoLI3uWR
uUzPffzydYHfdiEmnWLqxvN3vM3SkcHo5ueoMQs0K69JZ9flKBh8d/ZNfrlIemDl
TwJFqsThNDqaGLf0/IZ0fa1z34WSDDDEEmb80g9K9XMtF9ztPEE4Fnl+kqEbqOP9
PVQ5wgDdZPhFtN9KFVSX0yuLT4ZaJvI9XPusN810OxNoJZVYH7dA4SQw57U40K1T
pzSz0h8Mvk0d5RhTts8/v859ZF9QEsl9dQsCkZ90eAO/k32/QVKMMjdVHny/9j3a
APCOxO9aMDrQgfIjp9rav9zOSZ/6sWXfg3CFAk81GLg8Vagl92MVjvaYQAJQ4RpF
3xwZVrmgFZ83stoqqfB48419XD/bpsjvHv/PLmirBf0qHGuNHtyEUNsVupR25rNB
6OuHKCNAgedCYm0BaG9aqdz00bN9Y2j+YzG4+STsmZ3v/DkwuWaXG/apOgmMGnIb
PX9Da5uRbSSJg187yVX6bYm/S2U+NUANSeUDO+wUE5t4l7t07yJGi0ltCtH/ifZm
vTQzujMFwTAwkSEFJKlbHZnMLxG4mletyjsCV3rC6kjPxQTEuXLCyeRD92KD8BCk
sixLb9lahLPbI+kxTz2qVTTeTNMHITXHed+aKQ/W3Te6lXY1CwkqdtOGLzIqqBz+
kggsUnOqZ9NtMtzWGXkvLsd7nzZKd/jEW8Xvhkdh3A7uZurSkX4HiCpc6a8j/DY6
YoBCKfMametQN8i8E7uO4dbzsCKjJaKvlYYofjevFjT7CxH7bgwVPsyQYdVsJYBl
DW3SwnhK+HEsWuiNj+my7lAlkeFssRVhrcth6qPONS6vKZkp4+3zVYDLSIwIyy6M
EckLKbjYhTGB/6iDwzK29blgt5f/GI5f8tbMjky7lYfMXAJlXIFjcQprXOMu1rAf
iFJhZrNMq9ttNn3hfEpWfX3vmjB3o3EgJ17713fUtWamoknd9SL5IopUIwfJM/rP
1BRFgv7m1hiHX0naAas9bt9Hzwvfhn7KK4XAxeU5B/SUr1Z+YXnyg4P2omjapaOI
+JLiv+xTqhqmC2V3+4ux0+eAYJuSPTAawDuw7ybOS+DpOUDS3gcCvXg/ofOWYD6U
GJ+luIZ66u9taqaqcHDdtYIC4NtCtzsyccOzIHAQD7O4LyD8O1hZ8DwEJ2wsMULP
FTpUDcV128F6dC9MHbfZrCQc8o2HHsWT5kP02xMce7wv3SmIw09Ei0d6qvVWUPsK
Uo79GgjXanAk9PRprQEEnblQEzHBT6UbjF7LIzDnDbHwDc1D37A04i6vf9HkMwI/
hQzaM1QAZ9CLYkG6TYF1at+5MXkDzgets1xoSTo7kxiyIIeXOUdLHcBdk7Cp8HFG
cFNK90BZUwmWFrUpHiHaLHRayp1Ua3E4pqTIF5ot3aqu+/e0Cjr5y6MjzjsAyeso
Sh/JuXaOtPkAZtwIlwUyzh4c2+UnNid4+N5e3xlk6G091uwU55ggE/c+snq0i4sZ
54rCL2hK9/OOycezH+EtgDHXA4J0ijckflRwksaCeVzG3vnEJiNO2bJSmvcp7OOx
8but3ogDsT2+tg2nMNuIC1WMebrwGicJFFz3fmpc6fwB0zsb08UJb62/lm5huRb+
aDnQ01/crMogxb5PVo9KVKga2XYkPvrKdnFhoaCBik+BjyxbNFRqoztPah7VnuMW
za03aU9kOS/MrDLksIztkB6lDUvHHUvmNF/Sw4gzzLqbeuReqrH0YiqN0eFWcsmN
L4fqNPlQSuzfErx6+Gy/M8Ns/gictV8vx76oZJ6GRQ/oRDE66anNghLUl00ICttN
ewYpM8YvM6BcrowBrGhwZRetoa5vLqvXhaE/ytUi5zwO0XDkpD6DF0CFfrsLKEii
4UXrw/IXh5Oy6EtuiynFTPpltXLIntbJDmrw29trpszoqZVw8v8BTIkVUQzvoJkb
cnfsZbmMn4z7Q+FiT0Lq/YOZuOHGTGcJrMXkk9nBz6kdiLwu2sjM5jfP4siHWAys
dXOV/yYzApzcgoxzLvRPyarlZ+dXkg5IjP7Glfd5n5wnVJYr7GRyMhn0XJDuVaNw
4hMazYiHWekYR6hhyQpVf1uqobV+LBHlBgmhvdv5sx/vJoZbYJupSPHt3UyFIbs0
FWv4dQ+T8sK4NHns5zOiZWTIr6LzdYVKYuHaxd58kEulCSfCwzGqStsYPBhcatrU
5gAzB0Nthp13hIpLjcVExLSoiLuvcbVWrA2OXykuFUI6pOr2XPnT48Ssm80SUXua
18FdM0B4Ah0+FtCGKR4IYFhfqwVCH5nDM7Q97BvpTNLFd9ikgqGeHkQZJbUQaCOR
AZToOw4WNKzgmWUeU7q5hq8ouJ5daT5aS1Ol/RTp61UkAgc/6YfWMSAFfuFok1io
JvoLBXJc3O5zoNl5QS/g6px0uYW1aezWoopGQj6H3LxTr1LTFjulT0sj/RnI/N15
/nTntro05dTPrgQdr46KcPs6a+9YGoAC7B5g3u/yKjrxPTUgUHahUr55GS5ee4QG
Xkyqz650Ka/FQ1YOvpaEcjTc2AMBa1r2LKlpzt0wtWGTMU5nXx1xXXmq9rPXjHXb
QTFDWTl2VNSrIL/HtICmoFMgShnVAi5v7j7in7BX8bJm//D89o8zFunhgHr4nn7E
O8fZ1oY4XXm/ufRg440rrRWKOGdPm4JS2d2zn7swTPeFEuBHmU+Rohzpzh/Silvu
Bie6Aby3yLhlUSbuT7GTddfc8jeZfYa2JE3cM6xA0bsMUcyC6tOGe8c4r4+0qohj
OmTSayrdBKQuqSWPanAa5MQND7u500klOn++DsRG/1e3lFE8n7yx/V0+kLW5nRg6
ywFAWZ/np0yAuMj7S+5zLxZ4nuExf/F2alMnOoOWPJDMmtpQDvvhVcvlh5CzJc5X
d7ojtbiWdV5TX/HHTn0Ei1lDuW0mxk3/XdRuJ4HZdqcwgxjeAlyM79wrzvqe+rxZ
KJmLqLJiJ1g4Vy3yxZINpYRDUQhjZ66SYjBLPzVn+I+ZOEeZrUeI2f5OvZonDJf3
t9t3aMfM793Zg6bIHSRc5hhCPcI18kPF886jNho0OQdxFTjar++C3W0R5WbYJ13I
sFb3IaihBpswTRRskMt/qLVMqYAsX52+8Mn17rCXL7kQYkl6iKwrOCq0gYCiZJ6D
WSYv+l+vIv6zKD7wRKKSvH8W3GvoMsmKXO6DYpC+MPB+LHj0x+69HXDjgDVRXh8i
NzOzNemkKyx4W/VMJlkBpyDrAAOfs+nBljE7XTp/cJTvapLS10M0rW8fATDEJvE/
6ksS3bS/JACynTCO2spAdnaw6MD6cswiHeyG6+w4GkUGMS3dRb2y8yyy8sTCYgSp
l06Zy2GNRx5BfRG6uB6qk3hlpPHflLdv4SUD+s04T0UGrbvkAskYUZsvlQCAvqa9
2AO16nfNSXbKJgdB9yLFfcafM0Spl5/wM81AsKorojzQ9buzwYE8DIUuM0i7SSNv
x8zv/RezY3pwOzyfrMaN5Wv/ni90JeXNNKywfL6HO+mcG1m+cbmxuiLTZ6NmgqY5
EH5AJ0536Riey6ts/Iw6LUCv3Ch87HHdJ94ARatA6/bENNaac95s0YPjqimMLxFh
+QpaFQWbtfjk4po2AtFRCDG/+GX02nW27ZNWeobq7hTobQeH/b1WFfPSqnXSrP9T
lTb/9muZEyx+8PtdJeyRD7wg9c/sqZQiVXfeMpsO2HZ+0vjTgoCw+jIzf5UFEKhg
K1kZiRVyvWBdfVPBwPt16Eh6nwMAwFd0/YdDB8CrgL0Cpq6Z7/lobQQGwtsJRco+
9BvowrOKNtIA2faUW82JDHRygLz7XiHEIdxzSkj30+SqdD9Ep4rJFcDgpj2BOSfL
PK53R4kqbUskNc5EGdjqPXmUrdLblNiXjTyOXoscLv55pWo25ah4AalSIkD9b+yw
2bAsW2YnHUr35cjA68Zxc4tGllHkW0g02rhHJZhzKAPo0t9sJc4M0q+Lae3d5NqF
NvUc5WMxDhLapQHjNaVwaKrTvVxQD5LMevFTwhcRKsO56VeT3iwug7LdF+LRFiQB
nuVMauLpiOtVXt71z4e5hkE9QAg5axW1ZvnB+FqullXsvp2ouRF3PF9Hm93X8d/z
ISi94HG5pYyTrSnh+SAuFsg7fwoq2liuIqxJhmc+FPjbq6CavovMc2sYTmxjLXcY
OeU8pfGAnaWxEbYPMd3P10z6uWFtP75TR3H9q1RBZoFaFI7r+A85kf4X0Yyzk/Oy
S8/dVMfMUEHYrvjoeLNritNT1eYNkEPqysJKDekL4lAn04SF+A7NFRdmdsD/nCEX
IjM8S9oRfpCAmIdcbKylNDUKIborUeUUqGPRQv5HC/s5S61cNQ2Hogv/V8NTbky3
L8CwQmw+DD7eiH7Rc1vLJalge3Oo3nvQFWOE63/Y2bFlgAUMLJiqo3vHAj4RKQho
VI9yI1pkdQkvivByCZf/cS0dqjDnmU/UjDt1X7xWt2CkwuXiHg0rrao+XG28Vx7r
O0hMeWF4INzD8L/LjAg/lm4cnARCxtxd5SEnJgQ6yMXiUiHLHkTU8EpSpzHypFA3
glYErpDyy6o9DWVKMuFTO1BmSPQdXQJKQkYlJq2vlWmgcVlt+Dq5F2Mu29+ZhMp1
0BOavEyeZt1OPVosHLWJBGTi/ct6HKmrq33fpgyq/5nZsBgvIm/dfrELI6c+3Osj
rNInRqbwLTXVT7HfzOi5M3EpKi9MXKw+zqrhfRQ9rSa7aTVDwOygpM3nSPYRVtO0
pf+oQTknB6087zF44+5RGkg3AtYeZdi6puo85JOOhIjsRDbnh1VG4HqaOm9bvaDL
ZXOqhSfou49GLCKt6GjgTt2aEBf+V4BWqcDw81I/mulW+nN/v9cYu9M5psKcCdnb
QeeCBk7CLBfemU2GKfOu41bBl+O4MFCv2jaF4EH/d+/vRVV04DDmT5IGhi9wVgJL
bkCPkFvz1JutL2rqSy3zIpbehK8F73rnW0Tpmgo35ZP0cEJAEXgoKv1RSSqbqSOY
TheY24J1dJhcX8SGUaca6jsgPRzyHgKK/HQUME4FmJY=
`protect END_PROTECTED
