`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nHtiVZlSbuslyoG2O6kbe1uhSgKzYQtrFKqjnloPvdozIrzl61cXaUWtGo6bjRws
Lspz8KD/Sc9nrMmjvu1aE+hSlExLE2rqdrawnKZJUpAajKM/8pRryNUgGQMLwKUa
S+Bet/Lb5Ue2fb9ywLXORw2N5kVHkjfWusIS2X+On7yZE+f4G1XHWHzJNzfLp09s
9peIaIzrOjhCBFYF1v2BNi5VVA0EqUM2guwFpRO0uv04206J3aaKNV7yHfl3EWnO
I0ULBLqh9fIliZV43kl5UX8YvQGx/cLEABvQxtiKvbwvLI9pjk95+zPW8O4lZVwT
+krHRwd6b7/Yc74gG+kmcYxPpy5kNegOAXzawnq611u+M5wYW8G8yyhkTWFuebp9
WG67tHXvSoI3lvsHrkLoDfdk3TW3CneuY030rhqK0vv5ObFB+/wEIK3drZgC1HEF
XVGx/ozJ1Ugqdls7g3ioZ0G66R/kfOR5nJWApxg/jRBoyKT82i8+Et99xqes4saa
hhj0yz6Dte6NBXF5vPI7IH3amanKJ5DHh96AJXnvX6APqN3OlGN7jt712l7/IwK/
Bo8UreepBrYcyfBqfZ8DkeIqwJwamUyjr9vgkEOY+t3Xd1gak2FYY9z4G7clSXn5
QVbLO3HsKofBwu6icI7H1MSnAsUDG/XPQUaudBbQ7AbVOGHc+cxUuSFFoFrz05Wd
qv8leVo6W700d9DjHlFzzyWSfKfrXztjShmXcZRkqowVaIFexRgtI9ghjVQipeaT
RzzpIYcWFuqd9pgZ5gFsVzhKntJYX0FffjxRHK5S8Khf/I2kXqFP5FqkjgjJo/dG
vid6ESc8IaL0POx1JYk6NqXRiTvtL1SFIRKGFqkTSg6vkcNBIKCdhwSaWqRsoXdz
jGaUPBi+FJbtFgW9uCmdQDs0woqRTkR4JfD5QmA3//bS0kuA6lumhYEC9BAAyX9D
xzjy/RkJmjXkzssp7I2G+J4mDQfUik/Y/B7/pW99AO6LM/pk5AZQmCXvkLf1G7Pb
Kz9HJRxgKgzWAxT+JFMnusHV+dR0EJ60MgxRBwIgPUV3xzGk+x2aaxT3LYnMSC99
ZTfe1SGqRT35f7CQ3wtI32A5CNTJWmtZ8W1E8B1hmkzuJwSh8+INtAPhkXGQypU7
UllEWfDJCysteOBS9G/KQKcrRXbBj34+U/S/UBZ+qjIVMPESdhapkqBzDYj78kRH
qSGu3maR9u3ktQo2hHKGSgCWKXiuF27+4DFaUlKyN6Lx885TOpWds6tL624oESmu
J96xPFrqJ7Cz2A6bOq23ISUEy5394vv4vUv9T3yGWYAXpPCTKxjG/Z7dqshBBzCl
fB2y/VEws4dERihBNyWwsIELDTMzolYkHCr/taHGqJnUMT7watd3cpDhIUfm6e9x
13Mljih+maLxnLGAS/O9oPeTyBbmqygXxAs5l4JMF0kQRyOQ8mc+/dEJquLl+muO
FkKmp0A0Vqqn073J2oM9pI/Mw8SOruyMP5w/w4QLmPfmG0N7sf/LCfPzhCOtHM65
TCVFfQxmag+7DGlwWgg8dWTFul/kZymq3hAuuaLsuvepRrhW4qgsu5f2ImudUeGJ
Qm5DJgOx/JelFJhbU4DthyDPYP098lxMJNMzgyIMheIV5uU606mBVfZ1nonBx6NJ
7qQ4aBlXkZW9UIH/bM6/XG9zDVsAM1MaWkhHzbZCuMNarL2PgHFMLSNFKooGRHMn
L7Xq05XuchTXM6OmtcvOu6PmAkhC9C+4vpZO9qi+IwlvaE3LEGClZSKlukN4gxda
kRUEVeexJg/3oUKmUUOP/ENTou8LrRqYflGhR8maCR0eCoKSlj1X3EmqaMJbzxQE
HVBkwkiGcE7/MOQGrIvK61NhHaKGSOYc65pn/75iug6CyhehfkGok3A4pWZ3dKfC
1ScyzDxJ2nmtnVTbA3VOhd3ds4dHcrmBWrCAuGbFKRSb2Ez555YJdFac45ShLvvH
FURGLsj//gUDIQxXzqxYp6+gSA5tQj1VHMnOFkYCcnji1IMbIB7vpcUI2rKjAqEn
is56A22Dp12iQuz3uRpyO2PcC9E1kGsKUhrZwgYLE8ksTY7PjL6HeqZ6zbyTuZy6
DEWfgxb2DU15EVtAcFjkKB9v7wo48r19axG3mQ49nWx4TM4jXMMZAnUG9xz+EqyQ
RddokVFgFM/+koSmiaDY9/t6d79Iq62jUzc4wDIsEuOfZC/j8BV9ALPIuzz9goNY
+k1adjlAqF7n69S2ysnQnDPbYil4ONXDYJXUV5urxXme8VPPXzz8MuIMjrqjeZI2
GOdDEb6+ITQCnK3IduJuWWcyguuzNmhJdrZvPDfnVW4Hip26FYFpHJcVG02Vr/Gy
UEZlHoZTPUk2a1pF5jmegtlwlx6xnEmLgBYFpoh8sYQeDH+fG5OBHDcxjYZQYS9D
pEREeYSeneHY6eekMkVjOVQ5TVwans4FBBxNY///s6jJ/65epduSt1P0PP5itDPH
DCQpEhe5CTu53wrURy4txIrJLFrTynm2vT0YAzkY+r9jC+OOqQX47QLCe2u+8Y6l
FUeX8znqulcVHGr1def5ji6bs6mtZd/WUlGzQpu8UKIeFH8TxO57a1zaKjkuCZC9
y+kTfCHBCrAgzbPB6xlnD845wVTCrJAOpulLOnM3cBErrptp6pk5NK7c0ZHBE5FU
NpZu9FGeviGe8zanrwHviSDVcwHHaL5TJVxATu9Rc+eEmp1+D7Hq4yDubjHqr2Bh
BxyQk8/EwwWlDVrQAtfd61RIwXzavvrxlXaEMiSXNBBVJ6FnZ3elomtEn6OVikKO
gdIAqTUae+UXMd9g4nlj9VkP9OtZ2T1BmJx2RQZY0RHmpyBFRbBuS4x0RQHFucTm
uoyH8G+xGutkzl63QSwJjO4DAsU/t02F8oC8JVBPiG0JScuBkfhF8C3UmwrBICcc
NW7ba+LIV4Si/0aegoQ9glEfRQ53O9S74s/Wa0zHU48TjdWQJ8UgQ+Frpj0Udfk6
ow+JdESGknUFa8TpbKUGtRKWZgLHvTXIkWFi6NCq9X9gfO9Rai5XQKuQ7TOAuINf
XShgFbtYgJTl1rK+TIg12Qycf85ZtpbpZoTiV8FN2URBtab+7yURPTVW0Ltdu8Pp
5hvucXdUMRfqmqFlt/UYxkAPSxlChm/XHcFKk+zdvujUf27xVoCBd+oMH1Z4Qj+U
dtsjDKOWsDaWlBw3VaZVAN70fYxFS4PvjD1DbAdFpLVnIujENgWitytJuVdP5vaK
ELuAwwu/cySrfp2DjAjxTDXwFWH2oelyTl3rHvylGgfMPZuKFWSMpuq65Ql/W+p7
zzy+cjYjz02Kxt1eV3OyztRb2q65A+Hc2vQtdsiDhobY+KAngDFYYtfRPPShK8SD
ppkaimSwTUqAvfwfgZbVt2LqxuL4RDHjQSA8ZotbCLvQSVBjkJGPB5v8iMfHtGrU
8xDxNqe8k7uRQVMusFDfiG0SKL8E+Cw/EFmB/sevWWboiIr1Dbq+zD5t+G9O7sNj
+ScwknfjsBsB+hACyWKmzFNKEabF1xPtdi2vMyDZfueMoFdb5rEnU4jVr3zMV/Ki
NZLFjADYmEExsZlaEY/4NwhjU3fFPro48Yy0Rh0h/wxGWheMN2O1td2Qa36i4Ms3
DGOkNzaDgce3HuPsDgeFvZcgnyGFG6iLx0cibWWj3NP4/QoFssCD5KGZytBwPD8V
zV5Ww4VUNtN1Di6pHy8Km+xYyRXzRakdipO+zfXW9GuR2x7tsPgMESN71sUYAoPA
/RVPG2rqo52esEnzaU7CBukVHb+hLVtPuLPIabZUI+q3KDfAfcEoX2UvJBYdXZR5
ojFNc3PlnKaQXNLQ9Pac3gcCTx6ZYPk3F7/2yLp7HGMddL1DZaCPhR1DxhVRoEYl
sVbYVyo0QXi31I5rxfIjqIXxrpj6NVbZ7zAqZP43mTKJjhi3GVhO4e/X6+vp+AKs
mfiGGV6E72XCn5qCGupMvq5yR9DMa7ZXS5/s0kEErIV0dkZ/pfkNTRcwKc2VsO84
VTozRJkbZ4doozoxpI3SlKZTHHIRfsUhPfzn1a6/8E4c4El/0C8ujshlECqnlRuk
ftJWLk63o7kmiqXCxREjbPqqIG6UloVpiSHz9B2NtH3KcPVDLfReULToRsiz2IzH
h3F58rjyJg46h57Uwlg55X6ra7ie29b7CKlAF4RJPGolPGTjShhXAJJhePYKoNtK
LsQB/jiHnl1Vl5dFo8ziOQ5j8Q6Q4Eusuz5j8WPQm/e27fvIRt6otZCdGJLrCa4R
kqEXvB23kp9UtGk7+qeePmsWJ/1HoXdUvw3u5bW7xN/vRhG0nJqVX5uUQJnFGKO7
zu3CMHX1gVDpZG5tsbY8AAZnGzGkRuEChqLDHNy6AVMeggqa4J+JJYmZdfgwfQDp
T08Ogz+021o0UuQop4nkaeAsXClOrxf4/WBBl3RwjL46WJZOG6ZNwWLBCSfPfZPI
hh0s5nCPgbNpQFz39pU/I0pjTvpXjI3OHMCEF5UO7ZH39m8b6JLpZYfrC8PH4lV4
QBX99DWknETnRaGdJIO2fSgQabNVRAhkbaUzFfvRXkjUfS8g1OaCzF+NeaezcEud
wvGvebY4gO6MFrev/2cmrVyY/0O1xE48hvIVeFCfZIDDk0EbcwKtfy0WJ+uZC86b
paIsyXKqKyHXy2rvQKGAPYW/VaUIcBYobFXPyTDWDK68gNmudOkkKT5ml4ssLmfK
Zby41ajpCeB9pYae3Y5GPgOI/e1dSjux4iCMpCR8GY49895t0rxzIqECK/DkaL2H
E/AEtBf7dulJvUv1rh2XDvQLLOzbnwrjHHpNdZwJswOolUPGV7tFzjS/88Ufl8DF
3oXf7d4eFVosPL8wMJujiS3yGJ7RBoXw+CNkuWFrGChxvvJ0CvinuFV4LYicHB0Q
VdDiAoe0u2GAPAKGTD8WuRtToL+bkvTux45TwrcNZ5OzAUCTkSkgoGp5Sbdph4XW
HdIIUxeVPPFEvRrc6wUBYd0TeHK4xLfv4okJrO4MhXvDkxp9Tdex2FFgD+R4fK0y
J9LHAtJOnLZ3XUxFIp0NjmIiHOd3gjnToMSUS21l4a01m2JKHGAUz92dMZCqp7g0
heUvH7hvaQH2EY4YuuVsypKEUtLuk9qeuKrq2aD7UJmxDKkRhSKOi+3peIxVHkt0
nA8j0CfynfHEoBC/4YgupLHop47QJp2swe+8HK1f0gFm6t+F/Kq+7yXxTeAWwcYG
HRhVevV8Q6dYe82+OVScyvwoTdH+J1X/AvuRrabPM2SnCAU1zyaV6oQokpTdO1Bm
W8cBVQicbhWww0TiLoCCk4G4sXtLvd1OMNm4o1IIkp0/7PsckFwayyg8MiI9z98P
hMxjBJ5dFcJh+ZFyFiqgzNRl8WFjUJzCG30gqScLO8cEX88nGvRywK6H8oocalt+
19WNPGtubg0EBd6Xu3LPN61wZPnyxmblJghWCM1FUKdaVOQnkiq/kCzdJmhGsL+o
d4GmSVZetX2Z0vI203uV7wuEkbWETqD58P5j2uTTbqbGTQBux8RcYEdiWG9iLBq/
W+/pHJQ4txgbNAKTfXDeKAoImr//saHllxPFloXh0IAWkHtXZG8sOOYlsPnXN4Ep
Gb8GpqVMP0wYV0gP2tKgCWughw71On9zPy03u/WMLMoe2s9p4uStjXZzWiQFKB+O
kV2a9dzMJcaoVfFcrg98SCfyNtclFI845UkENFL3+DizczhirxPDDLZJgvl86XM0
gk4HhJ1spr7fNzQG8FwynWxDvo1wJzQEgQtOp4E4LEwb1T280nN4XiSesi4Qrcfj
CX1DvIYg8+80PyJvHTE8GU/5wGRio5LMDXpE7m2Gz8kpKtH+dAHN1z72mh/RZysI
TZKhKNfFEarQACqS3Vp/tg1rSgAm0v/RWvlUx3WTFa+bS1jlKOy+Zbfpa38WMD4w
pkNxgPfFI4Ceqf1QPVocF4FGWuGVwHBmDalV4/TNrVEd8l1iTCwWsgleqAbiq987
7mHIcESfEKcNwnJOZr/2a1WZbX/bYF4lW1ZXy2a8RbzG7pCP+6tTVtV1SZArxdq0
jvSOrW6FPQkszFjeAOqBtEuPm4knoXTqewuRM45a40LYZfGyH2z3wWtIt4VJ3u8H
9m69cXuBKAg9ItLo4kGPQtNX3qWN01vZavuKsRykhLA7rO5TRpxUa9BnaM/Tk1kK
mfUaDI9oKcUaIfwP2BtDKbpXxnX6G9cabp+7bL5HzrMd0X2YrT/xKlSNNyciEti7
VsOLAKD3FmjiwQZbZvYvN81O49SmrzbeJT/LnOKQmEjxurbJjOMF8gkgL3fMyqcf
Aeiqr9nEHs1tS2W3GnD5XCVZROgsQ7d+dFycXX7d9ZTdWcQtGzhvIs+/Pe8jCtLG
DFuDcSvbmp31zd7gG3GkEYTMAtHpVNRpbDC0oIiGOvlsUOfQADwZ38g5uo2cvX1U
5uTiy5xSyAenqwEax5pmrbnTXxJhlOUcfkdukbKt92tdRokqZLaJMU/tC504Z+zt
62WX82asF5eD9p4VgUKMroJrX0E+woeEi3CWjGEPTZA6567Ef9/nOH/sZ/DaRQEO
rDfIFvbb4r5NyH29HxeHN7K0X6YHVcFkVF+A7p2Dy0osFg/qHQEayXtd8+fBuOON
tnWmYgCHTDAgBD8sY3aDckvUAG/Te5t8pRFTayScXkbOyuBxtLqwwo/rRZ9V81Xh
gvF+m6UMj546t/rAbejCl0b8feO8oaMxTbKFmKT1p7dRFGmbo2u2SkC3Plk0KP55
7Lad9nhKjefZK8bue1ZaFely4gLgT/96uJSwapMJiZA=
`protect END_PROTECTED
