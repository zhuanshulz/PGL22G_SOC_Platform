`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6/NMYW0P7aA5fMzd1sOvOKAGscNcNDoOXVpq6G+5ZPYKJfxn3hpkd6mTCZE1j78Q
txAHxaL1HbE2YrrzfAd7obMNaCs+ZvZu128d6jMfuW9CmRCFFHwadilllir+MYay
htf1HPdDKH/9pXT9JkXqXx7jXVUXvi2JLTKiTxCuJpGP+PQUSaPlBxxk7Xyj+oCf
YGMjgyje5jnL6bExqHKX2VVL1lN9nXxiwJXfMownD/1fO82VTO6WYArKu2ifmUVB
RdT3KJ7DQ1CXg8k8wG6mWcMWLL3WGiQ6uOLlAfmn+D4SYDj1u7o8nh51Ut6fJeKl
0AwF6HecT1apeC/mR3OdW4+LLxkMD2cl8kZ4qu1In2XsGFRkKoYyMoqg9E4N2qh1
bP61MvvDyJ6HiobmTZoap4a6mKHd5mfvpfSXfuNY/lXp31Jmp/oEYxRMXfefB8SN
ihvIc/7WBjqRh0mdK2wQfhOElfcjJ/h7Y7UnWy4IhUzUva8ArjXBU3qnVS4Fg3//
olI/Pl+Vdj4WU7gwTLEGGTzJW2d7+jo55wcOErjr7kqDSuvebqCSDiVIWRJr7gIm
FhYPCejMpXR76RMbC7TAmfA4tskAELDmzGh16ILh0rGtFuxbPct9ebdNPAlL8r4w
`protect END_PROTECTED
