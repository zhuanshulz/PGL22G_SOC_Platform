`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hZ+NRn0wd6VY3SIyH21OAPmJ/9eBA5j5uQffiMWkHcT//yJQMKPDGhArLttMOtVh
utkSILJAf98qGEo6TNIVTsrTqcfFgVFnhmQVvAANMFFaSJ7nyU3V9CbAwum2TV3H
0TO61ihYh0o6m3hY1ApVgr3HLRaSLbGqEZh1FT5DpNrZut8ZtLwb9PhIB1xh5kRx
tPoja2wXxaqTSYH0hcAulE6nLO6OjfQzw1dAGg09+M77JawoW/B8DfjtgDDeok/T
epB7+XpQnTDpeIzlirT80CiWoJJgCAKfNPHg3uoxA04hScYIhwY0SrOX0/aXtCF9
B4p24PEhFUW8jTRZjjLqMd7YOHrm8kiXA0CbRsxkJpoIkJtXE8pAtjoTmdLONZUv
eZGsZ3v9lyLWQM3fhF85rBux70fUYtgCU9WszBpuYIOqlIVwwkJ/c2551kPbXROZ
s5wiOtobb1+pI2UnzBqe6MHeWaURXiahPRimhPrfdozj/rgJufkgC2varTxT9T+e
6N1zsZNkaDewQkqEKDxEUg==
`protect END_PROTECTED
