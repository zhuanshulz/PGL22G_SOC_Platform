`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eI7F1rAQaQFAo+DtwBLYc8hnb3tvI+PYrudrQ7F+oPA66p3p7J+0jL7zM4AGTFNU
aBydJr3e0xr6AtW6FDIT53S2gloqYimHTHhUV8feFSxEs8qLSKgCkT83aixFVM6s
97vDKuJSDswPWo/j7V1xr5BYIKj0PHLmz52w3W4gBpY5U3HCE/T6NnXEzkPS8Qjt
EAH/QFl3jTcy+eZuowE1Od/2aKtWYQ46GIddtWyu7djOaa7hg+4jtrgBsb+iU1Ft
W4EW3K59FBVcVPgfpMsdA5sHm5INEWBnwqOC3/Tq4Vwxn4cXJ3PS7iAhvADeasFD
Yqu6LysLzKwRg3U/Ha3rI0G6XjcjnfeLWjxyK50nOALcl0bWv4B4hGcCYX/SXl5e
2JE5rZwjM93NXaWu/jQSOTUP1UmpAJACKdbN6yEIhntBnv8olcxwGvFt+D65ClrF
WjVDcPKMfBR+znWjV1MwvUxMLgG38h8ODppCcf9uXfJLwagpAyEOgRHZxhyiPgMZ
/iL1GiPCR57Js0bFnrrH0OwDdtjBd4Idx5ox0O9F4/Ty6LmTv1TbKBGgJE8UrqGZ
ND3wgFNP4gg2cH4fMeLY9prHkG8aJCGwMi97RwBFGDAZz2XwE4GtRz4d/Iq4+HNU
bAtjbeSV0oRVhZx5FK6eum4b1rDQik3t4o/CQ7FhTGpu6JCFBWNRPcDRUwOvyTuj
teHbbjklhg+fcXUk8cnBVXYSJsk4gFfukuN1tI+7BffEjVNExLhZVV69P1D8rXFP
mJz6i4hdYiz9KxUJbWeHasP3ciPXnNhdbZAOlikZJHE969eCNZIP3p/Qvq5eZFn9
9Nbr1mgffy8MBAq7YtLaUAF+6zV2Uv1O/S69F4UMsi9m1XjdhByn1iOIY9QqvCrY
iu80FXNbUWGRSfZWqMS4sJ5fxwEdpyNrfOt8O3IEiiT9ptSzHyaYNFxAXCUPHEkY
mtUapRDohvsWCadp9hTWwDIP1d+pZRpbKD1MRYiy5YtQd3lRzQuZuoeTuhpfdU0L
8FAhufKZKIqUhC8FWerdZF9tKbioiu5xGQZyzAKBbrjjCrsBCsNVfnfpaG7rVoua
k4IwNFzYu2l16WaUu5Pd2rfo1sARnYNY4sKKW+x8Cl9azzAW40wadNcWei0DneZh
RS++/sP5p53W9R5nzzR7jn9ruW1PhCTJttxfj8TIsGQGPqt27FLXFWMCqd0G+XHB
UjkZZM4z18Wyn3hiw3P+BGNoaGtwSU2UT6vU6SFQjiC45ipofX4T0ajFFrVO1xne
+Toj2bKFaHNop8t2oyZkUSRy3dsuRRfTsSO5sYhpZ+FI6dGJUVoy96Bh92FlH8fJ
F81vuXieGNcYM4gEr+iQ2r0bo+X8LxQuL23D/iwc9Jgsc3+6jLNvPkyTS59D2h/N
fb1aozJTRXLh6JUyK5UrcBDvvHsysv731JXLtwgHxau/9OjHq/m1eONgiY4pg+u3
3CRb3AKzBGXzQjgiPIV6lkryOHZEDNMpk4tSmA/y1Q0hKvG8S3wf4OtLsCUU8Tdu
zxqOZTA6hQ5qbFSeqDnjYZbf6d8hWpq2USJSaASobeuCfVhFcBdOmw+34HYhkAYZ
DiS0CoE/YfeWvLdqL/zPkHsoblz23Fb1PKAqj0E2lOv5q/Y4Eny69pEmdsZi3HgS
NueKgNBDMQi8Nco8czbUZ+EZILkpwcLGSMrBPI0vMZ2JXg6LZ2cYSn+DXxDrjaSy
JGK86/jK3p6g+b3PQ07/HW6DziL2XZl5rMJeBAFG2uUB0eMNGtNPq78/txsn+krt
urnwg9+rD/yrccZ/uof+yskgSHpTqdqdM5/sIj3ScC6cY9ZhEWFgUzJB6ygwosan
DYgwWpNBDBvqjRZpzP9geKOolvE4wiZwcDMKFTlga3qm7ei+FqBtHHtSb7fC4Yue
gtotmXx7SGY3DZnp5cZsYglIinB/z8cicmZMlfriPsVZKzw3IZuswweT0o57ZlkA
PpkEwOF/bGXvEQSwwRmTPDfZefuH4hpbKUEEIVB/UyyzRB3hykQvHqOElPc72YXP
zhojjBBGBhMFBRMWHnySGgKWs0YPOE2N7Qki8mJBfEwS6KDCAmRIRSDSIEdXPrm8
RBnRl8xkd2j1sDpDhVhwrW8gNFp+jZdadL4iZFVOQX1zQeiWQSIekhZ0AUGkY7tP
vuv8YSl96APwfYuI1zouGfMMEyGbKUE98GIPg4kFPyqDoaRC3s92wKnV/zL+F/6l
eGLJdWR3L+HgcsSUw2yjSsCWpPrzgSafIl4AgGAC+gjTltz6A2QLlq3IGAqLUUst
+fH+/XeuS2cFeploojw9E4DuXAZ/VPtADn+qFLIVj68wXRh1nOVgbzMFvt6pzQRB
giHXwmqHNivlSCd/j0VAMkErzS2HRG8kDYyjq1KC4rMbE7c2EErzf2TO3SrmZDVN
0X45fNrsQ4JYXP6IM7R4yn5BpCR8TfKrfQJuZeiZKbhsJCBlC2BIrSEJ5MlI6nOF
LsxUOZ2eZbEO0R4uNf46Ha9TZ0qV2MxQBCIt2Y1hiAaaCcMYXvLqO7JvXfbKGshg
oNXpnhPZDvyFC0lMOuVTNSsnb+HUPQc58nr6BFlYS1RJmJYjWwghrLZl3CTYx08k
kLXC6GcJPLTPVs/2hLPjBPMRNuYENl5YEtLPLUM+hSWEoaU/km+XBgMXdEZEYqQE
OEHd2LcMBUh4ILW58/f1nCOfmUkE2r5EBYk6I5u7eQKKWHugU/e4lGGlCfZo81tU
Xj/3/QpB3aRspxX0G63ZYpfQY5iZkTNETFjnH/gvu+rzFvZUKqid6Jf0rsoNSxz8
yU4YYWFYiDwZnstQRsteqHCUftDBLduu6WPuLyzLCeoy2EfK8snQJ1bzg+3UWGXX
84nIs+1qQwgWZcYh222r2XC9WaUrWoCKBdOE3RCEy1OvzIkQoneuMwKLBNG9DD0n
lC5llUoA4M7FEM85U2Wjy+4jOkthnvFlfH2j61PjUJEoaZFSQoJGfPNQOAKShv9p
hyWPrqxecOUI06mZeInufRqZB+BDuiMykng+XmLl2L+FAE+tquBfJ8LC4ax6OPC0
RhYBWmISlQXgBiFxlYLm976mFvs9EFZm4DPs7jooa5Mpro3CSJVJFpCV6aLJ5yv7
DBr2dESbJb26zMoMPzUvj40W8yPYC9wowrBHcDFaBs0xXwaoY38Sta9CNnNR2q/Y
XMxK9FGCiNgewpe1GwYj9b5UAd7g7F0ZQy98j3LqSZbN/l0o5mPd6Z5JsHZu94fm
nz3TttfdEXi0Ti5SiHW0y6ihX03+eW0+0w7ZzGCPSBUKeC0InbPY79DS7CmyG5G4
y1ycw0Ar0vgO19JUZeM7jBc0ANsWpc+dalfuNNRCZVqC1rubciyLHpk5xhYrfeCW
3R7UoGmEYZzhxlg4iIhBvSTsc7mVMJqcx7olGXubtDj8vL002YdfUbL//k9/HWk8
8FGMIAOitWPamqDCO1dVRgGMSHIS76nLQ1n82ieCzuUkpZIkA5mukG4qbiTkF8yR
eMWaEobexvfbcEvlnSYmlETFRo1A1Uf7AhjskqX/KBniqJVg27XZtfPPnWkajhbf
lV4gGZmzOWXIDvuLxHBWVTAmWPXb/CvP941vvmm33AafCapS6rodwdRLznAR5i5J
4P54Fax2ktG1xN5KmaEALHLtrq4+LVH5XyDfJHyTcNAB2znGVhQXP7iO5q0dTcN5
JJaypvnhSRFjakS+IHKVBxdCGRk/GLSV4tiVEgTHRk/UGrNMtdY/yubHaI4DpN26
p8yFURaxSxZVXN9qZqpuLdL41S+GfMaa2REZy+Qu9MdN408Wo+Fv9h9s17rmXbNg
c8YmiKp4GS9npbJfoLXhJdNCzjXkFMex1Uh+SpD86yP/7WNkcCuZ0RZAJMOVtMcZ
SLv2t0apoMK1FRoAQm60qw==
`protect END_PROTECTED
