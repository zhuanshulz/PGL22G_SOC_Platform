`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m7+KCdCbZ81TUJsTXFZ3hrIueBmYHAqVKbxy5KTsumG/C95LOELIN7w1JDwnpxxp
OnbQ58WWB8L+1a3mrcx1VTIkmVnkZcVxJEYdkyJ9EBl18EBMNIF5Kbk2VH+5b701
yTeSx2nZWFX6H9rDTejoSj5nlgmDfHBL0XwE4e6g2cH4Abc9WZuYkt3ei7h1Ipj0
wBt87Mf9bmpGz53RCMDRo7LOQQNO4YwO6htUL8ehczF5gpAT5knsu21wIyKhJojm
ZJRk4hBpUcIc48yko9fb9da0Mci4DjpPDBKltE18UzeGaTT9mAQNAQvxIUJUH5Zg
4hmD2SVCtrcFL8XFGNH0bxiM+UZDyxEGMWImTFY/RnCBPQmY/4qMmstf71o+KhIH
S7AS7uAWou4ur4cn2qr8lGtduCBE8POt+0R6raOSU4o7fGR+Pv/Tg+Z81T9LxQZb
IQBzV8z/hRLMHOlI/BRYkI+EUW98IzXf14Biw0lOp1Mb57xVOZqCDkD/jXMDUwWn
Cq/H8VIeQnTlnGSOyjwKSUZMT36cVOQ5vcqysaw4xLPSOyBF7A8Sp3dM1Vu5w8Mo
H/QhGzc5rpVptPinjqzIGiwdCx3YIRPd3tUm+lpebnxWswnzILHTtZI6Ge0maAsT
ZFl4daKgCJnUJO94b0R1pKukm7IC6f56+iu9GEO8RD4g1XuCVscQAOQfB4DRceXx
6sRklyloHEZXjcDDbNzhj1kt3L9+krBphT/v7OJ0gPay1c7NOqnrZckWVxO7Kkv1
t8wxZwPPEyXOjnfalZTnDFuMqDb+RMo0TDi/LD/CF9E6nYf3lgp+/RgfbGgTWB0h
Hn9YjWmc4u707prd7XmdHMDavvimJpsYCaLlpO5/P+o4Xh7+nM3nUq2qt8brfT88
eDXkMT3DhjVU608+x795JQcPAdbpp+aPluAMTUvv3rqAY6Wf7vd0O5RedtIuN5x+
jMizQw04WhguUR0d6xvDS9jqDz43dGs4sWS0im3C/UAm3DBKHXWNfGwsOFVqRjV8
HqVuPsuO4OxGhVYHLlzRipw2sTFgVXHUCeoZeb/Jz/J7vYDEMBZJnFblizSKH6Bp
46oMIuisBBn9UGPjORlCHV//UvQHSphZ4lJsF5T/dth3r755slScg0dee4LM2jZX
OHOzSHkz2j2d75ZY/cjI+dQ9CLUxo0GnSzSqQYbigbLRdKlnjxZk0z39jorknJpP
kpwei/RMdxJE/a5ddSWQAngRRasP3eBPN/sGUfCiNyuLbDvpfs/YpSPxRVT67s1Q
kN/w7KN/zvhoaCeP1TM5hWCcHtSb/FJKtmvDDCIrmtnS63GVWLLWRlFZNmtOd92Y
SvTsRC920X+LwGjff+0v1zEKrfGmHroUlD3EprRzlearGrpsAC5dt2DBmCPh3Ru0
I+yL1b5Jqnd2T5ZIbD+aWd5AZHAKaXrVar1jW9XxbckZYSfcaM+wwSFWnPcBGXZX
DYfI6HvJVbYzLtQNG9IJehn7H0OokVbFr9PJLc22dUAgtzC/zbwJ6GNK/VFBILwT
/rBG1SXceyOWErYXRNBo2f2iUCQ3tx/1gT9MTl+UrqMRCG/vHVNU5Mrrk35mF9yf
KKsCXVbzmkrWMxmg38zkjnomN3jhtn6hgl1J5tGYlRlRofiLMy3mduuJRY7bQJj2
Qwnx/jSvYzqfUJkPa5nMJ9gNPEbS2/E8J+Xp57bLpzP2em1qMCg1i9vxmJnTMX02
OaBCbRxuDgOD4kBR1cD7Zp404jBuKL/diV6fT0/JqqNQdc3GYS75VaMzuIjFTWbr
Dw4L0vavVRyTnbFxvfqDX8g7aBQnEcDLScskXyYWnvSjZZgVNgxgQoA4zVQgSjdS
pvb8NElbB++bb/DN4sEWihwQu/2MRvFwRvdX/HFl/7e9a8gExMXuAv3g00OahaUC
kZD1vH2lqz/IU5nAluT2JvNOtZ8KGMEbWr2WDDsh+BDOWurGeaW1aihOWYcNynSB
ZKoPKPEqmk/y8w0qJXDc945peLDSGGU88/jBwVrFdmZ778HjNZJiP7V8HsUI+xPi
zAY3xECe/ry2wOf6qzpfQBeLudUxq1rk7cDsWt12RHTIthLkXrUCF5kyiFlCnFpO
PfXkniErFjCmKU91lKjllnovjzMzRi46S67p1aVSzPwYCKenTZrGEvwTGCh07RPH
1gUFsutQue25yQLTHbyPUe6MvTopAeg3Jk1ZpEFXvxcWgmZsZQRK+wwh17+tf3jZ
wtxmIZKsNxJVALj95w4XbhXl4aIs/4dRsC98alMuespV8z7DYCH0K0OpmmzY6Ria
OWr8HYe29d2NPM2iheZhchTW5W6Az4f4tEfCoGbV87IttDEGifBaDCyAbFxhKKkS
GUiVwS3IdW5J2OT+Yfe9zBjR3A8j97qEhXdChqDO0dbiLKJLG61taboMM7CstBS3
1vEPyndRL7fc+EkiFnZpCTds4CgJHz00lnUurzVyvJKYRavES+/XLi40mCQwn+kT
Cv0/B6F/JF4OWMoDkMx3h4Lt7lVLyoIth19ENx6DrnJwBmAL/N47mQB2rMtFxSq6
NDzJV5LOt5DidEeAxWzF5oVYCCsO8jwTuKZ++h4ndgalSDwRWP+jA9919aR5ZMK1
wjdsO+vnRlXzQ5/X6XVW40h5b+pFRfB3CJ4jV5UlAZV4iI0GI08vZAlrs8WemISF
T/IoN5qdB7yRACiq+w6rDautMWqvPcOLdiWs9sxjAulm374TKv4SvrlnCCR0qjUA
pMdVc+DfeVwIY+VNGpqCog7WzDpvUouBq+OjHgY54/Kr66QKJAeklicsStsExxBx
nOYtPVSnCyVRrMk5dxW+vrUEaSI2Dy+jh+kagcwa9733yqAmU2TyxqJ6xhC//tkP
ks0hC3ASQem9HuUyvU3BnZ9Cko0TBYJrNAz6gIsVQYisOLzjRVvRsF1y1JTaqucw
Aq55kSzg5ym+N/3RzveB74+gfIEjMWtvWHoyZWQhdXGgrqZ+oFFWEjjzeO9ijshD
dm5stwT2qjQ1coAhuqNgN5BfdBKwP0AiuzpHV4r819jcNwHhFWuDhU0/r940yqVd
xQtlN8U1n+EzeO/+QPCWq+NfhIRBuvlM9cRznzPA3WiExI2h6lQFdOO98LYjBQrU
1k+BA5rECLojawnrdwhhNCJcoZ+c5+ZdN1VBcpWAx0dMpv3/H/qe4ui9+rHAV8WY
SGk6Uzq4TmnRYh8mX6zK4F8U8OUBUAJmLix+o4fiq8FaM1eZRChyAifLAC1a35yG
v/ExIMUvDYvWastNl+gjSGv2ODXcVz2NwrARgLnI2w4pt2gQ/tzlXX3cVkGnsJIB
Me+C2FRmS3Qa9eedSa7cWcCrscC5ZTmyqK9nbdAcTtDfC5+YD8Z3CmunqnAsn9WL
1J8r9eVWwgK3M8jRMApPpuhZxC1DU6wIIwEJE99ymZ9Thl8sao+3FUqGhHkEo5Tt
Qp2ooubvj2BpWWW/r6IROwr1JlvPPkPijLwxmlyBv9F+ffgn99yewMEA4nrKvQi0
3NLzx/8/97QvLmUrRdhKe/nBun/fyipUzqOoP6Jf2uQhLqpDLyVzE2fI7fX3CgFj
1UEDWJsSl41e/8vHllIn5RaLMaBa5Ll2OzTLPU+HvUQulhuLggGXWPxJOZHb7ZnY
oQxmwzRDSefkRs/8yn84XXTMzz5BVNX9Gu7YHgzjOq8+uXYyUtWdiNfckrUMiTm6
+3+KrGPm+GtgP+/ugX8I6H1S9aI18Vq/8x3l2slsc1ETd1xqPmyKgZdbTL9smpNg
M6pdrt0MJ2AYxUnKUi5+7GkvZHfhtMV0wiYspHRmw7IL6XmDO7RAxV+GBx8EUh/J
RuyjhmNbFgVfqsB5MaZuSw5OTbvwjUtKabvksJ6JHi8fnGtN1jv81roHu+RL0XLu
YdHuST53k0aozCd6GY1XNw351111Xk4Pyy6eAzCjKK8P0oNojELJUAVFyuMZuXob
C0Q+v10U6uWWBcqtt7wK8jNLUKAKo9jeotymrnAbrDYGtitkV7AEqxvuMFWe1/uZ
EboFxl7/sdSSgKbbnxtPEyQ27RD3SVrVKaOp+sIY+Hg96rqvTbfAEgfWyIqkRANq
IZTqYxWaPFV9sF+HJh6paV6YJUfoiUH6QEXwnz3DP8UFb4W5cma0ivXFBN8kcDnf
P6VGnSwZnoBf7Mk6kC2hWEs/zZkHiKGZvJNtNkL8AnKH5JdfSDNPmSLpVG5HjtOS
vvSqcbO9F4KhyuUGjm4uDvqojakH71H1frTIG9T7uJNOktTxYcG9Lt5gFeL0Yd7/
UrIZ6vuP8+BKk82BclloFPvVAlcTJfetXZuTqC5APfF8D3OtnVJsGskU8rhcF3Hw
PsF/PMrayZ5aFtp2g+QD5aQw/QrajT+6vc3muDAI0v2cuWg61MvKygRrdb2k8sqr
kKRNAeuxDYxtbdjLzeQcNBvfkjsVFefy2Uefu57BFpFiXljSnzcE2RD3rncTCcsY
sIPyc32RsfhOX5nVFAbqwlUrzuEON3lS8pOhGS6+ibPL/34IPHfvVI09jrRSdvM2
mveNbS88BCGdF7inxRnurroFBUcRntIp804Patdr3F84E7NgJ4hZR3O+PYrKzTXu
ojARu8+/WL4HtBSnEPtHxSlIF67EhdS7fIZBMsc0s7ukLmO3Y2e2VymSUf2d0rOA
`protect END_PROTECTED
