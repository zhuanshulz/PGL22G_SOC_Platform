`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/JYWn96PGF/7sYCKOx+O9P7x46WmDtsN/8bAj+/bzXF60TTRshcF3BUolr9KKnV/
FqQiwYpPy3haRaJ/thPChAPBM7gsK4VTwNRYi1NW8dGl/Stf6TrGSfViXY+sd5Za
zlsvy3iAzhzt48iEafkToYXR3fM7SsLbf8uPsA0j+TTz+TOg/2ua52fL8Te1a7T1
Ff8t4YTEId28F56GCpL1D4+yoy26tFEJY9/vXRpUkP9QC6xQsxpRz6mvfbC2JVOX
r6B+3KFNJ09SKGask9OULdCW1yH6WPejW5h90mTbOiE2udWpFSg6D9MzWwSemQOA
vrKjpWVsVoLMMNk6FhCu2q64U6zE/sUQeXV+4mJa/zEStYnIwXBwAiqRGUUTRcfL
/8f+lcNJBRfGDDrslldpIyjOMeeGJ1ey75MzETlTyo/8/a+ihJZ2saw2Uooa0ps0
QkQ2ZJt+ZUzb8r4WcRbcoJ2wnjbIPVfpFz/TgBgAY/Vixy4vN5F9QfrmPcdXat1A
WViMPTvCE4X1peLJ7Lv5iTdpvSke7uwlJarXMEQP+WSXWkticHcM052jrCNAxvxg
FSZKR3JSI88CY9/3SwA3PGqI3t06qdAckoKF1TDtb93aeXuH7PXnOr4KYtOlXsdg
YCENY2VwPSLaehphFcjOZOHSS/ZXnuID9PaJbHXkbRwR6f9ZJVOWc/Q2SECspErA
QCsoTC17YqsSaIfys2/IGK7LgYoBqMZ2YH6pQvOdCiM=
`protect END_PROTECTED
