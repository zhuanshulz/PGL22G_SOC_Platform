`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
16fPyXoRItXQ87z7Grb5G/YFzh931kyNEGl9Iu3fdXzqI734LXk3bRrM0ICIF2pX
YHNDblt1AWYQ1vSHynY6FN2u45fU6mxhqddmdADU+iT9dgGSPcasEdic1Om1DQ3U
FqDu5pW5/0o5ey/VJheD7Zeo4SD3v1gdDJg9WXM29sv3egMqXk6vSsdCwnOzuMy6
u8UZLPGL01f8dP9v1Z1fTMwcxTz3Ia1Hv0PBIknIIFz71+FUJYTJuoqMytG/eP4L
WPaSJal6cgPVLI+lo8Uwbuo5oHR36wSP7v95m4VOwFgtkC4hHf6at1/w8KkcUUce
u39lHABoqoNjs4N8PFlOvJlSsRGkspq+0e5GiQQ2k9hCBDDX2mlTA/1RPqwHYrcz
8av6yABUvNoylPyCvWVMd/s9etunBtDBIapGS3oCkhZ1QML1E56H9cOH9NgnKDSn
pKbF7zsgpT63AwjROqILuCwjtAo+T0yYEa7KBXnWZQqL5IBW+x/9VmIh8elhXBPW
jxh/quHpD8TOiU2K7kal2SkUttwjsODsWaWlkak1pIcKHtfc+6v4eiZMXOT5mkg5
EZOfdu0KbV5wnN8DRbVlhurZUXXcNbRVE+CmLj282qJ/aILQDFu+EZixgKqgKKgx
9ZZrs8yExY93GRFT2tjs9y0KGesWvn+By3mAfSgFYwmoarrlrokclUyMS+5PVlQx
`protect END_PROTECTED
