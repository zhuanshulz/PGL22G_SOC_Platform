`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MW2wjUjRRxZjebNA+XX+gTOxTMhAwvRJVk7/5OeAS7m+bzQ4TgHGb4BfSvR5E+YG
OxA6MTtdx5sIRoXaIwi54DSb6mOCxUuQTkryOCUnWO5PLZIvOMGBHI8D1jXBkpb+
fAXN84BB3/kbons1ne2x04ZYsYCVfT69lQznuWysLekYTMJzOa5Y0qXArAQj1iKa
dPzu8cDihApKHVSkYG87hwzeV/iZ3JFTPBNXEkrjbgO1HGT65Ys0yUGiOEcV3UjB
WuwirWu9MV+WqkvzG5Yu9Q==
`protect END_PROTECTED
