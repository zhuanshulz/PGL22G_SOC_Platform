`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L4dU7CYbvlYTT4vuMkuBqJNq1E8V+ynrRn7PAOMO79qa1ZW7TMllS7xv4+FCsQwI
zpGXF1CTFHI7YXYZ/UhDHcivX6Lqr/IstpeUQCSnIWGNK3ZmEA+yzpFx54Cog32H
vlgoBjknhTa9hb8bj2mi/deKMQAVLIORNIzOd3PYa5wvX5Za67TWC1Pog3cMlqtA
iKftsLO7Gz2UPa/YQI9A7VbjfuIki+NwRi6g+NH1pHrIqFPdnVORv/kIKQDvFVvW
R3t/Hp/e6CYLjxVzbmh4UpLE4l/7uv1xbsPaanz4L4vNnULdDYTwMK6DTVtQ9Uf6
KFwL57qqUSzByO5xXQKYug8JjUrUAoFj6qV1cEwBKJ2FPCbaJ9dgqinU9MHiv6fN
G4DrblLloVMANL8sODlSozCQIEA0MO7Ynn9t1nAXHu2p/gl+YBT3xQnVbzCKN2fv
Cqz8wHS2pqPWUTeITc1nA8amleM0yGsAtFU5IPGLUFLd+Fa6MnB1SDOb3QaC5al8
BO+GeExJwjRwcHswGq7GBfWPX+wMOJIdZhyePEgjS+XPwY4TrGAY9Yr879zn+nAg
tO0RRYPXpU/d6DOpn4jOWWZd8hh3I0JutjPqAtfXumeqEIZODkVygQc5dkGoZiNU
`protect END_PROTECTED
