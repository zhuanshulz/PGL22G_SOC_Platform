`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UpF4+LiVfJU2rIVSOdjmI9YEBMBLRofl4Jf40scfpMulsCPokeciYB/xuXqotrDr
T0V2u/U2MK6xrnWoK+WvyIIUns0dTa6Ci5+PEGceOnvwZteRTfGIQPt/yB3KdqEB
52N2jOUKyfZ1tmTk2MbljnGcKRRWO6o14lyjizjclrc/z6ftdl0Ayb1dpOa0kXw1
NzL/kjLClMpaN2N+ssEnk5zdh6q32YM2dKs2LapcAXBavuLBLqKi9Ea1ksLz26ih
zCcZJk+6RcNaFXkCI693lwYTrOzOIwsSpNdA6Pqf30NFGxMwZ/UALG4hLPnhBK+I
4nsfe50FM7GKTBxYvX8j421xx/DGBG54JHe/yX0NPrJ+MNzyTRalbPs+iovVUVdo
vvpRR/KIPm4Qo0LBxQMdR02SjL5YyRAlQA6KwW1EsGA1UQbxcBiow2/zccbqlx4/
YKtgX10CTw8H1I8EpaK65f3DlLmkTAAABXZLdYfe6WzEC+aWZ8wXfyaWejieIwE0
hVGH6YIwZzf9WawOcNWfYw==
`protect END_PROTECTED
