`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1xn3d7lR8PtbweRFGDkirx2JAuQo//uOwVdQINkv9103PcNh2mjuFHxXa5nVN5UT
ANnkPOhRK9/bogIqq4LelH/SO5FzZ3c1kBrlNv+4SNlbiy0R3JZUzbv6UiCmIgTn
emNXIKm121elsqKkQZEVv97z0ZjIOXNOmKEKODNtxq++bmpaVmwgDRwVUrtK0tDi
bUB2HS5lCN3RrY0O7XSI9vUTSEoqNZUHFBAsXO5g52sb3Lvxen/c6LsQL3RzzT6E
Kxdrch7GyO0eX6mYUuruj6eDqhzn43ya/S092MgYX6XHlhh1AyArxTDa59QDVWdS
dJIaLOLF/9b10aWbE7FXNQnSUAuHpsZt2ifd7oN5osyT7hzEqiVaUzli/CJVBT7K
joRunYXhv6QspMzX3VASqZFzjQN8YaXMjvHO9SHAzqzHY15NjTRGcSfhUGN8XT++
kVzul9r7esI5DwX8EVSVBLObSsnCw2/fB/2JmSeSUeSSOGtAx22tkMskpoQgVope
aUTT4rStuHXcJFk34FiOQB52Fj8TCaCxQASkULgoM6qTb1rVfA9nQfLsdasIyqYH
Crw9zxK+I/hvYF8173ZhPtLbiyN9b7Q0xfSvGkesl7hFDhBsws1bZzfXEc1Qihb7
/mU27R/eaO3DDEC28hQgP17vYH5/gT5izgZB+xmCAG9t5nTFZ6ay/QjH5INkJZH4
i2GeFM8cyqfaodOS78lXrR66expsnNnv84SGhgyKzxmK9xw/SVpDdDoNvS/tPYxZ
gwJdwKW9MqE8fzcwoBi7U+Qy4lrSK9M5UV+1f9oLKGjkJbcWcbL1ltGA8SHG+6VG
PdEfJksOZmvT5Dx7yVA+JIvoNUqEV0NQbYUiHCB42qKEZR7rg7enAbsRMrBC6kWT
VEz4gsB6HIzsYEXHhsTB37XPWKW4A2Gdj+TN7pyvItnAZZY0hB9EpS1YskwJCDuH
RwAIFSEpqNkU8KLl2PON/mMXQf0KLXTsqpvqTuO0wjJEdFadcgyD4f/fKlVkJK0w
WrIEbBXy+XVrFFdE/1rVd4MjCSJ955jyT8VH/ng6sklxJpHtibAhGTR5vR9k1jLf
7dJvJFvu93d7gvl1XoU2mluKMP0ejOOCu8oIzt6E2vPYm2o4OUDbQO4MNvDjpzlH
Gk2WCWI2aljC7hOegc8MD2gUJHRWiWFSA9ReuTUCDpqJuq0u0lkXwaG45nAqmfra
oSItsbdkphjMNQAo3m6cFDbknFSgAKv9O3s1+JHx+leRBgkI33gDX7zgvb+KFqGM
jsiaO9F3YnbsGutLJZYdeixoH+IAcZ/lwGCOQNcBOQFOeZNKfRpPGZBuVdJLC1Hf
SxMk0K8ZrtwE2tCOn7mkUA==
`protect END_PROTECTED
