`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hOBaU5ve+TWhBN1TRT90KuUgRWbD4F/IxHi1te7aFI2g+ncZuGhom4FcKwWBvRKW
mWcElMzmDUtZcvIi1EYedx0iWEhy/EvuEiit/2L3mXow9a7VVkAJHEofRnmFjwnS
HvFCvcAH0no4fKVWM3nFn17KZtVMM/FeOHmpTKUUIpEFHxMqaj/ek/2k+ZHOW8Fv
onrsIuZ6O50xKLRr1etbRr76Tpa8gJpvW6BG4POQMQLzOMuFpGuNfwbHrvKIywRF
uCSgspevaRWprhe7ozp3NkmsuxywetbkBaW8uUMl+n9EUAHK0Igk7GBU4v15Hu73
eevwP+T4v3KzHkh+XUNEZmiepR+2QrDiwsvinpDZpRjNbQvnwIrJXPNKvdN3Mn6p
5Nw9OBI+tAiot3BkVdC8lNZHMaghzDmkV6bQKnJWNYKv7+SKeZi8EoFvBWNZKOCL
taAXOUQ0Eo/jbS15EypoP3RFsq5JpyxOFqfoAl8gFbfZBHPDJYJunu1ddOQc4S4v
2DD6Ojp+mk15wtROqGHf7hUE1bnFqTqbl1tfrCsjne/vZhWt0+T69d1HjNUhiIIz
tUaBJH3uI3462lx7nzMSCfaEvGq5yt4QWYpbeFD+9bVKIXFdsbcDsSLTle6FFipn
S8/ytWRynD7Ol3dy1ZBsRTRI4LxLW8IhA2vBfG4/+QGoASfs3cEnp+kDB+MQfBhl
wLadhP3h5HyF1ROHAZuuQAVX+x7UA0zuHXO7DyQ0ctyQWFIpaX1C3wHfrqOCTurq
0GNFxKzt9HG4tczYLMWQv2vBfKkofKkMHgOWubcLMtLdsbaSPgOME0JLzDjpwNra
MS8z3rPcB2jPGbvNeMi5coQ0ypHXufkVVbjcBu3pOQR+XozjLa6SjOYDnJ4g06IA
0JIvmZuL0XHgKiWlpsiBfBYNhsF6LmMJfun02SOTffmZxObSKG4QdfrJ5LOajxp5
HwhAURfKA1lvInwlCKg4+0qsIOz9H6ZcCX8ULyJd6aU/rUWCA7QXTymoD03q6ihb
fSbCQTt9+D1I0DmMuprjbAAoYTtNAGH8wZrwMYtnkBqFFroRGoMvhKgwzbjI5WsY
GPAM3eO3gzQXXii2VgyXq7RqEvLphqYjzpUB6LxgIG/e+4SwfILBhSuJSRc0yLwb
Ko4GY9PenvceBWJJ1tlqEqj3tvu0lKYRHubezP9QV+UL7knZcY8+VIFwffrWOG9i
eQVxgEipJFo3wELmxeabHDqVQEYPKL4zZWPRoyM3kM7XzTw/+LtzxOBJsc4by/Q6
6Ru4gJmkDfElR8n/58kUhSt7QROWiDOXJIPromzaL2SMY5WFrhQ60qxiwD/xfgsR
7j5DOvxjwWYNnSv6CDAtNYHEyg9xVlAfg1exFXB05zWgN675gEU8Jp+d6q6Os/+R
pW3+Mg9V2tkAlTmfWKH+ydqeFmsYInRA5wuXJ6qV0HHxiDbNuIyk1NgWgf/q/2Fo
pSf49kSQ2xwltrmZn0PNWsptlsLT25dpU6YiaAqGcLLV/PgnWZtej7wMzcHyqEhf
LTsTNxpOpiKg3p9CClbXCnH7/jCwEjFf751RJXM8Ec6Whz/6Cum4OdavzBJM2J5W
T3wmc+sN+e1G7DvKfZRcgJlyPr625RadTCuJymIzTHfFFd64NNm+UxjdxhNpJi0c
boXeicn8sOaPyOqXIkX2ibuhxyL9sGDnbo3gk7FJqryb3rPv4iSm9qCgbPMsxbYA
WLnFH4fhZSeyHp9uVPVaejOdVN7nUcMgkpI02bX58BT219HDHATfcKcKnpx4LIBI
FkL7Hv7nLCpCPaeAIZmDxW3mwpegMyEsU5AI1oslIsJmqrxQ+qvV7lxhRRk/GnVF
UI3tufQNwDDHFWI9CR+M9/Uo4VTUbNl8rzEchaFBz3ssWKZw4p0LqBdGHmRpXToo
3gPgqjiyqCrLqbQ6ZDUqmDflQez6evzS89zCdDIh/hCvdK2z8QxnnIvirWfIXBUU
8h3bbY+cZ+KrGqhElRTqZR+dHdmhCWjtNrPkbR43BbYZb5+AuXtl4qDh0xY8bpz5
dT8QN/WI6cy6SiCKkatJ9iyPHv5z/3LduibS5HuqGAHdqtEEFJzj/JY7AX0AfQH1
UsHsi9+hDJygSufUnmmhQM4g65fbmLW6OdQYbVhp2vb6x+ujc3H3doW/WAuMmEmo
ySjOeYYRIAjZHq1Bdb2+b6dPbVK74zTl6tHTYLa6B6FQR5Xq4DVbd4fY2y2Hfl2z
omemFhp1Z0aolsMUQlXjSKl/w0fkFWzTy/s4sTDvl8Lr9hpJ2d5gRkOV48/QDFIV
o2pBLaoj7P4nkmHX5v0Y26PMQMTsEvDwQbsoU17jYzYTvDYAaI37+NbHuxVykvfi
TV0UuSZNrDT0T1b6syk9SgzptmKJNFXkTzh/YMVDdPImSrGSTPeGHqGKH/FnN/Mu
qaoooxMgbUHI2XIhqlr926TtmohYJiX2EkJx+IkMT874TOoDa514CrvsquBoKfr9
Oaf9Jaov80jPzNMlsyvxgIByRtLyjEKmv0rmUJZz/tVHzXJX9e+NjP2xieSaC+IH
Brq90/xAf1wxY4UKKZ1K6NairUX1+9vr6rJXZognMVRCvElWXdKQzchGvhg7XqOI
`protect END_PROTECTED
