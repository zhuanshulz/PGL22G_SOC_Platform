`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yMS+pwUgPkRG6Ab/BTmPhS8GJ4yxlhWg1mZUk5/08qdaVSz1vl81oBwdr4A4mpLm
gq+M66Mi2BSa7sov54K/VsgrPTH9KPQy4R9kn0wejCnGxoMZauHu+eyKSBR2i6mF
h4K2nbkwlaEgfdQzTxShFFhwg2e3LrPzy/ZxHT+oeVALU41M426GUojxfgU+9SLg
CpPnvbKFhXnCjBXqcDihm1ufgPdwDqpPkeU834DgX60shV+kGwKAINroP8UZgD+E
hpFKDaFqH34mts6mAd9Wi927qtgoPoN+zX7jQLAlW/8kthD79hGmlUdCNiaePPa5
Zm/BMfzL9imI1a1HFPl0G4T7HlZGS+OYW7t4avwPRj1zFFdPN9q2gqPvHqh+pIvB
2PKs/XiKJi5Z3ILqlWs7jrzrS3Ws3qsHQihH8VfSf9zaD839s4m20wtfcntQzpUS
9PQnwht+6ZE7hjdbcTl5RM1TdNVVA0oBqz2PUd71dFdkPCWjqbp9iSm4tHNsIjuJ
sVcv+PXzQbA2hgjIQnId3FuUjKF2Fqpu2+KTUWPqCII=
`protect END_PROTECTED
