`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fXPq3jNrBybR7Jqx42G6Qy0l4XwjOXnalQ63aKG36Q1khmkH8FPeCmstQYO/SZdk
/wx71YNY9XpDSjC29Jbu9ErMhlKMqz1aLsZCZOx+FRGLK/tZTiJaUeS+z1domx6u
Ye2DjKTDHbRpnRYyoy14O+7YxuNgTdGOhwVGiBCoexEbtbutYvz/D2FR6m/oin7C
2Jbjz8LEvRYF30KpThZpTrqiaYTUBxy+k5Z63YgccH6yIOvjH20uLGR0OMmJRq3z
oOc6T/mnAEVdBixQSt63eHOCBQn34swoOAbzYreqgRhXm9bn6oitwYwkmwenlqQg
D92MltOQmG/2SWLoQTzNBqkhl5oqwJC8t6vmKH1Pf4NIBmbw9zZWq0TDNcDG72tO
fDuyn2h1rfkQrCd712EoDApvNpt7q/2d13fs/ZoNCUHO6hpROCKuNdn0VI6cGyl2
UmbC7iyZUGmcNcJPiLBTc/B7MisJEe9q85fBK7niFlM+hkhChVpVbef3Pm9QUHIQ
Df4z/u/nygtmTswvuASX7PVuiizH6gXcaosIlWI5236KNdwMJUIh8XSIQaas6ukb
oIIEf+gu4XRLHQcr942Rqw==
`protect END_PROTECTED
