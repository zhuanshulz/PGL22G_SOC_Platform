`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5VhZX/pOkvxGwMT4W8dsmNPEbDk9/XbztTEnwm71qGe3xkSwjCjODTHtR1zECpYX
phnX8NEf6Xe5DLCklIj2xY+VHgJUEey0yegmFFVb9uv9EO/D3Gakqz4nEjSczBcC
kyOcV7Vq7ajmDU21W5vHktgca0Rm1Wx3w5RK2Tc2Q0Eo0L2rfLjsicBzDVkv9XRX
SbsRTS2ascnwdPRBGeMTcdCQUolDXGevvHP8LVdPEQp+AEMSKsHe0B/QX7yynS8P
/FhLjL/uHKGOmgrO8Vl29Ck1WJvTZk1NfLq4ocQ/4O/JU7AWFRMDiffUzb+XxAIq
Xys1r4/l1ZF9G2bP5DPg5PTu1AJfxM+VnlOYufUS0pWM1VCvIk8zafh3fY/BvUvG
0IYbItz1LJpy6iz9UkULcvQmaAcfN8IL/Dj3TIFd2pvIgomCcFoXz/xJV1aBB2Od
yrYh/PnZ2NHdn139vQQDGoerOiEEPGVbQpiA2dh6Tj44n1uEGJE73ku7lQWdnCxw
HN290GYg4Nrk2lEPaFE0IfcwbyQzbb7CSD9YY8vLSR+mViEyD/NJgQieT7AkGNEm
dsIFhlJXAd8OAG/5cz+Ad/FIa2nQ8q9WzZjOOodeYzuoMgq2I4TEC+kpvG9S4xmY
1dBg3yYf/TUj2UqtS1J9tbIoFsW1yTAylwp0Kai55DWWBqkKC4P5qImInxF3vbc4
DudoWa1NxpVSHUYzJjME71LBn2xcM+L260M4JdsHgQ+CvgJjtFEzLON42guEArym
n7e+7Ii5fLBhw75G1YyOj2sjpmIrdxPC+Wg1v8kbTj+DL+KHlVgtqLjmwXLvEbs3
n9metse2UE/pqbjYcQLLv9B2AKUZFG2w4fEl4jG2rVjcTzGWt6gbQ/MtyQ5CLYzj
CPLBZoW7xW4QjKXMXgKKPL1V33UTWENbUZAQa9pVHImq2CHc5b9XYavfnJ7Y5Giy
TksVh0bWP00J3UPpHfv0Taxj5yqSe48B6sfGkpL7pvKdex6W8cDUNA1x/zYmgMUO
XYqW7eWdUNwnZkCdKog1+OWRL4Vb2y9Os3BigKpRV5+4LSc5ifJ6YzHHeSDOaaLC
I9v9lOaq0RqXqh182L0rLsRWadQORZX18p68I4vs2g6Ir6nv6hOiCWw1nf5RUuyv
Jjv/7aNuotJD6ixJyxacxEj8vmWEv/tlsojTC4kQXW1rHC7dYemZF8jIB9tig/3f
MWaRXwPwkp/yWB1ItLdBXTXqH/+f6fpesq9we3oLni53ohM14URaCkNkcVD7zFKR
D/e/evuDKgJ1m8r+YBZCq9ltO5oi52XE9i4ijcoj4ECnGatc7GUTVFUVUYSyOG12
14aenmJvTQZ6bkTswFzPhQeDF+jUke1OxkvmTgDDl0Cxmb0WrRIcbX2BXeATaIyW
tuaQIMtrAPlVsQ0TS3S5qMxAnsrK+seeMrGXFzjiZlctP7dGQemjARQaTuuwfUfp
diBYLf247GsSx3AccRT8E3AfJr1qnVKQWYKH2DhWnbA4RBeL533g0NBQ4knrNpMs
wuKe7p7KwBdTa3rr96EQf34SX7cZ1jJ3j4RYM4Bzr1Tq7hagfOMjOBoW9O/b4x6X
WmzjD9IVuj/t2T3NzZZAaTojG/GVkxfYiieSNxfo1pHqsxAizHFUaiB9NQGhQRjt
8aJVsXM6bqvwBST9km0yOFiMdaAeKDFla1DpL2rBTFUD9G4ptJFtU4HcMHK2g5ZI
AeeS+ltHEU9aB7HOwHiXZwrF8AiOkS8NzjMYC7TcD6JdUa3rW05WOuvy0Cdk9zBu
BU0UeiinIGs/5QUdfpZEWusBrUG55i9D33t8frCKHI1VGnTLNvKjl4Zak7eETEqm
5BTDfa39xsAhd3c5c11tjY0gXZzm6VtM/jTu8d/Of22t1hjPOGOkAdoZt3c1Ek1/
rPPsopcMGOLUW3KAn7+V98oRlfBvgQwxMQAM9Qq78HdVX78poS+k2x0QhHu07Xlz
cdYrnZw7JcorzI8Pr1ujonA6WvO9vXrzpxuPUFCGAHsMbuzNT7DoaWCI2aCqFzPw
s7+dqJu4o5xsnclBruTG3cfjQobM9Y8BQ+kBoJMfqax6gySFQX/wXpgrZgvYXwlG
aff5CErRlxKMmtS4AH6LPAfn6hLuihwMIrZm731vLVuG75fc077XlI2j9cegKg0v
27q1uEcNyGV3w1N0pgJ6UGVDBhew3FgPHg9KYrsQUHp4Jk3d6lVcRyWgvvrsRwWk
HZXjg5IDPiPpPKjIdL+J1gJaPoC88YFE86+xGTjUgpIpldLEJBVluvVVCk40NW6r
kgSwcJcGPDxnl7RAKJu2E2z2Oe3rDQZI55hm7T0Vwz8aRajSXj0HIUvXe37k4f4p
NbEMvPwJcQ6vTUrFdrap3tjwdyvHbGKepZWxnWe7riSz+i8ANXJ2gggtDshPPXf7
kKqePrlk+K2JqnRNvpRD5EGqe0aWk/8pkZrIQC9SbmLgIrASr6C8p6eANJc7hWC8
F+A6Gud9B+wQRixPgH4Euvd7vz20f0ss8XNDj9gUbGKA17TYmcpnIAVzlzDzrjXr
SjBuHR1Imd+4t54F5yjc9sdE5do/n6MD7EJdbOFk47X+oV48B9+djS594Ee4YFxb
R/bv9kRj4fpFuwijEYW87WOGkzhta8uYvopb+DKKiKZdfRqBW+3we08Nnrbwk42d
EGNsw20x3xlLdOm4D5t5ZAg6tuAQqUt9FkhWZV0JDIX8HmDxxWCgAroQ/YEyk9iG
a0wNHjSDaY/vu1yVhozVnhG8AXSZ09LYhO6OrY2guoMJ8YHQCaLN/EGOnroVSKLt
chIR/uvIoKb5a5InQPA9l1VlJt5v4ks5fdPuN+Ch8gdDNn8+u7nZM7cFji4O3WYF
sey9nURjpkZCvlRzR9tVmtvNr7Kgkg3i+QjqGl/4Z+Yy/ecynJq4lL14ou5Qi3ME
skz9+25f1Vz+nGM/5oOWYQc42pIABY820rpAbzFeCCDGhIXykjlu902ZEZtL463T
jMaYDpRRU/POyQYekvws1+mEjKO0PU8qQSvrm95E5ZZGIEEtnweaSMAeJlkiLTvL
LTA6kQVIjHtv2Q60o/ZC2Hkm9QXjCTQEam2IrHAv3cyWOKzn9qevviO0xVfujjKJ
KtAeJAXuUGDKElI7MUKGQep/BQloF9DLYtdU4tcqMHmaX+bAFIl9GiagO8/dG5tN
BwpFS8y0Kbx87X+ok8wwz6PcdW3H27b1c91LeK42iBbdZSwMSwCFeM3+WkF/qaWi
uO2K9MunZZV9diSKMJglfR1cNDtkkaUbD1y/Ev1jsVHMNrDkLLdSF9hCGVpt70Pq
OVJf62Aoq70VCVhGwoFIBiRh/R7Rj2DXKSdBPShj6JMLTp9mhS6n20Er6vkk6Jzd
0v6bXGrHbsDpNh4Ah8fPOuaJe4IBwSeoPauzMNNc4qVrB09ntd0wxXXLPfR8y07O
AuwIQS2oAneHSKNngOAI+7satTKrxtITn9sLMOEAnQi9zZOvJCLIyvysSPnNpdHe
pJYs2Tpg8ArBhLDkn+g4NpFia1/0sh59iLuYIfYJ4KMwDKVsg3ThVkhZcBlKKUay
DPMZD4grL6fudYPlQMUHwYSj6GkTfFXUiv24OX3TEuY=
`protect END_PROTECTED
