`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R6+Wo+GNA4nw3M2goelnCxySz4+q6E4Ldd2HL2UQlnd514wLGnd/2st8JBsezRGl
yGLShrrMZZJ/KSNVAatVaEAllYVEqV/chuiormD0OF7F15DUEMPeJDXdf81ZW4zI
lN1g/Zt71JrfcbkWB3uCuXxscofAPWyl2P43ZZCq5BZWe7e09A2NvzNVO3tREOYm
WnvDVRUWKVs9udbRQgwuj1l4cPFPkXp70sj+azXsHP3x06NmM7gsm2g9wwNCYjFX
TopQimw38CORP4blEX/zs6MZDQsP7gxWrQ4SvybppcW754W4d/CRS6of4ULs28tw
ALnvhL3V9ksBejAbC0ESEQpT4x+mdsFEAHSLM4CtAqMNxJQKhHy/dA9jgguE7pP1
QvUKUAzEGneYIckLLTMq0pP6oVEBBEXgxyt+keTcblmRfaPWPy0byKMPVrYcXpQ6
5uhGdX3Vo0UBuS2RZfXmRC0k6WoTh0eFMV5M+BjEsBRe/nF5gsGXoGx3UAOYwDxz
fsHHFLiImtKhRtKXnFt3qWFVLrG8BZCp8adX/KwaJs1wDEZPEh6cEnyahThhHNyj
pm6bMiPWNUZVkzb+dlovDuzJ3hIhYTx6kpzhwHiyVXxKpheqZZOf2fggiHWju4Rs
HAjKcl7bH85C6axKh+QtzsQ+gypNnpg5o4NNLdayoIqHsVUwlKUfAeoS0g7C2zS8
GECrBEMsXhBMx5qDTeVSkJNwsGo9jANkjhvu7w5fC+pDX0qWXwhkwfe1OTbLioMa
cSYyI+2wr9v6WdyuD4s2J+07sxLZdew+8rRldvBd9ZN96GQCk2zbioP02UsDxxRy
YC+tYdM0IPngcBG0opIrn0tZvwJ3/17lRcIBRra9ogyG5f5c7w+Bi9bNMCe0PRTL
UET9UUw/dPKgVkbHJhxRVJBsnUwohMYYP+KA4/mk3b7z9Vy7JlmxziZXNMrOy4tO
aJpVOVVCTrDrrRZc43lRr2x1AJlqNQPJ97OXXDdjTP8=
`protect END_PROTECTED
