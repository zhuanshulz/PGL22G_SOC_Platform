library verilog;
use verilog.vl_types.all;
entity V_HSSTHP_LANE is
    generic(
        PCS_DYN_DLY_SEL_RX: string  := "FALSE";
        PCS_PMA_RCLK_POLINV: string  := "PMA_RCLK";
        PCS_PCS_RCLK_SEL: string  := "RCLK";
        PCS_GEAR_RCLK_SEL: string  := "RCLK";
        PCS_RCLK2FABRIC_SEL: string  := "HARD_1";
        PCS_SCAN_INTERVAL_RX: string  := "4_CLOCKS";
        PCS_BRIDGE_RCLK_SEL: string  := "RCLK";
        PCS_RCLK_POLINV : string  := "RCLK";
        PCS_TO_FABRIC_CLK_SEL: string  := "PMA_RCLK";
        PCS_CLK2ALIGNER_SEL: string  := "TO_FABRIC_CLK";
        PCS_TO_FABRIC_CLK_DIV_EN: string  := "FALSE";
        PCS_AUTO_NEAR_LOOP_EN: string  := "FALSE";
        PCS_PCS_RCLK_EN : string  := "FALSE";
        PCS_BRIDGE_PCS_RCLK_EN_SEL: string  := "HARD_1";
        PCS_BRIDGE_RCLK_EN_SEL: string  := "HARD_0";
        PCS_GEAR_RCLK_EN_SEL: string  := "HARD_0";
        PCS_NEGEDGE_EN_RX: string  := "FALSE";
        PCS_PCS_RX_RSTN : string  := "FALSE";
        PCS_BRIDGE_PCS_RSTN: string  := "FALSE";
        PCS_TO_FABRIC_RST_EN: string  := "FALSE";
        PCS_BYPASS_GEAR_RRSTN: string  := "FALSE";
        PCS_BYPASS_BRIDGE_RRSTN: string  := "FALSE";
        PCS_ALIGNER_EN_RX: string  := "FALSE";
        PCS_RX_SLAVE    : string  := "MASTER";
        PCS_RX_CA       : integer := 0;
        PCS_SUM_THRESHOLD_RX: integer := 0;
        PCS_AVG_CYCLES_RX: integer := 0;
        PCS_REG_PMA_RX2TX_PLOOP_EN: string  := "FALSE";
        PCS_REG_PMA_RX2TX_PLOOP_FIFOEN: string  := "FALSE";
        PCS_STEP_SIZE_RX: integer := 0;
        PCS_REV_CNT_LIMIT_RX: integer := 0;
        PCS_FILTER_CNT_SIZE_RX: integer := 0;
        PCS_DLY_ADJUST_SIZE_RX_3_0: integer := 0;
        PCS_DLY_REC_SIZE_RX: integer := 0;
        PCS_ALIGN_THRD_RX: integer := 0;
        PCS_DLY_ADJUST_SIZE_RX_4: integer := 0;
        PCS_CFG_DEC_TYPE_EN: string  := "FALSE";
        PCS_RXBRIDGE_GEAR_SEL: string  := "FALSE";
        PCS_GE_AUTO_EN  : string  := "FALSE";
        PCS_RXBRG_FULL_CHK_EN: string  := "FALSE";
        PCS_RXBRG_EMPTY_CHK_EN: string  := "FALSE";
        PCS_IFG_EN      : string  := "FALSE";
        PCS_FLP_FULL_CHK_EN: string  := "FALSE";
        PCS_FLP_EMPTY_CHK_EN: string  := "FALSE";
        PCS_RX_POLARITY_INV: string  := "DELAY";
        PCS_FARLP_PWR_REDUCTION: string  := "FALSE";
        PCS_RXPRBS_PWR_REDUCTION: string  := "NORMAL";
        PCS_WDALIGN_PWR_REDUCTION: string  := "NORMAL";
        PCS_RXDEC_PWR_REDUCTION: string  := "NORMAL";
        PCS_RXBRG_PWR_REDUCTION: string  := "NORMAL";
        PCS_RXTEST_PWR_REDUCTION: string  := "NORMAL";
        PCS_WA_SOS_DET_TOL: integer := 0;
        PCS_WA_SE_DET_TOL: integer := 0;
        PCS_RX_SAMPLE_UNION: string  := "FALSE";
        PCS_NEAR_LOOP   : string  := "FALSE";
        PCS_BYPASS_WORD_ALIGN: string  := "FALSE";
        PCS_BYPASS_DENC : string  := "FALSE";
        PCS_RX_ERRCNT_CLR: string  := "FALSE";
        PCS_RX_CODE_MODE: string  := "DUAL_8B10B";
        PCS_RX_BYPASS_GEAR: string  := "FALSE";
        PCS_ERRDETECT_SILENCE: string  := "FALSE";
        PCS_RX_DATA_MODE: string  := "8BIT";
        PCS_CA_DYN_CLY_EN_RX: string  := "FALSE";
        PCS_CFG_APATTERN_STATUS_DELAY: string  := "DELAY_ONE_CYCLE";
        PCS_RX_PRBS_MODE: string  := "DISABLE";
        PCS_ALIGN_MODE  : string  := "1GB";
        PCS_COMMA_DET_MODE: string  := "PATTERN_DETECT";
        PCS_RAPID_VMIN_1: integer := 0;
        PCS_RAPID_VMIN_2: integer := 0;
        PCS_RXBU_WIDER_EN: string  := "40/20BIT";
        PCS_RAPID_IMAX  : integer := 0;
        PCS_RX_SPLIT    : string  := "SPLIT_22BIT_11BIT";
        PCS_RXBRG_END_PACKET_9_8: integer := 0;
        PCS_RXBRG_END_PACKET_7_0: integer := 0;
        PCS_CTC_MAX_DEL : integer := 0;
        PCS_COMMA_REG0_9_8: integer := 0;
        PCS_COMMA_REG1_9_8: integer := 0;
        PCS_COMMA_MASK_9_8: integer := 0;
        PCS_COMMA_REG0_7_0: integer := 0;
        PCS_COMMA_REG1_7_0: integer := 0;
        PCS_COMMA_MASK_7_0: integer := 0;
        PCS_FLP_WRADDR_START: integer := 5;
        PCS_FLP_RDADDR_START: integer := 1;
        PCS_CFG_RX_BRIDGE_CLK_POLINV: string  := "FALSE";
        PCS_CTC_MODE_RD_SEL: string  := "NOMINAL_EMPTY";
        PCS_CTC_AFULL   : integer := 0;
        PCS_FAST_LOCK_GEAR_EN: string  := "FALSE";
        PCS_CTC_MODE_WR_SEL: string  := "NOMINAL_EMPTY";
        PCS_CTC_AEMPTY  : integer := 0;
        PCS_CTC_MODE    : string  := "ONE_BYTE";
        PCS_RXBRIDGE_MODE: string  := "BYPASS";
        PCS_CTC_ADD_MAX : integer := 0;
        PCS_CFG_PHDET_EN_RX: string  := "FALSE";
        PCS_WA_SDS_DET_TOL: integer := 0;
        PCS_CEB_MODE    : string  := "10GB";
        PCS_APATTERN_MODE: string  := "ONE_BYTE";
        PCS_A_REG0_8    : string  := "FALSE";
        PCS_RXBRG_WADDR_START: integer := 0;
        PCS_A_REG1_8    : string  := "FALSE";
        PCS_RXBRG_RADDR_START: integer := 0;
        PCS_A_REG0_7_0  : integer := 0;
        PCS_A_REG1_7_0  : integer := 0;
        PCS_CEB_RAPIDLS_MMAX: integer := 0;
        PCS_CEB_DETECT_TIME: integer := 0;
        PCS_WL_FIFO_RD  : integer := 0;
        PCS_SKIP_REG0_9_8: integer := 0;
        PCS_SKIP_REG0_7_0: integer := 0;
        PCS_CFG_CONTI_SKP_SET: integer := 0;
        PCS_CFG_RX_BASE_ADV_MODE: string  := "BASE_MODE";
        PCS_SKIP_REG1_9_8: integer := 0;
        PCS_SKIP_REG2_9_8: integer := 0;
        PCS_SKIP_REG3_9_8: integer := 0;
        PCS_SKIP_REG1_7_0: integer := 0;
        PCS_SKIP_REG2_7_0: integer := 0;
        PCS_SKIP_REG3_7_0: integer := 0;
        PCS_CFG_PRBS_ERR_O_SEL: integer := 0;
        PCS_CFG_PD_DELAY_RX: integer := 0;
        PCS_WR_START_GAP: integer := 0;
        PCS_MIN_IFG     : integer := 0;
        PCS_INT_RX_MASK_0: string  := "FALSE";
        PCS_INT_RX_MASK_1: string  := "FALSE";
        PCS_INT_RX_MASK_2: string  := "FALSE";
        PCS_INT_RX_MASK_3: string  := "FALSE";
        PCS_INT_RX_MASK_4: string  := "FALSE";
        PCS_INT_RX_MASK_5: string  := "FALSE";
        PCS_INT_RX_CLR_5: string  := "FALSE";
        PCS_INT_RX_CLR_4: string  := "FALSE";
        PCS_INT_RX_CLR_3: string  := "FALSE";
        PCS_INT_RX_CLR_2: string  := "FALSE";
        PCS_INT_RX_CLR_1: string  := "FALSE";
        PCS_INT_RX_CLR_0: string  := "FALSE";
        PCS_EM_CNT_RD_EN: string  := "FALSE";
        PCS_EM_CTRL_SEL : string  := "SIGNAL_CTRL";
        PCS_EM_MODE_CTRL: string  := "HOLD";
        PCS_EM_RD_CONDITION: string  := "TRIGGER";
        PCS_EM_SP_PATTERN_7_0: integer := 0;
        PCS_EM_SP_PATTERN_15_8: integer := 0;
        PCS_EM_SP_PATTERN_23_16: integer := 0;
        PCS_EM_SP_PATTERN_31_24: integer := 0;
        PCS_EM_SP_PATTERN_39_32: integer := 0;
        PCS_EM_SP_PATTERN_47_40: integer := 0;
        PCS_EM_SP_PATTERN_55_48: integer := 0;
        PCS_EM_SP_PATTERN_63_56: integer := 0;
        PCS_EM_SP_PATTERN_71_64: integer := 0;
        PCS_EM_SP_PATTERN_79_72: integer := 0;
        PCS_EM_PMA_MASK_7_0: integer := 0;
        PCS_EM_PMA_MASK_15_8: integer := 0;
        PCS_EM_PMA_MASK_23_16: integer := 0;
        PCS_EM_PMA_MASK_31_24: integer := 0;
        PCS_EM_PMA_MASK_39_32: integer := 0;
        PCS_EM_PMA_MASK_47_40: integer := 0;
        PCS_EM_PMA_MASK_55_48: integer := 0;
        PCS_EM_PMA_MASK_63_56: integer := 0;
        PCS_EM_PMA_MASK_71_64: integer := 0;
        PCS_EM_PMA_MASK_79_72: integer := 0;
        PCS_EM_EYED_MASK_7_0: integer := 0;
        PCS_EM_EYED_MASK_15_8: integer := 0;
        PCS_EM_EYED_MASK_23_16: integer := 0;
        PCS_EM_EYED_MASK_31_24: integer := 0;
        PCS_EM_EYED_MASK_39_32: integer := 0;
        PCS_EM_EYED_MASK_47_40: integer := 0;
        PCS_EM_EYED_MASK_55_48: integer := 0;
        PCS_EM_EYED_MASK_63_56: integer := 0;
        PCS_EM_EYED_MASK_71_64: integer := 0;
        PCS_EM_EYED_MASK_79_72: integer := 0;
        PCS_EM_PRESCALE : integer := 0;
        PCS_CFG_TEST_STATUS_SEL: string  := "SEL_PMA_TEST_STATUS_INT";
        PCS_CFG_DIFF_CNT_BND_RX: integer := 0;
        PCS_CFG_FLT_SEL_RX: string  := "FALSE";
        PCS_FILTER_BND_RX: integer := 0;
        PCS_TCLK2FABRIC_DIV_RST_M: string  := "FALSE";
        PCS_TX_PMA_TCLK_POLINV: string  := "PMA_TCLK";
        PCS_TX_TCLK_POLINV: string  := "TCLK";
        PCS_PCS_TCLK_SEL: string  := "PMA_TCLK";
        PCS_GEAR_TCLK_SEL: string  := "PMA_TCLK";
        PCS_TX_BRIDGE_TCLK_SEL: string  := "TCLK";
        PCS_TCLK2ALIGNER_SEL: string  := "PMA_TCLK";
        CA_DYN_DLY_EN_TX: string  := "FALSE";
        PCS_TX_PCS_CLK_EN_SEL: string  := "HARDWIRED1";
        PCS_TX_GEAR_CLK_EN_SEL: string  := "HARDWIRED0";
        PCS_TCLK2FABRIC_DIV_EN: string  := "FALSE";
        PCS_TCLK2FABRIC_SEL: string  := "CLK2ALIGNER_N_DIV2";
        DLY_ADJUST_SIZE_TX: integer := 0;
        PCS_TX_PCS_TX_RSTN: string  := "FALSE";
        PCS_TX_CA_RSTN  : string  := "FALSE";
        PCS_TX_SLAVE    : string  := "MASTER";
        PCS_TX_CA       : integer := 0;
        PCS_CFG_PI_CLK_SEL: integer := 0;
        PCS_CFG_PI_CLK_EN_SEL: string  := "CLK_EN_ROLL";
        PCS_CFG_PI_STEP_SIZE_TX: integer := 0;
        PCS_CFG_SUM_THRESHOLD_TX: integer := 0;
        PCS_CFG_AVG_CYCLES_TX: integer := 0;
        PCS_CFG_NEGEDGE_EN_TX: string  := "FALSE";
        PCS_CFG_ALIGN_THRD_TX: integer := 0;
        PCS_CFG_SCAN_INTERVAL_TX: integer := 0;
        PCS_CFG_STEP_SIZE_TX: integer := 0;
        PCS_CFG_REV_CNT_LIMIT_TX: integer := 0;
        PCS_CFG_FILTER_CNT_SIZE_TX: integer := 0;
        PCS_CFG_PI_DEFAULT_TX: integer := 0;
        PCS_CFG_PHDET_EN_TX: string  := "FALSE";
        PCS_PMA_TX2RX_PLOOP_EN: string  := "FALSE";
        PCS_PMA_TX2RX_SLOOP_EN: string  := "FALSE";
        PCS_CFG_DYN_DLY_SEL_TX: string  := "FALSE";
        PCS_CFG_DLY_REC_SIZE_TX: integer := 0;
        PCS_TX_DATA_WIDTH_MODE: string  := "8BIT";
        PCS_TX_BYPASS_BRIDGE_UINT: string  := "FALSE";
        PCS_TX_BYPASS_BRIDGE_FIFO: string  := "FALSE";
        PCS_TX_BYPASS_GEAR: string  := "FALSE";
        PCS_TX_BYPASS_ENC: string  := "FALSE";
        PCS_TX_BYPASS_BIT_SLIP: string  := "FALSE";
        PCS_TX_BRIDGE_GEAR_SEL: string  := "FALSE";
        PCS_TXBRG_PWR_REDUCTION: string  := "NORMAL";
        PCS_TXGEAR_PWR_REDUCTION: string  := "NORMAL";
        PCS_TXENC_PWR_REDUCTION: string  := "NORMAL";
        PCS_TXBSLP_PWR_REDUCTION: string  := "NORMAL";
        PCS_TXPRBS_PWR_REDUCTION: string  := "NORMAL";
        PCS_TXBRG_FULL_CHK_EN: string  := "FALSE";
        PCS_TXBRG_EMPTY_CHK_EN: string  := "FALSE";
        PCS_TX_ENCODER_MODE: string  := "DUAL_8B10B";
        PCS_TX_PRBS_MODE: string  := "DISABLE";
        PCS_TX_DRIVE_REG_MODE: string  := "NO_CHANGE";
        PCS_TX_BIT_SLIP_CYCLES: integer := 0;
        PCS_TX_BASE_ADV_MODE: string  := "BASE";
        PCS_TX_GEAR_SPLIT: string  := "NO_SPILT";
        PCS_RX_BRIDGE_CLK_POLINV: string  := "N_CLK_INVERT";
        PCS_PRBS_ERR_LPBK: string  := "FALSE";
        PCS_TX_INSERT_ER: string  := "FALSE";
        PCS_ENABLE_PRBS_GEN: string  := "FALSE";
        PCS_FAR_LOOP    : string  := "FALSE";
        PCS_CFG_ENC_TYPE_EN: string  := "FALSE";
        PCS_TXBRG_WADDR_START: integer := 0;
        PCS_TXBRG_RADDR_START: integer := 0;
        PCS_CFG_TX_PIC_EN: string  := "DISABLE";
        PCS_CFG_PIC_DIRECT_INV: string  := "FALSE";
        PCS_CFG_PI_MOD_CLK_EN: string  := "FALSE";
        PCS_CFG_TX_MODULATOR_OW_EN: string  := "FALSE";
        PCS_CFG_TX_PI_SSC_MODE_EN: string  := "FALSE";
        PCS_CFG_TX_PI_OFFSET_MODE_EN: string  := "FALSE";
        PCS_CFG_TX_PI_SSC_MODE_SEL: integer := 0;
        PCS_CFG_TXDEEMPH_EN: string  := "FALSE";
        PCS_PI_STROBE_SEL: string  := "FALSE";
        PCS_CFG_TX_PIC_GREY_SEL: string  := "FALSE";
        PCS_CFG_PIC_RENEW_INV: string  := "NORMAL";
        PCS_CFG_NUM_PIC : integer := 0;
        PCS_CFG_TXPIC_OW_EN: string  := "FALSE";
        PCS_CFG_TXPPM_OW_VALUE_0_7: integer := 0;
        PCS_INT_TX_MASK_0: string  := "FALSE";
        PCS_INT_TX_MASK_1: string  := "FALSE";
        PCS_INT_TX_MASK_2: string  := "FALSE";
        PCS_INT_TX_CLR_2: string  := "FALSE";
        PCS_INT_TX_CLR_1: string  := "FALSE";
        PCS_INT_TX_CLR_0: string  := "FALSE";
        PCS_CFG_PD_DELAY_TX: integer := 0;
        PCS_CFG_DIFF_CNT_BND_TX: integer := 0;
        PCS_CFG_PD_CLK_FR_CORE_SEL: string  := "FALSE";
        PCS_CFG_FLT_SEL_TX: string  := "FALSE";
        PCS_FILTER_BND_TX: integer := 0;
        PCS_CFG_TX_SSC_PPM_RANGE_7_0: integer := 0;
        PCS_CFG_TX_PPM_MODULATOR_EN: string  := "FALSE";
        PCS_CFG_TX_PPM_SCALE2_SEL: integer := 0;
        PCS_CFG_TX_PPM_SCALE_SEL: integer := 0;
        PCS_CFG_TX_SSC_PPM_RANGE_8_9: integer := 0;
        PCS_CFG_TX_SSC_MODULATION_STEP_7_0: integer := 0;
        PCS_CFG_TX_SSC_PPM_OFFSET_7_0: integer := 0;
        PCS_CFG_TX_SSC_MODULATION_STEP_8: integer := 0;
        PCS_CFG_TX_SSC_PPM_OFFSET_8_9: integer := 0;
        PMA_REG_CHL_BIAS_POWER_SEL: string  := "FALSE";
        PMA_REG_CHL_BIAS_POWER: string  := "FALSE";
        PMA_REG_RX_BUSWIDTH: string  := "20BIT";
        PMA_REG_RX_RATE : string  := "DIV4";
        PMA_REG_RX_RATE_EN: string  := "TRUE";
        PMA_REG_RX_RES_TRIM: integer := 50;
        PMA_REG_RX_SIGDET_STATUS_EN: string  := "FALSE";
        PMA_REG_CDR_READY_THD_7_0: integer := 174;
        PMA_REG_CDR_READY_THD_11_8: integer := 10;
        PMA_REG_RX_BUSWIDTH_EN: string  := "FALSE";
        PMA_REG_RX_PCLK_EDGE_SEL: string  := "POS_EDGE";
        PMA_REG_CDR_READY_CHECK_CTRL: integer := 3;
        PMA_REG_RX_ICTRL_TRX: string  := "100PCT";
        PMA_REG_PRBS_CHK_WIDTH_SEL: integer := 0;
        PMA_REG_RX_ICTRL_PIBUF: string  := "100PCT";
        PMA_REG_RX_ICTRL_PI: string  := "100PCT";
        PMA_REG_RX_ICTRL_DCC: string  := "100PCT";
        PMA_REG_RX_TX2RX_PLPBK_EN: string  := "FALSE";
        PMA_REG_RX_DATA_POLARITY: string  := "NORMAL";
        PMA_REG_RX_ERR_INSERT: string  := "FALSE";
        PMA_REG_UDP_CHK_EN: string  := "FALSE";
        PMA_REG_PRBS_SEL: string  := "PRBS7";
        PMA_REG_PRBS_CHK_EN: string  := "FALSE";
        PMA_REG_LPLL_NFC_STIC_DIS_N: integer := 0;
        PMA_REG_BIST_CHK_PAT_SEL: string  := "PRBS";
        PMA_REG_LOAD_ERR_CNT: string  := "FALSE";
        PMA_REG_CHK_COUNTER_EN: string  := "FALSE";
        PMA_REG_CDR_PROP_GAN_SEL: integer := 5;
        PMA_REG_CDR_TUBO_PROP_GAIN_SEL: integer := 6;
        PAM_REG_CDR_INT_GAIN_SEL: integer := 5;
        PMA_REG_CDR_TUBO_INT_GAIN_SEL: integer := 6;
        PMA_REG_CDR_INT_SAT_MAX_4_0: integer := 0;
        PMA_REG_CDR_INT_SAT_MAX_9_5: integer := 31;
        PMA_REG_CDR_INT_SAT_MIN_2_0: integer := 0;
        PMA_REG_CDR_INT_SAT_MIN_9_3: integer := 4;
        PMA_ANA_RX_REG_O_61_55: integer := 21;
        PMA_ANA_RX_REG_O_69_62: integer := 0;
        PMA_ANA_RX_REG_O_77_70: integer := 1;
        PMA_ANA_RX_REG_O_85_78: integer := 1;
        PMA_ANA_RX_REG_O_93_86: integer := 65;
        PMA_ANA_RX_REG_O_100_94: integer := 69;
        PMA_ANA_RX_REG_O_108_101: integer := 0;
        PMA_ANA_RX_REG_O_111_109: integer := 0;
        PMA_REG_OOB_COMWAKE_GAP_MIN_4_0: integer := 3;
        PMA_REG_OOB_COMWAKE_GAP_MIN_5: integer := 0;
        PMA_REG_OOB_COMWAKE_GAP_MAX: integer := 11;
        PMA_REG_OOB_COMINIT_GAP_MIN: integer := 15;
        PMA_REG_OOB_COMINIT_GAP_MAX: integer := 35;
        PMA_REG_COMWAKE_STATUS_CLEAR: integer := 0;
        PMA_REG_COMINIT_STATUS_CLEAR: integer := 0;
        PMA_REG_RX_SATA_COMINIT_OW: string  := "FALSE";
        PMA_REG_RX_SATA_COMINIT: string  := "FALSE";
        PMA_REG_RX_SATA_COMWAKE_OW: string  := "FALSE";
        PMA_REG_RX_SATA_COMWAKE: string  := "FALSE";
        PMA_REG_RX_DCC_DISABLE: string  := "FALSE";
        PMA_REG_RX_SLIP_SEL_EN: string  := "FALSE";
        PMA_REG_RX_SLIP_SEL: integer := 0;
        PMA_REG_RX_SLIP_EN: string  := "FALSE";
        PMA_REG_RX_SIGDET_STATUS_SEL: integer := 5;
        PMA_REG_RX_SIGDET_FSM_RST_N: string  := "TRUE";
        PMA_REG_RX_SIGDET_STATUS: string  := "FALSE";
        PMA_REG_RX_SIGDET_VTH: string  := "27MV";
        PMA_REG_RX_SIGDET_GRM: integer := 0;
        PMA_REG_RX_SIGDET_PULSE_EXT: string  := "FALSE";
        PMA_REG_RX_SIGDET_CH2_SEL: integer := 0;
        PMA_REG_RX_SIGDET_CH2_CHK_WINDOW: integer := 3;
        PMA_REG_RX_SIGDET_CHK_WINDOW_EN: string  := "TRUE";
        PMA_REG_RX_SIGDET_NOSIG_COUNT_SETTING: integer := 4;
        PMA_REG_RX_SIGDET_OOB_DET_COUNT_VAL_2_0: integer := 0;
        PMA_REG_RX_SIGDET_OOB_DET_COUNT_VAL_4_3: integer := 0;
        PMA_REG_RX_SIGDET_4OOB_DET_SEL: integer := 7;
        PMA_REG_RX_SIGDET_IC_I: integer := 10;
        PMA_REG_RX_EQ1_R_SET_TOP: integer := 0;
        PMA_REG_RX_EQ1_C_SET_FB: integer := 0;
        PMA_REG_RX_EQ1_OFF: string  := "FALSE";
        PMA_REG_RX_EQ2_R_SET_TOP: integer := 3;
        PMA_REG_RX_EQ2_C_SET_FB: integer := 0;
        PMA_REG_RX_EQ2_OFF: string  := "FALSE";
        PMA_REG_RX_ICTRL_EQ: integer := 2;
        PMA_REG_EQ_DC_CALIB_EN: string  := "FALSE";
        PMA_CTLE_CTRL_REG_I: integer := 0;
        PMA_CTLE_REG_FORCE_SEL_I: string  := "FALSE";
        PMA_CTLE_REG_HOLD_I: string  := "FALSE";
        PMA_CTLE_REG_INIT_DAC_I_1_0: integer := 0;
        PMA_CTLE_REG_INIT_DAC_I_3_2: integer := 0;
        PMA_CTLE_REG_POLARITY_I: string  := "FALSE";
        PMA_CTLE_REG_SHIFTER_GAIN_I: integer := 0;
        PMA_CTLE_REG_THRESHOLD_I_1_0: integer := 0;
        PMA_CTLE_REG_THRESHOLD_I_9_2: integer := 1;
        PMA_CTLE_REG_THRESHOLD_I_11_10: integer := 0;
        PMA_REG_RX_RES_TRIM_EN: string  := "TRUE";
        PMA_REG_ALG_RX_TERM_POWER_DIVIDING_SELECTION: integer := 1;
        PMA_REG_ALG_RX_TERM_VCM_SELECTION: integer := 3;
        PMA_REG_ALG_RX_TERM_TEST_SELECTION_7_0: integer := 0;
        PMA_REG_ALG_RX_TERM_TEST_SELECTION_9_8: integer := 0;
        PMA_REG_ALG_LOW_SPEED_MODE_ENABLE: string  := "FALSE";
        PMA_REG_ALG_RX_CLOCK_POWER_DOWN_REGISTER: string  := "TRUE";
        PMA_REG_ALG_RX_CLOCK_POWER_DOWN_SELECTION: string  := "FALSE";
        PMA_REG_ALG_RX_DFE_POWER_DOWN_REGISTER_0: string  := "TRUE";
        PMA_REG_ALG_RX_DFE_POWER_DOWN_SELECTION_1: string  := "FALSE";
        PMA_REG_ALG_RX_CTLE_POWER_DOWN_REGISTER_0: string  := "TRUE";
        PMA_REG_ALG_RX_CTLE_POWER_DOWN_SELECTION_1: string  := "FALSE";
        PMA_REG_EYE_DFETAP1_PLORITY: string  := "TRUE";
        PMA_REG_CDR_SEL : string  := "FALSE";
        PMA_REG_EYE_DET_EN: string  := "TRUE";
        PMA_REG_PI_BIAS_CURRENT: integer := 0;
        PMA_REG_ALG_DFE_TEST_SEL_6_0: integer := 0;
        PMA_REG_ALG_DFE_TEST_SEL_14_7: integer := 0;
        PMA_REG_ALG_DFE_TEST_SEL_21_15: integer := 0;
        PMA_REG_ALG_CTLE_TEST_SEL: integer := 0;
        PMA_REG_ALG_ANA_RX_SLIP_SEL_O: string  := "FALSE";
        PMA_REG_ALG_RX_T1_BUFF_EN: string  := "FALSE";
        PMA_REG_ALG_RX_CDRX_BUFF_EN: string  := "FALSE";
        PMA_REG_ALG_RX_VP_T1_SW_PLORITY: string  := "FALSE";
        PMA_REG_ALG_RX_VP_PLORITY: string  := "FALSE";
        PMA_REG_ALG_RX_GAIN_CTRL_SUMMER: string  := "FALSE";
        PMA_REG_ALG_RX_DC_OFFSET_T1_EN: string  := "FALSE";
        PMA_REG_ALG_RX_DC_OFFSET_VP_EN: string  := "FALSE";
        PMA_REG_ALG_RX_DC_OFFSET_CDRX_EN: string  := "FALSE";
        PMA_REG_ALG_RX_DC_OFFSET_CDRY_EN: string  := "FALSE";
        PMA_REG_ALG_RX_DC_OFFSET_EYE_EN: string  := "FALSE";
        PMA_REG_ALG_SLICER_DC_OFFSET_OVERWITE: string  := "FALSE";
        PMA_REG_ALG_SLICER_DC_OFFSET_REG: string  := "FALSE";
        PMA_REG_ALG_SHUT_OFF_THE_EQUALIZER_OF_EACH_STAGE: string  := "FALSE";
        PMA_REG_ALG_CDR_XWEIGHT_I: integer := 4;
        PMA_REG_ALG_CDR_YWEIGHT_I: integer := 4;
        PMA_REG_ALG_CTLE_FLIPDIR_I: string  := "TRUE";
        PMA_REG_ALG_CTLE_HOLD_I: string  := "FALSE";
        PMA_REG_ALG_CTLE_INITDAC_5_0: integer := 0;
        PMA_REG_ALG_CTLE_INITDAC_6: integer := 0;
        PMA_REG_ALG_CTLE_OVERWREN_I: string  := "FALSE";
        PMA_REG_ALG_CTLE_SHIFT_I: integer := 4;
        PMA_REG_ALG_CTLE_TOPNUM_2_0: integer := 4;
        PMA_REG_ALG_CTLE_TOPNUM_4_3: integer := 2;
        PMA_REG_ALG_CTLEOFS_FLIPDIR_I: string  := "FALSE";
        PMA_REG_ALG_CTLEOFS_HOLD_I: string  := "FALSE";
        PMA_REG_ALG_CTLEOFS_INITDAC_3_0: integer := 0;
        PMA_REG_ALG_CTLEOFS_INITDAC_6_4: integer := 4;
        PMA_REG_ALG_CTLEOFS_OVERWREN: string  := "FALSE";
        PMA_REG_ALG_CTLEOFS_SHIFT_I: integer := 4;
        PMA_REG_ALG_DFE_CTLE_PWD: string  := "TRUE";
        PMA_REG_ALG_H1_FLIPDIR_I: string  := "FALSE";
        PMA_REG_ALG_H1_HOLD_I: string  := "FALSE";
        PMA_REG_ALG_H1_INITDAC_5_0: integer := 0;
        PMA_REG_ALG_H1_INITDAC_6: integer := 0;
        PMA_REG_ALG_H1_OVERWREN_I: string  := "FALSE";
        PMA_REG_ALG_H1_SHIFT_I: integer := 4;
        PMA_REG_ALG_H2_FLIPDIR_I: string  := "FALSE";
        PMA_REG_ALG_H2_HOLD_I: string  := "FALSE";
        PMA_REG_ALG_H2_INITDAC_0: integer := 0;
        PMA_REG_ALG_H2_INITDAC_5_1: integer := 0;
        PMA_REG_ALG_H2_OVERWREN_I: string  := "FALSE";
        PMA_REG_ALG_H2_SHIFT_I_1_0: integer := 0;
        PMA_REG_ALG_H2_SHIFT_I_2: integer := 1;
        PMA_REG_ALG_H3_FLIPDIR_I: string  := "FALSE";
        PMA_REG_ALG_H3_HOLD_I: string  := "FALSE";
        PMA_REG_ALG_H3_INITDAC_4_0: integer := 0;
        PMA_REG_ALG_H3_INITDAC_5: integer := 1;
        PMA_REG_ALG_H3_OVERWREN_I: string  := "FALSE";
        PMA_REG_ALG_H3_SHIFT_I: integer := 4;
        PMA_REG_ALG_H4_FLIPDIR_I: string  := "FALSE";
        PMA_REG_ALG_H4_HOLD_I: string  := "FALSE";
        PMA_REG_ALG_H4_INITDAC_0: integer := 0;
        PMA_REG_ALG_H4_INITDAC_4_1: integer := 8;
        PMA_REG_ALG_H4_OVERWREN_I: string  := "FALSE";
        PMA_REG_ALG_H4_SHIFT_I: integer := 4;
        PMA_REG_ALG_H5_FLIPDIR_I: string  := "FALSE";
        PMA_REG_ALG_H5_HOLD_I: string  := "FALSE";
        PMA_REG_ALG_H5_INITDAC: integer := 16;
        PMA_REG_ALG_H5_OVERWREN_I: string  := "FALSE";
        PMA_REG_ALG_H5_SHIFT_I: integer := 4;
        PMA_REG_ALG_H6_FLIPDIR_I: string  := "FALSE";
        PMA_REG_ALG_H6_HOLD_I: string  := "FALSE";
        PMA_REG_ALG_H6_INITDAC_2_0: integer := 0;
        PMA_REG_ALG_H6_INITDAC_4_3: integer := 2;
        PMA_REG_ALG_H6_OVERWREN_I: string  := "FALSE";
        PMA_REG_ALG_H6_SHIFT_I: integer := 4;
        PMA_REG_ALG_HCTLE_OFS_1_0: integer := 0;
        PMA_REG_ALG_HCTLE_OFS_3_2: integer := 2;
        PMA_REG_ALG_HCTLE_OVERWRDAC_5_0: integer := 0;
        PMA_REG_ALG_HCTLE_OVERWRDAC_6: integer := 1;
        PMA_REG_ALG_HCTLE_OVERWREN: string  := "FALSE";
        PMA_REG_ALG_LPMH_INITDAC_I: integer := 0;
        PMA_REG_ALG_LPMH_PWD_I: string  := "TRUE";
        PMA_REG_ALG_LPMH_REG_HOLD_I: string  := "FALSE";
        PMA_REG_ALG_LPMH_REG_SHIFT_I: integer := 4;
        PMA_REG_ALG_LPML_INITDAC_I: integer := 0;
        PMA_REG_ALG_LPML_PWD_I: string  := "TRUE";
        PMA_REG_ALG_LPML_REG_HOLD_I: string  := "FALSE";
        PMA_REG_ALG_LPML_REG_PRESELECT_I: integer := 7;
        PMA_REG_ALG_LPML_REG_SHIFT_I: integer := 4;
        PMA_REG_ALG_NEXTBIT_I: string  := "FALSE";
        PMA_REG_ALG_SOFS_COUNTMAX_I_6_0: integer := 127;
        PMA_REG_ALG_SOFS_COUNTMAX_I_14_7: integer := 255;
        PMA_REG_ALG_SOFS_COUNTMAX_I_19_15: integer := 31;
        PMA_REG_ALG_SOFS_DACWIN_I: integer := 1;
        PMA_REG_ALG_SOFS_FLIP_DIR_I: string  := "TRUE";
        PMA_REG_ALG_SOFS_FORCE_I: string  := "FALSE";
        PMA_REG_ALG_SOFS_FORCEDAC_I_5_0: integer := 0;
        PMA_REG_ALG_SOFS_FORCEDAC_I_6: integer := 1;
        PMA_REG_ALG_SOFS_FORCENUM_I: integer := 0;
        PMA_REG_ALG_SOFS_INITDAC_2_0: integer := 0;
        PMA_REG_ALG_SOFS_INITDAC_6_3: integer := 8;
        PMA_REG_ALG_SOFS_SHIFT_I: integer := 1;
        PMA_REG_ALG_SOFS_SKIP_I: string  := "FALSE";
        PMA_REG_ALG_SOFS_WINCOUNTMAX_I_7_0: integer := 0;
        PMA_REG_ALG_SOFS_WINCOUNTMAX_I_11_8: integer := 4;
        PMA_REG_ALG_ST_FLIPDIR_I: string  := "TRUE";
        PMA_REG_ALG_ST_FORCEN: string  := "FALSE";
        PMA_REG_ALG_ST_HOLD_I: string  := "FALSE";
        PMA_REG_ALG_ST_INITDAC_0: integer := 0;
        PMA_REG_ALG_ST_INITDAC_4_1: integer := 8;
        PMA_REG_ALG_ST_RECALEN: string  := "FALSE";
        PMA_REG_ALG_ST_SHIFT_I: integer := 4;
        PMA_REG_ALG_ST_STARTCNT_7_0: integer := 0;
        PMA_REG_ALG_ST_STARTCNT_15_8: integer := 128;
        PMA_REG_ALG_ST_STARTCNT_19_16: integer := 0;
        PMA_REG_ALG_ST_TAPCNT_3_0: integer := 0;
        PMA_REG_ALG_ST_TAPCNT_11_4: integer := 0;
        PMA_REG_ALG_ST_TAPCNT_17_12: integer := 2;
        PMA_REG_ALG_ST_TOPTAP_1_0: integer := 3;
        PMA_REG_ALG_ST_TOPTAP_3_2: integer := 3;
        PMA_REG_ALG_SWCLK_DIV: integer := 0;
        PMA_REG_ALG_TAPA_DAC_3_0: integer := 0;
        PMA_REG_ALG_TAPA_DAC_4: integer := 1;
        PMA_REG_ALG_TAPA_NUM: integer := 7;
        PMA_REG_ALG_TAPB_DAC_0: integer := 0;
        PMA_REG_ALG_TAPB_DAC_4_1: integer := 8;
        PMA_REG_ALG_TAPB_NUM_3_0: integer := 8;
        PMA_REG_ALG_TAPB_NUM_5_4: integer := 0;
        PMA_REG_ALG_TAPC_DAC: integer := 16;
        PMA_REG_ALG_TAPC_NUM_0: integer := 1;
        PMA_REG_ALG_TAPC_NUM_5_1: integer := 4;
        PMA_REG_ALG_TAPD_DAC_2_0: integer := 0;
        PMA_REG_ALG_TAPD_DAC_4_3: integer := 2;
        PMA_REG_ALG_TAPD_NUM: integer := 10;
        PMA_REG_ALG_VP_FLIPDIR_I: string  := "FALSE";
        PMA_REG_ALG_VP_GRN_SHIFT_I: integer := 5;
        PMA_REG_ALG_VP_HOLD_I: string  := "FALSE";
        PMA_REG_ALG_VP_IDEAL_2_0: integer := 0;
        PMA_REG_ALG_VP_IDEAL_6_3: integer := 10;
        PMA_REG_ALG_VP_INITDAC_I_3_0: integer := 0;
        PMA_REG_ALG_VP_INITDAC_I_6_4: integer := 0;
        PMA_REG_ALG_VP_OVERWREN: string  := "FALSE";
        PMA_REG_ALG_VP_RED_SHIFT_I: integer := 5;
        PMA_REG_ALG_VPOFS_SEL_0: integer := 0;
        PMA_REG_ALG_VPOFS_SEL_2_1: integer := 1;
        PMA_REG_ALG_H1_UPBOUND_5_0: integer := 55;
        PMA_REG_ALG_H1_UPBOUND_6: integer := 1;
        PMA_REG_ALG_CTLEOFS_PWDN: string  := "FALSE";
        PMA_REG_ALG_LPMH_OVEREN_I: string  := "FALSE";
        PMA_REG_ALG_LPML_OVEREN_I: string  := "FALSE";
        PMA_REG_ALG_AGC_FLIPDIR_I: string  := "FALSE";
        PMA_REG_ALG_AGC_HOLD_I: string  := "FALSE";
        PMA_REG_ALG_AGC_INITDAC: integer := 10;
        PMA_REG_ALG_AGC_LOWBOUND_1_0: integer := 3;
        PMA_REG_ALG_AGC_LOWBOUND_3_2: integer := 0;
        PMA_REG_ALG_AGC_OVERWREN_I: string  := "FALSE";
        PMA_REG_ALG_AGC_PWD: string  := "TRUE";
        PMA_REG_ALG_AGC_SHIFT_I: integer := 4;
        PMA_REG_ALG_AGC_UPBOUND_0: integer := 1;
        PMA_REG_ALG_AGC_UPBOUND_3_1: integer := 7;
        PMA_REG_ALG_AGC_WAITSEL: integer := 11;
        PMA_REG_PI_CTRL_SEL_RX: string  := "FALSE";
        PMA_REG_PI_CTRL_RX_4_0: integer := 0;
        PMA_REG_PI_CTRL_RX_7_5: integer := 0;
        PMA_CFG_RX_LANE_POWERUP: string  := "OFF";
        PMA_CFG_RX_PMA_RSTN: string  := "FALSE";
        PMA_INT_PMA_RX_MASK_0: string  := "FALSE";
        PMA_INT_PMA_RX_CLR_0: string  := "FALSE";
        PMA_CFG_CTLE_ADP_RSTN: string  := "FALSE";
        PMA_CFG_RX_CDR_RSTN: string  := "FALSE";
        PMA_CFG_RX_CLKPATH_RSTN: string  := "FALSE";
        PMA_CFG_RX_DFE_RSTN: string  := "FALSE";
        PMA_CFG_RX_LPM_RSTN: string  := "FALSE";
        PMA_CFG_RX_SLIDING_RSTN: string  := "FALSE";
        PMA_CFG_RX_EYE_RSTN: string  := "FALSE";
        PMA_CFG_RX_CTLE_DCCAL_RSTN: string  := "FALSE";
        PMA_CFG_RX_SLICER_DCCAL_RSTN: string  := "FALSE";
        PMA_CFG_RX_SLIP_RSTN: string  := "FALSE";
        PMA_REG_TX_PD_MINOR: string  := "ON";
        PMA_REG_TX_PD_MINOR_OW: string  := "TRUE";
        PMA_REG_TX_MAIN_PRE_Z: string  := "FALSE";
        PMA_REG_TX_MAIN_PRE_Z_OW: string  := "FALSE";
        PMA_REG_TX_BEACON_TIMER_SEL: integer := 0;
        PMA_REG_TX_RXDET_REQ_OW: string  := "FALSE";
        PMA_REG_TX_RXDET_REQ: string  := "FALSE";
        PMA_REG_TX_BEACON_EN_OW: string  := "TRUE";
        PMA_REG_TX_BEACON_EN: string  := "FALSE";
        PMA_REG_TX_EI_EN_OW: string  := "FALSE";
        PMA_REG_TX_EI_EN: string  := "FALSE";
        PMA_REG_TX_BIT_CONV: string  := "FALSE";
        PMA_REG_TX_RES_CAL: integer := 50;
        PMA_REG_TX_UDP_DATA_20: integer := 0;
        PMA_REG_TX_UDP_DATA_26_21: integer := 0;
        PMA_REG_TX_UDP_DATA_34_27: integer := 0;
        PMA_REG_TX_UDP_DATA_39_25: integer := 0;
        PMA_REG_TX_PD_MAIN: integer := 0;
        PMA_REG_TX_PD_MAIN_OW: integer := 0;
        PMA_REG_TX_BUSWIDTH_EN: integer := 0;
        PMA_REG_TX_SYNC_OW: string  := "FALSE";
        PMA_REG_TX_SYNC : string  := "TRUE";
        PMA_REG_TX_PD_POST: string  := "OFF";
        PMA_REG_TX_PD_POST_OW: string  := "TRUE";
        PMA_REG_TX_RESET_N_OW: string  := "FALSE";
        PMA_REG_TX_RESET_N: string  := "TRUE";
        PMA_REG_PMA_TX_RESET_N: string  := "FALSE";
        PMA_REG_PMA_TX_RESET_N_OW: string  := "FALSE";
        PMA_REG_TX_BUSWIDTH: string  := "20BIT";
        PMA_REG_PLL_READY_OW: string  := "FALSE";
        PMA_REG_PLL_READY: string  := "TRUE";
        PMA_REG_EI_PCLK_DELAY_SEL: integer := 0;
        PMA_REG_TX_AMP_DAC0: integer := 25;
        PMA_REG_TX_AMP_DAC1: integer := 19;
        PMA_REG_TX_AMP_DAC2: integer := 14;
        PMA_REG_TX_AMP_DAC3: integer := 9;
        PMA_REG_TX_MARGIN: integer := 0;
        PMA_REG_TX_MARGIN_OW: string  := "TRUE";
        PMA_REG_TX_SWING: string  := "FALSE";
        PMA_REG_TX_SWING_OW: string  := "TRUE";
        PMA_REG_TX_RXDET_THRESHOLD: string  := "84MV";
        PMA_REG_TX_BEACON_OSC_CTRL: string  := "FALSE";
        PMA_REG_TX_PRBS_GEN_WIDTH_SEL: integer := 0;
        PMA_REG_TX_TX2RX_SLPBACK_EN: string  := "FALSE";
        PMA_REG_TX_PCLK_EDGE_SEL: string  := "FALSE";
        PMA_REG_TX_RXDET_STATUS_OW: string  := "FALSE";
        PMA_REG_TX_RXDET_STATUS: string  := "FALSE";
        PMA_REG_TX_PRBS_GEN_EN: string  := "FALSE";
        PMA_REG_TX_PRBS_SEL: string  := "PRBS7";
        PMA_REG_TX_UDP_DATA_7_TO_0: integer := 0;
        PMA_REG_TX_UDP_DATA_15_TO_8: integer := 0;
        PMA_REG_TX_UDP_DATA_19_TO_16: integer := 0;
        PMA_REG_TX_FIFO_WP_CTRL: integer := 4;
        PMA_REG_TX_FIFO_EN: string  := "FALSE";
        PMA_REG_TX_DATA_MUX_SEL: integer := 0;
        PMA_REG_TX_ERR_INSERT: string  := "FALSE";
        PMA_REG_TX_SATA_EN: string  := "FALSE";
        PMA_REG_RATE_CHANGE_TXPCLK_ON_OW: string  := "FALSE";
        PMA_REG_RATE_CHANGE_TXPCLK_ON: string  := "TRUE";
        PMA_REG_TX_CFG_POST1: integer := 0;
        PMA_REG_TX_CFG_POST2: integer := 0;
        PMA_REG_TX_DEEMP: integer := 0;
        PMA_REG_TX_DEEMP_O: string  := "TRUE";
        PMA_REG_TX_OOB_DELAY_SEL: integer := 0;
        PMA_REG_TX_POLARITY: string  := "NORMAL";
        PMA_REG_ANA_TX_JTAG_DATA_O_SEL: string  := "FALSE";
        PMA_REG_TX_LS_MODE_EN: string  := "FALSE";
        PMA_REG_TX_JTAG_MODE_EN_OW: string  := "TRUE";
        PMA_REG_TX_JTAG_MODE_EN: string  := "TRUE";
        PMA_REG_RX_JTAG_MODE_EN_OW: string  := "TRUE";
        PMA_REG_RX_JTAG_MODE_EN: string  := "TRUE";
        PMA_REG_RX_JTAG_OE: string  := "FALSE";
        PMA_REG_RX_ACJTAG_VHYSTSEL: integer := 0;
        PMA_REG_TX_RES_CAL_EN: string  := "FALSE";
        PMA_REG_RX_TERM_MODE_CTRL: integer := 5;
        PMA_REG_PLPBK_TXPCLK_EN: string  := "FALSE";
        PMA_REG_CLK_SEL_STROBE_TXPCLK: integer := 0;
        PMA_REG_TX_PH_SEL_0: integer := 1;
        PMA_REG_TX_PH_SEL_6_1: integer := 0;
        PMA_REG_TX_CFG_PRE: integer := 0;
        PMA_REG_TX_CFG_MAIN: integer := 0;
        PMA_REG_CFG_POST: integer := 0;
        PMA_REG_PD_MAIN : string  := "FALSE";
        PMA_REG_PD_PRE  : string  := "TRUE";
        PMA_REG_TX_LS_DATA: string  := "FALSE";
        PMA_REG_TX_DCC_BUF_SZ_SEL: integer := 0;
        PMA_REG_TX_DCC_CAL_CUR_TUNE: integer := 0;
        PMA_REG_TX_DCC_CAL_EN: string  := "FALSE";
        PMA_REG_TX_DCC_CUR_SS: integer := 0;
        PMA_REG_TX_DCC_FA_CTRL: string  := "FALSE";
        PMA_REG_TX_DCC_RI_CTRL: string  := "FALSE";
        PMA_REG_ATB_SEL_2_0: integer := 0;
        PMA_REG_ATB_SEL_9_3: integer := 0;
        PMA_REG_TX_CFG_7_0: integer := 0;
        PMA_REG_TX_CFG_15_8: integer := 0;
        PMA_REG_TX_CFG_23_16: integer := 0;
        PMA_REG_TX_CFG_31_24: integer := 0;
        PMA_REG_TX_OOB_EI_EN: string  := "FALSE";
        PMA_REG_TX_OOB_EI_EN_OW: string  := "FALSE";
        PMA_REG_TX_BEACON_EN_DELAYED: string  := "FALSE";
        PMA_REG_TX_BEACON_EN_DELAYED_OW: string  := "FALSE";
        PMA_REG_TX_JTAG_DATA: string  := "FALSE";
        PMA_REG_TX_RXDET_TIMER_SEL: integer := 87;
        PMA_REG_TX_CFG1_7_0: integer := 0;
        PMA_REG_TX_CFG1_15_8: integer := 0;
        PMA_REG_TX_CFG1_23_16: integer := 0;
        PMA_REG_TX_CFG1_31_24: integer := 0;
        PMA_REG_TX_PI_CUR_BUF: string  := "525uA";
        PMA_REG_TX_ATB_4_0: integer := 0;
        PMA_REG_TX_ATB_9_5: integer := 0;
        PMA_REG_TX_MOD_STAND_BY_EN: string  := "FALSE";
        PMA_REG_STATE_STAND_BY_SEL: string  := "FALSE";
        PMA_REG_TX_PISO_PD: string  := "TRUE";
        PMA_REG_TX_PISO_PD_OW: string  := "FALSE";
        PMA_REG_TX_CLK_PD: string  := "TRUE";
        PMA_REG_TX_CLK_PD_OW: string  := "FALSE";
        PMA_REG_TX_DRIVER_PD: string  := "FALSE";
        PMA_REG_TX_DRIVER_PD_OW: string  := "FALSE";
        PMA_REG_TX_SYNC_NEW: string  := "TRUE";
        PMA_REG_TX_SYNC_NEW_OW: string  := "FALSE";
        PMA_REG_TX_CHANGE_ON_OW: string  := "FALSE";
        PMA_REG_TX_CHANGE_ON_POLAR_CTRL: string  := "FALSE";
        PMA_REG_TX_FREERUN_PD: string  := "TRUE";
        PMA_REG_TX_CHANGE_ON_SEL: string  := "FALSE";
        PMA_REG_TX_CHANGE_ON_CTRL: string  := "FALSE";
        PMA_REG_TX_PIDC_CURRENT_EN: integer := 0;
        PMA_REG_TX_FREERUN_RATE_0: integer := 0;
        PMA_REG_TX_FREERUN_RATE_1: integer := 1;
        PMA_REG_TX_FREERUN_RATE_OW: string  := "FALSE";
        PMA_REG_TX_VBIAS_REG_SEL: string  := "FALSE";
        PMA_REG_TX_VBIAS_DIVIDER_SEL: integer := 0;
        PMA_REG_TX_RST_SYNC_CLK_SEL: string  := "TRUE";
        PMA_REG_TX_PI_CTRL_SEL: integer := 0;
        PMA_REG_TX_PI_CTRL: integer := 0;
        PMA_LANE_POWERUP: string  := "FALSE";
        PMA_POR_N       : string  := "FALSE";
        PMA_TX_LANE_POWERUP: string  := "FALSE";
        PMA_TX_PMA_RSTN : string  := "FALSE";
        PMA_LPLL_POWERUP: string  := "FALSE";
        PMA_LPLL_RSTN   : string  := "FALSE";
        PMA_LPLL_LOCKDET_RSTN: string  := "FALSE";
        PMA_REG_LPLL_PFDDELAY_SEL: integer := 1;
        PMA_REG_LPLL_PFDDELAY_EN: string  := "TRUE";
        PMA_REG_LPLL_VCTRL_SET: integer := 0;
        PMA_LPLL_CHARGE_PUMP_CTRL: string  := "type";
        PMA_LPLL_REFDIV : string  := "DIV1";
        PMA_LPLL_FBDIV  : integer := 36;
        PMA_LPLL_LPF_RES: integer := 1;
        PMA_LPLL_TEST_SEL: integer := 0;
        PMA_LPLL_TEST_SIG_HALF_EN: string  := "TRUE";
        PMA_LPLL_TEST_V_EN: string  := "FALSE";
        PMA_REG_BUF_BIAS_SEL: string  := "46.875u";
        PMA_REG_TXCLK_SEL: string  := "LPLL";
        PMA_REG_RXCLK_SEL: string  := "LPLL";
        PMA_REG_TEST_BUF: integer := 0;
        PMA_REG_RX_DEF_SEL0: string  := "25uA";
        PMA_REG_RX_DEF_SEL1: string  := "25uA";
        PMA_REG_RX_TERM_SEL: string  := "25uA";
        PMA_REG_TX_DIV_SEL: string  := "25uA";
        PMA_REG_PMA_CHLBUF_SEL: string  := "25uA";
        PMA_REG_LPLL_AMP_SEL: string  := "25uA";
        PMA_REG_LPLL_VCO_SEL: string  := "25uA";
        PMA_REG_LPLL_CHARGE_PUMP_SEL: string  := "25uA";
        PMA_REG_RX_EM_PI_SEL: string  := "50uA";
        PMA_REG_RX_EM_PI_BUF: string  := "50uA";
        PMA_REG_RX_POI_SEL: string  := "50uA";
        PMA_REG_RX_POI_BUF_SEL: string  := "50uA";
        PMA_REG_RX_PT1_SEL: string  := "50uA";
        PMA_REG_RX_PT1_BUF_SEL: string  := "50uA";
        PMA_REG_RX_EQ0_SEL: string  := "50uA";
        PMA_REG_RX_EQ1_SEL: string  := "50uA";
        PMA_REG_RX_PGA_SEL: string  := "50uA";
        PMA_REG_RX_LSPD_SEL: string  := "50uA";
        PMA_REG_RX_JTAG_VTH_SEL: string  := "50uA";
        PMA_REG_RX_SIGDE_TTH_SEL: string  := "50uA";
        PMA_REG_RX_SIGDET_SEL: string  := "50uA";
        PMA_REG_TX_DET_SEL: string  := "50uA";
        PMA_REG_TX_PI_SEL: string  := "50uA";
        PMA_REG_TX_PI_BUF_SEL: string  := "50uA";
        PMA_REG_CHL_BIAS_SEL: string  := "50uA";
        PMA_REG_CHL_TEST: integer := 0
    );
    port(
        P_CFG_READY     : out    vl_logic;
        P_CFG_RDATA     : out    vl_logic_vector(7 downto 0);
        P_CFG_INT       : out    vl_logic;
        LANE_COUT_BUS_FORWARD: out    vl_logic_vector(25 downto 0);
        P_APATTERN_STATUS_COUT: out    vl_logic;
        P_RX_PRBS_ERROR : out    vl_logic;
        P_PCS_RX_MCB_STATUS: out    vl_logic;
        P_PCS_LSM_SYNCED: out    vl_logic;
        P_RDATA         : out    vl_logic_vector(87 downto 0);
        P_RXDVLD        : out    vl_logic;
        P_RXDVLD_H      : out    vl_logic;
        P_RXSTATUS      : out    vl_logic_vector(5 downto 0);
        P_EM_ERROR_CNT  : out    vl_logic_vector(2 downto 0);
        P_LPLL_READY    : out    vl_logic;
        P_RX_SIGDET_STATUS: out    vl_logic;
        P_RX_SATA_COMINIT: out    vl_logic;
        P_RX_SATA_COMWAKE: out    vl_logic;
        P_RX_LS_DATA    : out    vl_logic;
        P_RX_READY      : out    vl_logic;
        P_TEST_STATUS   : out    vl_logic_vector(19 downto 0);
        P_TX_RXDET_STATUS: out    vl_logic;
        P_RCLK2FABRIC   : out    vl_logic;
        P_TCLK2FABRIC   : out    vl_logic;
        P_CA_ALIGN_RX   : out    vl_logic;
        P_CA_ALIGN_TX   : out    vl_logic;
        P_TX_SDN        : out    vl_logic;
        P_TX_SDP        : out    vl_logic;
        P_TEST_SO0      : out    vl_logic;
        P_TEST_SO1      : out    vl_logic;
        P_TEST_SO2      : out    vl_logic;
        P_TEST_SO3      : out    vl_logic;
        P_TEST_SO4      : out    vl_logic;
        P_FOR_PMA_TEST_SO: out    vl_logic_vector(1 downto 0);
        P_TEST_SE_N     : in     vl_logic;
        P_TEST_MODE_N   : in     vl_logic;
        P_TEST_RSTN     : in     vl_logic;
        P_TEST_SI0      : in     vl_logic;
        P_TEST_SI1      : in     vl_logic;
        P_TEST_SI2      : in     vl_logic;
        P_TEST_SI3      : in     vl_logic;
        P_TEST_SI4      : in     vl_logic;
        P_FOR_PMA_TEST_MODE_N: in     vl_logic;
        P_FOR_PMA_TEST_SE_N: in     vl_logic_vector(1 downto 0);
        P_FOR_PMA_TEST_CLK: in     vl_logic_vector(1 downto 0);
        P_FOR_PMA_TEST_RSTN: in     vl_logic_vector(1 downto 0);
        P_FOR_PMA_TEST_SI: in     vl_logic_vector(1 downto 0);
        P_RX_CLK_FR_CORE: in     vl_logic;
        P_RCLK2_FR_CORE : in     vl_logic;
        P_TX_CLK_FR_CORE: in     vl_logic;
        P_TCLK2_FR_CORE : in     vl_logic;
        P_PCS_RX_RST    : in     vl_logic;
        P_PCS_TX_RST    : in     vl_logic;
        P_EXT_BRIDGE_PCS_RST: in     vl_logic;
        P_CFG_RST       : in     vl_logic;
        P_CFG_CLK       : in     vl_logic;
        P_CFG_PSEL      : in     vl_logic;
        P_CFG_ENABLE    : in     vl_logic;
        P_CFG_WRITE     : in     vl_logic;
        P_CFG_ADDR      : in     vl_logic_vector(11 downto 0);
        P_CFG_WDATA     : in     vl_logic_vector(7 downto 0);
        LANE_CIN_BUS_FORWARD: in     vl_logic_vector(25 downto 0);
        P_APATTERN_STATUS_CIN: in     vl_logic;
        P_TDATA         : in     vl_logic_vector(87 downto 0);
        P_PCIE_EI_H     : in     vl_logic;
        P_PCIE_EI_L     : in     vl_logic;
        P_TX_DEEMP      : in     vl_logic_vector(15 downto 0);
        P_TX_DEEMP_POST_SEL: in     vl_logic_vector(1 downto 0);
        P_BLK_ALIGN_CTRL: in     vl_logic;
        P_TX_ENC_TYPE   : in     vl_logic;
        P_RX_DEC_TYPE   : in     vl_logic;
        P_PCS_BIT_SLIP  : in     vl_logic;
        P_PCS_WORD_ALIGN_EN: in     vl_logic;
        P_RX_POLARITY_INVERT: in     vl_logic;
        P_PCS_MCB_EXT_EN: in     vl_logic;
        P_PCS_NEAREND_LOOP: in     vl_logic;
        P_PCS_FAREND_LOOP: in     vl_logic;
        P_PMA_NEAREND_PLOOP: in     vl_logic;
        P_PMA_NEAREND_SLOOP: in     vl_logic;
        P_PMA_FAREND_PLOOP: in     vl_logic;
        P_PCS_PRBS_EN   : in     vl_logic;
        P_LANE_POWERDOWN: in     vl_logic;
        P_LANE_RST      : in     vl_logic;
        P_RX_LANE_POWERDOWN: in     vl_logic;
        P_RX_PMA_RST    : in     vl_logic;
        P_RX_CDR_RST    : in     vl_logic;
        P_RX_CLKPATH_RST: in     vl_logic;
        P_RX_DFE_RST    : in     vl_logic;
        P_RX_LPM_RST    : in     vl_logic;
        P_RX_SLIDING_RST: in     vl_logic;
        P_RX_DFE_EN     : in     vl_logic;
        P_RX_T1_EN      : in     vl_logic;
        P_RX_CDRX_EN    : in     vl_logic;
        P_RX_T1_DFE_EN  : in     vl_logic;
        P_RX_T2_DFE_EN  : in     vl_logic;
        P_RX_T3_DFE_EN  : in     vl_logic;
        P_RX_T4_DFE_EN  : in     vl_logic;
        P_RX_T5_DFE_EN  : in     vl_logic;
        P_RX_T6_DFE_EN  : in     vl_logic;
        P_RX_SLIDING_EN : in     vl_logic;
        P_RX_EYE_RST    : in     vl_logic;
        P_RX_EYE_EN     : in     vl_logic;
        P_RX_EYE_TAP    : in     vl_logic_vector(7 downto 0);
        P_RX_PIC_EYE    : in     vl_logic_vector(7 downto 0);
        P_RX_PIC_FASTLOCK: in     vl_logic_vector(7 downto 0);
        P_RX_PIC_FASTLOCK_STROBE: in     vl_logic;
        P_EM_RD_TRIGGER : in     vl_logic;
        P_EM_MODE_CTRL  : in     vl_logic_vector(1 downto 0);
        P_RX_CTLE_DCCAL_RST: in     vl_logic;
        P_RX_SLICER_DCCAL_RST: in     vl_logic;
        P_RX_SLICER_DCCAL_EN: in     vl_logic;
        P_RX_CTLE_DCCAL_EN: in     vl_logic;
        P_RX_SLIP_RST   : in     vl_logic;
        P_RX_SLIP_EN    : in     vl_logic;
        P_LPLL_POWERDOWN: in     vl_logic;
        P_LPLL_RST      : in     vl_logic;
        P_LPLL_LOCKDET_RST: in     vl_logic;
        P_TX_LS_DATA    : in     vl_logic;
        P_TX_BEACON_EN  : in     vl_logic;
        P_TX_SWING      : in     vl_logic;
        P_TX_RXDET_REQ  : in     vl_logic;
        P_TX_RATE       : in     vl_logic_vector(1 downto 0);
        P_TX_BUSWIDTH   : in     vl_logic_vector(2 downto 0);
        P_TX_FREERUN_BUSWIDTH: in     vl_logic_vector(2 downto 0);
        P_TX_MARGIN     : in     vl_logic_vector(2 downto 0);
        P_TX_PMA_RST    : in     vl_logic;
        P_TX_LANE_POWERDOWN: in     vl_logic;
        P_TX_PIC_EN     : in     vl_logic;
        P_RX_RATE       : in     vl_logic_vector(1 downto 0);
        P_RX_BUSWIDTH   : in     vl_logic_vector(2 downto 0);
        P_RX_HIGHZ      : in     vl_logic;
        P_CIM_CLK_ALIGNER_RX: in     vl_logic_vector(7 downto 0);
        P_CIM_CLK_ALIGNER_TX: in     vl_logic_vector(7 downto 0);
        P_ALIGN_MODE_VALID_RX: in     vl_logic;
        P_ALIGN_MODE_RX : in     vl_logic_vector(1 downto 0);
        P_ALIGN_MODE_VALID_TX: in     vl_logic;
        P_ALIGN_MODE_TX : in     vl_logic_vector(2 downto 0);
        PMA_HPLL_CK0    : in     vl_logic;
        PMA_HPLL_CK90   : in     vl_logic;
        PMA_HPLL_CK180  : in     vl_logic;
        PMA_HPLL_CK270  : in     vl_logic;
        PMA_HPLL_READY_IN: in     vl_logic;
        PMA_HPLL_REFCLK_IN: in     vl_logic;
        PMA_IPN50U_IN   : in     vl_logic_vector(1 downto 0);
        PMA_LPLL_REFCLK : in     vl_logic;
        PMA_RES_CAL_I   : in     vl_logic_vector(5 downto 0);
        PMA_TX_SYNC_HPLL: in     vl_logic;
        PMA_TX_RATE_CHANGE_ON_0: in     vl_logic;
        PMA_TX_RATE_CHANGE_ON_1: in     vl_logic;
        PMA_TX_SYNC     : in     vl_logic;
        P_RX_SDN        : in     vl_logic;
        P_RX_SDP        : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of PCS_DYN_DLY_SEL_RX : constant is 1;
    attribute mti_svvh_generic_type of PCS_PMA_RCLK_POLINV : constant is 1;
    attribute mti_svvh_generic_type of PCS_PCS_RCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_GEAR_RCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_RCLK2FABRIC_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_SCAN_INTERVAL_RX : constant is 1;
    attribute mti_svvh_generic_type of PCS_BRIDGE_RCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_RCLK_POLINV : constant is 1;
    attribute mti_svvh_generic_type of PCS_TO_FABRIC_CLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CLK2ALIGNER_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_TO_FABRIC_CLK_DIV_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_AUTO_NEAR_LOOP_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_PCS_RCLK_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_BRIDGE_PCS_RCLK_EN_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_BRIDGE_RCLK_EN_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_GEAR_RCLK_EN_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_NEGEDGE_EN_RX : constant is 1;
    attribute mti_svvh_generic_type of PCS_PCS_RX_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PCS_BRIDGE_PCS_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PCS_TO_FABRIC_RST_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_BYPASS_GEAR_RRSTN : constant is 1;
    attribute mti_svvh_generic_type of PCS_BYPASS_BRIDGE_RRSTN : constant is 1;
    attribute mti_svvh_generic_type of PCS_ALIGNER_EN_RX : constant is 1;
    attribute mti_svvh_generic_type of PCS_RX_SLAVE : constant is 1;
    attribute mti_svvh_generic_type of PCS_RX_CA : constant is 2;
    attribute mti_svvh_generic_type of PCS_SUM_THRESHOLD_RX : constant is 2;
    attribute mti_svvh_generic_type of PCS_AVG_CYCLES_RX : constant is 2;
    attribute mti_svvh_generic_type of PCS_REG_PMA_RX2TX_PLOOP_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_REG_PMA_RX2TX_PLOOP_FIFOEN : constant is 1;
    attribute mti_svvh_generic_type of PCS_STEP_SIZE_RX : constant is 2;
    attribute mti_svvh_generic_type of PCS_REV_CNT_LIMIT_RX : constant is 2;
    attribute mti_svvh_generic_type of PCS_FILTER_CNT_SIZE_RX : constant is 2;
    attribute mti_svvh_generic_type of PCS_DLY_ADJUST_SIZE_RX_3_0 : constant is 2;
    attribute mti_svvh_generic_type of PCS_DLY_REC_SIZE_RX : constant is 2;
    attribute mti_svvh_generic_type of PCS_ALIGN_THRD_RX : constant is 2;
    attribute mti_svvh_generic_type of PCS_DLY_ADJUST_SIZE_RX_4 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CFG_DEC_TYPE_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_RXBRIDGE_GEAR_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_GE_AUTO_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_RXBRG_FULL_CHK_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_RXBRG_EMPTY_CHK_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_IFG_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_FLP_FULL_CHK_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_FLP_EMPTY_CHK_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_RX_POLARITY_INV : constant is 1;
    attribute mti_svvh_generic_type of PCS_FARLP_PWR_REDUCTION : constant is 1;
    attribute mti_svvh_generic_type of PCS_RXPRBS_PWR_REDUCTION : constant is 1;
    attribute mti_svvh_generic_type of PCS_WDALIGN_PWR_REDUCTION : constant is 1;
    attribute mti_svvh_generic_type of PCS_RXDEC_PWR_REDUCTION : constant is 1;
    attribute mti_svvh_generic_type of PCS_RXBRG_PWR_REDUCTION : constant is 1;
    attribute mti_svvh_generic_type of PCS_RXTEST_PWR_REDUCTION : constant is 1;
    attribute mti_svvh_generic_type of PCS_WA_SOS_DET_TOL : constant is 2;
    attribute mti_svvh_generic_type of PCS_WA_SE_DET_TOL : constant is 2;
    attribute mti_svvh_generic_type of PCS_RX_SAMPLE_UNION : constant is 1;
    attribute mti_svvh_generic_type of PCS_NEAR_LOOP : constant is 1;
    attribute mti_svvh_generic_type of PCS_BYPASS_WORD_ALIGN : constant is 1;
    attribute mti_svvh_generic_type of PCS_BYPASS_DENC : constant is 1;
    attribute mti_svvh_generic_type of PCS_RX_ERRCNT_CLR : constant is 1;
    attribute mti_svvh_generic_type of PCS_RX_CODE_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_RX_BYPASS_GEAR : constant is 1;
    attribute mti_svvh_generic_type of PCS_ERRDETECT_SILENCE : constant is 1;
    attribute mti_svvh_generic_type of PCS_RX_DATA_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CA_DYN_CLY_EN_RX : constant is 1;
    attribute mti_svvh_generic_type of PCS_CFG_APATTERN_STATUS_DELAY : constant is 1;
    attribute mti_svvh_generic_type of PCS_RX_PRBS_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_ALIGN_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_COMMA_DET_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_RAPID_VMIN_1 : constant is 2;
    attribute mti_svvh_generic_type of PCS_RAPID_VMIN_2 : constant is 2;
    attribute mti_svvh_generic_type of PCS_RXBU_WIDER_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_RAPID_IMAX : constant is 2;
    attribute mti_svvh_generic_type of PCS_RX_SPLIT : constant is 1;
    attribute mti_svvh_generic_type of PCS_RXBRG_END_PACKET_9_8 : constant is 2;
    attribute mti_svvh_generic_type of PCS_RXBRG_END_PACKET_7_0 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CTC_MAX_DEL : constant is 2;
    attribute mti_svvh_generic_type of PCS_COMMA_REG0_9_8 : constant is 2;
    attribute mti_svvh_generic_type of PCS_COMMA_REG1_9_8 : constant is 2;
    attribute mti_svvh_generic_type of PCS_COMMA_MASK_9_8 : constant is 2;
    attribute mti_svvh_generic_type of PCS_COMMA_REG0_7_0 : constant is 2;
    attribute mti_svvh_generic_type of PCS_COMMA_REG1_7_0 : constant is 2;
    attribute mti_svvh_generic_type of PCS_COMMA_MASK_7_0 : constant is 2;
    attribute mti_svvh_generic_type of PCS_FLP_WRADDR_START : constant is 2;
    attribute mti_svvh_generic_type of PCS_FLP_RDADDR_START : constant is 2;
    attribute mti_svvh_generic_type of PCS_CFG_RX_BRIDGE_CLK_POLINV : constant is 1;
    attribute mti_svvh_generic_type of PCS_CTC_MODE_RD_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CTC_AFULL : constant is 2;
    attribute mti_svvh_generic_type of PCS_FAST_LOCK_GEAR_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CTC_MODE_WR_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CTC_AEMPTY : constant is 2;
    attribute mti_svvh_generic_type of PCS_CTC_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_RXBRIDGE_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CTC_ADD_MAX : constant is 2;
    attribute mti_svvh_generic_type of PCS_CFG_PHDET_EN_RX : constant is 1;
    attribute mti_svvh_generic_type of PCS_WA_SDS_DET_TOL : constant is 2;
    attribute mti_svvh_generic_type of PCS_CEB_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_APATTERN_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_A_REG0_8 : constant is 1;
    attribute mti_svvh_generic_type of PCS_RXBRG_WADDR_START : constant is 2;
    attribute mti_svvh_generic_type of PCS_A_REG1_8 : constant is 1;
    attribute mti_svvh_generic_type of PCS_RXBRG_RADDR_START : constant is 2;
    attribute mti_svvh_generic_type of PCS_A_REG0_7_0 : constant is 2;
    attribute mti_svvh_generic_type of PCS_A_REG1_7_0 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CEB_RAPIDLS_MMAX : constant is 2;
    attribute mti_svvh_generic_type of PCS_CEB_DETECT_TIME : constant is 2;
    attribute mti_svvh_generic_type of PCS_WL_FIFO_RD : constant is 2;
    attribute mti_svvh_generic_type of PCS_SKIP_REG0_9_8 : constant is 2;
    attribute mti_svvh_generic_type of PCS_SKIP_REG0_7_0 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CFG_CONTI_SKP_SET : constant is 2;
    attribute mti_svvh_generic_type of PCS_CFG_RX_BASE_ADV_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_SKIP_REG1_9_8 : constant is 2;
    attribute mti_svvh_generic_type of PCS_SKIP_REG2_9_8 : constant is 2;
    attribute mti_svvh_generic_type of PCS_SKIP_REG3_9_8 : constant is 2;
    attribute mti_svvh_generic_type of PCS_SKIP_REG1_7_0 : constant is 2;
    attribute mti_svvh_generic_type of PCS_SKIP_REG2_7_0 : constant is 2;
    attribute mti_svvh_generic_type of PCS_SKIP_REG3_7_0 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CFG_PRBS_ERR_O_SEL : constant is 2;
    attribute mti_svvh_generic_type of PCS_CFG_PD_DELAY_RX : constant is 2;
    attribute mti_svvh_generic_type of PCS_WR_START_GAP : constant is 2;
    attribute mti_svvh_generic_type of PCS_MIN_IFG : constant is 2;
    attribute mti_svvh_generic_type of PCS_INT_RX_MASK_0 : constant is 1;
    attribute mti_svvh_generic_type of PCS_INT_RX_MASK_1 : constant is 1;
    attribute mti_svvh_generic_type of PCS_INT_RX_MASK_2 : constant is 1;
    attribute mti_svvh_generic_type of PCS_INT_RX_MASK_3 : constant is 1;
    attribute mti_svvh_generic_type of PCS_INT_RX_MASK_4 : constant is 1;
    attribute mti_svvh_generic_type of PCS_INT_RX_MASK_5 : constant is 1;
    attribute mti_svvh_generic_type of PCS_INT_RX_CLR_5 : constant is 1;
    attribute mti_svvh_generic_type of PCS_INT_RX_CLR_4 : constant is 1;
    attribute mti_svvh_generic_type of PCS_INT_RX_CLR_3 : constant is 1;
    attribute mti_svvh_generic_type of PCS_INT_RX_CLR_2 : constant is 1;
    attribute mti_svvh_generic_type of PCS_INT_RX_CLR_1 : constant is 1;
    attribute mti_svvh_generic_type of PCS_INT_RX_CLR_0 : constant is 1;
    attribute mti_svvh_generic_type of PCS_EM_CNT_RD_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_EM_CTRL_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_EM_MODE_CTRL : constant is 1;
    attribute mti_svvh_generic_type of PCS_EM_RD_CONDITION : constant is 1;
    attribute mti_svvh_generic_type of PCS_EM_SP_PATTERN_7_0 : constant is 2;
    attribute mti_svvh_generic_type of PCS_EM_SP_PATTERN_15_8 : constant is 2;
    attribute mti_svvh_generic_type of PCS_EM_SP_PATTERN_23_16 : constant is 2;
    attribute mti_svvh_generic_type of PCS_EM_SP_PATTERN_31_24 : constant is 2;
    attribute mti_svvh_generic_type of PCS_EM_SP_PATTERN_39_32 : constant is 2;
    attribute mti_svvh_generic_type of PCS_EM_SP_PATTERN_47_40 : constant is 2;
    attribute mti_svvh_generic_type of PCS_EM_SP_PATTERN_55_48 : constant is 2;
    attribute mti_svvh_generic_type of PCS_EM_SP_PATTERN_63_56 : constant is 2;
    attribute mti_svvh_generic_type of PCS_EM_SP_PATTERN_71_64 : constant is 2;
    attribute mti_svvh_generic_type of PCS_EM_SP_PATTERN_79_72 : constant is 2;
    attribute mti_svvh_generic_type of PCS_EM_PMA_MASK_7_0 : constant is 2;
    attribute mti_svvh_generic_type of PCS_EM_PMA_MASK_15_8 : constant is 2;
    attribute mti_svvh_generic_type of PCS_EM_PMA_MASK_23_16 : constant is 2;
    attribute mti_svvh_generic_type of PCS_EM_PMA_MASK_31_24 : constant is 2;
    attribute mti_svvh_generic_type of PCS_EM_PMA_MASK_39_32 : constant is 2;
    attribute mti_svvh_generic_type of PCS_EM_PMA_MASK_47_40 : constant is 2;
    attribute mti_svvh_generic_type of PCS_EM_PMA_MASK_55_48 : constant is 2;
    attribute mti_svvh_generic_type of PCS_EM_PMA_MASK_63_56 : constant is 2;
    attribute mti_svvh_generic_type of PCS_EM_PMA_MASK_71_64 : constant is 2;
    attribute mti_svvh_generic_type of PCS_EM_PMA_MASK_79_72 : constant is 2;
    attribute mti_svvh_generic_type of PCS_EM_EYED_MASK_7_0 : constant is 2;
    attribute mti_svvh_generic_type of PCS_EM_EYED_MASK_15_8 : constant is 2;
    attribute mti_svvh_generic_type of PCS_EM_EYED_MASK_23_16 : constant is 2;
    attribute mti_svvh_generic_type of PCS_EM_EYED_MASK_31_24 : constant is 2;
    attribute mti_svvh_generic_type of PCS_EM_EYED_MASK_39_32 : constant is 2;
    attribute mti_svvh_generic_type of PCS_EM_EYED_MASK_47_40 : constant is 2;
    attribute mti_svvh_generic_type of PCS_EM_EYED_MASK_55_48 : constant is 2;
    attribute mti_svvh_generic_type of PCS_EM_EYED_MASK_63_56 : constant is 2;
    attribute mti_svvh_generic_type of PCS_EM_EYED_MASK_71_64 : constant is 2;
    attribute mti_svvh_generic_type of PCS_EM_EYED_MASK_79_72 : constant is 2;
    attribute mti_svvh_generic_type of PCS_EM_PRESCALE : constant is 2;
    attribute mti_svvh_generic_type of PCS_CFG_TEST_STATUS_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CFG_DIFF_CNT_BND_RX : constant is 2;
    attribute mti_svvh_generic_type of PCS_CFG_FLT_SEL_RX : constant is 1;
    attribute mti_svvh_generic_type of PCS_FILTER_BND_RX : constant is 2;
    attribute mti_svvh_generic_type of PCS_TCLK2FABRIC_DIV_RST_M : constant is 1;
    attribute mti_svvh_generic_type of PCS_TX_PMA_TCLK_POLINV : constant is 1;
    attribute mti_svvh_generic_type of PCS_TX_TCLK_POLINV : constant is 1;
    attribute mti_svvh_generic_type of PCS_PCS_TCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_GEAR_TCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_TX_BRIDGE_TCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_TCLK2ALIGNER_SEL : constant is 1;
    attribute mti_svvh_generic_type of CA_DYN_DLY_EN_TX : constant is 1;
    attribute mti_svvh_generic_type of PCS_TX_PCS_CLK_EN_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_TX_GEAR_CLK_EN_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_TCLK2FABRIC_DIV_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_TCLK2FABRIC_SEL : constant is 1;
    attribute mti_svvh_generic_type of DLY_ADJUST_SIZE_TX : constant is 2;
    attribute mti_svvh_generic_type of PCS_TX_PCS_TX_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PCS_TX_CA_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PCS_TX_SLAVE : constant is 1;
    attribute mti_svvh_generic_type of PCS_TX_CA : constant is 2;
    attribute mti_svvh_generic_type of PCS_CFG_PI_CLK_SEL : constant is 2;
    attribute mti_svvh_generic_type of PCS_CFG_PI_CLK_EN_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CFG_PI_STEP_SIZE_TX : constant is 2;
    attribute mti_svvh_generic_type of PCS_CFG_SUM_THRESHOLD_TX : constant is 2;
    attribute mti_svvh_generic_type of PCS_CFG_AVG_CYCLES_TX : constant is 2;
    attribute mti_svvh_generic_type of PCS_CFG_NEGEDGE_EN_TX : constant is 1;
    attribute mti_svvh_generic_type of PCS_CFG_ALIGN_THRD_TX : constant is 2;
    attribute mti_svvh_generic_type of PCS_CFG_SCAN_INTERVAL_TX : constant is 2;
    attribute mti_svvh_generic_type of PCS_CFG_STEP_SIZE_TX : constant is 2;
    attribute mti_svvh_generic_type of PCS_CFG_REV_CNT_LIMIT_TX : constant is 2;
    attribute mti_svvh_generic_type of PCS_CFG_FILTER_CNT_SIZE_TX : constant is 2;
    attribute mti_svvh_generic_type of PCS_CFG_PI_DEFAULT_TX : constant is 2;
    attribute mti_svvh_generic_type of PCS_CFG_PHDET_EN_TX : constant is 1;
    attribute mti_svvh_generic_type of PCS_PMA_TX2RX_PLOOP_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_PMA_TX2RX_SLOOP_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CFG_DYN_DLY_SEL_TX : constant is 1;
    attribute mti_svvh_generic_type of PCS_CFG_DLY_REC_SIZE_TX : constant is 2;
    attribute mti_svvh_generic_type of PCS_TX_DATA_WIDTH_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_TX_BYPASS_BRIDGE_UINT : constant is 1;
    attribute mti_svvh_generic_type of PCS_TX_BYPASS_BRIDGE_FIFO : constant is 1;
    attribute mti_svvh_generic_type of PCS_TX_BYPASS_GEAR : constant is 1;
    attribute mti_svvh_generic_type of PCS_TX_BYPASS_ENC : constant is 1;
    attribute mti_svvh_generic_type of PCS_TX_BYPASS_BIT_SLIP : constant is 1;
    attribute mti_svvh_generic_type of PCS_TX_BRIDGE_GEAR_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_TXBRG_PWR_REDUCTION : constant is 1;
    attribute mti_svvh_generic_type of PCS_TXGEAR_PWR_REDUCTION : constant is 1;
    attribute mti_svvh_generic_type of PCS_TXENC_PWR_REDUCTION : constant is 1;
    attribute mti_svvh_generic_type of PCS_TXBSLP_PWR_REDUCTION : constant is 1;
    attribute mti_svvh_generic_type of PCS_TXPRBS_PWR_REDUCTION : constant is 1;
    attribute mti_svvh_generic_type of PCS_TXBRG_FULL_CHK_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_TXBRG_EMPTY_CHK_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_TX_ENCODER_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_TX_PRBS_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_TX_DRIVE_REG_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_TX_BIT_SLIP_CYCLES : constant is 2;
    attribute mti_svvh_generic_type of PCS_TX_BASE_ADV_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_TX_GEAR_SPLIT : constant is 1;
    attribute mti_svvh_generic_type of PCS_RX_BRIDGE_CLK_POLINV : constant is 1;
    attribute mti_svvh_generic_type of PCS_PRBS_ERR_LPBK : constant is 1;
    attribute mti_svvh_generic_type of PCS_TX_INSERT_ER : constant is 1;
    attribute mti_svvh_generic_type of PCS_ENABLE_PRBS_GEN : constant is 1;
    attribute mti_svvh_generic_type of PCS_FAR_LOOP : constant is 1;
    attribute mti_svvh_generic_type of PCS_CFG_ENC_TYPE_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_TXBRG_WADDR_START : constant is 2;
    attribute mti_svvh_generic_type of PCS_TXBRG_RADDR_START : constant is 2;
    attribute mti_svvh_generic_type of PCS_CFG_TX_PIC_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CFG_PIC_DIRECT_INV : constant is 1;
    attribute mti_svvh_generic_type of PCS_CFG_PI_MOD_CLK_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CFG_TX_MODULATOR_OW_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CFG_TX_PI_SSC_MODE_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CFG_TX_PI_OFFSET_MODE_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CFG_TX_PI_SSC_MODE_SEL : constant is 2;
    attribute mti_svvh_generic_type of PCS_CFG_TXDEEMPH_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_PI_STROBE_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CFG_TX_PIC_GREY_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CFG_PIC_RENEW_INV : constant is 1;
    attribute mti_svvh_generic_type of PCS_CFG_NUM_PIC : constant is 2;
    attribute mti_svvh_generic_type of PCS_CFG_TXPIC_OW_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CFG_TXPPM_OW_VALUE_0_7 : constant is 2;
    attribute mti_svvh_generic_type of PCS_INT_TX_MASK_0 : constant is 1;
    attribute mti_svvh_generic_type of PCS_INT_TX_MASK_1 : constant is 1;
    attribute mti_svvh_generic_type of PCS_INT_TX_MASK_2 : constant is 1;
    attribute mti_svvh_generic_type of PCS_INT_TX_CLR_2 : constant is 1;
    attribute mti_svvh_generic_type of PCS_INT_TX_CLR_1 : constant is 1;
    attribute mti_svvh_generic_type of PCS_INT_TX_CLR_0 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CFG_PD_DELAY_TX : constant is 2;
    attribute mti_svvh_generic_type of PCS_CFG_DIFF_CNT_BND_TX : constant is 2;
    attribute mti_svvh_generic_type of PCS_CFG_PD_CLK_FR_CORE_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CFG_FLT_SEL_TX : constant is 1;
    attribute mti_svvh_generic_type of PCS_FILTER_BND_TX : constant is 2;
    attribute mti_svvh_generic_type of PCS_CFG_TX_SSC_PPM_RANGE_7_0 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CFG_TX_PPM_MODULATOR_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CFG_TX_PPM_SCALE2_SEL : constant is 2;
    attribute mti_svvh_generic_type of PCS_CFG_TX_PPM_SCALE_SEL : constant is 2;
    attribute mti_svvh_generic_type of PCS_CFG_TX_SSC_PPM_RANGE_8_9 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CFG_TX_SSC_MODULATION_STEP_7_0 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CFG_TX_SSC_PPM_OFFSET_7_0 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CFG_TX_SSC_MODULATION_STEP_8 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CFG_TX_SSC_PPM_OFFSET_8_9 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_CHL_BIAS_POWER_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_CHL_BIAS_POWER : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_BUSWIDTH : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_RATE : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_RATE_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_RES_TRIM : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RX_SIGDET_STATUS_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_CDR_READY_THD_7_0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_CDR_READY_THD_11_8 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RX_BUSWIDTH_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_PCLK_EDGE_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_CDR_READY_CHECK_CTRL : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RX_ICTRL_TRX : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_PRBS_CHK_WIDTH_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RX_ICTRL_PIBUF : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_ICTRL_PI : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_ICTRL_DCC : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_TX2RX_PLPBK_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_DATA_POLARITY : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_ERR_INSERT : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_UDP_CHK_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_PRBS_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_PRBS_CHK_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_LPLL_NFC_STIC_DIS_N : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_BIST_CHK_PAT_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_LOAD_ERR_CNT : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_CHK_COUNTER_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_CDR_PROP_GAN_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_CDR_TUBO_PROP_GAIN_SEL : constant is 2;
    attribute mti_svvh_generic_type of PAM_REG_CDR_INT_GAIN_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_CDR_TUBO_INT_GAIN_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_CDR_INT_SAT_MAX_4_0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_CDR_INT_SAT_MAX_9_5 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_CDR_INT_SAT_MIN_2_0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_CDR_INT_SAT_MIN_9_3 : constant is 2;
    attribute mti_svvh_generic_type of PMA_ANA_RX_REG_O_61_55 : constant is 2;
    attribute mti_svvh_generic_type of PMA_ANA_RX_REG_O_69_62 : constant is 2;
    attribute mti_svvh_generic_type of PMA_ANA_RX_REG_O_77_70 : constant is 2;
    attribute mti_svvh_generic_type of PMA_ANA_RX_REG_O_85_78 : constant is 2;
    attribute mti_svvh_generic_type of PMA_ANA_RX_REG_O_93_86 : constant is 2;
    attribute mti_svvh_generic_type of PMA_ANA_RX_REG_O_100_94 : constant is 2;
    attribute mti_svvh_generic_type of PMA_ANA_RX_REG_O_108_101 : constant is 2;
    attribute mti_svvh_generic_type of PMA_ANA_RX_REG_O_111_109 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_OOB_COMWAKE_GAP_MIN_4_0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_OOB_COMWAKE_GAP_MIN_5 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_OOB_COMWAKE_GAP_MAX : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_OOB_COMINIT_GAP_MIN : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_OOB_COMINIT_GAP_MAX : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_COMWAKE_STATUS_CLEAR : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_COMINIT_STATUS_CLEAR : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RX_SATA_COMINIT_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_SATA_COMINIT : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_SATA_COMWAKE_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_SATA_COMWAKE : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_DCC_DISABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_SLIP_SEL_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_SLIP_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RX_SLIP_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_SIGDET_STATUS_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RX_SIGDET_FSM_RST_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_SIGDET_STATUS : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_SIGDET_VTH : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_SIGDET_GRM : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RX_SIGDET_PULSE_EXT : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_SIGDET_CH2_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RX_SIGDET_CH2_CHK_WINDOW : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RX_SIGDET_CHK_WINDOW_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_SIGDET_NOSIG_COUNT_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RX_SIGDET_OOB_DET_COUNT_VAL_2_0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RX_SIGDET_OOB_DET_COUNT_VAL_4_3 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RX_SIGDET_4OOB_DET_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RX_SIGDET_IC_I : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RX_EQ1_R_SET_TOP : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RX_EQ1_C_SET_FB : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RX_EQ1_OFF : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_EQ2_R_SET_TOP : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RX_EQ2_C_SET_FB : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RX_EQ2_OFF : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_ICTRL_EQ : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_EQ_DC_CALIB_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CTLE_CTRL_REG_I : constant is 2;
    attribute mti_svvh_generic_type of PMA_CTLE_REG_FORCE_SEL_I : constant is 1;
    attribute mti_svvh_generic_type of PMA_CTLE_REG_HOLD_I : constant is 1;
    attribute mti_svvh_generic_type of PMA_CTLE_REG_INIT_DAC_I_1_0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CTLE_REG_INIT_DAC_I_3_2 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CTLE_REG_POLARITY_I : constant is 1;
    attribute mti_svvh_generic_type of PMA_CTLE_REG_SHIFTER_GAIN_I : constant is 2;
    attribute mti_svvh_generic_type of PMA_CTLE_REG_THRESHOLD_I_1_0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CTLE_REG_THRESHOLD_I_9_2 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CTLE_REG_THRESHOLD_I_11_10 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RX_RES_TRIM_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_RX_TERM_POWER_DIVIDING_SELECTION : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_RX_TERM_VCM_SELECTION : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_RX_TERM_TEST_SELECTION_7_0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_RX_TERM_TEST_SELECTION_9_8 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_LOW_SPEED_MODE_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_RX_CLOCK_POWER_DOWN_REGISTER : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_RX_CLOCK_POWER_DOWN_SELECTION : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_RX_DFE_POWER_DOWN_REGISTER_0 : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_RX_DFE_POWER_DOWN_SELECTION_1 : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_RX_CTLE_POWER_DOWN_REGISTER_0 : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_RX_CTLE_POWER_DOWN_SELECTION_1 : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_EYE_DFETAP1_PLORITY : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_CDR_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_EYE_DET_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_PI_BIAS_CURRENT : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_DFE_TEST_SEL_6_0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_DFE_TEST_SEL_14_7 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_DFE_TEST_SEL_21_15 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_CTLE_TEST_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_ANA_RX_SLIP_SEL_O : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_RX_T1_BUFF_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_RX_CDRX_BUFF_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_RX_VP_T1_SW_PLORITY : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_RX_VP_PLORITY : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_RX_GAIN_CTRL_SUMMER : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_RX_DC_OFFSET_T1_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_RX_DC_OFFSET_VP_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_RX_DC_OFFSET_CDRX_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_RX_DC_OFFSET_CDRY_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_RX_DC_OFFSET_EYE_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_SLICER_DC_OFFSET_OVERWITE : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_SLICER_DC_OFFSET_REG : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_SHUT_OFF_THE_EQUALIZER_OF_EACH_STAGE : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_CDR_XWEIGHT_I : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_CDR_YWEIGHT_I : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_CTLE_FLIPDIR_I : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_CTLE_HOLD_I : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_CTLE_INITDAC_5_0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_CTLE_INITDAC_6 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_CTLE_OVERWREN_I : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_CTLE_SHIFT_I : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_CTLE_TOPNUM_2_0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_CTLE_TOPNUM_4_3 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_CTLEOFS_FLIPDIR_I : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_CTLEOFS_HOLD_I : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_CTLEOFS_INITDAC_3_0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_CTLEOFS_INITDAC_6_4 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_CTLEOFS_OVERWREN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_CTLEOFS_SHIFT_I : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_DFE_CTLE_PWD : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_H1_FLIPDIR_I : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_H1_HOLD_I : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_H1_INITDAC_5_0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_H1_INITDAC_6 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_H1_OVERWREN_I : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_H1_SHIFT_I : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_H2_FLIPDIR_I : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_H2_HOLD_I : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_H2_INITDAC_0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_H2_INITDAC_5_1 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_H2_OVERWREN_I : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_H2_SHIFT_I_1_0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_H2_SHIFT_I_2 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_H3_FLIPDIR_I : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_H3_HOLD_I : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_H3_INITDAC_4_0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_H3_INITDAC_5 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_H3_OVERWREN_I : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_H3_SHIFT_I : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_H4_FLIPDIR_I : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_H4_HOLD_I : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_H4_INITDAC_0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_H4_INITDAC_4_1 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_H4_OVERWREN_I : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_H4_SHIFT_I : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_H5_FLIPDIR_I : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_H5_HOLD_I : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_H5_INITDAC : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_H5_OVERWREN_I : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_H5_SHIFT_I : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_H6_FLIPDIR_I : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_H6_HOLD_I : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_H6_INITDAC_2_0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_H6_INITDAC_4_3 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_H6_OVERWREN_I : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_H6_SHIFT_I : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_HCTLE_OFS_1_0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_HCTLE_OFS_3_2 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_HCTLE_OVERWRDAC_5_0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_HCTLE_OVERWRDAC_6 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_HCTLE_OVERWREN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_LPMH_INITDAC_I : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_LPMH_PWD_I : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_LPMH_REG_HOLD_I : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_LPMH_REG_SHIFT_I : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_LPML_INITDAC_I : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_LPML_PWD_I : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_LPML_REG_HOLD_I : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_LPML_REG_PRESELECT_I : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_LPML_REG_SHIFT_I : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_NEXTBIT_I : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_SOFS_COUNTMAX_I_6_0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_SOFS_COUNTMAX_I_14_7 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_SOFS_COUNTMAX_I_19_15 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_SOFS_DACWIN_I : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_SOFS_FLIP_DIR_I : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_SOFS_FORCE_I : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_SOFS_FORCEDAC_I_5_0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_SOFS_FORCEDAC_I_6 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_SOFS_FORCENUM_I : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_SOFS_INITDAC_2_0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_SOFS_INITDAC_6_3 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_SOFS_SHIFT_I : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_SOFS_SKIP_I : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_SOFS_WINCOUNTMAX_I_7_0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_SOFS_WINCOUNTMAX_I_11_8 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_ST_FLIPDIR_I : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_ST_FORCEN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_ST_HOLD_I : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_ST_INITDAC_0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_ST_INITDAC_4_1 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_ST_RECALEN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_ST_SHIFT_I : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_ST_STARTCNT_7_0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_ST_STARTCNT_15_8 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_ST_STARTCNT_19_16 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_ST_TAPCNT_3_0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_ST_TAPCNT_11_4 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_ST_TAPCNT_17_12 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_ST_TOPTAP_1_0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_ST_TOPTAP_3_2 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_SWCLK_DIV : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_TAPA_DAC_3_0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_TAPA_DAC_4 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_TAPA_NUM : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_TAPB_DAC_0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_TAPB_DAC_4_1 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_TAPB_NUM_3_0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_TAPB_NUM_5_4 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_TAPC_DAC : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_TAPC_NUM_0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_TAPC_NUM_5_1 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_TAPD_DAC_2_0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_TAPD_DAC_4_3 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_TAPD_NUM : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_VP_FLIPDIR_I : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_VP_GRN_SHIFT_I : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_VP_HOLD_I : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_VP_IDEAL_2_0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_VP_IDEAL_6_3 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_VP_INITDAC_I_3_0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_VP_INITDAC_I_6_4 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_VP_OVERWREN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_VP_RED_SHIFT_I : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_VPOFS_SEL_0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_VPOFS_SEL_2_1 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_H1_UPBOUND_5_0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_H1_UPBOUND_6 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_CTLEOFS_PWDN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_LPMH_OVEREN_I : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_LPML_OVEREN_I : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_AGC_FLIPDIR_I : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_AGC_HOLD_I : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_AGC_INITDAC : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_AGC_LOWBOUND_1_0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_AGC_LOWBOUND_3_2 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_AGC_OVERWREN_I : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_AGC_PWD : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ALG_AGC_SHIFT_I : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_AGC_UPBOUND_0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_AGC_UPBOUND_3_1 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ALG_AGC_WAITSEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_PI_CTRL_SEL_RX : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_PI_CTRL_RX_4_0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_PI_CTRL_RX_7_5 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CFG_RX_LANE_POWERUP : constant is 1;
    attribute mti_svvh_generic_type of PMA_CFG_RX_PMA_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PMA_INT_PMA_RX_MASK_0 : constant is 1;
    attribute mti_svvh_generic_type of PMA_INT_PMA_RX_CLR_0 : constant is 1;
    attribute mti_svvh_generic_type of PMA_CFG_CTLE_ADP_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CFG_RX_CDR_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CFG_RX_CLKPATH_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CFG_RX_DFE_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CFG_RX_LPM_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CFG_RX_SLIDING_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CFG_RX_EYE_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CFG_RX_CTLE_DCCAL_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CFG_RX_SLICER_DCCAL_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CFG_RX_SLIP_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_PD_MINOR : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_PD_MINOR_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_MAIN_PRE_Z : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_MAIN_PRE_Z_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_BEACON_TIMER_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_RXDET_REQ_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_RXDET_REQ : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_BEACON_EN_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_BEACON_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_EI_EN_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_EI_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_BIT_CONV : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_RES_CAL : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_UDP_DATA_20 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_UDP_DATA_26_21 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_UDP_DATA_34_27 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_UDP_DATA_39_25 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_PD_MAIN : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_PD_MAIN_OW : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_BUSWIDTH_EN : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_SYNC_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_SYNC : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_PD_POST : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_PD_POST_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_RESET_N_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_RESET_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_PMA_TX_RESET_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_PMA_TX_RESET_N_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_BUSWIDTH : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_PLL_READY_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_PLL_READY : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_EI_PCLK_DELAY_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_AMP_DAC0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_AMP_DAC1 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_AMP_DAC2 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_AMP_DAC3 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_MARGIN : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_MARGIN_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_SWING : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_SWING_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_RXDET_THRESHOLD : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_BEACON_OSC_CTRL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_PRBS_GEN_WIDTH_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_TX2RX_SLPBACK_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_PCLK_EDGE_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_RXDET_STATUS_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_RXDET_STATUS : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_PRBS_GEN_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_PRBS_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_UDP_DATA_7_TO_0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_UDP_DATA_15_TO_8 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_UDP_DATA_19_TO_16 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_FIFO_WP_CTRL : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_FIFO_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_DATA_MUX_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_ERR_INSERT : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_SATA_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RATE_CHANGE_TXPCLK_ON_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RATE_CHANGE_TXPCLK_ON : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_CFG_POST1 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_CFG_POST2 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_DEEMP : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_DEEMP_O : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_OOB_DELAY_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_POLARITY : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ANA_TX_JTAG_DATA_O_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_LS_MODE_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_JTAG_MODE_EN_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_JTAG_MODE_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_JTAG_MODE_EN_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_JTAG_MODE_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_JTAG_OE : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_ACJTAG_VHYSTSEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_RES_CAL_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_TERM_MODE_CTRL : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_PLPBK_TXPCLK_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_CLK_SEL_STROBE_TXPCLK : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_PH_SEL_0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_PH_SEL_6_1 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_CFG_PRE : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_CFG_MAIN : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_CFG_POST : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_PD_MAIN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_PD_PRE : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_LS_DATA : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_DCC_BUF_SZ_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_DCC_CAL_CUR_TUNE : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_DCC_CAL_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_DCC_CUR_SS : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_DCC_FA_CTRL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_DCC_RI_CTRL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_ATB_SEL_2_0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_ATB_SEL_9_3 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_CFG_7_0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_CFG_15_8 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_CFG_23_16 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_CFG_31_24 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_OOB_EI_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_OOB_EI_EN_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_BEACON_EN_DELAYED : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_BEACON_EN_DELAYED_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_JTAG_DATA : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_RXDET_TIMER_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_CFG1_7_0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_CFG1_15_8 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_CFG1_23_16 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_CFG1_31_24 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_PI_CUR_BUF : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_ATB_4_0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_ATB_9_5 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_MOD_STAND_BY_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_STATE_STAND_BY_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_PISO_PD : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_PISO_PD_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_CLK_PD : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_CLK_PD_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_DRIVER_PD : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_DRIVER_PD_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_SYNC_NEW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_SYNC_NEW_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_CHANGE_ON_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_CHANGE_ON_POLAR_CTRL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_FREERUN_PD : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_CHANGE_ON_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_CHANGE_ON_CTRL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_PIDC_CURRENT_EN : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_FREERUN_RATE_0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_FREERUN_RATE_1 : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_FREERUN_RATE_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_VBIAS_REG_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_VBIAS_DIVIDER_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_RST_SYNC_CLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_PI_CTRL_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_TX_PI_CTRL : constant is 2;
    attribute mti_svvh_generic_type of PMA_LANE_POWERUP : constant is 1;
    attribute mti_svvh_generic_type of PMA_POR_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_TX_LANE_POWERUP : constant is 1;
    attribute mti_svvh_generic_type of PMA_TX_PMA_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PMA_LPLL_POWERUP : constant is 1;
    attribute mti_svvh_generic_type of PMA_LPLL_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PMA_LPLL_LOCKDET_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_LPLL_PFDDELAY_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_LPLL_PFDDELAY_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_LPLL_VCTRL_SET : constant is 2;
    attribute mti_svvh_generic_type of PMA_LPLL_CHARGE_PUMP_CTRL : constant is 1;
    attribute mti_svvh_generic_type of PMA_LPLL_REFDIV : constant is 1;
    attribute mti_svvh_generic_type of PMA_LPLL_FBDIV : constant is 2;
    attribute mti_svvh_generic_type of PMA_LPLL_LPF_RES : constant is 2;
    attribute mti_svvh_generic_type of PMA_LPLL_TEST_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_LPLL_TEST_SIG_HALF_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_LPLL_TEST_V_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_BUF_BIAS_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TXCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RXCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TEST_BUF : constant is 2;
    attribute mti_svvh_generic_type of PMA_REG_RX_DEF_SEL0 : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_DEF_SEL1 : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_TERM_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_DIV_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_PMA_CHLBUF_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_LPLL_AMP_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_LPLL_VCO_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_LPLL_CHARGE_PUMP_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_EM_PI_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_EM_PI_BUF : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_POI_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_POI_BUF_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_PT1_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_PT1_BUF_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_EQ0_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_EQ1_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_PGA_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_LSPD_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_JTAG_VTH_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_SIGDE_TTH_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_RX_SIGDET_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_DET_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_PI_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_TX_PI_BUF_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_CHL_BIAS_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_REG_CHL_TEST : constant is 2;
end V_HSSTHP_LANE;
