`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
agR/md3W4LC0pk/ThSOjT7cnkN4YyPXQUwsg54K25MW/gTSe6mu1iIp9DGHBjUTk
E2sUlKbRptqPPYq9p/Revd4lqo1/AdEqEqNSTHBhdsVtouWGUxeNvaZ1hL1ny5Yn
lujEnOoN7YnTlTS1lK6NQs/YSciwjdn5LuYCxyPgtpYONbo6wGJrfcB8BJNHkOXJ
4oxt5WOH1PUuewTASyCXoBHaKtpGY7TaTHvbdkl/8Tf96aFvs21hkvE/g9nhbySE
xaJG6dMg0eVPObJ9Pj+MN13RJqa++senTAGtY+BfWgKrplD3Lwve/F7xnAnWTSze
X8Pf9auPisGBDICxesyDFS/wuGUsNkPcRiYDk292SrpmrEESsy9/9phf5qskKLWU
oN/NOi8Zw6NF1AATE/C/jA2wgtzcjIAXBY861lptoTiP8cGXbgVcrh4ikEwkZiYp
R589+P+OCThkthR41wb7kBBNFwqMnsIMSIrnVjqY5eS+5nl76JxDWPvpeVkxsLjG
injkB7Is6rhF0FIVr3o6KoEcmJF/fZTvDOGqktuTVKgEH0w+g/x4TmHVOSKTaxoC
XxVFmXYfd6caFkIktRmIuq6TvvF3ZtgGe9eEdYdA4sZH5loxRtuaOvi+p4C5KLFJ
hkN63FYaWwk9CfSrnYriQm1aiIuSs6TYQbea4SFk3HsFNmfmsg8f52DllZdGwWG2
ADRGW+jg84PrjKFT3Jkg/9cIAkRs+mPsnSHzsaIzL8y8TXzvi+rdLOIUfCYfQbjF
MDXe2C/S+U0ULXjoxDuuhUiUbkb4PlcGE6gQQRciyS4=
`protect END_PROTECTED
