`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sFDmJ55Ow1pE+trUKkTLfwj4Rghus1nX9LO/XGX8Ab7gj36KSaT6u8ynwBEL8LYC
u9TVPmdvPgDvV1LCcS/mke01Z0BJE34O3brIDbiXplmoTEI3DkqXJ1EAKPUn/vbA
RQ9vkB8/0WjJOJYHfVmzMgzWqNAqSUtboe9YBuqlYueOqwVqjUCcWPEZ+2y3dRTj
giMMQI7x/8Bgla4IH8A4E8ZTQxcPNB74n6TDJHyE2YP7eJ1kmUBuFvhF0NJDLzG1
4/HTfiIs9uhxnYEbzzpSDbUgVHQ6+tEd4snXbtsqyDsOb/hpzXPEr7ZSgnIwjkSm
gkh60jwjBLERo7hG4DPrh7aTkc70NafZYyriDPqTcPTr+yhYylaYaY7EJV7DwiJq
IEscUMhr05L88LAyebh1d5YnNXiErWdRIVTjpwAx5Tf/AbHT977U/WDuL4u0sHan
YdPnh8MaUdgcSPRkCotbCmrpmaXPqzzkupGN6WgjU0lZAO5XSLdH187emeKz4DJD
noho2yuXxCfpjDubhSCWW5rp6B2liZ32wMTdEMXSeetDOWuFoBQcZswPvtAQ0y0m
f7y5qDPe4Vmf7e8O3fIQtPEA1NgWtCAj5wx+RsFhuzWbLm9OebayYf5mt6VriVlE
uVj1UEodOrfHNZh9g2ORolF7glg0OCZmZk96dzHVlhgiB5LyN++oX69UquYJVw6b
VhZ+qz20p7Z005YiqKTJl6BlPvycgVAkbcJbXeqP/uyu2I2nt7wfaHY2/gjpkcgX
fZtph5HWVgd2bwkNynjwHDAbC9vZoTJYJUpBt3tG66sFaxerWyco0VjDE00rJKIy
6YMdSxRMQhViqGAm4iC+7HaGfTtAYdqdtwMEhASDTYSxLOSLr8hrPc73TBk4YWm+
FbTmClILQbma5pIPzfoxIU2iZITgCl5PY4GAh6G1KG5U/TysDhBh/7qCJ/dKi+EN
ms+qiAFc1XUe7YEwhHODDNxOvBnUIHW8MlJucRmvengHCTkKM2Yy0EOVvCg3hWlr
F2arCTJ19EUCYVY5clmsHjOCZaLHwwO+MR3oE9xl3nadLhJm5WAhbuGsy5lhyxeL
IPScNob2IxEfsFukJmG1yWzunktbg1CTHQFDvHiVJmASyNT0K+k/BQiDlE6UWSSP
QUcKxx76hLwqGK/df26J1CLwlG98mZXY6teV6Gb1TZOGF4KAiYZed3BpL8bEtURp
ZazeRYOxfJmozdKZPqmWCeOl3fVGLQPZgeTyGW++t854vCxMAFH/dC5iOoqE2bw1
Nq6hbQtmjbOnRUb9ePf4sCBiSW5rAJCZcNVrqsUNPWH4skUIPTYWzFme7yvxaLHC
hT88IP4/YsVXODMn/FH0scu0zzff6/52OCT8QbkGhpDWa2pvi4Av4x3yemkbp/nr
oQ9ksnU/c99Uq6gW52AdSJ9hSRavoDiPR5IOTpx4XRJisgaDH7KhUPrrxrz3Wmwj
MsAbOcHAun0MP6igg4PkAki0BFA5iDp0MKAW1bZaSRf+KKpMavSsQ9VFoUJv0jxY
u2WCoiXtpVRtZuVG/00qN7Mp1l3vzX9oBAldmkdZcdIlWV4ToY+Ex0MSxMPXCv4r
8vkLMdpCMRbq9Wu3pF0s09VyG6+JjrPuwqnA5W5DzSZAN0lpBGG5F4yqgSYeKpn5
MgXPRdInUGeelwfiAk7MUXpqP9bTJBJegY5hbq21B4eWIBcutmY+i55cPrqdKoB6
O4r6OHrqTxTIkshzZW1TWK7DEWDbPynB/1FNjEP+IcjanfBd8KbY30fu1XKWdJ7P
vomoLbdjDhzq33KB9j+qN5Dz0I+3DJ43ncYOykreKsWm3TxkQSUEWXHMTxiBcjjq
sOHFeZMB8y0eh1tW9wgLSADyZTbqGDYlH5Zr92xiR2FIWkS7yxbf3XjaopnAD/vP
cni+3SnsoXNvqVUzjF8ss5jsKCXShFF3nfO/A5HN20+uev2G44btJJsYayH2aj0d
FvhbjURrT80kn3JJQxuniEiVdzHsnhfMAuf4CloKToVtwd4Rjc47DToOEOBe/nsg
2EMvDZ/c+8ddeXpVlp+Sf9ab9SnJlQ8we9Iszk9AmyxlMaEYeZxUuapAReAZM0fH
5xIXocnE5cnKm+jQJyQVX7nRxucLfdC1vKeg7Np/VeRFw0YSfw43Y51j3TcFx/ai
ZQg3aUbajZnJNz20AxC+waK+69FkILUcGOTGpvlM2tRckJFtr7YWkcAfNmB0ww0P
/LxgB/OHbRUdk8qVGtuv6c1HrS/Xgetm3YnN2f8TPSho9IhsOfxn+MBqm2FR5ONs
WgFKC9UTqW5vB8SLe725FTfWoKr2dpO3O/YiEniva+OP+gl640dmURjOni11aA9s
FE1cWglD8ui6RjeWvlxWvXFRQsYOGTlm6JI4EmHzlJb2EilyGlqXV7GCzrajgLBy
1YAH+x+Jpa4VSiX52Lv818Fxt9AYKko3flcZgre5LQBBlVWWX1mCF3TWjIyXRCUu
abxCkz96yt50xk2rQy73bKq/OR5f+874+bPtldUE/K9WWBQZdQJZ3cc5qNPxx5zQ
u7VwEyy5RnqX68K7d68M4804/VSGLl2hFYswKxg0fc6XK+Wui8Tn0fZC2pSCoVLe
FfQrpfkInhpCFfzPeUVOsSaXu6P6o3+uFBGh56GSL6SUyJpp3y4XsFvyT2skrhXB
OSqbxQ5fXWQH3yKkUIzF1zyajKfBSX6wLoPd9EY1cHBQMs0ugUjgeJ9hXWzMSQ3n
hWMVdcrQobdyIIhU65p5QokqgdqLdIyawyWsPou/lpBjQ4XZAX7uje2AU4EQUZ4G
F4cFdaWW1DjzII/mMLzFebhF+S5pgHu/hx48xdZIShpHVdeFr3R68NrWLFy/Tmi6
UZslE2KT1fbVVhd7w/yr8Edf12Fwo+ov6MiyoH05mByCVcmRRujCvTPthKP2U9T8
gSoBtobIvcMm3z8iMefhODJ5EUc8RBqQcc0SKYEb63iDH3e33cS8Xmatk5yugbYa
PgBF4uYAYOtLVG+tQfhJC/1Kz6Y8uKihgp7vWQBnDfkvYqIY8NvVkefAKn0lqasG
uuVKb2q/QBHEb+5hS5+EV4D79F37uHHoiKOC6fPBtztjLIrcOrR+DCGRjZFXXP7L
sQqAwL0V8bmw4DHipn3hxZNms8AZ0PTxPWmwVzUdrrUErZxOkCygAOCieSc2r+GN
NCxl8Rm8sXiN2bHIWpM/8zQPwlFixAJO4VBi48KSBBddG7GXuHkOKjJjPBSPZkFG
Gkr/3NJD9oHO6ISkWVS22CnX36oJEd8Jk0s3400IBbOHJesfnuMGzSghcl4aLaim
esCKEHN8znCNGsNRZyLzdZZe2pevWyKyxX/DbTw0eant1X+ZvBnv1MxM3dcSSHla
D9i59DhtEzQ5/0I+YTpBTbYM+Vaza7ON804ufn3qFJyBNxdRv1eH4Vp9YtuvdL+R
DRYRUXCzO78a64ybYfxzehCC2NQtmQfsFVLUcTzDEwFOC8gTSw3mPbKMtFDEk47r
iIA4suazNPKwDTK5RPqlbBYO1YnHXrqrohsJxCeZl/Z/Y8obVMxxFt8KUqWQ6NyF
4XWOYPLFdMZGDXvlqRKAGVSmfZaNFM+SseKsUz62C5p/QYu9oVSdvji+bE6YlLMN
oZ3iQzHP4rJWhXrzbA44qjbJtocx1cBY2kWPH5N6ClBUrSaCncWZe/C4/y/doGQK
8b3yAEnWpG5bPQP/XUAhjxazIJDyh+PFlxctjcDpp8JUUn334HmGO8z8YdiS9cHI
AVBZ6a44lmcPfB11MBWAHr2Ix2QcSonI3sB0OQea0nOcYCL8TnU4yyoEpRvrdDLC
nx9g5clxpfNjw2R4n+eOiwfpy5sF9QsM44a47d9XyPq26knCclv90NKL2j+krM+I
Y0hLauMzB3Yime6dnlvx2b7keZ66Bvs2eTRR/TDJSUoZqbLIP/QwlE1Hau8srStz
u6V3w7Aw4nREJ+1uI301JYhHAXC/9LBfPw60jCD6186fQS8p3Xkt9uJ55ridxFn2
Bt2RerlPYTzqQpsfSZI2zsusO7VBgt183lR7fLgJRCToU1H8vXGguYihYc4Y495c
byY3UFgBDpJZSCZHXmvi+B0OoRP+1VYAX52ph4wHItvT1m5UJu7dMcHxWEopf92R
U+CEkaUXlIz9qFDbzNXghH0X1RX86/AlJPbQ9s837ryGdjbPZkiu+4b0KbE6P7Zc
zoeKTNvlv4GIv6ziYYgQi2YfNeeJU5iRc5ct0V/rAeBIrrD5QTpZAGy0dzepy0gO
RDXsjs1alPfqiXD49bfR9UQaeaeRChwl4aoRJAsxLzPLZF3VO2T+k2ef4qpmn1cZ
BCcQ4b2Y55y15DMDxD6q15V6ErjEt3gqUF2X46XGlX+mFm0Iv8qhgAwQAts62Dc8
Iol09gXtWi0m/3Xmyw08Kql8IJyBJ2yvsH5momlHqvBGCSibX9JJs/8o2eCzWkiy
IPntD2chLgwHWrtsIdPOnRdKNo7Kvh8Jh+cxIfyQ5KU3ag8G7HsovhFzFhXZa0+0
0+9z8ZZauH60a1E7y87x3UxSJZGWZABpRJk0uDiH/4ctuq92XBvWJUwcuksiMRmb
bT6DOv6lpO3w4ifoOQ7lNELJLgORQQMN+fQqxZQQ2vBqk237QvDJjwesWPpmxBcY
ND6/HXXVZ3XIgwwvKyPyqtJVNcSwt2VUW1hBH1xP9roKnyx311DkBuaskJ1079JB
w4Mh+qM5mlYrJOt1Qddf2cW8B1sWyeusguvn1W6BkQoqW9eqqmhbHtTXnMA0IZCg
nTKH4J0ZdYEdlB0zjwx1UraEXKOssReEK0lVTsXYtwehGDcMq6rf5B6/wSSt8sIL
25ToA2OQF67YdgAqbMVD0kcK67LwkqYGPScNRGvyZDOLssRyXz+VjIKKGnZ3StYn
110XeVKsDLybghdA6FRaqrYHeDEIfvy5PXZOfMQpU8Lo4x5K/nb8cEKAhxDFLXri
LkOqjkfSQ0Xl51Igh75dKpPFtYDTml7+E0vvX191BnfdUKdGR0NVIlXGWLj+Iqcb
bSfzVeiQIGFLpTgcMTf5VtUQLAuYnyHFIN9tslN1BqqUR257jb7Wnq1sdX18ihlb
qWP9ex1clF8kQtJvBroWdnKL0pm1PEAPovxZlzvZ9/fjor8AcfU1jn1vXFL1QRl/
dvnHrbKPFn5CCxJxxzXQi65gCXIjSnAvgYbT9i5AYEbP+cvxO1zUQ/kj1QeP+YRC
n4ydNmbem4+ViBbB77PRQq5QIp2lz/77gsZ+zdkEuiJnW6ZH8lMxqv6koIpQW/U9
6pBCthpS3qNH3V4stx1rlSCf/j77Nxi+lvWHV644lAY1cmoQJk1MTYUAkQT/6LU0
g/J3dsuVbSG8J+/QZ9uw5Bu83VMUO91JJ0URvPHJ5yA9p9JAVKHpOsj35veKyr17
oIEAnh8x7TvOvywMfsNjP5asbPXBF2oZxn99s9wmbariWosDrznp5AD98Am1pkqb
GC6T3buHNEp7Hjp0FDkrMtSC7spSM8Bubg/QRP2GizQSnyIm60npJ4xMTd10jKHB
dhpcVT7SIyTBlWbRz/R710M7eIhQB4ls1I6yZYxzaydcwNTZEHRUOW0Uq80mJWgg
agf1I8hIYsgOWyUVxPB4229LZxzencNEuftBFYo74IGQzHqkhIKot0vPa1rXF0BA
IsEwq3ttL+d6/eAkY/CYrNEGtJAFjzre1whqxhkXjdnQqoFS57VdELj0XYrK/2KE
j1qEnFUBsobIfKujUxI/8tdiVteolvA/HKAWYre5EYIJ03/UuhuBAHCprYCkmD66
DmDalLWm0ZQ5hUp286mgS8lTT9Nx7hNeU0mZlhVSFvFRlQ7Z5y6ccDl4pScoSnlU
CEWdWIBJ0Kzb2UyA8TmcPqAhE9+/98/5F5D/64ZMc5BuQBuWgB1b2G540v7PWe/T
eeMv6eDV7ll6e6ETxy8lN2NU5eYnZiaVJPWr1PpvFXj0zfK0dV1THSqQpmInp4Nk
MxAYtdZUS6dkJh3z02Kf4Hslmb8B3VXO5SGM1nNIsFafTREdH4TkoYvOLJo2hEoS
CtS5G/g11lDEnHNHWnMCebrC0IjhrS+/MnFFuhIcbvTF9rYwXI7ecugSuTwOiveo
8OnY38Kfr9y0Vrig6FSnGUQOf8MeGBcSEc75MosqQwywYJkYqwZi3ah5yOD3Oo0G
yBguAwe/7Cb5KJAldcvy1n9M36v/sAX8ostCOXPEuFi0smsG7A/TSvabIJDaVq2h
HC5gGftRh3vH/6+tgeHc/0HmsgqwatdgCWsPUF057zJBlnunTq6gkYHv3BXFeDWX
3I2wGwDTV3aHzDF6f3YcNYvge9YCKUD+sypxwfEQiMSs3vE2Gjm5EKsDOlw/jFij
Lcs8dw9kp1Ej1vOjCoup2E/2daN3uLc78VkwGO/+fFQgg/XAa8AsWNYEtDygdGM6
9BY/0jb5ov0WpPseoJm/GO6Bp/weDsOAzJw+RkuxrvGw99E8OFZocAdH6HijphGb
aepPP0r8p86diN9z/8/QJzbE90y4Zo2T5GytSovEfOvto0Uuu7b7lxeJyhtkoEQP
+6fBhTSqeeS2kdp1Uf/CAbiu4Ky34gDrOMvaasiMy/S1RB1MF+PgGgIdRrHl9EtT
89+9sEwG2s5thscjR0zIJOu4FYThHi6WqsBNvY+43+J65pFqxt1dvwyhwTafPW25
gM2DYUa8aldvMkZB/DOSEEdkMzfddurtcwJhLXH2LsnNQ+i91vTqWN2Mk58hA4mS
D5TMHAQHoMm0AgNI3dkJuh6/cwST6sUKfgbmDUVDY2xVEwxOQrcBxHoh+nePCyRj
ekAtvvNU0WgsbT/65vbEJQ/MYkaSoKluuZuWyGOIHJ/gKrjwGo0M3TI3CCp+e3NM
YcmhUT5BlifxcEVGmzKbLWh/WkDmWp4XdRVAW35zziK4GopaQj5lLROYWDefh84f
k1HRDE4se5QJC24jVJqIWFRkd1CSXE7kcoWUbiNBJLyW69YhvTfO/LzHX6eZ44yw
0Q4zrFlo8sP89JHdzHFIJ09d8MxSzZn3h/li4yg7+4XmBf34O9P9Uc3KPFyGTtQV
JZKnKeF8RO2Q11q3IAepmm78b7o36Yp+sFGVHirELjxeNr/39pp/AdF+S87/z01r
FttjKLWmVj0BlWWmGn7Rw3HHUdkLKl/XdlZGBeY3PBrE6N8/CDOj/XwKR5yMTlBW
SWCpvS9jjLiG26LOmIs6k3JIuzsInO6GpGaebIVWVCA=
`protect END_PROTECTED
