`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AofHPHTFX9m8ScCOIHjaDCAiWJnnkFcH7MDWSPVoaUDufsiGJkBzZqF9RoM/Wvqs
Jaf07zfp3/B+f8jpLbk2lUXaU34aSCAWfLw7R/rQ+zKTNkBWsIVMjDl4vCcvgMcO
jxYexpLdZkysj6hpiwyn4EqI0eCkbaKrf3E7KZ/tyPbVZLBOFUSR3pMagLeVSlcX
bHQolP7eokmYd/lTliiJrR3tk3SwVeQ1XXRdns3jewKhQflw36OquO52l+Y1BWuG
O072lr+VasRxJ22Vfk41cBJDS1LmAjAa/ENOC3Elt1zn5Zs9MH8CNdo0odblBfty
mEhLD/vMOSGgCEOS12b6G74f8h1Z9+Skvk2UNXdxGOw8WY0o8+7ENtIIQLSdZ/1n
/ER5VwBg2LoT+wd1AbRhlD0Do5WTKlxBkjCfVfpFBpDDDm6lhOtQ6gULYnQp3EfD
pmxI+FAGCwyaiuABzNmhR2iP6G2/6OE9eVVYlwEKvamGA0ahjkNNIsT6IyxE6yQa
rI/oGFZg/TZPsXfe4VLETK+V/9YhSA6nf6LXVenMhSWujmpPFFCFGq4343nlTYG1
uqji4OmxAzJOyh0bNe0viQChoyQkpVwg9LtOTxpl4gXUNl285i7Kpg0e47zP7B69
`protect END_PROTECTED
