`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u6BQJvmIu02f3Yysf3EADF6qaUU1swXF2kjEABL8D2YnWReechUNxr7Wr3ROYmFH
UTU3KHZS+hcagbVooPYwjFSyHTamYuNjxv+M9mnGKLah0kSpIzsZll0Wx9lcKSdD
pLTBxKhge8NFAifN6c8zyGZAUEqWw3rVkfzvk7lkEk3Ir+YZChzefZkrc0DEuOiU
T/AaBetLkr+S7v1seFY4aqu0RiwPw65kNPq6u3u4EXZPPl4/cn/P22GQHUPcyamo
Wcm8m7uxzAlF6zD6eKJvX9+wZjOOhPiW9Eh5f/bnlh6WMIyWnphEeE6LFo+X5+g6
dbmBiUNaDr096Xib2L3f8iZLc/brOSqCW+BuloQ44yPZ+Pqh+tE/UXlwwyBUHozQ
`protect END_PROTECTED
