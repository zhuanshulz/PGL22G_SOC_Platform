`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bfhZYin17EQ8sL5GjWkrQ3I2ahL6Iiwn90h8Yh6rXaKg2fScxWAJvfqjRj9zxFir
RB5QDUPv0KmSIYUmUw+LlnvDl8wNnh3EX9s6Xq0sdei25Br/OpihIOkHBiHpW3GX
A1Hfh4fRJcSDxZnohqemv5OKJpX2oVbRNc9i5XTG41T/t+rYh9cShXFCM5Iyvv+C
3zx8UCUYRJLzmXLJStHyYB5tRBMDKzdMft0wINp2WFQeRKi++XYtsbYNYwuFroMt
/gGgu6dUwVP1YVt7KWKAVHWx2v/p+b6YN1JbEaxJ9oPrLKBmyqxgXEgBtCMNhzSZ
6qAXQUpULnYQlCBhnKWjuJ2RvqF1IHzmSCPgbZD9fBVyLRu4hUwP/V9qr7cDVm+n
8Ypx+3XhcwBHx2c+TYqwZkPT0VF8b9ikaPNf+bZELhYaJOPOiEZzCM6XTONM4iUe
y9cr8W+cG4FOYPHNSlVhL13LD6ctGp+sP/vxwdtCnwG5eSktKeOG9npIW5T9N3Dt
S34/oGobgU0ELefkUCfWanbnKF4xd8pEXwCxdWToDqSeMQyHyCLyp2DwRHCx5YJV
1kP8p++bQ2uMx4wq3xQ+/FVWcO0yejYRjsapkqY7t0q/9k1fid8qsJ9qHmokUv/S
WyIaIThknJd3axKRzsVTzA==
`protect END_PROTECTED
