`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NaNDZ0B117VFTgGs7b32eVOdj/brwG0e69uxPujWoRGM8HH69ORkGYOpGLwqmjH5
p4e1lmGCHis+qjOzxQLrUQcfqA3sxtNIhOjxQEf89lTR4qkRcFneTo3ICBt68152
Zo0kuTMMwDOiqiG/2byMSebREMva05hd96C3qbDXxLuqA8+OPUrh55OnfvO9D11A
zW0+W/Zu2pxdJkAFf5nYK4CeAnoVoloYd8z6B39TJjBGfz+Zdp7l3YFP67mIMsBS
xMwk0djUy9ojK51ZhXDM4EyR+WCBgGeI9gwA4jk+TaiQZ3gfalHlJ/3McIAT93Rw
soW694G869NRPVF2M8QZAUDKTRYOEJ81rQQ/Z9hz0l3MxmqO211njLzOr5OGhJc9
E1hbFFPbmQFWh9n3ZOFi94yEK5KYT4cG27uSIx4eQ5riZgb8TPtGTdiRgW12rrdX
osXgrR/HS/pWVdO21zYYKzpiIiobQ+y0q63L98xUQyEiomJ3bMwoPSY3HlSUG599
P/4qX6mh/++gTFj8bqSDYA==
`protect END_PROTECTED
