`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PytWVxsnS7J10QegLtCof3zhLBII0KB7AFieV9EfXzgro5SD0m7EbGpeNRc72CJ8
GQaCuBBP3MApWL2mW+eaOjBdTRdSrS9rJJlGqN9bqgjxcO71VU7k1r3vg3rG8ujO
15Gnh9gd8oPA84bvLJtwFYMTs+2zLFC2vStYFkmVtZaeLyrQiZghOLYEGgPPy5Ke
+Vd6F+RM82GjCDGD1GH8tAAK4qZuJyJOtnV4Dkmrm6YNFbHO7d7F2OFltjooRU+L
fF4naArJxSqacvcFmVpDgxs39CXCgVg/bbH3CykPV0D+tmrUBXS6bFI3llJsd1+v
Iyl++N9SAscWNzqcBOcXqhSG4YgEQTpHYXpT0vNB1PMt1iv3VlLnpa2C3KJSMMmD
POHpzkH1q/KwEy3mrDOXhFQCmPpN7IVV2mMXQOUWY8wAQhRvLxNQED8794aUJ1CU
DFB1aAwbWxYEXcNuL4TGqsTOE9dZ9kELxzDcovv7RiRxg56q/Z4at0EZa7sX1xAN
JVEPJvmx1TLmVWtev9zfx+5RodXgNgvhGkcuGZ50RFyN6sb+0HSqPZyBdnVxT9zY
nzcfYV5Tn4H2rsO0bJoabM/R9g0oIK2M7fM1l5IwAvQtJhBMCUmrSEX+XAN0081t
1Kw48vcPlPPkJRw/t89kapKV+HMM915yZsm086zreai6XCO/hPbgZqode3LkZW8y
j1eFcy5RG2NrskoGNK1TVAQcDB4H3B8TWwPqWVnyc7MWlhL4bB0i3YCQYQjVqEb4
n+YpsCS5bk2cK4d7LhAvSQ==
`protect END_PROTECTED
