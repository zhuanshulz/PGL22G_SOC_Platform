`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CCkYVPV8Rg5EvlNyzqMFErCvLdbR53B/4my0JM2QqdUiuqY+zQ0mq2MkBXpY64pt
Ma80LGp5IDyCVBmByPOh3R3lIquOBjS+mFqifIK3QXYVXWeVhiAC0KLS6wZHp1T/
mipGC2+sq6UUH2nAAYj/U9Q0c77y9X7cf4x9eLMl8ePc+ewR9QiS28NfSc27+pNg
slH+TlXGF5Lul7jv66vJT4anz9KqsKakVoBGcvBxKOER5aib8dB4du51LcgSO+zZ
uqbCEd8iAoOSICiW4nC9G+V4VtXRyVY6meLJ0itfdUfYzNAReAMT/fSwhmcvWq3o
SA7y3H0R20V2oqfiux3OD0QiDliSmO0+1merb/IhViA8jyEn+eUUCqjJLm1L6uo9
1IG+ky9uNA/HtzNiPSafP1BIC5OkJ/ZeCBxaF29zmQ5cjV5QDUGjT5Un5g2/6ynK
PSRaW7mh+QHIyhYB5txpH+kV7rPWswpHymPMW80fKYLMFLFl7vnA++WxoQBmEzdY
dM319bm1Ihq/83DzXJ9Lt1Et0pZBu06uE7dIeUVtNeyRZ3ELTc8/lKvdiYQB7Kqv
kH8fcZhsuaEjw/0vveVAkADusbrjhzExiq+Nhij54EMt9oGVH2VGPrFX04PmhsM8
ffHbhYldWvswmiSQ3Nx6+3sX/5jLLqlTwsg8DC44UA9pEJf3ftl2hNCpdUdwSpgJ
fbd7pmJBYowc1bV2z7JOjMBCTNyXRuNiNXTwThB4Kl3ZsjYkUmDdVPQIPUIGawPy
9s/JH/Q9eXl6YaDMPeJjlqxWYmGkgTniSFJSriZqv7bCsUXH417kaITV09/NN8fU
NC3xspbI44s0jud6Lxa6PWgB7wR/wZn2Ysg2XQWL3X28aYbzxOYnrT0+gBFis1lq
jaCrSPJuUdknF+3J+GgLoGmUP3k/5BdjneAtUJepnDAfDOOP7h675eimY0H5NdeF
zN6hf793DhSGyh7N36ONxm41NxKqBIg0SOEWQvYD1nMz8itE6CfUnFGVoh9OZ+x8
JRwt88HBkrHRwk2hmegDgHJdqk3aJ2DhWvMRWxQzuWWekwXFLQatXDDLs8sWjXgo
NIgZTrJlrY5SRGOMudlQl1KbeHaV/hfuRBPiQOb1eEDScZCnilUgR9abmxGQew4D
Bk9kz4Yyz1Ex4idCy0fd5GbOplA/RyMwmYsAi2qqTBSHhjACHnXVUrXQgFkZtgNl
+fI2RtYHuNzL6cpmH3GHe6XFl5fG6EHlOiPXirlotZMIqCiyW85+vfrsEdUwFNFW
1JQwwRc1NR6QJorHRFP78qA43OhPG6eQuvzkHYqIZu0vt2bgSF8ni0pGqRW2uJUq
revuPZUHr9J9MIF7I8bAggKKFxP/j+ByHRoExWi0yUpsgPOjr0OGlWus10HG/GGn
VpoG1IFG5xosDE1Z/N3o0v9l/Q0+Ji6VxNdb8DMCUSD6BaQpaK+5WMo8dNYXa+r7
EDxBEWcPziRrfHk2M7290Ry1UlK77taZc2QCNz+RqCAtGcPTu9uEWtmCBcTzK5oo
XX0W/rWN+5GT2TzTw/F4VtQvznLM3gCQeygV8ojQe2nQSaqq0+HXjClu1W10OHzR
gfTJZwy0pqrCLdBGUlPUB8HafmwNIaCRrI975Uw69PhqNAWokpf+hmJ71BhxNNaw
FqoDarhQ5Vr98uUfcaWpoS1nz7+1GADqt8g6J3FtcS08hZ9EK7KU5qEX9iV5JG6h
Mf4Rcqu1I0pDHpvoEEaiKW7ShtqaKc4cbXIXfbrChoYRbH87+WL8dYM75AOMw7pT
xA9lXhWpPcrRM8O0GbfckIjmlFutHDKLW7uiifJs8M9TL8qXRnOPeAxXHFZcvLC5
9p6b09YD9shPhgauY0rvGz54ea4JAwT7rwbUrX4knbTtdXIHle8pkcz1LnOdd4i1
ltdc+4qkVeRITg1O6XBfFF8Gg5kM/f5qyKLpGMG2e3cx3TEXSZ/9xepTNEhAhGR6
BynFhWFE4HsPsZ+eIOSqBAuwR3TYKRJDTt/2lU1+PBYOT+cdUdEk5ybua6mo5xis
r21Qvb2jRniyTAiDtvGD1g1c9MOCumKjFQmgiXOYy6vBoPP9/indxpdePM+7RbcV
R/z72wKykh7K0X/5JflZ1HngcQQ+UJG2fSGAHH3UIlfT1Vl//7Y5xga9gmTSnwAd
AM1Ooz/fb5RzZOt43/iYF2XBHrhcKPdRMFoIPpy6o/jB3E77yJZR9hBPQ6ExpyS1
G8MFNJC0qbw3uzlHC9mvmJxkqOWx2u1OwpGqKiYnUJHlaHcy6k3euuFnTqG1CO0R
Uypy9fkzYCbny2ufliqxOS+6wSsxi0zHO0SeY74odrl+i0oN/V9FISt1MC5GWVS9
5ag5/gvuIolvBDwExmRmQap6rzRusBwl8qQnWuWLOzsDfA/phi2P61HmEUnAUKP7
PZKKceKYW8FqKe+njLRjxv6Td0tYo0paUiL5T+Uhc/NkpRGRnQU6gXrFQaeM+b4c
0P/sJpOt1jYVun9yL2TZaez9iPjIy41xalnlTMIr85B/TqXYJMC/aoH+JNOgFwWf
E0BTDmC/IZz/Ay0glFI70rGOGZnu3VGq8mtLgrIw1rE5lnueQEK9h8l5JDiRK3GZ
wmoUf6VHJR+Sq1n83HwU8iyE2wvDokCM2bRude4RANnUiTwqllIb2HRsDUwt4fLd
dGNhKLp9FvX+CAC2DbwaWGJ6PaQ1g5Rj1pnKch8fd+YY1FEyYEXXNklgwQACWM1c
xVkF1OBQnNhXM5ziUdsMSB5AwHDsDFFP3C2+LICevGBo2XXXyncqMucH5ZS04/2r
XjFWa4Z5qUfD8UAhbizjswSpCY96L9H00PhS3T7mAJlEFP/gTajqTqMxlhvFBP9b
XxYuXGEA/FepzZIWmJhmJqxUqu9miDS+DbTvC5IsVfX/30x0BNNbuFeR1b8jDAKi
mcLjUKz2rzQhVdfI4HTM8lTYEW/KwSd35dMlqrDO2h6hW4SbZ+n1mvYNZoCAq2Ou
YYZlzhDJ+f4HcOoh+bZUU+Gli1bT25jN8I51PTcxvaIznW4mL0HRJSsxipTY36ab
7pFGjlxNiYnqFSx/Y+HgyNLlwsAgjx40e4MDESe/SxOmcBC0fExj3yApNP2+ZPxI
E2xxY5S8Iqo37mdGRDEhh/TKp3C/UsSAGsjr+pDv8Qd1BoEBm9A42TmKnQlxcmXL
H+ZkQOgY1e3YvSOBUYqbN3Plzg0MJ0a+UsWoFHu5WsMbwbJfE1fCCVFwZr8Cs9m4
ZmuvEomwxBOqz4tWxevn6dDF/5PiR39GVJ3VaSTkB9ipCbd1CZs46sHx6CrBp6hN
3XzJlda9vL/eLeLzHTt+z3bmQZZDf4bAGMHVGuAid/u1AmKwFX/1c25S62ghoP7W
u0sOFEYEH/VWdjGoEaID2au7HYS8Altz/6iZxwUa7PIkGGtNJPn5g06B37STEOmq
4izPf9EQS8c24t6Dri5DGwOg+p/UrhxS0TAQhlN9wH9ze1zJZ2H87BUk8vye9bok
KUxNkDy5YxdThEXgbcCMAHRgHft88joPCQzBzC6tiKrv7Fbr1iWcmDoHBK1F1YAc
6SrgEzGzeYSysnycUYwYk6M70e1vl1NqhCVzPUna8EVPgyWWJxDL5X3HAGu2Sipx
PzRRzYe4KDosDtQzthmBI2Jm5UYMN8kxbF55WeFyzrx0mf5wNUQQzfDf5PYJqiPl
Az1ncy7zevao2+FT9oGDi9BdoQM6n0lHPq82WrDSak5GrBgWYZONrCa0t8TAC9kY
ygEspdQ+I/EtoieNt2QVIab+5Qqapcl6BgpgrEmFiFdzKU/EbLnN9QxXXf0QcpSH
hfeu6hafC/pANyg27LqvxPcKBWPQl4rxalXgy4jAHVTSMfS/oJ6fVPx8Zm/2DSag
JzmFEsJ+HLBZUD4W9Zom6P/WccLbCO04QmllstjE/84jFrTTVUsdCpzVKsipUiDF
HOWzkpAAGtVLHH0Gf4vDVMaCybP0taFwqqOfxsRfOec=
`protect END_PROTECTED
