`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aDR6lteVeIQa11F/q5KhRZ8ffgVw4WPm0oISZ0Uy45E6oPRyhqUJWWM/b27WMJIP
T7wPfnNkrdzCWgk314yES7A/Zo7tYPmejvWKf2T2v/RoO38ozhhNiP9hwrPoL1u1
FfABTp919q9bZrxkq0KqAbuzbDN/6/QpuyvKT+1HHFpAxL8uYzJo81o9led7Q051
zFgCAsvDydL+IGDsX6DuDnnBo294F2kECpgxy0ih3elRwytfBiVnA3gPH1SMWZCZ
XwgSma4mmxvi6CPjf78PZusbRmgLTCF3JWyGMDCJQnzaii69KkbT/MRBAnE7rbcf
cP+/FjMJwfxCQZWpXpYzMx5s/5CTAGkdg0AQovO4Hp6H8LqcwDIHWkBJ0r/kHK5V
mDhMzg4tQxOHT7ngPAWACLwC5aMb0lpf5aOZ9YoGSKAr3gexOGp669R4ucUaWUzb
94TRbK6vyyPXS/Mfn0tbhfusvf4KNqXmm+obiEQ/iLhYB7mZFxNcAArdDrke7lhR
43fjJ5+sOFOLiBZF9NwMW9gazwTYze+0GZwzdwbT+7Ki+IX8p3iXMugw3EnGTA2H
TaincBLYwalMDbQ1DIst2Q==
`protect END_PROTECTED
