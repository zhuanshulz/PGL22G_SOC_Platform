`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uz+UOUUy7TeslxPtQ3unq5QMm6PeQoKMbdyLPfJIP74XfymT09ztOQMqcebwcjaR
UOknU9FBWVB5GmasmjsNNpEHguXQOqVdl4dgVFV3TXrnY6YYmPw4EFeNA/2U0du+
vpqx1/y8RPD9ewk89J7MZmDZaHDvQUJQ0Ff50IBDYqjsRzGYvLiPX306QQhHG6WJ
LnuayFajkXsPan5XWcRmDEQbZKHREsnUrWb8ePYmCrMGqlzb9T6grgUJHIkcssM+
/ko3a1tGDXWt1XXGvihh9S6lqj1pjg7rDyJGXFXM8xEPM132ZBbCBjeuCpCRnZkO
cWA/NK937pkjT/FxTA9rQYsKT/vtbTOUpPAP15D+6OtWvO0bAhCfT4tnZM4beoGD
HpgyMB+sYU+eBudvxEqa+ALAP/zjULl8GaOh1Gxvc95CD50MkClBcqTazxes8ffT
lTOyagAO9X+x4KA8l25vQNvT53SejAU8NwoWjbJobPdxnaVQu5NIjEQR4hxa+AdW
+t+kV4c/MRyHVMmsyDgS9m9DHHbgsgChUPCk8bYPgNABLeVUpHbBqAqtqujUscsC
jXwk5hFBAiUCD7taOm4OwjkhlU4n49sstezCAXuVXPkonowbkVOlSvZB/iDPmDt1
4ChF+J+3nyJ5QuLZYlPG862TqSllh7tUzyEffa1JCoFFyiTJWTbP7xBK+XSqEKfX
Uhopxsk5W3EmNPF6+wMvTpMxc6eXwVBAP+nf7cwhGxtHglmJm5h7qxBYWy/dwzS5
hG9HRTBvDEMPK2I4wnVY8Y1/7pmA++fbPJJvAJpusiCOnvGMlcubdLZYaK4litTW
iqg49epmcDFRPfuuUXvFd3TrMdB12UVsqTQVvYol7mwarCVT0YuqWep5H6EZn+Uf
6O+v7EpxEi0mDzrg+16qjy3aMpSEPARyYJEICDN6uNPZeugIYAvgbAnzVZim6TuE
DPs7rPPV2hE9oYj04+IIHx7BEPQcd/3gXmHgfTexe1Ew2GRr7tbj0PtvH+B6mOap
OP6he4Gdw0bCXwCBbHMlZQ==
`protect END_PROTECTED
