`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b4+GyJsuWkaMobpgsydoS1/0QvCkmftsaCCSvissrcLGukTbE7Q+jQkxmSY/pPEp
ZT0/mWS7V5K7ikoMouCSYVhQI922Jgf3izxCbn2BSBS1uQ1q4RcndptK5CGy/eFB
zxRT4bQZRZnk2ft/G7TONmQtvnZ4n+bO0fD2QzSEqH8uLqpmpCW9n6AfEslhGvxr
9/6cNJYsHio3dM72uRoxmPSz1JKGrqAdF468pyM+xW5fsgjaE1SF9XWSMLa61Vfc
f27EaaRU+0QLesyaFXnEXnqSMs9CPda9OqXNBBxsEtUhGwaxhoExOH+O15JFXteW
vNRaOGGCKnUlLsIz/+7ayx5RfxuhuoVn+BWGzqrnFBTMyEoZouFM0+KefB8Wj+ss
sXsdiwXgph9FxXldYDCrDtPRJYQFzZvRpsQM4IbtSeGFNmR00jPP73ozpWmF/wTb
ld22Xgmy+ksb2o1sdvH+HfcuxpL8P4re/KzybiXtKS7um/l0fyx/7CkQjjDbeRrO
ETUeadNDx7REEyGaaSnzpa5fUAgFAO5rPyj2UKeuL+bNyobXKeEtUSYDAR5OMQba
y9F1LBvwhAG48ABbVyZ1eCJsjq2SpCa6AX7PkHqRbQnWA2b7KcVTgfRQDS0vtAdj
aieSrpfnpK4wTNpopWTfNOlm6S9ypV9cZuLyPoWJ3xasFLHgr53C/XZjMogQHGxy
U1NSXk5gzMgA77iRwv3FQoF2ZIw+5JUBrgx3naqXnYwIMMeJ6Zwofp2EnMDgTx61
2RIKah8C1hXLildejAUbxvGGg9kxwgmg5wl9jIlqj+gSOuXyw9buPIJx0zw/iky2
7EnBaOIdoIUMHSsGe+wmeHWa9TfUitmtDVotHEo6wr/WpNAdcA2+gCkIHF6DBQOU
`protect END_PROTECTED
