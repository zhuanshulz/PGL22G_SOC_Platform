`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nfCunphoBlr//bxsZMe39F0X6+0E7WD08yN3xgwdESWjI+eErXpBJ8HVWiDjPZHn
2lTF5KyG58j9UFDL5QK1SDzG3Q9Yyo/9mCpu7HbMLkqAi3K2DTpb99llo4R+37Nx
q3EFEWL06mo8KRNJHmOWoBHd/kUYR1b5GGSJJBC9rTId2Wx3TwuYzJ2AwzPDrRZH
82GkwA+WBMPW/2sF05R3gLNtKFX/cxBOTaYaiGhWFdJXX4HdNZM1xfhagKp/FEoq
jYoOxPV+5VNLkbFa5ixS/WT3MI0mgRfkIm18ShH+a80Ze13S5uNQKTuMqavNjMJl
/zGqnmQdbCxn3XryKQZiYmsX4zJjh8ib+mY2bz3FTmq3pJa6TAZVVjnbapcRDOWI
zlwkZTGHc1uacFY3cBCGse5nVc/hfuMOsxja5TXeN2BSHXs/+dPt+PzssQIleVx+
e8hfVmcK0mc71Bj0wxYyuFCBLSEJxehXTAT/9pZE7C1zwVTqGqPI3A7nhsrR/K+/
lWdBzuWXpmixfo0DHjA+A8cFH624tp9leiOF8U9PA471GZ0lM8Q559vq0c/Nidhw
zSCXRG96Pt92aNQ2rAKjpWPnu13vpcCGqAV5enU0GXs2SL7r4n9GvFRxawxK6eGB
2pt5tFy/QMFU0TEIPUWED64EDvxr9bNZJTnknQ7V22wJTd2fbKG9A+OQsm6NydVf
DrU1OToISmw/5Lsx5JRjtfs8VwjaYPQkgGXRXaDkgtuZ0VUzlC7OFB6NH81oMfnZ
apGtCdp6rs1Zkyaf0BAnud/9oi9Ld/IqliDRu3ouuir+zEJ1cXSUI0ocB0+Qlsah
NGHAT+HCwbDtDpMRRfbkgbCFcegfRgFGv00bHivhnVxaZmvnrqgUHH62d2pprEOA
bX7mkU63Uc1FouNE4/V0+DqWI2JTcpwZvfh4cLkj06aynbQhfedmhrFWtRXPgus2
ctFC4U3X+bBruMFfF28BF0lf6Wwy6iN3aBYKBC+7CLAB1xfDpVifbA0rjawl8tNQ
0XDNUzRxrS2AVJBrQ+sUbJLUolyEmU9XBN5kI+g14Ad00JsnAOS+M9qLZRUW1JeT
KSADEE1uz0aIOuzowwTKT5UbqTDdzxUN3bsdJx6lAt+ulTMIRA7FJ0SHVvwpO3Jp
zBFylFbUieAXw0VKuAptk+lRyFESm3L48PPSyDoN8Bo2Xh8yTpC6kJSPVHxpMzOq
Y8j4YPcLSLV0jglXadvKkeXWSDXKx65o3R49GDfK4CUyEaPrwB7OzgL8Syt1ankv
47P3zPn3KQwWBOeX+9oTCzWRcDB6RTMORhE6e320IVLe+ND6fklnag3119GD+OBI
Jl3OEU0Kx3DuteDc/qrFKlZ+JR1m3c6P6OGPRc6GXs3fiqYwbae7+vNkSvQAHns9
IdphMAVe3aWEsWYmcQj4ShH272QjNm4MPoQsE34Db0spgO5IX6ZRguGJC9/yIbel
tDnRfAGkG43G2sby9G3d4StAglI+LTitRKiCsM/hnmgAYXhmbG9CQ2gJof4VD+KZ
C7Hz1I7viN1iB8B9mMNLArfs/OrlnX/Qx2y8VjE4pO8QUwvaRJeYqXb2f9KsTueX
1u7O9lRoqMdjiRMOcNcXGXd+nSSnCEmz+XfIeZnlzeLBMyTxCc1EIUzvjk8ByGsX
XjyZuNFpM/PKSYBO7OUWr0VFZWkqMVwLvyYzvxaewfEKWPoyyfe7OFkstEDJqeJu
N5++tHEVZfzqUWkWG+FMdQ0eYlYJoDlLiTnpdycYPwkRhCIXzqQRqNNTeWqI44VE
kgExajZcT286JUZk0n2H4GtJZNTZKda+CSFFMgPfes0Q2Yr9nWAc90+tEcFQ0Siz
A7JejfPuGzZ81mRRJw0vR2YvW7W4PPe1mUuPqxLEbI92tjOYbUBJoUA+oe299vqF
nScqbX/KQuL5xkpcNU7IsetdfiBLPV2UG0HhPSipQ1p0S5xQGUbcgYyga3RuKaGA
bVbgPc9hg+/3pXHSSAq6uBFL4PlEm87EzowQsmB6p8YmIh7OpdRpCjgyHJpMN1lv
EvJHhx2HY9qoFNJaAvsk0mmLHSi/Ruj/NtoD4IqToF+fewH4NL255yT7+yqDig7a
9jP20abWlcqyk3hCbx2fn6SaE8GaEApiXcpHwLvTcP/vICNJ9xpkLNf/ENs55oQ6
L916EpF8jOaja99tJ3L6z53MXjez2TcdCJQ0JF+eD9IN8jOoULLVmiCAq1+Qnf+U
fhTX7MblNVSqVUzI4EddhUaZ5mCIz5jmgpC8eQ4415YMiNjyPdJVwAeJaRmRTDyM
Md9XBOtmL8/IsBSuz42+MmAKwirJ/2EePYy5Ig1OIUjnDkLpvPfoWX06iGgyBqr/
wP1LHYGClYRYfAJ32crNfLQ9xbhqEFZfic2Uvp3XO8MHO0XhJwnBKa7i961SK46M
knPq7GebZFtDquGXTOZG3oWpbYuupqpMyU6/IrtADFtRzgJtfJ3ZeZguBkRA+WwT
zTFRT9/qrnrCzsvBBzCLOPgSkgwBa2rm6toe3UX51XpMDs7fy68IPhgpGNf13SsQ
5wa9yGSzLS87uNdjgBLOVDpfmcXx/a6aF1JNmKlEljzeMVVhaI3v5jQyXD87Oa84
ODpjZl4//H13ivAXhPhhDx5dNBHmGtxuydobjWw48qMA0NR1TW9Ly7A90xaGFEZi
lJcrwV9Q8i5JkbpSwNUHI+VAwMliR4QipBs9+I2rwaBo4nhebGZw/+k7AzgFBxko
i0IYimStUrzHulYx2v5J+IeV4YPWZX8BOvwA+/cAcXeSE07jLEfdQpoEmfpbA9AD
V/3/47ZfmgPgZbM4VjOEdwaIaoCFoVKXXw414C3FvNqxOsbP76SyMaRE6/IpfOdZ
B+qm5rXlp8t/YqmeWnJfsEB3mpA2kSDwF+HlX0EgqjjmNF1CFI85FRwf6yJdnzUE
UgL8Fcz+4xSsi0txbBMLgOEaBTz1wZHwPZn8jrLFZQNdAnX+wKTmNMleSPFxh/1t
8sNBbOo20E3i8lgRxl50o6JAnbry7f/XVpkY2MPWecRzWDGubHO2iuvBNoshar0z
wF2g74AI4DVHGrmx0oAVHSvoXhH4vLFAGTmtWQa413U6n8B52Va8VyjQMlU8b6Eb
cas9P7y1MhvVGs0yMyBZcSfmtuRsqeIqScYD63V3XkAu4vTn/szBjZAMDlsQ7nin
YOcYzX5ax3SPJcN6FZ6nrpUU80isFWJH5WacamOkD1BqUXvTZI10SgMLOWeDGxga
s9Dlg2mKKDpHqx2u+p2M/JOOcwPvNZKpgLx0ctpcFX53Bv/eTSOnuwcABhc+TBzX
BY5Oq7e3OCfLbA7tG4fDaUng82lnEat3gEd/SnFHfOmzeAZtqcRpCfV/Wd3Xf+Mh
yh5xFEHIYd5rgOt34m9I3PDK00zftrnLRaGtowhpnRcDirOb9916iwWcj2sY9aMY
hEZo8+2bC2viDBSSWxJTUXSnCUNj81GkBZHSeXlldw3BgHYrJMl6xa1whVKLv3us
lZQ4jbgXFTrp6XImANmx5ZqgQCnrV0yPYPSsgKIjTa7XpGcW//AohvPwWFQU0q+e
fkNpkBahbLgk1lycT/KyiTn6bD5zEGiSVNkAZfG0dlKVOQURjGTIkj+UdP9oW0u4
FTUY4w9OVm/fQpHo21ds9ZuGf8bXuwfcI/QvJyEZuRYFhcpTIseI+N22xPsNS9MC
FtZaBDO7UfymBdqfMl0fPDxy6D/dKNheAu71pyua3fwmA5S4nfxBTJJNaxoU2tpg
0O3XtgyxGGf1PekC1lTtrLnR89nRsI2LauM3Ihzfjs2JWLkonDDBakgnY+JCDCz7
AJQmqRWcA3yNHBkczmL1kA9mAoSuucL+9XNfxafLe+h53PTIu+Lpn0PYMyQePgy9
fgDY3PUULfgtymNnsuwNTVqD513I81DCW/nKA6TkN3Y=
`protect END_PROTECTED
