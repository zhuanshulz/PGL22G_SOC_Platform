`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U71u/1t2tZ59VBbf1OO3c3DW0NvxHyK4IDTpDTkm4dDdOdRPMg0QP01Z5BbfXuxJ
dubQAis1K82vMF0CCnvCSN6aZl1tUVyDyELH4w9oDy8LkcRuB0vl8Ib5Rskxj1VE
PIWGcFpYk5HrK9ifRvxycKr3j+ObOXnDhEh8mfhEy4Qis+uF1/uUI5YgvrmV31qq
3lsojxBt0J166PM62JI595s1p9ju5o12jCaF+UoKTPuawCb2RKrnzzTDflBnQqBb
1UHWKHguWTrHmoYShuhKSRCxCSh5GKUkbw6VyjBmbTiBZiZfsi9Rulc4trXzeZ7O
oS4zYLChFh4LzMEL8EM4smWOnb6oRn5HxwCqShc6RMFgFXFbtWe2CLEIKJQzFFwT
jdOysRHGJxSqW2hwvJ43ivhlHp+k/FOdt7KA6YHT/37AfnqPcpTJ++FhVYF52KQZ
OjcYAjmgxo9BSDg9gRR3XWl4te4hgraBzHCZPUD6JTDwY6AWCMoOSc7g3wCT3A7I
uiB1sbmetUrK63merf93QtDraMmfyMvPeZzeIipmwffcJUMg8W408mKAcQ2vAveW
wi5vZsQOFg2Ijf39SQis6ClTr02PU9+2hkj0EHSdAE87yk+revqxpADlpTMWinwy
Pj27A56aiGW4YQOdCO2OFWBsBo5mf7NZIspp+2pJ+lUJfhkMzqd+EKog6wUvO80g
TC+wViNaYSYeot9U3K06KsWIcIu8N4iWb038sjGX/lX2ImZWXGwl7ZjGo7hg68lP
UIgsLlsLUD4Fn7EqgTtN54Yes5+N89bb9dVTNt47AgrqKQ8nSjxDG+WM/yN1KVsP
YzWexN939w/+W2qsCSloEQ7wUOzkbnzaPenvUhG2SKKQrHjk6cHBWp6u2qJAXWgt
Dh5llicdefb5f9dNB549pq7gN82ndqRDxC1/SXSNseAdgCHV3BxVlM73rz0FI2VN
D6xm8RCXR7pFVyYLD6eoCsYQrJpJFTRiTVAHH7pBAz071rqfU91fuVFmycjcQH41
i30PSIEwrtrajRNJK5Cnr7NLbtHg5ITiXgL/1fZhhETu1zXmL7YTTfhQ1Hs+xLQ9
uziNaLYtwIRl6W0gk8yMQDgDDApZqPLXHxsa8NpHviWZu10VI3Hn7/gavWVLWYWV
pMat8l5FXLOI60rCzSrnF7EEDDdUGVZbTSa42QhagGMvJeP8ufYgSZ5iwDNjJ4Hd
izKllYcEHEd5fkQ1LUjFBeKw+N7bYWTTcAA09nAMc3gTEjZAYQkBM+CGGGVmjB3l
tAFY0y/7AuZM08ZDM+44HOkqUKoyiWkmF7BUrtSW9BqJ+BNEY3BaXr59FuEtdmb6
dgoaSlNpJ2uP31DqwMbIy7/iImsf2YmVcsmUiEa7M52+T9+p8KjLtkbxcRmmC3Fz
Gvzdr9cHUneN42c5gCR7gaX1J9vEVPV9ODuOjY0tv1LaBIoKGju6UCXbdGT5J2Zl
pqeZJ+2kjBgL7exOgCjyse3hrygpOm5fXHKOM83qJ9Gu9ELZd2OqOsOpc3QvXvzc
MpRCvbIiSbHRN/C1tXYGV/Z/bdrFlAO+dYGmxG4Zf3W4xGIPAUedsU9s8rV+XbQZ
N2kW8BWNDpwmtm0F2mfnvnY+AOKp8MQ/gWjTC7qx73uWNu4/O0lLKOUicHYkhVp4
CUfCn1C0p+VRigaW9n0ppsG05PSiih2CK5mA1wO89hI1oh/qRlHwsH8dGUPfiExw
8/B7VvtdlwFaWKuJOUfxHABFUG/hfMoURxU9UiGuwYDbGw7Ga7/a1VuVI+31ltSB
5lUbMX6S+X5O377RZxIvc21U2LYFkUmKfO7H/Eshn13QvR6f8uaxsc/Lp9bEFnT0
BVBbaFh3VYrliytUbk8rgLxU5POXpLu7Y817qSoo0gnf0aZ+RfwE249jJetsBlEb
rZLn+iK/S+1Zlzy6gIVtCCpnFEFlRwNzwrQnpz8RcyM90gnHLiMQrfAiz4fORBEf
53efnRF2YP9i6bUhdmg4Xo4ieviQlRcBeMZkaxar6gNEPNLJ9E2iLWym5Go+7LtR
DigXukbqrWo0MhA+haj5SzChr9bL63F7rhTTIh8u51+LqFmnz1iwvwn/gmUv/ZxC
HQrRb8+J6ArLutd1vhk+ysONpPsB6Pifu6NHH2GURpNcBBs/sYt4pzhx1mkLyNpz
RbI9/wzMLaN7MUAEjHoWp5JHovRIFQ+ssJLX6MWcrM/NPvGaNXh9gTHr5+Vwpqvh
aVBXfBaATLPa39jCpEykhozppZPClP3wH7TJu9OHOAL7OVEWuZZ0H0jH2XDa1kQd
xJcUS4v8uJvHnxR1wt8lcNWm7WH0MlMkELduD5xgqqdMInpl7eFoX1FLOFMDeS+h
Oqefuvhck57Ye52EV/wXA40HgtDaeYhnhYb7srEQAgUpXM1xBa8x9aMPS4zgtk/i
pQ1hygM3f1WJL1Re98zpT1jfxr1TEiSBFH87A3ldiyBhBETetv5wPxZzBVey2+9o
YqZFyVuyfSZ2op6+pV71jw==
`protect END_PROTECTED
