`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gX+MYQ/vBGaQWY5cVV47Y4D53eieK4F5Y5H/QnA3xeitgLq13EIPnki8f1uXgKT4
T/n/sT8NWP8NBTWOO30CzapTfFzNxu3+b6FFXPplbmhG4itc8ZvUpqZgVzHRJs0c
65V0Ogum+Ze5Ilig8qYSoEwulF8NRdvv95ejdZl9RcrsYkN2FcX0ppmArdNjoKHF
RuU1fi49CHGX3arV8ojTaIIoRjXY1D1kMvZMFMhyZ1Jk9Hntk9AyzVkZHIgE5bSU
at5DgvZXTUxXYTCmYn99WgJmKTa3oF+8x2asLZxfSUIoPt5tznk+16GfEYlqRdAz
OcelUXJFMTrbwa6jZuKc5qaWdveI/OG0vGP7wyVQGRdxBaBDzoji6kULEt5xhOys
iw4rZmuswxdUlzC7gShvHUm8Bn7Wtzz1cuxmOKVJwSvBbkMMx5sOP5RzIQNdIDuW
glTyOhdH/M5/20fGca5hcqjnUGzNmd+1P6qIuMzL9HBz4QlBakpvP1zjarmL0NM5
xgmWQzJ5oKvEnHFbFf6N9Oz9FkzFgo8Eyj/DS7gScxRRb6Amd8y+82k1oP26ROyN
LT/MV4BL2PThVpY8CuDVFB7PMypMZFychPKn/itDMHF0Vp7MUOMqdKWtAW9nBnMe
h+p3NPixCxyV0mcuJn00eZF0Am0svWxxDwh/X0naJMxC8JCRuiHmjYAraM733la1
Ry6wt271NHIE/YDwFIbqliAHoKjdZxovZZQesFq8wjdvVvG2L2Z4AsVEbBYRMus8
UKcHvc2+9U6T+YBVDTH2l2r+KN0DV3AYC7McWPUg/TWrpQpSMeLEGGc20bQ2SShj
TjNTySd5CvfzInOYY+QjG2JM2RU6ai1F/Opm5gBLlb5c6w7I5LhABC+E2z1P92KC
pNnBkFsWrZM/UUuHj2NldKJoaSwYEnOClZVoxNRNLkYwYcztk+1Ooh9qkkbOdmyF
UMnlEqdnbKkJeKVAaZxMCKICFlqqqcH4wmOsT9HSfN0Rvee8osFyVophmGoY9Xxo
tdgNsMbyKzk3rgpCBKy2QHIqkmfIG5NNITigT9vNRER0yLLWJUfkSVDV+85Fd8GY
ojVe7PKenJpSmZCgyid4lZ2yyZIS2tIbf8tO2jUVGxAXXnkCFvs8BYg7a4nBsdy9
biNwuicC3yBUZnwsEViSSkIHIt/wmuRZQFYj/6UTshqeivPQA8yFyavUxj1UF0IH
wCC3plZDmzHL6vQpJTUHunQ0xQ/EOlVizGsfmfXXrfbknkFhqHxXsA57o6MPVHtA
JgtTyKj086ck0E7OHgzHRb3bwP4Wvc1VlXjJzVOlPysDr5avdRyd1YStZi+G62bh
rhZrB63dUFlqkdXmNhJcMM9pnX04IORFdPXnoV7pgCQnD58ySig+SuO4Y0gbpE9V
cc//V6v+0K/9ZeSeERHTnWjCa1iaWue7nwQ2DqxK3kAYemaXkBR/tSJMBhgsLdzv
+QV2nKCSuh++C4s5QsGnNsWlvMucPy2YEhFt1rgoigg93Oe5FApSgX9s9vp146+d
c3QxZU5/Pp3XalSpnSz1r6YVNHdIFteTpI8QD82OXZ4Qog2Yxiz9sZ3GsqTX7erU
QSlvx3l8hb1+nEmnx2WTYuzHgmaFej/qj58wXMTeU9Gr8eVFyMVMRfKsGxfe5YJ/
sBoG4FRkpJnqgU50AgvCVtds3Rhc4rp/abZgx1UiZcZlGpxxnsNP6GfyiRKIOi+D
qZNiSP6HVFHpUmMa6VPdbKBVcf/ad8ydCIrze2rc3E+uhuGS2hpFshMZEmj6gOBy
l23q9Ye9JUWZz3ue1VKgGqZCAvR+/PKEJfTj1P2EzOCUHw+5SakxKabAYrG6Hp4G
1iHBjTWJiUDUExulpGKcj+10SV1D+F4GpK+0uw2PRaw2tylvWJKVRic1kKhMHkkd
801iYLAf9Zy2yB/Ih/xPGS6baVsVDK5IXHmN0Ks3f2D5AQzHgU216hLQ+d/XE8bm
nXd+GffjOuNw0+yagB3EfDtWZix4PdJIguQWq37XE0gyYS51Pg6EFmPVn0GhRB9b
QJiQgrb9+ywwrJLUw3oEGa6S4s6hhM+ixKptfij1uYgGbVj26bjeosBNQGDxrmhp
obvZgBbEmBpRIN+MyVFYU9Ay3S1W8sS3yrfdP13C+/B/E2nE6FqRs5RYTlGakjtg
HoZoPJLZUkezOQEd9FJIKCGM5cfkTpS96TQGiKFBIBbN4x7m75+0nHFaHbrO7oDt
FsnD/ZLi0sBkEnN+6HnHXp9nyQ4e/bKUDJZi97k01jT39yCMuDt7sUGKnLd/7860
OuTIJlvDPOtCSaGPQVoDpjO9tDq+tEVzy/jK6NO/3yC6Ot4H2r0A/ZcRUkjfD5lD
qQnSy9DWwN993a6qXDFGZ+6P6QtqoX8Ou1tHVnpaz+4pCT7tn6+v9DLyQBI5VAEG
GgFwJhSmV8ZF7EgdzfN5a2cxgqDjM1OOCKD3ugEEx22UmXTpqPnRB0X7CeLAmDTT
SmcBh4N+ZAt3uqjCFpr6Jf//hNmoHO4xW9fjHIPSUl7dlZuJZ7h7eP0VWvC99JbF
rW497sqjcbpLtOn2aGVEslQlXuvLcvRB1FcxcRnRfPZpguD2SYHWuxx1q5oNGz5j
KgiBzbjNnFbCiOntl99cX/9UlTfyfzbOBeaa8OHvcdpI/fk0DAQGToDCzoZAQ+Fr
MJRm/CtkypUDzPUwgXQTCLJzGSOkam54vWMaL8j3xl3yXGblSqch74oCgUkE6SUg
EqDaq6dTAGpr1Mk9DzIYfzDeqatkbCanHQo9DBjVFhe3q0Q5mYmN/q2Oq1s5k2N7
Hk4Kykej4+h7agdGf074ddpy2V4wKFjAfjl+uvrO79Q9mbDaZu5TOQMPt/zS3sfM
Cnf7QtkW4tbMdRiuC6djpCqk1Q6x6sT0I/4NqG2371JQKspnE7Gs1+13twQLr7zV
+S6ZXE/sWuiWUigncJZLeBqKLaIL1yRKdX7gCHv5U3dUV3W6TL7t9hZc1f2SvyUP
AvKZKlGdJaT7m6GwpZj8hYayUdaBGwDFmtYexkYh5PCgpnLoNGFzlhWgLb98z6s0
IAM4paTzNr6XlU7hOwEHqHxBbz6yZiDAqjYFzR6oIzJZYXE1Rk5f+PWPUYqr+DLF
Zz9jlMVcri0AXbt7aykinwJp5VuUaVdA7PP+OX/3/Q5lSnE2ks0/28I7UOuqtxBC
BUaYgM/NlCuE9ESYami2fykZ4dFuY4YcUeGavzXdGqjiT+D7a8OLU6qvXRQO+7P7
QsLSgUYQCnZwCvxpjMEO91l1Klg9sOxxYBgVRxx0z3W1FZn0659zXZ/TWMpMYPgn
hhZRQt1TtNIcnRtr+lNb0B4z8UkCKcfjMLbHrSiZxNOitZHg1/cNFdz1HRNc204Z
lCMu1EqFjg1CVUZvaGIVgTzsqlYbDUvL+GZ3mPCtpRCJKJ4ca8RYdY9FxMGq71LH
NA8tsY+46FZ0JBjhRj7+QeZPJpvjkabvmFTAi09G/2qh49TxaFMWou/SiuI5Q80g
a9wEFs3qxd4gtQh+RTAfCiDmVJaLTnPskNDNKzo8vXpzU5vfXY7VlkJ8HN4CIFQo
At6lBIfjhVi0d1CHUpsrO/b6WDjsut6g+A05NztbxtJrwTXzrCNj/0F5uuHg1Wbh
Bfu1Ng5UgHjtnWZIe2W8H176GHcU0BX/Syme1GYfI8tjvLak2SvujygUsU7ujKv8
7OSC7WbYQELT1bpTN7lSa8kyRaRUV8k9DjeDmDkrF9yKNTyaUjZRShiTZoZjSS/6
3VwOSCHkMxV185M7LTmqQWUq7MsEQMbKJkBJtK8fqPsdWfF34aZGBxJ7bjlFwrMA
5tOVBHXiTO508fpNWL0vA536OXNIJ7XDXBwb2cHxMgLNDhLSJ8h0ts82TTkxzGwk
L9UTGf0jPavDCo5QbId2HFfaGijdXVeJhiBYKTEorwos9M6Bm4NHFZznE+0I12Rr
RTqPG1VINPCAVJXafUxdW5TSEJvI4CBLSv4MF0nW0uty+zfAf5ezNoPDBf60EIH2
FZTwtFm/NsYamLS3wVGsfCZLeBZuWzwsYQ7BoHPtCHSUEOe7EmfmKiXNYeojo1F2
niC1Y4SJa/gkaG5ZMTbbrOe3EPBCT2gFyBNSP3CLmjT7DyOsjcFjMwF+nzpat6bd
47jDhwaLt+Vk2MauGUhLw1LJ+4AQ2LepYNifNX/KumLx2GCL6/rr6et8txI2nm5x
oWTdVGl7ZHYPEg6OXPfNKEY5Sfd14LfK+HSAumln2TKH8sVDwxpJ04Lhib5u/QjR
RVaiSQMb2m61UYPO8rFTiat4r50q05kTEwTv4I2uwdCo2nGILTVaPSFflISeBQhz
42bMNGPMYXlj76HNCN5C3CwwUiak3dfSbc3yCy13ZdTcEpiG/xUjCm6KGW5FUQuT
ehKuBYwJsVTb4h2cKK/USxN/ed8dDSBQjl1PkFY/SiTga4yLJAHZamIBJyav9gCd
A83tNrlWXvI6FNZNtwFX9Ck23MGyJXYl1yOr5bIOToaRp9pKv7/2i1UtKUc/PZk3
Rq8zH+MgG5hnWVsxT+wfCzNAlSYndP765Q6K58h/wMdR0SQKE0b4LMESj5Bg3yzx
NIXxdLuzCCAl6R+HM6DqD5gOUsWcl1OIB0Eby/nFF4A2oC8pqGX2z6EK5KdobtTy
4HA/DtjZBWI7oIa12/sdGPCXscxu2TywIWEHDozvhZN2q4Apbi6tN2tNR9qILfbw
biXtOjhHLSwcP4wGpdMPl5Ibv1wRGGGZVkCvQ6P6HzgVpxHUVIjRZ3Nx8NAsDQDY
kdq5PTtJlrbk+0TOLlHprHJX9QrUdyIVqVTkRc/in1ia1I2XDlUSOX9A3wTGwdE0
PTN+B5GjXLOX44aCnvPj3rZOPMHwJ1ySxuD2OzOinJhSB4Kex6RpsZqfxLpCiESH
friYlKIXL9GPEfmmEFwZMS9GuMnt6t8UdriOilui6fqsdTWAeB/1XPFQGCmPMgx8
y8VIZMkKADTPVd4sDMFB/tkPKu9Q/3tc6nWCIWimnRLyDGoLfsRhtyXKd9IRuEc9
0aggY5xmy/Qii3upg9Brz47zzuE6PDQUBjKXz1VROehZPMpsVEO2JxCZU615qL9+
yfbgv1RSveK8YvMsovxfvJ3oE5nCRk/SkO6YVVyTT3dIgm6lr8FQGhL2HQLypPTn
RR/F7N/XVPNzVY4koq0gFBzmFrMz2cc0wypBpERsZOvEUFsZXnTDGR8fJW9FYT7u
I/lc8MAKQ6RTL+P2HCgK5kihwHrBHX3IrpjOgiqiqP6qR81qRddvTf3b6PkWS+wk
29NjC3zbctmvOFPT2wCdpr7Mq+OsEUudJPcuQ+8RgLUKeMGb2wezFYXVap5kBOm3
JGdEzaNT7P/6ny18YDvDu1JbR1dbUGhcoOlgoeBH+wUYKkpjz7hKwERMN5RYevzg
0PVjxXDjh6wCzGzSyeK41V85ugzqpgSfAXpcCID8Vdfs3hsiViNcdb3fpEjB8upG
176kLj8l8lll2PWW4P+lGHLPu2a22x66WVtNDu2ybjf7PH+XCzd+Hbptu6EK15+5
E79JOnnj1QeE8GeW/zpBSUxFjsmqC3W3rt5LdBzDwYxppNW50J7L7sAZmPJKtIlO
hkHddlru/FBDegKl4L6OT+h5IQAONwcgY2XHXnCAcAwvwk8gpm1MZlTLuJXVMjLo
Isa4lXhPOMZuvvcnkWuqJyF+x0p/MvroVdOoBbRic3RrFP0v61mgrZucK4/SUdvg
7EEtZTpmL26moJ6hlEpOEWMuz92xAjfcmSQqkBCLr0vw8CEgJVwbEz7iMwdjkcFR
CviObzCW0sQNFBUhXJhuVCKoi/8dFayfug9OI9BT0kN62XT/ExNwP17DNbzXK7po
h5N3sfxwFQUDjCI+4Q6p5H8ejifOUb+r9p+Yw19SVuZtXCHthssNViM/29w5Vea7
U+DLAanbRKJYGjpIM0BJYp7J1ZaCZFNB2TH7ZFsys3BoXyPeDpDhsKx7FJFn0a99
OclpOf1bAC5i3a5dHBnBAw==
`protect END_PROTECTED
