`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Nqke8AybFjpgwTl5/HRgO9iZYtCi6DvN/8RiJs3d8czL0+uLpuF1bfK/LFOcUhlA
aFNMaBZWeusldCgiO5QRi2ivvRZlvFn0/OUF+JyE62BDNGK92rpx9PI+SejBfwiy
tWzbCXayfdA9JrEwq0QxPklPb5A8IbHLpNDse3Adxw1fWNoKE+wulHpEjCDGWbj4
85DLZSfoyGKcz59K9/IbARaBsofYMQnLlLE/wd6gHH7ooF3t/3AlFhCufaldMpeU
pujABOXJnyAjt2IlnesSwVIqMrPg0BX+0cOt59+9r/MA1wQFtsfGC6e//jaIY6n3
yKCjdZXaEwO+hXGlSfplBjoBprZqWihv9FJ9GFgy1WYjNeIKQZlil+EBC60/OXqV
Bar+9K0ZJo28v4LMb8dxgc4oy5XHFvIA7JT+HP8B7NTepEf+Ze+OCzStwA8klw3X
DkBdczITrTgZr2BJDevTS9Ud3bmZHUYhBQU20shRcEMen8uPqgA36WuLyATwKjU9
0dWdmiXHIcl1aEOdV5tz/zRvBMsg0d/2Uv373KqBwJkO5VGQN4KHZ1GcGP/SjaFR
pACPcYIGBNkIG4OOdsQorrXC0lJz4r5P2h+p/0zTO27sRPfUPIEeDT6Ic2w4rOfY
s2kxIzBbOQeXouNJuNOXuLlDLeQJ9M3DzxOoPUFEanNx0Un6BJfVY57+UhXwVpXM
HtxWd5Ap99yFEDOui+4YKDhHsEiheFVaYt1HgfDYKyv1Yyi/fXgSDyvYO01nmf1f
dBcpgl9iT4W3xRBx6zUdp0g7mCOWjxUVWJqatTH6fww+LetsY4oGe997p7H+J0yQ
agflKA9fVLdld/E2mdznSg4zSD1Swn08C1ZasVenwG0JXAi1+6sgIkSONAKfH69J
P8wJzVtuRj7RTlNOGj8STtbHDyo4nL3nijZIiiMXJs67ImSXi25jzBy8TqcCU5Oq
kCSdCPzV/BhrH9UJytZt8dsbJobPE8MpEE6Onk6ZxNyXKCPLQPOs3S9e0N0rg9yq
sBFCvlZiD2I8SaP9IUUqkx6vckInuxfauTlEjSI57EfPGBuCmlhu/tK50PQZC+ZA
rNXNARCToIc2UCJa6Obc+o98PAZ+KKyorkWaJr0s4SQQb7dNMNELwjAtI8Vslacb
E8p74/fNxYfJPq8sUaDrUtwVagLBtZxk/xavVMkVyanHTEx3qYLPQZlEStaYRpub
50yWMqsarR2vOhsU0omh8ZyHnS4l5A3Ok8jEJYn2etpspwZKYLrHDn5M3IL2+ItF
SkTFNPrXfKbTzkfAkZGtlmzKYDzm1qPTXYiNeShbijUwGWBHQTV+ney4k4stU0FI
bEP/ARj3cxk8XO1D1qZbwwDHP2fNDsrfl2/pUaJsB4A2ea2RH31S4agCO6rp4Gok
KCaX5agoLV66qLWbpfFW35zIwr4bScEwgNUPVyXr+oPT5pfyEY2p66lJ00Q6Luhm
JY1N4rdWois1GZZ6QFBuHXHec+HyNc5HEqgQvcSGJaS7JVUasCt8PA2R1ooa5JS2
L5HABZKe0lbF3w7LRcIEbw8foEXuGCiWOoCly2KbnrmPg2BOKVaSqsfghdocekJD
ZLgNl2Y/mGr8ggm9J0tYc0oNto/CO42FMvBQlahc3Vy+76ANbsIX6bFcbNvfqbHu
tZVIP+pk8BKljVN82lSEj4IE1gdwDEKnN3GlyHBp52631YhVyl05pc1vuZ4+nuPH
WGvxgu+8rw98c3Iu+ja6EQiFqDe3HZwm4ZmmRaNRmmavZj2om3RNAWYhEC6HTL2D
3/aC4TRqQEZkRRDpGF3qrxlqgR9YvMk2yenIkMaHTz/Alm5mNsO4zWhcEZpuXV24
2qvo7oVSWa9+qjIfkDXYMusDXWATZDVLO2YxdeI55ueg6dsRI/xtaMg7n5AdSd30
CdrDDzIdJzXH6Eq+wmSuwqAXM/gxlaA3yq7qRDla/4WAcK2UTFZQXG0gjzEi09o8
Ut4xh9eVIbKZuv6UhCS+vA5a8rmDjz+7OjJpmU2R9XHU4Lfzuyo7XxyAE40a6qhP
ETKKgA4T3Cm0OUDi00QmGs4/FfxV7uyir2HvP3QQL8XiKpc+ycLmAeaNqX9Vvzpo
7vzzRMt1398XuH5vQ1LI5eXVflfGN0MJ02Jg4g9loLAAHL6Gt9sFPd4lCipufpAu
eKTePKfYDrGozutsBUcMhn4niu2JqaCj9YBYvIEPBCdws6y33RmJt9QoMFlFMmso
HpKaONmJatS/eWBrla9KJXJiAWcnzW8NPj8x0179quk4ifxeY2Jm2PgJQ4S6Fz1D
77ruRaQkNIoUg5MC9K57dLMLMs1DkfU7+zmLzMmyrekAQQDE+iBzZxgmTcseLZaa
LpUJiLq+j3RbixpL6aohni+PBKbZMD442WnUaLwBJw1B2VfrbQp580g4pUhFclPm
uzhYxNyc22/Du1fdcMBj+QBonRuUnDo8hTr/e25AOIpy+LTQRQ9/zBZi1AUAvCQh
rX5TbnHQsMhQ9pOeYJroZaD7BEglIK34R420RpQy6wjKjrFXb+ujBX9GdkQ8CqyD
IOtmHIeKQrvw3C0ezvqPFTmTI/xCJfjitSGZOKb46wTPanuJ/WtFqNsZhvJsrBZR
F/bbqdDw9dgsxAtS3rAG6PA82+7VqV0wkZxXl4Rk/+d3H2TzbRg7r+OXcMy6fVuj
WJGmRXB48ICgVc1uRk/fTgARKJUJKVJec/Ee9kmV/JOjp/O8nWKaC+S/KbbOKWBW
JZqHHaQ9GrroUjDfBHWthjsihGbDDPxcfPonLAhA+2BwZvOdPqU7BgSPX9+EGvDy
TwSGrSj6rC9IZkWDclyVKNr+HhhqdK/dML8/AzlKwXofWUrpW6P+ZxjhhAMzt4a/
GKbR+kWD/GAXhICq2rLy1W1Ti0pvrKOmjjjcVn1YYd39xIRxsrEtMBR/5Ax/BcRq
3mN73n45fjF+MlGUsXYX5m1S2Zpz0L0rJJ39lSYvQ8mNsABWNAzxtlFTSkbaKTbk
OtNgK1mYirP2nRqDoEJtvH1H1TkyzbFHTjB9wQ6fdVr65TjF6JJTEd8gr0N4M2ej
i7ZwPhP9G3uicXkIiKYG28gIcP8C0i3RLUjdOHTyySBARRlJ2o7mIlT+rmHMK6Wi
yG4jBoxQs+heVg0Sc2uyKqFq/xJHrS8dJSYrzAkZUP/awRFOua0p/+N4MEk9dOOw
VAaZf0fQ/SDUdZp8xW48BZTFI/j4TF5pwuOI1ryVNY58ACv5PfZRLZt6AX4wxyxT
cN1NqR8PLJc6ewtWhD/AXAv2BU/IIphB/5wvQoHYlsWUw5lAKpiF8sZLpQIU0pV6
sn4e4uuRMd3saRfMLII7tr0Uphj5GuyYcnf7pMtLgdbwikwwxxKT5I+M2xHmvWgW
xNSc9sk1jCdAjayLoVlZAyc8QoZt9Nuw7aTmfBlHKCnJbiWVFGYvuSKSOPPgNinb
1jURBk9EzlQLOq0V7h1qgWXwGvXHLLaw09/lrGnBaNvPgFHHu758k9yKoTgsY/yv
G29YSLJmutDRdzxyhzG22DsRbhPusOO0qQtOgXs7gBV8S3ZU0S9IRDXt2aKQ82YH
p9+Mn7kMNN3hwskNeIsMTwlA/egEEhEzrt7mv/9lN33EkbKkVSttfPAyqrMLnadj
zaiUOH9ann/od95jx7zj+niXO3UqDRvkTn4i/8S+AcMwGBdXlNUKBYgZ37GksNM2
sgiEPrXzYeGy0t5m7i8U5gnX6ZOuJpxrkpWtW1Ti1G6/vQV3vsJ5qxE6PYymE11Z
bkCuA1rsrv5mkwR80gns4P9YlZ3MRLb+Ka2+tA6xJHCxlLiT7Fr1Jk5wQQ7sQDDJ
YeLfbwrTk6gHU/t9EqolrXUz1ss367XyGoGthqw6FcHjgaEsZXExoumSqwO6Kkik
ju2CCCk44oLJhRi9vJtORK7om0y3EHjIzcnFWBNF2oSKZ7n6bQhcQv/X0VEN1TGX
FktNdxELolkpVgZ5qSRDZv754rYHaqcOIn2RV+FMG0wH5Ji/Wnbeopx6NUdGgwKy
zoF0yh3ov7shxxzOgYTdGh/Im3MzXchzdPXgCPInuUbvR+XWAHnMEGkOH57+p5Tn
QZIeOBA6LJ2WoXu8Ml/Jl4hlEPxRxdIOiGsRANtbOSuXRyBaMtsLmwniY9fHlQCQ
e53fJ+puCu8k8KYrdBSB7DfuPfqVaIZwhG+WX/i3b6W0cmaVj5VQPlCALJysaLsu
RkdtVt93kAMDD3WHQRnt3aKRShNKRZ11HHer0VHNeBvQ2kOKn1DVP+jXskcceS/B
Dc58FaMtybOMLHG0oQHPZu/YPhLzSXvHkcvoC4BU0Dr3gaSYJk66gwSDY8u0CRVR
p5raknkARlf6NQOYMQJ55WpsnnH60oec3R+4uOnsOYwwFkjGO+iczjt83nOJbDde
hmuTO+yufphTOSDkjzVgkJDagFucl9X0Sbqh53ac6TC13zKEJTOWxpogHD52Ww7h
AJQh/pYx6DNjL7dlRgWO5keD3UgWzoOMcD1TOjZcrT3FJ9/mUSZCrKyiK/2MdDZ/
FfANlgvstVBfd7zz7qWAGdZuEpmUDhSybJZ9yKYq9jrf2mmu3f2Pei+/JL4Poke5
3f8dYr1GtyiVB/ErwnLuY6M6Nd1QG8k1HEMOFSdQlaJbFG3IaYfAhYyDmLsHUU3G
4myb0rQve2iFAVnj4pJMI4+bn6b6KYh7KXyaJGxc+hgP6s/Qlb+m1l0QI2XGLU3P
MRz+dsD8r+N8woEcxQCsoSk1TDk2TqP5oGaqYfUbadXTL6pJ4u1YJ2PHvwBUoXZt
rsL3Mj09+tRKdXC8HIFC+wJQJQk463HFu9ERNU7pt0xoPOvatAr8BTfAbNXeyYsQ
t87d3lRbklsgDjixR8tUYmhztNyw6IbMH7M44JKRXzSJxRwWjvOMN3OXT+0gXz6Q
v/gNYjlehHA1DlD7Zb7QOb8tWIpV0k5oryTfHVCL9b8rQlOGTORke176FgtLyDbD
U+RZ39ogKjFH6EkXDAaaJFRiHZxIVOQs0kzTPGcaYgQhzx2hHGkGPMGpBputvDJ6
L7TxqakrYGuhpdAXYF04pEEBZiVto+oHXRyYyrRFt3zPAybCca8H8KSkD4PcU59e
qUtYoDniUpTnHuW5cp4IU3Se5fqHUS8aNs8OzKS+obfcZnH0VhOiozAs+nqFohrM
y/z0CIRsBZ6DEWBRF92kp0MKXOE0hPd2b3uK/gUncLvvbZsjAcMI9hIWLtViBZlX
XD/ozxAzx8veJKXVfkrJ6nG+DJOpf0Jss7ucD3Fzi0XLR6t9JUFT/pEAkDcjHM3i
6/hS0rV/cgbgazGjXdDRRtuPL8PfAu1S77Vo9DLIp1b/Bt+4dlS2noj8v8yTsh7G
+kbui0Mf7CkkT+GfkVGuxm5gDKb9GSL2RhOudoyMJtZqskgKRnm3pxzopQG+5SbB
ATmemVFjhb0Yxlf4RSxhAhcFO3fCO/F3TSO4ucMVDVismHPw+Rde+C5CkvO39wMy
qvk0S57Grbl5g1M0POCxgB/GCSf/RoIQHalaVjFl3L9susckILX1E3GQwaQ6gCGn
y5xI19m4/g5z2X0+ICN0fiJrsq8iQ91IPempmfkN0I5bgqbQ73IfQrevDgmazgBt
4k16sH3GG0FJxaL4zbBfXjz3V2ncevpY1eCX+F65eg0uS8DnNdhfgqFL18GS9Dqy
xSw1/dMYN+BWppeY3xULK04xU+TLAngIefJM9umF/ssrrvt5OYYk+BcCD8X38Iz8
AGjAxiMhi1lfasa8D3GruoKhIzelMcYEZ9FExlAjBpdYs7o8O0XASs5MmgY/f/4y
uX92TUHruHMN8pOXSSWi76JDt/k8VwBG80X2l7Voe2ctFpvMKwJS0OvBXayswEt4
NWkCoK2xsvmxB40+oKV9qU7Q1HCJLOjBZeIgY1AVUcgcTANnrEaEoafJAHyJulvW
yZnU9G3wTJ2SJkh/K1l+DB8c7nXiULAvyFU5C6me/L1iHK43JkXnbMLPEmizIrIe
ZPOBuRc6kLcZNW/J/OaXVrhHA/gMEN1xGft6wDVbxsHduMvzBAqLkTU6HHHGEssx
gOxu/I7KOxkd0bD05XvRt1l1YqAB6+y1p0PQz4yApT1FjDnYEqxdxIkSFd+TbTao
7WlGQC1da6oOuV5PN/aFdE63rI8LBQrOOn6QRAQ2DIvLnOQC8rP3lr1hjg8YaPhI
TE6PI5rh/1Y9Su956dHEXnY0WEMWcD3v3xlqzZNw4xVF1s+b6jz2ILGAZLOVpnfE
1DYlbwOK28hOdZI+nknvxg1S+V8LHfvFiiBijx2La7X6GjC/M6CrBtl0l4+7TwGz
pHjR2Q6fTc45pn8pf6QTc/sX5xQDLZMI0mA6yKPSMDX7J73BJFh/BYQEFF9fW5Pr
xAPNtTCYBPpVsqami3GxaaIhJjcE9xQ+tqxZsiVXuh5liXIv81a0TuUKgaItUeTd
47mts0IDUk3UpdnZ+Nw2j7iZH3lP8VjBk1jtcnmMc2sjaKOfU6OTaOI5nOb9c1jh
F/S3RmOTOJjMyp1tB4w5eVCnGSBFbrNiDNbv4EehogaQsZ1qh+lsxjJT0KexjB+Y
Uh8Pb3WBgxseb4VvU0HfRz/G9pkWWo9Uw5UJMPMaHNWb+bXbWxjwsgWUAiiTFDEj
fZTqpmhnn7L2ElqPEzQsYNIka9MYmmKrxyRqPlMoiPhlm3PM4KsktTuVRyMPGQot
F/6lI2diQ812vusArg5SikADFlGiHxFbLmavOVkXKTXk8x3vegHxGroH0E4mR4cF
0QDCe15iZfcz4ivZtYLrOAK0hWhZgIwDpZP7A2ukjPKliAJ4e4LWp7Q/bRXA41tR
SfFbw34dpjnh4cbBplPevSk6Mz//pPmCyE1SU9Ri1f4ZCGdNVGqAuNcIl08BZbXZ
1NgyS3UHjtirmeEkGYSwbNvfH2ECy3Dv58BmXh8kc3fgBwkGC9+Sj1U5YGfGG31O
P6vmDhYpPGcHdxIX2YBr1hoI59moiEeAKzXaEdVxr39UkgjB24T/NLUwwrUWUkOH
K8f3GshCXhScf9tiDf+qiUHMifqXJqkOrb5kZgMltpSXyMH30FegZzx7u69nupJe
jamY4yw0EUBq5ZmfBvWC5TXBFgS8y6rGdBAR0o/VQlU50A6oaXxKcHdP8XlTZoVl
uStoILqRlMBnNufdMsUW5i0ng6AV+x1LiHonUNF+hRVIAV6QL+WHvafLzJojl/iP
As4MqNX9eQmNgH3gd9vPVcc2DLBTrfb+w9DB5Bry43ysltedmU4pu2AtlvYkOyjn
xl3tZroniD5/yTZN8KYraGxBsBgL2dZBUMd6x4IJTvMLDhjAfhsmr6ZiJttqmfRB
0EW+0NroK+XHaTEPjFOI6Q2vbFs90Jtf89e7/jjwfACmuEDEL0eUCy9Y7uJ96yZZ
ZMUOJWZIZwH0VXEbCTmJZNmMmoU99dVfjzsMVYnDzshmtRms61AK9A5KJNUa4dGp
j4kiSkzENl/xsWtSzln2wWuT9qgJ1UGOkabtCtbgPNuroqrHPGGJT5lxxc3A8ssA
2rcrFrrgQG0kybqyQ87ByfgMAkJAhTdKKmK8PkfyDBlluBSawVemzaVwJiDvDwyS
IQklo8d6wKMN0qpo7p+Z1H4zVjsKGn3Qu99SRqj2Pe/ToDCEfbkXapir8xS13guZ
Ko5+UFMAznjb5ZaKCmnT+cmLx9epEgckluLkhpfMJ6+nGDCBfYWFN5/0L0DQUP9V
Ir55IqS/AOL4bCOeas06exJVZ3Rrjj3AVC+xyNvg0stXbbYvpSdip9QAsNkXO+ac
IAG/+rz8bz9/xk/ksW0xocjxF0AHPWyqWfe2DGZilMtO+Cm8bmZ9JOEVsCrsH1TL
GzzhGa8qGeQIEFckvoRA+Rsu2jdyXnH5UAFMmZtLj3wEmNjckf+lDEEZ20Lfj7ZR
J7KSV5wvkxD+GoUgUZNpubnd00lF6vjL1rT9q/1ecJH98vvP2OoOQqcdKROJucmq
H4AqaXzlL2mnoq6Br+xPIBUDiRexxeyC8VIjzjCeO/z6p8JgSeVrAIxBBwzR/PNa
yiF6rMsOwedjM0tFGsDxgxqjuFGHQICJW5qvfAJ/5mJGm4sYliQ76oeGlMoeh26A
9BWJtxv9uzqPmLo9vg7OIkG3RTsD1t1Cd6YLuocS8Tj8XyAblnnCn5PZAW3IE8uJ
jD8e25VKO4jCfebPQmjeGX1NoKZoQIZunDyFXrTJo5PirokpPCk1Cz1tcRmAPiTZ
j7rUsSmKt1HXB2tosc+ahSrquhEud8iwwKmTR00x8LzXeLsrcGSbShUSw6B0+tQk
Kp3ztN5LbaxJWL/DZ9R7I8f+VU99I83ZQeQ4Kb7KgOdonWc+ivGeA+LXN92VvzYn
1xhpBCGgUzWTBseFuWKeN5VDdCinRwxpul+y9nEEVUwkxQS86xOETAbOSHDr6+c5
KtfMEb/sadUTEHrs85FWFFTzDwnZMObiDtTOdx8opoZNF2wiNVw7Bu/vSVgyN0NV
s4N/laXEibZB1R4QPwx3GT/RT1Lhzc3mHV+YyTxoqSvJzT/yJ1kXJKwm5YpnJkBE
2dJx72iezcpJoEiCoMjcQDZBEorcnegaxkJURzqLGkP7Q3Eb4qCIi+x14wfnUfcm
c88Ht4MqKsyq8P5vHbI73VdXjYOyTEk+pS5/N1pn12M1HpqmJNcmypkY+cxVPfh0
uSwuaha/ZrK+t+ptsr0oA9PYqQw/t+1knI8UY3xPNOD97Ts4Z70HJPgUXlICZnEX
W5pJQXnEBorh+CTXVSXEi/L9kLlMOjvgeGtQjYnFLOj3GV0YSJN3Vum4j1che8Qy
hJH9/NH823ybGOjZlhpqDsLV/AyAyu4l1FrNpxxhN47Lo1rM2ixdjnCo4VqrpiWx
W3jPAtF28d2IHKq8TsN1rgwzxVpVmym7buMaqmCIZMegNnGCrSSavi/Imvh9tLXN
sV7Kl9tp7LaMJGIQWnx1lrScxXu4OEPf5EdPs5MpVcevnTfzBPe19oH/OsTK9g/K
Vw1E/S1n5G/k46mmhZRsp81oxnqIeT1wemHPvLvgnytqcBm2S6+Y3jPKnaEtPnfa
JLx199KTyUX7wTu9vjX+RLSBcGDqP5+SER9H9+/8hr8p3owyAv5Kdv25EwQWwYQM
yQfhikxIWS/uaU6iUvB9c1iCMAS6vZ1p2FF3eOph7RSR8i6jBGCDcYurgFZcjBWJ
34QmaW/B3guBhOSRn+1z/FcZXCeG1lJaq/CfwPjL1Ci2YeVtIGESrnpbX42awaYg
zBBbr8omBO0w95W3l0m1d5T0hJ9Uwe+AW1EUYIoUPl6x9SN3NSk76jG34mUBywp3
ExLs5hOZBnaEced9E8BpDY3GFGkjOTxFrq/yc9xU6LM=
`protect END_PROTECTED
