`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bsV3l0UFQXsThqeh5m00+3Nu5s1VYZjNZVmjs33YYOJIGfxFwhzZLT0TIa1ZZmKj
+VMrgPyKy6n+awzzFmxuBokZrsyoh0e8shN2kSZ7Hg/umgsYBNfu5b9E5VvkxHiw
QjVyoQRERunBOuJ220DpWoUjAX7+sjaW6N3BOK+Wu7oeCwzkQvNVdF5QmBbs57za
5U+u13pwLAJrfQcfcrGy+PSKccnsAS03pihewjkmYmAu2zXmMYxHKo9ZvIhOp3RF
753Mt5AuuF1+ihq49CqjDiKOWGNwjqqZm1cC/VkPw+pvREIS+/PQq06raGCLytOA
g9QxdyvM5mJn8CV6EotWFz+deM/pJqcfau4+/dOlffkd4rjvzpIo4Bfiag7y2Vya
quwJwxPFAUPEE5gEgkXXsV1pu6AwzACx1dwaf7VYKmNOlet1OCGTm6qpyWSIwgNI
OE8yoAoTt4Rg7VlOQGNwURtSRsi8ygEEEqs8xWcg6U01qCm1EKNp/NBtEPMAP8wp
f2f6NaTGOV/zhySNCNhvUjb2Gvaz0xRhQb43jwvNx//dbmBHFvwnjxGTro+MYwY3
Z6mn2Co8tigHuON0AjEC5NsArYZqtcfjl3KZsyyHZZ8MtQEIKexLJAd8hYu6/3ek
LWLC8SevoTy0hTYn+8NiZFNeHFfAJYdVE4YlNGuA2MbasEdSiq60x/ro3dKy38LU
fDJZfozWhvTw/Kup61UtKeYobJLaFG0pt4tJvS3JSCf1Y/QTKBSK1wb/2bFayJec
kViLkrL7yAUgIR+aWQzz/bHcu8gzBHhOHZfh7EHe6Bns6wFSvtKodVQzELd/g6X5
feLLBV0oez8WtZvPCnINxWpEn1rT3o22sqRozTyjtly6hBWb4oZ59H4c29GRNaGL
ybnWXmfOew5HKUmve0U7ZSz7H5SPTNm4SU8A4QuOhFnnFLrowuygaqxUzaD0ic64
aFz/mGfzM8B0LWE0+nadzBGf1SvaA3nIx5xOY1Jy21oxKnZLV1r9iEtHxB/r/LRZ
3MStVuOAuBJmOV6BWxH4YF1gyAyvOhLRq/9j1kGOie4EdkWXQxFOuWsXN+02Z9sb
r6xazWfgbM+YL77B16bUE11tM0MUedHlrW4EuFTRUDSW7qesR7MH22UME7cxxKpO
PAMSC0uyT56axYz4pLmTB770zn7h8h4Jyz5W/3WKXfJtKa3PJL4LhB9Ki+qHdyfS
ZKR7guD+Veys474T7G7sZ9faI6FKscA1KU4FrmDtuAoTRKgzrnyKscgQF7B9f5gr
msXHHec0V19j71S11i+hqwG/hHZuUdq5ylio9PhQJFcwH9WLB19w1ZnVs6QHGkNH
thZnyeX9fmm5djmngVyZj+2ED633/BDEWojMKmMRpuaGlbm3zp9rPJ/5TR9oTaXA
aR2oagDFBiE/NvFstOj549hG6rPpcMaCTauXFbqyPM57+Xzy3AJjgUlz759VtFpj
x6fiaWoihtsIuTp/ZP2IqzfIFPbbizLNz9VgRjLUpaZ3q8NTb49JeDjbvs5YnyrN
Al1Am3tePS517NW42lvqTX+u8kRKJ3ao2v49J35ycjZBn+84KjX+IamzxKQAXr89
r7p/uekMdY5NLfbqnoCG2N/PN2zLn38x9nUG7DT2lLDkiWMjFLauby21lzuqkjPI
oIxcFSqnPtfyoZ+R3pxhsNz4U6mtXwo6gl9TxdzjfnhSuHUZxr4xhPX98KgxcIJB
P96b9hm/fEyaSM3Iyq1yLhiVeSN3MZXGU7aj6VkR3oTsminWvymiI210LDGPD9Bm
haCkI9KES1qMzCLUgpyQHP+oEtgRZ8GCTx7905khZX10AwI5aX8Hae7/UCx6RzeG
N2T1UI9UsQE9OupMfoE5ZFeCW4qjE4+zzkzjSV6dOCvXG4Swueg4bY84u5sIhVZv
JWelas0xCao9MgAstCYVekMpQf1aTvkqzJfaPFY5PXTOXXdDKs99WXsuBlS6uRj9
TJHU+4gMOj5QAUv4TSo3wkVb+eFY7dwnvJCN7z87DZDmPSQdw/3VSHZC6Xe6rQDY
aD57sG34uMiAsZ2BZ46wbbLRfnk9nl5yX0l1It8UKZEsVws7Pmzyz/rtMBwOHriD
tzN54LPsikJDJQ8l1pIO1PCGWdLaR9sqj/GbhfWpSHJIN5ZTX3yv/DLHlVohmO2H
XVq2XCuZZ0Gu15grBvitBBUaW5xNLV+aCXiks9mS09CH3g6W1rZ6MtpwR7zUH+sV
PNWy8mVeulLF7NPqpP2JFJVzaQK62uLhjS3QDDRk8Rhf9WJyb9wfxURqb5qXuEhM
d7WsW1oY9QSS8TovSLE7GmBHRANSqjJtA0wyJ2V8NhdbyKb1RaUia+tKQ5DNzNBt
6tfznCsT08N/Si3q6vyiIFG43XMzB2m3/0tmmP7oeAgayxtf0dWD/Qa6AN1ssZeM
TOOyu8KMV49V6Nuphd1pljZdbLVzy0ci1nhKgT/GvDU6VLDdcaU1Y+xysD9PygP5
UY2fuxH6i1X7uCfrKLBO5cIx/SWJiiaqAC5nJr1goueyFX4aaYftJZm27JRYCTEK
kYadCl3QBF1xAuY1DX7sfw2y2JfNyIegai9NMhqDL26vOFYvFyu1p4lXevpSI+wA
kGDP7RFuCXSXMYHfd+W2f+W2CuTh75JY7+Nsag8EOytHvBayN9oxKprcdw/EJMjO
ZMwHC299Ds/KegJZ2rXY6MaqrDo6kvPIJ3emnsTI/oHw7i+Ww8AN4MKQRj9dGBWS
nE+hb/n84v7r5SQb6HRs2/RUFaoGcnRlIXae4Jy+Scp2obImOaMSr6+91ACtPXBF
6ZllJEEWCIhiVdo+O8tEgADDDS4LTJXVpW3Enx/B86s428z1EVDRmqFMUIFv4Gco
vKCBNfQKR1XJ03/vg6NLoKbA4NV9sifPor4qOubctjE+GHq3fOL+QLsRtM7y2qsu
mlWsV8M1uzyDM5OY1Ga02xvmDu4Ac69DZIdH8OIOupRK2NDIZXSlG3Tqv/9uav97
Il6MeN3XzLkxNYwBX2K/Vb3WVbMpdySxXpoXw0bPr8KTFYMfn0hZvIxeJw87AIj/
DD6ANyZAen3ZV9mfNnKysTjjJEHmtyCDZPjw94AQ+ipdw4K5Mn/nkDteRwuYcu4G
cT8tqFVxSL3Oxr24TtTprk6NoeJHTA7X6Uxd4e3N+nEhSYd5DTOSjmHjPH1U3IOS
NQvj59oKsf47bM6uoSy2sncg2bgAxZ2zU+RmZXl4Rr2FiA2gNB3qIfS11wQshdnA
0jlL4CTI8/Y//9LtlnbWxQywZDmHV7rmGLBV/gPPAanzmn6WhRXVQ8dHTDmpp8NZ
DG66fqs4uHzjPmTF0KufGMoQ9wpoL1o6kWA2uqtKjQ1VtTwIy0eEc+8GQS8UUUeZ
QHbIhzHk6bqzna7t8j4GA+TTyodhYWm3niGBIahdPuK91Sy/Bl2K+dFnHyMrHCcF
vSDbCpX3yLmmZA8YFl4ac+rj4NG+ZRDEeNMpNqmjvSr2IrZnVNmrXhpc1mqG7R/l
R4CqTzt9mmbHbiCBS8I39vPpn5f28aB+8tYe+sVdUxDGwlmOJFS4rgI4KH2VDo9V
jf0JfKnrNvGZYOdDCbefQc6GHkPX+7/TShgzkw46KxL6v3ohgiInc1poWLRzflsq
S+XiKJ70Oiei44065+1qgduacQtvFTtAxeIPAvdQhildrpxscIeHYy2HsNtD9sCI
AXEnz+XHxfs8anEsZ4i9vejEFGXHoxecCKK0XnJKv70gx3eldtKRt7gqYOc6ntYR
MhUXTlUcpJSJjOD60SjdYiLMz6vAUNmMHoWSzl0XZyqJnv+ZwuI3vHs+Ew5WE8Rk
04AlWpUj7is0Ux7pA8oq+D3Z+MusWauOmInGCw/HYXE6LcIqvrAS9r+xKgVxrPjl
KziVA+LITLvoVJpK8dmfHX+Px3pr4e6GU3LwO6BlnoqsxQ6Aq5v4cvCXTMtcQeFc
0vtAaVtQwqkn+cZY0zIjchK4M1GwLBh4ns0lZ39cQ5nl5kUBrbVTgnDcn9qvvPvb
TQv6R1oOCQyMGhKTGqtPPhFGm8DampAoAnXyV+cEUi4bw3rHZrnuf8Y6SbG+TbYc
TqA1vnGhX8rqeDRAWuFgeQ230x+r2C+KeMPtLjQ1aj/aG8V4P4oH16NYMF6R12WQ
cyOAVuNvVpwxpiholKPSrYOhEp7xkb2tz/AfB+dPvD7Ejx6tZ05EwOaSix81MIAz
9CAlOqjRbxpwJEMFNhY/cG48n24NCQFF6WoSCde6tM0DGgxz0SAB9B6f0KPzRgPQ
ict2A7Xtm+sX2g194omThCGVfFUbI/Dk4xzD7qC+41xo7ltRp5NoZ04A+kN8bnUL
45qF6bS6zimkmcGwSYB7dQ2tgpWCWHjEB6quBvKnBBtCiLsjKgWQ+quXPjXaPWlt
NIxtAd9j02I/Rg+K+cEA8Lwd9LrRMjzHgcPvmXy7Lzcn9ih0wH02xFxTkyeum4Jn
7Ro841ZXPdBdCSzatbFsl+Kd6oXBiieXFc1Na8lE/dIEX6bp97FIA7QLZ77kCTIj
+vm4LMn/CtI0eVzY0RwsJykfYXjvWOSTfNJeAHeiECmmgUfg0gZbKDLJN+JHwjy+
8PxZiYYvh15elIMwenF+cA==
`protect END_PROTECTED
