`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E6WHUxUhkfm2dnDoUeSq0nPbyw9zLrAffybP+6Ka6lJEcl/ox0mbTmtKdjWdcXSl
y2dEXWTq9IkB/IgBboJ441WgM2Wwh2XPBiSOXHZPsSDkdF81wKTCcRYDTOAfkuoU
D6pW2UKcclt4i9kCpNN7M5qym1VyjtkZrQGlb3NW+HsNwcMU7tcDTDMvmpP3Nxlb
60CGxCslPvxQMEGmcJghU/ChOa7cbMGDdt1NHWuKh3rl+VbCTIEh6GeEOYIlzjwo
ob23yPA995PqKXu/HG7i7wlrmm7JULDJqKjdFsEbn5hEPgZ2R2MEbRLMslxYnuGE
hdU6XSBtzFtJvkqXqrcMB0Uhwcm4Rko+Fm8jZOOSoNlsz28XvdzPkVH27Ubfw9xn
UDa6yGnolw4ixpWyFUfTfiTFS5h0Zan4Ssav0SZ1hORU98/aMcJn8uvEVtDDDIsa
sUJ9RSors8lp76nzTH6bYEaVJ15G6IJecNYun4VGDnn1SFHFPwIZtY6XX5NlJbWe
RFsB4ftM+NgRaSSrz/ybC1aVjxoh3LXx10gXHnfgAjs5487aJMffsdbZP/2yTyW/
SDpdhvjT5BllHqkfE0HnE9q2dNFO9GFzVTQimNYPGVGnrQJ9+i10bMgNfzdD89Yp
b5semLI9+uOR/g3kakL4ZO5BMIsunRyXSDvlTzEsrIFLewhQgRVyQTnZ0078QEwo
edGbZ8aHYYkfyLgA9bOd+PIDIDqSnhJLQ5tlE6W6QaSiq8oardFRZV5wW8m9VTRd
xy37XiTf8Z8ZGqYNQuwpRm2AhvnahqYxQNBRF2pTEZQqwu4jbOlZIl8qpWH/ndEu
EbQHfyKn4QFXIalE4PZ8ADsIdUAfje++2U9oiTCRZq0VQby39OSKp98ZK3sVTEVh
BKBLj6Je4LluE6Pko/kDkfOA+rcgiMGXisQ/Gyajx7fK9P+30EHR3FFjZg5/bJZ8
M/v5qM1Bt4ROJc20kVpJun4Gmx5i8aQTjyRgDhZ/fsTAfcIz4AORYrY/UNGHr2Hb
bEel+d/Zty9Vmq7ZzUOiftF+tCoWeyNGFWRwCzpDtanxxGejJQ/VQyt6mK6JwW0x
luvQa2NF1tIXlqBMFOIqK3fSxfv7f+SSEAbHtVUeftVlwQupiS2m+adulLtbqcB6
6aK+hFLcO6eVRLmRqRcHsXyTGa5vbBT0DliQ/6Y6gw8EqsIHgb22sm9Q3bMyuR01
DA21kOI6JTWUR90V9IUmvn3Ewg3mNfMlL1V4B7mWgcKLM7L+t6Da++1lomuJfmxL
WIuSWy9IS+f3a5LGyD1a/JnFPVAkBLGUlyuqZbt6N0XkqU2Hfbj5uGBmYCIzXY36
6bdTyTUbB+QWZrMEtr5jhhVxGqgSJ5OND2t3spPKcEY2ulc8G0WqviEFetVMjFX/
+Rsf3C/yKBXqycZZx/l52QJmFHq2D6c7zup8mYmmoJw5cSrf3HDvDuD2iBYJGDsp
wy/aGEvXIykqpng55HeB5brwyc1gIs4wCBKqb6ca7iD/urIYQ73604oUYcD9E34B
LlTiKBIY0F38OsOuuVPKNSWCoTW9XkmQ74QpLxRbiBeY9AbYLFJwLfWIoGoaVP0h
090+n3Kt+B9C0XE1RJBEfGAgAnvDXfiMgNC+llunywHB26+Ahr3/9Z7ABUuifcaJ
o8eJcUAO/xWfoo1flYO3qOMJiUPtcORN4qVcbuHC8/gWmFk+/pop6hwGmDL0mPhm
qPANiBEre/7jIGsfdndSVIVJnHKJwiY9LzUnJaLPKaJyDbI+H4A5NTCpNf0v7umI
2pwPQ3hUSYN/8ybqgZyhwpyeUKOFx8fP+ZurcqNAHtSATPqIwq9fL9Rttwf2h3US
OW5hhmiIrZmad/kUJeXqpOkZLnbpGBn1e5z3HSmz20G5iTzLyedySO7T02mVzHt8
dc5vZeBRyhV49IjQ91cizqT3nBhES1xBvOTy4z3921vlY6LS5QWUknNzfDpD+zoX
fVHHSPRopdJW3W8iwXH5PXmp7aLhho0A2N2yy8DxteFReGOCwXxbdZde8hHqa12S
EdVXzrCyQMlcYhCi4Dsa2NL8JRKfYVXyGS7D9kSQjGU3dRTElFZtaj1zpmlt9Tzg
7KC3es9VN3ZFYGzpwCf6y8dBuhPaBGtcAB7iY3MmTnKqJPW7fjqwQB3Yi7WZJ/Uc
Np3fpksdf6sMPVSUrDL50jngcRSLg3k1ruzLtOJ//yBUBbNW3kDjaD/cWxbhQIeK
//G678nANuBS+VpkW34rnsfeQ1KB4DruDMOUb64MIxArPqJT73LwkTwiOZt1XNz5
0qiWqLhpxlQAAQtmRyPWe3vw1W6uNRVOXjRCEXNN/fSfssuk6PRgjmw1xGuM3m21
a3pnwFPjXWW8add4B30E4XNpa/i+B3DG/Z11zwIgVOR/ZsfKRWgwCbAwsV3ZSdlh
NpMLNTC1OdfGWFw25rf8v9i93ecGNFxS6s7c4IBbwd9Tuy4NiuB2UlAhhTSAIagn
020Xt9PhPJlV2qQ07TSWsNclG5bPNdwdLWTfAl7xO6a9nRtACdbJy58/JpTSFE9r
IwTA1Bdey2dQsxLv1qYoKF4+QTpFqF0ZCPw7Iu0izjtD6Ee5AieeduAX2cCp4xjV
d2ghH4DzRHyer7LrEW2Z5TF52eBBKwZUnNMpRYHZoQXpXRv82RW0cR0LaBlbaYCy
3+56ioiwD9eXMwXi9y+tVgh2LoDXMUlH5DHfY5hsaebSUh9w7BSxQe4RJYV11A/2
YwwXqVY+/AGuWhEvBpBhAV5MU90hryEoaC23tkPhIJPHKHsh45EPvungbiUomhKP
Our11SbU5TUqLSf5KvbR3s12YFyxtTIZ8CEH8SWNKMdLFO/4NTja/0dAq725BLUi
EQH2DglfjGDJtI98XamiInG+1Rp7Nk1aDpp5Fyt+3Y5AcB6HxRRtaW4Ai6sDDSJk
CGNXjcLuphKOyWCy64vgaIfbTOSZGi2TOY5o9PzRm8//bNBOXwtwjIN0qZnhIK4m
FKEDBj8zFcZZyb3swUBO59czXESAZEdA46gMxXn3AeANG8uqTa6gy1C9V4Itu720
KAxZUZNtv3O6yIKHwWl53vtXFbwxVeMnEr/DbfhFjMHU/9zpt4Dfe480Ht2sGUrF
WNyzupCuIEYxe2EILFePe4NVnViA8M7znNZyfPi71zUjE4GnX2v5hsf/cGK4Qw1/
EDKlqJB7qS+JLudyNqSc5Gtb+mQ8G2wQ9Y8wWhMtpxNLXe1PygOwTLsdSUpEbFV9
PT9RlRjYqHY/mwWYgDKglYa38XYlHUrAbAEOnGg4J60xrYCTWhhwmSyk9iMbZVmP
decW76r1wLh+BI8/mH1wo5AxzhAeve9RYgzo2Y48+yyqeKyVzdK7X7xgpPX/WDlj
pXrUVy28W2NlW8Wtuvym4NVuB0SxoEXR1GnGGudDoRG3VpYu81O1yb035HCJYxaD
LlFEIdBZD7mabybyT0qDVDxp8W1ha/BaZH2HWYvxron1kT40OKHYOR/tTe0OCsPd
Sl/GqTkg9uDdPt5HenY57V1WyASnq0E64nGVKsvNxx2VOJ+gGX4RXrlekBuiMX9R
rjP8trHpfoXf4WLPyRBW7f9ZkliocZkWxqSJk5mZE5uARp7EQU1QYk4wXpIcehz8
9UBFl9WV169DP2fIXFEm4OuAdm/qL0GBrg40FoBKveGrDYtnZ85ho5x/SdvCJXc0
SQy2yEVrpE3OMmYvnd2Er8kzs0UIcEkseT5u49XX8HTtxKzmB36MT33W2EBvRZoT
bCyqnwndfDt/Ab1S0ofioiR4Gd8I0Ty6sSrdd0v3Cf5axJbpnGO+9z77ADZLQaCj
TBqbWdwK73WE++yDA2LDyagn61KPVQvsT69wTYV2fjephImcjQ1ElP2z8iacvOzx
bvR/uZBClOCd00MM0+TegpYEnxmfuQK+71N8DD3FF1mJS/cGWS7pdmcXPaGPo6Hs
v2zWz0sn78pLWbzmHFDoq26ZPgZu7qRs1ymsU30OZI1P2vFa20LxzvsK8f3G90F6
mhL5WNyFcEED79+9FWxhqqCkCqs2MnntW/Cg4SVQzz7EOoA4g+PeY2ZL6gzBRjt0
Nn5ddsT1utG95MD6Wr4xi1Xvh6/z+5ZNLQraqkBySnkSroTFwy5rk96GXVrevitX
UTsLds2t5L0d00QlHys3vPryur30aIahDi0it3J0D9i8TR8iUFngLN/oK1APqtFB
9kRdnzvS81ZtL691doOgf+1Tqv/hBfAthuzqA6/N9PNdynGkY6ZDJ0reG6y71YJb
63Q4IUsn6WclFDqbmeCRUOSbnWmAX31KDle1CzD6XUi10t75koLpUnY0y4Ud/Wq2
COj8ZkJYEyJm9TtsGfgSiEeZSUEqUU8nvzHrn2Ntx+MlUHP1JTr+/mIRUMHW2mKe
CRzWv5GViQ6XAHycyT1zoeDkoPYGqTFCS2CHeyVx2VBWYFiS33LkHV50OWuxS0Uj
VnUIK15ejsyhCvQ/weBjM8gBdeWRILMz6kmzZ6NblBeW6WonhdjtvIaNgAI/QuYX
GSA5ekSO7VqFwfx43Zm8m1+eDzXuRJgcQDBrLaElYrTUyijWde5wLfUAG886HByB
MN2hohhdThWNUfI1Lp45WsTSaEDLLDpB7hIFvHL1VsHO4iIbltwYjJg6s9Ui/3Td
Px7QtMqsUoBAS+clJ5T0Rl/W10PvgIk5Yr2xbyn8vueB3ExTRtNperwl9/0N3spN
V73gFBOJ6vgkqtKw5Z/QjWhSryY+wpMpwrBhHc5d0+bNwIAwegi/2NGaf9JUNiIC
c2kFOpS0g2DG0RQex2MCB2YFIWGPZC5/Md8M14Yw6Uv1RDcIrhjhrXA4p6I3SPv6
kDpsUm+AezZFT0gjEpTIUV50JdzTakdn8rBAO2hVWjQwyWl0mDPRl+qUekbqyKdb
Cy+jZZ2Q4+AtiKMUIM4TfSjVjT56bA2v2kxhy4iT1tVCDKYH3UQ5UKcPRVk4eWPT
OUVogykgmFfKow30E+ICPZ6wqprjwFrr6F3Bws63wmed6iFnZD2ttpondp4tvTSi
NwFNbR1RS8uNVQ9y3ZgjAzHJbkAI+6MkWrziyPi6y4fMSsqjHsITZbcdebYX4njP
K4qgCIuMSb9Uu+A90BBkXjX4lTvm7FnhVrkjHLaHAyJlddN7E0MdCD3rGkpPN1U/
+UKWY/1SWoVtQCXkMZJioSJIfMdbTyxvbyt2O8/F4pej0CCDwCd8GtHECj5IcBY/
x0MXAYgw3vEBX+kRGuL8o1Jwi1KJ0WToy4P1PXdIiRALfEo7Uvd6uQbClXKnf04C
NpnqC0Pfy9klx8656Keb3d5ktgh9O790j8DmstenDXzMP6ChAyYCzTMnK/qpBALu
3NKswp4eksw/r8tfBqCPAVtrRPuQfHDks+Ymw1R2PP8OIo7+QI9OfXdM5EuAaGL1
xbmGNxR0JReZEuk31HVXrwcCCE7JKlB6+2D1nPnQ1WUwte07BWFgyxsbf1+0t+uq
locPXaq86l9n7Et7Xnp+HW1kXHCiIjdIBAnU+dBvJdG9DrE3MWmUII59yY4aGZkP
JIe1UAqawnxj3WW8iihUtnn93P85Q494S2X3KbuqQgT+ePO15WwzL0TQNxPOvAo5
a4KgJP7tbp1HiE/DPY5n4QbVZIaDfbws8SlZZ4LVQWv71ktNJ/KqLp2AVYW0Zbo6
vCBMZij/vCEYyY0H7QRlVjeydzrbm5rrzwW6XBg0TlmsyNGU0RuAacrEYYMyUG1U
PoxoTADeYz99CHXBVeZ7CHikQbNWxDGntmI6m4QVIZj2JtgPErmo89nQRlg+MTHP
K+qO4OXS03pk1hdW7T1IAjGMgAmgjnoEDFtKlsIShjE4jUeYAJ1CY/liPjdhtlxm
lXxwSjYQS/rzKUOXtOtayVIwpoIwGfMrQTM2fRXJX2lrGkg7ddZpbbcHNMMOPKii
mlbapZyVE0DEcayFVOc5xlt/3daon82L8JEGMfvUIOEpfLfEdGMmTa9Oh/w68IKt
8QuWO5WVuPltrkBeUQ7qB6N6fp6rbelmeCpZFd30JzSs9TgTOClHbll+F6zCRw+z
3fnFc2+gwBWuP+rjXMeEGfmoyLfSRp09kRRSxfUzvJWj1bS9jZQFJvXxNYuXAPw6
ThJW8PCAka5PvN8Ct/yGZhDIZscHDwJnU8nD53uZRxusDKZlsCrQetKJlY7TTCN1
zAtK4rfmxNFqjY4C3TzzttMnEdzjaAT/ePG4H+Fz3GUWbtiwm6hvRYtMjkifYvq3
jJY8fbTlXyAacZ8MRGElWJyWHicuWjjqhEHLkvShuFRu6U+Ku9RZgSuVQLBHkzFJ
/cncpGL4EI34Y8GWYN7De02x8K6IfG7NXAEqCD8g1K5O7lC8SX5F0TPrITAtnimZ
FsvFlhdg/IWmXk2sgST4lGX0g0GFae0mt3UEBK/Eq7JVk2m7iIadtVSzTGuPb+rp
He6PI3WInQGclq4jcL90lGe8GEdrCJ6leh1VEa57WEJakedpDV6Zs371lF2Lixev
7DjXqQbaLEVUpJvsCHmRY8kEjyNqt+jma2ufaHMdeZP1b3NIctZI/oyP+zBpG1Pd
tkyL8r8TSn/YhuxqErf4xM/w/AAIdJEY2rxVe8gkxRh2mLeq8e4SMA6KAOnKJGX5
gpYoQm3AJsCT9k+qZvRmiwP8QhLUPKYxGnzcI5Tvea4Wutsam8/1cDPOxZqr+112
hOWUB+3mxtSz5iT/Pyg+8J73oOCZOW9Mtp+HRAdZqKyHKlzbKxcL2bAJkrtfg9XG
y2lw3XZ+B9NggHyEKCSbaoXJcbo17dh+Fwkaupdxf74NHhVZ6B8E0RbYigSObj9k
3IEENhec8HLMimkPA1e+bmdnjM07JbV27rpFV/zaaheavAMFa7+ud3bl8iRZ5mNt
Ce0BrN3em9k6XkN47SAk7NjQBp2suq8kVEeZftmlCB4I8b5bgLLJ+TURzsbmVlz+
2ZLNjmqHeE2NqXkerWTlUSoZPgZ4rAXZl4/n78GqGO95/v5zgwKwe6gFHfr2LuPv
1wke+kj/NmnEyDMTTm+J398L882cRRqS8IgxNcRHP2bHL2r3ShUulkANdb79n8GH
XD/rOVkf/7qMKoAd1PnhYkskoz1dM4OpTYfE1/mUObyOrHKrEeb7jVK4O+fB9W4i
BQwwo2sMeChQky45aSghvVQTZCsiBUFyGox554rw3o6pVhrZ6ThsGSN0ZpBPQAED
w1ivYiu94ilwudB0oTXbixR9PlJup2FwWhRqvPMo7QU8z/gAOYpcBNY7hmJg07Eo
FqRsRjqgpKsQcMwogEMeLYmsf3rpHf5ilNLpj8vgJXqhJiuluXlEHL2cUQoZYpIq
1OpIxKFtfWOGeiPsS22RHNy2KtPX9GZpC2BEsjY4xjZAKpzlLsGA1itLUHfvLH6Q
RcVGN70M+EluSAl6yngRTGIklvZtUzP4P6TM5PmNYRHDSTszUHbbvBEW7qpTsHUD
r62z+R3K3IVdnOYm1A36p8yfrFrzdAYAX2sls88QXpmWEQVLOGWYXG2mZ9RlgWQU
gZ1jc01bRSDxvS2hKX0zWgv421rxYeIPWVhrmUwMbqp+hXMMA0QDnzt0uetwAJj5
EdJKm09QaMJiyEigmEcYgEsEZUOM2pSo98f6gPlMvau9iDLEFnBcmRHpDX91P2nD
ppmm1XNv9n64nJCCQ/D5BS9KNLKRiPIw9/KjJTc5lDXnyNc1i6q7mLSlvSdupg9U
dRdWLC2Q7Rq/oaOz6JMoW5XjPs/778Yghc2sTlwV1M2XP4+UXBD5BUFll5LHPucb
w5OLW46Sm5Kviggf5EAikCJ8mO3TSJy0uK5TPpzpnyioHo14LANxePfKtF/gfdPJ
otBZLJ1/H/hac4OSe7USELQ2TIcwCbzeraykFoCVkfiqi4pYQKI8JWhO6eLyBZX6
PrziAgFSbJOJg633NardCcq3w1Zple+s5CC8Vsmydil3LQ7uK4FbbTBVJgweKv6u
Sq0bhkWqzWIs+Vsnw0sRZKak2CIcuae00mgL6uSECBhx+iOPgV2TLF5zG+k2p6/P
GDY1gRSmrE9ySiLZGry94ETrAgECDhXcnL/i9i0o40/Cj5KGgDaRfF6lImITXIe8
760N+67KXEinGyC10xsMXvzuItxMd69KHT/hDOqIRkSuFegMRphAdv4EoKslqWx5
LlCE9mNH6n/jvS5/umLjHLFFUzkXFdrXWoE9Dn95K4fE4xEcFk1w6U4cpykiVBME
9dC+GpPK5OYE/G1NIOdKsNGfcD7qyoh1hERbAjLbDz8AJ2CdGr0EczpnrXlqWLWD
vRMznuMheUnPIxklizmGppAWK2s4m1ipgydM6JgAKyRVU6agNxg4HY6or8OpVWiV
DnncUEtbUbe7amhCDzQEdygdy1y2/18balFAH7g38w4rTx/vr8dPzIslG5bBRadA
ogO+Sks6HBBwtLWTGawaZO+wYaow1cThEwEnupd0SxnEKNlnQEzI+8waj2mscKyt
unNjOmXniFMh7ZZoC12EyEQmJxHOiDA/g0CPtrN6V6E/Nd7xiGrrydeHUJfjqkMk
enOpaFiCgGqpEKzXU9bZcXcsNd0pu/UET1/ROeVS0GvcJUbtHnA9A0yshXgI1q+V
urHTSRq5eXETxbkPuclmhY6hQpEwf0HmqdoQbADVzMUUJSd8mTG1Pm89wh5QDSnh
Oz4hiiejE5QUhhVxZOJjxTpYSApISNj2f2k1tdx3cZ8Hh76+kmTxI/g2NhUqKVHu
FhCsRJ8X2ntZCt28TAX40fte0M5m+AF2bYdq5To1V3ZEx9043o4tDvA6xbnDZrMR
wPWLDfWDUAcyWY44D2/E3LY1yiUS8VtVL40hOOSQ/i9Axp9lm7x2b3yBNlk8cfVm
leNRaN7RnwBgW+nekG2vV6tM47b886fkGpl/tVIxSOBMbjFfgxD+FK3ryPlhdlBL
tSRuReDuqvGJQ3Iv1/GqryRCiQIfPlcsfKmKxmZPX6IRdqy4ZcoJkMBfmi0ZJHpO
rpyMGp0Rp8Rgzu5r/0xbTDw8w2+RTe4urU4ntOs4RiN7sRKOrEsvf6KcZF/LAD88
kDf6f+fasezsrJilQuwH5aZYpeaKGsuWuwIJzQUAT/khvBy6fkFTVSeo1w6s/O18
pHoX8LEx3Pz8ZR9DI7Qot4Mbt3WQmK1aiuellx3GW1Dnkmob1UHZQVW35ZPS8GlG
V7y/0BBZwa/anc0DMOd12VeCgOOyXgVrsnTGSsM4XRENSvTsXOhG31N87h7klGOi
vvS9XdPYu4dIFFq08D7FuAv3utEXw7Fw2YCo/7QQ6uA72jc7LSoEdk+p5Zs73+H7
XKNHijSDMGRSuc1VgStl7lDUYzSrBi6Ss34uF9GwKvI4hjFOs5HjIgmVVJcu6lkc
sanTs/sIX9b8VuN3xPE8cgpwacQqGW8lUUrp3+1oPkptnqWDviiKofKXYQAMNhVF
9JrxPZKqAhQoQgm83cKTln5uxK5u1FrUFDebf8csqw2z++yhnGvUuJ3/6XJc+9rP
wTcOFOmYQCfASlrXMWFg0bEeVuZUswMIj6KIhOx7YgifAyFfQaK+v/HnqJl5Cwj0
KV6ydaxo1zUpL0LSpHns6WkCvJ/bkf/74MIW9zfj06Sq8rCFcpOFHiPiJp9xQol3
bKsyIxRllFI207MJYR82tnxK/Gh4xdE+mDUWQ1/PTgB34O4aM9n+2qIy0n6sVy50
Wgz57EGDpldher4GMHa3befQa+fq9YzfRJ9cyA9iP2hPnBQ/h0ISAbsuzVyak9DY
PSzBU0331OzHr39YxUT9csAQze/g2fPEnzCWoA8JWm/c5o+nVIAcqqUjKIkYVgFa
65emAgwJpdXtl1ArfPkQyuSb9oFE3IJ//9yESZ02oIgEKYeydwkxdT/VvSwmBLnI
dyH0dprQle2yjehikElmClX+zuXuf+VTMnikjJg0Bhq6wx7UesXKSf8Fwigi/vxF
vfXfWJ4BDd0D0jA94Q6UIUA/fbnuCeMrOuIdIm9K7LcBR8DKB+vNcMrKybCBQrQ8
ZskNgwh/xszHfJVWGjnZRn8hKsWX+jMJ2OInXOOFwlos4iab4JkoC58Up18E1Ml3
bFWwkFcmXz3+xD+vBb2Uh4xswsYwnt62xidWItPXtMe9r+1Hy91VdRz5e5dhsANE
MOYuGXz47Iplg8eXeLw9+4HiMGulIepHFfOKLVDpcdghf1t0vmb/JeHEg+7ZnaTk
DUCq85cEk1qIPMfQGN7LDj9Q+nkLybzoSOxpU9sNy9bGrlf2EQZILx3A1fqmPake
j7nMvUY2qblzpK2fkwzdDqs7ioI0MUlDkoOnuWuIWWtfPHWWWwyBWIDGRmsCxki1
t9S66442WEYUPo9BLjC3s5eGcdJdGtGg5bvbGJNtzKYP3fcKZtt+hgukkBg3Z5Zh
qC6g1MEPdAihThWLEXuwpYOUey+HiaMNkQIZM0Kv9/Vt981bWbN6n4lXjoIl2n6R
5zTBoaju5DfdIjkm1oki2rr8aGIoIjYHluj+rPFwz2jumdYt75aX6Ok9q+TelZXB
UbCt4h3TMIiWRxHAnANhpWsbtxv6AjTDqFoa57PA8OQifZKD1exg+zT4FpJxkFjL
joNQCwvbgBccBQSDnqsmVBwKAbM6dhhk6/H3VkFqbpU4DTNCGBjJeqjXFGEaEaLm
uy+xUugJDi9gDn0zBN/JJCGjnobe04Ht/aeEa0B4tquwXowmwnzEiP4uuYCWjWTn
EVvFc7+/KKtTVID9COQvdUpxrzdehmA72Ea55LGVXm/tncGYRms2N1xQBq477+U0
3uyMUrVPlVSeEqOf4LAADLIlgrrAgDmBPw7XTaWfJMnBTIXGcqQ2EmWI5Zh4+CV9
4kcJxm0Aiy6ujkz14UFnw85IUX1RjyXUO50pB/8xeG+tp9wzpsF8qwqzBEjSWrdu
hgDsghGVWw6Ch36dk5ytMuk8hhmNToIYmi0ewDpD3vrU14i8+mlRifoRXa//PFFR
KFqaSm5rB9Y/mtb0EmfbM9CcWB5p4zD1VgDBmY6VkuKBKQfKujsXQnT22g6DdXVw
31r9l48R7nHksHDBPUOI4ScWtp5HU5SvnvFeCclyBOIxcx9S7ULvtBmY8Ria6/8U
yOhFVH9foYRP4RO5M5Ui3EMn7er5Z3yt8S3roy7bKNix3mxjwySv6dGYxdKD7fON
0eF2rk5KSKy8jyV44WLpKT4V0cQEdHocacEXSYTq6KhOYJe1EoVacW/VB3rCrcgc
DD0B1CkET8Z2MrCk2tdUXc/xQBO3ozwG6Qo+Z3Sj/8v1P8I0pdli67TerS3TAbkK
uGNzp2hLpP7miotKG3hbaaGDFuc1KmUQk7jWvJ7lrhNFH8VqDoFswtpHkyoWHI8V
iSrbrYB6c/VkwEf6T36F46VVjnooxzdJB1XCeYrB2TJnYhNIvOpSKdCIAhHzMyfO
cq7w/EGw0Owj+7DNqzmTnjJUjBkvUZAnZXXNnEWHQKMG7eANaa1gzSKiZ3yyBIr7
EZVR06ph3S7RduKpRZUS5xFJsofp/GfrolPzduaNAnruN3W4HpakpCno6zPRMG6u
Z7rHxAam5b1qojfsqTnR50HbwLymd1BM9loh8JefLkoHWoSD7fjBEtVY25HrILQX
qPIqZZiGqIUKfLBwJMyWDFP4DCaqhvhQKiDaN+wNev/Uvy+w06bS4/W4pADRaM0h
j7tjHD40ZM3v4Z20zTptgFXPxvRPzLefjLxYXz09O5oQBV42XPGPyIStSBOAG+eH
8uJL5G3+bnGWcmjMbwY+T4jQBu2G8CCLuOopiuhaQBBNAptQYVyWP0SSM94gPYUO
Cxn3a8lCqLxLmKncCq8OExCfo25i93dfj90ctjMiQPEuQl2KXzmemAc/b6q0uHjk
NGBJ8G+1DNkxKNu/UdicZTirQOmxlm553TE80CneMO+ghRTTbVFBm5xOn9mEzlJe
Lc2+CkWWtxf7UbLJG4oaEAYYH59X0sT50XzOLa43LGD69mFpEv0Egy3Sr6Hu33Kj
lvbxDGwamaaiqZWmZIkL/r2OMJGjs47gmsT4UKdB2ob9r6+7YTk+4y9gEMxCtDUo
y7uU8yHYM1khTi9llpdpyeO+I0tYBFyIm+pa4VrGnmGE5O92MRxb5b2etka2xWjg
aw7sFs5ON49KjFTYUl40nTPRl1oDlvliGG3oQ/bH5feTf5qpHAg87s0ZhTxuCwAx
C/mHcWL+t4916T8Qebriio+oLBVXNrqUrL4tqElmvkopkUEfetOyEWvIdgGKwpEk
OHaj8FZDF60J4W5EpH3WwywcfVOIh2jHLR30XMcXTR2M7N6YAAZ+zi622zq6h+Xn
K+eZM5vBUrdqHwh3+k2ELVpkh3KvqlN3IBDED7wAMoUkX/58zBqyiyK+fGo7+/yy
mQPExurdZMbR08ryXEp+FtsmP+oRN8Xx3tqnmEYIbNY8kREC1rNizY8BdWOUwZ8I
yQ77AGCMjmPKZeYz2ycfgUHJ6+uM3g2hYwSjsgyHvnhutZxtRmZZ6cLRUraXJYw0
g0kHnTTsaPub465j6sKjH7LkIHNo699z6WaO3fYPt8y2U6BmTecu0oblczLvVW0d
E12SJ0YbH86ZbqbGhXMyvFYd3qcgdxDqAoGftWP7ZO8NeVeRqBBpRcNoTSV6LyP2
wWhjU3cyWmRTUdT7sr3kEtyi79oSc2OHjV0M2g2AkdoZpK0fQdQ0iJ+YfByS4lpo
BD36+/3mgbgzADBQdVuJgwedf7wdB1HnIXIJ9IHaVC533CepkKnyIdUeA++EEC1K
KscDFnN+oKSW5P4o4IqUrPf6aANfuVicmj2sRl34em23lYLt203DudkUyn78q7jh
epL1pdq6hMdKPISCzLuYM/DoaQVNTlW7peUdke0dFPUu3SsSKFyeYRvZp4nHnqQK
klYIag8YSUUnUYeKYmqER6sHUGogzkJ5GV5NzXswys84nUkoFi9Dj2sli8Pfq0iy
enRs5pEzFczYr2U0eVAj60VyR6lPkEfnzI1JLiMbU/g1XvMp3sK90to3S51bqsPG
0/0jGaQazDVuSBD5PwaqoI4hFBbrSjRUcjLkDvfvs5qJNXvaskP9H/j7OgpS0CPu
OFBgh06DBIEZpMqupS1H/t4PNyy+uFMafCyVepuf/HUx78dXjwK+ohf2HAyNy9d0
T8fGGacP+++dnt/CdPwDeionCantiGaYKvgedhUJcUayG2n2mhLlZOSGD8r8Yjw2
fOEmdEDq2uOudnyevJy8rrR4+R9eogZdkn0uepS58i5BGiMY1Z38okLgB5Yos/U0
fpkvd6RU36TxDiQm1zY94SunCKg4WhkUy057WW8TtzlGb/rfUBWTDqIpND8LFigQ
LBRo8Z3lWhwDm0G6n9hv9ZPXUmb+IbVbS1EiQ8ULfn+0VSTBf3LyCdUlbBNLqOHX
NZcPlUiqQWaZVUfP9n9wYRYcT040PXpNppGmTjFszW8=
`protect END_PROTECTED
