`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HRev2nAOFaDzQEuE/IOn1qvqQyiXb3YDD1On/mrDyN41VE5IqvqkZAx4Ti/w0+89
/wexWEq28cNtlYR8hW92vU5mnaS98G0co47CsMR74iFaOF3MjHhDvz7VaZO+pSU/
TBCgt1FdJOW56kYl3MTghFSLKjJzIUwCJAP7UPauWr9SYKJdTO3e0of6c3Gp+ZDa
GykSWfhJRNa+Xv0qTxDmoEQ/Kfz+XjtSFfgOpFerdazY5ebqcdn6R5qYWfG+UTo8
m3XTD42CeDVczgMACUHctjxUIcd84pEtT+36CPDCSlq84x42pnqP4f8feENQR+ZP
5lAvM7v9vW64QJw9U6F9tcO9Oetiubjk+q4xGMtId27JO9OdXT+hYFJsFr2TLhLK
cd1XMATP1ZbfFVDu6BdRTODq20IbyiDglnybGamFN/M75Ss9+wLRKHs7tmsAI1DT
B+5RmtoOiHuLMb0ewOTFqUTVXllcQ7km15C54+8f1gp9RS1fpOPjrTKHFQrr7Uuv
HIVtfwhplpNPbbiDHmphJurrXNt6sutWul+MDSxmyhRts8PmL0HQkavEivwY1DuO
PohKKujqWUgaYQ+9UMyT7iCAK4/ejtNGVue0quum2lG2+3wh2bN9ViAKhhgdKkWm
W/LOPTuEJHuWnH+h/SdHT0lOgY+hMxYroUb8D/xIgpK/jVTPm9gQWRhGJr31D9Lp
0L1JHTxZ+EwYsWbJ4aWEin5mY7MzgPYH2WXqynhlJNR7O5e6IRlm1B5JFuKddYgi
KpJU4UnfuCg6KTAFyUwtnSY9JKl3fyI3ZSNbxTZ1BCAwdtisga9SA70vNkiqU0H/
p6y+fX2MWz7HJRVHeFuIMp+DHKcynrAMEV2y01yv1qQFXHBdmVOJTI6ag9mI52pW
M3M7MJFnGhgxSigk7Pmsa2PoByEYXQDbKo0bRvkeuf7bastIWPwMZANXbjKhwNI0
Uc0i1lKV+lFn1Fh33aOMFZfupC2S2eSDIykRUecmGbPzNZNe4eGS4cu/KSUBuzrQ
ZQA5I7gLybMMB9FGx2oIBCAJyd3eU3S4EH/v9/GspMp9PgWPfvf+yKIZrDHs7Uq8
s2WrBvy0DF8pohj6nOtRfBzRDKzpdSx+V06msW9I0//e+f+GyKCVfjemKqnyqQsG
6KLXb+xJQsLYgblpYBPlIF6oBaU7iWwh8cdiL0uibWu2HikTpVvieJsYdlL7hdyH
aDvW9yPH/FcuY0QMupddspgmFgGdvH+O7vpkKjifsd9HdgMH1/jZNeEiM0ZvUcKT
Sk/h3Z7/A8jDfKWxeOUFNYvu3PKWgX/QrMtiZXbA84HxAK+/RG5e2q88ERfu1dqC
K2ynVOd0OO8e3Xh3Ml9nI32I5nhKKxOiHhnLfT3jna0qMj4D/VeKIRK+D7Aw0gFo
C0WBPzvzX/oYVYYUYFt8QVS2ZrKsuzSJDqir7lrrhIrfLFpUPIxPLNKprOyYt8xQ
+bB9vUESo++wUKsf/IkcG9gKVg6poMfxa6rM6FShr8KUhY1E/jaB4PcfBfiayaXf
rAr8/23X121cFg5pRGL9ee/jzJxo85r/uRGg5d5ICO8KM6fmVtl0KIPQqT4UPmyc
GP2AtPIuDKa8BfFt517XEtA89cpna4UdIZiLDl8C+V/zdwNBm86nH1HgVesJGFVq
LKt+asqkomWK5EDXJPw48IOdst9Ht8lFC1nSpbocdtmw2ZrLSNSgbb/0dPvV/AmT
6/I7VpXR3BT/a7nP10yzgVBR6MqnAMGUClw33Sly/DM2ayax1s0JQADePuq43kH/
+kI4XRvwf5FrAiJ+O5oSwLqykIz3vdjZ8/F6nq2zyaeqz2GTV50s8jwSpB+H64tG
XUZbMNDGS/pPDq2oRokFX6yAzc3Qb/EYXSyuueOdTmQeojOOkBwjTFIuoz3cGYyl
8qVPl8rCEs5bb5HM/1LvbR7yGmnNz/sC13Hq3X6Yztf/kHwBl8YaG53lrPhLcpCm
AHtO24mnk88ZzqGZDNQfDbR/vNIHhN7OoyJD2dNxzZGdd3R2AYEhCdkUEbJIXvva
O1vRFacP2YWIwWIFPZuLPEB5x2Le/xrj7CjlhGfTWsxFKWBbZbIjHQyJQDQLzBsn
MytyfzfkIrlhzQ/fRPr6zX0Aa8akFvUMhSe7Ji0vjG2likxA6yI7cx/BN+crOOuH
D96fUJNdVPZXwmrAR5aDzx9rqeHKZfSv/UxD5HIN191fttyMzHLvNXwUQWxQXfvu
EQAHsx3KhO53W5jMixWKhtVWdcwQjrEGquUf2lj5rqLW+CA9+bsDhauzDwHCNqVH
w+EUMg7534p3RAChuvGLD0mkVLLamcvwG/8dc7Uepc69v5ANCsX6GJvOOUuc7RuQ
BoWUxRnwbdvxOcL9XLqX/2jmF0+AtO/Y4Pe1GGFjlybFP35NjA+dNG9vk5YJZksw
EVm7C2xiU6qJlq5q+HYKJnX+bgi44E0op9rDvGYx316G+8mju1tL3xf50hU0UDIK
gPb9dN4p1fPstWZxy39ViBmGvb4dqd7drR2hdnb4p3Dgk5fsWhX33mex6V3MDgx3
pK67Eva8GMqFIhd3zSaDUZZCprs99MG7NqdQya2KCG0OFJ3K/CKTi+JYE9Sy5evv
tQ5UeTQQ0ZSkpp71HUaDpro1Qmgm7F9p6djAq9KK6HoP2CPx/1XXqSnvXfZjvUQ4
GBKN8spBiL90Qibnd8kySuz5CvkRto69/oTunH6OqwD2D+nz25Aseruaoqqz6sBR
G2ex9YHeITWJnCJ/+wT62504nXhjiTSgXjsDY+TAxFrIgnBLMGWBKlbvU3dgt8A/
cSjnBFwDxdIQagoPQjiXgRj7OtEaYsj81BppzMK6EMVfbZql2WM+/+5i6p3w3d+L
5x0M2PUzieu44EQaaB+aRmPz8EaB678S6er+R5mEHDsUdsuCagbe5uqxOfmeyhU0
544cL+BcpO71BT6nkGamTY7zD1k2oJLmySlUfDE1kadxGvOgngqixFlnqZ9ZhkPr
viA3f1a9hmdiJNnk4/kLhbbkm4d3aiUfukFRTdCkl6jX/i5DsS9k7rEkRT2CYdaU
JRNYt7vBpR2kYYw43TOZHy/+oCTVcWHiJxInjzOrIdLfhWVCcM2C3KWhQNb1JpwX
nQ57nhKOO2LwXOSJIBGfNTnGfj5UipgTqBFfIrVg7Qp7Lk0BVUEWzkLf7dam4yRO
MIa+FeOZLB1dUb9DYFXOP/MBhFfnYURx4jgfmcn9mnlHY0I9GV23w5bim1I9m4WL
dIs/SxI7WHMcPv22BR7O7QUUyLhAgrr0OA/XOFfyi87RCEl6th9xxDRe0LJmFdh6
68ntkKdc5DcB4yoR4u79bagpPI95yN6Sz3a7FBKmirBHAgBXZW7lOijMSl3TQKVy
FdG1kpiaCyxRsysvg3JO0p8/MrdF5rqbyzzsijCrCYuUSowqJDHnUcL4mM79dFts
bNY0YtT7iqxKfXtg82BI/maV0yQ+pJEDMk/FxCcatioAOhpiB56LkHCFGUr0/S1B
N2zcuoFhEXn5vGefFGqjHNvqqZ3qeWE0s5yU6BOI7yPHPhtSDOIRdAOGmwqoD8cq
/Y4YZK/GEJfuFwdeWM9juGyQ4D6kQhGq715fMfV911JIIjy/Z4Lu0ijV1sjxHMZY
J7TAYA9z5ajtkOvLzM6sOIm/ZFYCbaGB9uogKlnDkxxTPbToC3Mc3gUcDmymL23q
jg/DEA0ReH8K0kuWJe9EGVL7nBH0zzVhloljBkJRajWpwsrEz1DNT5TnIkohxu5e
zUbY2K+nGP+Q2EB1S+V2e5OYLjgPQ3kLTHVQd29DEI/O+elj8Dzc1qvlZpVua5lC
5QpPy5xnDLEPsT/p67CIkQYdTb8YLAU0vc6+7YJhx1YF75zS4yBOOI+5iT96c3CL
P3fRRIPkUIMFXhAEiDSOJTcWeUvggxDWo9qYHlABuPk0NAY5zTGd0KAoO/UqyMbI
XZdoUq6hb/ccxrgUYk+msB5myFBldbzZ8cSj7G/uz9g9ftmbxIki1Df1yYppo9tM
WP5KHZl7rGk5KSRYW8bf8rWEPzhiNZM/qGYVk2007ytgD9WS5FgQFW5JAaaNHPwx
bUuSM5fwZRwbksnnqL5rl76Ye7HDKbL1vKpLWOCqzbezBn7NIWW8wAC3zEPtPAZV
hIcZZXbZNVv2HKAWCoAnUWB2Yi9Ds26YzlIsVqNjcTShXb2GkNFkUHJ4hT2hautc
PctIp5GqNn8rhCuNKksx9vcNcHQTakLNJ8fEsP/6WPEdXeg8hgkTuPZYO0mk0jgq
Qs4l0JWR3SwQe3XZjJM6CyHkajgsGVrM5XZS01JWwcrbzmvNV/4Ab9UViG6e8/7C
oWdJhwgmeUxFUtJ/r9cqL5jKhX8bw5Si+CDU9O8jR5qGEbwGtA1jhB4VQmouB4NX
kkNWovO5TrArLFJvUAuVKuB3xbupf3I0rNm6OWyYKFnKRoUsstdesYDSl73P44U8
TJjD/u+XPjEMSQdS6GH+y1zmIvTw/50jtr6O75qFLVy9QnQkqFXO+z5rUlQ56XJJ
n5/SHOkpi7IxmcMAMEwkTz8j7OgMtODGQ79KSu9cHuKCqsK/UsYAdPPpTeB+Nqnu
asaccdJ+2ArPjkdKm0WclY/Q5gDVEcc5ezx+fsw+tZB94vRJFUyupXdNoarmDrgX
qqJCKQKEC5zDn6iQQgfW8PW7aXe8elMHdaOc6VRwZPLsayu5kXjj9gD6QCMMGu10
L620IePHuoha5p/4L1VgbaioLVGymBCN0NYE1lxgqdYFzJl8PwGADnIdJ4cymLpm
ehCI8gMDUYq0sYO2YJ7EwtquRP8s9qtuXUhUFiPLCjS/bGy1Jzwkm+UZRsVuh4hq
PqoJJnPMG6TSkKNmrveikKynNLCqeko/SG+JWqzsQ1ixFIbPhNirwiuNFhn/fKDR
os7Vi9iSeO7vJecuI6XSQRkhJnLO1/cqGmDNIv+8+Aha63CSG2KjcOCtr8GGo2+A
pSiJZlcDyU87FsmRbtMCyFYK2mfZ6zUt1ycxJqePU6HocddWjd+VrqLbdPl+HK9t
3okh8Tty77C8E+otIOlXup9Ss6bXOXSNNqlWBObc6+X7RTiKYICYH393z/xjSosy
241uMVAIXqTIc2tdfvVm9bd2Ws61cfZnXbqqrE49NQd+2OD2V9DtxslosWGAvOsi
MyW0ZqweUm889+esAZaVk2/0vQvzxa0CcVVKoD9LZPXq2PeqqVw54fMjBDLAxcP/
Zg1RsWQTtZNmNFg1Ri39yMnhpZEuC37XsKrOo9vQTqrxD7PYKnAdngzFR4dazcJF
Rbm1Efz4qESE1OabK1pWtHmaEdXSe6lhqFCafxJAEJTHSl74o42Ryg/kncYyAjPP
neyYCU7+KdXK4rkphjnGLrzL69OMpKIy7yE1riLopEZBTTXLTNV36LplF/pQmVhC
499+8awggQBTAHyzivAgDxh3Ik/iplxUIvzrGM4+x69sSokQY4XxUerpRnl5akjT
Nq1EEL6sQ3CqcxGTEFxAPWuLbgaC8qK9MECPwWOOcsscR9l3bdT+Xzw8OSvoj7Mg
+wJZ2THGCDSPS2mUaNU9XgTJEmuMQObHWZ1817Jj3lgcC2T0T+0D1XaRS/tpQMOr
5OVSnnk5tdRKWa2WugqAEoXJFTd+zyUUWhWXI3X2ca3KLsA3vYv+Fwq75i/e1czl
6zmgK1j0udsX3vq9CNSShkoBI+kSwS3Q3ddWfxpyMSzugb3dZc/UoqB2JSVP/kgu
CoLsNWxIO1vOP92TN+0s2YrgSiyDHRoxrN/MjqZf9Y+KnEeVi6/G71QeeEEuAeod
Ndxr+53Nyqtharf+0+Gw+mP9ZLePVptCxEZG1XUxP3xc/dVTzIFmVx47+Rfj8p/d
0W+JvKZwoe5+tGZSWwf6WMprXLAqwKYYacJIAkFmtu+fUrSSb7b7sz6nw4WT5jh4
SCxhApVZ2vTRnhbB5ZiKMZbSD96wcSR0prUviGWo0w7AMOauibOStrYl3Mur6+nJ
RAlWwAaACwKSN/yuKqgFrUbv/ikLS/P8caJH5vP/FgwAsWLwLscX7WlDjhRXz8q2
isLE/DUY3XEJ6MPcG4tKI7Xnbd5+NEhClIG8nv6dqpJQKRHzMByP75zelyjmMxV7
CF6anjByUV7To0/8aTfLvCKcS3d6kkSSwaJ4DGsCXPzpgCm6dhEqrGuuGXfPaB+p
HrYE0a4C6nSQQjBC6JGtbvVpXDHmbjV27bThMFo6J6IpEj7lcpbAq4aiF1evsHsO
WsKoKsxwS13bcAjbQhYgqY1dLhIdyZYV1VaG+2bNA7eEinwILM+NfTKej9uMOzbN
DlcpWnQJyirSEenYlkW84X7G3ovkC/IBY8g9Ufjfz7sQwKE6lubsWWsaTLmoJ65s
o+FZd/tPI0cAuTjtMyi2poR/k0VsIabZ33Ibg9yXGRKKkPeLt8ljn0yVufYMwX/i
TojkZ1BTu8h9E1ywE3R36vBUvHz+65jTLkk5BzkMu2ALLHsa/9tZaxPDlhnU54d+
kQCf7SpM803jRGgJkROEogEQh1njlSE0DEk47p6vyF7qgqOPSTpy8gbHFWz+tHR6
ePqESI98GEqqG7UG3rQJsnnb+DlZoUxFcyuZf7UtO3sOovzoXyTfYaKdnbQUcUWZ
9R4Y90VwPK8XAsUYl8yYOqeZ9SE6l+XkFVkzP9821CTiqBObdUCCLgOIGkG2i8RU
8R98S+53Mi9zBWfCVpH0n6DBqoPSeFovnW3DqOaEcJj/t0j36eft+NqghSVfFhI7
Znev6FeECd2YdsmDfuNADlJ8uHmr15QFrSpgkcftxi42klZSELrXTAhpxkeS5mHb
WZwProRd5BOKZiuE1N2w1OJRTRx71uaZFkPAfNv3gFhRrRs5vfJ/WWhO1FYUXNWq
HZbtp9YGwFvYrLuzf7Cdt/Fuh4gNrp1fByF4q9gsfTzYQqiegqiyRDtfNyv3uXqY
1Z7F4my2KNkMlp19vS4rx7MzPLfIAcsNvFdmmbfYmxe8rLbEWWLYsRVg3vVWctYt
J28izBLbbe9Yw5bwYuPDh7YrnGuIEjxl2wNJu1KT2yONgJqHWESOGZT1O2VXbiDT
TeQyibT3vXzmE1PdwQ2AYqtzYEoUqb8kMomIDJ1JAhRh7l9qlsK2nPl0Nv6zWNqY
p7cuEXaQ3VoVtwfLU9qVIqorfIlB2CFi6LeapH4fnUXtSjtRIx+/L5bB8hhFmas0
DyqM4ZXwKCkts9MWAVjpcxMivOaUr1E87TFIe4TjY/094PKiZLJ7WCFkp7WMmf58
t+BbAvmQeyCsDN0eLDTG2IpjqSOn+rq7uLeMb0eXeKFBrAhX7Iqc9+5J7Jw5xr6K
igjNjkwvfTQ6TRAzVRol8j17yLZJl/AUF4WJmNcwcaPaklq3/5udJNkiqcRsXY2x
1LqI1oM7iX3/NGGa3YWNCWGJWWArYMWylFgAYEqfM8WILhzRmzw3mdkAb0mDtb0Z
Rui91ZAoqYJV8V0IjYDw+w7mpCgCzvbh7m83bq3WmdDtTriZMRkZe07+U3oEBum/
VYzZBgoTXD0lv+ZTdRcknZbamJfK7jlU7ui45o0bx2YA9NSVLbg4P1m8MJndAPXT
3GJZI7d1aqfD2qq+BshUFQ==
`protect END_PROTECTED
