`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6M3SBwjDzlJ8Jqynng5e+/zKZcDWS5D8fQGqIfyXC7aI0Xq2CIbD8Vf+UmPRNys4
RLxl5RPU8oGPrl+QnG1ELW+t/4iBwRV9O+5jwyEpy9Z5KsvAUSkBXKsHJ2JyiFNi
4pOfWK6Ll010KAC2/TECJK16/qa6j1Fhm1FEvQxxM96S7qXxpMkhfIg803jhuacR
NsJ88BCACStdOT1mpxflHYLQXTOmY6XbDhPRJjVx1ETb7lixF7D8+321ho39huyX
nAW7eeA1D8PJfEk1Bc2k3lUYU/7P35Oa+blBpXaIOBjeWbiMJqjf9HkZARz9RUCO
+R+/wiRpGI1V/KyNM3ZsChbUk8uZh+qD/0mJQEI2DKFzF1s8zzv3QBAliOtUqmZf
U2B6wIOiqRnxl4uNPANRCol0gtCAaLjWsOI+Kt5jmJaF1D3sfxiKzni8HHHG6YvV
TgTuAG+u+c7hVp2F0jL40O0ZwxjiSh4ljZdQKZbXkwcdHIo3oegtEG6nerDreXtH
zA8ciJpSU7p/zEX5VLumHCb+82YduAWocieAsx/uXBFzmYmqKxp9STODVlqcX830
oShJcUMVANQ/Gl2GPFkAwA==
`protect END_PROTECTED
