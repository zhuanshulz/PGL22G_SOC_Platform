`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l3B1Wl1IlpeJTVNHB+hGeRuoh8rII9wkUMH5hzvDjru51Gnf4MubFSiKUii4KJSa
SxZXuefI75zg4QypMLFc6war/gwOP4/PELpB4TVTKjkYEPeF/VQo4SUV/b6HoLGf
KeEbTzrV7SSu8BM8xKF29GKqBZKlS1fuCYXKwgNBYxYYshmBdeFvoSxxzBtl13KS
NpwKYYHwGCXYoZm/knGK1DquyDAoEXPBphn61NbHZgS3/cJoan/3iWJHS2UMEVhi
UfmQwROQC8CAi70W+cLLPmaoWh5IimjIMzO1coastdgILoCcMirE8yofFX5VbZln
nAr2ri5wgJ63kDb0pE2Faszfqm0C+kmn06F4iZ0YstbWlBzzJn1hHgyoaw+yasrR
J+6BC5MnYpAC3dHZBOVAk9QKm1d2rrU+JjxnWghon/+9zdA4LVX+JENiPjY/lY9F
E3sW61jWp/R2KIfbFoKQNT+dG0b1VTu6EyUgphe5wXQTDG9Sg5GFysIXhU0lRJVP
BJDgw52jxNg7jhAix/e2VYMy/vljyYCOSM1c3MSP3RseBwVmi9juP38CPkhDocEA
2aq6+gfJXEtI3Y1cFUkIasRB0otd/6rvIfU9LPVLwxGKrkzXjJktHKMGk8JmA/GG
EanX6ltLyOsCDHmIpQuTAiCAm0I2kXV3cBRmowvl8vxkyshSHISd48O7sbDAMyUo
kIX+agcz/g5ZWlnwmTDKZ7knS4qeyBkWtFZXrK/GlYNE5kB7y4b0dPjZ4bXQ0Npq
21gbTs2+oJKwAGTQPCrO8fIUbSiuPDd5HqJYI9KuxJSCdlnJ405PnnvZIvh9lCRz
ro10eBl9RvFc1uv5BK1cC6cVStxDgUgUzWem1VIEp//PQoorE3qxskXX79K5EbJ9
l2LbzM2Nz6Za6BD8mu/LI7rrJ1Gmc7K++9ZkTF3skQ3S3p6VEkeFrtqg7t4oeITH
zTFM8Hcjwrx4nwUatKHxifTcfDm23o56HuG24FvvGa7WNziRCi+KJH4MYA6RBsIx
CZSYNhnvYStUUF74sgfLdNhUrfsE8aBohW9RQPxXtDAYc5H6Zg42fECT4Onae7PF
rjq+z5uZpL2JcJfdfbqPuTU061E/snmsxejYVVvxJZRztAXsd3ET/jlxbg5KwGr8
dgPnntbguFsiozB/BCFUslVzb7ORLSEdR7jU4NOTmRLhLWE+NfPaBVUw99TmiT2G
Srf4tBpL6g3DC6VsskQjozXfFXP63RVCUfU6ZWZyKamtRoLC01sBqCYb96GcZcry
Ot7lXBbgvPC5OMHH8Co6hLYnAS1Z2ihB1sp5y2Nc7LUxWT3Tcmyo74X6iRZKUKbL
jVYJ3C0sEywXMewpizQcAmCAiOYiKYOiXaGV0cqgJB25NlGLSil/CDIv/XY4BmCS
IJqNptUbC6L5qLWIovuzZr4MTkFt8y6NYTDwntKGn1YgwnWnoi0Za/WqqpAB0jea
D+KAr7TM9gcIhN2QefwnF02PkDplhF0CIDBvJ/ycMF0UHz/fM3teP69gaJp3vWxk
KN2ILf4UgwwuFFb9zUoL5IAtd++YyqGOk20YsIz0weQT1ZcjhcW53eddQWFDF8cy
FSbFjVXaTTUDG517+8oiqZiZ3/zqxUGQjnGt56jhyFbcidivdul+yG41jYd1eAQO
ur6NmRTcE+uBSl5dmjfh5tru5ePRsMHcPB5ghOTFJXh1gQxfKtHyDaIBqM10tBtR
+m0IGX6NP26RvK5ET/SbSGlMbHAQltf++FCdLAM4QCPu97U9raXfQ84KdLgWgKXM
C44DP0I03D20d/jwmAwzxjsVNNMgWDeJw6SJDMdL9PoHNCJb6Bcw2+IbIf1YFE+r
uMkc00wltEdl2R+QDPOD/IEqLhi6pdavrqUOZr0ToJq6JsFHqxgMiQz41CJ2VpZ+
qP+lUm8mxmGQwFNQvNHNDVSv/nOUS3PA87BXxHxQbz6B9U012uGFd0oadkWgouZ0
zrOBFsAZcaPWvG6U9JBzrYTqf6vSDl721yj+HLvPPhfHpDxJlFKrts8VTR6OagRp
OtXjVq+ZR8Z2sQ+J8+bYb4OWcXgD6qVE8TwBY9cK60jUVV6VoJOP4qz3Sra1t9/c
KQzPBqDiLEEy3bgKPfCYZ3Z4jq/gxADd7C53HvKgaHlLYFn5SL1d/em/Em252o/A
QeDrDJbSj3Md6lIb5S+ajeev3xE6aGBlRN2WUYGB17/TyI/lPYzAJTHrnQGLPI/u
o+mNNj6VQWNE37bDbxScEy5V7zmSAwfSg0M2FbCSk2aUtdsiST6+b9S7Te3Qcg6c
qOE4EkPRJ4SRVaX+8Pnx5I9eN14bbwFOLIX/XpoB23ofQGHR7VlYG+Dxt0w89UxK
C2HzNBnTS3KP7aNe4UYT63voU82hSU1mXQBc6QMckuACJV8aKSxkb+hEvK2Y1nVv
igJopKS2x8CZZU6wEyw+Z3DTgWksV0Sdv1cAn/iDnmKMirVSP/acyO07RkFHFXck
J3pB38H5kYhEfbvdd/RPgSB+V4SjI2QFXkK8DmBxLHgQIg1TsdFV85XLoFVgP4W3
LT1QmomFf9GbQKaiNUn1y8W4JkVvhRxv+5FRP15b4SdYH2mRJo+1zUY1drgGrpnA
cXwTa7eFZet53ZtydZyCipHK0kcDNA47wNsPamzYeY8vgpggBzWUprdyQWvGMk0Z
9pQd1GSV0rH0hWJY7U7nJnk/DPE/VMTiAc5T4KcgW2ZYoTexJGYurop6qYsSXRUn
fDq92O5vSwvxEeogy5osSTgNbRecti1MM4x2fmq+ReVSEcc0X2jltiM+x3uAM9hz
mq3+Gdxki2TCFnUuybKLYaueH42/cJGL6huwot4PGgrkfDB/kePMO4TIduu/qT+B
8710kpqjgfEl49BK/b3iHLE2qWo5To88C6vOPOShKmndfAq4Yjp4Tun4utnjW8WJ
wVyy8wP7KrexbePGbuDuyZv7vWl1IDcSC8xEgBPnmwg9Ev3ltcEfeFVpjrZrYPhB
E5mcHtVR8BuQ/305/cmUDL+kQWuAr/E3lJ2tjaEpSJQKSm1k0GqMygEL9ys5JrFF
bAsbDGLxpQnc4sO2miRTSbHbnsdENWksKjSNf6QKOIgdrXI7mgeqHhpOkOM1JREq
yl0yPYag/IGz1CeiOsSNmL7tHhL0lTuLYuJLx+poa541/p+LdySb//2d/r+OsRNu
VCgMS09CWM2mT1s8Q6954beT8u/58/fUg3njscuP3QkojlCYUetTAy2KQL7LKopb
4k1HBAcMDCVg/IGwMny2AkLYehNxBG95bEu7W3sLLtKLI/rI6XwXMXOs+1uoc256
hbjm8MNpzytXPtKJfjNNr5DdhVzQfMXwXxWIB9rZqBUAeloogzmDjkk2H6/3+ZlJ
TLUsuR22D1h0h+kjsnnaWEez2LIJmsNg7wXbhPkga1ZyaOcsCAyb+/nZAmHa/KRF
vPl3kuaGOM8ZtGf76fp2YkAQHac6DcylOZ2uFvjIAdqfKS7Vzbjrl11y1JA1hiRM
A7FpqQ+EoeN1UE69Ai/z6BiiG9TEHizYnR3wkibClk6YbZ5Tty1BgYXUONSsvS3N
24lvQQ5zeXr77WqY0EyOMuN4XG0HoMM6BmUv7sdBIPXj6HmjqN79SMwc+heLa2dH
Ga8Dr3y8oMnTxW1n/qAOO6uZ1Tq0GTj/pl7iyxsSNyME/c8qqHIaZ3139ebRQW5X
7lyVpsPrAMeD7WtWg24j6Ce8+4Kgijrb1mGoSkGflwldAbvXIZCred6m/WqQoVoU
eK21ECuo+z5EUJTpQyhoNyoOV4x5IyAUUhwv3ftddF7xjYTgHGaGNgdq3CRJTXt1
ph29x4K62dORQrhU3nGnRtl8Z2EhU36dIUSZK1LaHqLWqR6v8BnB9D2fi/8SVeb1
QIZuiDEU7ypFoOKkIA6LnLEmOoLmR9IiULl3nOpV32DUu82D6ROb7G9MLgaRuB4a
/BU5h+3vcthJkonMoh1zWBiPIIYTOrbJQwX7EdGbvnuj3W/6kz7UhpOH7qXOyaMN
SIlVKhGY5xBdXo1KY284TxoAgepeqR4PmJCIKDYKFVNHN6yKkGz2EmnxJh7WmyZ5
H448tlvAc0S9Cig7XFLNrbDaA5Gnzie3pDJNWJ0sSReUD0K7eAqw5srZTNqujK8+
y+8jNBpRSCGobmXXiVflg77cK2t4ELns7yFnYfCaXMxIBP1RkukmifHxv4XJfsNG
0uc0K1sV6ylDpGVpPLe/b+lpDGsV3TDTkOdmXfjiQ7+csTHH1A1OFyqTSQhb99o3
hsSLw/M+hkOZHDPjC6t0EWfSiHN0NZseA3N1oXsYtA+xar7po0qpSVOmKXCUtEWg
PRa/YFRtzpzBKjVfjq7k+UJTstWtuqvrn181B4W/Kf8nz4XsiOKkP6JJRTNAl+0N
GToJYESb7Eid89V4M4gC2y3fR6Po3Q0jKKZHqsemI70bN/P0r/rL9g0ZRnQC0d3F
xeWlTUGrVKT1PNUuH9vwlPs7l5hAACQlcg/07QDBER03xt7F7QGbAJN3HMb3EJKN
U6IIGjzLod7jFpS+aZO8Gx7wMjXp+PocdUBhU+apD8VPs16DhGCicQ+yztg9EBHW
cMMqdNswdpgufkiImk4PjbeQr0+3aQffcwQLYZ2X91CSh97ZvPfrEEg5sc2csnsG
2zBmKttvCC0ENrDVYmx0gvvvyYpayRjB7fLN6rJTuyPadKqbNSkZTenpO0uhxTeb
SD0c1qPhnNm6sS4d3IeFlGza58DWDH6rU1RmoRGN03kz4bXRq6xwNcKQuQG2+q16
Q3zUeTiFH86/e20JdY0lq6lBtZmYqrEJN2DOsleRDi4wdIvhqej5ZIGnKqScWuUp
rqaarwzOuc8txfZRMSOPPJF57w6lfzcnBX0gqZhs1XE6/yXUwy10zPrOwCf1sOLl
11KArlTg9o6lENUr/3b6ROLkUliEXGiAaq1fmTAKcqFa7dxFcJhGEtDNpqk/+jcj
td4t78y4jdqQFFmOkFe4jIHLQRP3tgI0qlXr7ijreJLxjSy8v29/oRyu5IIyUU3V
3fIwcN6saH+uWk5nJ5zDEbsz8yKaWPBiNemowwtjHS4Z3ap6GnPy0ycduAuQztiS
US9AGS6v22OsrGU2tfpNieDcQsVsBem36I6QocDsPHsEgvq7MRPBL833zCsBj9lb
4C4XXWs134uVBYRK5zxuw1fIDFM8kqx/8tk197pjxwrjt9tOqIRgVENOZrLddId8
L0NFA/Ol9FPuPSlSRtw9LksOlKUSBDYmC2dMeBSMYhNF95Y4aSRq8S3fF7Rb/1Fn
T6HqLVNLrQWmrS3mr6IPQuuiuyMasCFi7Xnfl0KuO8vs1D8RW4i4Nc1FlTl1B59j
nSbnpTo3qC5NYDybIBWU6tLDOPWA/V2MQ8ydkxmo1L2DLRn3JTJFSEdc1fG70fUb
nPiUDaWcWJX1OLl3PUqBX49Cy8lv5xhVmiGYvq8POukiVWgYDB4WwNnGmT3uXIzK
XwJJRkYrzUvCJZNfRfXX2IzWuyj7cfCptyKzSXpzK+Vszcmt6nkhYwBoY5t2beEM
lqv4U0ZZnfoScKvbTHqD9hqhLIFHG2q4VFLrbIXfAiFZ5SWoR8a3GY688OL09LrR
bhOsVYgTJ4Aaw36RyWHNLuVL/FgV3u/dy97KeuyAVJpQi4NkDQphnXI+euOx7WEO
`protect END_PROTECTED
