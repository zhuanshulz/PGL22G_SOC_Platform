`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/x0aaOiZxpjXOMnqudjzhlMZUcaltZe3FZe1nLeicEZAlREhZipY3UGV+sZWP+0x
4kyJfSbQ2LqKm4KumnL43IdUdSDd12potxgjVRFvcPv23Lv+u6+B5t8M5vzN9W0+
KLAydwT/DT2MEFKZZL2M+4hTusNMF2SxeNddL2dtB2qpUrcUBRICuuIWR39hog/M
xw5DqTt8ONfqVfH/svyBYiijq9LSUb21pIta6dHIofkJ7RISiJCI240FtMhkKj6g
H4qItXsltKAOrdt+SIYPMrIzzpw3t1PHPWaLBMTzVOlP0hdm6+RNv/dmpvsMT6wT
uHZOl6xv9freG4Xcgsfv3BXzK5XI6ttYzK97D0YqLk7nhdQopDu5btx2a3Sk0jvT
UCR0hxcl3XZzhwR6jk1bjZmCPspRzcDHTMUm+uW/Oustw9DkZdjJSqgLrSjTRBwP
TcYFUxnK/b+bJQlcKAfVhuz0Tq/WbYjSGufc7YdldZvcDaHO5Gym4dyD9SjTf6jQ
yfHZzZEfXtx6nScTI3g6CqJ6Lnv9BxVa05n2sj/qU9SfjrrB3pneY78L8kJGFmsv
AcmbQ3HLuCW4zXfgFaUjCg==
`protect END_PROTECTED
