`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LwGHQV7d07BRJE3oFz+Gp5ma0Dkz/DiNjJm1NX7xIqxbk28m2BibtRx2DrE6Zpz7
jn8FUqGBXSiupjMMx3a8jP4VHPp4VxuBJsniZQ0D0NcidfXFQ8SiBXwAk8Io+a+i
DMzo3DeZr1LaGuPbeX4PazLxlvyXN6NY1SFA2dqtl/mnH6LMeNjbYzRuUdoI9pYN
qU65FmFz0hB3MZoab8ngbyFIhmDsfd3BhBmEvtCk1yUt9Xpr6Z1RYtRqCDw1X6WK
wan+X1Z0W1NRUKHjEQdrgXldbdM6EkbJWZMHfcarGj8WXyNw8FOxmqK5uJsd04+R
cw4fLEl8PhyVMn5kqOggbJnHYHBTBGIBXOy22JYQNwh2EQbD+oNuBKl0islPEHKE
xZGfhcif/HTXpYII5I8l7lX+PNct4d8Ne3Zyug8y6s3ByhWI7rm5wdowONAeDYPV
vmhwu3tkt7dm9e77GyXKlv9VylIn+AYKjAy5oe+L06rfMR5lLoB2yj0G47LUcYzD
`protect END_PROTECTED
