`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zf0lMHpdn+dRV9jJNc2VTBKOsWupZTjChdH6jM9d9OLeP3EDePsOU//iDASxY0KI
Jl2dXdoxWbzookVVSzku/KbtMcQSxB8OZGBQ7DS672OyrsHOJm2dU29Cu5U+C8rO
wJqvglcBVROpKMhW6eHp4LYWMWCyJqUXCMD0zkvEfNqJvjhyVDcqPjaZ6jJ71jX9
tEfhbU/xiMIPTgt82A5LlLd/ygkwqfkPG/Bqrwz73FzVVTDo4mFtyKy5mYxs39jr
UAcBVa2zemiUimUZXszlDWsM+eV7WoS7ManXNzamyAx+3XHykNDEEHwUW2gaGepC
QptgnNZaUx+C0jAKLS/FI/YIip+1xSlBYqKcI9w6xqzik7umUregCEPhUBM3ALSP
r8PToeKW+ZcGuMREiAyaHWeNRSs6lOdshPcMb0qaPv8sKSZEkdIbjJig0dXHgia5
Jurn7risQKEqkn1rnC9iTtf5VzAr/0QfCo19uYA4dN40zLv4FnGPdMfc9AdMUwto
dr5t7zqZ51Rt5ZvGrWc5BjTUtiqPt5hdsvUPEbIPw+5CVE7/id+CiF172lhCk2GV
8rOgmAZRkPlQlQA4j3QPG8tsCQFW6Vpi0rjYqmqcZ4niVdocbmPbf9apBM2hdyf9
Ot0rm5PWN25VWEL0VGJw/vQjqkO3X+dAlGItfXV62SCChSI6YF96pzvLqfvhpVgz
Pu4kB1ezijLF+xPnZFk5L5bAO2emuTvWjQE6HwqFFAqSBg5NgHCC6YCvd9clowRC
q2CsZTNQ77D/Ezt9SLYmB2mKMELOPyGu6jyJd5Hj41cgYJcl4BHW2TTpDODUctIB
oNYdBFhE4JX3yKws8AOPxXRTuxw1UGEQmg1AN+XJp7TcTgvenJ3UTz0ymqmvKauR
DKps2mIqKqF2pmtFc97Vj0f6P8ZgLb6j02vVsZ3wMSjO9mjoEh3YaHNqWZ7Rzb9E
KxqGHo7FVRucCjtrRKx/x6M71vcJbGnDgc3V/9VZajWNFGB970dKulVipFsKP9yc
QHnHElgYkAtGyd5cp0i3QykcLJaQ4GXU8gUgnJOOEsK0e+KJS7Y+Sm0GYZVcoPkG
fWesNSpaA+d0A2p/Jozv1CtkztKwD/0EnrG7DcnQKQPV5o2gLZ7mfShHEoQK9UGv
9VqorGxvYUOpJZgIfD2l3Qwp7VGT0Sy8RV3w2jRHwXmbNzjN5nwOkf0JcTj4BqcP
f8T/Of0tE16iw1gtjds+QRC50m9n/3w4V7t6vRY7Chl82/z6OWsZHAeGln42DiMq
U6/i6YgGgwcqz3VILhm+wW6qaraoWblgCDjH/2sl/+cbe/24Gk1eoAMRWohTL/9e
6TLL18nW1drt2xFFZtZXHnxYEIgO8JZnWUReZr92EXm1GRm50EabIpSnEhOS5YcJ
abRhqOafSrcvlvmDLAEZDo16PMB/Pxy7OoaVhpf4kN+zHQ182VgZ+oTJgPwoB4zF
n2XbhiIBvIFCbfCQ9p3cWo86G+Zh4cu0LcuGlxilkohes6JeTdAioAF/4sNi3DGN
KAq6vKD7GgAsnNAAyLGGdQZpkvamWIl/i6ETWnX+u73UEvyW+g/BVeVMiRtJM8Kz
vD6t9Nz0gmOXzCa3g2mao5jLxxNe5+U79KxnbA3O0c02KbX+DfV8YR2Erp8cOdrW
5gKVUSUkJi5UXqodMFrpmPap0o3zdjYi7vGbT/3Apgt1Y4uIftTTd3Crf/JKvkD8
3eRTjR+5Gc1t0uiY6fx1bZhrXsRAM6jQGv5da2zJIu2aiyPWFs1rhPr167z+OUQZ
FnT+No7SacRSNlEIUGjOGidGJWM9b9olI0PkqFrDj6ttNnNqws39gsbbvwk8QDup
UwMMqlM6M6anPC1YU9i/ocNFf+u0xseGvkM4Q2loofT1rp4wwrtG3Set7B+MQym4
VSfGNxhHZAMQ9y4rJ7hdTDv/pLDWASJHfl5hHkXDs3s7nefFIkpSrbGqo7GtYBdd
ssecGon0j9pwMHDiFT0iCnnY3EZJyiZKSywWHVCqo5qDcZpZc1DpsBElopVxEPkp
bp4q1FFsWFsT/vsaQgRAQxePaCONl33OUr0nBsvFzlryewRYjm9nDIhuWMgDPRLk
M+sgjIrG0Y02BLMUNh11Es+UYP4ckjBhMFxjhKZR/HHch33Dhkw1CV10ZLhfwiyO
R+lqcYtOJmtWX+t06eRme+rItg+F6E2CKe7yfe5Mydj9YVXzw9QU1fBa4NmIK0BV
yAW4j+ULV4h52w6TZVPu3hJJfpMuFNwXaYqSc5SJwUkg36VwXDSGHW9VqQ+L+62F
RrKdZdDDIPT+LS6+esBqf9tmAwIQ44W1y8Nr7vQJjsgA+JVLTtZcCg5WSD5hBTnn
WU50m3ffRZTR2DvFVooM09a5q4DWnFGe4nR+HMcHsK5yCsfeUsIJ6XCEEXfnx1Vr
rWgXJi38GHCu+ZzYDAXeYc5S+UXMgMjZJdJOYz/SJgThSSIepBTe7aH7WYI1ipyN
iS5XBZLzYydwGWoeTRojTsmgMQ0LiuoOhM75peteo3jWDwFXQcp8DOyucY46dhpZ
6DGIghNpsT2xbbvEKmFXFPfxNGKNHLJvwN+HOXOAx9O9FPfJiPPNeiloyUdOoWVP
IerwaYhKkSp91GKWRykVqtL838gzUbIjWuuKW5AkjJiC+DTvY+5nQ2ei0MYVKHUL
lxZLbPoxrDtzP0ZSmvShmhbEXnc9GHyyAnPzIpSVo9ERCjZy9FXfKsiVzP0wNUVT
ppGaILH+zagwbCWFb9VOZ0ueJGuZleBQeSvjcHEJK2JGFOSrd2K/Ve81jjOz3Fq0
avJeku50ipHYyR6UbWZxqr3hHZMXint5GEiO344sB3DmrLrOPvtbI4UMFJH07sk0
PHptSaL67f2H3DDVD/jPV0uKwaM4mMmrJn3bVboJgyFUPRhqKFBDyc8rmXGgCAw5
8V2oJO1SNXhp068MuPLM15RHWr2Ax7HC6F9x/9URFFIDQnmvfGaR/ZwFPt4FaSNA
VdAz/xfgiw1tu9Ta6iMzBSfRIuEumJubbIQko6Lx8EKc8XixOVDMj/U8v++Rj0Eb
01I7H7hUOKc1QRnvnOXUOJ+3DHNiiFnlkFTt60DGE9cAbCbuxOpN1UGLSzcNobMV
iJ8S2svG7awK3WKdvH+HKc0MuV9HDt+ckiTYEHsi8GpmpzCimkd1E586vukqI9PO
oibnUSjbI11LIIvz3Iko3GACn9373pYVaJqHO9Q7yS7QIsmc/TwqL6EokyyYdaru
e98cZQSWDx8U3lRtmjXjWoghNs6lnqFzsIZR8oj17U581QY7dcGTCztBMsE5FDEv
jb6S1+augVNZf6I2q6OAjM64KY2OgSATTWWA13I3I9EIRi7OFczdiz3uiv8R5kr0
1Aoj+p9CrrEQc1avbFmHiu64YZFft0kxh3ONF2UIilHvr25kcpjyJKiRqkzo5Zo5
1mRVfR+WDfFdj3ryXCLfwqOVFA1CaT77VKuqpBTdOlVHJwVNXWWnfNVaJJuVCIkf
5g0Lk/6p4X7EDGlFK/8GlyxievqnA+nu+GzH7KSDY0bcwEVIC9tfm0kUAch0i7Us
G/LfmnSOtsjYh0uUqiCi0MbT2FPaSkNFhHSvbJYIUDHZShJitZLr9y/k+uoS1Z43
ZRmjEZzLxtGbpCYqMdY6oG4P5L9h5tMS2QWgkaWU6PYi+vHHRqtLKrNh0mBUbODR
pkPaqSmTeynp7/9hTmMSUBJn0RC6jiQMfcvZy9YF01LBwYBr7Um/NFmGEZMf3jGV
+e+l2GtTImpSj2UlydeCx9MhONSF+QPx2sG1l5xQ2vNSxeTrF8cU4v9yhjWvIrql
rPCUhu9JIi8KRTVNxQkssvryqRHyxUSK5lxyt17rd9HCin6fDJrG7WEb2ZOVV7td
7N6i6YYX/sbbyou0g/oS/gyyOMRIp4M9xkHiYD+bIDM5zyDqQDknmskopyZ0BzJg
0tG+ydkbGPQJCoZEN4piOE9ywkxO/pXcnoESdNVE6Ycw0n60q9ZsJ8B29no5BqDC
eSp3RNO4mIX+DB4p1s4Ujb1nDmH/3BdMW8riKk3J0wtZK7N0pyy8ogEbQziSTuhz
kHDWvkgMgtdYC951WHkErVtFK0ufVEmdjzcQnltxDXWaYMsleXPfCKTgbmLoYnNM
W6kcZlFTcTVEgeEevHC2VYycEpcBgVdxhHTDqKN+cLRgTf8FC/g9pjpSx/d8qEz3
PJS16Gf4IeI0QZtSfJQs5ItGm42jWZDySY7ipGevtsYEEo+DVi1RehRDbF6RA4m8
fnXtTyBQrhU0trrm3vMkmfqCIKVSyNHCF0lONCywvflRhjnPVKiarLuzcp3xM426
YbTNkROqPIg9iRPpnCXR/d5vw9bZH0YB4di1vM/z34c0fpnwfAx2er63iGjQrSkC
G2SXe5attjSBBxcq2HZqIVwLXiLflGWykofln/2AVesCBA35qHZgxuezS7PViXRj
7Y6tyxFEocl3uhaxl36S5BihKMuU0ZjnVioSH0oXu6xifQZ/RTbQ+F0hjhK6QuT1
quYDKtzuNN9OE5j7mZN1SDXFmXfgfqY2CKbbjGFiivVvIsKhy+jaYRSMicfJkuWs
Z247qncVpNPbuOy/p9hHz24dd6N2Wpt2wMVjURT0SKwHTFjBnoSgeQ8amPl2kvTI
pnHTDjzMIs8heM9O63Noc9tBaFEZYqYezGxF7YtGm70IaXKO0lPntLC59E2E4T4S
yVlGUyx2n0PoAeBIjkhAwK3I5cpzL9ik5QjiGzDxR9SgOCcLqTT58UG6HyLdRM+J
NWBVc986fcImgCYeOHOBpluuKj+BIg8KSnWWYZsPIvl5i4eaX4hm1ntXnB4fbnLV
oAJtR+a6ZgWaCQKbR2kD2z1u/ad9F2lY8KrPspEEzG0mlOgZI7Q2rGiUbABhdQ0o
YubX3lD/cOqIbEO1ogCIWO1RNIuc4VQ1bKfocNjPWL593gJEnZapdbrMddk3KrF8
dKB/WDoq8OWhPp4kDAVds32bc+ao1dudvQwPGbjfpNiWnpsyRGwpILaMOKYbjyhj
VeXc/8aJyzEVONrpkApH94jKD54jj9wo8CzJl9u4VXpOnbPoXhoQCn8DBTp0yXld
mbSY+J+wCUarpexVOEpMywdb/uVXcoWhiQgitfgpGYgj97OEJtPf7XzcVllLX4GI
RcOunSAcfgXSUxFTdpeLofPo4EIqCkdc0uju2sDd5WLJZrxA8J7F/IGg7A6OpmOs
zgxR0l/vz/Euj+XJCQ/s8o3mQUkns6Fuw4xa+acs0R0V9drY9LbstbI6WE3rEClQ
kE/mK8ItriY/8iGDVfktg+juHngj714oiHWFTpTwejKTC4KUaMHCBCTCGF8pZ5JP
Xb0kRZEPECJekfs/OJZYuhThXSWOCsS8tIwOQVYXCS+sRXNHeiGr7EvSlCqGCScO
MH1XH4e1pm8P3Mcf4ytf8KokuLmrme/A48CG0LWlKRnPPIyYLJRxzLQeGlTX5Qfn
08BEp3+JxO1FnlttJ+dUUeLgi3UlhgFG2bzqcevZu1BHjRE5GAmwuFyUgglyuS7T
rSIXQ3bLcHtCfsntja13c9Ab/OFLwv8T7/HvxyZV0UYgwEvLkVx3z97ncknpkG3H
ZioltZL6mdAI3JRokWj0sS1bWNyqOZW+QFZxKIQoOsGr4xMkt5aHFT9/baq7ARbD
mfiiyqI7E6pd9ijNWQ9pKFiiCQbCVuYC9/AcI4lhtcZHRHIAJKGSRWJ570qezyf5
mLTwVxpcB4z6GP/TLx9r7iNRuNTdQGygyewiGGNFZ1QdgU/K7yF/fAa2rN8v/Oth
X+Yml/hxduo1EtcuyMI+YFSq9KQDlit6Vuhib7ip5GKo/a+YxebGLdUDQF+w0Fqf
SDlRdx3ByeMBc8zObfCHK9RIXeEYXzTjNzf8ZgLCYOlCno09MzYIhGn1r7xhvex0
ETLgSEGTV75rE/ciduZsngqyaP5FmJ6GAjRiGeQ2t0xK7AqBA1E54S9wFdK2iC8o
brIsfRWYPuPJDtZuhQ8nvFx8mi2+pbj2SmRCIWNq+MTIcBfuvzQ/ypKytQs1JRGp
e3M1YE4wSR8xhr0V7oDcn9N2h9o/iPJg4tw4aoOuQX1OhHm3oTMaRjNGc4StPGGj
R89Q2T6xXG9rgMHk3qOfvxVNg+aMw3VYeKBedx9RjOOvQ6A3ZwVfrdgrUFC5926c
VfX8Ok3gemx13pLEHffEgeretuSO77C1fW3YRVckZfHKPSNgvYxTBzhXpQ87icE7
KwAWy/fuKd7WsrxDTR+GKKfyi491B2/UnycgZx3t1fg/1NyR092dBeGQpcZ2/lxS
T+bzVCvy+rgrxJ2R4pop1Bz4DwiBuaHwrPvNFnB3tjdMX9PDtqWBliPECtLBhllC
bxGz0B6yt9v1cRv64UMVSyF662S19b7Kb19+jjwWdfp7jKW/Gr+NlGNV7NdpgeZh
hrHERKhPezY6HcvbS2UL1+PFG8vIl0vkc44EiAXUo00EPS8vdxMEXsHRq5sI5B14
j1d9hvI3YXQoIHnXkZQALNvWLX1F4n1g+mIAhwKuQDqyOaVBhSgtgMKIcryzaldL
1O/4f6N/tG1FVp7iGVRms9AUbM/Pm3MHTHwpuwqwTRC/gRlRlc9+8OE6SsLfWxN0
A/0lpkABJ2xxeOls+s+hpW9APZByanCinZE8F6FOF8Tzvt3NZxaGNDKLAUJ3mZRl
pD3QBl0425/CH99yEcwp8w0fMiNUVM8WzMNj9sxAGssEZ/wRlJTc0kVoqvoMtfyO
htCWrgeY4IIG9V3STAZFYLxDsHYPpmFOedsZdo0VefCT05LZ+Je74e3LCJepy7nk
Uc5xw9D8kxDHmo9GOtJofaPUE+qah7Iwedt8Vorn0X5kxsLMXDht3V2c/ln1Gkof
e4/GUwjEpeTlQMc/0s8jfCY9d43YniiBZLuOGq8GT2eZuoY+BFExb/GiGbsYF1ga
3SE7b2MJ5Yw7P7koErdtxtuFinaciFXVxktksl9n2KJZa0ETlTfsF7uSMhbdwJ6j
PPKyXXL0JgmrHbs/BK5vMwUTbwix0x3BNJrDYZKrdtEue3uzaWNQbQKQF/lGWAXB
6mDKZm4Y1Obu+AuCd/SYXZotBSvJ6apIG3NIKsKz3qPFEEEc1JATf1V6vC+POJ2P
T3YtxXwR14LDtPOWP2eWw1mTndA+PNa9TNcWxVJthwHgUpGqoK3ruKbk8yNHHnxn
D50/9K/zS5ZhsEUDdg5IZEpaknvbOQnGs8pCcxSmYFcp+WsPOWmMyBlR8MBhan9M
GryDacH0KHhSCf5yVPjxr9n89bND0IsRALGp43h1uU22laAfAe1LMDrmCMqhc3JS
Xw+MONc+juT2GDPyAmtwqVySPIKQjCUqk0sHD3d0Q6/ABLPRVjhfboaBB6sLRaNV
/h76P3HU/3j4CSUf852lxW3pue/450SyqTUyL/YmQkgNDochLD4uniV092LFEhtq
V+HGTLlweXYv+/UTa1IUkAqCjZq6lzRyT5Qx6H4z0DjU7ajXTa62oHJTjBc5WGfg
QQthoOdeHwjoNBzZC0zTyOGn0D2/8X29ppVFoXzDxREdue61SMhI6ueewJri7nL8
ZQCb3hsQoc4ssbnlYO3QMq9RJFSJYt1YXcMNuz3i0l/xkSiBBltLS1zJ8XhU2DiX
MDJMapj9uSVVQC7l+lPpo07MomOan/e+aB2ExrFu8OVFSwwNHN/KeHSxxtCGUJ7r
LN0yTU4GZtIY3twQi+orWcSeyHrAmshr9HLogdEJrvSTQWOo0N6vdHK4cbGOTPJv
UnwwLpq13tqBr66AbON8o1cDpoq7gChGIzV+675SJZzyy+jB/zgu1cT0UAJfn45m
q+stLRVyuqhRzg/ghDQL8yXF94Ws3c6wscpuvMwkd9QluIQvO+CV3UMZslLuGpa1
YO0DfyZx2ywROWx2dNal3FeJwP1kYygYoWwltxXPy5gg+R8r/Y0uXFnJLjSUuTZN
Cr/SJ4ZtsRcaEn6uvTsxvsI3sLkGQcOMNoXE6KFtrA1KsIVoBI2Ogrpyfxad5EGa
Qs5ibh5HlFmAbhvTGn8QPvhsA1PP9n+oGqNOKYNXkr3j9e6oKp3TA9zYE+7jczjb
73bX+J9AZCHSixQ0cq81w2qJxUTpNklihkNmoHDL6qCO+6eNCe9DVX9ZUo3AdGJu
w/Vn5DPgTPgFjrY/yuo/19bzou9ZgQTzz7K1Hzu+UmMoypHf1OoSBfbpj26cITJF
OBpDqrPhiF4Dg5MfrwFDO+J6i0XuAebqWw1bzCtu2ercv4tvOZ+iHZhAqS3M8vvs
wO/BtjYFOdUSV2oM1E03uakVji/gdzpatjsUPWiPhtd4VTYEvt4hQ5O2duCfQ1eE
OWQJPyTNxRKem9sx/mRDfDhexQsimijz1yMEaoY75xCqI6/07DEE2/TOplQX81Sv
NzGWuCCbEFR6fEe2ho/KMR60+5CN8pa+lyV2bG2VtPQ++qZ0ji68JSjHGa40FasK
q3ACj3SFpZC4ibCjj3wpw/t+cBh/X60+xcvRDgkOpUG2IMy92V4kIV/rWWRBwQ4C
gobf3GBVmyUiYUQUeeiBunPdn71F1dqtbSvxJ0BPL+xkGvfuXI6WuZWI1hColDRe
+zs6gQ7QgBEViq1oKn9qet1zlgotjQSG768hlqgBiHh8+0h/5IsqqyXEIqCnlB/8
Dmanpa4TvgOga2hIOlZnwCHNFloJX7nfAOaI1Ay5y+8/YQyROewd+9e0+qvC0Snj
SLJDB6b2+xC/rgHwEuQVebC/k74oSUXBLJ5XzaTo63cs0Ezj57gGBcNnAZXegYKv
WN9TT5jkZuQli5FaRhOYzoxAZNqTqBpmfSijyQrJnrYv3VA0P0Tpaj/I9fzg5Mw+
GncdKlkfWzFQBT6qcvUNNW90Qa9/xfQOFzzMjzkUSnrh66me+ay0xkFHUao92gEv
S9/ess4+x+bM8XYzW3Kjh/gxJIShDvPbc1g+N9J/4ZKjkeDlfqQ9GFDgkXeMD+SY
B7Amm0ztQheoD/EwNn13EytPyOr+jWO7vMVmdYBPIV84Xw708/ZhzHrxFAq590aA
vOFb/PXSeSDFHRajqMIa0+qdoi8F5YivaLyHI39amYLuvD8c8Pj5/fSXPlg+/a0e
rf3nRbS/BwhXT8mRpv64ICDKvnKtMgRkZ6yznyaIjh4t5sZ0ayS/f27Ntq9nR0q+
n+IDobUc45NWQMohsShj2MglAB4DMO9AqusiDdCOeMuhAIF1kBKffX2eOeY/Yh8Q
decleYpifgTNQ7qNp5uG+phakglDT4BGwPr3XvGRXOq2bqEJJVJ6mwWa063nELrx
gUiJ9gAik4vz/2EgsVRseWD3o9z1BSop98q/POHBxtCIQ5UKnX0f//f+Hr/LUTsJ
ogWBkd3+HPG6LEkCLaRAVFuln+iHSnL1nJ7SGKgsP99KCCCcWoVyRTNagmZvyPCS
TWt7P93P9x7ZtpUU9N2MZHpGFpr5Hv2Ff16JrQJM6+nxisyPPZYGYI3Ezly/ipiS
q0hAoO1ryvR9QJals1Mg/v6fI8xOKVGihPU4npWT4LwhyhcpWj6z/WlKJ2HwTURS
mn3OhSqUmli8xE6q9/VpGAxcGdOM3yx/xZMn+oxbLV9tVI7kW8z3QBnWKDnQzJkP
GiTTp9iAAHHs81E6qMB84ACgG16Oz/A/7AlQ8RCECO+uyinu0BjslguDljabLHCt
A0uLXP29kltqzU4dnVnrTMjHIA4KyklUQVplE1FNmcDMov+Ndp+8DdGY7oAJ9b+s
Zf1QaoNPO5X2bPx/hCaHN7b4tJoAQNDY4yPG4nhEp+9kaVyWPFON+OjoAoehwoal
HITox26PDoXNNkh+5s/J7G5QZVzX6XDZhO7xYkqx3pr+b4D39GtKKNM5mvUHL4Qi
yhAV61DmjpLemoPu31yc86tvayqjZ9mVx+Xv2FZNf3l6WTm9BOS+4cXiAeltb1uo
nV5PZe7fgklDkzkyQc6VSx9RxbDGyReuSowYGbnuSd1f2OBGh0OZspcs1/yb6Xyt
awB4hjkIC+5edMnddi29TfRCFaWtPsW28IB6mn1Iq5lQVc0IqR6l/dL+TteaBBl6
CpIcF7T7DDswmS21KQ+ujD7Zkcm7N766eLekKIs/OZmlwFzahwmuc6NQ/yiCCML9
Z4XTZ7UOwPY9nN5Pj3/wPU59TmTHDbnv8gyoEZLQHeXK+lNdawAn7PLT0rML0gsp
38nXy6QsLEwA1YioFYl4hq+KfmWNrFq4mIZuwOfQEZIJBHxsvL4fnZrUSjhVHym/
w98aCCA6jzC4Xb7fMhRSjlmrNblGiBRpOJiNM/XBFPA3RYWap4tH0afDyDeaWNrs
uhWxNMD3INOBbOLcQr536Jkg6iq9wns2ghyylX2gYo271fyjw1OkJ41GHBCqyOCy
Nf8aTpum1qXqNpAFWY0opHsxTPaYBhpdnM8e6e2pP3F5PgS/FIhkEfld2WzvLDnX
7dmxHfp0u5ic2azr+Pvr8KPsB3QUpSTY5uE+IhaMYaSPR8fpcjEozb0EgzWjYTZE
bNI7OAQj+XwkBMcj19zxXW7mE2ADbdldyGdUWyg2DxA+jGZvuGpTXKnMb/qEzhFF
GmBVUngSGoVo+r7wU1tUZeQZdAY3ZyCm6waCA6enbYb688+J5in2eOzJNCHPzJv1
B6UlELixTYRYkFf2wPG8ohO7WJ3f2VGioRTAc3k9aBzu3lEcKnjnjfPv/K99l9Hf
qVJFkYZH8OB/6suHLXzW8Q4IQFC/bpfMgAqcvRMp3TsYq9oyhuCLvo8fYqmrwvRn
tqU4hVwWeM/rvYjkDEJs+G5bV1SsuO0F5wLyzlWUlUW3JVcE4ZDTI+Pa03MyAxgg
1lQGKgLRpBr2hym6Qs9bgrol7kW08PdOSPG9Ez33aAQEz5Je2GMUYflmDW6QXXG7
glmx7wG//lTlnyolZU7jra4ge257lWGrkmeIz2qZvh7ocYOATgAUT1uut3t4FOMD
3zFuktt3YUnPfAw3djDLg8p0G5ODTHsnWZnQ7PTXQV2PgtFgZg48iw4RRP5W/5KN
7v1VzAfQwIHqtjUzIQ4XhJxAmY7FvZBRvDAKKpF7Ad8UCkferxTnbnswfYA6EKRW
oRPIh49OEQ4+Nc8thmODO1RyOQx6dexwoRyUcK5dOLRI2Je977d7ETI2IaqxF0iP
Ivn/FYNA5xfWY96nqFwQhzhGrJJ+XycYWM0jCwqGu4vyyOsbAV5Ov7XF8Hca2Qrn
dqd9s6ncmIdmAr+xssQ0SqPNh0SELBw7A1TUyBx49mS74SmWGYtZvi8jqs+VyzHX
+nwfseY4a21t/iksotDEXVZLrAviHNsBoGeA3weuq3PGVyK49wlEv/BM58zUnce1
QNsc3CVJlkFsoH7WtxeznpVv6Vh/EFhaoxfTmf1wOdFFCeqRjdkiCw3nk2HxQmec
3RXVdR8L1OHemjxdK4auo76vdpYcl9Fq/YMTF1nAGPUO+WVQlnRCkXAI+UrUk8k1
o+/8TqoR4HJmbAQkdLM67MHR33qd9vWmtsqy+6T1A8LaVgBpJDoZaGeYWQHA4HFZ
FCLwVjLijBYUY66Qm/bzRnYMc8E+5o+SFYuGayVVfXNPAwmcm3iGnUG3VTjU9evc
NI8e27BGsokZi/Ytk1RkqbUK/blgZBZEFtzDSkYhRWEWUjCwLz9ieBOjMWrGTokH
oVtQvOWMRhe2cDHXUyYrwJydNWvbf4kKRgqy6z16s75kM7q45RMJ8VwyB12FOtiz
EBZkIQwIFmgc6mp9SYqaJpLShTdtuM7o8+OQLXo1dO7vcE3Pw9Qiq6NZUBrbNTMu
2ZZjFKyzz7vhwJVOa8jhWIzMC6ZbgqUZiM4aIUwUkmv9kBHRXW6lu6o7xJn6WqTR
suW24Q5G6aTMJ3uA8e1UgBkdVdQPiZFcGoa4Xmaxukg12c3CzyO3B8tnAFPUNygE
R3bY2qI0msXAT7x4JF1gM+XRrLIdMxPJCsCYNO9dcKoKWCkpYNV+ErFMOgo7FXzq
F/pGKUSslDM8ghiRLtv4lUBPE9fi/XTuPgXoS8sjE4sF63Se/TAAqMd1DoZx/gEa
2yPFnhuYz2bFCkH9ZQo8NabGTsD+3zNm227ovJhdSUZs/OkQAV90izNmBIBa8WmV
A2qDPcQYzITe7jBAxTGLTyIEhYe9J3F+GT27GTO/jLv1YxzVPDQPKfo1VDxSJrlx
iu++2u6yHFfhPwyWOmQMcph3fuIvx9lOukRbXVtWmvFPaPGZEBpEUOtBCkqzzyT/
lXoXh62UFabjpKqLVJLZG8ZZkO7y5lwmaAKImQ7LmEdhit1JABG5Wnf6898LASgM
ALPT4hKY5F/S/GLu8ZcFWx0kypeCTO++9GudIEMgx457Ff7W4I4BVQbcbw/Q1BRw
L1bMmlEkvh1EvlFcYse2cN7VFK2NBsa3UF0/CeDUIBteWd8sa0x//cT7wu801AuQ
z4ml2TKkQZ2YR1PZTP3kXtytjJ8TWE6/fJ2/LH5t082STVK07KN2Sb9FPJFpuni2
VzSTnp9TbN+b5JlMKuLa5vjvp/3uEwJn8Yx+sc0P+8/muwgFxymIkIS26PkbDQ5B
EcAvvqOwpk/Igzn66dBomzXUxcDN4l/EZ1nmE6zPc86Ou3IRpcxQLEmuEBRFIDKj
Tz/AZmWTcwuqdhs4KwnYdcMwDCQMpR+AuXV1T0Q22bsUDq5a2gNOC8dKdDrV1AqB
Nhro76bWEl6cOqQYA1z98hZTLYDvu75MmeR4k8TYhCcY+xuqrfQ3ieMFUbGz6mVm
W6jBUM42CPyS22Whp822jJT3GFxurMUsaJ8EQmpslBPXV2ETew2OuBGrcp0ZlvIQ
+bkX1epZmgVrNltCu2ToAzahTBP1WOwsfhpxgdJImHMotyvSd1nJEfCifcQTQPk2
TJwA6kCmnRw6qMZXng+jQ6TE88RdkxILukdntgrFfWkO55cBQUrW5UrK3M8HRGDi
Uuj06ZwnGc7AB4CnX1K9aq2aK27QhOOaszsvkMuUpPNAIS4Vk8N8Zm553lAoxfoV
UIpxVQ8gLtpflIKA1605YxDDLNEzDUPiT5S8ZoK1HZqqEA10zKb+gMeMWZ5DdvdY
JB/vkZHdWhHg4I7OpJxHu/E/XXdsIz1T3RCaLY+THOeg9TSwFve7JkSRzzTJQJte
Aje1zGkRf+lkOZ40fr2eEySi3rmRv79JBeHnCaqHLAgv6NpfohkzmrIugY32qKgu
LL6n96ZBLRjnTaZSDZ2th84a/ANNF+6pUUJUvB9BktaLPf2g+VBDaVZSGPoDJKWs
LtZ7gXXyNVMdJm3eiyL+X4425WmiVMPh89b9SlQVmtgPQt8LVLXsmqJ4+Pb8bw47
uE+gByA229ulQqin/u/GIyRi+mfe8poOklC/o81t1qfTJT/f2lVSSI3IizkPg4Sr
o4L6H3tp0PDv/kqldF7WAYxiakVQZr8CQmxlENEvImlnTnIm/xH4u7lc0vyS9WlA
8C1PuTG2LelHpoc9FJkIZD2uK25El8j08JACWV9yCsZpvKlurvwsf3eiwmrMPWtI
Vd+rFV2SeDm1xQRgmoP5g3TCl1opwPXsdvxi4tUK5O97lSgbPkUiiZbpQ7ICbp1J
SzKNvcsIjT4876hZXwVivNMHHbmZKPFFdbTK4GllPG81aTrHTneFZ76OEf2hooHB
CVKdw0B6mPNsDG//JnYqU5lHRsTF8qoUAsuwNIFgmhMl8cmdHG4/lO8c3t3yKOs2
y8/zsO2hAFOv5FECrRgG8bfTq0e7aBtgCgTKoyHX9Tu0FQCkoM1e7FYx0sDZZgps
BnMthdW2IVCGvjYLxZcY4E4iAXfgQG1AA/gxh3l0MiatKh4NYubBIO3oW/lEz/Of
x80+sN8uAEe+Vwsc8JQZs05QuKj3WQAwA1hcQotM+r7/teopAvl1KwRUQlnHHpUT
Rb+Aqh6x3ySFztQ3Zn/zzgtCH5hTEjckNjxZ21igC/Qi6J9nrdSTlsBbMOs9mxPv
EIRXL9YL0UbwTTFx35wyCQkEsByJYhk8eICplTFjyTye7qgcFxsNLGsIYXzBEBra
Zf8KVb7ucnkU46jnbYB+43NxuKuBbmlou9CRU14yWWl+1BTjBam2rdLnEGBXU+ES
V5k0Kre0ySxEs8JYkDSv4WPftpRVTgMRTqpNIV7icpQtQ/OY8G9NrKodSUaD9iaQ
1fShHcWoH3hS3W544+brgafnd33RJWJRVNJ1Sxu0rt4rdQSh2/D5gNFCygWCaNS4
4Ap6VdvUgsyF6wOYG7AqJfUW3a6ne/8c+xywPHzRwCKNvgOHGvyuBrXo6da4FyiX
hld0dFz+hNM/3/E1KEbXt9JI4I4h0nBNqZD7mSC3eov1UQeGX4ThaRudXLwAsFG4
fc9UQ+6xz4OEtgIdNP2jHmoppdmehoZeaOjDTlWz3S6okxUuqNf82FI7X9S2VZJg
eqhdtCmWm4mp1BF73dN7bCyw0jbTRAYQ+l2SmIAO9+rYfnzm2ps52LwupvcYuckE
iKgoFv8O0IJ6XZctsbMqo6QOFSy1T9jyJFTOhDZUx6oZ4gmfQWlPVntfDuXz5nKg
wI7virv2cAAPmnCZu/rZqkBbFPL7vUwvD0tryWjWAdI=
`protect END_PROTECTED
