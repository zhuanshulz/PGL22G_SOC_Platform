`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KpNBHadC//Hl+HE2P5VD5fYHc60hU/iIM4FV+1eReHkq3RqiF/2x53Po3mNkSH8E
flPMwPmKZ0kXRZcimAA4iV4VvVuh1fSC06XYH2TDAf9l6vmVa7kSDXBnnzHxH2Ze
U39/1sqp7kP5bN6dXjmNwFC/ns4LMQs+6g7jUHu1jer8ZFsruL0eL8hJeNlNxb0a
83BYCKHOcEzJ5odbND5nvb8tLRmkI3QzUOX/3q1bJ86wJFN1NkiHpXU7JTXkW74T
3sU43pCXWlg7wh0rkFhwJILSV0buvrZH4sika2j6Bo1cLATJG38SnEZZtmN2YNlN
ujfV9RqWJHyZeD3r5RNldZ2QdZv6VDzx9xBA3y+Uha7+f6hYqQa3RvNMsnmz7hiA
HQLAzKM/DK6dDvrncG4h4rYuTW2X2mph7t9LQ2CKItBB/a0xTMWBikFG/6ZQM/fC
Yr/eMXhstTfTCNGiCnJDhyh2vvs03mgRB2Hs60D9O5T3YFaEvEdyQ/SaLbtD6dac
xQQE+XmbXFktddwT54tjj81uVZdl7WaBl1eQvghBcRY2HeLiVnBJCsUecrhKtJt6
lpr2fYQ9OVsqKs1sb5asV8/hWksMYMQcWZRr+qmMmzLRkj0FIxJ0k0N+Qxe8IA9Z
CNOCkFLYNdIH0dlFHcAcZv9G480zsCDx0yyaKlGw+5pDFkozrqlw9PjmPdNemfZh
Qz4kSrXoi28hLrcPCEaf/cBu0mHcBsCic4Ov2gJ0Lox7YDZj+6hgUsRnEGrdqU7p
0tq84CRIs0iG8wL7jO3wVQ==
`protect END_PROTECTED
