`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ahp/u4ahsrHuZ0pgJNeyeW7Cy66VxsMoAErxJjRUQ1MDDG/K1cXgdfcebwtlqO2I
Zes0eHskWP8wRZNrOgj62ZVdn1nde/lau7GUxO+9WzGkTMloXa/XlwMIwfBiPwGU
mTo8pHgW5zvmyZNzHOTnI2y53cfBBLaRWCbK1Ee53OEHQ9+W6GeETV0jGtr9Vheo
j86ZxDfnAN8H5phqzM7HqtVf2Cw2Ob2TJiZu3FwyXzFJAr5x/FZA13Yx3cV+2hqT
s6DVFIYKiwCY2vdjUUt7Phj1oZ188G9eO5JG5EjXBUk4RbEN9pOO+QY0/ps8L0aH
`protect END_PROTECTED
