`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GE2QYSXNY6Gr0vn9rmrw3R0NXd4t45VLJhQSH2EY+mwKA9gprBKf8SAp3Ecay/5M
9fz8LYLFa4WF1DgfZpaibbYEHpNPI/BMzxZ92dc2AdEfgS02pIX9dlA4u7JjHYRD
B3wCOhdt+MllrOM2cCE/ujLVENz8MHNnZRuIgbM9PJKt/5tkrP9G05xd+M+F0gJE
SQkx9eitb5Al1gzy5wM3sb+62a0a+VWwQsM5tS7hirGUaKQKhizDUMtlFaltXLIp
0q85Tys1g7lpKP74JcI+SGlXnuwcquZrw9+xx94aE7+FBkHGtyuh+U0T2MtdM/rH
D5PL4wleYaT2+Krae8LT5G/gqO2kGJi4pjFO99PTYNBJPRcthgDuHnb2YiFKzcf6
Nvs2//9CVazVvJu3UqYtIS2uxmG2/4gsZh7Y3UgT9cbmDdjDwrvRq+G0cH70BL4o
n8srxqSlm11Z+GAiy5bcOX6IYoCToNDLBt65gL64GleIXAy/sEvy2iuvoHcwNOEA
8T2/8qTMaSJmiGCg7ELBpQc+GdwoOoASaGcFs4AZ0SR5GHKkuzlsVasgf6eHPdct
+HVQkPyTBwAGNw0CPDiZfIDK0E4mcNf/UVvg5zE8IY5RcKGsVJLa/sp6YtYBpLOO
YqGxn0+Y5rHgFjXf4YLn/Dtfk4A+5a+hAvayX7PZNIbXV3MSoLR/wRYUvSTzz6q2
KkFmdVL4taZGnuJ2LgbxQx7cirLfvuiWoaO/hMGoVEDH8Tecyb0i+y3uIyZUJE2a
62uymM+oHrj2IlsZnxz/50ftI7MDHTOK9KtnP6E3TvK59YzWzmqfFLG8hHgx4Bi/
ttsx/axAi90ohnrgDpa30zG44XZFrFwg9tlHyKVOCjyl5+DisG4XSZNYj1mr+9Pg
jAQD2kJ+eefTup4aVzmkyMBlx26K59l0L7E7D/4E+XqpA4dWHoWKck6uEXMbqhuZ
FaNGwV3sF95F665BcSq8WnUm0SFEVyAg9emB/yjoSIYijHcLeAzijwwIC4cZjK1q
gBnoTW8bIdvt1BQpFzgjcv8ehuf72IPbPWlbzYdr2lBBobB9HOavYFd0YYn16VZP
a+jSAnlLbvTRZYpe+IIfeqnHmAHI+3g53n/bxHrOc2qSU0ASEN/kZhTOHHZTNsP8
88ArMyd1h2jTiR11Z4ifXVWoTJt7cmbxyg14PGLl/wsBOqWL2J/0G6Ef7nnQccuv
Cb78t0Cb87fnTOYwEQmXFLpC5B2i8+p+B548hbJKjs/Y0OtBpgItNBFs0Fxe3P3L
m9rnvFhf+X3ZbS6gBcIKhpYczzNUm5/5/5fNGkb8LWzcFp/t86yQdiGPNGobQq29
j5IxEe4YhdP/PTVHNxm9b431UhdeypAl/z8nDVHLItkZGmDtYbLa5H9GjcP+YXXi
DksC+YjbHjNG7N7D7J75DZCTab8ufhXkar2jSuBmcLI=
`protect END_PROTECTED
