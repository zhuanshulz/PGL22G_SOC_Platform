`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ycLBAMu8Qg0cb6cVdxSHgktGEUuWd5/Q9AyBq+govF5aHSyAw4J7U7quygjfJ/uo
VZBlYZe/YFsYspKx2GL8C09ERcCzltscAczX9EkpmsPvlHK12+VbpEg3W1B8ifGB
4gemy3PulzyMmk+Dnq6QcVKyggpvnG8Dct61thBNmJT34E/zr7UhjX+kN4hUt4BX
TIDyGRfnBL/YEd4VldDJisbOB/VVilni2tL3rAl/XiJjj9yhdxtC0Zngpy2L7cCD
BuQauQ45gjfE8PcXSoVSahdH9lDrwpfLePkQmLEIgwnDKI5hmGGD93OOetj5f7rJ
+VEun+o84j35ypjbAW925wLVm/092a5pN9S0hlgZ1HH4vvok6ea7O+Phw3AJPQ/n
3dg9MQHsKkNnUKdqfcYUJQ==
`protect END_PROTECTED
