library verilog;
use verilog.vl_types.all;
entity INT_MULTADDSUM is
    generic(
        GRS_EN          : string  := "FALSE";
        SYNC_RST        : string  := "FALSE";
        SIB1_EN         : string  := "FALSE";
        SIB2_EN         : string  := "FALSE";
        SIB3_EN         : string  := "FALSE";
        INREG_EN        : string  := "FALSE";
        PIPEREG_EN      : string  := "FALSE";
        OUTREG_EN       : string  := "FALSE";
        ADDSUB_OP01     : integer := 1;
        ADDSUB_OP23     : integer := 1;
        ADDSUBSUM_OP    : integer := 1;
        SC_PSE_A0       : integer := 0;
        SC_PSE_A1       : integer := 0;
        SC_PSE_A2       : integer := 0;
        SC_PSE_A3       : integer := 0;
        SC_PSE_B0       : integer := 0;
        SC_PSE_B1       : integer := 0;
        SC_PSE_B2       : integer := 0;
        SC_PSE_B3       : integer := 0;
        DYN_OP_SEL0     : integer := 1;
        DYN_OP_SEL1     : integer := 1;
        DYN_OP_SEL2     : integer := 1;
        ASIZE           : integer := 9;
        BSIZE           : integer := 9;
        PSIZE           : vl_notype
    );
    port(
        CE              : in     vl_logic;
        RST             : in     vl_logic;
        CLK             : in     vl_logic;
        A_SIGNED01      : in     vl_logic;
        A_SIGNED23      : in     vl_logic;
        A0              : in     vl_logic_vector;
        A1              : in     vl_logic_vector;
        A2              : in     vl_logic_vector;
        A3              : in     vl_logic_vector;
        B_SIGNED01      : in     vl_logic;
        B_SIGNED23      : in     vl_logic;
        B0              : in     vl_logic_vector;
        B1              : in     vl_logic_vector;
        B2              : in     vl_logic_vector;
        B3              : in     vl_logic_vector;
        ADDSUB01        : in     vl_logic;
        ADDSUB23        : in     vl_logic;
        ADDSUBSUM       : in     vl_logic;
        P               : out    vl_logic_vector
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of GRS_EN : constant is 1;
    attribute mti_svvh_generic_type of SYNC_RST : constant is 1;
    attribute mti_svvh_generic_type of SIB1_EN : constant is 1;
    attribute mti_svvh_generic_type of SIB2_EN : constant is 1;
    attribute mti_svvh_generic_type of SIB3_EN : constant is 1;
    attribute mti_svvh_generic_type of INREG_EN : constant is 1;
    attribute mti_svvh_generic_type of PIPEREG_EN : constant is 1;
    attribute mti_svvh_generic_type of OUTREG_EN : constant is 1;
    attribute mti_svvh_generic_type of ADDSUB_OP01 : constant is 1;
    attribute mti_svvh_generic_type of ADDSUB_OP23 : constant is 1;
    attribute mti_svvh_generic_type of ADDSUBSUM_OP : constant is 1;
    attribute mti_svvh_generic_type of SC_PSE_A0 : constant is 1;
    attribute mti_svvh_generic_type of SC_PSE_A1 : constant is 1;
    attribute mti_svvh_generic_type of SC_PSE_A2 : constant is 1;
    attribute mti_svvh_generic_type of SC_PSE_A3 : constant is 1;
    attribute mti_svvh_generic_type of SC_PSE_B0 : constant is 1;
    attribute mti_svvh_generic_type of SC_PSE_B1 : constant is 1;
    attribute mti_svvh_generic_type of SC_PSE_B2 : constant is 1;
    attribute mti_svvh_generic_type of SC_PSE_B3 : constant is 1;
    attribute mti_svvh_generic_type of DYN_OP_SEL0 : constant is 1;
    attribute mti_svvh_generic_type of DYN_OP_SEL1 : constant is 1;
    attribute mti_svvh_generic_type of DYN_OP_SEL2 : constant is 1;
    attribute mti_svvh_generic_type of ASIZE : constant is 1;
    attribute mti_svvh_generic_type of BSIZE : constant is 1;
    attribute mti_svvh_generic_type of PSIZE : constant is 3;
end INT_MULTADDSUM;
