`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5EQunmjOIx9JmleHSlJGSC24ycyCtLGjXAPzKxQ24ZKNB74CVApJpDE1sw8XbNx5
btxTeMt9RoeXQdnGapzT9PYWNonKn2NvjtEn2ubBmZfbaCaavB7CC3iYhIPj2JL9
HWRQ5ClH3gBKqBnhqf8s0R9/j2ZKQRjhyx82mhhFHA/21lUkwOT3AhWQXrQW5iyT
oZx13dQSpBZpRNch7YJv1Z5t/IFKwQkVXOPYlTmndVWRbAHTEWb7Y3uGG1zRXr+I
ts8IlYMDiD1L2uYTQO4bEeux2vatDT5k6OEkbgQ8LKNnirRDo2qxg673mUGh88zb
Jy1Y/XVt8EmljX2zbrZQVP24BA7kjLn+Xgal1ALi3+HUso51DGPVFB2/BCI9et5B
tkikcGydhQbMqTSnrqYRyQbEFBqlr4K1EwQW1dYjv/2OKMHAPrDmKkBZQes/nDbm
dpbrSoTsOGfVONqHSEA1SjTz0W3vVadT3hl/1wf8iLWGY45Dj47BK1PO5JIOOO3P
tGYt5jQ2o5ZI7+11om0iULzwQ9MULfpPVaQ/5K98SA1uQOP/l/EeU+8SKjdOXr84
PIhFWJlBc4n4dmDKSdpgv4Mc2nJI3bnQHE9Xc4D830gRSSAlRIgXNTRY1gz27ixi
PiXz3/ugQF2vWu0ugbFL5AaPs54Y19lojWW/slb8u/bE+DMcKt0WW9QZ3HQ+DTdC
VTV/LwxOM48W7PjnnkhJjzVSpS2TT+FyyjzkHCpirM5mlPNF6+POO3RPGCIsotUr
wdBywj7B45za9pQAyTAaaVw9O7F3vQyhVLTYpygociY=
`protect END_PROTECTED
