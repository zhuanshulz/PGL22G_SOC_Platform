`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JIYjYGENysHgYlJXLHIrZ8VCn+3Gt6gCIfsUG29A1WwucpgWO4u3nyjitZmd2UpF
0K2Ms5wkDHNWZk8yYncBnC+AgcLed4W0Xq+eZgcCCvR+akAgWW5c7xl2GNc3OI46
Cf7PpsEqH5MWtYI6adeO4NhHv65bVL8MIimuxRJv5EGIrE4QL8a5c0Muv+YCy/oF
MOVqkMAND0UXG8t855/j1BwZNDp/hNXmoiHd32uBfuMdxJLVRGZWvWsbIv7UV7LU
Z9GAcCKeN0GBi0MpifG0SNKb+527+au1zG5S0Qt/QqSu/iiWFrbaPVGqdYMA/aay
NNt5z0Bo8BvsOcnPPDfhoYr3TMS9cp1wX8gj+hbUxj2M4w/6Ck8cboPeGmgo49e9
noEd16Ye5y4/i3GRUoGnBsz2EdKtoKiq1Ky8ERyq31iBQ8kzaf2NjyFRjgrLJTLx
88HtxKZfBhUpCFPhTHMItW+CGCFpxpQjGH4A7IkNr0/dZyBw+huSuOj7QelnK1hq
jWxLmFMfFCFC1S283ihg+mUtK94sfwGQKHjHp6I8Yu4NOBVZm/VvUY4ulAOm7sSK
q/tJMMB4zsLniXVQQxiCMy8/O1hWu3XHqJ427EMPW3v5SHHe1WWtOqhAicItCP9m
DlxW8oyYxTUjRzlF3NihWj+yboP+N/CLOylVTw7Hb18El7vTfc+ILVGzN7YDhB0M
I1h+nzRIDgEkD7k5lCARHcWYH5lNiMAHfJiwQ865yhUoxg4TEU+FYr2aNPEvv6wz
ncDsBh4pVT1fvXiDBRBofKqK9506Z9NhyrJT4tnR1Pj4P7EOvMcbhOb8AlXxpTMp
SWqROU3YlVJhLB2mjDVSrLnKQsPM340Gr9F1SYmHa2M=
`protect END_PROTECTED
