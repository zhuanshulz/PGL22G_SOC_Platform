`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Lwu0vuzCmcZCup486L8IkBBWD1vLF9gbByvySBl4ZOypnBgpl77b5XtxCROPbEOD
FV+MMn5tOXv4T+sXRxR7aplckgQIe+p3Jy69l3ykXMLx8W6B0pFiYdiuu72fEbRg
vMWmcXMItplFJeZfr71c/7d/I8DKDegHNpR25qGstMrdGBYqKYBS/R2GNamk+2rr
r2ciolHYzQBBeMnByqsRkd/E+2fWIVWDlfZiLv+koGAyXm2L1m4wAO2BVEdLUKHN
s1ONGHWDr3ISOv/LNCKG/rpPRW7VybdX39waai6owO3wfnkE1TQdBv0xmH3z9Z74
jZLF+feuYpvOxKS2AFbKOLbXPOTOmVJEhNvSehY/lFjPDr1RQy5L/2C/cyWcwE3x
CPh4hO1HZMgrDGjyUVfLVgq0HGiQtzt6LfVIcd+kZ6MPRzw9HqO6h1QLZpFyBXPJ
Ztp1cU+YrN0BDvjAbUjsXk/n/2Qf46K0E0T5QSbjd9Ox4ge4O7boLrwtZ6jqihx4
m4fiwMl3ZcMXTZI6xJ63dYdjZuSZvT2uUhmad3VrJwYmIxUMfhGZVhJOvj5vhYt+
+zMrqHqhTnOQJ+GyuvlH3N1y5u9QhQSOfSWR8P5Q0sQR0gIscHD+t0YqH7yXADvS
IuYA4FuULwFwqH0SZV4A5SOINr0Aun4603aLs0nzFKtGeEYY+kkImGzAbaHGexCJ
0ipwGJ4YQA2+fEI0G0mhdLJt4U2nFFTn3dQ066SX46fQjgPWoHZWrpPiGUv02Xg7
Cyg95bS+8hbFjBLDzk5+rA==
`protect END_PROTECTED
