`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rJAeDTK//FopzC1z83K70vbETBWXyQKSUTGsfkskdNNQ2yBuH8lJAYECLZvcZK1a
fuxi7Gl2ABGVCK/5BPB53V0K+fB4ZrK/jFVtoy2M2Gx3qDme3HmG2ydmLr1VMwuI
lOaze00G8h6MkdBSxDFo8ls5PZkzc/se+tFRd3lyVzCCigmWRHitlzUnw0rlzvc/
+ax2jisgyGQ9bEKLltf9JR/uh9SLmHPAbNXMHjh3ExjzY1EreUpZ07jK7gmRvfQ3
S6rXFesnl9R/qqrhqB+CCIyZ7XjsLN5E7JwiLQgOONQz+rVI0/DePsPdZMG38l5C
JSiGDHm74OZ3vWTYOKk4MIt8Y4z/VJWy/Jb+SCks3jjvd8fnGDdT5356jLoxZSIl
rjtQZKUgT3klM3PqIiXQbl4xVSIL7eC/KhuuKpCBEynwHGHX4KvVAr2BLh8RdhkY
3VUtUeRXTgGxxCEsmDqDLrmOgdqMI7vVzgleAJfDLiYdL4MN2bjizJSkfD1L0P5U
6Y2KZvzssmtG2aN7hi+wcHIP8MIwzV5uj0XtUFg17aWgeezru3cqiq4FzZOgGxC2
/FIAFsCqvhAzYQCoimX/b+26QltnhxjCBSFlGvihnto7rkFVF6VceHdii+hL4HSB
CCB4c6Nfu+gPMVo5RX5VG0OW+fWgloLxVinVZJHgGH6/2c1m0gaZmOLHLwgeJPQD
DacmQIsizG78u9yW53hbL63/1TAqCnvHX6QUNaGX0B/a6ss75SX/EFjPgTuzortE
Pdxh9qKSBv10dloYuKXLHgN1Y6XH62G9mpXyqLPZeKUndK2Vo7ZfkMsLGUQ6zptv
Le0lo6HOg75dIveLFLb3UK6qnxVT5HcAIpplWfa9EB+XKslxiauFO1beXbxoVs4s
RPwDAChto/klYAoM+Jy3RIR1bsLeRQwoJhgegNRH+PdpGY9hsBT3zJckuxXsuLmG
4Le8kCSUw2ZUcizivrAguu7Gwd8KODNoE9I2GFfvB3UZ5/xhkiMe2hsgx9yK0PdG
t3eaE2knlsJjMm85YneYi7kzhInmZ/fEX2LPXzLoz0U=
`protect END_PROTECTED
