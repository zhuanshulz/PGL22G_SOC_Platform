`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1CKfGbQH+AydkaYx3mOH9HWPpYnql5WeSSSl+YursQhkceXONHnWsSc38DFzKXv7
0sXtDo3E5rWVUCNVgaBXwzersJsHFRZeQ2gyXzSfnKyJetKpuaHYfCjuSy0e++Ge
T5ER8rW8a2rnujyQ5u2CRLlX3UX/TTMCSj6yOnIVFTdfziJHIVLlK4qOG8lRWT2P
jrdj+V+8AY7krqCQ7oC1RUe1sYKQW99UtxIjwY2mH4U1ILX8te3+pL+9JhGS0+my
IpymXehSIO5agNH/oPFIcRXioQNC13h+U6QW6JyL1Qf0HC+wevKmN02x5axr7Fdm
9FPq87i5UW7rz8BZxtiFox7bSMvJ8W/9dA6kPl8spSE08ctdYJDHP93uYz6afPfn
98rXuTouEOiclr+aP2WD/0+YlzIMst5t4vp+XoRYKHqK/QIi2woguXD/5f74ohjH
ftlHWav5ZPYOpIgvWGyU7nXEywubK34Y8cIM4eklN0FwVUvMLxbzsi4P0yTcnCVi
1PCc9eTjvJUGgttPvl4ALqdeu6oB0FPlgjGiHxplwnBOn9olEEYlOa5ESSsGJ/pL
1Nshg1QZKkqNxe1Y2TJRb2n9GfvOLLtruWfgMSkurSAF1Eq2ZRHkZAgsKc78cywx
8VpMm2VJfn7T9CPsbqhz5WTgF63ee0FNmc6bH83DnYZuWo320/nkujfLPl5CFu0j
A6Ke61nHQtdfAU+PCHNdRxNUUKIdZVmqhk4bk8mVEETaWTdbTSHrUuRsppD2eAJL
UyoeCbEaTqGstbAtqCAVP6wV0ZcEGSiCfvmPyqYfrK6eO4SeLY5H4HPvAkbCc4uU
kjFzgd2dzE3VCXWi2lUP4oZQLkyV3sKj9Xug8KjkYNJ0SP3hdsdc31oLdxb9x8kC
7KI+bweu9R3XTalK/hryRtvWiV49lA1F4fistWElqrQXVyrMm35s3biwfhLF00zz
dJsVAWoM/plFto0FjRwD1e+AP4HhuMhcru5WclK2TmD6DsyAhFLC0P6ZcQ3MjD7V
OAotNPCMaUtF/ZX84RtaO8UkXt0XCN49GdoaBpfa5vA8uE0O5sXBgd7Ycnaai1IO
cWgMFaRIt0VK/8PivsZnZsu8jG4WqJ/+h3Z5JFItqXZlNtrPjvb7E6O18oHNQNWT
S2PaiBIVm6U1HUO7yD+X27cJc+Wy0+bDUSwYHS1tfslGKYhZNF8T9u+TwoZdVF8n
Xbw2eaugJ2Iz7kQQ3awEdhU2Rb5GCzyKdOuoStJu5uYkXm1A4y+H1QwLCkHOexH/
8vLoVJZ42SNeTe2Ft0cGlZ7Tgq+7x/FJgMj+O3MXe9Fes5oP0ISKal+7rad6a7YH
ozL+ohVWPo5oO1wxfkA1HZf+N4Rdhk8WO/I+kTaIZ8Q24t/xBcfccqcM2zUvex9s
Z9BtQmnay/Csdx1qB61szORmlpOOhg+ENPgrSfZitTq6FXtY9rbn7Z/hozs5YRJb
uEfYqqXDf5H/Tpk1M1aiiPNLFbslneo4EHbPxHqDbldaLxJccukWCKg9kgImBnCB
NaXU1ZY6xxWaTaFi7kMgdd2SCBRx6vVEPzosTlk4lwagTPzRG5op4oI2S1AgKA+K
i7vFmKZxIZPjLG1q9szzbFYoOdhG1cMjZVxEnfeMXcU3HiD8FwpXv7dskWSAkxgw
AuZz9OmIwFcbdps+Lhn0c5YFKjIpI3hy0amXJLQkylH3MVc7phIndMRaL0Y4stoV
7YJhven+eX5xNvRBSmCKinBu0sYm1rZknLwYy/lLdJM7HR7A64+uyTYJTjGykJWk
v6iQxbPDkTHrodtiR6JEFkWK5dAVTADRp9CTrx9XPY1p7pzsna/rsBa9H5lUOQG4
B81BHBty2ucCiqxioqmm4w+79VQZ6Z/TsZ5Kbzrqawg/t3D2tsINfFnOcsAoHwzP
jGJMIB81g8U61OJgDw98bzKSYlOizI2q8o18htx3cOpHG7h66VpPvceYH9om5DGk
mbyMj3OqUUvQAYF/l9h+dg+IH2Ide3KwM1vjr09LLi2y4ougmTeKCKCSPRVx24jd
kTD2zgHjUtXRNe6NZv0+p/lkKLWWVCBdxsa+lGLVdMxFFhRa8FsLfxsS8Lq9xBDf
YBZOTbpqdAzDDcmx5nAkoT+QeRuDFg47PFCYZCU9joNMXIKEDMFYC+j8zJ83I4xk
mfGWM5mudhY8VZIsXw61J2q4Mx3mWLOkK+FzmKbMDcb0pcCWjiQ74aphNpJZAEyN
AfAdduuEjxycH8ONq5jfvsW1khIozzLkQQpPsN2Cq84yegrHGRyj2Cnkl/KULPvS
gtAeXmC9hRLE9rUzy+TstJXAQBioH4+p4LPqvSD6sLEMOTGxEu00YHo3C5waNUJ/
g0XxXHcVbN66ZbZxuNZWbCWeuwHDeawn6GOUT6Sd35k9BEdh5iBVZ2fxaivuUoiu
KGnmd7UkhP/n/zWki0wL1FiQGy+3QX8ANToZ5/lxQmrNYeJ+NPSW5V4RpoVes36N
v1+rDOhW8ovdUvpks+8exODRaY2DN7q8cuqQI5EcYCGSd37NLVa1vlSBKCPVkggh
wkOdr7jMsm49EoVj/vO/PVxrBUzqWQh31IhfyAa57lC+RZODwVALyGBwO0gT6I/i
NTkdopeQxpwvwyBjXeZh8loesSF+S1/sKoHyJOR7mVJe+YXKNfFfPkZH9M3TOkJD
ouuAe/dCK8ZVh6oo3+Q7ThRWJEEtcAn80cWCWudq00P6jv1O7zDJvR+MeSKiJtRc
NABs//h/kpwR3rbn3ag15F1RtkrX82EWpLhW08QVeBZEYiQuL5z/sPFmFGTAsVvk
oZx7jPXvPINNB7vQRQ6wecwPk05BVxMcqAoa6NbF2QGh8TVronh6aA5gWa5zKo2s
4A3+jBZpjRoTFTJCZ93I3YACobL75iILy0+VFNioqy9NjBY4Y+LhkUhEGi1LWIaS
51hEi+TxLcf233MRu8C7O2v6fWm52qG+MByQMwIh0Di1IKH4y2PRvrPxl3l2GFq9
RIHE6QlRWl99T9KpN4b0n1Jn5wlEOsbBApuvpXaIBKko4/vqHxjI0EK/6M1erS/z
TLVHpeWzY0Pu+YLP15/OyiXqByxvjW+cHWQkMi/dVaVsLhZ6oggWNGAqoPC/FuNr
0s+Kkbni+TFf/D5cePuIfd6uCGsd+IIyKjXhooUiFunX6KonYOYIc1gbuehR6x9H
mS0STMUrgjsCglJ8RYVh4MhL/iJ4wDOY5NWr5KCDp/u46T2pB7ix3cFKavMk6hdf
C9G9h1LrTmAx6aSqErhlJqSrpQ+lyupd/XP2pff3j1XNrJxVvH+jr8zy3MMwcVBu
V3GRslZXdlJ/Z7hkGpdS+1UP4BBHjitZRwLpn8p2U6PRZgq+aFBauSODXPTLDjiw
f1Hg2eWWDXMwbSTv6MLPe0V0WCDhuORVQL7Igp7cDVBW4lDNvRay40jFbrfHwFDh
EHnse+YwQLJtDn8UdFrancuyL01Mzl0WKhIvMKbXjtVHPqtTazles3VtS6Jisb/+
BAmKsFVmM6X/mJUPZj9CGtlABFHDQxs9mcJFu9AQcI0QnwBZNzjWF13xLHUaDbN+
dfhIfBYuS7NgNAvVd+WbrydxZUDkLGx6BgtEToKUr7kEbss+vkl7r2K4n19J74Yg
xHIo/8YoLk6YkjxuDFbHPy8KAC6H1ltmzjzxjB/bsh4+nGVIxX0Hugmo5Tb5GeBj
qr6/RtF2TU0tHmiofSkEX9Ta4w8mEAIFzUgsDHYTjcRRkR1xcpTppoeffBK3cQeo
c88gpzuy7qUkUvXoCEj1y8w+nTpmfdBBOcCGmt2z83OPuZHa4mr8Y7UeZuIgroRM
7S7M5nDRjTxFlInytELX5s/cQRKlRZ3HxqW4nC5xmQsiGcTGVAppC7NxaYiqr6c3
l8gAHK7ZUArtq1X8CqOV2zra5+Z4rHvHvxE39GFEeFrZ6BQqN21F2QZ1NSH1nl0T
o4rTAEmmQ3v4hDzV9lzU5TpuLljDyiJFmf3smwWhSMRxfYtjYVTtxZDJaie3nlKV
d2N//r5FUPC9KPeAKbeWHfMgWS4ehbGg8F0Tus+1hpgV6tFnJzZNlrG7PUhi23MI
CILkyGJBLaFCfFR8W/S7rVEfKIa9SAAKbXnVQrVHsbbbhvuRSX7dYSPnY6cOO9hf
U5eyqqZrwFDOL22ZFZNutU3IbexK77qAVNUBMCR16O8A4IbTaAPWDICjkHfyXC9W
AFLQPKZJv4SV3AP2OtXqvOhWm76ESvJBp47O7NitYryCBn+67qUr3uZSp1X7YhX6
fy9rJtPSxUMOVxUW8fZ3RR+Ohlsdle7lfYFHAVETovaLJtZRLFrkRNneirDZoEpa
SxKjg4AbWYsIDHs6g+j2aA//ESs7Za2RRfyk4YLOy3EvhJOZij6AdbehNVZb2ph8
xgns3Cm9lPFRSvBfH6xHYZCHPtajQ9ye3vDD6EloOfFn4WFtHrW5gk/oLSIARi6f
EBU+5S3/ypSo2ikScc20e5x6LHB2DkIHmslhfX0XFhjb93Zk9A60CAqL243O4YM9
NllbLntUqjVJ/M5H59g/dJHIaiHED6kiFkdG5xn21XTKiTTipoYKy7JFiNprNhrE
FkthCZboyh9lJAlyrSBjch3BlIhZWVvUhzYSRM3vBTvQnSS6yNCn6p+ygojitoAn
XQdCAxXFf+MkL8HBetfkIaK7aFbJJN14KbCgS9O2IiZfbin4wMaj7PrKpV6JzChp
FQNGj5WKxouYbl+g9m7Y6YQtkJPLhPSIH5VnSFGlB0cR6i7ssF5YA44hEMdws7ky
1Ylisacqj10Puxbe7KUJt8Xbai3OO86VLx9Hn+4OY7hZChj0x/ths7g6tf6iRdLi
zgBaLY2KuLOTgRRWdAZUl7Rf2f5C8+XcZ6I1RoI2aR/lQPqnYAdj2SJe2YT7QDJ8
qP3NAlJkO/j6+S78GGjmU9kRG8jQZ+gQMyELtGFNbOUOkONKjoSpZv3fBPUuCte2
Jz6fRchzNMZQFM1vX02GH0OMlA64UwctnrojTnmiJbTQ8RhICh29WLrOh4Mh1+th
jJUwEwLGGt3Zm6+J18SbHnd35k4eEXX6kvFbq0uMXkToa0abr3BsJC252xAhQwAX
S7gIBEVkjOQk6gwmwL8iin8joOMNYl0RwpmDIQpcDKdPxRGidq33xYjB11lXVWgG
71V1k/BXdH6/aKVm/O5Oq6qy/Y5FcN6yexeCqQmszfOJbasWybPKpdgU+k82J3N9
ZpWdE+kgeEwp9CXzG6A4b0urXTsz7BE4xweANNcdphL6W0UeKhtyQTUGe/QNR+lz
pNb1ES5jmB1xC04X9QZu+Kx+5hrtWR6sSQWg17eD1rEyyQprqsMFPuSRorXtnebx
z2KQ3bol0bXpOUDq1Cs8/F4hHWqC5PwQr4WgXbu0URIigA/lGiKrpMhf9w1D3LTY
xZv2v01iKIZj9lFxjSH9bC+9xBoRH6r8PsS0T9cQ0I0adnQ4DVCOPeSRmbNQPfzX
h7EmIt2Fa91fQasffOB4Aehg4sZoElJ9Iz8XMTXeH4Coftf7CL9yiV4FnFjZMKbx
ce6AdvU+EVTrvbbZ+XXc9xHuKc82WW3zShudykqolOG94MzYSagcMjmGErHWybzB
Brxj+XOQbJOT+jdj1jneJGsAPv88kQPRC3EvrfGkL7jRIKo39vyyrYAnxLWeTXy2
Ic7dTyBmZRBuK6LJd26lOm/Xn32rVLp1F7HNdzv+LbMVyJvnXh2DgjP1iq+IgrvL
JqMuOHAM/3oGMadlx4DQXA0oIfoxorpYsiJr7kS0un6NjuJenta9jObOmALNMaOm
g2U9POcK44vU91vX5U6b1qUCI5xwrbFENiI1YsFeHereh8H0rTVh3kxwpSdONCxk
yFppBxhFZh2yU65TgGNXR5VNkOCgd2imkENHxJoO7HEg1umeVl+8kPWNUD1mqoyJ
wn2lw3q4EbIR3pkTqJ5N4cd2BOq//bg/wtxF8Tty8JRvUML1vj9gSUdgmm0RLQDg
46d77MnrlrptlTbNURk2SVXpOikNGnHWLLwhfmuvDlpAwqAiuNQpPGMg+MDGeni3
ckHa5LNZeQQhu4zSR3w1Zl3cu5e/j8nxxUHB9ulWid/ju5KMKJQcoR3+Wl9ng9fS
a512bf49CVIIH6mAFUXb39d0jwiH6Sym7phsqBktvHv615VbdwuzRTOsBUl0tbTd
ehkhBqFXHXkXbtx+OZYbLroHOWuxBCzlJOiaYaQrG7hTLzx4fWaGkBOZ9ma/RdLA
zg1wnMl5yXF7wn7L3ZMuJq353ExkpVaQiHz1dtBduo0kDinJKCB0c59BOcIP2sI8
OyM3LBFoIYChvJNtwaKh0j3D8KMMdnN3Op6WAWR22DW569YORM6I5uFibwLQ20Ab
/PYX5ZG3nL5BD/jHLEtirEbgYkhYk8RLdzD1gB2kNnAivk/t9sIo7ypWu4cbGJHE
GIoMHcowMTaMnH6Kr3vZxFQiIEinQrf8cA272wMUBKJ+KgBobVsf2Y/vGglYZt/Q
1w2F/F3pcsxb47NO79ejRCvZIWU8qcOY9k++EzoRXAr6jPzhMEA6nTqk9nVvmhD9
bC8tEx5+NoOEZp+JkGK6IQ+5fF7LFMKEb4MzZTDAxhWmIgTajStZxsrJbsGV59gQ
ZCkFjkEilBniixwfiLS3K4sAg9C6wJ9bl27kZvBEZNsQ55FJGYwEVOBZZkCasHnG
psc+1PPeAc3BCyaysm6EY+SZVOEEU6YGvrKqZ0N0vz4KoBFuSpdp/uwjlxLfgL4d
nSZgVHTc3w0k0WUizjY608fvbBWaFk4j3EVlDVuaIw2FmICfAMYMUKeWMkC3rSz8
5eGzFbcIXA+73hWX3ulNAfFEPsH0gWMcdsU/TJrAMrGQaUnKi+xx+4kiHndRsHsD
31KPcYfZmrzxi4FN3Qxm0gtvdoR2Kr5sQJtVBdBKMSmjDr1b2mItNOpJVFhNe1T7
oC7hME6ZwLLCy7lN90vn/4bRRUfqDSj17JIVC6C07YF8URbZ7Gicm6PCab1fcRAc
mM4sa2YDfNyCxXlMgP2eh3To/HVJ3NaGfGQOphMIv1JWEq2WmRDy7esT6iIGOX8m
j/pvxW+kDBc7qdhMTvpRhP9suB8YJEOyOvaiSf0B0+l0vLvgER5HWvCKTVmecNzQ
8eSOenSsmmbElzfv71aphcdQRfgJirzA7iGGV3CMD0ALzttcN2soIv2ajXAy+lA5
JTbJH4MWiOj0U1tGFwVer1X+juqbSOtXvjauNliTcvYNNd4/05mRVjLzYiWUAxns
e6t1NcwNKRpjEmN/wpwSh8j5kWi8Gf1bwB8cm6Mo2+LW6WWOGXyRRKjNfnN8Aduc
LFGsalJyWWB/cJf2GYunnpFiCOlmAP355+pkO5ctluM7tcSagBIxwQACciXdeS+V
swSHSHPaVpXJ5j17N8eaH+H1LVSmZXsejoyJDik6JgUerNq2QKIDiCZfaHE4O8A/
KJPlH2+jfG9b53QEkUKtFzF2x3JYjH6x/B8o2m2SxSxku1+ERRrKvFqY2YLnxXW0
eNk4kK5dUBVWdqv0HNXjSNEZTjKqEvOFkPZv0fRz5p8d7Y91B9oZT12WDs2/qE/4
tTwqAZugcSTiPn5rSLxJsa/yghltzf4CMDxuwvuc0yfnLbq86ABrsKXMZ8aA9nTO
zlo8tFHGpAAdhVqz9V0ZjX5h0eF78JefoDFx9WcDCwE2MKZciwfaKfymP7zO2LF+
efN7pDLizp+B0y4xY70UVJLUQ15JkZbxNhLczBFQ141igDrf3PghpzjhDm+3885u
aY7BSfRvmIO3U+f8Li6mAPvC1zg9LSa6PXqiK+0LW/iWJ55xNzYcIp3W+U2of1fh
14Zs/x4D6A8Vqnfvt0NmloLbgdJY9QSiHBpBfsIs+ivUeAk0GPhFf5NQGQlXsehr
H95Woi4CUP1j6yZm5mo0A/LCc2SRBu2MeSlkAleXVip2k3ILZ7E4O4lHCyJwU6mF
jRO8s5M2JozvZwAhCshztbOI69Cq6/H19+BTfwei16SmWK8ve9v9RxSn83Wikwdk
zRL3CJDqeM+k9qRLw9oajwK+gYQr/zmbOaQawfcFIo58kkgbsJ9bf8EHKluziVH1
JjM8rKQaDLkS1YJ3d3AWouD61gkeFBvh3T5HSIlS1g7BqdbxD5hL8EyJh5WG6VAu
ltz0RzG5Z33bPGaQrsdImi5RRGpBYRHaN5Vfe0FOHo2CxZWg5CWKVMJFsxvPQy85
p60hvH0SoRxvWgqmk6S45j0fnSSh50oO3VGRvggtk5bKuCTP7/5mxg7bSAVPbj9b
fu59WLCKU+8qagZzKN65EgHJi8SGNnuyzu6ExNrOjfD37fh0tLoSHXe+wZJbz1ja
CRWcYbtKkk4cm4fU1kouwIbmgz3X4QbVIGtnv4SojVrAKK/n2lh+hLMGXFYlMRlG
3Tj7m89HY8MzFckp7gsNWSnvd6GUpcHGAMvfbLWmwMNPdBzCj7sJo0CnKIRagn3w
5zcNjrzDoz47f/nBFF/zrY1skd5nIhF4ldw+6nfO8WLSX48wnRkY0b9tEUcVHrjn
YYKIJEGl4AVy1OZQThBGldwlnPZd3j39rVwM//bcCK6JXLgHwVomDY5bxhKYHiXD
7Aqr64xzvHn7tMZgvAkj6on1ckyPo8TR3sHgj7JeQmNH2RcCY8UZkwn5218kbLCm
lZlNi4emF4OzyWXRTuKHOqy3PyezgUnjhdCSM7HeYYlkh7trjrZ5s6l0BNIREmC9
UpaBCnpNBUvHwwFyhQoFtBbstl2Qj7po8tcmE7ev0gfh9MdCaJP7jn+YqrmqcfS7
P9NVPCMJtw/lQHIxLp2Gil3uaO7nAYgjBCacXvu1ip09OLC1WQex8c6SS5NGGJ6e
KiUOgiw8einFgRcGgkbzZpdExkEL/uP9WPiBgbWPt8Fub54+zQXu/1z+xawEsqYp
IEUjSzyczUSNlE9K5s6jE42w5xVdRdfjmDPzpdVlkx+ucBTTbzODdJJ/RPajojTE
a+hP88yKb49gCf3DSq/z1RPFrqAQlvyz6OfLFiRgPlNSsvA7dSWYVjVruD7TvR2V
SoaVcegifh3xzfJr9+KzbPh/u5KNfpRSPzSSZTco85wVoAGGUde3hu6LM4NsD60q
VgveG3mqh06l41CnPOYa/GSoE0dSNWLXjOw5LeEVX10+92p5dtHo+0QdFlUrPGkM
3RoAjXHQh5zw2lSNVkN0Koj5LGQJsGSZkpQ0Cu2Al+WUh72oPyAuTG/yKmYjIbj6
OjOiONLahHK98SRNEXbIJtLmvjZcCE/R2nZ6jNWUT6dRWWDGrr4EvBPsL1j3/72p
zly0NZIdC6MxpELjVvziY87CaO9SsStw7y9iwKm7Ue6wfizFlCWAPcKep94qKPXx
b3NroCTwswU6SsFeWRWq64U2dsj+4EqbdOrh2P65VZFENSVfcylHDPcyJEHPu0mX
0WIgV8yXDa9yi6rriKaA/wfEM7QEVLH1q+GTZhL/E5+akCkf6lcWpPHAcpC1+IxJ
RQ3XQV/yw+UE+FP32/qkMNPgUYvuYWSc++7SIzX0kwE1YlzSV2LqSSASeoHZjXW9
FBq5btqIlVWtMoRTXP41TAHQXVOv0lvyhZ9EfyTyvMg0jlcVfSv87uLe8oYnEFKQ
LHR1+0HmgTaABxD+vaX6yRLjL0LBiaG5LVboHEsLssMB9cKhdodej5od9IHzGm9b
IEws8Fxws3uhuG4XH6iK3zxpoyWx4Kz+A9pTEz+wN1G05xV+ZKYHqlSO0ei73y9a
l68Bg6djoIKGkWnLUaNKQuw/gaesv5WMzheP6MxSnx33cOsf8I2k0lIJhFFwaAga
ER3Rq4IiNKDashO1Yku25aSmTkcipC2KV21QwvTj6gsFBgxop2ByM/PZsz4Fhj+r
TJcUoY0Dsep/GBWab1evab08VJfi7v2ws5rX8kXus4IL9ofdSnJ6UJFKXLLM8ais
pO5saxju+V4+0y4WTaOoH4u7fXIA0antqToW/lwpxnKdzqdvQQpZ7tlG3p5F8Ecu
oyfGB7eQxoF6yE1QS3TMiTA3udr4GSeTy3UjOilk8W0mOu+CvMOidzGyVdu5Lb+0
zhfw/96pcWc0pbJdCrexITVeDgqRH+YY/mV+3+oCY0IYEE7trWj9RtEAclpBgFHO
MDQO59wW3O3RMUx8Homem5ScvWijsKmp9F2mNZmdHajaIoGMy6zbrhgqkgA4xUFd
ZExzo2OWUBc88N6KWOCg1bG36ZLYs8lte5cRud6VUaG6SJAxqZaIEOUkPS00rcKf
S/8cDUjYi3X1sYupUhaW2SiMJSGx1iD9IvOOvqFNfz1m/Ez/jKm4ScoBQDWZFx91
Gr/rYONEx8PO6+mM9X/D1mPkebZqdEqHTgEBhF2kclSxFuVydCJLVwrMKgYHy1Xj
OffOlaEC0TpZPQWVKhMVs2ld5UBaabpuptGZ1NnI//7qZ6va6DykmG3d2k+h0axC
kV7JFcfakTz7xYfRCDURBY9Vpy9gH8nnPz8h8/ynDx3Hb+pwJIRy6hqvx7Z1VneC
zsWUg02Hgg+LzTsKr2MXQ7xD2ePdP4tpR4IHCZX4Bsad7U9Otvu4ffIifsjHugot
1YNb15F29w+oZSxwqiq/1kiBqGGmu7JM/BOqJ7sjA5sJWdz9nts0oahTnWFKaHEb
EYAJz7M8yHyegC95Z3F9TL96A0JlamYFsp8D1Zu7aTqQo/lWueCsjPT56DOYXA70
sV7BVhiG4weLCgGJQNgOT41taItm587XK44bNmPwVKLqfOduTrkpKJ3JcJqzT9Xc
4uWB9R5yOwBtZAX9P/Vb6pDEw7X+OYq+2s2fHU2xVA0JWr03W3ke0Wkm4XT+EMRI
Gvns91/d2n7Lm6mJFCNsur23/1MUsoqzCVXCUxP8i0y8RDwi6PWKfyc44+C87Fsf
5kc6ylpNpQdG7ABnaH9dKfrNS6//lo84KtKRbUgU+314yhIVZm8GfabeOsj4P7vr
5gxdr3Igkz+haSlwmYBH937qDY28kOrTmiBpFVlFDFEBMBGKw0guTXpSMtYiwtw5
GKc0ZYV6BdPe7xV/s9IqlA/JYHuRNA1eg3mz3sOqMBppWw+kQplNHanp+3TSNh/j
giJ7CgMWiIbMbONziQ5EE7Fj+EFVnln+c4z+9LIUbcXv+5JESQZtPudZF7nWVXxQ
VRfgdCcrrjxLBK8FiJDXwm54WQaZyte0D2sXOZ60P+vteQ+yIoEI2r8Jvbsf5IU3
fhnJwirT67n0y//f7mvjr4dp4FkgDH06ieU/zEN+zd2int5W+SzqMCxt5Ga8PcDy
qjxuyNBskpEQe1eU1Y9yNwwbx6pm8trA+OKq9JhvGw5F7qm1RQgtXoSjFvW4V6Kv
z2JC6yVXn8IJbh/J52ahEK0zDgcDNcViCmj8+1EDoUAGJgtg/94XLDPkVWRp24pw
BAoSUHmAJ59bZQp5KdOjJ/T426p1hvKT7MRwIH4SCatdsmYiLVU1rNrXsoUirH6m
d8aeIZFBrq1iT/NdUZvTXJulDx99CHujZQXrwjr3GV0SKSU57ScKfTCMg8roVg2t
GZ3uoILp/60eUm1E/hi+o6z50q3j3wcWOxBoOZ2hgZ7fwCRe4/9xPTcpuU12Ah2F
IoirtE45imuiS4FKj6bznCjdSFlubOPVcZz4vIY+ShzLB9UJiWo4oiMKVX5XDCa7
XdrNl+0Jt99xexVfQWFACZB2DsWctpjcPG8Amcl97Y2gTMiAXVBVwk9cZWmDL+S9
/dFC9O4a/4tiOBfKlTxE0UKw2rKwYBo6urM8d8C7tTsfw6o0uEa/LuQ03rkONi+b
CmszNDMYY+i2gFWKs5dl7lGmMYd8PH3rau8/62RD6uNPDzBMwKg4n2k0OMYYU3IM
UEn+JFb0838bJVAThTFWNwR/AUQShoroHItpbblSY9T/w87zwMKxcMx+1yJ5SpP0
D0LbhmQUhAytT4tfc/yZlOvoxM9HQFUONm/4VSCmxITiIS5OQz7W7kljsnH5e3AV
5YPQB46rn+OobyJCIIKonKsnB8ya9nA/daNb6bnqL7QLEPA83EqUaUg0/ZY/HgoO
MFMmR2sgjoHFR3HjDKuR9eAmkShv49lsVi+fDpi3OmEkIEPFrlqc8o4GIz1vB+eV
TdAOz8dXkJ3g0P+VjCfePQkyr4mGl/gmLRtR29LdyxjrIhS/8bwpqmqsXpvZa3FA
DX0EygAiC6gAUpkOCt0mhIKYlYSSYGJfmFMuB4ezcC+GbJs4FoAvish1J6PXMBrQ
khdQJOoHmd2I2TrhZBea7z/8a6MGcWdiTKPeO9cMk88GtSkbRZ8YBUfaq5L5azaE
DxycrnxT009BJ7N4AXksOYChRBROjICnl6vgD0H+iYfNa+glK72403hzy82/tJaw
rhc/RtwhQJ9FmQu73kuLT8/NEJ/+3/6Ihf0I31arocRdwcN1D9crkeRtgkbVvxUL
VWJ3l4+WHML3LDWKMlS50Q==
`protect END_PROTECTED
