`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YgL5HXgow7Fz4XjbG1NDJqPHSWoxHOelsuaRrhc0/AMPC7ExWnicdCYmUiG0dS5y
SbUQt/vK1VXhcZiolqkD+zv7+EvUlioPgub2a0QOU6jVSWB3asMxFKcI2go/bt/P
cPDhzBmGWQXWIyumV7kZoZn2nsJENXSM1Qe7H2kIqrVeX76WPKH0dkC7E52B4p1d
/nplDW21YtK/5BoGxB9Y0zVUVSCrv7RjaR+nXGAAA13VjNMzBbDsROVmr4AZ8Lrk
2cVBx6KqbzmkUn91MmZqHOHGFhGsJeNnMGoX9z2mvdXmYrsfzS02SDrW6uAepI7y
iysno8P+Sz6NVc1tOqkmv34pgtwuVT8ChzVV4JHSPK0drYv9DMiPO8wktH/t060m
OgHtEa+yCJRBtC1u7DXe+nrXWdmCj2QdK35mV8WlwBA+EL2Y+4JxcRUY4a5QvDFg
2d7cHSwAwGDHBfhAm+cZBg6a9Yyc4XLEmd7KbxfFkYJnFXJdGstKsTWHGhWFtPx+
XyoPYxZOJlR2pQ7Q0yRVeaNRTLuO9o93sdLU6GfRmvtcDqm7cjsoXElzDzU4M10l
7KMf127a6Lb1ok8+DQnRrhrOqGHsRJI0B8FmNal4S2YTGGx/A4Cq9OK5P4oMIbnS
4apb6Pyo92FKLSWVXnijvw9uVkjKhgPMiGMpsq216W/FX/000OWUN8R92UGabDn0
4VKErmxwiSTXODa+Gif/m2/lX22a5r3lZ9+zdjgXZIwaiFTGF2X0uQLo76H6KZCE
Z4r5vCmKHNzlhTbB81D9LsFV8e1gMPyAMkZ3P5vBMsVgvl4thZcGIZnq4imUtnWK
2jZSCudfBFXo1JSo8f4xm13LU5Wz9obmzDmWnu5uA85zunpL+oRNhJrwjxIFNluK
ru8Ue6nR5pOiQBJrUoGM+gZGVUjXcnwdzZhjC4CWRfklTpNueOG26iMdlArGL/LA
fCwfql521FMLzT/eW1DhVOMqKkKJTUMIIeEP/dU3Ti9LVaT6xmwKc3Yc1VectRuy
Cs5MruQoIv1FhtA2+8bIdRqDXFy3VmSTxoia4sDTXvdI1sVWVdjzo1hUbB1t/izZ
usgki29/6zpJGO3O0/+c0LSvtUuiaR1HqeL5mo3bF/fqcDoP++dTju8RGbBzPMLw
T1qeb+Q02mh0V4kaLCS/5XbcTlM5yP3MjNzMQKbNMf4GAs9kfmqGGqlwgdKzJKSf
hPmtxkOCPN+IB+PTQQy5HOtD+EITfcYEK72a1ngrZvki3A0rk5yrw5DCAtrmBnCO
U+hFJyDv4ONzgp/kFJdlV96hcvSAodm1mtGafTNHboAjqayup1N092rp07EApa6p
YPJ2KmduExAYvXLzDX+7iPxB/H9V4RoBYjwG1RSOlj8pqeZyx6aA07Ihcwvl++gD
BeV3h4jTPQqvjYKTBOC9ROxdS87lBmU6qsMQon2GqowJAXer9kLiTqUl6hxFzSfK
ORZ+9UTdWiY4lXksdMWfPjOKXUK9X/vy94qjJTfKqNwpr2vIn9jaRKLMwh8Y8PHf
p8bV3QIpR9CZD1kLQExTNfPlcWL4SAcqD1NTs9Kql+AxraHodyTfw1PQ3MM5odMp
Lbte3YV2KSxP76B9i1Fr5SnkSI013bvfwH/i/TiY7tJoMCVV0j8PuTe4VfqWt8Gl
rrurL6NNww57AqJcV6Nf38GuEfWKk0WGjSweRwytajl8h46Z4JfFoWD9+nFbzVMg
Vb1ol2tPj/DbZd4RBJwTNza3q4rGfdEoiBcU7exy1qQVX6AHNbMrhYfPqBPQTA//
0bfLF4sapd2CR07aOJPZJ0w/shWCgKxFFxOAgVgfW59DYrwunfZG/kba8TgqpEC5
6HU4LdTf5pxZfdKcOCCKYJeEe19cSVqtT6tbw+6TUty24dud9PTmOC2yeTxMhCiI
jvM5LT3DzfaT1XIDOGwgwUvsdH/pNqVfX+Z85daEjgml8mPPUlTDu7hLc+KNRBtI
HCTaPl4yLt5/6EGRVMY80cSpb030Wz+f0N5ABNO08WlFf4M/ucO/zIEG21G5S6od
n2X0fHo79NZEx1X4dAK/RVgktTigjNGKprvxMyYKJZj0GRjrMAbnEI5MOtMLE+jN
F9/8+OOlr2gRnvmqZSZdIaLutgp0aMX/4SOhPX5Kjp/yvvupcroLxXtTC7GK5kut
3X+MdPW1BNmLXk9mk/gxi/2Oc1FJtewZyxTNtq3c1Dv92KtklLl7M6YR5PW6/kx8
te4zB8XRfBo9gYU4qR2NLmUmrsBhAsxNWAuSlSA2j0C8NZbaEKAc32ScFwzihlr2
M31RebrP/uwQnahuhYNQw2szN5Nt6VYJBpR0If/4xN0zeVUVv5WJE0Dzf5NQ0y5U
t7nFulUisICLfqbVKtHU31s68ooViJKccLwARQaP0bokz2IW2NoAj/jSbcfqTMkp
LPirHoBlge5245IYVG52M6IcrK+5fFUBlnWl3jw79ft0ZEIcFBy7PgwVcwpVxxZP
pfqr5P7Cn8O3fQkeBefGfHoW1hC3vP9c76odtaNngpThvuQtM+9/HU7vcmX12ZXN
NsgZ+AHgRQ3id+tDQdprOObUS+vnenCntkW/Yoxoikue2+7kSM/J7jP6Uzd/503n
xlkpHbsd10BqA8z+7Y9bcvCzamiPlP0VEDGNc+iCgSRIg04+f95t0VVfOci5x8Qn
WZhvGNmhfpsK6/wzQ9xFZ7DXqIpl+QC3uio1H4ocyLjjafyu9HAqs/UjTslcE7Vq
I/yPsJYmqGBlyjXhRynRh0ZcxusVP9dNoSwtIbibpPGxEhQv8gc6vBdRpRJk2Pnb
MGBGOOWuGuVP62OBbok7k1B8sCztCVKHrXSq+MJwtEQriKgIud40WlhuE/cYvq+D
fpUKeEQvwQ5XByiGEgNz67Gtri/LR81ZTJtRO7t0X2aH2KUKX607ShWC9xcV/UsG
w0sywxBeBc3LXZwQSOvh4IlQIzmK0snFo5WNgB8tgeo1l3QNXslu8qAYXQlxZXG1
bpDct3in/EceMRQu2Bb0cF4Wj5NuZ/oo+dgP2DQ52n9u0gqQGOPdkhycNI6IKXdl
soHnPisQzhszyYVP8rRO6WoRphTyNr4LIBzlmyHUoGucVhAKgZc9KDCM7TZyCbAo
AuR/Mcfo09mT4lq2wT8cnl7jD654/kCHJVRKqF5vRcwkUxINqdgWinGNga+3BFPQ
10pYPk3g0o4Fh4cvxO6hpF3y68XuTL3CxYYWERSq3PW6a1wl/Na/FoWc2tomV260
hJMvWs4DYeLIBtBo5i1ONQLa5EZWFT2gUoGDbjO2UCRDoedPjQRPkKNQoSIOWhvC
X81NAn5i5U7cFOkUhGi6XoOw6JybAxySEKb6romOqcYQLNsrwy4BWWb0Dhs749aH
cjrHwUJkLtJ30zLRdMmi04+2oH8zgAPKTy3RCHX6YvsRA/MOS8EfhZCuVfyTajEW
fdbqBZz4KAEhTj/XY2uE23e3VFH3weDlQKAQkqLqOZ4DmzmbkIs2KeH7F68twWNl
9xBjUjkPPwXfG9SrQj6gz/mHNZEb0H9R9yWIpr0SAswMmqjmE6hCmTOpuhuQ9pSR
VoQ4hadWzXYAhYuSL6ibVOhVjrA02XfTUfeG8NG6Ziq2XLS9UMlkKDne5kA0gCTu
qMDy8eVH9rPo1zAoPXJC4lUIJNv7T77BWLjulvhMuTsihrl+EgJay1mu3CkXS8Qp
fb1RfNGH+1FxPJPp0WTNMCpoCOHZlpe9dce5nbQaDaW9g8b96h7zQHY0mOmJyA6Z
7tI5HQ6fU0rsHm64tXWD54nlI/95m2lgHDga8L27mmwV8yOqwLp7X8/KHALEsbjZ
FDN/Ntqzv3RNmp6yDZU2YXZtZv3ftavV3A076ErRStjOGlI1GUg2Yu3J4voFX4Gx
KFy746FJrwXpx1hgtebvuD/DjyHONd4AsyrkjQdTz/eF1VcPvpABduW4Sy92F+w/
MIyfd/VqXY1mcwme5wLl63Ov+I0tk7mYgFuoVU+/f66LQvmF3o8r8Ef0SNN2PwEZ
hAotV/7KBTjvxEhhhgo9cVeiGVpMAkot/Oasw9Upaa1pvq1oQc+i2+M1lyoPrb3M
lApKExfeCQMImozOnNL56MvnqMhKDFzPuAkw2uuQDffnEQWTHo6DyEgISFwnhQq8
Uv7NikUo+y/vbgMbLhpmYmWmDD9cFfVUxuaReY9cYLVCsT5HUgMcZIaXLjtHept7
hgxW4DQSOonJ4Wpca01F3L2oqHPgBXkhQTwXXDU463RF52RgYstvG0dLE5mIkb3/
rqTnldu28lJyN2jNHXXBjmJWXufEgODe/nAS+4AS8uaCGUPMYFIAKU6pLg+y1+Zm
FtuOwwmMitxs3NJ8uG6vmmDNgROa7bOTkVPLdONWyVZt7rQqMxT9M3tPVZfOitU1
29gAewFP7GbOb/SPgMl+Ka9S6e9eDOQw3D9bgSom3dU/9JWWQDRXb/9H1NqHLn48
JW/rrR15v6MeXXqzopjw4MYeKGG551xx1jP1e4DlxB+6XX1M1+vBkZ6qVXxpgabr
fmoqO+5sQCd01C1IMAI7BZqa7vmvlHXNkPsV/lDFv2aUf8ZL37tmNQz5E2wMJRfP
TUdV9OsNOoT3aV1JKgzRhBO1Ze3C7X3bNv3X+RNV5UpQE7UTMmVDODHBKFM482j1
K10smccv+HKFrtBsVs+KZMCfob+pvBd/SPKDCch5q8zIcSm5+n5Ms1lp61ffJ/91
DWFUxH/1MfOUooDVsH3PTi/2ktxkOKbcLgx3iQQE1stbeZH+iv42dqDJq/bqMo3e
ZKN3RUYVWNSne9rk8ya5IED49gMKe8OKcJk3I2qWZzo0IibQOkMf2fsDmJvARwPL
8v2G7FcxajcXnTuXWwDzjBHhvBBXudwSmb+ud4HvpXCJ2dpJy6vs/GHokllEei+u
eGk2UJR5G7/lOQ29/2t/UVN5A2tVWwCSIlJqw64ZGzV58xzFcoACM3t+W1oc+uiI
ImE43zG56azmqWG/ckbWeDeUFh5k5zbUwJCNxD7E2hVBSkb8ujKCI4bLZ1++X1d8
tlv7CWqHZURnB4Z9otTNJqLFOwjSXF6aQugP54pIM/0J7ZilUcGl63nwUb3ZKCgF
WJmN/2mGxAu6t/pcj75gjyLTyg6uuhQty/BtvV08NVo9i7uw5r+l4IjVzNB/nM/8
5l6Q+oiHQ7CQYJwEtnDy8JrCbSRsdb15CUq9DuBjcXY7O728lkXT86YPzEbOBAqo
SGsu9lb8f1d7QYxwKMaC7MRkdbHTHXJhGcw3H1ofg+SO365iYaXNfyaCYnwaKoNe
yb5k4p5msQv5nv/P6oWf31tkuyUe8kTv6RdiGaRPj9D8LbBQhd98QflVnYD3Ryqj
5nMH382SptHDig7jQQlOroo4rngCTZQOqNVq5mxbbnWI3YozN4n1ZhHfyHYYFkre
bKdTXwGYfZV9lE1a35QxnM7BvRTLqnlGm6x8d9nO3VClarmoAm+hHr+J/3w3nf+c
JlpwQCduFH3VkRSpt6+5MVnwM9oRIDfKOSZI6vd2zw6vnv397N0f75Ox5m5STQ5Z
BLi24INXi+sCrwmzqB7SHBHqKvyuI9g0qbpej6x08IwHXnNBkzXrBsstJYyWd4IR
ZEzuD9yMZFMgiImFTzMR66qXnMAXJA1Cf9Dbb/UuBKnYoyk20sVZZ5NT/1Pn6Fnl
HqSxTlRjmhT56CTgrEjR2q1aF+kMcMjwAI1wGO8p1IjMwju1SyepjF1pLJoAdXJg
9CMYL+kBZ2MmNJZUEavULDCB1RYNzFq3AXvkxT4kBOz4V28+N8DIP2N9hKPZaP70
sugylXADYHyKXE7fP08kWgMkmSsSwVZWpCcpRUoweg3j88E7C/xNak3zV9WAnRH5
zYn41FTvbpTqZDmU557w5D45zwL3aWXogo8T3JHRjUkmZHnPj4yMTrliKZdouwbw
cIVJyGWNBfHfD10S4a9lDv3d9ezURGKN/LIPT9SR8vSP4wB9hhQF6x43BoyJ91rn
QQFZikwROMeiDUTG9ROLfKCIHfmY1NJlFPjcxDp+IB5f1UXFJulQeyavPWRXQ4ou
tBArsIyKSRzro1gYn2EdaNI6j5ajdHihl8DPuNUTrdhm6gjGvfYpfX5Q4Gp7hlpM
PIbCboR4FjkiMSEfi+ZBVvJhyj4wDliHemQTI5ZU07ct24SOXoDjaSNU/UeNNdd6
bDzJX7aFvvy5VS4G0Yd4Z+GDRxlIjoGYbFjShSHRV7pxEVqz7xB/+eU9FN9jZCU/
5wC3rIAUZ7sw7Qru0bs5Nw8uam+eBUDIfJCMyE4qKUSajB6x0b8CU5u14TqXuXn8
IaW1HvPMZE7mBGUI1/QE9Omve0cal/FSYMfZaDTikYLtIET13q+T5hSxpGsjTxtt
MdMI9MWlzJ9SajkTveet5XLS6YpAKIJDmxMKC3notcDFQujfiH5WrU/aXcntEHDR
qSM58f6HV/FmGWBkVdODa+m2MPUpXPgqq5i8nbVhOodbhTIHCLvLfqxXWHOUDbbg
Kxqp+uva4tmi3LktfsjvCSZkuUjUj2klAGssQN/ljt2NYkz/ulND5GnXIOPyfr0D
VraUUQV8dbDsIPQKfKVQbH6cX8VvFsyP4b6kAbeBCQAm7RD0kgM+WUklN9W89HWu
nznqEWguKxF/YXmpHPSDfmj/b7rfa3uOb63KQ5s4hyfx+p8NcmorjuHb9VVrikZX
hTD6j7Hip0itT5IQqtfROqn5vwLwOZf3Va2XHVPOB+DSq9lEnBjJYN+a9taNHMeZ
6zSFIQW+6z1i+mJ5q/YMfQYSvvT67lJeW4T71fAcgJAGlkYRnrVK+wsgG9k2K8+i
siTSHMoOnBhLhcvE+lGxOUkwt4CmqAFZtrR3NBNxkcEk5fqwn3SmswllfNDAd/32
1d7zSsfSU8zTRpYG9Y/SnnlK/H6QL5Vv5MpfVsrxI/37gzslr0izHoEYd9j7/h7v
35zh4GBGh+Yo2r3rR9YNG9vaBU2+y/K6+gNpuZ08VkKh9C5cFXeDqxIJ2tVMKvR2
NFaSXlvacyMhnR/l4UgThYFf0e4XGIGWlicamnJ6QAYFeYCjqFSXW+tdoKGLoScy
UOld94+D3hdFlWpKSryJjCrGQ8nN9eab7z+ozZby7Xuoc7N/aNOMpXciF/F+Bdr3
vC4XuR/CjwXehHXIwOPIvd2F/Iu8D+R16e8WPPgDvxhvLBWygqzZG7SH5VPVGAuC
Kn1UvotqEhBRbp3W+MIxMnxvKQ+kDXGBCoIetpQzKkoThU3Qjg4COw9HBYb8AFGb
YXsnjioG2/bsXmDRriMkPiUtXjJJiUhdtlK7T0vRDEh1wQeWbbKx+QcyQVz1X1AO
OzgHv10acISpdGe3iGCO5a82nyJxp7nDHRUduYTK2u6qbcSlgn1EVMFdP5rix/Cl
wXheWI8jkZgZbUQY7jAt6XPKWylZIbCfCiw5LuiXZM1x+oyHloL3YHosfjZw/ku3
CrDalTlaFq2i+cD9Pb0Pqv3a5XnOfriVVxV1AZCYXPNglt+Aoru3rI9tmjMHXvHJ
mozh+B/6y0I9cOSnwQOqBQ4wFW0PCskaT+9DxPzDo77UB9XSZDKCcL08LY7BD+mU
2Xg3E0/AlIry8Om47wi5og==
`protect END_PROTECTED
