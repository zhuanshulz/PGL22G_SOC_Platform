`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jyVU6uK78uEII6bMHczTT7lkcYgK+RFiinqV+5NJpEUIR5RUD7by+NyvbRoaE9TC
I4Nf9w15itjztUXWSJ8QIL6S5RUCjbs8mN56GGnqiorKtRPCqp+15g+CePRgfsKo
TAGAxLm7x/96UZl0e4Cpdz+mpq9wNspA4uXwE3WuUx+ps3FIbPfhq/NvlLYZAQ9T
dQ0+H4jNW0SuUpeLqzrEhO6YN9fW+LEGt6bqIZoXoJkuXgOdPfRUTzpuGoQupXm8
hKg+kyZEq6J0ED69VfgccYiqhBBhKS3ZvmClEKE63/xj3tO4kpUS/8vzpvjiNM8P
yD4V1kqwWdOlj/ooDbI0v87PtrjTJBBvgQ2QSF/eqLaah6kaqHJyPOgpYrMaibSc
56SWIpdNn3agYfNpzQGgPTFqKjPwMaluur5e6/EW12m/tBsU6c/k10jIFxmGX7Na
W4SPKntVgjAbydGSxdf2/v0RCGbK3WMgYC0p7LFp4BcB5znsu/L3Fx5iX2w0CKon
`protect END_PROTECTED
