`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ASr3msLv+CuF7fubUqu3Hz0/r4HRtwzMEfsA3qtQIsSKe0j2vF9OErlvG5x+oDff
xuF67WOxvM+dIMV6RDptSpvz0rTngulIQGyl3E5YI1oqReMpp5hu1wYOw+6D+Fsj
Igxt6wznuSb0LFNjEqB4jrECS7BQPMbHaVR3FV5exwseCt5SawXTUeEbdB0oqBxZ
TSmVMG7NxiWjTVLFoTAX2OiTPY+POjcgu5kI0HcPwXjdxkygCtc9TMsN+3HFrSl1
hPNvcTYyoQakeTG87te0BeZi1ZLfucp/RQ/w6JfEwv05okD4sYbthf3LtEWwFVlM
GU8BseG7DqrxM0P4hCSNr2Sl3sQOFAP0/ZP5+Nkkj4kUiHPzHX4GW1BiipB/hL5p
cMccSgHmTZiAKJ+quwjnDBUc7W5HuZJ0Ym4k5JSihOwSZtv+YD3QtIUykgJW0jRg
WYffR2jU97mPqSaVdIozpkgdE3pcmCtm1hnKJX2fbZ0S7cDrBqlC5dnBICV3QlV9
xokZFGhlzzkI/w7Ya/HhliEuOxjIU44FrCvQlts593tcamI0Duaws5wkUYqWYh2T
TAkS6+z7rqHS63mhfQGW599rQTNnxenqWXU1DrHiL1d3hmmltZU1AMRJkNSIXdvf
4sfHFeQUBh/5eUN9m1dVWO9BXeateQUh2YDBV/ueL3s9+Rsi+Ke2X2No+t/kYMOE
2dXd19DgwiLkRBiDcLHu6H8BW34hSvCpIY04TiI8V11y3AAxi1b4D5kGvloAweNo
saM68Ckq2iMM7m1n9vfgAtgOTf0qgkN2trJTCTkgM78KiN4sPwhD1CIj55gi+P+f
a9TTWrp/FOUmS9me3cL7/PBoIMduyWHDIxPdb0qiG1b1FFuQv8p+Euxh5PKeZhc6
mJSqQ39xEuaSba2tZ5EFud4LuKmFd0MbNxEeL+PB1kCi7uE4GjCZ5qGCFI46nMN7
VlDsAobczTMKqc3fhDy0Ra4Nk/AbVS4z4YyyT3nN/8Ca4gG4S6r+6PS/pZI5+zWm
xrZ/8fEn49O9LfSQdQPRuOnUrpxZH2JJo+VC8C0+Y36i+CQrQT1FrmfRFQ4792Bf
Fa6OAunERE77nqEWRF8Mot/O/oZTUZjgh8zM02TNhoDv3pXjVC4BJHUdM7f1dKT7
iQlaZwOY68jKc9YrY/59zBCPUfSNIuZuy1L3sQAZ3clew5ULIZcdzadL+EgUCjKH
8Ul89U8NfD5VvHsolG0rRlMkAKtONkKJlZy07ftZ9En/9NP+G1kDU+jhfzV3mCwK
FyP9TILw1Tey4TXMxCt+BkmI/5XToC/Hzr8lF97ExxzvpuJ2OVG7+lcVq1vLC2Nj
cnHvObXDNtkyW7oCOK+cgyX2ptnETywYs0KV98frPbIy/oadsr6PMyKO/VzgYmTJ
Uh+bh7Rwj0+F5HQcjxmiDg3D/7VxeYbSrpXafkofClitqmHIYTbT4RApJFV9tZgr
66e6ta6vsqGBQJ2J9bwu0vzJdiW6Kz65iFeZBYSiKUSx7/bfAABnAAy4d+ai98IW
FNv/+/wBVtasbl0itE6DrwnX3k83h+VonBvGNrEUzl4dGBmY6dx/vpZy4ZzTphVg
37pwnm5oRnds0JuqGWsr5z5iqv/rVRQQJFYio/JGQe/wVdfgfe/Vk4T51NqO0wJO
iO+0zDiiBqsfPQaGksKNG20DJZYtdBLKPbrk1tUSVaCTPXB9fkXDarzAvNltT7o0
orO/YMFSAuuJ0krbkla2YOMyBbXJP31zaXL4B4h6FoeaJOCCno6dtpOJj4IkkCJ/
fWovPp01DAUailhvl/1AvA==
`protect END_PROTECTED
