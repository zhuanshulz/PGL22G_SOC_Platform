`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hLilTKWFi0MnxyFbKv7rnrX1ZOL/w4EFsB/TduIzEdhjhmHa9QKnW47txVS0l7O/
U7Hz7iZ29WP7cL7jFB5X62VYDXBI5IYWRzcK28tWvaK2yYk8xHCxiG9KDP6pSu0T
C0ykVkW6UN4Lbf0DeqSMpjt7pXovZOGi7uzY59+i1GvGNMc5BQ+vr879VmGcGjG1
RPCKjt8ZuCg+nxK7j6gl/pQEwO/YtxdPLSyQ4s/HrD8M8pfHP1NC+N85pxfcop7L
BJ3cXUWPNYK9kS51RD2A9RQPN6DKcVGerLSW4kebI985/DaHTyCkbnMKznfqu+B9
wiso6+3Kt9Kd5heaQ6Tf0RvaJph/bXVPPbEy82gLyb8VnGo6mrODBcpYLDX2xRwV
H3QePioINqihRauwqjV/PPNg3kPH9yX3AuQLIte4KbSh1lHWmgFqR3FIEldjyW3Z
ak8XOaM/Lr6DcoxPlWcwmVvz8ZP4Sd276pSWHJIjwGXC6I7ABLibtu8QttIx/9cG
+bUQguCIePWU9ahiufq/GJX1hVLc7lKzJqO4bo/SO3/2ACR1IKVLJK1IvErgX781
1nWDaU+w5/Wbpei60ubtGmD/MeVFpSxmJ8nwyQ2UPCNEed8niMnS66uE70x/0ADo
bGuTdfmFi9WOpS0TcoeytpHf/3vQMA9F99wBCupgdtsYwKANIaL9AE2wFBUhVIWs
8kQiMHkVvuD9uslThPPK6WW4CEfh/4Lc5EGT24cnZgnhno2/5me+cBt5oNLMBCay
BXhsfEsCKwyQ7L/YKZlB6AUwz+5mvfK+vFaYCOnH99mehnNS+v1poarCcKyYQ//z
sXaNwzJL4evBz0Ew+QIA6JoAs8D6xwh86CoCkvvaWauP0uKAkMEYJx5U51q0w0yR
/BTlziWxgdn3vwlzle6I8hhYGnSWAFNZHBegPMIuH/ApeGVEthflhp5szTf9Ukwo
lrc/1dwTD1eOpyU9+3hsMD1YwK+QalkzM6HH13yy5lSSZG2u0pEMELZgAx/VJWSN
CC7FC0TT8+bdjNp2gepFNna6Bnuk/li0qZFbRRKGaC6vsgSqaevV5Ni803lNN6b1
uqH5piUn1M0zJN3gHjQrmDGCRHmStNlOXcnaA3BkOmkwOutWrnfvYkR3dqss9xvM
OpCKZCk8aRwAwD1fDC4P5pTw2RSmB02/a9M8FVawojeWfjWeKb2zbtjF60fBgvej
oUXnRwH8nW/bcTL9aCNMPNiV5VUaGIHv7fXc3pPE7w/ThPpSE+1UcAnV4QW2+u5T
E/ddPYkZcwgolPXySUj+mzo45a0o1xcvva6ax27a5z7KtZEgOhiILLivJsTuScmq
zEtCr3hVKueWw7AaHJVmoRLCLLwmfqtAZvbbrcaS4jbAgthbNBU7eQfvOSlDZXhK
Yg4SMrnTxJM+Rrydi7rEStGQcESJ40yzZekNmoqpQzIxsEhWkzIvvO0aX0Jlpl1u
YLqDYErSF8NX4NVwajvc3N0c0u3fEHEzYYn/Gt3aqJlUdsjW1cvr+mW1ncXhw42D
tdn3uStMVvp3jeQ3EvUx5ZXhkJsrR3k3erbjeRWN6yXn+GXCZU3swrF96IG7WL3P
INadh02M7FS5mQ/RPwEz/lCkTQq5bu6v1Uqyw61JbFCH/w6yrHNDVNf2fjLDMxAR
Hv1NTYacFLiYNF0vfyIbKM6+OqQXsxhMB9i+aG6cYrLba5XCxQt+03fO8B4JETES
q7CUY7Ba4K1i79/mk/t+FavhUyvYOo38/qil5EvcR9vWUzyIUUPbdKN9KTtRyBV7
K0cc15OWTJN+hMW2z9BBCgdw1Zf5EoPHvVrxaOF5qudCiY8VkmA3AvwcnK8Dsqij
iU5xAbbHmO2IGt9n3YxlycT/LVqR6u+HRFC5MGbnoT4Srg5DJI1w6FDOGKO4Ic1F
jDxotdghDUo7IPl9ndn0vZcEJXvOThNJ/Q6wEA7i5+/EXigvgN4oWrYtpIQS2BQ0
H5Kw+72AVBdU/7VicSBN4c0VGWTcAIAyH9/2TqemE7MXksMsA8kqO0RSGdCC5V01
LjPpcf2++P/7cKeF17BxYPy1pAOykxnU6mPxiNPmTu+piS8zSVYPSQ2ysqfDh6ee
/oJYCy/bAObLaYlLbQmxumgkebIiXYDyhWzU34WFy9lgphHy9m+otlNRnw0lVHBa
lRyQS5MIAQJ7f/XZFIthQjPehMiKuiuIn2aA64UimcX0dx13in1iSYZwE7nOTY9d
DHwfr8D2tZKuyGokUC/TEIVC9Qy9ihopFNRE5gWut48VsAzBe68UnWXusFMc1M43
o4awPpQVihUuCHi2s3XPxTSzr3Id4OdL4YRQJAPtadCV0ghjQjXfdfjCprKhv/NC
qP/hxBz6hmFhSqC8n1SAk7fiE516jhmk2Ms9Od9+q3IpJQgSK9BK5uNacn+ItqrF
vW8uDdHfBG+MRYXHTkv6mlTBQJAW/BELs0xTxuTzIsjDMcCv6FUIMcDK4xOAq2Ow
QQ1JLIyYInpGRQz8kFuEA563+eJPwnI2IvuliUlN8/KsrJAflVwHt20k5nSoyt0J
orbihCWvN6p8NVr5JYgVcyRJaxihXW7r0d5ncIBuOZwbjTr6uCKf4lVe5hYPJdcO
h+T2U1Htlk2yAgLIY1yclqEnMGro6IVETcQBYo2IQvgzOoi6WitRh6htvWxy9gMU
XoKZnFaAEtjmF2OXq6joQeNETiyACrsfWMp0yma9Fk0VtKkkxj9VnQCKw5KL9u8i
anzOjIyOhxdtTr4YlX2q9GSdZeNVdE/gy+l5TlLC+czmgCVEM5ov9d84NvXND2Yf
0HLvXx9WiBgD1TUp6utrdnyQRKF+n3nNw8KixcVPuH5z0cI8mJD2WRvi4CO9jvvV
YwLKHn9EULalx6BTWI+kONB8fpVnqr514hJd74aL/ptwY8ZuzhyKT11s5mJmm9bu
wtZn5bvwnocNJmRxLKMzP2WqTGVdbHrYPGSzMC8IqVlD0JHvbv2k9/gIb9Q9/Qbd
`protect END_PROTECTED
