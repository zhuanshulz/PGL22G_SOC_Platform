`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GP0S2SkLVLcpcGPNlGrtK4bQL53WqAIYKCPYpCCBMi/wNjd40IqU55cXo9UZM31/
TpVFm0IilEKZyA0giSmKlWYBu3Of3MYN4dgsrCu5xEW5Ez1NjW7tdlwavLPzLJyh
VJ3SIQWN6zJxReKfPqeKg0OC4M0dJXG179b3thrWelUkYiNeR4/0nXlZ225CGbi+
LaxRGvN6TCKRfz8/8oah1CbQt2A7u268U4zmYk1hE/lA3ZHTQTEfId3HNDbBHErz
eJafkRY+wSfmsqjmqlLuiAHy8tLdTmmH/SSpgm/zdVnRc7XAPY2NEQHGUAXyZJTn
i26y/UTMeg/ZMJ7iPnaFWx9ODpxkIMt43jH9V3co8AxlNObfW4XYyo4ZLfQ8UTi0
gAjhAwM0K7x2cE3PGahpCaLJyjhnGnmWa86yMolrhFpD3slVTxKhIlRaaKS6GYy0
6b6XjHt2fHAq994OQp1rwoRsbp9D2jQodPD3fIr6nqzkNDS6pE4JBIHXv3ZnzW9l
MLiUhg89YvGHc/BdEl/rboPg4VYq9KsC+aGMZOnzKBO5D9aqIbyVkUpkkSwoObLI
PuNShh7Lqh/ei0CPAFM3TTohg/3n1FBl2q8213gLaiNU8EmLYxnyG8jV5ICZWRsq
b3jvY8KIarEHaNQhoc/Tl6OKfjE1Z5gdC/6OqqUtrFrKE/mM6y18ESORkxEg4Lri
ccKHFRhbjwjGTFX4NjIuG3VI3nIDaSGqTC7IEqtRIvt5pBBlw2+xqvgU/O1/UR9E
R3ue7AYlGAW7kFY0gVFb9gOuoM7TzH3e6mkZQWqhRzqHjR348qOzJGBaiNlOX5Ll
lJ6vKL3XdIEflu1K8HYwIcuN6V1o5yZSKV23Psw6XxZif0ZjH3qbyhfAbaR25GyU
dBF/H2FbKpgAhjNscgz74reX3/nMUgFfbK0ewsFYtpnvO3x4CE4eMxMzOEb9p0iW
dJwxueODXThoVTA3o+sI/C24U6GDXDQWDByCTJ8jkP2qD7HBjdROMZB0/FmVgjHt
Tr4B4lHEpMIWv9/4OdsM0XlnbD5a/gnsIr5Ty17zk4APr56lrKPsDbtA7QcY+6MO
`protect END_PROTECTED
