`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CKZ2FvGMe6benQgumWbB8L8xXSuCJ2mX7P25OvcP9p3QKMm9aqxPo6PyQgzyNrOJ
rN60MfG5eCljvTbOT70LqmzjqwVDP7uuFthyfmBaR79ANIze3pbwPOkQx5sizp+b
KvCI6gxunluoqBFEbCaR6LGRj8d54b25jdaFNwkh4KONuAgrhfjYcjmTLMs9HD93
GYMbRgSJrBYUQd8BuBgjxbon/4lTeyweoSGJN8ypgXFOsPpD8If1DwLA+oK9pe8F
Qu4l/1ik/Lh936v5YznGXFuCLHDInY6o9u5rE5LPkwb7eaiL5HnMG45LfiAoPLoZ
V94sDYQOYssl0+giv+ips81tp2d0txzQUH0kR5lyIFVpMmuNekWCmgJDC4zTEP29
5WPvFWdDM7rGw/+G5AnNlsIqfcZHjaEXzWLkCJSn9oHz+OmOS6z10PNRZHu3lfoE
JmGEW9RKrppjXQMeDHiwomNEViZxbsRd3lsW19GZqj6v9sgixWjD7OGXOuj83NXu
0YvOSxtyTce8qLlyHtvQfebopGgBRVDWDieB2XUZqoHOSMGFfyqSLk3sTPqjBPWC
X1Mm/9CgS3PyRvI7YzjV1WD1c5b54KYjI7kPsYjyMe9N3gFv8WsNvsyDXsmkjrkE
hJBCLyru6cKZOuY4TO+d1pL8rwcBQ2Sxf2sW7uzlwOTSLNZDX/0HayLHZyjUBdKs
lgsa3jCm1eCyoqIabVmqOArVWimcmsEGCDyMLFTQ/ayaNlxbMFuTJ9qTKcgeQdqS
LWM5dfsF5eJQ+HatQrQp5uqdVIORDuTEyOBcO6pT88HiNFn2xtzhLsoDdt6b+ofY
GPxi7lAuMPdooFvCi2yWZIUwritAoeX7dM1CKNzKQEwGcHJQ0Ot6Zr4i1dW2tmdu
b7LVDlsGdLjoTdjC4nBd/8bzCLtPS5Lheybr8Br4CtyE+pw3oMoxSiCSM8gbFKo+
TDG3drNaGxjKjJdbTUBhWt1/NPZ6UmTn0T9Q3muYgN5gXG0WI3QhbhDA2VF1mRvJ
sRiFvCiSc7VqKjeTrlTG9uaxXwLPj31rzEpLTa6juPecOMqiE40BeHXUwpgeCbZC
YdWUIykRtNE+T/xFR5zbFiL6YS4dcCfaDsigtmXziHUwypfhl1t6DQwf/i6/xSyr
j91y+sDgh/mOCzmP+1xbh67M85HZFOlXiaMLHWSTBER+uxa2x4fjYKnd9EYyNLnu
6BvBu/16Gr04kiEG/hyuoJ0N1LsfbcK756JhEmWn/5trxPGa0ZKG+W5DII8A9xLt
+J4szJX5Vsm3ZuWyE45jYhQVbDVgf+fHZIc7xADax/47JPm0PG3FV8Zi07zRH3S4
kKreukHWBM6873Cq5+w0lliOIwFx6PoFkbCdCWTtrzDr0kdOf4xJaF180wkgcchY
bvs95Qe8u9ldAiZArCfqEbX6ZpJcwNpuQ/T/ZhOymHqtP/zKDM65YknkverYJJ3U
iZlpIq/I5+Wp4kE2cqIE0Y+BUz7XwGyjvXisSWrj9zHN+AWt3SHuh/SmeWbz9NA9
htaf3Oz5tM6Rl5b2w8QlR9q71pg8czz7ItE2MdlglCBNygwSid1EyPVF65D9/ATR
ixYGCAESmla1A5X8IIxdb+wc/oYl9w6PMQHLObAZv67YfRhW27zAsnyp5FNSAU0+
K8ahLGydTUf78WE5b7EjOknK+fWCRaaDS2nElLaD58DFNjd4s9lU/NL6FzLjguRc
BONmiW/lgoPztED2gPnYNYKsMdw4D4uehSY2WqN4d/DF/ux5P1ghb7b5FcHVTlVv
ALxlAjXKw+EDax9DgkYxRd+gXaq1N+Pgg+98F0zEZdFX8rLwAwE3Up84o9aLap4+
WcSUVK5GunDx19KvsKwY1FdAomVKkAYwHGiUbI4GNWguIydNGxDVraED16PzuJhb
7EC1CPlvBDkIwvNxckk9TDLvLQ3FiH8r8u4gE52lBZ57DqtiUkn5gend2jC2c8kG
ZezEY08HfY9vsOQAaIg31SiC+X52fIqMw1JE560ZswPuDVqdGECf3QHKbEd+kSjE
hYuUFhW8eQJ9MXaAyevapS1+TGmH5g8aBLT2xNNLKDVBbB6TmSo4OXxcGu6H6m+O
QS5SCSAigdI8hAkVaI1VF5DG/eGIKw2cluKjyl4SgGZJbhRPPRndn/l+o0s3Iy+b
0QjfDwxGftIeXt5ICNSKYovdcL1wvwvK/RaqyOaebFDxVo9s+DAqElJbASyDtxAc
VtUmqsnOOPBAedqxKoaLc+YivjHA6Q/ygYmernB4AytyEHbGbp/anlB2I0/reXMB
ypkXnYVss0ocRqvUxhuJJjX8tpX47X6OotizPeIUJjzR9uaEdZOy1mPWBlLsJtTw
WwolYklJyEVShFECl62wYkHpKeKq/g9+P/gC2YDzDddD6D+YMRb+La0bTjHVWUC+
Wzawsv2ihSrvkluUf0rtCf7PbHi8RKeM95KDncXVqwMht+EeZszirxu4DXChoKjo
6kB9fpMMgnObUjHq4E1w4HXA5nyBqOClXpdLvG26THXSR3+dUy9MCMNERJuUmxzI
ZD4NU43s9SsMUG5WT9nrpaW+97UYstrHlv3H0Vbo0wtF0Iqzl+EsvMEyburicl4k
Pk+wG7Z0DEMP7ASuTOFXowBTKzxQxtJSKrUiWRQt4BAhPq/hxkE5Ez5D678hqkNW
HsLcvWOpxv2p3K4Z6YGCQvHIBncrMiq/mV1Bs+pwLjLmA7Fxvl5/MajPOtvwF/g2
2C8ctFerbGXhryhRRwJcTLB0id7MdxFJJsDCnrAEXRVJx5+GerUx6iAwycS3Tfa4
MEtDvVqt+xmM3JfW5GY7j/ktEI6K67P3N6qlcM0K7886KKUdl8EUBTpFF8zJFVB4
7S9fgi7iA9TUgwXUWY/c1baEjlJE8n2lSOXKaa11zxjFSKAhcDkBZmsYTCWIW4YO
Z++nSDWYuWjRhptZQE7MUkFrdqTwJBhW0P8m/K7bbJJNJVU5Lk7FyTjSIktcke+L
Gu38q/qixGQ2LL5S5IPnhGlxwuHcsnPsOH1X0v698K+LuG/twH/cHFze1KOA2ueA
3pxTcU4g0jDHuzbIPUpBgx0zAe1sKNAclxHVB/hbkorqxji81PcV9kXu+IIuyTAT
wyF7tEoTlEax9TvHUkX4k7z/EqXS7VFWPtzhqDNvGQctuwXe7ErPq/ger5pkERG9
jFZ9skVKLNXjUBz8J5Vwp7p9PLiImt4nyxiSECWM+ZzEznKkPrFeAYYoyDmM4jxr
3sPhSlXaOmoEN9KZ1qNwzjuT1BJmqJdgFGcdNE1IpiDT9UeM5JMX5KFQOBSKZbFG
IbyPb0yRdatP5aZuw89pFoSeWO2NbIRiCwxcx3kQy0eCraa8Jvx14KvTQ7Uq/nvN
Pki5DM4jZPmQzHNE6/xKPAU4IkyQllfsoQBa3JopX8PsQ0sT4JzJabHQbQH/i30Z
nbUZ3+08KriXz3DSfnw5WdOGpikZam9RAnvHg8tsjq89WMaiNVvWBxUWhf7Fcwnv
JndLedvuFnTWbRKR8ZrEIZtxH8dL/6ST0Pdzi9K27a20Hmi055Dcfz4TB6EQTOct
mgkSkxVG4dKoOUCcbPF1v8/2B2jjA6BWcTZOHXeNnZdLrl1SDWT7M9Fz/N5d2P/J
M3pETkuMJ6LEtOFQ7AxAoC1H1/aTKR1efqK8v9wT8uJJpxHfoaloOFiZgbBzbxLz
0ayhs8j7SrfAV4koUXzEqUltuJVcje1D0PIDZNrCGzniDCt7qQvvk4VEo8qZY9nB
OLdx1VSqEYdRhvZOAR/LPIElvN1ogYjNmHMVsBCgAnOvZ7Tqc9CbyfBjqMknKRS1
FLalnTV3kw69ct1fsNEmfMxEUycckCT4Csee+eIY6SDISJnQJZK2zIoMO/dh86Oz
BaKDiD1fnE+UXzU6zbdpyRjRW4miBbzRiH/F/uNQN06fDHS8VssWJernHQHo3JZJ
ipc0DknWA2wIK2hn7RxthN9yAu1WCf1wvgWBh9vCrSCqdpqF53x49WRtoXT8O4H9
HXRMeuRoRGAlKmXHt8nEpVVbW3GNQiP+XhUvQhfzg694F6gW8hPNs9YpqZOPcXsf
fBzBy6ABM3aKFv7TkcPDhI6dpNvwzxu9wmNykGz/TmZgFz2n7OlJMH6h2H3ZrpOs
0nz2EP4GE7HscgQddz+zCQq/7ujySq+eTt2KT0NnRVupoETMvUZxsmlbJePNrMFx
VufRQ1ocToLeDr72v/HUv4aPqRWBZtiADK28TzZWM/wOC4IUCZZ6QpTfT8umf4/5
3AyGOe/ecVUPjMnuSAyTNY0HAjh94/DRwyj5+YXGm9xTNzaz5kZ4FiXScBv+6edY
PyEtlO19ru4BiXcwEMYGB8dnQHNCjN2A1GnQ7gVTtHeJqAiN2w13JvEKfSsdpDfB
AY+Y8VUXhs1dk7bHa+gMaYxLE1VXFdvkFZc4bpAnQjMhkiLbXRXZe9F8vnopCB+L
5OMayIlrHW9S9bSWnyWgdEeFvNvR5eRu1PJ1IeiSa7PI0OyjlzUmu5o39LoshLbM
qA88cWq87wWGzT1mmH4bGItJxlaMbJ/dRGmjk1meD4mAmaVApYILhlKXS08PUpE4
0U2xS2ICyzU8qrA6BVNG12unZCiZlEgJvRa5kID9OBEKhtHvD1TIbGF66XR6G9QP
maCOOgNAzRT+m6wPHw5ZLimHBnWit1qw+073ova+pCBAB2E5cwrPaXOfCRsh4vaf
wqx9CT8OXVscvBVPQk5ce61lpXjars4DoQ71Y3JzHGU/KaEqtOFYGK5T9FqCJPUC
R8PNIy91qWSlzxE4t3p/1rGPrZBAyVLmiba5OeZkarLB+EhnZ+Yv1H3RdWQrlJvI
G38zUD53P5aUGMFJ41GY/NoV3FeOt22l7gj7UfrB7Xur2h1alJRvHdAgyzoAGoFQ
xpQREMRJMmeViqIx311TgzdQQVsMYAKhq4bV+StRWva0oieP/lAgoZR9dPkybSMY
orO4xJp6Na97WK/8Y/uWF6K/QxVwiGGNwWHLUU0u6xpDEPgbnAq+EWHkYbSxbta2
iuOh9mQc//fyGOT0RXqeQUHqXwTEyUxe8mb+MB6OCa0yquRY7cAOmRxX43njWikn
7foRislMYAdNh4SoDcJn56tfw6mT2FIIHMhSNr/JcIAOGTdL4uvb2N03kLX+d7G7
72Q15Nwg88Kl0tECXnmuZfuP2VRLddBsOuHH0dJkM4pXo5gYeEldpfFnLRRmXS/Z
yjNwgcP/g6DIZWXH0z7o2HT7HtMKIHguRTfnj0enxV8INO1NdIxm4haGRSOM3YRx
TZSObv03zMhbom8gZ88N8CFtDmW816NtZaMtMpstZ3RK2ymMwkv7kn9B1ktsbEiY
DkZPaamQEHbbLOBrTJ16MA09d9Ae69A4B+424rC7eeKOnLjd5GoE9QVyqMj5HHGi
kd+xE6blBBkEuydbtV4dGNgPA8Kg6YuZqknjL/gsLAOWZJ0T/vg5kcQVcyWnnZHZ
wLUoc71pUDj9GErUzB832JtrMuueI7XvsUK4SFRUboXh3EI70/d0E5TXxIx2oL/Q
h61UHRrKB77UKpH3gLtq+faucta/NJ//yYi6q7KlhC450Ggmm+IlxGWPMs/NBrZC
DYS2q4d5xrcsuczmK9E2Afd6DVd9RdqkS7b+z4VzPCUDe90fNnadKiY3gvCUa+Zk
rHONPHDtkZ4ewGxp1eKx7+/go0ZSMwyHfwmbQV3Jdxqegg3SEm9FI6tBtbVj2daw
YvW1XZlR8Gkkk+mxbKaWKztnVRUvW8aRM8QFvMS/ZBI3faP7tg3Tz8mKoBCQptoL
8c2IiuV/clh3VKHj19UKWRaOdl2L2TrliHdPtr+TDIzwKNMTRaX2FJ6keMa8OW06
iN0EFjeCsHJOvdHtrwhOIdUoZrPjW1jh9FFiZ+cT1MIo0xHnsA3ue5p3FrsYx3nX
ZL/Xl+2mG9+qGe6Qg1Tm3RE9U6kstsGIfadILujUUpDeiKKWAauy2j+58CFnE6zg
RpqCVuqXDpvSq5ONZKag9b1xYKPKXq9nwpm7of8BwyUNXQ20aQI2RnIc3VWqmM9M
DB5Ntquh8e32GWgxI7gFfls3m2FGSeGylquG2M/OgcRzi+id4r4G3Yp7yB2H6KRA
0PuG3UVbnqOWq/AaZ9PltiWH219ZEOWKCTu2w/8iGjSDkc/6BjeOFPJYJTmuAZVd
nGG9ciI0marUTfdrNuos5t/qkwOT1BuYBhZFBYEghCcl7CHiabsGek4s4KuNuq5P
GbMxAJ+EFRcephOOGcRx6Yg9BQ/EzMn5eTyhmUJfRtoNcYnSVGf/igqkVL0aa/og
rJDUEmDyqUM87KCLiVN7HZF2JnYmnxn+PNW1nBNLDfwLZOW2u4m4UZY27jI7ca4W
YqS1jnWrVfb29Cf8vsr6DZp8POlGb/i1TD/MnqiWweDgu+coDO/4tU/314eKDt54
cpDPA3Q/MEjtYEnvrT8CpfGo7FGYKgXVUUIoTFbtRaABzfT4k+UiYcPjURtZm9UB
teET/7Nfoo0dOJ5HWA4xMoz/a85Gx9453llbaPQomlgh4u6AyX5tunO9J2QQZ1sT
YCGpAyIIP+QC5sRN9snmt5kSzj3uWhUmEHNPxOBX2LqRS8wE2XqL6EezWsdGdoXU
iJtk2B4fCkjqyhKqv4qBwAXLvpDi7Fg45yZp8LF2iAbw2sVFICPjUJxV0Qx/6aO0
4VCzjISptCcNcY0cxlz0YsIa4FLfB5UBKiyLW3M7fv8=
`protect END_PROTECTED
