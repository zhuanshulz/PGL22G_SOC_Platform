`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZnGoF4DF+BG16DpgXVLwgUAdZC/79mWpcmh0JgSZ3Akqh5Bq4yQ0f+ye6hxugQT9
BZ7tRdB5kokPJRgVllsoQBsM/5oEF+bLcPWgn2+faNQUTWMSBeXVk63nkyA8ayNO
9M5h3K7uuPoRmWb1By8h9nhvKWjo20rufiN2e5yYe+iXfru7akkMySRovfXz4/aW
1FEnIcIsI7rzDmoAfdZT+vagAs4IBF3TTfiPmvRC4lgTonML2midx99Ebk2unz3h
M6lEhZp0NGjwVJ6AyTcEUb5CkBiCPgGl6KzsPSTa7a6HSqwwxeDQDMsaJsfjETjD
0PKOdOWvzlRHsojKeTdP1d6nxDWugXeK9DcWNPdwzR56xzn8+vDIvma+59qa5j/4
csFRhjBDmI+972+HPyZ2JGSjlXJEi9X1X1y5hlnZusvnERMKwNzXqj/J8qSHM6Gw
D3P9ij0t8R5M8IBb9Mz5Tovds7G4GQi2SYn3bBJ270GCYy4leHPcGki3fpSaYfoE
ljyzJZwzN47Sr1r4zJxjAw==
`protect END_PROTECTED
