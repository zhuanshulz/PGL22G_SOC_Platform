`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q4Hu5B6NuIOQ0cb1KrGXbWDEQaoWKXmH9hyzzh3x4O6cU6AJF3fJq2Vjn9ws1+1r
QT9+bFBSratehjh4OMQ/ajvYn5sUuqn3K+j6dsw0PzIBsUUvGBrVHhqgUhqEOCXG
cqy558azXmuOok0BuY27TSZKw4nBrltdskOMBsRL/fBbrwlM3uFuoKmF0gr1C9cz
RkljSoz5XZSif6AeVrOlzmPoyO1FCOlb3Ze2fGbJxG08aB/hi8DCrOUdXJJksxBN
JwLSbvRc8r8YShnX7f/bQkjY/IF58LEHa0GcDsnEbVdVyU7Z31yxNc3YIqpoYsVx
WPWq2wVFk/SGX9v3N06UirJRhr8LnPCjy/8G5xVflVew5flspY4wQOS6B1mGaImX
IYEmUq8V/WFOQKaPPSXm0zWdmLqZcCUTNMmMWFUkypFszcAQiRDdkN05KbqAHGhH
6cQYTH7jRTr4WQsqJ+9hLfU1Vxh5hPuOdHk6LUoaRc45uLpJhtPeZ8GsNbC1mUy/
Qx2Wh8rnKELeAHrtnSMGtQ==
`protect END_PROTECTED
