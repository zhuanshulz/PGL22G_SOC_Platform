`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fNxCH1e7i2rQhSOJ+uCUNrDHAIF+RxHCrqU9rUc8i9R2g84AvQMaLqlBnQWPx8yR
7oo65GmrbrwExSUuIIg6aVem3xup4ZnqCoFtq3QTc+TdUZkexvuVROhprzzRuGXJ
yztb9pt0QgslAoAjnqxptGrUExFkU3LPKQ4+ASO4qllJwvK6bLFms56eBj5qtpB8
OXW7/b6eGOUrx/lI0Z2mTXfij742U4krNi+bzUlxvLRRGKnpm80vyQeEtQXWVSOa
hJkQFElgz0xkNA0xiR+cxT2kAyZnDoJHplVthoQxwh+troey2erVb2eqZkT+Gaba
RkPfvBMVM9rxuoeWNNQhzSq/CAV1cexOny1ltrYM0989bEle0gs9ThRpjPTxcAjI
cX4lV7YoDeLrKMkO5Rj18tcJilfWlioBWy/vG4uUv9rSI7gbb0PmQIknexLew/Bo
7fkVJbRl9zb0/JTVyo55AbmCVtCOBpwGPocpLktP33W0ARLYNpH9PnEUJCOBkvK9
BqqpMLQze/nrrhULxkBK8br8zvUy+sX5v2r6Xy6/umLZUk4pAuG59OdYRF2Xsexr
ruowmL7EE3EEHOtP4bwpgG3RuDAqR7XqUxZsb5XiUCPxbM+pjeTZh0wfNXLmC5+z
iGCdhvsGaHyuhL5fX7aAY/WPQVcyVw8EFedc+EQkEETgLY9F3gaiI2cl6BLpssgO
GZrluLOPB7YCVEPm+B6jtlB4JBvzneOnXeeEB/IQBkzs5OZrmZRxcyrIoGXn/yqr
2B7jD1JUr4hg35p6KLcmymgxpiK4IMSqdBcBjoyx3AG6ZldN9k5ClU7rXxZHleyM
2tJ2V0I6fooVQJFQ4+GaJmuPw4TSfA27VgmYmJ3CN6bk9EGebuQUonqZ8+dRJBzZ
PoUtSiw4OlprflYT+kFs6PzSND0XxnSJRSjOJGhbJ+I=
`protect END_PROTECTED
