`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n2lMubn72K1vjMrcaNhPiEz3iLrtCRj0B1wLXXLCF5Q7XJod2HkTZNf7Am6VNHW1
Uw52Ao9r30Imkbv/yGANS5EdPxUiu9QO436wpdizDIU89cUF6A4HpijsejuM1seT
gOtvlA4MrUrJcxuVofIYHgRGRDfL0IhZy3wFzpD6jxESEj9GX845bqRPOznAUAPL
e5Nxm9Btv+1UVtUNa0KwwhenRioKW6EfaJ7CFBV3Rxiz2y5DtATmBDDIEPWQMMbx
67REiFLorGGxtuXfBvhsp1nAJBuca913BrcBgRxOPD8sO69hfMSa0PyxLp3lx+GD
AKBXusp+R3wnSaPRLvXmY5QZogiCcXSYyjv1Z+tScu501islJj+qw2eTr2Vx/vf/
0A5GUvbQ9fgE5J8/Cg1JRHVf5mRcEoInivnpN+Dd0LKJ2qou+Lu2ArSHS8nteSkO
NKhnB6+mc+MKCCu/R5SV3esDLMa2PI3GnewUKVVbeaWO9d/aFTbSmTrRWKqP8jIH
Ie29iHmw3cfzIBm8FvcKDmCr9lyrvw6AWX0qMMOqmcwRNdgurNpfEEYpE6jKTfn3
+Oy/9fa937CmJRU7pb4VUddblwtdARKhoMpxcdKnCe4LsD1SfPjXECSyjtU48/wt
FvSqFUoLbXgaz1hwOoZdwKqcIc+FLgtubow5LLMmbEDkXSVONwD+0dhdpZvkJAZZ
4smxsGjCw4UImtBD1ZEgmrEpx7a1czcAE6FtLGuQRpSbEcMrG//wzZ+USwL9sbYH
jmZ/PpxNSyVS2jno9GEkW19PAdAdL2n3JmtT0YQcNpDARIR741McNjIe2E80SDrF
IcC/3lyTc4eU0gJU8uJV6vilF+W97YtxoD2arpe9w68lnwMKk/TkdKM6EH3eutbP
6HXCY41WriZZUi/YOWkj8flk7wuU2gzEyFPNwYB/Dr2LS9q8DvWzPJSuBiMTB3fi
vFLIUC4KtbFjdiZYqZmgcmM6wKMhwDnJ6RM9MPqIPhsO39r2cZm+f3pBpQYAcW64
UwMv2OOGSu1RohO+EA/ZYSvgD0e7ph3DVQEBRcDzW5BLQbp5oEipzA6628NYV1BZ
XJvzwy+Ij/jZJoHgLxRWzr3ZEg/8P63rbTbC1M0sfP8m+rkj12b0v3Tdapi6sIZj
ZrmVlLeeC4XbCFk3+hwWOZzpheFnTCTleA1j7wQsw8DLiJgQ4tIpzY8BDR26P+uQ
HGClwLqA4KmVC+pPJJuWqKtbSBAWL5+8pHbIBlV2GhGFol+lpvfHgu63PKbpAa21
vqoCwcRsHwlrwYsw7umAC+6g5t473qzzake7Qc8Z/grq3iPnCLmPn7F0WIfzNb+X
n5pMbwEvt3uaxhGrNM88Lg6d/90CPL0qUld/XpvO4sOBwc8cRtiwSC41nCieCqLx
Nhst+OLnPI2aCWsVC/2ecMr+g7LN11+NlIqZau8mkH1XcbtGLdkcbigBYb/nlMlC
Ow99F51JEWRxo8lPxp5ZxPiBpE5OdWa50RacI6E839hiVsD5MVWUG2+ymrdTsMxd
2rRJGHhcN2tlPNdXPp/OpZ0Vt0PX1vd8+yNaU5HuUGArai+7HlgVff8f5ysfmpEN
OBqGrucuuEj2WwNraqkwtzYczg20Ud8LnwGFEdXCIqkoifApI6GuceMly7O32Vzl
CW8VDgQKNBxyBzM7U8RhyY0+82Zf7G4fVj58w3ndg/iDC+H6hcfbtCWJr+zRADGs
70Y3UMiQ2PuR7In4yEaM0xVe4Wp5QTk5pw6xf+pL5wlzJzBn3gvJresRbvuc3XSE
xGf6bn/XRxiqN/DfvkeP6LU6sljpCxrEBfFusMzSU+sajOlSdufDezUfI4//zLQh
9rXRV0x6C8EWRnkbuD9Lc0z3VBk8Sw2ATT62N+zR25/seimwp6ykk659GruU+qcM
gdBXXX5rhzbJeGKO/tvRywH54t5DqnU/sIX8J/d4gyT0ww1sLVlcr62k6//yAe5m
tsN48yLet0nY5gq7ngo0BpSfylhbfddWTcD5qRX/FML07xkFV8cAwRa5qUKoKSGV
t4xXXvQpjeTf20Umz/OmPrf/sFU+sc1B0WDc44Lcx1OXL5VYOMyltuR1nSZKe7ol
4oQ/FUAngKOimDPkZEGyr0U/+NQ1xvFyLxRcwmOaK6VMvBGo7WIimTGqgMBYQ40N
p39iE5Ltmo1i32+ktlNZYasBR3VEC9fYbCYrQKSM9qNJuT7dAUdZy6zdMGv/8xDI
gPKT595hhxDTAHCPSvWdzxaJqpf43HA8Ki4PMipA41Mt2ROjbl7HcL7pCIw/0A9L
2ppeX3UORRv6Qy6A+4KI87ZAcfqr7UYrx8vFbwYUaREQMEO3xmW2AtGT3rhwNRzX
QGe1B3sqt9oMGzNgCLOtvAmMPIX7/Rq/14IKTf1dyS0HrKGhz7ZMHUykmA4Hy70S
XrPT61YfLqxPPfB3skIItGZGENxNATZGpaajdO6Ie7Ivzh2xvRbrLEaAU/RUSXbC
YNYlw+3VwA9ax/s7pVTAlFpCkMo9nZs9Rde+vpBWRPaIL6ITic3gTUalwmOtv/f0
YZFmuAtfa7v7dA7Ib+gLhBr6rOgpqndAx3bFMFjuvd0Db/V48H+lpzAq7/L7lltg
ofWOyphDQa+egHc8s1SX3GIk7WAfzlu44pSYM63ZXm+/nK/u0NdqRKuJldeGvBOC
dBFFX7vMyPEcWyB5nayA0zmuoKm1HHmY9/SDQwQ4/E+v2ZdT91T5RboNci2LxoQA
N3w+8vJYcX9LmmMDNItkNVAS4n/sTThVewLRvX/d1Y98YgD41TwE0qWx2+xh/4ok
MrfCC84KV66tKh4fQ/PTWtGsSgEplNU2/OQwd8GEMWzicq19YwJCZsrNrUKU5WVf
eGS4SDf/kgpY3EPzOqUyLiYEc2rw2gM0NXcipsH3T9M1aGtxPuUP/v25UW2mKMKc
MlDibkthrYvAe09AzK3UmgBPAx9qx9Kl0/JPifizBj3H3FeLm2ceBmMtDoHtm4ts
mb/S/qsQ+TXrH8tzZKrTBN0/BoBqkYtrnIQ3/G96QGk5KFfnFZLcaluXzZ/5oZMf
vguIQFtRoqYE01geawdof++ukPlhL8AukU6SGzSSvAfH+tzgYOzTdOU0w0BvUg7u
0TjvqWbrMSaHJs0k3oY47SDgPCXmn/O/+xC62mDmlwFL/1zXTdhLxiHCkP9h1/12
QWh5xQyyAhhDpWHykK1bMBxi3tnFo+FcoJ0p4y7qqGxR7PAsENMBv7uput8sJ0G7
h7K20AE0gyr0+cBsq9C1+zcHi40IsCRFCOIUahIyVCIM8L/TpliQ91M0a8n4hxjn
JTXKbuAEE+4tfObnjYQx9PqFyqBEqW5WL5kTJEUHjC1M0fZtQA7DiTGxIn9M0q9x
BUn/mYHuR8C4OyVRzen4McXWutK4XTn5Ly+ytHy+D0TLvxOExcRBXzsgJy662pEH
wo+pO3pBkeDGqoz0A1VnkK+C0d6C2PknH5Z8qP+xPepOtOE+0kDaaCduDMDIA7nT
ybjwOHa+GB1YRmRTNkVcX1mnXinZGXI/TtMfI4CoAsY=
`protect END_PROTECTED
