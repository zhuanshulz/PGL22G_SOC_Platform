`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tno2Z8D/7pKHgKDlZDA6s6XHpK3cCSOuAO9qqfOiUDRdb0uZchMEHQwfvYEMyFq3
xI0Sx+/1zJXOam9rqUb1qh8WTnl5L0zF+cxWiaMSJKsa95aCE3NJjkorlVCkAfUr
kZ9xJTZnodQWpxfDzl6TXkYpbVykyh0MCzk3MlCMrfM3Qa71Z5HMQ6rmr6IInJbt
HClnz8d4/QQ+Hne59E9GiWHAvs8nwD7fVophzF3zOHl7qDTbo0bog4Y0p1BDIqcz
WPCz2HW6aMLb1H8k0FdC88X1qlvN8Qc0X7xIUiMUbuL0gSm4eZ4PRGpvZpH8g1ml
qRt8+Rbn6LUdNrxeN7cPxyqWpI7u/oYbPBK2xhk7E/YVrigpXTMEBWoM2QjcZjkz
HjTMuN8xC+jWNUjb/NOXA0IbnkbAGUneIE5f6r6slzYiHz+8ylORAIkMMGi6FD67
iEstrPlymVpgMBq2qPmZXRdH8fBGmF/WAsGSFQkgjXnNvt//PCJYLPKOy8KwqS6Y
pGmR3661i75tmzdiN5sSmgqy81LxlwUyzeAn94wcF+AfdrTvrsGcfc8BjM07DP7h
4QLMMPHNmqazjyZJW/0ZBpcS5XUCnAUeF5ImBYtEo8VZJGXQmbc2OlfwU+QwKM2R
tIENRKBRDs1dQCLPSLGph+OoNnIqPxHnah1BV0CBKaBC7Vo8VrKE43U/aiaYJtqL
MywFcjDkq7lZSOquRzJ68u4VahTf0GVhEmpaif9Og1jCq98OrZ8lhXpBueXK5bD1
TOHgpIy1yFEhymWnYDfJ+SRmFHHmG/Q0shhqN77wt1oqYuwmkhRuJwG3tRbwHF40
KpJlQy149+KB8tMBJ1Gp2oPI/rRqjD/cnCMvF7LIgnaBUnhh4qTCAaPzDFeo95up
S7VLWoeXsxQqMbOlqZ4EjeBTGKgB1cdIZR22jlKsUBIxlDX4iyFfEYfRj0cxnPT8
lNUfbyppbVzoLulGe1MTPQbKDR+QnopSUMW1KCaJjXqAQhsjVsHPjuFnHiom0aoM
2FYSA3X96y7Bx2UfyNNR7OmFhPvDtRwAlF98sFdzvveUnur+KDbd5whWBHUhNM3V
KIlBj8BRhZadrCjLMe7mmw==
`protect END_PROTECTED
