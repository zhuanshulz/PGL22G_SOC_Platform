`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t0S/faTcOnfi2Ax0wqZIbFect14dh0Ycmvn5yKDpC7/BLRzT0Lo2EfisCWjwplfK
1CJb6f3FyyyGzYfYBuDkUesvDbK5KToXRZsHZXagUBF5rBPIjE/FXNChvsUejQXN
g2rGA4xJFhMh+zz0Fx2Z2V3Pi4ThhAPn8LcrktxnMdZU4y8Y8MVU1sgteIctMCZH
JtEKDP4x2J9GZiaE2Z7OXLabKo+PmTmGx+muxaV37vd3nPo0BTDV+l5dTvjmuaqT
j2x7W48vB/wlEhx2NSnozb6ltpvm9bSJ+vhu4/up5iGjDArstTw1AZH1F10r/cQE
CY2m9YeYGyNdQyKjsanKRIG65nlJ+oXNRfdaxZNPmF6zHYDnxMRk71tCp35Vc3Bb
jcLKf8tga/+0OvbBMOkNqtjlG99Qk+0XNVzSqNPadIrvo6rVsU9BIxcq9GFT/ksI
pyr8mpa3J3UKU4vIMVXiEPgGAQIMGe0IkJ7+0S/mU0QJlmL6lt9/ESDKgW4yXFHK
4F4JDYIPljlNGsoNYikphj3vWbptrKTye5bOmvRRovttf/UNN96eZvw/A4vbiRuj
NZaHA4U7zAJu7SksadrSS/Ouhor6wS7OfuAJt3BD9j4jHA0ZXaQgyGBjlANXbxjp
g3ePclJV7E2WswVtF+dBPmpoZ6jY5MUTYax/cLrZvuTRH47tF3UQC72DRCvNQCVA
dmC6mhyJxXQgiQraQxqwV3n/dPGMLOYEFV9FoCsUnjvY+7O7qadWR20xSyqY6N/a
kObsOE69wKCYOrahGESzpSE0iSWjOLsKFiJlNB0tUgNAMjMLNX3tUhz+w2GS6tZW
HGJblgzQCHrofhDWeJWRSnF9IjDY3/WGz4FoRmp1cGFNuWhMbNg70DbDrnTnbG1x
FYBhe2Jpp/6tyCGkOUv+yBydwta8x87PnTesJk0nEar3N7oDxVOZQjeUjJjwh6gI
mPQV/Bi6YT6yUvxz0w6C0h6i1Svm8q49ssvoCrJWcRjtSK0p3Imw5VDvpbLCE/YS
ipIsTb+s5Zc8pU+/IK2iW1P/Kz3ppQMdhOV6M1zbkmovQaKvtrF6BjhhvSm5I5UT
WspuhLy/Kv6a8CnZCya4G94iwqGdUD+/4MnPnHvK/0FiJbSGpHSEUtdGwbg2z3hO
2HEimJOW+eh7laMlOioEfwWXe+ZC4FK5Ad2BscAcpIPYG2/2mnayzU9Jji8RSP07
dW5aR16qj1T1iGCC0xxoRbl+KH+XZmligu9OCynnLmZqnJSyu4Vcp4eTYc4/aRed
uadZcnT4Qn7TnFFa5Mi5LFCfziVh1nG5RJuMBGgs4M0DeH1IYOnmiaGUSGmVc0gh
SDYMZ2EEG6eIN6NlUWzAKqkPILNyVhiJjakv/8BkExzgmi3TI9h/Ww/TKX4EzAOr
sFMaIrLz9wMCKRm1C1DLcg==
`protect END_PROTECTED
