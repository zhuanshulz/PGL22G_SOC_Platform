`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fXnqcWYlNuaZNaUWuNy2uzNjvNKNLLxNJ/cCg/qpGDvX5AtGSOilXegGN7KTpfj+
Hz3nU0QffsbtMhVGr7PfF2ixt1RYJ35unvTZOO91il5q3VoABtGlYtUTUUkV5ZEk
t6xnGFmn97L0e/koNKRRnk+kBSo8lAchG2qhLeKv/Vl4te8rWglDWqEz7cCtmuGg
XtzCyFCfi2wSuiWYB7gStNZ0koWW3NXnkaB9W5y+1mEEZn/8rxKUMmP9GobJ07wJ
ORNDRgIOHxOglOm2I2fMi9rOIoS7wW/Ci/ij3EzOc+agegEKiaUqqygzjI0EEiyx
e/sPfBxGCHZlu2CSyVSIByUhQHGY3lbJQgOpFsSxgjfKxDhgK7+0p9Le2VkQkk3o
dj1hH7iI+oAt2kdyuEypTouTXZkF4JmqwTMbMhy5t57MmHOOZOF1lbf12h+tt1it
`protect END_PROTECTED
