`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g3H6cU1o8a5jleq05tCC7ddS4Cx62qc5WW/lbikurkk0z/uqXRcEM+QXCGZ8S4mM
oTpLCin+XGjrQOm+9+nfMfWyq3tIxC6ER+MjZpPvuvaF0V7t6K1PC8A1D+KSM2wx
Cgdg7ist0+xs2cOgfc0oNwDxRm+J/1iT0zPyzSuqplmBhF5XEmrv7l0kI4HklIZr
T7dD2jU2Ngp93fCL9z57kK2IVV17HgflGFRez4hlrmYWKF4rAZyH1p3eZEv01ObQ
D7Q55VdyqeZNuKA3rzI3V/nQP3sMcB+Qa+ZrGAuuOKkDXhT/rFRudQN2zIO0WIIQ
z0CFxcs4yD2wp9tetQkboKjxroTN12zDi8CCXjM4LoMg4zVQkt3m6urEq25K+6UX
QXakMwSRliiOj3JW9vUO7cXnfD62e6VvPlXV+9ISYohT3RDTYc3IEfr85ft8Qkcb
WeN3k09jphQAzBthVynBvdYGcQKZurXhOj9EjJ1jnueVtgEijfQwg+4Bo6opMgww
Dg2VXaVGNQLrglC2ab6N7+c7RgMoAX+Q6ObJkNDGJWx1OTXAlO7m+4gQ/RXmPrD5
pvPATyQVmz/+jAoUk8tRsqcCYFx42iiKWvwiQGbJiw13AewWnLAZQeuEFfhFJ3g5
UNUu+KqitVSxnEIh9AfVlDdRJ7W29bE6wOzyfDLTz9bbDxOnpIv2Gd+WrVh7aros
UfXL22Cj7YjpgGU8HJKuOk5cdih/aqFYbP+bi4Mp+VNwjUKLOiAQ0ZWcTC+Fivdi
8jynlpxGDZlCAZP0BcNFDlowW7xhzZ+MU0y05mROZyVoTwxy8ROBT80EPGHWjQsO
aaMFbZQYI+yuwr463oQ7hrQsdMY40XzZkJrYXTOXYcdY/FmxYjwnbuvjRWTUn5vK
XgELUmn0vkmw0VSYOy+0ZvW5XVuA6P1Wln+ooEAnv3s3TbZoyrFML8Mtp10OmqDu
lxWtWhHHjZ94kXaBX928BFTaSevTQJxGXMSHuuI9fAAesj2ndGlGHAT8aJDBaB6l
D9MNSwJLVRNfAvA/pkQBHKJK6AqUclDn0SBpW5BoIV6R/iLIffCWDtWWrRpooQBn
`protect END_PROTECTED
