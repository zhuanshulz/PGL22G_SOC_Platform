`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
grbqvu3EizkT1bHjNnjuo8Emwi+GnPcqyVpu5/mQ+/hWmzIeNkCUb2q0bI8fcjvy
9+gmQ1bwpTIs0SpaRaNn1Uza0MnmghXuhAFOECCMa9qzAJWmaKqP8McJRhE/hBQ3
kmQ32778u0G8J3LDS/WtqQ8gql5mxD9KhYm2p/fQNtsjIKLdEiF7IBIutiF/rzls
H8EwqJAqlNiuXy0NkaWC+qdzSVMCgKxoGP96w4KBV9dQeqC9f6QkL6ZFH0HglBUV
DrmrF1uJoGzbFXEREdL/hJTbu2+hh+RK6z2xa5NgSXjlWW8p/veTnlox7v5frpi7
/6eVpy/q3Nuudeh4DC0+TDMqRK0ezRka8+NAMpoVgIATa6w7afK9q5/8sYv02IVN
nuymZBYdc2KUyztLhinHcKYgR+j66RtJJHgkK5QTtZ9Bo0Ma07Y/pwJiyEEvFq0W
`protect END_PROTECTED
