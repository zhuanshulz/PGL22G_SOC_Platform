`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0LhEmUJ0PZIWORUVXyZ1s+vyWQ/MEzfpyxhvMSS5o0jWrZgdEs3Faqor/QiTimFj
94vo+BObfbGietETPf6DzXj2B4/JF1YNJPoRFQ4edRTs2OmC1pOGOCvdgYL2Bz/B
HyRXpEupdoBJsWxfQj9bUW+QyDm5Tni7F/5FkFx9VWMjviIQ3fJp4csQI7xQkplx
gCw4IEYGrlNBKsdknFxDkfQ9MJ0VluHDbO48/hVEtxbvN493s1gLwNdPuuX6RAHm
ATfsAdKJ0cDUF9U4tTrOyqy8u+3cuN1BB8QJM+VTxFNygfArc34kUkM8wI/1HMe/
u0aKf7yBp5Vf57ohfKaNlS1H6JYF2NEzBlGI5Bxofivb/7UCsSz2ppDz85hUfiBz
4dAQlEAl3ze4OY9qK+stWvxm0wUOvJmTu/tCcT6HtqCRCVNMb98H0EbhcZoHFwcF
XYNZQAqB6lc3LPgpxOTB3ecxKKiJTijkqiSy0dfC4uJWUMj88VN3wXu+C/4OgqmV
0DnnSGb9Kete3G72w+wW3g==
`protect END_PROTECTED
